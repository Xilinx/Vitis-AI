/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1392096)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9ad926fczzm/hbnrwGYb+EK97y0ccPFTPGljyVVWZxDj/maCr1Xk5RyO
nUqpKjzuuNkqe1R4e17MzCOKx6dLb0jq477QVBNF7/YVToE8T983x9KUbuk/M2axt+JauJ0B2BGh
EECyJLH9DXKOturFVWlDxM30PGfnQ/zR5tzRcmkz8ve2QGF/XLA5+mTFCW74wXftqbMQLD8yooP1
SSdAhAfkAzsclhfVgy7GY+WFn8n7znLx9FjyAeEsbcV4isIoQkos61a3woSZRJpiuBOAT7NV1DTx
nGWzr9eqnPsYhqdKjJElCWUXn64UNRW/maV9waV0uYIp3kSFg8ULIY6v32x3UoVm98G/eOQdQDiq
vh7UeXG6Y8Z89yKZL3TVohSQ+ThgQ8YaJ6qYwrNsTIcnM54KHzbgRJgj/WxVXOyL4rySMhL2SL1s
Hpko7Emk5ir7rmrZxvG7+QQqLgy/wYMzz4n2c+slkHvwvOgtGYE497ZAx0nTdJDTPcA6G7gAtfDC
/3um1VL8xrsaAWp8taaD6wNS6UiZxC4EO8FzCvAH1wx6H+iIcWNpwDCx804nlZWEtJ975m+lxEF8
oU/DqAV5t1aX30A3GkOEe+VFaNgnioG9CbMXXMjyb8trTXZI+1qc3sKdFolT8AnZ6LypEodVkzgI
mkM4uYXBJUDGPLlW2ZA4PWiGtxnFAvv+vUJUYxBZ2q3ub6dAFN/zSLjeMzgrVNjW8piwoBTh9qDA
Cy1SKWERtMZhdR+Zco2LdIcjeS1UvQ4wRbxziDpVG9Ceb+yxQzDudaaIxtZN3UtOOnieUaN3wDjx
f9jkYctbCDIeyY8eWI/nSbKTenWUVtbUG0V/aPGYAw5+Ph2+rRUzbCXno8Ms+t6basyheDM1QRXH
hAdhvNmzYgG0F2/ctlmIALuaYnMaoSCAs9+D0CIAdaakiDcZ3EmD4FqRqqnuR3b0w4WAYssSd1zs
8n1fze80i3mmIydljUNNlT9sbe/ZoWM7WttQJaIcXhnhlh0JEOpssz3IJSqE+FzjLO0pQUAFzLxN
Qaf1VpPRv0vavWrxHX+v8UKHKLu9keJJGMXXnsKp+WpwRbend9ThA+6DKAirS4QVxBXx7Hi03uiM
jp+jkI/vVgSSv0F8NlbeKhHK3MrL97WJRqC9h1rlB864LC6pdRToZSUXBbFJndtvd1Oh7DBDzTkO
F+b3jVO/LlDFJ1Od1+9MlDUSsok8GipHiQ+E6+3BemurcfSq039tJ9Qmif4q9m0eb3aGVXRN+SQG
4HwFr0Qa5ERRUyc+ZCyKFba9RLCMIZ5u0wWnJH1HWoELssEJpIwXZl4/ryLsqdljKhZz/crJDQ/D
vvd627mkKs5opC+dTPTvO81ka6Hu8JR7gbvLaVunKw60eqXrxybsEfSxNgvFX8uEmm1U6jhkoKs4
sxNUhBCqlIOtgSqls21aqR8cc+xQn8P8aBp7Rx6bxTEjsOpUMs1a9lCv12OGN+pce2F37FIbp7Y6
z8zSLtmUs/RJqLL46CcLggA7ipvr2U0ZE4TXe4PHCRXALTrcffk3/0D4Y83R14HvBjDQkrtkHBnY
J8HbGK82ftIKNOh76uByhKHKceyTl6IcO1MIQPqHGDMhnzigESCu14rGXS2DfpnppnUDoNvxeRaW
NxamV0xfTU+4Zc7OertoTyyv1JmwmVloxtJJQhzcy0XWMz4tZNhkaHIMy5MC0uJfxge62YMIOYBr
9bauAq62QFKE4Z3cQsV/2X2x/N7tc9EzfVe5LfsO24wAKko9lpP5dXLw2ROeT7Sa/pLK+wxbzRiG
ZM6YJZYh4bfOcgmzeBBsx1tjSGsrlPMflrRFj3lGsN0YHIYwql7SzxR/WSLDQl/ARzJYb7+u/nWF
sY/JjNs/1tiHnHMhp6NdZKHg5IF4lQB1SZ2swhCJQlPv0mgQq9FqnKheMyeHFaiYwhcfEQLkfdSE
YS9y94ry5Gfc/+SzuYON3Lm1fY++hlhGeRtzeEozVHXIPEK5LC7fIjBA/3mWEqYJe7GCNwW7FfVa
HOS36lOUjnz6bkjPOxOmKWvUTUnIITLS2XyHaJ/CeGDtqZtoJV2hS3OGNAae74CqyDvcqbbY9whq
lsMIAUja/n3i1/cZY+wlT15TpPK3NTR08mLsgTRqWu9uwIYJxNPMOjwE0h95wom5LwwyfwIl+KX3
qXmjC8/JT0UIa46rOcsd/W8jbZsGZ5VwdJyB55LrKooOe8n9SIKIpHYepJACdrBelx1HMX8uuiB4
dzcyPp+X7b8Ez595w91ZlJzNfmWHyFGmwlso0IjzkhOXxb07RAueyYD6P7ciKUAMVe0UuSGaKbgU
D37h3CSR2PTYDFsoHFKlO2vWWgC7yrwz/i5IQw57cD7DedEonZYMA7C6c8+dEApTB7Ljju2Y17Hd
drZmTmOMTbsG9UYcYYbqwrNsPrusxgNSdwFs1227QYl1zyPH8CO1EApQEnaPJl4Ruafv7MWL0/5G
715J8Ay+ilSyJknrX0qtFX+bVxIRwXO28oYg9RgzSET0M6z9xq9CRfYZ0xrj4on7vbCphheJ/bVo
Eve/4oPT40QlOKR72qOHqohXfmG5VQnzzMjwlihtYbLUaeIkKCvV97oZML1THpLTvzm5bi1EbG0Q
+UvQtGkg34rWSQKyebjMK2HB1e/pJ+r3vh6EkbrT8i8fP/oF3NXB7KFeiQzRTLV6JB2bpgbicEGp
megs57phkseaOurycejLheRJ9AE2uFH0xWoSZsZavCpzKoJIwNmiGAIwGfqhm0an6wclSaKYgClC
v7Z/Q7w+jnBpX70/GyJIZa23slCyT/hwgqyU84NdlNm+7TIlijratv5P0rk5CIHrHzeppzCMPXQc
Xxy5PQ9LiXQpClncnjLYWLSXNSxxa7JNtpSNR4wn4PQr/AMypUT97eHgjNbdDZdWXr+1Z3U67E7B
SIGVYaLqis/0YJgLnt99EPsEXV+K9dxN8qsf0qekgQvWs8mycGL2qkUG1i2fbxc7px376OxbC3qx
5UClxBv8ksVNp+Y7DZSmpAYLyDAzRmaOOKrQOtonjzEzsOOcloJZml81IrcoWSf7JWQlw1ciCfzx
PTHyOrk4g3kyMxIqoUcZFSTymE3zrmVQYFszsKQpl36YzFkuNaTpq0AU14fQLc1lERktNrvVhRKJ
Z2dBllGCkxF7fKKMJQOjloeqbHw5bn4K0vtaD14drHG/6PqX669E4BlG18kT2O1rUdm1YQeJBil8
UgfKvl2t7hmxV8Jy3CdZzps0uQl5VzdAldbq0r3zyM9Y7VJgfuR64Qpnm+eoLBe1hNAk0gir5Huq
7qvZilDHtICC1qrrxIzKI5tWQRAmS/FDh9kcqoSVcEjT0lL/VgkFFMMfZkbi2fioRkNVEo0tdaZp
vp0JySJd7FnhQ/xdxJ3uzZLjRB/2aD4fiXLCUKOPhL1JIcKsRwJjt3mIq/TjP6XFy/9xhxeemxbk
+cU8NoPJMtikbG0SGevH4f+XWy9DdhHweli+aPr2NogMw0VV6JpcJGQJTSqnukrShQ7OzafSD2P5
I/8o8/AZkZnJIQ2lVIdNPmpmqJTkdPIbI6yd2NSkK9Haj1l9lCEHz1tFGJZT23CP0EMJfSDZJSR2
i8vmXGyu8xlAhgimopwK7fUND/YKuh/ee53zr++6AJoAR4vWISUyinnNPM221l6H+HPLou6OjQDf
K83lLA4rbMLbqaCagKz8jOY8KpYXhc9IyDI4DRFSJrHaJJ1L6IRNd1WDVFxBCwNGaHfdO3O74/Zv
fE1wZXYH+y06J5gvf9KcKJhyLgkX1dqdWxRE1E2d7EBoW5Vt0cM1CxutWfuOz46tuRNJlACS0Ylu
DgZgcRCnobTn/fp7Hw/CcTwk46Zc6K5Mq9UNeiO7n4LSC9e07hNvwynWUrQluY5sT1th/XK6iM6Y
N2SfYfleULJH4sKLizeadL48AOkMkv24K2XO/rB7qzwAh4Wyuyz7rZuIzLVy7oEnYGInpBJcG070
IlyOy8coMAT4nAYSOBhl77t4WiCmLMUukIhHo04T66FINa4tRfXgFK9JWIEDOEb9s65OOgyGj3HD
oqSyGM4rK16VzK3u9mJSoA/nKjqoVAFB1vSAlPkZOCsRdp3VVEGV6G9GU6efKY+wmvAaNi6mahvW
ThjJHYRyL+Q/OZ9E0fMSOb68GZN4b9iN/B+Nhtw+SQNCIQtFDgHbtmOGgPEMGX36NHaFc/gYdBwG
8BkugIfaKydeL5x87slYYOa8XunGm5aoGeEArF306gBCYrx820YWHWFnRFLExGekLAkrcO/n/YXs
d+crWsdbO6HTZm0QoarDR4fPxIy/I26QU3P4cTy/LhpnKkZe7nOxTSC6WnBCwUntXz8h369AxvK3
vOFzboBxOOMXf827T1b5p/MO/7YZ+3y2OBxUyWLLjF+9G5pWmZ6ATRngtS7q5vkhz57VxR5yiwV3
MieBHmgVrRJVliOkrZJ+vXbq0xB/KSFcHyCXl1wl1yNEe18F0Ze8zRRuvpk9org5xg58fuQu/skG
009vlp1xDwJVMDJeXd8jyUtJ7+vc1ZloPL9LI5T5R3wQ5lphbHv6am4NC+G0KIVFtIUyWezUymef
g5Kolhd046DianJ5WcSoWUyVF4sdsNiw1dWw80juas1zNCt9my5UEnJ/Bu9Xf+zbWMcT/cAPp2Nj
jawk9zUc63RKznyGC+9g8NIpEL4O43Mxm+GoWDZUf6TZSPvDN6FugcwZowXZurafRjZThrFJMBFw
DFu5VgivN5DpTcgs+6UpdxteJjY+xiy8SSA+monr0+JkUarrxcH2ajfy9ysCp16Da0I/8nfZF1dD
c3L+U81vj+ljqFjTL20u6fC4R6tpenuRJgHhEVjvS6KhmMESbDej7/Jmcr/H0VdtZnIKgGQyUnlx
CEVR28kBK41ROGptPZR+3bGPZV8owbVBmHGGfMchM5cwOEOG4Q+3/6z7kNTN4di2Vb1Sb9Xc9vZy
76qdqp+2p7mDPEEsGNfn5QaCcEUvQeh5uHAn06zxgvjDPLMKrXu9fasJdGmYDpvkKe30lX2i4AQN
SLIjDlnIXEr35GEo+4u1JFC8gJyR2s2kWXDaOR7vAQkR2mxfBUPZDo+N/a5rJmCSK0oSPakqpnzb
UsQsDMvkmm8zQvqUbrjQf/SfpsFVEyyvbDAjyOrntn8KFT1gjipBZE3xS4WXh8eMmH/OjEuh4wo0
paJCaH88xakllEHzl1xjd0RlQWx1wuvW6rll/tJVsDmEQl5K2/JYk9E8H46QB4hHg0/wNyHiUpbS
7+42RflFmPtB3YrzBe4BrQNPeoIYeLmGBcrEefnFB6oXOv37ROIkP6p1cRJHysRZkNiAVrD3Uiqn
ggJu3f/WAEKmlQYtUemciIu4OkZctUfaBqZOUigI8p04S2ZPdckVwNei6NXUYqApG+DzYYRLUAoT
p9KZpMDtEZMddjRRIO+mptVtTp5+pgcE1IRe2mRGrE/9sDgbV0Fvj9VASpfaH2KLJILIVtkdf8m5
YHORRuy+2JoQdQou+qH56KlE4m+p7tvg4/0A281QTNqXBktX3o3byaxLF3jOAK0s3UsxNU1EwjCe
EqAtxxe05mghdsmAdKr/J3RM7gNjCBtgE8UvFDWufWjykrLgarWppFZu0R3fN58tb5ExkgfC8yvs
noLTA7ZiNSC86QRQCNPjfaHS8mhWfcC2S+8T3ai63vS7oIvjaOp0soiKx9FlWELPuWSleZm8B0Md
179Wy0JgNjFX1AqfZgg8ghau4ytplTGlJM7sgmNysJwmn6o/Hbl5x8apSesfjbQSim3UhKcJUS9A
SVeUygvC6F87nW7YdBax4Mjh4zaaoLo8bEnNYjl5jk3T1PvSqa+NdHdxrTcnZnMZr/TtzsD4omd1
g3ugFksYTXzlGh71Z6tVrNlsmcp2QxB4gqXbcf8uKL+ZtvvRlzNoWfr/NW/8/UAjHIvbPZwnon3S
8HIOYLUdQ4LCA2t6eAyDcR6/tdnfi3Im+URa7Rd3KOdRm/IaFObm8ijZh2BLkmdnkMO9hPhz2uiV
6HRNgksYZXspDsSOu+6vyC2T5oMJf5ZB/Lz8U89pi4BaMg9tNKdx2zZYt/B9Z+C23R0GgUhldDKa
Sve8TD4Kny+SPN4DmsVZVYAWsGLOwEzdZvoUNvYdXPfXlpNNTQSYFQXGuJvOlwGy/t2s4JNvbbQY
+ubllLjPZLrUvEWhISOZX6uM6R2VioUngBOYj4aLsXodItfRuyA6NmRsStTS+GgYWjCM9oLtSQ0h
EG7GvK45On18HZD5mo9qEWS/H6I+OS4//eCL3EZFByguF9qomKCxWvk3/67s58m8qIWFVTVrXtq+
yxM88DX00cTVfX6oF7z3kbP64wlyFk/e82W8rOJX6qNUIKT3Ybvy34+MPpqvx3j6uNDw79OnLSWT
0dIWS4iNsn0RaSFRCWMjzK3jiQLdJmBm47CUa6RbF1POc0YBdbNsi76tn96/eE9aS5smzOd99hFq
qXH6PE/vsFroXKCYP0276lrYMC11kxQI3fcxGFQH5KfaheyOPn2uWF2kl3s7q2kA5mtI8IngEuj8
fqQKFlwH5StboAFnJmjG2feBN0oQvFfUrxcDO3B1sAyr+WGNRCrwhqyuJDyWlymp9QACOGys9Am+
toWCRPrjSpVm/gWEXZi9jQuCUk9J1mymQMRWjc0MRtdrRa7H/1Si6lAiliERidDGv5YfgwL6OON9
iiB/ImQa1UWohIgDEtw/fvpCXcR7G8KqSSFhLqUwLBKCjpdW8yFzD6t+CfpGrdBp6/obxpoetVLA
ow0VMq1pGCOBO5HvWkw/iK/KBsnEPuezwGEAsbpmsr6Oklax15F34vkQ7QEze5kk2ZzUA0/YKMb+
iFRiT3xJTa+KUA/oRfaPP2YuXGwKfxjPqWc5bHAcBuJvLK7gPfi0laOieeCw3c8BbsO1CU2zBJWW
ZQwyr2UFhf4CpVe/qbfxDQbyB0wYWYjqa3AwcYw30PdxkytwUcnqjuUYRyumXR94/IPDGJphnV9n
bqnbvLoi0hCfSqm3kTqCLA9dkKSIYLg/MevQOSjjcj8BW0YadbTl0gFPUj4//3ubrF9+GOlPpo5J
IFmD3a3NBFDT7d1w3PbCGvgTu4Io3vJ3OvTIN+/b4PRtkPI3g8SUZdZgC2H279SkIc4NTqQ/5Xlm
b+mP0SElEBwcMu/PN+D/+BFgG+Q9R6vp9ND0bk/hdg4tLC7SZFUJKqNolIyI2sKmrYDpQTxUdpPl
18Cqicja+Xm2VXym9LTXqyMUQ1fU5Q5RwH5sUKqKYxk65zLdzlTVbi9n8f3f5B3WovC3UIRuUmZr
T56XMq4UWbhNoSFBiAtgKpumwiKlTvlwXtIQBnAIlC3/BxzYBW/eFBrVE+Bfe3LSAQFG+mzJfkE5
L42gadbLzPvM0dcMZg5yVkpinxxsQBlMe4ejipP5YcBQf/XTDf+dZyL7PhZrZ5ZwpIXByFKs5Aj6
CcVAZHpIRew4A7VZg/5LL12YYGAdDjLjMEuas5BOYdkCkTuXngyJlf7jlO2tsS4qkbFDpFVX/Xa2
h15GbX5CQ0a/OvbuXzESaj8eoiLDm85ed5iD5Z9uedc9/tegxZPp+p10Sf7tizuF532JKtJKLZg+
lUDxfeqNgENsgGuRAKknZ4n7f5Gi7ltoxy5pzppehyycMiClnhOwbrp3ZmUcBI8zCSjDlXrtDJD0
oOrGsV1ySw4ChdhiUt8BmYRXAogFrG8rqEcicrl1wYFW0WOgP5SUsBZr4m9rxW8Cps0cdRu3fieq
Ak1SYWqowcHR/oybhc9HR89sV+aTQQIi7h3qzESO3pYUPENdt4nz2dt0aRtNwPz8rWh2hviDOZbx
LpOSh8b0R7NkaoSPDkHi3M+qzKRXO1l9atWDlMe4CbKOwZY1aojbJtrpSS/qpIpEvc9otpguQhhB
zsOSiWHWjtEZGG3jYjuZ+ZpFKKBzwQ0RTyjlc2f3J4lP1DbxNEwEZD6UYlI/2w+08BpKY0Eo2EZ/
DSrYarNkF3k4aTvwSf3ZNRzCBAomea721CUkVq9rNuKqJ78FG9H3Se1V5JTKPMpfLuVbdWPWaFDp
OFjgrovf8u00uka0XEslEgXx/HUrVpleNrk80QavGyE0QYtBfC3BEajM6t2PIAMuD6dZfVYyjtmC
l/Yk7pII/TS7RjVfq6ckUo4uGd4OJmG4rHyuHMiE3cxQqAnw0LOomxp+aB9CKVlOrNWVg4zjyGlx
IR0j0D5HtIv+qPG5l0Qle4hCEzYZZxOcZIkNysTfU0zI8lMcGcoU13DiqnwVubm/3byoNnhH17rX
Ah1Zk9uIwjpHpQYjE0qyC7nqHuzkoyMJHX41E7/bzNlTK/JErXA+SBjz7tG234Rmi9NhT5h2UD08
ad9o1jhOA5JssgO5unGkZSN0wlgeOqxfkK4o9ikipLFxCTSnILNwrJpxNrodGz7u6kMPov1cAU0O
8ziebG1JwXWPpqcmEyGjNlIsXLscdyCXPmuT3rUYD6u1n4D7onxrIIBS2xF4CxkALiGTLGQFo45r
/oFuJ4cEeELIzdYlW7M+VA1I8Fc93Hax/8sh/kKiRBmLf05yz65qzinYqOp3KODQeOKxDT5/ulcl
fhYSvkPYoUmYf0fVJeYjvc2TS/ZM6o5+yptTUUmCRDsfEBWgYLjfB/yyKDT77fLwhUYZ+zZ3mYhS
Ger4BG0MmNx6gXLms3wKocxTwnePCfhVzO7UgaIYiJ556vfHJCgNEKTV7IbNMCYGKgBNE/95FUf8
ikpbA4KPkCttGD5lO0kQOKS2In6i16p447ciUYpkb3WlLbjLiaPuIfGmmqmsEw1Vh7Pm98f6dwJZ
2lFoAuOc8lqfP4H1khc9BclmacKOjuCebBcGCcmIz8UF3CRAuwHT16lNSU4NkwK1ojm81fBwq5a4
YvNp8DLkrQHNFTauOwggZ+kMBDi7qFn2PQ1MffpUc3qvqIiaJeHQjn4vK/j5wxZvgjUomHO4w4BD
KEeyQEtNgDCH8JP4YcMNQ7E9P9y00CdXUsX7My0R5A5H/Sxvnvo1BE8EheNpWXSPAUUAOzuAcFff
8V46QbReO7iN5YtFpT+bdVCnm7Xr4GQEjbFDvOfHZRKgmb+uB/NR+MA7fhogxRyQTQbY5u5QlbKa
IVMK58rBktVHiJx4WvnUQa7avs40sEkyNNl4o9RTLRjGtiU8EEPoGGRWQfQKrlTAgWL7z9J5UuHT
xSukQCzMzOAfNq+m5yNx9FrGGBeNrRDhFQV9R8m8G2Q/Haue2S7YhVHKokrMLOCHUHKsp6MBU1Z9
fDnTAolFp/DSe18IyOMopY4OzE9WJvH20R7/RIhQOx3ZHUaTCW7BKgwA14obz7+QUBT2qMUxcDUu
n2WC7rkKdr8ciP4y34wLPUqp+7sOG/AboPyADq5c17pUUd8f8RzQ6YoB1C+1GIta5Yuos3VAoaf2
2vAhk9re7liW6Bh8Dl/Zwcd1WVzDy3Xfi09WCGfqMxSbttXwwVKZXxYvhxkA2cOaSYs4AqGyYTZy
Su5fSuBQhznosiuNHAGFrBJGxv94EmqUBIB4eIMqFIzddJoxCBy/dqcdy0KHCGYXWLCPhKuw/54X
10IQmyndIc2RFHDiYNIA5JjI0ooXBvs1MloAy3akGcJj7DwA3ExgvZvVC7yrfF4cW7/uLHWpCgfI
WaY65MGH33TvDEkzhaIY4qr+Rp8tOhXbdIz0z7DUyRaEVlxa2GOR4LwDa4/z0cIHljO1T0uZh7Kx
A+tfQnikVQXjlcv2tUOTiePDLQXl12eahuc9X2ZzJJ2exN6a+jmtGD5t30b0CXNxDRyyscX15/qr
ePQRYJ5uOFRxbylVGSNeKD05aIPkBbZoeS2omewmW3FReLEA0MDRLmApI95r7UkU4PLx16sPWt5+
RyT26svqsM5CYS8LaA1u2lXnC+QCYggadfqwzO4REMjlj7PtRdiWCRNq0JqE2UCwUoZ9v7FQk9aT
7N5fjh5ZSdqT9ipVS52FzCnEnMPo8vj+rzkXVaojv1MHDiIfwIav4UyJdUdEwnhpYTqId3d5uLmO
a5rYw7Ak7I5d5eJCaAwfQNYuTsZs+VcOqezbBOD1zNgdcnqI3zFuvHJ9Y+9WbDNg3Pw/BDQ7ZXt4
SyjImYPILQajtewoIgqih5YpBsfIWqQjlhUdbFD3cqSPWNMrCZ3r7JMp1aXJjc6SS1ALQ9mqvZ75
rfva8mDpQ8RjbJtXBlISP4JTcMSNPlfU71JZIBa+pP+YxdoBeTp49vGHcMxB3ni0c90U7nRW/pqn
uNouPKoyOljmlF1iKN85yoIE+qjfVX52zrQsdbtLkmcNxMummVYtlk0cRXJ+Mx7ozJH/MUzuXcB3
2cEyzXV5qHbkpJuV0eOHKQI526z7jPF/YtgYc7yN2F4rYo3Wn4LIH3Kb/imww1FReFiTqZTMULXI
P9WIp09YSk+XZPNyQLxlglQA84s02e1OAYu86w17kw8YsoO54zOU1jBl2ItWDWX9mIpC6GmpdcwR
7yXmbZXkQKW0HhKNPY178EMJtW0XKfRbudGJdPTU7y5/aW4+OKrIdA1HnUeQcECejphks/0B49OD
UROeO7vKrQh7B9mrD8tDmcR94HcGnQ0rVUfo6OleAZwcitL3GpZV+NpfkFB+5Wjhe3aI8b2+PIp3
GDf4xNdwwInEY92iL+mU+VdZa5zJZbhCZizxCbLmem6MY3HfnIv/KiGTG+LPgjdWBRKviDndV6U9
W1fk0ghvSDqLXNjo2X0+HWOCxjNytTmBA9ElBYrWx//yWC15ALHbqOJSK8vjrlcBdRb+1zYysxcz
gJtjzM8uLerxe6WihLSOa2RD01J/cVSGqdECsDhRRoX671kO6vH7BS91FaL9vj4ilKCAVQCR5Cvc
7gquuYVqfHo4ti5gohGEDgY083u1qNKdxjmxH/38RgYcfN8JwRNmTD0qqHn1bcleU9NBYyj5tOIm
dvi72JTXAyuMX6hDoKmbb9MRICGN1LLhxM8bzo61Vk5ZmK7jsLyzID6eMkyzl83dpTpQGBvJOW4/
1c0SkGoCM/cX+cjm+8EsBu7U1w3ZhH8oueKV0mcwlrwr0OHWmMbL/25Alm+9vFaI8Q16tbvmPgM7
0kzFdBeeOuG1+zP9+tdiilAnGh528ETOeXsZtI3cY1PA0u5q8lwNE1Ojbmh/hOPsTDv53XuPIeTm
YZIGllawaUaTS5H60jAOeKscU+bfAM2VVtCswIos1TLnnEmIelhT5A3sqMbxM0b2tMLA3UDnRj2b
3G/lVuor7iVtMVeQNU3/BfZBCNwZGMcVf7aR5kR2rnIG+wDC1ji2w6har49Ci1S5V4UceSgSXtgY
CUg530FmXcJSfrGWimTjQUGTLdCjP1Dsqn18NKv10oOu8xZADeUd4IjAIuXSmQCbvDFXLCfbg/zX
rFdtPRSIe0qN3LPqSdwtXe1xO+RjcjQXiL4wT+HBfiixEWRi1EQwjiZULcQw39hNUdYINaQ3pktS
JyBHOvkWPBWXNTc86kI4HTMdm9ADEPjtFqeTMYUYG6STzYWBKcGHZYHyVaO1euU/62VsZ8Wssi5X
zXqH1dLtLK2buVwRmpHGSi5gKcuy9RqR1/y9uHkQ+njS9HUsEx3rmY8/eP7zaJkMC6C37JNwigV1
bQf9vGZyFCMGLamm4dG689Aa7aPbO3pFIKonO+4HH7v7mSlsL/2wqNF5Tn1jIXEZXg2V6saI2Lfg
W+RW2TVWQDWHlOONsF5KZguPxHOOOHhQkElQSCYC8Db4UuZo+cnSr9k/wKox6z2PKvtH11xmFTF/
wMPbx9sQWdn/rSmlo6NCqlMA5ciNZOqh+1S5XgTQ4uqS4/hNTdRs9nrpXD+BDy2VrcPceLUf1EnO
utxYD9drd3eVmuSnQrDfgtLnmIUAZ1cKeXdo9I/XYzGgGSad34/KsbLgel7Vg7ljIrFVwZd03xK0
y4dXcq+u/7wz9MF/zM0ocCOvAQhd2je0g5fZn8aoAmM7FZj/4+viMPpxD5eQb0w3gqHGYKFm+nth
V2JSWn5c3ecIYB6d0J99ISCjHLZ/0TJNh4ejvEIxBC5mV+P/rl/chW2XY9IhRP+W08JP3NiKwg12
VJyiDTAmqZHYa68i1k2Ws7Sm+p+SGHvFPNaueIUpWYM+oZtyNQ1BRQCv9DxXSb4WTCQa9x37JInp
c1X5WQvGjxtqCL1xIg31TcGYO/Ke9QJsHYGJKyyBTIe4YO1hPGiTKL1tmZ7iY8WDVOoUHI/yzcnw
6Hvu6DK37gS6Ypg85QDYE6cHBtmVCxiCLHikcmalFL1kFOTvdNUOxfGsSLZ6u0vohu6+S5HdNDUV
NxogBQ/7IRbCUXRuY2ZEQ5Ayux9wPQASmv5AtCyU/unlMJXmn/SYtXA3zROA2jpcCQ46S7jsmYfX
c56TSxNdr/JikSfKD6FNwX+tnEB7MctmNZObX6hw+4bxZvIVcg/2Yfm1GkgA/YUGIgZCbskQUMAg
LtHEOFPPgOivKcIW+KszzFx1LxM9GWOdeXawm8xKYJE+wW3eIec3T99vUwV4Ho0+K47Vz6eK8sUn
NnW4nA+XIfZ59uV4yqr+Yhy3UykVZlLUVNDPmdaannCBCfY+B74wq01OL/cyb1b/fict99DMSWu1
qVH4gZtfCvLgaRb0JjFmJbNHzaXg8tIEcpt402GU4Zl74pnrTnsRAGdIyJO6hqJg6dhSgA4OXQR7
NPr4U85sBAKjOclfzIQKel3TRdfQae79dqr6c8yV+r9F56KDjZojVBr+9crrvs4iiQaw8AhQQ2WW
90H8I/35xzmuD7pMJatO9WgMd797bxlA+Sjou2kKIRyywrTza2+EL6IfG2ZURrB0sFCj1HCmEfXK
tiiNDAboY5XQryD0IdFhWBJ1c1oSG/iARsapSfmEcsCgPVXqyn6GCx8dqCCGo43DF4BbJuKiZ+BN
32az0PeUX3NFrR00N9TiyFR9ntlZL9gfTkyxsD/8Hi2RRUFyoiOUYtu3/Q+bw9F5ga6fP37kNaI8
+mUtZF/bj8a1CKIaxNcm19t7INlN/enL9/JKn8tW0Fp1EnX5+nwTJ2wV6XEaXt2029DC1hlRXqju
31+3jcRjlD+LprOJMpJ+3wWpNLft6En1yykM4Dy35CxkBQOT02hQnmW51FfkW4EzPQqj+ugXder3
cMkFU3FTJcJu+cj29ZYfVSAeZFtPksHNvDH2M1KcHSDioYVQ3MZEKg4Rq+nHgqynJq8LPfVlC2gM
HwTCBSv0lrvt3O16X3nivBwW9vAF3pghxFGwCl/F6Y6GJFlZj9hcVbCNUzRc4ILEaiLLecJuIt0v
9CvzEWonVe9xHECzDmNHSgqUY773fnKI4A5S7TQ9m9IdPyul8aT6xzORMQzBvScL9OakXo2mSxna
047dXPGRwX3c30fcamY99duNxKUsxV24XRaY9dqBtenU3IXMwDXv5RxE+IjMST5bf2MZOB4Bilzq
Bby/KUKyV9yBYeR25ZR3Ch6DmxUACGITTxHQ3FTtonwVJkDi/NWyn4gfSnrcPHYx75DZwqNq1acG
Vb3ZowWTna/rvGW82epiBwU8Y2ps/OqZTGDx2idRIhX9QU8swm8QceqS0vzZQb1X1Ufqg3y0qq6w
LiIojMq3f1ftkyzku/LvhwgWpCe98gWWZ69L1rKeqoa9z7jp456i8esWaUHUpF4FoA8B3fE/F9/F
tI+cM5EiUzRXsoCeYf7V4UupN8UvXQrBnjWOgAxCY6Q3y6SV2eNAzY17nHYfFJ/omPEnJF8zU3/z
/GzWSKlyh5fCx/4e67wInSXMJCUuuTum14ardg+/C/mD0xp+zXB/KbRt9DNYGbqfX19lGnWJykOR
1p6ZZWYtsfR9nJxCbhbQQ9LUnVKyU2CbI3hny4LluG1fNUjz4LWmx1ooGsQvouISVK1OQuwJm04X
s2c11eMQnfYRRkCn7Jfeq5Ixme43RcMbDlbQv07lRkOVGO6krS/CUBgwl2lfaAAvVJnF9a0D7/Ac
yRX+PDSLguE/Qj0HaKWDmQHqDC+bwoPNUJQn911I1WI94BJDapl+tAKlZBeTzZzmhYaw9FGdPomg
4tdUJn6NRwDNuHUBK1qTwB4Y5Z9gLRvuWCzxUPbDO2ZHbGxbTc/5PfoX11jFhxQLD45EytRpJbcE
j3aO8Z6B2G38JKNxYVn5r7xQgN58Cby4Ik90CacvpaiYgv5wAUgjXPg+95HnHrxyMXjMpgtBW34U
p9lNNhQB8ABMHsY0XB+ILCT1kelbVaILSvMrvCmLqEZGuqTN8xPpQq7HX1y57TW3yE32QKTxDkY0
bbYMOEfECApq7CBK6xtlYqVtFOiDj7PvM/nq4Nsr0XvRmt6f7IYZ92eH8R2JIqZFlzGCWK3BJ0/A
G2MeqfkK7LyVe8Vb1jk8gvUpDx/QGJ1Mrm19g2GklQNsF9ooIacxpFH+6q3TaVyWchwBsSiOIW8z
GcE+No/9I0PA0Q9LVix1mDK18uhjOREGUr4RcWtDRkjMrztw+dHlcxl8k4ALlWYPjqK6AhEx3mBc
0ntl5Bvj8ikc0NNmgeHVEnYs06b0XbZXukkiTNy+Pmi600CGfN7GxV/o/BJchlvzvKSl1zOGMMdm
80/9haSncesgMY0jrKMvyltNKHU7HmPQoRq/XzGbA4Bccl+gzFKQZKgZQwhpUHDAecl8ASQJWO7k
eZ6l9OVBy3VZvMNtXadk2wOWRBnI82P58T1HJYCxLs27olaFvUiyWY1A+JiVHh/gr03Ek6NtunVx
c0aS4lT954dwrqiwIqt6lZAmIdJ1c3Hfvw94wmqycMV+KnjK6UPMb28MuxuGNy/ySWn+lQF3ZBSC
liGJ5R41LrQBmmfnagrtqVARXS9YpdxA50isCDXO3GS2m6xjph++iojw566l47V+lcEqk5qpn57l
XZglx0SKsK8D6jMD4AFodj+AM0dWrFPap3MtarQxq8I69Kw3S62tVq0HmKItIkxq8aFVEFXz0JiL
9Kh24E9xlKlQvQhWHtyeaCUEiRIYJKxhQq5mPLNc5Rz5sVCtcWS8C+jWRa7XUKJuHUWSNfLDOyqn
hiABbnJZq+CpdZLjMWg7cG1fxWXcHPNfGH/FN1DnH24AVwNpXj/vkTR/bGIXtaEh69AQPQZNbtZH
UOO6IJBfNG0nPjDY8xP4rI/+8ZFHFVUlvtJEb/Uhp7gXMZPU8FCDwY6mwTSH4zxjKE6rBmB1d9+X
HLJ6Ha2TJOgckRwNGfhNTQYBZYyX3KqE0ZyoAyJM0zQyHNCQea5yWssw2puk1LlChtfEqLAT/EqX
8wgVzrSCyOhdxQKeBGyvRHKPNlpyUzFyrbGdfhUwNuUvnJB8O7+TOhEaF7UPw2PKQ4M9SpRa/wQZ
uSYb7jHUqfRNHWnRnVUaYwao03rF9r6+9mJVHMxt/X0QTA1tnJG6rez54USE+CCorI2oDlbOrinW
gqANlFmq143/wSOOKDrwZ80QY5oMlSMwaKvWQbgkWZYtJebaVCJSoa2h0b0aYGxpZNdOv1je3oWf
FkC1pOr+gj9+nlKVbgufiWUf4JBNDV6OxLkF+uCleaARr4TgIg8j2hd6jIXMT46MBn4GKjJJH7Qn
WUkcj6V9CjVM09Emd6qJ1kfBdPF9XglG9W7v7rAdbDkiE75MG1z37hMpWxE8Zf04Q/AgEHFVdIak
e/LD9Zn1sADzHMJmhTLdDFtjOcFd2LUIPXNxGe97U/V7tq0K70/jE1MniGf0gkTVo0vPrOywD0aW
Su+I58ss2Dj1J60cLR3611VWVYVY3g1hdzwFFx6ikMSlUNeAvKTbzfTNcjvyapKEvXE4RYb8Pyfe
oJsz4MM6oWYm/o9iaN5wOv7daUDefguyUV5S6xTVO/RD7oW3ojEwuuPn9har0577/MPMywPm+GDI
mu/WFG6WQF6tBUo4fStIF2Qs77AvT6LGnkr2sozdbj7LaAjJf+wLPNpa/zo7UHQhBDdl03ynT57E
UnussSLJOkiHy/T0nMzpQD3Mbysz1oah0Z+7SWtuYI3LMTjnAHw7trPYGIJBexVPYQlEANC4zNl1
4OHoxFruBnpZzDeOWwShXm9JipfKgxObWOoyee+daYDAKGDyxN0Xc4P9JlPQM7g8GKuFH5kpHo/o
o85kUfjhaHUtpJ+HrtP0yVq1k4hcxb/kLnPG4A2x5U546rCjAjDmxP8/DKE2mtGaArUEhPuJ1TIw
jHbjhWnDj8VZcY3wM5ndL1Kz67hBrxMsMvg3X1xv4B3AnIMm3ufW6jah4GC+SNL7PWnsAjsOYsvs
VQj+yG7+KWvvMUCfQFTkfvKykakM8I1fb/yATqS5gLBQQT7Nb5YbFOnMY7YeZYonrYFKAMhXAfz9
hH22Q9M790BdT3MkoZwR6ibZvaG9BqIFCj498gXwrE+FOTg6nf2RHlsq16uVLYodxMZy+cOcvRIo
YRBgeGAYlErBYad3HT+QbK1icf/SgSPwRVk653V8ZJzvm1i47ITlkrik2jo0hZQ4e9w21xzwJwB/
46A+fccHbS5ghh1IQ7LdbMeF/SBB7MwuyGFvjaUUzhlGMlgs9t11hIrUhgUVmG3yRgy08N4jTn9P
OHGzi1vyqMIAe3Fex8CS5ZNK07xWxBXWaP3Txd45qQb+Hf8hX+TH6W4KAJ7BosQIP7tIwLbUQr4O
GLcLcmglmeLixNrpJxkPYDssOpfiJ467LZfl7Cc51nT/VVpYXoEpvHzxEPYJnJ0R8du1lUwKKqzd
6yD6rntFBA9ji+Fz+S5SIuR96zkQwun81lmJ/J9ktQ3vWsN/P4iSMCsJYo2nCKVLOYpcQjlxCR3o
K6Oc4rg9ipk1zKMtgwpl5Z/0lRmet/V6P5RGP/gDmbv2unU4+RRFwMnYUZF1oUw+ah9jyBaGmgCO
5TP0CuMqj9wRe3BVUBJMYNiedUaEmr/Xp5MIn8kmF+V9L4Q1oLs5NDeJKQGKIvQUFuNbIxkXgL5B
/EUhqmtfcROKhZ9KOMPj9+QsVrB10P8k7MXdhRjc6vEUSXkQTab2SZuPgcKwvYWUJ4yLCyrrTjPd
L+EHuxoxKpo0Q1u23nlLk1QReuD7smWo6A2MHJ0A3ui2pkuZ5OUYyhq2K0DlGb9OCVmv1zRXsCgy
ehkE/fFSRQF8/kPI1aJ5wUs0QiDIh8KYH7+Dco7PoTDZL9LWmg2lg12+qgHcv3O0q1MD89z+e9Tb
TBWyuuqo3i4U0kPljvg1ihjY+rdV3hZsXhmurT2kJJNVBgxrF1qw5Db6Sevh3QnRbuqzcL/4nEOP
8vw44QyaieReqsqg9iFjtsJ9h1KBqXfs+d0L225pzGenBes1sgZ7ULzfCGc0POwdHmtfkLIxoE+9
cDFbvvSABwZIGpRJ4W1+Ox5tYB0TZHYSBUar7xzNkprXBhEkSJYcRp1QUAExsfWRz+z0dGAF4Qib
XF4aVw/0MRA+vVioN13RrU2pWiyba3h4Bx+A/cyvAt9r+NlQ2uCo7w+8vJ/ORbis0n79+QliptEg
3PJ3PRxl0IJft41OiDPWSeBB5ICgKbgcnGmTqaGXI/cWPsaN07MyOf0bQ7Oznnzjn/8yFuYwFAmf
vGMGpktHMgX9bcpYg+daTdILDjTkH+pZgOuuk8K99MAh79XD34KsjaNbkLUmLvo5k44virE4/nk+
+V+Xr+Dpd7EJNoRkCQJJy14eLjFXVkONbXV05w/0iqdXtRL92CyBk0M/IXgcf0fE7qHIUOPA0ejV
9VjjeHuI7j3c3tT6N1vEIr94BOSfXsszlLmcHX42y9y0Z8FMSdvYDE6VxBf1CfYYMA4DVaspPYDA
uCJ1S038rw49amk9m1NrT+zFkTEknFEvRLTsbnwQGMQtBlzlqcLkxSWvlOR6MeRHjS566crC167+
x9gnfVpi6LMtYOrHr3DZu3lzNx4ukEjL5+bd68/yUQMCQs7bVLxv38xvmwkB5uydUzXpSRnTXWqI
svzc6Nk6/qSEtO+NjyQjZkJGKqYDDtYnDV2/MEqVMdADJqMtXFQSOk2dxCCb5BciJvXNk1sUW/c+
Rm8c9ftycOYiIYEr6jPWcSgLUGxf2MkMuuo4aKAtcn73Gapi3O4EkT9JUtrjPC7+fRJUnkC/RLo8
D3ja88JpZXapISdTLq+p3mMbw5ZHrCw7gPaHIe4bsC+E2aS6VqV/ZRPXnrsMRBx4opCfrIihE/mO
MlYJHLPs9HvgUhcDhAKIJcOJ4hbELzVQzlx+IRUFyweCCOgrq0lXy+yhavqjZKib+u7qfKbVkJXL
ee2tKerOz6H2vhwaQRSstqppKMn8WxpPMkcFZd7Ei+/Mps4BEhJpUpWMjbUpFBluNphkJRUY+7Vz
WCXlr5S1Hwce9hMNcgOpFxU0Ma2KfcZ7UGBe341/IA1GGGnKnlja95NtGEQqliHyKfC9Q56LlTlU
KyDZ0uWN6TgwX05CYymoXhMHTIbnqtOJ73uCZtlrMiM2BwzqWT8As0t82t39T0uCU4YTz6djYGq2
2gVCZ3ACUVC5IpR9IS4qOkVak7wgTi4Ye5nMGVdBFy0N/WEkaY2c0hDvUYpVtGFwYoNjbfYfQ8dP
XtFkhBwftHMKhMbzCq6dTcKyJ4Yl0oTbMVOsNBS50QYCu087JDt3X3O0mRsz9OR+msB2uafzdcIV
/bocXfn300iZSiHiWgD4UkfSvGwrHw9bsHXtj42geg2pLsUcVnmP1fNJfVHbivXPXDIn8LhdIcP/
LpVSfh2eA/Lr5CuWwatR4quY26uxqlaaKQFUaOoVq6v1shA5lBfMIoFB+BaN1ezVSnQfcM18GkL7
apTljU187BARBNa5bVuLyRAbOazo6xRoRJZk21EgjStxisQwzbZIeumcmNRFBDtZXR9puKDNaekg
6nSKji/PLgcPQnZ9Zedsp6LQEGX2+AAnUUa2+2NbEIgPVRiWtSJnDYCBsSTxoiZowBQXGgn5bC36
PIF+b3e+k2XpvLU8tIRvWrFpgW0jZ5/VfsZjS0Xkn0bpMFoeKJ79VHuN7CWdqCvVBZimimzTUhxQ
7hsp06vv7onUr4wMjX7TwpqjVVMDTmWF40vyq++nbogsltgn+FXuIFB1ORQJd2aY9PfbXDgrC+up
v6nuzljsEXq3exIALU1mxfw8MK/TMKX37yRXwVsUFWvJgKZ/Y/juYtDhQeQl3+xFAA1JuWCJkK12
PVI6kfxtFw2fJ0YCKKrjO/EmKdJqs6bFQZy0fqMzoiqymyAq7FBNHDmMJ4odddo3L9Ql2dN+llis
J15DcgJ4wuGSQIBlzI7mC/4uMp7u7xsqXpJ0ivTrr/xoeazAMu12bFZlOONOe2l8c9aCXbU6B/KG
rbvDWMYXxvGx6aQi0o+cMpiQNIVZFgYr4VtJlOcKV1P7hLnox5/pDXu73STWFBC4owT7V9GV583Y
Kg2qKaqTcxC+4nZ2+IC7PMXc+ArL9ueZXNDh6BXlU+t5XzmBgQXV6tSd5A4NPocC0qVDQsjiUKxh
OdUzBg3hmTyrji+oQHHfnQ7o3pnn3Y4snemU3W82dnN1DFas1rnQpQu3Dy94h9rboofrpAn/qDz6
/ZJplnUZVSlIIec3yqu7uty5wQfD4UPl/7t58MtzqyxnUGjVe74HU3UEeAAZNqdK+ytYrMtww/Jg
PvrPDsPD4plkH52xUD6hpxWlLUwDoEmhFcevTzv4TeRmBJfhX/WUnb2lGeuS+bKBiY4UMuGaBxHu
YwyJzmpYa/2xVPlPPFOdtF2N0RQtsuCWNaFLRf95u2BrIM5eAv6NojmP2h2boT7QXAlEDWuZ0e8F
u62DRROEwk1L4ihhS9+tWkh8IeQfUJRwVXbXNthWu/jrCaVIIugsBaukcNszUc8JbFydLy1pP7z8
JI4r8ljTNRecxTMCADo/AtEneEWQ5Qumb8E+ilFKE4qMlPBKVg1ifNKtuEPpeBJfXq70cH+GQpKY
D4gG8ie4e4jjmjh8WFhLuvhr6OnGSZqs8nmNQxJYfVYAp1B8DebBBYv5+BdK2ELwTw6kwumH7AAS
L2JMf99/MgnGCLwiHsQcwcWYKwgmKuGA8InYcwGxrVFFAmU0LVsRaJREk+Qs+fOXF1P8EhO5JA4K
yUoV1/yE6mDfe38cz0CBKJ3Z7HaO2WvlpgAU+iKmrokVSKxQbUQaNDTWgYdXYNl0tvKxCvMx9Xg0
noqFD3DtAWByMFleoF40VKLYc2RgwN5hBCaAwgtOsOkW4AYv1h01ZbhdXvDBVRCa97+48axHXljP
oiakr/JAkcYN8FU1KVmJ/+S1jZl+/26eyZ92C8OXXGycZ2gGgb4+D5eUJT3VcEZdjtW5fm6zn9Gs
J2+S9haF9o5Pdy/nZWaMRgd0nLL+al1RSkThQQyStUAWf/Clu+awHVE/K16UmnSTDf5Zr7I+jxMW
8B45sVH4kiqpg4lmz0iNBTPnFc7MVHIonMav/2YBdLoeT3LYnmEGEsxcYsEIGelgKMHgfj+GjULS
LAQ5xn1aKF48/fQJotjcXu35sFITAR3NgPSM8sFzludAKVOeXZ+BKHJ81XaCAw1IEotO/rXCNzQf
/e0E6/aAWrwNfFwsJlZ4FfVLL5zvm/3S+q+WKEQcN4/Z+b5U6FaYI7DhmjyRWO6eQk6lRZCKyAkZ
2BF2NkuikRkekKPmhumzMyjwYX9HeIpBykKEFsH5ss8YZVimiogtdTVqlX+ryGSZCrucdlG+AZDF
mEVObBUgSn0tSpQmdnfwj9OvZYwIMu+808dFjKoPQa7pBpH1Zlnryg0P1BLJ+dzyCfOpKSGgqPZK
J6iGVekSObPYPo8w+RhKQBd3J+u7HjVZaw2N8qLZBVN8scbEbx9USoo22UBFV5XDpUb3eNdZj5oA
Xrmm92IfnFEby6f8jMUnuc0xXth1OB1bw3/Zpxqc5rXuX9nEBNN74JMVjSpMTUUK5OLH+QqETSEg
QYY7NP6EmJRQnOKt9UvbWLBoR+1IdaEHa7Kdtqra5/ttZh6cTLK7ZQ3iZF9FMEZzG8PdQe9ZL1JU
nnP3anuOAf5jleGCS5Y2Lk9PInlny4wHt2k1rYTgPhQUTILKSFocTOxh4XsoFyPrWNkYtRIlzGgL
86vswauXhqhd6bw1EnlJXGisvWKkZy48eKBMBFkivg46a3QLtLU5+xe3qVbayaduPUd26ODzmP6V
y0QYM7VM1xUnQ+RCAfguq21fbvwMghARLzCYjWAst2TVBAgJNmXsX3RZ5TW+dzf9oluFvzF/eL8e
3BjVj9tAxEO7L5WfUAO54c3uFLZEsLRGTA8Hl7CT29m84z5/PNz8olOLePy+tO6ztYG89zrMIZzX
TBzyilqw3YcxpRPo0mAGFTDr4zLrp2jVXKZITbZMuihno2Uwdds9DcPYo3jIUSAKOGWZxn12QIdH
4v6h0JneRF6Yxrd/GaQyeMY2GMZb6ROjZ+ib1Z4WIL6evV67diPYiMg6wOmwiqjUdBc1DOTgrDmf
ZxDNinPs0Ysf5k1ghmcVd4uKoGRbnRMVPjK6KyswnDCypznqq1olV9eCRInPVh1Bao+U0g0YQB9H
iUEva8iPtxbGCM5SWHNtzUZBGQyRBL9XxZNeBO/nA0HPy97cQo/AAvNfmVUJpbRl5is/woTpdmMy
BWkizt+3zg21vJ/DlBWrktZDgaCh+L5iECo9Rp+st5fOfi4tKLoz6yfBKm13B/+CI1VnnjjH6iNc
bl2A73jqGdzdvi7kT0lADPiZU9kXtFxANadDcqTqqcoPwuRCD6tgh771fTCBInVrBWw3xA7LL8kH
7EbgZBrVyk0U9dyFCcWf73VCtWS4aq0j5BX9zawcSw+cR2ywKZ6/uJwgSIJRTuyx0UjS1FpwZ79A
kl9Mx9S93KB+OQubDXDcG/e+j73EGuemaq1QC+sYX4PHDDzdP60Xrfis9ag0AQi3zqziP+32cH+g
0I8f0inKGcIbqDuMrM3ESka2swNjCjxKZn4yrHBL4Kw8Q6C86bmBO0ce3RxlvSGmdOWXzkyCWjlr
vUccR2rItPaVN+jLTjbwo9naEBtvDP3LUO4B4TFhWZCP/d6xSak+e9+ZLVERr0kCGJiDT/snABSf
moOr9L/2iMXc26UuZdJ/QPuWLEVC1u+Ccp25ybfUd+p6cK7OuSPvkOqqPvvgxLIt9WKHnBm6HyRv
B72t95MgKEPzVy2SU0e5SV4bB92ropxNbQDW6x4kQrsr0KeLg8mvJIMKVs5K8Ui7nUOCfabHGG57
43rLHEyJa4yvgOgTnZj8DwXyfYoS4BCh1yYPxOu6sDTd9D0pCID+qpZ1Z41dw/arwPzV4e/NTEqf
JerTc8lgCP8B3PoUMFDI/PEzhkIpC5tjGR9mFocqFc/4g2nj6bYd7sLslQfJtal4ZEoyREkm5NHy
elnaZk9PkqZ1m3dgIWRX5nhYOZU/937mGmH24e3XiDo/nR9AZoCAPGHfJ/UwK+Z5Yg8Hit5ML5T8
NhD5SU/dMpO9U3zE5nFzR4PPrr6a30sKfA+0UXpeQ4cAqjo3suyb+D95Iu0qjUlUvKOe6n5ZrSJM
5O9k185AG/Qv7iSbMQ+GmXQESk4vL8BhqYewVyoNAtvTeecXaFh8XuUZFxx4jURG7I72luvWoruf
QpcHGBYEqh0hHcWfxiFxsHR06AiUiiYv41pum+hYBkiQ1bEESdDmh8p4J24VMCnkkihO5zSOjGyP
kbpNYN1LmQ391Nnj9mP7arEmGnVVxdlNROuk2VWOUxzLmfasx9Go+BKlWhMjnqFDTuwBapxjn4Qk
SV/CADReaF354ynSs6QMhGZKvGsijyUAO9lVLoJnPNXQalFuyXWeisbJXhteW4yvAmFvQudVpV08
DmRjDKij8qUc8cPUC/LB40KsAvJRr46xNvNJFgROYJLcJ+l7FsqCcOXXPsac0dNOOPftXRpyAmEc
QkoB74G0jsIrZXmsGqjBSpHtBSKpRBgn/4RIF1lTHlnNXL01EqtNqlXiuQPm7FyTfKbnZ6HnnlVV
ewYWJ51QAatQu1XG+NrtAqo7N4kTugZNXoLOzRXzOWBeg9m7OXFNMyRF5HLdYZD2/lHVi90npDVM
VT2HFwMUhb0mwkOKG66OYpvudZsnlBRHvnpiysbO5KyXJrGCIgtUiZAtPBp2TzFbB+IHB6y8jOAf
CijIhs849IAincU6knXMWReojjMbtmris2QWrXRaIjnWo7wkAIRn24hg2frFrerRBPEVgBOhpQIS
hNjmKbBNVgUsVCQTRjhhrGfrPR/H2uiOq4OnWIKK2UPwDALicISiOm+J/tGNAxvXIFfFQm8zXLAw
/VxftDHGE9Wu1pWYb3FjHFiuhUuZKRIcZybqbTXVSwbuqxCj/mmwHjuATkPaTAy8T0KzADEfye7d
DSh4lXAmHaWsQs3Oo2bUuHzWg3yseRoeq1HYIunrWu9mR/kTpA9D37Yry4JQfQAJe8y5yaMcar5p
CQJtZUOWr66ClorZCuQmaj3cWcDUuOPv6jisN89EAhQ/BhQvOmOdCjFmIwjp+esv5mauUC6V3aXG
HPhc4yixAZk52t+1Q0PEdEDyK6yz9OgdPumAHSMUxhBJcsIzDZUXWxrQOxM38zkVXdy6/ZjM5w8a
o5Fqosl9cExwoUhhiRrrSZdcMMsyYp7LBmgYdEWrJbbp6XRIbLsaEfKg2UO4RkjbwmjUYqMq1Imp
yH3jLlu6nAzwOyhUdlH1VNJkW0MtnW5WHhqJVfNNdILOOdwPtdrVF3FthFY9bgxOaJ38rKHiESdN
0nS/DGW/+gexS/qcctXh36d70TtQUGROwN3WRCZwKtqbqn41X8P4s4wMGuFm/JQ+1C1BcI4ixXoI
LacXgKQ0benLouQqNh7mweCpVGWpM/caLnulVGzSbLctGzgH/bC8kXAr91G1Ul1P2lBXcdw8jEyI
fM6qiVlu8je6rm8JpT0IA2KFA9CQKID0vaOk8qYEZcbjex15QC0P+Ol/bc4lEvoK7Z66mL9J4nPl
AAt4Jo8Y/rRqXBfz2nPokrp4AxxAVJg5H8CCcSUjZjTYH8LJxHf2a4oAqHYSKWynN+Rpk8uCLWs6
TyBXVAsoE/NTPVaqUnWNKar/vxqXOl2FS+u7CGQ/2Pav7E3m/P+u+kqvBfm7tU1urrsyDEBCZRzR
4e1Fx4KJmafW627FFtkea2NHFGx0ThDD4PBT0wWCfhpEA03kLwmkt2/lxhn9zRvoN7jEZnDFiWOp
Il6wpRRUGf0z0i9GtGwgtZqzp25qitUxOHYp4Dc4irVzN1BjQ+Ko5ah0RqvEEW4AUVEBkvw9yml+
iYBXsmricNEW2pFZ1gYDQEy1yrl2RMeCN+9US5RaqPf1wlhxRDfcGQG4CQovC39m535h6GFop4b6
IA+1v7sWjTlLP5mT27QNASWvw5nxwDFblziFgaYk3P3ZqCFSC+uHVkwqizS+6VK8TNEPjAoE/vQu
BwLmQ433afcGkJtjPw3fFNdXNSxKCdFr72U3ACCPMcsqpfuManC+GkDmVXdX+CGUpmwmgX/QOuUF
p+XKCGL5nB52KvYhFioHg8LFSPK69eKBtQMO5A9k1dW90ep7wgP4vVgzpVpSZFjYm5uYqMUq1zPx
bMdHNFE/aaWujvWisJYYTwAHa8JdNHP9jFOCJqZI6VcLv0fyEkbNvss1GSAQk6qRxJjFXLFIISTu
c7kPnVvMBkZUlBJIf+ZTw2WotxIlRqr/7Mj8+OTDwoTpzOfDO47PmBn99H4kgLERlJWc6NuNoPGP
mrebKoyF3SIJwBo0Ht0SrnwR/cSvob9LDX96foMfvqjT6fg9WXO4grdOxPgLs6GVn/2LyKYdLTU9
2BrrPIhBEU9DwUAvorhuyvo0LozSaYOv86Tx1cKNkoonnaKGNcLfYorOleJoUwZHzn7TQdi3EEw/
Ou+tRsmjBAZH7Ba0f9A2qL90xR7P9HPKHlvod/YrONZZ9jHnTeIeFa55JamGDns4SFjGkl4nB13L
Trb1lFeoPmqWP0w7QrbFtuFdukhi7JIV+d+WQWvm4BtbfUIYAsdEsEJdmHCJlVgmkeFYa2IoltvZ
N5cyCU66u+ikbe4QNNkTmVL5+BcVL4LRMtmLaJptFjr3Tzg6QZ9gvXUJHzcvCtg51b7XHxss7zXd
bYmkd9HvRH7HZ+WW1BDE55PfVZ4rr6lvWBHfSWt4gY/7C1OGtoZUifM4XUQVI8S/eKrROJHt6/h/
FyYYUj6tX69GOFcmZVj8tCibea75BN65/v8NVy7lnSz7r2m7p8xgJXwY4AnZU8MBHRoo/GPeNMMo
k9QvNHGaAwpeRgFdOGyFb3A3/xfo7APyLgzqC4P1liCuyB4eT321l/81FJA7w9adjUFUYK0N2Tgz
UeLeYpzVVqr4NK5P5Ih6YlLHaoSKJJwyNdWGhEyTkmGPze+c63T1ub8UzRn1XsbZLjewP5PYfbSL
mWLyrqYjewAm5MPm7c3YYZum6T+hBZPref0j4ocLcnCmcVHhWpa5trlSq1+N5clFPN07qtMlUNBH
MYve28d5vxc9uLDLg0NXfLgWcOCyEm+e9omRlnlsgQY5oWXBoJ7KVp5eQ1I55vE2Do69N6BBGEn5
MoxoAcXUrxKoyWR/LHRlnlBeoaqix6Q6Q13mP4X2oeu5DKGhSTxyY/lBkL7NHNq/lcqjqIekpQ2O
9ZogiMpJKuVxxyoRzKvuRjJA/TWfyL07ckXSuwZV3Hb9SD7Vewu75oJNd8MReFwVggaYeUY2+7/2
Y81oDYPGFSp22tjuahYIOzZ8REAQwrID/Q/UeJlmeWGbZuhuNjGjGdSaDvwPO8iCifhNQuyHCvH1
R/Il80fdnBMdqPdLYhPaqHh89/8By5C1FKev+rLPrC2NxwkVoa2zCWbW/qn7LdetoF2ZLr/noDWk
qMoZvh9DAv+bDkNg0ETWjVR48LTJVGMBe3eUgcVsz2wSyKeO87E9C+AwpjZzPBpsP1eTXgh/s/Yz
AeIfvo8D430J3/OToFObKTvcm73tDHT3D+/zriMhnDDJrt7LW67FhAoG1hGbJaX68L/xkCrLCBac
A3obn/nxH2MABPwDtu3InR7JLVV4VsbUTM66eyrW2TYmcEjEhl3c4WlivbXwlj0mx1jBALobQJRQ
oqCd2X1vyxbXn+dhIQ5+2kn+ZstXHEk/mBag4DeZylMEY2TGL/o+X2QuJ7YuK1T+i9m+mDnkrD11
HO8oATD3xvNdlNA6OzjLaCF/OFKe71sOafhR27FJRAW/iW6RspbYhg+GUNbI8LMeVbjYBOc1qbxd
aJFgDGfMVwUxAO27XMz6x58QiZ9Zg923em99tv+PRAFDltsSI788N/IQDhTDUSpdZwW9Wp6tJJjr
S+RDl/thVxnpE5iNrrRwBgDiBynsAsR9wt0iVAmc80i70GikJZCbZ0fwufFgNYo+0XfgufkEDS/f
KUwO8RBjQiNTsG74jQzG5ewX+aF7+IbGZ/lcA6fVFmF645BKW2Ae1V49BOn81c331V31L0K4LBnY
Ly13hW7mh3Ems+WxA16/DLHK4MFhAAU8xjklu8CONBYlPECEqkYSU8L6ZnAoh2CBMGu0f0w4q35p
35doNYc52akNNb9PtuB1JpBRyjPdN6e7+LbWYEAvhUrCtyef/Ol4AGaEsGD24faj7bVKNJW8XkR9
qlSJYHid1dD2SJfx67IdzMtC1Y8FGuwVk/CboPhYByniOzYmcPvy7Qk3UxQwtfbPHqXrsDRWZoO3
03Q3kJUeEzuOL8HcHIndnLZM2OCelghlLWpg1vFj/2DeQUIPi0ykWnd9f2vYHnp5lh7KQP6dBXfN
qlAT6NPxjj3Nm4/ooRug/7n7AFQ7zFafYalXfr+bQaJDAI2itWgE+SgH7lVMZEivvF5e4ycvXBvw
PiYtrzTA0j4pSpo78gu5VX03MgG553hwjWfwK54TbQydrhQBDTXWIycmDaw4MmoTTg16iBeO1AYj
cVX4WkXa2h7kBbLrA1jQxRSxQDHgt66lQihV567nUfbs/nuIeB0cTNjNpsBoW0LCnWV+7ZpsipTC
6P+L5987J60SVNAj/jyb8stkxKu+UqaS212Q4VNLE4OHRl7cdRnkbBlrbR7lZDn3kGn3/67eXVg4
LtAok7dSGFIcIxzrLZLA17ovRbhbKs3ugf1+kRQBvVYJK1P5+pmXUb0ZRS2kYvqY5oD9j7D0zy2s
W1SJ2Eqfw2GgvXKmBkTZBjxlY78tzAh8IohR6SQqxmvU/x1+ObxQc2sZ0+TcI3pC6oHf36Yb5+Pf
GnyMMvJ1CCRkFXD8G0zC5E79pdo7RDK9nZlNuJxsjIBu7kXzMzZS8GJcgy+50G4SAtHbs3ECDF9J
BSi316cvBUN3wDC1jOV/Qn51j6XrVnsF8KOSXFN4vMRRBw3EazL8+6drlN17zW3d7KWg+wePjaoa
6QiSroUfFeW1EgLIq19xyT2Ktea+yvSGMipYlNDB6lSm072YtdLz8UHeb5gHJzikUSnM0qCt+g3R
j3iQndctGqn+enpQfjnc8aNe+I36k7lQYglUFl31268QtHTprh00Nc2+FAVeXrZdkpe5ia2r4rRC
Kr4DbL6qxbCa/MJS1ESRAMFBBpOx+hgrqqg73b3v13lOlX7GEcEmhcTX4gF4PyeFX+HgH1FUUQvK
EanJHT8Palc9rSjzvFu5yUyt4+iYeuARtoEWev9EGRHh0JKMy3lpA0u1Wz/Vi1MfwMjsayAQ17A3
jz0Vcc+3USoNL+kQp6UvyZbLg5FHOVkLjS8eJC7f62v1GyNEg3H71zLQyKmybm9dXNQLz+SmhKER
7WwOqh0RDMAA+QXevbHHX3T0T2lJ9Q0tFzFfuyXfLW8t0ydkgPOaNDlUrXhGv8zfM4lY5qkPMsEv
QCB3fHJD3bGwqPkZVk9396Ejt9LwwUdTEbMpJOFrWO9syCrFcjuFmxDmJdiiSYvKbxgxlLInMBBh
tdU3dSqB7y73FvRYSgR5YrlJaqorAn/r00X5oyfP5Da0vdAbQ1W2j4HH+lubHsIj2fkFIYWzC6S5
vFDLl2UREXGwEhypHGSZRw1zdTVG8ip+H5Ke/+P3+sFj0FVDOr+mptb3lu6xtEg8ySslwFE1EmIh
Y6uVcV0y7ZcQxeqBrM2BJ3WwRYjNI1FH7wlYK9CITTskRYfUWiTmAvf4DFBzNspZEVqVDim0hhrT
6pXu+mBZi5+d1kBDIzFas9BiN299vTZfrJjrdaRiS1JRotPqtmCxj7hD0l39wETyhSpoDrt1TyPL
BrzH/+RK/oxh3GSHsm7TQf4rhWTZ1Q3qveRB4Rc4soGGHkzU6dNOLvcmuuupdMdoa4/RmhcgMFEq
6YpyMImJ1NI1VAxgJ4pwoKt8+NrYIhBHzVvu5zuPqUOUqjU7UH05jiiETcJjbPZfXn0sPgowhNmc
PbLIJJVLylKoUhr4t1hdIWkN4dkwbYtC88+m4XGljfmMHCxJLiKXd8vew0ZFgj/apMVdnFGYEtBs
h0sQ/+2eUvygTiu/tx28bcI+wE4cGlasVaUdtPevmbIOFPt2SiGRD0Hdcy4CZBcreb5L7Drc67HI
EnAzJCLcV62ux26ZzgsqF3NaxNumqvP6z1tsg1Wj9lePqaYPTT8Uba/jP5EjCH/BJK62xUxI7mdA
Y8pioAakUfo283bnt7vUrvoopE2Jh2YsOiFKsES+8D4wUNLeLElB9yRZ9EBUsjgabmD9qjlG1vYL
wDPCQsf4buGrKYo1LJYnHBFQbRR13j6xTNYQZoN2CuldEaOZPDgVNrbXMGJ4M5uVdet1qPeqVB1i
xdYB6moismF+wtObGT8mRuYpO4UjL2GW0+IhB44Vj9WdTpxFt6d8zqQqWiNAW7D4ZZFLPubhyAKQ
f0cGXM880TBm8xkxP1/otQrXVuoyeUg7vPRZKmFQLYip6uq4arFjBBWMLwdQmUVtOI0P930vYsl9
UN4se8OsEvAqyG8oqE6zCXysuFpoS6MNBIQHeCmUyfHMQ0ulUrYBVVxLU3ZzA2XmLq5vvPU75QTw
+ijoIcEA7+/IQ6s2c2tPtyOW3L0eSK4kBK04MaiywEEJ9Trb7taSGcDPZmZ+d4WnWizQFbCJcHZt
oM0SM0zbuxftvbB5pN1ImUrt4zdTDPJZ55VZPWBNM+uelo8NiQ/CPZsXYHpCtOl2WKtcSNMIDD2u
2zG/yY+r2NMKYO2wfaxITbKtNMOhZYKiemOehWcCE3t2AGQLYd+0lSxnHy9jqM9MvZl/kj7CfyAJ
elNGGftdM3F9NbyThjordlJece1sn58tT/SaMDBTzSRLZkx+m51FIKvJ4ivulJayvvTQpYhcoehq
aGl4pLBpkFFYtp0Den0nRcDATyrV8JeDjX5UKqpAMdv6Hpy8f/WWNG0rzM0PLUo5BmS/XilSwr6q
n36J201/h5mDkItwR+VHVLBGhzHM6mVlfi04cU5CyIqgMrlZCbYk4PraoyQl+quUDjYHPDdK43s6
fMdCPZr9Rihwd4fvkHxfpTd+UzVWMG/PKRm/C5wZvCkoOWQmcITNip8ymOrOOZp4OsAmVW8nOty1
iLecys+7Ab6V7+BcldArrokvsOlIh1KwVUtJ5IfO8xbjnRcBi1MhAyimzGiwcJPopwFC+Lihad8p
2QmhOtTLvShrqThlojqZLABTRySESSF2LyONho3Tj3FyebDb/LyWsI5ZBq2C/017bQLgn8d1e3lp
DnrEzFp+Jp5lKrKL65OUc+rJntjOzkxenuCdz2/8VCasGTXhORX5QIS7BQV3u5X7BIHD7Ud5qBzL
imZmqr6Wcd1/ryZaiAUpSPUyw/iHVcHcNUbLBh1BtPkU6c2wMAn2oeS9RHvPq2dH42SKJkGG4oFd
e0S4DG4aKpw1dS4066y0FvHLKGEfycx3sfbMfFPAvncLnaW8wPUCYjsOhiwxUC0E97DsKRLnzG17
agFM6u/sqOqK5aRp6Y6imI2iqMNcEuCjqKCl5wSjqMwnU+NFetml5frTof06g1VoSJpOtT1119N4
7XEy3exTtDopjlpdz2t1AIqrGWTlY7lYXZpn4EnF/mWYzx+Rj0XbF8btgOMNKbmcw/AyZnNDnobj
Ke8rAC9lHLVEH7/ce9Ie/4MQ+CtjHgfRHP2lRkyygNCzPZIDDNPip9FkbIkGQuFLC60IAknn/XDc
iojN7ZaTopJEobG5Ao19k4JpVMRkJ9SoJO6Wcjnhl8X8oe0+yRiRlim52apGIClxealCTUZ+ahrE
mnL/OrdkZBad7/8j3xRf34co2iivBxZDgD28urvmqC13zl46EBb4BaE7uztr52zWInzya8dSIXmk
kPWuImdqTeTOCNMV8r8B7ubnaic3QIAVaN6Aw4T7xF1ajwMIj8wipPa+gYaQ4R64PTG5q4Q38EjN
au2/vQzk9qChjOlwVwl5i3mH7ouL1iHbw3Sj7jlWB1+PFo25kHGmsiWr+gdYwhw1DIwreZsF1KgN
InNByF625y1ipjWshTm7CCeLm2wYosBKVL383wcuZQvXR830Gf7mApqksgz0ZUGRc0XUQswFwXNX
5UJBtPBEnQP4Rp1oRsTObcEP1VToHhHLx99KToeB6ow1YgBqIc9GyUN/Q9wsH3cGdcKhqwCL+KTr
ZZvgY3NaUq/QPE2SG81UXAzSaa5akKPk+skXDq9I7l5CW3OZ3tc9ooKb4yyEK+G6sdnjw6IYHFLW
1zaIOSDyn4Gv8+t78uZ6P4+yqXWrsborXOMJg2K6JP1oCYQhl0tkXESD7BA17rb+5HKgn47ZvgQJ
MqjNqe+x/cupJAVBOaGLFqxL6zyCnd/I2B3K4bitXGj5v/aRU8k0x0uGyv/AEkyPRKtsbYuTwiA0
NGd3Y7dA6QZyetRu1vpyS4+7z5fDoQ/B7Y5rF/ilpxWofe3Vuz+Axqquv6QGCqoA6GzzKVO1q7cD
ixE7SvDf0V8DU8snv9ATOgZcz4VlnZXT+RmK3L72u7/Vzupivdqe1cUXkNt5QC8kdpRvfUxUczJC
+5N1mz5c/AropJkPJX3Q8MKoP4SwW4K+0RWwyNBWvXqzNxnuGwajtHCHy2yojlUhIxSFnj+QAA2Y
a7xA45qUekANFEo4tMEzGIBk12XDIvkvV9yRESrt1EyWFA9lZ9a+rgEcfIfe9nBHhievalfRA3NR
zA82n4/plzE+6Nm34ysRjkhI9QVOT0rYTMsUIutkBwe4Y1h0qb/2aMmphINaC3cSAA7kG4fTXnDv
THay91DSuOfOCmGuZL7uv6aebjY3M+uumGn1VJHdMPoP2VORGAkwEqlmWvlDhkyw08Jmd6hMgUVM
kEeaCoBALFZnuJ0u7dyZQGUg5BvlgiomiVGUHE3+XATypPpsfWy4PTCnXb9i1IblHfB1mIpqyWKw
kfpk5fZpW3+t3ghPgAe2jLNk50wQ4t5wO9ikxO0K0PfSytAVVuyEo/+R5JG5CmSb/eB49pxsxcEr
Phjv+mL9/xb1525Ae2SeHbpJYha2xi+HDWOph/+xp6GFnblMeg7QvYosGK9QPP3wU8GHLQfHJkPi
6Bpfp5w4/zdawaS4cqXeD5/miYuDMFNZyFc+tT96AdcIWbwjJgC77zpnrvVr9RMBDQFxYLrHCzzn
XO/na0LZItaBRYYDFsy1P609obX3MkgQ3XvBhSGAGjO0udD5qrTT8eWYgo7haB/LzfQsrmU8om7p
heN6tFzAu5dqd6jrBovJfG6MWOul74ugRNbDijJjcNeFuYhbaXZMEXhelOr7MGCoB5FduUVC14lY
eA653PQb1/D8oJdCGg8oZ1TdsPUHeWrlc9pgDhNpUdUZMsa6fGbjV/3NHiuj2ndTH2rdOJ0lPSZp
sOAK6UH37u2WZiTWnFuPhJeSN4Jf4uU6/FL114SoW0EK8tX7XWxKJWu6pLJmqru131sfx+KYYT43
zDP0sECVCuGT2r1a86+XlVBQw1gglX1A8SWm/Lme7bumSm6dq+a8TvATf8nRBXnbt4gSNYqlTiWL
lE+IkRBmsgABmEtsrbs/brR3DCDkDmt8+UQWWUgE4WXbvIekT6WyyWk8paKOixEx0NsjhqyBxH33
6W9XtA96RXL7Vsv2xSXRwJ4CWVNYbhd1mKlF3oL/J6voqBSaPnoK13Qbw3HgmyCvYujXjd9DocPC
4rPA40/s9VjiNtR/q/5TdQSfIOd/uuQeFpB5rlEmSbrO98BDKCMp3ICtTPVG3reTZtZxAs2niGc1
u12v97DIgkUN108qdkpOjXyGGIGloXGDSrts4I4Ck5oOXW4D3jZOfZ3aZUPj/OXB0uYYlWKA0Cfd
bXAW/YC/f5iqd5pMWED05j2C05S0jeWkZFKA7xSvf5+Hi25FASjU9IbopfzL52GdvkYgdO6WN7A0
9Y3yXL8K7UD8iDjOYTyHP8KD1ljgajn1/dgafJkDTE7+UoWns+rW5A4ro61AwsjCfekOiqba4/rC
HqB//vBRCbnGNqwm8AKDQH1Ymrn3xvpiHbirgirJw9yr10JsvLJRA+MGL5YCaz9HgC6j5DYjMH/D
PWxSy8sGoEYoAw/KW36Mq++X12PXsBR867xGbWlDz/ZmcmI0IWnQrdZAX8cUWl0KdRULcXROzTT5
NQVjfRhFm7BsfH/lj1lwS6KajIS8hgfqqp/c/9+QMFMoyg5ud4vINzwREmDU6CDesq0s+tql57Ye
O8NU5mhfdB9XTbQXnx5L8rZC9u0bf+titztdXC3ZEIFniAhJGA0ds93yaG/CyvZ/7iUiH49jdZu8
EXfsLYvM1b5jB+w+BmAaFZXYZuM3W3g3S5c+lhYFQI7QY0quA7ZxIybvSvZNYSPeZp4Qa3JZSk3x
Unc8HaKPKdPWshGzophxq3dAdO3t4QhHfr091UOsfcOWYKaFdGQDQvz4ERovWF7e+Wb+4CajrYeR
RtBGPrlFRp6v4hIQMcKFLTpPsO3J+sDsHWZG1j3zI5y9J8miVhGHqiGohcw43n8lpofDYzzP/nE+
+ray8kGdqktnur6OHzxKxeAA3rHYc66lzXguEG7XCTzdpar5NZYeF5fWUfF0lBPCFoRs37MCR0yC
yHGnkvsZng2/SfT7BPI+ja+mwSZqxxuMq9IPj4PzcAqSi3rMNtFIzk24Rhr8cQnjEBMb1e8bZi9d
D01Np9X5EvvMmPuEStiKiurMO6tzvHLKIeqWTujK17SO8usDPPmf2ko0VT7AIpiMl6I+rtrStgeH
t08aTassSh6dfyqIvwRbd1zhrsEQCSa5ufMOuHgkMa6W+rPqloG94nhstwWPROtvWEk64UJlVHcV
BZqLWSFFXdB39osx9TsUU08vuZee5ye7N3Zy6J251IVQ3fD5326lCW1VjGsGZX+WiV3uCbMrijmL
PVA4QFWNrITFt/XjDacsR/Sj5FJ6Q27vMP+SdSDuqoQGiX3tp1XoVhB/IuLDRR81pn3oVEz4XOxa
RPIuEbZVh/FB6+3wv6iRDp3cZqSAlXgTUnelNNK3umA7MwF4ZnK9WaNDMqDbSCK2jvcNvrBOP9xL
XaV4s6feGNaHlcrOKP8sZsTmXaCeLVYLEtBzQRhVu/zdb9OjOdygI/ZtcO0pUqPOa2EjAai+IXwT
BlwW4pXKReoY0z11ehghA27l57vRE+hJh+YjDFsZ/XIHPIIAFo8RkWaqZI1IdttvlB2bMwFVVzIm
x4zQLmmTpabgZ29FHEthbpLFkFlMJDjQKBehEotyPdEkNXfHzvy8fcuFOZ1ung85iE7r8DelBvoW
NmD73jP3IiGpEisN/0vgsehjM7DkOz5GebFsV6jpRhM/7Ma5HfnjjrT/J/kL5nwQGZT4XuUzEOT8
qHppbuiJflk4rVGWZmBeX26haDynUYYwXBKZMtxU+6lGNc5szDTXSBdAs20VFQnqZV53i4VlQCZh
PYeoOgVgNFYFQByIdPGiiWrJv58DR8Q+e9kHnF7TgM4W/HpzVCgsrkNupsQug7hrs+spazUll+zL
mUBu5nrdKnVPiwng+/wLQuPhMg7VoCS6J4whFlFptwqi+1LpjiDE55um2FQfb5HOlE/haER0A2+y
v2wT2j1f8VzQMUxUthNb+8Vb7vyhOFYspWkyIEtEeYt2k6qtEKw6G8kGRHtssTIq3mFQ3je9KwJk
C/ioiwEE4QkFSeT6fjABrfzj7Oh63QI9CWHmxtDx2UBJh0YX0LTqLGQy9wXUi3a7bFAcwAybPZrG
m8PI+qLtUmgk4gJ24Cfx+IM0e5h+lvvuSYTMid/P3UleNKFUEVO1MbgIPQoWeathTiL370r5U2vt
1Kd0fKnRTEsSfKiHWRxCrmRpul2G+Yh+MftuTM5TD2Q3nGBgkJDmkMKvv6on35byzLMygupVvPp9
wxv36/J+mttsQ0N3MBBlOR5e1WHrqF8o3iCYl76ITJeSW2RqQA0WogMRP+RjUTmXAU54DzpOlLAC
d49Xkn/Qb3WQS6H7qjzVMiIHdH+h8Ndl1ctyE2LJfvOaC+p83Bm60yyWy1vY7F7H6tlDXblBHvGw
tI6BI42p+ouwo7xBUU9iXRdg0uIcO48z0MI+jZ4eqhO2WA7lsflR74f/k8GBBdwtpvTZ/+ztxC7x
5Uj93wwTcg1zvwYcq+sHcMsVtUYyoIafcT3lgkqTKndKGcEZJrE4mNRT78nOXQg/2oY53+bEi47Q
8lYd75zz6GuKxpe5FxvabRV1jumlXa5NrtYc6ZX7JDqakGr3QSSqsxhODhn7xotiyvUI3sEGwMiF
oC5t35LzIx5ok1fTreJYVbpsHtAVziuV8SFxIVzYBjaI+6KQa+vUIb75L3yhu3iHwlB6PB3qfuGZ
tOSm/A9PyGM0unun9CsxknUcSxgafZA+M3Jhl1Tuu3pP5qXwh+C+qP8KexOGiq7dSOtNX3K2LOER
/iZ6TxXMMQpeuMpILtnT6YH3dj13G0zfvUmjPEJ0x8M27ZcllOgBLOt8oBvxs6SWmoieXAVomk7S
WpMb4VzCv825HTI1Vyro919XO5txK5RRTAfdqbxtP7hSyNP7QzrYhQN9RpWQw8lRe8+qgTKC7PVS
h2FZ/gSWG0l7CYMaJ88LpWSRYp9lc2bFjfWMW6VCQT40H2B9hTtVx5JucnyCuZg/3q59MKmh19E8
2rXHkjhWMkgG9H/ceKcJ+Avm6/hjgMnOigcC5Z4Hza5R09a2gLQykI9DKtBf6zOGzt4taVb+JDy7
ePLCvGcgPjssahJ4GFUMzSJW1c8aErl0vTc/q+M4RUlmeqYFx00Qql32v4YThqk+pVCBUdqsnmuB
YGPJvP8+SQsbZwITq0l9NQNKNNM4gygCtQ/nfOom7FYYWrp/yDO5Es1E95YmLDqvlUBhDBhOLmQS
MlmfKC4xJOXIHA2LJ3im7WyHUG1hY0pvdXNAK2lGrPl5d8cLHlivaOIWW5LrG4HiKOy9QXcF06yS
cRQtzaNKPFLxDaKJL6nImhBDwucWl4h9qVbpzhglOPMMp6q5VbxHlXyZuHRO39PCjjGVGh/Q3rbd
zdeidihYVdtTR4RnCPW+BTuI5QjbQVpe5lybJGsiLT2pscwntdewXbM+XEF9OwGmkCJRmizEbknU
5t4kddKjaAZkXlyr5bLVNLQUzwQB6mZvSmaj4NnYgl5dzD43/CvFy+Y/DxSsY2jlEg6wGXLR7uM7
2xeDay/uzgxwmPSJNu0KKUBR3aSdfuM83HoSD3pmIk6IEkkxezlMtH9JOg3baBlbiP4mModo1Ets
Xy8dDVT+3nSA6KXyAJntGSSXbF7NhCeGmiombpB81HlC2V+2AC5xJ6XfdcTPcIe3W80HUNbrzzzZ
DunrKv3IbyX/L3qVz7bYnz5VYxLXQxvcvVuiV2RVOaW2ON1tBegLNyqhtHwLmoUT3ZVwAJiXARVz
LdFdosJ00EOuOZA2ssMgn90mi4mr8kNmSJEha5lwRen+DR+0z2pPC8QClHvwbrnrKE8kHY0vF3Rs
WDAzAOrtdvN6DYgeRZf0QGhFeW85/auT9Guo36XhRAq3BqtvPk7Y20TdlTcAoIuB8MJmfmmF4kuT
rECgZ1Hvf6LyiTXHHVQz55o+EAF5N4aUwdZj9u+nDVtULu7oXadQxe35sGGpIcK06eflM38wnauP
QPAkBXmmW5DQJAMSzTCiW+SRniLBCJ/A3tiV3seBVwF7xexvNr7vfWJPbaoZ+aF5XAdBIezlh89E
xzIdM0zFg6zWQjNHEpEF9drSQizUF1QhOrlY7DZ9y69tbv18G7MtAIjb505PSvoXOXdkwVdXefNq
mZBbSIgrn3nalm65kBEIqpeWGAR1e4IvQlBv0YR2NJGSQIEKf7Vhil0PaRukz5VTZ/c5qBGtiL9S
31LBrynHLSre8NzRDRleCTpBndX5GE1EKM7lbo7cRIYvwBP8fzShO9njrdSzEn7c6LLY0gpAGerU
hp8d+vLjGe24MD3+h1PeSGhBeYkKGa8qkPuz+v1u7IueNWlXAthQb1Ht6t7uPmkTXpUZrkIt/7XU
KmbZSn/gYOavutRks6jR1Eits14nzRlVcYcdx/9e2b+BliHmrYoAi7X+wmb59qsr56oCDYg0LEsN
DPCPJzgG+qx6jb+oVW4whc8bLWkMaTPaLZuVt3XTfNc3TtG1Qrcb0InEFOsEKxO7+KsBm/yBLm7H
KfmngV5jjWLG8xhgPNMd4R0roPXkqUhXmnB2ssQXRnDoP/rnd40VsiSdm6cZlKNLqhHnhId8vCph
hlSS4NfaloUWr8+p051SwjYylYR858UJfPllm7kWXfIa0ZHd5ze2NPU7226V04wbAv8QLUU8aTZI
29eSnO9hemkD7u0XMGDk6RpT+/gnoQ2a9pGb+8RGbJ4TrF16R3b7zxtjiVu5DWlXQ8N4u25H6oK4
PJzUHa9kbgkaIC0hRxnoZYSTLPrLKrb8O/elrbViQSR1wEgGH8PKsfU34LkYEvExXEbeZD4r41Hg
LmzvIpHJIMu8/tmVljsL4yerz6JVT8aU4CuNexKb1xqrX5u+x7WbDRreKsDkGE39OJh808ptJzJe
yfSw+a7VvWBxSouZfyQYe4M2uCyXSDLTIp1X+CUGiyYBOzooUFiD6M3iOmvafddRDfLcZXK9uvil
PCTXB6aVW7+wvHj7z713MNDgJnlja0BwN//Wto1pUSEBAEyEvxJtfaypyypzA66a8ssAka8Fqr3H
+CwNIs7oA1HJ2hUrNiYhjH+fTfOV/JG4h/isWwuvy/Vhu7Gg6Qu99HVF1rLJBn+DJhBpUQQ1OcS1
psBY1108dI5FgoqOMjDVW5SrEbq9CgBN5GzqrBhT5kRacg+7q2YE11w70piSxVG9aWBdCOmZHb3m
jqHLfYsupku8MEJEqTdzSu+Kxj8NJqFpCMY1S2m/jpP7/YVRTWQBQZTFDC1uUmYCMRuqjm2p9wOU
yqyWHMH0nWJczH0wNnOVUYPjFKLugq06+kWQlNPy6GilTAJySd/fR3KVwybtVncUf2zbLTgij6jK
CyD5W0kNE00A/BisA14OEBeB9kpntYgrHT0CZI5eOFcaH5/4B+l0QnGX4Fkz8FYxOr4jCJTbXgfB
KZ/ag55nle7bBbWLvs2O6Utrv5rtIVjAKxENAN/XEIWDIdqNTbCaaLpWGg9LD+qRo8Sz9P3PHp39
5BrFejB8wpPFKk8ijeMTbcdd/r3GbtLPlZAwFAnYS8S0AFnm/j1mtr65ZFT91GE7A434qbljBTg0
VoEbm44mqwwcthkf+sL18nn3xfaY/4fsmwZMHNXhDRofVg+LTAwEyDTXb13jZHBKPJznE4eUKtpf
jz4f3hOYzHt3CBNfO5Nbp4phMFbmBs00v3rJnTEBVvfQfY7/OHLENrMNpRgjeserQ4mR30hIFX+j
A9XBi0wFwPucr5OpazTJaYAUkQ5IFWFC/oWSB6AigVWiMpXPFVcHLUe0tFBgBeZ1HwxqA1j2N2C0
rZIGRamk+dHUzGxycJnkdM3edhCFsKPC7O8BROSWDWN85kMT5j012aOwkAmxPo5hYq54sm4Jwgp9
zXxqS78dubsZH0g6+CTXQL8pznqiLx/4KPXtkO7t/59uvoFOApEMGwSysLwfd3CpmB03J97iDrPO
ga/h6t/6rDrlC/XEs/kt76PmwNz71Rcc0uOp71sYgNHpBRojhiEfGqBMGUqS8+TWODSdr7Rrre8c
9s509mJ30leOTiUhBBInnEYz/EeUF8ocsO+daVqtWqD7pR17cPAhxNDfq3RGWPyjGPRmyNDWFOu1
bsYFROjK0PyAqCvgPNlcfUfe13QTGoN7vExfrIigIIsP+BVbK++ElmJd5wwmEpfYe7K4Yofxgxpx
UR2r73o2uJb+DDSBIkKDr4WcCaEIMi9MG8bh4thcOrM3Io2DqiJ2b3yeBcpa7XXnJe+TiCge03H7
5YhiQYPpocBQe2yQzyCa0I2KiOtLPdH71la0w9Tfk4FWhoEyHfSwi3IeDQ1ibIAb3kD8AZ7KsC1l
b/rw+74QfTMoBuLiVdHOybppguU82gZE3QY9iouE636bl+ejyPAWlvIZj9VVtHpPgqFHPBO1ds7D
FknIRz+L+ihnqnsa8mbt9LbxFselruzZ3kqC9dKzXr/z7f085vhqEqN8GXgG+S7NDGeam2Y28vvq
YgDS7B8/uIWBRqUGehv/Si6X7m26D2xof2WdP7GecQqBIwOlgRaxv8FRPutU2FYj4OD06kA2s7d9
YCikH6MgbOYN+9cWF5ssK4YmafXFUgLws9D0LtH2XaH/xA5Cv6YYXhY5cJqoBzIOC4O9cJ0ct3Fc
zORrlaPcfCB/hRghSc4Yak3OXOzgFePBcBthKvE8d8eA0EuzWy0t46fSbr+PZsmC95pf9uAS7WiD
ijtfSA4aYZSDj+bKafu8By/Aek8OojchP1iYIs2zWXuzPuZvc24GwSxWwhWSsWPu8/hXubLsdMrW
pFrgTd9TUSx8EPeEQ4kyQg40BljgS0uzX6hbbtGhorqDW4NLZiUpYe71YpzwECdxCf0d5NOknyQe
9vEUPHMyvLZSLm3el+1fcV9NqRP45BAPIzanCyHyGu4JlY95lDR2fMIIQgpOnWLVlYIVw8Yrb8BS
f6+Lx7u/jFSNr45cin6sDXu7TqEOxT53q9W7BQ97e2+8qcbbrVi+eEs0FFGwK1VGUD+1c/QvXHZq
O61re+1YkTx923pt3G/Hczq0RfWvrhYxhdXSZs5WQos1JRO2xrxCo86N9N+24PHgGLoyhn8kgqjm
rGj7rl0YEmaHujiX6Ld8Dbq+z9HGu+aJMJybHeaaifOmzfyLqyc0SaQjfKyn5XZw//eKiDFSckqq
+zROOjthedEDK5tkx06X46AgXFHM2OlfhnnjWWsEsKTjTlJwONyI0hSQdxg0KBxgx7Emr3gNJfdi
0Abo17OCNUldlKQuteooTgTY7S8bE1JKdn4+CdE0qkaRkITGgKjFAbUWl0fsHS9PwS2fWStGPdrW
uQhuO3rsyHpibFC/xMEVCwWPG8nYH9Plk0e/nR9+Id3sz1KLES3KwLllQxN40dnv/iLbuW/YXRwO
HFRMXd2CkvFD3JesnD8f/0B+6mse+vuseesfDMLSzvqATnB9IvD8CupOk6vojIE+1tILJIb7m6Ev
L7AShzK+7ySn3xnzVeRVARKFHEOe+cjK8KJiMn98OymDmw+h/CDhLxdlNTXKiUbYPY8GtI62H0o0
pcgpEX6v140TA3BS8P6ljffJVamTheeuquzgq3zmya5nD+1sikb3FcANTXVLEHcQvtZvtVT8dMxY
iqKjCDGAXQz79MkXhThm4+GLQjxleN4Ftd29dRA0WYcC+cfikJGFhnguDWgnEhk4BIMpVAJNG0IU
vTL68YzI4ZrjTEXxLcQtAu8WR7hEzXuwDSNcia3rkn1gchs6uo7t+jnaCjIG4D/amBJMgYuzZRwj
JTHwaxoa6RhDZJdh2QG6+wb0CtUgF+vuGvNQnjMxUrUmiIWTMBLYf8/mPRumuCaqD10oUDwpSQ7S
QPD4Kkl8WEAxAYvfzW38PfwYfRgS/L5tEA8/wD2tPtEPBmTBV5YTWh0s8w3nx1MFqIN06Q2FIEC2
9fx8FnppgAc9ffg6suk2ITO0eG6oNIh02dTC0LML1M+pYA7jlRSkyTPSesXty5/lEczZ57H+BRE3
J/T63cUm+hwJRRVebMMNGTfC3j1EP9iWE3IJv32RkdGuQ9h/5llAB3yTe+IMk8AsAD7Rtb2V3DjG
d/5qfuE8arc/wLGXegvDX2C885n5avP2/JO0jHn9tKOvUicH1lJeO7F8KbUycb4KKFnFRAr86V19
PpQzN8KWXsuqjIU6b//vk8PNuOz/egIAxRWv/HaZBKU+hfziyaFPiM0HpXy4z0iMHT2DkSlT/y3D
M/y4DNO+ZscSfZ13mPdHvNAQOGi+SuCbVtL+ysNLGZ0E+oqLh1SZ6JAth8TDVub64EFhnKfM8fnS
b62PRH+ZmsSH/66388sdHhNRfnjfZYXBtNvwksVrO9SKVLc7YPHVqYPQuG1txXWPfO/4ankq4QJc
gAx73U6nzkPvpROukRgmaYCjtbjTbJ+/IlWPR5DIRUm0AWs1BbSMt1HtGpLukhVvMkLkrEf0FZb7
mc0+9I4tyCzU8bAnAbYTJ7HGyx44ooqXkmj3NSjgan3oiopFRbkYIoNkjr6OjIpch1goIr3KICoW
Wl2hr23TGog9Sfswc03jvEE86Uz/lz5S7vS2iAF5v93ujLMI4F9oJ7mNxBTatYYDMwBdqTyxn4b8
WEGrier1Htrk73RvFZ8tL+qNdbaTPIu3VNVhdOlWB4W/8QUsXN1GoczGwW8EfSdWDcxVfou9xIJf
48zH1VeoSGjH6z9tQPw0GZTWyvtwxHg3QjFmvwqqdDlXPsANV9NtSwi9U5yzfxc6tSt7vZCLGZ5I
AZAjPHB+/QobZP+IlMX346mETAymlrYHNBlOgk4NmWj4C4rY+M9Ksc2WubYyZuLz2ajHZpO3NEh7
quJfo8VcNU6PJb3uX3Agouw36wT7izSPvMlKjEiC99U8RapWQCLTHGtonTzdWTKGWMFMUhYtlW2t
4tj99QvuTSrpDNFBGcTgPbdP/k5zOZJ7+5o0rZVZgDBFA5mozUAgv5KPiqV6BhkwS2Kbu6N+0A5m
Hk45ey0aYVowiQrf7V/25igI4JUZ9rVxM//I9V6zHfUrutcr3h/0RsNeVvIO3cxOqOTWPpTHZDsm
BeNc4ka/sUPsJfrmSYnaDW8czqAOAI8/ih3RQbl3KN1JfQh1epygKJZT8IhQnJiZjV026V/0seeX
PJedpjeJiKtX9uyVZOScpB0ilr0DPQbmd/SUNYZSZinLPg/auY1PTOTwSIpIq59ORZMi9MB/gZD3
mgym0vOLq9r/u71XWJ3doPUX6f4tY9xaCy1rIeyOgG98Q3Ovw4HmcmHaqE8zEUTd6L5ieNcP6mUv
Ed8m2fXLWMvy+QCbZabUJtIHgmZg+tPYZlHYger58cAtd1Sc9j2X2U33sI9UaTPH0JnJck/sD8tq
PCSJm9sr/37qcVWjodGF3XATBDhK9qOqh7jbG5Wzc/M8CvSSrS022asSZ117yrGgOpP7hoBVy36u
woamkE34F6Zb4hUum4VnZ1S5J4GkRCRQrUl8mqpCaDJt/QaDFAA4lagZ+ciIees1oplU9SzJTUYL
ZRFT5kk9ndYNPGI2IS2zmtBCQYdr2uxpCwSFis8ZJLYjE+tOAY2twTz+FteppQ8v/IyC8bloAAUW
bwPSLUqotpyqvhOfIb+8GGb/WjzyFLY7mmU3lqIYpCvzBv8rEjNvpA007ATz3ZW5vADVAlSByXJO
7etarCbzhz+ZpF5IOB23oiSLw9ICBT3REjH69xPxQWcOXIgq7oZSYo0TVbMx3Er+LaNClxhFqJgH
NssYz8wIRAY2oC9dtB2G6GNsBbANnuSoFPqQHB2ewew86Cn/LUpyQ7ZUURW8HkWMNBlDSaNsyc+n
z2m2hJ7Bn4lgRv+PD8nfdUx+izF13Oa4C1Ml1q6PlTh4+Zzrk0XfxV0pVdz8hlsEU1zD4QlzlOXM
bDWhnaogUVUQ4eYcgGGUXX0FJ8GRRAkkquQXpBGkui8gRQZWLTPUBk2XX1bHhTXffvdFU5jb2sFi
xfPv9T5IMrnM23codm8VqgRF41OEdpU7qcZTw/PfljKDOQ2J5yDHQr4BCHQHiH1jTqWXigdbrdeE
q7oHdu9EJc36cq0qK3sbjp6zDD2Ry8ONJFmb7IS9CVk7QWLjOGm3B2dHIJkN97W9fmXUMPvTbXZx
M0SjtrN0dyOsIp1OzfFhEe4TCuSzw/v9VDTBo22XJDpaSV9wcXaigmekXj+WYaHOGIEC/uOzcFeg
Hfu6xwafKzrrsxUCUMhM1EUfkZR/JgDa/5bHcp7OYc+ORftjGBqkumQEWJOT8f3ivW5TYbqFyBtT
Eea+zsUE5FRsfJAM1bE75u6dL2mP5/PXKLHkflN4fn23tRc8FlMTsI05kjoJDaf+doBDsqo5AuGZ
icYaYrFNgwWosgOQNTDgxHaQtIxOvYXgcOoAE3HJ/4eZHieMfp3rKGjcriE1MN1nH6n23YPJdplB
D7Pu9YHhQmPLgkQqnNCsAA+WoH8qlJQuGm6ECkoBxNx74FU5lfVYZQwWWk8UG+4JRYVn153aaCkU
qU4z8LENnQ3vgjpIi+85ipSc67F/ha1FnXTcaJ1xINZ7j9Hl/DbW555JLsLHs9USyhT9bEBf1aE6
sRKrumX7sdHKuZGtwMAvGtwAxaWB2HgwXnobEVexQ3kTclNpj/T5iO31++/UeQVfNgemuHhD2wFs
lhZCvR9S6pe9KxFPUbN43AEbDwPMO9rRYwVrunIdKPMuhQvjV3AFtGNtvX4TspFCETV+jQ0xFnv8
dt95yYqPdCyn8Q1iMXkZJWy0xZEm3H+T3bDJv1WqfkPxbMBq7NSGwBTifACG+BpUzG5WOIZfej+X
4djbvFZ3birZMDblD5BlI7RV1P/ocuRVXLAFC3myTRWopotF4DUPjNMYR5uwidLEugnCH+Bl2gAq
uqI5u+2cBzqqFTNGZoaksi4cXOuRJUNgRoJFcXHZnjnlusElC3QspwdbO3jaP4S04Gj6G+t0Hpt5
PCwVUzZK+rzxzanJmeNxT696Py48nOuf+jsFL4i6qIiLcXE4PwdkRkyVlhoHdsixGBKxPA3wyMRQ
bgrWhZFfhQ7WgOqPko29N39w1OSVtKQ1IMDME9nZLmKFNK6RHkyGTFOlvZd1mdGJpvvvxyGXz9M1
oIgvLCcp9MUVQE6ZlkF2C89Gx3ON8kcNbvnm10lOOmgHseMHhoDRc3IMTuvIa0s1CmcyMly6ZeMz
8vNjj3TsBOXsLTidAL8hTkWaGwlQr//LkHL7A0UqXz+URsX1AAlHhv4q/Zul7kzOprF5BIbGg/1p
Afuwq1geRkb/qSdPpEOcwrKP0n4KywEx8LkJsOr44v36ST0ixOfs71NHEZhHxOo+Qw2coEn3AB80
TTYaSyM2fa+4ncVsH/9oig6pi7QL3JkX3xrvCSZlCjKMXeKGkEas/NP+uPsdxB/hpwRUK5fCKmNT
ahJeuOv92dKQQPWxo1beORvlYrZsxT90n94EQ3WP1mCqJWIh6CJjTXnEgpLqQ6OZD14wq65n5FXk
IUjYzegbDNSYdAgYT/u/D7pbWwQIwWcWHog7nfqIIKlGW/1B5/fKG6XnDEUtglgnOOwtembzcAOJ
fkPhWqOsNtUpvRvYB7PiLelGujeKf7MKQ5ZPf6+zopT0Ci9XY32PWTXx+dtHYFo3bIFEh93cOJZL
jnk7V4uNKATVrCVUCNsxtuxNUKPtCeS5fFrooP5JB2+x46nK+DaKGFMR9JIo5mgxB/XUs0Er7VqW
VWKj+6EnVDaQzy0c9eHLgxx511krgGY5JIqg4/l5SfFo2iKCGwRQ531xHb+Gn1Xu2WxhuOpJ5Ql8
BucqlSpnTe5i7a/im6HmTcfZNlfg7e6jnqg2g4Dr4X+hfTSsgFvN006tWEDafjN5yVKztSTjSecL
iXy7ZrRzQ8EmhRneDjXMHEHG5KiYexbyVGD36SXL2iMoLElfD4CTUqrXiK9+A6MDxs/Jp4mY86mb
18OacoiuhV7cZsqtk9R6pUiN5K4XJoiiuR5Cjzyhfe5o81tAiNiH+Vj8BBLeEHTxiJ+HUzGxmxYt
K2h8dblLGBeuiEsg/O9QLkXdMDPTLWl7twzEwlaiyloyKscS2P/H2+aBSV0soak56n6lNBS9F7Sm
DXoJNAayQKoMyA1FJV1BemlZdhN5uLtIghIZooY1WYoQlZLYlf88jawV8olA5c/xQdBQtaXO5t1b
Z5xjIjFRIZ+M6WL5OttLp553oGThzBip8QOR84QLMBHrKSjk9EpCzPnkIDrgcV6msr+nHjC1UOme
Ep6W499lzPsveG7ENyqsThck/GFGqIIeGGHT6chryn8MEsmt4eQ8bWKaRlWmRMKoGcRIq6h2bdjP
6DELNTD+lr6IIa5TslbCMjvCYLXW+Z7Zop4deRt4msuouCBCowL+UB7o65gSeFWrSnPC5Obpl8Fm
56yGdc/YywaFaV+YxPbZ29+8yn39i91qnF8Jdgu/BlCaGesJO6rmxhzJqkozvXmX68xTm/0q19qt
Pm+yDELA+eQRerhLbPa7ALEj+wOMU10bZByQ+nd26Hwf9WLKemrIIwoTX+BfUEkCVwfk0dTPkvPS
Nkmo5LUcbe9RbOhWj7pxAio6vHeoS38CUEaxUabvGGY5b8z4ODC8c5MqdwWd0XCRpkbgWLlm2jQI
jKzF5EpQHr0ypCSNXJn+/OUZIsjWso0+Ra1aiXK3qjU2pzAQjzFpL6YqMUAFdq9gDVWUM1oF92+b
NgwEFOnd89SmPoFRD6nTgFkjJ24JnDD3gs841xi1UYvb7kJYkm4sFM090xHyztqXuABVnOFEwT+A
HMMywBH6PbKoFcXqzUF+DPMwbE6oveiGGv04zNMxi9LDfxOVrMNvA9xgztphxhZosPUCpwPiXR7A
9sBokt96GV+O3nx316xIAQnTGJabylM7dEEuIYSq4g6FR5NgAjPJHc/Kz4BJsJoS6kXtrVmYAXzE
1L5o0GzaB+F+viNKvv/WSX8mLdxEpF4AJKUhFqX8UT3aBGmWxSc+KUDppihr4xw/4CN4YRpE94gu
75jSYf1hP75JaPWjQ6mK5STdvpi7y3SB6A+cc3I+r9IXasd/3mPfluJ+DVieFN2/dYszdq9P3MT/
C1DmMVJMuHAZEz8P43JPtayLkPAnuMblGvD9ep+H8A+6zls7tBYkubJUJcIYEReN64grFEL9NG7v
FORgc+coJVVhgIFhLqIgvxFE437NgJle8G3FFXvSXQi7/2AkgsVUEpt2S4bEY43ss6ActTEMkfms
UMi8sp5ec90mJQj5VWi7X3u8SSpTF2Wp1+Cq/yo57iq4bPQ1Mc7we17h+69TdoFQT6sg/oMtRcaS
RHqCoCS41G6bpRZGGd7lKtBUrRxWyo0DxBcRFbNf+jCvgoIy/6ZLcdRuOj7L05E1uS/EIOegf1TE
q4AT+gcgiX96y5jB32kN9FiYnNId9oU/BgxKBoZ5K+66jWD45jNiRJ+axAh3r9TOsCcNaujphSdW
fv+QQE4JLuBKS0WeiZHBX0ZHYKPn6dXWAg3RfTjaCVN7nfGmnpbONSCQeFP0NAyTcADo0pXwiImX
F1th70zF6KHhBh36vBh2ss3Rm3tjbMqekU+WjZ6GZbsCw1WEcdBIqUAQyxzgCsoRoBR+cFwCpMxI
MYGsKBK5grvn9SMIL8hjTMvpSlsqD2EsWfZJD8natvrTWobqCktcd/yOtU6OI9TpQFJbWlvBXRnV
k34T9m9PF1a5wFBZnCE6jXz+/KH8KWORz3hZqydA2zTfBEh3y0AHSVXIcjaKPImlZw1g/fVszcrh
nP2JuzwwXC5aptYko2nOAjyK800XcshDaTGijqC/eGj/zoQNGJaqo3fytIMaB8R4pbfyReD3mtQw
AkWio0Sxuu7iur/MYiPnzz2XHvEnZBwn/OKSCwXDBDuvTB484P7U1VeKbKs/zlYyuTYoscvl2flu
ETme8o3md8mw1L5d7utgwG0SUUkaHEhrMvGY2+l6JTvnnBZeVoydcRw/ZuBF2kCJRy2J6SRYw3HP
PIIZjkQkAFYnzGnhfqgZxAsKJzGIXovWD0L/7FUOGYQWhKJ529TT/BlQnobYM19kPJx0+3mVMcpr
ATOaM9AeBuP8JAl26NVvy42TuUbQKZDPI5ygpnWBcdJtvRoSSb9UTsX68w5SLDj5GxbwZrcsy+jf
SIs51tR9jUsU1wkkLFWPGBBJjHtB61Dc7uf7oIHKj5TGymxbao6Sgq4hQHVcjxl4oVoxb6Y+5Pjv
vDPlFL2lcO6z4JtXaM7JyB17tC3kLXz8SRlhEBb77FstT1QHmsxRX7ghbnDGk05HrYyJVqtphRpv
4vN4z4a5qikQRtHtUbaHDKAiB24mVn3kGOBhhdN9TY+DknBda+6SjrHmTOK7+ZYCj9YMqmhCw4TP
Q6344pLIhH6wPjvb3XLVCdaB023cnERqEEdm3QbPAB5UyCPig5SfqtOHuzCZSx47xuhD4YvXI0dk
vUDL6IarDq8fTIER0lE8UtCbzDjg5YhJnGW8aT8XSA/pWpTAOiKCQ9s56/z4rcSanzj5yOHnKewi
8zr8zZGLC21ERWWnjNk6xszKJd1AQPIE4bmZQTtlg7wMHC5p+lvqKrRArYVJQJSRWVtyxYKnELz/
fPkjlPkO39RrziuUfcw5mA1HiCOhfbBmYcHxYGpYeIVR6vUByfr6R+CdTUP3fVuCGLMTKDgkzM5/
Z0nIdk/4XTePhL4HSUrpjfdTuFcMLKR6lRfDNh00ball/wglYBSgLqaLhh+Fu/UZBa5LOjO1wbU3
fYomquSn9NmEnioQ8lxkzZhXJVIeEx2mmhPamVphxXDu/BixHOc3RtW2MBgW0ef/kLxBQS0g1YfJ
Ogo65NsRw/RZlmvbMs/ikMf5ZspF/K6ukQFJX0ihQQvs46ZwLjA4mIjrGWZ/XZy5Cw9ydiIXdAH0
XNURIO8RV7RpN9octtO0lSePubc68l4NetVGih6ngI3W4pmBK0TsU4/bOLHs7pX/SZSZwLZCy6Zn
niq/MDBgRvCsZLOtTWwTwwFbBy3SPTImcsr/m233Jmctz7J+6NI6PyHFLerZVbeXMKiUYjNw9Gsj
d9LPFuY/ZNf4nosWWx+P7ksvJIDodHGt+sqU6ZFx9lgail/8Hj7Xeg3k16pTkANWs4eE6vGyBUd6
aSScT8kZukte2FnwZbtwRAttCdvAx0d/0Z3dxZOEOWz7wx9x6cKnrzNC+8Z/eQ/tJ8SRZMEnNeUz
uWvopiLe7wRY4lt0U9o6v/92Mutu7EzrGai/elkHvk2wTepazgWz9mqKC7R5QN+K/h/d3oK3yau5
vKN+Jiq3E7G5utWahGG383QjwqzdCNzFDwHC6ZVmQjfKIbSEbLatBjGAIAviziBoQg6e60VrM+ha
2HoorEs46gn2zXvQ/KdnTBawViavTL5Kzlec19sIeahTy4/P98DfjWKAzSOu6Susmo+jFuHxhOdc
nZQVy4nefijFeutQI5sVAm6rTeLgGZaWxsqU4QsZzSv4aLQEfjBqbrptnQLXesCc8SLK64NdAgNK
he/VbNBvlB4SBV0a+FwXE4wawam6lEM4dw2q+gIR32wzmE6XjFVBAl1O3+dRoAIm8PJo61wW/mSH
HoZLTHmJr/jQZwN7hlufnLM94yjUJv5lICWoWTm1OUwz6iFjDdYjZ5Ycgc9PaWo4BbCuN3+eoonf
WsXJbqBikEz3FU0/BF2j4dFHUW+rxqPdRQmE6zVsp3vL7qIuflg1N5fIfKE/mZOZ2Ih/0epY8UlP
5ll5omNYT1QNWSlyV7YffilKTIjFycAGfvPklYpCvTdQ5nZvvGXkTS2qP7WxpwmjTSw64Vj7+f2N
rpW6DJ28qODBHbmRs32s8hTIfHFlalFxGreWwTQ2UWABl0Vmh33Jo3E+ZZtcwq4vogHFLPya0EyE
AIcc4ydBubQDb7SzxeDJX69lE/AD3Mf4sTv2FpIKZFTmv7Cmi4Xq0lTgcdj/RM8xd5kp3Sw2n6Gi
1vCFWrlKHQPKAfZ4qMcPfumLiVN9yVaxwyGW9VykPlqT4+YNkLM+91tYvfS2vXNDsfFfrcTwREzo
XDFQupcaQYdgf3kU+YHraWPEIervvDz85RS00gjx8eckp4gUsNIbFl+/zTuosJjF/qEA5G7MuMwf
XW7xdzjLyq6Jm5LY0xKBgh+Ouk6mdxCOA+EChNdE4wlSuNU3hV9YM359BRGYl0t2JIwIrB4W19hp
d8RiKYvN9LToKHc+v1w4okcZNz2U/dqRuoPy0kPmyN3UPfbPuskX8xVUs6CjEI3tf0iDtPi1sHey
7rhjgL0NYO+rLkJSyuHI2q6Ju9aMoPsa0TgL07y3MyzeTpxQI4aTQq3244cHejPqRp8+aCZ64V74
VWmALUXC9+q/RkrXLhwNJhysCR9icIXFiUcgMKPjlUs5ADvJIU8adjV+JRGWlUm1x3mHLOjXYbPq
Ps30Kg2fUi/UibZ/u+uo/qV/Paz//hfv0mJ1G9E+7Ge+S4MWHeVJO8ZLD4J4dPjnYmKVRs0gltVM
6qpA+r/AmESUVOH2KiJpNk6oLA1LSkS96iVhyGzrPehirrrmBFNAjFrQAuoCU207XLu6Fb2ENyOs
dnns4AAe/stfj8JX4Qh6ebZr9gsPbMFFOe+sK3XDIwTeA97hU71v4dXugnNEML1z19gCQoTyU+z8
YtqztyX0Wt4CQve63mUp7Sr7Jpi7+VQNOu3nLvu43qzx+siOEy+hDtb2dbjtG+7DhFW/kCGkybwP
NPqDEAg2p2AS/JhskCSASI4WlaTbn64pjhPU4OWqb3pxA1Z6fNjY7yJ3Pprf2C8SCQXCvWBwYbDQ
LwOwZfDOtKUa/o7/ySiT9LImGzM+SGQnoJKJZbIR9QeeqqztnouMr/XbTsxx/wtR39AG90GVg559
lq9SAGus3D3V/h5NO8HNrETAYla+4hazEODlXIF7kYWqkemN+QuX+2ygsuKPgWdZ/QLWtlJlnxX6
+2w7IamHIBdh7WT3nqlz/wFkQZvDvP5zC7WLlLoS+x3ZtDNfhpjAC9TZOECto7SkOdURvW3/yv64
E+UO4zcZv9Tmz+ilhBwqq8ynqyH4FoD/wN3nhgC3smpsNVoxJhvS9xhvF0HFKyPaBt2IxTH3xct8
wwaWtFeR8w0LVFCQM9wnGFz+cVA8orK785v2+9TJwWopT0XpM6qc0oOVgHSUWfxhWXXjQHxaFPIH
C/Y9zhbXPELN9FWOdl6tijr1R11oowQ2kRvVOi1HtmkVXbHnXKaIhQFJuXQCd9R8lczI3CzYh7TX
z9ccIxY+UM6q3mAA8yGCYlQvDS8GyhGGg8VJL7ygorrY1taAIdTV0P47eJROjnHlRQNX7p7nvy5H
qRcU604OwvcAwcVgKgh4lsUVNPtpXTgzWzgba8Db0+KUHiVHwRVaAV6SlKAY4K0Om3RZxRDOWhOM
YTQ2u/DQOrxz7LEy+ezt6kCTxS3IdfqjKDTQLrgUWtGr6Oab8EHeReA4p/8eHWu44qe4Qv8b7Cm8
7hwEskQhcHqHrYQW1H8BL74Zv5fugQISmSTmcK7oxrp6QhefBqxr+mzuZyn/1gBrpdwJ++4K1p44
FZCYYmTGcWWU183qPh7UZhCxvrxndCSt8a8AWE+DxuANlrfmNcHFwSay3MjJ5/SR6R0yuw3/isJz
bKIlT2dJH68RFZFgXRBSXdblRZG8++eegP3eiV7VCZFa3h43hmxtVQYlf2drvLKRr2mH1sU8Zucy
CehFb7O9kcT13GchsrREpDhxHT78Ok0H+6vIa0o1CoqZFixSolVtMnuVMEJWs377Anjxj0esmQJX
OZ/uGA7+t8AmKJpteUjwtgOVypHMqLmP/coUXnubmfPHaYrZe2C025BWffaAFwuEiYepCN899cQO
e85SEV0cxqkO71uDrdIiw97Q5M4aO8qeIfdsJckdMFmAKxLcdQU9FklQiiDJcO/CWl2peU8Vp3P9
JjpjwsZ1J8tgxho3Aoli5GQfZuzERLeb0jvfN9d23zWFY5TFgIx1cG+wBnOfa0ABzksX3nF6D43L
ba9hRu6AVmIaio3C5NoGksrZaTpLxE+73ZfXJry+dq0x+bKba0gZW2SDUowD2fG4KEhN6KZK15VT
ztfm8fUNPYeP73sp51M+5WuXCiWmlsR8rXiXPed/m5PsA9b2byeA4nvP2463AeVGJqbDbeC4owtv
o+UDkDV8lDwFOxJLFIm0fPcmaWFeFjBUAOUkFNQHI+VEtKStfIVPYLf2aacA7iJnZE4ouUkOkpGm
+5OKMbCX4wYvIH8yavoXzcpuzFH8x3CzopNVcNVyP7UT9Q+LWxhG1DfCRqYsXtRgG7PVcOvEu1A/
vttOvoFMRf3Fa6BmTFa5hBEnz7e4dqltkiYksX34M7Ams7dRH0ZlOrPdLLeEkVwrOBEM1G9J7iEX
cJnG8zd4sG/SbiZLQ2F4qzqjpIiw5oWiISppf2kgErBlceh7jD3AITibmuog/u6R6aH2205XtwSm
KrIFczX81WjIvBj4uGZJrW4nMveCVilHzXW4OQR3QgVAQfSBbYkOCNHWlmGjLoIRhbsrdnti89wW
f3hSmySgMNJYsxMF3lQ9r9NpFPJ6A6MkF8nIeLw+a778PzOyGVhFQCkEzbFseSBOQ0TOgZsY9Qhj
yaqR8HtUxDOu2wzwDCQIOZ5jT2OcrkzHho6P9ERa+tzirLilRRtH5i5A4qr52z7J11NgQmV1l3Mc
v5KPKBR4RJd2I1ufan2gwyDpWHQyKNA9FZuKXrpyJJf0amU9hvJ37AO3A2ALFlGSSH3pNnoxoGwl
sV7A3Gjl2N1nNzZaVQEJb2K80zsW8D52IIM8W/9aVFLtTpkqSKVdP45XlpKBButJRF0uQ0olj1XM
EaANTH88HsFRbAcP51MMy60W+B5I8ExlpT+gr5sKdq9VipWwkM9Hhh9z5B1+HGmsxuoxcVyGqd7r
k83fUxmOlpxBh61aOXqUdcOxuwUCwvb55CB2qafQeC+oJpsOqSSaRI4tKZsHmzxbLH+F1I04C4ba
/trkET5MDU4TquNgeSSGmPXN7FuWdtRkbPLP1atF9DdwUi5rn6ihj7KetqqEvOLv8wNmjHRDB3kr
l/8OJ3SxCxUxjlltRz8ekDM4i9FdrWcgm5UgPWwRz87pi3XXvil/Ojrvbt3ZVvWmjeB+cqvf+FTq
2OA8U/kjp0F37vIh7ECF4y1NGPotjQFHF1lCdJHo2Ak00IY01Q2SiOfvOyBRi7VkF1q0KuuIrspI
8MjAR1n85UHwuFR4LwSCXLZ/roUF/b1/cgU06MhebPQyhiBkW4U2Eb6oxnovzoU0K5515beOJbNc
y9EzRWSRXipcGD1uO5L2QVACDqj1sV7L4gzK7btN3ehl3B96TbyKE/NRoFznJYTaPQr6pVIirG2/
OWt0cb0dlfo6ZRt4Nm7nbXp4ldgZpPiQLVgWaaym/FIIptovZUjy4UKE75kfwOVR6QXYCw2xTrgr
P1rd1uboVvKMdUF/ViyVwFfKGg3wLdVlibcPYSeZeC4yQ7FfcaEhADjpjwLWVXSakpsU11SB6qnv
V8gfSzmu+d910jjOd2VKiVudUvnDrPkJ/j8Qh/9SAfKGFnohMdo3EwWvwCgZBrxiZqH9cpJPjfvh
NhY4nMekqCh0EAd82tyEftUxVQCC3A/YVhZZjPBiD2nlJBtsjUqc9T9pWkzSq+AxjCbE1KJ+btFw
9524CZtUZoZO2wx/QXmWoM0tsoR/yxEunaejRuMx2azfGtPo4Mk8JlopxQ9qLcsZYxeGBLFBalWm
0BGsVtmao3eQXETGy99JtOv9eNqhKDav1jIRJRcIr/WNoWErN5FcVmZF+JunkhFy4TEb01JdVq35
Tpxt52UAFP/UL2DOGQckxrm5dYJplnBH115TTdYehjHosu0FwDYbSM4DcBkArof7qTkqTQm5807N
xNyPjuYe8JjSabA2rmhfRnUAsefS83Q/CLGdDjg3F4Z00tojtKe1HsuOC7v9KcePWjfIsOGH/lb2
/Po+Mh/jCG5rOc+bCZzMS3CQD2lwiyQbIqpTGlBk/+zmQZH923KfSkfYGq/ecZReZNlO1px+dFhq
o6UeSSoVbQ65BBld+tN25zumhgYfxjSC1c8gkvC5DN5NEPajiG6O3M+LNztfauSupOH0ppiuegL/
xEvZjEzg/inekuYIt8+jje0lLC4Zps0qJZFP9BGhLSPYy4ChDau9zQDG4qQUElHtpyMdj1SYQ0U3
t10Bn/xMmn5+7ugBGzlfGvVRKsCf2QXDNijhxmxHSSKce2yzqM96AYSYD9IaoLEEohRXV4WR//qH
V2Yph3wE0AcYkl8kt8LLkU/QkKPyEOJ2vTTpijB28XjiPhR179ljxms5jNydRP9X6WfPr+EI4FpD
Cvck3PvLsNSF08dPiOs3T8lO95klGfXBc+5rXZZLbByDLDHf3duxoiuS23FVwRuWCqZmUm+pfGB5
rK966aRcKbGL2gukrA8DwJ0DTo0x81iSo0sIUNrDj/CrjKATRYCj86Wu8lBPkfrWJJ5wLZrx4Y3I
AJirSutqOIQwbYCTw5W8jxiwqGx7tFVBaWg0Nz3dFA/JyzY2g39oU68Z+N6hTxa4iHpzFXwvIvFs
YGdUgHdeJJscxKQjWfa3LKmgx9mi32frv0V8Hg/Ziy2/WH3l5v4HzJAbThkVKXrtsU+JR2KMvELw
/ZES4SkG9jbNE7f1WcsnxwTtpkb2OAdPpGjrCsqnbl56sKdx9O6GjQ7ju20PBDzCJSejWrbHWvG2
Op5B3AnM++1W3FKGecb+rBJuHIEhKPjtUJlW5mSy0K/2D3DLZuKqsfHl2495riEwIOOYJ3m0z3rK
sjIP9FQuQn/xKgp616nOPunZqkm47RkHIlLSgHNxki8Hjqn1/zex+x8cEt8+KD2Y6kSAmkpQUwJJ
zOdEN3ZnP2wYhJhRM0PaAhQ0BLY9mS5atwa8AWcT2AsRmAysAY6W7LCp/YtJ26JLgYilTvFnOVIW
0KoIgwYmGMd0J+qoVbfRyIHF9PI5W44QqV0LBqlqYPjBaLuvTfFMzRcvAN2X4RuHEB1WzPBNqfsx
1uIqVN9WO1m5nYbPrFT3FW4dxy7+7SMcGfr8GrzE7gTASJFRAPHPFO1vBJuv8njLXRkoEqQcC2+1
3FIc/1KmeLxOjL75hJTZZllgn2PuLY+mETKYxQxORYmWYwv2DlyCRiIdPYIeL311Nf6sY2fH1Ioo
9Nk5dFZPDC6t9oRwkvBzYSLH9ywH8vQCrRwL+lDlnfqAuzTTKl+G/qe9MA7egx4IqdnP9jIxFjzX
NSdCca3t6Xbf/vu1Q31ahl9d8Wdtb/qKoYxtisbnJvpK+nW3Nd+7XM4YIYFiDpf423UwZ76l/GN5
AW/QGEOy8NnGcANIQnaWAYnk7pCSSh+XCysWvAdcNzex+i5+AmpOt7P7CXB0Us4prHF1GqVQNHR0
NVBomSGq9uXnECGWbWjg4uJUUYWvBaSdwdjUmhpZ+sl37WVRmzKF0Z6XPUYPLtomsMvyMRsz9IZM
pjH/ChfrPeHkbfo15RSjls8JcttyP7xAj6IsHY5DGrscxc2rGdzRhdaAGEVVOV5SLOHuxu72CdYB
t207tSN4GTX3aV2CiWYGM48fXof93I7oIqPwVVqPBK6CsGvuBUN01AiQqtKyD7ue6taksGoCfkdJ
JgktHdbqWvL1SXN2wc2l41AEkzIUUKo0dBnrXlFoDFvj4mBvC28M5uDxzhr+AcC1VWHRv7DAJvVx
ZoUNa9T6Pdi0kHvbOyVj4ZvZmh7bUSzGJiEXgyrSpvbmL5LpLJoEwS3H2AUphRxrNnKwEnIPGdI9
CHwN+aWAVPk0sMCuZeRXjS16f7HCY/AZsrzrLH8+7T2YAbaWIFR2IAE0/gjSsOJZeelB3KnvZPnc
x9/Yu6AmazVgC2YGhnY44XIxgZ3z8gQahSjLNb0AI0+aNhzOW1zWZqJJVKPCZvPXnQd6gYvmBVde
8Os2wW8oMjZ9seByNN6P7XKUn/rKATwDdzIUK3lFnaRX8q55L2JyORr/Ckq3pL+x4sjIPKiWCBju
cUZTREAbHWdcKaiLxqGriamPY6S9fpiJdm3dV8iXcyBv31yTuZK/J2/nGVfJC/HrO0XAiAAtAIRI
f8e1qsntHRPZezTEbdAP9GUJ+y7PQZAcDnORoJBR+378qY9H5mtVNxISvSasz/ErGV7lAam6NTj0
mAs//YVkKON4Mq1PRbeFn7Bg4M5Am4pbkCR+Kl19Vo+QuB9AlJVAk+lyPQtutK1owHkJbRlDRzrX
s6Q2+rrMwuaZMH68ZS4b2X5ashT5rj7C6w2kRHfvB2dEV5adBBuHQD+hOx2EfSIf9ZAYavwmjwyG
XQRJsutibi8q3RaOubNodk8N8bFRsTNHjWYFwv2CMuszIl4dcZWvklRC81eVbSL1L/57m21pz06s
ubQ+g7I8FjR55SqO0Ww7Pn4pflxrmuPMMzHU9cfmBSaLa41YVwoKY5qNe9wbisQRo+VzBE//rHIW
al+eFT4O8TQizwsdWDzMuIZZa4WgMX9nE1h10v6tRgd5/QP6E+kkJjWjMd4rxcOlbFuJPV7dz3y+
VIOemJr/wh5eHbxgh51oSctuj+cy+VqMjmZiqOU2q2SNfaTN9udvGraWCryiuYycUCQ1V8c9K1E0
fDfSrpdmdZPkd/LwEgezKWdHw15XFoQ83+U3Psbo002H7cjEYQzw1iHmNbckLfpSz/iKr1Una2nb
opiGHME8xM9REHLWYUnLsOeuQ39e8z/3VAIfkv5iF3W+BOaAQfesEddPi627C6sgRVEiIX6EyT35
wAEKGGSspvESJ0pEo/J8uHPEn/bGtcbf0NuKU+9svj85KosTvrXxwisdr+HhrF+lnDTHqojFHKQK
W2vRf31dUPa2DlX3JR8OSoBjaaJ85TrOr76xYAhutEsPHIO61c7OIJqfeF6sPmn2o5bOc2HAfAqs
xSCoNXkJZIEFDTDhjNHw+CQNz3/ichqHN0aq1A2BRmHS+i4Iwh7aWl20WgwaQJZuUhFq1bFD7ytW
qiL5PS1ZzZu6R5Vfpi2SrIWshB6dPUd1aTk06JRWhISWABsv2Hjj453tVO4u6/QyEu6jyNZHcWUv
7QspvQSZ75TTQxzWE5h1YEilfSHJ9tbGZMkqJa98zxbD01hVlbrswAu6PH5lIbPYZakOogj/7AYs
fg7FBO8Lvk12vIVvHOCDgJxwRKIr/QSTuINOdhXhWDLJ0gEw2R04DYWYw6M+BLcb3dWXfAahn/Q9
nqe4Ix+MuhJG1xdLdiVIest+282dYmk+TRcQ3SCQwhWdiCAnmeRoV72cx3KPmiIuVs39BbBtH+Sf
eYYZ62yZF9p1voDaDxxkvrayt0Tzq8D9R8Wk4ywOtWIv22ZcBvbxh7KI9wOvw9JKRNyf9xKJ8ygE
z9e/aCZz6cpqOn9bDpSu4cFY1IEymWjpFONdpq+3fkD7E5QjDbk0J+3f3NB6LusY88LiHSIhHqNR
CLIeVo2GDZAUz+DicYs3x7LSNQWURUlow0KYvpk0RZmDiZUUbIWPBj1xAiEk0x8sS/GkiQnTiZXU
d9l8IDep8m1toa/NUoGRbrWrRmXz9/uIsiKk93gqz3IVluiNYZK6oX4fn/kV323WyiiE7LddjEvR
bvAZRckt4SI8TVq3uSguzZr+7UD93CzcPriFYfucVJAe8YsHO/zLR/0pLyFle1Ubggi8wtamLT+F
iWSitA3W4wlbDsl7lxXYRshJF2YpwlTAN/ugeg7nUezKBz4RcyVqpGYWogt4M2LWuTDgWr8tsj7M
t7zSty4BXt0rdrzRzDOecfjdMxzqwa5KwvR/15UB/XGfb0vTBFm9Kr5EVG13PjiHgT42k0K3CzDC
IHG6o2FTy0xh1WaD8bKS8WcisaMWKey6cTIly3DOLEvJm5ox/GBT3IFDQvCA6CK4R+NCqKKiibvZ
YT8+nwOxgBpNK784MZX7HFniCgjq9gyeZB6zxZcEqiadQKZcliSYQ8n6FA6oYgP5W7L9CzmmGyHP
5TTcROREsdF6EvyygXCnxn5gW9s+KgBb0QsmXBo0EFU2uy1OJyLSzq3Rv+SL8kGGNa0/1OhxIhxS
wU8qdCW8RdogtRtvFUC0lO2EZlrf1HfQzQADpT6QDlRZNGrT/F4UBggnEKI8lJaRpxW2OQ+5mF5X
MofdiksVA+IQ6Msb6XEXceyNec5FHcyxfIYWRPfntCwaEdBGgRUWFIqgyy+qybDKX5ECtPju4GLF
QPz75rqb48RjfIsvbQDx8FjVfkMDoRS8u40sfaeRGU3Ce86VdURPeZclSiS8qNwIojZD9DHiM+n+
28DdqElj/SPdcy1QHy6JH/37wWea4XkaCAt0LuUdINaKTacad+6sK/XEWftHJ+EmXal8x5WrBPNp
CSATtmlaJqyXJBS4ycj9W+FbYpjUB70M6b0IYLSoONRUV2Ps3X/wc/cIwIAZ5lQ74Ldo6WWXJMrL
TiH9gUIvDPRNih3UJxhfKh42MgncxHqO6FrmD+rF9c4NFK/Fl6J6wu1aD2l2XmnxINdNrOdidOWw
qy8JoBC+7dZco+p4ocptYGg0z9oSGPmhgpfoHIcZAV3hbRVfy/7H9iUk4Gew1+oIEv6fURmVZs0X
WVZhGjCucNGOr9dPj3y2cUihDTnLWJZG4j9t+zu6tVQcyNnsDlG/X03OKK8ku68BwCP6OuAc2aUd
rT391Mn0OFZNOrOB4y+dFgUuenGm+4WVZ9ZLn0C6iGlx0tOHnMq+eFW8oXFuFgfI3jB65mX4AUTf
7UgTS6n3XB59cqgbKq0B4Cj0FWWImyXs6COHMtUPncFbTMAg/+mx8KXAzjp0zpbdhoezit3wl5++
iNLYCs0XPt7HubRZa1+XET1z2G2unmDdpS9oHbE7XFRbWaxvDMRwwzz0+OLmnfMdiA7spUMXTHhH
ilsZnnSeMP3ShVCRMcQIc/LHyvyinZfnmv4pKc+4EgF40AqCf66CgWv0Bo1TVob//E+7TzDKDjZp
Oq5hAO6s9Xibe7uWy82TwtMfuvZQBNBq4ThvQinSIqyqO91F2QlQateKzUMwQAmbpAQHfRxrytk5
Ofl6o0QLAmF9UwFrgrFb7pPddemu+FeXZff9FjXzUT99FfLf86DezbrlISk6TO8BwRlBuTaVTdYS
UDhIP22iQUJcBsIVw5lJ8alXRtbEgGQoyE0MD4FIoKSjdrOkGHbF6ZB9gohYRLiTRkjQlvmD9uZK
6DFEKMdL33b1gwQj020CKWgqkXfcSaY/i47VkgugwLeclk7tdvWvHIipcesza0fshn336IOo4Rzf
APXpVrbJW3shwoT2Ma9kTAtuB74ZheFStsV0rLTJv2NJrc0A6Vi08S3X2PLZM/MPQaC0J5A5Sk/3
rOIRM4XLWO5N0ZUFLJ7HpHpGb7tOOy3Te0+m+oeVdmovzzCbiBAsG2avHDcy1H8zzr9qziaTY71o
YygPivzHlmbId44WIycm97HzOX6TPzSsmb5RnR9KIhCMrq8ZQ0nggpOsqZ0HLQMZCFSntgpQz/do
5oFVG4+IX4rgHmDj4YM4AqGv0K0XxIhoRzJW2s+5EYdGbqyXv5q9W+BmwTah91nKv5iwFz/8Zwka
IG1lJ5IUT6vdFbHk3bMH4rWyGpZ609c6fNN1sdfGSpYofQLrf74SKqTTSefH56we5lwp4g0ziKWS
G6TRNNinRPt85njDujOqFvJHfcAmWlW0su8OgYdAUU8PeIdEO6pD6IMTCQdh83SGv5jlQXejXPvj
hT0ZbW9Qgjbp80vNQKLEMUk+8A6cWm+B3IMOPy++Wm8zJTSVrf9WINEjU2xHiVjN9lORhmwnVFt3
ox5TVQJim8RzgLmXSHqzQcEhh3FHj4M8Y8HBeXZaaMHnq7j5LhWL3fdQfsAj88QzQMirqZ/6+uQp
7gXxE1Ns+4r/uFjaEfZi1uLEVbdvrBT99Pxtb5RHRufY640ASW9lCQVHfwOZ+DV2UXV17V+m9XSA
M9Y1NICj9j5czS1k+Vgj9pSS3ikC0fiY62Hj1xByxXY1+MHzGbzKfErGNfIMb6FET5JxWIC3c2CN
BKhjaEzxkFoh6YmA8rYu65/9W+Fjq8tkr6v7caLHhsq7ycYMRCKy/z+2bIcxByf4omFaIriEdjvc
boDOMaPr9WCbcQXElVIH1PfSN6zJKRykla4JPhpNCSgEVFqwpH4+l2wx4ZCxZPVncwW2RB9oRtQw
V3XkEfw4qy3awsCjcf4zUCR7yqcTuyLnZgK41nCfszjpAcAo2+1HPFYTHjTd8t4PyYZpsJm4AYA0
ZnTT40GM9/khC5eoPUCSGdfmUN8g7o5WNy05WTavcPEn4gyPwWXdiTvXF8+kbXp2gA8nQSh5Q7PU
NiDjGGc8njGkCLAQKjQPbucIoyo+Da3gLtl5FYEXyta8l9I+pZmw+uNz5cR2Hs3nJrvoXkGt6vXY
CR/QLe9jMqgNXX8grSiIDR8G/f7aSABx3s1eAYemwpveeNtytjzgDunoZwv3FsbO7521EsJAy9rC
/bCjfUjx39raAeKC5uPbkVV4IP7exsAp8Ey+3qGpxhIDu429io+i9Ton9KMC2vkYvytsiLHSJ+ZY
JKrx9FKVB5flYhJ7MSynjRn5bywUt3c7Rv0fd5LuC7ye6VME2hvt6LRgTEG2RRzxesB7czDgYkzX
R7zYoj/1k5kPGn2sBwBsJGV7hL/1ZQoOFAddnHA0shagg7wgE3FOqkvpikNa+6GfDJ4ffu2rGe9l
iwqXyulFe1pzG1Hdaujyu56CeBmGTQXlV0h/zUDChgQNEUKTazoZwm/RmAA4uc1Ymh6Y4AAohFYC
njWTy446ETFlDSBDM9AO8MStd1OpaguwNQSGBySOcLdPX7aq1hEZHThlxE43I+/X8YcM7go1nPty
SouNgOCrc2wWxQe9TAwEPgakN8kUVRWXvuRNLKAhPuPJlHGkuSKaDK1630X/E3X1X3nT5/qDdYui
jJQEkGxYuk4joWUDI/cgX+1/NM9HpeNVEvy184dw9B1GA/kCHoiMvNyCSMweaOeZqNlC2A7bkRpg
ZtcuJikC2B4DJSq1VjDCBv3Zuci9MC+1h1gGSrzJ3q+Ar5/qZBYEA3hJEU6slS3Ij5vwr0qDwvqG
1UIDyjjoYN3cQCcCtef/Fnb1+CsXRJSrguYJjoFIDHnj9aVu82bgKibPuWiJwUlByDlpXvNDjY8O
F2Y/1JeKDBFxLtDP+wfI/IskIJt2QvukCG0VW4lUlODYfkci1ZYwuQACVftxEbZu4RVXZKlfEDQr
uvjU0CBiiUxIw2iKP/6xtdVckUXJmV+mP3pkxVbd9/QagqBe4SZF8keSkwLdkob1C/8dsxkBYrvC
QzRVhjqsGK+x98caCSziSB6yxm/nZJCfyqUgh6Jw6YyMW6mgCNMD5mBQoF6iQXYDziXxnFREO/G4
ZHknXJnY0cCw+kUCLktWTb/1cUOWYnPYMCh0gCEY4iQ+uuAB4QduSfUUB86ob1oSXetA93U96bjE
YloNFJWUsHB54cX6SomG0okJwdpmfeFtQW8Jkn25UncAJ/Qgm/lnARCGy8Jix3PPExFJG/Ox3JRb
DTzynkRvJFjolKAWDSm0hFhdDMMgfL6Z1ZiuYUDaVEATOo/6U7usm4wjHtPB5AqlvQf4hsi9EIcy
vZW0Zs0Gvkh8Hfx8bVQWlaZdX/zzjLZdz9LpPrHH122ykZaRfYOAn0PUJ3ZB3F3PEPphZG6z+T0n
rW5hfRU8ySEPbIJIUsTFajjRJpRDtv3AFv3zLnZjgOkTLIm7OlR2wcFqI5eqNwnutChScLTKYm67
4cr8sLaNZJHQfXXKGk9RN4foG62kWycU940MUd44b8ma6aQEqjyufRoOA8iDlpZegCqr//0yjlqi
r2kFcABvoUlx/rIlDOC5pJ/OP6i4Iv/X6ZSV9Fyvhb6OyY0fxgj3B2Dm8WPapKSI8DCivr8jKPMr
RTGfJhImftrh7fC/fibNq9SiDgeRD0tvCI0lrphfnoAYlZbPVaIehpRmj/GtXU1jHF8MxLJFdM3F
fmF+6tXt9ssfjWyE2h+rJsGnMOx7WE22QgejhNKRA6sBY0jwJ/C/88AX5ox+ihV7bvXJYIZvd3aE
6s04on5Ee11mYP1sDzulwYMbW4q1O7q+V5dtVBhLrsbceO1+5MMwmWHjfCodJoQUkySTgTdsoHpM
7Z1T0UaaPN1R7XrrXIQX80j71EYRuLTwDw9PPWObdzSqVk7gUwGx92O84kg8bPmK5REsH9v3oM3k
pXrS3y6ZwPRcimh4ktHkd5IAa7+4AXotdHev8UcGqPNIdsPcQ9a8zwQsAvKx2O5CliDtyZw28bRJ
uRG8eVQKpsyHfOZcOKLKJeC3Ak8HzHjMuYh871EjM8MaMcoIxARjdsskicrOmlmpbVBO2PCZ4Tl3
IrTimIah7LzSGI32zhAAU56c0xMuiNZUNHccXkIe3MlHR1g3zIkKgvnNR9CIHAcBIBFA8ZhL/q60
ogauFixsBiNtqlyyHw5kkAFR16/wMmocpW7A7oBlYBffWpFwpzkBwIE5jzbEHPRvNI8eSk1H9RWc
D0TCbdUjmEkZWLszfmxcN3th+0zgpLxbwu5LMZxf8r49aGAhDmhJmSS5lAj6/uGoninrBgo3W78O
s/y+EOKOY6Ep6bmfBRSpmVSpJK4BppHIZB/79JabyYpYN/W7tfHX5vj5Tw7/ox+CGd+oGiM7NAsL
Oz0JX6QYpmta3Rr9FnO7snOSjl8PbtwWIHTsD5GQoFKp9MyMNlV4H86j7twNUv9H8n1b2wkJ44MO
wMQseaaecRa2zw3vRpRDc61kKhjceVumkQbUY9pJP4ntKQB5Q0szcn/ayHdDAyVCar2PNRs/Uex2
18c5g3PQvLRF4y0Q/v/u1tOFDw5A7W13uf07mPSGh7psFLXaa8KUmSSXk+c/EJt7x/JOxXpfN6vw
3o0Lq9UPjD3cmsrAMDI4zxis0LDBdHBsndAgMvnsF4AHPCSyK+8KAYf1iUkcynJaZf+GlJNXd/Cp
/uaG+HTirWsWUCcI/usEI5UH2NOWgHkz6Bhgh77NIaRZVyQsW81JuMS38gojyFuHvO2B0519lmnw
vpNVy3CKxh1J6/ErDBedRLEj5lJZ/L//WsePOs2XzZuxPsi0omRFyWbb1Hz8+Whw8yxc3kU4BeJ3
piLcHDbA9+6aePyfGzBGzqWwIQNO3EOmz2KBI66eh0eICBX9vZ8dUefoNXCOzumPSN5K8d7tsd5+
LwwO7r+1dphT9ZXrl3SBo9EnxXFEBZ+s3RcZUumlJNyX/opoLX0zru4gqCPbca4Ra0z+iSUQH123
LtwTJx61jnm+RcnVE93eWlvoKs6HC/sFA3ahgBxHYO7eNr3+az3azlv40OYK0Q+/pu5sFvglU/4f
pIV1qe0xoxpX1gXGRdjQLIE5X+1Dab//ORPQCumMkGqKXHfOGeX+AaSaEkccxE7gqLtNg81uexEr
nGCuE+xxZnf6gtECa0K5TJ5vXz6bjrFJkXBo58w2tSwApXhshyZZMxx/JdsNdZXz8XyEhFMEeHRO
BP8hJUhyWvIqkGT8YFct+4C9P+Jp5O91OTAFVmHovwm1c8bu2b36+Zx5c7UCaQp2UGEmBoUS6kb2
FYQwV8brUrzXopMurq4M+e86ikf31zAyMXwa/HAxQUWShnPbBH75y7CLNlS2hTN14TKPkimkmaKW
WFtp77wTNnBLPMh+aG3yBLP4q6MSY3Wbq3gxONmeJ2pd08DusRDLi0GkVRzm83GkCsNZ515paKZY
qy56MZMek9/+7xD6LO01EDb25nBSciSnuTNWgO68JgGL+sKHCPcS+BjwNa+elUmbrx5T1iDUvyN7
BxpYyIh5wh7NBsH5hZt0Zx54/BLdUPwfHPxrWYnuzJ/Y7D+L8YsY3wtP6x8OxhBCRll/mX5II43h
/PtltccYNel/lW4zEOShZVbcz092LO6+xdqDdoNygXtVJZDjaqj1EEtM/bXBhKAkGfMnGlo5sUzG
OpUYxJBczENq4bD48gt3j+1Yp3NAYhiNFQVnPs62aUWnbb1DEB+tsQpy0zDB7RXNq5bE27JuT+0P
w6GZpHyjE9VG0F/yAVzMC+RC1HDRmGcjd4MW7Kn/3eW2pGVqWFZH/df8ooRRjLLR8n9xlEILUL3p
40JAsSyVQGE4VaVUHLRBhUTFIBLgCRYm37Uerfeb5LiGW8q+nYOAFYOf9C8yqoyGeKyG1VxArQ3C
bLEjg0aiir6vvQV9UP4mqlhEiYaWTHdifbg0Fuo5bVvl7ya7/u50Op4+7iFuerMfbBpLw32bpO1Q
wl3/V0iB2F5tY0VDLj6DTY0IvS0jtUDNZCCw0J0RRT30k8oa8HskuuBz/CEq7SeKpz+fxuZohVlK
lq+78hXpTeHveruYFcxqIojcxC/DuU7FVpGCy+/14pODJKM0PkrCWCRivXsqSDZV/HAeGkgpqKwQ
sfUNtwxiKPPQ+7D4xgWTUgj8zTpY72NVd2wxOdF47gv/SygCCGUNwlmFQtVtqnH2JHJgB1Esn5Ps
BBONBwsPqIZWBorZ6o5dFzS3AvYDA2m4ZNN3C3Q/x0kaK8LALRs1BQ2/AbjtmpiXdukdPpk+5uFL
bLx+P6ptkkjgu/MUvRbOwUZ/kVGpuUAlFsGUzSvcAEWjIT7VqQq3OYG0gwopbojPdzMVIITZdglN
76WCV+EvQ5qs0ofMoDIqkxJuDZgLZlyUHWZB/uuOExWTKtlrz/h95YyT3eWXCPHLTyhnHOjNZEjt
NPXmn1Fh+QqkJ7aeNGT7SV+FMCUOcN5xua5ITCnkNZ9gC4czklfsmZGwZ0D/7e2Uy5OSG2vRmZTg
btmCgUWbP2kJKDizagOSSvKH5NMpOpoeodv3/nYhVDmp1QCChB9EX3qxPuSj4cVU01sfLn4aL/Up
f1Vw+FdBfvJA05mw5awaIvAVwHGxbyXlOSArR3e2Ag08HfV4+C0wSp69PlPOCW5pss+Rwe/nhwU8
xOlB5vfGkdKDJvLiz9f4YyiBfpSduC07G9qK5IRoB+YfgT+9NphHzm2VjZHDZtiuN7CF6df+t/XE
tCbD8zE5kZ34UerNVHGzevveaLrckrnFuah+GHTsGxgYno8F7qgacFWePfnh0pZHSX9rMDIABr6l
uz5MGt2+MWjhstHis/4mcQv2hdsRjdJla/cx+s8/UtIProqHC0CADefEFQ8RfBwb+43IWcF+ZTfg
SyJvsNgNw5CWwB/qZRDnDtD/laOj/hyUeUcAV1Hw7bfyeCt+iGsGhHMidGKGrb/BPi100QYDs2ps
p76CRWfwCWPjTRBR+9+jgAwttfvg439o7vfNfKlRMDNCvRvfmopiBOZnv8zmM3tZV3HZ6zCRjuqv
b1pSUcWgIkthCHV2OthX57cegUzk66qEtr9411GJWDA0gr31ygpKymdejS1UoB9ikHUxd7nBUAlh
Otwg/ZmdVqAQHXwGG67jRnXFkb2M6dmfSPEJvC0ACNm1+1J25bUKsRLyfDmfp7e6PHr3JWmRAd08
Q4Fc2fiqORZU0shRCLMeEdcFlt9VmyAJk2R4zxiG0Dsi7NQXg2m2TxQ+PGTH1OClWTfuYbPwp3/p
gG3GNY8Uxie/si6I1ahsY9jgW4ZH+GaeKjFHHVsjj0UHC1wfgpwBjzarNn0KVh78QTvK94vpj6+L
btVg5OCFCHbIJW6qJ1ApsZ2lqj4Vxck/6y1XwLrWvfQLM3+DhbD8TlxTuw0dajyvpp6FkA1GJvBK
VdA70IPVZ/9aW4YjbYDdWI9qFwKy6zD46ovEXDZ4H/iDyshdquIrr7GcpMkeyvgNYa0/0kgIrHdH
wnpl42jl2vmX9guD9kq35XBOWfewtvtcg45CA/iY3bebLXNjPHOiQ8MUtZp+n5xu8PsUPHW33JAQ
lYDZ7fHT4NKvrx+2oyoGT/fGF9/Yy7WSROFIlgcZVqdWA39CfgAVkd3B/Cjlnffvi1NWPX1MKzMo
KY7ZE9ZCjDBx3mJBfthzFwxq5Y6o1wJsbLKwJP5p+E31LjLQXavR0+69wy8zh6v10AB0GLsqeQDr
ELCcy+WV7UghNV9DMshwTAQiBL+ax09lHplvYzH+EVtVVqI9PircLJXaeaDXFjT8qYFCNO/uFXgC
y8fgju0UPi4WucUGvmgzRE2y4WgGSG8dGUHOf6cWfGjOr/pckQBUciVrpKAemfRXQ6OSLJc4/v93
YiZumYztXUN+Z8cllSlYyU7xsKw07SrAoNQ5Zw9f28CJw3qSxq+wlv5IQ5rnWsoTpPr5DiZMl8Jz
3L3+sYKKqgaI3jwfXQS56BJzFJomJ/hMKSrIyQS6vra6B3rJoeB4Bc8IYOjTxzZVy3fy2zNUOonp
M6xP2uf3G53jcT8MI2uORegU5hR0sD2BlbExypxJUMlfz0n0oTKEITvY864ItHFCQ6daJa1+Mwz2
Q8SvuhHQPGz2PQdfu2hITOwmdrvvIkfN26c35Au0RjzV0jsWEOqT7PquaSzj1V0UPW9AOG0Gg/1D
DTIYYOfz6W88kCC6kbvy5MeW5bz9mSJTp8I+E45hH3hFWu/aLwR89dKlq2Fqr4n9G+/E+UjJ4Enj
aETpiJz5pHs13t98xJjQfL/9j2EuoB+MgQpQodvnWkr8JWak4NOUE8EPv0qU1jrqbhtLvFjacyRe
wLkIC0ogjxi2xIHAErzMLwPbmCKO86I9fbSMIoN1VMsndncZpkriOCA5f9b75eGheOQL0Ix3fXv3
hK3u46d737qTdpF/Olpr5um//jk39LilP0ZQfjFNWlt1PL6Aro413UGNvJ59xyF32vJy4dlxmgSU
D2KwnYh3ysAFyA9P4YykeUbg/54dFa1IPr3HTja317v22BIpUv5hR3JCdp2sxigJHQlYbQN330nn
RQJzR5JawMRyZlnmXIWjq3lZNlxdgQND3IYasd9th1tdv1WVRfZKYl9LqMg5K5dPtXnDlUZBXYPw
g8C5B0dfbQiYDdIGPhLQAublYdQmWv9zqWnpd0+3iCebmopKNdJiv5UDz7wO9kH1OZoIiWKsgJeW
Dd8Wz+0UTXn234X1e5CXuxpzx3hBHljE38C3WH4U8OM1nVwN/iXHZxEfEXyQhdtfi/Zkw84e4a82
hta8IfbDNsmPYS6BtSfhGpEdfpEL/zynbGN3R/H8OzfFe3N14YI55qkgzK4i00gF3sMYV43DwpTg
UnO91atB4wT4YaAwSn8og0jDrvXYhDY30Q2Q/3GNL5/mfDBbL0fGVNq+rhPhf/roViRS/fWXNG8J
L7HR1gi0JJzmauZXs1/32MZ11IslYQR4fSOKOWUrU48Qo0P7aqLT8AQhstTyD9lsnKXZlPu+xkL2
aH9M2dWN7UuMcphD8izjkzkFLXIrKcRex1cWO4zWdctplTayfslnvOdUAVLOFCQc7ZuA80t915Gr
sKw/5TI0xPmyu5UbpgLiWvFuTZq+WXeBlEaH2wsxXSIBE9lzK+1+qDpKXDcWS59wJgJe9vD0vojw
0ipX3DZ0Undwgh2P8hSLkFmhKefBagpbynW0Q6aaHCUP2P82ep+Yw9EkITJMm69DfzlPPntaE9Rh
OMf1UATqc8GnNR7VGQkHk8HdsomPjAIPudyu+en+0aYXzRZF1AAyENisdOebLy3VGs1JpxCKsACU
NU0UwW7gtRteTBKIraszER1HT12sNQ5hdvle3VHyRgBIwj6KVGPd3DCt6//cnit8JVtGmbxXqqM6
7NpOT4vVwtT5AFaES3oztvoc7HK/ufkv+9WoRSr4HV9qdWecdf2aWTXeZQqWclR9vmtpan0wh7ak
kRM99oWR3L277R9wcpZ21rvi7snOE54W6q9VtI8fzlQ8k1sK7qCD9wNXciZuQXehXdlLk7O+Jro6
+oHBTMjisapzJ3iWRG4mkA7+VMjVuWzib4vM5lWmijOwjZEWWFEkN1RAndHLJ+VkQBUry1dZ2EKR
K5DWdOcPpdLKG/0vCCudnrEVC2xGFf9sU3TNmGr7OKW9CytwIfHIGl0G260Z6yfzL5fgIH1KqcS5
CnszcPGsZm+xNRviU1MG5b0TIBQxxoYzOI3TBJicaoUiglW9JY1iQymczy8cSn29il3UrtveGOsD
yJ+AB7UuI+QR6KMIitxAn6kEQIU/e391vLoFtFv/H5RM1Z8ApHxcZaME1T+QpTPnSQBjApgTE5B3
NnJ9mSzI2xBddL8DuB9IPC2hNDPl7W/oiIE/B9cMw99qTnV3AlZf5B/t/gGD676U85LSFzCTpPso
7grRJE2S1XWn3paz09eZH4hmB16UP+cBbUHq7Qj8jzECoQjhScLNAtqjy4zh3+PqQbid/ixQkstz
hRzXWDzKOA3DO2zQ08ow3IeBlcYIHYPShy7Rj9I0Nu4hDYC9eFvnevkm1TdmPTmuP7T8EZ5LjjRK
UlxsIP/fq7JwO5IU0hblTqpqdhDlHk+0sJ+3nx/1PBhtO8vB0aOAh86pWDDrEAf+tilj3JkyW+qN
snXQr8kKDUNV3Usgv4kcy9xI4v3ilHPiEX4q18PookCEbsPRWghZXKGLVag1Fax9k6T9/qcwd74Q
/dhzYm++tu0zUeeLvAOF4VJGNAliOJk04BV3MhrfLNvIurpaw73cWfknq0ysobq0uCjRnzgkX+Yp
vp+Kjm6SKzWAD87MkUlK72+K8Ae5AvSTvJqnXo73pLYGkujLAHRFvAZ/vie0GQJuATnVLUJPb/Nq
67CpCQq0UqlsGmj+2OCxApk5ZoyQBTa62cKj6lkjaNP9SnxVdbnrhJr5xEP65wn9YnBUIJUR5Kr7
c2C9lQg3p522y9Q9Ar4tpZdKngaoJWbTxhwnDOYZWD30YqufW28FX0Gix/nVfHQiMFEvGMRoEFiE
ME4pKVIpQoCjcmydc245cfdZE6A4at1BwZjodSNWzyl9wSzlVDgUi4bMOG/wVlQwIb55hu4Hk7CC
9t8MgU7S4FRSkLn+5IV9rDQnJDOTmBERiesn1ZaauvmADSKaecEdRx8C5N30Vg/my7mommel1LHL
JiqCfhSjMK009KPPqW2j+lkThJ7i3igiBmsDq0cOVAP6tigoNh7dPFtxEKweHmUFr+UXRV/BsVkH
5Kuhx2VXdSGk9M8RO5o5qof7YUnsGkoy/Ngvtvq9JbsUVU1TTN8cEIyZEDOVbe8IgKEV+2dx0vzY
ivvEjPbIUzj/AmkR8eAlRGp1M45Cipy8HTdrZXkrDAXo3CbntMvz4sUP+BMbXVhyiQrxklVp8QOC
ANffp6dO3QRGEnB/BebCgFpq2j+4r8Nv3D7zL4+gAr3ruWAQHhCJl8crMb7YE23s59x8QDj9Z1vs
xOUHBsqBEYlG33oHWOKwWFzefLXvyxNEF/k/6VLi1aE+ejwvDmV0N26MQtBJ3mwuoTf2zWHUspXD
/LM4TFqLboNm+ZsrSsb8j8UqPP5Rni/NUPoqWxyZyCnTi/7KMgX5687zWmpTrMEsZ5xl8ygJRfPd
HYrs8D2MnU3SkGoShyBxm3hmfLzJqWLs7eqlTfwQQNhzdeD5ObBAw8/b2U/T53fE9O1ED9BDQDa0
AlkEVrwf1JTb6Yx5FlXekPgUuE1fQhD+oLxukzj3CwjRAbmRxCF8gJSrq6siepA4uzyi2RFLH12c
1WU2pLtdgBMIudVTH65YBsuzy7tzwzWOe6WzTaFyL/yb3KyYbOSf6M9Bu+rl/p3aNDzW7EB0vukJ
hV+udp+oUosJ0d0PaL9RzxcCx5L1F7TcoA3QLMXkOLl8ZQLxZB9XZjzTkI9F9vo17JmYKEzRRHDd
ycAd+vmLPmqtODudSsSWGLDmYb/f8okcU8kpykzu+a6T5XOtNoqlX6QWlbtvjN6rgTqrjOYakbAF
XQqOM/OGZ209nOX5uHRjaaznZuJRa9boE+dI1YtCUGRg4K2MROBULHm6EERgMYLYeT7H1LWalYEy
EDuMT+LtWzvQLNWpPxhfYLCfHPi5WOmDCAqEeuHLRG0UmwXIhqs+WYVQ0pIJy6j2pn5a3IQtbqWR
JGEN/g7eKrXjONXo5hADP+OGTRU8tVhAD6JC7pjzvx/vxLebJNqBrdPXspKthG14Xkb7dMSD4iD2
V0dVxJQlUvqcBP8f4fuu0OgXkk6gDrIf5b2HD0vDSzdKfVGYD7+5oeYN7kPP3FzGLImi+M3F4CGP
DQysq1gC9LvWLWUqfxIiFVehAuuW8vfNuJbFlKIOMEo937T5kleEbRs1B4Nc11P4YS5ce/DfXIH0
fUqTpuqrkmc/RZeGIl/jx85VQ7a7a0gjo1joCHp4N1ElzBS3VpBMiO5VB1BuxU8Bd2uo9GlefaR+
2/4V/LTIYMl1sOgQjladnUgL837YOJS7/T2AkuP0WxPT5bp+vZn1sOcW+PiIQoNfg8Fj+zel2VZb
m5icIs37BO/LLeEBRKkYGf1YfXTSWnK6AluXQS7VHuJq8VWSxexJBJpBIcPd4CYfaF9nIZdrggg9
Gk4EZzgwflUg4GV/ZF/A3F8/Vtu/mJsy/ktz+cP0E08hw4oTKG47ofcXfIhY7GHXYMWhX5baiBzI
s8KqJ1R8wMoEe345qyEPti530pBRQ9b7Pxv32vFUtK3tz2tqv/a2WOYV8hWC3r4jKraDBdAY2qYr
wELWHiqULMwvH1UF4+ZDl06DfkDmFHkIS+S5BvurnwbsQsFtxxbpX9Sd++Hw1PnOuGy7osIt78r6
/30RDMnSWXNhCq1bZVFFHosB9s+EbZv+el878IsYswad/9fRtFa0XHUs9m3RtWrp1iAoeMUJ3sPt
0IkaAozdnkVOauOtn9LDvbtQ6t8/wj1+2JKqMY9uJH1fiQLn5uhkQO5lIptrUcezaSzi8UVqxA3p
7dy8UHazCOaYNHxMH0zaZCm4buH7i1/Pc/IX4UpGfatvF7s6f4uyeWa7lWZY22Ae7x5nieufgnBt
ahqUVqUqO+MrlBQVsTYbDl8E1TBj09TN9KZv53rtYk/z+9jnpr77wo25eZEYL4hL/6IMzcP8ehDB
ozEPgr/GyvP6oO5ClrENmJ6x3Nm0tRpGoZKJIo1RUqoC+pLHGO7cua4+vhQ3x3qJ7nGpgOPTmbS0
U4g1nxhofXqYFpW1YNrkynRu+4WcirubstTjZlseyr7Us3sjRJ6ma365vTN781JtryX6gSTdBjzY
j2kv2qn65Z4xksfMFSCnckuyiuMOKvz4GFtZtuEHipC1UzXqxQsgYCimtz5jN1t8c976mpJPL0wT
WLyGYSU/01Kf2cCzH5wbLt7jTszGf547DXLWDhcNQL4qMoWn8VvUAVmKQ2Nt6s43cCZA3CrlKxVH
meLByMt6E6Q1W/I1ZTYOng9Xl9Yx2EhB1xHX85tqc27h1NqHpBdmnt3xq13UKKZQV78zJubuu9Ed
0k1/0BXZagoo7tar3bRRnciUfD2A/SSPCeYsfl7WXhxAe3Hbjl4RKWlkFJYonY/Z6Pb06OiNB6Rr
lgXr1PL99u7zaiteVsCvdt+5rt2LlDUjnWcheAC6C1j21YcbmXHKXMPUIr0JHGF8AVP1uQDu+fC/
8uXMBe3TWPbUg1SVbJK0XhWQlJ9RguXymXyzb5tcm14vwjVXDeOSnssAOaWBWADk38rkpjsKJHkv
cIohs7891w4UyLKzQEwfJSe7HO3OH52fWV3eYPcC1eNUKgq64+AnpyMDcCiRQNJKzuQzPJuTOCUt
ax/vG6Ylx1DdzrQfpQ9+BeMqFGgJeul6kt7bGP1pDOkTl8FIQx1/dsEnfr1mF+iQki7PkxMxL45Q
rGWsOGnfrh3N8JPqWzI71Sx0CW1ISEPrW4y/ZXNSUakTGfj7R51K8pVurO9VIm4XRuwxaSWpxXZb
qjrrt+np56ctfFmlrcRUW5U0fhc5HAjNABteEm/HXw8xxTE2Ze8DeHYkT8HJb/Nu3bqHcUTMaE24
cyYeyLy/8CRAKCxKbgQl5knk/dIbNiTTNEhvtlHcMzA66E84hrxWPLqEEqWbkDxTaDtx1tmytmgJ
h69MCriz1HSKkYCyXZ6mtn0olaQNedZk5rFFTBl3wpwZEuCNcxIgsAJaQIdCTokYtkpuVWoD1Em/
cDPjbk3Fngd02sK8PoDD/i2uSJDCDtKt0FeZc77xY2Lm/0cQcG4ltutTdd29BJF4Wz2nT8lXEqVF
s8dOaniXDVy3EU3FeEtXlaaDYci0Lv45u15Fi00OGYanx8xsVr+UcNQYmDrY5uJIUC5nM7BY28+k
ZkKciOPkXfjG+d6RwTTOflI09BFybzg5lytfLV3Tb7hQMrbPq3MdWzL9VzSb4F9bHEIxIh9M8y8b
L+e0SAzYwgntJEkczJlze9pcSocrxKx0DAZ3EmFXQxck2s6uFK17KD2nSXDk2wcgz8jFvgoaMvEF
zUgIj9YRZzIOVFZceNLl2WWRh7rVo8shI3e/Mumi8IwocWuKu11ImB4UEf+ZfiP4PmsMGbCqxmz0
fCN6jcnqXQVt+PDLlVRvydIOqJoAdidvDGqR0m94fUMOzFGjfUdgLqoERRZLZ8/dEP6pq2Sh9mt9
ULOE1zHsdLvn3xjnhMR0gGC0d5YcxjgwPyD0ROxB2DEIaCjXQnDeCBxlF4p/9yWyk/LOhRPli46X
7+16IIR5hwnlG+MJHk6dqWGzu4Ee9mN72KAZHsnOHu2zJ7sQq2unPIgmqfL7rdyH5tlCDW6MIu0S
4gU44gPdDOHiOOaXnLxcV6XoUPBBP+rAPZHz4gzQhJFGVk4BSVshQy9Ou6j2bDwa4BW8/ti7p/GM
Lavx4UGJcs65P+1Xprxgc7J6EZ5Y69DxK5Xz5B8Qf4OAAY+fUddvxbe7cQ3aLBWY7ksQUuv2P4mb
vy7xBrG2eRol3z2oYt5Txng9ni/VIy+DUEXyGgV36UVbVkFW96OqjWUZGv+3Q2j1O2tHbpPgj4YP
3yRKbA8u2msvuOEyXRx9xz6EbhKcBOEuuN1tlCWwAIPTkIOjCAKrTyheRJdFlzHXcclhFi77fVqY
Uo3PwN0CeIW/mGchf8/Pv6lcV7MKFIIBlKzoEy8iuhihy4RhEPO7vjn0WjfoO11Out/m9RjiMonX
J5Ff8AZbymSK/hGCBJ5qDobyz8r022tUrsCRWffQv9Y/0a7Puny1AClaVFTKAduddk0btccocas5
DS3P8WwaYjhKBMJcD5fiZjpm0qAGATCBHI8o5E1lNb7xcfGH7WWFnM4GITZ8rwEppy6PBt58Es3b
MJAUBV3UnTxEpwuh67VEyStFOujzW/18MK/bgMDtVbiBgmX4h+eWK9wZ88BQX2hpitAdsFfZpKSd
BIgdL4dFuETEPP8HaFMYHgn5de1j7sCd9U/8B4PwvOVmFyWMPgm6VMc4Yv9Dc2qTFHlJ8pWtldtK
iLcRNf/5x4EDiuxdOF1mtT1+M3VChZMKxM1RG24QAbksbNdhIzHUxgpdZNUV4FX8OjkiVYYYNrBL
O7HJN7djJq7irmYbGK9gZY5ObQdXY8pKyq/9ulQ5oHZVXdsR0JcodsDFicNi7hRnTypKlDaNcoqJ
FzOsoYYhIaKLnrBKi9ZQMT87srxD5K0F3zSiXFWcGGaRZwCqaJcxm0ThwkVJjpCtPwacM1DtnD/0
uYEusiRaYIikQy9MlguTg2ZtCkpLHhTFjwJ4vSLohOftmqVI0S/KLEFs31EULkLo0wmRsy03obNd
qX4RMhBmz7/dkaUxegx7Id8JikD3j96/cVbifcImnhYn91k+JYMAGOLg2OFc3v1T7HrAvzbJaLkC
noX9WILOeo34d//NFy5EBxpfj7fnBcoeHwRJi7sUYVje4rdXygwvD/bdNMLaOrzGIyFqhOYD1VqO
d9k8IvZsgtAcA4cfevbGAd5fQmr+lyGKIm4lbF/yyzV86bfRhVvSpFRJKk/IxTLX7Xp/WNJtfBIC
LIoLcA0Obvx1lpERgplE/PFB15E3Rscj+gHJxHt9wrSufI5cIhQ4cj6rKh+4RwTMiLx95af3fHCN
xp20Zmuce8F63Z7Ei2HGOnu+3ItwGvVCz+yEdKAosG96bsATbO/K3UTvaI4ojZUqXO0zYz38+Dp1
9sJfLyynTWG+cnw2Kkx0zevSX1iiZsePUQZyyxvKT0Vn1zi7fpt8X47Ol9s9M2C3xOilYJzqPiOf
z0j3xamuPdbfPQOuzJ/c4gXod7isla0hqmjU/SAKBWY0h/auDDrmwpaJ7C6owVB0xempwItD9bJ4
AteqMTcqcxRSAcD3nlOpECDYCblHudDpSIYXqR3FDeF5K02/izXJYsZdPlVRBh66JR96vstE9lWo
8VEvvzqsd19R7QbnHMK11ey7VMvu8/pexsD9h4mTzL1SyMVl16EJQ7oL2A3Us933+6CwMzk+8Vyw
FBAo14Hx3W/oa81nUsCmMut0vPLfwPzdLN6ZPPtle4+o1klHZjRlxb/qCqH6zRo6thrqxM4373Dk
hAT56nEe4Nl+h5Rrk6/RW0Z0QGabzcQz6bHLoZ7pYwsQ2mnFKmq1/+PmU6SN5UTHUiszPH1sSku+
KSIqa6HP/Zn5GuRxYD+FGX00UBCE4OjXyXWikhLB5INFzQvmZLOxyf2wcmeer+5tqsL7vWRMWeDx
mEBoHeH8+UBJVIdy98MIE3WcKc+A9xxTeFjqHu3WmVJvFBacnJzsBRj1VHhdNrxzxrsZu/wqEecw
Q6PNk/a5pFaE+CuVNoN98/MJBvJTkpIYGSLb/W4s7Gv8DVbNeyksuasGKhVCwR6CXGsoqdc/Fcn/
f3bf4xpygT3tY2QTEQfscNvpZact15Tb7GM7yDgoRTREKSM18mOKcKQUg7OmefFIWzP4GrPWkOIs
wUnlKJ6yXvGJf7Qc1no8HeK9VBTym8S+NLiVvO05ZHlNItEkht1e6L3oul/l6tOAkfW6nNfohNvV
8tbYEf9jXs1xM08tJLXGBrk/79G2g/hF5q6Gi0WI8w/qix965B4qycNuJdqpxU3ghXPvHlzDkCWb
4lR9D37T3gKa/5vpOvAaryaZdgTSzMPUPmB6kZNfmuOkfFv2sqJAu8BTSYH8X7PbaSWLPVEo6bKy
LFawGgUT2m6M6nsgxaHZsTzmQtP1dJ5MBDRP9LnHR+yb2y+jBAsOBhfAnGd2oBQbMMKaoPxXC6nZ
UGd2P7gFvIhivTrt3Ag+XyfqqCI6ExSVHFTOjZOGzihf30Vy8O5UcQHxgbqnwKJaXw+vjVeSOQ0y
+3OlKNsc3Q9rur2BzQdtzyOWRG5GwHDHKCnBTy0QpzmW73MFfh9UFXfyLJZii6S8ADj/TQzGBq6Y
vvxVozr0FxgBPhYsX6l3TX1Z/IIN/k3ojPqJbQzrqnvH+71tt0KzH3AKJ2Y38spumErcrUBK4Sl2
pQWTtSdy92yritToITSwgaod4qLDiyNv7MITVS0onQpC1b/64oeKzHpYT++ONeYOKbPZDZVUIUe6
Qcu12/ghzaQ1DdUjyyFHIHDWMvBKh+ix8IvspWcufy4LM+8UTXNbPYMIoEjdDneintKhaZsRdIz9
jkgx+O/19BeHLl4ggoQNsA1Bh1Krmps5BFZSNLIspE1hp4G2fPp4lkRkyPFSi7vM49ijS4Eji910
M06cLYIc29X90n0ChXNJRv8Ao1p9H8afdrYdGsIIWx/0QAq3sOrzTmGManWGPihyHBIaEcIbwjgV
UcSZO46AAAQO983iqCJFmSQFLyDb7O46hbjwRIvPwjrnhfrvCF7tA6/EmMg9JQjbQcOjmST57hhf
YaRz0JqPL0ikPAbeMHDhMZzCbf4Fn6Yni6gdUgixoCqccMoB8LfY9tY2hFpZiNje7H/GEt6ubewe
jsHUhMIHEeeSB3qK+jaXu24h3u04B0Maa+/vM5aLEpH2Fges+/wQe65EKGq1V1kwvnHfWsnq/lFy
cRP3tof1LeMyFWXO8/9Fo4MrfeoaqVP9IwhgAm8/b/JI3QRf/wCtq7K6Ko8Cji3tS2o3LO3wsKiC
5fGBak/Y7Z4b/D18XzXyE78F/a1dC5WHAI/OY4uVBFiGPKE49bxNfoirInXlcjlZIR2RiVtBr3hH
0t+rGaZVUS+/aon7O9a1MQwBr703TSoxHWWMVVzJm1BXR/9y0FEoMjd1yI8VOj9zxXrmEeyayQCL
pFlIp/sTCIBhartmCEaliMa6bLNL7w1pq0ydOEF8IcXvHs5ZKuGvHluzN3cRtmhDl34KTdPZjCI0
6J5hEwDApXBFEjaOcYzwfVrlKJY9WUoMUYdDLCjhrb0RPuRoO7JxtZgHWK9POZnoR81zqsQlCyyq
6bHq3ob/Z0I4k6QZEgnBmy+nDVQAjqb9nRdtmpd/ozpvxHeHHVw29GKHcclFuHhZE1AC7jMZrVsu
lty8NfH71xrSy5M7/JiYrG2ce0VRDgLfbfUJyLTA5vHPw8kam+Xe9A/94rIQ3/cPE+tepvDUuN1P
5uWMwahDca9gwWBzfvHSxFJLQFpkbBHtX4gl00D/F9tFbXkzuBL2Mw3Kxtn16YL936geeeFPs7P+
q+WSVOspyMbeB6wWLOGcZEU3CX9zgA2VvXU7g25bMD65EhhVrednwAEAaVl0Tjh//ny77nDlRRca
Rp/VzXozgZB3hbOeP/xmXjFBm/4q+u0whRGbXA2Kj62DZVXypzSNp9IuUrzV3A11G80hVIzWs/6g
mTq5EDJCafCVh4eSzYtGxMDyR0eFWIZbQkq41tvzfGSsvXrjQRrukxgaZl27gp0m4Vk6fPfiMsz0
ZlfP9YL+JKfe0n+sPXcvQVVmAO+Gp9V/GghuPwF9KHE8loyRcamUB1NssbXGCQRIlD43f3O+A0pp
PallYM00BCm/Omxo4aVtv/sIaIst5007uTOVkILLxHgs9c3dR+9A+lxdZVZAY+nQRF7yO2ze3Nip
e/Tsol/9lXPyvJWDVSHRokkd+Pt3fKBIQbxqUzWlhHz4rT2gGLgeSp0U5pCgWnB2zDrziBK312Oj
mD6gQ9dClBXosBWK0v+UfFtIdQWDRHDESmwO+HLby4/X58mVB1NMhsY/h/NkyL7oOdUxbhrUh52H
/r/gBPhityX3swkYQPymy78x+GFrRmlTHnFH0rPXMdVa5rnYg2MGLglqeyB7uS2nWkvynrV4azvG
fHIzHXtWaPQ/0XVdSZVlKzqTJVsrAjxXBmXNcJvDvwT1rmUgFl7yi1N8wCXEdP812dUqc8gsfZZJ
beNOs8G9i4qd0xxrUFBNMKRHaxqfmLhVTU0P449QRgfjqpmKrd5My3dUkii7OuiIm1vMDzPvVo9B
qaws3oZT2eOCuu7LQaTFs6TAR76qwTwU3cma83HOC7gVDraB+8cPd0rK93iJU7yrFeiXsRtti9Dz
T1W2PXnLLiG58s0TnvT/7rguMtNHgKtk1uwq8DGIWeLH++gsPq7PG+FpdVQ0CHHnW/opKl3tAR/r
/Fjmz9iLTAMwp9uhFx7B3lVuFwPZAiL3oT3rGtzTMW0otAPkUbqpFbpt8Q7XivD2YYE9a5E04oW+
ybVgDXpwUkF5moFdgy1MbWkoQmn5lEj2SlH8PYdhDWSLSrhceMuM9rgMZlm0J7Kg3rC7HnZ7wu/N
UOCBX4oiBpFgS263yd4tiOW8jthWymjuTjo7ZYDu6u44thDil0il34kz5AXaR++u484q/pZ3cVLg
67XtEiBCIo5MAC5HFfsPG5+6FuPwtWSnj7o7UQNGySDJ70Fagz6w0SUTzzG5HwauU45PIqqFBq1s
iTc81y436YdDIuJhlk7GBC0hz6trcLsMDuImHY05Jaykn2kyzuqTz4/uw2fItjhARyNVrVrMXq0d
AXGJ8ThtKcabHLARKtRQJvZrgaUBe3E1tAf+K6zMhTWdaSJALILIpGNn7IIuEFtd8fq4MsFXj36O
43r/JHjAh9yYzECM8nnsyCoe5wnW2MRebPqk0ZxiEYBzEXJkgVG8wf0reSRwaYRc2wnXPNakaoZ0
wn6G7kjM2QWieSqmBEFRMp9MweeYxok0+/J8QCNVDPg7dinds437ysJvfpX5Vsf+n9JSKpRrecYv
AiohS2rYeGj42BdKEiGl87xJNEBQRQxW0HZOdFxLocZ8/SsaFRolYh/XILirlMqXZkk2icQt9ltf
oQFq4RnO7p01vHPKrtewCwk4eHwpaWPn/zkqwB5WPkT9xMDHDryJB4+CPNmw2i81/XdIJFMM1XoO
erIY6ZYVvspiHWf9ftFP4jQVV17jDwCiZKxOfAkccc/8lJGPt5JfQw57h1ZLc8P46Hk+KD5sQ6pH
hJbnQUXzvk2fD6FbYioV3mDMSM9y6QC6saRnwIaFFAV0ib7tFLNbkD6KklXOmfQ6Q1xK3BP761pL
Sp2WSB64ygSzmnH/+WWs7iy6T8oASS7422leUdsiH9h1cMYEKRVSfxR4WHFFhQTdskMhc+2EJWAQ
bK8dQszAlsTcRFA0LJKWswF/6/VylaY1LtvUZZYRuPkf/5rzGSgcH5jneLd07BHYERyo57EBfLg6
E7dif4ffO23jEuQjUOhEXOa53KGcUiRtL0YOqvUHJ+JD/eh0WZyUk4X9EhXIMUVhGTgzNYffyZLj
k0mlhzGNgKYRYswd5FcvbRxBsUcs13X2oEKQbCJlY490sRkq+uhPboYjiq3nXgWvQMLPjGk32a2A
OOV56We/lrC0S1tdf8gyhLKb6pODKer3SlaFB+36Y/5qwyn0qSZkERBNs+aJ31T0MnYdD1XmgHRc
1Yn4Romto99Wi4Isa/PSe8UpESRaC1WOuFgMCGuCBZ201zmsPfhcA5XKDBtd4gjQ99oZxiTYJ0G1
CJ/owvV+8VTQTd7GlMCeNr4pwvzxMFLEBYxKnRdUS9XDv7RhewXRKRoCl7krNEYBVKBQIgn247kr
Y7+NrbM0WpID/0HB0ZsqlnKGUIIKeHh/TzkH7QV0r56WKPzkVssNJngQwwginHIVTpzCcrDfeQPi
pz3yS9wsldXRTn+pfVjYbvMJYr37nAuwdLxyJq3sZxnXIWslvfMGnH3lCJIK1wP3J+7WwcgY7WP5
aAoxflg+DGRWa4exr24EE5cNDQ9K7x86w0akywLMNieJ1fMLzv7ypt08tPb2ivK3WQyx9l/2eJTi
j0awzdflOARfjp87DF15B7PXBHw2iX7EuD/xEtUQrS6WyzsJjOou1hiZ+yy9P0b+NuOcq7yX0f0E
pBGpQE63i8WDwSoH9owu7VSlZxnHSFNhrtDnb1VCEQ2j4ptlVVib0f1yT05sOQKoxIOIddfQytrL
K+6mbe/8CQjGd4CXyxtrOZtkNAehPgTAMk395QrWDpIik2xfH7VgFo2xzS1dY9/+xRuccfWJJtW2
+x9o2ohL0HP5FnoyLqjY6rFRG6dsChA07JxNGIKCbbqMldqv8+QB/pAIPp/L3JIy20BScwiDykZk
dMh2g2YuvC+AmFBrwZlDNi8VfE3nh1wpDBR5kK0glaPuuDpXnw2yRb+9H6IDsPFThI6vHwiBVa/z
FevIlAQW3e1QLSddWs8Alk8hje998cSo8C09DM8f7X+auARk8eO0b7kQ8Wdniwr0RbEBqWQ/bRDP
CbUzRSBQzTYaNdCBrxOsL2/1tZH4Nzux3UDQT9ziY2374I0MVwX+FefZD0mr2+MBCDHOEs9CPQXj
VeKtc+CpGqL1UVt5NM1fW6LUkROpZDLpW2s3cbqzH5kRMpZ/pyAcbRyV13Taj2pSQsyHsj4gCRcs
0Nwdxy0GupeNGNg+2qIN2zkQL+hBGtflwvjuHMpNTrbrdsInz0gbGVREIe3JiD87vPwM5B16g3MN
uah98I2ozcF/CD10juJ7/G2OHpUgDHZskRXMoHIPgjPNU1b1xud8XQPPTYf1/YI1x4Xl4Udv2Tsk
CsIS7SP7Ln2/e/uIi5L/Yi+sNTb7tuKPH1BBif4leoqUfbmQoKQIJE1GXvu0r5pl6ohwimwetGJr
VK9wLzwlR7saj5Br01Pnvi9YrKu78Ic0gpFwuwbWv26ku+PsfQakeJTdwdO/xNMyWmtw/n4Gl8ed
DAXT4loNgDW/Iw4QT4IqRKPXkm/HG3qBuSi3SthAthQsQklrRl2doWFODV92Jjz0jQzb0vyR1As6
nuUh3p75UEY1La0Ifr6S9iz+p88MSU6G5Vc+DZ81aczGvZYI5YcRHmthPumUYcP7hVBXhbC6uGFz
V4dQVvx0/INhEP5Ya6kLn69/0ZYiIqyVKAOHo3Ban32xeRFQwWiU4LWcl8ipd4uqQhkxiNVtPWZh
Eiz9lovCMp/qanQ7apCipumh2R1itGlXve5md16LmsQ0Sj5Fm9kkFecBO75eizMwgbbgrzpnto//
wDNVO8M6SaC/sANaGaN6ILNJ/qKEHTNULqTKbqsecTyRkSBibNaublMo9+y6a8EEP0KI5qg5PJpu
uTpbM9/WX7p+Yx6yZbdiaYZPDy/ETag3jHYuqjU7FTpQvTMw2wqqsDLrx2gbxpQJQSSuowORwpx4
zAhY7x9Ql50qY9gh1Gx3/A06wbnZjJXVe6Izv74NBW4OB9vLezq5zu9VsqsmUrqCJnInIQKEzzJe
ilHDH4m0jGH32q96f4ylT1tK9p+gM9l2IuokQGJC5UyFLUvKP52SpX7rLR617uAO0Y0zRcR9Igkn
Y/HakJMiTWWIjM8fLWVr+6PxjW6dbzast8KKuQKIjDovkQ/6RSlPsfZWuPtFeAmyGyzntRLlxaiK
/qQErgXBUaw1hxxDMjlsUpozUgxTMlge7qOKm2ck7ohrifJwpFC149WJ+LjNWG0mraSIYPCTgOxy
ErWay2kmPb7YfPAtdjfoJfuLnqKZ8Et1awQPpRLiSBUwtnniv3B3IfCExMSStE/5t0MaI1L2zbHt
CVJ/IHlTbFXDY0lqRWvrmwW8uxOH9NKs1/qatx1BsqcB5/yeYSXFNGFMkFM1Kl8gJf4hZO5B4vug
IFE8ZUOD2CM1PSnDg9Rmv9SWngSkwSZZzoBd2jC03srVxwMqkKFyTVowBk6TG26x+2WP8oOvkyEH
foJyn2Tf3smsnPRpYq203C8625MTkSegUMrT2mpTaWv2AKGN/cJYFGPJInEQ76TKVOCPfBy3TbOe
kgcg2rcCNXhBACQn5xQnPobllTMgkLOir/Hrkdrp/Cv9EdhpvP/FhJ7bZaJSDVkDAVcxoKwCtSS7
TTv1nsf5wmT608Q+Who4ZlmBB7Wf4d+c3QQ5Vi2Dm1cIUvAq7e8yqW5S0ZHwizWyBHAuexnQwxTF
8Y6XEb/7F7CDxQMoLvI3AQkNwo6Qmb7/Odizcd5ic27Tcaqbqvs+qw0gmPLRZLZMBvYX63/zRZlD
QwiAD4CRaoDafUZpA9/OA9if8TBoByd2XeKK6Src1x69YGmjYmhJbh0sEpP0V3qivC5Ax0UxmEhg
BavLIe/ra/DKW0p+gpLmGstCh8LUSHSM0lkwW97awCexyc+WD+ArvwwHeym72VuiO/9Qs/K1A4XB
bPQ9Qjqtvb/bCbHxKHo67zucntKJsEC+zhlGWzoAiA7WmKCq9EIJ2FQTe3kddEeg4QQspU0No/VH
ESrJlE4rUHcJvzA5iwPPesbLYPqsmJvTRfbppw4PkZd4JlBFxuNfnTZdSFdxmh0cyCxuxCkJKE2q
Ux43H5kAejr2mYMm4iTsb8CK0JpPoOcT7TMDTDd+QcbHn9cq1V7r9ixkDV5T92L1FaB5GbiboaOJ
1Av2PoBEzdzoJ62XMcCms3ANhdXvoSvZkOr9nJJsLEhwUuvOdEFfIeK/mtCVf7vMUG4mQUb0G9DI
bv7TTyouGZ/blJVPqcB3bzDOD0EasDYlqhSaTg8ZRN7paOzeIv5gz5u9deY8iNPPCvcBEH2PkMdW
2S0mB/hCZu/RgXU7QLf+eqGQlHLgJ9OtgQ+B6vaVRTQFEM8ebtW7vRpsIP76zme5sGF2PFaNPOh/
DD1J++h44HxmNfbvvbPJ6wTEwIJFKYPBLuD2czTcxlWNEX5SjM7KcqG1f8Pu8BdaIQgRTXuKeuxJ
N4TAx7L1fnjWo5DFVD2tUOQDpJtZdY5AdRFaJ5hm0ft7X92jZlBzXacX7bjT6HLdRaZvBhAH4M20
TXMV3faMxmD9bncP/DJYqokjbYc7Xtj8F7IvP2AvxW7UJQY090PpmqqVaS1ahBUXDFtsjin3V+O5
Kb1isWUY6moIP+4TTupfBmAAusB6V96Li/JbpaL+2XZaqnGkovygplfLy1jQAwW0J8AdtW1Nyh/F
rYN5FfQ/2HLliAGpLXSd8hlXYBpng1vODJ8D4Sg8Pv0/b/9a1Wxd8cXDeR9luxU034fwrwV1EIao
5MC7Pn8SbZhITBcVj0XzPQnuFHOnxFvrHGNDPs5QUPUX2rq53kceQTMjQusWwDdYbbFCxOwr+7lu
MF7qXEM/vMJt7b0sDV3Lx4JLitUa9A9RyvpLRt/2zrbjigiL/WGjsXg/4o2TXBrN2vc3Dj/8Ivsq
rh5vhsSZKKf+iubUgzDUBs8mg9DVCgiyS4o6sV0brU0Wtvxw+P0bCOxkmf5MHQU++OJWhmXOstFd
jV8msSGzJCETFhEvhYNi5jARDoo83umJLycL/offC376N1lLsyw7l7M3oq1MTZOD/r0TfKV0cL18
dK0Umal/rxWNLnIrSdVBaJVHW4S94xj7LcdtneToTFd0zX42B5N868pDiHSPoh/7D5qmTP0MTIqV
w2l1SUftrqDpHabKmISQcvh/4+CL3Ruc6O0wdA6319xBxkmuIOnlosDlnSaf5CCgWU7UcRkWJi0O
2L4ruIt7Vap+GK2sdJC4SOa7fo+/Sq11YdqM98Ma3seAntiNy3Q4jgvrm+p2XfagGyczBhyOS07t
4ahHNi1jeboUjwzUtA8yKyTbgxSbLsEVUPcx+EvMYY+K7iD7FSSuHJWNZ+F1OI2m6VdCXxb2+Uek
vT45SnoW0sLLKz4MJq2A1S+upQcR3BIOdRpdclwHfI4c/aEoC0iMh4Wx16CFFyj5BWQExmjXWYrE
u6ynyIBxpAcS04g6DW9+I6kKSDE20OuBHMsLKI3r0f/8IDyVLrS4SZ6tuJJlYJVm5uCsVjJ5UBhM
5zIb53Fsq8FwIpwP4iR95Y0tUjS6AQr+EwESubJJbOGfX//+8Y1nM2X7jHXCfQw3ZlX9EGT9Jmkw
CS7IOkVLilXws0OVww3FTSowDmSVN6A/XI4NO1e24iGQMJ0zSTPyhhPl1V9ru7Qu0dK3oZv2bE7C
EuF8zNW//z7KDdnoILApE8a784rxPRB2MT6w0nRDhtkgtSuQxs4YGb5cc7y9Wbz3D0LzkeB7dbNi
D6ffbucKcSV8UmWp5PSahGeBTpguRd6vMyPHJfl17mkVE80u97CvJj+q8sx30BYLGfceg9kKUi/K
5Nw1t+gthJtyTXfWNVoSRLfJ8KB2eUhdJX4A5IZFX2aNxifBZCCcrknblriG4dscD+j33rWYymtL
KIp1cgjCnmvUznemdgqq7UJsShrR5jif6fmqQVVACvlt1uCCar8ffzrBxWVtd6O3xpUCY2JLLCp4
IJmyQc3ei32/2pVpj/qx/HzDpuMQE6fyx86wZJk/eSWOaK9v/6xLL3YSVHGSxcbui1AMhzLf3Y6t
w9V9oQwY7NMLSaNrdI3c2wQXsFG39oG/0RCbWoGlZcy9ss3845al1+0e3HpCdMY9pfF4CfZ8RUX8
bMiiLWrwNhK3PbbgrSybfeo+0N2WPXFah/pG21TvxVjXIhPL65a0qxvUIv3WCfiYx5GqTBkbCdRW
9k44pkzV3/wYZB4/3BQsWp6XuCQBxAtQGXTTTq3bbvAa9vgLp/wx/Lto0puGyZMgdQU0r05KMlb0
YiV+o1R3oLc8GDwcJNsbuH8RJuUj83hzqDv+TmQXz2SLH6ulOqh3jnqsWCf8QHRJ/w762yHcILD1
8/RWv/UlI+sxQNFY9aHzwiKpOz99gRaEA00NKvmWakOyx1pZ9Wlyk8T5U1MWxvXsn8VKFW9ueuHH
WHLHrZt1H0smEnhbgZFpChgd4j8uuIGhUnh9Wk3IMAY8EmIzoBNuM/eVGqLrG8BtypDrZL6ibGy+
D+qTSxglEI1GvlCOCObsDmi6+i/WuIwRgSgw6V8iuobsAt9A616esEinIdX0PwbF0Gurr+beDXyp
IPxubBjW3ESt0wYyH/oUUwNc9OHByJpLZ3q1wTFIDQR7OgXLxMM62XUP7BklMpTdpAgFEWqM9VS3
NEeywDL3d7PYlmpOySR8+6d6kooRN5M6asuTRixhXh+1aQHhUtxY7lzNWXCEcPUrQ0WfnjEja3sx
OWjKkdZyWiY8Elp/xf5GzODtwx8q9FlRGeZ3GqD9Tgf6wvZ3b6krJwX6CeJ0A+X2B1VZKXiq8FpO
kp0RxjUew8m+FoSUFpKaYbMLwBeBmF8K2Q+y135YJ6g/0uQsf57je97yfPNqiMT552K6HJtbFyif
Sp0FhxTDeonDr0TQyR3ScRbfU0X/HZqqgIBA3tmcBJZbDqRHdoiilX3CnAdADxkBQwBUM+gv+iqD
CKJBPVaO0MP/E95o9Hykl5adX0F/l2TWWE2mIYYWcOZqT4t/TwtSvI6zXte0vB7XCnX/wPKCjUsX
kJWDtPl/veZ+S3kaea9cbuatC7mLfFqLsi/8zYuRzxX7He/aFKEUMahJl/FxyTjPJFOlQCBgF2t2
F4FGdbaGrEKL3ququmpKpQHr16yVJO85aBUXAYxc3UUt02eYXBod7Vv89POzA6OG2nHVQkel7FIG
kkXSYLazHH4E57G5dsY+EzlJF2E0tJ+YZQryTdRjx4HL2mSe/UOTULaWNlYqien7uNChy2Xp8/dY
hnRjbfurCTx9Aq5dkBPwq4Mv/aVBDdv17beuI0Vikf2nt4s0mxnnWoGHY0eTdrKdqsWSu3hWneKy
dbZqaN1bqGe8OIBdMxb6V5rUv0wq8uro9h3dvPK5dR22cWcYdKHkauJyY7gI1k3mKGTsUWS7+vqJ
T6SLhQdvAl1KOrzdPMrs+bSA/CH1zDeW0AT7LIL7Og0hqOaIIiIdhvUUs/BAnq/kAoDzWO+eNC+k
wnOJmfz7TRnfOWCu6Rxq4SpLpubSAcNRZ64Lr82sUJ+XORKLD4jJtLhIk8H+1+35/HjE9Jsqbhy5
j/lZ0yM07FnDnhcK+gpfr6MdEKvjvTJ3drydArvB72FJcN4k/84rh09WzJS/F2ve3KDi+/nxfCHQ
4NfdiSWJvo8fCTXQHzJGTM8SNOEYerflbI5sOA1/H6vDEml3SYadNQ5hoPvxPAiGlVUJexhllkhS
D+kS3mhhFoCC+KUMMLAMbhNQFzIV9hd9KIeGdYJ5uVCedTGk1rv9H0DlCW2XROhpBmm2lmzKkZi9
T//zwk0Ga5QTUFfxKENnri+nSSC6l0JSyXzezWEDYTWatWHqbKsG2voiatWG6utQjXGtrE3Zhck+
zyAkahPZuyCewtpnUz2+dBIfhA8YhQPdLGxO9OGHLSZUGAu99XBJtgt97q2wWCSTRzdGHhZTwU6e
Rbb9/5b6M+a5zljrm6rAVj9YRKVNur33jE+G1lDERngB5JPlxMEytkCkEU7hXBkn38yRggqd34m1
YPsAwU5vSpB9aBzjqBJhKhQYh9XaUv/YRyWFJPNjxaoPIzB/D9r4sgl9OV5XuaUuhIOBK0iQKGwR
AFxGZ9IE9j4nH5Bl9edi8AP2ItXg0fxmvEEehGQjwhOHn/0+22iMHVC72l4YFPKGbnJw3M0z3UXW
P8hQIwALJrMIpJ6mzM+VIu7UXfEWyVK3kgpy/INfrV4EkpXelRpFUrBR6L+Vqo3GD7F879CXn9kK
bydeXVnf3ey3bk4P4UtdDxtl5lt1xnwkXdAOSjXNLAa5Rr5z3yCmLm/WzKFYvukz4pJRd3y7Uxrw
bb/xzslnUcsSWnGzFbONjObbuhidXZn40pjk6WZSpaDP8hnsIU20e9qRyTG55/jxvyi/IttU9AVk
YIZVZd4oNvmLcEvm7uCLzeuEEdoQiyuUvEybc8Sg4wQ8QKqy3AU6j2SFYfW/LIOaXSHD3zKQV0ri
qmmSumHRsbiyySvJtc/Xi465OV4CP+y7CUSUp6w1DgNpScuGmVnTxb3VfNx6DsNzjXXWmweYZ6Hv
l+18DULxBB8tpvYtt9+n9my1QnR2D/PqHzz5yNdLzpRNwhIN8AijBN3QMOK0l7QzpsLyes8s9I5v
9Miey6DgE6E1y+65dq5NjD9NhTWv3ffg1H7kR//dCDWiCnMenWH2OFVTCwtdQDxANgXgnPvs2Dzu
RGIAAObWAaVS8i4L8onYeCT7109cAaiw5EnbZ0ugP/wtSim7U44l9Pn4qkOZrc3hJGofZI7E1BhY
BQLTHHGNuI6T5P52XIXvFWjeCCbpKeETXi0S4ut6dEc08bCBe3ZyCKX4lUzof3yNTFXlXb9ryr15
FR/od29gqVvCJHEsxVw/HOuC/RJ7MT+zzdVSVZQiJpgnns6ml6ELrWimSjqPKiHK5gol40kaK6y/
IuZ8lIW9pYgDFWZUBBCQFRBwVVo04lDh/OjF87VAnt10pgfd4haa5TjNH6rPVb0XstPUcFQ785Mq
4fLs2nUNxpSb8u/MmuLI0Q+bM4Jj7OrYyJQwJLNgsEdyH+51zOmv7Xb91Y5+1UvgjvQcuFaeNaT4
6vAwqq23yJ+W2YwBM3XHu0EvUsJ/qR7+kzvF5mbke2g7suRHtHQpyvcZU7vAbtP6VDvFhubBD6jd
CdPiMhT2o2ydHqgMelapEUajRLxs/8v12LgKklYJPvdeFfAgorAsyQ8Btns0bZFpNdYEznKEJK7x
usL6RH+d4/PGgl+Ayneg2BEL7hJf8LCCoVKxyJlg+9c/T9JnSeoHmRqmp6PlFds8cQtTX/rLSyPa
iXUu2hfTXzMS/AuDfwFolhXtT4ApVNKj3QfwrExP8A4wRcq6oev3+f5rB7JTBleiAHgjHSZfMw0O
6wamw87ZOu68rE5g/U84b7wpPDhjBe5WJMRiK7aaQMyhKESgg+2o8eVZPk9Flk0Trok621+VTT54
8ygiFKVoav25z6uubrNY14H1EYBZmnGXytCcSlSgN6ZfI/RaxgM0cisslXjQ3pTafVNV7c0Cscaa
L9hnO/D+DGfBxWlQ6XMMCVkUxraD88L83KfqF2GF9ibo2mxCK+Y+7YRrqPOKp7gqVWTQ9PaB+Bau
3AjFgtQUA43XtOqonNERAfwiuKNkhLaI//vzlf7mcpVRZ5LpAPh0Tzj2JdRBjuW5474pbHQyLy2a
0euhrPJb8MyLihdfmZRkYqr/ZMxWaUF/MTYtEFDArIRXc2JQp4PDKFd6kkhQsBarQaH3Y9rCFkBS
JiUMGxY0c4h+iXiA0DUIUQkJF0XknyFxmhMAM/2i8ORQle1C7fbKs1QDUaItaEdfilMPrntHHqGl
V5mklkOLjxoWUh0ok/i/zf8iAGRATXObgvkYWpo7BbnjXdDnxc9WF8o4LaVbGRSiASFd7emjmwo2
TyU8BBrLCMu9ZIK55BxLI7REg9KNhXs89hUyW0+ebxlMAZxREsStOlq5YI2/e5+tV0+Wf75mNVGd
ZEwR0q5zDMxFxUQxrhWyfTFFUFKW4XvA9PFy5fy3JPymD2phEDnb3HJkPYQJPyUNV3dFJfn+nPUl
PTADynaxLlgd/h0xsbEOj9q/b0vD6bWdgOXe5D24dBfq3NxfJ44HzPF1tRbKCvVfLhEOOq79CkaK
tpiIK2ELzzFKgdOJ5sbdcpQQoZvSlIq/TdprQrISJ8SJMiCCGgBpIxeeuTVQRXyZjYDFYrjGjyne
fbSc4KI9fpERSm4V4sFfl8plsWmgyHhzOvENqAMwkiIN4Sre3tafW6t/lqBnaoJCY8PxfqhcOz5T
LJxotCA/x1zQ/HRtmNsV9CQDrnHNwDMM/wVJs+k8sMtEYWjBX4NtRONC/HShnbcM3UckFmg0Dt/7
w1XmUAIA2+bisM78IlcLr7bepObo/zjFpO01YPLmjpa/J5AQ/TzvplZxWqOMnaGWoSkyCJFllnzq
7yV6UDhQa8Mcwpyo5z7NdUjxLXuatDO+4jsdIYsEUR9cLRaOEgrlx573TtxaP1m8xUzoTT5VSyfi
OpEZmlUHv7qdQwi+Yo7/SI5v2I9akENDWA6TDhSEH9XqykkM/W7oKwtJLlBcxj4DTlrcdxJ1b/WB
SG6vqg4p0zFW6kwpjuwChGZj8oKqkhLm2NhSJxoQAdanGhmTKi62KeSkQMO3/G6UrUnr3XqugiSa
E9ZD5MkCi28CtDe3LJ8X/N2JYpERmOrNZ8TGGbNJ6iFCGsolZrrqFymLg5frfSPVMVqbl8XKFdOm
qy3Q6eSoB2v3lLoiGai3ZB7oFcCjYVvqqqNomYHwWjE15gmQYBNLUf01S837zANnlXqI+HtZFk7G
NQKZvZv2vlc97FREW/+0LS23v7Mr16xkKh0uqi4SanAoF2mzZcdtMEZfuz4FkgYarLI3WsYX8Tmf
DW2iuDnw2RunfyshfO4j49To/LouU8e0ryxztSHwsJbCT+V1cmMczQKE9AepCz3+q145p7M/D7GY
PT2M2QF244yWCF72e50feTFokh7pwjW276HljgspXYtx9DrsHEIKtFrygj4KPjlVsVfS+Ay70TPw
Y30Z1qe+imyr4b0YvuuDGyrtMIkrsBuOyvQSdfONCGx3/2Es61xIcrwGXQitbFP3/YLkRZwYPpX4
C0DxWoX+iVBcTSS+FOYdoHDFydZiGyrRfzf8NeU/08NcA7LJjVbzuDUVWMz8kk3ONoJ7V4lXffFw
bT1b1XsRTAgzvHWgJt1JwGh8eiP+QF2469Gt8tvSBoPfI66KxPABA6WWA9u9lMKTLavLlfRocSIL
BYWpoy/GovY6yXkVVhwpmYoOx979CCFOBF1KpyNyvsogj2nEffZPdMPVFoKKJ0eeuqW2k5mFAz03
dZ4URLI6A6K4MbuyioZRAWOB5Zo/NTXU6DJW+AWD+cG7kS97omRq04IBwCr5TjOd9RUs4s15zlyL
XH+6gAPlQCvLSgCHVQAkMX9QHHoMpnVuj5GDpJgNlHgWWKgacFijmuz12esIURecqqzp7NOZW8yH
AWqQFaxlM7VhMK4p4YBo3m8fu91a9bXzb9Xa5jcg65HLYA9cteyRsb2bHq8uKZUAAIw4tSOYK3rH
WVl77/Yn2UysWhnHNa+HVoEIQfQUmPYuZZNeAx31r3PcmC4AZalWNtzB55JgbfXrr7YFI3siyfwC
72chz1B736uEEqXPfx+UhyH868ZsndEYyLZa8Jk81QfYxX/p+UGXpUtKTYsQW2k7CUNeQcki9FtF
p2TEcfDkjHAJH+Z4j5dh9dg2CC0EtC6DTO7O7sLsS4UzM3zcU0KUN0hYyBx7K0Rl1Qe/LJ86+l81
Cbc5ng/UG8cbgRaS8NVxBz/HNesgacV+hJRgtiu7mEMMyq32GvuXS+5klVHt6iRzBM6jjnAn9XMe
OC74mIUtHMMro9O/v7R0bRK8urh+oP9tPIuCePGOIAKT172rTafTSE21uTCdMABjf+TuJb6oI2NP
3fVAUZGzyD0BVLTIRSBgLqquBf5QFjN4ttUibB3WrpZtWUro6eVGxyH+ENYH/nh9PtLNlceBaM8B
3walydp8+PKLqUE5kugZnCP5UWvufWuEeLTViRAwi+3Sht/M0w5/zvh1wITiWiAglzd7p1zf/QFz
Yguj9PMSGjkIiSXqodWHKNqCVwv78bzs/NPThXnzs6rpg8eMBHnmw69LiGMTWQpBWgbY5P/LP+dR
UPGYdVF5Rldy2napFWW9wEZQMe2qXEsKnfHWIRK5SY650Dwarz2JoR3NKVUYfXVeSD8OrXXszQI0
tgJWCaxhkV2rYa33rVV+CwwqqKpSBhTNtkkNuG6hlaRuikR9hDsZTSmY0GxAIWtFZNUZsbzJNZU+
vLnQgeATlMAXReKI5aUjo0JIzxiJF+v+BZ0JH2LoqeUFXVXb+1Atp3e5Yx2hY2fAp6n4nTvfOSRR
yHFC1kSMlXd5mozPIYdkHEvRTtnpYjJW8a0aHwaxSnLCd4RDGs1AgLLNLbuQZppjdVBBpmpux6QK
7Iu2I+NB3BI4Vq9/gXYuUQc/3njQbJCRd2d0AyAfOCheZgaM/CHEU/YlHvb51nVdBLQs+Q3pdR9f
PZCGO82QiFtoYrk1rsyRlude1z/x/+0KKj/ZUoiE9zNUlzQA05u3lv9NvXuVFZwcCftBJTRyxpxr
auwml1npDtBgCE/gpXlbm1cz4b7+SUAVNWsR5hJu0W2khEPonm5YNgqDX483KSWtZUYuPXXZHhc9
b/bpzzUhNzBAihFrdSPvSgfoMe2XOU+AOCOQd2OwOuoR3vGwuw6tm/GZLdpolQbaC3YNIfgqMfK3
bJ+ysFcDMBfC8H0DuquCTG9eFZDDITYABFG/kmiPdEtbgpa1kvfBjH6EpVMIavemm11W3iM8gKQK
t+V09QtU0s2tvlqJYyzkqpWbVhNL8R5XO4sBhIKFntppd5uib9b6HYyhr6oTApdPQ0kgd0NzxGdp
YSUkmcziruF5TWI+SrJvOxxZHIyFKtsbhEKl7QprV0CbqdvzgZOW66y8BJkHJAw9ZVrj2/L9nq5m
vG7HSSBmQ2BYu/zDcJLOL/V6nq+T9Ec7DG7aBPscCwNhAK1nd4diUsvw9R+stNTwibHJzHqgBD6y
0mJ6U5dZducQ+EkQs0yxzZ//Ut7hV9gS06eS2FsxbI6AReNK/Pp+x1drH4ZRHF7Kqrfe5U8u0o/M
jQnSx2guzpGeG3GHEnNh6yB+nbSMt9FF+5P91bn4nT6TZe3gQNOKetTF1Fi63UruNMy7kGqUS5Oe
SBAiWQekn/7zjLcGnN15PEgoZ6tq0XRBtcgHZkFp0mgTtWNZyx0QyVAVgneAQBq5RGShVMvFLJuC
i4OKyCQZgPqm5epQhgjgO87hdf1YFw+1Gp5Xnw0oFhQCkgwEcHGcDmWKri4JUnFqWPJBXkzyZOGu
G/YdPW3xrpChP84HINlCcmBEU6V5E6A2s8XoAVcZAfrTfGIxPTq11J7N5hVdCR54alVybMW/FWCr
FII/KqSDsAvVlBuB8toig0fnN2ENKs/vJWC9jrzvrU1OKcikvgiUcLSWldLWuhYzCkFPxIdybY9/
xZkjVYXODIhGnulfFyElvjxFgssdfBBDyAuvdTUods5WjiJ/E2OsQCj80It5WI5Qw+5KRUPuxszJ
UvKUyqProqsPdBlKtBm80LoNgzjzPBh+zowMd9Pn3n3ltOQpS5/Eo5OqqCXO0YfCSucXrlZrKAo+
RqwUKsaajM7Upw5w7S/DUQWNYqHUrwDBUftyZkNkjX2gpiQJmcWIOQ1UI1tf//NXEcZH134HO+Rf
WuolVIvBWgRv263S7FMzh1gs96ZvbrE+XhNa+IaSsww0qIxgbkfwBaJE0jIf0rGuWu1pKuakr9rc
xqmlb/OXC/jEdKUTU7GAmyzUndiTyt5BDH7SkHcLR4j6wp2oFmECq3N6g/9AyQTj0lcMp+l4gmoZ
xd15x1FV6D9aEhJgTYWle/V/V6M8MIPzPZwvevngpRUjdiCpviPB1n/1DVc+0rC69nO3BafucgtC
rYw7TG8FpGmDuZswZSFJNjTWZy8VImkXBOjUho4wO2v61JLdg4rCLvJ/5JT36diZE4E4wh1wxexU
Ns1OEFQlXW3P8MgCd167OUpDrWXg9HTvHBIqHdWLWG48EoZM3oZBcmzqK1LL1TGn38GRLBsdOU9Z
K7gVJ0wOvXq7hZvB2409JVl0MUQKKkTcs7At5HqJmU/Y8ot74UYv6hpCzGZBao18q9CT81gN0mJE
ZFpvPag6L63CCWIqnt6JFhq7bnY+3QlfGyOXCD++tlYR0Z0SAa1e4s4r/I29FzRvFWy6lnck/SM7
9dXQOf2NjRMCcni3YS8IYVfBhpB0jsYiUxl8gRiyYtJKC8HvRgXv06zjpXQ8EORG8dJoiJFjPWkf
0fOOXCNIDmSkc0XZBEHXtd51yAK5VgPuRA/Lm0RST3KjoLXunPXT+HKUnkxhRyM4tDUFZUixS6o3
m17k6FT7621xru2wF7h8M0ZC6/NzuNZJNIKUgTGUhQBuoD6ZiUABzSuT27xS3QcUuzJzHD+TW5if
7Co7oVj8ztFUrgZwa+flIuk5OPWqupEw0qfsGILegk71oLbzzbdbHkiCYm7B4lKDCP4Ae34AHj3Q
IIf4gFviZxMos0ghM4EDn5aGutnFT1sCG6Qyftrq/rAMesGlz5hFEHp16V9QEedOeIlBvM4TWos3
irIxegBFxlnWtSs8qxTHFuaUq9QegZf1qKKfCT2o+Q/d7mnbk1wICF7LWczcu3+/Bcb7RUYXU/pA
KDmz0S+2oHXkrxHzwUWYqLLARfiAPusmFm99jVH9UIftrv0Yidf4PEppd2KNtQ8FW+O+1oNlTwQu
NhRkZ2djifRaBbIOJKsUmXrCAJFK4xdGw1VqQfBrw4Oo9TCzZ5R2FbrR85h0DTJ7hkOKB1KnMznM
O3ydow4AXh76CrmJfTXHxWGT821LXEJdVZmGL3wbraURDAYb0fiQNDzdRxhghcJCqg6Yy0Lc5ztD
jiowqaWHGAhfnAfniZSbnSZ9d5d0Sdb6TlF6acq9qA4joXprfPfH2dln9MHWir9D+2uhb25FEzPv
bbv3MUi1f45i16/afhJl6wJAPNuYNHbDMTwllklZfi3Z5FccbaoeBU0kxk6KJHycsCs54DOFSCgM
W1CD1SHMI5dQ5xYFh7x3VEPr+Gdc1P35pUWCNesHMp4Qy51bfTb8HczDWU10Qa3GJx/JAjh4Ovk5
yVpiRrGpxRFxJ0fOexh8eitFG6QyWhCezussv67dOiy76KniTGuaRZNe59SHRAyR79Mrb9FVogFR
3+xms3ghCKu1mBsuRFZA0t8qhGz11yTpL4K9UK7bdansjjMU8mcX3tFohxi2vrF9XHE/HT1t+8hK
/FAZQoTuw5MH3suZM+iFT9V6N83k/W/43pywCSrRk0nww8iKLwW+SofHEXVjvkM2O/dZXORdg2q6
bXvC9rYzRsLQ8Me9TtnjCDilobqXxxfacjpE+WANFBdtoe0RY5IugqJUGdpHVmZWmgsXGWAp3iXS
WIHRb9PV+HfOpxoYywf+heVcK+h7nDK774MtfkcL1tzJSJvleuuMDNROkmnIFOTN42UDq/US4OgV
LfHiqTZyZWri22l8TfEyVXdzM7OGIqf5/19Z9Bg3gKjn/gtwKlc/zkwAeRUjh4VC96j0elWk+iCL
3dvms5i50ufrGnNf86PcPBHHmB9r4uYGB459ZiV4dUlK0hlSOvwHegSKPCffEqb12iL3rM1kGYZJ
+JhxLGsTYy0kkIcMBFQckUlyScz74zRe4fTQQ6n3Vu3vsJ7qt4E8GvomuIyg34Sh85BuWH0CEOSq
3DiiDAXJeI1dUh8iW+WAarpPW23yCGhAzC1QBmoGlY4gaheS3Is19yiemd7VGv6HSA3rDc0rGJNR
m53xZMrE8NKKmkR6W7eTJqRlfbtwZpy77xN8R9qHBLSJtQN7eyDSBGUIkybBAaPHlM//23knsSz7
dJ4vLC2W9DhLXGWF3sGPcJMR4wtHXywK/BK3MdIXPg7XO+9lPDpUj0V6sh94u18FKLG475HgynGE
dEzys8mOimETDLQwxTAFP6aW9rreg9ja9eWjyXRi4iPA7/ocHf/kpiswGJrDUM2vfZCNidSU3Kxd
36zfVR/lxCLCxfBxvUHMjQ1UFzJBFpgyF7k6Bt8pSc6D6HDteOyN+RSdKtZJHtrqUPhRJUIAf8i/
mAE09Wow9cLgcl6Ku3REj4YakqsINcuBzS9XMMEd+0a6Y0vpNz+qpvyb6prOe4fesGZpL2q9AyQE
u9Hx9ZF8NvDiZvai0W8SyOi6KHIi46egPw9ffoY3XMqLPgxmMVukSsxPDDv7JkP+xCwtB0HCWRyu
FipqOcxHNhGLkXmvUHUXqTc0/jCNH0//e+SGh5C7TLCbTxQmnZ6VNfHQxC3erz9H+WizD3RdhrIH
VXqDe4wqFoUddLLRBMDVVVtPSMkvHLxhS3rZiGp0bgJtu5ftXoSl01/i/JVerQHw7+XtiEJ3HcQc
QYaW8WoWg7w87TZFAVuDm09Cu8+jHviVFOlXTKkw7egPkl2bh3X3m0vbcrqX34jdmZHkiDo9oMWy
tl4nj6xJ1WvTPlXF1RNPNRYeVe9vOXMVlQ6leIAxT1nVuFz9agJFn4pjkEvhjaqNEblMYbHAMPu7
N+tgSH37iT/A8PBI2Y2+2vOP0jFApg6v/DBW6hBIw2bJWJxyddFbgXfDBAuw4+xKZF11jgoBGXZO
YDSlKuIb3fQxkui4Q34Zx5iQdzXRmYqCgoEq3Hgm5QWX6COKdHyxs8RfGLcnMbaMr+9HEfG74eZL
oLtf1sYnCcpRm0QVflhyoJmOLGgxW+IZaIpo1UocbMwNbTFgYUZozqTWyvyoziynp5v7MCJ4AnCD
TB0gxQYwQY6dYmKSud21JzjHYNhZBC9j5DoKDaiTrbWxBzk8X00Z5GIEjikoN3rg498va8SpFDt6
b/TZiTrQIpcolGTxwpRVr52nmKM/Jg3ucuYXIbBC7axL8aQOSRbna8Ec29JyQB+SRPeU0rlJc8KZ
mt74x/R4lTrRGVHcEMay/EokDJiZz7dmnJnRJO/+baH+mCEWRhh8uz1kECRniQ3hONCwDLqbgNSE
YUeLFB8biK+JOZPeTdV27hRWUlsswbmd+3Urub+ZRlist72Djybr2FcBDqM+kXF7SV1WJlxfmwgO
uRfsd86KMAQNPh63X9mnS79nV4xLMf6NR1dWnzZZL/Xt1mZ7eGePfcpY0EFUAcQAItNbz+0J7bWH
m3dy67FYIaAxt8rvBcaRmdqDg6Ev/M1XthvHH7AnvmKQg83TD2RHEvw/TUWsrrlLrHCKxBEh41N9
Tjde7UYLhnRTm8UADlowHtBjmW31VEO04dAdREjhRTCan5OEw3TX2saZb8bNVUDr+FMsftYzdPaI
PO5cU82R/vFKBtgQaO+1kYHobrXZTA6MuZW0LKGNpsdnsNm13w4x+LueIalUGLULRC5l/qYxYEOk
AC+vOal/LgP2wxHuCTVNAeVvSgtlpX1k7UoLIGMoBL7M+PZpVtQKriynhLIGMxJD9QfEeoLnCCPi
V+e8AyNZ7gVsjy18kBZduB9/Bo7Pf2UYe+qBGarOf/7RtTmbeMOUc+QBvXvMUii0nTuSVBiQBfCY
keT1OumGSpIVaMZRokFGnHE9U2Z1TtK41ID2dc1q0uleqvLbRNJJW/h/p9dAebdttsYBMFOut1nj
IoaDq6gIh5WZvdH3D0/3TciKnxLsHt9GQIFdnynmNOxwprjrIRPJXLi9YjzEua1MMeAfSa/ft92K
aim4bP8QM5f0WKsDeOkBMfvkPxV3ziHLGvI8LYrJ+EtqpDRBpa6kI/7yCvfChhGgypRV4aMnKPFm
UEBWM6E00q9VAODaGKp1FhC6pUCpoNNZrqlCVBnH3g1CgQ8utsoXk2ZxvsGRRFM/sKWm7o6SfrGc
D3KXrBbfoAbp9tUAzNI84vvGZNlIAH/k+4W5nQ8r1do/tBwzF6DznBLpUQPKQc5qwfYN8RnvZYN8
ja6iK7WXq+E/YeyyWMNDEVz6LQjZUTafe2zDIo80hrnoB10IRUxemifOIGfTmm6709uMa/9r0ybT
liSCaNgxH9etoHI2scVEpbVyiVjsHo+wTtNSeCSAC5eSKrBqSt4CaPCTIZTaEve8Z7J5lOaKq0gJ
GLeawDDjVwhq8cpRhqYNxaRmp52vMQTDwcjgf7ew6mEiE+BIooCEdIytQaSzwIdiIF39Z3w8nVqI
/pv0jq9Dr2nZldcse0m/V1WLgVU16JmP1Fifi2veEOYj2RPigVBy1NG6YlS0Vd7spw8/aYOYaTCz
JI9HU3tJrGDgvQu6jlt5I63EqnXk05RJ2LBhBUxbbTfyxt1qqGPl4KsWSLcWBdwkyyoeIkTHXyM2
We1AW7dpPB3WfinFD4nNbv5Gjrduo6HBvM8zzDw1d1pFbTAfhYZ+jxRG1OLeE6f7PJsg2GWSbq5F
7eB1wyLBt6mnRn3pNjfrtB2rxza8OW1PLmhbu/v5/imcyJcraOWIhBLL99v+XKibWyxvg12OtmEw
jpdT63LwYFNpGNAXnbgxgysf5GBlqvwUTd74V8mliBOkRGdzuljsHQUoQKEfNNVHVh3XP/izKNff
NMyRi+hp9BHh99Yv95n3g3j40dBhlyvqnN1ua3ZuKlQGAXdmnkpf7BoXNKCBs+Y8Js64O9zfDAef
lXy0jngQ0IRLDZRriVp5v5Uws2nyMF9d2pA910fPfEfxlAJUwW6qWifFgvUZhgC+xbrRhIkhSJuB
cpOuEsKxwKarsZoupSL48EyfJbMvNyGxEFdTVTOVznpgXqU5A5ZDjJm/nclooyNglfVJNzoVhcEG
3UNZ9CYVzNmyWsVXaQVGqMq+TPi3Zjq3g3dhdVB4EwxoLjqfiU5skfbBFtGPIrgMaYGsaxTitf9i
N4VkXHL0/BBjqZ7HLsIfizOBZvcXRIY32Xo9HuRIdcC3ft3ND0qDSBi4Hh5N+P/UI0QptUw+Ltfh
e0kFiCHwGc3jSUDL9hcOboCGnxyZIFopq8sEw7cudR+t5ZK1o6VW8BPUyQfQnYkb/42lBiE+fH9/
KR0tttOxcB6XYzahxmC2TOvd+IKFT7qPg+HPMYoLjLe/x7JQE+0c/ow/laeoU52NRDDOfg8OPbd5
tUlJn4niljy/mrKLrfPJME4vN0C4kRDSNPCHd4KtKjPhn9DCg4/WEfEdPm8WJROWPZ4LjcfBs4+q
lx+0Uj8vRdiTbcQFtqcUghFO4OxjtBlV9SNg+bzYlNhdzTUf29oaAkgab4MWHdcI5Ps73NyVsumb
u6XSGzZ+xa8gkMIm3TeQf3RqL0CzPQsUrw8WHwj18xR4YoILO+5DG/setGQbOZr+DJse2HBqSFdP
Jy7OsAkdlSQUbYTedA3PC31Wv3c81gVIHUF1PizQW2IMsihsxg7mz7pyCwkHX5eLOVqyGS0ZiLNw
XQlOUmntRlUENn9tvqSvU+G1eGjNN2QMPM64JczlKZUnSMli1L8pkWlsRC5qx7QhFilydjJRfnRT
vYLj91jkppGM14cIrRnH+16ANnqPncAJ/EWqyU+Kw7O0kvR0oooWT0EQQPHIAGvRa31HDN0Xp16A
BJja4GaqRcaO8ML40dG0tTf8xUiNUzNZNqHAb1bguOEVn5SrAhtiwxhD+ppiBg70Hr7qcHv0qKKz
ZYgJD4GivtFo5jwSi3EtVCeCPfJbd9ltYKy7jZSH3t5cDM3+DWO/FzAffJFke/yWPrIMkYjzTDb3
vOlwJQ6/9Dn9IjBy/1IDhgMG6P/JR2LJiN8mMBC+SLT0pEKEm6IPWYtIEHebk6KzaUEXgP9KDEJ1
zwrrJoyZWW7lKweiVgGKJUKFcqq6cZZheR2hS3KnNhGzSKtoOiHgtLBmR/MfBEDPxfYt4LCh5Nu/
fRxcB0froAny6xFOgx8NOtSDPKNEc7K7rUFS8TJaMRV5rs071shJVBT0R3mkC7PSG0fE8pHe4DIc
FA0O/ssfnNZU+h886+RuiihOE8CxAZZYkHUqAajwYg4IZttSfeDkmzOW/9Nrs1oscKczFF3jV7HN
ZjZdEBcv7tvgAJR2BvTggGCk9zz9Ql+USQcHzp0J7IcnPova9cWNgyf1/NP9QdxYbKTE3JXX1/ti
Oo0HvuMZfdpxK5Jf7oMTIiVBUhmTGPQ/iBUMuSmBpC9PwQb2pFYzAkXR72BoUW1QYZpfbnZ41W1P
kJBkdaNc5wpqFuA0dyLxeBKR/v+1orySPcUI0UtMN45nnDV27e4aJxeIAJvZDG+Tg/tP+9r6ERkr
MYzcwO9RxzDqzMT5LGXZD+RZY2hkAZsdU0LkBGHC3kJHLN82p2mmH5lc4oHgg/ldLoA9vm5K2RPR
GDcQK/oCFnTjqIvMsgf1V4AAPjWFiQxEgH8A6y2qWvvl/2xVQgZRisZJvverx3+bma2d21SRcSSi
csF99hnps8fcn8lR//j2dQOjztNMWKmc4W7pN5cgouMpjk35825PFNe/FFZj7DvHjovu1/vs4AWi
CMP3QcrDu2tSOmaC5Uz3IxudBjnJtp5agTiEPIgfscS7Bh6B0xYTH5/AopJSWKstKCRUrGfjpOnY
FNuAvXJkyFVqjhHsYMKeWUbEPnep8gFOe9kB7rgXMuJuAoi4SetYL4fwA6KjR9byXUgBEJihtiGt
pzVPeaYIqnUQ8Tlc0c9xeyc1EQMWRiIptET3QYmCQ4/3i9mfp+8VWJZflOxPKjpVn+eEHVdZ5fEr
bOyr9I59eDbuEB7YcQUwJVzjduDqln6KpEmVgU8F9OSLveO5COTb93sHv6FdYUkKHEwMFAlupoMD
8YoctgXAu1sCWnp3/jzqeow/KWlq/ddLwVSpXqD9W+iLHaefsTs0Cj5ZmH6S90IulVxjbk19n9FE
DhpMzCerID1Ka+YpklJvS08nUPMdZEXhbYlpnsLqG5QCm4cvbwgVIvLn5zbIk2UDcLlpGvzXzJDm
+gUCRT0oREL6HHusaos/GiAfidB5R8urjAN1jrN6wJ8i70pGpwKB9wcTxeNjwoz4yhZwiJ4MhrgE
Ub1j9T7RbUG/syzblaL0Iz+DHI86F8YFsDGA0E8vBYMPSdpDrssQTF/eL9WVL0x75TQ6eC6JRRUX
D436LAfIfhjbjrSjjzFU3MbnoOyAaVYKD9Fjs0XlaPyFFfraRG8txW8BO6VYgsyAMLbWuHvsfN14
vbhBYhLiG9dbQ0nGSEVkgtncKgjA7LSDVuIzJArRxwP7xYtwOcAxZI6pr9JEPnTRmKwh1vqayRLD
8sg/w2bl593bEdZKW/kuOCzHTn/gswWcTQDCoTT92bEAahiUkoU8zNm5bQGCpf3RbTyWs0id39bn
mHqzR8drSr64/dA10mit3pZHXbHiLsdDXiyovH8+AsBBf40w1xTmqrLbtemHW56mdcU8DBsrKkzD
mtdQlAIdUcvBA2PsQwsyRTMNMKJMI7HnSDFM86t2+zyqhE6oym1ln2YxXOol28REiOt0+8Jt2F1D
vzvG3QeNUartseQ3ls++2XDbXCaiNXNy84DlCB70VMEwNe7069evaR8fIngLiCcirYtudkorL3HB
26s2S9qdC1Is/1Z+pfSyMaXs3JUQnfr2w9EtSAFR+Ua8Q4OmytyiT3bcUOJD6MPkzBvr1Gv3eiWW
dsYkb93EZxL2dDHyH9pn9EeBKa/uG7Bvp1VeiJpq+6h6LnEPHmYi/chVM83UdAoKK1HFhgk9SW1R
6dVHBN/9BOqZ10nYjmpIOzq6L4KZqE25Uk/MBk6uBAPm85Zhon2Pz39Ba6aEJnH9N4lq4ElnMUHd
LBWKetA+3LL6vfDN5M4d0h3DBluK0axbH08+74WVlbaSos+k8NN/dicHgO0/FeNFs/pfwY7cbcgj
G6CR9OW4oZFwTldE+bJBlWW+EUGrA4oGU9dXNzPT6Q1H151RshiWd0HWy8kgXNvspz02DPF+X6Kp
7k9uWYxF7f2BJv/Jx/nzGOHzd+0G4g+yBwMAMgp5hHeHMShIRtxyb9TYdSGSh97ZmsyBSQmV1g+Y
Ouv635JocCfnzddOWkk5s01LFprap6RYqRKUcSl7Nqq9R0LwbMPP/uqoBtmbiOToxOZ8iF4gZMu+
k+xVVe6SJlPSS+avQu6Yof0F8JPcsxi6003rhAazFO6dHHAr+Gz2l4cEmxxeSXxma7/Gxis1dgmM
2m5Jx8E8rA2FtCEAg7l9kyEVE51a5GUOiqtCEHY+XDvfTOjGevGbC79IG3Crs/vOkE4cjB2qGZJ/
N1WDCOnk3erXEK1VUQvOPmjtR2y88zycXsBNPz0B7L1iLgqST0sAxnyGNnQZZQU2VXRWnTK9AKyH
HR/MsZ2zJ5F051QS7B7ISRZsvWRGtfmbK3eyHBE93SrPbGQifkU3PTD7qvUjZBK5mQXCC1IsDgDh
bAsgQiPpzXt7FM2QND7LUSn2O7rbYzA5JCBo2fOZe9KiacSsR84WfSG8tfkLbfwoSFXMVArmXTTk
OiE/YvwtdjIA6dnqPMqJPkpQQPQU8wP576refIAsRUtOksqOgn4s/UruJ7mCEKwKlo19+IVr/6nb
YwUaOQaFOrasvW7cE/T0yIPEVsweAR0r/Wje8sPJZXcpSfeCILC9xi0dloMkmHUY6J2yjTIDiMjP
tMF1CuS+Icp6abvcIWxUtis+QDjONnLt0byNPB+1hCV5ya42hddeaGEnKkXIe4ot6AzBLa7LHwri
HtDDrqlmMlbkn08E3/7VlOR5bJFiRfqIquO45F3eGM/qz56jEnmn9xj15fjtxXVbbT4GTFnuekgT
PhhXUjS3Ddi6RJgZoATGzAvYwRv3bcYG2A94QEMWah1NKl+DtvSbwjlLZxAhgw5Tevr8to+Rt9wK
xIPS6CQKgOzgZz6oz/4bb0GZjQhYeCYUYiP4M/djqHS6r0sZlFJl4pFN3a07g37vC6ySM4e1WOOA
kpnhXJGmwfDZ49BOjh1IuIW3K1R0x8FLTvuf+rlWUEj5EMIy5y9Sm1kc30Ri2EQE+mqleUwICgSy
paYVMUNZ1huyYzZPMcRlqKqkMwvPaUEuD+uNjUfLwZu/Yh1lkuHqtARDzROhmsqCDlBTtD3U8MTC
s77E98cztK3IOxilGjpkIpoCaezsJFoQ10wNUa5JtRw/S8Ojk9moGmA37yJkiGKRqUjWFmrzpyqS
oHJy3ChIK36iuy3bek2GTyEBntkPTCg2UC1zX1Yr6Z46BKxA6ydzaxNmXHrTO8OwgLfmgmMmkIFz
OcTJXPumr6zzSrhfAEtvbv+GhbKKSaSsJOh4ZMZhyI+E82SYnwtVzDoeVg8O6Ok8o4M+iz+qJkEA
whg1A4KStkwTkykCB8fbIdPtqUioho69XsAzAsE6m0mfh7YtFAHA6hd20FxstcqVDeOx8gYQOC/H
qcdngG05KixG60osQd2tAys2pAXPdmACON7lLfh8Gi7CSLC8a/wTta1Ej1TGK+RJ5DHR/Wxfi1l9
X9qGnQnuD8Wd51KvGIfj75iXAmhdpL8cj771PQAkb3I1hn2Brb/dAnDW/AyViGAN9uedmwPHkwMs
QyXFV2mfWHTbe/wgdmanLLIwUjDSjvlJuhaK6hA/Wxj4JXsafGIfCkt7WzgKFoV1ctkmEqOEeKD5
hQfgaf+fWsBSmJfPSgzv2EWBmWSI4/Alb0upfdF9HJRrxzEogZLOWkfz2smi5b24FWpch6h6ThkW
Rld1j1Zbrsy53Syi+xNGlND0JfouR43fV5tK26qR6zOs/OqcYXmInNXMh7G2yldwxl21p65rmJfz
0gc5yRWdjOOInMVe7q3BRLqAJVM+KQIYG48WfOPgyhclsRikbtANhIF8Cg1FlVTRQdgC6Eug14oL
192UhcHr+agkG4ueWzIENeTeHsDpWP3Mz3M5qXBfRT0V/TeDXsnnjoSumK4fbMHemfr2XwsOJZCp
7Y8TqJUc0dxsnCzSUAZD6hZSOa19BTgn3HXXO0MUSxndAnOVBdSzpuhZXzTz6pCuRWjGu1+1y+fk
9iDSbR7m26lec+cwyW2Lae1zlC5k08tmFeDh3KLAVfcWwou7uWq6oh50To2BnDrvunyvf87BN5Ub
JXQip1aEo9/aJycgOnXlWlyxKxTCgh7Lq55zS2/hsyY4VWZzIOEj12Z22wHmHvRal3D0CLLivlde
6LHu7cnEdkD9vELt0o+lPirJyvFJ18FZ4UaMvBCSdNRF/VqG0Fx3u3ISUFzdL5VFAKmDVCig9VS3
JkxZZRoQTrayD8+fnOGHfWYZBg0x/Dp1eiT5GfGCDYGi0ov8/bBeAn3i41ZGw9pvWEcKxtehoJAS
PNvePip9B82O0qkA1oNkn8MgC6AREr5aGPcNKJPxaFDYgtPdzWuiYTQC7X5bIywcF/ukukjf9yVT
BbXvGMRM6PVIWBXmTHsRabRfzcOJe6khn7iRR1+kAmDrEpMfC3qeBqj5e2iFtKiNlmkiZoUZiyQO
0AnzV1cR1bxy0aG1w8+A8u7hbF4C9fQPYvWhls/RcSDWjHQ86LWMg+LS2SvQlXy5GSESGHbak3B3
gsKAiTPfrneZrwCqS/RFh85tiMnvqRx3QMXtCgv1D+ahRnIE4XRCXLfvPssHgsNz5jaCNtCrQsk6
ASDeJ29uo5Idsek5+X93UHH7GRx3jOcdvRozQI7G+0EQJai0TK/bcmyTArKTDcVlaX0S0N7ZbV7A
Bx8vXC6Tc/wq4b1MceSNky6Kl9ngMyPGKYljyfXFO1EcFWNYXJobPLqiXDoGRMeLzVC1vgdClhiN
GjIG2eCMXudJTSPCLYVoejCxCYh6BbaFo0ScqRfeawEzW4BQ79K3TPuV6/Uh8O+yZsFxH5EE5eA0
pMzc9Jd1aNoCmQqArmG8l7pYFdvIJmXPV3SDwlpE9VpYWeYvGg3DqyRW3YLYXWl2O/vWkd3CRbKF
vF2FLCGefnxnafXNXKtD6f6U/kBWu9qHsrVZWpYexD8tqVzq1ZYcWAKODAql45n/nHez4+RqwTe8
bMpXQmkGrNmNTvJ/9IAOQ+Qvbja0oM1LJeznME1a+3Dj6HgvLpAoGu1XoGM1MqBAu4yhzKch4BhJ
tAHRZWK5lma5mc8tRbayeiqb8X7P5qrpcptpIdRIKUqoYathNfTvslkMNDKQhEckg+q7muHYu6r/
texeLdWWANrZ4UsvyaiZGsjClF8GLTC/dA9TYq69trXYCyNFUAdRFo1eHu0x5U37xgl85JJAaIpH
I3Mr7sSo3/TJ+YTrIqzGB/qG5JrAmu1QYQM8BLNkDBBwsqzaT8PhGYc1dDw679Rax7tfO6iYTmOD
UldOCX1CHqSjE5lqvTRz7PPKWOhvKFl1DBr0yAadzqWb9RRkAm+TSjQeZXRpq/WOwV0IN+T65f7Z
Pjpcq1qA1yCfUszarXFGaVM+GouCGlURLVmPtdata0ARXgX/z2x6DZoBq7aGw+16FAssIq/M6MsB
RIQWV/ULKQVIou+QcnHJA/MHHM+SVk8m5dFbO+35ZQ7j1oJj4L26dwuLpKH+LykBzGWn7e7CHpaU
XgFLlNXmfiSWXZUpeZLQXC6VkaGOyCTNXqP7CsTkCzCI3w1x+OKBvT9MgFfPMNHo9Sm/RTzpTonp
9saKG7d78fjxhaThG/oyz+wChQ8jZwrYtGFx0PWnbXLTyTfOYFfW5/RZMhZQ3zcEnGLNbKEX+NR3
jPZLKdra/6Sri4NJS3YTvibbt7T4cu81mVp+HWdiDM9FDg4pt+v4QFEQrYfuRisyHG5i6dKB3Vio
pZrl5BWd11yE1aVxvY5T5UB/XsZFTCmMb1zPmHvyTy6DPvK2vD+ez3JQ/yX9mC5U5wy6kwyXY8Uc
z2SHRdW6cH7nHtZOXa9guOmtRJAwPuREJ9BgZQTBN4t+Ta0QR0ek6WbchJhhx8KPSA0sIYWknAqn
8rV+zAPaK/0VfAKYhCyTTGl3fyk0fAP/ZsqSnbimpv89+8QehWyFZTcQRwtQ+t54rBBEzflxF+FH
Py0Q7WjiA/Bh2/3y/oFUrpllDIZ1HuYE4E1wqxyOnjqeA0CgwPW9/fP8iAZmG0BLhOQzVG+d31DO
gqRZOWPAPbUfjiLBK3zCk4a56jK+iYM9vZ7tH6FeJU+Kz0a+hzwlsDrzW+kNe0sU/v2PWsi8uJcH
00gaZYy2B1QpEdfEH+VxeQmnjYy/JrH0rINOODapOZAXPH0vu9FqaKOVhD5MFOx8ybaQzi2jGqYv
DXBXP3O/yMjfPqsks1PE0GhZLpp9Ef/yD+mYNE4SR5bUcYjDuV1hQupD02jJzIlPmcB5CZWA0TcV
EmQxhKD+6X2IGsyGbS5aPOY43uzeS2ZQEwm8KGEb5AYQ1PrLkTz8cMqQ6ONwPHltLgGE1ocnhxvd
60LnW75J+ePiqbpPTzOGg+u/XJKyy72F1F2CULynkM1F1fIf9R+NCGINbevvNMRsNgab4bpz059x
FUfWwnU1KmlJt6m4Z9W54jd+p5elU7eRzZiYpc6J2fT0j5hSGHUnHEoBGG+6EDGExntE50zXlrB5
NxegQpyDU3QcNy5QhxtJAWk1XbEnp1xUeenXD0jcbmv8g9JF8PIcA1iZ/ch5QyVGitQOcloUXsbu
LJ4HjC54M/X6klAd/MfsWIWAi6vY2eCH4Eb7B9iOE8jmrSLXaOGbb3mi4AVjDShMcdIakIMRSI/b
Mcr3F7lsot4xx87hRvTwXfEKNPtI6RoTcKFNGQbY2npMvycBGI4IR1avB9ylSgAkalCiTnxrZyQO
ZZd9CS6rVsGo5Kc0TOP7qAPm8LAIv7yhLzMmZ5Iu5apayi4/JOyJj29hklXzqNBfQRWpkbNM4FQ4
yhCy2O0OQiZBZ3tf5uYCPl3i6jwPq8M75p8KoeqcAYaUVM7/BPEOuqAxY5lz51oCd/i4mr9GyzIF
gl8yi74B7pSt96Y4i/bE1zjLkb5GksiXm52lCd4R7SM+l2VMiVm5GanJSLE5Zl/jAU2sTrB7CDci
BbFWl1qnzZlgX5fnwCXM2yr4iiARqPzKR9veAZeYlsedhHNj5UwNavQrSRmIwDkRNt7MdUeJMrL3
NH1CKbK6BcPZi7b7VR04q1IcnjuOtUmrSpsnAH1J4ap6iPNaiDNNyf7lk6GP7SdQIVdpdOgTZuO8
mmxTTB2Y70BuSl+cag2OCWemE/gxsTp5piqHY5zUvGU5XwnnZOGeXHut760QsaclB1oUKiwlZ8Hd
Dy1Sxl2cJrjiCBw8/UKjXt+3YI1Pe94vh6ZYylXn5dzLvV710KbAipMJ9Ps4V4mQrGM4cvj02ypW
xBHSFRCvF3v3JIMEfOKfr3+LQ5XUC01X2Acxv652aV7GeQQh+yYq7Lu6a+ijWHxKNcjzSVAmRy0m
I69s09mi4vJ77JM/aWb0VCFV3pzEvLNWueEl8oltSLyrjH4pEo2i8e5ct8xP7Gu9TwuTjBPsHFJN
PmMPb4b346XDR24VlzX+6ddcCM/qANYGCO0/veu5nHWwcdEb122KbKmZv9sb7esVbH1usmrKOEnL
zZIVRrBJOQRAFEisuuX+mhbdltrsow30IQs92iUIrZYX1SlbRGxKvV4tj2JhheVvZdEmOOPRzAmc
VmS2DGVpVdn/nWI93BxsijSWrXy5IKN9sVJZN2zJMWK6T8AawiutRLDTOdHn+a7fQLGlPqKotyP8
68Kt3zeU+FpynKvqpfqYJK2zBjC6ilyYTlXkYLvET0Kd5drx3iOrE23gPiyAgSLlomBFRAiuAGqO
JhJK7zwmK++ZP7LfVNgJyvb1iuzm0/jGnzW//1LAvUeBNVGRrB4T//AjNRELcfwaDdO8DuDVwRnu
kUF/MgExZxw9Dm4K8eR/9IV4uU30LsZygUSzRE40T3YAk3IfaUu3UkrRteOlJUg4hgLmfma0HoMD
pySDxqNethLFn1K0saBA6YJcGoXPvhVeFYrxTYTP22swU0Z4hNcyeSNoIYMfZgtCfbhmiarejZOF
Ap3Y3xHInfRA6nAQOZP83mlBB+8Gw89NCQ95nHMOK8UNDJZNf41EBSQ72kpOshygYCk2kaLRpBbU
VA/uxnypnGRDXCPS/uHbqTBBmpAd/Sf05URz2EGLo5yVkY2U7EWQf6whVOCMUoN3Q+zPMwDh2gdh
5znxh6IuvDsIKsKf2bJKgSamsNzMWdYDTac0j8XsaU7Xr85AyUxL9X8KBIeuHa4RpvzydgrUVnhM
ifFYXmzD0BTjyMFcSSVCd6zzEtT4CWF8cz07O+fRERgSR/EN6Pkj2o6nfzd7dDyPHtCP8lbFkiTu
exjodFBhXl5tLbmOhKJ2KFjJ3lkr6acX/45FKi3snNaTRzbvSHjJ8dquwerr2dMoLvxOnuHkNe86
g3rI/0yIWxZkfnxKSs7fRjZXEUrkSDz3j3Kl8xrvQXOQMrOmzhPK1bj6lmle4qJIK2pVaW2w6itC
8529FKNc/5hdkA/ykkuQhHjYdlstnFZtLBg4Nx8g+7CwFlIBnnuRUH7GFCT9Td/y/4cC/jUR+Xkq
UZQ88RPNvFpkS3H7V7+3oeY3ST3XKA1HCwQtI1Cph8agLb0J6VxMMuDLrggPir80k1Zi+eG5gGlo
nKFnBlZ/tHr3nMYa7OlQS+elXJ01XKTuexGUQwf/LrWotoAHA4lkzz+RtYoVac3Ff3g6cPIS47Wy
lOMnAIiuL2QBLmsrK81JWXdWGyB0vnRxLhzZScYTXBAHlTIQt4K5sFmFBPog9pmt8wnTKXqaYzsK
PgI7kljjiWFde2OPVqfYa3KEgrTisvlNu1wx2oFZZH00KqJUuu9knymdsLEqLbNzttuV8HaA+xwe
0Ixv/UE8WHFGS3EbpA0QFh35IPwW/pwL4MBNkYigV/kE2rNqHDH3EFIhPino1vfKjLurKAtxzqkp
Fx2d58g1I7KCJvgrrGHBA8Tt+vz5emb7egXnk4ClkC+cInJuUUKeYzJ/Nb7wqD0Trgh+Twq9jegz
RWy2HQ4dcW+K46128D2qfpm7ryHxL1cBtPjzGFEcQPDjvnKN+iMkH/Vz1Wg5OQUWVuqfLicksWe+
vYq3fHXVuYtEvR4ZID4gp2Y0p+BBfsQM6AkVODTaHJd55LxYXrTVPPfaieqa0+tLMptGT6EHVRcG
zCFmyAvczMGxoGJSFTuNDHV56vOMbjFsZ5oGlROEEsOjB57kuMQDDwvgzOVQbSj3RTa626klJl7a
S+uhqZ0NI7fpUMmoi48BfEEmXPoDO2fIJazOukejmq0u11U40Nei9RODyTqBF4sURldOdE+YMgPd
2NCmr730rAffCRYR/4sr5CPWnJ4TocyHT77LHNffCjTk2pUIcpiBWEU/p1SfNmKPNFph64/GaJqC
FkZv2iSTMwqnkSJvLbMhCWYE8jfnEvgWAzbkLJdF0SD8k+akk1B2urCavU6jlhhkzAS/+VHvjNVE
FkhrDVLRYHjSx+N6ScWVvFlbER7KE/od6xhuZz8MlDC9IiMYTf82XB9tKe7c+1GEfRQc2yqprJtv
lNKRi0bRgKKNCfG0vOpVjqeyHDFMK5PtZxxnpV/T5kOCBFCgZTuphQzgKFw+YdNLsPAgfoki6FAE
y8k1cmcvUaIGWjSnIATtvgcEsY8J5VG7v8kU5MhEVJA2iFFnmBY+Gi9BOTf9SpctFTh0YRPI5s+R
eG2X+8Vha/pQQPQmm59+Ru858YM4lHuBUA5CjnjOwfArSapdw3Gro5xmSssoDxfvRf8y9yQULTmM
6OBl7i+fqv8uwcDbfWlVl3NGeKW6hS8uwfOaz/ir18zvBBa4M47YIVR2DzaEfrT7RvWclEpMoVuw
yF8JFewaPOlv35oyrE6yzvDWQrJtOHfu/QlYkFuy3yCwJMLKkj6e7Bxq/Ek9b5MLZ6ZN4XJ229X2
1n41GoLYRdmAtQlKZwKzulc64RQruTeIijHZnG+YeQ+HoREdEBCNpmtDQ6OLSGXKVsOVdho4fCBc
LngbPsg9MEiapmwAxWaPFhIFM+OuVIk7LCLG9nBFuRvuSLlqhXkoF8evPM0Brku8o2uiJGbStcXH
3Rr+5MZessEoTDxSCyxqlYxvF3m9C04j1qZSUl4tAxSmWYO4CHokFUV/Xv4wsdHeTXLMksIweQih
YvqlA9h6sNZfrzFGJ4KnPY3AFiDZ2bLwuxuY3EhaSAGq7iilU0Ric31rFuC8BAsIkc9s56WWB8Zc
LdvkY+XYwz0mKTsoamhRHuP8Nk/h5VnuCk2oQ8t4VeusSGWfHCs/wYM1LExq17rkEKm6vJTAOcvU
/muFN6U8vEIl7DO6dUlYHAIVuwySGYzda06txa4eBS/5a/zOyh+fwJs0VcMps1fao6KdkcIMf4rQ
juyReDnZ2BrEZlynOu1dWiwBMg+59OZMZpY6jMNtzZvC4RZcEBDTWtPOSANWbafpKseyMrRtyHZe
0JQ08IHQWUhpOo6q081zoHjoYy49+8D9JFP31YONy779nh4/quQsVODPalnFTFehHsRjhTGoXnpB
pNq9mZ55n4MhjS2CyDWIuQD4Hj6VyrZrK14SZnEo/CVFGUdZxgvGTM9Fb5vZN+sOSxeMYK7EmIOL
O3TSzC0zsSHGQAETYPZgRG5uWWrm2+kuyUjLmNFESIwUlVvUfLwOFGVegQJ7N/EtFUc7RE+XcRLy
HqFqsMjWVWvFbIijRPXSrqU8pmZyLh2IbNmhYPGtBDs/5HkbdxpgrXrQvgA5nwHIx0RPfQbhvSBX
XiocxDepWlKSRlX3IOm6DmQLWHtUzyW5s+CQW2n+hZO9OPc60E4XGMvNkk/hBGRjYC7oIO6ab2Rj
GGusPRuJPDTVLqfdsyIymtkLhlEPJ4u2Z6QYgXwSgYvTb0ufBFbm8bjsi10evwrN0etIIThZNLRr
zn+IDa/wRSCX6UTemoJYUwt2Ry/ea64h2+ssyoVLiDOZaBJiy9mNiQZbP6BcWMZWcCVpbmPSc6MU
X6RqEVz7qk8xBLUu7/vwOCytqZsE/am4ft1dogmeLSWfkFIDfouYHEP696PI7HOtbqBt+uHN/1Cs
Zx5ZTISKlXXu3NlGwQkjq9SLLPZWH16CjJRvo3U1qSjtAUxLhPAwZCMHM/kVkKpQItCO4Ha0AVxT
ez1mfVnBkakrwA5XGo1yNvj3+Y+6N+1Xb46ACBzmhkmg7n4j3OHmmMdfre6QmXzFRoZf/YL/oD1U
BS0ZxJfmYvVkMLstt57IXpUDDGiAxS7EdCYGZOA4kZcH+QZNxjRnzPTiHFH5RvvcxOULFQVKzCOJ
1l2EejR9PxcluCcketz74bEqGSTbY28YH6lRicmAI5mdu7N2ZgVq9P3OwWYanzxYk4AtizA4Fwao
wNFXK5yfDiVjkOcobq/hUBeATj21KUmxIR+ZqOr0JFn8+e9GLX6N2cefqHok+4rpKpGLKw7erbIi
pv4cIYrDZeLULUWIvOnYs9jiDyUMUjpvqUs9HItK5ls0swWKEOlk2WH/3zmaUUcfAG8kxS+59KOc
jruIJclShSqVF5Ol6DOQ9hGpppOIZ4iXh1y5x1BwzfPchl7XJHvkK2nK8/aalmiTCp46IEYvSBjJ
F7zNY6X6hly5ATVr6Hsct8BBqir9JNXxQDbpFf34Pen2AICjI/AZavHpRSz6dgKjQXqLAwhVgFXh
H6vkLK+rq+86oGmD3zGF1vDWQPWlC82G9ahmDM3HB65+hSG3WgmnHctXA5NLTssbfNr5tcg49JnX
GF6BwgUua2mZi7LdsOHpZf7poTfEh/GthfrHZgNuB21jcblXY9/FEB0O0pI4hz8+KZPtIa0q88lW
uxTEYQAXleTPlidwH8GD2En3a04gHo9BfA5zYuGoftRb8aL4Eitw2OJmRM7udXdmdqp6dBcwMSQk
FCL9XZfoIaBeIIwK020gJPu/Wlyqs63oxEbG4gSeGt8sz6wckv+0xBav84/4djPUJTSmBdyWMBk0
0x8p8YsGUCRXXCOlSqsXCwa8PerVR6EFZ46NpxfOsHcmNuO2Kt0PaWaeQBvCIH2KUpUGsJ8zalLt
u4vRHLoL4Eno7B+Sf4YoUYGjy2/pUzycVjHFTNGW5c1lop5NSCqtViyROKJBzZulPuNvyyNwIZeJ
tOWR3ByJDiDu8ZNg860cP99nVQ2/3Nm4FpUv4KB4OTuMLb7wWUnx5pOKfnqSoVfKsumy0qs4FH8K
CGhTVZfhqrow9PrKVe2azJ/k8cclTJsGkKHZFzBZ3iaLT5l+2lNL3sF4IDT1cBfcOwH4+eDYr8GK
oyWHcivQLfAWlA6tArDN95ySsGNCJCXG6nHoYv9kapReh0g4iuwCwmhzSTzWhz8Cd0nLJ6YTY+pZ
FzOGS7pGGP6dGfBr7e1gMlgjmON2wyihmHtOP7wl4saJIcJDhiI3SYOhYN+dQk9Fj5uxUFVwrNoQ
3FOtEtbiZyzVsu2vv9BO5OZBpzhgwfQYP0DaP+FfmoeNE/m5jD4MNHJ2/HvYWH9WEj6iUpzt2zKP
72jD/rP3YLjFHtFkQQuHNDCNb5w/Uanu3GucugSAr2vCx4y7jRV7RqPXU8ghfeKSz2k79CzU7Pmo
Ge4u597nmuayPxi1I/Q2gRglXJx5RhepGfdni5vME3mEjA24LQj2fYoD76p7XN5/PmMK3uPMXInc
Li8XcU9FDMfsbDYIy/4tqMeTO4YrmTdlO2thf1EJVPCitVY9asZEW2JNQE1syXQ7Nzt3bc31MYoF
vKY6WasSsRZNx4GjmBN6eDSQ1ULMjNBMachTVfn7yCXWutpwCRilI5CAK8TJ1/oZ5afp2DkLA37B
fNf2UNdMtcMRg81lp+bNeGNMqssRoZrMP6EaE9FA96z3fjQGmbQzaq6J6VnCRoOxiTSQ63kI/K6V
BTo1ZuHZcDEtvjSfxvc6S6yZvz0ju3PbrczyWCJcCACPzRTQdEVIaoHLr+SKKXUfHY5jAy23vx+R
eN5dWKfDG7ijs0GFdgG2aFWgIAidsk/kUd4CWSN0rQy8Xu0NNPAE1qRZ4HQsh5iqQ1dbLyuA+WOj
FK2jTKQ1o7MBC+fvx7QHxd9EfQTrYTs/9oSDsNAXxFUO7Co9umctKr/N0VTIXzVPVQvCfiiJnDBs
nveqoWZrlDQqRIDaofTIA1oj8q3nv9ZTYmL0lvng3KyQAv2bZnlkQ6OB/N5NJiVITQjub3XXF+OC
Al/0uwh8YaFE+ux9KcwvhfI5NVF3nR0vWKFirxYfPG9jRI5tHjZdSJrYh6214da2DnQFFyTIxU/f
jySIVxI5FN4EioQnIH4KxUxQdMQWBaTykL+28kVLxhEIXGnqlmNPCZ/lbGPgRrDpvR/hl+dAQAiq
16I/Sk95RUIQmqkEaHPGduYzQJfj9OH9b6fZYi2YpZlZPmw5Q2bCC9xMa8JDyssNZUaqnCvQOwtE
99uw8LYpYDUFzSaFeEbMUK8Wkwb4pNrjsnQE0yCFUl1VZpNhnGbK4l0PCH5QxK5GGSlg0wQlpD7V
qdYagg4pEQaf4vkwNIcM/zDTnbuTqNw2CqsCkvXDZMRrys5YzIL8v5hCj+xnLKYuHfR1R5tCp5ke
IjlQJRCLGWr6M0yaxYZFm4ED6vP/FlQGz/cKluvVZ/hpEvgKtWZ2yWqIo8auaOxbCDKtdYGCyf1W
VEw8BngQyczs8wHlXrlbCaQNuLNZp2NPadLZ2W/ckHxoroJLromtaJU23bRkuM/eaNT0j9RQQBpz
2/zaPwHUjeeFMM0s5vY9I1HOpY0m8kFXVSyzb+UD1Mi2oiNbvvYA8uQq/IiKjqJX/7qis0NLFNYr
j8mSNR9483pTC06x9gmrXz+R9HDpTgvU5tl3ER0UGU1v27Pbby2k/KQx5Xe8UpKCtvlYB53RUjAG
8ZfZEZ8L4ZJvFrzrfy5agLUTTqRPFxKCWbbcCudVZCbRa9R+wZ7Rnflq7fvVLWAEWclE6mCzp4yW
Jo5huMx6nAUlibTM0LUXeYkqQiRekNFmyh7KR+lpep+mTzjdBdRDWXxI1g3BfknFDbK5qFgkH8P8
NDrHZCKT6AWT3w3TaDb05TPoHMAQWPvMll+K8o0A0FwIHuaHo3NMOIahMSIdXvqYLB62ydCVokTt
yYWaeDm48Q3HSGfQFjSCSSA+NjiTdzdjKqghicWQJNPJpqDgMQjlds3tnYDw4ibTpXMLKzZ5oPLE
GSQoR56tdJy+NX1sbP8vjmeg17+C+MaZaSjUgDDgKJ0zSkGmjNpMjWLk4/vIiCMBGQEbPu/ZtFMR
+UR0ATyMRcnklZjHEWwSZq2RrZ3f7JVi15+gNs3p2xOz//718y7mM4c69Lvtl+tNmBKlLcpbgAVd
HvZWQlQxa7lp/eT93ETjvOv5lVJH6PoddtYJtzCcE/WA+EDI7kt13nuRMPRV2cLCP9dCaCUt344i
bhnWzRjdI1V3FpBY7daiGkVZbSqgqYIe6ELWgcSi+T/qTVLtQ3dJrcnNvXiGlUsjD9RpaDs7A1mC
frznrEyTcXgkjBA7R46culi6m3VZlR36Xese31/8R1Gy7cNED4kdmdhtESe+Q2WuEnRkzGiwPYAd
yOX0uyptQKiCMogmx3Sbk+2it8L0yoFgqJg51A9Pxcvm3lVvCoXOOkPNt8yheNJYZpfdPOakOoHw
GU0NHcczxAhuofr9zH69dj4YbjVe08wnz13e6vq+/vm9W6K3qU8KBtznWoVt2PYHjfJUb5yiyO3M
tQnN4f+2SuvcLlHE0I+3SqAZ1TqhNsLCEf41IuBipQOX+XtqugaihUnFBi9pfYqcyQbvJT2sMJ5V
c80NzbOUklYPuzgc1xkO+wFu9CQOagVGIcqHsxDXvmFa8INS7a6DFcy4BVw2fAOzDt2X8RPOLMxG
f3UfwWBMCQctHxoQBsfgL2a1H61FaNTEvWgvy8USSkpJlpoIQAFefVbgoQOin28v4FgCDG70/4N+
rwdgoHnL42i7tw8g1ZlorHHP6Dr9t3kbRV+Yuilm7p7kgd/XfpS1jHKC3MvSnJxhaC+zD/5jhlrC
nCIaFq64q3XO/WNCRhA5CNQ/dlVmxUShXB2rIlMdHu3+qwskRsOQvGFGXyQsFv886GzZoFyxHUDM
SeeIxCmvvS2zN9ZbZ+YG/LkoIU2YsdihiJ9BOxS4AWnr+lbF0CSR9qv87OfxAFSdF9cSkWrxBC51
ajPRyjcjFM+ZOXDYnhdmQiDcRTpROSUwoW1qC//xluT1oZUccLtlT/6p62xnRNoi8dI4Heh/UCCs
AKM/ZaTKGNHNoq0uA/zAHy/9XdWU92QUx3UNuMrRjbqMreDQuiK2Ku9XN7LZHNbL+ScGfEKP2HWk
LRi7Ok5mPUSf7mI/NFexF+LhtjeJ92hCEaQSA8ObjxQ2lKqQ67kAT+lrkO7/+Vn6tUU2UPhBunxp
bDDx8HinzxKzcjuUJVQXC6WvzCGIEwE8jxrmIlnBt/UInk8ldGwleRqEVLkHhwOEAOPOztytB+9M
ux3tXTvcjlGLQ5ZwWhRp0ucNY4t+qai1S9OOFDZlHHWHNmTtSbT8da6WDaWBseU61XKuNnIEeSjA
JhcDfzdkjo2bnDyGpZBNKnAgye/tVEh5xhsLtqyZXsllAm7OOd6fwfgxKeaitYh+1mjY5JytPKe4
FPYcOZ2SxsD667BlWQyRJipO0ZBCbBzNJfLs8c5E5CxpyCS0jG6r7swK+/4SJP+aUILka+/Y3Btx
2sD2HNkucwdIsT/pcU43v6qYqJ720O0nA7EpjEf+k0UtmPBd3VjpaL5hr/GhjLHfj5RAfsImEUc9
O9ei9vUUM2AbwBa4tFgUkTP/2i8P7z/UJJDefdxIQN5y3MGluSfOls891KwAkAtOTHwzvxZSRwIM
YRLwcZqi1mY0qTE/J48uge4DEXL6+3P86iADHaK2qdB/btDwi7ab9o4DDQ+NgRaLt1AWEHSwnm8V
9wFX12iCM++ooPiJqLp1C0DRkqJHavihPyggGs8PSiHcdOpB9CP1BtVW4x9j0brfiYkOebllGxbu
6bS3L6OQUYohUy9tgHzI/FCiu/Zm9IQ/eEA/uQWKwW4YxiKMXPVA8Ameqba8YNV9pBPKZqFw1QvS
aZxnl8hlH7UxsOTJS8C/hkDtFmkgbH0gHAslC48jph8IYqNsEFCsMTEVW1r7pfaurBUvLv5Bhg6/
kkmD7c6BoXDGBNfTMTMONPBY6syZSKoGlZFlVDsVmWnvJEa7EoaqthMb4m0IG1J2EC/aBIvl74Ep
BzLwTDl7Sm75iOKFJOzSkTLKVvpoZIqMkvBur+QQkUB4AmNHJbwywypj8/ZPx9K15FT07rmGG3Qf
HkYbNmfXVLu5zJ3104KBMAhgUjV78dvBJUL29MaT6lyl7sW+6Z4Y2XFG6Xo9RhNcfAcsdEoJYzBx
6DVleOLUk0BPNz0eKrOyTMRduYu8X1SH5/0GYXnNZ0ZonEslrcBgiR6xIV6vRkC5g74NKFC9V26B
ftPI6tJLvunAPxw8kwToTQnDABvU3USzE1Lj1t1TPf9m9bNrmfBm+8fFg6WI7z7iaDDnla74XU2I
KPQbwxRpHfWcpkGkUiIxG2L0xC2WS+m98Hdmfwm0AJiPIgjwDu059vGyFrSQG8s6VmCXcZ3u8QVw
R51tL5ILC7doVfMW6lnVZ6ubisWXkPga3MEwq4832SKRWWWMP3tP/1wqpVXwLRwj0YCdbMVW0YSD
caYlqihufeoUoWMvj8+fqJhH1P9gFys8H4EzP36qCHPPvU3fFC9QicNlHNyMZZsGkm3moHccgjsw
c/JQeOiUDHOkv6sTLeafNA63xXl504P0sEHzLyzj0zV7PYWZNk0TkZQo7UaeXeTnuyLiQFk5fO/m
ii8zIKCXTxMfKVXCmGEVVmwb+ux2e5Q0vJG6OWkJ4aBBkbodNlVttYCUhnLYR+7VXmifGolegNZy
5iXizqnKjKXVEdmvi56PoSHTqZ8delmm81IQPcKt4vk3QmB8/Ivzhjc8JxYRPYxrqI0C+rPAIGwL
1pDh0kj3XuNb2PFsGNy8+XMImIXDV6H4OoiTi006bGQ3YSuNrphLdpdPjtQDNYQOlkr+YeFg5Dku
vQIL5Xfg00BDauks5hA/urTiU8GbQEhi+JC0iB91SyqCwYrmsL2Eao/jDpjdl6/cai6nIjA8fcYZ
5xePZ5+kIhj0c7xxQmr38twyS/zVJQIC/+5TdQdNBqtZ7Y5O0+32t5uC+zeMwCCXNVyDDDVCDIW3
41iFpx2fk91FiBhdY5HM319aE7iOTZ9tSGVUSb+peKvIVurkdDqkSQXADDbTk4GuC8sDLER8IJok
luwmEZJGOhbvLSdTXsOWhdQDW3CrFA2+55XLtJoe3A0KZ9fS1E1UxE9c/tB9Gmuh//qQ4J4ASV6F
xo9llQHPHmsTQKnneFMcqjGfk2g/FwkLibJVpqfY3uLx/3i1EL/wBSTFAjAM/4DZAXFB3AGj1iFT
rpLwt/fZ7QnPBAfsZt1DSDbeMFP9Q7BKHc1Jdw5gBXfS0wvAO1uIY9LxWmOxZmmHTQFQiRt8154x
mRl7+b1ID4LXAD+wOT8LTraap3gRSJztx1XQZlAVNaG0Eb/A8Ag0wjWeDgOY8BMsRNIZs+rQ7agt
gPu9vdnwm6ld7Xwqa3/kXSHkxD+J0wjlm/5C8orYPefVexUUZ5mJ8YxeWozRsELTmZv1kZdmv7td
PO2qPvxwpJ/KxL8r1e4jmmvpAkgxlByObI2VypkAgocBFHbnt7HZhr3QZesCLrP1zx9zm5IB5NKm
ov4PQkMsgIMDlnhUOQI+q9u1m7Tg+BAxfw1d8zAW8YmM5ZtMJ/VX+jGqzoK65vh0cxItAO1tnBik
fxrHF4iWW5fnTwOlaCaDdSAWNp7UAtDhJrtVBxJO0eb40OFwPOrCvj0OmGR5iy6aZrmpXhOiaHSz
EN1hjwvHk/+GTYnmvAelBWsqbmHafoUb8fAxyHuhIFL8LNgRgJCr2xVlRVHKkpJZ3t9oZ0h+BwjZ
PoOPWIJ19OvljQPgQjDYoWIzRht0uxzwPFQJpW/2IbFvkebIURWzQji5rMSYEIQg8OC3bt7OjZ4Q
C3V0vD+517pu67Qd303hgW9o/ZBhxvTF5zGBI8Jlied8cahyzxIBkq5AQo23JdZeWIRg0NCSl+zV
e5EtLO+yzaeAnCeBSkQM+F738wsCZCOHSuDGGRDQVjrKTp47rGcC0372VGafg0UYKOWaDdEGpULT
K8poLjlrA1BIdMrCGkbh2tFly/SM7WldUpxMtyO9++70SW1KkYxfgfzNThGV5bto7EqDTfAXd+Q/
kz8c4zppWL1e5PN7y4z0mSTcEEmqf/GZh/xso17PbFGw5YCTw9UBJSuPMNgmlkNUL82DB6atlDmA
4mDsE2ysIJQ9ZXjTewUHt6DUCd+qYIg616KUTxJQTxvz99nMnlBwL/mwKSjyn4x1bLU5uM7YInnu
17NxARin5eyrP5buFwwTzYuvSgAjaxPXZv2vk78K0B2MZ0qHtB4meeNK4hwV3geGSA7+D2UMfi9B
yaz9tDmntlX7xwDDRXCJwfcuTWGmoODPjxFxBdwO7EYLboC07B0ZMuBTIQN5GoaUe80KvLeMam+4
oBdttnxuk3nnT/fUhamPesk0s9T8hxKodmgtKSbOIhcn7qMoVeT7agakGvMX/RR4AkSMrX8/xhi7
m+IRLdhTpCo84oyaVcOrs59xbg03dokwge9Kg+zv3POxCid19ZNMD0UXolf+2LBzQ04HPRp+zmFv
1zAyymbLcm0BFC1jd5gQKi6fJNYcwx3C/LqVPHLMXWSNFdvuaFryhEZoHYNhLranuJG/FgUBrU96
EnpJsfN5r1lJmv77L6ZVyEcmZrBAxRuBnwEwd05WiCn3lQ3pJ5ocv56kKBG9VcEUxAl6CjpRMwK8
qVP79tnfDglcSO017vexkXsRE8rQu/rzWHb+YIRl5mgqUQwCscGmdGLJicDuMwIkdsLubWGU6hiT
Tpxd3RUnDa8EF16q0IrLnUxZY8aHBj8lyFrQgczsTFeUVPRAr2Dzvf+53jcv2XPZLAKqNSIwFBv+
wCnGoSCg7d8DPzq2HPLhwI2ZhcQqvpSSherrKpqDc5LzIlZxPoF/agiS1OYCZFLCPvWuFVfRfYmD
hvAu5yOijN9ZagkvBqWMU7FMj4G03ir/QPmySp4MMMYFsnfZLqxgGmOgj3BYm0pzNqXVCw3aTd/5
jKvK5/s5gIyu8B3rd/L5tZrnqZpkXGWQ1q8UsbqPqxTAMQh8vl/qazrTOL5BvevEWuPs6vQmYcql
3HrcuZBGyAfxktqGcL3GKMql035kGRr4HHjkVgsRPwOLU7r+7hvpIDfxuhcvdDXW0lkJ8XUmzvV6
onTvu5y8cFKUWCeLBwBM9Nw63/cQ0jT73+9G1nkxZUAaAiLc7ky85ZRnN5YJFFXRnAfN30KSW+1P
x/XcaUyVUxD/WSjzSlzYAYjiCGvx7CTi+3lyKNwgeZwH/Pg7FIzW4X4iuAr0SnuRPXaN35r8kCrv
eNrXfdZK2Dc8FwamCPjRpEdUd7qDwGRrnj/D4lWa0oGOMu2fn249sY4SKUt1c+mkC3eNj3PLXDew
tDub5KRh2lzho5q7mY/FVIgUG1ujUjq2hTKowrMALP+TZRX/PqV6dQ/Z56faeWmWZXZni117XYRf
XZMrOolWVii0xaICcMhxg1KkSKBV3inHQcwilBbTWloI+pCE/cC6E2jL0XieAhp6MWcZbzPXzPds
rn8aN7AxZ/SsEBlerJtc1tr7+rFDa/MgRVwVMMGB0KMrmQHCQg6E/NEBjY7LL/ZkFxyaULFKfP6F
G2h0jG2qILK/tHCa/POnl92ydlFlntzQAyh5jd9D0I1F8H4k8Wn4O6vfTn4p1ELEDpGlHq54zpAT
kP92pdrN7ZzttvlKiCt7AnHD5NoVFXvC9td0gXWJSarRvXZtmreMr/gVy7CIxS0dSTI+eIWe1oY0
8UQYIdHsVFDWkmi0/tPGMY5pyZfonW473EbimYvAq7gRajR66D2/gbtXq9Td3AAvPKSV6969gdKk
+yj11Unzuz4OP2AOo4iQPLitWuyREQ7S4xhq0op5+D/5UfojdOmDOwnb81HMZRK8RPX4rIR6L4af
wQIuBOyvBlmU99BNGrPNcM/GOCSdv3caBGFeE2N8/8Wrkwzi/NbZmbNSljE4q/sR40XoMid2GZqc
9PPIBxu2SWoLkj1eH2hDglgQtxyspYtsg+Hbu2rrNZ5YkPOHkv+SvoCBPNSQlIlWnwPzdMw9rIaj
p8oxY62gz6eoOXpgCWwbdG+BgFyuqoZC9DMKUcHbN4MXuSJYsPwdpH2L3LMq5acbdyP4fQB6FfqT
e5K1ovM16nQWvgEwq19mjIXYIlQ5O0Gnipeq6JsvRfyHAyMvefN/dbT0umbOGrMqf9idMleafu/8
WcpyKX2jyhn9sJQiXhkC69HxnDk8QDMYFnKmCvVM0DdG06mOBIPZxzZZful2HVAYYIt6f/zT4Psu
+g/Jn2GF9EJjI2fANOvEmd9NJEGTAAEUoabQsAx3wAv8mRdWS8grjpJFbCmWplRZQa1sFEuFfhI6
6XszCZeWpZGZi67kJPwy+AdfZrV+ORUYsPMdm3K3Ezd+/+9vhzw4MBTzJsvxTcmkA+o4rsIYVu2m
VhV/EFSi/o3rEiNECBG9dFwKplMNoAECUE1qkLC4+pRL68q5Kp+X2vPJ04HTX+PkcysT87JK3SNk
RlS+lhTKHyIHK3bz2UQBl49ns1GR/f4qFUBXN2T70rwy/yYuSrmemXAb8PXDKg5XmaNdbjSw7VcM
d2va1otxsN2UkEHxYb2o9Inj/QVfOQmV+gc32aVKqi60XeaDI54xwTh8kHD8YckArJpOhf96Fb3+
NKu/qUl0YU0df1LvZjD9moI97qImQ8pcgy27d2vP/H4ASIIa/6gU+8TBH+NLl4ILoj5srlMOUilI
ctoHLeD28qA7OXnYQQTsxMbCJcjc1SA96T2+cfDCcHqWHg4gvQWF4YIpquxbDr3PlsTR4oCLqFpE
Rj173A81ENeDjzbviK1rcEwXK0m300LiXCEcRBKfZEjilmRYWjarI2AXLqBj/46l/u7MvZ2AOF35
1m1h275cIdV07luK4RS593N0d7GD8V9UmwP5/HQmeYZnK+0mZi/DW8UcyN/uA0FXjvOmKdlwRfiL
pU3LrGyBbW6o0XgXCU0rHBezSs0EkJR1QpHLYrGIh3GmN9+2iCbhE8J5wXyYx2ozYxfVnO/X/3io
rW8eKYARXByGs7WZDRY+RtzG9uyAUIhLHyhXjmR9VHY5DLo3s3B1Yn/aONiYxajud/E/X0zha5sZ
wnXniMN1Z9h1x/7dzn1yrhC1ngBw5n/a8Bk48L1BdRkBiju4jDvL0pw5oDu67HUSRl0aXWkhiVeo
NuoHla916buiX6zWjyaa81StHlPVTzfrpIjPXo+R1HznEOQmMe2bSt90799sgK4fqBpbKrgc40p4
maCOr9lKFClbMcIQ7bwlOtzMNOwgyg24cNZ4+ECBYMF/6WXg3WFQkVCVZQ85RKKwSXAnVeIrnXkJ
eFZi8JJTIMUrwaCt7qGcNjOkYPQKeqS0n2qLVFgok4ln3eV7DNP/WNLz1eGXKyTcZp1GLEV5flGG
or9wjSl8pGm0W1ZxLfkePae8ZEetxe0FMTunh7T5rZUeDFttLXEwMLzA3WIdaTyOU9CylWkCYi8P
lqYaQWFw9nPpivkuRHbsjv28JnnnC5r2PttKqMMQl6QfGUiPC6AUjSEiXn7Hnfgg2qlGgQ2qC6qu
9HDrspR6FCXnQxiJZe6b2EZMZxbSy5vCVOA43qXFKxG2Wq1ZROm/g4PtndY14waNlQZ2Pu0ksftB
NT3lNy3FKzmRHQ+fRv+6rRIcq6hEve0IHFZsflZ7Fizdwiis+1NGDnqQjzt0vINO6uM+jBAUBczq
w+r04Ttbxh4qQxfrbrgm5Oeh+Tpxid8tP5LrwRekEPaZCZjR768gSTZMJ0WTeSqTwES+PDStxdw1
RNtP907FN+XdrU8wuib+oeoTqivoZTLNj1SJcYDWIyx5x18DXUnYUws1z1NPen9M2FJcBUCsg253
vFMkIoMAHhuBrzVOaRfYlMLYrXkRt/Fsn3g+jcujNPdllhpjzQbAk+6R2/f7SQ01I/VqtWBo/bH6
QBZz85MAuCmdRPKqMYnXjc1dsGuph4X8TgRY2pb8RjxmiYAAz+60wYOUrOPvwMnUKrDk7xN4xNwL
WlPjlAEu6my3Q7lfOm0pPkxEoQE4aRYq8GuL8poLiXo8CIduEfOriMXn3oc3/ICoD2S3UOaZKXt0
rP/+bJTBpBWUAxakQD+XcmiD7TKVT09aLFuBfmELG2PNv3qM2vr1BlumF1TNzBfHdlM4I9oonjYq
ZVRz/hAxN9jO8LvMi0SoPoERxO4bTNmYJddq2h/5gSaXeLOBZMwoT+or1pJbCHEnc2DhPgPy6xx+
/WWUhBslC1VOvbA6ZlKXl4YqnzclcwTgGMqh3Oq1rSl0Ra7MrO+M8JFV4FEv1CYDqZMMiiGBmUaK
TTzwWFGIk8vR7ZWbs2xvRNTfniYbztn9V1lENJXH6tDJvaOBfZfJwTrO41EmxnwlJJev5rsUpP2J
VVHTEmtP8W1tkp8Z2vz++yUGmW3jGfYfd0oBL95q+g6mvJApYRtsAzRDLoI3NhTpwN6dUbVAI4zw
B/nAwl0Wg3vrKyQqehJEgAY5D/wQ6ckSpvsvFqIcIfa+dYt2N/gGa6Ds50pzj5+8f6cB57i0HBAk
zRnMSYgZctiKlvjoHBcDWQmk+OJ/CvUaauIdgmMwBq7Ko3p7HUiw1MnYOpIOnyipoppDqi86G6bO
LGjwjg5p6h9aGQtHM7Wqs0SrYbK6NWJC0dvwEMid7vlNrtfCR3SIfPUHMplsIC2bXIge6Ghxl5O+
bjJvwkYOpfKxPuBmC8sxQB6RkUJtFjgGBZlFK26hDqEZikpnHSZEnTCFCPP75n4RwgdMJbonUiG3
SVbBljpRupvRMi5P2KWHUSX9kgx8wqy0KInefaVJ6FuY96s2QLfuNkuaPiX5egYPoRyh517+Qmtc
CXAuyBNevPygjgq90TUUpw8Cz3Bd2GYTewZMsLrIOoBoiAfk4M/mYFQG7XIiRpWeWojAev6ou2PQ
ClQEXFO/6ID6QP8lVmWCeHljQOnj0nvLIRolQdVkl/eEcWlys93dYa75/ZOlTn+1rzoEWFmZMI+F
0+ZyOeFEf0NfP5PN0IQdNubnfzXbm9HS5zFwo6jrjVF8lPEfPVdHEeKeHeyeXiRvMzDBUor7Stl2
xd/WEnhV/BDvJhV0QI8fSINCo4dQRHqsIQBElZCF2AUp424HRCMVnrYBvhop53Pq0yCallpFsMbE
Y+vNvyFn3Ed4ViL5uOSlBA3XA+LXcsYePqNmJuAYsqsn4mC1mjDUJ+bW/4q0kzs6ebsRMZ4/mgr1
OEFdvxJurYIGayOkHYWyktjhp0DEclIsfy3Sh3E8VrHJ07NGxVWPDTfQNyKfG8jX+JI6g2JFRuFV
cFcKiE7L6QC0gNy6A65X1OD4AHsIawWvyeDU9l0nIXvJ5WmiDIN0sVjOwOJBiJwCR2PFQ/ZquJE7
c//sw9jyJjSh3cDK+JGS20vZC2qak7TUq7veoRB4vooBiicEiwXQKLVOlY91FP2IByUDHk9YNTWk
FsgOV6NH4Lc0a/uZMQX/ZafQ2KjS6dqswPQ8sbXojha/9YdexwXYt70jQ1/7W178+RaIrVLvUj6O
l3m1AgIBX2mtA2iye0ESbB+k1wU3cHto8Qw7nHUONeQGbM+RQxv7Ifn5ZgtHHMoOwEdQw9doD3Nm
rgjnzf8f1CqydBS+rcxHALGuPKaNWW4o86u50WbOTheTvBgy2raVVkaFRs7qmL79ve/LPRgrrnag
JBcbxmS3yvbZ0MRtphVLGZCgQ/ajij72h9vLWSncr87ZdemlKRMshpH1IndxWJ8VCyfYGQutr+Y0
T5vd4bCuDev/Jy0oXdq/ps9G8RwcWUK//3Q59qswbEe8/g5tBYZQCEYxy/BgF456uQg8u02ivT6u
Vj78+v4mcQJVQBq1fDoQz+BFz/sqZFoXPtdvhPOi7VWqSBkY/oA8fpXWa8fW+uQv0+l9W4HTk6OW
gJKw1wtPYUdkDo76hxfaas6cLcAb3lms1xQr3RiiiZvFmTlrtxYKS0UpFoQ4ancNaE/ZVrFqjPqW
tMPBoEqZYqK7ynYWaeq6BdmnnnHXDEvXW/20szmFph+jw7rQv8iJi9hDzjLW0WB4vkSSghfCvKdi
G/UPRXnH5iF5BMIctTGVJHYCqgZ2GlzfWetwb1LC4gDKuLAkQYxBlpRH6NpI6fL1p28F0zhfeL1q
BFYMfTXqaDlnvMpwqAzWbrYN+5dSqOz5Mb4SkEztMV2DuBchWfTB7U4Wbi3QJjbHSBXJczGqYyiu
Sm8sSkmI+zR7W84YnFx2DzNbcVgINwRn0UV1hbZGXSAbYDfInt64Zvl5bXkJqCQ8zLB2HlCMm/ke
IIkdOlUbEdTutTElLuSGqeUxvbUlXh8m1paS2reo05Cld8fbv4aErT9p6BwENBD6wp5aAxCj4pvL
jWgt9sPXfc6708BmQMljccAmQjKtwmbK93E/RlyZnwb3O8le2RLjx05HAQL0Q5XY6h/KEHRBvTYl
KHPJ0wvsaxzLSk9M01wtyWskHsWbQGacidIAr74I7peWx3F4SAUu/LhLz7kJIbEHmuYj5wdT55jD
/aPPvR3vo/YOL3Q/fqH/YqMAUl8rRULClbe6Ohrgcetl0cBLzmsstLeX8WYcYghQAvwUNGs5FTFh
aP/qqiZTxXFPWjGppYFDAj2L5dK/CD/UIOVNaxNSXHFvdfQtQgUzytJGG1RFaaJr/6kfHM4uS93P
fCy1ozFGnDMLc7snIWcbM57c86yw/S/IvstGqHktaFeW/wDS/+MVIcCsS8PcNlYpMpvG11L1m5Gw
mF+Fp9hZLN9Cz0bfeKZ88cLXM/BO6fZoFUd/SUATh++gKecbrjmY96jRoxXnrZfXF+AmMFVHt3je
nZSes9bfGfO0s6OGNL/G5TF4OSBz2/m+MO4c6mclulTizbKFExdk8w5EolZiKtmLljqauGMjjrS1
HjU19R5nVsuiYYXbnUOoAEoMLiM/q97mii8uPZhE1JSxsEua4xrB1QHDX3izTUIKAJ+567vdALuU
b2Z+87QBTVb/SsKWGI5Zo8nqPXjCcIv4smhazKWIWDGElDUTUwXe9g57xwAvZpGiLZImLPgyopNc
dbGsRrI8YK58u8lqQPd0bmxaLfUHZdy051R8RRePzbtyTHvgAdsIxSi5JHybsjdGDIPsb1BZfefK
8LWZxRTqLTzUxmjWJ7JImdEore+CFYSYSKTOYMNy50Dk9Hsoo8kn00zDUo170+QkmEmY4EKFK0Ru
xlnQKBSHMUwFCZwNhqdg0AfZ0Qs6cqq+5BbVpthRFDyOH+xY4uZLPcugBwUJGQPLP3B2Xa/JwNVw
BpOCpj/3I6W5lUpraquitPrdqi7ASK5CD7pW2+ttvGC8qnrT93O40AVfTU2Tf4NG66U6yVwGO8Wg
/7+nNCC63pmmNhTfmDbZYIxEdCg2ygtBXB27O3vCLog9SWLExz8M6GCK3PT1GEVhF6fZ+Z77u5Rc
siLPyYiJeSZ6uPHcd+lRnkqyyqbAaA7WA+OsCH1iSfOvIGk+KGr0dxg11Qkt1TGueOV4wIju6YeG
aQJ8XM3fJv/OzV9ZAMJtxc9FqdUEbVRQaizBSZS23FaDejwiRWoZ9MiwL3wqDV6JxDphVs1Gp/3b
UXQ1HdJ9TqIxvOxHmTk54YYK+LVwaprr33QpviAa0KHJ9pLR5zPUd5iF1PEziSkPkEg9k5bagowL
K6DjYfMyZfeb3vT1iR6IaoZWif6NXdw0xSg3IfKw43L5tzm4Nmk5zoLhY8TfwH7Rt2zQPB4KfBC9
vZrIhddLpPw8vllFokR2mDl5sMMvr3ySMoQczFFnZsCo2hom9msX8BdoOcgBPgS1ou3b8ag5qLbW
TIQUQo9PIk9VDH2NpuUxmNKHuJOcyXAgqmytdtWgfB6ov//b5ntBvkU8nw1PFzIC+oP54VfNQttG
3geif/ndLOU+QfH1nSWWvGQvAUwA/C0+wyc9vSs4T2D/YRzWZh5T4O0kpgDxu0FhtqzRXRSoGLtz
wCCjHcOhYQTKsspRPMrAA95eMpgZsKy7+LiblXkm91IGrqcfg1O6e8WNc7skr0auVofKzleQLgHD
bQgggW7xpwTPGlcuPkjWrISnj3QtoHRKXqQrUeNdwiG0SfyPEMzPnQ81XVt5uQBy11ajV+c522L1
BDMg4O5jmhiL32JpKRM7UqIGCHDKv4zjqbPbXpHb1Q5BvK1CIvugTbppu3NKPhPoQWPQ+qFEvpPo
rWoo9TUzBgxjnIAZbgHt1pM324OIP/ioWHOVRwDpqMwFxlUIUxJnzGeHDA9K9crYW1NLUBcNdQnD
yN/SqxuFOBpe7dvMwSgdqjd2Y/boia8+gInkknPX9azm2NkYJp0YZZXtMcfIRgdB9XqSg+erF8Cc
LCQtEZaN3ABJiX0JvbhQcX7JcQdXFxas78Gv/Jkca2iz83VbpjddR4+gHSW+02Q4+DW/E/R1mhHi
eQMoJB+AuCwiKKxhWqHIsHEdu8QhQV/OpYiA7Wp6LAe+GCdliASCk2lCoNP0BlccAOz/hC/zK5C1
wlSyi/qXC9BEcYEVTRZi4YYytrpyUQmXt84/eXdh+2iv2KLU19+Wda4TWVuWuMhyWRcfvu6XMyVv
b8qzukRvvbIir9OPFgWyHCiGkDbBXt6g+s+hmD/84sFT5olbiptDYkEKDzvwL9AOnKe3b46ct8ah
YsRx0CEz0UuaKkVASG26KvE2WNUKcsMlF/0kXzmR3RyVUBRacwtVJK6XM2FLBL7TXRrj8RnPs8HT
WJCue96BSxCJNaPIzqMulmto4vFBW3ffoBuX+bgB4eK/lW6BgdOXsaSaQAJEfF3n5rfECMy7Fhmz
eamLvp1Rp7uUwZ7XpcMZL0W2X5BrPloku2XJqfX05rnabuW+PZjQvOCITaZ6JSGQyifLHLQHyJXG
Op3GnOcr7+9cJPn10FfJVtwXrvi8vO2q8LDZC/cFGvWnJqmyaOmsuky4b2wGHdtnox40G2TOmMTQ
N5px3i15dhr++mIArjlKAIQeS0Y5UIOa2RU7jguW1VR5cMaeTefgXuKwZi2m0sEZ7IqIrbc1mCTd
FfrgyodHL1b9Tg9KkZCUnTSPxtsP6EFoCZ7y/hdcQUsk1TZTjZRFG4NjEQkpjCvvX3cb9cuaXDuC
fE/8IGkbji4Aud1lmUdny6EcIpTyiMebK5gEn/RF6lOgHQbEttJnOmzx4SHY7mkST+zQjc3x9Rzl
jb8v14lrlT30zBP5Y6lfgcOiyfPcEurqaJeT6t4ezrVjxMAzGu7TU8Nbsv+cqXpN9lohUXac8/uH
9OqpBymfMK+A1vWS10ZePKXdxXehUHIBEbrpP7LKrUOfQhC5GUqTVvXxV9CBZBCCtMIWt1R2Ar8p
7of21cf5I+a8lcMTYh2HOZCt+CwWFGdMI3+ZTkSq1viZeqwJuj28WU86la91q18hopoF0Ag2yN69
cI380hs1ET6KAad/mBQvqYOasdO8L9Kz51iyPOBjponiTgNw6830saUcz93Q1HT4W70dRFBuTm87
vFGe+HiYLASqZITVZUFjiqZ1R6Ew5+7wxqzJdxwxs+EIQgvOtzF7/RWgGBubk8x28ZXkPwPSd08E
zZd9qf+xLQmoTB/yLE9mJtDZwprsSIVYXhE0M2n0ZkeQsIGmkiO+Udwx/oP4yxkGIf9jgcILMR9I
SVhfXh8kj+bdPrdnHWxCcHcMq6v6jD27n8wuwPn4vsXr3+62aoKwaZpKN+VGVwqs1YBOkW6FQhq0
EfbCwqCUSKwHuAWbVVJZ7TTNw+9HqmLhi/M4I/WpVrTQmGRAHIQE2PHFDCLdRqKVZCLFcHCz4LaK
l+ThlUGSTepm5VGYCkldU3DSuSi1JLmME4H6X6ymr1snaONqLJw87xCFWM+UHwuM2v80aGuyxNJS
CnKuGt+GetgfURJ8htO5clgag4QeCZT4hBcUaR2H35hMRG0GyWwxKO1RBnNusATQfmQgLWiWZmiD
aT9E5GH6xPmX7ObKD6W8rQMFIGzMQCa5nfXsoXnrox6a+n7usk+Ytrajdg3iIv3bAZfWAzv+cUxy
hPIOBC6CYDxM4Xk8SGqvs8iQmoC6W182mlvzzgN5/G5pdKIhM96FjliphgheyisuTrC9TQJwXuan
WrZxdXq1M0SyAR9h1hQirffRU6OEj47gS6Xl2aeUlT64+gwTGPo2vYmgX5wfU+kWD0+ByCfLXd+A
skVtJ4+1/+q3zawDKs6JDMVA3EzBgbvwk+ZJQJ/YYyvEM/KeEvL62KOu25+9l9KnfeRaz0+AZsdW
yvkDxDBo+LIX+mOteGF6JJcGEOtmJkOyiTyqQVfSbTLOUdLkPf+E7xS+3k+vxj0/2VU+2yEypDDo
jtuPeWz2IzI6mX+fyL8Kxiiq9g5f8eF2QJ93SYvIb2RAFsJCqYS4m3AL9iZG5XamwdUIoXsGdZ5q
GgwvwN0hDojOJwOsYtJguukRop9djKfNSttcOA/Jvf6c6hmtL9/vGcKNRSXDlr7+cvlOvN1E+TdM
h+HSGXWDuX2WYU4b+KEmvnFa45lAdboh+BFwj2cMWkIQuvd1etxuFpiSK6UU1xrYM/jxYLiyY1kE
E8epdicMeGZ0wQPzxBDgisxdsrCSpOZPnxMZrUZ/+OJpACdA9nzy4AN3UFoSmIisdiER1XxZPqzz
qw2tecKweKK0/ZgxV0fiMOYoimjYUiBUOcJclNymjUDd/YgfEFgNhoE1pzYIRlzcvC8EYC6oWkb3
4IZN0zMuqKgKH/3vHkcJ/PjcPae4AQYIvhaj+CG7G5z5R2XjnD0ZFMfrCc44DHBYLwIkq6FBBGJk
BJ8UMvpquPV+VmJaoX3evYtkHvySe5HwgppoNGG7x7bSsUPNIqRM5PJlxznUM3IBRTYJAFPHJIf4
hSMbBgT6Gb+45I8LPcTQOwHziFXEILoIL+cdNfchVaFS6Y7QipyQifSk/+w02jZlyx8HD/g2bu06
WdhzxJme3ohFOP4geNnGnnNcafFlaab4J0fnywo2X5eQssTNKspKvIRRLj+0TZIRux3+Jq0WAvgA
4kklG555RVaH7NPQsuk5q2XQW+VC0hh2fbWC7KUsQkysRzBMFVnuPOUHBmbZONo/f5gK2fJtw8Dh
gypP8bqlhenJTBL/zq6qgMc2IFadka6pvBC4mx2IY09CQBUKrCatg1K/1tKhpdXIGELu1UCLP+aS
gnRLYyF8Ml/rdZNzv+gwqR2A1dw21VzXUgazVHRcN76hcx3Bzrm8Rd9aIiad6kBoRe6QDzTaPimy
q/ZorjjA5SkrIayQyqqoCW2lx5Fr4CZ4OIOqyOLVKWLkndYdgvkWaPWgJj3S3gZvTlIS3w+mnH3F
8EHi/eYH3UcEV5H+DQutKR+WTfklBi1gJSLJ/cN0u04BQYE5nZwsHAD8WsQne9L5goauBsJhim5M
FjdnWUdgVa0/2q0k5EXHUIef7FNyBpmVEiIVYRB8hWQkkvq/7xAw0pu8QR6A0xGnl3vPyRzudnWC
9KlLPpZ/qFrVilktgNIVi3Pb/l07C8vfORURKa11NJkAR5u+fkKNYCCbWOjQYdotW1uR4CxnYs8K
Ty7NzAK+Pf6ZHBHiRWLYWarh1R8edWNjyGgQnWy/OdsiipoaDJQqixLxZX7RctuOpyWWmj9AE519
nUS63MBcWRuV1vJIolk3NIZOnxn9ChTWdmEZO/X1Ucr/WyuWvnNmnCQKAhKMl8NVkLZMtXxTO+G4
hJbB7nn/4jmlRZHWJ64QjV3nkZQ/q3YTiUphAeKSUIzdRyx7JyMOPtwN/7rtVeBjrEZA/vhi/bN9
ocu6wy5AGStHsQFt2h13/T7MiaJMQ34nmMZLd2MZjM6esx7KLoHYHlimQmi4Cofl8jPfvqk5zcsy
Fhw/e17v6w/JU/64kd/fNLkeYmNcPmQLXiNXGtuxY6yJbZy5fkMouKqCR8ApsfqJgq1xov9KOl23
nqGQOdiTpQgp1yVyCzIgl694Mw72KCT5n2nEkxFv9kCrqM2qovohRv6L+OAZptVHNGfe7Tx/Xuxy
qeKRgnSySELDkIWlMyAAaRzC56GapdCWlY80+jevGmvgfEtNgVvD/Oh4rD8sF/1+PV8Ol++PBwmo
orLehwDrfL2lZSJfUdeqdeO01MH2d7BT/1XfhPbxhfKAXJNxGD61I9zbtDBzTMmASSo3znozMVsf
6Vi7GEJtrTdrrtRnCja3ruHbKfnK4Ch/TPDa4PNSyl/YzLriKnUbMHlAhktnMRvgT+EoaBvVVa95
Tv/sb6qhqob8g1XNEax+tXl7u5BLuTl9npzMchjzFJq+gci9PlWTDy6VnTSBsRAmKAVkS6r5Eswx
7h2bn52CkyFC2mmKVkbqKcrwWKmWg0CTjSpfafd2xUsBsigMhE4WdGPt7KfhoyAIPG837+8oQ912
Nv73qR90kEXLZCzNrRzi1MufOdfnqegNx2f7wqoK8VBCBU1hZHakKc+H4GxXoVBbbof+N8lQ2nZu
2umQL7x2g6e71rbDNGGKkd2P47q4BnpAGfK98sA2xBobD0REIqN6azBCQhO/wd2cgx+s7mW6cPFK
Jq46qLHt0UVaf/GJZb7UfbqGmf/UTDGDWDdqyaNyGWyzTi1zMyN5JzG6zzJQIhpYUZQiPkR3uRb9
VutrfVP+qRhOr37CGBXy8DJSqdJC7GC79v2ne4yqGFvvEOsEuIY09xgUAXi3s/2DRKk3AhsodjM+
plYx5CsoJeD3yTbhud+VAEi+4yg9FJxhdKRH1+2rjlVGN2VVNjmXnPvul6G4VrBcULmrgJViUGXQ
tBp8ZKEO3fF/1mHCgsbPXXeyHkS/WSw2Bb5E8uup3OxwoRwPBr9UOShZ8X5raC6ORKFMg/QztCnP
war7CveBdcCvSFKfj0d891NErBXgZ91WL22RHXv8if4cSRAaF2grY1D4oF7ReuFOZBvyXB6u3/2h
LpnBZMLDlkbeXgSZ00c1RwBLJuAfaKkuvs2SjEpUWcSA3+OhZ8al33GbI7cuJB0eZnM2mw/VAycj
WPmZCtMIxTvVBiB8iPhkE7NjxbFLa6JO6Qc4fIp/7wgfvqn/AmeW0jTigRgIVgjtzkW6B2AFWvNQ
eWvnlLg+a78j8ngPYxp8yfHGC+3LzqY6v4HgIb1RT19vvZwylyOJR3gS5VpVvH4WA8PaWP6eJ69a
K+lZwrohuSVFXLNxPwgjy8CQGIPXVHTuMe24v3T+jFGDQ3qwooM8dZzMcSxCB8vVm73CfvVcAAK8
/R09+w8u148/lKCdknKrOV8z8oba2XodieucpA+EIqCBSVdhWuZfZcAMQpgegiYrYZS33qBY+rSh
fCzIS6tGK9LvS2oRScYd6BWv5O9JGlE8USKcFnkwndtySud8jSe32Vk9NZMcXqePLTPpA28r00Fh
ZzvLt7idPxA6bggcz7FAvh+d4B4oOk59vXMUtds5XWE6y45MIfHr3nFHBoZ7AJWk+rjKQ8ruwpDS
iER1qSwYsi6BcQbi3st4iSez6DNETG+90rx0iTKriacjOL7pgJGxwfbgVq0fX6gg6oqe2lPuZOYg
rlb7gSKJRcSRiEWtuTvmDIrLebt6OHydZXUtxId6Pik0QbHcF1S2fRTiSvVD4paDhvKHlGQlFNHo
DI7rUZs8eZ5umInXufgIgRtimnm/OuLYOBOkxqZmCO5r2oCwJHqPqkWEsDjYq/NFFx9OkIcvaGtS
YEdKxvHuy3jI8/tnm8xUkfCDKu+WFSa1u361IJFYtTld2wgEskUFo+1+OgfjyEWWrHShdTOtPDRW
23NVU6luF6Q4W2hW07bJRWJeiQhtJ5kbZUu/XqYwDPmQRHc2nq2xZu1kkhLFtXzbBkbGtMJoFPeh
cy50k7v+Ys2IVZnizCL9kRkvFv2kJNJ/023Ms97C97+zp53P1RJhRoyR6lS6/JT9O2K+6aGK0Cpt
dR88iWKy+tlgqnaG1Q8K0sZ3RJaa+jsvnWQGrSqmroXwnmvWJmYqu4cDvbyGb2YdXUfkSNQF5HXf
dDq2sG7AeM+6q94C2k8g/U45JUSq9BDoUDk5ifk2+4a60bvNR+IzqHGFwvSIHPM2i5bHuIAynHBS
Bgxbh/GwCj/Ku1lO4Lbvre6efX7dsdqYMpYbIa7yRhKaKPmLCB6W20Gx/0QkEG/Kdq0HBnC0D12j
18YzDnq/5g4ESM95lYQouDIKi87utUBC3wFFulreuyG6OiDuqpuV90f2CL69u+Ezo8AmmovBLYdZ
SajJsI/XMQXMwLfkEm+qz398wXLOIAX9DtvAzik4WAHYkJ7zc4Uvl9ZfoU4DYBfnU4tZfLuGQ/QC
X6xr/hDeHiU2pYRdGW7jjHvFM8AZIzyoNJDqnyfbgqO9t0G6q6x0zwxj83QU1NGmxnDLdbS+X7Mj
fWVF0TpH+pIkl9LfOa3lmSWEIgkwzBRKDazFiRX61/QxI/9/ngjqFer/UyMbp5U86n9B+Nm/LBKO
93iDkZXz8l0sTg1a3NOB/fF+vuvo8B/nCs5RXUjOaN5poUn3gyK6QdU8EHNaAvqo9l3Su2JY3MAe
Kgp8RSVaI4oYzRhX6EExvajI5XSscBnONrxW7ORGaaRQMBOdk26XyWa7r1uPhuNtifBSOgaen4up
9k446iUDnr1Qx9dGmgJoW1hjd/ozilJbbmX8l6cevF7uQL4aW7jFj3UGVqvpPPatliH+SFVdh0dB
dd6M6F2/xDWL2KU0HqMG3ldgws1/w8RmHTTQEMWjaQ9Jt5zYDY7iRf+VkHnpAva7E4s5281TPqt0
8WW4FbIouJ2MD6nYCnbnVpwVJe9sNpkUnyrjlb0STcsLXS/hN8V6SjwvmPXZMvmetguxGaDzhs5J
Pg7+Nwn9yY8LdoLKUGg6AHCVgxioB6bidpw0Y8bqTdDyblNY/tbrDE6vnv1pbDac/gXCpqpFCai0
lFnkhzO3AOR0ZhyiFwztBQyTO/MFlIADJVeahKyfzSJ408bdiC0wSXY3BZhbLG0UDBV0qFBHnD59
Etsa6/idZ5M7/LV+8y1gNiU+L+/SIquRk0tBlCVlWtYzLREOS6ehDF/srxu4m3Sr/ApvTKbZvf/2
2spYAQkF1KAOEUE1sH2ycLrpDQoqzzX9keNbBCuUFMT/tFoFixnzVANHtY3O73GQvo7AolYBsm1o
ADg5psnTeTSp3Y/g05XbxxGscgQmezA35RQlmH9KrmvhiA/8VMh4iDec4Vzuk8uO16PjUCagZSSv
DpfMb8peiZUAl4b48+xFPsRkipZH6NQfvUL4DK7+54ZJKicgeOPhykcyt1n1Z1Q52y//Jkqdu9Dx
FhpG9aQQ6FnhD+2xbFPekn3rmY0TqT12JyqgeB0W4mOxQ97ARc1+1z+nx3nM2UkjAkHN3WSTb4D5
uJHDFlv5pkuus63GjVEs8UFirErQGJ2lnm81hGyeLc5RzU/Grqoxb0HtQhYNG1JIQ73I13beR5cs
4/hX3rOZU1OOq2Lefw8XebZri5V+tfZbxzGCzFrwdx82eOt8+K5OjUTpa0+XIJ+MPu1tdq9cMPq+
sUx5+0D64g0CGsJjzE9RLJeieWwjxD03AcfO/8ddmA3+9RRY9Z49FiBGgH+NZxTr/RNiJeGE1n1y
yu5Pfk52p3rIO461TvtgB34IQ2j14cttlQ/YgYEb/CRbmBQ4SeR49H5YFA0++qYSrubi36DQWONy
jOiE5VQk/vbvMTlj7MZcB9zvztVUG/kzAw2+KG1c+sAHeJYcJXHqeTYQ2fwhjQZI0h/lAYK2A/p/
j0dJS5LLrhtlOdCMC2XUkgvi/67e88Rc6ipOzHb4RE0+0S2MLKg5NfrOCyOQHOpZGYT2JF+UeSIh
0lwHRlpab0kcpFG2bkKIWr7ueZihNhpGmfafhipvTKdIrV0oOwykuhhf5bz005Svt3zWLcsBJSpA
/RvEQYdfXKDZ+ndMWBZ9d4pa2YTTZHVEdvBS70lI7+EtwyGGEKb3KDztEOJKrJasDMkRJe81PSh+
w37e99HzaCRSftiHm1OeorzdnSqcpiCoKFkyMmyhyELafMIwq4A1I7f4vZwmkSNFWm1akkcbwZbq
i4719nwHUlfH8YfwlRO3VDMYcvFO5SQ0zA+NY6QLJ2g9DwJkrvDCIMdjls7+Vpxkb0llUJUMXMCX
8wpX9t1wNsY+tmkIGXSxIpNHrZJeqlBRT4+l/7PlIsGegH290tVjEoWOL5YR4m58/9WvuPg2ypG8
Jg6P+0i5/G68WWgas1gSMyCbOleOVFCX3h7fhw6jt3Kylo9wP5KjNtWR+jFm7hu+oGXOeZknBtw+
gevD4Dn57W80NZfNbMAhjMsW6kPHedIbwtIT3TgY94tRQjsKEEr3MozpN2qUGQl80DZMNe78+Ny9
A/CYP+HgFB51ztw//ikA7ttPufKinTuBOrnqw2c5E5SK4e7D0+Gw8K6kOzqmcAkrYVFKe6jrZCpr
oN+YWg2sSiDKvnncr7sobQ298bsVo2xZ/XS3zLcu/J6Oe3WU8BQZMvGZTqNw2iejrSTxQTWIoh1D
sQzhsBAN0g8zUEpyzc0hpc3lzT4Fc8P4YsRqdAJuVZzymqbBGibS/NRu/MrZ7g50QAzcdhZxF552
r9LPDY9AQyevhloTFFtrPnLbYo7hDpbYhMPexrq9cDYqDxW4pA6F/735TRb33xFVo08eEl+MJSbA
lYgxAcBGUaOAC97WD7c8fJQE4CMp+SM4JWkSaHmbnXJD0YMl8i7Nu7XOFtj22RXO4yExneWSF11t
B44D91zaSEp4oAWiBMEKs2jLw4usCFhOpzAoatOEx0NN0qoB1n5q/iQlrjOXFzG7SDmbGvJnsfWI
3mrLLQ85qaaU/GosZ8YKrXtVnnK4QFGuwQQlG1/1G4ZLTYN/rWUneD3kRJnePJS7HzlCq3xiABaA
jUJ/M5US33LpliY8BP+M6SdYJSPuP8zvsvZ1/wge2W4LvWmwzuWQPKNbsJ8so1RYXbp0K8uMB52w
/y0orvh1j4DVB7O9FroxUw7JjczIl6NLrbdc2Oz9bxbnSsQ9moCSGzHcCRUn4wg8STIbhEdGfcg3
G4sVCDNvWZ1mdBOAiIeLcxYePxNH6q9lsSTV4DDmI7ravnQBqH3z26wtfqiN6sYGKIYDcM1WguXC
nInbylKFzAuvd82GlzbZvx8J9QVngmVwb6ZtE4NypfRBpHX2THHgtcr/juJOTZb0Upm+eT1VEDr+
aaU+WVY+iI0F8MjAOD2JTnvFNFbY3qfcF9CJZJmRRJSLPzyRc2QWaV5UAf80nFRGgde7XCTSe155
j94Nf5641J3Bn/fZIUq8AcYdIU8THqNIFAGp2/hnew0mPJlfTarOANFmJYIo/EYuyO2XJQSZzXgF
3PEHA7vxV2m8UYRqeQLH1CfjxRBgVEafXMBW+rcNKr3lhfBiJoPF8QQ6Sm+ZE5A6OJF5SIEy1PVS
Zfbbf7PduJxSHV4LASJpdG9IGvimVJWxKB6qUgudT4nBzEi4wDknHnTwIKekvvzudyHa+Bx5Jlya
arqloHiTxg6AWPZ7dLYscouKiwsr7kmoZDfITkD9HKQfRo62Om+ema7fK4qBlpqxqxgDRxpIAaMW
aFjpsJIfjnWKAuXdcr/+MYh+SHItTpLivIR02BMlQFtsuocbFmdc8tOnG7XN1Dy2rsSP6yDGscqQ
Dsgvw6La5nxxHGVhGaEckB87QoyS9f/CXw06HdcWOpADzkNsyq2pqNyuHy3pjHxDJ4KeaAR9d96U
8JEluiqgIJiem5A4Vll2jGaFhV/oGHUvMenjeAJiqPGvird1/PxX5QwffcfEZ/ANwBww4lb3a9CS
vnKYblFq4fdjEknwXPQ+Z+lOozFrc1YvUC5srH5LiBh5Y+cVYecPoxlgtdO9KpwNpXAudDnWRIXN
ezW9Ug7eryvEx+p5SI5O2yGcRxUGeZw8yjAPqvWy5lRYDOuRfDw35sPnFeO2qfuK/qtHsQplySeZ
YkJIE7uPi1PKHg8Cikl1rwq9CC6YNMeW9+bAYzzxaBKQOxiNwMZ/ZfYq3oI7YaIiCrwZxICaJuPa
ldImv2C+LcfT2VTq256XNFkJqteeqtD756FKSGZOB351TBuCfJtKCOReBdh2ZTa6YxYKPUa2axsj
Ysow6P8t+nJeOuq7Mvvt80pCGk9ft3mMa1mNNw605or68Ih6Cvis3oT674zupsBECub2LSr/K021
4SjpaLxAt6XEMWQsHgZr2Yp4WNZG6X/ZmC/M+b1wa3gZsVZMTiSXEX+WUiOanXWiLpXXNIq0KZFB
IYxhtIDX60bWcXSqUhMxYCZKbl5rujSnAwX91cy8p3z7Uv/Zu3oc2Wu/+GPSOusnsI3WpdWojBVX
ZialOpbJfVKY1uZekUhg7Jo3C0CwJi2VdKEKIn2GBx0WdXpMuZOsoQWqBrsZUtqu9CeC5BjNNqOo
5CWYV82Y4U2GJD7FF6A7fXSW8VPZGtNrx3huKCCfsy0QpbkxuRs/GvQPZwHAyuL1BZIkHVY5FdmB
cW8qWhewcDA/4xKh2sILjwhp5mjabFTqnUKwH30tFOb3v80olVILz62vL0fCbPDYtghTrXYuLMnv
iROa/w/HQazPYl7wPHuDMjxoUenhXhPPvhga1Nye6VJEOKkl84SctSqvyfVRB/lIUz82IFQakpN3
xs7l+3WCRnQjxu0r1HTRdhqgAeH+OnbhfYfPAo/QWekHFB3S1M8p3p55JgSVCgd5Gvk6AZ7J0Ehe
XS3MMKJIKrynRPvRn9INoGQKiGWsC4PHM0fnFe+YQg4XcETlEJREJcem6aoKhMFwKP2iM5J0LqbQ
4qv/XvjoPV2Q0lKDgpa/AbGeKa0m5tQYMSWx47bB99ZoP5zN86kQfxX/zwFsjlM6JD/CKiFBzv0V
PgmK2PttNehTVdTEACy15ozmW1NvRIggRqCKcbgZ4M8M4wblWnlS5iHeDJIl4bCIXIdz+VqhWya9
YCLYWXVVY3dR60OjEfg8uhyNKE7rc2Vv2z0HRLciW2eyxjU8egQ4lkiZuBRTOPgJjt5LjQcXOpbx
E41COPBgZOhmhMe3aJ/Bg/v27HBZrKaNk+quaEA8CkyP/iukhTLEqPZvQb2Js1q7nb/OwAGdKypH
EU9vfKqfVc8okgmp9X9ihkUQwvJr/KuDUP/+bQ1E5TWggiACcq5kdIfYZq3zCqFdLTN7FfhoN2Fv
njT7KbcT8YiK9NhO4B1O9UKK/X7eReGM0oiawbwBmVBUrw2ia26HnAVxAudgKeZ59+UvUz+aAP6k
xuxEnQT1GZXYwZgxr5o5dnrFIsd0r7l0iLA99Oh2ORPEKo66dpbvqElrhqHFIlsj9rTDelacLBjX
NzP396+Trq11D8QmvPMfgUy1Rt+BOtXHKJG9iJkoJkI6K25nBkW3U7VNJJt+FYGxhBC6J/mvp0gO
g4tpI8HoVMyA0s8XSJKXOsGDgTEqHUh6fpSLxHyJIMZ0RUzTkri/mwG7FSdViBf02U3HimNujGW6
J2fWp0w+YMyc90c/kj6uPJxSSNK8I6niq5eZnKbenV4fulRvleV2UlL/7YpUMNznBzOO9lkIocQ2
gb7xZvdhzhQImqx8otbLnD9IVzFRlTlkIS8jtYk0Pcl6WfyQOqvs6Aa8tEZb1jOIJybHtG7auOlJ
2gBfcF2JD/jlv8L8QzjrEfeaggNPCtUPaBLuB3bcv/g8SFn0xRxxI1uDY2v5GIPKKUfU8WORZZcC
LTl4bDeQJRirGwcW3GwIgT9OvrjI8qt34jsGTJKzAcZYv/hmx3A3nBEZksOzccxOllFyMwpd6Yg6
V/CwXNCj5zYRWyHQOG5qVHP6v0I2dm02klD1ifF5D4MZZKJa7nNmMUJvaL3qvrPr2bVnpDJS91ID
dUXYyJl1MHtq12/wFOaYjo02OPKlO7ZQfxL5j12Z1/kOsS3J0+k9MC1kezwZaVAoToy3499aSH2p
7N8fqp4/GW95Wd6TqG+tNeLVRTQANE63GBj7lmjeMpy/QWrJsL8xQ2SQwSsku61qZ7TRHcWJnEOq
NDrCO9/DD5TGVpdyxsZHD+U+uoh3DiqnUa4LQn0DRExaXid6GZXRVCzMlEsULLQhNwOz5szmt5xY
c03JT+Jc5F9EoRWTjFNw/pJX3BWKsW9+kS1cxG7GlX/Yfl91ga1tNCVnEg+kNovFg2nTT0g4p3I/
igWdviTOE+Ct4aaeBdOmFU6lmli39CQxQguAq0TLMGw9oCmmQqyTkP85Chfr7+ENGP7dX+sPB4T2
xLcne3ZMUIF/YSZcply2Im0XqLvbuEz/QEAsYrhZ3D3hC571xNwP937BjASh2kxs4j2+wTLj45Wx
6nYzUmr29Y4fIr90nvFztBooZhUlrVB9nxhagXGOOfGbz+huKfQm4CLJImzPKU3mzR6C73tgHbCB
z1YTW5Z/xDo5ZW/h9rIAyBXTIXFwJfiKfYPCcs2uRodM3VA2YxjYtvFJnn8q/rj+O1fkpMK8qd1F
EedAwjujnp6+OFn5BQei/fhruIqChcKEI+8UN4AEwBZGqHs3rE3YGQ6SNbC5aS+GoT4ukuvk7UNx
0f9vs1ADqP3kE60tFmXstjyOUIKA3BPcxRlR5e/hYDLFQ5ZJG2Xx4fc8uUpZQ09Jw+Nqk/V+2FX0
Cm4W19hvDdRpXWQWAyF//2ZNeZdq3n4PFVgFNQfJVXR6WpJ30lHP/XyKrHM9iJNxZcvRIzKcTERA
xt2FKYiKX36O8r2742hk1E7UP2tSP29uAbKQti6VY4EyeagNN+G7aCs5K9+wMEU/lvcwmdyq28FX
ZsKfz07VrJmh1HbGOOs/CfJN+au0dOYJEH76NxbkZ+lStDicAdfYEw2nXRMZiJQkl/3uBCmnOjC9
Ek1zGnIO4fvg+YBGKopkwF2l38qaU7b7pdAg0c40Bb8Cc2H7mOzRpeLucUAUaErFSLRw3Zq3iwyz
G8TEWqyY33tj13XlVlra2KU6HLg7wyKM7tKP92ZnsB6xKRi1x7U20qzGjGnaJs6s1TZilvJkH8Mp
LCij6ojvDWkg/5C5hVzBY9KKsPl80+w64OVxdY33E8uUQ3dbcElzoDGpKhQxfY33iU6yWEjECIuF
B4nXy496hEe69sS/fP0+fii1AvzPcyMjZ65CBQ3l0k5gETUIW+9zWYCOTKoVdVcmRGNFCtKld3EI
kftBwfthO/Oy+6lUJctOboQRYJclGXeEkDccsWER3YwWzQtyZ/fO/R0h7cRobABHQGeRcJN8K7nY
YqE+lV8JgGF406pQadZR6o+bxXpO9+QwZjLnxfTeChJ5cG14KJ7NPRNVc1q4acunJ5QjAyzc/EjR
M8b+L2MyBs1T9XXDi8uq9Ujv8n98hkHm85CtvYIVxemIrL95wtvGMuVyZxEsH+4UV0IhcPX9hJT3
caFJ+sLwD74PTJr5qPXRWAufdDZfAUHocjpgf9pWC18glkgHKsjrqZbvD+d/2NrS5nz7bx5DzIiK
E4i2PlTebTyZW/YQc6W7aEwf4mBrpqRdLlrP2wOPs9+Al7hKo5Kz9nTOei6YUYY4hP+Hmyv6+Ldm
+eu6+GFGti8HFiaCbvSFp4L20R3M6Uu9xRxlo3XLt1eulKgSVNs/8NrvvocQVHea38MouQqCmRzE
sVXaJ12ubnq/YLJP64XxuiCyj0na+PdJuPq2qn3JAis6b2nvyZuoRBuArLOIo1Rctw3gDy3TESf0
NtsIUnCdmy6UIFTrZDnElXj9FEUkivzD5CXw5RgcQSSqEaTap2snSReqmYyTuAIhdJHweMjOs0r0
yHqPshW6ohhTMo/ftufUdzn4c0KmhwuBE+pjPvMH4EBW7FK88bJY9RYmiUwyKdA7grDS8curzmum
7vfn79rEer3IkPC8zLnn34Y40mV8989mG1acW6JIvJjccgoXHCu30ty2U1o4P2mG3haiDqJaIsmR
AJCZ1Naag6f7XjHJK6BEaz1rTcsaDFYyACFYZK4M0usUcqvzaU6T5Bc+31LBxWIuVEh60rurSyA1
Lx5WthZ+YIVtmj1mvWcmsHOtdYQIZk5V+m0lQ/b5GN10r0gK+mVCaCblov/sbnR9VyTl8DrKat3w
18Qcf7dvABVgQt+ZZZKfubpa9WpUuoLK5XX5jbELr89PJVUfcWtmJIdJ0toUd5QfTwKt3bmWomFt
GyKOJu53ZGobbAYRVxinY72OfX+VEefdbftAJlZgJHHaijQ/y8ds0ZcOHNyaONVB0Lo6tdvVMw7q
hhqfM/8pCQmzvaqbwNK4QjZ+8N86s23CHwu2en9Sw4QBMRswIJgoyo3sWzB1qtvtnIEvi8IDQb8s
n0DgZ8OYQ/iyU6HnxaAeTx1+EZQ/o58I2YmV3npTXgNiHB2+pERjqnNSwtTXicQu1/laci362382
9bAWamwlYKQ551zME3YJDlP+PB+ATN2EBGOkf4bbeq1JdwDFf7wtEu3G5WqwVqm1Me+MRxmyE1PB
cBKRIlawSQXK1BFw4nuTNuyQUFpI5tvu0/2URp2NqpiJfmFA4pGjUU+8zwNQxzL2YJQgbv3XyaA6
r5VmmIAr086oNgNrbMs7nN83BQGB4UH1eaHCHTMu89z/UR1OgAC9lXLRtKso5dPZsZWjsmOylQX8
Gb3m0DTzOs/f4iI6FopV6DpGMVPN9uC880Tkx18PvXyc7GuP1scsio3HnUmpMZP/okf69mK7Tb3Q
rapWFM8RIID8QcXdTffzPDqOYXHMqEYQbRMCkqurYAondZm7d/E82UPHPYKlaoGgzmHBs0czxmer
BLDHlQQeNYu4ZkV84KPY5X7fOFfq7FyYjJ4JHK9on5EoaH3NPLK6GTYnvoc0cRRX0hRzH97S1vIp
GAqrZlz0mcxra5UPToRiLcnVFd6jYnFqpIvLWQIIhQbYEt1+9S8w7Aw+UDCSnBdst3xzp4q1MYoH
raEc0S2TTJXZgW/ofw9Z82T47Z9KTX1C8d0citBJ74xTQC7QDthTli9oeTn/tYS6WccezbPRV4KQ
/bDbUDZ/pFlG/V9rt7xganPz4668XioOR1UvEzfAFRhOUZwj/xePD1QJoHUydVRrSLa7Of3CLTDB
k2LtJBGUj5EQWU3bxxvtvCIJR74LxfupXwuDsSNotguhcuyn5hOKZ9T4jHBoBdT1VN85Br+zMrm6
escSK/UoEiEPVMMxwrofUcX3RUUPUoXvESxOIMwV9y+QxuTOVi9qT0XgcuiqaEMbjqSJCf71hQ/c
nL8WmeECaYh7WNDuj1wzK31bxmUv5N3bKOjpryWsxruG43mYasPsFXkT+sYyweiW1KQ0F4i4kFt3
5ZT3CmJ0vmbrmurtAm/1l2OxzZJ8necOijk4c2vKKZ7n41XTMOTvQwd25D6DJA3RE3rgVSt732lG
pOnYfV8D1HPcDj/W+kZOstQbAEErRA4x1ApBFMQrh7eqXHg02TwIKnMlCt5v7s6/LKDa0W3jfzqB
6WMU1QP65KSGbEOwfscXbB7oigvsA9Pj3adBSPf1oxiZHg9K7wNpu7+2jz0kYMX/yzBxHxQyhmnb
pM4IqbBIbJyT9GP7s52AhUokKxyeTovfOU1A5W1JUKlw5KjjtBoKExlEvKV7a85NAkBY8j+Q0vIo
Vast0DqSgHlkTYbp9i8OH+s9rjebTlC4oT7W3uGxRSOtJT2vLXOixgodvf07rSHj+92ZIHLa4EoZ
TLNg62gFYBvTushmhohXeMmlLzZrG9dP0p/tiNXYqOx7Kr4wz+Axx8F0sZTpSHo+saBPA2mDGQ1B
EjCGEfeZ03QVvlGafI+MzSBg68bor4HQWjOFtobsqAUqg/8E+WggnJ7im1o0csC20bZzpqVmST6J
55fM/DIgGPOiTtIOQbCcsAK3Rxm2JYbiHeaz6PEkC7cHIw2g9pbIp/jhbZ6C6AVKJKSY+9GlS9KF
As0go55seVwnbn8m7QFGFDoCIlrQAYtokLgfaJaJ8WtHeQZT/QmG7mVskl9szDc57LXFBMvBZ3QY
05oEeMUQgUTyg7rXpgHZx3IeCg6W6atSC6r5+nrKhPFfZPNXH1j0a9QkDtW/Whx5Bujtgx+tLeSr
YtTCRTflZLf0j3t3LqQfmbJml52MnzDOu5AyZXRkp1JalF+Hl2UeSaczWygEGEgetWtShKo3zMYI
pNcDKuJpFOU3PpExCG2d9WyZwg7Z4bGSQUgX7PhHUSm6lznpQOdnnKxUMyj0F/fwLieDomIX6pNu
eg9wv5iS6gEkETRpCSbh28w/X/GdrGkljBxkqC7w7qod3NcsmggE9SKQcEhpvLMrJ1wtwgZQ48M0
8DLZenqmJdYH2xnBKX2xN176i5EzO4bqapkY2nqEw19lawQU/GGuQE8wVjhCy+G+55IlQdgikkgk
mho+ftD+UDeord7/fOUY+PasAN9dRJUK25GwY/Z45gQl8AeFBCXZsXarjbEK41X+BZn2pzCt5ELT
TLrU/gkStk+tY8jgZ/KB5NlD9p/42z1qTGOwYFntYyUuA8evfb8NyXMckEi+fhJpZ+hB/8VY6vof
LiLE8/TOdY1zMyG8b4PpSC+tJwOwyMq1os+3lQtOveHR3NQyG+ZSSE5XVbYYvk1HHMa7DSEef4/i
5zLTDNKAzHX60Urh5zZ3HrSBGrbcSMg0AsQXIl0V7YEMt5dBvlnCq+JPDwZwvN4wq6ezFnpja3uw
dO93ifiF/tdITLTHqcvsKaKjUPUl/zRmmVJ+1VvosN1JPGwEab7R2g+CPVGo/hi8I8jF8ixdc+aH
AxtLIw+tW2M0+OOR02iDrIGD4q5sn95KO/VzpC7KT3ugS32AYVW8T+7Vqp3oiUJbeEGqmg0e0ehq
T960QbXr5r6iJt/UHWdotu4HPoVpDDZyPeWw+vg8R0Lfk8sun0u4O1Gaaw6yhU7ZeShBHVxY0vqs
ucx1OF5ZHWmlYqldOiH3nRmy7ufBdDYDrqhV06It1Rxztte4dvjqC12BndA0D8zIzOawFJXM7xcZ
GEDMejdLaC2+4AIks4muAufEsPZdDHm9vQK+8+O+rcpCArIZp4PbSVpjJcvV5BnfoLOh5lXLpOaF
XiBSPF7yfw9sdembPKfPaicB+CgB3NjwhRun2rm5IYBLkjMOPJG7K/XPfygSz6G5599asZY4qU2L
W8o+1YfxThE+DMrYtLspQ8FSlPT/RCE1TxUk0n9LbsWyZJpPwi2mrXRILVMyRHRo6vfphGns00Li
9jsrpuaeUT0G/weVqIkdLNdHmoCaZCkVqVBQTzJFgrrRlM9rpp9Z/5KzRFYDLLmqwfTKs85Bgi1d
cZaBNl+roBMGygKtVeEle5X8r53a8D0Bakd//hGIDA+7dbzvjxdIJisj7Pt3pRaA1YIVOBt6g75t
JVjef8ikd2b4+geKMEulS5QCYTpa0so0Ml1ieICgaCGZFXQvcCfmf8FUEfAXmWqVeKSksMw2yjLQ
DnHFbRJH5Uf1ZTAcQQhMjbENVaNtihA/neq0CiucDHei64UWZvU4nSQt4diApbm0IFvk3gXxnZzD
7qD4yFfYeYGdPzhcyOvuCx12F20fyc9qVvgu0Xgq0i7a8YcSrmdSvU6DPIJG76UKjaSdsHTFihun
BgtprxnPersGD+QSoPFrQwPuuff1tKj4VE8818SPj49vhAbXkznx8GX1+4uko4V7ifsN69uZO9vd
jIjzPQqxd1XiATiIvmvjPpcLlZoqRU0/xzAXePsjI0VtvMA1eIZo7aR7thi22GM71uNL/iJuEb7C
XeFm7frXqBO9qu+J2knQJXGmbryaV7Uo4SXe4YPw0ZgwhcpamFBZVl2Q4U5TIMrX8fIwj6s6MSgM
4bp6TZSz18AXaCiiac5D/9Hnn+eDpbA5X6mqWtT+Qqq00vyTSgsKchor0SXZJyAVNAneU0DFY5mc
zY61xdCfc+adrONY+7wjMUXz2i2JbxTD8q0LE0q9TcA1CXccWaPlCLaH+bFUeb0pGdz2EApGTr80
w+DDhV2HTs6XiWk+J09tgyqav6TUvLTcwOFt5sec30yxzN3GaHnCF+j2dLq6U9DHErY500redrVk
a9JfFYNwm884gb+oIyQe+RseUhIvnD1cDmmXLv3BKqi8jpmF24kr4dloz7qKOIdRYlXpyFUCjBUg
B4PT130+Jk6656MoXgqV8KHjjj9cspf65gtPMOXo893H0csM0s41a6v7cDPqnITK8Sj4YyrmEOHS
H9Wkq44c51UEuXmi45hHn5KTrI6LtZiHlPCOuD4iUDZ8+uobK/Z4y65yjQ2vVrq6RY0yZoud6hmd
ihq6ZgDSm5l6T8JyR64r5nLD77nrFIaQEXMsaq/C5IOl8AkFU9ZeEzQh/i7Rc7Kn1CyPC5A2tL6W
jPwPdZHmp0tHhHA3ynhRMns8+Tx26GTV4RGdhNHs5PcM89giCUmGkU2H2xixEMO4iXDAkuSKlenx
VJ4C8tR6t8sFjIEh7wvvNkewaLYkFR5i2uS9mLG9Ko7yJV+5W9NvQ+r7Lf/fj+Pdgg1unombv/V/
UoqYC7NnCDmlTkicZLhVkISJPSh2B3QUn1tYqbR61QOX/c60qc+1xdtRLsqnInAYB8uHmdYvi2as
oTdJdr3wvK2jfnGSclrCa2IXPzFfGw6Aln3Tt3YP1pGNliiKUl+rH4lHEjH8ktEvZ2S9BTZjxMnR
tqGhFs0ngtrYmULTNvW/+NVP6xe/hCirU7QlhEze2EHOvhNDN6f9fnTL1fan8IsTk8yCLBh9lAPg
q3TuEQU006FrKbsO4PXQ//3wAQPW6lj1uQVM3W+V2CqwImS2V3ByMCwMvC6NfQjjNbn1zLQSkaxm
o8ydsLyYwvyCmX0Of/t97Z9cyIoEmD5HMKlsQdTPcSFTn92bPzVpOEE0crgjunOXStz+7/+PSt9U
ds5DCGuhWFtlJi0yoiMRRrz8swfqP/zP97JhUOAT89PmT6AapJUITvXvNEkkk36UsEiyMSwULpgn
h9RfLYhzpp1fK0A8EwJ+MnKKjPdOflhxM2rmji+nHcdvKUjtsOOR2KNHDgeJrgNDmfFYBlTbYKpH
sXhh9D48JVcwD1wLbSYim11KTg9A667QaF5nFtNx6NNMN9m0UzvS74HUomZoebc4zLJSVdYOHQlc
WZvpv2n1CNg2HqEEP9FRAm2FAstUKEOOP5rq5c3f0bqxzoQWH8HrvZz9NjTAnUofblvthLyRbcJ6
beHj2S8Q5ieX3cxYKmGpl5Vvq3UqmWPJl1+LiHbafLtcO+doX0FhI68pcbrnJu8oLore8p2jUSgh
koYuurGZ9Kw5iaf4agtGeypV5lWxCXuZupLispqujw8I2+H3oHDI8AZyKpjV/AavZjX25zyrWpWX
ktwWVfLddCMJ4QddJDTTAehfQDqUhgxndpVVfYmxJ8wLmvg8Hb318u1FRfCl6366+yQqzSlGbOPs
J+9F4SmDUXeB9zgidYKdfZRdIoIAJLhHBVvXANq1p8zZQjJptRJECsa2HaCtI3af2kZcHhTjrLtl
Pg59kYpQHVC1dl7GZ/wwa1WolSnevM5MvkdYqkHMjdn6MFf812fflKYjSoReb/APrXjCuFF0Zq+q
GCd2C4RiGOs4560XUJbOjKPk6l3cYkx8Qbt3zMydjE34ZN227dKAJ8kTwb/kSjWqbIEvm0qwWQZx
OdAu9PFFScV2P9Guyi4suVv14hZOZGmWMDwluaNzBeEqpqae7nzb6U5m21miwGS8hh1SOYFHjFWf
Gbua2mEhk6mVnZkBJWdp2GISQPErpFF7DPNznaMywIXTEk6D/iAnAMGlZ63awgAMR4C+6EASyPjh
TdiXLLjXhu5BpOeHou6o2F1+BqydHzSWXrXWm5Dw150ve4NduNiilKPgCGoNsQH6k9Uk4pogb7yl
DbDHmC2RNBVH3Z9kOq7TSn9Fj3UuV3244VGvHMuoJWTldU1fRshtS4+aF7OAq2VycePv+cwiaIeu
oqJyPlM3Js4B2aSYyoeqG1Fz0QAoIOVE3vSOXHPFgVlgtuFw8VL175MnqDrfCSlxxgHqi2wqZx/9
+KBvmE8kBOGZ+FylGRHQVkJgrfzrIyLpRPN54g+W8K4wAVVWy9iygXFtk/Ijp6QMrIgt860liaow
asziq2vbGnneuGW/0r1edlHTOpdfbPvOBTmwvLOvu72D8qpqxXrGIcVXmLIH7KojcG/09pHVzEL4
7Oo5osa+u9fh2YQx0rtfS33QyC42CYJCCEj9TtViPxlmzkv2SvNaQCixTcp7irDeDApDQ6BPy4vY
WpssMLyKNbOvFJI/g2hIKXxgi/HNDpCJ2Kb93GyHVWGTU3hkhFYpDNR3yBNOhRZPRADSQ5lbfI2v
aow4uuHBXRteWs9knj0s19Y5keHgOCzLacw9Eqnf3DYqH8ZwWkP3Oyk2zyZZl/ZhB7fNL1wb0sX7
5oC+82hKaAhiuu98RYGtSTffGnRfafR3yk4g09gaoEFBfqPxGyw+GZaDVMFuIsomSkpnAOi+ew+R
iaGbCB/pf0wMOpgisoMM8OBtsvrlc4cKgBIey+ndzQBeAEgyJ58N5kFVUhuYqdnoXR2XAmMponvX
eRmLu02AVaMWNwXg1kXayBASwaK/pjor0ifXcERp+DukRSxa/PPw4cmiBdtbu0gLtfDZgbC5z/C8
eaPzH81YOYbYr2MpMbRIEli6r5PH2D+Tkqg2WXDxHkczc+Cafc/G+Cp4fl77nYcr2kgsBQtydJmv
FE0Hom8eKUwM6KsK3a/5wQzJtEPfcSlsp3XiffheKinbRaWziLeHZud6uGIXxO/42DQHz4xYPBny
mMPWtKkKq5sbsnOOSROTh+8TbkLa3q8/wzAKg8pPD3QLG+cUL/bfeYDTCJ1vWjExmVvYbF8frQio
qg/D0aeVPWkEbvm7DztS5Zt8Qzc6E4Y4xaEBlid/Hi9x3C/+GdE8pRYlU/p2PEZ8TdWJZKClihNV
tA6dqg7fVB+KsNVQnE7ItN0m6cmbz/m2Fpb4umgi69guhWPr5EkT2mpbrL1QmGYtfcVJSshcv+sr
d5kVi9V5grsXGDqRWsHyOLflzxBe/JeaMryv2FeumiCBXOKsgEb45dqQS1FPMpYoaGBtnUKyBVxe
Sj0hLo/1y8ZN0J40SS5iG+dFwQCiZmhf3mtwh7Lz4oNI5hvOszKVTGd3lKhViWaF2687fhYILzfq
uS0pBASSpGcdYoQDHWP5ktdseIgrwmxYJU3mb3SZWfqZsugiR7XJ+3F+1ERSexbUt0QG8CSYzY5a
jwYxefou9DWghRLvhj3oF5LHyHTf/ToYrjQLE8qjG97DFFq75h45pJ/F1W/Ysc1lqU/pOjLf6b0C
JYvyx9jTWG1MJme9llthBasfLCWdw8HX75TVl9Zi72+1qgMKbASv17gR8ghR0WXgRgq0JIFnYIpZ
IhxQkVRZgD/RTtd3Q7dGw82aObgbgkzSlmGlDpfl0806Eas0s9SwbQ78OrgF9ib+fBxAkq+vpQXr
uGmm7XxSUbI5ssdV/LIhxJo4TbWf4bpy56Rz3kqAGRcqUYksaIVNCnjjoe2XiHLT0JTAencS49Ar
Uon/lAQPPn93bPPPdEmF6LTjSMAIybzeYuMEedgmJiAe9KNmWgojBOgQp6j2ZX7C2DZ2Ykqj+Jo3
rcfZPJSs/ifURsDXVuHmvUx+9k9Pa6uA9Z4hwVM56jjcUNXaQOzTExi7hcUz5tWBlL7QE/xgrno+
9CMF+QoQTar1oD/5a+WlqPeIpKw7UfaiJHytNowuwFW7okLGm/wLWbee+a513XEYdLwkr9hf85yI
+/L91ss9kFNfwzSYAdfcYqF2Z7Wa/FUcr+bU9n/iyttyFr1hOtiVtqX2o491TB1WgAvxGze9Rx7A
lwHbeRkpHXn2zpR92Okggpyxv7xCvpG8uuwc1wqvEhWijOy7UCZG2maoH87Zj+JkgKcBfSImRrb7
Udpa6HW1XrjHFA9Q9Xfd3ni0wX9dcJIBPJoptthHjPjvYUkrANxamL0i/26bNDyoA/blMZWyqhfQ
rcedj9oFdtHOOExctEVC2T3YqIIhPjPqwao34vsIEFDK2ti5kiU/urDPV5ET+ZQ0Ng6Opr+GvDTq
26rPv7tkgzdmz9bes4jomm+hO6+/zyo/rutdouvmWXKEJPfz0GNb7LYDHaAg5Eq6Yw3otu5IR+DI
TsSJE+nakvzD7e/TBWH3cOn6k2xcfQPF2SjeqhgxUl2UY+IoyM5AcRuMdCVGvCglllZIYuI+RR1y
oUaEmp21D/c27G3ICPYZdQTWwpXgYsL/jL40q4V1tPeqdJ8VCzpbqfTORDRefht/irLIFdiZAIGS
yxidW3gw49lxkGKFElh0+EwqXvcQMLfuZeNabSQkm7EmQ3Ai8rNwLMsj1nSOsL33c81lYEYhqdVb
i3w/RiMfSoMn0cVLWC9hUXpe2wIbUy5Dr7jwtyCsBnmgIqjq7bBGuJzRMwbQOWBpCoDO7tnNopnG
x/xWg96kPRgee6Is1/XsCPSMshe/RT8kJna6OBM7UVDUwMNUXp73dht4LDmWs5xUhsm5xdGQpFef
FmWHH4xnSdTlgnSGkD/BI6eLSgO4SvuMNtRM6fefy+ENpfKCM+A0OqEuB0wNXXOr7S1BtRIwId3l
2CxAKtOu4chdxhvwby+1ztZTP7wnNPqc/0iIqAYxsneeGwwWnQ6hcEWMfnwzjt23L299Nasizbhy
aUe021EQTP9V5Zv2FNNzo4bAoEA8uTtQOkOm3jV0T3fSjL4TVxGxWIKpfx9iyQh2Mqb0v7q7r4ly
xAGuEoQ7Ogwu6GJ9yp1TLfGxX3gMJiUk0eZWUfaefTqAmFbRSGr/rUrQPz1lbUTnTNvx41g8r5yd
7xcVGDH7yxCKbCCYfIeStdeZyqnMG72ioZXCDeLBZmat8qpW8sVqEUi42ZWD8YKPJxBhg59/M6x8
1dTG+PZzYOJq+CLoZP82HZsuj4S0DUJhzUobtVSUvBKvoYGsCS7ym84NK5jz3eQLCly6SZ4WJd14
heOLXXk7MdzDBlakYxz47uaiYaoVWZGnNbfUbmFR9cUpoKXFBUF426PiVYi8EEJ3Xj5Ua/5V8Xws
5Pnb4iM/SJV0DmkwX+sLBHDvFckSXZWRNCdTEcbWp/evu/lBX2b0mZ4XkpxMWSqO1Lw5Fjvm84C1
C6p7STiyyeb1FZO+JKZQQsnl7rp+LL/P23JMWBoc3WCYhk/XNDJDMEsubXgg4MNt1Sk+lqW7hJuC
zamdNheiXfGXzozIOYklh9mSNy0OfkKEO4/sF7LbUqCXjT8wAW64WvJY8ngDmGII9/0fzP29YO2O
Kjz8mf7/FnQfLxqgFzG0F5peYFDskZKpa/+CpCFQh46CSTWm6uajcKOAv4mnRsDH9fusGqRj8Jcb
E5obIY0agfSnXwbapKXZxRpfTRWYe0/9aPAHwWFMKahX3/ZyKjDrM9VnB7E+30hwgBQuzPWN9Csw
a/xHL1QH/Njy9gxmNQq+ydmEBduTsPJvdhv5GTlrDD08lw7VLetei7r79h5StAXKpRPuT8G15qeQ
h1vTC9yidyf1/03E5TzUFfeYZC56Kat7NjUwMe1Uo581ENXpBSQWDGMy6fi1u67PPKirTzy9+8WF
znPJp1sU4K9LSEzJyoyNiDeXSIYt0KdiNPYmrbVniohE48kkU8KrzUiAws2xZh/QdRvzHdmiIBgD
JMcXqylOYui64D1yZiC7IQLmsZ3GZum6zXdv5GnNfHWF1uLcxBYfFnxwVg4W2KgI0Gupk3jE6URZ
5ybt35sWqcIQQWU0HCXk6CvkCKo8S+bPWeo1eYuzy+QEKlBByjeFNoHgLrW0qiLdDX9CiTeSj1Z4
VTaFu21mqZvghWsEOmm01UTyuAmuHccaK6DcZjs5Vc1gsWeF5gDzIHmKkEDJsOww8r7yU3P3Nu7G
uWiHIs1EI43kb21fG184HnUXnA1K/+t7Nqha3ipWNiDkTEu9Tt/7TlWziahChPALY8ECDTMY0rCJ
VlFe2GxpMP2r+sfvaCgjaCNoxVo4FSqfHF75qXYK3HiT/gOc/Qyx1izoYEqHx1yo582C3RMWiB45
sXagzFIxKy+d5KILcSvQwWL1UqOQQLTY1oRRN1I1TfV6LkM2hpAyNtC/G6YJLf15R5NDeY14oIbq
VgIsv74qKVG5QlT5YuG50oa8dw13HNlLSkx2iMJUz0sjCT8y/ft7X/hBaw3cSJX9RfUm/lgAASCl
YekdG4hDZIS9alkPg5MPW1L+fNGhXFKju4X8rLqIV0jXjwWp9VKc6SYGkFMaQzOeQzTPyzjQo7iW
bnmilvRi4qMZEOvizzXIe5LTQK97idcgTgd5w8LINjS/YQt+R7PmlxMF+Gp8VUiXA+68s+bgsIVS
ZgHzg8Nhazg8WWq7+9RY1+dKf0ZV6IK0OLz5X/pedEMLnJtDI4E59DtxAc3U4CpG4Ns0b1lXE/1I
fIyVtB2Q3FbkcNOlvpC7kB8DOWjajkEZLOeIWfKao59lfccIrLrhE8iGiA7avCH3S+xV+lU+bMYw
QSlWmXtZE5o8Jw5yUC4cuk9JVnMUIaML69BX0GmAohjU/1OGYEiwPqA/GqGIdlNOMnAmrUP4WNhC
6NQTWCydgLYptURbOf34m6Y1Q2iljGnk6tdCho0WBtWdQtQLFMGGdc+1gdwfCAV1MdyqzJW/5ggB
eR+kiNb7o5WcpWWeABH1hlXOLyg/9vzniPWoi5tVfS4bR6dyEAPqKzbxGEGO18jwSh/4ZY84LFVI
P9IpVsrjS6YTC9/D0BGlUitPNIrp0T/V7YrWdWNCcZwbpFRPm6fGJF9xQR5mN95OP3kfmQ/hmxL9
xjcCpLJzHBruUirKDR+TlxzmTUiYXNvdWsfv4kKAHMGV/Wow74eByQ02n3C1d6U3E4sF2PsG9pGx
20L9g6PUaNbgzbqTM6V0ML1aExL4xoOXco1fLPvarE/Muc4rDqi3nPeB/Rvk9Zw0TTAugJ1mMozv
IGklnb8E6nHiOQVbzJQqDibLvX8PKHSZ7f9xaBGg4mL40LKP9G/DT8NsVyLqZUXQTvT9ozqgUxfs
iUXkBW8kNdUEPG56yq+azoEA9BMzr5Xf3Yojy+dhgwjvw5yhGUBYIfi/D0GG6Ry8DQpqLpjlfp0c
9Tq8/H7SXRA+HXpO/qd893kSFOUEQdwHzbD8uBoFG3c/8urrWsJmIFHvL77CwaGZw+bgHxUy0601
J/2+80KPJkRCD8lwSMd7dikKSOLsnyzgD7HsB4/nk4qOmyeok2FQlva1w7qHNYJ31i08vrektI/E
8bRn+BxwSYP1mUXNJzHEKXOb979ZTuLOC6oiTPPydIH6fnVWog6C/UZd2s1aOaUo0qLBnCnrmaAK
2etxK9YnPoym3PNZ4m4ex7cazWjnHTh6mx5RJomCAJs39WYEDJHdpiTjy96zlXHnTwKQfkiuqSU3
rqFediSY814FXPEnygzJarRp4kcfWF0dYlKbVWTcin8b+n/vZIBljRm4eCpWeuYn77I5KJTRThuU
nFkmlB3/emUy2spHoHbXCwnchbfzq35AmncTB266PvCG+g0jHZNuCU0T+TvXdJBAofk0+23hspGT
KR2RrTeOOEaxOJGysTRcPkRPqqp6jhfkjw8zYsmZnInW8iPv8pND41RCrQte2hacrwrAx/kmz3Zo
rikgNjkVHOZIuwcrbThwdhkeWnunHghX7a/OcnvRzPJIwxeI6r9gLwSuT6aiZyK19Vl4bJYUtaKq
7JpCKtWQ1Yup0zu8CvNyY4LKwc6ca4gpryXTdjPsut78XBbQzllmv+OsnLvoLwFiCkqA3jMb9IeT
OQv93X+OX4ur/UalkOprIST7RzBk/kydj4QrzZvoRqFJKe2yo/x28pGbn8ZjBbmieP+f6Aa1GhqT
YwpZ2Yn0CzdjO5qI05Zm886vPVZGokzBj8NunRm3DtZR8EO89H9Hxkjx/xFeIkKkkTMOevA7JY/Y
iF60B3KpdMx6eqdFh7w30A5w+wmXFWNqMPAA21L1UnBOG2u/bRO5K8VPpbs2FCDs0ONbO5jx4W3t
eYnpDnxQ9L69gs+BqJFJDlNAJc0OjsjAPiikC627xJVNXS09wecB9aTU0Nh+EyqP9X0Js1lqduTj
cLzryqyfbvtXAfMFl6i5pFgtenqMtLN+xBO0/CKKEDDxiqut21d5VzvDI+guX5n0wNO+r8Rr3qdD
PC7TLHNC75QeXdi26UV9OnSUS3EJRN3WNSDWcfLeqchMAFkPeopFv2Pu5Q2xhQ2yUVJVF0y3uV0t
v0+s53XMil5NLp/Gj9qW7EPlNOpMk8IokDNMxX4BOYzrKttE10+d34zgNDtzCcoa93+J4zyUznuW
/IlIByDHdiq+3zQMPedc4y21aJJxl4T8kY8/Rd7wReUx4X3GOXS+uz1gqtWrX/61JVrZjT2iWvFL
Mlq3PzkAkltpNixTItH6HGIHdYIjxTICvGg7DziSftl2bt5RlstBI0kx0mJNZZI3PMt/mbI+/Um3
rMpc2RfKODkm9f7s/qiG8odX9r4RCr5YDfTdS0YoZaoUZKJWnTf/I2ViokN+xrSzoL3wtVNBS+ix
Ml/oZtmrVYpUK1ssiTqyuZfCqYunZ0B4Towrg97+TS1PeWZbooijxjPXX0mgMWaBU8/HAVS/8iSJ
8nrf0FNSCux405uOAPRyAAjkKVqFR+UObPXaJONIBflzaL81PsnoIR360sEO4dHmfLq9GWxBaHoc
c9wqX1X+yEsL3mZwrYWSeJrGW5L2BQ/Mow/IZxKwxLrWuM275EhGrvGvzKdxp2p443K1KJ7E2mBn
CLrqJp5FBK6svOrbXXVZd+580WghjFHImTJ/EfHi67g9ipHrGgEmLGL5PI6mnDSLQ1ZIS0DIdofb
n8GBFRxzTIMXLwgs3uyTj+8Fdy+C8migvTNG08jTZ/a2BPGuy6WrfKqzPEwl1VIzaGEs3JJxNwpC
WNznxh/QSbyI2+mVUJcgZdNkbDdBYaUdyrzYiU4NEKgoHbQkfEZ6el0XJqQyjZ37O4FFBnC1NBSh
riGaCdxewoAb7yJ0z7SePuVhO4ISjridPdGZ+hTRRjFTMnpNA3HVdSQ7cXOP0w7c2++7It2cCVif
LkHRI5dz+ElNZpcUGYbizeLT3l+2JNQCAyihIC/BUi596Ltb4oIZioA+2Q/AgoZmadT5mb2m7GT8
KWzofyrG8trWNB/vFqJKY4RaICnfHNYkLm+F9NIeeOBV4zZNd6toU8uaOxxmVxMOJKs7JmrhtviH
puQfaqS3BGT7G3a71Tt3DJZvGBKh68PTEoAkicVpfOCQLmGnlHCQX6BuRsItRj9RMkBRoEN5oblH
4WjlQqtxrTTTujg5JJvh2yJJH0Xiu+zUHs2hoGK59l8xCt2tjCmXYyhZU8kRuOkZmDAnC+ifqf0E
qf17c04XVagQA2HFdL2kg6TlvS7Zs+V4nbTDdxFygH7dDTUng0ScSyeNPNCkIWz7hoP0BG4ai6BD
YOV4WtcV9YgvQzGOu8ErUG5Dyblo6ZvxhcwTXpTMscw8F+iJwoE0fCixekcT+iJQZEduG9nfFSkT
ZcxW6CoiATwGcP1VRCow0QlcHqHMIr7NPTRFIzZWsX6UXdgXzOks/b99HA8XdcBmRXSzqmGEGoLB
dwAcdQZc3vdfg1kyJJo3ZEIlu7vPeQ31wsSLiMt2aalBQXB1kTbip/1bIGjzKaDXl17w5esxUo4W
+MHEfkpMGdQ/aH93BjJYxWuFnhj7/xmnRc8TeOSUseYFMefStrEnMFfdTnOkBPoKgxeupB5Iwalq
n4b99JOf6EUre+1LZybb/JPGuHGSXy0CfgGAtb6nx2AAHvJCf5e4UmlB4V5lI/gojc/wia2noZJG
PgUklifaY90WrE78mVIjffreJlfOc7KXA0tqqnKdbuBgIMKvenIxtzb1DOfF4UoL2a1qDy6m2TTf
LXyKiiaNQFZhw9hZSKbYHwYmAKXPlQnwNWaeDSLO3GWXa5R3kbLkM6fdyfmJ8XFiOrydM4itkHv4
BT3+dW8PthRXjcJc6Od1sTvbHm68hlg+rJpw90XIrW0+k7k28r+Tlwkb1VFP5eRr3J1LO/ja5jLR
ztq5q6noQiSRK5wy4BrJ6QPIxD9NT2lqMw7cdIfv6g1g65L0+FLXox7Ds5O7BqoLM/g+vuGvs0+f
vvwMNRV99EbDUh/jVOpukwc7fMTWpQE+YUPrkZOBP1Y+WLjmoSdFied4uBG3ytik9RD0Akp9/+R6
6UEdCHTTHakmKbtI/Ei+VntQJv/JZBjdKhuMlvcIe0okQ9r5EbK7bbUkJTgnemsj7AlOtgV2xBmP
iozgslaqyL13ojWfTEAp8iAluYjRkCW701HbSsYTwJe1DUPCdrS/u+uoXmt28SAUrdtnRtb1dycI
txTN+ja3Eb3/c20md7++q5kHZQngonSp8YavQQ3vxIoQ9klqa0+tPr7vqA6DkrXE/nS7FHkJvOXx
M7Ld4l2qB3Tj5ynY1r4X67VPem8QNTm8Ayg30NBunt5zEJVyi5n0d/doWzj4aBJl+9iks5xXRPop
Upgl9AnkoCZ7XXmP2xDnYAZ2m7ot/7YaE0wVwOF2N51C4TVbmIhSwANb0NeITwQ6rls/xjn1eJ7k
8Wps3BQfWQWKYqdfIyVo4bsZag1udP8XsLLPGBbI9CsxXycVNDt2FJESm5XIm51rPrZIYdbHhxuG
GauhK0T0CvqioKoa52JO+jBTvTyQ4iAi+Fwx4jyGuoaNYa7u4mfpJrpWM8BCPJ3HfIfpdOfAhiOS
wHtNn+xmT/XoCWh2bmRt/8+sdOXIMswwWFAJSA7Ezp0QTCyjRQwnN/7YEuvyGepHjBF2LIYBXrEu
eXVdLzeHJPZZ/YDnWyiFg7WEnuTnTVNlIeoskaUBx5tWRcCekrMG8hNmhgzZPClLkbAEfW4xXm1c
qQExVhJxDpdOFm1yYtUinzeKtPd4b7YVKlqv5mYAWMXJ6vvVtf0e56qYZFUQzRaZ7KR5fIW5aKOv
HQ+ozN6jbVFKDbgRtUfxN460GY+WDOKlRJPW3qy3QKrWNGZzaHFXcW3+Hj6fOOeQ+Jy8o6n93XAt
gs3jmOQc6C5BT0ZedAd2ZP0g59CBRmr5BqnXwKNe2AjOxEhj9Np9r6L2M0E1KEkQqE/AUrOHPU4Y
CvOyVziDE5O4bkgLfgC/U8RW8kw39M4Wqma9MfjB5jlAsrSiQ1XHmuS+2rweUvs2hftgOiUveMX/
OQtIDd/ZnFW37wJggqweRGVzizYBYMN7DdTzPTZC78P25o431e1UpPT82lnVclUimiTifSP/lVrq
CDs17NZN3rCDnNJnuPbIhxu/XcsGwKg72xF+/5Dk2PmlEFPz8D5RCd1I1I1iakxEbezap1yBNmfF
5aGgFOCT0fa5vkb2AADblxh+5U9jjoywk0dGfxhxb4y7K6fXJ9X+qpuEsIL4IiB8iAOwP5ZRRvaF
KzTH2nSLLEIryUtQuFOikyygn6vCvQYVjnaDTyD/iaEvmT5C/Eu/OfUZsGu2kPwRtmW/5vOaZIWa
ljyK/V4gJvoqrj9VpoMQ36m6+tURDyFrUtyu7jrYsnlxhQqA7uGXZrNxzU+SRi7PCcFGAGyNOUZn
xjCM0M/g0Sp67XTZJAdqrYeLqqEoezw99XpR+12rOp0apcaWfrIzsVESZDMSMOB4KjXMplYI42BZ
juQ3xUXU26PIHYyX1bhA9A7IW/skdV1dhF93BkVWatHUGdfjL6wAy5FtOYkaTQPkNCF4wfliqG1F
OkHhZkginEe/FnxdbMRXL399SGtBoiQZ8tb2o92mi7LRmCNKLKJBjEhXtrzVVDa81suY0FPwJ/M5
jfebLnT5gBHnkIXR7mtl/ptjde2Qms3WG4y/HrBC4+2Jw7EtoWgv+r1b0Te61CaxaIcpX1oPcqfP
xzGcMOikDT0f/pBjrcjUlRNmi5916vdA6+Bo1CMuN568oUdMOLa4l5avMipMUnod7Fm73OE98+hp
dYal5S75X7eP60J+xd4M/soYzUUayeDeoKupN0CHIHwprr3NBh/Wp5XxJCQATDzl1FNhtjTLduyO
7tyhdABFGd1FDsyrqnYBzHkjm8R00lztxFnW0xAx/HLsx78m69If9DocvipGjKC672Dx92chwHY9
Q2sOvV8dPE+4TibzfsmLLIZAbA6iULUaPviCLKCPvOKkcn9IJj8G5p33tP3kbxK1g/570L1tsAqM
ineNBBzSsjmLd12mpG56m7oHku5c8ON5+YNqNiQ4fhsBig2hsgTsL4LK1QipSOS1ikFv/LHUeEuT
0dMQAFiTLWgnxJra607CDAkUDEH34hn/LGXjLKYWC2vB5p95HigZpbu/Us0mZRBu0EvH7HnQfLWp
uw/AIzymjvIkVW5+8yEVj+M7eruwpekW9MDM6qR9mzr55/mlVYKiDDNeT48tinQ6u1InuzjMwZ5E
Q8rIbguu+nFcBq+LLc5G2YT14UupifWffPfkPA+eff7SUGukQjYJu41/QU7jYrOtN+11y7Rtl1Gw
fui54x4YXl5fSXPEGuT09n3WSUNTJNQLUhM3fP0YLqHtLhB5Nil2ZIYSOZ8NDUBNdq7m2fWFl7aU
h9xN2njifos8AQMDCv0Tku+ahgYgmrk3BoGQU11dtwZRf3ltYZMqvLMAL7bYjF3eD82b4FUSiiOJ
j405cE6qiuLDjJ0vIazCFkQwZ5Mg12cmKbcEGPmKWYIalXf4OxUuRdRIBi9amtbEjQh2dOeLttlo
fi5143RPc09FiWsVOAOyPUtYU0u6dwNJLPFGeokiD7N3ozPTL+yFSTvpMHoFbWYyde6qBbTACs9F
6+d6R0XJrIr5YACgI9W84NAmA98p4U7RtMYEsvwDWVf2rp5nCECdEtIjh0xsSAQYEoC2/KZvBMYr
+/WFFvCXraeahH+wqrFdDf9DrMzhUL/RrvMcJbR+/DiJ8oZilBUh8ZbAgSfFNK+uOXF4pHjPoNZX
TE6gUk8TB6aZSKcOQesR1ZWLFpyN27rBi/twr91l/EsnA2SXeKIdFuAN+o/2fhVC3xmFZUUUyk89
pYbSAizmS3fnT2I7ve2FkAjHHfLPD+NdmZVY75yK9O3QVQa6a22G1ZozQaY6aR+9YFNV+yienC4C
TEkIIaEG/p5Zgf8OutNslfGMRUg+bjOZu6ZGSjB7rcFr4bseRRITF6t/Cm9UebIwu2BxJW5qnYZ+
f25BGvkxSF2pmZpoFWlFpIziY11vOXYtJEsDBQpSjwu8VuXLVGEXqMzAezibSmdH6LRttKSQY5ky
Kz23+wKTPLCOcHk5LD9eRxcekrsqIA+fGBmk1ZBITKphSQGUsPzzNE7jCN27EC/NNDefyCL4eNRE
uz8pR5XOUyzW9alsBF0ayFm61K8YflkeESeUPKCkhvnVgYCsYsyv7BG4Y89lfQQGKrK2h9j7FhVl
f+LXMrdgpDge/3TRnbGYM1BEiqP1uGh7TxGppaHwn2FQTQ/1AIQIXcI7zPDj99TB6iGdDEOTsDqU
NRanQwelxcp7FNRzPitbE4MFENHCHZ8wMiB3QXJZwS+WAYxxe+fTjJ9OHUpPUAH1y1+18t/BWu2j
jPXRqfNAaINE8JIOsiwarBK2pkgfO83qnJJX+E203Kkhe/bDlaedS2s1xkgxY92Is2Cti/WLikmt
gAkeSXN2mi1HSAmRHZ6UMGO5uOn18O26tCRqmy3c641wAJPu5WfdzdTBwT7fpDD/PtKj6aHt1eb5
iIWSzLBMZtXVVWeqfwk93N2ynSm3cl7KWlMl4i100/GCh3yV0psO/4oe+6sB7/oH8a286G46FZdb
B8niLRKk9S1Yy+i93GWlSUdGvyIj/5+2K5RTYvprDRmhD38U/5GIPvfa4TiY1UFkaMIXDsO3y5T6
5+Wix2w5/wVcfTtvgYnO45KrkIYk1/R62VXrDMiIteWU/2Wnc74o03jBYmL+YwOvB5rq3ExbGn0H
B7ExovSEwQRmNXINObQlf5jOwyaF4gJBGzWel+cbXlQLsLsZwTxxPHcgBPemRaDhNDcXRCfddZ0W
TOF7YExezFsHUHiqxmPGrQ3n4V1GOprTlbqU0lWzmiskvLyMgTsasnp6xw2Fx++w8pzPOpFvWj7E
XiteuH798zFmC5AFnOjBrg4SboiFaBmNCubf3a/Y2iLCxNDwwoGgiju7d1mIUHLO5+rCGXTua/h0
el0u0jElUeZZ+nvgTds/Jk9Qb+MLZXBJU+56xwy1Vy0oQJvnlbLBUtFVTkqa9ebno6momf3tUgux
2HaQuvuBtNpOTMcfI9AQRSO8Jr/6aZAc15lUHjI8KD9a7daxPO20wAvZ2cBgM1GPFG3GIx1t5NMI
JI4kVmkBXvsPPTI4Cs9kvkWtMCs7Ar+itfXu9UCPxTa3RzIRj2DU642L7MFJ1+TS33aF1lVXLLsP
wOuMnUsEXH+pP6OL3lC3tfcAcUtmTjO9aDSONmF97N3TpSVhzbhE7+zRlkdjkHMLgEO1Lenb0W4f
HbAmMyLi+2gYCRrTvaJH+b2CuueyDMBqbLla990Ehk5ez3aJaFCGm9US/Bd4CDIYTAqb5R+oGgoo
hcJY6FyPONR4y4xbSIsVb0CoapouEUlmTsxwh1QgMz1KsLWk+CzRkthPmFKRbAf41OQpC5u0Lipi
G+WLkh1hk5D81M0jt2pIACprXZGegugVbxgmIyCo0du60q6JeeOdhLv7MJDqkgFca1emR/hGas7X
6151KctQr9V/ZeHRkOJFTUlFnzlQ5mB6Heewyp4P9xarEbzhoWuIpLLNGoYY9zU61TucGjxvob5D
97EiNY+9FP5jJ3YTcdOUm34xEct+1DQ5LFH11OTdFA6SWUyjhp+UPio+zvRC9FFsV15wxwQ6AZvS
Iatdf9q2v6P6+ZYuaHHZU1PTMyeKpSSG5mgmDaYMuV8EL9Mklp6n/aIMsDbnyj6MlsGzUkfNI9zL
Q3wsJ994oM8s1jhmuZN+4tqGHfpEEdXTc8j7ldPzaGgC2cu64QBpZyMfvhWi1pH35SNUjCQ7LWip
6jp+tEayJl3fiBEF4EyltEdXwE9ZUp159nQx3tSy2k8o2qZToyrLz3AyeMbJ12KayrTJTyqzVeTJ
oGT3ZXa2rQWMKWiZaj40wCXvDRtm5dcHGaiGVbWPIoeaPVxmwiWOaR+IyBysWwbbv+64GfyuQD/Z
fDLnjdeclOm9WmgQRaQYruTbDEqWd51hPGX57Z7A9Ah5uTthbx1k6+e4IQxveVO8rjbe0ZVMQSHZ
/KJ1e9QXTcY1HqePYWJhoHz/GIjTfq02anTBNh4EqNx8HiYH5y3jYNg/CuE20wha8wV0tuifoRlZ
2wbccHOGqr3Et03AuB/qTz+0CG42dn87uMbaL+UEIoZGdSbNYz6W/PfuZ8yPjUuIHuaqgDaENW6s
g1qUCrUxlILKlLFAGAO/8uCgOV5akUTCrUdtnuOO70o0Q0JnKq50LcCXvgk9NTjF+IYSCbYXW60j
5E0Vt5diGXTZkeOfBVKrKt3RdVpkpD0R0aSQiRwhVGO94pkFf/Tz9jUlPdfwEmCukHxRzaUVCMWZ
k5Q24FXmZ1qtkh5UbPDJ0nWmfquwDXfdID2dWIXJNW+P+sraXjrbXrhWHdcSMCMPP6+IrKhdrdZe
ZC8QjN4p4tjEvBnr4CYPUJxDz581Ce+syp2z0RIEZ6B9DAMjVmN+CVl3U6dnUDT8fWSgj7bMBrJ1
kWbf/KCAC6Ggs8BLOeicMzBahZK/lmAzV+8ksJzUfYaUj+r1Ee8eKHircUgCwVfkcfWxFxXb5dzk
kbAdPZ6CNdhtKgMjc0NqKALH2dv84o1UPc01XI4RdesTAEJj+nI6oEscBz3R/C8poqy7tYClJI00
qgge3rl0htdm5Wr+RaH5U0GGUEmcuV2mPJMDOeoF9SAaTsfXJzUQNZIJu5mZuirykZIV7VyPFDYh
hm3lGfyebv6AJaOuW4DSLCNXQk7UFF7gxQqwA3eun1GSfWKnfQcT7R8PkETck2+Y4pzTd0AuB56j
i8U14YtLIx2ZzrcTMR44hI7RWNBBwGBcrOM+/L/T1e48KA5JNpMLNziKk4KXO3ztl7ifyAGMqkXV
mp5dpF1wc9kCuxx0HMk2PuLw1yRERZkoSyTboOWzRFsDjtZ0DvMdCb3azq335kLMcd12QQ8INQPj
Np+idJJdjx0aDE26BmHv2Mdtw06EqktJ8b9pHF5Bsvdbpf7U/sjhT3qwXiVquD29NXoFgOPHheG6
zQc2MePbVUZgknWuESy5uhT+3xWbgHvmK9ca8gWappHskNSKOOXu18K9OQV/VIHqklu9blyo7HEq
iw7u1aODLlVX7G7BtKlhh3ezz9FRkJtaluVJqSuGwGdJJUwOQ5grQUIzhFdLu0+q66M6FJ6O+qTd
7xeA4c7dTOY8rLAMxVNegZl17/xtx1dZKjWjgTok+V3swWyOEUBoxKxfii7JVj5gOQHTkJemUYyx
/LEtd5hSn7tmQdNPvFRQ2/sUD3tx1VCdg492aQrH+GASyNw3btoG3NYX/M8xnQfH79Oa8/NI/hN+
zwJbisaaNp/Em3VkrBf9j+c0JayQOPfPgImAiH52ZOxnM+YdvyAjM270LUvxNfU8qUnv1jLkE+4t
8xGBc/q7Ss2dG20oMgYcyJQXUSc6NsP/Q233x4VvCJ4+WfiU4FsmJEngdgjC1MbiSGp6L0hC80WI
vlrd7ZQlcjdSLg8qMenyfCA7SnpIiv4J6zyDeaJ5wijOydCUwzbTyDO4O/JvMSKrXRCtUh5+r2g+
Rnrw0PefRsFt5t/83FW/QMvGiMHkpDLXSkArFNRTCs4+ifmXoMoJL0NQp/Mb1GQz43wI//p7F9Sv
WqExO5EvHn9d0cp6eqrAe5Cg15XO8gtMpCy+8abZcO/I0cOLcAHJ3t1ZZdlD4nNjBdFPwC5v7q1y
NsnYOqi1Iw+U3ML1CPpyl4gXDZVVuaq+PN8hJghbJtTTd9b0hrgztVzJgC9I75yOlCLtgtuWueF7
1ZO6lfgP5MVDdv2gSG9gAHdb3vKT+Bcy3NTovdyonOKdOYFlHiLfdhp5Y3j+2PiXOoUqhw/tP4Ix
qRT6+2MQoSzP00YeU3QLWfLLZnVZ7K6TX/C1PBrtv58+KMcqPBAUqrqeWEf37++NVpMKtlsseKLy
24qZjVq/1EdxqduVqlPp8coH/DcDK3FQJPf8orH+qNPlUFxtIERL7dHmToez4l6qTMHlZDXJ/wlZ
N96r8+YjdiZw9NUBXvaBz9eJVOE3Uo9WOvTo1zs0c7jHrQwqWrTpGTtERfO52SbfxCRhQFoGD7ZE
eW7QR3Y3Ggj1MvVaWHzgZnvOdXg1t6GcPPBQUlV5hJVEArq9hLEcGy9N0UpAlQThITagBCQz0M5a
Z1adkJigIPYDlHKXBRF7Wg8+Klji4UDhKEF49D2Ljw0pOOq45Wp53ArzqahXS7uCW+SW1CXgofTc
I67/vBVsjqrKVidx01FcOlQJcDJZzva7KlHHv1xfjg7PJItbCuPkdyqKNQVhm37EwICPZ2emVyli
YsDaCuV3RNTQLUo0tOk4okoFym7gQctYw8YLyT0sWTgSorsPLELGe/5Xcfi1exsgZsCaoJB4KM6q
3JJixLSi/HHl89GxFSWjym2AGzJFd4EyN8/peJuARK37hePpIvNk+9jgCeI5SXYepR4Vce6oIopo
ioOEsswJPYOaZ4Ccdi7O8hNIMpNvnAEhOshF0el8Ew4fL5LYALfIdgx91x1mmvx3SI5Rv+0QYqT1
cDtYqFE8rzOgoZwVahvNyGz/y9lazCPWflGHI/GmYTwlegSCgODJ4ybKX1/VAty6RwUklz1S++nU
tzhknjz+TnJskT6mwEQoTxMUTlEe2UjbTYe9TUlMW9VAKfTfnjctWh5ezgCM0veUJNPB5Myj+z7M
uBzNguOGYjU7W4ak/35OhnvjF3RtQIB2x7NW2ck/0ICYDLh/+CJwwDa163MAwrIrawOaGR1Z7VqG
6ttQ2R5sfVbF8zrIaewFEopcoGdhrWEA8IxQIHJZnY3GLvfbX3A8ozxMDwFOTQycODPVMOkWiTBu
Pv/VHLC3ufN0BAX20x/10UyRja4vJ85MM5T8/diByRXTIwGDz/GlUkl/YMb48/++fzfowXeOraaO
wFrfo33ZWndCksDa31Egz5H4TTH7EiKcMlnbvTKEFlV4VkV592Q/DJ7p375qNGP791ZTuzCzjW9Y
SGUPxRNzpNCLdwCMXpeFuwTWw1xaid10i8mqNLH7kofxO9trvuk942lGTGgbTrgeoNThUUULllUk
WDQdi4wAi6SqLwbeNCiLe1lICdCeEeQ4q1DrLIUW47TYSaHSwUtCkCN4+i3SW3QXeDsqZhTaOvlS
slHfUvO5ob3M5ZIwjjhowp9aWBw/nZaMpi02wBfMxZ+W6NFPWAsrz1ZKbgv1V+5OYpQ+utN6a+IX
/0aXPqN/ScVbyBGHt6mEc0im3TzOIb//Zj7DFVXWWft639Zm0DDrVcoeEp6belU6992WYBKIQ05g
DDRFX9r0KTayiFsMoooT21B3ayMRl74wVzBs1SrHMeFWb//bFuuCc8fNbqz65QYZQIqi/I6OR2na
crMBYM/A14PMZ7RMPe0hArmcbFW+Tkb0MYX8w3dBI5y5daDAEpvD/tEi24/BIUSgiBoTzVR7RQmm
ZpX5gEE+huGTZEYwrfm5kpERbo/DR5qLcTzEG9RfDvtJwa6kIlPbScNvf/M+JgNwN6XInhHit1Cl
auxlTVa3LC0KQHhnANw/J0FkdJKco6oFAWcr+ni8LusAULbZyiYCeoHFwReOjc+DAzRshvEi1y3D
w0OgPd8SjgPpxeypT1h+2M1QBqsSv5ShccrxukpofyadXjHBXYxgyVrjAHLIObPux5iJGI2Wik+y
XKxCXlfWlZJRuELGH96NaaYiwwARQgWK5uCaJ3lY1uf0/tilMUM6gJ4QB4UiZVs4ACXyHgH13mOl
8YDN6iExSM1ybaOKM/cXmozGzHzgBWOyCWGTG2m6rktTiWlXQ2lUD1s6ps+3hfk2bBxHAMBnDTso
d3+2g93kSKzBxW1/h5rjpoUcpZiUwCu/d/gUTJynuoJRfUXOQn9/z4N/BmE1xQb+sC/nV8m6N+Oz
m66ycITz9q57Cu48jUN3upYUAEi89grtex+94d3hZ46FAkZKjCd/Si+jqPidHRNlkq6IpWPUOZM/
PMOq5wyf9QYv1dBAYm7zs/bxG2N2RA83T3uYy3wsiCd+vyPqCDHtwX0tM0dcRiEtgkkLQeg+a0JA
2eMDU4V7B6LWuSCc4jWVPtMegz/ULwXiimLflQPfElS5xDEobXtJHKKK1/DhIRTMwLtRbl7JaIQP
H5xek2l0idrrPu9wcEyI4EPGTFxu5ZQ7ZkP6iwuUAulkdRlrkFjqpITYrz/CZcxSgXGJrsKBKy7C
elJn7oDUvWMxiTlNQw7sprzqvSy8n5xidbawJ3CTjuzNGXKab5/unkuHWIRuyYQUBUrKCsSrFgQQ
Cf23FQsp9sOKwh8qYAhk9/MOSUfhOPZOkqOt8Xm1JbF89Cv6HqUVcizKFpeUv80WvvBUb0WallIA
8j9lOGYHsQe+TdIGvKz78WC/0CkHm2xj9UfM4gir0XSxuC8PCNq7X23W1jnLWuE/VXarnmCgKM4L
SObgxy/6cZAKFZhHmgqtU//A8EHtBqfNLj5zoaSjuRBTR5gkCBdlDtKoV11FnbDR3pN1G3kUJfbD
1zDoMnmg+ZSh+giLWt0VV5TPw35l+XkjXrOmWiaBjbsdsWqUO4z3H4v0qSOE4XvDjDdnWizwbohh
6uLDLdteynooRFiVa3xyW4oP1xaZsrHkVO2Z2FpBkjLd9ficmRS6DdKCI+NJRHy3awfuj+L+5zP0
TJci/7ZQKLbu/fiOXxvlXugVpOsTT0n21cUn+l0PizSDBN7ywVPdCowHZ/vyNmuk7uDtI/Sf22Yf
rn+7oSE/svv0bQvcu8qsipnPeDFO97ble58wzIGu1leO2yFAxSDk8XKUVbi5rd4WX4DRQooSB/T1
U4/qp9ve75iD5h8MYhqTWXxblsbN86uBAiRGo5QbxFoWiQQ/9/39zppsJQn0Q4b5cB2F9Hrh5KYm
CeRlymvQkz5YGjw1jjmu6t8hVfv8tvE9tUIlQZNrZWnvZxvj81jvxdWW6ByBPeadNQBaOAUlIb3F
ehXJiVTkt8IczUCzJhigdijEkBemvTKxAS20ffCe7HunbDoHXte6vwb8X5A1tFZr55rUG6TmfY7g
6RuGF5jLoc0CcMvHY2n8yhORXOaytuRkmWg12O4zFZ77KgRAGu7x5wPkjlYMMfaDyxFCzapT7m8C
e0m6fzb4I2gpqILROKI1Y6fzsUrBnSf9MbaLgFJd3SMGaP4G8ZfPMolf49nj62/MUod9tVANu/UD
g0dmJbgAqvoePyBAjh1HNAgCPv+u/E9uE+GbyjOIFrsUXzQV8S9swCsFu38wWT/9ApmEZORgHIM8
JExr6Nd3Ri+0kxBMiI/y8EfpOpP4722j/YQa4kIjsQM/cpiuj/C4H3UBe1w2jIv0JGT0GZDCLGof
Ru4LB19MBc6SUwqwqj/Sl33wb3mxpPQrqaEQY9fJ+QFeA9Zb6HOxb89f1x4UczY0uJ7NnZQ8slfW
oR3L4k1temdrw4F/fMjr1DlnP9oCyZyc6heqlyrEWv0BpgpPWjCq8+oEslP7i1uKE8ktA/Sbwa/1
e8tSHdJIRItL7h0/Q1+Lt8tkv76edhGq3yOzf2WHgXgEdlOMyTsEGsniIU+szS9oh2l0tjC7r0/C
FpWuHf8Tl4Ur/BDxbEOMqyZEq4uo/7AW15iqiV1QkpM+mx+oGfg52z1UvqWRIzgeirglft/2uJY6
OfwXkcbxBWrun1V3yN+wBwFGgw6W4hmP2stqQBwa3Ehs0IW+AoqpD96zhTf7IOhXG4PKxS+nk4UJ
q6I8QBFAUsWiR4YppnpxZi0V0S2X3XpPoGdQndNln4AHjoBq74ckywh3q4QtayZWpWpYaVrRMADD
Cd4bo9QF8ylBBRA6AWc6FCobPw3lIpuz2M/xEFDk0odZbaQZb+CsZVUDkWqfGDvCn5Pj887+qVul
ljjRG6jtcjiMvZT3U63vW6DnaRldYeDXfMiLuEGXW2tIMUDSJzDdICSi+O3qNiVhvGHXb6Lmt+wC
UwLsDErwhiFUTwIm40Ii3ERE7Lojn4SWN2gZb+VRV3dPu1koxaM4t+shDQYpCzqcTO7oX5cP7TJc
gUZVatlCyBIT68g29s1BbWNLJJfoEb4/ix9pQzszJFYHcngIlaVInfqzhzIZF+ZJLaqkwuAePBQF
bNtpobXOiIrbahGDjoDXzyn8pVdvoqDYYSPEwcs4IIw0H8RhVTM+4EMkR2ij77NM2ji0fsAzmSUj
ruSC4YJt404/mAVwQmjYF4h/+GscdEC4PY0zl3aOxb64l8vnRHKXlx29YyWfjdtlNRCEwvofGBMt
TIlT1KB9RJLcy9oR2xscLgpEDKh0dauKFpXXR4wgH4f6Ytfs/X9Lmv6a1Zm5ZJXmRU0oHQTxRtsK
RB8tM+Qdi7F9bv6x+WhUycnWpRdv8TxLyUrGD3OoTmFnmUrjTUN8mVOhiXq1IzCjqeZ9XZZ5YlZM
jJlze+IEZawYYkbNh55+PUqgXW70HD/2Zy1ZA65bKdkWnxF/4fAfYsh65hGcHwOCNXMNn5FSqkym
CXyjiuJByGF0DElmMW2rC5Hhmxr4s1naJrZ74xHthTib01FObuf0yLW3NE4O4OhVxVzXSwlYQ3K1
Mi88s4DQwUwBhw1V+4XfJtRYlwqcjiFxq37dMHwvUWqbh5HqqdtDVrRBw59m80XhJqtFDLVFoB0S
ntxFoSqnlnp/Gl5kMGgsM+ljPQDxM6hVHvvbfzhkimZkmnWXwrWwnv8Xw5thq4HulBcJ7KM3kZcM
MbznSc71LzOmQF6vTsz06QJHyUnxE5Ew6LJsJugWVAF7fcBxLadQI/QdE9tHpOuaT5swYTiWVaA3
42o2K4qYR6dG2J1oRBP6DPJUPjXjwtfOu0wRohNE9XOtIb/J/sbmb+kjEEig7j0PwLWiPaYGjuQ2
7iVbs7jwQ+slTSuN4kO2EK3dKJ/yppVoGvKEjwzLyyjDPbFZNQ7T8kUwx6ut/fPErzmATIXTaSRG
DDffCzlTL2zhGP3ngqs4q440a9QRTMhBrByj7Dz2FVtysQawjHHJUx7TCosksQE5olVx5XCvxsW+
TkGSnug1MgQPE85pxi3hDsT+X+ITtQYz7CqI8Rcoq8SSzJTarVKfiyRU2+Smtw0wLbgCecQA3eMo
H3VtDiTq9GiSK5UUbZQ00R9d/wkvp1nogrEFHZmX8384CccKhb5JFIes3I0auhgKz6dUmNFJ+Ubc
RBuZOGrhSkUQ1asjAFsiPhS0Ry0m6rqaF23sKmnbsmWdZbvSmgoBE9Zgax8YdaIPSkaYX0MhgQU+
gwrJ2Ls5CKMn7HA24w162SKrq6ElK+Fwq/0wyV6fQIC8rlarpMRLnVXw+eS8jjI4hrq2FjMVJj66
7hmbJCQNpw7ZynChYtbMLN147Nu0E3F2Z5JWwCqn1/VYqsIMIGiI5C3LB0z+SB0Jd1FP/OUWa/mn
sGPV/1P68RixEFhJEYxmq1p1WWxiJ2lFCyYrQwrCP7ciEqiEy5rg0lFJU5DTjDcv6+kuvU+Dunbx
7jAnfOOGPna593C81sWn4JbEu33BA1q8GtmNSo/P3qeqNFzjTE3+iMmfH3IiRyJ+CdN1XAYSwIfT
cNZN2Cg/vAKMVvd7ZjLDQLwhn3EAmxV5NWoVhq9JVeiZJps/7oLGtqFU5lKaKnSwwYWYDhGVDNfh
pP50hon/sYdHjwgUx4JV6XKHcaQq7aCMWVM5xsyKSTmgzH9QMO4pQgyoNwgjV0SezSHEiWlvlta+
DGgunAXkTb3RgptNSm8Ib1arOlTmKxVhxJ/LVC/0oJ8HnGfqwBNvWiHrsrql8/ZWAbuheKvc3XsR
OhsWgPao3yYTk6+LIn653X2vekChhmY2rbRj9TUsFI2yViC09NWy2usHoTmdUQmJiNpyXtfEbIML
JVU5wmZDdrqUOLvGFTD8fyFrphMmWvHkI8U3N/oUUrcCX/vdktw7qErhKhlz//f58WFvnBYpGLlW
YYis0wHLdMnqf1rK7+PFkn6q+i4502PiNDV+yEvjlSDqvHPsyj/c971lPwo4gwVpCnnMJbG+73K/
r8wpl2WGOFzPe05HOzNRT88OCO83KsG/qrbiEUZ1iXmu3Oku3YF36oqhEielTABjSZArQFJWAGP0
aKQWwMc2s9czxlO5ps1/rTz7ZFRDjRI5YPNqpIdmdVBiYzSN7FJ4MkdQumpdH8w0xc/vQbqsz6t9
WijonBqWNA9Xs/X76XTMDIWAI2HyDkbkJgb1FrizHERqn55tvvp7FDXETkcZomKMV/ZRzP2qnm9g
7x9xUDmBUr7uN8m963LJ2QIjSEWGmMM0iJeyDRSpxPD0h6id5lUo6heeySD8a+liTsP56DFnWfrY
dCElZQ4LKkNtmQAYu/dG7/3Q8FRsO3yHlrhc7LYKeyCj4fecht32fZmfVqt0Jq0xUlZxTfC+bPjt
+j2V1l4afrWa9dfhe20V8PKOUmNsaFmMVAHduLvqSzhLe+nC6OvnYRV3sqJdijEnFxktwEyVXc3m
9w3yx6+tn//HvgahUr3Yn33+HUg3t8UhejG4Dis2PPWbcq7C81wP/EKoZpHokPq8Lu2ho4ILF7wH
aes0zmmzOG1l9qJfjrVti/g64FgYKZKciZWCIQO9AKaGHrVIU53INy5/VEBFfYuo9202LrqzhSHH
l02zslo8AZnOWz+TnAbjsQlwkMFGNwxqq/6df3rPrhrvHgHUSUJR9eczts8NlkYzsNNPedR0khAZ
nJNPkEoH79EFswZey5pDtGOaovANPKTVWjo3KysPyZ3eWmlqXtVftV+aFsfbVEydQ+4Qp7ccFAP2
Gup9HmwV3n8nEevvp41sQP61VeAGRoCro2KFX8nJC/a63uT6oFkCZwyloiWGmac4qx7vJidJb1tP
nHBh3EtZSIz/MhogLW6txlnq4NWPFOn0vHFZf5NfZTT/C/EfUcGXn/KG41+5zro+jyPiHs71Pdcp
ukBYwfFduW0aRd1jedm5wdcCd/YecShhFPpmkkJ7Vdo0VKJYrEJmLfbw+mTURTr7I5v+CTJpbnrp
lJkxqnFYYmMPOmWPz/5BxzUBfLGHRUekt7fqouxsO1iUo98obBqo6d1DHdIR7DOERM3lysscdEtO
pvqWf5FeWdccbCE20Fb5m863T4a450CRLzfHNvNLJVLpesptXPZNSYS9r2m8ayv+qIQeWbQPNJf+
5X4TYXmKya8QyhXst/0sr6CH1qazcsQxYfZO7T/3N+lGoevbmu4EgEUD86p65OA6xnOAmk4/VvYc
CBY7fFPklDsGV1PkctQuiICX8SMbsR/4BH/aY9w5dAK7G+GTQjuSGOZJ50IR7tONmxIAeSU9etxK
caXf25U7XKjcW+TN+BL0IkWR067wCcFk64Vy0xPJ6TdGaKgkDIjd/lCOujVYS0Jv3pfep2GFjkao
ywInURiLUSgjUI1q2sIemL0T2yS8+L+TuxmnKb4K2ioW5bTu3T9J1v+f2XeY5N9clgKKXUPU3kUj
f5fx0apMZdVKbL5TEmoR5jB+v2fgDSvQAmlLqZmUrsVNvEn2FcRMpy1JR/v4RRdZuBdZ3f/3R7SI
3JQrrUT73UoNa5BfQkU7WKeTEFTgULXnBT6EHiNIaN+LE8sTkIRL8QhV+S+VNhYGCZsm29bmVxeq
KJh3D2Vaze0zXIG0mRrn2KZ7ex2qU+bxjLLvZ2+nOD6TVSfUNqJZ4zsdmfrta9j3IQAE7fjWC0MP
dp95DlpG0fmO5MqiBj1zPKyL0pdJ3y5Ykdo5ydQ3g+APLIe3D2l0Gsv2UKMmDQju2hjlq1JL+89Q
OGuJqUiHybrZS9GgAn4V7+Be40H5XKiA45zQWQOAl/fO0fvlApTOmY+6FIQZLSpML4oHQiOsGfkc
ISd4GDsnQX1fW2YmnTCY2p3qy1NMBUZylVstN9GCT7p6NvrnToMqiX+Zie6wlbfNc6woL/uDzvom
vVHokM1z1ybboDVWfuITMucwjJH0RTPIVJnvBobqw3rn7FAoJuJ81lEY4A4VhxTeJwhyeYJcdkKc
L8PWXBDVr4VqS8axdsOKcsvANC/vRgZ8ypRlRc9eZKicJz7ONjbYtukd0mZ54fmKitGQ3hgW14Vk
hMw3HGMPchAtgHixD6WO0sEVzdbOhPq0rkAfTqn584QQ4Q6L5J8HEFTLDQcgDRvlrYTMNeNSy+3a
8UdCC5cuG+SDrOUOu2Jeep7UJVp6d5ew/3+MRMn8FL0nendfvcHXBq/1ui7fjeBs644eUB5N3zLB
dGOmMO4EV4S2Wh+95SOfwxODUXy8kSBpYCtidMhbWeaaGXfoHzXR5xmM2fxxiwabIfftgLiA+ixv
OxVlVYYD39YgkyB1gbQ2cyXke7rOZVx2JWcZMY/9GpmnjV5DEV1knsfntUEkggmbBHRdeNxG9Pih
J1SR99hnrMv4WSJP2V9g97L9MB1szGY3qA3IpU4tOZulDRe0j0IQUND+UogRWTwyDx1kCpIbQ+RM
1z0IbivKmdzbH0/NTpYkzrrn3RqnPxbv6RZOEIH8YHLA1DUCZ8wNQXw0AUHfKk9qKDUg7pY2Rvpf
pwLQ8zvwvWKWJ13C1VUgrqb0zHNM6Jtvv7kZrQR8a9Tf/AyURx4xG/KQFD1Y0lMY8QO8LbhPvEAB
AvDWgJHrVS2+bDZzUckGHrPLrvv8fgAHmRMXSQFxr3d8PneqH6YqJpUaiGt8tPtdD/fYxM1d3Waq
qisAG7ANu67XcQ4IgHZUVhtBfGgV9dEX+HnhfgIuQFzbrwCBn8Pw1UknlnxVOkUVIzRrNnT/QmNq
dfXR1awluMqu65FdVmV2DVolyCsGH735vfXP4Yz0hSYNz9ePMgkZYY/4X0hZdtH+IDr1LfoWiQIt
9zlIUvitZpFbjIcOWzk5jzfi5km/CZ4fvKrc5r5xHSf6Zi1H6QD1iuh12/h1Gy9WeDz1MhcWy53T
0Ypk5uHc9yxZYpuQhZxCQw1768Fj5tMcADA3u4NC8s0uFH7wifB+CPcAHnqxGtH3wpkib14z6rMr
097al8xGf8QmPXAlJFb3bzLKVO3fIqjLWIAgxTZwkEqW4ZsLV1t8C/TlHi0ynMUBRzDzMWWXZ72O
wWTb223H76nBDMbfY8TLEArKyrPJ2XmDz5f878TMvpG15xs3G4NDPGXpDPlb/PQtGVK8vXDg0V+J
7bOi0jZmDSDgrx3El9TC3yGMKYE4+i3xASqbDGwsQiWgxRcmxMExpJHu/ltxk/7TSPm02F/uueix
xTR2JpgvnWD2GvgwjoihUpsvNO9YYebrSYary8NCQmMv4vrF0az51r4gER+GHBk2RHzomTFyE6hl
qGoxxlmWudL/LsUZS8mdZddz47WmilmLrA4o4/yK2Bu3GNpOpbr75wCtnrD3K9X3MkG9+lBqzf9n
FcrQ1+mUw5eq7bwPnRbhV6Alh9bg1A4XyzCx0/kBPrvZWsN/s4EYmq5GN3AiYs+qawCI/3MxObwX
x6GEHV83y+/8MQqTgcH+LIsZb2CA4hY9FfDw74NocdmHXF8RvlCIo2H5xKiB+bT9jle3NVIQcY9h
brfZ0upLimu1JxCozFMVbXuK1HGgzcxg+WqPJRBPFPStv/tyEuJllQabHI+X+rPPLD7fFD36AlYw
B4kh7LWCRZOu8eBy8rU9rk2SMRKwtxjjYykZeaC4tB588bpyTiUrncEfkudNB5jCoW0GmXPvGU9z
HW/M04cjxmiBhEoMnmANJrgba2GlD3WFIWroFMUzRgN8H6Cl7UtGXhJ3uxIWDFAc1zRyV4dRliAx
6rbIUtZvF9MqmbYAx1fpuBAbQGZVchTQXMx0hg80KNg8upW9Y+DqebJ7OVPSP5zomMpCgxVBhmCE
rZGwm0MWPS/hPHBVxC/U5KxR8sAUbzbW5e576898Mu10eQ8wjHVwqleiZ2pmQF2DQ6OKIj4gdryM
19xf4sRWAfT03pqtIdWLltIToUfywyFZ1RBCmjwv9Esh35OAGyfQhXNTQsuCSTFpuCQYrTphq+WP
u2+vf6NsQ0mIg6uwN/uO6EQ2Wp/fblhQl2SC0+Axyw1BM0xqchrlcw7irFp35SFNZbm7WHP/mlsF
PcayQNjaHu3gu2jP433z2IGzC56Um0TCUgwMYj4VSg/HU/9g+VtdZ+BiXR7FenRKIHWuBrUCsBYD
IBmd/oKq4Og8mt9BK9I3Y66C/bDZcbznCisvEiijEsTVU33KWiEp7Jmb9KkDL1hxnNSAoUak0jeQ
uUE3Z/IKgORifrEBVYxGmzkWa5fTnpi3MK4huJzsTmSFAzlGqfPxLqwvxi+RCvMsOR2kBd/Ghsfo
T2R8VqzWy8hO4YOpDwZkHipjgn5kdxYuxKphgHrzIOHyttT7oXePgUXZNdvD0OrUS5ZESUdNdLJD
O8fBTxRGhh+Wi7vMLRC8Vl8AEPdC+dAdRj0dFE7XlS6e35IS9uIoV4ILM2S/husPC+cmB/WWrT10
mmT698P8OPCSthF/A4IzjRg16MG9ncFMCauZQ/6exa1LW7TXnkxTjEjBMLLlp3OvyZ8h9NsOVEA1
AMjIdhZtcUG8ftf7XtQbYps/Qt/m5h9RH+q+Ucidq5VFgiBG3unjDx5ShQLIv6x1vImdUkBfGmOQ
h5pO1II7ZQEz/AvXh2U/3l/mAHfrFSxuzlr4kXwVK/wrf5Ybl5S++KDVZFzFD2dNBxgkRAhT6bgE
RSnVm5Ug+sH/+8/kL1btVbuI9ZoWVbM+36FuwXeB0nKgvsgHn8eSzs5m5k8iubkKEtqxUsDo2KFG
TUQevsDekpyte9FRZ08K3HzMGmdI4/O3dQjABK7LzG+oE8PvU1sTbzXzCSHD/E+1A2SdHEoDXryU
ALU5G5yxxnTgy2wempotBQqIL0VbX7aXol8WxlTGJRZ8xcv/d03Pf7wmpWHbj4rQVGpt8OZ7V5sW
0VVwig3pAjMvRt5dZml+I3P0ugUAiKhP2MiRwpXdkSr/HPmd4ikSzddMplok/byMi91kiHvet68o
h0Ywluu2FbnCsnxW0jv30G/ESNofPs28K+Y1Heqbv7tAMoN9s8IvdWM9G3ANH2Ne+x5aAbGJ8XmI
7+6qn5lS2+MVeQwPM0vOpPEt2tldmPqtkE96Sf7q/F3pnCavhYWaTZdkyYrThK9gWquLC7k7lwqs
qB60F+qHSH4MztSjFuctLqL+RjqVzsFG+Tm/k3sqJT6sf4ydQFnBWViX1hLXLu+m1/aIyefqG+lE
+1EQUwDyVp/4POc7Pj9bfK2UhCT2/6K5gRjd32Su853q89vlT6fmLU7HHavH8lZZtxXOH5WJ8b1Z
2Ro2J4/H5iBkdn71IJb30rLhFafw5khiucoj/UycJ22W891ZcSvMkUG36DRMc4xTzzIdg39YB0ld
Ztg+i34SHcSs/leUzEFlyi7uWZjX5n3ddzap1+R8EgoqO80uo1ChHRFbuybxkOSp+HHzckF8MgnY
uSl1qp1FuStEp7v/iiMkHGlMN/v+QX2VmGQTuF4Tp0/gVAJmq7/WuVVnaXKTIOnSdJMPRKqAO1Qi
Jkyxwcx31yIUkHge2Dh8IEylOWRBXAh4qRt8oWYolcQQPq6K/YJiih7nCxer2YMJgridEBlZcJgB
r0ynFdmDA3vp4sz9BN4AWdiqhge99wHNLWjbf558dckf1akI9j7YJkDz1WWUXM54+TZrp+Ni98zq
70pvv67SXHB+bgj7fPLNoP0sNxUovUZQ7S+ZTNxhRg7rTEfWTanFt6nJfcRAgbMorCJSA4oQQ8Kz
R4OQQfMmK8iAiO+nNKgX1ouGfUosL9zppatTUwyoiH/q2U0Ak2XvzIOLyPLOhVVlEnaIFxaTCsoe
Bshx/gsz01O4s4OJQBsVTRhbQj9X7kxD8Qc5b+3CuFO4xc3aRr6qK2esex+d57Kfw9r1gbzS/wrP
MMxGvEDiEzBwM8PMnlvie3Mz4Lb+L3reeyxorABcZAAQkK1eOBevgkUPsoivH+sa+8r530labqwM
CgULuU8WFkaox4tRIY65tiovR3IXCqO3jXj+eoR1XaYt9Vt23BgWLnqGasLw6iJMx3fJX24HcH41
p5WN6Y2TDIXpv/bEOoRxBmN7Pg6GnEbJEyLlLN+H2HSGgbUR/hBFp7eQMdxt9PL6IaAChgKTsYn2
JwlPJTfRKbDQ4mWwXaMSS3sf5OXpI8ABTRFeUdbpkK3umiwMjc75dThF24NLlB4vitMXM/u0rYPV
2pWeMCw6sFel3EcLx2CndoIwF0wnhd+0dzxw53iZe5X5CC7K54XHKRH3+lEMJkpWFqxeW0M2THpI
domFHAKrPtyiX9ST9gbJU/Dm1rg+/4WkiWXR+FXEzQ0ie5rs1jM3A3BfxfdEMxU3FAl7gEj/03gQ
z5XZDaHFTLHXMfhO3tVOZ8IgtZW4ajYbGmkkeG8mr4+4XjqSGMNiNPo11v7hAbMRfs609dwvsYmY
rI9Ehlui5E5Hpf3c0RcvBfiKBGADAAZMDKHELhAo8yRV9FdeEd3oNWvDPUzAktkFnHjANI51SnwH
BW3Tr2c9j/BiNRjQG+vCABT0ZT88kbHgkb2Lv8dwBvgs24IGseapY5KEFH4h2rdfuddJeW1m0hqV
PNwRTzdynHc1JfEg/8bKTYsdwjQZsV9Q1VeY8l/MdKIePmri8xq+HDewQznAvUoKyotN8meTLktP
1YsKQBQUPqXLWE06U2QA9SO1z5ISzN+LguA0jD559THrk8FB0r9V5Tu1HUwJDMb5cNwSextIBXC1
6O9Jppr16txuMG+3gpQ20+vE9AtW5LDR3DOelXpIWqaKBOnbJ42+ck8hGwM2u2JuKZxyJC9vZAOy
o90vPAyXaGNCj9IlnFrGaIF/MHwA3VkRLAD350kWXM47ucqqMVeKRFnn/Llz+smB/6BvQ7p5tMMU
Nmr5aR47FJ4S7LYbLPYu1nKGh20dDOlh2KbPZrKz96nk746dcIxMI+PTubQpsEPLWkL/Jj2pug9H
UQliKwIbMzpc6lfaNaRp4IYkLPK15Hi1s6iuocURCcjNLEkTjqMjhVo11WTkeXOsiwaemgrm9Jj6
9TQCAo6PDvWIkrS4hIondO/e4Wz7S/diPZnl1UFef0/Qnd7igrtqkJoHTqobNHzhaMqlojPmkgdj
rwqVYhyaGXFtnbkvXc48wDmoLoDkx11HCKd8zi3erKw/bRUJfiPtDpklFR88cMlbVnmnbzk2O4Gi
7IKsT8Ci4iXAMEA/piYlVFa4yuLU6SeGcx3c62MQUU+YguiykfVx3f6WM+ZftoaL+TXhI2KxqWGH
I1kotwYWZFpyyeSjGQ4cpcCNZcLLCZx2ReIZOcA5mjExxI8PqSy6TDDn1drBOvwhKrbAtEjQjwBP
nWcWlS3jseb+ndGUJl2eAutSyulWnY9e8A1sZeZG7lklCuxzS+UBiq/vxpAjtZNhleZDFIY7bzz4
sfcTS2TFa7/UiuTCM5XAX+zCUK9oW57tQh+hwb3QgXULWSTN9Rk320r3Z9YActf2cJuo7fRLJPu3
e8njHAWHkveR1n1BGhW0B1uASqz5YNzqIzm6IlpUVb3yEGPizPzY7GEv+O1k7VOdIHvxj2PMilJl
WunKX79b+0h8tMxeDAUBIc4iig2ZkEBRpRpxaPxjOYLWespIRS0kfOg00s6CTJ5HXZE9acfF1Wn1
/uOfaCJ75MRwmMnh37Kb2ipjT6AJThZNV7W6Pdr0waF/NZxMeuB28TaiZT6Rd5YPBnxfvqaCsovq
KNfs5Nu6pgEWxnN74B1C4iGpKxD0G8z/m+vhjrEYudTK28D/Ua53h/Yg1O9Mm35nbarhmV1q/Pe6
gIf+8E/uyCNEJw6lksMHlCtyaNi0cplxTKxuPjYvuFSSSINbO8lUE9+HSkLmIyCr7aphjZoPysln
D6nWLBFkF+b3SvNT448NhseidsDYLbs/5vYx2k+UXkam02BqspV/TS2etIzUdEOb472psxpz7aDI
CwMXhGjqPNXYxkTh0Hu7ssBtu3QTd0KYGvhMjgDXW/ykKCPm/a8Az68GW/JLDZbqvaTLzKnRuHUR
gJ36jRCKJ/pxzhhrutZ9Emh7EgJYwphEN+ZxrS5hDlnNmlMassvRfWzlyZ6vrBScdVY+UF2lpmyk
vj0POg6dq6OfJMYIUBxY/o1stXDeVPc2SpGrsizkJ23EqF/E9jsGgkSqpx1J6ZNSzc7D9BZZTVEe
8lMtB5BJJTalYGA8WOicnUAhWRF/klnSBqUp1QY9zM26XWwSkZeY3GY/0jirfbty4cgTOlwCXkZ7
Rom2AILEA2YIrYEssMe0/uD3yZShQQRnImvXstqPr/jnBVVrMD1N0Xbpi/EOb6P1/Nux603G2q5E
lxdHolCB25DSwmAH4hkzzS2m4Y5r0WF0St5R2BK8gTu6OfMRlJ3ThZyte0acTa1U2+N9wJlSg/Ww
YD/A3WJOmES33ufjHc2qhxXHTR124F+fRCBW8Qarw3oVtP3d8AGTFxluqfJZ0n8uV3/DU/dNvu0Z
XxAJ1c+YXRGOwr48Ry/+Z2qd7KltVWsi+mIwXWOkhwg65hE2uXVe1x7rbW/xmUpRxBWPyWqJQkHJ
UCXnHLKL1/SjmtH/kqtKNdgVKZgOSuqV9z75NLmBMzXL4AgojumVeiLVrLox8CDprg5sx9uQU2hg
AFS+tpd6wIJDewHyXCZM5RFA3sX6XAf9Roy2re4rabCwyg4bvq6E2/admaIyFk7411U0TJwKLL8Y
che8l5rfdSu1UYNSa4Z+Zm76cTpzrm9gi56kxInwKeVdTKy+WeqVsu57q8zprGtA8npMjsEmrzRq
gsbT/AeUH7uzEMlccM4pRXvwKSUGTT3ywtVQmQtT1G8CgHRI1z1U10HahVgCDSV6THAIbW8mB7ja
kSR/XFLIuv9sY/bD5OAzCT4hzJKFUM3pc9ombbywHoJBUAjZ6BH5PArvtda1ubhuNzrjzizsxKLW
pctaUMrCbKzbUzyt4/gyaW9K0eSoEMIHPDzORidUVE5jiR0u/ObLMnBq2RvEztbwl3PcSc9vgRV5
tenpU0xDPR+fLg9RpM+dLobBjVUTcnRLOGS+yTVXLQLEal+jFaQ57LYAi6/nIRHYVQ3RUmjjoGht
nxfo999/FHmZcw7AwnkitnDgsYGbb4i6YNvHNw8rNm6dLmG8lXxM/u/q2AaFvJOC242cnU4+u+Fg
dyofdl58P5R8n8sblI4bE05EXwfxfyF6ml+l3pGdXv3RPfE3/FdN1J5jG6ygL2/GC555RmDsUink
6j8CkrfUF4evVSNoBrnhJfVKdJu1MhGHSa3VcEZLVNJprxtRQQk8Ijip68uf0CoPTG9Mhigm2ewM
obrLzhoWKxE0SIWd1mIF97i1FNoFfAKwYwYSoXgqgCUe7B3r+6rMv3/FehY5+Qoi3wheho9xr6gQ
UM2JpjY1agKQhrlz9ACNFiyafaraa+u57nOTy5r2gw206XEhLJVtBnMNC4jUkdAwNmUu0IjcH/hB
ZJNcYt142TVuy0OB+usbW/h7sU6VDOPuvablNK+8HaLDCGiBBqLbHh07XZ7uOlP1cCrR5mZYnqLg
DQwCcjep+JNd3EExUCSM7pJZhmUHY/csi5NEbbsKKw8TTP+6G1CgNa5fh4WGlYfvJPX21DWGW/LD
A217/F7xR1x0R5Q3VjCOHWmZg8bycnxkGbxmRw8t0vVT96i7DkFgcFZ7DZ6G4N+Cp7HDCRuEkEDW
+5ynA6UFCJorh7XML0HPc28Cy/WAIrJdr/6ooOn7CxjglGuX9DsGgjoSBP4zQidB2v4LUewHxDG2
db/kdD0KUyouKvjHXg2Eq97R56bJeWrzP/g2onNCCkx+VJ9xWsYVq21fQqCemZl35CVKAhJwsevR
75r10EuZkBvoXy0Dj3T8IDmPur6eqZz69RJKj0wT3oUYwTJIceGBFVOZw2aDYnN2haaE9dNsTbko
ZF8NtxygEDhtEwaPUl3fRdNiDDzXvh7cV3J2GkU/NYKCcacS6YGuRhydt8Vy3i7GbPunSgK5+IVY
OSDsspRqIYx2KwZH4evb3aGEXuY95DZn0Cx8rEFtrEBDeHbp5Zt2JBLHrC+y8LWTgic4/z+oC9E3
yEPMmu/ZcWoB6EMHbdcToXuHUULiauWBi2DZ4Wcxk28OpJKnfjL4bl9DmJryqt7wNEw8BGSYyS1p
wDScIV8f4YuJBdNryAYoVHFEFkw0O9YgBiJ+TgnV6qcmj2rldwxkZ3nn/tIlq291CgXUp0T6ayHB
t/RWarv+ACU1DwNxgZjREfxiDzh3cQXzpHUav3ZmiEdLvxAdNu5rFEOJgQ5ZtYIxE9gN4GfEa6bx
SiIHbGv3t0NaK75RqIklxVszmYPv3JfapUgsg7Vy69lxHKhOQc/RHVQUc6h/L7L7ZzYXMOSGX0B0
fVU8XeETSxCsXgVfDmDseYD20G9qH0NN9x4M1JDJPfh7Gc8foOhvWbK6xPczdW/c7CIorOM24qjI
hCyw2iD4H/ezgmvzwKwd8n29B+hh6TcJrOjELW9OE/FMVh9rphi344hzzMot6Iq/ha5kGYPaVbQ/
CG3CxA+V/SOv3ksjGV0YuCr5iDvp7HP42kiPqbZ9RFVAFaahLH8oahiPRla4LRDZ2HYCvzuR6ZSn
0FxKbIwDxbjEqv+DFU71yS/X+CCdwfoZzg0svke2ENY4i3p77EMEclVFFGsHfNQSkTR9feUaBo4v
pOKjsxGnr9QI4U+aL9/nF9U0W56IMowj/Z++pN4T+J1i3OrqdE7MucXeCb2JW+ln1HtP9bzhuM+w
ylV37n5An7NYDo3CISoS4HEq+AIz1yHbh/aiVHXtSZ8FTRljNpqfGyj1qHKRtP+2uk+yvyMxYret
Yjhb0YyylCc+/SA+62eeI17JAmOzAO5bc1pgmWThTk8BZ+UtzvyuShBqd3e9PDAdmu6laJCq28cm
9tqPDQmaQ1JareW2C8ZQRGAgpLDdLeK7Ihz7pK1i0V2Yo+mzSCLJywyvvMehYOfnRpDv4bzLykbQ
YGM+gP1KPXAACvENQo4yDnIhU03OL3dPYgU18bALj2ypHDP5o8JwjneVUhFZz/R5bMsAqjuB3ueS
qMXczSCZrspbvzKKyI+I4yjjeB1gXf1uJW1H9eEYqXwL4jZ/DkVfI7xqzRj1z13uA2Qu56gIseGH
yqEfj237i3Ia50lDmIqzCNyoXqXFavDaYYj/mr9UWrUHrxddRDg3D16Fa2t2LcV2+Oe9soo64fg9
vwUOJj7h+8GtCKeYfpz+YxLGZwdtYYrDATLarn/W0YRruAWTkMvXDDuOoOf1IpkOJ0qx2Klmju3D
2SyVkaIVBA8sKV3959kcbv2KDZGp5QTi41+M6DmHFw6uJuy7I3gIYGPxOZYrZuZAeCHCwe8nlPtv
SsrSBEK7+DAxL/2Nib92LPGbi52CtDMQq6sbIIll1WUogbbytzax/Z0Tualk3qEVb/wxRub8rCDU
Xz1FSXdz4BM+1k3HBhj/JAeHz/Q2i6neNzt2jkfqpj6WYE2a5KNwUududTPyhouvV1ET8ARljtw4
ge4QKPWkzM+5/YNf+pAnCK1cWkQbN7yxhiqgDPAoCmxr9whyWMjv8gSU/5xr+h+pxZwe90BWZ37R
BFzNW5dcEdibyv+MFOZR4p4+miEo/sp5BdxYAvk2iTtvMROP/I2j7wnpkH51PGRTVIh9k41tiJpX
DwNtkCyvivzFoY/rB4ctobfdqak5hNDV/AhZQnE0bjP0dbRu9jWF43QxKTIi8a7lP4+bIyg+I4Ql
NY4mtL/l80vNOyEPjVwgyfYVi8fYhxhNuYVs/TqK9CCw7PKvyn0YAthLTr55/VKV7eMbLiVE4ARr
ryguFdUGNicZDiQ337La0El/PL0B3/xhIaDQXgosKKYxEVhfTn8pC4rkO0dXXwgRshwrECCzsFdT
h1hDcbbxyR6rC0KF5T5AMJyp5ML9CjU9gfvssfCmPbfuGls1X2WqRkF0IsfUJ7IsPoPdrosa1aPd
u58PgRAGPsHkmwv/u648xRLkU+M1BhdVtUhk6+SZzn2UjvDoIPg7CHrGMS0dwcwrQp1xw4LuS6BE
ZMEiBo4iPvjRvBTbPabJsU8EMH1KIqBkimYHGIw5kDCtavJtH/ccySK1370QwJJpyTblNa0rhP0z
3xncm1LVFpE1CJRlggFRJEzGojU5omnfyT3PGmApnJoywCktes/DYmlGsyvOYvoyfSU0In+ao0Pf
DiukSId7sER452vCOqjWgMJaF6mgEAgH76NNNo5OYtn7R1tkLOQw338tg+Jlv6AIlj2zkDqx79KA
w4ybCKe6ltuPLXi3dlbUF7U9SyXMYC/k6nU8oh+DnZEnkQVpVn+WWHuGywP4cFN6Y1HdSKdqgvch
EV27GvsO9a3w+0KYcZfw9SUIF+cognoFt8/KObgwx/+qjGhcMU7h1WnRK3yH70Rg/Kos0YG6sYBk
o/ZuD+yxux/kBqggnkP0/3JmD65vpOdgsvDoyd+0quCy/AV7coWE4FB4HjMZWyrDzxPP1i3KofUD
wpcitbyW8NgeaJ4tS8+Ng5mC9JgMuBI/te0KPDwN3tFuqMLEK35O565eMCItBs0Mf8uvVfcoVYqJ
8tgR4iFCQiB/7BQXDd8UONQYzLSzSt15BE1qxzZQccP1wj2pN5II8tmAqe95T4KCuYEs9eyaqKQd
exWY7+92PGtTQ6g4mX4rSOuNf3Ols1m714gNBYloEBottut5jFUik5MQPXgWnWqn3ncUm0TQR2j1
0TN9SWSYp+2X41W4bYbPt9oq7TpD+txW6Ff2ghVK5XTOVdiM12ztSJ+3qsZ1dwpAjO8l93P7PjEV
5HMEA2iB+FZ679hu4AULg4tPm+faYtUoIfgtu6fO4TMRrDQgX+jFyJqjq8zdjSpX1mN++IkGN9vL
GWI6sDbJqkssn44/2IZkn3+ErARZH+Vm+uRR9VxOStLxTSDLWAr2rbuA9NjzO1/shtcbCBkMNf8m
54bWZ1EWFdH7wVp4YgUyIrS8T0FdXoRqRinLnOj2xW+WzvKYuSrS+FzFpP/D3vglTbtvFNPOUpML
1zxd1yqJ14gSFiiw8FUBJC9o9vW3J4sZZdWBUKM76ISHpduQiMWIT0AgaI2OeKrRuFHBTKjr7mYn
zUsreA65g1Wf4o78HKcJ4OmOAurFrcYWevVv0ZphBdbLY5OZuLuSReGPUT0fLFz8gDq7s+Y45gQS
aMLsy6KvpKwAZ1lAad7h3X+S2Wkg5FTBYbHyQk5p8KpaaBNFn6UL2M4qU2i1WM1veg7K/26rmYt5
rVeEvgd8ByhdDc6K+AEIkRtEs1NttuP2yPHE2soYRVx7SPsAWsSoqT2kUfgEnSaODx2wYcKOqnBS
dXzht1JuQiX7Cbj2rkvM+SAALvcCZSErTgO35ZKPGrzrNUYee+6bobSM+2wMOSFfdpf2ugtVIT3f
PYY77DPswfi4bTh6MawI6oEvOxj7KxEkmyc6r+0aTZw4+PaZ71u5xm0btwgqgVcP4EHID8ILnCa9
ULJktIvd6nbJoYBVsBFYvj8Ir2xdFL6L+6ekmlgHOebzNBOIvUQ5G6EId6SmZsEVS2lWCIppxsO4
di7eAwiBxnzD6a/PC9KbefiqSWCXGN2hO2RY6URv7E13g3cILsiEJvQK7KofsI76tyU+a5yWXTJa
z89UcFjnch12K4qijGKFZ3Hq+omkmTNcn4rSMmjvemktXPdxCgEquCcJ1HvxZmPjAM9M3Bku2ZY0
RvOtglqTUel+NrvlQPGIuc61gbxiBxDBEETeGKaU8BOooF6XWrBdaghe7rzl4rZGUa+XG9HTIjCA
/uPTd4XFQu7+GTgDvUfMEZhejM+7SrhRiGZ3iqINoCqMEiDZSL/DXtewZbs08VxUxHjAUKVIavLz
DrYLQzYVkrvgr6RAkLYfTbk9OUEAo6PYShJi1dq85YVGK5EcH+p/TloSlkaj4cuGbjLuVVyL7uLA
OiGcEwyrr82wCU0uhSJLQ9XgM4JnLjqoW1BrUhFUEiABRMxoYE20okhRktrZOt7YESbPFGW013pU
vk/VRCAvq38UI1PcQJrGqODVL/atRz3GdEVKsup03H545vAXkOTRhKYcmF9eJG0MblbbAD9B3Mjt
mxr9Exm70X9/vx3ht3OH5KafnK1Nb1ZaBdwskK/cGH9Jtgsr8uGDaew9WKca9gGXlMdSl4F6ILi0
khMbzuEYRg6h57AsumgsJsYeml/22+3yOBor1FMXQaItpy16YHl2AQPnMxcpODGJhGgfaM4KQI93
oYPsoW39zxRFo9+/op5pD+mlKnJYQImi4cS3xOdsI9ftvqD80E39RllzkXpkwCLdVE4/8/lWBnOA
1sgyHgWvXINkOVXyb8kEF1dMSvdB9nOxHbipSzlNs97jXddveh0ZYYfdr/MD7Fk/nlGWD7cq8xMD
hI8XOmZ0yq7aOLEv0QN/Ayn+IYyp99uBi8ivZz8U8O/HPtKlZaORX8rkkbAIFQei9zIAwPp7udV2
wYMXEx9O+mUDWpmZXn0EdZR2eRIxMRb5pX9NxR8jQKQrGbpzgE1pj78MzPEl86azj+2xifNfHjj2
cHOq60cZK259CNrp9SBsHzpGJmY3EWsRufOKpZXBTTHn9eYnFg6lHDW1N9X6fXB+O5VdEJdQq+dU
VXYyJbwMY9cAsW5oy/EI3LULDPhb1nt81uaSu59WETZTklprPULzZHfDBknIB6GDI/CKpTY2tpoH
Ru3Nn8i4ix02TFBpwiE/Sw3dQjKMMwsDetjoxfgvvJysPwB1fEdfVARGRtSvlckDwMCNjghPEssW
GnNmpSlU4Li3Pf6XvLQaXAFTo+ljob5OX9E16qfKDwRcX9Nf9Ii2kecH5AlrRVlYpUk7ZoGQSbpL
mmpss6jIuiBuPXOpyt9iM6BgrBBZfqW/Quaa+2epLjG1zAl/ox9eLYRz3F8X6CNk5UOwRCMcT21C
TM1WRTodLMdGXMljDfM++tH94wotEXpeyy7ZwPsfSqXrGisKHei3YnOs4qUAtKbLfF/SzgptEyZ7
/Yd6QOeQ3b5Q9JQ/e3NgVcxVij7F1H4+RTpLHmV245GUcgauwUucuaIbwkpaBeh72H6GvdKKMECg
0Sw8MLM1uSDbJ2x2FNUoou0iGbIr0fjz1sFs0R/YQdWKLXiDDPVnD5hWrDIlsoTz0QKkOEm71Jrz
77O4w8FwgqDi/J53AFiOPF3WDL25Fh8MVu/5CiPIavtTuM6YP4Dx9QSMzzsYX54fS/Oyom0jFs6N
lSt2ZEn7E5XYB9vHOuWvU/uuEW+0J/lmC3PCyWGymDikVg38VeXGT0cDEiztkUsXJZouuW6SlB+H
Z2CCf3mYThaJXt0IFg477xtKYEzR5dxEWBZVYneP6kiFwODChNXWfDI1CgKvQxeYHv48xz9morvw
YNIfpr6BIuUTiCoo9UCZaU7wJVRdzo8eHW7pH77fIcGKmBpt1kZ/nb7P9RVvvqzclwieyX+voAVf
P+zNhp1MrVN3sfUn5BD80nkF3TqQKND9Z5+XyqgB039PWJWSNKxbdDr99YG8ZEdsXylD4KqREzrj
et6z3gFXZcU3CydHyT75cOjI/w7b0OOjbhFWXLwoNi8SfjZH0OIiEEj0H2PvJDaEj+t9KgDXAhVW
sSQIGkb5B2SssOMNc1aRP33kNnbm7xUvYYGTn0AojfGndGYBSufQ/yA+uBYN9o+BaTsUUs6UkDjP
xNGcsRS0eqJ4v+/4bv6z49okUeyFPGAQz3Y+4djcXreb7NrcI9551wJ3B3oWqtDW82TCDkgsXleH
GWMvO1uehuIpm/0z3E8r/xEAk7G2wVn6Gq3FH9tdA/pRJSWr7ku82oZhV5zIL1yaIaGPq+gYomDE
1u+D+bNFMm+Nc0YuaDp86eks8/jcCAS/s03O5DyNtJpWiFOc069lMaTfnyP+ASuW/S80g1qNH+zv
b/T2hff6Rc/h6673iLDgVnFM1UonA7YU/JS3AcdDGR50SWn6FcNkQWeH6sQD09u7vMZWZzPhimYW
IoinR35h1mw1X1BLIt+RnMMMqYrdpE5XOXdVTbr6LO2gsdBCrxInFzclbzGDONbTgaytm+sP+88j
RiLqvEUPL5MRgEEQ7WuswEjl9Uc4q3kNO8S3SbqG54gwcLQxwqr2kSezQQZEmeK46O2WkrsSs8eE
nT9yK5xWAawLCqUwHdSs5T0R/rYqro6hdiYL121OhmaYdR/hh91r+yZDWNPFtUP9GjDwvO44MgZT
fDg5Lk1iZaHOS2W4Vpqjek9yG+NLzYWOBFukTCaZ9MkON5+Sb1m+2TJy1rHs/64nIPL8W27wPPnl
KNYEWTFG8qap2IlaMaDoimqIf8VFnQHRlDrOmgu5k5n+wZKE28k7zE0TP0bw9g4MISbVWCrTiXAb
cPsWVZOH3hiKScGMIind45pUNoSpr2A7JA2gOjA2wYzwpGKtw+YuUbOMdK4f3t3IU4gJelDUDkaj
JQ7dfhaiW6K/TjUO1mbqHChbH3/1Vc3Acg3IsbceY4wdyHqJ7MdFX1R2xxg2DQ63R1NSXWg2nduJ
VU4LbxTrU4iwMV4FuHpTKh3FFY3NTLaeKjVpzATEwCaNc/V4mpTc6OZu4G8VwIzYLSPXjAY6m8q6
2lbbiOvR+nVIuLKa9/A8EdqTxd/exKsUMfmg2pkXLva1fnt4I9wUruDr4NVkRJbwTpFaR+ngZC0t
clfegnSGPYUtWHPFND0EK4H+onpH4Ob5YaqH5tNkQ5fc3HUmgkmZAHQpQlUXonFz8zk3ObppuoCw
qZf7CzI/Ny/Pw8EWEUgjZjAY17qed/46+Oi6W4VrYOnfjP4ZxOTP2/IZZMxSRzfRBCGFNzf88daS
F4CKH0EM4QGlg8Pd/bcLmmdaLsjm4wW3jOrUpSmw4Xuz99IFb+tqZu8cwEiIFQD9KdbMX3gIoZWM
vq/wndt52Zb6cSlWagkgtyz1reNTvVictxn6uINLxDbdP34Wi2hgpF8Mt2BI/AjGE/teX75Fjs8x
hF3vk5Xu9nxWOr03wwbrG1wbZXRdctyMvjbqp+yujznfmyba2KseXAqqEnuUukvRi0KoWcnbG9F+
GzSPK0UVsQZ4IWyhFztQPK7e3nE1RWXRW2CO66ckRaDu+7TqlrSU6VuQ7xlKcwyYtW6c5OYRL0B6
Sph/jqv9Yjbrs1k48g1R2dn/2Rgy4Z8BGrLUHUIFOhEEW8sg+qES5X+7QQkklkd0d9LI+4lWuZmD
gBZenf8Hsit4XR0s43CtZuhdW6ZkXM38pvexqAC6n5eHJ0rmwnffTlUFEJnwlTWsIifZ4YDurufs
hPTFMo6eHeBehAFBVbYxoKSSsQfo8lavlLQ3X81hA2HAz1+43Drn3ccBMRicwFkPYzL4N5lZ0NYg
ZG80fo6n5h/+BR9II9eMCMdqMkHjId+83O4pE1RVjOhmvGYuYvwllW415bj2WsP+3r3eNecOKGgN
HAcJxxmAqp5a/cLGsTj8Go7lqpffMnb4eMEz5FwrKnVeJyIjOhfYd09ZdmmMXY6dzLvOUFxkiTbE
dHOrik1fT13v2qyTFrig7/3ON1GSoH8sZDZvgqBfVh5Dlzq6xCrkNkpBJdb0Hndbyw5ShS3AwsPC
I/5MZNMexWLLV3FisUZiydNqg4+bQfh+RdFhwYoe/OBzseNjB4Pq9spOzARHqJjY71hBVrTr3S+D
isYQxdvQyYZkQIdDDrNppT9LM6skRSfp5MmCFPtYo2zP3AR8KpPYL0OlPGU7g95pMpS/gh91LWNJ
5dX9qCQXaeEuGBDzTJH8TNg/+AFmU5MhDY/+UYbG9IRTapw3uI75ypKuusiKXfwcH5odcQjF18vo
YAnlYySwrZOmtWG2HIaBpHfDfukDBnmuIR+w89Srl1QeWB8gkeeWC6IWT0uD6IU2RnH10N6WGfqd
lyXOdAhVtUSFTcDepXpbeCFIkUD4X8P2MGID7Z9uY+drbBoNiHixdTPFtKSRqOkN895zMSzuFKTR
np2ItOTFNLIThgUh/3RT6MXlforggl24a9nyK1NAh+Ft6hGABBdbfHC+/gUu0aMFxUE2u7HV7d+O
yyAkAu5LOV76/0cMCIk45/TN1pQEVx/UWXHZOw2Yoav48SlCLa4DZb06pX4XWSa/KXWPlccZKNZA
i/PlpLsh5nlSCiiJuMiiHrBIU0o2uF6ocV5ph0ogBZCA8Mqx2ZkYM/r3X8u50/FqNIB7gMKELFN1
ni++F3UDDetArUMK+kBRht2ZdFKhsf5wPxMiLRchI2zQPhMc8Z+K6o+zFs9HyoARp6yB77S9Yc2k
21mNaptYNtufrijr6WbAdhN3lzIVwFOR6pxDpt7wZPKpzs230q6xD8T5V2UMm1Wxu26blzV/AtjJ
zpdco5RBN58vKFF4GTw7qGOl/2J6v0EitqTZSjqPgCGw3TErJU0UQ7tpg7TZTHS8FoqI28ic8GSp
7JUWCnKY9Vzd4eNFXoPKTPbaBDpI6nUBOlae6O7SoMGTUSWu4XSvS1cNbHCZWEv9+EdP36m/dFB8
StcTiB2W1oiGTCHLHcUzTQvpv7ErCIBrYIbdb9CtMQL14iMw/axrHYvMkkYaBQyCRuqaTEALV/QC
hEbaYMwi4BQXVdP0kLMaUELvE5C6P1vxX3VEB9xGFKhIAJ3T5RbWPUBWneYsccCrGlerl3U9CoXI
VPX/6m7D/KK7n40d0/RXwdih1Otb20JkzWl1IvcgQCxQySSjzf4POM8YnLPwck2HGWcN9lPOU1on
A4cWetcykjpwrrqLY1K6bnu7jG3P2CeV3VsoKjUquRwiJMjpOnEb5NeS1onH9s//t0oozDRmgp78
46+6scNhNtins5L5DP5x29ztTa3EB8S5j8cMF7Zkc6C7uZ8XvH6uKQ/eZo9qUwqZc0oMVMMzgCD8
eV1v9BFybwj7c9y4FgG6Vvdek9UOP0ChJNMaUuyGWSoMJfZ7NSnHKDKGHvN0Dk5w9vXqYgrfVSFy
RVetkD372oq5yZZ0fF/t/o1xgoDLi6aEWgR9nMCN7PevjDZA2k8+ReDJplaL72lR5O94d5OYtXAw
vQCJFRiq+WDCOPfMC08imBn+1+lD0jDOsUtWPnN6ZtzU3AkSUusnRttPz+V7q4NGRg4sRm7e6GdU
X9zbh38xYMEIx5f9WoxThZLuQmLBlC2OQTKH1MW/pQhVQf+7AO3GNj61JJ/WZ8bz3Otw4wQVBlEX
u2ShNlX+5hExpl6IOChI/8RGcmVdEx0JBzFKG44nE8BmK44wC6X0SqqX4Vr3f3lRcfYDFcrTHT/j
EMXffktzpgLO5bPC3gqwLlVTpJtyI3vSzOaurfZACVAxtZP4mXPTiTr+aDExJS1VbxS68ivjD8Gl
gXWWn+LgAYpd+4xBI/8BiACp6onGqwpynpOJ2y3wVEGNLplY9l34A03+T5JcJBr4Pt3i4wKNYq5Q
ZX+YwvI6BuQTn7a/7qJZUux+KSLRLlDdxsZ+dFTe2TnT/xiY6OwrquNFhelBIgdxiPv0hywoxMhg
FjawWt2KIs/ml6vYLu288fyzUUKSMJSKOyzGs4uLCWTWlSfscpfr72UzwLeis5NED4RZRVCrx1HP
FDYGLA63lVVw8ZX5UT/gpQDs6riMbmeUJAYujSZGnOlWhFZAaaMIPGWOTDamQa8mJNcmnOBkTDU+
lb8X/NH2mV0//dNn1+3aPbSZCT5juoG9cmW2NNXlEoT/djxxxMc3c6vdlO+iPwvZRwUzXM8tV7I1
s+RCXN/yhDLLzDINunx7/G6TzgyUeswMX388bgy7WPC53D4u7qO4Snr4tXe0mgPfX+5LFkJ55H+l
SwqrPUb4301yGq04v+ouFVNS7ZnrfcxYbp7SKG8yTjsgfobWCjL49CR9+8dVU2MrTCwuaaZsvrvq
GLEy5abG4jfZY4gv/87Gv6KmPrKZItBGj2uqvA7SI6MTX64U2SqROH5mywAQt2WhMAScdM0/diIO
DUHufZ7C2LYtWxO9LEUMNFRQbjcQ4RVaWntN8rrVhAgDn6aY7E81/qXcVgsbpGQ42m8H918hXzrf
LsweQ++/S9ISfvn6r6t/12ztMDYYLG+QAZ8toPNA6Ohde0qM6v/RUjIISNvjystZc2NqtFRW/ITk
wXhFXHL1EZ6EbTTy7m8jowxKlzhd9FLReBbGht3lY+mv50tvU3Y1rljkjIMqsmlq1Dy3zb3AhxMP
PQyzpEbf0zo66QCc+mC7JEZyl6n4bk4YB+sKwfIVbufd7c5IUB+Z0Yp/5I0TvQLLmOBVCvfx200D
AMuOnGTJmRNvN8JYsTsUQVc2DdvtqDWsOCjWXGhHTQoz0rjLjvmIudj8IZ+6Nrq7NCTcoRNhTq9M
cOzyqoiINffUaqfKsqPu54mf3vHAestbGX/f3U8kVwdyaqjIGIgWfW8lOHyiFClSY3dAJvX1kgL0
7bMNMKkr3PaOfr4ab+EuBuEcygNgTTwCHrtPvJ884axZsvC3Y6RIlIr0oKEJtebz4ROh8RZp96gD
DY7Po4AN2qLyL3l/7sT6TmXsovgBzY0kZcyD7b0MnO7KObkrFQDmeXpV9d1p4rMPLo2Gh+AC0rPo
8mJwZoL8wGO6L3eKWgC9kQh2sAZ5DBwDLH9CRZkdxgub9nK0NFZgTVOGtP93Ky6jjM1mYATI6Xyg
tb9zDCcU83cG4oB41EMQzwa8szsACpgUGJPFyK229om2CBhnAA16FyqBDBxKgM1V4N9gGERe6WYb
x/NL4ACd5kl+nzQ677tlC67WdnxbDjuRXjl0T/+Lp9VFqYF/u2QMJlbkSHj5FSm0c8D8s4Q/p7us
NEkhpyhZ/ZU2Lytkou3QdoaliRb/dFoV8MxQ+++sB0vJrQHMWDb+OdSWpvwFD8I0AeW/OY2PjQS7
95mK9DtRQvzHswZxwvJtzWl9+STlXG6cJKQ4aQi/+1YR0on9Vq20w10rlRZuHs9+8boz4ZryV5Ji
kHjhouLH+fOkm51hRFeV9uyfkN5ElM8FAYl+5xqsNa/IAQtxsCiNNK3Q7zHtKzBl8a+r/peV+4e3
l12o30gQEvkRJ9dESzSQM9lEW8JvxnwmYDaj3Pub/DqZRLtp4GC0KYDrSuugoZxBktQcMJg7B1W0
ulmo3XGDuK5QP4dQwOMMA1hvKQdBHTKm8oxYFu0n+j4giWAWtGx/ED1h2jyewUYktKQzFsiiwHYC
4pInvsUX9a03hZSzm9k+BCUoxoBDgPWtelG3nK8KlpZPYL6oH1Z8q1v4eo2FEOfp9sAqD46e32PG
O5JvEemFOYdkBhcs2nI3GJBYrneitz6XzlQJSDLm97fgDANSlZl4r2GpAwSFw8slxpqlEvodawwt
9GB5MqJnDPUWCW6kFxIBJzXWIsReIWYaehBYiqCutRydfW4GwZQlg2rNM9ZA5wHwphTUT0exbZ7D
tECWuLu5NcSKaD9SsNStZuHbYvrBzCRWooPS8RYanS9s4Rc9/C5KiKBQGT+j6F36ZTI7qX6EqYfD
+RCQ+nmVDDhBfT8qVIpYBsvtbFSGDFNc9zMUceYfw/2VqDrmy5/dKVMzGdDGgMghtmpCIoozCeZq
bL77uZuhcwa11SGRQB4D2d3MoaUP1QRs/F6lO0L1Q8yOC6+t6yjLj5DkRmk8pzOFg+64MNmfY8mG
FOqWLDHTSIy4K9Z/ES1MxJ1eTfwOOC+z9G49GszoBtUxYHqaT2sOCsF+0/cwsAUO+nOMfq3BSYqt
RCWzthI4VDnz07GntFMuo4Nij3hi+8mhFq4rgNTpwnJriGjL3lS0tpukbIzgEqJjGgZkulmaYoSS
MAFJMrh6haCYVOos/BRZR0oUj9S382DS+4300/+Fsq91obS1IP89i+nCaTxqmcMHG6lmFJ7vTM5h
1PFLtaLvISvaU3uvyzWCdzOb1TIuJ+ASE/1vZQo3IsrOQB0ulqCWkfbzNqlRQtVI3U6rMyoT8rpq
0OL0zeILEfxMeKuYOfC47ksMgNj1m1nKjcI0C9w9kZgyqJ3TjiP95R0jJRuhucKewZf9sHVHIvEo
/qnNdWPd0f8if+feQrHdp2wfnPKSmr5kEnbQRrVuxmAvygtbY/lA+cc3JIGRkYBiHVw2mLCCs56B
NdEVs3oT9RWAhcIAcCU/knWypjgdC7eav1AStHpCEYk76UNav0QiUCONvoy0M/BCVqbzTHUztB25
741AADAUQ4ukuDq6l+gTZsRxsaD1QHQeCLo/uZaXjqPQxten/d6P++kKYvwrtJZUbYxEZNT+SN9B
9KlIjvYWNpzHNiZssOgl40vFdnElW5cN2vUytmepXOj/gRAlgQy4srIXcECSbzktmH6q9XUQyjHO
4rhftAYEz2aDifw4tm5qqoTu3cxGFZyqKZiJL9elulEMzaVRthj6fJYOJpEylsSy3hyR6/FWF7Qv
ih0q8h7EedXOdzPuxjhSIqGoPFyCX2yyGBEOFmmJ/ILLOpeVcrwUD9pBe9K6mwBGObfslkAf9NEP
4F0j2zM9bxj8XUGSri/Q3/Vg8Bb8TCfHmKrTYq1+2lUGjrCxi72WNJN/xXErdGxIyVrgDByAr0nP
gnpPmOte7517h/WaiFEqaq2YJ0dgoAmJ2YugTd6cDSUrjUImQPYPuAjLzkNMyzrQTIFYFGEZHyhx
UhsoL4AMpLRqFkVc2MgjoLcWayNnMLEy9Cw5FFgUBctlxiNa/Vo0ujPX8OUi7MH4ofCwLj37xD1G
5Fk9NGpziLs69z7SNnYbnnNuPjcPT1XIEhSUbmPowXiuxoEVEg91RHBj+DNPLxeKDDNQTqZg+yde
C0zms6zXG6ygNxhGqnxpqs0PJY5HItNN2I8M4z4pSoFbY6LAdpp7SQd+g2QfI/cuTbN31dU2T9Yr
KUQi1qhmeto8hgOtQ7RHGNzVz3kMVu4uH6v4yGyFQIEy4ke8ihwokCbAtd14ZUUtvM5+X8MTLaIS
P9l0zpK9zlKZo/LX3W/r/n63ZXUPOm5JdRUenk1kgMIqXbaJiezHJYzOhlJQQUwuhPNUShilxNe6
YG9YK5KKU9uHuqbcIUgACVqaK/HVh8D/q131TCyJrnk8tOHv/oHTAvRxYSi68NM3OrQvkBnd6MS0
jqhl7XAM/gfLPyiYKeAmCAHDToe5m4KlfyXEXlDlEJP/8UV9r15ncKhzO1G9SVDKWVEyJQn5Jq2q
gErxhVkEGp8RiB8hiccvUDGu+rYBDOTdXwNETuYCh0zh7qzP8RA2U1uJkqkvgI7jh5+7EbdDXn6P
W6LqycZg0NxYaICiDJPI4VNzadRWoDgULQCMVITv95i6Cn6uGrTVKn7yTRzqQCEZmBivWIWB1+ws
k3CKS7L6JilKMJh7mVGd0jKEwvjQ3Z+upgCI6wLy0pXWQRWzf4TRRcKqvI4Q5v9VzMATLHKf2UDD
+fbMEGIkkU1YMs3mQz+ztIJLtdZKgLX4bK1IwlQqVeJxjoyZzqOO94EnR5NCejUfipK+owmV6Ubw
TMLZhlk3lhOxXKNF8m6cH/M4Poor1NTEI8V44HBTr9YaX9uEnNIqNvLBZqXxFGOhfFY7C4byEhXl
oEMoTVlTRNdk85GFMloXLy6LPZUXAy2gpQ8C50wfJ8OYDac6tv9QUjSPAiSQjQqw9g90W72YtjEX
R4bXts3m/q4Ex6ule0ym2yBOxIAinAXc8eHw7YEaMU3/evdmKhj1iPGU7bCFXzLSLIdqzHPyQpp5
or9B9YAxb+dx4EFbeamuHPHhIPCzxg0n7bRVKRG+Ih0BZDLaRx+vTVAx/RBju2eTDNa3rnxl9AKw
v8bDJKpGoplb+8lbTu+IGvgrp4+f3vNdz1KoFGSq8aqLG4MCFxKFm6lX+armpBJA5f5mAMB4UEUo
JCYTRupkgPoJP/lHaU3e2z6DykLRT3wDvIYBkeqJp6DDyeELf3qCV09wZeHG8/pDdJgyBf5XkKjX
SLaMKzw0KpbyP2mzubX2Rw7vjR7k15C55akfnKgwNsRBSMxuc4j6igqZIbqtB06nDrbHzuwnpMmn
mRJ3PQNcVefRNn+dFXCtdLFvcKYHfUqwNaFmzy8MD1rmhskI9YuXAbf7NramLDZgkhseURmNYDy/
Ca+YDjGhxjMxBg7Nh1+8w/pm4RsZ8SWCdA7CfrGs5E4fCKoTSVH98uNDw0cehUetU2NwgIekR10d
p30kxYvFpEziFYbHHD4GXB4GCxrX8JJ009LbjwpLPalDe2W/hZF12wR1iSpPjlFXKQKa4AXZ3uO6
/UFR+lKfnA3sjgZOQ7VCvBViKoYmcaWfzbWtEAoVx8C5f+MZRkI6uSqEQ6Xz8tzKe/W5eI5p4Wu9
LNqdCM/8IjH/7InBLbxsw0Mo1X5HzNXFGLuMAdDIP8GGYzZaR+ZiIz2StxvK6yQuMzwc+d4q91BX
KCn9c0M/coiNbbkH6PWMjZzXQo2McosKazzvtUpaHudCXNEiDxG1KOhD3UF83E48M9JyCF+8lQW5
JWxbW3wXTlgQbBwAsKQRff9N/pCdYYOHNxYfB5TyoPI1HupnoRcrByaSz1aWqHEv1nZ+yq1aQmmD
oGX2dd+NgHCg2X9S16LRJ/Rey8gDx2jPA+wdlGEfybSwDdkOXNOtaSxBc5glo23sehjjTuQO13h4
+9eOZSLO78AZ7pJOY++hcanEfYjGF+hblr50NodJmzaSZi+nS+FzNL3xq+4llP04jF/e5jF04crq
P6QZwVpJ9QTm/MhKT7zd1zxhrJdG0AFl8XEJxjqZP9y03qGnsSZyBXHRndAR3NTQsIoW4CenHLYE
uyM5+UOSs9EbcQPqcyVhDNjiFs+W2ZJsXani/gGxwikjAWmYzihBHwXo4IDNttNhuS/x/enFIBoB
7Y8z8pW0M1+4NS8nhYH7Tt2RXDte5GH7BgdjJ7jzF0QHXr7fznWI5cD9mST1mjcc+4UR//vDaUNG
ceKkTLLRrW+EgQU1o3dHcTHR8HF7em+Mx2xukS3bSFgfm7KQopdfZEbvMzNgSuhy7rk4wbjWarIM
qJ8k9D16ZTeHBai4b119KE+sHIvR1p4ajYQ1OWtogn0o+xWfDKeHQqgjrPOruV1eA1gx7QLUllXD
mtFTMDthYSTZbIklkr9YORA1VyPHvw/d//enzMdXOx5qX/8YattYkmCvJ1iCw6y1HEq0hiLJhRb1
3S2p7tkZqG88YzYrcsQ507On8tBL4FkoOQ3e17pwdyjm+AL8G5Y8cJF9aTVPSH4CFvA5Fbvv0qUO
oDUh/wFj3jDDiWc1KNhxyBz6sVLZPhsc/SzudGZVASJu7jCTlBYeiS6e/LIgzGXSsqamvjq6wi3Q
T+MedudwKlIgxqzdq4eAXj/wHTev26iFWxMjA4TXtamf6+hXb7K1VpsXXYIZaJuiWBoTu435nwGJ
/FlF39Z4W8VnMLyiQj6OUuEqeFxOiLxqtg47cF+ok19rUy6TSerLlV0skk2OI8pD1aBQa4+HYnVP
YxWCyL/G4pW4mMbhiRadDrA8q+5+PGoVHQnhRZCLVpz3Wd7ClH2Tddl1dJtqVI1ge1KMz4VUev+o
5tMiANJVXp6AuIHnmpy+HGp1RXNsnbcKqXhE8/6qapv6qBabKHkrguf6RQNI9OldHKbaDq0cqBaA
2s66O3CGdnwYDhEGR5nour3wDJcPlMqwIBRnhKjXFGErvGOWhg/COrvs3QtA+MlLFyh3XXyM6rly
c2nLjVH7QJHWBRSIfQnL5HPnnh6GN0JHV2IHg/c2HNHOtMig5SPsuaGVoPMSgOIB7mBE+43k6Cff
wP7fveJEDVH7GfyMwsqdaOp/dEYpKjCtJFxTdLiqeTZQe46M/LJ/tgu3FPQElKKvbkA8s051v6BC
UT1vodwWLtt98umdpSmxxySnap7/d4/tzM1ub4KNxL18LRuj8QukpLdSi8U6wDJrmw+oDgRJczV9
VRnJLnY8hdWvObqalaFVpbXouJ2x4WewdIw2M6WUQZ0UO1nr0MtfsuTdQn09BnsuZxw8NWYW52w0
g/BdsG4o/HlqWnXTd8QFagxqOk1VM8cMK7ErkRqA6Eq5QSNFvaVorDJkaYf8wzune4mHYr9KTl4t
chFg4mB0fSd08kMeuSfVAdwSevWUd3tfktUST9mP1OXugJUof9T3PF7mzOsTxVWdX+tOO4nSgUvd
k0iHE8VuqhxtTDRSZFuBiSp2ozcNrDMrgMM+seQulSAsmfDIHQVVYxQKEbjJXFWGSpT5cZgBnYNN
k1DYASPTyCYVkQ6KI/qmnDzeOrrz/mgUXjAeszVvMOvDU8qQJKV97eTkpLaamZRRyX98W6y1kl7m
WAbBPPU7vMqoOslZqAocNVxzD9ENRwCd5qv5eRhuufcEW0BjXllAsqqqS7fiuiIBPnQ0F7aMhiF4
DLkYtNOKCucSn0aKxlQfgTNcjYsacCtnQvUSqEovNJvz0MrAEqkbNE7ei0UfF3oDGvKJb3FwZ/GG
MzUcJgoA/FZ3TnXugKKO0tArpi8IjyWp+jZT265Ymvw5geISBvJPWMpg/QpdUv31mcZLHGJHhi3t
BD7sR/HWMjDJzc93hGmTu3NpRb9wJ84cEZgu81TjmC0o2dqbzu/3JHNMGg8/5Hhb96hwxCYCakSC
0Rg54Bs1LHTO7eT6xzIJ6TMVNTPwQfHpSzZEBqtJysqSWMHLkrzFRHgPOT+iVZfEGb1K3QuZB2nC
jVk5ik6qoEaIE9fEMWfW9E9AjL1Ri2HPWh/5j88TiGaWqmA3Tc/qQFSiZ8HJcqUEpE5qDIWHQpDH
WQ7vsn5+X6SoihfQvMypIEwHd6WuktgwD9WjhzAh5WpNhvntK7yK2dOJT2JcO0rbeMIc0N4H+uCD
H5I7R9PQMbwzh7sQKvZw0MhmLtDsl3jiSnACP48iOjLczKxB6phwLMEa9PeySyb8aWkMm2E5hfME
J/bbROMt41gxeyaN2YvepW/cdvvh7V2je/ZSCxwWwn/RQz6mmCb5yF5Dv9NzlV3jfHyMNr1ANE7I
HKHu7q3V1lqgPBWkbDs9JZOS7E0qqPanDjATJLXAMZmgXhbKD0kaRWoDTmkNU7bkazd+Yd65CAWc
npDTvbYkoeOD3TVRdlZFaiubZCnEVBUktnFBbd/iu0CN10ixz6MWMdeALv+15KZPfeODzdelfbq0
eliAvcwwmv3q7r3ORPPlrhtS4O5vBX58jFGgLSyhflUq7SIW+p1FjsIB1aKxii0fLxLB29ZtVCGk
Ea9yHBBbM3ubPo2K95RwwNTZcZgO+jIIMaIuUmPgubu42Ula7Lh3ijggki3A0xWSSGDJUbzDjNSf
3E7OKyqhsugljv+uujCjUNYTy+0TzgD7612Kcd+t4jPfPBFdVnep3Twgzkk7wxdCJXC3IWrVpYeU
5P0Y/hQE/Xq0b9EcVw70idxD/jxcF39e8neWGGZ2IEzdbawjUr3pQccjOjryyhl06Z+TySyM01C+
jSo6R2HlkgdkPZhB4oGfKu0PK7WStq6Q2kMuP5m+UcqSIFusmmoETekfd/HasIYnhiicbQjnzufR
BfgZ5TimCCuh+Y9rN1fMu/gwUJ6yxVBy8N/7qwrdar3Jzd+YJOJ46lFI1eD9opNdlt/KZ6Pdp/Qc
f4ZX9dJXnewZyw08zDEgY+GF9zsQgJW1684sWxriOqdNM3YPqcSw62GfVxtQ8hOzaP4zJU7AdlT8
i9hSgtuibV48mFKSUb7Uc6UklWXhu+tzZNcim7sLek/QyrFJqN7rq2i2Ff0SCwkGuQCn80YZJ/IZ
TJ8jw6MuWeI+w7LEV3fvn2MaKJ/82cnzdSGMec4JVZHaKNbSECn+l8NpB7nbfNsT6g5kZKqMXYv6
zZoPzhOnZ/xoOE5JEsHz8lIhDNP+NaEwZrpwU1aHQq6SbvOjXYtSwqxPpjoZT0JPL9jvd5nJBcrn
yFFO8fwXmjDeFok4ERY8CLcQSSwzHpDg1mxfmSwXRAoE72pwBZ/r3oXyiSigSUqrUuzrrvX6T/g2
fenqCDlk1zIzOxlEeH02zflorMEb5YC9Ti/qIqwpaBERJtd43cQaWhtIRhcry+orPYbzt3q0Pi0S
erHivSy5NjJdJNQ7YNuiX1MMlTLeSLBUTytKo8nFrz4ow2eN1ElOIF6+QitzHV0XHeBeLEPARkvn
Jy2YFxcxg45Y1Hv6bbsnDxmSHIVqLULu5M+Rjg72Ja9IYhrHQ9/JqyqQIvKrBsoshqjf62KfN5y9
8MFplNTPfDUkiLN6QZ0UBZKRrtq/ydjgHIWEPownaleyu7oqoFUaPWxxfk+VXBccUp4dACm58fOR
nifJN2KWpswH0rmXJ9kjO6n8aJHp1upN3l3IQ1I4bCewLLu3Db2zSqZ8kvpOq3D0mNLeYkZ/ZQoy
ofQHWD5qoa5vOphL6/0lNwPpaOG1xECb1HBj1i1vegllIVuPiu8bZxdHlqkoSqfZI+a+Iz7GBdlh
riC3LHu6DjaxbSHHWYv+4gRx+p8rlzZnZSFZLlK+NZI9e1AN2VsyexFSvvB6rE2gtfGCOGAASkON
sjMdIjKwa0w6s5J6Jvv9JWy7JAakHGKjdqPo0lotdll+W2Tm2E508eS9p5txSeF5KJpnxu0UySo5
zk/TG0nUp+d5lMrlYNGoWNzBIz6QEJOqmBr9Lsq75JDV4qdK+55DT56TFDxnket0oIy88sUqyP/B
aiFj7j2XEIHkMyUb1zQHP3JWMjAPGal/h60sc2POYfUEtMOWYx0sH9R8PCEjXPTAc6lS4UGezcGO
ifG1pQlCG7NRsMBOQJvIfr7k/dFt006zC2I708lBEb95a6AbrMJ48W9YWNcchbssTmp8HmZRG5H7
OaaodVPdBG0CQskR6Sxv1MY0PkG5SIsgN1qYWJeZmblmWIxYU+DEKpAolaXqLEZsfj+4W+iOYESY
39Bv88y8wDl8bvLsC+YJZ/sSwLRcHJQFQMIgiJ8BZxqTrTO3WjjLKEUXz4ozkeGFyq+RMrPha0aS
2EYD/B+cUYNnXLzhRzSwyj0JBU+8W9uP6O7uVZ9Dc8tJqqN0wFRXn6wO3wHHKS9q/ChSH4dc5uQe
diz5dTcYeW6U7XEtHzjvYC1a2v2V+DtmbZFV5KVn3AGq523ShtokiJmgAasrAx4wWxFkkqQRGhIC
o0T51fFNSsI8IqisfbLifVEmLNOA1tNzLQed4dPPjiCY5+gsEPMaozd9N7tnQTzu9bdEGzlZXeSN
2AxXWJvkHygFWNR/0NWW17CXdnLUaHIQQVkB1z8El9nxFCnI4S509jXrvL/4IgkcJ64csVxMJwjZ
MwMa59T+R8hH1k2DyCeE5MiXPsYDDzWYGV7abnJ3XCurXSG9SToCYTaDcIG9SCpyStef6lxoPD/V
l35lfSonKrFoBu6kxKEiKBl6E4921YGjAc90xjypjmNiNo2f5ux/1EcTCLODyvJqVLA36Q4Za1Cm
Xt4GrRzJf/UoH0qMmScdG0E6HZk6quZCM0yZmbhA+Z2+UfpgcJ2hfXSmA6oQKiEUcsFJoh6C3d9m
YM/OkdbgkNcCLVqcgHFCCh3dc7YsSxjq687EmGsLHR0OkI6CbJjIl/ej7be8SLmC6OF1W+RSxT6Y
dGFBMw2D5SNwbCAnG0mD7wFpTopIYfIPiOXmVwPkxgLCoseQRWSK9PdkGXHljb7ob2Zgl1n6UNGi
9v55zFsiis53WWVEMmpBHl89QGvI0PwSvS2qVLHrLeyunxMa2HRW1OaWMormWlWEG//nBvo59WKM
w9mGeOd23LTOZeaWjPXV9C0I6qcPXIVn1HuyMcvOGQBW5UCDCuWJ+e4tzshPwvFoMzyP83/wgTaA
yfmffukyE65blX3AIUWKnCmdWvhLzcvQO4cKH3tMXqJBlbnLf7vShOc/9RZdyU552NzTIFLfgCnN
g/TO6b/6lh93Vp5VkiwXXGZG/8R+IUQOvR03jbK5MzYjQKkODw8l8IXgg32W+cqiLy0CgzROxtdj
1+eX+dp0EHXaecw3AvnOYgeC5EwjIguVa519afZvBsJvQuVkO4glFlrzRAXuGwxM2LPiyoPAlcMK
PEBDVvnEIP6SDF4ae/H2PovHQ51xmsRgrIMH97J/y8APHZ7CCiPYnyeVSOnVf2/KNbd1yW62pix8
aroqCOP2wjQZ2gnXb42nnkN62dqJCjkCXhQ9rIrAJr/zAmTtKmqWdclf55cmt1xco22fHfD4lQNB
OF/DsNK/LCLT42UopjYmonVTaqmVk6Lfe/U2TCWTqwYKUPKq4KOsZp6O+onxBaBvB9GeDRLqeCOa
oyVXx+TxJ64GxPQTAPSzqCYbiIarwsMns1OTWdI2HtYknIWopTFUD8BuTsotAMqQ/c2SKP34AMLU
hrGu8ytfSNzbUuOf3uQOM0p2LWSZZ6RLH96wQ3gKCA0tbbrqOdb6lgqy5tENelqyA9Fim159mqrz
6Mzp6JgSfdIaTvqvC9I0Za4WXBNgwlbmlNnzASHFEe3eHUMWauqFHXlRbr/09bIiHRRO8RZEGyCR
Q0LPnNveMtrWk03fRO8TX9jphecL/LfXW4erd1E+DcLNS+C5378d6cQgYcwXg+a7td74Ija9wtd6
c743x/RVALj7Fw9MyKKB3+kqPpF6GBDZaPVei+kAlfD4v1HQ83ZYy64HhLl5+mOL11GZrtWY+piw
RiSpQPnDyLyyhzWHlIOPOASSitOBK2WpR1sU5epsUF7M6PKzzegxymIP16Hmarz0hcjB+6V8yTPL
2x0h1yx9ekjoisIrXP92GVRtlkTUwsXcdjUgdNwdjUzS5tI0nav/zZmv3R+Nj2hCIbMkVDs5VQsP
LMpTlSHVNksIZZen5u6L96ib+YvgnjeIjgobG+LGui9FaGnIv32XP9I0w+O0SOvOGcbGDpcAQY5g
i9dhTM1CxRYRIQrreo0Lg6HtWrqdUHxfaTjbpLn01J275e7h5jOp9AesEeh3BYkuL71uHLeeZWtq
4VGa06MOQN6SFwxJ4lerq+CmlgOBPBjpz9C8MYT+Y5SqgW0CqH10QZPOXyNryqTwOZGzZtfz6IM6
k2qfxm3qXBx9+CxJoz+5NB+igO19sSZVHSpKV4k5c1S2Wv3uwHjbA2vfCtm92RxZzthFIhuuNfIl
iH3uFUd/KREzA7p04zZQHvv8uk2OZkBM2qzNpiCBgjqjdJbdxjbSPOdzj9dBeErj5lkJBra3B1xs
hyWSuDiLz4YnlWefQS87y9RvEXR7O0Y7JQKOFMXDXIlQIQr+9SMOHq4UWDPnaSXSwqsZXBQ0IBrE
todZZTmhZIDw4eYufXqYQ7LujbjUOGmfFDWu2DptJLSnH1lg4N76oU6/pWvc1jfQ/LnPmPGSe4Lm
Q+uAVsz85bkufuXLISfelo2EjsmQbuToBM5/QuVQWNwBiRTdpuvoFGzeW3jsClTBA+TaLAcFSXow
i92fUMW3MvPsjO9Cs1qO300bilhvIliVAAK80myLRYR9HFhfzjN8sJwTQJ/zF1rfJ3eKcX8NJOpk
3yP7AHQUnhvLpoWA+Wy3QPlMmM4luBvcQVlNEDN+Qh55wauiJkN9+lweaWAKTjrI6Aj1Rne0zDjm
VgjFSwYBeFliD0vI9gvJCP0pXDsGyQPoVu12VrxadVhg9ZLyGdF0yrDSkwNIUbFdkHB2y81jFl1t
apyebBQayJNGfDoIzr4HnZsWERfg5hysW7ytVpkpKCL0dfgPpQHu0RAbX7d8v+kPBn75NYTYR13w
CKHbaJLAaSMWCBQJ+NaQoZmA+tdlg4WnFgVHu4jEKsGCxNcy7JzxzU51T+UiRRIWRjuUlOIH1Yki
MClbz0hT5qWpLwDXoXTijml2V5d+bex8WsNvVeZtctmM9PYmOn1+PAVEzftKtRSv+Kl4Zttp2wMk
dCas5hJAxVSbub6OVuzJJyuW4esqsQXJisyjFGOAvf2P8aACcWwODTEVMZ32uwcxSSjGFLjhQ9ye
iFmWm21o5UhTUL0ynEJ3As3g7THG4scZW7cP2ruv2X+zIt7WXPPfEChIvwdM39lxHLAeIvxaiKbX
viADc2Vwr9K1V43GTcfGT1rjyFB9+lxkZvLVc7RpzHVafD6awjdfxqWP29STOsC+Q030OjvrQUHx
dZvG4YHye9YjKZmWUCFrTz/ZSRzTn68KELc7afgT5eEs79wbXMH1c2rfEuUzJ35YZooXUVg2CPs8
Gf+M0DkWPkgfBjCUo6+c3LEuKoeUWlhkyqutEudwX35etMiWchE6HEY53gY/cSRi04NJsO0gtlsc
/Kg0EcGlqzIExqKQBRQloqHfl74BNKaGer22RE8V8WEvLq2jakCtfI/O/tnymX8mzDTHisTghfyP
8ZBnwccr6Kpd5/4Vxa7nptyFlj6K9hzCJRvPVhq42Fu+ZRRGZbg9VexcrxfFP9OmaoAsFF9fi5XU
L3ToSaA9t1MPyW93xvR9ZHI+Efili6QG40VHHDPO9070m6iq5tzrDz+RqvvydqcLV8JqSmswWKyv
t2hK1bURw9ujedRilp1pBG6EeepT7gAc0nshB8DeHxW4MExsM9HFR7PXngIQI5gyOUAI2S1glnOJ
i1aY8eMXdDG2T7OaWqo8U6KpvAq/OuJcAP1/UewbGmhVudPmesC3CfgqDrjs46QCFKFAgo0/iEGz
Z/Wqe+1yvc3oThKwNkJYESQvlcBNpbCZRceuAsBheupjBjy8h8MTKYpBPCxOdzp/XTqXoxuE6s2o
uc7Gp6iUBsoNasS6jDUWp8Pr3Sk++0dcGZjcUDt6J7ETPH8XCTIC6rgT9mWkArO0dvyTWrLmujFI
+a5PJ3+grS8E5klXs1kTl5mDryRxkBK/eIDRfQuvxBRoRkLMjPelu2HSaGM/MVOXg/metIHpnzJm
4GvfJbibEXPdwly7EwogOuftclEIov7Xh7P2wqNP7FQsbDobk1CoR257bp5uPmEk4ZoaR9GYTWLe
n358sV95Pz9zkLbjLpwXDvWHkboXpvdg0JkE4yHBDYw3oI2etBzKSi36OlbkzHN8gtF86oQPehTH
gWPt5TLNP1QduMpBojqSANSmvkQ99ue0k9+7xT/U4rWEu9alHKgn3zlGPNVx0mfK7qpIeFeKTHE/
jOj10+84YPWAf1LhYO1Rh4y5TIjxg+rdRU+v4Q3V5UxX7dh0tHdXrycJQQUiYLwf/7XGr4+af7tr
Yx3o27OLFY4GbtfhQOsYLeJKVBzBdVjbGkgH7ziSK8aEChHBK8BmH/xBLIddR6kk2zUiPKrMLGd2
vQoN3PPUSxxDpI+QVru+Y89sr9vKsgFXrIsa5dFkxZYROLZhNNTbv/WTESpfuSF+EuRfZyHtN2Cs
wrbpw6nSJmKe/vqsEF3PKwiQHz+GfEygCCZcalbC1oc5aeejUi7jzm3toHqfSiYS6P0Cht5LhXnL
xjsqj10GHkM53DLWyVMhWXGueriByZ0OXwQYxG8U5cUHK2k/LitEHSCG+QI26oqWIhbk+6gBtZQi
m0cY7fVgawtbdknbBeQizxpvFExowxlP/XnM4/PZ70J5hx0YrQIRMzJKcE+pJFzQ6xm0R2+GE1Lp
NpJ/5FQr/i5dTnWeMobWlu3fDRrFGUw6bnKXmsyTyEgC+Va/6Pc+t75N65Nk6ntV+Q7rwvS/IUKc
Mk7+WLI7DmqG7rt4rAjhXeZXcyvcC1QlHaxvw/ZtbZq6+uqNH7AKo46xCBQ48HJ4sf5mf9u56vJ0
VQ4qBTe41VKuBCHfl2DRff25JpLJKHuG7B12LcuiZq0QajUWxDuaq/kuzJIryI0CVO3HMjQx/o3V
4NIcXw43n0/OBX3rML3wWxOOCsOVeZH4r2a2CmwH0fARGyddCwUp9mRRaqnVEjBYRE2HlF3mpQ5f
La0MQZELFzVH5PncGCExg5673Q7h61Qx3QG4JE/DwrXZ353b5s3R9QJHSHCUbIirNhZuourOmHef
rdG74xjQkI43uiZ7XVPHy8v4M4xLeLICcRsPSn5o/u3WVBT6c0/jF0QUIvE+CpkC26vi4yc88U9p
W6Es3l1g/j3/KdDcayj2x8cu3AKbwZgMf7SMYHDAz1ST5t11BmRPyfaR6hpEIoKLufTH7oYgWa8k
/N8PKIU8zVQ+wDxHFYviKpuTjNsPBq60mG25i6GNj92a2J9AX05ALFzkJfx/K01TNQ54bYyl5S4R
Tp/i5ukhWI8fuVPLJjGLCyU9tVh34xPbzfCnukS3jfuZjsdbB5lJ2mc1X5zhBUUFoYaO3GYGUb+9
eeBhBMhMXl9SqVz8Ophoci99IitlQwO9A4LV4NufPGWdvmTAx1EHKkq9NGQuzn32boWkQEtYX3wR
k/lomV9UsRcZ144riYymKKlru1HCrzqLUrQKthb7lNarqmYk3AkMki2sNOnRgOzQAP1EjmHWZr4a
FnmI2DEQ1FKoQpYPwZU7dVM+3aGZgTBugKZl9WujplyIwr8dV9Xle+xXEiXmcRmB2gVHBXqB9g46
BLT7vUX9uxitMHZJ4q05CSqy4D1zzOYQx3vorSCDy1ILDYx3P1fCWMaDNl+yaEV8/bNy5ZBOLXHP
nngRjI+jUEwJWzOpG0LkJQN10CVoyO3teJlv1N1Jaoq52cKCZgzeDKjXlPqK4vuiUiUjp+6xRIEU
BJ73ld3+qpFrv2sJbt1/u0n+DBecR7nykqIdk90/ubf61UfaAt2sSPHEAv4DOxcL86uJQwwTQB6f
sPLxbv8Dy3Ixrxi0Zpk3pMqhvHtBDU5tcbApiL8giikpFc3yPeUPWi7OCykmMCW7U4oJsFgAe3be
CCpxG/c36Wyf1a+ykLieFXIQQCUuoL2iYJXdczNTsVgpOE9EWhIzMl+8+JFZS71eJk3juXhNip/N
YSk0niUORU7BytY2uVkXuciutaI/wXtGOZX1MJk/Wl85g168iC1QRPca2DYwknIjRXdq/dKOZf4p
nF1YpzuojEzmyBFMqUFgPALvapV1KGJ7jhyKaw7OVal7ATMJM1q0xEVxJRhhhQ5bzLwiDUZzB21j
+5rnUOYOzVoOdPx5d/Uv2jM1aRPyc7ZEHnlvHDdKV0hTeqnTLcis4jVsTRwCbvzNCZJhK4m0iCNb
BDSB1GlMTXpD7tL5BcUvq0HYZYEz2sGSiTdQjSkDZnLi+s9mZtI8wxijcjdCNSH7YyD6neubvEeR
zVmRO9G4eWhda1l4FrLTeQMHe6o9NXsl07wQqVakhAtxHZ5zkOwrV4WLf4X67wSgM6xZ8ryjZqNV
soXvSesAjnQmb1ZxWwZDt9s8pW4BbZBRTtwVKc4jPn8bx84EQT2R9LsBSoDraOxAA7jIql5Wgpb4
/aTQpjU6nrKjXJxAce2Gg458bS0ncpGR5Q67KZnzZDQDLkuyWWQyuMRwwrHTi5P4e+TPEmGWgqU+
+cSabysgYxOdLx66YrbxsdP5SyuyQmCHiYaCRxvGhLLeVe1r/jORmkf9ZL20jolvTILgrf4DRWSr
a13IQCVPWMfgOT/YEdj1UHyK18SFxCfVTrcTo6VT9yIBPi+gsup/syoS9UuvWH4PCrvyWlN6xT7i
3BUTnfctL+/t1mC5oH4VpYhcj9LlD/uZ1yK4npxRqLzK/LXg5FJM56poIrRmLodoaQvYHOPHRlTz
pIc8dUlo04Z8S8xKN88D6hIarzEmAR5Jme76rGZcX94GpqW7mrF7XS59XFvc/+4qg4thun/rHY31
qbuOmeJ3c4rNti1TljWzc1j2Jh0nTh0NaKfSkfKUcqHKgFywVbsTCCU5yMcY9NYSVLuau9SHUICV
ZK9mTwwL9W0hMZHIROrvxME04tPBH4RLHzf/Y8B9xoom/G00jgD6e57mUsN4/vm6leH6ditFkKlT
bwWlVbs8O0oZQHaM/nzTAwUjN8PmgqXO79DnomEfZLHv1d8C3G8TG5tVmWTJ22lLV11vGk4y46+1
kXdJRDVvDVwM+tSHRWg2K5pt7nVyspm59XmBooYveXH6pVpoS6v2oMs390W+eRwUFdarCHAW5RNH
jVCX3GDVVD9lkzQgTMiIa55VGjRyIktCQ95CaVIkk7gG0eMwx7DS2NrttJFMEk8Lh/WCB/aA0qa5
DLy2GXllNaTO3xYyvvXZgfFFHrXyPABV7BrPri52zWKTyiCrY7lNGMezUxbP+IvuWtx4r/HN5/s6
mIqXsvweQKEC+jggXGxny8WBUYUTAKeL5T8/heScZhlvHMiGPlEuMFKg9LkkNeUBWfaatKTNy4If
fIg5Rw9sgMlEuR6OrEN+frDCROQeSqzZT2Nvnfhez5V+IpO5IeU1ddVJieCSAm23ibpnwBOFT4zL
Ej69p7ADtAUDLn6cNtnAaFRmPw/DmPfiX5OABeFocAOEgetdOq2zLFnM2OC6V6yLElVdMEvjI1PC
IiFE4tALmhY/kIxrptfpPoMVFr5Cb1HVOekcu7Vq7Wl+P8D2qZD4oFKng6lEL10nfWnS3IZMQ4hP
Ur3lJg2t2HoKaxVS9QtvBWLkakHZpztCadg1iuqC922qahyw4yJfP95yocrtjGaj0XqvzKo4x66V
fGJJeJm/qQTYZrPJnyzghidfOeEghh+t7emj/qI7K1FB0LymH2CNMqf3znCUS6vCaMT0G+d51IZ4
899TICrRrpKbUDTuDUgJRtA+tBCKQjlsY2geXAq42V8dLbrR626vPxxoO0M8nM4UHMnzWiXf3BbO
CH/sukD3T+O4124FztP/s7DuG3vZQotTQna3Y5tRhWbDKxnODorHbw+zt36zcBLxzXRyjk/qf+H+
+9a6q908c73JmG7YRiMEQYEW53ykK0Q4MQSaF57zS6g3Cm1aNim+gPUf1H4cQlKp3dboj+/UicC5
IEbIHLTcPs9aLOCfANQhe3z9pJtFO7ihA/QkSukLiCd5qfF6GZKcytmQ3Gxaw+MKxfUn9LkRts1P
pHKGfHjxSrbYh6kGH74ZU1eSJAJG699OIXoMoX0klw358sKfIAIC3AL6XuTsfqTl7nLAu4nkf2N7
Ix06khl4i6XlZ/wmhoKzFqXKf7i8zWhGbg9ktA+FUEf6+fZnm6vzsvNJJefVjKGT3q9Yl5wNstfh
mWfQhVGCqoXMlm+pxKH2fiqxM084RwpxMLnBwcv2HM8ODqiuCnH9SsD47wDBsSZ3Wqwau5LwptLN
XQnHEZ4cgG6Rxtw8laDIYQJSCUKPSo/W7eR8ZrsE6YzquvNq3O2UJ9k3ski3Kh8w0W+mML5d7FT2
0iKSDenMXgsUJelriDLKJOtVf8rFTBgfItAE8HL8n7dnAQQnfFqawP2knj1utm8PUtrmwfg/kmTC
siZS9J2qBioYjbCzwjvDuXAZNW9zqGXeaD3MqU4zCPjNbcYm9nN6mZb9Yo8qyRzYBkSjfC0N7332
oy3cShwSyktwUUsSNZSF0Lk28u+Bd1Max6yG0IcNWZeSOOVYHLomF7IX551cSrahZ6oWlrjSefM7
6Llg6bYg54bhKutMbMEKu6j1bQ/+m2mKKXRMISXyoCDSPQ7pHp6EbeP4ErFpsC1BeKphJ+prqINJ
xTxTfCq4/5mh2lXc8F++1JK9U+diostiUH0L+/8XGLiF2ovodGp0hBbbvTwvX4RokztUbz73LnB9
arqi87gh/yU9lk3ZY2htmfWfzMPIgkwMmpcjaSFfovzW3X8+qPUouHsItYS3Ff/PgeQpDLlz1Mdl
I8jueo6czFBdzb0dBt8Co0W2C+e7mZKzBmhs8++Dk1rORwylGWGa4VQ6zt/Azht/YTd9hR6QUktd
oxdzY7jZS2iIIoC9VdbR1dvNLeZLysnm/L5Jl8xChpgzUyWLNDyJPqG/K8dJJSuFEplQ7Tc1bOA9
+Mpey6EShesq/cOBxsYI4os1XZTag7t2inlCyM1tKNLJZKJlZPonfYsdPDbPmMsFcVsoHK3Gigdk
uGo9Z1bXvmKp0zolO6o0AERgrQ3qaKYYf+qKd2jRrYykjkMizPc5u8mUUKoCC91GJLP6uiiIXh6B
vF0EydKUaeHjWg94HlHNn5zOkW9vFyA4z2LwgBWFxd4vkEtj+zJEjPiM4UNu5hh56yu4EmAHFMQh
dVHIxC6GWUlQYTx0h4A9PwjHpzBLtx5uAKewIHyW6QZS8iHW86VFJq4+yn/zQbXuz2dzP86NUOJB
GsLFPqhYOXVLyUkrH89UBNju3tfU+nUxx5lnpXYq6AM1zz01Unh4mwV1GfqSJLpe5hxL8w2D4XTK
qHUnfnRsbEWXakxJnUScovZOCU89NUj/2niQsaMdr+n9x1MQ8cBnnrMPdbLVrcb3ioba3CfcIuh8
4bOLXMQPYRE+vBfEAfWNmKX5jfEGTLhtcutk1dlCkR7KT33s/nQzq6ylOdXCHM4xz85MLxDDCpCz
u0BeYiBltMvSegVN8HhQlj/5Fvk/4IJxg58m/hWZRVkYZ+NaGL/nUHV4uAlQKTedZEsrhEP5Lwwk
lm8byvkym0zGhj3fRjefWQgW3DY1SIXon/rlSKAEu6r7rnZEpOeavcqwgiDVcFvkAv4ATKX1D09G
MhOXPHx/gUpYyAlQvy6JdBuNS0JYWBOwCy6liNtjCezt2FjBkvuoL8SyQO7q2Wu2OiMoEpxPvLsn
7BxBQAvQRwTHyI5SdExMh/yxXVlTECkSsnm9y0HrC4LcnBBuo+TGQ9My0PMAnS7lecZounLaJQ9w
BfBfyS+OTjxyrO5nMbXT5XcWJBEmjtjchHgmuAxsf6LfOttXK3AT3GjuUqDIRpwQWnK4oSKdjdlW
/CMb62g5UQ/NwDXJNifYe+edtTmp6zilD33NUwGAHNaJv9GIfB4GpTTzqvcBFmOxHr1eoWs8hpqW
HxpecSTSKGKsulwbdaLqjJ3PQTf+Rh+p1gmdU+phDYAJqjs/hKSKtD+OFeecxLwV/ztApgnWwHJK
GlQki2tJHvCjVzZXogZKGNjuP3gYkAuT89JaCzPUmKasXtVvgf5r0yxiccZpilD2VVlzNNC69qms
64Siu+tt577XGJO8Av++z5q681C2KPFaypcAXHqglisGEtD6am1ORGZJDy8oelr+lRdWm/tO6uLs
Hq7bSQf5PV7zLTA9ojgXPQG41Gyf1dBqUMn9ZOkwFzUmDihjzzWFpEiULtidB+PR673WrNEImZxj
NdE8/D0/X0BaJWPWif1avU7L+HO7TSsp171H0a3n73sc1ZDvD5Xuit6s0DAWnYa7igVUmmZmmb45
SsU08iwJPD7Sd9weyPICXEwwFATo7fItFH8Y5yajBbANCrbNXK5Tas8zXqJzf4TatHk5G6zNPx6A
/b9M4JLMsAzotPZ/1FF8UB9vfgdG49GLekBZsIhEPcz70h1n9HJWkSQyHVK/9FAp5E+UXR/91PFO
Fag2PegsOtXVI25L9fGL+64CaJBmIBt4EplExSi3b/puVOd+hb22oei8a940ka8VaqcOG5fDdXUK
V5iCZbO7Yg6po+Nl9kyqF4TgEL5pbxkC4tUWfadHzDPKKAq/zlfhcppELYDByRJy91byF+OdF26N
gIUt8T74ftUl1IOOpsXp9scZLP989+PDhe4cN3Eh5Iy8UauW6yrwnQK0/hyZ6O4wzuFArplxrQsL
viHKdZvVsIqXZRy2wqlpUqYoOYX2dxWEhCDYJk9agnntFT6Fb/nMiiNJkAlnJEopVNPrIsvtmUqZ
vxlALnoZtYHq68TWfBDhLNNmCSUjGU2+rbMojWzaWBK6W3jmhcNCXGxx0oyBX4uTkgFJ5t4drSdi
M5YVCEpgbD0yYUVt+iwIjZAweSM8vf8Pg57qN+yi86DY3bVwbOV0mGP2pVMzQ+35AO1VPPfcCMge
jr7VZFz8ZTuG1rnJNQ4w9xW9lzW/ZI/gflwiuuItVngOIH3qEnB9a1rWn65XkjlXyYR6udlq209b
3VZsov1QcX0Jn0vKh20EXaige9e8v4PEcYnoICLqWD5/ZQ7srcr5WkgADe7Qc9CcuiiguCCtD7oa
uZ/Ai3iBh7KMRouv5XRv3g9ClSfn9U6u2EtXUIyxZnhxZzksvy2xlIELXRLWtGIixUeIGx5TxYkR
0ylhjZT0pTn2ukXF68dsQY2aU2bfKaNBMzH/laoK+EyAapVTZ4FhDemOJQET861nbXxCuYB7kV7U
eYKPq/nAt+o7YtuJrwWjuFCesk/+YLBOJmMcZVM4oADisxq0s4Izr3NRj7t3U9MbfOBxafOqCw+w
EBryal45uMCATKF/EFlooPdkzjCQbwkm6GFFXx9VxbPvQpRRfpPt9HdpqvDjfB3KQ9J+6stAjE7q
mfqGqaFEYBi7G4lF8v9WnvxNPqDlg53GChCF+J5vW1P1lVS+pY4RIMjeD+RYXEZGdurGu1R4C4Yo
QIVcouZG5xcHoIhzwPxGOUP4ILNAmfgFzZDAWgedETKCgeOmbADdbXgFajHr2T2bwOwm978qOcLs
6t5RQcjQiiGpWhYwKbOqFl6FoUpGSArW0Ogxv5r6sfcGK5UEpR+tS+v8HnKFqpIUreDZbGOPC2Qc
BVgqyjiygubrRGEKmDrh2AgEgCJTobPgzaGc2dBmQNHFMaVJ9o3XcMHq97dwvjIpH624QC7axN8e
XI4sRc/x1iQFXAmskgH7YOkXT0Rr7h246aOYlfDzdRxDcTqKJ3tYjQC9xcA4j9/LerY6lwpd58dz
Pfv5/IJArAL6ntOT4KkuRhte8alxuPl7HCyCWluTbd0B7DLKS2MS4kNzhmzLJOVdP9bdndGVNI6x
gYJgVpV7xaNIUpKFmajZB4U0ru4N+kxYlloSG8K49pJeiJjYlIYeieExnZ0B4g0qWEXap4qDThzx
k1Zz9vvdug9XwDronLRjOdtL1ocdcfCY+AOxgnDT1zv9Ttg5sTImedClosvWuMb/KAjD5+R/qK8x
1NrQazgKcF/SCfAL485WXlGnxc887xxtll+OMs6b4T1KP3C0TtqP2PLEV6lX4KTczBdkT0r6vhcC
DLLto4gJzR0QLNnz/83cP5zOc7cYdj3Rsm2M8ipd/SgdZRYJU5JewH1JvzcJJufi9symptkWGytN
HAjTeTEvdpqixJW5w/pjMtG0BEG/BCMkcCbY0U0i5oXm6pNhXJ9ElDfQWT9SVTS+Y55IiQg9jG1w
IQXRrN9w7oCmWvFFTE+HFFPvkZMwprd4IeGBpWanEGuCL7AEiFd/AW9MORPhE1TGow0aryAS0hVb
bQYSvOlnrb19KhHkALxoyzlKqCeaSGlhf/AqpzZPPSWaUXLncn3QOAmd9giKyMcNYoBqp6rD0tsM
9GYB1PzEbcrW58tABIgyjRQyFEqbjbEqA/aNJ3chuJmyzSQcpytRnJOTZxHmTzlMeXr40dlDyu7x
xak0YEV9xURvwfIFKCnffOMSSJTaCGR+FjHAmWd6icYUTQkMUGrm3XbtDLEmFCt5gqQ+ZmgTj40/
13/f0+bZ9k+rur3Cv+Az0+KzfVt4e5Xe0JakfmkHOAXbFzAA5JdAkGPKqKXU7LdxIg297Qob3rtY
sS0ybasemnSBpQ/LG/VERDSUmzIx6iBYt/yA9AtwAVoCv+Jrl8ssnjFLG9XCgrCIge5QwrAm8Beo
MPg2v601ISHcggl39494JHng0SQA99fn8yIdWHDlbgOMfFHwxBZ4/ollNGkU0EKHx56C95Nj6N6e
TnxpIrPtNSRpTddkUJHADO89GFplaOmEigYlCtU5LQz5n7GwRSJ70AhjSL299y2MGMjVcGtZ8Dcm
ZrDknXYqzfwuDI+OE8ctHZi+oRRI50/jZV0EyyhnWpd1pXb3SX3alalwg4yM2ZbK6pmLWwF2CudG
Wep40o12Ka4tUKm+bga6if5OkJiNkTAI8Y3vSdNDq6/2RV63eBMKgkUgTjP9I6ChIVGA1SQu4BZX
oSsvKbarUTptI5FexQZ8XEu/OkSsS8z7VXgIOLODej4nSn3QPVfy0WEsYlbd2qoHZrhgOggXZZxs
heFfMuKABCoCNuKIuaExbbmrl8ahyl8bYGU744v2ne18iiF8FPRwvLY9xfg3r5W1T9AHVZXa40Ww
K9WdXKbE68iNpIrZL7W77Sw+GiqL7CUwJ+8vTyMTN5T1MBISjx8mt/TWs44i8gmQaAuM8gtjTp+d
vHVbRBDzWYFKGi9eo2dESV1crYOA4117H02UDjXSTcK0okHgmKbbKK7vZ+TYFqRQqnzcVwNMDY7i
uLv8z/SEz09S68F8VyzWpp6wlHia1jgcsticf6KhCMu35DlRcIF4Mea2S2WE1/qRasW8x9m6GN5u
61V/UXuryQsjDxANSnfvRh1Flv+8CoEhtKfeb6bYHaAOpb2U5Ann/oyo2RIeTHOwd7Um1kwIYk4q
4RRgNu3V/+j371OGGPztql3qJJV+yWbiWctG1EckOkozY4UL9cAP3DDDJ3L1KyMKDD6XpKoh3YqO
kz+8orpEI8+9GgifXsISXBG/whZhmsT/KbG+Ob3SaGdfeAI1kKt+LhVoYSL+IXIi2+4QdFnNlMrQ
bfVKQX4xKC3uR62DLpqf5P4hkJbKdTTg2Y5oxaZUesSehujKrM40prXUzbkaO4Qx6dLUA4r/wH55
iJZDZ5kupmM21kH0tsSQPVPJiHB6bb0a6KeNZC4t27DHlbKCBM/dElLHwk8uXWHI4VQCakDF6r+0
6YYjfqp6FBUpJNbAtg/0s+yN/t25nRwvZuDKSswqMXmS9pLbDlBlf3OU4whKrOoR/TXFilOAtJ/k
r1RmedSKe/jzcCvk/vKOVlssrLrZ38EmFHu+E6lDtoNQ0mFAlxvRibRQEe+hRYHtoDhaifXUEfRg
4ATYcDOkCudvgrfQDzrt+TwlZIAhOFSevoUo81KGXKVzuwPEwyPN4mqQ/sLaSdHsjjC/JqtWUKvb
menA7hNTEP7Li23Ytho9/j8uJEOMXdLm+LD35+HZsqH1R9gMkC5xRQ0gn2GzU4JhN0781rS58kM3
E8vMvKkBTIZddP+jhNgI/pJkcNEjAumweLIrUBuvTkJTsZg+JU5Ib+RvuepG83NdmAi2wCE14Ko1
2CWb59FvJPjdvMJPjR5AUL4Tgd0+mBUTP1l1EUzsnmaCx3BPWGEzVT9KRbktaY17khK7y9cImoCE
W6c6YgJ8FCD/wbKGQuhjWIObDGwG1rCwQ+8SiOysASASmgPzuH5wkBMjhcYyRyRYSwViPxz4nncF
3AY+czjQsGhTvfZMN5gEbUVe+HG+GaR7asYTuL3eE2SSH+X8vjJ5tLje28ti1FxuQ9aaxwJniZ+P
DYZ4dLLoy1oCpOBlp4Q9U//o3B98W7Vlj1yDZKr+rv/snM8qTK0F5C0ZVMNydPKKSRAa+sM3yseo
g44ouhTx2qEemNDUGoZHE4vd5ZCacUgCOQowuzvv2dMt8TQ5fDy8t33wS2g9+hGXDDLzkCrWrF52
z2gi5wz8cnodCgOaaM35PbC25AkOTcbGWy6qrMfl5Wsdpc2tVJg77X0kgueE9ahtoOFKb6XR8RoB
s+uv2J8Bl7t8pS4hJRt7Vfx++Iv2RYQt3WPP/q28/JIkLXVD8DJb1kqpaTDSzc/plAFUs5kDNm/H
zFkN9kIBoeFEJ+R9PuGcGU5yvU2MtpzHSrESzpTvs46prXPSru5oDBnG157nBzpBMlPHreZCNOm2
/+cQS+VX3BAbZyQaOz5TrBglma18MOo8btWU6JIDMWP/Pt/Q//AB4gadVS7vAOryHb69XeWZxRUY
NunVDHjVIzvzy39ww5BifayK72AVkI2iCYccY+p/7nWqVKUGzK2P/kFXbmIN4KOqrQMdCNi3U1du
FODXO2d+qwX2wZ8nhHNSAhS5BSyvq559PaPxAJt4TWlMSbHo96VmrPXp58XAXjXDYEETUuylP1+Y
PhN1MTOltIZNOJ2fdW//GJj7AUe/2qQAN5HAmq2yT3gHnbzEISSWmewxtj6Mv2qdbQwrKxDlfEZC
kIyjkSPYAkxud4by6dVb748Amu+TNnLsBXPdRxO4O86y9+wxv8QmEvnHuLsKiio83zPS+9J5Es/R
hfBajr5vDxBsfWJAgg/6Ldey6wEhH3rCeS3XQifF56k0gPxiuG0V5Ho58jVGNdugA/I54e83wXLN
uEm3QrQR7YfdFFZsn2W8rt9KNyo+EcCsVr8bygCbVb6/4YmbFuIWlq1zrbbQvrmYRJ1M6lbdltWR
YK+lNf8I29DGXCfzO5sO/AXhmq36HtnBLoaJ8FN9ECd8Z4wg+2lB8fxTAWV41juvEmXItxhc+sCs
jv+hDNSA51YrQk3D/f3xZhZKY9HWGN0+3F0j+czAd3S2lTEtU8/ozKs7i+KptNEOLs9dRZTUglU5
WjDjG/nU1gn5y09FIUxGG8gxefX+fziDUEWvAcd0qVC7Q9X5ph3aoXG0C8vFRb6Qb1f0fk60uYCU
t/7F97DMk5pJdOkaqXEjOAYLpV6n4ZX/O8AYS2rEkjaCDJaBCi52vFqcZvB0QP8zWLGaXM37X88T
scDkwR0yoF7lQ/kuvKMj+g+uAS+TjjMuswujxMgBm+pUOsYBhDq9Mv3tFJw/sz19oR1N3FtawMP8
Ss6AjozGAEKd4pDy8jmbAvPsw+LATRCwUXC8gx9XDaVYe2j2I/ga42nKScFPCYaIF9/J2cK05UoX
BV0GOzAD+k9LwUShsjhqFoyAoXNEatnS1iJL9WiGbfazQVLlcI0OCOe0vph7+zbrDsRAlIkAMQsO
Tor9daF5hVZr5VupfQQwPNaCftizPSQyWG3tFcyeG9U9cl+gqthoE4dt2zerrkknI0PMWc1ZfbHx
kzF6mGgDZvhjvL/+0kiY8ktyMM+jJfVft5pj9CgwZ4+4bgdliNUieBsJQzxp4ya8Sb7EXI1fXafE
UG+MCY9xAraePd2eIV+7kTiNUZ60/SK+ho0ThfJ9frkN/hDoB2a1o0vYWcpQjKZ6tcYS3KtKq03b
S/lUpIqzWzFygeRV127GlADyDO44UlD6DIrl89MPZz8TU0c4vqaviaV2hqjThwqzSdwoLQ9s2lns
gnSAPs81Ucps6i3UELFePlA0U77XzJF8Lvue6sWrI0w9VMRMTW+zGIArzE4+29H8HRnudkVU8HiI
CW0XN4hySbbggEmsuXpBiCibRQQP6KSgILcAfNlvoIoLfhYObOyECgXwrJEXFUdP4lIrlWwthf0D
YRtOvTf5FRqIo59upjIb1XGmfAwdSGt5dzBgMTZiTidQe6rkQCtpq6ef3jPs2qC+YCLuhQInq4TJ
iR5aU6ly9b5/Agt6e4SvuZYVeVS5epBDodBNScyZ1IXmJ3MMFZNvmgIjP4WeKdJuzetXNBiZD5Ty
ro4Kx17FZwK4c7ZGjd2ei5cfFPromuFVDqtV85bn+rolXTeEddbbb5WjLG0ci0oVCWLmmXt3lS7s
0yonKk5/wfhgaaBcEx8zYuNW7eq0lzhwMMBbhkzMiH2zLfjlGo1ptKNNlwAYzGAzcBOFlPilCxOu
B6FhgiF8lT+iONVINYCQ4SMM4IvY37ZF3O9VxzuXXEFhdl6bkGaBxWoJPSW5Y0g2WB78EtvfllhO
WvSAQKYPn4ZNNgjwp0cBQISFzY44SjEr8HaEHiGP4Jjk9shBIrzpIpZTLasn5fESKtiDoViO2q17
YDo4IKdm+WDLUCX7HPybM88g0321EMKC/OT9I2lY+sATupucm/gHxDlNV67NfZzD5C0dmX/YLbOF
I/YRSagu2ZTC4blDI2SUX4AQ+obZKMdRXG++tsZmsaU6qqehTu0TgN5kmIXwwDkt6av/EFohXw34
F7XgGZr3YGjREGW9rXj+8ppvuV/NCDoCsb0MASX3OO182maF1ubpvLAdsiA0ufLCv0CGqaZoY7pI
vl1WAomQzTwDvB4rZhEAXkrbw2B4+1hIQx1HBbwURipg1vcx+x3OVOi2iLLWeg35i3X18evqUM+Y
FavhrHm6Jb1zqOfdjsO1pzC7y1YZ0Q7o6jr6Bs0rVsQvyw399IerqgdUQVAXh4/uBdy3kWKhBAPe
hncaVMkLCYshw96TrMyrt/smoeB7eOsy3AZClULXdkJaGvpu1iooB5ocZE1G+AdHJ5EQAChfbUYg
QuGp63o13dggniqlw2LjYjtZZbsY9CPqtAFCotUjEHKBBzRc2A/32N/36lLVQzqXl4/yfjsILXOU
BlK7r2pT00yzD2+hABejZPTUw6v0W7duqMqlVfbXerj0w7lGL3jVXxZoVoA8K5Md8pBaCrC6sdyA
3yMHREYg7Najl4SLJuuf0DpSgy4rwd8cyyIOvwKr7vJRoUcMrtRzSIcp7pt9OvuMdIyLqSZILgZP
GzhOmv3SACpS9ySSpg9I4h/HMmK8ilJbR3Di97qKG7UfOauumXnYYk7gR77P8YZ3kK1XjL+Kd6Ax
qoRPEDFxQEIGAypG37oV/wxXE8S7UFYgJMt1LR/Tov36an9Pi2jcX0yn3jfCiZZgi9mPQKzNJwBX
IaJ9POQ6jFQ60m7SVSKzbU5C0hlEf7UlnhJpnA/SFfjx/icNJqVIYFzG+q9kzw8m55RmgD88Os3g
yIGg0blr3aTT8FrNKEVi+ZhoQ8vE+sa1hjmzcAZGRNgkpX61JsQqHwy9Ti9AnbdDcyApQCZJK5lS
nHfIO1rnHova5mWZYkVFnmDlIqgO6yYKB74lmOPmuBGWWJl0CqMDEDX6e9QooSX/g3Aek1ADb51R
4E2OPXp2cNuiWuI1ugl8TSxExdxf3WaVpSS1Po/iXw25pgtnPm7E0rQF7Xt1E+gWw2CqRZngkPdL
72grj64qlVkwYauyWR3XnJINLGxPLSy51TrK7TJZPeHFnyxP8yyZ4I8ozG/qoOvvc50f4cnyHtoB
lzjV5XeOEBU6vZ7LIYqTJVTMrcI4LPoyHftUbWt/5kkqj15VpDKxEwadF8m4w+Du9x7TEnBFnL3f
kcQNT8NMU1zmxXnF0Xf8NIRpmsM+bZx4QWU8yX6c6O2ypibAfUZMGJrSbx7Zyfpe981G8KE9agwt
0GO+wD5kDB/IRtiRXPbG2/t5bHPfphIpzWpgoiFdiO4ApYkdz6eMUAeR6j4dHoOoSzdoA5XzW6Bc
lqlOoPh3WAGW890wCeDzUoSpe/2woCjm1KxD6FX0xnaPx3Uz0sMb/58fF2NfLreBOjx/285ck7nv
LXwEgC341t/LCYmyxY+laOh7V2Y3E0AdFtcDKWlBIyhl3mY7wT3dMIx7SN3dawgHC2hSd4ZkdpMj
kIDP0KX0P49HcRC3hWm5R2SXdqq0aQByGpmjHfD5KAGkpzQC2ssq9/MhkpVBI0sVK7k95oCTV2ki
kuLWfSU/xCSa4uoP3RXAQD8Ayl4pjizScs87a0kEfcUvJEeGHgLDqg0cwn4Rp8mXL5rrCl8DA6p8
1ByZCOgIdUke6m+QX/zMv5zpVJuPKKFqv4c9bJRHretLpG5tNh9Qf8J0Xq9ALVrIRNewxlI8cN3M
QyVvA6tNL+FDvfBjHr34o3uGddt0Mgjf2ONh2XOWcK04IVuopqddGw7tZaEok0RUBZHiSXvkXNpk
nlAFypJ+ZpoajXYZ4TWEmsTyK58rSMtj8IT9vghucy+5P9AD1rChtgPFLaz8OpS1H3bLYSYFBKLh
UgygkP/UItWxA95tzGwCJAbTyKvE1ccCSjXwKlapB9VWzZqLg3oco4W1pQUfJVtIC7/hIDWToUCF
Xb0Ym2+vlUsFbDhe2e8zZ1ScqucFIT9uHQKw+oiDbKddhPnTxFoRaajbt6fLcyqsZLL1Dgw1V2EN
zq2InsSln9hAcPqzuG07yh19k4qmQ5/CvpMU/GbbZf99Ki06kT13be4CImXsp6xcBftrkhaqLqSo
M42ai/bXJkwFx19Z19fylHSpGB/4XexiAknjq8QT5cNaGk5+f4YAtVDOMfpr/aPWoH4CY5IojgG3
x+BuqXBLX+QVIdp/KFGktkQ5a1s3zkkx57GDzTqbKyq3pTJFXuH73Gzb6kk4zA6K4ae6xuGzds2N
keNGo17CkAySfB2+1pMBOS5O6T1iUyXZXJ5MVmPXzvNKqyJYwgCt3mvmX8pdRf1CKQE7opaMflgh
ZxgckFFPS8JnC8IZg4IMaZa+kS0ZEXP6AK5VTZpobXXSAOwv0BQ5Wq0LxjF2eENUkQxBgNTb2M91
VJ5j1qxkC5x+SThabU5Z89CLl9ET01DhLzo+iaDf/f4JSH3kKhtHnCG6Cc5qncXewcfrlGTaEFAT
+OqCa6Tf2Tnmaae1YSb0g/QCNP/x0vfup2ysRzdt2bINkUdUnejHWqhl+G6lKVPLscbOPH3uf+Dt
Ra2S5Kre0UZ3q7tT6Qeu4xkGaCU3mzWbCupcnIayRs2HAGKNJI+CkUBerGhWOJzhV30C0eJhNxRE
tNliHaDjeTWBNUyigvLGRotkzzMGt9HtuzGK5QSryZc3HiRR8Jm3Oh9pZ8442YszjSajylMkw8jS
PMY6uPO5xwNsiApR6ubLrr8pe52uyljrSwdaJoF0HEREUOJeXkSiO5vTJfaawMChdxCQeHttdXnp
I3jczjqFnqhWcuGXL7xlRpM4wbsIG9H7cDO8fsWQxtn8gi1S2CeQB8kJsPYZS6YJMvA6QfbUc285
NXWEbgoFnxOGUjLf3v5NhBwO7ylC0tILlFgbmiZMzZfWVQ4johcOsq+rM66LsIDpQ6ux7cCwFlEu
NvCmjQoJ+vyvmCvVMhudgLssDmMyWq/Btc7XqlUny4gqXObTIDGrp2nGkLyDKIke9nXbq8vj3sqM
FOncoW0jG8wnwp/r+p1QCMFuiL7MYnrsGdGLg8dWkGVAHLEU3R488PVerEV37X06vrGpqt0TUQ/t
X7yM88TR62M38/dsqB0rjRBOL3YONx0xncy7brzYki31j/y3CVJZG9dCW8nyOJRyZxu8FTKaqxgw
aHexaXJVQTSgWMM5vWwaoOBp/J1LDYHuVl5mqEEPI2rCqM3k9YKVD/bkyjK4j2DW0a8Ut11Rw54G
FrIaogUNtp9DzAXBx+GgINbW3XzJQMcvYuclU106ql+JggG6niXfHp5mVpFVSxPwJk1r6wNVYBtz
QoQtKWkN4bsJLJclk/k4ANXms4WVBQdScnDs+2wjgCLvBIy48K6prGNTnCgWVgDUes0TakaaFhhb
ft5vikfFLvWeO2U9lop7uyyiN8O4g5L+jzJioFrnBGSmHdKllBZ6yhRTCjix6b+2SkVoXwnHPTAd
q8dPw496jD9HfHhTzrGLP5qbAoyRoY/bdB4DGkDiKnE6SGiH3YvOw2TZRgA2Gqmb85PIGQS0DH5c
MqXclQTOjmqsDIrcwbVOjcuWBpav/T/c04RA+O45T3MhWAUTWLl0xK/m5g1jzLQGWKWMzCHCNeD3
dAXLlvNyTZbYuNxV5eFLN6hxiBZ2VdzJ6j2FzrQqZlsJDYo0g5pkGQ0UswZBHTcBn5y5sPp+y58L
HgneAklPIcwfzPxaF4MlYWuBHbeH11YGeQKFK+SZpN4y2MSUItC9F6cIdPUp+xdfkKu7OJ7yO5Yy
YsXyM0+vY8BYOvMMgp4g9Fcqp6bMESiPOgZ0HuSMh7NQbLhbUctZY92hgVQNFz/FXIhNHceTNd9j
KTPU2zfvkUT9Iwkp7J1UFhLd9aXoeFWCQB0GB9IULpQWw5DzEWXGmoJq4Jr5TBifXD/8zz5uQ4mq
VcT3qrHZtzAuy7FyoKIR2nDbLSTjet162ijpFjlXGkBB9oWT0ZFQjimKTP2cH+hk1Z90P+toB//s
o3rZ3b5SyliIEG+YrFX6KerMwPzjs/LUeZM7rZvl0/yfGVGSQb+a+CvfWwV9+BZO94ENpxVSSGYE
dPxJyNahQHS38hEqKjedjGSDqpaTTDyLJSWvyXT45PZove++C2TYCWq6sN5ScuoEq8vpppP1nEz9
pCnZH0PGiLb+Mf5eIHPCzQ+7sJZiTF7IwphJanePMqymHWQyuB026rCqvQreDre1aT5NVG6vpKiv
s80GAczRTQZBx7ipd0zdvNtKbrr4omjqbUPr0viiqesOS0Lq40yXAy+0YdN7CZrLk847dbBnuRd9
17BrxL4yeHBlECYw/ytX1U3S+2vm+/lVM2pP42x53GalkNuo9l4RL8S458OcZKt32EQp70T27arh
5otE5AT4xS1/R/SSZk9efiOpy0+L5q0g4pEjGNzezXO+FU8p5X0Sy3rw0geodzWGin1uFZ0QQ7G+
YZue3CVpGw70ZIVEoFSJDw5YN7X+eh7KVCBEBCbF5fKWx5f2z66YvYoWidwRnfUSj16niA9iEYUN
43A/MxUAoq0QtDO46432/TNjebYvqbIpc3m1gS78mGS6RVniu3QSWJkfiH6lc2Dn0bTTyD2J8X4v
LOIp8b/q+rtxdST7zpjzIaXn3vrNJEkVLLOKdTHo9ANEgnxgAfhWpd+CSIM+YQQm70E6YCndpfeN
c4+jNPJg1jv11rH6HpItoRfGfggoCKpzrePfSO1m/7IsZA8dK226MlO2ldQ1iEj8Y1jjelf34fTw
jrWQJEtGDtsBklNKCask7u8ae38/+fewbRcoGhddEcI6J9EnUikSNxMvtCjyMG9KSniaT0Z+8zm6
r6IeeG9hcTWzkGvVpdpI9Hovm/+RawYreStZFkWW/eQPX3mjBxft8dvY1nHlVyGU/bnKi9MvibO4
XS7hAxRVc5cCXNjlaIsAqlDVoT1RILI1XnP6nmywNwvXHSL0QLhqRNyBNXRp/kQhSZ92VyvKg1PN
WOUaoAXicpbUgRrDK3BKFnVDLHD90gq6U07CMaovPQPU4/4GjYRYfCRN2l80b5im/9O/lTvqLvoM
sGjpnxsYkRINi9T8EnVV/tjqhk5OPsXSHw0emgXvKYlh6KknGnugf9dlPfhdkG26mHzyhLIqul9J
a+few7nZe2Swh/HtOXdTZRJcyW4VglST70WgbFeGqdJiiBxrrB3ieqcgfEJR4B2iFGMNAYTnksNQ
G49aMmiWXkGJwJXXOeHIOGBE9OfVESm5NyXZePZrr6pN9Hf7jL0yFVU1AGHuFSfvfZN46ruVx2a/
dGxdPbZC3lHwYVFl69JvyqaSG/87MBhSLdI5G9ekgM5KOlndz35805k0OKZ0PLAsLATormNwgjzk
i8QKWQndtxtC8Y/GQGVdE8XbTJJkpNXUxLI5/yQOi9yquHrRdbUSehu6Rjc/YoDv7xoflMDjk1RZ
YuNUTetDaQcVLbX+KVtx8GXb3IM1YAdRegsmx6rh5/oR7cq++Qn2uzmKpGizvjIP9z6XdMxZNBAt
JJOS2zlkHhA50VVoACVS1ht8msQx4/qROu0GxpCHFxXSlqL+jzlQtaPCTzU4X+nUWOL4ZKi939UG
gY6nlFnuPRszdGE7KhGQ3TlTD1e65yzZIHRPTknNIOJDs13v1MOC51tHM2SwJEO5JKFZarRdmDM1
eqkS4Oh45kvJDm6xm8qpeoxXO+dOjX7BlH6yk1kqeG+pw7Z3n9YhMytQfU9+EI+46s28zE0t2+2c
UtmfFbMJaV7PlfWdCEwxgBuG0RyRrxLiJ4RDKgBHxP3RSOqR/tFY/cU08Fn5hANVdR+YFyEYFJLZ
zGwUcR87TXDHCBzOB/JLDhSEAylqEzzpL7RXsJL8Sg8V7sBsfYFMlUO8kN1OXI510P8jIGJ/BP5G
1p7lsoj+lK64L+tr089an6o4S2Czmp+2CBGhNtGvN4eUfOwHgnrG/lyf8fiQ52vY0B7kXkEvjCZ0
AVR3XdGbvgjV7KSs3CKGKau6jfQoZ50FqliALlH0Pg/ANHJJbIAb45oa5wf7GlkST+0ZntFcHpnD
8a5OlY3y0nsa859osli//hwlhou37d5S7GL3TxvNNAKPit0t8CIyErT9SM0xdJG8zGAbFJIKjXEh
zPLSZ2jCakHCaxyRH6GwQZFALGOwu+wfo5pzu2CZYgVmAsNHieW3ZgFpISyb9B0QFZTCYp+wSwci
tfEcu5off070SaxtmvPC7wJT5KUuSDo4DMFY1j/bjPfAIrY+7SAj5sOyH+ExkIALTsFpohLFXjWx
osb7i2n9bbjXes9Gns9IO/CqtnOQ/8Den3b0DuN/OGTQCEWiPvrLBcZ5Irv4+KNRXwmyFNs1vozj
H2TXfXsbOdJ943eATLkjKODs0FyRHdfKHf/5Ik3Ah3ZRsYB/hKn4az82rW365qwxRwyPJtpar6c/
BzJtXhA1wdT86KUcz9GlGuKmoKhrVjwqgZe5807AsSMx6D/2xDBuG4g3R5Qcl4DMI+sMZJ/Z/izA
HKcLi3pmg3rdNe6az3B2vKFVMAq0QMleOxsEIphujIchNFExX/9iHApE7F56PAMzGyOBBLYGSa+z
kig4t7mq/zBaW1fCWRxZVTuoGW7fExjOpwDgWHydLgdKdn5rRkJbkhHh/mwOYuhgaL6odB8EyHQL
SuZQUjOCJiNweHbP29DjntuMaXlLgC0zip8DjDFz89kpQOvXiG09I3shRcOSAUHi+c3a2kIPKFvi
O3eZC0zJksmWNocyJGD6Nzq0Ab6dnUXQdw4WLQcNXxe34T2Qdkiac+v1hL8b42uBh9+ydZz3QmSj
VOlNNG38GNK+hgJc5RwShd3nqDGkcSBNBnuahJVoGnLpSd4Cz07VyeIvSgRKXOiyDmJFbTAqrAyF
7E4pu4/6jGd2jj1zZOVi5chHmkq8S0gfaXdECQvWJ1Y1U72wqrWyzeTDj4hqm3+vR2pp39/V85X7
knQnBYOiuoU/qlApTcADcZGmX3W1oQDSgaLOI1X++mQmeDAbMXZL75ArBIDg6bm16q5qI60IJZOK
qlOKVVF6UBFu7ZMDK1VA7EBrzk+VX0eNBloysSpnr4VhnEWcI+Yei18Y8FLmbkNKZOvEr9XsARYc
AXmolyoDwugoNTnDv7kHcBb5sVNGpNQiMhUFrKFLXrsftG7kbE2YvRKYtueEYTlSSp/9LTM8E1B3
c1v8TorXJ7q/VBEECrueAIB14wB38AsuP1gO34GlYfAg6qKZ0FKW2TSlRYIfMKhrPFMDLaScuthU
ZivAAEtmY7PXSNRMRU1NRmuoWJXC17/T1JxGysPjh6yDZUhYSWcPvrjpvBQQHEHEGzwMS/iIO+ml
AP3evKQEJzRpj6lcGQMcytl2FIZLdaQqCmcAfSnOeRq0HRt9047ylAqXCN6/ZsTDjrdUoDpEXIPM
4UzsavWzvCIH3yuQkJKPGyx1kwQa3yXcb4N6G3AXkPLw7uN6HfL1hKy/J25QTMZmzpCjseOYOUFV
Pljtc651jyHNuk+gSiZsFdXO+t0gwOu/bPDNSFUWCviRhMyCX9miufdIsvDxJj+vKWI11wIcleNJ
4kDzADR9LaP8ocXczwev/zZgQuxdoLCU7V64r4+STKbNT1WxSf606kiQpS7i09Yz8xM8z/p39v7v
QtNgvlXB/36Twt3SQZ+KH6VJKc0G/6azaaKdq4iMySJiBVIcduyosmPZbag8fGI6Si9nfVuvoUgg
+7lHZ6YlJEbYlhPqq+T5J/En3tx7TVrNGJ50T8y4UerL5jk9ZvQn/w7iWTQ1OkODeRzjtJinxYoj
7fzNm1PbclFNfOLingOjd4vhCtfL3B/gJX4IBdzOW99OjwvC1W1oBpGu2YBhdfvXH6VE2IdZWBsk
moyillAobGYfbQgQWQva5eJDuETaLmQlKKrcscvC2a19pWkxwO9teCRA2WMqfcZZsPoizoQa9EiD
fIAl2KufTlRe1ybd8Z4bvv2u3Y6Z7Tx+VliUtUmD/58MkB+A/Lzl34Nwjscr0q+p+YyGleXPz51T
lI4XJpVgEfRwB9m4hkxj05ONPbWzimx2IFt1qm7krz9xJlmBUEnl4n5Kgw5El9G0Cxu0iF295Afu
m6/hch63m2/3xmIIDEnblvwWDCL2ozSmbwIyKeT7SYD1uc0CeUD7ldWl7qTmLRcHqJTSGjo7IeZV
oJB9xRmeZtsisWBAMeSTjqXRNMNIAE0BguM9/ZXXAeeUHq9vlu37D5g8sg+V7V56rw/s6dm15Smo
/l7qq/cU893XFesx9fq21aG/CU9RGXomv+r9X6VdHIHE1C1opzbqmHbbZ4A/jURaS4hLF1lAfCPt
PfJHQhC5/5ptQDsW5links3fQfK3uHR1lZqRoZ8V3IPTyoOkpI0MJ42y7a0NW1eGL2pRdgnH81gb
lFJ/qejAbchdjlwRtrQkFHqNAGcJQH0GKLV6jm405CyadJ/G9XTsjirpVpKYx+nkPOVlrergIxqe
NRIPsL2vmIHahroN9cas0I2NeEgOfA4FFUVCcMS1902+iVPsZIzHuG92r7SJj9E8gzkb+Yh1L2xY
NViPh9GeL937dzGEYclzIf0nya2QjO+J3E0mXjiDd98MpBsSIF558IzJ07mcxYd06BONGEZHOvTU
RJ9ORIYUCn98QEcJYP0bSeMaj+Ad+THaLOV4y1HY6EVPQXyRTgson1qTiAQ0jcf4KoRGRf8Proi3
MuBr6Phz5R/yLa++cUbVvoxNbuNosOK3t/oaFJMjPkGuam2Vd9vkLVwi2xG5j756U6o5MoA0YKzu
b/gLYrBBUQbYeBzGN5UTYi8qFyHBYOkNaV9LCc4HE7+CVHYXDkO9AHFw4aPdnrU9TCyKfMoIDYSF
wqbvua6LhZ1K1JeDLpSfIVs9fav9lk/QAgwti4XoUjzxcA5fq7xJjmhVrfbJI2rHm1yRxJVvjhxk
DkbrMwRNKo3xLtpyrzb5d3MD1p154W8pbdJo0JSlCdaxXyomYvLlamKt/4PzGKFDsE+p9PAHngAS
A5NneB/Q98xRTLt3E4IsGjlKDCurl3jHJJWhUTkerPk/UrcNzrjfZMc8VleMpcNDqi4VxhEvogx7
BznTzieivbKGCtYiM8RqWPxyAgDCmv4qhe85uorO3p+2eBLYn02LyKi8i4VEuyKYz65vJ2ABtkng
daLRkxysi7jcn5dRTgAHSO/PQghIXyxBEbvkUDixauyATYvgZ480DLnpjsUjo8vCj/nIyWDb1bWh
zNYGH2px7IQM2vClHaoEBw1ZyR/GQVxBZFTNKT+cBpcvcjIUOfp9bYSU8A1amO3CXJt+ubkjdtQt
19japhBixzPnfs4DugmEgFkpB0SNmkT2ZWJ8PgqXCDt/0oE/mNjmE78Yl5+kaUO83AxO8v17YqCB
bsYZKFyWCaVd5J1ISlz6y4bevoHfLBzMK5Wa3dIU9NmD/67ZWNCLC3mBsM5Wgwh9/YcV5pDB4NZP
6Glv9dnfYCNwed54w3cRYXEOjJ6myJ4vSFhorgEQPdMDVjTot1La8MUPUX3tOzvfmPkU1xXX7J7u
1W6NYRF1y7bNManFUIhqI5NxxBnxdcaBLyEBeBAub9A6K+33Jvm6A5LxmUF4wSnvmpbijmGK0QOf
JkBVFHDKB+n8nfKQsT7jFFFDuYqE8WFKQZJYxxI2g73E3JC/cG52KCpiw0DQVlFaHIYmDNZBNRSo
ED/YL1BsuBQ+ibAvECRtsdv++rzruRcRJCxhlVtLoV+NOMv9Rk/9tYrV+Osgd86MUbiYR7/+f0Z2
kY1RH/LLFBsio3Ebw8fGPjEN7SWn7htFNnEmNRPYc6Az7fLb8C5fbuS+v+QltJ9mrdeOSnNWkmUR
OQKBtRr5iJUr2lfdcBO4c5rgczLx+2yylS2RuRaC/kFxcMW7KEW/17R3ExvrKEgWJBMZw7q4ckDk
nzu0TqOuMpU9/h5oWOPQvCMLcBiKkVWx7yNIzIUhHyCnLzS2fVRCYt/OiVSktBEcAP0JjwJ1KPli
A38/AyZg68sUOtYArq1pNmiQ2qScgwGONgl9nN5u6muwWWtFNRWgEwIFwIJETNl7EV/WuOYs57/e
OgXtRCel9i8tLuslc70nN04QA0SmSGWRZk2NFwe9mIgoRMq61ILE4TOaizfT08FHg7c6V8BPWxBI
JJ9dSqJvkZbxsS3XTrY/63EP7QNCrxs7r8RzkD4ft+cjbd7f4wucE2QwvMJdoWcvfMKtiMAhnE0A
tTXzwCQrbjyk691JE0fNRxYViXR4JXgsaQf3bkIk/OyEOQnOzi9ugwTC5D0WXDJfNN5vIVUz0+Gb
DJThw267ZqsprTFnTTznVouEwxeaJa70TpY16m+cdnhjN2loEjm6svd9ArzjjpDmJ2SKT0mNYkBi
bP/OUgf5qu7jw6COjM/J/oOj/Z665/vWK2oAUyi2cwlFZ3Tv9yJn7FwkKWspotvN35NGO/kBi0Q/
ADEnkI3jIHBvPm13q5JLFKMLk3S7Ng4cZnMoO1uB5pT7dhvbX2SBOYeilYgtE8f8thxcaIxhekEn
FU8z48ClJYLLf4M9iHNv4OUKYoZkhHcD7ArNxPF1h9UrgMFxjQkGbnVGgPnDTYjMwXtOZOoUuzv0
X1Nq7i/dcvrLAMARyl7zDVLoBBD85ishBqqEmsUTYhzCKz4xsWnZvqtRAwGQtOrpS/l56pCJvC4d
R24BPvw/EtXdyrv+yeaMONNJfmAgqHPnBIq4+ykEHEIDHnL/uOID0SwAM0d7pbshKpvb1H7fsWhW
gC0hGt9OwIYdB2fiAfmtXQtR/Y0asmY8RJtOqNP8miMK+EwAO2GR4uWHaB8cvAoXfl3BstjIr4WN
aMtbN70R5bwg1y81YyHlrWmmaPe9Z8ZSPCTe9TJVK2U0y5k6DFG4xFBGnLR82eKvhM72SRzx5qW5
jDWxTkR4e1XmKjVq4KR9cd3vRk6Vl2jtAFe+UfuKdFe1VMrmuoQOYyqbUCN7ampkPOUE+EQdSzXr
sWgzKdMHhLqrfGhXe5X0aIUTL955yshTPi6JKlKlofiQBqMr5xXZSuYtWr8xYQnsX6OCCzmdimTa
FGFySZ8jeupHElVG2WhreRaCrpCXoNleODp1l9EeKRxt/5pre6Bx0ALYbNcjdKfGsY0XPC+00cwI
H7d2JuClPGJlmzRiXGDiQIMIkXm3MgGw9A0QoqRjjEHG09nZPkpAKhui+lGkrPAJjVEEzNAJwhPL
9I0pdDHu2Nqnza08mR0MPYFRZkmbHCnJsWG8Nsw9KcZI82fMZOobEahca6OpYD3qGeFC2cj6CUuV
lFm//OnsF5CNTS39hRrB0K1Bd1vv860M5g22tuavWRxxisOuRkdXaS/DLX3TVSIaXK0HtRLEeHz+
WX/Gkv3VWhiW2Ua8G1kKA9+ZiBoaQ1MnYusm+3dQqDATgpUSjonJHA5YdPITgwVOtCGHwhXPx9et
gI0P0vslw300MceT9XXKgoan83EWPfBqNYHXKzcGajv2JeJqrLZlb4YKA4+T+Kkt4g48usCxXwG8
dXysC1dvfynTUscvHo2iYw0APPs4XMl1FrJyLqVlNlySQEbDuev3bnCmLSjqcT2uTBrSfRIZ/5sc
QfkupmEQyMxwipH+am61omm0kExDfJzmNR3PA1plyuuzGHl4LwZDjsx+WSWU2lAVlriEb0BTrMsn
lC807cSlyQWvXDkPe74/PwYXzTr7enmSDmXiw/jCj7qh8Ws562duIaMSd9VxVJb/4Bw+E3bYoKEz
xhmvtj/StkBAkLAB1jQ+nnuVZd4QgBNnBWu1SdQN8sCeeNIvIwyh+CrHExeiJMJ4m248iPpxE9/8
lcG58HoWlQIF/WDLJPD1VsFkpY7jtX/LixrL/C6yIKlzxgnCQrknq1wn3+iGy3jqIG8/2OOMlY0H
FR00xzVegwE2lhNDqoy84W4rNtLxYNyFAoCvaRRx3sfVTy5SNJAkYyn0j3xbvJ8CtWPSl8xx64Zw
oHBpzrI5oFH5VQerwayMb9SoPYa1wKVDmvQy5h3UlbXikfFsYWllu1sFx2MIGG2YN1wj/lpcCOWO
1jc+ARDnEJQf+y6qubtxy86LSF+pZO/76sTHhaQRqcNLRiLGRo2Yj+N4hhaPR0BAfNauEwSIVTOp
44amAcBUtj8gQa0ARFT4JAIZEVri21FLClTwRe6kc6+o/W5gmAXR0SFc5c4JgBhwxlQUlbjIpb/s
RcdSH4vxlgk+eYItjEOg3QZDNXsqIEvlNl10l4bMGguDk+RmwZpcqVqUnvxvjXtvKKNX4fkKd3fD
DsJNr5NrBpEBMhLMgE62Cxcl7BjiI8Zdnf15FfsCbrfwLuJn1emSFN5JpmXRuMqkm8vmIJpcDhfy
OBX85JffDS2GT5Ml9uchq6QTQt2nVeyJjF8hWmD7mGz2K3LzvUYlr9KirKOMw1AI7av5jfIahK+2
hsK1ArscSmL1B1pEEYyfq3CFoBs3sYYqxPrT79WNoHJW2MbiO96+MphclHgtHczy9DeTKpJvFjyk
a83c0IXWFK2J79EZKk8z/fgFmQjd7KnD1EYbJHBQafFV/q4GzDUYXSDMSwHxlvQjaVj2KPMOrJMo
ImJZS4pRb1iuL6s4KwKhGsg5N8CtiN0bEeD0U5/cAJ+fqB1jmvWYp8EfaeXP4aH3PsEfYZcsUCl5
8YdLQk62C7L/pRr9VY1DyfgBmqqf1QNKX7iZkTiUa1CRNfSQ6Zgk/IioKXniDbmh4EBD/gBZMv0U
lvmwJGxF2BWeuB/mxOJ6MaAniI46oJxHiqNW8UwjGxhr0ShemJFinF8gWNl2PztkRVI5LB6XLsUm
wTl/AFYE4sb0MNaRUnGyroiGcFoSzspXTX6HDZor0KvT8Ls9xPnvoW23T2ab12lEheHI0VjqtOge
Gnsz0pIGWeWElefEzzhlYCm0yvxMmSgT9CheLZ7kZH6Q1h70ODT0COUL9BSbzOs1YC9FEGWNWHu4
90pKskNGWtxGZHLegN1DnkelUDEydZ/dxD4fnsgTCW7+XOytlg74VZtWM171Q61qrTu/Gw7Jq/Y4
yqTGkIVofrY6TR3tA0vb7Oquciv5EWW9LY79KGSvkpbKSkbk5p3i3ILKIsWUShg3IJCeq/yjEHy3
90S5298/toXGMsQtKI1z9WRo4fbEnp527yWPyD/v4pbx851VoqiAILSD5NQLCfq21A3JSpyNnTSl
gYIrbzS+AVm8T92LXUg/hR/6TE5i00ZXbVYtfIsdccUZqIcp+li0NOsD9FK5J59+iV1zUQX219cu
SYBLgUVAT+O7NguupKWXSw+LLhGj9Es1t73GwtMaS3mZsXXVLztLlQDb9C5unTs0R+j0Arz5Az6i
79JPkPO68pqDD7doBpEvFwZy5rZMXjbaF7RhfqwQvlCQynJIVIuzB+9M5glZucxoXNOst+ZtXM1C
6vlaowGMdd7/DzI7gqJGONXyv0haVT9IuqwziBFUMZB+jEEb0rw8Z2ca2AicOL0wc+eEgMj28IpE
hayJw9wBGsTBFFKaRScOTpJgdse6ZfR4HC5KBl+Sq9/XAotloJt8+i3IkZWTwGXO4GjsyZaZA3zV
HuFjWQ2kzafor9IsM56hMbNM5GquW9PrKo8aQj2h2rRoVJZ8MxX98BI2iB8MNkODeYCJ/c/ERdyj
O6nqxWJdIXWOdVFYFUSx4UTIEAI3OPAbVLOS91Fj+ezYQljWGHLyr/EsOeJiAtiwjeJHmdQkyI7p
NOvTEyJ8NzJ31zheuup2rdh+BPWTuoVHhiEm8U2j7pTb2l2fxVKzWbZamF/6DVDzOo5whVzH5+L4
MA+T/dA4k/CxlNgwzC7FBctX32JLNtiH5Pec9kuxlLcW2zc9uLw/9+EwxdeywVuFJ0oHTKilv9RS
ATrFAoxrYPybsxwZUczJAA5PLth6BN7wYMAOJKHTHA7OAlQJ3/ORJnvBQLmHPnB7fYvymAhUweEo
phBrfzrIiMWg5Yp6eCz4GFZ6pNljZZiuJeE2DfL+UG5rExUNosJevDBA4rYiyS8eo+l8fkN9EuIn
7FkisETvI0rg5utGUUcuv92zk7ub4CFURmY99LkIdpKdNz8FE6O+1NS7EDFwAACMiCn2Pyy5jrnn
enlsgl/SiBD9fSQSnTAyelPa0SzKyusU0+WmXDUJ/MF2TOjIk6mrF3vzsXZhGU+i1rw27C+iGBc8
t03YweukD8WnICtNhB5Ssw28o8IaJ99jBvJU/ymDDnxKls7/QqlFUk8SsL+9FX6tgGwg2/vQePmQ
/R5qklUPRyFLbL1z2pAFt1Ah8vdCdl7YOaS2eBsdO13JaOdSPHPUR/nhfHj6eUyFQAetPYM2zUvM
4x/kSZ4OOPJQ/GU3J1fNortFKYUxHHxGfAHYNY9lWLbz6+q3+l1Kd2SyQSKqIXEoLEODIzRyhepx
Wm1euQB38wm2Nah4GUCLh98glK0Xeez4x6PlKhE7oh8WwVSABpTeuITvgsA5E0O9OUNYysGonw9x
HwomF1Opg6SZuVG10Wu8Q9KWayO0Fn8ESiPGoaUSECJNk0oCYYnsdj5Rizay/OKSgLBsAui8CnqG
Rsy0MIAVEfDT6U/RqXK1jwuMAGivyrHgtkwdkl1Ak5OHH1AmY2V9QLbNUtXz308AEaqoGJE8Uc7O
zBDWLCU2MjRzuFByjXBVV/1bSSZtPmgNcXyIJxWe+PHfqkbmTYpT9ohNYJw/mNmEhO1zHhOD129I
dPa7ahpc9s8buof91wPdDpwvz2cVJBCO4ihZtc/8k5idTnvn2m4QMvOFGR3FgUD8HHzzQJw+X4k2
0R9OO4wSC7tB+QBU76+8ehbaZYDwhG1Sq5bDz1mcFo7SfxIW4XxQm5zds/FTNEdBHhKqOy+AKPpu
RUHN+BA7UdWhnebBB+Lql32f66ReybHWErMyRPzIbKRxys2IOBYNeCZWOcfXFUVmSLS9QSwo11D2
4tY4ic2sXK2jkJbjINGh6sdIJiai3Da87kSGgXPlzYKCFyDcnUVJ42+ALj8qVZTW0y2HsQshjZEL
wdQE1l0hzLChOw2zZAu1hFDwRXbbHWofHMh03AP3OAS5O+Z8mg4tXLonf8ad0LGCW0kkc8rDdlp/
ms/pdV/epqAO/WJ2es7smMU05WQIgO7sR/1VxOAJAbg1+yXgmBf90DTfFjE+wvoevY9urjfGkTBA
uzXDEDfYUnc+zJUOdslZYQlu56yUyD23ug8id++PF7efD7JG8dpq/pbNb0+cUtwxiC4qhDQZOYZv
MDpRTnNbfRsEwHo6RESC9xmoKbL/oJCh3t+uSUXpjp8HmUA80OzPE7D8OFLJaDv9QEpPOyWCEDDD
ZiuEHekNX+Qj6RBy2F6zjmEvygorQDyxNfcqZgEGiptkzJ1lC1F/kryWrOStZDeqn0SJHWi+uMNd
xV4lqo704VL/KZvR6ijDK6r1G2i9gWsOu1Wyw5scsefykKPecpq5KOVW9bohcPclYnlzWs9Vaj1x
UEoRhzkPX+aw8PayrHHgfCrTiJePiFWsiQ0fHJD1LtqBW7QD94JTD551560VlvY7TIeuSOO4TfbW
LghapIvqwvv4O7ntf/+0f8wIvTu/ByCXR9bRb9idZsSyYM3nnXCH0H/7M4zgBroqOorTRkhM3QQ6
1Jom0rRAkAz0DQ2T+8ztsCpSB9nyj8tWiCjAKKP3G1nFQpQ5+exzZkkCTEwyroKcPmc0L6cMQp4+
UZQN6XygnhfYtn5d4+yfHudfXyM3jivLlqQBGRSKel8O9zu41tA/OZ9wKYjHTMwCKqxJ1pviskVG
6E87DHqlxn4Ile1kKaRWTVDcCp2BuBLqbcCt8WwvRTnX12GfG1kdNLMF+e1Wc58e0LpkypAWkgtu
pPY30uRlUK7qYrnX0A59vnLzF2zeoTbF3edf2rOJIGtPH/Uk1dueHQDx6pR63eLXuOhVOVUw1mMI
Cn+cozjnt0ccQSpCq051cbFW7OzuaVu1RYukNyrrRNuTkZYJuPKAkdJMv2pvmOiZSIgar/DIsXWq
TOKB/v0FVbZqRXAzszfvBUpfLBZcQKIV7rDBxQ7DJinmZ+QHRWEhBteOeVFlSot9YOLrcJeZZVyf
RBRiGkPn0oXiD58d67bjhcO4bvYW740HziVYdIpS/XvB6+lLKyBfd7FeOFKSvOfLyCayE1W5oa6Q
JzDNdpfm+smVyp1cLKQnrpANhYewogrqKXLem6G7nFmbdV4dPlcMBCkXNxwSnWLOXCk7HRUHAxqP
bCSGtwKmj5Sj9ui7PQnVCwYjA63aUcXlwHZsqU/iikLrhVpzCuxfeOyS0mgcNKuNkzdB07090mS1
Zn5KoijoTZfRYcHnccjJeFOmHEaLPlnVBG3pMV/AsLLgzMVVA4r4mfgdS6juzyy85316eV93FapZ
jswH7OQktV4Jk5HQPKNAx/4kc9DnXX0sbHbhTgI7EMJ//rLLLG24NNoTpxlFFZ3V9g3p2kre3ApZ
K8CcE4hZb61xo1XHsQxAV9+zGEu6J5W6wKCS3GV/ecVEa7A9LzF5Vq/i1+utZmkeVOysnPbRQnHv
ihSrvUIUHxYIsrfm7XfDvxQhVwKCbe4GtnmaHIQbOeFrkvxyl7zOxA/SgTfK0ceQLpww6/XSyVA1
x4+/EUVg6Z8pvO+Dw/sCpgLMsOaTJppojA6bful7igocoNFV20RkptUdvwGSQiqnDDVNBpvD1EkJ
UizNLcPu6cEryIQSxE/48GMQjAT5Pixg8kQXmcDEXTgo6trzoeiabHdk4hYd7N9/dFOBieAmlbfj
/rcts02lSziIxxXIctq/KGOlERFGXy8Ui5aynzGIJQyJnqyXJong135MmN3oD6X6GwpBKChC26Zu
ETHXyMSj+hSEE99msXzYo6CqHPeLO9VNu27L84vKsiBmlzJDH5tNIEgwxsxt8t4AgNhJ+mocqlb/
ahZrxMfzVbfXhQ1pBsb1eq4duYMcUtSFljVm476AlBsPJFnOhQcfRwnF4/20OUauhdVrfCgxir4y
sLctnjllWdL8Fk+khJfV2/Fyrfnfi+elJ78zFvm9YRVFSPJ/pZc6zHHcXZGMSneu+BRK6MBzUyFp
Wqkd33oJyFLrTKiIG/UyUgVHAnjzKSpn+giGwsA11ivcCInZdNcmnETaS9GcqIjrdSKLWsJ9QN09
b2g5daTNELaNFqVJkleHyTfcOVYfOwWg1h58G31F6hCmoSDoZuy/bYBINMl186+O+hNRcNw7HEeG
BGVVdr7n74MY2mOakNv4dVQf9KkE8GIoKgw7EldrdfkT7oWSVXnfGpZZ4MMqCs41TG5yf473duH7
yF7LaXTSZsZUGS7Y8TEnUdxnQdIC3ZrEIX1t6ie/HlC3iRz/dx5RZR9xY0fQh4bAUqWFIAjnerRS
I6MELBjO7EkUaUWkTIdAapB4msPrWiIekgOacBDdzfMyeBhokF8UBvIkNtYnAXxlLvt1xc329TBI
6zpHMydRirAxpGGQfBQcCKCO9oejN8v3V0Hw+TrkjIxL7BH5zM8ccMRlpDEYc7qUhwORd+POTrb2
wZ7jYXxY0eNNd3HzmjfTxLGEwi/VZyI2mJYTaTFLpge4b/GI3lbK4Q8zoUQd6o6XUJXzmRRU0inH
cgjkjvQDFTKKSwMib06hwGkT5jlxDj7gHUvpysPmeuQsp/XwD8NP6Pkfz6SdWe1CSKqXa6o2E07v
vQ/jpswVDgviK3LwbRlDoKci1FMH/5Zq0tON6lKyRhsqD7TJbjuAv7k++Yz8gB6CY8UzrCYDzuxa
hN6UKPiBbIpbASWVSk0oNi5mhGCUA+U7kCRta0O974UwEVK8hVT29ChfBsLgNyGi682t0SfQMIOF
+MoNhsTKdQuc+q3lxm7hh5jQIJ0FDvVNYJHLi24IDPZ+x7oxLnnSfHiKbm8mZn32jSYtIfFfUALc
HQ0sipGo6MJs5oniV9J2iGd7cMVs2Me9WcNt37HsRa2LdMQtHL5+KqR5uz7oB1yx78t3cE5Wjz6x
hhnmsdKe28aXUb0XrSBtdDhh92ZzVaAsEcybJRE/MhPfzGM2e0zw3yGyioaNXVKPb3w1E+OWpUdI
vW8YUwQkOVbD7zaSjvLxqYGFamDGUkAozpMJeRpFGPMMx7CTWqowu+RsQvLZPYTZRcxg3JCAJ694
jsxcU5gmJ5tSGPMfD75WT1zgnfdgCUOpE5RLRmOlo7tbR/pXt+Vy8dP/Y2pJKPv5Zkrf5B3pGkH5
2XEwLP3AIrlPzOOmAJ1uxSWaoRkyk7aqUvV71ZNbDIA/PHw7JGOlHkQUoTOy+B1pKOBrvciLY7Mw
1UH6+3mlZrF/quvS3pN1OFLvMTXmgqZ+xaApzjWvUEVMtsK62z4/AL0ZCjAuyNWs34JJu42PU9Qb
oISTr5GP30beOCUlZOM8v0KV+NFXtOBgDdn5KWtHBEcOl+2Lx+UHkb55YUqdLMuJgZ+hsWJOrHqj
+EfQpS2i80vU/oute2eASaVyOEo4/L8lAh9xr/RO8tO3mBGEoy46LwskwdrxjMXoxJVKv2aBNIlx
bnNPEKIm1nCESucJdEniExS2xBLp8AdEukm+ml2hE8ZQYc3kMFRSw+pA26O1bnfDGyxBBmM0hZzI
gDDEpDOTgV8w7m4jc0YIDTI7STA8oS0uZJZV0KM2bJOa/kB0DVxT2sFCKbn+LCHupPQzEnXn6N9N
NQ8ZMQgmsa4Ibx+8DOqKcXT4L90XZG83p345kFutrsDc4foxsU9um08uY9KECjdK1w29o97URe2R
gYk8jIiz1nSRK2AFyyfqHt9rOWMfSVpBMdme9WOnt9fyJRC6Yt8eTjwf6+rmtJpxZxwunFofRo4w
UXh8OnmCcpkfiwiwri4lWwLUy4Hl01NXON+6EbDkJYJYMau5fp/aOw5HnpZIxOYH4jrqHR6LXDNv
D0wGdKVBpStNc38jORRNTpzyn/JsyvH8osm4DYwbIiO5gcvBM86dXgBuYawa1vST8fBWG+rPOdB1
mZOH8N74BWoB08llmb5nBCuHcYsK74PsJ0K1oOhfgl3QwWPn0TqLLi607iMbh7HDr0fWJLmHqLlc
j2qVwleRDrYjqoFMs/BWkbX0z6+Yq/XTQd+TjgdVSXu6yTurxqGiEjt2Q7UFOG1N9M7+XnIUDCWs
xboTLNwlPNPgcaIiv0lx0yomAFaH0jWRFeAEkLatK+mT4Uc2AvscSP++IEirT/Peqzf9Kr9P2RiP
iOyvIuazVLOT2CgXNaj4c+MxKYF+Bs+nGT/78xd0kDaSfodWBrybzKLs/yqyug9Bqai9yemAGW1+
6+fHiPW9sLJC8sOI+J4V3Ip5YZIMLu/l2tOUitaSpb6QRJD6B6Uj0Ltb6L9qk3ZlHKitkl6r57Hc
U9tPeX8cZePrBishd4O27+2CwXiwMiKSOvhb1KzV0gL7EA6PVkSqVGIspdIebL1iBr6e/b8lDrIO
GZWIu7WmakqbxRDiW/yrZfpioqa3YMClGBINywgzaBoM3ubZHD8PyQT4qX4HtOZt16TlKxCVsU19
6H0oPe98UgYMFw7RqIxmaqThTQEgBVF1KZdDZfPJz6YE+6sgrwQrKo4ApxzqW+QpHOhOSOn15LRt
i5pEjUBYSFXk81lLj0w9eUxMau5yLipbkkbtWu6tWftRrs5kePiBA3GbOOP2cYUJsYinh9wlQHHU
o7nFTxih0TEg8EYQgukhY9WBJxDio2JynFwSph4A/a2GDMg/o/zGAwmFJn7cHUuST5NQrIlt0/fF
9hSQQ4GWSh3AFCvW9vLYc5HkYjGFN4FAnoLuLaEtz/s6Dv/I7wQmwkXy3rsfI5qwER0sGvMSZg5c
ffkZv2V+/7Nt7/fus38xoeuup2eDnmRtA01fLUe5eNCLVx0x+fhr3kKry2LY7THn4jjsQlXLDviF
LqEqNxMDtyk9lGFSAnlBMRNFuDEJyWCX+XWDgxZsiPeDhJufilTM548CXDJD+MmOqpnvo/t0aQ7g
RVzg8c/jmWCMpr4a2Hs6f07L5qLzF9HExqCy2WUk52nj/147dXufszDNXBb/k2tplQ6pcn4S2U7z
zRALweS+iaexupvj8E0hdnJqH6THE/5hhzMN+NgJB1oCmLT81Jm57G7NnEbaibNlAeLb3EydOsTf
u70+mMcqeCv/e86GLJ9TVyEB6MqG6BKOMbUcsn28E3hN90VUt30j3o+sTUX7TnlNnuOAMG4jUeYr
/WArDIH+ZkkxrkMBCRWsEXX4bhPWFqscpxGMA3XxnG0rT9vQl3/2OA3FJzCGH2YEWUmerkXa5HI9
+/9QsVABq3VHlfC5S/LsY9wQ/PgcgmKhNA3UqL8wHl0FrNdnPW07vD4nvzirNsmHh3UHPKj3ZlxO
Zk7sgrEH0+K0gueeEoehJ0wUBK52TIWZhLRgTyrobugB63M6FnpjdIKzynpLNC8BWuKQHAwZLIIP
3gdF5kP+FUrxDIB+TDFjW8aZbqFy5+Ss5CCUG+04RCYRel4bVWRGSRDv31wJEN4fD2RpzYblHkgv
PjEZNnFYoxMleFU0L1gT0uQivqWyEjDpDL/tGeXBXeKUEbQLzDujqFCPBxUmi82E4Hr3ZghEoPJm
rjgWLd/vbtBD62vd4kuOjw0+jh/xI7WWpidyII5u6TDgRnxNSY9E4BKJ8Q7Ukc3Gkk7CiIFUGYwS
RviEJWdN97b98ArqJOeeDbq9rypLoP+zhyM5R44wM8sn27HlVcWJmaqcayzQBVvZSJFv8/jBEsQl
3i14HxPg8WKD4h0J5wBseRoSb5Jc4+aVx7HwqeQZ4JYCbOVyrfnsTB+TmCbf7b4f8Il9SI8fX0ns
LA92AmWRNhUuPYJ5kAlfm7MZxcUmw56C92Tf+oqWiGP7vtlQ7BI6LKZorKXifUMstwDIKBFawq++
WWEWfZIM7UOzc32pcU1nZAey7+GAahYEgA76BUumwYWE1x+F0nNqExTBSXzGwAHGoOhvNvfWJgWa
+wdmXN5/EtGbMirAouVvT7pjYcnDxiNr+Zeg92eegZvbZqrNHB6MrUTYSH6fTap/Nrr/XyU9GC9I
D817WGGLeyLTud6WU+DYVosyauOi3TpSPGa4I5+pSt9VLUTsO/RYXa60DjUTYz8bqfarr91A1ItL
urV78A8Cz2OSfw2MbKaJKORDGRhlZQe+70XALUkgE7f5nklbxj4iRXmAezGuDz7dUf9rvyVVqzQe
X1LaDGhJ8yLkUcqRAXqsgBSmp0MCg19eiybixVngsUkQUdA+vRQoEPxJG8zjDhQATsQrN8nkDXBK
VSVWtuGrB+pHhwm3TY2oj60qLesmNVi+/Xzg8+gX2slHS389DQgn2wOxkEcDt1y77v4avpcf1zEv
53uL9WtMnGOCebD0I9HGgrM5vz9a8RDrAOJmyf47a2Q1gpeR2Fu6i8xzxhQcagRUKx/Cft95SAA5
R/8dtABAlpzqfYywEQLuD8SBu7YJmN0Gf+fF9CTV28NEwZy3LoXadYHr6xIbZVqXdyrZ0y6GGDZ9
p/t/NBIQUcCqsLr7EfXSy6aBNGN79shEwIgHoEGi+INqLn+g7TY3fFI9wdNRIZHQcgV+WcWvgGOb
relCkHJsuPBwklHAuHCJUbZV0f7woVqbNMF5cq6IA4WMUXgprWslz8YHf4xAPLTFhuvPSO1D5iRP
bPqWpKSZoYyCUrcsyMEhIKVoqqvC3fZcP6fHUClw7N8+RN2Oe/+OeMEgiZBlfgsocI5dcDpZd1UJ
IxetH+HCYiJmKiCxbrk3TfFOfuj6lk1UUYKIcedLhkvZkTV4M5ME/DOUTbzKv6uDPJe4OaJMIJIv
oQ0xrxFaPrXBN1tPbag9Hhtr6BLum1F9i1UYamIAYvFq96dcIfo3no52wIqUL6ySTDxwd//uTyX5
Fxp+Lh8UdWpGPucA0U+b1JwxAVHCtv9DdQ2oq3QqgHfEnBH3e9ACwwah3Fp9mcQkE3hhlZUrADnu
qRkblCxYp65C62FKmgnGgVI7PNaJcR6nfY3vX85cDkI0n3kErQ/8ufcgQdiDLgh35Dch0A2Xfc1n
ixDF5hW8kXXjcQKPPkBxAxaOekQLrWOImjZTA6o+SZaiWwFR8w7thOG8mHAQfxzRiSL9gAJ4pM5V
3xwL8rpSmRNICVK9p54iQUc46IE3T7ztO5GHgXBA0W+5qftyEwNqhCpVP0ltmgIwYWvdb4BG6pQo
b7N2Qr0HJIfjw8dGLGB2pAU/hSUee8yRdavVhV9m41xF2OdTZR2sERMvahVhtekSIiODcWAb5weB
V3rpz9yX+1gKN1WAcQme+SyKiXqXblymxnF8JQieNE7zAhlJXiJlSj1wos3gJ19uu3A0ArOR4t4Y
MMgF5sCKgOExV+ZSx53U0twbZvLf7VarMSlwdBL2YL/YSlkez92jQa92VYHid2SzA8bJ6TkUFiGo
DX0yt4GAcUJ8xynYQi4IbiNE6Gu9y5fKT+7NUGP6ivoZ/UQgGO5MR7isKHyMM/qXVcE0w8SEBRC2
eZ37mbXDk/Hi+gOY8R9hW2w96CG2LIXQb1yQTTl9Lo73utYlo7wOzWK8bCg+ZZbZef1bvJHNZhEC
j45L3qcEeLPbfdBBrZa7b1rV/zI77bfbaHzJR6rHVRHd9DBH7OR9CEzzxgs/od+4Dact+2G/fGLj
4KI/BQN6lkScJ+cM3sQKLiORAWidbM18/kS7cxd+asCLx/Vl0quJS9ZgJ1F/Mt6BsmxfbIXtSNY6
oKONMgpt3mi7wgRZ0oqGlIrUFqV8WUAMh3Nhg6VQcMia7gz4K0np9gFsZOf/FtMaWrfaxbKxVcR7
pBg37Hz788TWvktZrebZzPdfZHH/3L9v7bNK0PMyPW8P8DRSvTAKGBhyJjgPkFKTPQKGbVkyykJb
92sMCFpyOa+mZm6MO2Mnk4gj9LQ0VeOImVcwXdWNwEm1qb9aW9dMRvsBlBvwfH4XC/YRVlyIr3Tr
LAGMH4V9pLhwpee/R9Eh8LkfMDse3hZ7HC40wiwlhGM1IDYJuNcnk2dSNbFOGfmr+36JVtcieZee
l4VlrPqxY1jAdyDiBDaOnS1sNhJw9t4pRxsK+BpjsCBBVG5Eq53yR9NUBmBaK09gDNuqCm7C2A+P
xfDQXx0uoqiKLudvrAtUO2eWrZ/Y8vbRlEUFDq2sAKICaCWVj00fMcQFf2SKW8sNF+Rc8gCD9R5g
Piti3IrXPXQqTvVWQZKzq+Bv6Lj78DZDol8ZAE3RnBY9KIOlXycRjOkm5X9iVlX4nQ9V1tTN7l83
wNg/pIzexN4q83ieEGZbbClxvG9MJIesF8dDzDD4qLWeeN80BbdMnZGj1wuhrGivmChBLzIymDRV
+71b8RE16SVc225FR8rFtOnOanITL32X5Lb8/ZEmHvKWvhrQ69ZegTXMX3YlxO+9te3HMnF4BrDA
Qt67AzD4bmtUEv4u3c7uAz3T8ow1WCu4AIY5p8lPwTK7dzFg08Gk+/SV4cXTYL4Gc+mytNwunOEF
caKnMP3JHwoy4i7ZWPMhtWn8zNg4kDDy/PxMafLZUnkg7Al565pwUQ9nS0d0uGMYY8GGBJA/8H1q
PcYzghTyoFdQtbAcSnzPM3nbI2DvkF1/m2vHL/t3KLHxnLtaZH8iMMRZh/pcMPzYQSArXSP2vp9z
g+D8beTGeZqFdhfAFiDp0SfDK/BsrW7cYfK3Xzc4Zpb40KMXFOZKH78UmJU8d7RVF5qZ5EhI77Zz
xBrSEptFOwH0oQPjtfa+MYxt+LgmfwcJGPoC5CPrG8BX2e/2W3T6aNBwAJ3eO5jyA0Sz8gUeQg7G
iemEpj2J0dL0C0OfFMFZwOv3D1yT/3lg7u81My5C7zqQbqz8IaR6hOGnUDiD19FxNBvzA4XtPHFk
NFzmCSBGwFp8dwUXuKWYc3rm3PkGP9zgS4B4oHOp2YR2ZDBjC3qY1SxAszClG/HZXJYsYfy0Ya4O
cHD+iirbpDuVzEAQMFL7V3DBXFbw9bDZqerm3OHF7O/jXyU6/cqghK5z8bLIKbs5xDGujfklPH3S
iG2u464pWIr4byjoM2TxJmd1Bx1FxP6oavgwqHchss2OEU4YmfCFlWpsFoSk1JkaTJhwj//k1cp2
2YMHWqrOVLresJSQLXwG7U5WyyheLvcNrs/hqfOpX56lz+73xKGj1GVf7SeaXmz/aDcgIFwxjR1/
lJ6iJrSR0v0rOjdBUU3Iq/O7xZMJtg7EYQcabbIHTqmcxhQEKFlNacwHReubMbpvxZ6/rqaM3LhI
fzSi123TZ+ScFH23WWwe0M8lNbnACz3WKSXJUaJyQz6qH5epjdKi348Ovlbrn7n84yyjJ/8fpnch
8OCFnIUdHloFiXTCpwVdnV7P/uH7BMRPhX+tvSa+ZY7x8j5qoimHq6mq6LExkW2W2to9PuTiYS4f
fw37Vg5pQtN0sR+haewGcbT/zl7uwr+mEV1wVBQdU9me5vxF2M3cDQqLo5Hk2w8yudoZf9lhW8m9
CCwhkeypz0WaJsxf0/1h6/FtR2dOHG+vmodMc57mQHSMYzLAtFz79zySpTfmwkLLpEaua/YyzCKs
kWJEqj5P5jkDpasTWcxHAL97BlwXzW8bPurTmJuy9Un4zlLYn/cUPT4DXeOnJUsDeTBs421b9cL+
wzz1N3tYOmkC+ohFJc5EAKOoJjUzFgK9nIAWneCZgGFaz+A4wSeV+AT6Kz/Igmop2DorM02D/2qb
j9884v5p5zGHeYLVRGvcN8M+AxlGJUyLcHZmimfsyQfEByHHQtmYiJj+mskWbpbGyQ9YlSyzHpm4
APA0TX7QAb903atwX7Sgvil5iTY0BkIDB2WsYN3wqMskzSov2in08KWeICphHEx8Fs3biZ3OLKB4
cEdb8xDP0ej7BfSY9iDYJfSdUyb2FSmppqQ2BUD81vnWOW6gV+epl0yTIlqOnhLVbK8J9t5/4VYP
s0Kv+pZ4wgrWsA0l39zuTAI9i1CeR20L+k9OgDfCLP1b8UwaU7/+9LltX+J+ruFa2piIgHcsy5Mr
adpWRt3ZrxWKC8+S+g2w/4CrcuuRAC5jSuLYnp8Q1MVCb7bEnC9WCBhLtOZF9oUlQOyQJBrZhs/P
o7H91JY0iNhjaJh69GIRj594VXGU1RVBBE9Obo5RUE9M0kGWxCjr+EiUfZ3pzzS+0e31Aaq9Tpt2
MS35bBmcxybgXzKvYrf80Z28oJ+oSaPFwyH1Ic1I67ksplzWMj4gcUCG0jDXCfT1xB8kBRbWwRA8
RZStnJ34FpHYpmCCr/bwIhMaCFMMPv/WcYYZSgnxrmwpje0ea57jYE17y2mPyloXX96ivoCa2Di7
6Re0diwSZXvUP4nR947DPR7uHtR7rQqVxNn8l6TPZoLNSvObKwknoOvmgRZpZeHKsp4ELImtF9GK
9QsAN9fwbLdj26N+IMZv3vBoKPBiGK7rezdkgdNA7ujk/8YLAtNnygph3H3wcLlBAM6jJCktTfwy
Z+0NlL7edgOBMQF5chIm5U1e//F28gsBRFv4O/u4pTurf0e5HXK7/bULsifh6TBDqqn3eVzldTZM
l2ZFH3cNBU+R7HWYHfQr8olZ1KaGTsnGSx7EhCNlOAlqRipaJN+xFeaEBFrhLPApmRTvIg/xDcIJ
K1Dk/lFgA0ZtJE5aNgFvfCPmzfnHmdA9daue7HzUKdqdXYv4bO/yMUuOWnhNITdFeF2GhwF8br4d
q/kXt0Wh7qCOyU4mk0u+aPbtoXuEwkrVJskYY2Iy98ZUg5f7+2hDx63yJQF6MHdLlQLfZ6UoYfUm
Nl7EKC/3MNTDoJmmmf+YqDr1ywTD9+Ka4BTS6uajKgmvGdh95RE5dgcEKl0C58OiZQYUvUzysIMC
04b1zsmTUptP9W/J27yhGmDNE2fyRS1dyXMJ13dvNymuv9akVyDDsSrqr8adHdke878kK7ND1iJf
579c8sZlFO7rQHA8toWUEgI0Utt4UTfPuXKw4fmCRTJBkz83Z7Oqcl+rJNYe6JycfYk/OvsIZihE
W37H+WCIHJil5Kshf58q8oEVG9ULSrGHVb4pL+811Ny2R9SM34XpUWQYKoMZNx06dtvFZz54QYg0
eMBJ1a6jCxZ/atQFXnFZvhtlgepRgp2B5aW8HvMEyBHfm1M3xUmKFLHwrb4i7uSLAK21N2kDwihG
T+9f/YRVGDEhB2YObGkAvOjgiqntqQtwWxBWWHQ8+bGUeSNdPhWFRl/r7/GLtLOTsZLkX5QSiu69
1prB8xJPl/Lf575lqmiGf3Hdck1EHN5bzr7RxWbWOshbLfYM2YNwfZ+t/ZigIqD7mrmHoG2DGTHk
BZhKlr31pQvTWShYAwkcpYMeie/3+d9jqpfBvpDj9Dyswidjew1KuI5xbzopYd6I8UDlfVgDcHZ6
8Z1Vayb4RxyHALajHTL6MCtpe6NkRwq5/+F5nTCQmZoMleUv+AzzuuVmVcivMAIl2mrFe0h/cx8s
r94i85RkjalZwvSxJeyVwp3dhLXRhfeRhzyfodxzNU+Wj8cbo/cL7SGhpD6GJ6XXs7O6glAnJNpE
75hxY7fwC8xnlqVPUkVwQErHHXBNe+C4ovcHwzlqpqNwMRT9I2dfiyFfSt1UdDKy3xlVG24tUXqj
qTRJ+6nfHPdRwEiV0S4D95h4X4g5vqJpu4C4zELtoWWMeco2A5ml1GbMcVVHQP4zge+5vwybMvWr
4nCtH0opiGgAPctmmDKxzFWC5nZktbFlsPN4tZCBdqA/zHyjxrWKWpC9JP1pDUpxGtax5zv2tN1V
EiWkEpg0MfRnXw1fwLvmpg64Lwk+husOOpnvo1WhDmICELQp8PnqiEajx5cei6WCafPEjuIfGaWf
Bf5d8dOuYJXfsxDLc0isgBcbZQ0Qm7tw1+rdfQF7xKeMqxGV269tLTgSr2r6Wxkeif2z6VBOWuaA
YnHF50jAbc9UsNbSqBVwUfi9AN3TJGKT+kt0/6g82Q4tQh/ThEpqt/WYLuyVWp39DQdHUE19I0jg
i6Bj8yLOWKRZDGAshjEaZaTqmyldeZP7TvQG4aXNBewWhF4G9x9Fqg8W3LanweeCrAEQ8SoplHt1
ATlL4E7asSBcMGeektcwi+JeSekfId0urPaoUHcsHgMQXpSTkSMCowEbjZ2OoenK6psIFJ5/FLmi
HnqS4PjIFvA66uzaJXuibnPUPTYN7RDXfiBmeMb76wG2XvyxYHGizvbB9Yk0ao8rwzg2h6k+G1JC
V6A3goUcV8Q0tGMMD1v6/pIg7592ICfP8YdevQM2rvMlrXBgTU/wK4qEMFv1wYIjPEjCpNf9TDaU
SRJuA4Qw8/G0dslTDu42kSCAkokyiPxO+q8tkDBtYX0B3uy+nFbuThS/QxW61j/68p89IKDFI0Hr
SZjjtu9lJX9F+T1a+c7UxUgNF2p+w/C0pXFpoId2D8134BGrinCMEcG8bKMnjIAghHLMa5pq019N
XYkIcD9yoUyo7YAuCLmLDlIK+cBNx8uY9yXelV4+DFBLW9j9pi/+8W8JwpJ50qs/9pz0RpHm4V+s
RxESojLDKCtCxB/I71imRx2u5KgpUlsyza//e5PSsvgfdStUictUeVz7Nz7GZzxPr+hUWYc2HCAK
lslCmbcv6i6LQLD4A33kGl2l/7r0fof5RVHr5/T4EPBBhGwoQiD2nCzV7Z8b5Su4T2rlT2pAR79u
yvgMibNS7DTQLbQaBciEZvDTN0SIxD5Y9vaCPcV8jko52LlI7EwUR1XJshKfepbb7zEFk+6ePOIT
1Dhnz2p3P3w1auLMd2uHKa/JSvW26hd7F3SXkALxw5aP0TYXy5VPcRX44ma6I9P6lSaEplyiMYsq
Yh9nK53dBJoy9uewi6Gn+R+XFHJ5fFYb74nXn52tELfHHK3X9sebN/v1E+DWANwWIYXmztocExrn
EBdYT0oNPC/+YaKrzYEBsrCshqbGv81129jZoYPIQS+YGJsJQPxKCIqiiY7qEl2pCV/H7s4qwI5J
QpKBuGQOvqZnQb7BoA16woMI7mFtfT8Ol+lz59c44vkKs0fNo6VobwELfbxhCCTRDG0GnjunNjTZ
by62czoTJGeDVbrnQmyS5AdzHHQZAFq2KjPGPcFoJBR0NB5j0c6hlZNuE4cQAoDL36U/s8h1e369
4LrWxAm0guIsTXdpxfnQScb4bkbP5oHuaX0ZBlVCoLR098o+1iSCrcD4oLbreXnUKWq2QXzHWXQ3
/17jxXSZoceEw/R3OY/fi3XtERE79aL5bKFuUhC2e2SQXyigh99H7fGRzIytBxV9lH/AY4Oo/7Jz
vq724lZOP+sXsZ1bitU7GzMQ2fiWY8Q+sL7dSZyg6Rv367/KPGoETPtAu53cdjqXIkKej0u4h6/W
ZGEA4YRj2RLSF6NdtSRkPzBz5L3r+akjUQVMJ8bIecttIpuh8LrwpieRu6Dn5pd99N7L+v0Czx6b
tZAlRlfIWAUos0VLU2ZqC9YwTnN2SkMtP2LgpLBSmSxLWsPq3W/D97f2i+x8yJiaEDpqsg0sVK2k
okDtl8NEh1AfIaP8if/TXYn/GOd2QsrYzOgbIpd7tiYCD0fuwA6UfiiXaS5Sg1ukDzxmuKPZOtlG
w8u9UXsJ1Tvoa5EDF+TEg8Crezwe4kYuUox65A8lWPoqsDUMXi1Dr/O9NPgKHSpHGUpOJV4oqwJY
cChyRtAJoYkzPkAGU7grCF4HYWWpSa30sZL7rgTlc8uTBbyEN/eEZEaQHyts3OJ1mWbe8bTkA6dh
DmD0CoOq44NJM0rfIuESEbCq34CTZHXohWC80omdk6BrlyKWcPBwbZJr8CpH51k27yWU6r44jTkQ
8q1Q0JlnhR7+By+Y52DMSIiEzf8WxowKTbAONKTyuu7p6H6puHe6UGO+Ot/oFXD2HcVJUp3b306R
Eu0Jdf7Ka1/u5B4rTp/WkxM3nmM7HMpY/JEkk8bHGZhqNJGXK52UEUNQzru4jmoWGXOpGlGl9hX4
SlPWNrqTiotz+g/uj2ox/A/BhRNFzlL+zyUZrZiESEUqoslTgEAAqLVQx4YlJeD7cqg4n0j4raaF
T2GWFfJkRKVXm38Unkg1P7OqRiATsgTCmxXDb8GDIXI6sBukNmEPk6n8zGvbCYTocvjQg6C6dT1z
elKI1H2frKS6XlbzpMioxM66pf7A55liT42fe5JybI97owIkiG/79H7Tu2LqeWfUX2sIc+XxWuoO
AdfU09sW2dcG9Z1QL345YfOU03YEqilMpsDwadQ1Icqyq7EdPxTtgoD+3ecERXSC0qmP5yB4TdTl
IQgehd/k0/A/rLUmniSDpZm0x1s5OC99n1UAHEpOiNA8JQE+8DpKSJyUy3/s9t69jgJrSAb6wT9c
XaRENZZsqbKG0F5j4+N1jXyCey7r+wx4kohWyxKjqQnThKn8DOH+sXZbabR1aoxSRhcXNteuRXQd
/Elmbun9bbq7H+EFcVS7ruaaqRYqR9Ec5U9Jre4wLLQUgMY8gNlJ/xJc/aO6X1/q0a4Xm8qh29xU
BkRXROGvvmKQKzwjEIYiRSQGuBHJytDuFkIstvyTHQ2A6mz0eAyfK0PsTCCwJ8MOXXOzHR6VxGjl
iN4jc1H3onijQll/EVRD06cfvA+b6oRECIpQO5KIXPEpIAlS6imdGxyY6Z+FtVUVgtmLyhV1KmAZ
XguTvGkaMmIWnl5vTxD7JsElaXEBDZ0K/KPAXl8gwDEjeRFCfrbmOYzIMcVHjOfwRsm2z9cNfVi+
iYe1IcTn96tpJ77tk582nlqeK7SJ5X3704RD9fpFHUsJGE9rTGB4cfIeVrtkonTb5kthq1XJdcje
yW7A+kCEoUffTNkwthdzdwvnyk0BL+dsb9HrD1AvJG6VmM+xXt6rpZz8bnlvpe3tFRD9HXeiZipG
NPKHeUEHUB0ngIOoWZmR7jR0Mg/U9gCwf8KI1uds2HameWyuCmHPV512bhcBBfqi6uKmXtzDv+cz
+bYrikaaxjtIQOlL0hbfDKz52aAywT1Dx1g9EbkXAZd2mIHA63CHiRRAID1mQWsTunRwxT80Mgdy
vR3BOxkpxsgwFU3kGpZjZjDYJC22xEEkPFLvgqnl/LmJYpI+JmLMtXXe/6TzsVAh7PRMlkjBJiKA
q0bGeYPl5SdJTC0LX+wFqIOAXmeJcpyN5/AzgapnZ4cdfNW5WHvD17FXtPR8iUcC5kO88QXb2buN
w3+VwI+LSwwIx0JujKGqbL8iPrQyIoAJEACfedK2ajt9cqnrUI4MbUaqB1e9emRmYdpWQGctTJDb
OjJ8T5LTjbsglriFyR5uR1yHGhI4Gw6fyVRrSYMcEOkwxtcrsEPXPJCNNps5FndxZGda2puWscXC
0+2W2SyXROOH1nY3bdZYEHRmmhiEfgQLkofB2YuGnZf/og8ChSXbAtyzmEgZhRhMo538fjLIDkxQ
yCJ/tiqNtRfSTf3VTV9FYe0gSUB5MYVeCUIwpeayPn+4SY3/gFE3XG6bAwc0Mbr/jHeeuuKC0nhv
AAtQt5x5+6IrDCHohO5LjzUyeyAuLwYdKipxbzpmPiZjaCIAdvk17P76afM9y3qe+gHfPuhyTuMF
wZUCF5Ydxj05w/+b6BKa4DsZjWuQXyCULayhjdO/MXeRSamvjhkctDbfxgcUBnsBnaXciANw2ENa
KN0V+6/4dJ8v/MEP0WayecEA/m66QHv+WED9VxVgIEWyAgDvBsNEFTt/1a1AmdBpdzV7I1v4r3Rh
v38o45OofQ7yuZF0OUtI8hlkmSPH0Ur/cJZxBjKRrU551JJVctSr8xv01WFcKJmAvwwP9HtjUcE9
MfyohgIx2/Ttthozh/kamWro2QNbGYhmPZxOb3/4uCz9uEcoiO9uyD6mxPcPLCwMPo5TeySNqVZ2
tYqGgHiddDugfIQc4SEDW9B89x6bHTxaoV9W2mTaDMtVlVjE+NEzazOXbqEXatR/Fp5PTiPwkz4E
rVy/tkXXANgE1tchYtvzTLqwqhlt6w4wloCnoppis4wnRK6T4g/rqlgwO2KhU7UwHY7yQZpLWb4C
JOwJ45MHXKpXcBmPhAHXBza70tH8kZanGrxoYrPrJglGGncZl13nbtP96pJUBTwBU/VxHHS0D1Pp
DY3e4oRsNZ5MusQJflUqLtMHkiRpZxJOUDtVhfeFcoyh2rcBcwhsNpyPj9kFH8QQEg6Pr8qYaRR0
aw3YCPjz53kmfsHXXtxh0H+8PR0qfQIAjaHxxKvaBxRxL5QBCnBoUBuDy2EkLvmHgml8BMe6Arr0
NFUdrh1F7C2qiLulmdxsB5G+0fIvcFpnR4ckwRZMXLdLf7WpByqkRhYAQ79AeHgGxhcewusRriud
GJ2DxIxa6n80HL9zfYj8Tf0GN65arEr0DHe1cjkyUrRiWWw0wV+73BKWrOOiFzkZi/5ZSlIEuHkv
usR19hrXPPxF4c3Ple7p0a+3kWhruGl7NxN4+/1N/IG8gTiz0pKOICbBRaLg7e8GY6sjpwuG4r8b
W+ihpxNOoGGOB3ccAP3QbUshgZ62Rpa3vcK3iDiHSsWCRA9fHz61U+F7qRvNOIUogIta+Yz8lbU9
034y+Qv0h0KwRd+rpcOYypT+McKy8LOB47psXv2MsX2iVTJ43OBBXBcK6TWMnASQh/eY0cLgQ/V9
s2fo59VZ+chIGOaqqUp5vGn3sMoZp2UIfliF1oxnqUYnV76KcTVPg/VEOq0JIYFaP67op9KS+0i8
1BkvEZ/kqYYG9reoWNjHOEEljWtO2pxi/N/ENgMIksdkL4bF/wxo1LsT0C1S2OOfm0oi18mvTbsZ
WHzgsCm6dQDB6oMgqSDBiKrWcQCBQlrNHbGefvBvIht3XwpTwDsKX7rYGoVBdxKKw9gG4Z8SCUh7
nx+3701FPpctqD2woAJODHfVYeK4eIuln50xoI+8fdrOka54qoi3QMo7DDXbQZ7JyZIOGd/hDtEF
3FeK70qaT0hj7Md9RTwYC7+BvdZIuC1aPrp1ih5mJVKkpEMzodrg/1JvV5HsNHiZlk1b6MJ1QlVf
+5g0Ng/W7IvD7yMCZ36B3vq47VXtA2Ly6yEf/bNPk7/fI9+MbwTpXEr5CEI/3u+54yIj+mhuasHu
9i/Bq9hNRrvmVN2lmBPe5eCEQVhekyJqIgAORl/b8yfHdIUUCcOvEZtxPIhvOU7r2GeCucpnQumv
OWr4ic2sldbKku5gmnPL97QUPtTZV6ZA7nq7BiNGATd3d+MqJ82kZcIWZhYk+NMpRGGIUyxx2I5I
uwLQi1RtvO7uL0O5i9szrlRd0u2Wu4Sl1xELnKc4gkMoQvLxEnX0NmQZ/FgOhdL7kVhew+eJR/JL
lL+tPIpTT0+95RhNZ5fjH90d67qb5t08JD7kcfTBnhu8jgNe32ukdrhMbxyEESM88Wi3r3bfD3NW
tmHCuSd5D7B1CTX45aOxUz7WrgZxYepXidWivdu3zWzGBnbMSBziFLVB7isyAQEA21E/RG61bpl0
ft5kRLhy4UJDyjiQrmcly9N4b5Un8X7TVNw+BV3v6uxb5aPfC4yG5VZF1UZ0BnXfLWRQG/HEf4+Y
ak3As+4602F7u5zyuoWsVHXc6vlNqBlYu9A9JdgHUWUg9XkvEJGZvGI+X56/FJxVZNWszaHyfFfN
QDQQIEvs6V1DJSjezqlTYhpbP4vBdawmq3P0PKOt2czzaynUe8lR0FeunAJ+W1huLbxc3pGjoDF+
bGEhvuPXdq66vLyvqIHdych5o9QKtTkELeh2yAwLWgqdsePOoZXNu7jzfW5oiJcBCRFG8WWjLb3l
QSF5f5hqTepZOYP+dy9OwO0GJjiNk2D0+l4i6eny0sRag1LzI6ENsd0saMxdw49l+6md2MrQdpDI
6s0kpLJAEj23Uudd3avSYhdRBDR94sEl1U7RIAWtWIwCzbDSaFt1rPBxQEGZsP2lXQKV8q1qYLWJ
2Uvta+hYbLVAZGMvza7BhaG0IPoy8Yxtah5/zwk3JVHCvjRZwrnSs7qdPl7GqspeH0R4x0qfmEd/
ighpxmc2q5rdrTSQyuWWOSUlSGnAb4AXGH6sp2LC21IWLxUhEjJQd6y1RPOSkfQR0kJecBJF58z9
KBAQ8EXr2uSmRU9xxV+piobELjdIkxGWsAiZPjle8bbehTAigAPO0GRsFsSHSeG8mRK0ecciUW3e
qzFEiugNJ7MQwACdwpYGawUx/kThbzP/Idvs9Ceq+3GdA84mwWhRWhs7U6W8J+3rNfekQg720Kt7
Hr6x8VqqTtH5U2JwOpK7ISwt29jvikrNN+Tz9R2sRj4LjOXxr+MopNygfAICjr7JouuVuysi6GBm
MofXoGKn9J2/Lh4PgClUAugWnMWzROXh8INmnoyBZdVtkLGoz/fRdldT71+jufk3nEjMSBL5B4q9
/LrPmLxclxGhlEhgQQlzbJZE/mfUW+NXEv8FQoz2fuEmx9i9YlN6Yh0YeQipaNKNCGZi5tNPuPmc
LupS9QREAiJ/QOFKD8DAiRIubEBw5hmkNguYmaGjVqCLsyZiGsuMuddBeUeFgg5lYIVzDJsPztk/
nO9JxGvSml+RMktDhkgwL4kKmqkUyTemBXe1/NxhFULyvjB0k/1DTx5BD7tQObv/J69R+ck4v0iA
6RX0ZcKXWWuHItnamVmVMDrl1nqH8ShM3QhIVFGfpvF8mRGBpi6mJcHjUwkrqDvYi9IGiHFtw0Bu
QcR5hwOr24uweOwrh6XZw4I1tjmZGd9GQDlz3C/ISPG4+0x7YILdNaVwOAJMkrHe46b8l+Fvzghy
vIc4d8wWpQ/1qZ4OGZkB+l2liRobbXToqXm+kByOi1SbDce9MCzCW8cjoZ8UmDzZE63qMrceLWsI
tbP5MRAVMnSdH19ISeAalgUeTiWRCd8yXB/HuVKEUJbpiyMUJpHAMdYule2o2xzJnpobK2Vx57d5
GLrbW4OFqbXBbYzHlAkPA7BdtadcxevErwsmt2BCKuHqvOizc5IF2+PXhnUEBnANj2Yrzu+o/m+s
VYi4gER+NdtMYA2RNW7AwARI1/ukm4skhsv/Eu7EpF5FpiXYXvrmCjjcNcfCPAGksCzYu83oD4U+
dLAFqFJlcSpmCC68NF1eJGGQ2PzEO2gORIJBGnY5LlhffiLIa+6Kxn/pkD6VJ86Ti0COCfj8Zizn
kOludCTgBqw5NpdNeSwDCz/KyU80i4Fo7NTY+rm8DkXf6Je1olh81jymbdz7XOU1rCqGdjWI4IbL
aDGZrS+MMTL4g3BhpS6OtqPjC5NM2oIrIBSDbcg2XqZn0+rAqVHx6zDghXKLinE3wPrJ8tNHmwn6
R998QghYU3KmrvA2+glAFpalsYV/uARKCOt4RP2GZ+LLYWmCAkjNjwZDXuBy2w9txiRKP1e2El1m
x3PKPEomhd1j3/CptevL7HwQQTVUzRHPsAUVdDWOK+2U2nuArrDukpWtH49uFFyggn3r5W3B0LZc
M8Vn2lSIwxerjUX4z5zQC5q7WhVsv6FZULA0trPigCXIzrj8T3v8KBuHAXmM4kBjSW2n+bahDjPk
eT+EOcC7mM9GkAh7OpXxcMIlKbEOiFql4owy+M48PxY/EMw6/GrjhiIvpKOCp2NqB/YKkdu4ufKI
8KhcypYW4mcM0W/ZVoIG7Ut+ldd3fgcVvYt8VcIJnU6pcCCWCyg8EfJSK22zN4wXU7SKD3LQ+hSN
LGqpyZS5PGWKFDJpM3MKyWXCXb/P1wjwYPOZNWXJsdjBZv1HMI8oCAyg4Tqli75p8XdoRhhMltSk
vjK4i8Q+U1bsHztzg1AWubcU8pzYxIN5Vr+CHjjSlToZ4B4Wc0MavKaRgWuHpPx+zm3sFS/lDeT4
EMOr++i6IIY4q4xAN1fpL/BzmMhe3RWN0TbjPIRFdybxqPCcf9B51K9OopwKTf/TK9h70wZ/BOtw
/kzB43wdpSbYBypcpMi9bx3msNvz9ijfFklb89YmCfkiE21u2Ud2EkfCawflXAj/cL3PFxHyCpxh
jw2OzlCzut60ojEyuRfirukjTvuLvE+bSB9dRUGo8BFePwOoctk5nlp7afjuvridl5EOv+jHo9nG
spSomblNfVqnpO02v2ZXLRE9I8DVCmK9NB7xC23M0x43/JwHOl+mEwptio6Iz+TE1FzvB+L/Berr
Hke4H8UfHtM+F+F+QXdTFxeC0G7KMEYxbtkKXVxaaYexj4W5QWjU7slXvQ8+eejsLaqHwEtbK1D9
bqf6yZ/xrQJhFqbf2Vd5XuxNqUce9WspVsRqaXtm3zda72rPeh2yd/kDY3Rh0qJ0OGFekBnnxBgm
W2yvc3Awf9sIm/MyGBxf0KiDt5f/lAIxBBueLbRRnz+85fRGXTjtYLv/8oBCCZX2ZMmxz0n5PEwB
tz+1A4V4ZDFEfrFhph59wLPB2xiWGFcHX2hI6QVGnwXm16KDM22g+9GmA7Rpg2XybUBKTtSNPOnW
xdGVzAr9jP3Q+hjqHF+clcqIhr16UCxRJakbLUUuEEm9DOwX4L4OEa96V41kucbEIxEaxxlgKcZ4
vjpLwso0+yaoaOnUqMV5gkuAvWwKVqClPB+FU7bZ/rCrHkGE6asArAMOvAZUD2xYdhBkzR3KgvSw
3yRnLzbFjrTMhHnSTwtuMpWdlykU/RVHGYun2gUsBe4tlyIXRbVRmAUGgWlMl9+JUby6Wj5BMAGx
jjYK8bKd//wBMvS+r7+J3vkY/HcnYTJcKDjejnBkOduETxHTCqmBjOoyHCQC4Jb50ewWvkiEzBOM
pC+XChQfx0PlpIyuANWHc5Q44OjhiPC65JJzNWk7kaIDItSCm+BaxWX+/OjaacYHXDlcAord2bsI
c/MD7uNC9FawwN1NUa91HvG5TiapedDbhPdkjAI1EK9+/6c6hoUjDHXQChI4Pl3IGXOMVW7iy3/L
Xm3o1fV4cDCco/xLOWLlXGR9d24VY4dCfVIYxpR30emU8hO4MHEw5aPpodfHzUqitPzGiXCxDEim
NTEUQoDBcQUwvaQU4AfokMZSOPffcO8dL1vQ79op5qGjXpXJHYa3av1wMnpDt+yE+iMr+yHLCccP
mviFWH2WIQEouj7kR/A70iNlHoQwMGNA/j5C6OoDIDpw0JuGIMlVmR1f+fPmUeBD/gady2kdkHkA
WXQNd/OpV+E2bMT6VY+jvRdmA946rFMPo5q2BhGzEUbkcAzXvGQSo7tsnd9W/ALiPXilPvA+i3Fh
ntyGXHeIVtgb6vLORfhTk3OSargfzBtu+7VENWgMp7i/rMsXtNR0n1PUkg57HFLWJSasjsDzpOXb
AsTsCo60VfT2cLuo6oOV5Xg1hzk2/dt7RsZSqu/0sg2eJoiD0yCa6yiJeIqy6qBnQKdRKJKOrChx
J5uSuZSZljang7BF7wGUF+JswMGie0wIrEmThNrwDxBZ8XVp2fW+a5ky4/1bpLGBRmpdIXAcHT/2
sw7lxX0lvuamz1fHO/2WcIUkEv0V3LMQ911vKKKQB7DzMhzrz+/6eEZt7UzcFZty0JXqxth+Zbfj
K7BefDCFIImCHIRMwzNVRwaGvHU6M39AbGUQTxXoQtNFdaqjNngau9sVXHRfPN0u3FSOIAnYW4L4
6GsNqxI9X23Hzg0lGxjeLrRLt4zGyLsVILfFa8haCuHJVZM9r11XLD8JwLbc3g8zbRO8flDV9dev
+zupR0wGSlxHdwrdaaNpYcE6ePR75oEzXZeptZw+YUiuufQdfiTZBh5iBJbDpeJmfAZz/0sYINeF
QJlRBiPiu+q4cvZpb+qIR9P9m7T0ezCyzX0LmmVxT6fq7M8l+gwBBjQjlp/Enz80lq8sK12qb9ep
4CAJ+bZv4sm+Owq7mYIt6DyhpAQ9ifWvVwtKWMh2eC/9YwczrSDznO2TA50alxTHyOKqL+LdqJOw
ZGlvXmWdykmQ9/h+71rgd7Daj5GE/2rfx8RcYIQYyG6NHaCKqvl/3xyA5SreZD1Tt/9MzVWOUsoR
fo4sz6osZa5vbgBS+0vDovppjfo5nInT1IYVnhjghM7gDFdcOewD2NoKouMoXfF6po6PGx/Iy5mi
TgV6VIN4Br0e44M21G+xIM/GtYjXXMBjT74UdkkxaU9Wjwk16UcY6qZ8EtYFDhfMOWm2G3pYFriw
fJYM0Cxo5ZGJsB3+zr6Wirl5mk7krA5hNxgiZdCxNJRsE+QMHQ+Sae5v0sSA4w7Lumx+Bf31xxrL
84EJYDgCuB5Ry8DpqzptaZ8aiRjawUXohxZCHt0d62z/s9UJbH4TcVZsHNkIEEGBCly3NKsxxPt0
PlZzoWdAqFmrV3N2fr9YzHpuXyJOXlaeeBU+fwZrz6kwncEwWtqDHCSOr6z+oc5N9E671F/e2Gme
DR+cUuh9vfGrLKn6Dm9mbQVycmjyjDP21hJ2Z5ZoZIOW5TGPTSuSZQF56lwN59nW0Jc2XVLx1tmM
cHTHdwoSRWfkSBY8Ms99pY5hFI4BgbTrlAs4prMS1oa2hB2n4s8VABdlP4RAfjVB0Jvk05ais0hl
Gy8WNA4TK0uJq74S4kOzQFWWxoGZL8NTqb+dxBEwE8CXfhZkbsjTreeFJ/lP0k6gTPtdXccnqox6
O2au1D54OQkgb4pnpkucb4ZYBjsUXYoU8vRTEg6XUXTo2a7pOFnF+Nu9xsTIinBXvLD+fLlnhr3z
ghAayQl892bIcN9V5jmjJHLAiXOm4j1qCZFcWqcuaH+CDgr8Y5SCuraxrbAW7FfxYXUhI0E7J3hi
MhSb6sXfSdIKmSG4dHdDbvJgY0XwwqaZJtwtLn9bVSl6ZhhXryEsuPaXNYDSDWjMtAPP9C/ntIxR
kTYRD50chk01E5QCBULXK6/O4dS/ZrgI1Msltug7gyL3od1HA+mjbuDj9BvgFo41ck55aDuJOk0Y
exSDJRG8M+cWjGUTgeA6DfbmQDf98F2WjEm7aEK3PzojQ6qn3Ht2Y3gAPFSjzLOSUl8KhLB/31Tz
9A3eftOlqbclUcFKHPZjSHPgfESmI6PHmctknCVztZEPc45l+3SVFf8vRC0x1g9qAqsc6P7TKlFw
R9lhBMR0ULIaluyjVoGEII76Z9nIpZJLAybBgsqUWFijZc0a3gDhCluUrmF4bRX4bWFLVamxQMA1
HqPmc23WMPyLMlHkduogz8DaUBA6VPd9uKocpp/B4RrgJVt1usO5/rS9fVBVtu/YICdcptR3hzlJ
ucrqt/EJC9Mw4Xtn2NSzeylNdOY56YNRLDjo22JBbSKuXUiTyO1XzReEKF4LyL7P6eIrtW2bQlxo
CVwQqdox6n+2twqBamB2rlGQ6itO6NK9avKWLvpfI7yKGgXYQ6+4YsiDXV5bFMIb5XO+MoUWwFCj
PUBQwBnXR9oQ9hIaG4ULXAL+diMbrSkRL0fdDQYz0pzZANBAiwGFu1GsO79w6V97yHvYUUEJxs0g
DhETf/yioNx51FM9gucRpvYfiYC4kXQcm5iDkUqtYpuvNC/SEMmMbUChGvtCJhtGGFEhuvzaS9Nm
qRnm6g1tjzKMC9AUaokpuyiMFkcTB1ilnn1OwM6xpnzYk9CsH8ZTjDzqJqsN+UR2uhPEfVotHTAR
YPwjy1GUMSvjPmcJNniVKpRIq83isojejF2UrwvrAtB9NrSy4kOYW1YjirMIvEacFzA3y0QllXDb
L4Dll88gtkejg+UCK0o8dgb4ge4HVprf7lWvjqBQyYW86dYurPFZDdpVmrPvOIzMWiFhDSbw09ij
JvSLcIW16B4F2kGRFvD/8KnM2uMnuRk8tX9EFIY2nlWvbufg7Lj1S4qrTHFduFe8X79XCe7yMvo8
xUCt62t1v4vGBAj3cq7fdoyQoBhWjSjpSsc1cum5OX7mxh0WJbf3RoF4jmJikWGsCJt7jBz3aHgl
Lqb7NcWnRlX904cVJy4ELUKbm3yev6Qool55CmvHWHJhELvWI47DbklrmI4iAkBVaM4Kv4qO7ZvI
m5Diwji2w4Yur+eCP85n6+p9YjQ3ehVUKbLw9I4iA9NhwgkwrICDfgB24IiL8IpatneB1+QP8MTg
KyOX+i3ZYGpf+SoggG162JQLmn4p4nAYKil4XICXEkkLc9bgf8G/8p+1wLEgD5fb1KAZ2uGZGOIj
N5bBFjXViwX8SgpuX4f1Fb3FqrDqTW2He96kZ04ZQwU+zNyrhBK5Gph49rkXu+ZPa2vPMkALyiXf
o5YeAi8cKqzvigbnN6hqe+WKCpWnkPkCNVGY6KfDnfun2ldJ2DJGiYXIZUPXI+Tc5fQdouo7GjGR
Z9SPNVC3pglZPqhTBZUTzssrLqgUVPPn8ojA0eLjvejzTQ36zHc14dwXr8mlikbf3dlP6VqHYAX+
NrgfNzylslIfF6tlUTJDEBEcl91oWS5nDbeSYSFa+i2UeZKsDRY7VO1c1k/cD0WIj1fjUmCwfgS1
069pcBrZA3CHiDF5fsCJ+PANq3gtRio5+UVmGD4bRhQ2NZ6nMZ3dWce5BggJgwB2ErWVrclnfipv
nc3rfPTuD9QVYy4pOxffm0qTnWjte960FvfCXU61lSRyTccvw39dHJFgMicZ1/S7s0543vyYPJKC
bCFq4oDGCjonG0VrtcBZcBJ4JAP87OWU/uaEhUW4IPib/XaauNcrTVUq2Zhtnp5E4I2lXFTw/qv5
DyqwdXjMayESWxJ1MAAnWyQx3THQbdzsE4MEB2J6+jgAozcxvjOKjk9Koi9bKXTyisDkrFcvr19e
qgq1ggsj2/JT97AWc7DSZy/q0RVFITYdK4t6YqcI4A2BXsCXLtSUGGi8rMl1bEFzljI8oIisPV2k
aYxZF3mfsRoIq3Q0S2ahEuXl4fcW8dkkjK5lYYekN9QH960sNoIdMgiYEZOzsB1aA8DAYdfbHysF
OjWPwoaT6hbU44W1ddDkiM/g4u4vM+ZONGEbyPpfMXUdD6ReFzNG/X3MV2S/kAchYyw6ZdOhU1Vs
mPcRwoOTiko41H/frL7cmFLk69bUur6pFmUU8lQe/TbzKaf+NFXrB4JHYUn9wVV8P6MF943qOZxr
jjNcRjhnHHC+JNvsv7FICOXMVD8QJtqh5RO3g3nnagX4Cqy3XTRlbKGEOVwdxIaoBt+jTcr31vQ7
poPHADcpsn3NURJVOGDCvr7pmGICxvNf31DtSVwm0p1UsosDnwBB8p/Rk8riBNtlZt2gatmlhLg2
2ABQYhP9RUuZ8XUrd/BkuY6EDxjqne8fA56fsU80jzDjSLPSxnU8WjlNUtP99jhhYCIR1FBw4ydO
485cafOrS1c5py/GBEga9Zlg1vCLvaE0PTxDjj/xtJx/4kSowOTB5mej1+6wGdrn85OkBUC45oca
nS0a4bXqbm/Z5fisU8gAAsrkmG6YZnNSAkNrgGTmuBMPO19WMIek+Ff0GsjuWp6RO7PvQ8flc+RK
NzZ+mDrLM7xBsjh3P+aoXfSnXQer8ZcUqMZbxJKIQO89dWDGC5hOBlir45VaYPscCy8ccxnw98Xx
+vWngnvRFFcXZJ5tAUlEH538zb+QwWkV60mzpKWJ4HwfY0Sq9epmczhIy5bHAZknpj2uqGJTWMuT
7lDdu11TEFUpjlL29wg5FkXZAU2iygKC9SuFIdB88H315pVhY6qEMdEgN4E0B4mxv+fsl1y3Wd+2
VwhKjPbvxHJuus3v6SYfhWaQC9+FI+aQm8CX5G3WIlPC1V39ZLnZ8zcxxxPzKksXkZMy2zeSlTVE
WNXN7sMtW5P5JThnmNCjRcTYzEGNa0Ka44bqLNVzIVVIb8BKeB9SLrHob77pOGNdCaIBZDslqCQ8
F0LzJZNRlp2G57KkpuNunYnS3+Qz0y9WaiDpt3awb1wAACZwcaasujyfwOOsB8AlQDBEjaSsNpm+
i5HBFh2AMyEojWVZ+cvtfid+hZA8Y951Q++tfONR4xYrRgZWZa1qCAZaWjOMWAvLtjaaNhfeiBB9
aYqqasVPAnJ5EyVrrxF/DMjUJBgFsg3ye7uaXjhc4Ux8ETlMZe13ieUl98BWfKMkVKWeJdpzLrBC
IlzCzz2mPNroEtYXvub4h/hFZcHcMdptjVMOTRekylJ+EG5R66TDRCdaxCpIXg2mfAureelV8dcE
ba9B8vfpPac19hTTVE4RSOj4Nvuvd+jv2kBsQyzxce/ukmYd2aCqKMXqaE8A6M7sgOnUTUwW8N52
X8Ld7UyXMdwWBsNa+kbhX508eYE+3KCK8nFGEYP5b4T6emR0yxBkGAjN2mmCMhyYR6LHFUnhpUO3
o689nnXjnzppkQyR6pUZi+M1Lz6yIdxEe0cVCIMcXd8u16p0TQcCgquwPQ3p1rHmIXWP24fHzP6f
CncTGVQ3AqznUIi4NM5IfjIBIbzVwDyf3RTjkqJfKEW3LTVOj+mCZjjVx9uO5lg8mztHvtywisgi
E/9VUjLHSJgXTzFiIYNwnEAEMYrx9uauJKozd71NbbFG4EXUhJsFclVWssnaWWzguAm2c+DVEsxX
jlvcdpwQYUkzpB5L+cLa/XZ+31kHoo/jTb/sT2IOyVb3PN6V60sJ98XTs9PYVJxhJOCSiATm1uIX
QzJhe96Hl8DM9YGsKbGCeGWFs0U/UIbY2YN9rawtkFTzsVhpl3OOK2qtmTnssnx0cTNzSNm6Fxof
4aa4+4Gs7N1mTtxfyzpg0bO1kQyOYlv0NXsfRLzE7jgTDbwj/H5xvDw5QKWY6Up1PdZUSquYuqow
w2lbXM4Q4u1YcPQohoVzDUzAhihqWc+poiwLaIw6zfAilB1Fh80dcppMwmVg7FK8tQofNbu9kpYR
+QftrjCvzNar4zOnKkYi4YA31VeT6zIemKJ9quceHlnvdtSO5SCQHp0t2WbimQ8mImeRdh2rvdju
8w+eyvq+AqJ3E0/4jsAbpofdVmvMgYpJvLY9je2wiAi3KkBqrSXfQF3d8Z/fJ0QedEEdyjvXJLoo
P4w4DXEOi+h37XSolNRz1PXurPuiKDBTLNgHtXoVJzPN+8Hdf54S619ed+YgbIqf0EQOq0KFddWm
zVGmTN2BxlDVwJAh4Qb7sKC9Gp3yV3r6dzbcqs9JQONL6PPndbMDWMtUe1GDFastpQxloepbCPDl
VVfrkCY0V+AjC1gRA6XYZrnpBiIswnVcM6TwyJGd0kVVEzrRpzGgJMUWPu7CsKUa+H897BwySUUK
dvh4jHmu94ccJ7b4IR9bT+SBQBU28Pree0C3ltilPcgb3TqwnY5S8wVNroSUbcfQV7zgMnfTiPvk
h7Q9Ii94ddsnRhQY177To3o7BFWEXE9v7IsB5uryMDd3vjxsSrilPqIiKghaPdrbfPqjUglZM45Q
EdJbgozOZff3SoebYzRPXtOxhS5/r4F3Yn1LQmJlolGynSC3zmO0G2sUDQyR0Tx9qL03wd7e9xDT
S1SpxrFq1dhwJ70JgOA8Sr9r/lD9CJ1WyTcfQdTnEQbNy86ONgYwDfO2G+MdOBQeT6zPdaLo3Oii
GP8NyJBj8tPsqolCEE27p6LiBtRBx3omviRf7tnFgJBsHmbRbtW56MnG5/FfGeaCLIcUsO1OHllH
dFn1CGbh07GUWV5ZBOm7gxFDIi+PDws2SOE10JSNMKXoPicMu890QRRR/Ad7PW3h8TTWvicM0QH4
X4m4LbRhWgqDZTAWSmi50nebBRNFQFk+I4GEjBLDv31oYIwlyYbh+9n+luVeZqBZQsNN2VPzZ6wv
u2UNnJ/2xvBbTFfBW6wnjqD5blBGJG/6JQL6ZaAYPL/VYKMd2/aih84oXBpZnjcyEA1W4fbimpfQ
e/DOHWs+ugX51fkUWO/U5iiKb4iHvbvQtW2eCz2hNYhqGuAdMgwvXayooSo/Xqm2ijiYPsLezTpj
0Qg2rchZ4W3etVZxLsHlfaJmYJHnle4B2hX/xeC/7SdOK16FoPPdGR9/8w0DhNz521qipRglbkUl
SZhSpKEK1CHVyBjw+d5kYzr81CkifyC3QhSWdN0k5qAL+i24psUghNGg6cNoFkPIhOoB0rL/5KUK
q/4H82cCctl5PTX0p3fUf6d/g+5Uy0lPcTQMFG46axyFUI0PWuECPr/qk8iYGkO44uvFrosSgj7s
2Peq59X2bUbXruak5W7W1A4B6eygYDxnKbtGKv9LYRk4K0OMC3GYUjRDYKHxWJr62KbN4B8jtdMh
3N1129Y/cd802OIbjl7w6nEUtHOjKtaOI6ioyJmJ7tSsq3dvQciD+jzzWqat29077B49LZymRspd
lCsaEiz90P5Kah0uOUtmjH1mRM0beltwPYsY1Ha3M17xLRLGPR3wnvKdgxtJwiN5Oci6wZ6NBqPi
xDVBy/dOv7d0vi10zmzjalkUJGh6FFc2Y+L7nF2lmvLb23Ik2rwvWwN+iUX5CmJnySpf2xfa2MLb
2+5GC6ebXi4pes7gq0tKn02uyGzSC/1hRuhncX700cIEq6Hi+OB7zrbAG4mnUgigLRAQ9NrB0r8v
I2BLXyRB3BmwVSk+Cdew0CgNhsz7i0yi2VC8gwEpgcYyk5THVwmPqXr5wmKdwSoO2YbKBeywXx31
9re2vmeO+fR74BYbKT0yPI7dP15aLHfdRbDVEVDsLjmmRkU4E/MI+mQgHvjKt8+R79diGqgj9tbQ
1pxpVHQZU1YmBXwa1W/kQcxRLijXufImgfPtfCG8jrp7SroPf2XAFCdyfTIz0NgHJfj8vBB5KDYy
7wDoHUOmOqBs2PpEW3DvUdo4zQFcSm2PXZ+Tjw6O5ilveEJKAzVgNZkqmQVkOG0/KUX90Rf4GmGA
Qt7R232+klYiIEJuQI3qMgtlNUh/vDZl0fKaQtoBM9HkwE7MVlKIU4uu1de3VaI3YzZKZlxB3Zkw
KvM+wSapXHRaa+J0IFFPQuNoWMWdF+Mau46Lh5aBZ5y7JoVD8f/M3fx3B1zme/jkOr3sahcQ4h8R
a7kQaWMf9ow1LM0Bi6HgLPx1OPixzzDPyWQipPBXqbCqo0kschYHZT8HWzHYHr91ZeTf8Ra1K7tl
nxgGBTUIIXSdn8+3Q90Rah9HTA0t629ybjF91w15Drj4DwSoaHUtqOJswrQzVJwXl29xBZuPTGsh
t4If2p5PC5eGOPsKGt6DA9mLyW5PX0LCik9qDsdr6X9VJYdyAefIL3F837ZsS0x74chviYkCnV2D
XSAw+QgMfSIr9mFAvjSDA1lfpjnogHlYoIfM0DYdfbFNdyJV2IO/QIQxUDxy737W2+7RABotRFjn
CnA52qaCQ5FCLKUKI2B0wvlHyv78ebjEaRDRAXCXdhS9qRE3s3jYke3YMt/6zl/7OdXn+XlyXhQY
A3yWqXh/MLzMigp6sU85geUIDSD4uYu8k+rTDUSGyzuNZzGQBLWLRduEGIM4f9IEemp3LsRRx1Aa
QQwN+Jp907dwRFC0no9DXh8MLrsRdoo3T7hd0pT9UOnHTLiYeBanWd5UQrJ6y2lXzA8aACkb8YcF
NMRYvdKb+MVoUvzG2EZuS+g3CATEECEdYe+qcPPq+i9HU7ncQY+h+TJXW0YpXNOscYnXJs8tvchN
1uKqVWehQoIg0f0eZh3RY3vTPojij+YhTDZfk+Ji+lnuQDTC63CCX1p2EzikPFqgV4tuTebYx1/a
AiJTxLk11KYvkT4qDwesWf7peNHGA1ExBi7o8b/jfgT8S5PJOLGGcsXw6jc6mNoLxdG04VxKyjcy
naa+byA4fNygjgYsxpXbpss8JfNoO6WiH9b2MDjLRSs3p+EsRU+dxykFO1ndtz5vo790zfYl5H+C
Mqy8PQnuaPJ8UJ2z60n4SjzW1etVelGlE8MxSl2LnQAMofyg8J/afUhmmAp6OSeGaK2JG34262EF
NaY00QCj3frzrmHtou4VpYARRhPK8tMxHQjzFKIf22i14CTjWwMS57evGwgnD3sL/z5ijFMNbK6C
MsBQkqCRdBU5vO3uO6STwJ8lLVBG7voZjJqleEQ7psbCAuOfAGlYFPWn/9soQOU6V5h3HfY6eJXx
CfV9yGqAE9rV2HTU8HD7hsH2IgzTY2sgHgQsZFzz744Ec6gW8i7c+tp6Nm/W6TE9B9L6nbabbJIe
REu90eogDIN2N6dlzBJcdmw4esz5RHLU/wuXAjKlv8210LV1m/l1tdDL56gNiJcwuVogSTT2wh96
4mVDDbC2yDHWlm9n7d4cfUHVy/Oz5CJHQPD6oPtYng+of+Q9kRAPamRyA6S0UpHD8M8c7u7f7QIW
a4aOC17APnwzgG9HzGJeXUgUaMy7t1nWXD5CGPlfGNh34c92LpIByAJMNsE4DbS/6qa4tVIPOeYO
KoL7wW8HLjr6D0+EARAY4wFmdulHyDP45JNbz2QeHElbUCiRtb6MKN3DeJtZIVC7s0sIyKFZ9INH
dnUCVWFBmtNSl+QdHRYb50o2PvWg+C9orSOdKaXsk0/qI+2oMDU/qySkdWrnb6uev0pTC59c8dMT
KeOlycuwhnUbvnM6EcinZMfgP2kHAZA2o4l5SvYwYXKeXjdB0fEylBDKD5K9azYv+IwNNwj03KM7
xtf2vfi5hbWT9O66MTBTuAb3mN5rgKEew01NhnjR4a1rvyi9NyBxcBKF7Tifq/p+kdvFIegoOBBT
rhR2sNgu34J1YcqW81JDMbgtpt61MJWQEW/HOdRvk/7hsuTJKac+gxTyoob7eFUVU0mGAiCNoCuc
ABF6DgZI2wmynmv3XjyTXukhyqfNo+xrS+0X4nxflrnY0Duw0B5rXLGVmm9oUMiZUi1cwYPOTEPt
MsIbtNLB4kCSApTO3HZ66we4dq316k6m/yL7JulPovk4BjVFoekpJCl/Z7Vx+C1tO2t/7F5ZiCMK
qThIrqEy/UyzUp1rOyq7D80qJqiD6+YWUQcKRPx90m9GPVH1u/toK3E8flSIEGY6OFrd2wJX6OPh
q0ryKsWIhoyU2muV8/S9r5p6feJFdu7iXH5J6RcaRd6L1w/pD7rBXnzeXocbh73T7LFQapcfZzzQ
glFE+793zoPw5jjP6DlwQm5XpLzeahVMV1E7o9LEmn0nrM26vA1CpI/7KWDz1SPgC4nSlBWZcTLK
36xOugju7c15Wcb2oAbt8kIhiX3GvuYa71+nUFE6pnB2nVmXy+IpBn/X7EJeS5BM9ZewCRRBipOK
U863tvcKMPlh/ylVF3bGwEifJ4KZz8W781vW6YS9/uhJpboYx+es68dHDUbHEK/OvaM+2ksTy3XH
FVBH4UCkHNX17jLVlJO54L1BI6/Woqu//seqHTKmsZ1MyqQw4Nc1O7vDEPADXM+SJFdVxbicJ9eU
02gAnhCUr3enIVOU3YTzLGFhmWXvlZj5/7/+45kBH/4Asw85IodV/wE/Q9U7B+18q9LY7m/uGXJk
SgeC36mUxiguanVG4vUIepThZ8M1hco1fgRgtmetchI7BXfmhMt+TUFhqJHzKK9GZVTNicQo6nR9
1YpG4xu2KzcT6ZrMsPqf2XjUzjExo0vlUIVqrIgVFBaPhHhj7eWNnloH4Kt+IkCGmYAxK+UAbBxV
O2Z1ihw4XpRDZX9x7w2XqAtmcWb7O6z2Y2dur7z62pOt9vz8B6c7fVyWowlEXsRwcKC7Za6Wecj9
Qo7pdt2jtL4THqVbrgKignxdyIej8Uw3fAwfP8aysrJaPDLiZjqrJcIsp0sLZSGkkqTcD1pTCV0G
Tiwk/Lgvzqsm2WNbV8ZJApeq4MQ8qTkSs5yGqN225T6pesL6w2VmANKSR3mH1+zLhLrH2oXis7ds
/f7tCLovJF9aqI5BFYq8zIzEhr6pITkSh3asK/3PbsZHyJC1oO0Y/ob9eT2j7tnnFLc3UURHgaHy
Q9bExFfO6Ilay6v0cdmfotaIu+X+zKv+Dx5zDrjU9n3KdacZaGSf38lUKRwm0hOsRVIjCViRtOLi
yA5xFmiUN+EmFhLdDFsvxRIlEIaiEe/4IIaoacT4vSr+Ldz/IueNv0/qHE7c8yhGZJF5hc/6N0JW
jD1PwVHT/TGGFSxANhKzsICZOC67VIlIaBLA1WsJZQ+HzZNw04p1lA41d6m5EnL8B9o8Z3uhp3ez
EwSuF7K8WSuFKzyl0pSQxoaeccRlmA8/pBLXU8UuGTbdjMPU8/AYUdetRvMbt4MeRhNlrkd2+m61
vDT9TO2LjY5RvLpwQe+5u655u8Nzs9u2Mzv1mHQRPpQB4cmn6VHy5X0/+dEStoZ5HFnGmZ2IdEBB
zmh6hm9LNw+wtd09mWM00dIJnVQLZ3XQkGbPe3V2Xnln+Q4vkVujP5JvAs/VPi9Fkrb2k/KiAko8
fzldCpqjpxKgW6EE/eiqSsQSMxJehIO7tu6Jy+e6g0vOleYR4YWmJiwJ0cKnB3yvZsUk4fAa+VoW
BnFBmAN/3/9OI+UHQmVp0SHDIzT27imejEONlB+GQOqlZrJm4+5rwOar6Peyh43cXtFA6MXBiwqM
2kw7WT/wk4ELnvph4hq8X6mHAHm0j/+XHwK9NLPYIrk/YF/F//QLIruv69jjCUAdaGIJhjhrIDtz
EqSpXFB0ausGC621425o10YLdG1cHbgbuRTJ7j8iBl3/+AlJZzPhtYFrS74cO+c9fWkhbCd3yayp
/+NLJiLGuwsCo/oFLFO6rLVWcGSUzQUOwbVoQU3SF6RCx2yt6zfhOk9zyfX0rx1NBrMpySJZ2vIc
0ApLPu+iRJxDbdabnOODwT2m+LO3K5tHPVrYAZCbbYCtRflsZiFMRBzVm9obaq8oDEbfDO7y39fQ
iQ16CBviw/mtLkDK3sSjgGCIhjDUVAcDRK7kymSQgXbDDhfZ+nRetzEAxL+03IdS9yYcEqA3WObV
OTo8YD6nVw6/0VCWKPYZuLpPItGTRveYSzteFNPRHn8ot+/9gtgKEL2mL9ncAAqZLHE0s5daVe7T
nAg6GzGcmtT34BKuAtLFL5GRYP4aa43/CaAwtr2SVR6QJQLYy88NVm2pnDX2+cgwPExSIK6YRGrd
aMuhIgUX/Gwm2zrLRfuhCEdNY3IUuWTCYsWwT187r/uCclVwto1WGSzQTO1DQ93ET3Lrp4Bqptzv
ZoHyq2Z8XEogovF8UqhvNYWOGHUvCgT16xku4Ut/xSLwpmEUWkuHmJydMi1JqFVF65OXx1eHMrCG
9G8jp/1FDo0QaR4cUUdX+yGQbSWQXfjWJyG7zn4/4epxAYA4hHbrvbihRu3IC1eQVnfhYbPSU4fT
BQ5BsfXBw36fwByQR5XXIQP+OU0FCJl5MaV/AfQl8E+RZLeBt16JQ9mNTdii3ZPcNbWbSYWlMwb6
HhRO8XQoLtQxURSmdFE07T2ngBHCfOYPq9lNMesdPhqa4oGcq3rvcCMdIICHgEkQMCiACtdlBvQw
b206C40uf6bZTvFGHHg4VOGdycHTYBA3RJPtFo48zyIz8Bys98pg2xYmfJvmpO+aRW75c8bhyYXH
qlGNMGknkUQOzmH+NMQfPrbwAk19aM2swPM7HJFbHsERMX4Qf8lBv41rjXFh4Hl6iQx22Y7umzZ6
spJILsax/5z/VIWlaRU/wepQXgW6UzctT+19XQBlz14/1BDJZR/TGK95GI7gTv6Jf9YUKdnM03YX
IRuHxMQiwBWY9ZbQUAnmB0Lt2wF2rqUR5pgFIScRlhe6rLnllTfpqnSR4GZZesBFCOCwVnY+r+6s
yz3hPP+JMRmvwXiq2hjtncq8uyWNKhR20yS+Uvn5g/qBpW45FiqQC121fD9KZ3rd8kLk5Grcfpib
BWQioDWq0bCp7/LwYr9a9QkPOWrnK/iTgQJCOL6UF2BahyHdq8WbasGOJHrVnaBf7uUz+MasjFA1
oj0+BtesApFuesZ/tVXuCK3CvDOYpuYCp0Y/Af+QCqeIA6aRRg+qxAEnmgfwtkmYIaJg3AAfnxRi
tQQk8gU5brNkjokrVD+63+oG/9pjCZm+HMyEic1WkHtPr4/bydt772HImTraagL6o2oBOi2PF75V
PMRjKSZMchKmjio4nIwO25shWQSet/CulydOylL+kKLyDqhgINuVxUrC6wpyLptcQxIABKSIizAo
PrsJbGG4MAWvj8C6eUK0s7JnwiDyswotdm9jyzrySIMDmISmancHtGn46JPp4vpMfnKqVqvtqSrc
3TQn56gXvCtrbQW734WdQFZWgi16B/1lMBWzqeMG2a7NNjChaq3GZxm1FptUb49qW0j766j4+vrO
/X+6j6jnIqSIKQcij4hN8ptgUjlPnCVjBedkLdOFSfMaGYSPSwCMw9QILPPWgbBwgB6LKSm042/Y
YV9f7E+elPiEtb4QFtMZ2U0/i68UWELgbWM5F7JIX7fjEEgyFOzh9K3DFEQ1+/MrjkeIr0pqexHy
U1x3GzaULs9fogpK25yzM3Tjcj5Egi4htZ5pfOVNjlS3AHCb/wpoeHmRTqycVpwgd/XEz4ESQ763
jRdfNlR3omVGpCb1GYMDCDAJdSIWQYIFiY+krssFTCAHEf9GtfT1gGtm8+ciKXIht8UT+vOdR3+o
E8Oy7RO7NrVE78d2hdfaVIdClOU7P1221Ent+IneEbnBmLg4KX3sVGhvXvefxN4ftJMtNVju2+Rd
VNS9TC1fdku2vfMmmvB3TOBQ8AG15f9WZiL77oLtGA2A0hH+tU975KpEIhHlQnSGzEsN3jaPTcw4
BFuijKbWKqmvLltnZTZN3PRylet2XuUqvVklNyI31WC+E6Q8q+OoVbekDnr9qwf5+USf/oABlINP
dRlxq0KmwTa8xWHU5XI+v6CuqE/rtDzSKXueCZvlXRGcLc8CIKecR/s8R5n4fP7oaM9WRticwinE
2OV6Y+wTi08IArJz95ffr2jUEbRi+HLsq86sV80e68i7K3+FZ38vh/+7uLQyToX5/I+s+CPQBgqY
HNDCn8yjgb2kEDaEeFxA6ON8aIalN1gKP50iTHEMVAwbsZFJoYKbR1fE28o6gK0WYF6fGQ0jU1CE
vUtR53Jm7gwt9pJNHmT4s4muSMkBQLnLgpSv9ZEv+WfQAvxWRDGFBK0dAXSIKspg3IumHX77tXGf
mp6+4HorFnNbvfolthS2uoTKrCN71H/M0RkXTX6sKGfYfZeSAhSI0lm15WDCnrHOBio1ktrxhUjV
Hqn467Cwk8aqlAcq8iDdMhOTLw8O2qVBvKNtiqNpCvqmblvT6k0lZYbYwtF0XFDInkFHpB57ieFh
qawCP7sW0cVoBrkxUbDWM2FtLmHz5OHRovhnpO65cw7eejiYB0xfAHmb77aYPSrmpSkY3QluktS6
oLTS9N3Pdy+Bw3GXzLfwqTjd5W78TwvtJ1farbkw1Kfvh75/hx1gTAmGKKSi1zcBfoOJSSsnLVMT
bHHiikeKzy4GlzGxUUFto1nrqdlw6bSIPGsG4k+TYMZVNZGFb+vcZatoMtnIJmd+fkezu9lb+k81
HFVALpZpbqoyKOEqeUbxMkuVIwqduhM0yRnqgrGeqHHW9x/lo11tnckDxAX7SfqLUbyNXgojFDNo
zKHxSMB8UY92Vu7wljT1qvmXqjAKb01+xGl+/yzPfQPYl200RfRD19sgApOKzmTnao3Rxp1pIMOi
eQ5osDoSOjRZBGHbA0PNwF46ESHj9mhDW54Qy8VYG+ZLC5WgySATXn9kx6+6yCjky+7z3ICHKg39
xoMvpoyNccNjX3SAKwhPS3tMgQscfMhYVzq4nyj+Y3hQq3L7AV+Hag/SZ36oQtu2EAgO7J0BmVhy
7hFJPN4cueAojyC258iV2Rg5OHq15p50NRecH9gRZWaz+U4+X8Z1/MuGTYWhvyPOMHJQzVURnfIc
VLu/l0ajYAy85+9u+uwG8U8cFqG4b9gV1I74t3Emf0yUYnGaKEFJE9DVkrs3kmLwSG4Vt+rED7xq
7woYwIQMXMCrV1bBeLvUaD9wAGoZI9dbT3BRBGgJVfl7vKL/Ck4NEJw0vw+hpBFgd+wAKQ2xalI1
qBuqzC3MLAqC/EgI46GXQVGTMbhKRcH1AvsVZEWTlRKMr7u6E919ebIwNwWWJjb3Yf/lyNYmymee
j8rw4RrLpwLUteQxOKDPHlFVvWKZD+9R7yOVldr0a80St6nDTX7HT166sSKC8r1sEq8KeptgTjHq
OauL7LZMCEvQiYGM825jdgihgt4Jy58KQ9/eS4xTT6QdkojJUDO0xY3TmSU6zhibr4pLxVaYtnQP
j2Fa10bzgA7NFjTAFzwi1qIpUyKY59po6hM+VGYpvlzoPG90UDLgvZ2Pf66P4s9U1aG+sB/9YzOs
Jqn9h19O/AJN8DWGjv4vnVXsuf9l8rO0YtZD+tDEU+YS7yyFp215uYmDIj8rBVYDBkY8VaoLV5H5
y9wBrnMNtV3pzwATudYGRJPODpLMsij5m7WrB6ru9IK0R5trObcu3Qu3WSfldUGL1J5irvi6uqGG
iNkyJgzs6tB8OxpjfBuQhYBhCUZLKG1O+mf8VwklB3cyRj8Ww/5k0yINpwXGnb3KLY4eglbN0D7p
t/IPzTmJ5Y0mLulo2thjEXlFAMw+Au5qh3PN5vI0IlwNut0JGruCARBk3w0zq/voteYxwEakbTPE
1dTwv819t3qtoiXWYdfrP8xbnfeO3TGW9UOtO5q9nhklZhzKihcln/oMlUzJNBZTl3x4eJXPaMpM
869mLynll4oEEd9jXNGpzfXzjckCEBMn7+QZkqhdGDVDVu1OMRYMrA7J2hGvTtvawq5IC/8FY4bh
Q/h9zSVsrXXMEEZnifRxwbGYi1mWOv4dExhV0i3aWAMOzpXIm2GWpBkj8znFcubkWOrF3lUl3bjT
VOr2NYQk5kejjatrC4KITVfll+wXWqSlRvawZ5jViPJjNA3PtddO6wuG+JORN2CxsNJ5Prifiqni
Y13qXe0h3FN+PrTSX/uyf/lXVQlv80P05uj8zbscbyFcyCFsc2hWXyn4ToOxzrdW3UOoIGUcSTfe
SiNE7lvaUHYzfAMQAB5r+WSn6S4BkSYh/YfgQvXMhVfHSKNHE17WXgupuNCNTZt1sswj5/Wv7MHs
K6lZW63iPYJznQd3bneSeMFgws9hU9eTeAtTdklj0kIwv2QeDpEm35vvU2r6O/yccSm46JcCIZ8s
SG9PEsLUmr2TYm1rZn9+MFnR9rY34D7ThV7YRqgYGlaXZQh9VtWkQCPiaS/3rRUR2dVBNJ+XVlh0
XCZEI5rD/C84f7NEP5jE+9axWOFe4W6j8zu+2xonDPr/ePlVBRLy2kg7Ep8/TnOMxIOTC6cAjD3d
kfF0Hd9izTrhedKAnvR07tbxXxUjYhh4vOhn3ZyOE0mssr9godjlzsbfDut/TnjHppyHrt/iyFGG
ygNOySPCQpDseYTA+6AtFqzu9uO+eX/bZLdOndkW4ObDEr7qUcCv+f/Ly4uZIzKNfLu3ChOX/lfN
0iMXbY1jX9//A+HISMxl1wFDpfVeOFcQCbqjCtdod2BbbZD+pIE7BtXW+lGdaIPpxF5UA17GA48O
sgLDObiLtCj3EUqdFDqGrNUkspVp+pmrZXV/SqaeMz8A/QL16j3uVdIIN4oLZE9gL+CRp+20gs7y
PgT/ZpCTdz93nbgD3SZ0jc2qPjSRym7F4wYaIAHGa66uHem4PNVRsRe3pac+afdXJa9sTUEkqEfx
sJbRZ0SsLVyB3G5P2WDaxLcOfHarH3xjZpq2sHnMFSCKxLpvdlxKYYOqV32PShafq7b6vVXNJPs0
yDrHzZjO7Hh4YQAZ48E4KI92w/Hmtp8bAAKsjy15ier2424zOIwpmWkzyMSeP9kQku+ILnETqzJZ
+hzf1a7LnwnBZG0o2Fqsay9CiCTFt/VBS1DgNZnl0J7aQUTObLJzCT3SrPbNTjviWkKyIgYVA8ZA
G16TveFEICF1puPNBR86vS6CUwUOdC+UDwyfkSdzcU1oxuDx6NKJ7JlJBszGcv+xb13J2l9i/cDd
ZPoxMhnXl7gIR24gnXeIvwbN1DKlT10/f8zKhCV5QznzsNY7Bm4HLFV3PK3S4pneMRZGPYSeg/u3
xGm7vyPr+uMka9JQ357lxgu9sfkgIIP2wXPF7DzwwqwTUGn3A+kSALF3vUd/GFWm7WkWL3RZ9Fgb
KcIB05aAW3BNCkuSmO62xVv2q9NDzYKzxYY25yIVgVz0ZlUPFOJMCLDp3NlInRpynjKfHuNtZcGX
3WNVGJLQop3C6K6ipsAdo0NCoQeEl5UncTPnQIzpkDSe1TiqwlrJuM9lpEs1u1+ruM5eCF672Ukq
f+k1QsNKRAe2TvXjXuYtSys7SUjuab7HplQuhdn+WRtlWp8dCVAaeaIvjnFcwn0n8q41qhCML0XH
/VuSbYy+XQo5Kr84fYjP/g0cIJfC3MYn6RuoVbI63D2fzp1ye03dsla0+AUYQwfI0/BVCGQ6u335
i4Af+GT5IerYmL26UBRXPYscq48npY4XsoxnukiTOo4fPmsmwulqVghtRA+3UhYXzaFW94KhQyjO
7aikPR1bvpy26FXUbNaenW7SMf8GmsJJCXQ2MTiStSAJe1ZhhddpqhlheYW8JRYbpoqclEqkKsnU
TufYsZDcgiuOozibzUsoNlVDqcKcomhLz09E+h11kzjZO+TMroyBWdJlftm+fh48HdDA1d/99LTL
rVBV1nrslqyy9pTTgB6H4sp+IIgWSl1E3wepxEbrQp1veIqO5+WX2LO8QBXMaWWNwYiusI34PoWQ
8bGxKErUJYgRLCJ3GD9tRRFs7aJTod0bRYC7GTZ5XMoMwuCnjRBpYBE6aJDUWRguFnT4THQ4fb5F
gk4Ufpf3TE7gW/+rYr3BC6M364X8HWpkU4iZWbNOVUfx8QcZt4qc8l54tc0l4lDNM3RJqNUwbQXe
Ob4f9YJBSnb3960R50Pzj2ket1bHnM0YlHmMbObbxmts/YeSXlCiYW4daBmo2qSzxq/fqLBXnUgm
G8jx4Q1XIB5flfG/f0B8ZXabYK5z6c19Z/fYkh25zPK6ojVnPjk7tQhcvl0jRu5E08fSO+32cNqF
KIntH8ne5pcGmRXfjnyPN2F+P3iKfTLpkKiPi3jM5MKWuxkvk+ZRSwZGR7dmBTXpdXePwDBNC3xa
DSaqkjOnpCoYys61LyDOS4Y6gMQj2Qr4sIF7qh9rSizWM1heoXDO1CZIEy74stuDFGzr9/m+IOiD
ODG5Isfegpix250DAjRbvIiU+TKdXcHJMtFdNu7V7VVJhKQOHY3KVt9mQyKkwdHAUi2zc0R9GMs3
s7lNnfNPgt6GFzN0pndx3vdSmR235d3QyleCUzHAqnGb85Adm1Dxrxs03WHsKZdeGdcCpBhnDMwR
+uZbvgBckUu8JlKrvF2m+mpKIBn68t3NCYUALxKIuJDJUZbHtf69B/Mogdx6bRRkPOmvoE811f/X
YXxposu0mNmww+KNwbe70ytYVHeRpuYvYBOnlPlmBXTQAR1HGcHWBDJ7z3Dy4BoK2UwxejKSGbVI
ivpMFUqsPDFyD6h0bOWwgwvkwrEVxZIvDBQbqeEUGBEQOligfiYz/rzhIQyX8wK4Vrv0OROnpZEK
XEJJD/NNFkdfbiQiuMpni6Dj8Cuqcb3y/5sQuAn6Q0r49rf8pIx9pIYs/qMNjO6pX4uBju4FnUWk
8jCagaUWU+gYwBlMeV4hxDVfwheKU//Txx+trr2qf0QjSZdExf57cyDSV2mo8Wk8O7kTcu1rY2n4
RB8MbexGOOcneFZlCbMH8gSeR+4iPIx0+DchYxpNrWwzX15nx2wwfeW3pdgDghnMZ+vDZEvadm8I
zimK5JIza3qOZSvPFcsYjJI1pQKqKFNF7DmeE8aFKus9XIkzvoQqXfR6i08D16SDbTfq1vMu6ptw
SaSGAJ8JQubUCD8l538OHs8G4eYXC3HIqfD0mkcFRzmPqkHr1ZtkEdrnrR5zLPD/oEGl5UIgiefv
GjHMIhSKKAd9cRjQ0IEgcNeRNy0ZXC+VfVHgABKlJbQOoEDQTvuqnAW/r4Dem76IXuXSaLZpvVZR
d2i7Vgl4SfvOPm71bkw73MzAiWFtR3ErqP9f0ckUi2op7tsneFaAlAiuD38jn3BhC0lvPLIncW/7
7dKZSNaui2zcR16vmG2NKm7zoqutBq0Nx44ys685SlWna/i/bfNME379fHJovu6GBg9cNxthm5jY
+bOa6YJySwKJMrt/QOAukoxdG8Tng/y9MSIUyE2Uk5XV5cW24hy2bOyAgcpj90wIpysFMJau8piB
F+MOWleu+2ANSuVFoApZ8KWi2ptn73LeLo08TTkgsA1jHhMWcWoKe+CA3yu+VSq81sG6ZPNYxZNc
tB6LnqebmpFCMoZZZBMzqMKdbJd4Ou0uuPls6p0Wc35rqmPiHFJxkdX27A0MDomHrSK0dumriN4Z
vtYi1Z3llXDkhdNcAlDT3Kek1OZpux4a4hrjmf6c6wH20GSA+S8knbGMZTMZNpL1/ElVT6ZOKGQn
u1j4nLVE+iJrKUY/Bkm1Vz5OPAj6FYDfxeCwJmlL7J4vrX1phVFQgSp1doy3U8tIGSNC1w141Pnh
o1Cu+qXxFYspkgDorBL2QI9U4PZmPUW7On+hj/QMe8B5/2itmLZzKN372gzlzfQErCF+rIHsEHKr
ENIv7N72S1xcS2MffLyCLqXs1SaEq12+9GZzHDOzVhlf57ETIvhuRgw6iRQ2KsIGKuJydm931vPl
ILsaz0VyGlLTjLmxuHk0WHFM9bXS29S9z47vz6TAGLm006P6bUFMSC/+BNjhQ50HghtuQDgNkzX6
GZj3vy0+uU1nZNTsmpLfMxoX2qHwIifLX0B9+f4o7Px1RS1rV/arvhUdvr/yg+igveFgrOFiD5bf
wiT3IcB4iVaz6tgHgzTO2YMnNbRoyYaZc8tG7VKw/TwIO+r1rTB5QPNLXxurR2+YR6KUx/ydMmTd
lWXJ/OpbpMEzrF7avdciC6Xzm9zkRYLD6HzbTZ3J+AtD/WtlcB9v/m2Z4W9OcHilR8VCLSLpRUjZ
JHN3HZJqPzzpCnIjKQoGdd6K1dIcc5LOoSfroj6b6qRRAYRrz1l7ku905zehkr4qT5XhI+kFcwXv
em1jSYslyjzUzNEmHk4H5E3hrCuLje1fALKG7kNG5SxF4Kzn9dLRmA9tNedr53GUcgco906b7LZY
LRFiYjahe+kNGgoAaFMHyeKgBpz+KEv0Q0aGRGihK6B5aujHvhyFh4xAqbefy9Aj71JT3ieYIKMA
l5reyW/G6APPGgWL/VF5DVEyrDAUFP1nrF5u9yYbuSV9TZop9nw8FtIMxn3PLYpkNzHJFrfYFTvU
RVwa++roCtAgPT9CyzIN1Nappyw1g49UsrFoX6yTgBRzzorDdwZ7RJfyptg8xKZWnH2iCpQlFhaT
rvniz+rhZr4BGL55vMXinn9j3OJWhPVCJZttQtLn+4uopCMtAhyKi0F21CHhitNRS8Bj5mwmz6dI
ElvN9sR1ydl8wtQtciDNiN3Ubt3Xyne516iMLyOnjLYCyPZqnJX+l0BK3AbOFKg4LGVsGWVvDwtk
n+d7Dae1DkWqZFF+kJDrk/JHuVPH8mZeGZbJksaWxtJRiCPslkG7rBYaWpx9nnGdvYKghI4UtW7H
7L7WM+yABqvVPo4hjuwsPlP/Uxi9qL4mPah3b3yuNFLY/SBfWT8MHjb1WObeuYMHvpgqS3pmwU5c
JyUoZnpz8QMIh/vwbqaZBmYneC3xs8j3G9TMfJK9H5Rgy9UFgVqy4aoMDGLMHAYYJ0lAKrqXl+G0
VgLi4eZeYLaKed/aiPrPwq5RkNE7gWbdE5i/52rJgmJN7NIYdeJgCaseuaF3ZngASSmWYUqVKkWu
7/+6we8D5ZCxJqfPF528OxqM0E9A1Kaj5P6Aa/Nf5JeweWInIvy+ABt5GBh+R8gFCJp577ZMXOIg
npmmFwCIM8yKrrIARmY7rwJFnAlWMEBArYwGF+3JC/xuzI88iFZWgY0Ev5xi6fURYUFiXYqoyIAL
TEPfB52eoMPgzDDFcKEO1AXZFDAyr/Mo6XzyUlK4899XM167MnzVB1J/+OB4WhwzTNOfR/FbLnSJ
F+zUcjQShOxHcPyQFoWy6+5cVcx3mPj4skmox9MQlAtzJYr45cmihRgBADAwgo6kZ+nyvZA1bvuI
f01iukeBuoHn1OTNLVa1V2biPAPCZ1PfbS/HR8uO637E/7mH9gJJ4su6ewdx1lFgwDGL91d23h9O
xaknP+V6GPI6v4Nz8xVm/ngFKorz7RHZmIWNSBa2Qmr1hY4iVrj8zUMk5vgRhxT7Ih5Tdgj9HLEU
ZVOh1E+kCrcnQeu69fBGC9fC40tci/1kxqeBBHPd7GqpxnIJb5s3q6T0kq74F2T7HrQ29iQw+E4K
wo+HuITpdpa4ks4pYTmDRX2mV/HEFNLInbLTSCw07rNAf91j7MysflW/jJ/6uKmhUUPYcV7yhPUF
xkKeB5lKvVNYVH5BRfx3rL9ywottw+DYOJUXaSWoVMuCylLlkzpvwr92BcQW2bicl2fuCHr3e2U5
fDI4SLfsRUsABbGwZBVEm11hbFGtq8IfUFtTRzz2xCemZ9pF3hjGHYwRuGKWiADM1DzEYEgtP/V+
CnBjTTBP9QUExVXDdlUBaheBmG/mxShLgiRuJ1h6QSCyYQ3QN+US3S2bvSPlvdRXO4hAdxXNNnlR
hHEb6mFqzd5gzoLZZo3/on8xPrbaUvKsH57I2Ee7NvdCqeJmfocZ925GJBFdSOLj+rPZFawQ2oCA
EVF7DjGQ3RjXnECNqNbvrKdi0HeZkelf08gm+SyMSbkfgp+y59Cjv4sX+4tPlDNymO5X+sHO6IyL
dEVdOsFNdjxqixJq5Ix6ux3Cvh2absimQ4QRavHEoF+39iJXvjSqObBId00CdiTqSZjHbAaNZWT/
APJrBuLIlyWybXFA4vUJqNe6HlHk4cw4iW51fqYix1hMcexqVtAwZLTbheJe11g17dgK3jGPci0p
cZaUoeTfST/XuPkKR0mgWWAGgo3UTTtpAR6jAFxeCh6e2INmzMeUZFp0ywudA8bnrUFofFUlUUhO
IQzk/psX57bKBFnwzhB3yl8sNFaCrApazouiuCRD/gla7AkZKnSBTY7cJCJ4iK+OO1t+mtk2XZOL
M3KJKW/t4W4Lz0Vcq4hlFuclZMoapxne0FPanVCsA90XKYrYHB/CsfawY6N992PettgvqnfFtvPJ
O7whx1ePcAMHpOR+Pu60TyEOapyZL74bwbKgeJzhMCgjDqcsGz04//ks1c+M308u/4OPE1FSBCoQ
nazxbHGPZ/rV+XatUHr9uw1ROVdTArmf5jW40HOv4gkyWFpWHrNDo2pXQaG3T4VGZWtEqze62XSK
OBzBetRARH332WxJQ//3lgAc77p4QYk6poL8C6/+xLOmm6c72NKH37gRFT2GsNNZM4VxCyqSxQOV
HxkesqSSPFSyurPgQK5FssuRloNbtHWKgPMlnElxc9/nwiz8TU76X2xml/46HxdQb+ug5cEc/3xg
lgyR4Z4b6lom9QgY54ZutnC9QidXngIhIG1+8L4Hvu1Pqs7t7fYGVdqbyyTfVRo1dCvA+FtxXydW
1tXJwr6yrTttz/pRd3nU32Gr90WIvZZnnqTpd1oTBpaY/t3WTkPnkYTAtrfTxXFV5i381cHlifTD
lgcvAIGm7azb6YwgHw1Wgm5k2PjbajiXdykI4Nv3QKsEj0iQI4hT77zXEv54P/S1WLT8nUHPcGWM
cpcHVnyUHkbmdTxGUAOeawVWPwoTA7cEmakxAC4kWGCJpzK94atAWOfqv8pxZF4jVe1kUYyMig/I
OnoN2ZByUxj/op7XQsrHnRKBHEBKV1GWAXWWFl0SxIu1K550XlyQrYlZTDO7wsXwFtQ5RkmvdRmG
+K9VYQSsMFmYbrWRdMLQ9QCmRXig1IMYwQ4rlz/mUxkl+kVzkCTbQwfCIJofDp5DZgfd+L9Sdout
1ElqzpzK1gTvU2wgrEUljOJ1CXnnDRHm7X6dwWD5ikAwLqQ4bq912UfbG7Ao4adOmK5Swxvq0rQ5
7ebzVTBnnKVZZ7n2RaqVmp/oKyQqzHhVuagt1PdLkalcuDi2xrOFCiuVzKCTxkE5dhWBVi2ePUIp
b82zDstJPYEmwM3z9taL6pHiuDe1T3aN6+xHwrYdzp7B4gXdh0MFCV7NpXkfTp1wsCBBepMhOz3J
XoOM4xFs1fSmzQnTPxaXMTTv0l4HG32X6qLUWWj1HrPlgcdLjaoAdrmQ+eGL8Q5SiCa1sQC8Eli8
QhPr4Vvzi7M7I7JEJBQ4HjjPXgMPUpfd4D7OYvlkkmpZ6r6d0rRwbM3r7zcq2T0KsIP3C56utMdP
FuQIU0nTlr3awH6H12GODnE9pfFXpKW3N01840zo050k0AikOFfz044KyD5GLtEQURtS5gmuIQTB
ZydyReCiSIhaEnmnCqhRDvwNox/AXZEYDYIvZBaQc6igr5Hp0mkRms77NCyu7gS80Zs/6a7fHFNY
SG7mCxeP9FjiLyMTemc8axB7nbzDHQkNY7rPB9SxI5HSFboKoA/I05T0Oke+rRlNHJ+0ghyndICC
r9J4+5THNkKNv9pBxH1nAoL4WqKWyyozbcE+CA89yaQLu7BztgouVAic647dMrI1L2a4P53lpkd1
pdV1q8ZWtEa0DGIQoGV/28FBsD4vlGkqdvYhnxtp1W8lbd9YHk8Xg/u+LvlaBt9iksfZTOf0qoWK
6r0OxaFtE7PpkbnG3zXycgK/SFD7WfBec/trDbXBgwzkSEGAAzP2CJ9nIXdOOxXnssGVFswkQD+h
pm2UKYoF1ueO1IWN17AIyCs7mD7sl9dGonNXlHrlVkg4u3qc9Ky9oxb9pY+P246gti2hjhBbQv12
nTiyo9CLo/6RAgXgWsZaNFetepK6hRqYe3uKUEslWNznh1gZgyO9ptiH/Rv0iNypD79Fkk5bPhAx
1GzNOBDcSZs0yECR6jXDVxb416kB+/TUjkFZ9rhl3GQi7qAqzUVXn8L/GsuTLGSGMQ2skrRKvOBd
RiAoRrfyx7SMQdVmNgh5JxJrC3yu+XJBlvUKN9PFCBK8yK5kwDeofEoV0kPiVaPylwZDnLGEiSMv
62C2KQBiCj00Jx/0f0xFSX8/91S9UbjVPEtJRUna++cetnf/b3m7QBih/+2OZN4HOPFbqtlFtIhl
e4EhicgneJeUKfdE7gbRUPluErt8M5D8iWtoqGnWR/y+gRksdnGUnpRxV+B0IQ4VLg8FIT/kkxDt
4iPA0mMyRpmOGfE+ia/kNSwnzcSOVa7lGJTKvUleNmsNZCf2ahjprrKHfuL6+CnLn+RDW7JA9EVt
08+Hr6a2rBJ+8qC34KEeYsH4bGpx7HZ+3Qk5EhZsQXhgbhvrq50BbrZ5/6UAgZIbUXg4ZeBbvCRc
3mYyIv3bv1cqtQTGFuPSUVZD9jFdhpCZpYdQe80QJHLRLWngg9egAurjMgk07RnPvg1AuaJWmqK5
AYQfKvYoBDuLPAw3g141VAY3Paf4ppkDUx6b7qVKbDGN61VL4kGObNICeoH+HjpWqNTgXy0ddoXo
jbkMHxw/55TNvpK/83reOitkWmANiC3/i8dEy/+S9K761PjzgX4aH5QT71Eor0IV62nVYpKUc1HE
SOaDufE3s8FcZC6hYa6LncOaKtz2Zsr6ZOeY7/J3oOHO5c9RzvNJxY82s7ZSh/NjwPYnCBEq7zF2
k6Sz5oH5HsvGbvFzuG2vbeZ5WvQ/YFI5S6j70cqc6SK8i+Y36kN0YYAmCW5ktrlR6Dwb74DTc+pX
2WteFbkrPo9anPaLzTTor3J0mUZTYEIUVexfbYzeBFaMGU59uPkB0VjCLWYoMvE2giWBaRuHJKbd
E8EYWZATXrMNguASqH7H9JBoo/JurvRsa+9puS2yv5UUw+kzN4T2Uz/Ghsdo87SJ33/OzL+zZ0T9
N80G5wvC+ZQyfq1P+OicnB3E/Q+RhKsOSiD1PxLtwrCLT8tBPK6jD0FREpGc462bdI0BZN2Cuusp
ynKppnNyALo6b3W9dSYZO23JTmYUgY7uU0AGyEgyBWCNsMHYNjiefkIXS+F+ViyflYT5ZPl1ji+l
PcNujkI8opCCkGs73v0VgovMn3nV+AxIaQR9aI0FlJxE7dRVuuQTzDWpoiSDLeidn2SLGzcbk15i
msXTlJpdJZa8JgLzdQVOGUxC7pf9hkhoHB8bqCnoX13Kzpc84wSrkwleJ0A5QKt6F3AjJ7G4+No6
1DtCcR2rbaDknATST7mDOYsRiSXsfgzUlpGQH8CnQPS2TuDhZVcZhkqhWgdwiTOdEMNE0VFAJUll
CiEfo6GnyaWjEohOOvu7/837YR7C6ke/p8Ehz+AuPLmzFfu3Yj/+JpSyDY63TX0hl2fisT66PdBT
ZI01iMY/0mCayQlIZdoIpLxnTR3xzGQXNRRhzKx807AzBKA0lmris8E7K5WBgrd4VCGXQKK5hxy5
WkU+JVvfVGEv9fE1zmC6CKh8Tp3X2QX2uqER8hIjH0/x50XXsj+oiPSNjs4CmDZ4rOlOg4HgtMMb
wOxfI3KDehlf51wz4InuTuoadBBIHvacSTeHPCwO4B6FcL8qsV64mOLEfYPuqJ79V2Hl28gMvftA
w46Opnx39/rKEzfdB2wYkulecVStOAPSZ0YSJmXUVX7UqXdMrbrviTq0oiEV1RFuURqqarg1I09o
+yaBM5hC1XPJ7lAH+0bnZnAD+tntzez78N7IaYZsHKVXB2i1FYMQtIrClu3J9j/HycsNwv06H1a0
Onf2zI/TdskqMbnvxaZmXqUlJem8sG5yfY5/jxxTyv2le58UHXSYwzLOFv/FdcmmRGTtNImhiYCl
6QicubRzliB8tpcTJyupW6Ijt7FaevOvLco178nbIKNWSPa7br3Lxq20/DVMapfmweFq7BbXrRi/
883gC63/w41/FgOTp07+HzdmTrtXfcKB0NfXHN+xNYH+fEasXk3SnaboPror+cGmCJi0hxejfw9Z
VoGnlokk5kToLFF3hV3z61Hm6cWjR1mQMVcMx83pNth58l6P0PgT0vZJYnYpDuuA8c8A2ZZ3bpMN
eE5UxVJDXerPLcdpXFQ6avWV9xdMDG35PjZqNs3NuvlDrfdmhkpBpskiuM6Be1py1qaqBySwMj5F
pWQM5aLFDeDN8UqGmjHv6G/OrdIWcgw0+U8NrIG5/PzedG8NpEWqNTD91Y+s06ftpo6YRWOSl5HJ
TizuS0r2u/Do0joAHXXH9wPhCfQYZxsSFaJOtgCxHrpkjcvOMfUJqAhEcnmYKzp0S7Hv4nZEMIH8
IKpqh/4S6RtCpfAaxnGPDprRKovgWmK1jUFbx8kMEqTSBlq7sZuyt51MgjwmISqiPqt0ymW1tgv8
b+BMEHsKVx8YbuWBdaGQF9os+Q8bewWaf5U7TWPg5UFldNGrz1INVDHIT+JS5/Kh5tJvrkIBt/ZZ
niK6OGN3jdryYFd7+54eiD6xgbwPwYm+Pz4r9Ys1GKjK7jBjvuG61YJcuIAA5EJooZsi2DulR1QF
XAi8zsU0PghFxQ0Q0YHbLTw3lRhPvurBMwpSF02M75YZfzArS1507jUSnwe9tlzu7LrTJUBq/hiX
VyGJ54Tc8ukKQm5iDsOx1XlIgeaJoQFBKVsSfk4GJ0Q8nOTL5werhSwBEUkSS9l2hjnCw9MSM0IG
mId/P6taRX3FVAkiN6olnou9NidePRaWZQRffHOlPtWJW/2GW+U1WWgr6GjzpHRInGfe7eWZNQ2q
m04jS39mmvTrRZ+yg7TlkWppmwBbEpG2Th1MiUAQ8QRf+TZO7gbzScTEf9rJ+07PdJ+AyypgEiu+
PS16vNREgYF+f7/A3B2GQ0JsuByyQh5LzEkl7OEAi3T/CCvT1J+F6HuP6eBvQmwhZPBpYwN6k1G0
/xJSnO48RRIyCiQ9ZUaJCSA7CAfvBdAl+Fjs7BSOWEycx299or+1snz38mNF02lSrOkgHusOzGd/
oMPTtpQRwltgCeQJizQOLYmBV5/8AvZRmndhmaaRfmuKXOUaSjgMv1dHDyfMhl0PWQAc6HKaBVsb
dcPObJERC0w75SmWhsdj5B7Cv2RPvEAyXvW+DW8JLwdcrPr4wyRrC22u/3yMCRZygIwoPo/xJGja
1OaS7exFPEVYo+yndmSJZ77pkqlP79wt5SzxSfPlnwBO0YC2DPzkViy804y9Su3aqHrYFiG0UrF8
k2ieUyYfXa/fevFyEK90HSHDM46QgL0hH8vJfG/G+WD0p5ktjYqGQ9xMtJvZfAhta7Jw6BYxvC9U
JPnJiA8G9CcFsUaYsLcDXbuxK3HHpa/8d2Ltb/HOecLZuBpv1IqCbkv0LclM3FJxq4dYRjC9Lh3J
CuvcG4AEGuXuQF4x+PX5izilMybCRp5A1BBlUQR+LZLBrz5JQTpBuljA2S6J5ysElvk+b666i3uk
naPpQsukhE56SLNXYsqciDN38c9Aa2FJKFYhoip60YRZMN5sRzQqRh1D4DRyYfV2mvMDAIkqUoLF
7pbierf/DsWQb63gUikTYdZkbk6ld5h1R7q5C51kDLuKvSGRVmr7YzYLJlf2yaDEcIG5bsmrIAwu
HrXp5dasUEzJo4oIGMe06WgfKYSQXjZH0xchrrncrQfFI5Iqk52i0fZf5r2Wkpn1M3VscfaBGjDo
UyHuCWYE2YzPhUV8ck/hD8uEBjgDrHtFKaLihQ/U5ziBoXO7Y+0CVpySa2VbIsRgegkxXpJ9fZq2
AcqPYMKkjb9BuqwpMAu3tlCi1YtwXyomJI/upEHfPQmuMgcbfv54a8uo+UXuQ8/g6xwzMOjLkVj4
pPpOZ7JQFfOVskG4IdHWachkRXcdU3oLucsxvhEXEKy4Bh4HtZDazEPWN98prL2l7hPq+YkS7m63
msJdkfl9iXBKUlV9U4ZbDoTRage8/9Z2UJoFfUZPhdD1MzTNdSNLkYLEcsKGDMcktJxOJmfto7zr
1TGwn7qXf1H5qCXaT8M/I2kefCTuLyeg58pAFqJslY6t8R7LYE77b2PbbNjMf7RF8Qe3lKDJlGIR
xyqJLC2ZbZENT/Fyb0ZjVzl+7wZmacAYsZ/aj1OYb6zmWCWvsFfYk0Qv/3DlwPzMPNdlRG7yIOp7
V3/kIkob/4jNJ4qD8lkHE2EmZ1mFVmnSRo9Z99xtKXulVIe11jJIRhvzYp+S+oZACn3/I2SjMk3m
j08oPlsufOafNy2TEtDk1vRRUJhaiXmzXQirqKKRp0CFac/nXH7+QzQwmh2HxeClnemhSNGbMCsO
PkZAew5r9guwn/SphUuMnavzLORuuU/5WED5E3Byx3NIMB2UTx1hX4p963/Ikw8ilgjR9BcbxhKV
u/LGT0KfMQvMM4ZBah9tz8Isv0kEeoZ2Kzw/iVYxwOL6RfeWR069P6+X7dw2C9xkcy+awMjCBpb3
XqG67MnU5J2YNBDJviU9EB4wFnhLfNmz1+XlMQ/JPr1bsBPjLtmoqwsXXwlY/9XFrN1jvIzV0+gI
cIOaFzgOmLzZRsmGQdPuu4d2ucG3w++l/7jfn3jr4wMRYW7MnZu1xAb1sewDZik8ZG/NEOfKcwF3
CxsaKZduCQyPYcTxvGlg0V9z0nwQeMVJM3KZ2q2GjpxfW9dOXfaQcy2bpfLHuyGbqARgoUxdkTrk
HUQLyVH2+Minzr72A4xaiEzbsxb/xvIjfY5IlocaYDzgqO9aaga6OLrV5hAC6aso8x7FgBgntFmA
kAhogl3BodssDreG30TBQ7HMOZNTJUrRfBNIw2fu+OgmJktFzTG2HIc3rUXe2gQs9D7IHKguhAG/
Rdb2h7AuZ4Nsif7J0lTBMc0bjpX6vZBOwIE4yETWS4yvQPnhfZc7iCY7JDFGmdg+P1zwnoTOit3t
WU5rTNTl+wc55sW/LeEWy7Zx5uXkyxwxMEzrIWIIcnXD3T75ATlWt2PxeBL1oKrs+1UiUlWvi7ym
aBW3P8BVoL1EtDC+5ngESBxsRdZXaTOZiKGNHKtcFVlkwmyf44Dh0G07eyEj82u1vereNu1kL8/6
IjFY/Erb2ZBegBRKQ1FLyyakGRRS+WE6OIcKqiMr/aSS+T/7dxcfLdoTt9NXySv8+y3SgyDQ3Id0
krXkgkTzXwfdOkFTKBHJmatmgLOpZktV9wUWWW6oBb4qLkJxQgstZZ4muzVas64bBWfAOpW11czz
grxUWHZGN7tMhlVho7zSQRf8maDDPdJ+62TpJ1hZkXCmJ0vbihVbb/s7zuAqG+PTcKMFBNK/sDh1
54tUiUIzanRKW3RljMkY3ImUU+JdehDnXDgHIiMzMVDBZsgDy9tIuMEMA0C6TAknTgCQWdoohSXO
+kQ8h1K+g0qaH0ZM4e7QjlSaWjqows9AoewPsV7bnqABQYwUzhMlE9l6TUNN/CstNefwDGLIWLKG
HEtjrFYRuvIAYklsbaRXFdE4IVnk6aCL/+SHf9QV1uR8uK+t2AwUeAz5pc5m9GY9JPtZrst3Xgm3
8QUcHi23FrzZN209lvXEy1EIl4N6nuxu45qvVw4KEGt/T23da0KTgvEd5yD+Tj+GhWN4pePmFWkp
6qamQox+YYbrekPwM3uEBNnSGqae+3teGuWLide4N4V+c2yoLo2HDaP9ZWhC9geoyM0DdaOaevPh
8EElYl/AkWPpH6kteDL2PHFtymd1V07ezOBR7i8cl0fgHCe4FGzQusI2od6bpv1Z8/E+Kmk2i3sg
YCWRi4s1NYLJcaRhc9RrCdQQq7mfGaXsfA3WRyDingnJYEI8/1wTVtl709A9o1ZpfKQFVoFTLQmN
La80PaCAdZsIOImGOkJPE3EGazy3VPCMi1BITCV8vrT3soN5KNNsNnvZuGa+F97ea+reXWWk/yLL
D12Ht5ELzhskA+NH4s4xbtI9d9oVuf0bLf0yFXe4laRbfzrlPnk4/C7KSSmpl8lncv74W9jFapWU
OkBIcT4yuTzRtMA0jTEQ69Qorp6dUUXQznDtteoHj2X7GqGdTkYEgXREWKW/H8Dx7XlG2JEhnBPO
izZD1Dc7expZNDbKQaVl+nB/kw7z+vEUwqXnGLrhQcMpSelwBSqV46vKfQvtjlwPKCzi5YBdV7mp
XJzftqFFrGcSuK0qnOweZvS95Ez8ZanZUhO4nAMyuPad5Wg7ufAkluo/qdgBNThZ+BD32mYdAkxj
fC+0y9qA1Z+Z9EmrnHFCNAAj0itE6yE69M+1XvTM7bHJyD/9u9kFWVViDkU5CQeEjFJpqqUvMLmE
pTQ9q8uNlMoWUSUTeirtEAkApKcQWrZZCCeUBpRTNFbsnJkHmTAGCowIn4RCK3HRIGitThM4yKL6
XBbMVz8OGo1m7sV8mbexD+nOte6JWGK44FnncsWlM+PnnA6LcMpCgwnD6WXYeO1wGf6uq88oE+pe
rkfac/ILkHwTYYZISScNQWQmvbiKy5ywfzeAWsFm4U+cyxkkd41rLwd4gaj0DTm0Ty8ZcyLRxRyz
HPF7Vdt0CEEePXoZYZRpHjPuYlsjBQPHvJdUcfOcxXXjxnMagOAxqh01kOv+gBVYetoTL4HoNbIY
LWX/sDjwGeBMlWd/1diIycpjBPScBLqcrVEn4p//FgwvkIJUphtdRORz7ut+pKaBiqF3r+l/QbkE
vxES7III2OjnwjN0K7PE5KYb9lnxxdIUOvOHPVQI91h9x2pwq/8FOyNHqAFUYF4wAIoSV8w8uvkZ
o777zNH+n4KBCHLaW31aCdg7LRtHz+G+ZVa1FlwizoAyanULcLobDe1fb2IKxO3jFjMRtsB8Qbml
TRt/9ZrLdiald5nEZfOjPc6ohAePpExB7fzbswOHsNoDXljQXGaYTIOt0w966N5EjTPV5LEGdIKg
P7JooNWgIoxV0Ieifpo/lYpPE6ugQ2NgjVxjaiW/9FnlXhViHQXkTwIcKql2UtSLD59SQFIXNFIA
BMVX3UDDsdt9PrIoFS+qjrR/WrAWqXftrEe0PcX3ovS4bpv5n9iruaRIiTCJI75ZMBMbWhO9/EdQ
jNkVdPBcy4k2bdFIGDqWXWtx9onHP/yZzPyffVXr5i4UaEbwbLyqVxaDbfNG+nh1B0e5FxHAAeEf
wl9PRKGRgoRm7DPALLhfqtttEG7D3HnIBvbN229x++oFtcTUfM/JNxEqFZHeVjo0tnP479kCKHC0
z8mnVKz1Kcw+9Sm+JocXG8XBnB9Lt2r14KveCTDzkVYAG+XPZ7ncltuF/dnQy7B4uNjfskiBucA3
yle5QU7th5XukmfZ+5xJBoRjlDjbhQ/P0fYbIQ2E29Lvn+v8NdQLoBoZ4PHijmPANJTtnWW3PCRY
WzfOD1/VurjzYb3MQAgizEtUEfCPdQ4WIpdV2ue3QVESP4js5nveBlivgl9VVHFeP5vUA82SdtrV
bkrkXUdZM4Gn3JLd6gc46X75GkGOOQ6Cc6xQBzNTMyridMMakUm8m58pNTVD+XAX4RGZBmi50Brc
e+NL7ZabNAzA9vm/jMMawQ6lsS4McHq4hzjTEgFRI1AgVBl4ojrLE5l1ndEbfbCIlcZai9tpGrCA
nHUWGRquapnE/8Ii2zrVRpa29dt7eionn/BaoMsy/LHB60eX2Udwn4+Ll83vPHr7bo/eqAklGlvr
1sMpWQKHwqJjdr5p2lyugkMF1RP7ixFGvallvO2F0X1qpGhHdTODonA1x7myZ0gJdov9VmiEgIF5
d7V6LhC9SPHLCHrsBDRXwm5eXM+NLgMi3111cqVJcLgGoDsjlYJ51tRW+KHC0WWGlTXUwzxewV3y
qxmFXDGvOA2IS3U46jGX9W9cOTCVQI3X1EyWzowCIqAc8nvu9fWykvrDlMfkle+6EM7o4sIfvmhH
NS3Q1vXo94i38brfyJ0yWoBjBmeOm+IZ7y18MxNsCrJhsWK7hlFZv2FcWDqPUkBIClW8Q0xc7dGk
k/bz7JS7HtSzSqBrXe56FWXKjEAEGhhmpYJ7PneNpfM3M7svJHHVgwawJJbslB8n3c3JCJZh296Z
OnRuL/64mXNDKACxYkxU0fEOdbdDjnbkGul92lsmdzwtv8QCnJ98G0n/tTYVN9lecAfuTsETVTbD
V2kx2RQV7lE1OmDQKvtuIw/rHm17gVYRfPDwS8+ABSd8dxrJeYZZZHr4ZNxvE+3QNDewTxcxkWgl
2ZmEPn+Z8nmZu35LBJQlu2jNBU42ZNRtdvaJUIjhAyXqib5ApDdTGNz+qn9didHb9/4grPurM+je
WtNbbSM+NbDMkfRdDMrFgFcx5eScqhECIRsAHVwasSmiqr9vhbYMVAtTvgt94HUncJf/McdQJkGo
g6hHdjdHHB6Lj+IqfxUUBk6p3ETlfxABIVDhhe3PmFnBb6yu5uPYK/n0oRLYRpaLpTdzOodOj8px
q1GXEQ1T0z46eGYCbUMOLV2P48mo4YHLVZgMxpzA5VaPdNj4Hq4oJFGnvpPP0pBOKhmPd9RIli0/
PzGUDI7f1DP5YwX9kF0J596AAef4ZnntMnD+D0HJz+ivs/i9LfMCdXG20hEQjcy/9mZ5KAJN6q9i
hmUhPNrNEzC9AWlHIIfhf7ONvmqBhl82amd8UgGVt7HIxnWvYXq7bq+U3SM5JLf/pOjs7dSWug8N
fDaET4aUB3TSmlPgX2/PyaRnkSopf0bXlH7TJ9O99N/tEQ4c4KETUSwgyUw779MR8yn0wx2WOuna
4PuADEwDB3KSZ0ShMjexAeZ5M1Arnt6X2NGQg2Xd3qmbG0vHR1caWo/8eXugGEimiVcmehfh7rbg
XLehBMQKOIy7eiTU5CgEJMuybsKEPWBOg/RIQqi4yxT8mLr9Y1I4yVnkdc7bq8UdYwcovAZVXKO4
jZ06sL8OR+uDmuqlJNbHSPFFMkvL7djdq6VZ7iiDFuaynbWjlnyMouWo7mDlQOer6plKg8U0swEl
++/cua55xnVb+Mu6aIn025ylI7MHzf4Nj+bbTfypRv9r7WCWtEE47ReifsswxEyV4y8GUjH1EYIn
y5rxKx08nyIF1J4er/A3Q9quKIsiHT49DOJuNTzhiddFqwZhT8ylAKlYilQlSn2vFmLOo5U79lsZ
QAC3XU8KH09qMYEc/6MLlo15kTQdGeawGhTbrin581p1H/Xr3i0wNLrp8eQt5alpWInjrOLXIx7N
4UqsbYynI/cTQjG1fssftp4bF6g1bChA/GjCGmAh/whlBvxIwbljZKDprdeVIOqtBFMhvUAA8qcl
37umyjw7dlAzCIOFJyvazsxW5UxW4k083B4ujnXUhKs0AlfZ5/eN0mvT4gm2gCxNvGAbP8eihufk
Xr1K9N5VenQq3vCxwP3jUxB/KQYNM9JYkiVL5e/1Exdl0kpiBv63Ae7OrkZYhDhFlflhNCZRJOKz
oGDkq6sdteT4z9K3f/lnXzGb8+6EvnExGMP9K05jF+9gwzW9OsYWL6qpCIIczMbZ2Lp4PvUB4B/W
vidSb7v7mHG4DlVu53rCgpOx67+xqK8X4wVExzKZhyJqzDq0YfHhj2PxmJAgYd3jQLLLKplQqBgr
uE4sqGSFXWOpEKvsNCXjoLloUQlOdFZ4G5baDWVHjPGk6x0f694B6CzWycgBQGvQ9KdbRf7En0UF
+JvgBcgEzK05bXW1JCUof4RIOkCL81T1CwZrWHX45M0ErlU5zzr0+6C8VNNSS1BVy9oL8mc4GIKh
vJnaG4HEQP5eIk8eXAeTLA1LHaUlxNRJjMRP01kZ9N+Yx4S/R/G4jKC3GJ12H5A+OmGdqGVXAsY1
M8iEsPY8op+2DjH09fiRg2wq7intq4kl9lJhV4IMbL0F4YjOlEyY47wuXoSufu1dS4dJ/VRNtPuU
Acsyh/7pXynI1yIBqOuqmvTK5ipyUR6TRnErm+bPRgpi7uhJq5aMBCa1qBdVGHMI6yLfCuD2uGp6
lBiEYq2aOg6hO0fRZm+7fBaIdncWD5ech19PxQpT58ok9mGsqlHkY4/y6O1kikCKJvFL+DdbADLT
w3W3I6RSodSOQ4DzS55C1jrfMA4M721cdPYWQ5SPn5j8RL51hOwYKbNbJzcgsMOECCpdpSrrj0AX
EmCfTMEOmjJn2MFFlT34eqgF5WHs7RdXJyYe4aaiInJ3UA5IPg3vGS0IBspw7KP1bTB44V9ofJO6
0syOVY4XpcT1mWechL1h55pSOrUVf8Py5SsXNFxUMkxrRi50iTpKAj4zBDQTRVUdVLAZ8Y4crR/P
1lWEgC7vA/yeW2Vyh/KR/jo5b+Q2wyimeG6xU+5m4wQCdHwS0lB/pjO5UrTU9GA7Kb2x4jSzq+dV
mUJZS+x0iHoEWwHwGoeF/imac8T8j+Y8/W5/3VzQXXIiC9pU2deiyfW3ZGM826awaocAvmv1ZWXp
F4Vft3hqvtT6NRdQ4WxXJqmlucLi6TE0QKQJWbgjwuNG7Fo0o+GUsOlL7GP9g3dQp6tJ6Yi8FeOt
ODG34umdM2DGf5ZQ4HG17QVGiDqayCKAyw16v2qbomiQbrFDLrbhiv6lfBVIQukMNd9DJ7/UtVU3
+18cR/c56iOFUQJzas3nxoem4WmnvL541Znyc1kb10G1lRUSZOnAfZHIAIAdF0MsrnUzVoCcrdY9
4G27XMOhcIlrvxOhxdQV6eNpfgB3e21+ck29l5+lTPJ+G+cwTBCTWX2QEhxtzD1vmK7vtPkVBBn8
Rk2vUGRfvnisF4j4kQ0VvwXjekWFTKhpoG3bF0qAjK4AgxGUzoftunLGxl8hEmUMZKpaoE21d/8X
MGRVjIdoK0nQZr8pTrlKF5nybBBvnXK3AA66o2rzgwrwF3o+yOTWEuHnjO1sY4iAVRWMNBAc7v2o
IlKyaYlXZ/DneqVJdltANo8Je0w4LvbrgoqGew5ujorTxU8RmCG2MYvbKc27xPmtr6Kur2OJbSHe
CK5WuEnmPD2fgkq9AN/yueN0KSQ2dl8x9m/qDoknPSF1iJum/e33AGqH+ysEg8wW2q+7S5T3flcc
EW/3fstO8zud3+UvYQ9C8yxDyRH2x/pGW2gpKwo0IE4V5y8F08zFC4xL32zhxgwk+7zP6Ll99VmM
CqN7wWcNpEGNznPPNfhlEPqJXvTsMs8GpNVCD/TlFE464W+Zmh7imPeXhq2rvVe6jXKH5BoK2y0e
22X1ZDKV+44+gw5t90QDh3MPyn2n8eiGYqvWQ3lMGVIlFX8XYZ/iCjmYPW0Hexb7IbPV5EO3S5Gr
GE+omoL3JiNfRkejTExaD2XwHXNmZTP6GASLffsXuckhrFYOCplKNUhKO6YsuSOEqjWwpY3aNT+9
CSTUAYLR4sHiw4GEyDaCaabFwNNtyDXzmIShquJzyZ+TNpJe3lGgneD8AKgxJyO4yEBCX6wWuVss
RnD9ygGaiE4UUnYiDVNdGzZeCT2EuNkKDoHCnTxVgT3cJxpsKA5Hwe9qHYx/ns/yPFbVqS43hfYM
jKh8DvgjzrXtkDKxuTWm1Y75Hd3HxPyWNz2kQFKyBTAEG8rUj21POYSrwrjJzCemXFXkyG6zx0jg
h5nNw1RD7qGmqTxle81hnszKgEStOI83ka3FH/zR2FgJ8YG385RZNTgpOyNVWgrM4ZLLXkt3Ht14
0s1OEDlxXI1xxDlsBNGWT0tL8G7pSEZ6Eh6mKpCSPwqp3+SSa1factw4bMajph/w6jxYe2IkqZ3T
JZNu1IIG4ElHq3RT9zolsfv9SdYjCiT7Md2iwNiA38D+hjEX8PWoGgmScNCnvfYiJqca3cz1RBs7
O31dwso+FNA/MjZCx/kcXXgw+bc1JtMF47/SSWPsaN4zIZJKWAmdA/HN5epPrTLx4K4Js78Q6XGH
oVz8TjEcnEr75UqCfhdlYWu3FTfW+rybj8bWCJ9xDqRVnQh3hoUwmXB9sjgWadw1Oeem+fwVEMuM
j+ivKXdNKgp5/YI8NZc9yME4NlyWlwWCVnxv3gmoWNNGgGcjE0Q9iBvJUjprU2d7p0pt92czm+Ay
wVxRDCHW45Hp0XVqfD/dzs9VFIPVRkVVOs8EdyRB/RIsT49IUMFYXXUbV5aJ3r64k0xbf7VPVdw6
srnavFNjrrf3FtouPR3blBVIhvGLxWNLiZbm6Yt3UHGMaLRkjsQ7gTshEcHsEqxM7yOssaVujg7T
/LzpFZU0d7ZUQmqUEIcBCPtCAcT+QBtoxy+x50wogcUzaVDSkFkbELXcdeHTPTg+xkpimzL8qIqk
aCgp3B+JFJuFTfBRMU2Vbn3HsupSui/7O1B9Yyzu/4x8k9oiNS6ZvePvFqYKBRcElhMowkdR+kjj
YyjzjIwYjnbRQDoR8lhRJpmkKzTHjlIWXKsDYCGUZ1uI3RDhcIwj7xFNRAFvw/Gs/LcWMUi92f3I
4z35A9HKKd0JfE7SGMQdcP9Ykk7Lt2tmyDIlyH9xMc7XMkONgwXMfij3qWJGGKKkB9LwcErlnDQz
tKB1AZvlwRp+XIuCIhfBu9QQmFpKOt/+oeFyxaQL9qXNx5zWF8igig3in62ydCCEv5nIYjUDOGLz
YnAyOiq7/dfZPFtuvq0hy2fuK8WyqbS6MzyIhQIMFWXANeUtBNdNMe/EVC9+pz9vuQsM32Oxjjv5
xHpuNV88mlJF2lBJZNVd0TlxQnn+wK2UdzseBaBqyZCF0uisGevzye+FgF+NKMhkSiRjvZTKCjvc
jBtkgBq3xkLlFD0unt7Ml2Zoo82axvdwoGb1d0De5CYaN2A2t/2zpYeK+gLthxqEu4oBBUYc+IMY
0CT3O9usvv0TR3h6v8Ne/gYhMKOaxw6ZsXzLn8tH9dgMXrhd95FNZoqfETTz2MgSeBq3CShJNlAl
XpmLcj144yAWGb+CngP8Ju48eGElInCT5cRCdTcNdOC3tGAlR+cPnjnoJKYteyU6NlZzBBT94I06
iY5/tb43mcR7miVj30BHVVRq1NfB5RwNHt45CdvEQg81D5NZeW/xcBXCT0VoGgSyLU3bxqqfropO
ehNDiXAzvfNt8j3JpknrLnWJ0b3KDVdkIarWhpbtkzl6RqpthVV3VkZPEnwiWVWozwhQdKgxuxZW
Yiyi4e6NcWQ+STUPBEyijqlFIJM2Ec9WJL7RorxcsIFVDUf3x+5Kq9Fc+mG0xaooRFsImNb9YSjL
6/jhaAmxTSWglLYB/W/WZo6gm6O4XyoKtqUYGW2LVuNEyRIM5S2ElnQqfllqC+cMoRffxIkQDGmS
ngzaHDUjCZ88BPBogAVXuhFAsX21BVucGsPduSrGU4dMQAXbMc13Tq7ZDvlWdxH+CAIf4BhIKz+N
Jj5T4vhksIeZTyOspQADnli+2QhktVVX86jCKbuEB2rcNdGld+0dsKd7dBdhgPBywtdxR0KnygNZ
g+vH+146Nj2fjcNpmYqUPVKwzWirloPszSQS9ZF25U02wUX9gw5Gu3YsclcDokDMQGYfXX7fjHJS
zHd8qf9R8mibwYmBQ0oi1EXmCN4tdKQBkTY2fowUbtUSmiir52pm1xF+UJb/+s3Mjb4uUsgBs7g3
MDNdwNokh3RkA+K6tH1eP4gHatFBsB8QCVsgcYmBfxRBu1vQkIIGPtl7nI03g6N/GilEfn2JsuwL
FyerpY9i64SqNfB08XSEZ5QLfDXQ8GEhMeR3u+e0Gjk6W1b+tk+S++ny6Ff+Z4OkCBrYAMa7ackh
bWjON4SE2eirfayAGWzO8+gLIGP3afR3I1tEuGGk9Ye6k7OZkF7LQfwpCVuTz5uRWK0UdN8PeMEm
9hihWJ2wK+E+kVQRg3oJDMc5SByuOuqhkU4MzyxW1WP6+QUhTcPQLRTLWRx5NyrkOcPgNC2Y0df5
y34LEFvwDFObMlFtleTXjlYxdlw7jG4/5/LHzyXkJASyXyhUkjGbT7qBGXfhiK7Er5NZrpkyBGg8
j9gIXO+SLrHLjqd4caEKNT9koibxC/F2Qb8UxQHv8JN0H2H8X4GxXVhTHSxWMzJqsYCWFW7Auth6
cI7A+eV9tlBSsvnD5agxOC8Ri4Pv/gna7U+deE4k+HIi9nzWE70Rp2NRumuGM+9T/gnOyl7RxPnx
e991uBAphV/6kmdCFjRdM6S/dPYF1bX7hJKQ3S1AmeokRjyen/Ojdhl65IxRcBUl/+p2jcPY7QGu
juGq699eZZR440WqRlPM76XhQesF4zYMIOLVk2cABCcSD4gKndgyr3To4Hcrgkku3Bc8qO9akDpg
TaI8ZjCELXhemfp4QeAW66HOw9P9z0jr9JAFZXK+6W8ifP16ye5rcsTNoQBRJ03V+x1Hvs7Lthtr
mgTmceaHcCc0cDba4x9IgqmSDmtf+fvmCopbSE/6Cp/GOwBZ4cidnkGsmAVx5wiXnk5qyVRmPXn+
P2plHmbk9LCNn0ulwq/RMZSmrh1IWIu/SZGWKXThzTZZilcYX9es5MeeRIj/2/hqRLhq4ql1nTFc
zgS1x5FD2sV5bi8nzBEWGec28rDJVPwqY20am2lpfPlCwRfel6/xQjqHqn/KO5vTL/98nrzXmUZa
T0lC+agpAbUSnrSS+4A91om3avcoFzJ/dZ06udcKDN15f7FiFnW2KYOAmz9tLhR0GgjzWAsxlvYn
dM007raJz+iRZLCx7CtJRpIXCgzdyuLAm6EHKOXjz0Id7WmyQrxtb+T1xd3V1Z2fgGyTMvKQ6vL4
KVwIoiTsVUbdbrm6xfBZrzBlOjLLg4RB6HNODGn4o2RjUtsGHrzgzCM2OZ4yxGaElMkzYFbsx3le
25jVoe8QJQoy1bC6i/jqjqMpY6mjUKtbJfxquFm3WOxJCDqs9jdPMUmIoLjNyAC+MRJniSCqp5Kh
Jugqa/aUUPjcc060HM5zrSTlFY2OwVFH1zt0SFrgROd3ndMi3mUkV2XPdnZn5192EinTXJp8/5j8
HnnzxnsB1uPVQtSw6TBxr0+KjmdGoXE5lcT31hnL80NWjPXz49jNDBiyQp7akPnmX4Pa46xI8v+I
jrTc2TUHuLBJxT7hKqBh8NmaBZv6CtSyNIoFL9fjDIQS4mjhKIhtNrUoLpitE6uQQJf5obWMGr2t
5t/FE2A2dcXMMN1GG2RqI6jNIPbECYDrF91OESwyHuiNEvrf5o8ohn7kPkfkbeBoVpKMGQUA4cDg
3vMdy85QT8kp0Qs2FdsDtLXKHpEGxhrdIGVqf3XB3bTLgsieZbF/8IaF9VHSvv+0bSmMqpoA1aqh
OgBz8DfvAjgPa77RhtBzGPVHqmQWkG5NcbrWNqbwR7xiT2VE7YW3oV4HvzRdZhiAwoAwCuhmiUU5
q8gg+zclk4WJspNTRYzSq4gwYKsdgtMZtlWNFW1xA/y7IvmvY7UPq0EOGf5Wve9Uy/N9FSmd8xZ7
xbL8hwemwTm/zfkwha/DTuwxvEVC5K2CRLBjMbLbJJ21B4elvgbn6wfiyLiIVKrzYcxQCTps6C2A
2N57J28LOR4CBPuz6bCKs1s+sWi6afmqOzJUkmC9GAOEBOijRNM+o2Uv1WrrDdsVd7D7fMWviJkM
1yaQajuO6R+Tz5a84ItzOicfg0BMNBAWi9Ev90tugscEepXD7dGEV7HlRLwJz/706WP0eqKiP3yo
rjX/74k52k55ko+f+8UC990z9awHKfcf7BIwUxrRGNkLCnFOXEF1kXDrDf9Gv/dzYTvqYiN/BADH
6LpMPNHsb+eVbI9bXkDcAJ0kmXlUITkIoF/M418705yoBLGcmbLBU8F3fOYVcRd84+Xop6bCNMBx
SukNVwzNJugCuLyVOLLmn8p36L+1ipr8UXYKSeAGm2MlCWAJlrSGjdxs3OM5qwyFUwRd4UtI6Dtu
dItj5EdaK642VC/8dQNswJijySghdzWdftUxzquOkURSSiuzO+kmhQnbLD7ulzlwj5gFdzr/PZ1W
Kzw7ThgTOsomhunCsbtPfXhjF6ayqm0uPnD9Tk1fHLmbSHdK85IFqtt8Jvvs6scgOXbD/MlbIxhH
XHFQsJVaVRaix2CPJwra6N+gM1KaqladZb6GRYzHZFIRLcxkw8bOVJMq+1c7ncE/cbrjQzbWZS4f
6TlYq8rE1dEeLV3m/V7qbOHFbDjdLZb6pHqTLyJXn1C+1d8lqOZs6fI7i8h7x0LT1oGvxu6bKIeY
+70C5jzob4CNewFiTi+i5ZsUzF9CHHe94xQw1jNLhF/ITURB+48FjmLtVqYptjI96+8WU17hTOgM
b2zHCK5sGLI4Pzkp4mDpqaPZ7WLqeyGGxSMAIgOYQe5/V6JeSo1Sf3yZJQ7aUdxOHAyZCJ0c55y8
Vgqqfvbj3AYeDwpKGPgnMOE+44wrLZgT+TQV9cIb6V8dkyzY+6qlnWPkj0mXhH5JQhSGTXoucHQ2
r+1E1iL+/zyCEjXal6u6KEyLHPg/NNcSpwO6jif6B5ZXZGeilpgqEsZXry+HMcskJZqLh9fpHpkp
ui7Rp7QF+oz4pNzB+YwOrEHJxe1lIxclLxoX9rN3h0InaCtgXXbNZVlJpft9gPQZ0qhHa5brTw8B
+l3QmXKzV8EphdN5uPJkfwdX3gKNOg4mQjHW/j4egCzjnHwJ+rFXDqQX69TjV5y4ePKhumzTuiMG
ppNIERdGQTeeiCDTBvATRMAS+2kDwxDNWfJSR5C4ZALR4K4MXqyzkzSJcFxt2JnknLf+J0bS4Mba
0a6DHZwDfhq3C5ASGGN5UpX6mt8bsiNkor2H05J7aeInXl7ouICVqIA9VOSTsz43gGq6K5ZI/hry
k3pw8Uz670PRYlJIbgdwpaiPPIP194r8tey0vWDwfBF0Uoq02tcUuMWNFgpADpSkmGVZQLfEwA25
yqKn6udKIDFjlwxc2gFkWSWRUHvGADpHrYAysyNkST4t5tIgSSgLIzhhuosLX8SB6wbnLaAkwOs2
eP7jIiU3TswYRg24Nus3Cq3u3R8GcPAMOoeB7Kg7B/2Ccb1Q6H3/jhSJf6uGtdfA3AkiqRQA4V4t
w7GHRNE4DcFApq6Z7Wqx2qPo5FudCwoApm9u7HxPZe4w+f1YYlwCEjqrxtGTHNtGk6+/r2BYSbDL
Co21UI00q1GOGHOiYajH8721ZPOUsqt/E3nc+vYDH6JhktQZY4gMP49wcesG7MaltQmcgudaZR1U
xjE6qdoF7q3LsOPPPQGZAOAMBsdJdARACH6Thoad1RxPWYm6gYSzapQc7P+aiDWHICZIlYSevMnd
3dFl86xj15i++DuGdD5AiTXIyDx+JUC/HMVgafiEiK7dV8lEpM9OwfWlonshjo2fpsDFVJczpyu5
EZwpKyJLKcSawmVPkFNgy6gdRTv0aOpm+7MBIbC10NUszeN9u3dZ3EkoshkIE/2VWp6lw57pI10r
HoatZTuERTZIsEo1+IUG+XJ1FUmjnsQ9qXSg4QnxXvRdvhSBuiNmjhrMByNtfQp+VQnB8TOaGqD2
MVGJ9pzbiawnSr/BdNOLdRkoK+XQTONnGEgdbcI/ZCIEiNOCNgE4VHRTpJlKksLov6Z4VRCoF5dK
W3GoFFfvQTJ9khj1E6JmHeGuCRxzhYa+8ITAeSJ1Csw6ZB4GSDDVBDo7FGcccBcgIGpxo/MtBs9f
9HjWyLXUQzXGbSeI7pBl6o5UWlEseyVTjHyMcoLQEI4HLhcsTI4CQKJwxq7xdZsXPDHE8Fa/5eey
GgZG05jT4dXbR735sBzJe/nBboSHggEvVCsl8bJh6vB+VU1gLPl3/jNE/n6InlAJMjSmCHDXMhLg
8dptCwqA9h78/fqa1xSYKvAcPSzS4auzteHDzmGbFMt/Kmf7Q5n1mNpVfvH+nLuAX1M+FU3dqU+s
KyCpqDhnRWdS6PzUIcVM4Vof8lXMUKiZjq4umZHjflz0eHeQTt7+tcWniyFrcKBTv1KzHQrgvl6+
Hy5KKwQXVNg+/xg3CJ1a1eyn927mECwNmuzJ9lT/6uHm9rlvlYg5kqWIBJOUqw88G33oWiCCZAHt
0/3kTQvcXHA6dGAPqtj582sxPAZNyOVQY8yCTAkd6yGkMtGLMJ/1EtJYr7XyXbtAAutRL0F+Bxvb
B6aG/ZnC6ePsEArmYG7XJXksnM76zSjlaQOhyaRuqdu0kKzufOIpk6qAM40Zergqm6hVSsaMQT3d
lwXQy/9D6ciONpcE5xQPf5Sg7lCJu+260m+KFsVCrPlOWsjDD/chy614LlGxxa61zClYE/x7iest
lGIJIMj3ulV7hKnFvAk1clcqaI6J4eJTUPgT32wH3qfTrPDM7y+eJFHwBC4O9JFbm4nEMGsFAmxw
h+KquF1cm9Dhq0sH17Pf+q3xq9wA2uKGZ2Pxfim0LnpsbnvltfXHNS77E+7s7xegUXRaFAdfa2jQ
/FqqfknYvItYE7VDP/Wdg/h7t1TImFGKBbeSFpi7WUMCTsv2ZyJNhX20vnlktfJrq7UqPR24PL0C
Ym8spIHT8DAP8+W1108rJEAXhjUhrxkbvtoblkxX4omH8pRD9gCm83UC6dx98i4S+gRX8SBkYh9I
BV/6WlLrNiXqcoLU7Fc0AfCqlYnrvOztYBx+SN3kE6MaaUrXbh06PlIclf3U3Pn3SlQVBUkyP9dd
7vUCO3sOPmqPBvKfmqB9wr9MdkS2QlekA2fTk7IqYCrm24fmoWY4HHWRPluHHgtngwe4U2wxzNK7
7Ui+0rzWszeG7SNoBK7soDI902FjLC9+QS7XR29LWpGp04a98VUK9W95ISrm4S5Qcce5JECZ0m7z
fA4NAge4PWwaTEA1vC8Piz8+QQpWqHg15XQH6M84frxK7kc+aSecofKFWCult+VJCUL6d5FKz9pZ
ly9nRnkbRnwBZmsYA/5yoRFLg0M+OraQwmoRI8og6K3lMmpNhBNyCmYxyV0BFlwwhSdUS+DUHVOK
hz2PHoaRGkvHtmOUHKq4UtPQbhEZmRMxatXJ0gd+3uYlkCRi8xLa55UrsRMPBleM/Cmqcv6gijFb
fn9s60Ekg6it5UH8Z160c0jqAdwJNdsOIkDjdxykAYX0EifLqoHmr4mu/1uuj+TCnfodNyuxEYOe
Xp4JWibo1xBHejTS8/Wj9w1k0TmDUDSyKYdUWGBOldifaXkv8nEJAo9dI4BSdSdYkbWP6GlNvQ6j
gjd1/SB6hXqguoGo+Pcj2NzyZE45uWsXXBKllNTbSP5saOyUk6c6TKgNV1y6NHzNfDoSFKh54+0z
J7Y+2OD6CVqo4+R/wi2UKjAvd+1FeUTYVLhuMgVRypsr1a+8HeEIys3rgauaYYVxET4EoCcKYE8n
Y891e6S96C/qO97oAQFt7gxgd3TtQfpOgz0Mk94OEkam1pe/5XZ5bNUbVsxSorQwLJY0BtwmbiDb
EEDgeZ/PG8s3wf7CCg0pKDGnuaafr3fhFO3b94empTdX8aFT48yYH91nXlAJ4zPhUime75YJaYec
9S84Q+8wobUY7J1jAfLvZQB2SUwJPDmMzS1Fc5piLRLpPAMo7YscrYyrIBv30WXHT+IttwIcrviJ
8IlV5YPut0pxqgp0ixfR+EoI5+N9B0EKGjLuIOsuyEZeDGoc9kyE2h39HC9fxzrY1aPltdJZYEAO
pcIuzUsKP0ICfB5GNCRe5NsEUz2k9J+L4LvcCRBIsS+UzWrzHKkJyuYEeKGVZzhkLaMi+lKnpFAZ
didoOT9BBUTo/S0I5q447QHTikigH1H+Zv/r7dlQNeJ4uDqIMIpq6GXPxRVITQH6Ff+VN21/mI8Q
R5oB7E+ERLGHkuZSn7FAQ7XzzhqyoXWFYgyHftFg6IrBxhpUGley+girGPMf5FzQlo9vQPYEajPj
Sm2JmaEDYzv0QbPSBcDcxQXf4EywgozEwkZV4YobBzEkkzhMV+oCcq8CdxPl7ZJOCp6CrUTCE8ht
RPoENTCwWaOeet5DqR2lRcACum4zG+MQKw8ZDD6oIHbTj7Lwv5uJDOYcqWDBbNj51lUFaxlKk5Rg
oCN15tXtTRNEmxFJnh7NZSOXPdCQmx9ypxh9SJHvYp9m0txRUPcKtynZ5jfGQ83SRkG12JObRpX8
364pX/b8qPyVU43IqcZt+KbNbA2/9QE1k98x96hgtTZ27HGlQNHFkLqoXWpWw8RZ01PbpzDdQIhb
iCGEVAqOKqUnsoSLZhrUluniM/waY/S8xNT2b4iw6+m6wNbf6IhIlwyh/fksjDmcQdwm1omjAiee
SpMQDn95KVohULLx8cm2yqZQDdo9Tsq+1RhELVkRRHdQhkntL7/T6/UxbmDUsCXWg/vjkn+j9AEa
iIhj3igDqp+bG4vfa+vfbrcq7KXkbt/wqqur0BjXB8jXt9mvyxzdOxCCT4xpPJwo0/HjZ2aEwdrb
AfD1lNv51w4FbwRA/+UvnqyxQXxzF61kmDElChC+EplC3J2DDObnNkCzo3l2UFY/kUdAS7dzmIJs
u7Dpl9c0HtrCHGAosZxpEebmC+XUPgK+X2szc/sitG1hoeXD1A9D6oFFQZ/0djaH8RVQrqh4Tt8+
O0vKCdFmnO4+qfIgCo1uknOiBLIvD0ugrGotk3JySqFTUrYo9cCK8i+b7Thv6rfTWRZ5Gt9iEp96
fe0YNX0vkEb+j2FM2S9as/615D2pl1OashGHvYZ62ZweqIvVqgO7K20Q4OO1hjXGGIo0eZz0Ec2J
5vrom3aCy7hkoScKv9PU2p0+o5vvcwQHI6qeXHb99mqgu7oMEbqYnLxbj3eK+efPavMuJtvvt+ve
lZq6Tuqn8AwcZ9/gvGp/bg9ToSTs79wG9UccW1pgsRH8QLyC0Y9V+OREthG1Ts25u1POm+F5PV7Q
Z27Ncj+uU+Ff3wFfnNqA7Y3YQKYFnYPT0bUEzd4PntHejeXcvFTZmSZo0OqXhhQLLKK66NbeER2V
70cCN8ywX+fE6ApE0HbLFr5l3WMbUmTrnMqy1xfQn5M0KQ0V4HFJEVw3aWxdElifIqsDl8EjW522
INjR5PSc0dXCtFeYemxLqtMbZJDG5ztv1bdXX4bajsUsuKRdkUAd8+L4JLVrSU/VCoJGVXFiPTCy
xym4dGrLn2OsWzgfhqdUtIw4830lZcYH0+9DRkHIKniJjZO/6s7B8eaWxdG7faXDk3Ma96jilq1I
4l37FADYTZULeGU2ardH6rDnLeQwIR5eESg0jzHaOOsRF/pom3ajUVtZeQ/wj9cf5+lFrOCDTz7B
6PSX66/IJoktnylKel8SrJaslqR/jNhbko68z58NRwSH9ViKi4b740XsgBHca9MjADZxD+752XPa
NljbgQzs8cT3/LACBu1S1x8+0/LtsKLZfWFzBVC19cPhbQ1nLY1YuFzSNnM7HQkueE7s1MYfFnjK
8Dqb1BA4ieqV662ozYcTLSRPMxKufT7drakmlDbROnd0L1eK3QEM3LgDd8zVfkbsUXmMNOIkNZrg
VSOE9cqxiCcUPyQdlUrD42LrMl8WNcc3Fubw0vTXzvu+vPkCaHvHJ6dqeU0SeYSlJfMgXa135XHx
KUKFwOcOO1Bv/Mmyk3cwN65fHudAlupj850286hS8SnevcfGXVQH/LEeWEIw/N1JNUwjAozpnMdL
tVE8ET24gMG/DwKbazzjOnUAvVE6fIk5SpJv5KxDoflIeZfIFbUno9UDKMfS66LTjHSJNSKzx6a9
b15Ckg7wuTQyf3SRD6gwEgGSLhp3xWg+WCPDCs0v+E5J9yx3iOl6Ih/vL0xAdJb+rKbg75PMzoNg
094M4e2R9wYWveKuapFUkIypyguR9QgzCozURVSwWLN7xfRLddls98eMa5YFlTkY8Kbre16dQp4I
Bb9job/3k9fCu3ONsUvTe5cwIN+/ifV5IxwYJOWWj+hYVfi8pnawGBNs8RoLKEltuV/vqqw0DXHc
iru7mN6fsvAhVQZdm1PeJ4l6iM6pvs07Nk1vzLN2nNXVWyeuXkIKxqmUhjrJzZfRA3K/Jf3GRln3
9zZiiJX6ECYrD+kZCAUPWMK34yLvbSQfV3VVink+JOStb/X/BDojaCbIz0oyZKHmLV/z40a4v8v7
BE63EISLn5XSMO0i/I2zX74ysPDw0BEazEs5yR9m67w/PvEXgCoxEbnQgiNX5x1Thy4Vp7Iaa8bL
yD4mBuR1YeBo10PrIKzawpsBGERTXS046eiAfv5KZNLYkoSL1UAnVqKkGl58/09F+bdUiZiOE2PG
J5Hpi/kA3b6jeAmFYz1hCEuGzF+KGQpWvwWmMZaXjAlJXKdjBDByD8X9DGP7vzNar02Jgueh3i3Z
myLqiLlvmwkScR+QqHrl2gePHPsGyKA5gb5UzpcNSwmDIaUelN5VgEPgXlS9AJxc+h/gN6ikMn8M
DfYBgkgaJGb32V5gKUnU8GJ0SZgz3MJaSiboKllBPW+Jveu88Zk9k/jFbuSwwU5IOeQX5V2FMBmZ
ury81QJBIthOpL29QZcsI8Nt5e69/e39khooASTQWDLAumJ7neldojlf/vHb0lptIMJ2Oe+D7ruA
xKjsTSZnp5GHUqSqX9pEGey8b7eHJxH7VNjjuqWE5WtbLMLwdz9aqbwtDkzBEFcV853nYRYDt+6m
Y+ck/4QNL0eQRjYOdFK8SNt64NRVzm6QEHO/5DIQDRVnt6skT3KCyCkC16MEJpnzE7kwWlGEq/uv
jhbxb2SRpDLDWHu1/p7+w8dZTDm1xuw+6iC4eqSLjk65I6oubIPugR3XLSZiUlXbIAwklGFSMtDK
LeLwyZyPDA7jxCr2nb/bJANL7c8bA1y7Hrpvc7BoIvq/FbZjprpkIxQLG1jyfcwHaSlts9xnVtxs
HCEhQ2rjTxdR6QtrDKvyPEHvOETzpt7IpaDNY62W2CbLqpth/WdIrpbTJaNa/lAphzUvf464+xHN
+NZaV7LHFbriWmZdsniVIyzQjcfEAEVyze1KHMitL5bwQBGxlzyOBGnsFFeZdcT2pfSLOpAjxPUj
HnGXxWnpmbQVHFa8JLm/FXxcBd5vMiHvdI9YlzSIKsn0/GSjHRF5xHE2qAriv+w9qR/8zQhxq8V4
SucAhU3CLJEUxF39vQhKlSVYPJh4pUPLFYeWOU3+PUDmv56OzQ3SVx7R6rRiGyXuFyrtMtpUV6tZ
4pwH5zCTD3u08Db2Jq6oqKoW2g1H8r1XRuiv3dQRsS4Wj9vHe6CTJPI9Sw+TSLdMsmfBskYt7hbB
LyrxrsKuMKrhx61rAur+a7acqJinliNczr1cTPbHZij3FtI11LhT3y2a4wMvlKW7PC9avaMmCTwR
HGSCdzOLOP5yQoSQdi3JErC1LNMr4VMGEumx1WdpXrRXm1NsFJGRv0l5eV5jJg4iKu7Z4XYttmT2
2unxcSVjks7g/3CsZAoZCUVVj9eScjoYwBcjAeQpE4uY9onaUUroNuKumkhfJu60vY+bpSyQwWI2
Gl0grfo87GhKE+xvjSe4J4chdhMpIzGQPf+AFXBa+KQwSnDTJz6x3mEmRGvVVat05ROxmEt3KPLU
saPGTLsNwwIV0LBPmNp2ft2W+hmAOwxvKtI92GC2tkZx8ltDDJ47lcrt6NST1RSc6ZKmdS9nYUxT
F1D4ltVXJb8gXOItuDXLlfwiPbn5n6xJgfehbax7X8poLDbyplcaAc3v5VtG4Fx/lG9eKDzntz0g
98PKR1ZzRgMGsWkeiqsqGaEaQ8OIbvyh7NZopCDVCYb+sKseAiP1CNsC9Y0aIxCATt2AFPUW2cD2
In4T4ty8uxeeFXnhpigZPyTBtG29wZCtY4e/FxTIcPIVCZEayMBOPNyqh5bHXPW5Y256ROxS1bS8
YSWzByc9GBypIhHQuDvmUCR5Re28QGd3aEFOFhGxNaQQA7BT2n/SFZqhkJdldg2RbU48lyTfKmMz
l7ZQI6A6P2yNpA20eKxK3zb12v5tooQD3rpSZVsegZMDcn02hLMVJFTIToAEWQdxVsRbPIYvOPmt
AM7sqboKXoMwbtOt6N/+lDmHSkdipTqL12uVxqMn5+I1i6RP58GyRGq0xqK1MFv5ZB2QDQr2a3go
eQ57ecYJhjhfkDFQNqNNbt08+CY85FjhSjRP7lpQsdLamVc3cFCnmbHZtTA2dkr085zEqi3jwiEi
jPWURJgxs0nyaCYvm4xgnsNbmSjl6FFnXPKtps1dwC5Zi6k76fmlpx+ZFgaOz8FLImnPW9KcA8UN
b/px+iJ5dOnDsXmZ11TRQodkrziVPDi+nKc2ZNBcGh9JzJ5Yj31B2YAs5iJa+ydeewxsTMHuBPtQ
2Li/P8yYSb6hn68loWsXDoUOP9ds8p9cTqHNNWU8kbN9yChOmo3hsB9hL9wATPsFmESNmZxFRDgz
ohIPmKJWSSRz514JSficbxF5LgNMm9CXKcgwg81kBSjHbyLh7875pyRVaYeIOXBgQqzXsHTcB/NG
jAJcikMa0yOA7WHPoJKcnnwwsS4sGkNY6NGUdUQSu3yQSha9gmCEhaf9/mfsRzMyrmhRUAgQQ7B/
28Ok1GZdf59K99mkKxzVt4MHG89+vv1MdiElo4iZL3uYGVP+LaJ1X07L1uTfXR8K4eum8s2C8iPG
QDB1AcaDf5PCNmXJoq9Xabt32+e1R6qUgmF91IVXRST4qEhBSvj5jHMG4DswM0whnX982eqOTLlE
XqbRodsw2x4bJB+wx3CqkFpY71KukG5miU9qdEnw4E8UtXVT8rGDSvO/cK5vwlu3B9eZ2f+Jgg6f
uFtKyWIpvn/z0pxRroolqfZ/cCvbcWXXLlNaiei0PSPyBs/k8Yd6s2zqQuju8HoiEv2m71+ysYEp
UOjGo/VbgK+vdAgLgOavBCjupYYKVcFTO60HXcPrIjd0RQDxNcVvZ2beVFnaSVSZcKB2Yv1yjs3O
evpmEDINryIhxtOKw97yW744wrwWl8J8jPZpo5m7F1HgidLzOVj4TuRdUp8GcoQuc91aVGyVATlt
hqKbB96UU91gvcJUqZ0z+scEyNc3HPOcvYQiHzpChkhvl5WP3ep1/O9fdPU7UFUWvqLsZR64ylYX
OngUwvDNfGWy9RzZYygwlzNQKo/OYZK3UL3qVAJwKrEO1Ufnq0Tt+pwY9RyUDX5yQMEBCB3UWsGv
jEPAaUY52UuYWIg+uE/ND2NIzcRv0W15yBdryZRs7aLazuVm9ZrUJbxGIR4v5NOyhG+LXP1ppx+N
j1KoiVWip5BTxbPVCnMfqYA70/6E2dPTRQTa41tPf2oSNqcd6XWC3jy7EqyTCeXacgc68mGIZK15
ma2/FvQFFFlOG57J3Bt+WXP8P1nFupHEoJr7Jx1rnAOKeMHWU+ty82vN30Aq6efOyHBe/OC92K0g
U2a0iF0OQ/pvjlHbOb2zbMPu8l5lq7Oez/nEgjh4o2nCbFxraBwz3Z/4YTzt9iIBKUUCYioaZhEG
XmgNRnl5jUIQ6d/SqSW2vgMjI/EqiH/Hj43FSQ6FVL0AHo4q70dlAytQ/SwpdDdYKp9s0wnx/FPg
1JY6jcxdynDgpkcXjUiLKNi23B8ilmxN6otKUDAwwvC7ClOxUI9AfTSw0eejmkHGVgsyQUsbXCRj
DK/kSIMpo4cdia3hoSPRFv9GnMs5KioyDTNuI7ZWY8HIAlXxMbHd5J5jzxDCvxmcsiTLSSdxGvha
O3RmjKHhuOe5odko5GkZS0ynff1kFPNsmjEp5rcvKMKmhqVsljRWp50tKbaWXBzsXzA9fgHflvSH
Ttt6H8jhu44Qrq5CCYbGKaAnlHpf/EkwN0J9GADx+4Ncz5Nb8GeXRKadI38Y+YKaD5RQlizyXH0f
R7mneqJha02+P6xrwGC3xNZp+g76esTnQ7hLmxvY7ZTejVAsdwJs/V6YJeRbPGL019DSVqd0wu9U
b2/uEt3a+Gncvsa9oTY9pocFVEP53eleqfsUu3gKCVWh/eYBfd+KqhiEsCk4WOq3uWpnPDoUD7Bd
/Dls0SB4vs0xEFComZJVLDbmotzbHfYyi/jBlFN0v9Pu5eVwrP4LrxlP8yKW+AUjWQFrhjkVhtpg
RrHxLKinjxB/rpCkcO2Ovh/VhuxN4b9UDhcfpU4esLfBysBd6eqOPKGoDSJJBj126O5384xZ9WL4
SzpmlJFCujdeEk+Nb4mRKMB2g8PogsbNRFFighslitmF+Z2wQw7n40LF7CaEDbmyQ3l2R+YArnGs
P3plRlQ7d7QM4uB3jRbqlRE+infO1v9h2g1GQ7oKCiOJUV8VWrY6K5UvoLJblC1EUSOlqGdb7FWr
7f54mbrJ/P9ciqc7Q3mP8GiIie8AVpbV9lRXeTvI/QwvBOq3G/76wJcarlW1c6MRKrPFc1TRiRUp
5JLNXvYRNO6ETpmDt4RjO+xvqBGnbe7O581dVW9mjmXRa1yZ8DDmZNOrDL0DFDozisW1lYp2V7dY
hAbyErj7A0UDiAGIpYEJH3oAgYdM4Sa2XZ4QM173UbyQS5JNrOTeSGyOb0IeprE1S/94grek/104
73oLcp7trupkJnDbw0qZ4ATcdaTp/CkfzWLvFlCAn2ATY9xhtYBbHWMJjfznF30y0GMaX2ryJ8ok
PPEUgYCqYv/Ejnh1RQFtfvGDikAKakQRhA31mQ3nRI3+qJ5MlwkZU3qbg7Y4F2viR/mvwfk7Z2VG
UFfawpaI6EDpxOK/kf2kjpQPicaZMRzDVuRYMbOJWbpQHzphg+ibbpc+P4VD6MSFqh776UhDTX+6
1xlDC/qn3vZEGLyX2Mswr58fA/OanPNXyGvAxAoyhxPdnO17nbwv4HmETtsVzssyBBTYoMts2FJK
Pdf8SWXxIc9NRcnTHFRUx6iobmJ9eX5TdW+k4OHwGKdZkTXkrexwA93+taq3Yif7PArPtXBomw3i
RnduY8OMPO7MX4cDsxmaTG2Zhn1sia5fUXWJ40Xg87nmMFnFi0JQDDQLeIhHqLPtfv+qt0pw5LFK
VME0+ZIME/87F1u55l0CawwNLVUcJTK/9+JQolcYLFSOcNXW4Elp8AvwGvpU960xVk5BQ8sCjfgk
C9ucEdgki/R65+x8vowrTiZnOuzmgfR9gkVwnNAtZFn2ekkd+fcS2jSN1IArUgmXMApDJ8aAYCqq
jJn6h0vOeTV3VlovKWRyTyKMzl4hS6GJ0QzrEvbKlIk54EznuM+R3I+g1so6P0LgZHcfRDxtiYab
G3L6dLYopNi5BPnmd8Jj+OqFXPkz8MrOdsvzXUXihcTzgP94I6vM1T8sYLoGjNIVfnb9pl74CXWj
28mupfCYdWw04Nxn6Gu5JC+D4orTNUBqlYEF2Fo3yFI52hSdP3jYXNTcroORZqn82BMnqRcmZy71
HAe2in2GohMP6E/+16cYvto/IPZ8PtzIZ8RzT9CS8N8lYrbs1eR5kkNKThDPzfB43jjZ9DThLa/O
AvlPEWij2oIkkAWl7186LDYjL8cJk+qyPfTf0KJJlTXfR4xkwkHYrRETlw/joHLcvR7L34YKJ6nH
vzd6j09fivdQSc87tHdX4kJsw1vuM0yVLC1j5Cr9o4WO05AKKuYRTW3OUMZOnwWMktqS0Rt6B91g
gdclDCjm6kIXOoA2aEGak8RaIv7t8zTtOlrua8DStTvQMSEQQjO0oZ7xo3QilSpoEsj39y/2GnXs
tb4IL+0lh1JeTP2bpgZUHVfRC/5JKRRmBhEJLxWM3tlY9sstbFA8NpkGWxZ345ayOBukCJzFMgaf
Ff/xecvCN+CIs/E0Supd0ELgYuaBOnkzeuxwuDdG00NHwdwXnOQHO912CaNbP7bpoU857ltBDqe9
gIVP1x6Rk+fT6hgCjJa5dafcRw7uiTnoGY28gnvH+sNg3RV6navEtjkgnvXj5LZVlinuSTZ5wYsy
1aT9dfrks8TUtVIWgxTN6jDLsB6Ds2BuPz8MJNG0GsNJu2gC5tAq9W7RwIm+PdDEF+S82ZsFM/60
dwU1RIkVomyNLwL29tRafuXUL8IUYY+Y1yZyJ4Epl3iNxm0knzOPE9new2ybnIYqB5p1RKcD+goh
aX8Vytb7F2S3BOOEwQFfQD26Pb8NEOVXwZcS+EXn4G0SvyaTFXOUOBaaP55WlFEUmsSuqURP/xd2
bo9wH1DyQhVawZUxgskBtpts23uwvR61UyAXYySNeThbAHGJ83w6rqYKnz5Yy6csBR0Ps/SLN8Db
JenSRjJ9Ym3N8DisvyA6QvVQTpRL7eEqTqNLN7QRmYEt06DHkxNZSkDaKRvYFdSyrwiINcL1JG2M
5Os4BtIJSI6tOLnFDdylAUN9jENdYiACof/DhOMvQmJVXqj1qvmzX1tZkKZ2d6/EgQUMBEGnAx4x
jpFIX+9mOdRWvT8AFcOmv1lg0UlrZAocyEYq8Oq2pgpNez5VF8LaCVw4HUKftKejW2sbnqROkiau
jcTB4ANeuiuBUu0cKLsCo744nuizElSbaCsHeMIQZbj8c9AiZrl61WMuAczHznyKfHkn+Z26Oy0u
U5PuSfLbHJBpT8aG6zV3XOAAUFB87zYe+sx/kIBFFLCx0eVULVM6odn9GTlm0AMvaA1MBmaIyiJj
Pc1qCDbMjloDmSPUXMDsKCD8vROErMsCD+Sa4EmdU3GmfxxlUNr4UkFoo4XGnMl38FJP/CDyivEv
sk5Blf3HiRl/5AHeBGstXnpnnSWfzkHbn+Aq02w/v09qCnoYCxiSwfL5Z4DkcYV+64HGNReiGuuJ
Hb422dapr1JYgbDuY2cgCeDTK/w8DFnsPrqXrnsHPB+vD1tHUO3bq2pjlKb2q2ngRT5wTftLV++E
AV2v+jno7Bph9WBcpscDUIS7qvNrfeyZay3WdXBmwyO5GlUpzULrwiCOOSa9qBNw/zL8oUyvejak
AnQPflj0s6syXbcwGL/o3Ex5VHo4mluo9uVcdedbrVkYV6duwdYf9Fy7rDd2KVOFNBOJh2RWKiOj
RX1HCDnfqyWzVKxxKRpxmmS9W0fHJsJ8/vyez3s1XlsRJXN3l8OSQCwo5H+yr4GWW7Mae/zG+iQg
pjBW5BlacO9qOhz3jrgYWEzN1/7g/dqkjMkmNkZHJNJqFFLWZxZg4LwCKu3JbwqZuHat65GYXxM7
9RrJltA78bVPfjkyO7/DSscI4SjL3p5gjP3zBWZYPo6wxZ/81Y3ClCblZZRYdbr/MFx2ADq1srLs
vVPjiYB8DZbQojrv8IHXWajG0R0bGWLfWyVCjRs0wIs9zMEx5+xhtvYHiokf+hb+Ai/L1yb74JY6
EADtMYtWG4A54y+aUGU/OePOkRVEXROrZZn5Ehn1bcEGdTJtW5+BE7PmWJCeW3IMxz/zKzzrdhHt
d8Op4c/qbExcrRVgg6/Ood+SeTTyuIEBy+fxpYJ7/IM404Ncku8qyox0nrg33hPj+O1V0aB2jIa0
ilSwVhXGGfptP166kFioL0XTT7CJNbAb3D5lfVTbk3QC/Kok+CSYCM1gXUZz3zObfS/5/A4iOiXA
w0kqJWuD4l61C0BfCwMiIccIBZsglo0R3aA0zW6J9uGk/jFGMQXTBQybfD/qrdUmxmKyqpM5/eI+
5i/Ei688E+s3IjZXyHS5MqieSLAu6yT88/d8HyRzASihLmnOj25Afq6Ha69ao6sKFOlrFaix4CaW
K8ZVUhj4MMDENisjtFEdHoFtr2YSP8+i6Hn2y9d80NrBjsztzrK/t8Mz6mKBdxFw9LsKs/ouFYBa
anmp1qJ4jkbyDapNjV6Idnfj2UjTuu2V10a+Uk6K7FmZF0252r3Noxi4uny9Rai5cmJ5hF/r0El3
kIL5W5jFiowWt7nTVFi5zYI4lIxgbAJFnpTXWyL5kasV7ikNq8V8bAoGVXWybdvR16GdxPBEC3Pa
i8Ya2gusa3nxAtzNyzFFT3xPNYoKlWMxBWuSENzi7jOIv4TT9qo9rQngFFaFYs9J7zSTe8QFdXkT
ykaJAAU8Ct3MR5udxWxm/sgfgRe/miLj0MW13ylvw/h1xHE7IE7MfafF2sFao363gMYt8SLxuvh4
7aQmjcNQes3f3CxWG2bd77+ma0G3n+xl+r8dxmbRi0hVFTMGM+xK8zad7piuR59b2dSbTBfx0vNj
oAqfVL3lfCcDcunj/5qnWgdwiZ+Qp33PDClDdALcqL/xCHBcfkjaXuJM2WRRUbFUtgGjPrf8KiCl
5jgGJ+oghqFeFOCNCcj5cdyu+yXfMn61gyZES3hcKOtJgCP61EeOkRPsbgiifOugOOfu+tTl2xWH
8sa6zORO8Kjra/rILS4/mSvTBMqGywAbdPMp35mSyT7leyXLWN6jcBrt0USLq+ui2v4/VlUmEp7j
s39rrYO1li/CG3f7JfPDEq2bKUUMx93OnyRpfJe6KH1R9T5FysV8NfbgmdWP7Y9G8SNIHkThNiXd
LEkHXPZVLKnsjbrHjMHG5LSuvvezvuqr85WY72apMRdgGPtNNygkKHI6ELoPhZTsqPfm4gzhDrN+
p5mjuCShM9qnJWkiGrKalUxX0Q18fynW4xPkDNUPIrNkSSjwhY1mEIeg7vQC8wy5uz0Z38voShtl
EtoX9dt25TBJ1dd6gw9pud+jaLCvdoY9vyYletufLbCBo1uFgMIiTU3sqh09KA/XyTTeuBDNjB37
Kws8dmXUxxwd2q5ij8ZTp4QNQS31sLhbQBUP4299yvlqxnfjgeNJHZ3OeUaJ6oTkmufVTNEq6asT
SgHIxeYhromJaF6hyTb/zFATXFN1m/vDnaY3vO20UHFkt+nSMnM1H8yQsm9izyVFFz6A9mllZZHL
4yuyf5vc9wodleiX7YLj5l/pePTGO32E1w1fn7JIBOEziwO9RaYDcoLv2Dxup63A7iSQb3loqu8x
Jt9o7JOfZuy8dKqZysYSP24ecFmrrfl5QDKuXRhRCKrlskzfEi4k2sMu12Foxx4szpWlzQRECo8a
FzOBj4ssaqoz10ontRQh4n9T+/Lu5hxgAs1GeBMLNC+lfTDngTaCpLRLMkh47yH8aZF6PCmHjrbX
CG6F8RvVOuyVH/FpZiYsWJhIQDj4qjLHBGdqLMN8n7tmFkNIrlJySI7e75+O+j2oXRSwEEC9jVlz
F+ABXHcEiig6R+4T9R3MsvUT9FXknw1l4GmBQjFKvk3Lms29bIH3rjETqkZ5g1dYU1yKnxgfInCE
WwdihV1xMDOnleY3R27xC2eNqWVpIqhu8ZDkfX3MQGvBahkqj8eUP6F4V6Fy2zRtZmag112A7ogM
VySLwCkegdbTj2bJEixRz4RbvIJHJlJM2bk7t/KktLstQvoB482e8rHr/VDm8lLYd1It3dl2FynO
G83N3ROaLUExNwvLT3/vv/hZF0Tsx9acySsrbghDgy6HTaQ7g2WJdP3Rz00PV8KwK9X+f+cCjYEO
lJ8K0cLMIc17fbXmB+sUJZg9An3uyIS0XnqrEcJSEeSAcDfaBvmsiYVDxip0krTDUol2qp+GACHH
OgDGHmvZHu3dmJjfwTNZk8jMQ1pb/1m8P11J5DoxMBWNE6Fuv8jckdM94f207BdJSL0gLD7EPog4
XLrdTnjbFCnjWLVfEMdE+gxACniKDKTpX4i6zdlMDljUJbotXj7w4RXhB9t0nrJccUSdqBB7pwui
W7rputeSNx4d++MNcylXcgexw/fQpdaPQEwIzL/rduCS6C1Qh2HhcOK6ijf9tRfpjuYlL4Eohjlk
wzRtoA5BVsWUe+aL6YvRQjPOVL/T4OeeN2x3T7J0KJ9aE+x7OLvpjmXUG2Qblnmv+xS3+VlLQDE7
nx3a2hLIfEUv+1g1oKSvUaRtZgCVt7uF2wZZCzAZHtaXXzxNPU8axQxHzJ2AG/U0a+9j71oF7/Ve
Su0DP+2bqml9AHi5vv2CwolT4SV5JM7iEL6djL6bHf4riqYQwPHAK7uhIPVZgO3uEPOemcZMWVG1
bRdwZnyF5TvxyV1MFCwvxGg36TpBYLRmgzlagpexLEuUJbEMsuDb/iWIRDljWOD5AiQmJp9JOKC7
yCyJUKz0jhMjVE5bRqcpwEed8wJPbxidkuzVvMnwxYdGmxeo8VnhPevwVlqONkzu4JgmWycx5ztN
pQAPoK2BrHgYva93q6Mb5HfnwuZc/0QCG2ROAtYQRQ6ytFMceytK0eIf/6PxeapnI9Wa07GjjfYZ
s4YWw/m0rh9Th/yTc/VLsQcx9U6QGRr3/oAOzmM6/cN+qslNzZ7T/nli48XfxR5Jcy86Mz6Vsph5
0Vws5RjZUSoHryfNEWd1SvceBxPCTANs9QMeE2sSJRWDBthv0lhjbG45fznvcWxJ9sO36EVTuR4C
GRykxSQtj7jlV5jDoGNc+oL8Mwv22Ti/n14yeVeBAmxcz7HYykTju8g/LllI3mZP8GEFm04YKblq
8isKFZUAEGCNJopx5sZyCn+FubkeNM2ug7NVm1xvcPlRuMg3eMVkFhpBh+gRvXHEc1zleFyr1/11
dTleqItoh+VKqkcKBu95n2RN9clKcuifMWvDE9cdoTR/GltUK2J3Od2CY1GJJ98X7aU65R4Xj4sq
IyaupfsdLUNMa+D40Qpg8ChsWTpFUZ0k3X0oh8I12qtQK20+nShPGakE3/KqNtpr1Ugnoy4YqAa9
3zOUctm30D+C1gPgSgkyjw/W9kPboaFogjLUqgm4yXufNqBKJPBBZ/cewyLqCI6rKkzJysJerjro
Ae5yRqe19P7Ei3jDcHLovKocHoJigG4t2SKB7KRfsaQgVuhPNJ+jhsr5hzoIhfIDpnM7N6W0Mins
mTPVN2d4FheTNPSeyPthtJbNsTdWo1GYX3RQYqwg0fNw7inrzs2SX4HR/7WQ7TUV844K1q5IUvaD
+8D3GrmBm9IB8SSKlIAA2OVGdXxuLWd8PfvgDJYOl0+YlAqpu1uBaaabWm4VXij8+iTVZAYiBfuC
aKRS3HZgg23DasB2SjNmURTRBNnJmwKfvaiQC5A8mb+GxYfGh9BZ74dnp4ATp3/SVDcVPlr/P1tM
LNYbly7FzF/ybWUOFdr4QulDBYJNBMBOCQ6dnggw9tYTPGsaFfHLROqoCW9eGPAWij7H9e+Atsys
10X8aBp+GtxTZKkkNoz+RRC7p/GLSSTLyk7Yz4NUNBeQJKeO0x7iQRbdByCZGOMqyS6vYbCBUd1Y
JyKT6t8ZuGzruSWCuoXgooX9Z7X8mQkJMeYnIU98iHNhOOQt+4yw0/zL5Z0G7FBGX9v6/17IUc8M
kcC54+hnuBZgNYAAcJZzQCQe2fKCjwoxjJOKJeQl6rmdkHU/IqZaOD5snD71rqHdrXwCNk1Z9NFH
jvZVFdFwAj3ayohWHZ0gkhckwcFWmujGKM0cpINxBZ91LUPiMh+B1tv6S8cDv9iawQeLwNMzfOcR
etTHn3A4Y53tcYS943zndDvDM9PFylfy3X+ib08kTSls1umVQ9vl9MQf/kanRNTxjo5EoiEBsKtN
Ct1Ui0ZqASn5IXyVgVkwbdrdKugNuT1hNRZA4b/P0nEBPWMEsDlMNeFLo5td1Yibd4e380nTK8jd
OCKoVWuZVxnTHsCl5rlaffRsymX5Qw5oyEKSSdEYUVCyJH0k2j24g9CtRJRHKuMP/l37hA4SUi50
zI91Apn1+ti0HE4hV3hCTmp91hhj9DVSqga3dJK98fzA/RL45LfHIX7EyTaIsMhcVAvkN8UcDnZN
caAwH7Zy5t6+ugzWbWraPphgHpuv37igitkUZP+QDEX0P57mBfSm2Ud9gJc2RWMV8hv8i6uZLVCd
NOsmtI8/Cxt4gpDUQUF8sIAI784UREhgivUfNxmSfzh5gU/hMNpr32OACwyYyhDKesFpzu7OJtHF
23WkLv6kgWNIojyQBJnaw23Wo2RlUsCq4okSGBY8DP6K9PpVG5J4i1uP4Dl2J+KItRrriS0ngr/z
ilPBJ+Z5INijWGB+LlXrcJO5mGXhRaMO2EpI+UXUPAD+Zm5yez3WeY06QE+zGgKKrKfOxGayjoFb
EmoQh5JCRaziCPXwQob67y0GXVlouB2yR2czzUkUUMZyaag/JECz/7M+wSVDCuTsEObXvGoMmqvh
BaohQqJzGWXbl9oe8j+8lpbw6/8KutNUksEZdxeeB72ut8BhVR5y3xb4tPcx19F2A9GxVYpkVaXl
ktNci26pZ5h3AA/TQZgzUSSz3TSUWgZmhBYUUtdQgaLSwCVc+LbBX6IsRNmQKJo2n9Uz6O71m8Oo
27fvymVY07ColYotqF4fd33+3e6VdLgii2XqwbcAkwhIVmbpddOTupIUSoqnjJ1UjPRbTULsfeoF
O6CcCVqbdodpiGmOqrtLqe3EQ4XRHaH3Sf4NcaS6iXeq+SWX9maxAMwSHx0WE9JanUBS2gvaQMzS
7ozY0VeLHsg8Q3lnWuKpJDPeNffKTuLTrlIlwglj9clNMkFmpZ9sTW1vu2R4ta84j1dpEo3YiJLs
yG/7KW6+7wlv7hwiMoU/u14iXzUajSkQYqOUHQxGO5hH0h76oenuZo+i+ftXsrvG4PHAmT/i9PO0
n14n10Fj+QpK68kb5WRcZQNTvRv/IWMtx4Em6qUMPLFkxD1JQEOtLzCio9OfV1SmMJK0ipdLv/x9
ffP0saxgGsah/b4AxYjSNC9tKIjXIeIX51wjq+U66Mpe2eeLsyl8vvdXFpDekt9BasTxsqsoD7pg
pT7h/Rg0dJXXv04fQzpnYsqyTxfgoXY627EYWGGU/lbda/2ypFwr+N+EVFL/IPOttXV/xQNR+Qci
cHGEcYga/ezutIzAYdOCWdqiq+aQoFDnpjlSYRCrtGAwckEnfVHRgOIIwJ175BlemPVGA69S5jFq
AaZPvMFlYuHs6M9gpyMp0GcSh8o++Nsx/gchwZ8jgZGy35+JESMJhBZCb+gxveWGFmNAk8r2S6k1
QOtES6K617FxCk9QhMS0bzw8R/p83eNSpxUalkwXDkAWuX7tlcMw7951Itcb5x5T46NsTawsBntJ
NiV8TQFkM3V37E9jdHFDPkF7N8wesPuU9hLfjH7Fro8v/2jscgQ4K8IZ9f5Y2VA3DEYFSa00T7Bc
4Mt3AZ1bQfbG5yaFnosO1nymZD0+wX9K87Sgxg1NodvGsOZRPWh22oWZWUlLn2hQqgHtLNuACN2i
CJUn4tIfPPe0cVUw3RT1pFJMQ2cNKNfT7YUmuytLBdkFFzEdhlSqhRDIh0SJCqG7A2s4GxvU7Rpk
CtH6iJ/0EaIbgqnMSFR7dxE/vMaRLNqBrDQItIM0+WxhjMZr/i/pVTO2RmwaJpYrXRVJ4dSd8n8K
IeYZaF2hOTKY5C6IS/VgkktfpO75f5QDRwCnYlZ9mU25MoMPhxgcQ9XTkrEgrn/glxSid0o8y8+V
Z87V8ZKfXACw1C5jzoZhgs2lYhdmWdObXkrG+H0O6tanmhvvn8GEc6korwXnveyXadgtEBzfhkUD
c4kCFh+i2PL3/kzZlyw73SqODkRaePrOwjJN4ERbPV78Qm2Nw0ahAUZIk6tqxk7VxULBW0qcsA72
INv8h23MMttsj+LFVLP8tuO4hU03MbbTS2nqaUskNEN4hWbCeHER0dPCyapPPvAnlhBFX/IpKHUS
SzAEbzZ1g+u/wZHRlNjkWUbv30mY024DODzCIn5tr4p0FXIuyRlSEn/YfjAd3iboBaJOUEuvttiQ
hLQ+udTmTVpuLT1FmNbnbJ05/JYYFC1qOM87Xpe8JPeN3j8tgqaj9jBu3uNu0JBGaFjVH3XmU0zZ
Wyuxm4NMp8EJoKVDgvUbOWbsAXOiTE7G0q+A5pq+SxTJmpOaeQARHkXR7P4k7gPDLMdq+6yQuyCI
+cwoaeNydpFLLdc+Bq4rgkchRcl45BpbPANcJroKoZTJk3p9IA0zaD0H7WgiAsyyXjDBuZnvrmxm
kmjx5sc4oijyAy6XoDvDchFUwMgysg8kP9HOVZa4ru934QtUJAq2c3Hywk1iUYwJY3/FfeGZu8pc
dhaBnagUvHm84NkSzA+xI9wnAAdUT0sKPTjbnlFH6LSCboxwBy/0dWowPjjMek7RcbEN8C+wA7yG
X/C///Iy6N1QHwUoaAorLCil7Av244lwwwbvE2DkjY6XdpvtB2uQRI2pbyPAyWejVLwwpZvOIlSg
McGD9BUihsvVs8vAo/pzchIihcy4DX7xxKePNgFxFd3YJmE+XPfVVn0ICEBSdk02d8a8FY9kP7Ay
uoG45Q1ymF71dOWbvsRs6ezvN9kP3Nggu9w6r8dyaqEq6wSR5gvQ+a3sYjgKUamzgNh5wNmxPuF4
42L6BR5KXSGMaT2nq7MP+enYbAg6irxCW9D6mePDAgMeKbLqtzoyeDf3/kkz5+XaAUsRxaREJ10f
R+YX9XBzl0ZDB/Jw3hA5B/pxHgdtr7CX0RASQpWhVCBGfooN4wH2CEXchCIcLWCj6tBbyAiJU3T7
92M+RS33yu+BPbkLEasgsl09OhfXCjYUw2rRT/UodNWIm5B+B6tODdW5Mam0vGxjLALxT+ToebYV
KCDKzoXQyvOz1i9FbZgto1x79FUccFhy4ARi0YWsmJUuDUKh9kGZKrDb6i4rr+u95m6fdZoVbE9d
w59DiEAgIWn8ZSNUb7qSeeBtlJCMJFiHZFspy8UDMQp5bjYdvQ0/s9JLFsNuBDEmjFsr+uY8rior
f3Mu2TpvX4nc07hF9oUFSR+SqlKKOkyRQIM+zFJcn3zmgBRzuxWveMhyAsDXvBOon0+lrIfwheHz
V0fzPnLBiMNWaQtCJpMzqq78fRh6HwTluZepxju1TPipYTZEQ+kl9dgFYt9KSVb8Z1pZ8AMARzVl
QBQ4OUR2wCOIKHKcmtOB1QWo27YsNO0vNA6mr8HNTNGU98dgY0cEhSks0iQFD3j9T5mIbtWirq/C
umAQokU1RyDlrgqtVcXpGHQxwc4qG5Vhdf4vgmYN55RHQ/LXMEnQMM2hXLXEeB8CJSjFkF4ea+qu
ujJU/nnoCxKjDvICpEDQV0UWRi4lna1M7+x5fDfYx5ymI9p4Cboj4ma8WO5DvjKaHf3mOTrgCyTy
zTCR47NFkFwstMsDv0D+raVdMg2IYbTxsocNxC2EhXdmPcWOGIO4tk/JtX4QPTjeF0WC11E1Qfxi
mgApSkdg4OkWgZvW3RxKT2csdwVnE6+pHOWZ4Ylr+nQUTTN+rTQ7v/gob/hJmU4DOxnYieJRvWNw
PNUhn4SndrZzkVCz9ECYG89rT2CMOdaLN8b9sG5CEuIozLKXBD1gjZ9TMCA3fke8diVislmhJo+z
2nrLcu2kvljE3TTK+FtKlgJOfB1XJBHpjFlRkpe8YBb2fbTfdS4eW8petJF78y++qLC08XRXzwMH
oyrArzGseGrORJTF0/TPDxk1xQpIb+JM/KVR0KKgcw3I2wlEV3zlb3baeGtpl0Uutz0zDDowQbZj
dYT6Rb3KLOnqbXygNw+P1oZFakPWym6HwcfM2BG44ouaguyraeJDYntAFyMSyPPOdcHCFIVFfr8s
NMfFzuyWSM7q1r6gpgk5Z4eLsms9Xg1NrjwHAVC7RH0lBqDdwvASeKEnk37G1RmdgvSCEkdqxjon
jJTqKvxFnppKE5qJ0R+3f2d7y4tRzmIJQQqYckMyRfWrMDl1yZgWURbxzTxbz082o73CRH0fYve4
x5K7Aw0YVI4UdYskkFPBezyrAWr4nJ4tdn4DOzZSwILbf1kqowK/r4QX0p4R6wrrSm3HCaCaLL4N
lGIIIzh4ZebQD0cBm/IN6vP96C6Xqv2WAr3VLw2gTfvkl4ePZztHUPEhMz0nEDMApDgeM4bbzJ7W
+NLHhQ2OwWeSl3SSv2ds60CgUD3L9BzbQQ0v5K8tixH7/ZCEg7SAUgz8iqcy2Gr3Hj1WjlIgO9FF
oCDVnV+YYoCfzN24cGi+OirhlqtXwwjC7SMpiYW47MrDaqpXNzBa9ZK1xfacZ3+DiHSyOgZI7XqK
wbnCardH1SSlhRAsLJ6E/xxtVGrsYyvgZdrfopVNd8336eqaHoqT58AAQspSWWsSwJLGwJR0xaRW
pswKBmHaj0SnO37plVdFpXgHSThKlILPCOfh3Dgi7BkbTxo9PcaO2ET3rPE2UvpcLh+yKL63G6iB
AVpS1Ti0rTXO/UnhxP7sZ/f0FKfAsSwZb2/t5YiWN/UpPMAE/8nocAsykpch/GN4VCg56MU2sRZY
BWmRzgR4s4AAPEc8/0WIUhUL0qcgWI9Y0nMFB4xhIXByVO9g3ZUnj9K3iEG104VkgYcNsFZExTNn
rP5lY/sIt7Fy5msV5Qpw8hSSZAkK1nf4YILlYdG2jdJatCzTh2GMyXFwlbHH4AXNglFpgUXMDDdC
fzpSzLkZaQGnt7Gup13Uu6Ld7dR6jtgs8M7Nomvl776kjmQ/YTYCOoGKF5nXoAaHxRqAuOd1/rk/
lDYfm/noHRs8mvKRcDijLTyOZCaszEEy/Y9txx/oJDnmq2McdLCdrkj41fwSJAh+ptf5r8qY0/vP
IWV+r6j6jZyimlkHAswZhLDOLaB47/UIJnaycWMotLhM83tWAC8hsQkN25oadez8WGA7gob7WH0D
bjAKJJMNwJoC5QNJrGy9cLIseGTpIPoGnL0ngyz39VPbnlVlE9iiEoRZ4j2hH/EapLWdG+FVLfhX
4rXLFZ6XWzy9p7iXRk/sjFkPBR91N5PSxBIRvAr0WQolQcniN8tdhbvEKh6WAsR8DtN2solTURGc
OJ9fJoqBAWWHK0OMMsZ9NQQHKom1fqfhKbGeZGDTvewTdjMN1owRehZbBXuff7w4kNaKiiAy9qzX
R59cOu65068iI6AuIekYJdbHJcc7jq6ZfiUQ9JmhI/MvYa88GDQ89w4gWCeTMpLIXpJb+fIoG6Ex
DOPjFtRj/YotY8qjoNUCGYxeQFvJxX4vXXebWtdoBRItQPuoXFEyyqZxclOD1U5fqgPegwfCM9BB
Zu3vEt3gUwcnVpdsXFCUy/rvnZaYLJs+ERfbimrTNlke1UIOrFkaA55Fpzm4gWNfyHGkhKZqjBuV
7HcQNVceo71/iLHYqNnim+hMemG2a+Ni0LKzwSGiArJ+S9BFlgBnMCnudRqeEiKMKIhke9uEAhU8
Tv+eGp3lmc6OgkOYXtb0MQFnrYfp4zkvXqpTjD8Jxlop+QPRfBeSm9LAFLzt+jL8m4saerv77akE
sA5Y5b8QkbuVIFxOFRnRvcD4E6XMBIZVxAVRJG36w6tQ61pbxvkHD+LoWP6U31WVV0zxDO34TjUX
IcUpSo6Y2a1SYD4AlkpR/gepCu6al6HCuHh063psoWNpvRPjYk9xkGs2uNkg3EgGKkjqs+4wW475
AeXKIV9nda265u6z0vdJrHvfOUnq47TrOJFTRKnEtxyRWn1mRGH63KxAy2IXRbY+i05mSKe6DwJJ
fJmZYEMM/fQgutkriIQLytM70Sb27fOvcarq7FFwII7GyFF6990rh4gVspJncrr0+LoGNBzAVIKK
l8Ve7pypn8AjYmf9e7OPaccr1vzsgBys6BERFedkLpEKWMPVBRNmhiKGpN7Ridx/q9miq8wsFT72
58Ii6Q5/SYVf6rrcHjil6ybbV9B2WPF/Sx9/X/O2Gm3gEl39O0E71bKA6ubyrsf98rYixa3njY1G
TlO+ZVx1gN1+Km5PJxN+zGjwvZvAd8+qFrz6JshCOikYdprd9g+EPaUvEJG9yd5pCYB9zOQ2y1Eh
uoMt7O7YF447Z/AQVX0a7LqnYDNE6CUv36B+ffbSx87PcVcA+P0oeJIEFW3ZTRM7H+sXcARI4BqI
vVeROQ9Lf/73zrKvGJVbzza4fJ4i4m0WWweYXaEioruJojbP5yokkYVLsFR9S127n1zbapZ73yGN
5R88cEjnrZjec7hHHsbp0aWEkEC4OIEdcU+s1kdpGwGeRZKqvxuXUQi1XM6TwCqAKiog9W9iXOSM
aPSBI/4//pBcN4jKQDWskbmYttlsuH1qRHkrBvmeu4ngqbouJFKUN7m+hPiRP+ufN2eJY9RcCCtG
TUv6NLuAD0mezL+qbUb1gA+P+18ihFaVDkHiG9Do/4r3veP4WKNnIxmdgeiQfayUn/LILWpm6zXS
GT4A9sk9AST55uUMCWc4KeFxh3dUrc3omj72VBmBzsV2oVRm9/pL4YDwZ5dIWfNViVdjxMJ40bfs
zXM/Nqdrq20DTNmGWtGQGHEz1X0z5btneDRjuI65Muah3b4495E1TTd8Om9tI2F0z0ysbHXvuats
qS/R0fbixDEMykRTmkIs6AS1UiMuTOaCtycrJOAYXUK8DlMgA1SmwkVkK8kH8WK17laPpKSzLxBI
7QqMtz2N5uv+FVRJjxRAAYFRUp/z3GzROhu2seS/sEKJEmdIv8THermu4Zqt7UCetWibG3dbJUAq
BpMcN0n+nsfDb+EraRj8LNxuQIAAplyvKB2IpsnIkbdBVLaLOXk1mlDumJPMnZdRy1Txe9cIjfFp
wL0BdBBmtt9xI3wxilzeqluGgSeIdcxLI53z6i/jmpdp1GJptghA4ZFob6IAx6w+FmldBmNP3q9L
ox0GiqHK4uf1l3hoEa/VLBqw8iUtXLEav2IlGj/4ClACptX9qr1Qyro2LbMog5xiky9gvlLcx84c
EQcaoO0NAnOXVCVF265LtqF49eEUbWkEbgjJOKTg4ME+YXKFQb0UNosSrVxBYlxY2rnIOZ18/SiY
S8icPuX45/687zBN5c27Wl4Asos9FFzyv2uMKNAjVmAxjnikuxOKfoy7UsBABvHv0dmeff3oGXbX
EcPHjeJcOTFVtI5absqKpMji4NYxmWR7waJv07HpdV4Jgo/qxFcR91aNOFJaJwcSJpXjSbqDI/s2
W7DaPQIs5N3gTTzKWPLuKh6S6zkXhMmoDnZw+4gwb8uu0OyUWgHHkaTYmz5NogMva7fZsgDyrPfH
5etOpQc0U3c9s/9Ol1DtrEISVVsd90IyRaqyjzjYr2Jl8/ZRY+/qLJw0BrlixaBQybFsayvNlIY0
HikII1oAlKishEuGDbnMjIfMf9knewpR/GeAHOOMBfUNM2ox+NpqIX7cu1rPor4lIi731NZOVUoz
dRa2IqOtHa76QJ7gXBC8meiDHxia5IZjT8aqX/ZbQilS/2g+WIOFQeb0t89M0zm+mXbOKcxvK1vW
tStQZ3ss/tE8sDG1q29Z6Q123/yCEkLiJNgFBAta7xukVSpnBA/+2S+RZgnI4uMRWK48Mkv4bt47
jW8t3MfYQX77yqYarVut9cm4dM1DRu869CJ8ZipoX6MGmMdRhbOxbroBSTVml0vaz4rvfdFGDk8G
yF52lZPdLqTMuMxy2WV20oJOWCbe85j6ua0Cfd4DmZEfof4yzElJ/027ysVon1mJUZ67x3UjMi91
nyLinJbigxwaouaPGfdoc1P9lQepYxIdyCIFSgqJQk8pV6CknptsBHIR0YibZY0L8Qsewu26Y0ZM
1Drqyhb/T33TB4ypL07xgWE+9UwZrsvoVIkTYSQsM1hiM17N3JwKQyvHOCzCONnHgeO9Zjb/V/Gu
eFZzVRsAtK007AlUL/pfxnlHoW/l/MHvhHWt8D5Zl1qz5Z6rKTULRZHg+7jNH50EvcLGb2sC7h9g
NndpEYYA/BIitvbLFku/Ahz50QC5f3Ni5Uue3vZHnzajjZn1c6jUOLdxx8JqQKuewj81JEQ5MBGV
xlO7zEKiyR4M7XVFXF/4vQJbMZsz9+6fAsC5AxJbvjpnwhK5m4U50ke97lmiR06SkNwI/4pqRJiK
uwTwyFJrfZiOL0A1v9rW8CKMVtWl+VJZzYDYDYDKQjac7ZU6qPPsaLqa3P3X0ZqIBWUP24mbeWzQ
IBsdE42O2uInLXIUmA9EjJ5LLe4O+vSh2N6MLXmsRaWX7u4GF59AisZbBGbTEd5ZKAudH+pbtvXh
/A2izaJugBTniR12cqjAA6EuCyhTaqqcD5jbgO45aLm6aKjuAUsKhl6zi7SmZgKFXbR/G2IJV25p
j1D0Bg/uEpINSPYlU+NZDGXCU2bayji1oz4w+iOXPt9haqelsHhsNYniRfyy6wMbNO69ak9HTPwa
0nRiGdL89wyzgCmiTPVjuUYLrodonDSTCf/8syyLS7TGOdsvPWEipcPgkTj5l01XV9/wa4KyPeIf
OU3oSUS+OFqa9nMmviOvp/J2OduCDX16KjJT0x8jsZCJkcbESHAJG3LTCu0T+OlotCqAm8avfX/+
5eNpHdSHGLl90JhICtr182M6LizkSLubGi0K4jNZrjb3uJY/Agi8QKfEiI84lbfLqSsHMTRUB0rg
EZYvWpCTd5g8XEsSkde5BrbSx+WQiLOMOzj7LYpeMBgh1SNvbbWKZOdqnymENKo6rYhrW878+7zG
DT3O1TPyl8M2wJxRCpFcNdYbfiCDA0RShH2ZrX43zQnlv5/QMCIaP1pR13uQe9kjjCHgRVRXC82S
yQ8ck3yuG+S7Y23CjYfUGpIBDgXPfBkDVc1URljpyYE8G6pfKBAZGjXl8CmKfr1HW3eFU2jaJEly
dOHOKPwjKaus2CSJDchA79iIfTkPVzfb8JF+96m+LZCV0fMfszcxNp0sCfeLs3gzSlOBoVKshMvg
4kbHoeA01bHppIe98CZxcycJ+kcpMQ96Cr1SpGd7ENHbmU7ORIu6zRkBHNhIAqsFXyD1SMChyGW9
uNv/Nqi6IXP6wAw+dNR6pNxIcR9mVcEJ/j/DGHJmMX2ATnMVo/SIXfHwj/7XSXYJMfAbbmh0iZpM
hNNNTk/5k30AOJk7Khk2cTIo1VsKvNOULLtxtNHh9UmcOGd6KpYHrZ9dVDazeI4nL5AJcPQzNnWq
EGCutaYC28Yzihtb0+w/Tbv3oohf/4kINPCiWD7UetpCiq4RJpVl+5SE9I0fNpaVK/xdgvKpiHHb
ko4dr1oYNtgAqIzgLfBX/q4p28bEFE/P7LNmxsrURyfs8fffrZ6uyVOER8CyOpMBXjhoDIBqVnLj
yI/+GWllKeaqGFx5OwCn1RaxDGGFg1NxP5HDXhfvTz6JMexEdouUSlU7AhZ3kZUmUzFOgfqNNWWR
oinsdnRDrSn+nRWXjvAaGBDb7FJ016Tv8P0UFPMiFPlOXcrxZv7oyuf8ip0e8p1kSf7Jq0mkXyiw
DL8J3vOboNvxX/YsByRjn6Ggolu2KqP+6RFOoURTwR57y3/65CT5/j5RfS3v6lu/bytr/dVCXvSW
+CTbYEqimvaTAzO/u6x4RZiSafAgl2LTCJ4CFaqI4FaAL+RUNK7CP0ljMue8g1f2uFUpu2wyWS/9
ogYgAfMzgPIdNL5+0EpCQXPE66d8fs3OKgg6hp8Rdxh4oWVd/uCWXzWl/5fXlBZICROBTE8fYttO
MWN2SP3TBENfTDYyNednVk6RtDgKDDxI7H8zU+WXUo+uoTRzq3O33txOj99DBH0wqzxHf2asdlTf
m+ldG6Z0aSJO+FXCSP3Bc5+GxsuwQ3sG7rwzfRMYwfHkDo94/4kAADXZaOTnSCu7bOCFJw1ZU61r
ERKyjZGmvzazf3y7Y6vJCECyOs9KvtNpC62kXAuGOvL+sWEDpbTSOJjsSBUTYzXB0TMP2zpbu4wt
JrWLKxBD5rMI7o7vIzzscCtuJSIk9Q3+fuIg8TwlpNqUZE9LiI9baMfFIxVd/zreQ6gTUCu5aI3c
1c9ZA7QI+EDoflZyOyoCYSyz8HO0Yg+lISutT1I0Z9j6p5JdZ/3sGcUZ2N6S5c37x9O0l0k9l4xs
xfGFxbJuE5g/y7F0Z7Gb1iDLwg2Wt8t1tgKfWjZY8kWz83T2OcOBjD9TyPOMw1h7rD4i5AdC2Zn9
AbblHHcD4v3ik8ca6/gVvk0EpjmUZDlfCIhf+BMTbu/q9Q2/rf4W/QcXyWCcxuyQmedgHqE59PJO
IR0wwwjSLq9Ize/TenDqKwVSlBi80ExnQI/QZyxhZeDYZM8+KoTKOg2U8xzlWsPTweEwslF5+wsU
68gnyMXiDr718uEfmQEAspCyenYMrwooQRuy/WZ6CFHiFvqvpkkNA8qsnc5Aspj0sq7fq5BlU13V
0FT00arLcQlmXHDoB5DB96r9yjlEUlVpAvMZaSWZwZhndtMzs++suzenBrJzfwCVPS6hVBzNr1qG
K66O/TaLkm7obKNwhGqSFLLETIWFf/D8NBKuY8+aHQ64S8liiXLHAMidKjrW5gEjCZQ+sjS2ILbm
cshJ1Iung/GJiEV4QaNH20uNoOa4oVtVVX18t1aHUxVDoF0Dbaa4REIiEi8RuZNyiZPmPnysq4am
FxdxFVKuMppHaqCSglA/oVI+Y5L56hFaAOh04LfkhKOhbY8WApE8s5KYZYPZ75VK57IS3MzGJw1G
6idUQ30lkmq2KCgBhzoMLWYGAV4IfoEF77dNDMh7Paj12QCAXDiXtwBCzVvxAY1XWEan+ba6Hdfw
gK8z+3pcS7iW1Z5SZSnWnGTd6DIzsF27/PIat/8TCbMSaYL7i6V7MJ2txudWaa0KRq0aw9i4Bkje
AeBYyGSLFHfCveJWkJ6qkVC4OJ7zbKT9Xs40aaW+gbNDV6H4uB+pq6b9WFoATuS1v+NaGQGI3sGU
iU7GCpn1sRI0IKHO8DQwIg+Sm791YGBXgJgxoHOTKHlc0UZ7F33aPGhNcDtLUf2bQRnd5Qnu+cru
Tk2K1YY5JzfbBXuv0wFVoKaqgblsZ8kRY9Z3b23g2BYeSZPdCUXP3lozlEanE/jWBuGWUjagDl4p
1FXTSA4yHqMu862uf87l4OxJjY9cwQlr0ExEagLYGJn8eLWZiUQEZny2WbTj+I+r02EzOfhlCYwm
HbkzdXy55T4p11eUcD+MN0oO0czzEuBPILhwpAx9F1Ws3TxVILIbbrfsCEmlLYps895mgxIVdFBP
7WIeXciczsrgy/zfPG/muEsl9wHmmTQYq9SNuSnac79E1+hnpQansn4tn5EWtNGT9AwH2mxus3kV
3Suw1mNBW24gEEh8GX4Yu7nLTBiMn+yPAAhHD2sMS68rORrdlYoCTni3kqLXaWMZGZp7wkmZJ4J/
dcGtn70wTfC6UjKfcIwYXIhTxN1dL93maiJd44WdhG/WPviJpnLBHYW5wz+W4zYrpamAGDqUUyT6
JGHddyiePX8JH6Csnke2917Ynu1fqmIdiP9p3CwrHGGCIkEeiT9oSSlIAw8HSQzTa+JKOJTaZSrz
I9hbUHWB8SZvoSKXlsHX7wApbP6n7GWDvMKA9f53c0jqdme5o3u5AH6uxfgdg8Gj4BM/Nzuxxboo
GHiaoB31VH8ihMImbW5E9lW3pSPlStx26Xu2Bo8X6UAMgA3QP/BtlIUkl8Vh8u05uLVAa0NIqKPz
33wo/+7Rg9+phHSjx5Od6TQEgFbu4HG3GEIO7gSy5twtPjOATn70o5I5hu2vvbvDjLdIZG4CGPDe
9uZPYDbANSrsKGpWPJTIVDlMEEsai9wsS+7bfUmAwVPwXgUIPpee2YWH58ihLgIU/2AdlIWR/wcO
mNKMe2ZUVnYz9hsXdqwnYeiUWSrbvh3HPYHL2FlIjAoRQ6T7WkWoC2cuYSTY0HZ0MldyTuNW4aOc
W6TfPPvIysO4c8XAE5VLnkep3bQLY4oyMvgiLSFJg9u+R2vPjJrSi/4Qy40/Sp5BfhlalLYbwcmN
whQR4YKC7RRnoDS66wEnzzF+szVN1WGojaLwrQFJrXkAnfHQzSjj3fsJsOe4HBJwaLimA6aAZG+g
tEw2Ny6VT3H0utI6f9mTqYL3kpBte6OhmFdz9jwXQ4c7G6Om43pYS1rzeI8XIzlCE66nXxhFxVxa
Cl1UcMabZszREdt82QNwFu/b25PeurF9DDmi1+Q7L+njK5SsFVR3hshmBz/Ibe2L9cSU24jVPhp+
VNyvYcaoaZAhuqF90qTqhiOUm4TQV1X426ryvAo5m2ePNN2e5np3HdP7pmxPnAHP1lWPZjYnJNhk
WdRF47gsXHX5xRomJzaql1ABInLqpFzZLZ75U0q/Y4sDW+kIisGRZGlYIQoJ7GUGqOyrokxSzQMV
djrlB2fdesugFe+afHZJaRNyV4I5IdaTLCkLnzFV85GYkbuIcDmiWegqjCf9xManBUujVNAGC8jv
8egUT93s0OtkZu8iDO4iHOCfW03tK7fRdh1M58h/xsRwtshAbpALxkieA73As7P9e598ZPIPiJe3
3Wyv0j+wrRf6OQmLcKBxS3lZZmXUkMANuM3fVlnIGWulGY7q78nU/Zx7Yj8YKXoeehpPVbZcHFsn
5bjjJlJL9buvqG4vfEpbxClXwLVqI53f7oOGxoXh4Zuutc194/9Y4EibGl9IMwWXIVLUKD3j/2l0
Pw5i+4IqjKSVtkr5nLflr+00eCXkKzzeSF7dbrkqhAxJMZX6DUALAncWnUvxr13AoGNPlKnm2JkU
bnYqG2PRJndKeOE42hUx/4u7WJNXPJGZub7T4Ji3mAIb7c4Ziu6z+hc+5i79aoBzSyk8M47VM+pN
lCBQVjP6hYNZtY2rcHucMuYAV0h64r3w3axAVUlEIWg81zIkr2hG277SMpP3lUrtldyaDnxdA12Z
zjJNTR6sZBpPHkO1FAh53vnMDJzpGwq3FoKv4L+omVuV/Xb6GolI4yndXBgbLaxPCXzQhAmbuvTa
Kpg9m0sZrb7VwJ3gL8pwrO2aU5gWNJC+4L00COj0Go/aFN0A62H+UbLqzrlSIMOWDSOgChlTetyb
dUnWoxnyNEaSjg7Xytx3uJQtxmS4inBVXuyKwIqtYtZE+Jbv1FCyRUu4fxY8JqGI3l45tHsgz58W
smo2gdAdFAE0oQOUoV4tbtJh0yWLQmISfelaB2L4zCuOMygg75ATDdUC0KjSvjvd7RWG2P/jYSlR
FdQmMrnJJpZ79li0XwQAv7W29CYhZ0A5ssa7EA2euzW+DKD8ajPLK9ctFhxkhRu8P6u3tbwTVzCf
gBBzYFhrhZ8zijN4LivGKb+zu9Zrm2Qx/VzGEYp5cGAiG0gOzrKrRk++J9QIAIlQlwOUURtyAHVj
ABLQ0fvOl7zEnirGuMeqnAmd8MOY5BvrJHymR9C97rDDFxVBSu2Ozt/Dx9r22zjQuzkcKpR5/S04
0e4WDjyQAeSxsCdju35h3KkX4x0XFHoVvdIzjzYd88MNQv40Jimh5henEDdIjUoO7IIQbXJmDWhm
Nk/LWc2W6XrB0+N3/oV9+2scEzHcFX2KFWtceiinZq08vqboh8SrWPupZp2dobjDMpqVRzJwBFIK
XV+Twi4mIlUzEW9pn8M5wwnIvDLGD/PiJNKzg1pRKLgoFCSYGULCuO7gzaXghzLRBSR8sPFrIuFH
qfig2/TP2nhU6jcYV+REYY1aESTSpthZRUeYk0+DGbdftmZrpfhRROicvtC5N73bHKQeUcoaiEt1
h9wwwk9wHjoZ/44CJeEQhJOBaHYqVaeD/AKt+LiNSqVRxhySm9KYCoZ7+QjwUaqmoRT3JzqE7JPX
khRAi4QxdvVXXq9R0D6a/qtSiWz2F4bP40uKKAPHXSeEWSb4/XWpCn1yb756nbKqwXEaCf6xuE2M
FoqWHcUu+4YCis9Kjgx0V7eE0qV+wzVQnKtyzx8Pa4pTPPw554Gf4e6XxjJxnYHq+9Jdo1IDohEV
F2NAd/tM9o+aoh8KIQzY8QQDOc9PBspNhmVAXYGtZvYWMH4ElcLpRdT9jGsLSV8ER6LFDDiOyRn2
CPrvv9AdY2TjJMl5HyLvVkY2DMPogFYJ6qA322HM22gU7unKF08128FiXXCL7BQErZ5VjQkHC5j9
9KAfy08SOiw1SzPn5CIdRgDm51JmW+a+IicM6DF/lBGDJKWT0M578NZ24dpE7QofSKlKVk2gQer6
P4nnQ9lRCRoBPh096idlmuldLy263OonIE7hq7X5Qser/XTNev+CO5aV0oMsbK4arybKVj3W7yzx
LsyhZxbC6UCusArUDPMrY3n18AdFLmWCRqhK/waG2MsxcKj5bx+h/u0/rQ6lnvK3GVJSxSvKNEyl
VuPSRDW1nN+EsVgOATp0IbISzES9j5L4HOT6+zHF+ZxCuNcX1GTnin0HnwZxAueAiMEz4cfuav6u
3V0LTrUAx3cr4/GYSs9OlwXg4rMIMR4MzDg5fkac5+jTflQHMwpLrNlJR/7/IoW7CaecWLURfOeR
K89IXvDqjUHxTz8mOuMfkkYjpKUG/WM5rRBNaL9eiNKSShgAVrXMDOzuJLVacTNmZkdBx8szKXT1
VZ7yvsdqlwgZmp5Zyy6Wa8rwENTipFRXZxo2reVU0eZgPdmmQzoFu9n5fQUJa6QQV3usmHjmsJxM
DDXGEkgWuegtRfSPhR/BDqQVxCn8mQ8RH47AnwmIV3XHC/i2uN2Ac8qPmx8U/AEDqdN+kjnK/Xp3
Fv3ZWEwCEBF4vyNMfWeJsaK1FSJWS0JVL8tt/l0JC3gDjS1U/jOykRGHYmFOViX9HhWpEhTuNUZO
qJe58xp7ITH8qDUpxoN4W+LnIxqjJII1mqrrZxrLmyPZJOZYgiH25hoMpG/IC435We3d26AYS6rx
FKXqO3oyZS1RArkOLLDDJ8uYKKivm7maZO7sEQ3Eto77oPn3Oov58hYj8OBSF7v3spvkXU684uvN
3TA77H+g6O17zASchrcVt4lC29Yv9zIup+6ChUQW9poGU3xIhNDkOQYdH1XdP8+k5MvA7LYKd7BA
xovUPaX2wnI1lKSDxCd/rpj1wXn7x0lpIFEDIuF7eKtoYhwLAu7vdB62zUvyrLaKl4fZGoBCf5j7
mxlMuLb9KAitqTL0otllqW6B5dPpH12Ij+4+8Jf99b2dVL1IrxOlDv5xUSrIWhF19STuAyQ8UcdG
IrGIINQLbg1jYPNk8SMryylFM7Xj2G/t7MaZZRUreW6foZhISDJsffrQbvOujtKV7VwCPDYgPjc9
RJK23Amk975pozfLNw20NkXoazceXIdrN4bF5I23U/pMNqrppHDLVqpR6SbfuP5mPzT7rltgRv/l
ZSZtCFXPxHVKq8+EvkSVuMGpILu1ILIlyB3AJTqVyxa2eXdZgmEG+lT7pCprOPD/sOsVRX2r/6rP
QqCtn+5tets/It1dQfUPfn4hYbueDb+PIrMkF9kGU9c6fGJBOSfCcRypdvnhlUqXlxm+9r4gmTRX
rY6f/2nY6Y4kFHM4Py+JsAVowEXAABtB87hfbnIvhKeu0GtObqZKugfghKrZezASfbFKoduN9GOh
nEidFpJ3VAGXj6jjgQjm68RE6AWdh0jT5Dqq5bdb4VApVstFdNQR283A5qnQ3qH/M7WDd5kqP5iK
GcRGqb8/aOhOk7Ng9+becGEwjNvq1emMpkFwEI2Ff9SrZtZtBSBFbi+0pX2XWEwWLbuTgGZeRBHS
l+p74qfh/W1oX/oEggfUy6qX3R18eNLiQSh+Yc3CuDgCg6g1kh39E4wkRFEtFEPqVj3Yp22WWRRD
ZWAzFkEwfLxHNSP1zfcYLhX86Y5G7MSn/Iy/i8kp0u90V22wESQWedAs4Qk2G3MMrv3XaC6+IgDH
5zLJxIchFp4/34lB1HfkffGCmiUa1gjfg+E6sJyskO5AbmYRZKvQFptqTIyDKzEVRLj1PhGyfq3Z
10HZYX3yWprhgN7wzDa3OC/hDqbmDEsfPtfOv6JTTVaUkCmf8lzIF5Shn8oArpJH0qgXa8u2MlU1
mf+i2YpsCqhoKLwxuEN+tv2PUFHyR4WmRnAasPD7OdSM+XcX8VJIdTa1qOY2Zue+m2nP15oC+YvP
xPSYH9DFlWs1OOMOYqThjtczFFCXL13kGAOEUar8Y/k58yxWtX26R287rN6F6WN5G07xNRw9nG9x
6hKv1+U5BTXgTnTLSdNxpnwW+JTZemDPsL3ZSX3ERzg4630Kk2Z4dYc2BUNIxxrU3Khz2jUAG2Bp
RKA4u+OpXgtxfQBH7KNvA3/t5LiCpdEDM0Pb/zdOaWhMMJTflb5Q3pmYhq4JSsuY0Bggn2M/xXee
kzDQlMJcQp0eZ95wp+iLmXv9/jacYkrZKInI4aNVL7guT0FcP9uhGpGB9XgAZGJDwu31RQy2L94Z
xQwaMBhDpdVrDXPYWV9lKcKl2vYv4pyaaId1zj/j69N93dofurEHWtmzjNvBGY/Apsp3Znso8nQq
B6+6m2oY2PLC2sk8w1iNvhMk//GuFRwzb+A+MwYIirgdetnFBQqcmc6FMefeReeYmLJbCkYMblJY
srd90skxgClgogeYkDrBnlx/BnkCf/WyX7iheS4s59QgRmjD7I5jhnMDxWNPXi14RuMvWkLNb/ng
IDuy6oviIFMDSmsmzTi8HBYcTXwV8CbstEiV5S9GAF8BHk1XGoAyBoEJxVJTADyRMlInJxQJsotw
j2GPpxASaHPxvblnWNe9uUhgRAmC7J68HdSAfisAxudgmhDA43qFshpaYKhXu/qhnfslgaNjhJcy
1bK4aza/mcte0zqnXv3jBJc/RS1rfxiKMlJIlRP8WZZ/HogQ4UAAhavlCsvmt0uuY230LU90oIYJ
p41p/4pvn4E7UqXUnzrgWu8x4d9U3GPisVBVkDDEiP93lJCvWULDV5yQU8xAEcMTCHfHuQGN4zS2
9j47MDx2VJIMZUaUP2c6oo87UaF15qqZO68iMk9DAXjEGCH7VYbB6Mjfu98VuR27wQ4UfdasxXuv
G6yGTjddy7QOaQqmK6cFUxvFzjV4NxsUtKE2nEJdJ5U22KVLoJa+GfLXJYE+AiEnFYNi/KR7Mw0X
AqiJqARNxhaG+pGGtEKMM6txPP0WPRxWYMCoqMDjjoSXLuguCBY6s4ftCiKQ1HZYiMsUgEJ9ZaWF
XPtSaO9WbpWAo8UuCpD+BnDyM+Eoi9xVYNiF1TKiNmLWz7LNiq+G2zjeMlsdbfxw6vxguHgmYNVY
6xJ3tWrj1fg9LrCw8Mey8DfeCy8Zwgwv8mWBCZyQ8g7x9zYH3ep8yOLOedQD2PRqiryPGP7z/WMe
V5PYMN2PO+YMAeHz4+Q+nSlaYN36JG1iPlESq2wmMOjJKgEEDI2/C6Dpmid0/8BoPjMqeJCr66RM
3FOgo4/bPlCwsd8ogM6NTh4e+P5eQUBziyIdCE0yW3u3B23sKAJqjazp8rG1I0ZWX+Ff2arO6w8Q
grNo+HIVvjytLDkTzSo54zb0MuGAV13GZ8AcDX9qAzwBNaXLO+SWhd9Ez+rX2Tn2WzQNFQHQSgEA
RX1ndYyj+YbkpTi8KrEI/BG8ZG6eeJ6dud/g4U2JVI9QqJsMxdUbNz+1juoGWeT+xq0ct7uLzpGu
77LfHB+pMKaEl0waXcEZUAWuEmbQg14Y70nhutTCwszT4eJ2puKPYlkvjEyHJhyAS9IDL/hQjO7M
CQGIXYA3R03HkwtpE8Gbr+E/tSoMjPlkKn/28LPnFpel8vE9pW9/pCdFOeLB684H67lhsQ0Oqyy8
qwI4/fJwteiasmbnrqvZJZ7HHWDynP00GAl7m/ylaf+MFx33XbAq4VswenHxNieHFbPoFnovRhFC
5kq9THj4toPl5ACCUfogkXzhdb8D8p8+EzTCkSE7MEtPG+TWk0zxTIt/fSsd+AESF7EYyelP8jG5
czB0+KPh+hGNw9V5iY+Hl+RNyZMgKb0YzZmz2tYxeJlyQJO4Js4Nte/F9ZtXhEih7LPtqSUXrcX2
kUQgx6kXw8WYRPyZyEWrhL6YTA2mV4vhbRg4VUlSB7fZFgifvp79uUXatl4I6Q+rQ1UJOc6v/Urf
hXeva74+yzbUt3FDHcOSZ/M/vSXVXhV2U67RePL+4xfP6yY9ci+XSRotPcZ/cH26o9+82z3I5v8S
opS2YuwagDKiCNDeDujUWPYCrHFctsMoMnlztizb8GDYOooUZk2dD8XJ3Eb3jy3Aw7uHLjVc/T6S
OJJGu9nHGoLhgwGoHeohZpZHv/7ih0Q0YpiiuOVFNh8qduLFv4aj9tD7975pIruvPxcS7VLu2KUR
aufa+DG8niGZ6m+1nLXBVoeqYxjhOPsrk+A8OxctDVAKJclvSFKTLYAUSNTStOtoLENWaZM/ImQ7
iABElSJaQ00m0C3n8+xBt3dGK0nSQHrQVRVNNLRViYMCgGjkdSVmoMDZ4KiZ0XdojDr6qDab75bW
IEiHINF52aLfHQ5HjVNt/EhAAq6hWnUSH52vv3HEPcN7v7XOjTcpcKv5tcAiLrkXIEPt562jTMAg
ttgtM1FNqgmlEuXO2kc9EXnJXIXMeDXtsGEzJFL+Pv2fcjzNNufEt7GqwLlMnctOsjP5eb/Jo8wT
7KCHdYQu3w+ajm3oRVS4SUis8a8C1XmF2cxdZ1GiCdEA2NJMofu1hUB1Cuv4K7K6kovx5n1vkBa5
5HDYhjrxU5cFfovp6vCGLHryzpRFyZtQmRy5lXQQjV1jWLEsA/8Ef0U4cOFCf9vAlM0pKh6DU1ta
Qf7BE9rbT/ubG8oFkP3/xjPmUZJZ9dxf+dJA/EKRm/roHWTIpy4R6Tp9YanFCd5BhZ63fn8hQ1i6
yHd1eHv6hdsLS2r+h3dBJLcHwSc/rYiNFStGy6zVxsW1Ubht9paLijpfTgLXU7cdyr/0SLmew2Nm
K/Gx4fH8P2nrET1cr9LkfsM+mFge7bNpyqTT3qIqN/Z0zmhnony2qyVJ0uaa1b1JKTnVkRvGvVMn
b+s63MBVEPwCPr3rJELHNENs4CTCE91tu72AHrSP3KxG1ibQhK+htvzg1gP0YXTsniBIpxumIBEn
idkaGgXUS5D/VJe8BSS5yr9SUXVTUQBZcPuYDxmeu56K7tBF+kv7RB/wOtCr67WeC0ZGjryVm1+/
yo+nrvmYU92XQEPlDEA8h74uIpN9M4anl7PXRoWwC9UMT9b6WxWxo6ONfUEG771VdCxZa3bdF7S9
kYG28wxKOSeyUvlbdEqpura2ejphKDGQLmhDV9cESzymbpIXH3EBnQBHPZFbfM5O2oiHdjaf5JO0
NeZIpHyALcdyvK/VmAzqS3oujd26HzRxOVK2Rx/GQqdxWNDM7TC8xYXs9VTC5rJV8QeThW7fLbZM
6hGrIo13ypkRKG8nrQebo4CW/C3PEmQeJK5R1wIwFb7th7LVPHCE/MGPSXFOS21rI+rNaCaFDjKx
clIm/x8Qi7g+fqxy9t1kuuks0WPwfxlxM0bPsSR67lAIRJw188cvKYto4g/jMWWDVbnztpdtA/CP
V0GCyRoiBVeF92R/4etdiG/3K4/0YlAIdd0leUBBMBkRa5DsPeaJel/tBHyKS7aUr0LyOd5np6fa
jeUfyguT/9yFCCuXphVZEO1oIERpInpW6CjIGQn216q03FO7ovUo8ZPh0RgZ3wnZWv4kpQQw6Izq
aqOOE2HNP1aV9Km1jQuiWMQHcg0qjOzOplMMsI8iv617Yc0mn06WMBXNkM7btvSLs1JID0m6tsQf
vJ9ZyXKTSbFUuJn8hZYEh+BwBQPYkJ35VEhn2RgUDBYlxSxtMWOnIDE1e82BgFQtln61jc0xdqd/
CXtL+ihmXZ8ySFObU4RoOJt4H6RG6dfvTB90j8fHoO87ZDdrESnw3No+3YmbgMSncgPIhimpQY3z
jBZldnNJryMv4Qov2AsXM/5+dUuETeBaBtf53WBGeG3872SUG2EDgMz0rtueMnPrwqbTC2KvgP/4
DEWsKy1hW1CLHVTvxX517ydTo1aPSrz4GT1XB5CzdntGVxiqG9TFmhgcB3pkt/0OaRqBGszZFEPx
rJ1yOzLsu31Xm+fUvehGBB2govo6gdSrHcCzYZ6vJpva8teUp38NoqgoG8eXD7a/TvQQQqf8ohiU
YUeBPks9MW3zZzP4yoh4MqvhJw0BjzVG2rQ63+ARQ6wRyP8yCoJ10t7DB6J1mE2ZMPZQnY+EwEZI
mweHBzNG6VX1hIHMoL1ECz/wAnyKwdOzwydLunpWDwJZ3PspUZzcNBjVdh5xQH4aj7ygAd4fvG7k
Bjsv8Kl9tc4hIWY5DeQUFl/KhMybp/nB2eg+EDabCiNTVWsJP/27+WBLVYc/kUM3lfGv80jzPlDC
dAN4EHU1tIcpcuZhEnWTO/TOX7tba1iUfNAW4SxMOJP+A9eRNAk+imKpgPxgDNKiPd5psGaqZ7kq
CZKEM56NVMaE63NOc7QCIPfoXMhG14/nmYIDeipcTw0Aftlm/FCVbV+7qvNGaY7IWjFzIFPNc8Jp
AIufAcTjFKAl1Rlwn8cIbqo1Z1idRjCB1nMhrPw8L74/jPW3673D+Spjh97yKeVL1seS6BFHnpv9
nI5+yYW4nADYKqWltQW4yfLd96zqxSsNBBX2ng6au5He+ukbc4IT+HbozSgObxA3aRgQ2Lz+W6IJ
EI+p9DktNKyxXbiqNMhg4igQ5PyT7ggFyu2cqpqziXmjVRaTo58evUOfqwTvSrfoT5ep8qCsfFlP
2G8QQZpVrYCb42Uxv5j1Ig2eDlripeNg+ahopjcLx1m7/v+ZWYmHQeSX4YKymYOrZObTj8VO2WZz
aIl3908pP4kWmSH4qYvveJIJTPpt3ReXT60P9cloCTXfVEm7CzX9jxjBVxjyi/xgryvGRmn/5iq6
7CzfhXdVzkBMMJ4nyvPif4fcWZobx5KZJFmGQqOICPGhzG1o94m61UtTXAxgWL5X2b+YB+CE+5mf
kpyKXED+85YwLA0mRPwLg5VGtDLbveHtPf6SPwIuWmTHdF4raZE2kINV6AIfQovNfIJFicX1H4Q3
ezFjd7NcnuvBybRC8E22OpkOkmp68w+PiuXQI0LCj43K4UO1ISBY7C+/9EanG8pRMeatiH8BPWOA
+sdMCWKdemtmuK6E3yE6Ji5Z28cT+LveUA5ylD9aggxTA3W9uvsg21w/7R9+Y3jYyjYBB1OF0xkJ
yxqI3K0O0pg7dMXgmDV8c4aexbUk35cbu2/c3QlI+wXZXmG371GTwMnMRXALsXWnThrP5gNELrNH
IhHwP5dDM5M4ciYqNb+FR90180VXx3utrRi/YenjvoIAvSgWcxdEwHtQo22f8PRLT4CbckFsBLK8
ova08ZfDVcEh7oxNgb9gBzLo6X6LgGwaGTewbbLb/yO04w62prlxUwZmdfWxyxMZcSct55LjKLMm
pSXDdmd7TM7v7TRsnlHNnazrIJv55kmLxZEqLHW3QMY1hNkcCcIcVcybNWKnHCq1iT+gByMFPgHL
oJ38L524zmjyRSx/2iPPXHJPnhGC88UtHZqnHRjhBiHt77M1RI9Pg5IVoS4Rp+xetNx24pcIUCLT
X4dam+jbK0eLw/pvsFeHfpA81pgT67g0rpGVmZ1e3uKprCorAChZncGVqQFyeLcnCP9mxhsZtYcP
2Ya5XHlfB0MkB+cx3j2K0/S6o0kkOdnxTJhv8bBlyl9JC92/amai/x3UvuThi+KkuuNH+3PPf/Ys
y7d6BdOy1P08Jx29CpudQD+Rj1Qjt+tZNV0eUjJmS8McOu0Cu2lCBNYSMIoTIU2iskcmiTf/t/+K
N9PmntNoauZ3rP8Jb64BSwB+HrixDMb/YJM0PAWNS0CqWF1G2i2853ZBcu5l32PzYKrxU2nPdGs7
PLi29f2XTs09X4MTQc1S5Var7chwP6oETaxfAfq37jgD1/W8ZcEX8Qht206HmUKivhH/EQ1aaxL/
PSEUoKYCR8M+gaKPug8pQOO61naNuliiAn9q0TsoysWuBjfbzi3NviVu6bG4wkXtEkEoa4swyxsZ
Cf0Kfp0f/XAsgiHB5uZxamN1ew8S6ASMDsM9PCIrBe5nA1Ub/HAcIo1hcgAbPOBFvSVinw/gi17l
2uDDh6MNcLh+3Q0Ry+aUnXWimmp9Ivt8PHdNXsEMXl46524mp7PqfXG95omhb1sPoM3wZW9I0A4+
+djJ4uVUkdtTcLIGL/3T+pxeSr6Teg2kuRLYlEy6Q0kt0eMz7bkS50c21uhpLitlOXMaO/L/QVqM
arCFIuMko6e03DP4pwDwvw/eaxUF9+3QTThr68OCUl6LShvEZqi+hLqefbYbkmWO6N3eRaPAR9xM
xOiAMLlEKTImzz24N7m+yN/MQPbQDkNDOnXJ92Jgft8tnsT2VQVcIAgsLcegRihVBA1SV901eAS+
4WYvQFx5k/xh76RqEY0hYyVtD5haCeGCjpoqYMRjpZGqFN6X0VBX/9CDEj8vwblEvErMo5rXp77f
bm0pcE2gjVyCBveuscnm4tgh0Q7q8n7UIGX6g2bPCVzwjb4a0b4DcUMqGzUKCfWJ3wAP9p63J5on
56xfbDtQI5wLw71IWb6fnuw1YoLG4KbbWygn67CeUa8pmDOR7Sl/wB9p3REtRU11HtBToBUSLuS7
ITRzQHzcwF0ZIr0+hbEBjyK9fL/lS8c9O98TlWz2iDWEpRgscnMITfaMDGtNAHs5gyWFVtaPv/TR
LJS7oHk+RVpnpmuLxiZNetJdGe0A4tOdf2WWVinDZqg6HkaFa8FfODWf+rUHoLIjW6slNA9D6Fn8
VpV6pDXLBhI4cmyadeZ60r8bsPQ7XaGd14D1VNum0FVwKfYLnXGIizLxYyQx4Ae8KVc+jRfd+rsL
wEqDoWzzTKlkPgrKPuPgE9goHikMtI9lkxnCrRTaxtX37TMBDa0Wiqz4nkdd7A/1s8CjFaLn1KJ/
RVxY40v7Vuo/l4WpIUkF2fOniMjc2LYDxueQ135rosL8rbKCgZw+ZDdWS85Dn7RjoXIFoup+GTEX
CgVk7Lwnt2pn3pRG7BNL7ZAhYcE/n5eveToQG4Ie4UNvvtW/n1rZB3UdqpALPl/tKZWFoTFk3b2N
O+2pSYoLfDUwLBlZJNNlUWk/CEjDOT52UQonntkiAOO759TqOw6+0GPgd4yHWF8ey4tyQEF60PHR
tvSfHIevTmtq7CubWtqYWaPTMkmRFDx10ihPwcJp3z4YwLoAMHL1VB+LCdTQqP/pnzOwBr66LIsN
KJ79qYgRFyKvipKrkik0E8XaleDjzFY+czbsrTpVisMuUsdU+rAY5C9BJCaZm4GRFgCqRUQcVuM2
k0yQ8hbt6mjLOiOTKvnciVHLxR+jwZgAkPp8d0xAc9LK17EptzRsa+O25aidGpxzcXD+JvRjslFH
RJ3IwpllgJKfDS1xf0n12UWB9GysNmvizjr/L1jH1HKTczrJryGIwJ8Ew9UMQvZ14jkPNEMLsQxn
In/2lJ7MDnEVSkli5hwvsGBkPwflmOqzAAtMT3xed1bszlonljxXUx9YY6I9Fjb8K5G4KIHKMY/I
Uixa/BuDcywUMtA0y8xD/llJRJQj0365fs53K5X6uYscptuqzSxJxZvosjBBxtM4SdDyACh/sxd2
kHN3juN/vr1hWfgOJ+QVdl9s0j5HPHgUWplDvxIg8jXBAWXZ5HqN5ATICDD7+wrMYNuU8ogFcsuO
NwGvuJvigCHJrjovT09qXnn14TVGz4ezt+hB7q8XglXjVHx0mG676aQkxdK3J2EsdT4oZ7adjKnJ
ao7KM7fnkoeZhL5OZV5E0srjf2SECsxcP9cq4Mwq209UiLzLN39VcGQNULBzbRT88PYTKTqifdNe
ns1zu5LMyj6Uc+10CrU4mIJiQyyVebIqMVeq1aVoRH3gEYjeVg2anEj1pxrj6IUbji2LG3G+sr2I
OdRT9nckYuopcNSmaf2lg9guL8A7Es3wj6JQrLWRrPxHnpMvvmgLJmTrHDVlFcsakzkQXtbrUbU9
qfzptAHpubNXS7Ex5erFxQn27UET4uc23EBse0TtYbCA4+VF/WsaZwO7gl/TRb+JhTovfEKFuXxK
+1qh3+pk5/54wWV9nIq8jROynYdRUHZ5q4Y0w/BiLVG3rw838AItnM79EJEk/kDcI45s66EeXtrh
s7iwKVKn8AI7YSdbOZzFMTJ/AEviV1ErOIhPnZi1DPYXxcdfMZf9KVNH8mOOOnPA+OyAqK2LSJer
kpdK8S/+pVx8kVV1GpQ4o1gR29cxmSeAmb0/rIbjC4ErhQklmqLptQBLNxlN22AwZXGkGSFMZtI9
CIjY7uhcCU/tJ/fzDeD3i6lbEJNtEfMQXflIn5z5mS4kasLb6PGKEpqB8pK8DdeMRAGdOTKkwD4d
axX55fOP2UMHCb+ZH0TWYwVIDdA6RAUiEyRJGDwWw6YAMbFEUIMzreX3BPit4Qse3UheBrXkKO6m
19O1ERIfi/XnM4RKwwuyYi+JZSlj9nE2VjwYYzUWiqkhT7ZSMNA/mFCrcoRf4hg79XJs7iZhcCQV
H4xclfEon6eFd1yGRQcVU7ip2tjcS7sfWn8TpRqK2EISJh46re4XbyH5zajemO2SA+v47mnjhdd3
wS2aGekeg9f5PLbhJ7bfnmUQRAESwrx24R8fPYkZrDKQTMIqSQPNkWDBXZvQajmyU1l5VPBDKOj4
VZUbv4EkILZJcz8Rv12SsHg+QsOZ7D2WuXDiM/JObTJS7tazSKMS0WpqXxM+z4+N0q2iCS/7BW/+
x4TR1EqhyRuvFMj2b+tpNUuuBP2a/M+Qk3EPoamXFeAlMUBp5qy79j9NBmkuEi2QplOVVTbShBbT
IxjJXgCr+mKZn+Ul2agsKUNK6guJDZYqpDSRgaeGKa8BUd3hyZ/I4kEfnWBWvln0PHqhOkiICCMM
5UK6SOq/xctdyG+iWJGZdua6/Sjd9ekzKOoBhaYfh1xNWgxvROQjGvNdYYjVT+A1rhgcSXykcbiS
DGMt25RH0q4aLuobJ7NQXdvoOZYoiKWoc8Wwufn8B6m3cq/PMkKTE5Bi/4UaKkk46e9io63YzAVm
D9TXIyeZZZYpyiSVsJQpnClgCLo5Bh2lJvcPDBx4QwInYIlBF0flHU+TmjvhWmeH3s5Aa5z8lrvG
GhUKdftL2VLJCaic3ZZ89uuc5vS9Qtl+Mlj8BfpwWmGHXKEBnexgN8wXfoYMCsV5iPQTBNgMGfJ8
ljEnMKdCoZa9VgZEBpad4LGfXx8tD2y47AfZSv1p+BLGWqYvMPHL6f2Gmwrd9Z9m87zoKmj/4PKU
fi+KxNNX7pYD+jw5Anxg1q76cUqBKbLm3XEiWj6XsLwwsq2lov3g3uxkE6qKt6lYzHygLQwOSt7n
6eZ5YQThuAkftwX3ebiRxLSZHZyOeAtettqkGQ93P9E/aBExo6ctXPHckITUGKCsNfgLHfbAUPHK
RnxtsRlao8RqxvGBJL/7RRFAUx1EmJY2B9ra+ZVyRf56VXL0D2eFNSCqgbmww/ejcI7aFpr60XRp
ABHaFBDk63INQ8gR3W/+1IanWZV68NvllL2IhJDt7lElVvoZyofGie8s3zY527BAfhMD+w/UdNsy
xPDuObelplZvvTXHbGXBAFguFp2TxJLvYd7yc6TmCNlkY+r2JrIGVuWhUOJZxw09CDtmtSuTkF5V
Micvx/DWmpibQRNCkIYmQzh7sTeW7NCrN9Z8pkUrTolPFbSVtC3gPvwZZVMnhvWiWHWVHOArtVcG
FZiEZqahWUW2vJiHQ+6WrfsQgVB4bsgwdc/NK2Egs3SNOM5NZYQaX78123GFF8OlybH/Kc/xx5TG
FFlNfnOOxLV5Zx23Y4A3bk40N/QCTlG3YrdSfkwhPYNTbvQ1u8HMXMslbVudJC/g4aifkTSBXPV4
UH6+5ENXr0IX1EcVgIJYmjpqxIUB/WAHsF4wK9lsIZTLZhrh7vaTZiqG82TOjr3g5lsfZmRe2WP5
X0F93wcQTpA3SO2L9GPl8rWAqcvN4Mp+YAU/Nj8aTOEcJ0tlH301yzWdDB/uD3FKHInqVyFq8uSH
v3QCsx0ej2mrgJ7mlBrXQoRme2T7ReUyD3gYcllgKdpBPRXNzcQXGADUMV8sI4gIsr8RhV+PoFwq
FEFwU3Vmvdm/lk2tlcAYYHnTPx89KbX4yO3FMzBuWWuhlM8bTNnKtJEaFxNjskNwQWBI/4AsUpXv
Yizv94NFWyHHnp3BEJ8tPxBop7eI3T1nzck4/urGt1K/0JuTYOjGmhUDEb5s/r64lFtvCklSxCn2
jVX9hXq519uhQ5hlnBSLvWkwse/gvHAw8IbgZuDDZ/wjJz2a3hC5wwuUdYXz3DCgK8+zmo6vEapw
IOfiveG09xMClfrBJ2lHvySAIGRc/zW4XrJOeJWkRQyoZ9M2WBjMH3LCxX/93W6+8NBsioETe8PI
FHBqjdmCubPLJ/xH8ZFvMCHvM80HSNakyUHnJdJB54InsX7SlUNKSnn6Vdo63wZMqVAfIxZgj8Ey
b6jhPPFB+adEv+eBS4YX18PAf1s/z6G+rejRGPByhor4RizMSPrPsgXxbGmjFGNU4EGxBTVUxUhr
MlYou75n/NRlCtDMIPZi9FfwPfwDttj/nRD+hOT55svEuNIv0ylEtLx05qllZncwfPenC5LvNElI
SYbePCLPhQeZDngkGU78++zaaYnwmVH4CG0lP9LUU0VHYJRY3BljaZUPnhT5hkG3Jmsfifvg5W8G
CTey8v6oJ0T0/ObNcTtk+A07ybIhzGCWM+srF/CaA85d7IeSEgGDlwXZUknS6uXal/xQYvYg3sp+
zIESe3gS8drLabzDtUHAsLxvAlH83Rcn4DINy4ePE5kkYCGv1J021d5KVZp3ev3oZMyq5XGVGPQ8
rhwDzIKGv03LVGBuOZyWxmYmpeLhC1L5Yd9UF2AZN3OcVdmnmkhEONO2m229qLoZgIRjDxyQkMVb
6l9g7DRC3BIRNxa5AvHUYV1hqPGKxHEps1QiD84nWVvdRNhoj/p9sNYX5bZMfQhYsRvo9TPsxM7m
CuJMFh94ki2Ka9TL/TzPsu7GDYdOpkPzbe7c6qHbLJzWjxWjmzjvWd6wtBSaPHvZQm4RRzC1rrrv
8vursnTDxNHP9rt21tRIDVbj/4ektcI8XsqeogEmVk52nBRwCr2/kZ6zh0MWvSe/akfRyHYVfI4Q
+P7om9U6SDDQbKUTlOPWTs9bYZTtJCoz/G3DOBRQsrS+Ae608HZwoQz7C0qCntgUxm8i+G8rL85v
X67X9ukSyIeiHrt5NnfvYZrGhNqlNFd/1A4/fIUxkZYUc3WQTKRHnMEpy4pk2BOTNtFVK3I8dJjo
w7/UfGihxgGqQABrH7Tdum6JRaD/gZBQb8LCXVLqiTzgdcshYXqAfoqSXpa8exCvLQTUhnQsl/C7
RCVJucEP3okqqN4Q+FOQx7PdDJkWcXkkdmRNUjVQCSrNGf6EioTRulGlRTurD1i8rFlMmx+CSl6B
KTzJoIfQZqxbw0EqK14+649hOtFC0AE6n3c6D/Z/kPfqHYe5OsK6STIBMs4o0dAlCgO4K+Wyrxe3
uPrcy3QdrDlgrHBYxsG1TLvB7p1LHTfcPpcgkDBdQxCJpjqBEpvFbnjHTPJOtsGluv/W1gkfcea1
CqaXiVrGSNfAqCZjeP8hQHk0CY4k8aDq5pE8txJjmDqxKsynE+e8muqXShX5/Sl4aOA29IQqLwLm
w8aaVU4HjOm6VwYD3zDoYp6qnYuR9BvzlhE3P/s8IEB1pRAbVtW8hHcsbNPGZc7FvhM4CnAemxQU
tP1eZTFxU3kgzAUnZbrptKNtn4V1p3N5rxhwCQ7eTvrSvArC7ypLnofKNg3XkRwPMbxA8QWnIFZ/
KjkW8def9obDSZnr/Gr0RhUe58qRNsdf8wLfv6CB5pTCtfceWmqdcnJvaxACD7amrYEokwf7vZou
ZQYTtEq9rEpoWhSMQOlZDtQIrsrHwPc1ukAXbLRdytyN0kc+jS6SLGNrUYlbVMQ64sEhICNqok1m
4/LulGNynHXSNn71FIuALALZoz5k1FRNMa1ZIS7WjCSMbcDcLWKUqVNGSCMBN73UCMOI4SJZEj4O
hRpqqb8wccwfMLiTrBcSi720brI6wTf878u/LpawcwXADuGPjHrW+ks3XeegVH/SmIEZu2/XGi0P
OkScm5wSDSfEZR79K/5BhU8jgRXMopfHOGRtERqgXCHJlHyqyzSWD6DBdqk5LKvslLrUELtRQY6K
3jxGAQRFKuPyjvYmelCh1Kewod0U65kXgUmevXnCE3m2VVE6a4Lohuw7boG3jf2o9ZVC0QQan3nl
F7qVcFtJHwRYzLf7teSZ+H3VrayoB8bLKzXfav/kvEiaMvLcxXy6nYOsmElEspxd3IAT/W3O50fV
1zDKvQUIiMq0LizMH8nGf52APrpYhm+G3JHXqC8/Id57DNJACCKOVtT+2DlHmQPHgrG13Ni4aV/5
2Y2URpujSDE4DYEdXUJhw1ehoLAPns2iBTLF83Kb3Huenpe5tg+Onjb1ucNzH0+CDrr4yMLKYo/v
RCOp5448m/tE+ki5kSijXb7b1+bUnDlClxg8bCQwxS6HXw1hr9ZozsQbOBKngLfn7Wfhd1WMTGlc
9DdGk9RyHYKNy6dBmQyMeXkrga6KXzZc3m+rQayJ7h4p8L4HmVlOqxvHhAlBnMPzPnAJ0kYoxAc0
WcEJK3klNagjAJ3x4arswIAs0qWB8oFXJja8r7b+pDY9sE191vaTK8dcdHGFwBd00612QPcW8v65
QQm/xonsIEM+l7aGBqq53xt+v+hp1V7X8v8YsL6R2IkUdCiZ0ZsCMJOLk0Ky714xIFOm5ZePuN8A
2FMucSFybA7c3m6R6Vcad92OWEqz5E5jKWFF/jfGhFlj/G9UdLN7MO2h8xG8QIarlJBEDPgg+xKQ
pp+RXD6luCp6J9EKO5Hpn0GXGlUBylsmlmnDlFea4gmT8GZsmJ7kRhD2hX6lDFeLD065wcYGQwSl
9biapR0tAf13pA7f9Wwq3G1iWljbQabwbW7adDxH6/h8Ds5nWgi+uzLHFLwpqAZ6whc0nttbBaKY
8N0MRW2yaM6iYDT7HUC9WCzWGHXp/SvGoyiZ4Y6IFYxMNX6urbqe1ja+9qzI5mkoMkRTbk5MNLZf
edazlFO58+PyaFigIA43NK0S/uy6B/iXhBoJmv4jylQgDbZtA1D5lxyCKUfJy9wc/gUcCFz9K0UY
rSc8mrXW2AAidtuf9/bma8nF6O/2ygtCYmCiAwN8S4jrvV0kkwAsOfixTY4x6efZd/cfwx0Q8NPl
n9kqKrJ3K9LLQVEeYaXOZaoqyPbDtliEHdZ5zP7uMp/9EpJMb6XcRNgXF1hDBhNVSlWXB7489ClR
14W2XJBIggdOSdIBrD6XTep7khb+SJSdmwD6nBSqovYzfamFuyqRIwE4QQ4I3LkPVJcIvvdUIgJ7
k3Ekuglv5Wu2sQVA2jw5g2+lziex+fL8+g8k4lZSn20P9ve188WeI+9z8q5h7OD/qt2RHaelB7X5
QBRiB/IMC0lsOzrMtx3NZVMD8FIKRG17b6EoKjWSZ3WgnbUc95iwjyYwHopCUprA2nQEfxkWWobq
acfdvAhwlGNFDsugfNUy3xs/tK4XAjJwoYPtFBBnOapizj5Ercz37p2RlzmCnZ5tDbIrmn9NXCM5
KVQjCelzjOqpxPWT4hSCA08KPZ1oD7HbcHlD1Eyxtz+UycCPvBf9OpxydBHxx7KqSSIrCHGfqQ7H
A9/mAaHFZARklvYkUgHmt46GLpX6RF0PSQe0m1XeI9U7c5A6X325urR8rx5SaUGyyYt29+ELbOy2
fgWK028vrHABbOO6m4B3UYhfADXRwXVMWPbQwl4lxj5Ue0RtY0uMpvP9vCCBiSzitz6TlzZdqntX
u1fK3AEISdXsnaN5rNA1vXE7athqCI43Fp7Bl5sMSLKsCNxGWOnuvJeMZNnVY5uRzW9t4v8sqGPf
4XNlRWmU7cvYqkK1o497tL4Owu0wMr5W3GzR3vjQUoBpF3nEBfJ3/hyK2cxHjCCasRk4qMom+Xce
0UALcLNDWSxySNymb+b8zXIfH6q4zjTaKZOfDNi3PYwTxqSZ6tLf+4X7bPNXXa+xmpX++CefJA9m
jrkJwl0shtQcyg2kHREi62ohYKo5v2xAdD3bYpgODjgxulXBoqKPg8qz3dtOjTso/LcRrtOK2q36
rt0hY/ObD5htKUuzH9UjP6p/FZkLz+W5aGqVUrbx4IimpO5bkOd1DVf4BlVq7YzVMPr2otoH4Eut
rIG1sytyblZWqalBBRb5hAco/UnGEBVSG5MVlEetwyQEETBh20acv9t6x73003PBl2uDp4DfvmC6
nWgR1kpnNPUJ2ixq9Fniq/V9ze6G7AaNnRSS4RkqvZKqR/IlELs89F1D3THioujDpU7y8v5JuVl/
SMNYKNnKC0X38uzBYdyFO91KzwXSC2ie3cO3ap1wHMyCUiOWN4/I+jnDWn3AW4E88ZcwIhIr8wuS
ZOEsMt+iaHT6DJbC01ehMULXDRRftbL1FrWoEYXonTaT6hbyppZLaJUSZKxpc01ds+rEYhENXVOT
0nYOBx2ob3PwYm1JeQkEQlQxjhm/Ton+MiYYSxLhXD7XA8B3wf11d2qa4snPXMry52oRgPYRx6lf
6o0bYS9/rDzYbNdhM0p+c4iR2rDTB62y/K3tNMiD/C5EuJsdhdJpzbJ6Ir6UZyZAGWAT8p5JIbpL
TNNrTSi4SRhXJniruxwg/+oHNP+Txe0wduwZv9Ej542Q2wSKglxKsHRu39aWiOyd9tbVbTjQdO2B
18FT6/34MUuvEUaA5ldsmR7zObgmEu3on1N7DRFIG0NIOumu43PdpVxac6Bs6rx70FPa1+/tzKOm
EronKrEywvJ4FOj1qKl3oRp1Gd78PodvHwgFTVpS/7YQ0H2AOMyzdaJ/PrEj8K37Q22C7Azv+Qgi
OnNstJDyEXqwoyoTtXCIvxBDt5ebo/rrdyG9mMEZH0PxfcTADKLe4PiWCsfELoBGkhvaBH1byG6q
garibDIv9gjVeU1Zhu4RbORASiwxLOM5KEV3iltkGvmT30xSSaTm1hhoFf1YNGBf3Ac0r/0Zg8fF
4lRTK7dXvjL4QqXvTvEaxkDVlCBL6LyMoZSahBUhYqcAA3sP8PtW2EMVgPCtYWSM8hHFGZj9UAUR
BdqcVTa2xJQc8yx9ai6oxR2aQKq0uvCmSX9HREGJXE2UJFJHqnQlr/4FsiCC+fAAX9bMe2iXuV2S
jrmpRD8KRrKGgFaQNQM0RmbM1329BWtNk2KDlYDVTUQCvPj4kUYbh4C0jk+FqPBpIvZ9xsWp6wo7
q2oDlVXZDwCHR/xNSMaNLeMy1lD99Mdpf1pe5f6Bf9s55WMrpniv2FBy+/fkm6UoE3WxywxjtSfM
b4SxrDF0pFo5Nn4znOdAT0fW3vzcb5xL1pm0zr7xHXOmwXZqI5Sa04rjkmE6TG2ccFzgRmV2DCPO
rVPq63HBOkvyNAcQjkuqr3rRF6GHVpv0N1ooLjHlPbzGwZKJlYdg3aLtXz1gN16fSR3aS/rhureW
k1P9HIlnUh8KRCQG2XR5TiqNGfDlUOWMDAIGQ93r3g3fm7fyYCLXCRWiA8pAFPpe0iSbEVUp6r2F
IfMRkrvq1nV64POsewKO+9Nbxu8GLp+01kmKXxb7a6lrh0+puCuKkN5FiWZk+s0mFJbvgc2yl7T+
ee3KX+w6s4Cb9QF7zF2QaVk33gGDUaLwL/+7TmX8lPu0U58/C2LoFI7dC0jCOz0wRfX+WOcn/NRk
alHyuNiD3ZxTJw1GyMtl0dwkUZNTEzEZsK9wDJpyJVLvq70g1C7ny1fj6qaLFenlQfTh10TqW9cL
Izxkb1NH6gwBUJiIbVbe1TUWBjSiQjDuAk8KiM1Q7QB3a80OtFobggWUk6c0W36eRiSZhZ8ftQmP
ystVU+ZZI721SYZMvtMQopGbIV177f8Yz0OeRTWLGHU/KU46bQljh2Aa/xftF8aOgEOkD28fhCrs
sw3OgXQ+Mexr03Ujzu4mkZXSG3hLH3o4851F75WIU1b3VTu+6rvHn6bgNlgv5VxBfMYP5jp2oKKV
L+wOhGr7MWDu7s9mASrCCCAQSrCtC4bsX2oqR6mi6w/BoLJUXql2tEE69YsKX3t+CoxmcD3o24QJ
hkFH1jI5VpazpBu9toZxmatIEbURnLKzwmItFDVfj/lB/uynN4UxrTFxzonn0I8MvurwqsS1Kv+f
mk7c8rnSqDL7o7LWUXnRfxjShFc1qUHwZBMuir1tg3GwR8ElxFP03Gi//QjNMPaCTzdptHOu+6u6
ZFAtLl8oRc+zTmw30yGzNJQngoYPRezF5m/eRWv79Vw6J/CM2ERqf6JuNYYcDC4jZfu70HdvZb45
ENPc11baJGD6kMWXjwPpEwhEtZb2/hOo2QehTKI6ToYyP4zSS12HdG1XoQBP6HQx/rRNvV7nHGYv
/V0vGB3gaon8pBoAgpRmOdM4ZNEpjGamaQqq+VS+9Wsff+fUaBzj7IWrl5DHIbJvhHp6R6nc9I7I
1HwX8N30H3AgMGwizqwiI2NHyOWPSxlWwwlWtJR5RrG6O0FJ4JNYCkXdOHXFVKfJIK8sZpmZcRB0
lEDamjt+/rMDGauBkh+WAeOlLrpo1r9kX+XUh+g3wluErz1YdFqW5VE3weMPu8cq74BIwi/f8U4T
t2ynmokXs5ggj2k571gqgeXHJoMffvanyf+gLUTeerWpLfVg8jUbh/xs5njCj91pAIlPEGWFTE9d
6Psk8QlSyXLny7A3r6OPc3xHvBT2eHFTsyTp/X90OuHcZznGkuepMsQzpUtPrP8YspoLJ3/wbo0f
8BDrCJTFut6K6zisBIe69kQVUqTgVrTy8m++joSx9ewxtrTZhGoXB/8X23oCHREC6OU+WMXRT519
C6tabdGHfxwvPGyPLd2j+2VWZ8P9Oe2UgyhHaudO6fDu6+zgSrBZIg769rpRqV+AjMjxKe4/Vv/U
rw2LIYB7ej129uyB3JP2o1/sDqcZUcnKgoQIXGj0fP1RJwpOMr7uVWBlwt2ZwFqbClgZXpTeY/g2
3kqZdXdwqhuGCY2q4uc8Y2JeI6n1phOrTe0ih93a2Uvc+gIHlg4KiFmvz8W2sFnYtYDcbKNCBVyZ
KkTwQJ1M5ppRWiOdYki4Ek/gZ9qbzhiVyw3iHNoUK+q0/h8SeYcvVGMHfC71l+7OauRBl3OeJDNC
I8NbL1O8ooXWVJiue7VsU5R3vu1R3DSuwWuDfIE9t/hoTXRRzhPkqWQ/WRZPn0sn7hCYoYwHpOes
DenmRmZoC7ogVzZb5X+uVKxrEseo40sSJaWKn3169c3sdFSkqxWewFAUAgei//+TiNKcB8LJH6aR
PBHNoeT7Y0Y2Q/PLTNZnaRJRhEeIjd+P3E5lT9TWYQH4WqJ6/E9DDZh1RG/MfAnEnaY5YQlgPZ7Y
pOr4UtZ5lO9a5S0rDQJYbuoexwKhheRuNj6YWwwr9D9+j3U4PVO9imaMNUhYPsJ6GQoMvtjO4fQJ
zCaPwenmSCqJj4zt8wyWUMsjUnOgMALWYITxq0IJInc86YN3We06iVECLMMwPraNhEDQEXtBN50l
hzg1hex0EtIXJE2zvanAiP/PFXdGt1Xu7ezWLPAfjwkONpbfziVmCgb0rqMP1PF7idq6McQ5Za01
SUlUmTsJrhyNp4k4JFOkqDAiGpMZ7ImfqB/xrWMENPiGMaaLE4eFOBqh6op1cpba02OMDYLcIysE
uZVeYTT1Q4J2YsHmJ0KROA6M2R7qjTok7DB2yqWiJeojrWslGyaH2/5DBIsKB4dlrsJnBYqE1ZtQ
yibsec/+KiZhS66fgZ8fRzgKsvjZhbzz6wC8yl0WADRBInv1Goscrg8YlkONx28q7TdyGYrIoovu
KLtqyL9shyyb4e3U6DF3kSWUKfQ6enRH3zolZbDWuKtf6gCPpHXQcoxttFtMkwWPvL4l+iOuF7x8
Yc5aOEVjNMNxnJ3R792tHrLl0G22X5ukVQsSCNKyq55YGi+Z3N/RuxyXn8wECKotfW8mltP01xAy
r5eHg0aEc9MegquGUa+m8P3dKAwlAhUpK4kA8r+24f1BH1hY+CdTu22N/gHeFL4ac1Qyxp46/pkp
qj4nPWBP9jDF7PWKgz+BAC5/WgGWfVgdnJcvAZ4ck6IcbWmH1aiJ7V57DbAJZavzn2h0HqPFV7BF
PO/Rz/ioaQwhjqFUbUEo57ZzfuTSKpfB8sxT157wG3WeZQ9F6a9bssxll52dk8fhBdzmMHAwZTr9
8OiYpt0uY2C+BnvhdK4/T4yRC+3wBgR5SZ9Hpt4Zbr0EOPWVsKNoCL9LJITjvqO7005TGA4iGCZc
w5op35ixXGqfwHlmrPyuaS5bqzQVA54X+QRKb9xjOGRTXaZkq93lXaozb9SycJwx6QVv51w572hc
ozFmP+pWslM5LQaZPin+/sUx6Fa2N8YnOTM2xdRPVChIKNVA51tqHl+2HhaZRESoFw57xVL0/NJM
vfTKmX0YBz0eoEohPI+9ZzOBLSbqf0Lz6VDStsCIZvndRxfPQAI23s7GxVlJu40o9ySyLE+i09xV
4ci9FE601lkvvbhkr0m1CQ7ped8qusRi4I5BJMAl3ky+Awr8j34uk3Fb4SpzUWPP2yozf2iZJJuu
D2+winZI/zdBI3H/dSeyufMOP6ZGzLPrRnk88yJion1A9blMpwUHYpYrSjaWB1yi5rsr3NoUndTw
L+HqJHbG8b02b15R6gC1zL5RCBuef2bCEbJQ2bRKR0vhh5KqnnlVrfQtfxlgjQMX9sNdRx0HmHiK
20tlFHT2FuoAn21fyblYnOJHWmzclRwwTytHfyvhyXP+yiO/wrVAOXhv0R4g0b+3AJNG0Stf/4Z0
3wPpiefvcGlUAgwKfiqmXBYlPpzU0yyJKTSE4S/3rWgaog+1cPjt6xR9/bfyGIJX3MCCTa8sVR1S
oMbx3sWpeEXn+F0BFyMhOuOy8pi1W4M0JuwoAtwabI/b+t0SN+nXRfnN9H6vQAePivP5POHWnTRC
ig+2gumtJsw3q9kHR6USaKnTV2Uy3MoHIB6TXtRVkX5Zx2oiCOL75Phc2NsQhVaC0VELm0QQMjHV
UTjYMbDbtPYmid1Kr8c0Fubr30CxVG8LpFAY/wFQ2iLfsnfArVA5zkIvyjYOkBHolaWNW2T2SOfE
5KXwyIti19RHGF5urkZhCan27kfWwu4gxUn62yxQ7YtqWYO8JfUnwwWLGBscY6AJyIEv0u1XSD4S
wqQv8GBMNzzPov/49FAfwde2lY/90EZlWeN/5NFQv0dQF/JkQWrVMJUax2CkiyAAbSaYcajhcV4o
VSdkFYmyG38NZHTyJOgfb4At2+9FBMqoQYuWHoZTKEyGMhgVn8gSGyZvG2c/VTkvHBhwkO1ai+C3
xx/ZQWwB4R3JoaPe8epXCB+eQaKDoz4e96dq1BMZQclDu68FPMkP7B+lJftyVUZ7jYA6oDoAGuI0
e9VaoU37xT+Grs8w88FrUN23S1zdEQZu27OhQLRYv/QZcUCZ/aIJneJqUmZ74JzZT+9T8UhvFWH4
Pk7PDjyvZP7ktSlEWKLZZVoz3ng95YxZy3HtYOoU5qsU0o8voTo9nCSjodRIGBO9wdwJSPViPqO0
OxJbafm08awMkikvBan2j+fDZMhIhaugk39RD0bBvWIgI4elxlVPNh6vNXs5VuDexkuqYnqRGmXn
PXtABbsei3mU6F8XxbqEL+CuqSy3EvKGaH/x8w7rCjgiwa19AtA6bvC2eYISmd8rGdd19jC9fjP6
wGpjF2x+wjWb9q5CBPb2aL86K9yye+7G/KHhgIySo5ejngN0VGlwazGvJpe3sH9RB4HnCF2nitQt
8w5TtN2rjpHNtG/DC+sfdy+sOTAQw4WtD9zowkXg3Z4WkyvR/VXgHdUxLVLr//DDDJKAGkwEYWWN
AJCYb1QFhk9KxwJlA0Cqp0rv2/zMkg2OpQLq9sxnZFy8t462+dsM8Y9KVwNaRqqz1C/zIyx6Wq1W
OEnobIvxUeiLpD3kHAQcU0ccDWk75vEzL6bKE4spn0Obt/x2blTlrebfn6ZLaUDA22e0I2Mxq0PT
ExZbjtDx3AwwljGc/E1bhS9vDouvSHJcpUNWGa91T05kfBufL5pVEcHGHWI32nkJo4q9QW/gAs8J
yDb2GtnpprL5d+7+SMxcwj9IR8k5l0qMjrY48JArL/dCxqqRHCQM/A9EaTDO5UZG2ZvJgtR0gONo
K9rzUBDOyMhkN+Qu40GebiGPdCpCAx1yHSeHfcWO8+JEjhVeyBxA9vSyjtIgcah/6bLMK92DXcsf
3Yarzon7tcidpvEz13x7uOchoKWpAkqzo2+/MWFbJDQBJmKibhFkNo/PYWxH/lR0npeEBxznF5lw
rnf1vJRi5E8vo+jubwKlEINjSwJlYqFRgW5zvQKRJ9DoV4im92PXZGOTCI0QlwbOUR6PCtRlPlOv
5E6NTLLP49z1vQM8gEEb7kBNT5g8Zw5gvp9djTb9yc6De4kKCDWxWmzLpuij7qQb23CVG58owJ41
683UHuAPX4/8NTEZ7L3cgL64cDzOrtwmeUmCbui6rqp4JQ2USMa+yzBeHXwId6UgtEPB4pQsJg2E
EKMz3oH9tgExNWI4ZEGgouInMOvmKJeZQumxZfrTJDdaX80H1eRr6wdALV5Huqndw7JzDmTIqXn6
TnepTroMyzFTd9EHPBpCOWqztwVUBcqO4hvrV6eLZFAliyHRpDunQKYhoo5VkJ090pLSQ28BZIy3
OPylQDelQ+p9ckj3vFgGb5lG0SI+SrK1bYUi0j3fRGoHtwzplcG6/yVfu5kmeE7tjJdlICes1Lau
bXvRm35vp/NOf42xPiLMHctsF4iXV4pKcwqNGXdJzEwG1hrE1gzGfnovF5ESdnaHE1F/YLdoyYSV
JOziKQxaY1hboc42UaF/pa4YV1vjzrul6hoUZRHQoT2mco/5inIK3Cml6npip2Al5oekiH8a2wo1
77qJtTT09hgQjQQv2qn9rOXu3qOT7Lpk2IneF4gw/kMatkgtoyTAsiMcdFpAFgAAJGWetVZnG+RI
Bv3pcA4FSZkMmMqGUijsnJoP06xmZ2ekrUYx3GMJAWAwfW4BqskS8y0VqACncKyZePvXjsqUM89Q
71ZJtGzkhBtH/PFimc/OtuUUAJnKMsqJDHHwN1cnj0j8ytHeu6ecP2hWy54rJBqcToK+XkSlqAUs
jhcNqPG4XXafksE5JlLLiRDedGWQa8huYEzP44jCxaE2Rv6kgvxR11f2oFWjrBrZUbQoYdLRWsej
WROGYFEhVw4n9gcDNHo5apYCgTBV6UxAuAUnTiJTuYPdZT2GTR5rllKcM9MRN4zsu4TsktbhO9pw
KjpVYhcUkFiuFqMmt8As+OmFG7twozIdbwa3oNIPWWvfupUvNnmpINxBtstpfVMZsLD7XW98Yg02
D2Us+O6ECzlh0MbBxxhEm9SQ2J5czE5WOHN9PowqIRfRAJALd2Cag2dt+8ZEhNdOP4nQG+sDauxJ
dTcZRxJg6LPoze6zhVbogrSArvEyU0ulZHSDtYLWrAFWMc12wE5BXeX3CzHfkJ6TYCFTgP5d6Y8W
3bvAr+8BOvDQutd9439movDm949zYci7Bm8L7MMM3TMGat45QjTDLV7cQ4jbgazqvhrbsBkgaG7j
3s4gKdf838INNv9Dmbbz0Ve54yztMYgyI4Y5SXPm6XlAZCxEDw4xGnrmlWmjVAPsmejLYs0ycLAE
WCCx6dix/BUl2X7QWIxhvh8zMbCMOBFxJVGqp+GoKh/XQOdAWCFVCNjTXNzkO4ytOZwr0F78pgsl
ZQ33no7TZq+Wh+rWOocbeqTzGZDPkH9Lh082jAGx++fm9VHcKN9MnSlyRD/J6V0BISOE/3ZvNbOz
U+P3HnC1IiJ7D/PVi5OFHtHRxXaOjDy9SYTDl0eG6gPjRMRPWt2ZVZqdGMfcqvoaGQJ60ef+J6D1
X69kt4llZfLirAfmr5CITF2AmWjAAFFKK48muEYlXlA7eQjq0mWve9h6nLslpgZoXK02h2ScrCXT
sdjKL4HGRGXJRY9YQQ8NgMTX7yK/cpqLQaEwummEMDrz/UNzkujZ/1flQ/49YB/stCnjbEJM5dJ/
mYvftj10kZewsmSKOsDOvcl4w9/ISz+YKJ+2qzXj+RdzQMd4XVCukua8VUV+IOibIlKpk4pYl4ry
2F1qKRaiyueNV0+qbPuYnCbQXCxETKxk36V+g8kDIe/D5pp5R08K4HI+oiknaEEHXmDF8grubmRV
0xmrI0xrXYcFIj9NjaagZJ/86i7ev22dasUCMz9vgihvvGh45vVhzLiKO+/ryUBiLoCfzzdv7Kkp
yxeX+frt2qsVL/GyLtY3j4ZqNdvmHSFsbbNTEfrPAyzhpMnrtumiRexqfmCRy70pkS8lkPtbKz+Y
OaQCn3/4ZjRr+StGx/lzrAIeuVF6dpbzjmuQrkoIqUi/hEylh6bjKSKDMd2miLGVsvtEHQz8F9YI
CI1OX3pjCpg8F4yykuO5uSSSYZ7S9sli5HF3mS2xkhY/aF1S/OreiREoI9ZvIe+OCJWHPO536lD7
wHtclmBOHKXR37VS6oFH3ynXvOTwQ/e6yZDISdBWgSImC8jWP36N6DrdIJaTiZKJigK8LS0xbYT5
/ayCDbcT0rI7JgUxJr6/PRltQ2LBHQyeJaST47wzEIuuQAjLmQbY9bGgTDRySsG43nqlqeTmAD/X
gJYWysqr/ikLwSRGrBCOpIPZT1DiPKFtkGfG0mPdCEr+wQ0kFeGM1BqmMrkPEV51PlHzyX9Bfzpz
7B8NqFkwskGD8m/J+H0oDY+IkesQry10dqT2nYaD8Co+SCX2sZfiSaOITLR1CTVf28jC0GjTh2BI
MGBgIsfvSlinkz+C8zYP/zuJvjAy6OJA60FL20B7orT0fKrNjPRmehr1jYi5Dd8SMKPWjONwFWsL
f65WQF8LkyulZo5tw2iAjLLb83FHSrRAIJFYqDHYpeFxtVm0Morgt4cQCqfRJv2/e4rleHtn62mU
0zXNZAwflFhLCpZY7exSYiRuREJoHpe2kCf2jEXfXy6E543zDFBMbUklrv69FunYWdoN2aSoIitP
yX8bXgQVuPG1hU1NT+QuJlNlpjgQXYxmAKDUzg5Wqrqoukw/j2vaU3QBmGyB+U5RLVG06sw8q/te
pYVsWlmyRHtOLYJ4/l0zW5Ur5kNkZTaWwtQP1r7CElf9h0/CrE0+wgzcTybcepGw9fQQScckq2i3
5ODHOOl2asSuBOztSirnhutIVjU38wh+pFJ6plqqPmEyutUmDTTgCxDzoSIIVPvQuv6cZP/YhJ1L
9WighXAU/NMihTJdpz/Vgo8hJGt8aUurjfNoAH6XDRzfwemI0GZAAfhOrSxJIipLpw0bUcBSoKSe
DEFMS9ZWL48ngfIJ/GeE0TRYwEaRKTOAoG8aKUErP8daqfvDhMhHU5Z97yRLGDoQ4ZTgB3qT3in6
//vgclunV7mZaLAYxJ8vnUOqwV5rZ4rwUdLgu9Vcu5ZbF9/f9Tv81E0SQXhqdL57K2MSCPMpMt6h
pSaWINCclwjFD6QEh43r1zJrl9t9y0xIemQXaPmnps6z6c7JLzIhNPY9E6lMARoyWHbXM10hL5sq
kd41a8RrsKyJYTe2BfT5bHnWL7sehV3FBaOv2ho+PISVHj6vExKr5VAYNnnZcO7KwkZfxUBWvAXs
08ZDeW7dmTYddNLVTirWxIwu42djlS7O1WVVY+xYOhdltn0JaUMaAeJfgY4IpmUTN1//dJcJBD4e
qMRLI8BKAe7aBhhGKBsPOAcT2RTPZcaUK/xZkDz+rBKF+LjvVQYcNVr0MTvIrj2wr0WsG2tP1bL5
GAVQFGTttON1ROLjttjI/ITjBZjPf+Fl7X6GaHxUHUv5XZrDAF3KIn1JxOxPbulSoKaVf60rdZAC
LJMoyXY0ti6AmlRtlg1tKq/9xmCC59hBX10eRM/R7kLLNj2HNwnBc3ryYaiSHDCtpOeEoV2nq/Js
5PDsnJ1w+HKqmmypvCJ5QeLfxbDLXeAe+GcS23BMSI9PDH4LLSfEdXv9F2ieMleZobizurUyGYOo
1/68y1Rum1fl9QiQu78b5uwwmWB+GZtAYyNHuok2szse1Hq1OC0UXf7743oCSrOql8hJQCMCJ++G
wGsPICpenPSqPJiupQxH7APVfvop0h3kfCnoHOY8yca9Ja+1N4To1I8cQAikJQE6SUt33WHhMoxt
HCk21/KAQXleOvpS+hDqsnylQnCONOpwUMGDCorGDb6PBurAbDDl+k0dRgwSiJCpoWC5PLo4ouA+
O2mPleuzrV/2jq5FtEKw8Bm9OiF9Oub2MNiR9tkY4nmAave4kjs32zMuEG4zz7TP8r1IqbFBJCR2
4TlnhM6vfaXZz+7u4Cvn/RVT9gKadhuUsa8fegq/5kLmQFyzFYXMehdnoSaifQUxOFa18XGZkXC5
U4aW0kbZIL0Ok6EX33boVDD/+0F1tSmekWxd8cqapBLk2u10R66z4DFTX+oiXgMmSYab2VW87LjW
vCVr3zzXf+EUdV/L/O/oT4eu6GSSzfP9AvUV+GsjO+I6uBQeYIo4N7yBTcrse6UJWnc1iyCDHSNS
1U4GvcARDkbzF81QeYPfE3SQR21HuAS4zHWnP6kdAHaMnP2uF+ntAimgIcYuPWKpdrwFHBqzpu3W
hHPj6oTLbJpi0IA6YfYlVZyi1Yi4xeHBFCioVNRnu+1tFPPn8dnRgytt+DU1rL3nIlkd0+4QvvaT
QzPEJOQvY5trM+qZIbUXw3jpWaTS9nKRl1tb884YZRa//ZIqe0C9BEGDhozmbvGzXf4E7dmStczV
9FmfwXzUWB7r7h1ZrlJuVzWJNu6jsKuKyxpsa75TGhRysWsVVZ/cVZV8tCWjMnYgZOeHYASQVKAO
xwiwRZC72yxkLuzcp/96CVu13m3Y8O+6CSeKqJ7zlkI7H9R4WPVG3+SeVfgnhnh46HInbumKcwXq
Zkz+LpPO5jK2f1UYd82I/wEp8xBq8PlEUXtsWIJi3dU8J7Vp07it/rlYczErodDxkO8c7w8K6nvW
LxLnjpUAT/Z6qZixjAYv2cZMevvpvC5pTLsyh2CiF/epKsoZ2v9H8cHBQ0C56hauvf4dCiSh0i2o
KGsTot1ITWlKoN1e4+/eqsrdXiETE701Q4eKs47KueKTqzH2EsSBgRrdMnVAmKFnThwIHPANyNXa
NlBG8bt9J5AQiHwV6C+j0LiiJwBuC+FHRk6xdAeCpnbLiLRp04yi34i7ywIU4NPBt6QPV+xe3HaL
ftUccyBU5KgjU1+6woRnm8FPWPnZoBAckU5vrSnGUAYOICloyjMglrZGgrF1DK74C6BkF6hAb8GN
Q40+8NDu/zwCcOFwHvjwa/oZIL2ObVw7VzfWvpc6D0HrGQ+3qh6fTKpKlYBJMrU4/BOt0yehONC1
CZr+27sWMC4SgsNQ04X3cj2XS0e274yTxdYSHi9CYYnucOxMg3OMWHGi+gT4RZ2jYyNDD0+K8Dek
metzWvtLdCkxjwdEqItjQX55wjDFXa7WI6gxjxUvazDGTFEUsq4v6LQ2UMk3rXwWP//zs7vlrCz6
8oaRAmgHoKKckKfKX+cYmoDJZy6PULI/HMIA5vFvKg6mGQpOJQvoZduow6RgPC+umt16h8+achfI
aQEMexUGCnyrrKUW2jm1c6TRY17B5IxPtnhVUh1OP25XNwRXqS6WoZsUo72kGrRIIfkhMjy0zJVU
OJANDRTJ4Da5KYdsMvcmmJPErmJsrlr9o8c76ZOs3DQNgUojQ/Vp+8lBHf2fxevDjYOBbKUn8+Yk
N16wyW/58piIC9Xi58tRFjMVyS+F0eXKFS7fnW3gUJ/bzE1iesNURrelbcPi/BZmNEjCnqBHTZ2G
fRaH/ne0fxzFqBmIobLl5HCebw7u5qf3m+wLQ6pqG/1EXnI28BBTpP684rRVy6IJ8Zv7rRsPtpVL
wD6MEWlSvhDe+FJeQm8zmgC/NFZamQa00ur29OI+BHpt6euEJFGCEz/1jsKNB13wyxdOo0FK1nc+
SPbQiLcmBx/t0k4i0GnzqnF7ZjrJ+tL5qQPvasz1oDT9TP19vbS57D9dlKXQ3jR0j+3W6YOyREHK
WH1fOVSsArobwgctR75SKaKBqAKYmxTore67RZqlrulSaHYzO0KZefZrJ4l0Swx7q+vtEaaqVzOA
QQXz6qhff8rHna+on1qtIACBlEIaFQUxM/F4+SxE6nOpyS0j4rMbmctMq6tz4BQ1erTUv9ImA05Z
XqiIpCtYeOH+ZRvp87itjYFYSAa8oDi+kAprE1u+kRTFW8wQ/aSp4lYQTTJlnix3u9TPNoIl5y5j
iZJHvM9wJOcGeQ3IwyNvibKKU6GZ66oe2YZu1l3gEOa7hp7G5MfwhFTmZLeeM102JVcgg8JroM0K
9bmvSxt8aWdFZtTBIhn6/7vK1JDgn+IP4CgGUk7Sc+/Sh+9KujTXk5MzZLfwxxUSbHewiQmNiA/g
emlllxVch3lJRMTJV1PHO0/Hz4o01ycr23HKwx0JhzP1JoYGklsqY02HerujMQ1LCf36cdQHVk1V
KQfmG8JXSnx+JiBqNY4fNIqeseCvWEn0KHQkzu3B7O/ahi1NBXfBaKkjX8KKJAimyGCy01fvHl1M
b8C4ULxxbp5BKcWeORPtI4EKYdmIY9ukIG7Cpt2wCp81SZXW+GGvvm34QCrFxReyJerPsjd24dW2
Vow+7xbh2tREtJarfcZxkNoDs8+84Gd3CZwzqyC3Kv5yOtLsXxH2HKhUdR6iv6wXJLBmvMRJHXiV
rPzMDzV17NgOdxg5WwQkyl4ZSBoFoYSe+8NhRBp5BNbVvfanB1lVHaXXfDz1znnQCcbSrwQ8lf1I
vQSTtrPPqz267i8yD0MZLfIenw3Dfx2zJum/KCqjJ1Z1s2CQwEiVWx59PBQzsUavL1/ikTDQ5edI
GUPxyoJg7VIXfRgVQTVhDoVXLE3SQPBCRnGg1wkHGMQbq2B/nqeK8HQWeEJTxnqKw/t6ixDsW+Hb
tF/vRT0W8E/oZjMNRd36x2NWPVS07oSRDIXnxDq4nz2JVIxjJ7rOZb1g4rMTmf6Sweq4XThaKGMI
OUj5q6B/BJ4bc3E0aowow6MD+QWWLFSb6SXXXVqn29/u5QcuUOuch6SUrGAYuaaATQKUAx7LV6Et
bdDwPjdGEcjjXUUvxhiDzr5CX37xEmSFrkEftUeywRsCrKpy8c7oUnvHPAwQAVowsjz40ZDm0XTc
hODmwX5hhlSWZFQloCgPI2w7UyWpcBQ6CY3lk/uyavhs5eNlvkAPHccg3O69VgYd8bQvOwkt8nxd
IskTlx3QQCFOCMiKwOB6XyOz75nQTQgwqYDgpvTO8NEVYfKwDN9pSHS8Ehtozap33n4QRWuFDpWF
v3gIqPyiXu03LTjrT3SVTlSeVWzlVs+8Iior/UCkVghyq+qQlpsRY0NIFZRx87Cq/hIMWONiuVdW
+PJNaNDX7s4EpiwoDWGdgKp2ejsrvuett9IKhTxWwkgDtclVkzGnPdYB5B87ndKD2AE/BjgowEvd
6rogLyXQGun0XYKA1RoewlRAWdoIeKHq34TwmDNN5tOaDQH2uMc21q+wwS2v5BiTN1OBryMxCvy6
IbztUatwXEv0s/unlwVmOKestuT8IZaI+fUtGiEUJWz/f+l2B6yjKDLlv0qyGEOgzonYD2LznolD
y9RsH14KkLLsCU31S48Q4ULCGO8kNHyvJ/XrzS9/ZmFOvn5bymxqgREZR8YEoW4yH9RezpaKcXu2
7mzXJdxwDBskCbskuciYGQHbaUvOZgPhc9yL+wvr1J/QBa/JKiAA08yLb675C1Sy4yYTi0T0nmL8
x8C5ZRl8i3E9KeysYvtNwBKosZ5p5xHb9dNBTwF1tOxTOS9XQUIig7Nv7W5AN6NSkmam3auObml/
n21L0AWxnNO5qArHMrOPPX7y+MMiyL83NJsAUh4O+c6AQ0y+To3KZh+IskqvFKCV5NGXbF8LO7KG
6MKgBHFt1J5tQovDg+lyK+5ptwChB3AC52lxsNtrRIRA3u0iQ/RPR6VTlnBqhXQhOuuiHuBQERNL
KgQ+AZ4p+ZkfFoSdgeSqamZoGmL8qypp9Z6oSc8X+uITVCsmLTgqd4HYe/pKwzC1Md3OkjsEO9Nu
caggO7LU1KuYez7b6Bxpluteqtuoce4XDhzcpWb0JldK/vHqmV37jfDNbZoPGBM0yfBiBEEzLr6W
kyEXww+El1aQs5ckCeS0NQB9Ep43rHDh13FMpRG82qgEAorV2lxVr7k1CsSxj1OTWZXA/b/vQZ3b
5S2vrpxGuIuq9phwr+jkgqJmaey6zlVKbmrZgW5ZmWWV+gxyjeW6aJGeguD6AsGxFb/MlDcPCo2h
1Y/MYyfckYlUKy2esJT2Ma02+eXC+q4dlYcdWqHm+LT8Y7L8tGXH9IrcmHwteT4E8FVi883D59Qw
lnWVvS7wsYutLDkASq4EHfKpLUZwfq2/HSq0nk9dXahW9A+gJDZcnDG/yDS3Gixuyk3c+WnQCl25
twMrpT4UjioQrJHEW3bp9V5Gc7xFPPYBUxvs1aa8BE//vfvrUEd7vyjwyBAvLNpkWkq7fLAClvwO
i+xNXx5KbKdXy6YZKHRD9hGw9ZsAb9vw1/xH5YLCVCpLtCTtENpdvPa0I1o9bEQqzVtSdVZHgAFW
vxGUupzgSy8DWqCHmkmMfLUHXsm5g4Lk9hNM/9vAj9ybhJdeA79cbF3hlfB64aPippETJa55zYCN
Vk565rrkPT5ttS7cRPpWbugzWLXedXM4e+q/TEjc0vpkYLDG0kQ0+WfRtXIeen4j+hVXZvNfipRg
yiDPPzwQ36kheWh9DFTJy71pVoLNnKMFuEqnDeGvXcK72p6DgFAT6IJKqbwVnqzEJUyCbvIMoa/Q
hOAv0TTPS2cgNRdBC9bADmPrJP3D5BEEV01qLPSzqRTA2NOmMeZUJdR/gDWXZfnOgpWHXc6R8QTD
UAlmEfGMNa+HT8TM+lHP3V43/GsapIB5OsZgqp8ynUxF1eeKp7ePjJXh8m5kty+ovYgFUWrUZTex
C1ih1T0M2SnX2512wOrf3mNOHiHDvlW045W/9cF7Yp14vZoZji8lS8X0ltqBO20XpU80zgR3tqg/
1yT72kiqtyVDjqplgqO51VuV1afMzp6CaNQCOnAPSQwJjQeNwo+aX6fsJL/NQCOiHgLvjRezGdi4
+MY1ezDXLFKz92r+io5DFyBcW0ObG3APToXhzIQ9yPksmP8nC34d391djspO4//498suVYs8KUjT
xgODtzG/fI68NASFVZn0G5y+vn9A0dUaMlz6HNlJD7o9x39rr3ZOpXqMnzpW1ig1PLCSaYk9LSu/
gSl+MTiXgPCLOgjljktPg6x9aL0l+Ju0lxJfkdxd407eqPaNvTJtEDzWFLoSm1we/07QIUEPw0A2
z+C+/rTRz4QZI8OIdiGXwGpABQwpZRLT3cmJVTAJqz/4eubd6LLVBkz9Ew6xv7sD2WMKXDhSlPyd
DMes17vFROfelS1VafGCioupnWYO3nhR1ezuIVoQxplLNIMjnC+aeWDz+PVE5CRgA72GtaP8uIOP
zRdUVfX5QJ34J6oPVwFMIOH4687BvLtO7vu882sMZqRBqQRmGoab0xywQQjQdZjlnhTChgrxUILj
97C2riPqrLhQm3NUC0pl9HthtOxWP4LrvLCV5F0TslST5DD4DC1w0VdQo9tLea1Xrf2qapMGr6Vv
7cHFAq9X+51mYyJ19NL+v5BUxEuLl5qNRiK2++n1Wfs6C++/so1sgFo5liVz/wsT5gfmrbzNJXf7
NlscXB9dQdkZxsxUGqjjkEm6BAYQWWamkvxh5tdBP8S3+FoSenkMjmp+qI/5sAh1y3BeemGdkXK5
vpS3WkFeTu8td38qn1e8vciRuNPEj1qxElcHcU4D+juhbRfr9+3TDmqnd2OvIOnMTwShUbb55e9s
iuyIoCQ+tTvoy9IyZ3RjqyFqZmop2gpyrsOmQ7TAs54+YLpyvMgZFAeUO9qb4j2Gb54OHWdaV7uT
9Qufl8dy7Ia1uwCAnHvXtxJtTuhsdtxMZ3MpoQCs9YI0Td+cWkPYHztWI8x+6v+j0lgQKDOk4Gvc
holpez5iip9m+rCexpuOl1mGaJv9xoR6LxeNeDxQ1ucW+puDPZ/O9vV/+ZRF6V6mKD/VzPt2JxnZ
o0e4z13JOxC7q21dme/7PkIYb1TtaC02SenV8k8oeyp29yL8psqIngVmE9oppVjWoFnmij0f7myM
7N06/V7n1eqLYLuDGd95JgmSDlvT1KL4gKSKqZ0DhH6TdT8w8WdkRsYzosjdn82IZuZQAU0TNlmJ
TO5lZPY81R8a632M4gSue7TrQMBx0tuS/UwUgt5CnJsGiU4bFYeSrHfF8TuGeosDW6KGzXGTZ+GL
4Yi08R0mX7PeNnq8UfX5Jf1/OCc2gbFMc6kElp3TabcRgEU40gWQNTX2HrEHKpFOtWBE0LETp/Pp
vlV5lcoWoeIoC4EKGX5GFigY3gFY8+nsZ9iE9jMNv2vD5hqFGWk+sKMqcwCCm1tLZJjiqbS95jmZ
j+jCmyUefoOj4naZo/eWYzAFGcz8kYA5ackrJDEct6/+AeEu0ERasVdTCC62Ntz+L8MokyN+ZrWx
rBPD8CA0hGXwDfvu2vzu7Oj35WfQ+Y99I2WUQ98y28VYaEce68Do77milhs/XPv3Q9Rx5YxD2Hxb
uPDUpnoMovUdftwOtUcdwhPryEx/ayPrZ3wSNSO6DTEYwwxux2I1QsD07BSDbvkInPuYrQWFpba4
iBuqLGN7H+CyEiMp5JA8/Y8T7wFSvMtRlBsOcZHGP4zCObzw0FjYmiQgLguPZmEk02yiKrUmndsj
qQo+emTKK1BKKeSfFpIXPtCzw+q9TIAD0+JxxbAyzMZaPdyhpZCdfuS+WJuCThd2yh39zUVztGDa
kpGEHFHdp0z3/Gh+xK4mWaLZLCs5Qs9DIKC1e4Wqb95DRjU2L1ZYZLd0V/T2YVPnlABOrRIRWK+o
SO3dye+OcE2mzhocFXeQN0vbHpcGC9KSwo689mJNaylGThgzCQ2Qb3LxWqyBXjpt0G4MG9HlXQgC
IilXZMfj4mz4pJscLqj4UUG5kTvOW/XbS2G8iu2wHsh3oXWRJaWP2SuypJBqPq0gZvJARhzs0E+X
/VN0Cg9pMPMGGHvDjtXK1hgRSbQeYfhETGn8OIDtvIA8CDXo5j/hwuOhaBsFD6JNoztD6Yv85To0
3SPRrqU6UntpA8FjdDEMhuECK3JZok/xOFMwq5P7bKaQSfzNkh2Y8HrXPsD56Ta7r2WwRsR6Z8Ox
dlefcyAskwVCoD04igH5AKsncdM7rpYjjmg5ouqVSJcqTo85zKbHnNuMFfBCIjZUlzzNvVhynY73
ES+PHisiLftAhjtPk9EyqHtiW3U5wSXFd9NhjOIRcHBdjq5WxsoL4gSyXwlw6jzxQP0K5NkdXOAp
Vq37KlpZv0PgOikJzufRORAKnkss8a50z2Sb1ZbmcghfD1GBbAazvQEIP+vMAX0xjRkco/FYi17J
NQQFaPvPNwbwQ48b1nGBJaiUCE6eXYsFa9M0Pi0wY6EjxuCrBE54A5tHqc+w7km3pFfEfG9yKT+w
1PmxrlmgoiGc3CUhID1c+LhqxFefBQFb4JfHcwgKg8m1iT1RCb9A/vmW6WkdpJVQgfMhqUIHA6US
Dp6hw7Eru+Xpop+sZdT23jYUYn/3r+xNODog6EBE0EmLVv6dKt5XO65abEP0aO26AJiWSX/+L9C2
3CO96p0yEB4TGmO4eouvm355p2vlJcXln1I1+Wkfmvqcxs9p7RHTCVNcGRTvh8k+bmJdhc1qKNkf
vSWua4zRFXNz63EIy/lojvvFLgWZa25dTApNW7IbQdpgDzMw5X3jsYEpkDpy7z1xMMEWN8YqkSIy
humT89olamMHWqH4zPq8Xv1PkdopkFK6xfXBJEfeExdnlGf5Wv96y8ltWQHATh/wdfF+ZrDAdaco
gNtNHNJJcgTBwGOLFq2T3uSoao3e8QQphJIDtmr7f2DDObFfr/ZIQhV4Lvwrbd4Lj9oDy42Uf2md
ndwlQOSKbfQeEckJrdW9PtlAoS1obMuGQvxQBnTDPEXJYGsv1fiIympqpMSqjNK7yK9Y9o5s3f74
rSj4qzFOng266xl9yf0udGxUctzwFDbj5lw+bokNXyuB+O9Rp4/rchl+oICSaUlayFooLSavaLtt
9H7+/Koag5QzoPZc+NKuCvKNarMRKXb1exSz04zmZAu8bjbKmKTlnLNDYCNJ3BqH6jbQ9j8XOWcA
/MhOScc65SZ8TsXBsee+NtMl8KeyFodbwe+KahnLcATqpL60bAZN5wzcZHpfxpc+oiEXB9aXRd0e
xyUj1jdnejEYU1w0BzD7MhlDgZlo5qF+hMFPjH3tsf4E2Xc4IDIS6AsFLLX4OCN8YzEa/tx/RhQI
PBwA9x0QzaKHwNdFcvzd6gGi+gPA1gnp65TOl8tpVS/t0wBwf7EzpFHDAB90UIVOxs0GIJfDLz6T
+Dr00Yp+791mmENOjBw4qy+xf8rcw/CQYg5+m7Ef7PAlkAfAenhcQ2aOtHG3H/0gkr6Jl1SxJ9We
eIfyuvV2yKGQeEVPjtCzxsT91s8uyiNud6fG7jgty65MBUkIL9qwR2M7wsx2LPaNvhZ1yfPG64Fo
ZQEW0YNZRW/gTK2n5rXAkUwCe+iCW95v/JDs9hXr62WVk/cRhTzAK8Rk/FgNMA3PzrO9KATyfkj0
OTDBcQVvYSqmZhtPYrS4vSstIver69egzQVTaPyntbWE+UA4sdbEPNB1M83SjpOR9W0mR6xlS2gx
oU+ZHj5CgY9a/DL2LLOL9Ek8jykM8Ez5bs+9sRa9BlGlIy4Y9Y3HuVPLQJvzIyJK2tSpLfat9CUJ
/CMypTG/1dG5TImFznFEme1Zfnef7t3j3lXZ6J7RgKBJEcDbgbGINaVucKMXYbXFY+U7PELBiAby
vTSoFv7PnZWVP1liEPug9RQa/oxlBnJGjdcQWq1ES0r7OnCo41iS6rUqzu2ihkuQmVcf6xQd1shr
qw/yHAam4Jmkv36aiWUrJd7jIL65UIYQk2ktd3zk9aSilPaf/uE0ugH4CJnZdJ8lK6T6+czvQvoo
Y/jIFjUK7Qyi3RBeZ1nEMRAJ/5kpNl8zv4ZEsNfJOT4h1hVs4DUI+BiHbXAVVz8HgW2bb464sYZr
zB/Vm0ejbDAqx1QQVtWDVr761bhhfNRWj+GGgv4fLkPFwYqxgPM6qK9cZtgg0YbPW3jy/xku3ySY
FeTr+ryqqqnxhna4SNI6EnCUkLWorDVWr6o3o6mq6FZQnwVo9B3J2xyfutV5jqCwFQCp9vH+kpZ0
ysni/AywbrIJCiFUJKzpjgDCrcUcIjXTpQDtmiDDaFvHUK5GPUMfi2i3HkVf9mXghXuql72gbnuZ
/VSmzxLTdAJcdRwl+edtxAP6D9mmC4RzePvxyGRHSE3B3oDZ5LCfRTh6HNgcZ6CaG+4zBpF+Rxgx
2zf9gJ/5kGZNkgqZgzdXjSrLEz76aDilY39SRrgZYbegH4kHbAXVRLGEJPRyMoAcKP7w8JCxlpkY
FwcQ9lKKVR3DkYzAGgBVBtjhNK7O1FEvTidlO3PHLWnpQsfcKv/mllpkS7LEK4WwuwF2SALND3AB
8vfIhJ7+0IB3+5rAzuiedsw05FEUgllCEQbl1wE7ab5gXFwxjZJrmrqCaHS6+I6QPHXAKbwkG1+6
T5aqtZNqvTn0ju1hAPSpuEBwurb3JhMoPWCTlLHspRl0fFPpHpph7mftCKNVnFtxoiGFumadtW43
aHpVwdq12tr89T/Hr3KS8m62aw/L/JMIr1DUR6zpZ4Y5eZ0jmDSzHKouu+qZkxX3auvDhbYyWre+
FjSugGp5+T7IvZY1R9K4DlE9fb4WzrcXCxeyEYtO/X4tWymFzgIcF6v/eKbXuxbO9d9+Tf+/ojGm
TTzcnpDP78hUxF5b5gJ6ulwzCZY0ky7bO2o4gNGeLYwRz0UymnC3+hVMNQsUyS6PpN8/FfMWMLTB
equpkiohz9rZ5EOC18Sn4czweapmcB1RuTtb5ThRWat59Cx62K7SVoyeE9qa0zE7U+fXBAuSUE8n
lQWMahqZ1qjudoA/w1XChJbdEbtL6Z74oOgv/WinwFJujMm2YaPVmkI8k5UbJj/IwgYLrbo6hoY2
svLEC71gPaguvIRy2SWYG7Hb4L0c51XcbxybCsjzLV3bTXOdRoBkZbYcxgja1VxUr3KWdX+5NpIg
I65LQch0nkog6JS+JDIIUXwvvr+VGaCJ9cKqQMAnctL9sA2IkcJOxhVd3pjGjZfSX3mOf4NqmIs2
/AP/Qx/oFXou5TkZyOVoWNDCUr/cxdMqqP+ANL885fyRtZ1eIxf3MsVVEqQLOIg/cMSeJhfijDWt
Wjvj6EXjWTK6GjbhajPH3jIBR79pB6Eja8z4YIIOCQ+zMwNQDXikCkdSDvjtx/oL0LE1tN/svW8t
nwuo9WiXMFqaKSknQtmVOBKET296bqB4O03gyi3Q+Qek95Ek0Q74bmzHpxWIpffm396+wLIvDHql
DfE75JJbNYUy0ceWMWCZdEsjnTMcymcdSDm6gmmnXumzpKVw4Mqe6hBOBkSyWKOWP3MX52DybG94
19o1NNo6WghVdSy7oLAx7lkOIq0oVHDLeoasNfAWlGflfItjXhEl+7v8YHN+y6vrBbappVT4/8kf
zDsWIlmIUPQsH1+NhhDXOchlC2vefJ1OONGU/AcDm9Q50jdOSY23po8MLTlJHSzfdrVeh7Tu4FFY
/wB1Ud419G0GoDkMpseYBY7Of6b6A5U+JY3Oe1jaFw7BRVtK/eMDN4HkPZ5FGlBXhkVi1g18ESFc
j0pGdFCF8Fu8/yQmamOKKORoAx00RJC1dTa3si3SQBar/jyPFO2xD3ujtpOAtuF7ymPVGiliFHEM
AIAnM0LrC2pn6/vthyQOEBO7P8Ps0FQuc27bgzVEc69Fm1veicldXzdVW7XMAs8M0BjeI7slkuXk
ewhSxKmIr1S/iL4hFM1oTzfiOKG0vy7O4JPq4WPjUUw6DGxfWvjY4XrokV1H7mBEY71raTck0Z+0
rULR430DII8kulTOh9bhRrtfCPxVhBRK8R03DCxN6dVbTCeE1LOnC3HDpmoYFYpegGoulCWSF55/
cvT68LtVrXtdQCB2XJ5AROdZCZa2vbpPRDP4+2/zL6C4WVIoKUiViWp6CoPo7jnJ9eAn8U6FyHhQ
uErgs36Pb2LnDnxuOWstvWa47Vuhu9s0BUAVEj0h7Mgsvf/LRcBYU+Zd8egHCH+x239KHswO3jGQ
oZcO0g7Gfr9+p2kGIZGsAIppu8rVWqah1gmhsE0R6yxANRjEvwdlkSw8GAQXcaSHvjz3eiUNfbfL
COzEYu05TKP+WFZA5OoLvwdt0Qb5ZOtl0nA+K8oZTNMcC52dnsdOhtXNc41JtNyWvTtcRV9oEzxU
+P9qCde5YB3Pn9X1yQXV8WWQgfQ0f8ioqpapNjBw5EA9awQ4jc/k3TsMFdVTRaONxpWQKZXbxDce
gi/RQtXS1tE4i8vqWxUc1i6rLk+hjLC4NgIMTC08UExejaJspiI8TJiycHEEzw3Lx35NtODF/Oc6
UGp9QtoN42oO5u4V/9rq1FzOR4Z4kpyXaxvAckNJKE1Mx39T4ZJ9WtFzmpZoLOEgy43PT8oM4q20
emPNl/Wei7/M4k+3SfXWmYEYIEmXDH7YQhqNUycTheZHF18MuUpNYUIRA6dyWBzove6fOiEgMJHT
h5R3WwM+kIw3PA+7uN8NzwmiN0vUcmydgq/TFyNnDjGwJbHq4QAaFfbjW81o97Dt9KyFgrPzz8eh
M+q7dh+7p/wXVeUOn1lf+YWWfHMBycpN8MYri5SGyRtmgH1f9X2qMSU6fCUayXr9g+ZsLLVGK4d9
KBvKt+LG9szhHKupQ6DcW85UsCTm3iLgArdsclLH4LgtbGkFJEVQ1QzxFz3RdwusRbw7Uygr8Vpn
Y7WtaVRCdrj6+xIOVAD6vemuM9JAMxrbQ6TtG5ObM9RqSohn51n4eWOxBk4Fw0EnM/BQfhImZ/BD
RZnJDXol/EvjJxKWnATBbt86WFoqxbN5vhgcG5byqIhSxaqEUBLFFg++H/R+K+f7OZQ6hcwGEZO2
j9RKxB7+4UNaEebbT3UYi0XNSbG5j8xGZDokLn/PcI4ViS1nAVBzySpQ7x4XwMuqZLNkATtIyZJ4
bNUoEFAm3r6lx99Ru6JNYrUpCCWKAILHDm4SWvQ1Nc2ycy1EYn3507zzC2P0X42TuPR86ThpD8MI
QlYYDSKBZGCQFSqBCrFUYH77RZMcQrj/0lxsGoDSGleETZhfQiHYJssZoIPorELjnUWFjD+Sl6Co
9IfUeoQ/yDiX1P5HgiKJ1oOCDh8UWDULGeqFGdRzWi2LevL1BkMDFVqKRV/rL/othfKgWqeozm9B
NHPrthgBKsOTB1yQjZOKz4zYJtMm4GynorbMMAo0XOoqfmC9lV7hV/5kcjqKA8AQ3Rhojvku7/fp
1xwTfPtroFvv+BjWQnCdzvrgYve/9a7LxO9xtG0t6CVeiFhtTGdkHjwwd6fpfPKiIU88d2r5Plg5
C842WELmadMHbgpRpqGuGpYU95M0B6LyYbqw/h1Pw0r7BK4r0nR5dnAREemGvxa2+uRRDCpZhni4
Fm7KumtS0qNnDjNVYQu2rVbIkK+LYFa19dezSDO0CCYXyZPW9x3UfdMG0dCllBGkA5VGjinYzA4x
pA5y3AzPMyXH3KFJ+3S0SnMPHcLIMJ1qSWuxj6sFSC/G5tmPob0Schi+gTOOKcXiSmSt0ake2ouJ
qYjWTJfBXWEXA8mD6OHWzc9TXxY5CPxWBnr2ldr3E+i804FtEnU52RSiUY5t5ScYhXYoRYbSvMtA
Saf/v2/go7Jl+6Yo0nJGsEV2B0d5dOhK2QsDhaqCaaVpyCdCoCGLcT9/lIiqVFrALTyAfJ9Z1ukl
0qLOA8F+uqsG5yb2IiHBHct8rm16+u1s77qPJUK9tdsdEnmcFTXIbxJ+66SX+G2qZ6ohoVIDCz4B
0Rw00XyfrIOX1tkk5n0wJNFg7Hx9LTXl5cp6RJe8azomQmlVH22xtdXTXIhohdMd6lfsveKrFfSb
Dn1nxMlQmF3aaHmJ3dogRHFOLjeK0Xq3GPetMjhTYbQAfy9C/7rFwtt2z+T1VK8KVHm5bPUKc+b9
OH08gRCHWGklnjzSL/shf87SJJiLLJUsrRsF8tECuSPTiVdLC5/f4iwx6TEP3jtFxqaCdZa6u8uZ
6IkuKMx8u/obO+H7ULHUXHglosQNIoDKOeXFMEAmnvQLUYRuSQcA69rqoQFyiCv2Or0VwNwTgdfD
nPba3ntmfonTfOaJuAE0YvudZmlp5Bsp6qWvynsIyxEIswlPf+p+3XOtIcMCmnqJPDcMd6bMBTz4
+woYD039+tukgdX3cSz9jcmtuWkvqkrgODTkFbpF6nc2x1SEGcMjXZW0skgeP2y9w3MVSmzn3uzO
gYHskfFZ8MVAHOlRYJVJfuq/5mDybP7rRgqgwNdrCnZRdMYFeVviEUK9jCGiGnWRwwASIllU5XsN
p9ayzF0aKuHQG9uxQSzVvlxm3hlw52ztUMHokQ7mQOex0RvOYcQ4xqWP5lLBjdvtjsbH5qaZCw3Q
s8fFNdRgHa1xNOhJduGgNuxnZ0YBq6BVa639dMf/t4pK3hKb0GvjwVx46egHvjugq1+dIfxn8ett
s17GJvYRxqbcZw/qgrLy2eYn5IZW2Nilp5rpXZAFVjiNLhwS4X7PqDoGB6KtV/KCZfSS1vsKwb4x
XCdUfFyNXKEtSB9KJAAv6Z0gctVJxtG+EW2nVAfgHsrbiGNZ5tpvpnG9ONqQdFtq5FdLIFNceHty
C3wYoMJ/8KRofmZgmmyVDSF74EpEp4SkMMG4H2QC1NUebeUufcXduYZZUtXDCSw4RZ+6lDQgqcwv
pImQElK29vNo4s7wO268GyGb/KyTxwyvks0rf12LT0poFJi8T+u3ptB0pAO5RUIzDhpV0hkxfy1j
kFOKJSWD88hnqHkOW8qKYuW/Mjw9b7YBhzfpRd69n/3jbD194w+jKri7Q47W31DanTfXfw5lN9eJ
S5qn+8TlPP6XmstyTE2FjyHO1FO4QsqmA7w9JA8P1QcR8r1K94X3gsemWzg7w1rBEbEvBnbAFH+h
9+53VOGeWKU632UAm6ubeDcNQJrfKaZ2xudDZtSYg0V4hc5K+wEnJ2zrP6xqqZP99AVh7XiRu4f0
g6pSxK/peGpaC/c2LG2yCBEM4yZLB4LTEoSQNgXo6yrI3F08xEo2sQHQsr/PU2c6fSNnlhx/Y21u
6P4s5EK+lc9c3AzE3ZwC8MguXGbP8NXMbWDorI0IPss9iXcNPf1/hJSiyRXZ4f4qMxZSnI3C9l5l
6+EwcRmfZE3V6GMriFLCCWgF+4MOi2oL9B4IpJpuOYa2YqqxyPcTmyPo/gK3O/wqxZb1DFF8Kl3y
MGCoxfHM8uhvp7omYD1wKK91JyyRSRVdnn8l7DCkzv6CLaZw0hZpYLHppPLuIJi5qwXUAlRflkeL
PacQCXdJUwkKR18V6UjTPHIZl0G82AGjksjPUSVFXZpIARI4c391Dyto3LS27TAdI22bKktf1kf6
en6wRzbCFb9YvutRClacqhII9FwItVDARi+IwNZYpvDAzzEOe9lpEgLSnPudI87200LKDVPTg91n
dGI8AB0xBv4PjZXNDpOs05+812fex4U0hTibfgNMvq+fvFyRAAJHtgHKz1EXdB3DYiTFJQRn5q9d
TP0GU7cUuvbG0HVY0bKMCmfGAHL04uTvkYU5xEopEL1p9HbbprQnuc479ZoVN6wF27thBok/CJKE
GnKYDX0jyBWnpIwrPiQx59uyhnrI0MUxEhX4hUj1AsyFa4QLTlC/wl6Wx6IAM8zdEkUx7O5t9vlI
IUGLVV9Wo9pm6Djc8Yf/cIh/oEtLc8j3ByqUeockU8sRSTvRDb5NuMfVlLy5byEBVOiw9DMfPiY6
jtNqHilCi6vp4WhWA6nPqrkG2WiVew29UdSkojnv4JQRJSK0hOHX106RsbD4tZdZc/yd/TjGyBwl
87lgwgi/911J1+j56qeg/sr+HmiiMnndIlrgUhToXV+S7a5sjVNbM4x8FGyrUKIaKDgwuAxYBd8W
I5NGPiKbBoQv7yRU92YLFYjwtk6vlWq4wzIL2f/yTjp8XzXDQ5tRgkuMmikGDoQpVtB5t61b2XgU
duYZb0WkAKFJ3VQSakaV6CQfYU0GG7uTIlxNbgzzu3cJ5tIFDv2zbm3gHU/4j7+rKnKp67Xz3Djg
RW1P6GqT1UqNcfkCC+iXvFz4QcYLXedpzAJJUzcHX9rZHqR/mFCQ5ekpAJau54mnul+lhP3UEiTh
X9Raw0Wf5luseLOZJ+nUFaTsZsURK6PGNymFqYYCkh+gQr5ZRbnZxIQiPR19HDusw0322idHcFiT
M0O7xxBiIRnzkICNEVlfrkodI/sYir1HQwxJYwCxP3cYh+9srF3dhVywHTzhmC/YtI5NN6m6BnEK
qNRzocbjmqfyVWqDp6EqdeLgUjTtC/o27fPy28o9LLTP0JvQYbcHainBD+rFWvERxXdGPaa8NPBR
m3WeBn4WLAKwE5Ba8lkL+GamFOpWwdLE62/RInKTUrsjweHku2OpO3PVeN5e5+v6mt4/r90Nz3Jx
CnQ0cn1/MaI6rxTuaafD/UxU78R+pLT1MsCe4ZQq+ZMo2JVlyabULb5dRYQRZ+PynX4dj1JzVOr9
OT7o46E8Mp/IJcqzysMjluD5M8UJUBcR1W3+Rflm6/JZ2yHplAvnS2n1St2hVa1mkUcsXqtD7bCY
1tyhbwyQ9awbdbXskPfeAo0f8t5qqNrI1p3jT2OKjni9VgBuwTuyjgSKA9WziHzNBHRs5iKIkLIW
WFx+GbiTuoeJghS11MJEc4tbT6PinqXuEFcCqTBorLxwFjf40K1iq+Tu4IBoE2BsZ6uCaxTJdIou
5KVGwD1L0N47ny93CKVo0Z61m0AMvMTQIxKZK8lLDFMQxjncDn21qmSHoE0ViGTY13/D5sbXAfhB
YWUr+cqEafuTy4t+gjbpiX6kMTirkKFxVMdy8uavn7sxZJXlQRBa8/pWaMGwtGl2nWF7aMZRC25R
3QJwtSfBTLv4uH3xEr6npFwbk8SfL356UUH2zWzd7MF/s6kb0WkUhOzkSH9wKzLiSBYFI5kZSMCP
vktYzFdE9SQrhDl3960+FBwSKv56pb96WcBqeEYczZMYJvTIQZ9uu4gft+APy8lhbxH8P4w/Dq+O
/Mvi0dsNxmAHYjtkxaiikZh6zGBkzF+9DTGbo7ks1MJmRdd/WL/gmZOOiHAaVYk79hYSqTYxUcex
OKx9+0a9lL92rpTd+maj9xBEtPRZo82r8ZnbLDdC8CTeG+CM+DERjPvBba04K6VoO0m+fYpIeTMD
GMyN8XdKb8ZCLnG72mPHab4NhykL9xCruUrziklfYCQqw+tiZ8I+VQYZDKF/+kypY9uC1+9HdeS6
/ypSPARCLTtfcTWqggW3Eq7zfxHurOWm+TqSXl1GpGIX4v+aXtU0+2ZohAOPP1dpE1IsHeJQXjAL
WcI9wT9yjXAE2srMyq3OprDG8+H6MpXruqplEJ1KpIHRL+jVx4iMg71B3N8olIra282LTkicgPkw
/Hk5g1+z/DSm2xUNYlEJ2y+uYnviafrM0BF+Z1QEmGelvuKTUKedTnGq7Vs9oFhS6Xh3brr/5ulr
7Q/nt092TfLyxnJL0hbxOLi/FWel0BRozqU9oQNnjQ3kALEY3ow2Dh3Jkv/vBSmemteZ9hY4aKy5
nFpEHOquYIXXNY+OAgpIneS+D9CzTZ/w0sZ4GBqHOAD4LCuXvzfeeMWM1vhAMJ5PyB0NDHzRIQaM
YknB5E2eN7+C0YhSrX7dll7zJ2lUiXge14IKcYVY0K50Cc3DywU6KYozzOZzLEO7U2+Y/Y7beHaR
fqQ6KxCbQhRw/JzT3mMdq0UhemLtvTHGr6j8emephn1V5ES5fPTgm71u69Fbt0P/58ViDxWPOm2n
v61cKc+BBe1CPngHNBxT+th19B6EgAJTP9AluENB5eEROgv38TBEo12MfGe1Bv6e4RqDLRVKt0Xz
QoYD8XT+91J8QQYpvOO+V/fkpxMlSmjVccxMTn4Gid73J0qX7ySHYm0AV4UgkiLWv1nBzCA02cmJ
QPqiz8kLJ+BRcRq8KJWH+Gm7+SevetIrTlEy+QdaNv+8eizHP4iFQrk7umqxuJZI3iwvpAar76zZ
bIu/l+I48RovKRNjFyc4hClBda1jOBiVR5W4EEl5H5rfK/h5IXTwsBNJRe/OTBPva0JG1Nj3+SBZ
EPJHcbm+xTmt1tLGtzsIN1utoBfMDRfwjK43NagtxCl+mDrw/TGrLZ+rVFkCkoCvu7qhZEZs2CG0
/GLtvgtZ9ZvW9s7zLxWEeQZD9RCG2PnEjfZKAceoK0u1qM7BA+T+cwLTON+tBzrCUiRSYgKmVwFv
HFM1LnDvo56le5PJ7sS/Q2UPROBgYWPEFJWSeyyoqoCBfzc9KYdeLj/VzvgRBxEWggFS1EnaZRIx
oAyzDRNlrM6pLnEJOmsfJUvNxYvdvxV+lnw5PVfW7LOt9bzOuUAUPT+YVf+ojC4lNpOWaK8J6Zi6
wX6bLCNPANrBQDfW4m35YDXrsfzuQkOVLcoUlPynhyw3akKKOO4SYmD8BzDxWpO1M77l6wuRQbi8
tEWoI79pjctnrMM0UjAC4EPON7S2S3JtroSM+I7A9bJvpC1hfaVXtQDy0M+FLJ9JcXNWOFsYthaa
LMZASa44EQBvCeNP5FyszXhRaeHPvn6CWc/JnL+B8Ubh8/ZfoM5OrOgFREXPzvl7GDs4arNqx/Na
Ole+CL4uKGHQvu6IdYyvem9i2Kl1yfm9okcAhWihJ6PgydOseOi+qyQZpGJaNES/Oqk8JuZgNk6y
gE/k9wabfyA46yNBq8b264PTTQw7QlY3Z6+jokh2ekxgxfkW3TPVMoDPrPQd/EcAZRaVKF7lyaVW
T+1TLKs4VxL5oebmDx2Gv7PVMFU8vBxIsvLx/fcnL1FBnzt66YV17Xdlfk3yDjM9H3wNornZRfDX
6N447zOyVK7fAqjD5u/+zR4k3LAj6ibxJQzcx2GVB2jACmf6nHyORejHiLCm02DadPSt5JWL5/ZO
jZNIK1pftbY4iL7n76M8vsNwkq8REp1hWJx8RT+5xZ6a0xD/MYHIdL0bBz6UY+0DGPkX4KfMcDa7
lscLTTa1zigtWg/w7dywOCvPmwcAanhFDgBqmOsN7bM5Nm99JbHuI2J0vEcDnFP4fEtlaVGYa3CQ
MS6peLUaCkUzhKqdhVjYGuujn0BMUjudqm0VaoQNHxosMIg9Qu1GiZtE+sywV7DqVLzKya9ushqJ
JBv4nwqgWuB1qQGrpTY/RmHX+abKrAye2Aqc/DOaOdpjYX4Z4faEH/qJAe5DF+sxwYoMSL/hL1XK
58SlxBSNNLiWiTpn5o/SRRLt6mdDeJB9qknWko1SZFaJVauFfbtsRhD5+0PQP60OZ2bqRfU2jWf1
X7z0xlxep96ZjGRxnCU5gdxmAARF5JXayjf0HR2lglG1nJrExSBmHT2fNTOeM723Vi3DggKHXWS3
uMYCA6XzgZ5q49L0koFl35qrQRShgD3r1bQfcYtrg9RtaYLshm1Y4sCwhX/mzYjC660n21Hubsqi
4HeILseA7sI0ZBQ0TMJn9N3BmaqJ6Nx19htWUdtO3pX4wiqRj28ftLbpBMsJhXianuZWuCEo0LOn
b2lS7NEgdzFZvLP3ofgwXurpLK4HB0DjCBJ17JrU/4hJ7PezZeWCc6BtbBugflstUG9I0prAJ9p5
x1sCbYgZvE76gIJBIbxvCB2TspJPrj8dzLeWqjAhg6gSC2KsIdIM88MhHX6ViWwSx4dFav8ox/to
3MfuoBnFM0mWXTROh58lEjJ5KuoUocIb5mgnuWiME19MpcMvKgFf+kXyuPInGn6+Ns6CGtvtyS+R
1oz9AYKZiZ9/YW9mePAqlwUbdTTc40njEnAJQ45NeVCngwFKyLlsxoVb9W95QCXeEB+BHjpeXKIY
60PaX1eLHdGolbXv3gLooHHRXedxb3XuVRB8xlcdYucTuPabkBMe/fuTHmQtBa6cPLRs8e7Aolqq
en4HAU292exKThB14Jj3OwjLGYmTbfwddWUxKt5ajn1onoAJ7R+Xu4yG6gsKi7yFbQKdLYhHLvsD
bzefhZ7fpyA+0vlMuzPYuiVNqNSmNTHEQ64WfnNOr7dHYcbvxmANmItYldBjbnMB5ME5o/xcYWg7
CgZl77b1uH0s0yjYqRfRRSblmUV9iQUFPyRh/TcAImou36yJtyqS23daRpRl5edi4IbDNjybBpek
TOne9qBKQQIsfYYKoaOa7o6Wxl26RNQIIuw7VsHZbUqA7URu6r51v8WC10jZM5UIaN6qgEy60p44
tRnH0wCwJyMGdwsNoWMR6T8CoNnRFqttRAU1eh+pj6g9Ae0jbMKMjrqLStD9uaNKayqUC27vB4O7
UKPCqwyTlJvhzoRqrH9h7n5j0Tx/MLNvaKizzvR+MO9dUd89xu4rLI/7wSq0fHyj1NWAeaAX2333
u8mT+nT0V7Leoj/PxrewFSwqULXi6G2g+DpzEeGRUWztzfYsLHc+S2/0A2r0ny8QC1LPGuZkIiXa
/tikljh0nt0aQY/0LIjDtXaRGdhyBjJRVPhOJaGG5zp2gDHJBA+HRzFsxu+O5gXe/+fwFxWkYjvz
VZcb8VTS21rv+OT50B0VJEmsmpKQ8RBUgNFcz4AVmBYcnL0tObjmKMnMC+Q299pa/Ll4BHR0L3UY
kI70CbpNYdUnb6joc/6cBSs0KE2uhkU7/nsPulvjRMofCPLljD5xDZ+9ii6bTXLRZX9FF1vJkY6p
WFRDbkX2O5r7pgQm/VdxXBSqM94Absjrf8i0qwFUCHvie/wz9L0TLb6W5ZOjPl8GdVNSvSOiqq3J
gyFZGvBZTWzW58LS9RWaXXO42atUuj+1csAnsh4Vytxo2IlOL3Hdc7rttAU+p9JJTXaNWM7P6shj
to+WYZzorC4KNwuGPx1fLR1YpRtqP98wf4+zTCJAOQQ2QNbTxlB/NTjCfq/aWnuOiklry6FHfV2k
5yxuGxt3CvjmZW/YqlzmL8lVYmYhZOIiRKdWbrIYjbxJLUVqqgmueTRgSiBg/20Jt9/1T2p9F406
zJfo0H10nd96Tur7mHyGaiujP6F5etqIIBd1+s26u0ccug4KsBScl5TZguxGPKkOF2LM0mIVhq0e
vtrrlyzfphvAwI7QFlz+PQP+bWZqT1yDmwQcQeHqYoru8vd/NgfVBXub6C7sZNK+qes3tmfnarcV
pJTMZIz/l/q62edpOJzBrv7v8V8Jb3XLhSf2++Q6i7/x7m3Uo+jmrknx4OuKgHA/sZfUKPtciAFk
OjrRqQi+Bc27+rrBTvwgx/D3znM8uYpVVXUWHEBfWdD9SUhZiy/G6E5eXVdDs6EpBkG67+urLSyr
EOwB49m0P8Pc+vzc7RctF+xIgeRXOPxRpD0RoeREq1Ro42myai7vJCPcGZOjIggknTXUKXKgu3aQ
RrAmnx+S44G0soUSphH4xFwsKRcwDlgBul81SWIONQ0is+23Wc/IBrXJRuOzK5T0cKOz/EusNsO/
gemeR2K6g9eUPsNYVmna8H74iQfGq/8/Z8Qevx3ZhWy3nDHkD3O6Qh1KuGE/98LxZzwPP2C/UkGW
wnqXffAeouANPDkjSioSeWV2Hi4D92RXgPEuDYeikzpjnsPa6ZzmEdbKFfNsYmJohjaJLHwFLRZi
nXQPgOcdUEcVJKkQHfnKkUjgwzevQAYr1JJ/TmTO9292snlIa7o8rlMDqjyMLKi5VYoSM2Y/CxLX
Fxp5jd9osBtYyENXT2le4k48rEIAHY29gT2t+Og60k5dY5+2YbuLJq95Q2SEtGuNzdBdMjVd3fch
zvMozziTV7LFyCZIayluNo3V/IKPl0Fh3+zWhvErwkLdBsh3xPvukq4zGclESBRA/FOl7WRfjTbG
g1p1bhq08qy9MAU7fstEFEcyghv7mQvTASk8CSDYjIiFT/BeNe0LpTFaJyWdxf415oihAVJYWbr8
ISS6bWRoWT4HT50T3M7Mp/nDGc4EiDj43Nlj8PJ75hYrz/twcJJoWnJtBiZ9ehjsAjvqFmTkTUnb
UckTHjlkc8n8Cn9Um44+b8ygO5kT670fxL1ENDvXexQZdlWZhn/hzDTNPUUqnmssTG//z4tvRN7J
FBHtWW6HES8MbIb984cUE5Jy5G/Vhm+D+4tSpU5Z8/aR/mzMexylRqkA3OmmSqMG60R0P5c23sZ5
vTD77BOmlytRSSTeDudzuF3fsOypDsxHhBlemh5FGyeYBQisPELt1WsrNTEeZuThuxcchi0IPstT
ysG8V2bl7K/qMFlAXPCDXN6vTeaVXZ4PQToFrnaQY9G5IumMflzPfizyMcMPZnWZWLsYZOsujbqN
osX48bh8ebUcj0JAg+N3kQ0Tm2URU2NyGKgyMBbwxnNtf9h73dbwv3IThdIConsDbNiXhp1MRvh/
4zlBVRscBDnIw/7SKnFIXXoAQlm1rfeRQt/YLsaxtutfodxxycxxgDeqhRkKUgE3NDn5GJhyxbUE
qEulEdt37JF9r8Gk+x69VvuFwmigv9hWWI9nZ5VqkwTV6z5QPhkmgojBe6h1O16kwkZBnqcYJdFa
LXu694OKQsWZB7LjWOOR1VC8gCxGk7Q2w5IYcNJ5DIBe0g2dKe3B4p2I2fhhQbDxDFPVoscc1W2L
OWj2VYm/px5PSfrHIomNXHyrCRtLlIKRvhYgs5dnmuLdafiqUcZIX/ZUchQGe72e0yPHvia+LT10
iU+Ko/uaTcpZuQCF0wrx3T6aINQOo5YyXOyzijxg3ZbpZBtyb5XeKhZFuZ0pBxtYcxi3vjAirHy1
TD3SHokJCKOf8o9+/rom4L9W79TLx2g4MXjNpVorR6D/e7Q788/Upb3q1pgb7vNmsYuneXgbQKGu
bkYqU4FGH+WbwVQJDkBA7zElMwttcuhOLKsXT2py8p9QsCiq2MT+QFMU6OHkscFxSZ2OScgS4YgD
0EU4lGdqPlKBw2SoxX88yq88OqGzEIzavJMan0Z5msutlNOieGIrmlj9bFOKrMODY6/diykLd0gU
PrQrtgmovBSlZ+PFGV02Po21VR/Iv80/6f9TBmzajfQK2OGqjFWa1nVNHd3cW+chBP2vaIdJv97B
b84qTJlkurWDhrOOGrQvLh/LbH6zWJTDR+CtQRhhqsoCU10ygr2shWc+4dmDL9p54TLtevXl0wXw
9x6lmwXr+263w31EOVL6SCRLt6Wg3QK4wYX6Wmn6CLtuPL59+0u5vUeCnbW/Md7fm2o5r46I3j9D
1wcUx3Kn843a5NBktOyMxHiQq/vETJe5VQ9T/MX+6Ajntx4E9hnm/rbWiqIOlOaGrF6TbDbr1KpW
18ABCwH8uwMu5vhhrHApp1QGAcv/RKqlMcTtwEDg7KCTmJvs4ylo7tj9wZTYmUC4BPJD5Du/oHpe
6xyfuooaLw2hsIHm5VKmbEcIo7WoYLZz+KZIb+9DSI6w/bSiH/TVze9FH9rAC/GTPZC11Rekk/Xu
2VD8K6fyUs7q6ua47Di+MMNpBmSrjyDzss60K+iSrZBKE9wSBQefz7HGLNr3+2w9Fg8TPcr+tfGV
yVZelY77M/Iz2M5fP+jPjMvYlqb+F2fr+wQkndIfwHFkviBYC2JLPS89YTjc+swubrmGE76LfbnO
qXXk0Sd9+2nca8GZCx4PbTSTMPJ48NnfQSovQg9GcW9JdSVfXeqIm4kel++b0NtxFcpTQBzON+/Q
svpY7a5GK3kHiGaKmNXB4z4zHO9wbmtutg/OCCwM2JBAzB7jp+9TkHNVpQFldinZOq5//oJca7F2
Gl1S9Oev1+skfzw4J4l7XYzcxdkKDCIB9uHHQCcfIkt408AVkxM3q1fdX1sBF+fM0QiDI19wSJBu
aTemb/lGPnrcFuavs+Waha4jTxzSNf4FbK1Fi4sHldB4GLvarmieby2nF5ScNEc2ani+WRpBxRSF
5enNJPEtorhiGZQpAjlwFzG0a9+vwFAbjtKD6rXZNwJ2ev/ORLUu/BL1EFleC11+E3W4TJMSRr9B
prGuDmZRSDjZqJXIxeYeAvdyN96y5Np24XOJ0W4RvS8Max420jRH2AXWGUO+MIfcAJvcrx7LtAA/
hcYWF051agUkLVCsf+olo4hiJ8NZj4K7Ue1LzYk4VfHoddIc2oK3I2dpcGoUpDL+WMPblraCpVjr
wvb06fu919iVykil9wXQtl+UtLrjGwjP1J+L9qeO4xxChADPrsAmZBqtFkQIcISkJ6+J/j47xKjJ
V3IuA+3MP+xla0Qum8PGdtlXnawD03UJqITm4xYnvSsproohFwI/zdlF20I0HmRqG5k5U/xigPY0
oYmUrOy3h1UQDjQqyjUEEV4gWK6aa7fzmH/i+f7whnjm7x0BzLOklPIfQLS4I/44wWhnZ0cjvHgi
VNec5P77qXheOjvdBc5WnldXTj90bT3XUBEVNbwajoXt2gPGl4hDpo0BmIlehXAnLAGU+DThNeyI
kZ8hLq1MCHHWlP6FbhKr0g6rti7xVWS6cAT0rbCH4/xn85VnVbCx1Ob4Y5OCxCICPcPa8NIW4atK
aguNcphgC5j1mRRVUGdlw9AeCZII0t5ryXRiD1pey/VgvunvhE/on5WKvDLqRFWHrN2qN6PGgqm3
Vlstf7AybLszTYkq/eOopmeodDOCoqBNNUBIWeZw/naWZQB0s6kjM1S/lgX4A9MmafygroYsF4RP
5cvyTG8wlhy0hugsvQH30ZQrtxFELcr2Dzevoebh36+h27Da+tyYRgDNlJSLGuaxVrBVWH7J09NA
PIXRIt9fpENqhchF11vrjkpt6PQ4nUQXkKVGXkU0pUrMUWmlBmVL6q+SiAy1/l2GIX5S8UBwz93s
SI4Fc7uC8oROm+6DCmsz08g2EmJxnr4sUGShqKBn1ElrQ96mBRUj5GMS/blEJjVY9+H6EzK2UaCm
qdrwMpZqMNDxILjXm4Mrv1bg9wUTWcVxwG3luztyaDqqF1OIOWlyw0S2ZX3YYHDaplbKb1kFkiOk
mM1ebHGAGka20cmJQL/ap0UeXxuhbsxPLo222VgSxkgqt5LCBSevTHlRuY7SBO0LM2c5v9K5PmGn
5FqNkZMGWsz5jy3huMbdcZ/MeeaJukpecG3mGBx93iIjpIipHzJg1x7p7cNZ6BAFIlCpfLyeBRPQ
KWKH70PxYylvBf1sXXk9X1j1h74u3TBR1oYFlnvvN6zm/lrwN3PXRQj0vBNrXAXDfE4ZG7KPBWGB
jsaWotSel/rQ61Dk6o/eIW1+cgqtukQSSWhvDyF0fhv7ULPWuri5GBkgFzEi0vnWIuuAvLspQf4A
n08nGXroH1BJukHM+9el5tOfqV0NHyyBgQmkq+Mq2wo1YrBVhzt0n7ixBDPaG7a47GK6lIRMCOH5
83irfMPXTId5Xcg2Ju880tVr/zFlq3kpNY5v/jkabnrWfKoQoZe7DxWu7YZg43Dsj6jto0lMHYCK
ejlZnPVLggClH9oSIDlVipYts+hs7p3tCjfG8Z1If1FFMUM4pGVyOqYFpsnWrb63qEVAyEyMka0y
tbNYSPPGdk13xSrlLb8BvejyILRRG7znnL083XHVmxyx3l9tMlNR4YYks0ptwEvpNK5h2Gaf4nat
JtDQBpdRNCmibWdeBY6RiarH/WGO7hVY4vQOBMURC2YvvWdoBwEwQulDdOx7MuCjTYcQ7Lp9DTg5
XX2ELrhOgPh4UlVkAZ1v0OSkMulAYZLV7YMgjnp9r5uCZ0K6wUZ7XVgb4zp6nfS6BLwcqw/tdw/5
yVhgRGhIOo/vTtWAHYUoZLR0t63qOY1eTf5Nn2tClN/6jic+dAYsHpneGKxAJETZSTP22RCncU8v
RbUgxIrDJQ5wcQF9aAU0sWnhiboTYoDf3ZsxekZoi3fes1/A5mKedi9K08b+J+uqBBX/mH1pjgmt
G1lqO94pjBIeJmw2raZNyqXBAkLkJ4xGUB8NHfWCtx2tCy9lpuo36Nc/9nUq0Ok6KKKblewi80yi
oraXdBGQxRDUpAz1xok+Lu5a+ze+4qBSJr3qr4h9GO83TjDGi6kqiY0mpxY6q2ow5XE6D/cXReuA
3vT5VQXdDEYmCCB46CODIWqLLshS1+LWzWrfPv9lWVuuSX5U6qD7LgnMAc7oAyoREAGJm8DUCjXg
YpWsFvx/5Yg9O7aXqhKcJipA2wREqIzrXKkl/XXkdSfVhJ14CObY2WV4xSnsKHp7Zr6rsn/qoc1E
oDeRKW6ljsscVbzlKZpBrjn4n8etPluttJc19LpTs/2zGY7E12CnmzFXBBuKbBEvvbBEdhgKiz+F
q6teuAEjuoyfhr1J14eTBdDY5kloyeXzpPKmKKb8r9he9Nc5MoGMFZiiq5A7OAsOpkUbAsLxm+Sq
zWDH/ZbR041H/tulXzIqWyzHQ9q6bFsef7yGbVqYenBdFOAidMSqL0aqsBAUYOhf9Ov9ig/DjI6S
6s7FKAuav16bIhI8PHATSoav55oVgHyADI4wxutQJHFq8KzCi/RDZIxz5QhR9jdMZYzLkP2muWcI
zi2MQ9UCP4T/ukcwCZ+cFhhAnJKKTGSD5OYh7olm835YPXd6wrLuX581xjFBaTCHEcY4/y+tKxdB
D2ba61q5W/+lkqZBQzTFk9plQXNKu5qW+fWOtEJ/xKhwvnus4o/W5ZhV5oOcpUynq5lMMLVVkDdq
7fczxTUBsAW8QYoWEk9JjfJznxObcyPaCC1l+MmUPoXRU2bysdzIcOXYzHSe8CgAPsdiQTPquzxs
ml2t50//yqZGmTgMa27aJz3xY4Dfk4fSua2TiaXy73YpCrSEC4UnV0n1kew6ZH0PV4jXdnf6RKYY
nbKE/Fd4YIexZKuJnPgiAllpgnMHmfFUTaXw03qYMi1350aQ7hZmz8/+Qh+qcAD1FpoGjR6tmxKx
p7GLIDRhG53aL14kS69NFRis7n0p94sCCfPpjolY5gmbwwxqgbm/CrzdDscClUpTx2qynKs4jgp4
hMaT2bVPK3ZfW/QHdfm3+gJ6CTX8uRMAl73vbeOHhHIuMj3ASZXvCVpu9sbyzLRdIIayrkhMKZxv
MnLaGp2FCuikeBZNA+0bpufbuT26rFGGzBdXCHNj7NPGI4sorf8T1YyAN5vp5SjfSY/H5V86F3Fx
voVLxpR5S0g1w9anntp3bXYZEfyNY3ebRPmmommAYRWDRk4vasE7bWFWbfO6Qfiu++7izrtypJj4
6fFOh/39Fs+woiX8CBZXxdTpmA00lDuaWBZWp53Y38qngr1Kpb9DMWLsIAlbkAU/aKWECUZMSjy2
hSxdwrjkZbilK8pzrpFNgHyJz1HkvqCeCZW21iwQivWXhELOkl46Mz5LbcpUIQyaO3+egVJZuGvr
CdxH2UvPWlb5I5tg/KkWAly5FTTA6yHcDPwSxytdVZfvyLnJa5PwNx1eISKOee7zy+HyP57lN8mL
bbsN/pWFNjzmoSXK1BAwT9rx9LN8+JYhMQ9bMYxgbJyYI9t3q5rkMnPHs2DwST1tu/b4nePrxWml
wWnRuRwY06X2rtg+jUOxHMJsQcXa2JW5AGTVqdxuXmCGx/WyGmnswSWJYEFCc4IFHpqOPJmzHmCj
kH554fW40QLy3oCzQKhBw6JAJiVlShR3o7X7y06uLzsha2e5fe7dx+l2zphfdHP/vHvcrKoBXygU
pKBETm0J5uPVLd2I9bY7ZWApvjmn6I1rE52XFcgED3lqmqX8LqeK04rEZQ1mWA0tbVHrEQfjux2i
p5TdPe1f9nyO6il7ckdWHwANGyVi27GCwALDWhXTOjS5IWnGEaKQG+47fxsjLzCAZXtK0TGgbxcD
faGkw2+58julIEdp4/wVQ4fEnQZnk435kBA4K7lLHR2hz0BFZz58SB29NVkso59VkB5R1VCVfHtY
NOgIZGACzo6Bf8+siDLMbOInGqKe9BnMyPNJiLVAZOmRuyiE8LiwLhcYxuYI5STKZQPYuNNCJ/6h
M7OF/X1YlNqvL1shhaoHxVzaDtQ5ATZXNUCsUq+OIRQe5dmg0zoxedDkNwTfIuaz4Awb/COmPq1m
UWWH3VQsMzkmU4qX63CoTK2t+d82lLoIh9pSKdbAOV9gnwpoImekY1sstMv/QSz1GmSkcgCJfm79
79wPdpkIEXZNLI3OKxwGYqJ5ecFb1eBVLSoJ1sWRq8Fq0Gld8I1tE7NKLpW+qK+8ym1txe3LAYox
5SQVG++kYCMZKSMJuE30rd1zoa8yL3UzRSPOoppVI+1NxPEuxLatOxBi3tRGCemJ0LVgdRQ/DpTy
RinR1KRcbQrPQENxEEOqFhGI9K63QViM/kZvFZDLp2UR1dyK2kIN5uZ3JnAT4Ly98pWcb1y/UVRU
Z0NDnad75SsjxkbTwdEQ/6DQwaWK7ugnM2YK6mwcIiZF0y+innl3xwbsQiAD9OHsoNM0aNW1nJTO
WNgl6dD6zP1eW0UpR9MlIslefBNoWQJY4qXg9XS2b3pvxdC8601EHbVIxmXsVooQLSNGTzvKCogt
7qMuc78LWpw6UsKYbnDB6TiiRQ57BbDe6YbA8qZyH0/OpRQWdvRgujHGdKaXJGb0+zrUvpAzIrdM
iCS9ZJWJP9QlwyyD2jIblAkdFnOXeLqMkiWCWGCzrJGXQLkykojnJS/yRXYgUu0wFDbQrKO0mjXA
L+KhzNXP1JLKjiLQq/CDYX0TfN2Nkodccu4cihlS8pFbF03XgkR/0g+KG/AE8WU69f0VV7fTnZN/
VU8Ym/hxUQfUyesEC7xh3zIhdjkWErPNYFofMMmdIUSU9ffED08ZXycw5VroYFbswYFF4SgURDbE
uHhb69wNJZ3i/ENUYF9mu4YFIL9V1zfUjQgleDkvcbFULf+A8g2RROTeEqe29GiiEzvNZWw5oGjJ
hV2h8Id5/mAJCUkHlpl1wpO3f7C8Z2aG4BUAXEMgZLFoB/MYYDbOywrV7deBQ44g9FQJW1NK78A4
zhPulmHyA+H5jI5Q/CTeiD52Sl1x/4TA7HbJzJ1VtrznfHdN+0bz4qb6/F+JtXqoMiZzeSZ8UzfZ
NtmT9nAwXlj8XpDhc+4kWsviJRwbRPIJdwub99tvPreS+8RsRt/gsuFj2nkvEawq4PnvSyEFNIIV
UwSsgGp5w3pwyDppsSp1/PiUbgUggTG6LLkREuYfBdg1+/Wf97GJrLjtQvU5SADZyLrZeLKc+Bpv
P8+/mbWiqJP0hW5E3YVOHIolUV+03KlAcTHPoHde8N46wAIzGMMyHJM+l1kAdOfdteCDGLJpsRfb
HyOR4WRYUnl1+MRUe0C5tAd/2NgtRB5AXHOeCL5+gN85k4uh4n77dbxNyUDIgw2KNknpiULynUYd
mPpoHNqhNfLg0MxG40+j2BxmssKNE0HYTaJS/zwIG5vJJqwjrWSZ6tBCQ1Jw6ZbwBWW82XAReGRH
dr3e5JWLikZfE4+mhYOIJcLd0ixG15GdHlwnb74HIFFP09w/5mElAxATCAq+AU965uqSFu403Qwh
22wbeJerR01Rb0iVNgJnFr6dVT8dwwBPHI8iAcsG+s41lUb18F9miBs6rfwVJoxCjSf7N1dJwbnK
1Jkx45B3g2qqepgaw+hhKMsoYI9DEL2CA4DJ2KojShPjQSKFF8ECp83D5vQ1DX/F0yQxGkQ1VQvN
zB62LO4B+OoUPEdV6pIY0Rnrx/iOW3YFi8tCaOhWj5xXSNMWjcL26jI++0Kk11fpQvIbmcpOx5Ka
bi9mhF6Y1rwTzArTnJUSAMlHJ7xvpkvIM3/9jXdfxpwLklQ8+naV0+1wOC1jYo8ygl9YDOXaGFBR
BmLImZ5/R5juOBv7c59oV9gY8awvdRb1V3v/RfZMu0Q8e2LIOEHlfGFN8Fh0PyLbWhTbgsFzKMDg
agqxgX0sBsFdkx7UjRVPsqYkHQN7At2DAhgs6J1hfSro94VMzdbPlmN+WgPimBxzURYpnC3s2sZ5
UVuClDbTihIhgjgN5thGinWp96bKccVwyd4uClpH3CFrafDuMbP2ktgHw1yLILtlaVNgkuyXDuOj
0pMuJB7awaDcCG9fcIaaGIsmw/HipGG93gfT478XAR/XWcIR8JyA6A5gB47QJ9QFmXXqotTZGv8S
10ItAuETWx0siaff10RnnzzrnXlAygvN6rZeN7VVsuyeqUfodrF64STG5CUbxAXhabWBME5K3kKC
K7OkiH12i4xY4CTFz5Qs19XWNWWAPbUB/ylq9uBmXGtZLzg4wjzQwyqjMAxiDSwOnFsyHaV7Xw4y
mfvqnESzuu65sup4+q1tA0/ttg3nRoX6NNW0SEGzPDz14iC8C0gQuIFSacL9Kll63e97GLbIpF+W
LOcCD09RYhakBIFSL7u7gU49HeJukIdqzpUxCp61PHxMXV5IlOIIdQyCqFebD3GlaE1WcHjy48Fx
gIWwLq1jl5CBuMgfNb9y5/chPbshzq8FpdnS+MPJzoFHtaLPGIXqz7oXIhpZVJNVmPQNWSCLnCQH
F6VwtIk6y0t0WADFRrbyV4vZ60hmF4IR8au3y7fI/z4Du7A2SGGeWKIYKucnK0j+6Sst6RgCrjVW
QrwPUlMRwv5xOczoisC15D1wksNchElhuRKaPyAuu+C6GBQYbURGEoxUQb11favA2jHwstrPbyNE
zH56f9+94BZRkq5j9lGLYN+4X0Bx80A+u/vafq40VWesvdquLYjg9nfT63bXYstU9HLvtO99sWjC
gf2yxfewG8YRcefzKnTmiZeg0MNvoKCxBRV4+UW/gFLM0a1R6JztjEXiRoR2FfeLjuowS78xLOSy
H4r6XKOU1eqtA/YvzSrKKr73CXBZhtn23t5C56R0kCHQiqhltAbjVRu3/7f2WiITYszijxpXc9d+
WQ9DekWTffpUqFtYJYCqcnTEXCkySCL5QwvU2yHBteHXg9dh4YySFSGzdaH5c/1QM1XI6/td8rbp
bgcGtnR6acmtNt18y0Hir8AxgXwQwaZ78GyxyB0YvSlDTcnlSX3PXI9kBHWwLuos8ODxK8Bao8Cq
JtqePSa7oeNyWNzfoEyPszrVeFFCDt4toluyPdXekSBdeAdPrDeYmZSzQZvBLEnMwAp9dceBQTiJ
gEPa+8r9pPashoZ8nfyOktOBey7UcbUcZ//mw+jlDyYGLwV/j88GhY2OYGzx3JQ6EbuFj7ai+Jrh
nmUXleY8Qai4IDbcQkNbwP4LtBiYEecA1e5F1byX5kBghCJOcJOt8EUEygGAZDnRN2AilhALt+Rm
1/6ddVpAiVbbZKoo13bQMxnOi4RyFUfpvzYl7COqIAF+0xuMPRNaC8pjjFn5gxiOjn0wj+gGiqT6
RLgWXOAGQarrc78FXR1TCZRQ4siC4f61bffz08TJuwIBEPtn2qN6UOQhRb5FB2jfzEQXMZjuTe6y
3PPLrSCF0jaqRc7Glzm/V2jccnIrIeojKebyPfYWgpKAC4/LMgevEYQff7zAugzrskFnuofXskkc
PMUk4UMc90gcieYHxRD+YP6sDzJp7Q/QGdanx8QqMFYp6SEr1UPWJWA05YRidXmRkXmRgVL8Hjxw
BOcgtC14SXxiJ0CEIPOhENinw+IAjRTki/tif4yCG+UfoSCzoMgVrcnGo90JgxQ+ithPm20W+iLp
s7Umf9n9vRvth1kaczoz76Kj2Fuz9BsHOe/lep7PuDe5ka69l4qGBLNV19Pqd9dqvXI821MKwqLD
KYIiFrPV+gvL4YMtVzPa+T4NWlxEWDWMb2DyLKQW8HnAE2GYGabgY3mK6h1ZTnZF2kR+H6K58PGZ
DPyUK92Hx3oXsrP/jNA196KQpG79S/a/sAb0J/tfFvrn+p6iRjTv3QL78++INJS3+4X1sGwQDlPT
ZAWYpcEubLCdayjuNL8qerYjGPA7T8HVX+z6+2vtoGVuWeJ2fsiU8yj+m/MCKi4NRw32PW6Ckdq1
ei5Ral6w5fpFWrXXb3ZyPyUEA+AVUasWelsNeMPGcWltEgkZm7bKoRR3ETN+spsQE+6k9NWaFZ8U
etsFADyv5hAv3iOObc4fZvqtJrpR1vn91uzyY/6C08Wc5WDFtWfa2sFQn7piiET5hEidHczc0qh3
LSpHgOV/qp9Jnmhn8cVit+lIcmvHBkgUeKcJictKc6rrtH7rwV8JQeesNjiyO/VYVXo94UNk7plu
hq+ZoyMd4+3ilvzDwy/cseT6zQX2nXjK43P20HtalQLUo6PFnFKHMK6TSBVLkY14BuaD3OQweWaQ
1sRf5L0+0yY+I4cY8sKWidlyPIV1KZaQ66oEkb/Pn5W8+yIuCE57m5EM4AHtx6pUf3l740nqxGkT
Y76EvdFRMMa3lwpGOu/B7yLy1pChKjquerarGyK9ZpSR4N/kJLTmoIYsq7lTF572su0h1Xyky3Qd
CHP8Dr3zh0pevh8SWZO5XWd58MfGfJ0kYOvYvsl0kudZAtsvJOFtYmtPeA6wqBFvyujJGU3IZbqf
+1v1ax+F2uwmlQetI0HLl+kEe4uxh8+C7s/OJzInFwZrz7Z5O0nxFxtL07f4HWH21hg3ng6oVNl5
PmCwSSEk+bP35iYxiRZSV18egvqOfaaclrphzscVtn1Dkcuon1w+3eO2goP0fQkO3wIssoFQZSF9
7h84OrnjCnfZlGlpGIGqEs4JGmy3Pl6tclQoBwvz3njvQL4CFYuRfOxzhep/mSmwCLUTYwVQYXKL
ulr+1oiTSWHPh2EaHpgFUDkfSak1QFNV25Sx4dEUS/8uuzVVR2mutYIywjhI62ejBgpbDxttj1iT
xsfjqb+VAgwJkxQWZ6hpDuYSWkWS3VRuZZ47Ti5IUoOViKYViOFdgs6D6Jlq5RTcRSh/5wY9zsqC
TVGmngjyNiukLl3z3TAXsMvEpw4AjKZ2TFrtAiQP8HU4xnliTcl2dVzvsJfX/zk0J7/Hib0C/guZ
FjgFOUAx9IyGd2DQdR3obOjeM62e272/0mNFbuwcab2BKPwaheIQ1+7F4RFcB+4VDxhKc6EufUO0
fEigS1KCb2Fr1GBLLbxHlIM464Rv/zenbEkzJ64OBuWvcaF1ohBI1ytmfB5654hPtbqi12iJoTTr
ajJIs4iWpdJEf3poyfdStnJwejtTqYzwSiGTK7u/7mgZ1QvD8KxMNdkMbZnpesRok8w/bJ8zUmdb
Wqv74BprB3HGU83DNeEAbhJPPGFOOld+FLYV2J2O9SEaUbkMJ8rP5CtHRakak7TEySd3g9zrp2w9
PSL5iEqbw79mX5Bu60upc8vQrL1Jmhx0uaQQKjppvci+3xUGPsUARZEYUsaIbgNQHyRorvplXd3i
hjx0TT0Ac6rNqLv5VmUPTMqmPJaCAY5D/JVIkdWtUMGZba9EmOBIn8lkZBs2WMt3ETzkK9PSqFR+
fTv3fkqKGUMLhj6OoFx/+g86x1ltdBEzVJJZh4qQH4fAkxKhWwzjJKFsl8HIJf33aX/2fkLx64nm
YgdKChr5USCd4d55+gt1PTHsqxlzUbJk1ohoZ4b4dwIjZ/g66C7JIFH14mV0jjXw5bEy2rvyJ0hY
sgknrJrI4XANZ0aZrZdhvdoZfgAhIPhfEJvlmXkYqXvPs3+ejeUFOXho03kv1mkW7Z8O822BvBV1
+rHTBie9pd9vVT0EpXZZhl3DYulty8RQCC/q63/GoaVgWpVd6NUFWc3zdUkSncWP13YGFmspPs+A
E5pWvSvljHDvHkX5WRtStOLTFuuGA/0IhYZ0xickcZlwzyy3p8FLzuhEOLbQWzyhenwL8kNFDJ9d
vrKKh9ldmRp02s7PVOJ4V4rrEksWk8F8rWcK00Twi4Qc8eOpgzQkiRDMuyATpXkaX6M+GXO9sAW+
k3heJSVBnc4otdawQAL687y2PraSCU4CNY3nqfp8dla7o9VBDHh5Qea0cAoTJvWsZmDDvg03Oh8j
EB89E3S5thY+MbhJ+g6PmW6B+rFARtDn12bzBT5UKMXRa2qF9l8OYNqQO1DoLnmoVC6mUBUutJnw
sKfDk0RzzphnElKu9EYLVtLE44oQNFTHj97xdRO0sXA480kRPqjkiSnGl9sxYrxuo/j6M6JtXR71
F8XtkD01tiayZ8t7/O8urbmDR8tLeK4Sl3Kh6ujybG9UIdsxsvNSQZmI5Hgupzs/sTyvdOhpms6R
a0nNKLrUM1GPr6kM3rwFR+NbWhdufqmBq3d0F2G/mDSi29x9cFvoh26YT3turQ+PFgoKqjwTrOy1
HwMDn1BxV4+6eqQKwjAua1bCx8xosZvMWVT0G/hf/ZGHX4biYGN+KUfOiDyBBPv/Gfq9DkXV7OJe
a+8dRjdFDCI6e/jUhPk5eJsllwfFPM+mBgeSM9nDbAuJGfXWAv7Lm0Kr3CWG/iYconGxcT95Tke5
HEwMTLyZBvCY1cWRUb7skQ82M4ppm8He7qW7zILmupuUfxv2oG4rwxvEfeUnWQ6LQk+KT3OdDTJ1
Jc/cOCSkLyJ0qPGQ2ySUIjgahWHlo1xcOKNVcTv7ymtc6HPwbzeAjyky0Wtc30Veg3B/tu17wHBY
NMOMQv1A4jEELJHMDJ1pfUKh1ahcrRqeyEg+sFpujbfsqmUJnva5fso/qmVTXEeJTTihu8oxwHxv
nPuKp/9LrAZwq8krdV8tSZxHlDSazQfvpcW7J0tQP5LR64vzkmD6LwAWIZQ1d3sdCEaz9ptCARlz
P/3NR8MRo568O2rkYvST5zOAqV03CY9Zj9ALLL0Z34ikuSwDXafx70Xhz3SHJ+ZtRGhzCkC5YUho
kVB+2i9UooE7RuKPtdiXi6eQ6ATbc6EwLTiWlgfNTROficay8G/UqsWx2cQrJTYwdAD/xsf60oVh
9a34Kb35+Nt1ZBSngaZ+4kp+a0+8ah7w1sPEKx0CJpk3Xz32o13b7ZbN7+GCR5Qob7H88kBLfLaR
YazecqdKFI2+ZPggBmnGXTsjzBfJiUqM4/wV86p0bHyBGDJTPeyd+lZjDDfeLLF0kWf0BB69SWzA
Vw6I3g/cjAVw5OW1f4vzAcdYPoqSmDx+x7GQr7DkI01bLSUDCPlOGNOfW+TBYCHdfbevNPEayyPf
NMHRL3EKvUgv8WWfmC4O58dP4WwTHu32lP9g1IT28nIrWJ8+mEGCMNrL74eRz3QO5+FJ7N/6dHYb
urgOI2Rf9hYP+zlqokOMV/Hz94oCUw9rDYG3JoCBrR02dxw/8eMSSizCdjm601Mt11DZ1fG0H1Gh
r3fgDk77l4AZ4p688C1l/tpzkLcQ/anNiqoaRhI+k7n9/vaj6xtSS/yctp1lYloQJjbV+pjWl9fy
KbZq3o8NRMSVzkQ6Nj9kS8WiOjn5sqtNyMAixwD3WbsfGJz5xFJHyEP2cXB4yO7Xz0ACWqZZNIxg
tAYeGTDuR/dYHqCSB4fQgsNA1kKQ/ZuMPaEyd+6nEvZx8AqWniXnbnqLVggqGnCSkoJ5iU3tURXm
ZZghFztDkF51/F0djZkQniOYcQRP3dS0YfqPPuDe4KWRUF+AmgFroGWN+fT96hMhJye6jtCTvuso
bzROFY8gZJEHYsTors7sfYuMHBb3Jt9Id1sf1JMHxtuGMsoLNwpI9rLX4Qv7QZPMEsoO0bzFo8F1
QZh81/tAAPwt6S77j86PCdQH+iKY0xgWOWaBfSjofK4qlTwfScbIkzDHltYd+ssOREWNly1bQsZw
3pFO50BF561KpD1IEJypj28RnmoUogDlRJJjBnB23jJIfaHwb6ytG+vjIQJo4DhpsaT8B7g9OjB2
v8divkgW4qay5fx2hJM4cwwguqJSFCI45qUoio7G36miIev8ukQafxnYuepcxOzgXfR72sPv1UsE
nR0ZkkuI4/8EUgldSYy1tmmbhoRHXcLKeIGA5GxFU3NIleGAujJUCJYE12ShD0jzuWQpPoiL+d5u
fEaLmeQfL0hZP2i2UNGTSiuizrr0j7Gb+4z5oU1AP2siQhQq81mp9URnYqZZpzv44U0krA00V4wI
w/NubBEamwkI0bvpy7kU1gZx0mE7mLUh4sVCEkCpDmKBBW9CFaVYoFX9Xh69cthNeiEteZ1ksSTT
biF0Tsg1cjgLbbx6g/8mPTzSiDbws1CRMEJKHaUW3oDv7x8UtFqnzo7WSFMXsfK8UHOhLTrDcx9h
tMnP/XUwhJ2imtIP2h81iF7o8HGtRhX7vIfdls1fyB6OGGEV+ukIYXfSrdt1ek8U+TSnWnK2/beY
TMGK13+SIbxln6sLefsEoFS+fFwnpG6YIf/9PDtlZEar2EEMNKqiTRyHQ6hdZq5i0cn8g2dkvoFT
8l1A++qm0V00zOlaBDMv9tMj1Jg7Qaqf2xrgp0n7QUBqY8qfNQBUnLB3CXCdDHZRutpu6F9W1nCb
EvX81q4FRcBjRYf5boa05nV9fC3NvpERYDJDYwsQAZAXaC+JitHeorr/O4hZXWBNINm1kPep0vCZ
2iTRVlVhuD6lcNZuPzQ0E8fQl/KuzpKwOufPwJSH4VGifwZTNEISS+FsQhhJp1Zuv4SSdgTtjeCa
rgxIPo3iDfu/O0MQphOgkqo5EGNhFDSaw1KU6S4yUDhRV6BBtbOpHITybmoQ9SVGhf7EyUvtny+t
vf/Ny8s6o2Els5K4wCPbuWomiLQTlQfRM3yLWf3ee68dNddyWZRWpx5PWUnEHze6DKmdXr7hUV7z
OTWgCuNQ4YadpeGA4I++EqIXdrYjJGBRyq6y7OUWpVTS45s+ufGhcSY6cRWhs63to9eTitH9I7ZG
7kYj5wBjzTui8+hurMupjjsv7fbiZlsIf/kao+Rc7NVHMYXvLkK5F4Ju/KW5u4Ofjiiu+1xOw1sJ
stGlb/Zo9nzxYhXRcysZccXsjZfy9KddnNl14HA3QwuKysVGirlIl0fBEnjB3LcN6iOJzt7yOzcn
crDNie3aVTjeM2T9bcGj/OmRU7kYIM0ebDCUnhk/YDYQeJM2vk7Sc/iWb0ZY13w0U2wAR4IxeIZZ
AI5tE00Wsxqif1jXh7I1s/GxyjK0vW5qMOjQ+ghttVMTOBPfRCfDOH0CLdTUSbSt5UCk3J8DBFzY
skGDAiUld3V+5wtVRsaWQUYL082FpHtHOX+78NcFP1TQwP6hl3GvRbItmQ2LvPrrSP851ZyMsuH9
hA1vHQI8NFOGOoQK8zGOlyQDskS4zh3VhnZW1QESaP/0ITL20r53YzxQ0nsml6m39Uq18kytvK04
jgc6RXqZn9F/agKsllO3YjtO+vnV0Xf37GPPjsAlXz1itcWrNL1t7kuL5T9btKQMAJ32SIW4zknS
+NWKQn53PrM5TGvOccik5YiEBmsQUAoqz/T4pKj8BJT8W40co/Qcubx+JOpSCWKTOC6ktW9MxiKu
pY7kqLlWdyF895BPL1fpjZV6txj3wY7X0eQVBwzuS+6KnD3AoIXWeqlbVeV5/zz5+v0M1xvAVALE
2rfapJcopdiojL2n9pNvTUAEiH57+51oNME4H9WMMFB7dig4yJ+vQWi/5Jm88NLYNBw3O+Deq/e+
jWpTJBXsg9+q5QGaUL1Zg67BzowRueXWYpQIcqFHH4+HL3BhNmqpdNAczpJRtLSfZ90/BzKF0oyP
O3v22cIN0Fw3G4HO/ZF4Ct761A/OeZcqnEiVBUUlZC0BX/YS5HbU78tQISfEMMnRsNPc50fKf/B+
NJ7o3XXl2SArWSVnH5m53elkeghFYSZjqFBpXhb2n2pXAQalB0bvr1WmoWCL+G7wz1A4FH4/kELf
wab5HpzdMYPVHCbheqoHgfc/4pof3oe/C43Vsf8iAF9CWZ9IYU3pXV9lxvPqtvnBY3xbbnQPAEba
fuXBaAV6lOvFSeqM4sjTjL4uSeVpMJIT8bnfqltFeXrtwaq17riRGhQWkAq9Ul19rNrXVZmh0wYN
JGjlHBNweZcsiDNBmVZlhITQlHuvb8b5ov3Yp1bGpSASwNRuwzfMnO6DerHqBsfwguuaAPQU5iDD
FXETEhSsa5PTEtlVSljbnhyQrlNeFS2iAbrzxKPa+/vgMjv7kt+KVbLT42+3qF9ipZHuuezVpPU+
p19d671u+Xcx7Dm3ney+BmiMFLxTOQmOxh6q36+bGQBxxzkZ0c2f3z0ELnG6ugls/HEprA2rtzrf
ffcccJBvqiYmdJBWqAajkYSlWKvtNNlRqSWo2rb5IZmsYiurD+R2BEDu08SJIPhr1g45ZDfc8A71
TjiYuMNmI0ZQVqCWNumNvX6r5LfvoMUo1HWYkMOXxAfDT8yDwW98jK5k105OJUoskMAO/HUEDRJc
NFIUujpOq0IP7eAMHpTmb4uTRduxXj9vnQRs9Bi0CbiZPM9jjDqu1l9ZdRXlMHriBXxrmfP8A1A3
kC2AAW79B+g74+8HTq2lknEXw8Kp/9UiIILRvYmVgjdPpZBzCI9jhUKJeix19yjp/UZTtTs4gK4l
5Txj9wg8666scLBbib8gw2aoSbrey4JHPXnA+K58lW6fg4AYCug6rpuqC1sXrI2bdCv8L2tVwnsy
mw1GKJEl9n8RqL4y9auqdGyFzuxBJlny8Rydbzt9khRv9SOhA1bP7o/RAzb751SD84ztL0+pPhxc
YWBPRFDO4IQLcCtYfXNxo94xOinDaQrj1D03j6RBUgRUmEXdMeJWbTLf27pNEaf/9iOft0B4UGv1
8P5gmJn7Xqg9tH4vQyOblVlseunvfBpAU3ZbrjoimSEjBbC+QKRUk35s1ZVn+uvDdlp7uWYMlFVs
JS3uI7zGS2gMld9zDJcfxIzf0WnJJb4Su4JZNKbq+jIdn2R1ZkEJTm02MImxGo2tHfHuFqWYS4oL
C8CeoIDqVQ2RxeXr33GOaHN8XX4gwuzlQBLzitP6o7VDZN09a4CCZlT7dJ3G2gNrYaZYRlHW1Q0N
zS2/l0s5D610yZVaVepmPdRc5c2DVHYA8318eskKTbmCymC6FuvmoQY+gLRj33owQ3j0wVZGAKeK
K4+KjoQBy+yDSGTIbGUUMM5A8HOck1JMaZNSb0sIewuNhVqzqWc9IkiIv5qFbejuzFC8GtD+8q13
Q256MT0ZEsRDVNhOn1/Ge0Z0ryX7ykdAKkb2LI29EVI3F4hAIuu4n5rhewg/FcW9hiSyuqG37VzV
qGgriccB3hRGOoB1W+rHVLJF/OHlecz4/7F6fz3qEyRZPpQBITPWWTx+nnMkXQg1vgUT0z1+Xr4p
E2yK7EKlUUwW1uq8i23kIcEqtaw1xhQXILND8LmZwIa/GOhtGdJPwdyqxOzH69vq6ON7dbJv3YEb
ILdz0N84NJvj+vANhZEZ//6CKlmim06enPMqsWY7/+qF+BaZZ64SnU9mOjK+3dvrL6apIsFEez9w
WDF8wJhYiFVR3FCl9tadW6T/Q9s+9Z9KD257ZmIjTAvqwOQXJo5P5zvqBTtnfFRR4rn35yrb0XLK
ZhchuvlVNBmuD7eEaBES6C46P4LNrO71lxUa82CGmYZZzwxUapn9Ai9MAfMgg1hMu5ttU4MNeKVZ
UBIJTtNsdH/BtjPjO7OX1kVikTGXJzeb1BRrgaSrNCy60n5I0JLisupcey58/FhSCnQhkVzBXH7k
Z7lLoS5WuAuUhs96LVKVXOy7tVmuFQcZwSSUKbwnANqS0c+7haRusTftBHoUnlauCRaQnRqb9sa8
zq5HO9LbCRWQKCNEku/x39r7OAMZSxHGyImdiCVB7p/U/GghzPjBC+hGgLAslUy8zFnZ+TSj2G9v
wTds63eFAYjWJJhWHteHXa6k6TuWVtpnUTs9hk7LEaAZJKMDfjORw48X1Rs7BsWLptHCdvzcF+gl
JdfKF5g0mt9Yznkci0Zb5zVgXOAw9HDfN6KGKWdPc9xRGbDQi9tzZfz9fyTLWeuj5Lz3RsPxF0YQ
HTCvy7mC0Z2y/z21cZDjxPIq4qiz6/1jn/U6oZkXW4uxThM3ZErZ1mxU3LaNbzyEXmSnx3vnjGW4
e425NExm4CZ6tja4DkxqedyVFJZSuzPOD2edk6cRlGZCzzjBo8jr9rJdgKzjNT1WsCQawdl5YUjv
eFAMAxlUm+zao7FzR52s+DYARNxmoE024FXJZ9zFqdY/AeS/oGk+gL2iFxAexVfbevdvb0UGJwM+
9rWuauPQb5ZUXzB7fg6KUiroP5rXx8/ZHNfxWNIkNk/Cvp7L0seFSKTkNZ8HOYdeydcJpQqdni7D
utQSITFkNsF7wHvFE9yIMNYEkNAKXUoKaFciq5tdUQ5rEySviRIU2BSqjoZMRpCpOCl1EqoNuXwo
lNez/hdslqPYXuPW7JQeAyxNuDbrZkVeSxSML3HAu6zS/3N4CXvW8Tm8bNQLGXxU3z1ZGf97rFjM
R/9yOFFW6VJR9dFuIA3OY9KGA62dFYX3jng+86nQQFaKL4YlDTDFsRT+wcugOZfY62eRl+RSrG8N
hsSD5Ndo369MD6OE640pkJdoXZq2vzFRwPwSYWtKgWftkQylHbeKkWFkfcQVLvyBn0sR2kR9/qAf
fUwntqfjE+uObbUdyKLmxta6TwLSP1PbLs0q5HuUhMTPpTP5yZCC4okke44zuRDMI9BRsLgId3gV
KFHrH2Qz1bj2iz4tbk1i7Cx/8RCHRe8dJul33g4whIyNODO4Osuwam6IFyxhoPdc1C6FQHoHfbbw
U551XuxgKXD1DLyJPv69GGEuCkhK05LpabnjOFYJ+hgS1EBARUHzPaFRKXYlT9luZ1PhQYEaSeYH
VTMz64xdYSMDMsyCDe9QWNZZuvFEaW4Hd8cKXP094JYkR7gJzWcFrFERW0Mgrfx20ZzrhSLqYnaL
1CsBGpcOOkvsN7033j/aba4mnZwrRwINLk1EHNsnsxKDF/QkoUqA0xKYXJN6qOZMQd/rmHJtWe4o
kzD25U+uKQ3YakVO/aqoHiVgyTGobr4vpkxHZmMW+fXG2He33D+1cwQZ9ipp7bzoABAohydgDF+Z
9ZFp2jw6j7E9Fv+T/FbYYdkTQ2A6ZXLVoQYv6uKDtsJ0smHTIw6Dg+q/QvhrxlFExQN6AdthaKXf
sHdmEQdwBcMU4ZbGDE5jGEX5twTiK0e6ktibQ1qVhIwrGsr7UbZzCNSNDRWOAKBGTglvCpUKdel0
utYot3PgijyE2nyupGWEcTXln0ulUNffKR7mhbth62gr9iyEZ91864ZtnG33k9xtTKDlgCW0P/d0
JqAx/THJVuLr9FtAyuQlmPyRPWwyYCsrFuf1Pny81J03wzbPd+9UToujlfMMHkkkimOCSGn1NAll
Qy5ZQuN6rHdaZ3ucTQJ0VIaQ2v2iFgn+dogBwdJvsRFExmH6+JoQbETVha12t1WXxG5d2Ig0xVoX
DX03d0H3mH/SN6gHRhCLYRX3yn6TJKp/Ln8abRmdX+fFN2LjzG2ferBXnHfQMBMfnPAE2izLmX00
mePxWaeZC0a1CqUCvrN3oo2Fes/F3tiJj/ce5RhMLn5HTRnQtaOsSzgRTlFEqJcyTaOlqm+K1/x+
PIBgPjsKmabiMGLB5jSQGVod40404K+Hz1uUAPGeRC3a0VfnyPUx0MJm7XZuVsjAnLBgzAJIBQdY
pAXXUfySDp3dpJsl9vpvrWbOD1eeUia5J4MdTI/Ynj7kUUfk575dGZA34bWpc2r2lB/FZkztpg4B
P9NQ9zJ4uXUHNwgswvAdmXlnhitgqd8CfQxpEvUIRixG/CMn8fpyEoDstgbgFF8ehyLuJPOug9+y
+Gtk1yA/jRtUbK8+wNJbrPg1enoegk75KHqcfODWAxujnme3zDtw6bve0nQz0A3jaZGdQ1HN5qMF
x+JZ46HLARuOmFIasUzaV/XYHZpwhw+K2CgVNNR5utcxUM/KdG/0rZ1Vri45c9czg4C1iKbiGAnJ
TJY+ecUzjiRTYJuhOaQWyjlAeyqMzKzy9y6K923UxR+aQdmiIa0JkIB4J/DVSEUhSrw374bTav67
GzjknjDH7kBXVuwGEIUT81tJ9FFRvqOdxEOPl3kuhmCz/GV4CBuQzkfQRb5K/8GiSg/beHw9MUWH
phV/S0GcuvX56D8ez+f4A/GyCOHyJnxfW8A3qjv++Bnl6lM0F5RneU8P101kPwj8OiWY4WV3PvLH
4uL5xG0T/Ww7YC37+59otLbAt2/vVQdHXI72+XIDn0+mgtyepCj1W+wrOY5m3FqSuLItwLsCgcDD
Br/rfjaAa8xya3aAJW4Ddic07gSDCENHbYXD1dzhf3db8iZaNnCeJ2GVacHoRpjHOhZ7hA+Prpg2
q0ApgcsvA+B4Dz88gB+O8SanvDwM8NnZbLdovShjJhl2Rnhy8JXU/czOk+2/LQQjpQjXKjfsWL7F
/Q6aMGEoohQM4gxGPPyvoD39rj9748/MrFExUBKaPNvv2b9Msd+WCwg21A+EUpWnSm2/wym5n7A9
k2wWLFm1W7a1SpiNPARXHmnI0K3S96UpZEXLFngqyvgl4MdTt2EhUdfeVNaI33BCPGQvklc9JPKp
BYJkLFShIwtNXFa1Df7aEgXABn96BCZKCqXLx9vqj/8Udvb86ZUFs295assi1tPprdaDL8cDsWiL
m9Rp6eghKsV2P4zqkySVPeF8p6clZ6qeBkAVgsTizOSmcUfug/977JVresiuqYCFjhXs8XWmnukW
QF3VVS9xu/j8uPQVJdhr6H1igOISlko22hLZkt1J7c70OCsHOYdpefE5g79Hnvk50hhldd3g/Llj
h3iR8Pef9/pNthLEmcNppUrd0K48PzZsjdDxJtTgiKg5iwRlMTPiF4Tdqg8Psj9kRQP8fdd5xT1J
SvCXaa8r2WNAQCjenwjACc0AyPDtQ6uQNzAC2/Ir81vyvtpJBS+bjkUErdnFrMAs2OWMZ4H6gYOT
4eYKBJxTAenbRrnlQEHu2Zhq9Sz1cl/pnyEh1kEJ0djdXyC7vDOO41WN8xCtvGCTcrlVb5W+cc8K
nGrVq47S7eQcp9Ox1WY0K6bjffDnc/Z0WZBf6oTfme0zoE0Z1MNzqTMlI3dSkqxBcqWP2NqewanM
eWiwetxMnL/kjDdIDYBEmTj2RCNCZhQ1gyl4UPerRGSgHkpOdrHhyuP/YzJPdUtblokPiGPS+cGv
Zd7LIuWG8/KkCHBJBLIgba83yPU809ZIz/MGFjJSl7gHtA0DptN/62NPIqjKQMzZbmWtCslccKh9
pht1Amdr/83mZohucjrS9YBWt5jyjz4bCyC4Ecl+f8wOJTINMBzMwlDgbHIElaAOwErUnYwZJjHC
S6zbSKyx9HVslPrhCJXF8D+AcjY49Yqabb6bsAbOp//MEKQ456hrDcsaxFrOfMAZnOlf/JQrhD5y
PRmXBQWFfoL4jXxzpg+/SaTYg8ReCrVLww7jCNtTbt/E8XVMtl26xG2GdPubH/XH5mfTRv6fBXnZ
G3UWJjSYGcBLltW2px8WuZekqnUNy0+P9j7yA9PZNYrJya5o9mjz14stXE0dt8HbL+RZrgrj84lq
y02QR62eERJdoXXmSvbA8q0DKMT9Q6XW0y7y+n7hctnXGeOipCU3nFKNYi03biowLtbFwj1+poHm
LkBSdv3a7p0ro0qpd0k1k1y48Wp1UFZm0zitiaszZbALI+EfT97HbceHUha7J29w42IlBa9+a1Y/
9rOfTy70gh/VFd0eFWPS5LeEoUVJ+Q5+r8UfxMNgg4Ejhsru6Ou7eCiWZNTs4g9IOlSVO8ReFWOO
xSK6gPkySHqHxLDdSu343QV9GWRDGPtHJDW6aZR3xgI6pEjZhefZbrPf848n2c3lV0jsrVihM6fr
2nEq2be8a2xbeJP1TSYRrEwA3xHa1gqBzONjjebwg8XasfBz/zH0mKQfCvDeQJuaR/Zlp5zLhawH
sAOYdwZctNr5fsrO3+4qomXR/Zk/PfbLGWqvqHJqOOt/m2fSmUViQqnRrSUaxR2fm4EPqxwMUHBX
pvsvhqhKNwsZkMvTr6UFywHtUyZk0zRVkgqAZ/UwiFAYU5oQ2P4H7fNcs+FNGeKZOkH7uh1cikr2
A+FvkCb1mKCJoKkvyHKTgMozoeglIcmkXgDZoxkOK17Sp92gjq+ZvTPT8ELwJGMdVkhJ8bpUPoE0
1JbQaJSQr4UdzgrfZb13q/6x/lPfuYJRFYDVtM8l8B8X5fJo8GuYgT8dNHRAQa+04w7inCvNfras
9CIrIggA6Wles0zChwF6IZu+JsYoKmGE8xk1vSP2MqRw8yf6R037W2cRukf7nMgoGD9uOWtQw/zP
QhYhpBTXBBYhuM6iYHp5OD8n7c3BjeInEgM9zSUdbpXWde763DVpkq+oUgw2Hm29Eu0acvCT+kxM
/BtoMuecpupTcgNWKS7Os5BTt+0XQzYuLMx5wb77JUW/U2hvTx0TIR7hyL72/Zx7/BG/cztfJGKV
mISh9XuBzNpkvubPKAx9+lm4WOW3cjDmLfoX0+ZvgBY9itWwBcn5K+1fWVVHtGHLO2PLsGtYVa3z
QR96SktF1SfoSCbAvWvQ4Mzu8grZY2xjub6lQLvnoO9TSuj7G9qP+8zvGQmKYOfoChMCC/uxab7f
noDhpuLtq1jO4x248x+ZAc97/768RlrO02MwJsWrrAG3kvn+WF9IDalvbwEkvszL6ESmEg6Xpg2w
1OkgNrTRWjTlOkhrdDtjYEnmsK74T260t0YteSpSpvC3ho587wr+YlFjIa/2f5xSyDvy4klVg/yA
2WWprp3TyS5AGKHM08m1VOzFUhgGs/q3WFoq+7ANEGiuCK1HVV2EqVG4mHgsJ4ZEiHPEQ3tLy74i
SJpvPPPwIhSJq4Ycsu3ob8q7swixnPEU/vtCYJXSY8OBg2WLQ3BmlE6cdEOE5tvvQBVDQbiCQS4V
wqA285vY466JrSL9vpf37jAnVLcMz3O6xPtCMW0gg1A6LVeiTrLzTilPX7ioARFDb0Il2WvD5P3c
E6yf+xzSlLUS2CadKdwj06V/Bh/FOHgj/eM3jrBHfh/PbKwgKxM1fPTrFDd6YutkMebSPn+9zuaB
2hfTxCTGK5SIGTnZzyWCPGPrWHzmiQCA+SJY7aIdLRliAn72TgH3ruBrm+mLwbDaHypEVI9PINTz
CCw+uKUD2hgYnYZlMQPOlVOUvvr9ZBDa/5J/CbgDKkLrLG4zUwVvZMDNektsZmiUu3uPwHn6Zei5
IqTcY5ZGrezfb5sZijWmr5feFPke/eWZN/8jG/l3vQFDfE1n5PFuM8y8JbZ+593jtB49nDq0Ba6F
dQYWy1aqVrzofxZw9xwcFzL5vxJbujINXcjVhfJVEJfVvgApjTh0yNS5Fs4ZCnoIBp8KIXgPhfwv
EKwUxTfDcPwmpH2TGfP0TxphOxVjQuUfTsnwRMPDyTAsO0ri48HJqVpFsTl9UnTStiT7xiQsoxpw
xK4OvIawDiVPnbmGwhGxrzcCdYhnqlx8XWehnmN/Gpr/QEss1B41vdlr/sHzzhl/IOMGcFUcmJKs
sIHWPfv1sCOYCw2n5G6/LE9bir/6wmG/M3t5GNXshIRDpvW0Fy0398/4e4XcgYMyGaGIiFaCSHJ4
PbG0/OnSSOnuQLZ2ns6saHMZefKLuTWbIgxjQ4WD+FRUIVLe0QYF9a8D+9MzmSAXG3z1JmuDcYX6
99ARbACVWN9yfQX3CoBRrMQET/dN9ZvMkTZETYoqn2giCaAnlBNmPQpfEv4QDFx9bqmn4OjMK+Cr
7SZZd+ChTd+K4IYQH4xchPO/sqteS6w/EMmMQXLbL0uWtnMJSjE1mAdTlRqBcjPBPxV2fFsmCfWp
qAEEImMSlIa+bPXUYmuMe6qgpEGVleQqg3eMwSqqj+wMf+GUmpgFgWQ9U8PikrVbbU0tZQgW5yoE
Ibg7rbxb9ydy3VB0I00U1fg07lkG5UX1wxk/26Zebo970aT+xmnhLnUudKEvaqSyjlD+bd8x62U3
8Uf80TI3h7xPFyNrqc8BrTXSPzIOVtsqaSuDG6KOdwdYQKoHgaQD4wGm2PctyqgmFdi33povIhSb
wGlJ7ODEIL3jD93u20EnL1NK9sGcZTMiZbwJO+NrO/M/1yi9HLwcEF1o6o9pHOXUhtwrTJqpaw1K
H82CzKVRpuHcZarqZJeqpQq24IvNzdWPRnRp742VZUSxN+wdJ1kX7B74e7KR+gfUgO2fJTdDr1XO
kYCXcPYqplpJ+LyoQQ0zI7F474EJiAz4lTRo9U42c8DRKQkDC2ZX9rqR1xwDmXpFyLmRd2mw82Yi
TufDd6qxq07BwY4eNV2OUixlACo07Gw/emgsa7Hq7YfqWUvH9cFK0O+QiMy2qpN9Fd33PlDftqYX
n9HL3lSgXFc78h9MYm57lTtdcW90TmV0+ENT1NJCTCsYnl8qxNETZO4AMt1q1OXBHx5bC8sZRrsC
aeEyoUDOFW0+OM3Xj8M9GSEOyJQwQnEUZrdli2HlitBeFQOpUhU3oWtNFyysqhe9ntH7YBbOexMG
2J53BH/0rls5HGXQZTTIDyXwJKaNnGUpb0f7lH6ZMSfZo5PVON0Qk0DylsZ4cX13GKhnZ5XT1zEa
XNNFbksL5cT3EuFJG5YvMqz+hpDOnuDuoXKIpgcJrMP/spnbp6st1HcoWeOvkreANNgIt2ZuGyJM
2fwzN8pV8eN3pKeraBIiVtR9cCXFcE1JKuBVornncjKgcugFyHXFymKE5qIhPaOEkVhyp2jO/iOx
7UWHqvtLMhlttXtFVPj8V6NO0R+hi96QqDu27ZCVfTt3diomQdBQEzH7YePlHSPVRiEA3wxHgpr7
aCCcdqpO9/3VnEhy2ERn6+JquhwX9KEiZsBM23G2uZyuGVQVgaaLN/S9K6FfMOO++IhReX/usMdk
vtYWjEDBHEtKudYMw0JLnYC9KErh2r/8Uapb6jBhLSPy8iJDNoaGZ54EwdKR4Q/FhsU3LiEnwG4/
9UcG5HGaIeZomJBLLXzOavuRvKNy+L21xwBjcEy3PVybB4ik4OEJxVl0ebNWvKBfKGb8O7zwsGNG
tZRnLnjTcm2O0PDnZ8gRviJQep31OpmUVEDVffxAdd6fHpav3tqSXvvJOb58XZcinVAaSct6GgdR
Ku/aZMhD0ne9F9mmW+Du1Jn7oDUjnklatv/xiKbr6tmx5tsvh9Wt1zrapGLnPF4PUteDIYXwDByo
O4TXEGI2F3QsezAxtTx7lPt64r+1/nPLTdfJq8HcZIt6Tw+uUoMpv//uQcTcfOOe4npDJPDIlkkt
+AjY7+XQAiR7j9kG80fO2gwiFKh5/exlvmtOx3KiES2VigyUUriXF/GUExXL+42imm86+Hy87D+6
Q3etJo89x/YrUJDQuYMDvWf+ypFmZ/TOg13xaBwUqkA4/Gp5tVLtddCpuQbXRS0cM8xwFI5p/5ZI
LSDISassuq72qDTfDFiymK7ePGdMFHR59Tl0eEWfop9FdK0LhIYBZKltAjV2GwObePeYO/8s8YE4
cfF/YXLDday10fw787QwuwUO803eMS+VTOhHR84nKSAdKJr/CvCAj5IbO1q9Fpfx/D2iS6N3T8Cu
haxLbETT55tqspD3TfUhfXQSnDzU5Im/6JgJ3cdxtKYyBYuuWkwcBcOeCi0sRIp4vcrzQ81Yzuyd
7Bfy7GiNJ1zAL0/FPmG1SzRpcvNkAOfti2ZoWzMsGsOnhI0DFoF14Nlry4MbPF4GWth75M49hm6S
jIMq91GAcms6yT/8CZxsOHS+gQMqqpkwoVSFb/ec2ZgUv8LQ4Ytj9b6LZ6gTc8IwWP5LsJSSf2O6
E/D3Y+fEiYKZ/3YiQ0/t8LuzepYl7pq6RWyn20ujHbD3K32BOPJo4C4UxlmaPX3N+N2oG57bQ/kw
75R+RGawrV7UW3k8koD8A2gfBjvPa8NyoAsGpobCM71WSXoIRwMvQd5dIy8DxKoIWnracONJEuab
oqRh2N5UlqjdwhKjWew1Lw6K7n5daKGDXns9OkY92zPZAuKY4upKuXxCwLcLuT6Xy9aZCmKSQiuf
1WDmsq1hrPGCfp0sjJHQeVQrZz3LnZ3nc24UDj3z7SB/BkohOYRIK9x0Gxpr3BkSBKS2wdcSoZ9B
cGmncOY+3YZ20pt2VLEQQKgnDWfCBvNtccYXr03k1kPX+F9T6+UH5jgxBUlOu2OA49dh01WkJEPJ
sQKp6A8GkTuxVHpemnFLHekvS7IvDxTKBiM97PdGRI4vwSwbIzYGlfo8tiboXDFAl4DQ8q53lXxK
0bMVWoHMfr/9p7nrfjRWOEVUSvlK4DrrsRHB+qn37n5LAy4iBnA5eq/bLigPDIZ63KXGao96J01j
LxoTSwhNkKXhIDtB5oWMoAViyK88CaazE0VN56i/I1tinBOWuNElikb+pJGmzz/Hq7EiGV7cyn3n
a3U5WLjPv0EkiHaIGZ/8lGKhCZ6GQtz7OvEl3LmAQIqm3OfkmxePxNgu4czWUYHbmQdOGYthO2zU
pek7T4NioQFuapFNt/yEz4hBKm+1nTa5UpAkt84OXTzcMXl+LCrS/nuNm6X3Xj79QDkPwz9mTZQL
iUiw+bRs7cn7I0zYoWdsJn5a+O3lLhqChA81RSkAReDbs8FvaDlAA07KVnHpwucNFII4QLIaiqgg
Z4tS4WCsRgNMbjjoDbTXmmOd7lnL5FV7Ft7eh1yvukH57KcyS3t2QC+OWfE/TGEE5wyYhQSu2K8r
p9OkOucBQXxW5gqeQOfqG875jnw6Fys8l+lZ+AJs0UpQ9K7sJBh2V1cyZb33bzYSzxxSmESNyasJ
9T1OjVi/DQRxHn+LPKReab8H8Zpu9nHcHfRK+87sYWkypdIGhTVJaY32uvXzupVsw90Ma4uPKVss
mPh3b9QfqoPFBI5lcoxwEJx6c18BW7+pvFgQ6jxdgOqg3JL3bh+UPYapkCxj8SeAz2gyYmpWgeoZ
w1AyE3x0Sjg6592+CODynjJKnb1PXajiy7o1miw/uX6QFm4tcU3NoLg5haLo10zouUCKJMyMVksh
0mNEdlvTBXI6u6bU+62JLX41scEnivE0kdOJHL0zgPOoj55DR/g1vbGbv0k6L3lCHg2uL1yZ2Drw
Q7L06Vb2tR2KcO/V1426Fcp+fqjiOCwMEYeRaargURPlPdTNgvD2qGour4Q7ehNWs0X5ykCpQ88h
5ZOPyzMEmtGEFWfdqnCXK8kFmp0C/4ZYxD4Y6Izb4hFM/lf+AQlRwn/nkjVabWUyXD+e89hq+fJa
PNszDt2otUMwDJhIrfZLV1qWjykuevef3IIDzAiNbTOZz+Grvg9sk0A1JXQORnbVCKPmLhm7NXm/
X+lnqBKMFHmvvwqd7YtmTue2kNjY9bKZ1an+bOj1Ik0fPuzbHKuozaiLZ2Ana94J8GqhMVOsLXXx
TMMDcbhWW0lacZXjP5DsF2T5QRpMZUNjNwf5j4I/6pbRaB/C4eRP3eOY8AMr8faRW52SuVsHauFy
kUZ1e3ScPpAweXrM1g1oFB2/mZgEeCKBHmliKAhr2FVCf01We0Y/mHUJ7kmiELKsY4ozlPlbxbXB
6Kufvu75JIofPL94bwXmCRZghrc8FJJuBUofXwr3VQ+0p5eWK8COVMmBkJF6y5u4+fuQpiRFAt7C
7qGrSJo4cAluszZ8V4OQEhc6mzdYd2QvfJ06ppydqbvFgzwuJfkKtgBU7sJtlFVQYZ3V4PIOxC11
Iq8Ucqwa2Tf2U8wXH08hDewKd0aQQYv+vF2+oy+9Ch+wiATd56go1PwZgXZc+xxSVzSGcDm8nIOt
ox7JsxOfmFuN088J6ZphC0jZIe41bSStMT5Lyc4hTgjuAVK/KTSzgJvGm3dgZWmoKtmKCQVJYSbL
AnXkGKvVuUN55Wpmnlz7B6zqilaZ8HC2/KqKAetaCW4i3DLq/8EdVk52kC7X0vb3Y1i7wSPusL3a
o4IKxzw6nBlAI9b/3XDRTCmHT1hd0CkQrWW0wjBN/m6prmL5M7GHnPm73QrDRUhP3fvuEc2KBoOW
4Ux2gy2jjaxF+Hq8sy42XEH+M7+iBmMqf0qOK2n6Ge3KrDRzHRQuAPn59kZhQVsYylwBHNNUW7bO
gLl6hA+fXyY62/fWkhbBFIrZ/6mx+W0h7+zBUgJH1/EuRHUPtTYCGLRY6HQEDyjGapqDWZXXiRJ7
bAm2v+qknFAOOGRp25NDh4QCTboVH2LRVk95Jknn/1+JjmMjQNCEiiks6uz5KAY02G3Vsb2gjMV9
QiGbKW6Zmp55oSpJn+PGkfvB+aKB12ql/V5xTRSQt3WQNdCKi1n3OmYP+qGz7NFVsXN1qkLJafKm
YebiSGaeAG6t8AoCWdjjES0Bps4kxQEHrV7gCDzvBXnCvNrHGRzL7NmRp+c+FTxopVc5rLDwMyVA
7tijKvHafMh2HkEgdKt3gr1ylcDJBJyel4AzSEnXtbC5Tov1eOuLMdrAv6h7gpbRoW4zH8NqMW6i
n7ioqWeSHz+A7GY701FzPkmVXZ4ZY1ZSlhRrqN5uu2jneHTLN3FUiSDCIQvid1GKAOCW318EZbwo
vvGjWqFTP2lzoSNtw6z0HaTkPf0s8HHUJNoVTZHiI3dH+0tq/1FGrJfMF6RUVMzs/7tIw36bCFCz
lIkIT7GIrCawTkiCuhPbvTnPQ5VpGCX0cadBgZZEiyu5dK/mavkFtx1qTgh+qvqGKXoA2DOR6xNe
NYBap1nYPkCW6mbTJ/1/yQ0PhusY9Wouvj55OFRmsTfo0RAxeoPGXrHDdo/THh35h6Zlubri6TsJ
M88ZBeZfHCAk1PIzbrkILk/IfoV9MOfZnpRGXo9R1y/5NN5m36HKUAsmqk2gbi9z+qSnBKLUuL8W
W3jkYLGAXGgfBhOFObpNXnNEX2MaHZWm1oDxokjM55Esj2rI3PaO1qe67Ojhql0b25I1rzcyZHJu
GyTdsVcGyXSrh/afAeR7ERslp4ukpYkFOHSPruqt3nWHvFseKeoEcG+eRIdzDj2w7mkOjKDJzDrk
lskYn7FSUe70W4yqSfblfFcnlPZxgJguxVvRJm5PbQEjuZP+3PAYO0gmfq+hMNPqWL4LgtWOJsZe
yps6xzP0nmC+ho2qwam1dZQl2OzUjeJlbefQ4SBbCaRIpB8+kmfXtdaOGjThmYnNPYFrZUbN9MOy
ZBdLQys6+l2NGPk1QGmVBIxvddyAY9j6+Sz58KvvMEb+JNTP1nnzgkf6mDzpUTLTu/V0CSryoBd+
hX3ztlKNTiL24JbxYIBwbxUyD/yeYKyU5+jn31hhDAro21D5XIzeBoxHbJMsULFOWqBjKz/otMej
zjDhLkeiQgoE6lzCNEVr49Me9WIpndukPaq96NldVIeG0S9H+zf1U/MZEqOcIrs0kzyN1G/MssUI
qewa7EazcGt6KXEntcaMJvrcAVLSWLKbi1B3FdXV+B/BK2mWta6UfQCM8DpCznBNHN9q1sYQo6g5
BuDY3neRlxc3FnMFqQaFa8avT1GsS4OuMJiddx8oJXex1kmg+/GdLGhGX+1FYT/3D+bXH2Id7Ech
wlXP3lZTrsC5O4X2Q0XMbk4dUpl4hWqwPEBOXdeRm4gZ+siSkmhF/xXZMfDYf1uzHBYs2z1HMOSW
RT02iHjfZQQ5EjZflBXxz92cVOsrog8EYVO43DU58e2kFbDhKTS/7aJaNwDcJky3KaVfgZNbdpgy
hMOkXvCiFerWWSRcZsiiv1ltZkuq8yczh4sPQSX2HW+ZQXDGqpXt8HyQ8rebD0EbmeDRg+U4J1RU
VG6CZd/gj+D1b++XIkEE3obrMqg2MLAprMyWWZqcHzhLnEC8/Uu8aA4QDdRFhb6T0mT9IHna8GfD
Sj3xPwgTUqH0JllNpmaYJ3C+CsIQxBsAJ7U3tr5NU+b9ttY4yLcrseP9kFvf9MF6VJmnp/gd1Z1z
2SYmCbdqRzs04h/grJbcPYwbHQGWap/9se85axyGBRMQaI2e8Km2JQBUioXz2zzxnNpFubDKC3Yx
x8PF29/ga2Zdp1hUUMz7fM5H9u4VYhr27Y/7neUKGaXU/m0jXBTj8g2m6iUoWRsQJASICsAeWKmT
yh6TP3alCNQpA+7O0CD/x6jdeJfknwaipHqeHnbl99ZIx3ajn1g2EVm3ua0R0t2FHbErMGQkcooJ
+hIlVckFuxGqK2FzbYtO/te2D3YVYJ7ilnHXQIru2Xz+pK9W8Q18MI7jY17T5V3bCwytEenYu2yV
AJHw9xqBQ4aAhSWPJ83Hj3GqTg0f+VfF5xoxGaOpAKgWDicC1j6ZmH2ZiTkkAjV4xeCnXgOD6xcB
BgW6DkT3yUABPlafGMj2PiUsZ/f83CF9hOCV+LGl0GOy8tkJjcvsVUTPzeOU7lNr3F0kWWQ4vGI1
xGcrHm8MusgqCr4C1/e1IxycTxJgtjStmH3QX9CxEddNxUpMl1xmZ0yA6y8+iJjDTpOLXlDfgQOJ
s0s2aCpVlfqNRMW2t2qhYVU9THsrt2PVdwzd7eTYWLxlAUGYC90dK13fPIVkdPsyS9LDMLVdk1Cp
ftr76DocA3hCci1c1/O5mEnnnKY//3/8FKtMO5JXEVvdEgBE+uwyAaxK1nxLwuZWE5UBaLF8XkQ0
7wAKd209erGIJUZd7Q3oL0BzrSkWko4rpGtcw9b0Ay4nyxeCIBipOUQsNbiLZOVXGx2z7ZbE4M9g
xpsQE0TrVzp5UG6IAjv16RVCYawOATPKh0BjgtXLizPbRhSBMq77ApxmJEslem//8KevySu6BXJf
zJqzTZwgTV7OtpwJzohlgw+THmQgnOkX3ZtFEuQ0bz8OtdwAWzxm9C/m2GpMOGz0z8SC5ejwWrHK
XpeH+uczQqr++l4Z9E+eAUqhleExDF1g3HJWLSBNKhgdsqg8Uiitqn0CIq7MlctnSKgcKv+CVEA4
tPeKLG+7hgAq9eQGraq8zQ4cddZdkIr89GVUC0HYBdZTeJrdtweHnfrJxiwq1etUDjA4Lt9r/9MW
0YtsMuISu4yiHzHJTxPADqfDXR+M0vBb3Ex9JbRlmHJawXrld42mIBShNooeCszTESnob/weRLtW
cx6IIadMR1tTRVEnJdmSiyQbpTQJdr1oG8lzOTuJCefRKi6HJ3y5jh2W3/sugqE/2UGWtouUn48y
0MxjlagJHWYaeOGSE2VjuQMjHKK2LMgtlAyrCUKtdLHgGg9WfWuV9Egvf8a+ld9XRQbjX5vhs73C
zHfk5GOVpKvyQkUWfQf4n163jz/tz7y+FJwW3400w2eLIjKfvBsFVEAjgBV0MgLWf9WZdhvuNs0u
Jz2PljtBU6pt7veB29/kCZ+UfPnsdjU2iSZT886JxywVk217SX+2bH9M2pODebhGs8sFWz/GRAaE
HFUdjXvGXTSkuW0tc8rc73V7N225mF2b+dd+UabUJ6O0927tngBB9GuGhjQJC7a6zLvxEczsjvRr
ZIVzGhaNC3MqYdiygUCv85so+BXTTLj0DIvZh49KpPT98/n980R/6FY/wWRGxpBJP0NsxJ5pOf6r
Ti1MvuBi6uHqxewH20vCzO2zagWg104CtosYTnle6JAWKZX6k3w77ULHMycup7pxbw+wA6zySvz2
IlsACKpkX/G9KoTuL5q2mT7azmAjyd7Fqh9wdOYC//r6ZQX7Yqw/PVMiMpkhqiUy17OIB3fLNZyr
kEcEgZ/mYmTR1gejuD90cbh1p2QuD8j5T7If42BBKKCu3iXtGaBTR2wpLXCf9OAZw0cDOOfcmkQE
FswpvhNsA4F2nFsRfVISNTyoBXGb0GClvWKNk8DiggrT7ZQL5of6TvfD+YEYGTeXkdmsSo/JS9bJ
IWSz4MZpL2OOieBVlSd53/q1mEBiblCBeq+E0abuv2u3pTzEjue/qddWWSWuhklLEGcU6zdjKnU1
vMBy316HXIquX1xgdZBx5onAPakLHZg/JYVzY5ouum4Bdi0u0GN9JXEHsVj6ihNTBtkes++arKPz
2S6UCrSEtD/Me6U/tM7tid4WNPWeKN+iN1ip00Ek61Ga3ntbc8d7e6YED3KYazbtNOvfdGT4wX8S
p+sXTr0PV+rt+xTrJDRL81Eh31lnWUH8xPBefT6CGU9l82/5EAtCc1Wi54Iq0k6cDzKSAWlfq61E
f6slCTw40DHsNTV9X2wVnOiw5ZOzqz+GRq+k98a2psD3w8wnL57oweGWkQ0h+xzJFswmyxOZOAZ4
q8reZH6r2YY/EZ8L438deDlryzITnayABGIZ7yyNvWHowVDN7dO0xHBe4e+zkEwtaj5XiO5vQziF
u0C27OGe4yQM4jVUeHEWpv7pNtNXhuKqVNM72DUdRzW1kx2ybdmziS6YdyPEwjmCBNERFt1Fl/uc
MYK9ZW3oAVsC9bklqFSD0F5YzYvJBmTlNjekOtgU08H1AyJfODeweCXqZIDsJPAyZ7pbpxgvog6G
VCj1rQ8xK7mZy/lAkQSVK7XZyxlKwqiTlwQ7G19eNkA1NvKGXI7vjOEbh+1d9C150jaLrI/+kyPm
l6oWsgg0EWBIZn8uekrOhHlwauOQptxE2LF+8jorC/oMhrnvEQbbZPZFQ+V8YONmn5f2D22IVfTK
Jq98ICHirO2He2EOC/2Ff0C1Yvs9A4scoAvQypbLVaGyevIjPVI3nkAePuPcNCvYU5EX8V/Dv052
fGyi0XdXdMWC8TNaY1TE8CmPSrJNwOFCFCGBwOzEWqrfVPuAHPulAEDACTdD8iEcqPBR6zTpC+gv
gp+R9pUevfnN9W4WC+yH0d1YIUnVimL1XX2gYe1bkuAcqy0SZyp1qlohsne8JeW6br1+1ins9aaZ
3sqRmgHsj+brbvO7anu2EmiDTY/l6LoTQRlgJg5T8wAEC+gVEeYUGoh0R5uVXMtfecOfFCaTn8B8
rXs4imiBmFYgbByAN4DwWGQPb0BbZ/39H5VFoadX40tzARjO+iODJbmgrkw1wZflSTmY37YIB20d
a0CR/DLaah4RMJpm/aDQt/NC4fmaTHMy9O7k4lVt5SQ6FtkwtUoL1x4OwP+BqvSx8Y3ZapaR4Qns
rmlxZZMUet9nHRJiZSJteCUpMNJL7OWLdtx7luLMojB+ak51DNKD1NkNi9vGjlZ4wZ+jEYxar3ju
C/4YG7ytZDuGRv1eqgHzTOaEITEXjyoG37vHalyhya+HzlHjg/kPKf03KxuVv+BGRNg4UlFRR7sJ
kztJHVKkSgpMaZgm1gdlXwgEeCWJCiLRDJ6D1/zM3Hz05/IPJTejx6ZSfLMwGIA/xjFlPirhNzkw
OXYF2LBrLZ4QND8v832OE9fO2Eeltg8qEXCbOOVl70wHi5dmgV6Z52FdgBx7g6Dgtu302ZLXXQGv
wqLAefdGBIlZoiJS1ajygpPnyGxvL4Gs9UPUYgHFA4xj2un7MXCwbMNj4fDnsIfUsdX4kqf81cIC
zLq4/xUb+Gx4nFw+3ScBPtkgJ0UvaVrGiwwRLNSunvMbex7sDpPSrzJz6l5Wd9ommFjZerVkW8QX
aSDVzmi91e+XRJYfptodEVjaR/yxy6X7aWRP5IM1/bYZm+5oEmHhNLioTuwrrpvwSULsS076nh98
eEGT0qmE/nVJ0Px2mPVQsC3G6L2T8lKoE4to7i1M0pAS73WEscBmMfG3cKJbplp/o6ucHE/QlqcI
RwQizRq8kj37VPRN2tsUOd3P4DvD2kLKEtdPv1N7W0/I/Vu4ZK0z63+z8sG05iXaDFljxd/d4w6T
Mz6ySuGivG1aNycPm2rs/NZ/bO0UbQ5AsuiMAhC/La4qMWEB3j4ioLb6QQtG0LkGZT0LJ7LHvWCa
HK55Lw7K5lwt6CNsmQ4mxb0qg3n7p2WwgprHC9WaVpljd1OpkQ8PlNfPibAtjn+hk0ge0otOBAB2
7M44dgeKEzrePOiZjJXdEpJTgRb6F+JChQNwcq/JPB4h+uIhNRpdmMIVXOnYRoZk18N9c6mPYK/r
WVADIAiDoM8M2SyT8SuUS0YQyPfTNViVJ6+oxoznCWg5SqG1Dmz5CODcRvo7Upt8ULdrfUp3ZIkm
4A9PHYR3Ivf7rX9keEuUW+uI5rsu5pjJXpPaIuSO4fu0h3d8cVozE1IPOVnpNyDLQoSb0BCjY7zI
WYPOjQ9IZdsV+FbJYHJ9HSv+/STDq2yX6l5l/gZ0H/QqHGOhUTQhbbC2/mMVgnl2iDNmIMn9prGX
UCSjApEXbJSpg30H9p+5PB6mfqk4PGOwKOnhNI6HNWCRNMWi3zAKPyDUK/6UIHFBRn3RouSP5fwd
Gz27gBn1rsHwPQA57WVc2MHglWb0iyOwUvp6pkTyxpOUirm3jJsE34puXn4jso/fAI0jULEE6NoK
59AbUsx6RscvIM21K/jR46Z2L5PQAgqTh7PgZQ93OKY9Wnfs1rrRFn/w94bW6++kfvLskncM5IAU
1CNDewiZeJNNW+5SEBBy9D59rPP0LePj7ipgdomKwFGWrdtZN7X5l1XGaRLJtZJ2Q6wZootXJUyp
SZ7yiyxS/3SgMbU1QdsduFoEM6+NKEOv1k2uHBq1Y5ZsLVzXtTf2vINqWO1RdjBG8SHYrkTgw3Dp
/teot1NlnufVIkpkUObFLl7sZXnJNyj6UdZND6hx/VYG1GZMXTNIurVWfjP3HZQXZ6dkUhwYscJ7
XqL9TJih96KlniGle2K4oZ+A1/CCqglCOGBdp6kiKb84xZgB/P2je0bqWna/4hp/j2fc0q1hrZRo
t+u1Ine8PKEuaZrsxrsl4IJUgF5HElN/cxjdOtyJh2pzCM09ragDOaRs3R5K8jUExU6y+c/J4Ae+
B9pI0IDFcY6k3j5wHrh5pYr7tkDB/yuxYAeJ5WFU2bx05iTVsqqpQDS7ZlGqjcNF3+xFAr5+UTeo
rinRQtH7tCF3yP/ODMqS+nx/mOJGcqvjlNS+bBxUf9UX87R2LlYQj4G4sLV9Bs0WBN3VXaMqfvYv
uYO5OpOFxSBRAyZyGaRndHYMToOAp+BIXlO2CGSoNRGjrImIERfef3JeJF0WRADf2w6gt2Gsu4zb
smvW5W0b8G+2fb7bIVYTcBgk6gxqG7V5c7sdamQPum5gA9oDqupQs/6AHf23L3WAlfua4AQ0dSkn
WRhmoL08qo6tZHPBe5p7+Bn8iYLdWXKAQJi7JPEg/YahYSqjQls7ntceegFEqPFdVFs/SPV+ElVJ
G2PzqPayS0PagL26NhgkdYNVph5I2GlAcTpjvTxHUHklq02eTwE6/wFXwCN0iPm7Vl2Kja6Le/TS
uz79MWw/eBHeENyGr2HtdJEmrFmzZYtjS3XpIrREXLMKaetkO5c+hIl0hBW/cuB8R5P4hYMNIWrJ
BoHT94DvD4DQIHFnYjlcCUUm1ur/EPvrs9WM6jvayTrMcHl+/Uwr3p3UYOQnMB7rW+dK2h28MFje
q+yFBt0xYIR4gzsPgUxtq7DGdlIWFrwvu0FryUGizWEF7jJ/CZVxr3xreJHeTTmvuQyJP42zd5K3
B2OxxxdjILFw916aaUVY4L4i9RN+Y/1oOS0Tf5ZeySEBm8q9am/P6sYGXDuuZ6PQ+itHVxS2e9Nw
0yaKuu8aB0CtdOH7LlqijUqILCEa5uJ78Nk1PvO7nW5Ch/aNyQQkMHl9/pBV59g63kCPwDU9mG2c
HR+1S76WbztVFwKCMmzTGLwT0nPpo0IEV95mvfNvRaFotA7K4vQsjmaZ0mxxeqX6fvRJmM+onRcR
vMalVNuq0JcAsvJ7uuQ0tpbJdmimD4ijXqth1aHVc7I9uHKyFy4dWuCSH7bHHEiKegueboATVguQ
tauvttSUivR6ZLOsTYxCW1D60RwrTHyMFytuzxzTRcI9g0+qm9S0U/a8nCkIHYaS6yisJ1Q4joJm
9O1YBFndM3Th2Bp5QL6FuMw2X5Testahb8Q4QLDyhPp7FBe7+jNWIPa6phm1FihJMBR5c+OdVojZ
4YKDK9XoUtgwcAFzGOPR0j1eLw4HO0cyOs+n6SN5JFaQBKtUNdW0LStO71cyUab0wvYadB+3aSKw
i2x6/+1ExB1fVIX6XHEqHv5pF8zPnmcUY5RqBZ58S/Lw2grn7mJBzmXtG1mk10fHcyi9HXGlmJFV
XsMQ/dZNTiFf9Vye7bfuunfBOGgR+97qJ7rtvgNJy19BaZQut37UzGcdxL99DeMi9WjaOSRFv0VI
jffTYA+FmJ380IZCiXB+LIq40fwEWsFTjPMWDAk2je6d+46pyEpT38Q2Pw0f0sCFhJ08Fj3O1TNU
wG9c0WxMHmIjDgSqwbGPty4MdhfedxQxQjLSVIimnl04ZelGGqS0wyg5bQEaxC8gAd9Q4FfdQifI
jQzLflj47hQfJ7FQjpDjZGtLlJ12L5V7kbiOpCZnBQLeDA51MXTyfJ/GudJ2WbPOcyeiXs9w8kbF
as0nr1YG6pnh23bS8hspMC02N/SPrUrxP1IVABTaKBDCZuFQshEUvGRD6jfc0ZXfPmPVOZxXEeyX
kLYJmwLXi5XjfjyDaZxRyEA1oabEZr+lGkyZr0R0YtoHiMon8v9UBQXgu37geQGTbHBs5JEfqVOK
0UT1MjXbA0X+Q1Ja/mi4Vkr0rU10PeoI+YsACW5ncwr335QM/MSAJ3Zw7vmY0cqbCB4BGBTs0qD3
MZ5d+YkgV4OD82JcBVwAjxaS+18JZBIC6qkJi4URweVhRDIEvT9VCHy//YgC6eImTiHpUecmYfiA
ohr48u0wiZKSXWhVauLunJciL5hAXhLZfMgAxYjRsVLuamf+QcSdsqBabMRaxsebPcOi+orWaV1G
gq3o2W8tJbo/r7FMGBOZ72M5Y9oEWaf642rCt2B8T9pPv3hFtFaYA5gIjkrQh8wjC7qZQ1J5Szz1
sfB/1K71Mfy1uDE2y0ZNwe4j6z0fRrls15xJHA56+pXYolCAZRcg4qN+lU/5j8G6dpJNfoIaSCSe
bn/apXunUyc15PUBrYHwyOqD1Bvxlp3AHQdhC/kbACMoxRvKzj3yUpMOGDUhhItP8ck9tu4emSQn
FjOvGOvhFu6XnL5WMvCHUncyLr4ymzSEoX24++3Cm7hFQmwlNhfFUiLa2HJdE88sCXMMkvm5VjVB
IUzN6o+UJL2+oQPdYvAg98UCpUrexFgKOiM5GXCYhJGF9XVK7ZH3zBnRv1EUgbQ3Oeb0wi93oOqH
3PqIXF/RUej2HvGBmFehIuCfH9M9MSnyh5CnUDBs8HhqjsAwNBJd5UgLKcg1slHx4aws11Mw+dwt
Hajq7VZrHmywWbcMMYP5zFSSQBDXUFUApDZrJ67zewOu5+hYQGNixfDt0YcyF5GIO2mooW/6JTl7
m5P/o09omo9PFSW37prcOGdS0tMgxCeE7eUgo8+VEghRwUt3wmVdeIjA4xbrgHehsyKtKe9aQJZe
T4UOW7qCEj16z8OhAKr2j5MAxdlsTvRtYaTIQyMR6GymvAsbc9YM9m1k4x0Qd0P2y7SqqF0WjL+m
9fcY21z9zmCBipg7SyteaFY2faP1A1Lpu3SKzSzNDinecgrjqxwhVrGAgpZTS2ozD/6im4AYYnq+
9Jd27Fxr1vH24GYX1Gd98jBNbG3bP0q/79LgPLHrJEETyY08vcorBqoLV7dLLVVVhCQuTcNCJA+t
FhJE6wYiRCnvIVGWEVwyok88bjZ7f6Afen4mUIEjxIDmcDjYgYM34gEr900Q4QdO2Hv00dRqyaAF
sQtMr7VTnRRq7ihOa+cZPMFmJPIKdMBiD2FMqoZJMhGY5P5rD5S0RbFgdEQQ8pcPjs4gzRmZ9PyV
+xK2q5iajSLc9Nf+rJEqgl//UY31hNykli0uYP2hAWRIQOuxz4qdCN362qlWigPYnnnqtmbpTgYY
r0XBhllYqIg76KWVr1vsjkTvJ0ngjRdGDHXkwdgmYsb4VGod+oo1Uc2ms8Uj5zM8mSWOgzzTnW3y
CO+ccrDQqqpWEr/J9NOkigE/sSoIVykYUMff39m8FOvSltTXh03ogxiG8j+8Gzu8CfM+tZRjfzjV
CV2sjxw+E1Ia4/FgkUKCWm3DAIV9rzC9TgxLKd4vnf8/p+TYIVXSFr8uIlzVf9hi9zAzUOVndXXR
PY2JFy5jAPTgisOyfEtad+8m3fVN7MskwlppIYjmt1Q9AjeMd9hA2jg9MtrxNbgU0pAwYxs+cSlp
vaNsVkPYd78X2bV8xSrImFnpvBtqsO3jll7T6Z3mc/vzoywKVFSxm8MSoCS5ndmQDkATWKjg/xiE
xTxV5qmWlmF9KOrYSUOzzJ1xIOHCr97QOtUOVQux2u4Tl1WWmebLHTOzrDxvt0PUV5AjsS1qM4Ir
SSPPFWmwwxRdTRGaCCfCjqxEaKeOn+wBv/QT1JSj3PDwh5sRQ5trrk9uErGCwNvO3Zdval7CJRzB
bi6/cV5rKmO9U/Xa6cLoSOvYDwS2ojImm9+7TTOjDCaeZR6dK2kEXTdj0b5OrGB4zKrjEvwIkiTL
M7gqZgy214xdqCLX0W1hTEcg/H9xs0EsmrdSzQEjL5DEwOr7yX4YaixSoBbmfgmvYJIf+1ZREmw8
xGvW75q1ZAqU/MK/68g/75BLjwyKQf+9w84SqoPCGGZV5uSxuX+UeaJVjfNwxGu3yVx5LDhhJJWa
6XC/j4tojKs8OyGeH98kZMG7nnPcHCnQRJ3QMbd8PEnjQgC8Zg5nC8yNkH1J1+1CHiUPxCqPwRnP
GMyIPtfD9LfqI6YgnVb38ZdpdDMvOhh3hvdHu2DYZkVaVzVvk06CzGPyQwyBuBhNWqx0R3louyva
4vDkrqkDXGLyivboVy6KF30+Zes31TuaBdxT02rdJTGmrh1YOnIt3T3C8PrORlTTW7JHTW8r3nIE
lbPYeJTmxihRSgGxQS5lqDtP0j+G0xD22WlAS+P18U8Vgb3vFEp6wR2XnqZZojYFRrWCCboUsFSD
x7CQxLskNSmGtSqCrDFQYk3O+HcISrbJM6snikOyPjz+hJW0NeNobCP5+l0h1J5Wuc1K1QyaBoQl
T98NAA8azvlhXorP3pyKQ4w/xSkNrmBPxgQv72qAXw/vK39QkWiqOjEK5OqVcv+pf0HeKxyfm1Gx
bg2+k4zaYLIGB5yztbTcpQIUT9wlRO2ffwJaP/3TzgJhRg3tkfEtmFTmevb/nwQTuCN2YsgQhj+H
KxlgAmKSei+tym6UvYyGYsqb/jAT/b3NEqRNmKkqWxUOwvmw5oQvksMlH633s3v6ZYe7kLgfa9eT
3apVviAOrY3PbJPeFrG3Uu/q5G22Nh31o0DPUFVzp9D82kHGtKcUGnsbo5gQ3qdX53gD7K7+Keqy
TC0JtHC0j86rHj3UDXr6k9DXBtNr/6RT0qlmJe9XpGUcfMFDI/MQ4lTZQfVhp4bq9DHmueGE2xlC
AgYyGI5uS847mObsaCXg7UrfQLXFXtJfDhaHXZ4F9Ev9w7G1UdKPDVjltD6N0RlWN7Gj2DM9ktkg
ck7uGZQyCVeR/72w44hYyU113XiJ3ISPZqfaGp4sPeA+Q8qhHc3t6EubXiyhcquNw3YbqhFaFu+l
KyNLVwrgXNLSmXmn07RAgEdDioAhttRHLvDymjA0E877yutIZKTDfAJUWv6MShj19re+QsREtVYJ
o1Rxk7ocVWMyO4JMJz0bZqgbGTQND/FPeVW3PD9exwm26Ea4PdFM3ZonPzteqvM5Kt6iT5kOW0qF
DmkCCB6Dz6Rx6KzlF5/9s43NYkbbQncoNz8HpE38JMDsW2OeBhQLx7f7NL1+5L9ktph35aqYS3Mr
056a+Ms6JyaJUAe0km+5MiAPSeY9sXzSAe6ifyrbsN77TJYr2ppSarE1FpsN2D93R6z5Vh4JGobs
gg7ZASo2mVy54SFD6D7Osm5W/6Q9JzvpfmKiibCInwtkjpRbAjPFDibLma/xkvStBUaHdOEiqdlL
WXoATlr62N28LtXbuY6BUOtDVwCV7vaoyM/qXtRH5Tu/iyeE1X9sn6PjFiuUdaVdnwkJ4r+VBTkN
fB2AOuRSecTBEDjZAk/6LUD1bxrO5pAEpWqwStGWuLXnjka+xFWczPozZGYSgd1ZJroy0wXD6U7k
YGnanhudp0lf2sKMRVVahlWQjeU1nd1tD9koVmLA5lvoKxesZa6xzmPNlttfG2QNq2POuPoNPxgE
0n+ucmnOfGWxhuZPYxtLOiUJuuj8RmNoIQxDCI8u0ICeV4xzl4jEzNdxByvv+M7N6/cE8hEUCixM
5uuF3VlhzuVfoAqFubSHTQ0vr0uOW5OEID4Ro8D5TLxPoHyYSj/LCPZHbfxkpPPJMFum6pYl3v9o
PyQnCFaLcspAuP54lDTxFwHGqSj6IgygiG1QMInKnwgFBbWiJiPokVFqd1EdTZ9kFkc9iPsZKU2M
s7wa98EvcsJi0n3eoqQ7VWQ4F0fCRglJigy1m67r8SgxTfhBvxundVfpBhv7AkUWhAKCQBDigpEY
P5vEzI9XbYI6fXrnOre36K6nWHpHGxtY/htnfj1tzESn6kw7MrGue4FY3jBrJxcN1Ibbhcanfcvf
3hEvP6O5eAoEd2J8BqQUIlitumq91O6X/HXV+MnOv2M1QEecdSLee7jx9t0z9KyQjIeGOvmHlW5J
Ez/Il/Ql5iRQ46s3HvVmebJz7AzdJk37rStwX1sZCLoa63WWD6I44eYNFtk1eq5hUKXKdB145YrZ
SrOIVatlUq1U61eMGgJ87w9a6hw0eF/zG0SWELlIrYRHQKqnGS9HWM3z+iPYJq/Z8vYUOdOflK9O
0AW4jwIvlzr+QzAXnHIWOuTYhRQhRGp5CwBZH8TNsyR20JammlKl3ZJ1dAZHwy1WXTC5mbOmez67
CQFXvpkuQtGjty9LWPf+BdtxPr1N3njvS3av1KFPCd+T819vem42WDDkeeyD9rcRS11J3pPn4tDN
ot2gIooDHiFFU0fJ+J8+FAIT1ohixh12dtduKRQd8jltsXD4V1OLib7R9QT4IIkGUnDpV8OKakDI
usQv1t1wJadhkgj4WYPOoi1hFtPY5rn7qGkY/c0ht9Wb1aW/7fqJsw98tH8tbt6xRFLTbt2HYw1G
m1kiWXDUml/5qzuIWM9UqgHBgo3CJpguHtATzAZsGa+MI7Kjtq/EA/g104k21AzsdY0bWWa/cqtc
U6rvw7iNc4c0gEOOoH9VGz9IC8tswAZWFkWANhkpMVHbUoPhGcid/VEuuDmrnfnSZOXEvU+4lZEk
7+7QGwqw11/+xtN4IDpsYjHwh2nUGbOBCEjuQYSfvAZ9Cc2si7JSkSfGDkpOyCkIAk/r3OlmgQjF
jgYZugo2HI+lsQHKY8Btcvb7XrP0+l612qxOub8W9qMoOEo1ecFWnYQ/usMOPBd1rGCFwvVeVTcK
2NKuJjwDjQTqM4Dq0MH8I1qlzrbSMCzzHODoJAqBMcm96bBVPhFliyTXkKL4zi0UTC4Q5gr2hw0z
vquKMA4PcLoGLUSd6+RWWZajeXePCuSwA9tKKKrcdxiQV/SiEx/m9gK+zE1zQ4D0+W/LxPwRE50K
z1ZTa40yAeHXS+tYCtIiEl4R82MBWnHxJuJX+Tf8HYDNdk0K1Fmik2LddIFGT3YJpCHu/YDABKe/
3fekQe3PkZvu/fhNoeopAHZULrHTG/vtE0dIkA8NYDa4NzcS2N1j9AZb1ANDKN1B1jUcMqMIjg9I
JOUF6wTx4TiIFe5YJy669Yr+pu02apCQRbXBJEV2ELaeh0dcHweXu2Uty3PsXS11/I9yZfdpqILq
3zqn1ui7OvJh1UYofXWGR1CZaSVg3v38KbOI5imwNLT9iC5+0w2GFjJ1W+shs3oa/Bng3vKCnbvz
pulnkeamyZ66pGUDLYjtfT4Zg6KBp5Y8O88qELWRuDkNXuxG0c2k4A9ST1MkcXy8ldpUnRYIy52A
1CKQwrLKC49or4LpDjgjsv1O1oSqmMrdUIOEPhzygvZtkdolujyjiUp75xNCaNxDndmLcbL5SE5D
Xlv78oYcLAx/JE+SmMtACOjT6kz8hftaKzFFLdry65iXumwPVCvyidvazfPsThQX2qnqFrL7ya5j
r3Vs3po+F+GoLwEY7oDGExm+s29n9mldgx4eaJDEF9uR6O0kQBPLlaDg9tbgBc9piL2v2PMBRFUN
LX14HoGgO5NgaE+ZMgwMcVEYHBynAtqpautgJultgUbHc9Z9V5F828NaNAeyiXJqWjazea8t+g0C
1UG32BhrgHiLRN/dvhNL1vpW6abckEsQ39N5cmozJgT38Zrhd+S6vUMQaJy3+skhZJS11gIf7nT9
W4qKhhfudVei1X3s1zrPfJnn+FEXRLA8KW0W58MfW1kZ3bEIUVTyYq8wV4+JwJsbd12K4WXTOW3a
zz7WD+j5huBATlNRCdPowmu3C01UwbIqDzSuwfoJVFywbsPA5umYfzFBmtRs13nZz9L1U96REWJX
21EvhxpL2uNbVlgBQAsC1W+CY6PsZ5pSJgghpzP1Q4SMDW10qDvbJnzcZvsAB/xBfK8L7N8odM14
dQ7cY4brwty3N8agreBKr1AY7sT9pqzLI+GsGH1AjOwn890nc6LPqdivRR+xSNk+fPkxE5qJpfyD
SC6it03WokrQd2xNI0P+qiJE/SK3swStyqc3wpR0+LBqKTNBAjIl8wmZZqquO7BYPDPMlPT1jOq3
TUUmECkikfbFDIZKosqn4p57MQrbv9nvYjyNqBduBEuOi4ReJgDUgALF5DU00wlu9F0D2lHO48CO
kbDF4VvkdwAb/mHz35LO8YfwWf0lmHP+6DGrQ+F2wi8x90Md7SmW2edXRtu/h7guHluES+p4dkwi
zvU3epCPLStfk4PdzBa0BpvavTg/Rr6nqkEGUHUhciWUThKezREOtw+ojFEUKc0bD0QHNgA3vZT2
BpKOXTAUBPEQglNoy3TltEp6UyGXWlXVe9lEV54alFzUHhiWDD4/hz8jv2wRYSuEt8vvppFqKXUH
eZNfROysyy4bV4kG7TE7MREx6rqOMErhewV6WJThSnIPYB1+gRTY5src5TVHiZDbM6SkIpyj+hc9
z8VDk4xKNSU7AHwn1X/lGPR10yTH+htGZI+S3aMIsTINeMlKIx4gd5eezUgFFMgN0YLc4x1t6C5L
1iejDViXKl80Cu31uT9RknHwSO9thYRWv5xvr6mxzjNf+45XmGZ29NkZb1BngLUxEumZLD4MQax/
02U8EcDS/FnZ00SDNomBvuwdAKcBxhnWwJidAxmmj7x7LUN7TtdmsLEgPcK9wj/IbfTTg3pMol1Z
OEVSaZ5GzBjhyvuRAZFp4AE1IBS86rkG8ZD+Mcs+reve+vFljdYw6BiVJ0sXOEKEXDSR548SLCPt
RujD1RyHqqePapNVI8sY1F3CD0Q5j8VggwgY0UhlZF95pfeTngaFVjCg67aV1sMJnZRi2dTyw11y
FJcLWfoxI4G4MX6RLpT+y2p5Y6tgoYaMSYEPyFOhVGcd/F6rBli6XQX90/MuekXZ/smokiErvRZa
GnhK/bLT25AAhTUNTeyfVhx+FPm5SSrE+nZAy8F/7mK1y/jLuIRV3LQtZ/GPbjNZFWgY2jjIuLiz
qCEIJLDOS6gBZSE0RM+RLIKI5uQeKB+PD8UC7JSCNvYxPyktIxxVOOB5AWxlruOklYGd/UxteIqK
YOQMWrPMVDSfRj7Io1Kp0T68e3xnI3sOLDjEdvvPICH/2gyELyZdkfd1jBSAvbFN+iUX/L7GgR0S
mSUWXC8flUpTqFPN6h+ULFRPEaxaIDHoMXHW61/Xc7myJCmIClo6Wa6dpnkRv7II1U/JtfAJ6O1J
pyVJwRTIDGvqRghgYKcEg0Lcx2V9OjillibOUlo0M2ythYvgNK1dfq90VrNVpYPJp2dPb+98M1Me
WF/OPWiTjb7fr/oZaULv6zZevZxc0ANddOR4scmSfGE4tPOG5YsUnXbIg2Qg0RzQt8cRQHKzRF1t
X7oiQE3ZAk3fUT5wwaLA/uYpHgh8ic+kQmhWXpuYb2oCqqjCosGCSn2bQKdRip8JFrdtjYK0V9xS
KVYThGvYmH4riRKGS98wEEstpno9mLhRcQZv7gFCAmwclw+leicax4LIZstkpMSnHPcQSnK6fjSM
E4W2RIfNOvzVWELBpYsSiDMq6bZrftmxCz3X8822NwgpLle+TdrDDHmbXIxg9gyabyDt4FQItMPA
UsR9MM+6b3hGOW6aRE2wt1y1WlbKfM2jyQcjl2Fl2Esx/0Wx5mJNdjEaff4H62NIu/LVKF28tWlw
KhcL1SzdtWcEF8BnnCulWI4H5C7CQl+JGegyrtxavPPFr8MZhlygg4pbLxc1o+0Jx7Mse904WgjP
Y4amt7LoIbRbZ/MwI0UBxvGhUmQtvKx68b8HCzp8CyrMivgIXBNyc0EavszuPzyBO8eDXwgAn7Fv
pJazhcZerPQEHMIf02WsTk9QxnyG7xW4Jn5E10Leo2Akr/aTeAeuRvLHoIhwkgr5MTOz3zpiYtT3
fRIeyih8OQW+kQoFoWbbrmKXoJKgrHdUZX9h02jTM4YmVGDvziyjClMKATEybVjFIu9j9T76UAHD
/86U0AiwuNHcK3tdas8mJCaWjXrJPei2wxmIaI5EjQWuTCEqQEasbvNezJVrndJToaB8xkrdmlQh
pc+m1q8OEwgkRXCTEQjQc3/yUPupNmE3rXDUReer0EBgDUs/Akc2rmvOulAbnhGt2P3166gRhA3h
Ej1SeLNuh7bBDIDqSzoZTQy7f8w73A/8RduhxevqZYzbD+eZ7PPPrA8Nc4KOppby75PBIuMDqNik
sNcdLS1TZjEQeGe3sI1AGXjeUNNc6P0K5sN6g3qDLzTJWs9ZBvH6rB0QbGX0eKxdd7jqEUZ3mAKO
Y9cfm3sxPflqbNrFqY+14RAEz1oK6UXVPl8S30xTv2ye/fij6xpGQViaUM5O8jgaYN5AgtrRohfj
xX6w8BEmyCRD5hLEv/+w+KrG9D0WRuw3rZh5ygbKI0vHcnylC7JdkcPsMsyHzTmCrPM/Y6Qykdc1
VlSA9tB5FmDGIKgftqX/85ofuzx7Q2dHmnCzfSeJ5SuTYXqrALqIg9Dg1UcZN61OTUVDXINLzI0O
99TtDk6RBQH1zxk972bAF/HI9mZtHyzmnMuINxNYvmmTDcwxhLdYz+fLGKaZZPA1PMpz2Zu02Sqo
H859gxYe6OZFZ8/DRVkNxHZ5uV3h2JW5qsQ7NZTiTHDHDQilRmCT0/Sv9VJ4IB+P6uT8xZpjMy6h
QPFl574+hz6BykF10+NFSAl7K3tpwJ8nxYN3uWikim6rL+lGi+19Alzl5OIc0NH/Z1sQ9q2zBRYY
Sv+ow0D71PQgPO9ZuG05KNXifYNmc85IIDMWtXg0L8l71IeFLHDiWpxfH6o5/Ma0usW/ALeincSP
Qxx4HK5xhSuwnY8mr2VVNP+q4dw2wOHP3TqpwKIRIO9mqiokUnKRYUoED/HYob4zJzHV18MY4KLz
kxVoMtBjpWIhOXFGXQ7FZ9vnkJhYhLYr+CSrXaLMkRLCzVx6DAwapXRioWivdtqTU/NEfA1IWY0r
t1E5y2pKBtY7uXeIrVHvoXtaBYqazYGZRN8X6MLIsEdP1XdQVgTyofUyAQWz5LNxDjs2CK5iolfp
ROfF6nt3DO8F03aLHgCT44DrJc1m9coiXOOFwkSbdkW/OZRp5LUBiOvzza2oeqzLzT5h4AMnp4CX
3GF2ufFSXybV5LoXKKgRMzgppaWZdnjDGaZH2ooNnPhc2EapR9ePkYXILOOmom2TZXe2QgaFSqc1
DWq91C/2+6dndtzNnk/yGGUb8pKhTJHDOaIYEqZ3tTUvasON51a9iSFsPOTSiRm7YJFg4hUvJ0t1
3HeP5z8TgppuVUT0yk5CDA5NiuNyUV7+bl+aTWtl+QTc9M65ZtL3niUHyOkCFoaDzS7tdKtwX5Il
D/App0IpiXqKJh89uLvnFmxPIhB2VUvW0Av8ihlHmlmLMHvU4HqUAqp58fLsvX+l1ptJhHeW13Sd
tMJIF1KQl59bSaSmYdg7aVyC8mfsS7mRVkpSKXPr+KizZoTBkJ6oF/A2hl0Trs2yMcGftGLrCFFf
DE5xWJpZTDGqwyMcNibQe1BLgGR0Hp5S6GnsOiji5LD2pE2U/rgttSS8Alo6+YntTUxMfI85oa59
bjA29cX9JbMko/6nsU55g7yBaR/vUyvjBO6ivN5mQk8i6ekmObnxP4Qr9GpQ5GKW3/stSKnlWBkz
7xoPMifzE1RzcKoxpriuQGkjA48HwlU6MT0qklA+MvsM6k2kM6Ek5S/Tw7+FJecsLUMG1ELe/l6J
DYN0sWFQ/gA58Xe5G8ywHLsl12N5dHDQpYKSMTMXxivPlkoHld1CuDO7E7rStX+XuHi1mSdCuEQE
ESSAP2zH3gGVyydcD888f3XWuPvWXWXfnHa8XhrwRzrWRzXeR796URlWs/woc567jkJBSly6XU4f
u5QApJNAD+C6d3VjqAgIPv5YHGZN1BsH5tlrRxgSCOA4MClPdqocL+V+8TZvd/PL5xAHDbWiVCXG
3dveHqq4+cG0TlGEuYIXHHkwUiVjjswRLR4wJsdtPJH6REIZnyeGjLDh3tX7dqt9PBwOeLzjHepl
U36mnZPrIixobbCkhFVdZNmTkwe2Yetr5glnCoaGgcnKV0qyZX1n/NDQSN1VhmpfrH07o4FuElS1
H1EJfMBlTpRM+P79nL69hKIqDqTad/FzS51B46WBplnp9T5O+ujZhJSHgwXnlYGdH8YfFh/NBQz9
l48q9rgupM/jm0wqX7i0+d78rTQOJ5s9cAcDq1OR7JbZLGN6NuKoHUGTNrFZeDoZxHy9j+azx9OE
Kl7nR/d5UOV7PCumEMOWaozJa1NAmGzbvvstAzCP2s2gfhnB8GQdmGxFKs9ogIkC4c34QrdRPKRE
mwYccEWjt0hAHZqUQ7mw3WfXM5L3EPIOUVolNxi/q0jyKfoYr66ZJOgQz6YTul8lbMhR1qibt6n3
+QFlYUbs1d2ekETBVqgbgBI1bn6JpvzjyOa5net4W+jYxnYyjViPutWGC/PHXjJwafeV1QMF5qnr
4flC3z4G94BdhvR2Aygczy3fGQDbfEKzpr/jAsCEGf08xuUCFAKwCvX33Mn9QLodqwMdqbq9P7k7
W7FyvOzrLNAZg0bTpdZXfZ7xvsYiqckq9+FF58XD1aTY5qadCL3fdO5nkkbK6SgpUJ/oQ55FAv99
OGycnH4blfLqa3WMObgQc6WRTLij7EpmhqLGJYlPu3B9CSYyoUMcWm2yx9bg+LAqUva17wDUcRax
NnDIl0QwKY+oacxja2TZKA/KTMBDzqdZ47oRoq+AnEKdKj0DKOMXwxLaGMsxAr4prUpK3l/eiWHt
2MmNZqSe+pG58C/yOGSZ0lzrhpy4NSfob/1/B8omDfigdHUGdHjJ51dhfQ/Q5Fh+l9WQ0mbBBmdt
PcPWzub8UStIK4ARt26tFMWHtpadm9rRTvEZIWaX5KrrHtEczW5Xu6w5RV1dGTPs5mo2J3WFe6mb
JyuDnkcNZlnf581kHaXO/wtT3Qcqf2w4CrATCJl55dFuy96xbaEjCCj1uNF89kqZ1BGs29gpfKcw
p7E3SzM+Me0NNuKkLu3mYEoCOwdoMhqrOUELkA6h7TKvSY3xR0VkyL08kXJ7HYVe9HIIlVSrVNQV
QALIQsze3JJagByHLJG2DwHM7DRFyaARxSMRLXb0LECUxBCjnCPxfthQGnD5s0dgHpA4yYv6EBPt
MhaQxaIpjWd5wgySeTNjmxm+3+kgEvHPAKcjW+SDqLBhYHaQzVV80DFri0xIARwiRO6Myp3Q8K9n
8tRkKN4M+RM9Q2aCPsJfNdDokrUpzlPKN0aLmEy1W1JEib+lWIerQyXkemLwGfoWJHm24Z1vRC7C
PZpC1UHVs5ss490Fvsr3Px9fxRTZEHdiDs+wZqimBXmxllYwpkBf5pFgwlWee0avoYy8cQhZ3Wpw
hkAynk7Q6cwdV8hVNLBWFydTzaPME/L8q/cIT4daG0XjCgVQCfigwPTkKg0w7U/1L9qyOybdFm5M
5gqUth6VLyr30z0ouYEolundGzsmtvIV0zpQmPJ4OVZAaWGESR8k2AaU9qbAmoTW2/xdwAWsXV7p
ihBaLoO64xPDI6bdtZS7axK/K+yvIqeuHjemrWt4lA0EUcmX1DVv4LYNm/kZ8tqVvfR1W2hb9UK3
jPRbkEh6B+O3h++ETJ54pgDzrCBdBbY8Apd52sYXtvZD8fU1w4kTprgdVe39N+DNGsfBvWrl7sGF
LzVn+sVuCuxgIAKFSD7CkGi+o0xtWV60Ip/9frHTaq3bQc5CWyEBd2OIYoq9NGSV0JwFN/7spbGh
9IVKhEHqdqG1/Ly8MS6Wp9BqI29j2l2XsnAIwR/yjJqt1ksSS0o+ji9ye4lv7Eot3D+UcoiKJZgM
nv9qApaBEBAv28+G9XiK5iadI7PwbC0xyDszbukzb3ZHHqdFaC2+zeqoBZjpi8F9PMNWzWcczfd+
jqN4qdSks6iu6uIwx/9OQ5SS/ywiHbFgTQvJpBsTdeMh4aBYr5Ufw4O6an6FyNgK65BrnU8Ey2wi
i6BC0nIjtiu4iKx/P2cZh3nzr/9n+incTb72ezayXvJ3Lb2rdJwNnSzG1RyBe4Tra7Wmm2aPbwLd
yZO6Ro9AYTrQBczdXqxHssRAmwfkHOYQp38kTvXhISoK6jErSGz2LjF2LLGIheqLQe7xYDk+N/XA
KWgt9uGqDSvyr0kEItBOjC8qXQiy/oF994DijrI3NakQpio2tj/QLrBgfoFgKoOXwBF+XN5AkPtm
F7MrzQIgc2MlUmYP6diNstHPdenEW3+mierg0zRwdRMmWimE07Gnd09V5Ucv1RqKNOa6FWgsujoV
SUH7Jv3uEDBC2oj3LdmqNLXpDlLEzrcRj4XnmEuNFLXpq7jqOrGBE0jSfz5bWJLNTDflC0Vzwm6v
LDGiKUaCQ4yXVByNW5NmOzdeIxGgXSHURB45zWG+zVyzsuYkFXF6tORfFM85V8m8jaumPLtDofSO
V1FPDGVoyxzXZSCUk6bfARMCWG+3kW9Yo/juJiTUWWnQGpfTtysU//pcxPcs+lvCAHXtl/e3dF+0
68Z8LTjYKirii3tl0tw0ruArjBKcWisp65/5mrO0Rs3XI/YYpxyjeMM1hfZkMkfQYI3CIQaJ3eB8
q9CzErM8xC01UfIcvVje8N50/jF2iS/ctXJIqnG/kLirNpVKejG0r4t869xQUbGQIb+9r/WRQlUb
+Gt26UUsa5PIekWcQYaiSpLDXVZpYsfidP5eybm6jEhBO0EOJo9FVUoXnLwgIB7HDTOCkhNLur9/
8Z59UEvncG29aqKx6fAknyo2dYbBvo8R7Jk16hJp0OBW7bdjula+AXwK/RgqJsG7/I41leZeQqm6
FfmBvnf1KRfayPVSmmg4MERsn0SYSDfl7WtpqWuBrLj+Yd+L8755SoZUZ/GciyRkcsaZSZh9VC37
J9cl6oQlL/9uQ697tHXVRfhwFOIxzsU0P4Wex0w7BIQ1ey/RNP3eA3PEa5f05cwZZOCWbub7Dkax
PGwHM7xULDjdqSSc+uzXHZWwsdNuyudYJxBAugzxXjxPl38J8+umg3RiShKo54T6+SFkY65xyz9B
gi5x7isBzofK1drLVVhIlZ6Ds8FBE3GjuiXm3X4AteXpQyJDhyK41KnZJWlsz3xN5Qs7KTToD2zT
qsQUFEOOmdo+xS4eLilSxK7cuPFclqEXfInTJxoujOtBaZmhexxuDZvx7KielJCBMbW257BQxJBP
/UpwBhEySiYWidUwptbowjJpcXL0TehLdttxF/hmLUJOPIozKUvxJsoOjoXTc2lUWcLwGc8vnV6c
VjrRZuibv6WG4kO0uYVLCYLy0EPMiJMSORqkiScjnS7Dl2ymTQCjaccG/pW3e90YHebUKCPdKQ2P
2Nc7G3sHhhyW54TVHjHMNpVkpumn2Lwv0XBdIdxypEhrofyQero/fbnELikcWE4QqKvYiZJ1E8TB
+G7BRE6XP3Sx5rHnel5nc446l5zx+yb9L2H4N80mONy9Gj85gxy1qq1mLTmwlNdg7XDNPPX8HpV0
oUKYa8908IpuWDZFDeKOr5mB1I9D2GEIEW2k5bbsGdiQiiSIz5nYm32a4WD+j1qlkObGW4NrR5b3
Jv+vcgH42Ido2aWyheNOb4ipEpsfdnolEBDYMIP9xlP9A0QRriBcRsRxC/o4Cc0PgaF5PfvNYum+
rm5ykpkvgiEzaS6kUd8nGlRABIDdkpedA+6gCOWjV7YJgiGMdl7ffyXgnSANAGpHfUPWXSr1Cl06
1bqbPmwwqKIdWBayp9myKMK9y0m0CFRRXpUst2K3JAXiPI3/kty7ZMBpaayi9ZMjGIJoIqQrlEph
XSY1xBYtJ1mdbr5KAVA2W0sFWOVPbK09Lxu9UW8c5L02a1DwtqNIWw70jpG8JA2ky0Cr1Ncw/CX+
9XCRshSxAHN3EyyygX3BvpqR40pNtOXePQMdKcbmgrjlZOxXC0VgwwpwvNksT2PXnhiSIcjSzorI
CejDYDqZLqUyvXpT1Js7cKNMILSinP6OX+eAyjNB5uttHTytLw7xJb7u3/1jnNpbV9eCqnA00ut8
nDO0qnqca0GT7pur24wc2UkadZOSdLm76Pgw+si3trLVHYBBosaHTnKVYrRcPQUSLnozMHBEE4wI
dt1bX8eE2AnSIb9JYL40Y9f+ajmLzJmARRN200UfdNlX4nHU2gRnupkPySrlx0RzFU4O+VDMtuII
t4kkgm4kO8DxqptdaO/JeGOyvutUvKyCfJEXMpFuEw7mHPnWn4H6scs0Ypc9pu3eZxQeRaZ6Kh+b
XA+LyLR2xikdokJ30ce9NlT5D6T9wSWhxdKVsvfbK1xA5l1mib9/rVC9iLwQlDNvetSoAZ2kRBJi
QoldnsA2emYkeSMELY3rQlGOXz/nr6LIBroLKc2M/tRLiIA7m2KUNukPfm6qdbWJBhsFyZSO3hCD
Q0vXiRnSOnvxJNYNZ57fR3Mnh1Zqo3PeDaFcIgagAcwrfhaTPuCVUqjqjGWfNWniPRqWDKjhiQKs
QZcWhkZRP44ZaGUWLav+9QPhACrybKAa7m+Hh9QlOOyHkdtl2kG+yR4s4i5tEJTjB6O4bP2Nx6aH
2s1a0K9kV3sUAWHB0XL/fBud8pLUYeYaX6VTduOQ3GmSno/Nzc7Xap+ts3nE3sLKan+qwz3FKgq7
2jBStktr3hkQ0fFlnkgjdvIG8PwCEwWcx3J/UAIVCHdQzjOwjelkm/FyrMZYUf7mFa0MDZGUW54j
wyBbTnnXVqm0vaUXxJxq7O9Vo/jEcZbBdrXBw5JKGX3huAcy6hgIzp4YX5fHa+kEQQJ9I3+Vimvj
XZ3NYP2w4NOq2CjCGJ9UEfqlK9I/LHDCdneiuh84HYuwl1DrlH7TzscOSL1EVh9mXbBMmQ7g6FH0
/JT49tRA+XSh+EaoLuiDb1q5uy5vTYYEpBxwI1QeYH7zbmVNFy5zq85inH8GNtVMMhegR34KuAnB
/Rnrs/V7w+508L6dNGOb21RUdYvFswpvmhpxZs3Y/ICDeyVot3RXOJoy90wGNGk+UIhG+ezUrI4r
hiDgBu+5b/uNrKqVc/5z+0+yTU3HZFwoMDtyuT15EjlHpGC0OapQ+dsu6MtAAFo7azssBK/Vin8X
d6z9JQ12+UjMNirrYOFpMBntc7Ti69PlTOueKE5EzuBCHyl6+yId6otWdrYr8pNoqGECvTEUowH8
CEeUXzNxJRXFlJTFUbKzui0qiAe1rWGcrcbu9m0lUa0OqflNqdiluPQdHUZYTGby1lHpXI7rTuf9
UMFKhWDyHj9po5mDiz9iQlr/FHLTKkSgLP9TMsU/fCrIOviC/jkGDcvlKB+oWeWZV71C3GZZgImh
4zd5XmKU7bOteXnTmuHJwU+c1UOS1Rrp9GdGDy6CBjCoqCHenwIAE6+hV+JDoLxodL51mEIhAnJC
hKQgjWILy/6cAIhkGqA1czrQNoJdDdxkg0srwhg2XDleHWwxzTRgarykpFH2vPh9HTUfWmU9CsQ5
vfj5LVXQJbW220W6WTa7uS59SgFXKFmCg6svfBeg3Y/vVGMCn4+B+xXWaBvG8m+eTkU2jXIdzFLf
bVwP9GwukNvjvNpN6mBzsR3dPR3YwyyuJWa3R3Ux7X8LaGQXpV0DuyDFAALyFWussngofbIUV7Xt
jiB6ZOxvmSKexNgBoJQgtOUpa6nczXuqRRkrXgQZswzwsFZa9JcXyY3ldgsl5486XBJk6bsx9Q5e
PJpDjxSZ5shfPSG1nnBhZP4yW/a4a4n17Is1YEIRf8x41fjYtYAuN6bM3Xk+OaCI6kX3io2KL4YI
eKm2uu1JN2czk22RL/Sy86zIe+O8tmVUHeWV1GadFgIBH5AxJMRT8lo4jGv4m3l/QXY8/4JgVvcE
qK6yUBEyZ+5eMohhnIFHT+W8jeADO+JCZI3lQ5Gn6O/zAr9tXJsrI0tSRMxgLzE6TY13TcWOUVHM
jrVZ5VrZOdu/qM+jJV6OKT8AEyzGTYJEou/ei7C06+gtaY8H82nEQFEJYu50xWzoOFJ8OeiOZpgz
rf0W43wjMeck5aFYpTzB6e1Oki/grXWf4qVYWod8bNnQ+YdnHJYrc3395Y1gzdZaJg89/m70RpA3
fkfRNDEEGdpdhjCK7Ec4TiWkpqAMsmjimfyiCc8ZHHXk05jNeA8hVB4dJ/Ouaryd3msWiBmhZb8s
F6ksfq005qzyo+bx41GOEQY1LHUgxnm9n0yt+5ji4J90ysC4CF6w61i6zZJ1cwsDUDXcNku5hA+S
Tfq/nbpa6pF2oLI3z6Q+URFTkpR5l5gEscIZ4dgZ7NPI60cVmtA37oSIWbCbQ+KHfQzeLOdL+zHR
iXxTeRldpp9TKUw1iJesoXfE5lTBD0AnJpRY5+d013lpfJzjdhLOgzWScjen0p94eetFGvJwQs2k
MBwrhl8TUW4vrmrByYH7v7mapSNxiGsdveYK/pQvMJ7NpAdcK2gXDihChffLDSTUGv6gwfgolLz/
aTjo7qy6JUSdRmAL/mZwr017lf8DZ5H+uoDftRbPFuKcQoDtBfQnAzkUMS/QNB0OVa4U3BXOMPSK
jIKfwjBjLKTYQWoxXOgYGzENtB9PKAj4jutExzBADiY5w8LpkWaRFxVaeeO3tfET4SyRBhkhHegl
8M09pVLP01s2SGCsggIec2ivXLVa6Jttuh8sPFw8/F4Ug0guSLQqS8xhcNbcNfOqcepE84FaJiyh
ijnV4lxN2l0wUuLBgVlg2JkMFrlGaSwvRQOXVjXfkbH7dBKOBIjj9Z2ks9IEnITncRO4iPyojBdq
XtlWyWny1JdxFVvM/IzAQSSxQpWv85aAlfI8j3fpvByqt+bRgdTBHOtIHyAEoYEEvoYT9AHaQeF+
GXDePreEmepqpcHwCpOlaUbUlXZA15e42+pNwjq/DhHMYXpPRJmC2mqPsBCXlfQSB/xNK7JBn8VE
wnb9FgEuV+H+5FycekwnHx/3tK9HMpSnUXfkxMFCjP5nF+jY4O49FxXrcIwDIqZ57G3421HT27FP
SrXBpI7KKvD3vV5Lzh0p+nCSqQZi+9pgdN5v0BSK1ysTks7ZNag3AU2UNO855BdFyAdcrQgiitcP
3DxH24OIoLU+z/oknOnG00KOLgTQaXymMQwl9wOznDZ6DNQBmULokfNnVYTetA8U64Im0nY9vKCJ
ophgjITDw7T9goExZs5+S9l4aMKPxm60L6JyibqJ3Kq68d8fQQ7YM5Hq5PFcuGWHaiROsmC9yXI8
vrqkq2s58qI1zRgLaiKYXaoYxAzGm06MdhQ0wz5z4WO/skIpd+KWyH72vDehQrgBI2ke1HRqa47w
KV2QTsjoDeY7FDPaYDrIhYAchhUxzynLlMZ8WFqnG5/2dCDY8Kh2H9c3oufT+iBzFM6RfvTdGFsb
BGQJsCLzFL7JMkY0B2V79reDqf1oRBJi9n4rwUZYd9pdQypx5HhLg44EAg9/fa2pPgGPpgkXXMhG
KbJLAA7ZpEMNjCISd4j8SpZxUslBxuam6rnfpLCvZ2+cZ3HS6/FiyY+3M5JYbPqArjgUhrGb4XB4
1+hKYjosg512iOjjNdL8ryDHTvcQ+tB7jYL8TtlTaijeJiOkTGcIjJO3nPmVPYM69ZfpALjkakRk
9w9IgzAr6KNIkueXsBGXVWFFB8MkPoDZfynFrfNxmVp/ROjxSYe+m21kzLP/yQ5nOaoolHpJ1PZ0
nwOFWwsEdJq7fgmAUmV1XPmCQflD4so6LIYmoXXh0Vy1K5R0gtW9n4bpnoWV/OIKb9DyxvyfT4Lh
Ic2jFYH++mxhkj5FmoY0UVt2Dg7VbNT+H9BIJ2YiqDkHLkhASwuER7BR7UTLNxoboLh2+hM1sKRD
qUXYgI0IMRfE530KuaYOUYCICN98TC25yYZdAXfdDZ0h8gxw+g2cpy+zhsh0FEM6x3fsOOcpK4cs
M3WBSZ4wZhbQFZm7BY5o0uCRnSnFE609D2iT7aTi+kwr4N3SBfq70IHmntVQ8I5iOxT+eD9wc8qC
fYUvcy/akGT15mv83+25IfNCjRuR9uGI/jS2KGyCRqBpMYx77WJbQY6W6NBGT4XL/8HU6yF1xlM8
2WQpzqz016rioPxZoxiLsKlgGfQBE7j7P6UVLMieKyLfVlyCOGh4SNhd/iVRcTJcpJes6QwGn2xg
sw7T4sWqbwSEupI/ijdKKgsV98tU4uD3DpG3NS6q/ewNpO0/ZZVYxV5kFFWipGNSvfzxIIQzqih+
mADVG1pBjzCsl0fpXYe/Sj9PQV9ryj0qNvvFMHVjbMuEmYpIp3PyjDkhXmLELbdeo8pFbR/WxpM/
A1Q+WQf8k1MDZU2ZQ5NZfRN/jJRy9RMAKwN5Q7kcOSrRRBTEz3elV1NmngfLNtjwlfvUEBOdfoVQ
kgpW6rcVUByJi2B8O3nwie4tjc5hqq0o655pnH0beBZxK6jG1YFPCSxnrfAsbH0NpG+K1WJqVohR
9mEZHDjrirr3bP/oaVt6ilhGXN8qFkyh9CLt1w/l3XZtL9HDe6bgoz8nrlSVAJtn9ea6ayjZkDAB
qXHi3PvrBhHPLYyyh3NqMNWvxb+c49nFzwIL5bRg9IjZ2xPTfDgJ1zuGhwlXWVze5zbjMWzQvtW+
YaAZc0wlXi010ig9KGPT3vJ7wYb7T0JaM1YyIwFpV0CrZN+Er20CIjHC91wwg84QyW/eSqKB4tLX
vBS0NiOR96C1M75KNck1QLhqtbBz5AsYZV44IsrmXLVQWsGT278trGwjvbFhVQUD4j4X0nWMus7n
/+MIrOUOlhN9ME7kHD0MAqv9TOuacI8COAmIh01dq5yVF/scvvUQbKpGPJxwuwuaPeHmquYj2Xb2
4w+6ZLCJjo82yi5ZGM8xC2o0O61IRUbGDLBtbm9SVYs6XHHQFROcOVjdnNagpeYF3DSwve47VZMW
xCdcB+y9zMLfX2hGGZbluDX3SHReOXBXu+a++yITBf/EwgyCHvQ9mMUVU8KERdKY3Q03/4pRyQhk
IWk+BYrpd5+kk/jPKRPuB1AFnRz5IsqZIXdGm2KRAW2rbugL57XJoJ/f0KBGoLxsB6b8z37OdWoQ
iaLrpjrqN9zDUnzxYv2qg3uAhnR26m8MgNvLLZ8rVYC66WjEfj1CDGxX1Il2dYXzCqqFMjrs9W0q
YumeL9nOtCdyshZWHeeh3PpxhxJHD0TU1RpmIViE0tNPFsGBFJz2GE/EljWrhGtP5yzCTBjCAzRA
Z4twa/IVUlWC57QF6AG1C5ZN8YCdPWJBdHEsFbB9qDx+HYe2TpAhplxktfCfrv1/bfSMh46pdoEN
OeBysqoAzX9W1ZruGHB8x0RzmmmvmRIGHgXtWTQVg1GAzZaSLp+nxGGJfLuqTwHOUPWaM0ZDLfJN
HL01rXPXvUaucV/APBjUmahy9JgVMy2QWYMXdIPHShJjZhyaHVP/zlp5X4mUGEoatcvx5+WUadZm
QxyHyaSN3caD9W0tUWWYL27FNelWBGHykqdZ2yVzGbBAU0BCGuJxHrmbS44lZ+iArWTL7D4wrY0H
4LHq1lkcNrP8ph1YIErNxrQF+zw9LGqnwk1J+D0lW8Rd7QQyCT1AJ9MsPfqQPwHmZ9se45lpfM5b
n2Qqz4+r51OxKUrG4o0k2bIhs8a1afRQNMFrrBXY52mit0DPnHqkmMLIqcWFvUAtnMcvl4r8Kdwh
pBAv2oyMkq2T/LBMcIkkZp2uDTBjxBwAybibr7ddehD37ZNAf1NE+ujJpzk5+S+No9xmbir6hzoF
YzZ0kwYehkUQbs7aq+MuAIjt/XGGkCyEk1O4hf+xgMma4pCpcmD1EnjQpMMg4eJjrGhtpNMe1Jn4
wBTxPX6C/nUzkuFLZ7ZC61afhRxIJ2J9pGYeKortDSc9KuuFp71ENPh27XEiPjdjMmPdLA8bW2L1
SJdPcW7LDAD1exL4DbJI+RcsjJjQniYf5XJ0IIMaTKgMeplANBsEk6eAz4TS5+iTiP1R0wQMSmoP
+tR/kYfY2J96XUO8x82tf2XYrTtq7QlhkDUs8yX68ojLP9d2f5tNeg5nhUgnK5bCebdLamiEyLsL
dx6tfcJA9X3Q4GnbrBDVman9ae03oDPVNFrTbwBH+1MUFbwSBYGQS7YMoHqlL1e9GrRSPKttd8Ww
1kDlZ3nW5ot4Is8P4Ay466hFobRbGFrJ2N08wDn5n083FMl3HYv0URXQJt5tCBWggmuK+OSjaNtu
nkBoUag+S2z+bXywQFvf97YcMzyGIJ/LCcUlpn/Vhf56Ot4TUdF9mEcdbQJO+GnyK1S/xo+YIahA
shRJbmD0TDj5hfTYf5iKasWhCJfevcCWUbNQzxfpMunmC0hGhCl36YcdSDslkQFuw9oz53SsSB1k
UMrPMq1PSKthzhXLeNXM/LZ5LUB79zbt8tQAZOl3vsUFgjftqFXiwYT1Bc46xOSVjJ07arEi1Ke1
uVCIypIVRKWcvSMdmtM1nI59eWSm53OVAzsouCAm+1PVIx3tq9rHIOymA4dyaAeLzpZg7c7UMFkM
LPpDz6iRC9uNeaPaXtK18TEWvIc93mvvsivo1s1+T6mVeMldedyCTwEFOUNxftkX5mHJo6oDqrMT
3B9KpNr5nBUlY/kXlTWlHNLEevpnDqHdORtW2oyGzrVR5OzQLfUt/eguOun44fuhgNN8F+XAb7Y6
QwWeHqQ8+zKV88sSG978sIT0qkEmDNff6XZn2IR3JbyPZ4BOzAIGLNTg8Hlj5LeAEoLe5yajpAV2
ff0vzWYupDc9eLKWXsOZHURbMe9mervomi/Q4mdXkX8E9daNTFEoAwYfRzJz3+zs7nZguoI0ZtgY
UTOg4PbW6ycnVe0JWwagpH6yKx4YAkizQXZtZo2SWMxkTyL+08EbYRcPvMR4bLDnE1PHL9a3daSt
cZjNbRGTTfJk8A4976WIvQa1yN/ArH6FBlPF1IlZVj9YtRxd6Pb/TWcNTx7bWAQUUtezmVGoUT1C
zvI/LYTpKVa/zeo5vu3hOB2qSgheOeiYysNR9tY87uCOZHdUiHVOfkgFWkxKxg/rlOYyeQt/dZKr
L1wnv6NsK8M4spdhAex0aIH4+5Q3L/ebr3wHWhj+tm8n9zPAhukot1xnSyiYK2hTOqF1ze7TrcQ+
yDGC+3ONK1dhl+E6yTnDB/ovFvnQAuMrtNBFGu8QrHQtPzqd5NF1OaF1COwVPOJhFMZdkxEyez7U
0gzMPWcBdDSMyjWhc9NoszSva62PpEpgljnTdxHoijiuw7b6Ur0mIFNypDlbNkNtm8k0W0U72hF+
Bmm+CEn6CEzRdtWByBx3hAKvS7nclCFXNnn1jqe4xjFwAAUPMfnuJibESB9e1X4MgfHp+I3JJDCq
OGFLVMDAuFQatsFCeow8Ajxir8zpilN7iORfVpPvPg661H9IpB7AdcYevD8kSOqkTJB4KUCRhv3F
y0Wrdkn8KIU/AOgqtqPHfUfRtTMuO2fq5SQsDrkc1+p/T0Gip4O1rGFg68itROvXLgNzcrGSrjqd
lCItvHckQgIvkA/O1JbD+PA0SWb42+8uyiOShhxX3L+QMgd4pcYr8r1V3B/EGGuMubPm9dsilfwW
PI1FM5fA52/an6n15CuioONWpRoQ0fEKfswN8j15+xA3j0SXMwMNov1dtPXzhgEkwtHrbklWJixA
QQE+6YMKlKyJ82RwC6+b+2je6aeR/IhJRUi6EZwjLVw+p8b2CT/pPnMFVDZH8q5OPEp5ZFqm/BOl
g1E/+YnmHaE0ajSfAEr7AP3tuQ/FnlwgJ7iobRNexbcYcwgjwjJLSQsYr5yI1is+bvfzAyC+4Rak
w1rLFUT4czY/I/KaLzQcPSEE8/9UHIOF/FrhJDL2pdIeGkYWmccn0TSlylUpNwqWKct42OOMiHMq
na9d7/QjQn3ApEbnfrXqyZB3jU58dmXtYMnu+AyIQf7pn0RijsDqL2+uH/9Twjwwr6r//guUI7/n
VaeoCZFAWEtsqwaGVXB2KNhUuIB1ekGle0rU2QukIcvzQqhXbXjS/stYS0z52RfDM0u+HUwVJWyO
dk45rcgpTpZ3vfUTH6VGystUEhGUe0hHpazSlCq72yJupDz9YKXDJVs7mCxpEtZbQNGrtfXRov7G
bR9+rWiryef2PMDUeG3zLIPpl9dkq2/lo5LKjASv3yHJ2HZqS4W+kvGTppcdkJtD6aYl+cPKHk00
QgMdIVLDFIfXUJmzvRtA4f/gwotujH9WIP/N3dB0yBUNg5nKjS4gBEAr02lyNNL2G4O4vIq06F7J
P6F+VVIYTbH9t7tVlKlQzUq3dk4GZvsTQlbvD2skEgGhugqqTr/E0Yg6rhz8U8t3kipj4EGWl6j7
07H5hPnoKXGIoV03pulo6kO3VWT0buXd6kkRv9JdM/gfvzlUlklIjld4Yncr6MYGmeVW5Sjd+hkU
X3d2EmSG5ZwBZcZ9hSGG1E7m1rAQd1GuZ5MAeCXbSwQ5/5Bgt8zS2zz6HW5LbtI8SBmHraXYvF6E
27U2V4jQX9VXP2cAYj0Z/9FcXTp8QSA1FTu3U85uW39IdaY4KnMD8gEwtzSCOGrroOPhAP1LJsPA
PdwrO8GHf5J9iV3z8mEYMyQgkvhiLOXdbjlt5yjH0lkFTLZM8rAx1DcdyhSC+62OmoIAHGKohqYA
vn9/pSW7Igefev/x+Wfcs+ctTTat6VcbfVTeZFuhHpxkafzdRP9oVRNFqWoNgqeSwOwVL7HL0MG9
SC2bem9Y4lLvZ5HVngHOg52epQakuZkCA3FtI2DVNaWyy4J2tgy2KEa0LYiytQSvLwTXMSnoeaBN
JmOlH0mqXuLamK0cPc/nYGNU3hgup+cmjX34fkf9+8oed0MRIHx2T5OVYBsZIeVIzfd5cGwR/r5E
D45ehxSffLobiaZVTMj1JKBTTVknfjF5lK2QvZffV/teDItxjp2B4HfgggzN7M2UgABc3S0ioKqZ
B4bnBBKMrkX4P63+RKoF1l3F75X0fmQX9eI3V6BoPaF9KzVvxLwE3OIjeoJpqrULqsNEwEpJqH1S
S/9NiZBHTfqHUmbWjmdvDLFZbITMg/naoatPlHZwEaaHWIHGXXD9Zqn45r+dF5TBFgvKTxqMfMr7
jbxkjeYHInszTi8xNDwxoOIdrILmJJcQeen8GH+ji0BiumLMWZQ/pAKn5L7B7GoRQP+Y53zfZh/j
wbDfauNs0vQcypCY8d22BkML48PAktkRG4MG6fBa23zYMk7j+gsrUsQPJwjojITHHVjxsDAetyFR
woOXCvKHI7fm1uCAsg9aynXGbPqDcUsb6kq8pZKClx4lD5AfTIgsfJko3bxAtvTPBFZw49p0kwcc
8rb6rM4qz/tXOfx1rtmQk7kdfAaTbOs2GwPMQ+oqDFs5ShohWZjM2fvVkg4E8RR1bsjgCSCqX9sE
chK46LtjEl1+W+puJ9frUkjfj3xKxGaku8OC1utqCYRqN3vv7+7iXj+FbEPs/ThUXr6wk1msPHSq
JPhOI4rnYKq6Te/cgf6UbgT6MflwocVAcuuU4EB73qP8pLG5k/fViZX7jpfvV3cylL0TRKolZj1Z
kz+XQhdVVCt8S3rzwPXYgkrMHZWEsAG8SDpD6lkrh5fJ+5tfMVcsFLCBHY5sNp4kkzMDtJR6lQKN
9n5Wg2ojIk9ZvutCdgOdCl9hCbFPrWS6XwMTD/lxo00p8k/Wmwckitib6o+NQMcBS1tHxmZ3GzS6
j9ZYZeqsmHHo7JWdJps83az58E4kk/3jHfRJcB14PbRNqCBBSpS0Q/x62eZLx7OUJqC7Pc34s7Da
O+lET65wHUfFu9tS7YEih+dwvmdqwDKcm2D7f6A5FVS0FS6wERWMlM5MRxh/ixxeZic24DA0WH1g
+gV4w5qfkxUGkd6Ufoovxs0X/FjzWsmlKnvKkg6f74aaShjGCdV6ebVE/Mqq615zp3/gDeBoH1uD
KjGZWw0EUhlQr/g/7Ff726c5fcbVj8pS3VFTQb76ehGn2S6zhtVSKraQbjkfBJUzhIsKar9kYs3t
UUMf7qeJdr/gF4fvSj339sEyuz+NCtREpLeyTJeCECgIO422u/a7Mf9OFmo14UaACMO4VJViXN6K
LDiRKn9EWBaVRC+TKOiQHU83rBrgeC0TxzbTf3Me32Ju3afOm1eYdzqZzh8InRJMkZROqUtIoMw6
IgDa6SB40RMismw/AGxL413hr8WO8hxZZT7lvAPzTS/0hYmyDl4Wn84FGC7rYYjNxBUg7648JQf5
2u7HLvpHfKmQWRBuQOTsmDgEfRUFofDENq4/EnlNsgoK8ORED2xMeXvXu4+PBNAMf4RLJGJzreDz
F9jBgW58Hu2O6mXauSrWEo1ZFoqKzFTY38wGUE19IgJSkv5MwhkfNas8D9UAriE63Oli0YxbUmoQ
+E5f81E/xCfztSpLK3BBA27xt1p9QFVdAkDZTs0AjrMII4oIMPWtu48ttiLC2SWIxWeZXmQucrpU
7m8nQMrtjcmn2pBB0Zx9AShzC1qXvoe3dLUy9XUEKKjUXe/WuuMQ0v2HeojhC8GAbYsJk5cN8b6l
SIX0M14xhaN/dDTfOh2b/I5NQpsUY0c8pob1cahLhi4rDpSL/qK+hE+1X8xuSbutQcMP+EtnPc4j
Gekkw6JiamfNi+WdEeVNdkgALE4bL2gs3hiEW54n8YzQYqPqU1xqHtHqANs6bDKfAmqeFlBTuYk2
uifaOhBhXQNiqCYjCaGncLpe6nUK3p56RGJBqyvdtp0I1nIEA/dyVRr2jdwchRoAffqJygFGJKKt
ko8wnLGuOcez289pkiOrXzpqOEbcxBqTZjJ9x9OXxAyYxaUIjqlCwQho8fOzZgdJ1GLK9e+j+Uio
p6YTa8VjluRCrJwdjiq6EAAW6smDQhXz1o5WdMl0W13WNcUBkNL+9juD17VvsXMXuNdFSnkOThBj
J5CN4KOq2Vnc6CTrtwwuaUuUhXPtycbUs8m8WgNHK5BA2l9LZ5SdXjIC13CfSNoUCSIjkwB8OXnA
Wq3M3ivDIJVW2pNSTOGNDjlHPBTEUZMTqjF6fcgsfMNBLgKLV5x3yQtTKsV8G6W8/XMrMwlrRn7b
pVXJcnAaO3iwChLwh6qEJi5G2IDIP59K1F2L0utYYwd8at4DCk7walJ//XwGUVSu7aExxpswOe6d
LqpD+fhiKJua9ANgzVL6DutpVRF83b/SMb6gBuRO4vbAElCaZ6fGJBXZipEjCWzxnH4Op39bvsU3
1dozL42yDRdo8mtfvIByK7REPTh26L4SYPyPH4QlctmrAjnAnYLoO1NtP4tHUY1J6gn+1W8EckP1
Gj2fCLZQuAP3g6QoDaB6TpiLHRooxw704DFHOL2qknbDFwDXwZEaI84VuV0zl1yH5wiGGUdofo9e
MgJS9B52uL3Ks6IsSvEJhcxTx0uuXK4JYkF9LzBYCzFEe/JYhH4Dta97vJAuGWOv809pAhHGBOZN
CZDG4WkJIL+VJDvfvy+VLfMRELkRZ/pK6bh5zMLG32ChP0U1l7mraWZFU471CcD1sj9/WwlTV23D
IVuRMoU6eYnli5sR7o+oUg0TF26KINfemdT4XJd9whwTb4WFwxc2+efk/am+C7DU6fa6gK61EXaS
bd/L+uWtGx+y/SYRYljPvy1nz+IRsuCI3D9BLp/rci/Ey6XHkYBcD1ckQfQKwXjmbqooXhb6dJRM
hOesq27Fzu1tateCBW5WNyn3/psrmE9rNYxirSEl3PZcFHhWwJIEweDJjamykkuVZsw1VeJb0I+G
LRYgCQAQseqsm1t5nYU+nRGwe1S6mVT/j5hf7ZxFBrMS3wWe9zkLMprRPahB7XQWpf6EN09v+j/v
8kuz6IvTAidqxesof2OhHmWTucMLjSTSV44dtUVbbyx2cZ7u6iJhHyolVrrrGvtCWptetmEhOD2Z
WM04yUxNW4yhRj/1VRXGfmotNl+LlDPOShUHITIST3RNZ9pqJwVR1qboHlqW2BWvn7NEw8N301MF
o+0qkgrjHl55ZTsXYkaOv9mXwHuELhKcNCXHWIuOpM8By/dXQdsYT0UBJwwtTk36mS5FIZrrP565
KAcozJ7tBippImj7JlWqT/olUn4FNHh4R392iWBdCAE0li4TdPvreUOLp5RnJP6EvhE2wLaEeyOZ
7lRSCt+vdHijCqK9KzbBaaArdRnUfSwZtDjAhTEGhTBCWSh904Z5Jtb1stbkkQeC/2d2kt2by9VB
3Oaxbry1QghXZ3VilpOx64EZArID98PhYnkQD7eQMPkGOvr7w38v+BKuZOcx4/qbtNs2qYPuglLc
jwUCJzwpLg0e8yW2o6ERBJKGxLsplCTuEqS5+N4HfMC7KtgWM2Xikc10WOroMAkpowCSa7KAw1+d
oMIZ5uLqG1mYQ2FKnw5hMVokmAWV8V5QUTqpE6CZuvxRA8o+qplDEDWS7QUCwFxybPaB/hZNeMVK
wJyebDJejHhsbj84KAedYxDNefsCBDxAdcK3VJDEoQtEAafRvJ8hwX4GD8ywB7FdvWrmuTxI6t6G
OMRXzhNC6ppi82r+WeURFL4Qbd0jwBaw+UO+tWPixBkCno9k9kCWdS7UfdOhlvc6DajlHLEkrp21
jSTQirO2DzUWbh2hlN60L8MweGPKDrHu5XNSkEBLMUk9khAV9uhUxLOe4p+QEVITPsCmn7AI7IX1
cJi58MyBI+iiXDl1fD2hPl2uOjyf3NmeCdkVEi6ProPvMml1XRTwK2Gi3xwdWmsGmm/R3tFVviAZ
84pJ1MQ6wCCWWvWKdkZcaK2u/uBwla8jfvrffAx11/g74EkvqP9/7ciPgkCqNpciCqSMo953MCMt
2VC+4MqWkEBDtpu07KrSNZe5wDznq7fQ5WVncOjuUmktawxU251Z+4sBz22+lCh0U4v3ruCMZ+XV
+6tfZukU7kmThkdICSvuwtx02Firq8LcFWztzVCPcm1pEkyXne4sCQxoUxYqLPFLjq7+nFXMz05H
OzRua11DejakAO/SF8o2rVqk3pvVGSPoqcNiJ4Pwj+JIQo3lkia3T171f0FCdZFRwBdrWi9/6nhL
qWoA/uZPC5jqH/ybtvuttjmKzVoF2y/0VuVYJI3YGk4RfF72tK2uXkjP8ULU184wacwcEmThieVw
qJkWRXYPJmn0SJA4ZHETe/nHSIGX2cdx8CtdSwMaAQoaIMWp67LTpJ58BNG37RcOlNmDDng105Xz
U1he14RVwGhFkcA2aPwTkSqTsXwsTb6FFXYahUugpVtCeYLHGMEIZDMv1DQrSUVU+TTI4gcp8QKa
5uG2DmOKhD17vAaCeFV8sJCDXmh6sZBGZMUipAIr69QgwkF7rw8RLmnPt4cfEepiefQJ2Fuo9JG3
/xXSnPRkyPw8rymKNbYYGei9P/sAMD1YebWcCDfllSk5dwWCAw5HNwb2dRTzZURm5oYiX+8EUvvK
M0xh94LmMq7pUlGV7uf95u0XavoY5B9/iUGTkWWkrs0JaWvgzTBBlL9coXXzsGvF1SIY8TsojJqj
0XmgEJKzYZjHtVXU7m8OF0nnraWk277G65LFqZYF3fOfnSci7F21SsXv44BnexeSbxa/9+aJuS9l
nHgs0bV5drhuKZqezRel8WFJdwxkTir+x7r2sJ2EQuvFzZh0/KGshNp3Vfr33A8OxMsQPbhnbcud
UCTOm3CIMXAXoQNFNOruGV6CGYeabV5ayb6uOAE/na2bkC6ggYW+ZqKsxQGcW+RAylfccEOXEH53
DwOaeran6LH86uMo9adrS5scXPRn0I28D/sROWlE11TYWZzWHLV8GBsrey9IiCRGEiLXoEIOkPKQ
x8dAxA3orvjcMeRgKMkCdlU9UvRsnEu6NOInwDC6ib46iCCCclSZctgOQyHliByr/zBUtoF1FhZD
Cs8fKotr1FfNA931cYac91lzmDqupcSNdY6UX5cTVvpbBdDUFoOPnNVCaVVu7FSAXgd3xfc5Nplq
TOXJi9R1IL7lqUFGGSkYSwDI1H3c8jH1mVeO8UgG9aApulS3mpyMycxcSyZNgzCEJ2EoT0pRIXPG
iem0R9eWz20d9TQNyEi69qdJ6md8hLMbLRkjcqHhlUkklIlxO7HdBSxvz0ut73YF1Ph5kIkwPgZm
S2l1FMqj4HkUYoyJKnZ/YK8eWguxsHVvHnBBNIY2hcxMNVs6o16xwifNKPtERYR8KVqZ9KLIIw3B
4XgnAppN4NRO6ryVDUjGkZsmZya2Y/CVeJ2FZDdzirCTG6gKtYXXCiCxhQ0w/TWv+8ezZ2P3H+4R
cYkCVnJbiM1h3gYQbCyoJrdY+53CrL07Balnr5G0NcJlAuet9tMyYnXYlnkgwpU6PoH5u3RNB40M
Jxb3bdyfeUNLgaBk2bJKeSqHKKFMbW+nMYu3YH/HDDQPPM4sqQdl9zDw0/ngsI6DC7rtve8ncvG1
T8xpFD/W81KvUSGm6dSbVTGSDnkyWHM9SJRiN1WsJQ02JzdvcRxnM08hlboyNfWqWwIQexk4f2Vw
4/s/pkaSsOybxNKiONkPPUg3LbClwv0QsL/HHnn3dYlEuuK8XYYrwjbolyjCfuwHztQCBCXGXC0o
PvcD8MLPC99iaf37ZRRtBGXXsU+J/a8QQ557UMsfRiL5xB8wDpnLBBQTbXom6wkFf31RsTQS4Tbk
TF9ZbJlxIW6dv5T8CpnaN8kjApVe5t2OjMMBwHzBOSRLvC+mfo3qVDL6fnLcL9+TzljTGJj2k8BI
JwfoxFBmK+NMtgU9Bl1+gYTHskhQqSlL4ufxOgeV6LUfplOqK07HV/z0W45KVWh9mMQjXlat0D98
6NCsa5RDVCZsqDA0wLe0pY7jJqrQc2NH0FRIM+TQzX3h0lhiPLb/YyFjANjGKMlo8PMmxWkAFd8c
Zyxf4Cp4Xk9pkZ2dIzx1ZrwEWIE761Rboa+xU0iQSujdm8Nv3tLM9Bp/CVU7TJQAIt34EnwV86+A
0N50UVvcLampVA76/mJ7GF7qSdmv9flusfB66EflXWw1zPCM8NSsOmvAYafeN7hnHa9sBSzeV91f
UrEe5ehSuUVSFZ7pXzc1KrCnz6tk4o0OqobJoUzc5F089m4Ghreg8f171YeIXaF/Lv8EVJ3Jy4/V
IMM7mBMfzXCJTzWyGiGlZ0WWDZIcaU5MqVECZR7/dLkYWdToeUXZIK4pe1oSp/Wb4/VgHuUzSXa1
rQMkWmAJ1xWA8TNGqW6G/0tEV+wzh4EieJK9SvFO/O6EQrRPJ4bKaWLW9t47KIf3ZoxapzW3cSXf
/U6MGidmSsCSxy7Vb1SQ9LhovP8lfI3ACq5Ckj3vUEVWlvi+XIzN22jsROcll0Zj/9gp8sYLT5on
p5lhwY59IhP2uB7AN7aMZ0wJPJ0ONNno7NWctPTPaUmRJmyih+AUEysh2N5/HcCdsi9r67M4GG5b
MPtGgbW7e9bg+xd6Lz8PGcZbhwpobttrC6Gfd10uFgUPhIqxBrifGGmdii+U1aSZrmoY+Y+zZ84v
N0QyplzpTb0olW0hETdrHGy7ZvPdSGn6raFp243/yJNh12uYazDui/f91IpwcT+0yfu6jas5EKfI
zFOlyepiXb5OWqJO/A5H8GWDAV0/+nkDyzc0Hiq7oYCxVCpS6jlWizuq41JNBcRXYlBKVGRfL4ge
CIfTYuJ3fxwMu3VyIhXJ7CdjWY7wpNQbCJUoeJPIymRsEUlZX/0U9RSUqhtJ2FqpSTUtUwwcJHyz
gKBYgHq0soSxyQsoaOWWy4C2HEkZu0tWGput/OOzRLfNQc+V2wiIjxttML/hbsbGbdnU/8XXRfZ9
xqkk7zXANOu6p9319X3WdbAZVGL4Hs3hdyxpGVNkHfdUhmdwURc87WlZwRPglA4F2LM4cTBvQGwN
By8q7CQdHegPMPH9JgCZdfFtbXbY7WGXxhaWMEf3Odh/MKUHJ2Z0wY3Z3za/+MlERMO8w1rravW5
7iJKF+cmS6K/xJXL0sSedAnioZLgofqnAB1cBxyst91JWnK3Ru7Tglunf8Da2oCoz995y2oeMj46
J7kTtJzTDC5y1KTjXpR0z0RpGYMPNEaFzL5DpJ+3VCHIrTpgleOGFtk4dku1IyShWYmY+8nd5ZIf
XOVxy4cKYXHbnuakye0gvYHHW4BmSHf7HHSqyZ4bjJF5hSfArh9YQWlQ5eT3gjxLSs+NRdA+0T1e
dAvlEKrM76aNOQ974TAErmqWsXVprZiATHeaR+OOuNo7JnZgyIW7hw820kk+Lomdw7yxT6+iObdL
daiexfU4R5RWOq7UvT1pJ1uDgW0491m0FotHjMVvNjSNeFmFCIGzOxxPtEH1BWL4Gn7yhY2a4ocR
IlJH2kRXogUY1Cs7YBcrB+2WVXOqXf0mEeCzM5YWmhBAZSZATJArHyHRCfY/PAfISCpvpxaZdRKs
dlpHIN/NQL+H6BfQyhDoaHPhP464gUig4MG2XqcP+z/iCSRcKe9PDuqOKoqYWgLwwlUytRRboI5m
IVTsR2xlvgtqdJwKULu/upEc3R8zU238jOIgoTq3FACWx/hjV/LOmVERcilCuYcrE0UUV1Nb+LXL
Fjsp6gJ2PPzAivLGGLMiTzqwC3iCh7MKH25MdV/yI0Yyzs2Keg/crSvnFZ7tgxtPM3BZ6kCTcqq9
kOOrwQS6O1l1HinpuyM2X5Ada4J26HqHhJKr9wqlfe3+fCYlUI+mOUKRQoyUjkTl9BNs7Sk5CmSx
t5ScRhzR5W3SmFGqdm7FrHUeKgWXzoWmymcMEbHijl0E5HjEW/kn9CXG6bUbPHF954zQyMjBpnz9
rn0GPm6I4Jeur7ii3gULaVHwIOG2HNjFKcHQzPiEInPqNCMjYMbgBywSeE1oLurawru+db6fRcav
IluWuT8OiBkj7YMTZ09uQT9oSwS4WXt+KTdVNJ1+mXN9lBNQsY/DCve3A+JD3D7uMjAo3XhVf0+Q
3LGsPRG0SjCO03gsTLOeDqkLbEfXsVxrG6I+H3q23wiCnMKjAZxtefJn4Z4AbzcbIKzifamvda0f
Xu4HiS3+SjJLCBjL3Is59i1jOHaN61qH/l5orfkeQWJEMhMkA3YfUsImZd7m2u7oCOlhTV82PAkx
gsbwVVykjRElBXgeQcmlHcDeOHaDamnEQ6QkMogQTps7uj0coPAJWhiBWKLxUgGOeCQ0zZrZ/u2/
LwKLg+CYGeZ+j3xKlntGEtv6latWo5kui3yleOFhlVh1VRl54GovjK1DMDxJO2hjSvMjkjK+cZc5
3ysrn7wTj7F7xthvYLqoXTg5eFiIrVmtNisIDLkomF6j0Kuz4gzWi/ORMvw2fURjEv2A5KpDAUvI
1CJEq/mrZKj90UHK4psj+nAXO/v6ORFRMArRgFTlgCzh1T8PB5hXap8GQQWo1XvjGMbsEITNkU2O
1hnQMfMMq2hG5rdzEmdXDFvad2BFuKC2rFztzhrYu04A8RK2EnZ/KPfr3UwzPMrjIN33nzIanRwX
1xzzhyXuQ0EutsNNYS6TlYAA6HM70m7gVuh2nomLydP/oSUgANKB1/wdlwKsuwgKguOdh+UpwDcE
sT5lBbgA5/ATH/VUDeZfR8jTKHYMzN5K73hXf9CdFQX7VyrsNAFf1o4J/ylYAtpWCJ4DJAK3fN9W
/S4ek7TRPeGulViub5imV7nTaa5RfBqtyIwCv03hsGWk3YsrNTn8Y+/OQIVx/32H/p7lztHhDWub
K0CYYl0ocCtc+D3YqMjycas8MYqkPPp8RIoF9s0S5ldJs8VaCXXdDBrkmA4xIyOtVgrQJ15Qddwb
ZFvm/ADUzMx8Oz2k1ooHwRcXXOuhF/UMrHH/DWv795OhUQbNiSGhDc5iu7Rxg+EBaF/+aPyoCWG7
kUCEMxYEVXBhPKD0sTSY790FiJ+2L7suWVy0LTWNHPVZK+8Cjl/6kagDkXA9Ohhh2BVPbAfy4AHG
1aO3n6EzPUc7LvVu5aT9bqJfK1h7+92rStlkYuyY5gJlWlY9HM0OLksVrD1p7BGLDfH+zqE+FJxn
ql5h8m3VbbTPKUnQA2cq1etwVkP4bGTHfJiKW9j2oyy6IeHKyTE61Vq1Sokbouz0AohrfBkiIeoQ
r4WZ3HmZwAI7k9o7HpjjJ1Iqe+n+qcV4xpDFTDBkJZY316zxOrIWvcTSt87OTyBzPua7EFwouktt
bDxfk8iuyIf+hxb3bNVXCnU8ruXA8ZlBLECjXYZiCXL/sD6b7hmVI/GCrvEQKeEcpnc/Rd/YfwzP
4eimH+jDpDu39M6JpHyfo9zcteb94rqBOB6Tw7fG1sU8XepP2G5B8AshvRcgkQ/LiawcThdCMbqL
dEzQQbkQYvLbO7laMztVQ28uCZjRMzSETMqQnz28JtK+dR3BzqZnGZE2dFWffpTJMH8gRBoe5RFl
vUtJ6OGZ1pBCDMhdHCXaJFKItO/mgQTWc3TO+4SbbgvtfpNyzgFJGj4Qfe7PbhFwR+1qRk4ohCd8
RRdCrr4JcAkj4K5li+mrg0PZAtId7CumkctORfeQnv4MKQHlnNe7oLzyZ/TucKlGwgCBsbwrtSMV
RRGk7OnHrqmWWT9i8BpL/QVPPYbTW3s3c463YCckZduXk0FnPLnqWqfxKly/s3DnAVlaw5rH8Fiv
wRNW7PZGye5AHtVxvLNFnuvYsnd2yr4FaxRSvJIQ4e2f5LYK8+hN/W6PO/gampkvq2JCMpzpnIlO
bjEWMxORhkapixxxPAHV1d45PAriTX4e5pJlTTEeWnDTGS5gObx342SAcliidyqVKx9GVzRy8nzg
JhMzlXOwN66YiILi53n/vsqEEeVm/t4FF9pZBWHqtDSrtpTeHoQLr22Go1b/XY+Cb6NeMnaMQ6NQ
0D56IEqqvf+4PF85R7Hw2pWrYnJqf7KLByUD4kro6D+y2b6O5j02rU1YZBH7bTBGqKTvmq7ylsh7
LlanSMo9TRTbWe/XkXj+gJxFQvxwQ8aPp9AsD+RUHHy1DeVHj+DoMs0tXtBfI9i3t2AEHzePyTIm
RYdOQsh/4SCJyUsKMnZGBQEmXHVaVT8rDQFuwKuozktbfFV6j4VxBCmkmImVuCFlnDQORoa5h2wX
MK2Y9BhmrLFGhPsHur41YjcQhEOX2uad3mJHPbsf0AJ6/VeTXyO1xeeyX99DPQbzxqUitpAKbLWu
LtHP9t71a95hnqmVyPX/S5KDVAST3zbbzf035Y44jFTqedHan8RfdQii7639sC5rpq0SLPGRUTk8
KYPTnRbBNtUzWI6vfvGUOsaQ8uktfkadhCMHEC+EtqoNNHonYGmh/MUnnP0ZRtk9uCTIRfv5v0vM
lcMf5VFp1VPT5VuXAoGH+zZXM1JC6m0u9rBeh9A6Iwf/L/SXcfllhU6bLOR6TnA4lGRwnAzb8X6O
E9fLr1R2D+cpkPN2QYqngU92/KMw20erw4AXd641LTSx+iD+0pO4XWXZsTBNPJH0PIfpBpbmtxWJ
nY+YbxxqbRVBQpdw3ZPXZimuObXyS2CbwZcVbS0dh+7+HOILDsZQnnHOPGFDJluMD9yleVqBzhtB
LZxqsKdIXWDLKk2ZT6J3/E6kYZnFw0jdHkFYnbyv936GdTnF8fwDqIxwpY+W2G/Tj4UOc4aucSJf
ZLccamOsRSqD4swcSpZUdSdc32PvxfC9RQRYmhnywqwxoBvWq31jKZwxkGC6kybOlO1RQiFLwaWR
eJdVVLHcqI3Jk8pdD7bLkCatk/wXXxMyPtKXpxT6pSiT/BNcMolttpQPZ9W0NIarCRwmg1VpP7YW
dh0uoE53OBjEIClXnmyi2ZmxpJT4GtSWfkNs2QCdNOt5VpW1m/8bbcuuBSxcH5WcDnGZ+tx3ZnPF
KI4G/1vFyHhIbQtrRSIN2EJgE852aPsdsdairNTJ4yQSHPLS4h7tJShcmbbl/v4S0+4WzENfOco4
gNElt8ZaY6JMv7nyl8Lp4P/qbb3Sy0fU9HqmG6DiNSoDrnVHbg/widzlbflqjtqgC/N7ZZx5Wuk1
dQAqV4qjFgFj+QvzmRQpqpabnBJCZTNOROH4jCChi1VxZfRAAgk0IvfTwp0j7PxWMuuann6xFyGz
0JGM+UROhGcmhzBGzSZzU6z3jQ2tlY0EbK8J245S3TtEWbjpKhzfNNl5IuZNXlLtHUKmK8wwqdK1
i0wAGjhimS4Ns7AgYevR8lSQHgPjVKRNJ6V8sID35/haXQtw+x/CpkgyU0yka0V8dFA3xw/Cyeq0
7rwFTVM96kwlDmSZqfswItI48nCIOJfUM75CgCbYGv2njAyxECAXd5NlpVA6231DRGB0qU7dZvUf
eD4p9ZNXuCVllpZ+EDb+aHP5s+FWOT4sNcsIaoUZmNoXt4ESj0I9DwxnAV/fIg8dActhuAqk2NzM
diCr3qnhOeBUuJUzrri7gb9p75Qqc64tZCCyK0mfKwjnzdogeVAXFM9yLiS9094tXr57o0X+mDBm
LNtITpFYURwRgIH+/9GgZiru62SQ9pm5jDZgocZveXsDNHSPDavDB5y7z9TTLZjfpV9Tp7fuD6JH
szslSILNJS9HCa8yV7qwCkZGrhCQFIkgfYFY5xdEhSHvvKKu02ePjQ4B19VK3YzUs9LdZH9kX3YU
0iW+5GN0wYxTxinPoRiViATxRlk/nMkescbnpa9eOfunqPJ6pSHyAdqd9zfUGmshTame+QIeRtLd
jxA/JBEyEb7JxlVgXzcIyZt/tLLrEuxu/pWXZh2BFibqhERLAWTmmucqG0Ya1yOLa5eDiP8T7V/T
79kOHIc9QaZlDfl88ek1dxliWxOoUWdghAJRfTaWiDUl/tZ/pomYhP22/P9fDxLhD2nJQsUdOihH
gWmGDiPYWMYz3pCzn+IZpDWWaW4G/bMUcIzvpVD6tGW5wRLMQ7yQn3gQBBYpIM3vih6Kh5HjiKKe
E7qVkK5aASCCWZ/Gj4dzB1KNq2NJ7sTJMFyNHV1TYjQhFVRhMSOIS1Fk+fZTtgyEllVpgfe4DSiT
jwVFsZzib55IQaQIHvAo4jyLR2jyrJEufsXy1DUl73qRFXIuPA/AnTQVnIaB/PaZdOMd06S/vdgV
0lnU2MAjMprZy/2ATTOcEQI03eWmkbOccnshd6BbApY+fG2U91NcVcbfIX/sc0UEGYCAl1GKAx6q
f6iq5mZj77Xl2Hn2IWN29Z5D/0VXVqrB6srf/3bBMc2TetWyoOx/NUBIOZ1NSOVBP//W66lkWCga
jz0Ja49CppR++M0Zg2YUEURKIXelQizKO/BaO33NZd8Manlo7X8pZEO0r8603HohEAfBAV8cYjxy
tZ90s91RIj8YWogGU/ByLLyVjkDurgio4SDPmVCkU6acANDrlwzPJSCwlMPn9DZaKSTHOLeYUsjX
7WjBKfHFy42B4itDYDWJ81XnXssUBSRUc9Z2qkKkfWln92KdRmtSqmp+DNSYknYiyHyD2yjI4drQ
ldDvVpe+UK3qrDNNVvPYeDdurhTb2LzfC9XfQ2FM2xb5SQwKvFnDSiO6JdptXxjO1R5WgmUGQG0S
nkrTsopB23o8wXKQcDXekgtUOXBfyuS6Gf3E7kBOIhD7aCX3lZq2doHVbEH9nJ2JxhlWFcCRvBVU
zd4/1STEUz6UGvx0xnB8TpFgoHPMsveErEfkyy0pY6igaiMiAOhx6/t8KriSUB2o7s/GGZeE4sRB
J1EubR8yx6vrV0N6wWE5fbhRNRy06xQd+0p4Ac/cAIkRncqRK/31LRAzRLVE+y7zr1jt7XZ9lD4W
2rwRq3LiyCWavI2MtBJ1/a5F26i2yCOKliyJmLkUJ3q5YJAhyt8UVMjXCjYjE2QjhHJe9zd5aHFR
YP8+S12blfgyBQoIwSgBeQF5vYj+iFhnmT5OA+Kq7vFWOFJRhai1u1SnJKU0kDpwMbSbdNbzuogK
uoYKYst9axVMsCDriG5fXV1/crtRT4xcwUfTdyOvHdZt84PFl6QhBVQwVVQuS+8s4Nl0QdmSxgYa
31/fl0k9W8HC5BIP3XTWAJperufK8s0JUi+z4IPiNvJRtNpz2AOYinN4qZasXyt68yFNjZn2KVlb
Brih4KpotnksU9XHt2F7szB72aYacu1I0WFtfEXi527BSDiwHzlI8Kwfu+R3dxEbC0ausU5Z2Nxo
N4kzJvirS9Jcc9sG3AVCoZdX9Zj3utWeyxhn6SfPnGKOxkzIf34WGkI7M0S408G31FglK0Y6YhfI
UenwWQTZP27NFFk2BSYv2SKvhn+xvUzPVMil+Il0CJh9i8U2Jr8h8KYNrAyZnrDm5lJqkaWxqBi2
qy6kTWxUaSOpZi0BVmduTE9UkWDhO3vOdGFq3QfZZhSKDYM9aaS6ShSWAkDTKt9PwtKVdb1szzl0
tA7pL8Mwi6A1fSPsqqMgzg5Hib1GycPvAQsZ+l9p9q8Vfv2zNf14XRJ5McLfhR8KD3SgRcxd0Ycb
uk7rbv3NtqvDcloXmD8M5dk5HkXgxekiJ7u/+TFYvy3teufImfNdDvzCy3yNe6/R10ceUB3H6QW1
+K/FMlC19W9sW2ZAzo8i/qqPemD/7eC/lF8uFcERnk2hcr2tnGJibZob4CziOtVv3AlL0puUbLaS
iA64aGnF2U4M7//S2fglUnGdO2DEB9W2jhT1IqOp90yEcaxLdvAiq5f9U+XLL9vMPVzzZaoXdGuI
s5pUChxqhWPLRH3uXhVv5uYzDig5FSzHgXLMIS+OIr4k8EVF3rX5hg4RSIZVhyNbxTtz6+lyTe8e
2yNGWl7a0LR5x1oPHyTfTo8LfF5nTEmjufZV6eqccGRTnxyssaJ8DbpBZVTQ51NN/FCRqAm6Hc3l
6mxMeH8jbqIaYPetL7eBGUJoRiMT+w+/pA0c6YT575zUKRruA81z4N7RJYDVTnVIJUdTqcIbA94k
TQvAySRC/THacwzK3voDebdWzKNQzBUJ+Rq7JTSzaA51KrlvPZInrkOi2361FNgiJLonnzwJtomI
Wh1zpLveTxvlPaCGrdEputoN/Jusz2IsQQJcgj/Mrvt9rqcJ9S1UXsr9B7lXxTZ7PkH/zDyfbDzg
wv9NC7yr6kR3GHC/sY11GZfT3Z/g/6OaYhhhAiFtx9RiiYAabuGFEHIWQOjola7IzJZ1TW5ZNNQ0
bTftiqJDjgLrHzdKkdkOSHxOyePjcRXV9oAVSpPbZL0hGaucOyDb7fbgUKc1NFycrkFzWX/okTOZ
rY8SLR02kj+wP34n2ynDC52nmK3x2NUt7bpO8ThEIjeXcBCseOE2RLUO4rbeefpCzkZNmecqoDHQ
0CVP0VaRnp78Q6xw7ZorJKDDDr+rDTOpFP/qHoe97gOevQAMNChnc30x+rzn77rq2J1BpUqD+P0b
Hn0KmVMhKUztUInU1d0YRbaRBYQXzX+DY9h51Grv3KD8DJCHW2izFABiOmqPDFkfjLiKru3zLACZ
0ENMtbJ+dpLjezCXffogGtxjbk0tbHStYlUFystGM2M+8sjnLTIdAR/Kr7vWuuO+LV9Srn4xJYwv
GiN1S3ne5WoDEfoeDqyvPUH4UUTbQCaHxcUvDdj8DMzCeMgmxVJt0xJto/28Xnbd7k+qos73BwnN
q7KjRoExQMSnR1NIylLlGcMP6WqUauf9hT67EEW5xFsMt5e8PpiQUGHfT13BSzlRBlgnWgR7ja2L
WnTQWjPPDn2Wy56Be8p1cF5QWn3PUbfiLt3pMYQ4a+659jgJqnfb0A93bVLLh2ZoTSEEPI7PxMIN
t6nashP2uVT+Hyk97sL47kU24fo0ouA5s5hzIInGdCDWoIxmTu1cuq0w7U/Jh3GO0sNzOIZNV0Bh
pGeauQAgoePjvLqbN3UjChlV5/QZgW3f3NFzs73WOf9JxjA+0upbH/hdZCXzBDnGFhsTTrMWq+Ld
3HAA6aeJHaZwfIrzM+EpkS+8EHewQNjc4fnyV5HtkTvXFz+qlJrBrKsAcE6YvhF7TPEs+iqE8eYK
l8F7mgfkJV/LZWopt6W/QtBotkAXM8OcJitiOdpJaSfCNAGarqf4XX2vA21S8gVtYLeysdPOp+C1
J+N0UgGGX03VT4FGuXfG6hzS9VhMQsXmzQsvB/VvysHxrNYDWZ7omkChnQIv2koOhgoSI8meHpvD
4w+29iNNhOBM2Vke1WRO/6xGO+4O7HDca8QB4oBc/qJ6Y3tpZy4brcMeAQBb6V/oLo9oZQ+mWvix
3gLa2KZgQx6pARvIzuM/4XzX/bgl9gRsZFFaZAuTL2kdoie22XSEoJsWyT8tTMyMWZ7Q+QsB1ObP
SlAw4UULxKQsdPAauUG4SAOsXds1dRI2FkgwSvx7X64UrtxfCCnnXFtW5kiJOLsEm1zrH0Nkr42B
8ykTwMsdvgQglulY9UxAzUIe0ATLQ6Aqd0NIOSQfUrFgx26C8QhTV9Af2835K/HbjMHi1QRE4CFr
ESbLRfTjIJU8nip/32Ls9JSyy+PwOoL2uoGbaClap9SdDejc+jE7n1EMoF1yW0SyJsD0KQmbw3kY
S5tJROokRXyrc2lWvvwQ6/2sWZx23BRzMRlHlhGoSac8fZvhpo7RZJfEOweg8jJjk94GAaZt2FBl
zqsXjPIUNnaz4UNE3JfyNEYieHmMVx5qUdrjgjswKl+S5M3CCCAhXZ4RQVW2ir8YPqScA92f5RjK
xJSftUqz0bzvIhyO7d0gqVEqiEDTQGv1UuxstgS5p1nyic7WAjhG9nuc6CVCAaCIZDGW5D1hK7Vx
FzjUbNh0ccbl5QM4SGnZlgMqHD4PaYuyJLaLt0FuFomTCY9nEiN5BH+zfoyxc4aMHGOq14saqZBn
9Qi7s71qwqCwiOEB01IPdGsmMa6j90HtnEySMQzdvhnpVYem956pFWsHfp4VGxwWFwOJi/z/TX4N
4n+V/VTXbGQxWntmYf/jYRnUcrzPQ+Xiz45ABYu+8cMEiEH4XUi+1x1fsTcnGiYH4101v/JnHViK
1H26uJMHkVwCUonEGaUO793kUJziScBVq6Pke6/3u3J8Z4x6D+Cwf8XwfxtN7cIBuEhfvzzmGfU2
1ltkoF4mADGiTF4op2C+RrVRsqbM23yJp8fJXUqOLPu+FgE8M4vKF8sJbT4IrSSeNxFuT6Ry7qbj
kgzP7yuIr6sAKs8qg8h1v6Lz5jDXDD4QVr9qdvZwTP98L1V3YMTw5qUW3IzbVwgJ5pUjxcpmvf6q
JOYXXTDY/kASixlOrTR6cRk05ETaHfYe1akFKqmYGb5+7LDOjKGcj8ZNKOiai6viYuM7W9yitvlX
xypvEf7us8VUKgD3NwdEWSU5N3cdpjyo88aCPXZwIQTydHNdURa4AtVDtdqSdwLg3q4TjKIiK2c9
X9/Veizig7vk5aMPtD45b6SulBcE2bcYKQMoZiAAxLLoOeJMOukpgIX0sN00Mn8HN3+/zxoBnYAb
D+kmCNQS1PIXs3ZAM+JTL2x1+NQkSh04tlrxG1SRQ466fjiCkOu3TxviEjORraHtv6DQ/UkntyH5
3wV9pptPTexbWlk7AL7XZnX8gJKIki/rH6yNY7+Gt2VHhvJKIvOBCFmWM0Kv1guI+qbycjp2RRK3
GMISgSfXOuGv6m8A8MMmdB1+0760DAJAtn/hJgLoZ0E8jABAEG2vYZ22d2f9cr/FNhzpZ0C6WJwF
hildq+jcf8LCk/falzw6n1jCFVl2axE61g35udgS8feHMF7dhoduL8YL0M3OxII3nhE5YMX8rDhh
OnMoUGjvJj3T7HlubKoMlxuwRL0U/3w9Gnoi/ZjncYDo3piive26bXjYFWBX+djupKuGHyriq867
sGTX/rq5eM4ayDUaZtD94vkQhPCKN7+M89XCoYI0J7/0pPyFp7VY1sJyiLJJIjmqTBhPaO01Lj6S
1OxGPlXkrm8gEMFbQ/8K5F9yYdjHbJcfR1ipNq9fVAUiObpq/8eB7D/PdcQkljoyTXIyE1pOn1IY
Q5y+eZ0D9RtL0jGxWTD+hw13iZRTTubK3GsE6YyFUS0KaFrAd+MogeSlvrHOi8x/dOBvLPxBRX3u
K+87h9q9t6EW0ZZKadFxDcsbdJHPS3KWIRqJiKYIF86EU0tNWnZTW1W/J5XYnmUm3RMNKgUh38zT
wckiIYzz29a+D6b7/R/O3v5+89RtLlzQ4WT3ltOzQ0oYez/NhOz/c5CdgX5UHkqEwTRcjkw4AigU
d/refW0CKnS0zQrUMi3eKLNVrFbZVOaJKMreGLWY/SC0eMJM+PecjqWse6PpIaVHGKYRjhxCmOfx
h9u7NMTiTQskQpj0eXt/aPIU3oxiTV8Wh4NsR9Kokp3b1ZivSaaCjsBBOvuIwPS00jI7nuYPNrhq
AH1hONxaah0HivX9fREXzSlN+em6P8y4uZtRx1dUVtHFANhv7Rc03R90hjeexkR4V/25GGaU6qKW
xZETC3u3uHhl4IAN9KzE0FrmuA1/AuPhJ0l4qyiWfjbEdkBx2ZlXonT2Ca9JlBdI39c1+MN5iZuV
A7K0GX6aSdPVzVST4r5lOVJ33fMEsSBtW0hXkxXpInphxzOc0W9Vk+D0gpz+V3jNyz46b/Yishx7
Xt3NOSUjtW7mDsSjJdAImGl/9WXwlTXMmOPaHIFS53uTDlqJKQ8DgktQzGWlog4gj00BGdbXWPh0
faWrqo4OXhSVkpgq37oyU8hPzD/e3Up8PFarFafS3oEFtaGipXuj7t8FPxsvsSRytoL+fEwfvJcf
xxTcywhHQ8LtY4Jt9NZf1rbnTB6RL+yGd8AokU641vl9JbG51+VLzygT7vvVevkOMSbQG3aL3ahq
brvB3mbwCio4gkSee3dbmBtIbAIyWxPGKE2u5WQNjASYHO1aT9ciouH8Hw6+YtdySJ5f8WeVaeii
zuRz8uUaxfw1GRXNM0daFeJNsIm7FgdqudnwrY8Hssd9UrJDvQC5/lE58RBduODT69sI0HJgYf8v
/Uj+iFHWx+r9Kx4xF5dU8eWIHkTrF7iJWsVUe3nqIacFYAXHj3b+4pk4aQeTaid+bh/OvcvEoq2g
rqBeLrTvriVysRrvmSVZaPDODLp3tYXCzEolry29euxIOuQyQFkaoc0jEQVas8ONxdQhHm8DuGvZ
4pdljtgTJKg3midRz//ydyxSaweEzAQICpiuWW0Ag5FNWvaeNJ0xUtG1kgJQZaMM6qWFD4hLbGXr
Xky3bBT3N5HNkjbhXBIXEviD5jWpQLeCQUAX+NxoDa/uwEQWhviE9IDfl+jOuAYauyR2RDJs8fWE
qIKPqJwws0U3QJAclVMd8XyR1DHB1BoMDxhH1ZlCYPMxRXihnQCCuEXfHM8RC3MFIXzt8nm5y41U
MH/2wgJRxXJMTI5F2F7i+p42jxgR2TCyinO0XIf5YMWydn9Fz9rm9rGxlzgLVWmyX+vMUvqivpcj
CYhz5UVQ5sl3gw294Swnw0O9vJT2hTC4Md2HZcN88j+A9lbS+bJJWHhW5HNf4r/aqsVvNY8dnJjy
EP/u9W2VuTVHviI2b2ekQcUAfANZ4aPVlB0vI8+w6tz4PLW7xrfvRVNfIdPN5fLabA32/qM7tizk
pQ11+9YzV8phuGugV9MkLrOfsnTMN9uMmbcDmhnBoGVQWip8r2xTCjlkiBOAPaJaLZYn8C+8KeMv
mYlBanvnvn2rhBZTY2N63I4J3VOTtEmvixRZBFsfnNwKmkBLY/g9vKQ1kG/gCyfmCudrsA1pOMvI
SIFdYchuq38ZvroCnsHKIXtFqLlYFXR+XW7I7YLknw9pSy5u3BCi6YxGjJiK4wOPyxdebWDLrsmp
BTUpx91BR5UBu55zdfPE+y9fPGBXkABi2u1WMdG1MVH/1x7kx0PqcQ1BtbJ3tA6pMTMEl1z0akbP
4jFhH5vRSd3yrTffx8/aiWc1J/aiQ04zXnI6Gc8WSxWlWyLNyKA8XIx4/IkIFq2DeOtYcR30o29A
MnhVH+Q3pMJPlLwXxHkAWcU+TTtjWT0F2eZ5moHKZHy71JeL4U4J6mmiUGl+EkItW92AMjWsJqRB
OJPifa912Fm3qcBp5TnGFLw1uCXr6jnbS7aqkcu8Rm0Zay/xLTmLgzUh9XUnVIzyAAl53SvukORG
4pH6+DemIVLaERm5oyyKclLxNyYqIupPNgtliNMfsQx3YZdT8vUgRRP/MoZGitM5tQyy2jfnXhJf
icdRrtRovmKEI3JpsuWNogOONqQUA983F9MlX8/MtFO0qgixVDlT+BGNhHssCBSzOAyzurQa/fpJ
e+3Wlq5yk0d2nRuTJjLGEjtAnq/UDTTfW2saKsSl1jclXvJGxC+3ErjGwzoqynEDWdSVO0kZsl7Z
sUcn2m7GcSW3QfMLAg8FPlOpPMU1nJiTolNmcHDRBe6MkbNXCN02oD0thjai21Hc9MAPCK6QFtin
Y8AeTfeSfAn/fQNid5l0oe17s5nPxKI8TuzBfqksduXNkVI1W417JjCAGqV6y0xu6l/AfZ8XkbuU
WGkOt7/BWmyxq23cJf5ifqw59SfKO3DwzW3iET9Ts9vFxAx2cBt3swUPavXBar1Lw3Bz+G5z/tDW
hdPLBjlDLmM7JvnTYsKlp8Kce8BPjiRZ6TfoyvYZFEjX6aqX/bIFOeVNtQAi2w9FJTlr/co00Qm8
1c4L3Znop+OkgjI/OLbqLDquxB/S+JYfcJe1aLR97RQoSsj0f0G/vazy9eodNjlmUKuKG8x32MSy
AtUMw0/vRTqH1VRFIDCvaYkPTG+9u17DUBk0tb1VQCouadzfEHZdBum+Sz/W4wBJfJlWWz4iVNfo
Ng8qwlvCbIbm71TbK1aNz+77zv1zMQ8Et2c9+EKNVZi8yPETnUDA9D0xVvPqG3Z8VXRppX8GUm2h
U+ekzO7/YC8MTBu5ud2/299OFAkAdlZ0+6Ob9doP1Cd0E5XRy+X/SKAw+VLjko399+b3vSHIr2tA
l88n7H/ko5aEUCtM8oNEDX2sVifk3vVNRJuHgKopQ7ozj1PZA2ICmBZUNb4QVnz9li+OCyjGZwSm
DajBAPQqYo9UvYfZ3yK/YhRGeTaCc+Z1xF2qmUc00c3qQXTSbEntX4lIbPBhAVY9k+mEdmH35HSo
nDcqzSTPcfHHtdJiEdBz78T0ufByFyGIt7UDOhZs228+M4hj838ZeF0rPNhPCx6BpnD1n+j4xyNG
niw63lMJsAw10SzuxagMgXi6NHKjko1bM4YbJ8IqjtCGBoEZbZQTizxIc9R+AHbuL1AI6B66LXxg
fSNiK6pM4atPHTxczOxwMdob2hvYGTKW3lv13Lb5OoVJMtknlAG4uX8Xk66m7zDUo8jQq8jpfQg6
MWb0bSOSt1gEDBhhqX7GQki2oKFDP7k05Q4HOCfnGPWZLgyDr93HzKqRpmOetiKDlGa6BsRwM6/o
GLNb4PGRnhcK2hqxhPBt/dN/H9vNj15kIh7fmbJuxeHbbIDkvVK1LzbyTUaCLQl8louUgwuuvvgF
JQRfAusLhoHBd6z4qaTm9GtVgeyVwV0K9H0Ra5/+lNYTtBPjLyoiawQT/3kiDgeS0jz+84U63NOx
oGlICnoGTtQ4VFLa+dy/7lBvSM6/nQyT7y4E/LXDS+zZIvo6BT9VE6QhWpdR4WssEVN7/A189JGR
q4jlb3pApDYeYA88JpCwffPyZL0TshOXNq5Wr94mX/JoLaFyTkWffI7WKtX92JN4MLa5qYPMtPkM
T9bD8p9/ZOPOJyynxs+ic6f5ASsE9Vj/5CmETJxXmRvoq0770U5I3rsF30Bi4WOsvwbNDmtmf5e6
vGC9PVZn7kp+8kwdvDPF+uisg90005pGUmp6Q3XNfCKrEv/mWDod+QbryoyFpIaQONTup/RP3Ppp
m8IBZpejcfkyiQYQnhr7MR02iKSdBZaSwOI3UWKhD+uo2y26bI+wCbDYxuxKngafA/JgAVBZKQzP
dgMiLCo/oIv+V0UOddkst0mgtA2b+OITtxxeFjRwMoJ/0Bi5dwy8LjzEqVg7YMHQawQoUNpqjAh0
syZHlm4rhCxf52g86Y4xyMWuA0wInOqnBWEdVrTjp2phkIGsBLGFwDvPPtP2rHTxJ916s3eMPubh
RkAF24O6+tUXHHORWP1WSnhgEOCyy4u4tm7P7w8sNHu+5S1nPtpl4tPr8fIHjYEb8ICm8kBv1mdw
7BW37USzxQmoPw0aeF2QhTq7ErVkaJPSWYSXJwLyinIy0OjGU6/p7/uXfNl0HOFYL7lE4Aiish1s
lJfKBBwmrq/KrUG53xVPVMAn7igCsoHqKXYQd/m3MlCpbqcTh7qQmd0V7ony/AxLE3hmToyfysX8
ss4kY2DipGFqtfeLJDczxWuOfVtN/0vh8WyLZIjNDsiniqxwStSnZPnj7bcTvD+I/yslGYOheJRq
zLp5qBVal9F7JBb7TbbEkx5r4qNVYzyJTxTJR/DL4eZmCtX27v4rnYssLT3QILR6aBcunTeeMD9E
gQx74x3SgbsqoCeUYqizrdE7EOZackd3YEhQm8U6q4Ux1Fdzcmvinop0EwlAspcu2GfwFTAdhEiw
giWnMhsLY01PYHo0HeSqo93QG5UkZvtT4pUugit/gbaqSwmz/nqtbF3Dx7EciYoEuag8VmFfcrbY
y+rWSbC08XpiX2vCQswJOqFGdjvaSFfykccgDbUMQj4ggqctnf/Jml/3jkbmCclQynDI7Xoszm82
2lD6CfDDJ0fAWbZIuKj7E9u8aoMTGjtmmLcF5gNpGIiE5thehTRliZYL1EpBtvE9/kEn87nqm0Yy
xXucRGinqoTB7Nm6lbPbsTnEXnNsPbleSCahHwz1JrFeJuWkaTba7Z5VQ5vCvbx5rEClQLJ0qxzS
ZIVoWTnHl7ZwGPDxzvQAXYzbC4+KegaGbL6bInOvN35nBl5nWeM5m35XjwmDnvcitEEv+BzfQd1m
BvkPOGRjUTtMi+YWnnizfJ0w81TSakDBVB0an1amng4Dqm/QGdiLNTPkqukmXl35dhPCTQJ7jfbL
v0VV7vE13V2XZG50gEpDyD6dJxzm4fx67dCYMjY4Ue/XCShg6pRjtTxoDIeOCzP2ZkNd3ntdBcNb
U6fYQa7uU+ry98DVxJ0z7kClMetDD71yXiDtMJ95iPNEBW+/I9Aq3kdV4MNbOid0662XKWoMW5KD
lbtiBo9JN1trWoFWzFPs+gcIZOs6nO9TwF+3XUNXjIafkf4yr7+0b/VtKwVpy+dJE8B9B4lszkIP
dXMJB4A7APVJrkULi9ce7NTDJPhik4KQFb4zQxN/7iN2JTw+5ZG18fw+sFDkW1XJzxYahry125WA
3e/EJYpe6KmqZLSsRQqhjzMy6tg2wogJ3i0EJTHBUgQyWivP5k7s11NRDpg4a80vqeK4BlvpoYKM
GxA5CcNLJ00BgEFG0EJD+ZyIv2K+WZRp068Gznzn3M+KWDIkLdvoTM9wK+cG1PsCjmWrbymqBDOv
ok2JHmkt7UyVPNNh7wcGhdAddnhIwsZSzlHeV31fEvZ+aCgMzR0Ck7JmikgPfq39+8Cq+fX56omR
B2mZIKnJF/roTcVP4iqrOltbCrNwVCiticIS5tOF76BF7OLyMwe7OcKs4syICSZpK75Y/zod2XuI
lWL5CmPZAzjFLKwQHsRIksyzC+FXsX1/fNqEnA5k+vKgGcdhtnhfCkLzUsRs3W3avp0czid7eJnn
ccKWNY1TFcHmXm7Ip4zq+ttAIdLf6oZeaSxlhaOp5nOyIz/YPWiHZmjzB9ItmOHCBK8Q9LhUpJNN
ywnVUxWE0P27nGBdU3vvDBrw3NaPJMNP8nh/lDD6rzJyRxur5iS2sJcfdgb15PeuhlGRrZMWCChJ
Amp7Qar/am0NMarcKmmu/iLkNosNVrmNOYJWI8FMR7/Lrvh/oTYqg0VJMUKziMcgO/KRNAPNCabO
/dx5k71D1Ulz6+yCh0G19LoyK6iURQ+qd/m2zBON4rRLQZ+JvSyuqLzDq/cfhUUmkYQ2bLhniBnB
YRMAF9ZAAUz5iXGoMg4s4/2twRQ/Kvv9aeGEX9eVz2RwBuxjUUXX8+0Af0NZ+jk+3J6gha6NgN4n
J6uF87pm1J1wy6PyMWPEvtbTQkNWYt/vXBvBvZvk/v0tvECDBPVsuoNzIiNCT4sqbvPa3Ee2Qyka
lRYckvRbneIjaKImc8qvMtBg+yJ3fGwtXqxfYv9PcUWby2nYI3/zPIhZBjuohzOiCv+IMvYX5Rtc
lDMNjLPLeOXeNZq96Ya5trmHF/4WxlZv1mNTw7IblguObIHyDw1bg2tDPBHH1Vw9zATLGPgvccVd
CdZE0vVCPKCMR2J5xL1+xj2ODC2bn11AWcHKQWldcQcf2Dda6BMisUtpd6p/Bl7s9+LkbV6FcZFw
wUp5tP1QSwEJpV/hxQzun3KWolWdMlk/cFBLXH99xF0zA47Bm0Si2lScujXbriDOubKwQ4pYjzs0
v99DClRW6Cy+9C2nHWB6zcEr3i2B9HkjIz2ff7lFDXIooDOczz1touSPFYnlUvmkF8mOxBjqHLjn
bmQtys87LT4H/ieEHnBmIrYdNRrL5xgoJcknmQnYP3TTysygnDyLJ7Kne9OkP5VM4drqnAMYqqUj
Ot4KLVPk4LxIa7q24QZcjeHYwR9s04L0G/lI9ATa4/EOslUrWucAmQWowaFeD7vV9wuijkLNFo0N
zKPZ8zgqDWsErN0mLtawCnfJPif1Iua4kOAjWNuFdaIdbv7J7ogglE2hk2PihubaIdz+RdhVyas/
K+K4two3Fzhf1djlKO9jFxUVuUz7LNYlJ3kXwd4wEkF9TlUaOBqyzNICeRON28m4ynwGD81OQNbF
SRFP3lANGKRNiR3mO1F0XGJdaQHjCMD+34ROH13jK5oNkq/Gis8eGeM3yLXuRBBAC8SJb8fPpZJQ
cyDkSqeMKVFTYpfYSUBTkOUUpai/jo8wmWJam5/jqfOjR4zfVBdZma8Tqd1zoMZ2txpxFao+p+NA
EC2lFbYVRz72SilnTMXnA71DHrOShQbO3ljF1oxB1NWGAn087eKMkzKjfyNPINfLePEq7szmfexi
zD/uv3uJPl0nlAl6qpc1ctTVv2/0Ds05jsTMBMtt5dswFn+L9bJDoc3H/34v0Tufv/6NVDTOe689
GdnyrTa2zSwRcp8F1jArH6aRm5IFzrGXbNH7bO2V9zcRCmgRK6KZmGfcnof97xnYfgvGd+VypYYE
f+hAhWvVQhtVTOjSD//MIZci7EwqoG5O6PLlC6FtkFTwi2cyWfjX/XJZJT4mumwoBhc12z28ilRu
8ML8C5QeoKuzqoEK8j3TTWFkxU6rJN78iQA0tjLoMQmLYgGOPCVmVY9hKsfm9JTWGneo5FY20NWe
ac6tR79TDgy/fH3z7cda78YKv8l9EAWXAynAuiSzuP4aZ+5cVMbZu2XjRPB37BqEbPgdvEc9/fZs
sBeCEIvMB3iCcuC2hYF5hYqEzBibElK+uzGL/BmfQ0gX2ET79bxC5dLV8PJF0fSe/oCnbSa+YQIy
RjdPyolBnuGSxKoLMiRVLuSjXighUqzI8vbXKuPdCfWaqovCk2dd4Y4CPpQkpEYPn1js8FVyULzH
D1cpQWwOoD37Ab1fB5xooOOBC3yby3iCha2U3rkUaluoCiIuUreTQ3L3YAmOVPErt6iQDC92DqyS
+98vo74uUDKuilHNU1EvPhuBXBrHkIJo5s+Pr/slAwC0xD+3Rs3wSVS6Yu5rU+tp68tR92jMEMxR
pPHrI+Lw1RttDanCDlLxQHXhYBkA+CN8Jl3NXykockCoKnsIbwSqCzr4xoNqhy0Ird5KQ4SdU0dS
Vh7JzJVI7tFnM+4/CmXaxV4zVIuCb40L0XHaA4dNfYx4F1AHn3Aqup1u0kFTMAqGPmZkszkExDKj
YFt3ESZTbid0Ifw98XygmAqcgT8JLRKU88Yc75tA0K8VUM+UsVC3ZTfA4T+5oYQ6yQMbGwWrpN6Y
+DAJb7u+beuBpWh+uexypreUdJzhrLYaqx8VGJbW7BV4PrAgScjne/Jin91dlWOgqx4glPt7IoJg
srTJ5bfzMcG2k9gC1UORyboR8fHy66bXByYj8PXFnki2bWMJ/M4QGoSmG6227IQ10nPIMZZC68hy
djz0e6KqdFkwTCwaFj2jhL862+aIcwKlpcXbhWlr8XMKOtxrrjnFkM3lQ68I8R21atQz2gEVt0ka
2xoQ1vd1ZArVH6kApAsWd8nBRx4B7qU6LBVVE4xGyBxvKVDKFu0HeVw2TCTd5THBY6rxl0byskrL
B19Dn/KIZrVuAkLKTxL7pdZdctEBuN65wsdmd6kDJWFoGguLbjDRYieqCZZgZpT+WipGzqElnrOK
QDIEnUl/dxW+p1FV8cGgmUi6lyo6RWPF0zZBtL5VNoRYM54h7+yQy1peQCDd++6y2o08fRa3y2m3
pM5CvUhob15Cjo5u1gz7RV3llCEGOAMi74flEhBN009s1sCB6CEs5xJLpHYFrFvvvenvGEnYRjOi
Xb7UTK3Qv/rtvJjukCAJnJB+WFGvA2C1RqBEce3ATDyuCaQT2b4Nz3o6Wzoiy4wmaN2qDyhaKmCQ
yVQwAqatbYgrmzlcEfi3mb73de/FKUVRaA1agc36SC5izG0GFJb/ScmFKkpCKUABxl0eu91NJ/OZ
iN68Aqf3ND2GOs5+SY7z8hPoS1fEvEsLkRMcJrAbw7/UttuPSBJ6HAwlkx710otG+JpxyWjQ5so9
2bU5UT26V3eZB9kqHqXctLq8MQEwbtFOIlYvyjL28gBoQYlC7LXCES+sB2EZM14XDSAqxgU+1qpk
UQEmV3WeAyd14ETV6iblnLGRMoXkWLXmAsP9EJf+SFaVV3zLGbMLmOUdwGIfggu/WDq1jTdf1qbT
ikEBCUPGRTksLm/Ebt+lS108YNAewiFKc/xtylnLilU3RNglOgGw8qcUljln5tJIlFDSSDEtfQST
isVV5VufSnqEuFfkazrXyfqeObT+SYBkqhAMwSaPjmUr2zogQ/6EeHq5Ba+ZeOy4yskmWQP291pl
iwkWDR+gtUcS2Z8daTQtK1APprQX8dTRg2NetSS+GsdNGWIzTi6XeLXapybyDonYb3QAMU34oypZ
wV4PXYM9GLuHPwDlfrYgBDdO2UHsnHNXBVtJz3B+d0DC6ivuydxKmVgXJz3d9mGGqICz4zK8o64f
M5F1h5hPxfOhYdVMSdzgGA+Y/Tb5rz/yxaqB8DrbrW0P1SYTIL6pndiNyKcdVXHhVM7YVDnjn6ip
IcBs2GsakFJmrxbcdTE2BkPHmMjY3MPOJ1tPqUYAR60B7QdwqijoM9l68FvU31KDbgOurbpafeJq
oRLUMwlcUdSPmsJO4h6iAUXrqKJehj5QOshITVdgecI3zj+L4MgKYbLaaWF6FFlpIBDOCFmJjk6u
f22X0gTVvJ3DAKDmZYSH2vqgFjTyd9EK577+kIsYod0+FoWq8FLV5Fb4SCIhqX1F/xAFeFLM+ja+
iu34lWr0kOI2ohaoqX8ItxRErTr2HkGZOOp1ot38XmyZXdL5Q/BUqyxZpyX7QC1uXZQ4iX0q7TrN
eUiX3YrN5jMgBYODU+wkRXr5YdHmaGJotswAQ4RNj8vusoaWneJjgUSCeSUTJx8+LxQibNkABfSG
sHe60lmoJpNs7AF4K6Lgj2F/wC/s9+g8jloy/mp662wK10/m77x9Yki9QPB7pI8sGKTEpxqBtuHO
skD4Wv1C9aYHv7PDk6HESgZsyrv+kgLLaPVIjGbnQw+kF+hGMYBaLbcB8XgVNHPHUeKqv5z+W/RC
81L+qwskXVpmW9qDVrz07WQ231u0jg1qqI1okYuhEegBwR4YmLnhZbl904iGuKVU0YjIkoBxmjd+
juVg31YZ/5AYSJA9ufuBLXA4B02KvFuJtoIkpByYhiSFbHd+JJTd0LixfaTFr6GXsPJEbsYwGj9n
qS9NNFIHNcOOq5FGkvCjnznpD1AFGsWzOKbv5eogoU/3y19IAC3uuyvyeNLQr0Gf4vAmoeRVvzG7
IKeQTqaCeXJQNkNCcPSZ9j34rd2GR/3akmQkkmplQ/YqWto5njqSUKzI8RRbI7Yaow0hPlOgCeaI
ea9Ew2s38dzDN7U5i4A/cRufVafWY/s+0lKp1bPcfczVWReyf9vpuPb86D66FarIg1ZPSv3i0sgA
Mqxb4b2fVwFDm0taB2Ji+R3DtEc49YEkzgDUA42nSixFy1rWMmZiGWk9nQp+dS7UULpWf6oJ97AH
eJQPkCeXnTCP0OUrx5kEJ5nCUpXgMV1+SyoHF60lhpsEzI83AaDY1unAyWrZQUd/dgIVNTnHWd8j
CGDwBNv+GFHkjWgD+28X4Lo7AagotigjNtv5YA/qWRcvrd7dyfoRv5HJZnzMCvdXrwG++VU3nKnG
/2eEHEi+Jv6DJAwhcoN40Z3DfA8fF9/OR0XqK9BpHEV8eCVRELeVtKFq9sE2iGFbYg+oPbq0QXEX
Phh4i3nBdo+ZpdNG5LkydKlY/8kSQxZqQ5FeLYFHKfsnhJMTrg/Yd7eaAdBd+Lxs5xibrbdln5hx
NTPp/PB/HSJhJHmnuGUBLZKcdwBp1wWkUPI7Mi3sFRXz3VWvvlDaVSgvEW7JLQxb2EKRIXRGH50M
Dew79mEhy7+aldc33FCU9Zy6eckxG0m7/nBgE/V2kXtthXzNI5LhGMS44txSUh3v3SPyvQm95UEp
23hQ9bGBO4W5bXxJZm6tRFUUUNf6FgdrWRdPOYAppjPtY1kmHTdC4QzQ7jXJomTHqBiBjwbZdMQP
bOPR5mZW4/jkse90SGabR1fMgD91Bb3gvy2oVi+xtCuucTubrbeYEYfY5IDZF2DOgqefDQR71wtA
RAMmuewV/WytJBA+LcC4HBBD7Jj+SleIz6vuCDdE6brbzE6BzI+5aRLkbd/rJAW+BzzYW1Bp7Rz2
YKZSp8JKYJ8Z5NEquQ/rhsNosXxzQFzd/dgxu/7MHYb2qHxZiYgRRAgqKYB0MNSUO8Vs29RZbLPj
veJUcFfzN3/GNFw0hXt2FugutI8Kb1JFtEQFcP/aFNkVCsd4xltEF//SEdGkcbhfPl1EWegtZHp1
YLy2fuCht6wUZSmyvJIWZ881ttP8pwDrP0eyipCCGAxSaeW7bokoSCP7yPvYdTlio26JmdGvY5af
i0rKlTvC1FbdpQuJNluQOmEI0PSDkvo39lWRq9XK5rwDuWDZOqw/JZ9OJmqnxMQw7J/GnuUncdeR
e8KTajDsCVl6AZgrAAPQHmlOg5fgaIRL90Y9uVNUf9PK4Iy2VKFvSH613rB8umWoxOrLPv0/vBKc
3ndWsPTszj1/erImd2cXhqBOm9VlPona4JZP82iN8T0ScGZPGBB9m+kbHynDtdsWs6ZgbVngRJp9
PZbm+Oge0FnbgDEMP4LSM0Ski/ygKSawBFlwoKoVk77vuWzvtLBBd6oCEtTU+1yZBTQzlROc+Ewy
FZEBSflDydvKW2TrL6ZbCQB2dafWJT0m2/7hupsyXaK+34Q+oJd+Qwua8gAF7LfeSGSr5bVVraN5
EHj+LBUr+TkfP1+UKqMAKueXri+24LQYJz1+yv0FawqLgQfI4DRoRutoFatF8zSVMUBuvbKx3nK+
uyGFk77PegqE6GgtKOPIBcd1wP24qwK76Mmjflmz7hfzrLAclntGvJ7Vv067x9muDfb4epOzn7p6
E5K63d6ekMDpqaMuTFZa0pt9sXpUqHqBL6UadkiJ4oDVYRZB2DEUo/e9wczG6NprHdphQ19AU0bD
NbSr1SKzVgE+qFBSR2Udt5xCjwLrrqNB3ue/YXm5RRjafsmGd9dEQ9Z6IEh9L4aSNb2Mw5j6Rkax
ijzZZWA8PKkG+AbKQeQGCORb16q1jbUOnMjRK4QGG4mD7JcqRc4cg5BruGu12+9k6MwNQRrEiSfk
ObJbDsuU0nnUQb8m0bwAG2uR0PoualCzYmDGROByUUc7GmlhaDD/1vHafw2dl2D+Dh2BInnDIPIx
T3oSnvp9MNh+BtgRNv1pF2QK7mpsRIPLorx7NDWxCf1cifSx7KIUY6Yznv1p0n/PHVR/4ckZrVgg
jj5Abz1Yt6kbyPU4zHRv9uNDyVhHIlYhmkSMSv7WtK911p3Q5wgPg3sCOBtkaw9/vKMMPP/EYsEX
OKgN9goXD81Mnd3ieFyshNY5sBYitb5iCB0xlDY5jtXLEOJHWZzEUb1NS6bOG47JC736OXVxgqLz
ZdlzfvaRyADUAzgYJELWqBcqVriPn/olpBJmVT2yWDVn3iCzy2/GouEYo5f4ygyCDslbfFCf+ykF
VTFsJeDOECbmsyoDAvrs1/b1CFhyTrThr9cn0WEQaVOcOJLZc2ETQRz1StB9u8Tw4BOAZLtGQxLp
pRqlrjHgAEaxUwJXvYCgt3K0RCor/fxouGnYThHclgt2pf/ond1e3CSSatiLFNOD6q8wsL0P06qq
4lXJ2BvOwH42bmfNa0AH4PGOGrnMbo9/BHhUVv8yl+MTndWgFV2/Yx78BtrfjyB+F5Mgwx9Mb7ee
cpjsq1uIOY2GKbDXYaTE8n/SycfQDy9TGxnXzjEHTtA59bOUi7IO8rf1GhLdlAfodmEoRdgh31lv
ZiFz9N4QgzL7Rkq6TwUfacdovtMTDMuQvwL47Bv5W4DKqL+BugLZu+Z7fGCC8QVz/tUByPmwvpQc
CRi6H8/Y/HS7R45/khRA20JERRJkVlEMjYNMd2pnSe2PEST4ZFyd2fw9TTzYNNJRrqm8T5b6c+l+
xxaVEUsBWEGLTIycg3ySlzuI5M9EVJmI2C3BdH0WOPRwlO8eyVZ0NK4rEYy8kh9bNAsEw+qb5rx1
W7W9eNrlWRLVfMF8p02ealK0nm8r8s/u8De4lFMiIibAadJdX7pmgySYC+dRheNn7zBckEYYmqZD
GCO3EGLJJ/bSh8Y8N6IUh3iqVC9VzYURO3rgw8SzKHxlVlnjG0hqE13Icysf4q1x1AZXq+DmL67W
mhBX8tmeNofiX30/biMisn8sGfliWXWTTh/hO0tG0IvVeWTN2US/GgbaJrRSafQ5xC66JdiGn3x6
BfbU7F1BQQShtHsXIrOA9HwkIGXNNXuNyqDVqfBB7xzhE1llMXquiKHTvmpCRNMSMo9hkgg/hKx7
d+F91pPSK2R7Z1gCT3YWXVkwwk2pXfnarploXaqUgsVBUFFR39dDc3HhZ7scaeZQkF2Bhk92+mba
Rh6qbiGtm9EFXr3e2PQQA/9EvKanAwe7CPnJI/osfxP/F9R2srOe3HtOMHpnkGyLnaTgP1W9vH+s
Iw9hG8rD+xVCFc1xJo3R33qYiPNLdxfsIJzmPkeuikE/eoeTsn+l/Qthw1+SluexWTdAviCNXSqh
u9dNzK8z69p1jflHBhqYaLsHg7KTsZ0a5oKDyUYYqHz14o3bOsHGEjeglDeS9AYsAwecjucF3muK
LdfvHA/TVO/eSAAceWv/JoKJmD35j/IJp5SLa+k33vmCgSjMJpe2X9Df9FvYLlJh+rPJB7xTlLEX
8Xc4Eg/2X8IyZc0c16u/0iAwT9Bpm1FHLPkdbFss0K9dViri239pppxNQuyGIjUj0ZGC9xn7pn0V
iVb61pBb+dTUpDoom4zVk35iLKkKJQM//voFQ+OW0UXgfN/qxgowqckx2EeqrGWxmQ9EjAOUTxv2
zSaXtlgBS+3RKkzmKHqH3Jk2hj2WQGskgJ9/KvNAfd6wt/1F2UEtvO9QzJkCtLeRfuf5HztRxdND
EECkimtXx8jcxaUxe+UpznuQqxh+/hpi8W7+NEAvQQYR5A0fUvhrq6dS1t/FByZ37b/6mBXUwUIi
ulWx8eZTUF7R7QXlER034l3OWlo0WTSs5NPqiftPquBtLDucn5XQfZNjk+Iew//6/5mbmelujVQ6
u4wK4Ssa6mbn/nsWM9FWDqMjYBS3a8UeKbp+/pvx+YrcifJxU2Xy7nbP3IyXdLQEVijIjU/+k6sb
TnWUE+DA1ZpndTxr8MkVaq+nX86QThB/qceIUGbwlr4Ucnxz7aBRdHL7cPx9mVLpmL+ZcFtgca7Y
kqkTOJCjJeWM5WjBTP/PNFurPoACjr5eLPndw2F/xOi9M1oKL8KWegA4ZC6vcevr3wE6nSL9mzYl
iPy1FxPoR6WSb/VEdTqKcvHZklAmR03IO6jSU8mVmYdqL5ah2HpK/ogV5mVbAda6WbeRhQBCxSdo
mU+xQX6BHxfWqWpuYeiWuY3XMOGcux39JNuaE+BXJD63xBkaCBV6PADIsEU/pn7Yq6GUsKH3oy0j
8Miu5u6Vs5hWlQyhF38MzPisG0ogZI7yo2EwvtHQmxJNKmcNp/NLFvv2MFp0nwzaP4rd7NXtNIMH
aWxj8mhtj6wpaw82ohum5jvQpsRChtsB0iZe3ECvCvits+uJC/IU+1PHXUR8DIIvcDJF0Z24P63q
bjcDGPDztTwNvc66J/HOJ7kR9VKJXLceFNIW2cYQ1Lu2qUZja6lHBUO+sZWVUhvlh8HATe4dN63Q
jONXfjVL5YoHL+sVpnEXuvd74KNIMY+6pFw7wD7kJ8rXpwparXqWim7U8eiyCw4amMMnCTgcORMK
Wd8Zrmgf1gG1uLGP9bXSF5cckbGp4fRok5VwnXhMZ6q3IYLIrAWrjX5cMnxHgCPs8Ri/W2riOc51
C7PbcWH9s5l/sWrbf5biasOtOube7KBC92Ub7sL2tnbbNQMa4TMU5Fcavr0MuvmBTvtYo20yU8LV
ZeqvuR0V2yejvXAM4oOGaCdNIJgcV+WLra1G7S55ow5xB4jmL4HFzdzoZJAuQ7h6JlnwzUhlHhii
q5FTXIPIxoiz/i68iFIKOhzcS+CZsroXFnChBCFU+YjT38MWcwhLlNkkTxnS8DULD9iGk0ll1xzW
wERnhe2k4Bz0G/bCGan3Xe43ASbE3Fi9fOFCYurwqKCbilleEbzZD4opw+AzLB/SLaQyLvXl25K3
L02OTWz04hOEWgkLINPkZOPaV+5SUyd3qGHiW9bKSONOpGLtNTyZcZmh4vYPJ1UefHB4ikHAKFc6
wR5h9vhgO9OM/j5TqCsxL/AjjiVzJC+tuwHesLjebn/OAbGHNxSMPzeVsnc3HSrlK+foREVilLZQ
OEbJlc85HCYhuOn4Z8kITV7fQAjiEN8AomuAc7R/tJYzouvY3PRi/Lg+0KLPQ1BTgfbSizAojmDT
eC0cEhbv0sMlC3PgOYrKmG44Ml2HCOUhSTGACQfTgF68zHSF39nhjRm47/6UvFQiL9bpqBlGXdbw
1Y6QoWSxkaEN6pdD8ar8/6FPrBEO8h16p+ByEpWEEEV62LTXxCcqm72yhvoppQqa/4l9DphlpoEJ
DIOSsjehIz7uNecQIFGcm02LS3AKC/aVo+v1STKRqLaQWBiEYXfYCgslY1a0xRD0dhX8KmeZu0v1
RhiPmNdhmfdeKBikeLBODpD0CotYWlbaVuvNyYc0AiDTeM4pk9bPQsB7OvI2Q9bZ1Q9rTp0sdbgX
DMNp05QvA06wfr2DQ84W64AjYuDKMHTqiAOmKOpF1hIn/f8lqMBJOLLvYBSgwCHgA23J19kk8yYB
HppZ0tQuT17fWB0TWnE0ql0WuNlgrzk/xgv7c6r+4Z2JU7PcOqRFXeeiuI/fOj1XSFv2MC181JlQ
ZlaBJr5jKFr0xw3DuavOQf+mX7RGTDaOOLAmvxxhKxmdjKImj1qbhNPhL9j3J4zY2yNUSDKLzmC2
kWTzN/NiuYx/Yo922hZqk+/CTx6/yDc1DlCZl7GlkTF+Z0pXyd1BgzKc20i1qwBQSjG9kfSxMivV
nd4VCTNzXUppMfNHazlUrq/dQ9u5VPAmpi6HWAnCUbjYK1UljPtoY+l08cVuO8ov7+c28FxY3nQf
nIeXpHXPag+PTOhBuorI40UT9G9p4q+QoxL2fbrY6IfTKzQDBQWLTLFz+gHy4YSYQUquXf+tz6Hq
ySuxIYl8UauHXYOk5m++vTokSfsKZ6OPyAEwks/FM7JBGtYLcBu8ZqIQHV+jDIjknw5GlpxH289D
bP0TVQJrMa6IC8sTFryrliEZow3NSxjOC8MgUH1cCbGHiZICxcuCSyrRXsw5bpiEwMaJ+/uVrXUa
i7N5Dov0OPiYCHNOF1RwQf8kDjL3OppgYWRNbJWaMeTR/ETGn3LEDEcCgenyE0Rf6MtQgrdtkiTo
hoYuMX5S5B7yewUdV7DGBLtr7XfKPDnGdhWZnJBgjN2zd9wuJ4xNEbwFTmD12cSltEsZx/7XNpcd
y72vDCsvdkraSXQ0iMj3PynQ+l08bb+5kpTNvQR2ZeIO2rGIJ8annlWzZ2/ZHuJpnWX19c1Nb9tk
3F0o6MS0GO6fzqviyyiMM3q5MmZXLgXPFc1poeqQ7uGqNXj35Cu/FDYSe4nXQF38Q4VoGeedeePB
JHLASH2Vc8eGfRsHFiX/SkJRVTbK3bK88j9H11BnC8WukC7yjSxsBhnDkqYmmyCxVXNF4aM8djc+
IWONhxuFf2p8AlphibLOWuFrbMtKfDa+zMOrk/R9TqxehQesTiFF8Ba1To6dga3ytfQnj2dI/gss
fDlsEkXAAKyg7IA4wP2ct6fXH+xhcwjkcANL0EEgQOgWKOdAmjRpmsL7Fec7nKFR8Es5JA3rQ3kY
KdHTqBu4W1zcNce+k9AGnr0BNVkCCmzNaqXcsve2ZOZ+2bUrJ6jz/mFjB4nZ9sFsGHrJoDvjQ+3L
5L/ZzY1QzBBMcr/yfjRBRTatBHA8Eryc21psfNl70cwv8NH5DZzxh4PIPvj6YFPF26o2giyaRKhk
Bpc2s+W8OZmKeQqje9GKuLFBn/BDwGdHuEnol4XWNswqtxDfHUlxzwdmMkzN2mk1g9b5Yv8zpwm5
3RidCVyhwn7O7nyVo7hhZTesEFFPe2Qp/fep7vZLKMEjAdX/r/9z38P0VY43mczTBmCEOddLiiza
JEnU4j5dpbEjVvC95x3zj3bQgh7H8ABK1ABVNHN9jtv/lZ8vSKH+UcPcFAJ4fSGlfrNMTRRhJDFf
qc6Y8V0/b4Zu4NuerTU+dFMjIJM16beONcfRJLpUeN5x5+SV+zSEmbfGjWIk4GQCr0v9vRPl9uJi
p0d+Ij/N4tHdHdnoxJv7pegTqRrtdUpepjvfG+n+LbWhM4RLqFvPVp41GHsj2Cth90bNPneQj2Rn
1mohviadrfH8RXE0O3oEqtpG0N2VVnXWnrOgOyF2ZzUnrNf6STD4QHEHq5gker4uCeGxNqR6sDOB
WdUvubRfVfJ/GgOxK/lThXjSQRkjVEZWgkG84WS193HCcec/v9GGe2c9wA7JXLPlECRHWnxB5p0r
EMSau6FCazDI5Ap9k8xW+a9kcHR2B4sykvaJEs3kiukdoA/IZnLyWLbMo5V/FTzYrsgZ+9cxEtA+
Nj//I14n+9733LgfLlQIganvRT0MiDz+882DbUXI/7XJgJQuWC/B5bX+3L3RIv/NNWfTJotx4qti
krpJkgnoNzOuQYI90h7/Av2xvK4WYon0aPIqhTscGh3vZkiUvzT6Td8bmb/5qwCu3YTbvEl0WphT
XGbG54st/MAtjVGLyUL8S/RnP+kGUKAMqqI9DgRFqMwa4NB+aqSjfUih3z/SP4uZNpvjlwy2NVR2
+LfhF+ekIHH5Byf6fG2YfibdLNPUqkToi48otXRNjmuwHLaMD2pIsOVI138ReCAyAYJD1EXrcW4V
aFH5a3RY9aJJUr0JHBiYjaxx1oAfG7XY4cCwwlsJv9AqHC2K9sXzhVhaPlZ4J9xM/DshvUdYTe7g
wtvr+drMm5JfWEt41v7WaDCASJt1WnQX6JjXFV5nIxuEg8oxyJkxkAlqao8rF2Msmsq1rMIch9w3
OEPa42K60kmtovckf+e3Sqt/G3ktSwD6o7fDu31gUN3zekqGGiegjw9Gli2x8Sb2D4LU48fd6hsG
ZErdapbxeRm1e9wgw880yt6mPDk/0cPCcAYdzEd/6x0hfUNsXJhLq2dROeLlVLywIbiPxsBxhrKb
46et1XukbH92HHhjxOcreOaCr3qlTLT+KEm7RSnd5tHscqQsO/59RcVGVmWfGOsYrDRxZACxZJbv
84cnt2kkhANxmj5C0tTiIntxHJdjSGIndoH+AGeaII5ZHGKTKyDee6JdPqOjtI10OzMl2T0JcuwG
xVi27p/OL7elemsG/ekKUpVS12TJsFidDnNksy5Vf2sSnFpYV2JMgBiLQH8OVSxZxklgOaM2nqRO
vVs5x741BOeXL0G+jUqJH8xAv7I+40w+bh/G25+SCIBgHX58t/GwjpNu579BD/Z7JfW56dmtCnfH
2cOy70JJSU85amAkqWJpBljk6YiwNDJAKF9TEH28YtJApmaiIA4yFliORjm4xeRhVgnEdUsJy98e
TEAP5N7RMKdl+H4MR0YNqH3OPieAenzQtFCSJq5R+bboohNg3bXfvXMdHywVNSU1fmPuWUn/WqsK
dR4nG26T/PSE5ptxMjp6eyqiFGzyYrd/WWSIRPjQa+bcc0+Si9+0Acszn5tErslQIISaKSg995vG
xmCyuP7B6PkR8JT7BBjrRRKrE/1GoYciMRTh+qwlpbM3nceyd9NwLWIX5BurqgYwQwLO0rZnKKDv
wlgwPv3dFFpsn4VN2W14g6BJ9QZHO7nvdR2EcuTe/6FqY1OzkSGL9qWyQkSBmRXPxDQazt9C63KF
oNuiWFUSf55crlxAcWFP9FoBw1YMuWeqffrc95A9nQP/Gwd12MZG5ySy8GZik9AXuVfPfL6aocNO
3TjbHSBgjS89Mm9AgMR5fMCfyHE6h9s2aXtT0+/KCZrUEow6924YM6SPVTjUIXmvXzwXfWfbdIp2
aVOf0SSjb9i4kOQ6FyB7JPV0GREdBa8tJy7xi2yaawFrWvth40n/FWQNXpV3GwKFDdv3stpxgiLH
39jqesu064KiOo06aDKyKaNIQixCQrZoCaPesXk8sMRmJBZ46Wn0sJ7Ji2exmgKnWXxChpyiXKC4
96a8P6AE5aKzzW7VvrpO06rbxmsZQxf9otYXBu66v4WlaYj8Yl1mql1jjLSph+21h/eb+pnmxhBg
bgnEBTarD2ZGqwX20qDpM4pnfFBpQMRt5WDgl5IQJDc1hIoQ573fz0CP2Ltv8a4jdW2Ksp9mMUiZ
0/qsjEV+GV9URLcVl/tdOoh3cmaGU93EVEWsXhkd6d38uB5JyVpnNk3H6buRIZfoKLuNrnvBUXH1
sOWOOVV2tseLM6KjyyQkmRzj7eB1x1KSiuYDRtMfr4vCbluPkfOIvJ7xLXA7aCRd81VllHJynec/
NpyRbhznzoZu3Rkygqt2gHPmfSlP662yIf9TpFy2KJxde0ia+s520BWS3Cl5ik5EzXAwcjI/gvEb
uvmzdakSeEPHN2wGH47sIJ+cdnc6FChK6Us4a+Qae+3Y8RqC0X5aytow/XHYDHyLymbMHkLRRtKr
Pda8gEYEREkNUVYdUKp/SvqrkDzHSWYSdEwDv442bqk8CeQ9Gob/FLlky0VKZQfrwIpIFKD2f4Kv
ccvypAWGNOfJJ6xsXQFT3FVYo15IzNUpXzAtafQh3SmzzZjagcMVVp4m9Whh7gce01PYOYxphTJX
4L1koL79FE9G5HkrRD703WREBCTPQm+mgDsLw2e1XK3BodmbBB/demNBJ2H+KsfxKrgRmMY+D7Wt
T9b8QunvjG/dxKrZA09VdNP6hPqIRpup0214t086ttnImuq8o3tHH3Om5wWLxZRD3IVQYwTIgGJe
jOssib3mmoE05dG95fsa/5togkFyBwyPMiC6BDhXdxentOh0JY5XoCF5Tg08mpTwOVAxDm6Z0EoY
gt5Zo8El27xikKcPwQDmbU3AYp0HhxwKxdZ5Ex9/1G6bfcskXE41amYa45x9HRtkcJWJAgPhnzIX
d0Ga6+1vXRxWRRamUWExyZ/FTEh3f/LymKi2UlsgtTmC+HZSr+ApO3hJPgZhQkNjxr9DeKUleRYT
TpgBthTbOTlXZ2PMChJk2I18lHzv28+DUwLpKv2CN8l+wj3+Dih0/zYoF4GPxQ21PltqH19jI+b5
CIuy+Az70Il7xaIEkeLolX9SRJNK4qBJTRz7aj8aCtaKezxwEjhrf3/WDBQRJABumMMZWk38B5PU
zVwoNUOXlt1fwyLZK01a95vw5S4R8Sw28u44G8gXvqXYjUtz+idKFbsJDd1zXKdkDie5gq4PTiqL
cupYthqBZD8nPNl5Rs005079QQQJJOrRQhvkyEvhLXKk2M2WdXAqTf5FYJYSiaye2w4XAYcc2HT1
R7B4D0xhOAxb82EA8CoVm6fCT7OUXu+EsxbKbh33pIoy2X3DTvB7sWqgBTjEhSLSGZPsM6vTYX10
V5jCP7KZlkvlFaaa/hAkU7Ch2b96Xv2YQHr+3TcTnXdET3JB5cATSoplpxL2yG6lt9LTKr7PMA55
Ni2nfZTXExF94m/RfzFO3MmcKW0rU0nW99B/l0KQ3Q5czNcj1QsrFlSZrRbKOXpogbRmDGrur+nr
Gv4szs1XuiLymqENw/JY3RA1AJRuE5obU7I1Gg6KiDdTFkNZwET8R2bcd+Ka9Er4lFsG8uBfIgcu
Aq8VeAVzxh4Ue8Hn/AbImI+gVYlmO0sU/aXdzC46NQcyHVQV9O+s2Pfk3+KOywZLmwgejdnau3wK
vTQTqIzGKh8kXcazFC50JyJDiQ11iISgQRHpiPfoeJVb+cX5cxy2spdnk8kWSnlRWRjDantwOVnZ
aB/NCkZxLRf2O5cOwN6FSwWDGwr2BAk4/3xTo7uONlpau62BUWYIFWr1GlgSOhuXaaLpFF9WqLZk
hdkAgX2z7ZnJ5ORjss6mHmfKysIuX0CYPebu55RKBJ2cRC/qQfz9I/7Ip+LoS/BSOu9RWn7lrTHb
aWnrZY4PDUiScuOWlJkiSoHk2Btj73TK33dpy4B68o3y/6WfglKf/w+kB2nPcsfGoROaQ5r/McUK
cSh/+/hxsbwzzzRp7StzMdmrSvtX9MK/hXfMDxu8iumMMxpDlWlk6z9S4W419Nr4one9AtpnKhKA
mwK9J6L1NUmGvBWBxlvRuK1YM1UAG1xU7reGWCpBG/9GkUuGXyF5olmAQLpTgPQHJH7r8nb2TOLK
EL/bPwFgz+MsB0c2p5KQljsF5g/W7wGQrPDE8/nnW8zkGYhUoSJ1q7X0a16VWff15pTOgQbkQWcQ
bxNESt0yyU2nIMZhZT6+QJwhd01cXawQ0VgRzmWeoTwAQEbBTW6ZPmONiERzJc9bGYGyTs4iJgQG
55rwQpCeDNi4Jj2GugoIUpZWP+JMkzSwooz+5PLMPtYkR5viX3cXDXbsFhlG2SJAfKofz25qdLhg
NvUzhb2Qd8n36oxIO1Tb/JRIjX6cdsLyrPEl9sTocxEBT0h6JOOwvLv3BTgfpJ5vKjS2tAYH/v/f
g16ocI9IhyDxLP73q3oPWIGh5d9+Xny7WFDmcDyYAuEV+Vp7qf6cEvxSFmuvA7xCgWFmMagp3unk
yEMGH4tFdwDfB+fYu6h+oDkSp1jfRp/E6WUTQr42pvMZFTfwxmhzstOVpMg/+xEzvtAVe7unFrZD
MnFjU1gyEnTUe+wct37WqO7HcS+JzFNJpMOR0YEiakZWEthcCsCJ9y+SpPOEhy6W9rLhP0nVI9ZP
DwQ6gYBOLYCuyY0yMde9h9qWXC17y13oCmXokLxKOMkhRtzGl9EWLCuqCYagk+Fww1Y7vc4bmZSY
A4w/JOpYgsk1lFO5+8A3V5uNFS1B2C3GcLk1O4gzxsK6Tu4UU6fGIEZWhn/mIhdgtyXFym2R+a+0
0mJitW4YIRfsFV+kb5CD16jMqwjt5tP746gNGxbmrgBgpjGPVsuz8hACADv6U6eMbOIIR1m5we3N
UJ/CpHw+GziwpIPGHXZ3E0hU39Y1vdZONvDyAhFvEn4Wb9FLdHBY+7X+i7a8wMfohAvuRpy3O/3b
27DxxNjeRCY+UmpMgqkQJcgH9Y/JkG7kRBpcewcwj2srg8ZFXtIb1qso13+OenHpvTaP8RbiYQu7
LXTZnUOtmE5YJRa+mgUW1azs4HI26c0BhkLshrv1c7F7zNmDNwKeTjBDea+RFqTqfzTk1eVeHWdI
G5xSEO1BVxzV/+yoQkiv99ak9SiU1+I2I95nRNp4UfdAoFbJdkAuMbGobWQKf85PgJaZB0/bi/Ls
y6mmKNcyDfIWmV+foC0auqPYzy1Lca12RGBuJ1XhhVBm14scrqpBa+fudy/VdNC1sMHXW6LWmREg
TNdukv3g0e1O1LHr2VP6NzSaGoOg6BScVJUNsihJmOmt7rZt5KQr0taN70cApetN7cTRfApVKJeP
m9v6HTiYTPbgCnsdlxIEHxiGgZDyCrBWIpxUYAEH0RPnQ7T1S6NO3cXEwg03CskKf0hhd1LOczWF
8DyiEDZfwNDkXFwDGPt3d0EwtWCHfoTd4PjeN3uh0GnNvQbsZ/N+aygPYDo8oOIZSIDt0YhkcZJD
vDdPJniSdklpUMunMGFMnVIRDVrvcSC1Uk1veprWSIX0zEwTmkYFEni99AosEwM1Vw9qomsNQJQW
+iziJwXOT04l5PTU04KSiagEPzM6BOgitHwbk7e6kL0R+oEXynD4WdVdS9b0Jfgqs/tWWariiGN0
Dm4BMy7WtrIV5dVstDhgU5kCJrhwIWjG9M+4U83m6Niukq+sCVyqq8FOEync2pHj4xCI0UsT5X63
54GAiSJD9oxaFYlMi3ME0W+OmTd7Wonb5WHYdZ3CUIppbxyBbo/AUN0/e6b9XTifneSq8y6BfOe3
66SXiHD/wubkX+TP9uMoByVokpP1isOqYe4m79oPr4iNv16+rVsbK/GF25F2GnExB+6cICEit89G
KIwKvHDnym39sXDAD0IkgG3rTU67pZR3dd2QC1r4YxOtrW2kBWAuNEMaznz6rQBYepAu1oLMRjlC
jVvjoMG0ZqhLUM5d/9vZdFetLy+abgizM6WBu+avh5Z5KXJf3hxt1c27miej3q1rUb/9H1A3rO4G
6yFWjsmKASU1fvawSQwSJPhIacfq3wIpEGB7ouD8eoCGLEmn86I/kFiflBn17C4DUqYAcf6OKVvJ
RzUy2fkWDRnEuTCB4QOn9hMaHQ2HR9QQEZyWWuqVMhpkHr0CJ+Avh14pkWOJCpZFKugkAs5yIZL7
usV1ZXyQVAar+8NCzSz27znkLp/TdC4K5uoseec9vAW3PkaeDuJbPyyN+UGI9tTHL34illE6xkcL
ssQhsnOug/92zim01NckMXoFvdEONFUuo//pZ0xOvyUl56HfvK9vAzUc5Mv2LGoU9YGfuqUGvJIz
623d2axfAxB6JUAMHL7f0MWWigKHH1wgE+aj9rRmDBOL3QqvD9VhswvpmrCAcPF7rpVJlO+fZEEs
NAeKQBfmmmedNjoIu+lsUwrUyQgpRQ9mj9CwlQd6qCAL8DqhBPkhIueafYRGuhg5u1lQgDSxFZIt
ERqmw8GUa7XOJ6F6oIqgBMsLksbSaouazP/BCF41rkTrCvu+XMQ/tH1w7I6eD50XgEIr6AAXhaRu
L/gX0uXFMJl+T+l2ZR7TtRLUom0Ug3ZA3MOIyXdmC5ybOIVZcSLLlV5WICNhUw5EGdplQSAr6voo
gOyddD5KpaSkaKy94ZB8sWO93/VHy/wYmH8ysomnX7osv/eFCDXPf4dF7fwwERHfGWPf2KTbXssx
ySoKJPR1yqo/K2n83CbZQbvJeunIO5JWPPGGnQXCg95pj/r1yAY7dXA/taLIKgUbz5rC2YWnAnS9
8sNtuNYbUlBHU+D/WJNIUfJn4ik86tX3PXK+JofMMgzVX9Bzd20YLMaB7RHXbUKz/TzbreaxsjES
Ua01Q663hkAFGj2NyZ61tSdPRcwTaMHR714T/YRD+3V/gadubUExi4+MF5ZsBTYJcxt/qMYSLQDe
6AfSNYlgd5VWTuH1ZokpnNqQKYSjPkT74yMsLbfkXGVcy4CpWHJYL4tKHV//pJ1vUO386uULZtmU
C+rpSvpE6WbfBmu5vTEw+yiZEkdad2/R7bho4tzBanaJR/wbuC2d5N3XE3y7ITPJ7wMQNOyq3QYi
WrQPl5Si4B8N4GQiomgMGCbqIaaqmaIMAxGf+xdNEzf0AoB1P3ESGP6KOP0L/MadMLu/vdEQ7F7y
9F2m76nTGULuZ0LI9kpYD1M7OaGBrBAnw1XgF+aUFcJBQVb0AuA9zoOduK1MOcs1ABb3hX/TAZCU
1dIH+yHHEY7Bz/zB9umEHKqbd1vZ88yb5SPZmbIAusdshQNbVigrb8PeQiaGqOBng9LYwR7M4NLy
hz8wlTV7KsI9F8G36Zm8oNj+Wrmf50yzgMgJlaoWjPGHZUZceDMrme8AhSUWHi0T+xgIscDF21TY
WKEQ9kozgnu4S6+Cj6dZ3j4T8rXoXpl9/YGqvatPZqRrpEjzB//aMY8fNypbXtHJKknRlg4+eiV+
AvE14r8UZjyTgDzfSN0mmwLmWVMtl+CJivrvvxmPpjAYdLsyk3jynAiLPT0tcJAvp/h5FWO/Nmx3
POLc4UqxR24z0jPNOqCUF1eXmCvc4t7/wECEjJL/a34pSCClnFdG0DUXn9eoBPYT2eJyViBpbIOj
2tY0XMJU3dXBnN7KG38/AI4VfmFvSq6KEn1jyxhvehhDs3zSHF0cV/4ArO7l8hMoP8g1fAKp1BHX
fYd2j7g9Syzf1zQAWprLvGXBSXqLRn721NFAf0RWBC8o7KNgh9gmr2hzXd27h6MpZFkS7XoNbLn6
PE47cD60IJP82JRIfzIV2mLune0y8WTd4wOjANTkRagW3TOOmXBPGDA8Ka9mRP4S7MRYRuXceKOJ
/OO/Upil6ebzAkWY3D/5F1d8z/225eNq3X12nlxmtqUEsxyfOKAMJgT/Rnry0tE6dbF8zEWFEGv1
A3VBFe1guA9UM8F0UHGii9zx8g4SvTrL7ab5+vrHsH/GYoJ/Pyr0RVdA0c4jWnSDN1em53vvQJrx
sKpRqHfZ8MDmZmKGPGm7cp43A8lwPvp27BnOOZwiL13SG+8j/Ju2nmKOjxfasCPwe54m4exGuWYA
EQdan2nDpPSl3Ck9luBBJOQXozKchDrMnI/VvGqO/YRJTET7PXmZ00jH+Z6lcV+bAgaLpBtO9dn1
RrgnZYLOlZIbzy+bHw+pscpKBZ2ErthClSZSg91YP7J8tTClA779F0BVarNfaxQ/VLvg7DMfT9gs
jJZX83fv+Rg4gJ8Cw/nWCGU5N1md5ZahsOymQ1llYvhoca1w7DSZ9CP589OOU8aGh1vx7qMBkyzI
Z1PYEEbZMDytHJz2rz/3aUARV5ds1TIGToh9yhmwHWuX2jPBQjfnnpEQ+rd5JP9GtemAWS62o1hK
RkB/ZjhcYhneku4+C8pMmtzl1lFJbzuuj+iLvNAV9bWu1fSKZUv9MayNv3QJfTcVbuyZYQi7ZKzA
/eIkQ7QiK+he3OQKxvXamNva8cfS+tSfJRmTvu29lGmp22WfKYC2qEoKqaG0k9JeVP2hhxzqSJKt
pa7s9GC57tB/YqUvZivN/5kXgsmuAOgf8JpsgZGAwtJZJZoQO7OwwHPtJN0Qv21M0U3Ka1+PxKxu
OcI2ddTiQagSSsvztALsFkkgZLlEVkRExZ3h1lHNpnr5b+1L7ZVjrNwlYS9wOJ/u+e0hCJIrOUPA
iTT9xWcVpE4UHKJJHgkEc9QxIISeFBq0RN915GEspM3O0BYDS0PQAHYnKnNfq55fh5QF7/XM17Oi
xhv+yhua0LjPQcJq61h9xRdVKhR+5xgwLjr5WxEUbBJCV/CDeJ6qG77TAmQYxidbYb+PI9ETt9PO
ryqJqQWxVix/l9Ae7IzffFA5vVEX/MYOhMBUIvoc+z0ibfM5mueQcYUw0tEX4FPQjfp2nVt0paRk
vqYTVEAYW8bfpyf5ccKsWjpIK1XYA2dIkmVBEOMaaHOIZsFw1tcAXvEYzP/hzDrCxMVvE/359QRf
inydwDZBFb4t1Xp1Eee0lyHJxYafUEl8nlqqOONgIn3hc4j6rdLZlOrmEGRQw92Rd1KZVE6IQhgq
FFWzZ7fgfgBNfqbBn9n+SVSGIkoP1dDbiMJGIbSqx3Y9mSsIfpjE90usa2bq956OOMiENDDHf+hr
aS4iHvBq3ijKfdPe/7HWJKz5x6ssCVRd4HEYnU8+cMfxdT/Bf+thhHeHS0A14QDXn7YOPZfooRen
oF6sEglhT2hIdIW+baOubrVMC5Nj8olqDesSSF5KbfJsB2jOLPgwgGHtpAQL1ddMu17UFcZxdw5Z
k5FZIZB3vHTKXz7e/ZJuRP4n+jjnZFSCsX+rIVLNSFE4TuDgZmg1avQyslbad8mz+Rk87PXxitDQ
maKmY+TMGB/W662M+KpEqB9wWZf2T9cG62pRw2NJ67yk4QJhHz/plpPGuGWxfKdHKJIXt7QC0wtV
r/aWfYkAnG3thqo/j8e9+3NzA3cos7Cy6NA9MXeFu+gd5dy1j3rWj9nNv/4J8BW4gCXar8jhtiGk
CShL9SIjkwxIDfJShToQ+n6OCZMysTmnAPFtynhaL4O74fGhgLTOlnf0YFlksBO4JfJFYPgnNk8o
d1VWmlCgd9oHDoOJYoWKbpJaYVSnXKc6DbZ/+7HL8CIR0VEfNZdbTwGzVzJnrftPk0uIZRRRZK3i
m/yfs40NWm94Rldz/DQ5bGQ5KuhcfZth7sCRlcK6bSCyPjN68ffvnjgDfHya2FbNJTTc0y3joYoT
c+aJAbIIApiFB1MNM9kZacR30DslBVT+3RimKQJjCl0lRXlV+UE1HjQO0dJyPqyv6LgGRHFTn1VW
NVG5qbg/T2ItaseRLOqm8s6zhJ3YU1O98RcUbpJqItOTd//71lXDMN/6J6K9eiaBNsC77X3WbJl7
I3WTL71cUwhdWfhQuUgsYu5zVqrXx9MFRvPROqg0P+EsW+f+iyDIp/l2JiIZ37HpkpGqUV/L3UvT
2F7JxznD32mDem3EHnUUbVkhAAz48QSpbTkx7PUb/6IXNXxr5AqFqyl/cEAEU6ko3uWj6dR9dq5A
h8TXHwkbE4qp5dq6w5ARPJcgt0Cv6Y7FDqwVWDwSuK0RwTQnwTRRCmUoL/9OWlOcBwlqDzjJZfEG
Lc65hOt+G2zy1ZP9ScSNuDnlO9MitDhd724ovzhbh/mSrxUz6nHJl9uGfR4XMWifWvdQSvHMA4cG
/eUXGFl7QKDtXy5gZVZPZq7GZ3i8DZk40AWaYC4oiAVWtbbZi2XFXoF61se2P/GCS9qW9CxNCxC3
tEuT0uRv/MdMJT03km5u8dizEdWzd1WOh25D4lhPOHLfwxECygV1j+Ci8p2UjJaGoxpbaUNsr4d6
/ouaRQtnU/gCRGvqL/bbdd3BCaFBNYWtaR6qVSNe37XF58hJ8pwzYA3Zf/SzOX8ErwT0UA7MGpMZ
GLMEAqrdH56GkwbuMTm7zuu8vMfEKGByIR98htxa7O3YxXYHx5lUiInigfcdWX/6CWzz2ktWmGeg
A3f5Q90g4vSZlqcq5qzWj07URT2xfgcJNtpv7FcftGGwWfuPPkk8pfeZyk6J/CWRoYa7H9xgV0Sb
KPyEpfLlWhVsKdk6RYux++B0vSSuZoTa88ly4OpwG88da5ucjae+iU3iAKFMazgLe04veGbrCc4h
grvvyXyn77nk2H915t4uihQtyRgzjlw//M+uXsbQFSdxl8nP6xf1GMvjHX4EdQ56qfYyj4kcIyNw
apvK9vVDrCL8KwNIv0BBWtDjtngNylWitI6RcYn3/POsr7c+4GY6TzilQGkUmILH7RGeoNXAudAd
hgGdUCWZjkZ+jhjJ9gjPtXGZ6ya1aZSGr6osKtPfQVx7yVuNWADFPJ9YHRUAqJuj7iGfNVGKwXRb
iu/m+5vkAaDEEfSvDlZxKbgkAlVIMNfSyrDAfQav+I7IeRug7pwtATURamRvSwqAY8JQ21wZQ3/U
/A5GPsfhr5GtpMgC5dcfot5XuiraxfdkvhrRtFIrTS4uar2cBFoueVJt8+pqhhSqVuDGJrkq58C1
ySS4C3mmnLE3NJZbXw7mJ5ToSuBI4WO5Ouj/h16Al8h5KuA3ud7CEI7Jre9v+z6Yw9FpPrszDkA0
I/4z6lG3N2KOVzOykDE9uPu4/OQOPlPiVoBPwuBLaErugFGGxG750FiWaWi4j45rAfjNllOJsbdb
ROYOmL+4OwD4VwkTtm5pas6Jg7zPENTmvHv8pWLFGmog4CiQjkjWHOhcmljJfs3zdO+LBNk6PGoK
S+6ptmrTBz9B2kjphxh+z5Ggq+NyyFK6UKwllszOoJIxEZqjRRdnTUPxtJj/VourNo895JYQnX5L
DHAymVULCiJtvEqgAtJTkYy02tXwSnzlUD22iYSnvzvW/khTLxt+GG1CISLfNV+H97LuRQxEimea
XPUjHHYBEjJx30gPEoTpCToO8kybQt6OYMhHGuDz8D0nB8ka9TVGpNWWYmbyT+vzIBRCkYwQyIFD
taafxF3X/5lrOK2ETWx2gwWpXjZ5Utu6SjLcAE55kPhDzDG9xMXqkPv8vjXbwthkILILUqHFNQnc
jZZZLcPTKXCP01IVKRQTaixgYq3D2LSP9femsei9Dv4lhl2PkKrRWu6EWdFe5RLQUzA5hVFkeYVZ
O32203twi0LTU8arzZrUjJGof5DHT8kbyBJOBZazzHsa83lMqY4uJkci2bHzc6S0fVnyyXGcZD7t
9Uasmw5+BqiIOWF7eq69oqzDkZQFt9xGVTboJbv3zjvTQutGiOXframGH3Lab+jTSdvcB26bEdTs
+kmAmstgAqEyxiuJgy6+eKDfLO2qAqs3V1mRyZ0Sq5q0yWKH/QXRfoEEy4NCnymPSC+RSgotWFjO
MUfnCEflVZwEj4/4LZarKnjJQBVnq+Q4rSq6QBR4BtLtOsESevVJxpPHakHcSFW7oVorrDHA3Dno
uuXgBHNSLuDc/JSIwSk0Dbwj15i62HkbBfkOZQu6nRkK+3XGkozJHreZWlhIMoO7n2JWIuGxUlDV
1ZLIeLh/zqlu5QUxlkI/OWwnd7NTxLyv7KCJ0NBq82UTHR0047i7BLsGWkvHh1Xm3gsWBEPEipXp
HCuzlOJZHl4X07mAH4dzeAKTR92AyJQIYZzTUCiYm5/z9snfoMZ7yrWJ2r07az7F3h0ZrZlRJoSk
K80LdD3C6LfNYZ4JoNOuQTEWD41QOYUIivCOrI36NpvFZu0xr+17FW2xSxdmJ+f2mkVf5P0+jkbY
PjKJsvGOPrK0Kra3PDZpMPFtR1YOBZWGMNIc3bw5zm1MeKWTTTeV/Yea0VyR2WV3KhC5r1Os1F6H
VXc44EnLthFASAaL/97/TP7Xq09bFLvscAVaStmAuEalUwl2abvWJOktDAZ8aKbdEv6aRVxD92JQ
vB28hPumFdwWGD28lEosnG7/Ip3rvrpHdAVYvPFFDMEY6TM8t2vnN2x1WTf7ZNPkJ1Kd+8R9A79g
SMZbBY4IUQqgy3YR51INb3/OEU4i2l9XXjebeovrahgcdDrJkwg7u7bBlC+r3d6xtVQtFt0URtnI
vMzgwErFMOJZIYlDSoIxY+YvLCCMlm33RRFAQ2eMDYPDs+4UF5sE30XDXdjhG8obSRQUejwDHS6s
A1bQYmq5cFE36hbovlfyyDpAGtCITEse7cC7EAfy/l2zLiE7mSzcbV/SPigtVogpR2F/i2eb/R8w
ebz38gmKp0dG1DK80TAUfanG+tZoPDhc+2zRwHufMT6bHCkPkIHQmHwJ+d4SWYxXs154xV00eoTt
24hiOYZwayfJA9NzgUDXsT2y5TV0vF9KEMTglneUPXEYQq1a4mRY7LnXUqXQjb4WqEmVeutw/fTb
btpQF0GAUtjPSrE8CVSVCluB7ReCH0N+WF60Qgom1hHH3GfZ8PGwOgHa+3jMIeLqJ5TpOsCfzbua
v8Th7wMe0LXr1Yh08WoAEKIBTI1h+FJgmsti52O2lmYdabZck/XobSIlb571ayfZnp4fjBqGeQ9v
sE5R7kQmJUEf24v5oNfPKC0/Y1KmDgcUCsnkENoiiX+aO04/9qo0BQPFdCilgE4prGJpdEwhBN8T
Y+yD3Yux6eJ/yRZXzjOVlCNTIvUxf+aS8UtR+g3RFtJAjccUQxnLMTRfx0wVPuu2d+KciqN4WVus
zO9GKrSIEXssacYagCKoKjuZFnKEwiJG4h+y1ot3E6R729lPgiEreMFhGa6hYkOEI+qO6hQPaVOd
WXRPNq91KzFe1umqkv7VsSbZ2bV6YGNmkcT2IXyi+wtRQ+/JRczvYXRyD0nYjArpP9ABvH4dOz8u
qyZ+602lMcLbtmvLnFR/fEx20haMVMCGK+YeRh54JBQzFND3vLugTsRwlM8We0TgkbzUjfZMadbz
guh+rasa4FOsRRcp3OinLyAL85gvb2VtQ5EnA+SQauiLXerq5H4w3+SknOZZ/sPt31q1Whl5zTuM
ER92cL7F/HXOHKyEZhWaNsywSlG3SFqHwq5s+vb5cNiqfLSokLWvj7UhGbuI3yP9sVxGh6mIymSS
qK+sDEAHUSM2cnxOuvfEPvxqL0ZDQRdCB7k058ZIWFO65D16mt718uwLYyQ/hxzO0eNV8F3Har3M
MlVBN5mEHQZvtDXDd3E8HixYKEJcJXfrWq5NKRyOZZeW4rZLLijzkJ2810Z5cPaVM3lX//9sLu1V
08R7WTxUzvAHG3XijoGWJTZq4Z8YXSzYg0AM8ne8ZbcHKfhTRiO1+UBr8ib8sgLvMPljxStdPqXu
iMT7GdOgbkTQKeJJQNU7zAl/hMJFBzUrcCWmPQ+tU3Bx5peak/dMCrQbRlxdRbqyo/y8dpC31idD
CO6AJNZWFqxjKv/Yn2nJmq7oVh+q/AcWnC2y6qczPcPyd8yEYyi6/h9vX1almL1959GKRb1dc8F0
Kp1P2OW62x6Yzs3YbUPzlzytu9GW7hw5+LvBi3+46ofPERv52FBCtKMydr0rNNmyhAccXEVfdBgN
JfRFqunNlVqXzxNueR/iaBpjhkpIwU5V7nVyZR8tFgDotTslDrDpSPFHp2LRL202kX2A57xtx0v5
l3UpJfMGKRBLFosoynPttdQps8zsSx2ijr6jvuR5UI5Gcj64omN+KaA9mwM0LO5mfAxjk8ct759d
0carHekjrrare088YD5GZAyjx89wUyEhZn2IDfQsJGO85qMlFgGJRJrF+758mosZAgudrlsUwgF2
QAyJFoltu3U0MJJQ7gz+3/6KE2VYsmJRzRVOGGi+F1o/iStV2S72KWCqbfzAuA6xYpbb1A0yYhDm
JzwS5phCPr56+iGoXzXl/Wstwi6FVhKbIa9e8yBx5J+KPe9H+mkRCGHUBqeC3vqAIbhlIANTrYr6
iJk+l3nGVeqzG59lnAjC0f4+WYNrqK8WgjRy6nhf94Nm5+6XQEJVUJ4WIaI06ZvYZGfEazVSxwx4
dE73ERxawExuKPd3tkMaYCeunQDx4D1V97hO8zAl0WbGBKdd07EGpCGgS4FBM11EZcSi/AEDy1ZF
oo2ODXyNatEuReqAvbY6yH+ajEJEUPRbShruiRzrNW0dpn7KG8zPtwPuJgBm+dnPE+IMRivdjobY
ypPGOT4bVvmLCnY6yCxTiIY3D3zuC20BdraDkfnMPR2z8btVEH0CGjilFUGO/AuZokl9iHAjQBVa
jVCMvRboBR/c8KnXMnNCE1TszUst3zvudbsAaYo9syUsJNhJH7iDdzDroizT177b/RjLJ4ybxQOh
BjpfCGsHNprsoNelEDkBBXvfEz9X5NeFMmV5FtP7xPuOstR9nW3WHirjl5M4Upe1/RCAqQtveVY9
7njmnZW1OkJerBFWBe/OUvS9N9fnfZh8XJnLicpEvWKp2VGbW12alTXUUf2ulbtLN7n1GeN6nSYo
av7X15/EpJTcPujwVf/CCBkUxjH7KeBoc9RF1dKMiD2+MOLUNfgaaojcxED0q0S1xaPHr4joYL/d
aGe+WnBR4ThHSbmOJDCLHvInUgh3JAu++DbtgSO2EIQrxBpf+enVElErgmj4urI/9jrhwMWpKnqZ
xed0caH9XpvHt63wf+vMb0n7M+RHRWll+cUPb53Q8iuy4E/jkrp93y1yo72UAsiDGHS6/zLxY5Js
jO/m8sizbrMpr2Qcacwwf4JvaqUXoYM6+V9XkSHyDJTHgJ7f8ovreBPun2ZsiHJXwDBUY3GgQ5Yo
Bpu7VfDhu/fXk/rA3lmuI2/zQNAe2sUOo6nRQStIvbuc3dRXECBQrv/aYGHE9cENbduGCOBMxVoM
BmYm9ba/bLe36/2rRNl4rdFWGN5snXFY8rViFBlb9Us2i5almtFYgFTkDNzoQyeGA3G4mpCs/6P9
B3eJJHdOLHJEvD6DLQJT22sdwPsWRiMbOV4VFr24DjT54Ssgjz547Q6V6GijMAW2zEnb4ueJQb8F
TeDQwxlLezWxCnj9TBbI8jKoiO7QesrGkSC8XZ3oRsQa6nf5c7AZfNxkTDpI/q+UC1E07BhayrL4
qFScYQskmBfbG7xWi5dbIG7HqBVIHzDPCvsiMRYaijDoN759qvNTNNl/+BYtIPjdmQRdqm5Rqcf/
rU8i8jZrR/N5+tR5/+xcvwJF/ghey/QMBnWdPErMq9P75dzNd+6YM33362Wyq5jg/B+M0R2pMjTC
KAI1IKQesrxjHDR+aHrNdEqkeYTTzWR/nmJnELEPnWwsMC4Ig2S96cItj/aQ6ixnlk5VP4hgmEf2
CDLNltOlRVFQTYBleYPh0QDZoICDIwahqN4w0182uHuKMKTjZah4jY1n7rjzGL4MxivoP56Hji/a
k057fh/x+28eVm721fWI8mP28DhuYvsrSuA6qUc9lS+tMb6noNX8JXhAP2ir+RBtgAY/1oHsFla3
QfSrdkkTqzJIT0HMn+I5UmHtAmKaD6ySfGXr54EO0qqiyE3gmcjEG7pGNF8f2jyzt3S37pWk0uY1
0UGtYySa7p4r8ptLdx7ysp2ynU4VTjPJ41fYwnmIrh3yu7XBZkpx+iyGo/QXFCoebv48P38UeNAu
PyM3+iOgNFmhlxRvhHnf8NFLOatlAL+PbC1Ye2c2m7eh9ii5Daa1clmw1cGW/2R4AznIz2+m+Pgy
2mhx3/DiHpSGyrMWUHguBUevAHVzhJqgEBZBoe+wzabRphYg+dYP86agx3+fRBgTQFHM8CzWjflg
WmymJ/A34SO5JlCcN9AurxvunU5OaI2tSO/ggAI/JSdILTR+GMhymnTm0vgKXm1pCssrfmY9SSoj
2YsKmzACAzpKfuG6SM50xZ0y9cuO5Udz/EvMVAgunvenhvr0GhAK4VMcUW2okGBhQj7BeAuAAcSS
EH/4BZsvp4eUYysgcY8e8AYhoFEVpnplQgWEL3FNQIZFqrjhuB2kh3u7fBQPhBsfq4S8+eoTlWSb
zWQQ/AmCShNMBSQryDevyIbp7iGGU2kpu3XGuR+CFt+UzTwnlWfbNL5gQXGEKWerMlrFCrmnxszF
jK2pfXVFGAvpWtaRdTtC4quW9p9QJ25Qg7PhHbGGDn7gBiIPkmLxEgoOjmhZulBaBQ6dLib2MvHF
T/V4H5TjX8Hz2BpgGDXxF/ykRWFbya5h3HNhkinD6zILU+WYbdEdvPyT50WB/GErYipX0LzsIPui
V8Rro5P4oyHvYO2pqUfebgvsHgzZY/nJz/tJL4u3aZXhx4lpDqaMqPAHZC+MfhhoxH2IHyydyfPD
U75PEe+vVQnWEX151CjY3iL47QdvfF/XeQTKPZHCMpV46bQN5iRtW5rwxcjQtqc+RO7PLXwDC5FD
LZefE9Dv5XKKQcZrafDpjRdXBksDsS4NtyFlqEGd1ZImerKQTYvukaQMiHVWcii8pPgLZpSve2Yn
yt911xdCMiQxvf/gQG88+E8PW98VXaGAZptSLFlXqvs0JcYmI4AtdI5p8fPzdS42Yjdd2//A3I8V
NO7qvFZ6sq9g8lMqLRSXIunMXMTazAfHwwEa7K2rWFarhXMRCyrMhkAJrnxb2QvtgFnVZsFzEz10
rzxq8xv+zzKn3gdPewBJSZnuaMGIRPRnJ/SD8dCVZkDILCVyGaKe/eFYjXPckcnZfC7og9hwcbEn
IhON4Gv6+Cly0h2Ib9+S9gCi+Zx6K9kysta9008XGpHfnsTlEXpl9ON7PQUVmyzQU1ylunyA0S79
mn5g4ivp2rSXspsUoCoW7LZh4ExAv20FsqyDCCwDCFUgAjFuJz+FGihjeEvF0to6LE2IAm1PESDn
4khRSnq8TqLvRlNaBkWgxP5s1RtEVBhejSM0C7/vCWeK3G10J8c/LBrQXL8xWaZImhdofQbkNh0a
fGn0thnYxsMZdGp2TjFlnJTJMx9GixgLeulgJNVm8sIBJDttGhNR9JdYR02mZhkWT4V0Nr+ARJoB
RTaj5LAlcsaOuMlA6537iIToSymXRo+GURoZ2t2Lv9yo4ZKilTB6JSafKsGQhUp53njXI1i2ZgO+
Sq4kZvgoRwi6ywvBfzdtcJ38J9SvhtLy5TtQvLP1Rb9jhTx/8dYD7ZLdNivWhNVFvq35ZlIXeW5m
p591dsfGBs8ivu6j4g46ynCBewJAwpycGP69k5hjdtvdkaY5fgOjjbbGEO/AytXpN3jovb+cyA41
lXIRTFy/t1wnupVWZ28jUfCDyDz4cSkNwiq7it5d8kB/CnnD0k8n6kykFLuHDeke8QDvxYeOPCNl
7sk4D+qps75EhNOi+ap7td3h5AHY3HmYTqSWXXb3F4QDjiww8SkU29mfmhWebnB9qpiX1eunTADx
TvP5cJedEmitRHwxutzKd3uxZpIjKpa1Y+G3WPUmye5nZfmkFKVLd6qTnfRUVKj4apWOFHhJh6mY
T7NtfezdmQg3d3DTkpBTRWDLGnEcvQ7bTHSjKhP0dEDaL62pJmNLVrm7qqmpdrJypTBprmNUA6mn
TfKtoFf6P+SUZvmpRIDGsPEWeATUTMkxLuUcGaxJV42tzrsv9qxDWonmMsF797fITVPUlrqaVPfe
JPkFG0I+DrNyGyl0IBxNYuqe8aixXh7sfx6rMoQ7xeiWzsdlVVrtULgYGSk0pi8TNxUIO8tDs1OK
ZnanGUfuRYTW8q8g7ahVTsSzSUT5SjQeWOTuz2cBcoVYQ1BkvE8uZZS7N21vU9lxpiQ66asUPM7y
hKlapa3v/WKQzYt3jQbSMOi8yBkMU6jBPHsjGwgXCmwgMkxvD+wTNGC/DXG2tKLAPGJZR8ZW+KD4
HY65y62t/1ILmKh5SOeJopVpEwdqWQdIJe65fHZ3Lz9pcDdCZuJg87AcUNQ6nh2BxFhbdZQLiG8r
8AUa9awfzCuXimu4hRKuLiK+XZCUiYUeK6I+BcqDs35Y0ERVVKYxuiegIZGJoNrgM7jiI7VVj/1C
GaWq0q4raWkwzH2LTvJFvZG5QDOOmTBPLR0K6qoNg992mgKeW9zIYlFBJ6OSIh4kSj5ThoyLtQW0
J+4QIfE5Wdx8sPC9tiGbNus0VjaDiuAHgMzAE8BX1RrFu70MgiJ7IX8ACsIS39vdwYxA2XwtG3Xb
XQTW70XaOl57larLaoGuXCk2yzFaIhaEnMlieLIUcNgOt1SgDBnMMHNutkhf1BTUnwCxdgf6MEnZ
mT41PUNawvOwNEdpWNPQgZFYC7/gTe/s6EcfOi1udGiy1iuCrDT7BoQBpeieX8v+YRo+9kGjbnqE
N2LM5wJ9QqOJ7nZm0X41rPaU5IkiMfLABuGQogYPUog+gwpPH0jJ58OtCkUQ+W+5giQYRBs1OBOv
EYubHWGHrTD75oqmZlfrtix43UOXT5nD14Uc6WDNQBHpXHmPinialtYMiHQAbOuhU/Tyc2E8EK5j
76LCFkZXPF0vdzxr3uhU5xE9w/aQNzCv/T1dFS7pQTSjwQnObI+AD2RDz6hj1TSjPHZDgahbVdag
CKNZqVcL15/zsawIAotHHFPBehamKfuSTiUdaf6/o2wO50mNKOpHkeIWxUThquMoZ5FvOOfumOgJ
HqwHac4WkKWBFwFWgg+yQZ541Thbpi1E0somjXuyumuFa6doJsdsv+zylGl3bl3VJKAct0gdBSVJ
ZPIITD8A6ybJRyfH9GClI2tXv5qrPF1spLfyDVd64Z8NgXwgOYsmLssNU0KH1IT0V8egU2EjpfMU
aca5NMRQbJrxcxvHu7ofO/EA3kNDK8AyyLhmzGcY48UjmDxkdVxJZUJM81o8Jf9kSCCMQrbgT8u3
Ny7a+CUKDIX7DriPiFPX4GgG2wWR62xjMVJ0E8QI6Cdx621p8HA+hJXeURzJGs8urf/AOutJkUMN
vj4aqp5sXgr3pzu2kQqyQd3NMxlFJJdvqEt+3qoNjYCbm8Xe/QW1NK84p3e6GiAVuEmjGCGKIimE
yuWnpSIpIjF2dEt7tUOjsHZsZ2xL0uv35rWaKbGLqNVV3OkBqpZ0zzRBw1/5eBlihtAMrHbr1J3a
OLOpugd7n6gy9N5fPC+Fr2n/I6KSq6wCI1Z01STAkJnb1XzH4e9MSJpduQClCIR5IIkDU6G1FrND
8NoZCE5UF7cKtrBIaaVCEBqtqVKh5Tp8QZP86BT+2qfhraeB9dD8qFr9XC2GEWLmIrAZFUxweuc0
11Flxj1+7PIVt6D8+3otn8De90MfBja72es7bNgU4dTplva+7N3iQ1MUT22QVzTfYwXkVAWCq6uI
A037HQfSp136aWX9+Ddb+C0SOXJ8ITttwXlDpBEUmUDng5EEP/anUIOH7MYMLB+SzKCwjVy+xv+w
VNzNCIHoU9svIIqVuT4Id8waNxC68LwCRiszP2mCKMxZNuJmKLV2xIKjr7uK2gZgJNLIYarExdFm
L1Z/1vmQ1DjsOvZva3uCqtGPC3JLO3H6fw4IDtEOhVDwNFyrPhfbIyA1wU5bOO3MrTaB6EDlHwIy
wioNVElshRZpI002wagHlnhAfsJYlyBukgnEgYARq7Sr9Kbz5/49vTdD69T7pn5XIyikZZwJO9TC
8O8joXbw4kcGRLMw8C2/JpICKCrcpwlQ0jenPpN8Fwp4bjUpWIeaTPCCSLCATtB0kU8faP8+I9es
bzLPOJq2oZA7zdOS88Q1zXlfd2+KUbgfOjMUmesLwqrtHbUiWYjbnyvU9eY8nsnTusSmXu1Lj/ia
BsseOXbhekjPKV8E/2ewZOCuOHoHitEiQzRby8a6UXxhc4f+vVSfGSJ2QDmXqp2w8PZl12peslbi
HGucyZWDWsRxHWly6pC2+EwYwesxBgxWqSh4zKsV477LrlVVnUDPI4Qo2Uj38bKh+eKZQ0j7P9J8
N+6E4kCwOgeI63OH57FcxQQ4XYIxCWnaoI2OHKmSM5d8HD5FWIAYU/GSxhA2GNnRNSSEb9NppPQd
ncKvM8AnV/DHJSiF///aIB8PLjenZrFtBkHkE9j3x1JUbm1ph1qwh931B78V7ogHrE4u4y+SewiD
vOSo/ZW9HPosnGpixeYYmlsfgBSRZuzJaKWnzXyUfNmM3vwT0A+Peuj1Ut+6yKcthASrZmQOyN5c
pwyTXDl2wv1Ie+CiSMvh5HyySr46nIcRyExNx3C5GH2GfaROzBUeboF5c+Y8QEEERTiM8G3tmWCp
497/6HTJvQ+DFPewO+7lQksXHYxDziOupusazFuURaRFUNT5C7mzltuhNH8hIv3w2dIw3tBWCkCV
3nXeZpPOj8HteScOrku6JUf16liFcC1DOfVKpAdT3FAKqKihA4CsH9YFFONm4/KneLPLCwSEfJg0
uCTyxfElEc8982US6REkFsqvDiRypIYooss26ILVkq2PmYa9+kPhj/t92G8Aer9u9IQygbdqwqbr
KfwkZqIyW+10Uxz3NeqqptmIFj9SS309i/fohJli1TUMRKPi96nsOaxkxrTSg50zxb32omYmIpES
2mN6XdsQRAfWBDDVc0VGfcBR1Zc4gRk6Ib3QMPwLqfF+B80YthaY6mAtu/+SjtNzaPCWb49tOhTZ
vpLYHNtvP8bSakj3S6KFC4/gx+cTSYnTNSPQcqgEO4r1wY0sVeiI73r828IjJZWJoW9ERo1Y/+N/
HQtNquhXLbH9AomNx7+/LapAFQT8bVFFWhzmZ1mo+iv6SbxUBXy9O5j13t8kUcpwFFkJmbxw9hko
IROVhwA/vJeOIRwO4Bmzqz/0WllzTRSjiiMlw6naf78jUWunCElamUsMk/Sdat0CRU0wVXJicqjz
YTGHe1+np6SlsDBnPLYgmt7lIbcyC1yT1pIIeYVdW8ONktBS2X7rr/3rDgGB72/d2xsh4IqmZcru
BpVBL//kAaLjN38q8VoSSECkECbDtvQLHK46c/0dKXcMVWJWcdVmiFmJ4k6G0577L2FPvn5Ao43Z
DAh00vNrgtsd1hbndYv7GSOSB0LNmQyO5IYYERrhz3GZlmko/rgdkWQs+XvUz4uleJqEdVKKhx0o
mtwa5PFHLzq5Ub9osqEUrKLc3/+U9G6cQbZNbBwsWnaozyAuvGu5rrR/0yDWALvJavYzDkJk/HKo
7LsFq4AE+s3Yv5Dup//r/L8WqeIGY4HvPAuJpP3YKNFwhFEZTZ50CJl9puxSDBQQ8JGr/9AYZrk0
tFPczzuyiUNfGd77OMJc85YL2oX10QFHH/ve7+BkmzHIuR40SO8O6IDxnpUK6kqXQlxTWy/lnr2n
LGOBDfS2JwpeloU3Y9oIKEtqk0ucfhSrTC02lz7sdS6RlZsxVIEgJku721KMd2MwvNqK7807p5Rq
5YrX9Khw8K1aFxhZ403X0IQ9QpAFxCoxMW+P+77AhfsQJ4UKwQz/IPaRpWr3aTO55vWW4Ic+jjYc
drIlOZ8EYgIhln10xRGdEcEyhJrtCcSEzkARNjn/DZNe+o8II5Mn2Jp0xC/DvSYyj8PusOAadd7J
D/GkbS+kF6YwTIRLlGvKW3P8x/9Uwlkrg/mVQExCRQxGlpEmuZML0APJjbkTQ0FGEnhqq7Xaa6LB
R3mGX3G0fLybC2lhvF339oPjUMGjLJr7xLsgiU2X0WwqAIWhsxSIfDdyIE8hXSDmSqRNRxxN1O0c
ZqshegbngZD511OWkbM5FvTITdIiV2VP/5P6lqVG2HB1nI0Jq9l0G6EaaH8EX7ZSXXbAW/zvj67k
RgLC2WdshzgP0uT5VW47+8NF3ZSDwRWAmoB+4t7npzgMpdRQu790foaMuu9BNE2xqZVMj1LeUwBc
Dv0wNw/K5MlFTKPIoEFX6Is2annqaJ1GqhSADD8kWAYnbxKM/c5maarxCpKeu6JPs7ZBV+vDDKgK
VCCBrviA8uqnBwlhGbcUaQ2ZNw27ApokQlavYYdDgbpBb6onGDdVxEOynMrOOWwIBVswkcN5nr2A
f9xvvplTco0u2uark0X3BBMBUZBizdvjySo9ztL4/A5DqCtx5f78TmZ1RaoWWU4CUIEDAusJjA6N
V5zHcOyUDFz+HRrq6Hwnn1OpMkJaQLy0pE2MB7Ykeh5H0U7vMLkGxDyHNV/kapJYQ5/Uxykjci1v
MU4ox6rjJFieBKaRv6BaoiYvkcX11wOxhzWAPZVtkzYJ5xCpnI5MDto9TQ4ZQc4J/iMqc6qBaa5W
YjwiJImzyzLjxgK8AFyzQoAd3k33cFmYpxxllUqkFBhvTdmzqeoFIeHRCSikkwRGyx+IUwwZ7hMU
EuELv0Rtt1rs0DnMfmBZ16FzxFkAhwyqx3+bChFCMg9e0l7JJDeNnww81y7/2vAbNknN9ItxTuCX
KgF00lcnp8XZ7WXsVu1gr3+N8XAXhQYUJpeXo74HPXg9OXg/2vNO9lAiDRezu5keqg6yBuuEhkwI
jGdp2jtBB9DJ5MrZdPfYk6bq300VI6ODxsAKDVNApzd6bUFIaM+BhJWsEmfdKT5ZT/oP4Y9x3hCR
7/BT83Dreu9PuK+6fwdgb3E4yG83TSotAjcb7H+9j3qp9v8RmT37UWyXXE4q/VFgEaVuwcvjZybV
0r0CUl7O8NYew6gYSFBzgUi3EigZ7muJeScXevTTI/DgsBS76E2hUrskrs4osK+13qZJFuhZn8ve
+HW/F05u/dRCYPzOilVwc8VkYvi6fwd0qHuKcSmRcNvi6UT6MUZ5R4auYgHxGzFF7IxQCZVHyii1
qLaoSsC2jDOxRyjfHCQxuxt7BBgtM/Ej22KkLi3QC7u/Oe2nCjMBBtbMe7SFJAwe1g9691hvsOrL
ILL+kZD/YlxYVHVoNmLbK+FC24Ib0V43Hm3G2gF51oFunJsPEZgU7VGBqmdW8AckyPqnwVfrMciW
ag/vzbjfNAg80VskBpYrlY3gE1vJH0YjvEBn/UayNsVicnMeWWwnSZ+XRePx9RJlBVYopCWBgvbE
E8NjWryY0e+eWU6a9fny1XAl9ohjW98cSEvg5UDAkDLS7Mp5vADnICJyDnOBWl6PB6mqoySSojo0
22V+ZP7c76lJ+3ePgUc0Q0gua+xBMVSkcd90noBy++w7m866EhXzWfsJbawMLtlU/SKDVgiJhzNZ
rQF+wUDAefOWBE9YfuKfxAegzH1PNNgBSYjKOnbL/mfZHm3p2r8VlNpWVOMD+yTJp/GbX+LJOvka
GdAxcSjyboYj5QUsLZYSCIzIWKKlpJTPY+/d8EULdI8zzhbOgm7xay1SL5Wq+DHh7spUlkB8tF3h
IjDO/vMy3wg5OZXi/Y4qvvs/4jC1DpgcTWtHNgVz4uc6czG7rjBwzqqdmLMiHLnIVNFNdGASuU2x
h5e46TD/HgsCwo/o1rROzWQx2wX+TZ/7b+h+/L3rVJ+taU6d4tMI+nR6uQ46nDs+XzvHGSKC6IJm
QZtukbDXjPRqaEwjNiPDQY0gxoOXQ88NWK7+Rs5UpXPNuSrWiZx9AyreH0dVX0vNWqopt5wpAIvD
z6xVuFg4jLx8DB4KA+pVSo+TQPV/MSfDEA+BNf4p6UQ7kUl4i3umGDbHZqxrXIOHX6yz9K9ICKGv
VOzOQvtFpitDRu1pY8Uo7+gDhokCVVZ+Nf3d/zYtQE+7d2G0y55Y3jMxclX1+fRz2HiL6RCERfIp
hzccf0AUtZkiaD3VSocQloJ43s7oYLditVl2/oHaJt5M/XNOGT7ahcUvgC4TMPxXMrWDEpMDMq7y
KYfj3/uRXDCdcPOIHq1zQ+q6pQcEh0zho9XtmlSXas6UIqK1LrATSsiX6Ck66yUHV8BGKCpIqJEC
wimaMftGM0FbfJ6UX58xXmL73u0gSr9/0qjdsTIv/OM2kgWh/q6ruNtd2SZYRsGOfZz/R+knvacj
JUF3QLQg1pOwmrz4chNstcx9XsronhSQ9ioZHw/Dk9jpJRsJwbBGuEn2ctj3b7c7yiVKf/5pqkhR
ndi6GZ1UWjtF+PmbMbwqfMQfBE7LFtgBZtfm+yG2yPO1BNZXSJb1y6VS95nl6O7KYahWB+YEjd8c
mKhpSmjuXT8D/pUpuWIMx8sL08X3uyMsyY5uqxL/cZeFs2wIpQbaUfN5YGyGCzvdTADoy8BQa/fg
8evj1FhxCLd8K/V00dkgYxjNT7Cm/h6E9GRgg82j6+GN8rQviIwK2JHQIvKwoY2AJ5zaQ8e4n+mf
PBhW0iuovj+Zs+5B6ri6Frz2VU3MIQDElBjRwzDgDaNRtNziMbxsN9PbUe8gYTBmlWefx87bHl1o
aYi3JTrzTcucDoEZITP1h2einQ3bkuev7f3lrgkR1dn5hZowUh+eXJwI+cwc5froEgGRigdLDqgz
08zAemvy8MD+EjYO7AcBp3Uri5FGHbR2IZg3A+71fI6k2jL2/TaO/Ek4rOApq+i7C5q2uJD/AICU
EwONEl5rPXn8zX9a0vxJ0LpfGvcvy3Ct3O1zof1BuJi6nQU++7ZoMPLJkpZQjrwNcGG08iANiXg4
QSLFjaWJnFERLSwlgenW91uNt25r+PVXI8/k0FDtseKcAyAI9LovIQk2uQIyVYBy9vnFERT7gCtJ
3Ix7PZ84QBArq2JqsD63/AiAHQ+rXBKP6tJe71cMLxL9/oZidi2yu0lO/SpEIQn1FIY14cExV7Li
O2+BdDVe38aAjUsWsGEQdJ01uVsfyzRgMuRQ232BoExSfOduM0QaLoSDBXGuIQErUTuuNrNpwXOt
JVTpK7pTkODsDeNoMrSUZJptFPM0yAL0XkHeQv33X1bDNixb9CHMuUr63yMTTNxW38bcP66nos/J
ad7mTSR3tj6y0R3oroZsgaMHmlpXPNvEfDjOodgvfceccw+Gb9D5kFZI5BcIapQry21jZzv0a3bE
EvxNz8nFdhiMN0hxPM+WGglonf8kXV51q4mvm0+ZBTFm21B+T8g4bxzEYcwCJFDhKhITtEKH2ASa
PY1+yraJy9h1A+vGUTtxaVoo9HE4MpDsZcx4Q4vADI4t0krF7t8fePoFStobWkb4KNmc7KoZ5Gww
qH9w9DkR6M2B8GspABXvkEkSN1T/BcTUrCHPHIzSvZRdzDj/SEyu2ouklD9lrpvtwjSPf1sf6rsC
Vj19Zn5qRRa1HFD/pEpcNsgH4EeAQN5bHIBpv/IKRA3DQ4BE6XPDm1k720LAcYV6PfeYufZGiAdW
rVG2lrQVupDyUUUptJh4oFzdWeZwMOfcJVuJFIXDg2Sluq7l+XFpCPSIGF3RAVVtBh38/yDoRLz9
bKGL41GXUhGRcWXSyXaUDaLGNPnROVDUE7YsF8xGX96yAv989AB2RCqOhte1j51Qpg2s03EQ6OLe
6y3BebWPwNe7PgU9dl+AGA0Sgdcsv3/vdTVfLueZsM8IvEorJnY0buwESJYZ7OtCrGHKHqV5jLZe
x4tfBmcPUUvxeezUO5eAELYxMi7IqciT7vHo0KN36rpZdpAEjVeaIgJdcCbpjBe2iQpVb1/9GzgD
Q84m2mjJA2EbOkDU4KNMzV7smaT9NaHrL1esxsqtEdJOpSFYMTzTPBCtujjQOcDvegRBY3ZbH66b
XUszWUQZ32AjaTHPZbTD/pKfQh6Fo6dlTdndg4k0H0zgHyBGPKVIn15x/g8d7nIsmm6tPmHHW+yZ
KeNm1GfbdueFnFZLvsRUWGAPJGidzR0UfrkmUeKNsbnGJA8vWnTNyNzksHyAcxcilPKL2/tr6Ngd
0HslxNHL6qRm+jiopKWV+EduZJUiwI2XJyKd0Bq3oXJ6TpA0qqeOilrBQ8m2smNGbnp6bOuRW5El
C6XqVq5E8NRfumsX+6yQTZKYxU3EyWUV8HLOX4sPYpu6OQUs1ZBHE9pmPbh5fym7SSmjbXSB+GFZ
g4asjOqD/WiSs+a4+LP7QAOr2LaZU2QpyqjSSgao3N7j4jCzqGDCk5XOZUjAmBzFglS53TZRB6JD
nMniOJgK4U4D7bJ2mmIT8Zbs6AexAyu1FSaAQhO5lbAIf+j7oL4LW0yGV1LtxTZnn1/UYyX0wDej
MxdbNEwbzPvV0dAEiQwibLG29ak1snbg+zxgU1pk9UquiCIfyWCTiYZr4/jIoyVYuZ8Ai87CNsne
c+oLSAAVtfjjQa7ynuEmmLXUg/5ASCF9y4Fbr49KjaFdEslLZkbfSKj5KAUliVU8txwooYfKDeat
9B1D3qeDKwcQ/um7jKojQ9nQS73oJG2V0gvzjT13nwOA2/tO1w88+0B9I0on6forcofIYfbeKNgQ
BsHY3afgs4H36XTB76bDHVdXjzggKdwlvaHoZfsBu4P4QiTp3MNC2L1tTnBueySoO+Mf74UC95jd
yBeSRKcSrkfLETBmO3o2A5p5cFNP/uvesNDBYrzEw8fxIg0YOwwc4P/3LZ6jcHGcbLXpqWdDbw6S
QXjtdSGCHwUFyGhRJlUL+KogGLc/sR0CqCV7LFaVJHRB6Fw6NhaB7mcmjESXdQLuThd/kxolsmne
r3zJWuCpngxIMEAhUoAGHceHtVnLAtxIrVUUyS9LtZG6l8wbK+sfy+WROvu0cwbQJDYbb2PRAc+7
DT0TERBx1coz6Vn0R1vcksh6lsqFlT85iLZ6HyQgCiGpWCY2d12hGmog/4SKxPEFO/AR7+OAA3Hu
LYFn9VFjOe23x1ldgKX7tq6xerFtGNJUYqINKFPIArAQy0GMDxZ29fJOH5QwN/3+fxkvMSENTRg6
iySstD+C8xru+2PLE3Zimk3PBAJCpYp592DczYHSqCcztgrkc6vRBPLXXtp4N2Cg41Z316z8pTby
ZgetMYVT6J4Jyr5dneFPg/aLgRTGDyD4IbxfiznGStNKb55PLYQzHLxGlXXT/+du+EdXMNKRMr7I
nUVOQuFUH7d0Qu9Rs6TCQdVHTaz/eVLmSUW/dKrwIOLuAwiLj1Ws2tdYJX9Tu5nfQlKfXlpJtcLb
/h3awvqtzEfGCu45GKfDkwxuPHDoxb2xymR6kjRfjhZaKjDrv7yyFDu0vPZngKjjdmqNeE9sS5XT
0uoMDkuFHcaL/OL0nuZKij1NmAesNVYXChzZ/qGAV7tFAJ9Kj8NbZ9HVdwwGeWlYCupAROraVmEg
bDttJMdHCBlG8OQwHdrWHG63xleFK50TLunbjET8va4LP+shBcYrIWL+gVxAt+q/C3vzHia8BvJA
fVzwqVN6hJmmGpPbFiFFwhc3Cc2CeClymwXcr+aN5JUeVvr1ytFt/8wdRwA1Fq/v/fIbuLXnbIV4
7Xvg6mn7Ww2N+Q4otmAoUyy10wUxp+65qQa0SKvxC7ZW9Ks8nAPfPpzNQGh7GZnQLdJsNt6JShNJ
4nZ4VPJzXNmZRgv0Yt2iSObbuVUCkrpB0UdFwEQvsj9ZHHbjXybK8r77lUolhYYeN08RnURiDZFw
gmxbWNT2zptMrGWkIH5ylLXWYr8eRcQcOckVcf3bA6e9DFu3XyNOLmHayI7TczNo2zBWlQC23M8X
OBKn+5K7d1lnsRT3CLzeYCPRUQICvtWZ3Qsk+6nlkJ3YgTXuZv+yY9Us/gciQdNmE0yE4HxgMSOV
1Pzy43S7zM5StbH4CA59BOlrxD308YzEfaIMSbCUjl4IbYUP+lEin1/wk/7ciBFxEmTnsX51gU6K
49BKjFAEtKRsUSsK9CYrd3Rm05UxhHtAAiuCKUwlTMSA3wOhrqI8et7kmfYuB3srbptpQw+9XawC
+RqbcxJEj75RwY9JYWeYkZf4M8vd2pwkD0x0tuvOeKBElFrF7OVoMG7NjaDAeHqL0zXBSRoDIB+W
YoSwakcnYS0Ig9/aLFVqCRBYvXVSc78l8GJKAeBfNbYvM/5/iPRgq9uA1Wgq2QVB5gmHIOWIiHKz
Pl5+4qSsOPzM6zdXRDJRiaAaWhQqsr4DKVdl1c6W6KxX01KVCIaYYjd6xPuvZ2HRYbEKCocl1N9L
fG2ZUwINJXMFP/N6AfgBe3MYxTxTH+1LG0R5os5FQeuT+jbhQLkD3IYExUbHdEcyon8kBXzvFzda
BFPZMPvYHkUlY86EvLjCfKElN8qeEpxg49gt41kHyQw5yQfhl+hbDyi1vpLZwBZVoQL9uQk/37AI
TPKixpADlIkWUJIIhxdaw2uB1Nee7I9xWTI6awVT1BseMBnMSzvX5ys33QLe4fMRU/jMYlgedwkR
nVCggKZv/Qr89DZpL2nUc+PUTUFjhLX1KUhYNkRGFLdXklLofMuLF4yIof2vOoxuyX7d61RztGwd
eF+W4jEVANGEkrh62vtNQNOGE/zMQD+nHlawmM8ZP2BLm/nqH8osfeFz/VsXSIsbzw5e2Mk2eOfP
5RduTNQUOJ3wNQO/g9v1PwwW8Ya8QVXdrGZhy7b7CZ+4h5nsaFhPeGm+QWQkB8gBKp987Jtgkyv5
eAVVr6vWgWU9yHZGj1C4cgLiu6TLULvismRiY4gFnD/Ovtmfkq1zSBc5cVNc8kkisjbKiTLMeKE3
K78xJpG6ynHQyABVdR1rqAgNVpTsy/EDEMEEGdjUOcrin7nbToPyxj9hDmuVg5Ee3MESv/sIOtsu
VxxfeKsyR0nhflE1cjxkryho8vOGP6lK2NJXLf96Z/yYQnWdXATFobiPncIVdfKbEPJ+f4BCQdPj
DDW7ZuCz9mII6c30SpZo1SUFXLfYd3KkfpVp7nvJp06aW/pe80sSBv1gOuYf8TAoNNj29gHPCQmV
aVVpAq54KEQUP57qfffFsRX9lCl1SsnEt7W+rQMoZJNRLjRi15fvzsNMxkhz21SSH/eAeBJliJ1T
H7eCSzSEpvMCvY+e9R7aC2drPWCvLZFC7JREDjoCVQvoxcgPDVuPBz4aKen+1/5IzCjHBcQkLBS4
OiAIoQcXLFVC2NfHfw6ucUvS9QlexOsjMFu+/nMkPskqRgCDn2E+JsOMdDhkj5il/o1ktqdTS35o
VCoqETY0Mz7SEL9TD1X5cvFwPIOlfT7xDG3vC0KkLb//Eb3cAjOcWS6PtyA8u4RTj0fs5inpVyjN
c6RkA5WbLE1sMV1Wo2ygJVFI/uHGZVS8jPVPN3nqYs1FpKYmQZdo1ycoyc+J/9BhogwQqEGGVVDf
H2gWSpaoHz/oFZ4S3+TnepTIrOhfeQJ9kngYOuihzxZsqh3MFkZm51P6GHjhB/2XWEo53lgiLTD8
aIqtGce6lOH6m2N1pZV/o8l+BXR7MA2Omn+G8E8TXaS+J63hOoxvap0dGt6N4Qyq/DmoW8EwNgUA
34Wg9tfiv7z7G/uP4qVbiNZy++0tWZwtnFvjbiiFE7jWNSqpf8EsF2rsLRhkMnFcPOANwPnB+SbN
wWUGxt3grYUv+G1p7k0vBWzdlbn35AdGF/5kI4ilV2XuiPGGEkikAgUrFcpI75ucVf0pGbc7RoD0
sleKA0oxMJ1UPrDdumMQpHCYlWOudJpgAm+R/7tr0SpeksKkrHVxhMG4PHoB0BIIzzuk4OUgip8D
RkHPfX2HpLMUIRGY+u7o5BL4qIR5n/5F2XavuPI7FHjDMxiSXo7ijG7O2vuUskswxmNx4E/18YK0
IHbfIbSaStM8+VJQjnZE9CN6zpmFYOJ+ketDRaOmqjTWdrp7IRmfRtzAVPh30hlH1OaS5pUs1zc/
eCqNsq4APk7E1CIujGumlC183xTd2mQQQ3fh+0b29b7aY3ph0SPurBfBRjfNBS8MFhJ+1i925NeD
Vj6rpcoJD6d8nfLs5rR0EANryJm/qrUzwsuwfVSvVyXn6ojZ+SuWT3ATRwKYLpFQq3mOhhC+7x3g
YgHm166XZ2XrNfdy44Z8bSWRKJ1h0fJVklBdtI7wIVaCM1jjIRq+6WrgcwHXEojwnAIx0CpQpADP
wEStTezPzuuaw//6frMgXJn0rJKWX/3nq6CI0wb54pdfH+iSpq1WeXp+WkPBWIA+UX9jEXK5St9y
0ksk+YGAL5NvJTl9+5YQaLSsON02iqL2Osfw7X7oAbObei+NPccy4fl1VOesBD/EeEPSn3fpxTOP
FOutJmlz2xNGG2lr4ZIqZFFewL57QxoT/FsP2d37C0Kl6uOjz9mrcPBqApOEjaujS7jA+q8Nu50b
lIfNw+VkPY+61Vnt7VB5baOepjPq2fAm+nHNqNvQ2pWp3sreNj96Eoand4b+LW4kWbDEmU36FrcS
lkutYKgu0e9jfkahB4CViixfAVoQdOgGLPxAuRQzgFg82FS4c73ZoC7ZR78KRTD4k3NB1zv2WWw1
C2mPAP2xHE9x1Mcm6DWHl5/Nyx0dDku4S6pzNHu5GYcY2WrjUzHSDLuqMhrFY3CrhoXH6NWfqa2c
g9HeF4K8V0bvUvXLlJ/N6sQ7toDNJfIyuJ2yfgvwPN6m9XtSJ+qREeIkj9w5hn75btzjEULbRYvm
K2ZcbdqTwDf7Aaxle6wTfh7TpSB2at0igoC+V3dzuzlVPEW/Vg32ICSas0HP8T0dPs6oqyFnvsAz
mPekiVRQnslOyxTzOZGZ4xI5SoU4kXgWaocBpT0O+TB9qR3xpW/w+gRM7Jx/kzNT3HSe3j8hL1jU
zKxPLPaoEbWDcqkk3TZwHtMFJlVJMKfmQTa/t9Vn2ndBDykDjOA1iDV/n79KZDMrK0UF2M3keBoB
4ccRJjmCLlbXBznfiuhpSj5T8Rxl9/c5MKJncvKY1YFRdL+Sv2Cz13ddL3GEmuKOMPCCgIV5e5x2
PujgiS5FddyJ6SoImXyND13R+gPByySN/MYj8E2nwXdMLL6hqh9U5fVoJJ45BkJNpCU+kait1s8I
QsY/Uo5q0ThH2mEtZIFJM+GhopPiGyIecfMrjNfRMgvX6v90H7xDICwse5BD6AIMCT+RFr4QNP8Y
VAALw7fMqNB2mcuYtD0W7VdsFOkhQuS2mfKrf0Ikc501D88oYTRx2icGK3vBL/e9r2IjEk9hur2y
6Q0V0CBut0/XOQrdH376VqyCHUEkOSgUXV+YVP5XJccSmoCEIEbt4HpDHXaNxwvJHXs88v0TJw0N
Hg5xCHG4RA6G86MGFI0SaD3Cy/+IRThmRG8sxeVy8mgb5M5yl4PF5QaIZ7RM3j7KMZLUU+9lAQnI
uuEgrcSfqZPNbzrDLv3+0fp6nQTZ+k2CpOw1XTeqtRPShFnCcv3+BPa5zEkZCmhDjLawxfD16r/u
ZrX8feY+H2Wu5+wxXOoscsK0Wp/uIDc/FcjUk57A1IzqsnN+FNFcRhYL9hPfrC82GeToSA/v35At
rHuzmJAuSzj9cU+EjWtmmG6Hnn16PlXjg1xXfoAY0jku11CnehMmeCFFFAmO+eKs3PbC12zBlkB5
fx8aZLQ0jygdX6/qSj5W7FaDNP93jNxb7ttqA1mhi8GLcfjbefMhBhtIwGL6EhMyrtYnBIwVVb5b
KDW6Jaxpa/syds3gHd6QdLK1RtJd76QGYw940U+/NVNAd6UeH8b9RegRYuTqeIadUpR/BLfXE89G
ExXj4cRopMlbqy3iY13i8Lw09Wsu6zAFxyxLJUrT8OqEnhXalKIh9iL3VfO39aZoXtKqQ013JIyr
dF+jQ+tay+I9txGDm3pfTxXzY3EHJufdwN55mliMbtWO/u6BiQfLvLnFy4nYqrPE/fS48v1E5zgm
SG9FgcEPt1PDHLJi+f+hQ5uRzRiuYFVf4kbIoPAdPoseqDofIKPoyVN8g+mYi5EZXINBDt3orTML
T/qia2U5deaONQ/xW352kcKO82dFYGmSofDjU6SSq12L5b8kZsnNDVXqr886kkFiCodXASCdUjRW
/4fQMDCjcOlO8xAdZ+wvpKc9Qb1DDFiYbXj6Ri0lGdyAVopzY9CmX58uU3DupHmMviyrhwbTHT4o
eDD9octs6BHo/u+LYkMixH8QQBNPsHXLueLiGtcXzetFirsWMXrXbywyfJjj/0/BI9ylPWrwZ+WB
lnCBL5+Xl7P7ZmenDw9spuhquqqiDG2i+LoMdxF8AW1yhGAbktTYdzjhQU07nF4s4L83sfVR0FI/
Noq0RL2VeSR+rmFfJFUJ5tpXbqoOlXU+GdouvHTFAGtX11mPE4r0TId9KJMCPWeEm1cGNCOhOi4C
s++pdGy7gk4xpzKRHsggtvoaW7Fh69Kk8mEVYVo0T33j1w9J7Adns0uqTVt6XQlQY7zA5Hons0G4
WlGEShz6juKUzZRreUPqpgBK8tgezccaOGOgHJSdJdcBlvg8m97yPuXlij4kYovLChUBkxy0O/Az
dm/Cz/+mMF3PCoeH7YQsVCzlAioCIWsDKqP1iu3QTsq2nCSAfrzRasEU7/EmVPfqZiYB9OZYjTFM
cz7DEejbRFeP6g96z9GADJqgz42/Iictwc/jGPE7J4eA303Ny9k0FxNh3TJ+KnIIlFKg0+AfsPDn
stX1U8K9cZZiCVrIyVFMtElaoOR3HY1UebfiUW014Y97ZrUZ9ySj4tHKZlhektCcd6MO5VQuETBL
oSuyV9IRuUekoJ9+5ZAmCLzyDqOnJjEzPVjTwlNnOaPk5wh51xFAVgtW1nuwrfWM5/w7q4z9+dSu
RRWn1RRXE68xXAycz7BxohKyehrSjjZAZLgQjDp+t9s5rtSHuba4PyEVX7iFvDc7sdWOhETUiYIV
zoNmiA53cNdzJB1R9JxBQyNMrjym/1TobypbM1q7q+yWSn5UKcf7PoYcIVJ7Cx4ZE/rNlsRGZfEE
QE8G9RRJcTMYCsu328nzuCD51bvp5KmnwJPy+branf4kAehYzCS/CGVfFHHkrM9hWjEnSiobSzoO
48L5b3kTEXwAPK6nMN3PPin4mjRtUUtAo+V05x5v62abagSEP8jirzdukq2hVh1FFtbmau6T6cBP
+cOROC125g78svAfV59lRu+uTiad5ELgR9pSRqtmsytyBEGt5l+60fXXyjmcRNI24qETDCB0P4eB
8/OgPbdSzGlzzffRhPVV7XBxQivyEuPFsXsRYHtCs+OT53V2+/s2KtoSV/WCSuDeGjyyiCw4LDUO
+2JrixbIV1YUHISCknfg4kurQAeMzwJScMPHCe95Te8GLMHv6jiwGPeCd2pHJO1L8H/sdCyiOews
zNZTUdpcHUGOoSY/7+hPtPb/q0/ier87mzkws8beHGbIOB0O+1S1wIW/VvH96AqVYq9QajwScj0u
blPpSDHRruT37ZWFQpGJFvxeo7kH4Y8lTHYd/qLAyHJw2UwHq3t2k4V0RfxfSddPspHMDAiwLZ17
7QSxar+/9kF1rBgwlSZHoNpGB/0Wsi//8q3Ay4Cw3LPDvsnUhVFr9j+A1paQZQcNUQAeiP5zzScN
dpSwBVRb3Gv0Ps/p+M675tM34C3k/R6sdBZTcYK/HZcBlS2YdxuRv4+PHBbV7DILjMkiXXDZetyY
D5o9p2yYU1gQyM7LyQ8D7/ElZDiOd6lyOmUsnl6KW/WGGZvJlG2Mm4YOTeu5f2sknytKXGa3IkOX
vAtgZOf0eNkoMEjmxFNn0fa9iP9ahwwcpUe4h+vtJi9WswpAS2C3ctr0bPKj5uteEF/Tb+k1/F84
iOofjuyPW/gz3wDGXngdHEdVo/7d07E1OFqXu2Cw+WE//ET/2l2E9eBDs9ejNiAurmTicuQq0ld8
Dv7p85Wrfkk1vDKs6LN8+ptbmtOdZcfvS7obMi8SkPIUjI6+Hc1F1sc4lWK5rNeYQhaoyuvbRqx4
q5avWekj3Ywj+Gz5J3JN7CZ6a/JdkLQFroue+FrOD36lOQ49RfNR1y9fSmadlTqFotv/rXB5vtsF
t0tMR8RMTT2iisFxZGIITIkQ9lIwO0fUDVDwjrpL++UyLqUlRyqrunHg8Acak8ZssO9Gh3Kbd0/s
oGlhZER8jsgbmeI+WaH8XmgEX9L6UpaTVw6Nrgt9FWzgYpEYxmcoaw2Ue10tOhoeFw4a5NQr6ILY
7dRQtQJ24fFlLchkSPXg/aBREnisD2wIwGU6Nhh+MQHmMsSllQ1ebT/fJ3TQSUq0THz+9/Snc7Py
UfwKJ27Y/v76B6YI6t6LhnjgVx8QlRV0JAeOwpQ/8C6aShHvmqJh3854cwQ+wfyZbg0yLsZbjmze
9n+HbME3RIewc6LsaupA2XA0JvbMoSt4mqbQRoaMASWcdhck41oEApKcXtrzBNyrJyyJ39hU7Y2i
CsTp8XW6+P3HWABjk5lUhuIQt+1eDCjltPeRWIDdaP3QnMjRQOjsCQouMPjq2n7daAp02sWBNbgW
k6IPdFx8n6ZT8zqmhm3xrpc+PFjQ51JvCwVB+bXDzb+yERrjasNigYobeMNKNlUSWghRawhzsr7Y
nkpROcHxEzHoZXO32CU/6dtUgmCuK704vDvWsauRC2PZT+mfCvKFbgORRwGvUhjMMpQibQuIP6G3
WGecKiL3DLILNFty089FmjpCLO38mXXlLuFjCcfSE4XkXSV8Nps5/bON5RMTfCo6rLdlb8wmDAc5
QHTKZzIg0n1Ysi553DidBKWJLCgefI2yxmfOOLNqt1E5eVOjTDhianB9etPVngTf+QcALRay4MHN
vzfNBcjn1smA35MeANR1WEDL5wDjlosOh+rTaa2n1se3KNwXbs3MdqzQBFEDVTVZZTFOkC3ZKUze
jzf64mafJgDKqGn69ClAfFSYP/Uq1jYliK8ZTa9QXqST6Ofxq1mOmI9xMozdc3ZZ36k3ypjmx6vU
D2X7eGG8hU3KlF7bqJt1zj9PJ5gaZlgIzQ8P87eGB0/MKRsFsSG9/kWs555j8nHXTFSAjy7OyIac
LFn3V7YrjpB/HDirC/LhVtKrFdpvMdH+dlnZO6CtMfyznPkjxbDqoaKP/x4l2REuwj+j4KPln5x8
tIwHfKZduJdtdSIKrZJaZGHaiChbWZqta+P6U8DwfpIWWYw0KK7nOTpvupGkIw2QOOSYLrXX6HSz
LpccZrElJTuBNcxy9ZQ/gOgtP8uEKWweVnEbzCkh6D+zh9JRlq9q+4Kru76FogYvFajXN77Egnfp
BTvnprHZePOASil0IhkreJrpgsCztVfu0MvSgvMlQDwIHnga8U/XHJJW/OSoLGtj6qfrxNFbN5OD
O384EYCNjHp5qgsV6H7OXrMMtA0wICSJXzVqoHs/QjX8CV+r0L/V0g/kj3KjHh+6aCPghHZUYSgX
sCKwHVZbsQAHBlSGpN3rGvLKhho8FbKrPsD69oq061udGFAZQa5DEqmg10zv4ol3NNVK3y8a0FnI
l3tQv0MeIQ52xAvaXXPh75oFjXTjBIirZhHWTHuNGj2IOTQ9zHjV6QeJcUFfaMG8vvsiRZW/pVIS
8YJOftRnd4oDbbYcz9jtz78kqWNsdSSOZWoUh6+kahlvH9iUavvNwdoNyUM4zvfKfFKjFPJh0ypb
zFOQHfwxY8gQexf+iJ4bcMljNhjKEJok6H1TYcUu2x41dP4FmdSgvH5grTLKRxVSaD2brUS5vR7X
1YGJ/rhgEjUfE6VId55Vl0XWcVhXJB0DCP63exgL6iJh5bIpDmIFbURqPEBKrTv81zLhVXLMyYmX
0mh17/bygDqIYjVVMK2oAzojwV8NnJiAqVXI0CghilGwxiRgVgQPPwA0ruyEjS4GlpOnkcACQIob
qJbOmFjxd5881VJFVyeEb57S5TLpe8Grt7F6PUyd/7oWAv7yqmYUXVJ5HxU/uJ5ttJj2S0NN6ADv
eUmy+uu2432YpnAMMkzbxmjMLprF8RD+08THgURjkrWlX3pCaX7wplez/+bH3xKi8mG5t6TvL7jf
CfiFYL6yUPNNPAVnoL0h0BG6MeQR1fiiqGLkiea0TW7Sx9R82EA3CvdAJYT3fNjArDIbobkWM0rU
SKGCDXZjU+rwdF6ozhppMeb8n4CWw/BI1uOxGL3v1jtDgLF8ES8focFi8ovppVURlvoVePCrrwWL
LequOlgLMIYEknNkPm37NZxgJjKX0WFoacXENRmkXI/VtL8ita91XMW9YVoZnjSvfTW6QaJG7FQF
kdKfDKYTyFKocb5n5rxUocF8WCb5u25kmRtLwNc5SGS/BXJRVy5soTAU6LS/QPaw24BxXEmb5I9N
T6RJiXG9A7H1bOpzEBE+NPbDBCCe8VPc5JXjwjnVfaRtvBV6cHsdgPrk6LkMqoCczMooeiB1N+NE
Ug5nRQBQGk1FUZREvJaJdy1uRMxbdpVK3Fe1IQE4b+k8IvS/xMSsrJUMAy1s8eTdwVDwzZv5R6/T
mDjkC519lGCYnWSr0u5ifjjw7eM2eyivzdZSdeQABCNgMYGoSLlQDCXYN06w2DvLnsvfhn+vV+Td
Z5ima4IoD8wdpdTmk91vp2oUVym9U2AiwRrXkdKjBYNE2EHAnPpzvxAgCXBHPk5trvnhacGfQC8E
c/qqfYBACrJ1WmMVkcJoM2a/aXITug7CdwHTMmIqxXxKrlpIxAH8TdwDex0mJm51ud/DPrLxPYdS
z74K1Efi9JYlKmBYLopg1ujaHUvyZlH/ocL5e+olPaQP62kAnwDDuf+NV3g5lntNCRfz2tc6DkpF
bnnonx/qaSKJ4XIgdB528FFyAycUN39YmKxfmEj98FdN8Wf7Z2CIw5At1TmzgSzaMyIV3htrIojC
9p3xQt6vM0bX3IEO9uyVpftqyJ449fjGUUws8nTFgw/qPwF2rGF9AisEIBFhvjFk0B0b7OmZtbL5
+d5WPS3+d4emMDzjCfb+7hO0wuYz5CqWMzoXDVLphayEaZPQ8oXeVW6fH/gq7vvcurk+h4t7mGTE
IgR7D/F7eQ+JxzyqPJQ9Ac4ok5q2TyFefop+F2AL1Wqd5o5msBIIizBI4OYLe/eLPfUWawfeFFKo
o2mw2WJpwCEowy0KQbQvM5u7V8FKQQcj+JGi9v08RCl/xXPCEeJP+/TZs4tqYQrq0MjercpFRmRQ
/QO2LGVyzaDB36NYFZvJVgca5UdGv1JwfD7QYr9ASyAwg1RFjTEp6iG2LLzA7gsvXP/z5pXFfFZU
F7v+UvAEiJFTTzsMnip9wyW0ELyNwU4+L/PME4bY+QaKbwRymRi2GAIM29zPI7wbLNbnEekCVGDU
sY5NZ6GkF6jYBKXmhIH/eJ1JurkepuSUbMcTHaogGl5sG8aFi2iRH7uNVHo2KcXluszB0WYUnfpN
O00EvHJyvMQKY+rYEFDmg3fIxYJ5dH/w7PwTvWbCsaQVgfZw/3QaZrTndJVQ6C36/w3T9TjzaVaA
po6w0HnHWGaBOeU0RPXuMECPGg1U1m4RgHSuPqk8N4AF+xLow/XWAJDzWLgCJOPIH5YmEMDvg39Y
D7Cqr084SDL6GayPY+c/3xJmz2r6gxI5KW3DWPb13trboAJPUJnLl5NTm94ytQOULYrfoKG+rUM8
DmxM/lDwqUq9Z80TX2wZHR00nwb/brbSai6IsbbfWKj/pYF4WnfOpo7wxEXjsgrnjI+esOoEHhfn
HyhCaGtHvNFiUQW3Tlz0YNAHUvCPvcyahqQfGuK4aI8a2kwM/ddBc7NMcPCDkv5V09oM4zTViJOc
5oNb+2t7THkvkkNS4hkOiey+uDPBjLY9iX5zPDFPpnexSyVBevkMu8Ty77LVSjAog2SgV9+sXJNG
q4OR1+ImLS6FfrbMCuA4V0u+gSONbD81ayDxE8AkiQFybeYTNPvmgNdBRBVo2hiUc8d5z+NiBVwG
RY/umaTvL5AlhcNg8N/LhMdRtqQ8TE49Hl/wNMAAQnT6u5OkOS6Mic9wlEdgAzfF6O1ZEgX2Ue4m
0/VuffKSLjJTg0UFbacxBH59x0bTpZG6onS3lSiqtnTfJHWYoG4++kxAaZvymru+dMtP4QJ3memH
oEW1P54eITfrMWVFdyY1PFIOHHX9ojNTyc2KgaBUb8fFBxPOFgx4WUqkv05pEPv+uaSzd9ngQzi4
k2JppkGjeKWpiAorjdCvHBCB+lmuerFlE/9mpnW3fPa8UJMscYrzTn7lixlnvuCcCPEqZo2EoUeM
NCDgFD/fxcuWVnBNS+AWtIWaAu0WvhQ87szh/tkaF1b/m1LHX1/rVnKCGbsZ/RiEUHvrN9ewzsBZ
eaGUZa1mYwkDZj8gl+g8/h1uWrvfh46L2svAc6Sd+Opb1NKgoGXfnv8cJcA27PQtKZcMhQ00ldLp
uVPS8bmvyUCvS9U0oCadZ2z2/ZYbYO6j+aVh+ghOXzu9T4tegjpCk2Pdhy11L5OVAPrOyvvcs7dS
reoPUMs5O+WoAQcGEfWtOzqaxl0XwNpopuGMfKtZaHf0DoUqqkFBHRNKmYotSskYug+hgyybLYGC
6MFRJBB9dh0kGCasFMhTNpv5eLSfaKeGonluwt7YXwMTXkybzcgJssOeDt+Wkj3xZorVwuKp8C9S
c4TVt5DhUezoAuqlGw8L8NpzzHcGIw2bkIGEvfDT5c50Shj9lP0SR4h2AV52WEdZRYeHNTA5uI15
9kiDkFCWI7IhIyYjRw2rpiV0v9OLDN7qgGdNJw5hwY/KF3IDD7AzpT1SO7fBkNVnnq5Ci24EaUxo
zetzG5BbFi3IfE2c4BSoIgIS24e9Lr6FK6yuG+jaTslORnY+lC03xzhBjKMJorDaRlOAJNd4b+ea
3015hXiG3Xmb2weNjTayDX9KcVFzasNy/da66f6L8LE1z9v+iatlRvebp9WjCUcxvkVyea0xmJTx
8PMlrAlNA0gb4gIIgC6oSIGjK0yg0/FW63Dsj5NRos5+IGGUh4Iwx69Qgppe4z7ai5s3QTe0bjgY
b0R+ymxQejT1Ufy5DttuCfIskfUHefxcYTfAy5xIsAm2PsVgClBZKdET37N83ACYMHim3x5TT9lb
tD8iUaxzk5f9lEFd+cDdp8WnTqvxQEn45t7fdPVemW2rDlk5rwNBlqQL5reGElem8VLa0wHP+p1y
y3i4xv64sBBNY+LNkQ2rS8HVgJHWRwBezRcG9xddU4mRCN0CByxtAfQWHznlE0kUFhfsamhse637
8OFDNH+WAJhIFfGeaILwyFdqpAh6MXw07sdwoLsiO0lppidUgzgg81+H6IirdBBJbtLwJClXj1i4
VEX26wWseorW3p/1/+k1Mz+czOEoXN8SK99WtpVhgaawR+gypodFCsHu+oB83OpwcGYSriHfY2yj
sRMu2QL+hqt+peelf0hD4C9gKoIp8UnRgKW4ERQA85w6X5uxRfrwo3v//0535FeeAZJWfb8QWQQA
Qek0kY5ORFLqO2ftSCURoa+35audCCVSlnHe8tWFDPOx+K4aZ60sOek3kibvvkXHWjwNtkOu1IUz
CxipJ/ozr89rW01yzn29YwO/RRTtbcioReuBgFgD7QGJKGBhsvni67HupgLs3q/PKdnGw14CWWeC
C1GiL+j+7qx+CjcOmGK9kWcLrKLRY8IdsloJmQaRHSUB2CSu4fjVxRFO2+YxVoi/1Z0Df4OlTuNl
WUkeXvJpB7yowtbyFZ6nvdQ0FcqFktw/XltihDMGoiZM6E5g0T88f7qToOTG9eymkLfik3cYFz4j
dSEqr1+NunS+1yjXXmOmTDSAq0OGUiDAIf6s7RHCnR3PzwQXq2+LmCcXPFMhV3RoXpXcDXEaxJD/
BinEhb+zIr1pfsoKRi7noBk5S4ydyqhBdvP3rwZzcv+ltsB/R3bX6hrXfyrB7WmhsOT92xr53frg
72VIGNVWb5b9sVhPGwhcBRjcZ9rT3ZrZxHgCX/u+AWv+CbBVe0oSd1Hw8Y6Cc7uWDF0nWzQq7LA3
CZRBVC8Hzv92sp3bZY02a5tLGBqIKUkWMUuTa2KQycNqb3yQYzDVp9D9qP6jg1cAjDrGZL2fjmoy
WKiM8SQfONtdXqnyvNGp5qDjqcEPRj2JmDJPELEBPlPtbGbLEH8z4BWQlEEDuz/ZNPZd5GoyP33+
a/bOhLuEbNtAsjf52oY0KaOsUnfIzScvGNLXuZzAEzlA5gk16dI1hIvU2tW4i+nZZ/YcxJI35MNZ
dNiHRgxkBQ2Br7N7V80lmjXbeGyZ+3rqpNZGhpqpFoM1Z5IgymJGvzuRYy4pFldh5xSrSHA7+diu
UDwsTbINXGpbr39EwxUEtAw7nOiMdKVtS703IGvTNseGO0PdIliV+l3M/A9AsgQgQOb7vXM/lijI
hbl5dAeFWmuJEa/WbQlTouajMcjQ5KFUBffl+tc2JM6w95E4Ay6riUrJs6xlLbvoouTcFcRXsHAj
we8yZfjZP3JoUQFstYIJfM8OOQZrLMmxiQ3iXR4Ak5NjNNsfiyHzDycf0HC+08COD8c9xy1tJu45
KXVism+bQD/81Ux2ElJAt+slS2Y+47id2EGT79HvKds1rSK8Zdop3kRNOH1WVYc9ESOLyn70OPjZ
eM5XStB2SX7gFA1xpP9UsyhiyhzWqpd2BQxvTYvFW7mOx/IYrcgeHflwAKsmj92FaEOfl6tr9Rfh
vL6BrYiip1fZmjFbEmiobGa1FYMQcYEWT023Qjrpby3pJ7MXEfj1KmuCfKteqNOTMOfGuktPK/gm
iTzmfHZ5Ko05P99mIShlndvdYD9REc4zsi8J0jP5F+ltbPg1nDFwhLNbHCGgzkKODwJBRYmhwjsO
b1cKU55y2IPni1uPjZdRCNzMpZPJx3udN1gUs+WUrKorAL1V+t48f81Rsjbvfek3cATQk1DCk4Ee
c46JAepCpMr8MFBchi7bAduMFwlA8uojL1xB2Oi6biU0F02q6WwgWdUIqzD5PtT1NW2/7eEO5WtR
LcWYEflGBKlxo7FHssrgk9FKIjBkaLI8r3YulJW6I0wg2ZmZ/fWjCYcRldRdkCOad1zxV8Qtwv7+
nGVcWSLqx4dhrQnruGJmuBO3EIGVQov6Qljr9B2FmOVOErQSAtE86YuS5dFAJQXH5JEVoXVOOaxe
1FrUK7UxgqMgDXRTGFGPoZoCQsnYomOmqMeSOZRFubUNKN1JVtoCme+skybfnZVZ2tJH3/aHa4Sp
sN0o2UDvEtZevLLNCZWaQlTnZ2aJPqPFJZkl0K0jt9K4tXYoytbQOLMI02zx6r8+K60DvIbCRVCS
9Lxq8I+jEwoMmA1Je+E9sodYM7O+iVDpWIAAWYmJBpy+gS8rpVUDHX0wEbI53dQvzyOtr1IJol+u
oPoZgL14swnEATp9JZfNgltRKpEgzxbN5RZ2hcXrYdXbB7Pmt9pqqSebGUqLOd0jXw2+5Xtsf1Kf
kMB2oWDdpklJo9CTeVJqrlEF/GTHlugspS/ggSWrsLZ0TlSwTtjtnV0nc1TJKbGQVu4Mqxbaep2u
aRvwOFBlugPeY0DyY6bmlQ8YM6EO3PSqJiW5VpNQZW+CONwj9jZdHEjjhShOvtT8wJF8WXS9OBH4
HJWvfJlmCqjL6mHc8Xz/WAVtE/hZn2i22mFXdcSYBfy7hYITRn3gp8w8mhxrdvKSyKaS0+jch/KN
xWySiszDKr0CmlOiN9j0LKVG1TbelBo6UzrZiqhNChczb4X271gU27FTaNvmiAv/8Q4HfRVOSzD/
yDej25IzSYYpop2prKXdI5Awub/KbMgKLW+vcRABLk1t0uNOGsLR0EtXTUrn/f+NiYnjZnCeUZ3c
jQ+fhMwqv7X6bhoQ4giDZ2vxynqAwMRO98A7heZTYsrufZjYN0MeYeFRShZS2BNxFoRUpyDvGo5s
5nsSUe4Unqi3N4nptbYOatBOwF12+roT550Y0zOXx6o1KLhu4D7C83+Mh06EWX5nTI3rRAeox7WL
uSzWa5H5uU6zJUrnoczYAghUtGpRgGmQEOatSUqhOOIclTTf4+za7Cf7dkf9yJ2xyX6LWnFEpie0
P5L86bN9kF5gIHJGjQxEFRnOukYUFOS3ObyINgq2LnkfAtMnizVCnSmozp9XgxtNid81ouTH1q36
lXGXzq6JrE0clsEG967g8vO2xtaD7VjOTjrktD8q2e4ei5Tflqt6yz47bhMGnzfgEh1U12nFkDLO
n5f9NJFdjt2tUKMlyGxZnHg03EebUTrl9Jg1c1VNEb1x6BdfQkbUqDrq+Z5g6ivr4ZL8AZGTz87u
xqayOHcDT/bN6HO83Wxun58Q2ntsqfxXXeX02shlgDSTTFFVcEjeYwD2L57t4KEzEvuQpyYTLn98
ApKb469HuLByy2dTTWJ0bpxmK8KiRUOQ+j14QWQuIOV/ujeD6bkbTbVgY61GvuC+0QoQ6hX7l8AM
dp3+XGdnsoy1ccd3jMDb8VYNR47FQcLbzGnW65Qk4SdgmE57GW3s178M7YqFyR+5+Gu66BiOvvLr
GH33dxhJbibd+xgQynRQywMW+mIhzdRWEOq5p5IecKTd1kjcK6eAckbuQ/4QOcq5CIKnXmrwuKw2
6TD3iiGQyuLUbzp7AKkxqlntkOqsDIdVscEsRBkIM0JsdbRY4jian/cmzM/9zo9kOZu/TwdL6KL9
TfU2fvAyHeZ1nmoqVISGnl7j6s6q7YWVdC0MxaRkrHSNcGKYVmpiI4OmtJHZgtmTg8HIzXb6uenp
w6Ts2uZnj6Xk1TWtUI05rf8CTqCnykkujDO89QuhhTBwl2zFmN1KOQrYp7SmaZlZjBuvRBZ/NGX3
75xn7yeCF48NTmiUy3/XCeeBXe0AwghKG8qZdsSYipFSL0wBu2yg16nf+tFjlBD+Lh6RwXQo83hV
VZDxAAMjkylzwuEyxTKXD35T8G7ZShNGu5jmYuKnyolTAPLar1ZUD+OFfQCJvbsACdNh0WBOfNqP
t8OwGjHMmTUI8I/PjPXD0RTJQqLCvUwmRYrqK8HzCI8yHpVLOwUMH7x359L2ERgl2wgjeJUOdaE2
nMA6aq8CMPVt4urJfP0xBuw6p1A9om1A7zuVqkkpvA8ZoeP0b2gG2xahtpc1t6ivCyX+7GuAghRd
Z3Br1pMIEoVpwYQMQ4bj+RVVxglP1uHGT1g15Q0OD4Hw6z7TNgRXgLqTn2N4eJisW+jADxZMYWyk
MKWwlNm2m57LwAXTCTLq9tCvzuwyO5CuQ305LMp1SOibUOf/v7HAt4WnHE4m378dbcLUrzzGov/8
GP7lqTWpTP1q4JAzcz1CbEscFjLjd/cleT1nI/4M2dqy5RV4nyJAlpuFS5o8uB60V4Gamlv78HbI
ZDqDd+OP3GOn5ZymfJ4EQwDuWmIJChVVn7+Nfaq+tzZduibDbFRdNlQJ8BS/n8PZwLfPHXmP6v+G
MIFmMOI0He/l4rYXxbBthazf83gUMG513/OnYZOo83I4VHS2+zQTN3hGMhzAK3mN111HOmkny+dT
PyawFgNWuy3Bhf/IQDpg9V2VYyRVjjR0XOvPkAyjHQ7sVq95ofBLC4G4hXdoAVz8pXXRWTh5raOO
kRycrUVDqlIxomIdyBwDJqAP/tWuyh/M75zlMlfh99PSCChZQG3L+tSuaXHtkgdEoKUxe8RLxdfw
dM1e5PgVtR83CzhmGmnGH2K/1Eiqie0FyirkLjMPJ0HFyWxc+O65p7UaMhyFMwwDb5JtIo49N8Ic
X60APrSuWcoAEUbkhE6MZEDURKpIvGEpRAXRJi0zq65zZR8z/lSXmJeTZxizFOJTTTHMlCTgX6yN
MddZMxCd92a5uZdbu81VPJmLKEtw7OyBG7Nl8a+U1YWk1qdKwq8xC/LBywfaI/DFM4aXpeBlOZZi
1yjuAbPsjsejssBPUdz0CR7r/MbSelz4QB1wCNNrQXcuJEA6tHNwMCzSp9vuL05gj60KmR4bzBXp
Ok+S4823aO04U7X3J7u039fyNjrw1DGKeGGjOspWVnRejIjfMEcAIiq/0X3N6J8jc3AHKXjAZVma
i1jERlsDl7AGo6QY4SCElYIPVUg2MJcBngrzQT7pi5YcYzsBPZHdd7aFcgEr7kxfhjU8xExCzSbt
VJOsIbsk0jdByNhZi0xqxaNTvqev8K4ixcjZ8NNQtsPoYggyJk85mxG0wvtKCeFu0VenmqCXoXnv
KUKyhu2fHt5UTEhFqCn3L83iSuTC8BJS9mWGB2Cot6pnfG6DaXh530hWlyruK6fz1lugGxz1svE7
okUbaJ2TPuliSsqUXUnDl9JKUON54hPk3T0mkUEDOKWpGVUI3ou6/4xC76/oJkQdYYkq8Z/k55Xi
uERudlaKJC45hBDaFC7QpAFnRzVEp7AV/MEYPiJSBAJZbmoF+kvY4XyZ/LxA06OM/o800hbGErmG
3ddKMOqABAa8gizcF6YadPu3uqsA5ex2O1cPrFA52bugrww6l296/UvB/T/P8574WXHEm5aWdImM
KKOCzccQ7zMebx56F7OCszMAvU/3sxgJZIg2gpw0pMU7OF1mftx3VNzdy5iARfu6WZRCTOXt/e1Y
qlepVWBJmaR6wNo9274jPYItNdSEA8LA9WS5NuKij0pIqpOP+ZVt31YcABeC19nuB6lSS+36Ll4t
Y5FAc/yyxWzsSSqc3pQaNf2677Yy1QXxJYpB5gIAAMYroX0r+rx6yA5MMNcPgYRj7K8HedNwlm+k
7ukk23W8qAm6mwTjvY3m3VcAKCuEcsJeHP/kVWKdivsVPG8jP2v6w8lgPycWvef3GIJFivHgtS6f
hz/aEXIhi4AYaUfJNAHyHAOZKr5XtMgMyZtLaR6h7GaH42eO3VLWcQ+7n2OKP5FhYSVQciiwy5nt
0Oc0lqf23a6k1sCF4pOJ5bAVg4v8ryYQoIVMufdkK1i7wn5IV9L1P/e2Y47V7QGc6cuIoVXNmc8r
Zo5HXCuJL4o4e+Itt4PacK+Ht+Qbibia7Ui40qvokeWuReRnZBE6/3zgeMQ5Suxq/LcJNNxxC0k5
jdWzldBLFLD1iblYDYDQWmfpfpfFffNo4ljQy6QjAMBbl7N1oPmdPDUYy0QGChQQN2y6URFO+ZL9
Nj8ex2wI/FA2dXM5J6a8MBH1zntlZRdZlmpfG4g8eX0k5k8b5e52rkEcxCwjeXtGA/OTUDN6+OPl
8HbSuHYO1jetC0NSJ62v2JurFoV5upgd6HUD4Xdc8P2UNL8h2GDG5c9uOFLTHcw76n7qZC/zwN2D
JGFHkkHoJCojOIu+B8SaDynrfioUp8cqKL59UXR8xROtlFd2zfYExHj/YjEBau+/yJhpZjrjKp+G
Xeby/XzmioWGDO+WxvBo0LZVJ2X6lqAj6j/6POl8Gf7gM6bAIfC2dHCy5ovp2Jb5TIDakkl9/vse
dzgMC7OUbh3+H2FA5AiIT2IjYd9g9NDFJihnm3ZZPT0kqfCsJFxEhSr1aXL+pXwJ0m6GawRzyEb6
dgyBDBXkIuid3fHLB6SFqW/QckAqzxzF8Vn20VfuQO/B0mWD9TEpZtp8wJUZEbnrrFwcY/pzk7Ra
pTwjNVo10l2v88XSieL+m7h9ahIKadlBfpBh+hWIRCuxdyki/hmMl7uCTzi+6onDCp1JwPN5o8gi
Z/E6XIjxTD2WO/YHywQs8hmGgcYbcjHthOZArel5qDeSdbaX9z/NkRXg3R7Wiu7iCeCW6qzH/aUS
li+7O9Pdox4BBpLW/Qlp5t2P2PH459CBCpWKtTzJbUHMcLpVLu/jh0Yo4BD0GpGwHMcoyJUIwF1U
+qFoSU0hN5eYtjuMrksfQYUPvS7uyqorpqoxV2SSWj/nNUeN4wN/iXGPr22sm4ewgrBUSgUeS+pc
cFWBOz1S0Jhu55Xfme5c9Efq60Yy6+sSDz7KNbXbWTpJ4N758k08IYRkwuEJzbAo9T0BKkgejFLT
n53busuDiOBq0CEqZpThyJ3iwygmsmRUFo/2dhcHf9mCp99v4t/VNVQzp4Z/u8lCeGGJVl7JKY2O
wyt0LW8FhhTURkld0uAWHiF8260EAl3PbJS0c3xKtOUT6CIuwc6oDWWRjiZbYYpIZadymY63FUxY
kDqSgSGSN9P4N3V9s4S84RJ8e3ubvywBwyUixlBkbJ5W4VUDO1/2blXpbTh4Kf5UxLrLy4sWbnAl
FEzcBEaV7w18vCFXL6rA07BAKinsbZnptrLM/iLsMa8V4VCkQIygdYIwZHb9D3JqoPNpKLQNemsz
Q9C3glePdizRJaFfWDnTO3OIE39+PVfqHalZSG6xX3NC/yjYUA+R70GYcby3CV+tRND4dmp81ya+
ClFunLiPSrhq39oQb5QMDBr5pnmuJpa9+fFzBAcpgXoShVizHVvjA8fVJhyv4uvt7WAw8hPs8qTa
NkfcnGAcHGWnXZxqtyPhQla6PNOgYsP7rnjsc6fl18e2nbXpnLnCmiUG1INqC3Sq5CQroJBd0Dis
vI0EDTn+gM2OQ7s5cRMZZZvJetdOgH9WeHRhSRodpNUlQdO0vAOXi1LbJVNEbK1vdblLyj3SZqlI
DvIqemsX1Vozn4C+ogtQNXU3lek709JmcWQ05pH5BLcoxx3wtRwoO408mUAFSfGZQGxlJrHN+EvM
LmMxMxnCZXZP/Ec2go3n71UHc1fgbnoe1IKNexD0Ws/1LjU7bC0Myg+XJO87PqRRn+oZ4Mu44TEm
ZyuzAZagGoiX+VFt27bLKmrBX5Q32cHfim7y1XgFcXvc94nZlBgO5yPodayrNOaOfJEI4mBgczkD
gK6BFwUxUE+CW/G52tAx/aQl4eJHX5qps5TZp9L3w4U6H1Q/CnUxfT+DShgsKb079eAXnXR09Thx
cFL8jy28EXR4kCyVoneG/imD149iD2Sn14L0Yj1iBMcNm6s4IPhESHWTLQiQLnJT1zI/v3erTj6i
JPWUpQD5nCxS9BOwESN3RHsTKHdwdCUyGw9L7DgGMkr8hESwSj2t3ZJf87riEAxoEKRYVzMHePdC
UyXsSkJaDxjXJGdepB01FhWP9jwDkyUoVGVtYKTofD+fiTk5Dh6boKXgryVDzFp7NniMno4x0JJF
synvvVQ/MtCunZLImMiLVAxz1+yPhOGnOIVhnhQ5rRAtZyC4V8KPId8XUgf41SWb5OosOTpQS10j
dzTBSTPqXABjNHmnj5pNpz+YAUVCNgfTYUxr7IRvum6PQmt1Cbeb6IYrxVD0VKaCYc2BuNPAGbDp
Afdp+qoos05fwiUlc8Odaa/3RNpmuYhYx2ARhcDp4tBiIj4QsyrAyGpYc46zkdlDjzcAhLMd2O6p
U1z5GEqnuOKJXCLkc+7uxkNd+i0BxqmpAJXM7+eqKRbm3RIxiR+lOju/ImnRJSJSPHj8J5T2M1wi
1j7c9Ix1zP2cCj3fpLY4CQQk/ozcRYbUqROknT+A/LKepP9qduIyAF1d6vFub+HpSZ8cwkZ7Yqt9
1dBESopAaJ3/bVfGhMRZZXrS0OthlLPKokJmb60IHdh3cPntWCgs+UFzB7Ax+0vSrjrqe10XBPXA
No6jIe13//xyil79R4vgLJL08RrO7EcLZZ2iaw1Uy+HPsBC+h+yMqVZ7/hRfgEiRked/Q6+KRqj3
weo4xHx4BSHdu+xZSHoPqnlWY0upQXghOZtJa1AC0eajLcHhUyY4289HGEV4WVzYxYf0CxSSyeb4
OfQnMmIgh5KU3ykwDeZ66MuxRs50V0FTl317dnKqeITFotwTKjc3f1I+A5Y9ZqbxiHN7M8wMIIfy
3Q5wO/qQSR9o2iNzdckk+ZhFuxvKuVl45QbZ6PYa6w74soGAQTBKh6A9SOYMZs8EdFjgkBEhtRi/
Ylwo7RGTvbEYkqBbZrWZ5l4MzDW6Unse1/jYH7FDj0kqzT6vb66xaAMRE90yMHZL63V3J7i1tjHZ
GQ77GAmKSXmQ9V1P9YEYQbGuelTlOtNLalZpLcXrk36piNOEUvsbvVOXYdv4YAli3s5qgLcOJY8g
IFXtPZsvEYPOZpRPdDw5dz3uS2hhTfs/InC8KsOh4bAM+ia/7p5gA1IMxUQ27V4w0lIW5vp8xiJD
D4iFBBRSHOL1XZuYNDMOSkVRvfyYs2vtKPIksrI5YxBKlAgmHxK8IwsqKcww1g4PST9lHw1X9ZGO
qrt/zskfKRUdPxuw9dy6HMV6N2COiSCBQSHMlPGab6Vh7WyM6rOM3tocryKFNzsaF4bsOq8htrTX
fv8wtbNZvn/pdiDhCHG6jcSiiBq1EQ7odlvgRpZZyPLeWK8K0p91jMaVyK2pxhr1pWR4V0JYeRUj
uI3QOlpPwUpd6nmtbVdVW8ISL2/zhFqGZNXSO7PGtvznuEV4ybATks59tPQBguRhY4t9WtlO/zpB
8OFGLbLROOoFgT/r30i51Al2Jt3PsvOxUhNvuV8RIXSqjHgwz5C3jGQQUCQvhXUmGjkVsBZRrRHA
Z7tReT/s+JEAz12C6JQ5aTBoCc+XDyxMqqItXxJKBZPpVEt4viw2L8cDRHezHSJGw/SpQnjFP5ie
tLcB9kVVhpArHGb1UCkz5oQjsJs1NN8rfKYfk+9VV8o5pYMHarfr9BSd63+N4t4CYNqSMEb6ckr1
wn2dRyBqpM3VZe9WvTpaGrwbCQXYja+kE9eF9sJ2PYEGFpATaOC0Jrg4HglNBbK4fYBwfVNm9oXe
uT/3uQeSjeySEQH9EMqrIcKaeWvIcOgwaeM3rJKs+gaoyLjRD/an6qhUk5gKxfioaRSFsjF/L6E2
e1L5/vGpBEQJAvi7itFh8EpkBKjliprjvgnxRl22Pv46zhp+9Wkj1+f+UsJu6Ce2UATcTl81V7ca
aJ5x2jaLtDF6twkybpF2XYjffFZu4UQwVPCIbFS1Ct5z7JZFtzmEMODEfqDO4Cvw826x1kUzE21h
SgPxILil5pRXc7+vjuIYTpe3E6HSzFlQzztRi8W3GRS7UjPKfF6Wt2WdgAeYSIPcCwf5njDF6v3c
vb2hQ9txcBxIROkbw38y3miwtLaOFibkvjkttmcZ7Df+16a0wSvBJYKCHZpAN9Sd/+eUYGGfTT3n
NG4A2lSWFRUONgazb4DPi4jnyQbevPPcVLLPwSDziTac6z/TDxPRoVJTD9JkX7f5hR/jfRiYIkty
3SX8bLev3qwUc/D94S97ZHf/7htgIIUqi6PI8ier2WFSDVdVIpPIMGS0OHveae1a4umput2e+jjd
lkX3jJE1yr17SDMU/0EpX7nA2zAfDJ0OEVPfcq6G0Bbzlb+FglSKw/x8LhNY083iRX05qH1FNKOa
vsgpXTE9C/zvn1/W8aE90YYoU08vFusVgOO2l3DnjSWrmcQnIg8W7GsgiovKsCF2cD8YNWR5un1P
0nHfxjj7d/qyQ4agoDMGm6eRR4BMls0qS7ZHQZtpHJDSICh3BqStPe7iZkpiZV9KOnZsFZF7oAeu
+OF77oPpde2mJlCR0QZ38fgvBPHb/JaGV4UZuQFgUB3zKAL7h7IxKJxwQSAJlx58bvOMw0ULFiAy
LEuI0qtkiRdVEBBu67FobESn77pYX1+kSRHAQF9AIYsaI5BdSGwgCPngg08XchBD9Pc1KONKL0hp
xH+y6iD4MFoBFOukycHx2uRcG5XySH8uvKYCZ5LhtPKbQFeyK8ItBqmTaBQjzy69efIb1l801P3L
Qi0uPkHD3xBozArH8Hm9moQUg326J1hPa+rjL/h/tZMBxUbHrdXYJYoYGIQXdcWo1b2sgltHJ9H9
scG7X4dBGJoAa+CIqsTW7JzS4B8CcsnpIfBkc1OlfYU9Qrc3WohijY0i9Wn3ttxbcN7+h6lM5C32
bGMzwLufpAGkL1iuVSzZKuRuFNcZDeNTNTPEKNU62SwH8G9IisTnNVUFeYYnXNlpobtaxGJHFmlN
rqc1Ey7sEMgu4j5LQRM2Xz003vg7nQXR+7Ugxzj4s6rPUysoOapg39RN7di9Y4e78yVZ0I0aktwW
IMRNPz6SD6dEc46qQZO3Lx34ziGubb3MirJYJzb0QyrxANxURPo/tobe/3Kx08hkgupO9Oyg8ExX
2ielw5aD3VrdxJXNqM9evfNm1fCNI3dTkaHFnPVokr2WO8TPSavcDKlpQ/ipqYqGzTqvCfaJBXpU
W/XskQ6in8gRubQzoD0hSktHHa0+dKD94/lvBw3SgBvkmqeGWHdr3FTwvmA4P5y4lV/Rzws07lIm
tD9yr6e6B5sxthhkl502GYSSy32gmpB4v1mHzQ18QtYS9EyUsm0m374yzqOzkFaoYNLAk1I2zZpq
FUFMU1UhXb11KlHs1v7uwjAi2/dFgysDE5D9e4IgHyjHFORUNvV5O3gK6WbEDB2YNYDKxz58ise9
fGNoTY5GaXc0HNnMHuqiB+ZvVKFGgF1RrccKdLBblRVZjRSpfTQwDpatf97MFw43x6KHQ+fQLl8G
n/VqUEkTXGWp4l1fjiQKsfHwACITsEsUb1leHttvt06XO54Oldq7Bnf9CUfYm7k02lUMqqenIX9h
aojaI7FRZagWbUr8FBjTKaPMWF23fQ6EJJxRSliOwQsniuXt4/qhHMbAjuQzzKeThCRQf80rId2d
pO8GKWmor2o7kEauhoqCMBeaet8zoElW7nfu5pXBk/INdNwAtfHx6Z6HFPXutsNsdRwUCqa/L1/w
peP2AWYmSLeTTvBtQJifpysM7bAp0EQdkPT1xO+NTMWKfcF7vuPZvsUKP2XrKYo9GAnlj15VGM0z
8BwMSKHW6+rt1BCDufEY6tCqRA7rNSYYgV9XEVvHs2WmtyXlyPWCzBx0pV2VQCtWR28KJgl0Q1v2
Tcv83M2kha1ydaArxOHuVvWUDWH3a2hDQJ/VxEEWyV2y5w+HPORVd7v8PzESWt4rcfmYktvc9tsd
Ch28v6prstP3JMTrad4TKp2HaW/6RZfaBAIyOsP7L4lWXd3yv0xLh60oBZlDn2k3GlcPQuU6L06X
aUib3RbLGp4YOO5rxidCh8M96nHSYat9EnmazBBVHRVj4zax3Qnsb4FD3Z5SMsAoryyBIqX3Y/Ss
lJFPmDUCjfN7MnN7mDJTyfvaKtChEUSI/ELdGfChS8RLQnuOHcngg+jvkYywYvBtkx6H9VI9MMmF
TXL+swy/0spCeYaPw9+IIr2vud2eQK6smQI70tNhXjBhEwT4OqRxo/hZxSi3sSGnqnLAl5xB/O/p
anqC5i/iU03St+9gs9BDKUoGEjYPDvS4uR6RYAf3ZkMB1TuM6sSoq1hZsSZL2MateEiaqqa/PWe2
HsePtj0zlwYDizZuZwMTrnM5RQBeVceokzaP/746YfptWI6uN9xvnuyB1E4yzNkYNuTvbzt+aUe2
4O6uRh4GgRhYglN5jT5s/1XI3taAyExvLzMXyxhHS9HRW7EdUaG9+72BCK4B+cTFynPuM2PgCKIq
g523g0+7e5lhZy2SlnlBbdfXPXq7TdYoO7iFKIFW1ES52l+XYcem5Wukw44hN8oO0Ah2IP+yPa5B
Lwr54wBKf2W9Alna12x9zivk0ikB1g3NeJjlPJggIjW0vT2uZyojhw9RdjmbbkZMLRZdEScxxy79
mT8AkzJPC3Mg8dzYSM2I4pibBVYtJiYikJVcfCeRNxwsqj+gz/y63rJ8dXvHnkVFfHF8CWgBklax
m9At/vWTXcQG4/3n54VyiAp074KdCKK9+EgXZAQJNVvKGIet5AFsAREHaiK3WLJtEjjeYFpPD6Pp
fyNRWGxWbSCIXgQ+muPRcCvWjmZdrXjPiazbm553zjXtGq+35lOgotO9smMgL7tKzixHhcmYQib7
9vQjEZwwLPRTYz1t/9bOdxHJ4FtqFD7VhDiVeqa8aWqT9ci5GuCSfTMp4bsXt4fMhi2gXBccAIwY
2RibclCj9rEjELLPvtmv+TegmD9hWc06RSqU6jwY77QokdRpJw8e/I8LQBlmAxe85DFJIuOVYgeV
WFZ6buhdphBOFKEOybcMAmWjy8Ks1RqqnZuzWu5UtdpE1FxPj1sjNRM5HZY3dPTYMnOteqqa04Wb
5ioc7hI7BADxzSfLYqBq4CmjXYvJKX1jnm+S47Si7VXtVxfCheTrTvOFZBrnhjm78p88GaaL4LKd
FH90Hlymye4UftWwdKq5n12Q6KKklGEu6PjILYzKAIYnTPHsdHql9IyUmTQRYUaBQTwdrr0QnIVQ
NCmPQDwwjEYhQBFK9PgStQbF9WPrSeE2C+MD3/jaB6+FknJWqs3LgE1srrTUWkCOK21HEYGb+Ott
J1EEsVVdjFt19tPhT3Tt6Rro7nHE00ONznvN6uwNjurwy51SDNZGbNaQHBwp+/6KU3FMVdfAx7FP
KKH3pDC6WPP8c2HVhEVRxkmeeO7+tqUrrY+HnFo2vzl/4YK8wCODEhlvXVIxShOBf5KwyAuODct/
w4i3bltUkSgJVBaiZcamrQk8lgYSCgI+4yAPeqzHtrPgpqMjSLcWWt0EhW7VDj9OkYGckx9utFdN
K4OTMTodemowDM6m+3iQ6LE5OMGqp/0m2hjfMNDOHrtwQoxYFRJmK4tfHOdLeGSohAunCWJOWwl6
E5gh31Lx6n7TCSjGx0+QUaJs4nFlYUpiu86Jyyjhmo1bQVFnhlhwarPWSEx87qNZ3RW9K7tQW/3O
drfa2mReLOrq021Q9WhZg0+93JysV4XlMBuc6hcFEPL4dymznC3mpZ/PrUJR4isgKB7sdwsIFeEb
N8isJI1EyOdlYbVUJ05LDldjGSmfp+0nc0Zp/J/mTPL0IhYfqLt34OOFrOPawUSzhLf8WWsqf3gR
+RkGmal6kDDPa6Z72D1iE/R+Ab0QhRafFqC4dJ9kvMv3Aen4lRGEVYYN+bOf2eIJCbFjQxOKqA8/
zNedRrMlDtfz8YPrhcp3GQw0QMerdylM8iHVeBrpyYYOulogkRAa/pqcnA0UasMh3K4Ktd6+tLSO
ooVQbSE034UUtsGTJN7xGYeyQ3j3ZmjHwGshVUYJu8XRx94T/3yBqY95dTfk2mkR0YYxrVOplMLn
kmNlAzwLhFyoecDICN4BI/tBjLhkN1AfDGa10uL5c6WEbNtD4Qz9YzUGozCutWCkOiIcn2c06U82
CbFlKV91AhGwh0JWj4zPURxI+Clcq67t9NACvvjhTqB+7lfNGupkNmL5/AT940K30pDP1saA+2iX
tI8xFZoPWzU85jpRahI5z7kViIx3a9u0RIILa3MuNrY/LbNHKoUGQq42oTtWj/AkzJIOWdlgRClj
opb4c/5vNycyRXQ7nGh0vpAjtqXdRN3/eBPgJVzMo8hmLztqdCME5CXgDIfVAGLYIrBqeIPIbfvS
+gY5o8KMrg65z5FKDhL9RYO6UlF8gKsf8EXglzWzAxgN0uyXTCybWgJnoXq649sih1YhddWmtSdY
WcC1N3ZMoG90s3BghfpSMgwn0CgfdGHiZmJ7XLGmXzxS7i2RaIEvEsDHz29B+UVTei/AiGZ+U+wo
L5exSoP+jLSA8I+ET5EL0kw1iDGqNfVkcq4E2xbeKR5gsNEz5PtSTVnM/Bkd4e6mUUN7h6ODAtjL
np7aOjvCXmMXx/GUGHfEejm1js6DyA5J/pq6nzim4C/J0IDS/ey3DYtrUa7uITZ6FcE6b9ZYDQ2N
TIivBv2+CeJshWr4CzpME7gBD6ZQbYcpCyHCyGw/OjkMUyej8JpfIhyc0Aq8Bb/vNdJt4cgu839p
GlxdDTUJOFmUwtLGZ61VSn+G6sgYLZJVGKU5jPE3o/PvortTRBNBGMeBZ3gxce/H49Yms/vISTJz
IWFmwaWrM5Mm2gZD5yJJNFCsZmTCKcsIExpk1NqA7+2rCazsoF4m/vf8jUaCqEZtNAG+FMG+hfb7
gRbfuG3RfGMOHu9Ptam6QZ1eU/D50A56Wiwi+zx2DGrmrvMK+TdG6AhSO/sZS6cWLeOeMtpjqJpM
vZpBMtgJMNVv6fBsO77EevLCVxD0/VmKgdr/vmRLFsis3ETuYxaa9c/bOv2zYxMO0eUeWhI7xQQ8
a9NjwfuBOXuDBTSR8A3s3a62emMcFo9nks0nR2YH4DWsFPbAYGYSxm6L7H26b7CmnUbSFhQU2CBc
YTdafmaVoMMrHduQazYIEDi9caFWTSHrnduViU+ByZzmOFIW3/JJGLBkXbbwLbzy53ijgZcXtVnh
tY9qpnRKlk+d3UtbzdLm0pCvedboIQjklJlC+XgKg8LgtqK7M4wbJpuVFWARXjLoeADPe16YZtZG
b/5fpBQ/XH/+85E3omBQ8KTrJoS8GNjVMAQbRP2zixkOuVDH9VjAgfL8eRaPPzxila1ApBuEtA6G
4f7rvv9ka+QijLGhIm81iZ3QAK1oN9ls1hSEBcpa7ztw2B25vEk7jl3duL47yCSpnFxLArTM9RoC
Hh9MJwhoOKkouSGao4Un4F1KS7bBeSt61EQ4vMnuZPjSNfbMRx1uychq0Y7BmTaRUq9vm7UWG3KO
eMfSYBaglCJhWBzRrv9vYEKCF0vaOR2cmfxoq+BfrfmDDJWS2TknaNxbTwR7pzKSQoSs5eI27qML
d9+mytCp/6yn/7Gbys2uQ8o3z5lwCjukleUy7+t+fLnp9OeBWT8RhlWIgDelbuCNbQCGe4lAbkw8
VyfweAwfMA1g20Y8FFWqUaonm+UUyitnQZd0Ztmp5FMtWxf1vG34RaXxdO5JB3Uf6RQPj0AFql+I
w45PA2+90mh++qypN/QZuYjxpnQmK6xYEMdoyGXocgIeGlVP882KwvYJwwFT/gT9eiV+mN7LE3ph
43Am/yq/jVt4OobJYJqhgWzg7qX+TrQt9yB6Rf0XKGN04pS9LVixiGzLrK7dY35lTexUyNXURKmI
dEOcyVyTuAzcSjZreqN9t8d0dHXrTFLW7eniSsBZHSw12frPKzAKdabWQxkfrDKBlZ844clyTAaa
EdXuF6P89onPJs30G0nHWYLWNeGKV2P82Q5FdSjOH1zANzkd5qR+Yg8jzm33l/3NLQUvY71d+64J
PBCrMKc7XhGpIZU2D9wYk2L7jYGti3XykoMKnSIDSgsxXmzFNeENjLZvuBBVJPBZL2qhwU/0HLG8
pG7mypkbspiOLOqiG7Vog5PLd618xnaFd4QO1u2ODl78C65HTSSLlBHHYCB735HHSY2wJLmRSzYh
r9sogr5oFnwulAcWQR/Sg7dKT0YgS9umwxmNGu2xr7FNdEt716Gkc0xW9bRRP3Iasg6+b3NZ/uIz
D3sotxm3kcVAjpj3ikWDh4FWSoznTuhkA0JPgLBZDGG/PDok3V6PMmUN0hL6odLZalOyQDNb1zgO
j5Y54Bny8OGvu4zkvXwQwYwcu6D9J/1cijvwXXhD68+7zQaPV/gxKRsRikcBtXSPBNkPqW7cRhva
dWtSTIqznLCmqjyBLJHgBL1q70tYNIdlHuT4NbccEMHMng11DL2EoTLUXSQ6ikscL+qiAlFn1m7r
Uz/MReN4kWv1F4Qtkotm+jSMSxVNR1YRmh7uqYiJATwdzM5PJ8R+AopzaqhvXUpmZk7rBYomw0EL
dtVdbcjU+WAgXJd6zRHwntOU/sxnVHsSxLgafbl6R1zD6A36GVFQH55wHr+Jw9HJc5W2tl1VNKL4
4EcJDpDgKG9TsqOEH4RGDhxc3NoWoiK/oHLSiWdpGTXdj9qRR5o2EGyMa6mMhRLJGyyU/1MOBKQ4
kQfUMCokb6jhznHMzcAeM6jtu99x8rQ0U1fsMm1BDvsZI34Q8b3h/PZQZTv0XnCl7oLtIaWoQgCZ
5CFyIXrTFade4ZrkJ53j7Zn2l+IhVRVzn4qKD5c80ah9Vt0w5F3rZc9fsLEjRf4iDJIMv5iTYTRg
rx7+k3aE2a8Zll1je6QAeIwiGq5wGhsEbsioVAGjHoRXiYTrLjIcwGS7oS9jdTBJ633aMMaSF2Ni
uvfkNyFpS11dm3Km23xA8JVeO5PPomR/vO1Ljl3ERw3QB4Bo7pYRfhU6fdtGrxQQjefeAGK5GSKe
vK4kc86W9Pxxmo3GUacLVWVqHTd3qJ1+VXlkgqCYpEA4CkZLOxsyPuvB3cMh7wq6jWIq9tJn51es
JPGv0KlnCwaAF2qWwU7idDW9srd2j3Fc/Dkcl1ohFFkeVIGbr1yNvzixlnkO5z6klTyuEqeDhFH8
yMEezqx1rk1BSpCtgVf6DRKdT3Liei5AYsFt2euE7skZiiAki1dP3w2pUn4ex20hUfZkpk3PRxbW
LWH0ov1jWTy9nKGolfB0wehPqSXe03t27f7cnpfCtqZpST2Fa5Ctkcm+zda04BhEskG3Vs6yxyLX
RCflQDHhGhs503ko4f0c7b4OOFGhlp8vXBofxlWE64XfVNIH1ObPrFyiW+slFgMLdmCnGz2h7++0
S2kX2lWR63FNQ8ANTJkEFkUHulI01/cekoai0NIE3ZkFT6naUI8jABfbaqoA3+ILddXfJUlCCM5v
iEDSrfLt5r03+i9J5pHKWH2igFzvYnsJCPYmQIuSi+Y/Pz6n2/GBQMGB2NyhYTyQS/jwFns2Ot68
PxD4fMdbaSEA4Yr+usSA7tTT7QlnEQqzXv+NA9GBPNArgKSFe4O2ofL9mIf8V3898/rYLfQRUhqu
fCFJevRn8dUkSCOBXx/3HS9vMuYT4kKD3zfzqFXNMfczCsPxrJuMSZKciOgQc/FnzxN5i+Mp0RWw
+geYrL8zGet8FMtN/stT0cyv/rxAp0+7GvyiOOiAkzY7Mw7l6FCglRDOyY/hZaanpdhLqf/mBKXj
RD+JdoMXgQeDDTTw9YpYr8Wmrf9T3g0h/A0p7E76gagT6+Kpl7hQc92wCdgfcnlejSCz5ccA/BdR
C0l+D81SII3Ev6KK34ss0O1K50fPtW3n8LaChotxsy3Gv7IYcyF/B2K2ICp8kw2GEP3cInQK9Z+1
np5O/gq9ncs44273fo3F22mP06vWngs+hFUYaSdWIKM4GWoFiv41eD2BlNA3t8gpPui5mk8BPnn5
EFa1KJ7ojBRlysYZ8Rbq2ImBhJdGpgtBNidyFzxnHRnUfGua1yJ96mxeEt0KkrI50rHmVnYGZifw
Dyj6IsLg77Ds7ql8JvFB8GK+fWMw2FuJYtX0iIlkQnXhtBd0ZKivp1LZeVWTxKG+huSeuUjc3VJU
EZ+9jERHKvX+DPGpYmHmwVLYV9RSWEs3ad/irrDcYjtFN6fJ5BvmVLwRTdBRIXlw5QV+ulrJ89Sk
GmxDxmowR81kUoM4+laNELnwk9W7WN4EAK7LBSHTbn074pYgAYHdpKgClLp/to85cqJsQ4RkDvVM
AT024dj8E2QP1FeBo/ZzSfu/Obs5WhYe02N4hvheLa1K4jKZDVPgxmh0YyF0D9xD2G2JhKWXnoNT
KpyT4wKby9VJNsJWNO6Mg88TSVZDrrGKKk1352bCDSekArPR9DzLXACWP/nf5NCVIlfO0ITr+el9
rV36pdlYjhohutEh1U96/si3b21R5vYWz9Ofbo9q6SY65sQn2RAMopSXxgrF/vFlyvTkjLHkwJoJ
OAdi6+dPJ3Q6JCKgOIfqVmORuFX4sEp0woCm+A3wCeFQN/qipfze9PR971wANqD2FCudLA64JY9B
y0COm5BKqjbnBvUPfgmEhU9bVohxM7fAuA2IHw3gYBKDulJjp2mTBWOGm05QxhYk4YI6sMpznqjZ
OdymG7G8UUq4beWMT0JjyBCKzjmGDLZwB/y0TQxyN6DqYNei6TSNKeT18mgljvEbwXHpQDgooE3D
WLAGATB2fpxTQppCIXmkQrMm3PF9PXUFp13izfBM2p6Bx4Th6I8G/a1EFx/G3vjRVeP3zICBZ1qX
UXCmby9P32azum5rcp0Ji5akgKCDHJ9qYcx9ZlwqziYIpZ/IhT2xoPdIiZt1VrLJkSR9JX/iBE+o
iAusgn6zQlZZYWPP6FFtAwBGpHo3Wkxl4CtIg/QOSKZsdfH77yUPDZSDlSVQKE3vrTKnjjwV9XmR
YghKbZqrGs2Vv/rUNcRvPBIasPQE0DNId+ayo5Sk/qLxzOKgECPo+0pCEaUKKgtne6c1w+3Y9Zu+
CKlqezmfCfp9+b3EOAt9LcoyMA60rSOtGkIroKwaYVNnTDgi6V1vfqo6i5ZvAX4Tt8eXc2M4DJIc
WnaCA/r+DIYlZ97NevNTHWQ5CpLQQF4zK880FYOFRfk+n4ISPDYV80EF3TdAfqHrFjHMyLxsIaUE
liKopZOVg1HPWymFJAp18VzVyw6n1+ZjHILKXJCWdbLknG7OxXI10rzcB5KUsxYOzaMZLM6NUu7E
hm8MGKfUdg+kK+W/iZ2unDl8Vj+vVo0X/J8E2+JyQeYyM6NkBTakRl+my/wX5SqrQCLUWQEfdYww
dzOg4GOiBNg9tSYbOgBiVfGMD2kaK7f2hrH0N4ZiEZRpVftiOe9Ax7Y/tAJaQp9AJEMiJcU46go+
TLyW9o+PUDIkRbNYvd5X5r3mU/NG8I6w2CFdIW8PvAYrb1ex/a3TlepsfckNVT6iLRIvyapup/9u
gFVsGNCi7QnfGWg8oCwCTzBX1MWM4Jotg9aPisYYjGbpGjXc7jRa/Dep1YLIBgTQqeaZj6oGE5P/
+tYeQjAy4I0nTYL8LfgoagV5C7S8MGXdUuUFl3JPqNUC0H4Ayx1fqK18wrSyFtdvV1sY87X6HiHD
xfQS9JTMeKXCfK3gkoaWxHPqKs70xov+ASNK1UvrrsQvWynSPsRB0VHIIg8k+37W1IWGD6Y14R/C
6CVRGgxzbxtX4AYvbgEk5E34yTSNNmo/bzdCtF1aE5Cln1bQOjyJcnw15YvpXzf/MvhMx3WvHRji
2u1JmHvDwd639Yt3YZq5XRa5iL8km1tgG6EZyxgya5mOWSK/Zx0SiAMrt6z+rt8gNTdhDm9dKcMj
ftW8ksBE24SJiDnSIyivVG02d+GgUqyvxz1NvHDSdXZ/3oac2e1dY3CjxxNEtBSRP8uX6vQsMlvL
Vm3cn6cODWZ7UECTWotbIBrE+ldkglQVUDAxSeceyjk4nLAFB3PhGkfvxkWV+muQYq0k3ZRh0bE5
XnZrJdAKMnjIYN09QOQUm9pf6hiLu3BpouS+GGRd5No0e5S+YCw23bLprkQu0halV6CZJaZoaD8H
tL8DdIiqsZxlZ0M1/olx6xOsV5W3bKx3cxAdXeso34CoMJNTLSEBoA+ug0f1OWDBWT6NvWA0uN2m
cFwkiir/ni8+TYYw/1isRwTaZFXdh5Jjt6GTaKhscUxrxEm5CV5IEus0lxMytLACUG/AVk3Spumd
tveA5TtbS0YiNeHgtJIDOGtbS8fQz5vpaNLGhNNb8PALtVqNjJjnffBqFwQpd/z7XOuqZYMtJow4
on9aDndHmUcM5WDPJ8FablwTmCblMHrYp+OpvjBOeyhUS++t4qdq+0fqLjLWjmtTB3Tqjjj+nLHT
g8zvM47UK4PwMmTQ8L3Skdt0UOtGpwJTsQUz/9H2kuU836ZCYaasqrc/Ga5ArmeRS51Ry4k+DbLr
+52F2jKeQBwH5jlbeSdPodv7uHfPTDcPb907hFKuTBEHxCBIaQiVZmwSiuYH5X12q6B8gAo0tYzu
F2cM45XF0gpX5rYOIWo0Ue3V1Ii2mZbOJ4a5bTuw2R66pQZtcN8k9vZ0p6NL3xrvGLNVz4yfmL1S
1IRlcuOv/SF9weoKwqRVPKAmwLGdaLdzr1ScUpb05kR0ikRAubERV3+6bSuZkhVj+/8ERR/gc5tz
kkvpjRgwXobt2NuqTdM9AvUg7ui3WqWxefnJSkM+c5EbwC7sy6lN4rDYtRvC2s9eACb90nhizjHe
XmH6QhADadFK6zhAFgr8fHWKk6bO+Z9cGYeWcJ2rqltyOsxCFqBpjihZKXEGdBhK6CkNFNV0GWEy
98eQnmRpwLn4VjEMEEEb9W0QSIZ/CfcOrkiqYsK9ykLM3eYmgy2Ur/Bkv5oyCTbD+JvNNfKL+ixd
MtLKimOBxq4u6VN+V60VCDD0IYOHSz7D07srUP0+ALAQRQCm/b7gS/UOokV30czBKgYO8DaJg0sF
gxVEPW8T+2qLj4CkQ8HCx8vt9ANA8vFCu+ofT/YB0VQ05dxEaVIFPOHEaRwHbGIaalhSLiqmcRkV
9fBleJl4WTcsWdk1ICpTRMt1ZJjLxBMONNV6/2Yi4Qji4Jzs3yAfD9InF1EX9XRqG2nwdfm9hrdX
ObYc4yfwzmhF5hEcWSLq7LrxT4ycgnN6WPmNTFPJmpmQn0Atpq9wt46rtrrbPNI1xG71vr5q4ZZS
k3zpWcW09E5FBklWw6tz723GwhtGzFyPn0ogr9SXb4nu3blVVmxAMu7Ulu+K0Ij6L8SmiXdno8Nk
1/LPp5jceKyKiAhZPyUjBY5aQb7U+3HWfPvwqcBpS4UgKdNubVlX8qSY3SB5jFkr4SDH8YgzndKm
cnuembbYa0MRwGptZVw+2zvx1D7cTLSA/PZAKAFmbXQgxPgPw5k99CkCLqKL0UHbA67f+zSO5zv9
WknLsW3OIPqlwOJU7YtZ258qn67kEzegqFZWWRXjLa2g8/vGG7WGMGtXJdR9U0qs8/kgYOXgofOj
8BIRAy6jqO94guYOIo8Y9GrDY4HPXUGJSTJZGGKCLmFs4aQJOjimbRY08/exXcJRj5iSeobzjdR8
KkQ45SBoA1DpPfUA5qR51M/EzYd/CfeTcE+z2RBlu6AE93rpscFHYbPXph1oqoJaI4MpAwet6BDH
NHnxWyWiYNmEmxWZOGhy3WOLYxlUnwTgPdIHZcNsHH1+cgxsRbrJEzCzYWwB9XaNAARmhPRagBv2
L1K31BStT6rUyJC9nYQGqHfbsxzkO0LePCyyvuULeLqJ3uu2WnqNiHxqQfQ16e8PqKmyMMyDxbWe
6/VARbp6uYfi7PnjOs+xCsaAwP6VrG9CHg6TRCUtsAb9v5yDvHX+gglfMpFSHSO+CtzuEu1PCiyx
84zzXvHmTi8z4qCgq8u7BnssAQaO+44PQyrS8LEbpLcu6HK+4cY0Mon1o0XHmWtXxl5tqoewaKau
oyx3rrLN50iqSzGBM2zhDHPXDPzKDN7RJ+yZKo6pPvCHrdjudfqnXE3cl5xsFDZBkUG+blgqfQdC
meAaKK5rLagMDScXL124pg66nED0isfco/kUyTw2fGNz5kjnjIC4//+DMNgat3Vw+ky/RU5MsZjY
PSFe4IaOnWHEVI3iDHyBUsS8kta+AVXqRK6fWt57BadXrbk+g3KwwYac0pMsfJTX7quUxlFsWgWy
QXtgp1TT1Q7YmfHEOtNt/HXLRHumI8ZnMdPuWWBosQWZTgad0SePQJAfdfa7QcMsK+WtPvhzeymT
DFuASUZyyNLfCq18eU8M+PivL/762c2JJjAq1USqaIyS94u0Nr8OmOfmITir/26X62OtnpXMRT+e
ynWWcxzMOKi86QQXeF57B00jQc/r35jRjJYqeqdYrbRpbAkXgefWtbt1eZbZKgf2vjLQ05UKTd4C
4SyH3SRtEOXBlvVMiWSGZmKhHqhdJjaCFlmClrpPL6W8k/dKyxQbHkTbm7LLWQgvNkYTHoP0yVfL
TOZdAPQtsR/j+STky6fK4p/aLY+ghnsWCqIlX/VTMFGWqjDL6j0z6A3T2oD6JXrz5CbRh1kEnXvg
aoZ9YF3GE0S4E20ClJscjJpgxlGcHYbDFsveoH6Bq7nCycxGC9yP1my7RxAcyAMwAL+yFQaOBAt1
44c9GvJD48fS/aDy4RMUHnzNYNBI41a9Gi8fr3bsVshIlmsg6XQ7oUxELddjA4YtXjncUDI/oOO7
WdR1GVwuS6MfH4jSlT8psusF9WBMD+KW+l/ENiOIrdlQF9P147GjOpsdTpuqGG0aUPRZHs8fhgbk
U02IetsmNjAqNAyKO//MYzc6XC/2HQD6YmOCBLfHu5c8L+OJ9oC/uiTPQhAg5c2Zf+3GJ31cfCA4
SoLCh0QB3jh3TY9pYOoY9c5jIQHhSTTaY2j80mY7316uTLl8i2C/tCeBc56aae7rGCC9D7Xz9Rnt
XAvic+7HO+ykQpvlHi6SZTdYCEJw9QBE2C1yuSQgstFlj6IDcMFsIA7nnAz03L5Yef04peGpKNwH
qtC1vPyrjixLADkJNBKtzBtt7USibHTdPFSVTWIeSRy4SF/5JwC24UQOQvdWnu0xQFN0HJ8BsSjy
5gSHeCkaWJ/KEgoKWMcU4iV7J1aDJqOlMu5QV/b+6p5CuxQ0WqDvd9Ke/AL8BDBi9FbLUhP9FtQc
v//OCkyVOlApW1tGFButF367EjiMgKVxiZFfaDRvWSKsiBjDbFHpcWoFx8FAW2/CirFFzi13r0Ps
jsqDYpBWsRymPNdCEkaApy2CBBm+JmK/uFOvdG0svuq7f3EJkiIuEVE883LlFMT0mTTZddAIOMT6
qkuHtKP2gqctv/Dp2pgVqdb29aED48Bo0vI8fOaAaFQprhcdGhHy90xHTGF3j1tplPC9Yc8OyMIU
e2sELrkGl121UbsxU6O076rJien1xqhCtfdPLK7MAsehJD/bNCSZsvzvVi0SwhE8yQxDDoixvWwV
SXGTanTiguOvEcZmsLpPNnOPaOGSzeJZJZpMIhgNqLCIBI2GUW6EOFIK9/7+CfoxmDsvihmN+hSz
1cYf630pxibXAmAniXkcoWpXWcg6JhoivlmauvBpgK3qkUfoCnwJRpbLlN1vNM0RaKACJlcpxpva
pzE13m9P0D686272SydvZl0ws9l/4ItyLEr/WzciV94KjtxE/2FcivKPZBgUr9RlTFqnSi5B6nzA
icUOznB4qiWUba3cEbYY+DXjrmyG8rfDFWpHmYOe8VQZSy0psADcMEkEfurwVH2meqtAbhnMC4nb
CzKVYz11uHgzTTUtW2BE4YDDig+1KfNE++yQTOxbr7e0OdaSJP5KjrmJ9dNqhvqT61fSmmv0syEK
zVlSkU8LAOLCFtDGnvlI3F0IjAUoGM33Z96ImEy1G7Y2rPJAZUOyYKa3KVBFUW0VA8N3e5g0aamG
JGEXL8LHLfQOKVIarwpRM5AGeTp1oK5dPpUySB9ILtSAGIgSQ1cIl6L4y/kO+S/r8mkJy2u7SPr6
W6di3/8Ioblrwe4ekRVF/CgD7dCtlrGmTWvjJjqtJnR+8kyUQfUY2v5N+anM6LQuLVlenX6qpG6u
94UzOPNs5dUnEgGmXLsUwFj+snpcEC3+Q1c0aam/IwJCs8sWi7X/jEMAKzb9rTKhvBbl0De1HYTn
G7GISYZqsYh7nhqVkg96DUs1Hj7gKJw+ZvoeGofmLuqZlFLpqIeJprsgZ0P28ca1IQRMgFIWuwuU
QRKGDgJpqejGGSkVvZ2kI+32qAqTSf7ghmZsSi5+xVq4HdSnLubFyOa2hHxJITP/MRX3VdZ/SrNy
e0+IualEdno8HtYvsooY/cP5dWKbTt176Euy7+sHaE2cnZ0SUNS6xWdeK8WeGmPPIrH2vFrtw7y1
TN66R025m3lq3sKCLmCP43fB5LwkMsgGOUlTtCik8Tb0+f2Np2wy/3tsrtcKeO0hJCGsy1veGfoB
W1zK3cQYE2NDe9xlK6hW3W9QYX8Vrb/ZhNiKB09YVXrkglrCC4ZxCIHKQ8MIFpEG2MqBF3AhSn9V
0T9bWXdAFqrcINIgrMtUTQlZENUNib3g4z1vZaZW3gaafIUu3nCv/DxGdCBA8MKOlM8UOgflcD4a
qoOAbk3oRwwyfCNvg9prlxJbbZjDvZRMx4NKHCQoQvjZXOdbpl5l4vbxtrNNvzeOjJU+umQb49DL
IFvYVBNscHSNwpQTc+lJMSZp6VIJeO5gcwmmZvGeLdJ47rRn4ilrpRn89waulAOvk5hsgCZ2U+wo
Fqm6q9HPxXOwqg7PZ6Hz43UQLI1RSmCDV5ukUUUX3XFfckmf2ZJ+lEIk5v3iQakD0ws9sNngf3Nl
YZDB37xFnqU9B16gXII/dKiIGBbyhXJU/QV+FkHpIcoIfjd9ta9qrKCAfMVpCAXh3CFG2/HTBZ58
oEna/UrnqVVv4W5GsTkFjUkW9O0z7ILY/uY0o2fYffiYhjg/l4JU2KeW28h2CTnjyl8Q0oyi77Hw
araE1NQFw+QubxtM8p1agG2fMnwFU8NJapKuSzhk/k3DRdiKTlVITyn/XWguPc15qo57augPvv/h
+fP3k8r/bjVhjXGySGcunY/tI3uPJVq5FsBGw1AqsGeZL7MVpaXbbVEVsKlTp4lHHj5cKLjinYKs
eMRglpi2tGA6vqHQNJ0jpv3LnYvlHz1qdPNICmYl5qKzqw/ggQ6tsh3wl5BgoBgj6bwvpj5K0TjO
88p+eB1Gh8vuqM63mcDT3BGarh4+WGjMKe2wc6VTw86NxnRJyaNUxyNSGZNpizs+RO1nUUBuGunv
lfnPNz2hK9lSpg0vTfflYWUcB6zybpVWFHI9zEz1kFPKQ65QEkiWHSHFEF/CJzRVsIZVJtvj7HZ7
9c6r1Oe6wFb8MNo9U7bWL26X36LoPiY/mcsG9gSt9OFLO3Rfcf3M0Wqr3gp2PlFNDAE82Ra9IYmr
O/LWcUuf913laN/NtGKK8Sax0eBcnPMbRF/ozNFRAjyRJKDyhILLNouQIT7c175m9gWLxz8KpEK8
Ht/cKT0zlTUzI1WITkQuqhu3AJtND/czLYjZIeKZ9QiUnIPdetF47iiRD7Jj7q/dsUIMkbauhG9B
/vGeMrfXsTEMtgqhjdGyc30VdtY5NMiu1l4RT12OnWHqd1jeBSPSuhWK2rFsNuDcy1Qp5dtNPiDd
UdPhVHS+5FiEO/I1sQPqboudtmH/bv2hciUkTnpiE4+S13Gq0Dr5nVIdqVIy/p5Nnn2j++HasKcX
5NZqJHhXLr99ZVbEsp9s36PdjR+gXRcqd0zoLyxG2Z8BxqSPQIn3S30gqRX+w27xsC9Ty/Ey4uns
nBMp3BaFSLxdd+BXqJ/u6k96i1mF1kSwSQfZhHgW0dghjpovsBS4lsRarEcjNwFW9mNcLmeV1SEg
kCu5JCb/uCrz5aWr0aI7NN0r//y43oe1ZeLqKzjF9G2IaAY6rpaeTje3jlj0HYIrwKf1+nM9KUQT
PyVBRky8HO/y2m5KjU4xY9MPbJlKl7pT9Y4WEEq/el57OCAWhdN9eHunBvHHlNkaqNEXqsvQrRYU
OM81QTVhk7+QMyT9K+zBTzhuGMkUoksLDyLaEhX243YVQ9nT4A2QXRq6mfOrp+ysRohHI3RpBdD7
uWhXlmVhfWjB4DU5S+GQAcbDVbwe75DM6szU/bXM9HUH6jOdWUtUVE7vxK7MWQbfLoMMe6NZtgld
6x0OWdpEGcsHAxWJRzkkhSu6IqNiyMiACXwR2psc89GIfOpMUqsPgCh+Fn/sBoG/Iqx+5j3AFNwZ
oxC1QGf59hYii/UDBR6FBb5M40UgR0Op4GW1ovqP50+FR2+ZxjAdBYExf84lS9bLxfyp4chg6ka+
we7y+RV6owqTIzJdoYCsVhgoEEq8tasABX24PMuS+A4SZhuSzYVmAWHe/8489ptxvzYC7ohRDp/s
J/nuNeXrITAu4SwOU2m+WWRvW7N76GZcA5qBUzqPzabMiJmReIwkf8ox02/VuF4S9SwipWuH2dSj
pVddgLZm3V6COQ/1BkI4plo6BKELov5o/0cviyif6bFQKneWefZcWE+97kzdk/5hX7pJ4K1RC/XX
i0qhEDQaIt1id0H2Qw14NwZL3VqtYh50/YomGDe3eb5tgZJy7FPNwZ1lY2EDGjXekROCTws3LFDX
LnGusbhzoUIrThtC1CMkSRJCLZGuxMp1Rv3nDgDjf3RiQNWSUEPPi4/HeGydalAXEvSyx892bU+T
6WXVz0drLBRxkAYzscGsuSa/h3Z1ew+sdKu9qaY7E+2whX2EVo8YpAZgOe4nF94IQGVuy9/QkaNZ
X6oSOmwo4e9464Z9tjD0yYlF0b8oV4DssYjnCsu2ByBIDQyLpaFOjdt47f8JQ3FgxDJ+UK61yAys
zuszJjOwOBrLz1JNKBMCxa/BfJMY5NdUV2s5uiUmB06QQPfEjqZAwM6gHyMD7JN6+TVUQDoK8M8m
1hIk2fnoYmJQ5IdAOlVCJRfj4ivhXW9kWxI+dMLGYBZBooURIx6vIxsz98+PH+u66tT57NQvi0QS
iQoqn0rXq1qWpPK3NOUimVy2/oFOBRWui7D0H+OmPswX9St8hWPW8sh9v4zLcBvnKQhbpM5E9q0m
NSmfuZywm0WMn5MysOt8ZJZDkF7eCqSJ/VjpHnVJoNPC8W3/rKW4MbJQeaWFjva/g6Og2pyUgUgo
+GkDPS8ScLE7DJxI6iQwBtyR19sTYcApfUqjZ9zG8Bx3CKKR/Qw5Ti+5CrjLPds2K8YKtlemeffX
yHI26XtqbCcrRANNB0mTtBQO/55JVGdOLSI+6NOv8uhSpdjZteTH2fDbklXmNdHd5CxdtpWHlnwx
qfvdPKuc0RZF2Tqhf6l2J/h2Q2x+SPpxrR4q4Ic102AKFNUBhSfWy0P9tr6+rqugjCBQ3NkaymNE
RuWlZ7FxBOUECrhs2fRz8Y1IrISB7zb6i14HHPHeVwBQZREZsFbXTESXjlJ1zGj4qv0cSEj+qZaa
6bFhxJnKr8WbjdLblmEjW3T9+bZNZE2Dwj1oi1HFdVlas3LoV1wDz6Y+FWoS+5jWjIWX41SfEhaD
ugvKsqLaEbUjRTi6WvFj1gnVygnIc/YBXcddn/giPkpkHcSvUBopLkfOcwZADHywvFodSsGSKKM7
A7dBrOpYDn8TqhHfbKMfOlCTzLBr7sTVkRZuktLHsj6xOJ9intDx+dEnjjyhqyZZajxwQvCor9LT
8yZoxE1RIzMR+INiccBtArA0u178lG4dDDWfresR7MJeOYU+bL76fa6szyQZTM9P7Kr7cJnSW03C
1Y38pi7GzWEMU4QqF8B14ITzcf6xj0UI6ny+NTB0WkUO1KxmXSj3/mIq1G8d4YmxKqDLGvlbPYNJ
FV0Vuys4N+yEpC6wSbmMnFonJwWMdnapR4oBFFxQ6XOAbU2JRfQfzSs3ZROT1ei5IORqYQUuHQ98
DyGr2ArxZuP4HsErB7YVk9wqhcLnRhwRnjGScrt2kCOJs7iQ8O2nRPbS8VvhB7wbz+38YCDyISiW
57rkfjqETw0DsFcXpe+9aW4rMCtQA4D6xif2oV81ZUuIG0+ldSq7ao1TlUdc0Sx2M2dr4HWziqqh
ssSN4DFR3O6dGYSNlvPXN+CLvmvgofYLVH4iuFGboFE5QyWwjGNWDwZX/QtyNPuqbe6tX18cStJE
KEF7VsRbhy0Ek6UPWzWS8Oo4nyFb9zbIaWpRVLSSepjHmqmtuA9naxKr//BiCm2bS9KOaoMmV22Q
MHRw4UOon9CljuWA91mt8C9jSDYxBbJuHfOJr9yKcNpm8JfKLLsWCh+dk6YcQlM275F5DAdRgtBJ
MHlFTGToVSoYD/TestavG3fKL9dgtrTEe5tCC1cjamjMEel4+TdRka8iIXqhazKBj9vRpE7k4FqM
r6rX1M2LCWjZ1bWaHITEg+xce+XcHMgEZNHkfgUVl78Cfu48dtMFGHffFBeft/0hNw57OTuudppX
WRy6gIESwGD3IX6z/CCBrMfqJ3h4paD0PSki6oqX4DTWQxF133y2DJ7QsCiIpArRq10quQSZCTY6
yPfTkWjQtdqPJdnQL+uzulT7VEToI3SSuaiIEpTluD5LtRt8PkmxFXg6pOE9VkBN/9o+i6ma46yx
7F6tj9nCl3Oid0CyS6YsAu5vVz4WdZ2nd1NPNCQXppjPPlfh1QxQcRebDZDJREv61xSfa7Wu1Nbu
57OLXRPW5LFSt/LI9VGpt/B9BY/EwOpe9cHVy3XC74Fj/GbNE6JsAdYyzuJKA0cHUsBa9R63J99u
oNxmjuZ4mVb4m5hIfW+9tkQAbDsaaIpyo1zscq+xLbBw9v3d0buZmDK3HKr/vOwsuEK5GaQ3cPWf
v/bNreh6xqmHbe/kC9+K4c7+UOalxIo/+sH5jypRJcXDHPnJ4YokjZxY73pEqd8QDSGP2MveX3dY
qGqEpYyuX5nr2iJZsQQkd3DGyvOzPzs07ciaTjObjb6b+kuPvRjmDEiD0r89wEttrHWCJOe2dB7e
q+l668l819RQMHtQMdyWAXpSkx+ChhLNEpU/PEuqLGtj4F8Zck7dtuduJjJ3UfTr/39yt+sML+ta
66V7d8p+AJtLixBz74cIlVIJIt7nKN5PEs7MqGGwjQTWkgLBj/Dr974DidJRpYXvOp2Od13xUV0U
qUV0dRMl1AycRZyg/6lXj130hIp9bHtopm8aTlNkikMICXPvsUewUboapSvpUprWmTQaqN6yWCHW
e9CNaF/3xOydXKBI7hIFkWuQXvHYpRuRKlyFcudglZzRwcNvZc+HUNMosXcanShXoQodsU4qSP1h
p0MDWnsOOHGg44hMh5fLa1Zwg9CKb9VcD9Qf0PkRqIU1LRUYFE7FXRGM2+jhF3M3xcwPIggOA2cH
YFRTl+8EBIQh8ogMcz7UWZXmHPcABarTTjwt1YD9ZJc0m9FtuuZSMvdPV/kwZvZZEnR+UzEls6rv
+M+ZYpVtuip3SNtdc3KSBSDDHkiLd2KgGWtBdB7obPJ4fq4j7oyykgLBTewPtzPqnzXAzzwJ/mu9
6od2nLoe9bJ5hxRMno53tNx3Cuj/p0IoTOXlnVWC18b8QEZsruDx5OOUGFCbm1DhaTOF4Fw1D3Le
amod7OB+t5LfZ2AfU23GlS2lO3X8RfCAn9NafilLNduCXPY01VW1WKRyLb9ma/fxeG1e0bIuSWTF
oKJMivhk5V+ojn024UOmh0MietcP7HAqkL+ukGu4HBbc9Tp4dQgdSqogX+L5ucVURsHWgUjkJADj
fhlrIFt2Len1Ewv8/SxwA5IepZjAmjf6d/UtNXjNQIy0Y/2/isyWQnO/Z/8bgS8YLEZ4cdb4oSH7
bzZqmgRWyN/ArL3ScWweX3g8Qt7lCQRDVpS7UO4DHBgcxTVMM5ZOFzh2dQK4Z15goZfoT+WQMSY1
8BK6LNyrTBR8/LK2py2YmaKVgA2iYaxydNvfG4Np4vc/H/4OadP/xECT4whvVQzQCYFpp8tqlKty
rfpHdzoPqCfFH+hiO2DwrSHvhzBt8iU4ztq+BQPLmmtUzFN2wXL/sDQolohuNGzF/t4NfE/pYOqX
DfLU43iljZEeSHsIP8xm1bxkbp041BfiV3pZHUfGBS4BTgbbDnhhsS0QAeArWmdz01BAd+l/JO25
MJ/6qNEKqxgMmh8w1IO3OydhpQTOeImDmeZIv4UBbwfnfJUwWJs37JoVq+rVas6nEfbGuYzgILuY
6BdhEzZ79UBJ2tfpeDq/7mQuZnSmT7XIIp5IEJ72lstVBebUWkTpdnfnM7ZiL4dIXXHPCaleOMXl
YT1stmCSnrmjhluslZQ8NlW8H8C/xQ33Vad103JVRmwmNdrMpcLyX2L50bOPSUTNXoM5WWHRqfXJ
Au5qNi1zWd/VTbghPXlYd+A77XdVaXy1wtEHHtXDhO68ijE62G/xaewwVl1w74OTlRQgfHsVKzXq
HB/bqx92/l7dmKrVZL0L8I7RgZ0fkR6qQVOd/3qHX0DPhfOqw/gkqmUYDFEZUBqT7G89pAYjiC7/
uc8wru+vzm711yPmUGsMB2thxdkC4N2ECH34O6cZjB++nZQOmOq8LMgFkDNUYK01RZWbuupDwhUl
rDnilusWP06G7t7nzY1NoKjNrZ2/+Csmwqhh5O5SM6JDmkMjLIaCeqlRETOxzH8v1UqNMOmHplPE
gLOsyUz8W9iftJxIPQzi0LqTHcoeYvAvArOhTuZQMpxDrYCezj90/hYhpYqIEYuuRKXlQS85R0qY
yXMJdFSSW/+3u2sf5nJbzb/pLOtO2O6AgJG0BHMoYG2jXCbE1SoAEJxEas0dhLQplm9KxY4EM8Vx
17QoUwA+4hF4Cenks/7442jQnOx9oIM/L43X8w3oZxFIg2h7Pf+A2ryk7TE43lanSRwvt3/vyyx/
+c1vGVk8DXwUjKVC2r2mh0ZuVNKdL7nx8XazgF5Uho1ZGQ94PRzF77B7VxB2Ul0WW3IBUbB1Sb+Y
ISotAPvMozYuJm5OPReZfLprVknmp6jVcEl5sS3XY2KSwgfIgtmdC+/wCUGsxB23X/vdbpxO+aih
b+h149WOx9QCAwicSqR4pSvQRXXZpbU9smd6yTLkwd6R/pPEL92Psrh+HzpgmDxZYHXWotjF8iMG
s4Jtje5RFEBRvnGERvoDN/+FHtZ2pcMGBPNQ8Pu7sOy9yIRrFWFaOMR+R7ty4OMmYRSgSEC0zmwO
QDvOF6GptX66n0hvAWsn7cz15F0+48Bgb08czvlkd85D6tjr9Y16+o47uYJPOFlMRNuUQhkou3Rn
Z1OvVLjzABIWyKf5g3PAK99MQVgmEQsbceCbkNpGvyjAKTmHbxJkrkXGkfWFo6KuWiZXl86SB+Bf
M+Uyr2BNWtwuHR1gHYCI+3y/wDT/4uuyJoCI+hPWTHds2nbYCwF6kSXTHyVlP1MUGn1XlVk0+bo7
Nco96jzJk5a6Dab40EZ1Gp7t97jILLv1/bI2C5rSBEEzV9oOLXc4HPaWCOcJJfJaU7hD0JeFCgnz
nNmzyG7tjoTGBRhVEzhYgee5cO/Dq3cG3BSH/BrHY8qHRmNAvKX0HLJ/26rGvhQYe2hT5a+2a9NL
iujo1ZbubJoOPtaCL7oZw5PTA42hozlhyWWYDY3pj7VSs+F6Jua38At2ReR92nY+kfM2p5FOXici
yHNqqGsQ3WDhIvG1Y730fSU3x0ufBOJ18gPj8nCsX8qcery5SFnzEzlpNYXj/ODAFwMpFWz5m+G7
w0XnVj98iTgcA/vg66f4/1dLSg5nETJUUPl2yN8CvDcj64nTQVK7t3WCZ11V7p9F1R+5xQNYCEze
FU1BAl671yRPo99ZOd7niuVGDdnIG9dN/YEngWB0jAFs3hAY7Pn6UFFOskSNI62bxdScFw6jhIJ5
nbTlielaWtE9hWShhYpfcxFktn971lp1bnCLFwn2KwOt7Z5KdBbELPN4CI5CBxDc4NAHeJ9sOu+e
PHqWLbHW1kbz2pE7CnU9GFqmvt5JMfOIzpqL5EHEIleBo5kNvYBQvSlUSvJjSgQGaKehufb69nYa
+6ovoU/lwUEJSIVyOj3Tg/Wxlr62uQep7/j3jJwj3+3ukuUUR4V0aFg4USWqkv/8qr1izPYgsjBV
8BhRtCoeZSc00ePev6+CN606LsPrI1h6zpezYMnMF16bxe0S8mLIiKydmJw8obMjU8UDezto0jyd
T9CTCbg8S4w4Ei/GaeTU636vtLZq5TXmDZMFgyxcdFDSPSru8EaJXMHIzLyLTwOSmp/PttMrNx3f
UZhEoJQFssKHhuOtS/2P3dT/i8hO8l4K2jkS7IaakXw7xCZ1wyjfHFo6vlWwCtaRJPMo7XRww/GS
/SyNn1vJ/YXMhDVZFJ1ctL6R61I6MMtQnjEsnHMCniDlezGms9GlcTC+f1eSqxvbSZ/4RNyhFkjJ
5UoaYC4GdD3pqlcIIZgK3BIy/tWVG5+kYfs5lYNR1zSBr++n1snokt8jvJ6eeAjL6rAdauRWlv9g
e6cWFf2Lx3lQsHuZ9kSakFaE73vc2X9TPrU+yVk2Zcln2SKozU6sbv+Yzv+FSYgTxKPUw9DA/CMt
CET6ys0CXxnzKfGn84whYbpOvLC7qWGQI02qJLjIAXqoXaV73FtbFJniNkg5hVq0tzNCSVVXQru7
giUzZjbMYPHZC8NuAbHaG0VoF2rpDv1ef6QFMYAeCW/fLoJ4A/3konz9h54/euIS0SbGXJHpMEwh
sBV0FDiYklhR6RfqHkmxNTkxMFAaw2ybEyC+8L6XJGhfcF3F5zwpha7Erwkwmkpf4iR3PuRMS4wB
ZPmQo0S8FhFBrpeIgHTC3hFAAXhP8eTzvV5HZUIOhxj4+mEN3ZROYRifrHgTnsOB6n5aUrAzs3am
ivDyYPh9mliblHcLyNHEBl59xNLWMV4SjmF4K6HLquF8OwEUpNXdeFuqH9XUYa/SxKnTrJnvmMlv
WdO3c696ogS/+4gx0Toq7lG+ZGoN8/9EuBM6ZlBjR2h0j+9tZ845BBf78iC8m6qM/hcHQM5tipiJ
5kwni0wKvStFiLmxd4/COQetbfQTDMhFPM0ZgKH0kRxfK3mLpLbn4JqYp7nVGEQGmRZl846wAn57
U+RMekXOSJK35HX18pQfC5uw+3ROnsgqh2A8EVSWxWMYh/SwM7K+O1oodUYk1jYhhShWeBG38rKc
lqSBava44DVP+EBSIpwWZ0pTy+rhUFpgGGmiaiynL1s+LNBjQdoZTOiBaGSVmpTXiZglieMx9QdC
bo5zG9sHIN9jxjY1xXDJMHO9s2rgpD83rTA1ZrOmXF/LnilA1iI28BYY3eaALOEF5bCKIQ8Zclwo
aTObXp1IH5ob0LKV7SYbsZBuXxksRMOzobaNgKkbBYMVATEsVd1DcOnHaFswYatdsh7LQBrYJXhC
hza5fvT+wFgapOEQ3gpOTMhv4dDEHPmTnPMfos7T1zW2d4Y4RcfjN3/hHiLoNcq5UolKtJAaQNT3
IxYzYjWIC3N/bGhhEKPKj9ojPRueFUE5xZyQBCUdhgusHm5JruDGifAI5FXxbYveEBW9mFVIpXge
bxeK3IKv7rauwIlYSTN4h2tdJmKFHhT0uzTRLlENRiN5aE4VAfddeegQuN1wXh13Pn+3PvnUdlQS
pNqgOHJkXs5qcarhSMlI+HJsLWwwEGRBMLFseHUqGC3dDWzbMbdNvX+hcBLZ8TZbueUri+luXmEq
GNRnZaphlQLUcDVBt/vJJP3vkPIPEUz4hYFHytrZqhGR2oRzToymnms5K9UccRL1f0Z+TqxHngRk
ti5OcCTzTMoiXoeteC3CQR6iw7BPYRHreWcJ189wPboox+CbgYmYo1fk+g+Q3fnxyfUKhIgw/Nhi
qAqffkgn/s+pUawG/iL+1oR3d/ueOftUNxlDvVvXntqOBOg+dGARb10/Px80Zh97nys8AAUGW9ng
KhhoGpGll05TlkyMiI1Juh9Qxz0cW5OuoKZtClOqBfoNDu/Tde57YF1zEXaMY4cjV4uBC2r/6eNk
QufueRQbdQCi0E+Plma/DNl5Cq+Q7FQ1aw8gsgKsYcTD8Uok6x1RhPyTUrcZOTGjbM9A4rGfsv3M
W0HSZvNvM2ep+5Ig9fKRHDYg4QZDL2ctddCcckX/XvheMRdYzZ0C+522zTQ2BPVSRiwvM4/9SxFQ
Liol3g6D/7WnE6fR8FOUpQndzCcMRu15e3MwzJ25qj+g0yBxIc8/7hqcv1eKwRwLBKVP6M9vOcIs
kxsP16wEiWN0aBcn7MFXge6/6SM8QHxlwFUt+7hATXf2mfo8P9ofBwWSTBXuITPh8n4WbvICjIqg
DLQAt58I2JD5dS+drQrP9ovHr7CVJR3EEaGstZpH/0IJoA+0wzKG1Q74o63oXtPi8fXaG9EqAoHN
Osl2O+zmGf6mXYwuuZZxbcJ9ToR47jEYBPN2WdEuf2OgEo5gn3NWSG3z88dHLEorq5L2LQU+Vn+7
1wEVNp0555+MT3HJPLYazZ5yTX+2bx+F/b56uIB4YON7Q+jAApv4SA3XOBhB+nkao84tE+B5kMXW
OZi5YsB7HWjs86YUNXEKjHSgxJboUVpCZ4pu3IUGFwDh8SYsX0EtOxCBk+vlRovnKgsfrBP0yCiZ
nqff0NivNr8fRRVisnF9MlETtU86gecR/9WjgeENXRPuTov7hNhX9QbkGxENz7peBdSdn+VHEklU
HaFiBVxTp6oAdsrrDgJ9WNmx7LC1ZRagcoewQxYaRqfziGRKjsZNeU0cjg6f4S06q719tnnp3ElW
/O96bO0//adtJr2fNOEQeE5YptaeGKPvmNa+9EYxSPHN6ePA6dEeQ0+0KcDb0XKucVWAqigFShgf
1FQiGtq/nJCRHMNYYQXFeJACu5XWSIAwpOWLTB+IqGnTrAZDjZzuy2jh1Qgf2KmheooQtb5dslAl
NvJ+zgZ6F+F+GQn9uYBXFgyGiM+plB5UjstrayMpqA1KQW2eL9KP/qwEGxiWmMQwTMsrn/AHmSds
qtjYfojRwaPuQ2WGaiwz9AC1X4lhc9tdGg0laoqU+6bfe94D0lKiODx5AO8WF1O5sYHZXcPt/qtL
4YkRmn2+dj4LCGYJjpvZ2ozTkgWaToekyCUnkLd35i8f932hl28GU6kPFeHc/UO+DMgl29693w6q
BR91pmckaCtnvBVvtHjAuZlau8WQU2r96Za8xOs1nKTPzKajesw85nsBHeVRVrG4RQ/r6SGOcWq2
531vWNaI6C6VN5nflwpsqQGADQt4U4nkrz76NLdc+6U1A9sZdGnNf5J39NlrLpGbcdsZIXyZnNMQ
R55+nGkwFIczQ33KBpz4GrSjzpkI7nVhp587IS+8BVgWePdpIef6SHosP2afdgJsmhQ0rnlyWGEH
24mq8MboaQEYh0Bwpx2GveYsLzaEiPme1Jel4xRRLBoHLeTDyjMNUM+J9yRLkKsvI+EG7S1kBu4L
zZF6EhATLq8ONhq0ymrKRjRoEdy+lUPly8priwgIZnhEup9KgWpQFZQChLF6UiG1Pw3BKB519y8T
hMzIMi16JgOjO0Yz+77fHkqOSKjdPmVhdVYELqtOPOqgy4ga34Mqp5m8gQwf2DN5retmIxeCcA8V
Ysu8Kjqp3FNZrXX1uLjgnb0QtgS1yWu0Bqgp76NuEHtXq8OeQElwvpfDZ9njKdUcoqTYMlBI3IFe
Al4ntLpuenPZFDhD0FItgPJzKyu11mUj3ZPKf75lW3u6Xa0aewTPns/CdOOPTGiVfXPjG8IQvGkI
FNFl/2x8wsUFXMdlYxuXOdccVSWx+AeFn2G5MhFdWvr55goo4bGu0X9bBAEFV/eUVeBzLjGaXrRf
tMeIkKuIpIjzaJS+43HN7xvVy2o1ekZTS/L4cjnb6Grrn80xK+OnkCoSd4tZvbrOGqiBHOOb20NB
UJ7TJYvJc9OtwIGQ8VUcq1yMGlcxvOQqsIUgUEohXNf3Go56HeJCCnhAtSlrS48uf9w9CvTvykF/
XMyucfQm3sKBWU4GRJxfa/C71sJXbuXr2XUAI4EFiEpDjhRJd9KfGYllxLwacrrvcVhv7TaSUvee
n0W1UvdBay+8ooTfUngb77v4hWib7S7bemIoqjWKkvjyOHwP/bxIHheEkK65grKbDe07qxV4UOgo
nGQOkG/GXFws+QXrq0Eg2stNDFuliGTMR0sgdYJp25VeuY41IVfJozCVbZd0JIXtclp0CPdakqed
LVBZtl7B9/Ym2II7S04KDfnD5pXBOQFwvmTEuoJrTaYJMirQP8a2tcTfcHlpBo/+Z/AUbEzniURE
dYJaODsxbfyW9xfoG7n6BexYargkuGiByYbiZPTIuiZXSqp+4v9r2xBvaVPv1Lu0wWlW3DzVVWU8
8D+7LeM7hQYWvcwkFyHQbdXE/A6505crX37teBh/VKdfiTxfQaZ5gMs/HtAyQFhU0787CzPc849a
emMckDFdk1JElaAi4JFXL4sVZap0Tu/XHrNS6mYcCbnpn+8+6agoO7YFSxTFkIDGcELQGd1aTtD2
bnCqcAnOykRvUBGjtHnUyoXqySWdYMjnjUZsPQbTMWhUUh2nVrzC863u1i7do9sE3eqy95lO50Sq
Q9hXaHHZc3ojBv+ZJs8L6gamDuUKT5GTtyP4DMFL+Pis/jFtWSp22gTgXf8hHYUfuYHzrNVoBfLt
OxeYRObZ4PgYhzS4f8+RMPhcX4te3ERZfvwPqQCuv8l96L5mH4jXeCFoxnbbMj7ZbKYhc8ZvrvYx
x6tokQlq+zlU1Ioe1c96ZLU510ID0iRa4r78qd7TGEs+PNlV4b909qMPAahL6RylOE4n3sGjefSC
hNu031cj2m5SHETBFToqEzC4xia1Z6s3MPIOdSd0sVN8RmxVQcQ2HZvJb9l8d9o3d9yxdnx09H8W
xekIvjBzaCdk45GzV8rQWgAHQeV1PBqFYTArgPsFxd6Cwv0LcyX+Hx6EPW3t34cQEH+Vd4sQrCf0
ERVzjAW2D77HS1T0HwdXj6kLLWpTnDrHyGKkdkxxTtrkYKRODcH67y/koCt1NyDBZnirMD7moFIo
jnYbWBo90ffazA3lXqlREpqI+Scl/DvR8K5XuF6KW9De3MBEQlmiy4aC8ujh8V6/rlNh9RQVZhtM
9N6VVDbods6VUjgBi1YhMZSDl1b4K5mJ7nGZZUAJNVIph6t04nVGfxDpJ339s8YdLeRSqUuCm0SX
A2Xqic4wEREci1FLFe3nouHvjsK/5M4flDMdnywdZRz5KA+857rFBwxzdP9NW26ayAHi4uE6Z1EX
ETAhpvwPxe0ysW3w1AQngrT7mU/EoAZPnxl73YXtUDySAsodl8hbaHeVFZVXdlZiecPzRKll0Uph
vSuCdVbYtzx/CrZaVPC61s93neHjrys6HVwspV8a2+b/+M697GGS2NnNE8G2AXUM13LbeaDh+AKY
Ia9/7+a4o741VxxZiDY9lxnzyFIz+Y7WrpTd4ARg0yNP9G1lgsK4oLsW/hOH5TWWTLJsHxw0p3tv
uR5tDwh4XUtIB1E+cVh0oDP9yIv3VF8CZJ2GdyxbuR7ZTlAs/h5UQiw3Nl/jCFkLh8kErBlYgjxT
yRswGz17QWVEPErSazkVRfaJn2wVfZZqCrtxB2VBBVFvmmNqLVf+CIqURDgAcqY3g29d5uy+4BOJ
kL/Bbx1ngU5EEQtrSDxV3xhgMiIh0qUpesjdTUmnlcZUMBK6cMMG85xWEuFyC3TtJx4L8bBIU1MV
tyQPbgS+0Ew6uz+UxGcQaIRi8+xPkab75EVefQ3rgv37nGR7u8oyHq3sXisOijhmEtY8RJ8ZS3An
6lN0dGU3Lh5vkw0Q3UiIQeaK4atYfZQqweJr73XDzidaqo3AUDy3fsekzu/H+J6QHkvCZuK+H/vs
dQLJgu7i6emqNxKuhm8LlqppPRG9F6C+olzIc3HzaaW44Xl4lQyt7pQwxrd3Z0KnPGCgDFILpWJQ
jwOWVCZ2LSZtl5TxKCCsO/czFdWjU+mQ4aI0KpIqlOkTB5lus1d9G5TZFl0lU4R3tjMdEIePYFAf
oPPAmkjJtQrQdmrFfMUM/xwrs6RrMmxElYMXVzWgeM06D1tfOQiXIdADWPk4oCDo9fIVegNsJO0V
XhJXN1Z8qe/FcgU2KteEVvl+bxrNJSjDmG9vQOpxFPs+TxizZng5psLGe9i7mX6h6+dTRvDaBJj5
ktX9GKwvB4bfTZJeNMyT7A0/fGBM+lH038n1zsr9qCqU3GXIE83YZRTpJJ14Ymrux138izIS/tjk
a9LWIatFDBvYXsBhj9p7FYcqFoMQRdOURZawkT6o33jmLuMd2WA+jhPB+/9zd/smRxfE1dSUXfXC
1kxP6muIK1eXeuB5UfF8yWIvEaZH4TG+4Va+vdPZ69RDIZamY1ZW4/V1y15OCfa0uq5eGpAxnx1t
5uSnaTh186IIkWc5yTr0mTk0wHGiRqmJV0pO1P9pz8DiqyZCizlNJ+aRjDcLwE3h2ZVQeVCrFE46
z86EwQlA497AhkryGzvd8YpN+1r3vI0YTieNwNBfbYs2ZXWbqHlV8oV+q0hN2Z+ogp2TM2qEJGH/
gO0g8tR2wK8XtfXiNXKf4nDST6js/yBfySEYQm2oKWY/PstMwM52racPQNl2T59Y/jRjwjLx4hLg
hJMfdAGN3cWcCQO5dUDPWoMcvqA9q3mHL7JJXAaxhzUC640rZnAwrdOGC4LzjcDMdIzh7Kp17uJm
7MGBVnw7O913vZ8+tFGADvOyg7/dDFCtKhzpUY+YsCs6Aba8tP9JABnh07s/6yhaqqMNNAl4NyDE
/jdhKcSigr3apbfQg48ACPc5NF47VuYRw67LkYjT/l5yXczExt6rU0lXlMNig/+tvp+iEBeOi3N4
xiI2luGK4q93A9SSSs/VDkO2yCtQoAi0mwPNgMIEjkRUD4K6wT52IoRjT1g8m5VQy2wT4XAV4c6y
SdmaM+ew5fsbFK+JgYMA/r26my1g3epwkmG3xCzP0cFkT3MhHG7ilXd0urI66UloaHPnb0zoHNjV
eBXtRci+5uryHnke3cZWkO0cxAcjjpz5Kdx2Yyy9OqBrnfn4OL05qL2m4XW0nl0M6LGlWrGnkwe5
MlpPrljeX7NR/BeqnkBeuK9yrLDJox9ARqNjoA8kM4GMCcXuqHUgR1Q+1cDxg0O8pMrXAxief+Vn
41xeBDZ7i2xJrBppJDKqFaR4ncpSebi0u8MLkdsgHi92b2EE5Ceomtp5j+2FuLvz1PDRV+FsD3sM
l2RaDJcHPR7hnX1chRDtdGEAdp3pdB39jhmgKVllQ6PribPuxuQLck0Dxqw72vTkUIC2bddur/JY
Q3AtDKdRJfWf9bBEpoFE09f8dEEJi+Cjpnsg/YSLo4wbTbFf8ywpgHZquAGpq3vBSMuf8PuKjpuT
E02joDt0m6ugYILHtkbupfCENusQAiLuBMk9Aef59L+H61y1yTdy6Y1IVvgl1UU2ohYjL6zOFoFN
xuyxpBbnVyh8aAk2AjUZOi5nz3dLFqf87ALzOT5kEbeXYu4zR52CGNFUZSyljl33GzHMbN3L3d31
QK7fwwIWVtpdtkFWto7BvXNPI0Ht5BfF2CI+l2c33TJEX+Rf3k8ixLBO6uaCiXdoLb4nzg8dQB7L
A0C6sqxPhedlIYNzgA6S7H5VZp2ziLsgKYEzr5we1qBHe0S675ru7Y1+c0TmK+FbtRMkyMRJQZZe
LgTeg3VnvMYD2Y7VaG8w6hlEWL03cO+pyqflo6zFTq0XMH1m0JuKeJQ9oKps26lKubA4Ty8LyWyJ
ur5KD43bZnWcKhGCCsH7E7LZ05lLr1sFce/DRfqUtg6Li5RAP19iwPpMKq3Fmyswack0OCiI+dIa
Qj8jM6cmbi7TZNqKy103+7Oqcrjj3SZe1oVOBAcwiIp+hDAR4i8S7FUlmi938FeVCrk9VC+XIRMC
DpAjNZ2gFeROUghSZ65wEmHQ0WECg7wG4nZ+Y+RKJVVnoXGOQ6waBJF4LyJKQnU0IHiSINs2IVhC
hjmsrSiM9VW2Vv4/2XinW2Hp/8IiU/oN+Iq7ww915CKmVqGPaJk8Nrxvs2bHkGIY3SAQv/EJvGay
B+PdZpkuc4BfZBZUFVnspgO+XrgYOCqqdOhjQYTUsFzLWwaQWMQe/f5n/bsL6qt8gGqIXwsUjf24
wP9MdOrojEpavoT/s68GwS3TOmb3cVG2aIoeKGVowiRBuFW6IiHOR052cQ8mW5vy/wSd+fWUnkl+
0fTdAu6MIXH1ybByp7kjAT4nZOqRDSKc5Z9Qo29Op4h0sPA+FjZX1vMMQXxFZusfze63+3NCZPax
/Zs5IGxVPtT2sFsBern7+Z0UYSWZg1OJyL/le49gogFaDkrNKogeZqlxeaAKwecS7bFN1xh7kwMv
T8htzcZ4Ku1K+K4GFkAmD+8o7wT3HkzzgypWMe51tTHhX6Kp5HVKvDv2hHoTkeH3DOJSfVT6wJkr
Peh6eKxFr4iuavpXJY6WW/09+ox1qm4+cj7nYCSqX7yu54PxnHMFFjRalxgZLuxvcNeanNQSqKk5
dJWO1ElY+37A7YPYfFblJsj3yIBtC/fbWy0fMB6/MUdiDD+kRHAXpbQ0nJqaok1j6dgbluj4+3B9
29tjxZwU36PnhYH8ZS5SLTHOXz2JlTQVTktLiC+vrnuEKl53nFga1JLv4niYSTszfgiYl9jdRhkF
kOWWZzjNgp4ClM1a16UxQyxlbyWiOItC2saJS+ynp3t3qBVx8ZUnhcV4TMOnoiANpZT3yvn4ai2A
olLxKOnwxK9ivJRWnV0eZYoOHxYsh8mGFkYiUqYM+eZEWmDr3AnmDuqtgWkWkzLivZ5ZZoqvSf0B
4h+7tX0XT2Bfa0aPNiDK8bM2nO9oPAv9XrGgbn0ya/MvLKvtSf6VwHGyLE+EqGbKqzsYeyZgcCsH
syoc4iRoUYzGy9xk6QqZelNVFFu3LaH/9xUvTbHGMvXpdtTU6/bEnz/Im+/Pzns48fbEsnLSbLrq
A37DMBuHMN8JttMQYN4CQVxqxqbWacKMKF0RDnzj7AF8tcUMcuo+yYwT5oRxenFB2oNDhZc7YW4/
JzrklQ0VR5wQyYDF7uHfdeR5H8m0WlMOJihGkXPg18d52oExv3nvvUDXTwZj3g7cr4r8lFGW5J75
GPtsSZw8axe7ddBuNtCbsYTTRDHQIUU+tawlNnfFNZcgWH5PhnDKhvz8vlbVo7gM4HubweZeLcjo
0+IkOhh7xxxFChrI8lEj5F1sU81yH1wF7S2I1L3w8BuM4zWKfDMkyMevKTmMA/60NMFKtSQJYGCA
GBeYap30GdXtLZ06k+8l9EAScxzPLcW5cVlWCGjB34I7T/bJl0g+RtalfcJJEZuSCW7qRwjiXVf0
noqQJcbyjTHbSrWYCQZmUF+xZKrf+ssAYPBxyP26D+JmSVie6aeggQYABibvXtTzjWqMsNU4Q5Gi
Eqv9KcPt0JtVyTRiRn77phjBzeCVM5vZWor7GYpGceFpM8cW0FNRkq6uiGSSn6AkVijSUlf+gEU6
sWgTZV8igTB22zZ0DBgiT+RLgihNuXQkKx9bZN1E3v7R7hjJxSu/OCtSPXAdmneLfVeE44Kv0rbI
yoK1BwANAfvHU9kkASm9RFeYsgL3Ul6d/j+5TpLDQfGqTYAFM4q5iqcSJCJGKevBgBQKUwJ2lrud
XEA1gUoDtaqXUbUgLywLak0tCBPXnBWpPduOMW4Wg+LoXQkw6cq8piI3tzoOPYxH9vGeZUg0BxW3
OFOnkagwU6DL5O3pyRWwMUcIF17ue4I537+W9G5DTzchSep31TGo+YjpAbik2KC5otOqdVpCdX9Y
JDVgPskQZPrCbKP36GvaVzUsw/UtjpKpH3EAfJoUk222BfPTZiDjxmVrE7ZpkFQOHEUt8tI9WRAn
Bt+3qQmmb/QZINygUQaGxJTHI6PA+2s5b6QrSjiFOTkrC5OzrdYh91MdfKBzDeuHvso3kWm+ejdY
iqHQ5arElI+k64XNjBjzu1aseuEbkLcxiKgSiKh5oEVk7FPK+Gi0kDPKoZwZxU6++nldTvrFYYNP
Qgf20UseTwYPryJXkJSTJBRuspM9V4Os6KtfZ3wVJA0ZEuTohXVj2YT3II6GxryTkSstL/4qKir8
NmrSWCG8OVpMF/LRRM3URLiXLC3ofIh4SUcUcuIJN/QTU1S6pLm0rBJcGrhRG4SxGwbWrimLBz47
l80hEMgd85S8oNXYqyolKDOQNToIU+d2VdnjapXjJ+D/nIcAvLj+6CCQiJ5QQ5l9XBarWioZ+loQ
iUcl3Yhv/xWaIJBQqVczW+ekQpdBgWq1lpR3ArgT/hZSsVDL7sAY3LbrquR1C1OVs/QTLEZ7yCii
w78frLoVJF3TTbMelIdUwmkOH840dB9qDdWbCO6fAWQ8yTSDMfmaD0sJ+BpEO8W2MqFXJ02znL6x
gyh27YWx+P9NL5bK9eHC9DNLJRmliJUAl+XVSeMkhuB1Jpazi9i1JyMAGDFuSn+XoEwIanRDEFjz
7ApZRkELY0+k+IqWrLVFd1tW74TBFuP0s2OQx8LLTpFFsfAL/AM8ehQ1EncN07kHRDUuRwx6f1vw
vOIOv56yesY+EmP/b5yqwhnXZUGhG4GSln07OzFnLvZRv1rWlaIhSnnSNRnkU6iwOTmB5aua7a0R
nCXqpkTnruNAAuS2fMJ/1+CENtcXGI22mNCcKOhFYg6kow/be9E+lSAZewmfLNEJlEdHOCmJFSL5
0Igne32PpISZ1Ioxc2tGXAIKGGPIlJoaT3I8icNudWs8XoXgJ3N9k031OjgmPJAvBzcv+emsyFWS
ckEkf04SvFDcX8j1s23J14NAL8Q2c2XQ9rcUosKC9ObylVQsn9Bgpm5Xnv/jlHUae0WgM6bWk2wx
mQq9je5Z4uWV7Z+wwgvpdTps4GSBc8eBe1HLygwJ+/HRbEZ6hmiDgnQx9VgVnWwpCcY+hl/J7/Ci
XO9vbOksE1nQt0FikL0TYoqkk/VF4ItwojY62gzB9qA1f/YlnTnGentnb8+72uSEsp/slx/TfPAe
DtvtLzxbcuM3C+UiJgGabNeOEa+ozbW96HkXb9jqfkzV6UKLI+qf9Yi4Bqrh2Ps1th1px0WTEL1O
fOSqrVDmndzZu7blxgoYkybkQVsGQqAaWbJGnYF6yy9UQonV+85EDiuSEr3aBVdsC33N4oZ8puRV
N/NMwPZPqDApig0b+D6JviQEq30n8Lm1QzbIh9KcGehxobUOEtrLdIGD9LsWbtPznPUfSZShZas2
QSvUQZN9kP9mPkwBjLLpFrU313rW19CQtu24HiH7KIrgvVrGosC4n+dg8AhhtHMGOH5utkcqdmFU
m7I36+NFMA7XZCZdZA9moiCQpKE0YA2Ue4/uKamBwvYubq753W9ZgQeVVep9mBZeb8S7KhvFolzD
q2EUgumSLS7j5MMKgMH8hMSISKx8P3w8q6UMzayqX+Gy4dO8Wq7nI0u0xXbLscFBK98l3O2X+YjM
Ul9LuMMcymYX5sqDSXDOAiGhGR/6CUOe+pdvaFyFphEM8057tKqh4uJSvLMAeF6FvN56Rdy4hfmB
fYjXqnxZJWv2+9dlaDB4vEbrWH79kTNFSagO+m+EftfHKOXaDr84TMABNpIFW9228G02Z8N0Iim8
o74X0BED7Kd7Gj7PnFQp4U0tqWVJ3/igMKv5yV1JTTJTSLQc7EMWIxrYLlYepUjQDoDosTpXH1Kl
t/OOGRHsnlLERkaCCQ/NgsAJkxuowb1XrcpHR6rg+unkOl22j8n+vW9cl+xP4rVNgFekAufZFgdU
OiSq8R+XGbTfCE0gQjxuR3NF9Xxr+2/jKHacGaeaodOQz2GxYPbj7h+4fb3zPbem777m8kgc6Q/k
N0oV4BBIW2lChxFsBv59FC2mQT3kmCjpi08/hGCqjnrGjMBKDiz4DoES9dvoohf0IZB1EjYDmrun
s34JxXYQzePna2f4AGi27+gRNjJRfo7lfOTJagZl0LoeaA3YlA+xJfx/GZymc053ygJYSMwTISXn
vzt0h88tjKULd8GVrGaGaKrDFMZk7DJ1HniiScVNzD46hpW8tRc1Povg2Mi/KUEoO7q4sXHIflWu
bOurGxN+2bzU0IoizhxtV3dFP+vZHWbedJTX7OGH4ZZZ9J3dzk058dfBCCuR4/X/uezMxSoca7e8
CkCz/9qYJwrMhJCobImpZHtQOzw3NtvL+0dSkgqAHnANf3Ob4njRoGVlGgX2psxw5gApryJK+ZX/
ZbLF+Bq0Jy7B39d+d9bgEMzq3OpI73pGbBasSBfXBor8P7x+R0oYh7G7ET+rjrArM7ED9pIdwW+0
c3aO8Vmtu8XoozotayID8YDkf7yxsg5ab6dHrzuTKgarTwD9E+thx49cIS7CKY3n4s3SnWroEXMl
ORxcZlYXitUF89vTupyu/zE3dOnisYLRjLXHoR/vcMc/mgtN2EbdeKy50NHqT8eO7bgS/N4scpPi
+kH7bBC8zzNOs+nQUed2FMEAj0vAxqC/xTTl1bg+hyy4e6DtwFj821J1o7HbEEbcevD5z+72hxw/
uChvL4xdepH8o6PTN+oHGzYFGBp816KUL3XzkqyKNbsK0X0j+ibvIyMXBIO4PKmtizNq7H+kiJiB
CAvXjdEE4CC83siqqkHg+JAIFNdwqBpv6278vdlEX9gNwcSdVfM7JE87tokPg+EaAPE43immzNG7
PEDGt/uCoYzRzpYErjXUnGpzpwINYltVgNGcTRbUNL+YIcub0wemA1VCZdYX4giCPLCiKNIkcYHG
3j+GX8NRUEcuikYwXqY2dI3nHWKsOpZUsrcDdJs2NoNpSPWLTEYgvSSpO7rQkQiXgTUqDL+RIK1d
VGM0UMYky6oh8yeoVPDkbPOmenIhnesJWwh2IqlbkJaepKBhmh/LjWQfjfV9tZV2DbwW01ucX93s
i6eB1nBIWhmMAlTf3BTCdQFn8IKEzJjq008OO0hIXfWBE5hq2nwGsH4kYaRevVYVOpg0XsvkDYiw
1Mo7VhaXUobfqggF/JS89ppEXSlqEJCKBrZM34GrF6EAqhxsiVFsU2b1FsQC3pAKKnkNUyQ2EzBQ
uGFlqSMe/e0pwa+WSsCvAEWdGInqOOmkmvdGyhs8ZA4wATvQ1Kig/xu+saw27J+SjmLmCnkVDjO/
RM9rr0Qh+NeBfFpz+T4svrf+BxnvD559jonmVVA0ok66ddYi9HrULlWv/HpiT3DlrWODkSVzc0+R
gmZrlOxGbfREOSijW7CH3xwh243OSYAjl2DZXB4sE7GbF8OQObqHxfhmHDxyw4MspUyPotR9If6P
pUAUbR6C/FnAyp9MM95Cdzo/qXj0B28WfDXpixWvgizIm/0XuJaKHMpnsOpMpRQ3V/Uw3y3dBv/9
mpDmfY2dbARVv72G9GTteqqb4KOXTzHqb/uBg69jRx08doDUHfAyf+ZCuDyXfwoSQdBbziQiAVl4
5moMzw1Nzqtj+nybBWn3pmP93BP9HF7mbG5WthPrXOLcWxhVOpE3Yi35PwLeV0/P/gIQqIyu6MT9
Sa+UwkYFW1aC3Fzvc52EfUU1RsYhGR1EnljNNQEqDPxvjxgK60xEyBBY9bSTW9AivXOTGK3yOPfE
zan/3E1Vu+GFqRMYOluWLKGnGT5DF4If82XVUWVGgVtE1Lsbjo75QSY05Qdq9Jofg/vLiicHsnd5
kM8XSoxZoIjtPhRmuM2s4hU671rcvzFQdffMH8SrvuICAtIPt6R0/CEznhlVTfuOCmMNUnvJVxSq
rfQOQthFCFADDTeNOS7b/qVKHgh2/b8sl6Q2O47XzjWE9O5zIx0/iHOLfcI4HvxLI3V7XTuA0751
grq+2roqI3t9pL+73yi1WbtLVl5ZCpdsN39IUxNCI0GcDtA5jMDok/SwbhKoTjT8ATP7yBwWJpZu
dvAdTxSjnXHXC/92P2SY98np0faZLEdWa7h+hl72fgrK86Z+HdS0GMUUQpQ3b0r9frflLHATlK+P
CZOfteYrRw7Ty8kgchURY3V7O0dsT105rcAfhI6aCpKUv2CNkjzX8+YF840BvukoYUgCNYVJzl9o
O842t1AQfKO/QpbeEUVSlS+aBFr371IBcWrMtKdSRYhnXPlzb8vNARRodmuTOqVNvNpP0U8xEDJo
vhk8vA6R5+9KwhGIhxyU76A1jHv6hNi3lNxsjd/KfuVaoJS7AX+xGLhGTdmn8UxsMjrnsV1uGItP
4SLGddbSOl/9WLTKhIN1nFz+jmxksvENVq8oUyJsps2cAWIKtaFVbCdtLuZFx2lTPMEN58GCpqk2
Bunoi0K8TpvJQOaxEG4lV77oHMrDJKiUWjkO22pbBW3aGke6jM/s2jhVPtqRz6ZPW06PJR648Xsi
1kdxDRo8bSeF1vLUbuwKeftPciwvCdmBNWhu3uYx9kBuuWKdXue4NCpA483MA+5dqcvAZVTfE1L2
qH4Z36PQnsnjCwmuxcjAQQbe22z9++5ge70LliwiTR2IwsPa18xfBegjFbRA4xnwWLQk2AniC5k7
41yvmg8tfnupH/o3cfXmY2bd/5F51Qg2r4URhh4OQIe/7bJpk0A5dKiHz4xS38krp+mDsFw1NgIK
pYsGA3g28s3dOjHw10SkPgfJIiFYDmI6ehYCgqmCuOxko8mcX2viPoYV6uyRvMe0LOhs35mDoVUk
IJkjC+74lpB5CuIlR7QQHC3soS0LTLuxKR2Mj6PDcV0Yhlb9m/qn2eY/3fl8KsvQwyu+m/biD5ML
s6s2hrFYx5haTG7NLVrUCSpx7BmxLeejBxtQQ7mzF1m47xq68JufJcoemxjn2/M2uIoGCNcIxzVq
NsG2GLs/lqRoVInlg9NahxuFYvDgBbmA+lGcXD4b7GzrlHd+pe8rVkC2kliUhD31XN9HzaLDAO3u
dc4DDqKhJlmJC983ghKJg4nWS+Zx060vOK0MWQBs9mSn4wfcO8DyneHEG8CUjOggCXkrgFnQMxcI
U/6WpHmLfipKqOQ8u70baxHVv6YzKxT+iw/J36Gha80si1lr1Nc0sU5Zwu6x7JzveJV0/UgsGMvW
ktdL/7PizcFafHXI1+REraHq85GWhL2u5qYHUhJ1585BcloNIQd3hT44svQOOS7vwekMcQBMH9j7
9mnoIdGXFRpq1tvUURsk8+yGcJ0hC3bV2rKrH7vFOmLZd1k6ymY3cYZsj1Q8QvpwlfZMwJc0Ikny
mQoMNNcDTvZZvtLbbONJvcxYUPn7xQkz61PWI/dKUXh7brr61yCveUBDwhOC8lYgOnR2ZZWelF4c
MbTr26sry10dme0AjW8CuvSyQzntOMCFAYlOUkBUJcjPegHnoIBG4Z/IUmDYxVO0CA4pvdXM1xf1
HJfV6XEy+VtBt4a1Em4RT+7bNVENEvsil4WetGAx7g5JDSWdvqIKh/6t7EL1XgMfqJ8E19lC4Iy2
4hnV2KyGeDfXnSDaCOjhFSWlEjlSLjkrny6BKVxIa9zwORsDoGJo1dH4/u9/rs5i16vTuHj1XIKS
r0GgK+3V43hihKykhkE6Z1ZE+nvIS5xtPKmH0/HY0wwGFdBhy8TXa83bzpR93ty+fYYwXV/Vfd0W
Pc4EBqeCrUSZp9pez8TydPh35y7PEy5+kLZZD6bcDZYuRj+RJ4CzKIXiwdaa+xGe+A/OTWNKUwc1
yxFGaSzKtjtPmjEiD7dszb8ZTtSXYbMsqF3totWThIdxpQDQO7yDl17NH2kW+qo95eE/g3chSlFm
iOg/miCei+BqWnR1G9+s23I9wTc68mHJp3AWtREtZ4DZ7nn9XuxRG9+RS8+I7G19CltZByK1WMDu
0zbbJHGQLnZEUw1721nvzHUo58jQrvwHogkSuas9A8RocAe76XC0VsJTuQazXDF2KpVN4MhNCHuC
RR+sP9rCEwh/hJ7mj8q/8O5S1Trru4U8/0zRO8RAWhGqxYt+EKknSNjvvG0Ea9elEoJcelR1v4Qh
UoyH0iw/5dvjupuKj9ZTdZhdYYndAK8ePVVw3tVscUNuny5ZXI25+sHqnGAvZCsVmQUbVWdUqTXD
R5n9qrsYNrUHRpmAXAmXCKQ/scthg2scWE8+6K5P6olsoTxuJwZEyMSRkmKCTRoNbOm2/FMkYXot
SmvQ0hH9gRq9mxK93zWYcHxc/Uq761NXGnM9dF69mQyGNTRu5Dzs51ZuHsBod20vcTRq5f+nJAaz
3fO/Dxy/xTYrxL+dIEBn/0jzNicyWgvJEs4X94sTWyCXDjKIqXdG0JKGzG6VQXLzuPzvixLFB4EQ
aaS/AlxXnKr6LCqMJkyTe+p1c63HKNqWWCLfFcm+Y6gktkeP5g19HczSp3oGm4FHjg0t+fa3MDrY
TSGmMbpuyS26y7lK7cicXvsJCiimIBYXfTjgHnKwIlAVHSy8Tjb+66OF1dHfCBduk7f+cb6eLeNx
ftXqXXWTyJEHdE1vqF/PjtvbMI+Avy6wGm5+yCGdif1tNEFB8rxOQWp1g/kuE2d1ASQkAL29eOX+
P2QkCX4Fft0+2Afzgp5AdDxj2sFSL2HVk3DAzyfM7esNzP7Ff3iqcRAwkJf2DTTudmz661BOnFGy
KgRE+FcOHEAqgcdQ9r5hI84uiF6v33mJj74pzWEEf6CkvBhdbceA/mIKVRcECTeLi5PzZV5sRNXw
3njsY8M1lbAgvEBoPbPIGg+OHIkh4+vWMVWnztD/4GRpcAkDms936TFCB2kNUutxwVw7uVEWcbn7
ZPVbEieBzGL11nR41y/wcYxKBvNZjZWVdbHSaILvCet0EDMnGBCUuSxUbRG7v28UXkYr6VYdDmkn
b0rOG56KbDUvV49Bf+3STLgUNGtU08Id823v0Rlc26XUKacPZC6/yoEoc/y52Rcpp4mhmDBMFEZq
VmPLnFHK21ki6LZV1vnnPV4gOj5GJ2/uoWIXZDbeKyzk62edvv/hh6FK0KToqa1KwU59Uqr+0jDt
Q/a7LWnldS6eurcGgvvQN6SV22mj9INWIoUv+bPRWApuv0xOmOenjq012dvBI9nR5aMcxNB6kCIV
qbjLrmfsmZBiD3OP7tyu6PxBRZIzEP1rZXqtWv1cGNp/5YxoYSWxHtaRO4PufT+6Vg3kQrVZUDSc
Gj/n14u0gpe8m+ZdaCn00Ij0JMhfO60Bezo45/tJpWsCu354Xm6N4IqHW9N6quH69H9wo3hXfhDI
ChfuLwMsodRfHXfyujvUSpgGObBAUCgYnxBC/h3YqiNem0hO6axxBtrtokq4f0qjxzNWylQwjAoZ
d4UkOAYOYHYMo6I/bpW4NUBDXFJy7ZSgrQ7DEfkfWs6WNX5uiXdrPlq0G7+yAdfT1u9fBMPjv4eP
RgUHNSNUQbFdMSNwab76TSA8g//wxG278bWOWPpIeSLv/fRvCtTLxdnvZgOlQknJl3m88C/ofqrf
BcAhr40gHVkF3Jkf7okx1QWV8gcg9jv/KwclbEcTtFCihLeT0Wk7TC/uN093qAnG+e8KSNjuzTcJ
iw8s4Q7DdrqE2U73bZ8OK4ZprGVy2FGo2jRFMuF7Nl7xHcqsTdk9jlbYmixAFqmncOuGmcALgZ9n
YLnuQ5tzAQ3ACFV0DOfyjrLKyaCFz4TAolJgHpSQoXyqKcO8Hz++hfXm1oLdAnBfY6t8zPaxd+6u
NbPro1LSjkwxyAZl8EONfW6Q8sBvjjXd629CDVL2xPJlm7kpSTSl9RNMca3Tf/BkN+2SZ/PAzlxe
pbYn6t7cW0erLtWZshhGFZAo6YrTm8zExG0TT9s2wl08p2bxcxi2LUZ2WTQ3WlzA3R3N2jsM+GXS
yfhY9b08houmKE7AcIVnVBlCFTGsubjXdDyGYbGdUhGLweBRWsgfU4q86KnR83jdLU2hIbCK351N
6nu6VD1FbPhR0FxXUPxs0Z/jEwuMUrffPKDleJxezeHQOwZ4CbE1G/n6vNePpG8om+AcZkYyzY5M
dwEvnuj+y/OwRECYgpG6d8qyPfawpauDZaBzgKPJNsPm1Y9W76j0IPzFuA1M0S7LX3YBxag4m4Bj
KQdyVSQyABNfo+XH8GdVw0WEGPlVoDS9SfLUZTkahT40yhO1x/YKMqhjoc9pqURVV6MluTTsVnhu
zGsr5nX3S7KdykJyyYheXHFVieyBVoNBhSn//hEch1gkAhc+bo/2GvB96aqHij/1DlvQk29HKQQJ
31U5u74ND/KBGzssXbK84oPsbRIO406Nl5rnitlUHxwjiNQL2cqYmCL6sQ4eBMoKxomkwP89SnF1
nRpo3i0MkHDHFYwFRd7bL7B8lyDpnbPBy1/p8n7CyOGMxorY+s7PLTccDTAjBMHtkpSwqxfM7Hd9
HvPPx9WipcT+X6S7CxCTAhec5wgSLQXkZFZlyWXSUMUEuX/Gr+dqmT0SBd+R7XGlvQfdX5DcWjZI
GfVubvH6B1EO9ct7CFYn8PTYQg3JCxQu+QqrVCZS/fwJ58jEAHDmh2w7ZOipqVD0qlEMPOqI2LDI
kAx2v+GAWiKU9hPMkhDLj/jiBQHG66//Q7vMkjb2y/UEnDg2GNCmZmCmr6GES4NeDJ6qKiprHhHd
u06z9hv/fmJ5/h6K1eQEh2uZOiPOFdNd11ujwE2QsFCRVj1JOV9J8dUuciUfODCiX1fvhjw2qk+A
XctYMRbpfqnZcpuP8llZBNgWx+C6L8o2RoQzBL4fOW+WMGqC2b9oiZeAD4jnNiZRIBAwOplOp4Wm
mlmCT+k2jR1wLO+DBtJadJ6ma4YM6fJgYat3RPM8Gb35KW0X6//fPB1Od9F2FlAb2BcKEYogvs9Z
dgV9g5O2uvbWp/uJOv/5D5bDFoKQrhwo87DZrnNIGo+q9s2syTJRubtKZxXc9Bk4RFuKvOZyPoD3
NceM0/8w7SHDKtgLl/kynCVURoQiRH4i8SicdsgsEjJ2sgNK+6XsJBYWOh5ZNZhyqUdwsmJ5/m8E
VZx/ZhNnraDIZjAfXqDGhRMt7tiKo36gz3S4CVc2p8IvvqatOzb+0LmLt3AJsgPiRHqk8n+0Sy0H
QSsnzRZvfQLKAbNQksX1Jk//10bIRKsnhNj2Orry/aJH+GxxAET3YJ5fVTv017qMANEcKrzSsn4A
/8Tgdl6bq3rJoVzCLTcpnToJxXeeFqQynl9wZFoyZNB+X+dOQjFGdUk2pEhPuFFnAGwoo2U4iL2e
xZ7RMHsrSGZyCw26tVWhvEzy3ZlduZ/djfkW67bfLg/77BiIV6c3x9owYbmfwxgURxHHZuBjS+3i
wO7+XAfmYh7xtaaxPDPLY15PIwuwJWAdZw9WNB7CSRzNW4E71pwoq0fNLDDqnmTtSCQd2Jb8U+x6
8rMgIlIN2KI9WtNFLt1IENtY4ucEkgc1NHfxOM2O8ddaTpt0CDPvUttywaKIYlElLJg6GguILgy2
DXGD3EGh+djcVnga+of+axEYnc4El9zcKdFVzSMpqRrgrbYiHGUzctJXdNpIK7TrgsYrGSDDofn+
cCoT0Mbvi/P0dZX5I5yg/qoWJQrPHyW/KTr2iPG9qd3mj46gqm+tzxVK6e70hdQzDdwkhjI/J66J
W93y539ObuqoyNREBPLPAGTbi2oGMI/5tdLVKtjKAtEDzCPeykqLKt851ggonmsxToODZEWwI8ml
TxzJCqV8H/djNVkwyOy1SYrhsEmN9LkLLIxyjJa+5lAjzwHZ7YX1Ybi7c8eXJlK08GvwnG0I6TRp
7WjkmEBpJyzovtalccVFwuGty6eaVkTBCU6kCS94Rb5jyGueD7DG6GnTW9e4P4Hb+yL85DQytzpR
f04E849CjQxN6xFkoku4lFVCqg8x0EnoM42B/AA3tdxpEbGhgzK+wXKG5eUK8Fzj/MRftnhzUnOf
My7fPWKnFlXJyhYkOLzYg74MV5EkjmD6CETYknu3RSJVDUN0Dst9ffvCbiijFGligOwlIT4474qT
3gnU4vxWt4/s2fwVoGEvx4TVCFlAGsdlaDyflOhlwg9OwmqbTdEn0O+77z++S59xF5IGvrafE0kA
cPZSX2FUNXaYQLWbgKMSHVwOrdhMvFajkoPDfRcpdeeR2ldenHHJ8SwAIj8N+O7hOeYbohca34+m
9mKuEce+exiauOm1R4zTyMqdEbm0UA8mU1gYb+M//KaB5xBlQ9FDJwB2JAiNZq6DV0e3gTzEjmFE
xCSsw6TSWL6M7SdDjC5wG+4RxuwKT8JwcfPWyU2AnjZC67SeAgh0++93ZiAkQOlYNwjbBfMfQI8Q
wuLKA+olJj7+vTl2E9W74SL16bItg2602PATEhry1CUPIevbHE2Bqx7Jd2snSLh54H9mX1O7do9G
LmZzKpfDtF7U0GMebMCfkYb9EtPzId/ryZuSBSqcBiBSPGLSEZh7zdkMwwn73Sr+dzc+SWNVK7q3
pA/4TGfPJtwccxlAis33lbBdaSTQl5a8sthn48v6NPgrNOXRGml5VOq5sUYWE8xGSYD4hOSKVMqJ
xT8FxPCRd8iKAEKptjxQeGm2IkwW56IOowvfCI5JsYSW1Z/Yc6OxuF9RX9RqCes6GdsNnvFh2Id4
gPr3gy/0Iy9SkBKQcxGPIGZMDj41ldpSXq5C3JjymXatFupILLBWwvIOWViv8UtCAaKXs4F6ibM/
lDhMq0CAANhp8YXzR+SNefAqUp/t/P/03tN4eOSeV9r4KphMiEndUTuIRilBRQw4AZG6OT3suyNo
SAA91RdLT/54pK0qOjzj70hPG07tZeJE+QTCAiUoDNzJMPTT+FIdpcrfrrBruP3g7J8IyGXAE32A
0d29XiLsQK5c4rso4ia7jc7CPxn5enNUYjzAnLgNGbWNevdxeNALNQA5swgdkmwmgTIBoP8viip6
wbxIvrLE5Glaqlh9K3z3CSo2oeGYYIuNT7YWJGjHO5JF3yRclECUfarJvwf4YaeXxbR9XzzVuHdl
5pKjjHQX1zgO1IrbOq8XznzJqbTuqjmHkjDWe81OwXrqSgrL4r9Y33FlB4/Zic6QT/lTKFhYQvre
oIPSfLgjU06SsldCfJtPmDIuTHTmHqYLEK+Ggo8g2viBtTR1/NIbGYmf413hXO7jQuEdacQ2zQjt
olr1SyGP62QCdCt7dBlzuMVTDcrQpIx+ervDkRweGJtNpveuq/iq4ErjkbNdarS5YkUGyYVwfNrD
dv/5ojqP0DBGii/M8rBdf0+H7CxCnofF/L545qrryvp5uQ/GYEoB3oOy/8+XE55bORtX14j0042F
k/27cnF/N4vJhfZyDVu0aR413Oo1i04D1jVn1mlJTpMCoX+PTRueI3Up+5YdhIul5uhqS2WkKSRQ
dJBlFwxDJg6vJCks42OAAoXlkwh1sJhgQLN4P6hoZs/aS3j2yuJHyD3qoIUMyj/6DbNCc2lLzPmT
ru63A8U4CGy+HMHFBrHw6F6ant5qxq0766hvL0K2QldMXAlFMkDTq3h/XEtc0QgIUJWgbTh1YH2m
MyU9RBCTXMCKHU/91o+K5ZqXQU0jkjJV8G+FBdQ8CSA4OwWT4+LpWE+IfhaAkqURnHFZN918FP04
TROAcCAthil/kMipr+DihiBrZygA/qo97wbfZGIgVvfTkYoABbljF1dOk259Rruuun42kBw/tVBM
4MXEDAr+r4zlZvvbgHrzrhcoy8dw1nHKVxzHxQWk/bnK/DqJyXBNOmMBZzz817dCRGFvOu9PWBjF
1UxUtK5TvBM164QdBzx95zoowCZyC88FW1tZBRxu2xk5wc4+rJfCLsYb5tDYwz2sW4gdK+MxX/fP
BT2NPpLO6NYF6dqW/c7y9ZsVWVn0HGxQtUXOTNc9rh+FV3whH9gFuYEo/drS1QNhJdbq0O1x56e2
FIk2UBD+mSLCnLFPPCNBBGDKba+vUDE1QSckrVrihOyFVNFrprQx6ozu0J2Mgl8nciBgywv4901d
j2/dZCtgXyCo9SZOZJAq7rl1SkmJz/IiE6sQS86B3L+EIEIJE7qwyBLrxDakgMqwiDWFnNMtq/Z0
xV7mZ3HFBu16mMo3PH3CfkIePxPVQDbpRWORJzMjjKIXOCA1TA1f0WkrK5qruxECbaXj0YJEHky4
6+l3xdCZP3WP98FZJhQsgpY/JwSEOVG2Vbso7sabtYXQ8RB/OEqbEXAHknlfefSgNFnDa6j1yHAq
jo3jBs19fbOswkLdjiDnZMnjs+6gD9yoQdVE+6D3DOYGwhPmOX0kCvg2qshX25+uNNH8hD/JUxkn
GN+o4XDHFD7rWqLT3B0pSzhVP78misd8/JziGnhwhfYjFs8q9s7i/UuuNqoHKMf7vZ50Fwj8PBYu
3W/+cwI+Stv8WQm6+K1a4jcgl8+xvaDp2QEm9/xa3eU2lNkxn7QLPRM1bK1LIBlgSoNdB6lWLd6X
wXK4c2yoV5LmA7StPWkbziZ3q2aH5lJEkYV7hOiE68akgjoVNuOWutR9edqaMTVMUGPptmDNvV+I
AGbaLd9gq/ta2lsUr3owLaxrImlPJaRyYJ/mDIoTrEz2C9S1RB0xSnn3WTNYYbk97EdMoZrMhY0Q
OVJSDqqVwu4fdF8rMcpzcFJQBwZs3KITYcnHMoIsJ0rp6SBJMKLxLjJynsvf6W14Kzv0dG22H+cn
wF7wyqnzmkZ1QuCO4LC+wY4w0Iu+XgnBZovB9AOqm36Pq0lxHmexXfxSYsmJxhA/8SEWmMMFho5B
JYb5P2stiJ4epuDeYI5MSKlrVFpvTRdr1SuuKCssaRJxnEDwMiWMa98be3QttZbV9IQDfI6rLnmL
5Sus6zivhQr8rvu17Dai+0/GHXsOV0WmieBtO/P6fkANluFLyDhZh3vSZ8awywT02pSducTj368b
WghlQZHW/19oJdX14OVnW0jNms66rD5b6wJEPpZZ9jgGj1hFcreiF7M7taLvYGLn6OFpRcEDXGSd
85iNWhcGD73ulzKO2aFob9t4OSv4WJmMjudEvaSrH3Bheq2KeSwarNfWBU+W5HoN2iSHak1tfRBK
UphwbzZgnbJ1UqnspGNrQW3Q+fpxzIjxsGgFTTOFdNui2AEd069BE9vGCSJSvX/wCrNbb1MACNdq
4cqbjJc9TaUaVlcfEKxV1fYutwRYI4kW+B1Ji0xRqAB0S+fCCdzfedVx1mjTVU4Wz5Za6QTm8E7o
DWoW1Ypf+xeKl1P+9UJIXteH9+339rW9rolhDDcxLGKJnb8PJnebnLqVnkgRq3igrH2HaL1stZrr
yVX/tP+Lra4D/o2VPoNmnJ3C5JJcNbAiLFZ5ZrFAIt1ZvzUbdrUM0DY4obMF0mufjnhhkAYsqtGZ
tIJZWVbMaJJtAgQ8WC46AFhTZaUhuFMDjluDIfxQ7L81IolAKV2h3qeNfxOuUVEeUQaUuRmk+fzl
Onls1Zc9q1zbAKWqFqdLpPAhc6ddTaGonk7tdivyP7mFqyI0XKlxcwLAKrLBlA875GH67ISiMKFA
WX0u1is7VthKB95tfcuaQ6slS+ZFR8Eaece2zuHGL+5wuP7u1JWyI20uftIgsIgbRDGzG6BtH/09
3hNTccp/ghBbpy6txB2NBLxnoZ1ylRILfuEwMinsEaB6/DxC8XBzLyiZKmlWP4m5dNfQYzYoswr5
ZqeXOZ8HAfFMkTk2POhWP4UUYJ6ROWCW/1GrhqFGLmN+a161m2s8Wni+SpkURK3ea1oa4Foef7J9
3/r4YTRPkwe8SVqlgITEPyMsJxU/ujJ7zUvKO0qGRrV08daB4Nj1iePJCM0F2BX1/OkhGY3aQSi2
YKU5jqp6lltlgueKD0RJDWgtaZlnou9PWFaShmCJi+a2aS/Cer50HrZeEt+05D+ovdKBaOCfQz8i
AmBzJvvOQu16dY3nlw2tzl30eP0I1lqf4lpuW+WP03Vz7/sjG3w5Zuk9zvnaJ2H5fhQH/Jjo/h+j
cl1UK8O9QBAWMnFjraHck46kurTnObHWhx4UsiwfWMNp7TnNFg8GgakrhOwlewMhPcBmBntbCslw
jzPo7Qkv84RAy60ndCot5iCeN45YjTHsiXK4AGVQwTOu6YbwbgWsB1BpoO5QbarkJF2+V6SQQ8CU
v27fwLOVJ8/8atUYzgjHOWy+hOv6UCR9EqiNHXscCZNaL4mU1/XM2AyF7YFovuUOzkCu5eNTmzd1
FoNRD8I+MT7BRSCFWJIRq9Bb2j6ed6QLFcKUP4umpB6milOK93LIHyM5IjP9YFLK1omeCL3o38PV
ZjqWxuTLeuQSr/dw2oTP1alNorOTDe4UHPEkPLxqRpAry9X/dyc9SJG2BvcnRklDzKUw8H5DyOvM
8eYwiSRll/8Y84r74cgKXFyTVQzm5DYkj3tuiZA5JOEmqToetYCMNxzACSlbd+guGLgczcC5DsOq
nMf8aVt5q+P+teU2o9yl2ZlixCrEij63c14lHKDl1tKqRor6n5FE+tEmWN7EXTF8yAGOZnODOIHu
gjmbsCD6xnuFj7GgyNhrvo4TnY5xuDgdrQtVFQMlaNKirDO00BF+CHAbEwTeV+4bjLFndFRGw+2X
C1OKF+zFNcrtfAtUp98LctBvX89TQzwTBaZVVUH4X3K8+kupltJvHw56toAxWtvs6GCXkYguioCe
BaDYztWrE8m8G2t4zoxC9iQwciVOjefbcwlBmoxUbGpPEUIizOnCoPKDv+G6WWv8AjH3hNyP/T2B
i/z7Z9mDHfCdpBbNziPFJkz4Nce+sVXqdHlXs8b559hVUtz7vXVfsA57GDvl/L+An9a00HpGjPhQ
10zLavMPhQhWLX3cKc+287n4Kkcw4d/VYUNuYaN2vt2a6kKnAXFDI1ieAQ7KPNiJekJJOWScJ7FU
sIqYX4CBmMhiynh3XzEhSVg1fgptAdD6cyskPTIwah4jnlmk9nVQPdj37p1jL6gxgWBprfVvLBkH
R6FNjAYXjXhVSpur7llHnCCRSucM7eD8ZFf5Rbm7awXL0V6k3oZ1zn9TezpzNwduOEV7KkXrdhYP
AOMgA10hP5puDs+fR1QorrK3tuuEBEAE+NzJxqG3rmkISTb+zoxc739KThgSIObqiJkE3+TOwMaR
gKTXzCbtE/sGIBcMKgBf8cR9yX69tmsDWO8VMAVQn5RDefT69sNT+kpOMukYOoscvkYg8S7GRZPC
wYta5BSnHZ4RtkGtf7KiKIVgDez8JtfG293dVbDvuWksJ4gFT1npwSt/awvtlQJHbk5MHBY16cQm
cZ7BMXEVyXSrorikNH4YkwaFZCDeEBvHA+0VJarQ8Y/DKQzBgylmq58AAK116aTawl2uTGproARc
3U817Lm4RHg0cJMjKBiiIvxZlu/SMfzS7zrQU4pynXr6I95m0wBMagy1WhU/wAGuBZzcIex26i8k
n07pM6F+5I3JSnrm3N6QcFkRGyrQ6cVclwB8vXogQlqdPbg0TruewEfcB/nxgRKZPXGh4gm96v5F
0CujiKsmHnGyjLNK6xk2Vm1lycJXSY1Mzgw0oOkRnhCPu6+QNDzdDKBHWo3G2SaRDE2SRVbxFQaE
Abgiq1S+wPJj9vmHj/IZ+y6iEC515wvow5voydZG627iLqxPQY2/DGrV5To43x41ESyHfHvqXvoE
+TlaUYJVUy5MOeTU8Qz6307XqhByLkOACkxEPNWlOq1qe+fd115e3hNg4YTlpk4fwZzP8u/LXCWt
kxTeVOWBBm6Jb5cNy154JZ2KOSVbdfE7axlBkankhZMugwKW8SL91UT0lqs0my4bhgfqeGbEPV1H
g2d6PNrRItbKH571ACC4HX7PEB1oGW/53HNzneH752/YDO5NrzgZ9969rTraSLLu6YYrjXKxeTtR
eaZpNp84p3+Qh5BHgiWs8ljs5tSpkbzSgtXF7e9GK4tdJE85iDrB79y06nO57LO9pFD5XfWf+KpT
aScg+AttnyVAo5/zlAdANeflodR4+8chJTOSwxjA3zosnDxqIkcI3XRlqnaoFyNO/cyEQPThn7Hn
6BwqYgEatZlMJcMbKBCKYneJ8TCfMEkB4WPCl0KFPJvd8DSiIMgBd3LjECQp16DR9XzHWSHvUQ0t
WIQmNjkgTZHmG/xuBLG/FhmsjI9GakI8EVC86qAbMTvmcmRFKHJdq5Ir+fcH1uyo7jpSAMS8ssMm
gEwRnSrIiMIycL25A/1uj1J9LGU5nlFY48ZIs4mEuGrGKSKPsk4sDTwJHnIwhzbx/9sHkwSUki51
uKETGxVtNXx/ac85aBO/Klr7DFXyMSGpBLvHiM9qSGG2qs9gABt83pSGNvjBjgQ/ZdGwQCI6LUi3
pHwYnwXcedKodqOXZts6G2vHjC+zMh/7rpYoSQOs0R+KrCUKSrbtJ6Dqu1TwMmVi6KqKTI/s1Iuc
ifVk2yjjb3IfTy4oq3AntWAXTF9ohZVZCsZyoX6s9PVrWy+K0Zif1VVphFf6p4BMTyiDhKwr9NTW
5NmSqmlx/fN7jYOLTuOebO7uXsnKgq1MzP8wqwxLjlDx3F5+MPSyv+HeVTmGoecjjbuzQUPn3W4s
7/JWpDVaRr+Rw7Eu5f6vMYsDHRcHDTERUgv1tG0ch6jppdIRgTzMTgLAopyMbWI+fOWddlWjyZkU
cVlyjD+oCPHWC+O5I1EbhHwPYyA+PrykkRji/HzsmhbHIc+rG8TmRxh7LQIt8/ssbjNjZ6JMcQao
9+xmkwOaIeUoL2C0l57SoK0x+S/MII0e/yxA+7mGhvZsNMinUsndrWFIeHiHid7LxZYAv7RqRpZF
AxcAxOztOO+M2sHDOaPsPqt818zodTERx5HsdsT6AqOgvCk2iqwvSMnDD58Vk7gJ4HZU3dm0DgEM
bsvYC9CiesdggQLtdk4xfAiajpbInmR4tIOPAowthYwHZEtGhs8vPh+93p7MSdZDdFTCWF+vDnUc
khzyfaOlE6z0KzdqD5Y9M/Z3Bt9mtKyfutkIUQE0CGA3610tNbT68+atAb8TciRaY+66R+c1/wey
jd+iFR9+y3Q9jI24DtCD/hcTkuuurg6CLFtIDAl8RybcZ6qfu2cTuyHwqh1PVipD729V83sD8c+1
tuTsfk+FW2TO+3/jfHvMBkvKH4xxBPz7VYMwD84EFWJGhmt6OKjhPFqxsozP+ofgA+u25vvBJCMd
YGtQ+vgevQZOubS4iO8IluFZGI+XVBTlwhE7s0fl06CSZLeWdxeewX5nJmlAX0BB659LczNMZEGC
piTszV4Ajt+VsoEJ6I3PXIUmZ3mUvW1Q3XMemV6v+raADXdAyppXZNJAmSoAJHSr8RmwCsUSToei
kQBPB6n/F632fXK6erQWHl/7X876MEm9EyR8YcjLyD24/889q8YLCy625PtchwzQOqP9IcrCZZz8
9FMn5wHBtziOSbJVWPjOcJQnux2sdGxTpZdpltKnkohtxjWmsrmLJoGLPlI7ut0yKvTRfntWxF/9
sZuAOHPnOGiauN98rm17e/IPJo4emGjmww74JQCNoGBrrAM9bG3LmQujbQ2mFiC0rurxTOz/Phpw
+CfM//R/S0/9AG9ePfznT8uf31vHMaNVTUyiWoL/iqaHD52lCPmJ5SKFdvziJJB7w5kcsgvkliT1
xSFhcJT0fP9YtT9ZXZOM+lTu7rTkPYhwLnhlZOMW8Z9tmqzINatgogPmGYR6gbRMpLnPyhFwhHtY
Cshgc5R+atxnslDdhkaDbafU2l47QIoq0erPuU1ugbiHyEMaVW+RCoRRlueHpeB+LRdt1sME86FA
hykNIrWl3YkMEEaBbhUV60WnUo6nRfJ4xqpD2NC5pmRk7/Oi1Pvy6iXNZjEF+RkfM+S7zm27mXhc
YNaWRUlXdHTxbrL9Sp0tuIzlcHSAjoEoCyh1aFxPKnUX1k6CB7l2Q7odYuq58YsYq0zebflPHa2Y
iejDKzTcRzKAiZdN33IVFHP3yhjUb5+mIBX6tvMyCogrxhnNVdVR6+T4jb+JXyS9Z5Li6pyAuvmh
bpAhGxg0jLuyHmiMdmW44WhCCM4BRqVTyghgPgL+QqWJeXib3cYxY9g1p2DdS0P6Hg6gXwIeY9St
HjLL02FJnnkTAIWCZCxa5VHg5c6JaZbg7pD4S1PuWQsqtVZCfu7A7W+EDypIx+ZcYc2jP5c5dOA1
OKllrOJxw9jCjA+8NSc5h75mVMXXBrGatX7unVN3EIFmAzEm7lBiUpmw/aoM+hhrjYzycgPV9zON
NrhC5X7h0Nw2lqfaCHapkiTtYKeE9EcUBVYbezGbSxjOmEMn9uN1v1BE5P4+5QM0ou3UllQojnbL
YRnuWo+sA0NRcZQBHyu0sxUpf8YquLtW22DC2iUFsxLNiVjpx0Mu59SLmVPfw9HexLqEHDdrSOJ5
6cQRaILME36QKzPYTnJ4Ccgfacm1wMf5ytkNlBbpUwn8Q9fWxeUL1qFaJBB1sKlTnWb0qO8HwZs6
FrWwIVZRIbLDqv+KiO/FM0umYy4ZciYNUTnJYofjfhbwHECq8IA5l71Rfz77h2VktgVdtVd2Q1hN
xlOuYp6NSfEtKoXSsO1hrddH5GxGNIHuLWmTbKqk5vd0PgvpjOWGNsfnurjQwpwRdgzYJuu8vz04
1bhOKiDqAIEpwZFlgxbCjdE/yIx+cgmjA4VaVXhF3NfsMD5OVnm7J7NpEFuUeuqyWYox5rXNLp+y
Lb4OwvZSWaGB344FJaTYmPAXmpi5t/QAzHoTh54Jv1gXIgAl86hYLb3fHOf4a0MIPSnV/KFqIfGm
ahk8as+ke7a97+LFgY4Omm8kReGjQxrkd5Gz89511gHep5f7gXljt/8ibE7Im/l8mnAgkFvN4Lvg
EtJD2k7UmQ5kytHfyiec9x1DVp7E7zdcGxQPj4OCsOoDTFT+N9/LUpwLPI6W2Sib36EczLNuY+M9
+FSI+5hTgHU/ZonWFCRG2WJzNQdjunF8HI7HsGH+VKCBodz/2OYDJkzB46nnTSgCaYQjyFHolIzb
SmuJ2ioBcHDvSt7gv8V7Qcg+5+M98cwMxxwfEejHvIct0UVUCcVw2bi+D++FYrAEMofHSwgUX1j+
xKszup152dwMM2m3lta7BfYq9Qu1UxSnODrwa2JVIvzzqcdgUwIYSawNqJWnBQ0Sp66+WYba/cdx
HY4afqA0/Tokd2Ond0A3gLbSawuA/mNuQhUwSAo2J9egGSpWld1tDI8+j3AOHH4Du2t8N6K6GJ29
nRCWbT9DZyWJRvPwVSSrPRaCWVc+q5wfeyDj09XiBt7kvDuuzDp95QGuZ9kULIV64KyOvibl1B50
ewnwz7g0Mz8NxsJRo50+Ounbon55ZlXpmEdi5yW4V3Gzys7fpl8LlpjlT6mtRqYVCnTqqfjb/BUp
NC70+bdu60MhbRoPyY/DTq1JW8Ajf9sfKfpRyx/76EH0yToVm7OgtADC2ysradTiNuXcwyx+d1oI
PpDtvbvCmzAEx8K0Do0t6cJwg7gICKhLoZeRg3y+lvzP0OLSf+gp90IdxqrsB10EhAE08B9N+Pxm
OwTKRINPC6gqsqXXpEcMgVOvyMGtqD5991GcfgHPEX62r1ZGNoP/vkA1c20tPCyKXutPqmoE6PnU
waZ+ADXze9E3QIwigAbUGofZzZQr+CaGY5rirPv+UIT7nrLEVmq1NmQqHcr1elzqJEL/Aa7MK9sI
Fwq94nZtYV/zjpxMERMRxXwvnokJvQVQ8vAx5O0Sic4AnhoSnP6CZ35aIViSqactDssxI/WxkToB
C+30TA2Kec1yvEBQkCRdw3RD37NVj7J2M5nByI+ZiscFmPa/pE6I0J4bWsM5nFnqxlsoxCckNh0G
hjqIbIEfQxF8ISdnB8lurD74a0+BI6fCWBcWeeGAmiVyUC2bWAEiNIXazMJCHYS7N9e2ps7F5Ybm
rVV8cealBw+zh95qQ8iakm7VIQOBd3iOWT7zMAUHFTxNLOTJYqEc93jMey88buSgpYI9vVdmYooz
UnJtn1aW8/n901cFfl/A18Wh5D7JNUlXZMKH6NImqiayOS4auVdEF4pDMlp8BjigMNf2doEw0NUY
z+4Y2J08nEYesUCvpMZBmIYfZRRJlKgTZ+Fj0pQJUbMS7eUeua7W3e4+iH5qG5FI0Pc73XCkErzK
7+mFWEQzbzAf2zQ1PfYVXwiYb9g78BVBJfOcTjLg3RRe0rtpW8FillZFyLKRx7mFhMyqdjllFdUy
nhCsV9sTaqezC6XVK5DAK5KNcXGBf0XuBSmC6xapjiYz7m8oGvLPOGAoSCbM9l0LjMdu0OpRUVnF
PJgRiP61jz7Bmoc7HgBEp4MQPVCgZS6e9z+d5nUaZJz5RBI8kR4IKC9UPwk1eT7u75ickGCfbDEo
tQhNWOrl8lcxMzRI0GgwVKU7MyIKf4L26N3s1TjFZyx+lAY0texmAUvXCxfI1dfiWG0CEBrG+OAZ
hIIJxb8fuBaqHsqqkaHqA+lJcHbzxN/pdDWBgd0m5fnOdqY2TyV58X6656JxYemx9nNzrvTUWP5h
w81z1QnKONx4QnkKGe6/W7RSg5zj7R0J71CrNgACwqJ2fkjnE2Wi5scLXbDfzSbAN0KglTGV/R42
Ocb9xbIdTgqJhRHnV9KEL4GzVFsSZky/yMrTGN+W/k+gUUQeB/Utt4pfSrik9PN644Ed+QtsEBG9
47g0wTk3qTwowJ/LfLLEfp9ziK5++dJPv2x9olBCt4+CQpm1VfqjsA2PC6gorzQjNecCwBPauHaS
tSOKO3jgtqDpjXcEE/9XKmOa45Mkk230wax3coTJwTY9MCHZEcksjYxIYwHRPI0msjykMywqpgKz
RpS0CUwhyYA0nldezCCSC3uBM8yqMe0z3cm8n+E3syRvjJ/JUWT9wgx/q7v/Lzdg5Wkcm5T5KwQQ
In+nlGcn8Xx+Y/5QyWKaMagcNaYGuVEa2BqSN26IA1tkRuzoDHujjIj+SxWT8fe2yVWnSlsRQuUE
nQdzULAzPjmyh0VTdaSD4tJaN4nqXL55g2Pn/gtt9DEL/vAruAaVCzT/F9LtBCB5ZOvgCBiZ+DG2
/milyKtJZd2K3HMO6FOFKDlRq82pCBSBg5oL4mCNNtiSzA77eqKp85RwqOVrwhl8vEcTtGkmkLW1
auuD105GeNYU7wTnDdoy3M2/BjkK5w64CPJFQadIxHbo8vl9Xjrtmv9aJEhIwdo4x7cJMIyPtBQu
yNuE5WM3pBi9PdheG0NQUFBXT0cyIlZwHNQBkpmbCWG4bzzzY0yEZd1UO4Yjqwb3S4MPyktQzVbe
RLwNHmXhv/rg2kkW1WP7jVnHSbLjhlXgGG0HFic9x2pGyy5PPWxwIYSG9DsaR0GMylgIKEl7cIu+
7U9DluumuoyDeBFjsbY5T/0ASQ0wbmX7ZrlOtGrdGfcDXJLPbUTjtC7mLGg920LtGZZtX/OrqHm6
/7JCi7edv/1B7znh5y1PNcpKkwMkmj1RjpXP+5SnoLYFZFU2RwiMGz/6c27BlmyhUoXFDPitJE6M
2gagVwOC6o5vIMP80a7qwSvnp9vsF2uc2YJ3u2p1AHTtC+/uh9NOZXUvIGcw3tpnXnWdbJ4Rxp6t
ShoVP46bf8SYutuq7+hXc/Tn1IYQphcgSz3EOrMx+ppBfBSsgGlCpp6LCoWVH+NvCP43U/lO63yt
P9fCA2LydL6SIkChrQoRllzWkSaPd5ANR+qmXze7m2y2+juOK29idBvqe18tjB2Zl+8Uou42qlFJ
uoaEsGJSDKl0YO+gNQ7grQgaZgo0J3QtrpOw5zLOEuV1gyohmq1D4880KMmzQE9M9ZQw2CMy5tuS
hkqSLhK1ihUSspgi/GU223eIuP8dWBbVv8JJGvBOLqFqPgXR6SgQu0TmwNigReDNWgMaO9ie6Lwq
WgdOSP/mPglMO8XP/yyycRelDxzipkllcgsO3RHRGspipIOThskQfr65M7Tfa7OXTpGEzZbligMf
zCMryhUzfcZYwfvCZi6du+Uhvs4AzSIocYO4B/Sy4vK27dZW39gQuEoHXz9b5j4rYlSnYVATNc/V
Agsi6KgKuudYi1a93b9ZM1ayIahHxM5qq+eEjQnJ+Ip/y1N/rTyf9UpscMD1L2UuE3mTlfLekavZ
+YhBydHCGjDlVoMYhju0FMRFAmCBVvg0hDHL/HMHdQjKM0hxXDS0QKlRxOcZw2F0/i83RBnMg3rY
yVzmGHb+akQsmfByyFrgGdioUDUy16AnfZSGTCjC1qoNJjBbLwzwRbGbq6Eo2jDDiNRBuaGuzho7
VTOQnQ+7hwkbGhyevHMXO1cpiTugeAzUHQbCRmLLdXq85FGOo3VQeDqjbhGv8LJs/bHY7r/3/Cyj
K4Gu+3u9pEFxN9czVGpUBCFwOZOxum15noQptUe0BBSAbis7oOFMuDhVhk8BiQwypdb2bbKz6CzG
zW6r8EF3ISrtB+Il8tA7pdCDbmysS4Ud9LUYlFVugD/RxlHpTZD7cSiyS6VF8mIalo6KfK+VU5bc
Ptim11UPWWPtNm535Azx/OCuWGUv7RIyhw/deodHdvjJGnvJbx5u7QLp3Xm/iHnkBohrTkwGVydp
6leHANvzdO8NfpWXUeNANvexwRd2gSE16TmbbjuC0Oe9eTuaXEPGmBdgUrid/L+Y3XZquIYexzH8
PSoITzp0bPCTvKvZnJ/I1dqm/N2H1hldV6X8hm22zFeDDvBvKFHyb+GV/cLBxstvQtR6scdHdu7Z
Io938YivQnEDHX5J7RnOsvoSO2YhueEVsEo3K3XAfT+kHGgw/zR8y8/MCXhyYtK8DPMuN9wQWpgK
0wBAiPiGRqfauhkYG0LTxKgNbPQQslSoWo5gSsqFxgTmjxaTZMnp8MxeVAEwFH0KoryTxfnv2agF
EGoBn2DBdCfU4pXGfpRtjKPZUyk7GO1Hyo9vsNVfWQQaxYjBXLSOoGu4cPuA7XA0doimpR/dxlc/
Gu5t5JXObGZXLn1MnpIhIrZ4eEnVrdYDyUQRH6zKB+GCd/H0VJm2NBNHnEXnx+iaSRNcsY7CIKMZ
6Ndm1IE7ipPK2NkUYTLAwY+B0L9+PCN8fUotQYTnnqCaddsqnXWqAY+BsoXIVHkO+Yg3/Q75wCoW
cbTkw3e2aczVav4IbFp0bd1G8OjW+wgy/F4B/a/bMk4oJ0a9rhp/HkF+JMZizaNUmo6BAbBg29OH
ULBexWuzXaAPNdOvZMPfxZnxy75gtUu0jKDU12LzAakG9jIck2LYKOve5ebVqYI+xak3CNZdZhxk
ddM/PU2oNdEuUaRdOArkfHzeEzSemKzOd7UnD7wwTTd2FhOlFWaz46q9atRVVU/q1yrR/V4iH1rW
O2P5FFuPRaiGPSOPWiywR06wqt/8yI7MOZxo6xksCuZmnpbMSvPDDm09+fr+dk+96O6mu8JZicOp
fr8PsXJkfPrzPdg2j1bbey0qun9NVTKxVAAROov+mN6VWTgW35AAfLRLFGDcoekIPAvahTao/wzR
L2tIlw3GQVSK2xNWlyN3lL1R5M9QRGfeIDXNaigQ9ANhtCSNAUzVCgwR4/xMomyp9vYUgjcR9Et9
5N1NZJcJfFJEarz3heO1/UwDzO+4NuOxnZR2iXefVkmlcAir7SjJC1Zjddcva63JyqrFj0ZJiOhZ
+lirzTQ4TB363MOnSqoOhUBvzYduUbBj/+RgDtwjJPZ5tY2ittWsxAxiCrELc/97VFC2NjevHIMB
3FC3XH5ATiTLQwt2gwyxNN50EDyhVtVqzkXTIQn+/aOJ+D/wCcEeTtU4Jj+K8z0eam4pf3ziBjSg
mkSA+9Oj2DOSe9v8MtdTGP7T1c6kD1Ud5Q91NrNs1sLXsT4qxMCdsQcvi2DkqP5Hqol8i0diEN40
0BzicLtH7VaZobM05ks++8hIR5i9QOPXWrsqLN4aHfNS2pBQGrrXRgfYEBheqimK9oaMR1RVxT8P
kYEq9oT5a7RguTAs3prqt9PeTdcPA7AlzmoVYcPZ9DmjK0gKTvC3Zml4/4LZFBcvH/VmxMbvRgMq
R566VnF6Lwb0oOqO8gD14I0TxEVV96AeHjrY8cfMOrhC0X6hAgeHzs3digaCFpiAVgRjX/lprq4M
fnJOL1uJQz7DYpStbn7E3kdW4GIvuyCQjds90We/RWALa2FUpmPLNPr+0WNeM8Ln99lBz4nfitZQ
l+ai0rfg88gKjfNilCjTANatR5AEwGdQExm2kA2+N3mWI8rIOhvHkQ15PizxfWyz0yz4+ww3wfpb
mgnEYXeHCbZUiR188rrLiutt5MOoj+qwm63fNV2pRZzZTaolbn55aapsZLgJ5A6THVKHTJQ6xbZN
Fz4NU5V9oOj+3QjSZv50h0NsBOb+3q7/TjjP9fEGWH9pzs9wMPFOl0xbCDCA7ZkDJiMQS+70fJSI
/rOFk9yjDo7u+5n6/KnO9JW+BoShHgTbsAYoJ1rhOBsAMXxYRQpSx1ulbWoorEdHobplQGtCYzm9
h7YD24MISpb030rZPEZgicxX77xLxViO1X3fKgHm7K4/qFW0vy7BlmtomQ/gaftz+uVYGvEMhBHy
HzTJptMPxfMTpWiYtLGHxAXOq2BtFNL0XRcKZLk4/JDf/x4i2GcsBQsNsE5Sx0iTA6B8OT2ztjTX
D8x+xEiSAxRlWEqsfy+97L96u+Kp/wrR/EmIlgnfzujMOM5jNPXVIW73XSZKDOPfNJ2ZN+xjkkjP
WCpD44wD99fe0p9ayqty7NB6E695Lis5mmnQf2imLs9t/W04Q/Qs1K00lJfP/gwEdbNbOLexN5bW
AaaXAwVB+iFHIPEz23zN59WRMPhbX683ZcTlnCPIzlVsszC47X5RTpTzrm9aSIOa5XhuaPvuqbMm
FSbl4WO6mPsE0VMBhgeeL1ReNC5QAYVIILZuIlqBWxl0kSNA+OXSCW6Z0uxhi5/4s0o0DUWovYDQ
Ng+Fr7jBk4N27vWKA3zm7v0tKogWxY1y9aU/nBwMC2uNfhQorUDv6D/yHCbAafSgK29xo8g1hkIS
eRZtBy4YfBzINp89x1jR+3/sJBFmEBcrcF75OoZw2b/QX/+RrP8paXXUlNAERgsHXJe2vzl60kNL
NJZnAM3MDvuwt8OSrC1WZ01MBjM7wu6Id0m7WeZ4KteEzXjpWfc/o7ucXSN0NGQWh01XmGEbIquK
t/Wtx6CTB3oEQd9GSzlgjx5cpiSLp8rF8L9+VYwvpnxKyUamUJn1PJdcpeuNetOAW0n/uqNA0aOG
mmTk++Y4hW2dpXuHe2NXntMWzmmmWUUJ28hT8LVTBU3MkXYeQyc/blsXpI27PA/7wIkt8FfA1VGY
GCCXVTGiPUAefucmerGswn2A2TfJY+/6Vzu7fipXHhGpaMRTdrPOMwU5zXRfHeHlCK95wZ+O0UC1
3Vv078uCkNdbV4g81LM59qZgLbK7AyDjxf7DRV4XmijZgtBR6zh2xuBr5V6auUhpEOETfUwW/pam
UuybWK3MIjI7EMgoXjo4lmrs25XvLrxXUFbE6sDSDg/rKhS6sGCrr3sF26MiDfWcvsgwdiFTM+LU
zHg/ch61jkATytVEKHD1OpUjfjhlCCwHh6tqwAbHRQ3evLf0hx3AqwiFHO1wiXvw7zK1Y25WKMC7
hbebXkEc7gdAQt7+caMqVwwRJVtjTKOGFsR4Xmdk6i1QkIYiYEqKviJbotyNT0c4IsBu+zPKCsbR
TSPuINcqfyrCLgFZOMb/jR64DkfA6anbJxQyOYQbxJhj4y9tVUuMFLDlY8Kfh0AG7J7JXZHrVIyO
CeSZoItUBITNirCyvOB7na+hZk+AxhwacpP81afoKZVxSmBQl2g9b+QV8XZ2JF9gz7iXe/BQa2qf
Uis+TssUJ7sRMjC90s7xmC+gPAS/2RNmi0X8bE9rMoM0qmxPIv6bjgCWIHi8u7yEZjDBnBfpgBaF
Weht/aCKDfOcw2jWZomawNpxO5+naYLp1SukXanFpMzIOHtSKmhz3FyQxgPHBqwvk6DMAXevrSef
R7LlsS+wcXyluu9P/7GLzp0LCI7N4boBKyNwOGWePSMQ+Z7brCo5mBFkVksbP5yOGeicTYvvdWE5
OFQ799jJ+qvIFwS/QM8OIUOwMWSsSuejwKzFjZ3LjF+KVSG4eAfIHeofIEvkvLOKoltamh8Pq7fd
jTgVJlqvK6epOKp1QZU/fRooNkVmeoRyXFP1LQ86e8/oq47AG9ZXR8uvbNmmyffd0gKjf5gBJUka
7K5IuXximEzmxJW22Lvdqv7H3XSq6CU+GAnIa4Q2VAtYcupPbas5/tCBI/C4h3INhJDAm5fUEV0K
no4ThTigs4lfDVBKHZ6yieaCBSQgj1i8XO67dlm2Ia7j/w57/GMIqmZwo2N3M6GcPryAXobvgeqF
Kd+pI4jwl7OD1zAZUd0V/G74WtZwagvYhGv0qj7ru2CebpdMdM9KVde6N/UMQfOoTAabXR6ZYbi1
drXzSiPZ1RykScLGa44pT/WyUfxhrzk3+oxcwrHcZiP3Rp6ktarRBauMMNheqmUVpdQren5K74yz
12Jz6EesFCC5vrNvrvVHQk35t51qLcr0CMLs9ciNk+0St9APtGW1V0CwGyg7/AjmTKdPT+Us/iCF
xKOlSEM5OvXwMi1FOdTgqsPKWBuIkL8lUjrnxU6eFzoCzQ9NHgv+04XIdfhBoeQgVnNw1LT7E21K
facwGU2LpT1cKNJw/LBjSWb/8bQA0QLL+RxxTxicEm8OCHGxMmRYkDj70IEiLOy/X6N2u4rpEnYj
WOorO3AAkjOOjhgc446LD+Q6f8RSfxa2BSquJmgbhz9k9v3gvY81NYKy5K+wr5TgKK7/xijnIN9g
lMnZ2m5U6AJldyl+NndwVcVl8KxaWnokgKsZlOGx/5ejYnIvC0Mc21Kkn/bjtR224a2OHBH5KHSt
y0Qc2PtlxTNZDSxP0Y8zmGudfRlEOjVEW6DCxJvWDVDqxuwXsDoqyEB7BDKhxEw6Lgrs22eoWC4G
539xeRdJcuqgQEXl8nHxxiiDsoxUbiI0TTWkZkkx6d3cYme0s1R5M/sXucCc4bF6AvlV6Ng3B/XO
qWhmtjpusjCY7WTZ5GYMEI6ufp6hT7loZDfpD1ugL6qXyp1a883X2kkfWoVa4Rqn26GIq0mJzcA0
WLwmzLppSWsL62RpIa0mwv8Bg/Gjd8Rsxjh6v4oc1QN9FhVyctzxdI7LJLklaUzuokHbZPANa/Td
28ZFRweD3G0roT0vG+JyA5KLQ1E6Iih6LeZ8i5Ss6OcQSZkdiNkyOy7xC2UGAuFuFBdAXUHw3mXv
2RUBKie4Ne+DhNMv+Rinqdv2Gce49G3+ZuuPsjNJdQLTRYvgHvtLN4il+tR7gcE5r6hcBuwcmBnU
Ser6hR6gM4ZI+YEEHxoAAj3wD75yqcY5DhEA8Bi9Q/FVbuM6krfeQe0qvA2i75rOlZyZxiv48f+f
5c5DWhLwaVp5L3UfLRrFumO26ePgV+qfzFI7jFUJUOj54s464oUhNm3d28YvA0UuUTvVpJssEhbw
l8ohadntqm4asyLkgMsRO0z4XDNSDUm/Z01DusTAHQarXQ+z0qjivwxJPebmUrTsVnvRvp+WXnBf
r8BcSS7w238hZEwkpL4Y+sdsm7E/9lznRsQT+QEuewOFdlU7bpwAcy4Z1GL243H3txuA4V0QkIeC
nGrNHBCH/Lwnb2/29Bex30eFf2ZVS17RDGyIWx0ELLpIScyek+/100WGEX4RO8oEnsRjFwpXmiiU
aB/o3FshR062drzqMwmQeW6wzUS50beKF8fkD9E3opZa+w2lGY8XMQTV3RQFckAWdp36qBK9hEEf
oi0fvBXzNw9Dv9rHYuSqLJrBfR8FxtssbrFsRbnpd6PVoJzkZKVkr4aOQ8/KIwtFYZ2Ewzi1UeKo
ZQkVfY7dBUkp0wtWl7v3pe0tGinIsbRC+wdtxrpEV9fzCDuhtGhZqyMYd7EDWF2yAyF4czYklGGh
vHgRiX34NZFj5/c987+YVi6D7ifiE3fo3UhboCd4Afo5R3GYSA6ZzVFZTUKXgAGtZox9hk2eDauf
W/eaChIpNtSlXGexRmj+7k1CTH3XqPkMjRZ8mIgsQ9AdZ+nOaOVfvF/TKo/Xz5S4Nb+Kl6Og/W5J
+4oMbZ1/CeHvnB4jb0vcRdr3yiKyjDirLMR5IByVFTw5nGbNSMBRMr1TipOgAeB5AECIlQ0lDHXu
jl7SQFAToXbOIj/qGi1W7rlb9lXqAl5DfR/pzq6TrC24h+aTCY/jVnO5k6VcijBNijR1yYqpRNvS
Z37WZOE2RBXFcFmUPxk8xVB8qjR/Zo851PYKjw0EuwhmHfgLbbetELzfrqPyNHoDsn3gaXthMU6H
sarH0OilwS8y3PjjoqNQk4HZRfMdJPGqa35IsCkYZU8KJSAl7LoukcXZ+tJmxkGt8f7KSuFj+erv
vOhHqNKu8nP+cGnYvxdmXwfkTv6lMpQQPPPJvIVWtAaUOwXpftgkSpNHIXDGmi9t4I5iJ1UPrODV
ajonztnt4bD2lCeRvFV6XqsTcWk7H512uzjHaNm7+NVXgoh7FMljkRbJl7Ki4vtktLR+wzwgXSe7
OOWUhFGADeP9YpVRRbk9kOfti2ZgozIAAf0MoHCv00jsPAp4NWEugN9J5eLETglm+F5XcZSHP1Js
8dplynkAlYOIeqmPSXtJeh3sCtIFhKDlpoGvMVljkjZxnowG1CDh2ctEfdeBk6SMXTe082GkU7Ql
t9LPw+o/uCZenz4Js94XpZgqftQW/cH0koJh/LI3VOH6cl4/5HSWiaZ/x4qWqoTaddRiEoth1ftE
4jz9hXrBRzqh/V4YytPkxLm7zXvuvouy2a2F5NX5D9emmt/iAxeroyxgw1/e5iYlCJCFvebUj8VE
goC3oaUKnD7tUFtK3n5fMeo1zR/smgqDZy9Ti0rDbX0o/z+2hD74DZY+ZxLJSzpRSQoP2avuEedV
d3PNoxe+EvmNch6BQjjg7hMmOibWjItjtng8AA8HlO136l54kh0hbxbbPI9WPb/NZbexr+4+mGMZ
PdeOI1QFUkKYLew+Tin2agWeF3keha/hzNs3D+ISnlbnwYinAtRVv4///xhEht8bY370HVIdB9tC
muLFSOSZPS7FFmt+7sgFoOBV560eaRRnLue+K8GfXdg3sFR4CW1Ci5GnLoUOeYS6avDU6+LnHCMk
7gQj2N07pI83PmLMasL+jgT+TPlg1mWrZsbicL8aD7tMxSDSho11SWnm16/XzDn78pBLz7RhCjKY
g5bw2Aa9PfPOVSBuUpiEY57kCBC4A9QxP11LKli3yKUR5MqsdH00p7oNCeNydwgMuXgW+NNsqCP6
JPoV11UeCxes/yZcNmeCDpIv9eECfe0wjL71c0uGvs0y1VOtnbCNsO9mZQEA0R9IZ4TmhFAqGR6Q
5EdRaZUBXR1poSGi25K+EGTTsbh7CTkHI2d3+v0gYqw7gZkjMvqtCezil0jjdx3ypp8/JOmFLqWm
Tg2gCR18B91QIrj+y5uL+sMmcWSYUowQT6+DPRkBpQZlyUmxrIxgI6F3FRPmw3Tad7I4Fdr3AHBe
07AjFY/PYsepjEse/KIUbkM8LS5ZF2EXAFYpSlLKT+VMh0P4mipO7hh4e0KTyygKT7KM0foOG373
PNmlFD+9lentVf76WLxTVQK7eavtEeQHTbhXyDjF7dkWv4/qpFC0cOz9m9F99ULX9ylGEK7xr/Qh
CN0wVt2FwTl1szrYvxYZzTu+mDiX7RaTkluqHBlzQj8DZk2/nXKZunB/p5rTaKI5u7cHFvgGuVTL
mMqOoUre1MmcxFHdviYx6c77tJvnefZoSbkIkv3AkeZ5aNqcBGwJ4LGIL/KqWAJ0inWKZQsYeHM3
+9TJA8kctoX/p2lML+SpwZYX1T76qJwrVY6URk9bNn1Lo7i6iTH/XzGXUPsH3aYXEAvf5tHdcBJ0
Q9ckgCUYQPjZfGOLGUqqVoQRU6e254ZGq9zfaUqTnJDTVAw+vOa8mgoCQxP3EMX1vi5HdPP70UfU
GeiXho0At9q70tG/ZAU9Y92zL3eAlrxb2/sJ+CnQacigcpburnNhtOqRM7uBOuDhW9tNu3TSL1rG
pJ+3avbd8XWpkoA0u9EDRsC/VhiUizfdoG2RjNyT3fm0CQA/uZSe2+qkij94dcoDu3ApFnCibiM0
eXYEnq2jodTIH8pQIitTSFdzEKNE2ll2Wu+LMUVpOCzt191U9dejJSXt78AxH+SSNrZZywTvEHJJ
3qL7uA29hOF4ROf3qLQn4lcMAwu8ZMCS/aZTTPF6qv29hjFdrMqxOcQmwY3G0RSliVE+mtI4RwEE
q99G0x/MXI4LEmlLveXF/+77z1/e1RUUsgsSJb4o+W0q4HC598FBu/f3pB5ezkM4feUrTSvqj11j
gWIR/v54FFq8Yp0MQGI9YxH8pEGpjvecq23cB1IQ87c4adPf9hVVsf8lCuhxsZZ+1Yry1c3s0Hml
8A7bQ4s3k1ZUbJ8i6Q0UaDg3d+S2tEslm+WIrlUua3+H0HRlSxrsLUjjWWyRcIkrNm0SrzxmH27Q
AkB/FfP+gll5YNGscgqIw5sfkGgOuxDP1gHuprV8sMKtbxeHuCym2zLZvIH3MmA/hVF/GomgfwXU
hDtWY5Y28RzCklV8dZdoHWKP8xQMJW8np1KoLznO0zcAIZA1WGtwRHFvS2zSLCF5f1QqSZ8sXSvH
ZRo7C3Dps0Pa+J1QWyZz+BOWX323DWWge+HSE6Ua7cvz4FSVPFomHFGWIfDBsXM0A/dHNc/O8sEI
k1CxbDoJfDVPgTRUB9PNy7YaD+dxbmyOBPblRw7sC6JZYYZPjzwhmdzlEjIGQLQh7mCn5h8FAtRN
5d1oZ6LfXb9Me/0SBJ4lhGcs7JCozFForv2sYxZtDoYkyBh/0QeDJMZvSGjT50lPzCKc0PXZBE+x
dvAr0dI34nAYsxoUEocR/9QdIHElzDjIN99hRmc0E6uwE1ZUmQExirTAOfzgFGelYVEpZAp3NI+n
1sbzwarKKGEKEAhGWyI41e2h2lMI3LYeXwnsKGDvE2CkNDRA27Sjr6VLy6BmFIGrvLwvzcCzykZN
e0nLDgmV+nfrTsAxM0et31+KMKuxWc1hc8I9e8+EWdmbE3t5SywavCh03QTz+jrrly9GtHeBvJfM
Zobv7RW984leO+ycg2ddsiucCLA0PiSbDe98gQ6+mo7G0TObxq1Gj633N7DVElS1mfs+nvOxHhfv
SianQ7Yntdcx1LdPamUntRS//rbEMYbiN6lHt4DjzQNiv2+E5wVBe4/kLTW35+HqAz7zJTkFnXLq
h7z/aKVQlEnomL4Ywo04iCXfTsmbCEoYx1dKnIrieDIZemAmbC8JpoMQ2QI8Zj0u1DWSnV302XkF
HG7pwdmUy2Wnm7e9wp5+eDPBCnSw1U/FPXpgYTgSDHzwqdB7DHYJxrmszqTxxRubrOyC3196/bqB
baICYokUMHI6FgR3SsTd5NnIe28p2uDXTNpg+ofDI2nNMxFii9kkD10aOGoaiQ+mLb6Xk6InShqx
7zswXQkwhCX31ho4Pvm4usvrFCOIlVin0i0AtklO5FKqYiz6Z/s6gco9Np3Ux2W8Tnm1w8B5Spj1
FRmdrsUhgFXYfqr7dcKmcvin41zxUjcEDU3diXjEnIS9qcbYEwWYrZ8sWoKWKeoKrPu6f9wJwe6Y
jT8TumFlC6f+tJ7qlI2PNdsTGKOA3/TB31fyLBpziOj3evYMOv7+xf/sXWhKn4ghzIKrzSIwEAvo
mTjtUXO+d/h5wjrxoDXkKRmqshX5nsN9KAfw8i+YhwBVq00Sxmr8FySqPvxKLuxxjPVAo8PM7Sw/
FoQ9guyMInVE+ir80NnLe4YYul221PakY4GTAgfZqnj58VbryimJESt6s5L26wGlBrKZBtaaifT/
76t82LaHjPFZRzJzvxW3Acq5d5lvmHoLCziatwlcADqd3Zm8kQDcxqW7R0ejck+uCr13S5Vbbw+p
paDFlZytpU82v3Fj1396OO63rztdyINavqW2Q0ig4ZqcBOz615iilR40hJNIMuV395UdIVfXoIH8
DwRgCu314axjZpYiOU9I7u7txuYmnqaWEgATj2KIKLU6T+n+NBOYGhomJyBQnHbWh8GD6xFAh424
uYQv39CRRjwepyA1Zy5vRjZhmIwJ+JpC1aJ1pTjqo5QtOMzOSII8HPF8aTK7cioyxZueXljVmlhd
aG2ECt+p0GcLWZ4t1uszkFNnFMrkWhFfd52yrPw5KDbieoJC+UDeiHd8kZSo1HGMfv2wuy7/Bq9m
aEheIKZ3cy73CDM0HUhigtBBwMgpeAmqRoJKGhsHa72EC6lsJ4JWAohAHqYuy1Ns5D5L/uyLJBA2
ZwTWSN6yaW88x+nnMh9lX/MLnZxbQk6WfFhxuAmdXZuBTv8UnSxf6eL9fOxTpGsG2mv/FDBQW1Xq
cjGNWrGKzwi0I6m882ymAZK68hRUrgpxZxyqm0DDhZTpLVIoB0WkLuBPhj1P6uIVjQQAevvt17wB
+DnABRMkiW05B2oOPBBotZLWYMIXWz7StAcElv5V2Vp7qSnb6mIeeju/Z5q+NTn77Ze22/b6qiIE
h1dE7W+yrzabXcptR/wlaamcN8jQXUGWA1NixmlR4bPlGBf0m/Njrj0SoOQqpzD6XV/GS/dL8E2/
uJmCAyr776+SvmHWii503a0zo8TT+Rx6srqqueJHN8HD6A8ceNpBcCxQmxXlQjtmuGy2uiK30h+P
qe9kDTQ7tjO3TJInltR0OHDosj5aSSPNw6JUHnoSEWcNiRIKYXVxc/2422vYh3CcfWZ30vX/6Y/D
NyNUBnF5nJgRotmfSgxb8FbJcyeWWKSUB35XaViheqiT1ZMauitmX1aIEJrqrd7OxaC/EoTb6yKe
acXa4xORf25dC1ZZwZA3zeGEjto/505hRaZ1KdaoKtUulz/lQr52VA+FeeSJhyEsELzJaHEvnoRh
ZHchsvyptyuIEU+lzRGpcmJJkYqnXfRbOVWE0JAL19YTCwUNlQAdz4lbJ7EaiyFabT1+emM+4a9K
+m7bGKQYaDGSCTUif83NAufoXZvGb5MUJ/NhUEMWonaG8ShDW+O7OwB9eyYhQYdsDXKw4wkM2PnH
fskNMYVaUqiNt9YLBlanDztfD+j45hEVgORFEYKFAdPdBVdioTeowY3QITDtJDsT9UqBW957q7Cp
TXIgrfdndua2vWGhd/QFkF11VJVhv9CBbHZBBxIhGyN1KnhKQEuvhGJi2ig5ov4M/mjyhtlUlEHA
XUL7bZ2n/mAqxjfnYedVugX/qDBXPaqQlBgBL1X2XYgx1dIRIrnjIw3C6lK44pcG5bKaqAHC3EV/
KBuCXu5Etg0Liwk5rhR8Gb3agNeNyXdC1Lu/ZDHdad7Hkc/BYHOm7dkhVJ7b5Zyn9oTjedsbLtpj
V7CyfYxX8R8bQXnTfuqRS/BMOAF4U/eZxDtdGwF9QymYesrAnp1SB7EixnNP0h0TsH4GiLK5u601
D39TFJB51yPRXU9FkO5pZ0ailpcBuR4DzwgEpvEJxoo5ga+qamstDZHZBp9ZGcyCnrlwuPI2UwUF
n32h05oDNiMTvtsVIwN3jtUnvyqMQ42nvO+ykJNLuFsoKGl5jBWSVQKkyFnu/vL1Y2+E5W2LHLFi
gKCro3DEoC4aNCtPsKqUTpNpdn/sVHzz7+DD/OsAmEjLJcfd7kYURmwkEKDtK2CIzGkujJqytssP
HYJwDyIurxornf/HblzvIX2DnsqUIe0JJcOUzgIMxqYGQHQHXh4BupTJrIfyv7QrsUYOdCYUjugH
PuG8J3HV6yT78/uadxlViJJA6sbOkqJSJWYF0Gz32iluIqWpR2lxZZwFHseccQmgkHi7Cv+4JB2l
KkRLCbvaa83pV0AcTN9kuJjfyxxFILGj4bicj9y+fYfTMG+Fv05RcSd1wUeGJaCoou54HW7q3KWC
I104tkVP4cG4UnZ4KqInGL9ZAT0Y+ekYzql00CczLruJz4QWBXZqauhvOMBkI5LKtrajw9TCIKTw
q+20jkV9RGn8diLsw1cbequSiYz36AoCQnxD2YsjDfk/aKS4o5PB24f3Cl0io6KVpjnL6K8+w3zr
1rj3Og+BxNu8H9GpHIJ6K1uZB5nprnu5hWGWGwpFrazFeN683bctbHR24IwzY9RSA8V5gNj3qKgQ
KECpdbmsoFIsKBvG6YhZTovDE3GPWMn2brUAqrQAJZNrc+CZykOS9WAC4IHsiclIpRgsW2vdE3ff
JgTint9FUNWc1qKmA7pb7dwGw9dl9Xw3yiQYsCzfuoBV5VLmpV5u/wEXyU6FoEu7dem4mIJyghjK
orMb3gh6+S1+gAWtKFE1M1K+rZRPaltV+EqEjIQoUmM4TkYwY1MS010Dvmet0642TMh7t6AFzBgC
W6O+Ji4yJt/TvUeeVv5/6VlCHYSPv/1WGxpljFxafiJSqv1MTua/ExwHZffXCKup7Ad82etEJfGS
Aai1lOeT8ZmDcBTYvHNbJtD4tMiWHpuDJhU0QVL65mYWfboZ7mDL8vmUJ+T89I/tu1ha2MB1aw83
C3YSBIm1Gt8mgwLvrttfL0sw6aY72w4UxuOEDWut5xUCCBw3mNBq4yw1HPqJzHD5DPUeGojLcMpq
H2H1pvl7+5Xvdle4xn8q6rctT8VUtflMDU9O1v0Xe0PeBQs9jNbHFTEYyooxhiYfao8sOD6m+qR/
TXtvCRavvAiFX7Twe3z/NRjYoOvsaJ0/dOCSmLBVoPYmSivqXeRm8oMgPy6EpM3dF7wDidD9RO67
VHkptYhJCB3l6Ya4S8kqCNITwGfeHoNSjHS7eRWzdl9SDWz+JiB4IRBBPC1Nq0dyJEBdEwTdhboE
444HbSQVUPD/s6OkDS4aNbGHKP2/GVAI8dB2SekD18mzpLir/R7TeFBpjD0LVZJb0NNiKonZP4cG
yEadN2M3D9W+EQ5B7OTn0iFQ9/ufokcGhAGoLDOJuPG+r+MrRxmWl070oUWsKGA0yhVpeB87WptF
pwcxYCXP+wdV95TBkDfPY8bVVbueDPPn6xN0f3h53ONexJRCDwKGO7TDGMs/5W1pXjxDpUvKJTBh
2kGfKJKa1EiR66VYUzLjTv2E34J5e4c0bg9b0iRD0IWatZAdaXp/z38NHXB8PokRFoaDzBHt8Nak
59HMH7oSFPsUW6XGCq4tuHI2g8K70sLnMNrw0DhegEkEIro6ScPWza8CmotiVan4GcpKNGBZt8Uk
+m7LIHk1aRffta+SXGCAM3PIN7Ae/y8XMaTGv93eJ+OQdhklFwUa2rtgUXRS34cdZhPyG2RNNn3R
sB8Gas5vMrmoGAF58pQvS2xZbXaNguHk3uJVExhlnx7JoZ/Nuyr7yF7BqbPzCnfOO+MsRzYYMoQd
hpsO9vz70NlkgIW7otHbqMEhIHmzkBnJsR2jUMe9cXQIIXwTXaxhBnc90zV78FjjCcKYrGeK0dZ2
N27bmRgnowpXzAM174iVn1lcR1vijyU9JPcexeTmue+bvc3UiU7QDShN/CuUddYrYiR6pxqzqDlP
fEFuG7VXsCLesmqvE7AieK6Ps99zTFexKqrLzdAFxuTeJwljbK6fpM5zFMVPHNE5A+eHyK0y89lL
uhKy5OsNQcbkJ8lykBXTW8F5cRKLoi4diX4+5tdJ8K9nhYbGzlhrHFDkLFpy5QVHKr3D5BSP0rPF
wDSgwV7tV7p+R1kPpMTX7wxhuj4EyS3AMQNuvMidJiT/KW9z3vmxtVCS/J0nyWbZ5GPQqy2fSEIT
2fy3dOXi3lO8l0JWeUpZAMZ1E+3izfGq59aB+sM7UvdoHu8FkZ1t0DZ7e6s4eQyyh/YOnxD7ppJD
xER1dBVeG0N/5ymn22tAWJYqDeedja8ofrDsOuf/UTFvCJM9qnYg20dEV2e4tgMSlaxgnBIAMy4V
kO01HnY0MGFMSxsvGViTcq6uj0y6lBQIgmh0byJwydBA5s1wJ36SihlYJSdcvzqxhRUp5StneomD
xb9asmsZmIw6hfIyE3M1zCvGYsbGbeQIJ+49aLjCo9mvXXlvS0bGbUliFKVxBRupHvXSDWlOyz85
F3RmJSWo3c9dLPOFfa6YXRuECSldseKcDzDp3i3g1J2ga1dTtIgmhUgf0LctNrFyF66C5bzhBMLW
mFoFdbDQNH5kLq9WQuv06OnPZNbomtj11pAQJgGy1PSl4SZ9/KFXZrAN7/3XHxqF4+d9W5sYQ9J0
Q2hpkf2/SIEDdROlfpuCmgagwKDM0UpBPUdNyKyl5yPsFLH/yx7MW3sW6rqVAmA6ZVaGWHA6+xwv
dS2LSA6DtPsROwpPNzBLCn66NeqrTDbZAWl5oyU3G/rxGmPODUINOveXJGG4QKy8/yr+pGqTKvpL
IQEXO9bvgc8PoXYtplpF+TpivlNtGX3eIjZEWyoe/uB3uCOnFDDv94FN1jHpyqRaaYDfrRs/sHnm
HdC95UJICLpZ7S1CBgzF/h3dTgSEmtyXtSNbnEbCxBx9vNO6aL9LGUhji9a83T41ME7V7sdhPrhx
XBS7G5h4KYNIw20/DcroMQfoqpy6o70PnBD3srwgh9APHPcCOKHK4SbnIyCnVMPukDaz3dHquD5R
Ydw99xds5IlN521Da7OQqwAq0SFpqEuqVohuquPk1ZBALnusoqvBxkZel7Xz8We3gvNTjn9wwnS8
2J2eseN5qqGKhN0LGBNRRDtCvoxKKaG15Ki1Z2h5RcwoawR9KKzr39vi80vmUyL6bmGy9QhrrgBY
rgGW9kDlTV+kM6uS12w4Vbf247HtA91cFbI8Lw4t9729aliDtxImFOBiEAftoLw3XC3PMUg+ROhk
9lzMZNEdWRfPku0lWwoyR0RUegfKxR/gOykWJbs0DPjWz9/oCiSTweC0huFj1ie2/Cb0mr8pZz9v
rrC8LJU+6LiJ/XmuQyPtj+1VHj8Ms0vOBM8F2ZkJPOwYLGMpjabP2MwXm7xzYwj1PDGxCIkDMij0
BDtNF4Gwi3Z2SpzN5b+z1KkR9y+tW13fXm6d0oLLEJ8cl/yVDBDhOBHkpUFoqwJYDI31Fpmwua/U
PknlAGxSwpsfN9KG7PAuJTZGkmG7u/DK86/ubsh0NovDFwP32y89ZthGQe4MglhaGwEQ0Qc6jjds
6rz0BtkNcFG+TLREG82MNLGdwg4xqjaUUIh/pfxyxQdxG0+LVaYDFbEqyx43e+N7HJXLUTIqOhge
4U+nFetcCXWxVrGCwJtmY8ippjKMaRf1GiWDIy1y3iT7/WpM/07uR99y8M7RZibhHjnQpKVzpfKA
IzCmVky+Ve4doOLdbKVxHCGzjpc7KKwDas/0VrsAy7MhZOUES3Nkt9+EP89+ddFIVCRUAi6DNXD1
XQgrfsfEEFTjWx6Eoh84CwKybft+igKKm0lI0+kfIH+hXhHqDbOYm8PMTx0SOFdRde/SoMUu81id
Q+quyGzeca+WxSBJ8vg0YmczdrrBC725MNQeRRWE7QSvHsvsn+F/y9dtwumhSgD69KiXMnT9paPS
FhTNShmWHjpxyztyOwPt4y96OVsU2qlYKeV7INAKlf4JD5nz4MQ8gVrm7YXLo6K1K0DEWmVKVy97
d2xtBo2RwQnTUMGEiQ01+P4g86X2rTN9ItgyaKq9X3rva8OE3OXVifBHle+0glXEw93WWqGjMCx3
afp3vJsmjGpgK7sBsJcotT0wj5XtfgdLLT6THjJ/LRh10wTAHLGJMuloGLxcZngeMAh5VItnVWYW
ip3T+fWFnqtCx2ABGr3PyEarX12TnZMe915N+SRQ0fD2m2JeUayu4pyrpKsFSdqgTWTQGQ/ebfm7
VU8NAHAPtpqYdPpCAY2Yjxsep5mvk4ugMjNE9GxQNh7YX+YE2f3oRPW0A0QuldY7zzx+2fb28Iu4
CffnCiJPlEOGjSfoBj2m1DpfLUirk/bfLiiuO+A35BgulYGejtS28BVhaw1DMDtnOXbyrRCaIsCD
oSbl1RGBRAKN4co9NuwBcdff8ngXlkqVNH+vA50DAF/+WWA9PGv1EuK7g3j5LyAshyd7ECuFVID0
730qQWgi645FpwNex+NU+DTlOvhSnIoTYofiTh61i2MxD5LZ0RDiUW8J9QbHklLD5e6+EClBujVa
pWLW/Nig3yWnN8mT6Ywscu8YrqO63JHJHLkIG2ii+PD6dqqLKYrqoxEbeN1p4gC0vM/Sexo/NvSc
V5BEwxgz7RGGKo5DakUquS2a9cFGGuoUUeIEDIS03gzg+4WipJd7ZPb+q3CNwTTTxdgtlXBMsg6F
NeEHDjXKsz3q5Z8QCeY/bRm1sxcVsRfq/bigqvVMAMRG8P+VQT0TEcIpVg1qJ1tNCdmaKa5IEC6+
3ntjjCl5KKXfx0xxRBIXnBtu9SXkiAQkXnbag2xRvdb8xFrat9+xclCoRGw5lqpNh0XAlzmE1Jny
7Yaoj+5vNE9wR+qEJqJbk8WRuqEOFSeQlOu56cPEqCoOfQlLadvo1Bqoycih4vrCS/rhJDx+w54b
dts0+nzdsR7s5LHpwG9veqHeOfqb3UMsfO6vc7GcTpqZIlBF+wJB6UoR5hbS/OTTyQjFMGToCKyl
H+wlOc4S8TujoJHC4UJX6HfhLW6gWO9b5zIKbjmX8dP7DHNscPqFuNwzuUR31BP6YHLD3qfHaXjM
5ADx/QzQ5DrLCV8MJ2boxicOyJ37gIEcrV6N2e1Id4tyyVigQuKfUqdskQelEa64FKsxYYbMqY/v
gvwhcD/JAYIlZ1LC5bGyQ/KmEJ353Q+AiwUBFfHsPfBD4BPvv3JgIG9dhHLHZJHicf1gvvG/i406
UR6T16pwI9Sjz0PfVbSnUPEl5eAMjGdn8dHxNaiQthswxkVKeMVjXif4rhISgU8gILbVWqTObkaZ
QRRRl2z3wkP6GyADk5dmO06bBowbZiGYEY7mpWIcrSYvij+ni3ChKpxBoGb/ZApCyLXbyNyDlM63
T7v8cfc1VhMTgOED+zZ20BOgYCkvYQhmlv8ASewfA8pDJITV7La9LQ+0XhZ/K3/u0vc1QxaXd14V
lLk8vZ5MyFzt1sXm96mmCVvtCF+uBcYKlClHfd1TLh7KXzhzThzh6suG9BSrsQOV/zy3+CjGu8CY
igkg1qjIXFD1S4ABPqE2vvtpZUrRuk89XPqdCjJrDxaOTr8Ao0jM/vATpbctFaOhNio7BpBvrkHP
glo1K60WW6SL8fWgML60yEUP9PgS1+FZso+U8C9vPU6/fRsM6Q3Ye3OdXIUgeK5QcJuMirRcxu7C
BxAPGb5RV8rSE7ZJLeRTp/MD9wQcp1i+zKROsz63T7LwwIVd0TuYZ4tzBf4yhQ3FH3G7OGvTrotz
TWtxLDPMT0FuRlzYmbIJ2m/sdx036PCUZ7Ay3XIhfdQtPghYAhLhm8N9ak6TMz3qpSYhw7hDphmt
n+b48V/JBgb+zeEUwErWnUEoCRJlHTQuw/i5BB5eVwGVA5asI15ZaPlU0kbc7D9w6v7DEdUIbtg8
CZTl0Q2plJ0ggR/ynOQL5jFcCf1i7lteBzsQ3hfCTvHILM2QLYB8kX1hpa/Y71eMtSMWFFKV8Sgq
EmerDUPoxE3wgvADc284gTgNpzsJN3LXoK/VSwRKobxaPbEMM52EYy1kAGsb/+FhnTQ6RGv+mq5/
7+wflfe9cq1m4TvDSfGzDhnbB38kjE+Gv5V73BAVhstRlqVULjbG++s3+DoCUNA7d+/4nwC2Le8/
J0cuiHc7KN5TmeLY0uTQr4bJjo8E7EU2nLKBAB6jVGFvWYk7EO9+U5XsH32qJ9MeRMjkTclGJdbU
Cn4BQQQiz8cYyWZy6fEAt/S23nJUs/JU3N2fLgn227hCbCrl0i4TuXtb2sGk7jOg+ErDwHCuBOf6
FtNw4lueb6h+uOFsZ6THnmMJVniTy6Sv00V9FffZx4RCSmrzZym0fIqXh5wg86Z11nlu+yPB5Z+m
w6+A8OP92rDBSw6cnGCAkcJh7dU51TO+f7JpIewyVf9uzvWl4k4lEagYCGifthjMCVCsYhTbDw6s
ZriaFIxwXudbYDGIxI+U0FmnszUWUDsdiEMfbqG2oKeR0zsidS+HiN/6nyuMrUJSmh6arVOcpqBQ
rFuMYxqOy6loxjLEL2av6a3D08/RU5RKHlNj7U2QXRYSQU6gyJdD9X1cxxBlSsj2xYdYq/fI8Jy0
LysC0ozWMaYFD/MaAHZVworTq6+jLPxt59ZiRbxy5lq8+VE0VsA39nBQEq1jJPOn/BxYVk4tH4mK
PhCIB+qSj13yZgGlUVKakDvrCrRjvjSl2dk22oGMdK9ZuiI0bAGvJ7o6IOVr07I6eZ+PP3Y2+ql3
K7k5anF52REum/z9EAsVRFE5jLV4rexPFj4QYjCCHBjHArtYiUPj7nRACK2vonCisQRDl5A46rv+
qmELNtLXkXD7hoy7scfEvb1rziWPcp8nuFsLhGuY1eNHtgJBRxPPLj/EQ0OJ8n/SOXUp4tSpJLSC
6Ty2trlJu4AFQsuBnJwYR1V/lTgONoKHMCehrzX+AGQRnqIY//BbhYNDeDCEADV9dy5N/SuzNKSo
plTpimenYSovKT7dE6kg6fFfNqSL/3slfYlvl3F32INU2sEjcvcL6R/v1UOrHfvUfJ3s2cUrdOhu
ByEWixRAD5juuQEivbTG1C/pFTfhsjkcjnxuLOoQPHFrqdxa2HmCn5tcWzMYqh2bEGy15/9rWQCw
8cHhejbQuSlcbqg4Wg7WeqNT1DIrfS0INfIhqN1rEeaEMRkcP2+QbAzYkB0KDuoRx/sIZH5Du2Un
Lak3gvMnzXsuICiwV4QBct2ofoXPkOwq4rmgxIdAPDPF9vt8iTJoJp0s6blmGdRdlPEEPPWYopCX
oWUiZWMgTJGmRpUwJ9339G/E1gsCA/eBiba2GIj1hXx419DrsO3J6PnauFLzLc5NdywJzLW+RvVL
u46VXQuwMOwjMvSYY+K6VePu9uexOEdlPGVip0hAHv+5jrpxv//XMPGTTbLNczTep8juhnYQtxQD
nPEzsdL8zMQ6V8PSapqyfTKYVHIZGmwtVPqGIuJ/v+CXaaRp2MWTziAmnp4xcp2zc+TXCcp2Sim3
mIU5EP90u520jTpZFd9JeeEMIijtfbmyVjOjZ0/m1keVTPqfXF6ccGQT6RqVImNTmgdruwDqEQYK
TXV2QGRhMU9GDXHuOa8WJdXeDJoWWjvY2eVpAvR9f5/+25HSiCWjLyy2O2FDIQWNFfh5Cgdl2nbp
p6ZGUwCsKoif+ZTZX9Ux9Y5puD9Gn3uipjhvwClwyBUFyvO+PR3IWi2BmNYe8o+AhICkYjIB4gdG
9t8fBCPNfu+EamqTNqQj+1ris5Bw+/O5h/W8GlBSR16jas8e/R3F2A5iMAif4L13WUwZ2Zu8Hg2A
Xr0J2ZtRuPOZtlmqI8BKA2LZw6CKd00/S8ZMdrKJGBBxmIZ3qEvUg4EHg0Liksfs8l9N4M0gl3Dg
mfKN9Ku53IP70uxNYFulgkcczmor/LLtWnCuAbXQHqWkmhZGgey2BnzsOYPrj80JnJoVKF4yag+L
TwUhg98b+iPCvX3wLquO1GDyjdA/MbhDF/I5F6RRrCat3EgtoCg+Lq4Y9xgDYxKieh7QIIfvIlex
Fv4zvB7+aupZBxN9nXNaes5J2Xn57IxJKQRVhNdEOtvVaK4ysmRUpfOqYI64G+tg4Po5WY+RiIkj
fLHfTQaJbkRQGPR82+8T2NGYEFqMlNhDlLq20ODvvSdu9n0ZJ8Td0n8y+3ho9TmNvKL7Hn+QRh6a
5CgRWMBw43A9JYN3CGBnpkdzCvHW6VRtZZounyVGVoINQJBFo8iiQxqEi1/gPX7wCy8BxfNwFIq5
8sj8NY+a9eVh3opdRbqBdJUmD2wpdU3WD4lFTnSkXAc1lEWl8AsBaRE0T/95SLU2tOdHbilgTz/E
2KZM7+IJkXFUhOuKBGckdp9+CQTpl/DYwoIVcp1h5SQTl7Pc4k9Qk/lCkWr4JRx2GbaWG5cr23AI
/8yTSw4aSnEX2OQycwEJB+IZNCGhgr8JqrjXZxCc3mtyTilmYBVFnZ5JiNZd68yT4LdAWEOeM9jP
KmP+Z9H0k1uU86sT1mH+1zzFVOb67nHzF9+nLH3MN0pm+J9/KUrzj8EHUe/tsOFM8Usd6q9iHPON
1Y1xV7LDq1uaHiftERMdX0jLYmNtgwwy2qMO3yXyt/U5Cb8HwxaW490a69b9XJ3lcCoTf9T1v3Aq
4FC3yRoOl9Djhdu2V51WgSR48ATk9hSKxYE0vEjN5mkU30N3Rx/4LxLjKudKSkg1LkjaxGl647DL
WsS8DgOvOHOIXonm7huNhohsrQBSQnAc1XbIbjL53b9EsrkJZ5L1/mdpiLST2Rrr+nIEY71v7FNc
NiKYPp+xAcRcc4qQYUgC5KPES/Ga7WOCjqsT2oAmImenjEh/TyLV4E7cmzbTAT19NRTzRqpx8GUz
CUFkouEOgPW6YJHfljOauU9gjtQpiPSprQ6uaIFK6JSBx3gad2eAMTdLor2x454kbuELruQTxxHV
35131LZyeixxqkUeYNpJk1vP2X2OGBdJUsdOrzUl4/C4l6kkpVxcE966nEbJElMKOyPq4vIESY8M
XQ1luDblK1xyes4a2vWYb3TSHsvP5rM9GUC0Z59ehu6E15zZ68G9prbW7mw0tBeuyJh8EMgHhUHy
HSPY00CNYOy2rpnrJhyhqt8UbdYMybiAd/sGIpDFmoJs8b83fPvZJn1EOlorCJnWlX6Y+QguNErY
o7ofocNrjT5C35yoV+C2idrxFlmS9ZV21AzsO1CFoShP1gG5XerCgodvUQZdmb4YnZrL0A8LIqgm
eMn2Dabulp0h6HZDZajtrANjx+hPuJyCSsSHvbq9DESMzUQDMOLxUOcNGexvu3CYhuvSaxdIamjH
bKMQ7LA5rN+TrdTwfJq4TFPj6/8rfUw7yCCeK/vJx2ftKPgCqzJnxX7EOzSgkbzJGifHnga7VYob
Y5OoDs3R8ZK6P+1tomVmGslXcozRmWeVUA1/UM/Z0udUadGQBdLjK3VS52dkp2YA5WkPqg/qMf6W
AlkA01aMzA+xEjnShEXeSk9bk+uHEkkb/Mt5a9DBE75PHVxOGVNVzKf0rKfpXn4NeiElp47WSuBV
KTTKwuOjechK6gOqmITEm1ZARHkwLpXh6yhxDcjxu/wuMYFaZvJSQ0TFvJaj/p557e7yELjy/k9A
zg1d/Ns2QZG+FENle0+frc/ieRe3TVzxZcK2UGoOpq7/48d83+nBFstlh2nmUKGJVp2LYap3vTbh
RCe5qdfftqM8lWcUpsWL1IbSELuswNVFDrL+AsMbmxzLeKkRZczuf7FhOo8DkBTsSzlSi7C0Rh2E
jd+mVD7NfKXHGIjR9ulhLXHkDCSHK0JYvqw2Eo2FnT9IiZxaTfacdShhKhfe4E3FxXR5+TYeBMzW
JlFs+R4w2MFC0n4dmztimsm0MqK3ll0QNkhwHCpVLhqNMTsaZ230haejnXxUvIIf2c/Rxu0jn8Re
Iw68jXh2yvTGefKhG7zzc0/JnDw80iUq4wLpbBFPtosUPTIF7cLmFO/GLOoMNcOp+NHh99eN5OB+
Hc9VJEQXHGL/L4IhJLQeebECYS2ZmwAtEYf8MA6NGoK8KaBdfpwvFsoRjbb5H6q+uhBRxrMaViM/
iQ2gjqQ36H1y8G3MJOSLEZEVi5peyfGvC6/DeEjfwsrYYJHEnY4KnuUJctQurDDUquw4/EGkwCr9
fU9jYcWUQj+k0ccD08SAW5K9Nnuf+GkmfXMx9PSbHgcI9v5j1IHUl3lGHR6JBqYI1kj2H3l9pUc6
umP+lxMzdupM8hiveQQf1nqVu7eHCf9YxOaTH2Z5Ea/36NfpHtHrwRUgp6+OOmNMPz14rlB24MfD
jCsbUVycdFcFfZUZY71n49WLz/6ZkFlLMBR/M1LqfOVBLcpWZGGNGidn6b1DqsPnKh9cJ/LhzkXT
WXhl+tErhDqy4StiOCHZU1P0xn7MB2waN0PouIj+tIaE1Scwk2Szj32PmV09ONm/DSdLvKLr4wrg
Nj7qjTnFPR6qr4ApXZLz5q77qnwV8hx6cF/Rq3iMdMJyCuaiu7hRnmt++HqA3inTyGCmgug+SZE/
H4wx56EWU44sJirK28aj9axBfsBGXji7WlMXfYx6n81rjl5Ykwc6/szpwoSB8mBLOAypYOKc2DSN
m99bVdYDzBWk3RP4aAYamaNjaiqNJ5OKUi2qfhJtcgdq0fBQ0A3Atd2HIDhAZRey+X+ba6yGUS+6
8g+08IaFRe412dY1MQkezq5KZktpp9/0G1BA3Gwi7DRe2CWaCWpdlzLuvVDqoc/7QkDJ894F8Jwc
OPegwWzDYs7EiaMow8pRZDdho4+fEyjeTge6IMyaCBkPFu0URG+FVskumWmmtm21J00HG9o9/sg2
/Pz/dSnBz37/QK57ZZ+LhpKHrztKpsW+Li6H8/J3+p2SHcGqY+my2GOAsfbAOFDTSut2z+B0O/ge
8HQDZRjhPizG5Z2CR8DcM3cH+T9IzBtSaal7DI+6uucEI66ldJqFjULiU8HZWBmh4750vs5dtsgR
Vvlkhv02Csq9jtkdXWlXOGg9opibKu3+8OE1D7yKwFQLl4KnyLePEuQ2/PQtb4SRxXe1Dym5KX5r
NRROvFJHHFJmTwfwdc8ZN9kBkfmdzDhLGU79M1wVjc6q5lAnnUCCqKHayDoKUApwXbE9nWyTWoC7
Yef70wudwFz5iJX9xdEnejiwJ6WN1wRlokP9sbo4uZfl8FVAIEJrQAdalka2C3KrCNSnHg013yIZ
Y0U8HNzW9uWGLdy2mXtkqDjT8iq5NoW5pMjuue7NwMnobEVBv8GdtYcGQfTFLl9E7SCIPS90ovdZ
T8ecuf64PNCZhhj2CeRfqFF6+r09PYWXr5rnQzo7/wPst5nG3DhZ+koeSowaT3HPyi9So9J+hY7q
he17z4w7AwydGGITMYHmsDY/VaJsnTBhRob3CqIhTzZ5MKDpaLOK6RJCZi04PnBfVQ6b3xmY1Oih
9TPSg8fsq89yPydAi+gKO5+Jfm/DSVFk5ae5NrhqiT4mWlwdfqED/DVuz3fUFHloLQvY07bqUw1D
SshFpcu9HYx3Da3eNcPl7Md9f/vL2gsHluRxjGAy0+Kd8FaOkPUP8w0nmWSjLybbAvU0ncnbNvDe
xIUM/FvXc+UyGDx/M/3hmJt2FftGNlyrNPeqpaIaxUqplGecWkysS4yxod9jSecQqhdSCLUqrQsH
dybFsHmI1iWYN3LNQFKKRqPbPfRtmVBsMh9JUsgKCtCoFpJgx6uqQz3VR2v0MirRttAIbtDTj/b9
MGiY9uTucwa7G+HP0wdYckgOpfRKSauvsz4a5leYnTMqMnSoGpCLw9m2x+o6pVbhDLLKq7+elMHm
AF5EvvtZ8AaSXnTBtRYJiDOny2TImzFi9cnjxVP7V16hkAMXW2bHa7myvmNk7PpFJMkm4Sp7/9/7
9u7ZxvfnlkLEV2LH49omZ0umit/vUqKzOIHE0lS2hN6PEbU/cThzkhU8BxGk54E0/k4c+0tY2kbB
LK36G0em6Dss7O3UJ7QVGgvpGpPGUgpirq784xZYKXTDsF+MP1brxDAmUf6JqoYh7+e+JdpfwN38
TH1zsNPWn2aP8ftRCZbVLu0B9W5ijv7zPZUxKWJz9UkvAv+6/vhJKH8Ov3AY2YFNCWppTN33FTOE
M8GSNHM8zM+QFVPMikHYE5ftQvHlNUY5G1Y1D6btnm2Gnlx1mwvaAHSgQxQ46I7LYaFBObqvBiAd
Kavr3ZElsas+iDpyYNott+JnIdDD1KZDKV9QaL9LlBQ56ygyTTPtpIvGYeMikaRcTiph8lM85F4x
oBOAJxse5qGn4Q9rLaILTHMgRNjrnape9fQxlADR1Sod7Yyz3cbfTIxum+MKnLQ13amc/Ckp3+0B
B5jk6G3T8p7ZT0/KKCxGF9P4ghiM9bst5Na8iX4vD9SndaG1+vVjH0tSmgZYHxXprYXsbls3HGdu
H78HBZed7gj23P6KzZ5WKMVmoYZ+ucDpd+nKporstZcAdENqU16TdnKFe7kF05+n5jMYI+9rDP+o
9YjAZ/kjG4uDZyCxJ4SdozIgQcCDDx8Rwl4vokNAqwjF9cWScJNqt7hfqF6MV48DQc9RHnJDCxl3
dYfeTIiBeFyqnrBUbltdxLrn4RXjS6HuP6LfjR/xdepOH+uwRocqbVq2MKvXYaHkrPS2/4DbNea3
ZIh/M5oNnI24VesPZLF3S8Lwlgpk/tsxMIu+07zBlX2FeOrZp+rrbo9LN8ATIcp7U8FUMvxFOB66
WDIN3f2CSHdRcrYx5wiM8zkupMvCpql2LIUUitu7YB325ZZrfazqZuqshD47QACGZSull3BtTYjM
mRPIwBkfIP+b+Tv0xhoBnfE4K98+E+obnMzugKUd4qTdFN4rW3moq4mm95PxuIC8XjTgUsHKgRuq
OhRnjK2GZ7CkQiLv8LFqeu/IxRETNWNdk+KwGPAXmVIuijQwEd1ZyZIcSHoG8SAmYukxadWydm0S
X3so5tUuMqBgn9mnSg7ofQx95IADbHovoa9CLJz6IOK2aADHxf/GfCrL26UzUp3AMnvB5oO6WEcy
ozyGjyag86biRKXQoxGWbKWMAkjveupuoUAVskYvjx1qcGBXNcyi7q9N4vgJ5WxiukK8QqddPFu0
p4Rq/IjhK2+AXUmCMiiHD8/i9GRwLdkXJLGkn1mxO8dJyAcTztmsemExZeA96IVYAvYfwZXXR2ID
gemiCZUwGlCW49B2IYLIuN/TkbD4srULhGbb6GMmSSE2XKFe3KCAjK82t+fP2qxxoRvd6/mpQwyF
aLxZ3qR2Zwu5enHWuUJtozdZnPfS9m2uHlkHBM5/QeUGnjgHl6Pi/kzRm8oCqoQdbwbmuapb6HhW
OfHAo5E7vA/iqbRLpdrWNiUFblNan+IcNt4Ho0IVXAvzY+L1ObGZQhJ7YfCtgZ7agR28crrBgNl5
iw3PDDes1hbNNqPvDELqF7zXpWWaYfuieTMwi/79RTEqDNiAqNbAs0ufh8qD5pG8MCRQ43Es76nb
B0xHQ24kHU5Rvy6nIHVO7y+Z+ZZMz6kvYIArGcngl1AtfBvQK3VgQabtA27Mt2Js2VO15BGQr44k
GGzpS9uiGFrJe34oRJ5Kp6u4WsNaBu6jAAOg81UKn/7WOoxNx9/dIyrh55wkCpZE8m54Z1A9kCcR
TKZfoFcCyMVoFmcFH6q7x6gj5uVmKyQ+yQmF7y5YsDNw7TcHW1DIez2ittKsZR9wxADBYxS0us0I
vKvNMlKitEDa7FDUKdRFsHS7KkJ6PCQRRAHH/9i3lALDLotwHc+OZ9yEJg65PHxr1TSmtyl2/Q8P
mlo/EKwD1AgNE/FIePjmpyoTgcU+XnpWRdCiTKDY9zfvuWaI6TBav/u3CvmBHv191cOKQJj0gdc4
59F5g4ARylCaelKyJn1sAe0inq2b3Tqhsc7FdNz3SxOVgJlDnvSL+RHsGCb21UW6MAYJZ222S5Hn
ffR1zXzDZfXsF090zMjNr5Ym2VGK1D2cE8GyNOGhDvT+NubeOPjyu0erHTO2O2zlMIoJEu0fpQlR
boWqxJzT2eYktH6hc2JP+EdojUiHmyMNeSw9RUgAiqH7uA0r5KzrVkRT8aFYJbuZakvic85HJ7KD
oAvmX8m9wM5A/zwxZPUdmUwwkDhfI2ZAnjlHA3wZvP38vYd9paWANEroHXXKe8GnAgp9Tw3xnkvD
CKEz/SQnMnwa8/smSMCsc5zAkqGuHqmDch5/E7tFUxceMgfSjY26BnKZtb/d8sE9UQFcP8kDBc8U
4h6MsxTSPSqL64WtozcFR7CDxyDWpmhkikBRmLAWaERaYvyNq84+HuejPFArbLZO6JZksUWjrelV
FyoP4ThAOehMO2BCM8ODuCIUOcS/vuGq6hOZ+Ex9lYu+JQ18PeXtbYXvsNi/ojJdd4vO4P+cN68S
BmKu/GCn+5lwCSX3gg68yLi/FLdzbadGqGx14yJcNRgEovJ9lsLQvcMG/LAv49bQPMhpcrQn3JL9
CFOb98Fm/6qDATML1lJYT9TgdzuM1g1PP6yveOj9BOeJIsGobVrOr2Liqtn7acjZdr7jAfTBE4J3
cO/H1o1aqTzAYLoW2Z2XHQimcI8tHRtO5+w/VudR2Sxx7ja1Qde/k4J7lsVTJM5OmqNJqks5LKLq
qjjTlXb58vRsmKHVeYhZGLI+pw8GtbSqYjzp26vY+bn16ZrGjRxUjygF0dBK1JpNBYPyBp80T3UM
8evJUDZ1fjC2QjSV1qtPmMhjTrziN5EeRumaly26RhlRXN7+xKca93B8+HpuDv9DFPDvcjdZbAz1
wbQVhjwOo8ay7piNEWmmqf3i7nw1Fp7MhtVdMEqFeZzK3mq25D0op/LBO7Qi8U9J7oWtxInN/BkZ
kaW8nbiXNfwnwTrUlvRt0C80l/iqRUKEXJgZwxY92C4jC7/UlD9nnlkkXOze2+hW8gOBA/VhfX8Y
XOn5lYtBw01QV/wWNfkc5jHCZTcJ88PFNxf412Sm52wI2cRqGiDAYuDptGNm81cq8FL25LdWhcdX
lJZMH1J2r1fGf2HHPqGLd5NTY6j8GGuXUp/nYi2y9zczeKTsYG3E+232ExBduUBHr9KYVmfXW/EY
yE0CmYLN7LHi69pO1IcugdUAmqdTXC38vXwUnxaAy4H4cdZBKQFmKRDFil7k90iQza1R1+I2I1yE
PwWpf56QdgnwLxzr59Wzob/ssGZv8AWcUl4lMK0c+6mIfSzjyXPXBSC/3tDCfER16BpTbKzuZQX8
hsRrfRHLtwoivZEDnnx6WugCC59xAH2DKIOjz9em9hgYPOivHIVIc+Jx90Ow1FxMU1TzPZVeFeu2
c2KBvry6wFz5JuHMvlJnioWg7is41rMvNtiZtBna1wtD3H67WNB/yDdK91oUqRK+xkdTUCshdt3I
yLnLSZjFxhMncAGqKCVijT1886vxMmet94l/D48tjxL8kEYoF1xvqoF+ecSr2y2zlBaC7aEx1kA6
P4A0BbcIyp8BQ6oSt1lGbK949QrAmbWkr73IJjEoDN/M/dxaL8vZej6pzra1cuIHfMWrunB3rb53
W7u5CpUwQes2NUTMIWi7ZauYMt7YR6FtmUaStcjPi8x/MRc9YmEXesMzSy15HxwLdWkb5jUtbFLY
oMKtbckkSIskDD5rTHGvMYf7qzuemknES6HRerXaUWq2V0JQI54iGWU5fH2y77FwV9d4ANP8KFxt
gDtbCs9FteupSJpgRSla7UhktQRUCoVNchY0t8VJFuX2D8mdVSft/OZn69cv/s/zCQExNYCLDEgm
7kjXBxiEKt3lR60tilWriui/Cz7GRkFq3X4cP8Ze+4zKG1ySaJ7pTcLZR1TospaU8MoCwzyybfBT
nf5aIwqb4kKEI+f8Cvngp2i87Ve3dd8aqHePabGgnFiCjJ8xYq2LgI4qD0aNQ9b41qOj876qBNA1
n+gcw5ozj7oAJ/yED4BRB2kU89SmG/PsiPFt5u+jaNuCl0wRuYzz0hcoJF3FrL15BRHtI01CjqMN
3QJCtSU0bZL5Mg9eBsVc/KAW/8A3SLIjRv1C+XKzXT8bp6VJjUwqrsvgsiXMmCwlxR0LqpsYkZlW
RritKVIwlVZ6lrvbfJCGFhetpgIuhdDrixMgXrKlfBbOpu3Sgsp462BvPTRT9mJqa0eYKex3lSul
KDA63c4qaWmW7slKTtSfZ3uITKHpnMYfn/RvxmBPvlKY8R2sHE/j2SNI4FLJ6mV1FgOVSdWmVCvI
nGe7knobDftMhReb49FfgVOSzNfpgY6GafpiZU8ShhoPqUiQTiEzT40SodGB8D1sFS0iyxmH22w+
8b8L0M6ESBTaRCk23jrSh/UOLQLADypBadHUiVs9MyhTyPXFdHs1spm8M7sAk3uf37D/XCgbHbdQ
ATiwjVJ5RAIYLkF2Y5fZhPbfwR0zZkfUgTbB3qVC5hV8w9X98T13mFl8a80ONewvyuqOFgAUEatN
XgaibI8XipK+rxddhMOYUCLAvR74rbrS9Y7dttKFKoJeArycNrb2UYu7x9jubUf2c0gLA/imv3S1
Sk0GEfCbbdBBmQ8G+6b352i++DiAVtaIW4cG4LC+W0ceBYrAlqYQbTaCL8ocPLMsqUou01A0765K
s4sS3N9vM2+izzrVkKpniTuDaB/pEF0d8K1xDURGmkdP4y5JpK6rt5HOTfRJ7IKSxwES4juf43h+
hjB6cwt+TChDHnODNT0SaNZ1Bfkur9UWcffV8CdQpPmUU7AhtHwWigP8IVvHB8nqFbTQbYQ30JS6
dvZDjd3V+vCGfoHa/SaxNdXl8VicDxv2o60aTmEJ1TQvJH2ZOEEh8/ub4p2MuGbBu3UAe4UGNaaE
7NV2kC6QKbj7qskYYHrrpE8mWtbarOBNVF2VYGN11CrpWyRl5/HoCVKGkS9rIlwJEe8wm852/lXf
qnHfUChywxuy1IWtf6bh6LYhpbb82Xx1EL09mBZDzFB8h7+ukSQbe4lexbQOkV7rQnEU7wezx02l
lkjr3h0p509h+oqwI9yZq/yk1nxEQTZIFXQL//rvdYL5gHkB8940Dxof3Tg75ArO23MiN+5d6LR+
Ke6Q6OGOKWuJoGs1zhKckWd28DHRi5eO7UdhhBKI8/CtH3LLfkC7H+K1OHDLFSZm+iMoDSTsSErT
eolKjBRs5RE4BpngVbI6Hb1Je58AuQWsde3GYC06byAlTjfgOekZgdQv8mg0j+eFApS7TJlVm1Gz
TDHb9iu9YBvep8i4Hhu7p/KAnPOda1gCszYTAYFTP9H9AXtMIQ70trtsTz6UzbgfQAhVyMoglEex
hleIj/z+SFOMKLr4sOgxmOBS0lsrcgvb5jiksZSXP0t71EYf6S92n0zVK6WBzBnzTV8Deq041RZQ
p2juO3EYFVPZ/Er+lpgmFNwNEap7fubPAc1cKbYibuooaNHE+ujrKExs0hgvbqXL+qE/rXqSR4vF
5GgRVzXij3LbrDD6VPHvKwuhAfvIh4DdKokHvL8XDtddmzRTe6oGqv+oQ7jD2VtZG2FZiyOAa9Tk
I8m1GOSbaTS7+rusZ8GzlPc9USahQJplcIvlagY6FUMQLLO0BSM03zekGCI409wFtTHcgcJBj/K6
dJSes0caCv6sDVa7FvtpkRlodFyw2tXNvv7P2xrWDTy9XODxnlrV9ecorM6+TYH0O+CHxkVi11of
/2UhQF8rACWyq/+ynhDnbXA5O9uiNZ7JAMgb7GaZTZzupzOqZ0B8odlgq003l3W7hVNmyOfd+81l
QPhh6J5Cf/D2QV6OUE+cOWUpLFxoUc/FJCPwHcntDrkbwHrfUa0AHAeWdJcTAbjDdfz/WXkwZOPR
g7iaxIq0JKRioszxHBhLzdIy6bnWrTAMb9xu0mWdNNdoZ5HzW2hL5oHYRb4YS0tNdqP7jICimOdo
tCce/QIPC+hyij0z5Yd4eM5IeGLvScqmNwrVPfUD7jB8GP16FQoyWDhPH2L5MPzEJValzuczDNQD
734n3fndf1LjdwC9+7y+0PX3LqgC/4jHTcdRFtIegCOh0OxSWmqT7F2Fjm9JYz4JDCv5QTw6iNyt
lrb50ftw8Ici2/jTg5uQnGbFqUMUvjsQarLt2nzZkchA+lkOPsiuiJSEVMbYXFW/tpKw90JuRaLZ
RZeibunLdaFwu3FDP19jozXyVXr2nxzcW8U3f6gGFQjfpMpLry4MoIfXkgwGX6iI8LnCm7BNAbk9
VA0Emsvu8K8o5Fh5zQmlMw0Cu3IxWRM4+unExCp9+Gwe91iu/8z4XDelGLDEmggZ3ukfSaZ5n3Px
FaVo9/AAKeW9FzuAhVjKsXuqBWQva9LNh2Cka/dPaOn4X1A26A/0+J1J5mszv/77kXLey3ZmBfj/
QG3XaBbTrzyUpFgLQn5JkAb2Rh2tk4RcFPpkiLwEHnZQiy+pO3ZjibWC+acb2Q6HgospfvqiGOuZ
I7w9fwL6atWJr7VE9QUdcUZr+NnXuiG5mhJL5QjcxhnfMy/53X5sM9X5IvgDfyJYjRtYLtHTxDSt
e/zxQVkQCWlfSkXfLQT8Sv+SDw0fLhp1+4AFk8ylyK1QNacrKSyTt3yBrmFN84FbIrKRnJqtvKGp
5mZYfCSALlfwql3KLB5YhDrLMLcto7JqreTcZ5KRhCb5I0Ehw9QrwktSNdSDs3nFZaHihQL2Q+q3
apdtXy+F1wDFLwGCkL3sM4XCkZ8FLBqa+39/whGTwTHjDAuIk93IAXsyR297GOkusfI4Vwpg7d/P
TUNiHW7ibEVG698PpuYe3Kx+sPN9le2xX5f0UpxO45doZ6I2ztbHbwP9cPyKOBuBhQBVi5fx1f4G
8sQsTeeiyZQUzD6n5y1PgwLJPfRm6nSOSsNmqli8iaxV86xD/mt/3IuaZ4Y4WrZ88+wod20UIA6G
Ajd1m9fz7bGPIQVXoBcK+nESSyddY3FY3FofUrD42qrhmR8fDTtUaPLqRsQffzfTR3VmsrDsrFLI
CtlsJ9uuE3iv62tMvCpqOPOme/KXueYFHpc2rGBnbBMLbCGIZ8fS9yG9tAMKxxapRpF+/B8cE4z+
FzbbTJQV02Kfuz45Pp4qe1rZa7JWKRyZRSZqo9mTKdnNjwFTWRIHBqNeJNFKpURtdQeGVfKvdua6
D5hUi56aEX9f4afnzD1RNZfBbkMku6Kh5lbXqyouIToR3SPRTt7yTuvLpkvCki308a0V2xWmqHHq
tauNhlwZmgQhA5/tpSiKDVoXyb/e+AjgPxRZ8CvXqIO6ObC2j+74xRwi25B+QF/JlzcqWiYfcLV+
mUtd64xm4gXhCkpVXqkGuVuMnXqjjmTBfH8WV0HiTPoWQvEFaD8JBFE0YNV8Yfmmlh8YcTQf0rv+
n8oLNiOD7C3bUjSPLIiQEW/Ohjvs3mqbQ4ambPANor/0GSKV0u2dVp+iUqxsLBhGfSMCyNkb30Zg
h1Wd9MEBySyZS1f3Va3rzw1e4zxuIgRO7XeQpBrB5F/5O5bHhn0LZ6/eUKjBePOTgIpJZGlzbbfN
5t1PAfiTYcVRtqz+EjaoklBUku7yRmLrK5Ho3dxPJHZ+VJce+hJxIClFYzqa3pMSz2erGqpowikK
doiO43Ws5yiNgRoHCQg05Wro5+Jf51uR9/PyJu6kmGSQqiufHsHs5QkDmXkNFoPX1US2oH/0/PAk
udrPEJ00zo5hYbJmfcjy9V4tpxJ2jwPLYjF6caxYJTHDus8szBReJERm9U9IPbAQwZrpgB2brXd9
Rfr2dl8E55uhVT04zi9e6O4p7syQyV3f2Y4bhuRNR+BOWLmBf2N6VjwGhNSY/GfUV4bM9lyK49MB
KF3EAAtmpgAYZqnu2GxlPJ7OXVpzyOL28qR92eUGtCoT/+C6869F/fQ/M1XrUAqsonoYDqkP+xcb
qdw0z4L9NxL3NsjkyZSHMueSlg3NYNhvujJ7HQZ/pBnvOLA5Bt0Nn37CsN0uxZ61dvFXYIafJlZd
WINOu3FIGCPU01lKUzaS0rpqV3bVWKJW5ajPZfASePDLjQ274JtlQ1uDaKz2yecsJNfiKqN9pvpi
bgDKOhgiGphYoR3bj1xjqpN9gY5KrxYrwUO72Q2NAGU+U+T142Pp9TdNEQnMoLlpakSnGGissiah
rY9FiAMt86kJgHIEoeiAHhMd54gn9Gl1KiSd8cioXqPsIQ51eZXaHje0Gq+qMwiVfQa8zqGJsR8B
GNUJyJaU5O1bGPzrmc2NRG8iyIdmVX1dycWeXv4gCZdzJmK4IWFFEDcO7oRd+X+DFk1ME7GksPhe
HYMvwXqp0gvCTGu86vQMWZATqt3Em1yLL+qarbFFCXNKMHiB+Rc/HKx79UK6LEvjo2XJziTipysZ
Eqlj7nfMZ4FeLkGMy1TU9B/pmz/0TnxArBq2bF5rmVgWKbZQme4C7ju1Zh+aaj/+9HeLKlGGGNiC
66dXeZoV6kWk+hM4HAN1MpZHwFSIxXj1T76Zf412ZAAkcM59TwdWB0C9L4ZSKtyeE4TUhoADsRyA
Vi7yFfnYOJJkAk7QWRZolPZV8+a6SwCN9YguY4XPOrhcFHx6SSLDyoNEWTV8R73hllSC2Sszs03a
u4iMrWA56v4595KNTvL2yme2hjHyjWJh1uLo7wfvW5T7aHkHmGxAesD+LbQQqsUl5yGMjQiB+ClT
91Yd2c/m3SnTnp2qIGIAtrfxRs4J5W6vzlAUvIPOQ1Jmg6kUtD4CDtGY86zH6Joxalg/4fh43jV8
tfvr0JDY5nTOArVbb2fOgiWQ7v+NojrQwxLZDgBtuC6rWPlA2gJaLCPCSeMH2uzZ0EZQChU+Dx7o
GQrAiWEmY+2Z/z+UWaRY0vx63PliHNS6befrEhfwp3SGjVP3HxNKLo02h9Mk9WLXDvNVWZFhWD59
AsHULwfjaISWN7ImyyxFJEwhD+ES8YHtSYVRibcg4fGj6zR6VrMERgdd2IpU3S5OKWP/ARNkZ3mx
gt6M2vr7MDX+gkWdNLdszKLE79KAVnczQqq0Mw4qhl3tF1wnzhBwzUI7rkgY0h4aTL+FAFGY0NsF
6Aa1ZY3qZWNxprP/74Rjn7qGzA0McWrqrjzR3YzD/NalbhA72R/GWXeT70h9GMJ/bO4uWRCjC0Eg
7/oZxaIJ/a0EJ4y5rMbBSY6yiXFtkkJfDRdPv37Ie6H//yXDXCl7e4NOE91JdK3aPrFxDy3wbgeU
e1+ASgNCxUwyAWejR7OppZvfYNU4NFyxgUI6BkTQImlH44MdgGoNtiDs5leQrnTKQtY5oVhGU/4Z
iOu30rK30zf4MTfv8r2wUYKRweaET98YMq02kU73D+B9y1uZ1JDZYLZpRuPx41JcZwRhMZV3t+dW
FCePamDoxiKRajh88QCiH2GxsVT3SkoIOHt+gTU8ldWatWxTJe2fYsrppNujSriz64kbF+86bxWf
sNqdzX9o9tTp4ZGi3nLJ+9Y4aZYaiqu2seqUR5ZzZEh9l3wVyHXdBucuCMyiTI+QE5Gik/naJ4Eu
Ca2la9r4XZaL9983fBrazsoujrEqM+t27NyZCmrmGwkW/88R6X96+6b/J5bWnMZMP+U6DJAM0VcU
AevaLU3ReFljCJn6hsH3bWx9WfT8OPpmXwr9bGFLBO1VQbUyBOKyixMW/5yoL5yJGnJhya9wSUYX
7tq8KfFfbd42IsfjYYg51QgVgtaXxvYvi90gwqRqT2YeqS99V7N6jtlkba0bQrMjk8DodM55weOB
BN0M6z5LA+4Ociz0rdqFTjotatXqqf+uSCFhp4kp4o1Ivr+znLhoZnu6I7jAMEzea2SvoehSwlhS
NuVtvNrBERLJYobsMf8ZmSCsMcSURZR5I7+H2U5fy7lfO+Chgk90VMqdyPdMJWe27zZiRKWA+YJR
ejs77BgnzpgsqRzSRlvIZrJj0ZpOJOcX+nvDqxQZU5oORlU92NZ29qUpvftH1d8EQfGppMMkfY0z
X/rfe9Uzq6TH/vWI/761fRMDI1cFOzBlRAAZ5IgqIrdSO5AZJgxIfrr10AjrDZHq2a+WEBPeae9K
lzSmPXBCxt6GRdZLfvGubnEAYe4ebJJt/aytqNxRBb8Yh8cYnXcwg4VciKwHltTtZdosxgBwoyUV
OBUF/hrzUX++QHIrjJQk5HvBsk/hOiqEYKkHGMeIEL8YoqIQbnWJo1Ptlqbpm909OordTngC3dHT
j+ph/cGb8SablEvk1pNoNm5eivU3xDpLwsy//VEe4nvEf8k7Q+aGnGuxs5BknXoVpZ0pnc6EvCA1
XijEf9MI3b+gXikVY2u3wfle2DCXgvkICGJJj+xLza1/nH5K83IUCDHi0AzMq1pYC7dr6WsEwtMO
MkFBiV9OcZetfGnlCfZpzHZT7FBomxTv2xg2jFGakSHchAKhXTvnrGxzn2tvyBZ2XyfkqiFWqXmd
0BKZ/pJJ/6khWm2FHaOxPrZEwLlWZFq8hPZjKKUgFvjMiA/1XBOEHOLr155ctKOwx0bVsgvOvpAo
QE7hg46teD01H044tUAQPaARx86rV2OABloXAW6POuHYRXUUtvlMfvZC+IA3ocSDe3OKwNLgmjYG
GbUUsP15R2R0s4im3sfijpKynwLnH+5B+pbTMkwBgSANTtQO8Sk6IdwAWqyfv/KtGwtXeyoD3D4l
1l9A2qR7bkM/2m5XJPTCNwZF9pDQMDLIFplLelkttdB8p31W2n8FKvyGd/Jnql76+hV+qk8paGZu
HoUiYvccgXsiYkitGTpg5w7sKLzToHSUF5OaAwZV/pEQIW+W8QoEyTaG2ii3MRNAsA017ShSwv2c
BTpTlo95MdflWl7w9tCV1H4aEiQCSPqwXkU4KHc7aK6Tsr1yLF+9qt9axtgciaXWm55OglNEF+F8
OQ5MUmgSctNLEbDFNaUlM7Y02xuVPTeA2C2DrYyjCzVCcYEPxF08mflgRtMBPyKany2GdM+ILVzv
AL38pIFd3DQK4K6sCpHMkfC+N6AgM9JGUPCTlxU86pqFTQVdn14WIHPyexUI1gM/jTGzWF/0ZvsT
XTp7MATaeQ7+7RomDdyzXkcRd2Q2oEq8w1ix45gbRPhOGBUOe+rnZx4x2OBNvEbs3hJ61jR4U+rY
afTYTfRI5eKuOi7roho5DIQ7Z8UdYEOxfSCp7ZnaG0x2qZS+REEMVdqkUMlfBaZtOauzZpCBGqlf
mjUKOWqjAXCJ+0lyyY1MDsXS3N+Uw4lgmzXjLz+wcNrDTr2Bq7hlwE8mt5fKb8paMIS/7JvV9VSU
9TEQpi9lfGP3J62osK8Y4JpTFarOjXmgZwUrk/V9ZVDkRI0Ev6540fpstWLxJtLHJ3qDKWiakPKO
bDsu4Hs9IaK98LOahfVJtxhecs8wr6/uCcMI5pm/gthPYYppI0TNmi7qTnHg5FuxWR3mx5Zl8xOa
SqXcaKfPxCiTJO2NdJNEs/sZ9b2tStBSwnv8OJn4+LTUe69unYHB0t0s1+4VtDyGHFkh65KVDs68
1KoOWHpTOaJIQ3qqsF79xdp00QSvQ/dDMo9myYJVi8D4MAqtsEJ4WAP0f+XCvE6/HEN8MjrBnm9a
UFlVWKDahGzPtpYNfoKYUmVFwG/StC3O/TUz+Zr4xHc097Xjqk+Eq4+8/pUI4PSIjlvfrtArUCcB
2CEAP29efY6spKopAQ9L6un89ia5DqO+JsI/AcPAR8jWLbuSxTF/nIxxG5xQjPHRNnF9mE9JySzg
gqqikNQwDObrWGAt1PmWsV+HO9Jjrh1Ri/jpx//qKaFta2VZtToImQnALLEQCDRVZ5Bu0yZuUqz9
4K4z0iCjoGoTZuugvp1d3fUcFesYgr9wAi5I51/bUFCPiIC9r6Odc3MBbMKvhlz5JfMDdepy+G81
bh8X1yYmlb4NpQTdfLHlqQRK9evXuhuZxU9tVQCVF6LFw5ZmxT+jFdsqxkrwGZkdJGrl2QZAY3OF
NGC6LNMMVmiJjRim2WYhlw2ZOanbXrEFx0GLT408Yej6tA7kYCYFpCItnqS0ermyCyQW3Kc+ugp7
0ufsUFD36qnugmxTU/P4/HKagLTiPw6avr/VyYO/sSlIzXT3m+eXFhs+9czzPl19eHPDSYEVjxhN
yOn2Szpklq9mjyzCebQrGR74O5zEtzUDX/89MZdMV4ck8kQAb1f9oPS5ZX5TCu5VKAlnoIyT9J2g
7iBdYjusJrpBbEnK4hhjgGCBph6ZLYwe+JV8A3if/R/E1lrvpCJroxnsmZzm0gFkNRmlEOrW8frq
Uhp/iKjJ/Dfl/NxB12Z5Pb9IcWzpJiIzcytLLk1hYQ9SWokbhrebrZbrUIvRMPp/JiD22pCOmwnt
PVzsvMsDPjUjvL60pjJQwYDgq8vIoHlIug1wH7hwBJQimUgW2kg4MjEssw3Hg5kPFs/gg3L3AVi7
zNxLLQRc6Bauaka+7pM8SRMigUQDQmMNLnL7Mb2fCH/XEC4+CBFBS5KW3hkWUzF4H9kSdGuqD19t
YQGBMoLHb3wiPN5Ip4wYhGig2wllC5D+L4ffYoTVpy8keB2Jkg21a2bBHypNFlEZ++D36y0lKZaK
rmruciXvi89fMxIFMT0UzP8i/5oxDLfNY0m7ZtPfKfXILsMJZQiMOSK4QhIMxX6DFz0AnfVzFhN0
7xZndX8Xgqud5ZJJbFxNw8GI/Tsqy6/qOjD0XtWdIJXw5Dn6+RgiOEt2LAOoHLzV8/u/4Jjdc2fs
3CkchPhQy3rzrwpq0n8Slrlx4CJ7FOJD9kZqNctkNpntSR6h9z2lXTA9L4BsKFaZS5plLcBVrLeA
KyrB6nWiCEsznD4k4qR1J6O4UiOPdZm1VnOzujBLRtA7SV+Tf0A/GYSwaP/7COgEL32tB/8K9qmS
nDSnXfxpqm8IoRWxP7DHEom1gY0MYJRzovofFUcVfFmqGqVeLZVxfXlGmE9CWFDHuMnVvNcklxBA
UBrJ7myPpppjYqWmW5LW8C6js/0DOhT1FgDIClFi/wImgk1evdoYdQ2Lhk8aZELY0ZuKNHmmFKBg
liFqAVzhrLg8lZbVmX4xv89+gf7rcM/7xSYc5yo9S3Hopp95PTIY+y9rMdSGA4lq7ucUAp3DhDQU
v/AW6TVSy1RTrO5IZy7TGdB62XzVVfKB8pjuxTf1z+uFNkbsfqpU8Ye0vLxtcXhG/j43h71c01ju
wX3m/6hb+NRglr8zF0+N7a8WiyJSyNP/RQ2v6jSMyITXhvIe8xmTyfCNsUE406nMKBWD1inbQAAd
osfRRgNmYn6oxmvYuJkJvEC5q+vXNsS7hfp2ApZMZtztEUeFWvqvOEaSM7zjEseCLkSwEbswaq9r
8EEwrBM/Ptrdu37WI62+JYI06qBhcE/gPr0CMv3NrbCHKrnZty0NHtzjvV7s0Y0s40es/FJXdkNP
1A85GjOqowfshlGQRvZWB9Mh/d7e5d36jQXz6nPSy2j1hQZ5A/0rRTJ5gvMjFocg9IIaiEzPbV1A
EZwUvIcDJR7QsmR6LMM19lOVdaXMWnDFJqaCRbYOB+GeOiXO5S0XxhuuHAEGaM2YDZ5ytpc/+lmH
hi8B234euXXBbKVGqbF+KynQdcqPFgAb/7DxdcQ0OZ8fgl/kHvfTtPXzGseGv+YFBWB/ZldnNwur
7qVpT0aQueHk3DPjariN8Sh91MJLNlZnM5TAUAkBNRYZ0uPGVbHLz/6gRkEa4Man/XCP+nY2NXHy
2NCdQbp1bUjW5+h9QqJWvAbKxJSRtMErBiaQvH4/7CfE3qqItEGj2p9IJDcAkK8gtvytr6FSfRpC
USg77goFKyiQMy7JMIXrXRnK77uMMVHpxuzWP2XmBXZPPUDn0hNSRCMrEwjKEY8KJU59SZObd5gV
Sjf18W9Qinlx+/j+MtERGV8D9aoOLxGR6qZPuglJ3NVPT7+IwLrIj4ujtigdx4dI4xSfn0A5+ycR
BlqRoLxexEhVV1D0h58aJmyprECki7e3F1NyH7Jy36YnPEC5vx28nx6L/72xPim/swwONTnPFH+7
ob4sfQVHeEVmo/GAiSBYmkcOof/goTLN53TTPSDpx8Ogb0Zf8VMSIFkV9355urkNZwrFlhmhazn6
SxM8vaDJzOi8zjnA3/XenbdVy3viIIBGiaoyAPCJpiKwfvQgA7O9XzN4eI8hFe4fvhQmziWL4Gy9
cqxIvN7VGkJ5Jo0m1AJeul72CiirRCunitaF3rms4Ycc3YFqaB+eySHXMTzxEOSNCmIdO42Mh2NM
Aijb6AhBjfqEWBGoAWZQGEZ27Kv5Gp/pYKXrhjzhIMFx2mFQSiYaFBgzB1ihqYQO810OPs9c+xOM
XKgHCg76ibbVdusM9C2MGAToUtuKH1jFHNQCjmLMPfaRProFBSPxjfmyiyyeH4D679BaYh371rpT
iCMeeo/NHsB3eU7LHq3eOpcOdABMpcuqaKzHrsAPQpUGkxpl6qngrTs4sNYRLSOL6qA0lPpSy2km
2xM3MBns3gOXD7w7/3U+ZyU93VBKv9F8SOAH69Ng1TatzBn5Qlt73JvOfRRJTuBAQY4kSI7Yt+ZU
7mOz7TETe6tOKPoYmd9bXElh+L405hjBiY7FQj1Q+8AtOj+pmj/e92L9f4e6X8DGOO6zzB3XnWhC
mYuYI8XiaBEUSOsZG8IpNkVT0Cagc9nkAT+mDRFonEae6VHkrE7BQ+5fZ3MEl06+4DBD+WavYyQ0
hqjIOwKCkMBY+Twe+KL1EIpOUliYJYXzIU8Js7e+E0Ru48k+CKU/Q624ZP/YGC5dvx38QqVqPiMq
ISugGPrTbicAkFmFt8OXPGiWMVAoYtyOjAwicJr2I9lok1lzRoHD8Pt7ll3SmwisM/hE6XRi5lXp
O1KXu4VtVu2XucHzGCB3wQJHW+A+jro0GVbOrCCNgigeIQ29b3ByMRRUIQw/XPHHEPJs7AcKRS1C
iHs4CYeTK/nqa5W0KuQoC3rIt9wsm/rx4j/07OqhVz42h3ZKeQqkVPQ874y0BuBX83erNzLjm6Aa
vMf3L9ReNHLSj2aRgigrv9D4lTAsTzBa1oLlalsD6u8yBJZL+KOeL7AUWulfLMPTYEfFeAFt8uJO
2KBfHGZ3wiEmCfAW+vFtFbmQZf2px5DeUXYyU1AbfOHli+pAFUKLC0jtoHbjXk9bJ32uzaoq4cv9
MJvTcPTa4MhKBIPYxcBS/xck2WrpeHnWh4VJtSxOgUY/BYspzg81AnLlyc0WwjCHz66PqnYxIaIX
4PVn0Rqez7WmuGgUPvFHrfPmkQ2v+HE4SPMJ7jozbyd822XvCVY875GsNHBnRYmGM1WBM5GIhXgZ
h/2loNgDaWzf42a3kr8X+mpQaOq5272Qi8T32VvIy7401zd/TCQfKox7+n3xx9EUbcX6KqW14AWA
SQpq72HO3j8NaZH569K2/OabsnSvbBuiHdz/7AdrUWGXRJALkd8AG8byqGTLaXc5FkwtkZcUa9c2
9BVbjPjETtnkf9rrBmzXtztV8TmRfyxCzv2DMotXRA0KFSiuyMOnQBCPnAadD3+v1O+KFLCuafNT
nOvdw7b2b6eHh+izuZ7Lam5HknyXNHv3qfuHoVyZgsUpD6VH4WI3zglf3l+Gz6Mu4HxMLL6Sfraf
eYznukwS+yi69IZBXChcM5EucDSn5qEaHQSUGs6GRimT1pVwPDtRaBndtqDaWGJ86QDYWzE4qXHj
Go10/h4da4vFdpHsgbgHLy8yb+Nc5ZOzMgw6b/NigA45LTSVogz487cbOnknSH9Ochyzu4aYiftl
iJuAenKM7CCTPFVDnrLFVQx2NSNR3kc1mGrrxijXRm+VPhjmj6U+ot99eO9/7XR6KR2qZ1c10/Pd
UfV3mMzhchuDHRH8qWYtBZg7BhmCjb+dooAwvDtQGmfAQhzuyt2ExIvsm6quGX5J3qnCUVpsQoxf
4332eg2qzrZU7z1j99FgrXAOAvTSP1NcN8h8he95EMxW0/2FAAJd9XFSjD+gksjYfsnNfgJDjmbD
V8UBsWF4xlkNF1FZYuDLLuP64hqlyjrTtQ4/FbpDfVSmR1UI9y+LMLlaY8Wy0EX3Tsl9s7SLCbnT
p1bi86Ql9ytZsu0X6PNsf3fMghBoWNTwpck1AMNe1zg1i3WzcZ2++D36mfwTRpI2/KCJPlQTPGPb
aWoWWpLTN/QaO2KX2thuNvvaGNCPwPAAVieYF2a9vJrf/DpL8TqKdTANqP9efb1lait1csFJPNoq
0clVXUIVatvCLNSarEVRsPIj2BCL5crRrNFoJL/C0PoNK77GZZqjADroudoRmMp+ml1dFWcnpDdA
F2zmgNV0GqhoRaqSzNGBsHlOfGsp6yGdcP9vxxP6gSCg5nddhAtbWmhcpEmCjDKm18PGGHjjJNpC
clCIK+P6Fi97Kf566GtdwoBdrqKTqEcO4WfgGNShsOP10L93RUbjETvz1oTablsadKZYIdpz7MAc
LYdWRnDaHauEjN8TeLk85pp073X45LP5Dz6wiW2421Z/h/ocPytnkLgpv76pONxIJ/1TSqz+ih40
CkzcFqFl49WHMqs7h1ZPuZrQY1JuTy2GkGDNBEbGbXOzEK3GjoPWgE6HXwIk0BM9sULWim6E2kAE
RG7RDkPbjCJfnW6p0axQsQGvnAyKryROtOgM+2ul/xFqaAldvw6cuSe6S+6cIaYBVT6mA1tgmCiM
Ra/KVOKHnrDWpqVE3wEHC2FqUjUe/3EfCM283HS5ft3AQrX1DyZnntWfJIu8jMi6nWZ35G2ubxtW
pLOW9koxVBgF6JZ5jmJMYgWb1iiqE0dE/TJQfIXD1VMJY53EIYTOwx3JLlea8LV3MScyfjuFaw/R
ZxO0pBi57T/gE1xFwofpvZUvAcLH8bqJwfUwrMA4vcvVPgH/JpI+EupjxpR7Pqgz73s28agL+X3P
upUIKsv8wiP+iebwmvZOT0Nc19bX0kycm6hIY7Dey4iHZH2F8WUFWJWGQsn13yqa6w6Jq7cyp/wW
j1U3EBO+0rmYN+eLd4MnM5FcJMzEKLc5ch81iXfohsrkXs/Qu227OhYmIICRR/c5+u2tstyQdQjE
Vouja5dC6r+YGe5cNs1CiKjZSrxs9/4gOcWtnSUbtVnhMNAzKk11TuIEBqBX03gsY3nBQ3yXKMG3
bFI8sKhhRARFxo0RUFNhHKafsCK4EWcGMLei0wcvc7LuUfZQGWltiZ+Ft0PKLelRFfSJCzJzFD2v
uNSZ4papgJntG9PLnQsz4xM8HFdCuhey4Se1+crWdbJL+3oZ0Hl01609Hbv8yBuoHCMj5wMN1eA+
68dRW+o7wHjNU78STXfZtod5o705W7/7OV8MxKCyUOuzcRkKYVvjhGEGEy/0ly1y3rtSXkYqQufD
0BkYshNhzPGQyu7JUC+6yGBHgLsXkY+078/W8RwfqhERyoLCEoCPaZqlhC20a5cPetMkYbxlpFQg
B2CPf3jpQ27Z3HgCcHno625TMT0XwKdqxP5NV8xVqUHclF0reT6mslKl72iWVziI3Bhy9KbC17vE
YqszJntABSWiwsCHo4Hutmdp0mcrUxILuaZbnogcLTkjgxwmZgCfT22Fk1YCcBT/g6QtMH8+w1ta
VIeyK2exG8NbeTgbF5bLduxDDFAA95zsa3UrBTv7gdOmeeGXURlKuQXagu9J/siscWohmEQVp6JG
5NwwGJAgiGVuabe5m64BPK59H8Rk0FRqghoEvXF1duwygbg8bTOVOmvoiILFNNpNfK7A5VCAUCTX
58x/xxH4GtnMTayCLxxqfO9Ko1yoa1ergMb1Fgm7hTaU5b9GRJqi08uMLATqBZAzT6CSHwhbue+c
ggamawtTBWNeHSeHUB3SI4hhYUfg2hwfRDmmB+zpg5CrNy3Ke942fHogEzoeb42xm6GV8CU+3s3Y
wBBn6fCFGXnFceoh+rFTGFcaY2m32vBMsNXzE3A592HEgtKVE088ZMnfYAjV+hhgx+pBPN3sEBNE
1gnwmM82a+jx6NGoJ7cyE1mckplI1CF2OG0dA4ijOoTuEYwuj54VVNPrtKn+8lQGzx4jfae02dlj
6LKdN1BwLZanwgnEiPhKHwWEGC0XKhhNa6ngU25RjucL9lNy2oY9eXgVL7hwUMuEj0jz4pjXUkjn
Jq1DUck9SBP+Dkn3BnU1zV8LG3DudOicT/uxT9WY7hE3Gw4eb8sBRwG7luZ8sYtEn1CqU7tM3x+V
DwlzZ9DGCP8ozZWJf8ICmZ5bF6UmS2nSb/2lxVYHpe6B8w946hKAcNF9Pg0eb2EtnPo7dr9j2zkB
X3ATEy1cdA6FM6tacYB0+z6ZXKVWD+GTXKPgumBwX6M9CMZWMjJAyO5drFBeRgyzLpb2dCPqixKz
PJXo51XzXyAAsH2OY7sHP/lO93BOVkQwDcNdye+5fNQGv30pDC/aD7rp7Jg6+SKLRlrt2MY/AJx8
wp+YHi+mfjcgWQhF9CeXkzAtHntyHpZyS/7MdAZCPT1txnoesjyKkkmbHrf9RfYoQDnhqbvt1jGr
KQrVk/COyHJR067D62kND0ulva67F5+gm46RbiamNOWcSni/WlkKyO1wws/2uJ3NRc4rXMSivFOC
kHWJ/GASzeCXsfNWT++e+UR6RZl7M1t//gjkAotIZR+AwKmFPy7+xiDfrLEie0Y3tZSjENOr0gha
U+3UfsMOgxaHRncoFMgECewkwtLln/1r3ujDqaNZYRdTUdUphEECRMEFv2Vc3271N8DttcgJ1JPx
/8JQGmZJNfLNgNQDu820ONeDGcyRLzQ1ejIsQHjWQAZnRPvDlwL7h7gbmfH+r/quch2Ad2pBQ1WL
velbjFEa5Znwk09yv8yfduvkip6eCZamK8u+tiSQCx7oE2+gbTCRLP7whRIWJK2EFnSBktdgUS/A
NyKhyS3kJA7kF/cQ/WjJ/DLlVMNqSTyZMNP71OXcVS8Fk8iYZjMu16XBYy0lfdWMZSeK0APJa7Zs
Iolmj+AcGB9Uxp5USilGOk0/dc6iK9FF1A7Zh1XmYOChbESrFfSgpJTRi/3E7IYAbJY3c9oW2DCs
llJmZmK9SSu7JeEziGYUqheWpBTUm4VesVnHNz0vKsFjUV9Nr50BoNHRKbE+K/Khg7p247i3Ovi2
aQzPOhhP73SuRy1qQ/9pokfoX4JmTEwYtcG9k6WGv3HMQNJKfJY0ysozcDlmJSiBq5KFRnIkqxa2
vsbAnCVO0g5PedBEdHYAXPXG+xWd1Dby4G7K3FSZfSF1QDrn81NFm3RMMQ2/fgAMBYQyMU1kSBXI
mAMpU0z6kH5PFAKYSiqAnAdMcQbu6NzMYYXS23B5q3J1V9p6eHx+S+aYRHyVhgWbzUbCNaEunMbd
V13YwXHfZsJCJxM+QmAx7OCVD9niGIhgieZytdDSwYxeuFUg0RPu3TCBKhpDM1c6aY8LiysHZ4eb
bk/AcVUoI7ii2HqzSwHFq/OhrZ99z1A9g5TDef0mwl74DBvCZtIgwv7k/hfkPT3SUjG9ShWU2nbr
SZ+QmCqX33piYgqa3TPHowWOR9DOPJSIprpNXsQ7LnviISksBP8h+iz5DTlWc2xfiO9nM9LHAXfS
z1Bqb5cG5NCtqvT9Ab+mJVAgehc2GpA94Tnl8Cs3IYXmk+OYJrz/LopWW+PmCBFLDZ8iKOittC3N
KvuMRlN6RouTNI0A4mSuiDRKghUWjNmsTaBVJxUstbpUZ1udAxBrEiBM8tGH2Hyt6Pc+iCfo8Hxp
8FaCZZnSodFg7ySkC9cRByVZbtry8A5s/6hNdr2pl1f2JmzaDCVRIKPOiGrDSWX2gLJAEQBWFzhW
KKK7PN1WUnCfImo6IT0h/728xAymGqqy6QGJ2AlkngAKUtzfnR7oYxS77qselVxSkOrxBaAcZc4J
5FGLj5P7FgKXI197uUXevS6BKjjh/7G7q4qieaJrvEFGdHC72vpF8e+0VM1ULm7X7fjr8mnVfmqz
24QqASk+N9eQ7vJBCESfWN6nhBafM9fFDd2Y3EnFxPD1qjVdW1naxbMS48efK17RxOcHOo1FN1Xz
958bzcmXbtZDColJ/DuwyaLYuimaoRe0cJJ7FZDNhJvUF9CGMPKLMGlNeVKboh2F/dQU/qD0BqBl
/FN8VqgTh84mxLBd1GT9tsfeuDIG/CSf94i7sppYvA6KjC/NUq9xUul3e/iQmYDWmbo3x7TGS8q3
jgukumopdYpytjAtVKDCqe2FDYb4UEbFTJKssYvKPIQoTuGjLyMtNm/tVJ/bcSfLLscRUOzQpwht
ihKBWiogYYM1cNXoc9Gmr3VFA6kFmy+dRLjY8ykkagG8V58eo0ExjbwPiGglqChsE0HxZV6pmpPx
wA5f/WZJwTGa2CbzFYfuAiPPqitMUUgJ/C8C8OF2CUHtUW7eZjs376Fw36LJ3bcKWuJcv00qybdB
fTqSfjN0PHciHV1y75tZxamiqSrBcKxYEc0MtEmyU5Jv/qymZWDQdCu6IhpFh0UT651mh+YSrkZz
uYXgI+EahKuTDdwSL6haKeJXApNggmDdG0W10jRLsl3jvqCHMWftLV+hxtK4/s9ZDFuMKw7rKF/U
c5PcW1+gFy8gak73W4ivRptES63t0ACdLaMjVY0+04668+H4cdedSCpNAeA6dGOyfKlbRI9jABxZ
R18DwNaVA4ZSaHCvBoxxgBoexwkdOG4qnUY2m8IaelLGJaiSYDn/Kanl7ds3kPP5EhhlNJ4p0Xj5
VwXYcRpPUXqwRx3/xtN6dt+ObJ8DHA8GdLF1twLsfOkc9oL9uWOGwR5AB83EyTUGmzRLW6qkqHyD
X8vvTf4LRr5lJp8rtfye8i/vnM/ef66XIQhv6E9umBaGbJptaxXZA1hPgslH82BnlNXFEt8SbUkr
4bni2bf5lXkElRgJ8KyIgwLAHAe+Tc0VZbrYBCQbTRGy0wsDxRUEVCGkERmYXVR5FSd38YUgGz2w
82uq30mUwUTOFa+fqac0+2iBqELv9Pr3Q/6P1DCre/v7JNFWfbo0tfZMo+JlbNdpsPOn7MMVxcMk
Sj1uckvTmGuRKMR5mrqa3ZEAnuI76Y32/UM1te8H9gKzIpvJl79Egpwq5Z7UDCYYJMrIHCgxJijP
njBORbWp3d1CqMzl6oTLipTR4xmHNljh668lB5XrjGfU0+aVk3BMyHnm4lJCj5LqZyzDuusqtH5r
av7yx1D6oQ6nOfG96yzx9B+Ju8RJn70wtuM1QcIYOoc0bOwVz5rF0uwEZ75IPMsySYT8Z9cc+22e
ArJAYeTIWo/+AHieVLsa0lf41lHD1XcBGZAFF+wr5hlLVVC85+CfMEwFAjii8RtEznkZEYOt3AId
pVHkHVr99xxA3x4Z4AViUKnbuMc1CkF0auYX2cPOMw4tWGbcIDtBbo/cFBchl9cSIi5jJRo4rHSd
fJjDfCu/1ta5JZgeTWpXu/EFaGx4p3I65j9WbTpmKOBdkWXXmA+wlGnY76C8aMrAT6ksVDcXgWrG
kFUKTe+BCTweJWm1vYaFD7CYEkbA2IhgViKuqzM6Mh+sOa3qNeLMFApc4qN6T+1hJ3r3ickD2PVe
vO053BOHydfgJgGeVjvYTCFQC6l9M0uPpGuM90/kbJxhsNyeRsD7kxYUvAAcnTG629UsMYp+HOVR
AzEx8cYBrVTLjjRmyg6H5mShFCAmUd8ijmDp+Oz+eeLWC0v+IFpcplutURgGlYzZ5pVBB+Vyfp3t
1b6d7y8ZBJmEmx2wkA3FPmm9bl0/nHiwtWMUXB8UvK2/41AVhHd6Uh1sPxorYbopFe6d+j2dFhP5
60i/96XxehPRWfintHJOfqCwww0UZa/v4NxBlPqs1XLElojXW7hONM4fUfQAwq/h9R9w/AdFtFIW
31cOAhD2QFUo2iYGMHnn47WZyYZEjM5tlOFrdtlKMw41QlXtUrEodYBN+NNAkqS4ThzJsFCT9BC0
Ni3otdz45olp1rRdnLG7ACMjM/5UB8QcBl9QCSRjUDOyNF2EnsxR1Sy8RSIp16bt2cfZBA9/Psxk
+PN/PVWiJpowCAUCRUQJADUsb2K17puShfUE2OroiYx6DFz1w/OZiy6iXUkqnHYA3179NqMJ/ZfG
ZpUO84X6bTNghiJ+HKY6QoCuY6JAxRaVsVWpmlsTcOGrhCN43Nc7bA0vQuHgWEMN9jFZRzrUNxff
uPD6MEoKvQouUGn1auZ0Rs0ACgmHfz6CIyppKn+u0uv5V+DPmmmrmfO2yIcecq65MB83HN4AOf/M
hoBQCeQBfh0vdJ1cgezMrry4Z2y/KaTo+/QUj2KXrAWLbwGhdofNcTMHSUlnNNf/HWXZiqPNhwYs
qCqds6Ou2ir5QpCSwqFMAiKlyZAir9p3j8vcSVsEoxYg8ExGcV/PeufjD1pHErrNV+zMznhFW915
cEmukfcHYpbKE2iPvqFUdajYqWa3TYNBxbJriIWSXb8BsMy2kAZ7qGFCSKkMVXZ4AT6g4FzFkZaf
gNYhFIfeu2zVFCLXMbNtmpxonIDvxmVBF+vcC6seQt0XcEUvplNR8m+I7JV3OiSP9Nz+B/pNtbOL
LMHiYkmOL2f8jfhoA5WeqhAl95cZRKiqADeoL7T+h/eMkTLEDngKtrU4pPTg7SwE9JkJdkIUNqyh
OUDoTp0pbOVSMBs93EIN2EDg+1PwiR2bGqNekTM6RF5SpxwFL/yJxtTWDsbeeaOl3p8I/55akUCm
3wdi7H6uXOZzd4dpy6vuDbz9KJxXmUQ+qdaFYFBECprFf8o9IN64PQAVFooqjWDt5aS5+J3lT8fn
DsFE1yjX311ILnrAhL3Ja/QKLblGgMGvpnJVxV2sPZUFOG5DLU0jqbY/CTcaa5foxtqvChaGmkhy
3Ktnu1PutHv5CSUCT/A1DxTMotVUgbNYXbIRJKllc8k1lGd7kzQL24yf8xuScnc170xYSkHOOPMa
qECItnnAqEB3f4YVZbOVPtJtqCCEPAE66DtotSBArcX2tcqyjF04JycDD8e3oPPNKdpD4cJvRnwu
1ax52AgWWw4x5LcETu6aUYWv2b4IFULEmm5Cqfm1oDMFhcbLDM9w2TKfI//+Hvz/dyH1BD0cmK3b
y97DvPyErw0Gy63WgZXOQLFXuNYItNfJIaK9CA13HK8ouvqYG/4QE0a1pvpKVJx2Au0grzK3eFXw
H/ASMPaYprBUa6F5ienhzboeEfT3pNeIUtvSNeBcwFovEZrj4mhLOw8pb6coei+9jN5b+1jdGn7D
jdK+L2jDgUQIPovqmAjP/Ocuzg9DdDv1wnX/ZBS6Un6TaooQs7jxnUkZHGs4wEcaae5VMH6ynu0B
99RU8KxRYBdLlmZpnWwsP4C6OU3jzTl0vo0hpWtvlfvlBzDQqkkNsuzaisKM7E8/uHkuAuN/yUcu
3iI2Lg6ykuyoN1U7W7Aom7sL85Bcs1TxMBkhKYsLo1kucUj1nIZRjAthYuQpeKPI+9jDbx4SeMXH
ktKUgAJevuAVaaqrC0fMc1py2sqDwZlK5OGdv0vjYoh36tFtbnuCrLBroVmJ/2GrgvGUrc6wH/t0
yOayShiFnCppVMXsM92yRgLOMpmIGCEKJO8nru77J3DOYOWxs6rw47dLWpmwtS6w8EpKvGC1J3VX
XKnmtycT5SpEsCDU/IxWcHT+iCiryozrwm2DM+ogvjLa3hKa11YHVGF6pT/srFtyyVodYZv6uxGl
SFT+Xc0Tp0xRBCkmspVfBMEIvYnWQNuj0kMcpQDgxlAKRa3Lzre31qgugUQFMwaoCOVeOmHfqgXF
Jco3QTVycPpMZsS5llB8Oaj6TOjh80+r4ss3wEYgRPkEKFa/TInzXSKT8Fq2AEGXbkhU2OTTEcR2
xbnF/rP7jpiwHbwtw/+y88H3eLOClpUkEK4IT9YMHnshZPkfNw3v9GHIXrVTJYX9+G7hayOu12de
0IwCCOKtX8Kofy1grvtY7iK6hA/hK44VXgMZkHnN6tG1xLH2D2HVHaySvZ6bj7kBUk8uQRi3p8Nc
o+XDZE/kMaqdPAGKJpAL3MfnK8aepNZFSEJirAlVAJt4r4WWCOM5MmY/O6DgbwnJi4Gp5usgIE+/
7sImMvZ53PJ9VYnNQAdqLnaOzJn5wW3ncdfjt7LVvIkGpU2W5j5dKQDyIvpR/H6H7yZmMeqNFBoH
40c+DKSkqQnLdblui8fYYd4+nQipdirCngByX9lM9emYb5Y1q6MAB9E7fxxZYFB6ED242H0tEjmj
tYiCn5rh52k25zlpEuZZvWWOfMXG+W0KXMRMPp97D1ad/06+abQPCpzeg5XbYarN/qlkOW2kJPRa
wYneXX+Vw/7UUkJEMQ7a+aNbt1/tvG8nnd3xKnLPvZiQh98WVhlLVHUEkAuCc2TiVpTIb1G23qzE
YDtqMP8khBq0wrILR10uu6MUPOPy/tonbFd81WF1jz0PrEg3EmW/9mVTNRIxCB/BwnnmvbCf52QN
G+1bRzYUeglem5HFKakBsn9bsrHWywPwq7aH7SXefIh5DHqG4Fw6C/6mwVfe09fPBkW+MxZwwb7e
n1IXpfk5oAs/hf2YmMVZYV0FRfTmwPkfT1ROZAUeZUUN5f2/3bqE081qM+boa0lG8GpKaWrPr8F1
rExc1bAQHyvkxRaLcROixpLOIZmVdHPPaO6JGI+VLz6biWHXE7GWBVOpCSUc8BcsxaJ9K1ywetRW
4NQiM0JIGuyAYLSV034ezZhlV+Q0+pCazkd0u/CLB0fNv5JVMNP3K3jk/NSv7fzu3H/2/4+PZ0Z4
dX7QUpxzu9eA+DYfVSufOgY4fXGzTroJiSv3qzRUF19BUjGt4OWZqGShog2Cc9fCrliZxqFYWEhS
LJgcXCL1uyHTDETZCwPWnWjfZkhsNagbZFg7fDDhCNglXfy777S2Q3B4b8dB6zEZXqJgKdcwtnsI
pdlurrrD7Uxyis9eygHyi6OSKvwMfpQLRrmM5abnTJnhrCHhWkuXQ0LNlJQSP8+d/mqww/jpUsDc
9q6MTvCRqfm/kVVZFm7acziYxxq1jwYDjWvtPotlZy3uAFvj2uZvPSK/xjncpyw58us+OaDCU+SG
cwKvV3pU4Y+PvDT8wS6buGvn4Okd2y33wkbOnvIosyon9i0ewZXVuemuIp7ysG+YTbKlga2zRGTU
HSl+KzMamUkm4cUmvd9my2fWr85P8jyfD55aIZ7/wTZmbrY7hvDxp32eiC/ei2iVIApdkB31dL/y
Wl3qJptq1bdtXXqu1WfSxZIW7PCQNMk73MeCsAXD3A99v3EAie3d5cp+o7KSf8S6qC3+XOSITDfs
NjiX0fleiAti6Jijcwl1C+5ABZmAAfo7fIfBSop7HkjdzMy9jrAv+kW1udH9FnbQSrWdNv5Y0t8/
Jl6IE2/RQxdBb13gxb11K4F9pUNt9EgZLAQSuubzNWX1z/MIN2qyuTnal/OMvuN6MHZqK/sUYcRM
Sc0MuEi1j+NxnZBgsdvJkiFm+l7b9+qMBcO7uJ7PTZdVDwjoLRd8qd9DhXaPAaitKb9edEyEtGiO
tAYlOQgGSxmhrQvE20MjHwhnMyRB19ZSwxFakma6bH0JxXvZwl9f+KhBtDnNxElo9R5TzyGVMOgS
urxlhnzcFfJez5IGeI30O5HBDwoq/ouBO6vvbk8teH6uHJ5gNXJCSprq5+mXEWCIP348X8SVNmbO
ZrlMFrZWemMXlyPVwZRZJQ87XOtFK4efqqDz0VP8m7u0lS8n8FzFsW/BBV0gDK8OGSVE/Z3qwM5d
IUmOVJA6pCxZf4PmJp8Ikp5wUHGcVQL2GNgc+n3mf5+hPXs25straliLDbXYjmXamItplG6AXwS/
6c0MfQsbndALOv17aRBF9TLF3Deyuzy7lS1O+Nf8CrjpKV6HXMTheVU02YRoO71XMutiXwq9k9NK
qwi7RHCnJ8L1fHUiOr8s5Et+H4jabbn3/R+u008D+2wVJuUZPFK/rHl+bNFht0F68dFYHBEuNS9L
3QtmYDBKy/MqdZrFNv4Du5I9+NWi0cGYl9DgT58/IV5x7eGnti8t4Ic57Az3+PRKKGb59U4NfAY1
M9ck2nTfLtWzZEUWXWtXbyHd5RJAqods0QWWsD4d3lGPgpmHB7TS6fUVMwmdNpcw1k0TcIXUk38Z
sd1TTCxBHrIBDl/uLhT1Q+Mi77yvuYv7GEQO49ffL0UL2tRlxFpdLUvmXPKYhDU/tf+oQlBIZj7Z
nrb5jTTabs0jzGuk8LaM0vRXrCOE5MMITrjO9PAT1GGgNBNzAcHRNZl7aC5HAyoBXfsteeVQY/Fq
C256KJRUdYCUhiQU+btA0NlzOEl9IibqvDNAoyEoM+DGYH1iqQdUkMaeuJsBOHNf2RxZ/MyTHJYj
1jSvSKBE9aIKMpUCg34kwZo1tPrCUyxJMVhCykvX/oykdi42bBkd8o8l4fpINQJ8ERJU+euSzaZO
3Wr6CuX92+s+/hO33X34WGFz6+tWgW6pEJYV6NJGV+yd3eywG70EOtP5D96vk1p+0v8X1OQh0R/z
+QS0znEawjBeUqXGyUSEKIZWaIASYD75raG3IjrNnDR1SEKT9DCbFDzn3W3ewwwawx+8tXQD0v7b
/awQuSdnPI20xsQANqEKoDDsKoXGl5Sot7I/qSv+6s2aP1qqwq/D7COdnKnrgA3ZyAIPZZLW0QFd
CIfKdEq0GTlj6A+ikzOZ/taEg+6QvVSih+JBbLxFJaqiRR6K1acVjI+0B/o9YF5whZoydreYLTDC
4fx+anr/XsGN1+oKNOnWmmVrlzFC9gU7WwLgdM9cfqvxxneUGU4EfFHfHx36sqMnTJDWJi8/bjat
zzgIXhmGJezpGUiG30+m2Lbi+QzcWFETZiLudO2bNxQBvQZs7RRwmIRhTi3Iyl9xwkjooBDwEh21
4MIYfawmIhRai3lMqBx6Qrse2UqSM1N1h6wIXzu49f13vaEjihfrDl1ja+3PoYg52KKjjSpRdojy
0/S1ldSWJHOp+sXTlyvFYWWZ7deuufwfteXvP9xgF1rPgqSQr5/82b0CxeEHq3hmPoXXe4q2VCBq
cD4YQLtwreh6/NKAcK7Gwxwl2gY1iR2EMpOngvlqLgePzUQXr/Hl+ol2zTXnIfgQCIMJKvNAI39u
peo0R+QrrwBq1VZM7PRqGQJ2cxmZudU30BzlOye0z/+qXGw0lIwIqisTSS9MOF3qFONTvNN15cBJ
qd21BePRjyYbzYSRjx3bTwnPZc7gWTOUuZE4qnxd/m/U40ig9HgnxpLXojTF8T8roz5s0d6gB1IV
6WnfjSiR1l9Ldq8sEmH7lJPOXYHsCanZ45pBuGHEG2rvNaSuPlIixFszB6Q4KDRZkqgJlxcsFtdu
ncKMl7r70DufUOeHLWCQ/vlrZbTFBXYvo0cMmi6Dmd9Jm7AYRnzvC7ThGz2rRLS4SHErv2bGIw0O
FSid0DYrJX/qJRNgZz4UT1AXBt8qFGNBcZyHzspHmUoIuL6YAZfMAV56iUhYRVJc/Z9TvpnYlDKI
J1R2f/3ykKAuZkbWSwgefqNJqRgI3IaXiy5puor1wpH5bL+c3eh+39cD3+xfc0ln53G3mTfF9V01
FyBx1XOE63VcYeqkRGDSPIkvaPdzUeVqwKj40/V+DYqU0Piwav/HgxdBkdlnk0v2JIJyi9w7+/wE
QTDStcRvmn5QJczIMwKSYoiaTGfq485VLf1L5bTZq2kVBoSfoswwUQq0EJ9DsEp8yXYWZSKO+QS1
fd07yzFItpJoY9ZVXwSNcw1XlJFc13Fo+2jWM8hgTM0DLCPAupj5XRXvLx+dix2QqW1dFNrEdhvN
AhV1gwrAw1BcK/PWrh2QkLWGU4fJMxAGbhMDoo3tsJEmzu80aFiZRR5jTfNAUBQ1cBVXf8KlWA2B
CWjGogd3ez0sVeOAV/riFJ3G8szP8rSjZSGBRjHTKDYhJhepMOvHufXuwCctI9BqeZtnns10RloH
cm+Twl7cigQ+ks7UbW+i1iXdFlhnwYnTKCh3lSAIEvN0bFUkTEXkkuXC2VKofo6mGwVHGmOKjJQA
vaKGvKbviOFerkliNf0YrhH+ONcWbd41P6BYwp8De0uSdJb2dLNOHL18rD/7l3ljA3w4OX2LU4Pd
wSNaBKwYBB+iM5re/sJoNtKGQycspYWDJLMLWc3s87QwDWsDiZNORrUaTiLm+h5oHyH/bJTQhnz1
27unDvM9DWLnydA7vN9VxcZfDEZGpqOzycHCFEom9bz07Zuz3lf644DwrLraDYSESr86ZAZSXyMA
oIkeKuNOPDa0VwQToJ/A8GZAoPuNPXhqchT4WPIFviy0VFbRgk+zpoXW62O+vP/iz2wzOlv4ykYf
FV+2ihPCewwlQ8KoLjM/u+OgpLpZ5E5DUEcP0eKPkGrMGvBmBXng3jFvzdZ9YheY031qdHJwG/8+
NTByoOIqe312GKN012eOrQSXcotb80YD3l+cCnAzvNurR8m1eVuG5mUDl3H05SqQB25p+1ziSebS
4VI8r3gu7k9/g6qt2JKzRqmYiEbIJ68tI/wUHzdhAYFCwvtjzV2NqOc8H94TGXIC1YGCr0/SDJEH
1d7Wv24KN8uvMoCQBMvn12i/yHvWkBNXCizkuZMitzfmI5OfGBw/vHp9PeL2TX+mFFEcj+/5tEyC
oTQb0n+40jhMa/3kTmEO5Rq7qA6+EDTCnMp9DtuNL0XRWtTQB6YTusgkTbnD1zHJJdI/6YLsOlGh
BHVX1mB8r6f93JrhJjKN7Q/PNOdQEERb6aDRCEGlkMXS0kxTFDsk4fOPEboYTY3P6j8QmEdUXSbu
8i2MLc3WulTAbOZ3LzvZ6+D/wuB38ueViAhE6I1KdReaNTrERkppZcCJDN76DdI07v5PXWzp58Sh
5PJFnZ2sxHgB7ilODDaiEsflMNTeGDcrIAHrr9ihfJMjpsYyCL9LO06y50mjaEO9hMCJiH1dBu1g
FkuqZSQjkiWb/j2fAWiAtiZiIOZee3oFUI3vM06FnpH3JXllA2SB4Cpv9J2NuREW4V0IRWekC0UO
AU132c4zcBxsB8p1pl9+7D/bzHr1GcDQTJkJnvIZMnvUnbqFd6ZCTvBWemgIECjv3ijnMnKSE7Ea
YJcvSCig5SsTq6wp8OC806g+3gcCPom7jUIjCGncJNtjsqadPczjtvqaNZ/F6LgTI2sH0ABUX2KT
Igvw9btnLrS9ieX1Lhpb4LZ2feoYsvqoSR0Jx9qElVCN/IrWhTG08NJmsN5Hp2CgC/1ZLcxMarfu
Cjb5K86GjUOlvLc+YFEklZeHjj1Waq4HS4P+xHxwGQykmXJEinmKeDKSnMIUl5j+lkg57aNiHS3X
HKFkTSw345bc98Q9XuM1AvFoiGXR55HHrRP6D1K4GBu4h6iS6L+GO3CDzJ1Y0UT8xzyu8FmxiL69
TaQVizAI8yZOWCjPAYwsUmcCF4SLaVKy2h0a+1uQodi6PqhxNV6GVT/dagnby5DbuuVsDAR1frho
VgiGcay8wE0O7UIudyIVOhAJLxqqhKWkyg7uPnrtEWq6rDvFKcjSOuye5MF+ArCff36iy1ZoGqkq
d/iUDMj7Bk9N3qlNupIbQ8jkdSddPCH9KPspnbwkSGjNkKWYOsg06F5Bt3xfwJlupAS5nOgrtOxy
SHUJkuydUAz0nN21XDCi8TZQTRIZfqPcaS6benp+FQ2O9vlydU3Eos8x5mUaSyCTrEXAy7Czze38
YVaU1Y8xCndSHJTATdNamdFDUsIWTfrH0OVP3rooc6P3qRzCqjgUSMjgTzuK8T+rxY7Qj2vyC9pa
DO7/sHeVYmVA5TzG3dKvNjCOm9DWQe0m0EVn+oEMshsz45euiB+LpgvC6ZV9u5UrlqsjcCdfbXGB
UPKM42Nt2+9nSmJpz7lhzVi8COocyafg2AepoRuA0ZcjphWb/iYw4o+9bK8DtNkKqPScK9mBNRp6
rWtA9zLyy7IBAv/h8PjvG/zKvhMmnKnmf/aDHVRlHI8eqgNYZCnBh0G4+Y5t4cB5Yj9lsY7uswBm
0cgh14Ih8IkPAFkRkC1wW1ONCxRfScilHWnMaaYzTST7Veoo3PhizfnjOpavGE/XPdAbpWBOYJNl
EZVvyw9WuLOv+lS7+lUX4FfRXbrMqYke6Zj4fP7xin6wQBvhyUfzdL1n4300xTI1I7Av0rNUk9IR
fRD555NRJ//ov4uFWFsuCq4ycBf/p2H3YbhrDu4aYahafDd8ms/fz4s6tqXWerX7PgqXZSxQL0YV
JYFPjY9NOGhDY7ww2250WByKELT3F3FCQILk6RP6fvnlFRr0hKM+9HRN18sz6tGWczdB0NAMZCA/
AvrAeg4Ch3V0CDx2hMVSZZU3p7+zeYsIjJNFLCIUfa3p1p5Z9Z3GAvia/B/pW0DE/BpgWCyEBlOS
tJxJyZTbolfquu5EWq8izM0A0/JK2+4z/Ys3joJdnudZbVq9QWyO5nr3oR10HRML5vIG5oDvS5l2
jt+2Evv6O5fFCo2wkrxydRet8+ap+xZjPiyLZQMyAZxgO1u701Ohpwb+YRTLe0hUWarwoDI6reVr
zgk2bjSswj/qKxY3Wj9v2Lz1RKcXJJrliSgLjE0EV36wMXdCAdLrHNfpjCkdL6diuKEfVUQVTMUr
qidSeaPIFQX1bMSAOp4jUpBlPqY79m66LbnMEcoA28PVy708T06ZLXIXNWWVk5dn3IEksrJM7ino
bD7flg+AZuW3kx0gBzUUreQ/zYu4kAeNmk+vy3N467B1+PmgAExWHtYmPGevshKOXIlPdrAOJp+i
EHJH2Zi31HSH0wGbGhKrq82xOzOrnwIw1DgNATNrkWGDNqnaqNhm87PGUWyWJDgltQxEGxq06tUE
+bRuR1DlylJ7fMsykD+/P8zmxqS2MEvFX5Y/RJbCjPkiQ0mJlNOFQO6IpOSN8A6KUtJTzDk2oNpC
mSj5Xs1/s70rp5VgfhqwHZlQeYaTElotHQfo/mw0KNuigScZr1fvI8iwivqXXifn2wlUaceS+o7r
f8QBIoI8XeaMTiv9MsfvGzuhkOpKoX3SdVMOXT3cwPMDkxJHVDtBhqhvYf1/vHmUskq3vaLF43Wr
mdKltx8e5aHQT2K2RgVcPI5wCm8ejwZf9cAd97Ssib/LR+M3PXd5T93lHonvEQxpAoGvZv/5C0/J
1Bg/4b/oG8GGBB5fjbcYoXBKACX36nt4pqbrjsb7Ex3qPwXaj+eZWMSakkolqtBT1hgQR15aUrcq
IH8loqqqMYjybmMsKoE0nRIB8Yz/QDXdyKPLBIvk1/FuNd3c3nGXvcY8Y7aYDuvFk3wYX+VJHWYu
+/a77BYJipcv4DpHeYs1h2P2/yOQ50Kn8MsbF8MC2ba/y2rTiZNPpM2MNsoaT63gXxwDOTIO91yU
RXRo75iSb03C3j3kgjUXA+/NHqRFTDbejKscgBUZff2u8cnZsqZhkNiU1EEZR9UWuwZdRWSZgAuA
VJKXlM32SWSUbGkbb5xDyB7kNLDdlWIaa0FgF8y0/qKBg7xZSUxOg+xwMVe2W4tONv3gCcbeB7Zi
Rkr6datIJ0Snqfy0YdOnV+etxCvW5Qpj5uzHfDumxLLf5yRbn9hJoV8yAgVzuPSI81SdZj1O9v9G
f7s/KFdkANycKdYP4nl+0mqKY2qA0BbjNuE5WYC8gXdgSzEj0vLeJXScq4OwZ9SLQPnHzSy7EQrD
eBJc77t8ZZlNfYEjSny+mdZhabkv92/4aFik4e0/8xK2QeWWaeCEiru2xkDV4oAdXYxLk3NUWQel
yKFJvyG3q/JMT8oi/U3RdfCVqmHufURWTVV+uTFLDCc19z325EzFr+MQUrwTDZt0pR+Eg7Ox/sLH
1r/tPI9wra/EhiVHBMWAOi7GyunFzxdaPCqlFBtiNFNzUh8IuZGWz5JMcepqrzEcdnMPn+Wl0D9p
ECltG/D0US/RW9RrsUvoT2ak0qxz6FkrWJXAsWw093VCS/FQ8vdWWT+5QJ+WFk1Iel+Ws1RIj9rx
P/nQZmHSjxp4NGun+CR6L9fm8Hxu38WpJzrTt+zR1LuEnTKdkxZg58gAoynZBdb/a8LoxzIeHajw
imri04agT9tBHozb8OLDIB4PfU9bKh7I2s6Efrb49eb1rFg/LsBdC4VR/XUgH4nfZszMOwYzpXPJ
QCxWtK7OWea7bkHHZjUn/qIVAtzMWFQLYECgPPA+IT/GcrfKTmdry90KyUDSdMWUVqyAYz3GM9/M
J5+kzihGq3YftLdi5z+6kdtnchkiKA7e97Vz5FKZpSjq5yUlewryyK1HeJ53o6j5kLpAYtqCIQPP
RfDwWzezieoxHejox3zhSJPzr1E2hQzheOnP5j0ug/C/+iQ/uCSZAxRkAAxSXfVNZBe7Eo1oUNGE
BWWrd8ruVbuBtD3BuKt1xYhT4L+rhw4YvPgtTQSnXCO7Z9dTIkrzdKQfOqMw8U3mxM2mlbmew1cf
yvCOGHLTMEc16TWyTj5lKeDtnE0ofcz5sRRMtgAhQghZM5a0G9KHwPkiV3fL/zvC3HZcycrlgX8G
tej6aPwQw+br1sHb/BJQGWsUBRuLm49De6na69hi23CJWSEAMx401LjXzoFRE9gis4bfqCUe4G3T
1c2oQNrKmZHXJbQIDsirAZQPp+CcWpaQ3V+jo/eBkE6EWLexoEL7iIv3q1kG1YgGKIZjptRIWNN5
DOtS6CcOBpp95ftPHQHUF/YuUZrXMv06/r7VIFettdPeDDENrsws0EPgd7YjdDR4L2/HralEGQnY
EBlx8NFfA6bNytze8+1MB22nUSke//z0DZDzkkUpFBxM5Y1rtox8tJX20wUzD0MZH2puNa+kjRYz
QZn277uQ46d5hVTajj88njwPwCbkZGvdXzdwEpfTP7kP9JDJAro/Zv5So14eRpsCN2jiOSyHrRNG
CRHHq8LHvSSLZYAvtYXkh2ctM8NfcKAOoTBbzY9IqYQmg1hbIlpPwK3lSBJszAUbIdDnxKwZ8BKU
suNWIjYhtVRSKnYHiOBBiB9N2KtWzDgTBPyBMtcwAHpM+5iR5I0JLRvTjiawIdRxjTL+xv4CJ9Xf
WGdBWZ+Wjjp6s5/TEccEoWD0J9OhawlVoPSodJVgrExqVgYg74PozCONQcf4/w2XbFpWyzbdnb/9
BYINEY0E6jE4I0G1E1oz7q6TbCvkyNFXcDMEKBQ7COifuwh+gde+aVtRrJHJJy3BpZRN0h4W5GC5
1c+vmDUb3UFfLvb+BjgOSTzo8yyVSl3EbUggLlv1f+yWpHo0wVO4P5uepRGdPT49QAUN3xDBUnWC
RpW71akqBNzTBmy8ygsDP3fFk7qUHXLRLynSmrvs9iyYr6/jP8UbPnu1Ts6fnpmrxp343L2mnsB+
DjyNs/qY1jdW+XbB10+mywc/gpzHwT6yT6MWQ91U1Cu71o/Gj3H1BPUeEYvgHDOS8bOpPj/UXpVD
Uog89vYMua1ATjHzyZFZmM4iHQkMfYQoSxy43H26aQftslv0Id6fbUQDv5A4JUmh/V9sTX7d339C
eI3/HuYFlzWDpmmDsqNW3Fo/6QhsDzk5koFN20yYmSG40nnNqisByrIvnyl7ZhXEqe2V8GK2lH+t
/RQRYJ/EQBRLjHQLRskXdTSc2fSRC6VGRbJcBUpL06LtA/dIzDJ8EbFFbwMrBkLRBMa6xAf5zVLd
3dAmhuMi58ypAxP/jrogpsOPL8LWxENdTCEC3sIoRCN84oo6b37UA5IXe+BF4aycUkAzyq6vtQmu
174mwXDXpQsbo4cqKAJ4YbGB/oJwa+2mSfV7TWG2gsfphCce9K37h2gfAbgMW8ICzwCoCDvSzr/f
5gMkHfOwVloYhwNbsZJmDV/lVmo8vnrBFQ862rdPTgyQd+ibHgoeZw8q3IzXkptfVXSJkVpOUU45
4h7HDVzjjUEIWA0r9apKEYoajGobFCaCiFzaggE+UamBHcpuHRfuALk2kWKbyeOcsecdhUXRbrtn
rLaQmizZYDw3x6n2E73pP6buk+yNh8LJf++6LYHsmXMT5k8xuyEPMEj+7mNFym/oufAjSL3BMLrl
9z4UGGpTig8/bIvMU/I2R19l7q/OgIUC9tWzGE0zT/YXuvj9RIC5liEX3n6ldHkN1a5HvsY5j3y3
ZdROeTL7WBw7WZoj5vrK4lezHqqXEgSl5jtZq93rhymlcS+nAz8H1jktkg1SGHlCp82vs56Yy/ay
Rmxny/DFW8aznZkKVGw12WCZWOz/QMYcNlyP3ND887N/HTEW5YfWS7z87kVafjuxu5EFyCiOGhUp
r8HygiVLAXtspMUyDAjlPkOrfddX+0zci8YOaLkMNC6PkI4xeeecuECo8OxImj2qqsw/K7otJxe4
v3vQm1EXZX0BMAQ0thG7TFDs4OfIoxTHvLeI4F3C4IiI9TyxnbZYkStwpXullRDgAbDuvZCQjfRv
ZIgf5eKB0sBwphM3/5X16fWTHX+qbfNfKFr19WnIGWABn04IyqTq5lqZISQAACRKkwXJi31WFL+T
bwZmZG5iORRvAnyxScWBertW90fWtLg8OB/IDBXedai6v8vG4KMf1K+IVg4sJDPJaUI8lPQ6AgBy
fkXiAKUVRGKCbP84mNbjOKp3hbsMn0i7BJzV2uaxNCzqJTddSGBhwgW0dWoQk56jCzr2rNva30Rc
eab2GSVyNyBwmkrhHVycXcaiWMpjvU3E0N63xLZRaZoeLt7HARUfs1/yRu5KSb/08zfzaVVV+NdJ
M2Jrkwh1GDUldxh1T4Ns3fFDRcm8vYQAnzyX+pOl27s2b1w1+no6yj6zyFg3KZ2PzYSiztnUGogN
GwbGBgEDyIBpNZ/BHWEeOKZWnwN6aW4XNZnKQ9O/d/HUX6xQ8jPrVDTpt37UMON6Z9l8p52LtKuJ
zcMKf87vzfE/VlqCpw5r1JgBAf9MDpVcmIp9PUC+zzrUpNDYqd+y/tSFVFcjIG2xKkCbXxSUZhy5
PJWKBOR3ICJJ0tVHIHNjE6iiMI5JDxQQUPw6VccUaC4KszTJxq8ZECQ6eGu3a1IK6aXC3QJJJqwA
fdskF/XiufAF1vxEmRRWqQ7LxhxIW0CNZ7wjysupjDnClwOdKFlbnl8gRi97+8f5WalICODI3sLz
s/VTiHOZXNkObJvh0YaIfXaMhOFFoE8RZPKld+bIgqt8wUwOf8s4hG/ZhMW2E9Mp5kwor6WSODLf
4HDxntQUDwXzl+f8DXuZNhuU5MKYhRcbYIxeBDOtuGdANHDuiran8cPLSmHZxatDubP/PUZG4jK7
IhJbv+6p9CSj14e1DNkLkBhnoRC9OJJaQHBNmCa+J44VN2f78C3QzZZdzXlc4d7jH7DnNnO9z1mm
GJ2VCIBnodJEnVH4vqNW7u/z7B6FnKKyjvj6EcqNl/RjyDMQ6ilsmYNu/MZ0mHN4MGnctu55h+Tz
fhblUV6DkMMYCqLrZ9GVb0/hr/SjsGaEFXoBbP4pYc9gFC3Y+G8akuq2XjlZHsds/5P0nXILgbZn
bdL2GF4ZfDEYi6QLTFACwirQfnbLk+GTKuYHkjnZPD0YkZ4TTk8AMOA/kCAPf+vjMrWsBr1NUQWv
obdp4x8NuarOnFe+56pHN25GK9/JOEnFLpfulxTlaOc+fbMBbM7GeQYn+rscM1mERZmUz0xtmmDr
8QlzLZIvCqctahx4eQaP2pyTw4Fa/rMdW8FzpQuULKtA2Cfg1jyIB0xKoRk5zHgcXSs5vnmKPHV7
jNYMlMdafidFKma/gfWGouXwHxZ9bEdOaLRZmb6OZFrZofvPVdS+v+oASTxZMka1QTWaMFRy6MPW
1RXpUmxPJxerJg3vl82ISWxEUmc4efTw1EVhrUPSzvJ7IVhFfcI4NMGcT3tpj4Eb0rOYfw350o+x
yX5w9+/U74S0aUnTgDXGGEC8j2iSRPU3Th+4MNLkaTAjB6I/uF9VBVc1JCDYCD8hsu+u/zZTV4Mr
+9ic6ntwrPNh0WVqGATCRWWh55Hye+RdRY0MFoSiA+ZH5R9piQ4lh+xNIkvBfnKcCruo2L2PBSkr
vBbNo3kP9YHBeN8RyEKWyWmPMDhe6vObVew86oQv1M58lZGsMXrXPXzWgI2kVOTtrKrwWO/x7uDE
FxT9urva1O40bkl50+2GixiPgQiGRuGt/la8XicoOisbCA3/QcrrYpvuq2O1peDeBAyc45lsybgW
dfhF90bS/Ug8maXbstbEoMTQqGQY3zSURYEA5ELJ3DbrmSYDWfqGEoDdmFtiI6GedOuYERSrlpIo
cxWr9yjxjXEwt0h7NdVH24aGgJ1tD1+/SEDT3cuKrfDJbFaKv6NZ5xe04UEnJhp0JQK47Z/Ny4gF
uHaQBAa8hor7vGieGjl9yZ1wN8jz6K1Pb700EFeSy7zEXuvzo8wn6G2xjPCxvA8/VkDa229IWA9t
NbsEvQn7WFE6OyI0r4hnuHGgPkxr/l5mub7KdDxVORjWf8EJuyvWBOxcEdhrrcHpO/RwZ1ueOuJj
ft9cpf2pfzBzc4Cg1oeFJzrwoIxalxZtw/K5vORxqyiVIkx0+zBFQtnrqrgkBcGxSz7LIlkIGV9s
E1yFAgeeKSVxyu6kNQVt68D8y27jDpo4FLq7gvMp0o+6rMVahNctcRUksrzC7hf3KJSDq3eGlawD
2x254ObJATO+wAhemALjfdiB7H807GmpbTupvuVSdad/vPM8GX6nEicsSKlfwbWcwE6/Wtk77BLg
U5MDIUPEnIfGn0/LlDlxuqpEDRzqXYOCOsAc4diVT/7hPMgZqQxp4B4lbxAylnthPGQSF4+PQfKy
Dj+ntJ9oDE/9rlG/kjlJIbJlo3igmgB+MJDBC9/At/eMU5XAPN5SmsyUNjJ+jHfUe8SRx9nEZCrc
d/1T8NdTQfw2FWLCTZTnPYkdBy42T5vGd4yvqgolXvgkrJmIctwWsec0yzNXEZEw99eckb1B697b
OvYYG5Y5LeQMH66rdZj4kPi8HpaKeiOj+myON5V230I3zCCBaPKFK6b/L1Wqy0o7Y4DeDYbdNWrx
yHPifE/jNm9yGO9blhd0Jj5Cx5utGBhf+hZt0ZjAmqbXwKU/o2Q4iF3Pe1r/ruUQw2ei5Jshaoch
R0ATHqxy4IMKaImqtd3VCPNb0YU46/9bsE4BY6c1ZfcaS5Oep2oJGYra8iRizrvWzwPCE/qONUaK
resLnhkD/sxzQUrCln2Ep2wl7q+gpC39YdVgzFutSwq5MIeOwV5saJPHvOVywdWmJSbFrP/QYSLs
VC6RGkzuFVAXs8AZUK2sCHRCbSZKHfBRyTw+sFZLgRM/MTnAb0zcepMuF69L95q5WPA1Qbu9Uo7J
dTR8Naxifll0dmNggDYih/p2gfw1OlbC5+M8Yf5JyWXifSQNKcTvHs/7j9T0OHymtkqqiFoOwKHx
Un3zOTi8ETPb0Jf48AnyGxpKTGln078FBI2DTdhfZWwT0oBctmcREd9OVe72zL08vt/jZdqKQy+i
bHaFeuWnP9HaC0NN4WMkQCRZ6jaGuCK+8PnXW92oI7ToBAFhCsV9ms6jraATq56BidMtJoDioYGr
27mOvH3z0vC34kxH5VKb9mmiA+kNodG+wWgcXE0nzatfZAN8KM6Pf0F/Sb3lCyN4TnnAXKfn1ubl
JvMzQwMFWEPVKcVjjQPCqRGtP15ab1FDmT6sxHtkHYou4eCJGXbgDhW/PrsjL/ie70f+eogvrJ67
mewcz6lDnxiJQ1gnuFknPKqd8Ata+VF/H9CMqeBBkH77EMdka/rDpgn4UT8fDNStc+qMYsMrBTV3
sEGsY1F3yidJAmO0tOEtUVtOCsWQJHMe1/tndE6h/9/MAWNAmRNd5+BKV4h3cCRebrUHeLPfaHYq
W4SxdW0teTTE4jaSUJE2O6DUcnn3IiaTC/wpRXtLps7BuY6HXNcbWfj+vwx0Ge0F+HRN9k2pz0iV
lUP6LmDt9IANPpAoiw+7JZWvf0PMGphi7wbtIoOxFgLeBY5OB1fZtYIK6N/+3UbL5gRg2NouHq9o
Bk+MOcP1/VPvcmak+29DVrN23HWGdAXX1MVe7Jt0Gkq4duU6Ug0Hna42IP77fqG3H5wdXsC4LD5z
juKDfw7jik4m0avHt08JyFGb7y86IlkQiq00JadTPJxO5yNBorwPQEM6N+G2NBy4OFE/deEmrKgH
ZuvESm29DlkPCx/OoDiQtHbcpp7QpbMZHBaFGplIf0E6847GRrn0FGSjsuhxwQdgfh4VKLmZUnwW
EoQUeUXMekQFBxM/bZbwabby1w7WDDKtz//gShuF78KxonrFNVMmEFpAsbwpAW9rjw/s2pPWhtal
e0VEPsNb/RZatZkSyuQFp/c+wOVF17zuaxGQR8oi2L8KaY+z0/ByaIQBxUgJI+VBQ7X8g+Ky+OV+
4/xV5yi9qhOgn5XOlB+uSUkA/r0Yn5YrhWUNZVbz0996rUTxlD9wpSMsK6+k1k4/SihjnPTIW7fV
+0cRpZlDOq6RU42JwLW+bgqV/YDA/ZtxOFmJEFnQQ3gqZ4iPfzg+BwxSWX5j4wXYVKpELaJQfqMR
SlF974WgSku+1Dr+re4dI5lhcaQajvzpTIIJHwi+aLxTYwzLsnGGPC7r1pGmDHvj5M7Q7ewZ2cOL
c2e7TLyMjwCSUBOqIZggK6/revkcGK8LTvpiL6fyrssDiZMU9M6w4mBADtGVGXk+TN7cxlir5dNY
3rXmLnA2ELmwlmbfrG+qQkBem2J+wzzUk9rA3h07dy6eR9ekkFwLvbzRuDR2w5YZ1bOXXkHmF7tA
kUxfbkDgI/2ROZbzgVURv/E/gXV3JJkkaN1us/VQU20HEyfMOpcrNF/u12F8X55rhTH3+MGv9zBB
0Yeul8ClYStlt6LMsGeR7pnuH80gQJ3znKSTMTosdZk41mVtS0hBzusVj1DCGPmsDj4LeTMVQa/a
9FQSS9hJb6ztncExA3Ol9Y3TeKv12LTiTs2uFFLoQ34oJUv1uSGbEZJh/GCrWQn4IZYuyqji9rQr
1PZ1X93RJlR2m+JabO4QriJqn+E5D4AOj1u727quwfkOOJxAglD1GwwCZCsuprmYCMlFBe/3V6UG
l7XyECgCI1rEa1yQ6l06E8zQFxe61eRnyfSKOkrmD89Uv2uo5RBCluLH+0bH2Ng6v8npArSth6nG
kZKIQ6MzFTgEif94rXkwKVQpnXUWr6Kw6BLtj3+e+D+tpQg3TxBU1rl/nGLYwmsLMt3qyXFCUeA9
PdndlvZoG7J72S7Dk44XQj2R8N3lLpG4LH/34FsyteE5DFErBNnWN3h1X6j81KG6si/Ao8SrWl/9
DykUOSS96DnZY/QXsmeirKFDNFrJH9r2tHpygvICEEX6RDbNjoz8q4F1EnDZL5fOVQ+7E6ruS/fS
w3pUYx5mFxmCPvTVrnf6037M7HUkmK4O+qKVuDWKqF8qiXo9YnPnt7nEtupnij/PyjMcWHPhGX3a
x2SlhiEhJ65s0JlCXxp3E5iaCRhd3xGl4qpCfxe4eeeK4nAIQoP57Ctbu4dfbTloeLNWjUw7CSUm
woZdO6NNyFvHmjvuf+qPak1z4i5a8GwKToImp/VAnBD/vLuyw7ghi0+Wm8dAXAC2dnF16Ill2AYd
eWjrrLltfMUWPZ+5pa3BJQsA+j7iwbkaO1W0TZ2WxtN+eqglv+TlCLOBE3BFp/RB0n/g8Y9ZGXLk
9oKhiw0ezSKT9TlN9IWpMLaUfwl1xnpnDv08gWUrFcoplIy2aLUwUTXtrIAGs9OW/Yrav2a8UnnB
JG8Oj/byPFNa78myGNku0/KxLK9Ew89HVixf/YYzd+3o9VYdw9vmles4PdYlpjsmf78HYiGfFqTH
4kRn0WbTToIHxWg/qdRMVLNKF6/TMGRwLka7pyyeSyueQADZ6oOj7mm3+KdhvL/2Qd0tWGBz3Yuu
JWCHMUL9mOnLxZ2g+nTmcKUM87KmvvAPbfXVlJgytjA1UrDLKqq8NgVCU6E8IJ0mPdyGQWterpr2
t+joQGe9tA7B6ZnQwrVHOup9/hGkSM6Apumihujl0nwAJEwYUqY+qVQYUgf8NqOtKZFq0/bP78WJ
wewB3H8K7o29xAVGHs6RUmetoHtAadkLWj79XNUpN01XieQqOZB+Wyw+8LMgfxwBBBtwcPtGNCD+
mGeJnivZ1jwtTfwag5qOWy87efK41ppDty+3gF3VqHFvnxNv6xUmfT2oXuYUFKW6w9zJ06ana/5N
CQE2wcC3h44oxA4pQm+co3kSf333gf3xkb8ZJXg7E19m4BqN+BzjITCVaWBXA8gOU2ANAVswtvjE
+mZP+HLQ9Gj/pKEs1YTn4Q8yRpOzg14SSQsPVd8iLScEBo2M0FHLXTYFAu6QGLamjsiLXDsU0Ey1
ZdytHvdU/h+8EAGn8qiKND9TeIT/tw7eS7nT3S4WicS4R5K4OaaB2yDXFVUOGWwHhIPbcHi+pr5z
PWJITZ5/V+rFbCtkjRmp2rzinlpBQ/rMDO+NgLx8F8+lSO+K4N5wMqw2RG2N1i4ESFGkJ8rwoEor
El3lnVprBmigAv7/5VOezirCa85Tx2eNCn4iWShijeyy5sVyIl8DMpx4XlukxWtbxDOP+I8k7uJC
2h1bevLoquF1aGk2nWZiJWiWr5tb/ngzRgpVTZu01G8n28DMU/L+M+rzYVRtgTMJoOTTsoWrshjb
KhO6wDTWnJAGNXJKBE6HKgDXq2xZYxcWeBkL/uobNiLNDEvSjHsqbv6hT0draih6SQixXl/qqkWN
7IJGE2ga9kt5hL9zo1fWtwFwFOcJmVW2bWqGW4L2bUpCS/zUAYOkppKCkUBPK8lHikAEECjr7GKR
Lz8q4lhWLvcHcZ0s5CF7x/6i9U1/ipjWRR6CpXU9tsCGzEP8ZonrO1Uo1p6Mk+jNgTuNvQ2qU02x
dGW41/m1+JTa2e+m8mEYp+UWpgSv7BJKTi9cFV1nZQWc/oIMw++ZuhTvvTH46wpW+x4cSJd1jPU+
hmYtJDUR7obMQnrQtwPHarC7wo4pofwTQzK2pW9v9hsQl6KrWlsjPv2gvlsBk26usEn/GwlhO/3I
Z2iEr533501QQKNzVdoaVqyZmzTJFHgLcmU0PzldJVVXi6jwts0kgdtTi9ESlp1eNZ1oQfMHqXMS
gSzKjI3/lBgh1HsOrvX14HzVxgRRdMdblarqsFF5pmH46ElWus1Lp6n3841M5KViFjPFl52HEvt3
NZ5DBENUcAlcNRoQtDSSym5cvpZIy2l0sTtFkxEIVXcjqAjCGyCEyoZXvERMuHpQQLqJ95OUp63t
ZzvtO0202TAA3MfKaI3SDYZvH+Vjtl9bqBR0lmdE5DDZBzT0xzxkkil86r1xQPEjAaJe8FDRuA90
pgxBWZgemXXPIFcQQZS0IjOJwNi5zfpDP3Qcer1lNJAe+msLBGnFy4kxqbN9I7/zmI9X9wl+dQER
vZD5ff31eoEcyLslvX486cz2/zAMh2oDhhEGEfGCf0phYtLh0dcRgKyEEAdyu9aesnZdB6MwnAEU
M4lg2gaOK8TUZcRLO/3Kmm+HKDGIeWESIkdv8xFsy9wcvgboj4nFbfvpSUJyykbmLVhOZ0T2DWlx
VnT+MEbFWPaKLOzQw7DFUq6iR/FMYek+dfCwon5VPMd2cyLvjotQ5s2nTQ7Tpnn5Ssk+RucMOAH/
c2a2dCVG/R1DpEpELrnXzPMRyYlQBhgukFfZP/HwMij2nYf6QhKROd1adyYdrN6R9PKnSMzR0AwK
SGz9dPyVPOmdfZb7Tv7U0GH0gnVHIVEjyaq+W6E2C4lmMVzwM+gkTH1OYB397ZuMAEpnycMbZl7K
1XKox3vQvjM2h1iFcZDrnuZSpGA5U18g2iCI07e6hoa+b+nEpQ07X5IxXEu6V7sL6i3G07Le7J/W
hi/xnBhA2hvQreqiCk2VGKRySGiezHw6PPHp8avYCtWO2TtLn0SmrIwevSU+EV/b3fH+cDU2vErL
2O1afJ6LFaovuzG4yrvJoicNFVLIxhoZwbI6NgbQgYBBdH0xaxnOq9O0DLZS/SqnG+sW7d9dcSmz
wAb8Gfypwde6vIL4KPdZ0fmxc5eT6ilYappJ7Ufci0JoGKNa7Wcgd+1qkGWU3heqJYIdliJE2dWQ
EBb9okWBzqU6qTA0ViLCA+YsdQ95xXreTxgGedF3uEcglIs+SAUsURYrLHrPbWff/0+c3WcSso7I
F4tq97bVd4xfIMQlZPojcgAkc8hi99MSqZsYPPwn0PFlo+I8aP+pUDjJYrTgV11UKw/2ktIuyAwy
0vyEIzouEgeKA+LC/VM1ANdBvVQfjs/4+FZaJEsYxZne5SXeIaiRDN6jhb7nC7yVGhkKwAtc/0RX
yk79ljWQFdAekoLHUvJH7xvARHPAO6ZL7ghvlhwdpFh2cnGqaUo8/mcO9KS0RLhMjL41xo1Tq5am
2HNEEfbrnSnEFT+X2z2HfqBzj6F9/XRhuZKEaOleJbiP0N41lqR21uA0lkGdNLSd+Z6aPk/x/oe7
q2W/0hu+0tapO21Rz8noNxubBVMEFIwEOLlNJkkrxu4g2J89pP7qwBDILcZUsnq9JfUsrPus6kSV
szlW/fxvXVoEm8+p5q7eLrMI4gl8BXoC5WGdOM8jBJ78XjrZu1SMgME0qUhKr6pTmlt7GgI66vv/
qxQSL9fkrC+wC97vzme8KNAG9Hd7BNLEqmVHCsGu3AmS3SR4jBjy5JsH86Ojr3yeWObiEE2/SGTR
73PCiTvdo/EN4OAtghkdqOvvHT4DChQcEZz5u6lBlGq+LDD7V6sJMO0eQTjNhR394IIC7aQD6IZK
iJPogEqSQJB41cJJxYgZHcLAc5Ij1b9jREq1MtDQnDoXSW7RFD8/4ZuZAENVQSmniCy9HI2QmDUn
cFkWgB85/zssF8RmoVL/1R3jyrxOSrWup00PM4Ixczsx9SU3EeJqw3QmE8/bnm+AHmlwsfXXjQrJ
Wid/IRTtIwrnK0Pw7P5T7FXRNrRADGauAMA4gyLuVAQ3hRsw52nTJZ+kNWL7mYi891n/JqUpRAIs
gyT3uSrq5opIOwjOYpJ5h2qUiBkAGGrHHXW/ryRqn9fDEokm/0SXpfbZYWyyq189zVneDo8/Hwwa
74EejzLxa6hH8LZHKZfseegVeffIhRv0eItb+9zjuFGgtpcp8Xn8guMuWQc/cvPCjGeBo1cwxRsq
OqVJiUqBTuVPkAzPfRws4qs6xlIscczhQalYvJXCNgmq4BrJa55ilOo4sRsDoLUfzAtVBvFlYMHf
EEIYWfFyepOIvWLtTJnqfRyIitnXXvfAQtMvAxxtUK4muVoXofz4vS9sNOapwBLl+wTs3jBCterv
Enbm8xJRq/ZPKpt7Mbk1tA5tB9lFgv5zC7NcEoWSeEAXZvjHu2rXuKRGdiixidKo1CpTsexNgoDv
/0VjUTftWlFif0/VU2NcHXKc6R+Jv0AHEvsLpKlX11WFgvREPbBLesW72uEK5jAn3JdT+Ls48wlv
8romnDRTfVT5yitCSO/iRTFFiTBZ/qKY9OOvJuDCqB+8uLqksbBOxomj6Y+XH6rM+QfD0YwPk+VO
Od7YZhlQt8cLMBV2n0QCoN7XlQ03j6bdMyeiTPKAoh5OkzQG2C/luEzZckBKi/WbeD9a5vMInS6Z
jkbUUciTuZ0+3yNY/TKk6GO3ea1nlhpsAvqrHyC1GZUTDW0eor1WgpgJ7uY/qXcxLCYe4qfwuZOy
pPDBkwghtMdKbdpxmu85LevBXn7qI+qhA9IWO+fZWaq53Da6h4XWKKHjIAqO8rdHB0Rl+vykbM1q
g6Y3qwh4tuEMIWMcnkikQkuPjLYc0zfcalyYLeAAOUOuocad7grWNjf9dMlrafQ2s5ATbsWXes0A
rhXlklX/JSSOvu0OmUaH8HPc0d91idHUnz2zv5+bMhalbu1pGg2a+V/PWDu7Nb22HdjnTjAMx52R
A6CuT3CDe+I5mPhOLMR+L0nbfGEldjIpmWxvaiJeuITpX0liBPBr4HoWUbfHBwwoAc23ZuZwLDyW
m7W2BAWkVnzowVu8FarmLfYDnbAjHwrUdxJxmyJzrfs6sxPrsMGSwuRfODhMM2uiBlnXE+3+xkSN
wHirx6wuk7qFI1bmrCqQf4Mat1WAZPl+7NRdPP5HsFFBcSgxQW/v3M6AC0Kw6cZCgWsLoICFGwVV
PWKnbfpwRkHt6unPdsGJy4UISn0O175KeuNI4JsBcmz2iTT8mlqpzFHK0xQo6SDcRNflKVQ9fIVx
7UMNBlrMnF1dYLvvidL33keAnNICkNyMo+IqH1byQav8vf0xJgVVJRWkIWeM++bknqALqCw4O94E
cggUX3aM2KQgqyt2lHJnP9dDT8rU+EPZqdM6zzIT7sT4PiiNOgcYk81nlm1tGQnX1rP+Jtp8m2He
fOTQQ7rHnN2J0zYLdHdueip9Hz0q7HYGIcE3ZHO6x7tDQN8jyxXf+cHJVXXwZLWZ+EBWbd4yG5Fc
OMqZYy4ACajX+aq70/B/7corR0EiStn9u+fqsRxhH1Cwj6vxg5amsR8gLO/klWomT8VRS+zGa6bE
DBsSlaCrW4iDuC0BcL2cmFLnbr2XGVyg95k2stSBgbPjaik3Uhecvv8td1YeRWVqfungx/JxTotW
k9gB7cdKQh69+f2Ye6k7ezc0RvDb9eF2Xwvnmn08AhmxZ9qmUK23O+blXRO3HLjYBKJ4VUr7FEn7
1ERy2tKTyvKLJiYJ02CfFHRU8G2XJINdRzsxhUD0oUkjGaU0CnVtgQqZZgjTJB7b0DcMolHsBHRv
nzV3LlzO/G2I98h/6I3QHobsgFYTihn2kliwEIJuwqHcXSAZVAl/xeR7enflPYj+e4q3+ghc3lEt
naOTPII7bSHMNiJghur2cnyw1hIekjdGPWp0crL7WSf+4fGBFJ0902JINapd6oD6wiptqytZTIr2
tzJ/NQh7wldkNR4BAgSL2nK7VtooA2/6PfnDBGwQHjADppRIQx7kyduV6pfpw6ETjvo53cbXYQPj
f5OArClU8BF+N5lX3MD9tlImZ92t1vnqJeKMgT9A5s/yFSCH7UHSLIaf654EtOh0VlsKBH4wRkEX
gNbgc149eQqQXt+5U4q7YXYNWLd79V62QOMOls7fS5UFIuq43woVB1nXX3Cur3QKNbxqbJRBnWAr
uIyI/d7ReWdp0wperj69/r8dbVe6lEeC7HkeviQQtmzofu/xJEBfMj23ZPHvUdMDktF1l7vbDVab
PeF9yFD/yeTWskh4oncOT3QI7AtKvgjeCzJx2tZ7Zc74mhwLy+bR8lw1+P+GTsG1loFPgB/QozD2
xDC710R7JSeb97859qzASFN+XxzTcX8THTZf7WAuTBKXGDkq1xuDk8witkQEmgG4Acr/fHYvnr8m
1Z7MprvE8L7gPMAuOxW5msNgk+PqfVcKrDqIRL3m+BR/m97Ynux51w2G/lLU1N4Zjmm4xcM9EyOd
69MpaaTEPcFwCpTmP5fxtXwwq7L0H8ShyHAeRgZLhzt1GK+Fqfx2i9oHZsflR7X6Z4T0VXZRgU5Q
SFDwvZswyHtCv30BNwsU9piIvUNDuwcr5L7auo2Ym0dKC8eSts/HooiCK101GkJdCw3pQZF7SRKS
aOEHOd5KhvNyJrLDgca7n+5GKvLBMV7gvDhWa1QRObwf79Dy6LjVM/8KR0Fc+9NEgIRd+wycz4iy
Z1TI/Bo9j8ld6l7tnsvqZu/y4tLnMVFwiLIk3WctiJuQvnLGCfzgZ+1Aw61tPTb/ovc9pCvVulcJ
IarmeaCfNiZsJRdorMtARe49vWxizvNb8Rp0WI2ysqeC1IBoZ6d60RRW+0O1NTc+VE8ZIewPM2pT
pbG55gzvy4KzhMNerBrLRvydXQYb+rXj+gaTc8xIZCHefTYaR9UFdOahuYRRmXKQs60VF0W3KWQM
8aqzEMMnatlr+diu2TWDQDKuNClmz/Qx35Dm79ItKazJoCTpOS5BF2s88xj5zt45ZZUULw2lU71L
GOO5SFUEgyvMWdeWAf/4S1UFI+SCupj3xLCd2CZKoiTpdHtStTNDJnXZFany0VrhvH8JrI8WkGjs
GWgJylN6bsdBmGTqnzox73NbHJL5kYGN4nAzmgswZ6/gME03XPwPYgusdCvXTTGWXpDT4ypX8GLp
rqqvl6PQ7eEFd/GgZlSQ0z13ptpaLMju/AFmgkHWj5oqTFhFXr5oQARFNYUiBiMjfKaRy+qozMf/
XGFVe/kTfiXzLfl515qbApIt+K15E/GlDBsAcP1b5Ze5dDG9+OkUisaJEsEvfvcMkFonh0tt4wlw
W2F8VXgENNzBSJTGqcD/gQ0+0vGSlk+zDaBjPWgrfnnmZ96bJ32QtVytz/k8da4KoYOnPRG8f+xD
XZxcrsuu4OWPMldsBFDiwPtCgseh0vLGJ2+eIlZ4vvVcJQRez2RDUD73VRQgb+pjuC+g+MZxQxBu
Itw3cPPW4AsC3Kh4HSxSLewMGXfcxZNp/oeet2KpCJsZ2Q5nynbm6Md7OLTU5iktlriPgOHzNmJm
M1ybQiH9RG5cbwZ4SzE2GFDC5zhUX93hmdWgiRsw0BZoWI7oO7VBGlqYbGQwHlkRmzemZlUZJIWr
IiDgLepR2+IP9NzOFjLVE/Ob7qGJ/fEj4Jf3e05oCFCQ+C9f4niPz9vEJhnQvWabiI35MtBnLjFs
7V16D32KpH7Bd7G9+Ij0vBU5/DtvJlWZrz1axXIJdNdJEyC6OBWtSrh4S5f8BCEBTYihvCdfGQZt
mxFpRx/xWi8H2ebOquwOjxizpmQleekBjQ/aRHKLhJLnboFqy7UmktEfnw482RNDj8c6/o8W6yxC
B0JSrqYFOCOaD7Uc76bZScAiWryCEqTodirflhph6OC5YOOPjEqEZBhOzo2hgdg6D+rb6oofHq2Q
N1kY1mFNC0BWN9VIDBgjlLNgfQibusC1BV0MbsFCwNz3XYcW2nmK59XNr7//ftdcP+EfBfaKTWlS
zecLn03Myjva5FRTymUmHGRESR458IIqZsGWbUCayIHbC1g+Oimo693b0r5cAR6l73KDLl22/etw
TJ9NLBln5m8LPyu86PQtwGvB3eFXZDWJ9d9qL90nI/s9vF1/QZhCJCCuak9VK2jmQh9UpHW7+roM
LfVEJxaT09ZOmKkdA2xyJwnNiqWdoJhprA4ixKz7IFsLpzWCrRziA/UCPqPSnnmtyPboJG6VDFok
y/rjAwOA+pCOHhAkN7qAlsfywWbowRu37bARNHfX0QongYXLxgeFlU7ArFUy+4GsPZqLDmTaAEzI
lLbABK1/Kc8n2v40ElhghKbs+JOwZKzX3L0l7mF7bTZlfHbBd/sbqecYBY30E12yReNmYrcDHaJw
LylFZYFlaLj29anbDBAT/VwBPDAPUSWH84NdNWy4qstq3kFPA2lmsSp+drfY5ZGKLI1TEA7bOzCA
+TmM842SI3Aksj1a/UdLNqc4t/UfErCclsfD+D1enn0ZxlAf6eeD5xgx8c/fr+PNMLFI5RhpkSJf
DHEjKBiJcnxFlzQwgQ7sjFGkAqhKOWeF5CKFVHXZlDgg2NA1YPK8+gcULkWJCy1lHMdLFgnx5p0/
9V27+XhfM1D/jSq7QitaBZoTO4ANNwPXgPl4Y6RrNHRwbuaJTufRFPQl+nbiLPJjLpbq4H6sgqDJ
sfzcOxlCqZmEVfB5scRm2dTbguURnDfUlsF/aVxQKvoj1kFko2zHuUnDJxaKptZdAn0oO5sbjRl6
0Tq8jzfoJ3iF14TQGgYmjwWkmdTVfSR7Z3CZyzPIB0WWxxLFKOrZjVkBCIerSQ+yA425s2red2wi
2iwvEQ3hj+op6E7AQsEft2U7aBuqtt3pyS1n2Bw3gL1B6j3B7zVQVXgYCyfWcPMmLb5DrOL0pgSd
XBCWmAQ8SNDTfYZcj8Lsp6q9xRjlYbqNjew/hyJvsTnKg/y7EsIEe4XdKO8/mSkKfwjk2r27VIjb
dcxKcpS8F5ydyoIS/A4mquSQNdfaceTUhEHxeXz5yk9bbZekntJUSSw713FqJJge3SzaZ2QYmJF6
ExDwoG8vHfXZHCbyqHfc/kFxDgdQJcRb/9z7mKmlUDEzE/rairg+pTJnnNQMMVvHQZ6Q31id8S2H
2GGiaRumJIkAY0ctiYGk6R7wSU5OcySTFUUohser2jtJU+FCkukt2lHMHkOlJxY3uqA1Smu34QJ9
uY5M4asSK4I6BBsLniv7yFdc3Pd/6IcqK9UZR2F6xOqEKxrNbQ9SJGXE2jL48e0qN1S90W1rz2jU
C5HIoAIpAOCGSUaCN5ktyzzdyG6sOt2L77GsrJacnHBq1YXhv6Pn1jsYBcgEKsJFQe901S2r7DQd
N+BJ0ke99hRikpHuVHdJOp0lmG2Nb1joAR0XPZc3wQ3VrlTxNunrmW4Kuo0yh+j5FztUnezgnscV
zO5jeLTNq4Bd1Gv0ApJHGHMXsAtC+IBw3I0vzSWBURJq+LVAIXFBvAOstY8X0J0NiqGT5mZdF3vk
5vkB1o2KSJ1R86k6Gejm2aiQHk+j7CKq2KpZ6aTrCZE8XxaEt4EOe0h/KyzDRF+wjBLUfvFsjgNj
xyHxfCouOboPoShIyo+JAJj4AQX9Jzm8bDK2WLIIZpfBqHsCrn67daCqjR/0nBWu/O4SsEaAoRqV
rUeNmjgK5BTY53Gr7F9bE221QKZrWEq9TAvYdMCsdFqjKIVs6XqYQhq/vDsuqET1k8DfgcqzY+Kz
UUmHstE4iUbtvQUoZlt1B5w6OXU+jV2p952BrrWsPuWoaP68J0KUDZm68J/8bGKK3riqfMzrGLxu
Ew+sY1KlSCNcT9kQb9fpbaWlK71L2cZAOEyyaSH0BRRlCUyee5EOBNwTWprU0JwTA5iKgFbZlBTa
57VYGzMjOJ9uIPAXiytFf/Fdb6wdIEerYZJr44elTgK8eNGXofNl3iHh39ypGZf74y0pp4zVueW0
yrHeV9+6luQbgaqWdELFCKWPlRPBTAiJ89/q43t9qQ+6F3ou6kUkb5riPGer7hv8OTFbp2rNhBFJ
tIRAm6S1NBNqnAKcnQuyhvsXU6rGKCaCMj54tB0gL95gvSd/5mGm+M6DKeCozab6j2nktl19RpHK
rYeGnTB9/KhbN3yo1RaTlf2U/audEVDlUfS8A/B777v7CXnmUpADFD1FtLwtXoXhisKSP8xhWUeD
HqE48iv4DWKv5MdjfNi/5f2dQOAUpm/pem5muTo9oR0fUaO+Z4fjw0XpWk/KxTD53gs1NFV90k1a
b4vzrBEZz031Wnd7vDn/tZhfccc1Tqvh9KH3G0ZuTmIbrvxHSa1aBDe3tCiSuMvRwavR5/CamNXr
zZB0Hfod2f+5f8ZtaZ5PrAaurYSiUfzA6O4DqH/jKZTkhZbB+7frcRKuDlyB15i3LlNOKVFWQ4ow
fMlQG5I9DqSrsvmWdvmItQpCQpQsyFVkDWqSqU6nDgixqN3i2bgzAY/dawp7h1IWu+1RY33pA/gm
Fr6mg6ZiF5MmLN/LcxgRyoeSe61/Rk/t1jgy/tJO2lxoIJMEqk2VNifgqB01k4v2AWMslpXjfjkd
r6nWDvDuZV5PsOeMKYzooO8A8LEx33r+1Ph4yPPuUZIEhQtZSVyfnK5x6RYNaMe2WgAu+k9qgyks
R0uJzGq8mWMliOKw6aytqwt0Hz2iuBA1YBileXHNHS6byHAXgflRdp0fkkEekw+janQMixHitP0q
TQ76mmFz8gVSNwyVX1X0zSK8R5AZZkSaZAVfjmqNNcqmVou8skLuoKMayvW4S4PuHpO4Anj3PlC1
+Pv+IvcEv+yc58SiTTUKqxeAoknX/4lifopO0SLVQPqGjUpERB9d+XBGjOYNpz1u9fCDDgQg0X5Z
9P5J9cVlFCUbhc3UKpTGUwgd5mkoPWFjSpIF876F02u6QoIjvbxJJXPsVSrp8ObHkLXwdvILHdH6
EmjP8M3giUyYrU1fyTcC0dtw7bNSxuyJWWBhEcV6qp5dYkhs+K/4INY643INSACKqp9WQcdIh+Dy
/0fd4g4kh1gSTInth6tE3EwiILKhwHpNzeaMQkvsL8MlcwmqXbeV7UxOytaZdp8UXYaR5nc6V6yx
zRuAj5INVHYP4AouI4IMHH8wSPXMo4x1fZsh5CkUWpVUlPJLhfJ0kbDtjuqHWUU6mI+Ltq/s8Oqb
yhT0RcTYM43fHNv7GYwCN2vfEbdEAqXnnLZct48zDd4bdVsMJA/P5m9AgaZp4YdNp2wWwBzbYNT8
Bd74C5b7jj6/fUUAYoqA5Xyli3g4pSR8JyVnjL12QSn7/EUQv10JkaOhgwnY5GelS3fUo8FqhSBE
GkmWX8QlkhDNh4RECwMLi+W0KGA9YVYXPHL9KQW23SZ/gsNw8C+ER3BEsrtKSXTj+gGmIzog3b1N
tXXLNJEzhTsLWu7GHK8L2ukl2wxLtv1Lveg4nhpzpBw6AJ9daTKHwSELqOOU7weSzLajdA2bOJv4
EwD0mFjzlIkHMUt81tvSNwjp0QECq2RhLxg2KbaVdEEKXqBsP7QxomYGVL/iOtU/P/UP9wqxEMtO
edcp5GMS07EIQv4oIBSWPvPBwSjWiIckE8byrWmU1adXkr34WZ6uFYsZ9CogoobWvL015u5DbowN
NBU8i19LIv3mKDoVJI+YNSOg7io0mUmkJtRRdDwsPQbZS1STNQLmlzJ5IeJ9FSsk2JeeKS4BFCqR
thQqAFpEKXUPavZipf4EXSuH+OFQQAIpza0CtdMYbRAlEnBgPCsXjNUG17GTf27WiEkrRnBYuAsV
uu6wTEUzxfLlK1SD07plvDUoZbT/lD2L6OQyjvE8G4CCzuUPAMxVDsGiLlxYHBTDBxsBIxIyVcXy
yhDa90UMcy69GScAze8dRrcuAHKWx+rvz58fMEFYfyHTdrefoHQgtOe8PvuwOgSGjxa4lx3gRiW/
12r5yN8fZ0JSUVhl4S56FxPfUdonyoKUG26gC+13iISPOb43eIZLV16IuF88VoFCCUhAItCh9SI0
T5mb5E0O75tke6cqBlJpk9JmVo+BLjk0RpwpdoJiqlxs25cmEZ9iE+wv5pl90vB8iF+H+J2EjmES
H6x1GBdwKbG/z2KNBgtn0aLF1wRaDJr5yW6cDSn3Pbp7iK1mgb424SITANQiN5N1EAhZ08Pj4gf+
VGldOU6Q0Iem7wIkUfRgcGZYuS3J6CieUlSUZ/Hu8/VbWSGJzSqD4Q5HBKeWiYTdNv+8ufPXzPmy
tnYVsgzZBQm67fHPUtHUdPt+FW2A99bT6mv5U7Z4RKNe0TmrnMeqfN8flJrveaL0c6yoB3v9Np6O
LM9bbatqvd1rcxS3wLyFxeKSxETbJ/xle3q9g74wiu6sLP9PYvU5bFTbvsUn9/g1FiYxZ298PT1x
EpVWm4uLhGy8M//xTGM1lqkNCCPoO1tvq/+V3r8q5sZaOj7f7E5MhCuH7ma5zLgTz1oEaqrGOPL8
K8EM6kJSVGg7ZAVYEqeBAynfXC/H4z+c0XQRANckbbVHpPLOS1CAT0kYrLrzhrWNVQAu2yOMQnhb
yFUTahqaGI/PwVT14MoZSXfrerFUUv/wk8VhanYI8IS9EYYi01QfF3qNHwbyYWVATbtYePOd+2h/
o4R27zVLJQJRr884B8xZET6kb1P71uhwpBvePKJQm35gF/BpoShBcIBTzPLy5AlobCchHDdsNCEF
IOw3op6C8EFAqPGelwsN+R2BetuStUkhfklc9o4siZ5xKQvYv/ygiTRtrfM8vMD2DZPCzFHRnudr
dhLx7p7bHoAc2clUwTYr/gzmffDrCIt0z1ASBOERPNYRyzv9kgj1U5p/Jm9QooZhSL9SOe5lLsYy
iGE+G2qSW6mtxiMs/5QZn4fGjXYgua+19VuQ8oGFDXrIcqHHA/8eNVKn/THwRDWFSwXD7grt1dQq
3vJJ6ZTCQ646K4R8JxM6j6A8RBwG0u2REMEpRXeDowW9J3qOk30cEJAcrmKB6T2wu/x75484/u1r
Emb5KedcxG9ORwIhyPbVTg3UBu0AxVO2UGOlwTHPbjiY6bWRPN6I6rzSd7PuC0QEraySzQjj8DgP
knnSQNGnc2HpgZAECzOXdM6zzG+r+loHjicJFbb0ecVLOgMtStRh7dt80EIIuyvj8oW/Rwb6OyUa
nRGjxGKuo1uqUXYVPI7HYg1lsjKKrpvSYxmWLyuOSKpJncQ3TJzxleFW++/ENZ4agrBKhJEDnpmw
TlrpHb3IkS8DGlX0ttoE0rGmm0LqcMU16sbJtGILxsU6rjAIYYcjAINY+ulouUFdKcbkyZEDgIiD
hAZf47DSobEMXDr5OIOck4Smd0rgr69qE1lLgsBRU38gWAMncbfMNDmkZLzE6LI6/s9npWQCf4YU
BWHQM6PxnkAovDxQKhCnNSuikix7YSQyRI4Ljmjia6PtTO9XodZIL26nUmW/0mR9oRA5KvP+dHTc
Y9+iGrwyVdA9Kcf64vw6UIM22KsUpIvkZAmvANVlK8lX+AmNcwRNpdcLu9WlHphKEx1Mnq4jf5Ji
P/NPGLVIeJV83KWq5pTHSC4nMw/5nRzcuo/nShx8xRbMn7I4YzEj6/NYJCGLyidsyMrlALXEpTkx
MHtiaYDjtjPPpiFVaJSKzIpt2zmGvWkjWyhPhTsS5uzpB15kY2gcYWrKK4KL+o0YZDytipO/evuR
tWNfQYmobNxTU9D8jiWQYZginxcCefxplmK0xXqBvILmHuVrLAxFCMuw68+zCwoYmFl65tz8oNx8
xp/yt7avJx3B6PLi4KElQ7xFGeOE9/l6yjXHLdoFPBHiFw4LwF/TOBzzq2LnWZ6P4aPz3Qzev2Yp
pglCnEi4j71cOeUgkHLBoj7O48sX9/FS3u4a0GSlf6SHhhTFk9Sx1/hQVWbpfF2EtbWTFgiuGaim
ocxCjtz5wY/Fh1w+55ldvPwP61hm9Pyxv2s5gWxtF9p8aX83dJe5m3FzSk+7eyoN7DGoQYsZxrvX
q6/pYxFNGkhYZSY1k2T/N1ml7cX28Vmnji9j9HX8x0Q/yC69dauKn4egLySujQBoBYLcZ5uKn238
6J88dzlxt8c0FNkZ2vgdLLbzaLi25KNitQ8iXdpGTsJiZO1CdAhJysly0GQkEaaBur7rNmdecNJE
KeGJQb/fTazfE8rLyYlYRjGM4doY33rVDTEOksahIB8xat07G6vtDtBbOaVt3bPqtkftESHjZANT
x48vhVXB1QNdBPuAg7rMQ0MkfBAHTsV6Mf/A+l5HMShYkQL8hvm2AfklA24kJ7Uss6+ufOC60WDj
5tM48MjhHFJrrAN8IlRe/W2ojBipk7Qwby0bgOy9GKTH0iif3gbRFUHL+gXuPDBeqAesnhvLdKVJ
VyX03kHCRigysn38e+3lLXMOXfYWylxUzAUKLUyH9wmDd80xRfrYNPwF6mhqLgPvzxc6d7EPa+Wq
AxBdndQKd04P8iIngyOA4NR8FyebYhJcnntpaL+ZmxuIuwrmM+N3vXszYGZx0fwxlg8O3TFhFFhV
Y+/sRAWAEiPnh1gyb/O7qTUonRVOcQD+nCziq5k8D6N1LVw6Lp2BLa5EAaQEoX0NnQ3gR0lBcDtx
yz8JXWo5/P9uWp2ewnSb+wbL9tFuiG0Ayj8XujYkaNdBJyFZp4AGSwn8O0snTxktxWMAGIux+BHT
KfPnwiMmYYIwg0h8t3bWEfu5QzYiMbDdK0s4jKNCAfOjBOs25rPHy7oVJQlEAEHBrc88Xh8bf4HI
/60n5JyoAToV7mTz+7Fw78cOhLURXwqV3TOoEGDbobjL7tOHDaPxSM1/OIqPc4iyskAOy+D7fGLa
tbuqjVhkv02DoGumo6zxEoIWRi/c6y3/XRCbPXFubvsIp2qLtgUWoO3L547We0bpXOf+zNq00fPM
nWifwOF2bNtuSeccLp0dZ5JtHG2IEEaTRb6GpG8PF6f9uDv7NnYI0zWFXr8FsZw20aD39KoDct0q
jD3TvROMNfy4Eeb12aP7BICN56uWTFBGnx8GDnpvsSYsCw63hLvJK+X2QVDUnqdpg7cB7a5Xoux/
i0PBTFzfmsdolZqMDwKPYPhsAMtpQ0ONZhJVcpPOSMW0k5RclsrGdqHVcUDtlWQspkEw+vWKIEXq
S7y7kBRg9M+48zRJaEflXmqKS7aYUaF44n93hfokTRGEJctaa1LgCb1PgRy31An+TOZ288Ty6QwR
C4p4ffXd4Yt+qr5k1fUKP4Vm7rwXqmA2PwXdxnsEG57+nYztcGsd73GGErq6yr+2dDUfqf7OmC3m
ZzLdIJHsGc8QnSbPUSbvT3KOLJ6HO5WqaTrdhkLC3F4R16YrD4onHWUp3r5OZoKAJENPgM5sVjmt
3a5RukbFDzDH8PGpZTI/zIPx0fwp81c7/WPhTFltf2DvY8qplPxSnM4S2SKOCGGryXjX5lJMhXF0
f4fPljXEW0VvKlm6dwPQp0pvt2HKLLsjjdexWOeZoEAkv9Tf4Y526on7KHoSSIIvKuoUkw24+qhB
auA7Im1kraI8/re2sqN5lKhLWdx0YomwEbfGjrGNpnRPoqISg0dyhHjjq4nW3p5xycETE3GDVh2f
0fTSq6HoKGDU9G8WdwWPsnKofk4qjIH0OPGXxBzGCtQVn22xdMjibcfV8Pe0h8EnSCpkyOqr7sw4
j7H/Fu82iJNZue7+fRy2VT4mii8pmypv/A07SEmbHaAGZs+JTL8y46Xb05fMcImwQphoQhu6/kRz
U3aIb17Dux6Wu3zcOdmt1YdQUlnUtNn9ZhHx+GeIewuVmAK7zLdvy/F7J2LH578VUrA54xXZc0MZ
2dAEPryFdw+ssNU5Xu72IWhldu8AEWSTHxXJ8v60/t448mIVXaW2dUXFLKqLXI6BgiSPNp3Anxg0
xdRu8+Jjp+NKdZ19zN0EACI/gBJbQRxzPoMbaFuGD5eKjP6FSXUW1WcOrgJeoVEfYT0EpPmn6rVV
92Vr+STv1OX2iHGHiCFwT8auU9ag5/aW7dlUo2U3M2DUuTMPUFKi1ISdbkxZIk5/SECLj3uzaIkG
puz7bqOcQE1oU2x9EdkRR/F/jwb8CeTbk7Hf8Qlui8cASYSP5cAFJAdVSgr4qSQBjNzDL9+UEuQc
cooD07hZ6qhh3BqfMjYKA4FTW/ijthdsyr4iOgxRLY3/cCtkaHQNFJKB5VcfK30zNjKya8bONx5j
BHVTO37885LpZHv876/0/AbtDfo+tKfnlsWFYHClovEHkocoWi7TPQCS0Kwlv+q1C2pX4oXdaskn
072k4B2W0Nc8Kp/iHGsijQGDZ4nPeVEPim0v1zThbFNEPtTvFhb4suOEPIYvXd3AY0uo2DxVSeT2
LjtQmp3QKEK5ADboJcOn9QPTgaElVNqoLoDA45ASntu0GwHDXCvbiHNq2FNJ8RyrJkIevz7FER25
3tg2N5C4F8oxDFM96KU6anTpdLDgxGNAQHfcCE4lUliY/7qiPm28pTVjU+KdBd/taDk4cz89qOeV
J2yKL8GmkuPdnWoxa7IUoS6RCdvTMZIXkS6jqppUF+wnkVybhzkNMQZt8Nu4ucspDMXMoBQcj33O
AzZKGWvm9ggu+nOx0IaN//EL51e12zdCgr+xBJYAQJvaofekzD4KO2Sj1D5Coe6/TCatFj+C7LCB
s3FL24e0DoXYIhBg/9Nb/sKcoQiiL1lNjs2N/rP7+ro/8i7dWWwfP3LagUcy6SntUmU1wHvHgEx9
LFRa+iXdhEXtMgIbAnR4Vsm27uejBBzVosr8dN5J/1Nn4qjjoTDm64tGU8fmg1xpnG9MUMboINAg
eje0QRcwv81px94LsUY4nHBxFSv/LWe7ysaPmQfAIPy7cnYu993uNT5KInaYoR9grkGE8F2Kcu14
Yhz0mESRw/PyvB6cmNo4ECVPU/4LVAQIe6jmiP7rV4eWNJj7zhVMT6GnJjml+l6p9h8BlGplZBvW
xju3WJF201yCHlJaXEHKLkQzwW5Ydcj3ExNKQnfMkWKs7aMGfTSF5AX9DKo+hehj1l9QYrU1Opl4
kn+LfE3qOV5fqBFOWEQB4LQRjot/kiWC65hjteFNVBloTdO//thk5iXWvyqzN20T0x0iFdi/5xOx
XE/ADAC4rhaKO1iAssnNcH1mBAf/W5xSVRFmW1TIO7WDzEQM2KeMWYlT3sR5+D0mjH5tCaFUhm/7
e+8ioHKF+pB6u3hNlU+LHpamrI6vDDUE4fVlJybxrvig13HiNaKuTyBhtzpu+/H5oViImfiBFi9o
89CZfdfOXqEM8s/TatT/lfEhKRixAkR4nKopqhRODcgkwa3cUJpncdmvKcHaDNy0HATwqVjiDkIS
aErKJ/QMq0uHjdfe6s7P+AC7SwaBloYD08XFHWCmxjf7KmtTJH4QEBaEtoJYt/zoIfF8z/hEd34E
VlTwJdiE62Xf+ulOb79MwVs9W9ERDD3CWomR+A7BQ0/H+OiPmDruYnFLCkyeGoQGgAXD2Yc8nfkR
2jEcKqiEcdTMzkypkkHv0+/a1s0U3nowra0Pht4qXEDrkNoafvQKCWvohv2czbqGIeksC4nv3pVl
7NUyWg1zFII9ITNAM9G3h1JdMGNFDqhXgKu5lpAQ8ldnxPAYZmCUxliJr/3jI8ssuIPUqAA508KB
K6n2TaDvQbT84X/CmBSC/wXjB0DROyJy2Eb1MNHvfIgVtSlE8g7CILYdX+5vo3ld0zcpJv58/dl1
jKWPXMFhmv6mOQHj5ZmZpeZ7tMw5VSuEHnKuMhsoohntPKUlMi67LHX7qADRdcw5+2G9apNoiNNI
/29fRRjcKZms1X6i2rVrDzXMZ7M35QTf4YzWTcAG7mg1mIPsLLYl7o7KN1mRf3Q1nev9TIO/Ifzs
zW9NFKr+alaZRE8qfzWnD62BYaB+J5rvaEYi+wz1HoTkQpPxWtDoDjH0dcd4jirWIopkwlEUa8/+
EXqfzz9FIG3lUTsNkPiI0bwDQGG5F2tmZnJmpwP6DVLI5N9brGzGIW6aLVSviRSImwSO/8O5CaH2
709B9pHZ9HBvXXkOgKf3MVAiNuqIejFkx/BMisUwgcpbdqwY6bvmHCjDwQV5M6fwk43ov0N00EU0
f/aoSETyMNAYKsSv5V58FNKDsNLKt+ffscKtwjM/YnMn5StUztTu26dTT/Y3MfdkEzEthPJxvvKh
oA+oMWwdBmITn+A6x87jbG3pZSUBF7i5YdVYHwJdYNQRVzjYQ7ahhOWGqvVGJwmXLoZbSBh0IcvO
1k9jIulgyhyjuosMFXbb11UQA1lPwfT92ChiKQODZ1D+lKAJlGgeVxW+0w5PElnCETzSqv2hHfPN
FVCQ/dtlWv92WS+/dIcQL3D4N5PXU9KFE/QF2PZGVxCLOTP0oQIW+jWpOx2PHq5U3fiiosOx08xB
IRHy1IKwHxq5scTL5iNZvWzX7pv4EG9o7BPogg4e/7xK6MkXQLv3wCvxNfOQ/th1+dXs8OxQXrGY
M3Mph6hMG/S5pNlBV1pp9YC2wYwDL9VTuvxrY1dRuk0iL0iwB5Gz3IZDECnQucyT7oOyQjvV2795
/4WgbB5nrze5iLxIjVnr+Olae9x9R2pKf9eb1ViZZbje8UGW4dER8iP1624oEUJvzDJJmRY/IBP5
TA4o8TWDMd6tn1UeKGeNfyO7c1wKSXw4Qe+KQNOQYknlkz6q5Dij4Pg5e5YQxdKHmOb5w4POYsDZ
PY2LVzXFO5d5lQF5lCATvklfrEC+NblD5KPnpywcq61wf9NsaxpLlEizDnN9p4twfxFUKLNzG8uA
fqn1FDZq0OXZ/W6vq6X1AXYwq82s9ZnLdp79V5NP4IIUtKCxMhcthPChajmgXEkNc4UmmBYXQjvO
Ej6PG81J6AbXnpDKdhaskEqfibYqIRfuzKRiF29IS9nLNqHJST2eKeOzAv+rp/dsz5K2MZ4ldmZX
7lWfmuDjnP3kz4NaaoE2j5D2IVXaPIQmd8bE9HQpu2tBn5zd9UoeqPeij7SXbo2g/hgH2iluDIk0
68chu+nZBnjmL792MsL7LizPToB/jI6mwVvyVXkPznirpQmFnW1Y7/zA1Fmvm8YWhQ2Y9JOEgans
688X7UW/blXLxDOH6DePIBGq0D45QRLzhjDUOi3+C0Kx8BT1D08ZtqhQrke4SEN0A8/b8vUkThnS
PF0kHa0ysKlACEnyu4cqFsiVN19ZNcz6xObCyYly+eIvj+Wtq88/L4vCsAA1ew3JwhfcLMrhGJQx
9Jge0Y3WrxKfVodET16wrfiR0oGFdEWbf57Rbu66R9kh5lFzZZyRyBbFN42uK+nZsLMrmnhGCsNx
QuUp3IJPmx5vKn854H7lWJ4NNQUEn7+4buqQqSKpIFjXunFex1teM9rDpBo3y18DqZ7Xxo6ohcTo
emzkrJLIP7iiaJNX3LRPIuicOgVvMDBRvaDdINsrSxaIHVGfzrsNAYpFuqWuJn9qgUNuWDaubamD
L0J7TNSDT777IAWAkj5NRysLv55/cyofO/jjbquqjm+cfTBXgmMNPklbgddeutGySOj2rx/e5Prs
35/EClErviwpsLdIw801aUTkyQ7gqmHS5cbqRAWiitXP24+lFl0BUiY/S9XEfVYEbFLH91CkyNej
sn9s3O971swcQ57n49XyHuEdeeR1AfcErDoMYHGwlkKw2zVLSnUEjDbd5JssQsyYufNa2LSF9Ww6
HzeOhj22cWkaJV9koF867HE+euUiCo/ukKfRTOHil8O7V3do8++sChYAbWiJz/TZlXoCbwxaFDWQ
UjR1JFeJmAHqapl8nXswAO2UirnUXdRPI1au9eu4kgAsWhOSMXqu44JPYpaZ8cgZ8itcQaJywn7K
y3yvVSYH8tQDn3+Hk30uUJy/bzs5OlLUxIdUs83iihkrQPmJfRyb1OUT4Lq70ne35V1y9WkV8Ii8
cDj2SJAEr+FNJnY6fy5VnX7hUB1ArWps1Wn/H9aTK6TzMnf7FqqhF0MS3SGaiqYrT2WsY5KEUXHX
1ptJaHwa+iSwrYIaYLE/SwCV8F03TnUos8psFfoL9Kyh1BkuVPcQ20duJ2chH+nAzy+jPanqYkS8
fgPhWWUOxfxC8w7Pf3Qw/AW+ou5GUuJXvjJwVt+maSMF5RU0uBm1lZsgKXSqkd/+Eh9MKRq6pj4L
FPdp+D8ZrRPTg6/OXDG/zQwAPsuIUmfxiQ9FM/ASGGDDJYZNF3wRXDAU+I1FJ0aPP46/OliuZluK
GrwlTW5uXAURJYOUGyMI2fKRzrn81fK/tuuyErNqB9cPmfkGKmMq2G0+jJzToqjhPSP5pXpk97Ci
N65Oy4mK868N/TKGKJgtzauSLSj8RECPoIYdK2Rf1FWO282dkHy1J+oAowRstK7/atHArvU0DUlq
ww+gqZIH+xute9LAVMoNB96U8PPzhlMZvjTkIvSPurDlTo3gQnEAoI2xk2oFENSNEfCmBd8l4kxu
7pG2VdgsSBmqQWKqNUspHWso0sgURZktGSTfrf42ClfuPjcanXLEpCjhqfbz5btmQiRpBuGxhKBx
k0yvHC1XzXsHSKWeLPoydM6h9fajik2/ooUGjx1RfQe41je2SQjMk11xoB2ZtS9t0/nd62ibsufF
a7/AZ38tMmlrGugBMKagYYAfJkBi9PJ6WRQ3adJslCDKvBi16VQkfePFA3XmUJMqGsxI3TuKeOwc
Q6O1kYx2Uly1GOZwwR4y0FKDwgVofZWlQqXzE4KmyKg45B1XndD1lgvznRxFfIOkblU4vBAfNgDs
07gUQSVPr9zGT7chbq69o8xySal/fCMhgMNfd8Kc6sY/OLF77po8E/Q2z5CDDi53N4OrZFzOXhCx
+mtfqBsBEv794UNAcWYvUsNZzRmsOMLhcdxrB2gbQhQ3RrePug5zIwUOIQ69Cx+NoAXMXSgSkT/1
wU/A9dHZiMFetJZYeLb3cSwGEiO71qCbcvyUt3JMuGz9ZuurBnt1JvlCZYfW1AO3J+CX2Hefvo0z
pLuory0AVrorhYzZUIyPh6fYpscmSla0dZfTW/xpFuAOx1ncJX0aobIIPEd+Zi1truG1H7K9+Pnx
5XTAorAX/SQhmFViNxYonUzy+Qwe5eKGWle3yER42tuuuECiwfugubBrO+c+MmKNDOAjUQSyYIuM
AyVgrhPuq5BDZvIbfbJS2ktfjx7wTkKhntdoAGLH3LlpVfFkUfcr6E+ox40F4HQ+iW7bmwOMjhYo
DAYgKZ1sI3faFfSVISDDr9ViYsDpk5XUKR+OVKTcT40jid4g9/iQSY5xbg+eskjA1KgwGf0DLfOI
Iao1m9Qyc4qMvsaJ2/pBPjU20jkv3MJ6KryEbwDzlpO8U1HU6fBNmiDzQgXuW6YmutiJ5UujedEa
Rg8d+TbNC67NCLown9M/5TiagmMxWwTZGQRilpAVUhB/t9epA8Ua0E6H3fSs3p52hvps9qcrSTym
f7ubFkrTVIJC2Cw0c8SeFz7+r1Et2SVU1+jXuPyqR8tEqZYgB28Mew0IBHUh96GV8voOyD6ekot4
/HNBRlONJcquuI6O7XMEkWOvcjS+Dgxs/e6cyp/8BvmQtx0RNf/s2hiLiAy/74odGxPv8+7ztGh1
N+bpHB9KBBkfaaURk0EEGxGT/1weR/26eiOLSj4aR8nS3NEvw7el3XyUboS6uV5KWDX2IMgZY1fe
LZOHWpWdUtAD7Vwmjo83jT2AqD1fGTnkt0xlFKCsuXJtemclA/8fRjC7k5x0GNhJYXpRuLPNPm92
jiOfY3Tb6O0ING3RoAMfc3aGhzkWuAOCMhSUBf3mnppmF9EyGprszvcEi0nC6To23x0VPFU54M+S
edQWRLD9wHmWIMw3B5p/t4QUglr5yBeua55QXJYIXljtRQXZEoiYEJ4bLcK0fOJhVoVsNpdPse6n
7v5hx3dj0lAZXi+QHRIjA/kZ5gK9tExNJM3ev/Gac2lXtb2uyhmuAF17DxLOsJtqt5maeXmbEWK+
pcA6TuHWVJ0BaSk0yaxI7u4tars7ql6x0D9IrsTFlXoM0taSpQHaptc1nUWJH/660SoBzU5oLczP
LpAErMmnqfxe438WRqIjhxYK8WVz+za7Gp6d+S7kxXmoUn/0xUFs1yz/aBWisHTeE+3WUvw+Jpky
gVaBC6dGWtX0i1caidD8jzjxNlM3Fp1E6fnwVyKect2lFlVNLlHRHV4/aKgba0FJh6lKwWnH4321
VDWNLDYyXt01pv6IdTe+16rL3tQzvUwHSuwg9iBwKkKlJNNPWp+Z2gL1/XTF0+t71WQ6UBFZ4ssp
TEzbxQ2J+g32TeXr03XtQwZ2GQyxs+r3MOIWUW4CR80jJ9s7V1JoRIPn5MaGjkLEHTQiwAdqweOI
jQaJMZTwymlV9qz+ABxpzRjDJHh7v1uvmTGqITiRAQG1BjaJNFY16xQ/cHqQuuh8FDopdnrPFqSg
IyJy8vCouc7+kPEV+wB8zMFGkY3B01v206K/WN1VGWo9bZnVrTgypOGaQspiG6CYgtDefPs4S2xb
shx+YLRQBRC30jGv2Al+Eez40U0XilK4fHA1hMWyyZeUdhhG9eMZoQ2zGlvJwC9nZhoDN1XBMHVZ
AykSz4s91oQoICLDl4HEoPRwWHZGXHK00Iwd8IqyBZOw0VAuHfYWNmpRIJnQdQRxC5drmargcyn8
LJmyfpRZi4I5dCiUNB3AomuvgxeOJcAwXV+wX9lDYntSmCT23jhWInbptfsc8UJ4wyE5W9kha0Y0
STAgtXtoPcN2nVfL+2S9xxpyPzfcDCeLAkUO71LS9ZBp6BrcYA0DyYrNI50oRrdb7e7/Y+Vw7G/E
X9kDJh3ikEwZjH5d01wAGxi++0jlSH0P03nMsEhxDbVhng0QVyRWWjiorK2oJAaeklrvRfKovW4W
UjgCbSw5Axpf3QN3wEfNxCz08iHXPqR9iqAcZu8RLKZz9cVKBEFo6DnI1/H28hGKGLoafeb1mTAg
PIr/C1S2MpQdNyGvsIaq4uI4NJKfIDl7rFWL2PqMlcxUtObOIVpTRHxoo7+c/S5l/EOoxods5nC7
iQ0u1CRHHPpkAFLOJRslStpsfK/mLPc/ZATQy8VnSERJmfFDV2w0OVFjBCWbVyT0s7vB9+KaCtmC
8TIlPqpUBel0n6t9gJoVvuicwiAKMVQcid9F0C9RyiqSw1+2YCLprppckQzxdSlyt1Bi9NRcOCPE
bOLkC55B0h0JDPaD93lmE/lIkn8JUG7ObVVdB5nF4K0pVNVdEV2Rgu7w3FuOxCrg6qafkjWTjsv2
DdiZFCRpXOEPMH9zH7jXttc2FdPsQbaA+D3v9QoUhSbwTVg+RCvnO4frB/v3tA9QjdYjNxmWIFS0
I0whzDx5/Cgg2oE2Th4/5m+vR+WKN4fW3RaWQnpmHVJSzeWehzPNx+rMMlVpq1SYC1M8j4Xn7t//
jtN4Le9swq2iwduk5aIBtp8+DjXYj1YET3gi2xofWDYfu4UzdkfPjQ1nlfByKTflzCyPumP0PLYI
RzCT69gvBelI8qq0U/g0hcazZpKmP8u5MbIzghW02Dq4TjOWv0LzYmAVp30qcfnbyX6zmY7v8lgX
ZCSViTuSxR7WUXoxgma8gO7cmX6T7Yo+8I9s+JEwWT4lmulrq6GgVGNBGllI4dSNGtbRVJHqCGNp
0Z69lQ+7U/hfiMeXz/F3FQkzbuB1/rSJgWHUq4Jx24KS5gXwy1aDT8gA2uPXCiBY63g22v41G50n
0QdE7/mH/tmzHRtp0Gp6beGD3Ana3RqqsFQl1VpMl1JIffPC3arIQ/u4Zrngzt6uFz62xHRezgdd
ZcfrxcQRsxXdp7xAyH17l9JCZvzXRXzzhA6sSkzqQzKrbOuIHWxxQMMS+xaQH6IF/yPAKfrBeyws
ax+emJloNFE+d7/WQyQqqGTdFzNHryZF33AnvbMT/jZ9WhQr5gePu53tcn36dDwcIxfh+rF+BS3o
AHyUvvnHknSBaNs8oYeNgeHSZnp8G1OTnCOqd9Wcd8ohtHylhLT8JMPpF6oHI7KScQWzD577n1gw
uYB+49vkUd58r79D/R6hr8zSuT5kCkMFZyGnTUpxkdrgtZhVdgYzibRNCSSHrE7IEJMJWqexg5bS
tlMn1NkeaP4/iWUqwjISlqhs9TTI9kzcQiQtHrrMqZwR5o0Sp6+2eiTqgra536ifY4DTkeyXdrXl
MEBn3uKJbjesA+oZ0jtVFEyAHZI13Dvhq8YCNt3kduCxi38MTHC0MIrUGpNw5BFVxJiKqQX86kz1
jcO/Tz1X8nr0W5zAfWHgCiNOVg6ZzD+ZGgVvHgovpxDilb2PRWCYsn+9fGzHw41Xy5vrccNbDvMx
5I6Jz7yU7FiwHahbKkCpBS03tYNhi530SSsxIgs3BOJZnSIzSMDVZfa3oCWQYwmVRx29vOiaAYem
eX4k+gU6FeWlWd+WZZfUKIjefJV6vGDOqkfZxBK1sP+LGLtop2/gRmrxYc8vI0jvm4jY1LMddvIB
g6Z7nZkG1I5XpsG5zXOz1yJHTcrlyTppbGBtuojy99Uh1OPa9odlySQuw6i5AOqmj/JlEduocTrR
HIy2SoThW7ndjuJanQpF/QildE4i27Tp669kHNAA/vFra3V2vaNWazWb/eOkrGiEgImtsKTA3I1m
sj45l8qxA6cP4IhpBXL5y7dnD0X4YcZ6O69IX4xfIrT/zOazNi2ms5FQTcS46twUvwTUOHJkxGxw
cxopWwE1GGXbsQX5aKvWAomWgRu3DSE3nepke1aLdFTmH22EMJ4sEkyYZV/ryC2hUbcjDMCmOTnp
gIOT3/e86WNopsbRkMEY2pbEnoXJzr1bBBTi1PZDqeyhaFGqWFl4j1NxX4e0Y+fjFOTkL3bJyYXv
b1FDxuHHKBMfnrrDljavYJvA8TS2EcPNs8gaDYh+5WO4UgtcnWvIrMmSOGGgJrh23zPVKsA7kplz
kbloCnr4NY3tSCrVYfTO/TXE/yUYzChZRqcTTnZThPgnLaGHM0W2lsqYLv9BYB/JMX3pb9B/iFjI
pjAKCVAJOk7+NqEA3mVWecF7r3kDMxMi3iCt5G0pZNs1kUK6Jqp5um/k/BGGmYd0DOyXbPe/NeJy
qdOg2tPy3HHxfJzKuTx85vYDc123DpA0u/Uq1c+xjjS6RKCz12IJMPLbikSSxJVxdjKFrthgj2e8
FIm0cV+nCRNYNdHVpbkBMs9+nkHwrDXpQbJi4TSXWZJhn6hVni6RBGnqvIYeE2Yy0loqe/F3ZrEE
buqYor9lQeuN9PLu5V+FboYoG8CdruYPNJ9KJ/XrdEnLgzJ/4vkpk+Z2CqAXuC7Gw95hbEYDqj5+
OmvHjySUPLgJwGM2vpAM7NYJbi7C+7X5JiMBQ7U8ZfM/ivBuUFNr6LOcxljdGHpPi7oORDcIFGn1
3BxE4qv90y8Zw6JDfm4HUFAWoF0u128vVlIwX95cokk+JR4S2dGSSZIUTtQaVfPju44bK3AHtwB/
rLqN3xjOXZ7jTjDShxgTKzb5HMbfZ+/16N2QTcXNdXsyoGzU2GEVRn4mxit1LDVDSaQXAerCY9xM
odT65ADCZPvyPChqdzVXgr/R8E8r2Vbtl45XTkdqdCXylhNoCMxFJAE7d+X5fvmztF1+C1rKhS+7
5SfA6RcUsuXV7r+5BpA97b5RJoWdmct52t0yq5H2V2N7qpgl8v9qkltlXhl5X7dX9Uy2HLElsYyT
4KXtCe+rfQ6QqyNPf1gsIKOr6d+Ou2IpRfiFujp/dcLMnRofHpEpjvHMu5ixjIIp1gsm0WDigF26
JA9r5mWoAe5+3dERavxEnT2ZMRz+btYjHyv+4wTDihsB3VJveVzYzXQlfPm2wWzHYh2kQhRrdTxk
KcJF5AWVESA8CqJL2hAhjvJu9ZGRJc6/Gg7X93K99p5As0EDZkddjHkX6gHw1CEIjhTH6WlvtR0b
G7GghPluTAZsunhxmNFGdkd/caTk3TuKqA0+73ZicFGKuuLxwkCn7M+u5ArBPcXsDTZjSt0Kz5uA
5jsYH8XN7gJr21XPkBssLywigj3Xjq4TaWGv0erwOOKRWYchXHsGwqjiuJcBIM/SLJxpuqWUHg9J
CBNj63ruycquJDBnpaZAuuqPGCmhkzsb5NybcOQE+obr8Pqw5iVBMhRZkCjmc3C7kDpRT6okkAfW
OKsxdx0jxXbXX55Dheps79PscBWar67q/KIcYGp/S3WHyLGVesVNpdToFgGJw3piJeg8s7yGyxzw
JQ5pUNdo8OFUcf+oEJ3QaHjs+5JlaazXOat+lH3Zdj1s3DWVhBc+Hr2cDlu47rtVj54OppnH6AKy
mfwbGw7sTF4gkbILk5ejvDjuYPMax5mcxXpe7GZDY/D8wWSPnO8C+ITovps+CRdSO1pT2gqAKuiB
R+06LAgWEWgNyWWDH0JPOg8Ke2bjuMYx0Q/p3HBTD/CeS2c+yERKRnPlori1BEuW/jikwrWvqwEv
mrfY5/DfJG4eRJivrVXMeS0B8FZQw+jmyPS+XxknXlnvX2DdvOlSXRi+1kDnrYyACZgsOwa+ZQs0
eDiCkhv/wgA7y4xyIduIGFpjuJYHLgTaC8dx3Yc93MyzEfiufjHx7P/hInVKlktFJ1SuQd+c7IFU
NpD3o54nLV7DXU7jp0bU+M0annwuqg/qilebpoXM0y/j5PNR69UKa/DZIuWE5hM1D37Wn8/1ZTS6
wk79AbagcuNiKaAnKjqMOI+w3+z0GMfP3+Q9fvnN6g5JpWLlC4OTuU8owniw0rth/sEp9cdqLDkL
m1r9Y3E8DgCkHkx7Iqu10O3cQuuY+KzGza+47i2Yb72mFwRNHoxqwKCUSYrmM/ufLSOn6OCdz7Gv
iJsW00jSXO5pTbUESk2tI9igR8wBM7wJK/Vtj9ZlyTpNBOByXdD1rAsGrcAHJCCKbwKH52XMsxbw
rpbyCYQ96nSR5OT8TUzCPNZ/7yquz7JBVdjysGcSRPiNxvuf+jOyiaQskM7hKnIh7IkcR5oygrkv
/5+5ZI5maz10MGqIScetqrLSrsyDXbL7UDiR38ipDVdn8Q0KcfCgjVI4ifYHyctxzMDVhJjwGrrJ
jINpfxAJBXoVuxivNfx3L12clNmPkiuXU0IyK/NG6N8SesvZ89tbY4Q8MAAod6c0yQU31JV7VmAm
IfqRo7k6qMtIG/gsgbHBFgfVnLYRUTy1dHGAb46UC9FzjAgK9HwM5ERnrLi7k5tzUNe0YawU0iGw
nlJ1mH1MxcnP85EwVFCkXo5Bp4WtV8i8F6EDnH9keCjwpHpmpHe+0OoYKwK9t8HMxYR8FPujYDuA
ycCmuUNtBqCIJGwyezlS/xEVqAs/KA4JxLrG6JNRE670gTHP1ym953eVTQmGYPmt0TCX0gqC5sTZ
RgzWsy3tdVBIYHD5GPHS3f5pN+KVoIkhuRjeVIXsGX6ifg+LJXAaVnb+H3jaVLjTgKi+q4VylKCz
jguP1I8VI1Ax0YixwNlc3/Ku7UOerWlmsXIYXhgA/XaxuzkgIgdetUhhZnj/ZKLp0NuCpgCw/26v
2xZY6HGfFTb5E7THrmTyeRZM/symU5Z8WfrmphIZMQ5ixzRYtYMR/0zwku3MumH6Dl+yl2ErqA0O
pRc4bqd5Zch+JN4dVhkerwKrYZp1663Na5VA2KEcAFgo8zCUxA9HseWjv0NuIIPkixl4wnYWPrfh
vltAhxJmfpNpgE+1XMDZUZKD/4Oyssl0QcT1Q9rTsVGa6RMjlukEsYJTvy5IEQMxbWotBlWV0cZc
RDxiUOwb98hOy63DM4vGXqfxT7aGtmQCeOf4Q2SFUak90+w2OKcwwTV0Jdd/o8FSeqL3afUtTXw8
Cj32GriQp5HvhNGkZbPRNRsya8ZMHuMH8G+yXi2OQW0ThxGkRL/bkgB4JPaBcCyje6kQXH041Yv3
krNiuO69BBGl5CDgeZaffE224I0fhxJQBLz+a8lCrJdFmdHg0MqbiZlAlXavuuQ9vwCa57CtoSLw
gJ9vsm3x1crrqyvd0Q7E/qN8S+jXjtTqw2kKv9/X1lc2NQOVdZY/SEidk9IDVgAF1ygU3246/b86
UWz2faSmgMetaFj8k4G7rEXij1Aabi3ErV5TMghZiUezHr7i9mmsLpJoj9/b+wjE4OjxLykS1tKt
0m2zu11gGKncNLt/etbrGdJCib97iQPhZe7koUkb2UVkchj8WnB6AJxid5Ss0vgytHm72JHDa50w
7MpZTfZ//IHadlx4MoJPVfCk631sIYeF3PBE7XY6vESnnaDw3T45+als73MBtoMa4woDileRwiOK
5qceXuDfe3hwRqxKWiFFYDOmTJ9sNDLiqNcaYeJwszM4/PS6QApsoDee5HlwfTAyUtFUqFpoHufX
xwDsRxlwubBynZTOxugZFeV276tB85JykrUzW5uvXAmhV7FYW56pmtgA3O12iHAX25T4d9Is4Y6c
QMpnA29vxK7l3OTF6Qu6pO/4tRQ4+juRqe9Kfg7yhwuFGfSccYv1txnO2oX66p3nH3n6qB/Wt+wM
c6yi3T8AyT46Vs2cn+y/4w404wfQRuf5hxM1s38NHOz6BpcSC0QdTQvIcXrTzVMxSPn1v0s4wCpm
Um4ZtKI0uojlZ5OpdPkgWbRiKBw24pwwl6AuJJpXKJ+YajhRg1F1N9YpobC+R4TwQDTGmuWGXBzZ
1z1lP7vKBJMSwNoUbzPuSEcz0U10SWTgbCPilMlgVsKNgXLc33j/IF8TihZeydwM80XmY6E3EYZu
bbGxiujuSkMowN8gda8AMUoS0fro+n92C+ComWz10gULzqj0XiJDp2eh0boVz9YTIHIkn4s8e0wV
df9L/cKITOqHI5ctfiopnNDeKCD6rAXmnWKksNDyYSjvR6PuSgaMYbvxhyT93wCu78mTObt8jWEe
ujZbCTLYnSxtN6GenWa/7snZ13yAlS1XJ7fHJQyeo+ztc08KXzqQsXtiApT4J4B0PIvO9vEbSsmu
F/CtkNoTgVCAqTGHW0FKAc+uMdaT+cLqeYuK8i0YdMSXy2EwHH77OFKMjYxfImEU83UBCacwITNR
1/Dl3WLr9wsRNvYx1XpyG6Hp4TnGNTKKoAnrwWux/jIvvM/0KUQMgJ7kEvnW40vMhjUy0iSQQCPZ
OtLcVvCSPo/aVZrV7xY/Dxp9byZ9CmgAFyWUi0s3PZWuia9mv6CWOQnJ3T89QlWZgv08I7LW1vic
LF+Qr+LY1j5K9crGgcIBolPw3Sl/LgZU6R+5tj4Dki0wVsnn9dmEE/xByomEvIjppKLDTuMNxzqE
4ChTBln53yWCGr1gepW11l72brhwUyNrNAtVpYS+epJ1A8a46ZevC5d/jTr73Jt/qO/UomuFCJ4e
m7fEPw0mz52eZQHZrLs3fc3n3+2mIzu6/Du+1E7YjfI4c2pK564Wbuq+CuAHBGvJ6OqQEHeG1hQb
I0P9IFD4txT5rZ//kbLzhAZba6bCogHO7ahaQvgoyytB0FLigdM8C4Mv8xCu6HqK2/3etPtsw969
S556187koGpaqbwy87segEBYJg2bHD/YottCp70uiqA8/awqZP5i4eDG2bT7f6oz4DfhlqW3+KZS
AtKDAKG+FucKfoKv3x77Zdzz9KvbJpYlYAP/vtgVoZ6Fz7SKMG8U7J1RxWeiRPT3cfKFvZMuUYFT
tvBKH3jBNJwwe0DVvHuukL+vv8G0n5pSBJOKpk2dvmNnvHOPNyWaq6saTV2zC9d+8+TLvc+zjZCC
RcdSUTH2O+EZWsQ1hUh+XFTPuHO7g9xdnYPx7S67ONUHO1DFQ/BTi/N+0mQzy7g2HR0S1sXeDMj1
v2WHbQ8C2YBOd2fFU2QcVcX0Atl2b32qCR4NAnHdQry5md5+fk7DwoMYxf+AWaVIhjwjirKfTRr4
THEZ+em4feYyseqT+pAoISxMLEU7ZQVeXfk5SlxAXZlxJNXN3MsuGFmTfgNJuvP4/tnZT3/Gy08a
42Zi32uR0MGP6AaB56EbQ+YregIj/a2BKHvgFyrah5D2eHbpR0/V+UMVhaoqxOQb25TYZp2lnpGN
4MaTTr9bZCYBYGfRuV6FJXxpVG/iuVf55ZgZMztgeDDDZoL1UL6djj9P8WcQcf3NzpzF3eVdxL3V
Q6yA+Kitkgfbt3nBdH9QxlJNMEbx4CZDuNOZqgJHUJv4Gbj9hO9Q0JMY2INtHNTE1syRPdQbqCl7
dX7jV77dmEHT3lqK0BGVU5SjRqKtE7u45nVh3cGVFFdPKHgLkF/xV0XdFrKVqu5oqMSG3WZ1sOu+
6sFRUa3UPze/iZQP4dy9TKyAsN6lpMVoRa491x5cpETaBs2TbMdB7qoQYInIWLKeppDmlUmEoKYw
3Ed+DGDrH/prLhUAcopPZDDy4vx39vvVnqsVtEigbkrj1xIC3JFNHYpNhovm4y331xLVYtYt6+Jr
qu7r7OZJIUmZ+lHzSnv3LesFo910rTM1iBTp3Uu6rMYbsc0wFyHm1Z6c5skdqvMGINitRDYAZgRZ
4VVWfvPJaZQekiwPDYgK85vReJ2LMW1NgXT9TN61ercOkdqcTLqVCkmtY37HQnKIKDbxIC5qQKkv
vnaNc3NAM6pGluO5mXJnjRLRsD77Ky/F+KCn7YT9J9Hap3KvaJ/6X9jBxZNY3y3xtnHDDXXYw5Zc
yd6a+vYnTcCbynPDQCNwAjEa3fr084S3QgjE01yLbNPuCcURsb8apYM+kl8/vkt0eAq2pOVLhLPM
pPakmNwthBBrmqdCCNc11F8q7Na7KPqI6aaU3mX12V4oEh+melY7otgnuwbCnnR4O+ln9VnKWIp7
QyxE3nTZGt4LiYdijUZhuG58tBLcii4M+QDQ2BdIDlgLWOCGNDnB1Rk+TcRt+cKrDPbF1KHr3oy4
l4obPuRnry15C6qtBhNxzWzSAQQTQiKHTNPE1l4Yqu9FfrNnthVpClzKoHmqZ/7mJqjVEvxp81oN
O9+EyH0uOcotGRCYVoJfbjs5n1ce93QRJBfgr+BTRmNAkAOhmM53MiIJ9sUUntMqFLDXk71dEztN
dM5jNEO1U54G102So2BMSuNRpCdeMUrU6hayj0oasJ/JHr1zsyMBbCzFf85QhfS1u8W6/dr5hnRP
DQ8tkZvJfR4tbKb6Dxy8e6NOwgah3FFACqCIK0VKxwtVc0Z125O6Ha4VZjeB4V7hMdiRh10hgmZ0
faA08SAlOpKY9u12LTZ0J2fiYfrSUJGR5OxFVxH4kI8vqBmStI2v2mbiDrMoO607bbE06MrH18k/
s+wFSEMbJ3jv1Bjk6oAoNOyTdh1aBidxIDm6G47/tquhw7/xYvUUF/l6dVYn57cBrymwmR8SHOxB
hNrWemR+RxT7640ymhdNWNy/aX/zwW37EWzicSebjDlh3ChLzf+eA+jURo3drw0ntr1Di0OK72WE
083Gyto7T+QBP0Kfz99EIvJkmzOxUZv00k58DwOxNGAJ+ruB79Ru0vaI6DZ+wsfphSkzZFkbsqgX
Aa5NXlxBgAGgeo3/nCvKWTU+G9QPgU0orbtWIMbTRFeKMzVKsCHKEIrEDEG6eyYjBIZ8Tz3oxWGn
5ZT+JbhsBly10hPzrgTZfhh0Ll7OzBq73EVzM3UWsMMqokkOVQj/sfs+lQFcAhTGapxQTcEJNoSe
564yX3Bd7oW9Dlr15ijeVFq8sWO+Zcd/sZP1kAJJQPj5uEFNRYslDZIU9rOeFUoNoe+etKoXDn5R
UN91gr5jAt612wy/thkfGtZ3Rb9COij5P3iNaWZr+hkC29K81QTiRywjyCq/UPKRG8kKWHH+CmHq
kdKSWprslW7zqlgvW8+j1zrIX2r+yUKXF2AZWpSm2ynh37GIgUl/Vj23OH3uTDuPv6j3QSpN3uVb
tTym2vEMohHdEmAD5dwJgnIGTNyfF0NLgiNvvZBH7lGKxyXW+Ezrf9PpjYacBUsvvn/rH0iGRzmA
qWv04Nor+LbxMt2Vc+y751t4Lmlzciry/1I4Fwbe0rptlqDpQF9PMoLdIMtIKAP3NiRRDwIB5kHw
nMLPUcczGwTVjBmEwUWlxMkBLrYeqO1Fuz3x3QZdxF4fha5GJp6FfY3akl5hskHJwrR0sM6Humjz
3hjXBdlxMj8yys9xNfT0srOao5UJU4STTxb/XRROtLlraz484gWdQ4nsikeKIT62tt3yugiQeLZq
6gNMZ4pmYDj17VWJKSBm2w2hf+qrctcK72diIxZA/mfGgor4x04IqiP53zytQdKNyjMGWsDvFF92
D1VgHQkeUzzIJwkQl9CbgLevVL7etB9jvNhB0oBH0q22NPjfwjUFrSg9uRHvpJHXYTWl1I63PAIz
7oEf/GegRNT/nySHYCGj4oylMOVkZa6t2MRb3VveaQ+CTr6V4ITzQVV+VBWg1zB3uOmTZjZiGbsD
rk1xdLdUM3cq6XYaQZhhVnt0z6c0u6OflaLACmgEh857yglNDl/3yNklvJlgxl9QRZJrq0iYFj1z
CIuZdVQOeY58U5EoaoG2t3qg9RQKYS48qHLa/4lON7gF0UmeFQkMXyKIIe0ACzjS+xJxCjaRSfUL
CCPqaVcUdyS6vR0ZN4Vtr1z907kp6XmXPRs5MWD17dc7KKl+oV4DsdzEvvkCYOEZIBz/W080YexJ
ZCR04LPbMfue+08YRXxap6o3ozXIDByfsJpvL+blrjJXec8rg51ENW1RCgowWcSJI74p3mixy9FJ
RC3cNkGgb8ge8K8PRc2/2miLH362pxDfZ9lscqJ+ChyYcrtBNMa64DSXFwHeMYuBvVlBp+oLuzqv
7KTxk86fHjkDCZW9UQ3XLsH8MNdSlKjZJMo5Qpnk6fL0b3MTUpVqjn7vI1GTJE0105+8ZvEg+N8h
vsR0rJQAkT1Eu22YyBw5tuDYy4ibzHAbV4Ppa0XpGNHRXonszRc1e/rDzyqL4WmRgaybm5BFAZSs
kCv5yfcyvli6r0dQDSyYTN0Ok+GPTu4cEJwRTTRNqT+0/Gkk7paqIb/vvcZvoAXAzors+DJs0kry
8NnZRR/Vli0VPP1R8VNRD8URYfhR5fLWWk8a8VZ49nA+y9imYCmClADe5C/6X3ozoilKErwBgvWt
WL/Ga+hErP8KetGA5Bbqj+CkGFJ13lsM9BZ0KUBea7smBbrU0X0BbIegyiVA3KYwUB3U0kksUzvr
hw5aEhT7UHEwDxmjPLYMZdBHn/z/2fAcgx6fsg//LR2WMof4Dy7L5QUAn4/zPEm0EQNduN3HjNfN
2Rh3Ze5jDsmND2UYFa3lsEYtzHTbzYV9+MWolixoRNeckBckqjU5X4By20JoL91GD43bNmSap5s1
Ilix/+afgi4heDOESkKO1dSAucghm1JJ2hS9Yfu8PgEsa0xqx2dh0sxqKeTF3bOzM8jz5kLsrpyB
DleT5oJtg1Z5faH7jrc8iluXcvn3u8RSivsJJDmlyiktPJJkZ/4g3NFZ4hNDjfKfcrFelDzCjCHq
qTVfNvXJif3UnWrhz68KdsYzf+lCVbWWjvIORmUzhuPaI7rE1kNkcUH9Ue9joMzePiYgL75yaq0Z
QtSMiO+Z62z1d17vcI7OPFdoIK0QNCVZ6wGmypdKGxbSJbZvkwYKK9zVQBI0Iv6bl/Gi+gbxaQ2z
E1wisy8t2bQc45wTY0sacDTi7y/opsiDrvIbEtbdEdGioQh5PtWPc2+gguaqj0/bLdBu9Y/hK5mZ
kXnx3xaLHTcrRIIHrsnga/4EkinOcZcq0ZKuGUDuDeW2UTxZzEuinTdutO1cCzb2SaNIQfazngHK
6jVbIlE6NLTFeYXP5mp8xGQ5oq54n0v9socwVzYgcdySummwIlvNbnJ4Wezp2QRNO2KGwtqFPLTg
TAEo2Lv/0811bIYvz3jpIwb89ZPpGnLy4nb8YpER1kY2WKrHyVlG6c1/i2ZYwh3TY+42KDerm8PL
ONp02RzStPwE4WiBwGRICqIqtjNRExR+cV8odlPjwi+89XRd2QkDlrNY50KjVOXq2i+EDr1uUv7K
e6o7jOT+nskF3cH7kxOxJrII9ibosqBFMD0EVgzC1u+aPoxJhyGIPUazdV84C8z1EZIGPDhn9oPX
aSKgaoPYBjLiPSBrRvS3+lr4hejAa7h0OYWh/PEZXYMtjLhS8CbO/rQV0jQhRU7seLZ/rY15V3rP
UtC/lEnyEyX67x+OYs+cQl+ljlUgc0W4Ckeh6OY4oJ9RD6tpJTe+cfY/b5c9Qy2KvJSAre32b+3c
KLe57TVp0qPpZgndd312dZvqH5rkSGLYBZKuRh8KmFJ1ShOnZggrsnSIUa6NpDCo6nPVRSQKmB/9
G+zscZIKKKBBxlkXqHRd/nAGvl4WtO+rj/Zav7N5q5fcspAeyChB35+KdVKKI7kXhmpdtXkmluRP
j07hKQgsfrkQKlj1TulFTmv2vVJxctevqTUvike5WmsluweP9qO4pIv0FvZ6MbhyeI9aXY+hUJ+1
du2kmjPJ7WZoR1JaoDVKnguWDhpxWPSjCb0lygbnUY3u7wWn1L+90XskfJs9BbTXCHzifnfIxFXo
8YyVDVXBUBVGGZI+n7axyigepRKCuuGsykyzQTRH+nYefty/Z82icpilbPIRxHiojKLkttFDsDUJ
KPEM06rQY+gF/vAwfV+stif5WNHhOCn6hwM3VDDQ6hStapxhNGT6733eHMOplCHbK20+JTi+80ct
Tw3FQeD5KdueMS257fQUoQ4gkP1LoJ07Sh5RS5WZ2k15HIjI8mBToglBLqA3m9+70fymq1sHy7z+
UkbfMu2PsP+Am40F31cDuOo5hO2F/QQyVaS9Nt5hv7hNYzW+pKIHAFAYluyEJ5bAULXhmNrv6J6D
eA9zzkx5vTr5ergPsbCBqi+2IXgTrBtdy2GlhDlDfO6LQK6VrSlJw1Y76OBQoCzM/BqVMJrwt8I0
WWSNzLTiVa/O4YOFmIk1TmYj7yEyC5gSumFcu/Xj1WsIjtjgpcNVrES0BFdVpClTBKbzthHcDidU
6jDkVh84gtKBRN8EniBHysMGu7vBywZygW2wD+9tGxQGKaou7CyW44iZPUrY2X+l3TruGn3F2fir
8hTd0vL7wEsa1dtK4Kf/rSkAfDLfVgcn1NBhUl2b93YRJfvkCbPheFVHyRu2gF3BiQ/pc1S+feGr
fTncd9JzePxqprsf+vZLCzy4NwYXjeTuZlK3ai1JPPSqL3o54Edn7n/zcjKJit5fQE/ZYrNFWU3l
gpcAn1QQWPI+tNWJZBw6dG1P3w+4jc28/oTox0EYc6S+OdKCKvuplD8NSbmP3yqCrdoaV2pL0+bG
L1Hqe/Po/x5BI0VB0bvcWh1wJu8c50IIYfAC8HxhW5hNdfXPuClP9voo7KUKibFLtORVrXX8qzVI
Y7uGRhzim1xnPjSSzCvioYjMIepIW4Dd71YNq9rvy7SBOwTJQZId0qZoqFo/nnFS/4awMJkIOG2a
dZg/pGYwmpXOykA8yOBzJM0boYyimmQGODe7TRq4rTuDPOqeoNyp8UVjOmtoTKCb8z/m6J+ovmw/
Uv7g0DU+lr4oGHoJgL7NRuAI+jlbyIMlg2hBDjGA0iUKEoIY0CEMUHRLaxtyGxJswPfFnycMfu6r
4abYXsXPkTdOc5pLQo2sagNh6r91JuBvq0pLhkJ5aI/PNi3u3mi3LatN8HkQa11SdPH8BlHSXeiV
w/lTxSjMy214ccCMY1MkLh5kXPqFUjw5OI1l/YvfLa4q3lyFhrVof2KVDfeUngBNdMBumaMaZXOy
nX6TVagI8nokDuQqck5nBEkvUwqoJSwuyp684yG9DwLoX6G/R2wtn0lhe0055wb0TASVwSXuSOcp
6537Rid6jEG/enVgQ/sBXQU2WVCX/emH6W/d7T7rQ+/Wyre5Lst9r5yVdvCuILfurgtmlMEJao+B
5wK/gT2RhuG3hW6oVtTl/2yG+rYtWeZqISv4A8lUA+txym9Bcpd31iwPAzJLzK8tjo/ErtcgabmJ
u5q1KDtlmTJqZWPElxPoOI0aVivpu560N8ywksLo4CFv3Dod4cjT3ldCjkMwdUSU16j5Z5JaAROL
EMlAUkG5A/qIGHnJHLy3mFzFwARCIX43rSVsDO6rWy7izaBrYbCEz15FG04LLz8paNHtAWlLyDs7
fx51rj2XQQtBw/kTAe+v+35TKQwIUjs6Y+XLM/EcC/6Q5+Mv/0FDM3vO2RE3n9DKBHmNaZNIpRNa
WrZDlwGDc2qownb/j13MHkTYb1wUx7LXIel6Jf1SIgiLO0nFc1ZeohJWUYEi8QinYjQeAatcr/H7
OfzKf00zYbaVzJ3AkFYowwBC6VA4SBwcJ44HduYT5wIRQbVCBAVnNB4YlqPcOuPkPn2lCoq9IOlB
WLOY51nXeM4LdvPwoCo3Xger7lMX9Ne7gXzJEFqYZG2wtdHoFB+6xMUeYTtFrDIDF6H3BYpdSNf/
mAxZMJKo45Kz4a4I6qh9MCAaRZHwqwFfC+qO1ujbwljItPJ+Mp672KI+/7vj6DUZZ1V9QB7Igxgc
EWDDXLsF5v9QDhuyZY1HAWa9/xfuKK5Q6HqHSips4r3Wi4tk4MhtvDCpszzFQka/ZrJ7khZdciEP
ZPN1MksV0mLCqX5E5DaoC7auebrEZPQI4Gvcty52KC/zDdSV2+4rUc6zygW/Cw+fXFr3oCfo25/2
MEKXMgqV68+oe2R2//tYIrojSXlfVog6ry5OVJTEncmFcZCqzd4IBOWXf9Pb/K2bO6ZpSL5YYql4
Z7WheN3kXeX3vsOj6F5mGK8Mk1KPUXsNzM7BkaVLxtcyQhTPIjR3J2iwF+SnCpeDunicSXIRHdMw
3jAY0N19EU74LV8fZvcel6FrcdaPXdjk/BKDoIifEroS8q63gpLnhgApa1BpFLey8whNKbTzkBGK
+pqcsTzyRyzWmhgQ2SR7PgtpjXKVTV9EO31nU7P9UPFGB5ky6qHffBpwlbk/fp5V93chvcapUDzz
eUPd/6Ux03NTt45y+UQJmWhxk0rok+NvxgUNoEuRSJpJS4rYjF83RyHGJ3m6PgXl/BpCEDlbTjpk
51gE+3Z3AcDTDdBAvcb149W5YJ31LhGOIXhD47nPvHPFAHt4bfOQ55GHqYyAdmvWW6YNPefePwp+
7555Q8GQDSq41QMMQBRGc0WlGYYA6eSu8L4HLLvLlgfuJHAraxSPQ6ffyGCcCQSfrIsGALvqfmI+
S0R5jWEr6klsktTw+rp7cHytf7vMVNXXeJQthl620j87TtOFMcFqiqBbySDvCLHTA0PVlZTLOg5M
tD4yrhsxCrsykFq7mPdBW4AMvCgR9Z4cglTIQAWN0dc71pTc0c1Tt6kAN001jpMQmL58hU6dk2cW
mJ8kHlB/2OO/Skr5Qob5CjZkCdgNH6HfNrGkBWuo25RndXXbd7fRWoJjWX7W+yVeyXYMiiiRtGmc
ldwjmcoLzWGBqarhVtXCNU9+lQ4mY8r3ttT5lDPdqlH6gjdSjA7/6tWi+MjUEEpJ9sieltFiOoWQ
eUUcVSGG43qstGqwnmuZkm/AQJAnzvIBpUyIHR9TbfCqIVwCiIXsbyQFM7b27xc4hVp2v1zrdSfb
XY52KQfncYsZntoajCPiSsPqlsDFZW+QqejMyHodMXNBsM+0gSQ53R8AHxcq2yK462sX6yE/VDb5
eXJqEQJwKTPqtGdJ0HZye3abuOsU/vcnMgB8bfO0g+7eIg+dQJrI/xnE+LPBw31ylfTWQeXxlLeE
8MCC/tqsqUJU8FwqokgW88i0H/+2S5bygUDRkpUh2qSJ71e8pejfmu+s8V+VJ0KyK+60DhQeRDih
IFW7+U/8FeEI9uUdbaAccibvXecDI9HJ7f/d5sh2zuaw+uxqrABMhgFf5ixDb6rSKiciGjSJ2FD+
SfwqL0IEnTN+yy/fRBJJHE07DzOtoNWwuYk4xrpmoarz0iq9utLXCWJDazJjlYGB6I6StPD/3yr6
9cAkTtKezMRMssC0s7CsrwuLjOUUpIJmjTZjzu9pKpPDetkzyHOMu/qbQj6bmHUTOrlnV7Ftk7OG
LDHm1Z+dgz/d1G/DvWfyup7nlifg7pWbuCr1JnPB7OGIWZAU9jvQYOpyxivkvJuAOn22KoxtN2SZ
KUlp1C+nNKISlADjGeF87TX3RSmKfzmFG+cUfaKgY4gbLB9Ts6VwMd584VzhtOaJemPRQJOwBG5a
WvuwmCPaN6XpadfAuAn0wX+kII7pTHllzHuklBXu+dMA4APSjGJ3NPuiIDheLcTSaD0RbkyOuc86
EQJkYBy8u/KFYOSA+2+qVjnZv1dHvABTWCV2zATDQhudtTQ5F+BKychWOWNqkrbTgB+nSGmVPzF0
krjR+QejuIx3E2nfPy1PKInlqdE4gHJBf/SDcw4tH0szqnX80w3+tLMK+UveFMijGLDdFSeqzJ3K
2U6CTkpaiYf6zCE3TaLOHI+4AZvdL02EUBoIXuEftuo+mfFpnsvd0xVjGqAO010NQf6/33lLnsoH
+dpAbqIon4zMmEIvKJrFH0y7SyhEnauK0lEZne7rOVd/YBWt+3STrtgovoM5Bvt3bUWKFb6HZwiD
8qz5d6ndtJSGPjIimN9bgcX1MBA0rWITT2vTrGfcphQhffQVYAckaOxtGuBUW6nelRQpjFmSfpkO
gDgd+dSFdXAAOB7U9EF54lZSvclTRrA35zMDBATyWdJCvudXDEYkiRzKW4gd1SR2JuAfErnnRoX2
yhYPf1ul27n0cKo7OISU1zGM1pgcYYazx1gOWyiorHseyN1hMp9OvyfNTVlyVR10QDJ3WnJAZ6XN
ZUo5FdciavFo2Ukf+jDQffivxjWqtzH/CwA0hBcAmzYuu31064J3PpHc2rX8qcEDvyyFb9JWoPwZ
F4yixRjpZ1uKKI0ijPJMSKkivB41VevMhyxkIFr2N8yPf5PSnAHzH1+sYT0NJ7Z51JL04MxiRga0
u0VcisbVyE2/3f/eNQPUi8MYONOC6quTP0hO6spF0CeytbzNADXxJmXCClHAsB7EBVX+I7sVbQzR
TeanQQRlwLgw+JOaxmv8xdBJ9NBtTyBlucW9IVjWKV8tU5o3z2ibOSwt3/1w7HHK9yZzETZ2RLih
GIxIspmEU7Z9E2MwWoekKdpCtt1MsHPzaotCrREb3WMElwDE4Zg+ok8hX70wWg8HHG+Vu3oLYO8X
KsX678zK9wL41goV21cBPj6a7/ktmUmg4mBBEYU1p3ZknjFeAbkvW4HAsujUmcxyu1021+7gZvoA
qqcke7QA5W/ev/quxr7FvZaD3//ST50lilpwlfnp3u9pPS4foFUC3hnnmKKrHtdPE6gyIpLQBKSP
LpueE1+zCJl0kmLoe1tGKyJUQh3mNYJuMotPzlEic/4oBBtQscuRnhLODqJejWlilhOAaLMKOfTv
vxB3dCFmML4xu9mvePk9Y6vuC6WsBfJKz5DiOFEbQpWmtZSJo+EPE9nxTPmGE16S0R6AonICthe2
1GAtjQuRnHsGzBDeYJfFSBOFO+52w3NoEr3ytPb8+ghlj9IOUMrNoVJqR3+8BFKNT97MIcQAp5hm
eNIkhkbidQjXc9laMvwDvBCMcHGHfylUE6UrrUCg7opEgEKwhRxaovF4hetZAH3upU7QigXS9uML
OlP5ItMD/wQxSAhLpQBW0RA7iiAGi8aU1qIth4IgEaX/moIqswwccIMShAGV6O2ytbNgMJiW6Jp4
KDJhfVFhlYqgcX+2QNpq/w+KWrXgraiqgCBv9G2itiDFPIsW84oj2kXt2y7oGDym2feBFuvA20Fu
GmOsap4BqfABdPjLNnN0jiU8QzAu+UCn2l3NR27iXqD04vvNHhSNmSgTv2nSjesjgtvmuF8rxLQ+
F3GEdWE+2V2Upt8BhFdwnw5Q/cFAiMkcBXUvjq9DJVeqXnn8edPMURRhVvlkfqrERE1MkGMLAM0y
rDn0ChkK/d42pxB7j5XVCo0Ls80isKDItTFd/tsOPG5pM+FMtWjXhWAXzD7hlRgGX0inS5rLt995
s6jCdpHmPCY4TvWn5ITQVO/Abz6TKYyc20AGtPSCgGKpOK7HyEPV9t2CjMun4azsQZhDaZ+1nuTR
XgrEDyr92Tliknc9iIMIaQoyoRZxWxntHvWpzFhOZZgFGKKW4C1VVx8YuMTUbBHZZOp5Ke5UnAaE
eY2bb5OZmtugt0eYDjAdlkVcFW5h7TAYUfPCC4/jcQW0U+X2PlHb6qZEZQD+FTyZPstrpCwvRAHc
f6vZgnOEbedigV0L6IjVQeJItUlciMiqhK92Z+5R1vE9zIzF1QRmc908Ij6OgtP1Tiy7Uy87DisB
ao9/hFYcarSUFfWDteYbHiR9vD9WLWp1ksjw53i/5AHCypw/fFvIMAUEdu9McjDfm/uDKXQGGmiK
X+XLxcbZS2pC5IVdIV3qRfTYEWE6iqIRBSmIQiOI4kxHzXkNOOPgME5fFUsMmA1bndR2Y5f0ndlQ
dqy1b/UuG8F9QcQdgyvFpGvacXf/fQx4phw3Nm3BeBCPqr/IMgAEbSLHeyOJJ9zZpmgYbHmOILRu
NFg3Khb7gNKSa+YJgt6oTuuM/GlZlxZ8gnwrtxcEWfl9S6nEH7gAZLlgSj4VhXjNVbFbZqXs8wVP
N+2kjIj8Fhq3Ldb5s+5mXpEWH2yRp7eiuyYHNZoHc9YxgW32j4czGd917R25WZrm6n398fu9rbs/
pkBe3VsxrNjq2BrFd9S1lk/eNgHFbVOB5qPzxFuDiyVh4gnbyVLZeGQis5/VukDTNHp8P2uNlcGm
cgXSKrwE1RyNX5J2BsDzH47rBrpeP+QIo4YbSVcsjwlyjHqIz9MMQfACIE/P9RApRV+8IftUBEwj
i3XthdvcamorK425l5IDXsM5chuVqXVvjCMa543EIU3MDFK66Vruvb3ZUwowDyMw9EnM832dr4Go
kOUYoq/dD6Pfkg+UnvblhHUyDI9pkOZAw4o5Ez7vkYG6RxOQL4dA5DpxdTc8T8gfSB7AGYsUYWLw
fwOl6UDOI9pY+zC5vDI4HSLnR6+WY1o1+9Anz7Z4XKWD2V889GlhYFESKlquBxS9evTulmILadRs
cIQAwtp4Fq/sqNx3+uL4Q+tvkDVmaVZxOOxh3QpO4MZxSi3q8jxDjQId67Gz8USOmRS3oTXaKuWB
TiPepJUTnS7QRfu0V+dV09ni/P3dKCGCnxGMyRG1m/4+R4lhyFqcmtJwUoR5CVQNpP2Ay5HzYrAw
xLW8Ym1gcEWqAnpf9fkt4B59pvHKjtlTFAjSAcZD2ZbuIdARg0d4SvNjUMdXI+rzPWpKAIUHkV4C
DirvFx/jsSxYnKDipx1/N8pT2X2I3Dl5w2IxELNLCrnEMu4tOPpRu4tgA74hXmzerBJWgibF5daT
ERXRe9KT1dNrO+fjRnSjPoFgdt7g0V00RFGVm2uWnT49skl/7SRUNFJIlfT2VowUFtiLKUFj1RXd
kmeecV3exynS2Q/G9JfEubdOla9phUJKqDw75FtNirWlmz2+7mnl/ls+8xTMUx7467Xo8hFMZjD0
bfnMVD4iCqt8iY1Euk1AJPxn8BA00UBQ9utdTc9ZDGALDjXvwmViqoHRLuasN7vAmqNq56Y7qkJB
EXbL5QJAjcxKR6ZIGdl74o7rq8WPT2Bi82MSLOjcC7b6YQolLtK/uOFSiSERZFSQvSSh5+mrD+Qz
pHAcyNCkgweIz78nwLpvyyK+bCFrNkD1t+i9UCkMeEf+lstPw9aHacJJK9gom+RK7mUxW3WU7qpU
9t6m9hWEm5hc75NVnyZJ5nBQ0+bHpSiKCvIqFiVP3GDCfNIiRV6PjhEuZSNejZqTcUjwied7rc02
BbV3wY302MJ2etcY/4/odlXn3S6hgRJrd0tc6auvqUTFd94ncjAoVMQLo9Ro7H147KaSRihhMcmq
YMCzRPkeii6uNn3wBhKdsrRb2ol+tkY4wL5ucnCFpqEp22fs3asPZrdFbT4beRZyFfIqP4I/EYUY
FakAQlpHeYWr+G6IOguaM9hj/zGAVmxWEgsBHqDfgQW8mEadEYXB/qmvgyvV+cuTGTG2kD/oEUYp
/aCye8aJi76gYRdxPUbNg2l0B2CPxIJ8VW92kKxigyZ7KOSgKYyGX+AXzo2YdOwgV2XLprU/JVIu
ijVFCaN5cm+UBHAg1XhDcqVmoorBZbKkgibXGklZJ5ODopv/EaT4d5tnicnPgRD9Vs2jtp2SxtTk
D9xTXKfAK3iigWyMaPQDQfDqyUPOQo5Szyo6EACDd01PUzT+1IQkcz8YJ34BPzrgGy9pt7DXwTGM
SzPkq3hIK6uHNO9TClcT1+ikgtIWSCCcUmfAa5edAzZqxZdQMhBqgSeIckiEW8Eft9hvyEykadDf
NexaxyblNOXYL3Fb13J7fUXB/JU+zi2PxFOBPi255/+8AchP/rh4Orm4T1AFiOtUaMT1crgF2lfj
/LJg4ToFNKZP5wIBJRfBJM4qL8MllumhO9rF0TztwnA3A3i4QhHMCyictEVROuV/iA9bltybVajv
ShqHOR0gdu1DMuQ25gexorQddqfuNm3aVKJugQa1iRa8xHFzmMIpS1PrdEsIW10PKaCKmP7Z/Eos
PqPK08ApeLTNxwp6S40ptdyfQ6ZKmELtGfJhVxsnNCPoNHjPKEGasfGTnvwXJqyvbbSHDLE+algl
n2GLRligN83XvG2Kg/FZVW/QuRsYQrqymRvkLxuImqrTM4SYTaQRDWy7iBAPXYckSICxMBi4canj
uVUak4KJVyaGdw2kjULyeZfhqOI8W7rkLcnaavBMXu1fuF5GKXxZpM1uDuywF5sVNFtvQjGwZRk5
Lh5jzuWZ5byyP3wyDGwl6HBb77rPgQEVsHeyLudCHnDAFcuS/NVXkLu3V1FuvEYdQcw+1Tr7DTT2
x55C9IS781VgMuaTSaPPxq0h5clagpTPQFB2Q8LfhvaHaeIsC0fH/ZpBxO7YpnnLwBvhCErZLnLB
VUcOiZpJY8bCifHk74wMi04sywWJUTI03rGIBjW12WB3br82HTTToYSDBSYdVptJytfTgIiFc61q
IPpn32I8WLkMjiiY6UaiepQO/l1RYb/ocgEj3oNCVUYQFzRZlF+NDlAhr05OoypRzFdQ6idfCW2D
iyFurxk1xUN4l4xm75mqny7trNk+Kga18NUZUGlI8FvjEriT0c3FIEPrJjjg3AFyAfQETVNPRVbA
UsgpJLcQxTcSCdo7j6x7pQHAFj0A6NbCHKYJbbIT0LSdecU+Vth08ez12yXc5OjPsUi3GOu+PVQU
TRifyYdfNajWWlkSE2SFfNYWoEctjEOJDUWtJCqQiAmXBzQ0QGo09JdbqX78ZFE0O492z3LIAyP8
61MRm8fzWK6JFNkOVb9ttIobxnDbnV5Y1siS9cJKfOYLmvU33FRoJnnuitep6ZFas86SDyIqzbya
hdSJOPHu8zqsADC6yZeP9Hy/IK+933SmqJknT5VLsGkUBI1sIkSyIk4r5h90D9UBeqgp2bG0JxiF
pwcOjcULtUB2GXRR/uFNzhA33tJoprhd6AQU+X7DFyKf6bHoFmLJJ8iNddXtfDHa2XXek3YN8802
vGpQsZW8+WG0Vum84gAZX3wlGMs2JPA9OrxcIg6KZvwSJ04f0W4OXDKI/Yf6H76h22xvKHTJaMi0
r8B4Mqsn1+RzEoSRrz4n6W0veLmjYsFjzAzQhZ0gL6mlbCgiTVcv+LuO1IUG/2sY6kDZpG19fJVK
xLIHDwU+A2iQyRJbmpgle8k1cYtPIVKdV+yCsdR3w4wb8hCK+bnxU7IKaUQ2IaAIMXY8AjB7Q4TA
Gy/GXO8jHmClJR1iZGOs1jo1mzXXocgo/gH+rDNNOUexHg4giYHP/bUn59cplhZUWH/htWy3OyfP
BdiZMOz2R2am3nQk7CRXQifZ2P+Ep1Y9iTNnNbfjFPIZRlsLf/pOJY7bceuI0CVUSGsPE/svl6Fo
lrFIeEdyXADh5M2u6zlbLNiymTKTedBlD+q0Bd7g5DsxGH4QwkJv4y4xCDM2Ju79R5Og7a5sWbLc
ZcUe1Yp+CD3zShY61Jd8WFFyeiH48LwCkB7EMOWoczTSilA71pseXTP27NeOrk0C4DPiFQy8XOMU
ifs6rinZ0w1PTdwSojDAVx9Em4Z6Ps0KbWqJwFVKRyGLCju9yuSV6OVj093gV6UwHdJw8OGFFSPD
bxRwEn4zp1st0QdzAtT/flllqFVMH5qVJYAolbmmgnnf/LpgoTYU5+6s3lQNkNoqeEMWKpI76buw
j7uTkDtZlwkCHNrauHrSvfcTWSzUSVxzhIvUTfu0PJ3TuIkDHmfE0ajsdkP7v2qadYd/Q48tAycR
upl6EqLp2e5X9m+M6gKidwBTPsjzRkQbcpSoz3GZXtHwQCcGB6C+SD/4oDErbvQNIp2f9PPwQXaV
Bb39aAlVDAJIw69NQEbe2V+v7pch/JqD1hBQU4jY3hqklfeP6AFbhJ4YcYw8cEK3hIyslFFL3Es4
ibRyRlBqOR0RLUmAHlE7E0atvu2WBwrmNUvQq/EQ3SfpHIk8XZnhfmglzaxX3zQB/XEAbeXPzoRb
KYTjOC998tkPCaTdnSHDqn0j3OaDx0KkGhJUWe4vA+Ekn5PWJFcAHczJuvVTliU2V/AILK9l5HJp
ytBVfSiKx2JL2oHEEk2Cv0zyQmUedj2+UNBTbvHp2ySN9vpGuQ+arg1dbHJQAzpZhwKuUmn6n1tj
l4vs5y/+EZtSCnNEG8IAJGkYIC/BJF61s6dXbFVBtVtFO9u8jDTKkEcL0yRcl0VhuFu2KXcTDDUA
PDxfztaCkNwK6ECU3sDT85a3WhfW3+MgqpYgZlJOKLq96OPiCkd6eRuME99K8XpQH6m/OqjINhoN
yeUfdOP79JsDobzZvqtD0JX8yYpjdKK0m6jMpu6irg9a57yC9aIf4NrBNpLhrNmxL+jD0+N3qsu4
G6+WGv61SyLE6412BQyVEQ4CAoh2iP4f0cdu2rvUobnlGQ8VD6H1Le+HP3CxbZJXJoYhwdzP84/3
LxglemyHLk2b6eD8iq8DbFDPVvlTPdrZohY42ktG91ilTUQHyOE4gr2ASX2O5KXrScqW47jMTuca
9/X0++Yd3pzMFhVg4EqiKD5L9RkNG6TCgkYN3+C7QJyHeyG39QEaZ8Zk2Y8jiJ03pu+yxsu+YRyb
/MzZyTz44PgO+/onGFwKMVW5cxhDGO8d633Rrm83sNgoeQWRBmb8AeIgBTL93B6DFYbUgAuPHGix
DH6eVyqiL4ZKfDGlf6zeLeyauQkAseJvgNGteQUHP5hlIVgbbQLPWcmDcA3VoJsJcqsE9192clod
eB1dnv3bP0KQ8r03IOxnqvV2gbOCXUWe298jy5SEKg29MOj2BIJN2J2oUUsv6ZTbaXEKODGFBoL5
iPnbbNPS8n1rkQhle4tpNbGb/bEFIyXwRa9Vg7xwQO4sK/Vc+tBTJ+ZZoRT+Yiw3qyD5p2u9CN7+
zIPNHr/tjkw0lcpB3ZGagueiI8vB13bWgKgkuB1qxFAo74WddV//uKwZPfbkzWUjAZR7Ml3rtQfD
PbnVJ14IzuL+dDhgXgWFDn7oiqyk8M4mGJcnpNHWNAA/wlbW/ertebMLesASJRbDXNftcWkCLvhR
fLahNv0fbgb7y2mll+oGdQcAKaGwuqhqD+av/TTzdmM/Wl0KXKFEW85EevMWsZ02gG0reEq2svGW
8Ejl1g18S0uae2voI8SB9Pkqw9K52KdpMHJ+bD18db2RKBOBE9D5YbnyQ4ocUGlLtTxdxqsVtSVg
+zJ+N3eiybxkcAwU7l9tyvqcmlkMzvwxtYp7HW7XiVn9stwBuGZxObFAIiRSafzM84yGo/T1Njlm
0g5Z6mJP2DB76az1RAYJu/0MrqpoHHvqLCDcmes18MDrYWtBxNMPWbZ8B6tjb/7mWzZ0gIh5wArS
E5QjIrP7M3/7s+NJQOEJcpeAo5KMBHG0JRklQ+nPiSkl7xZFBvwk2hMbSE360LJElKASSh4CqiaV
WQD79A6Fjt9d9PdsBCrxY9lM26J4SXHNd8Z2+mZKbEl6mnxkl3YU6OSHpWmWY633BO1RyGRcDtzc
GC3ZRy5iRTdLkONepo34a4lv/UXHGdWkeMt39y2HtxkRDWxbOeLXbSpTtnoEi48SgaJJmN8EjAit
SsTVxCrEtLNc4J6xHXSIWRBeWmwEIejpflc0DESey38IuWMvgzQE5jhaB1yrzsy7gN71giErJmBU
D+Szu31DnrbW8kf5e3zRctVqmA3OtwNyE59+qeXPqWLT49dElpvtfhBY9/8MD8dl1zOjZEvsj6kC
3LCe1ZjY+x/axh8ZCzdM4K6RAEmqCFZAHwKGF3eNnFus8eAHyw7q/SZnWCBUv/gxEQn2ssj9b4wC
V9HgHdpWRjxF8Crgvt5llZ51ID8xezp2Iskzan0418o0YIsqcLTTfma+G4f9/AkRiDEjbDk1gwx5
7NJzkkddmvXYjJPKS7TemhiEFuQlLyibAbodbqubIele+37LXl8xvAbVagGRP7pfoDYoJeVcn8oW
AS962ZosKpo0sp9eHNLcdgvXnjyacd23lXkE19rOiStDUXpGL1sE5ZNQMlYRNQJI6jdW8ZMSw61V
7kzo6UlD1/SK7lgMzAJ3OLVmzmmSvmDhl4QW/SNGO+VzeXvuXh59jG1cS71y/hYpqe6thf3r9xr4
JXHM/MDuOkeB+kuTtTLWcZBilGTN2y8mrIknVsWOxI7/OSIKWq/rYcnEi4tvA9H+42lyog2ALu22
9NFQCPt2wuxV0qYwDer1XVRcLCny8p327UCXXhz5vSSuO/Uy5JAt9NiN+qAuUUB02bpgVSiHaBjX
Ut5N9sEcraN5cipJteuw/3K6FFgmAhGFUG/+o+KkeLTKxKUGIIbIcyrgNUWOcl5iIz+MKKjDj1UU
LemYv6fVUN6sl0VlBLbUc+EfKAot0i6QW9cAxcteAAF0JKy+8F0gcjE8Qt7FH+xpSkGDSozCNthl
nOQQuDiU6MI8DYS7xYwEDYK2yOYxtBcp+JckO+QDjlA5cEIuA3a8eJ7xILmVaRjxlNe5BNu+SnFs
/53KXbqC2XaCBp6QyFIbOwzX3CPowo1sHtQglZoey18xb7BJbr5ABtUTXmFmsZ4aK+kxaxiCpvkc
a0sbuHEy+lmJfkxLv56UlNHdA4N+mMU6o0cvU8AtU21SOLrdzI2qIuUcZQqvWKeyu7LvwNw3eV4J
erPKCj6gUpnDfjI5G/DwQW9DTyU2G1whnwmNEgf7Aew7dqGN5Mu0ttB7Xu/FMCfh+hc/y7x+me45
1wMphSLQxKtUw96EhX+82VcSS4+nRcSK+TRejP0RU16Hi3YPZt798pwT8WvMAIZN8fGzLBpGAvsO
rDG/F6tbXkLKT8OFKS/BM7o20McsgsIgJZ4h3JHAddjs/WGX4dsusG4aRr9w60BKCVnUxspW0QzY
h7JubDYSp1Ms81fEdin+kNBZEk1bQdm6/nsbnZSKCVXb+RXCd1p8C1H2V64bUxP9Kf+kFIw/a60i
6mp66a/LAS2Nyr5PPbDztuG6uW7+4lrSdmnkfAoUexLR9tXpx/vmkwBYhvN0z1K9x9t/aREGwkeZ
kjUw7xM0nvBOBrLtfcixy1/9T3NMcnUjXk15xjSslqOWOqEuiUGmipVd5Hpwj5K+Fq2Ad/XnxBY2
Tn2y1H2TD8SFuk2HfS7MZsPB/4y3iLr5eEwC1ByfGAbKdxTBXPEZ9UXYGNQLiUNzLy4tC+PFWP3v
5yuxQ8QIZlSljbYmNJSmCTlRVxxC7EDzZx1y0oCTGWAoDOL7I5sfM5Q53l/xOoIacjc276H6GuEF
F7TkyzjBkDsZ5wnTmFa/cou4FDx9kmiAxdglJAW2tPS2ZzG56VDT4N/T5Iou1rlhnEvkfKyh6H6Z
jmkQff2fTUdsIheRwfG9IpV9hRD1dDXE4Tsaq6lHN1kM5Bw0Uhdcc8b7tMPHvFEyRJ+XOFLNeoUa
aVhnGloUDsQrEFF7rg/i/HgJg1I7OdevEFwpgzUKrncsI2x1nErHb34LmKVPdXA/2xupiGbXKw1A
AdrkmJYe6X+p5oLExsuAmM7dFX33mWFTKay8W1CFsyb7sPc09qSCBl3aoEYUFnA4MRFpRFIc4q4M
IY/GlEnUpl/Xh97EOaZoPnNk5twSIiaeJ3FrDApxTH0xF945vJ2QbC06RemDxALb1qkbgcWaVMK0
IUjkPg1xCrCr4Ai7RogJGhW1e1+GbubsCzTZhN5pWVmhgAMwFYZj9U1SSoKWwoK6Hk/gLLH54lZ5
2TqcD3tm+zONQRCW7l3adnR+w3Yzrh8mIEHhTEbK+yAEsXkr1yzyAxWOtt9EMZRZlIKGfjScLMKG
FaSDIwFuy7WxvfRfA3f65wPzfWp0z53m7xS6g81vEKxznF7bkIBA3n05EsjZz+8A2iTGv8Ys3Udi
IK22bHBBsT4zsTaI4BE4bMj31Qi6MTlk4bn0cAdUKEP+Hkp3xcbOtOFhhWJB1i/97aj8WqeWb7/t
UU+gFK6ApYz3WQxc1J1eaiEUJBl9fgsX04DTLLpsN5RObpMe/98OPQr2X2x5J1U8lnU4upE4KNfS
azP+D3hluMAudy8gasyjOIt37wvyYqUYbQg7EKk9J0IowydwMcX9ADusyyrGr3+12v72T9+4fBW3
sN/wz8lBA7YU3IELYa3BxXtAmnikkEyB2tYE/ZDdgO+qZmYpEOBrMEmXRkhWplIaDWolgc3HiCyL
u4OE3pOlEHbWFAh+JTkBmEbs3oc96xPUilZmc3J/gB49pHnRLZYi9w/VcCQQEzrmX9Cmaj+JuGou
Jv/hEL2Z7TGZdRMlZtKXEcHMHPOrOITi7FovhF7iQ9jJNZg2ALtXMrgp83SE8WWfX6RQhDHwFs/Y
MoppAVp2vRMia9gj1EJJTCRn2f1Yf7ztgpYeQBQH+7+hB05XGfRSRO4VaQ1Fq0elowen8/uaSww/
mANKBnAbUNoaPrkY5wX0LiFnxnEVQGipN2rdHjc1359AWErRSFjZLTSlMQL863sSZMu9SW0VBuOV
uI76mXsmEvkS6mV3ZTp2UTNzTvLEaeNYf4YlDMsP9PnlszIZJHzwmJNC8Oba1D8cE3velKHMRKWp
hS4xagpeML5Le9xt48NGaA2MwSrymeZXIMGPGHuTBs9+SOCsvYbwSmJ57WJ1W0E9Mnt4qLpZ2uU2
QmQUYfYaKUFDQxwwaoq13vvE8mmFVC9tSJ594muRAxO5FSWJPBHKVFrLEYj8nrn3UZ3T0o9nxpBz
6cda5YDVpjITfeek9tMnAfM88tzv7pF57IC34wURSKx0+Pw79GN2e1TQY4KKgFytL4LM8F/twmv3
JKUCZKpqoR5ch3yyCjKTSHBT6zKBb4v6EFICAKrgVQRdIkqdgA2aPZ5a/utH/rarMYlm/b3AlS9U
4477sNS21e8mD5GW1RRtwOcRA4YQcB6k+Y+w9Pb0of9v0NMlQMF8R/eszY7YHWu6z/55DUyV8rys
a93R7RLCfYRA0HVLizpDWSyduNV+ZjSRDV6VBBctNJrZiyaHkroceVElgjrdg1vXfatoNxEJsVS0
kk7Jujhhuzf9vSTEUKaUReaMoof7traRlW4UxDG2AjN4MAEYh7wObGcUMyCNAsvcTEUVqM19ySnr
esbgcmChu0wEiKqg0ffZdGH05/+kSzzWaDj/UDd5OztJybGmvxmAN+XtfkBE2TF5uky6UrlC9OBA
3BC2PaIy9OXdZsqwcrG9o5kgvaq773wzdnzjd5ARwSnmbWuS30GLYysKnib0tOXzMXw3DhnvIYNJ
S10WynUr4dKtfb7tJSTc1RcaJG5cwFV82TGEUW4vIyFAKPwitsGbKLIqFy3p6bS5K1q1kFjQfxh/
4r0Fg3sMJXwu3Nwlf6LODOne+tqHb1N0y+3v07fOpqvnf+p8NdkUDAqpx5e8V1+wDMkDkfXKK4bK
/A+xErPdJCQGygrpl9Rv3vfqv+JtuaWWB+zGN2fCUHkP+8UU6k/MxCgEtlbtp3DsZxMJ45LS0wup
5Z4ELdM7RZ7sYEaFnDMkO5rNbBZ04FphKbKNkEin7YwdNme7oiVIC0gFJjDiMbK+wNNLnZDOU8b4
+PDozXDgXBGW9+TCF/il/H38i3sBsBQ8UV1u+qj0fkfX2HtLMYb7EsfOZd533VNHE7tn2+8wxcFB
F9oxB8RLQU0891sKvNSC2MUWnbxUvNc2N/5jUkwrQOkhi/G2oHBrWWkRct+/QRUDQqOQaTCVv7Ap
fdTsk/t2yDUNLigCA1c22xeyZacu9m6zQdblqzq6uUN335af5cOypccTRTmTvQ1nbLRvPah+qs+8
jMG3tsQcRO8EYpnUhwv/9yBqIi6HJwMw8ZDRsVsrMkXQbWnDJdfW2/KYc18ZguBvPTZG3uDCUFk4
Oktm0bEzsyKozr7qiPZncZHB3Ff0dokWgY3ynCR8dAcJE/CO9CpT+WMuv3O67w0lvCoRTF35XxhD
0INisj07sIsN9c84PxLCV6htj9cJPCX1tHSrG7wlKXsJ2E29fRAM/lHCXkrs9l2QQTwGNmBdVbu1
O3FSnGwzJez4jQxtzp7LlA57E+VlOJ0hZd05oWZi/njlzePOFkG3NlNOFQH6Z0OINwmrKLoMfB4d
3R4gqk+9Xz2w+zZcT8nsFKd2acKI3U7qPphCIULvRDEmravpiCIYqgNs7Hmq2jIQ5VyqPi1e//SX
NN8oFrXNfJOoLoKtceYe4At9XZdD+cXnQ4ZQUVnZXN0U8asuveyI8obddGvAP7uUhV/IexcV+V2N
Y2s8F8zVfKYPGP5kF9MYVsZVqoSszFSkHS7EkqiGxyIJ7dRUqLeOWqcjLoaZz8yq1AWim3RcHZW0
vLpFEaA/8Mh198iXQs2BKsXl7vKH8qs7F769d6yE34f5mJ4ANXYwVEQzevteQNZfTnDqAkw8Lp2+
W49RGisIu0CZ1vgcburccwENFlvEKIA9gOUGjS9gXgbzaNxpyc84QxDH5Ivh4MUVm5s4slvRFE5H
FlMTjo7CN6pYL7kNLwQ1tZQSfBP0qfJHAvq2kenbbp7HvoqtoihW4A4qESb2us+GqdZViKn0wbGS
oDaKhEnngXbj9fH714t4iZ2nFZn01Ddi+D2Yxd8NAHVtVt4PeMCjo2h3zLr4Mxr2kYwbmnun0OSK
n+xzV/i7DvImAcV/L7wg2k9zSpcuk/WFV0bJtOiR7e6uOtlJ235O/pTqm6St3x04Sd//T/Kq5YAk
nXl3TIhaw2J1Hlrk29ZSMp978Q4Y6hUrFCovig3J9qdXS61D235dAOoAZfjDIZoqEToAu1uh1LQd
HRnt74jkMxhiZs5h9uAgzVyJ8TEVG9n9B/BKiIsRFqcbglHuxx3gXoTjkDR/RkEojbvROmlqU6oE
Pm88unhuFU1BVUIiz92YQqupzzQwaj0z9UliZzfOttQCm7S9AQdiKOG1KpNndiXijH6AJOIAP3kb
HAEq3I080opE4o7kcSgCjF8MZiWYtg2NxQ8af54IGP79PlIvd8hGLLUB8U3TFg/L7nBcgMP9Kuex
upAq059Mw4M0mF36e9DehjCTjxy9Nh5G32V2uY3O/lC24yoHBIZqybAWSwG0jG2U7vaZbl9a071m
0q2MkyyKGSo5DAz5A3Iz0k5ly2VcO/7j6KBsBGp/w+pPxdJv3qI8UQHklA0knkADtQ3RrRCTaTVI
1PxCnQgBkz/bwZSSebnqLvW7DNDN0Ds4b3YCDjSD02ZGcwY0shXE4vSx+YNZ7760bLGaz7u5JsE5
bUaRg81c3itrhD7xsAtfGktFiwmUBzzXh0V++xhtpToyB0IbXPTYIF+/ClL6O5wKJaZgLSLn1U1I
vClubJsCRxP8JepjJPlbAyRlv2yec5q1vjUniGFZBlZ2KWU/yZ7NkObEYslibwbKvANRB4fnsnjS
ke2Z/1PykSNkDmPNGl36EqoiGgZy0cD5Oz+ahbHatbYmbbMN7TkTlm+PjmO9Yr5n8DqzdiaaF8hm
JHd7Za2tBeLw2DNJyPbvdjehWlxIK49TOEP69Vi0FX4RntkjC12cdkFVan12PB+g6T52m68PjbeH
/VpElVDblVgkaXbSDwFTgd+A5zAvGmIcR+5/zEaO9sYzz+SyVjB9Pqe2ceSc9kiW2Te3srsMdBfz
XPhq2+cprhJrtI94GIMFu5Nax9cHBAHCkVHbT4ZMd1uu1RQOA9QiZk/04iT/8ZtqeGLawp3fQBHG
NBo4BmBX17Av6d71R4vQtudHTP7+NQNHoyk/x66vfgfTL3hakbsdNLR0t2CoZp+6QrtQlBE7E99f
Xd8Kx7PvjyqFnUrELb3Zz8gxAPcAr+jT5XSp8D0cGgTwQUyLSqQOvyd6I2nQeHzgl07cd7vlT+ER
j8Yb0nrqsuQlT1M3F+vbcR0OmR4sjfeAscI3EsTmz62TT/NoMRMvc9vc40h+N72B7dFRJQZvTXw5
6zpAqvxG6EEkry07AIE9YM2X4x4Ez45SuxDVy+sMSGCIifAlRtz+rrl7T4sv2vfL/RZyVazUtMqF
vkLth19SP5bElhhXYb3RN1mPm6rSDj2YqUZEv5tJAm/obi2+7Yh+Grfg6yzg2g2q5BbgN7u5dhqj
gQVXqlyxYkS/cwHgbKguUSFWyqyOde/AI6fBihQ0dysRbmAeppCRUa44IuZ7XwUaxwQE9BNEh38s
ab7rUB0Ve+azfFTHm39souAk1R/mcZs5pDROM1YhQGMnwqnojJwGDvRupNZLYS0GM33Lv4DnU/OI
HmgMEXD0JG4kPqXfHYB4JwcvSkGk4YxxeQAoLOR41ckGIjoC54LQwNiV2f0TVmIb2CveGottHAHo
TPt9D7Gm1NIWeTLQDJKpKn2fLPlBq2n4w70LSsmXqlAYNhKlTV9axBm7CMi4zJ0YwgsfyNNm0ROY
lpt7rg6zXpbSpCAr1b9M9UHp0eEfvRznTNA8nqBi3Mwq9zGSCsKJT88CiFvVM2knfKB0bUiz44Cx
aNRpaCszMjYRkeqfVYR7RMaZREfPcGZwcPCHJTIe6ftuCMIh2jx/FU5QVP9a2J93yODia5PFx3h3
5vzQzUhncssWpSMaTFBndzUjCAYljpAyl6uoQ8Y6QL9wlz2JhAcus6CI+GcT0/uWmSW5H0Fgb4Tc
kYi7xd9vmXWVo3x1oHv9N00toJ2SHYCC5VFZ63vXgTBsoYLrA3u8pzPfKi58mfY013t/UNQkbZ+X
5qkHD2+h7KnmRgc/rdhF8KIOZMBsvayDC8lacY00/nOmCxjog5YVa3x9a+qFYK/BvA3ukoXkG0zK
zCOx07/KtBFIR5SCKOvGJu0AJXD3WuuBd5IcSXfb2b6/tvjnux8xBS6OzzinsKnrwaYzlIWfPyJ7
uKMPI5MykJttLJiP0A68NJxEIbSo9sQWP3ZpFErL3rCj7SwStDvzxhxzo+f1M55nIXUMl/9qkFOS
FIJblpYSIcice9NOmiB/ZpAej/6GuC53td0K/09x32j/x7hKQ4ynndDpOvxM7cbYJ7CghckIxtQB
NaM3rssVdjxrg1Ubxn0LKdJ/YL0xLn1Esh2GwX530K6EhMAAUAhG6DRDMwpaaXFF/hmn/rbaFjbZ
MxGOlvXAO1xTZIEyUJTZdHMrnCdSi7hUv6wwmH6vXBi433uJUVZ7/k9eFpt9Peu0qTBRgNpznzpu
zkf5+xWwfJV5DFJ/GURU1Lpqkm041hQuK70ayaFZD5vkoDUu25YdBs7ytq8MZWKRVhl4mNiHKqVh
d8/Vr296eXfFyfQ7cu7ZJf62TH2v9f+Y+sNKnIGAcubgtbA8XtaqFLuF/T+wteK3CsURUOJur+6k
rN/QvET/tF+ClIyS7hl28LnW4kJhx2nR8/+Up8aflkXbGPTon82+A0Amn699phcW2fx6WKH6iqe/
QXSgxK71QiqVCkq7prGNSXpOxToxD9L6+6ggYnKCRlsz5mUoIBVwIXK8EeaHrSsPQP6frRjy9620
MlSPorTE5GEdjMf2assVJYEIxI3rzzB0HKPakTz3ML/RiJPH6R+rrQ99x835n5wq2dkbUhcyQ3K0
0cdkfdcZoWw+2rmT2SdIifoOMXqMD/HwleXR5PN0oJ7Vy8HDwDO2o5D6jhCouY/nk24mROVsszAa
BCg9m/vTpUJy5nz2HLNRjP1SnPtUd1ZOtv3oyYPpn03L49bdZqKKYxdRPqh3Cffj5BKknkfnThFX
Lb0skBS+aOO1InoWN6TH20rLXmtgFPmq5bFQTE9NT3RKleyq2RCqntdRYTsFhStWmwD7ErkPJPIc
t+TH87MBFN8SRZJSOZthYZL2iODEoIJcntAkfX7NDNPBd19BQuRKuECmjPGfO5Pr+kSHF968Hqlk
I37kUI08RIy91NnQ9xoREjPhl25hG9yz1wK6c5bqEilXblyBAkwSDTLrncEjM3d6k/EVe78PaP0d
FJjiQvy4F9PtbJrwVkVBB2o6roXqukjJWnowj3t42hQwvVqxGR4ACWFOt9VJi7OS2QRxIEV2JAVd
zl4r3WjshjH0u7JNQ/8Nju1YKrfCTgsH7TBPwfSP4T+IEb6aWwQBvtkDe03ea5XyRkzepHZXdD5I
Gbkq2AILdE9fIeTRLiAGbljmnenQzZIvkSzMlN9iP1Z+c3JuMrwDyqPwoo9jhSg4030mYiQvtLRt
Lv8fl8isicvMT1R10Wuy1MLe4cleyWUUioBrp2mU+IZEbRLdHIfO6vcVActCm1Nafa9j9dF3oZH8
Az8W1gnvdkeAu32Zk6TEHsfgML3R1SenQTJkocYPTQBSRB9NLgz6lRNgXeN48VfEEGApxUm0ODTB
y+IYZ1JMThPLaqL5BErRkz1os4SNvHfbt6tiCVRRXSgX7B7yV1gZnZxkfx8kD1FvVa9HxPCU03Vh
bGZezfQEJe4xBOpRSgbo5N7ot+P5xr9ubl4QQPeVBrAUTlS2YHKI7yciHQ2Lel8zYmQRN6sObjRe
rbM92HmavUmL9T3oo7o7YXhNXQ96lu9uEHBtyJZB+S8w+mnJok2rcyjaEE/MDdcDAabMjrqVM2z5
AvlEo9em98SkznUao2l6v/nlYU8FZBDQ05JqMGuU1AiL5voLdEMP7IjFp4DmkbKzmI6aKsUVm3r3
BdgaiCAHbPhm79Ci5rwQ9XUL7rV2gDvQhmqslUUsDOw/Y25F05AS/kSEz1dE33woXST1ihCrsCsf
ioZ5kIkagPfSmYPoh+wsToduRZUzfpnnds1UptOdi+8h0RmaVhJeCdE2gmmMQ+nv6RtsNCmCGdST
zQh2B77aSjp9gEGHad/fCE7qpU5Kym3bpqbzX+x6TGsMEkOpN6wCMiENKShx1AVPCW+rXBfhuN6v
A9lmk8J1xZ19QtyX7tC07aCBXil13r3wY8JWzagik8gzpXrJM6tvb7R2+2EMEzeUCGdhRI4r0AjA
G6L1uI+oOZ4eizoJxJi72QT/jORazyAjElLVYJENgL7aIbcyNWIP9b/qTRuzqYvOsnMk/wcN4YtW
I1x+xWTyBfaUul4w/fdtKVg9mUEm5XyPfXL2nINiSr0sWhtPczPeKjsQ7SWlj/up321hIJumQ/bg
tIoCKivV6Xc+UuXPHo7Q7bHPUjIsyRSnyj/dcFhwC5lXe4khrkyOKLRnTBXLZxmdoPxXokIuO6LM
Nruld/j+K+7IaL1GH4Amy+GwDFsEgpttvyjdRvTrWj1vwgKV5XfNgf9ICQkTa0BVnMBGJG6Jl9JQ
oN+lHt2c3Yy7MmXeqTNZH1oMzrEVLO4t2BHI/KQpHN12Sv8LzYtUXmLRKlRF/7OgLxXCUfPjX/fY
lYzFFR0wYsDwNRS6qJ0FO+M6itINI+/USjrMiVTAGpJ1jbV39DUGUZEd93EMwLuq9gcgQoahj5og
ZPqXQ7osRzL3Sk+3jjThVgkfcvdazBYK59dP/hO6o2OaX+XGCFLJb6T8pyZgIGJYPXO0yGtb+GlB
/e9vWR70q0eoa+K0c32NzhDni1mVDGhXZAjxuKYB7vMXqaLn6QyTi4Va8giraXVJbEOskvgWZJXl
Voij65uqibHn9/dELe8uhoLvO7M87X7SHDnbBx4vw9QWSLjAkb7h1z/YTqV/vvejc2ZF0E5f/UCT
FHQBPvfONA7YTSGjCkvrOKIjDxTjU103Ar4/K8BQ3DIvxIUBGst8rMfWbY1ZM3ufDml5oNYqhF0V
8WfX/MngAcngyPB2y8d4N0e0hT3d35bM8ah3Ng/ufZrjrnP3aYpaKBHmyVnTpTRco/0yFqOkaDvZ
Q8ujKIb9//j/MWzN/f1qhuDP0WISfjaGh4eXhHveXXD/zIqy4pEdna2t8Ypy8Rqr38oSj/x0am/o
yzcYLOLwpZhioe5RcfMZjh01XZwlL4wABfsZNzARS/NNw/c6PQ6i0MzfVkUMKkEK1zvwJuk9YSRe
Br1rLeVoqIMIDzZESttOWSmq6mLpLFXnD2nDmyyaJt8fLw5Lf9IeQpINUuJbE7EM6+ELK12XC+DO
9MN5h97VlprJDzqGAtWTw93Zt1qQOTSOFzP9QfvRk7JRq7T1aKpUIlQB744uDq2PO+BXg4jTe5l9
iH2CT3SlhhCKhtX/DHqSamZvSYVKLQQ1bBEkbJaXyGKIOVdgKoVynZt6+8aTNdBT6j3cFJtw8d2q
8jidaJgKgWXljPj+7Mf/GUBxuLK4o/JFNMccuRAXsIpLTyTgCW76XlDXumHmqk+5fLBni4lZ4f2q
6XBBg1HToCLmRvJ+FhsxQPgiOjQpW2sEGLLDWh7JjjJQ4mV9knE7hXM4Lrdv3PisSwednl49qH4q
qwT/M9gQTJ5r0GvayA5bASs39Ep0GYECiBNbm+3BUW8CX38XfV14iyP3hU5WdeMxS4/IRzNtUtdf
PUtwcK0/ESvLaUBPiz8RggD+YUmXcJ4J8KTTYThQKUxt0iRZpGkMJ6ybA3maerMArQwK/SOC3jYK
BUyq4ymahwRTpXVlwhTlO+APt4huhlyvwP/Qz0dEjwz/ORORqxA+JUX52gu8CM00cWJxMe7w9Kpx
OY2GlI9h3t0Mz7GgLUsbPKT9ymrjWlTttoEvupm0ujnqE3xFs6sXaB46gqBTLjo+ggqbjCeco8n0
zK42h5vD9WHhBykMk1MWAOHmJOfzmcVlEWaeqifnZUbTm59XJdge4LwZprK/wlWlWO6kiY2ggXF8
fwRm3RfyOS+5x5AuO0LQ2IZUUxIcXu0I2odoChainLtSNWuk+vYAQyRb02S836O3r/t1wVoT7FAp
3hqNo8wYtpgsYHVuhJGMPMV5MDdrHeJ/VSXoYX7/ueYaiGuoqXWGQH0iEyN1yGC+g7RENlmPGxug
Tllm222Z0xsqETYMKVoatxlCLFY1UeSSprE/48xMGV7CW+sXFx+2tjQ3qxVEnnPxFlv3RMHX1bBM
7LY/qzOJk47VCbWRnTachQQQLZNspZObsEkN7ZYff6LAwwNu3QXsfbIKknHKr4b6G7XQEuC1ULC3
E/fFunlPwg2KGfAGXPQlM2gBFjFOHxw9LB3F+p49kwvUyIP1skkxFKZnPShyvolWriYcQTgfReMY
pXLWnqyjHjF/u0vVbEP61RkjbTDsGLXjmdV/uziRfy1cfcdIcuca1ZFtLFfr/Si22DQEwkx82QnM
HiSV9jqDVltw1rkfFsf6iCeP1lbsO614QX3HIPxiCsJSjDTlIJ07yyrMf6Bq+6vZt3VDLOw6J5/K
oMiR2aOLTHMzk33BWdgsADLyWwCTDfVpeqCBDyPRb+3/eHGYBf1M/UudSCeXgIqIFVLEEe02yP4w
9z09shlUpkIW88Nd3ANkKNfouDIvQn5bEc7zGM3pIjz3rRTiRmKj+S4Yfhx3yNA8O7SlTIVpV/or
zxt6kBKsJilKpAcn6gjLY7mf+HIKsCJgJMn3mD9mCk6GCizd61+zx+6YSRYKYBr7z+i0WEW/9+23
8SCiP0hD8fUjOYJoUhBIdsKsCTFhWatxYi7SjBfxyoMH6XDJ7XMgHsX0N0xdqPNjgcvCVQ5OPbp5
fH8R5MVjNdwJi/DFezYOLFbLDD/e+ehmFpgmdkpgCHqIveH30/UifD5PQsSQPMm4eL/G8UbHP9Vf
/xtOldf3NtYLygp9wlnLL9qk3gg1Aql6tklAilcKylrFbvXDqdP6zYH/KiuvR00eEiPX3DvSm5fh
ahJYbZxty8l0Q0ptNAoeq/KV7xPm/8p55D2PmVNjUWTaK/0H8GYdZnoVsb37wmPN4ymEH9CsbA0a
VrIFh0bIjJCHyo3V5cARaChd+qAmQ6KCEg2Iz5mFRI+vmmu+jUKYNORe/2IAuPvDQugT6NtvglbS
DA5bGeRbrxWhlTZGKE4268Gv9ldpUqM8xauaqAl6IPCOp1svYQM5DsY9FQiLucOAeCkafoLJI9bW
gCGM50C39IdIjgEQrW9/26eREBrGHwAxisOjRTVhvl6hhTYE9+B2GNL+zBZAAn0F4CGMLiViEu7l
Rp98AqMCK9lu22oahrWAOhoHzflgwEuAYxnB2dFMJBfqqi80bn3558K1ddjOzHZndwiFd9tg+9u3
CZ9IgGIjoMggWBQKyY5fN0prHUuRfvDMGOfeoY8ekO537qCiXk7v9SukoBghxrg/zuYyNrgQ4TPE
oM0G5fOY6miXA5F/rq0zmrWJxp2miouOedlRbIFxZ010AB0Gogm4Le/CEs7sx/f7rm42wOLgLv+6
QBNvoZXsXU2CZE52bUY59yKhrT/vZh0/sfngGUHdE1EDH/0qSAq1v2OT7XpcCNyFH121jNwHOzGy
OUd1onoyI1tz4NFiZLKiAz6/nSWWMxedsVBXeRChkuMsOvIjhfgqJI8FsVe5aJp8N5wbu/9uHZzW
cd3cG2wsmH3zcMph6Y+p/Sqbw8NOalMWxRHVlijF9ZSY5o+VbrYioAe9uWNmqVTdNPjc8oO22fde
VJLPCP837r2+oz9OgRw2vpb9dbMfIsiRorbvwFsayBU8rIjmWtWu0IwrH3/oPuGu8OcA3L8z0b01
i1isqaDC3ROVQNHGXyYqEKAsndM+T5L+ZGdWTnYsh/xjK5saBD4MMOpG3+CgM0J+fL6A2JBY9UiB
N6MR8ni3DgFkm0GHAVNj8SDnQZ2wffl+MdaB3qH4a6b1FrKCor63WaIwuOGlxhQ0BezVD7xpBLd/
HQyZsb6tFxNGu/BNuN2fDgzYFxVDybRPBD4q+fGP+cJ13T+sWnD83cmi8tXNxhoM1g4576+ZkHti
SNJifl4N2EcQq86nw3a908Qp5GkEox+VPu2UUZtLvwpSojElK/Nz/m97ck1aA4RJ8r7eaWCg+Pv/
iB59ZVB/BWXb/9OlQwDLTjUgteEJwH1+B2c5q7aYzkOPON5Bw7A5hgE1sMqPCG41A+VE1ERLZaCN
xz7RvPk6nf8eRJTR4Rn3jiwpcbiTBKzyabjXW46MaMdzKw1hpAgstZCDHhga3bRdh1RpsVyQ7RBV
DlYNzXfDydnIQhJDMw3YxcuJ0pBkWZE+W9oI54P6M5KHbHHbSi3M88QCgQcN59bsa/SdrEKiVLK+
7d6Zc6OwefhWYGksayfFRahLpDD4XXVBxxa01o4SFNfnTGc3K/toVqH0MiUFnUlMEy5YXqQVoAre
ZPRRcdN3fVb7e2bdtY/VCC/EE/aFqcmfavDZCeKtJQIIDevzfi6e37YkIsj+2kNi7HGZdQZ+poDe
kO1yPskjxKiuM3cuXGAtnnhgeGiFqhwX3EO1kylIo/TjZWnJwKE9LkqaOR/z3xkLCHmaJg5xN8xf
vg373Dk7a/MChbITiMteq//oq+eEtkhhm690bmkdzLoBqlceouW0ADgYsFq8384vIYvUDbSLPtkc
ura16AtNxZoCASBkVVNiQmEsLVwSWkWjyHTr0vi+/KU/2idgiO6MvWXDtvp8dcjIXg731tilcbg1
iwlPn51emLaHsvlkLVTeLVl9uG+5AQ/yc6oYklFVKRPj/NCI48xAtNMzPQaTEUCds2BPdEQ3LPVr
OGaeGygwVIBc1YG627BDFzNz92smDfGEHjrDyCwBhgManU4OjimHu+cCrrtC+0bxgJX9vMEGTkb/
zat+zLv6yktXhJ94XYw6PlKESI/bHwXG7KG7qy1OMGsOX/R+V86LZWBHF52rJVF5iYt0En6JwM5c
20BbX+BoJ/wv6ZIxhHxus61AC9oVoUsy6I2SM998eOgidpGhqsRuiN2I9eYguIM7iOS4XUHBU6zn
L5HKC6BTCnuSlhu8XSy2Q74ECDm7bOI1MUvojxd1U8svQ/mgbOMN25blABmBPy1HVOYHuEmsCnEq
2A+GUXXfGUtr2sl3bkSrfql2cYeBGzMwJb/e9t7zzLfPh8cAACWwejSVAlSuOEPB5A9kmEdm5NUj
IV2FPY+vb4FKiPA1kSE2qkQK/slQlnzB7Bww48zyDhhP5OBTibszjKOeeaEsIxYjX5tQssIqpCng
D6wPZkkGjyNgkpQ0H0tXJBOo88SK7gRRa5PSwMGHg3tAwVeBFai/cLP6rMdhXpgRdJhQvU4dL5Un
h95kEY26wT/0sDJmjhFDcdVUx0iNTWVqWkuCo8bNnidhlJ2MKmwdW8ZRMZIIJQxw4VFlrQBBH1/Q
CmcHuz7L4RbNZSX6aNv88ALXtJ735JgFsxca5Qnj6DNbu9/4H+JavRyLfS0wtKryN9ZfS8C7Xdid
+YkhJ8BI9swWaBfqCRCc4v7jZLzLHmDDhSFP9MTbB7FUvhhr8ie6xoQoZIvxy1Agpq4cXAO8g9Wr
XJoDKkxicsv7TdfGYGyqqT0FXBinSXdYUtKEGqwVuvH6iSnMg7/EiBtFjJYWgkK8562Qz8I8bZr1
ieD0Eowt4H89m4BZWfx3SqYfXroHv5U0Xs24UljAMxkCHVXujKa4Ydedj36Jml0eBNDKvICSTwsy
QXRHMMo5c91e0Lrht1QTcnt7RcFKqs0UtsrdJ0shXw8nZVVXshthuUnAws4ZGb5qXJlkceHtSDef
y0HAE3WOGdz1rjJzv94QacmsVGR7p0KuQh4UgycDpAgToZ+NFQlAbji2ZBJYTJsbGrtckVjet+c1
caiuX/Wsz3rtv6Fgb14BfVSULyKC4bhhhDsM+/iqBkzBNhwGbukNdsAPYSYvqqJ5qsBawsCRkWmZ
tunS8ZBm1slnfSswW7+kZnOHLfpNeW0ZUva8sskZHGdI09VFmnzpAs66R1RS7a5+1XSky6RsLeJ+
xFmZhSCflzLGkqaH5rsioxOJkj205ffkiZzfKZZ1lUyb11okGUcAPDO7vR8ETT0+bwEn33GM7Sy3
L4M2AG/cNNdE8nMiwKjzttbWG4wnw9ne23KwH7+j65CFrwIinZ3H8uhNQXjVMRb8CPId+P+bQ9So
PXyqiFytdBO0mcRHbx1VasQ+uUNiCnouTGBmhD/efzQgmVUhLCJ5zmoGDiurYf+95icsE6FFPBPm
31a5RoHmMn62Qira1e+btPf1PuUmhWzoMhLKqCxdXi5AHKxlVOOUrBHj5+2qhkbQq96cYMgS5B+k
2oONHdgSK7ILm0fe71SsA/9WMIUpMR/yfEBseKk81DjxOxU7nQu2Q7L7Hu77KhQrxsFciE9dHsdH
D+e/HKHNkJTy2HdOIGCoS9STDenrRii/jafe54cjZo+lyQbZfP0VvUcQqpnyD6RrNH4/2e/NtzrV
yMJh6xTlsIQeFP7PE1Ma80/2ba21qDQ+FaUA1Pvwb2kNwWAjdJ3u4c+9DdNOJhadZPsbCPRBctZV
FakO73uwxLKZVuW7ys11h5Ms7HVVJRFqkeRLo5OFTGQjSjKb6I3DQWHx9ClmN9+TdpX8s95UCdzf
l/pQkiqElp9rdDp768B+400LAENpF9hTtf2FIBkDUppJ4GJKmdK6/6fnC16XhGIHxr6r0JFFBqZV
NP45rXOVu2eqXUr6nnGyyow/8B7pBorzHlIyHMrJ9dezC9efUOu8J0voT3f7ULUpskAlA/zPCLbP
4wMPxrYwLI86ngyyh6zAeIxq8o6hdUpDQ94ZJy5AQTj6XIbsgYbURVrPSspiuoQ04Jiiv4THsdkU
+NfwnumVRICq9qg5oXof9uF/0jeFK2YPF7y/YjAPqHTsGxYq51f7ZAGgoT6FP4DkoVqbACla8hbf
/ZpBOwL3V/+psR4OyNcDYzK8SxdppMiiHNph8oXY4JPqeT1XFUkSI41CPzmMk7gmalMCKB9agOwo
pi9B72FnCsdiESAcRZW74+46Uy58fUz6CKf62lWOWDDV6LKNu6RclD4s0LFAksNLB8WEhSAf2lnc
C2LCwxUa42xHu5llJvGQ4sWH/d/uiJHjnUOtmVyu5EZQdHUOQ51QEaYC7v9BEvveEzFW2xjSLIRo
6S3MAC7CQ75MwgBzAciNoslU2liuIoXl2vItFUGSKXFaX452zMR0HNOPt+93cIxWsOQsGE3ajYFt
PqPckvFLnCbLyJ8xlv6BhETDEcw2e9KwuC2SQxhckU+MoFEDdalmPB8/gzOnHuA9ut53YaQxrrWG
kKIXCGd6rzgnuHM86Kd3y0O8mBLOpFqhDvL2yhu4Zm1h9ZHCSF4vkznb+TdyILwyiuARVdMbU0yc
4qv1mocQQB4Jle5LgVfHZUvPdRkUbyVjiD388MsSyp01aplqM8iZ9zqv/rCVAUxN/cJCnpt/ibD9
CJA4OKtpdQu/iJjC6flApOFrwwSkI2C2GkCnrZtzFUVxGPkpR7fVs4yxw9tBd755SLxzNoWICpy5
W4H7Lsmxuqd3+uSdZxJEjHsRKPSfKYOZ9xvJ4lg3NPLS7n0IVz6fThrDWCSyjOohSjgqvo+YLE7Y
wMXBzcp+WJyJoJqzSIbkF4y/6yCCXg988ckjhjHoZaVIeej0gzuTXVmf0NyF0E8jZnt/9nFhPCYn
a+t3heqhehtZmzP3nle2tZRaLwr0QB7QLetUBewWZga2HvjjXWmvblmG4DU9MN0o5TflPWCZVUWZ
q4JjFv+iQfk34KhoNUTmBp4bVpzqX8HXWTq9AZwZpr8ZXxWn98tG6cbtJTsjs7AUZroKdLrdTeK5
TSm45bqoFjfkOE6/6Bcyj+h3t6GnO5m5ERNW+mJHpSLg0vAq/d/mfW3XoyNiRVjBIMNdLffg3u6d
NuULXyWHnfHX9qSjH/rVuX04ucwG35KdzOCaZXlX19hPQIRnvXjcmWAHNyYg021U5QhsRGsAVwmW
7s/qAlDX1VICdAn5X2H2T2Pb+CHLqIgUhr2zV9+vD5gw4CKEGLFAHk5UwR8NsfPf24WR5h0nPp/c
pvmqzwvTRCh5+ZpmXxitRB/0hd52M8vcGqsG7u6ZAslPwrD/swRqOn43xICh5nOAaUpj4THiacB1
Uaow3dwTsKgYVFLoVWKuw9X7q3q4+9CWoo9H4pQ6mvGKRBWgiA5Jp48UTfHz4nGjO0R4NEXkIAFU
MxLdTxn6I9Zf0uACbZLLPH1Bh0kRh2hZEMKkMlqv5bJ294I3+52cEkg+cc0CU9qC9mUa7QvRMPbW
jMicK/bgr7szu18kJjfRc/IgUECrzTciZlt6kgQiQG39xI7ScjAanlD6GaSHTk5TONT/bz9Ygwln
GO+pJZu7VNWqLsF44PhdbGA1sVYUsypaVl5/opisXeqcrsBNDV8GlO6GlNPMekDO3fBPw8UNSiDC
Scr61EJ3VETSFSSP/xiB4zzMdnCPTzHb+5K2yG+/Wcyi2yMosaIXi0Zb51vZOsmXlpE8XmUU8yYD
YfyuFNwO9s9NBNzH6qWk1b1P2e55XhGhhzc1RRZtPKul6F8zWZa2pV3kwLF7eiCWojrrIt9nQ1OF
WF8NZJ2wpKK/9RAXAbKzFOodtC+d3ySNhj1sHqFKkcmQ0r72J6dIHab8zlyx0s66XIuMb+IOhVv7
n3ArNwpyb7krC/9fqHPyRLdz0RwfIO3y7La99b3BqbdEsIWVRPeQHMTYWWFAirD3SuREFHnx7vdD
XGk2rryl6LkjQWHrP+X+oji0/kU9gn0ifnLBl3MJ/mJkQpVf4dmbAhFRTM7vmp5vJ6n1IJDiS0Gf
z0q9UrLSrgxBJhkHY5eEuRoHr7TZgLlBXGjkh457WA/qsgGIh5qTuDn8vn1QV0gthy9tPrNpLGRI
BrtYOEGK89t43yqrOfKJVsGxuSLk2WBKKwje4G3zS4vG8ebKQjW1IhmAwR6XQ4PdCmDOrO6gXtNv
InroeM3VtKPbnXGlkM0Qomjb4k/FM3moePm0MKzW1dqFBfSjYYXox1YVcO2eDpG8tSbhwgFDwgiG
GstSKIKvinXcIasXuzs4s784H2aj0vOS3Ak2txBKSJK4emLICsHFGM40MmpI1/8ZBAXRobqorJzX
3pzMgBI+8c4gYsqQVhVrGnVf+F3xFeu3CcMJGV3JxbJRbIxdZk0c0a1V2hiB2CDq4K8NMM/MYa3v
beXKAF6zrYWTA6MdNu1oz2vhL+LMEB0T2SeEN38cStupwEqDdYP18JIZDbqkVsOQzx2Fd7YFhf9O
pdv9J1cXrX74gP85C5vsvKxJY8eMwr+w/Cvdu/oA/ZuOhsJgH2Swa/lYB6lwQrVj/X6/1WCP0cOG
3sLGInoFePj35QsSxtOaMFAojTNtTgMUc2KHFjY8CrmdOG4p8xbZzha5Cllwl2K5W8gsgi7ZhAgr
LldLrYL0VP4gdCKDXCbGbrVJE0sJWgCff1niBQrr+7z3XSUTZohdpUWON6l6pT5fON5FU5kCCkrZ
xIO6SpimbffV4qA1KGUHUI17HAjAJhKp9y1nFyY5HseFkX44KpZNUEoGY656WMKd46c9ZD6JNOp1
SCcwEIuf6hyiMNYSO/ZEJy0kWqCRVfRr9JdcYAbhtWR/a4Jvk0r81Paz6j9qDQQXpV2TFVvyzTEA
V71ztMHTfOVEaDlOdtGeyUVQmJIsfwst/EnRB61N95pWJwzFO1m8hRFUck3aZEDP9Nvs7JM2Ur85
CCi/T18zYCJEQWmjT2Q8bZj2oqJ6GA2FJgX7kj89zmiHZfKlKEhNSt3uEheAi0TSqOE8QJ4dylXe
1NsV1JQZFQptk9+cWEw5CeUij6Kt9x3OFsPA8YEJ0O65HMQnRuVk8KhP0LpXy4rIFozzSsWOT97y
rS/Rv2AF/q0HMogPPozuEnQp8g16zJS1YbqywYTwIpANd+jzoIca/rIqi2umO4nyB5+YmVBP1nZL
UucIXWrE6pS15ZM13UJKHKhOSbpzMVXuK7bNaFzDU5q9Cg98BM4lQ7Z7n4PZEbOcon4F/hkIgWCC
vyWuA/1LktZ5aaM3JV7c/GdJrRTSSBCufqT9PjSYoE3LKR6VWZ9Ffv2i0C5Eghxc8BFBl4NNTCql
KGgpVqKfuFye0MFiAdYDvuPoKG40CQxUUhUgEBWoOdSLP4o2VxBjR6UxVkdWg2DC0681l1vOF4cR
UKf37cs46SLSSMm0nGKB+yHhupca/cvWL7FVOgSlSL7hM7z4PaTRGa1gm1PENA3WUZK2DMQOWVXQ
QOvl/QTEde35y1ddmCR8pqVnMxpHvQqR/5HSVXEy4KD8DxX0FJAX9injjKq2G1c5M4XbefPDK24Q
Q0Y5YoACgTQZI4wEDGqEHOOxldqqgjFNy+ICKmXCdj5ucjPZevlgnrw3pgrJfCJsjdqVABRpn38x
qHdVvNJkI96l0FDTEKmDEw5GiaG5IuFNGEu04NjUNVoWBe+P8FuO+0nw0vbj6k1xzw+GFbbQUSSY
898h+fTB0RxKIjuYqYqlr/I7ex7w7taXGwSWdbbiDvJ65uyoyJJ/4OiIHZ3Kb8nbUaSm+qaN54BC
d2OyI7gMHGI6HF8vKPecoKo6Q6JuF8cgcki3YgTKvfOUl1yf3r0WA9fiM7D9TMgDhVsm7O3kEZfg
R8+OzXahsJQBdVH3lR9vCe2WX6uFqbfBqDx+/M6K+wgCJkvzU7MxKs6WcqYQJIfgZAFCCpl7w1oE
6oJf3Uk1nHBxBD1h6Ps7l2R5q5clrNKATRmH2sLmifUtBNeQIIR3vszY8Eac/IqGN7yKqugSMALq
ZD2jb6+mCFj+Ad6oSImXAf2M+IbpGj+kcC3KgCLDh+8vBcuErC2fbYBM/0U4spgotMP3xlpuSq6H
mv6AiGfkFI1wzn1vS1E7tkXQkr3wCTKwglmRdoTF3M2Gxd7+YToLbxXK+l5RW6u12E8xVWxiMWaX
xgVrMEwpKahNIUMeLSbnORF1/vv4yJby7AhiPeq+msGi9gbU3ZN8Q0qPedTjlIuqxVrd+hHZAnZ6
KFyu0otsAcbc0Fqkua0Dx97dreC7RRxP6yeTU56SgnqRCozQuw40c3A1YkERrv15/QF36SNqddET
hOY1EY2CKv+hXdUv9tDw5A/RygxDuMaNJiwDu2Q0A0cOEnNXkattRiptwqpZH22LCXfi47IIWifa
8hPTWdjxc0QL/aqNvjilerMKl3odJSPp89Xzr3JjdKC+YLl3sltdQC6DluRhO3uotfy8d9QF0MZ7
hRdlVKpewqj6s2Sk+9eqmAJ8N5NwTgXfHmxZQeNw4M+Op/DKySWmqx138u8rHKdaqGRNqUaRxsZp
Wr5R7x+DqwifTbW0cKwzxgOyogPCE/y3T548tK4Vni39ySUZeh/yki58r7UgKT65iWei5U+BgWBg
OjIQPhmhjEXxan2QcT3QE8kLLYYece1RbIOWxXCHluc80B1iynIdweovkZzUy/DxYWuaVI0i9Y33
loZ/nEygc3zn7znex2XzsFGtmUkzCPeuVLD6WGp4VjvPeF+GczzXlmW7BHF/uTKtED0OD8Dbt2HI
XRzbUtoEC62XWPtGUfxFR4ERzTnfgd6+SQ2GRkpU+fkw4fo6tn6AcxIsxlqKiftXj7QlAcFKDz7Q
Em47/KQ/8+MvMtKa0pHFJMAZ7NhW1lutN0z+QN/LqfVenYAZF6/oEjZZFVPSQPka9HYTVzOiWFa2
vNylBZqOaVRecT2+qp+OsDvws73Az7m6yTqM2vGj2UjN7YwTspVSaLLMd17XCevYwBFGfFLq/OZ9
hkdTqGGc1k4v4plIw7NS1IiXO0XWp+Cjkz3Cgy0QPceSiyGEIF/kibrmozUUM5ISfRAEOy6gYySu
sc/A9FwIbBT/ofCk+x8+tBjrJAo0ZAaTjRB/QlXxKx3qYBqIMXQSpr60kKqFJeHyvkQiAj0DtdcG
f/lLhNwW2M8fW8hEEPwZWuI8N37n5CJFWP4pesfTcboSXvznKK0q6fLlZQ8xbJU11zVTmMmOfndY
m26usV0XDaV5yq9Y3/rRuE6P6eexUXMoYeXZ4xLAwipceAWH8DVqKNKaqDX9FqYgKKjcIDkYO3um
QxwNNcHy9HIUW6SUxTjUVesIl8J7/tnxCxCyNRdV+/TJyf7uNkCTE+64UNH10byP+2VBaryqiDlJ
zT0PnrjHuyBZzr0KEipqmneM6K7DEJFTxgOFMdRHUFTLk4W15x97JhfHxL69fLtc2XZHuTZU8stQ
7sTf1e0ivP9GV9BP8682mXXK743+4QUrfu7rCp0c6ctBqXRhf/Z6+tZCKw7H4yRDBkxcIUQsUugC
W6kYQX7JfD+MPCbIzpPudlss8erYlYY4o2veEpZxRH6+di5MfDZPeyjxFTE96QNGjHOhl1ParkLR
2mEKXa3KZkqhAM63nx1BG/sEtwsd/XvsbZdFh3C3wq2KxC2E6MseebAsuhKus7QQYPdyBLdnddFd
OEulJ0HbBN9jb+Q37Ua0IDH3RW8GOOIjbPxhtaiKyytPH3J0J93kJF09YwAd642PMKI3SibhK2Vd
4XvL9+DLnvQ9tI7kwzLISND6PuxZ6EztreShRiSWX88MZgTdH3N7gzzY6XlxVL7KrRQ6ygqsKl4u
FAuxjDZoC5lUfPVXOttCuEjmuxKzRIemZFUDQcTawzXnajersUdQIiLb1rHUM1tV4oujU5bHbV8/
hyTjAREHKq1mzf454SPITkCr9Ni6ewvONAOxdWXSYZug3oqZu3EW/bEeJZzGhcb/jLRIAj07hf4B
piu4YNUr6mIf1pYQ3FrJ+Tq6ZCnJINuOhwbf3A/bAo50hE3qENe4MHC5U0k8gQhk7PTQTzB7styY
Bvf2By19aC1D/wOpxJHUdGCWAI8iZX2v5MB0WZGLLdZ43iCh1FFg0BAPu+h5uZ4NLEtRKrcoRps8
kUptBrG/48a73AtpU51Z+WZi4CT71FhCvBipoSYbfBZZJUtEmdgyoyrLvHZfx1PV3ez/0TeK8MR8
Jc7IV2PEV68e3KjuspVbuCh1XYoJrGl+dkh2h3STossLa7lqn7UikRG3X2YSoxKFBpdpQ1yCbdii
PGBZtBvdpq45eL6A2uZxtB6IzAfSuiwf6zpuERUkkl/2pE/lHbjkz71asV4/sjklaZXAepdS4hhe
TiIIjjaepGdf45CqWpoTGDlJkefFDpu6P/WtBpcIyPLrlQ6BLf10nOXvtEddBUN+rPHin5TnsS69
ecLWVMtBoymRPm00Go1T/6JmFMe0EHGGg6mRlF3PR0z+UeS/rOTesZBQK4Ow1nFCmL1wYNjIL9Xr
p94oe9tk1JNwJprH8bc1Bkz+uc/YdxLb9huuhtY05CxUWD6BnAL0DBdGb7M3nVv7q4gZp86uxBQJ
L30OvwA40X9TUZupem9QK31JlGBWcWdyG1GaGV9J9oK27GZNk6UZLpd0HVkX7ZMGU5hHk4g5EpXm
YrXptgmzdPsuPIKJbMXnWBiXFf9zj8P8srBk/3vcjI82izGV9oNlt4NnFfAuAY+kEMeouJvoSaN6
gynt4kB77Qb0gG7Q3vlV5pq8RFYRcfxbreVKJtUzcY1sflk3sLC49yMKemW1NzDWofjNZV6uibQp
eRVvF4wzQ92+A0zoa/uvILGWPxUxx4K9euSHC/EqBnv6jtaNnJ03hOE7TalTY8I3fo8XYeK2G9Df
o8WnOItSbmaxiJ+Ws1P4XvPEE5EHs23tltcnn6EDikb/vW7f9x7BReW3U7IWpw0Q8DAwb4ULso/u
lHEPlXFIfyXMyhnexJRRk0zEFTYz2zBHEVEv27jB8ukC8lq8M861IWclCUS0YZIvfYYaxB2R5xZs
qv+mUYO2wdEPHDOJlqusver8Am7PhgnRFIvgOjq2tNzWF/I54i3glfEH6jIlST8wHksFRMsQJNku
n7eeyVkb7HBgU3Z18TQQey75st8Z20XzzGk58RCsf4S9oqjW9hULtK57+azkALmx5//TCWejyHCF
wzDaGWYWfMQ0WVm5C4zdOmQZvIR/OFcrQx+vOXhSaY2MnI4oFx301+8f8SPRZcCVeBbs0j+0SVli
6bdPHIdIdqMGbvHRy2qPSPlQCUEstxusGjkvHYe7cy3LUjgye1gj32r5DshnPCb8/siv9NAJpnnG
KjSYTqy/7wd5RM/eeXwsS2mB0FrnlPD1sc98mT1KD+pleWpZYjAVQYzOUTZOKRNSJNrAF0YyI3ql
aHfEYly/LpFbGtyPJOuj3yG2oXYH4MByEj4G6+B0UUMLgc6EBXzdQXld1mAOoEJLz0/WNA+r+2We
NHit7WtcJFGc+8qRWb/VnZCQu1F7YXk6jzGWg13ZWZ6Mr5PP7eXJPK6t4R2CzV3SVd5uqZXF0Bpp
+PT287GjAIOl/JYXvY3xDxNZnwi9ZwvsdCUbED47XRf2LQYuqlJds5UlmeAKp/i/rL1J/caU72sJ
AUKyqbjka4n5cS34XAb1qxDNo3mR52UPT5cXxUJk+tsVJXQ+NdWO9W6sPl0NTvhxKa5rWkDMOlXF
3B7grYohThB9ykpTzmyP4iHMBREaKk0yCPrShdGe+Ri0jTgMVuKYol5Dsh0mISGhedEoC4kQEGHl
4RU/BuFKR+BZbuojgCBVhaQmCcQA26x7gaxaNRdPy/gZkG0n1c2o+hLtjYmQQZ2aTQtE6h22Jgpo
eDtN/haDXn7r9VvHCfzvqifl+PIL3xuIpHLEx8u0Slns1nm8GVwGRxeg3lQ4UHKrcWVUMPG9aPoL
ytrDkWn0JNyz8dCMftaiTjoaMWO58H6ukworwa/SVM7ANwBdeFcY3HEQFSpLAE/Qr1iVs+hrZuiS
W2iGB3ZK+twUVIDV2YIEguQkt3yact9djf/BL8wCgpK6HgRaicYerp23RPK6duKLb08v9fh3n5iN
RIx354xb+hrPFXwLTTkmaV6e3C+uNL/3ACzpa5yvujDQoFrG3hzUwyF7C91XJ1aMETm9+0vb8MyQ
zmL/wzcmRnNMZNoYXvud0GvM8Xrt4iQ5q2yuNgkDg8rGeEuK1NgB9n+X+WlodauQHBPsMSEdQ6l2
51nvxtKGbnp2+a5zB5QUXbn3fFb6aHQj0K8DhqDe0EP0KVLGynFMSuHIhfjDRyd8VcjOYIZSdDgE
+deYasHFmKf2s1Yc1ZeExC+mwBKHR3Qf6r3LzIQ1yBAkUXROePCkQ/MCn5Ns3T2hwO1Vj/ZKYxWw
VHj65gDGlssaAPlUECu6SRgJ+e/zpw4CWk4UsIH3sg24JT1VaHH2zfwsmmzRg7wENnUbrF+3a9Jn
Kb1u8rru+l9aK3vrYwC4kD2wJw1KAJ0iAUIALKtSl6lVuPRCs2WU3j7zjxQASyM11nWhKNl9LbCw
AbCvUqOfrWBk5dFzAHFcafj/V8ABIFtTqrHSp6ydEajDv3t/uW2BN7Nygn54m5akNNaYcnAv8FML
KiuX7uhdpKJ8SB8heNsr2Mq1NP+5G00S+wktS3mJ8IXTkTFZUeXpQLxofKjwDAjWqhOsIeEkXzpP
xVaG1R5GGBcqXiV4ZXat6ITScBRgjI4YaUi3SreOlGUdCMH3Hm/TQozsnhrgRWSC1XMW4IB2DcVG
iEHpX2ASPHsRbOaOJaKPK1EGnh8KeafzGka8ae5/ueL65svP0JVGlJZQip++MKHAyQ6+MV9oAwGN
5Zx3jBnyBBkWrAUrZ+DkGOZcLdQDueshU/BD2+SC+COD0QG81ZFNwGV4Bz1uvZDz7S8JpIi1ATXZ
EB30rJ3ldSjaaL5PKdIT1oNES2CQXbLIDo8Ck03eCNnAAYIAFS/eRbNkbqhqYHrOQ1SD8NfcQE0I
0+1NJQDmgl+lZWI5POSeeyVwf2KILuUjbutN8IZCCSaSUrjmYVQu87cjr3Cf35u/E0sJtX+Vdao5
h7r0VVA6wAwHkR7F9OD5mkSf79bp2jgvzp++ngOShZ4MX4wiakwfC5j+HcOrO1QDcaU1u4q2oLHk
AFSLbCJPbJsnlP9JOYiNcMTzxaR7F3zsNjWC0fNp69UmXSyjHp9PmPkGGAhjMsQdKfBVfOP3GUq8
A6JVouM4DUb6DLYTH5on7n0R3mRMwtajNBrmlLbr7FJc4uhCpR1bqAnzZThtZZ4CSCVIzleoww2d
nMwxlDlv2WFi0ocy3XkGG6d5s27CV6DYZfrKx8FWditPC8fsk3KbMlbb2ov+5FFcUVmONVlrnTje
T9gkepnIU3brrgKLt08xEdPswlMBeTwSNUnD09LbptXLC/fheSOC9Hva4Aug1T329sa3duEc8g6s
pWnMa5Ga7BBmbTTc1K6sdyrEvALD1grwD4hUc3fhPBzeRC6GXusazuHtPxbBa9qNMmi2gY6MgNbV
d/1ei5HpMpBMmQcVjZaD5KOHoIqvoB31DbJ/uNz3S2oklr2aOe1Uzc7EAQxTiAtzdtz+mMkteSJw
pib6xMi7n3bJbLZhbOH8I3t7kOIT+TRd6CYJVRu/P9Brg9yNDqLvtu8dtRgntKL110UQYzhh78k1
Fv/ixrp4ihCaPrL3WErPPloe068VeKy2XFW9frlROzEJV7C98JVFHZeSpmWBNEH7yf8sETTtuYI1
+iTpqzBVZsHnbfB7zF25vF8avBcyv2a25bmpbsjOEeUX49+J4fOqznMC4F3eMCByoohkufQktZVj
vE+C8iQYI+IYnZG/nhT2k8qAZuvPn0QXBD6tsUb0w15gMsS3l0FD5f3v4vT/lDcBUbpcPeQWIPu3
jecbk1eiwwJvn2KOulTV4fi1lwZCX8YhcktAKkecN3wUywM57WSHne0r4rqSavwH4irjXhXU9/A/
7/vyKvrpl4AZ5E2Evh3kJmytSVTVsQm9n2WHi7vHJD72x76b7kwLTvmyZzde6+LE9UKOsvIzSGL9
EVdweo0rEBItG64rSldAk72ikIoIC7DKCriW1JWCtiPtANkD8FDwAmosijILNcQppK3kiPhYBLAc
wOHfkT9ATyMwhuZteboUo4WTUj+Z6durhPAbXZsWIj647LV2y25SHyy9kL1NQv+BdnDXzCimSRzC
NPk+72rCoDRVkKasF1dEImoCXVCkmS2AzjaWngVZTR99G/9zG8M5d6TzZV67mvUoimRBVFuTOoIL
7mgqs1rpVkJWotHUz66jofMHuG9z8KhVCMwNHizUAfG/f3D8fmSCVEwhBGF92Rkj4/nkIsSYztSD
tCKO9LqMfYkD4Bj9rSUPEoCDjqkObxgA+FvYdZeHp5k0R0o0+EUzT05IFy6xuUs8zLEkjIRi7Yf6
euDU/eojP7a5m7aKVChlYTwuTP8bZ98aXJVE7jL/G3AW0a46+F5K4lukR8V11nuiLc/DQN2raR+V
ycsM+1uQ0lmrAVBNGJ5mAtOJNNzhFb8nfQtKryucb3XUbRcw0IOULVTPeRTHTD5/4Q/zCFeENtrR
Mg3d7tQjpBNwkzmPhosLKaggEimwW2DJSNHrXzKLnBGl/7Zo+Dm5mo6+M6nQX4kGi2vLwK6MeSBz
BKps/G8CT89aHGTMPabM/gzwpSdXwaHVPajARw+ii0BF3JCpJYshicfhafww865xwMWaWPKYSiuQ
OQnxx6omSLyj+te4Xk4JPg+rkt0P5pCIjp//6rUShdkQtduNeJyEYskCjD0wb0gRpX7sp0ItPReF
EXlqtkmdAqaHEEsj0AUJqXRsZbvJwxxJbtf3hith3AgzlnD0yW11uwbFsnpdaq1Md2gVOT1abF54
wfpAZmHojDDnfDCAMgcECpkD+/HpoDULCDoTQcsrhAn3kjg0UqLupd7Sy0VSgxUIj2NjBkpI17hf
2CKFXFioEDNND/bQn/ywsl5kxZWneFecNbRMlvWAjlD/zDsTB5wdBeySVRs223zf62VmqdoiD7oX
pIkaGxwuVSjemiMn1S5WU5NRJx4QEtdgOGMrn8ik7X7YNpHLWp9EqEjSppmBoLOdOz3m2+mSb5M9
hncE9yKLgXSBdpjCIyW+KWWTBztAE28Cey1sUlJlW/rVQ9q1xlUdPQOj944qBQ3TS33W4W2etZey
Pei0JoBvr1C9Tv5O1i+SsvRhfGlsjLfgyMD5kzuJMVxZntE1H6AjrDaPpdjFXv9XnA0CgUiqodls
sgkJruAAa9Ct2UshR1PGsnr9sLakmQmRvUWZASsIx3z8uZul0o7YyxKfXdI7umTbH7iBX9pQKrbP
S95VFOWlx77oQceb+DZei3QWZ7D4OQydWTwz6wkpoSsqmCHRluPPVUC6XhG5DE/dPTjnE4vG3COf
Rvn+xxXpSIaQJakW0k6+1mg6lUhuvK7uKkMPMXeQHZCB1BkWz2j8qTMpQ5D7pevxFOhFuecc7EBQ
id5SYTE5/DXhzXu09HKFTG46STHle8SwkNqYZXTU0AE3f6feIXnRd/iXCT8c3f3cbndvM/NHxMXF
beb8un5isQ1ai9oNNT9UYJZgG8WcB29+OAoYJ122Tvex8p66Gx8Rx6Wp+JGAF/nQjRoHysHwGzEv
ZyQJEl4d3qEqSkefcogBGyvHjVL2Ac3OT5B4wK602RJYJI2BM4/qJlWKlsGAPLLPS51RNOGis6X4
3veTCESjkOk/pRLgRk43NiyHoGOFgA53yYnaeQ7TC/uhprZNv1t0Ky4WhuUi0ipAMqfEmmpd0gMu
NSXDZ3r3mpI/3cGGH4OGGI5pSqiwCrvLNl05rWFKysHRHlWfr+OI0mGqmjzTeDWgGr7+51l9Zhls
cRCC+z6hF5fs9Hd6LaW8OWMtqtlsUb6QF4IrXA/k9als7H9CQOGBZP6zQJRZlHIWNJxTBxM+4ZM9
aMd9zxTLiH7UDOTVCHtip7837esDDzpVR8yMK62V4t95B+70Nmg+DEOlZCLWque+YFt4RIc9Z8Dt
HbCZ6HeD3HVlbg0m/jwInvrZILwugdczgDsH1cicQ1wQUEhnl7+sfexeHyZSKigoOTTtUOARxBdU
dvKsh8Vio8ODoA3WqYygo8u2qCmGPil8MXJ4qCyISg8/gIwITrBp4LAbdrhPo1Bv2qVzYQT5/U3h
QiQWSz+NCxY6vSPc1ozecYEgGo+Y/xVJWTA9V5qQJIsdnfXcWYgMDtdIlnF2aLi8mgfqHvP+JKMT
uWxH+pJgGWmpsNl6N4wx029eLEs1r1Oc6eT30k5+8CHjrU1gHGM8j/oFD2rg6/zYYkhODSwKhqri
ofG4xQBAAe6IcqN8cBsKWe3XClE4ziVVwEczcCE0komHctbfW/g23j1wxldcQad1Zl9VNHtv2HTk
gRAHOiRSwYSo0fWFAPvNqQdG/LEIKRrTR9wYiPBlcNiP2piH5YRS04AG4Pn1rGZjbAZqi8A2E81u
Zcx4vpYG6/xZPNaOck02IiA0nlgPoORnF8dX2HDi2brMJNFa+JFJJOh1M4dYjpQJdrFjNxiSODh4
n0nQheshB7kaqM3DJy1b5S5zYQWK6S1p9YTxyEsjyo3pnrLdIvG520BjFzH+gxIkLOum3oZbnVI7
3AZ/4CkEZJSbsF0t9bM6xgvMoPwqgk1OSp+xoN62POs1leLb7a/FZiE1KW93eSJWZkf8EbGlz6o0
DPmz75izGKB0U0+6uPXt8tBQ1Khr62cSgAb64ixb0ScC9gZ7oc8Z00zuz5w7gAGIpKt6ZmYx/cpK
thctjGg6Tmubjmgv+XTnK41lGFjX/HG2rUzyCZd5EBn+867z5cbtjj1EFrwz8+aES+OKpl0XIQbN
y6H3SvpAd+kXa6jEM+0I0LyEgDFF3cVKYf42EqdodD9BGhvj/EGwJIKXYAa7++pUJjqjUv7UB8p9
aQ2KpR9bP0BkEIjWqAVqpXXAGfheV6k3lnSoCedY2aYtCCjQmyKVbc7gawwMlzux97MdZm3VeVMK
66YbxiXPXqL9Tr3ykYMo4OvoMaqZXS1ksYE2Q0ebYvq8mve7tAFvngj8HBhOPl/H28VqFS5tFigW
LTZuoTFuO4HRW4NUI6udCrxAiYLGB2f0QRqN+EGmLqAyx8JvRPmgNDzVMg8CLmMPUZfKfXHUAMOp
tHCWE1orR2+fQGpnIFEh3wnjTZn9F4dId959nBHpenZNJJQ1LtiR9Cxvu+jg0XhtwjaHRd+VbTh5
uf2pjPrQliTUz4OAOABol9nuNTereYlZ42bXuYAEVSauYUXcbi+JgITj9gQ/lTo9nyRw86LJD0Oo
+qSiZ2Hp71WTxnP1qtee6qjbH+Ry/ECs4Rd0S+zLArAYpxjsZdOS8CTIdmYhvncseBV15HJ9+M7d
5zmeUkVYq8kwweKhwHHcdcGD+dqdIm0o9e8ZCIdRQrmEoF95J6jq/gRF+o149FDpKaAYBPSSb1YW
eHeD0iQVwUjUEbJPe4kCNsIWfkdd6ZP0Zy4IOVCLSjxDlsC/KE6jXKU7T95OiJgdKy4XMDOZdojP
3CIQxAz6RHawK6uYpt0CTwaoOw6tHcphfmx+gCSBQOg1AfTSBPzsrIpzXF8ZN0fOHwTJ1fABaM1N
fcHZ+OcqxGw2scBCzUPYnBaNHs1ugUC8AO64Q+jEdoeLBtY0YyRUQqoU1FxpoG6WJCGqkptPIs/K
BUMyIJN1qZc0imcrUjvOlPe1nGCWMGJoCi8Cr0HNoz+ZmZg2vHbk1UlpZr6oUDfvwuvYO8EkGsQ7
KuODdezeeTTQI14omYAqlhtuUAVmnxkZZy9xLzXUY4igl0L5FSiBmUZmrbHsPy6FVwY994Rb8i5A
f854OXtKTNxM7yC5LT7CaB6ugUYqTv30ArMCkx9maTb80Nn096cBuXpsXFlEFqvF49d0uKE+ZY/J
GRfgoroZCFs9kWXAvD7UYMJwEVTZ4yxFfNZ2/01akVZMwoM85pqh6uoTDhBPyDw6ZVNsKP+zArV7
tfuiDitOmiwMXWz+9GBO/Ds/lAU5AkbAIw/7NuGl/7WxWkQai9b9NJ0gIcTZ7ZGZqNE65gQam0Bn
vdL+fooAFakHrgwZSEvU59br6c1npjdCEg1cBsg57fA3r+KorSkIm0qRM7hbrO3qex2MWPhQszKJ
OCXPX0UAgQkxeTJJouYFGx0hDWzjlb1sa0zm0LahJ3AKpm4pL5Pxbu17OR/7Qbt3q6xJNcd9FUjD
POSV6Q4t576SoZu5uSr3jjzlMZ78bLeppMvXTj8f2SptPR0kahlYaIfXeZdfoL4dzoPjbkNOEuWA
AA4ZevodAYMPwWds1Rv6irkYe4rjMwRofh4J8ats7KejVSB8TMf4m6rrcFMM+BmiN/4TxylaRcPS
htaj/vgbg9UVlECysXGtW8PoYA+cofBOUcPpRFQvADrwz4ye/Ews6mTw0PM0ah1Brc/0mDqVnqMj
Q71J5SapDWZms8QAdl0xxUniPAYyNwhbEg7t6s+KWLc5cxpTVQrlb09xifGiF/4Iy7ttiaWcttyq
bd3/8fuRrFWdSdpLau1rC2N0fYD+PRPH/BlKQVKc/Oe41XiOY2smFRGlcH33Wq63oV00vxQydpS9
F7/ttt8FNrOBg0ZdcATm0JBI6TW58Y0sxEPRWFCQvl0b3mohcjunBYZwDfwWDJw5hzDELvIZh4wz
fkytOUTMmRtCtff37YYG8q85u+zjRMfwRVw9CZgKwkM2zf1IZyC/QwGHgeFXwXsbcsgpW332ld1N
OiX6CEVPIycG/eoLzyOGi582KLn2HQqPKi2zojYw0Ds+fjSyAMsPI5/yYcK1iTFS2bQFDFSoNWDO
b4efbYWPGY+dUUQD9G8Edy389jqwuFedXj2vFKvSy0CX3H+aYQU0v9/I9XsnZaWQyt1oc6CArkj6
R/jxEpkWvvEuSoc98PYZpr2hZ8znSBO3WHMdUIEeeQeVSA3DEPT4vQg9yy90KK6m1MHvulRl9k9B
aXAXU70elCbnHaRNWFfXcChp1zmNjqorFOdxOfoj4uz4uqucE0bujrIQOw792fKfn3Utt9JERezn
RG1lhLgMuJWF3gCnYhXQKE9wAi8WGr9fgEtoAhrN/imaFqUzFBRE3MnsyISf9P5or5caQdv66naX
mrK9sBXzU7DcKPAjs5g8J/jYyucgddckatf4PLdD/m/dztf8DtiVJYPrQYQrEB3sPINQztucaUBQ
8V/ZLt6noMlEdPz2uFetpMIjEfEJBXoG8QlAb1BBvagpCxJBqZ8h6GqlVNp586RvCh/w4/qLeVw9
Sr/PD81nVTLNRYtEDtLzZTURCdWAdknL+2LzK8KFxRkMGNxYNE79nOzqdb2YFP8ZNM98eBoG0tJv
Ju11PsX1DtpQwHXu1+PAWLdyty5MdzokQK9E9uwGVwNZlNBw1AjrMse0rAW1+KYA9faQ5x8VF3+L
ArL27tlumPUozR7evvTb0XFOs+03G1Bv6xMHcdOJapCxCPphV/6dRds1ZUybDyPRJNHWBPdIlG/u
C9km6aBX8bDTPOBfCEc2O/Asgf9e8buUsf/Fp9RWrMT8wa7r5vUCFy6fMbzGyW/wPKfWWm8Lkovn
Y3PmWjNOscxD2LDvg0V7GeaP6R7hXpzop1IqVMdi0PAitYtwZe7GoRwXUaXeiXrIHI4pgvPwMt/k
8a/441lCDICF2jewRsNJ1sAm3MgjFKUP67IYTsnoz3RERFJHK6eiVl64HJya8dETyCy/Jfo//zQg
CmajV4fWIwXiI009PdIij6kH2iM+m49wZuG1FNqyyoNr11SGylaPU4F3+vtayLhqB7cVdDG/XrD7
MqJZlxwyiJmxDfTUOEUdSFRYVf8N6GR/Ls3LO0Luh5u/7Ys22Bcv8uTinGQ9o2tYcvNaiVK/CuVQ
QQGPO1MsryVugS0uYmeABPuRQbfaHHgnZyjWYLZyzaj5qgSVmh07XNdtgRWpuC2ryr+ObMvzUqC/
pIp6cTxcRHSRI6RSwkCKIx4CySqOwUpOZP1OvYdR4nfYVySnX8BQvCngctPZyz/8xlIf/edPQIMp
pa+6xL4PpFy1HNAJyN9I6VkGdbhS5bUKSjNohyqD3tJ7pCP/pOBk7kNN6+LOPJq7T4APXaN8T3pI
9fsypeEf9MwR4Cs42YDfP4fp8CUjmxuaMxsbCPWuuidSB5o1AAmCdlBgVTZcgD0UHPYFtAx2mdSH
B5q1v17Mkp3JHJUjkHGg1iKMXsAWhptbHBtjxpQ6uAX78xTFnM4xojEboBcnpf3zpJbjwJtCSzo6
kiFle8XV7JcO7meSXdWeFRo9kyw0SW6TrJgwmFdeVzBWYdSrHp/jcY22ODslmb0VysoMQt6LUyW2
zYG8Jt/lmaawdz5m3NbB+IhrkiohZfzXyQerqZJUetbnVIQPCR5VSfthHZDD1r/bqeTSK3sG6HYJ
PObze5/7K6VUpTA4IVQIkUaJWHm0CyNQq8rbb65o1EuI2p95MOXlBdrrHCYTaqCIUsImk4Ybg4vH
LogqGpAfttpd29PdxNgHCjtOMYAxSPOi7opk+cQyaNK1h0KkwpLr70HK/ngdAbuwEg+pMsJaBT+Y
H0neoNYpPp1Oqr/sTyIhOF2O2G+DqzHBzsgIFcvkLlKmcFWUjiS/glFC7HMTUZGuqQTQHAT7r+FD
dHDVDbLMOVRpUhKsMcBnCm1KbMTAnQvcC1N4VJVA+sUz7HVgPbrAi4WNquIXYXTrrYESogtfyoe+
wSBO6rxR/oGug72KOHC5qG+t1/D6dhz9yJ3ZeQGPbbjAQTsFKj5CbFR1nWGN2JjzkNhGmIZkT2V3
YFLyKvfPhdQ1Wkuoghtw0GtqfeQOKV853dloFRZ7Jm0naYOqtpqcLHFLsiL5NVO8C0Ih+fKDpogx
iQ/74pr3K+U8GcCZuFAMzVCs+AOVds2pd77EHaUscqOb30abKwniDmxej1c2MB2BGMUSBxZjpiuB
xj9Fgjo7dwBPxxa0qxsepT+IAx1zOukV/DdbgaGRA5QyYW9nGF8Om3vv6iEWqLatdGXoKxfe9GIL
Pkqjm1b8vGg1yManNFj7/rmn+0mGVI6woTgUyMZGRuSlvBtu8E3NT8CNO3BdNqjcTxx9PJNpYXPH
/yN6RViBy+Vi/anHsKvwXbX54UYnG1SAj3AiwWkDfY8KuOvMwgBLYn3Apl7GQvsoPLxWOJIXFC7j
goMRKIU+cL/sV5mXY8l926g6AF427BgyLvk9zbXCXy4ap81myuJ4GUgags0mhXlVcUIoeKMjU9cK
E8RpRsHRwzmN0k9bzWXuyDXmpkZuXTl6rBjzn7XrasnKQOaLc+I4n/fxtVpZuD5xe0vmzxDd6v36
4mDUdRn2DjgidsBuoyE7CsKlJs54YFBQgv0zbI9QyCYxUSvHbA+LtP/81fBdsoeksgGkRCnxUcSf
for4WkAe/OCw8UMowg2XDB4CWrQiCDjW4VS6Ql+QSrArSMxzx7XCe7BEdjk8pm+klwC/2Tb6CJrp
rVrDPb4rqXlHcX0+EqqflCdIu4pUNxGrLx/gpaUZogyx7wCXl0zVKkF5U8J2R19bK0zVkrcBBDDd
i7TJQBCmxahWoO+7pWG80u2xp2AhFsKkM8HihyGlO+olDJhSao0T4Ri7NitF653Uq2VwcIoxVvqp
3FToYiEoiZAb7UTkXwIH9Hi6dBhTTehkvLmb/82EARJhkxcZDla8tMJLpyb0L11/3Aj18V9+Avbz
cwZPZa5eWbBHHckY8Iy3ebUdd1Bp3u3Zv1zW07StXYjWB9BsVrudfxzbK38TO91xPZBIFJcWlGaH
TqNMOrc5iAXF9s2MdmB5xyMRVx3vc0pxz3obvPdEvrXMcKfyW8CxdlrTUvEYqJWymW7rn3BCL4ch
UlGXIcHgMwb8/4oXeiTs4fD0XQz+ivei0Chxa1iCED8GZRnrmEzTwA/wlO3PRtKxH9fmrXx1wPnS
xY/cbwbco4NayabAwlnFdjyONRPXg2ED64tVSWuA5hx1ccm0k8qU410VG+20Ce6QOZC5Ucnniy9N
8/LUCmRbJI6CqvCOjrkfvLU7vmyomcl4uu2X2Y8FmyzgQKKWn9jQjkBjW3buLypSWO9SNWCRhJ/r
7KMtJmn5YMDPsYKaRLbuuek3SJfj+i7FeaACiQEuzdP28eZAX56U++sWzd5OaL+sbum60LqST9rI
vmxtCbPs8kMwv8KXACx2Hc1Qlhl9CKWsKghkkYsRChct8jIkCLdiW/pNb0ID+gwgbO3O/AioyQcw
7Xpjw7dlrD9r1qaorcGgDfq6N1zCq587yYKYoyvyivJXAn53kpI0UlBOFDl/Ok15XXxutzVWRH1N
CjXB+A0NtmV8AAGBE4ZzYOQpakgAs3yN04jIZMwcIzfHZ6OgwP6TaZ08L/WxVS94Gu+Y09axKI1a
4OScLvl3ATwBf4Cme+p4tsUZ60l+LEpksqiSmTU9f97tiDkkO+RmkoELa4nLHOW6kF1c0PQ5uzkK
MC5Q4fZDGqw+nvWpK/aKlFRU2cdO9mEIWRjCylbNPokoyo2oxA9FfkMhQFpGfO1euou0ZyQcEyd5
YfpTiUyeqExbo3/GCxeYpJotWDAym753cvtuJOhWt56wEpn08xhP3Q+ErcgGhDmuI8WLCBds1XVd
UGEl5SP0Jk6mfLTxT0YWyp2Ic5YE7wqVB7mnBV1fjKsCoN6T+nWJMDuAbj/jGdzLQidbSTHo4pW9
POTnujZrzsFmNQBOjijTctit/NF8LkD5C/C4k/pMWJPlOxHCz1mf0Ndq2liQEzy1vJqxV+E1Na+J
CsPKB/XKkcFTMa+sXjtjMpz2zVBSoZGq7s07Q9Zeas4tVhTUx985Wvfwh8PSyFYbaRdmSLtHibeV
ticAVy7XlK0UUU6Rso0+P7pKP5e900Q3UVzcZZdYkBjvUAfSF9H6MKzsxfcLZ0BktMxoUTkc1Uo9
jiDmTl/ggsmmBg88PlNaXGLtMinDcl96kRRBBkhC1LGmGHgh9Jz2TJpKvQXGJHBIn6Z19CnbfWev
FiOWNnqs/+jLiBfEs0l0s40jiyvFlrnvFnylg0wvmpGDFn6oW3CnUss0HfohG46yoNk5ByYTOe7n
oxueRXmm4TIaPrOMKZhOKSu1GxS/yfiVIOQu9dd5YT2HJBjGl5WZorOKDIJ5UmyZ27Sxhjcn0G13
OCd+O1ivrlwexfHk5ehFeKZCx7XzIj3D3xuI/T9HIm8cJGCsfrABCXsAaCYZRLKtyi1dWcLOUrE/
yteK6RCyPlKLwFWk0PsiEA0bxKijvfsxOnEsCget8mjRkYHVfYc0BRiUhv9w35hlAksD/0Vf6wml
dgjAlIHPNNMTbSYzcF//nisha3iPx2a/7X48P1jfWT0uIjuC1ZZzb8EVHZkaZB+Oe5YnYGc8vwUD
+aVi3uJdkdvYGMQ7L7Dj6Jg0ZBd1kOP4TaAtVid5knNvZZWQKX24OJVv2CRlaaW7kUidJPJqRxN8
1TPT/1AKyYvJt1vpLy6V9a5CxTR2KKqaBu3dCWz6WWmSNfgdBZJGXzVv+iTPNKbieMYZQyuoIslk
ISN7YJAeZ4J8qXJf+w9bX/Twff4/DCVG49k08CXGlWyprP2weMSl6ESB2M/RO/GrppDnnwkToBIm
BkfdJ9Vy0IgTylN4iDpuRRLBw34ZoQkDep4hbsIm5KZBbQCMb4rFtGEi05ss+qTxQDkMc/POLT5l
B3sYhGkG4VMWHurNKPt1uMbYzr0PnKhOo6T/cJxOcOYKthw07ENCY+lE0ThCYKuuD5GwZDQ2VtYB
ghndrnMVMdOSQVc2SAMJ63tLXnhWcdbFdK9zYZ4TWQOnxEN1jLSHE14ZEWzv+1FeFBwObXIpPWZw
d/Bc3OZp2EplrToy+RwfBn0QrzVvdDkAx/yqBYDgNGmHjiEfVjv1vjSogubLdtCigwtL2zQaruoT
yV+azFLLFdmmjMypk62OcEcBAP7LA0TGlUCG1Bczs0aKftG0dnxKrl+PkSgXCGouAKvpkXXdqfrK
E5HmbtUlN/33IhdTRc3x/S+xKiqdeDaMfvh353RMnTxHYz4/5wDX7HWsBdIQLQf16p//Z2nQPxA0
RR0Yx9q8+Y58heTgPt8A2zJQdlZk2zuIzs4tJMZ2/6Y5QenLCqWqeNzB5MhZ0OtJCwv+Gh0eMNe5
qvt7Z1Ivht2RulMwT+hfL52JGLUcqswyG05CJF8qT94bf9CQZDsimWCLPix5SyHtzXj4wG3JKYgg
+Gd92PIsPCJPK0mKXwFrfZhZRJxPCk9cQHtq7dGwVDYnrzxmDWfu4GgNfTg39WiLXR2e0csXedbQ
cDjJLke1XQ454KWU15+jzKp8KXwFmBdzPAbX4A7DHSjQTiPKBZQ61QnrWOdk0mTAbdHPkLpRhIzb
aKYS7bIH25s9F27rgMriuJfmiTzcTT+LSbGxP8RRMEcFqr1oxdY9FMWIE+gIoRM2Bb+pSeKxR6LJ
uK0vUP/V1O/MVw5B9odaGIsB3Iwnc9JJt58pLosrjm+hJ2ScxJ7tiI8QHZw8scAwt7LxkaG3/1w/
5zUVdbmtn68guTrcSbhAuiA5+UySO5t9UX9QXy7bEp6A5wTqrIoxFINnBY/0J6j44JZBDWk14ulm
zY7RZHKJ8Weo/KsOpXIKwww26tRk71TJh/FjUQ7Ye2wo6AoQTdSMEWVQkAMCe8mvDKX99cbuDqv9
wqf6CDOhsTsiVBKpvoQvxyYf8PDQRy9Ib+zPnvDRb56RlgSxlJcjWCNu6h4ddQiz7vai6zYMDJNj
IB0/iO/rbmol5Ar/hv5PB6hccWyMMI7LLwvuACF0T0KvDXcEGPRfi0r7lmsOBdzcvKKt2/dKe8Sg
ejbbc1RbkND4gGunWccy0i7g4KuWzmgTuoLBrSqhKeVUI7OTnjjVbBnIkgyRHZMXTpkWV8Xc4n31
1xzRnU7rRZQptQ55qBE4g+pF2qHeqa4OFOzVY132Q4x2do2Adq4mw0cJusrbvoS9ClHWwAqkVOa8
eZ4+bPoOB1wHiNmHd9saIZWZlftSmdr06pAFhP2fx6LOX3HYtxFabAStw+WdWQvf+DbR8aySqLcR
rJrPjq23l8aI3LXLAKVV9XUijxt65B81d61Q7Gjomx4T7xZ0X312Mvxcdq45rzIQuCKjYTn6kgju
cxxmx5M0f8tqeZ3zOvi0vywjp3H8gg7IXtIUIPLmtBqCAhd2ScdjbJXfy3D0JNMy9xprcQLljaQ5
LigY5KjVw2t8qahCP09tu/LkOuDXJhKBjtjzn7uDQ/0POu+49MI5jOI41Fg+B6jZJLhzM/URFw63
x4CXBqXUlr6m9mrLTkifV/HjlUVen5xzTZnoNzWcKxMyxFkTeBXgcffOwJ6Z0pBOPHtBbGwVfjfw
3E3DslyYDkDd0tZE+cDhUNPfO0U+uO1wGVDUWlTPCEyXmt52vk7HAItjZ2tNW+Zc+LqgSSO4nwOU
+Gnx0L3QZPEONkH81fUHszQKxROUf4JgUTrTD6pqWnPOHgu/SipdG9uYROauCFAUNXPrQtzSh8Vt
weeOgkQBHFiM3o+rNaBvv7e+phTQ+yl5SfiHTSGtwUg5YZOkklx6ShTNH5GDsvAtP7sY8iK5EmHQ
KG/CqJtUxZu9iJ9A66mEUPxLT+kOqVU2MkcIfDQQx+ubxKPwElqKSk6qvf3U/7/s4hj4KRmMgm/m
vCA+ZcOhQ/8ltw6yWrUUM0Myh4bg0htw5bG81KH63vcaktFHOw1B2THUAKxcuFJhA2Kh5cbb5l22
pkBr3r87EyP/u+yxji+wQ9XUjIvon6f5vqmyEocUfAxx9VDyZwow/GYMy7Q1KSTdw34sy2tmvlDD
E3D1Ve1QQGD2ioQSN3w6GvsgswLV3yPn99S4sw2oNxpSRcQNsiXD6gBpekQgpjAFWvGxuMyMDW47
qhsewXQpcgN2Qo5rCu3m+YhdDroBwJiAMKRnGrDu8F+KCrzpcJGv7wscHNKM6shrHQwRRmKO97aV
tcNhBA+1zbJiZu5n7l/Vh8UC6FByh4oHQWAUXUCOFicddw065dirbf7OOZ4Y3mddGX2NEKQH527o
7Rc1dVbsHiglcqsTA/h35a7NurLl+KGnCFnb8ly4MaWMyjCdZmzSxEu0OlZRTnXdB1RuIPVevpA0
yDacGPJ/PUUsPykhDkwOi4AcH1Pf6TwbC2KipLPKh/YiAXLMuQQaUdtfxHus9kwfoi+PUraB9YYo
sqb+z1riWcQWThK4rXO21uD/1p8smnmHbJE87wMp3d43I3LucOWYTXlHHgCKKYBs1Lqp3/7DIFQT
hnQFR48edQ53/+55vyjAd2ost46F3sIaEb7CXybtWBu4JqeV6wAGT5aJfj9GOSQVcoqHF+H0vjnY
XjH4I6+VRvxAXqEm4K2V4DpAvmUIxfBZqYGp2GJJ1qcSAzoXLG2MRXycv0cQndygnGijA+bKSBt7
qlMdDFpQrmikxEOAcT5KnRboGGaJnYnRmjtIJwTsUXg3G8tMypoFKBlcGAyImr7EqGNvwhwSdnGV
Xd0xvqrobat6fxKgP08dWh8kaIPpiQpkcSkFOMtphtecYXXt7p3ZnRrGZiX43VsrU20tmd1kp7OA
hLpEC9WNKAED7s0UjntWAT+iqtA+rlln/ZZcgVnXCeZ9lG5LyJNxrSziEShrwz4XozD7f8PzJrW6
r+eaQq7dxHFCcBh7dgakJ/bqcvUXEVgauozfZnmwn9Hf5lVCzD3UbtGqB3BxFTrL+W7vQvxD88DA
YfVvM8eChmbfd1HV1zrqw8bPtorop/+0aXRz9x7IVKlfeC5SSLYmeTLLRUGfIpyscvIaaXPJSgft
MZfRg1E+kFrsm7c1/GxAf0zfRIViWIsm548vBFbeaeQQi0HFXp6yn1TYZStg4WZsMEhF89sBWP32
qo4ZK4hdY2itAdNaotuQMOyvwN2GwuQB4apIQltsDWNU33ytz6ABoivupZkJcjM1wjQyFr+L4eE5
vvxbdTwIEd8I7i4x8YYkP9Id8m3Xa5HxVXY4KIq2XPVfn4+k66+LfDtXcIVUD+AlsQ+ote09PQuk
D4Ekx7rakaPc1D340klzLyMjjRcldxr1eJGwCy+D/Yc0rL3aWqbzhm/iPR6XXmXMQM335zwYy32X
g85Uh0iBlr05F53ehB83efroXZXGMUQ6D2y05iWZ9wt2AxuYviYVWvRqsub37M7nO4vW2KHQjO20
j1Vi94OkjUpUblFG3kzbXYFTw/i9iI6hRl9MwrW+rVXQC15vfIisibgwDWHEcvf8gHyJ1RhyeYkh
E4QHnQWPh8rhA3pCnhZQMOXmJmDhPiHswJgfbtUDixA+d97K72MF3ip5Kpo+ypYUBDzG8I2o1vvM
TRl+mUNNOvaqwV68a6Ymz8hRB0hIrKzT89Aoh2RAqK6qmtbEOs6OhruVXt6dcvCMXcLNE5XXASvm
P4TY2v/l/DIj1SvHiq4/hEIHDYPKwwZcrQhV3YXbOz3XE54RgHy8n2ygY14SYU8XbQS3qUc215gs
2ydt2d5vXjboI3fTaeJrz0lvWyDSX6sg/iu1mxq4Sn2Bl3DFOOYk26/uJzd5QbiDVBNlSw+yORzd
Nx4L2yR02HfULRQKM/2WZ/VrQzV2E1w9hmeVfJa+vAr4UCLjU3z2jG5wwPnMR4PeCA+raTlKAkDU
DAnPYnf2FowM1YpK3ePIWL45WyhaFvByOS46LGMEr2iqc0QFfvLsEVGJ+9SiHH3YSQs0oUWKnlmf
W3AUJtYA2Wh57/b2WEinaKHBfqMivWA+aVyIaqTw98l7a0sA28B/5pICbftkABvr7qdZvEvHvKjT
YQYoXaSxz+7r+eiQb/102JFxMvQqalYOc9+MrH2M/4ToxnuARg735Arjr53RkZwWVpy2Cec4scS9
w3DEux3F+R+SPEHqokn8hETary8r29ATf0d36JJbM07s9vx0noGEtPSBOPmqMAJxFFg0cXMzY7hr
6dh0n7XPM9Hy2C9tBMRmfOniWwW7OsFWA6prIdbG2on0KXWTUcAg1hLV4QKpKaaX7f/zdBWTAepl
0hcKxPpuwiOhUuEhL+yuPweuk+fgiYD6g6dnM9YHIf5/VWB0fdcLJ9VvgeTJ+qHX6ly6e7mbS3tT
JgIEihSOaUPEre+cGoPEv/OYClK7cpay60lgdtFg+BCnTjAMgUWGWmNL22JIliNcXKAEUkZ+Q04r
gJ91JBx/2O+r5mPyRDOn9vytOTOVXNJiTy4ffgrbjgKzp3sTVSfvuZT9KJqjwkdG7UngMZtaaNu7
r+yvsTlEOR9ZeIvMqvmxQQGEGbpMB7fwGfBQrv42IUEcJ9e9dRJ/q6H9FpMAXelGUlAHRUYS/3es
q6z06YUadptCp9J/3ogxZogv496AjQd8TauM4FifVdU4eTT26KRS41ikUQseAwgSJgxTMWCzGNKL
xMS5i149cC+gjTXa9ONtpY2+XHf2Ci7qHNngIRQS1GP6f+kjH/nJwF+1i3bnKVbgYxRZlgCj1au1
TENkXFr8qCxgW1Kfdws6co7dIj9fbnVLPKFtKjBRHf/ZV1lVku4g+LPSU9TGHN4KkE8pRY8gIuu1
JyAUuX74m4HdafKoS1WkvovAw/Bq+3XVgfgFlZ/oxoMCqeIwUY6jkSz5Y8rZXRZpIBvrD+Rp+87y
AVOaFJ+F7Z4nhqUx71iP+zOWYiSfQwMb/y75A2u+fvaINpgnVvLsd5cb5Y30I92AOPYbX2zpSRXS
3xm5iThKHXE7dzkz1tTzYIr7lem4KzCqiURKSPt5kqpsp0Z6owZ64ID849cjtKaAStouqyHaYyq0
MTSpJkE3w8qIW7BuZvqJQvaHhYCaWnXCnJLPeywcnRXsWO3OHaZ4YWGe6Tu5+5gWMXvTigsKu9Bl
m6ft65qfQC0QwyJ4r8N2Zyl8TU6KElKG9TMY3U2wUhYYQMhF8TMhDFUuIfzXMFOP++aA2g9IqFsp
0di4ttDB9gm8Aqx7JlwXojX6anUNHiXarDjWMgDmcZ/305ZHDz3UUo1KVdy0KgXzw8zEXjwN7VEn
+iyf6qdx4kU6Kqf+0CaOIZMJ+TrmMNXx1M0O6H7PVwU2yWQAbrNWFQPg5q991e9aS/Z1aJNvM0Qb
YcUCJX4YU/Z6un056YGoH6mzNdQmBYsVC7DLHvIqoa92I7NF8QS1mD6XpO8Y7aHi1O/mneUq2N3A
kqo+2d36abH6EWpDX1x17ZKgDWzebK5LadziYEiPAAXZV/rZeAH9h/BBYIMFw5J64VVO3s8cwabc
9/X78QJXe/efLO8tGEDh4T5oZilxJyPHhFC1cggMBZBoCGzCfhDKrdGRWRaKTGUhaAVttf3l4swV
E7qezpwntn8MCJt2kmgvZdDnBR/uwFkZQ94Dp21upaZ6Lv5MMbUbF9j9YOqbbv/OLNip3aJT4fo0
S1fY7EX0JJN+ztvxIS/lMO8hnlZlQd7ET7Q83KZd3bhhOiOuuDxPA0k02Efbd7iXjQndH94uMWl/
iJRG6bsHeaqy0Yw7pMYhSgTA9CjsjhMONgfabDkJZ27beYvqaik57bUwVMLMMIBdfpsDb6x+vhw5
CjLrIaaoxr4cqqrSLTfB0QJ8HuOs8G9DtA2WCgu7kEdPtcRYryRVOcmt8WSEcvXyBi+/vy52QWbr
/dEcAauhUxjUIkY1qems9sRrv/weaAciG5bi/HK8vfvgbn7Hv3zNe2kVaPVuDVcbpvJ2BGslalCf
gsCpLoZ2LMILDimSM9dWrlVW0zSxg9cJoAQa+nkoctflAAwR2TOHpz1KLhB5MDFkF74El8/AvLDi
eGPFp8w6fzCbbQJnjhGiS1+h+vZnT8CYqcM5uf848UKjcTBdr8MGxvi86xl1QEko/l5nMQ0qbF8E
N1OcrzjjXaXaBpHzrrIvMXYTZ+B8rSxBMgpDWl/lJLTFlk17dv/pP6HYDbDu9FYaFpamhxMZb9Vi
dbOqO1csQI4hKWmcYWuMKylR2p7CmkR+eZfV76InbWxMwRZeZ9xxRaI7HHQj2Y2hDR2ixx+16EGb
3XoPdrK1Zvcmo/hCnJdPfli9TaSGEHxkZBAAUiQxa3pkyTQ2d1x0UHvCcxzZn8dhv9KZPlYpahdr
0La2euEUdY7snCbseMuhP+l9mPdGq/FqGeoH7eysKw3SE7QxMdvv5C0WQPKqtx59PfdPn0XN4uRV
02bgbdYmBYjeQkLxQlm6ZdXvaTIdYExtCCgcsM/irRg34YphGsGMNk7+ISQlmPsJ+HXAQNi+FTaD
w3Wop5ON7UTREG+6ypYxv+LSzHfUuEm+192VuXQjtFZVPpxlR6uhssTKVOzcPDTxMVebQ/8hzsNL
4ixUL4Z7FBZ/7iafGgHGl3x+m6gWJ9/CQ2w73ON5i2mIugNFJ+VM4EIEv3ML1O+pOUvYz3YuqeR3
7VXy7oylhcTAIqvTdG789Rjv1sFydbpdSQpiwarheDBX7nkA6uJ7TTU4ld27xoCM4NMwcaQ+ndum
7eT4Jd95ugYVcZD7SbpSROBJGtDP9y4xE8ln9puOo7p0PbKojIlnpf1hzU6/XqxYR6xKSHEdKtj1
rEjWwBdtxNJf19VeDcZtC2hnKuxvg+OwBFfrbxWkIAZPsmsiICRYGpuxqhCALAwrudeMwhIWVVaN
K5sjW7U7WfWLdqHSPe99GFLKqwwvD5dGBnOy/dLi0T+vn85gKRSJhatgn24juNebgL5ifVjfKZtP
ddNYTfFpAZGS1bWOco9AteyP2sBEei7a2cvnHO7pmN4C9Pb50rWkVHczspfIvYshjnwVQVhcnErI
5VXWBZdz2ctwPcSdIbSPMHsNnToV7NyUCXO+W/RJ1Oe5cPiNSvW1680+kDmpCA7aUtUW4gZJvXjO
ntHaeMwHnC06h/fvT2XGtroayZ00M6/W0l977ARatO0RRRifopaCQhxnTdUkbumJJDBLkk013W9d
8Io0t0b+dxofL+/rM0+Qo3EGsVcy9KVcBzIKJlNfJSITlFOeFHOHP+ff4m23P50iJZOG1O0Sylei
9w7yybdjlYs44F60acXKtUY4E6RBt3549Tv+D3nhZFOG+TzjPtSSXOek21gq4RyMtoTJvOiHXBbZ
Uv+dFT1NyK3M5GROjG3bCOZlIS96ltnJbdRPUonK6gmk2NvvzqrMPARBJFSKCeYSMMv3StvS2Ylz
Lzo5ZPGl9b9/z0Kqc6mK1HK0TEEBpmnlxmbAz0lyZK0cgim/Fj/ni+Kej98ZGquVkhBM7QuImHdB
VzSkcDD8izwEXR6DA2EPJH+jFocUJ9PX82xln7fyN0iUMYe8TbzBCcrdJfrN1E64XF5JETlObkII
mPiwR8VYYMR5gHnonUdVky7sKN2F2EAk4y7VIH84tXrIBxvaasApZU+DHHXHdxVzgAryRusmjsFQ
0bsuG3xFojgHU1fOTl0owYhofRE9T7Xp31nxdKkNzWWLm3GrMQm8jyN7rjLgyXxn3Lu7YGOTsA98
YNNQwK5PpMqTgMY+2+121zbl+7Ga4Rj0FLxt+Txg9ARXoLu4yTq2dn3ctZkuhp0/aJBV5EuxvH9w
qdbyEE9dJ2ZzrgglKtWiuhhokjah5skU3JaYeP3PNY37AW1rc92ZqqgEe+8Yy4tR3MWItGECSwej
w7/NEmCG69JJKmzxDp7l/PgyU6exsZ/visWHtyRG5Coh/+G2grRXleqSAYixpyNaaezSmOL1M7VI
uCNRDv643d/0HyuLB+0mJp/ByyQighpS1B+YXRCGUlDQnY5wBHpsIb0vw1fqcBqTOWmqwtBFTNAP
RScrkjr5SuLrxp+RBiMJGV42aazImm3LqSNAhaMYDKau62aVX1pl9vwU3UcM03/0FaUD3jjp9Ghc
1suhMH0OXyuNVkryEEHjtcX/4SpPgn3b4L9QwhPWO5Er94pjmQswcUxwzvL8rWrFDyC8ypb+wJY4
4Mr9k/5IvPx6RzfLL+rtJYOitrkCUGx9aWwFMLh4Fke+7APwQXXL8FSEBNYPLhqQWi9EWaE3fZIo
5kNey2yD92IjWzVbrnB61aee04JDtobL9/xHJtHOKdZNt/oDoH4Rt06MFyUz4aDqdTbZiW21ccO7
7V0rhULGuJdWNfI4+zYxEckAjNuTU+79kDjbv5i69jMAEJj6Pn2l6YlncizneVFbbmDDsSR/L41S
Cl3dXHJUV/TkTZjQ5/auGdinnjV1erbtTLW9KOVdJ/xWaAHqrsj3mP8bv9NSUCIfG/dNF3dmXGFr
CuTXrrzKMZcxmmDjZSZDQL2EREpxVZHyVOKERVESNJ02D5/ejilInw0/VyaRdal6bpPtoK6Lqf0t
8Vs/BkQ9Lu2u9CiBWI0O6UXZfb7cBwBH8xHdYxeDrwL9zGG+iVTXWU/8G8nd+43ggPXZbYUdvawa
Se6gCVNKLSYAdOPjlklevRRJjMe4sWE1RZM7pPIesKnTrV8F/vzv8fWWXpIx81cQpeC1JY0pwbXO
X3iJCKvYipwqrXeE6/pB0l5OlRYnSLAl0Ka88hmLzNC0ehxfHWBjz3l2DqL3PmTrTzt3Imlpo+2y
ODihniOnN7s4UBMmGNYBNvrjg+FbApERY4dOjyw4dOYS2MwSd6ge4bcLjY2+FeE40SVeqCCT/4yO
u8P2YuobV0973dRtf61T9JWYmVc4TSdwwCUkru5n8teM//iMW+gIO8rXxBdzerL5xE9773AxCNAg
D89Lf1HzlLlF1FBeWVjffyK4MK7nugzs7HrgVqTsLCPNvWT/lSua2pVr4EU7fPBwmXiqEFC00sUe
hdNBMeUIN0xNfUwdtpSvCpIrHPSMfhfjD1FVhZkyKr53QZgqidznAn7AzH99weSMGZB7PIPjJSj4
lacV/nRcO3LbRSjSVwf7Sm5eW2p3GcQJ08jM4Aza3+Tpekqdb6z+rud/ieIygF665hQ/WK6v02ty
LRM+OdpLR7oANXVjYkycE25IyNJdIpO93k8wxMQHCzx2z94JneZ8bZePNt6ZiM7Es8YQHerGuzFv
76Gbt91bgiGHilyaqyfPAtfAZjZLM3yGUKQ3xGXkWTWMD9IxwdUQ5kxXkZwSd6OC04uGkoEg2lyD
EWShzHkgl0uF3BWcPoBkq8TQlCeyjOXUIOU8o0O8r7CZFgCxqQ86zwnRfplmE4bmH32UHjZZYHS1
Pj9lD0oeOqBKuCol2kY77PG9guFqGxCaIqSCh5Myc38LVHLPbrj7qoPDrEJUd7+cPRDlAhcAv7QF
/CLq2kqzbqZt4aCwAHqouK1WroRiEjxQR288KqCu5Bkt7C1qq4CdfC8ZkaMhOlXwuC+/MGAGfIf3
s5RYFZNZUyFkisWsWmUN2DqAaFw/JobsJvmQSgiTVB+kxJPAhRkoI4y2Y3Jy/qGQ56tNrfX2dBo5
cVzByD9C/ss2X+wJHBkpumkhKI1gObiDRa6zQ20aaSrINnpplfFgHGQo2kWudBxAYXCx76bDvsfj
jryzoe2ZFOs9FuR7rXnEPaUNKumMv28uoAaEoz9cwbg5lykDE0PLb14fBXqbP5tySIxHofy9Oz7Y
eAAZjKDjwwfwdwa5l3IaTqqQmms8Lu3y2/H5AVG4aAMsLF+00WUG7hZEoPfnPm09OjgpYWCPgceT
Jb4A3+PbqQvukKdAa1XxYlSoHIl3dH01Y282bMft5EamJbHR0YcovPntCLzE7s2MMyxbeIFMaSva
TXAny2lzJeLs+nRKg4wJ+UmCfYNkQD/U2NFXhG7fOy8v3upKeSFFrYuTYZral++qK4F6E5WTlrwM
LjR67jy+7qdNyB986qRDGi6kp/W1Hy0PYXjZJyWW3vXzSJRPnvzgjpmCDaLdxaN2C9+rBI98w+fw
0YUdvJk950uc166mIGI8S2IO0K6RZrTYPI7PJjP7J5S5V1QWCjOhl8Btx1mUOjQmh1e3CNVontHC
oTXS1+oSgSK4bDtuxcPaQLhL1+TGCwvcD4mEHIkP7OIVKf8BHyGkb6SHMfg91QU16iJMsNOzNU4n
KdBFnTSd0LIzfTweuUr4GG0n6wMUQAxRQxCeU7cWFQOO5pH13BbP+zB4eIokDRqrVXJfc0LLWsp9
BNlCV8wZhwHdd3h9Z+rr6OazSrvGP6O9lAW8MqeMjDeVrudSqJR0mAHsNRSTnQNDWMQpxJp6gggN
oc/67PdqWho2GQyuNJG/L980qTIlcMtIC+nrohc1L1Fl+RVSKvjl+PaKxc/QtjPcVH+RgxTg6a27
8/dD/3O6GZfhv+ubb88YDZKJgB04Up8yk00Z2lwlstQjjLd0UaGTqsffmCEDkEFvMHHHfvjLpcEl
bAxdyksiiqOFYq5QHVgoFdgQhjmuqcK/MgEGHG96RD91bbIYhvoYddpGYkrMeWmk4PIt2PEJEUl5
4r0H/rpAJtkVTKEalef3QYfyLNdgOc1eL22OhdNHii1fmO7W3tuo0OywHA0c2Q+s9s1iltqr+pfZ
yu/Lc2qZz2yFBL1lJK9rNCpe8vK6SzEI9RmVbDpY/zdbfYI3ajK1qPf00iCASq0P899YKA6nkQDk
pbuO63epZvea7WOcyng3O+u2QXeDTcKmRIRw4ATjws8dCZO1uWUbbTgCsrEVGgGkeTDy7uWhePeM
eKJMmLmOYi2HsZ1JZ0+++2UFG6+5jot3oMUEpQ26IkYHxlWytL2RpPHOo7hrcb3jFyPiIWeEPagx
vyj0d2XKA5UPUPvw/SenTvdmWJ69Pvy9zYuoiA65z7hC7H0W0oCyRW3ePN0i/BPoz04egF21W6Mm
p6VWjQtruXssnwnQdloczQod2S8J4ac8mD20PG3YXLK8IEl3yybkow1rZB9uhvTyyadxK0Rldjpn
oBzrTC1njjPy1t/EORHPyo/4IfDamsnRWa6V5lXCYPLbbes2aOnRZPUWvY5E+iUDR4PFf7jqIwKF
4EcI+2mzpN/WCaaKJyD59aDYaadesoXOuEmk/9dwHVIw7rcAUtLdfrRjXJCxoCZCEbYad85TvbuS
it3Pt24LK4QXCe3/A1BM3/LBlE5BhGCeKaMwF97AX+AmXpE6TFvj6P6t0w7hPiDYBYBbh+dglGSC
kVwPh8DGittexvxD0hpmoXD9SsDrwwHF6c5I9G8eEUIAITVv8F9vSdbMajSTssh3JvEdPF9LJBP2
k6ffn1KNA84lcO3zZMAz26RkH+zavBhYcdn8UpRFkF6T6L0J4wad4qll/IUSzoiYJ6zlAUObOf75
IRnaeJXQudMI+CNZuhaIesTzBExx2NF8S+WuaswbZTsesjAtjMStRcGkSjpAdhMRL9HFpVCwEGi2
al4jaYKnTF6tvXrRQ0alT/mWSMG7UyEsCVGeKSfcTRuwp2eac4++dIe4iV0nufe2ADWWiqbvZcLa
xCjOlx7nLU5NHKVFNvP0jQrdiaBP0WV0wDY4HNHwf2hNVtfO4fyY252cRu6IYTIOVhgYtJ2egh4n
RxnnLZ1IK3CFB4B/QPMAY/QHzVuKIRrhT/+kZjFIcmXHRl0AKAxNV0lAyRKT1d94/TethajOTTN6
KxbSABupUx5n3kc+bzhioou0WcimW+ufnUoUdnMkMbKVcP1sjcMCtIDPBto/zxW1NflUhmhwwFxy
VN8Xc+yePl51ovDZtGUtqIMqM+KlPY+pZPZJ6skf1uiGSneZpU1yilBpqDiirdzQLQKR2za9y3GU
ottRqrCbG2Hz3Pl+8NxaTIdCMl2FabSt0Wk9Iasq2WWQHBDEdXQckexYWu5kThvTEb+AODDSeJkI
F23EbzNBlp5LXOI6tGR4fpHovV2DOJc49HuY5LNmJ+uxcxX6NgXvu8lIzS9gjl2l43dwLZW5aSOQ
si7nDzqu7b06+YhxnRtmKaBHvKhT9tCTgv3t3BLtM9wxAXgAfyF4QsI7o9cNk7GcEMVOiUGYX8Ow
9oqKrzoKAfg/P5x62tl4FMZIc33ySOHtgziN4MN2r+w54xROLqAvcO+/L/S2Sla5Z8tiyc6pTNUo
rzQHSC8WPgcYD+SjRpA794PFsGq/J3aZhH98Z8E9aYO5MBd4rzxIoaCL+B01dyHPGz2reCamjApk
9QFH2YK+ns/6L4ZXifj072POivB/hqtdCpiG95BD7HsSwU1FgAnW/91xeuV+elbyI/+xSC9rBMs7
Fi2gaJdyJAxPrvdZMfvi1vHQEJ9jUOLSZz8gYHFEjoxcY5lj5Fy2VU01KfFzkCsA837AZk03t2cC
WxI30G4fwf2OUGNlwP0jGFZriEo930nD30r5l7dZHRajl7ralYmfxIXJJPeQG3KcmMjY8/5SVjnJ
Yt12DiylLLucN3dQnvJQvWYIS2Ou01rv+Lw25e8L4uRo0zIxp0Xqi+5/adL8AD7poCrCjZbN1ZPq
NMp2jhBkH3WMo8rgqHTOQ+PSHF/tPCixlunUKF4+CtcA1R0Sw5vq8I0TuZy5cULhpfaPlR8LbC+Z
OB5nbQhT39CwiRlpPemjwo73I+j/B/duXnIyPNs0a3jNkjNFqMB6M1v17J6Q5EL7RekHFwCtmNJc
TLB8TNuns6/hlI8YNHuLl7sLqR8yeKefEkOf4pWOuoxTsUrnv5BUB1DCjaX30MC1/vZsGHIfEO6A
HM0HTgg+u9Js8U4WSQD6U57yOthrYcM7r644K07PVrLmsPNbMZrDSq1nHRTPI10xQhC0Fb5ewUNl
X+C2TSJlcIW2FSXyUAzTPx3/dD6StGpAdTSTFUHEFTjNNXcNZfAE+G+AbEuqO/vsD5ye3BvHEtMp
WogH4wpilceARxCBq4WoPnv+eW5Mk6/o3S98iNQ8BGXn5qxHoNXY2SDlajdrpthJ/wm/9SYoqf+I
yz79LpMqZLs6jz8P3wwi/kZ+lzJGFFGxIpXVSUrdH69pKLzsg8QCv/GLpp/XZM3VKhe9bKnr7o+c
7T3mlFI4bJOn5XwjNsUmMmBb121uiqiwx/YWt6Y9g0N5jEh+B1s/nkgOQzhmcRfJtukoZqtgzbuk
qnvQj6badg2451SZItxcY4wbBCKonJDKl0uO4b2Mtj9Rnpdz+0RmApmxMBgQJ609GxF9nyqQaXr+
DaNN6LuA/tOFD73Kh3AV4EN6HF/I/Bfh/bY2XSEQU4pB99S+8KjkywTn78J1faaICMemJeJ3kJlH
TL4XV3AlZ+RAIGQc1ELhk9+KiiQ7AAj0zJvK7lDSmD4gTxfQk3Nsj0+tU6aAfz8YVpM9/nQE4Q8K
ogoxl6VPIl0oWk2XbQcu+gHB8O95kiyQN93jZ6vYlIqWiZ1fhQUikzyiqr9TkfMz1s8+K4FpAxxr
d4IR3dY2AdurOo5+TlYD6H5cXpOQrv5mK+Hedt3PSl6Uaujxx8NIxrxfQWn6alH18sZQz4GvyPXT
VENVqxWTM4ea6x3V71jcBMcuDtUlAcjhqh5qWZZsjsIN0MxwLtR9a8gOyF9onXrc+Bdp0/zLFHnw
nMjU8WpadVezU3CQs8SOuNm+j3fEJIh25HX54NyPo/Xe4iuRo++O8hCUg286J4ORBn9IaE5MeHec
bv9gK7MgzawGASClSlbqaw0YqlamngkuxQBBnlNjkXRU+rmK8edIHes3MHHAvhOyJKq7toRMUwdk
Y9MZLOr0A6jqf8s60bkVDvMJwiHDaAXQR3lzHgTt1PkLEVBUZFP49j0mdh+/pcYUCeTCSHre5s0Z
4p3RZos9A9zSW4z/ODpmOD/ZWskOtOMppLagkOoNWdnWyx5SRbYrK60/e9RfT3fzogsYtIc2/mu8
xSk2HWG3QN0iTpysFRN2tyRV0sVXHqelrz9U0K9dpGKETNV5xwXIlrVAfW+DJfHN8VDZr4C0Z+Nx
nm17KClhbRldlRTlsBCh8GIfc0d3Im5K7jdvQ6ubuMsF/N6CQAmY3oECLlm1FEmH+UGsXGwzoTFS
zADNaj9RxW3IIxxiYabudW0RyzLOz/k2W27DNzXGyrOqcNxTCZCBLyVvCWdTmQCmAw59oc3D/FlB
QnTzrvQgZPcXS/+bb7Gc2XiKK7l0eTfnyJNy1fGaRnXGCabCOtQuiRjb3RQnBI/7HUAH+wDt0JVA
hrrr0ZjEvreXJjmNMXwF8HQRsYfzK/0F2055KQnN2V+l6HO8r4tabwC4I2Ij2dX8j7IZJXTaA9bi
wryb1NUIm+2DSmp9lrRKfybldZhHUbJOEvI2I+PwzaE4DhV/MrjVSDYgIvcqQixWkI0Kip1gG1Ec
tPONBRLiSu+nHykuhcZvJX9GZUDJRTdaJNcmHMLXxO0a5Aur7kCjDVwwXPVZJZwDkJrxrgsSWInl
QopMgrnGj8uHotfMDBmppy3kg0eBGdCGTazKuKnQGlY+ssYG641X38pv1YojcUGz5LqiePGe1Or8
k80h4oA2blyzg4hq54MKSiMYBod0mA4YKPwm9xkzHktP7fMKo4dUli14WSJ9rsGjRPoHvdQh0f7W
EPc8/f1zb05el4fXa03lpqIxKKm3ubX7AtUDjql15MPivRXq7g5xTVw85lqQEvuPxg3Jt2chiNZk
CTR8sv7MJRB+5bT62wnCl5yA3jUllZMDcFBPaBzndenofKwUUSOWYkF3iMWnpRaKoShfHiz8cWth
4OadSH4xKPWSVhF/YWAWXIHsPsAYMIV1nDqZXz0o3Dq/aP8ccS9iUrnVC8zzaS1lOVmdEX95m+ZA
wVSWIAJL+dTpKUQDtXSTNUityncA5YniKoRNeSRVk7H22RSIyxHOqrBcCFqM6G6zfaESer3FwutV
r7abwQQMYDDEog/txhEmBQoU4P4nLI6WI3dWq5jMBVHyGZTt2Zxzkcuu0eOg+LgG1qZDk8QnnO86
M7IytCK95HWNKS+WcomZtHgUeMUEAb0n/MiM4e/zTD/wTOsmNnDDlfDjJPvRwI90QZlCF+0gHsgw
b3fp7ylTFEkTQWLO3PieQTL8D3wXzdeagD85578jpmb+27N7v9zshgaQFq5ELdBC0Kcm/HDuwQoa
B9+ryIjbv7x9t5/c7fL/Hmj761KtYBz+WbPr7/PnsbFOI02IvXQuzQLAdbZhzit4fG9QOv4lqvil
ogzZ9as2GZt5gGV/7BJSiTOyqEbqauNNmCDHmKpz6msYCnbwxbuuCDpif3LZcaWrmr0t92A4cdmT
lHRPjxtFeigi2V/aMzrE0I4szw/mIBczhhuP+5iWmj4tU6xoIClsJAIOVxUIHJK+Ujhacia7v2me
iL9MfulK94lc1nRV70/FlPQz5Cx6WXmbSM6HTwaU7cB1gXKA3W04Z7Hp7BNemdVYP2coWaQvhKA4
FkRsbv1ReHkbrzNZVvkLfqgY4MtlkrRpfJ08EBKDuqsLmaB/gvmrw3PTlfbgT/P9hxDk544ZJJ5B
lBnd80cfnuHIV2ZN6EYV1ZrmGH/R1Fi+xvd0sW3zJuxTruhZrzZ1T2ci8/dkFZOIQerK/Wgo8bah
MqhB9srYCf0evEYiMSN6ISJXLdgV4EtpW9ngQGC4dWLgI0rJpNoFpOpDTA3PgwXHzi8t7HTwJDwG
+3AxeIJgxBKMxxx4rnwqw//bBvgDNF47U8xxG/9wHcuOpsWsvtno2S2VjiGUdZKw0SNR0/sUVBV0
Gb+tpbE1pCCqvGHKEo/i7rFoVNQRI788BtQyI2U6YKJHmsGAmNL3yh4DtgCP0VDxjC9lK6UNqdZi
15UkzPypMFeDVFgYrDrS3WcBL8ff5Yx+k/OyojIh0A/ndD5u4P4gf7YBAoJsxPgSZPXlIsPGKQu5
as6WaiNNO8c8ffsZYYiNPxCJxCWJp7hvaoUcqGYWCySzBJmUJVO8F+GwbOUo+e8T7kKKcfMoggde
QS8PNdnY/SJQxylLlW5Xtk0rE7+hsQY+IYhpiVC2Sms4e/IOHJTPfzLeReKozZSkmYcDzLhbWViY
fQuPUbVwMlQNSR/njgF6Jr/QFqzh/W+JtIawp8MPTHuMIqDGCrsagnP5tXi1URnrIFi/wqX3/4ZW
US7q77sptoITPjztsk1I46NPpRmiu6SOd2YUJ3xDSnh5onTT+k4y0cTOR9gV4+3EW6ccJ8pea69R
NEOizykOL3ZEz2I1X+hLqtGmpqofARmxYqs7+tmjYfNdyPWWFfp5d4uP1e0FY8GolXXepxIaYGEp
duvtXeCXRZZk5lWpjV8y7TvRHJy/l3rohZ7otRViC27aF3XeG3lawceiY0R3/eNMrKRYd8sYhyzJ
RBF/I8630qE/2hv2SKZ4Fb2Mg/50FMtXV4NuNqZjbKUooLhEYuux1cgGRalr4eYb8Wv7/oHXnXS/
r8rTNl44dAN56EJ2lVGmfyDZovSG7RakpGq8a3ZVrn6ZYtRVdtL1QHiL5ve6GyULVy7MomToVRFW
aufVcyD9rYk/OYUFUXzoPzUY9Q/teRUGKdIAowjECcIt6FmM3PblYGrO4HSMjmt3nJZFl9FXFfnj
A927Twuii/fV4K0PdqDwVg3jGQ9KxZ0u2KJBbwlZw+/0xl6T8zn4zLKG+U4id4gHsV39VST2TXwJ
ESXk8QBF+bIWS8gsOZBOYtOwLv71oeU6rZyCzChGr6EtUiJhhlVkfTVB65gzWqrae+xZPXmjt/pC
XIik30tzjrlRd9ilgSK/iNzBKvxABvAzf4r0pdBtsXL4rfzyjReDBJa9nOFJFr9dmkVemeOqcuwQ
Y7T0+STKY2f2OeyohQ+zKCl2ti5ZDzUnHKnLjtVmtyms26ecSantzNSb5eNmwJmD9UmGcjV0nZES
FRjNUuy8dcuAS7JbHTzx6KxFO2JYj7UnsycU71kZle87GsL4DsXv7ySTeqVul0zY4x/pgRb9tVi2
1VgEZACXyaLpbDBslSL88LwMCVTTiKiOf/VGqkJ8xbSAOu0bI1fIqdJhD4+2nV+x89wct6pNOdyS
7YlVX4QaIYdnL1MBHw4OJ3lhU8SuyBXhCucvNLiK6n+E5Z3g1k6zDIR3r4RUX7VFikVwmuG/+wiH
f9mUl1bZovwcPegEPqgJe7VGQ/mOWjNUm7nyooHbZUuBODuOKaizDWBOF7IzE+2gLyZnSsE3IOfE
eZPXuf9TPAgsoGayUV1PxO6g+bCBlbu4QXQHPcxAslbc0hhQjOUG1EnmigrniMrU2PppyXQCQNbg
deKAvTS7WAcXxM1UcW7UoPzFXJq5mcW4iG4yurl7V4opMyrxpjyzYk0OukLBacOw2Bi51R0P4V6m
g+pK8nJ10tZ1BSdzXWuoNcDjNNcoWvi/nf5ro2FcfpvTCle2ivOUlDGrLkR15fHGmhqilVU9W01R
CLoyZksy1Ii/uo/Q8T15lF7yE5uPtx1UnBCLgJLyPwC6stIXEDc2uNkoTQ1R19jGtJakJHGSjJok
KuJeKwHYoymIIuSbW0vNKEEineNJxm1JwkZCSfsTsIvD9UmOprGTjJFBhjB3wGdYYCzQmaluH7a2
4iEdda8EAGAccXv2JgK5MmV/EY9NMluId7YIuwyzlcYvgU41l6+9QvCGlbe6YMsH+OMcVPmqbRNR
2XHEWa47qWAkHbFODC+QD+ou/Fzy/vLuZmnDks0yGBsmtE2mdiPFsknz2sIdjXBVfrm5HLi3BYqo
RhanwwWTWcxbaKQT7aeYsLCoBz1U7AaZilWxC3Ju/msXSOsOfxp71nDW8itC8PHauq46uhWRyhN0
xNlD7aOc1ZwS3uXTwoSe77YBtvhcpS8e9DaRSJ9OHsRYRq4poOhKhsN6vrhB+aWCF/94atuMjYbe
Z2GkQgPJxGRSsBc8+wCDEQOHM1nUyuGCrodPrPTBkFVkmXZDlgKGYLKg2nSsEqyZkJfxF5qK1hxB
WlwIf8SsJQcBG5dJLDih8usNL7emm3VIGBKgTPPQ0OTlBNS1PE1RwQFoMUJUC7cHhgcdLFDVOlm3
rWTYJwh9e7iIWP2+j8zFuxuHUUt58GJhC0gZdwQeyeKG33a0/u8XnAbhegSZ93qEOrMEQ6Z5XD+H
GuKk+okbKeN2BgFVxZa7pU6CqIhfutNIdCpA6rQ2AtnGQ0xELAtoN0ksZ+jDSfd9dyW4AbF39fXG
sA1L8CU/LjqY1CokSypUsWx5SaUUjdrduUcu2GOnoOdrVUI2NShpoclRQQNpkadPaZDbTyFlyh9T
cPlNK2KD3YUwCTCE4EUg7wQeIm72P3oLDeboYgodEtC7BgQYZrRd6HnNPSuF0EZ3cr0sTp6knMow
wo4UiwaaQPU+njh/q5A700I2CBhQJ+odApHL1/RObhOEZq30JLMGGwAnxfEB29MXsEVyp7VaqRVP
BCRo5hwilxuA1y4bFZt0SbabX6blXJlKOMMIwPlUJjWw0dBKl9rFWXqJ7GOvBQpvFdRQj07Hc0Yi
h0JxAsfmYnO+LVfbkIpzDSDyVwksngUPKEAouDMjZthBNn033Z9IKPd7vN7Tts8OnpLvT0IdJwV3
M7JjzENZpOB80HSkMW/Kr6okCf1EsaDBjvb7IPfrRstK0aOkqKzExORiQUNkL6nxPXjwtUxa35Ey
lXK68UJhNN/vM12nRbmFRrItJfApdbZqa+cMzdZUZkNOXmlY3OiMwK/sTUjAdKLujZSPFQ/Ct64K
xwNBKdU2nTL3nhbuZUfjCzOZA25zNkZF6cr49Eh84t0O/ZrAwehXO9uD7oI4mA2TfPClaS4q0Bei
z8pV872VUZHcc10hUMkDlMiqavTUwDamzhQSnzsTLjlxhJWquGp0EzAqXNavzggUI2QbL4l5ou1Y
gn6VzX81vQuKjx3rwxHm+BmscSXx5aDTymYJFU6zmnhXEO5CNwHu+/20dz7fpM4OUbX98NReZ6XK
zAV+QCt6DLOlUOu/uGm7XVb1UB1b/sdfsoR23F+uOS1fRn11gRRPzNRECgNIzQ+wqrH0suX4ciam
NJXiqqF0F1KiX/WPX1dgkCwdhP45hibL2YhigvXoQANCEN1BhSUxQt3o2ViDpRkdUZDcu7cl34AE
fMZ9k5FPgurDSjN5dziRz2K57RWPRDan7Gz+65SenSxEp3FbDAWiRgeDx9e6luBr5faJ4RI22e/A
kryT3+TYZxPP1mZVeP5SMLO2vCrOxBa67/jBdJfKdIjYSsjnYGmEQEZAoGP85hr5eZgtAiXs/Ag9
79ONmSkyJADN2jK5I+52zlWHU7pRW2G1jKwsrU4pvPBi1jUO/RscRJWbOSEEFzYscszlCf2p1ZOw
oiwgrpF8kMBaAzOkCDJsQYXHvUZwJLVvOvlnakzQ/z3Ee6m1JMlj/47LCRMaEV5Q1t5bGE/A4Eo/
JjvCiVZ+5q0xA1iwxDdFZcGFUNbb5tkl7Ujw58WLVKGntWH3urb9w91B3zBGDnlY7hRhFE1I4KZt
FubGWf9/ryIXlsNabEUw0ywyhlEQG7ZCJHTFYcr9g7OFnUB1pbIFXfJdwk4UGKDARaTX0uInxxsV
FbNBtEKpfVcdZM3GG+BS0MB7QRl07sZt2ZE/LM573Pn2C4nc9YhiXBewsJmTxDa/vGfd3+QmWfWn
d84B9SI2pAnDxdx+AfjcvgZaU+XhqYIoeomMXHgDzHJe3iNYl5a4APs837S7xkUufktJSAPwSKOb
Us1b+FAhqq/0tcE1zjT/mABU3WtYBWNAXDq8FEWVxYbSip5j31TGmr5Zn6v/cAbCYZpqImI0TVs8
CqqMZ3tGtmlhOy7cNjF3OdtFAKKUlaegF1IUw4hrWIChKhSq/r9E/2HuY3XpFua8zDv0O3AqAia5
TU/Q6XnP7BUdFX/fpXCrbZm1nFaK4x8S+Dt+AqY5YmtgkFm9pozSzmBUTH3hXtZ/jdoBhZThF0hW
v5EUJWo3rewMvSTKDVDU+0gFmqVXozvQyyCzXHWPyyVIJezdnrNKxS9dPcj8txaTwKHA/Fl4MyyN
lLwMu/rK/97kbLP4jF5yQo/zb6jJiK2o7NfY3kJdub8iP2qvD4WxoYFaEQlSfeQZV0QXUpEF7/Wx
Kd0rwNvUL29T9YU5Rl1ExlUg9d6ZYvRiPNqGLrM7RFkephrviePYeVoMjjSLmZlGaNThx2s0ACg+
pChbhhddmvGQY5VkLx1zNVx3o+7CAgx8g3I1IfeiyglVM6Ot1TMwpPKK23lx++hyiWecTByXro7m
RRKVQdD+nBe8D9eiVa1Zv0Z1hpVXJgdk9/dljayiriyoSLiytE9+lVyM09iVYzZg0jYltBHinOPA
9COBb8pFBk/y1g6apVGc71laTkYm0g8ECnmsKV5vBpxDCJAHWnl4tg9/TtdjhfOkt/yKI+iD2W1c
KWmOqLkyf1l6DVvRjvcGknroUchLMpMXSrS396wCEJYLpg1u+0ipca4hST1vnFko1nI3K0uG1m+G
vV0FO/rb5bcZSmxfM3z6p7Ql6G0zowkUl+ecrTE/E7jmKpc/hDacs92p/PBhDET2vEKr+j2s8m7N
6LjCtD99ZP4GyuR25APGG7y1eZAayStQh46t1M5IS6dWLawYBQz0vLFnyze7KUap/JrmnPop2XU+
tw2ArtgaRSXabXhNCXqgMHNu9yNxmB1Yxg2rki9z/af9f54BJ9K6MfOBNPUGk1c2wtaFhmixeqTx
OAPZ7tms4IJuUeMYK3p+0MxOarIcVHkHyHOuK5/70f16z7+iwjMHgQxPkQ1TDRn5zP3byXmHzuFd
y8nFK7ePT0XmFvDHu4ePPhJkkG9d+oNdKWjfwa2GKlfOOu/Pwk6grvljbYLQzqG4cBZUTecBFb1z
RRW7K4qphz0RNYF2GIwRUVg1JK2m36XQjlcG2zhjngRYP8Ed2qQmbaIP9x0AThSd27GKy8sZrLrJ
tuBFWtrev+xjyF3nyEa5BwiXl7n0Cp8c42FkbD6F7fNjp/a2V8mKRJf/o7C5p02Vmb+mJqSeS1eI
pa+cyYUlMIkTBOB2bH6ALUOaBzUaFtJkMt26sOBKU6TN4mIJIKvh0V3DJLyv4wmwsZotQOLjlQpm
szJexETChSn1K7fHBvz9b4aD755K0VcLgVKDRKV3AvNHd3gWkBGMIBjsRm7Wi1tfEoJDOMUAg9v8
NjUiwuGxqSk0iRbMMrZ3puE5QAIs9/Fkc7uUCO9Z5/uLINm9j+FlYY1iP0b3ov1un8mQyJCBTAhK
wFNF4BB5OQ4nFECvD1fbe8YHleo6YYsozOpkFp7dihfGc4QBhrgwIkCOQg9pF1aa0dZnlpA7A0KP
278Gfwjr8SKP+4NYIFO86xJBoQmHzXBvz3AH5fEBNgEhg5und4WcaQIP498BPskexRkQNQLZVBpK
j7l/ELdDCWl4Pkyhk8YqZXHk1r4P0jdfnWO0OUtemIs1+wPr4YoNa4/Un0EFnDseiM//R8kkSVTz
ONLxuO7mnORWhxHbS+ZJOpPAfvU4bOaXjdQT27nqLMqZ9YuOtbkGSXiSQv496tmmlx2x1QlEEROL
NbAzgku+LEQd4X1ARF4EUTn80IxDh5ldu85fl4YyK74UTdY9M64Pyx08deNqft1YXppX0MoLEJPO
VqnthAutSu3pfZdRganH7H8aVnxhVV641yJD6fk533XARvDR1dvYcjZBg2S9+hCBYu0Uppn9gxpn
IaJ5mppavEEVltB2hKY+FXyR2sM6JY+RA655va7H4Efc05GoRn6b1geVFnALG/wJaU4PSDEuvYQ2
D4XrjHBW6C89Ey6iSM3ymFSHtPmmwLys51MJeBOSWOfZZCtVc/CGf+P9v3L1dNrcyKnjTk0RXX0/
zv97osuvwI6Qyn5kShs+5LkCnQtr5SHcfDRjp1S4D40kVfrmnElJJmZgtL3nk47qnp3momf1EKEb
tlm6mWv8uYCTtVkAP6WH5JYGIp5/PqszsMU6X+xnldYv8XTBbane4XxfDBnANKO2W7u5To0mGpT/
Vw7lRBj/5m2+aXkDV0laBUWLlxB6wuiN7BbdVT8G8i0WzntCFpiz2iLPogMwrK6BzJkFBJO2SXnP
1VYMaexalTsp0mM+5G4jPWJbtr+nkiPM45usdDCjweHj2TBPUF/VGY60ecyvN5ueBXQq44mQQ0HB
mNUNvc3s/239inhAwWBqWFecU51NGEHFVHhaHWK4pmxaEzzlmptiyHC1LwLUpn6lpj42dGnNwH9u
lTsV85/nZhyCOlxca1P8R3okH/l1XeBkvToPtUHlOv+Ca4o5eVNywXB1/MS8DjUpeth+LP131Ua5
o/8MI1tvP4UK5lptcaCvpRDH1GK5CTL+zx+6+WJXGMbMjOK6+yejwlNhXe1H4uVdLXL8jS75I39F
t7kQfqi1SsAgbqANtQ2TjoXR0dxbWmZxUS+MpwPUONti5/FrL3zRcIWWPzcZRI4ykNqeJhWBgz6B
ExbOJqoTdh1A8bjRn7I5TvR1d7pa84GZ3kNKirJ7OBJpFvDGVpN/SqzdWrlsQix1NWlxAOe2u8vb
6GMxXiWioyQh+V0g1TRpA5+hvyu5YiFdoc+3t0l7R3z1U1xDCG+POBLatn0rjJ+KNbQouFX/eofN
IRtoKnFXD4YhrOUTeawl5lRwUoxDxkcnFzR6CeSZBlF9Iz8sLaw2g1vmXX+KCepToKGzXo9hAwPJ
nK/9XfhPuBSlBWyknESUMgq4/OO9dnELCatgnUcntlyicAgn29akp303cDaPHJx6UiS5XhGYdlQp
sF8zVk2uUOIfcIq4SqjN9xOV0rJley1eIDySQi8x5CKwjCMCNhoZDWNDEe3WjPFMTFlJoCeF5F46
SZm8nmQ4H3uZrumvKugfvfDyXCv9Sht44jr2LZ4rbRD3CGR88cgp18aIgFQ0Hb1E3rCd1ASYb3Kn
Fpl9+qVU3iNt/HJeVdbCz4PZs5WNahMSogr0NDmY79qP9hHj0gZ74AZgNOlxTf2Bb+IL52w2Y4eF
cEooSjfURWAbzSznUyK79FsFw5m0vrGABuoRYM0gQiSp6X9sS0WLIGcBV2Obe7F26dKQM57zjKkH
wSab4O7DD6maOvvnxrQe71nfyR6n6cd4k7/NQMaaSKkCAAfZQOrMK7dTuFEL/rsM57QOeHp5MCGA
UXPzZxd8Cn2HHiP9oY+B5B2zIug1XPvZgB7kN7p8yl9me1PS3SE7ZhH4VYAs1nIlcX0KyGBFpanG
mjHyzgekLsfg/SpWc4c7+gaSBnGC//V1SIB9P+gIvXQx7nkpd2OdJbbJfF5m1hxPsgawi8FI/G0z
sqgD0FxkILV8zThI3bwEnNCUu0p/Ir39Qb3LbDKbTnScNcHcfBSXKPvILHrFQXUQ0sHUuyzA85lh
/46Pil0zODvuo7yycY60BLl0Lnr+GQT2/2GCm+Rf78kWGazATMRveJaAiaYxlvYmnbUm1jeoPbj9
f6oPtLB9p+FlN94UgTMCntbKG/f6BWE3HrZZNs/RAcjR7kemR9cagQrtzhsAjSumOLGXZMNe95Lf
64wlqH3R/CFyI9x5VZGV6S7n5FotQ8QcRkD0MTI0zJke8QtQo1hWU35+iFnS2MZN/NRvXZfDDRQ4
R7dZPtXHt+Jb77tR8KaZKqOAssnGOmV4XraHWADucjNMeKEbn+bmQ+wzODqbTHnxfStV+txr4RUu
3kl1hQomPeMtWUKO99FphN7PJ02/GDVXCLWQKLZ/VOmtebnVQdt8nPMptHLlEqSZ26lPNlF5aK+d
Gg9OlXhsPsL14gX9IUEVMwKhhZSUIrr6yHqnFKewsYq21cq9Y0Ku4fZRpRYSCO8pVQXs+DNfBF0G
2BxkC7dtQ2bwkb8kjVFyIXb/+fpki90G77It2AW9h3HEj7/kkDxDF/w8wOtHkvAx1AlbHbjr40rF
TSbeCnsUmgDPkBR3jycdrAcaJhdr2poGIj07Tz1aDW98xH5L1CdZQbkb67O7qDoGxfdh5CoKVN2J
sh2lwsVWmCgA3167QWqfKx2fxy+RbCrva1tId4n11Azo26MdULaNXpp9Rtz9rx2NTZk9l3nNsbH9
nO4P3ql5OzhLz4KtlzUGYhPD3qVNr21GzmVCGGrKHCnRFioPhQ6At7xqSiBe2yH7WgFHQEpnujlH
Emyh07BlBGqtwSGD3t3bibd05EIu9hi0BfAJnrXzyctKzoY+RPhRPPVvKXTJhbbUd+0SaYIJiYu4
9XUpy80v7qjITcqaxf1GYEcWfjTGgfsh68CLMHgutk/+0mRc9SGxxvJUflNBMMNW6J6p0EUroP7Q
vKmGe0Ahv6sYSPTSlUsiu4ti+8A4WqGiVLnJFMgQAgbj/ZgEUYuvqO+gUfKLlXRiKFFgMdJkSY0J
CETOhGQ/nudpQR5BxjY8uIjRZ8tsyDtROYCI8JsKmud1QiGEgEoGO/DuQL5irXgDeagg/CD4tzA9
9CL0YZDn74XUbv+ZOq+BcM2VZ4GRxMU/mZ8vKVvMz5i+ZH2n8L9JSUPUX0/ZnWwi7H3C4hCYXuMq
F5E91sxLBNnQmFAT0qRipo45r7qgIkZViqRrz+TdURgtI0ZNlUwnfPkis9MN1K+0Dca4CKRkFfk+
4WuMPyHMCHFnVx+v/hW0OSBJ+xWGE4vVrc/7IWaTpuRKNFH36dR6B/7P5TpJfcYxuwmfVT7gDaQZ
G1RroLjSb+930uv3JVTgGGkZ2i3dCb7AFzDHUbuXWseOJeDB4rN3Yi+Hu4QSi3ycz3fgxqQMxGHD
rMEEL1PZt9Rje1bMCi/I631o2H8fBiIb+0fuvwkli4+z4MhgDWBwygXFh7SafNs87q4IUw+DeJCJ
wGI0SUqv3tYWSlOLuF41Dnb5ySlpWX+8CK/CZzK6hAXvdw/lqgwW2XL5kugiSeII8W/7dL6huYfq
+4bR8YaGj+JjMpMD1wbi7RxXv8FaEDySG7aWJOZyahDatL2iH4D1taP5kplvmuJQWXeaRy0oD7lT
Jg+z35domiZM72rY1cJCkIQe4byyqeJwLZuJCpxhuowoV9lRDXY5AIjfietKCkEvCDf4PFvVqN/V
yjBmB8rqf/Y5QHVlZ1vsSfurZvmxcab+LR6URejTrkcOyrYQmrHGkWnmh8ermwm9w7vWHDqJfbGF
uLzh4ibapdL+tesVWhC/VI1p4pTWVNZv9vcD76PgMvycUFEGnTd0bFz33ebf/LU/fGTXUclInQMC
gfnu3UhG7JUij/jKfV6X3MU1yQj6HhaLuH3ZlacMAsrz0y50KowvrTJHOs0HLIy47vxfLNXpAfBM
Bewv8dI/uQGl9hx/aJBEmjxPplNFs4P8mDLReyAyAX57Nmlsz8zN4uE0iC+qyEp0K0jFoE+mHLBb
Qy1FCXRsTJlcGGA4TNqJj3kfZxNWXGUWOK/7CNtsIi27DeyuvjLFKQEzE2QJGI+ubav03dTJixz2
PekD13B4LidHYHqm9mtuAhv+YySpwXZGCCHXMCkZ8jjxzbMNYUoKND44XT/A0PtaNQ9R+4ZFchfk
vmQ3NjzudRuptOhpuOkuRH1wnDtqcvTlp6gu0TrxV6fMeG7NJDDYmevcfWRSWfBhz3VG30PjNA4+
/6KY3Fg+eRR54w3jV1U4PVG9RUEPKXNygBMD8j6TrWu4Edkt7xFbBlq/29VX2PoaW84XBWegaJgq
BI/ZZ4ko92iShe4cxUncS7ubWpZXMO9Wb/9wBJtABoZOFV4hqGSlfsaUCWpVr1UczuZesjDptosA
GCRcChV4ESVnTnNEhnkgoU/jmSzeMwhGb7/ML1bYNxrPRuRc+oWbfeJtmKvVWfNZIcQkzCeZu8I1
L8cNIRkpWK98wEsCrrHshE6SBe33y9bX4PHLho5ysRMIloX+oAjUYTDPQY5vIUpY1J4LhlGfqM9s
tOSRh7Wrw8PHsP3QbOrWraHMw2J+z13X3sILwCYVSuTbkPganjT4fRBo6G3KoPYCOuEDRbW5TspJ
KRMfDyUJvBXp8CgpQ8IURPbp1DdT0kUJ6UKu1/s98cKe+R1Nx40tVU55JZr4hB401tN9DrX27h3Y
BV9Oke1BPOAOxKgknQ8w6p+f8w4kqeWLCNj6hQti3v82K+XTBvDGwzlWzWNFHUdQyOMItmco0ouD
tdQC69oxssqiXaXs/j4U0Ny+wSPYASe6ysAyOyDZqZ0yfNbyQgvkh039zz3qtBDnEmtlAGhXAt3m
kdm6Sd3fUbLVYaKgYphjJzstZJqe7HfDwKqHKVceCh6SGQG4DQyQB2yxrp2/hqozEJU2lVmuNQ70
2wjnq0QPlO4+ubaEPvtn6YUOd3pri1+ICGhXTOHbqWy3IsVReDs3XKHdZwE2nCbI4SRaLHbhu+WS
DUlsonVwpzJAqwi6VwaK1sskvleK3ZHeSm67ER+QHBQVyiNIpWqkiSTgJzfTI+GGI+fqyj7ie5+B
bG2cK5Nk1EJ0/ilGC/SwFdu4uEF6m1j7UBt7nB9uedSTbDvyycRKHx+T6vRNBqW6EejaxafsQwzp
NtiBuuGHt4OG9+dBK9XHSfQhd7tUakiqT5RDO8exp4eIkCAvwEHme1QabgNzXSUzGdSleFw5FMp5
TBgXRyFXcGZ6WOeSzJ+WUN7DfcTRMvrHChzmQqPP6VjQ/Vj0w2NXu8EbuCR6mGDqVSZczV0FkZU7
YXE5FDKRextROCEKW20nQj5JFaJ+KOZy1GFuN3dwWlvZGdoeqGi9FhJOZ6d98VRjHzTf27SIHjnb
bw/i0DdURbavR20lng9uzjzjydfvAAUG5JPbXf2eo9CvmPRZqG51GfsFCnW4JAn6x2FZLbc7ZatZ
Sl9iDMPZrei7eU3s8QAgw7I0WPoPfR8iuUhI3q/5eivhQZ3DDty+IeV+a3eqytEIfw4GuQsDGYtv
6mnk41Y4yCD+dTanNiZxkNoV6Xyy73nSTTI1vTM6ZPG81moWkXpTlIme2An5CsA+EEsakkox/btW
EwpubW8z6PeolmEnRFtse8ytsYsWrziKy9ZYoEYPnFnOYxlR30s8o+N4n0eDMnmhxUXZFXHibI1K
gM79c6Q+3uQnYTPtAI0a4tAWBrtW084VOt97tmGJdMfbVC5ly3qKGVtZdK/UsY7pooGPKfbuDQQl
SdmbLOcq4REfYMnGq6Kqm5tI5msyDczna2aK9DSqONNGjZZ1i+EMoEPvP3+FncTWPEu64oTItd21
OhqQxmZX4bexewcVyvc7xpKx2y5nHXlUPQzHvcuuj+UVoojejHfEtzrEKmmd4Sqa6xmILROlB7/W
YqvpLyNhoPoYEGkZWA162oSs99LXGZEicQ1kTG4EqpM4fFqRoPDrChpborRhxcKpjYBhInc4uWsh
W276I79+ap1J1mqgRrKnZsUjgBMeRmkdBT79fZS6cDdvpDP5DVsWEJ4YldBhJIkgWwbIgz6rUvTQ
vjeVDLNSNIrfl2RT4adVKOPy+4yVUPZtA3fWZCS09zM7iMWpPGaKhXxXMTQbC4a7YWJIe4tYGcoC
HbYlSxEPv2oOLD+k4COu0JM3YjVQT/cVCRdwxjB1FhhQDEuUZGZ57ghCWPRFQu7wuKtYPIQfwDtT
8PpVeqcbyNqU7Ax0RmfJTEttfcCn5zugDH2lMGTAgmV47lrmNLgK/05LE3K66kOEMf6hrPTsct+u
9YAwYLeD1XS/qDpJ3cr9PjY35lCpOEadb/74m1iqf/G/gzpO0eN/lxxR6UaWDeA2yoI8lN0u+1K0
YvGk2CdZKwsJy1Rto428CEFPS5bRG2nrMRkjzFOnIcgwNjkE6lZppDSq874CrEF0R4+rxxH6wsAr
weSTO+ExbdkAcdc0Yn76Sq+ndrHuA9rkoERw5I6xD8tER8igyTBGpZYFSN7CVFgBm1Br0UNT/EWd
rlYli4UoYoC9V4vPhzHeYEcaZrjT/nE0qqmK2cn9HHmrLGDRRRDVV8soiJ0oQOCeDU3s51dFObwO
4rPdycJvvU8nXj1QGeyFLINcEiDHpGcjOMRtPPCZTLMSuYPYwKeHdS+daM7Mp3cxCW/Wn9PWGtpb
8QHUMa2kGvSU3EGAoCRb1ylGtnRF8cEbGMnMLn31G42b4UYb0t+IuH42p3lv9DfrFkClv+83LSpM
mZGFRsikrlkFYERQk2/lrXa8j7UXvReenquYejefUqN9nL/8VgWijDyO7tkdD4NMsif116Z1g48x
NsMF5pAsLKWvODpVyWYcoECIZC/iRnUN6sWiMKJ2+rjiWILJVg1aKDi5eugmkXOqaauKwTRqP5tj
I4zjke041YQ5JHqjZ8YEdUyOVF/BPR6OtCdZ7e74iil/XiOnzqWA2Ldftjnr3Nj7o0dQDjgfAxE1
17xweNSVGQxGkC4UNIbLorrtNVHPVEPqFww1M/4iofV64o2LsvBW/Pmg7e2qK0cc5GQfjmhAotpl
xNuxAV0iCJpdROCR9r/4USPt6zAB64B7ailJsKM9QyDwiy6yZMcg6xdbgHj9c6EwsOuUzt2FUZQS
LRG3/xejTPmEgMHyP74NYEznj1cBstNyR9jRXo0AJcHwVMQiTMYtUId1xMJooA7rVzGC/Uxr3uht
RmoBTJfkOIFhlFpEuuQMJOrHpLvQMKLlfEPaa3/CPl1OWFMRp8i5NqSuYdxTLW0/EAh8I0wy+foe
MsSg+wzFt5U4R+Q2fol3XgH3Hqo+bKya032I9Bo3M9zs2K81DSfHgJuHKLwploFEQFTX4r3irCeF
cR36qKoqnEsqSqelAHAU7D8T13W8mOxKURaKooNwApVVTtcefsMbCRP/AFAualYdsIum8TpPD7iz
3Z31f5EkUFrMpnjE+ivXbZ8tXko79r+NU06xoaHCPheoclpygjriO+fDoV1iGHIIePHdBtjomcQU
sfxXSZP7RvuA3R42yUR72yVQ+S0JalfERw56Ucxvd84FmmPJ2RdvcT1651fA06VTlo4p96kkCeTQ
Hw1fPuhBdnlUxf3zXIwx5cedjASR7hByJb/ZChtk+Pc9TRaS/5I/IwSKhOTFQkrDssOR8B5oYpES
ACIBd9rPMAd/ASnOeQKKIOs64kw2ISSXYJXiqQrGfmh06doZD7GNceaEuoBPBIONtJx53I5nLyqs
HDEZqOWMRLvTspf9tHPFONi7OjUzJSAsnOFpAHeUyiQUW430M5X7NY0RsUjP3es54MfUqswwL8bE
Ldz1BkHyDt1+V5Q5Y7/0kUqBqvogPLH+5RzrnNKvJxg6VP5VnZroSAh2+b6pwaiG8AR4ZqQwGJYT
I6cTkOtO1B+Smo9xzOzSCoz6LI9PUTQPfqdyFKWMPUO/7TOcXYI8z3QWLcNiqZB9LRIHQhFWL/A1
A12Sdzbo8XK44wZTZDKkbkt6vQotXs496OV/J4FWn5dDom68XKkioRyKbolhWqhTx9FOLnewO7Jy
TnxfK38hR4Zlujys/jzNK8YioN8xlPL4DbeETtbUFhzqsisG+5+juUi7Bo98tQD5mK34KAhYdNRX
0wR36C+PlvRJpS2yLzyviDDY7qeQ6DHLklb90SGqOrxMJP1ve6j8qIGtJX1Fh4eEZ4QlLdTNgVQc
hAT+H1OyqAAImNgURP77xbaaZCW7o1sMZuqbbg0iqI4TsnsKCiSg63zVXwGRcw5AaHVWg7TCMh1G
f2hXk6QHCbtWy8uTb0EjDi+U+kPszc4IE0ov9ADDbsXUqmMhUApP7SYRsDh3KVVGcyp0kFsok+eI
5Oz4Q/cOYBVmqmt2cXBbCUHJMFVxks/saPrWT3TGHRh741veWXogb9ejLXZOkS45qLeloKBfvlEF
dl2Jo+pyR0o+i6M7fZMrKUhHXZXdqG584OOBNlI2zDr70Fa0oNI4wy2Yy4e6nkWjg6WAWm4Vz546
opPBi+9kSJ0BSxBYRrDAgYhMRlxFjIzItuO473jq3IE8GfKPDKWRXHTFJggu6HiSZDw5nSPwtYgE
J77q5l3JhDgpH6Gmq54GoKcRETqIE+EnMlpO6Ev8/r6GcTAcqMjV5LigjwBzN9rAHRkkKm9dGLQ7
/kXEjD9eDVx4jFh1cryaKRK2tShkdCnx5fGD8vhCZVi3bj7mny6WScpK7GVwcvhO4f5ILH4WWYdl
d/i81oHGcws3tpuKclpjOnuGurERIUk7qDVUK/fApVX1CumBQOQ1J+HhD64a8La5NOKiAu4V1TF+
/jsanCulhkFpV2pClbSzQ9fRlU390p7pTIF0w/CcWhhnUvK6vMfD2/XXYSYScghmz5nWmjxSyyNP
6yItLe7TayZA2tHAVSrNwBejWsPW8ydfsk6Vq4WpifRsHxZV+FdY6ku6QcKQutzagPoNk0Afiacd
AkkbM/ft/0hio0N83d9RJHO6mVoV+6QyNuOuTHOR9jh97l0SDxSuijAV1VslmDAEGLqTW9KBJH7s
fWB47IP9enwlxldkMNsVEhV6CGc6fdOEnDwXx1lxf7mmf1yLp4ldi3caP0n7AI/lkfTJUEaJ6kZM
Ag7LOx1ovtMTJmF7cUfXnTGlvz4rVvykYDzmmO2To3Tz7qactKFLYW9Deemu2AGIuK+asG5nOhSZ
LGT6Fql7nUYRC/KwY0Rv7Tj7XcvknIvoyKTObRfPVh4v8Te5HRh3SeS+85PVTUYRn86+qfPrT++E
bVF9wET/mHVrxbRWJn4JsvseHfJdfkP1sAyDFbWr1m3k/6+mnRxvyZC6l6QBZoaVR8h3EqLThiKE
sXFQnds24qCwwcjBDvMnIjAoprBxWx7LNewIHHBoGqZ83IBcOUPyxTbwtZVKvOqr2HorF4lWfl0X
EorHrXzeF020tVc/L0JO0wUdp2V42d+slSSn673uenydQAXZ1AH+Gx2agQOOtzgGXE3ii0tuUYZh
MX5IR0/p5q1Qmpom7Aj6QYdM+FDYq9DMyH9QnSEzah8Xt0Qiltas2pOHKbfwv7ckSEW/2vVTlumN
40XaZLBavHaioqlYrT3qTJBsqE4GN2xXXf8Disyd/K+W9HkeOREv8FTlcJqakPcc9n2Hrj1Uzv6k
q7sNBU0U43RgkS70VfkZBPc93oTXnMIPDWFu5bKHjtMRI8wLQ9GIKJji98NnCVF/A/GJ+Uib7yaW
O34/yunPKiKzfCIcdHto4hprzUvETh9FWMC3oCKk3ILMwtXM47fM6Kn7N84if6JMa3zVT4cBiKJN
TQuLNH43/yYcMfmqRV8ycDD1BJCf6q1YTPnnkSZ8vlSnVCbt4tWlCm2lwteHA/07+eRzOpZjGNCH
ZVUlQZH/cX7faZ3/iJDa4Q6blmHcbOUxfCr/0+GGEZIRpU1a+IM3lXr9da7zQOA8AtZwsozFDcOl
nPLyKjjvcKgmoXoUg1wGiw3VL7IYefE1ey1U5Wdz2q+usFMu1Ma/JwrQuUz1kiLzPqZhdAgitHMl
VYDKh+5bjd8SZrnJlfPzmuaz7W8pXjaK2F8BNr6S5+8iiReQmwVIkqSI78z8EVmyeNBEqr+zhtkl
e0LmZjw0Qvgk9GLFJD8likjj0lwVnC6RVo86XaYKuYcunUHJaoE8fA+91Tz9lhitJHdEXZmVjJ0F
VjuKiZiUAptLphp9UhOfJMefYZdjsXffbvRQZh2O+wnFlxxKoLJDe5a5eJ1sHXU/AsxhPaBiTo5K
ggn/piUEqGzaCxPxc1vSFsErHrFwns2yI9VgPYXGQPW6BQKnF1nCv0EQUB/VEcKRy85Hfs7sdOel
/sRhfLXToK2sSVdwQW3/8SbuD5JecbBzCt4K4KMzVl5QY/hliBiTZdMnVP1YcFluRrKAPKrYJVnj
CZipvUuls9IuqkVZO0kJECmALbyDf/j8UljrG5iIs/9MiSwqVr6lOeEV2yaNnaIragcklWsEWxKu
N040I6yG4N14jKyBg8LNkgqM3yN9R8EE2mk1bMPG6t0gBCXaaQFmAkwFN6jTtYpmwOO6uJwGl5p5
Et5XtE3FYICM2cJuJV72g6Z7gq5j7MmgmNKAbL/NrvCgckdwrxlv1rzY44pwSRR/eVOJg5/Vzu9G
EvzyU+TrJl8AW/O4rC7JXrkqC4j/78VsneVI9Wf72NsiZtQOg3uacTyJuZxGTGx68BoXBgsEoEOt
K7Az815mM/AR22CmCjDE525JEvQToz2qZLTTLbXzFbmvcGETYGdIQlpMA+jZGbZGVc8XBE/oR69K
uPNXCJhgV/nT/GfAZvmO3Nvhi6GCfslzOPB1T38O+8PzhqyYSQz2PHTRVUSnudIPi0nOySeg7taT
c/2G42hhmRAxKWL1Vf2n6frWyQ7ZgeS2ondn1zi55c9H5IxcZWJOq0N/Uw/vdMT828CyG87LXage
fgTwZhZO6w4TbgZDwXJgS1zcqCPaRlOygYQcc9rOkVwG5wNJETp4QtNh41sTOFvLNkavt5rB0LQU
fij9wvMtO2bPMUwVtVe5+3wOSYonTJzfq1PsijGKPZ1iNAuRlGFv7qYidg6CeQ+TZ/mj5oMFPVrq
eE9aclTl2nUtdlim6+/NAs+y+yghpX2FgM5J+yCKAcKnaDZs+qHWU/GZF/aH43jVMX7TZ09KhWGs
THK2P1rpLdbiPcP2mSUrqnIQEjFvROKi9H4e312IXko8/kUKor/5GxUKIsPQRhURGPUThhXF44Co
cNGqb/Hq1Vqr8+T6HJ/nUtupZCm18ujbGB9eXRmzU8AM36xwKvx9SIGD3LN+8bvpCsLQmrj8lyPE
QtWmzQ8N0BKc1FPX2hpufVjYYR7+EpAMLKfbMShG8ML4NhdHog7Yn6vsmI5tJCrRxQ393VvTes70
iKe3rDztxgn8sK+QDQnP0jXvfbz+herjdB13L6icyUkbKyvvmdazBBXQt3n76T+ccUpm2HhWks+S
WSDOKFewjm0iiFskITbyjhwK4aQyk3A9/ajura4AfQTuiOjmMweFrtjqoUS2EL3qUIYWTyzBBQdK
1YvGEYoQKOp/GeLte21rUE1KgT+YTZihI7lx/nKGSCLehFFjxSTPcvFv907zSTqbf4PpLpBKG8yB
W3g3z1HhSWVu70ephhtYyRDDvUJ2QmZ+AYYZU77GgElaQuvCYccpfppNHE0HYmPX0WSjTRROmaFa
5N4KKjM7fl6QNftfbcr/y8sDb8/qKCPIBCAHZts7WUa6v/FRQpI6yO1JvEXruOzkIyh8PyqEo71L
c3WeQEfvge2k1bN8gBZ/znjTUWzaaQpHOSdY3KHfz/trToLrAmxtalkaMKpU9W56zen/ZY2BAzsG
Nes3C3S4naMCAzr8xYLf5wfz5xUlUl5lMCSgQNw+3dIzOfOjyYM0DHgdlYJKHBgGEJqHfOA1HqSs
P7hnV4g+OtxHCSoJQurmB2I4Jzq5mEFVTUIQSZaTd4JhjLdb1nRbctvKYMzxn/7C3pol8hYaNYAi
hI9h0sEraS79noONPYhsUE+X+82XRckDSQRGIip/jzMUr3l0Vs7VvabcN+NPINXGUbkG12Qhg98a
983gXdWEeMgextFkxA1b3oNxpkpNKK1D4w9Qdbh+vsKPMTuzHEZfIqT+OC9T7QW2MpClsgaEjhd5
Jz5di/XmN6hkDMczlZNo2klsZOqEc0zK3ScpvYU7d2sSYmHUyfhXy6utTEfj850kEhaB/FeSJDLm
OcB4W3LNNj1LkcbjbMlrSkRV86zmMDT9Ur7gZq4jIRph052Hhh9Y+EKND4DYCt1AI7sIYP1K4SNj
I+yekgyUMmabk01nR63gStWtgjX8cJZdKo5iAnWEtM0XJ1BcCAgWAM40SsxKdin27AT9jG/kEBu7
t8RPP7YNCGyYbKtPK70yvwxZLzXkwX74wqRbxmaQd7nsAdYr9b//SeBThqlKvojk+s304KNoKrmZ
hnc6gJIkHeui1Xg0Mml6NYnmn36FgIWgwnsrTYafWuKBV5kE9ppMQhiWxiOI/uR3J0n4Ytn14N0e
xheshWuy/DCY7baut0u/Txe6KmtLeaNSL38xCU5IeUxHYBws5XWfTi1WMgynqeht9FGhAORPrKAo
29YRSvrRtKPPZ99yL69UEwTS/jdwsRLobnpw6NxpiTzwJEOONQNqday+TR+ogfJBavS/8XM5bld2
n+eUliKFvwIiZaAOL5UUA9LmsZe3Sospe9JwSM51ygQarOSbu8m5Q3oAbUKN9aI/GiJZDnMeapnx
44oLw+YmjGZ/9gh8ExSpqA4XbRaYfCDPikf7jE8853a/12+KDXuu+ldD6u/8S1uxq/csGuVNPoXW
9egG3M/otGACKx3NhlitUtK4j0GTokCN6JpHUWJIO18y8kafB75LXOSanZ0i7OkJgLa7t9QeAqly
dxWXc8y+hTfPd6JBVilWSsAtMJ1jXnP96znnnKtqrrX0754sSjZvPXJS1CDYQ47qHBdQBOVfpuXy
LTmDZJzD/tc85VzUsnO7weijI/ySL0S2SiODpLw9bsMkSDBv4wjhh99upjLbWQZjLX8k6gxE8+bs
kydgwe7dLW8u7MF0jKPrhLIYN1kJKjxQ+XtWeB4iI0zV1fdD+9FSUnRDz3BEffvv+D52iPqwm6Vj
7/jS3/VEIPHIKwbKb5Uf2pHLPeHeH0rU2rvj/r+SfQ2VNO2KcJvcRJ2pl+cxATyUtcxrnOqkQzYH
Cz08Td6aK7MrCvsYGb9GTmnBKgUMgEk35UIZc83YBkDHW41vhPu8Kpadj4MTSqSJGVd7LH0jIO5c
UxWtz5wFdwY5nOe4kJMN2XtX0xqyWpMsUmO984q2LznatsCoH8ozRDkGX/iip6cFSrEESqp3WYIJ
S4pjIT9PbEhBGzzbycHcx3tjFPaDgwjXf4D0zEhWIDznLSSvbtzTYbth1v72dcsXfJGsICVJj47r
sE4I0yhiI8+c+Wg7bePyVQvhoswCoUALKZQL70SoZ2RgEzdJzB9Imf1AIQK+WknwznFmZyK+Nb00
f6xEHWjNeopQnaEPq88BGvjewNDz9A7r+X6qypAOLpr5/o3KibgCKDO2l0gJjSX3OoJhDrwgNwLZ
t9fLtEeVdP/pvON9tmtbfECAZcl14T4zBs7Zcz+NL8i7Z0lOUg+R80qBAz6orO9he1OgHtigGYjB
ciZ+7nrn3C0g7iY184COvER6gefIlWEbSx81gUzJSapkkT7YwctYjIZRVhrcxosvouUGmCMAgKGc
YfvUQNNFZQIQstkuBLp8+G9l8KYYVTGqeRZ12pf2Bsh8kDPlJlc+tfCmSu0eLVKSI//2LQJZ0++T
AWF5BPC06UDPZEAOmjpjiDTYD2blkAIj0eCs9+CD2T1w9Mr+rXoy6ym6kzQKUw5uWTEoTsjU/xPQ
zaHxuFEOVID5OyTueeUEHjHOVSi5sIfwsxeGKHX8BDBYDlxCq+q4LOhaV87kVXgvivVqOSJvcePy
SGq6OLqFGq3dQfXo1KNxHoghdrkKd0hYeKLRrv1SDnob86BSpHTWzGpBVkVKoLMgxwa4u2zbpVtZ
Dk7lXep7yVS02ODJJ9AR0xaIHuVjnwzbELjng8EbqKA72BxYhC6rg0PbUt7Ryn7utW220Hj9ihNs
bGT/EaTqXyasRdIqApHZ+sc+fWSN+udk9xdaJDPk6788Mws39jMZ/vz4kr4ZCPJe4SFoNPQ0yHmM
OTaP4zMzmZf/YO948m7Zzori2O79cyjHS4kTWKFrPQ/Mj7IIBIUKsQygEAG4IX/Eg4PYZbK4rDtZ
UeMFUXMKmLMJczwGXqwBu8SV3Nln0F10sfrAujq07K0npYD0rRLXQjRk85tPfqKzi7BJbEixzn4P
OlfnSfbtjuSmPpa/F9Rva6IkgPTknEjFZYlBz88xI3/yrccS3T8SFX4a9tGFFa27Q69i1Oowy4A5
XysmWeSxVmgsJUkz3BHM+mXMawu7LDjJgHkJcBU5jV7A9IK6O3kx7eUpBfvUvViu413q2zUZUX6q
2O+ORmIh/80RUNNIFY10LzEYEeUqXjG50CAPlI0MiWrmFj3lMzCMLLUT/BmaYiYBa49qD+0hKjrq
8k9vxBoZwF9GBwZUfq7cw3GDktlWOOvBVEeIk8FEqd4HxrK1A9W5J8FuMgKppdnwEZpF+hn555Gu
us6PX9KVGDbMnaId3HpVBi3bUgia/16v9YD9Tqufc3eRSLWShLiFGfWdezDDuPaxMSuR8ZmYilcW
8ohE4YzfCDGFI53C5wxaQQvdeaOyJS+xk7+tuGv6NOX6Zpp0hRoQRLkXQYF+RTzByGaywlzYI/jY
A7QPbfwB4EOozoC26ea+h7rywRY1uOpWbVZLZVxe5835oF3qPNlHQ2hPZ1JOm/DGZloHGgrT0/uR
rFR+AQDyLb17s3Juo3x9fUFyzVmrDVag59d/0+kuTR3iR/fyN6vaYZgYmB0gZphYp63G3dZUbFKu
TLGjd59c++fTj5JYfZUh9PoHHNJEMsauFI9I4mfazXjhV8y911iTV2yoJ/TM8InM0lgUgyq31ylr
0/xw3c6jGzzldIQjF8TGI+GiFDDNpLjRIN4nZ+E13y5tDINu/hRB44M2sz+eViT0FddJtXmeIYnc
Frduz2NAnrwuq6h7FWBncwLQvYLBfgFN5vzTHqUrEElmL5n/87rKM7IVr8ELWIllGLNOte7L37jx
bj1V0DEQU9EJcPuyonrRTPd6crqbCh4M4W7D1Q9vwKTaR7oEQ7qO35QbGOkH9c3hwYVdeM1X2PWG
fjHwgGU5IAYn1dkhCVk5P/c3pE4PFNScd+thpj531CL/sZXQuwTxG+RlPDBin5RHSI1aSDXNyHHW
bnlD7xRxvU1oMbw9wawreHZBzAbcyOZrN7DNgaPx3sOG6VHYP7IP2cfMwus0+V5SqZI8rzf9WM2H
pzSBugwiYv35+QudJJ044hAkahal72L4mxEKf4SXX9XkBmEjFhfIhQSVx9XmN2gcfa99cZQsfxvo
HTJHcnSzOHqZ5cCPW6t8pzt+C6rTEafDFr1rUHx2ODle30oRSF7lSo+trQz3sbpdsNap9/iWEDzO
gPJ2On+kkaVWyeRKE6q5jDpD6xkle7n0Hh8wctqPstn0T0gj8lI0aqECazdVoVlIMAVHMlGXTw5e
K407cj5m1K5njOLt9yJoDP1G5aZ5vTEjtg0LTw4RXHa4To+VHLvKwDevQnVN/cPN/3FCyqsEWU9j
+dd5vBuLPsqk4qmH2o8A0fjfZ0PNxKXbgQuDETzF9JXzuxxlV+Li0aEIrVzqmxt23p9JoUwBFKbO
qYZWgZTnLs5/YThfjA9y52g+I0RJ5cIFuTTArKJYnZGxPZN1DyxHCJypCgD2pdOrnA+ZbhG6PDQg
aYEv0y5X3sHWjaqVmU2IUGwN6M4KlCCCpWJDLXFBhWHhmnF402L+pzwH6IDwYPnnYdE5mF4sdqY0
yIuiI9mxEYpHg/X50v1tQhIp6b9x1BrFZvpBaPjxUP2WHy+Z65XzWcgdyyUZPnJcROrAEXsDiCQL
oeXpe4cFbpwiCrZQZmt+lC5kS+3ZsgwVBhZEviwIXSlPl378/LJE0dxKxEKWemmn9QbSXspwXPW7
ags3cvRhvR9dvZuLD2cwF7sSWps6LTuazZehxN6hWa1GBOpN6OQb0B4LZnduE8QKUhSqEnXXvyT6
Qypvdygu9OQp/8yDrYdOtx8M1ByI3A6NeSyKVpq36foUM+UztFrp0mFq+EQsIXjBuS/Kkq1gSmhX
koeksspwMJ4PacuKZ5LxyJm4xPe+AYMMrX/wbTZXf3ogBH0Y7IBjhE8lBSNuQJbi7dEQ+K5nh6e9
9AOKDRmGs6cbPtRRoKEDldRRuFa9qgwe8RvGnL7FkHg4DhBKpAqTRYslN9BcCrLFgsmQuYUYhsvb
impeVHFaioAT4yDQ3rcgRQu21kMStVK867ud6Mmrrrfv/LkhscUrqHyyznt9Wlwy6m7qGVedYGT8
AJMddetqbRZLp34HzXWkl8e70q9rhIVQHvjoDJtKEJoPL1/bTbRwE5MRkQDuhbLGjwcTCHSanGPr
ixAkqw5nyfEcnpU6Z9fHIx+tVNA6deAQDypLQ1YrH8YkKd6yL+1IM3V9QZUTIgLY/4Gl19iTX5w9
i0QH+yFqeRWqbg00e6+ZV3CskisPyt5SM7JTs7kH0w8vsxc/yZ3lOxA9v5kbCyytY4RzpM9Q+M7L
vyuZ+jp9BjbjsRmvlx/W0qg/HtXz0ZCWx+rxceA2AacHjt6N5d2I9VJEC9b4C1g6OyOpUO23Nhq6
nZfVmzJuEcFLbIn/KHpjs+T0oqh4Uok+Y/9PohVVie8cf9dkB2+FsXaL3VsQwDshwi+kJkEWNkxy
waEOKtnN+bXuDrec2W+RklE0gJiLg9O1LfBD9qFsl06bmR1SMPm6gbGtm7rxFZpN1jpnEtP99Lsu
MeJcAGNLhIrMn09d3PLZIGwXuuXSBUfdSN5y11xwLQkUT8h50awi+sTqp5G4oO9CQrbJwsnvjy/W
52oadQYjpjmPTi9UJHeVAV9+UrHQZcX9HDxbHSEVCEXUCk1JctnOJ+03oZxmXLPYHEcilId6FL9U
p1VkEUQDQRQQeXSG8lgQGMAZ3u4+HB6lUXgNp6314et9Y6BDkBuRSd7+B2ZLoy3q7BRm9l0J7K3g
NwVgP+i+eywO34265Z+qyBCCJluzFCl4FGKqHwuhTSSH3yl9B6aI7ON4fzHGnVCYKSiK8XmXxU6Q
CxmFPpFUf/+g2rne7OcCTfDPBVQxc8bJzCoIFfIeo5I31IKRIgcyDFC+rcal0p0kLJx4CZBYY3sb
RVFDgEAd+ySUgtwTjnRI2Xbnqnw3q8GaIHubgYniwZFcADe9T3V22nLAG+V+sC+pz1zfHYmGnR6l
vhcJw8k7D7cNBE6i9+Tu/GsTOvR1ZMTlg2BhieIvmW/qxEj/B52YMMisQ7i96Z3yQd/MIkg4+aF/
g4eYDZmSyKIGWKTtxyq/lHW3V531S2r0VVxKn7ad5FdyESG45JbNe/x2iVBC0cx+2F0f0AJWFRYt
+qO05yvbB0vfiETHq0fV1kFH5SmFtFz6PsMEzeM87nHZDVzKeeH/Dkh80yaaGyT25w0I23Wlh00K
90WFJLKHn45AAKemT8ojdinx71mEQ6ZEPCXl27YAfNAj2yubmwYAckyS6+NB9NYcSpKFr2IcNnkC
Kf20vnQ1KRWKuKDosP+x2TuMPhuHbwJhv5Hzxhiq0ktBZ/zhXPhbVUoLV5vObndMWDDhxqqn4YvV
DBWHr+GG5i+wzK7JUR74iIBllGPpqiHajfBzHNw2UFfxaZ+7R+OPBQCi8uLl2fYVgmJlNHJD6U6R
Hp3SPW7QEsUmO14AQZHej4WDrbj/8zGg7smBLLXgcFZkGoYcIF7KBhRdKRcdw8R8FigjmSyJtf8F
HPUTrtNCmQrYHy0gcvQun/eZ2LFqMmFdFiCwzPYeut2pzahZwAiELr2jgeRvy2I+C8lbyl8h5hk1
kiPWonakaiUy44nHdDpC+7ZqAwaEiAED78W1OU+0VSnPR3kXPZYpwsRkR+qa8RJlycsUwMyv4Zh8
FKGt1nxsKSkD7FyS6fXJepRHHGvjxeL+ymLJQUajI5KzYUY2WzqtQ306njQKhUHLw/mSV0hQBsXv
LZ/ygD6Btg0N0AIWrQ48yKt2FGWgcW+3cqX/gVi0ijxjjMnrE+XDTV4bgnW3nGumZcUPKM2qcEKL
U37qqJ7mkdi26+JDxzJgbz9uaXnR+n74638L0YCBZzZG4NXiCCcgYXDVG3Avs6XLYCF6bwr1r7Qp
le4Q5St6f4EfEIJANlyv5gim2Q2GPIKPKFbZw+NGQujMPTZKywSyXBV3k4aVMjKbhhMcUo22bdHg
LpPQc9L85U+FG39lElKQsE+AWp/kBNPxr/GR9FdFzLEa5SuIOWVabZQV+4rBlwfO/bYRykSyyaGj
KKb6XJHxUAQTLnD6+KMhdoMZHzEBMupjB23r+wvtXGww59KMy5H3ntIZ24DMlDMynavrqYAumUPj
2YxdZgK9G1f6uVsOAp088YGAVCXCBix5Izbb663GSRDzOCVOUuvYUVKWDh4Wet9wGMtZiJl0gGL2
2DPPFfw2GD66cHA/RCg0WT6iqoM42epEGZaabH7DK9LXC5VvKuLkTxlZSeyapFnjiH2IJ7ABb0wV
s5L72saym/lAAmYVNvyFGD9/llZVdPs8IgvBY6loetQyrftWKAA8kycSibRjdw61TXQf13nAFvvT
nlKSwiRb3B8Hne+WKweLzkL3qJYG4EH/EtL9FC3KL1ItTH/56S/u4YaiyE721ELuPEu8XU11spBK
ueWcN73ESM/dpyVDR1md271+RN2Tzcp/z0Pn6agHnkUcT0pi2mAm60ZZ3uA5D47fASb1W4aSHNq+
CnChNAaDsKnB/IChOI378ckLdJpOLYUauzbh0vEAGx6RL4aLTn1Hn3a5q7ACmVhJKsXjWPD7v3WB
dw9K67Is9V3Zj47og6lMhq8MtXArkIygPVhYLfUebH7/xZ86BMEYIbRDJaTzpjOtcwzBkLH2oYP6
wOYSJe5yT8DmVf1n/aHI4lO8d/GLC/DU7OtyOxfAPtGLdWLmWUcFvz1ZSOviuINyhjoRz7Hq37Ok
+Pf8G59zCKFcPJHYNOoEGSDXtTZVXJvpHmBMbntYonjJoP4qptmRUP/Lp1RtK5dtgLSZF/HOGd41
tsW+2iWfXUEyVe9Veuce8+Ln2XF/sRKCBbDo1+55gOfdXvPrqv/CMrAuQkNkm50OquuRGWfpYvwr
CV1+sp/wHJd6VYG4wJJw5aNSYCfV5bigmcg5qwTGVn80KXsbJV1QchYEpDh8N9y4zYuR86/v+Qwk
ObwqNebk/wkA8KIh5A7f8xssuZR+V10j64RxFcDj69F7bUPHibB05aPHYxg7p/gqDI8olYyqU5P6
U4GPJSVWvBMo2EBP4mwV/isf+kdwYkkvjGfDdOefIF+4ZLk7ipbv2I/CHvMSIkipqO3WxqVfO2Ju
yxy3ANZP5P+A9LqvhCPZr+detVMOYoK4579WVKP1vCqcLuNaikZFNrkMUmCOUHa+YjkxSoj38Baj
/5kmd35xSsPud7w6rvBlh0GqdFAIeF5nwFZGcUUGe/sHv7gLVGm9S+EYbSDEFzL/6BBgYZ071rx0
kz/VPQLQxfu6kwIfLYWBndg+Q0kZJqFK7nlBUdDJGoJAlTjPHI5pRlrhP2ZzMIX6NQNvgpy9vsKu
MMVzIC6NfvH1CXBaIuLRIcu65j49H2Q22N8twD+72514esQRCqCEyrNHYcMwbtyCqcvAGffz07oo
g+h2Cy66g7OR1TxqVyc727itPbnzVQyFgwuGwV6+MTNhtN2C/CuCboUVEvaB2vjoYPle+wx024ME
Wn58jUmKdrsLQY3ZAzk//vHgto7ZBXkrRdBh56a+ha+gw6N3n//W83iHC3U80Y3939Z4uNxjzCPt
wS4qseGFICGdqhGZdqgagK22jT1dN00QdFmFdTqbneGkLshaxSwWhkl8M7I66sM7QxdyXDdHvD7t
xJJCRft8QHQOlQIGvX+7DYJB9f3ecvDI7BheaQ+bMTEET6Q+nhJUB3gRaqnMt4nChC5pe03jFOuI
MGhBDKwqXkCRL6IZ/RsAGmJPV3Q9fB8WzKtURk9DsN51jDnyhQzTvYcZpBEkrXUySs9ouEsQUUEr
dcMBm9OdPKOBrB4x2lm+yct0+UuIIb92814a7gPKM07OSWb+0u2x4sinkTx7eRzjDhWRdWdL41cF
wPdhyddDT/1aWAOUGkD/M7dgNudTM2lJEozwOFbzg/UfNd//nFX6f+OJXBZPLuIg2GgcMjf3AsoK
OkBaCpZLYTWio4dP+cyFZWP5/0zvoa8gTglHCQOMyqDlycfyxPcvJC1ESkmnry9+L7AMpshzqoEH
hzo787o7aeJdkaiQVpZ6MoikFWsRjJ4wq04XDl/DjInz/BUBhLWN+niLV0TFVfjEth6JjrkTxdhm
XPGeA9iPtOVg+po9KKnt7OYX6Kyd7/Es7KaDUyNWtuQ7rmDFph8DArGoovqEY9obdvPkXtUlHcIW
1eo7VLAQzZ1lNRTM0WTbSJYPDygwisuWA5kFcCVtpnIfXUIXmMO80t1S6bB+xaC8oU1P1NM4yFrg
WkDNiSSYf7gFRrwOqtQS7mZC6X/8jTlO4xD/Soma9pNZZ2dmXznnv308aKAcaJHM9hlzXJLLX8f3
5eC3BrZdgEzw4T6t4wACJ5Vupa9Kf/CsdQkYSMZualwmpQVdPDtDWjTj0z6EasGRZ6zj4Fm0idQd
8eDLSpdF0kfpUMTddCMoCsoncmt2DmEWgAbtYoehYPiO9tn0+d3PhlTrhIyC9wVAMNwuTGWM56as
EzT98ZDNqiKKRsIYfc8cgQLhnpd1pR+ZD0Y0FcPglIobKQBbaEl6v0w6W6WXpHclZnImRlhTBwe8
Wi7P2kUUp06hgs/lq2FhCUNyTlNErydYu6I2YELzil38ctdIAl5NOv+RQUfWS06B6ofRS9WYQlpo
JYuQuvjnPtIKFneiWDgUmWUmcQAh9+WYdZuJ9YOVrA68ImTH9yvGTf4gH/U3+XCBcdw6K5fLNDCk
sQt9zWPL5yQbb/NacSHudvBwXK3n0r4vucVzqBswNFTOESkSeJzi/FUNWeScHofQnxpRvpW78zkA
dZG7pz6dtX1YdvmzrUmeV/fEs8MIhSM/bhQf0SICIkTcg/sFfOSi4nhy6AocQilaJPaA01ZiHu5X
tioQEzqJL35yhFkM0MvGVQ0e+LGyBM3Pu33z2HH+Nbb/TpxqxpU+m4xTTgr8N5SfRfD8a+pROfzJ
zljWGs40KZiRtYBD37I7YQRAZBBUBweXEMTlaN2eHcg3MMi7pFvV56eliOzPFqzxsu6H2g2Yno7s
lEnWxS+dHht644itwckgoejwMlxlbj2jUyBeIXUoZLhe536roi4OPD3dzAQ0YJj4FacG+dEAGuYB
Dd+6Ru8r3EYxEtywO3Rw08RzZxPWUiMMJrxg3Ef/ZSBpR9NMxoR1MrDtp1KpEHfirOSQJtl4AhBi
APW0U5sq+PFqgatF2iBwZw/WaqcaAkdH84BDs8PWRVvmJGIbH+4qE41P7hDV7Lk+Uyi72AEzXRUX
yStY/4NnD7YXmJFKNv32d4G3Dd2fKPKDMBzd4Pl9CpGDWCcQqCQnYUwk4K1gz61dvl19o/SuilVF
fpf+OyvgF3wvxKUXPyeC7vnAb+jClGAybaBDfCCixgRVi2xUaMcGSifxs0QDrHTiqbOkQN2Jgqw9
C7N2em9TxKYVv3NCTPeE3+iWT3eHME+I8kb19MEXQwZ/iVwlHYZmYh7oShn+sfSwmz1t6tpkVcu+
X54A3HW72PtNHMCarZu5Uf2AmBVUKJmJAWON+sh1p6TnISZxbbLr7q9uIUhLxKP10cYjkHGJdmcn
EKDnMCUgJF0PYRKWVLuHA0tt03wQF6SBr1QD+tW2azhVX9/tHAh8X+2zDOePsbvnO2FksSfIlbVu
fs1jK7MGBn1/cbYnKqY9t3z0P1YyMybwmi6u+gqgHItXQFOdMis9e+fJscEbL7oobIC97iSZyKRc
nLUOoTSw10TnIIByVlVZe/PREbP5j8egIrG7TQqzaCqEsStS+U6pH/rbcTdjVAEpkLYczKpI6Wex
8hNRHXHq7fovFLRHUT+kDpF9JqZivPcOrBo08vI8U3WBicFdDoOB+a//v6/ervQlJH/3uH7ud3Ol
Dj2dGbWKK4KrjJmF1GV0z/KJa5uaPMQNQUajwSKb+5Mm4wMihusyuI6XlgpjNuv4Umqw6wZ8yjyO
m1srNb2Rmf/o0Q9LWLib3RGNdWMqVx6jvvVbK9EyP/ai3LaLJCCJFWQ5fAVKU3u9wI5RqFfy+QFU
AUuQSfNeK7dOVFhTOiKCVF7X5xzNtzXCAI7gbqjR/bjRV1Rph70xbI23iv2CD20/7MGxbCgdBig9
dyNj855SDRX3JgmCw7KEYVAi0i2dmhSJNyeQ+gDPTbs1jHnb1F0QT9AqmR/MX+yeoBM23Yae03Iy
04+x8HtF+QiOgCkJ3VLt1hYm1oZXTGnMBjm4PLRwzh3WzD4R43mn1PzWMpvQ1m1AGWF5jM4JQOe4
V29K488wKpJf3O6X75myk9Fo0sxoKaKp6jgU3bm9AGtK8bCjOfZNwe4aKdcK35Z4AFAhpdM643K/
dqOEEYx27fKErn4si6m6QvWqe/G8rn6+WKREwP2vHrn+qXfYOxQQ+diTk577YI5Hssk/MrI37gs2
ZYZwzVdLKMecwkuMJgCCOGaiiuYPq+GHskPaIx90vvK6u/mkdrhl0wGepaoyEbms00/aLmeJE+bn
bSUGREaTlkRbaMLS4L0xga7R3nJkceEtGv1hz8sDxuXVMNIuG80DfGu1p/J90k82caaYAKuyVKX5
MdGPycO74j9C/R9lZL4rXs6gdeDP8al6NLNQvKLdvT4/ZNOtYWwxYWGdkj0JUtYj4Z65Eumd7z+5
qPt8WuOCo1HyBji9/Dfl8FSNrVETmb09cHiInxsLaig5muX2ywyHR4l0knCo9ElX3RaTwlUC048p
hHUtDBRZyxQIunUG8DIvSRviXIl5M3H6Hh1Y1SWY7KUqFyk/Hf+SssM9wESXFWDeb9DumYZOfZNc
4FPQz4vnb4UBONsmkLx+eRhN+R8cIqBCyyXa2ZknBouO5/HY52wmXs27f8noQqmdPR0clzDTKPbT
oYSLmVdQrY7lzkoTqg6IkOHiUc498JtcOWHkpNmZ5AaYFLSTv2Hhd5Czdch1Gmc0GJvJD1jhxwIo
lOxulkiLv6PII9Sg6lnm1mI9+WFWIWpMeF1OiwMbBZX0EMCWcnduU3MFCwzYnxePrZ8WUxVgssFp
mwFEjPrXq0MBJEAfjFwsx1xSmtUBSnB8A0vcZB3C5kMmEamkpvoJ4o8emkjJ7L4zw9Hp6/UmdZd3
isBlX3U5fBwXOCXZMszTg0Z0RX29LSSq03ERlPVT++8qff57br5sAZsEr6XVMoGXXAqjqNI0FrDl
I/xG1he6Po1CVjOwaYNmxSzbfxGKFGeQT9UR6CHl0pXZDW8v2OrG2XmXr4LGf+48vID7JgsvdeCd
E/Mwb+UxwYBkpZOuyrqjnAL5KHiT9IOhx2ipN252TYWBLndPKZNFOjl84kU6KgEbQk/aZGqCjOK8
fshIsI+8sQwIdyp7ARuWjdFHw8+sIN+pswoYQa0uXz6AYHFEF833gfeZ7/3uUCBacEjGF+IJLyGa
vww9a8AKczuZoPsLzj7gN+Q4sfSO4frJzW3QZGZcqlWXP89BWLdqMnP5wcwuVNUPkK1hMkHzTHrS
7flK0cKzsjV5WRwNftNWy3WZ2Q9GV9GhK1HRPlWTnhlj0FEtcvyg3mhtzUvG8f416nNcoy6L/Wk2
jUEMTRP5huPO3hpuTQaLFxfR+dZdZftFzZjYjMkr5uZkKc2OwJPYIdbx6ThFJ/8CwmlcrxWn1O92
65WvamPM/2teWU9TKY+ZJSvR1GRpQTUZQbmx3L00t2+viB2vYWw+mC3HG7w5n4qZchy/thhoxPEl
rZSKhqRjRft4y3KjAN38Kcv+K8BI/awijFyqcDULfS356sqxeeVDcECaTRX7+ST9a2/3xzZf10cc
nfFJJ260Bl/USre1c3YbdBTrYzv8FWO1AyPX0oQByycM+dMIIxMr7JCNln1cRlRF7lofZNq+Bmwy
0wBJOznLucVo68LEMELgsbwWpRc0MffZdIJbkXumje3ockKaFL4mD/HMFDuIVEDvx4tI5r+dlHnW
aYR4v5XaHQfL282VIv9a1/H4EeoC9BTr/ALgbfLQhDKip41Rccr9Z1CvtUsXQbthYtt9chVYxy4o
Y863bV7Ov6u4fO2j6t+t/dSM8qScOw6O4B1NyjZFJtcOJS1wDamDyTRsPFgwomaTQiKkdpjdB7pc
Ay88ksyXdVVT80P6d9kJa9s/efDexrSGv4cTllUhy91RyTNpj4oKpo7k6Oftn/pBw/dP91wwSlaA
JTEnMF4SnDWUg9GQjo6RrNgYiZTJKyAULZyOwX9NZ1RjZ4oqP5hEXcdgTuR7MhcpweuYmfwSSZn1
E5SuN09rK715XTNmHzeUSd4LPFnUE3GGrOJc9aAPkrO9kKCaawtiVg+rW3rwdbhF2PIkdwZmVjAB
Db4RF5V/B0XnmLFeloY326MHSWRCyBQIswf1HdXWrAMVOKER4HL5474BD3c9nH3pAfQYSH9wWA9J
QYVidMsLA46jaxn+QgvxlvOafeeNOUCJtsMlvgDGkjgPuQgi9jW+QOoVnhI4bvaxAlaHMnyoH/e6
xJo596n+qiaavGstSusLn9ii3/3SlLeXyg78tmjLrRSuj9O9ed8Q3dAUaXa722wenmsQC75mUFRO
xAF7Tcy5z78KMXuqsQqp7FPVi7HSsx/2DgvluzsISM1B2WQSa5wT7z40jTi5zUKfrE1gUge7ASbg
HyLZiVmVJxvyX1j9gGHxgK7+3S7bmHaKeNLjh2HnHcVubmBup/Q+4BWZjd6KVSX6MjT84IlUEFrp
SPGRfaBr+f+KAlJIXfGkuYFHosAEmkPah7S+kqBzlytNHvEbX6EkAdDU+ZlpXl2mzOqqXOd68iyx
+y6Ex2ZTzy9F8MQGwG3pqjRzalcQwC6yPNvJvPfq1xmsXAKp79NlVssvkmS2jIhHXTz2tfwCthhV
4aEHsOeZ8V3KajMd4mFsgjAAven7xhK0Yq/EUpPLnImJKbAWDKsnFWhUpJwaTZh1IUuF4QpFV4J1
5zGq3l4IaOjsuyQzztEsqyqD9kjsNGsLtXAz4tV1tHkdlEEgoxegvGxpRiCBpP0C/3o8Pu1Eh75B
S0e50dWKeZh6KBhiEgMG5gpAfikduJVH6lC/PK5HcsX53HWn2ALlnaz/nW5IXQbaV6IgeErwWmyM
LxAZ5ICt1Kn5oeUWQzB92j7LvLp0OezC38x/XLdsDTYSDTg+aRLRsUq82b+ZbgYHhN23020ffiBk
JlAfG7P8iFCXSPRlwPHhkl/s79yIQ7jY9WmpwDkTHScKTna+yfXe8OxCpKw8NzRggHoK+cHCSxrD
RYhxHEbBy4XYg3IctwJWUNCMs9bOC0tovuT85wUI16E3kCAX5aCh2hHvWYLBgfyZjwwBK9tUlSlz
WbmjP0L67oyvhIDy9VYW6+hHzwgBh3n4SeP/uqDDMcoMNt1Y9rQA0fkEf/GWmsImAF6pE/tgOGn8
Q49sv1aV9BxRbheLPEHNX9oBsMhKx5Hshjp6Z4ZJYM+1Ss2N6jwY2yVm5DzfgjioHmV8YV63OxAX
uyhFbQp0tBmgXBqkVOvzeYbRColtnbgOWyVBzrBLt1ab4ynSrrQ4bJOzsuRYtzYy7X4VJ8r0tkB4
Ue3PAGTnBGGjFT3lxUelG8mrZfNeQV6I4mFusZ0B4EYetWcGCj9PCRo0j6LALm92Y8QwjVOm9LeW
RedPh2UzuIIO1AJlskjsVeQlcUauWgNm1yYuVaQZybG+N5ZwAWgAt71uPrkVeSKMptI9C++dP+Sb
ankfuaNXCp9MWLN5kbrCbrnVB6bHYDmN+zNFgkaSmx8s6IrVKoiJk6ScOw0q/ra8l2IPxEKCUmf0
fqAuYvJN0p4Bzf3Vq+EMUHwPI5xhqha45oqmJVIHp7XZeWhkDWJeIwhzo/7BjfW+3MKJfE6c5lNI
Tv6RUsGQ23aqNjhgdmqbgjmCQS9qqqIRfEsn/DooMLDYTo+Hg2SkiL3/adAtYhwHUdXM9OTbF2eE
gFyLHJlHMsNaN+jVnOgZ7AN30112YNcM9pIr+9NABcHk2BqtRwW42C0ry2upWvp/uO7TrpbNNbub
Z8lVPDQBV1ayvET7eUvxahWYMXiOF84t1neVPHNbaTwxDkHLRB4fdQJv7she0OCEYEWtVlUQFtou
ExmvY+9dtVIZtje4do9Qop6jOBW7O9kuHrkXAmUQlAIP4lmqGndwtLo57zCkW0I8ChpMD0MC2xg0
I7d9PD2f0vVzOXLUE1gsVKZ5ilfXzmJsVhpbpbFQBeapziw2mED+rz11TM63li0F25T7FScABChv
moCbf1LxY51aPMoaz+/MRRi8u6cwD6TvEB47RtFAAo1ByazUNzh9DU9vXdubFlKh4wt8eYyRYQkn
50VgoMNCWmsLhl0UXMdWHdR27rAgvHWz1L2vQWtmbcnV6ADYEdvNBQVeRZh6aZ6v48u/G3m8EA9o
tG/3kK/iOMFNsNODUEPDB+RklxmOPOHlwFAxCFQ5N8bIX0RKtFKHn4TAfGI+pyXNd6PQtZUyYzc/
iDg0+5L7g3mBcZoT9KHam9Ip2x6O+CQ2jORP573yhq9lxEuzhUB2cYQHg3w1FBCXS8EjTNRBci9L
U/EVN4ytFkRiO6Ck66hm3OR4fqcUYZZ71ENhtBTS/m5qPuNUIChmIFVAeQZK81CofKLr36KKjVZM
CPx1H14qYEPv+sMKRzD0wLoHsGJLjZ+NiaOYJTcO+BiKv8jCnc8LrlTYWVefWqYAhqO2d2C2FQd0
8of/a9O5KMUorVXE8WUujsAv2goKh6vQUIPwNz499WjdV8Yq708qe7IaRUqPbwabtaLtgnkbAszy
j3zgJih1EMTrv+7pFCkiIQvYg+G4/UV1aq5MjvwOdrft5XFHaZetATH0eh22NzitydCYePH7HtQc
4lJDC5+J3/+t7NJjh7B97Xv5+IGtd1wQzHnXc/so4KIlbKDub9rnJXEYxeoHq1nZCd5b8S3tgbsS
3FEW4/ffLk2X9+akl7YTlUpjPzI9nxJ0OVMs23EB5cYhWe/x5JiwD0rsIuTT50m1z1NMp73HyELI
0BTO5+3pYognO+CNutO4TbBlt7REo4GXpsFXkVDOdxklsYeP1m6AnfKQ8zxmo5PawPzYe0Mj8RvV
YJxMKhOrB45JVKlx8O9R+ZywC7pEzDBdNfw1eG3b62rUk5Rk7tUt+WoKD9tP08Zw/RG08de3tBSA
kwm0OkCItMxw+DEOuYK5nWAtSJY4+rvClGirG0jUKi5s7M+VmpoBDWMpSTRS5YNpPtwlBsuKI1/e
sABLpnpwhP3ikGpPJg+0oEJ6PZ57v72SDnBFTIWcYNzhUptHJh93E6Le/7UpVSFJEb4xF1RFXKm7
skAaYssC4vUVHuOAN23a9iGZ1FEZPEWWvZS56p/mHdhyuHc8s0wux54LfySIla7rKSTUDVJF/5Y3
+f5FGvvxovlv2ZT957RUvFL2xR3ttKvBipVQcvaGKALoEexUDOO/Zrzw/ZGrsL82Cbxx9CNP6PAZ
prXdyWJGiGvbfZHKK2HoK+DZcBdhrxWJj21uKPQczfYr94lhoBYU05IpE1MKOajepMMln7wiktS9
hvdUS5gx9hQC1XOP4+uWbvwxfFfBqaPTtsdSuS47yN2o+2W7zb4dwOcnT6qxbsTNlelLv0CrLXqK
Z3aZiFzEYrB7B8YYAaG/WZmB4MInJKhS8NwTwxdg2D2bVY/IPkYfkC7lVqMkMn7I4R8QtvBnHcn0
MW2TvaM7GtIUvxnYpYbz6yn+Z+HIZRMpgrqYCufvH3l2w+kiUCnLE5S2MvVhMhot+VXHN/IHAJV2
70gg492OHYDGj9ssXpTEOBtOl7zwx5VFRxsU70xchRp5/XKyX4wEqmxV+PHKfsNFjkq+nSdw1a7H
+VFvtMHtSyknFgYMyCVcuVa8KP4SCPu6mG5GSlUHcgjEwdC58ZTzrj41fgln7o8oCDD2Xc9sfwH1
2oa1d6ej7SkKMkLoBmq8bZQKZPwmpBfNGYMwCAavMcru44pma4J0OqvoxHX6iyA7enZIZjXoZ48W
OxmS8ENuDCLUhzXGt8hoJKytqPxOT7dboXABYWLyBCRZW4/sak9qNmeNVLPwsVpiFrFXxKkxVHpC
m8RONeGYA0KGcvJsYDrFzqG1hoEKUtgRql7jggMJhBpsAmqh7cbLhiWDLPvvP9ZPP6nvOcgbTDP2
ruG3oIj4xDMOj8ZXrxx14Wr9Tz1uAcub8IJKKUfymqXCrB5Cdevl87Ie9gGAd7XScATC9ShmHFLK
7pkW60iz6GBBqAt913VmpJv3mpvUIZzhObuFiCGphlasB19jAOpcRkQRRFlEkvVFMXPmmimn0dHe
HcMPy9Ts1+Yor8uPDIrO7f0TXz75PxdQoigti3zq0CVXPh4ABPMesxxK44KrF8KCqdTUenaqJayp
ktUIPKGVCecEqsegj4qYV1yPgHKAG8RpWQrcoqvF8Es2tHP1HQs1xIQORIAS4WAwaNJ5CWOmhGuz
a6tw0PvBt69whhlOYjX3X/4lChDaFFqdafyOpttnelav/P19plC/MEBNysHyV8DhOiprMO1YpRI7
gxNsUgPCbOGi5UrG6WtNYJz0E1iOBj01o8cjKNd6ZhZXMwnmSPXYv67eROgYX1Nbdv58+eYvDvoC
d82ZesGr8CB51Aqx7lhdh10AKmboJ1C9xLy2LK6iEdWMqvwkLkvtQDiLAFkrZ3RVGV5AShrGNC1U
tjjq3QZ2rqWoYrSxNOpLZlacFYbuR0qjzO0Bb95qgx3r0LGJr2ZA6cwGxbKB7bcdlk4ffDYEayBt
SuvLHbzNcG7XpGKwXYun9OK99lxftBAiwNPQzIxImZbQMn/j0dcKAgs13gqSs9VMBngfWaQPC69t
ggYKNY87U3mW5bggZ7n4dlqsNfDHM4AqJL0gTHLrDmf6K9WJPOpJO+fBIKhJsQ7g21DSOjLqZEvO
q88toLSN68P8sF/3eH6a0i9XnhCDhPrcB9uU+YWHPmE+sZmPwbXX3mldMzXdp9sA2SqIG5u3lnb2
X4hZ5Rg9yY1sRyTVLrH+2s7lOtIHK5tzHJ/9yzsmS1LPwDUMD8GGds5JGwPNDcVLeikYOMSfU7ko
rgfkHqszRSvDlgyaEbl2gDi8yY+ED82MLOGJ2RdQR8WZ1Bo4/i+CJ3TFtID6xhfoW7vabvOZX0/N
LgMc+hhNPLph3MqWwHZyw2ZVjVOmJ/UAxJbAXs4HNUxoYltRsSvk8FUNjr3pSGul7Wyah+aLFtrF
fptZN4+3zCFFfaCaPwhLREgK0VGjIawjunMNxbPehsLkNKtJZC/zhsa6HXLp3R+N9Uq79eRXmNAl
Kvzw4lGOHkygg8MQ2Hj7ALI72Zrapp60airlZWJMMQihWvyh3EX7Z85ZH8BIqF1ZB9l/e+K5I/Gy
N4B/QoyGfbVg/piGgOlPes0CzHhGlWLKy9L/a/d+JbzVCOr/2G9wBrrz1uLVhx5Ioi8Sr23YomBs
LGAzl1GzWRS2ED0PVBE38i0tOzw/acPWb4OTMxpiFotUA5BXtbE1aLmk3MHGCKHVgckVyjELqOmp
CHcbSeBcBPbzXsNnUK1cgN9yM9JvXzgn7ruVCJwtRkhB8UssQSdUuh/bjjGQSf76cct2BYLPAh1c
MX9+aHHQA5+FtJwmwCHuLhAELcG7bk6DC/xA96mPWUXSsJVsJ6pViBLjNZCv24L0L6Uq0gl6y1GJ
kUPjHJygF+WtCJ+1ZC4daz1mcEmzQK4X3IapgBJgRvRp1WukIfepaA7tsFrZqvkb12d27LTP7vFf
gJRxCTGjswnp/HE+m0eI5hjlXPYrsxjaOhlnDsFpPMeKtlwOS1bLP+4FK51J7peESf7fX76+DTbL
+Ojgg2UZO49WOJHDhvdvpMvcvbY5OO2Zn/+t1XC4E8F9jKwveJdEzIze+Wm8Y/jrX7m/12Q+Wy7t
JB/W6VGn81PPyasyCQBzk83EQTxGQN3J0DpcHqokeXJ6WHXZaRzGeaYq5WaBc+/2QFnzTpSD1nry
kRKlzOkQ2ez0cswXoBU2O1RHdAuYZBoNK4Sx5kxt5AIZbQrwJPJNUYXKvdA+TTR5IKHKhEC4voNo
hnBXRU7QxSlGhT3rFAlQXS+Mkj3c1sSgO1CCJyYV+uGGQ+dln89jgClRW077+VwsFaEk9XEMK3XF
W3pVJxMOumBiXgMEPSUDy03o2ZvLZwhSQr6jcyCIcgjkF3GUsHvCmA3Tl1/NMUdfZz2pMoHKlPoV
cupyxGWf54YbAN5lc8XI1TyXTkbovTK2JpM3nhEbfYeUloARsFH6V/E+282a82edTKtBDyf86aYu
Poq0K1OPL6uJcDxF7dFgRu1u2sweNaljfBn4gLi8UhwyOq6B91Nznxp8z3XtUTM1ZoRxokb9sFeR
u1DcyCrxX5eraQU4uQKzHPxKt0vv22CvYKj2cnb9qGlLpvTjzC7rGmo5x7n8bOhQ0qRS7sbpOR4c
EGKTo7nLobnpu+fWxZPtUw3tEusQwdK55PoddrB7AE9vwZ0UE8oDvM2CxMR1Q8gYCgPdAkBMeYPZ
SKGW7uodaTPGUwgW629nNsNnML9tmqymU4hGu7Ju/YMuT6dMz1CvWDZ6OpEshNAwuEIhE7OWFNHn
VK0nqagZdhNbnyCaIVBr1s29+MugSWCpzoY5ItH3uvEfXNbNnRMeBjnP8PwqBclHNO3Cy21cAnwV
sTtxW1JT7V5KSe96i9UPkcZqjPb+s1o4nfDMSiXRABR7OvCjSKDh8b+xVqagOWcqLWcpyPn58QJL
wpcdgc6MQMwU9/D6XZsA3NYxnk9QAL8lz9tmh+nV4oSiGdzBJS0hjkKsYadeajp+WQBy/CCL1mHe
wZTGjdAKVlmmrb6XFLcVL4g5jm8yyyffNfWoxXRbGtWGkA8swgMymsb8OFfb8W0VrGngdki1d/jH
D5lIB9wY1rWFji5JrqvjG6gf2uEpqLtu1Bf96SWa7g+mtnmfEwc34GTwvm4EBoWL0FUJBTxz0RSO
Z4TPc9jaCESMP171oz2Kp0EX6AaNJ/1DwZfxqvFgoFKIyKFTotKNR9VOa1bAsE/pKj1p3vnqSV7j
j+xO1C6aiXBVKXoSzg7IaX+ZsQnmPXI++AdusAt9ef/08ciI8bfpJTehsqu6faYYjdzxMt4vYjLG
SwS9vBvULY9F3iPPm1OjPCiWSyJssNy1FJooRb2HDrv+jcli284+pI3xpYBp7FFt3CL1Ur1swIHx
xt9tRRQC1Sf06Eh+PVCp2CHGsVa7XV6weFkGqrxfSGFu2MmOV24n6ABOcszlliAHMzdtO9yhaN4I
IhUZfhV4L7oTLrGnCyd5VTNle2/xrFtaeSTOhm5N+e2vx+6b1bLqAOWy7KfCsBxdSt2YFn3EkLFT
X4nJQv0MlZltfGYeK+5skjbF2QXUxBcNp9NPlH0/DKQqNd34bVnqx0UfPR7H/Pm2JW/hNhmY5q7g
dXH9Zyy1wr4LGbxLvoNoKlaWK7vmm7RxMXia1XiZO+c3eBOxjzTIq1NVLRHWnt+qa1koy7UQxJMd
xP5nrZceb4cU46UGyXb9KYsTrEafIC2sQRznU3CMXK/n2QFDXo+cr3Ouo/VJO2Axl+Mf+goLPE+O
D4s/RRgHwUzO0VoQpwEGbi1qi8ZQledW7SZlrIbsyM5Ko8CXB4P2NuivAhmYfizubk2aWet/iNUg
P+P9rOHuuvDkkau53DslhRV203BpEviy4w/PwLX1rQ8w2/3Lu0neoGZoI7N+Cr51qEgjOLLSmW1P
l8DzzHXLGVWvpPwH1PMhqjBrvTDRMo2v0CwGmsumrtOlRye+E/oFlAshnlwONj7yEat6Is7ibJMe
lIVoZKqclNdqlKAOsSH5GCvdJq/iDoE4uGwaeVPuuy10VPt1KxY3BZWB2BYEDmiGGxIhAHITPuth
zZPNhbMCECMB0Xbb4YeSJpj837RDq3wcx27pkmf8dPfgG0JSZouUXZkdN0RkO1DbyvucCCE/XXR7
Bm3mcWzzIdW5nSWEGk2Xl6Pjd8udfe/5rdSlC0e7BrN93ivkVTHc14MHKo3Y7NEtdVriCVf4dJVj
NZF3YP2mTCmKCdnEtzZdA0qBfHjOifldfMplGsdnHvBJUu+DAwmUzBU42pnEhJj2Lzhx0v7SOouk
aHCwTBln/I+RAbf5hw2q0qh0z/Dou2Vv/vsYUcICFtQKYg99GLH9MKC6bxcmVDKcLFjKlHuoGwYb
ajbDLtpGGEOmePiRdjofEDoFC6ju8TMzc7M5QWIIsBme/M3F4dxRg5Kj8Ru3p5afdta5R1FSFxm+
s5oLmf6tp+VJoOV32h7zhKM7nRdke+Pf0cuCrVO0TiZwS2WZmSt0BVATmejBTNVhWsJw2bjPv9cD
z34vWTlfL9dq1C2Cg6y1t5wBrDajQ6q0FNYBVYmcSXTpUXD8qA2i5n7BTq1TIxQzl+RBRhtfHTWS
BdkmJ6UWINCDkod2PeJUElKvSEeXbH5uTQQtOzkC3m1dQtJDoFTtZVZWuKeLVnrldgy2OAzpK+oT
stNf4WkIfpKC8NjITqFZCdRlRuomc10j0aJwKqLXFI7s6dAzi4F9bqAiE0qy5CL/8sEDPUpOTCMD
JrhEOYUUbzffBH+/GfoGjmNU7zoSd7hMGvjrM3KW5IYOLjKwjj1fR6uqJRbCPlu65SEvXYTsI1Fj
hT8SZOXVuXqvEWmOq6LM6Av4dRZXsau9hqyXFYyPE0i9rRVAd/QEa9qOgm3VGUPdMfgphspss4iA
aKdDa9UjqAnpmKPXxEk/2OsyRnnofHhmpN17+1Cek0Ro+Q/i9QDWiYQ/new1m6idgOT0OEjfaMfE
/pSboJn7E1ujrlK1zkLwzsDTJnUyOqFPFvtvMUuUeFdyV4G/09MxBfdXZleImGitG4yWTFtVcHEC
eeS+8Wn4Cas6395A3msjrnCI9ZdPQ4Wdf9INg8tWBqhtypt3vtumJgY8zF0pdVhsuKhGzEFgfjXI
VtpsgxKSn9qb45vIqu8JASfN9B2hwFTMvVQgzP9QPUZSOSnuRUXP6FYDl0egtiwdSKKKVbjm13CX
HMOkR5pWahrLEijDd57aPTPgN4W/e0iUwmGYNyUX4K/tnzWRKYQ2HaOzNu4bUs1fJuLp+9/PJsvy
MBf0c3X8wuLwHQw6lxqRPc3cQ7mZBUMUbFFfO+hhGo9A0Tl2t1GHbNEYmOodyCElh4Z+8dFVyyoq
10dLQvNfPi4sgtnN2xaAgQdtO1jTeILIHAo69fSAU0Spw0B0vxBCeCsv9IPme2ykHLeT9yTxAEtn
VxisQ29eeg3A7NZoNjdXDgsJ/a0vSFne+K86NZ655vboXzf6gQdgzIIii6JfxZnN6SdoUbthu/dH
9D80Nb01xWGZxCppFz6jbQ1o746KC5QLUcOxYVf0Jd6xF7E/fKO0RLB1qbh65VE3Xe0Yip85461a
Am3EsbxNRIp+zZjMfgJ0csKGEFRfY0cnrry4lXm1mhQrgZ5q/FKN5QewWPLURWqnZqFRlmR+28d1
PrNeQ+jsRRhAggVxxPBlSZfJoEuAecibMG7QYep9cMkKBoTnxeuTc0QfEj57Q8a12hEyKKD/Q/tz
HGDrGP1Y5pJql7L1oqsqwCq7qahhECk8uby6/0PEwSt5jPSzoghHh2Ehm18Z8rFDjWAGztMv8QqQ
lXm9sZcDo89tcTiG0NP8OWns4tulK6rS6Zb4OGGBS0r1NZo7FwC4Drp5SAhyjov5NB6m3t+yv5No
sg/DXgTPIJIdOZm/LgtA6gPUQqENURkWnwWVIcALzmKs5upboehgiIvI7zHGg+kgdcniim5T2yWg
1ZcD20CTNMClT3lnEN8/8sF6zhdMw1h0tTWnqmHvG+HuLy3iVw/QwO26RONERmeB/03qX4w69wqK
/6P16iYNgJb+NxR7k1/8MWCIMNcN5NXBWb8PUwf7ioxFh6rZtpWRfp+ON+RWT/1Lh3e8s2u7ylSn
4gXN69tqgEjg3bXfsizxO4kt8MNtG9ICIj7/Kt7ZKROzwK5M3AZbvCeoJKL5tLzd2jRo+WQf3Xel
eBOq77WWrE18xoPnpUZJOF56YyGNZUl84qK9eJPkqSqh+dzBajsM97Yypa9VE+vS+XI5pMvexi4c
mgr3EhcZeFF2CUt4xo8nC3gazUVirNjgVS+8+jSqszCmU/ttKpQqnu1/0bL3WdFgSjhoj3SU2x17
5WfaJU9dN8cBo9HzCNRsmIywtLlUGoWiqyoIfPxshPLDJ1QkS9Cp2hyNa5i8PFmT+DAsH9FwLuv4
fZEaXqKUUpCv8iAnc2QUy/H5HgXny0OJRRs18f5myls7r/QJDYe/dBV/BANUiRKFHJ/a/YWDG19O
p+spNDeUMHa1ddd8tQ+LxoxjYyBT2RglQ8/AhynGsC4j8I/hh/mTH9CrIY0i5xBxhW65iTvTjWwT
DxNiYPPCry2pLHZthsDr744SevSQHnvliDWm4hC0AGTifEbBq7kLqQrawjv/M/RrgdqhKPMGbr4/
AxXINkzQX1sy/jTMbmezpWOWqO2V0jMNkCa/sqkAOncqf53TRGWNtdrBZGKASIOqtT0fZIVsURmC
kxtujMJF9CfcJ+d6P6QgeEc3p/ihASrQsdsuG1PLwpYKWeql0N1htEmAxSAysVF0mTkNiKWSnIig
L5Mrexl7SAmlJxg8jmQqeumgRW2K8GZjMonEzErvl10cPX2TTqOOoBpnLcbRuQKL2y2MKhATvVQg
FInIyCD1MGkK+PNe5wXL2y27wNGQ8Sut6z/2MBB7hd3s/28Vm2vz9+cTnyGi4m2M5itx1CCc3XYV
8sR84cw1q7eqNUmUVl+ylwLPVQFAYKzLgvH07T+/ala0DbfNCv1wwryuvOuRduHoU7DHIlpX+gFS
kizwM1KXjZ/ML3ZXC9gyQUrOHxoAlXrvoHSwJDNEWbLQ82cTjdiZqrRcfT7tWu/rQU9zeT53INTp
cyCIkF1lbyrlfCJ1cIByDq680vGTNQyKFhkFDZcOJPEVnr4LQYLwhW1bwhueKnxTdnk00BjlzmcY
2cMwNgI6+/YIsKj6pnuIUPLrdniXG4jR03zBxN7IXeYV2ER3KY3zZ3wYwPvHYYRdWzrRzegeVzrs
4YirNl3ddxEk5KworCnyIkZ9vjFw2DXG5oF6fMpjfqMklqpwWZFD8iWT46LM+IFvFNtDyFwWPHgP
e8k+4aj1RIjSAHxbfVArgcNb2vFTT7ZWxJqnKNi6hnMphrWi7tOh2xVG/Jhg5Ddpb1sbcmzutI9G
CisHY3WILIZAiHPbVCeLuFJU6yFLkuKIByyXmbMQK1OfEma27ExViKNrACk7HoJSSzVrh3iyfhcH
CC3VGBjC4GkqSTN0W3yBcbpyPDuYwalu4CTg+H3hOPadfA8g24tA2S952tO4cndg/cu58n7oBKWY
KStOJJ9s5KUnbyIPp73sORgaYN7U5q2lcMuh58IxLHyfyk2HzBJJD6N3gjc/3J7iQcZrDELF/203
9o33RuEdsngasZMqrTiPVi0+7H0Iz2bK36pUN2gTInL9Gp1J5O8Tdtw/6PVrl3z+xmyWrAwQub65
so63997bgrNUQQvItY3/vjF9oLn7032ChSKEXuGVxMxQpt5sN5vfzTAicoMt3o+0GEzOJoq4D3/m
M3JA+/VU4lAGaPuuQ4isVCtPl/o2PJAODg6RjrVmyfVjyPw9R1xTlUYdlkrgwSvY3dwDKnvqBq06
Dgbx/NCMPWp3FW7FKwvspILW030qEWtP21lgAU8UdZePX+B93istdgnEhM7oR2WTzr8M3wiCBccf
MXvNYaXWHgkQlWGe0xLtPJ5pPEM+yL95Uvto07zwnM/qGrX76OByfAKC6XU1A4UYe4LUd1Sq9QDY
YbZtMMXH3yVplbcYyV4SQ4YSGdEsQSwKL9b7/2JIwx07W0DxgZl2F4tNib/j0d0F5kfZ4A+H7niB
bHRy8ueM9AkGDHpPFINzobttalFGp3cIrnFtMNufQHDUPBP/V17+SmGcFSU4WLjsvC9sOb0CxD7r
vJ8h+oNKbXir4g5rPoJVvQSNcOSuOM3gF7Kxkd+qMFtw8cItmy7aGtEq+iuIuI3jx7srDymqhMJK
VXZCebU1clczkSarUkOq24YuUtrV7SScvvbf0vlEFnykVT71mYmLAsCwUokGmt5hcQtEz02Xi5aH
scs//CG24J2d5doQTFK+iOo96ydTzipCz2RZha3yD0JnZmT2aYTpOMgRJo/5/BNlqEob/HNbM2/W
/8XKcFoeuMbP22tyE6IbcQEnNzFo2DqEekKidvzp1aHZb9I2m9cRoP2VarTcK6ziM8xDQBo8pfLG
o3VRmaHd0u608//JZFhbwG8s2cnwi+Uo3ncYIhTPdbawXQPM9Kr4/5OVKk/v3Jx6zVJ5lj52zKn6
8UMGX0zXDf/74kkwY+Q6evLMOxc07e/XfzKO47Y7BL8olOVW7gxWqwDpAbUvvhqrgXAQ1xl2qKhD
ZF20XvSdL+knbTciCmY/sM9Gasp++OUe00dQtonONsrut7pVzMRr/V5EP6HcLicRzgOdJiFVgZh2
vBtFzQzKA8oIwC7ss8KbcPhfwgzU4y8Qx8sGjrmYRcF9rD3+H6r0+7AbdvxdXZbYnBgK6tFmoM7g
cbaRDq8Z0RUTNh7xLrFNQUO4gD1gnMkwry7LOAaa8UMP8IIDP48HX20qgs9pofhBQuVs2Xg0ElZM
z3MqH9bSi3NnyYJmeLVRNiaCoy9vJ0+y6Ynn67vmBdkQMPKLT8fAWnOGn9s9G1VNi6hlO1163RsP
rH5IKcdLNniFjbMSx9bgPa55YbUBytM6cbZ0fMZZhejbJYaonLYqELkqcMvn22pLWATFAjsyXVt5
Nuts9t1ItWNrRB+cVjXhsRfz/MKtedfRbA4vHET70F8TG81tphsQQHbzAuNAe6M2CBLTuluShacI
TvykxztojK/mUB4u5cBIcgCkiCgeP3ttBGOGTdKPX8AWLH2rAoHUtKlNuxmaO0YuZCUWbQKoMLdf
YHyiHD/S6tdZV5jzmUnq5Zqd9J8/n4Kv2aU8Ml4asbZ6PAuuP5FFCRQnjbMdUO67dx+FyYpOA9v7
xE2rKM8ZVZ9Crb0+wfU3cqNSWdb6qmxzpW/mDvayGnf5/jlVmoN4oyEDo6nsN+hNWiOPwWBgYbDD
idqVNHpd6gBzH6ybd0VXS1q/LzgKsyUJwbZEXBTgYIrFBvdz/dot1rlmgiaJRv9kvuNTweXTi43v
WIcJwU4nron3JYA6cj2SWfqXmeq8gGxFENvL1t5Ux73uXIOqdBKjBGedk7XEZ7aL0/qcC5AVdbLs
lcRgnOcZWRvjj9NohzXMcFsv4Kh4bnm2siKjREsAEfyYB8pO0GXts91CN4SUS8v4AmO7GGwwqws7
KzAlv9dyouPLAJkvS9OzjI9cYbA91MJpVy+dTUnvQnMfYZfTfdKDHDxeuYOZsZVfdtFft0oa5d+q
jW9uS2ZSpWZzmJSDf5TriUMLUw34IpMijzGfUFiOZ/ToWHLDQ2EeFvY1zliuRHdmdBNwd4MSfXI9
9cYCdnAhAsFTQ1NvbSW6f8rtu2IVB6NzbMMGjQfiBD6Oi880bpcE2aRH1bbEToFoPU8ap6aRj2RK
K44q8LH+hD02rre5sov6qs8keqFTl3meoC2d6+zCLFxbUBAnuq5HeV9dvAYzRH0IQkMu5EPtk2Gr
shCsc10FKb0UmRMU8s5UlBcZJHHNETk9HcHpZIBPpsB7NVTDJWDl5FTrNKf1CjiLezidcgxbzPwh
TfA6f/dsV1e7hy2hFnOs4nop0HJw+0o3p7dqAwCsUe+Lrym/ycCjfJz3/hVJq0dd2IKZXyffPwPH
w8AEK8YrzJXFjkT8Rcau3dLXix92NpWu+jvJww5gbZgbpiw6Lc3RGIJf67R6rFCf8KgmUbnuRGmE
fB0DrPKMvvq04IBr9Tbj40vs7Ht/z8MGsE6frEvR7WxZEOcgoLfW979dhOQp5lrQ7/9xcPX7TxR/
cVQ0da8baxmT/1EzM/TwvtVIn78gm43K7SosjD+sYXXdwEIfA1L9xjiXhU//AQZmgpsF4i0dWGxL
HeG2m8XSYeLDe+5pdumXHf6zM3UWZSSZjY1VRCRvskghl1LmmK1uEvJ762es4LehY+Zko4/0Gw+W
m0ntBosyDU/gbZrBVHQMGSkZAWYc7fC0BSH/J+iPxNErWKVlpRicHh5htBvanxcV2O2BGEYCGsuF
Pe7vnGIOJ3KEKnwUOQ1nTVdeHKuoefjxkSVfomfuFvteEnkk3bwHMuv2Nl3W1t0qEbNir0cdJYMf
bEgO5xZHaL/Fv5sHqqdzOUWQPrsuMx2BflHjiyK+b0jWXC1rWX3oTyChAjstFU0rm77Hy/fnHD6u
actotQ39ZeBB+KQq5RusJrGEDIqiQdBLW5G0UqMtqMupRihSUR/OOdEbc3cHAcqbkzgbpZC7WY4w
uiwPT4L/OYGuGoXf/eGcDmssWugcNl4KEStsn7N2rlx98tkFj47CP49rIrKpE0gpo+2ZNt9k1zzn
9v1zr5EzEA+z7ZMFL8qY6juCxx9/jRLE1F3yfEjpvdYPnl5Wrn2jPKriyuUws7h+916P3aybl1xN
wF0SgxWBsgbs1bMnjOUz1+nE7xP7o2ZNqda/uOwpjAj/e6MvYo33PG3oSov95NMBGvGmE2L6L7jv
0RkNZDWoQQW6msD+MmbmPmgMxT4ewIkDdrb21gH/SlIpByWO6/MsfOwoi93E1xkM6Ix3ft+sL3i+
901fuwB4vdIYnkKQp6vx6ka+zYZ94jdo90QHQsueMDCSSTPKu7IQzCCd2FHX/dZNDbVX2EkR6x8l
N29LNnJirCFPh8fpdFxUyWhYvayIx1WMogJxEGxOtvrvUnLfhJOB7IP+kRpWHJBsusyVrujr/E/0
pfIwogG5Z3LeDuUyKW6QSGmvi1OdtA5pUZxr3Vee0kTzdrB/M7AjvQ/RdsCpIF0/IobjbwuBlUwf
GLD6cGJYD/Cb5AMX/E9RPPmzeSY0qK+rQ7RCWIkDh7yp9hCmmxxXHOHcO2ok5UTQWt8CP4ysgR0q
3naHUw7P/zlcylqiukmVMyCkQGKWItGUtC8gqeQosHqNGA9GqB/9C6bMZlY9ONWommIvEqBsUL9s
3r5gwLmPavnfNVIZxxJR42cMiWR8zW3etr/6zr/fMEFjRfXja8f0rudqJLec2bAcl52B8EJWpKTV
nbOBY3hqUkXHEJbJxxeIUlSxQehQsX+porJg977FvblsO9c3cYs98D0aNAJHYiDt/GyyDxcapDoL
xIrCzk06nEpDiCGy8bC0NtnzHkSMlebMlRQ6rTEjtKS05HahHy0vyBRA7rdHCWyqnn+kGTi0WdR7
GpO9W7OvKss6W+jpNVlsNvtxUReQtbY84EbYTnugeIwkiGfhNCvF4i3fU/enSCntD4T/PHKG7Cr1
JHfxBkZXs1gcp7QbGtsnmsCmBDuMG/9h3c+p0onx1k3SsNCZK7m/rN1KWz5pMWJ8rOvAU6GgyBhS
uBJVcvPJlpf32aRF+xmUS8R+eax5FmEA7ONm6+6UPxE1O6ueAZ0E202ECsu3yoVSJx00XRK3c2zM
LGCIGlHE2NHGSVR0PLKsX2AC6ccKNayzLi1+gp49er2JD4HAOP/qZdzvKki3w82pU1NIAsUZx8HF
XfQEYfnpwbtkCM5NKbpFsMuhV8DuCowvHhLEnPb8C1MHjwO1fLSrBpNAwogaCUepRIymvYYUSDw5
LyW8uWqYUbDYK6NIPW+hyJg2jj6oHNKbeQSAC39Ote9ZITJ26afhU1dRrWxfwfo+n469/l1N5VJf
/n2mETSTNyz1AQ35RU3roexQTu8X3O+0VNgf0ScSCSJOuqY9MHe1KSLQeFtuJrx5j0191oiGATB1
E6UgI2y8Fm1sHlhr6Zxawoj4o9Wru3k43uir7M061I+4kTE5g5hg+kCwTr/5ZXGHkovR+E/V4MZV
78ieZcdFcI+wGdZbm2VEuU/LkAlZEYD+toPxL78BTxZYRH+HCoUgydyEYSVYaZVPaKodqOFse+y3
Q9SQLqqBzRKdY2/kKeYIYHHBilywh0mQZfi8KapcpOefGXXh7Fza8ijkVTkAx2sS1PZ4SdwpuQJr
lM0Z+5KLAkr14GHgFEKItikiUsV1QfnTJ46eRdrdtUcm6X6370As3Fy2UII1JsxXbSsxNbgew+LC
IxWnz/hk8a8sA8yR48tiGV2Mp6Ln7eKYAY5BS67mxxEdgi7/Cq/tHsVPMPbO0qKtvYQ3qx3Q6vXc
GA+gvM4zsN2WfOM6MC4nsLPTPN2PswzR/pbcl//YdsSsyi0RUXEAmVpwDyLxMVtWq03rM27h2Xxd
pMZFktGd5o/4tQfROqngGQwGuwSuYZ0QgElAroo6aekgYuWSkRLi8kOfhi1CLCM1WTHU5pUj4oaG
JVnrH8e2BThAQxkTRNQQB2bVT8pe1Mc5oM0BPY4xPuBn+9P/JX76i6Gd7Zb3r3njNHL9Mh2/wCAc
ZYEr5u8vFUwh1XTppgeqlt3AyXcD7vXyv4K+/GFfNDVwA2uhc2b6obORSiAlj6nzW5nBpinmncJI
jyBiTFcSKkZvXUU3RLdzpGA5wSh23iVui43Ke+pyuVa6hv+4dbWQGPTWgpBx1eCe7pI1WiTwNEtL
VpOyAgex5yuex7YlM0xxi56mIw+wLoEfB41ing6579PoBkH35TPTYq385rBPH6oychONtSXT9FCb
nBg4YheI8iKThE7XFvTYoNt4UOi2RJ7hNJ095P7BDPWs2PqcUMoR42xBGi5cCQhyyIOQXeumEmrD
X6XyZlqj903g9jvzRbGXb3l+NcgdYr2+Q+fufLaC2Qw00F/Nt0KumcQnIDTi8a4dG3iuC5aZ/pVa
iHVVSNWCmnXRSfbaHfz+4kZRwSNVL/DEWtIWmHB2t2ySC40IcAjU6fnYSJlnbofwXOuh2Oe3nDv/
YbuxgA2VZ7M4dEAMMvNg0WaN8OcOgZ234wskZhB1+rAwQUMaI2492mybtD960bXNk69CvA+B8Aek
MlW8VRqCVABjVX9syUjsBa/BIuTVsrV1AV+obbKlBYFNO1vnKfEPPVE/3JaCQhhsSAstU/lRw9Fu
OUsucDXRT4TBZ7RS1v47xhSacONm+SlURIu2DNJqr6u9EBG/aXAhjkcukFQS8Mq6xDXfpF/bECeG
a2RQX8hyfPjoj8UMJ8++Gq6CJf6vYQiZrhz/zelZxKgsIuzJCCqAbe1JfMLMYG5MT5zVUfaBmYBA
JeVd7UW3rV4kuoAayCC+Hl3WA5B+HIEflyr/JHk1NrCGOeFbk/sR67NhXZuYSVKdtHASZsTCRfaR
o6+cLBUJ5JmO93IPPPLXXvdHKhcAXtgrjV7CXsvuDwJ5UVT6na50n0igr8ep80mIqbKxXybiFRrI
DuCLpCAlUilHuBLd/MuK+4N9ydSl2Uq0bdoL0LSa18xcHPENoWwwVGUGmvGP/FSaaTp4w1HKpod3
pDdnVJV6rJ203YufDoawdxdAyQx77tVsay1jXzFpVFkbAWFnULvsmJ8cb966Tq6lPys0sdqDOwzW
rKsgxM4bxXhT7XQSXbMrEd/ymWXdkd0mbEUUwjERdd+79ZHLF5/KeHWcSKuozy20xH7iQnuQlmTw
wd61aICKM9hReft1oRsD6IdYz2SXQ29aeJ4V1dcjYfSziAIs6C5nC1xWlE/a1Wamok6cGrMXwFfv
kAh0xozVZKmtl3NPg1NpGlo9O2EdNM+tNSf4O0CGEnTCm+Doc3rS/2U89rqoD7C2vCCVoCebR5HV
9EdgCeNfEI0GMczehiy0QIZ/6fPAJMop4ZykikSOWq6MrV7raguWbEznGTMgh/xacB2phm3WQP1Y
QsfbDPXR98peazKHZqRM6OkclI13hYH+pe5AbVxUx/f4IfHSxMlKPietkaAtNZ3YQadkbxmDYwX6
4HrjKUyYi+oaSj0YtzNO2yVdw1ldrdFBKCu7JlcB4+PNR/XiFBCiq+UAi7AYIFiH7moiS0D5f6nV
12m1H+zknrZtzs5/plbb71+/62PDXQrsrLoOckC7qKsjI9vn5sIDKxg3q5h6OnKGB0sBIFKG2ysL
CqsC4quU8J0Ws3+mdLlr1elDvT71q/+Ka4ppj7euiLNkO87pqPefj2TCnmc2jbOHyADZvpyQW+um
aRXWF0bth6drIPQD9UPgyEPgX4X7SR9UCq+uepU3pixhsT07Km/t3jsLe5XaAJAy2YheitkY/qcL
3SqFVpZN0y/iMdXJGBj82xrAdJip+AvUI9mpNirt7o3Ir/tkFHR+zGoxjZI95arKA7mYT9LVJA4b
FfawnpjyPuCGYJg2W2fqmRI48tbDM5m1u1ONQy99IRYoyb2pMZ+Ijy4uW5CBsp5GL5EWfoLIQvsF
8CMGrFtPHauPeV0x/aSjUN4PNtCjjz6UgRlNJi/6f9a3bsz9Gs4cOb7E4WwOeNS/jIpapkR2FnYy
uMdKVi2TjOLUXkHVOxipRj2OJFvgavrZLXSR5DwQf9g/cjDmHIhiCczs8AidpOGoUlOQjTx2pQ0C
nE9jrsmMnqjLirbwhNHYbJfsIQwFgx2aY79v49PckmtlA+c2IhyeMufUJvWw98YZWP+URDPiTpQG
2Cn51zEo5/+bfLBmWmsSs0R+dVZomtetv3ISTLOnq+h4KqRPC5gKIPtgREofWzR5HO20FR52Emx5
890y3Nq2LB7qmZAGxvi0V91py56xz4txbVJhAyDGJNlqDu4OxVCbgsG1FaMC6C7FwoF+z6oGjmqf
Hj3y+71w7qvM97SuVsuBPTxH1LmHmcMffg6HK5B92FAd+xrSGjwiW/rkvYCDOj5d4dJegV37cffP
8Wce7Rpqiqh1PGY93CB0cXRHV5nvYhIqYzwLOAujLGUn7EAJh8IbrW+rO3QJnkM/kx6yOJDhNwUw
YOpI+Z3X3neM40A4Ar2z/IIBIFwE8os69wXN7j8R2+9gzKL3YZLKSDjxk4hBut2sT0vwLqA/hIDj
eMF2IelA/wVtNaIUWJw/qt6b3oIslw/94nTxg3fs5Xu24/FEks913M0IR/5WwjefmaNU+iXoXTI/
9NVFLhZubyrZrenco1oqml/o5aT/rWzRUHOG6fO9wu0u2ql+m6MJc5pmq6vwoMgyXj1U3wP7kbBt
hSkyln8BKk7XZBlLLfGf4SnZHL+gy+qXDqPq7pTMTjQe5QhqADjG6FwXFD86WLXsuypsEGY3mnGI
Ugh8ufl4OkOXwygOQYdRuUGKdzaJzHiYGjLuCpS6sC++bbP01EIWxg43BPjzVvnMkRu3/htUl7hc
5tXJXWQP0YI5Wj1CiScZr0YxJcUzvX8VPOwsB2r5BN1Vzarw/eWNFNii9Cn2xK01O39KC8srkNfX
pA1Cd+xP+lVXdd7cW30OXjEKc+zgg+FOLIVb1Gy/NCezRHQZfNna2wfSmSwA4mCLkPFfmHgCggJJ
yvUsqUVVbrKRoFaPDFz6JUWHSiMcONW2zUYmi+Mmmpg7L4iLPfH8Yu6Xf8G52q30eudi03qqBOf9
efq69ols3VWL7WiHhp69GIUC6x+hYo8b5z4unEo/DSl3cOLrDpRafHXfP+Q7uI/zILGzy06AgGzo
QemXssI/zY0x2tkfaOHejtw/MTjRUQPr9ef620wEQNiLl79cPVsnLaU3vb89fX6+LqN93/L8AGPt
ZnukiF3HWluvmwviVypLvDj6CM6LCkGVfBXwBUpN14c6w/T3m8gegSdHcVaKkVw6Mu9T3K4BRY7c
oiDBY4wKBTR6lQGGi+Wsz2mJ9z7hsx8kYNVqCHY2PBItcKxwKoR4sSqoCcV1Too1JcI82bmsNrpF
WwdzcVit8Nk6n+71ASi2yCuSD6RReshH3QpH/ZNC422g5h85uiEpRBzw2QKiVz8IXepfnsYa2PN2
H0bts+vtFt/jhlFnlXGQy+PeNK0JMgzjwAXuOzPCx2cQvqnWy1FEct0ZUV8DDvigPg5zr29ZxoPU
pXASjD7pAWcoZubQ0UB1L0yb0w1tMD+L2uL827MePvlIcaEtyHz6Z1FjcL5Rj5Yfk76EJdSgMKqg
Rb8KuunUUR3g9rV8F21wBE0mUC/ZZGkom2ycRqN4+AgRF8IimW43yTxuEKoTeG+v4NW48SQE+5T4
/I9puPQgnVUsduSeYfRGr7Itbhkb+FWEL9FiuEK9INFsJHMj1cwe3Lo/ZxDcCOp5vnrfynTxicq/
GwjFDoqrdGMz/+pZUEjIXtv0NLD/+Dub7KNGgkI6MGMkeUK2ZcIrEBre8L4GASdmEbUoVldRKqGC
U0n6pm67Ru0yrF6pxvaPVxMyMCGjyInpARv/s09W55uuOJrf0urWO9R4Tj2KrM9J89CL0u5nJ2kT
jrDX/v4U7u+FnSYWpIS6AGuncCaTgxr3KS5Xo9uZpjJ9DnyieqK2ACyOSMkHHc0R8WnozCewHatS
Z8TehNzqB0aS1XV+CMi1HSS+8DXkZz8KRS7jMDrJzEaBfyRC6XL0a+WecUJr+eClFAMwbpbPyZvY
4AUQj6zrQibca6dMo2k88VrRnhRRmhEdyffkd0a88gDXBrOUFp8ihOYwR4cRaXGV0bYc6r05U43y
cDwYLJwQI2XYyOm+OWXJdilRHAj+/KcWgOZl20CI/IO3ia8n5zmIJEIU2FTaWSjNiBSHRUGQrFzR
XxTbHNIZGy7YtteNFrVMdDA2TUsooV3+sul1IYuUO1NACX176TYzCf0spK974mFIFj60/I7YPkPx
k8Ub6pSErUMqkk2FkSY4vDQqfvayXOLaanxTuQBZ+dcst6FrcW/PQqotUhGUFotE+1UhDOGTmeTe
tS+ee8P0cxynXUO5WCgBaeq3YUsgTyPnoXT1/T8FQ4bazZv4ihMvw7NXbWtYTFw6/Oz5oXOSeptB
TM3i8aQb6WiG69QuKj/qrjhfyW+d/R0201vvn6qJOomOpe4Ow/zVXdHXDCtUFj+o7iIFrc6dZbNp
eiVkCrAE94sVuWJA6TEPTPb53jYudZTzB26ZonpqDZlvplqdNmqlSfXay+/43+aycuKI1Zl/yx+a
cNw9PM8jUyVEMZcilz9GPhVkmCNVTbj6Sdof+ksNnxzS6LZusC3LqF2WIpTmTT5XTUC+eUYz0MIc
FwI5oYdNXZSQuSZoSz43VlkQJNOSYkW9Tea/cQi/AWrTkn1NF85W52petAJiOZWqnr9AWBddVR1B
ikBBp+AE3rTzF7aahp426cOeW+PMxZxGoNzFEa+OLpyoR5MEi061sTKmVq20/ApxhI6Do43smqzL
PgSgjmNOgH477Lrz06lUutyO1VM120CRCzkY0nYOqzR5g9n9Ihl/aNTP7ZTH5iKsZYhSpM0x2WoA
4X4MdjD7DOYB53/6E48kwmmixoxj8Q75worMFerrQkvo4fQ4LMCSc5IMQUwrEmeT8ipeTeFN2hol
ChLhvAlgoyOSCCRXMaRAfLa/cVAgq6zUfqltipwB8Xu956mfa4uGMgZsjK8F3Tz0WaOOrgGusXTM
zuPZD7bc1ylOQCzZlKgQHetuDQEUCcscBetg8VyKe+TLQRFOlCmkOIxqfnsP/D1LZHQpIeW+SKMu
WOy8K4+O5CDpS8cu1hbPNUufDIMNNPBsiNz56tBsJsBqnEEsu4+vWmB4BN0St1uw0gXY/1rBp+qM
Qv26RClQg3gld0SFY3U3uFa7XFWB5LkeHQVWS/Qrm9Y0Cx0r67lRmH0vpX4qWsHdezPBi/eyEQ/g
T4fU1OJ+nOcxtkoFXT6DEiERrmgcH5EAz5Frev1DgbE1pUqDC//dYeEKcUu64zjk7B+bYjHoCJ17
Vn9gYMMFCUvZ2UkMhA9dJHtm3rE0JzWh5IcyPLHzCLX7JOekvw/XwSM7R2Xdwdh0thc0MDdysjv6
xcy5UVGNI7Qca+iLGJ7py0Rsle1BTk7LiYQ/vvDT/yjMUh3dG0/Vhf/0iqlO/0Atr4ALfTf4Rz+D
qlEz631jnOc7sYUnkv21ak37MJ7zn2XsB9xqauqh8HeYaZEfCpbXQE6K7LM+wioHy5duOkmlBuR5
X+r+Bs2CsP8DfWScPGWr7ZzjK4GxYCBqFY7vTA9sLOG4MfiCbhaYEdeoqpb+9NyVmSk07EGVrWo9
YI6kxPdnFUKNyAFCedhy50sb50799nFFvn06ZroyxIxPxpokmTlIVE58RXUfrHku6o9FemvPxtAQ
taBAHj31h4F/2NmlwifhEXnD/2iBCaMcUFjz95mnS+z0uoQQ/rX45EFouZYjGPA6ciSmd7FYsoWm
8gp3rFXb9/WnQN4tj60MwCOJ46UsgjnGUAqaIlCajtdq6oWee2CwjNQIfW5Tc/rha1uJsGx0EQEw
lm0Alo8CoN85NdsLk91N+00w3aI8WUCkbk/DW1o3q6+Lbj37LwvKmy+uwe4nQUldzHKqULrtTQFp
g65VYOrT27phe+zppB6kA357VPZXIb5fvIvT1qQ6m+S3rb64qO2GhdM6hNTctqiTIx4yazAW5pCb
dp3fRh+WPc05vsZqZXpb/UieYO/9GXCQOLz8aJdgByx0UZnfRtaG6AyT6cdHH6U4CCcSaDQqXPgY
QSTqGCjHn9K1sxLSCjaSMdop64vrXrO1FPY7kKjDvml18Ue+CMD87Jdy7kILVT5oJxS/19icKM0t
4W4qh1eNzw336CDAcPRWNkfEUGSdL//J4RMprptLxsJs+U5Qv1aBqDllOv968guiSptlvIDK0zIf
dAtoqdN2Kro274CAWdyeHQR4erdwYfM4QdkxiZCpWFzKa0VYXlbih8SLK6TIW7F/LXx4qOS41kNu
t0ZL4YSOKBFKA5zqx4AFwMeMf8J++lpkA/Yl2DQufX60h0uzRkC5QYfzf+770Qtha89KTUdxRC1z
AolATDNppXHlkP+ka/sH1BgVKZfZVKjFDzWFWCPXdn0JuT7l/rw4AItiTCkOtbn//jxVKFlesFJ4
gXPPsV0Dy/B9lTK2+7ky5UY4GrvJbIOnCrfafPnv5p45hZQSTg3J7w59qPGPaghm1NNwCKxVIuIi
52lgDrCFqE0fScJITWi568LQt/lH1s3ZUCpJJxnpV/k7v5IP6LM7+jsBlY7Sc3wV8jbAq42xA1ys
/g9in1AVCibQNgbald5kBrsBARD2CQq4IDRbueTD7qpw3bupH765VJXV9NQrxACSthCHThTvMEbl
SvTm5iI65WZVXy6L3vEMO9dg2+OfuCvFP6UIW/Lb+bK1c1q+egwy6GdNks10l8gsLMatRlVn2Y+J
Y6HRrU+aDJMunVqpJThun7wTTu7ayoqLuUspgZ3ZxJyN4P6c2kQqEmlBdGS4ygc7QZhrR0bTYSG1
phTSAKf0Q9BHII4ZWDbPNwPGZurDVQb5q35p1vM7JvruAmw2nCDgR5X/8VLFHctjKg3U542XVBcX
ilbp1WCzUcVv7Bz9VbxOy/NVN1x3oKI15LYwkRU0VBKBuXZUWJbPmGukMwSt+jbcIo0hsu/GK0yq
WEGopjvPv58CHEjmkca66B31W3zSD8pdWt5SqT8w+ikdYKZbmXIhoyAjK+c3Dq6ES5tmRLB6Xz4H
vHvfTMbC+yOjzziYPS0zSbOXX8YKgIGyXrBv7XnzVcZuogv92RJh5uSo6rXqYNQmS7xORksYNMpW
Ib7jeLARfiITEYDOWexv4IwQdxhHzED4s5OXMijw1+w31JvIBysjPm47cw8SRlvuhXxqmqpyKv4K
7kgiWR6xSr5WTfBBCtV1PDqBmU1UI74YgB17X9xoGnrNIGEBPmXFd5nijItuhKp9bRmUKhWjEywJ
wX97AOLyrRKHqTzb3HkCHY7pp+AfB3+2bMfacuQd8tUHnOiroR1UAfcuIeP30UenPOnkoO2pTeVe
JBgQN+mnSA1TMWdZ4LK7D8xMcl9sVySL4qkA7T/fiLDrF0uA3T9+Ufj3L8mv2I6Z6N9qr4aQnnLY
dwBEPBp2EGgvDHnfx5he2BG7zH9mqAZFjZMTxZyHCHuKEX0odZGUoiS9FK1FUoAzFIlyO+oWCbyY
Sqm/q+6GIeE6Zh7BkKNsKoikhrxGhMhWbyVqBqG4JMQr/vcnahL/obTRCCxU1lXxHCA7LFnwEs/k
2r7vcaK9TOj/DOXmWqaGxgpTwcbQmrKIBLG1m0tFhGuPvKkimyErdlcF9qKQf6c9t6R2RYDdNynt
NpirIAHyPD+pERzhAlRaiMRtZr6X1sqlXdFLxwaeEA39QFiIwbtbuhRMpKvilAyzzWW/ZTP/DH88
Th5+P0fM9fNEZSGGLuRobnQXcArDvvR6SAvmsrx1eIyEbaw9FRFmKiNyP7+K/RPq4N50mPWuHFVi
qswWwjDGmF1OC1xW1QB9mmj9BIlrk+/l793uqbYpx1mUr3YKtrljmnOh7LmaQNEhXjL9inDWIMAp
pIvqTvdUO70zLnf3Y8OslFAI/Hrfht9+45wMQwkxW8jgvMgvrl9bfw1I9Q1Gs8JlSrYmsYkfBBHS
ayJCR9hlTAbEnh0uE3zSV+X84DRTnxzxPHcby3K9AzbRl4XawGRvxBD65UvjUmdTrxg+x2elAeHc
/nYL6aRrHzsr943GYwTaXPNvz59qvLu7afSrynQDJqQ4e8io7T1TwUnOdIjPWYcS8O0q+isjCly/
Ost4rFGfOGj4m3nRtzRa4jLTyM1adA2JJ1p1RzyEC23bQSrJop0L3wijpO1gO+0ds+nd1L3jD3T4
cP+EBjhqu+o8CeNL25nKeIhecq7KpqH70W+LqtVVLqRgomxYmIAjb9VY1JJU6oq/6F2fpegBnYKE
FlbodjUERdEmGdU2b0258XA54fN+bmQuoTsXP40/0NMfLHWy/2HKnqatYHFRBidlCwCGsYUz2GNI
HnhkuIdfHg03nLcqL2mb6uzbJKvL1Ntav7eG+dtqZFuiTyT1zpTVSnf8GGEkErTJKcblyoNiRFDV
xV7SV/prBWCXJ7UyO8dG5RfEQJbbM087j6Jp19cZzF42WgANSeCNEyXqBHh6xcZIKBAFJl64rr6n
9PIWpxwgaxlI3yXnmEKq4cZySjy7piDJYyM4qEtRTUNfzxNNBhLoTqbBLau699bmL3drExw8BPXP
bBDxnTVL2Z2j2lU/GoVxtype8bAeum6peHCx2lQzz3Bq89uprXv1Ss2pT9vDEXWlfnbqMrP28Ot+
ykm4LzjKEWEQg3y+eVFVDDiYT0sZHmxov4r0ouFUDNoHMPoZfSADTQZ0bitnbHRH+EtwXyuxEGl1
Bt8LUot9wFrm46t6FmwWuZxJ6n82SnrWefFAhseMV8a+NnqMwJ5IMru63HgPGGDgFkrBURK2bwmb
ZLr/vl3WAXQQQkaClRcmHrWJsv3jmx4PC0KySdH8ygcXYEQ1dWghzSQqKbA+c1x3VHVAomNDtOG4
zhufLslWEr6obOVj3v7N/1d8z/beSOBk1yDZycvQNTyoi0Fp5xoiQbUY31+05EGosmG+p6KTMzHv
+goMZpbIifyjObfAP5usFUwcPDyRsfwHjetKMKRmuzylKGc0efPqrEVI3p82al5/tRqDfTG/ZanN
8GCRmj9NezoHsHwp20ceGS+vWqv7egzp2D7X3yrKWcOREl3/qViPXv8B1faBt0+2xCCKHU+W5jhE
HQbcZp+UrOGGZCZPlVwfNkKNrQ2SZZKfJQPlJzJC+BMY/9lSto6dEjftJasPi7Iv4sA9XH4nStSM
WHzl3q7FR523KSovppJuc0+MfkQGj2mCEf8a2PquH8CaSUAvfaF9ePPcs8mWLgbo9ARZRV9+m9Fs
d4iLiakdVQGqqoBcSaLaW7nxBaMJ7hT4Aw74r/u8xGLHSiJ3ytxJO7POWHVOGxAPjYu9qjSNnsar
Rx5vCGqXn9SbjnIsYmJzlNe7VgsKWgqhNLvQzgEFjVsajme8Oopc4hTcAki/yQD2aoNnu7/cg/CS
RQbWzctQ2RLHbKrLmWbsJ5oIvywnZ80CBVW7rbq0D+CT9AN7DUTmVSoo4fi/79avwbTASc30WJ/f
t3IbaMMKWONq215otYY5/GfY9o2NKU9iSsiIQpjCztt4J66FFGHdI4IKV0vuDhRI+LqOc4d1L0Zi
PzzwDKRD4ehr0XvyxLQjnpUBabISUethXWOLOwyqv8YnipZ175IaNKvrHNALa1SdxWb0nswrPUs3
dGWa6Yoooz/iqio9aglBoAUQGG8lt6D16JrPym+h8PSwl1uvQxcYHC4GTpiyltNjT2NPKpfarV8b
yscetlgOfGmHmZ1xmRWXtsaeQ1ivZf7OXnRHixGUB8/z+qCDUH67JIBTAGW6zzLF46A5Cv09Eg4q
4oc9V02zIfhLQJKG/FrKpJjHfLLv7SSDzX6od8DnK1MjRWE9ynNGsdjCvGdyQsY0dz8jUuRyGqxC
uFD1hZ4LRPM6Mz6Wmt8pAmGAFJSNi5ZqmaVK3wnIMppP0hWiO2ycrwc4zUfHUtZFKvzB9aTiOyBV
KezmhGFEOKot/JSkS/0NVF9jiq8nsQL1giqSdivgS+uQTCS3SL5ixuPFVI8yM5/JMEcyMh1GteT4
TacOzlraEOFMt1XrYeX0rjxCzoYlL9Jn5TivgMHrqhOb/10+ANEQW+TO6hco+Xm15cQSZh8uSxTX
Ppca8INaPJHO4oab/toeukCuyh4Lu6Xa7Vqd6ttgpw7JIY4syVDjOwFTtwDuKsapCq5820L0VpN0
0v+k9HzIoJdUNOU3XCQULOY5c0spYc8WiRwJNV8BmU8AMGi/s5Y+yQWCZ6JO2CBKmO+QHvzh27/i
rhICmDPOIG2DIlRFKZ8Q9ROqN0ojUmBwgW5kWFQ7/CFZDzmekTk1v2GE9I4HHP2znCC3oBLX0qeg
tIpG62xGlQwo4p5AZsHauB1YhWQfnOftvlgrqjhluisWdWLKQU8MwoBaBkHyzYFU0rJdVRXTIAp1
FK4h2L4ltH6QmsWk6rHh/gYdPXfv2VtMDUSsyKCzk5V+eY1fB4J2n8G27VB4saGpN6PFWk0EcM8a
vKc1JoPeye0oM8zbQ2SoYT2+hAwJ65tWlkjB4OtRBooXHJNLkkDjT1TAKvKiob2GToAyMHaQXYD5
sOpniunAvRBr3apg/fHTd2eI7hZ42NnI8OolwyRViI9ABb1yCSfPi+31pFlLq1a/oBThHmXqkXsg
nkVa8N5gcfGTFG48KJf4Ex9M5wU3zin7TI6INFDA9rUNyieAqJYnfdlpGaTK2mVr1YRKf8rJ8pI8
HAhvRAEFDHAKLHE6wIv4JBJ1tNkIKeTrZdGcGjMzVb9/SN5Egabw0zlbr7zI9Au2df+6rmMhzffW
0H2cKV9/VF9BBPLey4AB3ZYALFS+du9Xm+nE1DUggmKnYKMu41/B4KsKHoVn4/66vMjIX4Jx/09e
N9ibG/9nOsZLEBIOHXtRBUBey9/ZN4MyS09Kwo9oRl2KshlVGWLQHWlpk4LHVAnwYNsl4OZTi8Gq
EZzMPUUvRsn6JMV13O1+5BKtB8wUre2otZOIg6TGPsBqLMOherB/Z7KllSTWju16uxQY+Sy3o90v
80OQEa4quE2QDvvQSPha3bBY3zQWAy4QaiO8lijARhuAiWq4GUe5urvlSvEd8GlZgkZmSIiqBb6R
T5DsTBpK4Bo9VuTOXb41yN2Bjl/k86CUTVLvue80gHy7/TVrsVK11PpD5nZ/jFshoCrf9BXW1fRM
TcCiVL3F087yhPu449tXla2zNx+GEw13/yWJET9rNy962ndnR8/JLNLM60gHHGum5l9RBcsjPyWV
cAJwaoWmpQz0QMUS1z0YJfEyocULFrdOiYmx0RL0q3LM44qtJCrw+ayCcrt99nyBKHGSXPZW/HOD
pZml/a2aMYA5ffneXTO0ZrUb/hf4tr9PbFS+AErAUXmgTeTw/bdDZb5uQl7vHW7qz4OhNZhF4uJv
MMIGRprg41Lpvi750ErxTnwLyT1NjCcwZEsv911fuwD1jkXURUiHIcJgDNtZKg6Czj+ipTX5qOEQ
PJSayDB4TRRjhxymNmhhXOnBPj0ckXXK8ocrTq6wQeV0TI/vqkPzsQBsZa5fgdYCz2XedpPZWzpa
JWZZyH+bBs4Gy90ZB5LqNdnF4/v9wWO/W24qE+aLJSfGzqUruWTTMe/EXBgM3myCWasYEoKW5Gy8
FwOvXh1oIVzGJRMJYWAJ+g3jbOoTlK7Pj1jN0ijz3nstmMtfg3MmKqIPSmH433zWhqEI2mIsQzT8
H++0pqXnXutEEgAPRayCMcofy1l/GnSeyXwf6ELynn2jRfuKpTO0JALJDKGLEc11to/BZ0ajlEQy
nhKU93FCmT+uBVEDiNQ3JMp5Nh3o5QrZ4tU4ALZzZotO+NEaN/8S3PFH4W9cZtQYstelfA3Ykugz
ijJ96cn26LG6zhNmQ9y3qsT9r3nrbrcZgZkKIaV8WlWmvjd0W4jkFVwJZEZbt7kccAJ6QOyNoZei
7DlATjh/WXEv7Nt7xpZxAEGJchygOw2FljvxyBMjW5jNR1Mi56jJPIX9InidQu2mSRS80we9hKyG
lbJd20+6coYYRB83bB+Lbg97qhM/kXEsbOReJLbg5gV22J1eZ6HDp42KKiDL8AObvtAPSt9uPPpb
tEYAuoivklQoSCrUfnlelxU4H240b4o3rkar1cs5E2Wp+h/rogB0k3UsX5dhdTFFIW4kWDJszqKo
AyiJj0jenXegXk4mzW5j7uC8eIhTdc+4y1Obnl1i8ZZDse2FBZXTtR/CnQ0W5a5IXJEQ3G0f+Ghh
Wy42mtNxxKkxuKYFuw8pfBsI8ry/dK6x+sUWYUf/ZcrIjowtRKww9VaCedjuDDWIUEqdkRIxLKsG
xuABBYNjEdgCSV6s9MT02c1FOrTnvTkEDsZNfrlgn0pOYjmPTFmlUztGglc9leiuXHyNcc9qrXzt
UgsMPHXCP9s9KEvmzD3P0pGRYFWfg6+vI+BZXq1LC3Q/oJ4x56bqlUIFJf5O5SAHYBHe1hdu2b8u
YiylmSiPNGUPgXDSI2rBWgNv4MhZVFTgPlu0oEmzjs81oe5q3TPrE2QZzDqgrm/TewazPq+9YYcK
poG74cvr32fOlZzynavtbnG1vif2SDVxu/TI6wvW31siKsN/8y4LBS1+MTvB3hLE3pP2qDdN6NgR
ANi2knUDdJVKL3LdTwDF6Cj7Efe1SjdFa+8eXNpKAzzcJSJ1WFRp1TmHOkhzr6pmOWHAC3tWpfYl
J9NEXTHuQjY/9zJgn16NEDzw4t52VM3pESa4MLQK7EYKPuTYh3cN4i8v2ec5uxzvvlbFYSBiBLD2
M6rCJ6b1eKhcWs0SqezeAEul4Q6eHvo7iWPQfKJXn651H2zBspXg19baT7Ok8ioN6vQrqfjMMKdP
Ra16p5JHyoj12ysVc8hSB7cqnmxlR/xEWVWBq7tFXuYfJ2z5dm85rLbJYfJjzayP532W94JvvjRz
MxMRfetQEiRp07mXLHiD1WjO8ICOphx/MZyFQYbCaiJDlwTGHz5mRmzu2XRFtGqo/DsBVRuDL3YB
rwySfXIiz1EggLKYFfeSSfKOR8ktl819QL7byh7YJVYuhKeEb/DQGjucAGHbbjGv04z6AW1GJ/ax
JJ4no21EXJ8eJd8LUq8UBWATyar2WD14DIMSxeGNLtUgJ290Rolhq05SHQtnT45ksPzgO8KDetBi
ViiBtCnhz/Gfq4qeIujuVucdqbt5uWUjmDFOqc7Ho4kfUJ5Ow4HzfQHH51F5KOkWCxrH9j2WmT+q
NUi9LPbfNV9Yn1lypPtdUxiAMGgi7vl4zm8Cc21j7di1V1kq0yStAS29fNKOiMLf3Mcj4qOovjwc
4DfxP9BBzQLOjwkr3b5dGLTJplr90taQ1fXeFJzB+Mc/cfgZ3+al5/39ANmt69Maz0O4rA45rSPw
BLbG8IIfarv4MftYXpHPXpi2dkg1gv0UefLlE53YN/osymXcTqWn0fDfjOzRAX1x5J0nFvtOS9yP
lbcrvf308vSLH84Z1if0e5gVHpIaamx03VQKEdLBBF8JqseudfRxWrmy/Dvy4cLbvZU4mp/n6bCu
3vpHAsVFOTTQrZEjVbW+BN1nLIHzyo39jMVsk9wha8YzeGTSlKsJ38HxKtkT314j5LSloJIX82CM
pLNxXiR7nXRGTem1hATGP3mGC9Pd/NG0wHDRHGtnqLAZZ/q3iel3DQzet65SBn2FFygsEAhQBYfV
xTULX6XNbqPGC9nR4qTUHc9Y6fOqt18PwbX2dLPaES1sXinZf/UQ64XGPhVZMmuzOlKha4GAP8Ve
qN7IqD68Y4Jglkr91Nf8NmtvGqbz5MuWa5jOeebD5Qrqi6cHy6EZWaAFx6BX2cbdP8lhug1JjxMF
qDClilzytDn3JLXW12d39zPlITQXG4fVGIKIy9n5ZkWXhCYPFft+IegU6zQsL3JghwXut3OT+5It
bBZelb1bYmN5nLfLTtgLG5Y0K2N/R6C6SH3+Ap/2Q9LYUlpD8xy/uCC+WeQHQ3I4a6Pzk2++dSEC
xY5bfFUzjr5HFyzk1k0YJXMBb6nr1aCxGMR4miTjinzpjZKdbXZWykHbdBb/D8mDCZAIjvGDSnrx
kd0DEhNFoSDXHjq8r+rNLtQmCo7eCyAZzoai8uPfZGXba5sWdoB2EmJFOcsvDChXfQ3G6xMBABIk
5nzvNt/rLVgLW1PokUYAK4jPo3Vk+lZQjkJFDhZcG7HB9ym5l0EZ/JfbMZe1d/qT5sL83aKLB+Rk
lRJZiZj2Mz+pWDu8q7B0SdIVlNvDOOAweGBYQlit5g+jAwksy+732VBCUIHcTsAgyBx0fQzVI885
7uEXNHYt8rj1CJLgvkSkviYeYzbta1jMwIdVwseXnGe7Z6OCLkVnvnYwbDIHsB8BBnvwno0AwGCj
FmBCiyM5+jn8mxw/qsFgDRqt7wmJ33cBzIpoIeMlNn0j4hx7GTMFxqAAAHAvfMbdAffzKIH8YGdP
Iqj+wFKl4liSsfm9LSVNap7QzIKVYeAPkd4aFTG7Ddyjn0UDDsEmxcNdoDThTL4FkxhgZnVG4pSc
yRmjvOnghTeCWxr3nk0EvXnDxaYgO9ujKKm8q/TLSI024gqaJ1Qzv4DrrOBMNUfo1fXrMUj5Df5r
s46qA2KPlgdYn9Xcv/vqSZMamJIVzAEbPI6ch/3OMlhRx1KxxiSRWamnE9IIZ6QxVDyRgxiIn719
RYUXcGLwrIUkip/D5PK4lWymvU6fcJ2jAfzPVyX1ODqUW+8MwP1GIQJq43miJihxcFDSG3+RiG45
SUYgJURj0Y+YZIjUwrsmfTXHcNh8IpCV3e6RhL+/j5I4SGArX0OywutRdo3Q8v995zZeXVjnac+q
BRykL13t5Sx2E6RH2VLvp1IjkkSnbEQF5RaiuWJaUvWl6Jox1YNIg1C5HGQZ6dE0qbGm87lki3o1
O8sBYwWJHz9UEd9eGIS83YW4MhneQgOMuVXZf1QByT/GdFSK5PyPHj36BUwc3Mwcxgq0ging70RJ
2cCdb2nCNNBdHgj64/u6/44oYDifVvb96PgWwImCe2V8Pdlbq567VJMwcHJpMYFC57I/AfPibHGn
EbbA86uyuQqAPbHzUpYo6jIvRtklnUPNKli7LkYqb4+3Uacr0eeh6s/qgd1oOlk7AGeLyMxGUFID
jFMMAcRhwmXpMVCQBYOjyRxGjw6EmlL5CoxZMsvVXX/FEJj+XsM4dpBWDzAQkaPM2MzK1LzilXoL
yup/UuLJK8g/21bOg0iGUPEYW0Au6DEfwZ6UaCbmXkCvgseJpCbFXMNpfsppzpuO+po4UKLevS9l
LmyaKT9xcTbXcc1mRBNKlOJfEohmin3Q5gxnn8ZWSogP5iDfJ0OuH1uLkjb6OqGAYm1VS7+4Oa2c
qczNIoU/Ql0WZFbdOlNPZfCxo7WbqJ6VYeEXc8kMiuzFDD8+aWkvBzuOwSFc3qXPmlGhr91HMjqo
QIbjCgvQnC+5l2JUuJM0jZYHywld+sJ2fcv+1UBj4wQD1IdsYJ+hN8u/LbYeClymgEAPDjyGbxDE
7eDjIrnCU+v5tutr9ae6F6cOUdSuwMi6DrZEMu3zM02A2PfiLYKAM4jnNKEY1y5p74bQCj0MAKx9
hAzec0d1DbnjcP0+2zOU3Cz+dbhiMOBEZ4t09xoEDU4BpI6cpNjQEq36bSW/49E+AcUcB3CdBb7K
e+TyrBmN0WMmjwtqHRJSGoSG4muC7iQLD/tikvCTdFfMOgXFJvoxEzi5NzGdvARoGdmrYSs7rxWs
pc1htQI6lWFxZtxjr7CSHiavpAjYUzRgAl1R9Z5w4YZgU6cDGvhSGeYfgLnOdwXJOEqoKlazCoVJ
toKC99SwyYYj6nHd9eCettmgOuFf/8MouzjAa2v0t1bilPMyRG7F5l5HGxr6MXS7iJyNr8nudzsn
Y1ANKzPBPPxzGT4K6/1OveAItUozDBeOjNEQDvWV+lN2rEJs205nKxpvDfmZ85UDyVr4Zn9OrM4y
xRMHD44yXKoF7NHYEONou1NH0woXKKqTRUAUrSTKdg7F+NPcsZUWWw7U247UlTsykS7tqHDGT6hP
v0K/KH/9XZREF8iZqIhcVYdrB2EuDUbhbqbxhNsVaTf0MbyzKsSLNi08THVSz88NE+Ip/igrMsUj
l9JNPUbBkeCb5ATAfml//c9Ep7EsQgYXbEWiHrP6kFpQa+BqbauNKgA0SbO6JnZA3vh+tGVaLQup
TUP4LryhOZlpmR7/GDzfD48o1+wQMdjU9t1VIWxGvUOujYTiqCiHAhkHEDx+HP/mIyfqm2eiB+H7
3eDKHwBVXwjxSuQWjhsuyRj2tdsz2aIvahd4L0k/UduLR7LpnU9kKFtjZTB2giAy3CHkhTGCu3F4
aWVEsAmrgiwK6KkNmfjiy7D+o85lEnzgqLh4BwB5GcatU0gaKff7FoMsOwkMjtXeQcilgukw0OJp
qlhjtyq0YC6WfiO0eJK9WMZWeaQZC2+mpUnUYq6X8k657ZTMWOJJns1ZcDTcp9SQqLdVh597Xquc
1POr3L80mtgCPXRJ4NgxG8RkA0rgzJwCHx5VL34iqxDuwKXGHRYqQ658t4ZIUSkSznM0UBDt46bB
S/8mq/H8YxREt4DR9O3sLnMSDf9pELJ39HxRjXSZSv+OriVSw0AwnUqGkabX9clcwliINW25m1Wv
yvD/dYwOg36SFagekKdnMSwJIeJViBtnMOoG66gllYiFD8SXe2PHFdNrGR7kjxEsMlJsQeyd4SiT
B4zEc1w4msvnDg9SnsBTISJB/InB7tqIXhMAB2Ra49RwLKLZsE+Csm+p09mbvDpToDqE0mThWOiq
kqQvXcKU8NZx90QfM72qinS/Ywjwx2EECkyjuDo1Dwlrt0FZ9CaXSHBa5Z+zzMPfMTuaaW5KbEtF
ey6XRYacVlxfpg+r3czR0+wg7lZ+pyVMiScT8IoXuQ4bR7uEPNbF95BhL5mz98OVmmkgaBik3XiN
JQrVS1DIIlGZhvYWCf2wihtWEB2JBitvH5CjmKvmj5IH7fANL4kJm7F5MzYJoiRV7JiMCyKddpwH
guZgic22sMTMQTmPFq6DK7KZMstM3d1b4EVCNX3O+v8hwrTe3582pdbd4prNYth3s62+4wOlBk1u
gVPHw5B4AUCsBB3T864JsBqeRjkQS1Wvq5AD3HAz9xTYCwRSR+hM4ERtJswj6pxGlyWEchh2DNwQ
BpRX2c6uu33cKwQHHWEzTJMX78qftkQyIfZXutrdWtac8tBRzrtmriB5sNMhC1iWAjAFoEIBtWyy
II5fu39PD8iJAN7/jHG3JgvNvQSJJmIeQN9TCMgss5r8D3CR5LR36QAUlvAZuzFMHRitJ0cqrJBW
h8U7hNdF8avSSEwM5eBhZMHIJBX/6AQnUzaj+LIe6kLaJiw+5Y9R8otVVUs6xJPdpSsOeCpQhIau
H7qjhFx3Y/SmW0RUN7Iva7OOtxh7++cgFnEw7zLNNFRfObGq9eNFvljrJxYONz8aUTB4lDxGnPqN
2cyskDAg46Z4YdwifVndlx26vL0ig0LhMEh7YgHDK5vnAdLPf/3jfDTICkmFjTT+8TE0uij1EvyL
MNJMCWLH/3PD9ws54wZX3uZv293xFwWVjl3mDe171/iTCDG1tecA9/5gGwgVQxX73+k6SM+6g6A3
v7A6txzDqc/gvM8XUG1gzQ6pW/aIYzQ8+fuH/Yc/e1iBuXbUip5KcVAVanh5E5t948b6+Z2OiIeN
SH5Jif7NTBQx+F4eRvIUtod1cmOzhuIICbg74dfNVofM6aqirwjEZIKfKLUCfaYnt1OffzIuuhTZ
uGUO/5ydvbfl9zTN0QszTaQxjuEFn5DYngDePlBXpGQod5bkeOGgEx3GJhgG6Uiz0YjDcSRVTXkW
sC+QmvIqC1qLszNFIG4kAtBtc79LhyDNb359uNB4ey6qEAL7Ctn6g6xyGbtrEfHhy5xvqSvPkqf6
4IiHoptd+/u2vFh0tUhvi0ENwE6bkCd1FvNsV8J66hX6yeA2+nUw71ZLw7+5TriOsDD1djgIyald
I9rdv/Uaci7MHs6YHoRcp5xAvnjbPHhGDVPhaYWlxoghygaMmQt0khyLwb8S39wJYPrEa7oTFckl
VQrUZEZyRAlS2CYlmJu0ZYU+QlCWUrIbr3MCpcBW8M/YvT8DHPmfk8/lKJz6gJc1KPEm7vcPVTpz
v/CK1OOomjrWXZx+lD8mbVxtFJ4uKm5/3qAsHCZqLvV+pVX8DXNEG4ozLGvc/fFV92GRZxSi0kv8
Hwt+/X96LGc0nEn2fNcQ+BAh7pxx3Epa/5kQ8mxe98t8IfW2YsRYgXJSaTm5qjjOnNLbIctLyA/+
CHHRdG9LLDsXwxcqpf8a/2JG/jnxrLXcmDew5dF4KSyf2m7CwOVNIbcDO3xqFrRL6NrYKW6INDMa
LxSdqh6o2dzKcmynrmvmlUIOFMNgPRNkuvyLR55iyLL8YSu7Wgsmp89yubtud1fuLP69FRhK7VCU
CU47fRvJ6CwBTRW1Ky2oGGnpQQqFkgfwHIN8bVUkkIR3JUY5s8eKYCLyBPBc0qTmlqFPILoV9kxk
WFV+r5+eXofERl9xkLvxdjSdwwdXmCYRpeQGU1p4yaK4aOsxjUI6fxf4FcNOssU3LExxzAhoJGBn
orhHuc91yUEdOG8gTDIGkfTsnmx12I51ypgKO03vd0mhpd8Qg+O7peDWO8limY0CCmcEgWHQtqDG
T1JMTyKi+o0juj1B+nZcNJ4h8f29hXNv3FhCEGDKHGs8MytRFjVNCojmf5TKwjEwGqJagEu/d41a
Jqiu5kFdSOe/fxV+VcZqg6abArIUJNOydm5vPzYnFei/g0sNVXNFKTICCMPIgDRMCS3ECk+S1vox
Wd7idJ7cc1OrKpQAamIUPA7oDspnYPZhHHGj7Rv8HTLEBlBqp4Mu4g7geDQ0SM1JmPLdDJdLwTCc
tn2oYGI6GSx1A5alDh9idFzh+XMn3yVCBsVG0c9GmiKhwwZkbxc7xB49KXQo7Hp8xmukkKQQSFa+
uyfS1RuLzm6N8ocmSw4HYeFB1fRBCMDxxIWfpQlg5Wtde9Z3jgEpjFZrOrLvQfs7p3Qkj7HhB8Hs
Qssatgxt28U9XA4gkJ4/aZ0cBPPelbcwKWRwmJAr9hXkzrwZNYR3D7fGJ0P2yowet0+OiduFtfva
t7q8f9PfUCrauaMMMIUagKu7M/K5zm2IuP/Ybb+/gwowra+l5auYuoZuygVNJ/HAQnbJeoU39T3i
PI4Db0oYL7HYBhoJb4nzNbknZqUGaLUYUvod4SvW964+6Enpv7jYm/025A0rR2/ehlVbzeRoMK0u
OQNi76VpB+qZcIBridnq91dtbrO9x9XlE26KIPqy8ZnrZKJhLSFVHlMnDBq1Z+9OHChhtBAabHwl
rXwyAHh8P0HbnXq7GQhezF4Besnu6yJjE9heXsnNA6DgWsfwUMvAI3Wv4WjW1hwhNqobp6WrcbsW
pQNuUsfk96+krEEmN6RpAbBgrOEQXb+NSnbwsUPWJ2CcQSvBbeJ6i+UDknSXG2eM7mgcVLULuy2t
os322+uKQEST4DKLklDw4c1lMj+jpqNey8Sv8f3tGU/QX7wboN7enhqoKxaVDcP94T9sOrwn9KB+
cYFqfHZ1MKlODcXsYk3dmfGIZv0DcTM8G0tXiaB5WUjv1Y0Y/pcliNdXS9G6KoCiwalNnCv2TX19
lndY+KYyRpodb3XnPrD1Q3atiDHuj3Swg3NTr6u+Dpo8V0HA79puynD4BQfb7m+nkF3njS6gj5kL
cRLgXlc0ltZEYFoUmV+KJ7X+gTLPLZQwgUuwg4iNtqMNiANA9PqOSUpWErEHV1rYaoxotBl5XSt2
VSPEqO8TaTTTK3GicfyAYxxbbPRvk6fF/sYhCseMJJ0KNKhx7hTumsnrYjgFiTRmt+WQqq4iKWcz
01xiJMbBBReB0R2CWW5+IppBz4M9ko+mMxbhTgGd8jkUxO/aHgIuf2c2mo1PPTmsDvJaCa7sN9xl
Hsskp13629JF0E2qRCehLbT/JmBmzePYgkx9f+95faaxy24oj22D8g/A63dkwzRaj1HgmufcYuhI
Zyr7v0J6mAHtnTIfmKsGGTAHswYS/D6W/kvDhrTC4Q/7HfUY/5HdJUew0A1lQwvVIL0OVT7wjYUo
BhkyOPQ205eYfGqff5aJ0c3WVRq89Xm3jVsNPXEolNGRy7BjDgjbDw+rzchXUt1IOomx6kB19jXL
4P7QL4sfyKt2lYDAA9ePqhyIPh2mAgRq5zklIVWImMDU4dwmyRTDh/H+lq0gsL1qGdwqOlBKebSW
n8PYw/yIhUCEeY+XE7C9Wx8oFmOaxI4Gyev0vRfXfRgBHirUzifhoXH8XTkUuS/Onk2xbb2DGHst
5D54D/TZcjUi07sfHbVVwvrsVqihNTRMWmpwgMr6oDswmaXOJ9aH+JLifqm6gRudbcwIG2g00OHe
4r84o7RqVdNLWA2tEhHhY0r5QWf6doZgHqZSrVSVa0jXVpK2yB7JbKnHrPI3Lai70NS9zbT7Ic6c
zlk/LupnYz9pMpI4tPRjdextlvd9HUMQX4U/tuf/vh8CGfFUstdu2GciqKuoJ9C2axJAjhE0+O7k
VjcOVM1/mn0WBf0tu6XmelG0MINIKl1qlYbcmFVVDj8Nj1IARpne+642bLvmyZbQ52rE08mtq7Zq
VhsyCAABdvmzmrEFsBlsqTPhYKzDm4BP0crH1jyJeXGTOqd/Pn3j50g8y0+XSnm0beSpB8NBL6cT
UfRUJWMS4WncosnwIUDIKCqtIsHJ4fbDC84dcSwBsWJMlvWBPK2K8wDkFOOvpBUOk95VJxY3onSC
bNM4EPCyKmX3Sri2pFgsGg4bzjIHB8k0xJKOW2/TjOKHAeUrgH1AdDYmGJRrmm6hQ+L6ESe1Dr2W
ZWMEqHxMfuUx5dpJAQHuV4vTvsIGauSV/Hl0Iz9kg6dIn+9VFVW0zeB4HIsr/EVXDLrseK+Bi3GF
IYjXNYV4aon2uQEaW9z3P6+8oMd7wbR28NJlNLNKMnzub9h5sJqZx81i74amjTB6aypfjPZmoPU7
AgOS+PNtcdW6y6HnQccDncGDsShP7bMG3K74SUL9cQugaigK2h4t+PIwrpRQqTTY2dA6MaZukfJ5
9ug/H5zmyn+Tt7JR1CmCftxyQn2aKmuca5JU+cftBF2DrWy4Xfogx8NrF0eEuHsQdo74FKq42DCp
e3X/LqszEauTokZlDV7kS/3ds3fldrgyTZB8dSuh7smt7cZ/cKi4MUkkpYQzY/gqATHQNRhwLKlv
CdmsrHqSCrrOE1tB+oRkh9wmmnGh3gklSuI7ptNgfy1aXOnAE6e5WEvhJSrv/770Oy1Gy0q+oTwU
W3CS9D/juexcfQjq44NYoyb8AaQsbqwLLmVCK2nHCnrkJIy/5seeez1UFWJ3gN1D1KBxT1gHEVrO
ZsWYAGcYwksFuzRsFN4SuS2SGFM9RzCWFpNc0xWJ5JVzhERCnNNqvyE3/zxVSu0NudRN5+qCReow
HW3BSWA0b6MyfOe9FfLcAGUoxjIEEtkgN4gbDAeBW9C66LH3sRPZiMPCapMu6GgrnYrLpMndCt4T
n3S+21Fz3Q7CO6x/gCanQd3ndYyJ29S+Q9TrNUKb3C5AboDj8chxSsA6qrl+pkpzxDxFVHG9pnlJ
7GrBBTz2J7rnMadJnDjg0oCnr6UdogSAG6ISqKwQMUrowHHws5o6v5O70VenLO1orklYBaUQVVjL
gfYa5OySj2SbBgyzzTOIr7v9Z4SnG2Ha1vhVAJOuW66kuukwaOAqxn1ztgfyNs+xxrP83E7F4tz7
aPwTatDWb9W49d198pP3u0ddRIIlE8wGI0ot1GSiiRk8Rntyl/RnLpEpHxXkn5VQ8K+3514AlBLE
k/1WId3s8QufK8BPV2cyCifwDE/gAhjeyT/m45QRVLi6XxgIiFrB00Y0198J+6iUYiPhN3z3hDuE
l5A85tOvYSQZdcOVhFViwEaeEzuYqcuBLWRT+QTMPNAAr74cN3oWmP6bb7bDIn99Q8tVEGXCSp/c
kGTkOdZRxDPKVtJcwf7yDOi+ZivLTHRScobjP0n3vQF8ymcahdxIHC7OIAncQdJ5ueR4xLZPXMRU
mhjSbvwEaf/92/5viogVOgtJ9NJnw5ahFd5A4EG+jE505YS5TcZ1TL8rxyYk5xfmj5fOrElnb4Dk
SUZPrH9/qaM/PNPqYfbjIVWnrXSgJXh+nCTkEuxNpCMm0AixwIr+qKcbVoclZBEj5/SP+Q+h6A0K
Kfo5Xc4xwojUyOwYqYxB5LB+h1chE9brScT/fjlCyYTV4G3UhhrsPb22u5k4cGxMYeWUgchHn2u6
eh4pqD/lgrLssfwKljOUq+wVzAoLqiXNzfj0Gazt0WK4EJaEDaj2aF+nwRt0Ls8LezwmePp3yZVi
q0XfJTSOtcx4ZZj7Wh2prnGECA8BXC9QwSPPLnLRy80Y7qXGhqZCwmQeKoHWyyib2msJfbBfeqZY
fe5+FeVEm6CRf7nUB5rTWTER1nG4Mh9pg9nHJQa4V4GlD7xyqMDXN/BDijcLCfQ3yv+jPS7BEoei
9YhKuS8nKr2eCyg/4zzvnYyzWY9yaZNhIiKyVK9ufFsaro3QGWEKZxXZhUpJe0DeO/hCTbFTtTHy
GCRrd7yKRXzawLDQTqZJR5VTMNTynP7iYCDHcUOOGfWK647ltNiMpP+1hyvL4QPnTQBlk3duXgN6
eYUs4NOgk7gKgEcHs2AiVh7ZYIS1pz7bZX0FATNlQOCQedX5vKF2DQDqCYasivdvilVpSDVhJ0DW
/w2RSnj45TwfJ7JLFjTUCG7mMDFFyJq/nQtEoWOqJ05FeWew+3AhfDjaqz28IiNn3Jn1iDzk8haK
vz0RtJyl3vyuXxN95Y4dRrmVr+s4FkV6o/LYneAM8tedQYFnb7J6/z7TF9+Xhf8yulUig6vu+kGr
zEUmh2UnJWkocAXFOu3YPGtk2umBP35DFn9oybchH+gchBk8BIPIrp/Z7CSpOlVKV5QXa719Sq1C
DY+WbRVKKvPLQ29BXjEroTuIKDmkisr6myRpVhA0EBMxpQP7FzU7GqmPpFNrJMsFzcllSjCzE0vo
gGKkr5yw3EAiOBt1F3eEIZZA7EiMBzbongxmCrWd+bHyBiLTp+dIN0SiSW5pFz7hTU3pBoDO7Dlf
sOyzodv+T8+pZQ5/4/jv6VsKgucBm88jkvjWiafKhv+AWoRU13sG/qtN7JNkNxBsDY8HgbWKbAlB
bbbl9hfRDmIDD1cNRwienkTi0/eE8p0QxUr7KVK3wqNgrK0M34MpwN1x2LPAmeyn7ZdW3G4QAj4F
U5WVJLKUc2tLAy8r064jxPGutz3pc6WU6uV3kwRLcZkJE6L7xHyubjl3vauSoGbga9mWiigy/+FY
6mtCjmeF5uxrjmjSG2qLzaIr1aWBHAcV9m4V3HIxdmFE5diUCsM8jehlQXnpOb4rBf762AsJlLun
LApbczXYvZIUPtfYfz5dWh/n9ljEajz+UjL3mxAozih3FjYKI+7y8NVit8tNPoGNbdtIa6HSFrAW
Kgybqq1G2iXG4nxcgyVRggS+MwgBuGRJ09X/XN/0bs2OQkn8wTcWDDtQRX9PUyM2ih+0swwzl5E6
JOsMUqe3fPx1vqGnD+5XfvqQf0jhyuPx0wKhH1SyBJGANRE9MN6fOBI5H4LUxjr3y9KcE8uSapn8
Y12mob2iiIp7iG6dZsTcCkmF3v3kW6Tb9kLGphcYUtz4WovJ/L+X9AW/XHjoMbotvLHphoti9aQf
7EvXPjE7ly6YLZIa+wSwSDqFnp/gSwB8ic1TiAqyxqChwLLyvp/N6Eh88MzD2RTjtdr9wqEr9Kl7
pwjjY5vFutW5llH+E+nnyNz/V0uP5Lm/bPGqugDdN7E9Gx0wPqa/fIUhU/XELPVsjaDEtdbEoWJH
7nO6k+35k+vdElQ9e1TycaVbg/+qbT9ntj4I9g/eBQv2W7LOb62l1QgunkEyr0uJqwUBLum4uUhT
qWcFOLCoxkiAzKZ5pgpHMT55EHeigcG+rEm+5W2D+FjxkXiBpIrP8UJ694c/+vEncpUrRsx3rfZm
cuoW6rLHAvbf3JOR2C/rzHxSlPRumUt12w7E2tAvaP17oBg21NYt9sqnwrZiswy02HFvCz62E42F
vu6J9QCWVDXrJyEVoRXgY97aPp/n5HGC+2y5HJ++CGVyNBzbod89U/5ibcbAQ1Kq/puQnyHzyUOJ
9UUinunWmBiGqPXhJ2GRAT9CJd/IsZDLSfRtubYiBU76i4Fk4AIw1e5Ak61AKB3yNhVIc9Nndxx4
Meab/RM5fmiWk7zEFdDgDsbaHCf8apn1bzc6w/bexEAtFhKOmXmj444LbsXfphEKUDa+rlFNfapu
n0qTDozOVRlfoOSbAeDBw6P/q48zAhKyc35Jx6nB13HT07rSeZD3nRVvwOYunlIsRUXZZr4SsikB
fEvpBEu3gckxby6OnO/KNbvTu+sx22t73icpGTrwZtKqaIitVkz+WdilRCFZYTPJPv/DpNakFQBr
5/ycMEnpqa/E7Le+1J6yESUp3jr2PvJXrLbegfgWhZKxH4tZvN8Ta80PdB4ROmpKV48dpzQl7oeX
QKSe5CvU345MYbSYTu/E17jydc8QoJy69gt2va2vrCxhwT+9hUGjeXOdIYYvDw2gvYSqeAnHk1Kh
1NtQu+UA4o8oQ9jGQuWMyWGIjQvmXlWHAFluQ1GhigwDF26q6MxToHzUCxiTPX1eZOTO82TFn3KJ
qdGSTLnuXcRot9zTEbK021V4vdRyO9DFDuwpXOvLcPIpkPzWRfjs88kCoipV5q2Oj4csf1slAVaY
bvvvVhwCM7Bu7NrD9ibzfZcFXfcnYUzBQXvV3eO4kZl2oLAMsObJ07yg0qCrB80rpc1vOENDrcZM
ox+ITI9gnt79+JBSbpdHeFvNqBZvb5qBBCS//jIXDo66n4xwH9dpuL9UuOHN/bjvqg6brxKzb7To
N8Qd5YEfSG6QlvdQcC7T1wWwzrhLuwDLXAhCPaO2+fNaT03AM+67j7QZSJZJEPbUeTZKBFlN4on/
UM25dPH6Sozwc0KodC5mlLZObmqg+GiMaZHniAY5G/+Rm3+p/hSyI3xf3L+o48cMxkG/ddDsTX6J
ygsnNuGOvc0ecPVfyhNJMJTUVPp01rc6Ey6E2UCoGPp/4ZrH1Iae7YL1BFa5MQoqeCcxWrNOPVDy
R5u7OjBEh82Vnp0IvhT7LHLpz4DbYfLxMl8DdKChkaYJMDFenB9K889fBcbHTgQlee/vOrXHxHzG
QHyzngRr99Y7P9F0rA1wTis+QWmx08xl7Ubnxqeo91BgL43Z4/aELninCNsKI0YayAfeI1GaqwmY
5cLZVPc//DNlFi2zT03AiUYtOvkxt7z59CpWygn40Snnnc1y5RoIW7EJ2oNs+Gi+dYQwyShBaa+h
o0V7IW9IrBZmropMiTX+Oy0PmH5vWPEIEMtRSFehMpX7ju/Gb6g7foIjC3zDm1ugqH8GHJkwE60T
7eh/7xv+MZRiXSbqr0IyGOeHb9WaOD2vYC0WbUnP4KSKgCaJvQPZYLhsbHoUEBGPhsxfVhZ4XioP
JYYPaZ+7sjY+InEhhFFOHf7mlGmYoXpUMMzq0uiZ2EPbHzafIyBgDEEOddN97plrwE9sSicKtcUt
Ng0coYOxNsz/jyLIWixSJTEoE+3gLTjkWNZfejfOMtsQodUqNOnPz+VKikqOdLxTtKDfTF+GZFWg
tSKzmUWbuSzCVl89MV+sxxZTWZlHVipX1bjoErq22p0/M+QYVnxR/2Bkp89jyh5foTlDC7AgX+gy
BgkAXJ9ZDDQ9RPAfjrzuc19bv3x1brRolRJ37CCxyJNBmzViQDfG68IdCyYYqzU1XdQNzCPC2tNu
/NroE2OMxwHbyoarXMGippO/BATcE8P9+57L5qBwK3ZPO175EinkXvst6YKhXHYDFt4ybxl/b3vI
aClqKAGniyZJdzpdkfKZsJH0hznYX9EyGIrN4ZupnEmuav4hpSvl5+YomI1ZmDTdQGSQW3JTO2nF
BlWKkrFtZoNYSLYVTXgsHOyEWTMpI0brXgGKxmWGDzfKoilrBLCgoI8dJuXKUyGfvDE4wfd4/Xsj
txJejH9RR6JoiJQBNKO62ftP1UxTAQWj4xUhKUlUhackBHKzIlw3+heawAFrF9KnYCNnZP87GiZs
gmYv0VIr6/VMLpd8DfI6K+ISjnyioow3g33AfhGxCF0q/jJLUJYi5+XboZAhK0cq1LdAuNjk+YVl
ESFvJX429l+hpFev8+uwSrjNcGKJF/PK/B/BM5Z6iEZGVjeBjHctaZHqec5sYTIQMr5ycIRoCwIa
yhW/kl8yp//63VRNXewWmpVO7yGnU/kIx1eb5n8G3iedzIRPJp5u5M5hcVkrW7OuU2GItew88kVY
AxcYugcIyT+VH93Hrbumu01vdjjYZa2raT5S9d3LL269ItTS21jFcC+4ED3KQHaVIVgXvbMh4zML
/VTmUsQwjPmnZkFqj8fn6uUw1f/Idfg8Ml8+rBEbpJ1Ctt4WvTSLJljrbLqfPtGTYIhbieFS5GCK
KUYBzVRgzcUVpFohC+zH6AZ4JsQpT1qWMAtIMbqZj81H6/tB3l6Os37a8tRSLjNTMiC+uwr2kXdH
IVVZoQVwrZhipgVoWOpAICdAOnlYew9sb35X3ijOrUm7cD7pyiR+KhPLKIkmA/9q6fUMokonQ16D
jW4PRzZsTpGgOyuDlNsS9Rdu8F6iJ2XGVeFiiWOqy/hSrqasepbbkfFZgKpTh3/GhzrQV/d+Q97h
EvF5+B+uYTI04MXSiylEJX3ynUWNE88wQ9iVqHQ2UwS6SW+t9OkRJFRss1Iwaib2YqEewQsQrh5j
v97562I5KhgCEETRd7u3rkXGnUVhR2uuXwcimaZrFAemVXrBxUt9lGRcV0dQvhsg1xHSc3KK/inn
SsGNHZtjnKI+Ql8T1D1inriVSEJ1RrddYVXVQW7OQ4xqpHzyu24F0j/cCDb1fGYzqZ8tNZ3r7cb6
3qmvaPLt0BjyRPBS2astv5QFsFgRT5/XeuRigbPG8F2jJEgItgDfWjKxpTe/2TrRPd5UcX4T041j
7sfr/tWioelJhOXmn8ZG6xnypOFsy7dk+9SHOE8q1MHg6FYNFFCI3qeqMFGVV90ZVo+WM80Azkzb
j1QqRnX4yoLMI/eIJxWY06R2WLpJOIqyu/6QhCNHYAlrY2/ewNXMTVjT+VDPhwZrAg+Lf4YjfVoG
02nyoB0i6gnyai4VEwoT29sPWW490mvvyfLgYoZ+jYoTvQoV2B077k0Nh2qyW6WHWVpQVwTCRTYw
yCtHsd1+ygFomn8AkVNUDdobLJyzuw1VGldBM6msxJEEszzrzn9NBnSU/8MXLZILqWY8vxODJtx7
IGuqBY8ZUjCgvftoKHMUyX09iZ3aLZVpbh1M8Krd1lAflXzBlnBwEq0ou+izN2g444Mw7gCco+QA
R+H0kX6uaMMxf4yNIAYgGpmTmvRdxBgiANlLij4z8JYR8hzkM+p4rIp+8r2cus/0StkCwCvSxXHs
E5jJF//EnuBtiP1OFVFY9X23wvC/ryaxjkhw8+Qu7imxytgHiL0QRt0b40wgv63xerXtxfP7lFqV
/4FeBmM62wGA/GAom8hYuMWJZrV5D5gkt7eSadrFHpvrgTzBWU60b+AlwgrCuIqdM0cR65OmMzxb
uFIGLsIRpMy5PyPf5d12PjzcHpJNKrZTXnA+TjXgMDMIDuSoUbejvOn2h1iqh7m+7GOidse+FlC8
sFSBKAKD90B/Tp23lWwwXA9Q+GCFy5dLs9BKzjh7N3dYVA8CucXNqUMdkt+KwytsOns6eNw/sbSA
RCOIydJQkCkbNNTlEIVV4/3beOFzxQHt04EiYB6boDOIM3q5uyCeVJmkY258lJuUZqthCjvWiGBg
Dwfa4fR+S2NC5hjUszrCJMFOiNhAYWyAkeTUNfWPKq00cMKdZoVR8QlSkekPHqDaH6kyOBc9qt6I
9UJteAE5EPGNf0L9sIS0Scul2bb2shF2RsAKvIk5R0SgqWxcFCliQrwQVbwjFsmaCMMBj/XrUOPE
rRTCJ5t5WxT4THQqkjsV9AUVwyDDDOb3sL85f7GsZHMnmuBbwFaArxIZzjRYYpwilomXKlIA4IWY
5XDfpHKRMkPCAoRPuEOtlj70HhPWnq6QOeoHxN4lIhcBXFuS+RIV2mPl5aErWo65GY77mWW7GfDc
uN9GJJpPlcCSnb/LzGstuhJa68fXc8t1W49/vlia0bHbDV9l+EgMTYRyDympFiis7f02AzIXf6O6
2oblgywFdb1GY5Fsq1Mu76/sWXYrRFDnXsYcQSByvUbWjSzUfxd1VAIw3d6bt34farBPABa+fo2C
vOBodll2AMgoWk2mXQB1GMHPpAYWwVyUThBmdgNkQL8RtEPMqWSUBqChepEvIsrlF4UHgKKKVYti
p2jC+TITspTRW2TP591Mi5189GtFxDaoAZ/uB/g3TF2Fq4Ks3WT7TThWeKQAbL7z37UAasQgf4sc
nFzk2QpLVu5YN1ioRpbU3P6M9bxRMIR3P0bKQrKVAuWKU80HezGetMFr5gJJdnr05zTuFljQ8oBW
CThq8GZ1XG+j3eflLKYDWw7OGgnWOndGYARETcmZdO+mCM6MoEzFctgoGkZtxEC8+XSywYcViaFh
SCDQ0KY6MW5aBJ9NmDQ1O8FAEPL5ZWPJPGH5M0JuEjQk89FADNa/ISsqOvFq1wpjjUOOgCQ4wcWc
3UPPCpbU0Ovq74akI8HLhP9BPCLXT+nI4XecxA6djO+A/+8qMoS1gUKu1Q6oh9Q9HX1WPKpt6ysY
hheoAf6ia6X3jCVX6zeX3+PhslUiDyLnB9XIq3oO8EKXz7ReQqFmTbeQ7ymZC1HVf41Kqry+MKuK
55ik6M5xh4RaNHD/E2iReH2jvRzmRbNnicl4pE+34ndEmt8MRDUv6T2j4uLvv6cRr96g2U/6HwCu
j79kg4OSlcbd1VnWPbKjZTMkz9k8QfYB37Jsr8qAfMIRZNuWEkOIcylHKqGeu3n5w/Mi0celv6FK
sMvpiSGeLTCMyrFWhrjXaa6AbzRqMmwDcGawNU3SBTxteH3zgCjgvhgIpCAo1uYqYm8hCbafXsSg
IG3a1+zO/9PFTjY4r4pC2BwmiWdYFx/T23iDlOJlFXBX9dbnaVwVRTY/5y013jfH7+aL+mSCaRis
oR3MmLqFdlvZjfJjyUmVhh/JNsLG4tLa5jxemIKQgLVs/TNMnMYMJFzVUuljxLdlOQJPoizz2SUX
3PPsbkfKHa6jrg9jp6QF7r9iFVF2AILgxqGQmkQD5CZCxBLYy75fTuIlgz69CrzUtT18aNLEK/ZP
Oa9IFqwvHqXapMyjcO+23gWbpGoAwnBCLOyPolo5ATkWUCLKftdqjpjGGmZZK2f/uECSIFEHKEpq
RTHK2dfSD/pYqciFEDOfpdwmWX4Kocz41hLxun1WGcumHHuogMPARkHG3FVl2JFOaSYSN3Y/nqDb
ox9srLpVJJVQF9vPftapICCKfGljOfjcNlAYFuvkDZwtoX8abRkZVPZeXJbrfGDISVSfh9e3vYqz
vjTMgnWGsjVfOk/HTAFkfPAdfp3aHXzUc3n/Ynorr8ZAGjTRHKa2JBZStGoZUj8rrU/vdXnZ0kxO
qXxSVfjhu4PWZFLUCHHI06C3iZU3ap58vQ6DHCze4J7zWmk4fVCYXpdTdnE/nJ/HDO1NJrLEJzEQ
A3aXkRK8EwN0uJf1/3nHxmieakeTzneUbmM7xGefo98hoTkPE9pPkIQuby3443SWieq0Diq83xq3
zI88GfpQ84rtz7eUggx2Yc1XuIJC+D0UMxUwqCBzNm+wFAiQCxwoC0Kk5cvbg54pX6xY25EWjxOj
wanOqS/GrfvXt3yRZRBCCRPIa84d1LrVvIUETcchGVmbB6LAVf3stpQoxuO3QP0g4FHIPlpTQirT
WVQEharDxHzQhcczqYY8OnV3FyPTXdvFfETlwG2CsPkrym4w2TwlyZO40/LhUF81Ab4Ty5kGOSzh
pnEQQiYFTZAOJo8F3CSf9t1V2YSZ17E+A+kkEIDGtLMI0zxMAjNEvOHnZYoNs4IcxVFz+mD5mcev
3MbOaHEJx/MF1II4mm947Sn+P6Qtne1+ylQ9fd0GXruvOZBRCqBidqK/vFoTCKCW3Brg+UP4GjFX
alBBwt33MEgpMJSuIq1zl66CUpVZhFiA5QrK+6f53XG5GeyDsahV9Xa0OesxzhwZBp2L/FER1Lvp
oIjQUj2zAd0+5ryXPqkaRPZF1YjxuRX+t/a1yBgYWFlpkaKsOmstTvNLlomqZ0s7VYelQaktawm4
LAJ7e7LdR+H6oGx1jD3VOIRvpBfdOPyzHuen0oRqP3pbeWf0ejW7oEpwz1vI0vo07ek8AvnjMNPF
M6oHLN+eFNR52I0+cT6FqzB1XblhuDdc0vLVCj98Nvk2KykDbgOc0D6OtkDRuRePsL2PqeK+XWZV
7z7F7+D91rkba3C1uiUnuvb7WkgxRVk9I3Ej394pJDf17scrVdH23cUEmdv1Cpol23zUlSvQgg6Q
mXrpWVHM3iaoDi6cLEctZy5gnMCP1bCaWL15HGWBXKdhPmUXZ97Sl56BGONDbAUW8pXEh3sfDqfg
tZDI38ftQXp3LkzpGXS2x1v8w/Jl7KiGBFm2p6jXsmKxYmNV0Fk8hu1y2+OoUNj/Fq2bdBLHlDHC
D8P2xHvkYSKBBMrzEQz+3T3VhmqTFfZMofM88VHHAQLC/Q/UGkzpHuRxoCj58VV1TpXnAH448Ih5
09eyxIURTekbWZl2t8eurXmuejxDPRKKkArYThBtaQgzAjQGoEgjhWw0utGleIEX4NmcU8Wm67jn
YjU+lPWFTXPGv708fa9eZU87AoNrYdrgSN6qbiByGYSIB6x38qGjrsMEOu7ZrwFSGKTJs6fDwEmy
3C4a87wk5osPEW/VZPdO8T+faPDIGcWAQacpky+pmPZewCLp18FrVco/gC+Rr5lMkVZ3wrPbqT1v
/19PdGS07WR1zEPrTfdmE5BT6q98TQvOqXajr+G2NZEB+YjUbhCXpWTA+nuj4HY2cSgkdMT9F+HI
TORx5QNB0Xb3qyoonKf5X6cWnqB6VzIeQJs4PFmVUpcSo+sPshlsTtygdCPydttnQ7B7BWiZP8Ub
sbI2xYQIfCHB/JYBgjc+7llEFdzObz9oZgY2mUgguU+VQvfi3L2RDFXOAc69hpEMhpeO/ewo4kfS
2KAzhNQevFqP2zP52POtbRiPUfPtGjFMPu5IIaA2+0/PNY0CPA9J88Vz3JhmDaViXa3U94OzkaVh
BfPo7sfE8OAPawO095BLQyBnNbpxAmTfFg6TLCnZmbweQnw9Oiz/Z7R2kwim39VEYS0fmiXvRPv+
zL6Bk6E1KXST2t33BjyhLmeRjJpGRNrbUsnmtWnm8MW5ZKbww78aD7FeUPO2+0sN7I/J0mFhulNL
4KO0nsmp1vxt6oKu6/oVLrZil3M6Dy+q9lNHSIlz2xk6sAgbyH5/yWZKg0/EQcGuJvTTSDkOk+E6
DQw2Snyu0zREueXqEALPn8U+mfl4bqgtrfecISCA9e7n1DGjk2LucCUJrzXzncbj+0mTdLCFl+qP
p3iJWdgyWXwfI4Yox90XG0LtYyfjxadPGswP4hIQvdLksX28rYD8X2hBNtRN7XKDFLbKw7TAGstE
nGlCriK9hpHNmlgfkVU+ma/OSF7V7kVxk21tb0OoH81EvBK4FwyS74pvnKDV+UYECesmYYkew1vL
1hO+PHETsAiBg19q9UikIdCs4zQbbObOsESGvajMSLa5sVwC4AeuamvA3YVM+3Y5mIdbJkeHPIv3
25TDgZ8Rviemc29kd70i2LbnamWjzW2QsN195lsNyZWKVc2npJbRaGkPkJdbfz/cfPBaw2WUalrS
/PiO5XVPJiAb9o0QWOhAHPhlduKT3lqOxaodouYofXtSCZwM6m/xybM8rWenjpW06+Je/iZZV/SZ
qcw2R9elbcFrIPj76yXpid/YsLaWkuofBWSy2zBrpeF0IlsAUvgRjES3tAMPBK/oc+t8XM6Xj1uk
qCKGXhxH0cNwhaNhpfIcvtzVvzij5+FK47QBUH20m2Jqupp400n57cHHCejs7qlkrIJswaBwCZ+6
44js9D2iJfyUg9jfWwl1vp0sR+FrFRZ9yJASVxyMjg4JcjYZOYl2QXUEALi3KESIxlmRog+cnnbr
a7b+RBMoW6GNXhgH8/eQTEDRevIn6KhQx8f47ygL/eP0B2apX5XzQPhSwBGN1Omaw3ILboTeh8ou
/cSfE5VnNJfQ4H+EV60a/njCbKWjFrO3jtoQ4XSYvbfPMP/j4uxCy1NR5BUSYIwTVF1KJGaE5/Vk
wsefcbbhX5as/ekuDE8eKixHCEdrMC7JBb8MPztF0otyQKYhVQSEMPN6c1SCxlMJyjPu5jLk3bVl
ixOgFpW3PmvJ6rDetJCUI6wf88ECwbmd4m4Aj6JY0/uikqPPAyFEHFEVuWIo8twvStCt3PrGsQ9a
eZlTuWAgcJczi33T5w4mAptJkPtoDXgKoSt//uuJP9P1GSha3u97AcqvN6r6sXJcStN2GCxbO6/y
16hP/60IXiOEuMacW1Jn9DIIzgoi164JnEttwG0pXjtgDAvJbnd0V3RVIDphpP6DasMW8AZketS0
pKqin/UJ4x4fS/8w4CE99yPjgJibV4oSp82kYsaB+Y0lxaEnOtX29AtdcTgY1xOXAk3aoAke9ZmA
5dsRKOuOWYEPT6AGsgcnjo8VlFABUH7Lx/r2LIXc+3Qqio6VRFDTgC65mBQBcxLaHb3jwpkQa/8D
nsajA5jgvLsl01j4psyA4gTxdzMPef0MmorOghoGFlmFH8gdx4YCE3zCa8IEa+ZNGDo8VRFq+kBe
uRWoxFC46B8dYmocEj+W5VBECVgWI89qYI4cLp4fxUKPHrYqNtQ3t9DOIkHndDBVybOI51wSWV12
raNlz1i3bwNTPabJiuARGdUq908AqHK+dn+3P0+T4uTUw+aUgVySu+6SgoQCzpUvG3R5g0eSb3HG
+WlAahAkohJq9i2FlQSbM8yPaIIv+hQ9odxBDa4TwV5QEuiV3r9SJYPQY2xsCX4Ul7y4toSZy5DJ
FCaGPMdpU/ju+j6zS4Ndw10uLnEwffU0LCIjp6odKgh0tukA0fr1tO3SbBtS57Hg46rVczms8UgU
l64jWDy7gqDok7AcF5/OsxFQm2hx4Z7H5pZL2gpQz7Hx25vxdJiq35psYgTi4+8YE9ypPSKBvPea
eenuWtpztlpTe2M4Kx60HtM4YqdHSCQpo5N2Pc8tqMyJJy2OcwnUpbGOeTZBxBW5VUlqKuvFD1c2
9QorAtWl4J05bvSY55Q7p4/2jyt6kC2hhe6MsO+8FH+KDtsioKgSt3KQUo10oI5qUiuTrUlpIBdg
J5f9dp2yaus6Fu1eDpfPvB8Bil+Jnz/ncQY7znMp28X9cgeEwSYJxDy9fUZVCNFJyqJ8C1TsEe2R
4rXpFpBiqaeJjb19JhTZiCyasYP/fR9h0Pht9tglLuuhChuYUW2J6ylmeU7Ilx69S1EZgvtLOzL7
JMUNp8WJTkKncp4Q0LjVTHnbWHk4HHUMP8cZ7O3/0nEspqREO/pr648/+LLYkkgIIVVrblNhOber
xr7kr3sHqrULHsrzupi1frC+dYy8hX8yRJlvM+I+q2j22sHd8JMcmyxJ0rLpjQyWE9/KVzQG/1Hf
YTgXNPQLzMdIK4+gMEluxO27Y6MpqDSAh5jqIznQv9JrhweRuUCmn+bcIYBdQfqs5qkquhcEeGtA
lrHcuWRw2PZv9IYnAW1XkZW8F1x+fEXP4Fr6bzHtexvoVHcsXvLgvkYL88QdbcS9WE8WixzIfDQS
Vi2EYzk9C7pK7PD17vSKdZxG8elU3MbeOje8yer0u17kqAWxA5HsBqpltEE2iJgWkhQjkLKWVYWB
Qtigbslk9VXB20VwAChn3OgA6uAJ0BpFZ0CYA9ShtSn4VZ6fMwLjqb1wSe+HAXHKq3Ob/ZJ4ODOR
mCJodfk7iV/TlFXHVClPqFNU+nRv2bpylbDbhE7THCLVuVUUiHwc//Nv1Ko2dyZQQOe6B+iE12SL
gB+BEroU3u+BqfUJ35nNH7DWEfv0JB4plgfEFNe3+UsloOE4NNRAcRulX7wU8VZJfZ5kr7x8u5kg
Jt0zJ5PyUUBD0zziGXAikHxundq+0h0gqTcRw3BosW5d+nw5x3QgQRZIzxkcd6g6PW2K250J0sz0
R/edoHPHwMU+iV1n8LeWqCg7Rg4fiGRtIpqlabDX8V1JpV/3UUDczGhHtxuO5Gva/Nr4ctTsAWck
ZWXSePP9VLH2HBjUnZLo3qGA5kKk+Aw9s8cmntEdXvPPwRzvRp+wTp1MxGsWM/W6X6BVKIK/yyor
gVw4RSWq7yT8cApzpP7H1Gxtp+GKARFVOrnnDEk2dtGgToA2L9fYjX/PG5T+5NmDbRRyVz9IBNoD
d+igeZretMXpSpOtFl7rRLAr9sAcbqu5c3dLCivkCxh8pqjwo/1Chs4X1SFVnwI69zydL+nRkpum
YKrQigPYYL7mZIFhusQZMA2RDLa44DfIht9hvqsU8CvH83qk3PzNWh8SWCyvp8j7cdq+WHA2JOe5
WRV7H7q0umMjHP6DJ4v1HzNY+wyDMKZq+awqXrRVrdxTnkj/aJz4WtF780kixHz1sMN8Gnza3FlH
xPKGm20LAKmPsF5kQA5PJHpbVOcbAQwdbco1PUCoAHxBOyzOKc2Qot0Ea/260ovwyHyUkjnpUVER
8WhU08pVZtF4dIaOYQtvM0RZ6f5lMaPOrFRxx9siOrL7d1swRHWQ28bltOECkJ8wIRtb8eJU1ZdJ
x7VOHN824xe3Xa5kq/pCeye46s1Oo2Xrm4tt9a1JjrM28Y4c4YAgQeuPSWOnNowOJSRSwpV5hqw0
HhKsyzxwjHj2qV1ppS0q12/90mUoiHQYI75Y1Q/ol5s+eJtoXN1CX03uNWwCNDr2tfr2Vi1xGwD1
13Lr66z4SBPnhj7YHg8ezTnR8aUm7bJEkdY4m8l1yrxTDYV9NDqu9/NugJYOSHcol8ZZyizzxJHh
31322jGyiDuqjDWwOhFKKB2D5fbPGYJEPgsvcoR3/bVzVasM1DPrWdg0CO6xRgE8DyybEJ1K4VAf
lKTcyf8qluRchEA3V92Af7UVy9pg+Bkwq7Ttp3kB+aQE1oMcj41XJEJF0h81G8QtDlFqpog6mnH1
8KN1LtvPTj7MUBv1F9fvq/vrnbJCnQF68v0uWap6Z4uzMsMWsjnW9/agOrA12mVlvS5I836/yYqO
cVI0flsDSlNeCrPCIZQ1nLqnNPqgE3Iyy1Wxo1HObG8TOiAS45DtnoFm1E1aSnTcU2UR74i55QoG
Dqap14FwMhiIqLWYkKIHp+23ncrtYRbuwXvcZg6/IxIGwYxK9BvWSgacTUpFS/XEJA3twklli9tT
RYZoWK5S8jScMTH3uPhzBIVdi3moKLuXb9Ez7yuih8ZvOndO207PqI06aKgU4dslMgxm6ZDPz8Dc
UJbh9z8ZWA9nZwhqdFKTUm7DjaMgCzQsiGhsnAZg7FK1Q6FWFspVENgE38zlkWaHC8X8ijm89OyR
0pZo/CpBDsY4VjiTSsbXaUd3WYW3y2kctcd9AqsC/KBobifGisQQ7chA9JgEjRGkeFKN/zkup7Te
ODCWoehUmrZ9ioavb2gKksqIjrwVvQOUOoj7QbUXWSvbTgtuMFZJUvUcAGM1eD+49ucW59pZiPMH
mim++8Uchl+HgTwIJIuEMXfbO3RjBa+8G4VE3xMrAbQKDP3NnjeVcQSorLZTANBemwJg7cv+berS
nVt6/H/fZubeeqkjW83J4ivLfHdH3RafDhmAWFl7AzXa73mtOQDNiGOjHWb2uYaEnQhXZiB1XLNW
SJNQsJvtmFWjVS8BlCi3FzAPM0PeDjmUqY7Hcv9OT3wAz7hx9P+XcCVm9UWVxJEFLnNTTwPdcoP7
aESZYp9iPr51TgyUTXPjs5ORxwxrAxVUwC3w4xrErLfLkOKq1Wb7jpdw4XT1xscU0BPcc9X77Lzh
ykGtAJ1GKqyHkPHWrfAJoeu86IJYIKO/EQ5qJmrSjXminTtVRhWLzrS4bd/uLxIUqPWkJvGU4Eng
TumM3A2q82PdyJnI6lcz9qvC+nZsjX2JMbFav2SMEWVx2Om2XpKtvr0cFnP2fQaYU4klYCPsE/Eu
Xcnty8CIgAOXC76xujg+inL9Vsk4Qgb46+bWfvCZ1Qdlh8bkboY1QFjONmy9hB/FxGcNhthpX8RX
JHU2ZJ3gK8fl5wp9JlCdH/xkzYTZVFSFUdCtfbuc14xoAwAZdbnZ1MVzidh7AAOYY+hGOQluQCDu
mEjnmcYzv+FapoDSmIBA2iBMD6q50DVohwLsG3nB/Chm0JqVevfdmWB/wOBSdNrasOZRwMhrvhJD
DzKWJ7rZE7kxQ77d+4U1GL7ie9GYW8TS5Q5XzrDlC5JXaBEzhimq07jPDhw9u5aGWOI5BXKYBaNR
zd3xymdOYEafY1lWzVetRU0//BkBweKPcYgUylR1KKC3lqRO5hBIlTmt1IvosHwiR4w4+QHRvuXC
aehEwaCXV6uG5g2kJ0cPX/GvnLKUedtL0bvsyjMQD08OE8ObuS2INXoX1Xmqpxm5aiZiMOpuzR76
2XPFRqCijWbAvuz6x33bHVN4vNXnaISbZIgy76tp8rlvF1Fxd5585JOPvMdz0jda2BjKuPrts99T
ie9IqQSZDsnkT//S4BWOa2jS3dzz4KTDJUmOGc0nzcF2aVda+4EHxQmpKENhpijD5Pl2xTLP60OG
MIuw2u62TuEnTVAtpL9pxkdzQgVJOOjDFuhkqYp/pWysznYRavwQBxzHcUBQQdKZYNaHWjomYrSl
RgjlhIJUK7+hHYPs2VN7EJjs0GJKccKyBUrPL64HFV9ndX8fU3dnAIZLiHChFoBm0MVKNWIXfuIt
nuVSseO6h9bMlvY32fVCGjotqTvo45jnTn72i0RC4Tw+PceHiH53/PJLzf75TouIJrQvCFOob+Ma
njN83IuCpF/yI2oS2+Ch+BDB0mGKiYSJdnH0WvEqwL3pF8V7QNfK59Gmi96ka4nHS9+5QbIH937N
iKF7JtIJgfylTVm0L5pWFTdYq1wukDpfSsH84PrCO7WTZVwn7kak6H4pdrbAgJ6nYNfYOll7CZoh
y5EYVTxX/c860qbhGzWVVyvdyn2s5atwqOpexB6cg6gfWVv0DPOUlzI81N5mZSwLqJW1bNlCQ2lE
mrh26uz6xrxg66/KAt8yuQacAJFdTcGiJ+kWwemg/RwU94jtM5SaznUotbshmEIaDhmd9tGLftVb
fGdUHyI/VKjAeWw8KoAwJEAko28QOr9V1AiWDLzLE/fjXnDcysZFNsuRQI+Wdp3OmlpXlYHi2hQI
/2xDinZjs4s/RIwJmYMQJ6j/YVQuMlqAVk+gAfjBVVi3Cb/Vt785SSvdGhEDvSclkz9dlLgnXL5i
sI/vfSEJv4qHJRo5JyMdOY4T+pCLdglv5gqxzp+n+ggX5IZopTHgLTebYdFPqkVAtuVXQl0WnwLC
Lui9JCWuGFOpIkho6MN5z5dMy8WhjB8MELe7EC52fMt3Sfej+e532jzeTNtgGkHiBnwKLNARgNnq
C6t4ue6dnHgt+oGfK6xMAC7cs5hzhdOkblFiDjs+e+DLXSqIZaqc11r3A0WwRZ99DuXMijWgoGC4
s6fcOUIsCdNu1VfhX+v2BKhy57jD1QY12HEKumMqZ5FApNVrt4sfk8tdR7ssbInWaQsJCwVzg/Zu
4Q5I5JdfliXJUEx0EdPVGFFKZF3XmkQYQ7FJ3tC8fbLLQtbgzjIWKsA7VcV9P6mPileJT27ggOgU
5mIGXFvbcKX7wm2N5thkmGJjb8usRnu+kzY2m/cQsOX/UJbDT/zjf9ROySpACxE+2jRWp+rZ+Em6
p9GjGwzSFUtfp5Y3avgRGX5dFmrIrRb+05Z+tgAwQwvkTE5anT2ur9EfSNhOXxHZlsKV/9uPUR0X
MeEwvVlA9ewlKu7/WNG/FTcs9f3KB2abDYWZVdO/3GjpfUP26NztHB4bA9Ax/6HUeYqREZUCbgcs
d48hwJqN6cDRW5MSBBemBuwDJRjFXCWjhChU6S1/x9hJI/Yvi4IRFhLwdQrweMTgvqjYYiOvCPzO
L2olA6LFciAkrSU36zgLgtuJlQM/VtIAoy4WfLxtH449tLS3gEtXZ7uidVzCNNxii5fDgSYuMb52
CriTtrasYPTensgPd+qTLHHgAOSQmP277OH2oCLtuREg/n36RfGJVTw+w9X0gMC4rYW/ye/mtEkt
Oed3n9Qdik1bOEnO9/hQYlK849sOsD70KFdQT+6GW2JG67CzWYCexU8u4XOxWWAy76iqKFy467o6
UI1jScGGQru4IVUVRz3YUlzMhhHqY4KvDfSkln15ABc+sH2/pgRpU3sr4Q0gD8wP5FOJt6xXPBYc
bm0A0leWfYsieAXIueBm3t8RIEPaJQIWh/Sgd/a7P54KKkZFErcHrupMLTH16h6ItBkbJxix2PRD
+M79rQVorGzAtKRATAqJnL/9RY59sx+H0Tw4vS8fLHp6KEM5X0kaBXsx/8PQbgKeKHsxKSxvITkR
o5b50Z1vU9BmKmcCj2N6QQrVJ2ZewICAP7U1/ANnGkLJCvye8hRwM/A43GJHTKsjkrKyKFvebxpL
YXMzUqx1rMf/qXf6XdlECBh4+e69wp7yKo0H0rIhQZToT/o0s06HmNgkWKnfMEr/YNMgv2jqV8c3
acsxM6cugHCgx9y+QKzPGeMdNfDEzY2GCP0hw44Dj2xpoIH3LVmCY7dqYw/fV5fxK3MxWeu2R1vu
tzIrraaqkjDLpi+q1jqNqDeGQzK+KnegH+xYZ14dOrKGbMLOQBRz+x4lf4z2Ft1/xqk1bqKjd0+V
zXReHBARRaBNuS/R2jWpdq1xwSiOjrwa0oS0tUf8kvC5Y4+w+0bkfOWsz3yVbshqkcuXGcFyNFUY
PbzRQgUAsepn2x/FV42TzOal4nbPovHbuix21WglQccAstcTi9YZhv8TIX8KBxkt2xbW62OVcsED
MyZXE7p3HLEb+NMGudehPL8rSoXiUnciNKKcJy/XEbdb/JZtUc3nKIvOU8QdXYn6gX+mdxzbdWwA
hxgvPRvLwmUqIAPY4SSQDmavPSaP8z6WnaOCXGelJOiDEVxc6btLG96+LW/HNFK5U8OS/WZUpUuV
UkRdQJCt33wKEfKFZT9pYvZSlu8liBxlyo88CTMQGUdHzzOi/46/tyE7QOe6/dPk2SIUZpmZuHBw
W6UDgF/frcDH3YiUpc3Ur7bAlfe9w7vLeLL3qkUYnK4qUqEJEGE8+qPfw6TgJUvSn+dfuqvh8vVy
kNXw0Do0jbiWKTZmRk4HeRp9+ugostS3ExNp3T4SsBodPVpjsVVXONZ3axmLZS3oDqBXQQ2UqlNv
5J9fZOzjIz9j32kWarvKsLs/eoJDz1lZbW4tzEcdAq4Kx4ebNQ7R+Xkdh0DF54+haS+tEOdbZYpw
+fSvxzvl/xZS0+0gjv30fBjx6YyosDxD7HSv83BfRp04EY5Kxxaf/I8vnnfe3SrlKEpNvaZPTz09
xK4fvqh5KS7b8NzdvDTtA8nMJW9qFGdDUf+ArykYdXK1jie2x9Y/O16ahk04sECLwxzv+sYpcHA9
BcWHbY0dOexS4iW/lsYoupq7W23Df1iXaxQ8/UOFxvwxZJVcz3Yg8l3R6qoBAlkTP5ufxBdros9+
eDtL1nfE+QAD7eeWglss8GbJSK48dPwmXb7mv+Sh6XPZ9WRy+490o/F3ObxKbLkzRiMSCoDkkher
47cw1POhzDRf+iaz0gt6jO/mxtEyXh1oC7l/XiSC3shjSqj0TRN9ikVjfkZX07YMw5S52YM+rUpr
NWfmsv59K7UflzPLhr1ZBftYICD+CMVDRnCsZJF3c/vBLA+jLuaBtjIr89hQD1o7gTtbvW4c0Nib
kakfhKRKfyKvzUaqnPAKNXj41oILnzciOqxNs3T/jXceDhIsHkGFGufvFITysMvtn2II1x8RpILp
ue+9PYAQB6i9LzY1H6AbvGzU/+SS/wq76g5XQIBgAvVPEARS+K92S36usVDdADygHQsBpIfiuYzy
HlJNGpgrFXGqdmFvZNr1P3A9cE7mc3DI4dFYtqoS9BD12SJ7BRGVhmdar8nijCVt5LCIFOD9fmh9
l+AkaPEl0/kIwHXVE/zvHHXb065T1Wp1xb41CmmmnfJtQ/KO1+MTV7AY4ahjl+fWgRqITOEifFps
smGZcBhwNfd5q9wXKEll1dsxQr3DWXCRVvVUwRIBF+w15W4xLWGk0emnCss3Gsd+sNQK4L34HZcM
PVUCMT+wW7HibZxjViJNpvzthTsbJh1fykMot1v/awsQbEtLMrtVBC+q8aQcu6KbN2f/F/QIPtcC
MA+B5EocPOhbuj47T0MlSFVwUun5KFWoV9jOg60nlIJIO2pKeEYgCtnauq/Cse4sSiqTkTjtz/P9
t07ZdgnTbrKc9nsZUghFEt1GKHoeYQ1Gvxzo7BMj2arAZznh8RGw707U3TxJJ7co+SHRe4KFoICh
rYxMOYLpRgoZBcaPCnVJYsRSkqj8qFhM7cuPArxi0ctW9kIN7NlQ7Ll8/ICUun+MEK8RisRrdngg
9DnHiIdPzAZFjBet3nk6IhsaUzgtCxXDaB5J8tYRPmLH89385QOShrP+5wjNNOcKn2bkmRkBRDLW
X8/XEYJh2DdR1v3alxRXAb3mH2G/3l7w2KWrwLPzxC4jcEkBU4NO50j7k+eqMVPmhVn/YuAvo6oP
4e3adnFeJ9/AoIfyWHTaq2oWbkKrdxoEC2mKdGgltBe3iZHxvPerF2xe9xZXcFUYvKaVBjbI+nxI
Nr7M3PgfsOnpmnyw/mHtL82fSadTMX+8nMJQ/RyAFhRb1ItwpUjOeJ947NOBScKa4fa2hNBePWoY
8jBBRHXMJNgug/EczHCcreR4A8vRPpgpixO1QT1Nv9DQivWEua5qO9cUulZmc1uoTOE266HdlmYF
CcP7529jVLQaVreaVEXC21Q/Yur8Dj9m6PFimJDteIQSF0kdLOZvXHpvSPgh7k1ISv5E7gZeogFK
Bajrf41ZTqn9LCfnc5bzhfJg+MKBb0E24JBFHKqQdEBxfwLLtZmr1jYYPCF2+C88p66AfbvYBYy6
WTStY+MlxfxpzUhdDENfysTLk5VzYBG8+1bv1h2L8sEufaLYJ/7iTtQ3yp/PnfHJLAc/azH4eosk
7dVZ7NEr/dRRKG8gAG/njX43QLLQZT3ATqYQIxtATlV7vnYnraPMYbghUMwhbTG512PtEb7GIG84
HcceuA8726utW93Tz+kE8mBdi6/tUKKkGo3nZO6f9crj+fm06H80rjWX6P7A6kebuc+TqdyJSpMq
gTf6IUZyFr42YYcNo3NOqtnJGqflynh67xyW3B1eRtudwDVS+Op++y3Z+ZofojF3CZ5slXUkj5SM
1ORsMq54rJlW/HadeNVZzzJuAgmDg3rL0p4ke1YJAKtI0+NJ2WBTesSMkxcoxzg0TA5BF0CL8c4P
nHetl7JB/z+1sgLjG/ppNcz5SVj2mDS+eqwbC4CNG/KdWeE1Cl6Sda24FoCSzxDVCONkn9SbgDNW
7MMG/Z39VsqtvZFeK6R366+c/AUpXaqV89CPJaFF5xE9pfM6eQ+XsFW1mn2RqtQHDRfrnZ0B7AR7
sZEhlPKUggez2itwztixn+nGHAMdiZzuSsY77559HOuYOwRR5kEZYGjCm7KkN/TdHynCBYnMkWtQ
+cY/6DIeFZQL3Mdovnjpd7OHmcWdBwD5T/5TdR1Oe/P9NJZcoO2mh2n4flAO6HpwPgwqG/h/NzOC
veQVpuN5FBo8x6VrsSDIh607ELDqeGiCmQ8L5t2/UJERFsvWGV6qljW7ioKMHomNPcBMoxP3qSSS
tSpE19nCV+wKuqoXBpwyBO+aK0PHz4bI9ZCQMomQMAfRgbpOHKIVjqohOK50PQGx0j7SYFoDgxsj
Njhuty5P9dJ+l+BxNTzmd/hyJ/7IUwVuvvW9O7vGj3D7o0RAr4y5NnOkrs5D41044WQ53dpdWMGQ
MU5/h0GJMHcvBi4Pdq8GPUbAJUYLeeZ/dXSg7dCr+jjnzR8eBQaEwVWZVMVLDUciv/H+gDAb+jVW
vhF+6z7NXSB5mCk1q5OoyhbTtYBP9pb/bVp6aKy2gtBUkZqnArqAMcEZsyXTIrwoT8yLN3JcrLfj
LHgnFR69Mia8ycv0K43w16RpxLvnRiBLali1vv0m19TlKQ+nyIUCcc/LsK2YdLtaDJ5Wl/2e9uKE
lSsGy4SQCsj9gTh9hyDrMcTso93HT0vwoch+f3F2pnY7NzYx8vkazEXmLpwU5d+68/rmyAFQpgcF
O0Dlv50yzpVq2QK9WMmmU9JXbTfm9y/PP909WH2H+px62KKh1xmDiCFLasylUUOGjhxqWrRb36Yj
15UiE4xT2tRE+qNztn4QAOiSxsEmCT88u1oW42e5f6I7u3G1vWmZjrEYVjwgS6kGeDL6ad/sNWI0
8EvgyC8KUv4VJY+fIKOjowACu8flbrt0G99D0kRyJ3l/Knexc9Np76lSaLR7NfnAiKHrTaPszck5
44kOMx7sWWBJt5O5CJZV9JMa1XjnK48I50OHtymOGFsPpIE2ghbN5uIWDnz4+lHJdD0j+vStHJaw
zM5lbZaQYCqCpipHCr5Fr2ukisi7o/i2ThHfp4piZeI7tb1Y1ZLTeHPau70WLLre8eumfkl7C53V
T7wRwSlFG1XpkUtUNWPe+r4ps9SKJ3rDQR36JQMdCNg38beaMxf6Uc9/Kymz/hqX1o0QGukVo+pD
JelkIX2YPMnkMnqnrj4Eh/3IQE64ST6KHjEQbofBHVFdD7UIiahstPGI48w+bk9RKZon1xzZnps3
nEkfDC8m/roUiTo7B8F0A0r7NYAh5DJQrMhMXh76VecoY9sPffmv0+/q17snPohSTMwHPe2YP+NL
sfasGIwYn3VRvvrt+zZ/HEMcjotpvTjpWX3y2UbXJTK+fuRM3NlSjwxctg68KjwawhBKdphazDzq
79jDews5cAkCp3CFtGoqgnN4AqwDJZ279FqVd5exYkRYOMlqzU6HaMSawzqYvcDtpUCYBHYfZCYi
bfrKcxLcTnK81SEA4Z2x/Y7Mw61cJorfyQlOsTTuRHeEfOBX96GB0hieEJTj4blQ5tbMenhDV0Le
Wp6bjb7VtS3BHL9oZwXz+epmOJCaVL8WxrT/joyRuMAEEBkgxY2crfuG+3pAzYjdw6Tfs/yf8V8R
IO1QRnsXpMHXQtMUC+1ogyxyMRnMZfPDUp8TOM7rvrBjpmS0BwY8QwB2X2hJEKMersraHwaBy0H1
huzDDjH16aX0JSoQ93e2TrKC3aYm6gKX2GwRBIa9Aq0NoSj2jOWxQm+t2SSVi8IQ4z7Gvs2/MXb2
oYk9uykpYCNSdM8SW7mq99WjSOl53PmNEVGOZ40indIFaRv467TI3mUt5OHukmbri2TeV9xiEGXb
NKE7tEKib4BJYDc718GAV46Wku3IpsvPhtceHVNNXwQXJHnpk/Hwc3F84T6cY7uqj8nF72whlPXS
BqALIhPKYDVw7Cb2t85b4T+hSsbC0QFYxqc03anq5XHokx9SCOBR+yY7TPKGg8gkL7iH+VI0k6Yr
Cjc2GnYdlDEWhqTFIjX9+dtFfDYcKgc0UwWpSQuZvh1pyZyqOCmBlfzPP5tp7qlkLPzZgDsokxYe
31Tuc78R4pEXkgcZBctsbb3Dx3vRy6KXVlEV0FhVLwL/6UMRAhQBgEpBEumjXWv6Js3UFpHF72vF
9HHR4XP90ytDrvAYz8Byc5SyGQZW2UfeVCheolZiPge/rS59R7dfriV7/h1cSyaD+atQEFQsCPbe
YbTaLm10OVKx2+zTKUXzk92NSXWhvmKSESKlO7mfRcTvAOF3SUGdvueoEuIce6kDN7UkC+mj71tz
yM7Tg7Wez3K4I89RRx0HtMmMnnCX1Ue8WBuSkkIs5Adp+YwMNIeSZZyUgrhViylelpMd76+8BbaL
FngGHyWJ9tb0WH9RB0b981me1+dyW/VIbO/TVDVvrotX4gLmjhSiNaNMRXlxmOTscWqJ9p6Otm31
TdlOLUDSzDm9GDI29J6T1Go67vSylQZYX+mRRnbRYfbOx3OMypR+oyr09y9U2u2dEN5UUW2dvzlM
gxs60yzY+HEafVjjtPwme4MJknOoFDnZfeV6B/hADp/J9UHfmdlUrtbyMy4e+2yLEweRtLWPtdIc
8jIReRTjug9N2dKJtskePTHmBJU5atmB8cjDBVE5ndCJJYBMb3U9QbtqhHJsIsFZvyG2ievCqVXe
oPWmgul7A2rMeYCy/BDYsFmNNF2qiUPErTkq0W9tK4xEKPWB98SwJ7YPjp8keWwTQDhDTiVufgSC
Db/vWChYFqCMoMC7TpF2uxO2tbmQudOS97iurRHwQulREib+jJZKUXGDlBNZaXdbOETqFJvfVGVY
ZXU7Vn37PMNRNTAcqeBnMKA217l1+jFxPNcUzlrtOHSkydN0+poY7eJgpzksP3wDk4cdAr8HAKZX
oG5nuHbWDOxfCzJyWwDbdwLVBB3wQozQKVsZzJTAzun300Ho1t2kYwtLLFV/xhLnxs5IwpRmxf0z
ettmimqUmTFJrgaRbU1074ZtYMyrFv/U56oPgh02FY+ZNqCXp4zf4+kjTzdEJLXMpAL0GbB75fAY
cCj/sLADZkPaSCmwRDkV0Qfiw8Tya2X4YCJYA/N6B+W9VGdR/BQP32EOJ/XssCkdms9ClwVip+Qn
u/MjgTpI/fmMjt8cOHmLgA4Q5QgsD4P9Rybf/1q85Y5tZu2G2ducmaLdy0Cais0BgiTKKoQ4dSua
Izj7iMqC5mY2i87X6SSD19I0Y4eqHP9VtOCruKLdo1VNy+1j0wOU9C6VE83Wl3ly9jPventpumlK
gfHzGFSIYVNjGfduMFExKWO1zE8aIDsOdokXyxvTl2C/M+9EvXdn0FGnPWLpl52zMJGhjGs78Z9m
Wgar2vU7RkRyqtqLz/xhKtBRHND5Iil+i8uH96rxVdfYNIVWKgUZqr9UtNvsLi/Ejife9IjDjh/P
8snT4/VIhKyWqxmP2v6IQ5rIQm/A6naAaoLMrNEq037cbMhLah/dyn6nRDM+VWiGXAWUvkQX/jJ+
NoYiIf4jdKwnhcMUgfAw3drxZU8fAOeEttvl75WOl2EQ7rcAiYuiGiOScTwlwr4lfAukX5ehGmFM
zEHXAmLvn6jls0nu7Zo+oe9w6gA/NY1bkb2pbitu0UnMAhM4jnUSsrGcHMBrxsRHWaFPNpqsMvhg
zE9y0lCGJgMnnBL83z0n/EUWtnGaMXLNwIw0Wgg+QXd4zsNNIGPUMyW9bACcvEV1B/Sk3B8V//vs
RxuKijjFLrsZvJLI69Lt0e/wgcmq5Uvxqw+nhPmI81AWFjBSX46VM8+trb5a8E1aDf3AMGOm/Y3R
PGRLok9JTHMWI1eyYcL9LriU3YjqEYQRFibHjFC3ti6NKfE04Bopr2PB+p8n+d2frQDWJ39e+7i+
IBG9NgHkLDgogVYpn/61a+J6XkY9QrVPmQlmIS2FNaVVxXy65vWLoFXUif4w/kccyqBcyFRV2P94
jN7tBmmMLFAdloyEgur+elx4wa6P/hiw1THIOAWjy1tiC/qFeTBiKN/J9NXkdThx6mJI1lfUWXLa
nHEDLIhQynY09uYoY0GId+a/Yhp4b87D/fNrZV8S6qCcNnBXM6U/NGRV1pvwZo1jdYshTM1auq//
6+azo4ZOsGz7cFfi7qv119YgR8v5BfE0V2V+dFiOLAc2P2W8ImYZM7A6pRtDF9cPFRqIBqahaibU
+RwiUxcgTgSoAirAZxV33BcLms39P5c3uFSNeox5z+rvC1SaQYSZs60TrAxWWwNFdV4qkijzlf+q
epZ3PLv2Rn9LqpkBQ3Z4wA0f7AmFasbmTCpo9hAzoJ0PSeCGnJzUSFzgtpZl98y7mq5NhrMh1a16
HFYcnCZJhEGtMH0+QP1g7c3u4nSrMriMILlyj5iuO0cq9R6P3Xb8npnfSEHfjYUgpc/r0ZPIAB4k
foegZjIVVycF5r4m52LFm+bPVbCwxtvD9adnhzLOvdZKks9BHkvtynVft59/STjB8sw44DzXbdQ+
iPyfILP3pyxamZD/C3SyOi6W38lfmocMBnrwhPfA6SIEJR6TkCFtftEc5s0JDifDZuoK246V0mtJ
jAyI6GNWLaFZP0y/uq56sDc6j6GRLCvbNjLVa58seEB5poefpZ8nRmMfQepU+/ElGxerhLmB54/N
Y8NFvd/CGpQI26h+utED1kaILzA1LD3dCAg1T5C/AZ31emZlMDgduE2EWvKHbWfiXO4YFwfQD4y7
gVk29wDwSxGxbMVGML0ny/Ef1aThhqVKWXf+QdzmXPf24gtaQjbMcDkcJtD+Msoza9O9uEi/5r2Z
MIiNUgeKIyn0hXanCviDlKu/W9CtExU7a2fm2Vab/iEwETEEJgqhVD0feBurIk+7SCM0a2/kM6i7
m0F7Dcs55O7S2TlLjG8OsrsmdYmVflLyPjvN37066TfeF81MDPnI4uVuc5FL9VLA1ak87Uc1ZFQ/
vaNIUWucnwhflusgPhZULBxVFb081jGYRZF7qpe9HGZCJlaU7091rrnIvdX+EH00kqIIs5PIWO3H
xu1xt1Nq0LyWqDPWBvUJkTseVshHI2Lxwv8UTd4Dwhyax73KxbV9oPQ9gqae+5cmCZgL5eUu5dj6
Kh/GU6D6Yer1UvHlCZVnaPOV1bfpz15BAT+ewl9kixdC2yhjIDqqoshXF6xYitCI9QldiPJOz4Mk
sxGxyfqQHvtU51JcN+auX++nc9Ul8g5HAHEuVjOnUtXWaPdjimWCSShi1027VN08RjZvVm6Pr00H
IX6FsXYdSh6KFFzjOaj3aqL080mTxovx1QvTwam5q3Psn40MY0LCW0FM3JNf71LRQYGZMbTtRoKY
gQBVyRPMzAYQkJ/4x47Jmro+ef5OmV8Qe4fc5Bkb73wPds+dbOcixwKTvSXpYec+qUrTw0oYku5I
lfjg4ct0I6OxSxkFudhN82npN94VQuPIuVnIrmVCC74vFYyDMMIemPul4uU2YELbJ4aIf8DSBBIA
YySPFBwFoyIWckmklldCdwT0jMvj4f34XurkSrJGXG55Ni0rp/QbIGKsj7DknBGahvqhOnakZGNq
EIkXRb7lIHcy6mhGwMmYBGNuMS1/6eZmi+W7DYOjulzvw9gqg3isRx9llK+Yr5UTAmeNoA92I8qW
8p2Noe70yKVBkoB2ybbWKFLpQ0p0KEFLlD00qZ9DWAgWmqPclHR7mPB0HTuratIlUdEwo86exkmj
+P4dqHCdpz1mwpYIfDkvIP49dfqnRyRjDojIx9Zzns8uUgGSRlNwgjt9Wy//Ok9d0DUbOF0xTRfy
n3uYnpSAesNwVfPguj7pz+DNyfb+Ro12I/9ybP0crOcWTKByFJE6tRvJ6Lq/0VBOgVIMrw4phiTD
NT9Z0+yn4XZClVputJ14aoLiC7okcFDsvwWU/uAo+Ik86DTG5FwLuHs7oZt1vNIPjBiAmwW1uQjn
Zlsp1cyPWOzx3cjetUUWBWia/q3H1o/8szcVx5h7mdmCYwd8yd8BH5pRyGNYwJBkMgAXDD4nHVFu
u+0gsLobNLJjMg+33JzIzwKdlxtWIzxuqKbTfw61du7ECBBUy5CZswzseVmmDb+jZlUCYbkc34Bv
rEoSRGhFr36Qq/ZhEfgZxPky8xdhZ5uzu/5jnilWErT/maXpAf8Ren3u879KqwM6WXQqQdnqHWib
aIYlZ5Zer2nTmyl82pW5eApI7wxqhvgiIYuNesCN6uivDZtxbnbhZvd73wkrIPkh7+Zgyj/By22+
MUbWPh102GXn7TUZ9r9iVQWL/F6zdQJTHzZrjJyL+BihIv6jmnynnG/1MEEcR/LidBYEwCdPUq2y
lVt9CzXnROo0VvOJUTsXJDLmdsuVoNIXxXvCCY/wp3CMpXe3B/y/RREsoOk61O2SonUifklB+WSX
ONBPMKHE+CTiv4ImmAASm87BWX0lxo9BW/Pj2589+JebYmAtn2/KaXk4d1qH1kIrl/ha0i+AajeE
dI4rK6hq30XGnGyhm8PPF1Np4YNL4QytG6z4gxvybpq2M0CqPLzH7SS0Zqqx/KypcXYzsTfK6VVQ
oYuAou33uuZIsrMBiTxzR735C7kGEOf6830w0YNDf8DvGNBI1w4TYHpcVXUkXkZD8CZb+Hs4HzG9
4uf8HVcHbFnjTQwJT3T7Z3oKUhWtuotDRdH/jtg4XkiRfXImRgj/r9YhMraClTSok5E6GWyx9AsI
k6ioOSeU2JGruNv5vzUwSKa0qmncyXKWleDbYm6T963ll6wYgp8Fn1jswLXQQTl4L9Zty7QFyFa5
LjmoEJ7m8eYy3Ab+BmjuW6+CGZLlKXnIzawBOn5of4+cVgKXfFdQKXCtfb3BHW7VWwrNFGLOiwJf
jXmO54qrTO16NrpqKqRltcqovI7ZSGZzAc+nDRrN6S/U1KJyGP82aR/objg8UZXJQQueGz3p2GbI
1tGYI9913i5eI8b9hmFJ8XdAQVSy5qY4VdQdL7DfTdkPzGSDr8UrkwpDktd9GQjNaPiPBmLmxi2z
RLvwFEFhUXO4ERjABaCeGth7aKoPgBxUvacYagzc7vbsalFv0bzn8MKu0n9vkbEq7ssRbi7dhUFm
wsHxbxrKONZTy6rmHfvjIlJTYUrz70YSWcTc00dHkwkOUeWbSvXwMZ7RGPaNiITCuoAqSTE6+nPi
fq4ONNXVa0JhpZB41A7/Nb11kZEdd3bdkds1bBKzdoRy1FcCnsiBR+KTZUb0/NqopuGn51dEFGWF
jv22R7IEdzbqzZPg7Sp/AO9G+QeJyeHaF1TyBSCyFNyfwoOg6Mr4pZCx3t5qlAl6nvh571c1okMS
EsC9DFu/CqKLOpmknBo8fqJfNG4idLaUy9jL+rbE/JDrtVFMdUJBPFFtYEfVf6B/uSVxcjlfSnF5
x4t7wPcvOApvCGF91i9vKbx4vM1Q20+Acpof6dq5M3lqFQw8Y6mzgXRZvWBsybFAS7o3x+uYtOCK
Mv2JaT8QQ0fOQm2GpiJ5HzTOD6/EiQqrWWoNp5MZZOk+EODoqwxO+T0ufWgMlGIxmSTG8xfMkwPt
WFIo7z31/6nCyN58w2VrBwfaWQugrtSSJDwzcdFqUQRKWPX4JUHZOYD7CqbU/bDfWOVZgfapta+5
0s3z6P/xyVDrgbYvqYR295GnYkMdd1mlJ/hSp/NjJsoGU3sCvSCKL4VLTeXLX9WmgVF6NwK4+76J
obEZmm9Dqyt72mP4FlMuSn5syrifGo7PDOeUCu/xeIYRwQWzW17bCvE+Mnew6xx/JiYdNlftSVVH
nkTtuYT55s0xKE/IWQ+dAsFZg0430zhmAfdG6D0NtLwBFsky/rb62DKF4iSy1XfcnthBhZV9o1uF
MTtKwm7NwzwcPBqTQfin4VbXeAF9mTItPXSuQ5GV3im2NX4xgQdQx+UgG8Zoh4xfXkr/L/RbH0Zg
stkG6VU8cLtOL6Jd3GT+kbhF/hZdF6yA7gZwjHm4B6iHrp0+/OHpKBD+UzGL9p+IedaGlIHg3rFy
8hW+HnnZnujdz3cNRXu+eXaSOfkk/mRwjhDAL3PH5g1dO+k42N2PS7jMatnUUdN36XegnsKnLsg8
UStruW37c5LVyZ1YPabax6u+C+ZDyo8opmtwXRyxBAblYzSfJzDcPuIqgj/Fq6F/wjV4wBG29yEc
FvQBhi8id392CpMLiYyxRbN+odaHGJ7XOjN6JfRFv8c1i/SB68XytIKb4jTfjkao+x4Gi/eECveF
kcWwRPXT2SCTP1bgeQPNxhOhmOo5gBZVmHKRnXLSzUuEQEdIPzEN+1VmISjbMlXjDPTCmyJviGXL
0wrC7FZUMIYCTBaCKgo5XC2GBfy8oqXAgqY9AMPCsYdWF5JP2LgVlmCDs9je0iOb03dGq1nboc9Q
7wVshMGuh48CxHnm1p0N1TEJ9g3cZ1Iw4oPTBv+SaEt+By0MpmUHDfTmCUjh7MSPbo3Sja8GqvEs
2y1rbIhJZrciVszel+oKP7izZrzKCcNoO0jRgL19KV0iiaHXpyQgZz5FrYXiC7k/KygAKTTvUPUh
tkl5GNnj00nyPF5E1LjrFGqd8Iu/ontNV+pyy5g+s1SismESZAlnPcKaTdz2BfLUcP7smJvencrP
24ShZsi3bLbfEvbE/W0s2+XP9KWUDVn9JGQEBrXy8r44rGGxRYJbXdC9gQ69Wa+tS3vHcALqGBVL
fsT8i1KtXJnI9Mp5L5SDuRb+UBD1eMTfVz5VycH99ft+qs5PgTcQGx7aYFjTswAR6zRCylkNc1k6
n0CLw3C6DRu+hBJ4MpV9VJphN2XL3mCEyUAKnxmze1iqfaHS0JoFUUYrJUR1+kMQ7KZLn8DDCLNY
W7QZI18rWOYP0u+xnBLOaPIQq4XT3eseDIFMe2BLOmZCp2wPgtMf9z8fqQIG1wjSBgI6nEYHc53s
hvcL185ZGy9ULfH+B3iOf1knJXOgn8QOq2b+LgO0WbUnF3/0oRBc1PdVHnyluoa/fYWd/JZoXLqA
nJ79GddziZIw5S18i+y+8T9XJqRtRaUxCkwUyDLmQM4cAtoK2BwSdVRXXqFfT+mOhttZfI9nwY07
JHkMgWC8x6TbMlEYEcEc0BnmApahaetXE9t4Jr9s8ULsM0qhxlKEhN2LTrgAEgNXmK1BfgG0aQ7V
8pvyU63GCat22I/+8PFyTdKvtaX/DDx52yra17rsy0P6WHzIz2+NckOj/a6LUwWmQ8m73BXGYhFg
hPhGVYM9GleSlmi5ZqhpzCir7m7EwQduVN38Ve9xrBw/mCdJbIcGkQi+Pf10bYxLz+SHCM68Zybp
czjAmI/eNUgKAo5tI+nHTgUYR6dNXd0LWy58mSwFI974LsSdm0j8LrE6vZcJkzIcmwz61mM0RNrJ
aJlyjxlB0hlOPT5YmEz+n9n3f3nszMLQ4g17eplqI30FGmEaCKTQYRGR7R319qxWI76E/zt8I1XZ
/7kZrgyoN3oaeDvnpbWVfzuy6g7CUQfGJ31XY26ym4bPfEjU1MYLz05O0yFut+Fck9ud4nh74Ica
I4nxvMOzku/H2D40Gp7zHCgjV+LInwOPBxngqsSywgWN740+ymdSnnTJOD/HwiJ4qWTjxeEULE4k
5E3+UIL7hd1uNpSMjt5bmbIM2RNeFoahyJ3o1cGKzVddpxWHuPYAfa4GWDwNDHwooZaSFiw7P9sp
9SKHiD/zvKRKxe2cQj4SnUhpw1nPFAhexEA5Kqzpsyru+gEEIkTbv534uAozeKcVxOTiIrmRtWnE
JlYhu0SCdnbkMAPszXm0jblNsEV+j0DT7lPb0oa08y/a1U3sgDWtK0avCPZig4QFGSpEWSTypWSY
e78K0Gmv6l1FbnQUOdh+ujzXS8wPRtZZs8hqpOkqZ8FlxwQeadGfMFBANWcOLKR+M+7qJ87WFRUD
/6D+LWEc0GNLWc7JAKM7zPGjKifmrWnAGPTxEuAV/SsrozfxJ2ssyU1224/IZvTWKF8fkt/0mCaG
wJ6LkMjMvu/PJP4yu6839A6mPjwqbdWj5qZoWOcV7n0wt1syGAYhOL0jMkTYDcKtqR49TiECL0iT
c6c+DKvYVV0zp6c5x2HPR0C8EYmaFQEnTzdOhSa3O8BUVyhmolZl9w6fb1I5sFUt/vLEzqBfGCkr
B25E2FieYk/u6s+CwdDla4oaHraSQJycVUSorlFts6smP7/9ieiYiQ3iqCM73s9vxpFw6PNninrf
8MNF9UIhJOvmcIiEi5uA4/YksmdVjqf+FHitoRvU89H27gslzvEpmAqFUiOWSIW9QfiP+fp6b8Mg
HDq5icGjuPWwsLetbsrs4TCBLjdON8DdyXwMyd4OYZkHaySHIqx4pOXri7cV7bQwlZRvuC9lUVha
nGhTYscW+ZbQWR+eF7X5klMPNQNp0227OdyMNz18PYn3jCCJK3KudqlRbitywodMh3FapY2OcJ6E
CUDwXh9tkWuE7nLdD27rorHxJgal7tshA/Zdd97mh2vg29IYCuAfVVo4TC504B7Nkvu98Y8TWdbn
p31KOJVW8T9xxhpzACaBDPF2vgM2Hvik2VLFZEUzAJh44J+O4zmnKIk5L/Qtd0vSZ/+fyci8jLvA
G9LGffGQ/lurqanPrY+ObXWvp+iiOlC/NZDtwwKk1XEAInySFxWI5K/74Z1FzQuqonLfgvPaUQxW
yBeZzcNFniDsnTJpI0tYau4t+JoY7z7TipdgUTbbizhiMACcVtmElXwnuGVsTN0NmR6y1n3Zr16T
3u0KUkoMNAHj1QIG5nuuvmqHjmF9ocTtsEgIVC9NqBvVw1z30QEJfwX5EtbIIDf9bTVN9u6YSyAV
OnNqCNp2ZiYCiXqk840CfPEI96VCL4itv4X8zfmwKvW8Df0uf6VfBV6FtIanwaBrEU5Iz9dlA6ea
ogubHs88ex1sCQaPXv0y2emQxQwErgz5fcB6ua6nZuwaFQPEBB6305vduKvL5jZD9phXL19tdnMw
qV9F+RQYjMlMB06odUiP7hTFxYirUz3uPMC8JXXKmQ0MJTk/jphdDSGQgMgxkbKgmeTwcnKZhy+p
LkSRDySqRlb7gJtayJHjE0NhqJTtIbhvmSTxfihtAvPpwUckfEbzdKZBdlHEOBY5n/HX73kQGkKT
F3HdEc/AohewZBv9iMYIkAtujOQFCS9PKlJjht02G0TUi2DTF3BT0XAdhYdMqgpwmrFDlBDPHwXB
+ACaGHw//B4SLHSms+LCY2K4hEvincTNhtch0dCXJ3vwCvrNzzgTMd/QlAfMt+ggkgjKGwBiF9o5
JBzjKw5Q5Z0R2RPORI0Aq+FydDwKYs+vkpghw1vVSseN0XrD4EGJ1oEUkA+HM47Y5pNr7HTBpQ29
7vmUgGMXpV1BjiQ23rA02NlyFT+OK+CRKaAdZBWSvty6lkQcOYQs45CxZtF2PXPV6sRewNog5bXV
WYnJ0Rqz9rnOTe9BUUY5XHpMV9nAjrgxJ1SPSsAX2K2FOvhFgaQN1Aon1BoQUjSXHjd7fZ/lDeXJ
WQkuVm5gi3p0tncLbL33KRdWaASYBfRfo8px4ed4/Oq4eDk9Ifk3T2NXT3ynlz7F0un52czavTUJ
/HoTrRkjb1DMHkNCcN3lBuLc5+ZSCAqKDwfK3c2EgFcugDz9BMOJ27anjpynmdbt7qOUZGVAeBgf
UCEXEyOBhMWcZ+n5aZE8bQnfqjTuNwJ2NYJVRBxDAVFUU75OIea/OEVzjxKSC7xkWVV4yiTWbBvC
ZwWLQi/f9r9kKRo0Ult8IMKr1lxlBv8/VgUV4D1TjWpLR22Pfncg5PyxucpHZw0n+jhTNZZpY8iw
8AjyTFZEtQcgdbSAuOA96op/xi5EIDdWNUgsHYE7Bxis9wuXg16zklvBrThd2Awhj0Fpv70pXA61
zI7mz6f20qg55gZHhrVS49jF2JAnSDNdZSxn3ki5a7/Lo54V9E8U2aRHkShqa66ChnFVgRdJbP1v
sZgbMc0ofFqC7Zs0DBAWYHM2xYkr3tJ0ZEaUvsXowpTRUVOIWk8YQoBBPi+2ziToRjtTxHCmOPU4
/Q+OalDtYH9w85E8bDr0ZpyGJb0prQ+YCSHusIn8sQRlUO3AiwMO0QucuYTIOPrwG8Q9iuGWOLoT
bVi5x7/ujOlMAYQqoBapaum4w8Jg0u8EWJ3EPHr+4NmuyLTDVMWK2ll4jdiI9Qt/bA0D8NMXUvBy
gh6MaIo1qfyND+IVIR7gO5Ncvco/ko4sFg2YjgE/YR5mfI/9YI7AstKrwT9wLeFhZ+dOlLQHtFqV
mzkr17CMZP7k6CehAYUmQNFuiLEWds5TvKBaKJhZdBpPnaL/BR7K7fGSQanXDkXYBJN786FTNwxK
+a11t5RLxoBOn8dGCTGXYtF4LNSACEi+hG89GqBHMzrgaMn//LpHWgl7nQ1BiqcsF0MyTt+c25yY
93a4g1vDi72Wuh7UctgYB46HtSQjNVvPARZ4mHlflVNnqbNXjp8YHPV8ZHl1B+QLvX19c4H9AXXq
fbAJjRahYjOYVxM4EQTC6ompudM7X9GrPt4elGpPgHftkfffKtdMTzvLngWCCY5ZT3RAuH/Rs/qV
/xeGBtwe5WbPjZyTuUexsQ6BukzduSDIU39o3mqz9PZMxB2h4p7RHTqvfajibnLAkKccKmt4ZWhI
+rIkcXoetmhqYqkEgXeQoLVqaG7Y6BNvP+3KLvYXfI8zIDT1UrxtC8Us2pADu5Mowiolq5BG8YTA
j1sUey/QNlbfD/G41XbeE8A5xlUbD44wMvLKCrbKkDSUbc7lYzWPYIZok64rG0fCdUGlElVCTLzI
16SGiGVNTXWHpgJudG+O3l8LqADxyQodJKnIx3IeZZ9vAwJBdXdvKLmOShv2360byqd5XrcrssWE
kP6gQk+WM66KvJlbdv9KAHk20ut9qOTNX5SNaayUS2oeznu97ctk0lDdS+FFJFdXUEh79m94QdT8
arZoiOox4/HhLTs/TldoFZ/FaeFmZXNW/iWomudBQkRKnWCtJjenGqxNRclRTcLbLKv22RA+Dltf
RpeXKQlJ9kj86QfIqHszZwK7uDvRdFX9EYbGJfSdKj13fPPJI1L8aQVjkzCjlRtflOyNhkDHz/hw
I1clj2Z3US6qYrOUKnf2c3TvBAqLv8o/GTMUo4qUsEKa5pVsLF/9BC7965I8dsIn2vzqQwIV3O47
aN8b2XRgKuNCnymOrIrCoMsWeSXZOGkttH21tMf0yEBp+t+WUHnOMwE9himWW8Ret4tf8+0y5irK
acO1FNNl/bjnNP930WDp/wYAqgqDKDbmSTi1LFyzZbbQVe9oy/BNcMJ1e1RntIa3I51trjQ9arIX
j3S+8wMLCT4kSec6U0+RmsF4VvKYyZXJuPkmhZcw4FyCrRAB/65BWOCnaMtp5KX9QkbSjZsIVGlT
6GPVAwfDwzfaej7BpttcY+pczEz6ewo6ppmMRfJPgTFCge1rDdTi2sVGjYKSXmwYghuT543yOPF9
ueyn/0Cb/sbc4mIBGFZ/6KEGsFvKeL9k+X1+ASctEYb6UUFj83FFnAtJPxiuLkvGgEkQ/jqlAMI0
mFCCaZnljeWgYn7ohIO8uFApvNSlNoGmkP7iNnc/PZmw/TZGQ9x7pTFLUvp7Q3raRq31wBnVtCv6
ElLrjpPFmKiBB1o+Jxx1lr/kXBqzD3pmh6iQ3998xhZZtovfI8dmtUrVO32maTn4Ji/snEa/U51J
puLIiBH2k0Z46EzOiggDp25iuEaADThaZBjyx3eSQv7HUtVTd0al0Ao123BwVJ0EjHIbPZllo3dj
7MIlW7uXrPMQzA7ZyRXLj9n0bYWQVlpounsDWQxDrSUhmZADqKmoE3WlVXAGyPUASLUQ5Jd96fs7
Zssz0YcS0+1AwbJSDDHFrQorNZCsE03UumVgzlgkQ0EKL/TBbOj88ULqsDq1cvBhPCthxr2aNOSH
aIwnhrqiEDewLKd/qFv6wFQJCtTKgRnep/Hi4vxqOkjWkAY2mI0eMhd6K5R2D7ZpOTyjUG1GB/nb
7+IoxV7DzCyVZEfzxy7LG1fo5n8E9k/kLdBXhr7aDl6OFkvHc1Vh/ruwBYPrh4oo/E3C3bZRo9ch
d7Aq/3fn6Tpq8mF5AJgW4Y5W4HVNamDk8z7ON8Ef6aFb+GZgkoAgNkCgvfCMa2Lm0jFkLcJGLa68
wkZxMfUMAMnSz61FKAhT2AKc3fESxVkpN4oTxDF3T7zcM2jRJX+1iJWEcuuOSGqyi3chfLFkMt12
byCgLcBzXocwCn6oTugHUdFs8RxtTPj9QZHigwYx+3EmvWyySyNNU6k57RU78+BMH/lfQoSFSCGu
uyQ07e8V9dba2IBDsHU+49T3k/Gtu18e8Qa/xcescd12eLpt+aFvTe3oos7RWvKq9QczQOxX0EqO
2dWIT/WoOx7gNsgdiVAcYhgfoC/ujjS26gkdZklPhfsg+TlfTpa8WOADmneabfjLcnTUDf7Zk1WN
GAHPbhswugSCO8QhjXpgzhaDNWZqWYQW6dwReqAH/Ka+wunjhEx2FQ8OriD59MRSHW8pZXfjCUoe
jQmzd6qld1fQpeiOCec08YROCi8hQxjmVg+2eqOBuGlrdJ3JPldlOE/NGtco4UxMia/TTau6+EZk
Ek+HWCL2zTtTF9hwDawemc2QF22qmYQlv37BpLD/ObQ4VMHqQmoDPaUFXWBRDKHRRCcO0Y40iFdz
wIZMn4AFDl4ZBdnEnhnjB/8e7uXdZlR++X17nafz8+8W+m701B1buUQwOjnzS0oowIk79/wV7EQe
XJQ28vuC9BjdDUr7z4l7iJ8l0ExiElTX/0J36RJvFuCtJ3F/h3Ozei3WzWMCv8dEnpVExSz1jQbM
BdwwovEL2eM2wpC0gmZG/2xn8EkIVgM2GXc0npjT3zfIWNGynsDNRcv+JhOysBWNt8bgR5I0HZJW
pOGesiCV/I2r8fZbi/o7THAx2vHugtxlTYbrJglMTW/GtRWFuqL6bxaG3v7JYjEMJwnjTVUqANND
6SD921KkKSTygKGXeGjaxy4MIz8wsC4ICYVtMmFWu7wxAA2egjlU2rVJWdPgliY4m92Ao46jJln4
gejUqe0f/V7XyfHYBgUheAHfZLYtA2kKBvndP/Zcn2APCn+7LKdNmZndZIitoKyjXKjRd19QqtMn
WEDtbcG6OQ+Nujh56rw/NW9p2r4itWIyMrOXE4rrBotbPb7oXd3GtutjNHlxPwH5Bhb282lOOTD8
F4rokXY9k9T450eR3Ma15LdXyca1So6p7RY3dbznmKTd2z8mFHPb4mXKa5+dkKYYS50iBrRrAK0B
how3O/umcYIC4jOATNci3DO8C5z6a54zggFOzAUaC2t9fM7HUGaI33JSJr1RnWWRRroiSh8R3YnX
K/G7tiEJfqLqO4yi3CXn463G1oaUtTqRmkjgMwEWHhSbbKNuXeLxysr62WWWk9mybl7g15kOsCkL
Fz68cGl5+UoPme2xU4zVxIc3ifKnIoJRhIh8ZjBCeTh8XG6I3plNrfm3myKQ6p68D0J8iGcVCJMF
uyIMjNwFcSKHY2apI8OVnpyuL04EJ9lrPlDQam1MSHKTnNsIGXaqjh+iu7H6jla9LrMpMpqXIHWe
nKADG58nlatb2tUNo+T7GWuEVHVCk89ldXr5+tq5iimDmRjvMPfp8f2gXdAHzETZjgR5+SrPszP0
BK0EirLPuBaTYT9n6XRfZ+4LcLd2OsL7i5SxMK5+XSDGeyvTpI83A2Jkwsgx74hRzKv1hb5uhcmx
8ZmN6zcRqXH/yT7XNETpMmLgbBiNfkXqrJe8EpUsnMaUxiNmpgPQGG4VagBeBEh8NPP9H0KSo/Kx
JLXm/GzUuDPZIl3IxXM+zeTzPpgdm5SuRRQp49AHAnczDYNkzj8FQGtPvB0meH5hNwKJLwQVMrM/
lW3DDZtqWUD2YiaO1cL9Kjb0X/IHYhQTw4DZXe1qrgiLdXKyHns7Ygy+eRK/DhEFOkPIdKM4QOfH
M7brQWfsyIsx1uUtVUhHBvBfRX+idsOi/OXUYpOBlyHc4QAl88d6P5Bg+hLf58jKozpqZ4lxQmyE
XjXIdCHrLGDjUqIGEStypdvUtMvw6FyZOopKCrzNa6MpWQx1iXobAEdFojk+GrcVDZIolfQeuGc1
xNp/RyB2wzf8UWN8DYGjcwJ13eGl3h7dfMAZ2KLz8UVCy6v6oIX7Uv7pswf60uJNW3oVa5aFX6jP
1Ze0x/S9845ef/zIbd2iGoGyN5w+Qz5bV9t/o9Gaeh8QhfY8ajlctbySmoLa9Ihofa8zX7BcS4wi
eReRN6sLu+96exfYFSvdx3Ws5yHV7Ogfc90nCshsNzIewf8jVGUIsts+3Bb0IP2DSGSWJnMg2b2y
bIp/elky+U9AqnSRWjTrjusJTOFhf1Fw5J/2gJHqyMta8QM4Xj/8hCS+mxJomM4Gs3FF8Q4e32Dv
92VvzBp7kY4OJ7yf09jiYQqtMp/nhD8ANk3YK6FnTpbt+e1J07SI8y3+H9vS3tJLLKIYwvKS9eNX
4umKYudfBmoV8rlNqC1ku6Gqysc6EZ/fRw9u3nQZt8asoZSh0+z6Wp5idW9gyy4uUCsppS54w50z
ABV4YGpytfONmfez0jbhuHIPmrle0QO5aw5sgRFCnJTiy7pnts0/PDEBXcwxvtVQvj969eJ8BSZQ
6Ta/D7pCQLIlM0PGUfD++uC6T95C7gFBVAJp03ggDT6zOjnPEp/6PFtZKEQgwYUWkPxur7bBudRk
4ojdrDzTH3FBvH72ycC7sBXP/GI0D7GKmd5T9c33+R34hzrrPEmn/CXnpl0WXqJ54KVDZOPXgvae
r/S0eQJg6JIjGWZiaFgLIy1SbPHTUyXL8ure3aWuJlzQmutysQcXo8GXlubbf2XkJ0lmEhKPzy1h
kLgqV5/nKEy4613YL+lnj53CaUjNg2uSd01kb2O4ArLs1ZG7nsq8JOf3kPVDXNzfZt8Df8DuaZvx
pOznl+D2ZyUhuPVCMq3EzlpA5x2nNwmjpGppAnrTOYSmLuB+YfPL4gn8X8XuoIMdo6P5itzKdmu1
tsWd64ksy6TNvFhqQlYOTYMMSGganNlj8t4nLdTXyEjdWv9M8wu2+LAV5xslU2AxTJ216reNTsN/
SvexsIZ5DcEH4S3QAlzr4UmtNewXPtsYQB60yjv0osPMDdiH6uqx98BHZr0TW+uK6raLvB10lEzt
s5+f7/KcNJ6jZN4NLuIK6cDTR9+rXjzXhwtWkv3hdMvLIoSwILpna/WUpuOsvS/ofVk4TbyQC0xr
kyguIIK0XSkQXarylK1ifKdmfm+W6NJxjB2hIuvKj41/vJkrWIH0Mm6aTJWKzgN/VAGBaKVhJIJP
gZA199wKw1ZEbsemYjw9o705Jr0IC1o7eqzDbQLjDS4x+7f29CyojzGw7M3x7JnvmvQUXCJ2ExuC
Tr95wxpB8k/zcGLVjcNJ/QIl77Gejg6lW+Ff/y4HkL81plCWzcuHWwjImtsmXz3RoV9C6eHeSinq
1XStG43aozkowI+kw7GnAHbefxRXzweHVQVbGtBk6Tnc79Mk8MrEMp9EhaBgusbDYunLepbReIx4
XdSgvyEcsIxnWFMWb0HcZGtTP/oyHDkvZx0iAmstCjBlDHxPHlQrUv8ADNUq9LKQMUhpReWFrEYt
uS1yBuBFkA3V7P5WiK7I+8TZQWbLT/M7kJZTqJXyHT3gnK+xT657kj7gz2sX02YrEKMtFOHSBGl0
voeCUhTmRt0WGj6EOa+otx6laY9j+ui6m5tQmcKEFtKnOHxVol4Ic+RB6nB2gWfyGzTkSkzPLkTC
agoA4XffdQ8NQSeCBVYrbvqSA+ihnO7JfXpNc0+2CjmT3Hu2UREJ0iBHvUtxD0orq7PT1s7uhO4X
Wuz0TpwPabW6SYmQYSdSSRNHkJ9WESqmzsBYL3moieZ06M/tsuJM6MKtABP6CGqflSNwdl3cNFAg
5OKyoXAnCFibPi5AUVxnBt2H3SiyDyH08eh0yq6fwOtL8gW6djy5nFsBFoyOIuivjMUjLba5lavL
GcNbNrZihR+1KkN2MOtrpPArettHF4zTpNqNdYKHnI+59Y8eTLZREkDG6gywBlMwfJHr1zq+Qncp
90TGvMk4WUYgNqG5ZYHMcj1R9Oq8nqwkA7AJ6ZTmDe8+3P1+ZxRNNj7owPJ+Epgowig9CHfKCH8I
2xNRCBTiqF+aCMwf38gU0a1HKA6f2cWsH9H0vFGKDH6Ile1tw8kUrv1q8xCcUSv1FsDD+8FiIJKT
vLfZZWA+1/rsQ+fEt363snNHSOYNXrLUp6jKVmRfrrrBOcS9Sb8JpKfGUFWG5pLxctg34kX+wLuq
m/IA3Nb+rgWllVPVDef107Yii5KEaHrJF+Djb/2rEXZ6YzzI0rCqcdNLPh8rJAjmPV3NB8xK38k9
Tr88CLIx88vkh64kzY8m9zZdXm+OmygK+9KGv5J3GtgyLCYnvz70GPRZu/7jgyX6OA2e4nUg2gXd
nB8/Uo13oCYpVV5yDMblKPwK7Gr596GeRSAf/bNhHvtFx7ILW+qZDxWJtHtEDhdF5VVlT3bIqrVS
dWzqbJ9Am1dYSb8SbTcqyluKmub7W0CV/o/3/b42wOe/co2iS+Vz/UXaYk4KM6UxEry5C6njdgT4
IJ/t3JF7ul/Mrw0l99bzfhNbgkEZ1iakEQUYdGAzRCi976//QRpuBvi8Jx+s0HpGGff1MqsE+1VQ
xtLfJZWOkFRMpZOPb9q7v24awkSBsuFbwbhCxhQG9xyUVmwNzqwnfVrQI4+6OS5ZYgNv8S43vfby
tWFEuyKlFJ/OGrid07iXCG/6P1EagN7ZpIKsDlDOm7P2B9gGIrOLgct2mngSro9TWvjORIfvR5uy
fkQcx63Ki4bhl5/0ca4N/QXt4cZ+Nuh5MnUz+cH/14bmyE48wyhtmri/2+WqQ5FNfi9Bq6encFnq
j22h5IJezMtOv/FYWvIP3psCWDRRGws3xgzQKNCe7YjGbBqrvicPI62RtVLsZpgjHSJvTorq4h1F
U5TwfpDOLWYmk/5sRUHNUGd/ErIRlmHDCP4Xn6fbWqitt2tx4NgEXMmW/jr/d6PQ+WjUYlmGSuJW
s5urBH55y+vjVol5pTbygUf7AES01wXG3qES1XGBOJH9PWH0Gc03VoRM02w9VV4+3Sgoc9Mfrx4l
H0u92hPcN/iBW9vFGg31fyB6e1RROnSbtCUQRv9UMiwWWPCC1FJVoEaID4qIMP7/9vH6qv1twfDU
DpknlHAGca1kzvJLgTIuNToo0iCHW9D+JHoNxXjkBVNn3gMEKKIB+kk0O4Y+9a+0IifAC45hUs0i
yjedZVj7o6zZIv/1VQi5z5jA58QW23z6eP3Jx8nfw/nVuyvzFQawlmPdqD6o5WfbJjZauEoNuMLs
Fq8mIsRmMBW+aGkHvlJuX9mb9mSk7Ctsj9AVCNRs689sQzcwWljA2ckUGNEvf7WJnmZGXxYkDUOI
Az9m5Z/D8zsaBElJaDi7iXGnjn4shzA9pgYZ+k5ZJrRjCIPdpscbP5Act8n+2+VfJskXJYtOUqfA
OYw2cl8uRIzIRJYy8jm0VNeEFCI1Y57S5UxsakNnfNz1v3Gb4tdEu6GDVlniK7rJlXD2+DoYGF7o
o4uOEOstzZqfT1cf208ooRacRUB2MRc1AB9sM4evgpxOrxGWcBnes0fAsy4PeYhLSp1WwGNFX3MV
Ohhm3z3Pjia0JT0Zi+yHt2lmwHGtRb3DGzvf4WQEtSMs4XBbQmZEQ58b0MgKOwlIJ1VfgYM+Xi7m
X+jSdUo3ozh7rOYj9GAqcs/rdEYO3fa0h9OiQfAizawEsyTKzyYEqpxoHgL/B6yLShxv96HmLDSZ
2lI+kl8VnR4GxkStlBG08wCLCAvThEivUILFHq9MFwOis2ImZQENhBl41k7NblWjNT1xPy5m5f6x
ngdgAA74LMph546/blHfr/1pkFrsJZZ65ShANYf6+saUen+ndyPLSJMKRXbVPCDYomaQLoBFNU2w
KeghOb41mdBUrQ7W75IU/9+vJ068oXh+pVDC9QD3wV/Xbnh+3svykAjex97+nrNJLNThMDeaj9PN
qyVUn4NRM/T4JkDIsO5dTk7ZiJrHVoZBchLR50RLxSpnDy/nwLJYkHn4JAKODiILZL40Q3aGT+rm
ZFgYdyFrKZ2ciuFsUTCvjNTTiTHEt9ru09BRVM67D4OAhGRQtvwuSdEVL4Hs2fyQzs+A/uOd3YLl
40NNF37dnzm43N9ABQoA+nSh9i8nr/EXqG4/Iwt0X7PvlR94o8a0Kc0EG5rzTbJVX8P8Qnb3WKOz
FSpfB1F/XdejugN8ri9JQBN3KeVxhb5TY8+v+h7gfhitl4vGTOdSOFkgth4FnYLxhCNAjHmnkt2p
Zq1Xv1cPuYpCft++Z54IsUHuNR7AkjIEYFtx1r4e/w4fCIcRkJSFUYGGQsXukRPGHBbo8v8J2oaE
1VV0Di7VY8oBg5Ew3QsTUJLvY70HGlWHxliy0hOr0vqM3zLayJmYxGWKCQUPmBVUHUI1g8XWhNPI
X88o33HLDwX20e+h0v+kBjzKGFLp0MdK5uTxb4Ecb5GA++OzjlfQTZQCWOhFentz1ZWxwUuriOhu
7zFL5qHwxR/QxiiPTUOERy6w54a/W+LRoASUolM+kRwgdZIibb0TAL2Rb8BSWDGnj37dtBXYY7dQ
GIIEn4iUoVbFJurOpb5ckZNzqJXfb4BhCIqFSj3XpOUOY/zU9Vtu2WOYM5BFPVtlX1aiC3Fm+apt
yR9SPxYlGrowMJnIH9HCSKEb/74lscjj9xrd2qbDhdh4MwRrCupWiKiYrvwDxxpSnVzOjiX7mxwz
NcfwMCrUxFdnPvmj0brCFy40/zn4KXXiwK1GATvZG2g5fPffWzKp/pALfbPNEtD+9N950ejbmRwD
WJ0Grja+mI4+KmmiQctpMhDeD6KJ7cf3CLucQKWptGnmcbwGq9Xi9QFBlcinoKXzaoBr+p6oXJ+4
R2h1xFHuO9HmvLwsQSv+nXF0kSlw/qY1bFze5eYN5PNnPSu5aH+NAl/KVDLHud7grcnlMsoY3gEn
sp3t08tflvjEC/Z6GfgTUrLMPY1s3ygPiP5UjSMtGm/pKJoTADLCzoyq+2kT2WR0sN6YZdGDQndL
apcDH3OxwUFs3SG4D9DGYKLEC0Kn5hAnz2Ux9+xkcnIZKXGYJION/BKgtRTiGwHIXqLrnKqfWejK
8x9gN4/VazeZYjB4TGp0lU3F2VcGfgwMNKAIYGMskb33OajVp/FkH2Zf55SUG/t8D3kZGvIjWF+K
dufWHMxnxZrkMMp47s6+E6p5Kd6Dv+bM6k6NxfQEKO22jysK8JMA7YaMuZuCwucqw5YQc75xcupF
tF3nXzr5jOcpUHnfF1SJOmq0ROJfOdt2siFCRKR+40rAZy9tWw3xel84gNcIAsuC/Af7vvLK+klL
Hz9pbvVyZhVYnwmzYF0UK+MOeszg2xtvtRrZV8Ch0sjHBoU+nMoXvWrM3XAjFNdW4+LeUGiXYYQF
45Q/Ar7ViOM9bGzhyV//mRQHfHvdInnDJB+Ww3BZjXaGaQKy5r8V0VpPL2UVT3Z9aUkvx+vfHQMh
Bx5YzURt93orq+PWn9RfvoxUk5wRq8YNMWkY2KucBNSKCcP2cO5hpwS0FHpklhmwrXIc0gCH12ym
9EYDaZGpqQjw9vVdxTWbMTdpi+5C63oaVScQUjsRHk5whTaiCqYa3A/T8mWCHpIHkmLNa8va/Y7R
eDE3I5ZdpZTPhIN857biVovGC9M1yt3FgbQwAh5llTQ5e/wcupcLzOgiPTP4BbCEN/hKO5JzfTsy
EcH6Fv+0zlYVU6mFUqfW9pQlB8fvrQFqJbZQ7z9vohsMcO94iRfOfiYmh5UPPK7gss3qMwfYSDRl
NJz7xKi7TOhOTBbxcYBWAQeke+2mo+qkkd6/sfAN5zCh8gajYbChtPtpT3aOvJ9y6KMVRkhf/5ms
ZmGYvZJTkA7IFumrrZZldZtRycDTT7Y9bkrwM7/WK9AoIPAil5fUrUOVOm97dGJLK4o48DYewPSB
Qzv7ccBiU9CZo3BThtwZmf8EVUPaFKWiZvHll9Nfzj1RMxqND1uu6epKAmrMJ0hkcljOUiWrF5Az
qAwXBBQ2tv2UooK7Eywn6ehPsOdNsoI9tZ6/uE4hEBIjNkhCBjNU0K/s6S0HDrT2LyWi4MjAmyZ9
mt2iI9POsEhiOmFCGfAbMxvEpc21K5knJhE8n5i8M9SMqKCik004YEBf91KbO4vEJmDCS6t+aSyk
fNwJHvcGMY5dPKBL94DByq21whHM0ZsXeH8QTq790g0L5A28pFObalFGcggCLO8EiABgoadKu0Vh
Yi2PslxCJZJreI1FZrRWcJKVFvISH4CZ5Dbv/VKIuW4slLJnmX1OlwLLtNF15Zlddl9fNlQaX3wD
ukZVXAfl9NKV9AgrFSqvGhz+h5uoxwhL10sN4baNLhup2iwJou0Z2j/OW92INPDayZ0FDShupz+I
XaLec5ZBSOedDH9QZw79dUI1SEyeAi1DbjFWV+YnAaf4W/ECn8e62jA/v+VO053CxY7/Kci2H1K8
PMb4r6TSPI9hnmWpyo1FLAeCBfygHmTkY5OHu+QS7uA0laPu0BvTZTFvjdRfjE+Ff4G6XKDDHCF4
FdIq7qEixPdCUMxq3n6yZ3kL/UNv7pw86mRAhpUyd1kbqayHzbFw06kZx1vHGcjDbSIMJApeI3cD
l9g2k6kq5Qy3CFOG5KlI1y5bQOiniSwtaS6dqZP8z2ZA9xI2+kDOgovGNBsQa9guYzgeOERSrnxb
ktR2jQ3OZ96lwbGAaf4cvmWfL00bfgj4V6A7I7Lc89UgIrEcGB8khD3KJL+IuweV/OjIjHsADyxI
iZvtwdYS03TSUuqRbRuJziX051/AJMkj20l/SpXRYMgM/XCww/q7h/K3J9YIVfThSJvM7EENzRru
gW4N+fxDZn02DJaHknJ69JbOulvMYbJXXwagYvlcvgaOJE0I+jIgnyOYY1QvAVgwaD1qjuq+WZUc
HNgOoX+PlNh9uS3bKKJYoZSA7kwvXDDl00WjJnrbGWcH80eGU8C55lSV9DRiypGkrzwOZzsEsgAH
yEJoZJLXGNyxWALGd6RI6qIl6m4SufGYlHvGxxKfnsZRT2g199D4X+KYdeoo39ZGbnEVDCpbz/Cp
XPtyaQZ9s1H3kJp5YQHWcnIpsT0O5/gQ/XZodeMc1fjwC9Wn3+SHK2c/6pkk8ZCUcvkoDLe3SxyV
mDKBqNc5zDMllOj4GXv/Q6Bvg+yyUO/S/ANrHUl3idLgD+F1c384L0AaEKA34N7LSoRzy9UeKjqc
qRaL34XLmY6MOkSurz8eijRd3IDFM24znau04SqYasZ6LCNtaXTDmR7ypvtg+v7N55O/5k4Ot8Qi
FH/HmBdlN0F4sHg/wbzR7h5Wg80wqsHE6FjN5F8i3OMl0lHiyQjJB9YGiYbSOZJS0V7p0JZulryr
b0EAr9V3+agOexwyz6HqWl01rcAtQpx+Z+DLNyCnKwwyecRifNwkomhAPst0lzjDMcRIF1MXlOvU
1BFm/yCS/rfZLBZHvYeqxePIdRguFX6nGllQP/9WXHzX32GxCvGkoVC/aR3AwGnjII1zP+GFQ/j9
ziG4TQt55O6JMTcyF47eHvJWyEck7b5XZbLA48Bdt1DmY17lOjbVNTVJdPpP2XaZpC6UsO5J6cds
Svj6jPSCp07LQrxNpRbCSrWxvRxZEjLYkhIJvqn2YJbmW4H9nTjkZcwG1vVS7eP5BDRms3Re7Ysr
XcjNX4Jth6ujt1s9RBNzS6HoUEo/4/5r64VuXKtCizrlVW/GUFLWHJdYaMtePTdssFjIzv2Dd7zG
63c9kvxerrXZDrEOuUyD33OM7POdsWNZhbo7D3JAhMKnrdUCui3NUlJkmBAZx1/m41EcA9m5Djoy
heItcmYqNTYWryCKcD8tBXY3efKN851yyQBAUIYjcWCN7a9oKpQP7O2YaTg6EHsQ8q3530C8bJTX
iWLDJdVWN5JZJR69+RgPsfrXEoOTDUXrjBK4jS1JrXLCkUpvEhQ/cYV0KQcuB5xUyOY/DY9pX1B9
XkTehCLBywaufmJ/tTFTH01T3vGUEwcuWTjTuBoAk1goOXycKcGQ6ugiLSClzbQYT0t/txBk6Fp4
JZZ6BwRtkmA+l9ciqM/twT6olkIYaf3K97hEfbCFSXplGh5PT69iC0EjQWVmXnAvTqiWG49ny3Lt
v5u9vIqDyPstnuALyfKLrJMyPNz8Hd69eMWs3l5rNiE5iJUBVyzZMYspXDNyiYUBiChM790yHhay
3azo44IM9EJpUeC1uJTHkxhln8GAt4xeBfqVoqKTNP/darnz0ypxxRS+v2/zSdZ2ZmKdWigtFT4o
2QfkGefxvViHUtzdJxt/c/NDO2l+wRkipIf1Ym7x0bPDpuVIjPG7bCuROqgIGRWSG2pOS+mtIK1z
RXkSDpeXuT76yswdYx7baand6gh8Vxbt54US2W8s/BF04OuKfoZ1AgZDTzmgqL6mbtUzlww7cQgM
azs2gaqjK0udYpsIKqwIhRy1hr1Or0t/JAoFRN/x557+QQnXQ3ivp4E/A+j93zhBfEpsI5mRHb0q
QEfSy9ALzaknAlWcQiJsXNqX7lphIn+z+8c7SnSQHu2ph2uvtfSNUfjOY48LIkALEpdnnO/cZC3j
jDVy2XeyEZP3yxMTVeiGWCNbw7W8l/rKV3NqwGHtvPP0oHYPbKNFcdwr2RCm4voTrWmkfo0U+e8L
hK/Q20QjJ4YQuCvJ4wb7pGhj60gKZW/YYD6w7Xl6CcBF8lla9ARqgJjKjk9AYr5Qp+WoVOKE95P2
+2Skco1PW9bp7U79AWQ7NhjyCiKSIAwV0EhvB3PURvQwR/Gryc7XLw0pZupMJzb9tNT+2ci8oui5
/1ugPPfgiaGxMbdDlBx8YagtHBj5pvEfLNWIGlnefwi4T5RmKsUE2CiBUBlNtoXOCIjM50+1Of7n
KvkM2kYsAjj0IGVE17V2Igg+ii4UUvFG2vD8mRN1Wmg+xlS8ihd6wITiWWJ/LkPDjdJb38O7GXKs
uglsDhIKp5qvEyjpTE+2a1xp4Nm0NXp6C1W7M2cwCw5qC7RHU4nFgaf2ocSh5FvQz4v/ZJYC4acJ
LV+ltwSD3TPi3fwYNRYuvPySNi0QIPqa3czUu9BM4O2llDGt2MUqpLf3ZgTI/5LTKGrCU/A02Xqi
+V8u2Gh+mRtiv4BEyQ4bAwF16ZKE4ETeCTIgPviMREV2QPSLfvqJYOOB30EeGl5XCBQjvab+42jP
tDsp0w2pT28mz+Ioch3wp9A3sOku6t+JkSuN+vpanJyXZGq/Lnny7YhRCTmSrPmhURONVIhSCSoe
DAsPSvQeDSxv8iZAJ7fz/XTE9jwjLFCzi7DF6DRBfsimNkDxQBaLq8ZsfHVExrCbr2pPnF97+FS3
dPuIbXk/s6g6oD+FmIXkQy3BAApjYpE6jR3Mm4dQ2vef15YCQ3WMg6Ct6lsZwJf2M78SSKhc4mGL
sT23ySOsi4JyRrqy50wYRx0RwSzOjVK2IXbz+FMQvK3Pz2QcewGd65Ag1KpWTsyz8EVrpzLliEDe
7hgKSRf247vhnSs3ENogKWRru9daKdC8ieJAN3Z717fvq3J0o/nl2uJhZbO59rdl0AEJz95SaKHT
FFbzPPSwqmShoH2XpOKmqBCSFJmAVjYJ9pkVZXuR2eeP4uuGHuLWV4/92Hwku20g6neF1VqbUAbA
+ST3vY8Jjgkh9lPizzoAU8ggNAvwvwV2XFFmvIm90SB57Uf7Ry+KujTOJz9RFrrfzWRWYZsDntRz
+JZaommGDrYmJsVjN0n7CQ+fWkeDsx6sz7q1H72Zts1TGSfrOxKEM3eFypuqi+yHzCGLydH7igNw
0MG6mWuj1kFPS1OPtpt6fo8347ccFnY20llHFnxt9Y4UfKCx+fsDD67Upid5OW5NGLoR9mYEX23y
xkCpxlW7kkYsckLxPM/+aRS7Va+dyk/X8CN8EE3YAwvo0Sae7Kx8tHBzWR4r+Xk9y/D85wgwtYJ+
5Ijkyuvcg6OY11lNVQiLoCmhHv69w68V4h+GBcE10q0tqUVMAXk/tCiFzbI7UOODQiMizHkdJrm6
QaalmiGMpRVINpMGmAw5a0IzCiLM3HPuB1sKqv96mUkMB5ABsK65+SW8XsHRCpEw9vbZsPO85+0T
Hhh4TlPQohqtkCBKZJmMFcaCUopskvhPTNkvv9osaXWPurSxeJCmyYpHe0JOdRbOEsAdugWjOMgu
0JEYmTG/hG2hhzwIO0yk/+p59SgPxIwa/+awFV0mKSW1sfDX1dTAcVIuFEbQOsp4PEFOFTKQIrPN
nGxLLuB9R6MJZJ9s1SZg+mf+EcXS+GWoLH3q7O5xn826J0la9QvtpaGQhiAKGQ8b4o1XeXG6r4h3
2PEI+wlGc0tfREJh6rpReOlfakGgYRo1KvThPrOGE2OORU6s6q8zeP3OeaTsu3cfwBUVw11Gag+C
5G4fov5dS1QZrqNLGysAYfVb6s16hY4pfzaR/FRyBzGUT9XgrIOFXugDZv8WTM3v5YGgZfOo/awn
aTPbTHMTbLsvJJ0DMbzCuXQC9KWymPpAH9089Jr0R8+Z2/4xanXP6/5u1D4hE061QnL8xjaMcai3
c51bNaSnueUZl4gZfrSet8PPvnXwRe1sZKDlNTQLJU+ypOr5EWLh1oK7GN0j7e76BE9109eZ0UPz
R9V0f8Mw1BJasZok4ZErgDbJQUcSnCxNBg54FkVOutWooq74nSuP78SktJaNYC17G4LSBfNdwBs3
rSwUF1VqywLS49fDD683cRP1GYXkmMgNEjfA3sXwT6XGQ0kpHQfBhZ9p6yzQgI7DUgYIM7FujtZ7
GXWyLR6KZYWF9GUeXs5Z7uk8A/AuR7xQ+64SqQwfSbRXgd+Kdx47IpkN1kov098yLaviSs98sAbG
sA0BZanf894HSmXHPJRNrpfHaM384YSwWC1dBc9j0TExRwlKHqpeIvlG+FS+tLyyisQPGuGWRjEL
rQCkJNZUr9dAgFIlTLLCwKYWR64/FIsZY/S/4zUi+a2/PgBehUnwRVWlmlj6i9h5n0jLozw7Uu1U
txTz9ewEBo4aLaKVYCQTQXD5NCNP+W97KW/Aj2x0hhD0Bp51uzL90f7rhHavxQViqr78CHM8zq5i
xSSpTkmUl1l7alBteO238JvAehZ/c2c1XT8deRwKAXofhElpo0B/iCdKukd6b13n3kSUDzPG8g/B
s3Olh4O6A0Ey+OlRMNgk6Vuuw7rUZMBfWZT2Stcuh4soVpAF+Aeafdk0/I6KKA6JHwDEDdOmqBne
wpSDAb4akvzwho+g8tzlOwzh9mBhefkx53rpGdzRr0RbIl8SReT5KqnQCJPEv5CwBM0bV07QIIfB
YDBOV+MBmbujxTx4zrpvbopl2+zh0rRqOP1WWY0oRmArtQ7nHIyg2hx3xxNApkSMdBdyoVv0oe1V
0B/NPldhIMBjLqXGSScvSKT7ROU4QSlLucuc408dFvu4E198Q7iQa8gzegxTKi5HOFv0rtt7Rz15
frihnV7K8JgGP+azxh7VC/GSYZPTPVnT8M/1cGxSe6k6ac0aKvsbzsDhvNkR9RfB9NSH2ylXmPOj
VxESdvVmP9k+A+WGDPpjybRGScrluxmt+LGCYLMxlDqg0HnrWEpas4QKeoaflffPUL1UR2eOorkk
fxiAbOApjHVy/nst/lyvskPafBfGo8vsCq7sGbUuTn28wgPCeqFMIVm1tHRvfwkm7A6b4NTZFEbh
Zba51rT4G1MLRmCmi7X/PP02DSylK1i9pSkoHSQ0XqHr/Y94GBkZWmjTeOE50cqv9SC9MNtIWP7A
a69hGUAJk2sEoT8D0yILZY8jg6nyxbAy/ZSrfDoquXTZOQCnfMS0ECHRef4AP7SRcKW/yaD9oOzf
t/KV9ZqDljAcPfhU8AGDKyrCIiEypNAk6LkQd50htDlvBmFnZKSudoLFlf9fgbdTF/QOISba/IbO
jJLnOkgFz97JKBQmMFtHfDkVCpaAO9SfMCihqA6bf2cjk+c3TyHqVsHI1iDqyKyq27aUySPx0JHw
BXOQWv/vsmz06Y4aeNsNLKdoEIAPbOqIU7vMRFdZ31VYOP8VbWE0i47Ut3h8bbwSl/1U9ez8RKrB
qlP/0Bs3ge4Gw9F2Rv+xKTq95G7QWczuFTQK8tyrZaRDPdJEWZ/IEZ0uG3Mw/53jnvLYHseR3QaF
MODb8QbvwU/uTttq6bhIlMJVn/Y0jCPZJ5QsIWWOvxV5OL36NS6NqaNafm9rt55mxT+nrzOnukbm
1kP6CGCbNXJ23KBXjDdC3bL1ZHJvcf3Lo/CLEai0rEwGbljB18/Qiux66Ory21iflyPfetXphckl
W6bU3J2B1AeT4OU5Ad30VN6/qqruDYBtzTR48a9R6zXtl5KZG4V6CZC0Zva7s8hhGWdhoNaz/m7N
tu/cyE5Mt3WdE0JsBw7ePdGo4zlfdCvoiiIMk84JouWpuziQbNv+kYIWWjlx5jsAtcmpDGl52G4R
H5HUrYa0cMInkEbvFIW2P6B0KJOtYI1MJt1ETJGPWSLPFDdkWg9wiJdY12MlUWg7Udty4hAvIrSK
3gltTeQF/NczQfAGvptHIcx5pbGbGWSrPZxEkHdYdpfNzC/ZA/MHQW3lnMscXBXujTw71ziPyTY6
KYFqnAYF8EeEoRC5P0rcaz9zWJ7yvWgF1tZTc4X8qd7bwCHuRy9uhQ0ltLyXWxgyvnKeEBwEI7RQ
iEU4ahpD/nA+/GH5Jtu3pukSOy+r9elNupZs8EEPS6jYOj64JynnJz234vCHOa//iKl5rLmKgc9b
KcM+1lNfRG82m9O6EuCzsBHeiMVedB0iNaYLBZCGnHUD+tvREvBzziqlQ8a0Iwf+dVL3AXrdYR8P
8invR5+2LGg0DmO2cqv+YlAcUCxiy1w4hQv3xWtjcUsP+Xm8lfQNSpVfsrD0hzmVbCo6wVPXMrhl
AJLpwVhcXXqne4XC8TodbEo8Dj0xff1IDcCyZ/+dhvW/L5qe/rHPlsG+gAu8n1tg9wTm0wMrRju2
Z6t/NeGcHIAjxLbngNwmkfiji+pTfg3c83QFzm8efaQ5/2xzTuUqLKfYDc6gDvfx3E+tTfsqzq/W
LHUpWTAH8MqHur8eN/sWFZVEkdVB6ejObSWt/iw+R4H3CFSYyM1Jolswshh8vygcucKbPPJnJsII
JW905rXmeiu++g96IJHrwjQtOjC4J25yzzFY8NVARNn1/YuEbhMtIIGpoA1se9roa3BlO8/GRQ5k
i3Ut/esbyvjHHkRLg7AjZp9oIKs3sJHKt4ddiRNBzKaAFkP8+bd0djhI+/NNbc8tEFnQMJ3/J2yy
hCLtr+pJnp73QwYvFUB13qvzvgSsXiShkhu1gfFF4cZx+Cy9WC0rpkGSfSs5rvAZ4I45iqT/rjDW
X0NXZMQ5IP8Bxdwb9kf3Ar7Ze1i73vo8eOCiGdcZc3t6Qf++TZJfyL97tWevQ4H3SCHcBWWVncy2
LkzJaIaoyqvvvTbUUyiAHWX/5hzj37+DR4a3dQlkQr3HgueU8rBN1ZHcX6H+nyFwYq4PDLSfD575
WwAJrnTbNKCG/1LxLRaviK/nXLad5f7NP27lk58ZoUPgk/BLzDeM+bmiAnN0DgewNk5SSoYUHDn5
Gn4uUKSOpej7Go8SnNg10AFwTRwowSZcbMGkvoCtuPaYhAlBw+ulE4edU5HRmdurUqqeFSwYhImT
B+1enB6kKcUyc+QXfC4Cc1+PYcOOtUfd8boHDRQM+3NMknTY1hwI4nxBTAzDiZqPYautRfqLzqtI
N4uvhKCL5ZFLtc+HdXI5R7L5WwNFMHM+aULe4qfgE7dDf0LqE0oEA+d5udvPgEO/2BBzsNiZspDQ
joE9UWQv/asW9HMMaPB3EW27sL1h4qhipmueBQNXoXzi6igLNBqLrcuU4tZ+vFERdFsRHmKGznzg
3hwXI8KNCtuf/eIriPV/zW3xquXMdlZJ2QBmKwYjpv+mMgxRAJogU84PxCqkvb4fFFWdGdTRRXY8
AVkQ0Nx5edl47ZxZ+jo5D9oVR5UTOi0qdKtFouLX/HeBzILscq85Tf3LxamxWo9zySCnvSsN9MAB
Cqf8XEBF7mL5wOIV3lKNgmyYH1LWlhkuZZjDuYK0dLWYji/bY0K3M8P/ucE0qTySh6LOv9tsBPRU
hEKOY8grI00bItouArur4ii0/ic/DC2I3DXvU1od31K1AI4sJX3pF1aHpX+RM7tZD1M+dWr9iY7M
0S9kHPbOObLuyVPPEarpIwk56uDmjJF/iWEf89yHuYtjQJ63FDw0wEM5j6sd6Mmszhi94eOIz30A
nF0p8GW2EVmYw938HLZoVjAPEJCTgr06J3QBVOxAMUkEt+odKEdoOX6Ygz74V4Q8579vWIKtXriq
IdXX3qV64hV4h2PR+ErbdDrvRT6DdmL6Xj0vNwA0ObfuNosHeTh9MOLdH2/aeK+9rJs1YiloD0fL
vXOLuNrxGDyAXlxpQ7LV85Snzc2h42nCRUBWi9aFZlgW68SfySKANCqIhMKbrU4CV//oAwN0xIDM
gxDZMIT8V0xhwuhIFUJ250veNQtoX2Otc+4SaiPddGRWlJMhOvzkOKarFwrqEkIrxJrllRiVk+Kk
bDA25m8dxOZ7RuNUsnN1+7MbXOBxfTbzLKRBmgt35MsEqsCG8lmUzx5og2jE6ImB4Pq3TrX0evQ+
wMuI37hlONfOKmFI2HLTPDqGDXH9jCSgIaZPEcjdotiCo3+OYTxf+grKN3JsIYgCIZZ/a9UsyrT6
T0xv9oMbGZXnga2/a0AvOJeAUao9G9qjaVNdqYpn03D9ARhJmf/nhpUFn3x2nJpKxkPHLgdFP0cH
oLlJk8BTAIhUQKmG7trikl06VlmwnFG8lnx65tj1pWao3cVKaAMEcbwV8rDJIjS6l0bGpseE3VQ7
TwEEsKB4FkGJOF+q1MRy5sIv+ee4QBkt7HcL8zwQr44jOyT6FyINuzA04AWMysgM5K7QvDs4Tmm7
uh1kyXTL8Aewg/95GG54N+WoPz06oVwUrPULHVxFUYyxxIjo0fJmpaSczmOFuTRcMggPhOEdopFe
3QR2qj28bH3oC44ZxHYAOCpcAl2ihv4DOWUs+/DrI0GO80hYsBfyA+vxjNVmCFx8NFZpTmoq9MTM
qbwZnk+XBVKaBKuPzUcHx/Tx/amRn89TNIJKkV9H7sJ6asp62md+J/PX+zWEKUgO0JGWfKzHXN3U
4m5t1vB/H8pQ8ZRC3RCBGAAEao8gStCgC3SX1sin6l9lrGU3XtoYGVd/3OcWF9gNSoCMuA7dSP+V
SgDg/2CNI5+coJ1Lg5BzihpMuAAUDXYTXIoMcWeVfjOBdcTOkLqGJQalZO4T/D6lgZxOLH+YiFHS
7dPtX4/3T54ZxUBHLvmiVp9eNZCh0ibhyWW8jcPQ6tVOWOp5Gv5dD4sOG1XNZWqhPwXf7kXMyPlD
5KbYdSPTE/Ab+Atfrs8kQ/lcTNiTKnkH6CezOckoCqnZSVf0TfK4+reA4SmOlJIj3oD7JHqgF4rn
5rm+MALrhFWSaQ9gIPViqaN7vHPjOVJLRDimcBLO8sKdx7bs3zviJDDwR8kIVPXlBk/gkskV7NPK
2anXobmnMQGey1hSk+IaU+MvZTXjaZSeBOgA9qiYxhioqEYAYE6p5FMJKb8gV4y0JyL21A48UjDL
qv+WEIhd0tA5ue/8EBkNFlstrOsDAs9RNfSrjQ9R88AAreBKh8zOzrn+Yh92fAy7YPHkHh5dr9e+
jMMq26YSN7JkO+YRPx0AGYfA7WVrVnTMsEMskFIoUQP4oeJ5t5tfrtvsh6CT+s4xc/m3dwz5KQe4
NRbCtoyrsIX/4hxvXGodRmPbPSIvl/OVinsEzX/8LkOc75nclSLaQ8xYQj0emBSpNmWjqB3JNj9M
4Azg9Gop9sVYqWIZgRt86Sfro5JnaFUCxrcgxN/ov2ALwf0tyTIjjoCqiGt0eSNTrl+q14GejC6T
kVqj0AvhplBVQS+HE8tp0jo5nqxMqV0AFa/vyTgmuwqIL+X/W0JjOjoD67uFplaVwcxv5Ak13SZW
nSG2h1leR0YiS6sDehAuSIvsRz2/qoEPGxjfiFyBESaW0Ch4F9DYIbkqHN795PXCnSINWwOQRZLO
KA5Rg2tJWI1rXZsDQBOG9h3fRnmDM0i7a3c5LOPMkMLpKqETTYbMrdyfPQPuOvbHd5nSp7o56CjI
+czbbnCGya4SOJeLQAp91l90hdz4X3edApwxNFctSFZM38WGZOVy6eKHYsjqNRS7h42hBZtQBzSl
ejAjbWyQUhqYZLvbRU6U5lUdlTwESdpVejYIBvASJ0lTMPMNUccsbDC5CjYRsq+4GHf6QRMpL4Ca
DclA80J2uIkJGGJFqkxi1kltTTW8Sq/eLSIoCsk/cLLKkvzjpIAjW+TL1zyJpBNJDaVf8o433mQT
HtZfTSGxwqB2RHSWvL7q7k2wFLvSe6X6qxXljIef5XrJzTs8jERzXXUdCMmSmFsIyCXxbKZgZKpf
MAws+cBYIU/ojIDOo+1ovbdIm+r9qLwznIP/ebmVuNEWqOAWFgkOkp9lxS5whqwGl8nouuZ4TTx4
jEnIkDKYEC1BwgpbJupDGulftL3ynO3KjhZNjPlcZ6BZpkUqIY2LgxTR+BPXvi4r29Jz2rerYDLw
r3uYX6K1P2uwbk01l6pPJH4P+c4ACIGdMkTgFgu4E6vAWagbssWOEu3JYr9H6S+QDpuWAuuJfbqG
OHDuFLCScU190uwpn5+NF5PVFU60bs9l33V4I/q/F5JZwuQfTXcy5Ddoew92PTA2jQZakLlUQPgb
h2qjIQ8Hc+pk19X2WU0xsgaCaWNAe7mBtL6FYVEGtRHxODg7HmOqUEH/p5mW/DQQsWPfBnawdziv
ftfK55mtxc/TIC+ukG5jhEvYP76Yfo+hZgayoTaIscUCJKMItgVWsNL4P71WGfHumSgV6b6yuIka
eed9E9EV2ljm5NS2Jtc9QFCLdBXFouTOQ+pJLRXkRrE3Y+PynCgf9HB6PDNdKHU3hfcyV/viLv0r
7Vbzna8sQKisuCFVV5R8I6XDvmCo7rgMhcaRdiDKbKPibComD9rJIgC4b9LfQmrsYzkfnecZCeSc
Z/rdjQo5Jlmu220x/LoeZl2wjmQbMUxwihCwsgSLfJQZ3ecJhZtr4JqO9OGaXuGYLnyXBZ6UjN49
qlQmkN8k3747cw3qrha6c4X1bRFxlvKWr9MEROKBEx5+JLSD+zt0cqO8uujaLvzIQPAzxKfD/alJ
LINXEEyjpCJJafm+drMKmiw25HswPBFE2e8UWj/bVCrYl055+2/yRjcHxVEUmS8jVaWpegpeNpZS
b69WAXJA7WInF9qgXDvST/92yKEhyCqeqxvperBvK/ldn2x5H5vHDEVmFIn/uvRT+uUs9cL10+Sk
skniCCcBtwK1z+DKNJ7ToNcFkjt9X6FI6aaba1GlDYIbv9qTiyoadp/pxcKBPiD6bQFhu7uDFb6k
UAB41M+2+vPIvFfNf0jpuxKP8lrKViGd5Mvfpxfd9uDtGeL6vl/Q8out+vL0plwotDr/nyzpeLZD
O5w0kjTdIi4G0dZ26W7+YVbtEhgmGGnI18O6hWNbB9clbutmL2++/1VUAVc3jOQciwrpt9Vs+XIO
RN2z7DXzx/TBq1XyipqNENBbSQiF/z3a8K/0Hv0KvEPYxpjm0Z7U8ZOeaujvkpY4cYuaX82sylj/
1l4yc/HOkwBoOG5KqHZaVGfkzZGjhAwdrFZDwMuW3HJyxhnjGQVRyxO6LIbqAayb7WA5QKolHh4+
H3TjA0JVDUqZz+wSHEjlRlOL0CrJGBp6taR91pVtzs+8RbHNrxl0VMWALkY96Up7fmTp2EMV5uzF
TXR/yjifwoGKVOn1xI7IUlExUOkhNNHuMpuTjNOtMppy3H/xEX1MS1gh5DOuQrG/aK/hdxdPjt46
fodqWpa63qzBBmP4/dtHoqNe7z7j6wFItGKIWKioh0CCRm0wC9lgmpqer+pA4eenvL0r4h5br86K
V2B6uMjotcKX3x0t48zY5zfvFFKEONNdVLxydOY2qXBfUg4SiL37Hx9OekbRScsIDj5Qzv3AV2nI
2/AvUX/kfnikogWzUfd9TxSAugN2MsdxZoOoKkp8aUBaz9ViBLzXd+kX7+Wcy0P7cHLNjyBiug6v
y+uNl5wABH6UAq7YwD7rr+elUavLgbJIAcAnmx6KFTpHg+EqJM5f6eOnW8/ry1d+j9wkgYumd/5c
TlYKesiYhbfzMX7z0wAuahLGrcqxY61AldtyAVjvJqhAfz0sQ45DHv1UVgLmlqNfeKM5UhcxGmU9
6sSttHK5IEfT0gHZB+fJmNc0CjtH/dsL1gW9GKX9je9+sk6NvCp933TrEQdCMnSy4CdkDqEzjWaR
Q7w0LHgWIH0M2u7StCTGf7IJvQ/LFrjvNtIyge7XV1vz4s9sKjwDu2Ge5bWG0Z7OeVI7fNcKFopF
2jmnZZMmVfmD5z1SCNUgZWU3gHA83eLykLN97YJ1klIb9A9ws8uitGwMw+dIkgiI2YL7vFK9Hb5n
BpX2OeILCW7dpIBjRzmHE8HZyrv3ArY+JpL4Q29UTMxITh7Hf6Tuo0C6QRjs7gx2VLdwwq/lbMRR
2IryQRdjgK5IOLGxQDXFxNsR5jJ5G+tIKGLl9DehbPkZA311B4jktHjJQ2L6okqNMgAS+s/2WZgD
0OTvN127zjK+JXC9bP4q9NOSnjHINQA+vuZGEDaF/Ymcu55zH9/rHvXZz4E3o3YAEBMbGAO52ywn
OC7dNVZuK8cDp1qBhi8QmbYTz1l6btJbPAKCM4Zqk3O987hwzh4smVdQl/fTKrxsEitXj0+uhEaA
OaI/D+IKbkyrOV8vFj9kC7qvUlukzdQIm4b9q/zKuAecq/y+NIE268zID7Cs+0wabBdj3L+xDnN8
n8iq04mMVbcKRK0k8UKnfoYW+AstocCPewHPp90k+z7MwSUQlJjzgIiYFRNKu3olbGmpzFnReIa9
MafMLAfSLe8MKgQa5UE8QTf7ZMZD5k99u8TR/PFV/iJhq1LYBYKxEIWt/fD+plio0xWe89v5RvQ+
XFRaVqm9/oVbENCMtyc9poQqkfCDT+pZrwRYBJQKmSvGE6z1CL2i/F3PhC1BjGhPtBYJvA4KMV+L
SBATfVvnG4wRoGaWJqG1zm9npl/TzBbVkXJc66UHdj1FqzqT2BVHYWd/mDkE0Xb9Fiyk47jHUhDw
PWNxTqQpAZNSsn7PvD5smOjAwJQtIuRXUL7iRTgxa6iu+nsyDVbhj+ej51i/wKif3KXBJVUTPoJ8
CDVTu8kSaa6elwY5YLp4CyCdnYkCoheJiNL8s/T2/LyJSSP+bfI8Ga+bM1lAhbBjnkk8QI+rr6pp
EIKSHeteqtluUJckNAb6cn431cM427yh/9Pl3V9C6QFnMbnV6VN6dYwdqadPNjC3Mc7v95zMgT50
FfZFBJAeJgxD72O58LIdUCPxTe3WhIoE/oPMuP5SM1HOE7D5JaxxwcySk31HiBQJRh+AVc1uG8N4
rNbedrwomjCWcwBo475cCpzC0OdYsEq+XsOjFwd3kUoCC2wTtHScifD39SzcgZr+KZu8u4T//rRD
IigQagIcf+R4mXV4uqQPiVureoXzTodh5JXJ8Ujdw5e8jefrLIPCe8HzjwDNs0C9ws8HGBwE2sfB
xkdFeRn8TzTLzqrmGdJtCkV+EGxcX8ohij541cN4P6vDcsRlB3fmgkm7hqU85mPZ/kbzXGjXjgUA
Cc0b2WJocW653omR+XO8n5FfOhTYGN9T9x5POvsEju0JbrWysY22iPd52gT0c04mIKUDJ5hQ2/bx
hvXydcA04WIDV7ua8yYf1i7QlNW8Z2d8noe4Z4ITJ/fBZkWGpKnNeOLCFPIKzmULh3UjLnq/Wrl2
nrpcpmUJ7VI9gofnoEkY++U0ilh9gpqbNrrJtWaLpcblrZp/HmnTlE1PXl4DSAxttAUWoMfALL3V
Pzl2mo2EWf37p5ha2R9gt9Ts1j8oAO85DZsHPOjnd/goud47lfSPOPw0q8kG3XqtkzmXVom/tICw
qtYbF2itIcUzUOuaaOKbQQyOJUXjUfXBBNwf3qiCMhmQ6GhJLbdJqBELtXAQm22l+xtAtNMYWeh0
ZWPWpfXUgcStkDD3J6HOxoeVJNoALiKi4bQhhtgFmTuO7FB2O/cltHaN30Vp2vpwDjLRiZt06sN5
jKYymY1B2qjw+J/F2CzST9+5Km1ytGxpux9VVcSeKitmLhx4ZLgdJwyY9EGPQZPaO+QhutBbQo5s
IFBUq9ATo5ZkqN9IO8C+HVsazuINGisss2+2TiOMtWB6llLVnbxYkD3zRtVdRkOGyYD0hhdHCEAa
DkuBadsbjuN0kcc92/IQtyOKWkI+G+5Q/p5lHvjwLtezGX5kMopdx3myOuEx4YlE4q1pTu0LnWcp
eoWa5grdduuhwNxLiih70Ce6ifM3T5+3925RFeBuDY0hwpQhuPkdxWNMT+vUgbMO5YtjVDIJRV92
OZCrPN5KXwXTgZyzY4oBCa06rHWgBjoBDKoisHU5u4zNjLzI2f2+IL9dA1cp/kvqQoQFbk95A/Xl
M34Wck0e17pxLmKssozTOgFIqRhSCrzQY4nw4XCfTZM/Uxefy/DhEu28meP6Qq6vceji4ym98yqp
DHUx/RoN5cCp8oDjOUihzmQXrq50Dx5ApKK9bBkPD4jcpRcXJCAMBDOCdigzyEMZAmeAg8SGVF6D
w0rOQp3zzgEmIwpilxqpTQ2SUsJhvCf2z7aUWoOA0hV3LuRWx4OlKYKz+bVAvKsPjjeceue/qTkk
ZYYE5su1Ts+c+auaNAV34n4MlMch2Fb7Xoqn98zFPn47ZpOMhQ4ZHe/r5PUUTJ7wlPyUv2+InX4/
AecQvAdalH3/EkssLNIcTBYY2AFTHIgo92T0QV7V52W0quXKdZM9XUosTuM6muB+dvXU3ggUZQrZ
9iB6O5gzBwisQvqmfmWdmyaF66mwLe2XrQAkOzxqgqsWv44zOQkgNk/2RbFYiH3K10KZ7sL+qDTf
kSWH+BFql+zhKZq94YrAzKES3KakbHVyLKbZamcRdCu3Ju4scIsB2SJHOYwY1RwIC8oQeURVOg7W
V/DC7lcaKxRpk3tPamCmNAfK4ITz9U6Ynd/Ye40McarTUz8fUQRRRJnKmREiwgG4LwlLMh0jnpGZ
JNmb0wS74xxOnujPChfwhk+F44VgnBV+MXdKgOGgl0XqzzLe6cbZi8BonNgl1F+NxzdOV9m80lUX
krkYBqHJUBR8LJUYfBIgmmL7rqyankuk6i48wkmr9KVJufEYRlhIofqQZ9GUZ6mMbw7EbP/IMaUt
/Z3J9RveAyYA/OQPf9uON6y/3cE2f+qVKNu5mgfxhE8fuxNzPoDO/Z+PCH8s1qEew/1OqmAt/tF+
vaZLPtPbMBx6XJgej96+aTuLGFLbmmH8exDvPvjAqWnJ7cupITKbiXcVh4/1Rm/L4IjJlv3FnzJp
sRIzXnTd6GEllaN3oHFS/UgC7F7Clt2W1d9pn2jMwZWXpowN+cqhTuUtD3XQseyOph6BddqNotgp
ZvE+QNZ+lh7BLGyFHrnaiKUKlV1UNTsAWTO8HCQpoqAen0Z6KzNjZqCBkb6JvCrAuM9kFxblchKc
xMXHJT21P5CIU3bgo3g2KWe5QToYfVWLivlUlgfvMyeE0o+5jD0cQNaqOybnOy4viaUIXiK8ZRa/
2t/lkpkSWfwOBu47FrtPigc5P0BZ0wYNZsE11RPoX2Won7QHMmE89cL6MxRx+3nkhINHDUfO30Mh
Z5LjGNHwoyxA85gw9OTT5eSY189z314YgWsd92FdLWpoXQMYdUA4m5QGIKzhDxtkSgxFbVcIBHa+
Vy8fFvnbA115RnatDLsuyuwt9LxPsbj7dDZFB9cl0sBcimx2arhQ+kK9GQED0zvO0QWmi05AYcaf
XiwMyNfHkOCUSMi1Kx1YokT7IPoaDWyJm41kqq5pIk9y8zGp+L/hmPi4G3Ix3/SaSxyxP8PapFXd
UDE5mbMhBCT8DK+DYv6pkJl1ehvZG8OfGwIuSozgwn2jgPzHJPFaKlEbPiudPBWB7eLKbqvSlis2
fb0o61I0Bbg0HNIPck04Y7QvBylrFXrNK0+rSeB+aIcikJBI6TvA+5a0GlBZ77aBlePiA6cFULHc
o8VDQkGTmN0phITGZpE7FSwJSLLZhbCEgJyVpwV+imGkqa+tNK6RouShawJKus+q6t1Zq7GhFQIE
8ikgaWZ9q8H1E1jTBvm44tHH5XRBvNjjbV002Zo+0AcVv7aDBsv3OB8iuS+QIyqGj0YULOq5bln+
BBH7x4wtnkZHYDqh7a65lX/VBB/MyhGYStGTfryA0XOBupqR9yEmktmhmDIElXG2+xKVkP3wUkrz
TseOqZ4aka+kwWXJtCpmdFaiJqv47mPlGrkJ+hBiHFgKG3AO/NKCQ2RXhOAlMKd1TLCGCBddDNS4
rDRWgCkJTrNj+xHwMhilASKRQSo1KhLI02B2asLo4JwP4CIhMaEFp2MFFtr31z1S0NIr/pzJAPZI
lBeCgab8fq9+xkw59fnAhKpVeAFiC5g5m5QTcDR4ooUH47vIpjlMmv1gMTS2I/zm7T/n6NCI0SFL
ZbaX5I5HI37H9ggr+Un1rJaykjGyxrnI/xNpUOojwwDWU6Zg96nXXMGus0H0Sb3+Q/8KsPVAV9z8
+PLtsxYpZJPFFtpford1lGBsMA8ldjxnkvPCK5PCEaBzNmYH49SHR5n7vl9EQ2xe9fX43UXJ3aPd
WwJWz/4SqHesh/iTTeJrgbt10Z6jK+P+V2ojIwSq6Et25Ur7lo4oKwJ7cb9R7PquWzjRAWryUq3n
NG999y9rKFQfWR1sKY0qpR1j22OiOGTWUPjP0QQ5Cbwjcsx5B57gzROM+pURK/dTM1I+fq7Krid6
P0MiwiN8W3FDjaDWs0LB7bwUs2IukL0vvBs9+eGmdjh8S8S88yK6BMyAGIW6dhutvSVB4mU9MH2v
tjvCEm8gmPKyhFix23ARN8wJ+DhQnZCjbRYsQA/E8FrVXwuWbLOj6gOTd9EaAbEVNX12i2PqgPLs
41Ls1QvC4+6WcrdXpp3R3312+i6h5FrZvz517xHGToZUSroUwdFoXPpL+OFNFqGqgQtbt88MauEo
TIZiPMfZkdues2dCbhUny9EB5/lGm/csWSYZHf0BRu3cYR4khq/Mv2t9VysWRbbUrzc02/W9O0X0
eJndIon4IyXEO3+fMTdhi3BnoA6StwJyQr7ahqUcyncbjCf6b5OUZuQ+7H2o7WnoWYGXkxjtRTEW
mLhTMVEcyQ0W8Lr06YpQ/CqipzBiIlu6J9nIZcJS8TB8Fv4p13uv598NUb2csJY4AD3SX20dRl6x
CTfYtoi7HcrQxIYygKAlAI4tmlM7G1QeA8Op+Z/tG1WA2pf5dfKhYOSPAjEagVg4DmxkF7GV0ilh
hO/YFibf0pu8pXF8JW7+RjzA45U4oEGGLhms2TLqh2JARt+rnNNeu+rd7PHGZW8NfQy15IPGCDvF
EOWuHlFqghOARknNby/7hj9B/JQkRwGR88R2AduZRnCVn1ttbDXR5N9019Cb1zWW6VzqkXOsft0x
DFFbzWK0XOnDYWEbItnoRyG+3NFZvneLxKp9BYg/IYdZZ5kmTa6u6qm5wpaif/lX7g7M2qmhigbP
WjR4b0p3U6u1kHiVh8gAKTQPTOu6fLm/WoX2ZdxhR0QjocPrSC5yQixgRbT3G2YFll4d/E6pbLYh
m4kyMsddRsyuH8mCR8k1umvY8qG+YaQgetCbbnUW+VE7LkIhBSaXWvkbqtbssz1z0//w7YH3MkBL
BwfWve/aIk55C3/PtwnDe+ObwYWreISx3BFyv8AOrcu6YiT+Jj1C/NjKuWCDRu1L1x+A+xmKqB2i
KwyQ+tpQ2FuffH6H/ZgBJogr2kfOS+Cus/f3KHm7Ue36p7Cr7o2x6dEayecOf+EE08Jpc3cpBq04
vmQ1WDixhoJmXbP5CdaFff9JGPpY0dNtciHlaQOb7VP0C9M/anMdrnrbd68Zx8Z5mepGP3RzPHEG
XN9mt5o98hNri0MskXdZW5jkiNbflrA2TIezvtgJPXbGCy++r1HVm1NN4HXId5mndfjjgr6qxQUe
8ys3f13K0WWuFsNk6BiJSwE+V8Rn8OwfY86Z1uL0HgSMrfnPigSDa2DARUZoj+Rpfe45b6YywiTL
l1zSmhby/4YheJMyTSVzIszzQZc5P/OhhMForR12KS58ji1gdpOSqM0QHit2kbne0iw8WR576q0e
c4RCSIov+Ql6kIRaY9bKO5TzFjQaDUkS3F9CAQfZxuKatWGf65sRvqWF/Ketc/fM7ETTmc3WlB5n
br/JV5EKlbeP0sf3xlrIZtdx8Pb5LKo6ulewHxQuFQ9Tjq1aH/Pnxo5Ad6hrZ0vzP3Ns5Sy68ktt
KJPww/yPh8KUkW18B+/K244XSmvXgvTukBpQerYmmPjz/05cbtf4eArWLxZTZb//VZqxVs9ckfFo
QrGt8mutPjLL0G/z1u/lT70vI/xIHHEM3fazLGzjYRm5AFUGLvzu3ZctUFnThqPbSgWx0nvOz6ub
Ka7ppUkRNCLzEppQGQOzZf5C6pWnP9kdPVXm4KX4/oTv7YBSffgbYaaFFYCDMawnWTyaj9jdS946
eD3YiqOoBZsB13oBLzAJ83PJeG/K/rrp/YIHrnq4kkoo5CQcpWtr8R1H4ulvywcOAWPG8/TNGo+J
bRqNxeabhOifECKX1GQcCMdoult40R6/xBi1h3Gw3sZcRu2lcA0/6vqNXhkzcsmczUoeCsnPKCnI
yjXi4MZycEekw64GyfeX9oBe+gcmu04K2rlpLW6FlpCMvMdTG43ISIEMiKi3By5bJCcUakI9vmdJ
saPkpj5cEipiSFpbK5lZ4MXDk0Dp+gkVfo1Az7DcvGcrIVArbjDZOdd3+93qu4bFiFUe/cYzplxo
m/E59zn47lnksqBHbuQawDno/CeF5r6baYjc6VEc59Ukye71ATjpcZcd5SGO6dCMekMcyP/C4Y+W
PcCJnbReOP658hKkoG+ETfVAoDJfrmLmllwDwQV71kYBY2PSt1W2k4/TF/7pnH4QQhuha2+9YS0/
Ha+4I2bzqjhOarb1CTJf1xLBzTpKwSVU+EcnrZw42k3YszzkkIZikNDK3DVYR+mBgtYhA5zEu1zf
bkx/Sg920sQRc8jEHVLdrztS34GP926q2xOiDdMaulk1Ij07VKVHS3cjcO5+vyWvahZA0GwYf+jC
h5tFDyal9b0jRd2cibi1vBFfG0/ZRex5hdy/GNn/l0mpVJHIWIQxadrjwFA5Qosverp6HTPYKNSh
7nxFE4spZYEAfRTHyoQLE7lWUIfMmjW9sYH2zWN7xJUDtD+r6/1LbPjo9cf1df2nKC+fVGluZ/ul
xhLnpmTG7Xdloz/D/rsyRM4S6kLp2h6drwC1ZpYdnd3Q4G0G18gDyBeK5kZCfxFWXJTLwV1e8bSV
qgj+dhhBuJXjIxAhXAOtMuFcCKk03SdXPXKFzITfSSWRmJXX6peWuagGhG/kIdXa4WWhV0vGEV0w
r3tEe3jz8UluGrdU2oSPNyyjamKQOkHUzq3aSoUpTJQAMlJJdkPMXNde2CjEMpiJ/F42riUGLbBj
j8WnyW8RhJK/Y2GogAYvvzX6TEk4VPQvGayrEoLzC/2USWLscX7S2J1hhAJBxb8MR3hAI7qSX9XJ
EyuQXkGH94FrTvtEzrERVLLK1jmDr8vJ0Cq0lSTfHdP8rdyq7UVODYj4UIO/SlQLaLW8vGWE3wqL
cH9S68Qipu5AQkbLfr6FLd/rBwd3DGcvz0XuWBtvk5nB+CMp+IvwOBv6jO7u2o7QV8EEncHMPinq
cb8pBPFvH9Fhj9IssLj32mqB/5rAb4AQqe9LrYbnR9ZSv0eVvxrmtUCW8AbutNXtQA4Fowjm0V/S
OkIoNSRwHlIDEURlqt7zyChgFQUFAnEgXGX9zf0vFe6y+xYY1C/CYjJDRXLHpMbN0lLlrgrtxg6C
b4mTBz0Zsx+I569sDKCkeBmGSm0Wpj8yLet0Apbj1FzP70ZH7NBt0tah72Jd1cfzLLVECFtlhJK2
lYnPiZWrHyZVDel8LP9kJ9gZju6efjHoJFnzTi1d00o8QnfgiV6cuqhL6Kzu+lnwtilQ4lWKrTAM
CamT/E8W6+ZzNpVFrQ1FCefW3HS5Q6ZZo1sVFTJV8mRhLGWTvtKMsJhHU0H2zb7gytaZueMlwhf5
3H3wDf1lZXIw4stm7vH7NkJFhDOpTVMK8roze/zcqfUlnwg9jao2gdLn0n6C+nwDjBQJqDo7KC9W
uD1VbIQjtw1Ykmfp9DmW+7dEWgx7mvGV4fDFvcPzVMzG1y6ZfB3uqXrLwi0DkHI/YDcvHBB7Pj8A
4RLw8JUUNINIvp3FxA4sy1kPAfx4aRMA0sI71/9QZnFGBy3BY1wFUrZCVqxJbktwq8gacKjL0lmk
oGIymygwvTr0mM/Cr8TNlEkYpJy/yKLx3pk7syXXepUh55KwYol75ED68oGbVXZPwot+Kc7wSMoz
hV602a0TisWrYi4rWwp4jxesQ8Mxr2kzRhK805JKDx+nCsq3FhNC4c1RSVPjihX1YcPgjgsiBw6C
xHQG0A7UqXhXqHKIDAofI4+9hotW3fokx/sDi5kfj/X3YGL1oyITkqyoSWJSO7/2fGxjLABGb3pC
EpnfqJoTznAZoZrg4iLlBpVbFVtktNimcPGWpqssWP9UGuhqghJIc1d1NQXPlk4YzuYqgUBMdM4M
75mpncO1htPjmJdTOtlrPybyM0jBbT/aRLbMfBBRjXj057MfZBpVipN6wzMJroMf7HB9LsjiX2T0
srY2ISqt4rLhXRM3tCbBKfv4/HEerrmEAq4WWdWL4Q67ft5gJnRLrsRgGUhUmG7gAwLq8dzqNdLm
Z+cwGXBxfH5XOZONc3vzG1+wc0FfzqUYdIRqwMREQP7MboQLRAMn7xdhbQ5aCn90Z18+MaPMQtoB
kyejeHvfvEpQeCR5HawAUrkYhkUJVly289OsUnBJfzZfX63mIS8qT+FC3izIAZsWG971KV4QBXYJ
WtuK+Ith5zsONXi8lqOHUaHTJ/tuxzIYt4MtkDOYbFJyPEfTHEsD2dUNpUnkFIxx4JFEyVxLsA6V
d+vrMEXaXsP8aZ1FR9kXuw93LeYjENJmP1CpY3j26juJ6z3ZbDbE0/PQ1KFNDpPkc7wtqE2n8w/s
H1x8frSJtOg6aG0IOPcARnWaqUkneQhdYteCxiQRr7Qr0OjtHe7FeESNewmc3VctAHmIb8lEpdi3
P+iW0XFixlEwUd9q7rPWzyOh1mx8nRyR3KZCrZfPYJu+XY/vJmoOMNog/fDYAbS9203hXFLgCseg
Rx5F4VmUZ9nlQGDVdB53uYVA2lXPWruofrftfSZ6AceWkMpyV+Sb45q9U9iHImWs6igaTp32fj3h
JFfeYAxrUERUOBsmigsLJuh3BcNKsk+qLKOr2dE9aSFK4BomMkXJiJBThk50iG7yjNKcljZns61J
iOP4DX2xSbLfkBxE709mh+wqZreOsYI7hRGAnc7MlBk/VRoLtYRcnW0bYdTAaAAfzuo1RnrkPlVq
5hPVZCS+5zlwh0dRAhLoWpPz/H6rDMfjTJAVQKVji9j/kVdraA2+rHPfqkvVkcE1zGXVsty2LGVE
gAB0MgX9deAdivpi5oSLrRFD4iO/8SEEd0b7TPRSsCK0V2D3XCqMq9UZsWazMxJ6gtALECh4EcO0
toE9R9ixad0f3XTgKyKsldgD6214oVhLGhKO7g+PGMoAiJt46DUkQ9vVMqUK0OuJX2jZdj4ullCi
RuWVGbx4jzqWpMzL69W0bWk6CVE160hOVXYI0nJvs6GnoUj+h0Z9KBjjpFAF/g4Wa52S/DK+5Dsk
osj1FhmOKOL9OTBeiYQ9efanVbpiHq3nHHGlu+FrUKD8ATM/YiSwVQ/0cdzIqOJjmSDYWjvj35/j
AWFSVwROnzIE6iJ6dPbtBDa81EMHjMaMrIlCjH2wASEpwu+Y5HTF8jS4xllP6xlD1FGTTrCF3YfR
IxSabzPpuq19vUX7PElqL7ziATi+nGOD1EUO1/9Y2yFh7/hc0r4Zf23/Eh4Ujs535T/YtSNR1G+r
RSgCB+SKQY+lQTbDlJhrW4833imSO9zhWPIBvdjZKZzy7o/4pVJONnx8Noy7gEmFX/YZYOod4ywy
t0Y79IAf68o+xgagYLqPl2rnPp0YZLXl87a9k5t7cgN3v4AGXdS9dRL8bjv4zch0hcCSyfHYdojI
RvwbLjpCSoJeBLI5SZK6ZPDbfqJFxfltAdJ+srujMjOD+3joaUdxxPhCwZ24umot1gByc23z+Ag5
saEhrWfVaa1EzHkjSvYWWMRJrHQGLXVij5dZOl223EfpyJTME/KMAigIeNoR/CtsZmec8DC0kpXD
KMiuLGErAsluzarF4oynZJMHVKJYw80e4aBisnhqZTzkrdvm5jgQmhxNGM5tuvRZWvfqgzPAsGug
UU83Q5swW6xNtQQK4wh/HtLXNfEzZFKFT4Ox5+rTaf9UD+Boey3h//4ZoV07v1ryY/VlMLYXiBK3
A6j8sxC7tOvd7V3WdsdR+k6Kr+TvhyRQ0iVO+AnXXKAg5IIrORxXJ0R7J4JIBCi4GZxMqQmjVd+J
3LXHBQ1TWqXWzxm2tcBb97V/AtGidpE9Tr1NN7QQKvZJHKHsruEKZuh5rdxaR5SlrsK2vP79WtYO
Vzh1T1BjyxQj0UE32Ee8wolrbsAfZpAv8qzNeh4G9l8eKmoMsOfr+j9R+yA8C9gCwsvE/RaJVnW0
y5We8Osx05572WVQqRg3xfrb2Z7MIOcbeTgb4y180imzej8/wIxC8Nfs9JRa8bNwNA0gyddO/huX
gYD2QWpTZZk/tDzMvUKFpTsDB9mM1EPAiZLdUl6kI2K1WawUJXWC5FreUcJJrO63ywUwCf8+Ld3t
fwNhUaWdJQKsELBw2a2xvOYNrAHi28vOVRTvf/5Oau2NP9C9HcJkIEugQHz2F9cH9XaG2e6L4fTa
FjCYQNjpuvp/LE+UuCjQPyLVhbTjwmT47UzAWI8mLNlvRF7300rdmC7hzelkxs2z6Ftt8m+B8XAB
3epC9nUhjR+yd3AXrTObTrdu5ZU0tV0L537cqBiJ6Vp55vNQRNqqYwzm+T9HzCyo+EZm1bYN8e3g
G83cSVc2Wx550K+6ei2Xpdmm6p22nMuWOZdWbp4QMfzAa7M3b7n+tHCJia1A+RSGRzMNfZVV1dbH
+/3xJ4JhVAmedyH+lKakrjfx4ex5t93MWFXDcd/tpTWx739uXeDumJNlT7yTlGUj1tvCOVu2pakP
/HsdljKC//PBWv712OH2In9E7WK50SfShy6+iB7h84JAEBka+S0ULNEzImmX4qsiI8ITW/ecxszy
YW0bxeVZSLI9G44kECRBbtkGcjqhhIF4Pl6BSrFI6mrrCHMwAotLsQTfaSu7AvBaSgw573PfqKJP
sRt8FRqjK0rTJ3H+zSn4eLn6feNbWWbJDLFvt8xERQdfHMmwYgqvXFQexYVqt//6tUcPNCJG9MyB
PHx9VsALE3haIwbPyeNqfaZhnXpUe1/YIbuiC4DylqcT2kx8QhB1YKPtjLrqZsXTMT7N5YRBTuEd
QCk0EYwVDKvK+yG+dITgUHGz2g5Er9/FEa1ia50Wy5B2Ketavxf4Uj+hkfgst6WGFouEhiJ/+0Ud
lvBwT8PWS4nQppOiCWugLtVCQYV5aERmsOYSLzPWIMHWTr0gnP8MZL2wA6GFdoAaRWBwt3KhBTpw
U/LqgXkXqAtpvg7hv48WBDoPh5fIzLkgWsk/qGZ2BLahrVKWWRax2ytB6YObiAa3JFnWLhY3Ip2i
MzKsbVz5DCe8g1hUxrjovzp8++vtmRKvAoeqXyrnG8eM0Y9Wr5v3QK1a/EBeBjGl/YPSBezGjqhL
A9tgEYgY4MhrRigDPov5o0zlCdjlM8sgZ1nsSrKxvBlr0IcCurSIuATvSl9wZWi88mSRhTvqlrBN
lVE50qtTLyRmTuiDQWlyOnefHaZLqvKWr4rV/Ylrd6cEkgrTnwcW1O8HoFc0aLO2GuYZT0NkNxjK
WBDqVZK2dPzoxew9YF+jKX4RFvEYld+CQQqGPwl0oUOuD5BLT8vzpytXtbF57Ge8+S+TxqYxEzyW
5NqmGMndX48IUa7uXkbE6lFAOacW2y3vKXc8KMJxVHOwDQ9PKfi4O98PN4sFFawkE2nFo8VjdwJw
ZMawKN+qjOJv8xHj0EhbfvKM/pC8Ao3KP80eKehz53LRCYkmvHRKuhz3P831WptMx7IZxXxgUdkD
mNitdrQFRu8gmYw+EgoPQJkMT9BaXpWxWM31Gk/HW4VL8PcLxzxaGd2gvepFqxoAquT4U9k3G0yh
e5WR4zaSfxRyZ3I/yMu/6mdd6Gd1v7VS6t4Hvd/Og03Fadz5zWzSUjpYQpvtQDzf39+lzJDz5bL5
d0TUCEmAc2XO4rZ5nyuTt7cNkQDHDfaL56c9u+w7v/O7NFcabOBANUcFb3bPwixIyZ6Hh0cS1vDe
S71hNn++8OrG7vjlMU4bEi+vrvawWeugeLBD3GC6f5kXoYg/MvVfOypF9fVkoFtWJmOCViuYwGdC
7jaMlqoetGTV20SRBTEdkWgTf3lu/Y6doabEvilQCNwV+fkK+emvKCVWDO85XSH/meqBfOw4HBXE
CCd8QVkbwUto4LuOm4iGpT2tnDP3TUXYjgl+gSuXiolDeUjKH6bwES97dM1lXcwA+nhBiITR1U0X
aifEh53fLQd0WPev4bHtVPtKai544cKGg493/SvijBLLfBZtKKsnHvEsmd0osb9KPto3LOGrGHOx
0ThEm1at1fgm13FVa6TYHF5c4fOPIzPBtkdWA4zaPSKpVTOCKNuulmUFTcUv0uPfICNi+LkkwJgQ
jphmJ57LxTpr6g4cK7Z4wCzvPxpO/w6gymUtCE85BHtrYgA/go+1RxPCp4sVymToDiO2wiCp2ho5
oThrie+BV0ERdjllG4D66Ywq+LDPSCYFItNeNXuq52gcKi7kXvT3PgrCEb670MdV/eD/MreOY1rt
sNsdBZ979R11qdOaHEFoYZx4rFvJKttVi/BfHijFPpHahhQjjlaDDK2n6WrStb3i1+riXe7PnSIx
Hfpak1+NhZUNNQgpd9lKmCz3Dw98B116VYaRyb8RTV3sORe+aVTm5g3iWX/Bl71SFVH+UmOlWIs6
fHPlGOSUneqanTqIxBhDDDoQoOj25Y4C9kSp/lSHxJw28uKHhBtWmvvruruJTKFFk49IDyuwofKs
G11WNQkO/Wi6VK++tCY0Tj48Ue5Wf9Y5tmWMLfe3qydpGSu0q+FXbw5v1RtN9Q5c4T/NZvJlFKQb
+dUF4KuJghSLAEPOTVut8CxCZgI6sDffwqwh+4qPaw340UWeHMKUH+b9aOO+nXIHHnRVlr5Jpagp
jdWKDyiCaaPCS1Lva4XDQZhhNjplVyDWqbqF+a0ufKssLKcX7HhMJigt+8F04iwhvNBlsyPSFfbF
EbhsrjgJ5sTODQQxdRJsLtyXQ08nGy3D5QDcBmX2Xz7NfzH1j2+RYzc8y5HRm7+GHzFVcofk3Xyx
RovJUImvKyejsHvbrQA3qkGUVfpPXJhxBr4AEBcDaXNbLbjR/n0jm6KIj8H/ioH9xBrNheY3aHMz
SJfIj7RQrV4S5aA3JPS42E9HcojCBljR4HmuTc9UfPeVTDeBaafkwUiKtvj8lk/1VVa6WIxXxpE7
iGpprj99UObCuBkL/Kc76a/3Rxx5TcAqQS5naaQCRN3jj3daTjH63pDZChhMg2dGdK5RakGNDBDP
C3wkn8N0jeHQByNPnFWsVIOzJbpNMnKi7pFumP32U5et07zvbo7wkWKJD7iTxqWYRukI0eYinkat
EgjeU0Va6mgHH1nYX+zLzLN+iblWRSGky3mkGbypHf2lK4kLhVU4XPRQS7cPrp7C3WcEu3T6mOEr
iXH7YAybf8CC3SK3MeF+lTja9njOr77UbDAwN8Hr3CFG2UylkvaWLc02HDML3/F61BxQKWuTK5LS
LT0qcqYom5IaYxpEi6m3nD4QWrCK9CyauT3Ir6fgghNYl/LdzsDOeGrAKFXYHZp+iLNwPc1DCfMP
zPgLc9B8zwsMFXnxalkuh/DfhcoO7BJjBXfLD9tOIx0a8kqnPFEm57LgA6bglx1xDnt9DjtmhsxI
JgTZuDDTQHJxI+TJYs81XEva3FVVUXeEZuGLUnBdJ0/vFVFs5SbHHwQ8Dyh37xc9t33TkEbaF2dJ
1KpxO9/KjcEQ8ZSr5sn2dqAGp1NB9Qtk145Nv/P8YPyxRuzRBrgtA602qs2NKKBYap9uGcXjHKND
mRhtHrbRd98NZkEbvJYi/4IIwRHDn9HrySh8D9uu1tfn/KyE273P0Wj+zL8JeGH9paBFlFb56t5S
lHWh77O4TrRYIFrzv0AgLgTj1SgQNkNVaSvGuNHsyqhCIDHVE+6rNDhIehwknMLzaOCg8d5fJcGK
p5u85erN9XvEyCcH3Dx5d0NOPV15FrOaBAYsMqlGrST4XhoYE/G8QgxNWZAmGZ90E6PxTzp+yr7q
+QS057cI7U3IbAg/J6wJLDdobujx9uhxN6QgQAnigI7B9ZfpTQWurGg1LQAKoWYb1khw76sSNpiE
YnPnYf85hTGoxkqnnOEIp+On/Oj/Qcw70PfKD9+tG3zpyWf9SUNyLKWmQCz1iiqSGtY5oxQtP8ZR
ubrzhe7B0EnW0wpRJzHCWxzYv3dSNe+SdBo/rWt4eKqDskPIfWlWrzZkX3tmAy7QCxhiJ8ONzy+j
hzQlAbAX5ZmunlcYkXp1n6+xmMzlDwwIKEIjgAOLW5RYHDgpawJGnaDHek7GhiMwKBDoadp8Ci47
Nm8JaXTPHSPHOf+CgXGWTM0ZzPyveT5r84bw2gIau8Zq2S4O5kkEdqu8W8N4amvG3zXP/x8J6kAL
QUT2h4eL+JLxBmPzCYgqlccfbGrzCawmJReRog6XirV5CQPtYyqRMiqZyEN4mg4/IfcxhEtQPQzL
g1JdutAs6DqgBTb4N75qKvHXtBL31XO5uUjWRy3JXBuIXVG10ARx88U786IfMRtXyJtQRjRfTAmI
7xlUEDxQT+MOCYfzBJ7WDyX4m4g3R+DeMFQJ0cGz6dxag892lRMLRK+ognoZe+FbRhNCbnAcA4RV
Ony/bbkVs0prdGm0vCn/p3wQ10As0/7Rx46RPs2hdqa36KWMP26AiPSDGir7MtbBelwxoirAytiU
8FJH3RK8bkhr+Y7oPVmaAfJPlLrnuUxZ94DhNIOzddsZmBFAqPy4lhJJZoJQ5BXAkUveFxmFrlGB
F3od/siw4Xs22LFTg88wfjhFTlPh+Qv1UZCXB5oO943UQhyOGyKTTD9U9ZWn0ER4yJ4rigY+PXSf
U9PJ+BT/0qrIoyj9FxUZaCeIgHzYWhhLuKHyhS96Xgy40h6BZA9Ffj+d3U/5vNEkaIsNYmiVCDpo
DMB03zLQDqrFrK2sFlO1fy8rdJVBdLciezVQqmseMHEthuCVAdZESslRvKYgcCXo9dO9JGbh0WmK
xf6SGe8/BU2TkKSXYsBKEEQmsl2clP9BtJGGfDLEw+vJJJMxiX44GSM8E++YGaqxT/GBjFrSer8I
vo8Ywkbk+biVjs/X5RyIdQ58gbI/drLvcVbDDeClFl4rls9tDMx2jDaFHaXcu3hAiT1OS1db0+aP
J3jctn/sV/xufW3LSy3zLFgtehxzqa9Vf30DiQe7VfyIsIHdxU4sELzQOVhDu6muIrfhiD4GVY9+
LRH00A2cqWA5+jmvsVoqNTsUIp2C34Ar1JyEs7ZlXoTVjFD5KL0zGpu6M4XON/M4IBhG3lNyIc2M
57YpTScVMDXieEuGBBTitmHdAERGyVf44wruAgCs2/nFPRRNxgMhqmDPyRRkV9CwEgP+yTdXqupd
6bapRGywXI5En0RAuZ0oTTYrJ0uQu6VDVMDq36DJ8UVcPlGY1Oal7MhNxZoFIHShpXb1afCm28xT
mWZsmOPu7Tfnj9uaQRzHimZeINez1V2R1y7vWljWgw8ZQaejKeld1PDGspVs8Obn107Ca0JW5O2S
NKO/MPTsneBsKV8uDLDtJ7l/DofTvhQTAnVBEjht1r9ZP0543PKsfXZX5nVBxZc85T++y4ME/au7
n8tWNTimuad1ein2qPbUUGyIyZwAx6NGSp0BOsILaY299sU4LinWCepMxpVOOqa5+0Z2C+LC0rki
Bnfzv9Bomo0x4gM/ak0MbNQ9/Wvnvq6bCPVs6unU8qZw3udZjcaKmscoHtjfCaqw7pcc89EisgLr
GNRnYdq9CMK4844L11Xm0gaCwhjv6E1ZuwiR+HhZOj4vkR29R2O2P+oWLgC5RLWrQDtDH3ucc+r+
wolsgn6RSQV+BB7hMKxwFzIa+CudzvSyoNvmOTAVBgXqZqOXCZrglbz4ZmuDAampCGapizBkd2eQ
g6ej5phsDFfXnYPRzRUpJn5AXlyWfDkEOlf5fMOB3f+zxZLNqE/ZxzTSzy7lPmezqPi9FcTfUOOr
l4gEazkT+QnzIoBCnSv9d+zH9Q6xaEUdj4Yux+XAlHO0FIOmjagMZgUdsBwrk/9CMJanItUz8WwT
xRbZlheUlDDtNYC5OBt8ZUlIA+SxYTBU0GGYlGPLarEbvOu7v88D+LTrqJ9L62Bhya+nCqd40NPC
9jRBbytzHcaSB8uz1N3LvSuBd4uhJpJF4wfRub/YLPd4FXZHB6KCeGFEV2J0d1Z+u9NGGvEKlwAz
PC9bAgx0lZJjLmuneu9g3pcosjS1+PDUJu+oP/YXJ1aQwyOo9YR1sPCm7r5tBZaMBDTQxb97vxW4
UghGAdj26vyaNBN/W4KjfLsgwkAfmbNlqEKIPqbHB9Pft5Pd6ldM96ikK7Xm87TmlMmXAdzDAHwF
youdtIjb7BlMCl1R4ee13PswHkp4VnLKZSpyMSaLW1Rt0JgJNU3he8AdmoDFhBZKvpvCeW7W03eY
Vu0ZXPQf/cHObCpyTSLd7CtY8x5dcI+p4y8q3cAnwxSkNVRYYzd91503bruKasbcJ7VhhfcjgjFv
K0OVOyDusizvQHYOaZKUDqVDCjWRd7VeKDDg2h6v6NHhOSXwtbOYZgIoSXcH9q5mZmi7rJy6ILY+
75f0/lhXWg8SEBrez5tVmGS/mzI3pRz3qPb9HIakYHBNMXBNChB0bS7ciiah9r+Mpe0XXFbwBpSc
rZEgN5P835yvrF0/9eHTZYMmebtjvBd0/ZRS1OdcJnSJyGK3MJdjeUnp8YeRzNAqUEpiTP3WcjOL
DQn30JGmnpDZAHUH5/Emvv+VIR2RNQrhupRU0jv0mcDVNbqmvLbS2Zj5DW/PKA3GSv8VgTU7kPfF
NydIFOi0NX01TSPLpQ4kbGF8fTvk8dl9GOKStjtCXsavcHnKsvTKEodCRuVhkIe/i0nPJ7UhznXz
MjWNRt124RgC46MxWAv/eg5tIYH9b/P7+bb0xkSmzQ8hkLo53n69Vrv/ZUDmOM97MG1sRjRAGdG7
KglJDRMcRG5ywcCvnhAAGFfdHaE0LoyiaeV+sS3uF3qp25u4KasvctqzKDcQFF9FyGxW2dKFhBBb
lCw9hBZ01lh4loQ9acaFfdx6CnDWJ++Rz5ABphTAcEWfkOpk9GhMuWLI0YLC2fejzZg5meNs3WfT
K2vdDuQpEHiRfRiYPIVj6FDbYESgTv1toW55lUM2ukF1b/fQuQvvlaxFhBBskMGyzMVt3CON++Zp
fpBCHal54QxlLbk5RQKeNVU1bLslrCD1s4xQd70OJl7gdlURG4JaRPYmk04bXE+4yFXHyeDfYdvx
5GLtbLjpl1CtBhz+0nOUKAn5fI0gkn/fNns8JkIeb4M6jqemjQVG5Lc4QfFl05POACZPiYGFf6JB
xbWjkzrwQV08S6yNtTH1jfCLtuyZ7MClU6SqKK1Xvj6E+LRtw2hQlpVqFQRHz4V7khGtHUZ8FfF8
qcfOMZ9Ceg9THCDS9LDOU6nMO/+QNqYIZ1p7N43Pbhl3T27PG0TOg7V8ZKWsZhF6ngDA3iyRb3F4
LZvMA5Jp2BPYVPR3euIJvOZZNk0/yd3yb/y1xMHpSmJ80DKrgz2zYiGUWXt8YzyUkDBpVKWqHZYq
J4bqAhKWe2Y9QyqssvS0efOjs1wtLGo9M/4m10ZW/iELQ9nkUnh58DvcHOHwWiKCu0k/alf7AU6r
brbhNqbAUtA7u6LAuOuQIpMh/W7Zd4fw3UtNxXyuv0C3ji9MoF247zbDHoTA3OKwVV5t6qK303+q
I/k4ExrAl65CN/ukpb1XH9KhN+3ipEKpeIrXXbhUYbF8W4e6eGqi1HoWSZVhVMtQnfDcj0JbMGOW
1LYIvHmU36HBB9ZHbbwm9XaKr7NBjQwg6P1O+9TUO6I0REFTeh/wr4UVROaILCZyh7aSXQ62Psul
7rZI2PvyvR0TDuWIBPQ30fkj33p2Lm0XfasJMmT7BoYAQMlT9Vo87AS23Du6/3JI5YncpAYaFfRV
wEBtGzABmjnSQPFC1+O3XsCqt/pIzK55t/BF9t0qoGRLIW3t+YT2i2fApqQuphgyOPXafvn4RAFO
c5R81WkRQXkL0QLETIXjPzUp6XM44vayO0UwToZae3hvyVgEf0aEfQ87JUPm1RYWejHHQLFdI9+K
UXJuY/1pVX2s7pCEHzZC4Fk1YIk/A4R9BDtr4WSvRHLsi9kJlvZiWvghbxaZfr/Malh86vgFFkCL
WMVRmeV9KaPcbwgG5U32yjAWfAbtDVfqUfoxFzmUL4RkQRuv6gXmPzqqCnRpIrm7+BS/QzmGutSm
mBjeWwoJ+sNlXyVet9UXLXFa8o7zN9ZB/shcrXhfpCBpgzEr7+r1IeOzOermEqOjH4kIEa5ez3VA
Br/QDIujlJT1mRAJxE3+coE6vXAi0lqrJeG5yPXFszF4zz10kx3GytTj8REkHEYOhqrixR9Jd6bM
eerae526FEWlSsr6DsXwUJQ6lxif/fBd0N+rsp8BbE3L0yQ8q51XYl/hOqMmiGqBvCzzDofxZXC8
cps8nx6T6nbWMZNKHYymTHyYY0/o9sVDXhGEgBd/iMo1y1tCyHdpBnV1Izl4ZeHiZ7B/p0ZFYW7L
xZCVIpCj4EKtfuMAySepNU2QixST5EgzQRy4W6wpL5232dJmw1IXZMof0RzD70DV1FEF759WISAh
ZZ5Ozjgt2pNqM2QoxJxP30JCcVVCaokFRRIC0Mw6q/lHk9k9BtYUXt8d0dJ4VXP95leaczA/7iEV
SfW45UIJrlABpU6V7T6uNqwJ7bWbwyT60WI1awjXXvvZ4dLTOCjpz6kb4b0fd3ykh7Pdr7A1RlTa
7GS/yQs0bbTOQhfJybRPdc0obNPA1marnwylhfnwxaoJ+ik10lqJBB1R4BqlfLLdwts1P8AX2jSC
BWujdqSrMk81OcVPziSAxyDJvPpBo7C4DhiO6Kg/rFZB5LU9LzwC4Mmlvmd0jYL07Y2hACr+t2EL
RVRP4hKlykhNhtFyi6h2tDWrSwZBIcsFisnkPLdV1dxs4GHpS/pIxuFjlxRw4RELJuY5Ynl5LFBy
+tl7YYdhu1NZCJUU1yINfMFWz6LRyLYcMGnBkvb1rzW8n+NygzeaLQf3wraVcSeV1N7ltwL1r2Rs
7oG1dXXKAZoUM8348rsqJw2WsHnZukmqdBE1T2BEIjPYJJBnAZp+b56cOkdwNDNYWRPgTI9vQbX3
RQIVA7LmBzLcMkW00aQPJIPuH8gMm3L8WxffgoOeMsSShG/n5nBOpm44kG1EsseX1hs0gopNzxK+
IQotI90xdh4sDCMoZABF4wcKnnze8rFIya0quyK39yiO+EG6DujkX746CZl7wUtbH5AhbNkZ7RXi
27EzXSqUb7wQ2luxSrJmIGwRcAGgCWZJdtCA0V81aWGZU3Tv4DbiQKfrzZIJR6GKEkXdT8wNy4tb
xwyaTyeTkixsMtTUCNBL807ItEiLYfQDeOBOFVWzGfnlowwdUseY6ZKeyw5OugE+HO5o86kM1A8U
nIcpJZSWUAiDeor0PjRTu1W9fZawyzETy22kTqr5FDW/HG/bbd9bcDk2iDqnKp1UCeBqLtYVlfg8
71SOhR4cqhATsosQe2Dxtwwrc0TsYg8HtiIVrWJYQmhGM5m/EfTY9Z1+pI2zSdixAlr5t1/UO9f/
O9Oyb7XwfIJv4ByL7PHiPSLaOWUAf9znRahsEqamBp977EazdD7g3PU7IpIazjfedVCWATbX9doz
ahfModY4Dgcer6K/i4N9M+1Vz9jOGH/2vk+P/KyneHlNzCE0/whWw26KBALV/HwA848YvRnqXK7u
i+y0x2xQ2e7Z2QQv7sKpGbSLF2GBhzAv6HnVJulWZqR1o3feujM4CEP1z8TLYvJXvYrzUR550axY
uLxblZ9XaNEPptJKruwt9asvI3xSpPeSC+22KfCqpDa7bT1kZw2Pld7lHppR72qMibKqEgW0blba
OhNOdmW5CajsENDroJyKbVeIyGg72DtPealOQ3ZUUuzJpX9MGeqq1GmuluFhsmrBLr7bXu9GgbPp
4rbeTWVCpV/ezDPHGL2bQi8qFv4pKJEwCv8XzuYMxqTfUe9qBht1WT+ddojJQ+YibTunrD8W3aGG
X5NDo7wetwhKQVbG9WJAk18hDX43y6bXkjx6IN7etYtULoZ9/MY1bclBG/VUwY0bKALTi15y23tX
yO51BrPO0Cg4NLaFO4cx/tSIiFHu4B4arDcZmCEdBnUKOd+DEfcOqqJwFJHW79UfiwCZcnYwyBLC
o+DLdpPJrDRbcEulUgfv/T1u4tm9OxizapAAqD5lOpJDYPvP852DIMU1N8Ze/s2Zq44r2FyO7gVd
a/nUelof4aZjist6nfivT/iCdeCIOVZulAZa4p0Y1YJEJe3DJY+AZ+CUmWQDdkfsAolKUyoj2AGA
xZVQ/A3tvcY7d7I5eJvK4fLd573/4ITtKt9dSdkAwofj2f2bGnDUWx0ck1DMXuKCH3ixz8pktdtV
kdJYhTJHNiK1cbyKrkpRH6+gAzhqLDK2H8ik8OuyWtB7ls8oZlVa29ZcCGbpt7zGcDjQOJRdHZLr
UT39rVEJNX+XfamHEGieymVpjPZEhT+8y5cwl7v2j1xAoWdGC+JfpPRYPx6yI9mmxOtP5B2/TgqN
KX/5sIqUeTaVQ4liJxmPFBDak77AVffULBm92V/BqyJUh70jEl/pUadFVZTTOXWgAQNEuGz7Vr9E
NbZp2hZPTRjAlR76cmc8RuXV8d4XfSy3T0X8nZ07u2wZjnjABxnYlfkq3R5N7p55+i0N8NAnS5fK
cy5YfDkl8K4z999fCaO5aMP69tC/fX6CVDoNlLvC5Uzz6kgHVgDDeYsUsEcHpgNMy7PPy/8y9DkX
Em0xKLh3FMDPjLaMo1eavU4TaE4siYxGRLbKrQMFWwEJgCVjHfZWIEP3ZYl7UEha82oKALYU/PEZ
mWWCM3mI3ClqUlILHHNF5hoxdLzr2hx49kZlCBP+afyyl1Gt4dzk0egnVoqocdIkinxSxJjzyN1a
OFtnpRTOpJshipgw3znCBWqhEe0IpjX0DQEDRHlxhcF9fDAVBNfEKefKU3kYulL9WpjtUdsJ5s6u
ZalXqo6+jCypoi0ZUyfNMUtPozdKZ/G9p/9ZeQy5VdHTqct3m+RY1q8XI1gKIlr0TDG/h4WWYoGW
wIf2JBOPCBZpsSobBBblu0wcNrwphhtuaTlTGCBV+WRn9QvvhQFVrTKmlqilnEzdSrneYud0nbBN
IFoy/ETogPG5IW2HD82GykCqe0/BQ+oxo6Lml/2O9naq5HLxqJAp8MBcWv7sOoAVVaFZcXPCbCyK
f9Moq7w3sGQzGBNf76iXFJreevBqQJdVoJXJIJMoXos1aAkNcljA8gimGnc+IUs+Vyfzm71LbagI
fOYZEnNsEnmVH3rmzbrZom0kbAKV9BSZ+PPipC5UwDDgUucy5ylh7vsq1v6GjQW6yv9A4vwp1vu4
6pfL2YypqvLoauu404AkqLBd35TbZHSF9ppQKJ+7jn/kvbia49M+IWqQBZorm3l7N1xuscbnPy6l
b6dn78346n3rnHfjKJgVUcHWZh7Q3fSqgS7yjhupt6XvboH9+FKxaDW+SKlX9sQiz+n6/Riqyogm
k4Vgdn6icX3A7IVQWosoRm44MVsnNYglk31RRJbCEaOwba7AECXqtIVKtLeon4vvt8P8xYXFkzF6
AlK9ZEWqrgCFKidAVJv8N2WUsqt13irN4uKhpeE8q+7SSB7Eqoab0fY5QMgEDvxnuwaUXIVPWP47
91B1stA2+z8CDz/Z+4Tj6C6CzcmnIkkcw636i7f0Z2ESp9HjGxGPGPZrTGY3SIWay/RH38EEEANG
0phsvU8ZrjEqDXBCFnkgiQQO53xO+PlG/iDAC50aXySvgPOuifvd8rDZT+9hfRwHb95jOFmI6Cf/
svPQ86d/toWO5mtBXVzJJrVaCuZ8R6gF3CAZnYa/XGFsytVQr5wmF/x8ejs+xZp4dk5eQDEvnbKm
vtEgTILmmix2TuQ1bG573bX3VGjDDxUWD+Zzgl+bOu2SCTrQFW9O/Y076x0rIqOphOrZCFrlZ9k7
ytlCijo+XyRGqVO/1kNdOvG7x4E6WERNZYFJp4T4MPf2Z2aq0DFa6RqaywRIZFNgRTkFMaSqJCKs
mWIf6lCI7eezi6uqxGJBcqA30s34rZ0nxlZFtT/Bru9kI6db24PdKy81Zvd37QNUgT6QM1iUGLSS
lzWveTLYyPMdGPAtA0WerVSF+V1HhGvfb86cTx+8l891WGcQgfvBQ2A5oeYZ4BMgNtCTn4v3MhQj
XB9ohQJCrIFwnaVWICILTXD7/bXrijBdONvPa5Q2s63OFdwOnE0sgrXnGEJ711AZlgWpX56UYWUV
9MM+YbzmOUT2W4m0G0KxWG/6SjyY1VTqp7MvRxfIWSWu3n3fEe0JQiRQMGfrbMfEwcgT+qry4Z5t
ywvSYforT21kAkv5kBdJBG8qdeqERu8AKb9SlPbWFhHklvD8whiXzqfPb6ZOp3UzCHiguLpaWDtA
bRE+fgPKp7fNh7pkCOEyaSDzEsZx6pUDin5nukCYw/XHQyhqsTO1LVavEo3PGhiEA26BoSvvAFUu
uIm6QrRdNyrzTn0MuJZOPLcMOqOfsZxMX0DlS2fOITStHxLPhsCesAxHemnDzDlyqU4Pz4oCwkD7
Uvgg5wvxh4o4pAvB0OnPpk1jclHb8J9EuH7aUB0Aj6xou3/YqPynbNa9fwQQcN9um8aHbvEsPzHM
ShWxnbuZNmwnzb6sXCF7KnJXBsd0V5nSRF9/olRck9jktniJZetvASxif/69cJJRFGmwxoDIL5mN
UWlwze6txkkfkYuyttU9fQg++S10zwUxIMvqKcgDjIothxbppx1LcESS/Swr/pg6WVrs9/F7UiJ5
UtZDwHSMYDGRcUJl8eSSuLs6l583nJREOvNdnSq5mgYE7Xl4dt9exqKT+1Js1s7/876sClvndmlq
t61DxhksWxY0H9n7cgO/kSOz/+wO2IDeOHk7BBi1QdbnBz3xu1HCb+tU8+8mXvJvckfb2pHPq47j
qFGvbbj1PY+EzT85NUHjmWKLJyhskFXwSQIJ9gr5miWLWR9tGUCUkC7UJ2Kbfh83Jg9WtJSSlZyt
Qv1/rYG11mmnGihLAISLdk17XaLqoli4HSJg8HCv+KRrCzCBamKs6RirfS7CyL9DOqjfRq59rO5d
Koou/4z8ermH6wqh+FdV1CuSUes7EQ0TSvYqfbcjc2pMJvV0Tqjg/wekL+oOwqjR7uxCd/J6/Trs
TKIbFOUa0CYjN7hFEO1dcAjmQy0/G+UbeQJnwmD8usZ1R5XswIo8mzvaADJlYg2gHRO6Nu4Bqib9
p9X3vGVBDPUCRN4UdFflz1V+P1/huctqxM8O0gqpp+o7vxUJDFgnPUsUxDmEEvu5LngbtIaHaQT7
U6kls7EA2A4KbHHPHZhkrMhHx63x7RyKix1mXorBlZiHzckZB6ZB20sQGvC+aiCR8sz/genyDaTT
X/x4TUHHVWKUuBls3D5mt6fL93laap57eLqxFkLeNN/Tnroe7yPZpgKbqcVv2Kbz4CclN9nb9aTY
NJdgN6Xy7XdOysLa+7j6mkGOlrMUqiqLGNXbjtNHoL7Jw0xV1pnkFZCTTYLs+6aS4jQm+itBwg0l
98hJ6U15ir84HxyIxyLWVt2U05A2uXy9E8kz33GarbfjP6Ewpjt8IPbTM8Wl6d82RnJBV9yyqzrZ
4kqn2SGUkxTpkkcY3itSSQ+aRZ+f+oy8sZ8y9KteVMX2nv/FE4/LelpGHMAm/Xh6XXAkN0GxYteX
xIlKwC91OAsQYDuvQgDisP8qA9KZ6w93V1+RjMr+JQSdRRUGKpN6gmZFuZVc4eJtjA7TTJUDYYYp
3tXr7gnN2J3z17us3SbJVEt2qxv3j/U6HZ4JVO67a0YPkTo4N1L15FoNSjz8bUgwLISzehKvf+m7
0yFCdirrqyQpccAmBDWTwR3tm6bG7QI0GbGb5GQ6mcTihxKKLQKvNTvT+IfhXWT0bV8JBUK8BykL
gscGudWlgghY/wv7CFkGq6ESY6y42wpx9XA8nvzbAByxCl+dvycoO2uRT36/058L6/9idz+WRUpr
Re5L9Ip8YrX9R+zOYRboME+0LGGEJX56pf/HjkaQJ3lexDT/xcskIZ52o1K/u26yVHnfbJX6gj4Z
0a8AS3t1qeHAciKT4ihUWSa/F2F4u+2InxywDRE8jbiWtvKJ1e9cj9xkiMoRC+h/ndJ5uAdJL1Ze
VJp+nsUSIPxTv4QzoB6cOUIVVfmoTgFAJ/jixSqNsdcgsz9/9Veaqpxos9coU0D8ZSo8mrCX3X6B
eudW2yPoLiDfO4shxWVkwAjHfdWrM2n6glKSKlPm936yWZP8CHlwFtu3p87i2koWDeTNPjApQSe3
t/HQYH96qG2UWmhZ8Cth8uEhF7ZTm7Mh1Z39PDdbFiKMtnAztKkpg6e6+v+gnWpW8hp1AvkXLi6k
yrvpovzoskKVIFYbEqpWDgtd6Oj6FtlzGaHwvzdEqsgQG9Vxt3LqJY35NmjCHzcA//XOZgsrzuuI
36XE4LcTdz7R9NCbV6kOp5pkWlHOkr7dRlCZt1CONwrqJuidzc5KN/i3/0duDBdDtQSJjCJlCObN
4WH2n2pgelpBOFdboyrfdFYGKsAZPP/yq0K3bJnaCeuYP/VConDFvXSda2Yp0fbw4crcHkzaRSTO
OI8K3vGAxTfS5fTOId+gTPcvREqFQ0h7Ms/o4+KuPcbLJTwaHXz9r2Io8UaFugi6uWM0lmdoIESg
cT30mnynW/3F95VJlI2O7qIvAhSBAPFa6qxzOayDr4hUnl3iQeUdPRI5SidOapeRFxKL4cto+GNh
e9EWTh64SLvA2iV7pwbpLmetcYyd71dukCFIPwN3K1I/yAGFk42V/0ItBXxOPKFN5XTU9ayFWCJl
gpZtgxV5XDS4PS5hhKadwUGcoily0MNQgX9KUEAWt/kdo0PMIu4VZOqR+f/dAn9o1wqXnDpDAMPM
ZaLcjz4UBQNNWN4eBp99JDrhDnTBLSR914gfWAm/JNG9xzkTwX/WZGE0lCBgftxKDX+ZYjAxNx6B
TmNTdm/HxyzXNp0MnxYKYfQfBrR5HdHXHgLQMECg//XB/X0moEcgBRYAbhORV/Aq53EMYLpHel2K
4jjX+Nf06zX5Dpj59iuNRlsKjLi58BHWsR6xfiH+pxjumfjR7jJkyPell6C3T1dmhJJynzyWEvvs
EEw9cJMTcHdFlWHZcHQI3lQzmqJ3IRUY0lTmeGxbQWnskx/BntH4w4NVcpUtlrzZfZPS29f6le8F
RpmkGJSVioDFiOJylEf2VyIgWAeJzlB+7NXrfsFyrL/M9+Hu9Q+j8BWg8LhlagNOXJc/8JMYUb9O
q/CrbEb3sMvk7JYWVAQk1174M6uh69oOMo049uuN1Yvu3+zPEqIhsqZwMZijXssEI98sH+8BoP4T
GQ6xoYNt7L8598XWW8LEAXiHqOhmbsm9JkH5tb/pxiRTlXe6BDReh7q1oWFWj6tTxfw80ehoSBdl
yjN+09Hbt+TB6qTJINZZZGaiJTLW916xR5EimMy0pLhSHltsULzR+ukHPJJWg39TnnkGy3Wk1Adg
Pugtf4yqrA6VJkbfMUuvQuzWmbeFDfmqe3y87eDYcYDd4+rn4fa36PeERwucDUTevw0gN7Zktbe1
/Xd8EMTQ7cqzPb1S3zSEAv5NUQgw7cqgg2Z9n5x4cH+I4sr4LJjh6VlydH3AK4FGNjCf1t7ExTlq
NM2YH/8icVxezDjXwHwiyt2KxBvlwwVLZfBYwb8LHkjzUKr2/Y/nBbs2ePTHdEtLY1FAX6rrf/ci
rA6BQ/4RAvWbbPf0qhOqzpHgdCMCVS5KNC5biaq6GyEZWjFpxJStK1GLzSCokHQliiltzQtyunmy
5yOtE7oQ467SqKKbxNhRkY6n2sE8z2Kk2PTIgiMTVGPx8QdFM1hmCDdECH3DrdR3eg288I8SGGnF
toQrBBwCWt2RhoUDNgWyxLaEXQPuBILl+P1gsZO8hRZCD12Fcp91yIiMOHARSvjpBBLFff9ON/CF
/pEttJypO6p0whwCIkpAERvcfgV68aJeQxSdQgDcBI4HHPAk8AYMjTOe7YUXNzHlv+HYaDFSKyEd
tP/bw6L+eYEfct6uhLkQPrXuDrMFTOocv0BDpILDa2UX+eEbQ1t9NoMbltAyqvP6HX3jonpME2jQ
gvO+pI/6+4t/us4V6s3fSy1Co/jmk7BKzYIleAMG3BATtPyTLWBpJe3ClWz5DsuwPyO9cuu5R24v
Le2g75yC69UN+EpC+aCT6Zh2tcN8HtNr4NOfSYwfHQg/2r8EIPfm+U+4oh62gD6MAVSItjzpXS6Y
kx/VPOptyPGN666ku428e51HW+LuGfqwZ5M32TOK2To7AmRsqmH/5Vks3pNfkhcnPCdqj8BahiQP
K+um14hAlyOZy0XkNcLghoPWByWHxffhP/mxNulX749IEltmJUCZXX2YwF7Icrey8X7H+TXkAlmR
+efzlQNlaui2VYlzg4vl+6kAEoeodCpAZ7CyMbqQe+BwIr0iY2+pB2zvuGUetL5sRKDx/FQIn7O/
v2S0EPZUtHeNexlcKrclJgdhk2QJkTOIdF9qqeH3neme24klLlj4xGDzpp9Huwu9+nBX8Wl4X33V
1S2XyfNC3QK7EgBjlTj/hfjMFXGfr99W9KCs2mIMlBkQBWkfMIDoJFn9fGL5Yrk5h7EZGLauBmed
m/JfCg+C1gsKNVH6O3j0i7odISFJCSdevzsbfzKgAMlm1Q5U0QlDiwYT365+a45LqlamhuaWAGgI
lnxdH5vXTIicXzHfKysoqRKclDLmNqwmFYRPWTPjptplbnmttxX2LLCOO++EEbsTzq9TVV7o6Dpv
LVa4cu9JzB8CQu8I+aglifftuKOdfjw320YnwCYMddvYytYWIPYnrZYw1wKkcJi3E3vBaTO3sBsG
WDF61/rWCbkEiT1svA23UvTofgk0gmvsut3WHkGYXRHSRFDcfqyW/j1yZGTtTK3Td3ABMNeDi3Lw
GLPcCrxgPLVH7ePhn0xkQoSgrbG/nIm/CeIZXo4IJH9n2dwqhF/hK9SaVPg50TOgvRQIsMowb4UX
jKBEelWIZs5aCnfOavq5CGin5twfZoNT+3+I9/U2bh6PjeoAzygnVgGgrT06sz18ukjq0inEgd40
PvtNmyqlJUAXbcy+8KZ7s1R8mpxpenSOijnUdozd+sOgx0OOX2KTy3rtBs5UyPAcKkhAd25T9Xfh
PmJ66ZOhFdpewzL7wglPVDrtI8tf4bYJ3iUHB2PCSg/0VpEfjm8nTGNYZvS0SdVqPni6qx3KDnsY
ySszvzbkkFyhElxgxqqom4MOSJJVqitkGoKXLIo05Q1GlcTlo1BV4c/VAofQ5nKY+YPbmcBwncQ6
+VJ9q1hP1GVy8kFGEAR6gpu+fzCsl4BEE4hEhQXwun+sehfUSc39+hsCPAgz98M2458nfUr6fSfH
yKqPSZwgyFwy5cvGbYpCQVV5AnR5HYur/mNXo4G0LWJNm5D/1uMvwjUA5IpZfcb6nCoI0YqtyVxE
4mrEK1e5cxQJEHwC9Vz3sHWMZOixa6se5zTWIaXAPXuvpzTCU527frOjCbGUt9/dkbpxC8mFsPf0
hMPJuwdD+zGL+HlQTwyZxsz9FBnHESX724ZShT9eczkgVwfnhq+E6f7wTpNGQyydLSb6aanulbSg
RUDxBRmZpG4ylOY2KBqR6TlupdaFqQDjnALNi7b9/GsTgLkU4hiuktUdd1idO9CfekpYTfK1YOFk
CXTjrEAy5lVfIPiYjUu7w/kh/myxObOxdeD933RXyuniRY9OurclAbA+RnNRxh2dP90SxEoKl9RS
cQX3l3zNzSW2rytyYNTdMpEm3aFKDYa7T4XyPUrEGuSyLuV8qIWigewe2+0UxbxM9F6PX/IN5IJE
5Osi/My4LylchShQByhFQzbYp7KFUSfqOA0UPw7HdbVOkmPUL3RwcqNHZ0LlFBV8DtZbSlMX2nDn
n5RdxgvwHj5R4MmvHYt/egFKZyIWRveAM8hhiaBv6l0iOOM3TMV/CiXg/Xec6MKGDKIgfoSeYRk9
bwd8yeS2FnJEN2t8uBBcUdmypr927LwZJxb963nCjDrx3H5eXliPz9AWvFBF3fn+Ll9EJXT6oat8
ZaR7BiQTvCduRk7/pqSpJpErNkBs86DSAVnilEFXkFVAPnxtcEuuQD6SsyPrzxX/jihZ0paPrxIr
f4BNFHiWac2N2CwJYYoKyRV4A7NRcdusU4BMzTbRD0FiPJTbFfA8AfQZ5Jo7vgOLeLL0BtHALEPu
CKVYyIs47XEnSSo3hIwMNqNXjJTclwFP/KebS5YGuGdtTiEsAEinrSbQjBF42QxqE+U2u+psClVp
tbtYipqwAkFoHKU/a5Ybr3DJDYFkUIGZU4TY6xeUWSIKm72Sd8EUFtDwxJbSzTIBGmK+WysLXdhW
ZyEs5GVtJGOE6NN1YmanxQotJHyVlxlYjs6bc2d3XsCt8yQXl4bfBw2I6UUurHNVSAxktZ4HMxO4
NFAUfkMjhUCNTMIF38tuuCjfmRQ1IaF2gp8/sQTNb17I/k6XQOUMPpdwJ8F4Po/C6PX+2w789hgt
FVV0bLc64WrN/F8r2AUkYoPF4dB9ehkTPOcfI3TD+0/xQolSH7v36jYFJY/hpyj5vUZtRvv8xjGw
sLMqMzVMcNXDZUfhc68rRUU2oweJhHTjiJx1/dE/8lJ6cYqvj/GrCusdlW4iOJhKrB+2wVXKPRP7
13qDsj5Mdi1mypESSvls/sehLmXKptAQlYRzWymtjypKX3lZ+fIfD+lDP7+1OIQU1g2IoEJRQ6cS
ZbNZ8bSC3Vd032hCRnuCbD3XdW+I/Y99/pcKGyGBnf7GLwm/qGrc0lJhlJZFdXF6GbpLW3ZXqXCi
yLUVwEEvSH+VvWwMeAgu8qBBtjIdJC+OLIzN+7obcMUFAqFfozaPdlcL+1ER7FHlQAGvDluJbxua
Us1VOlefin9+O38MT2KlrQojwazpXyuupJOUNJKB4j3NrmDcpWJAO19qEWW8rMhy8afYyIhPzXsk
kmf8zIOOrDdHDRa6YxuyAnExtBQT1LaG8+knwiw8+OPivpjCBS/8RvXrqyJYXr1oUMbL8Yd8ufNB
1cguGoJZplsj3PDQfzfhcgoOOiopNA1brizJYiC33txN2CqGAP+otEFybQ+ZA1h7mJIP4K/hZDsb
ENajBhdI+yfUmjeJFFXfUw3OpCsRRA28i26aFgCgrJFm8/pnCGc9hdNlt9k21zxZwjI3ev6ywIXa
CKEZHYGKUP21dNWVXKcJtKMghAVQmKpT6Y6lz6poq6AKt29SGG0X4dM0CH5GW2XSVpUrTHjph6s7
SkQg17k2r+3iVD+JVn3fnFillW8TYHR30T0Tpg7T7awKbyK6J6ZbtedDOorES/vR2fbyzrmzBA1s
FgBpxea/qYYm84NJzSU8l52RjBHsuQJVHTvaYFCeQHo3QnTKU58BXT9NQcRi2pFGWgaN8MwXQBjP
gCtKM1rE6XGyts7J4QgCSzhoM1Th3hgYuG3XveuDKFvOT2JW3EZrFM9qhEZrMKXgaBfVeHo82Mei
8kp4Sy7KRuZD2yP+xzGzEPue+hAIrLu7uM5TXJ550dW9ONS866v3lfKTo2MZe9N3DkWbzzlT/3v0
98qYFhih3av+8sg3E1fYQy5VrstZOYh2VfKde+P3KZT9qJidpa+aXdVVsm6HG752A76dxzAHXpRR
mJbfftA8OGIXwozYQQwWhrrs9lQXx62ehkGtjnOar+QwSJfQ3SzCLkp9yGn+foJkqre2bxXTmGLW
2TyajEUQ3Tqkj5knhm7EEe99sYWleiY4D/1UAT0J4sP+wI0a9ZDWyKmCZU7DGd5LX4/4kF0Njnhf
H8N/gbChLz1dtlMLO8/CIOpKIvTdjFVt11P6ddOGB+lifKsorIARwxgZ1wQL8j6S0uAShJ0ybeyx
fEE4R97k6DvQoWq0Ea8WQIwc4li/9+QBBDh9v9u2ZVrSZU+z28VAt6IcNuGnYBbmhsRAq9UKRYTX
QA8V7nVm7CGCyIdgJJXJM3zX1NN/6FRNPmm9uPx38p7/A+KD78vyaY3p/+a4BRP4MaDHk4N5fVMZ
uMfv3LnjCjJWiqqgWw4ssFwh5X5MiiCMwlkB9662PmkbP+opBVI9ogPfEtSs9m0kLLSejUS3JEBM
aLptojy0S7Gx7ycd2q/gKOAUj2PI30Ht/BUyING0BPHy7n6jaHh1XOG1CtRDukOdEwWSZFXdS2SA
XnlW2U5eq6A9YQu6cBIDPV06QypwWVnysvD78XQ38g3xCzq+sV95EmmpuRG2bIZdENHUiFKOFhNC
k0zulIgin/y15Grlgu9xWVFsR9OntA5hF5uRCrjzmLBPZF5uQl5tNo6QnQ9/eMvzZPXgnxYOckqE
ZyUWIzR7PcJr59qhjIUkjOd3MBXqjWtSxXXr5pSlKUYcqmA1PyXF/NeJNQdKdCKHqzE3tPJyog5b
69rMI4vhJqy8Yt8lOPCIu0iW+U6R60wpb7ei9KSTjNF4GwFbLfljsrEU+AB7Wnh25VtIqXxUg+5t
QaEOmQzlN1xJP66u3/OE5em09pkgntxrq/fF6ZQpMDfbNNsv8CVQBMbxOiZGBw+vhufrc+pKC7QX
LY2aYd4c6yXiL58l9+9ADuz+b3bd44dJIT9iOQVthJ/4yU+I4/Vrs9XmAFkAaP6X+DthBr8cWt3A
kE0b6yPnQweVHtsDEF9tzEeWh4ENmoMoP9cYhRZLD8NhEy/vi/8R2SO5jzKZYkEX8cA5hsSaONkj
u2i9zb8tkleyFszqlK1JbRRZeKHqreIDRHtrUGYmN5DN1gkqOeLT7Ci+mILYve4LeH6BDlrPDUaM
UKWh95BD15GZ8YGwoDP0uaQtmQar80EYJGlSO8qb8unXca0IyeOid8j84JfQi8+QhY82WXcRXKwo
xWlJE/tTs3Fxc9cQMBrd/B9C1NJNAzfwpplO5odMNLigTEsCcuuFvjTpDRc4kxOVqSKPQ3ozQ2Wj
5UvAC3PxoQI4plgdjqbET8RFGRAEpjFv6KhTSR+5gEWZieBkxpYCCltwCTocdvfs1FfVPFYSuZTo
mbL2u23gA9ixUw9a27y8iItGCFNkU2LRvoiwNGIyILK4+tx6ARE9P9T/gJ9JgJWDg0ar2OV+WQY3
mN3Z8cAMPR27tVKGhG9KwoFjcMO6WLeseftmU8ig9AxxQWSYKdLWbId/oFRPfUL3XkSQKY2jw2up
4Bh1ZloFf4Q9wZtBTio13cs+QZ5TKM3JW6XLgG8XyoKnD753rdiKCU6oKInrcNBTC1qCxRpVgDsD
unbbZdgPW2HglBD6h/l/wsVDnTqSZhmS9HN88hFbCRS/vUF8nAk4K8q7+g3p6Iu1ZBn4X+bDg0XP
HygFlJ2mSTDAeqfz7sxCSmQ0dQE7yKXxdN32zBObbIKoTHGcLveFeUGxpq2PAnY7Q26SWkUxHFcu
vgCfpS7nrldDhzU8wiIBfZIEmxchIenPq1px/2eHmqs32uPOxsSlAb7cxV9Ib7E+e4ETez/0ke3F
atPG5Raf/7aeF2f2pXUY2/WFeUwBzobVW3VWKrlrHY4nEG4YTLBlm6qt3ehrmJSQqTyXU0iU1LLC
wZH/9sIeBPup3p0P2q/InWG/MO1U3PbzqCM1wtI8Gk4BxiZkJQSEEayppCL9Y1CjGV35cmTSqmf9
b6X+8z1G7uHCuqtbjcbN+Dt38rtdLY59i6QGImcCb4Bi5Z/xeh4NcoBSXqIN6gqX2myKEF0KR0Mv
00NabiVc3ZNAva5LD6BtjLUIkvqd7MLj0nLQWAe5qvdXpTyn6iskQQVlaQRsl3xb6rtTawhztZda
xTb08S7XmnA6JNxvzkum+mP3yr8VXEQzH/rsSOEapdkQWh17To7aYvJMSaiwA2QZVqUsxxXMn9FG
iVwkRqtW60RdacPP7xPSa4+yw9AAf5ulcd6tKT9NW6nKr1gHDTiryb2D+aqc8IaAFs1c4QNKCXhP
Qhc3hMlWerOtISlDnwB9D9IPi9Px08JvOBrhs9iLUtAakssRe81Pmvq6f/EtTp7E5ZAIoTrmi3/K
HIQDPsFYkfaXFqUKc2e7K4sxdmdFdRTAcvRCBCnToYcVEOj40vmqwygQiyo4wj2pXdcUs8bZ9qq7
8bnYUHyIHTvr57NXQ3uAD9XudN7jHmK2Ew183asNzdeGZ5lTPPD7ENZoRSCMA+awZwFqWIjjf2Lq
T5rfpf7C8Y4hb0jkHOw6nZeGD14cBe2bS2Kw0HGhBnOf0s+r3PPtUOhBTKvmZB/AwlpUFi06S8bh
ik1+ygk7klp+6hY0Klr7WSf5RA9ax/E4/+g3xx/vQLnkwok2WTErVYJHHYtrG/tn5CaR1VAKvU1m
VrgbHjUNyo2VGp3K9ZsVRSVIqrmFJVhTmL5MCzAkPNz5Hq75nQF3rOR+YcYAwxs5R9I58lY2GJi1
gu2DDW0j0/rvtBmIWF9Jnu05WWRpEzm3BMN5ng9edJRI8hitFRN8LiyljhlFwoBNfD5WRDy5qOvn
zNL1EpilBKg+OzPPpQVY2qOYVf+F08O/+oDQlZPhwPtjXtCdCK0zqrqeKSj4wFn5riceImwfoI1O
gWRBmvLqPOKtMoIEa+CtINmb+7TYhiZeo0HJ1yrUYVjaMmZHXKhWXGJ/QlonmzGQwWlHFDr/xnJ3
4FXSKlmrQb2oglpg4YBd5nOVrkHq8hHoDkmwPP3FgUEb0LNIv6ULLockhalUVTD5s4mP+GMSIzbO
nlSr/glGSt+IIsT0t7lqx7nP5Kxn8LcO3IYTvevMmnDYfuFEaZM3XxPGYKcGZ4np1JNxGJC6BZE8
3fe0DUX1ljk5cY16s/X/OanEB6BdURKwg3RrbtlowpBi6ktpLr7ksxrsiv5GNBBzY9TK2jliGkgk
YY9WMST/32xf74uE3SmHkhoHH+VSZenLPMPmdEgv3e9HORrcrfAuir8utz956Wcq4FKw9pRSyLVy
8UE9FeXAI20xXRM45Ow0cjzVeVSykad2xlYlQO50NrVqywP58HpqDdUvhA5iIx3sAlH9kECT14VS
luKCCdyh9sdHkRvuy4Sa3CaZB5Fzbm6HSmVZNMczaXJPn/LWnOFEkvwP8Ky3NyiZYuGRWck1Ylh3
K9LlxA56oMi8bYIQrmvWNkwpGkWC8Yv1ycW+mn5j77GqCVH6PjwgtsLKhNTvpsCeqkhFEzU3VjRY
byCB6i8lWn4q8ViGtRank2diIouwfok82hssvOf1aNzSmbFST7yjFe1XPLXIn+J8qiJE0oIcwgiD
mrE2FADAjQYFuyxZD2cg0XmAauoiO+8YHi3Tu2tACB7+XvKSQRjWmsHkinaQZx7sbeijzuegGnMh
N+Ubh+O9FIxtMyA3uE4ATiSk50Y74jysPszx3N0gkys8MjfxPhdWNIoe+FtEBm08e+rCDU1Sl4fA
3bg9F1DGpzcLF4RXQXe9cPIMunZglHUhQ8+QonnDCNakfbI/2aLae+pns3fc2fRBqsYUH46woaU/
NSSM9L80DCG14JYeU4rrzj6N8wY0mzygCqCGf6Vftz0rKAQ2OwUD5ehtWgFowZMGZpCDqvW+N4Ta
bVyiXJ+uzrpkm0S8k/elqPOyZhAJUTMY+4Kvb25A6ST2/Ig3Fqw/sK2NPksMs7kxCMWkKXhak1nk
xvYapZKidmYRvBLgbpRLl+qK/h5RYAmJKHdeEo2+egKr4KUsIBKtNI3ci6o8vvAk1OpscFIJMAUj
cWCHO7k2rOyGcPaMB6c7F0ISpblSe2Am0hWICTceOo13hXQyHah3Z18yoGATVSm6q6lqakxe5fVo
UCukgMSMgGH5sXANB/MgnJqFdIXomQKOts4fQfrSG3bdGLmgWSd28/6WLAF2B44TJnka6V8iRKWc
iK7lpd1vvKmah8csQSUInWcj43sEhzk5ci5XK474wNqP0cL5eEnUvzb7EBpztVg9A5q2AAsWkSVG
zn2yEWA8jgiVNxSzkh/oVma4SZz0/yZMnUhGBZrp402+uQXmMxuFrdjLtECTRc5rGe/pUuzvM+x4
BtjbJTh2XAC1gn6VnsqhiQMBcDBKoayS8cWJMsIoNL018rUBY7FfZJ9eu0zrsH8e44xoTDHHV37E
nw0z8pwT4F9uDIoP6K0EUAObhTXXfUcDWLSwsy40a323j/w1fDeXQ/nFTPbcT5PB2Iu1ynQt2cEr
78ngAcAsm4D6NEafp74eGT0Vyo1bJq4xN1rMEC9hMfRHDj0LQKB78exl2V71Dh1be17bKYZ3Kfjd
+X2HqYoR08Iq+3AaLWLJZShQ47qxL5DIfVoGEQ4xPkx9Kxr6ILGbFpS+ZxtDRHgUkSVu94HV//Gr
hiUBFmE+Id0dQZO+ShCVLVLWkqDbOsXfYCPVocdZukyyWvMlkYOnblvnqhNIpUzAmaCXzHJHg8On
7ymhysccXhClCXGL5r+cds9ZoP9GjunK2YHQUPYgDrkraMfWOnGKv9759IP9JqCFqe/gX4D+qHyZ
H6dyfOYy2ktIK3BH1K0WCv2RXoaPwdebdO6sKnQ6xKsEEiXRX5m+exXYlLn07S3PBaWBeljsjbNl
yE2LHcRJ8Rq6sdbOjMnJQY3sZF/bj64tpm+4Hsu4OjQ6ZplhtvSBcwFf+dZr2bRo+inPaGDSjvWG
1cHyCOnNJIEi45EX008siaeFrM11qGJrQTLmZhL62fpmMypwydV9Rmyc0zLdSoXu/HDsb4zxGd2p
DUojcC6VBx+VxAAumXgrXAne8zFXqge9tzbRNjhWJCr/jCSGVKMkptPDFi6PiL1p06piBgHczetB
tXyjLhdHExBqIsivpJHo82BM5eSSYX0nVGmRJU1VtGGlTYqrkC6D/+2C3BIOvLWspiv04/9vNXbO
SkFMgzEbzuCx0pF1MR+nvPut8vQHAOxTv7APiAB9UwojTC0DerRWJsGAOcaEVkGPY/X3P6hktt1w
aOU+OJG44/8KZMUs7NjwfW/X+obv1El+N1W60+gxIvtuzwzdWzo3WIr+6wb4Bbrrx9bxU2ZcExpk
vKbcPw5OX2MNZnVDz70rptqbW1tuDLPhNegZIa00n7PL15gsQTz2UPqQDngLUaN/R+uJU5oh5zni
WHlC6fVg2v/GV6uehguAaS1XgFjdLUroBOdfHFkpfHX7Ys/PlIb56g/vFaZWYnsmmeqb1s1s6kIJ
q3x31LSN1X553xius+/MlHE+VWz5UEDXIlJEDBLudSkIUsGKec7bKtKT+qKDfzcSo+Ro1AkQ5Qg1
Iudtj6OyQrjfXJLPRmUPbwETtFj/UnV1xiSeg331ilydLR9cWMRfR1kMhXMRfsb45AZPiKAglWYQ
IUqf+Igk56D0uHBzKMEQRjT7RpcdddGQbJH2UMwypk8/0LyXY4cKhnbf1M1h4FcBJrcztvNyAmus
PTp/ujZVT59QWU7WFoIy81bLc3lmah0u9dDm7jEFYYLNiVvuMdDKxikxo7JoZCBRS+xo8l60O566
VdwM7Fby/QyHpPwJbG+C3+3/aanCr1+HBotYCJqzDd+XZvYw0E+rQGg2GsOCss24PbGOYziTgfGw
/TGY13tr0VRloAQyQjRnEFuNHmUMRNrw+oxrLNC3fOYgquIwd62qyyV8E9z5yzwhTwr08MnYLijj
ApsonibPiT/Wz3QTXMKoQR0QLMne5tmkk6BxgmVPdoYdrJLNes9szPsXhdHxqkLYD+dAX4bzj4uo
sguOu2d+jsRD1xnZo1pKK0HSTr5jWSW16Wh3I9pNsGHREzlLHKe5JQtGqe4VuB5bkLQybHIXLCLP
1SqlBmD7ByzWd+c/AET6qKW6LsBdUoQniwlRRFu6A/gxwXMUQMJ2NGLM6zXwmCPKFgmqEU4A7H9e
lzafw2RjXWde99wuiA5qVN084W4Kta/pWWORMf//CCuUcxti+bOEF6ZeG+ZjgQIhQZSsQIUKs2lP
joKh7nhbgEyqBQa1yMQ5hnqoeN3Lr91MuURUF3YzNmQNAmQNpejBv3SEUKj7RkudAbI+Xw4nmP6v
wBGe/vgYJLzisyGdI3VVjL0gpWWtu9E7J8jwT4vfkRLX5WfYuXsB+OAuz/oZz25+omg4hpwi8LCE
aXh7Iu22nTo0lbiL2Jq9FIXTtXubvLFGxdKw2fGrLTmimrkuL41Hqlms5CBDW8qqOF7LxiYPu1RO
TWiFBbgdxOg/wfNn9ohOKHGEAU8H2JLcs6eDyMLELYOg4WTAiBzFZuvb9YNHDWe/aFq3Tl38TevY
P/cvXhtKCM6uxZZeIRf4d3lo+lM6HbtfferbBckf5RxqOY3Gek91c03N53uHWs9+JZSNbaQ1nsSa
fFV6LEsTEM5qIymBypqchTy/z0nWfhS/PjN2vUhCC9vCxneS+mjmxVbnkQ4XMEFD2XQn9v6vYB8k
3ZZbGPKkxeqBkm0RH77NCQy8g3KPDtDuT0Y+aWabuwV9p1EDjJ1+djL0/KnjAxhXvJS4uPIJIeQX
xi+Vxb3BUqT+0vOUx9AOcDW7NZLuZUTFS8b1/3USr4FoZO9lmYSd3AYE69mtTFFL1Qrwt9lQmJpF
cJmy85Sz2DJ48vBHqRjtMgle6uv2tIA2DYCXQ3d74fS3Sexhre7XzasxLph1fs7P/GC/ST7irV8y
N7Ve11l2zadvGsuXAPrURqIHNyjhfQFVR5xKz6srNC/XmEbT/2L44qetLlCDRQ55d5I/ODYQyXvl
dEFofIUsgt/lsIfDadoCfiNpRZzV/sTw/iyiwBzkynsGr9scdqF/ha4q7Rn6U2RkgkjxEHa5o7S9
YeS1y89LvD06jpEhgO+cb0LTPr0jNj5zalWTa+ov3xWRuWZ4PU2cLzMrW9lgJZ10tanh0J2cS1/r
+2w1EmKpXzY+2jRtmW7NU0t4/Ia8TPruZYO+PmQD2hEAlfoyk2oURYv7kH0s7G2N0Re+iq+OHHDC
ZgK51erOQpn/Mwq9lPFfsC59PM4YdQDxWUrnJdGZneEP5/UpZuw5emnsRUaLXJ/edwhkC1C7oGAT
AEh2tLMPsOVk19eKYAviIa4ZZSikiHf3aNQJWT5U9K3Rehp1PnECrUGTizSZkOWa31+2tym4iHmS
0maBjrOrD7cOq6BsnI0+036Z2BXJXKsOxN/xAnTltQue4yghiiZoN+p73pe4ZXt9h+czmbinqLEN
KD7wsJYj0AoYa3/9BxvYlEG4DWer9Q2/zS+FFQ12GYn/C8Yf6Hz+LaPMOKvCc6WzFf0p20gBm+5q
zdeAzAPnrpEWDh7iMFwHt0PjkMcmsYpKh/y9848df/scUJKxWsdgsZnZQakHErhkV4LeEu8Syt9r
6SJuThiMgJbCQ05iMZfCAsGTn3TUVtmaS2HZEvA9sK9CJfIGYCXsopHlrRiJUDpjEeArnwnEFVKA
7NmkqGtDm72EP41mgY1jWABfOLh4q3/4IdvzgBow28nawws9+16f+0POFflxTTGQp8O1m4gvm95N
lbMAwzpH2+AkXCcBQqvgSw0yWqmMPB53k51m/Md9O5YJHyUvXHiXhtiHdko+9J4heH6h3dCm3BVh
m7XOEQ5H6i3I7dl7J1h2GUeeEUtnihfWbya/qrpCt8RUjXPbxASArkAxo4UOeyEon/vAnJKs/Kt1
tKKIi79kVajo0IsVCzHItx0TpLOv+1t87EaK2IJcBzt4HwU5/euCDWb6xHugcRE2IYYmj8xI4wnd
Pi3/O8fAbAdwaTJ0v+8s+JHEH9bna/+SUSkTIPrdc9HL+9pJxbodHz67LZcrU0vinW+hpV2VSra2
7Y7rAYbwbJdoNPaqSZ7O9RHtGCE93BU/xgyE+suAyu0wNnl2AGUvrtXcA7bbYUWoRX9aADUBQYGz
hujnZXYHOWIpsNpFIuK3gKURlGf4OYH6mbqUgLkGIG66foaQZvBoyYZW4y/SLnoyyuArhE8jv6j0
BxIgJ0iV0b/gnozdJf5/DEU66mxVHLsXyLLBUIhFN5dLrhHx22WUWpDuzPMQq1fVZiRyI3i5+3Sg
YwZVF31aiALdVzUn5Zy3HWY1Wqto7mwJ9LxYTor9yWbpSgyUr1SgX+xJv0kE1rWgRkbLTlByet4m
FlT8VOzivEoVzJPgCImjg/Jztu8nZQ7qd2cpj9CYQuxoGEeG7fuvyjZiUJY/648iKusM5W149lf3
gKBl+oFpAYlkfSwjZA/33MjLFVtLDfv59tKhn4P8aT5A4znwiPZvceM2BhShoMIKi2mqV8cF9lPX
8oaTzm+W6ilu+U8kiKdGKxcjmxkZcbhz+I3LL62WX5wNT9PuLu9ccN2ZWrZVedmMMkljWPf8Mu9V
D3tZvMjRL8xxjGChDUzHgt37bLStV9q4CWzHD0mvSYs+5ZdUA//7Z4vNQxEItDfoWajvdbOrCY+U
mcaCgDxAhw01JX56oJA0HRiKg0v/QcZoYDiRyYlCSpgIQSciti7ADajqKu54dKxRMc/hL4na54Zy
BQO3f86haV8vVPmmmlgLJpRpbo+5rJbYQFAzJlIXPuog+P9bY754ryf/w9XvX+xh+up/zm5w2Xec
RseVI1hY6QX1miAFE5U53URn2Cp2/IkqMgz8x5nNb4qXGgr7+SqFatXvRZjAXcKcW9UxTIv1ayf8
ETl/s3UqoowPS+60b8WPJYsZK8LkIgcVAg91ZlyTmEmKc4V31bK5taRcWng7/zo6buI+6nmlFoRk
kbfCGJo3A6DemJFeXy0yHMg1UZl0bNmVCifXrrilg8GTD0VHvzKdYkNF6xDaABgKDsLjIJpHaZnN
12SkgtbqQuuzPJHgSV2yLuoshHSjVk3IvTHY8IgbIgR5RgTp1v3JAxm2WIRwUAvAwwbydYCR9tq5
k810TIngNVLLAGfEcd1Xb5ro0cFsByMzwCAGvdKO9SRWJu1JS0tm0XsNero67o5JqHmaYsqKOZTg
uCNV84QWp/VXzvGjsJhOeTjAu9aHRhaX0CK93uN1jYH+BuPdZR4ieXCoP+C31xNiUaUeK2UlvkU4
/S+z5RpY20qDbNoJ3ALsrV+NmwifbWDQT6miIN/6r8YUvuXT8HiM4TJIJTwbxOgXbXGtnhgv4NWy
qyTUpH+daUpxas2qXSD2/coQ+UR3yRNiH8upxOLAo8D3VI7uRc9W83gdG/xlElvQ1MASSAX9BcLr
yfu8hRru8SJWJnjNMhag3f8bSLcDwVrkP/vYcDp6i8wpbaPmW8utDTv7nuLGWY9gyjSPXhZHCJRv
I0SmBpT48nfclHlqrI3pvQoRoYNg8lMbEkEVq53TlrT1DEDhuVLdnJyKWB9YiC+Wvl/Awo3AL/gL
3wQHiEnlU5NPcvFjKpbxH70m/2qNzd7fY+PYhf/X9TR9c7dfoVtdobUholVWAVGowM4hWOCTMqFI
NXT4b6M8AWNq9DhCeP64GSZDZe2y/66CDLpv1+zV6J0pX5PoAn+/ClG88mm0WOywhNuvqJI7CUrw
m5f7YebLXyI5d8/sy2zB0XUJJBAVbtCf/0t6ubU6oj++kRBju1fuirTiJDvktMh+9lI9VhvyXRm1
5k3Hq88dwM+bIwvwoYAk4AFOLhJcOzAdeKM3PotBAv59zBDHFMqOd7KaR0wBvO6rWbHav+8MSiQe
Uxh/p6AzA3UBaaG+tK9mcH5e9/VT0z5cL83PDvuE3XtO0IyUZjL4wfNlFEBcnz+GF2BP5fVTFICB
JvESlmAybiGTwYpO9sO/S8J0pOgVDB+zGYED+XW33DP5lS59UYarV3NPyn4Mp91CCgkjbeWoL3VR
0Cco4oYkWw2rreT2ygIN2LGeQ2uG+n7RgVCcqF3gXk49vXslaWjfCdD3zSrGMNHESZvM7htUCBS7
ZPZIws4qEwhD0LddqWqbPrtw2riPd09IrfIfrx3hLsZVuv6sZET14/5MzcKGBP0uxBv1CZ1CBzgX
LHnueyuVqjDcbzUzI9JeeSo94tjJJbJZsBi0VNcTrEesE4+YLLbHqf71cPzDH1CMvRg3IF8pzMRK
rufKwHe6MxzH9G9uoWc5MxMDBQIYiYo1MNdSinsL3uajrErUVRdYzKBn/Vpq8Gdn36kZyWj3IUiZ
dCP7rpihTHIKYFsWIugk7seywNphHwjuOCKmbkddOdjdYcCOl22ZC+73eK3ecqJWe/olmx4jgqUa
usxQ84+UoECkuTftkqpkyj/MxKry3SSnpCXDLs0Es/mbjF0f0ul54TDVYclDCipZG5N/R1rArc3S
q56w0H0KX8+JVpKHOwgZybAj4AQ8/rK3bjm898UGNfJmYyY7aaFPj8JMy/QYJNbRn03xaa1H2486
0qj2iPguQtVoFDpqEV8xOe2xFH926LvQPnY3+X64Rd47KgqIA5ACFUw++Nf3qxHsijzmn8rL3IUP
L9mqZqV02HeHj109roQobghBFjB2G87n/vXpTOD1mtmpIlMnXb5arfxCCMO9Q4xX9wWQKS+W24LW
TKacswtNH8MLkIHHghO1AOxMiq673CTNsG4fMhD6qIiruCKFobPgGfmx8w7dzQjQ+wmkySHBUngg
F7VTU9kwgt3tXricXLM5fmdA0tGX0ydDwmDXVcuqY5nT4DnLY7YNelfxI2uQEaYUsA8ipOf47GuS
p+o4/LhAOcmvbcu6vtSbasSb061WrWinExqK8yf+mkfgViR2JarT8mrt4NFrKUfVip9Kbs2qPac2
LyQHl1ACc3EwsqJ7yZmSuZTHTwdgKZ3YdO9Z+UywGafpD62HeKsTVtC9BfK+6VLNeYvGzNBdTSg1
a6Wg8zOWjwF2BTZRa36rXjry0Va/5jjxRXhU8pCIiM0cc76dV7INBGdkqvf2MeBgdOJ+2qrzioRH
MpPHzfd/j13jyeyb1G2i3eJQMdjT+aKk93GiY6bz2EcGwjxkAlX853bomRUUPVi0pis7psZ8LZQJ
IxWuyitIv1mC4CZNgJ2Bu8SE1jOfspxuOAlvnxmtxMn8HCUSW/NE702RPYXRXJAw/Zg0ApGbsA7T
e+WJP4b+1zyAsW0uDqVnQfXCioFdtjElIX5+gKHbuzKel4j/4DoFrBfYZ1XZMBy7Mxk9Ah84GKCi
yIgDL3P2VqZtJUeas/l9jrByS673+QIsM42Z7dPvpot0CdZ94ewqqHUZWydi3t/zBVsc4VxPcbC3
0ROCE4aQRiJxNNaxFL/jXFsx4qh8aWZJCfs/Z258BJqfYUvurrk77XepcPhQ4QIs8635ohrbtG49
MOGaB/JJtvhFUGuSP8lD4vyEoAy0Lk1DoB+b6NbsfChfNUFJo26OWfOLqOuV6W75RgGEkqBmoc7t
rheb+Oo6yvQdHYeokEbcgcBl50Vrdx1ONrSpovuWe3w+eJHkRuDrYzRRk2rHwh45cig6sNaCtieI
GCeQ6GXglHWL2Lic243ATciJSzR7iP/ENOKQDKzUdUisNOe++g0jbJYrAvoWOSs1aD+uLGgZ61IR
9snL4205vAg3MaTk3lyJAPONgE1CtoD+ws3lL5HYZyD8cQCVTc0yl6oRKU0NVZtd0X2zulpkv6i0
P5NYVO0wA4CRhwMzXdS/eqglbX6lmSznrWStmW7BHxvRE+qpgyOdqmmqh7bztmYfzi6WqZCs97HE
lJLE5YOvAoe/Mvm5j9yrSo2+oiym/2HNYe5Hy5GggikRL+xbpHZxDRB+2M3fuqpAsAfYg/GJwRDV
SfVS2hVJgvyqNK9uSV1kMIG7fFc6L0mZaRC1R8Kg7kMJOEcEdBga00KPcCwArqG4vYUvd06zBiWV
sOhbSSqE7UkqYtZBsnNB3+gtCSQswMznfBrazGbVKFRnKzhEOalPXTp8IejIcOFH1oWJFSuYzDEs
ahEeGLVkJdKxIFgi9b6qYUaUxS4oImuHW926GOiWynZ+rHMMZ0gUUI8ghgD45CP4WKWidd6FRrG5
+vf81wdqwBWf0kis28U/I53uaSXfO5XOXjHkq/NqjlcSPCldrseWbcD1fOwTn/2xwRhzXWT5fo7F
3RcS7n2pzcQvzRnBfV/A/jVKNWXU3nBNt4WLbHJGRp+PkaMkJn/6Fs1njx3j/XnFnkhHhv42kyDS
fe95D9C22zEvbbQdKkLjx5RKEUDT/lc6qv+WlUJrLuC74Pg9h7n728CewpA+qxPWeSwo/GDBXurL
jKACFcuEeMbLiFnebwwjb9oMvHtbcQ7HkYpl6hCjTNoLGoVyki2Y1F1BFJz6NK1VRIH+82IYjAy6
AqHfUuN+m26QkKLqqEOSP2qVExooGBqatCe777OaRP/Gw5gv2QZhd3iM6CSXTyicMs2cnqDW+G2S
x+aN7pVnpPB1jTK0ATo/PEt0hCZy2syTdPZOG5IQW7lLHnicloWC71czsw2VWL6OJhbGc+sIQTLI
Iy5wHQjY+Y8b5sNiaID9Zip4yD7qe5UzbLLwsVIATnvoI+8aTCjlae2Hb4ha/nhHNb152XfM4CAb
ebSt6t/qCcoCgXDxmH5PvVUhb8AB5PSPmiQN1CuEUAU41x0kh4x4x1p5luq+IExL15OL5KoBvFtB
RXh5+Rlps7LHhEB3aZxE2gH8/EZLkGyNAmW1mj/QHT907kIearKzrrHLCeS39/9fN3AgDVSY/AVD
6s1oCokXyYMCNdUX5TmxR3DEMiLk41/IaNQzGOUpaIiGqR0Dgd/RYK38BWPV8XOib2WP0hmavEUF
4ALM5375AOojoAVFoYxurlMhAbt7t3o05BK08a/SYRl4XG9VAw7wSwygZMNvOkTbNW8BkZElWjyX
/RUfUrPRwoPQVy65GoixOtMdL4lnf7DmS/hkDSu8RsuNogp+w48r3p5zOCK+TydFmij9jYoiiOSI
Z3M2rgSHbNJymwnverNe9SEKP70xmrTrMuBNiarO/edwh+Uod94vEhlclkFLbQLPUVo+coLRWvPe
Y4prau2lGn3we8cglxplKydv+HtDwFJhxuFbuDN1EBXY9QDqHEw7Uw0wzNKc9gyvIM4ZG0bcs0w+
fK+y4VPFLB6B7/SkFpn8BOWIwVLKR99Wv9FUWM4Mt7o8MgveHLU5920w11UZxTqpMAQq8+UY+4KZ
45KO3BkzPa3mIVc1ezFZ+ClyxkUdbvI3DOSQaJeofyET0Z1Ki93/joGRD8Lw2q3ieASA//nFVK8F
Cn8ZX9KXOaUKzIugAB6arVx4rFFN50qeYRGCRM/CG2qG6hjYVHzAv+fPaleqcEwRjzh+9uO2tSiu
2u8UEPQWPSlBKPl/3vPVfVVnCm3tBq0pUZc0JPN6AsIdLEeRZPCJCVL2eaOR5McJHaNUNZpLgk2g
R46zhHTy6C5FPqmMf4GsgHBiI+O/27QrqMcWE5SRau+T0lvrW1SHzn1moMGkHmDm4OvZxxVRY7Zj
698Q9Zv2XoI7Z+d3ez8D86cHaZlXH8wq45fVhTKekpm3V8+K/kA0Y12vunE2Pk8UX4RwWxslouBo
ZSG2ycgLkXwS7YwKgCRn5heJDYX/C43xRcIyDPHi0ZnvphbcqpRuB+v5DElCJX/hxB5xV3lHH7pZ
o8N+MUL+HYFuBk1GpO+8E1nArlGurn1kX3mAXmTWSDoFHqtbUU79yF5GF0fQ9wkUt4SgBqk1cvcm
3w32MA7lqKJCZW90JTWs+n/Mg0k5XDwbmK0YntUT3/znTWBHwGRlXq/+PXKF6vl6liAJb73fxSQa
FKkrroRCto1dE8WXrmyzY9DiancZyd8Q24HuQ39kDxEKSXwZOCtcBhh623tYTN67ZtA0tG0L1cwe
IK3qpWTI3ALe+0xEIk3E+Tsad38EHWHzLypaFLsKyjBpoUufu5K+dOHe9NquFS0Do35i+GwKMv8G
3k+1CAFLG6Gxp8WrwptG4MoiJPn6JmRpbnS1H24G7iiWd7ENeuiApfst1rMiRWVjYgYgsYVnrlZM
OCXNx/I2qv0KgIl+8BGc3iikj5/ZFiAK4PyCvnw8aO/93FEZj+OsZZHpg+zTMNoCVagm++bYcBYV
mSSqtQINJs3kgNwGfb2Au6d1VB1HDQzczFbACggFOrUuSDqnVm+fBO1DdO4giLeARnwAcWt+Ty4O
ZY0XRxWaU8DYaWoa/fnCfHEmXvawO+zvL0bVWMPn3PrRoCh1w9s9hTh/eFSoYMdJz43Phl4GIlkP
kkFOt97e3Pu41fVvVRDqgKMwWOiIIOF76PrWI36C+RD0XN9vunJrwYskI2BRE6eAKloYLnHPUVGa
rH/NrSPcj6ljXZ83YARYvYgBm85vpnlusrwGw26Muu0kRKF0C2g4UIeRKY4Cg/6x9oXePocU9ygs
q9hgv7q9ysRJ0VDoYbKiPLn8kdQKDjaDp2I8t8fI//k6WsHEIu6nVzozj1/E/7414qPxfTDAOXaZ
KYxnDAUdvMbXnqCznmJT4ev10HebM+XozbyazVJ7FOAf8TyTwdIecIY5xvUsGWyRf/bmR2S+rMoN
2WxEZYO0t1WenGCE+UG3L9LRuTDIZ/HYyL2aJY6wFP+StNVQiftXvwywK3JtiXbDIQbTjLn/2GWi
e6hMTBnsEsPvOauIHaa+9bifWS1v3218qS+t2YeuJCAWN9iRSjP5x/cWzX7WkjJLGXDXmAGMjsF2
6Jn/hV8vVQIXURmrHrfA2TNso+9JvbHjEt7eOcw2Kawd/EhMDGihmS23hedzodIxdJEVzPbdcU5j
tIHiD3xyj9hlny+Uka9z18RPgLpTNwWBa9uBqrSvEaBKxaUOyAVkf0QPO48mWnAc8cPUmF+EyPun
UZlh/7aNv3ATieCPivjvwyudsbGP6T7V2lVDO5aNMxmhngZrP/8J1KufNoaBQeVMe8huiR60Jgh0
/J26nxCIoehBdUVRuR+56bUU2/J5mGXBzvusoYez73oxm8ZcI6JLjGjHfwNg81k6XnCiiM3/HbWo
/M0YFxb5mTIR2nlA7xQXaLwSkwGr3ccUm5XSSUFo25T4dMOoIHkGafCbkSRKYbzF9wPg8s8GPzHq
YhMWJ841lREHT1CayWgQcqVzT0YcDn4lwNmNk7FRd8/XhQFW5ISqY7JauBqC938sRUH54CaZZ/Dr
CRZeM/tHgNVWh+thIE2P+6l+sqklVQvDsz5A4HOKU3WAC9sxK1w9DV3JHaVS7E5qH6oryVb1zOWN
3lbf87/XQ1K0yhbEM3VLe9JWGJzlWAxg2bTNWFT7eMgCfuIq0okxo1vMyJHbCLBQYiun+5R+LsBL
S7OV7mCbmXuUwpZnq6L3qwXO6wp+l1GeHpH2zzWqsXBdL7NW9XoPIhnguyWxj8UjemDYJ6Bfs5+h
CwPw4HMSzrRkHgavz7b+0RIFS5QTDOyX0iS9PhOFBAWXSQnk7jrjSnV+3jTiFNg7LCWHVxnDpsqo
Tbm3l8OXtwBYH2pV0oUKyue7ZsE+pHbPVbJ4MjdGbr5zqfBV0OUb6+Q4ouUt3okVvaglDXpJU5O5
C2LYmbxzEb5smBf6ime1l0lGU0G83Hr6bUGgYo7hD0X+puUzn9CHHLxLZetWBTvDyBYbm2ls2cqH
olUdSRLTb8wzbQUkgjltbU3+LgJIn2sjp5PrJy2LUzNMfpxlM4eVk2AJph8uoj0ISe3zBWEUnGrZ
GU29xplQwGu0QJIG3NJCJtDkhNQ5emkNjM54t66cTle5OwAAFK8IPkZFyiw6Wd56wT5CQLBd7FeV
X3hupqnZPUxtcvAACiqwNPJ3tXPaTkcnd1DREt2H83JeCUme7lJAuA4Ovj7JUAHwt/RWL11I1omI
I4nGT1C4Fl14yqbKBENsPMue0LJ7KpJWvaVllFxICA4md5KvjtK2CsKbQyieLzAXchtPPxj5PqMP
EOb51Wrr9wphTeXn2KbMpUaKNTgcAXH3TUwNpf0O7WJRtet4WrWp9gzbW0vEjqLkQMiDW53vQkvm
NVJz9XmWizqk8kpv+s6PKcwthY0JOzQOUcIAoQajs3DPYjdmDirKKSWJ8vur0FDMFHXpd/Y/8w05
Z8aGF6c6LenqLii1sSmGRZIKAVHPGxm/dB+rRrZrqjIKv2pqpYOt9/LDJNvojueesltwz1I4tM9R
cqpJGsUkUUH4kDxCcDF8lDmVddiBhsA9ypjL/+DkWcETIx+1GIa3wQKUExF+pDetZceKKZhFE+VV
diS2LvGax0OvxtQLj/4hSBMc7IKrF1TVGmRXmwcXRIh3mnIAJTinhqssZXtrnZASA0/RaihNb54C
3wo7HFr+14RFJcBIdWju9uVPhWD78fnCodnmwg+1XbRFknfxT/vhR9G3EHW4sGTVOKsDVJmPXT85
kyQVMQ7WdI0TNc5c/Yk1NMdXXu2dh0hhAZjx7HmcI7APqIO/LJqAL+W4Uq+H0lrMEsCWnXi1uXcr
V2TqMy4ld83xq+XoaQssxt2h3T3bKDhK3F9HixYnayAbjitzo4yepu6RGAFYJUBHYFOESO/+6HkZ
S668G9ZFtnExurWwRNlfq6brkb90tsLElwDD6L7WkB1ItarVjGuXE8yJMqpxGrxg6jsx87KTg1jy
PB39AYUw7blKniYM8I2bmHZfSHxm3Tfl7eCxiAVxuNdWTY+95NDzMLZVZRVR/RNlxebCRtmuUX2Q
THIUxfuu8nXfds3xwAaX30dVWSJ+TBwzM6FIJAqDUNdlxY7pPkAPGxx/nH0zsjNTTymNoDuP+CFt
c/IEQgy6rU+LfJ6mg/5p3d8aNTywOBzswoHFrg/Fw3yrrBQHtJyYn1upZFIYXNaQhhkfsctLFAR0
jGdP/6d02WYkYKgtY8VetDwc5j3Awf1yIC6trnmpqa7TxU4jVmZniNEsvb7BCT6NpW6+D1+FurVX
lbuChNsu9C5WByeEaFES44a0u/FE5mfeAwPuIZIyrCBcU+7Xa0+TP/nKFso7kAJTSIe6XwCb3IiQ
Afyv6AQtuWs9yp2NIF/Pdt2guHbrgXn2GIpX+lqEAdkdpev73FYjWkxrkb0kxvi38bVNJ6Pwv3Ut
7W4ezR0w+acEq7v8y31d3H9vqKrZ9ThEP77h34kuVV9M4atWrF/wrTFwVvGjwb4puS1gqT7PwZKv
bIAkTSO8AF0nyH9dTqTrRi8H6LivjQcWUcjcD3Go0wzNdOwMW1uCS0LEiu2H2PM6rLD4aBqNPUch
rHf412LTgrQ7Trnap3hg9IiVhYX79J/HkxKqizKkJ61M8LA1g8fSZwOPRxivTzpnN7zYFZP9EzMH
BvS3Sdx0SM56hN2V2g8PLyDYdVAdV47HJweG5K1iRPxmSwWSAfHiFPU9BJHBHnnRln2xq4P5RZWP
3lxk8RDLcH1QF9x3an7O82BEEqGZ0SX+ttBqtY2Voj1kyWETvd9DXCHZRW+9swvCW6LXov/4CHo/
g1vOSnSbMM1Q3zevwSO+MHU/QqkMSrVgTze2imR7Oh8XEn18zuolRFCJ+xrps0d6ddbFkd+gJ5Ct
ZjAjxxV+1wBDFgWD7edjy48KBbrh+/4aGyfrwFtkxg+vNsRlGy6csrw1Gnq80TqMEVxOKFI4RYOh
IlSUxpiurwuK1ZJ8j1j3mkBgzxJPtBv1kgshcrpfjnUQabpUmzDuoYuvAE/axxl8OOIX2IrbgdA4
h7xX5vAnmDwtrSMUtLt5kNoEmUo8ewFM6yvqtL+NEnAVFr4Fiv3kEMSiRiPjt5X9dWcj0FpQijsc
YZbzSa2Icnc11NRRuxQk3b4zSyDUBtArpwObJfZ85OtXHPLDaz/JBSvhmvFY4XWfS4oXN/bHigeK
YRPVDghQCia/Ob3Fg40lx35a5J6Jm2PB3lbzHRbR31MshiWz8SImn4gnso0Yaqlwtdk5LtmWuCKv
PvgCDUfd62Fg0RcrFEWjdrxQDpTuqeHYvpKp3m5USq6aFdnfRKqsZ/EAOittouRF0yxEpcGcJL6c
LmAXONktyRqzwoPdidFzxXGRVKkEzgQVc9J/2piiRL0/Vg2DJyLg8EcgYMito+55NKDCN1yorcbo
xrZtAkmoc4Q4uyqWDhto8uPhNwPXShbzfsCd1GGArPqrErj+lPlJfCaad4Bp/6hz6Dj/VoUa6ACr
z2uW9TFkhuVcF9eYrrVB4Z6AB/SKY0N/M+jJhTI3cdJ6K/MI6ULGpdIn8zl66Zn/HRbLqvrO6Zeu
ExRAuJvy0xkT4RwWsL2yGlEzrbmnk741KQqonm6qwU/kMhuFkfRCo57nZkYZNRi0IIKPtMzR7XG4
HGTgCrSIMx23J+QzY6yVfL7LCc4H1xNh4VT/iO1HOh6vFTdWfLBQF/WstoZj4ow5Nnp7t0ntNkZd
jvnyQ90e6cCxzEf7moUQkO8p0ERdaSP4obh7pfCIAOqNXFebOENXOVgHcA1o4Y62hOEyg4XPDfsF
AGAxb6QkFvOqNl5QiMVQo+6LrwmqzHAc/g8NmZpwr5hU8eu66ChluScQkgmxUumKc0ic4a0heUm4
rLmCEVRmnRr/748YCS/xZPShM78nNO8LukzLE7iVhWSVp18L/O3s8tKKTL//KpAN3L44gYxjmrPO
aTyyNPkvHLJOKMRPqM4dLJV4ZcAaLkT5uCRy7myyBrS0DAnQRTqrhEZWBvllz3w5h+NP+XkskQs3
nBY0eBPCYP7UAZLbP6BDURPfLl/Hb5SYI2j3RDDOTROOx7qBVrSKb1lZG3FnKsLt8OJVTu4JYz1D
z3SUwD2VFYpJGzVSVVNO+eqwBMyVP3XU6rVuLCRueEgV6Dck9T3knFMpFIzu5YqaLmmcuqP4+DxE
pSQKxJ19haCYtmZGU8q6ASISlyQ+nnLUjFuCas62hZNGsV/Vrh2HZzNDfwx/CIxntsX5cbae7z2+
f3e7XWaMCj3bMVKczMLtdGJk47Lok9TpQiKiEI/ER/shkg4/txfhpDneaqqjmTqMv7kQPw2IFxBW
t9L3P7zoGNreE8nYejEZBMuldOKl+BYZv2sbwc6vKxu7esaC7K8sEkHDyE/zSd032AivuOfHIIJ5
ncQZg/W/uIRO5bx+c4fxQCOMwqknpe2P/cGyFYOD+uOpN7AEcLAVelLbT8ND9wpky9SbTTx04M9I
4gQ14FW3djesWCL5GAWeh5CWYtMJ3v/ir3ob1fUXLiGLUWdnDnkcW5Dei+TzE1zvqQBDDG62T9p9
yJh9gTbL6b17uIiQVcFrbR1Q0XJyqQZxRW7MZIEpU5LMxMt/5lbBcywDYIs0KcNxETMI28/xC6Fz
4TGnoNF9YolbnO9H0lNdBWEyDqyABR0geWG++mJzGNF+tso+22z1oVn7lU7r1FC6sm2CM0JX6+L4
IqmmBEHlE18kD32TsIbp5Kr+p3hvYNfQesUTpsF0Fmce03X7LteCgm5RK6Z6uRt//a8zm20lXu19
N/qAcrzmLz8t7nW2WrkVwztzdZ8bMcE5Ars9oFxLDq/8DZ2Ga7vAJwfVZr8lFBEWgOMvDJemh38L
rdm6hKHSvb228PawqQ2L0z1djLmmc4TFLuEOY4DxbcP3bNvtvS2YDlb8w6PsC9rDYbVFG4swnvPU
Qc/s0ii2LsorOYMl4oxBq0NU7+EDvti3o/1qUlhIX/NzLaFq/1QSSRoM8PwBlrIjFLYLYDsp45lM
8GY1Nb1CIe9HxzGGS5rhJ2CLQ8/7fic1yXkyMH/dtAaeJDSQx/lMnbJGSU3+y+3qFjLZ+NmvCsUY
OPZdxkc7za6r3O8ifDg0LvR8/xeL2hfs8QtLj8tDEeK0O5jCR4TJ0CUiqbI8ZgTOcFkHmI9nqFUN
1mIhXEKlDsSteWWQmZh/ku2jmhh8dy42pVlSxuijv9jZ6GwXVVTRdob25B44kUnQE1ti1cjDSofm
J/iB6LQQvaG5HyhLB1xKcMiRRmybD6LuvPGIav+8deGWg/L29oFdmxkcXlYM4BeFYypebr/JM2ZZ
MYFeYe+Y7J7BgINnqy3z/ysRmIBhxnpVasxxc23YL0D5HY2Y9AenE9sL9vrPaCx6/pL1rVHSrqlN
uWEj/Zx+J4xqD4arnc2ESlhXSXF2lnpiZzPyJTsMhEj9tzdum+fO/e8Yt0SI3bYjinn3d6i0FB4S
VY+BdaUrbxisrTd4RPDBAlZXN+E89/URb5jG0EDhNUEF5QspsAFFpv8hcZ1pqAlih0GUHFBA6Cjf
UpsJpz+kpNvtY6deDxP3op8Avlp6y9xZ3r7cRKXiFw9sEeUA9NhBvRCWm3tmTxBpBlHq76Morsva
yOf3E9tTuNRrhUZdFLrRBPNZh4hgknoN/pw+i45RVdpNt7PV2MEVY6Rkei4rWs9KPy08+Yzt2iOW
J2CLcX+yN4vqJHzf66HxYm6AFZGmpmelPWndURFPooQP3O7kCiIg7yIadWV/dQhfOQqCWIwIPlNN
U3hbDNYqUpVKVzntCqkiIGjlyTQOEiSob7jEEONECUo25rMOJclxkDAsaS5EKTpXd/rHoP9Q/SYv
lHG9J+A9BRA2MxlCr9yd/9yBgq+IFo7g6to6jFgG8nDGzRmf0QXgUHkDwTbKe9fNfKYoPqtrnmN9
BEDuw09cVF19SWY+Hvh2lQ22nEGhcOzP/hrs+Wo4G6UaFqLKiT6NVdB210w2c4NnM4Lkn+y8IKLX
JarmiQ5/j8tbUezLjRnT7nK59wc30STvo5Kk7xnt7Sr1903fNdjoxb0e/8WaR3vSfRwu2M2KHTJz
rp7bZ6jb7ovExhVw2LTvYcIdLbEvlvUolmkD/9ofQTjvqm8Molk4iIZm/J6zdoeDHdn4Zv0AJGVH
fOcFiWAzefuEkzSb+ODDLR9ni5WwlsoJcHRnw0mlwoxwn11zu/C5WuYTLL8t3ItnOoKRxIEccTJA
Y3RCs+g240ZsxDAIpm0xC47HDyUcjrC8Dj9aovAB8WCn9kyUA06flY4UwSeAO7N8s4ZKkJ9NyBs4
2rYQImP6Josy7IYG7jdj9w/UAnYli1vCw2zIuumB7R+eYCF/271D9UxAPOWhE//JhI5afxv/joS/
KPTwhSZyGxN1hE25CI7QU6gaomMrFPfGUVbmyqhKsNsAUhba4I+yON1bowdqdtos6yF8933ZXhDf
H0zM3Z2zn03stKRCfXHCYTuMv2kruQ036LJiwvLwunO4qJGmfEQOrehwnGEN1wptmAAoPQK2FGpr
E2xqYnTiHB1eE4Fp8zFy05q4uS/pfgoYq8xpjD8/Il5fPBy6xCPcaj0jOykGVTJBzLbO3kRFnXu5
Nmr8uzLRvyOUtQUbAE1mBZuF9yZuY4pYMKbk7VzP9JHAiakdWsAoPE24pDCE65o6/vXPqPHEV3l9
CS4gyL9t83POhB7zLjmpOaYeNumu8JAy9CHdX8LNpK8qA0LEm6IHsTMO53CDt1BeRigSbHKblmGP
iPsKWbdVdd7/kSG3C8WU8NdIIv/+ILDhhjbl5MyqoEOEkNQRcgf0MH7LQeoit9Sn+iOujOSiEPg+
SXNb511f/PNSl7RS2jkYVWmEE5UdrmWsik6VeP5rORZxSnlDcZWxn/fH5UEFr3HpjcqUMml9tFLw
rSI56bkOTD0T8+d4XeHwsK4oIWL+1UORwg7yg5elLJoulFe8ib9N9bPF64km8D7U6en8UY6nSNcx
JKVexUajuHhFS4YZAQjU6DmsG+x6a4q4hTEyj5gr0MSx9UNetgqEacC3mXbpH0MTF6jPbTbjHJze
sbhMUGGgUBoFL3eOqb8uzUk+RNn7neUlEteGgWNrZAUUir53Jfpg61F9+66zcSC5DW9dLEd3N3wL
pL7RP8Ckbf7NCgwK/58dxorT78PJ/obNy0RJra4jJcHVPYbSTV7hn4Gx4WqCDmDtvIqLVrAa7qJR
T6nkZO/YKPse42wRgw6dzCn3lxldXwBJ81T+ZHPMpjiMG9OyZNvnA/S7+59mwpl8LobJM4+7fjQI
AUl3lBASFbKjMB8WdUCyCLaH83mdfIPdSbB3HUih7JnXbZerIhPtZbxlZneHrF7vAgC4UUHmjvye
IgF+7eKcXclTyyvko/GsSaLvqjufW0/C2rM+cN+QgxCnuU5nlCK6+IFn1J/7kHNA0nJVVEM7xj18
/ciakq3ejqiG93rUxai34J19kF/mG7WPPikiaVHKJZJO1/W4BPo+2IjSl7sRjJQpgPF3qPOD01Fx
qcZGCRW+W/nfw7cUIs629weVLcRMWC2R8RSu0pd9CjpXRMd/k3wwM2yn2yBIUaLmAwnP0VS1nVul
F2H5Qd7pNj8SjIFiZ8/tnwihIgFWBPighn81SbIgs2ltlgc4hJSDN8h2lbVIV1cDM15jO7ubbZ0j
F4Uxf/JzbbPOmGsiUSRTGK9V9udWdYRk7Md5lT9GEwIRX8lVoWld9aOsK4+0hk86NKrLyGPYCQKl
5F2C64PEsZuX71xxa2sTQ3j1tzN9edznieH32KGBEEXeweS6/B9NI9iGFGSmYlO9H/SoKrTX+orY
JYGpK46Hz+B1aEIBynSiE6C8hhPUsOgLhFrYtGyX1N7Zldw38qdSkRW3pwOxeoWjswLZFm6etD9z
pS2QXNoJi0HPK/1bbaQPOxGxYin71CKOew4m65Xfjy8irGhSFARHcfANKR74px03SymHDJHIs4bg
RESsL2fK7qjZeSIdqHZRTNKCAC+mhv8l4OEpvr1TFLyaiNzYCodJsnXyAPHu1TY7GTZRQLWx3jpk
ompH8mw++TDhPF+eKtxyoVU2u9KuB+ZwDTTCOeBL/5ksv1sIoBZTytH/LxbrWFSNjRO17nN5+CbB
0GmQ7L2HhZnrx58nrKPDDQ3Jjp1J1taiRry44vxROIq85FycKKzvdwmL1GbBNea5QDm+Nc9DrWkb
I8xDF+VDr8CZW707wB+nKgJHeMho9VoymOIlWAYq0iIr067xOJLLVNLiD6Td7jUrLMZQ7B3xfJkA
7s9XLYSmaGR7HZvPQGEAMA5BXBFf/UHfymjdaF6bHIPWD+E/fbUwjOA8+1VJBVLbkfUlP55Tt02J
CEN0f7wtK6n2W390JHF0wBF00ielRTj49bBhp9RJMxvguj5oHiG4ceJoQGzpqJUGdRYcPJ0s+L92
XdBBPyYELE+4aRk9L02LP6+eRrXeRRYQ0UdoNnUg6M0+kgdSwPyjKQkedZRMsnS6+G2fYecKaVNP
KAnquoAgjeghnpkVr0kKOPiHh/Oc2UFS2gEDG+pKhIq1a0mx82SNyCACSZtL8cn0cRomIYQ5cNlH
3aIp7juE0YyM+40Z8/ARKDJFLXzfXk+jO21we6WukzwMmI2Od7xrS7Rk9KcKuakbLzEWiUfLsb7f
75yVQ27K0mWICWfq/E5PxVyAaLSJN+9c+DPcAA6WKptEo3KzySdyChvhKyV1PkjCn3Lo4LVbMMiZ
EbechNpw6EKsyCGCCkHIwSwTf1VC9HbbDzehClT8+2lWqoelJCvac5wbZafCsC9QFYsRzzQAsk4i
psVk06B2dnSD9s4UE3E685xFWRxgAcaflvlRdcLqH6iJegQqXPoZZCEQ3fXG9O1zBjhjiDDUfDhy
ra8l8kzv4fgPfu2TENNbbOQxH1Ws7HM8p5A7GgEtgbs94g9ztb0Z1jA6qJ0Pq9UquzHI2IWVunAg
p505Mly0xx6DkY2/6G97FIU/ysRM2C/bedxQKQyakpUWG0RBJ3cV3sLarKHqZcxsWk+/sq+kqsdR
9qtBO/czAbdcNymWcpN+bbEZi1poDxjPeenaehAiHFI/HItsSOfNgpgrlJ+M/9F/DIaF0loWYURw
ETKnP/IrrZ3aPf0n05ua64u285p+eSC0CfoRIb8smEuvWsv8kPFw99iugzxKJ8w5y8cieUlO4W93
x48iA8kGmRImapoAcLoR/ZRkBQC4JCo8ufaz0UOozFP2IMJADkyWD2vK7rFZ0c5tF7h1NM8iEZup
CxoMRByhmnUrPz6WS2Qcv1KjrLRWlytLadtivBYUkc37jO6ADi37Q/LR6Mh4QTQUFmQZejXPk6Kk
k1TwrYyL4k0LjpgQgRY0QiQAlooyBeJtL/J1aiFviBB3hYO97MSUtBGzyWm8kx3Y9GFKa/N0Qzey
T2uEl6gjTvJiJFLYYq2bX81ar8xqcfZk9k0bcjTk8SzK1XDV1N5kuS9oPEZU27e9Em49bfTeg+5L
+JTvOhmiCDavBZyT3L64BsvylL0/3OMorvnzSBMi8eJgiujOoMSQuiwfYG4QVszS2BP5odllezGO
FvZphSMO2t7POd85j9KDcnWEQO909zRN7T4iyTMRmB+CmoJ9TvQ/uGIqZBytaBeszl+P1CN5kb96
gFLBNHBN+Dpf/leF7wK4oPGu6JnfNvkKrxIscEQJqkdpxisLLkcU0JPtm2uNP0usaIW3lWHwrNzw
2CwMsQMg5h1Dz2angDc3Ou/kAHLBKA3BhkL7qWNNcBl2G6aqAFiypVTrwo+Y3KzLUqpjGKZvhAIm
DC1EKpQ1mmr1KYaWzlQ7ukh6LzXXVyyrL9aJjLmmIcraIJrRbWfvWO4Dgb68gXsxSCSjVntCIkBd
oOwBI8Qkdwb6HYjPOcPc4iivd2Iv1wQBT+qclue4cmOaZncRNqj6KRdjExU+v/Br/BHS9zakfgZH
qzCqs75U4TH1pd/+FRW8Lc5W1UzOSkgBGY31l4YNACyPT6ybAy4u7mrtZFI/GSYP51JO8J03k0em
yxNJXY2kpA7hm1Hk8uJ0+q8EPQLuEjwW0CBWtUPEAHplMMpBx4xs0NeYUnwHnHAGdJtD05hYcIYn
f4Tv59Iao8uXJdfbsJWzrvmtdszwnB8Lm/yICDBqub6mmopxaDHpGddlgxrhNZgd1e3Od9JFzBWR
9rQj8vYQVDSkvw6tI4PjNNkiyO7CTNgn9ZXNcBNewn8LY//eraKkPY5jD1ef8RLQLs1iHeXadw5C
kZzpze9gPRZTxFsvJTHIKw6Xh0ex92T60QL41IZw6clYVz+cXrvxYgjXz/K/ywfqp4lGWmh7/vfS
vEQYV1dhtaIn8RY76dOPQnY6628wR8mFn0PRvGSg5aGjNEXPxl9DsFiQ3NHOOTTp0u5yJZ7Y0d39
UBAQaxGLWBS0VyWVUrnHhl/otdCnOAMYKnfEaZYdIUkXvZ8QtT3hhbI3gYLaCW6p8mrW0H6XcAQx
a4HWXbKA9Pmxq4YT/X42p9Is1bdepWEo/NrHlMdGemzPpWuAG+F2H3fVsxwXSX/7g/dFzPXbL0Z8
vBPItAa9U0/ytfDrWpc2uo2nmkHJmP55rXa/krA07UfYmWVBlIwt369g0SRUDlJcu55CMhpbfikW
OIyeAYLqKkZ9qoAXVYO8uWdW8XTPN5MYK3NeGPV2jcpNS3nbCwWES6CwE00fLF8zxETpkrOhRpjC
xGrWpuLFJTq8bCKone4uBSrUrXm6dAVL1I9hxHzafj9jjJh4ojzKsUIXqOypeqwb6LDMGIA17/47
ZV9G+Xrd33bZvn7jB3x0D5FELPz0FHUjEpIx+ntwdzSB9JMNZa5h2l9Lnui5zcuw4VhrfistHWxF
9acURjwaMKbwhv1b8LSiQXzUrsbqkmv4ZFsUYLSJqHtzUO+voPYwqDQi26Haz5iyqeGCRN6O+58x
61HQJVPLmQpirNsX2MrDLso61o1nyDdgo0gBO7OK2nyqw1ePTmQ8MYR5HENaaxhSgALRoN1dofx/
M2N0kashajR3lnPucDH7UCupuBlogYwBuZ2lcIhAEf/18KS+YPKjLGhi5cdwdoLk5A+P4mPYkiiB
fdvAJINBMqkfmdjx1B1JCEB4HB0AnGVMvw8VNXGbDUQ2vMAF6JaUGrYkLS+6PH+KWpsoBlLlc4wi
C/TBsQY4YnW+NzvRlUIUB4Nm28RVDktHCx8Og+pu8Man7GZzVnizahmzvbbxvokUiJQ6o4+r2iwQ
q6tLtd1GBcJLHOIJYo1s0gTbO+cuVWLYHdC5zq/uI5jftGR5ucovbPTAdpQ2ltZr9VBCgQ0b863y
9GAIQ1xBaGOk/RiMyWI8CD9oDo1pOd+HRVa8BP61g97tu+fZqFyIVuPagFKHYjRRPd/m6d9WdUcj
eBsTJ9crVEInuIdjFPQ9DvRLSRx8fhH1xybKwWjT/qAdHnTiZ1/VnxClJkbF/IBuIKYyHjqq8THH
HulDNYwfVnVo0Vt5Jvl3VVnTdQq1lhGxtmtY40AdSzcBgEr7fPPV/9cGWJu0sPZKHsS14aPhQOMo
WXNx6ThTScSyfGY0aVtBXooeMKEhE+L6x5/63fSEoFhC7vSb7DRvxTg2i1171CNF9xYoebN29nMl
/GqzDu8HWa7zbQrRaLBUuKgGqOMiYIjPjQdK5Y0A+6tw9uDijdp/uhqQoEtD5pZc+QLztEqn40p2
Ps1dasg8OnHeCI48xES22W4aw3h5kU5eCKiUDhEY+f52C2cHN5MYcsX11kidy5TDFPglv8igaRQQ
9Xt9dBnLlMOhNXt0HTWUSeAiTGgCuAsQvemQJa4eTMJvOb+URcsKQ1JW0I0eKczPjHhomI4xNBZR
5OVJh/SZctPLutZ7dEaQ/Se5k5eFvWOHeA7w4eNgSgM+AviLiDSywZLaK6y0uG8M09XRlx1oPbKx
NX8N6UH6H9srU5bZCd4rh0n3dJkYVno5J8a6yWSrzucELFJrhES4/rjO9usv51qKwdZmscFrHkRg
DvBVZq4FQ0wGQImM02naWTEAYkfZ8p2+tkOxzoO2/270rMrCwmBfeVHpYs6EA/2synoIMVi//w7S
tcKw7upZDzRoHXpsoBvqu8mipcUUL4e9T2XrQS31vrtn3uGGvg+1g8Cb6Dz8wRIngTaprJAPZHBZ
GZps3jI3z6BY0gL9I8lAE6MfDigIlp7nfB+RWEFiYhRy38JVhJ1vNCPKeAgAE2LU1xuhODJLNLOD
7xyxYLQY+FTfTNuyxrWi9fzgB8X/OzxkOW665WjDYyJ7sH05sZLrwRm5Pulza+WbvG6qpAcBht+0
pLf8d4ZgwlzWiLGcxoFpSCax/8IjI5HQFYROwuzT1gLYgTd+ZnbytLvRbAlTcF93sj5cHExmfoWt
i9/xEXYv4BtlRO+Goaqepa9MUu9Y64f9wappqUwMlpNC/TCza+3G8+EqnF+oJKW/8mtnb2tJIFB7
g7nWlIxUHrbnCQ6I4QJ9ibKkkQdr8pwDXmgD9SJidnqwVP7ncCHm74X+dHj/dSmTZUSLsE4Le1iS
uoPoQNhJE9ekA2RJjgYKI9Y/vsr1rfLy6BPaubGXX0poxq5UQ7hHzhwwghBN25MjqbZeBydixkPd
36JZTpljbTnv0K+xPqceBcQBvVF7miKQIDpTR3uD41fffIY3oEy6eZqGoRBPOkgz4Ci1/CWmwOwg
9DSDcW8ZGkTV8zV4p2BrF3Bi9j5NTuUVLbPY3kdfjvrijQWokNfq6ZplPjMfhmJq+zc9MLouTEDD
AQNqYeP2U+v9Ye2KUrJd4djc0c/8N5NUCtfuvEr/BHZrsoXHbIm2S7xXed+IN/LU562pb5YAERRI
JKztk2uHX3bUsbvG0DsLeC2YkTaa7eJD0cgqF0yayp+OsQnraS1AVbmX1Fqs7rv0cLw+DIeNU37N
Rwo72TzSQo2tqoVHr6Kp0RifjbqHDV0r2YaWboh9Qyi+IhyLfIKOr0Ns7Ss2dcRDUx5zGG90KE9N
DWwXzcO9bC9ECYpcRGXWL+pzA9A8+KyYwv3qDWYWqmJ/b5gxJmzpM8qSkaKIB5ZMhnfXUkYLWdG4
Z5DnPvrP2/nLIdjkMu2ZqdHtE3xXgdHRTls0HVWVH0R+3Jw7EAarsJvO9PIRq9lI9Er1jVPUknes
AuKdc3LGd3RSJvRgaRjbwgWj9KXhM4ztKcS2PkbbYMScWGmCrL+FNsWG8rD+fngQjIlkTAsv9Uih
0v4gw9EE9l54iMNGkz9g68fiibGL0+zMeZaCkcktDOSN5tCMSmSDTPkzN7AV8xGHEoToG5zH5FAU
F0fOxzSb/XIAD+rc9cdvKsL9q+KbguitFZ18bXPlJN3LpzJj/4nOpemvSkvAEm1KB31z48YKZkrc
Y0wGWG24qWWq382srjf3vMgXrXw48qncYTz3+j2WWbIYUIT3f6qJ9fSzHKuD+VTNmpzZkM4742b0
6jMTMzmg+IliUNXwy+i6B4B7EgsdeS/icx+oHcylDsh1xBIyyDn4qatjz6KAwr+nFLfjiOLM3A63
ev3dYXwEkCe3zpO1WnWkPN7q0Erzrwr9aEnDQvPjlCAzYKLUHjtrP4B+EM4xE0ZcRSof8WNiS66H
Iud4OLCjY2rDfgfG9Zkh8/KyAAajNRVTKTiQtlLANwTcq/J/bIyHqMePHRT0iIsTipVGOp3W5Vlb
xC/JVTOgE//N1IiGS3tUgIfupuioEnMua+s3eoN8eWftXLST8nMMup+RzB4WHuNPcQAipkkN8TX7
WTAYcF+SCHoWFLk6nYwo9o6UBTB32b7qbNCR+8xlCC55shXQ/mWDD3dChdRJ0ElJdn8FXwRvykHl
WXeEONxyWhZplBaiTdaH+hPLcWHgDMmR9z4BS+NgPsOGvSb43MZId0JsjHFhP0bWHzAFGi99o2dY
ZB9Vcr10pwR1guLcZxUMbx9M0B+Cjmgd8V/SoYqbpt18E3JHnSdkgCmcq2nkSLpgLxW49NKBlXki
MvFka1DaQhjJl7JoQWbbrsIGfyEweOJWQg4PxdPXkBeC1ST0vyUd3DPha6Tzdx/F2RbmmOsNdnyG
z0cS/evVZqzCl7oBKZeC7sAajDVMj2S0QnyPBvbSoH4qPDpM79OZ667waicaFDVMa0Pjw4bk5erU
BYt4OW8Uk7Z6mwNxBZOLAtWX6M4kk1X7znZEjAhCID+Esf2NiJwbj5jL6EgCHA+G3i2mkzxc2F25
74seXb+6xvuTKu/sHhBhJtIFis62bprXv2VJouc5q6/EauSFCHHZtJQzLZa6VuGcvSuiM9moQ4+w
1t966odzbC+tA1oSaf8i3h3v4e3ENLKEjZDAC7bXyITqc71uJWJnxvmUlTjM14LURaQBIAmjaxKV
pnOB8+zk4gBZP+3rY7k3ddNWC11EjlOVBOqssIX6jr3OiA58hntDLnJro/JLfRlSoCNJzQlbXRz3
Sli3VNj8JomxZsnGV6gOytO+xdn9xAba/s3hJwFW53zlaB/UUm0vMNds9H1aqgJM6HWWXbC02XVY
H++q0hP+leydqmoPGv/K89+VmZUPfk7gaRY+QKQT4k2DtJgohXSfwCt4kSCQ0vKao3zzLUey/emz
o3E/uP85n0NMLPlSYUg//yf1mE0IsnTLBB98p0f7VEYFEAbZxpClYkwcmOCxIAEyPyOy7oAhmgK9
gsOY6RHP8m0Me9sTqCmIC4O9vVvXJFOFLwA/Vk9/0VJvLAGK+OItC66Iij37+ESxHyk5AadVRNF+
C/M9EHRgFVMAL7Mfxu4A5kBDDhD76dH5FjNQoMA0naAhvh3QfNlaCJBXOTFkHhTNft78leeAqsHj
Gq7vmWz8JXm0tiHHt9AqZysk6q/cc93QIMaWvLyF5ZAdQlZr2aqJ7rrIXXUr0gJiIeNZ4lxYrnj8
NKt4c1S1rwOLUgJrw6jLkvyj7WvWcqpa7vPPAoppCWvrbVEjVfQPo3upLn0lQQqpZrSJ0YEJ4zH6
VNl7RHF3j+yyVwRM54iW6savonoXddcys8rWATa9ZFaKKgcI6vn3W7jgZsk3A7Z05R4nid2mj9RF
GV0jH9IKQzcchkQmxlKlxwbLUQchlr0j0ETN7pmM61YGSDrIoHQvNzJKGf8QiN8UnungSfO7lVNL
UWMAW3DSS9fAv2JiMtWhe0gsvD5xZS0dn4KfE0z4uXjQE4p8Ed8vVFGM45D0NiiFKQRT0WzvGQSS
Q/vVEteCJL42Ycc2WgU6c1l2TQgVHRhH+Kl6NNgWXBpl04zLYGpNadthjImPD0kh6YldVjpxxRRu
RYPpsnVY+ipLPqyD652B8jGBt+7DqGg/M0ibzycL14Zr9SHn2pC1S+9/PkNyS8A2aIzm04LG3tEv
5DryOk60EM9AZODzPzcgrATfQimLhc/tX4JPRR8ryPDx2TI9v39HOVYhtAlFq8c2D8CTfTJqU5Ps
32/iNSjI9sR0S+xh9uhZuqoRqo+PvO6lMIA1gbplgbiWRXky0NwUBbZQKWTM83moRY4Xv1tGxbiZ
c6f+zimrPPyXFkQ83ouVUO4hQOLnMxWXpAjF/xyjHu1PmQQCzpaXGSaFzqjbXZcyhLx6jB14BNZU
C3+5dl6/Hm4y5OpSyre1mXWl4ZcwfUBko3LN65LM6KRcgIFe0naxmps4DbCUlcw3HlcjZGj6isUJ
KxdRAJloDR35BT6TN/NBXRDfvi0LiJ1bsbE2hIEUa7R0Lta3hyEKmKz971gdYdpGkJMYYQ/U+qLg
tki/50IKjgCFGS1ME/hRkNw3K0WrguCUohDoTQ8aEv98KNzH1LC45K7MHWmJtJkLVu7btRXA7dea
VKRnqf3qsjAkkbTyw4zvkqc56YmSv4XmTOBxVxBnkYWv6QFKczsm8CDFPs+YJVpLAC16PlXU88CY
PJR530CrdK8/H+gcfM/CD7LpHu6OrrjjqPktNEWtPUktM9PzxaERDvJeSdC1mSt7pDI03dcUOKMj
IOoMngfL/XTlftaLXqpsCWffY5nIhgZznDm4whiVMdOyvfE5vGI7ADdlkkK0INKXE6DlS0NjXONk
fKe38B9FTfSoHYGnfv8GBrOJVoV7oojLqDr7LUGKGvxmMXRT0mPlHHUr6RPwcG4QUiAoIY3vMK+w
15mZU+4I+xp2aJTd4Mror+rZg82AsNrkyoty77/Wh5uEgRiLYZaiQBN7XSOzabSgF9h5C+zs08Ax
13wNM5hvS5bOnGaQibSoCXWtO/izEGHTuPAlL6/0UcP+YcoZhM6kGHN3vf5d3XWyND6TGG/Llb+K
a2S1peAk6+HN40D22uMR4leozrMnk66BkY//932/2C1XuJ/6tvlnCEnWd+ZQe7g6788TJKARoo9f
QpSHFM6AD2fgo3hITEpzq4JAF0F/5j6zoJHYw8d7PinDmiASiR7KEDikVes1aH5YxY65cdUOg50X
r+9o+B9/7PHvPHz6I+HGu5xfZahzl9MaMmzb07GBX9iIUCeKJ3/gy3lVoeGJrBrDKK/u3+e/aZ6r
wjmmhLwUN9n+8rCo2VZ7XKUNLfz7mQhB/WwpyUEb+89UFbZO0Ah4Po397SmcPjCOFnaVr5JbQkEV
tqv2KpxewUIp1zOigXie90x+dNfnQ6scVNRi3eKoIkG3W4KUBjxfM8rDWsDfvsI7NXpkG+UXX3Mx
cOxAxr3ET5jwaNd4ig6YePOO7lfdn78fnhT9HWTN3zRfS+EZn80hEy0Ho9XigB1VkfOq07IqsZff
cQwAAAIf+TXT2MaApDC64lshBX1uxkdK4J68lZPxKoHB+zMcXkXQGfHwym/1tkUwgOF1ump6bC3I
bF/DM5nCT/DBsh84H9Nk3jffJMvy6gcqiGc+0V7gGjQZMswCsyc42nbWmYto/GCf0hGc1gJgbF1Q
sErYcGpTxZ4Swz+GjgM9zlnSK8TvgvP+ZhiN+NI9reK/GlttcvsGoHSruO0gM4VQauTOum+HrE90
AmK9uFBdH+SEMrrxOkrUBxOtTeF6KSHorgMUhnXGbPXRZs+gb22O0GfUUOLbSXFph+maRfmVfmJ8
lARgs3a7wZUXuLYAvAxYz1kc0AAPXHS4i49V3TdkreQmrXQT7gSEeSd83ARsc9tb3mFkYSTgFsP9
7PsSFfPOCnA43kNg7IrlU20i+qK2sC5uZ5bWDBXTDIUvEMtNLTdqA+bkHWfcXTSSG/37qCZNQIqw
3D5VQInbLTbt9QODJxktu8J0A/lQgCNWM/LYu27f+tlqWE2Es733RZJynigYmsefl9KMD58NVRQY
w96QFDf/DEfZzgKkWK3gW35uBqTYOp7iwPzynkq8horraN+nsHOfZX+l8oI5k5TvVeH1829U81Yb
cEL7PLCkZ11vqSRodf+2scIrsYn+VI37unjjIBSdXBO1zy5RgIECM7zSqQ4cCsXLQvdMBlL5VlHx
mjIkR9iAfIF1DZjn3UdT5I+QJUm7G59U8U7cgRWaMsra10kgDI9098m4UsrLOsiwglWkZeJK5GU3
A1kpnwo38n44DRXcj7khu0vqmXcupbe9gNE/vE9A1yMyfhYukVUzV1xXymBRKX6u73533pbNSwyL
y5TdX0V1yntttpDvhDGxBCUsaeboxkTY+bYQX4lwM1iayoD6paCjc5xVJbgvZGWmUuZYlLbnWoFQ
TqBMjRWxOgetWoQW1QmH1o0DnAPni2Fg8/01xRJTtlnq91qPl/93VOdVKWhjdCS1yTtoKoTxwRZf
4RUtY2sMLsoLCGciA6/UPFf39lCoqD0Afnvsi8KKC9vo7ZWCevQ8NkbMzRmPQPnsEnm0slWGe7qc
j5qZmsbTNkA3tztfunxyFSEWdwgUmxE++4fLWbBaZkeigYpv9cwDw2OyOzb8/mJ3kB8SffDaro/4
HEpvLpkHTTyLzdEWC+7dAkk/Tuo2V5af6z2dHGEOC9bE2cXBkzuiG+urBdzafS05yZd72PzgIofQ
U+9zgyySAPYeFjNDvLbtVXzPhuflBCMqpVztSBTiAxiSAoWRrqZ6p00bnhAIyK2Ay5xD+hNbWYhB
T2mqEREzJU5/6wERwdEC9vNmghfjF9YO+F60AV+5IGmWBsAI3iP2oAZId4v6l6P2QUwrXktYnnRW
dWzder6XYpk4gv2eU+VQ6dJnPk9cxhAGzvFJ7lAk9ObJ241gPDcPoulWfVqjmdx+qPpfD99JZ6xH
uBOabnYxT2XWP/jK8fnFQRe7bqOxa5vVCtRrP//vpqE9EW4t17Z0aTojTDRshv+dSnoWuB2xPxWK
0tSSGL72kCY1wkNhoJHMlpvkGNik8druilw0rMwfHuiqOqGzvKir2jZGnZBnj8+GzozoN7rVeMYl
h6iFofnzDKK9BI4hGv76MqRVB9S/Dp3m8kJN+B6TZbUiTs+cJIAKPvaGgTNcWtWLi3GU2xgLNouQ
7QfocR5ALDWxsE1cCaws2iTuFKd0/Ev45r6xH1K7T4ZfalOdEJQ1P/zI44ggHbjP91upuPdfgsbj
sG4IcShJwtVgVoAEnxxlutCKWwp2OnhTIDg2EdmkZ4O2sQePuLEa+C747x7EpzDv5HPckjZyaQ4v
YByM4dzYVXALEV01Of12xn4mVrqKd11d1P6vYVUsrRGZ5s11Co5csEQF9wPRSLG7GVl3rrzPU6Yu
aHZyu266G48Lw5bttRBkil63qcSaXEW/0pFBohkQDxkFax/hWiWtAol7AF5MHIt53uIc4fKuTV6k
/MgIOTMTuUGxP7MeA0jeLKEc/9E6N+KSt/WTVDe/LmKQxdUCtsPoUnEsPmYopN0NumaG/RFT+yk8
UDWexBKizfAWB2NNkcwSs8x89I+p2dNTjPivpgOJjyeMLFquUXR3Xchu83s7E8LrCKmZtZxLCXit
mbKuu4YOTS0sI2nOZ3dnPkk0SMTY8xwb+g4s3LMvQlsZG5c8aVqXgrkHtZSAwq3LlsnQJMKtZ7iT
3iQjVBYXZi8dqIwIpQPh9fZkltI2neEqAMzYvQw+CJI/gEMhsa7aJSq0snXz3G+HpECTVWD03NEE
HeBca46Z01BUQjz4kw3gHKMQ0KR41CiQEQ6WIokeOxaR7nzVSivWQaEmn1TgogxM/kRIpexKbt6O
9ZvCqph6dCL4nahddtWeIeC90e676ZwM1NbtNpupdrlxeIcafeOchIi7gBaMtCZGhaIoWjnOx4ip
wJcUxY87AGrSfNLjaE61CLIQj5xlc/LVCwG6oun8YgmdrHY6mdJVivJaII7feunGTSLAj/fNcfjV
3SAu7q+y3xfwYYS1Xr0LphVKcEWnGKUL6DKzuI9SPnqExJezQjozriBTNTmQ+4a77cgOomlh6CuH
YSPUmU75Uq60jppZzPJ/tB1czhaEf9hOf2DPC7Vvjs3+EaXtk4m1nI57DM2SBsmUSsWYuT2DOmmm
Xld4jpZ5/gJ/zDeNBtXNhaRVJx/iREoxObpdBEfI38yP6V/sgHOMB+vh+jrcBMF4z1fhbqFwx/Vw
1Yo1f4S9CCTPzs7/eOUEpcp3xbiro+U4Ftz0Fpy4hs65FEsu6omZTd6qR1qG+/T9hoMDvKdCPR0q
ScfQ3kPewnzehya9nbdkQ89AAuNh0QX3aoISvubcSxXD8/jI4I71KCHOZWC47BzlTaTpr06xdFTm
DEjJD3PLybMSZGeWlmd8ZXMgB5QF7W7QbyIBW26wyoBd9B5AtDXqgL4y4aKMdu+qDhLq4Nf1TDvQ
GOXW5y25sAaDeO9UP4slL/Y7QVvBVGuMqBDMeZQ+KKRxTbeXqy+6yv2FW7WvnshLGB67at4qiQm2
nW+3gMsRml/tZknCWscANDvqts7gcPAVhQJkudjE0uq/K0bXCysEfYGAyAi27FTj4qwMREKIFF+q
g3h3ovGEb7wiJafm5aiz/aSrE9hcD4995ZoIXI7BkQ8gG6JRChtguI5q/nVOfowSuUT3TMCJq3KU
y48Qq8lFCE1ZVZSyvMoTxz20IpaVkTkRhPkzjt2OVJ8XR6jqBDzhFfBLgzARNFKmI1R2CMpvSjQZ
D9+V+JbsNdCDno8zDFLh+e39PV9uhsIl/CjjY52VvAjHwBYdPUM133gyn5zV//7ZuvmhBflhXcF0
FLOE0cxp5BwmSYedsbPQ5gEJczoxaMMmRYKIk929Gmkc/G414UYlPPLdGNhe7L/RrqhngEG/3nNU
kYekW7Q+fOYu5VXWQsTnpBztxKUXAjkfnnTiIG8cU6x/bOBgco/1SmP7ZyhhsmdT5wxam1sq8+DV
G7guPhaop3TeQ5T0icsSZ86zjaC9jDXxo04K2pYUGBYXyK3qZJyGzcqFWvqLvhwVhHS6ylbWDJRj
uUSLD4py5k+KFTlOHuJpe50RH5F76S+6ktN1NcE7u4LiM7RakA8it5GFrxp8p8Nv66EgW6I3/1wK
b1+8Ea9zx5/KjNI4MMead9q+6rAVYVBALGROeACvVXWpnI2Deg42jg7xk41CZX928VdSO5U8F2dL
y23Tou7bhfVnRVzO9ubaBDowYAfNGlYOZs4NhM2JRhKXVEVOZ3Vvgo53Eac/Np45JeK0zxL4dz0t
kR+a+h1xdD8epRSntKZQ7GOuexitwCNOL6KpFcC3SWiJqrJ4uMYtYFFx6FDgV6LeQYqB/SUJD7Bu
Y+3JRXuSsp+xnRKIUhE+N2qPFM2K6aF04TzYx8FQGrXWD95JyFkEnqVT16UCUPS6URHiwGyKoHnF
ZXUInzAXcZF4tHLwIn7MvnRWNVZau3F7NgBY6OGVmaZrZ60HJTr18Jx8GSO6+zwX5T60C+WFXGsu
lwEXNJ8E/vZNPFGoHZXa7ct44JkmPvn6RUL8g2MVS8c+Zsm8zcsrlWC/SrFf9LWtPwUgHGQ0e+5k
gn/JLcqo5Hnxu5b5bF7MdtUrFisNAJ/km98G5DvXpiF+UkyWUY4TeXa8bRrNSM/LrAahzfmXQ2og
CSwe/Rzox8BjwHHQeVfn7E4xzSlFr93P1FmiiYtRRyvyBAvlcdClJIeeEaTuTQ/8xJjiuwHLDh6n
YHgTVXcoku2lydt2cV/EWqXN+vT5UrypQ6ctuh+xI+lnKZQvAQQ1gnLGmzuqgDdsR9Zv4mFtqqf4
nmOZnLa1ykWqNMLvTdC3OBTZzXCtnBF2FdKNGfLsTlbxJGhtWbmoElPs+94AYLoOzXBEwoY0AsBd
GjqzGoyAd8UWmKN4MP9KNMuglhucdpwFUgGiLiCtRpu7y1FfQvD9iFxDstfaT9LEutuwEKgGeBPK
FXGv1+aXEbxejjWyd9Ih+8i7cFJXxiPsBScsUd91ZGcDrEidg0l407+u91rIjmsx6vDWqiTqj9NH
EO6GyXpOZXCpku7JPIgzn4/WTHE8j/czutO8IMpYubR//SBigN+aFwsizi2ri9zVj9RCWpyd2JpM
FSPGrcB1AFoud6kFEVaHdRkN9ZxK/nHJqsy4HT75l58MS5g2Zn/BAIcWsPdM9Izyjf0muf0s5WQV
JwG5A0ZjDAs1AKUlVyPrn33JSB0vRkYtYpmFa2P7+Y0L59mvOjaHvGHB95HEakl/NTTf2KoDNrwu
P2PQsqiQiB78FqJLBnTkrBlvRpXdTfQDwuYAhNFNkSZDkI+54YoaFOLmetcLI95OQMHamihlUWSJ
z0ev9ku0hbEqmlMtUTQkRocfhT5VR52C9qplY9svn4vZIvQYBcahKF762JcCDmY/+VkjrB4hVmGL
gaJJLfQsWP/mWDZwmKpZGV5NsICPuORqfYO9TR5EpPW227gI2ViywUdCE1cPzH87rwY6d9mxgEY+
h6nnXvzRRBexHxr98wl+Px1hRqmISjRsGlYD8T/umQH2GBiebsx10OmFp89UE4SbpHYetIbQuxNN
oDtnaeFmC4rrRqojQjtyVCU4dzpeN3ihzT3hocpJxCLMsObLteOwUkUJwkopFpGaw/LMgt+vCVVT
FPHRH2dUJPolbdyE6Bi1ZmS5GWMZ8Hb6G0dOb+mp5RmmnYic3J1cBlDHZuxsKwOvq+e1D6Lulzde
aUQzTx4nwKsdj+VPXp6NMnf7/IUPDk7UkU3ns8+0oZkzHcBFJSxwuym9SAtezzmeEBjITNAZdLJD
WCL2xWPbfzJoNw5XMOgdckKV4NSFMvrffaOtYERTA29YzS8oM9EiVQnu2ddETq88pxe00wSGCINA
jXPnY7vs+8z0oFhm+h55Ghugr+swG/z2Ad+l4AjSd7vuiPjI70hWHAepKtVRSlix0D2QY4birssR
CjFRZ3SEFJS6KpJ8A3tNHS9VGR3CNoTwqed7WTgrRUFKaL6Cu/ofFNG68pX0aTXddMBYFGUNlSvc
GMq79Tq3pDTwRlwL7KTupKh/MmImYnt8YrTIA7OMwBNgF27SyoYZKjQvZrCAsi0+MhakEjlOVlhf
djhXX7kBCeYD6KUMPcs4agMbmH1wyiJORoMEJM9Z8qb3W+qSkw90kZ1PxRXSAIPoq3eMXv6zWXKx
H3uiV5CLtEyxIo4fsmu8Lma1Jc/ruV/D6Vsfv/TaAw5yZnQItp6yRNsUlUQKuzZiLvSUtEwTxn52
f5w3pws3wAYYR1L0X5H3M1cWuytwcKPrY2ECcxFiNes906b6MgUBd/0ZB7CnLntf9b0VWodLVMtr
7+VluiK2H7mGn/KSNTS3Rl26ZR041lAinhikEqBl1pzxsZLyMb65edwsEwE6rFnU7UBP7rrPuyi5
rdUNRtO1XE2Mg1CPso1kJdnd44XLJgG2CcMM+nCnWIQBpPIt+XIzVAsFv7P2w3CZYQgrIPppq6fF
lnX5j6ed5J7bmP4qxWtguNAwNhTMip1P/L3HnyQMOOWVgbang3ZeUmzTRBf23HRf8z1kOAYbFCpg
8qdWoub+zENadvgKnC3GRxyJOYXqL5TYsWjpXUgIvQfwwp+8wfmRDkNCeTBbSuQYp3LI179+fW2h
IfS6DkQ/kpoJsW8+nfNDRoyW+T2IeILvXuJVY2bYzlX6gCteOFVquxs/0W35tHLXqinDrWd7twkd
fQ2Z0jr9Q7hj0WmjpbWnRIHVkUILD8pw/IF+Ap72eSOXGaDgeMDDnS4wx+U9gC1O75ePYP0r1c/4
5KZLK1kJO/dCKSSkPknBkCuKTlMA2sGyUTq656r3r7C8v0U1S0FCtzbxv1ED6p3BsqDEykOZzLST
XKCpwnCk8JiaUX1O+6o50vx306vo/J9Oi999WDPEogY1GtgFieVols0QBuV1W3+XO0V3siW4itoi
SL8MFiup5jNYkFXgGWIfZrHrODOFY/zX2xYtkrEMnmXHpbLdWJVdGfugiHf+Wx/o3vCpCsLClhsU
f0jHqsED0G61u1EsrTVEnDvFbE3OhZdMGHfGIFmMWdrNFC+afj9psLdAq+eDpNlRRolSdeJz6NgC
RssKt3b7lyCqvupbyvCejG2VjjFtu/1yenPUyZ/uZWnH9urf0agRAP0wXXH+lEgrLTVaw9FDZEpI
5qSCdXqBaSJMfMT/IxSQPRGEj9VwuGjbpc6OKv3+49rJUEBYiRLtfhpNzw7KlTPSEvN/h8Jbanm5
b2xMRx039pROGKruBahZ86kawdt3913TO6CzyMHiOVE3zEncY+fR+WbJOaQF5fZSoPFSWzVJhHcm
KLbDThQY2AxTTzxQEe3jdzw6yXrPokjr1LQUBg11Z7d43pNMci9+sYwQdQg1QAAviFd8WhIu1SI+
B0qLeFS00fhda8l1YlCtpimDSW+Jj5LTFNHQN7DxwQlGj6l9lzfNrtrhz8n1DEtRMG18QCUuhiEY
UgDycyekeRUCoyOeIiuBn2TuMVuUaF3eICCbbfL20fuKxcUelqeeIJ0Rrh+1+W+/4e+XVgW+gTv5
GmEAocOoKm9DEeFEpA+TX4wygqlSkHaAY39HzMBiDQBMHHc/16bDKGPF7FxqInFQuWjl/BaAuqOq
4hAjyEIwP79+is4/HgF0UgY1CCh0YofbushngiZ4CNn9+qhW+Bkg8RdyUR/kUrEa3skoesxQ9zEb
XrpnCAXRPYOwuYlrTNqMvxQpMsIwgVNcM9nsW583Bd1sxmNM66xZ6eM6sREWiLiklFrcC6fhK0Ua
hyB22qKiqEQRcO8PEhLQGT2m3XbvjPrwj0ybuYcpGWgck3VtjRFn1uLlembjyiESUgvhJRqg9VYR
or9hDVCEYJW6Xlaj9837tS0AwiSYJzGJ4logjl/ayxcb2cGAMeXOx2bLmGfrbFgNnFv0QVsBUsUa
voiWhjirsvOIsEmdXp/hB/hWHeSNa/DisU1s1VMWx5ODqjWtELl+hj3yaLDE7joEZSPQ5CTgoLbZ
zB6EeQ+eTSNpjEKelfzXQ85TPZ8pdycEajZiBQWLG1PKHJxeTMgMyVV4qDibgGAOOiKnGKWSFq/P
Ra2bPIaJd5ey18ut+h7bF/PtfnBLwx5rM5NJxK1vodkUkVvzPH+Sqig6w5ImP1+qYjnd0NurJrN7
PoIoKaK59J0SOeviHdj5HnbGAdgB832oZNiuzYNh3tyFhpV9npirCdth7Zqc4BLMRoeHpx7r3Vq+
ToknbWFylimyFOJMhDDFbSS/ajjk9Mxb9ZPU4R3zp4RK5287NR3kXXOngILrshCevgHT37/A7T8z
gjN5GrFNXlLtjqzcFRil2/C5NWiTgrshkDrXikpojVX0JBNqwYnZaKRNMGoC7rVUnTY5eJugVJ9Z
yjCGBa00lTH3UvZ5wDj1yleNA90djNwvxsyQfGbBAS2m5Pm5dXkTxv0rPt+wUWs/m12RE75iSpxN
Jx8nsTYKaddrMyZ43BffIPQjlK3Y5YUAdYNVXrWO51M84z286oWjJ6+7gPsmF8GttwGbBsPgSQdn
hQJNQLL7OF9dOmBV9aQQyOwDKIv6Pa4tc2nktVaDfnqglbGmGihFQx9jnyn8ZnU6fTxZXqIFmBhF
jZ9psiheLwUHAygwxoXvYnBLYgc4lWZg6CDSPov1zi07SQWsTMQoPdNn/5ZqcT7JQQA1XqKEmoPO
gPCgJqnnKbtFiyMiJ59ikCs1U/9R4EC64fAZUYP6qoJldwNj7acfZAW7TtpeMiUQSlm5jFegJ4rm
C01Yd0snUEHu5jAm1P0Ss0oWXwBZKlY8YRAA7GzZ8mnt7yHiWw1GMX09dlD7zrX55VoRxAX4Zute
5YeV893mvOoJrP1xJG7jB8kG6TFDdy3kAxvHXkxu5s19kQnpRwNBTYU1x1fJ53Nh8x6ItfR4fzkh
Jezm4Ar5VURs32ovkcdm+yyxBcb/H4vVEv5tz8yU64MrineqrIuQcptMVdx2XDny1fgy5doMPFJa
ivyyOYSzvzlr17yIIZ+9EM7JkCIRq8tYXJZHVFlBo6er6gGM2P+vwfrzGJAWUvALgXCPdsNc8AGB
Z0WM92ppyCd9oOnEhE2xnQenrhbWykzysze41ww7I97Ev5HzsDT8NK3KhuwZGva0GkNmggh7ecOp
JiUHiAyLCdv/aws+nxIZc+BS0YA31baLW8KrXay8u0BlW1KrFpiDubGwOq/ZUz3va8+XRJWqFMeY
bLod4e+qT0IeeJr582xD+CBboXFv7mJdp1pN9B9FaH3ktFWAqcK0FUxhAcvONK7goFgBKoLerpph
BqqpfG52fSEQ3j5ZotawtoBgtGw0HA59MhWROcQ1tbebnbN/3dMZcDs9xv0UiFXBQ11p+SxQlcNh
WsCpWhM4/mLt+ync7pTFYl9aWiywT3xlxoexnNEbx99MTuISjHl0aVpyujK3RCLtzEfE3jXS/Ga9
pdXKRmnvji2u5EckE9P3Rk8SyYdxB8mcn1kgmDUp2nKtFj0IkbxtTn7wO0mPF83orWqKtC/q9dUO
v9zTV2h68ETg3S1FdlRUHmQdjFRU2OvjYwcrPYV8Ymw0zN/FcoXic7/z5XsgaMQ8W0jwxOdAydZY
GDhZ/HBiX2gN0nM0nx1frabwY/PrZUeDmV4vkCF24Ir6pThkevZucpO+wXI2nG9zgQfKXGOsX3Rc
kE3Ru2qktw6VlaP7WXATBiQ83sXjlf7dBm+GCwbnD3XxWsXdQBqeHeKShgR8/IxpIYiv7D9r5H6z
Nho2f79yHKXhUrt328+P49hvSPg3PVoKfO/0k7TXfGhMof/2px25TmKK8OLl4gAggknLoh2pCdyP
yNJ2N8bF15vDZfqJTVCMMMNejNOoAgeygKen4ordp1I1is3YOBDxGwmKycGsrQZg/1UQBDTTQebI
3eHjW2GTlNhogptzlayeK6OYW+9GkawWYbShEhn/fBahBIZ9qDegySfRQ+9vLnOEdywezxoRL6WQ
FR3rD8lg8U+QD0X/7MeeOADhd1DkfpVkOoLm0EAJjRfMEkNhHBNXgXEqZSy8UDVp5seFSu1IFXhD
o1Fds6rDljxzWVQEqo0d6CFKJGAVhJgspyjOkF5rypYCbaqWGvB7x3RsMIOJgDYYizNnr1Ca5xqS
1uTxMvWQn57hFRABreIqDU7rTvlqwW3LpBQRau3wjOMc5aw7BMv4vXY+rzoq6a0gwTp9Tf+77aRR
eZi4zdE00HcRbFTGmmDxT5/e8XA6e0XXcDgHXslZg7hB347HOmzc2HPCTup/MBtQZccnn5UH8xn4
CYz/63tVscodHY1NaznWfeR/1fgULKm6/9mPiOFY+CUqs8ROE3fRBZjINr9mwBsa/qmqIQPlRIhl
rkCqJ9wFellrvRJO/d12nJMaQUw/3qIuhrx6KzPkrSYCtMlUe7yjecr3BBVrp8VumRfAcunwzasy
3lHXWcGqPVsmrtEKsN8Dlpjx/PJ5jpmuEQvgcrF/IXEg4xO1WwHmk3dzGxCpGPcrDUZ7w+FbFJF8
29OTetay0Qh16e70Xa67k6IznNAfetao8WwikieTcYjxAWDTmbeClc3dbLzlemiLPgdy5+MEoRXR
PCm1lvZKwDOOAF6kGfC/Mg7hKmYgaSvnKgbVO52iDAkgLSQxAkkENzDTFIc4KgmCMhVJDuXXfa1I
bxdYcpU6Y8smOy7WfkfY6ngMQjfuTG8aszWl8/1xH5q3oTbDPOo6lBX+6ClMHpO/2VLvMrAEh1yf
SuhJAiMdq9bvQmiEa++Ly8Vq5e8mpQyBGjV8Hn4C4BZaXr99mtu8qmXrlALa7Rh9x7G7Ilgzy1XN
hxj6IiIYZDCS5IUvMZ9vz+BvWMAExpD1y25SmUebt3DpD7xhrdYy13rYek/+vE2aD8O/gxVNjSAS
krwQTe5IKeGYvM81PMw9A8yzqk8lBLMY343Ti4BDailgqZfd9b/FPTQJWbCgp9IXgDtxbWhu6EG+
hu9b/heakfNA7Ops78pXm+bLFD7uPZYaKcO0GxCapI2kSd0nTjrXd/IJKrZTwv68hKWQ+Hgtw2aR
9rLymULt8vGv+QsHEI+QpOFrJ+ieQI40ko3eIupPIfv6qkvt3BUggtQTgnZaNcRy24sIuUF4r3Cl
xOy2Lm4i+Wek3q6au5VZHA1v0eyLYM2yZdazTKPPvPkY8k8ZZrVZPRjv/iPmWWVn/R+qmZKeRf+2
EFiiYQcyKxisxTecbZfT85NGkITnGROXB9X954UjgbyFO9WzE43ivrdpdGaD71G9Ef4m+TUOKoQB
63jy5QwXeGsXs6hCKgcT2f0xFj28T83P2NjzCRbXARl6yLMkRtg4FQ8fI9NuX3jjWG5ru1HcBPrp
ogNZNmYWetzHkO6IxuCEQBbvn+97FPnPAkHQ3UzcxJDTv/VPNzo86fJaGuAToFOLP7hguyPEbkMo
tnCiceA/egk8depGXB9tX40o6PFqTKDDmWh8cVncgK6WUkni15VufzK+2xbdHvBbFNranZy9US5c
iCr+wRkfrjVdl9jnOqmED+ajQ6UsugU+TwFi/W8DCPRNcXjYbyPSnh1DnHpidURYsmRvYzeROBkG
uoQIpQmC4mMwM7AyDcNjlnrGo1KhQd3m/3QVGwzWYyTnfIV6kENLlry55S3lT2knqUa/k1umY2HV
m1URNFAeHdqfpDSbVP/wqokkt668/aOSAF703INREx8u//5kosxOrl3kjpM3vxxD4YyaPHP1z2WJ
mzko9lUiTVwhFQFPR44y/WDT8x4DeglrvtCpPABmPfcLJsK4a9PMZ0di+6eksqSplsviSnD3eUpr
r/N8pZChsz5faVklQZJNkbYTtisP3beaVSDsftwtzKxFeM9JBQfWsE0jAkhEfNnaY/oYZjb1YPZg
vysEEdanDTHNPO4OKzhYR253dtuRURh48FAPe1REHmo2jjPLSvKMnMcnk92ByKeS1Xu9JoSAtAgo
cd9I7gA94meL4JIC0c5W9YoT9eixvY/1BiUCoVrxUQBoUPpbzPgsFcBCIdwPO0Z3Vxxtul0Qt6HV
ETsOQu3U6NxRclMkMt3UtSYt5FmiQzpjT0/nFXX2dpnQeYWOAmPED8YcRzxmNfh1300KiRUYuniK
JYPk0Cevu9cbjZkdvIjU7icYHrnfU0cUQnU9ZEg/r9yPYIiTWdNKGGUt9oBn70PErafqqdOcROc/
/zWxjQ7w+kdAzD4p/x1+4bHrY9Wf0y9myvSMDyuzzIOeuSoEODQJofxaPtIe+rzob/66qWrNG/Rm
m2XKkmBvGLjltEL6WidherygJ54MsQLcqUCsqxcJUB9qMMagy3YV/JaoYIuBxAciVXbfjtPH2uP7
b09Wkq/pyxwDJUhLLXi61O9+3TMSLeE0uzSxGgk/9m379p0CfBaU6+I7eaHBh4SLjtTaOsJklWwm
2OPfPwMPomYR1g1urK6k72j5hT31cQq2wFn+L8KmkLC49Owq4sOUKxtRr8TLu7oeQN5IEe7Ix5kM
LU2DGvDdyfdVqGKwHX7bFEpkPODgmO6scT3ytaHVTTz5AT6moFPn7K0e6ZllGrAoXAbiWv2qmCkw
T1irzNtdvy7Jd4xvUxBtendDdbYDiUbvWaKmHUfsZ9bFXorR4i1iCbsx8iD2ikNwlGFSCLJyoxDm
1UQgriKBOBYFl6VrlK5isFCtA2CluonY8azrL8GPJycf8cpjtIVhT/nByj9ZbHk06SE3sHmRW5g8
Ku2Vg2j7CDbAWj9zH5d55RMutAyA8MwCHhm+FE/1OMqI/DBCqo1oa7+nv2e8GiLI8o0ywyJESIqY
UXTrHiE6tONdIn3K7bQTvzPp6r8SbfIrxcR/N0QIUO1Web6rqRetKsX3W6oYQy6KAzydN1My04b3
fdXwDJjlTSL3+jIRSSRZJcB58sw0/ZANOClsXylqvSGO5SgWOx69mLogHczGrX1Gx/AL5pK1jcpH
9cXMR7Jv6oYxC9+o3A+XzDiIuUHlWAVxuhboB4opkztZphKuRhCRujLVjtyDDzK4EniLCcb992X+
OM1cYCJSwK4X7dLzeMNuSONm+XDtRJJgE0T9DhsUAQiIel6XdhUOFGhMbTxxzrkenPjIMM1SfI7r
gVNOr6nzZ+TI08zGtxuvkoBzHC7yenfVHqZWnUa7ia2k3jIvaAtU8Uzrl/LEYFq7MJAhXfBsAURl
LEaqMvrjYccZJRwCIKM3Uq9vb7pAKLItCRe8+63xSFJiD4SBBaFq50OzBGAmGRuD2uepscMv/mwW
wUYzeMusA8fOTOAjidTvPw+d5F7YlRhLNowZJ8ii11HulDWlncgu2axkk6DPeQXWqy87PKNn+Vpz
1PcIiupupKW5rNh2gpR9WqZA6aONWlW3RhRTGXJVFXo+oygvjmeZOhTbPTKdvUAr7CTEW5PBlxhY
XZSYgy3RmfRNz63bKJxhK/HHx3Qo2b8U0rGu7ektmTT8uSFLYuG5fa/1BBLQKVsGRLdwuVW2A3wb
bLY5vrLG2ZVDduQAwD/1oGqOp2V//Ro9EvDsoqqXW9LpJ8j0hX5HQSQ52R/5a4sE8iLDW0hARd1H
3dezuatOq0IWSHEk765skwRBumEG5uRL/w3TVexiyUwaQRuQnaqeeNfhH+QZ3E3nMKv6VFW4mnzs
k3uInipdIEGiAwqYB702mMePSNJGSgNp2h2Q3qhNu2mbY6pkVU0r0cPpUW6Wea0fJgd253/zYECL
VLCvcJYSe9Qui8dzwUNR5e3AqCSHgfXDk8kyqFELtqTx7NyLBINMmpNxI9OCuZHxYd9RGSQBLVzs
RXHrjvE1z0Pj4YjHFfpcr2laKDaOtjVHa41V8ULb24d6GmbzeK0lFEd00+xvrsr8wuexRT6AStJy
gZRMtwTX8cRVITzMprG6+dhTcvP4pxtQL4Mq/5bad4+Ektaqlvgmb3nVPVVXPBJ4qejxfrFdoCaF
Ah4eaN7GhUA7TGlI4K0ZFPQfwSka4Q7Evz3EEuJVMryn01Cu6RX9PwM+3RMNOU5xDhI/kykB/Xu1
Mr/Ee3DDHsbHGVfZg4ZaLNeMd/kjeIUwG59PeeSo1/V0JwHDLnJFbxGHg6RltgxPiX5TjX4OSDbZ
pL8W3PTOVCrenuhqrr9yZWvivL91PLaBL/y29D1LfNbYBI1PkXGbkZeQgAPgxhFFmiRH2RKYwGhU
iR1DaNvjasFEZOBjSV19+nVbgh1nxiSrYmspfM17GQy6KTjENnfOrwl+OxbVH1zjQUKnjTGSr6Xm
WF87vAFWn/XCxW5ce1UGaVPc37ER8gEoA8QWt0uyAEMnst9IcgWvXPGNTrap9FK/82Tk2NJb94z9
XTD4yk/Xd2CRGmBwtE8Y7hKRBPgfr/tmonSltYSWK6q7iT9Y3+ZxUiLwBs+VK8yW8ap1NgBK1zfQ
FLp9mmG6h6IhlOrqnjpd1UCOP6ytRGeYbQ7APdGCMriY163oFKvCxEYgVYhDZ2k/KHB8w2bC63nP
rtwI/f1eTO8OPlOXD6YTSwEwPUZOrnikn4Ux82p2y/TNq2t8mqJipbBjbnshvQKWkABUDcAIYgB3
k7TN1hWHcTONGN81T+UAh4m5IeO09KRICKIc+jjdsDI7RGOmvwDJXJUsa6sw0L4euBIafm502AWy
CZ3IXSlz5M8PRZQan0hmKpgQjutbZ5d5DumZPAL+c8RE09m2Q5YlY9RTKMR31dHBMh9GFyxsRG/V
IDa0LdMnHROlxa7WP+T73T+bmObu609JVy7uqfioHULAAxRoL7lYUdkv1Ps1zgIo5WNtc9Un69T+
jkQiQ2zwhs0/tLmQMU77pDJ6+h5wmaUNNd3/y5ufzAMA+PJY/wxY3ilp8MaUy8O5YFrAh+VuWPg6
c7W6jRqjJ0XD/j1NNqcnSPRtILrtesReiWJlm23pF/SRJCt6WyquTk0nX6ajthcUKPqzORBQWqYy
KGdnF8kOOQlB2ww1NrEjyZwVbarO+pLsnhpV4V52Uvr6krbujYd8jxmCGWHSoj3fWrd+bfiimO6G
x6pUw5uKeLOQ3pIW6/MdFobZbI+MSR+IvYVGy60VspHjO4ZBSIe6l+8L0Agecp2uk65w4MZiQrX9
b+OXzonQkVtktpKS0+nM4P6n/ssmWvRT5U6gccOvms+rlKTYBldnmacGhur2BOnA8XTX3PLQz7ns
RMWkTZfGKtxYOSie7zv9S6m229+brAt3VxDLAFDtSoSJk0StD43SvT37wR8+3iHauqqZAg7Asdgh
RMG7CmQRekhaZrMFeiRQ4h+PdgxHbDWJJ6GarWCPeToHxghfMZ9yoDIVHe2BzsRtr8Qefppq2KoM
po8rbdynwfl5hsu10/3WiFLwrfLG2CsYZu7otoh1RIPaj8gg6/n9A8Ry+euBexEp+rUKWs6wKZ0z
vZ9M/3CBZuIyUsb3y4g/lISfX9GbOX7xTskqamjdlnb2wgBZmK7fMw4jx3zRI5pRTMENLIi77XQJ
Kd8R9FP729O60NI0w948xFKzo6n0Kfi4FzNuWCIiaeA65fGO0eAMINMQ1FP7hUWDFOeEjUuxOiuX
hhAFIioXByC5WtYPu0BARpaLyyJfw7a9gSTqVvxgGzuS+5/e4l4DymYO1CE06/m0qGSiwA6TTxWI
XIUlFa0i1htd8pqfT7giNwxWz1GTXOtvkr76+1M1enyNe7s5RhTWncMVQ16mz3Q9Eq8IddJ+ZwPQ
LsQNFTygnqXstbJFkTDivc5qrrudrN5/cHeBiqOgEAjY3dWIuv5bzb7BNht7CJp5bUTuD5GMzO+X
Zr73we3CbhCDq0/pn/8S/yRe/BZgH5QL3jsKw+9mZFeDV3k+VSqD/Ye0KuFhuWymXWfCocl2v7G9
qcfH+2OYDQ/Xkijbok1k7hNWkTvePNQq4N7nsBqfyMkijc53GCZJJFzZ3XKfgIf2CDm75vJLA22f
Y6nCXrGyi0MAmgus+UrlmagUpDNre0z5giP3nDxuVPav4RVttLISWQt6LbP2MaQolidOUevAhluI
O6V9mZFDmkawiqSWQjraCn51u5Pl4VrE2Z30gPa14gihfTeRHnvew1HU3UfbFTIv6rU5wo7QFuXv
qj94Kws4fPiAk2d0GWCAzz94RJzeqq5H3CLixxeSu9zckmqZICl+/Zz04jHyF4YMaVauw9xJfGx/
2uUPOPrcwIy1LWIE3K7VAZQboeZHa2r2H+pRuEYRSuY59MAnx1LqTL8paGJhvJ+39XSOjlRmieyQ
1yssLSYENGYtCP/3UOUJtYbo2BVNNDtYLIOamFYYwm0s194YxxDR3rcGbayihWA68S40Pfm9L8U3
EhTHDcB9Llb04Ax+jFSWx8Tz6VDP+LHruMgOV5bT0ywKXRB1HpY/xaUe9rzzXK2j9Y6aSFGoyco0
5YNcccAJTLUhQyUYOWSK1nuj/5/OZz1pwrNd7zdPTPQd8AdUX/xsHWIvrFZ2HBr0PrzaSDCw5Csf
5Q7/uBqES0bF9veDz6FTCkWGDYxyr7Z4dTqXh+aktZSpDi01qERgEqVh+1ezTNeNY928+FwGZ6o+
OUszjqlYfCygOV3gfT7uLaFby8qKO9iAGE0VBLtOAHGuLWEXF/gEjbHGs2URZkOppZLVv8cglfw+
O73aA+kTn9EkW1gn1M4yW70m+uZAGPltzmKiCwActDAqd4z5vOG6Cxaa5mNEPppp598tMSeosrzA
EoVStijCxDLHjpjsLs3pHw96YwD15KDLo7juS+6++icHRET1wcG8hPaQ9KTFNCv0OsJ2Takte8MF
p8+OpGXWazt2z1bInMl5VZ0St6s21dvV8aMQDcxYCTrzm4jPuzxwVunGIboF7zWrxTaErrfyiU3i
v7/J5ZiEgfl68DLgYAY3Ja8NXnGXLQ7+2dKK8VeGoY/q1QA+df8r6VBigig/nGlEKoMpJLo+rw4+
D5RECSNQB9xW/E7A9SFbAQ7KcIspHQe7BlIjiP4XOZTUoyvPVEWuvBGivGcd4kyPMg9q0yLzujh5
QENvqjUycBA0FZSiRu7EizzIn6AOBntQ+9SzwdP+MH4d2/SYR13RTUG5HaF/dMWLlCLDmibpflV9
lFn123Zan/9oVJ9O03syNTbX1wSjtiA8I7oGv6zFueBzUGatpAl0TVIs52NM4QD0KUHodNbyjBHP
fnP6oJj8bKgs056SCeGyntMXhBpv/x3yx5r03BKDTQ7KWkEHa/wpPcfxhGui0L0Q/lbagSXlSBkD
RkCKFpQ9nxffCCAXKvLbRN0DwaZ4P/uNi4zDlc0qe/QgKlnZzg9zJhrQZwRPulO4ysQ0QiLgMcNH
JydzQR1SclUYmxNs6jmm4BuLcXSkxM2cYVTZ3dZPg63TrqkmXLLtE7nLpOt5UeWqoEaWjpUzIRpY
8VOg05l6/cFiD5jP+SLyQnwNVnNOyonXP7D+92tvLO3GypHnYIUyAOhG+H40SNaRnv/Lmg2h0hgn
Dma44KVBmdFW61N/68GwmHT8zSQ09ECv0Jk/zwrtU57sYTSwp7aEc91TUsqq9LnpyYJvbXQ6iRDe
+34w5vXIMo9wdred7lBlgtywf0etc6+Kw1w8qx0kmYw/Wqdqrg7q1QAHrYREbSPVOH2ECaCntBbU
/iso7t9HrB0x2bgR5lZv3XmE5p/mYtAG2ihEQoygUxbRRyTpXom5+Yhew+KDPtUKPlKUmxraxXz9
VNvMWumIARWi8Az8fnz+kziuO3iTix1lEdZ8N2g6x1zQGYNFHtQ1UHu2tfMiaZfjlhEtxRKEVK3m
u2uKDfAE9PIq8X1CDOvKLXAUSG5YHxV+Lcql5xM0Cl9JMtwZBLQhIPyyENFlfPEz1iaZW/i/Ohfc
h/y/vonirMiOkuluTMFEJ6g8Kt4zJ+MJOmX6nYA+No9wGGWvj0QxpSdNFGD0oxO8ctN3Vhtz+fGc
p3CZ0LUrCc/YjKdwFlvJDU9BXpAPTapNAV568zBUBmQHmAY+LQ4wyrSPY6+KdGV3qMhjY1MoI9Xk
lx8LIK1P93SUGcBFb1gfQNFo1Bk9Y1mUbFgSh0DC1JKVcuSzBwgR9q7DoGBdbr5Ao4IM5tUmwAC6
EZM8WVmGNTNPXXo/TDGQHSYeu9snQx+zaFYZ2J3LLWl6uV8Um+Ix9DHPaQpcQrcOWYaA/mTl05We
joaI9RK5wjfe45C8BdNQ9Z5BCvrjRuW38fa0pbBFpeoeFZLO/l4Tsj/teoPN58EVKobsE14WOt4y
nTdeqALudRMe6qAXc7YUWCnpgxj8Wi4yw6yVqatB3pCSJvqQjGTKJUDTD6RxN8fQlu9afXEYKY3E
tIMFMzj+iqBeb/vwLCKdhpuNLMLQAc/JdyFXvMbgntdSGUUuDGe0LkpNplzD/MfNt6rIBSPJyq1S
XBTwB1Eco65PzcjkzQg5rvX/IBJhQqbG+fuwwH05jTAaUQFmzWI883Ei5DYLVdkKphQtc6nwruk/
0u8RnWMnuvt2QqzmUoYMXcGLL0Jr+Ck7S5c5RhKQPyw69le56c2kg/IxwM1SxRGg8bhnRBpiTDPm
Pc4rtsCQW+s8Cnvi0SoJJ3GLsgeUB40npBqgBovcKhz9+rHAzVZNRr5Of70wRVRBQ7q+iuBDDGXG
ki1aR/4I962bTr0tu8DNMV5oKEHP4tUcxQNKwi91OcwOrDH4st0mwb54L6BIVmkMmvzVYmF8Xydj
s6KQFF/Wti6BpOrCbsF76u7OPuLQdPtcEQzcmjyDDxNURoXSdfeNQgym1/cjqmk4MCyhHQhJeBzW
13Y6FrSPnNR0Ix80TB5uo/mDxw7Mt6fQUIY8PwFWgjA5BTqSgaAGUFWo4mol7v6roEbBN0NJA7rr
GO0TmLyZ67U65bEXZnYzAC8r7dqWZMpZPQDMTpCAgP+hbP3QvpC9QDHsAujLsuOUKuRRI0LJAYQO
xQHg5EwXEjGWMmZTpQutAvhMEMislkECyO8F7rAUt/QBbB03I+15nCEjq5DjVk3NVe6KAroEkeXU
Pi7c1m2dUt/czdl6Ynkb5SD1u1zjuGJbqNMQyX3S/Q4uUiukT4yrP12PfUt1vwQ01a9HYgMay1NR
SdMbOlCU1NJWSt9qpPlsKTYon+0m1J+kM6iDIamYGnYA0Jke8HTvWuRNtbFhKL/QoiHCDsuF36n4
UwraTLsghgf95Y0Kgfw1qhuKBaLYtjc61O8LTsCoHIt2SGFVs0pZ33RPr7/NwP/fMr20PU0mZ4a7
npVI1sMRA7SNJIyp1tsT87dzZw/tSSvnTVaIrjtfDKMG2UuZHIm3r6vdFqS/Yr68eyfD9NS1COXl
pqv9qNoDGzjsO4jchvuiitzGWPjQI3OxJt790TpRCbx5PO+QlWFE3Wlnfm+6oLWj0lZMs2LOuERP
1aQ8K3R/AcKJ8OigTwRuCvLPhlnC0BIhmAh6Z1f4YCL+rkaZgUuh1pdW/uL7hp84FhusaG+p3H4M
Ud+I2p/IjUZ5x8LKvWMneI0uB+VEo9FhXugMzqTyzDuJz09O7sJhSsRaqNLFtMC1urDr4ViHeVvC
J35GMy7ttk39v8IJAcDmVdK01IvdAC5dWPT5pk3Rd7Oa7dPkKXKobtEHQvl9JgbjkbOzHwSdvl53
xYbZTepsdxoXx/V+rQ1siUc4Aa88So1OBqgwS+JPABcxU3g170qcEb1aygg50u5dIBBdI0knyuxs
uPXXqGSGYnAxEMVvxLhTzhMUKaelEnH1rzRyTb2Tn38jkUOLGOaEUatNCX1hqT5qjtKvU8nBCCYU
fMHSi3WQIwPimNzr9lnMOcEwuIfnCPIFt9yqdI6gDcMUQd+v8tpRgmkzmChqMtfU5P37e29exO7Q
m1j3kUXCYVxRPV72/RPpqCHg3pKgRBWX9ES/FoR7+eguHe3HHI3Gdq+9QhHQ0W2qwyjq98H3cTFM
hEPXvpPMmkqSt1bS+pDIKfBLIVJxxZITC5JTyWb6gx63ooInC18IvF3v+iBR0SIfemdLFiABPGCx
+tHohfw5TogXMFTCDCdhhC97e4ewE5uStDLDJrigYZZOCXC0XClhiwfNa5ymg+iD5IMP6RZBC9bG
v2N4YTUDe3JMoVJ0TlTk/ZBfTqRAyv57v+mEjb4H1w8L8LCRTujXpExIsAFUJGEHdBwpA+5km7o2
Lhc0WPuNNplMRYmPPyIEC3eeOJiE1M189ImJ+1qXzSH2aVFOegONTOj3cV46Dm1rHnIvf4+Kbyi4
JGJeDi7/BfKQYMkB7ZPX6TGkDcBXnzvJT7DTObMFo1Ep0oI+MIibKO+ibxzB7GvE55znmYBnOA0u
RMGRGv4XE+muAvEEZbqYD2zYQi5K6XYYK6NMCS/c+B3u+INGPEH9cZT2Ryuz7bae3Y1YsrICc98K
SgST1iU/0q+R25k8/E14b+JDFK8zl5fWlbfm7RYU71rgKWxBwO8QNOUUoCk50NEcCGjzYcJm3+X5
X8oAEG/vdISDI1IG2fxpsdnP1CixOsSuOrM030h/3QS/zHdbh/0mLw9j9Wn6ENJ1VAVaT0AAsT3G
1NPO8eMON1cm+cLW+XMl12DCQr/Nrr/VPccn/AqEPGtrzvMSnPXGLMXK4I0DsgyHmKohNE10OMq2
oK0YUpFWAQ87vUlnnfprS9BqcqL0kf6G/fcuweEN1+r53AWHuZD6+J//Pbx9Jiek557aBa1MTM33
yUb/CMXUAu3osvlatqbNZKMHa4izKcrIX0Ng5yqtrfF7GJ/aUmgbtHaDOVY6bBIXvd88K35hE/GJ
wNnSzm+0h40urAj50dmcfGpXuSEOAPCARvTqtZVwIY0N6yeQ0ldJy78DWFbB7P6NfMgMzFEzk42u
fRm4CFw3JPwiDkWQIeVJlt4oHDHi4mE1fY215XzoFioGQ2uIuU432VNHoKuQ/Hk7raNP5BW8R8/M
oldSR1zwHoDOasXqMR2WTqXXMVG+C5/YkTLWs3pngWm0mGztDgHqyNm3N6W+MPlX6xZ1ynw7t/uc
yDwomqdkJZPC5cFxxWDjc7edhaGSL66TSHGP8XFGZSKH53EAQ0azv4QWPv4DhanNx+clVFPoZr0a
dpbycUUx5WBKIr4ayugLbgdcPMk2hQ3IbESnXJBDRNkHSsoNwyUUxblQ8aFKIxr8DCLRdO/xKASg
+hKQwNnZuyMUdmPHf8HhMpuWPS8YvnwPEEcTo0RUFefAZETdozHz9Qfeer7lm/i9CIp6W0QJjHcz
4w67nEYGzLlMDB9WaXQi8/ptuqTyohiWwKNvCzpWQYJrNYrTpWenu1n+8LLgSI7LoNsTMEGLFTh5
0IXEsIXB/9m9LM5qmJAaUr8jHWupXB+CwvHG1La0I4VO3O1f8j7zRGQvTMpQQV9/R+Ldvv6Lkeby
tpeRQUqY1aB+dQ1OtQuQAifjHR3fbW29VPHZnvCmyreugfbj3cEG2px3RQJ5Ra4X/imWqbLAVO2u
bWnGOMC/i8DJ5IPGSQ5tWkIcv6T1pBIv0Mq0NMvlkPhVvT02tHECl1x1gHmDNPKC9EL1U6hbA6IN
LbQrTkLet3mlOPunE9/+UlH10XAPWPEy4/IQFQ8Pf6ykEZ2lxzhM55RW0MDYhUQ1PHWzKmjDV7pr
zbw20uPJrkrqP2bkJnER70/6k/GOaw1ao6JWb22F1RAShrpx5BzWnTgED5FABGAvBzozm1cvhlxI
3Q8q+9uUbDDpCnaYmUr60sT72cQjnBK3GYGMykmSb/BA2oGyhrPorQqyAnZ5RfLS3Prwt0FpUQ7E
SmLNiiRad5EGhn5hl08kV5donaBFE+R6tZfIxbF/M1wJWqzEoRf0yv2z/2Xg2rZAN3JYjgRLpHpb
Yp+nSGvZOy+LBCxcVslZtd5pn12vp0sxJRd8xrLDY5IxC0H8umPQBM7gtY8WjCF7X/rYwlImj2gF
h4HLp22KcKSGpp3kyW0xJUQhI5bE+iAdG2bWBV0krmq+omh6tAh+4n9x+CXviVbcYM07M4biRUFS
zA9/Yar0pqgUAg5Hn48KJVypSQplxvmr3WZ4/PtvsBFPg52PkEB/ezgLKwIFAZjzexJasjnbBp95
1JpMWekiujI0I8cLQPm8mmpGkhFnFFMC0wuuAbQcb6BOaOT25p9Oxe4TVndswK7TPVUwXr5wESrw
L0pDV4saGUHxytLjlM43Ay+/VvroJHyYgCNYdfEMWW2WSJ7i70GIRsyxK2OFOPcxHeXuvizmC9tC
I6DwEGRNpg653GsG0Lx9uVRTSHnyLsJqdpLxO1i++I0E0dBtkzMj/Ooivoi1Xzz0hyD6YDRqICLl
BE5TcGHuavp/C0l2NsiSrdot9mumf7hs3EYTjAqLAIwe1bR5jz3FHJT5MnZ29s7pzrvPVsmpEDuX
O+tl1A9lDH3bWPSOPotUbX2tdGtmXhiXgfAV4HjoLkT2r3meo1icdu4vcCRF6Mqg7FUcTWO/r1JK
69SScqf/asmdJaVpuq11FoCxkN6BT0PRQb/nrklzOvQjFoMOs3KA1xMlo9vGYBgloA5T+oWQXlpi
tXq13ZZkphcmf8TAm5kDBrdOUZ9mvkm6qvoi30i67HGfrjqiLDs/BNmAbWddhQtyzH/XXxus4jKE
HwLhRiWUmCALhP+c2JfdpJ5XMbqPOTdRXNAt7HT81DsZEeQl6qGBdruRdJdgmcXnY6tCE5s15qZR
VXa5779XDe7FVvxRWKZaeG7JHmq+P22RMLGPysFxD/X+ZecsR2XiqaHxfBoqZU6wWeiUsIHwtOG1
a/vklZ4Mpi5jo3WPKAsQlRqnSff44yMYTC9rdWWPm0narKnp09u7i+AlW7nOZG7gbqcDRBMHTUYC
zIFzc/5rfiKhKEArut+qy5NZxhArdkQcbr7jUrUJ4JfAYliekg/5Twg7MX2DzMQWaSgdB4r9TXUO
icpu7UhNaq04wp+6LqTmN0CaMSCl5VTqVF1Qdw3tC+qD0d/N5GwEFXw37dSTs8M2Rni20VN+blpH
U6yMA/E7k6iVqOV0l0pvp8PvF/pLzbXd3GqZxkNph+C2eZcUj/u2hpjkTrfePcIArQ1rQk/6sXdc
cIGQI7KQOfA33emqlvmQcwyembhgOZU2LpdJFpj0OHktmNwSUjGUbr3/TbEH55w9gs4i+L2g7wyA
PkYW/NUEKCdT2mRUnt3Lv77+vMldO8dxPVFXe/iFEBdZJAXjlSrBQbS1KS1k43g4NHtDPul/FQ2L
8JubYHzEMoamZxzGzTGd418rQKThxNJE0KYEuH7UYX78hwz7DuY5rzMpswTOY/1XHVLhr9rccmHi
Wa0XJWf4sGeL5uSS9l2SIZKTg7OuZ9I3Y3Lzt862uHJZT4NKyPtuXxFRC3Ra6rvrq+jAfG3BHA9C
nanehqQ8TobJi5O5THcBWgdOA3zf1CNmPjmkbNu7GXFsbjuGEyXDMQNH0r3G7V685yCqWlW17w1h
qN7rJ7ogFucKTxXOvmg+mvLzTTk6DC+kQcGmvhgwz+KFMyFxwS8QN9SDDM/P71MyNCcXqJmT4FOV
rriVCUqiTpb83p8OP4/AfCHY73/zbra7assJTZO72gnL729LExWsi/Y475NWOpPsov6/4zBr7Sa4
FU0E2KPMBfNHAe++hKlPvdJvsgRw3e8fKqDK+hUDAEiLYxK+l4j0KNVF+RS5OLEZDo9mV2EyTswW
TTYv4Ne7Hvz0m1wDY/vMUoEd/drjr7Tp/oT/QGoJCxkUK5aEz7nGPc0Gr7XtqzV7qJk5aw/JDcSI
dcUROhWXz+hs7J2m5rTCXWa5IshoLk6nJoG2+9y4CJf8kMGA8DWHEVMuWlHUcRSB2nF2wTebP+Ac
4r7iUFJpipnKF0lPYz0dBenLF0XN0brStP8c5oTL0/pB9btuYZ4z4oBjwy0oe5SYGFku4nbzX4uc
oDzWCZGHPgEfcrMBJVO4pj0WMxNvmY+LYJYRUSL0wAYU/in/6jHsW6otElWPzcauxFsdJW63MVNb
mzcir37ySnmxQR0EvfXWznHu8c5gdJZ6D43yuxFdsbX2GpHNUuoSLVyuvSpUFqNaNwCMWTl0ujaH
z/83KO9D+Erc6aiWd+3kAnDo3+wwpAeLjY0vvYCmKAobcrkALnPWbu3cRV4yVfkvqEtaJsk4E7Y1
6/iGtUiL5pF2KoDHDzClGFHjaZ+/R+20W00pgmzveEFdQtvvp+qXZ2WT9Zw3L+tA7tCeZ1YL5AOq
hcDSZNh5ByMMlQgT1ZCi0dMMl5WWKjK1ZTqDrwDbli8N6fM/YBcMVsVfcZt3zcjBNbFInZTa52Pw
sqzaDm62MfgcCPfiX24v/v1AC5bsNLQtdNApSRKIC8Qihgzr9UtQS+pCdiU3p1gEp14bzoCmMyM2
Oe9iS/osGtGnGRkwM1wrYkfxOY4nrVwd9DchUfQTGPR61Bng9ZJw8mFlq7fmvNo3QeWXObIrMPM7
cmNxJZoRh/kCTnaZdizrSQsA296tQMOiMos+Nh6vnu9ApL8zx+nd46yg2KJH6fmwPDumZWX2Cve+
p7iuGSK4aoI/kuDUKQvAG/ew5c4nuFIE0oitcxx99izHk6IMrb4wcJZWHxFvTSUaRLZyOfp3bk4F
kZnQufyAVp3WIeBoBzkh/zibIjsNrGYNrdGj1lDlwtSIyRKDg5Sf2khj+DAiSvr4PpaJ0mqU6hoE
z8/Fv62fn1sOA73MwR5LEjKr7P2wwpuS75l65LQRCxA4vj36/zRXIb3Hs+oPZWRamAFtJSlodD/z
EGMyi8sOk+3RKsJjlaAjo2Srsv7eZdfBmhapVs4csiGQYtOhNXre/tpRa0aJGccsH4u9taALhT4y
I1qyIcMg7CldjsCJ4gF2TC/8a0OE36f8dDu44eI4NmD4gbpjAEf118POB6FADM2+sYaWO+JGuokq
REAAKqiK/0rNDMHymDq7vojkEsHrjTXlbYybUXAeh8y09YLCcSnlHncnjwQEm+NY3C7xqzw5TwO6
BIWyCxA+zfuZDsI44KzqvIjhEif47bLyYoyPMSfrHlApmAvMy2/hmmX43NVnqGROarWlGA2umSOV
5m1iSsv2tqMzX7hAfRra5u9+uPaS1bZ3hlSYPLPzRBAlx8DjLJ14G3P/ddgi4VONCRauhXU1bkbu
t3hACfTyfyay/S9tk6D6Pa3C1odDG6C4QlzctBL0EL+jTZkbK1BTJkV7TmB38Ez4+/cbRoEyZYr4
XNNobK5oGfkxa2Fsj8GncimIiRCJvKVVdDCeSpF+lfNQwaVn86QGU+XQYUFWeXyoLIw4Zy3a89Pp
X3ZDVTyUnUEaeLtKQygCFlNisyKkEzl/Vkyc8alX/YinTBoSqsY7wyP9nLpbDnPMW647U/n0igGe
rRcQyO2FEezsIGSsIbck0SAqOB0uo3sTdGk41YFpSbsHwjL4dqcnk94VBWFHIhKhpdA+vokScK2o
Kxka1K2j3GWjwQERSX+APhGP6z6ENYpX5NEmvubKXaNsfdzBa3ViYhVEIu9ODmre+upv7ljdIuWd
ddh9Mj/khmd0x+S7RW0HueMUL3xTPTKRTpnzNAwn5BycbD092YAM405AUmNa2ZxDeegU2HODUm9Y
jWkkd9+wY+De4tFmfGuU2glG+oJoC/VWInr4nciMvDq5wV4/UW8xL5unzoHxD1isumTlVxOclAzI
y3EjslbKyjCYQNPDKcT0fbV9Qs4GNUsN/apKbT7fUEVGaRVXB+iwI7hacUg00scZ9Y/a0kuPyd9L
iyIA5dUJr6Qm/GSTaJtddB43eRnMOrUT0FhZHRGyqa4+0E9aHWUGwkStS6fyI02ZvbSMlP2zUnvm
Cntz8RmwnDmyS5rPrfqxm/qEvzTQIp/VtBv1/w4MrK7qjzADZFDwttpjw5XssfB2OcSrJ5rNMjpZ
sdFxVlKq9jrIKplsunEPBgPbWE8leeaVg0vTqw2mupoQt3xxH93EdGaOcn6TRTcdxuCFv/xFyMgx
6BoheNTt0EfUa9F3YncFcyZS61gk0vmEiP1cAqQywNSCvJU8IBbxH2LcviiROoX7tvTdv6XdNpCR
sroFYcYyZ3H6ep+dcaVddhbDRCHmChagN82PxrrJrcXhqyi6kcCiXEqCXKY+RF3WT5Ub1ZIAs7QI
+2KXOQNRtPOVdxRcFx0zNIOCT7UWP9JUkTJYSDU+V1RoUJeSTG9eJSzV7RUcR9pgjVQftstAofWA
eAuybbWHIcdInp4rbpTIAAPHiY+1Bfu6XkjojOruFjSgpfyweuvnHcO54tXNxl2JGZ2e5F+DID96
gbSl83w8pY/GiVN/vMbGHfPLNi1Si2VSPWr2qp8QNTs59WCNGN4NxYQAkwNgqyyKsXgijDZ/vC0E
DqSiu5piFQsDWbSYdZTABudiO/05Om3J4jdWMR45xt/RjOfELPdg+7c3nLYnfIwCnPTUyZlKOqIF
4BUlsOjva2l2AILt6zSWgr6Vibk1wVd8LET8MKjm/WQBcBOCOF3aGphu2foZu3Df1ask1S/W9+8J
KIbeaDQA/3UWEn0igb+9/YYIFtpnvyqvdcdhzimOoynNewb/dW2pg3e9llkDN9w9XMbwYmgqa6r/
wH/429PCLZUF5Zhg0MvTdEQ0bvq5bgjlNtmdza56Efq8/TZKzzeKNplJ3eTu13CFlhDdDhD4UDR8
PdL81JeEFNJgcAvR5ayl+z1yNHaa6TIeMPzYQk1yF8h2onzWLvOcPURkQBfI0SD1TLnbmJsPE0kb
Sh/P15aWzYIK5MpPWdwO4wMlKvxXIRD7HP8WZCm1baYpS68ImuhAOgKW273kTsR4EGSX1xo08ycs
yqowiWPK9svNOjg2lFkxcEU4M2yFZB1MhgTJ/0fJmC11xWFRfl0/UFRt8rrld5NV4h4IbFUaP9FI
Ti7vSPushBqcSbzg8RfAokxjByCCT1Ujnr2qkETlwP+4UyDnOWedldmZoM+J9nYGEg8nLykvfEkl
o3uiDqCYRsa8QjVjEO/NlHf2Qd1ZI8/VwMoFGSAM0rqVsMzKvthMCSi8Lr0i/TUjDXnr9nGO2Z0Y
JtztlPsx5wBuyWcqQRCziDzWCD4AmCKKCKEH5ShO0zCNEx1fR7wXBHm4zBu3mRbcCNPV8bMDf0+7
DNCxklhkPAz6CJghnGaEUoaXmX6gETjfQtEpdg+9yQU4SElAn1usJCnTmgSdOfIDvWMeNdn+X76l
4uK6SS78kh3oIKVr4Xt3P6yrGQZiC8X5aunHx57SSMx4vvgKlsmvxDD8DaXDeeWHMm6oahTlpYcV
s2qvPDwo6RTVXrN1RdDWlpg8C7RttgkXcOo/OnWAdgrtIZxERrKPwq70DueblYWn9acdONEMp0Dj
67ZNb5L/cSXOsVIIVU76QpzFgosLDBXoB4qVY3x1flNwm8QxawP9b5QW/tkrr2klchhqGxJj85cD
Ut2A9N7nGaJtDrX1DUzGwWpMKv4+VAVhONnsXQqoFM056fCFHTmClUhaTAD6len0LrQwA+v5OE5r
8cJKH0IFaN6IXfq9ztYJt+cDpO8mleedSatD/cxCvXK/+wE4/aupobgNY4hSMBJEVcCyIkD/Hnwy
YwcmrTJGTtRl5C57g8oFC/AZfKohfs78FkJqPrZVnfzpkCTm6/iZIP/gtbUudY9VWnP1QAmMezQc
47wIsWGihF4LsUBLqzNICpDrXy6qennVDwe3xo9UwYEpT3VVVsb6WgliaIuCK+6sdiLGvWeLNF83
MmD+ttNDPoJ7kOoh1XODMPs+aWJXIFOgr4u32KrbrJpEIJi1QYaqfmwF73pIYF8NR6OmHhfnZSII
7X7ePqFrKL1qn4kuIQ7Sgp/g53hAZww67PCiBLI6QE0U1O4xIl3X1VcNjpsP2F2IHSX0gJMvn/kW
xCxV1QHOU/tbwKYjD1B9DXUNPLX/+9tb+0WGrm/4iaqlPraqjun9lYpfJ6P2mIB35kRq/a+7xLo7
Iv1qkxiJlf5pjmxlvdnAOzql1dhYSiH+g9cs4awC5Rda6wsbIjQroUlCdQC6gO8+AbQDa/E/mkDP
xB3RiaGyzegZH0rZTGNpvjW9Jn17C3izlHsL7N+brgXWhCgjE0ZfVHzrghLCh0Jx+C6GXNLNPt6J
n0b2r+BIB22KNJe8JnlXl9bquWEArgyf2mDgbOfK3url1SalvNp2G9RuMqjZU+Yf1mw02DJGvJlB
ZqouvdRf68uBblJdZWPq6YrDa3fVtN50pypiXvdXL/Nz0Z8tCfCl3X5F5DBxvGqT2lCTi/GwZGhW
llaSOMH0dfBTy0vvzojFl2D4rD6Gl8QqIAC/cWO71IMn04sBpFRCMUUio81ZbiDjQ6lWs72b97OJ
vzn9Syuyryg7o+Jh3wz188qjMsdN818psEW2c2YYuTWY+3fBk3ls5DOUMc0sHkGMQm3LnF+BcUYC
VJ6W1XBn61tPr08t9Uilfgg+qRUjqKVqkh475w22n6nkSayo6QuFof2Ou00BZVcmpsaHinUcC/rH
V4uE+2Az8GB2hP9a747PENYmuN7e3MC5bIkIs+uYntlDJxmUsl00K/Q1GhvXsminzmOsnCjx8V13
TB+SctFm7m3FCwas1HpnBXF+ZRnXBOqEtp70jSIY6yFbQV5gi2nyDK1CWDx/OeGJZPfPJRGZHvCx
Qh0jEhNiC5aDXP8D8liNOutJuRpAeFhuWeMnJsrGDkFsI1ewSIMuZW9aybBV2Ot+ar+zTME/BlAe
Sy5qytMol8KvbneztfWdv3heyEH/8Dsau/8q1IhL0we6gkOAM1FPbSBYZzkiVk9Q+7MUyTisM5mH
Dy6qccgUmoZrHY8mY2mMeAdsxk+r4qiDanLrgADLDDMFU71ixXAexFuRVJjBE/pgTT4dCLDsXe5z
/pcWymooz8x9bucM4teMJSPXUBm24tQg8mIUujV0FalHFTMeARu9GVtIgOFyj4gjMX4zBckfJvR7
kSKn5CT4QmwMfpNArXXbvjWhwPTKiXf/Qg9q9JM55H9lw/9Wjd3zuIKZBTSAh460rJTdLU51Mfr8
2nt3NoXxrYt4ZWzf5UlJifUjYg0vre53h+WdjjWwMXKnk7Opt72cNA2vgc9RFVeLC42IDFuD4FRR
PviRlYaFg2TXhBiosWNHaECIcvUM2+jeKzKaeALygOHbK5zQre+DR9QYlBSctxMyJfoYwTaTboFC
FyRdqUpKlcVdWjb+CXTKbqiExH1I1wI9QJfxkIHYm/884nyt30YNMR+8HHiHZG4NozG+QIRezBSI
yYzh8zRc4vbDa0twjObDvXZWDDo6n3MEPa1tNQapckAu82stgxZetVblLpv/K9GEkYEMxhMn6Tdb
2qzlJu55bInM1P68YIW+FmVsFfkkul0KatieEeKcfEwzFdIGi18xPQTf+9hx2ld8hPx2vxEx5LJh
g/3e0hetJ0d2E2b2oUKbuhi04V2FqXobBUVLdzUqdb3cjYGdeZ3povXkN7QEIDAgaroMuFoDuXBy
RRBE0Qn48q8mjRvJzDUtQK1FDKPqJzZd+FnK5vwfQogM3c2c98NS5kiD4X0xCp1Z1UYpKBQr3BpE
D75lyt5UIVt3yETrtUP9LkqUEkqjMGUo7Zu/FjLWSFZl0B3YGXbI0Po4LF/y/A22vo3iH/5+71CG
NiVZDtUYqoGHO4zVFudWJxYMwvd5eApI6tqp99ZKM7Jd9hNmF+OrF5XsVypJOtsQiFeq8HCjszRJ
87ddizzW16bO6cU2E4jkddM53kVnu0KTNlLnwBpzjZdia3iTwpMTxTalzHkGUDNzLveuMqzqLcAR
XZxmNOYJORYnUKO3RvNMUxQvFNWbVWZ3mmq9zlHgLZf4+VACMT+9NX5K5eSfcLogZJ4cJAjRTQ4+
lfx7RWPzaAYbMEBDutvk1Fr50i8ARlBTUGL2XFGzlU/lmBl/gGOTmmXtReHX4IWm2FOuHtJMFnq+
bqgvb5Y9oUhmSpAtow9ZLdg16/jQcBJF12dys+yjbkozsiNJsA3SsjB5JImNyIjhaNayDQLouSy9
qF3wBuSnyOvAmBo3v0eMXwGqqGTAyvqWNh1pbv+KZd694378JH6LYjKBnQAQVg0sO4cyTkropZRV
xumAdqBfm/mjdAobq9SN2qqV6ylWhnKr9qr8sehe5KHUbIPCNqDkhZt3SY+w8ys7NazHU7jMbHeG
DGzMECmtIo+WXFzOrsG7kJDZ8Ogr0YvVs9BTdkiF7dCPmf8OaByEoHJjkqY8cXpv31xe6l4yxztC
HM12om/Uo2QoQyYNTMgLEIK+/WY41mT2m4fhgEQij5FVmWrBQtXv19eqbXzVRMHILfIvszdRHI2c
z5PHTnhNnqPgWlOg4QiCp89an/qPgQXq2VqSgtpCb+2sk/HoV2QcWoSS+Z6nVdlNKX8ZTQHPihI4
ZXnbSx0I+efaBVb1UA/N4n5zW8FvbB8gHgxiHiyvTyce0XptirCWeQYg/EOnzoPTKBdaRUp+LPgJ
4jlJzTcXKRd8gfw4PwalgxjrxiCvbCBcND3JZVDd85t9w8R3u4CSWvfkUBJkODJXxbSYv9ot8Z1z
ou5UvaXjab3j4qzHyP/3x+agMAvyj7+UeaisOlf5zZI9cCuaWiCV0jupRrrQAeHY3OEbHbNe0326
4x1VpOOOQ3UcfA2gfC1gxF9U3sGmj8aBMiwAGJAQhy7vScCrR2Narv3y32Oy2pHybpKxkjREf86a
V1l19wWVlgypiBnucBkQjavSE/C1ZXc8tAYqU/Qcncax2f4Sb8hGcN9bMpB+Mhcql/LWIO3OhWfk
gGE7QGJTmAULNBEM23o8eb1wAccD97a9WvofhFbMNa9La5mq7vWuQ1wAbyiGVZN1m757SpkwfzpL
k9+5JsZt+VwcXwUlnSw9sgthT4JlJb2+4Q69K1yBOB84ldYPxrcUongxuMz1b957vJ+Bx6rHI27t
H0sE5LN9X85ekUetLyGZaqx14G5khMsdktY/YvX9rwaasaWaCXhWHFAxcqr145TbUXSBpvrAdliR
0Olvv9YACAdcJ91GDx1SJTff4QRnpCrOAWeXAch9mpym5NWlTHWxCZ6mEXQkYsKcBPEudSJqr8fT
tnSNt89HfY0DpYdmVRyCaJqu8MhK7cDKUiiMtLtrQOjEFYMgbK7Ui86KF17j4DKxkpje8Dw4mhmF
vWap+80stN1Qwb99l6kSVHWDDI35ateR4nenNGTcplu40/UsJZp585Jxnzdl5oV1hzc27iE5uUXd
T69chIcfclnStQujTZiJbAS/yv07iRaQENmAPqmC4LhiAICz7R6Zxu6RLlL1JIXzu+X8TC36Ux+D
dNUPznOb2xSBmNKHq0SLmVD4BFwlw/YaRrzzvTpNh2N9iu9wxVxgGoU+VjsloivwqCY/73iSHzMv
/sV/DGqrF8bbqHjbpwFI2yzDUxV5Ymf5oq8zuBX6PfIyBS9LTcKYYbiwL0VWna2dLuaQxBWyFdzk
j+c/UYpxzF5W2L6pqaiWbK3PDDm70M2wXidSZmRiS4wgXM3KCbXL1QsPvpnlFSv2tp/L8+Gs2eru
CbxHRra5fbsR1r4o9bRuugwJPN8y9GeCSxIDUmvnZR8P3BuNWUXbQ+SD78+Dk2TTtJVifQywm0At
EQNPPbXJRvBantsTgdJirF2zMkLgfFadD5xL+uwGq6lEgyjfJ607F3DohFEVKToY5Ekut0kYNt/U
QaKAWCvhD+0q9JIgyfunuhMTM9ei76KE+n9RxdYYD0Qw4x3jDKHrbofGuHWHnPcAAB5I0os6WVwk
BcesOjThVA8dkvmf27hbehLIoUsLNDKEEojKr7nxHxc13WXAhO9oPJThCKu95WpM1uObtV2RCj0t
KoCtQwkuqTc4vTufRUv6Fk0TaPPraYEO+3HqXTAHDmiSQ/gt159rZGHhSW1lzsbjBTYd66kLdcdp
wXYKY+o/y9N3fbKe799Jl2pG2fmCaHHW9vHG8j02KeCnaD5ZjM5a3rzR2A5CC/z6XMJc2TLgBTP9
DkCVVQwXu1offv6k9yXGoOgq/0d8PMvv6m8vHrAPPUc0jzETTNQSw6bCmWHgFNOOqoGd+WQ73xj8
3l50CO3IHDWqRO3OdZzumRnnU0xmAUestB9nynISfgMPj5i0SGbvSF/LVUIBGyjK4moeV7ey3e5R
l/u9pDovSBvzc/S6P4lEijz3HuIXYudZQjK9nmhF5VELnLNEK3kojJ6hinKcYqkFdp6fOLr0zqct
uQFEgtNkSkSXtuFW+g93/42jfgyzOeGPUPWdbF0NJ16h8osg0tz//W5uPY0QbFOnEdk2T1tsCuvd
wYCQrdlnM+MYw/ci7cEAn5dN2eKzWcbREuMSk4CU2THdvrTmOucxFkINm8KWPO1mQpvvieNhK0Ee
Ya/+UPbP4k81HmOYyCTq+gdsmed2+zw7EtBPkddb89Z1K4c/qtjaABshkNoKQJjGeSKAZF9qK4bX
/Ok6c7Yh0SS/FiVkh4V2yBUDU8n/LI6DnyGrtEfqE/ohwrMAa+JY4h+9I9PfdU1kigBA8sCzYgB2
0L31NpYj5ye8l5+Kjr7Qz45mr3adsoBc8aVm7PnQIl34zJ7ttlB0pn36Uhs/Wn/5u8zLwizVXXvz
zSqjHwoNfc2J/JEL7HL1DTzl1hL4ISQWQSkrm7hXEnEQhgcpWeO6l32Vhdr4xyA/p38qvq/v03Ip
lPi5q8ETMevFH8/J8TcM/eWdH+et4nVnKpvhrob64geF+eN+ibtOa9pksiPQ96xKWVB55hENPUpw
c0zS5mvUSdzG54gRI8NSDNeSXvcZZ8diHdQbEGZqv/db612zWGAtsvLwUx43429MFSzxwlS7PSKc
BNJGNs8J9j1kI68zyQzl7qBV0ErJ1qAhxQYK3EdULAXmg+xaEECSxtJxF9DdMt+gEkyaLNA4PKPF
0qYWLI431bLKoA4k0pGjaJYBbsw+pVjiX5ybUy9B42ktZKKF4wgfbFirOmtv/mSK/c7eIGk0JM2O
2g++qAF1u1950FDIj0W5FIGy14Lz2IH+kyA9AD4t0y3gHm7R0WHvgF8qfv6t3JPyudigvxScp3J+
yhVuNdy2eGaJ/El97pTJfGvU2e63JQmIYVB92Tx4fzq/7Zb9y82do/nUnGvKMaKCjwbxEhjclWC4
6XlY25L6O7qcK9QRdJtYdtKHatCHkwPUU9j0F/mLlFWbUidW35J4y5BohTZxmbT657jmSwhvWajH
2O1CvxKDVh9MAER2XoeLJLCUtGFOIjOrrCVSAupTrHG3PX1pxa0AYmgK6zVJ9DdVA7m/gS7dtNIW
UCHRL8xSP4kCG15NZVzXIQGrcT6ZyphgPm7zG/vaHtE9pdel8+7Z6RLaiIhX/B+yot8fmH2RWpif
v6DgM4q82ZbN8CdWmROlSIbfME4X92WNqr9YCqL2TW5ZQ1hb+joLOFuDYW3Fuwgp2zU4kcmD8LyN
T/iChvb22I6/59aUfnaI4FUwN9IHho6W9NCzwsbyDRg1pyw/hUNt2c60W68ZkZEnpKF/TaHTspac
jXCAUIG1Qm3NAg8fmeAK4Cf+Fck1dSPNbLTHTo1GU9nDvk1W0yz/28HcWZLVdpVLSfdK8NtxN06X
A4fKeXOkT5LePpccaMgjGlCCHQYQULcfkCkzT0ic5jxgG9uZK/I9vfHfruSFXbaFmG/G012AHG0C
5LSgllB3emXjKE+x4USGeX2jPUSXC1iaeBc5KSXZIgaGnG37w4V4JvuWn9Af02OJkmDmvK3jfp/+
N3CAS8r6+bNajpCm+498sH+2O8At/5Axl75gMD18t1amlHK/hMFpPkfLjDg8FQrPwvW8fljwnr1F
G32gbtBCmqV5wfcaVzhJ2UMdLM8R2XXCeLlwOh/qPJHIsLRINGcuBGwo9EC2EC4nKsxLB54/Indy
Wyez3dfYdIZy341sXXGuxFeBFrfcwi0LUnB8m9Bhv2TLKAKcTrT5i+JHAGSdRAOH8lnumURQvwzB
cOOt90Xa/otBtMNCak4hgJBtaifM86jXTGCi9ObqfoYeEtUTjIsGo41QpZwInd39/TZJ/EgR+xda
5ShyT9aQGOaYRvNUF0vFfuFt9TZS93fhy1LbkLhKOHFOtXIUBeOAQKBbg1On/2ApRbHBCS9YGnKl
G7XNWS68eVd7tSq9S4eIk0bk10AUBF3cujwfdP4MIPmiLlVtYFlUU2QN4UOi2qNU9492ZlASA81/
zkr9XNZ1h3ow8aSbpafOBBKlJJgm339QaVXxpZ4Gz0v3Qto2PA9cjUxwztCj6YhO7ngOe6IWV58I
sZaceEH5SiglmTBbJGlZ3LlDSvMLQwiEsIWXtf5buStH6CEv8xUt5PvFQyQdPo3e0F1uT0Av3sy6
4fW7jhzQKUG8cCns9Jy1CBJvx/8moqvwMMIHKfHDTH7s86Iny/JJKPENPhtp6+cUP0ETkc7N7cIz
o8ljXaeNzM3qpGERuwPTRPq2gtrwdwT1jBEGYEvrzbuXUqih3iXiDhZR288DHXYqUQZO1c3ziF+q
vTO+WfpsUth7lKfZJvLuI+bdkLYB0aKt26JlQY4Of9pEdtnS4HcKn2fmrVz38EC/a59iYJDwL05Z
XlkGOb0VUGA3H/7un9Z/YpgxUgH0l2ub/EI0PVu7lnpAxybCqgnFDA96igJecUVIslL5uQ5pCAdl
zsfJ3XiW8yt3/ijWVzD9o/xcQDK8U2PTxrjZzxpnEGjPenkQkEScvp0HgSnNL2qdZxZxydmSe0fg
HZC+Ct62R05NjdafQ+0EH3sNIBKvgok93kX3ceXnmiBNpyYHp4WnCEq7jyXjCdiLVImAngeeRM43
HPAfbTgSCrG6Tln6V3x/KgHhdXvACKE8DbrJkxzdKTA5FN5Y3hUMXmW77/oLYJyU1arI8jb5Degp
DD45JSJi8LBvxgLI1wGH+fZ19nhC3iR/abr0QMkQKXvBxqNzP543kNjNFRI/dEzyBrkaN0I7Fes+
zg5w1qfobeAQdUGELZww/wj+O2wuFIpWczDmyeNwqI/bEh0rIS2T3P2JtPo/N8NArDN3lym/hJP9
82WbszNjyRm+RXt+KKqdJLS3CbmzXcsvP3Mm3/+WFlb1maGN8bBKL5WEZN1N2ERKba1557tCXVVS
7h9qiB1IGu1xdpR3uXR8PgHsYiY4M7/Zv7iVbkIRMHKSVLTdXQuFGXjBCJETvHVUxyLAkZYVpUPF
UM37nmTyZbR/WgDyqRRr0Tjm7b8TMwkiV0QSeM84Y7W1GiPC13+W8w1OLvjtNRVe8CTaIp7wcRSs
Wbm7Gqs9HaL60EtJW6TLQ65pocUGvFnXmMyDBVfj97rbVXRrj3a44EeKL0N5BEDcnvjC7WNBSUCf
yhMvPi+NW8q8nnLgYglE9gtGtcEun75OfpjgWzdBoYjxM1NTr8EIJzRWHqgbkuzvnCi1yT25G5Vd
v2Xa0nFUFcmeRm6m96KXtUSCgXCMnKnP1o2qS0buJ5gLSe976BeMdZV4J9BMLeTfhF6/ekzrviCr
lH5Td+rIDZ442QdmT+3RX0edLysncpupB/wGUvRA5VMD14LtwXxSq7ChIL6cdgGQhdo/Ody9a102
0bAfhp0zpWYrUCrIlWttydFGtTFNLR4FBgImZLxPbVD11B2tFhPv9mr5O1REdq9Ti72Nv5BghXNm
mquB3YFvAiXtRTURUW8jD5VFk4HCgYLyyFfQs98nkUingiPpz9lvzO7Zu+uiV21b59kJ6oahCL1Z
6SPDSXAbHE1OhzLW++c3+zJkONWho/99ZcYRElDmUvJScfejZ/nwsDQUyzFLnvPJK1n/kmNaxKpH
8exj4DpThx4QN0785O/Ucdnf6oIqK1CzpI+1sfU51KIUJWiGUY44a2kROgdN5wYrnU+2ddPS7KFI
r7Qw5OgsQWOFhXwjKQ4/x5Lm4IxPIxN60/ro36bkvOhIwzClwcel51s+W+xYn6UOa5Kgz9Rh9KNL
mau861EzC9qF4uRMXvA96k6qAn+iqv2MwQ5Shz61hN46cGn3QhNnhi2hruu0o1nhz0Bzseyj3CXr
IXUbL4Vig5+6yrfVqWEqEYBWEVUgDqOWEUsNRjUldGs3B621jCp68NzsiYb3PRTe/HyFcuxG5Q47
R9oafHhrGIecmyOz5Glx16QiqQiPzdCmeZ2QAA1+O6vDVBm0Fj8n1OeI12TGg5BN4i1PBVEj+oEp
l3wPJGnWKlkT2EE9ZGxAxzlE1XvMrZSPPejKsuWAakT9FOujfbf3z9wjJfMW6h5jr8RmNnNOGQ4N
GBr0phKAjzQ1gYfOhRTZvOajZh2tNlKHH6E87Wx7s4+reMn79RCYmIoWQNNE/JQIJHduYdAUovob
cZ7dOldDSLFnA2iX7pTZ2GXc9iiNLy4Q8Z8gvwqLuSOycKxeVFWAf5sE60+TyiRXofo1IXS+XU5u
jQ+0PzMZEuEd+2dlzpFJ3F7vwtKjKsvSmZLm9dFfxknlWMW8T5zdfUodlBFAyKxEhFev3l9kMhhd
knJNJohgnJMSeLHOEDbC9PMT69omQTSOYLr5GDhChxrdVDEBNOG5t9bcy0rX5D3augzBzyL++NYb
0sXpZH81GeRr2lG6JDuMlohwHDO+JDiJhAMu3VMZyp7WQzvmYMoTiVAKiZ7gB2/HxSBX7LNEPv1i
wJhoWx9ADprYvL344aimr0Jv1ch8qpa2Sds1RZ92pOfz89KBqcIm4cGe9lXyGvKzc49SmgM0wx7p
GX4egHN/5UrOMo5bdW9nPe5eAeNolVnT9gt3qNy34B5VkVuuUwsmPtj2l0bOUvFHlluskFiOwXxf
vagbqkAhkJedjPS3jKHJ+6rlNe/ZETODsvXxsZbpnex0RB9zu/XqKmonMtbadz4KyJDCqFhShg3z
50OpWbqLIOe2eox9EF5NV+KCj317gkAnMZdgxQ5AtEXiQPZ8zD+DFesSc/yXtLa7cEJWV5GLU8k6
frRSKbOV0VBR+oWed3OQBMghuwThK3hnhuEGaVanMgHtn8FPYwyI0RqOouvyxxi77of/xEGfNdj0
JjNTJkMyTxc8afesWlfvCSThFOmY9x4Uw7oyJerZDS2FZksltQE3z8PDeW35L3Sp5wW4TQW8Pgvh
JcCBfdPtewf+SbK8BkxZOaSbaeiDUv9U4vvhqxgKoDRe+sq4PwdvIvCSAHGsdv+zUKlNSBSJYAMQ
OOSrxvoOcmqUHJR+muMijqjMg8KVqTrWTOHsDHWrvHTIElMLKa9gBM7pPBcrcfwrjYQsir+iHbLv
grKBjnBzcdLJNH3XxCAF0JUorIRTppzS2TP2LHmTmJ+T4yzA3DbOdVCtzZ2jZBdWNXSEC1GG9YSm
/QxXDJj+5HdEGYQeWI7OOr4pAhz5uoGWzrID4ofck5yDF0DAyx0Rz99X9sylNQlGKh1N4hAGgb21
Q0sRznJXrbUvZOcsMerbuoBUd24VnXqKj5cLtIeoHUIl+0StZ6rcsgSSsnj6lbvI2fr7U5HiW9Rz
tHcdZEKFJqlq/irLNdO56Ve+aJHfwUq9S+eS8AVpmlWyr7LuuflrDVioP+BfLFpTlwBLiZwBJfVc
UDLKQ6w6Ol5hGyqSyl0qFdhGGxBiWTtoO+obJTpJ27Pdazel+OWqn7qL+rNvm59V+ucaOb9BEwe9
t2+CsePrlxbc+lfyDRNZirNAtLaAR0SGaeoewS847WuzWfmfWv4d64nSXm0XEiAo90SchJ40PONI
s2/xmurGrDaIcuUTRLAOz9LRBLc++JnHq7iswZb5oJdYPigo/WnoX4ZxeW4msfvlrlUvqZGxwXHc
2LIM6WtGUxSorrpdMpQyt2NKpGv+Qi8masR6KUjtoeP08iv5HMN04GB1tbVqWpjGvximyFPyNWqY
w+/0hg7RZfbXbi+moVsaky/Z7b1xaeQ3VY/boKl+6O4Nne9uaVhpZLjxUzbzeTd/c4Az93ZOZWTE
mD95X018ONSYwW1XDvuxPSdrmQH6QOE4OBp4oeA0MK2kXR3xbcNRrHgomII3HW+GxjnknSLf+fN1
9z7Fc2nAFh+qCs5mE0ECSfAthX2FdZaSSPcyVhUsr8sSiyTbMygd0PlnukcGvcj04hrYRN0zSf67
7X+EtTAUyUH6UV84Wi2SNw8sSP1gdkxgVc+dRDYTkUYtH+J7D1nB64TarW4y7BF8TMbhCs/Gka57
fUvF88EXW8+vAaSAMcz+a3zoPBHriRfmKWQfGP1ckNCtvZhphLamf9IIFl37fSIN+YGY4x7Hogp8
qjxmmScRke1/G3xDRHX/d7Uu091FBpaZRpCRHvbekVKNPPBlz9/HUamfmuFiiNn2A/5Lcs9kKjbs
YoXT7pjj2cTTEe7OVmrhQJWNVQrUgyY9cFtVsUAPove8wTWSk8GHwRT33tKDCMKYnQHajzAa8cPd
TyPBBT5QDz06YjIN5JjRHLjABrzW8GX/44y0aZyqIfwRzWR52tWO6oueRH11K7ABb3ofmEhSmaSF
ouUBVbmvg/gmGtd1VCwBbKF2c16YdFUkuyt7fpo6nfsIURwOuaR5m27rdYlkRrPpNyvWWx9YSQPv
wOJHokIkRDVTVdg0U4Na0bgQekTdDUj08rLHiMVoR4z/MAoMNGXtKKSChT0HLJh5ZPetLgtIIc8h
EhD/4DFQOp7g1syhDXRIb8di2oof0InhbEPTSLYY2IVH5F7OOOgAifyQQPYTPpjQsg3HPBWMg0Ls
Fu1BrZwpiCvh2wMQONdThUL5XluGOy/9zg/3zJcV0MrVdB/jTdsGKmxg+lGCJ4GbXPYEcuywx/2r
EFkh83NUhA9hbozDRSU7c+1ptXQC7ik3VhERz6n1xTmAWcKifBT27P5n3XlOq0LL8Kvi4JpbDe2J
o5DPcZVZ2yetGkDqPqdViE3wtjpBQNiytQUUKlVvhDk1v7hBBzUQOGKbHcggKusw6vgzlmvyuIzY
hnk3O6JVY/FTTGmaySrFwPoUbuKkJwH1pcUf99LTCJRCEuCgagRcCjdTaer0Sgr+D8sJr7LFttel
dfw510jUX/XDCFElzPq2ytN6Pw7n/RuWSlm8/e6vfJUOc5P/6OR5Z+JwtCOXe4APqQLjuz63ic8c
TSLoyypwsSNbj6FtYsxQlzP2sK+WwPKw6r1en2vWH5ZdVOkFJDt+cHRQtpXOC1fVoPNSAHhzzzgZ
KrKLtbdh+nV+psCVwwIVgle8gGIYvCiTcu4j3SsJYNEy8Sk8ezwUmxKwGE7y51M5zA+DtKuKR2Gl
qky3KGlbCaiQvmQlyOUblI9iD1GnIbDd32X9hR5VJtA57zWUj0Ji0++BX+LAwDreElmnBUpZq1SZ
/hbo9lwvjvN2Wg+PpigHPjTi3h5/1Ej4IDGQWueTz/R/f5AjxU6H23aoIheqdZHndFu+A0ni10BW
U0poTBXfTqkeBSCE8Lpw01cfaCOUjVblIBlgZYGb5cr86Ac51Eea9kZMlUdk791a60k4lZIhcpvq
/l+Hqo7XnfHl8QoN0flnrCyoFNVktHq6VWjvaq1DBoZUMPoL17gGexGH+WKzB7DQe63zJpSkHI71
ZT1HSSH/hQaQZ6DWuONrzEb5HJOp9wgaZo07TtKj/pJBJklN9XkiFP+5ySA+6OIV1H2O6Rwv09Rb
DeJa1zsp3AKSE5hmmw2JvbLD5lv0bDek2ztDu68zpprLF6+yqB3+jeX0bvjawNx/wL/nXHtJWOj8
lTNPH9NmFaIgszfOcioN6XF+DMqaUqe719I7+wM2Ujc/LsxkJAgT0jyfe/3UzApJnuV04k06Gx95
7eoEDIxu6TbCV/YN73tImBnMmeRll/69Vr1YuT3T7HIKQt+EAyc5WV9Gub7dYUKYJVktoqBIk+Rw
HxUxlBILGU4vnbeLTj0Cw4n9cTf0jl3E92aW6MS7kLCvNU9GMCa/PlVt2p54oYKDGVb4cW8fAx3o
pVtjcVaY+6/q/cl2vlWFl40VgNSGgiyCFLlTamxc+tFextvOGgUP6lXOSSs76Kyk2SaA2zwP2xz7
9sk7Ad+toNUlRpAK8aZzHdHXeNDS3R5mjQ17EykQGKWfm+0Fx8FXfbLnCcS6bI5nbl+tw1uCiJor
lg1rqvrTD8qvU5SN8RBTK5Eq8rDMhBSlN/ncDahztNbOKKdnYgsWP2N3X2l+E8F9VIWB4IVJxkgc
Zh9W+Tx2e9Gzslvqxb9ArOTdblmxIvMZ7+wtRGjT2L1yJ97DcLqJRMcpKiraH/BAfmLh09L0fpAM
7iLoXyrVDFNNzBVxbGzaCCymyU6y5IVuPOpRjVqTli4WCRKH/oui7hs3nEinZtguib0Y11arUcj7
DWQaxy0fk0XHxxCGHlhQCDWnngUYdWXsSAJ2BAXK/oyF9nrg9WwHG9QSKI6FEcHNEIr0ttioOjcO
RB4Y98xSh5f2e6MkTRgF9QdrZSPu9L9To9DjhHJCcqbJw+7mJlkkayaTNELfzaHUkhzWkp5MS/pC
TMCasJ7ZYlxp6zG1C3luhQYoY5IruDN8HgsJayudCNqC47mB1iI/Chb7BjChXJSy3l78ujIfOIdH
cpY3io+FDiTSzv/U/AiHAq1Ldpye+WBlr6aiy6WWrUM4ar+ptCDzaGX+0Q8uXjnkfebln9Rhl0Ab
VBm/Vf5T/AX3XHjl7XoQia2JzCSjHWeUZnVVGGgpgJHxhrPO/yGdKjwQjVX+gje8AuYoBfapgvzA
eAmCiIqTYCKA5Z8usGCSW3RrO+SsHZ11ooZq214h8FYUTMNIohujggcaBAIOpGL1jHMuA0JvEk9g
9+RduU0nxaPZWgEnVrIdvkZqB9NREdztoqkYwoPnv3E+hxeubZIpyYxoWKdhXgmy++cJIcRhZuG8
82tLfRa2Sz3/7aBvkc/X+RUfn59vBKLMryg/kvp/+0lJIwKXN9ny0dEvXj5WeAxdUV3bcp4Jz53b
Gavg+2UGFtRbCTo016ddTrU7Y7p6zqLKTslMtD3on12zFJ07UrCSDyN2H2U6Of4fZg3ECehY4pVu
H3YEa4HV9gezXstzoPmN1o2oE1xv9SS/3vgfUifVdgsYSJ+Mon4v+xSAimbKPSmjfdfiMwiEMJwP
Gi2nTShD0ivG8ns6EKDRl/sV72l7xJmHLDyXPV55J8w4gHjxC5WUcgLFAC0jpVj5OhAWTOc/u01l
hV9Z5Ao58XatvYFVkqrl+QcNg117gLQymbrW8mJk2i4p9pkkHcxZfvoQdGvo607iXdsWXURBlHVE
/5MDWOI9I+qJJlDgfvCzF8XSfOOl/XagSvSWiJdCnRg2FkdmoyQspx57npgtA2LTBMtMGy67HiTl
Yl0D+duEELIzHtyl4kZ1AyFNWt9ptmXpRF27NPBFxw8VbWN+cS9SruHuliXTtwi0hBSFjE7odsey
gu9jNpXH9VFqa3zyVhaCXfnk102QiaEYgyLtnzj4UCOheerKsPYxgPKkB1x28aeEA40clrAWTKhQ
lcDwOMB1WRqwIVi+RnypNEwqk6Dbo23tX8GLfCWoTYSVnrryZt1NzQCNuC+ac/I3Iv8BY0B4dxRn
3d0qSFDEMZr+sFZ2nEYrfKM6qwFFnyoLiqiaoQHUc94EjjFPAAYC1U4oAYWea9UXDjtgJWqnwsnj
M1JyrC9eb2p9g7z6gKrPzJLDKpg5Wgg9FQ6+CmRnNB5ArNNNlh6mIsC2Ly6JHyHMobuqJUGT9Kyk
TfjwR8wKnBZD1XVioBJJeXs1ZqCyYYitOo8l97A2DnXeCs55Vdsil/02f4UFyOKhBj+sfKINmTz+
cZidHKiHmWSPTzYQpnAj6TOMBxaq9DikbR+wgDoxExqMn8NPKSY+QW2bADOnzTaV1T1X4ckIrxvC
RrDGOEJ08WNqf7WQ91LLeic1uNfZ4L5x2i8ItYt7+06OSEjsVkZe24XL7HWBnmhvP8xI0RkyGpDN
EElx1jCXsUgMrfUYws77pYJYXBRvCruAIBmd48LY+KNOB8Ld9ypagrFIRKD2Yb3ZFmYLs9BekkCC
sONs0PE9WpShKsP2L913mXgQ4wDB4Znu1J094NFQoXXJDNB+5cq8dbqjuAXzzS28AGKb9YhCjEjE
dCJQ1JHmh/Cckrz6630TDCqzX2cALbCytXXEzaY4VO86DinPdj8GDMfXrCUBL0ZxqJetvF2HpRE1
bRr6xFFkmzvjWVWv4xuDtPcyEyOwLGd+tkvrzaKT953y3dpKwKGgAjfVnQCJpEfMYnoXiKeVD9Hp
E9iAtfkhNDWbAEJgd+4oqb1FJBHTK4CDi2s1SU9+Hjrb4HsGqmYJIk/bb6sjy8cHSSYQSsAr2L1O
6C1St0f37rADJvln+0rxhn65scheKpSR/ly2EaOnjd5rzLKnKdDkRFdUdg3wgp+qvjCwNkEw2JC4
db+pUfK8v5ZUhsgMAxb0lBfXuXtXLqW+YHIFyjO8u+yqx9w6FKcP1vEeyYFa/9k89mP4YEPKKCxp
5yvzrOisdVVSwStdMv2agqYPXjXDlE3rv2n/gqFGqsZAfXH4mtzOtQfBAq3JU/5Y8s0MQorgwqY/
xwF42/fJFWO6+PrOwGeRMWqCZwIBDiTyH/7Hl7kDpt02j+8E92/jJadu1ewdNTegHK3htKcLBdCW
S8FcfFc9KNpRn8vGqUvj9iHWj32ydveNeaM7R/HkrZOe0GM9EWmWvNS/KNqACFhg0pGTTSmDZ3F2
+neRtW3JSYmwOgwN4FpSkYYZHwZ4dFxnKifwBAUQ7/fbRu+LgrL2G0RSXIzPqqjotFVpgmX0MmLP
xl4xLiYRdtjW6et1xPovcMVtUc/cJ662N5OjX/8uWa/PA3tfPidY8QAKxV3dE/gYeHw1bUDFS8oV
k0Rnh+1s+4vEHnDmnoS/uBSxCrBYf4UKk5M7e7VMqTVYUj7bReL1s/OZyuMKmK+ffRO6VLQtI4hP
pKPm/72PVo87TD73i3laFbW72WrKcXHMPJNnbYMfrOBRfFLcuuWm9XYfwvZz9MSi/osq51QY3Vlu
RoRxgYxhskUobVZfI2TCOq9O2NKsAoo7zJc5Rd++4NKMkx8cIa+cHAeAvp2MKFqVwQz6RdjksCUE
4sVoIhsQAGiwSadKtFV35pYwdxLncDBQNrl+x6vD4UcI2ngsdp4+eWUixc7NFVDbV/3g5ORRLLs2
aUDvSFCsb0M1TUI/nv0Ln+J4EpQ0av12gjweZ2by60D0oA3VaWAnilL1pqOiDI21gpBZwc3C2Vdz
Uv+E/9fsBynzXeg72m7VgbH6PqtsMfoTQTV/OwewiAlT51gkAr3WwypAAzqb/FlMlJir2P6+ZGU7
olNXaTjVCjOe/IzhxvG41IoHFnfQC1EA+OfhoppOjz9+VhoJ9mVqxS/5MO1tP6IX+zhRH4BNvNWE
paZHDItMOQuVqfcWsMowc7bW042jSs2IyanYouZEAgIvJ8WWo8s+e5sKlMxwoCtNYFEaoLfJY2pV
Plu+kfsoG9cCUqOWjNZ+kxx/zgFO7BKq3uFBPpIQ3n63cQAkd2DTMJj1Abf0AKp7/Dq+mKeA0iWJ
hLmPRQ8n4PsA0N+4Y3YvGanD28NDFHJ2T8MEWiwW8YAlcdpyczs6ZsxSFHc7I4OqQn+N5Wo/9oQN
reEG8xXRMiSog/Icr1BFzNfb6wuOY1fN7vd8T/rJSKfQN+0JJfJzjwRvxmrc2awqJzBJCDALaNet
WELGJC7SyBLNbCAeqtXVnQPRNUtsk4q872ZskTprkR3B4L28Tii1KmebiK5K4aFaLpz3PO7gQEtI
4qeMSm2vqedD029DTzYv6TuuVTVQkFTAyvG/Tl3sfpzKlOPPHUTucr9OXGMV9DDquSQJxRmMnNoa
zdsKjHT9PIJ2CJkWZh++sRL+e+HEoR6eTth2JxflZb7PNRhyVzBteJu8VvvjGLyMQ2BNCnDEKSbE
mTiaqd7JTgIfF0GpolltnQNQ5wH83u5dtGirIsnTBuTUkRQDzT/EKJaDxhIG1kB0VNhMy+YJkcU8
lEJKggRpvTr91LfIOqBUNFMXR5mp1LgK39eJ8SbMJ3wyf5WX+qzVGphNWqaw9+JlvDx/AKkCYJy0
533V1aIHLbgik16mcox1MhPlyzK4WXLnKLHM/90aBlNVj3z+93iH4vTpimCOG/5twF/lOHgRgTWg
4AJCUZAa02Y3DECrG17ma6mGVkcIxHCqbInYFoTSsthF0Y1BQdxFEMXjawN88eOmL8aHwr5TikfR
TRUHIRraV/ngwkKWFgyWuQQZWpJCMBPAprbi701AxDwDVtENoWr04xf2jZ5SMVoARwZNXAgxvdCo
OXANxhA5IGyLrKpczJYgIm5xkOTD01aVG/G+4lhh8lGUxftqZ58nYT6rtLouFDyoTdUmRTDg8h30
/D6Xrf9OPt2bqz/MlMjFdhsX0hqhMp6CziCREwqbxfvWyQSzV6NZ8eNbJ5AUr3z2gskC0rWbCQ62
bD8CTi0ZPxBeGos0cPFEzc+s1CJQo8XQas8L8ue8o9/eOEREzfjDZXtQzicL6vGPCTljQzbqRgGI
9CDxFtt9H3Lfgiz2ibSJOcNR+Kvlr3AsJGdvxPmZK4LCK+HNNMx2L0JNh7c7/ZRqwA4EbhXUjq+p
m/M870cg4cEwYuGr938TYiD/c0GiiMEJRVWbw2vXR9DC4vfw1ZXD/BS3XLTdCt9MX8JdzOKW0lWW
MxnFwxrocLUfKoO4S5d8ifc0VYt0bViH/KXdFN8X39gummTWsQs/5s8yffhpOVim6S6BNL8dUyd6
8FbIiD+qrtV7z2oUi7g5b7OOiOZxX9FBBur42VNmBLiTkKb0l9Q4ZsZhRVzHjBxOZB52UplpI0ex
/xrNIL7gKDd/coasQnozrjOWTpP7cbZG+LjBEdIn20VT7NEPgeMTyJ7ZEdmuZ/kO0jy6cXn9jbYK
pFpPEMUzDciUuT+D/N8j5qLISwKIWXjZcAbc/A8e0wiYT26sOtmDGRFu81b0934+qK5gGWUZsDtF
sPt9gZY1YQ40kZgBS6txuAvKPbkai+1IQ/SRB1c8ejLL9tkc35H1nbAocLVUQBJiUteQmMTWCe2j
tZgeIfs/a6fbVC0tKaYr1XFMyNhS7rHP5eCUS/pYNK0m06r74IOyyEkRjrcKSyb+mtZ+Q9bZbFlY
XXhasZ7S5OZSdOtmRs/eKPtjXRatdT6cmh7Bf6vN8GeC+ILhMcjQXqoPOUA+2AxFwFWMY1v29i5w
dcDKPtfRmrlxr1HaSbMeRwMwC2XT9k2ytcehIlYJJoCVGfJZhYO06HZeIhOx2Bc8gbL/9jNLJLPv
tGTgjuhmW5A6tx44fOXVoyZ4IHGYT+TlZOJCkZoAYlBdlrrLnAXv4//nXtZ2qjTanwNoIJztYCpj
rTdfvMg+THjdeAV+m2Wq6+y1zekJB2/ZbWcjVPgighpiRN2dpeIiqNsP3nRmARpP+TLba9UEHg5s
melmaaNTHAdUM5ekglEXCXm194slmh2/yON2edTBM/AgjW42c9WiLGUWnmRXj+FyOaB3c+K2AdVc
dxL8KAt0dF/BkO6qxJxujbLJuMf2dbZ5PscmbtAPvTGq2VfYh59QSa9SiDRiqO4gOsP3v2feTad/
eMRYHInWF0ehQzKOwkTscDvSxDaFp5Li7ExzYsCvQ5bLK0lAVm+v1jBXN0Y70HP5eZKR1nYoyC88
t/qahMj/vVoCj18oWbhgvyNmrOUTb9ttra0zhmUkTsW39fxWTCb77OOEmbT7j0pBvtb7OsRov5vT
PvcoqMdlmcjIEr+t6xjBDAV5Bp7iNgzCe7rfIbnfDo0CMPNT+FxLOOUp3HRiG7kIWnbTBbBFKHDa
4EE2THVccFD6lOpTd0LJEY7TjcEAOOSfg6TRuN/9/XSfn5piyYwYmFCoH6GxotLRkZgv+R1Pb4UO
CT+NzMFhgC97kXmVpBKCMq9IcklymbjJPOS5atobsgQJpumrXHUVMaz6koS12aEvspVcAsoqtaiT
044fzAuYxh2jyasVd/Bjzu+Tn7q9fFev+hdvRnBknEHEuMW0APIL/DfTxdg+H9Savsj+sOjHUcr1
n4zQIcP9U4cij8tN6SHnSc3X7WPaZgJtR66luw86hGlg9SaSDyOZ5lWSOC+eWR4A83Jjrgvxmhm3
cTA+hdhwTDZjg6HalTjsJbshEAlsXnDywH+GBde5zNaE55QeukbFlKcCgrL+f07GBoXqr33msAFl
pFuztGIGog9bP3ZPjfAG02swVuxVifU/plNbit63u0noNx8HI8JnsShfL/Pxq7dRdvWF95681Mqi
h8xBrbFcM3ZzPu2dGBT1QQUzEZlkm8N0KFgp5C/yeWYybLvD8ExBXnNz06Yo+EaxbtGZhmpoNe1I
JVJGqA/ao3YRbFziODmYshq8j840Ybc2/leS0KR4yoq4UM+38LSSt7O6CXucIt4P9spYGUqI/UAI
lf2YxZkDdoI4MB1FdMj1a8fUyFB9kgyYYZVQkK+8vmd9RufZGnFpGni7LlXMD8SsV7Sdcyzwhn5m
ZRZNh9K+ZQZq1KCs/mK8vQjl6Yz/wSkCwA88bGcKDVF1OQpegEDD3vPX7CwNw25oJabDBilHIHUl
rGcY/2FlIIEirh8thrJ7ShTHaCWCvYotkhoSGZC2W5zMFC2hBlJ5RUtQUdWJaLKL5G+RcDr9kTmt
G2pBhyCVUVAz9eCGGK3Vl8HSX+83Za9NhqMIUygLub+3i0bzV3pwRzVPcWAaOTnQ2l81iiqkevmU
Kq7I+h6Jwzuq064DEUpRjcgB0dKhaPd517KdThKcF24oSWWH2Hq9fX0dQmKiI3qDZKWEvOPsE5KZ
hgWIVYSvwCMwXkxU3AP/zlxgLUy9k11OzmwPw5+cX1Lhxq3kKyQoPbJtiU1cZzTPjJKJtiwnQBct
6+6zc9q0of6mN/4mlvYo9q2Rzn21pCS2ViwCDu8ANe+sR326zycQb+iEeemEKs1UvW4h4P7h74LD
e0V600RrhGHgWNFr1f/mAcmQtB9nH4+PAVjMrmvsm9BX89HCkv+kxmwVUTpTcgNFqSY31cN6/0Du
cGi6QD2Ci/lzeRWB1KOYZ0iUKxJXv+anliToZivFK9c13/SlVQH54GdgEvDbRdphrxH2XHJS2/qV
lr0RtcQcYlF4FevNryh6RWyLByVvjRPJUZ9ZTjFPLd2TaGSzunWPw0FaEcJY0VRcslVdOGpjXbJ8
lyQARtCf6BcoaPEzCZmc+PJkDMIp/LIxVm2k5iYekrKsamAocrpGZLLHcGwX5U6n194WbY7NXeJR
/3EPFkFtlTxJcdkK2Bmn3rTFI8Q6wXrIMLcygzJaky8XcvQrc4KHqk8E9aj5S4eX+Xf4H93ZZuYk
w6ZfT9wA+OeFg9KXudpVSAcHG/YuV1u0LFZ+b/asmfg6w5Z+WDE9pydd44ARdrWjPe8SMOoLVmHi
Po3YAu6qm2P+JXtJ3TwXEGovmKidyaP/xhNGlfM7Y+IekwlDf8eRCoOIHYh7DIUMwgNdPN/bE6Er
lsqrqWDZkpSbHmGWkSFmG1jWAzBEPQ4+4UZyFhj3SNuVDjXoT7YOJNIWwlozjAPpeqd3yAO20kUW
92Zuj9XoTjuyN/X1kDECOAkqbWkaFV4z29pzwIM2MWkmHCSwsp2Po/1WmFZmXKwgwqJKBIBk7Wi7
9hPMoIUDISe8XjpgDPVaieMZDFc8HOtQB9G4vUWkzvmFdaMHa0Vi762868kCFQN+tvs1rYJ08pGI
v1PqGxJg2thRwL8SiZHs+sBAIo0K3Xc59DnBkXBkIts3m6FJJO7zHxAkD4sesjA8FKmj02q0bl6X
aGpF93UMAjYBM2QPVaZ9usrFgXXwo3HFVIIP2ExJhHPd0iZcxauedzSGWxZO99AW4lN2PnyGaavr
XzrgEfvd3FIy1B+lJ3JSO2Rbq3usMqSEB5PRLbaW5tNAk+VRCG5uq2f/uB/4EeQfZe488obDJdyr
b1Ec9zbdoI2BpKbs7/scWWxWHfcJRRhv3c9XDixrUAbO7WZ9wfEPLOmXhMxZugJoLW+Ws4CNY4U3
bpYSgWfktI6jk61xgXkaHwYxt5qLkc3PwgyCxMySsc6KQ4lV5ojIcG/erCpEdA0RDNgeF7FSbBpC
96xdUNdhsBnjgtC93YMAugvHaF8EhbbhI5LYv/wBEdQV2an7NJPf0bvmwDlqJSRyHgwVpECHIaeq
KOfk/ikaXSPMDbBWT7kPpXNxUvjGRbw1T9waRjG4h74lLaz1XOb3OuBiiFHDATq+vks5OiXCCeyp
pdNVthz4RkxCCxqUKXx2eeDyQQJW6cgnCP3Bnk71HCFY1+mS8GWhujEW6NI4HWog1/N8MXLCMSBw
Iy5CRuM52zTFo1XxVBwsZQcgtV8q5LqNkDR8dmJQGV/fgU4O9UTMvy9UDt43XIHOxqfIk1eR5cyu
Cs8mLHkYVgqWZv+PryOmrPny+HnTL6CeNtLeOYqq5E9/rWSOlerINOpveihaXaXX1FPg38zFTjS/
J8uzB8Lve/7hUPL9LrovTkq0Qx/Rrc4dV0AwKcjjULx2eV4e/6/tPsi8F8pByMSw8Ek4b9LaLPpi
hTLk0RjIJMWpuCEk+st1sNjPoNn6mHuaXXuykKrU4JikZULiOGfJfpdfNZrCbw6H02U2T/OyJSrU
ZopCj2cC/UasBzaJ1T30DU21YljxmW8LSIrw3KL2Me9piG01n4HyVMKifSRTNT37wXQcLpeQObG6
v0DjDdjyrk/gNAosBNkDICh2JQR7im9hogzVnsw2U4u5ElgApUyTgGOX9OFnptLWy+G0F1iW/cQ/
g6Iar3n/+0lXj9JNc0dtcP7uN5HaHA/HaaArrgz3xP8S8HtQb040ksMQ6heUc4jdWWV0AS5VjdVI
L0jinMiAERuQ53757ojFdnr3txO4ZrftFoh3lB1iV02XnFV+Z26E053g2JkDplDl/BaSGXSuWq+7
ijtXvUMKb7BCsUVokecc7hzJfTktPi03IpJbv9rKICcNOcIcuhZMD64N/i901ZbloUHb/kYnA6ry
iFGrogyVM9JZI9J0J3BGx8K/DyHyldD4cFXz4Ryqx37UioPVG1JruVZ69GkXAWHeZlbU7rXBtnCn
OsPjIVlcEiTfir7JJKa2s0TC14Coe6227uTfEvt8ZhulXS9PWPuGC6HWu287+4nBTDsHPe3bSSkM
pfR7b38TeZZr9jCOU6XZ9lGT9BT3mE9B4tSCLCAbObUvzH2+AzNqLThZUypj0imxtopEw4oZiDZS
Ri242T5Y9UL4nFZbGM21pRmGWu6P0o6H0nwx3umWsfkpXbBm75yJacLVw/fl1hLTC754UAs9CXT2
gDlYhbpxkHUShonC5CKzV6ArXgMIksilXj8YPZsHOR5Xq7AkdQ7k1ihUgD7WG4yU/Y2Wyj50K3S/
vbMkdu3nyyAxJIywRuVNrFasRloJEOuCdJ4wpJ1Ce4MaX0W3Z3um0wlJA9e8zoqkUmMCZJHLMJrI
CoK6QROBPzzuyIu5a6RW2e1uRIg/AvHotzs1H3K8u3KHOQmXDVej89CN5fijJbOpqU+h9DTDkRmB
PP/zltorX+BZnWlPNiYITq7yAxIpKWKrBs16n/tUyFdhVpK/3lk9YdVdX88OvDZvpx+p4xZLLMq1
t33GER8CP7y0pXUN7VHXT/qFkze33nLMY7sSrlGkEN/VZDBxcbF69kOy9l97A1j4MbHSGuFOg8Eq
AID9uhgNn76X5P52/WDStg/W4oXJQQC2ydLt+uJTMCqPAWY3FvZJHVaLMA3XfwDWFNzxALmcL8VQ
x6kkREshFql/VUKfzFqzOBjrl+stzvZ8nz0kUCCLUt8eLpnYu0NxmX2mY+GCMJc2cr4gUYltAuRk
JZospk0YAEdUIRjDngAKP5rlzjv9bLtGmF/YfzgABR/VmzzQ4WqAWTNxSskQPdi5BgFjEmpTnJaM
w4I4Rus1cOhPKfFMRig2kZ5bE18A7dOrvq2QUzyCAIsNRnw4lXRi+xBx5TyU0LmdFhgHP8Fos2G8
sKr23bUoDydCgH0P3omLZ23k9bE1tOnymi80xsvWInXuIAaoYtbFVfsyRrmyWKDvY7MyXqdgoqtL
wkIZeFL4Xk9+NmFVRlV+lzqlCBzhkplY7A2gXnzTITHJlgOQtW2aXXWuep1058EAVNee/SsmGvDx
TrYvHRxFF0E6bS0uZwxnr+vbMkSd2pM5FzEOYGYMLFw3Tn0F97+tEcpij/uG+TmBo/8pw2F70WM0
BMZa6Bx5OHZKiUi4zNHz1QrkNkMPWdur+UGXzaFVKjvDLrwPZgdYZ7k0LleqlavG/K0IdCuoahmt
P3DuoSkG8O/HZTBQuqVZh8zY4szNsSDcNKANU6ED1pOAiqo1hzu7Smq9tUtx2PKmVQm56+8RVOI5
pqUZv+nwqqr20iUF2O6sBioOyLX5RtOS3JvCDAM31zZ23nNK7WSaS91YMLJLtqS7L3SeBYXSw341
lcVDYxVRrQeE+V+RSYmdaTCH+XwkQvvjJrTKgNcmQefG1fEoct66Wjc/VsYBeiOt6AxOF8w/LAv3
FD9cMNfHNXck+Y5eT1m72Ob8MXGiBCONougeJhKX3IOIrMRRZGoXcS27YDi07poKmhjeTDVfylXv
gK2r6xBmejlFHriQpja/76N3QyjoDD7TjkR5Oglc9/o/ETGXRn6nvB9Nl67KiownpJkxy1QtLLS2
42b9dV5LUc5UnppyXOuxtKLmF/pgtyTuycqeIRRtfJjUcHxfsb4DmiWsGs6G6YHyf2T5Uqpg02GE
l75p7pAJQ11E/bkmQVlIuP/xe53LiUGUfOouVwiuw7JhrCPchegdwJOXdt7UIbhnwYmfxukaxutU
IUtPrIHY+U60z9/+l4XyJfN7//y5xgC250J0j91kolWgqL/Ke22gQyYtvBe8OvJ38PWr6GF3v4w7
fOjVX5PYfFhVZfs1bfOTnNV08NkTxqL7MZDKg1SrgDXiDSsCHX+IfPAdL02kknNy8h0+GRyzzkSJ
6oS20Xd6qROYpLGZorYP+2vrnZgADtw7A2Exmsvuc7XyD2KDFNjKGGTunbOs+RpshhHoA5dh6huw
Wl++jReg7KiyizRhAFUDJGRcHTnaAxrtecEq/OA3uweEXjddVdQpkVByQns2SSjV3rkcnsOtpcIG
/eekPirVXl/L6fNZXiuo2kYIn7bFuSd3sIAT092HmeAcpVDHmu8u6loCxtbIzzDNgUTaBLckFS62
tUVh8a1fTH/+NLAie3yzZa7FJMYD87Ov2qNh5LU8yJ1+xIhxGffuSNvzHMynwvB58EH34UjUMLXf
sbbq+QY9UpWvErRQ3ZtRAhgtxWt1mTUfmFzAIs1RcPyR6ff+p6/sgZPn0wje5lqZcTtDsM6E2zFw
nDDWmomd8RNQZZ+oEgt4eKD/Nk6TzEMpvIui/B/XaYnAUQhDNLINCIMDXnyv0EKsO4Gddvx7dS3r
1UiqxC7hUwiU+xfNH3mRh1XyUoYP0wjkUFMFshiMo32nrx6tpBnD2A/ZIs2pAeB94mRWFAwA5mKm
E4A9gXCsBhY4/Zx9nTd17+z46B1pY447lqlYwUBU/D9EqvHRDIMcA4dKeLpJNzb7LPj13Q3AzanP
rKficvNRt6nB3xAIz21jqSQ2+eS0ztvzbKBiilwEJlaDxcU0N1+PjOSzx2C0C1g0MT2LlIwp4XEq
7Wyg7cQL4tIECR0PWZY454iMBPb/Q8FXTsR2JOTEA8IeosDbZADbhrmkE0Q0R7WvUKmekifYjl7a
hw0N9gF4DFnJdspkGaYiEpS5WVHOvDHr+xrrDNXtkOR45k99WySjZCvqMPcMuPTgTV4bhq+ScZzD
tgA0UJc09NQVD/EoC6aAyAGjR+6ntVw07g7rwcpQKiKuJDyU3XJqqAicP0XDWToNN53waUeK91Ns
M1kF0tHoRN/pt+tkJxq6i5tXD8gBv8upixmYXzCxfQuDiBVBfrHi3Yqr2Pn/fkKPl+Rl2rV7FIw2
Q1NwWONaMV8QNQAO5MBkTep8qrybft6zN3hrqJ1fkupmQy5roOh1CdrH+QsFd+T6kXnJerRc/zte
GCo2N3jUw/BNlqYQ/G0d9UeFQ5jyoPcGxm/lz1ON83HtiUoSkyUtcLp/Zm4pZmUMBDiK1srCz1b0
GXMHZ+TOP3Hz420iyk9CiSxbDDUjZBQo1CjpEBSn1cGrYLJZOxIs6G6B+ZIeWIBvXoR/MnITvw3c
o6qWJDfgvfkc8rSLdv6jwqjZ7Mf13T8HliNr87EkAj0OyeR+03Z8ovWKijqOPYmUv/mn0olEesDn
0XNyf+DA9ZBuQjBevabIWY3V0sF+oINs92fo6MpIS0gUAhAuCuKSMV5TDOltVUYlfmSTA9/sq1N+
zk2ZvvBTSL8WKduAXeDwWjMTRQG2+uzXaZIeIovgU3GbvFilvch86719+KvAo+uIMiuZICLVOZxb
ty4cYAa10LerTbolt3nDHZ7BHpD+7NhgZxhhhcZcPd+JIqj+7sEC5tj6FojpZSiYxMAcWCGCuCz7
ZhL7VJ95HAwP/sy5+B6mItqU07s4NN4RgS+jolgVNt+XJVUDcgen4SChVZRtLopp73EDtnRv5AYo
IqUeYSg3qA0rNQa5pm/EvPEOYolai1httKLj3onefsDtSwW+J29CjGTFSU9/YuTJ43+ILGaNN5co
VdsrjqAgKuG6YBECIRJs7oTh82ZaGI7T1UCaCV1emt4RSlsk5dz/HNm0ONNfuz5lg4Rl/YFgMoFN
yyFXIHjVIqh8Esm8fvGzwH6iGSDzYTNMmEu5Yadw9YtD+4YmNWrYmqmfSz10g71inFjMb7scGBVy
dFBeQBOuiiCcNAneO/FCIzIoq2mOchOzMbBhPT8eDwI5eni6LcWYhXogv2Fk5BSkpVXSKC1H9pn6
hlmw5yhL4HSgGaDvgqoMDX9U1441B/JrHJY1Xg3hQQmuE4nagcD/acqi9AXc1UlbWnZwIURRrHPu
VdcW9AxHyuqEpIEJVlLj0wqMMYuOMwPgq2Ud/t6QfxIBhMTHPwCynkP/3L71Y38s85jCd3V8B6TX
+yKDSmVX+qsJ5GwDxvOmW8BzH5T5Dd5BOrQxR9lr7fZxQwfeWwhVxZmYDFLVAOiRTbodUlxuci5z
sCm8/9hOoGEgjJ6W4twdjMbI6qo60pmtra7nPY5l6nNpnUmcpypzkIPJQqeFiEV7Or6aTpObqASI
Ic74e5Raa93L0OlsGUujokdc8Yq+ifj3Np94OIA6S5AiPzsR/HaUk6/3U5WjBBOlh2rPalBQMqU5
PvZ/AQ8UozGm7y2o0GU0CWUJZKLjLMa1cjI3IYWZtrIM5EB5J0RLuMJXOPPfUD49vl3bRnkZiTmW
qFGakbdWl2PPfRy8hYQuaackcpstxmpupk3pK0A6jAUcPxsML0ln2CVLvozpWuym7MeSSFEqvR9y
5OZ7SvdK2Th33IheuMlNRnDj+4+8iJw57EVUhuEFK7Og4qF7usu7Pp9oJGb5m+scBkZALa98BZax
4rT0dMTJh0+upiB1hbNMdczDo2cN68l+jIx9L4nnQXEmqI/ABaHGiMlyOgkRa0H8RcWTjOdDRSXw
UFylhijkF2r5vtQbHxdrJSPrYPy+FMsEYbe18UXbb/NC8oH4jXo3rcM1z2zM3AJpUlV41TUB9i8M
rde8xgcEOinJ89Dsm3/xBRv55bfC0AUB86UG4AZBPlcblppjevnaIrXZ+AFJ0xH//Ew8TmS/tvra
JkacHVI7AQTaaPwbTcogR44dn76SURYUxW8oo2C3Oj7yVLweCIZSXxEY1o6aWcvND7qsiWG1RRPk
Tx0gjhJt2ePrAxaTuodDjepd0LLTOBKgUKjRMsbKwON3cwWZ9PnmujW+lV8p8+2j/BuUR9fcQCGF
jTq0M067sQOOdto7ME1CFBh25LQlWz2/n+In/b0jPHAxEPCFksETt4WSNfqlrF7ZttY14d0JxBOL
ZU3bYR/j3KJjEE6FvH2D9v3h6Q1mpdvyNeaZB5stW/kUwxq42GJtGLzAHjiHr6HED8E5Zrdq/tv8
m5ajBkTtqZgBT7EdnYokFdRS2K41lUhZCIaGjledwkCIJ6Oxzlivxb/qK/aX6GBWkcVEkqIRt9is
pY/g3LCX35qEt77CFwrpsZxnmAsPoYGehf4QjxpgoPjjiZL7Il1UmgQ8d1/FOjh1FCQNgJO035oj
5Qb+SmkiXx5Aa9CgHBbV/OcDJ9IriQul51+1gL+dtS0/LphjfNfunuBPYmB7px7CoBZJParLYjA5
7RkqZwjPNHYENBvKZ+nz50aESyoJ6+gUx9wv4tV59WKmCyHXNrabgbab06f1Nhoa8yG1El+sOO6N
TfjbdvvsHJST3CELEJl6azBPhP56dlPq4BxwWJnosBlAk8kVxWaGKwQUK5mlyaD2drm2GzQ017qe
RpmXnLhDEl0nVH2580Ax5oWX7SCbE4ZjN6JtmdgqxN7C+tKgS4FmslEV8ReVprnJCTP03n4ngouf
8XRmDJo5E/BsIVkvg1a6mCbyF790Wgy6IcKjbXMghWhBJOc3dqG3dnFe+mj/obOEvCREPzpG7TJh
ltq3wPg238jnFVI2M2qhI9tz9h8usFHSJ1qBhJw+m4KAsyYFWfuSZdL8H0KyJO24IsETIdw5dYxW
J0qRuommsd+yI1uY4sDnuXduzLYTbyHGsKl/PZq69vdfqcesMv4IuA8st/3cUUERuo7+Ad/kyAdY
JzZFSm9Isw66vpIZKtqMAdELI7wMvw+xyAaKwwfO5VOvMx6vnaAE5u5TEB7fUFVsLHs4Z1R3SmRb
DbOnE+5cwb4K4CCUUps8kJZ4cf3ni6jxvpfHDiu36S9ND0QBcdnXwCwVZl1D+WmCWnP7RuRkWM/H
VepNyQEFHTTMyexIeuvKK6UIdNyja781E7tjdUGuTxr7Q3n/m5YH4UiHXgJGqr/JvOfAzqVcPSMk
HkvDA2A48ssUvYkCzD3n6rpTS01rFwsAgHhUJtMeLLtBaDdcGUD/EIADqr+xOqqSydSS66fUiYwi
faA+f4PxgW+++jdJaDtK2gYBWCkhMeqojCi39MMYhnRnTNDQGmDBw0wr9+VziqFrYzM9zg0vDYtq
uPrvRXT7X9K4mkWB1VzI/bKcmBktsiRDNZ4oGmJ08tmAqAoToVTbg+symTFKrtcMhdXFRhSmD7XQ
xZsF5cPxtUBPalfSSUirjXeCwp1vD0Xwc7r+0HRM45EKF1u5CMCf/EtMXiVBWMK82W14PVJdLE3D
Oxu9LjQfv1ENo/uPW5tuQMCygl0lWGa76BE0Juj8Tknu4Ntk0FESS3KVcebdDgHzz0d6a2OS07ls
8WZnNx8EQ+dGq3bNi0FE3SiRXn7sW87z24lPn9uq2U9R6lIlMwd+4EnsMpdCDQ/Zhui2E+ai4UUI
UQYkFV/w6kqRijKDoFkIkgtGEW8kfxQjOzowcogUlt6GUbmEiCmeXZ/lIRBf3ZjzngnTJ7tRgimb
a31hB9dcLhST2Z+h//VXRm/m8BWZbZnTFFSnp2sEwplUCvcJg+PJYwsXoSi8E2fJUz2npY8WwDYc
32UXfRnGYS+ybBxvWsMmS57MGctBDO2cgm6V9IMOz460BlE5qbazcwmA07hnfKWHRdsMAE3JHQoB
+JJDha6GwxS4XARcQZO5Nt0PO9Op43sokYdJQ2BRRa2F+xN+GGJHN5EqlCRqAj0x2BlCdAnxvno1
OcToAx3eNCZoHQjX6CZitsAVsuPI1sKfzCAK+C8G+U09vyBOXeJwf+0ndqJEIha+udotMszFLCf5
ht/WQTWM+wlZMvJSDW21go30FcNEeOdBj/VeiHZKoSxHnzd/HF72WG5Sk4RFo9n+S68UuWP/BxTJ
vfYVvqRGzfv+yNGnblpgyn6jttQ0vYsSHV9QyhHUVKJqn1vhz9TG7o3OAFXXIlv7yF1WRfdWdBkZ
R/a+l/xwd+iLhCrRB7vBaXlJNFleqk07AmraWgi+npIveitLAhvgn+lANb+pxKg4K+rfEmLLa9Ai
tR2UFSk8AMSaWkl7kQjBGwuQkxwonrPeD2e7jDQa+VknLhHvZQSJ1zi3wNS7vLr56c0CCF99mLJT
vwyVWn8REf+Y6qrAP8QWIeQWb19j/PeYEZQRcdtlfq8JJDBUyg5jEGono+dJVErCciLUpARltULT
wn1pvic7IV0LOhNt/w+SMlIhbGg/shLdM81AhuBdJMMoXXlh/HgPOrh9+5APkiUEzqeAKn56zQi6
kxFKB2KcnXD5jL+qZHkAFHGTcw7EQCkTPnjPSuxWuN4DOlZDDKi696Wz/uFQzJUKu6J8nSIWF0tK
m5LsHUdJQiIhDa1iu1epNsiVV64N1tX8R5hfw5t1UkmemlYzSRZbMEHLj6DEt5QDBPZRNOVLZiQc
elHPoZ7WGtNtp/5l6VOqkzOxi/WreLupJY1lkmnqOhfv2yL7Myutr2BUN1NJGB4JwtY67iJtkJoQ
ptre5OuGnTSGjv04lROTKPwZt6mVImR9QKDIwlQFWYviXc9Xs6h4DXKPlb2FlCm5FrzuczHCV0du
ZrtEn0JxsUbQe1asvsybCB063N3QFstUTgbxYkhU9WNofxTY26lcFCaigJHkt18VcWdTgBFAbOhO
Uv16ZUeBEBxlzQS7dF0sOjRlEBnT17kEACEcSOFyr5d0eRl90jk1KAIQBdak9Z9MC3ew1x090Jv/
2kEwzJOMuXyPF3usxMfLQ+4enoJs4oaFv1t7L6evn/uAS3Z5ozmewqoYeXeq0mtN+t3vk3VLdVq6
7LQUgCzB97JvWWKS4coEMcpVSLZsls3uiXkUiDV5fwHM1Lzq7QZjNTbg8F3Yz8/L1/ZC/oHY5DpE
TWhc5yzMK0s3HYY2mkOs6AMu/Z35I9mYo9+NwhFGa8FDkQLNuxNW4uAS2BuVaE0NC2wPfgUFzFIk
mN3AUj/G6IDiFuemTRPoOSooTG/oQ1wELp2kFo9qtwFLkndBDT8VYvTC//p/LuL58969WQB9H2cA
9NbRBQC01zJgEDqk4vEfIQ+NFHUZmtpPmHKk/vy7DWIw6C/8Hp5qYCB2RCgVzixtWjyS1j30Qyly
odjsVh6JCq4G1j9AuW3PLFWuEHqovS78FYt3X1WE2mxt5BqpIGig8us+ddpokbcPsApIyCD5MpkH
/XzAPHpGGKsq5zWxbQkjtoAlDT24cVHNG80KwtVudANQiRUZTStTA52nvPuJkufy2xQnghWTM3lK
RxeuWOKu48khn1VP8+34XL9d9v1E396PCkFd4WQ/1Yl0YLgSdC/k2NAYzapvgI1UKpwlMLynWxNp
N30U3stkes2v8YMU9il7uLj3Rag3ubZP3+SaX/YhVK7ZUEPBkXbQFnvRv1jMklHW5VMfiw6tuZ9c
ie/vQnoTmuEhJtJmeMFhnZXhEDb/QwT+RFS6PGdbHVGUrewm6EIImwlafalo7BNI+lKsbwPyx86d
FoKq576ab90zCmDTfl2aLsVcNjpz7lw62ElD0lXUfdxcez8s0vM6xFHp6ZJOTIvsY2U1CBKKMuui
C0rXOqq0G2dlruLwUMcC1IcCG4cuORBcyWqzSqfR9ZiF4xr16jKapkT6CRWoSKiJZiEE/0gGV9d+
sO6ff2zLdLfPYhflN5EN7fNNBvrnGMbMReHMVLOzvOcphGLxQry2HP9UFtpAcD7PynaPS10heAqL
JmqTAA3Lb0eppqk1ZhyvNnng5LF/yViPDA1zmpjT3J6FoGSb8sA9gTGM9Z5fl9VeX4MXc3O38GJS
r+5vsoyzIsR7ie93ZfL5bAZBhLUInBphFMlpp/2DsYRSaanEARVcritjVdQ3F9mqwWk+nphXY2tm
kDxCBWsUhVK7qU0EwrcxB/2j4qbHkdAY5cy7and1mYqFDquB4DErqQYFVezhk16g8d67DWfCGRrs
t14woq+JT0jvSHo70snikDAzapjlbeuLwkNM9A6Cvg0I5LvIQoWZKzYfpNBMHIjB3WG11/pVZDZc
WEX1tE/PSq78h9X2tkqV74+EJ5K0bfoGmnD2g4highg+r6sHWlojIz5tZirChYtssPkZbY9O2jBY
5Fqqt1V9lRYZ+oI1ftx3Z2kgOBStFAxAlLCsf6IGHOgkufL4WoNBZBmlfavrHuYVAGHPPuG04Az9
1uQQVBnEJtg2droC6dFecpKHYJy2GfVRUHF/CWAAGhXftP8BQ5vKqJA8yorqOZj93VeJSBhnBiV2
i8RP67tHPBq+MqnPqSx/c2HayaGV9V0v6W4cnY4fmltEKwS2mKUu4CRYgXDCIj9I6c+yo2Ebofzn
DlebvdA8SauLnPqtKjHmCJzETQxti6ZnE9Q8nAKCy1LAk5X7ONPZctt6nfOd9eqEjwnzcmrUdrvY
6HGjr7edmp03+1Ija5g+J4QzTh95usi7NeDfUief5cmKQI1qr+OKONZd+OVMBfJHzmKlgrEuJ8qR
uSWptOf+oblowG/cRpbopC/+AI5AFcz0eQ9x/Aznix6mpkWroHxPJS1qpJsdOmdMNIAmPuVO0L+k
qGW5o4M2ZnIzNC2O1l73wog9gMztqkHWBuVGMbf/NH/UyJZW8rs7eOU8cDPwSfGYSP9c0fgKnMqF
z0YlC0k5XPVCxX498GDS3DZILeE4sJQEMdL0qQ+SxCDOVx2MZLX8sJbjB/sUspBltn9qsTMbd+Pm
jx5kUoHmcYJlNo46OuKMLoIURoPB3RPg9f1Pj5nBNiyIb2lNFC3yl4l6gpMtJMcOxnufzrWalfFn
troJXxPctgl4r9rOeix51W5koL0IUpx/PiuSNnCSBHq4Hq3cPQKZE5NZWr71QDKHuKr/U2dT6vtq
K3oziIw+NkNBQK+WNh173AzHw1rcxj6/O9udU2qmE8fdSennMXfvUOiNpbeIet8qVMQRncrmDunU
Q20RzpTtdwuOCu222YCyut7xMDP+oizO5MFVyey4amJYs23U5DDSviOIj2OnYXY8DKbE15NnLIQW
o5/XvGBrFjNg9YQH16qfZHkj03Vcf1X2KbEAInXR7c/uytXw76s1ViYpTF9PXXqXdWYmEPB5VPmf
ZhT5A3njJbWyo8+xGvJxCf99EH98DT4mVIPS9RytA847JqgLfKGlakJPkXnRw3yV+aft5CW7JSmS
HyfZMcb0fOJxR/g00aMq94YVOotAH1IsDSriSsGetmDF/xhOMFUV/vY5/m48aIearBMl/DBLBMKu
r2HcW1GBiFlFifsvy37qH/F6jadazkPYOz9pmxo3sx5QUaparkI20QQVXkerUBWzJbvKB5eDVal7
4HcM3LdmnLqn/3NvbkpV1JbCd4MROSHICqBqAtJNAr7BbPDMEESAaPwgxK0Qeim1jCTcjsrw97qn
HSzFt5DeYq1UP328qRRmUz7B9+kgTCK4uBrobLB8K+GX+uPORl8FiYnmnW8kDwNwoVWpA9abcyST
ZrjwiwaqK6cxJmpw44XyY2yg6TzMpHI8E//ra9o/gBOkIJqp9Ht1aWGULk6PhQk651Mx4VtCvi4h
za7m/8Q8uhdEn1fwl+6oTuCrkIqNZM8fFAzyUcHe+1KMLJBupeYS9mrirM0UGPc9XIWViUFq9CUY
7RiSm/Q3BcapaM4AgLSvAhoryz80qUApaO7u87k2lpOdp1qQ9iZP+nsxJLXbKFEc28lL9Cz+shFH
cZDOce5kSBH5GaYivSNmfVOFMj+p4vngDrGOzZzF0T2sMgjL51K85q/vl6jAYGx5GA2l8YM0++QZ
PGPj2nsKLU90IDBGpTXqUVmL4G+v5UrxWRFJwNbpI/DACFFSiBvGG17stBwM9JX65QuGdmnbiWjS
bHa2A5WjLiSYREnvZzXIKfzXI/+ZnzKQ9JcN+d8bm4L9a3VZNdH4GcHNNTZOgDUw5ffjGhZ/d1wk
hrvP2GoYjnqnmNqkTgUuA1QiwYgg1YrE56zKdgWNiB+8LbzkcIyTt9xuZIvxHhdZk2GpWBuczgQW
lDuVBFsHZY9TJwjl8ADd9mGvBls0Ruv1p5XvZ+uxTHiVFZoP8Ae0tMKhM8whpls0FHuQ02IokLux
AUwRh1jnUocnV0HVFbup70Zn8TgK6etOGVI2rhVWx/kbE5xpFwBwmyr7+ncKeuqPOt9upEsJZ2l9
UTEl7yRwWM9F0UQ7T2YkfOwuLPQScEPyEX7gYW7o8kGE4GpHQBQBF+X0ljfo6DkcU8XI8ZA2Yp7A
15lh367wv9n5XNylqFqf+PTxVSJFbfmEdfqlEQZmY2d/pCcTNTeHgzgiSwwgGk7Rq8hgSpi3SY2L
nrWR+gRvJCd8TJJrdZnw+vCR0YcQLLXvxOBTYYsz+cueEbw7QGkNZPFTR1TkgijNInzRIxM16QHU
Q5d+FeuOkhRskUQVapL1Qt3BnLbHWyxxxHymmk8r7dfc0GFRVR7EuTNteohwCxx1R3dJx6mUQ105
tOgSp8uxwRWsQnQpvv45tV1Q3pNyNlQPVVgt9iZKTu43shNs5mle1596HiAq6Ff8E/cgbTnBNeDC
be4McYZNEWPLE37QmLf+OpCJMOWKUHd/PbGb002M4qJucGiIlL2fEGfmDh+nP4MyzqyXmJNMMkJS
6TPl87RqsnunmCu3rAwXngM7vtDOTXvTyyxqsm0NNQHcF4M9uV2e5GIlt3uCzfV6MvzNOldURPns
5/uyWEYI6l2Q4N9oH2fscs5IT2OUGDEL+p5gcdzUY8b1pmfEEid1sgzIpQD3wEATnu+ngOMPd29I
ShnHMwYfwBxnWOYXpYqXvRBhNILTUfltrpWUOS2hWQVV5hyZEQ56rRV5dqx75l+VDELH0TKlirX0
FH0ahaO85woAGMmiRr6cDzanADf+V+WoNa9ek6IbfeJaxfSDWVV+beR0EJpYeMoCg870peWjq11r
CxjZS3aVmc5J6dTRVTis7bki1l497FtsVhdDWpRXGSNjCCXw4VfLUN79+xITmcU1Uz1XIe5rQDNe
KlEb9AUKggy7cB+rolSfRVO6n7IxDF148D+2I6FBBEStl84fpvDLUZXJuPswaJYIGdUP6+JJMSC3
wFyliLLq5WLS+nV8PnveZy5cm7ZMoLh88BDLrNuA13wm4p+BBpgZLy4Sw+I8bQbD3YccRawptDwc
XvqrlDd7R8VOJvwSO+Ia9PH23bred46HWezK7/jdSEpvq9FOaHRMsbTNI35J7jWTmPrKcT9R9UUE
68GLSxfSwAcXq1wev9GE+ikiznbkiKGL2aKoxC/HEAxD9nX8tFcUXn1oN+cTuRZu1oxJwweShENn
XbbTlalm2/bwvp+eGtMUfAXfETKQLdXnCrwG707OiZ+V86hG3iJBYr5NtbNkq7S1FSNiZwPVa3f0
ArTJ2Pj1t7LzuCruHVOdNXtqVAXDPJrxXLbWKnQ/Kv99Sgy5fc4CQDFto61Cbpf4nW3mQndYmmLi
/scA+/wJAJz0H1fhDZwSt/48/nsqylEZppsAR6WvFG9TvruLuaQnhn43X3EJnWc6IJfUnZO2LuzX
KYfa7+VMfDPQpF2OejmwPEYPC5TI16PZm6zaWl6TympinNYL5Dw6xmHnGZChkahJII6JJ0yiyesG
sCTq3ztceOgACUwLl1WdrQsJZ7LgCM7BFOyw/PX6+o4RaquTWcevLvfIoZiW1sQeukYrJWipHDi5
HrfEeX8X9XeK1QlRayw833TM4MT/8rXEAY8fiPWMvYznncptJyRmFGVx8uhBYdVNfijTsyXpNOh1
VOmkxJVcv+5OqubRBNRmw7xHk4lzY67wvZmXITOzZQ44kETcnv0Ptx1mowpZ6OHZukg+nASUe8ks
UJQuWhFJBkfxowOGeaKeIgyXqZvHr4olUeLwoJVyqqWAW/FuHd+lYwTS0bxXVFc7CA/IT6wpRVr2
XXwNuKTJjEKevcyPVSnqkLsNXZLoHgyE4usDzH4k7BcF5HI+uJRSIc6E3cQ/ogX6R/xq+v5pwR8G
NbsUoCVr9ay2DVxVBbsbjsfuBJkA51q7VikdbUAG8AaIoE9Bge14LyjjLQl+JTbvwUAnal51A4tJ
1815WW5sG0/1TRrQZSRLG/h0D8wrCPeJJe65e7EQe6mVf02c20FAU25JxhOt/3+osrZbVXf/UUlG
GSUU6Ep3JP+OeqYvvnTRNaVFuw8ElCRn2XblRJ3sOu9pRyQVz+aIzWTp549ABInUv4jlJfoxxeJ/
D7mz7fiYgvcfL5FBsOfwIoenRrBm4OCPHPWDw0VJY0HplmSkScjF2kFwaM5xYp2QM/pS7fDiplvF
v9dOZzCoGIDlFr7bKJt8ulF2sWZccaKnKeZ9x5jPdK9cBBMDfagP/NNuDqa7VJoOEgVxy2TB1UeA
LpucyghLV0Ts/6YgaTU2QzvX5Z07a9fCg4u+psbEPKqI3vcftqp50cnhKx0PNyNRNT1INKlET6/x
ODbfCCzSJHoOC5c6qJCkmjWnxSsN4fO0Y/GzYpHAg3Wh3VWUHPNJ41qm+MASjIzOQxah5B4PJOtp
W8VlV34hWP6MYEwvVNxDVkLpQY9ep4B4WC9x//iOh0xbFn9NNBvJc7W356z+P4d1hiuIe5D2311D
8B9/9rxMp7Jniio0BuyBbeaLz2N2X43MWabnod0BJF2yMsfzSIW167Wta/Ubdb0ihu03TPUdaxHx
mUhz4GNa6FbXSue7aQZgfmXnxQ5Ik/IxpP/bCGkg/4xNS1EKplb5mQ7Z9dPKnhd8lh10ZgzvJNHz
Z+giYE9nrgNM3cnM/tgv0UTHH7g8bHIKh+x0jj6Lmb0AMf5XohMkVR2inPZ+IcLkfpnohH7MaHen
Ru23aXQOZcVd/5g8JUo0cy8z7W6bWZHZO8F4lssq6HTVq/0JL1y7LNKmWkGs1tE7qxSMTI1WGGUO
8fMOcz4OYYr+esHk4B5RZl5Hf0dqAsWFAW3n3Fnd5o/tj2suJAz04JFnOx1DY1Fuw1VzcTCV1NEN
5s4SoDM4s3/glkOdZzwzPsGIBkLq9d6EnRCNSOrty2+M2+OOrdVK0oikjEL/8Td3PBf4HBFR1Cim
30nevGatQrCayEiHMDA6qCr8keF7R6XZDUnt1QY0sABk3fgZVWW+2N3uYjC/qlScvgOyFbRSbJrN
T6e+81rqQk79REo/FgQSTykjXslwNe4PvdAjtC5zmhK2oMM3Lv2AidOdJYT3ETC8ZVYA8tzpNB+G
2cjv0YvSK2emE+MEXlc7GEf6O9O3HJhRbOwlZ4W83VP/hDK2MTbgQXa//RBg9GOkZQ4cfjgN/Xqa
xvLRhslHw4XQWV2iyk2WRofOX0W/4xxU4uwyrFgVSpWUnI4+Ad+a1PA/CWaamgS5HEzUOKQe/URy
Hv8oVFEw+aIVAsotEtyWA4ZpPCqhoiChLO7v3Nt3e6ureUG7w4mdQDiH7S+BXuOAq8ZPPb9i4y1s
0WO5g5GEb8IP5hwnkBChkaiJrPuzN1zhMDs0wiFY7Ymv49BZjUsdDqqg4yZfi82WAgFT/Fqjhozo
sKmsuvO6ewM3aus7FrxCPfHRATaEeUfOaJk7+Q2VZZkrygpB1AN4QsMeV5nS+37GJBB/kv8uVf9s
btxUMllZyilP/5vxSqMLh/lUi3muSipPdIenkUkXnWvyJk7gUTZAbFyK6ctzgBUqqKuIq5pjELyQ
Abjp/299Isfec18fjVqTTVlpBuJvktHDqgRSNRLmo8G/KGepO2NeKHpapdI4lnJrcwY+iovmZWY9
V3Iy6N9KCig6qxfA1M46dk6OaGHiTtiDsrZtZdfTDa26oTXxg0s74RE6p2zLw1mT/66RHyeBsF5p
dr40VMAeQj3wBI5bch5ZhKaSRsynbvOnoCRfOhj5d0D+q+eILbJWuP0kHrJLgjUY5AEFrRjGWESP
I2Xjs1y/ag8xwQN/PoNdJhob91xjKDhDtRqlFWSzdGpR2EjQfT+//ah6b2+VKq3WMQTs7LNK/Gty
Os8/Bm0nrC4NTHdhCRP+9fzYXoPA+Rdw4VUePgVNBAPD48vNLDka151f+XbBk+ciyRXsxeJMDbdi
NgWSZknXCRovhSsCNL+abIc7t+c8jkW0RLjGtginOuTuWGADfif7S1ImsPXLYbeuAHbxwqMWYI2y
CDpkM5/KoVtQnY5dSupI6Wh+UT3GqlOW/deTT+u3XSAte2YZiDwTLv5vbckuFM4VA78AZaYi4r/h
D3QvDV16WtFPDLPos/iNpnTZ1hHODN3AkPrZF8nndpKn6tKpO/nzpjKJDrZoq/fRbc5smA4AhUfx
uH8q5e8CkOwnv7rjoGIA5IGlWUwIejcjsLUfQp+Zkpe4e6LrdYqOF1UEyAZkDcxnPxcUePCGS79W
3IRaTKTBcUh5210ZiduJsCo24D+pRk5OlyMBva4qO8A/d4vgAxq5ses+X8F+Jht8FKOX0c7R1tXK
BCYxbyYeVYEcoS6rMOPKMbWP4z9bBceIBUAbxH+5Y3eHLr+H06W3LmtxA9tXfDxPymbztgBAcVCT
EoCemXG933u2lCY90KmlR2cHuNN7gtGECt5H5J0JlTFNxPpvHZVy2gznaiNkXMA8LNPV6nQqSSmq
pHF1ORmd94+DM7PU9voOaG3E54XE1PgnvJhcKPU5kXjZTTEkWtwpvSTds2jx5UXzkxKurtuFy4sY
MP5tyYefd9KqBMBulg2UyD/f3RTCUw3TJijTVo8SRS2CouLCcCvl4zN3JSbD2Gbjzvs8WT27paFr
C0iPS/UkR5Tnel4yiAGyMpfmml5VzHz9s983a6qmbwtYujN63dNI78DKATyFaZWpfFi3s6TxPLqU
XCEev70Uarn9jlPXXte9vfUzBzTs8JKXI4rKOlqfuCER83JnAxvpxiI40VoTo9UDOzGwekU/BZcU
lNZyZQ7emZBR74OsfF2cIzl5JLQmfcaIWKal1suJCFgSalJxjsto/LA3Y/YR3qHDTWrFFsxG7vpk
9xioys97EE1x0fhPF+2y4rWPFguoXHYAAfERFY9mwAuIk0RHjfbgToK+vR3P9O4rdsxBknjBgzdS
Br/K8fcx5UCiIzK3P9AAnnYzKp5jU0Fz20mpLzHU5TQ0hXY6z9GtBDDmIRZT+xfgjLdYgJRtjZPh
XmdhKWBxH1e1Q4/Uqx2w9BxvTYIb8blp7uDGdOaKpwmD5SZvqmhA37jxXY3NTpKV39KLTVYaecrX
4NTMhFTZpwZsN8OnG5pemWN654WfIFKqcQNury3mowKEoYUel3CLx6P3uhTS240Mq0Y8J8oQQLpy
OvofYQiZpWj+ri87MnDGwKs0T94+5eTkW9wuVkq+rjsHzuITu3mhF62Y1lBhEqcStqtqJGwkg0O6
lE6x1Ia7HFStI72whNwLB5ke9oT/HdQjbzE/pgkP79ppFaTwpvhCyfUZ/6O6P66RDLFY0qD8suDd
n8TIqo8DGf1D+adtZ1+zN2GR4AFvOfvePpIUYtar2mpRBAg569tWSJu01KJ92tFGit27VsUF+BS2
QpvqM5AqnoWt1LQo4UQ/ZmzUAMHADlYMJZgA/Sonp7ylFQ56egg+Bfa/S5nQgCyAgntS0AB6TqbX
tziMTcvqDu66iQbYyLypIlVybRdiMA3QzZdxv6CnOYto9WR6mCZ5XnCSjlbnp+vjZHl7lXXB8kt0
+FO55Q811KNqoVX7KAg+OdoDLKjVaflJrGNuemXuhk8h+oXnpmlb6fkftfmMZV0cLv5J3hRccy86
AKz5cY8Jwfy17NJPYAJH9VQen88+igWQAk0Vm1n2r3+XhaYwCbs0qEYcDNCxsu+fDmRRYq+HoB07
lxV4g4E+Tmb4DjhOt8SHlP9YLMmNqfQgnKolZ/SdyT+Wy6naBE4I7/q/xeSjC4ctczvtv3deljui
GMLhzfQk1Q5P+Tg1PbNNTQnjsCQJVb9bu43P0vxpyradtvvElX7f1z3gk5auxD71vbXJRLfcp9V9
g2mzDPl99kAi8wRKM/G6yoMw2GMqNoP2lMJchZrm1sdNGXhRTOpWAEhE6GIY+dsIBziBY04Bt8vt
esVD5jEmMrL1ftDfhjNjM+lvefIthf3CatoNfpFCRIu8j+NxnR9F+RXutsC/EQRaF3E94ea6slf/
0+rFCwqC0HU47h2J0F7Yo+hXzkLY2UAJnYplbUi1m8fSF4At2r3eccoH3X+nl6GvGnrIiK33KQ6A
Zs6vUu1JQ6roWe62AeQw8iGn5BgClhHVYCTZRZ7fbyv7EEB5juVGTN7UM5qdkKMYJSCXzZDX7U0r
YLmgZtxKFLhOKyAMpw3E26LV/OINZd3iEzTrZ1B8BMe32i+sRTkn9igoRwYOTBWsC679MVg2pYT/
/RbGCSTZEuB9Fmio8zEslkspXHJWFR/8yygqc68Bv7GhlMnZdh/JqzuipEcM5MIv31lUaPn4HuaQ
4gjrtRK3887CY81uS5d/8ccMt/RepkVB/HuDU7AHvjXuY/yr5nX6WZfZDBOP4XOo1TKqmTjEkBU2
K0zO8ZE+d156hzooaWeOfzuVq7n385N5Wi399jQzSDhPoSMAkUnaen7q+OPaEAlgxjAZ2SfMkC7a
tiEo9+008SoAApWiE7OhXKeNzh5MeUSmxKQpFIbVL3OAiB6bn9WgFBd/d5CcvtCegVGtzzCVaNdB
751hSQcj3fdMJg/Hh7eimfm0pSHaHtLPE1xs7xvll9Gcu41G1t4zktew5PglCdBAlZrMaMCWNItq
UQKGfEBbwzmJw7FbhXHZOVp6LgpV+a8emQMn0w5X8wsQsXXm2sPkSGiVTVgM2lB811OkslWFw2uM
4QJVM9kKiwOSylYl6xSdwgcOVaVsABSgVideDTWuQYsG0IXT3vysfAwXbq6cDehtJDmnJ/XkJTpe
Z1cnCiWm6t9vZucEvNHykQLWUq2GxyPSSa/reIXkjHUzqgWB7cnbxmQdHFCat3lyfkY0Khy47t+L
iTY8JAXDaIGn+VMr0fQNnJuEGdMnO3tuRSVmrogtVK0QSHOU8D+5HtBRcHJMJk5CtCSkpEYqXdHk
OAhXpVFcSyq2CWaVzngIRqHbCUsHS9cBkwyECBs7XbY5jHomMTo/PwCKaARBvkm+Kui1sH5HgvnI
6FCbsB5POuFx0DLGEnriVz399IVlpSnxgfcvAhwojk3SKxPifvoqmyHwJx87DoEpdLhpjMbP6u35
f4jYgDDpwO7hWdiuDeITgUdgVBmfPXt6YzGNfOPtHUfkiMxstDy+Vkvy6ZwrY2xiPrvd06GnwZlg
aovnb6Dx8xGxbzOl7k8dIN0v1YWtb0KesL9PIamedz7jtJR2NXSOXFIfAPIzY5rpvXkcto0juo/n
VSLAzttQ2HFQiO+UgJrTjI+xQ/UbJHqMgUXn+M9urU/gRBWrYcTsqatOCrmUIbrxJGKWGpWHDhbG
U6f59N1dgxAwFv6FW8oqsOy9lE9OnnCYocbSE9xHzAi2VZ1WPYDINWjw38/OgoWEIPqE0M4PtleX
RcaETA7wvjURYHASk3SOn7ZHg9dPieC1PfyvEjhnp/LPfgvjLoCd5H+AZ4IOgzv9LKG+Z4GiNhvz
gRHgXYEtJoJAv34Dga7OA7qv6fYDLZFMaP16yCXI0nZhb1SxBhvayoCsM2eUjC2fB96wwf8jxS6j
Fo084Oi4ulYwmwdcgtiimjwbTqPcF2UxtOGIjO7kzyYv5zYa8t5LZXtJ8zno3PG8FGWWnBYAkSbg
cny+TAmb7yZFbxif1bm/Spy9ELa7q/s4g4a86zWmJVHkW9ujR49oqr2knutAI0xqNG6XiAL7Vxua
y8I4XEnuQKrYEI5x1WtNMA8QKy1W7+BE40ivLtudQrqEsi8XuzFbr5UT1iDNmLpInFNuv8U/hRfY
bgockhv7YQWuJjytl3v1/Kz/CU4tY037KebbyyPM+ErBpYqkkTtygWlcSo/XQhAdXsGTL9jkkjeP
Xw510ITAOw7CMePnvgrak0KxWi5iPwr/7tIRADk46y8PHrYWbA7iK/isHjlIwaql2Tqzb6ehSz2M
DaGbrFfuwv1xGVsDhqlhyUreLtPZzA81t2YpApLjLnQeMQzKttf7+1nV4vgUVvfMQaqW0ol1Lb6s
RqDlXmiwrcnaUrKWsG6tRkhHXU6elgvPC9WbS64Wws+UoeyS64N1HRXDSHwWJkzq96XjqBQfxV+n
K0nEfvoOmt5fz+9A64bX8lIeAhRcs5aXLYY+7GJgIXBBB2qbmujcEQIcSVEqoseIbpWzUoEptDYE
w74BG38blKHrjHGuxdqvCdzC8ylMaziSANkvMkOY3j8DvdfiT0S9Wt4v7W7QPPXlZYyJCbaluDC0
dBVWXVrwMKuEUZ9m2erfCOxeWGLvuUXWmIm14UUdu2U2IVsGCHoKCnpKm4C39UeCGo5qYyD1NZVS
gH0N1+mrl0y3lotEgJbASDy5YIrEKAOAqOuWEWQaxZuv41PBY1oO7O+5gqwZfQ4bjZNlVxi/OFSo
g4TZik72FfxduFIZdRkYICrJUO/Ssy4hvKLa9b1XcrNRHEQ9iOVQkOyPiqpVQSfnAVQjPJAQRt/W
qSTDD0DL5qhwhOr9r34PKTcPsqjcHHWlkoExsoeUpecfmkD+InRNBQC5HCMpTnKg8WFj3X4J6VOm
Xxcy+SUUdxDawLM0ssvSU4i+ip0/EAAFFAk5tEGIlsCt8DMtc5HIsiZ4XQnQumWUchM+QEIxqO6P
e2vGnMZJ3+T8zkmPAX2rWmRWJkA88bWBqL3s4ZeePQFyFevxfoZy0SlOKA3A1SFnwyq2lRPqOJqC
LKyBpORu8R1TNvHVqmoUIvfM6QQW7G5NWucpgEt5+BwwKXM0rTuqrmBOomDYGA1icsgZbrfNY940
HPxKtBp4PXg3KUlysllByse1kHBZXCRQrchR4/zlDVMUbnXw3IcFDYcL3xbsISgo76n3v3MBIM9z
JIBvVTPLWhgjLrgisZHC2F565FffGWY0XbhmYicR0LhEjyzoAmxTKJq0F3WwLvNgvrwIAKmlD1fx
kpDp6jmYMpfTp51+a5ikb9+TT1K6AJXRkj1d8VBZsZXIuRUeTkCeCUuu7/0CQKkTPEphhRaiS1bl
0mbg8UYjtYORok1PrKj9mBwGGcyS7OkQkJ/BNQ/2IkXIkE5UhQpuDRpPfx7MvlSutyk+Y6GwJT9c
MlsLl9vfMJt5ZnY2nSNnjYH5UPy91yUA6jrjPnRu9liHolfkNfT+9nRqeUIxUMuWVrqJ1kP/RWIl
Vdp9mI5TDblZ/kEkukPIyLE2+C7wC+MGHUVVcrexh9i/4vTR9hLDfHKEDV4ZuYMujcW1Pzn8HdbC
yBHcAWZ+ggKQepvNrMNgaAlCHhz1tO9/TehWwcf0/nA9e7lAZIL4EWGOuE7xySM9U8xbf4FWv7aE
lQCdlFUyUwJlF6CqO13JK8EDI/GzHZ4i/7uJm2zAu3xhlB6XWZqJljFB2dxIR8QsNobb+9A5cuEl
stY57Ajov70Ot4HjQb3XxPQPYzyY/Ap/gkMqCwzh7q18mN0uOUfcS9C18ahAwCMzIyehPswJ5fiH
v4JASlb1OmSpSs3HXoa+f5bI/X+o52Ct9VfRYqdEOk0136ARZ2sFdIz0iynN+DMIOG29BS93aDCc
U+HKpUwYVaBF5N8cfm6uLwjvwo8UVvYpPvmnMyRaSavf+/qBMHvX8FldJrXMCTiv76HzPXGEYZp5
IVMbSXevvxoUfJ9Ub8UjGqB+x9HUqGYobjdrBUVd1zCWoz4/oO7o03P7iS+mEIHeuKZ3orCn2WLZ
UVwMPnrn+Ud700qquR+pPmxXw114FylDqBZMeWv94JXaYEUfP4FfFmfxBPH996JF7a+yuC97oC5D
biSYPtGW1cqWeh5RAol4FKg7f97kAy+mMLA7A3+ZTq4dXxq5W2DJtDP2R+/HFUn4rCEq/j8Dawe5
b+P1kS3XdQYgCHWTBPr/sbL52gBLhvXi2ZVrrJJDtCMcoBAGKOjXA16iBGYsj7gGGn1vrukE3t0s
gCBMe5rrDRS2/xtXguycO5I7GmRpcN623dD2LTYVk85bBVHNbkp3IUu+BR49RjLQ4zxJO/vCUXAh
uL431eMMQb5MGxtClBD7KvKHZ9d25dkcIPuVrM+rVUqKSwla/peEuatblpFVRQqy9ZbvqG3tSTRI
7usOAbxTNjNGisdWhUHcPEdQOmyJLKE4G5B0VLeT5oNvEOTZWa6lFPotArAPGq3EPdVEUMP2s4nu
5dqSQM2UHIFTaVctXK5mIXXfabihMNaNwwWksc5Ze0zb2uD3FoqgMRs29OjdMguziHn6hHmOzxnj
tNUdVp6d3i39JGihSNHtvPoA4j3KIQo4AnhZ0y/iS97NvSw8rxT+t7TOGg0rH9iqqOjXkQ5fH+U0
OYLzN8evXRh9NRK6FQ42Dg6gVsiJA0WZZY+grTY1dcm//MTHI/3ieP+31rAsVEcrGs7V///zlqpN
C+0l51pKTv64u4yr5pwUnaacKTFRqTnn+l4QzNbcubtbxE4AuUli0Yr6fTaALRjj/6o3v7co5zzK
8av/ULMvOgug1QkaRNpeD/3pAkThMpLCzxegULS07IJ8v8nOMtYQTrLxFCiWfvj+puw7QdS4gGDZ
H6zhb12wykDLStKP+OEcvawFvABVuveD9GCbPgKeF+8/g5ELhBr91W3mDQAxoIONBF/8fcqSApLo
rpKI6+KycjiT1msJbIwxAMO+gwkZlALHYcUo5SjFClpBmk3X70mqI+0E7ROl0GGHhwNy3GlqZREn
cShbXAG5aIhCe3oqWKRrCRncwpa7wIOvSRMxx7YjPYuc2zZ3ZeWVkh1ByUohq2ImKr5dTXeA2xo/
HKvIs5BI7UmKwmQnoGlHwhvddeO+IkKs+FhiiyUfYpboygMaIzqcKbc2R3y9CS6KDi3pIg4NnKEp
BUtbiZ+qKh5UhbJABc9tOC0snKo/RBIjsfaNIDoXg/pph3JcblwN2XzpRWhxARxZuodK8gnzzp+s
C5Jwai01dw6W64aCsEonLuaWp5+9oDTCnuYYUwUvTud52Ml7j/2DNjub51s4TQIHPVa4CA1oY733
WaeVSEXerawOULniqSotb6EJ/pUXQ2HYH/RktBKIYEtO2ma2oKTj5djESblk59udmb6juZdA9Wwm
kmsIlkHcPdzBFfyggmCUeITS/0fmqLRtlN3VIIVAUpw9uKdM6aLR/GSkb+/NiG2LEExCtFAlYx7u
ZXPBw7TkfFubosrzZaXllwybNwHJsdoqPxbKY7FhvACw3cwhqiryuo/I65rvC4o/3fRBoZqzf/ul
cOmp2HmCalxcIJojpt6ZvvFkDtv9sgT2AC6D44pD1BC6lIOBQw2uO3TGJumw8Qhn9WZDHLKj9WQ4
xMEoQttaXr8jkx1GxCE6Mum47gxOY+XEnm85r33N9GFtyqGlkeePmXTc0zp+Gbcz1SV+lKK3733A
4PISZoQE8qGXN+IkbjgtQ5l8b1f3v3fBU1syRehYlVuUDRLm8kOzOxqeVnW1kfpAhvmpFW7NnND1
hMlw9HwwI3Am9FNksng1Ti1E5SOKdvsjdqoFlx21VSKUsdJ+nyE5PhZl4w7DLzICSteZ5w9adpee
e42K4T7F96pT9tgF/VbGi5gfnyrCJEn3s4PjDi7M9WulMAvzyhvhjEWb8dwFOOIETR4KkjEFFlLs
Aq+k4D1RpZy38zgSOX0VbgGEBYzCwpTSRKEcIMxF9rkMrb40gv9YAbN4Ydb1IOFVs1op8mqR0isb
guBwwtN5MfqBlfAm0XuXvlw4qaEnRIcW76bM3eduRLGLhFDlsa+pIuTuCslSOA2v8dD1KTx2jQkS
dzF7kGBg2A3x03UppBtR35Iamk3l3VY8nkxxTOD5G6zyEN2PfNwTSoAjU0WlwNCFhZw0lZ/1U42E
A5U6cw70nGquReMMGEfC0GC+nI1M+yxhz2b8bPwasApj4Qm/b04qWGpd/T7NbU9Iiyy26JtyT88v
a3f+yOPg4/BQQkuUMnyElqeuqGBGBCwA7j8tUCiuFoweauQ91g+lbIhoFOkuBTqGG8QgYhtYV8lE
0UTTIfyIlE+Sb7pFtmyEX9gv+8PHca1t19LE86rkNrIGHIvkLaWTi3w4OVeddjXgkd50k0ywEMJw
NlxnJARJSCYCVHVdGLLFyLtdKZ8QmfeH/J5oQRGwiVeD+c4+BmEhBKgvD0CJlB6dwiIXKUVbqk26
sfQwjx726XdJdiIhQNaHv2YPCl8pIrpJ04WYS8anQxTykw6JHHDM+g+ypxzZ6zKs2mB2f0CFjrU7
7v8h2K6Kq61XKO/qAfi5PFFufZO5sH8rqVIa3JLZbA4JET/s+qc/4tZBv6KlbRxm3ifyybMxYLnk
FGjzE5dUjEH0prOO89jyzCOuvgKcvwvk5VMS1UZq9J8tEvPkyoE2FnZGici8W4Q8e1VqRkMUpL2A
fnx1t1j+TpdeuZPOQbyBanV+8ufnDvZ6GmnN1nwph2DNfS6yeT0Fzf1Nb/uXPJN/lCwyJJ0avPWJ
Oq/AuIwFGxa2IuOoeyyFs491c8gNvBqyzBpHxF4mKZ2VQEdvzZMg2Kh8LXMd4LSnhu7RP8BRTQ00
49blBycEIz6h0C0v1/MgD/FUICO1u+fjaj46kVo2h6wvGcR+IJOquPyQjbMvJY2hb6g+agskeMxy
HM/1O/41DxBHdmqACYVWrDLeB6K0DcFbliVGOUluGTPsGUHx+HvZ6h6Cp0wIZ7wEGJujCsjsGw6J
w725rsGsUk37sbwbj9pJktd4floNFCPg8c2daTeaR1eQv08PFx9wmyU0gParEcUPWBE3ubqN76XN
plWmpxRnogk7ehVTOQjaTgBKPDtXUZYFcDyYn+VEYzTlIUE4W2QVtXcKzko134c9FsWr/4/w786C
a3t0exzz5jXapYkwueol2npSWO3uX4K/fXm4pwOgyXjBuLj4V8zSZJ5ClxltydbAUcrUrk3VyFrh
9cPwUsf1vdIEszlIhjYyZYZn9wq9VeHqq/m3j6Ym7C4Q5EqZ9uz1r6R+XF1OFZpLmXUfBGrT9JlD
Pm6T2FWhHvEfZ3AyY05gbgxrSYuCTcorudgwzeb5b94R8OMCXTwH3G64Gn1zH92rQf1I8BIF1YBG
xB3g6e267C1O0WWiyCe0CwwsfJ6JJfbKM/tnUsh3pLL1GlIngjT0tneiQLe1a1dUB3IKEHfQlic7
onIEiLxW35AzZ+5RPO3UyE6bLNgU8pJu5lATCrj1C3mdi6ThhYi2oHa1R/DPr60JPz122db1MK12
zwCO3cH9DmfHOwblSe3LMH9SWFuz356Fl/kQ6hqfYMW7VxJ1LizgK2r8mZNl5dhQqT6ZqIzIN1AU
GOk23p91zUFSGVryRyJxVFRPBFKWx857V7noUs/K4ZuW0eMoTifbG+rTUIgempGcIBWp0vANiOzO
7mH5ld/M9+HYfgCg+qTelByX4aKYbEtHUjFE1DhcpvGw7EIFZKpwUQgoZJQQ7zXRueMEusTFC/ew
b1EqBI+9yywL266zUSLlRBB1/RLXm9J/QiC3ahRjIALXAcC+No9miNmV5z3yyuD/KlS7Xf/fCP1G
ZhDIDPeosnZNhDBYxELqSRd8ZhqNknQTrl33MD7iO6oNARU1N54hFM1w9TVG+zXBd/RO1tjyXaDz
+hEZldh9lIyS0b9iuSkGWx16fbCcZP3kdbgZYPDeo+KRrPfmw0DtytjmVc0xU++XIsHI+hHlT+0Q
2Wi/8/AHc9k90ZSIMJiE3GWgnQSTnprRd5GPLieinIrCSPmHepmKlk2DUBla33JGmpm/PXx4W9Ex
EJY1H4g/3iuTcbI2YMzA1Aasq6dGtzMeFKEwf7kGeUuC/7ku3BKAoGENf1lBmuaAMArCicPx8grt
pjwT+8Z1j/ET8obAwhsXuLbdqmSlgZR6zj5iZ96CgbCMRAM57gj8TQg5+asrF3xBCwCk0ZR1Rl/b
eVcs34l41X8XhAWXPwingf/LdSVbHXqRGT9Nd9EH2IVASmtUPueM0P+Hju4DwrRmONm7Qmr475am
JXMHoGt9HOW9jnoSa9daa778DrY/7yymmng9+OI7aNpLggspbvyjC73vNl/SY0/bGT99PTA2Bfmx
g9RN6JK8f4hm81taHS0PMBGqyIk2MrNjx3je7xMZFKuQdEsCRkIDlaMoqI4CK7OJw4TFHC8e+ZCQ
2FnDvuKsYWNnoOpcbM8vT4WJ3JCrmMuWBc+jb1+3jYxzAOvh/RF9gtlVU8k7zSLcZHsxBZQaA6hv
9ae4YAnlvy150IkJfv00Tweaw39HqZlJWoIUhJU2971oFa44CByCyLAuWE73F91/H1xjlfRNqKFh
RHwRJ5b49JdZiAX76DJAiiQHZLsInooAH5w4w6AEirPm8DdeYMDirW8qs/CFkRqldwsaE7C+MArO
rgkTOqRs5HitmhKMsJrZVTscfwzHNznKY9lUoFo9Qkj2ZXoJIwfLHCh93XNuXl8KopONONyyQ12M
pJdfmWCjRBQ7FUm6zv8PJHgObR0vN251KKW+ScOn2+2hpcwcDY30DeJvUxIqin1A9X89C/pBF589
Y09aKkps4kNUdOiqn756u73D91vVSahNcc4uYSjUCG5Jj2+/09j3XGsFmxlAYp09GQJgVc9vNys2
7YMnhPgBrv/Hp3xXumMob1ZTFNPkG2eSpQaqtdBR9PKTb+t98NguZqJYmPjBJOI8egTzDm7JsAtP
/WHVz7LTsmEMKjbrVUXwhiLcqBn/AWmTPe+rNa1nvKTP8djiI6YvgUuRtpaxhYP9QdtBcqJNuy7y
ijp49C6c3cP9rsBa6+4pHbymdrmh7vUNzf1W6yd40MlNGAU0eTOLOSQYvOuHkS2UU33Cr/nfHkK4
HKR8UGvUw+rZ4HL9cUFS9cpaAxTr9P0Kft2j6s2PznlsFxSGNeRI8NePsFzauwxUCqUProCCQkpC
FOQm7nBLrNr+u/WZGrecOHOd3cA3q73lmKqS5jgbIeXx4eKdSsBbkB2ceXlJIG4qPSaMJU+pFVZH
ekZdWqT+5zU/lNKLOtXnialZTs048o0n+cj/Oy5ycaUt7uLymVRNSJMzOu5sMlwnM5TEAeoFuHJ5
OAPALRawOmPtpdCqXKMhNBWiZpHfmyEToFI8Ys69OR7bTNz/ZmvTi7gvXldpb38b0cZe95h7DSsq
mMrOeqnzn/LDhWdI0aym2EzVif7Qp3e9VnvQSLNTHt/vzJb/TtSaCxTpufLot2y3EIewToF+/S49
Kt3+IEOtycFajoevKJw9Us+eueRFaetoY06/7JTSpQX8yhdfVL0OqfCmZ87UGRzHCX7xX7hu+GmS
PEGmgo+89DO6OC7AdTRghI8BstwEAXGDndrYork89g5D5hHYip+7BkauxrXxcfqhN+Hu1UMWQ+42
kQqym24cBDWtuBXfWTwVpR31yr4sMP4ZEh8nrl5v8e3zPK2q1aO4LOb7vGjKzeoH+ZbE59VW+Gg7
vSnhVdEofOtLlg2xVyO6yBWpBTz58JYyadMbAIbMWaKISn7ceyyrivjUTwPA6HzCznzKLYlXGd4U
IUcTNfJptONJflLHbdGLPKvkEc9Ow0hZw7fMFEk5M2Dc7Qa9OqeVd1FahiO1Yjsj7SkNA+x6cu0A
PkJIvQc87qCH1c5InyupQ5u2BEBO3ItjUrX1daJaL1f8ZUpQesRwXq+5fWJoIz6VDId2a0KYy+kb
OYGqiMFogIlRbTjygXmJFHLuFKq9GWM/pCDYi1ArW6G2vhX/SHvF8mU5MFQqKqkxaXBQi53EY5AG
7GB4d2W+LdGD4yLvoNL/b1w8+oMGn19cnkJvcXJO7XKmwOmYN0R2jISvZgOsL2OpwnH21ZxYXzpM
P+02n5rzbN0NXFHkEBajkrRvUhILdLtVhGoi6T+1E4sm4yYn3lbPQ5UUcH7KhaSyQpXxvjDSh8NF
fSSnkYE4xwOJ/Bs82dMHlTOcl1SmxycDTx+PtcL7ZgNZZvhkvlLuJsoTA1VpdkuE9vCQUZ0Zul8S
Kcm9xCoY7Cl3IOPGdaGCzbf8DnIzXCHoZ9jeD2mLyOSrjCOwbt0dIoETbUBGM7hGNSyYn29v949I
hmWl7+t9MTmur49RMd+LdhgJMyjifiICRj5FuBy3+7TaMBR3Mi7t6+CfDKuN3tDC2VaFjPblbSMX
FtLj/RT46MCOA3+XrDenr90Rn8StfqSy2MBbbKyBxwVmmUV9trRKkMC3+YnqR9DbxEpVedJjqqdr
YKk/gSgy1NdhedCZnY920VXpvjKG8/JY0q1WlovySaLjsvxXpiAxFG8IY7SvtWGdems5UtNAFJTl
iqPhJxk/gwydL55VBGhYs7rfMB09Wvh/NW46FIzclr8EV9tjP7voJZE82GzX/lJyuhKjPniD7naZ
LqQXj4SFUzXIBdBUjH67P4RGdfTV42GN58JAraMGIUJY9hWHx3ZBfovvmc5Wts0xB4L7jufRwWXq
kXGPhjsoV+zI61rEuETpQsOFEzKERQLh89JoCGmIjunFBcdJ/zDlXRF0gcO2iRCablv/fCUL6aIi
OYHuMclJXm9/EIi3GLyfieOHjx7M9NEEKIxrr8vylaEtEsoI+vMCpvK5ONts8COpmXjkb9PMB0Iw
P844pEAIaEw3BnqHT1+fuHDp27xFZqR6pTlcx489c7MAFA8tT85D0N/dqMcAFJGei6edzkGWyZe3
n3qrGOJyZLmFCYSCbbO4YmXyqVyfZgQ07aaaZZ3vD9uav7w3TWj5fjuLUdb9Iu2BAEQbdL0cIxCZ
zfZHn+/VeKtV9O0pNSOgEb/FMudIMEJw11eb+OsI6sAiUDr9HLqsCzqjbLfG8d85PdU6LRerp4Xk
U4Bbld5boJQ3YGA9F2DFDaPRPp5/MU4eCGWe4AB0ult0JcQxxWi/ZULYkCo5VO7RSfRvRGf5ffNw
Bqn5dUdlU+wVTpFeU8nyaJwXvkoGZ9DHQ37ltWChiPlG5RDswt7+oDrH81VtgcEKlaKMEQLL8GFy
zqOwBq0P0uhk+wNCFOD0c9gKaPOzSx8Lq8WrF616Yqo4JoZpOlEAohTNoKBUhUN1uvTnWnvxFxHa
Vbyg2zxKegYtJe3VWdZS+EwWAPi9cIi9Yx+0mITbCTi/ofasDnkvTzCWew8m3N/yfV1TozjLwjlt
/I6xQAiTRdE714kxcMJDFVQYOm3GLFLkT9GX6DFirMxX9vJqVBfn2vxuNXt9klJL4sclNxuOQb+S
3NKpBGZ06Af/okBsptcDrV1+ssBAVVZmbvKgWkxDkBB7uLTvYV8Lp6tDV94ks8ys4D5ecfVKipV2
oNws0vhh+6vpAoCfMVQ1720rJO5cA7ABCxcyqCMFuMrz1JSsyi7V3P0mJQ4tYuphYtqgG2XmNOV2
kG7NkI40uCpuFEnVeonXh0tpxQMFbSldfn2xiVe5VcthjI3sjBDE7GnPPZx+RBpTDeh9/jt1B2TS
DJZQ8snXCDHnUgOSIWIdko2tT1RrxDmsR2r5ZM5syiE7oab0+VRAGhC9vhwJYx2jqXRkYHJdOI05
ZMdk6pD8HbNxcRm5ouFf/MWdr6fBdgv4SBpRCxsLFzXebd+HhB05zd94UdiBmJXuBgBJUyXx4XTv
YnmsTUUvTFlRQWtdlqpWIACR8HPisWE1PAJHyU6QiMWhrB28TdHpO4soyTq1dYrTMEhoGhg6Zg1/
ooF3OC0MdehYuimfRy700d0nQjZ/mEhOzP/Xk+5T+bZPbo2T5oz9zeyTn6fuu/lfCHiFnNTMAKGS
OApDTeeK0E0Ilu7J/F4F01k0vgv4NvMRB3UNd1pVtVwqV+zNN5ltH8uF9lvBOgBQrzt/2po+iUaN
w00Ha0Sp6VmFOl3ZKPnDY67k6L4QhzcXgc6yKUIZzf+NuWmD4kzcudjnLus5fsFpjXqRAfCBdlEU
nN2ncgAT9YaZttyVSzIsG5cGRaCSjLcHRxIG9cBuDK4lvmM489//U24ZIdFDqD5gyfuGrApDqQ0d
f1JXKMx0Y0kdwf/kBDFgLCItLOuGz2mjlbZzTiigFEiUH9Ga8Ti/7zR+oWGv6DzAH4IQ2onvAFJN
GrJRTcvq4GDey1MMbzVsuezwPdOyNyYDzRSWJ72FRmjOyBzDOdyaK11yyWcIqrmVByCf6KSfofd9
eahiSYdz8gHaFr0A4DLlFHSpnXAsvc0K+ARGoaSuFvv/Zc1G0LCO/yQcEsAvcPLhcp13yzJ2KpKD
OOtSgVaGiykac/3AG8XX2EhI4IL5ktOz67/RpTBfrQ3U5SZcOYZ3zN72yPkl5gYvrmbCjXZ+nFqA
mtsQcHzZTHWscDG1edIgo3Lzm/1CmPle2dkMu2DPt0NTzzaxgMdCTh6U/HFrNsRtuxBkQaWQtJcm
GvajJ9N/Sug/dE8BJOuqXMK5CYLLlNEvP6Kg/IZDoCame0qbDK7sHRGbxNH25c0ubAq76UADW75Y
9XpnRIct2CQ6+WEBiu7XTSRwQ7AWj+uWSR6wIPG2W4k8fXaNR1rCoHm3ZgVjm6METGSrGtpqqbXG
bFAtPzgByw+Ni3ErtnLsmRL2UAB/XCFX6abLV0CIo2HrrfnoKr0b4P0joPzRaCO6D07EMxzGqDwW
Ihqt1afZGNZYEU641zuffJiw8k3ZtV2XKtNEJixMMGdGqx0CIGFuxBlu6eZ3k+mgf6iDHfxxE9Kr
ZuzTDVZFpcub6Hl1z+7ulQ/fSML6UkGT3lrjpRJMxoyTwto6vx0WI0e8Z5asX+3qvn/m5t5lJmmp
tpdNCQkmxo3hocgikRVVKhWqp6j0Sb8YKMImraYAH33qgGwD3uFr8zpdGqFQ9gWkeHyf/ssKXSnQ
mdcDPfovL81+nw0SgmU85BK71KnPduryDw4xfgE9Bo5jAJyt7By+gFRResT5h8M1jZNzxKmADL9e
xw2UIhuiSjDEzttlTRQOLpCtVrbukbW4PB3w7QSIJNN+4fDRXekvBCpiAe/zwaqE7pBrnxWn9m4t
w4X+kpvbOxmIsxtaCtwPSc40cep9fPFlvEYg5hWSb+oLdrqW0zetvJ72nIiU5OfZHTJpFHXwqjiD
nN2P3GXr0MAJabbTPwinFjJ/SkKAC7FyZwLrb4zf63fjyhqwk0aOicSHmLEpz0A3sa/So1YFiuBN
nX/102Ri7k23RE16e/WZb6zdKv9OyyDVePiUuMEHpIWGDwSK5iqS5rKjC5topFHAcOQZMF1I0bZm
Ai2S2nvOZX9oWRwR8eenVJi058DoAVpPdEJr66c2Url10Rc25kNGdwKfUOKiDAAJkdInDkVQ32N1
ERnGB3PbDIoAwwrRepzpBjJ/BY+f0+GYvtscXOQYmqM/ppE7ydDsoGgjgj3STeRxeFX4IiAfh0jc
VMXPvRyPbZZ6LfQwlL+BNm9LXF/lIE8aAGxW0J/++ijd3lTn+jaZJN9vCc7uJuk+9O4Oymxw+jXJ
gF1uMMf2aaVLZdmpiK2llknpxIEQ7/74StqIy/YvUOpW7bMy+VbedXW9ZeOpZLJvp8yqk6uwKTtD
EiICEa9mJIs9VNtIywQ+sIgXU6wPsP0/Gs5WPoIXfAOm18G4IwtOWL9Tr4lAY9wm8M6ba3QPUlHc
jZL+PuCHFOhtY+0u2ceA+zCFvH2hYgwGc0j1p1zADet0Ehws3z7HjTECCESdfCpGYWTTvT1HPGoi
KJZGvV7ac3pvW+y8AT7tT0hI5KA2cAvOoOFOV+n/7w53stTaaELhHp9EEihyMJl00dQrXNiIERTv
SsLvW1U8LeeKGMYCqJxK5gr1l2Of6OyRHs30FeCM0C8gMe/jgm1endvxHNc/s3wtcMp/evqvnPRe
lnrKMWdQD+IETDT8/OGs0T3zCXW4TW7d+SOFh1wTJ3m026TCFnDLfl3RNSyrY+ZyvcjvMqvuOGSN
8P4+8/crjZOAiKmILB/h9ZNhSYHLC6AVKPO/GLDa2+WhrG87nc+0wbrQ9SYveuNVUcph6VxEJdIu
Jua1EZ864qpuS0hURugV5/Icl2zsOtpJj5pMqQ1MHxGFlZdvCMB7QOoLfdBTdcBUdBdFG8eIli5g
tI2LmQvh+zb++R4AdzyRSxVM069bCWay9bPHw6/hc69fMPkFE4NcH9AuIo22J/bdN0Adfaub1IKi
zh6BdSJbPzzlDg+j0BUCS1D7crK8ykPs8SA6PjKB0owVQA8phrKRregnTsu/06ZZ+ofQ0vvcDbBy
kxtIssSHoaEP7m/0IO1DCD3oFgAhdCadKrT9jGb2apVHLXaJrZnFu3ssjX97LXSmGr/D1V1t2p+/
q0Ii5RCDyR5LITCjKJn6WBioq/nb1Hhq/GwhbjRA5F1owoDDi+R66pMitV1+uo+RF/bJHdjkbIVb
Yer02/zJSMsdqaxryHehSDkwaIsDIncuPrPmsVSyxrs4k4YhdxAcvdevmoanY3o/ZFLucIr0WKSZ
eT591PgG6RJXvuqJiKilEKOyD5SluYFH+jpUyF3XgLbfS40D3doZf66+Wsz2dxe6EiwU8dVRRSeO
xA52BjqFvzy4koICrijBaDPXOs4FGaaGef0Iq6rDbHGlmg+PE3IxPTWFJN35HMl0uK7eQWZT4MVU
kSh+GCgCNdLTH6BEKVogw0heMb3bppdoXTh/ISzi4hyze6MUiwVJMJKK70T3xIrkbRelXAUisImo
He/n6C8OEjK7pQrqVUNQb5cWo84YHJhhQgTKuza/H285ieqfBE0Ns3FLhhxKev8n/bD2JaIpTw8K
bPry5Gzk8EoiVdih+krlI6q6sCw20cxnP4HHRfzxsIiTI9NM3Cl5wwH109JXnsEtuBwetFCI49pu
9LlfcorkplA7F7tx7NLNihElRq+w8VRPSdyKmO8hCBDjAa6KvrR7VN94XG2XxSx8/HRwrLGO4eJz
O6GsMaCCwTnOzSicOA6kfaZQro8OAyovBC3e4c24zutyork8Owog7DrQ61Tre/bxLnSQ2HTMZCfe
yR7KD9IpIDeESNpuX9VjFcssrgOdxwfDeGCAZpkQSg5ffaVRIPSRWJTwbC4NNqmYbuLAXmqWaIzr
UKgo2pcEFQoXB1ponUz+9f95BnM+alMo4HaSGo5NO3EnmNIxdVW5pwrJUQ9Cq70v4eBQdI8BVqPM
7tFRR8X2jyNm/ZHscd+fhCUh2XJJbP30szY+aKWCzzp0tWi57GVsIoZXV7Jaur4EJxkaBizO17zq
UZ5OxviHTq5URDHtmXT0AUEp6SlMgl04e9i/8Vrwxi0mOQLe29Cn3p4A610VLNNYSZT5/LC/DTuA
F98xyvluXbhPeSuADX6gTTNwpJdvTgFRT3l8RTjG4r2Ix8K+9nc1ACYPL/mWU+g05tW0+NH8Ynfq
Y82ocDZFlFIG73xhwr0gx2SduB+knMZW//MGiOEQq3iinDfEVkGyPAjHdG/Q+q/Q0oCUWlTSdHWH
18Qg1OQjTxJH93rqVlw7+PFI0sz0FtQJGod0rP8k38SRu+BRnxfF5AU0CQWEByZE+BbKN+BZ0HvE
O4Qjz07NvjUw7Z3P3J4DQle3GemcKx5r19Azwi6eC4N5ADwSpRjWc+01OjBWO1ecJvEUoSHWaQjW
tVhw7JuD2z7WlEtppi4C2xdgsxTsWbW9kzmisNba4VKAaUanx2A7WlRSDCPOzc8x6cLUnLRQSxWa
A0P3HqTwTlsz4wBjL+Enikv/0Tte2pSVwdJubZVfB6d1a63Sq6++lbqx9UVYJelMx3wcfzejSYb6
9eVyxUPFkafCFyPiJJzI/sdJ6kUsK1XCW91ZCiSRMif3/Vz3NyN5Dh7VPt/V63Kx5aT4Vz3LNIq1
kMhFRcKtY3cMpEd7T+p2y+G0xxTaqYzxxrell+29btbPnas6pYC6tpqUVnf+elRrb6OjWMTL0zHT
Nnbuv5pGzEPb/GUsVwKNeWbPajPwTbmPQ92b+ok4nDjWhXtZMwK61e+6j+bl3okSihvpV8Jg+IOR
L7tkKrU/tVScdCQKysj+r3ReSNgJTf1Kp4uqWu4mmXbVaA5XX5MsmxfNS+ii9urCWTTXfXuD/4oX
ueekPlTgXjFzIa8CbY3yhAb9xPJZvcGBrxMGbmKawQjP2XO63PWOeeR4PC0S+sROzRZKrA8iZPY6
3R2tOFEX3OcoKjVPOCzMzI0tGq8AukFS+/z1i3WHF5v8s7joOHcpdzGGn4HBK/ilC+1WfSvTiPCT
2je3oCt16iltz2qmLVKYHutUgzrLoAypdCPc6IJt3IkGBUWjPYuP6vKd6lVRvM//dVg/IPPt21d5
9EH7TN9Bvtt544g6S4OdSPSWmuqj5oFZsHzDF7vgQ2hLUb7yC/QlckqBCl72l95FaqAKqoVgrGBt
VF2Nw7HbeBI6J43aEIClbmj24quPZcd9KUYRCrQ9JfV2j3LmrmC6sHonPhY/x5LjopLRiwTuH3cP
2zuEj4wepp7k5/PUbHKaTTbiLS0cAit/DuNMpf5pcxbXwEPpglappjmyFXwgwbpUtO4JZ9Z4iD7T
mOnPjLr5aIqObIjveZ6s3H7+FbvNGWydc2oU+ntROGaxySmNxPZ9yNuVlDmon3qTdlkBDge4vPWJ
4+RZz8yjrVIyICzf8fDlgoAAPd8PxOIOzLFUcSmpyNfyVYcmVBvfJ2qaYcRIb3/ecjpoZKumI/WV
5DmdAJZ8xnWviOd4+Yv3+XCWbJcCO6x25tm9xf8tQxhIYZiEutJcGQVxOGodHa1koFt9s8QkzZQ8
ZGC8ecH4/E8bj5C+cON0Q9WdqarTFQMKiTg5mBdac/KHB1xfhZZ3rdPCpDn81I9XPzXTr+QszS/V
jJrROwvnQW0Bn5PV8weE5uGvegGRIuQRFD8t/jVMSdGlV93DrarTVQT1epUO1fJl1lDXmR1mOboh
eljHNc5I1QruNUBGfkrqyDohxtLGb601OH5lPXHJNvLp27G8PqifOM78OWdM1Q62Lcqs9rHJEnUw
MT1tMwFlIYDtJmmiJdNCmNH7XMujrXFRnWn7AHNP7T8U1PwcSgzz1w4RHJRnqGTqwTpGmtMO+bRp
7dcMQAUlr3uaE76StWTh8KJXgJozGTQCXIv4bxO2RgOVses+hRsA1C6W2oAPoRhgXjpqGmqh9BQO
W/wr7DXVZ2TbQFWSr58SZIWS2FF5Yny29rZbetSUxN79xbQq1vqrr2bV5JS1mdWE6tJ3Vw5Fvn0/
haWW51pzxcIJAnEyXajZTR14SNITZPoBPnnFKmWaN7bWT3JY/vDDcaWm89Ek/l0QjnX65GVYE5Ps
VTi0mw9Q6E88NpE3l4HAkRIjYRndFqTf9PH6OdompjgrUSQTUoZG1sC4KQikPLgR4FWKCdSWMkVW
kTwvCINZP8yE0t6S87B4/rUmFTvqVpbmce9T2ZdoxfVLnXRn+a7KOWe3QFcYidH83DX3wPQ1j5Cw
MytcHlkBGgRjFNMt+BKP7yKfwSp7SBYi0DaQLaOUE1lnXzl4Z8dMZkVUB8CsYUEmpRjDvUealVlq
/o9o1j3w6UIcwNgFMATZkOJzrXlhyPwDexynnkf7FbxaUtnny5SBXe9VQ0IgeK+AnTXZK5WfwDSP
DTWXLPH3zmUanbYIA0R8N2NxnKwbyPPv/WReVY0d06DzMKOKnhPdsj1MdqxzEO1lK5lgmsEAY1yk
/ZoCUJnykuHqHA0jmx0Y1bsblD7VhV2L5EGqWDbhAs9XTQdNgKpPqobRdsujcTXft98U++5AzVFD
waWGLof0JT5VMPOq8ybI/ACgU/wHvgaQC0mlQpchzW2IpedEx186dHcW+W84IK3aYNedItovl36W
DOZc3GtGggvvUPQk4Uy9qEguaDcotqG/NunblN+3xw14y+ZRoS145x+TbsaMD5YI5IxFyqDEQmSx
FrZyvL++66sCMuzgoB4gWjj0bhkU1rEKDUJ/CaCH2eT1jgoTk1grx3QUqJWyDRhGtPRb77COBS6I
4yxCpX20xreXH3mlS4zsVNeq1ApNZrNO4/bvR9tyjparcPYt/LX7WEUxpwKCbnuqNyX5I6llY2tQ
IyV5cqZXt/NUXr6NY+qQzeAWY48DOHl0vaAbmKitq68N1EdmLmUmJGqQ91duR8xUpTIz+nBDyAOj
pvwdWMm23QSNuvmQR3zN/ZYnnUtHir6virbeti/tC0WG1FQRXNY0wrRxNmzqW1jm1bABKF3mguMF
mFrzpN44gtw163Wflm809cQTNkNIGcEI+U1GL4QWCoICPIdPMXhwZ8pm62JhZAZ+FLEQ8Ih0/iqB
/UeBgDdz56ZE4sr1pkpxFkpdwTtgTiAbvhr+xNuzT7SjjpdtiUO7a5CGYV7/CW0R+gubDBv7se7O
ZtT8xL+9voc+7pa5YjNOsyCnP00mIW7pNJSZw38J0M9if7d8YHZwBZoYFHR9vRASJ2XfOdCjiEla
PbjbTNFTjTEatnLhAc97iHXVAQOYzEZKc6xDzP9AejJfvjlLh8z4ZhsUpZTVW+R8xk8fJ4Nq1dxP
gdBEKvrx4xMnNPE6BcJfJyYM/ohHqXoLcSU6AomTNcm/+hinptizB8SPQo2+2jmHBIF9/7wcIF6F
kmuHw2kdFsYovMWGUOY3q8JOgbmEa9uUXymhCjC6fj6f/RFAzDKLsX/swJxG2rd3YdamSjnqgPJR
ZYjkoIV/PTI+r9aTuaTioqNnsDn5EgbmHAm15HeFgGevZvzhBZX08ZwlRWQcZWMcWvFZvd9+dPX9
UNxNCq14oKOvHDmMxoOdusbXf2JhZmjo4Vs/bRB9w/EoxO0YArxULvcULBc0PYJK3bI6Aod918eJ
aehhSZcI//q2vFHW4oOh5Iewjqd+ZYbT66NQqVj7riBdtcFUSPTXhMX+WN9unQ9BvI4dGk6ZIPkL
7ik/GVL9+HqefFpJ+YvKYErKRQjRLfflictW6eGELcnEezYixBEononczDWYjtz8Vpk9XKHr3YO6
RGTxsrU3A6PBhk0ANzELmjOXjAONyNxzPd1rMrqb08RvgcbbvPjexZ8r9LkxUpqKGHLxuBnoQUkq
2zEXN9hPJXjq/HCuWpSD5JODYXZfoqPBBCsK7z7o/hnQ3oQ+hVpUbvYMvHkzWeMIyaQIYYG3LMKX
vSUHbBqWyz0ZO8hpmSEx8dfbOSyM44iQw8SdtbXqkMJQaqaG4HfI3OGmkyKC66M/mkhfp5yocBnl
P4tY3Ao6HKaGnYdvNKMlpusANrpqsVFA6DQtFQqL2/aSCkOgKUckLneXFvaqyEBDlulPqp/7TiDS
PcrPSH6fMZUdUctAgvETqEiZD9ySgLOdo2yzDtlJBIPnhzAWZwQPCYqafOa2sZ8uq2MqGfW1rf+1
9POyV5oConEkc/3MaFqwy5gTAnkRDqOEdiqncNobfNE0qyri9bnlFWHJL9v485H7deN0ZIBFYmPy
QhVlQxtWt4Jp2Tp2+R7BIWbEnccEXRMoZLsYX0MsvdCbXtAcE+OcIWzpUC1W2RkJyesSeXLfnYNP
0IO5CEQflb8gDpaGbjs8On+BD5j0LODhp6wkcxIxWMRzxZYQ8BPvTUCrhCisLsTv/9uV3VTsbHLJ
jYjkYqTzKv8WopTF50slhViubADWMW8A/St5YNkaZilDbOQCADry84DIoPPDZVi7TCioQF8pvfr5
V1MVkZHHK79M/gVaKmCZfZwV2lctxXB/oeXGMshYUt7Xh7BDEDm8gem8C2oI9rqkjdzHRUhJi32K
r3x9dSlvWgI9cgiFKv/huX696hcKbkwAuj3jnZlEUEK2iwZx7PZ7HSTGnXT5A6ZHhcn4rrVHSrjJ
ouf+k+/IWHK+TipXo+FpBz9Eo/b7aNSBBwAJOG4zkBLxak4pGv6aFzgkkhilv+fZ5n44weaFiUaF
+D9XlC0xWaMBeeKYt/aR42rTYskQSoQmu+0X4h3Og4WPyY8cG3DtD8zYoK3ilNrwxS/o7BIr4RlI
1OK58FJJuBeRbbGe5xrncoYMJCzUCzsEMzJyGLj6oJtQkK5s6TIfuhE1RcT+ujcA9IKhpird49Bk
slCZKDDBE6IxHkjk6Iy8ENHfZjYf6HwQnWF7ie1QxLzmfpzvL+mI4jiaR6/1QaMRkPGZouoHf3qg
o4ykjF7/QpYkpvRhgOPlpm63ZCSzBhRDAMHFy5d2yKW006IuefKvjBAcqCu15UJMmONAqokLjJ7p
HtVQDDfKmPAnkGy1M834P61QT37YBtmJy/sqjChKz/xsYn47A1CM+F7N7qqsD1azJTea5WLrXwgk
TPmsWb67kGdj0eXOjX3k6nlc9/qzjXZq8YexmfiZMvRR9JiIVp3B60FHJ5yY8rYu56/JkxTmvLlD
wJIDl6koVNIXTfbsKQP+AV9PVRaEdgNlRmV0Rl0U3tHuL7ObcbDfnYP3rit3iutU4oYpeDNj11e6
/4NyBIlFS6NPf4cDlYuKwbtPa3t/+4AQYJgGC6FJy8FoDmwGOqdnfozsxXx3HqqE6gf4XHlTKqHd
/4uq17mOLoMMYnti+ma5tU7rvqik0ORgwIzktDyjywQXpf09qhhzDTQm2BUTGkjCgkD4Ay8mj1iL
WYXdJpm4DJ5vLRXjQtiMizBLFawwFW7+sKiDCKA+liC43BJnPktq9xR6074NKAnNOgDcA5a7CuWC
sLC9W11zAORCmEaabr6epMilb9+wMkpnHoNyVn2RhJOyFDWgkApOXRJIObn4QHqC408LPyGqPsPl
0OFXbAG1/uj10xZC2edTMAMd+Zr+Kgj3EiYMkFwg4TQVKKc33pT12JvkTq1vcEFugxKJeW72BoPV
7ebwqsaworP999308Uws554jbWexho3DWKShNh6cWfKUx0+WJUW2NX9g2Tx4Dx+BOJsAzB3PrGhV
HNEPbhSLN2itlN5Ezn9eitq456z1v/PEMFZrDzxH3WcJk0blvyEGsHU0HLiAlmfDaWFcze6bRoLO
b9WBMToUPs1tgRoiyOdRlMBJ7RQgHmY1U7nLM3JJyrWyfW6E0Z4Qk1CEwUOr4uasu7+KHVoenxVn
M3uNRi7QYHbBs00Lyb9iwaW7uX3nnw0edKMn/N3KXAQDiF2YMqldzwTQdS5avMW9CJvBIVX7yr7B
Z1zZQJHbrCgx+1PDTUGp0LBTSwsqY8ktJgNnnNSbf6/1QM3Y0I4oAdQM040cRxWW8BSUVl/Z81vM
q46rtf22nr8LpFWLPjLNq3E9zh9RsEOtIgc00f8MzI32hYVtro+HtxD4UWVqYs0BMuzAQIgLpUqg
6Efs15bM8LvJsXtr+fNEXSYQ8eUhyuTWOEc8GqOqqYG0nByMKy6YS8TdVvI2ueo/Hmx8hFLQaHjb
U3a2ozvv4wI5Vc+uRo0CTNC0VhHJJWPPGnDd8fhJ7e7Ps22FvL0pQGuS0gNY9kdlPhzx0oFHzobw
9Y1Mw5s3bPA4vAkLkqm5RUYsYIGQCxcMBsgbXXh/aOX3oP25nUW35a6Ye704n77+JVq/yAGRWAEy
lGtUgUBo3+HuAm2fsVIm1cwWXjO1VkrwR/8DCurZ6+Vpjjxy8FRQDPwab4+iENSM+NZFO14YS2aV
S2VV/csSLHXDl0Ps3GIswfdCSX+BKOFvruw9X04BZUgRD4Fkr0j6yQZsxyDHAODT/NzYJMLeIxBU
/R13l/LPOZzqRxA49ie+7CHjqGgx+JYBspvbqLj72ORQdcqDpSpk3MK8+iGiDlE8MDWa7w/QAXeO
60IdvfWFy+9A8DAt+JicMZfT4EQxHs13OszLI+ysxkD/XOAdCVPrmyCJmoPM/LKYWTD21lPY5iSC
lZSp249m/hOyAHTSdVCIRo6P7u+WEKBOXhboC70g86XEzi+BqJD3fNr/jjMSEFf5Xofvu3lFMjSs
OD9OjBqjGiBnIpR/ylpgJpbm0NzEghQIA1/qczLD5LdCTBV9JffzKwhNFcNvFxGJSC77tE7TbJwx
QtRV2I4HSj4fg2i8wSDLbLWVfZ+C2dkFrKHXF9xbkEiSk6lUZc+weEAR3Qh1SzDhysv3LlB/2iUw
dIfiXXiMEyZYJ2gND+TNBJVRPUj16Uos8rT9szirRzotnroOWCToddF0iOOfB3sgIhM5lavJeZ1+
I8LGA8iKqCZUi9uTB5jesUhk7ax8SUw5K5cJ8xZ1a2a6XKJXYx1b/7rEwXbzViAloP/vb/SaviVx
T1MqAH0tT9lyNatTvavzT2HmT5KbC+yL5eelWRAzlOpewE6Z5XgrWLhtnPsKyqMixGWFlrxQl9V+
B3c3XUPwhxp48E9CCdTQd+WY3LYo3R/IdPw0F+k3wWdVY465hbd6BPfv+xbOiVpxpfB9reKzO3jf
GwowzxbnaFxYvVGcXWIvl/QMyNtxRK52sY2rLFlLkoN6nqy0KBz2iNM3NQaSvv/eaIXAzK/N8YD9
PgRasXA9vlnVRkwWFZKk0c6xYnSo3IKBeRYvOBGcN+iSrr76PX/zBGjaGvuS4fCxz6+zAP8hi6D7
UT/Jystkf5TFJPOMRGFy62omAvZ4tkPHOvROYrg0mMlB9BpxsjbTqlxTKEMZMr1S18RbvYoQ6ol5
9veW1OwDnE4gSDu4QdLLSFH3V0gOkTxRsPBXfoU4WatIToRefkWE6zQIQjOv8rqN68sMqHm5t20b
ONTQw0clbdw4yCat3xl0QEd7bb/2a6PNg7f5+qIS+4mZMA2pYyrvh3gz09kePglaQscWBO8r3EZW
OAvnaUHYVVFrmXdzDpO1VETQMvGjiIFLdm8ItjdeQb1s5sfwkfiDwkjzNeAEOi9zBLLUPGt/LaYD
zTW/3ZP2gjerrjXTO7ccEb/6WEkdlT49lSSzYawH3vzA+3k0tj2BqmFsW8jApu2n9+NymT7FuvYl
MYvuzuaeSKtTxhLWin3cptwRFZh9FTEkf4/sXGtTlKzPvl7bMXIN90ZBuQ2ME/lc30NKI3FqJiG7
GbWes0/VdVlFE4ucfSe9BDdNIyWefVcr3tPuqnV/C3tI2uSE+PTM2u2bGtfj6+YS27nkZUDyzn+u
ZRsywGTxqWIhqvRFj/i964Lh05wNbkyHcXVSff6KkA9J/gh1aNC6KwzNniiCOhQpDZQez5cpxZll
z3EBNuUacVIU32TlHfkNMnYaoJuvl6fXaMoqrn9qO7SBVk/n557F7awcs0yEiT5c6mT5ZKxw4zmm
P63rqK9QKjA9SK7jAZWzzjz2/vrybhnMl+znmcvtaeEot+5P/t29V6V8CKPsB1zHcLZLYJW4CwtJ
Byx1VxgYM065Nke8e198E6WxYjm7IyxrxP4iK0dKTvMastaDDRec/qGmMUJ8xXgxjSjrLwuYUaJY
o8FQPx1JHNW5bqE5TyvhjDCD280M697SyOAepBK/5BCrDy7NAb4vK57doXJtqTABWgGaDApxT1z/
/lMhewHaLgKsUZ3Xga2lYvouuaDwUDA3ZRbAe3I2WUTgdkXOYDWxapIpKsf0XifvthqW1b5JVFCo
e4zokNhIGsqmCthbuo9aPuZF8/dR8QYGJSzLqaO2W9u2x4zmyRuzopwyd3nYZUshw/aU7QgbNcVS
Wy4XBkC5wfd+HnmesaZym4TAheOe8tozAL8dkCOlUMgSJwXRd96sRP+Dmiiwrt9FwOdt2hF0BdHC
VSfVriCsx9BC1VMfy/HUx4YpXGFl3zLkfr8qudD3M7/6ISwaezgYdExUHrU3cIgZVIFEaXWFHfJX
NiodMrj0998gGx2yIvsQPTvssM2ytIrPe7SWAAv8JCSY3GBvfs8N8QFDt0ZwXhVIpZrqiPz1LFXQ
Zw5Hit2SmqNcDGs92P3pLiVWjAvVkCmpH1DsQ4Qbr9gQ/Gf5TVDRaFG01k/s0tIpCOli/xF31D+v
cYvf59G4qYzUQUwEwQ4iXK2A50QPDJe50vU5pQliEJo1ZiZtpbGVTkut94ylS/sVi/fVmEScoL0I
VBG2gZyU91Rzmfcz6i5Gd2j4EAw0dlxjX4GGq9gYpwnbN8flr/JMlfkiaPp6TDXuLCcSucfQqguX
b2XCPV9tiMPyL/RVh1bkcKGrhR1v7lnKDEC/1eIXpXh0shv6hg+6r8C9oK2rqdR8ZDK6JfAsR2K2
r5W2WzDWZhOXwfax3TaWSTl3YX0xiLWbWp39z0pwvr3d9qPa0tVWIRqfprATJhWNCycKppzWGvgk
ObmpN81VovwnDOHmQc6nzjUx9ECNU3c2UT7TKO1ECqIzkFO442xr6Q74nRAxNvTK+fafCI49DMiq
cLAQnRLq3yr+p1eO2pcSSYbCYtizsyXNiZa52XAV9W5svDSMvb8MhoB5+PoznpfZIZRltkYgH60u
J0WWZudpjtVH5LmwVo3MwQqufqk/hxIKpwVYbbdc8z7oshPq3IvgY2H5fl/Rt4YgpWGbBcei9bqq
zjq8Kj/ZnZKNGMw14yArZKt61PbzmuE3YVeGb6TZiW6QkcMJVLQsFMzRzCReGg0XFnClgdT4FHO+
ypaAC5FG02m136rXLUqUU9Kh2fhZGe2Bp0n0WyEK0g2gJpEq1lYHW1XLY9KrVR7D3pQvkc3WrPo0
dqWMFoUY+3oZvD++My72LI9vtQd6bFCyJZ1fHWM7vtTdnVDC6Mj8Tjb4WEFCUiPkwPdMkeRzNXJP
tVZBoz0EPfT5yZRyWu+yCRsP6qZUmhbpTfTy5r4p2asEhg6W66J8y2sv6SrszcKazfGiTyX71rv7
YHkVTMpq0SFCAk5W5Iswt6T+41+hMi2T5HfbpPYbnhL6hPyYZ9kFO2GW0TzpJuuTPM9Zun8EJZwC
yGw6TE0uJab+r44x0dSgNWODNrz4geUx8MmzQfsNIp7M+64UTQd0qIXYr1nQwYqaVCpjGBnFpZLA
5JsfJU/6tQzDXGFMW4AkrDYhVDF2oNFi2R9ifoAp7xl2eZjPEn9jBZuCW17cRqpK2lTT9ZqUh9AY
zc9J10KH+qrPms4p3PDuv1+ZgMq2OuXfN7O1z01gc4mbDDT+0t0t6VZyRpFLIRpiWoo9kycb7fQ1
KrK8KU8XaSBlQrOOAHXLwOgXY6fdunihIY4a8B78AxWAFHPlBZug3OhFBFsd4rmWoNGexBiUEYYp
dF9jCTJkLdOYETSiKVh0oF62nPbm2jWkwZvb+rwhILcgtzYMaJ1V+oQZxMtAyQ343TkJuMBsM7yV
QxVyemMrq9BE9etHyWHmMNNKKm1RYPFB5C7WBGpp7kMjio5K3qCn0PxFo/qJ5CTi9it3pB1fvDpa
PPsfcq9o2OKaMFZP/7wKOLw2mqJwZSsK/QeD2tmC4TmsSIjRUnO15AZa/VN0r4D8DtW/IvZSlPug
ofked5IeaWtRWFw/ytjMcN11oUH86cC1x+ARweMxa5w/NxDfFifMbydnGFVnBfX9LvO5/cClWHng
kt84cmKqcZ5g4OlATh/KnmwpFb/8dX/IO4HcK7l0lMNWPxC8/2buSqv48/bXlMmApHvc3KZIrzBt
p3ZuUyu5bCzHv1dATQkyl+dy5f5FAWkah9vsCcLZodrIDJ0ku2EMW/OJHKSNBhggZIWlPSumJBiY
9bzCQlSWwt0hS606MzkNRqQgDeQ3bn5u950y6SGFAaBbCMKdAZrUoji1JfTXYfMFcTs3xFThS0Iv
NyeXVSlLrZJXaB5yEcN2I2pLz+jfwd8PKcfwjPq/inLsSA1qouY9674x9VClZkXcrNMpVIKDNcwO
WsgXy3w8DgmmMIvGGrGwCbU1LbS5Ya1z4lBxEpQ3SxtVSs5LCYURcdOu5bjkdBovHM2GpT0DQUBd
Q9L30mroCKt3YJpXHpcr4Wvmu1nQhahT5koGngCOc3RNOF9GCP30DkDx2ZOtn8xVm2BQ2uMM8G4Z
WQYBl2XMRIK2k4aRLgJrQZLc7cI88riPwv8LddKf/A0swbjB8VZVFR3vO4Ac3kfA7Rnzj5wra8JX
p24kAZf6U3XvLW2+9+PudtGKNR/R4DiHAFbTBFlDXCL0o7solCsFEsdBYjQx2lvxKeEDZx1B1SY5
XBumgyMn0ZU7VgNRi0xhhe13bQnJHvVYQirtJ/CzjvsHYLx2UPl7eQh2+Jx85H36N3MYPRQFy2C/
lKp1uqxyd/5jF0DlROal4T4PEWsNlSv0hf5efExV41XpV52BM7nKMXpCAJ24OrFVnKHtkg0y1vHc
mn0PscovuT/cLIauoXHgE+hRxjiUNU+J3GbPBelrk3mFIDARJePlcIqGEPv7KOT1DxSClyOeCAfC
d7zo9EdlIUbntMgHMENnjwZMO/OoFXRngBvgKzcZHisyvvFBBfv3B0/m3S77hAwrDJ6rSIdeKP6y
AUNnEBhNpGuAMpNbRhK7gL3p5Y9ADihfzXh1F2ylsRjjlD9QwMPVyCnwQpCTu9jBBqGdT3VH630R
L8vPcbcCGtV2vY12QiFAVkKpaRK7FgPGvNn19iO+DXtfXPu85M9rmx13xxwtnjO3vDQ86goaP3XP
Wh2yAFOFs5/Xj+hgHWxaHKPAoccYQHeM9TlbaNqEXzS+ZkfKYrRwv9mPDU+qOPaFW4RCbnJuASfk
eVhdIETKan3xjsHIe7ZjQJJdsbKcS6+wvg+EFZ0MghmQEkkPIhBt8v1UklSodxckReTDaJCZd0lW
nHaN8GstL/tSEfoqIu2e1AB7l2dcz+efQPRHpFuKm3ViCK0sxB/NE5B0N6Ree0C5a9Lhoe8QGZxB
aYwcYZI6va2nVoD47vxRlGi/axcB7SqhxDW0vIxDErcjTCgnDvPgde+y9YoOIQmUTndsvKvMd5ry
bDj/GiVtWRLe3qGojm9t6fXnHDCvxICFESRGA4sWaprBtzOxym9ElUqS0Sr6vrKfHwjrmtPGDImZ
yaRcLvNic4ulUkcGsboMb3GDZ8w8silrwx0PR2XbFacsy/jH4591fG2ZQf6aL0spRe6FHiif5jCH
+ZFEXC9mbF7rBF6OziJ4L08M9JLZ+tYe+5rKfLMw9g/NeZ8PtmMylosIODem+ydOaUjuDUP7Hery
g7E2ZV2SuLxeCiEmkmRJutjZugRmkpwywc+HSbTxwVfNx5SeLs9opW0moBMMT9XkqFfSEYQhZj3S
uGAM+Kvvwe/WkiPze1kECaMG2OErR4jCJDh9Ys6tayRaeYAJOQbniGsQOT5Y8ye+vVrLkkZKw+IM
nj5j02rzlrtxONhEXTun53xJM8eh4Glu3xukA366uxTHhEgU3oRLRuNk58+N9Xt/J+xrvVXt8HMZ
cTbLl8jbfUX9LcgAwzytuo9htnPt6gkGGKnSmDARoWabUpYG+4jAwO8Pj0tx849/9QGSD3m7Ih4N
qYAJFomC0dEho936WMV6qphMUU1iEO0BPxfYPcPh2VY6exjOG9uOjF6xU6KD8txSDo7p+vZCNIzI
sKzjZLJTBsCE+BXC9FaDHVMPLJsyoIyYeMQDCRlFOXrDRVC9kFzzLsJfrhrIpabnVnunobzpP7GX
6HlKdHUFKA4ZN1tIaEHrzN3KFi4rfRopkHMYnEwuiQmkIfzKjLkY+BvjSDo96CD26Z8P6hwwZnYK
b3az652INiQbnAtbfHTRA3BQDLIsy9AwZEPV5m3XB946eZxASazeFvl6ZbGPoAwfKXcQ+Ds6FG4q
30aOM7NCiTsg7bpoAGH2oS4mzmKXCJMPpxoS4hKtiNMtMuL7l+mYK+WB4mPLVA6o+1tbS7ocGsRh
dBTSVGsuGFHjK0hF21xK8iNYJjaKv+qG8kaUYkycndB4r2+qynU+3/XdbGdIgeG+mbNPsvCr98qX
gdNjt00vQ8U3Tl16L3Mhde8qwqwUtqz1lnC5yGJSk1Zo/KNH5SdfsMzTGOw+54PSgTuK0AvhvxNy
LIvaFvVjJtq0iDyXz+qo6+J6PWlKyfKZ9IXnuA92mJ3TD1kYXAIFo3+CO6MPoHVLhjV+GnQbqQbT
N8aXu+Ycyz3tRJioGZ+IcylfZV0FBs8jG7lfazcRYpVHeqP+92jKIiPf7IaGvhstaSjmagomkcX2
jQ42zi3/xNWz8SV9a2Dg7OxzDoGva6t4TvE3om1Q7JrdcZNVrXeQ6hcRFM8vsBOFo2BpqvcQGcXe
wJW3uiLbTS+BJA9GbRzHYbqml9m8zEmH3cfOKuvOKs57YY9hijYGYC7Kwron1E0DTZVV3wn596Sr
UcwFKDVeecDNvs+ttswl0wqB8n6at9Om9hptG7RhYff6eMzYPth7g4cvL77oO8EVa50tvlB9jQRY
jOvQo0C4A/yTc+Ck6+MshTJibTIjCDnPKThIGfdN4kkr/NbnRrEiL/9bd1fBQKO7j7+IacMXoAJh
9pgVoudB09j1W19x3igEEM1WhVaBMWeXwiFeCXBRGWuLEk9iSiqq3xMWCYz1dO10BJdeb67Wb/bi
om9XAMxccXHVhR7jJGXyaAFynyRgrVREVjQ1VZrBiZQzfGA8B3G/FrrNPXwdnSXanzPxp26cyxiL
kq7jMrFIH6YlWbZSQEAEITs7J+yPI3VEECW6ERClck0eRTV/1wkcf0HE9O5MwgIyaoOz2qr1EW8I
MVgO/ofZ6oHNR+zt1ZFoA1J+2bKSbOfgSWXzq2xoBsPFnUm2vYzzDrbd14YysnT0a7ffNW1RsWML
oSR54GdsfTi8lI7FmMpuRdn41mXj0SCNbRq0R/rEzIJMtBqS/1hTJodVptO36iTPRjzG9sznwMvP
DF77KzgijfoADan3qmjpBCWGrS9lhLKiCHRtv44zT3DCqiYYMez5hR7ooxJkeRpSQXAc0BN+XoDr
/CSQPqhq1yImopguRMKB7IGMnFtdZH6UIeH51wKe6eYZe38jnC1vYtrzKZIJk4DzikKHqPECUUus
BCVSJf0F84MdT8B7TNB0aaf0QCnrAFtOczYGCAXR+aG2WQGiU4xCgUvDI4yLIcJ7VP7j42TpLYgx
m9cIdZPaoLeNt+cAFCUFqC6q4R/xVDc0DqAOInauihaRrx70obrbvRKaVlMVqyqp1isc+xAOMgNE
iAVsMiAMx1gODaMzp/Er72j8sdmDz1w914QtrKSVtXB3k8BcIbHwfuAQFlL59UvLzhgVLP0e92K9
DsXBeJViLJd3Uv7bNdpVZv6r3/d+23nfa+YnT3rrxBCMMoLWYFvATpQdz+x/UmxnGuq0UEnG7bXV
iHNCHW3J5yupTxJPaz3j4VZmtSQ6hxvbP8wSroOHXklhRPN9z3sXM5yQiOuJarnPk9D5LG4z78iR
xV3XPCXuYhdAvUUO0tXHKIf0E/wny54IPjm1gGWF8Al6yubYJFn8QsYfHf2rcTN/hyoSciupNsbS
nYmiVFOOaEr0/8rLliK0x8oypA4+3dFMK9z5UlDBS1zGD3bg7s1j133Atd44E+gVuSJfCGmdH2mG
QQFFuTmZCrTDYAPKLMgkZ7bdeR6jLJz7DEBrr9X1Kx7ULf93uANGaQugDbVepLPah/QpUYFr124t
UvA8pR1cIhLxuhRKVqM5cyh/yPwPOxmJ11c+rI9fwlDWhiTiVPEdAYDWDnQvq13hW4rQ/EwYo80K
oDr7RvhS5J1xuS4zEQh3xrp6VTvP/G0d637RMSd6kJj/PayQzuvuphzoG5pRjYp4+GRmVsuBRD0P
FcT3EsllwqhprxwjiJ9XuVo3QDfLZonIlNETCTzfAnzTWiYRnI8ZykOTPIaNZnxvIPRjs58fzAWN
A3uWW/2w3DMp+rDWWCcVT6SZ4T1rwJ6/iOPUlmkkl30jSslUlW+ycij2IqSS5KqywoL4g7hJ/uFe
TSzvzuTLGEtKhzXK3drrtHtaHC4kV+aP0WnA4jg7og6kf8F7Lx+NgccEgo/tS9/hUgSvt4ufXgQc
OD1m0cIv9gN/z1dp+HARDdVP0inHuUIthfu7ffpwzKgw4DhH4DvZsXMhMtHim7aZJjfj9KpTswwf
88GguIMDGVzk55B8gid6v2quAj6RJQ3DDVq0FygN1kEHz+d7JEM5r8YPyHlvOGpxJPAUZYioROrC
ZWEZkyE5xXlZLC1lQkwDOXB0BahaVxYxj6t/L1KjECYHS/yKOnGVrB4MlofaqqJF6s+t4sEVDz9f
r8Dh7Y6yq8w9Qe2G6+n647lxVOGGybACxNtPksdr0mRQFiYGpN4wf+9sAQ4U4wyuZo8KUKG2jaYH
FUqqUqAi+nWD14vHoIUBBe2kVn9Y3Nz0GB52GEdhRsHl6FpX7pgM0cwqBGooRwQyhxcMsUrmmJ+O
hEHed9RaQvRUzsSNDlpCtBivGvg9mMTBFjhWz2D7dEj/4EH689dcQRKSUET/E1uCf8PSC2HkMEvS
T5opssEx7EAToiBBiH2vYvuZHZvKHeQKGLJeUzB/u22GjPqiFakhaQfLYu1/eKaFeEzajToS93Pq
1H3/65PRFw3lDUaYk4+cmfQw0h7TerV89GdYzP3lAfSZgL6mPgTVMKbmLbm4bRWCKrkVbLcBRG2+
MJ7PTnnyTK23nDpzMm3Px9ghcVqUJvAHCvuNZiM0CxAqUlagZ0JNcjoR5a/I7iAzYWMkC+cgS2ON
XGDeQsN4JKW7ljbXwfQEd2zyKKGW3npVyG9+HyfBqsmuE6lbJsIZQBa2/pTamX72/UPZ4InHvQHC
WoH75aNspDj9zThToVUohn4oMaQZ3fQ2Bq9W+OEbNDD91rtSOtIkLGtw6SKCPOBPPYHVC6x1eX1T
IZvYNIO/495FsllnSVbhG/84MeoO2yC5/EcGLJrcfN85YVBzOtbB9R019nqk2qvG6Tvz9yX06DLq
EB0x+Tpc4IoanBMhfxtEobDgbLhiP6Wt3Dt7iukkBE3tM/gnBoKbEejWD/MSA/q/Z0A990M5kaof
KhhhFSZ0nYu+zQTiFnyiePiYUXs7R6IisVmvuYW/kyDtDAQlDLC/shNHh+25gVf9Vtg3rOc4P7mg
XO5tibscvcenrZYysE1tgojd8Rmz5jMW/vx0Q3PcoFvihgBsCNa0atTp1j1OgJA+NaliGWJ+WNQZ
KKbXAzz6sD1hVMWGzApjYrjT6hatQ/rbzgyIMjTePueFhSebRha0UnuMPDDWt+0Pu7lyeeQ2FxCd
9C6JRldEzcM4JBXGqtmGvufJjgm4E2KnzdMNlETkmol8PG5WA4QR4WRkiRioRXcjea+0a80W/4VY
M3S6Bb7X/FhkTEeszzSE1TplLGB+K8lj+FMzqn9yew8ytrNMCLVZuCDgGLzzI6Z9u4akp7RNf/ns
dy11CmgHfXEgd6PnU7IZKebRtw83EUtqMUqFINtu72DJfkrmUBIe+oiYkBRoXxIKy/AuPEYGsMAe
/elbXKVFx6nrZI1o4CrcAYo9AiEsTQfd0PDqBs8JihurUUe5zlBIxxtwrdfpAFPj0mz31M4s1FSs
Iz9v36kDk612R4F22BCCX7P51VU8JecuSHMx5mw+eiYH/OZOb8KAAl005ce1q1vkCFsp4lD84kzM
7uKHU6qHfDMYwN1/BqPlfMyMBeI2QWWAjFjbf6WSKR1QtsHnU/j+98WSvD9ypWK7ETi2LYWkB1fT
cVW7iK229+pQlGxZKWrvrJ++KSfkdfjrspzvnj4yKBh2vYhhhkVt7WbHkzcmfrlqeqmYkjj/86T5
h40+cptdipEu5Mjcokc3c8ZkOix1DHt3A2/C3BmKGXZTYqRj8IURaDNFr7sBIGH4LxIWaiW9ZuBW
+WNeRwWioSN0ZkkC7DaVopWUUDJETnTSMzATkRfSHpUkYOd1DmJB/d5dFIJEsnV14o6GYuVAVARU
Ga7F9PqRonQa31AlcoCS5NyYtoU2Wg51c3tvKAiApXbwqdQhVyH882WFUF+1tQuf9pSvtGBGYqRl
awotMjpbVS9dz4K96fuswToPGH4+2TU/KgoYLrQkRwmlHQvsbCR5PpJdjH3aRbXOIX71yXGg/3uN
u0b5ElCyDiTTu2OURarl9qLwQtnVf6zHVhNHJyUGcV2njU5KK5UCHB1bjlkAjNDWhRsbmU4rhUFW
rlCAUe+zUkI4YTOFj1/DW37AvE5FXl4EubaNluEU9q/qu6zR6mGDlBa4lV1mJOCf57vpKDnFL/pH
UCcuZ4tr73QPgTfDBJWKKOmdF/CfxrhPm7r5WvuE1nYjcMN2eV66Weoyv0ycDPJHg4TgutbcYKC/
XVRKQ82kmtIY9L4rYsao/t5vXta5gjoW/uQgCzSduujDJtECRm4dy4hoVPCiqhdV5y6hbDW9esSn
N6/BG6o2fR3tHiDGKJxrCIVa/YGqrXoO7szO42lz1lEa823VpAfQgh9o8ElIPFPJkRl2ZdhdJn+w
ZCYSFzMu7ODyFX0lBnKcZcmrrOB0lraM9sjd/QuQCPDzsglCvbveViJAGJE9jDynvb5PSQx/t47n
7bbuiP7eOwF9rqeYBNhvHo0g9zLfwDn9MOSsgwmWyTuwxx/bOCycGle2rfp7+iR8RJxe7e6GlftX
k/IP/WTGip6w8zjsh14P3kbylgugJHuHTDu1A072g///Edlv6ZQiF/zrd7eoZgat//VElU9W4zNC
YL83zhXu98BV+bTlgXCVIziBZxXaupfXsioCfW3dQjra1jFp/PPz6ieX+YaRBqoyyIdeUeMxz6zL
AUZoNkVen0TP45tYy+T1pFbhivURnyrSImWU7xT7KKj7FhooBTJMweOWN0aHtb0i2JBGD5A5F8vG
4CUidehExE6TJaVQ/6YGJX86psbn6ObpNn7X6nNV2WHeAUWP9fIY5DCK0E+xtsNWVAFYixn06vWp
OT3o8vZEhAj1XcfooxLtsA8ArmsBga4YdfSxnRgiEeDXq3wCBweMGk/V1c0mR/iwIjJyewf/XxmC
ocU2eHtpeOw+5qRXayK1H8OkfUzaXXABl+La/gAABAEiCU1/OhOPWmuheQPq7GPvIClsxx+jrh7C
rWxaNwEun8ZP9guaazhiFSxsAfd9WzT/iINO//hvKblsFYVbi27YquqEWC8ttfeNDU6Yq5mjy+T7
wBrJ3eD3Tv2X9wJTgsI0+aAraACaPHF7CkTQwOCk6J4fp6qmwWs0DUJtkvf7vlbE8xUhIo49giXQ
Bzp8re45XOXDFlmTNeniOYR6za5SFCjZIAFmJwr6mMu66EdwTnf3gdrrwx8zcimbSlUvduJtu0KE
vFP21Avl0mPn5mG6iWcvaoRgOE2FEzZxTKYHwm80zYHAfzIdJRMzCyKW1lZ5jrpESH1kj8Y37C6j
dEP+xNb+wPlWEOYZQ5MllYhu6UuBW9KqXjh/rztSh2PbbgmQgVYA6lh68nlGSD2TZtU0Pugwc1/R
M/r9s6LMvTNML/Kpa6axgnntaHlRoIb/GihgmTAoAoxHx7puh2G5oRLEKeoTo6uWrwkBkob5Wy/I
JsBdmBB6MeBsmvBp60NrEpuV+FdBioC/HeXgsJ4DTCt4J0Dc7RKEntlfPzUI8lKmDk1jQWRHMWSB
99wwaJI+GYY4Dw/ibniff1x2bCg2CS8PUjYSt/0/MzxUrJhgMuFpG/ykjPl1SHTnQGOnLZy2C0We
+27LFOUb0p4WCvorHQrA3HApIXWSL8DLkJIiuCD/S8pCqBJThjSVMSgJqqpuexHLU4CeZ1hxgnCE
NI4Vh1nCvESzkdmBwt/0i7xhiTLIOpq2huOXKaOiPSHtjE0eKd0EexxwUyqQxWfX1/XU/o+5lATt
O+nlBCDCZY30YCapVK8ThU2V3sRd4P05/zn5sX/b7Tkv9LL2NSR8dWcH8mOMqnAkedYSMVwBLNXm
+Pmsm1ZPgikMn1Y7OwaFrBHzFVm7DTbwdCE5uyeAlXqQEnSbk/C2Id5LNnMV+deOp5BalhwQ9EDH
yQvTCNn9Lwcrp2zOd8uv1eadWFOoqYokojN96qmHDwBexLmALkUgUShQ08ZyZGBQsRweBrGNhVhp
AhKOwjMxuNWxjL399Uv4f45P7C0jQgHmqRauFOKg/McIdMJo3DI1QaH28Q7oP8G1pa2g7zofgY5l
YPzewG6Yo5YjHvt7G4BD8kJEZqK7QRuQd7GTzcZ2TC21FFUA4dERI5WqySNewB9fIIZ81IfBtV6w
8i5Ph1XgEUHa2IdF/r0SrMzO2/6kQzkNF4tFwprhj1tFIwuNOB3zHQrg4e3cCerqx6kXDXphqCHs
zNuj4RLHnMy9Daw+bFfPpGVXO75Ut5lnu6da8ecME7BIF8RTt/lOXHpacOQkAximtbkY32FEBdie
b4bbZ/WqmPil9hwbu7KeSzL3vGqbXJpc1UkSV4c3MS7oFVMRJ+KL4EDlPflxgk4zFlnCGc3GREKU
bJU6FPLYR134j5uKk5y1iY9c3MK2bep9QY6dDaakzaZ2C1pa6r+xZr6IyMxIUSO9tFRfy8cgyyJX
Uf2gbs0x58O1BONEaouT7xnTbO3fPfRlj+blGRjy4vEyFHvTIB6RLvEhX3ypWLPA4MEIk5rsK3/I
ty27bkobqNIjLg+6ERl5P3MGCli5ItxNKEkghMvOcfPuKgZlj+PIxUbLyp3W39fdcwusTb7l+nlP
PNVYfZxtTl9jX/qVlP7Tteuxg9bou25e92bMu/AdtW6XgxgueG1rJhTulrvUCsq6ttY6FbUAxt28
MTsa5NSU+CB4R+Wqxual4ONi7PYS2YfTetN8hFJowicqTFs3tZdrtbP9QTudqfkFRMdJFDgtTzKc
8WGzFd+BY/K4XzPhO1Q29g7aNf2MupDdCI/N4qci8vG3C4OTPaXXmWKqkq8n/ningaHD1P0Rr3Er
NWXldKqpk5ZF3YpoeD3m5xhFAn34jvJ101hH/v502DQ/QV0wzLzLMwKxoxmUeAKteyr79Aa1hxlS
DErOoFbDiQE7S6QHRWpiUErz3a7xyZwQ8nLtucO9V7+1FbFTLvz9Xakf2aMaXvamCoT2/ARBZvPT
IH5ZLBx8QFhmaBGAh6KtDLaLFEjOvHepiBeWn34yFnSN5IFmFeR4yTAcg5dyUZIa1tBTTGGCIksX
lm2FbmtBlajJA1lYPK5o294Y9588rde7rwaGKzG60wkDryWoTZcI8r9vwkp8cba/S+m/mbxYh2h8
oHgyhOH6j7r8lvvvwKMfg0vkPAED4jJkBRvXResSfsCc8ne9P1ycbB16QXeW4jrCRzBLv3hWSRjD
2w3xcWrUhnTV5ISUHGxpvEXBTmtCy7pbCcyl8y+Lz60iLZmGuNWKtakvWToe+p78eIOUejFAq1e1
33IaplXwCSRL9N/WCybMmm03NjbBYyFCGONQzcHu0sAHg0a5lF2ukOINeDQ9Laiw4vdOkpgjeWtZ
7dkFomht5SB5e4edM+MW4ZUAX8XiZCKgLcq/83/Ds0rIzIr8iru1dWrjbZEVGdNOO5C/pLR59srh
e/eTpvAkiLM8B6gLg/etOqEFP2xVd5TersRQfgjA5wbFnAX423I7TVBG2dBJs5i2f8KEa0uo+otS
p8ZIqvfZjZX3pRD06clM8pTALhucyvCj8lVdYpQAu5j2YhT4+Ml0NnfSMiM3UQZDHW5uyl5X8uCk
aRSL+7lR1Z4Ee8K6q1AaGsHVDBQJXPG37KlA8N8W1DAEGyM3k4z2dlvsEZ4RQ1tFrnjsjgzvfT2l
M15ZCl2C89dDGtfvMZ2jOQFgpbUKlUHEhdTIzQnC2fQ4aa4gUd5qtvIo35hVCFwa0XStk21jhy4F
bQFNgLjrGG1GYmB9csjHfWrM0HVQLEUnzh5b2J0wGC01JflBwLzb3hq/QtT9SV3K5A6fG0hs0ukp
Yf5cIaBSLsjaJ9m3Rp2DmVxYxVqh4//ltwsOSSXu5VwKEHxzCUNTnFQL+SUn+V4MG6Ebu+nXu+F3
fnUWBC0ZTopymYmKvnl5fInuurdkVwBCgnobMKxzbhZEVd6cTetqfpt95Fs0nPDa0l24AOsx7bvp
jzpiav0+pF5oHWNrB/f8qDNthIOqahHBItk67nysOCXDteUB7TB186o54EeMnL58F1yhTz02Cyry
MI+TtaFvgjt3VmOqjZRFxFzRWFHkIv4De+Y3AqtJSdL+lmMOFuRx6BZiJJSWyfrz3TCUp68Xob5W
uf+MsZJfcnKpJu0amRFfSM3SMMwhnQVpxU0UFylCvxEaYgJ1+9aQO2Tgop5LQvrEGP6YPNs6I2GM
v3q7FNCK9L0thUZzX9A2uXXdArXaO4yrHVX+BlNio2hmCcH4+r0HgcD8bjFY3WYIuwt8cQr5o3aN
BLeF12jNhyx0QK2XIBjpPsSG4Vp91ljHOEqcHRFfIQD/w2OxH+TaAa4fksNnKfttovbTbPGZP0lf
omCAGSs3+4O+MI2GRzmEZnL7o9KoL13HBMCAkCOwJz/Ym/JUctKJcxBO+mGGiuPwIM1IOVeuxL7e
nAwxtsLAWQl20KB7i7ctUucuUY3C6r1/ELO1fOT1bbdk+bQyOHAkVairTAC1L43n2DN1UPSMH8aO
ANpzQWSgO2Wm6Jahnxi1PsjShhfO17TyM4xZFQ/v5AFyMm7Q43Z5OHom7hdp7jFICXDWt9Z2DOdw
Aa90nlAQr0ZokIORF4MuZPg3NeJP2kRjkOEIt6efnGdPZLFnotCwOv7Df38WMx4T8Y/eCE5vFEdj
iz0qRyOS4o5EdV21RJJcGHJuEX3ewErW5lVeIFlNZ7eYMn8dP4EBXkxAAO3dkU4Qe67wjkKyfeEg
cptPVrolt0oqVt1lokSbwyu98YHo2kH/xYEglNo/NG0TU//9k3+16UjRmDWNG7vD7DwhR5m2Nvur
Rl2JDOG1YZ5t3lRoeucUVUoOZCbKSPNz7u1kHOkwepnbyvM7b+XlyZgPDalbpl5LR1u0PyTAKUv0
yZxSwD8GPIiYdD2pfHdoa9G2PcRczQdmLJHzX9+xWPwTty62XwpO/LbEX6pGufl9YQ6P2eRZDpty
ZanFo9Y3scMqKqbTbh38ItO1+/fU0IHcp+Mpbn7z7SSVQ79+mMyC3Piugos1ahVC3qJqY+Lgc6ys
9Y7hxy/8F0h6RwGrQk+vq07PJGphNm1MAcceOqMKNF0KXW5jan7i1ZM+Ia8TzlLF9+FEfBKoD5yn
fs2uP7PM60xfGZPeTUQU/NNlUq1RUowRPEWOcER6VEfqq6loRQKjWkCxTLYFWCcdLgIRcChOzapg
BQuKNA2MwcsSyYXTP++dMPvtyc5Dp9fKTRdLg45R+zO+5gLWi28uDSy7zOh8+N+TdAgQhqEFfFMJ
jLNeXPSoTTEhhcruPpx0TMkHRMhagNG5ybf817MvrBJhVSxqWBWGTv7e3GBTa4OuTl7Vi95jTDjW
Ard5AgOzdLEghAIbdIoVIq8gcwan5kYmf2bBpBPzNRQtfT4dnGQi5UrZmhuTXXbOJYVb8kS5Jd0P
zcM8wAAKGB+B3c+uXnT9Tr0oqaFrg46qKFEBEC6OblTgLdCap580pAD1K6JOgZh1x69fpYTeBFwn
w/u418OIO1LqlZuTkOQ2VgYxpw1czTpxjCi+zKBMLD4ctyJcf6a0SmQ+D10MLvjCKrjOGJRfI1q2
svm70kE74vYguDMXDm7iAmc4ChizMtMzlxGcETHKWLkoiBhdiNUIGnIJbHDhe2DlOU8ZiYQv1izW
hY8R+FotOVv5sdU3CDeDRwIocWLNvSUS2L7rMRbwBVGWRPaTbHVck1pAxSyM3m1cEEDftsOxwUda
aHo7ErubH8fg8U2W8+Lamlv18vZzxkFIDiUyc65akdsKGwzvXdH3zEqmPr5HQj4hfE9eeBsY1g/e
lzBXlLNSkTLdnqJJJPGR5gC4IMkqVEnANgQE8zh7U0eoNSnfrvyM9Bx5b2zmxgD28JuHBLaPfwqY
e1DcvJvWIUr9Mlo49B9TAmEhrvyAssyJCOY1CvvDAGiVFD95EJbJip7K8L4cfH0iOYyR8Y0WChnM
HZPEZCTk0Bqg/bcwxoP+rB6QEEhrbmCwuGCzWMa9TYT+MdsHnfRKXg1SCDk030pzb4B0Ip77+d2L
pR7/aSPOREWBppqApWcCpOK8FYhX/yB1FAP+4hhDApiFPmBw94792gZ8l6MGyHRmccfNGpjRtyIh
RiIaTjPh3cztHgau0bOqziijrNT/828HnBZqCWHMjStsDki0XWzn4vs7Ig0AuTXmwE7lJb211Km7
vAHElpjAZVI1Xr3BUSVfK2wObt91iDtmw6Pzq2g9ozPxtsrWmVRyM+bJK+cv+TUIomOCwLE/6i1J
QlDPUENLp9zOejCXDLgidwLmrBxoXQxOMFvHx4dbkizsq+JTCGqAq2bXVK9uc18rV2ScSLob96gv
lipQ4tpxOB9c8gdyLGcO0spEvvvqxfNt/pALy5QSTcFt7JPKrd8OavwiKZq2mCBbPDIz2V614UqR
2Ojg49RUudHhg3pEVm27T71Wb1LQe9EB4KEo4pOfINzxaBUrrpxtiHOx8MdSVhGw30QjvkBKO8T9
lTVEyQiIUOrkhikoi1NWYqY4jp42WljOxx+eMnDep2PZDMiauSUO0gXNBWe7TZ3HSP/J8naHDCw7
xmfHM2BPPjahGWyjbOiwyLYwYE/9kSIkMLUhpbWxeDHa6/bq8Nh8ppR0l6+GX5r+eZE/ob8Xaejj
uoFfCOag+98gZbgk8hb+LB7fy9NCRZ1j7kPOY9QBnhQ0MA6eimOPpHmV4vV+P8aJf+jEwY4gborw
ez3o/dXxtH+7BgyQuccSHWfqtvcqbYQMvO/mCXftaDIsIBw3S0wk9aSz0iQ2wkqMQtqBV77ZhHVf
Y3Oq3id1goQYvBnFJc/9tTs+rsq0GudphqasqIx6p8x25rwy31kdizF3ZPgJD+JTZujLQLxlQjhi
TRqEPW0pPYokmZbN4zBV7Wjepjkmmt/ApkV354EF27rPWodgKes9AKQJTo4Pe5w4s4aSdNBbFIUj
0pBQeUIL6wPyuvTvtUgdZycbklEe1zH+eHVZUyvMwBZU+snx0V49J6/yPWIFITM0KqIfkCBwAziM
Xq3gkS9zLDzoOMqeWy0XnlaHkuqhrepnUOsix9e3wzuC0dLsnytXkjEJEJ2bAiWfYer5q6hmWwfZ
umeeyQxBKZgI/fubBkh2V3yRvSEJTUSP6Wh2m6Fjpxoq1nalwb26zBHivwSjopmxSHWzbPSUzeO3
228kDGdDm/V+Kqnzi0bJDQFUMjGE6tXm9ZpIZp1gez4ElAAiz1G+aDLNRaOYmKFmTnuuPUmP3Ls2
qVBJWpC41y5tsRsbD1EjplwXjXcFJrIlrfXE9cI5ryNZLvLp/hWXYanblXzDF1csR1Et0SRyNYbX
L9U9wTkEdEZpgMNNQG0IayaoZ9mH/uNke+UqKRN/1JyfoxCz4XlxygvIebfZLE2iM1k0TontBFQI
bSYQNl+BhPGsV1JpydRBVMdPFjGjLYtJnlNJLgB1JEu/JVCoIDrQnntKg0QKON+odhptPK46nNjZ
KiXm7sPtKCFsYnIsUyGLzJVJifaFqAeWjZN/AI+Aa9BTIzrIlqbu6ALmh9yFVWB6EJ/j0Dh/N9on
RZDAj7Vzya3LG2EbiPvB7FveY6jQc+yiI1pgxzMuNivt2+vXk4vRgTKQr6JBaFSoAmZgjktCF07m
mu9qxn/B51ANJZm2i7VFMvc1hVH9srAEk3I5YRquEDi5UU/Nle70mHAOvyEI27XHeTN3OuetZsXy
9WUIGoX9HfCt2WuLuUOPO2x44Rayuju1h9lAtd6kNl2kN0kflogCPeCLYEKqCKMlq+6Zje8uwQYo
sKxoJxoiKsxOzcvAAf9Ssza/1PI9XxqM8WaJRq0J1IDPSL+H3HqE6tonm424xuVERAEhBdMSzABO
wI6MYTfh9/6RiPSdpB0Q30J/HbdwEjiOPxAlSHReUtjJ+wxfLMkwaLCoi/MlLv319VE196+K9g79
iRuVOzJgkUR1eDqd/7Fvx/2WALJK4qGTek2JJgEgC/0yKqccgioU+5eZNRgc2NaNf9zHtOvZarxr
hx9x5e5p4/k8c5VQUcvfDDy1vQ0vSgjnH3RRQ3xERsW8IDfZVBChmmCoalMqIsP/xTSjj4OCsX+y
4WVtkuya0iw2YQNil+ZgEeBD4EITZ2UPBYNVzXjeK3xuk5z5yqvJV2MNkEQQWTHOemym43ge/0QO
/kmcq4dAAPeOXtQ2+leJi+yX/uybZl9CJXumnBuw/EEGVZ7xdJG/23e9mBsvt0PBS/f4huosKvmS
23aFmk8qgt852ZMOGVtFfceLlAguIbZqZDJvcIzw7oFcUO49UpVpmIicjt50EK15/gd0tep02hip
N2uR1/uVWJ9ONzDo2f1qd4MadzuWl0aDCoa/C2AwbkOWnWtFvw0MXljMc7Fm3tglgqFlLEfMvhbi
gH5FWfWS35P6gx2iRLGqbq6fWE/4z4n2mCc9MDbNgUKgroVuymf+2Koou0Zl/aEq8DvQ8HBqH7t7
7dtI2CImS0fWZE4BR2L0z4g4ttUEpW2/OlRqd+Y8EaQ4NBuVWqhi8GnsYUd7UTJ5C2red4vZZ+vY
hBd1qgHdgM4ab5C5oWabzP8NVJAgIeZw/XTGawKVo0h8bp6u2RBlAX8HJ7qFo5VcsthsGUzEWzGa
SesTwqtnwC2lQkJyGsOwh9wj69u8j8BLPDb+LNh7OX2lOMaxmDbuplR5hF7zo/o9NywzdO0A7R4Q
euD4KsHioujeGIagx9tulXv2zwdd9nD6F8wLbJkoel5h43wC3uONm1HTQ/lER5bAcvwt3zLUVrId
K/1XJkI6wjEqNJgUz684LhfhUSSOq3CjXHL8WY9wn1HBDP6EZ10G/r9+oMEgy/8L/Wr2DWT+sSGu
6dcbxXZQp0Z0mPEmCDwg6ORGcWhUb+KZurYeox4W4x8ZtOI8Khra71gL2W3gHGszqLfI/JZPWX+9
vDZ0FiGepdIoAH1gTJY9jHLvRYXX/JGXmy62O6gd5tRl+JeNwTl4q4GIxLMMluYCOdjZWgn07Qhm
D3R7ljkvuCBxPEOhmsyYgSygj0tSOMh0l5RE7zRERM59tODI3R+x0pub+XygLTNs0p6FE7tRITWe
R6sGdHqf8jwGGoEJh/HncsVYrpW2fPKteLKUKQnm+3ND8CxGrHUOfiJsasQyXUeCVkqh/x72oRtk
9gD6s5Q26Ir2R2nbQjuVmCYK+HU8b0dNdk94LlcyyNkH6V2aOp07zErgHLk2B14e8Nv3KpA+e4T5
iWiWw13IY6MQj8uotVxn3NCoHL86lULNNV/75ZEPvbr7g4oExbXWAr41+HTtzf57KffshbOFzpO2
j0tk7NLFMGipgjdCia3AGs6HGPNrjXvKrf9sYjr1RjRuP6vIbN6eT2EL95F03r8UUcpsi/1l/ZyP
yjEaVyTslOIZbkFSbO4XREK6MWkje8fmkaye/qwkiHc1igHHvK5Nz5GMUBZeG+IcJaO2aoJVWF79
x9lOHr/1JWKNKK9DupfHv9wmw4niY74TXOKTLh9dcF51SmkuMgsheQp7EbIChzAbk7VtphJ/K2Lz
14hjl1Ab/fAodJCbdbsSiikNijzxAV478kTgdQMLjl8sp1AFIY36OTN9CtMVGtNyprzE1l0f7DQ8
Vts8Nhw+FzWFynyot7CG/4euuYd3TN7ooO65sGzGCy9U1doj4fyDGkQVMzdJOchfyyC+C7qftp4/
BoGFUSxs+BH74KVlHwRGvRg+dRPfv8QTjcXgpj72H6eMVaanDCDCPZX3wZQTugHvvmLQn14YHjbl
CVspOlMgtOvGV8HwNc4Kb8thoPZslazKDVP/rSs90NQD8keRT/zvhrR+4YLvAHFkdQKcDJXHluul
O9PHepXDM5CEt1w2fjA2ZKlvYDXWbAUsm63LqUcPGmJw6ENV6wyymjPal8ujfNuCFuYg6n2dVYQy
yklawDZwqDaA04JvDchrghzhPWtmrFOYMxCRIbGTK0NjCrcBAE/XaUiPhlc+dx16RXza/HXjtocD
EW4RBy2L+fJSk5dG1xL4XjS2Fnz+ml4M9fhRbYmUuC6cnSnbx8We+/GMFlm1vNVPVgprezsdIbEt
p6vko22Q1RYHmU5sW5mjgWjo9sFOu0aNKqoypiq1dOi2BY4fqFCY6G99+AU/FExMAcxmtBvjYYUH
vJmEJy6RhSL5+hN1Y7Sf0clzSmSSG1VIfMCk78hiZqqzGGpBuCCRp2EoG3oRfdnCacga7WrjkyMe
EUDt+CoL6Yvbpa0KIWeDyY4dYHVJdhXiKtkYyNhZJOt1rNEWkqsuD7rvQNavsIlhQidlHC0s7d9y
RUvLhOY/TxjhNXNankkxBk3SWSHp1NRg7AQmH28YKGGy1VD414gRqrS0CFAZXr2ji7aBz4Z1yDsB
Ola8NXXuPB3pFKiUgE6V+XSMu8eJ5SqDiENP+MacfP1IHAOfqImZHGorSgkKeSaNX05WZWxaLg07
P5gU1Pv8PTDqltYbZMNlpS4QYIOb81XlWqy4tKoSWhgGuG73ZjdKluLZTa2xFretjENytz45AHQ7
7z9C6zceRJEmOdF1hE6t5bXPK45He0yQE3kwiZEfuSbsS/qiyEkWuQRmtKw7QuTVqp2EUNmSfO2d
UcQFJJcWMQpcSuEWxqyLCaqpSaVDmYDsLBjjZSn7sAbD02z8Va1zTgrbnM8+dS6QGzUJYQzcvBHO
azDRHW+7Dgcj4c5es6pwEEt1FiAfDAk1SwsxpIrF0uFHDrPmw3dsV86KamM3+bQfliw+pUw/Ml8Q
mxvJpIlonn7rRluVResbAvaLYSvsRNPfK3LY9mth4x7nxwuLWEdiuDnLudbPN2h/xFKqqVLCdZ2N
SLRzVh3fknR9OjdBAb2sSVu8poDjZ7kLMYZIQGMzjCIG9YlWfv6IuIfZcoYP0py49oIkpeF/yqQ3
O6V83GOpZVHIsrzU5bQMq4Z77z0XzCaa2xf6WmSRsPhG+3lAbAvrWs8pfpFZfoKXMy9g/kHj0OGB
hPzdqgRcp9+UW40CB+RHTI2B8F3MQTvH4Nh0yIeqEngE94zI5YIAUwuPg0speSG3w7r9T96QsWrU
0lIodvpI8X9yu6ucNCVncTizIDfVw7V6cabHYxOWtnJH7O6T9/kNL3Mij9K0cCY7kW58uKl1yQMv
5XvsHlc+2YkZEwA787hLhcDnYsYHKYWkaTz81btBczBqV1DqyzlP1YbmKYCtTtXtqNOQQo89Cao+
mWWag3QanDjN55qJh4lELTqCJLyLhfPtWl8XxcKDqG1chUkWGmntqfWO9ar+YHhKrBf5+IplnrP9
APvuf9udWUkiUvAg6HzhW++l56wuGznfzon1xSURPRv8GWJQykqdlpCsRRYGauuzqBNXTyaP7kNk
r/ZXkwD2DdMlo/8w9S4x/0ID1k8I8o7TwpPDSouB3vNGL3TjR1oCvMdjMj3ZNdhzH2mRdsHTiG+x
98UxqkN8DyyMkDRPUEL/5sE5+1grOR1fegWBwFXVR8SGCzmbFuFyZqhSytge7sy2u3yqxSQhu56X
qzFqJm4YtbM9kJ5FneT5EY3vQm/f2KAHk0KbADoXIzJgWn5YObgJdHXuyuFfhno0oaq9sF+vA5ow
w6b8iWkprZ0m+hMGk+ZQ7li5x62ucazFH0WttdAd7lvexTyZLQqGMy3q8czMBC5CyFQ1t/q3XQTl
ifMh0qm8KqngGUeFrg7ck/HFmItb6GSP9XgHLeB/JnC69O0WFPG3v39S1vRp/kbfbR/MIHQQTcfT
bSccxNEqodEvQmxg4yFukvdCZ7DALW8+/leeHEDOmvN0j312pFbFhDFTXEd4neVsVR7BO4F1NOuQ
zypgDlFCtfuyz5s1bMeUERk5VdrOlic9HJrGLtS+eazvNhgAsb3csvtW67Sroa8AWzwXGzEe+a3N
icxxNR2icEXOPJk4Zhq/c2g2cgu/0uBdACw2q3fBOMi9ZdygCSc6rgRCHqCpYtiGwOjVJK7yAB5L
cgdV2GeSrvneAEZ7AG5f92+Xi7LzY2CI1ITiiw7pfeuhwiz9m2avbZnj7CJbqkWQah19J05VM25c
4OhZvLvTUAdLBkrJVQnQS99aExk32UbmGchcRECOi5KsyYEtjaaDDqTdTN7/LkAz+sYCtBUocIWw
Ggkfs3t4xIUjw3mpDlFSKM2nrdgkEseF16OGYB1LbrCzU6LgvBqX/2Faulpn4qMhfwbXBZxervqs
PleW0Yiqjjq9GUqbE6gN+oA6ppizsnrObYoaLqXK4qj9OkYnV1zeTn8yoYis+Q+d2/bHTasTDUjc
a4CfVLJvTra0gF1usUFoYKq3wr3azWPQcGk3rr+2P9unUp7HATkqDvW9hyCsNMDTe2r7dG75tgIM
77Ze0ORojhKt1XFhiLfjQSFDLaBs+h4wCJ6rWE3fdXDyubM8GMXmohrxG3E+rVlW+c8v3N5lDSEN
fBdu2wf6h2XcuZJZmBSNb058DOCDFID2Ds2V17qB79gXXCKHKWMnCZDJ8jpE7L0uBUb/xNjsm/uT
XUA0NwxJccnDwNWKqfjd4kUvdPdD3c5JKW5CF38jsPr1t4AbP/pZDCOYfxHwT4pronGmpusrLtwe
8TJDSFJGipkSjIb9GSZ+qBleoBYooV0ZalcHGtJYLTyk4Q54YxI9TBMsbeRhKvnYdsv06o3p5spo
7YkfTIazbQBBleth728m8BLspbNgA8Q9hMaUIyZzusPT/GdMPD1JNIU3jpj4ashOV0EhLqZEZqvt
wnkh2cYDkNIaLzyuTCUJhM7SnGXzOqMa2/OUlfEANHSYb6slDNFKC1QqZDqlPf5eYhCEtGw1Ul22
3JqklusEbJnkSPbCIMKpzFbIBeCRRry8gL893PJ+u0vXwxkLOSrTIUIiQYdbReZA/yepHjksgSDE
G/3uNbxkqYhIV/HZ+gIkx90qqdDtcvFKqI5EJCz+WUW0sbnCAb9SJ2S5SJVY036bERz+AG1YZ3f+
+QIMPHxuYThdQf4PDqUW+S/KxTQKeexRADmRMoSYs4Ooe3HO6brpjLUYAPjkiotxR4TrXYcAOb7D
ZexJOMr8c+ZMqdLzvQzaGGScJXjr13BtTL5VVFDyILQXkVas0Uj5UHgBS2Wweun9iN8vNGboM17b
/3vcnYjoLKu2Q2uPGxsxCEVtQ7tOq0gLN2C132y7GhlvBt9lIc98/04Sfnz7JsUbA5w90J8k+Czy
7sQKBQJCBymJNZWJuPUEWi6X1grAkj9M9gP1QKpiHTxowAoWhqaTyNS8Ec13x4J4xGZ58kU47kZV
HiCxbJXYJWOlRa/TYt2Ckxsu3K/tj4RtynAWijOLe5pC5V5xB4Htm6epDu5uhr4LhgBWJLEjearx
iADWApDFAeYk15aCvY/rzEwiv9Gpr2f3UyYs6Xd895JBccvZquREck7mexcqK2rLxHdIq8cmVhDj
DLHkVeduiY/27EuZOPrxkLnh5AQhoILoWcY4JoI/U1XpMbLO7lMbo+5Srj3vT7UlViKxvzB89Wbd
ju12JHpuVi3/3W3ll5OstfrdjPiVRrRSKcCvNlgWnP6pJheFxQ2e14QcRvNy+TK355+UWTqfF37F
2CBNTPw192Kij1nqVO/CD3t+eYB45zuvmXJgbKo/QvEprY6/H8iuKIDujkgT+IENCyL+KBDgzIs5
DQGznepI49MNgdQhz3l2M65SMIHsQoQqFe0N2cWfc52CmhZXeVJLQcS4BGCRteNt8Vlu91aW9Os4
pIpRoNpD08XLcqhQMOQg0qF3H2OY3RFgzPLDWMyowqTCwRfYS62EGpII3Tk3HvJA+n6+dQqkRaxe
67ExE5mt6UJzb7nf9dPkjqZ8rvWDomViE92b0wzdsgRNgLrefw09NCblstMM5o7cVHd774qjjZiW
YYaoPfOrOL2syhMvyAoQPU343zHx7oKTGY0UA2jDxVrGUoGxY66s5YR4qnliF8S9+OgwyEBaJsNi
UHorS6pSNKoxRyLpgGq7QGhTONYyrG6b/FL5rnRo6WLlxsvz1vLU766CNy513C/nO8UOh7mixHBK
VgJ18qdLnJ3LnvPK/DQk8/55ohi22CvPCd6st+ElteOBexTr+fZ1lpaMnew1DtP94lm9RRWF9jCE
7L9XAhKbpn60363AV7UVQvoiG9iXrFr62CMznZ0IPqBqUXixwebJs5v1dBHepXnqVG2BfMAN+C7J
riv+/fvgIBpH1E7Akpr51cw1ibSAfQGylAyRCQb6d/JYsGCq/6J8/lx6ld2PdEN1Y1a4nl7vmENZ
He2//Mrrkxzj3Aiv78CUB2GPJpuUlw50mC1JMf9PhZTBg73H+Lt9d8RL6iRGBz3crnY8S1a4QX8M
rUdQXMAgtbeTHfdqwSP+N4MS6JU2GPeebrHBGGoAA+zFCPQ4YczPB71SxnkmnEKzXtlLNvlsZXCn
ULRh2dEzBG9gVxIldyb4X+tuOXBnlxgdigbfeMXKaRjF642j9L3+a3SDZ6YTd4bFiYl2uzh1LAAf
gIOXc6XQ3Byu4VYaILRO9+F/I9GtxZSyGuIem84A4ztuelonf3l4ZYYoHQ0mBe9CsmgadzDjDvTu
w6fjA2KjV58sdyGxa9LDM/lQuTbpXNYwptn/AjN3Tfb1w7THbrm5PwIVPo8VS8aKEXCTj9zMuQFr
7/+PKichpgDEwLfp5CF4JtDIj1+Nh1Mitq9qimIqrGycdfpIDtR4/k6CwZnrBWvtuFOV/KaMGvnK
QkF3XLwfL7KOhQALql375g1/y54O8SeEdQQmtvBVjCprBkGWTkkiu+MWmnG4g40B5DwW5ljXSvyN
s8Qwe6CPAvWFIlC8I8ZYsWoEOPFIj4bMx91xLAzRc1hCSHAokFgjaCO8EuOFEmzhHWXZZDkEsd4/
J3XmeiBJF1ZIA5ImPszwEMn/uFvuKtvNjSZE3kIrydwnbW/Q0tznaJi7fvT5rtv1fPF3UglBhpv/
LdRl+R3nE4ukGu4lPOS8LGyFXgLJkatB51Ot4gzFUVdxZaqcL8DhDkl5gvIkuLcI+DWFLU0CV948
udmRGm3+JylPdYBqH1PDs8fHeYX3MO05BG/eJuXIibyuTM/cGblYRY6e8hD3dqUxIdgpxHglaLx2
N9XMvFI1XiiuxbxkDHqknXko1OqHBUldPndvOEUYOdR0cuWK0LkW5mbS4UPcHA6xNiExWxSK/9+I
nXk08GZtDdsTUOqxcFgUFcm4IVxy8MxJdxuZ0wEWt1MAfkPC2cM9aeCKgBJ31ynJqUHDuzUXRS8U
dUIEn8N1QZU8YY9yioMDEkMtYYM+GzpVCzje4gPym85muW5cD+3tjgHqnYckZ0MUc/TSPfIZwhA/
XPoW6VaqaXHlJ8pcGQdeW3xRQY2EazGf6Bzj+/CFhXmxkgh1pLmsj0o6rbc5dZIddHiT79eY6/RK
FWaHPZWsaxfsnfp7Yg7+LqtoTkIoZutYWSO3v6dNRI/rQd9t6a718OR3L/7yMiFIJ3FLNR4sdSqU
E/zn/eDBJ2A1g4LoRTQgwq8qP18Rea3wlS6ajftxUaeor3Y7uRNSu6SaPYlwnLnjrATgCntJRjie
OLyn/OsCV/suFcKU8g5D9du8vsiwrIlkvr7rGJnOmOrpq003+xacl6x4weZqCrc251rvA5u1aAJc
EAy2jjAv1ZcM2TGMw0WH6VWOYSlgqUriHcryAajhNwnpZD0YVIlsh0AtpUFc9Cb5ynMVMkCo0n4o
Z044jGRqC0LvfQ0Rz0oC0/yEP2ekIJ52Kr1TA5r76AWMPF8mvy4iQJyXOwWq6LUdk+Yl0CLGkpMx
iwtcLjoe0oAHtSmQAYCoCZNOEzEIbPOsbkKxFlQH29lySfeZDjtVodmaHdQyzBqieuukZekTbB1g
fFfo4wcqGExfjFT7XdhUZ78lb9LV5ub46nJKgLpAwnvC9UHzZHzwu/3f3LgWAxXiieaY/updEfMX
jtqDun8fazymq5Kc4998gG3ja2YwfZEGhkqKrUtTu1MPOQiLNMHfwK069iFC7OpSxLP0IUvNpQAL
0abz4NNcbVZiAd887WDUnuCRjsEonNzJg1LW78p+wy/eof6rJJDb4qE/EuzzvQ6k2dfV/xgY/+EW
skNINbAs6ILQkXfI1RBpHUvpsnpCFL06OpbxhGVY3yNLqfmGfvU+a4c6Dehn9vwSCYsenahTj7Lq
oDtTArrp90R+0pNelosGTMSYZQInDP6oj88Nvgd181goVam53kQJcItoildKNpmheMwB67RPHVug
P3n1ZjwfpcfFu5KBqYuuXz489tZ1uzlw+jFrKKK9PVT898zK+nJ7A21ezxVuswEhy6uF8NVf37oh
9lO+PJYj18eH6EdIZKv5l6+R5Xkt5ncPLPMabKN7RAnpEwwKlsovd4JBcYFKWeXJhRSm6RoDbtq0
mgiwSKk8agnshqPi2XWFV/mXLfRnghZ2luMaA/NdFO3usvHyQor9C+dwm6kw/EumWXX21Jbchvdk
IeJqlfKNgVDsZiDLSmvJwWqarKAaYMyNjC1t0fBlxYs7OlGFX0eSxwJgXI3BFiu44fLSyeZkjVK5
KOIY7xVtjxllv2QkyNSXy/kShk4q2LCGxKF5fVKZFBOFeg/bukN/t+JA1G2gLDPtPsNj5FyP2m+b
EjJu/s+QW7VSjd7SnQVPI3hc78mKjFut9mxAkNTrYPM0txkBR395IjrpRmKfUiA+Bds1fjPmz0N9
cgfRkXtZN9HiR+7IJ39EbdAp2vgE1vt/JE4CvYwlTbWlvVkTODHt3Jw4HOiOtbZbFtc9hW8v+oJW
ujZ1iOX1WmrE68Hz0g7k3kWPeZld10n6oOzKOhHjq4yF7dLM7LK7MBZabGIU263uk8DxZgu63F4v
JU2EXvV/rZOAWyeBgz6oAQGGu0XI3uh7AbkSzSgjCm0+tRDUszO8qv3GBT0FpxnJMIvjreNB7gLN
VpICeVQv2DMlISlzLz1Tmg7kbePoBpSdXvE52k45xLDWo8qZgdcnxN3aX/JcxuuJ01qcqFcFY6uV
L9z7RwFNq43V21iQ4Ccj80ZdBRr2dmPuObtB3VhVUCHrhfrYXhWMVO2xUvSpTpB56OqeZPYPgE0i
HbiGeP46wrdEsO4NH2PMp3YcbPJDb1J2pbeLKvE9EQzA4rGQTZ6iCvZRMArG7Vpy75ZyhjAjlDvj
1MsWZoYGXMlryWJhlVQ6Imc6R3FXfcfajzSybdBHM2Q5Ee8HWAhsxEQVJpImnBlGLc6Oyd9EbWZv
7ZqQI44wx7utJgbtk/3LYErM8YuSOl8Fomv3BrhkbIga8T4O6aK8CF6B8wZwfO/W2YHqclmkRY77
TLLYIgufOL7N1fO29eFIfr7s1u++r8EGbdgeefkEaPeVkFTBgybosEpjcU4gtqr0xZJPlEPIGP+6
vy3JruviF8mikgbckZy5KOzamW9W6JMrUysSenLLLI1NZIdHdUDrb1R4VzwfD3b64Jcdo8y2ZRmH
7VhYbB5vSnLOrwjSbKvvjZTf6PR0wjcp5bysZfz6o1/BHgQMaK/HES3FPdc4MAaJ88UeGlmWouv1
iIHGT8BddCPKflZMaTFbC/rJ+EspdUeqHUIkdykVKLM1+a2J37nlypEzXSNxGsNQKZxwgHayJhkv
BDB3YKGOu44NIp3wKMpD+Enwc9psayoyGn6E3aWg4yRf2oTrNyPn8IubhhhiOVW6iQtKxNnFDGwC
/gIBQNtatVFu5413lZoVb9dJev4fDHJBdloXnpmOlJDk3+ThdbeV6yaAgbS+wO66pmqKFkk8BZPC
U0yLRazI5f5f05AxBfKHlhJod1UNXQYZstWJ4jmAPa9FbPAxBJM/i9lIxDYRTx0FnYV6ZiuUS1mC
I3+A/o8WL4z1ADCTvpawPLpfCD+ogr8BHXIUPXk1ilXxGnrfcKz9ULSRoZujKuatFLfslds8G0KZ
GpwxZVJVbznKNh/xgr5UlJVzcb75V50H3DSd7ZbvxVcAocVuWbfo6CONwck0wDPfo05v/dmOaJ9L
hSe83icq0X28GvkOnTkUT2NYATxItoYeCNVsKC1MtVuQy2mEZNkbq7/PevGA0Ggbh/HXL0U4rGs7
W9MCVDYugdQ+JbvVwo6rn14Zzbm+nkmSvXP5r8G/CmwPZVudyYRQC8neZYj0ymf1SkCyB8+qSkBF
rAavwtHqttpTM4j8swq+Wuv7br2eSTo8eFE5IDCwi1/+xbPuYY+IWtQlQo6HlFd4ZXBCHsIKAzrJ
5i1Bchxts1PxoSYfHVRLI6lEk2KHuKsf8mUFQ4rZyEUS3QguQejmG9A8uydrh1WQU4oYjihk3PPd
ZYTEuBHEnmKsVwLxwXJR0Z3ioiPB7ih3eXpzWLCC4AUPcnF846svXm3qcXGpgUu39toYRvEQBF7f
DSV8ml82klVhvLn7iHuZI65VKgfaVaQ3R1ioR0MQfGZLMTO7n6pftNwdGIFnEWTo5L0b6ssnpAwZ
fmnrJPWYH3TcnZWGNSCOGDCmldG/+CpvtqFMr5la8arr4vbuB041qAhYhPrYcRin4Q4YZesXIedK
v1Qmr5co1gnKiyTKTFXD2KQ3GgR8YLP/9mHXMkGc7CpnRfKd8z5RVssUklgpn19oCc2O3d6kd27s
92HZLzzFtzn6gKyT4AQfLUzMn37XELFk1NM1Wo7sExvU6HPblZTHKXtvWfq0igPEYaZTvbf9wnO9
eCyT6qY3PPB5Xl4AioAtR3HRA+EbPeUmEekHBZnLCAd5yKR090FcCz/xnEyhHJyfW2fe/LYve6B6
7eGKhNNb9sneWFwB5JoR4vxlrfUt2PTX43wmIhXDtwoJhzJ8CqONRMl9S91WEjFMhuyKw1LqAEn9
II/e7hLp8+fZtOLxCTA4FJ3miL+xFnEkgke8iYGzcxmtXlwWY9B9Z+JyvxZDB53IZpNVsxJ4714k
SziXZOjyTCtedWACa+nxmDaA4jrBCZHyIblnmkqPX1i+hwXcKRF58B/RPyNasKH9EZutYRCJbSEe
r0fJ/ErzCmKfK9dDwlo5HDWL4dQGBLYjdWsJzWGfJDRR6NqWBcbCC/pizhXb+e5u9/xiuPZh7dKc
szFxshYYmbtM4TbVO8rWE2yd5+g/Ddp0Kpi66Pa6Hgb7uozBO+I2UV75weGiXjhiQFa1i5dm9g7O
N32TzoTeGFk5edDXm1IyaJQvXXnb9yC8a4tISzLO19NIIB6PO2H53gIDq8gRAgo2ZjdCW2sAPGJP
Jg1tipYz0mdG1KqPEmsbIdXs30oMdNLzY0OrhAz0z0ISZ5gJvM+dSuuuZ+eLmBXZ56kvpZ6cvEJB
uIIKDtTsezD8jwBT7AhvEqolhb5LaRN11G15H5xpPzznlFmA6UGytGAP1SQlBccGRU4/9rGo+v6l
XvzNsxzPfRA2ddAiLfX6GooVwpOZE7yiE+1EN924EN3jbWVhQafuYo0rzS5KZ46UBdrA9l6/2FDU
5YdZgB5I1a8rTmUrxBPvMlGNUWE+Nsq1d0xz1gWdYBr8T2bcyzdBnihCPvs1b0U7cDg0yI59Td9E
+VX6dol/pdvMlfBKto8g9OCmFbQWPyTvxZ79veFANhe4eoHDUV/FV9Wr6fGb4Yet8k0kvVLxcsLK
dfX499Wm5xfArXbundK6ZoSGk398GOlUBKWVOwEHOdKaHbMDYBlXvdzWxGkC7o73yKEBwfuizPpy
ZmuW/x/KkzJeJ/Yl+9Z9uMeG502w7HDk/nxSmURvo0qqbTQsYlQVgKFUfVeQjosUVbXQtQqYpdcm
QWSy/kHuWzHnVXoQnJk8gdKou+Mp8ac+hecIcsWeucY2JZMbOlaIxfOd17FIJ4ZQ1ElwpCv7xz10
Eyx/tAOZJUTe4XQqwt64mgmpCDcIzU9pmQYNm8N77e3cfRBMgckFM4jeccln0ZK3S1N1LF5NIt4m
YP5RxOkyqbbVie5TNafj6D5Mr/5wWmXI+704horHXIOnqI1m86DlTfZ4Vv+RXqEWfQMVvtLXILYV
zC9bnUlpLVTk0HMGsJ9H9hVBaRbwZuXOYy2wI65lr9z+0NkOnuuZsJSflEP5JThXfZ/nOhQK8xJP
6vfh3sqvtG9+ZGlUxJ9iP3ZMcZHPKe4oyyKQkU53OuYqAOqPLOqyE/I337vK0BnzTl6t9rIvhIm2
mEQJN6ucWvU06XMRLtBvE6aMQ56hiOoZO6Tu1E/kS7a332jButiXIkjb+tLXA0+SOcsxP3kftXRH
TfdP1nPl5TtrgKKiURmZ1L65iiJNR2g/+fvO/ZTQDJx42QGY1MNPQnVREolAHLavz9tBJhuwpD96
DA4MWE88Kgexvz80UbQR6A0wEj37UoLjbtPsz+S8k6qqeUlLKyPAbizXQBcpIY25gkki8gKdIEAG
Vr04vn/YTxwHlpeZdc4RfqdqFgHpHnochmiIHLSOhIUL6c/31hC/GJLZ7V7BsLv9Rp8TAo/c+gw6
HpYC6pgd5harGGHv4Ah4sqLWXOSuBPz09nkG66V8Z9LikdOlZh+ar3vxkgObGWq4EOBMR79YLlK7
jY/m20GH65q9vqfuwDfleagzChSGAeuKLZnsmh2EzIOuNM1jw9PAoaOk+15bjqsOJgZaHl5qVDpy
Op4rqDmjwN0LLwkE9CKRJ4mrVlnw+D6NkthiXkxvYmVqgk6ALIpLHLNhuLLT5vbmIEm6GtK9rbyD
jMcXiUCwtoEmOPxCHH2A1w8HuP6y7T5onXHJtSg9SU6ce5br9360u0OZ4IjJ45NhhAD9yjCMKQMK
Z+ZQfIj/OziBfQ8GT8cio283PfJDmN38KMC5n+DiTVY8aCe1iqd5v3Dar2HV/JHl1IsalAj15yxP
+cfLLmkbqn3MozfyDNKd+NZK0T/L05YD3uMJxgWna3IrLpLYAOrJZdafS8VqWsz7q9Ohtx+2x9A8
ac5zaRmdFAFv4PcMl5uEHaYVuShK3XiLqFFjc25lDf5xNLxKZdkznVwHHpfCffh4OJ7s84gF9DVu
Y423Lppgp5FdxzigtXHw1b2GsWUk4wMFxdblC5e1LouR4Y1tg+FktLEicJBGysQ0MoAFy7NzluGR
HuOEgh7dz3Xax8Ccoa9N8HyCpRbshyCwpJYzZpO3LcWR9ujqUOav/GcnvO8ZHLgIYdoqhv8hhnE8
nZvE6+THVBMjFNkgnBej4LeJGHH6IUhgbUjNL79Ig8xpnRyTwUv2EdbMfF8ylb8hy/OkcDnK2zVk
iVCWHkzhyNzr371eVXSfyJLZCHblMBnN1cj5uw7MjEmVcQQyASiR1B5PccDxTyDZjW9KHRopIs+D
j0DZIt+zdN5lTKmVq7QthX0qs6xLxEfU82TG41srPimPYjd/BFjTLWLuYZHDhwT4yveso60ZVi08
3Te1/VNsBjV/sgXXb7X2I1y+Pn3d7oqT9iiTxAOvtZy3E+CAXvJUIGF+D5alKf69T76bnipln+38
rTf8rALwHp7kzrHGLK1uHyVUfH9K3V1m1JmId//sEyFuNA1BRQd4cLn5brkasoPiP5mbCP2Utt75
uYnLXWtcr5iiB8DIdzq/8x5YIbCVA+7Kq+5YJROqzFgkFlB8OY2JjgXdGY6Q4iNwdlwi8a8c34S+
KDPVswMiXtXTb09eyVyKQupFlPYgCtDDqp7BGmzDtTjtCsH82RjUkPH33RP2tGfW70BX7Ak5r3fa
+dUoeAYO1fOQ5Utrd7h2+6Gq0Y0TE2lYpwD+P4nDux0Tfjb4hSf7n5E0y/sCcH8WPzULL8c9nqdE
JYL+rlL30HT+EzMAxHtTknyVdt5PeOXso452ssSZYozpEgYXcJHb5/qyKAzbcI/5MdVoAIYMTL+S
1+oxzUkNNXyjfsYUAIOTTVOT6HY1r4xQAa5G/UhcAbSMpQKLkh2CxFmjF0fnQdhFzdEw7H/o3eYc
xKSswiUQG1b+YZMpOVarreqiJpVx/Lod79JFccACXreS8SauEQ4u8+O57ctzKkUuuTXSlt3OEAjG
80PJUtOMZ91VZkt1uz6HJdhKTrdcDigqFiECK4CWuf2qv4XLl5uUf5kCJKSgB80cMZtJuDMv8ZYB
KS8h07zzSfbjrDQwAWxZmJzmECw23ia4UvnHnsGhnlNnDv9+WBhsTUYluwtOHTC6pcl3Tzw8TSkg
JPFAYphWxPifyt4p6if5Kp0m+BBY+RMxG4MItAm3UjT5N54s3glsIXKGnXGCgSSTwboPhxFdMG4Y
u/dY4zgK/U3ULb1BYWEG7C8FXuXxkBhP5PA+Ovm7UJOtau3qINARTDQLogK5nSRBc206IlVj7gZo
LHOK49SwLHtWvPIRDGpx8EfQ2lIQ5NzC+Ru6wecCrd95PDEq+I+goFJ6j9M4j/2HM13vGuhcNhPw
DJyvpGhoabXjfaJ0EYr0hZm+dFXEH3A6sdIkvzaEe7z5bB6F7c+mMR84bpbiWeXC30sd7PGxlC4S
W5uB7XgsE7R8niAQXFeKrDOWBIfHBh4X4B4FZaixy7tA9g3bOO3BDp0PYRtYDNu5JeDtAZ4f0S5J
+xDkW80GeXy6sEJHSGX7lYNCj7Cr0fGgAxI5YOBp9fmu7fPWnGCh+iTN+Fhjbi1tC1tQI+GYSLiw
zZJGUGJNvMEEo6VXYRYv2uy2YcZWqVZUOCGGs4cCA9Dn9chjEtLOqFb32NuI7anUuAoXuyen2yTK
eyQ5w5Frw4aFy66dxXpzqAfajD/ZSmVdK3okVc7AmjsZZFbigLkGv19h7DGl+C7iIDnenn5Sr2/G
yo8nolazHFbbL6DtZOK7GdWzTlLYtyAEvuYEAwElKuaPEvy+jefM7iS6BKPtwubNc0IsTnixGjqH
zgjmUXWQbxIYcsB9iEWyo0jwTC9vPn3KmkQWzkJQjA+hU7Lpox1ld41jyBqg3xHKrtdwaMOYzVzO
THNDxEGH3N2nEqZCBzZScvqOpyKhZs7Dtt//k82BedWtDZli8+4Qr6VRCTOobQV03SOApKri6rMU
TmljJ0it78htiIwiJpEWIpXmyAKznHp6W0qkcYF+Y3fuGFLRdH2Pc7FY/2vTlvFT2FSISb2f6Bqs
fQwxHTHxzKH/1kGTrwysFfVx8NrkLXSGfb6kCKzR/pvdxYdQOL1hqhPJcDpX8EVva55ESBApIt2f
pbyiHMbjqW5PwsgPcpGaqYGyQjpvDbiUgV8MMu3ShIBVoj5FDU3nyjafNloM5nnjHR3BwM6dZmSn
zYwISovFt9Wd7lNlwbzCwlwnhjc7HFQ9r2U9ORKfFhZaMLpW8FOrKe8JStDC2SiBlwDM/ZUbd8uq
vw+NgMe2sHna/cNp2qHKIqiySbLkxDbpeYSdax/09AvZejzHNJ6wIiWIDpd2llawQRuoSYC9lpls
LFtUsaKSSrJyTxFc0TgZDOBDSkn2kfZBRdKNPajWQIAIm5Ck1jU+5E5oL/RNnObUAvdSA2oi/774
OaP5bwAc8lb4Z+lWVUJX7pmrS8eW95E/iYbDMQ7qRyPgnQnQR+/nsAnoBl1JKC3tGkuYHeFY+wa6
gSWk/OEXjW3RbBwDp3pKRzvxPCH41l9JC4gPLh7u+CVTbRxjDtSVSouebHu1n6fPsb50gGIyUc17
T026uSCjtWguVnc0XmWoEE0/lir2fsv37aqWWErv91xA0sMaYvhtoztzBq4eDrvoCCeQtKeqT9eT
9AsZ18qakPmnquu6npz/ohF/NHPFuFAFKgZ7xJ8I76HWhaLbjDU3PzcNWrizzW1hvdxJCf2fQKHJ
cTy7VIp5V03G7wht5ZYyel/QO8Szwjj7KZzJ15TrYNxD8RYjkFOcrOxmy6SoUrqk89r1J6+TlWIv
ucS0q2kuyb2Z7sGa8KBcKK06j9fVcSdOCJ6gaXLx9sEZwMmcCTp+DhCErqa1dmL8gS01m2IRHUmo
uS73uTZkjANqRoAeU/jw/u2Q2C7iFNpSrW2laNcuSkTZkD4pU3k//OOq/8VozQufQ1tgHSiRPe2G
q48Wqv3dUUzAz/KTtEKK+UzcrDxke1zytClejUyKFveZQKe+EwHrDSx0uZoJa4qqWYG1Ykv8L+SO
AUOIn2ZT1qP2x/M5QIusngoNW23iQ0b5BIKfkEi19hoTegSw9dPjfkU4q/KFbarIWJAAiZiAV60O
6o/Mq8a+WnVGjZDoaIpYi8IM4WtB1IOgax8gOzHwkOO6RD+co2iA5/wS6slGkzTTQQ12IrYt3hWA
VCjjexlAq2i/r7kBSuh/P6ctnzYDfb4W7A6c6dQVLcBGWirqXkb/VQO4Imo9Up9mJUgHQTQqVM6+
TrINqcffTot2E3oGgJvHuJoal1lUMPSkc2wR0w2bM8aUAtg0znNdNbp4rtEoV0AgW40iG+KkObVI
4Zv+RhUN3i8nUswS0A1Qasn2xwbQfp70nIV7MsoCiWu+L8/RWNjU5DRyco5uYn7Woi4enXHSVIib
KYjGhLk6XfeR4JmgoyMs9AElHPh9lCN3i+R7ShGS21SCYEgSj3Y2P0GE1cCgx+4x3MMt+yDW+Bp4
eJAFLOllG8hhEdT+jc6W9BwZEtd+or/DQE5KhYMl8144GkPyvfWC0bj8iYLUo4Hsp1AoO51aJKEB
ZSJYzqhkVJifgY7GM+oL2JNVhWjCUe7J9iaIUG7WU+taSJKOC25oIG2nHDUH1PoW+Un7dnlgBdWc
76srmHxx0ZlQk3tS2fEYHMXnPe/vK9Q3uiISQSrNphmucQnpvUC+W5cug9byQpdtSSA0i6qkuNXu
oLAxG2I+89Zb2rNGc25locUl3Q4Vhzd4oQMng1n4rOezU778Z36rvyKeAjPvt7Xlb9cPvgVKjyuo
WevJUeUO7+Cfkmy+Vbxtal9E1SdsA0YMdsnvJ8185C4OUobGfZtq3zv5pf/A91BNGXmOd9rj/hq5
2hGChw9DxQlUn57TlUDHTDU5hj35/JxEu8tA4n/LVTtHO0Vmdfcw0SpBnVgEL7pwJyPWUyT5QrjR
cKETAtBQnksi5GwWRy2YLpqQK6ZFd/y+Xm1xnWpjJk/UX7rLwbLzYvHiei568Cf4RgZXFwpzYJA1
heZsgHmjnQemeEM8gJ6FBfyTaRJr2Tb9Vubyu1HPD4kEK3ime892diBWJQh8aF3dK8TdX61xACRz
By50EdeaJCLDBjHarGhN6L1Q/cmzG3oM+vZBh2C6KZxvmB7LogFo4M2Y5ovZUwAkeeKGEPuL8pdt
vAFqpUTAZ5VvXwcA7UERUr4iqGU4TIfk4Jtzgq6IwLqkY6YiA2J7FMYxl7JvvJENK83b+USJI/WL
YM0tLeVEBfNlBWpBFlM/nj5aMRYCFe6J9L9Q2fkwcCAiOmKT+BZAQOWoVPNeIeQ4EhJvPpHb/RnX
4kxWTL/HTt42iWvZAOilwAmQwkR8bn5BPLJovg2mM3K2xIsgULYlz//t+gRnq5VV5jNxQ3eAcvba
qiNtJ7X9kpjNKDYfoycQbDFTG1WRCG0b7t1lCIYnr/j14jqlXdty1s9FGgg3HIj9Snz8xvy8GNbI
qhfIdvBTG4vQp2b91gaU7/K+1L/c+dRP5AtBtFKHOB61sreHHkCvudvSnkBTcAAoQ8+DuB6tNVlP
ExxEyWqbeIQd0YCOn5Yc2geGbiInB9Bzw1f++GEsPqCErguPhGS8JJq/nCXA+dJyQWYZuH64NaW7
hg15SGq4f6zWYGQNHw9+lG/neEz8ILzbBvu+Ls7181JyqVj7+DH5q83G7s+9D2BnaaELlVuBX4rG
9prhVO/Nc0X1tAvNFJpl0tzUuJDHIGaE8GBD2zubsG+KiIneUPlpWJku4l5w2I2D3Qhh9ul9rfVs
1YPaUMj7ZE64nir89KSXfa9j6O+RTKHECrCYNF+yvoKXu+Uu1cRbddXcyglLGRoIrKEd8O+5WlK5
zaSKc3KqZ2nfTk9XlC/ueAQKeT5I0nPkcTZE7gSS+H2nCvVyqQDCeFDIaoX6gUwDCY9jlM0LMTOG
fGeO2lQ0D7T279K7kD48SY6dNnZRok6LDc4z0TtvBPisrdhwH5FlVJSSKNvJlFdWftLmD5Ip/52P
KZjLIEEWa1wPUeHJxKmRcJwiSzSooH5r2GRajRoItu90kAPMTQcEQr3ePtFdISc6NyA0BeeqycZB
MZ07AjRn8mxGkWU7Mq9qY5j0y5Z5r152hvipXZw7bTU4BDkqhr4X544ehei95FWxuaykMsHRLrIH
5P88bN2hki9ptXU2j3k7/KNFk6CTAwqlwQIgxZ/t2TyTcEj4Flti+fXmBbIB7TiG5aW3+F/6nENW
tNXR2k0rkTR8iWNx+ZKXSQZdH29vTAkE5peIzZB2wkGrxjrm0VFcyFrIBIrmh/n2u/IVwaVsN226
lnSdWDclZA+EZIAZV5ad9IT4bQEA7Op3mvEi/Mr2ed91iGpWXNin0qWSZ4/duIDaS4LhemGtlTIV
joFxQaGGf80vUMuNfSNAl7RtaLTKNzP6YWdMzE5/3tg8zsP3SkgbzdSndy/+DK90cZdOHpTlwJfb
cWxuEvZacSMHqsq91663b6Ax60a0pcYyDN1hXfTk2mJQEva4Vd7ASNZ9mqOMQIyxlbtuLRAsGV58
DTr2ay9Grpp7L2EgH5iaAoyR7zfl3mQm8aV6tBvHXh3GGk77wL98YRrkaJ8rxwgflcTAnOkWSz6f
2N/XPoUozJ+z1T0BqrQjg0HRkvG0GYaURQy7Gw/S+EIocevKumihJELZ0AZlSZOqfYhlAF1OFxTl
3STDe4Pm0UeznP8TQ6+hoaZ3M93mqkjynhHkTQElroaXFT70WQXVHXBlcUjj/d0Kc57CHWoTg1dD
TOOYDRI3Sn/zMct3x6Z9INf1oACYbSb/TD5SGJyY0+Meus41Y57R0zoPGBnFF3PH7mkQNH6RbH1S
HrVJGAmhUeRp0PBfKcyvT/oU36MTu+OIG0/N/rII2ACfktnHY0vaVTnjQaU1/4mitARIpAnX0dEK
l/5bdPuZx+4g7lafKwkkbrjOochkuJBXyQSoySg/dHoyw9ntKnzxv8wRWQQqdsMjqZ2fOjZJDBX+
qCHZLFcNv7GzxsFuL2mQyEli5lIOCAxLDG4I9DntI1YzxYSHF6GWXg/ukvs7z2H13ztMP8VdVUH1
0LdasHh15iRqfMjOppSdWdidjGh2uFxvOCtljV876ZPgNXNFW6w21GqI0v+fzgK/iQilUqjB4+rx
jTyw/XNxsFRBc4y3NvURVBDfXX+hqF0jcBdabgkiSGQdPNdvdVC/lSdd7x4imo3N/4S28hsgM9rf
efyz6tLIMmUgtc5av5wBD3vPO6qxqHNJ8Cihzexo8DnVtWfTGm44VCp+qoS8oSQ/LdWA6PBljsi2
gHk5Zw1+o3hsbJGEOTUUWh3xSB6FaTS3YMAMuBn05YRb7fMkUjr5zUZ1itl3QKNPi5/5GT1ppseN
7wLP4EXEu3q+7ZDJzaLxmXrTUwB8JcRVD860Pe4itr/rypEwrr845RCdu8y76bMJxciBvqJ3tMd5
ctdp426jqPE89Sz9Cz6CVBMzke3uB7mrtJlRpDIefF/6ctE9q+vOn6xMTH6Mz0Ux1AyA2OG6K6ia
ecIRfL6kJGSqgz4cKZGRyPbCQ3Ove90qqzglu5aocun6GoWhev4kfWVJxiQ9KvQsIgSKFTxmYCgo
NRnNB4U4SARvZ41K11B68l88tAqRs+jRIPITpqWpfOOoWajV62nA7SKgTespv7Qk9hEH+icQj94Q
9q8AD6YnLvXvElxtBlLIvkg8y6a4BHU8YL/NeYpuQVhU27PFRgx4UfX50B7uCKc+G5xVq1Jp/ic8
xZBhCiZyqibBTo/NEe9Jm0x78rS+DlhxS80K2NhsOYcx6QYHIgnm2qq4UeCBrm/OpSYdoRYfcVm6
qS1+rnU/xlbRj7MUqkMnAimd3T+J3lozjYhPLLsX+AUWDlFM/EOfuy+XDQeLtIl9NyEhgjaJ7o9c
DMB8QvP0FVNH2XlO5smEBR4CV71p/k+WI5ZEAvzCVW1UpFv8YJDJ9aQr48DmM7HrHZ8MISnW01V2
XQLqokn0A2ykTQf7X1JIxLLshUNiKuZAq+YsfAT80nBeJwS6oXkO9uidzhSjyAx4D8wwcaQmj4Nx
v6ib9IxmwfUWX9B6gAd6/M1XAoYL3WA6pyM/ND/uxZrDkHkcxWiwzG2bXIdgCKvAhOBLB735eSI8
Z7bZUKSTpinzsLLDYtCrikweqg7Y+xs7MG4An29ICn7jU3JDbtYPRgLJZrtb2RfYCEbQ2HZ2hNQn
M38hTakJDt4KTcKdbv+d5WNzzpRTVjzvIgrtbjmaLL2wzWVgC4agyM7fMwrewwt3Czw1N0tUEtQ7
8+7VPpjnUs21vD1udkHzyznv7G8gYz+4tuSJ58W5AN5glDydNUdF+3DIX2M0as+cT7msYvibWwpv
4PC6EabiPXmwrhRi0OJSMvbv82dgcCBmkmIGm6mTN20qaMynw0mjnjmhNuyd3PPYPDoxSvMvAWqO
GRePdq4XDkVMu7r85AGXhM5fi5b20Vhm26Z/5G3KUomhO2u843LSbQbRwg1zcOHxKDcs2rI8uYXu
N8+MkxtHVkINC4i9MQqHDCLIq97rTYuBYBJXFfwcJ86/+KA1vtuOJDSWi4954lGqOnKRmIKSbdoY
5v2s6bd4+FTfypjUqzv7Ax2J3laJMniHK/ZZJ3mg0uPd5+M6P6CGFc3iEZ+WU+j44O42FNBmOpyR
dArPV1pKl4k38BCbccqrNTupaa9W5gY8xbaclXYAVj82vGsUFIqzwvuMDQw7CqozJCmrpgYDaVbK
DhDUsR4aohQ77nHH62T027DHdRi8aq6i6EuM1C3QueX7dPkOZAGA7iMDoJhextf8WBS6RzPQPP+S
JAEVX+wR7iUQoGJhYqeyrwvJh+FmFqx9kMBqWFIGABEwO5FLkT4Hfq0kOf/O0+Y1bde64u9b55nF
eiOFRVaVZKYf/TPjOEZsHg9ufh/N2qP9ZnrLS6hltiLqsB1YcszspFPqG7EwPq2yU6hgSONZuTbP
Oi/5TLsnh+7ajYrGd7DET/2pZxuoiynLt8zHmk46duXz3zmmWRq1n0VuZthbFlv3dnLF0d+tyalb
xzyUR4rdAPke52tSYfTV7ncFmUuoE7ljij+WgAGnWEU0L/H6U1Cz8MRrKh2E46RomSSB59QfRQh8
s3+uDZ96HwrKQs5sSZ3Td+XdazJSnvrzx4DUGWvNyqIBaLVyBx+4/rCwPgSvGm723+d9jGbe0bGz
rt/IrqqbddTyKP7j+97bogJ3GP8o93i8DuTugkvGX+DcnIUpboDszZcT+niWHVE0NKtgEvam40DA
nlB+mSs4YUftyXJZDQYyvqVnmw6AGKUHJMixNGukVFc6Kkp/b3o9cuTnrfbEJX2+JlzENUeruMom
s5cNbf9Gi29JW0J8HK1qzrARn+jlrL90uN3Kz4m2dZa+pDwIxdoF+JoJlpqw+RlWly0e2ZrawSXX
CsMUp9L18rfdClurAkv4QuUcf+hyC8m09IxLtzw9E2XHuPJ/dZdgooMREJ2pkg6Y7a3aH0dSvwyC
UGrEhA4EsZYM7SivsGRKdSLtbjnUc5svimXth52EuUZu40C9n4YnLyu+XjERBRqoBmszbxnfizUU
gebd8yJ4NBVg0u0MOxuKZH/4wqs8ReqID60yl2l3yXeQuAuNKTAhDoXmJnP5xXBTe229ZL/Wpj3n
Uw7wS6ijxU7zKcaxI1LkZTSorxiPmfxZteg45X+9UHskHp86u5H4tl+lJFwvTHJH/LIeSSezynoa
E56F57ybrp8+XvwrHAosOqozxnT4LFSxooLLUJ+9YaHPNG7lKDlQ13/dgccwIfs7Gwzhv6adMcgK
VwYozQJ0LBYak6FOJaVh/0n2sLir/X8/Qfo5pBUkX8+mpvPwP2JKy4MSzCkULsA/qxhLZ3y+CjQE
iY15Yr/XYYYeL2y73uIR6Tu6M8JuuaGnj8M2oH14DdQLmZjAlTCXsBYqHRF/zxbZq4femjNRAuW5
aMs6vmGhgrOBstHoQ5eVpnGQ19qIS64rKloncfYtJh5X/+bV5ZV8oO+UwegsAxymNXMxkntqyWfq
rNuH4nxb3U/6maGYfJtkdtIQvixpXEE9tU/OE6M0eLOLJCd7KGEhswJmZbP8ovgnVzYcfQpi/NzJ
QHMIEbpTsOXzb/ypNzPJv4QmDpQxz23bXQFYk+K6IRheLjxvn0hZkofqQtyXckZru81b3F2qongn
GNf38gS1EBMVTiPIzmDOsVPInyKrUJkRjPrc/Gnx0PCxUR98Dh6jmbv2mL8R/GmayvZreO49KFDV
uqhagA5fApCgLRFTi0l2DhH69G87Ug6hQfjz7r/kJThmneKUir/DZn0jB1jBTu+R72g/+3zD84HI
mQ4G6bk8U9gu7SzguarxB6UYNJMAfBi+ycuW0XHstDpy+oDzVk840wSO+wQ+mcFwI+CZRV1XMrxv
z2yH6PHB/HZzl5v5GiABP77xn1It+599tjX3F/0C2DaOWwYmJv3jM4Nqy+wjgkfDHHkHNQLCpd76
KZv9nwXVFkRPUK7FQN9UDckpfwoAxuZcUOK9+PHMtWDWdrQz30coZgyxUx+Bm4c0bN913zSAQJT8
n1gaeJYe3FTSmmgNNvVOD23sMCY56ka1XTGueqcTAL1mmSzchXdLS2URatz1eax/IJ6vdjtNuP4Y
gew4FIlNsal9hFQXZvP3o4ZdA2buqg5gwebq3RDcr56RGAA5TkIPfOjfvpBcYkponFJkftpDWLx4
UJx7+ovH692bigFYBOaH6nc2hR36NFJlr4WTz/loGNYvF68LM3WTrsyoS9diMlzoKO8el4eGYNGR
AZg3KFoFeJmqReCvQtVhmdjBYQiWeOepNVa1LHzHwDvDM2vQWntM8iDxpuKgNR5ohNdDO6hPeS3O
5GyZ92P0z6VNh7CME0uOwRLP4zPIQY9/J4Sjwx/0trnQBP+PnCDHlSZrfzhVcWF5PA2cyYvRUUDz
/yfXqoBgveFrD2oVWkxAU2D/nLnt8n1g/9Q6JOKP3/3hR98yM2txu8bljFPxC+EikVLPAZ/24d14
Gg7JBxGrWAcH8OWieaMpOd6hfSv3uZdDg8RfHVCn+1pS4nHV+0wHpHWl5YQHs+F4kpELBTSh7IhN
JMbgQl7Q/I5yg+5Nz+hwUpLNlql+tvoMUMe7pfPq3baxB3kJiEmLeNcuFkS6zWFZrU2haI7rAmaa
zPfGrN/zM//ih09QlOcXqz/OLfjR7yAk+uItDR5rUkUQT49LdBwHsE0ARtyvre+DLKPv/6EmvBhn
KsqJEAdTd4BzehW3ZNaf1TSVSVrRlGQ05MOGcV4pwoQsN+qVTr9BX5wjH/DKLt20BdxBiRGk5ORQ
/UjSvh/eCMQssZ88u9SwDtd187QBysApRJcLpRlqPm8S2NraEZ1dOQJdohjSrj1uAkEMHftPTVs4
mC/d5weulcKRJsa8LBIZEhApQDQBUeZRLUjVkJqBRva1+U9+YvXXIgmIM4ICy7p4abL60EZt6nUK
28dwQMOUYdZdl4j5D43mqi5NOy0RQv+W30q1J0YU/f6MR1i/u9tmlqRYd5nn1NnBSIL1RMVPhMPU
9E7mq4+Y0Ue8ilRXycHX2WIUFoP/s5DN8Bsg7hshZ81FxT3Wok6gY0FviVcRE61c6/NzF+WFRSbH
vYfQcj0D26302FCAoyg+qTdRy6s/T8Z3RVuoGUmd5/npdY0NIkWcv4bxYIcbR0nKdMU0bATLORgj
JB8pwiBbtSVfR1xIj8hP2RpMChOxrGfrPcXTqnhrN26LCwbgPW1dniNJuArpcPXAD93NN6nHrDPy
sFMarzBm//c+XMD3MjnIisqaQ0cCtiEDHpRfFooItWhphRG50a3N1bKoazysJZllXwc5E1QnuRgI
8xhmjoEPTku6YEno6ZnYE09dRU6JUI1Cs8+kreEnBc82wY3r+5z4MEeXSy2KLi/72xvGhMjlmfA/
6WPSr92BU59z+VU/gKG0SfP0IBKXP0ry0PIamgTN4Ov+4zg3OvUrDiPkI1WSvnvfmHgROD6K8fuX
Ha1QcYDHXtjprPY/KTc9ZdlZ8Dj4p9C3IZ9+xagb+ZC54wF7zCLd14iAloT2RIs/Bn/tvxYJHWs0
QxAu5JRU+tu6lpjS1+7FdXSS/uV9E/ueu7E9BQobmUfvbKD37bDV2QxIxplCjh0NGg2+ZzBLgpJZ
g9cGbrbXYuVAy3Y6BLWUAduCHOS8bW0Xh9nyv+Ux9vlwb6bTtv1vYZIqt1+1V1psy11HjIuDqVmY
5Pz0XgqjGQdanB5twwPf76/sS0RZiEgf+dxs3qiYsPGx4jG15TcnkbMQ4igrHC1ve8Nfe8hSi5eQ
FuiO5iKdc6QzmAFZDsuL8KIfAxmEgtN9zq08q4SJDU4+0bVOTn24Cg9cWTiJSfLWDvWo3SBvtvJF
BNTk7ZepHajelyDTCe99v7pKg6RS+UJNMFU+UZwNPYW1iOpVoJyoKDQCjoCXtaIDzOLlrj7TRBV0
+AITYLyN2p9iqrP6jVRJ6x/Z4KlDd/KJ7wOtZbAX8HY9UVMZmsUUICcuCH9+ib3uSQkhcKPDx8kX
F/pctIOVxsDaX4xTDOJV6F4JZCNHhSFCWE40oVGGnYsGT8whyhzRX/j+49SRrucgxhKqLxEhIxME
w6a4OAiHhxCf22Z689fWzCyK6qokad+CvXoi4hdRPa0EUrHnwu4GRi/D7AfdK18jaNBHzrccMzdv
JdisGZXCZ1XDhzsnz7Tcz5bjGpkDZsFkLTaxgClTqLnDRwexiic+VKXImNH63Qrsp2EqOMc0vZXF
Ny05k426ugKBXFGgCr6JYrNzRtUUUYYvDx496+jgQYVQNdL5padHwPBC3M6kiTSYpb4iSFvBhsKe
PkLu8lw3wnOTgGBf6ADuGz8WxPDwb4C8ltFI46wOtLKpmBFnQN6hWKvIguypR2FMHONPGchl6Fuj
3KW/xN5m6uzgys8NGFmMcDn2BNwi2zp9onGs9BBC+/0quydgCnh6Kuo2MSflya86uXgwUGNBeKMM
AwWAJlhBn7Map9p2QCkqCpYPTokQtBlftsrt8qiWzT7L7eD9FQueoeVeDsBNzCmQ9UVEEMz9K7yU
bJAEwSnIRVMh/SpA0m992omOixhtOlYLyIbj3smi24fsnYFtlnl1d3EEt+d0CfRiErCnaPo+PbQE
ZFfn9ROtHYcl+qnwyPZxME4YtTYvQzFVsD3J7i51/oOd/Bau9x8wB9/PeS1m5I7V3sGuqcjlF7nm
JMLrSn2ARC0sIyV0lw3CosE41eVKTjAKpIi3XECZPdLPIgfRC5eKGKOJUeS1rOCvYYqjXY86UFuG
5yZqeegPcy6LYqGuLaU0TkxdwVWmhz6X+HDj2WvQN+pOUQx7QriMKotKY55k1AEg9ufk1wXLRbr+
AFCBoUI9/lppunh68/+MGoinaNNzuZ5zwnlzvZsW8TeLv6EfQ69M+XdU5eu8tfK1LfTviUEnWh4E
PUJ7mMfKJlWWrp8td1MJ1IHvHmZZaVgAGD9n3CVUXpq2NqNOCBciCRh8WNLhbrDtsg+Nl0WNlE48
8G+Kynq/s3TBiSzxdbke7r5bRtkfDrqfRxWXxMEsTk8ex5wn/2V4d7rpL3IUaqAuz5dCkRmh/WHx
cvdp4cSgAta+81B0BN9nTfxi8LX1EZqCPW5qAzQuyjhBK+/g/EmYT51UvoMfNju796X/Z+ktZDcp
Q+oGZcOAegjFYE7FG/pqmdsrM8IXVP4FnlUKW87zeeF+gp9XKvx0F6RDLZtG6+P0OCla7y9oY+YQ
Q8sPxk0n8gFPJNpXMI30uQRdr87BMTNwWu1VG6pssjHimMbpT4ReE4hRSxoLwaKnVWinYwdhF9+z
9eo/ya7Y8kGd2GA6etssdtHPfS36aENfkHTyDFuUt3ONXfSovv3eBhlcHv+f4u8kDdAOSNruVMt4
B3r5d+11Dqlp+Y0Sz4UC2LPMjgXfoYGpeAeaLwm0C+upDO5DY5rBiVD4ntB+eC4txU2W4fq/eMNb
UL8d040gg/hYkPUYK9FgxrEYD7HKRFjTbLqAsQ6x6pgtGk7R64bpwaXrwZix0ERm3eJHMHVb9RyQ
PhwcMXZQcC9i/lJZXfJsOwTvmcmKQoTVHnmTRemL8Hx5VrUjIC9Nh9aK9MtMzRA40uuDHBtqeuKa
23MArcpXlkiw47DAz7PoicMoNEXklZqPSEqPssNHCV+X1W+hTIpuv3mt85geWtKWrpd5x3bZbYfH
Q5jR/6eKVkfur9WLt6wBQKJa+l50W9aC48b99eXj9DjU4eYG8Up+DLb5lJeE+L+ZTT8nxPavdU+e
777uYtTlaHV8/7D7NbRHV/J+s3woJozsFLW8iYeAZ7N7KrR5RnyMoAqqPdxslW2W8dizyN5gVOXl
k1S9TpZDwgxBwyYCElnW9Ym1XYnt4SoqXqScOpU0VZ09Leb0ZfbCFSE6sA7kdZv3eqTambS2huQq
/l348ZRYS8NY5SQXbpFNoTFp10wdAKFK/g31GexpXZLi15VJEfBZq3GI1AWhZZScd5VoGF0v/osL
ZSWn1/bbjGVOgnoSQoOW4A5dIhpB+rIUrveyC/Xa8TeT3vES0Y/iZF9JQRIEXQeBHf+krOKZQkKE
l0F/FwDlxaovFPz1cqGjl/7kCVfxcptNz8UMZLrScxROHexL7CqSfsmeZFKikI7+heeLAf+GyQOd
Z2Gzp5TjRjpZdHX3nfWQRyV1tJafJ0Zm/XoWXKMTkak3na4xwqsKQ4TeJjPPqaVl0x3A5PjBeOoZ
hRbBZilta0kFGmt2V1LoEzJ23L5qiIdImNE82N1Wv244zm/+a+tyGbitEHGUpxhZr5XmQyfxvtqy
OOoIl76X9RhXTE+OcdE23UqWGL6fL1TeezFD/zOI3ORPLM1lucUL61FK8JyMbmuZgyfDbaw4jcaD
jD9+ESHo9p2MxRDazzNVQ4x3lJOaxr/Oqlv28o2Kpsr9XU5/FiRFyhNeKBJ/08heoUC7TDcmM0Lj
KaEdr7qM/qF8KK+JcskKg20xSgP4hR9n4KG7wkg+vDOWWMbtH/0pWjc2wQIN7B32uDqd1RGOD0yt
wfFmrJHXMa+PwwL+eCAGP+HVpCiUwxxO/oVhWYPdLbDHUnO0veJ3tmm3MUJBtTth2ji98+9Rg3KI
acNNDbqXum0/DzvIggLKHcUVe0dN55CgTK/XByJWqdba97DRXCJXjFSI5YjRYRnVv3+oB+TpZPWx
4w0bM2iuLy5i/QWHHxf1jzqLE2ExnPSN/DqumVrcV2DP6KKWf68r6BSWpBscR+JgACBdGqSdvoE0
aeXkfgmDCrmQElEc7D6o3i/PeOEFuQwplboS9zVPtADBjnochJbgqeMGVW1//qtP4Q/mb3JrYkwZ
WMdAQUNKWltODWbmS5bMnRVw1a17KLeRXXukY/gQHbFXrH1xe1S+LjJrSNcIHyetR2bwhIeHBMvF
gQBDk/5v3AL2uW4JoyRvYQ89PSAyZWnCYHUaPE9W/HCeHg8e/P9jaC0NjnLFOY77JQkhAdbFDTQJ
5msUTtC+zGcWIw0eEmVJO9GiUZ/pIc419GME3zBOlDeJ9g2BnnQtDU9rfNAotru88j6lECoQrud9
/vvq2+AFwtZQRYqF9+AK1vNezgdo2LWEpoiVhrxRqfspUVo9DQJerc6wD66UzLmzXWcJfnw7c+1o
hIgyLSSLRrkhJQdsafdQA24nc3RvZXn85N+OAAp/7aMLUUS4tRcWPBThefFn1d5inu/gG2S+kPvf
kaqp0sT28V9qykrmBbtfESQ7Y6ogbMrme6lfRYG8j7vJHzdEgbmkhH6qzRcpzZ5og+PcRlDT2hWa
DJT6ht3+6JQLKYt9EzeWH5TdA0CAjYEmV4iWNmZGr+O8Jf/1dLLakx/KuNnTyIYfaHm5e+IrU3Sf
6Hq5KLVMne7sy2pNj3IHdmuCAczhrSNJYSgREQ/yF4mFH2Z8XqJiNRdJFSKquk+kqeXdi8gu6NJa
sQfnqDN56hKAYzE1zpbGuk6hvhXTyhHcjDTZjQyNSnF6VrQIaAXG8tfVYga3xHq3n82MCy23sMoM
avV9wUV0FDK6LsyuMRLvgYRQfdtSTcGgOXcPdjWkj3oh4OsTkHTfJ+0G0A9Sn4Je+qI2kSGKDA0V
uk7vfvxcWbDzoyqD4hsA4gtTXZDI858Ao1UcUt4Jbjw4e+ZwekwDKaEhi+RIXwnFfXHxopY56bjW
D+vTos16cljFMBrhMZ4MQLf8qXDfxNmRg3Tw8fl9bJVTLel5DWt1ok7C+TTZ+Dgrn5G0qduSfEvh
6Hb8O3cHekMmZDZ9LSs2LQFHQUwhZhuqAPF14NKMEp4Z1yp8bsYtCzEaYudlCrVmO2/UbUdFh3mp
QjupKUfSWVWzbSOiRSRRWiC9D6fFpYOETDIqLWGqdEzQJA76B+r2uviNeFLyfmV5L1kRLb+N94CC
EfccObxj9X10qHLjBfFR5ylfl2WbHFuocSLvTKkG/8mzTYJ/DBk99EP58S2tQ9TaxwFCAwY6+7n3
4CmdieOZLOv0j3XpiqL41c1tI0V41sUi0MVR2EfoHKPcuF8Q35mciPPbE0DlwbU1lGU/vEH8xo4I
0yWhU9lOybMew2Dj8kU2vpfmljxEBHXXxZvMzsSIiEfOp2+MphTGXFiM2Fb3OOqSVMLfa939OD22
8Jl0EF6Mz+FbTd7kIHcS4ioWz+7V0yaVJa7f7EkGD5L3cUlbPfZNUuksRH4ycIsKX1LFcREHNkfj
wjQmw27gTfkW+djDDxHEH+0ZLUb1SpgBl/vzq0B+tfScVme0hrC0imZEij3SRo9nDwGpWq2Nd/cn
+kKyLJEaZFseqDzFGqmlriMj1j3g0sB7IhyEUv2KI7ykm73a/9eM7rmhtnAF3USGdZSfazYyhPSg
2+BxQmBAfmO/Wr3lvkGoYOknE4nqJCP/Q9YaXlxxAMOqg/bHtmnV06BQFdkG7NfANCFLIrru0/KH
fjH+80fKjAn1FAoe0aPcAdCNGtoklITPqhguophApf/Azwpn57BV0YALH2f5tNn+8UjIElwyYLJ+
4ASZOWaPq8gkuitdb2vaXqRanQIgteEGh0WHvipg0NsoXAJJ+DLnQy+f+CPg6dy547MciT1zV/1I
fVS1tUZ0hgImTG+1u8oFIsda1lIJzLOZU6sF3IBSlb45RgF1KCi52mAUEcbThZ+vneBz7mbO8EaP
afS49AQUIWRTSKdmr4W4QQQXQ6pzD6G/rH711zTy+ZMslaXKkNMye1deV5YkJ/66io7wfwPEQBDb
boG1YqSAwXUPE5mxbj7IP5S5hkUhKUbKp30Vj5uj07aGS1QfZ//LIrBQ3+Ax11YGliJN25UDGeWd
7mTrAwIhC1wj8BcdtWtd/58ap+Co8pBuaTFc2TUImHqXfefIkGplER7PgsvL2KXp1c8+ZfPhWrve
1Mcxi8+Fafp9JUh+q+o6miAOkrm0ohG24AuCYXPtblx0GTZmE5nknJzJEokAz/+KT9u/zWb+qQuH
xwkBdw42zGv7GK99SRNed+tgc3+FPUP9Dc6TV2T1LfP5RRFbkcpyISEHPX0geFHtwkwvJRZMm+Uq
rVTiuuJIuYl27uaql2+igMpmmAT56udkeVqxGfITS96bIXYmN85IaTRyMclqHPPPwoLivz10+1qe
2ulXN1nkQxwEOCm5099x17JtH8SuSBrwxaM4NTdUJ5YbzCrBeSW6F2dhQ7WeklXJGPKg8ps2wRse
Ld4RaBXvfEKZOxdOFdlUIuz0qzVG8vRvKhMwQ1ankcGEZBEwuuIE4kRW2BXUtt2gbTxKXqFASP8t
wK3VFgO/LoMShdxoOw0W77VkKgDG3LcIZjJVtgvKVyugejAFGidZyCxdOcptjBiM5os6pHYHRIRQ
OYTekrJDHaUKHjdlskaNLYhzpWkjUNdU8DdmjupXxDZ84fhcYarjcanY8kZX3vlKpMhUmDOjZ8tJ
2o1XY5PHgF0XXwYunwJQaqRcWwO9yQ7r6PMi7IoCMtHQsTMrEZA5g8TYUdhQNFJGuBs+0aQDsz0L
nbc+ACoUEWXr2x/4od3k7d+6JmQlw5GCHr82bGfKdrt3+YkDkPygCMk3a8lYPhuaGmkztxXRcHJV
vajaV7+Tw1qPO1t1/gze0m46eC+sFZXGweUjpuKjQKclJ2XZMDbZQgfnm3HgBeinogsJycp7kI8M
pVlL02l47pmYMEpv8NE3VphxFNadycwLZ7j8tFlQGvd9/8s66bVXcHQvGZkXOo3I0tRIq2PIVFf+
Fse5QCX6BvmFs8tp7VPHb0UEgyiE+N/cS3UXvDpBFeKnMsNVvnsrUtdqrJvIBL7NZhptosLNfF9J
M9PIRbuTUCAwrTggTS06Ls936tuFBL4gbVttl7k8ULJ/pGVjBWX6B7NsRzmHFuqDFX5ImnA1rvwN
JVZO0tjTrvySEc4er9rUg1UdfMuydJ7vongIIhJXG4wrerbnBGXZ1d+ODZ3gWlISOp9DgajvjQwh
3cZ8tPhSEQL0mcsyb88cp+dL4b8pRHzT3J+Su2PQe7zxxsl0CgrGRR5eEwWIdV/yrUE2xjMQVzIN
8mzZcdaJMecoYseoWv84aA6vC6k7H8RWP3i0BcuHpzggpMNLm8p66fvke8g9CmLl+Xjf3W+iuRoo
UTw60x8S6Lfx4xgYwx3r9QFNHzCRzjIlep4J+okCymQQn1Y8+g8wR0wJH+9ZHSFhIXqhkacABh1v
LPB19wZ5ZAbT321yUjSVQFK7Vs2dlSA9+TKQY8JpC/aoBOgn10Y6VyJgNE+TdT0fqDnclzV3EC0e
/fH2bKHQhlQ+WOkOOigbYX5MzaCkM7lAwgerBPhc0rsaD3THgQ8Sjp11oj+dDtWtuGkGIwec9WJ1
7itGi/wnQ4AamSlYzDsZ6tUuPBj4eEMepJBi0A0eQAmKi9uUphhxu8hgRK9UkqEI+k0JSvp1Lwmw
qvPvyiFDygXQQgXHihfjbgxuVtoTNSaC0oedTL8+IUpoF4TSy5IhL7mJ3YLGU9S2JFI5PDtsv19y
9PxZl9DXzb1wI4sPLIkJ+6wi1TssXd8HwE7jEya2CKuxSHjRGm6vqwNbMOhrDEW/VPj9TePmRQ3A
pnNldGsQmo01A9LvmWzBDERCqKJm9b9LU1Iy9ecpsMWKLzAoGymv/7FW24GHs7lTgswk+k4WUZkl
GRs3mvW5Dk0zAChw65u0n8yWTK6BBWfQUNoJ3ef6HxMMe1g0a9zc5l4YfBVydTJX9X6J2zQtmX0a
ix81RI03Ne2xthRVNnikPWiX+2UVxBSP5lpDvglNmSf3oB74A4kejSeAoK/uKGGIEeDNjqh3q2QH
2n8o5TtoJN2GsyzZFqDHt7zp33MDL7IrojXWvOzq2MhptckledMty3QxjKPw5f6znNubLLTzgMCY
IzlEvsfAlQufQspSR9g6Bm+BNyxuVzQgDS838wwBDFSg38nFjnv+BjC9sZRVXoQqsgUthKjF3tyl
o6lKScGFpU9WfmYKMP0zWH1J82QBwaWELIkNMk4HzQi4t50unAJcDC3l7Bt/Y5IGqs7V+Wgcteo0
ETHvzcArM2LdjfGVRI637lP2YJS4wuB0yVFrZvMmvSCGx40W120r3S1Zlq3lRTNV/kWdvGOKP5OX
hB60zqut/vVPfonTAFm2rkEuM6jqaEbL5JNE7ul0r/8ah9NhIRhFBPKbAa1YRm3lz7js2Yw1fMUU
mhKgpVYwobmP5e1+fUfhYJs6dokNX/lEojfj5nJ+V5MXUCHP1hPr+npTqXo+PRyum3iilofRCxK7
tbnlCwljWt2k9TnLAyCKN/1407m6jTI1Vpzqg6y2aNoBVj8ED1H4T0uk1PTNrwbH+ajWb6IBMWqO
VckhEbBC1oiCX9ieOgX/co1G0H0qXMWVfKNSDBPBjN2GR92XU+aXH4/DtKMZ7RHps1oiTyh8l/IX
J95Iy9X1eX5iLwuW3s7/F/eLt2b89z9MvZZ1mlEaDxD4NjGYYko/KiY+ZJiA/h5haAft9RLuj0tS
nu44NjyqIPXnZffxK5X0tctnRI047f/Nba/rWt0DIIclgUuvtGdzSah8R11PL1gQRt1np/XW2kVW
THbauCSSSjAYbGzb39nfEjwyDtJ1aHPeA1p1OtdCWlGSH15g5ToQ9HDuef8N4HJEKfqTkb8+pMsC
hPygOvwOTUHcrugzlP8k2UTtWgMUPZ6AkHzrOJ/ZlIvsRnO7TQFJlwFcBVQ1JYcAczP3HOwWDVi+
9U9mO1L7vD+kzntf24mjfKTiRzQHjXHNRec1y+nuMvrdCj85XMGa0wHb2YlUqn4V9OHOq7DYIP2/
O1r68hfbYIgsApXcGbeC+Q8ujDeGuRPGlb0rtBdiRPnx8zYNSE1iPKw1MKUxu9WepfYfwRuKw1f3
ihHvPUYWTDcH/dhD6Z/Ck7HPsF7r6ULZG1QQndNZ4X3vw8Wrte+8UtnNn5M+K+lVl8777pSLc+CY
Rm51Xzg6EJeYv4Ew518FZt692zijcAAOmGNZqxhv+M3GQV5afgLMN7q9sq8TcaDEbUDbFWCTp3xv
Ix1DYuawBtaii2Fg2WKAsCE61qeXzbjBRk3LaYiYCQA2FTmqi4J/TvZPPhZ1gX7JgwPpf46Cb9O3
DfDcY3gCRB4ulyUE8LT/FWOOKmusCpjoMhJBe2Gij5LbUwg9KatWg9f9dvB0x+3i52BlZ88hZe1F
z7BMQL9Sty0KljaE9CVpcgfW0dnXj+wVAYrlL0Gn6JE9J5JV7DmeF5zEqBaF9Pp9goYuGf2gY36R
R0Yu1acQfUuPHq0jFUTgZITH4TjcZQKOlhTtjzI8cAMVTkjXWGhJnPioh8Rwt+pUj0MEDOAj4zza
mocAldJHyVcPXqkFVYeSVXMlb259HfkvxZKVTPdG/KDypL+o0qVZaG+vVpYBg0ORY0VzpcG0MhAd
VXLUf9QVWBR03P5FHmqyXRwXo3IwFDB3JQa8ZdiyEb2ipwGt9le5VTtnrzSo9cQ4M/lIMkBF0WuW
ahqXgdhNaE68hPfNvUGa9UHbNjCirW9CQbbsEu1kQOuINaJmkN8e1nuqxGl/ZOPFRNYWM//Hv6zu
RuM7YTSHK+cRrH/lpJgsLdzfn47F21rvZKf+HeFPBG9k0cKa/0HuqQlIy0RJHAt/G72Fxj4uEhyY
oENhLo/Slz64sN5Ps8fgiRdtwh7cbC0kILQExjqE/CHqbo6/hWOrb00Kj6ZnvdfrRqdonoZbIuEo
Lh+9syv0EyzcfXsWcHGY6M0Ev6B5GLaPIDCYk2CNLwt6vTrh03CHaaAkKT1SR6TFb9Rq/ApZKnoi
ivxMV5AZBRYhh0N19CBwVnzNdg8rZ03PdXQfURRwhO6H7deGv0Foppzo325A5L8KluAGon+eb/nC
kSzZS+nTLLrnEdXejrHREqsN5jAaFXMOeVXXMpabnPO3ISbliKFS5iWGgGb22DhMClZvnQ2j2xVv
fIlPQmkKrpV0uyaK+0Ehvgo+f9pgGkYTQTC8hfQlkSZYMZp5F3M81eFChnbjtJfZ8Arcw9/AVPoa
V38J+wUNht/gOiBgcWiJpTv2+c/6p4Ybd8YLACgaP9yo388s/2YylC4bks1/ZP3dpVnqr/6zt9hv
a29vbqs5FJIYa/V0zzm8P1Ftheph9dzK81J8UttaqNOHDPY3uIDNx8zWL4NwmhD3snjMXRzZW0Si
Bqapa15W/+itM6Y7cquxmRoA3Xyr34qt99r5DhtlsaNrIgcE1+6yLnnz59wcL5gu+i4GU82OHZtE
p0wXVqNth0h5Q30QXpuQm2y8JBv4HMNuNCK4klkwrnwRxf+79yVn4mJrm/WFsR8Q275HDEU6wwsN
3W6PsA1LU5CKKJqLwY9y7pZg8oDS3BPh8BJIjJ1dZP4ZQsxZ98TjILH2AVyt5xncD7K4Rom8VnE6
hbm6j3/cSUeDvxZaF064rP+7rctAPe2GSVLeeMHrkmQSRywVAPdZXZ+LG+mHPt/6DrQluMU1T5XC
8Eog/qaGZ+vitVdNWdJ/oenvsyjSySamc8xQo7zn/4NTK+sPUSADptCrzF8JEkEKARK19WTuGmNp
PR1iFQ/YehF2jF3rP9ojHlkUG3yjFENAPTw49dUJW+hpnX83EaHKefEmampoFcayvTj0EPRlPdB9
xwCi2zqBCdSQmo2MbJakMCgJiHQCtdWojHWTIh4MIWqDZ4wR5AM9lUMYeGxTx2ECyJzlOrIJILFg
C727hy/WjOeTJJiH5hjnujZgp5qUaDRrsqx0TgAjP+hbVehMltxkt2QouronAAIY84NThWbKdUo7
cssvOvOco+Zm7HYdnHRgb4xD+5Qk01V2V79R4gm/iX1hnrDCbzsnDG9xcKqCWm9FXoFUFIdaobhA
5Lh5HT9LSPm4YNnpVZ9awksB+D7YNLoPeQWNIaO+jTckNXDo00ae02PggeC68dfNOW42k5PGqs80
/ZYtWY9+fncPlfMqhsz4uIL8R/kp5cWZ0e8Ot3MXef0gEXrb1NT9bW5amhhqy2OY77inywYd04Ji
3iAkTuGTEk8+VkJ2zmMMJ14G/HE3M3vpveLofVwSuVHKu8BLTWvVoYcCrjGKMpd2lGr20Vlq4X5c
8vxevfUUkO4gvgT78IYi2sKqDySLtyg2KyW0k0ieZfJKlcycc4TQy0m2Xuk0PBtwlVjRZNuKksTQ
YdV27vREv3LVt3iiKrAZoiAABu41JFYi7QtNpgFo68A8JxRNfTAYpnzdfOw11arMshLaMScViEGX
SFLMBYFsSg8nxIawjKfuCOyDumJPobFK3+ix55Q14+eawD6TKehGogPHz7N6AO26GjE0KoYD+TN4
CCzqbhSuPtJVS4LMIGfP5SjIMTP22dm2E9yy7C8AT8o3togRZHwXagPYeRrLb0IUyG3tX6awGINo
B9Xf4GtN15XhsA3pXkWvfzPOXE8oHZ7DuBKtOdojpg/oIBVNmUgfVmg4IiYqm0UsiVByqhI6RYrs
gFWUQDePmdOW7ekEuoUlKE1+2RGCoLvRth6rnOhiGaX7aEPIGITSg3vcVCa342gO1ky8i5Us0i3Y
r6ipjwfEa5q5L56XpYFY3c4fQV8+yrfw9Clx+xg1RfMfhMtjQdg5XTk4r3o95+JQApLi9N1Br6Ut
bo2lC8WWaW4ckNJrSI6kPTs2c4EtW/tQLyKDkYUUcXnNjEAa8ptnDAXDzKvjVhkEUoXyGCPKbpYQ
kVxepnmCxh6Lio1GYH2tluyju+LCXf+2X+RyKSgsqh+kNiDsh/DFjRvc5d67eQR4tm6qy95LezeV
pUdfHkPmj35oQ4QcTtn/RZ7suD3ykKj2SY6ToHHn8EWgfAMmonum8nrDPjp9rt7FJDqo3r2kJaW5
LAGA1KmbcPEeq6tNo3e+JnjE1uXdxVK9YTP+xQjyalEsIuxq0yVc8qDoyexuM26o8Bg1VTP4efjN
f0WISP1yHZ3Ilm3CcY4W3+2HjZYZau0mWhC3PDE8mJX/At8gJ6cYzGak8lIDVJspzUJU8CH0X5WU
XByjzlI4yDxBSr6u4kOzrF/LA/heovKX6EQkF/sH+DEpvKxVxmQvd+2iWDQPx0Y5QYqClr362jEJ
+oA+LDBphfXSeZpOA4sKKVcydrt+uVHzFp96Rr5Xd6Yj6U8m+pO2QRFg1JHl7c268qZ6epjfxZKu
ojRK2lOA0WH576y6nv9Cu6tFxwg00BRi9bWsP5fiy76+qauch4weINFyMaAbk+V9boXbxjSAVAKj
hq7EPbJzTC0yaHTXCQdf8hTwkmjCqeVoAugJLiFVgs/otVahXH0uiSOA16jyYBxdxXLu3VgD0P3t
lMAOPwgDCvNIxJA3D/HU74PtvHBa3xIGl8wxUMn9wrVQoYsuNsdyG7gxZmIrTcoVPw8mdJOj1vmB
Xm/Lgb8f9iJCZSjBOjqvxr4AZ5FhVnaCZqLcOJa76o2hwljHG67OstJLpvyLjCWGsDWwe7Sx/Uzx
6kLwnBKQTbFu5+XxCJHGE9PjUvhIbJbg4yaRjUBQmY0OneUi7k/EfFGt8nhDhNdReCXP0jwnYf/H
mqmyMkGs/mBk/oJIh+4x9C0MCnuqs1SadGqy6FQeD93W5B4WBWssNy9sp6XSMZvp+WkmlYwbfNDC
XIFyRpm2+8ZE77fVwGBdCv7lRuV1WaCSk+ONUwas6kkyqkhtPNegQpN1FFLHm9P6BHmmMJbJIPxa
R/HEpABlogCnrWxqtRW0Hv3rh9mcM7407aKIRFtUmKC9zH8S5dnaUlNLDqfMTL5DGcqp1uw5yME7
ZoxxyjaYhMBMzMIGsBCyzHd7WYApDM1taFvGlHXazFRd10161j9kDQuDFUKuwIXvMU6cOfLpsT7+
5vw3gqQguIBpb1JyXd4T1mnZGv83Dne7zpPiDLnOKlfU+xBK4FpV6iosaD0n30z3vT9as32jg9VR
9maUmahXQ3zGBhe+bD9OnjmijeoCNBRxjhAjVsLnyzkdePT2hvTTS8vzAjYHzFs91U+jOW7C94JD
RMlkAL8IQ5mvzhoK1CCMXgbFPcGC23i5J3DwI8dHrh3LINLoY9DCtXKDXrruLhHHZ5crPAAegyMt
lCJVdM5YQAGZeDSpYsIg0qLXe44M1WV8NlJ17LBc2m0CCkgxBcEhmJX5DfZ6hrMOtkYH1KBm7fcI
OyDffCzX0XRncXcN+WCJlVHioZdVMg4N1LBNPuzBET6uSkAJmcr1qNRq9mtxMlJOpJmmYnaPEGgT
T0K+6puml2fJIrA7UKg8mLbbpjl3yahxU3wO8nZSHG2ygEGPVRg9bP8cFoMJEaaAVfDBWXADscEH
6w8/mHsSejp0G6NrsfA3T7QlKA/B9fUDRcu0tkCGvMiPkbICda0VueeRvUEi3JDIfeT9j+czwSxC
7RgPjDLKcXbgzKs32zi/dI+futspOD8jbJQ3x/QUS2uH/1UxgTchMp5zj9YmGPF2WdKClDsOXBGb
iGkHlk++3OP+jpTfejtsBM1tDi8x2Xac/Qv1AVslPh4fxSYdwQakIFLA+z1/HRgViGXiJ9bPSOAw
HjLTD1crcxCuK4UHIMVbKjwEW7/plsGoh+NI+R2fP3coFIH1j/OpIjsG05Py5W8E2b6MqnO1Jyc+
s7/PlSogpihYIqa4ZU5A2wfCnIvTF8tvyM9MyVoy1TmJQIZSOfIhycnzpd0hF+xCPBSZgLJ83HLf
BPsJE1uQgdpBHpXkPGx1rnDpA7vGpNr5vI+CbJn872mqqrs4tKuWlOW54mbHDo1eorYIe5AXlNTP
YmlvfTXWRe9V1h+VIhQO1DdpYUrmFXr1e68cFDNzUFyGW2sPWgBvE3Mh04chutW0cgDeefzGnXJV
0juGriJEYUF4NFLg5D874+NpTrhmHnA7UukgObKq9gWCsxHWEQUlsfXB7Yb49GK07ZKRxvY3YQtq
8HSZyndcCH2r2oLO5XP/K2StAJv4xsMLRfAkLwdYpjsplVFfmrSdsNg+vtaivP5OaN2JtvjysI1c
B5Sm6o17xTZevyrA4m7KnzxGVuxt/Jnt/wbVF69LiKAWDeFQAiV1hM09LMUIZZfiYCaXQtwg9lhN
JzobbJ1EGNaaLoxiVkmuVH3pXw2JDyXClLnCzlBZ+rOLo65haJIspm35468LDNEWKQUxui9RMdB1
WaWEmMHwr7z2Cjujnvy1OKT09fK5pmL3kl4gb/hONaINeimh0cHGZI+86mBebjCe/00Ohs0FPCFW
8yvR/DNnudkW0rTtdi5wghp0tFHWxdyW5OJepFbzrgX1IacwVbK5O+NxQWNQs/ozNSBSNaQSUBd1
+FMEXx/OXTNltB02P67zSnV25R/wGThg4CGDUPBdTJedD/d9Cu3czm1SDbA2wQiAS7H+45IyzdoY
qvx+Zx14aR0tdx6AyymAt4lc+cl3Rg2G3FnBERCymWTNXpNBRyE2z/G65yBEZNKrFHLq2TZhOnzc
YUWWLe6rvJCPXrhKuFQf/03xhen2WxwT3dBSPFIKc3FfcI74JpWWtkX3PLXYCWJVQwdT7BwEg5IZ
TikSpOiK/SwrGrnUN3NdJuTG170psRFt3Rm4DY8Y/yuUdAf+fN/sFo3v3Nipp6DAQQl6lkPuRSI1
toWeJ5nFMPpzP78oowXUXDCY3Zi36JXdmYyxAq//t1R8jhDiv95D2y5rJfbZ+wRLmu03gGdESrWS
ciEVATnX3vukoGS0M96Xn7aMa8rEmRUK9QgFizgARFsA3BBeeNpALsmvQKNQydA6iwDjAQOnwYfJ
zDMG+bdBLcmPa2AbH6m7zZNNVe03IF+fJpl0cCxDArjj8UUIPLtXEKH/lgUVe4IlF8362ZhnjMn7
ApxVKOpHAzXql2mYia+1xU7Y4H+xmn0KjOUGH1OGSNACC5N7u6QOoJkyCiJzMoCXDoACCWLkOdny
+X1ESCmGc8c9XdI9eApFNxEzDl4ec57P32pqta6y/fA4po04ROKh9dMj4+f5jYtgoopHAF3NBlO+
OvryiMCjAuUhR/cNVYnxR1VpF1bz0R+6WInu3MjeWFNceZhuTiR3QgSIxsM71BPwwbTrbHiw09FR
/BO2ipoSQN35bYp3+tfgK1voiiqHeKx8NXhjBb2n5v2p//+zSzANnxUbgtq864e0srfJL1Tg5wbr
fXo+TX3Fxn1Um5xmvlKpOIj/iuBycYxRnOgVe71tsoPlfraRC3y5PVkcRIrmfSKpTY7+MPVbjuDq
jD/6lbIcWTus9cWlPkYYvgVAQ2offbKCZ1D9Zmlki3srrMjiWvFlz6lfXxoznYSC1LjCTKbSHYPi
MOtq5L6ZOp5BbrJdDdR3+BOWBvCFKomCG0NPXHZkOPiIyugDJKD+Hgs1OuVhvWC4TpmhCs/mq7z1
VEX69vP0Y4F87VUGmQJYIh08lyBIxG/LMvC68BGKfIG15ZL0FFRqELnhfEuLtIFArlQWZzh0MX+e
DGf3GYrQAoLro59U26FBKurfUxcQw3nyr7SyR9lieJEq8PvWJCwf8x62XN4xRqFPr5Oyx9ed7qrS
depKl6lyAmd0Gwv1eeE8oJi//9pF7ecTVoHSU7gauG90zYNt0gpaFyiSE41ijOcRFHjtZbfBDSQk
RyIsmSza97JkVa/hPZSpMu3jypgoOlUM4M1go6kJzwSDSoIGhkmT5JR3i0YlgjDIjvawpLAPf3Vv
GLxg0BqM/QZOgywHHgK7qEeH4o0N6npHxAa/DKg3fQBwNLI1zf3vet8PTBmKczaoxMBft53EcaBs
UsDQyAMMFIfXgxhEAjn1df5/n9t1VhulWW/VFhTWaX2pP+WvXDGWjI+SvndawWwtNGpoHJ1BDweC
EMAhJX5zx4wgIJzDM8Zl+H3rsrMlRMjICFc6fPpESo9LTTqE92mh72VRJSQwTJ0P+6kNt7lrRrdX
6pSNnGmHHI0M+o6k2uhNp/TA7X5OT4alJQLwi9/a65kWo6NJJZ3MIF5g8b1r8kGHelWGzozsRZ9/
MV+LyTyd+cq+vAfsSFOS5IBOQ3jD+JExPW2PUjtqQ3TKMqUqd2vqKwdJyWlFbIm+Z9PwoA+mb4Bq
bHL752UhOhBtpxlVlhPWTqnDIxR78GP+taRX8lueR6BjYgWkY5eVEk26yltMA26g068vD9E+75hU
t8SNrcx/nCFhw8jcefxIg71IECM+9lB7mUjVRLRnqEZzQolAixnr3h4XADEyQ88NXGqrPFlCYpYN
/INY1ufSSVWpgfmoJmyXqxeNblmq9aQI9u8YZlb5LNY+UkfMjIsURaro8F2a1LPycUnxyn/XHYET
mqrAlPxUKkyknlhmF+dB9vkE9+eDYMkRi02hT8+WPocAV2BIGEm4wSbJjvPwnuF5Po8eLJ1piwiC
seUgeVfxL6kK9j+TJtO5guisIDgXv79uSycQzso8NzsOWwBjR62UhC6BiOHhEmkdYLRvEBCPSkv0
j9ekQcZ2zvbPmFRNRa4WRpnCIn0jJ5//pNN77NUtA/A+gIxnHHw53OLTGEhH4bAqpcNZk5CZXrE/
UaI1wKQpqJqKdQVFczKOfDa80+YBuj4OUZbyxc8qiGdcRl4xQFEmWw4hJdQopTQZ3OzxyPgLGwfG
4Wklf535mbjacSU1PAkK2GkArxBQRC+iDz08kbl8PQHpsfx/GcwV/tHSEF4Qc3ZkOQYb5LkWC5nO
aS6fVHATF0RCvXdMjKv0urUPXK3arnchnabffE7FwkrE8oNVWhwzbtbbzf65Bb8/w55QuxluIFXQ
C77DAQ0FMTpKT6D2SJ7cxTNUuVpeUJpSadTlVppvfMe2IN2vI/0S4eGMqG/WE7+dFzyZSo7kFBF2
aoCDOKrsyKc+VHlLYDbhfhXYDP4YQJhOHw1mxdMVTDS6s/6A/etQ7xZd0VRhZhcnheX6UY4DF021
p8k7hjRz+3g6fHmJoWRdjFqRt6Lj8CxM0dQZTwcmt0SuI90SaKJ5fz5xkG1PYwjkYqQ4RrGqQujC
YPCqXPwRgUhJ+sLCbxlscqD6rYaReIm7ViFZ/bNzIH5Zw9smL8DRlaUuRK6ubm3pz6xlcwt3N7My
1EDIxUlNdaJoZFWZFuMun7KDnXW9dUQblu8HVp37TLo1CyPuBIgWE5monnZ6PcPM6P3waABpnE5r
dgOn13kZS4PekTUxqkg6be/MoxICD2tfJFYFvWuU+8OUM4ixT7PQfmZ0MA2M8IXuUYd9GgbxPqAh
PRbPyyHZ3Hzi7ThVmzX8rBL+j4wFC+TAy0paoWbxiMN9MljO3zvXK6a3HiJWUIKT8+D/BfGgiFjA
oul9RAnQyFfq0rJ6ofiYjUrDWHOip7BNW3A5Thsb9pHlAfdn3/Xqiibc1q9/IcQVQ6TiyNkNd+6U
8LP1ZBB3M5GDDAPvxds4qR5VmBRSZsZTmaDbn7G/CcbkY+YVEkj4JgbHrGYfaP5u7MxKeNtJkO4b
iMxBfYJdyNYeSSAnMTDjNZ7gvOQGa+0d1xQ4MI7LUtF2jFXrFhvcd/VtFN05ZFlGkRdr+ShO72/H
XLgphAnONPSjHUizQWgir6eo2ylOYs1bzu1JG/W4B9goOKoQZRDvSKuWCSHgcx9NUrr13uT+tQ+s
jTPH2dD+wkGm4uaoUsacWOT8C3M7LnvuxGDBxYl5YmeCoNHKZZMmvfOyJwYw+HJTxEfSMhJKdy5x
57yfbaOXZSSVDjDqxcD5Jpt7HvPpX1HbalHNTJp9JIoGPfaBOUzyMi0XotLufScUKzWDlfpzFHPP
gN1qFkAfIadVH3Hc5AgIajpKMc3c3JSKXv2NMHTr1XCpXAZ4q8W3E1cobkbJJcIPdkXtN3KU1GDI
qTJDQpjT9+ZYswHkAZ8aKyjrlqAJEfVXnQVSHCTWXKNrhVxRsGkomtizKFbSE4bsWAVKHPspyn5G
GxzMJfn5C2BMeaLdk2rnrGLQdh8Y3TTp01ri8xG0Bgio4oyOitkPAEKRqXKxt4Ch7uBIz1dz0nlL
3fTggzf5pB/kfxB//S+PZH0RUwwtTbwKdnUdsrnZoXl3YJjcKmif6gTq6lO0B0n061IqWKTAjtEz
oDtQTF8tJcLPthVx9M+EGANhijiLlAOvMfiRQ530y+b3oFcmLFgvkTvWS+LcNvyMva8Gf+uWoX9k
E9mh9IdiiNndkSKprOKuDv00Utzlz7Wh1pRqR8tEZ8eAkNgKV31xs0EjTR1ZwjixTAcjbUQOuloE
MKL7OSzR+DSVdkGi5I47N3v6jWoLhzSLvEAn93HUcjXI3UmQRfv3mgP3vo5MOPVhbU2oHhrTwz3q
b7Jf7A8tpWz6w8c8FIomx/YEwm3+F52YiK/nBpRDVgNFYZDjHrEj2nW4YNghqjbqNJXtDwfupb3r
fNIpD7VgI4TsvNSzgNGq+J9p42RV9vWXoWUg45r622/yTQsmqhH5ac8CsdgBGDx2EKZzfO59JmdX
9Q4lTbAdR22FURlazWNiPVqm5nkzeMq58WEu5j/Gc5KawFdMg9J9mQctUrs6nQZdgEthWP/4PymX
Z5cyWPAsnq8bcmYrfeAvQu2Ok8L5nvYR1UuDednVwpovRbF4iHDhp0xjlS/epXvps0kHCJO52p1B
7S81F6PVocZSsnTLauc0jHkFnDYvjL0dmjfgztbf1qCtrfRMAyy6KS6Xomg/N8BvQJ1W+T82tL6F
u7ylLSxDKRZjP7pv1wrOtxSYjibcUhvJgSZ1SoJfbwtEzZ9aP8hp7Bg/Vb5+NDkGH9honazBgONp
bzXILoYkxAK0t3STJPFJgnj0lbmlumxgGkbuK+Qal+wk+9V6jA00+h+WF0/xMrIV2hEQzuQc06ts
jv8J5MVGqt0keiT/L1ZH0rBeLm6AEbO6Mu4mATRH9XdA8VpuGxQ/+jLKpWPDuKsT8C0BR73c+z+F
YOkGOqth7W04CEpk+nCvoRoiH4JpUOcNJ4EABClG/PVyXPFymuVaO7xVbsNl+R+2Jh0xq+w8BBcL
Y/foovZ96DnjiXLXSWmTLnUEu175DEaNW3SeOV7lbrRSsr24G26Fic0mF9wm4NJTLzg6NDCV0JNc
TuMhHbOND0l2uKvDcT50oWpbpKMlO0OqZTknCG5KJUPn+Y6ZORkoJEpX06QsYP5BNYzlILEhxsY2
Kf0mY3J0uyMRziwjQ3FWwMP5mLnbrkkmdLuADn/4KgncYNAFnKeONwoWQuaFmkLnYzO/pH7GghkW
Th1qmNsBgf9C7hSyPxAkGkkytUTPtOKI1xfCmckNK8TYsRV6//ECWEWYoyDfGbhHf0gLJRiMLj4h
ztICNiJCCgEA7famsKbOduwFLEQ9ML5HvJz0Uv7NGPtx+xr4f3H0cguSQnRLni8a57RAEUzcgbpL
tvtZB7FeZf9VPHTt6WJ3tNr7hEwz1J9WhLJK1tTMt1NFAJ+lX22IWQKkG+aA2qXbsnNfBZ3iaRx1
pJHd5SFEqeq0m6GlfrI2kCmgcZCXcIrmnA1HHlpfxHvJjxSPtRRo4wGpzGtNg0gFlg8fpqZhkbMs
VtT2Jm5z7iGGrXfWJqau9h+n9rjZ8qqxC8miL2NfGkzVveR0oeWfZqGeg2XEpF4IkFzC2LQzmhfh
w1wai4YHmKARwdnnzFUQQxg8yxbX5QmbWpcZiwQYPBaaFOC0oJ7s6UQb4Klaxaql38BwlUTS5e7C
KqrYcHQyMr/Iv1sN7px7UvyvGg85MQLOC+7V9kWV5ilAclDXXaFgFGfiqdlaJMmcocZlKihWr+9Z
wIxYQ2IkKOxjztlGAOD9yyxR0dezmBNHkkrYkceZ5PAqCl6fNYSeG0hPIIji+4RzLvxrvpl9o9Nb
QfE9IDMLH7YDQlhLsuau0U2aT3q7pNPCql4rHVkQTA7M494aiBCTr9Zr72w009U41Otwl6NI2MlG
UpKB9rrvT1cUzR6oy7I3I1F8GLy/REA5G4lW+tRVFEJn3FM+7fmlHtTpgltZlnEar/1IbiGVYOEU
fl2MT5N8vDtOaa4cnPdjrECJ7Xv/dpZCHfzuWpuH+4oNqq4yHFn+tFHxQH3lM6+LP0EvSdTO3pi6
sXsq4vjAk3zZ7WN9utlxoL+YMSL0hQ5eN4+zyO+bR/aw3RGQXA5U4Gk4NsXnCyAYFcI4XFYHn8Bc
Tv6cxC50HryNuIXxG9ayroz66By/Hzc9rU2Bp3GSesHwL3V1hEEzFO3W/JrgqTJqF0p3sZzzLp/1
VPmmuUoLf1wKX/dDhtdfOk6G1+b8DaZDbi8igDShjXyschgsUFqDfTaP2LWBv0KvK6Xjilclhgou
u8UU4SfGKBFZkvqJfgr3WXivOwro/XrW01jP6G0lxNnBOJ+rPBXnB5blUJmqAIRckMKeTbXYeo8z
jZ8JMIzVFD+FoiKhhxw4AkIECvQmoGWdXQEQ05TKMUYZxHEASewrVkifUezpZO8tVekWhdmQHWFT
FOh4rvZF/nli1w5/tlrAQ6BvZV0dtuJroBDc5YMdldo1F7q6UTJUXvYG2GuaByP4LXZqRBiRvluF
8t7F53oc8LfHGdlp0cpanGNJ2f+REVsKzsVBxuk3lwP+ETY4wtfa42fD14K9uCS4YnqgJrqFOSsj
n/qswfOCd+Nxa9t3RK1VutA7ssTohmtZGGs0tDqbyPk/fkPL3AKB3UKkypCjAzP6w7FdYWHQIC0F
xx4TJ/UuzHFlPaWp4aHQoW6eKMA5gT+rRCgL1oAsDxGco4VvjrRrmLfZvlU952S580zhZa12e+RK
WwNeEYQDVsATIbhzBPVXSd1SK++U5XviQaBmPO50Zq37fX8w5s026CDjGNqg5en9oyu/srDBZ/Xs
iwuR3e7UUzaeJcUr+LfvylR+8mEHVA4ZpizL9HxWQ9se1kOy/gSGKsF4CcYsRWvXNHUGRUfwWHF+
J6vlCJQIpWLXQ4z3BqJNRJ8rxN6vT35eKj1S1mEhxUCT/7u6zmBTmzDhePoXns7ZKZhH7vPWTxC8
9ff00BXN+8LexluEqxAQK+tiDOzUvy4LNYjMkyG5QYIrC5qgmrq7QpGTvlaUXMy8zvpoQ7MP6s81
ehoNRPp/yR7/it+1HGEom5Z6s3ehGYr4gauHdfcQ4Sl/eVp+fyYy/prtwUGAILnu2g7hICw/1Fqs
AP3kxRCcnTaq6f+AWhWoElpW3BIuRS1bH+lOvIzwgusDChkQD1V2QwaXvOsxRZS/LszGFID03+uz
G123Rw+6TQuCZBZihrN6vf6b4HhtH+sgeslGe3UTRKBLGb1H7laPyg6I6OoURBacRyX29fMrgUGg
YnUAnfHLEUOhqBw7Fma5WFHIiLBbV7TXWvDooCKPpUvH5nfaJdlcSdZmusftlMkxTsovam40+z2/
co190J4NF9o13CdSCt3wCrDq9AbmVy89QNOchnrxFNkwd47FJdoxz9ARdMZb+JY018Dlp88wRSmE
Qh1r437ityhPNyqNWyx2lfYJQpQwpPPLiZu/XYg+AeBtZXnK/zf6uUR3OPwkVFzGCjmgeS4lC98Y
AgKoQkUe/SGdnsQFH4pXsO+ZQ1skc894so7Bqc8QA7GQ9O+l5sM4EnQCVOA0HDWCDxba6AX08G/v
te7GoWl7wczJ9qWZGMrKkWevZv/LGYY+hhJJufOVDMHjwee6bld7FMuE5VlC9uOptSIazpwhkuMJ
aGxIAFDzFb1NuL2BrwQC4BhSe8NNlmtUb8/wGwBKhno5XuFK4bGjYVVW+flDMvWYFmS1n+NTTRzQ
TSz2Di0PTtg7YSoZ8Evqo1PJYi8SR6zn2xGt60s6MnVQs0YfaQOkzoet6l0/KbsSgmdDVEPATahK
SVhRdzSpic4QbzOhe5v7uoUeHmUvdU8dkMENoaK1D3bHyEH0RPsBRezzu+FQqIFSHcsLLMCDy4e/
Yt0sexp8CNvlCTss9ML71NVdkEOV1IpAGDSF9+BAEoJyaTdJjO+FjRplWUQf6rWdG4ftHcJXdo2c
vH1Yv2wDBTzZNDAY0p/TSm4QeNWYCKpA+eJJ1u26WFDus6nDaMZY03Y6iU4rvuoQ1FxQbZ/yvlzR
kHuVbpV3B+OvpZA5brJndToSmLc90A0sUuFyeXQ447rTEQ61wRvP8CWaFdrKj62xmOQKNkYJzOGV
FiXRMob9cuPtasjw34dQQYQy9hb/NCHAJREO4azNDFLbmyiQnhdp1IPX7ui654MQpMIobCSJtFgu
nukAe7jiMIMhxhWTrUUP4xdkrQRkynvsvzJslOy1Wujb8HmtSKzg7Aza6Cczh9G0ApcNVEo3Ltcw
bEX7VtDiOPq5gFhNEjcSUOE2UqVKAbgf/rXVIVfuE0IpwlFQy7Ok3EKEJE2SGZLYYjayZ8VdEVAh
xXKIbjx8wt10mKko8MCnzonb6e1nz7X1nABu9V/YGXKAAkkDjI0/Gn3wnhzRP0x0aTBvmSYS0CCD
lGgW/cbYOYVdOn3aCo9vYHYHAetMBfXFKJI1LCUu6xlYV6JHksFLfV9vKmis4e/btdDIMpQadbIk
JVu5gyOwSl18QEKV68asgFQJ0GpEmo7V2BM73RuCtJ67GknJgWkuuQ04suAJykQN1uXzEPShx17h
jgKC5IWLrFFiP/+KpJo7eFFXZKjesxMnn5+pxDS1nud04CsBquOAXyeiK2ApTu7wWH+63xEngue5
pkH3B+wy8dhnV1kUlyoAXkzsyWc+NpXy7N/WUBPv7Gbt+TAXArCuE6Tc085COO3bUqAVI73bvOpw
C5HVZ2XlGePmA4s3MaEDq54QekBRkEtmuwPspLuRLcIgecmwbOPknDPiLMTGHVwBgGJ+R1WWHdBS
Zxo5JCXyh//N6SS11c2TSSj60JYxiiUcI5tUMLMQRJ/Ue0ZQBeuabliljERzSMQ7Zlax8TcblYm3
gOnURKoOrXlR7hKFH5MSeXwUMiEtWeFpaLAILKeMp9QxQGEKr4FLOwzNHP4/axMbr2V2/MR24GYw
aQwpLveOBvqTDa5d+u3+BWsbZIUlN+Dt7CBQ5egAhPF5hzg3dq6b9I9cDWxI+GER1VLwvW+HzzSD
wSHaoYSgifzsVIuxsMHpVfdf1kFj5QiCi6TltWundIzWl1Ioh6uLUD6tqRvGiSOSQEfIKDx3dWIG
I15WijFnkeBuBTJMdLzoO0q2Es3oy/Ln4n7j/47PGqrqu7nbvFj67a4ghJ3k4FVBPJoPgu5ejCbD
LSdFHgSWEyC8BEPjHnkPXxxUU0fozFbZFLwGE9ojXmdH7RDdzcB+y+29R4V0RRlUT/hKAN7L5Rkk
C9YmAFGmoUmqoxhP8pPYh90aKCzeB8WLvYVJDeFX289n7t+LMK3FvKuqL3jWkXtvRwC6p6rQQBlt
arXC5m481cLoXktFRqSkSLTfI/40ZVToYzrkhEHQHm+xOvIqueb9HH1Yj0Eiu0507A+5aQHR2T0g
0lCjHCOBdn14c+DH59MHLlXe6CNRVnkcpW3M0pstkLpu3WXMwunh7DyfTYgfMIwW9kdJp+PTqw3t
G/7pqQ95jw7dX7TqsIb3zSt9qNDafftD45Rxz9/dMy5WCspb8AyZl31S9gV7GrgbnpPJraPbvHWJ
kJaA8bw5QlIW6LRSubp2Vw0X+jSAXvflmZx8aMcRXiMHI4yoZlrJ/EUcF7ee+i6mv9CKYn4SLxgX
Go34bPRcb3+y1bE1Y0x+BHg/o/iEiojjQXBlJNgpQ1t08Ri4eAEv4dgXfpMeNtcm7OPWDvAORDNN
WFrMkn3NC6YFe3NkIjsCSGu2gfRzRGw7CPMXs2Hm1fpRFQBkfhDfknktF1b+GVdmV2x4HcPh+29q
+U+TPDeB1crLF3HRP8TMbgEn40oYgnlir0ZT+0woDayf5WO2mdhiFB5pwXhQDWVzoj6I/ticnwbg
l4KrDOJrYHQm+SD/yUgGzST6oP4xDYk4WakfC37bQQ6pErwmd2bVjuk/KD5SHDYAYxjkBaHcJwxi
mjmh8gw2pDG2UNqdSiqQCmRVxayMzJHr01WLyBnOIjQdolPUG9DYrxP7Okcd0wb3D0IZcv1CEFe1
P26EF+ZrReAgMGDfXfyzz6L7mGpT4+xgmPAyLgoDzJ7/AlKevIiaMGWyCbk1EUMrbMwJGKePnE4o
NykLSA8+HHef55sn1qDmgJsHSpksK1Sc3kj8YyNtOXCaOiAw+/sPq7c4AjmKVoQ85V4Iy0rKDXLt
8cCtN7EJlLW5BmV0toy3tWRiFD68XuA1Iu6WTIX5s2H2MpWO4myVAtbDKDgrpfehtHcrbgCsK8lr
PZnUwcbNPseozaVqea4am8C5bHEcdJrJhsYfPdO1ZmN2Ko4ARSlSzQ5rg0+X9sMSCltpws2pRJa/
hDN73NTawKn2yx85UO7Gpqho1qtqxIILBnZYoCosLuTiTpiswS7uaGqqewKyNnytuv8M+3/zfv6R
LafywPjO0/UqtNquiXpOyaCVFgpzV4H1rnGLptxMR/oExn26vRHGPBC/nL4LTsFl97cYnvEtlNP3
CiMBGullM9gcrv2Y2YEiI1c89hPppE/137hZLgwgE3f41O4QhVg6qd3Ax4G90J0kbeMN8Mn22XAk
Kg0Y7q24/oxNfHJ63W5AbDg1kk2MIP9JamnaJ+iAn055fg1VCoyfLXqN5DEuZbBiL8OINX2YGR45
MN1bUiy/XvIH//sirei0gi8m/CZw5uWKAVwO6v1S4SQz21qOTSfoFFWahmWYW8Wk2PEEV20cSwwg
16x3EzJW+0Vm92DZe+Xbo0dcw/vMYJzlj4ywsRyu2071mIUzoyc0YWdc2KmjyMvVl88Ja7EUyn1p
oOm7oB8chtp8/cph8jQh2P++nUxBVBnITNiwckDmo80QsQ4IAYN5kEk6zDyIFE1J8pKXOJCrpRNh
+9iywtnh4F8KSA4UxEV2HHSQVUe9hzpGx2qdVnP+7/2tjVbfuikivzTEr0rIGNBL1yIfyzOuklfz
pHgN6Sbw5o1DMD6h1E340eHGTijB0T1fmp14jvCrMuXMcr9U7WmQZ9hyiy88G6ccbSr/7Yqj8reL
lX8snJIp5JEIYww859r2qqTlHJdibKjt/630MjOOo6lXzw0kcWO+UOcF5GLmKHrg7obt9N/ktD4q
zsIzQPQg9eg0QybNI3teeel9EQHtxTpKODhCQeJHsmr1qlDe53ILpk8IN68dfYafHW3YlOcP+vSD
ZhvXEgNLNZVXSg+8ZZPXeTwKaPiucL3RWIVKdg7fXO/PrXvBwpl7O9cpBJYfIyi3/KGE/C7uxbIi
mSZlGcK54ZKBHc6v13hfOqcLJ+ls+s1Ok73k0XyPg4nG3h8I/ARgoeOF2MgzQN8QLbG6VYg+i40E
J2UZIqrrRPdxUHnPAVrG13dPpiSuyTLvPMBzEEWpjzSAHkOahdaTmukOJ3ZHYOPshK+2BMaXO85w
MN4kYESqd2r/TORzazRPXq82QbymAJR7Xbvi1v1/mP9DUyjjG9IJFlFTMIm1iQBE9qJxlcb8Hloo
bneO8zY+YiTTXYjI+eVCeODN0lLzWCCqVG59oE+eM8BRrfuxhHAK8Tiy/I/aOY5hXSIzC4Jzc4mq
ZG92D8C/s2Zfzx+7WzTGu7afj4K9QpyLW+ZojK9ZIG1YbsfQXpyDTSsorjCpDKkUlf6t+S+kn5WH
i1fDePpPPeG8h0xltY2bOogdZIB1VqXVxgrayDfbXHk1XIRmoifpkSUMQkIO96+4vMgbqfB7ePTE
eJ6U1CdxJngnCYX68wSYQJs0E7DrZGPSEG8MUbLoJ+4CLbiMIsNvbIA98kYT3u33mMmI3MgHLapE
3mEezbgZcMxawXI/3ffGjTuIhdPgWyl0XxuRNp4jhzTFahNcx+6tl/SJAFmUNSXHM077GwpwIuEr
tvlzpSCtovzNvlmTE+GPzxV3FLzXvSgyjSm/DQXGOitfMslEf0PSBKpkIGbdJrNixoLgRwJWmysY
JH2qtVdtq3noOE2IXOMY/qqqWBRGmUgmznuqkLZGMumQyOKCSjFndaWvgEdTCo86D18cQfw9V2vU
XwsYNjwTDztQ7U8sexoNxqtUTlLeGrTiYky/3wiGfBTuMSzwy1uXxsjYGgRShR5dWgz7pcDOiAtS
7yEJxrnd8bc+1SLvGSPDVn+rWOIqH+BP5A3W+WSXDiTBaHGhOPQJH3tFu43bPsjtsoDETGaz+Rlo
k/uBPbm8jxC1+u89jvubumwncMqYuacfC1l/Wm4ZZ9Moxc3e7zO+v+BklYL1IvgJfwVQtVAquqfg
oZY6eVv++JXrLCl0xmDWow7O2iUcSHncBegRghx9E+Dt0vPC1RJiaEfaOasYpJDrUEvEa+R3cEEG
X7NYCHNce1Nb05ZeqXoT9hYLrqneJ5ktaHeR0jUlLQFFkL9iRyWw6KYj74LKSK/+/T9AmuEk7cHy
0SqIsY/ttbteowxWK/oEiIQ9wiEN1SfWyexMVRNyPM/Xc60IrTFh4WoU3mH0bpzHSAn5tn1RSmvf
x5WglL5dpQajGniVjvhs8fjuyqM+acXzcNe4VZHZ7IuBqFrctBUsLnQiokenBIEqP00KcHzfu6XC
6V11FP+NUVERYl+1zJUi2ffM9Kse7zAeJOEocmEm3OtCXLxMkzBaKqkMazeHkeKNixnqRaGQCMpt
rbLqlEeIQA4JTF/83lpCV4wYBOLlhdiLtlID2cjkAq6HqjgnNz83RuE5ybOihmEbsAVuB0wmeQfy
Nf4deWyf4lthW9G8j4r9T3fVjRnOwhfj2/yG0lO98MycH+wY7k+B1YKSolUtR2MA+rquVYuJhwEf
T/Wa29/xpsWfC7qWIWncZUMzhxTns+J2XaaQJc5hOrcXGDIfgiaHFookhGXNn563GY++zJwWeY/7
0TGph1PKZT2epV5GmPwdEvopifegJrGtbHIzyrcmbYHvMiLVoQJZYzUFYCC2zmn9lje4Pgs6TYzR
WrryrGMrdT42R2HWp4nj+rYOrXwlYJWO7RnqXx2D5Pce512Y+68oDB1QK4+0jiUstCuSw9TFDuCm
C2KplnAVe0C7vITsMTD1pr+5WbTqFDWL9UVVlcmULbD1pJR5DNZ907eVoHNj4hdbzB3JQ6rTddC7
z0Su3B4nJnW7QZU+tQC+AX0aLdBEWxzetsHLldc4kq5ikleA6q9AVAv8kZR+Hm6GUTCJ61NQZkqx
fu1qkWobjZYv9+Dn439+yIx6VQJdbBPKLq4SPxkqmBMLay4qNsXmba+aJQPdQsiKZ3enWtRAA8ZJ
Vv6sAGmf1goYwicLjQjStV8JKEmMVfzgUUmjcrdemxpExizXa8qHs9+rBu+DxMiJeVb4OJkW065X
VeT+5W7Y8KU8sxXGM4DQrf6/w13BUN1/AJzDt9i/nYexYh7RpnBtHvyRLTurkK15wB1bmdDf2tx5
8BwT3swWXJuxt9DclqPqTmHB5g4NXQI8y8y/RtP0geSJBU+l/IS5tgNGauCM+iqWNNn9Wo07KMd5
tuXZ0k15hm/yvHhPjq3yHiML8RPbNtKI+AaFV8iw7TlzEVbdbMn3xkfrA7ih5l/LAXh+ggVUg51D
W4qzJkiJmYoxDy1TyvSbjlU5vlhCo5fAh3vN8CNqGuITOLVEXCzwddZ/5XGqHXesRD9li+xZ1yng
m4iO1CTRLVV8n18ZL1hoVIYdYA/E9OhntiKPZs+i0dm6/tmFOR2kCHeSdxjGlCcC4ivqDZL2xnrP
eR/+QzfFdKgSQGdx66oszgN7DSWuV0y9GEbfAtGGRXH+49Gcjp/NHhSFPtAwTTzYGefhWKtXpw22
qXHJpb8HyOrZet88wIJ+/bsbMRXT0m9EbgQ3sVju7++FfYVHYDC1Tgbs84a2rzfPmCPmcuzgMwUd
AHG0vO7ZkRvGSeTgOQqdJlIDDkYq/1dwafocEiQJNHR32jcBiA11us02jHo+Bw5KPGNUAuBW+WEP
CjwjxtNYUM2NU3Hlr74Ksv8B+/F35BG1lMgoAdxFSWVOKEo0QRLWIBhWFnSXDxcBl5ZWeU6C7dfj
lNio8CTeTVEkmkDsvHPF4NpJ4+tUv7IEiDBgoS2LyRXq33W2Xbfe48qU3AyC6L44Qmhu/GDgpHrf
5wawy0coYSHQNFbCW/WfJ1qzQT1pe7GI1uWy05qjF0je+yoRuH2Nc3trnQs+vBdQGD2I0WKis3yn
GmanqOsan0zWYhv2bXrbIv1cg1jeCFbY3bDMfg9/Ef3kpxAOQt+3kWvVO7DGTXG1MagA9LnYJd7Q
PfnKxwNmJkONxxf0zQu+kjt63/qr2Glz/qDvmviEekOF50Ke7WEl+STOndirb/yXFsT40jTo2mTZ
usYmakoZu8PjZQgAd+nyCWBVGgDZ5s+7O1JfQKuNUmLJzNEeC60n6Mq9vzV7VOjmjXWfT14SEqu+
q+bq56O8BVrBMCatkCVKYvL7/Xg/3s8Ly+nvtO7mye3cWO0SQBSr4NCjT16FMhv70Tur+OWmQ4EX
iV2ZH3EB7GsTqt4fuv6VSPS0dyVd/dyFDYpsATcZFEwDUcqAheFElUTheQllEyNpERnCrMWZ4XP5
KRZpcpx0Jz6gT0uryHBH0WpLCdTlFmQwJ0g/Ulr0rQ1gbEUeUagV6ehygQ0EZIzyZ47KoKy6PFEg
CRjgM63xY7N87xJSLdAjQcRpoU+R2TqrJ8TFf9WfbH3nK1VH/nYdmEctvBuvYDmfLXcgJeJnVOtI
97PzyGoteq7hnZlLg8Q6uWzhkBbdU3iVFD6ILNRvHlPlUIGHrKjwU3qVzl+oTX3DawLOyYsW3GVh
NMaQGNIAVbtGXR+i5UlgN1vsqev41vcbPA9ywuonlYkOP2YPNtfmfqWyLbKDqJprHTXhWgJp7+eE
aOrj0mhegcanDzsSyORZnJiT+Honx11PwVk+CZ/bY/1DsGdyo+rWI/VgXvxgOszf9d9yjX5ReNT3
jaCJRCh+CQI4bYHBSFqrmaQpI6pofLrnRQ5RSQzxdKGQfZXWKgcZhlfPzE2GpEPQzngxZsqRySAy
AbXYKaJZ4CrMg0TMmt8KQOwjaWBphdgH5v4aTuHsIJIdEmfN/7dNZ/pjqteGwCnC+Viyq4aVKOH5
c3F7wHXR6ijpwdxa4MkMD1FT2lVMNTZQtO9RZyUL5E+76kd9Bpfm/+lEpPOeNBOTrQUpRUUkbsYs
jBV2CLY5hlJEX9ki+RxhJtpCIqocNghown+85BqtOFIgQqDyzJOwOYxbmn7r4PPPR4suWGtpZPvY
29VfmLlbn2IXxgJsxeRxGK2CJqityn4wCUaMZNx7kLg1qF8JqA3ep2ReNnwDU/0XHVXXyOStAtaC
wzONfwFmngbFyHQFe7TwxORQzGiv+TXQlcVCPyF2w5NECh62FCS01BnJ8zVHBrsO4wBx9PNrleo2
FAv8tcFHMu2I6lUUJfloMyYbHMXRfWJX8QKSv1+EMBHRLi9gd+1ANqP085LfDstRo2Lo3jhr9cl+
IAyqogApQqt0FYexZy6XiLRvAiRHTuF6uj/UXmUYCI3V7W6z2ouC7FKeNxc8YE0llvIMddeeT9UX
AWT5EEwlHH81QrxE0MFYPEvNdtm9faUgRibqKCEtbEVFacrKbFA/sZ3bLEj7nKUmbkXGsVQbplYv
OicfwCayysZt4YrHTXO+iSrsKYzakrud/OvVKoigs50dmbyrdYzj9nkh1x1r9WfAkZ24uexYUzgd
tVJFMpr8JTcbprCRe3fu8OxqxKpSpif/g278Vfoq2jyfm7aOr7zcKtTtxuedAB3bhxhPoxFgcTjZ
CDPx/NqySJURdkWP9UagX5cmI53/+GwC6jv/xdHnApN/hH+bb22AYQYUPrpFegomnXe8apGQRR5c
n2MMc8EeQCL4yUxINQ7oWviSTK9zaquDQ0sn+3hExRniq+mVabYGSaPEVbGQwpbVKze/Jnj+oI0y
L/Oid8T5696At7PX9W1c452MRefqL3frxu2XsSEsSHyeQqNnHAkpVBUyMCoMiqySqMXt3CmFHQ47
PePP8NUA6w3PoT4SHgpOq6iS59O6RiGlGni4613Tew20evXSMzLx/zomNPgxqdXBY5vDdrEXUsjs
7nbDdbbQoTO0I53o7sbjVjA5PZn/UZR3ymRz/C1QOcZcraZj+yMqjLKIuqIYfRk9s74KLXzzIhzn
Z3zdoGhoR/ziKXer3dwugbLJa7YY7BgD6eqsKW3mJprtwtfN8jTYD1iX9zxncF5sZZ5OW8VKGao5
BhgqKGMCNzPfF/lo2gkGs64/MSgyRP1VfvnNHG9KYuwPwtqDWiWs69xzmOFGs5mDl4ybyEHYsfSr
qQsfHmfQz/hjtFgepzJ+H5ysPvH+3FzXmAUtgHAft+E7NY6WKaVcRu1lL7zWLJ1cfZd7BOSnV9t8
zcPDK0XEzCc+JOZkIzgGPBH2e/bXkAnq7vYOm45pYBGgDoNzSHkFu163tTBqtFstUV4DPYEVK9GD
otmluVuk37QXZgDy0Q9Vpx4sF9pbCQ9ssusjN89UWGDfDd2AjgP6wCRWX6LjnOHxppcEPlTm3j0J
mASAHQHJk2k7Eafaig4h2JNtDsO2BX5ZcutnF1wjbMe/tqso03EnV0FobcVUrKXw2Xervrq9KWEb
CdR9QKrA+KbdTgScmmHR8FJTrisT8dLYjvxL7glUb6CvGE+DFu3vYrbgxt/MUIHRDrR+T4uW3tVq
5yCGc1DuIHnEgR14l28Gv5DqPyyKmeuMRg6c8n6/WEKV9i6hdmujunBCuKL2VS24w0yZmE6Z9Y7R
51qB3EaQZgbJQW03vnFuCP6Y04F+3sqVyJ0MxmAvonizBmn1U+X3mzzdMhHtG6Eqvwh/xr4+mlM2
j/LsmQxmPUObD8ovOJCw9QTZVMJ4kohWCAMaIFTQJTlBJUd5bUGgFc8N/s0BcLLPs+jI0RAZZoxV
sm9jp9qe4AMTow7mmS090NaGmLkXGvZYku2guKwahcVs+FPu0FbL8LZ18LAe0DRNzOT1TUGtvmLI
7WGNFiz6RxF4LH8TTjPd14jFcwqnMU1pg5s/WFboOE4FgpLL8naTMVsk8X5m0etIJ293lEcNRoFP
SeGKq7nkyW3noC3ydDmexdOqj5DY2le20CgrBEc8bsc6glrNw91quYervSwBaCndhhtGpJafV7yF
gaqnfoDvmKI2t/5W2cPl6Lle+Gyqc7x9lGnZG1z/u37uTFh46BAmzEj7xV77Cak9AvDQxERo64x2
eScKUpnIJ2GVgjVCOXYARwc6fR37E2rU/BshifNLRrkhoRTTxHCXXVsNFxoORDN53NUfwqcuCHxS
RHvSW/9W/zRvlp72MbZWxlpIbamDCjg1fuNFF417G6kE41KdD3pBRevGRgh+4TbC5yG85ucPCQOn
e3JQbUZnPqztYPYCQZ9q8q8UpWUjTr6rBAkxnEkomiBMRQ+jos9BQrzoezkwWdNAk8uM0WqqlEJj
KrIgYaSQxktlCYJVcwwAO3P6knfbYl2+wnUQk1OXqXczzgIeqjFjltSi65MVaSVhOqsF6UyN3vsA
YhCRmB6yGbx54BCCPcxeCuR4YNr+1vkj3JRSTw6TUVpzvSt8JCddAzheEWNZwG3hMu1Sb+pk3yeH
Yr9tMJsuUzzZ6iFk9b3VbVCJXNLm2sNXq/NPVtiWHb8n/TJMtoIdqRDPQYju5j45DQ0frDRsTrql
1PqJAnKCjC4iNWx3FTG8yKk68pT5YNrgNv4rNtfg9aT3e+kyApnpr3KmJ1CnspIm+JVS88udmDF3
kDvAxtQevrUZImqrNyPfw5y0zmK9c75iTYruStxXO1P6DhQl/o80PSG7QEmujL0xsOQN/ykbNHdz
cnzVw1JCCPi5WlzupNDbuPnQBTEiTB0Kl9u6EpjbxFoFCryBGjaUh/VGi5wtYaRlIbL5fc002+d4
IfRNbhdwSXI9HFCRYUBIJGgQZBJhsACK106yd7Y0FQdGx/AicVr8Rv8O/Bb6IOlw5+mFeejamhuA
69CbV8oX/M3LyLlfX2RizOXtKSWUuPyJrEhnNBQZZ+s2GYYkcMyOsIdnimyw76SPof+wzTiq0U1T
bjhrNeWqjUeLj3CfS4nNXBHZ3/ZQ7iylKWLis1i+sElCvB5r4dyhjps446aE52KaKkXH2u9rKmNl
VsYniOGdZK2dmrRkmLXjyTYNvAysIE3XCf61Un4xOG5treAselel2ubO7GPT0+Gn1EBjiN42Xzo+
0gGhJ08g7cEWinsmypKLqggCghUeVwV3baZLFWDr5tivbxVS43myc1WtYw3wnqwsI+mDFADUlFCh
AAiinQ0KR+U5GkkDL6CHNoRqlslEEaK4CMhK5b5BjDOhgQvPBXS+3aZZLZ3YIszYO7976WYN4tnR
YIhtR558VUSnwbh6zlwvtAIi9WYsTc5y26xVPwY5xcodHZApRr4D9WGZIy7A62Orq/17Q4RYxMYz
Ew+1YZWj9eiN/43M0MjsPJcWsHy+EQ50tMn7LWD8j2qyTQDwVySYpymk/o/YQumX3c5/lmLZDfMD
/xhGbqnoqZ6oErMjCvDC7UWRdsjuAXxQMUOoTUkRtDDCBdCKPtmTTj1WDc3/K0gNMUney6F2jpIR
iD4fhiapNu4DPnH9FDDSWWDWziKfrqYZKNhBzAlUBTD04cLueDWzgK6/oPq/SZDXbarcTn8M8iIh
0aJVdnMC0OVLEX4BRXxwacy+++s8wZV6+jzaiVB/2TXrcLRFcpLY76SRiPuCGRuCit2yoVD9FBq/
3ln6iTfq40BDyIuFruOHE2ZNYIsI6CmdBPTMhKnX9m2knY5HPXnWk9w2TLVDRqM/kgjVS1wwF4II
+4KPsEftGTVMLVEJyvSLnRZGvO6paoNrxnBcVNIYkFdm+3YStonANUdROV0F4bDh67rVObS6ooCz
Xm1w2SC+HvOY8EcSdlZMlTWYufD5fT5TSSXdBOPOeGggRsrdP2rYi9J6WoEplfIIHTd6T8XD3+Sv
AJxI2XsQ0dkLguh04wCGYu3dp7Ea8/YAjysadnC7Ff/2tZHWi6O6+2RB70uYPKAuNjrpZKmeOmpR
4udinquI5913r4Xoq2/+EWTQVQce+ehX9jhOXp8m+HiBOXM6+jNCTG0CxZ7do1ILiOBxnkC6GhQr
1bEMeJDDFa3f/f5CpT0ccu1ZvjKK0P51ptDydjsS/IPGZRa9YhyaBuTx7bC9Mt5OHtETkv1vata7
G5t8dR5DbSHaX+g9bnM98hnsLkhoVj/2o6R8GifSiVEGjkJjpZtTGUMpu7992RynF9e+MGeCrNdk
fhAPkU7xELhHq30q/gEKvetqX0tMr9BomHk+0CM9+FNAcXM21JolSkH3VKZpvqAw0VcswID0e0WR
ufbeSom8jjqJO8gx6K5+YxuL9HDMcTZM4tWiZSXovzh031m/9rbfQdlG07Bool+a5zGYbNA2o4pb
Md/YGE2/7c8rT0HI5IcO3fhKAkY+KqjqHcnOnDLtVnO9GNAqLdWuxwxjSBtCcWEyo+6RZuhpGVxs
qWm4jK4gZ3Kpr7hWHUTifuqj7YS5MFdwqlJeBkRDEvK2lQ7WY3Asro8KcFI28FCqUs+JKiUi64Yo
o3SE8uB0x83oCsD7lKexdU6drYS3JEQX4fWPh/nqwaQX1iwSZeunzcxz5PvhWzzV9bKwBbxquFXO
bfIk9VnxofBkJ3Jy0u89qFK3ujzBp6sTHRc5X+gEd7N36HYwLY7q+YEofneK0hHjIv33ff93Ftz5
KURrUOtHw3Yy/m9x6l+4/gG9xtuCjyrLl+SC97fgiSv+QUMJWKCoLCQWOpjURFTUdIz/1JfAfo3G
d7bkcfIt7jHxtRXmHyqJKPLmTZ2eiOB1AvdAQ3dcue4g26Nz+IIcCYeUYvB/r1rPlKXuQp9pspJ7
+jt01EMZYy483DgvrEdyTb4CPMQ5nl+DlopAH7b0btQNqyDwEhXT0Ezy24VZ+9x+o2sa2mlwsmNB
8jUWMEacQANT1CeDNwxCLsa90IiAEvxTJseahRyySVnfdeYag9w1j5fRUEJpB62XuxkgRRoXhLtF
UNBKycxxz9XWJ2MVvW5Fg8mJDW/AXuJJxMMFxvZt1mAqKW5XNDRqMDSNUZZ656HCOwWo/LdQA5yQ
mzRyfIRFAXj5X1V0EuhnacuJQDUAHaSownOFzQ5yRO9IouX48oF3N+pzYwHPIP0m495Oxlzjqwyu
+JsdBCsn7J8AzyXB2mCtOJtITUkGXUgLvZiSyvQZe+lLP3gxBub9OjCIOJVcLvgQIPIW8ekrCl9L
9Ta5QOKqJ0p2S4qmhLJ6WeD61FkWiU/6FVWW/ie4yuo2mdbk8yqJlm7tatR49QSZnD8hQuR1vzs0
53BlL1FTkSMdRhTrGKnX3OUJw/zsEiNlphRoQE38H/52MHeowsYV3R6LzK1zhxrFOEERmW6B5Ciq
/r2xm1rwf939HQUwGwdtCLcHN7GltthdP1J3SXgxkO5fxsERYAkhh/ZKlLAC5y+/uohfNKbLQV8v
pI2I9iIJwnbddb3U49qXnRV5gfSoZiGsnFMOUOhS4q8AOD8DZ1t8ZU7YUpnwlDDtE8Q1pVA+08Su
CM5WTrTjy5Zw2HCDfQu+eCo6mrOuyCH4wme749uT+LByHqBmrEwFHDuLDMWsW45kuKv7hiIPvWGk
HZjt37xcQlxG/CAHAzl7suJ+r9cFZD7a7dbc0dPhpv0LIM4mGA0u54u+zcSnzMPNsJxbJCV9qfJb
EoLZmOnacScQowaQwRhU1iMXe0ENKooABoI31xBASnTj8YIf6ut6QLT7SwNfKK4cCgmh6Az/XE2z
FkUsKEpLEfWL5L4A3pgyOr/GtO0oeqST4Zz5/CvzEn3f+mfPPkAGMo8U6cEmkcwWWNkWo7e1ZbFG
qPNZ4HgVl3287T1LKOZDBE3C+dKF7t0WdxloR1lgMsiWS4TPUDNpPIEgOpc5ULlybKQViOsOIW0m
8reLUJC9PiQ+a3jE3IvAH3blhnzFpncQDTcY2cQdqOkiYSdZD4acMBzZHQXjLIA5hKXvfziukNOk
9kdCiMcuKrL6PQH2UKhxu1KeUmI+IPwQAcNPUpZV8jb09SAkLXM2ToabOFA6BfX8ZUZSNxA+v6Xx
xP9alLrqJ+j1QqiASAL4XFdaI51bcuZtQiCxrsotpKjSsn/UWZ9/DKitlvLNyr9bmvl+EX0Cho1a
7LPdOGz4H0kurPlWJ1MJ8oFkdV+TwFsUMQlY/ySxE+eJA+dpPtaY0vFWd5d6GXhVilT3pf6qFXTF
mOjPN0MkGGRSiJuknc5+h0k8wYAVe3UTFHo1WGqwXFbrecMSsy3/5wf9+E7uQ1gXEnZ/cfxmjNd2
dP2t1doVQSdaQUkMDN5cnTJo2NVNEIb/JoOm9h/logeXxt84fPVyY5Un905enKJXhfcfSA4jLdLb
Dd+C46pMQ8kunzt11yAl9bHLECwWyR5JUpE8YXYJJ0Rhm4fFLssriY+BBRPdVIKgAZyknhx+UjS7
QuYU/eunzVqDX5nCs/RVreJSCX0wSfRmtOpf3MY9UQ/QtH5GJ4rtMxDiPAcQ/93ON4mrHG8DE/ty
tPkGNj5yC7R8Fi9uEL07qUbY0dfAJMtoq9xbC1ZbvaFC1s4zWCKRGv5CUEPPr8Zrw0yMjQKTQMIi
X+73ZGHJ9K9oVu9xehSt5K61WVDg9zJd764+BTaNLS7taRmEtxYQz59IzQt+ZvDZcSe/jbGIPS5s
Ce0LcXp53RoEmIPpz5r77dRej/oFanb1SE8ImPLqbJu6I43WQ2vYTwg7edGJKhDSpRUYh1LNi2Mh
DFv/UGbMD23uae0d372gOqGEVEfQWr7sA17uONzVKcnZch9V6LiOVbmLw8PpI+6fe8HLf90yHLhC
M/vVBrOKCoYps6Sdb3Jssy7IFLPhwi8+csfGEi0c+1J0H1uBx6ZL/MCyT5BIAP27kJ8jghgK3WoX
C0Wn1uS19zaeWK6gXX3+k71Us93yldjQnDsSN+Hm1k2K3xdc8Scet19rJq3bqZZ3fhAWAwGyw2f8
zMdBS7QcSYsAenJvr7dhjDgGSfHhH0PkAp5tB15eWHqDVlAbb0Eoad9OEAZ1oAP7HLzkNrjzthsf
3Lvqf3LXQnZcuRmg20C658odiqkeYZpGsWPpQlP1MxOR72Ff54hhJRrMsEtN5E07pbyU0UnFGxnE
KMxDoflimp1GJxSZcrwjRmw6KnNoAyYhQp1SmYtvMqUZ+qvI/ASy088WhKNdJ7CYZBeEc/j6tJdY
z6XotmZbk6Z6foIrTaMilD9DHje6tC4Y0dqaV/A1rj2OeqXe8+RMlwXOml+R1Jg0eWIpVey9GHNz
+4sVudx9Bh+J9GMM5qEoQ+oWl0yRt0Zkq0tkkLsYWCCjxWwFTaSti83ZrwZM6Cip9tIU1TDHhNbG
Ds284PmySLdSx3LUQFytOE34df8m7k3WLCtDhFgKjxXbGvcZxzD7dPTbBvKBxwql5Kfge6drk/x9
B3ZkpIGxyvN3EyOmI+VJXgZFOlliMKdIVslgZJWsTloA6KKNu7tht9CCj1EbcIWY1c1/wVYuBnh3
dWMuvt/clyiTRvoW1RCh4xfTY3F6fygEM8tW70aNAqMpDx503/BjJr2OGZ2HRDr+ZPcaPubU+Ibu
WkAi/b5vVZH724om4QxweH/XXFF94++/ic3t4hVfSnmzCREfOl9dLHS61og7+9fVG9zHIvm7N42V
7vsDuxBFiUtdZPgXxtCfB3IlVikC0yxHrmfOcMzPdpgKnLF0xSmv/7K7QPfH09L+4i8k91u1PAkr
DztqN7GCqgV83tCbQ5o6vlrPDcumQqzW62GDVgv82M6b8m8miVWwFw/DcCVpDRYpN1td5E8grKTa
DIgnmLBM8jIwr1OU9exUVSxMOGOg+CLJrGtJr5G6/4RBbmpjXZ6x1tzroi+0rtByLYSYbn1937/8
iJad4Dh26SMukUfD7IJ0bVepGDeqclRf1aPMLM2ScsY/8FSTq2Wqk9CSGNAVxagNF5t3PE16HSUP
vlr8I8SkPVqJJhc7Ji/9kJtx8izbUoN64APflBr8eWJyzCPKkxdCZh73SdVBVkaqiFarwS/wnsJ7
KPz2k3MOuWYFPuXiAiyZ1cWwihNNLMBRKEREI+Su8/rO0qNo0bYfpeWhGfe9WUeTg72rodKQgKlq
dnCwiBovhrB9GSzwjuI2rFwRF+jL4lxiyXRHrvAPne6Ki+PP7jXrI/I6UXtPc5t+nMuV7O5qlXRq
jTB1Xl+DrUpGQsqBye7ybepraKGjkp8usXYVNhN/FPWjN7HjlsWrP4JQFjnlsNcXWgd5yVasGDxa
sZ/KiOiqv0VddtrFdizitpfBPkJmcpV6RMBVK5h+TTrL3P58WJqKfHBrywGNBo9ifL9dlJ4ZyFiD
cbA3eiX+WXAGiDmrS4g1cWPRRmor7CUCzY8RAjIZ446lu/InKD+r646wC9dgRJUL5CZf4sy1DbVd
HZhE/gZfq6aQyHmXwHaAQE1YP95ui9oOQMUcidC7CAtgQxuGo915l/woatyh5rxqBFAFrqzlvR2s
7xDQbK1zX5nYcWSvRoFembw2e4tIn0/1pZ6OhRJmx7qdZBG0i3X3dzGjFD+q61G28y//tOa16Heh
EtT6MVqY/3yTPKzJOZ1MMcKal8+5+9oiQDk8w7yU2YEAOWSkUPjzvTS/m9smaLw+Bxj8EuSyfeO0
330UaPO2hypsIHRF1OhHlj+rRDfrMIP+ywi0GvL6uerhUq9NTcJXa/YQAZZZCwiItFFIH+rlSEc9
9gL9kXKudP2VtJYir6BouUPcsNgn3JWZh3d9l+KAG0EhSF+X9xfWIygTazXZMal7rJjdQP/qvRYf
C4e3t79Ow083a8SoHzM6mJbau3wMGj+wIqT7QEdnSaFlk7C0WmkE2ZoynT3aa19Bg0l9ytYwqDXo
J/lwmxFT+I4PMu7ZWwJ5YgyCH7/IrqP2pWxYIBlpfHtoSSRpxbvGagwDLRy5yFRtCimASno7+GCM
Y65S+WpNWQX5jfllggBnqsW3cb9rt9Gwbx+D2RPFgmoVTn+Y78EA/xkMoWivRVruM4kHNr4v0EiU
LtaPCjGWwwsPXZH1wZqfL0+8iexJcFhNwuytVPRPiQhFrWzpfyDyl6Q2Vw7LbtiMoE0B/wPCuEWv
4eem0IN3om5lI96VpWPT14CoKySbjyTitf8YRU0qZJX22Q/nUzHD9NgX1vmXiaOXVvO6buH4yqiX
gE42vIOXf1OA1pIY+w8+xP7kXw5F+Y0MyU55AliLnWQLy/f0H9SO+RvdDGBxTbuMX/w2SGTViByg
hXETpt0H6THGr1EbiG5u2bGqG6tcfvVFlYTpkF8r1ZaNoyzXdXpPgFRB/04CvU+q/9l+oUWYnByK
MnxNR2J9+wASblsQO5Jcifhe7s0Jt/vluf0CPdyTOk0cJV5PiD/0qeAY3faZq9x3zJuw01jU2mvy
0gyOc2c1rrDJSpSjArjFHxipIgLLe3ASjJKrMOQUarPxel0CuK/PaFY/vk0wHBmzXiOyIGCyklGO
MxBD9Eos9o4y9N4h3bNk/c9qWp3AsS4BsvRcJEJtDI3ZNerLeTFjoWx9eBerFYtZ/AB7P7csTnGn
gymx5QYHdkXymQzF25ddmCrNg2GoOXecDa4IUZUhB1C2o2jIjtZA/EEM9WVwQudcsbsCqHf9d2/Y
733u2KVnLdheZoEBAK/lO2MXequTxZPe4PRt5qLvyGt5TA+8lrR1OePKbhQ/obBzNxG8fZqDY7lK
izfgLM0bVk+Ckx15jPwD15obphQdx4NOVpaScoG0tPX5HkddV6Sj8xb/yObWiADI+y7NSckVd1Go
n+r6xT1Qqrt2Cnyi4NPfD35Vv6l7WP9qKy5oeBURbbZZxAlEAJZB8eLj6ZkTULz6thInBwp9v8+w
AKsA7CHIi+WYKlWAXFL/fM/nfPt2xIVL3hGDoICW14UmrMk2slWBbHNM4CpR4fkIEZBFVH6SAshG
BfcoCMXvZctaZ7dEFXYECz/dJG1aimC6tcEfcO/KyzJJqGgALN0nPCxVj0uenCNwr9k56ne5wubW
Mvq+zmkM2ekIZVjt8fa2IBjskme5gXYwHXr8I0A48zguIBTlpWVpJm8nWCBhaOzrJrozJ9fuH0CO
bT7GmPUIVp2MWfwrB8ROYG5f3OZWAGu03G+QRWChN0RtZ+MbXtfRyLF1mwtdXI74dlYAzW+ZBS2M
1IP4CMcTFjcElWEARcaQF/wjyczLF6YA9x4ZpKnIWXBspLvBTX4rG3aXNaZP+W10JdiOb69Kdm6r
rHqwHQbDjSaQ/WX83k/wRRJZaKBrmWLkS59GZKw8xa0rW7wWTKUCwgxKyfkT2izA856p7KF1mikJ
81+z0SpA5IL5E0xY1QKM33a68xjXwKWK4zYD39iOXif5hlNw1C6Uq9orP5Qt7b7Vu5TRMcZOrg56
XBnZesfHed0lQVtjy4uv1nxbe7cVjVWNOtONJ0BGQs9LfvLtcooDJHDLu5zmXO5z2FZw8df5NKMB
8WX4VFf6N09uQcb/0Tfsj0wnknU/IP/8dfsvyf+sapXUY6UALFUxMqQV/m4WOaiL634KzRVIYoTv
OWMIJAvTbEHZmWUMZatl+PD+ZXUlgMYtU/Z5Y8zadr95QFdJPxeyM9hDAtUKeSFVLnp8Eb85w0j/
XeEPgL5UQLU/D2wR/Exo5waEqloutOFEQTCZAWk89I/O8z4yjSqzz+mMah2xdN74LPYsbc4jP7UG
Ew4cW2JbGFxAoj351pfZrCwU2DnxTVTauu8LE/zNco61CbE3f2I2xkWfW3nyLWpzWCnK0X4WB4Nb
6Egyj0zpuYSeneZe+qcHjICHHqr+sG8n1kr2ibRYLbKVYqTSYGuVv9VBD32zLFk3n8+dxnixXrVK
yf4tWac///bjdvf63G9ulHZz8MhO4YOyNfkEsJWgSkMUuPws/MWfF+SxhIgwj/ts1ZGfNX+OQ8KO
Td1/u46jJIYhyiYwA6Xnco7qNLm8OGea1q8MXiz36c2OUeTitpOHmO9i0KvWLRc+1kzf4fi7+1QG
KLRQofzaUexFf16zBAgpM//qPbtA1aCLPNYB8ocpmWglJnOkYo9cmOzS798q/LWzewa+nbXYhKnU
oXzvLkgC5x+L1MI6HfcDsTbYSX33K3HmZku526rwUJcACU1UxtPOq3fhprccR15RmJjgFvcpjABp
NWnhtgamvj67Pysui8EpOlVWjlONQn9Vz2OqfIG7rW2B7syGaBVu0BqVGSZZgYNMcfAJOOZOCaE6
r247fSotqlTdQvfYdVnxeGgp9ea1+QUsVIVN3hjoBPIOoRSkWDj1Djoy4HKRMDvNnD0tFVXBDXxt
6GcfB25AQ+2dHQPhknTIsCcSVWQ1uB9P34vGCmSjzpu+R5W9ADAZ33VRu9G5VoTq9qc0JnBlJzyI
Gz236d/8+N7ify6SIazxU+2y51LotWw2Xnovin1wEXLW8+m5rpLY4VWIhXX0gpx1kA0x1DgFtVnM
qA1Is08CL8osy9EcZdl6ZexoLL+cRUD4E+fYuQXktTLOsXE3yqIKhMJIU14D4j8KS2jw98hLW9fw
08Z4/yOF0UqeaqudQufKD/U2/qAHwuf+xdLKLyAC8a7h/Sw9jsTZS13tgaPil6v9czlJs+603lR7
xwN48bK46WxC91yloLmf/avVwsNfq5iLQfMH/tcvGTlhtJs14gSWzUu4AsTPZ2mn/wwRbadCjvLg
E6R/pr5yPacOJEAf1kSwr0pmcBm2IJTcOXOv7aDqSjXQ5q6Q4ymVPGUtNZlmOczG6duXMy45Ux00
R/aq4hhaN+SHQFJ2QperydH0KHoiMJEKt6kekZn9t4pbSn54J51CaPjtY7CLSiFLc9s8S3hEi02Y
DL1mut6QIZPtZUSQGLYqfcWoqc8xWA4vwRRS7C3/uNSB5siALCh9jH/IYHwavk7hqH0PayRkeDOe
gHBKt5nTu/hRSsho+r9nf0ptPCVTHgPs3dbrwNsAo/PpeF/UNuyEAtfaOzLZoCR25PDY52Pt4mlg
qthQC3jD4onanUPXW0y3+2fWTKlIok+SJvxxw5iSWudFSm5EwyGQ4ypuJgCWkmZfxFNbPgfruGVQ
upQdL4YyTfeYZ5mmdCYQrLGGbuW/QE92Vdu5dgY8NzHiXavERekck2oux3VMctfrhL6vJN5ehN3F
5IGG5Gfi/+n7U+wWdTgbQX1jKk98DfYZY6054+umXeoEQ+J1uG8O8n+SgxuUS5ANW6mcfHpzZQIY
7PAsDE5aUZd3N3QBic0u/Jcj5J25iW1wY05k/a1KYb95VhZX2Ddn3tR+cqcEtgkZCroaokHjukAR
DTQmIM4WpkltQr3b4AgrjQp8M9fwIuCyvswEO/bfCaA41pRmgSZlEVwtOaGuT14k1B2/qzqomOnF
cmOyMAlxO0OYlAdP6GNYRx5RjxyIpklpfBZhNZ2swDSIY2oZ551b3hSRiCKUhhGbr++hVCEYczwH
/iUH7gt/9kE1WnEF2VbuzzCcsHpKRhoB7RbCuA46ogVSdRB0A3rNN8dV6ucLxWQ4155rujKsYhYu
AGiNa12i8bSblvjc9ky1DE8/UapzKoq8+Tcb9lQ+UXoQJe0z69ahw/x4vXqCNE9tZp8eQLk8xqfE
tlqJc2+OR0pheW/fui0FKYsIfpzppYtGT8UFwtNeeuWiMf2JdDleMx9oWE6WpR5HDOIeJSNiQ8P1
6aJr1maOWqqRbIsFCAkttSCTHWrfhCiILozUWDUVth3iEUwb2KVfonP+jAR5l+YLq2TMKnRiDv94
G7WsEez+zWTJgmqcYNYl560EFidIsLdBeoyp3dMuSNt565KblQoWj4heugMDGCKc6B9Ncw1hEHkU
5E/ltoKswjZTuAelN9nYdcQT6rd9A/Y0VZtJLBuVbIv8C7Z1jONHJTQ0ig/yQz6ktPLjAofosp64
LXEK7QPoguLwEecs3Ie5WmCYdKhpwTaW3F18BtLsXNfnQksqu15E/p8d34IUQIDAmWYZWvWj54uV
ckzF3UhqVxm9/n9mDbUfJHVZ+bPNmH5kSLbocStGbyvindSzogvzgh9e0H7F6LvcDFZy/Oi5WcM9
lNtq5PdMQReUVnvluCGSPGe66ppcjaw6Q5eyz7Z3Tz0NjDnI+CuVjLRD43XWc6UJm2GMsyhgVgeR
5nduJvdgrH47VkGEd/LkoeIXdBp8VNylplMnx75ZGLs5f3UXWXkfeP8sBtfmQcMoBaORJkjHPnv0
wA9mP6diutRbciUKkWArXMiRbrP1DgdS7eAJliJ/k71sebfaT8JXgxcsWjb4ASm7/r2UAWhGQRbB
khRKaJRn+0N/lRCH3bapzRQfv+3EhVmXqs9h1q2KT7FVVikNRJCy1LytLb//iUSpvNYZZf7WYEaj
vSctnYsgjlzj9l/Vhv0ILVm4By9CGQoG2KTmXlYtoiZbmTfVXEqJYKS3CflTgk9KGg0572U1k/zh
0LO6iYKBEENxC+ZPGChs+mOBc4YlGw9d7d5aqaOOt7lCR8HmLH+lPHjfXUDrVVNRBhqXhvoy8xiL
LgAv35YXY+5SeeCaVdcHCu3sgzk6txnjjeEx87ZbZCa8+4dK55S5+5i+ylgxJ1n+o3OeU3vo2php
tfd64h8rQLaMi/oDD6GQqfYtHbEh2exBHjrikR2TXWDaW+rjkaKJI2ffLWOnZuN9Bu8Q4J9g2PLf
k64fxP5DfJmfW105jCE/xZUEztzrMieFh408WyKHLESsP0LieK7xY6jT6oOjf9fdapbrzmU/FE8V
Q/1bM+1/FgMvsR+O7Z1gyz1ijd5tp0APVzEqT8PjSpvq80x0+8iplG2QXqLy3M5/NTU9iLKoCfrR
3dS35JvgItRQK4OivbReDR03En7Eg1temuFhvEVeTB1+wIGpN0ItrqGLP7ewyMAbCdUeWFS+6GFW
P4/zvkCnh/0LyLn7YchneLjp861ia7C8q4USFhKyBLZo/LNSLUjbWklPYbsyRU4f272UuASAnUtC
4SCdCUdEfOQhVjvTHJuqSAzQ2I4J67kkuNUKwSLwAcCNlFwl94NhJFYl77/17GEMe+OxERIjgBj1
U2gGd8iahK93CFvtjOMO47GStr29Q1gBngdy87fBuvoziczQSJIJmy0NG1zhz/4Zt2J5AaF4z5nE
gg9i90q8QGKb/uNukUwkuI9VreXjU6PjxwwFQdeLUk2Ybl0nxdJkxy06aBXMwuUDfMz5WshwxdES
NP96JntQMoDqUxYQQOBf/U9DD45xJl50R6RHuBGNWgJk5Tz+179QsX9vAkeNn2ClT218Zoa55g8k
2rVTwlAKdik72k86ERBYKXDw/+RxogXYLLFtBT0fu6MM1Ued6cX38ob8wUpxl8AJ9sgBM7bh+b1m
vD5tiFk1/IHy9T5w+ZBLbPaDDnDKddwaXPbmPoGCovSLnJQiExaFh+QrdchoNJUKOg6dDmdbA6JF
mK6pG8XovOr0klXcU7LtqPSy00gfFH+8F0Ua/ByiKKbAk9qsV4bIVXH3R61XXFyJaykz+nJvuBWd
1Fc219CHErTVqo1LieFNttRDE33zyttGaqPF3zsjlw22yFiXKauuGvx7rlt4nNqUthVfe5hxepxr
H3DbvNBshm6wace7ZmGsp77fj/KB7Y5ecpv4DpDinkaUcFnEdlhMtS1ZzWzzVfSGmuXsHLvUOqhW
b/56FMbQt+vD/ANrz4fckneCnSMsxPq+p2RWXJmhxOv+uxV9F5ISQGbjEM5GNuwCzx1HMuZyCFZ8
U6dVCv8Om3GDebsFfr3RjKdEczBnzs4Etm92UWtvY7V61JYW+4EOmGNuac9bs4FRYfKfgNPcGkby
5TYnoNLEGSQMEiLzeeqDZnv7BkatG8mzde6r3rw4RawYoeyEWlwAhGQxuugwBoXRf1/BQZUyunyv
T1aRTMisrg9n32T3bALhkiR3SICRGcV10Rs963oGcJNsMhYeonROCLheIFOK/Sc52Jr2h0GG+ZZN
BuD7BWTVfXNxg7rf0e0yNdWBR7purTzN3HKhmHpj3C/7zfcg6dM3HLMRCf85+EY37b4CfjkCITb7
lcHLR8Owu803gGPjDyVJq76MzEL35oMCXIuRadt4Dja1t5KCG66WBhh1IzN23rs/qslX+f28rRp7
taZiP4ynm3VsdxCKTPLNPdbz1cRS9qTmcHo3Z2EoNroUicwfKSC/f8hD+qSnBzMZDrcWHcaYKmjH
j6mzzbvc0+uLPu91pf1Tv0ovlt2gZdUlcM1EDB4ObutGv6oEFxazguqIZyqMwng/Zm5NVbDdvSN7
Eq/g5mi+3UxE6CeXLVnXEKXbuX1TFNj1ABLBuO8gRlvMf70LFm5oh1H68TVwJcuaGFc7aKFF+286
ICfas0nPcYc/gidMM4W0qGXJFrBZ97CwJ//SlYjU3qe0XBoxFrYm3BOGMkTCKqWYznvXz7ukSvFC
/r10Or9dheipvx+Q5mZIgzRcnWW9Bf7NrwPsEr2S2XkTREwSHY4RfMucfyuKNkrQQwNIo/JPf16u
yFXQitcpMDLrIv+lBqM3qmtDhXKd8MuUs+Se+Qtsd2i8pIx2UifVXzxVvSioHUi3kx6GH271uojy
a8SwVdeSHIZVKero4WaLWov6o2wwRTK8K4I5/QnuNXpMzC210lx3iUFaxVSHIzJPzB3ixsk/TEfi
YEx3yWasF68A4tiXno35xFUdoCNphV9ze/Xb+tmOSHKdXlIrb77rq+p/L0KoDECZrj/7uAG+8pKN
HSxs2tEEwH3p/189dLMgMN7lkP+QrRMfqVPkl23WK/TnF7goA2ppU0RY6oVJldW4Q3UnoCwbmHN/
we3uuL+QMl9LLzz9VQ0vOxxqcw7lDeoCSBhqpwzOWlA1WdlRahTZ6+hBziSFQNQotXSHwg0OJvB0
IBUt+csUGn6GK8L/pYWjRgkViRqxX9Uz8pisWeJ++SFrs5d0UVtxXUPsA2y6FI7cYiOS+uD411C6
+ygcyGX+IfFtjp89WLzHq1XM4E0LNlV6ABOFjEJ/QOpnrYOo8RLqmKaG/HZ79XMmEHcfAaEp1FuZ
1iqNBreszHONzSn7vuZX7Ghj+QnGU7gZMB7i/jLMoKx1SzzaFmqOyrsQtoPYS9xIw8amySeZVUOD
hX3VCMQGG1/63azFIjql82kYruAZPpLuNsNarhQNJ4CbJOF28h2JYzTvrVY7ygfiL3nqxeFC7DrE
BT4v5VDyEclBiYjzG0zm+6WpUgp7UpANNhpD6BGSM1ZPYGKtFv6yw3VrvSoZh6Yqu393Qg+z7erH
1u2B28b5P/OBFyTGzI6cIy2Yi5udmpw8++nZQ3tJEsQGG8x0q8hLOK/oRRYeMadFlTTypBVwWpnR
iUBkxOGWf3C6E3UsQciDBYoFrdFDjH70UvLK3kuvFIzL/pcx2DLrIrCWR7jInxoKDEDVeWzKvm0q
Ac6FEVesWF3GypzVseexUAdp1hUCmJRv0hJvzRKsvWArBkRp/1fWppiZSzi+379m9dFXjqUpmGxv
gL3TteRWtBF7pyz5QqKSKH9PDYwrRi/u3gzxrJMuJWd+zsfeMudr7+J0Um8SAUkkHvUnDdYdqTVx
/m3+fOIBYfxKw+VtvzpyerJd/k67qpS71jtrlw/9pM6hx5iojfMYJFUylzntfX30B3U7CroSfY05
rXhImdSmQz20Wk4zv37itZxssMprco61FpERh6kba89t27DirZqidLoKiYpZh7M+96df2pE/THBO
HBU13cDVh2VQE0Gw8jF6cz9vsLjkLwQTuXQJDLWKIslG7XQwUwSWaKlT6wgaSkGsUAs3W3FL21v+
I9Bqvx2x06Ch5fOq6ZCDkb7k9o9wnwa93mtvYAz8ymVcF3g/xlodpENuEUm3WH/cr+AroNta1fAB
8u1kD1e2LBTzhOnfbad2ihICe5Xqe2J7Xkti/rDzmG7Tg1ziFAKickqvGsM0AyM+zLbYNxnJ5ymV
UDbxwNH9UKCbBVecfwq1biSsH95LHZmI9xZiq1U+IdVGz997HtilLS1SC6amvTfMZD0v4dzxghrV
YQTFj8IgRKXnLU4qHqqr9WvOKOEDYY4vANd81c+ZWDawte+x2nhoGVOl8VqUuddFb4IPqWzbFAaT
POG9eybij6MoEbLr3fjZIHn/GS2kFvCp2lhxDDMgZjgbuocAH/OrLwtjf9myAnd2b20ClbQ5Nipr
BJVZ4LgZkcr1ggHou+XNVny6SlUyeoD5n8QfcTEDjghdZOPGVB5iyCik8CEDkn/1ScZL/PJnMYU1
8EPS7iXTH4Wmq5gc93TmKxZapbIXVQnlsduDZrJuHxyGmQ5fsdpkq3YOivqX+qGjBGfgvmpAKgr8
/phFtMjZoqR2JfUE+Q/KpR+dI1/6nb0D0T+B8PIdYVuWT86gcpkpsp499vBHkT/FOBUgVBuwUIoW
oySLVwT8WJx8pCC7W8jYamOyJadB8OvcTrok1PbV/0iw34CK2QjW+C7WFO9DJ4lTZCLAg0KHL3WE
kM48IT8JehUjQYGr1lHbkrv9U3jNCfMie7VHsVrXp17Hg+RS/wexwMdlsrkuwRTf5NLtvSwsDIKw
9rQGQrqDNifLqQxs++7KzF1xXArg5gAKCAw/0o7Q4C/HvBv0IkZ/MKXIAB8gsGAJxogVxYI3eram
N3AAC8DGCEZ+XTxA0AEtXhfrW/TqtV7lKZxBoK8zpAOpq17Vewwlyx5kiZ0Ynr2CDXDm2EwnZWf1
t1q7gtH/MDJz+vQPOX60ThTLyz8JKmoWisf6/AzgQafPpE0L/oe8zjoKdn4rVCnJsBkiq3ihuO+Z
ERYYbCm/olavSznEgfQUXl8iHAAXQei1PMEN6FONZEKb3kUwTQ79mnL9YrqlIczW9weKD/U1/ofi
Oe9VZkcUnSHZR5SbStz7hINLNeqtvb8invZuPjl3fcVPaMJR+5BqaYpsBM9I9KgyxbeAPpVgFIln
vh9NMhCnmiAUj9hR2PtlCOVFqW69VTQordeurbvU1KtSfL6L55F98oYcn46E6NMfiu+iT0SnFm45
siZD5YcaO5Gt6P2erxpbJJmxHijxdlQBhW7rdehGSaZRxFueBnsDikF2Ht2bngq9YeoZlXjrTsGj
F7CaNE0c6kOPpgypEdtReQbeYEC6zariiGv8yyJjhlr0ikECJ5vsYBe70Y72OPsnDU/iEMHlP70c
wONyr8Q5yv7suG7HUMPO5na27vpJWK+DawhtiuydfkUmAzxtoa6W75qhU8S0AIjQDwm5UU5yYECc
KkREYrspGFHhgIz6VATEhF4x7NTlsp8CAjzJVaoF6tf9pH+H4oY2Hjbu+6qErTBaYYGL7QFImzOi
S+DtXTAUOkGpqV0YtkUQWzbh7gkS/VsPrCytkpj+C+z+I40Q1QNuBkD47wGyaYtZoBNkBQ86XeBz
+IJUKLJReUetBzZ1eBX18rerjUk/SeMY1YROFEVqjzSqBSufBabJhby97VPtEnj5nsuwenWVPeTi
8xxIOhFTkfW2rg24BNBhFQk4eYTWyK9U33aISgP6lD+20XB08oEfIIdvrh3Y/mf5BYE2ivFzOPST
8l3r6lSUYMgESDotrtxCq6YU88Mr8WrfvM84vBf+O8yERs8B03v0h/OyaRgthGGJ4yekgd2f7Hw6
IER5L3yLhVlZthqLaCQJ4FcOtcGoHTHojevAbuyEPNhIVzILKrHMt1FRhtaTH7kMemeQHFOrOIu0
sIGQDXOHd+8M5mUpJljdhW7lxg+DW/wKkRd/h+IUhNI/Rz4ARn9Opax7jKtC6qvx9hzbCGoza3ek
ALaRjU7nE8p0co3r/U7cBFBD85spONHo97WyjZZ7Jx79lhayPhqFuEbjnrzB8iyE9y3efKAr0ImZ
Ltd68e++vcY1uaPS9x4WqXJvzLYFwiwp4Oh3acMnZsaX1IAei5pAmgbVEStc3kFXw4b2P5Tma4Ze
EEs54V+6F6JCnjhlRdP2e5T2BYVnVnhnDD3EzpQZVkVPIw/ppoL2hGPXe90ioqyMI8om9vJqPC3j
8dqXI+TOPVaXHLbrwcBri3ZraLDUU0372yERXJ4D0sr8S+T1pqRCJmQdGu59PdZUrIJDKUDBBBlF
8zPk7JLky6caEftNg9UNmk0gNVOnabdtjN8BZlss/76yPmT1oQgMi0hd0ogRh4guIkCc3ZB+4dbb
n0BQuL6t5jkqfrF/YW6a5b8eryBGf2/nyVtz5Z0sXf8fN0//hWYS38b2kn/kSBP5JcKhBD4lW+zS
mmJN9kYU9F2kGt/nTvyEbLCMOPHc/6UCOlTHv7+QP1q4rcUewaePLwaPBj2Eh4aqNEfmXUI1kmWM
IW/v+byEomsJxSCOvJl5Mb21hswByQO/tAWXibtqirCbUuA3Tmm7uPHg//blkV8JgC3v2Z0UN2yJ
uqi4vLLBaUQEPdgTjgxFAxLlf/wuu8uvkeUA5Gsvgour7tVR0R4D+DKF856kTicfTTLGp6VhdNTj
/Lw4nUiBY32KF40kkM4JJY79V0x1/ceBLH4v85y9ahOVzakS1wbiYcYebi3f56jUHhdq8LjGVXSy
+HuE6aJKLqifpXMTOGIliYws99R60+PPPARi6/SzwFkf1PksTKZ2ZWtBlh5tidWIHLX0+ltcBSN5
oZmti540Y7A3iELSqffr2s4QYcUlyEONhO32zhdwZaiOzZ/HstQsWQRB5LvZLVNjMCXyk/vNoiiy
EsZZNr/Nzeud72OB49U/rakyObTZRJyKhYFiVj4T5MSS4Uy2o5F3o7bjjKStiNsCsC8YiUB/OuoJ
SzkQghuf9SUzaI2cBylxRUgf6fUeYir6gNMOgOG6AlYZ2YQxVoA4FrMwQkD9VY/H7KjaR/n2t1yE
cCzWWOHqtGBCTf6TejAqvq5Qjo35LmuEPvUwgq3EKlEo7HgzjXz01pnb+BCYP1GsQg2zuEAtXLLp
Qu9n2zTm5CgJnbUI1X8RmBO4QujX9BHm/5hMH50jIU5P826ynrjv+UNhcexVfa+R0V0hw/3MHXuH
L683QEZpLrvNWFuGFlTMSOYGyqvM/YChxw/rfMiUa/DjbIDxL7OyhnfTJfBg5PJ0hZHiFZmN4oSf
sAGNN/lan4zDlr9ar85rhJtd6qVGeCFcvRJUoSaIYOFvdj8lA49e07Wg+aF9XmoeZjwBcaGQTfSA
Ys+FQXr1mRJseeZ9fnHBcxG/VZ3XZPCAc36fTgrErLER4JIZNCbb3BrnL0ziDKKyQx9ys6z2iTCi
iUymHHs81AV0ZyvJvJNncxh9NDa4WPzUbl4s5f6BDG/JBsI8+PFc+2Z04034KxHkqF8mPGuqDKWX
drns5MMdkaGMKkClVfcAPX19GvkOt9Jt91b0h2kBY3c0l17B6/2pE6pJ6dyz/pmFY1ef6KX9jxZ8
P0KVJTiXIjvCBQQHp8blygsTIr5v6s1n7F2sIaWnP7OXzUwK+V7zcSnWlXcYTYDBk8pVn57Ek23W
DbUWEqftV0wVs7IGdy/jR4iDNGRpmVruPk/l5TTffDeEOAI6CQUZ3oXwfBK25jJTBxhCog2+6V0H
p4obz04qAXY3S7IATIrve8EpFs0zFOwR8wnaalqD6HR7l1Y6xqlXa2pQfQzYEopxJdpEHtx3d4Dy
FKcNh/XdNAO3i/c8UsjytVyw5RPsqgm2ANwrEP0G8sgrdoTjuI0yFc1XA4YPeabMn9j8LQRn4ucE
wAZDWmA+PxRGnJrn3yr3J5Pu+a6FP+FQwtcCTIJBRFYHotjHn8IF+TbzqzBBCXYbLGHAMRTTQ9J+
hNkgLEEPCbMZ7dTItCofZ0s3qkL5V/NtLy/TrgBP41ovLqxBfbEz3/3uiC+snfDGIySqx6S4BIOe
5+ywEdY9Y2evD++lugs1ttysZENXMuCp8lTLDiPyJqZKSlpJS7BI5TvAUCFygB/+pEA7rcCZrGYZ
3ciiIFljQWf1bZdtNjGTKuqRs7Z/767Q2/iZKpPG2DyEVgt4n0SZGG9Dv9RHjtxgYuKUoGVX4xrM
9TAzO0PphSSwjPy1s7UG9y9q0q4ZWFvSGD9L18K3xlHmnwFmzfrmReA7IqMZrxx/ccpeP9UTmG84
VMQ6ozmLjQfjTebRZd6xeZxcvobv/kEDf8FbPJzTimcwxOi/IayuNMZKtYVWJAdoa91fc/1wo9Cf
NN3tqHRBxidUu9uZ+8IL4ZrcI9D1NIvJOBDzT2U4XWchdH9fLbaicUb3JB87RGr7TxHe/iWdaIUD
MTngQzezAE8P2OutDDV8XYnLMnUqT551+aDN2a4YwV2vWupz3leVtsMjJobCE13Llp3Pb8gV7/KC
xwqWqj0V69XnnqFSmlE+FBilIx1hHZk9UIwrFYzDd6RFwjyugPjxSPz79kcZwcvGBa9zgY09R404
gF8h2Kc9a6mwsXFO75mVNVIwVGXUkbPOsHUg5y+dJBVxN5h6Vv1P15j+qmJ8eCZM78og0S58svlS
04483AxcDRJ4nVSp1OBf3J/fPKPGOPcnMHO6IvBkhklrpgVkMTLStI3jKrmZSsO4f1CBfXqVTp63
hxHlF/f5wzEA7Yep1j3N24QujssZ/vIj67v3Um5xcxz318im3UBTWjbkVAyZVC68Fqf/90so0jpJ
Yobtu2WJQzig1ByH6e64Yn67Ycbsb/MbJDo0YqYdyn0H+ZumLmXP/YqeWGTq1lKaRdjOnMJ+ufYU
I9Xm7cOE+G3U/yeV6VtZUUaE19S4ECHKQ2KiMAfPu6WBeAnaPjJwLILbqVNhY2GIu+udq1x7/LVv
3RK0FsdwCSjI5QwTOsYNu4+52nNVRNtKfviDy5K1QzCnZko+8g3jJWa6tTZj6i1OjODdOT89wD75
kJDQ/59fUuCwftQNKL/AF+3xSbdExtcT2mO5Q6vabK+5oh5F6ghHYQT7t3Q0t7W/Qle/ZRhGjRv/
DwupQW6+NWydAtM3+NgCz5pzBEWQ+3vkrImV6YiDKywh24m0B9yUTOH8/TLBXMxkqAsbC6//Retu
4WsLrvpG6QyOGi+qhoC2ft889CgGGzGI54DmPZK+G0BGyVQBjkB1idFk8hX+U8nla6+8tznSfQgP
mUY8E0uHYWXOu/bbMLcVMKX4oKOCx/aM+LzfKbnXMXQbcrat/krnShD0oXmJW0xyvHunvdc7YbGn
6TVL2jvN2WKxZjViHd63HCEbS1yv0EEyKh54RjU3TNZ99jpBP6ai1IaN7W01Oymx5HzvqLYS58/i
nqkIF0gGI9IKSi+IuOBDwpLMdwhlmxij6PqEC9ikw9yPZOf7PSCRsGkB2eGjYbpbD1yziAqfnH/j
A7a2Di1WdLfbuJX9m0gsHnPmzedRZAtqauLHiVL60DeVNbB4mh+nXg2nPayYhBdR7/TjaKKIJXAZ
7kfcxj0UTZrlrbuFpTNIcdH/xrWXXrTtq5d47pgj38wd4Q/ACj6rMnE7COMWhS2CrgTCOOB1LvTq
9GNUt5gRvsb9vkEvt6OmXci/7eZTxakbBEwZkwIimagMKJzw30l5NgwDgRpcyh2PXbhDdcr6x+79
6NpyVoF1bl4h0bvWBcYRVnu+VDBEzY2Cfe09babi/R3Q8c4MJW6jcciVKGkrllTzQWqPKUG7RDu4
ies3/1a7CLjjSLcM1do3ctSuYnuARKdy6F4o1gGnU8HKv3ZNet4nIiKuh/O479OZmbTdbQ6XHBCH
jdYW+wkP6SG2mib6+oocaBxrOoFjDrjMAZp+iYiPE/Vc9Gqq2B3ueYr2d3PKRC7RucIfb6cvAYYT
P29z4L0W3MrBW/0tyT1W1gln45J19mLIkZ4G6SfjEtwtXSLzwjiK23XTWSlK4mE92XYZNNL4T5At
EJRyy41nrGycNzzWWc0+4G1cMBmEJrvjgTvi689Gsq1dPs+qaCYsol1+51kmROL7+J/Z1cbixWZl
VeOhMndj/UoKpsroLMptCPeuAZWxG0G9wNeeEj8hJSbssO6bqJ/yqrpsRZdSJVaIpIuL7f31zXgw
+nDLJQ4KjQGr8EVZ0eshzbo09KOBl4S1h+hP7Q4QScZCskSon6aOl66AelHhZq3IbZ6ENwZJegRi
9QjtZJpTWeafAfvaZIjm00sN8yu2zdO8CBTEBddfMWyJkKyfROtheAUL/R8ZZoib8bBGwuaT1uI3
S2lz8A/eALKX9yO0+egPF0uNRUf0ljyNangL0i5qJmsNoTTtUF4jR6tR84iQQxixo3TFxKiV1Hmv
71qB0VPPN8nuKFI6MEftOA1WLXaErNym2JNU4gZB8f0tRFG5dGPPA/gMeRQ0RtPqE2MuI/iyT8Aa
5IJn6qVQ8y7veB/5lYSc/KM5/ln1i4mTKEEBEnfH2AFefu0vjzmLc1bl5uPUpiulSdg3F5/ycGT/
kdVfRPHcP6C9VLs3oJnIU1cltrbxuU3uuUYBYQWztlgQiN6Hdg2Ad8sXx2AIbqMWSA+wwKwrEjtL
8opbCF70tfkjofRS9D4Hun58BOyjvAPp2A59tl17+2ZFtGs1nRrjenizSZJeB9a7QARtDm5VrkBr
7lAwQT/hQ9yArmMEclWplz9Q1/llzbVpxU7mPSesF+fFInx2srtfSNTXZiUcVbz5zZQ+u+87309j
KqOucsnG0TbdDpoATsrL0cgIvEHAcONsedAR71B4DroDdyUJEcbRHyD7XL6wV59N1yC9urxfAkMS
byuPySb098TQunwl+lJRHIKc5Kr+U8n+/WbE3T4kOi/Mme7AbbkbjdCMXMpjv0zcx3AR15ihB8HR
0ar7mSCK7EEWJLM3pwH++3kgXCpORLA8lzIt/tBUzWTd+Ygjy1lP59qBMfljXTmS3g9JAsH63TFo
OsZU1bv2V39LinbIBAmvD984y/NqVv8xXoIapQAts/gUwARUa7KkhJILGIA3/p48Sgb7G94FRDYD
sWnV36uYz7YH6up25mcrsDteQejIchlRSXY/5W4PboYeahyE7wr0ued8NgRwJKGbKalUOIbJD9ND
i8wyLp7G88dnnhzYjCojzcqHFYn1DRFcW7K2DMweU/8xYHPoPV+0MXnG1vgBuF6sH3leqq05uqAu
ZwiKmtgRmmXiDggEx9Kx37QKyQLewRSKEKC4FmwvNMUGxG5/Gr/SHx2b0PKvsmE8/m503gYlufEd
tAqwXqrfrQhsGIJtvlsFIOBS2l8/VUa1BRrJEM+fsESsuZlUkvdV62tixONCAR1D5StmUw41BHmU
oXDG6rqqm+CDCiuA+sKFXhHk27YkXIoegqtr2MZlQMzQM3MQUBHNs9FIXDBy+XOAyR81tK2pH2nN
xHfmw6Ri6QAhvfbLlugCIUt2SoWWsr8L0hiIY1LLrOg6lFlnXtAnwfROyqxBAW6FGgE55r36JOhP
tVTFrGYHmuxv1RBhdFhwkQQ+7zV1HfrR6k+dLEQyJfEuHk2n1V+aj+FHJE+Z0FJRv4lTLIvCe0+x
bHQEuZ/Q2UBzV8dyrbd07zxl19Y3H2YTeHYOD8V7afb85vE9//p13z/aEJBtwVXf6SHI86NXkCo9
XrH+sA8qvGzXpn7REGi/rPZQjmxgissPSbu4Z9mpsBIZlVGgGMo9MUWtGLub+o1DahsVZ7pEWFYF
bfo29JJ5LBTnfzMWfa3eNm+J5eBnJthAVBKHXp+N+6D1AMAnPXP6zxPe6tjnaxrPKjgB02uv5B2x
BlURsW6ks08i+/xD82+qVC+LQx6kuNsR8y5PfRadHpxtoXN+045OV1GT8SBOtdJo1t0/Npu20WTK
rLc5312iwdbeHpcPQjXWdFRyx9m5YyqXOm94WGF6BPmTMdqNxYJ3jShF27i6Z/1twX151Am/dbLq
6yDp+gZtaUZH834b4TXAv50I4uhVgApDM7oVb+FD/zo2f7a7GNalEGH5GawXrNdJ06M6uv4kQBld
mZTqNh41F3nvr+2NxDjs5Pej79MBSpttYhLM5S1nVDGC7lJ1/+XgRys6yC83cI8Ofjc943S+EL7u
tuep0AiNkFVHm/q0l4HCsZY1gkKjf02X1o3cmCLnBWQHcj+/yzFzUsT1zQ9cGt+7A052o7xtewgI
e4o8RiCx2WmM52pcM36hVL5DjIcaDhP5J/whZW1qHUwvdu73CBvhCh1BZGrRsMm86d1XilAGx6Fr
jIm6agwn33MLDHzbkqEDRMUfn0eSajV4g3gPXLBWL7rWbvMMXoeMMwCX3EC8rlN6bof5l92kplT1
MxFOKESoIn7ijOJc4diyxfzG9AO/SMCkdLu14wKinWzSbChoT5Cz2j2B+bzip8HAQIY4VCk9+Qxy
1O051dUUvOZy5Bcaj+gGnaHgi8Yl+9i2mTRkBgAhDtEJnghkBWNXAtUH1/eDuME6XBGEoocZ8oNc
vU081GyfHCtCXPZfPJeR66K3IqbZovyETuMd6lo7GDcL6gt9dIbgQ+57g1HgQ9MIja42CDb+RW+V
en1xtaELoV13+C4srpan95A81Iln6sRgHg5vsAAgyel155yFnCDl2RU/CUusUQWp89xKKzeGHxWJ
TsjvaSo/2fkhPmziDJSnvqslF21Kt524jhflxupCi8MUCMTpyi27NAUaViaPDuDQq1kt/SRmAw4y
/Lofxdd1J6E6PGqa5DTu8T1LxjMLDnOQrCxq5x3brEg+kNYaZirEh3zS6MH+GRgEdLtZ05GFOuid
Iq6+ZXJz39bmlUwBR+bBIrlhOV/WV70YzgLFgIT08u9oLE9gsb4KkQgoQvYgnkn45k9ILgSab4jp
GydXE3TeNuphcwKrkeB5d8XbTlPWjiWRevpgCwcajNp1Lzb9plsy07YXG08bDk9cP8xlF1ujd7+1
YSbVI2prFzNo+YZVxF2mD7vUGCCNvWf1UGEYSbAAuiQB4VjozQ/gaVCktCMpOeZVetiatSqqNT09
h/9nRfChs0xbydgcm2QfW7kHvNq48RzCQZ7BDmXQmTHJHMvpez+4iY2WLAaee8I3Vt3v2wBPam39
3tUubvBOspXYZhmDouBK+eYGNfoI+9/fDCRpoVnMlt1laz+PA4JoaPGqScrpVF1p2KCR+FX84d8x
m2UryIkctlAx6v0bs0jMMagRG5ttIynjFiR9IAA0cDp+QV69BoiP30j644ZmP2Byxo5mBjWFG6G8
8SlpkeLPQO/VpmE4fTkeITe5kKk56dt7q1AxeznQRta3ncCeXPU6WfuOpeOOJOLhfBAzhljxtXFj
b+paCvmuTns8rwahDcSEW6a8aCBchKDpS6okEaMpZk0QQFUdFa9fNZdv3uSqOoU6UxMaWieoA9+s
etODtsftuZ73pvTePVSs86RdwiOYqiIQZT6MpK5WJLL013/l89WXLGi2MQiaZdaqsKVg2GIhNsY7
75a5dk5Ho44+E2afksvOe3Z/rOr42TL2QLmwtDm99Vbac6wILjtZ2J3h+Qv+Ic2xxTpCkVHefrSX
ogu8NvfZmM3Hh5tPCpwDbgswL03ahL94xN0IblyQm1OZ0cVZ8IG1Tq0En1sPN3IHTL3wR68hjz1J
8FCgWgJRHNBhv2Z38YJvYKXf/uuU2aEG2BfRjjG+B7KGR0f3bFz7TLypktNiHSuxdrEf2pMDWygf
PCg99n9QdoR0iHZsD+u1Wdqu2oJF0XqeN1dN2sqev4S/+olJ7DCIOJi3rYl+VhN9RpuvI81JgYD9
iE1CQ3AWbXCS1BArseJKL50aP2iKDG1f0I5/hEBO/ofuLo13FgLZ0vhLUnCJWGV8HOKMmqRdil6/
3A3u/E695KLeLlGpIm1+fR1EEZr8f1mi7uhuFTX1o9haKYheMgGx4lhMGTwhXfumLqTBBHRH7dAV
zIWrugv7LaCg1NUUZUU9p4ZA3MXob+dBOe43KnS3ApUqFfD3MMgmGulK4geKszQNDuu9LR87Z3jX
VHn/h0Jyu6kUmPDKSEiTLK4udehg+PBv3EFqbkD6A+q339r911Wx+d7yM+yTsydldR1AHFmxRmix
x4ps3FYrkG8s1I8xd1GapFPNznYvv84AAtUFazuOcR9c0JyspKL7vpJXteGkmrgthGD1N8rUHBgE
4q+gidANWSDHLrfYQM1JLq0Nnx8j6QnCXSNbyywTHR4WpxO3gHJ+ad5VWSPNmqXlmHHtKblVg+Vg
OU0fxRCk3rK8xf9b+Qn3CLUJru7snlH919W6DrdYgrKlYuQ6g71A4meGh+BqJWsrYYnKB1vXjn8u
NBIibC03IeNP+C71XGZTh694SX+5edxSawx4JxvIiX431e2Hs57poYZphuuFIldiOCmYKVNaNIvq
xJAM5jST31RPa3MkcIcklhQyRgsSCd4ehNBFRvjLMy+jncbXvDuXgqEUslFhqS8j1gktc303nUrN
6Zq7cmM75FqzGEqkEH7NduK9/Zcd31YlXQBzpRbB8NXtyE03ZrhonvLojnzIFhSkBSU7caLnLHi9
+tJogF3MfHHsAx2WjLTJlRBx7gJEibeEZs7IKnD3ihCbuhsRdjRTYzctvL6RyEtXKvZYma+XGNMR
wdaiRzecY826LhkSPdWCiKU18wk145odW4wOe8spZQerlyt4c8umEnK7EVKMJ0Ux2nWVMk/XgjNU
Jpn4TkatMr+W4yS9PlZ7Jv0yK1ZsuUWuRVMM5mXY7bcqYUT6Zg5QyG1zN96eW8tOCwQTd2qfYkBD
ujI5xF92ISGmO2/CVkeqdOPjYtk12v3uINmagfM1m+G01yrmY4gUZzHQVGwWp0ZB3MW0QyqfvARU
IMhehPh/JGA04h1/Wr+bFWt+UkHG5Qs0G4JUN6AggoT112Qzks2IHZyvB7tgGL0wWWn5d/pgmKOA
xxBv4ruc+vc4HfJ919L9/XtOdvyyVNQtqnzg/lLNvSrntXz3KJt3teiHVxjFEDiiSdvOH+u5xCfA
/xQzNbQdtoGiRT23koPczmECKrHnrKG2wfE+pOZnYp1+0Qw97OHT8qKrIA4Zu59WqtfRjbs/ZBoD
W69KWpbJiADLMHJNZUIPC8Or/ELvOJXIS5Yu9/RVsCoBgkuh0PbycHNmqAx/gYxEc/r9RFh3r6/Z
dSrUoq4xhfwrfz+9YPMW1v5ar66U1XdolgHQQSOf4QXCGUlfggXgXLRzqfexe69NTbdsKPjK6TmV
emHXP5Xqk4nJxVKr71QFkAXs1DCbhYdWbon+eftT0RRnBoEHkV4R60B74osx4Csm+Yy7gn9eePB1
HG5AzVtnQrKnrmYJF3/dTyO1Wu21hXUedSUuzgO5H1cSLUrKNz1a02ueWChX0NiU02PG23ZaB8r6
oBAF6LC7x+crm10esEQHLYQpiMAEgcTj/5QUYq6GIk7t3ReFZ0nN/PqQSnWo0YBgf9zU/isNUMaF
/5hqc9BHOzOAtPyiETI9/QgQXVgj8wXNba3X6XRCYAudtrN5h2cnuzBAUgzVftnkdO3wVXWtlnQ7
RKXPs4B8u6elayJZfFOFtGfh7XLTJGJnnR/lMxTiUmmYSphqUv4L6Gb/lg1TkRmdS4aE2CssZjBp
Q+xo5opFUsJYjKkmKIRe0qztRsJHRF+0UDmGkVVPVgpKJ5V7tdgM7tsSng6Jlh6DuOzYYoPIf2wR
LcnQeIBibP5aNSwR/EF7w1FVn4WebSm5w3UoOdwlMKZWzsy9J62RHnrvzReg0nm48jvWz0viDiyV
mxjZlJ2w4UZfpoaVlFKurM2Yxi1P0QnEHcDr6TxOFuY26G7bwYEEOPWDRaairHlpILDODxyyxh8p
hsdXWiUOsGts/Rcv7aipXEv6TxlVu5UpgcRZQv6f+1nmrqD2KZ3sytFc/+tthph8cIGsvNhMW5A3
0lqE3tUNzNQpbE9xW3koEOH0QAs1FEUR17Fwx+lkkIFRp2G5h45AZdbFKHCbJjVcn90uMplYxgiN
tK4icIwj5kNOQuT9xFOTepL2LtN9eH2EuAo77/NHUWX93KPnTdPxmZq2rWSH6NRmP6ZSooHvj6Hp
l1lLxV3z15+w7fTC4BIA8mjZCFnHnM6JRZuTlv3FRYsnsqD8WdrQ0dBFBxZZUfCTbreoZYAwsoZ4
exCawlUhACGvUQJOSMtwbZw70roCyiAa5NdOIqKiyGmuMUw09nfxun0qkqbuyrzqSwSZu2V7Qo7N
K0sqh0cv9pdkM+G4PcLNzkuFCeuym/2U0f8Tr4ZukSMCjMwa55T6xdvgDLU4yQx5YPM938xv/m9+
+8oYA/FL7NxRc2ajk93A15e3KmsOok/xmmaFRpFQr92uTBj2dlSLU2x7DPcMj4i9VGaAs18VrfGw
zDO24vvS29bqlHM3Ym0up+tgFg3/T8KC/fThN4jZIl6NDWeYcuYSg0u+D4jCJbCTB+2dch6QpFSg
WfqBlUYQ1odoW+2iVmsRcNCRfYONFM8GmxbJVY8qYXvjoMQ76vwumNY4/sep5CFeUYKi+G4chbq9
d4oWgfRbPYW/C5g+JK0hvoXbxUSyshYlCGfVgyAGEl3z3fTGx76SGOHAdLX725XsmTgbpPPo34xX
yOgGFM41YqPkNLVOtt1aZPf1GVi88fvbSHnuLDGVpSGa/S8O/w3XgetJhhE8rVKoHIB08jhHw1hc
l858nLBkHM8mvCW8hK342SmdUgfbvnw4ojynY9BaLp2JCHK7sbjXOvgExo2YMznXlwFPI6FhPTbJ
2KXq7MGcQjHrZWOVkDHshOLNiYCDrJl8xWT0itD02WDILx2WmFvonizyuZY18Q7IwnwVaB6cKHGx
HYqLZiJ6daoAW6+ZX85QV2dQK4EZfBlaZiYm7zo0pyy+rpFS6I9CxHfvTtRUhdVIdDqCJNiSXi+t
vbub+fEd1T+l5TnRXgFfiDeXGRtoVfYDjm/FtHda3dmfDCzGuPQrjj5xSsyEYXYVBs5Ag9pXAFxT
nkbF7EYCUDnZ7augxkVe/V2DEGuCfmRkDX2qY2bL5zYKberOA5Rv3yFHIpSKnE/2A/A3K3yhbcCN
DtRM2jIqF+SzTRnRcjJP10kJzVbjZEpWjIZsUssFjhJIvjmG2sNsYmB5B4NnpWE3+hbxQyQftSwK
ByS2dTHMiEQIk5mG80slFytevXEY60QpwtZZGNA2nRKLCBT+VGFCUMzlzt6OEpDlPgGbe6Qfz9ze
RE+AA9Gmrt4fJlxENiJjQZKVjqGY+i43PBBePEz9eY8p47aELEdM89uzd1ZUCFppqZAnX8YYMha1
fMN3yPQ5Xo8Z6xGX4yRu2LiglWUr/6yZ27mQRlTNxdqO/r9gaN0SeiWGCRq2EUPonPdNI1+UmRBw
0BAmUyvhjS5Sa/Tv3QAraH03por9XOOjk7CmYvIfF2wYTZ8N/+dSoWIi8Dhy0GRk+yhlVCkaOh56
MsHZVsqzBcBI720IHWH5AgMxAzpuMKxdFe++dzHgevhf+jmH6IHfUfetMYF1B8h7UoZE3jIAdMFs
INp+hkzKr4pwPnkMlJWqd3ktY7gwYdl+Pl64+N4oIgsPeSW3+zmB8dgtCorY0/XD7gwBwiS4KSwh
wTwrzfRmEf/EfDL7gVxVvwF1uIyj+ZVz73wdKKqK9gEuljc1wDNC0ihrIxCtmYrHBUAmP7wJqhiR
aGXUmpBTcNCCTHhB9E6S9ZWjP7kJMCb39T7iRU7SymSsYRyUzJhKgnckSrxm9oUcRw8Z47OciFSS
IaRCZXFCGyMmsF/cafbojAdan8Pn4Iidv6qgjORpJMeTD5mGxFm1FnRKRRe8ioVI6SelK2fFD24b
iG0rDGCokqhjyzwZJx0rTSE9BBPcDUgWW7D5HoxfY62F+OwnC3GGB/Fz/XTh/HmqUrbNLB8HfvD9
rQKSOLy586fjl7V99t1A0uTNzzF2Kkd3o/6TZZpnX8skMymdGOT1TI+pogptJD/v2iStEojYrbJO
x1pvg+KfgBYkSBtcRwXxbAL07OiXF3jg3y11Mbbxst9Y/CQtJuZheJqnRazSuScNwLatzPjXLfWU
QY9QVLYL0rYEnf2e1x/Y5VsNUduh8//n3qaLJP/8OeJkUy6FgwRwZsZ2E/NbQAJRMzntjL6BHlCa
eV0JAf3USxM/jpMs0HYvfxvgO92/Cao6Y9Bb0KOtQTgSFOHpIgBKkUCebNKpnlX0udoJifsTGYAO
6Ix9GfXdLjuji+TkoG6vUFehZSSEK3nioiJdA5DmQAr1xw+fkJWSLfUx9/b9nV1JHbPfW/hlFn/o
rpf1UnhvdUGKJm358YhZePvWifiksNE0uxbQf8U+qyDq9hGst0KvABPmIZkpi9GQ7nhK8YnvxxFk
iZQSn3jqLyyIv0d5BrA13UfGqpAUv7+P1y+Qf4Bmtky+4CwHsyjXgdQra07avyIxrUq+w3OFxEkQ
B+ZC8aFyB86O4aOem4svenXFSYRj3dJEVfCjdOER5kAciTEZ7ZYwl+uY4+wvB0De8ZjcAYnosY4A
4Gz7mqeOQ/PfDWMIWnICBuM1miTUsnVmuA7kbO7vznx6dgYlKjU9F9NC1740gTOoCp4Jfw9G0ozU
Ff4cJ1mdfpDtbKfpQm8umjd9Kmadeo/iVyR9mQcbfd+S72+MZD33oXKR7KB9AAnlAIfqfxZhMi5J
lKTaF1S6fGf44XUrve/Y3G0r41rJWS2n9ZRv9hRwTc/hVmCIQUpJC5SWtTwerJPqWIfAIH4ugvsO
B46U7orcvyNgjtocozcHLLIjx+5VD4LwFYuz0uNT7z8POdce1RbolBSoS/J1JAcpjuk4Cnz1CGhw
nfYVjkY/6r2WHmxpUaxFlmpqOOnIQIIkLGXPi/ee7Kncy6Ug6om1hvISzBhVjgId23AbVMP90Naj
azZjAqi9zYIQkS/chaZKzkLGP7qI5DUW83WkghoD3vqIVVjmee72bQtAwcwwP8g5SSpXEHWjQM3C
OF2zZt+McPZgr6IEDfimt5Z5+kwKZjVFoZwxBvBqi9FGonyyNN013LXQA56Ed1IjxN2ZukZ7XZ2w
4UPocACrpDVNFSE5gjOxJwnpd5YxrRbpiDcx5+Cx+8TNmUrKQkDRdJCzQYIN/j1uuvejxb/4UusD
4mewJjTihnHCKhiodoRzbuiKvMficyFuJVfK05Amf7fgzO9B4TxsiVY1vyP0ZLVaXfTcU66lYiF7
Z2X/+kTy7zruh/H0Xa0F69ND9+UQqEI+GJ5AYlFgpex/DFehucj6+by7vszAyGdMv0BZwan7EsnE
KfBRHcqB8LI0INyI+OfHxXBGVIIRJLtWiADy9/o921E0tdy3SN2G7C14j9MBbUTPRPA/mekBFuKe
c2h+opLwaKbRtDHmZEiTY4JAzZktQQP2L6rJ2bwI7HSzrU7fRheX1ATS79hYjfZtuI3uuLopco/k
mF8B1vsmC5IMrULGHqNwr2VsZh9MFbBdjnirnhcmCqDY7VnG1gluprXLYq8mXoXl8BvEi9LY+5dG
di2e+CuYYPdraqxj0B/yeNRiGPrJ/kMDlcShrvux393nbyCOWL842hP4dIgfN50gTSEdDDlr2KT6
/8hdJnqK5bc0J6bCD24FgGD0TAL7SD5XtfMX4S7nxeKfN1v5un2MAt/MA4xvXGc8RImlVQ4OYsLr
HZCyDqrWDcgdUXlNhhC75i81SrLY/oIp3yJxlBC5pGz2ewPydLepLu69WSRwSkzdOSKOH+2oz5dB
3EvYMXeo9ygga5ep6oK5GOpus+prkSMZt+Ej5k1AEApefhyToLZz94whS+ocmiijf5EpsCbA5joR
SPhQ3D1ItvjVKIMoB2EWOTojxpWuG3UUjtOonxnWaSWF6fAh1LchOHuTgWgJWedoHBGRYNF4SiRF
+xqYWWco+VF14GK7jTUBrdNoA6AiFVmS3JAD8+xujMVXy9JS2ntJSKTKVQp5oxO+97h5HDbWTlDF
4/A+9AmoZ5z7iKZwaBIAzmdI14NCnKAJtxYdKxCousVzzzFMxzuVzY2ZPKRBq8tzBsP3c7xovr0d
xRaworbXE3xInFwDuesSwvIOasfDG2lc7GNmb6GaqZ92foNOcEQBJYQRj9WhSaCRI7Uv4AqdnkAg
BO3P1/WbCVwFQBO5FZp709SuCVeUvrbd5S7xPm2Jp4uDIHOEExL65DFU6HGUTmPrnV35vALT0VpV
9IJCPSLUUek/hAeL29Wr6cFDv64hg21SXt8Kq+vo6lkKhn/UGzu01/vwzlaS5B64+eqAqCFLNx8/
vpmx/Xa9GegINVCcfDVdITn5aTGVxTzdt7AJu1wUYaHfvE2e+xOq4MJ4/wPIGMurWIJQ8BL2lci1
zMSYohS4SuTBKpRXHWROGkaVgqzrT51OTwZ/ceX9m2/SW9LyM6WdUr3s7eCAUgXfG27nHw5rVjOB
MV/SEgZvb1PbijbCQlJTFpezLE0ONt2j3x7cFngDJy8ggQsiUIj11YgsW6MKbvJTgacy+25PwDbB
XC2i8pXntQBFiQ7l7yRd+GwrgJD1CzfG4S0/lHH/4JjJHvI7T1R2GTSY/I15YF1oBxErwcBY2Ebx
Xbp/2yV9IUeyVpK8EKu8NqyGeZRxq8f+m0XsykAddE792gxSxqgxH6UnfhKGIQjeStzUiwIIpMOt
oZssktp+3dU2VO8uaOGviPYMWASXS7+ciSTHpXIFlQX3Jw4AlKymS03A9YTmO4jwwAvl7ECZXXO1
PQRfT3k3oZilSGgecAJESMxbwlpKx38IqgDXVyrz2Fi8fQ6Tg559cYoxd/lIXpKX/aKsuUz0IsJa
UUGlwxx04Sur9J6A/RR53RnkkCDLOeOGPCs1Tax3ISDqhRQXeR1Mc4z3zXK89glhvsHVjiwKxoAw
Hvd3T+ap5w29OWHRMsDvY8XhgrLez32teY+pLbC+QvQLJE1AkUAWukL8EfourHI9H/XProkHs5Em
69Djrelm3nD5w6gnfCvpDIIPQ6i9XBqirqTvNSjVZfgyk3jk0rTA6VXsbwA4kcFkcsDkCAlb011C
JWo+FfF7x2NkLgqysJuUfwtcn8yQvK13i8LqEWMxqB6vpklHI6eQI8eWnsfts/38ya2cJNOSbpma
+8DGHOoPVksUPSHPlkgwgTJ3KhX5WMaZ7tristswP0khAMZrtQFaCUtEVpM9bwFcoD2DvmU/XW23
6J2LI2O6Fx+SZoQ4WslSLiwDRNiV6TV6akXyDoy5FW/IVuBUrIbqXTId/czD1UBKb1lvJGH3QnfA
+jzvJ7NJmIooGQGes05KExS4MykHw6F1yNEqW6DVAcfHGnRDcQ+eQ+AiKvozNcBv79UIUWwRZa1A
b6RC0su3Lku1DrUmaZz78rtVtQJ5NSVTrSfmSkfVhQOFCg4GjIam9sjNIde5LY+W5ZrzMJQTUUNC
A5X5CTc33zhUCjK6ehhexCcAS0BG1vUbP3BvTdkec7mw2gtRzWWKfs0drfixdKguZ1pFv4DZ4nKy
EpcbF7uPYrZFyXzZuz52sDLEiES4UcyFdmWE8yUB/Xucd8f9LRBatXGzpq02H8aynSH/nn3U6Vm/
uE/Fdg4eqZEX/EnSXPVtM4SklR+ICMyio4kiEJdSOaK2ORZHculbcvNn4sAKw3h0B8pZazDSK9Ly
hSsF95tCEOBdFdNeSNUhq3+dMyubBFRIqUXmA6WekiLIYCEiJbQApa7/i/UvWrUn6se/b6SmRWmF
eC8bHT1DmxtFqvU5lyMSdRHZXn+0vw2YPJyKiHRoPamiY721cY13SjpZaPCdHSLUmxxsy6YUT/L/
2BUCAOtYGeSQCTbi3EJZEq+fdlNQ4qkl2Wo+WKd7tPyU/6Xm9gSMOM+qTCZi0bZc8YKhWXX0W00J
WlQNBjNcQ18pbZ5H+2OKyE8chfNj7qvrLWJhtZa6QLznp2o1+wPUwee49DcPgTpS6D7DIsxOMURT
I9vy8ruGFKxH7AQ6bB6aqfnD3vSIwlTvtcUAm1H20UW1aMeoDFJLcx7uQq0or3wKsA2DJ90emNJ3
vAJahNtdb+DBoMUCRB1GR9qBO7JYMZ2CAVlNgqElO1nAUyYdwkZzMKvZFKf2u0I51uJdm+te5e2G
WlOGW+C3XYpssgpNCQtfVF9s4BdbEoccNbP/TT0BYOFUG+MhZ5Sh/TZDW8hpFVJevbrfyFYqHobd
+CvJlDvd4Z7WA8EbVTmhfFQaHcP1XjrREyTWdKemssOpVyNFmfrx9M9tI6dfdL46AxRJKaeozukr
jlyK/9/fNwSqldYUdOn4maOt5ng5ouWv6+s4DYU7dzYeUZtzDDrOrTGWkwvzTAn/H/djTxwDNO5h
bBzJD+EjDkPY7hDUU+m/iQTuzfxxyQn2ehOo3BgkHyoKtWth5g9zNyYa9p72J/I6HkUQki3OVlG3
pglLJ/RtuEYSvw8M5PtmdRE6Gz1YEyepjtBJK3cCtAfMl2bKX2D+XZWTac9mOPXYuUfBe1/KVj/t
IiJrFawsC0zcIMIZGTtor4PNif4wojZ9Pt/ykmI5zBgBz1MX+I8zp0oFmUrDZs3Ps1JHrY5JJcW7
Fn5VXp+Ehq4OCMDmKQMbyjho48BEwNw3eWEqSbeVDahOWANdmKBpcPF1Ys5IA2p9/ZJlyLUwThyG
JnXss2AgtNnNfVsQrlXZ939tGNbgmxvXI04SF7NMAyES/fZQ8dlDUZ/mZx+gnBAcUVjcbzmBM2IW
egXiOJywqHPhMXBb99ylz+46vNVJ0wzSp49sUL6oZckUGpmd4C5tV/+2AGPG5q9y5bopTrEihP6N
/ANXOTEpJ7fFvKNzWYypd1QoYA+sxu51+8Kf+ETiZoDbnxQkZFS96yyPVxFM0oNM3bBwubgXPBNa
CyOnViCGLo5uFQmGURXPxriWKj0AkYHwO9+BDX60CVGEh04rJ8jk7OJAOz/ExFJ3DvKAII0+SU62
sZrsGdb38opWqQjLZhZDFnOiJtjPGmZG/bpSgUrZox+/RdRDVraPrn3XZl0sieNzdVlLTLhfQ73N
8YplruNt5vQFrjCvLyGzB3WyvTqr5HMmdMDc1Q+e3Ka4mYD421AdI5/uMpefluzWekd2hXtw26Pk
BtvvioG26IA2a9iJMEW7N44XA1Zn7PH0xee3PWe1r/Mdz3wG6qqutX/SLcoPa0n4nKbZEn924H5J
qsT6bASKZiyAejnQRBI/Pztgt7lrOZk8uH6/rw8FH0AdztdzeG9ar7gWt3MCWWZQqUNbRybZNPnT
V+GxfKc9ToJODfmm+iLhIehRYNAu8p0tDRuDCpq2Y3B4jurqUXvXt/lusidJtzBzGt3W+gXFGIy3
oNc9fYabKdKeF+tTVPDvhEUf+f045dFZJ8ICe5y+f3i3Rk/gCLUyad+YLt0XmgCHSLtXq4yuM9Jd
2/ZJT6cvr2++UKVw/uqqNhbrgqxW+BDoKWUvPkmAGsXmTo3KTUfwaKFJ0c4tDkcXuvQjAwwVi6i7
bHw7uKvUgJk2uq1TcxC1OC1EPjn1liEzC8sqIgjrybW3lVmAuw1N/yfdeAelDLjwfl3LaKaANYF3
ZcOv4vMM+D/SXhoQ77dN4Qs5YIKkhLFAMmKJ/wL7wX/IEhkYWy33Jgor5qz2z9gIl5cmSFvmlSgj
e3sMj/rl9g7tBYuh0+cXLm1MC1ltM9iMC9qoEn+kCpMnml+72fUVL8jrqaes1G0JgLdBStSRdXCL
yV1IklJDzEIiHgiCX2NCcaP5VMbxifm81iacEG27HEjwaaGft6gq9qMbtxSbFY5dZuZ4Np6Z3zDS
sH7soJTpPvgPagS9ecsQvHLRCovHEYw73M2O0USaK/cKMTcA6Kqf55TPoll6/rV0SuhP+feuYuqS
4PwiK5g8tgWZ/4msufoqfZSAdebnG61at86bdoYoizcl6ph9FIRo45FPMIEUmiFzci9IepJq/iP2
l5RlQXibIBhyGuGFNrZPlwPQnsfg0gv+VglS233w7bWBdUV2W44Ly5Pn5uR5IsomQD9XZjArevGZ
o6cxNsO+s7OnVS0T2IYt7hu9HqgTXBi46Dp0pcD9uEjlX4JJcQ91jHiUiPkAxDoHpg1jX6S30UGh
xrrn3iZ9dKO6aOteTx3/NMP8kNGq/KBuiC22s6ai+mkY8jr7ddLMS7mPQfa8rypTxzMXig1AaHhy
8QU5ag+xN8OFZXc0ANWo7ahVF6E19yDCB4NudAuUVW6EESJImlxcaVOQv/i0uxasJGtZI2J6PW22
NFYZOD+QMYEXoXcDPX2ACEJYsI6J/WcvVUFynfPkWrTk+AVBFhKDhfjEisOKgTgcX+uR3IOMWjwQ
XB2vglzRnM44tFVN4kG+Cyltch4rtChpa769HWPt8nnZam2WgUMYIq1/ga0pr+3ICbw6cs58UiVY
DYKbagAZxJGSi2bZvyF6l3mIJA92vejYN9bP+1hS8hsZpZtni0Z7RB19pEwaXDQhJ1Z6+GI4qD3E
wRqg4AUydfw1xorQJKRZDC/7o+x7CfrlkFM1jb62U+r843TP55iDsq+Xd3wdWHVrglQgSgd+vaqJ
OuoyRlUGT0jZkvS5xdp3CMdEDNPAMPuKhC1uhcW5JchMCuY0Y1QwFQ13+QPmX5cfRWRcO9uNjUN4
RK8zMe+lLNqOcx6Yh2y/pSn/8sazlIJ6EeraTGlwG2LA3WdMiU/yhGs3YbIjJio200MQkoI3E+8e
UYC4LWOpS8jTAPT4CIMg3np4C6fC4sQrp8vzqlipq7YNXOZTH4refhNQRUPc8BsyudPjHohqxYMx
881kYn1OFPlkClJf5NXFRqPGD6Ce3Oh0Ym1zmBhAF9KFzSBqIdgbTm3lWtePFDZ6+TEdePAf1lkS
qSMtQxJaNbxc2eu7WUc6e1Ili12I+wRNbX9sPozFpYstLYapx0tRWPgc18nmFY02TpWc0fmMvEXK
Y6drSx4yx1Se4683FejPb8NspM8kF7W/7nNevWhGyVGgk9BdKA/IqmXS3fOMNSg3RPY7YdYgvG1h
wsxN23/cQYZxi+l4yNgD4Gi7Gq7oB2Bn8kazWCgS16QsQOSggz1TaUw1AZYdhBKkuNqijR1JxWCw
CUnKSs4N3Npsoai7M7gj210hZA7qNcVpxuz/wnjLM8HsLHNQApKzgx6QNKGJwuew8kYBXP7D1hAF
Rq+sIVG3tH0pvggFaoaOAQngWBATexxlV89NuWAoLYFpyJLGU4qPIM4uJanHOFmCZ3mcn/CIxM50
koNz631TCOCVYZMgndlm95USOvlLsT/uqSoMOk1csPmVllmMuQAAZjzIMFuHpQvDK/J+kmeepAY9
XKuJBCpumJMFmDBCNTjuwakkPazh3WhT3nsUU3J5h1ldAdnq/s/uMSJ/k3gjGZcfk5hIvPEI350P
yCoJdc0Y592OJ3DYD5yqzOSUd0e7ClqVeVlg+0usiYsPpOY16GpvBCejvEp/O4eoSeLGYycs3Kus
hNEQiSNxHEbKuhnomNreLKdLVHPcVawjsGdW781OrVvmuySAFKs5qP365reGBDAY1GSgABnOaNaD
9MxfsEYBFdKCRgtAREiHj5Ipy873vEz4VS7ggwtNZ/A3Ihv+SEJuqf2cHCL3y+MY1Sf0oGReRDn+
AmXvi47KuuBKPd/a/SOAPx8XKgpBU1bhQf0xv02wOlpaxGsoQu3a+F6bkroDWxul59S25wASzGYj
ROxVbkMI8yJodAiUZ1+9yj1m7agcF5zVcdatUga+1JabdI5JBTZvbgbybbTeZ7xQmUig8eDYZAiu
ieVZ83tnWaDPCuDelmvO+WOy6bQTInBHwCl8ni5x7Za9zDXTs9e/NG87oIz8L8eawyUoVICn8zmK
qaHinkA0GNAf8/QrQcb8v9RFzBNeX9p0gtcWemGbj74JSHA6KOu+gSHN77rv2NVCUdqSqQOOjiK/
KwVLarhWef6vYGV3KC6Rt+zTTvw6sK/0yKzg8KPs2oWRhoTcjQ7P+vbnFlNdAfUzRiPx9gE+Ysy/
6unuIRocI/y2FPakwrOEr0z5W1N+xCb9FokDgkQs0XsdcVLa1tU3qb3naw7eM/FpA4ODyZbKfYaG
2kbMhlepTiOiFjKdhmNLZ/3UTWQwqG40O374FKhQ4Yd3EzHVxwIxEb6IxmzZTcbvTQyjQ1mK8a09
Y9J0EmQMHqYqhpwvKBuDlZImgt7SmCgkKM8kdpNpoypgcJwi3ebGwmnIUNpOPS27+q/uoPi5btCT
rEGnOl7EIQWK/j/9BOR94Ew5FLoRd66gNgnOg2xv8n3iSN2C8SyItCLgAW335fnQVad1LvMwdVVV
pl2dA2yLDjRJlQknJkw7ElM0UFcYLmAefmsex+Md05oBFSWT1F8hOVZKxeO/Aua3JhAqIMWdfHTe
TYEm889bL6cegFAqrHtui25/mm0rAs9fwWqO1hjzTPydcP4ltJOjBCuELMN21MeQI6LG8AcU7Fjz
tpRv+VjyGNVmNs1nqs153bQ4Xqm+Wbm52mHfhD+098uqG7Plfq/qZbfXXoGHO0VYrPYcaMWGYRxP
ALP008kTNOYx9OjRn76fI2pomG6YmrrlSfvxNv+j0ZA9QmvzMKHM+AU5kSmcf+pTWfJbCeEGUX0n
hYphk4QXe5lwl8oyYuAG0ty70Q5mvpmL31ixFG423qSf3DqqO3xDt12xg6fg8FJmR8Fa/Y9hJXNr
fvzpstuiXoTI8Vj+pjoxrgoAtUfgxnll2DkLpVLXCoSnb7pMEF8Xkq6JFu4TPYE2saAA8C40EAFV
+5w4OYHKXeOErzW24W+0u+SneT6QmmhZkBpkIbd5xUWfpUrHFhIdg6/yOy/MGcWBMk0M4+SOOCbx
gn8EsOTbX5FQuQKVZHqk3vVofAC77T59XNv2BvKoFdy2plqnaN65T07AxLjbIzMHYk4cpujQ8Exq
6XIAmItVLystYS0Cs9fqVMcCjMlHrsLuPr0/s5D4ikpw9zQY8r8yBfWADyA4hUrDB3Mhn8ItkRS8
oBz8b4zFK2xX+SdR2KCJAzDXnG9ldNWmSYFE1JuW0vLH2JkxQeXWYVy+tJr7VHOqbtNXOu9OWuad
N+UI84vgVfzAc0dE1x86az4/OiGVCsn0UduGxsXk+D8Zlv+PqOzOfxptX0QR9sduiWFd9cfvkeTp
zZ1OHFok9d1XadFr8Rdy0W68G/V4Q0FtctiC4KWbc5ruu6Wm9SedInJdgk6SLnJWYndLyv1QsZpT
P8sHcF0Ct5tbOqVQr4MYA+ImBbgIQMwUV0CH91//PsD1wcCNxLxzzjKWmRpf7PMCfs5gkVtdP2V9
cfcnRhqOgfxMtc4dD2AOOGf7oh3/oMNWD9gPHaBWzKri1cL4v30h0nFrAU55qdb7JYMi992otxYf
f2q5ewQ1xqYXESJO5q1lA0xN812hPoC3pAY4qRoZVwFCRCD0M3Unt1yT6d8rQ0pJXvq42i3hQ0j5
7IcyX5EvUPVMpivjEPXPrpC26uUOSAfza+dvb3lINSO0DZqJdm9AAEEe6JPFW2AU6571dYLk75FY
t7h/kn3BNpTbY9nSEfbbedZA2Y5M//3VXZI9cR5skclDmih+vtR3pIOyTXVA0yqPvaoT+epwmYy/
CxAtHN5n7BOYRSCvpSoQCqonwIR3oAja9gc5cs5sZiW016s79BFpcKhkJ7Q0PxN/WAlZ+VkSDPui
/49+JgsuKR4xVrQ1R5BIe71igXdNOsR7MQmn+zQ6g9+RDf4rWtTQOMmagKyhyfrpSC/IBjLdJPDH
Mdk9tygaUx6c7NNjViiE0lTyA+ZZZtRt7HoF7C7uc3sGEtBdanwSgWBu0tK8DO3KzhswByEtMro2
JlvIqJSalCeJUk28A+iF+4bWsfdvAmjE9TNCZvEoVep+Z6wnAyVegNzN7esfGtR0RX6Jrn3LmYyF
Tgflr5Sm/vBqGtJ2fhxUDwU6kKnBK8+tQP/LBWVzwmiSccFlTt+JnLB3VVgpkG6gO1RHnht6s37b
lUuLE8IduE+kCb+xcmP3licQ5ZJrT8TfsK3+NEtbP8Vxb0qqUnV0gk7qeu1IR6h2pOa3GgV3AO5U
Izq2WFMpvhHey1aAWyQDrQOYKDOp5dxmszP9X9hwKhXogycQbqx+fpyxBYSWc4eB26VNiXDlTN9K
nvHbEJR1vT6TwXA8B9QUNo73FPocH3pBeFvFWF4cWybCN/yy22YE/La5RaflXdyR5bxYEhpCatDn
RKuY0GE1h0M5Lfumq055zsdg1k6cGwlLcwrFoEOs7cQuyWFWABSz21YYUPdZI/WXRaFmXCgkk9k1
8209YyrlQHkbRk7KwgN+ZkJ2wwbwpcsrydIOwZrdlh2a9BWsIgayTwr1d9p1pgZBTBJM5//bD4/Q
M+Sg2bmPoC2Wc6bIOrG35RFhTekkH0njesTGpn5o1WT3yntwdrNj5b0LpK4nYBaSqJhchTQ2ffbn
pogni53nZh50UpgqqLXyg/Vfryy9gll9KUeBR1hktalASFuJKrFfT/zibRrRuu7cLDUzpmTg3F3A
lSw1CgTogfoAcp1Mo78ai1UgPr9Xp4woHSQDecUTkkxhvoakBvLq+kYyl3e0Np3+MZ280zjHojun
ySohPw22nm/g8XcApSqfVoDoRynnSD4p/K55/Vc+nL0WNJi9OLeuJd1GzRrSN7+Sqor210e5FLdb
9J7N8Cem3MVNVt+jLNjxmVhcz23eA3HWS//fBI7gbz1PXs663r9j65ZWqups1BFqKP9WKkiaKaka
h1uFRE1KueT1ItUd9mp+Nt62uxx+ZQALN5eYjTVCzzdjHon6jvnkbSoVOfHzpYDOjvHCjJG96tDi
Wo8F7D9r9UpcZYEi2wA6bXJ+8MQatirjlyZtTcUg/PSF5Q5AJdr7rfuPNOJCPBKQzwzOvOK1iOP5
VmVjCjrWdeLtRIBF6Oyw+rDmnOYLc7K0jAybA+X59udyVlyBCmyf2EB4rkXQttaQTbfbMu5TFpR4
lIhsxjNWKDZnNtVFjy9SuCwNo0MrUW9wSUr8mYFjOMhVvrt/s+2Fu6Rs7eX2od3w4s8TYwM2YjHE
6OIh51TmvIKdRkjNbYKLXQpiNXgv1OJIYWEQ4onZRq8Upk1zS41c2J9kKvS1AiplUP2bPxEzWsD5
uyyQtB+vIdEg86y692XSkRr/hmj5XivxJlapn0jRKeEuktRa2QYNRbHyXIRo0EUuPs7ISx3j6HTT
LW3m/2DyTLNImE8jfxg8U4sQ4e744XwEONI1bOfV9XCpbTsNbGhmSwA+h/b77ahnysA87B9TSff6
CE5QL4+ylzcAoCNNzkMcPNtcHWUOu8t6Dd6oaeP+8ERB5OuRZaXMI0Y8emwGAsx9tX2b79yoYuLq
RzONNj1JfSp+6ZyxRXtO/AbSf5mdSX6t/be10gVhP0xN2X9MEKVZSQ5dkXMAeZILLDosZnljTPXx
imejLLALUNNDUHic+DfPTEV6YzVfb04UWgQRwlAZD+VRgZRe0ArMjw9gIUxo4oaIubPXOwICFScs
fwVT5AuRRS4jt3ceqrPNfhEQvFPAyNGvDVwtbC5HH7uQjsGjdNniC4KYVQxOWUTvnUIs4OfRI6Cn
rpzAiNJIDl2s3uL2di5IvEYIdK0MpB3iSU/5qwAErTc+7A8P7YNUCUta78/1QE8kXe6gTL6ydMoI
fC/mXhiFbKIQQ9lDkYF9DlFkDuvr0AW6T2uIoE/778gZbh4kwDnRerZzXnJAGAxh/1vrbRq3w4CV
TNYYFH9X1ppqNMR8H/Rcnq9welPA0T4or65fIgsvOn9LgiqexTSuAsMatqr86cwhMnEZcGalkFJT
Rkzb6jiBUkrw+ZfptlKrPq40a0PH/DooR1taG0Zuto6NkWNf9zJCnKpQQmdSWQ2VHgaCqNbJLJOH
QF1EJ9LwBGxKEQv9JGZCvUC6lm0hmjAD0CV/kn588pzFOl7H1z9BrKc32RRnncMoR9dbPaOQ+Euf
5ey8m5TKFWO5xamFccGW2nDvknxT0ovQbLOLsX4KlChsP4C/9H4gmGXUwNwCZeFudld/tGmwIhAB
6YALrxZmjty9KEt237OyGcpB1IrJegAF4XLOb4RQfv52C3auXdytTzDkuYagd+WIg+/MC2CElQJb
6TPSh0DBkMNufclxCDcdOgHzsfYgn/1jvZIPGlKw7SaptEd23+4InQz8ExDamAF4CDgEJhkpxnis
XYS3y6Un7KfGfCOX8/xy1Q9/MBig7yOp3TeEw1FGZ5T34N9KBPXdDdqDCmFRLbdBtl+dp4GneNsy
N835nB3wbO9octt907UxwnTwLMH8yHuMSD17YKI3b+xt20kmx0ByxsnU+TTsNtINZX2f4IpfOajQ
zr6cKFGuuQ+14lm265QJj5xGk6SavpsHMDg6VrK31aUD6ZHiXx8cj+7PepGFFpM7FgC8/fQKm+Wg
/mwPERAMFpZgSM92XzmTNtEkwjOEUn7O9/4cFcVvKHcx0BGyWKGE2I3QZQ0OGaZJv/An9WKMpNG+
bO5nj7mQ1UZrsMF41U/A8jdKFI0QUG6nHz0dNI4nClR1DyYMl7viabDsp/v3M1cnrIkWM7S39SD7
upuyghYkKg8QiKcCqyrU6FYHo54V4Fhlr3Dl+ps3TWWa109NsePf7CJXbkynyam6n2d4z2dtT78w
VQuizvSD0YZf0zuW+SsSEstWgzfB1wQJX+737inE4+IfVyJle56e4nLQRoU0VIwrlSHGerQu1oD3
VGGhfIn5PW3ejvtnbagEvzhOMaD+LKBMogdnsNxUDOtZI3ivVdXpYwtHF+uumZgG1GfACD4tzOgU
O9PaiLRHIGcoSG0xvvOnrFeGljVBzHIB0KnvfRxukLHX/khIDm615nal5sGzDAFLNrv3vxXJYHVj
MkdDAZvYZSpy0FhWmj/5bjXOB9j9AYA/Dab/60N3rx4Yx3eLTUH8LY6xwcpVlH8YOm+lDizL8axM
OxmdGNnE8KI/ixuWp6B/kGlu91bh0eTvy9T1NX+Ae5Z5RZ88YOL72ufnVd6O/bGLiQCBilpnaPle
GjDGfv1QR2CW3Ht41OfE1Xu0QvOdiizcLHAIBlG3ARmMyvcqLzaE+tHyfR+aYvFY5jiPgT74Ej2d
LHq+li41q9h9IFiozpzCkg+gdVnpp8X1h545c4hPREGLttOZxeHfW5GDqQDO4pZJfix3tYAkA/Oe
jl6eDMED/2gCYSBdzLcmMKlk8qKCoLWfoyevvYdUEgwExe9qIGdP6daAf6y1QAJAID8+i6H8qZH5
rgUr9PTMMRWEujfHqAlFsz1RzCGGtJqYI1xwHMjwKP3yyUHUBU1nAuI2d9hOAEB0Ic7jmyZNfXf8
00jgM1UqWlPTGQyFuPDEmPXwoH/Qi1YxoEVdMlJeXV8dP/cyUVKSh/jWsyKksbZtDIdd6qeC8eNN
YJ8L3xXCDjtZAHeR87s10BD/2bHjxVJQwzwzIGyKcgY19R9TkCvRq2JTNpXooqY57S6lCWpiWrWT
/Xe7gQoyOEMWdO9+bcGfuLGyy++awCRC5naUMdyOEYrWKGJ8Px1MAtS1v2QccmXWOmsPqmE2jWff
W4Zg4wiIkJACEGfBU3oyQnfd+jLmbLdSiCmt539qT76yofrWus0jE6jo7ONCjZYVoxHjN5ExE5j5
iOqWrvmdxfZVZMMAB9K+jCZ3jQi8xu5ONS+V02p9EPpNdY8XGJZ8PswXc+WTD8EsUaeG97YwIRJp
nVBuqds33xUvuYPdbsd+RRUp0ASaezDA+GfJhK7EH7beDfN8LkZILJ9IXl7owfqS4W15KwL+/1KC
VYM5PRmjLYoQ+nJiDUR8hdOifcTTwWPmBoaBQAL8nsx7zYDxzioOAmrwdM8ZKglNiKYmj+JWJc4w
hygDNF+RBLPb5zz8ptNA7zaaU+EuEhgvz75Aozqq4VgaW7wxRDFdAZoeNwQmX72v5TiJSrcmtdr8
hTxMN79zXTP7AkQd8kXyluOhVzSDyIn+j12xxf5+EFjfQgdlbhpLnGvuWqXUbfLDMQY8XQbmzIQB
OC1f+yjfeXyIIxd5Bhu3N57CMdKPby+ArA9ON/OCHEj3Ohp87CBWblOD8bUS4IiqA1kYZ49By8Vm
1x0DMA/pkIA09FU0jDk9YAwjxhYRzWiDIRB/Tc+clgPu22hwA3Dyx8GznlBR20SKjwkGQx+DrYDC
fQUXDEzqLstQDF5X6LTNN25iIi5Z6HQ7N3WkzEcAldn73KYsWgj+5E02cpfi0QG1hS+LQ14K7ah7
FAOiVUJWLZem7JSOmXwelVN7BFuGdJeLWURZYca2k8nMLIHZssLhFJ3gi1WUOv2HZjGbVaS6oi6G
NcvoFYjVcOHUxROKeuMUNfWQjcaorSDkEFzoXby0G60KkQMAlwTPqgdoO+lPBSHxX8gnIv7nQA7+
1bh2kiUaB+xuygMbrwe9vPoOx7EIK3Kv2bbdtpVr6lWMlkZJ6fqVKH7K5JV9GqQyNlKIzQK4546o
QwavTHaz586rLypijxbechhdpVDLzXU0GBSA4uvqRr2jZ8zXYJBmyYmpqbeVHcfQTmRXAlovs5Xt
3vXsEgQv+v9v186m1B9i8ovnF26iyTK0wamLsySXp7E4KpCkAYBo1UsLutDmlY/3Ctri3cWUsDue
9t3oHCadGM5RDZbYgEW9caWmfIgsN6WueAHVZWue7AT/0Q8J4KHRuBsh3BwKSFH8/t0sPrpkhLLQ
zHldOBjoZcZ0ih9j3ZH3hG4P3AlWzOGjMVLJ1j3/wVQxHGI6Rs+K4+EXp/nfL6MTC48mBjKMYwki
7EFiPxfoS6st+LnhtprNfhkRUFnUahjR87EVcfqW9zm5gTrFJQjoWsoNiVohQhsJrMNWlAQ3+LZU
amw7Af2cCO3o8CDlwElXr5tg8c5rdWQX51CrcWyVRD0LXO+7OPRdZ3ycnRqkG3GckERtr9KMqCmi
3Uoa4af5n+LJw5EFq5WAvKpdncou+tyBp0OnV7/zrrQ+43KOIWasmeAaoXNYgxthWS+JSbQUARqr
ySSoI0cWN/Io4WzimYg1sOdkncp50fn2pYBXEoc8SgJinRTsQ+mUqzM8Cc3HdYf6BjIZ6mLPF+kr
1ggrtUkzLK9vC0kMKzi5rGNllHgInw0LG1bRgdv3+8VpL4GvNKYYWdF0NkHWEiNVPoq0wx8UmsHQ
K+qyQYSZFhyaVukyQWnlWRU/O7z02QPrUbn7iDriuKfFw3918d+UQ6eSCXcDPd1Ey8e1AY9ocFYK
vZCNnBfHPBoIyVCDYAFJeTbfJB81yPJT1XDVt5KYgEFmNiAkq2YvlXL8BE2n6nJl5KTKvpETmjDO
HPGyWt+0d+nAlfkxiEIPAdlSMahc/pgwFPZSyA8Oj1jBqpXzKq3rz9CS+xMwTVRsiybeRrhKKEE3
WYNBVG/met4iilyJ98mL1odhlCTX8DRyqyvSVWIUmNR0kLxPx14ObyGAe8O+QRLW2xfsLgl1NKSC
6bxoahsmXbgUyLADbm33Nuqhd+ijkZIB6KaCwhQ4Vl5kEfpmnQr/Ygx1LvfQVmPwU24qWqNyWxvi
q0i1o5dQy1BBDhhgULpF3RKfsnbhX1PjcPinviIwofRP+Y+u/2QL41QSfRpD0htBYIPsFrM51vHY
Zp8wfDEGmS7qa1cmTfkYre/UWGd+MSzhmntBHYvxmZvqiNS9V238SgSBKNO1ozXLiMi6bGY44hW0
IYMqq7eucEJ4tu8hyTzInWKWQv03TdQna9WFAo8rYKIp4tqgpRz9CP8EM/8QtYHxP4+RYCUizvWJ
1vn/cbYvDfGU+zBwtynMjYs7OAqOQaMVH42nkLQr7AVhN5HfTSJpKDrs6Dbl4nrcn6k8IoklawYU
7Gc9FxFlJ8D9qA0mNTD4RiJvMAbmNJRrI7uKupc2wBmKwHaMp9PGVPIewPi5yXnDtg5Ef1yyeQcn
4zj2X01VVaXhPe/pumnHlbJ+yooTb2YwJHZd3O/M4W9Ppp08KxzceG/j5cEzpwc/zj0uYVrxgzRK
pJhZ6NSEnRNZLs6hItrl4XxhTUQdXIUcqAhq38FZrfggPPHr8migRJIm/pPJvzlFQMLwb19p4Jrt
FAzDVA+T1xI7gV4M0f6lgsIYS0iwbqKM8KkxWieRRCKNKsth7WdITGCXGpCNw1zTv+rJ6eaLkDIW
doTGwzP2OiaJ03BjLEGI7BqOMYGeOeurR0NqaPi6VzY+nRtbqBR+1aRASX3ysfsZVSt+Z0kNZsxO
Caa+Zh30AVdGKAaajGjhm41Ie26fD/y3y6yUPUlJ5n1kwpuN7/Q42Z90Fxwzl63/k2Z83m6kTd4j
bdJPpujQCFnaNL8FyJPehMJ5NmLeYBElNieCe4VwCFT+O+DlxBEh+xEnMb7G3D1SxK76BOXBdxNe
cW4sm8gc2tnyi7WMzhsxa5lkQN3DMPCQLgEcAzzEmEjVGh0y5gkLQokhh4XBzrXoCfsN3jOPzHx8
6qVpWD/4l0raDzImmFHRmq5bfs0CqND+emAFM3DG50ARHXTaKNQcbw6RIH8NqclwddH4b2OBBci6
QXrhePSb0KK+jCC3WrUdtCGCYDKnKXrDrOREmTq8Lr2BTTzqDY4N9Y2licb6k+Hb3jDiC8sRfF31
HSJgwPsg3u3cmaEOXtkVT72sdMT8pSY7x1kMBYm//qSqUXPovT/wLXB+h2dezl85P5pffvuP2fwS
GkSxD6i0kBbVwccEUhvcwRZJZmWGDtpavvgOeLEHNMLT0+y75edENofXOTIFR0s0NAIMHkS90aCi
nb1wlBpcp9Jml/A7bDUkm9QvCZ8x1H6CPve2+TNRM8uuAIkH+KENoyb/eEG1pYH6w0Ks3MP1+V/I
T4g17WpyIK+weRiVmuR4QkfUIaVVXxvXrMmm+pGN9I41v3LaXtnEm0JOjn+X943TR/7h5uOditUa
NTQkpOiAcgNehxGUlHP1H2aLHlsXQLA2KWF0NpzIYGYEiLHc6w3pEBnmtymMuFxZVGZ96Pl0X5FT
c/IKxsOw7LPmI/WWhdcNY7BhJvfjQPnGwsvOGl8r0T0YJRgrG/fp4hwPmtPaZQnUlDXoc4VTdhkP
kjB9seVy67UCAdAaxgqYZxm12t8EaB2GnOoayqI5w9azWack73xt23tSLcFiTJ6HFZNQWO4JncvJ
m55h+XNMsIEw5rLZyiTwnReWQOAKysEwC8ZlsUEe9td8lkKeoWstNhkiPtP4EYtcrqV5xpy8aRv5
+7GfzfCqPTZ6EJ9Lnw6GNDgCNgw8bukdGwPChvxm8g+c8EoFOFqgEFia6ybsZyEJVNAFg7YZPh+F
9n0e9hZXEQU8t96yf/khCVJb3UinNLV+rAHGYZWXLjccsNEoLDnJ2BdbKlUVYGMUFgyWB9n16xmH
0n7U+JD5dFZrJudAdFMBB8ZR907zXpHVLRmUGfXUzppt42GhKdWKWp+6jY8FYtgvMTchB6756imH
2IGoek1KjRyZnpE9rNEgCtszrSF9cZJqXnW6kS7C1zNp2cfwrE1pitvOxqNhhFKc0UoQ+29Gs0vm
v2qu9InlncTuyHdluJXoj4lj1+w+P0rJ9FXiN9c7E1JW6ZX2jUf9by/okWN9v8JO6oqC9z5m0tn5
Wq9Yw4w5oNMNarGkAauEAU3Lx9wDFMz2yXtlCjAHmb8qZs71AFZhF3a+k7uHUpYmALVweVsYK02Z
+vvB8xaHUg795y+zBAZdvhXfLaQ5j1HjJRiuZCLp5XLRrcBrV0mPalY3aLkYtwLeJNvAlpnaZxf0
zvHv88OmnlyiXBgg/d8lOcNmOtC6HoWqyJc8Qy7ksQK/foMiqQ8qWDVFR4Oc7i5Qvf39M1iGFp/G
MfCyRGhJJSn7wuuO8MLdN+Xzoe8B9PnIF/w1U5i2lYWstNydtd7ufHR7tqPN1ph1h285HgYluYdh
rkCkdCBAmFjaKkVgqBMXmCfjpS/ghiwQKC4aWBuTaDzkxJXJXCYoe65ig6PiTwbccwCeaeifa7rp
0DNVFa3/pPu4hDNmOUpLmq31TNzTKwQJijU4Ccpvnj7YLstZIkOK2XYZt1/h6xjayI1toPHRNf7v
b5uOqIE1rp1FqrgnqFpSDlYfm3R7+Xe58qSe04UKl3mPcDS75uIzYa7z5fLor+rJo9wXd5Hq7Gio
V62/Igdx7Asy9baal52c2uerVXQAloMYeOjdupyshz06DPdi55yxbMXFunaEw0mphbItwLRH6IRL
9XBX1nYLKgvZGQQiRcOJtvrBH5GLa94cy0GemHAFpDO4BoRibvDKnQkDC/bk7pAXJjwCIr6h7g0c
BL4t8BMByASExGt+pej/VtmBBBosco96XWAcmIeZgftJZkfs+3Tcjd5KpqyQVLBlOYgpOn25AP6R
NjWiUqfc0zRai8uxwJusGrHhE1MhAvimwON8xaAtwvZjLJYyTvAygFKoQUod/8P2L+2zQgFfoiM1
YeWda4qskyBi3XxbOmLmbIkUr0Ac5/1lVTgK9FLwuP+Beaj3MXGNG9Kt3qC6x8LtY5VooIukt97/
YdYi34qUt97azFigFVg74mev5G7rrtqQYHxGVi80VQM0iWGbJOLVLtXUEog2me2kBDZvxl8uHGw5
n952Amft3YUOTlW1GK+G3Iasb9wgNCLLYNEHlTvDc8vlHd5GSpBZLXFqrsEQtRiozJjYgSwalXcy
tXZFEdN86dZAkAkOXWnS64qYLaa6PxLKIceCRIyUxj2efgbGOC9s8OA9It/AENnlGWC1Yb6064DS
iqXzFbPEr1F3phcDHztqea68FQ2g8L7aK3IstLKL341zEs9zRK8ncbpVVfejNyBwZSNeU5379NqV
UAvx2k62vE1MlcLM7PgHQJYmaYg9wJUBiUYguPfpUAk9mNTZVP9UULn7tuRKg37Y+3MUNR1yBeQC
wxxcWm4Nb4RwrPyn230u4JTrQfnsilq1JT3r+jeoc8WJgDqlPGA9WWuQqdXz11Nzup6dGnLKVaDp
feexbF640QysHJhNGrUPgUxbITm2/1xWOP4Sg0pI866nDP963dFS28dKC7JfZHaBOkzrAqmm5gD+
bcYbyL3oGePUufFKBsAgw+DvF2DOEciUIP3Vli3Rv0GuBi9NRcYQPTVgxwRVg+Mcb/876Rn7fHdF
JFaBg7aAkOO3p1JwDXECh1To3xK9ShlqLsrzPEOJSqbcH2hzAChB0kljDmYwGj5W/rRBBtEGjKfW
BynDeMvbvadnponUP/BobZ2o9SSdtVfbmTRzn7Ol5yh2WpPbAmm7LnnF5K78wno7jCwr2BBmefC4
EtPyQ6FV3/Hs6zuxY5rmICVEAyCzse2IHfq9sh0kZlNWMY+ck13uoiDlu4lDYpf2JbkqXjlmw8w+
Aei3k/X6RWYFr0NPoNBhPSeb8i2YNIEOHqS1gCOh4N4e/CyDGpoV0ztfUVmB+VONV2nXDVeEONBS
J+b19h8BrwxiUS/SobIuslG4caH0f0GNSlhnYB4NCox4PV6UNGE/vKwmJQXCvHc9WH2y264x2hg2
sbvn5RXVHB92pYDXtPzF1xX4NSknxY7EV/Vg/Tl6O2XDS2uTogZ2m6yI21eXivpt1PEzaq5G4YzW
ybwyegfvv9wzcQrh498HKbUI3HIhx2r4wAwzPtBIeLE2JZCspnbwwfTQmMBMhUA5IG85LGWondTB
8qkbtTYv3fbSGlegnOTSyXpA2YkmVYNCnu+CoFqJFNzcksqsazRYtWYmP9fgpgE7O8UBYPazpfEg
vf0kuZcSAq8dOiCzBoIUMEScuKeIkSIj2PO5TYPzPvuYgR4Y6UzBJMTlANgjdVPNqEWd1Af28qZT
8QNISmm9BeaQCnZQ8rJekewF2RJVIG/XMFesEJH4VuUUuFJObiRVIkwdW571xkKi/QsWB+L2PffL
4Tna0WDWKEXo7b/zHYFxue9mZGN26c5jrqB49pwru4Eqf0uPVDwOEEOc4/hP916MjFZapwuIp7VI
4MAhgSklMsznwMOttu9LRHoZtr0Pr2H72IJ0nujLAzc3QjZW/S2rAHhhAKZ6bilmUI0uq5n5Rc+s
hpjbHvPucSb76OyNn99xCsWuSl+Z9kuN6Ttcb/H6SJRXVNFz2OMl2rfsrFcwopBSnZuUVWIRdptC
z1XCGDl/m7xXYF8lHofqk2KaRMxxQgLi7Z//tVKqS7wQcVBMItQeDu3czV1VFS+CQ2AvFnbT0UlW
AhAyiQztCj/ahpwlgfiKHCZuKfbSvmPqZWYMm5JbJsEKmT31Q29/6knWtwbaj+hlaWWEXNkBVEED
DyXpT+4cfIIAHvWKRDXX5gpxGQNgVKnw8py6rK1XyolLrJOMZ0nkPzEkD/WfIfH4sjPjt7+wkKq/
rIIOSDXv6SGE3MLKHL/QvJVmFaosemmDnsu9e2w4smh5dRYn8hJUpBePPM10oUv1QjcMDMA1VCux
eamvDsPrNJJ1p9uMfb4zdGtjtoZdEvfb3zpi4xMYpRvZagRakMb4tZMGu99Tv3+Z/dN1jaFz/eMv
ziGzqb62nwrcTdXTHmy+8O5noEwtDs6vcyc/Bggs66KEkauLC+M3cvKke/oXouifDfxA/EFoCLmT
esShHMvDfriVqb1Gy2BM5GfbLaKOR1ed4S95k2obpKQLsBy/7t+fRwR/nVSxl+JypHlrqynCFfpC
om/YLn/EA9P5FTAHDWYvyfq2QtSf8No4DcbcaEXh8NmJfVlPnCOzz7GZQX3XbBSFd15Te3jomb1F
zRtbHwP0rdU+gCjkifSG1easSKUE2pBSZrqunkXFdpokYh75ZiwAan8Pzc3BipCiLXzYPcO1zhek
EamBlw2P1eAR9WQbVD94Lw2bl0MX9Zo8NgwpjcFUA/PPnk+53kUf06cnhwM+dgCqhv1ZWUlUXKa/
6KN3yfR+QWXhq1t/tGC1qE2nq50FeiU+3JOJsKh0n746cgUf8sNINPee/W6QiCh0eJmwRzeNsZHW
RK9hUQflI5iWyepr/icsF5hTQ/fUweJ7sMs2QiNKgOBOmDAWWOya7tAZatjVHd5IgmXCXz8bdIn/
ZiEqoxbx2eNHDnmYE3Zemj8GfyyJn2Sgpb/h8uKLhMlT6RxX5pLnhMwjCLN7tQw1uqyV/ODdLx8S
32pgrnKEXpeWWeD17L9qRKRz+joGiJ24az9aqct7XzNjLnDvRfj8s8qYIU9/UXLJBd8JChfMKXvn
cJ3AnIfZqFhd5XZKj6Y/2jLY3AF9SXKnemeb1r5vZL0Nzrvo1qchavJA6jfyypJmXbHWOkYV2rGh
J5HlsJlWVtuC92hlBUYRLshvGxK5BrmRcl9CRwOB/xGQhj2+gmqpit0MIE1avVjzZfZtj48sQaBz
SSyuBLfN4j/o4bwcJl8p7LyZY9lHXrIQy7fnUOjryzrlBGY5hJl4757oqb55Xf5o3UZxJrjcdQ8X
QESC39l34G8E/o04YujVXIF28N3fwGKOSPpJhiHKzd2M19PAgNB+YZFhkOgZi9LP+DcFubUxsbsB
er/89OUjcBlQzF0CKLw3iZY10sHeNpHFLj8tS+qxZYBbYDP7MFMCvy70Bp3HClZkAadPc0DY3JKh
4Qzr8HAZbwLY80JQOrqnegYuF2LFWfggoRAmZnPWn7bXjPrGpgGRNcOSV4i22a9/uzDs3x8Xlvfa
QLcGGeDrtZb76oMiJkwmiQxgccdaHKVtyEGZag1NOQKz4Z7Fta3CrPpzoiFQAbOHiRGJB9OcZS+d
oCmngtMd4W7KjIH6t/+21PqqLe0hWoQykegOctM/LpC6JWafdwfzE2CQijk80KNUKQJqxfK/GFBK
gplxOn9/CYpxv/eUKsR9u7bNO7C4RYOnq6inRqwqr/2WxgdgqS6CHL2kLmhlazXqnkXQDNfIdZUc
sr4q5E3rzYbC5IJrI0zQ1Qc6HNQj2I4u5Jgy6LJGKi3DsMuP/lTrrzyOpCoVouOXRimvbFsAkid1
cFRWG1P4+OUIRvVoNjlVmTgvFPxMghaNBA2tidoQWQ970bJevGYW+6IdaBix1R5NC5Vk+VR5NkVy
tkAQ34A+kkveQDpsROWO5IMvJUiMr0R0bsAEnnnJQ2t3+XOVB0e/ofgUN72chOxb9oQCUj8PbVUn
Cr4XEjoIFtozoG3rDSE3gh52xDXqm2LQNCQ1e+iFtYfFI/HxK/QsGURkLseN/ma+K0y29oA9tQup
M+irnx/LhihqZtAynNIBz9IoWF2vVchSqNmdA5ygJLdDPGrsKOYJ5dxS+htegpjdTJzSw9aMUGbz
SlJ0DYkEJ5ISs3am+K/tVWGlUShv47CrmqgylvNqfj/tZaPzXMk0GtnJrKlJXUx7de8L2PwGomdE
iKd6vSBzaUEk334YkwTMK7up1Z7wJ+sz9dsJxzBqcrSSlxFe0T78Nng4q9eqgYNIUPyQxNIqSblM
5WRfxotKn4P3u2swc6XtDWjFtvE3nrKdHttGlGRkHQ99OcI5azEMnnwpE32ipgH+XDGxd5BpQa3D
PDWlUlrBaMd6gB8w8fgMCFb7UtNZRQix0KQl49dK2rZIKmwywPZ0hEn8aeOY/xw7fdU6UA7hZIHk
dBk9UdXPhfhiDKUcigtT/JGUP6qG8e+gQMnCMLDORcdQ1MZ51bRGnvAhCy227Zw+8SXjy616rdJO
qhTcj0MEEVQPYeU7tPVJaPEi5uvcKKD0rcICbfQigHbxbdWMBjAChV8z7iS1T9bY37qnMq2rxjun
jN3Zv3aj7Zc4yzk6PrxszidvKozPjn2ZRg/+EWEqIA7xyYVLFxF+gqVpCy4ZtD6Oce7rCdN2Vz/w
v2mFBrj/GbZ/QXcYGXkYkttcL+fbTRxhI0O6ec/C9MTshm153B6i08Ds9xfh7O4BY4W5tRjIenAE
dr0lgocQKs16fYQ93dxAxg68V2GdEoQMrY2c7Iugym05HsxyqXLcF08/Y6QS1XCBV5xB72SxQEsO
vbTsQ1UHCEkhj65U/U4p4WUdhP4sdGeV++h/+3krU8cUknPS50EDJUpCMiIjfnCLWwPXdlGhtPhH
M3mhilYneKQnlX/tHGgzWlXytnho7tbUvl6Gw9R9kb1aO6qunIvl0fj8Wf2yeqAIa88O7X2FGZqA
AsYc9yfu1j+UVT/uzg6Gp9uzX8eTpnCdfwclVgaH0QGhi8hyv7B2A4jx89b5RhpWWCSN7VwRuxu6
OYb/t7dal6xSbHnxF5oNWuPUYZ7WVUT2iBjikAxOVuX8tN+Zl3wxTSF61jZao5Ur2wx+XiZ1Wmnq
cqTqI8EzPJgSLin5bD46HsoVf77P0/83zBILLKwaA5qd6rQ6bdGWESMKhxc8kDkRg0BiSzJl4YBN
ZtQZdATyJaYZHEEL7I0ZCztWSA4ef5gWNrcsQw9OToIKldUoSdtGnAZCOE8ybeUtqbCPWRaVQDfV
3BgH3C+QuYp4vFhdDqYIQLbpPEjfSSTtzird1onAgw36SoYbeyvC0PF5TTY8tiRb5DaW14WNkOcH
y6cSeHdvpbhLVwVZ9Ns0Webg9qn8BbW6QCfol65w0Prr6yZqoWiPUnYMc4BH2UQcuWM8JqGgCGet
+IkswK7Jlc/xF5m19gA7RIVqddgRIdN/jqEknvxOo7NRkIUDfZYNBaAi/CBY6sTqOWcz8FVlgdXI
pdreVmjBnJptYlSb2itXvigE5SfISJRW1YXrT3qbFwLN3Q6Xba5MJytH2EbA5w77cRcv0ljYJPdY
jtaa/NAfwhqPf3Mu/iheLDMSnP6CXVpWcj326AY8ptD8f85zPSMkTLFWqlx4RGtOImTfpT09DPi/
R4AZ3zD7LzrQwN34SzGUGO7T0vGWGwUuXcXQwafCkeFDkFYo4ydTdMmzjGn7W+jZOZ522maEUPOy
DdA+qZTDFxTieBXdB7QjD4+sRbjBLPZWtQWShounVrgRNgsxNGRZZHZh5Moyohm/Nqin/w9MLEtc
lrK7qxFyDFVXUYKHo5famQ2tfKnVWRZhaVvoduXCc/hiq2R3OscvOWqt9LxL/O001slWOHjo2UpK
m6B0F8Tj/NnD8csUU/MqQLrp/42CYLZWoJcJB3ylCt9AYFTK7xmCI+qT+d0044YsOXgflsGxKyFd
6baQ5pbxxlhIJfe+ru638IRHH1hFn0xXlNIEDjvKlWIp8sqrh8PgAtZh3IBghuwn/hxOOJTxKEc7
PSM/GNGnjoSgMvFYURVVa1yWBDITiuOB1bTfX8h7xQKfMfEFBMj0liE0i6dupR+r8cIYHAX69XO1
5ulcRpHtzkS2xnxbhaPMssyDkwfZ16UBTYIKNuG3qwsJBolLqOx4GyV0MrMs3SK3uBnPy0iSvlgp
302qMGxu98lxtb63QPCnd2PAi26e9If04mWubEm9FhYNAyjDLGpHnVW4jwjoN9rW4GSc/jxNgP3R
4CXIfVdS6sBxBvSmKFRxwQGFMZnbw3O1J+9J8uxFNbls8GrClVwSwwHxAnZZRxQ8HfnPzkMFTHQn
1nLBIr1R/d44aWlfrena6zIgY/Qlnwo7Z+u5SwGFn0mnrpZG5q9NrxFM3CtWlc+cnuGVi8kH2ER9
fb2EB89+Ykoa4z6RaAbWDaagt9BRAJhMsplAVrmO8sO32K4HSPsTzHj0Wkicw3l0XPtOlRvd2gK5
YdCVnWE8BDnuzfPVR2dKv4EEH1bwQjqJph9NhILCqhTe0Eb62R6RwIoqqExlmkB7TUvn4vx/7h2s
kDG1RPGWqXqwnhMESjKzTbz73aj79SLZgO8m0fI4v28f7k41wapDCjE+XQyza6Gg+gkfTWoL1EZs
0RlNX41mGT4bcO1x6fsPLzGhZ7g39fheZJ0/5us5x0gREZg2tgvMgJsfIZJjiBIC8pvEN5H4LzD5
7dPWlqA/YK/7BiZSQZMQtAbek3lLmso3eztUyUYEOkXpmo5na1yJoIgo94/pCa9/elKJfOkScMWT
cYq3uCpGk901pFIW7SHVi0Wp67GMDIXvlNyRIyBl1T9GRJ/xEqBXOuyW7eDNV6FYLp6HYLu3WX97
IQkEBD0mK7ZGY+WHEhMwxaJ19lM4TJ631VqRe5V/iGSeny+htEx2jSuzJSbFd4sEiuO+QbqWEcfU
c29OZsNGcJA2SepApQA/SKRQN+897WfxAN9vGUhF1zXrZ1aC1d1QMOlbI7R9KEvFnqavXw2CgGiT
dYkaRlTtl+SQXJLwfgITCFWOonAVkZTtp70zPI/M3KTxaTOADt+o42lCpl3radHz9N3yaP/hHH/i
/UX/7uctxsaChFBS9ee/e1oOd8j3ixZRUd2aTlmhZkhcHSry1z/re6EMRUXwbkulsrMpl8CUOfuQ
ZdorxhyIhrffvYvvHDYjqOj7La/CA5vv2oIaiAQsJnv03oBUI0TYb89NkW79MxZQ6uFHnAR90QLz
UATIaEQvNpoAvp5naVH+8N928HAvP1pQugzr48OOv+xP9/+eQXkU3EjyI5iaCWV9D61/T312CLmn
DXNpUBaNuEqmo+jQzvmzomoJjQZip0VkDvO5daaiw7Ca1NkAuGSkockluG9+Pwy9Ps/fpF9tryhe
5Yi4dSdwZw1ePRmzH9eRqCMP8c2P8T8pNcu1/lktGXIrlGAJPUTaEUnS35Ux5N4+8XU5GMr4pEdd
4eUJ0Cl1kYYKdraQpsorCgvEgi66uk0K07mK5PRDA7yQBhghGFyssMIpybUrHDPA/KCg50hokifv
3l+fhfdkUIciq7UWwZlTKDcuEZkJanshWdsSF6hs3CvySfdlI8kwMD9JBKcNu7CCXnxUF8jkLAtw
lgc90W/RL3MguLrryuAE4jdpdEdP1wU5OZKibYe/ACOiK0vIOJJ6FMUG07ZLyHepZDhOSeCL79X1
dMQAVxpnrYOESPdPQzV1KuEzhHA1AbqF3DbDTmPV229G3oYoeBHOK7kxqumCQbow1wNCcQVGXDZk
PzjitPeJyfqjG/hSILt86WISDUJPNeJzkrfZhL6lb1vTGsgYCVVeKqX2u1dd1HJS3uC2/SzYEnMl
cBoWwpIxO6FjLdNs7hArWyQnG1ZJxL2omTYt3XPL4ARUqTjxo2r3HEH+fJyCimFmc6kArATvVPmS
fkhLCqQ6QBnAaftXS+3P59rAcvQVwhL7bSj+pK8dsSE/3WGZz+opEyXC7+qyLK/ye7NUqeFUm/v/
Rzn0Vxh2sb+XefPH7Rm3m/p2dpsb9UBvlxNdTcuZGQtv+JR/W/X5SuRYHYyGrYGciWdv+ybMdpXw
B5BqmrDpnyNWSGlz5omX7IKXlmKKuDxZzPaAOlwFObp1dTpgndamwM8OMYEp8aW7tXibmZZL916y
6Wh7E1LXGxrd3VBSE6KDwMtgeI3raq82k6mEon8HeF8HBnihHyS7tGD3WQrinO/fOTUN3Ruinwc5
whz1eMJJVjU+pTH8FuLkLJg4+RVXq6KRxQg1q2542tkTFWbB/b31p8WGTcOfMlYezLfwXMOZhzF7
Zvgtxp0cBb/3ydI7l9IiP23Yg4KM0ZEZeS1BqAKJcIlygCYuy9zo6Iz0/MaHsORXD5SCXX8yflUS
s889si6u7LQu0+3xwchGeyfXtgXqNhul33EqcmQioE1NjkCuu5/RehHJBW3X9uIXllLLgavKPyiH
UQjx5QH5E8YMzub0E2yXL8S20kJcAgpko18jTfTaSnmuJhjOIGqNOHgQP+TLczlu63ObOK31BciO
+kx2Mcko7LgEU0EtER4FLgMFRvOLT1hpFlk/StHvTxZJAQ0vwsvu5P8rfP5FAqW6lO+tSE1wuNBJ
lGqdhUIWKRt1voDKKKTHs/MgljB1FBN0HawtwkscFQNIXKdFh/ZEYcJlSA789ihnDWBPwI+N+vcc
0fVx6YGYY61Lp7cVjSmDYEr5WOBqKLapfjZYigU/LRyAum/QiPIqHfCp+hHRpsPjHyh/boIDzxTT
OttuTIxyO4OXtgVUPTaHmCLIZ8J1A/9Xslov5yvgDAGA0+PbdhKeuBuFHNvZ/R+U1q6F2hWZuXZy
koeHcBOwfWEF7lghVevdr9LBU+wrEFppeRyzrWssHX1NQNRmiI6B6RBDEyUDP9m0aOe7/Ps6B36c
RFuQ8hIkk39SEkEJQiVZhI+MwD4BFko42lyWwMEGvVNQnlQ6JHNkkYjskOBgI/ZOuQRDhkvgJswF
76rCa1uA8/yqF7+g0AWywXuqnZdhn+navDAWz2D6sC1st8D5E6XYYk/D78GRQWvQhfklKhYITQw1
cOUdzJliwxT6GZ5OH92W40TiWy7MsYyXkTPleXHMP2vSyz5/3yOXzN1YBx+YsEXD2NKyHIDh4P/A
CCct4RVwL6jppF79hQ/X84we2aasOmChUJX79CLtyS1FYdVtNt8t9Qjqv6e80kLmShdDhPswqxo0
GmB4k0PvQ7DmCEKiClERXRjVGnEf3mGR/36Dgh3ad7zBOAxd9HtTcvct3a62CfyCOxue6YAE8moi
kWBEZKLiawFBzfLiMXWF1kTHxGNh6aI6RwSI3bMkftdTn9eOn78q62mmN4zwJIHky0XgMAvL8QBh
+uThvI4gKnqfg++yaaec7Wr5RBJxOTudf7jD8Ml1VPgyMqsoMyvhqVNx6uebcTolv/MtThZGypDF
tSZVVc9fIyfTvli+VmZ7sE6r1YMFdzp2xT+qUKAMsTueQJpf8T77tHmTtBNIsMb75bZ0LdSt/zoh
ZdZ3ke6rwMoEvBNAZm6nDbbwhAz5YdlyBzmu4/mQyWJQBLKH0kt0QIiqVT8GJIgHD3UU3LqrI3BN
6rzd+zr5ullI0N3Gt1Bh7mV55JF2ytIktGXqpojwxt3/z3rUJihAS/a0GUicSZrzN2evxMf4ruUI
nqw0ODYu57kwKLpUJ/nx46G1CcdXLSJUyKyCNo50b+7nSOxINLi2LWZ1BEf2qi78v7C5xrzoCQSB
bb3/qEseOIolKOiOnQT3QyfZGstZaE8xOSOuc8B87WndBuvJ6y4X40XuGOGjDk5fYnFQpUGW4rqW
+J6MKuGuDBYD0Ulj2W4W5e5Qdp8vjtaamz631U9zzS5N5mdyMCSDRG4B1KO0bJQR5Y4nCpj4+v34
LEb8xO+lj2BXaD3EG/Hr3YGAQaIJU6z/QW88u35G7aD7IdZYYT5xpNfVcFrLC+3rfI3oyuOUycsm
Hs7j6lxwrbLlI+ebXJHUmIlrGaCBjZ04ZxMPu2hbdAaTxwHyicLAiRz9qHP4I+wrxu/VNy4fd8VM
5DxySS6uQijUdGDVijW7lwDhhJ2pOLoVacqFkNAmQDxTJ9twoAwwAbWILG7jSejaKun+b3B1GJlc
mqIt85AQoxbVpwxclP8EkdcjGArZPNQXWUfWZZ24B+L7VV5Ji2t+GRxkdEl0Fo4MWoAU7HNe/dZX
Re2xTJWYSMnbmjotilY62KxO1qWHuU56C+Q7P4lldtY4hes3q5JuOajpyvBvmgeyfnufjNe7O7nC
x7zl68+tCZGHJRyaGXW7Kboe2+Koz6DsuxPJeixZJriuQcyZ21RQq7HNla1+uKwgRK1CVrHengQW
vhGMeIrDLA3RY5I3NVvD9UbGWMpEnLhsONHrvDF61xKzY2fjqIkNp3MXTBXXOr+dEGIgjs3uevBL
oJOby1axplYkDEB+/GkKiR6gN/cc9GzmZW7I/5mlpxa1hb0vk76j75DMb3hGmz5Ve5iL6RXOCyKq
gOMFW+3YG8SBWTha7YMeIzSr8bJooI6zrkDFWoDKCKQywU/6XTjL1ibpPRrLlnNQ1vdEUSevx/Ku
Ok4zMe+hpgrRgD+OfOJQUparUD0ih0HRgYnx8Ynm6kcZBckaWbhw6+6Xznlax74oYXPhwGJiM+0n
IDNxeTZ3hikSAYliCcUw21uK13UP0mALxlOLD0Npb0AKHHAz8+WHQRifaHwqn+cGc4Om5I09u9UT
UHCZBXG1s8bsim5fGmC1tVa0qPBGMFUTp7tQdxWEOIu+lbRv579/rN/Rua6kR/KaFMGqFlaxxRwx
q2s3ryFjjg0vI8xibtWrkMNzI7BlF+9B1jyqLB2T6H1kCM9m5MOCd/YijYKwYYVR0JqQVTrnL+YC
vC6FIrxKZFbFTzCHdTlmpwsyX7d/oamsUf5EcEYEC7NCcTCUywAUWGAovicy3sy7GAt8ClHH1am2
a4gLEZmYywnLBK0F3jIjZ8ihTD02uWVFNttMvD0l7GmUMsfi1nqRApU8//o1/gESW4vC6K20HJcF
LUb/DQcLL2Z9QNIR2piYItmMsZKKCdyw3B3TGZGPhDVXRkkbbz9K34MKKfEuIVd/Y1q/+1YvgIT4
aU2IPMl+WmK5d3+Q9oakau89NhJ8ECjCHJCbq4RULfprvC4+YkvjkGfYDvXNwUXKHL7GG2ZEIdO4
XhWCzg+5wL967UUg7E0HJwdtBOq7ge0x3lH7zKnAiALWoCiRYM1nB5rMVFvwlBvKc5Cp0Blpwqrp
Pl1q6Vgf7xKUDuUdVrzMRwFsSds9fv6dX7F9TSUfZK2v6077IZQFmEATuw6LRBNEb/KucUYimNln
3akL9UpSRCRk75eiji/N8dPtrfY0huit7BdeeNBY9oQk+MsvNHa32OToZ/8YLb7cWufv81YfamtU
TbTlGfwbdOZNhQhTOsCWTp4Td5SV2HPGm4Tr1xEzGn3ANRQ5QkGgYq8JujG/kA5U+P9JQKlCsRCw
mjqu1rmlBb6Dr30z9/+uuVPUOz0FL0/RO7yzYaZJ1o50B2aDpFBMOJA9TpUO7joIsgFRHWaW3peF
jnLMKMAsDCP+QN/iPZ+7IXmNCgkedPZOMkTn9NtM0ijIny03V77n3xgTh1MOtE6mp0HiGxxWKdmp
CCQDfDUqaQdyv9oeC+npKVfskemPalmbkH9dj3kjzjFv9NNTUVCDq7HXVhoDYXi8/0JB7DeOW4Mo
wMBgTao2KPARJf5y1IZb3BENu2q0ot/pScnYYNyXAVS+XYPIIiG1Nw0qRd7iYbOx2C6l0VEu+i4b
DeyEW23waDpJYRDMG/GEVe3O0dJXkhWWwWp4dCMnKUYFAUhxxRKWQPrPf7IMgQaA1z3DnmGFqBNs
/jgjcT3m6wjOUlaFJHuUfR+f78AYW9DQu5zgS2iVfTSV/CJp9O04J6vMgYirs4q/chRHo0pDExef
3lC+XVMZYuX2yJ+xxzR9zo6XQ3QHL2MhOKbLdMu6BQJdtzLXxTJpyzcol2bDm0+PtA8rFIzNG+iE
zIGwgH6wNJ5PPUTFr9os5k6/mgFuvOqwEAl4NymZ8B6sCSmLMXXovmbHSNqwkabGbvr1qRytosTQ
Aw6Aak++92GSVxKFwil1SkQYoHM8n0y022P3DLar/3+f8YROBDjFjL3Cx+wLyu+pkDZqJczqyFA+
o4N6oYNQ++lu/094Dwh2psUPSp6ElvXokuDXvgpIcSSvWLUlKAsPIPpoSP/vFKru8W/ZVxK4CoNm
9xoOZoaozHEaQ+hrwyP1oGme9E7+UNaR9wfnduy4u/VUNBp2rN8wvbG5x5+Ei23vy8O6ssYU7ldW
bpmorHoSt+eYFfpFLpa7PsiEwlOn+yBwYhMYfyLZt2PhN+t/cA8b8fKHfJn8wddNWgyQqp2GkbM1
hv1cxzfCpGXn0XFDUMx2HxI53ZahqGjg4bhzN1TpzGStQg4UB7IyDuSbDouNV+JhwFVh8i7kXe17
jQ48THG0luk5u4D37tAPbFE19pEKDi41+emylACa0xjtoPA/ZBRk4nK+TOaUXsnftPsga7gHd3kT
Wu5E/NVT011qlrDyq6YeKwvNES8s2mF49ITQZGP0f3FHIQP+h77NF5MnJaTt0h234XakeSp965D7
LQSZeGY8fTHzXwv90JoPs0iTEYLB8lqxpyeohBuE0ztHVWRPmBpjarMypCLUbO7K6us7P61Jxv43
fGVyVd8yMadjFfJ9Z+yoIHOllEje16bHmSY4qZNGA1pyC76gzZL6r8ucY+4tbIABX2N0ZbTzRUR8
C8Y6DWT5yAtXAHJZFDP+ObW9G2OF9UjWEj+NWw+U8+V6schOtaxhweo/1G0HqPhhPUt2dwJmxtnZ
IPu9+XNh05oe89NwAjHiICkHKzXeduwopOP2243B3TFPYjmqMUB6lmBKxeui5STINsdY8UtzZKoH
DLSPYnskYy55NlZxlhhDf9D0tsCTTOBffZ1MYjlZhYUz5tPRkydPhgN2Is0itGgbiQkpXe3Vfhj1
4+RYy9zwOph50Yd+9SytJBVd5RCeA2nXMBkNtGgYaEkwmSawyLpWwoQ3lXegs7qoocDWPf3MH+Dt
qBGreIQts2B/Ss/XeI0h5jwyObKsYpF/nrKR2EZLxmGq0d4WQokfEy6GSX2g6zOTnijkQ2U3mhaA
Urna2Xg7JomKGYAGwYd1jGHSfXt+2HOIWBycCVKOvHI00yRp+yUFYDnzdoXJCHKDuyPeHgbcnS8k
YVEY7NNaAEUEqpLNjFLf5/6hHrvWhkLv3LZdOH9llIRboDrVbULfOngq1mN7mtIKCWcreVpMkVmB
BOJLIaClLdB1L+8scXEGhvxHE7WQB8vY4bUdaDL5ujHrMVoIC97qG1NO+9I2vNxCNa8hdJaMGMiI
w3OFwNjH5DYANoFTxNeG4F5mbFIIgumheO+4ZR4mGlW0TaTNYKqXqJlD727HaMcXWo3YK6Ng4cw5
fmrxDQqJ+e+8O34gh6AuG7Jo/IKgRd3tcyBoQM2D59w+U5l76lOV8lx9Xav8tb3w0iTyWTQeGHLE
qfoFkCjsBjIC5UD5U9wmvJyKQQh/GVlj14tiHtSjIOmOG769VVJZ1hTcgsG5Hm6tXHjd1V+F3lKE
75Wq4azgYk/rjlpCv6jEDVnZYjG7tViN+Z4+yS+miMsYAWO5obVZkNYbIonIn7ozizyfsoxoaA1J
dAnqTatFS68/vtc/swnpMpJWUaAwEwfzDw0P5q6zqRwBrRrEdLUKgewSAfhxiVvtRByWbY0WDUks
toYQNTHstHKH2imp2K2RB3n1vdLXwwMC5ccXN2sASk8o+DzlHufo8tI/JFdxSSoX+VSvUeB9P8Lw
yEgcXZ0cFz1maVbxYN++s2nul54toXPTJnR92dwcf1wQbUtqUQiWdjEL/4Zc2rqXHbqhTi01KZZ1
/8hXX8Itz1SQdWvC0MDd1kC0ix8VOHrvqzSeG97K5ffMrp7docOZ+be+XmVRmS2DzMxxaB8pYZBJ
Z075bDv0lKOvSKy5qC9h7GRXdAe6dytIcORHcpno6sLQKP8eRG3AVplRGPo4C8HCwh+rcBTZj0uP
D0EdFya39aPUAhlmhOu9hsXPOrzBg6CInUVOp36LvfRSvO2bAxjwPm1Ztu4mYr0WQCKn+euM/1wa
ZoRjz7Rsu2yXmP2fPrZUaAyU7BTjYUaV2zPiDuS6iUf29V2XpkPbjg1TxJdBlZG8HJ2aVjA6LLVt
bj4aege5Mk0LTOqHNtQHnQYJ2b02kZ22bZnSQ7DJXcMHQ2iiXhUFM0eKtRiaXxXNzL25jkzRxq8N
NFf3ar4xmhxVnhhzrQDeibh5mT2U0nNWi0Uz1dJ5pGpPaMf02z69Tq0CwjJA2gE0GV9EnoDg4HHl
tgYQBqHokbMvEbV+mewBAI5KIywmyXRtyYm3EawWYuvTgRlUTIQMsZAOHkYKe7Y7X/+i5GYf7qyE
yQoOxYTRNPHrQo1yGLqe2AQBwC5AQdU5KF4kq+sn5THrDJB/L+xMSEiGjq7dideVPRQQWvB7Rf/n
5e2j32eAaVKxW1jqjwCggBH0pRa1ni27FhLwoUF0OKB5DGxkzUiCL7xrXe2n3IUkjvSo1fo4/vyX
MR6EGk3N25+RGlkBpQH2ug2HMSAtYa6LmoCp4AcNvQL+3vti9xLFW7A6WHq11VQRCgKbs7yh8KYF
w1bfNNYDS9RSNihryan4/QwD+n4ehFA9gfQLdMp1l3fGOO1nLtUecLtPuhk01TQtdmkz9840KBPO
HZ2z5tr0RbMkTNGE6p2EiCYD3LKSjBeVXM+fFpDDaxTdtd2/m06UqO3DCCQttyEe2d3+1vqBz5Nr
yYjv1hN5wY8VR9Z0Qf27dK6dyiZzFaeS5f2okyUgd+mW3j02S2WtuL+GWeqd9OdZkouuPV+G33ma
4YL6xa23dRE3pVKtwLbAu3CNKklt7mXYigJCDZqW8iy4MX04A9yecd2ui3LX7bpYLHVDcjQBhIAU
G0uSPLTzWYYJbcsypbU0DNq8xR5SVgGHokUNTzVgKMYtZ+CSPppKB7xV6glnP0WftB+nCQBFxE+K
gbAFoZpmhePsGiHyLvwyeDIebAD6PT46/JqZNOeRXqxFYiWY5apAdcXXJ7502X66YW/FlDIcbdBa
6Oinxd7ursTg2Xr3JMoOr0LNz4QuMIieake523qbgPYoPZOKxbU+H4uU+eD7O6yxFcoiEEBk2HuQ
JuFGtQS2kmmTzPUFvDmmdjqMZT8XjZxhJJhIR4C7n5SomDx2Cc4h3SdmAr802foEInSxOtVQ9L75
Jj9NQnQtfMYGf2xLr81LJjNrJqM4xfvXuBk9xpFY+EYaano6Voby8TSDn4DFJdJs7vuGCPAR137O
HEBPF5pPfrdkIx5LBe7Zp1QzTLMMqzTtoOXM6fGGtkPHCg5NO9fmxYPS2uOau/IRgSJLvDSC7AZa
NAsQH75F33cUPK1uzSXMjsCaE5l/YJ/sRCCAJqTIGzzFTRaeIzJy72TCpAkzZeS6NypMVarQeP9A
Xf4EFjKVyzaNL4p/ce6nIoOpPlAK75edJ2B4z4BAQK/Iv1xef/6BV8ohX74tFq8LgBFXdSxERTOS
NvKIcksBFGjmnJHWWEFMSKFtrKXEdXQ9n3oz+GI0H865E1MICRHoSXWAO1Vjre2Sl4od9Y6hrGxT
ww4KeXj1VytlxvtsJ8suOEWGtKks/KXx/khZOFK7eza13VjjfKCq41TK8IedWROlcfj9tJLazdje
VBbNUBU0EMF0ztge8VSh7KXSZIw8TEj52A2p79JEtgJ8IUhKm88wXv67P1u8h/D+WSxYtFQptJq0
gTe27Bwwfvt1iAIFn/brM2fV4bPwRaFTtX5ecCpwVSpIEuSptOXZz7dqib9SxXyLT5zBdtCM4/Yu
b74eCj1yJqmTGne3TZsk6067Nb0xMJ9iYR2XNfkjhe1WYVI1qPlqzZymSAZEXkBZW0WmPJduKkM/
Gx5e2LZLRtxUb9SdQ58t+9elNh2a5uPFBgr3hgBkXZxYFpb4l3wIQA7WQKF4liMc8m6zpY0uu1P6
LU4YIBQL0LQyMsNWunZ8xAygGNK+KcOOkiNq97Z3TsRW9wkgoU2qHoY/JvOd46CrFZjUIxvaTjSQ
EiLm10iPIBrjzF0ninL4vhjuKhU0Qv4I92Hdqyjn/Zp7Herwdw5vk2vFl59EHLq8NwiyiQ4efAVF
DLu89ju8kV0onm0a7EPQ+/cdSvA3liSh2QhQSujeWcwr0Tp1GSkJKJtZ1p3INBsRJ0s2mplfnF5r
miPERzSG3bGKJFcRrkYARXDE6Cz8czHwcZ1jeR/j3avsn1/vmclVuFI0qkFPEKNnQ4lx+sG9mrBq
pbQyl9DzI1AneSoSRj6V+Chd8Go8+AOziKT84vREuNz7mcadrqcs4v1lXSY2h6efVdWHFPA/O3gJ
fUS7WOcvm1csfxw6Vja42Q+5O8D7oi9Pdnt4rgljXojX9qneXLbMGHSphs51jOyU1PUAZ5I1mYnT
csrM8U09EhaNakmVKabEyVv+y0D10F4wYEmj8Uw8kKecnaAbupVqG55GYYXmciVzxfOIoVsgwcK2
bgdXXUY2UNbZQpwCWR+fgegzs6YYwklcM23oJLasiPvGVjhry128VjmeQeXGXuMU76g7RmBC1Gyo
syWyK7Gdfa9BiGkSZd/xQKlMklrTxG/cRoS+Px6MkbC3azen6X8MrXKgpy5n2MXFTuPyHbSjgtct
4LF+1lr3Xii/CBxx1OMHQgEzDGUvt0QJ3VCCnnWM3dKA+HY6Cltw2XOqFNGRWvmjEnsxeob5/+9e
HXsXnpHPD5eKVHaCp49ZBBLCks1mXqwdd8lu7el7fpHatyTRj1ooljc9qXxEgaHm3ELb+B49AZHr
BOetmQSEoTF0p0Fiao4YYF4vVFUWimPHCqbuQiMniZcPTOkP3OKEQ3vwco0ZfRJpDBHi1EcgjSiN
UwEePGygmLQADzn8QFGvEBmTNa5CMal52Fbub0+89fd4buc4nIsmTvv4N9m4Jb5htfWBda63k8gc
+6QF6IRmBkEsECW8brHRavCusyqUrCidJuxWKvHvZEi25ZWmbgHHlFX2/IQW5/Aq5ZH1A7P0JT/G
v61qAW/hyIXAH84/nLZ94Xy+Kr8iUxsRUDJLp8KTFW7+1n/ur/um+3UqaKnh6LEhxRjC7a379VVg
mqeo4MflmENMLK3MwLiACtClgzd3e5du+QnkHlTusaWfx7UnTrNW0bUJDLjzDIOd1s8fb4JFEamQ
eSkLP2gafE1Vi5wRLyOBlPnEA12bgInOu5aJNTWq8aea4wLcSi3AE49XNvsIrYVQoykNYtfImlMW
MfnX1G4figXM4EUsR3y//UvzS6hgI4av5xNkraKMe+6YdCoIxqz81G6gTlzDQMZkM0mLSDCwbHbZ
Z1KvZzcszpNNl8s9bj21qgkaFMSvM93qjlHYx70rBAQQQxp36KxTw2E9iceYhcYaB+RLDLWF8R2Y
lWnhW6j2QqAgiTDcsqEhsZlRUnYC3lN9rKXG0xKW82oCqNFSzS/+tnKxJiCX0V8lR+nc9QB5shoX
DKzFVHqFHchIM6DF5SXFxYvJvp13UWh0XcS6KYowTy2ejQFw+xD5E4saIWfA6nYo0e0+sqK4pVCp
Kim5/53+dkfIqkK17qBwXrerDULNUE6E8622P+xyShL6GfnscFv3j0Ia84hPiXy8qj6gfbMA/twZ
UVLZmPb/kqQcKKRawGMxGwhUj8LhcMg0L0Or9tFI+UxfAg/dlmsM/NvFSehP1CcwP4A8yxFkFqsd
TodW7Sv/Nnm7RooIEBqDZLOzdKZ3KNRWF3vg5eCnIWsEj2aYDAuRHj5RKAqbW+IwBf+tdI2yUEdq
7jM3sBmMtk/Pd7G6PYLm5KSF6iVEEyaD8uACc8PQVw74v3WZlcL1+sBGWZNoyRiKwrUR/axw8xYk
Ceh4EEf8nq7JRObFQjDm0JAHSRbhQ9godfPtnOTTF4lCdzDEVY6dk7t6tTGN+I+EHuZrAnPmn9sr
IpdzRIJznIopoR+AwbdYt75cKdM+0YAMWN0WNBIQMa7YqYJR0hd2QziL8UGdq+LeeJyWPUt1y+CS
VhiIkudxOL1EoJUQkAjUqSu7qgQYulGnU/RlylKdQxFLlUaftn/4hexsVZS0Pfhw5qBkRLLmgYOy
t0UarVb99oFwwtmkz7yPL2qeLjIr0V/5OFh7yB+oo92IUgg2hBiulx2B27CQ+JTXBjC52MyiZYqd
FGke/rt/tD1DzG/zVZpHF8BOQtUiOCpd6YI97rObFmoo1iUCM/IWR0MDNcWreeeF7OmVvRkUpTWO
qwXLy6+RcSd0CmmHsdJO32cBpbNp6Vb4HMqEQ78bb3P80BEMoDu1JRkvP/cKTlmFP2340Np3zU1/
wQYShOhIh2aNxQkhWQDr2gEp3qqRx0ZPS3ChoYiKG9MprrbV5SC0gYXmcNUK0GGmPfxYXJqdSkan
Yb89QDzyzeNf50f02pmnmfGuuPXDWBGUeo2u9bCGtO2LarqDBaN84MojETfCo+Pd4/aCiT3mVVCw
fuuZEfRnx+S6dLs9XFKs9ECxDOYqg9feorll9qCCwgKbTfXqOWrrtfVQSPMU/uxt2WXMwBvB4su8
pg48arZpaF0yXp7DBTKeGIQRdfvwfFcIBFGaj9VM7K5FznOktH5zGV0tbzoNpIzShkSSwfcBz6zc
tmoHujrPBc3zMCxRx6ZSQ1yyvgSHVa4INZ3wGNmoyenlMOqo6vRjQBS1xnkOCEWKEVKVHMKoGS/+
7eUsi7rwdND3p7CwVjAukXVIqn/OKKb0ySgA1OPs8VCkl04tDCQu3N97aI68bVt03hoKuCnCLd3b
zNe7SbeeSNcNj/4Fp5qzP0upU/1fkJ4XXVpFQjkF6lCuWBDjENyvcq41nEMYeMpJtpQeOvgX5QzT
emDsSwFQT5ZxhTtRQosKsYXX16AblVeIiAa+ni1juPTZxQ6R/pkduKmDssL2ZCbgS9dial5atdkI
9sesbZOdJWCyn6JXi332czZeTDf2glVO6FQv/KucBVtBE9o7M9YGOQlZZDkyen8Uj5a7uCQ+fTBG
g0r9fWserDFwDTnCAkd7gpaKYFGVt+pcVPneLDBFWg2WvufagaiSExjKUkEe7C1YXQM4gqaUD8z6
7kSS0iiM1+a1ZWSvs5dkUqPO1M7VsNw7NKVxeF5Iub3fvLkfxPiu0dMYZoJXKPzkgvXjwCat42fr
kXK3dpYvzUhL2BjRw6Zsv8qOJnYUPWhSPkRjq6dd7463V8IdiqXEVpUbEFuMg2doRafxPEX+w5fv
uiJqySVeGc9Ed8s+FlxsU8Ryq7ouodR7n/oRFK840FCE/B4HZXw+yaa2yWsxhB9KfIfwgYwmX0Xs
Fy13zD5rrMnuDuLoIUT5OvlGVmC6vMZ6WRr9Tvwrd5Csr07gsCZfwtMerI5KlOtnPDAZqj18l7Kp
wr2tUQuQYOuT5JVuyA1xmQEUhLkUZSoHgV9QlLfAR+mkEZ0ybj4KHH4rTfzsKnDZDdrxeD5Iyftw
OmTcuYrk2gQxWKxCXXoAJVke10VqNQ+1DjebsUnX42SKxsnKC307nVAFBqx33OodImpp4SgVoTx1
qxzwtSPUMO0uMC1EXzw9kK3PI4vaODJFRIS9PUQ4KcdqUdEzAgHbUKGgLT4YAkRKInhYmLY/p6D/
shJ+kFIw3tOrS5+5mvb9UGjOQjNSA34XrtQ0otwPNRwhViAW6aCE8ZV+ehzHvVkIOlWBFkVgeemK
yTEIBmwd6aYAtCaa/BAXSMmJ99eiCw8G0ev0GSufWmOGYxn0NGpHA7u0hM+InVuKyAyru5gM6dXE
977rhNonBVcr6+09QLNvPB9pITIlbgyl6QwIwVRyPsqw/VnM8n28unAna9A5CLdKoRfM/PrgJ3wd
O8KrP2MRyW5A4zmPF5w5S6RpgzE4XFkwrSf0+I23bg/liPlDT0GCXM/shvosKFv0rzal+gzPkdwe
govab8neNXnUttl43RAYo/YEHVSwTGUQChOyTdBqnhWdzLT3Af+eK7OS5YMydin/3fecupQRCxFY
KrECuB8zJz9lIJmbNVWWx2SSvFPNwPArqoWgMcZRybj+d7Q3v5FuQJd1Vm/thfMPucqxckIu7n3o
kupiIhm2oXDQeuPl/6J6IIHM8/01QsHNDKbrSzli7+X0rOnOTW8qfoQ2b0mgmLUEhX9LswV4YB6g
tuslujCqsnOBhKYfnpuuoLrvDb4Im+cGNV/dFb9DyMuMpJOf5GrvpHWY8nX3NM8dtW4ZAK9/5BWp
UtoH8R1IaQhrf9CsklvqlLz1/lK03MD9T3E+23sOTaMegmVMZZEKuEsxBy8zMgm01g2SZtBaFoW3
SUSa3G+gmB51Eoioe6xwvH1UoQ5hbjnUQy+b313SVXCX42U83SqJrdVezbhTjZg5DFt/pH+nAAhj
ux90u9bxl2SsWyl2Sg3Ttw4pxTbFglpGA+jKPmCAvNA+1/Ihv/nABXmI8N1kahhGObV5CHOPmpaV
zD6KAxkq3EFOunT72qLKIY04wvPHrZ+Kv8wNtDCFJwkCmocJPiE3XWW6bKxojpQvxCSCELNeY9mB
EcQTB03nU+bHSubtDcDxeMQ1qS0C1R7fpTRn/jR2hR9arnirfTAHcMO0CsG2XjMz0Xjdm+DhC0pA
JgBVUpedcziY1OoUEQYfL/kJ+sFca4bmhnQpIgE2ycyrcemLAWc7tCmjL8Gy2oq/aUHLHEcmjaf/
A+9IRWqdIcLozfFtANT0TTioG8HUbb94yDV1Wxy/Zxv0kjpgM4rzg1sYb+tjkavyRUvinDNU9oce
ATjUQ/tdO0tYorFuLNMJK33R62RQv1/yD/XUSdS7W32Z5KTm67p7hFjFVZiTq6q0spLu1Vfdgx/7
9sj25inERA6JidFftGV7vkEuLOEA3fxrj7WRWR7VRUYiCOqidCifUgo1vj9q0LiBOxm0ArEVEJNy
sL2CItUdH+AZi5Di2e18GveHECE5bZlfVskAVqTJvKZE8y/1FuDsmS0gdrYT2kq/gfGDw3DogFsS
S9fXyXFcT3mvHpIn1DQg4Y9a3vVu9gsuK/5hVS/ZjQAc7pN32v+oQWHg7VFnhgnDIg+7L03/YpCJ
69MM6/WxGsPmBRSU5lAj2qit9ydpCdn4l3iQ3MdQgdP+3btjH6OcY+sVZEOD/bmBku3BqZCq4337
KLMPYdPXeewOTvTpjm+XOvoCZVG7AOlyuUX6uHS5rOD3HaPYThTUX5wru4CfKnaavej33xMjYIMF
UzQoWLweMK3ExFyra5iP/6z04JbgS0wBvxKy0LzTOTlc9FQ1gV8uNw1wVeVP5nNOZooHBNd/sPiC
Thn2RpjhebdOFOGGpZCASiAT854J+aBob7FvzOpwai7TGBjRBa0iJOYG31wqv3BO8RD/45Xrkdr6
+yR4jinAv6vnOndfDLjd7QKvGU4r+wTWV5nNykkOOYhzFpA9RWZdzfI957fnJb4Ag08RLGPUx6XH
szz8JxA41bSsc4gRJCbIXnN7Wj3rX15RQ/8nnPiksV8dn7SK977Y1/y8O5y0YzAklZbsB3eCvjQw
0ncbxvLL55vo56iDFsH2qJ0OHl3qfkSnV0YOBaWOXiVYYFXU27VPsWfPhJccyri1gK8psBqSvliD
jfZwVe0/07d/VQ/KAuXtsVQ959xqki2UdCVVutFcF5/s5jWzbzdUDpCV8e3kOz6a+pjCq+59ChVH
P8c6IfVonn7K5150yMekD9NWprC0tOCE4wEAJiqOu3vP8JLJCCws+IrbtJGZPGYTWaVRgVaKmf0y
7sna2YQS4JepNiL5zxCM5LrWZWEmlnuK3zc0fNx1XhB+a2AnVbTw/WomoLXjUnTOB36AFvCX8bQL
l5Q46uZt2qU+ItUFWO4cyM5qqqoAn938F4Ykp1DLu8Zk/XUmgUlGzmxVCrHKDSJgwD75iOeF9buA
vZNbMi6+9bTUwnKWHe/U+LhRSZiE37fJsfZ3agqi1VXLiqubDB31Vfh1Rzym5zAhePNQIIG77C4l
CbGR3WBNPrPs7BjISgxaoBtfe/f5qv6QFzgle7VLRr3A1BvgLv1XRMhkTSeFKg9xaDg7hnl+rTet
/quJowI5DiW+vCntCfhrY42Giz8URW3stza6mwzTnXYhSis3F8SH+IGhlm4s7Rw178B9ob0mu4LH
iTHyO/f8mf5FzAwSSSeFFZuFy4ht3eT9O4KtKB+J33pm8zwK1jVPaD6WPR6hXTO1H4nXSO4/XY27
GGdIwkKiVKnNsXaMZltx1SKANpXJ2zpyCPWBbDVQ/2I7Rq0k1BJuc+Wrrz1uOMDmBoGmU2jkjboc
1I6DAM/VeylMa70gYKthyq0zUFiWFcC/QX7lxBe9I4eNyqn0jJiawbcsP6ufsuYFv4w68NgXyJTJ
PMa7WinS2a4ORiEEGGTCU4WkYHFIIXRuTWMOZIN+yDiofBYGPjWYCFzj1LQYuqPPiGa/wqO5BDeO
k2HMVbk575rPPErR4PWV8aRuBJr5Uduj8p6TxXMXqTJUa6qk9ehT3mGcWL+2+f/23opwhEJH/mFV
HGH4geh4gYgvu0wJp3yRFHp8V+qd4TJKuELujQrdPnjBLbeRDVGdmeTU/PSI/rW/jL17Kl/6eL8Z
6YcExDEfx5sPQXrRbiU5DtS9QuKXFypx9gciZmB4fsUSf2Qmd0rEIbneWDgy/l9Ua1j0Hjjm05tb
HLXRU/9/NecpoZQbJWlDEiESt3Wm/73aSPoj7du9KoqIHq09wZQeYRQKGQmQIXxAqTdzNUA3Yto8
qrAKMbIYLqUhAuxgdTHLkHFrYJWrhXhxUzUfa9JBa9rxDktn2lvGxb6qleqFbfKV2Tcc5hvJPv54
USyDWfZU/Wc/JnbLcJuNs6QtRyXeUR6MM6zYUQTVKQWQSaIf7s279lH+x0I/1FKtmOrJYta1I38g
6xUp1o9U1makV9BVdpXpUF1mug3EK91xkDaOVge3Ffj2LSa3+hsN8K8Mdss7L4gmjU0in6g48fad
pLP4i4vVps22UCiQJoHqgJp4QPeC6RKIzAgD2eMMv45V3yxSMgSZ05xCQl4bUcxh3dtakE3jzRI9
MnKi4RRgqO39Pk676uR/q8VD9D3fO7vEn9vgEOmnmlQFoFKTkTZwUr/rYFUVmyC0Y6A3be/S28J3
5LwVv6IxMkLnivnjtKdxtJUMAB3T0QgKE+Bs5HpWsgm6cZZ6LlrQR1KbmhmGTNIVfcNQfSkBf7up
EaFI6lYGykgTmYOdDs91otm30ojLAO94qe9bmlNvpaP/itKakdHxa95tfUkUbqqoEUM8kmKc5xSL
NbLYSE+2wo9qDq5RRq1uPCvorJ5sA0U3LhtXh9dcI//Xw7aH2nJn5wva9dqsvC2UbwOWl4kP2pO3
zLH/Gq9WyTO177GCvevXtXEMPguZD45bsv3TzMH6LP0JSn8d0l8kMgbfPk1N01dKvFAnmd9Qr+Mo
TP0iJgjV1JPza7PBOWNeuT9stOa3oAiCVasMxjfMPYDiH3ZbMkGsHAJNKNeQNieRX6fsLK7xXMe5
znzON8TVyW1PITGabKCAIazvb86x39fMriq468bVEg/5Utu1XVh7i9tfOqSWmVCpp2jPDsOgZuFZ
ndqDP7SNW9+nn5D2evmlr8vn6YVnmdKKCgh2euIk8hZta18kRfPkTnwa+pCkM3KHhjPPNpeeo4QB
jVlbJM+mr+oA6itYPMqf5NeKWcBfLnzokJ8V16GZec1PjSO7X5uzGMaRXgg4e/y0XF3duZxHDsCH
ReU6KIBAKj/xiSeZxBIDdQA+cTsHJabcHZgCLWKtoZ3zcU0uU7o24YXyYt33IhtrJvJcwdzww620
jy3LTyqjCSiBHiRFU8FGNdX8FiWxN1xyXtwJoX8blZ5QRhhJFgPu8tPfP3vTMiU+ZRuQQzwYjZc9
dNk5t5QkulrT7afjHK83z/SpKnvPAGe3MV4AO4uf4O1u1EV5irUbXv5tTrs2E4LIJfiBKd2IyiO8
u0Qk+x6xLUNpK+GTEK26EbNhgs4SvV3C8J0MLQIbC+JYKe0AemqS/GDC5jUMPIeNfGfaukQP0KWl
CetieshK2TTNPsakkMwojPcEp77cNypG+DCOCNKDIPSg4/BsN7w7z+OxaVauUKk4w6+36azH2IjJ
OQRFMq6vMlCHYfsY/bY/W74Ehqo+g7XAIZVZbdPBdB+ul8DJzDxpJentxAkbft4tLOV+y1SC8DbO
bSAnbkZ0vsanGePOsoAjhomTnDg2pBdyWbIftC5cZimTlPAe2/Ey66e6WSZ+rQ//eIIpce2rvisX
I2r+NA0nCkVyMBeFWA+c0DPi2WmqtkYzvbNwrzT8Hv4ncbrgH/LKaT9YFt+iylziienOeK/p5vWI
JTo227MYh8GtjXXBZKly0D3C5+eGXw3GEWtqG4Zo7Hh82jqTrq39SskGYSO49TnAcHGCfqK7AXuG
UTmW1CG7GLM6GNQJMl3SDjJUG/8L80rKwPi3khle8Be1g0BhdQeQ5IwedUTu+n3jc0ipH1VfxIdf
xTpN15Rq+QL9qixr1CakPfgPA9D4VRETvVACYzsSP4eCqElxGXFId8kuRGvNbhpcDwtA5X5wN9HY
EnY7xGCsNN9VcqVw3yS5bWhsSelX87ph3XtfJWR53KZbQyarqFNdTVBPrqcDjbZ7NPlal/bXpWaq
1II3GFAg0Cx32LWaqENuLLYIAtaL4Zyyd89WcLT/KcDkCugTk01FLH7cT30VWjiW2PFD64hoQSX1
UoIGFC1mf7KAaZ6wbaWnB9FW3uDD1Il78v7LlOhNnE1nVdaxkn/x0c+xnrmWuDsapg+9+ozB9nqs
VakngdUGKVhCaEtYdmXkbiZ3lgxiNy9IMiNsg+A5O4P/1/74dwiKkWQHgpYRnEt8p4jyr7yYgN3J
HoF1jDfXJAGiSUn6I2Mj+Is97JJhrpCqDJvWAGtYpVZnND06PNUWdKb0ejDtEUQ4d0ds9fVSbOfR
93YLfJ1z3YYzRWGBUtRhp9UbQ3Ivm3VlDsqHruJPnBlqSsoOKePauJocAT2EZKpnLJsfoInc9iJ9
G2oBDggdUagt2D6Xr++t3QUaofRXh5+BB4oG3kqebEfS/KbiDbg9McHgkgKvEAKmU6kYRg6QCUoM
bAjaW0qLW6QNVZH41ghnuWFOVf7tWejZowd6M7LPewBzG2RxOdEihk/WjufRdo2laJOJe/wwbyhS
tNTHHibEg55djlXlQikZeSHMuKCVHs2bv8C57wYCkdqM7asExiXVuOkQH3/o++kfI9V4wLjNR6W+
B21fcl8AuCt/3jxpU6irvWD88R9MZxtLl8wNgnS013jt4MUe7FbT25MZDLGMHkDSXgB2WrNbwr0r
ncsZHVTvOGPGAW08kF6lV+HQjFh5gGL0Hl30A0aIAdgMIlkQna6USACz7Q47UnP8O1GyS7GUr0sk
88oIZsZatt03bKU0UASyuN2y3+tPYHb/6Q7QixhFTn8EIMc2E/I+tPgCpB1llnaMZWqBp2hqVBUm
2hJoceg/5xePnSvmORWJOwwsxPMVhRBlkCoFG1PmGKy+svodJu9kYZVnAloOnzGnU/gICsuWmD5X
nSGhtoqGBcW+S/9MCCDhQxQZQHARDngGIeR7DXT10ASPDLvj/0kWk/Za3c0Qtdow0BNWYhltv9Ft
EPjBC89kNWDCYdPl+raVbQUBLOCjDm6d9UsC+yhJy7U5aZQifSH07udzhefYg8mY+u1mCdbR8QUt
3e5mpz4DYndpP89MH+pGvQ2fz7lhchXCVqAFx2h5/UBoyhMQQ/QYolb9l5hz+8GURxFzt8Q36gRQ
d9+S28cq9J91ygOhAjJP75ZfJJDXH2xM6d8oAfbOHXrgR0W2yEpxJ4wQfqs4bRqqGPToQNbLsK3b
iA16wKqrHlNmiLLFSr1zfV8b5rrdymMY3RCzogkX70e1nsC0J2Ue6Z+lcvTCEUVpT6lb6Ud+5+FY
v2bvUodi0vSEEmLJgo6k4eMWN7ycnJ9JGHBF2+VIjOnDoOvcORdmt3d8mLLtD9pYUBWqZkJD5hk5
8zrKhZWzHNGPubbjedIwyHbRujXrTPXySHjdzOfqzOXFYz2263Etu7lac14cx2Ofemd9LnsyuBCn
QRr22p12T62/3ip4A6LV5em1DNjn0qwbluzqDnCjaeLZ1Ri4IRtFti8WP1IQD6IwY+O5O6YGxdDC
QVKpmGE0EnzTmKnUl9oaGJFfMyf9zbLMe4llRDvjrxdKdM3Y1rC9Twf5bWEY047jpm2g7b6BVUft
kG2iixn5ZhOBE41D0QUZ6JrzH7z7gpQI3o60wkw/j1sy84CCFKqB6MOh11crtB84qq03ia8dPGW6
8sbQ0iJvzmmSBAzSqbONHZ34SxOU22rVIgrhqlyWb8FBV2GXV+7CR/EW7Ta3xsuquUgPLbT/01LP
UpBZ211tDQtArRxPUvWtk5BC3yTCGX211nMmWpG5ygkCg46NpvHnSTKiojN7KxjbmY10cuQh4WE1
hivtx2yTszG6tTRaCRG0A+tkrRfacw/Zdnab9/0bu8TYAzXGxzBX2Vm6YuPtYWJJtnqOguqEkf/F
IFfewRxcINw+pkId+llTw00gYAncWvTVt9DrxKpH1h9b9PoCl/BVBrdF4308ntlB4Mj//MfvVh7C
lmhmRTgllL3wAOYzGPqcqE9/u0pfcD/Fx8zx8hN2Ke6Zk4UMkMCWWtROwEyIgCrEspMxid/o5ZqM
E69e7dJXr3JknS1Lo4BdypnyFOQGCpLLN5wSfa0qBKUwB7x6r0WmOl+ySO6tvKKe4liNT2sHQNhu
16zvRJQTcWzZJzhW7MK4DbIeXkbxeU4SXNxN+1VG5xJkf+zNS5g3uTv/4bW5DKQTjTYQf3vP8m7B
VTTP6mWBjCzPytskBsGPoOoCeraXiBSUU/fS7pfPXCAPCYJxgpWhZlJUCEHhD5jX9rjAX+xXdgaa
aOrqdT4hBpekSkphxbIxz5edHSfGrxaPrkMgHXgcYSbePQdZQjrdIP9MWNbaRuf2wb8ZDiF74AXX
FAE22Wd2AUMhfdr8ga+G5Kp9XLSwVOAgrz3o4gsdvNl4D8xI2Xd5QS46Ug52HCnz+WdxB6R8x33k
CGv5e5cNwFgTONK9GuKIzDAZ8jeQkTWgnAgN3d8Zny1qF6VHl5u4pSPn5ybrF/UbXjSrGvLgIULC
Ts7ZJk3eXSxDDCwpOGM8CwwZLkRW5HI7yUjcQVP26WG9ox/4BdK01RXk6+4sICFsfvtfijiT+K7I
mScEd+dLVXPg3TFbecTsNPZFEScgrjMx/oAddDzxmgJsWbCzTe9tIeIh7kSaX19kbeJcz73RATl9
azigqyz3xHMuCMyk9Apm1/Tbef9Bo7WpUzEOTDDrJ1A/vAGQaSXBOoGXATKBcGyhHcnAXRz3PabO
BYayXuPrc4hnJuzHbUzO1l1nYA7HOD9/UAShlJJuosMKNQmcvmDejjeffTpdxS+paQoGIHThOtJv
bSp46u8S6ZQJ8zMjtMxb5hSD32AIxlIzn33y9y+mtflELlo4MSW6uLnQgy9j4JZJ2cSiumKX2Vwm
cslad3G/+6T2aTephtXkqryXtquArJbsE+Cv4AxFugHQP1itQgJlBuL1U2bCEWUWkR4BlNz83YeB
2GWzxdCcEdCN9bLjSGbE4h5KLrd8zeoUqnnCW3/tUscNE90zOtLr6gpNGXx2MyUopDMTJQ7IKXAq
gZnNhN3Q5/0meavP5afP2E8dqHuX59RTR5ZpZhWz8JTdtfoqPiHBBdKuFP2gi/ur7RgVimdfjMZF
1iTjGP9OxIirv4iWvzXwYrjkasW0RpfEDifU8cpYGa53XeHTioMpbPZvHJmPQfGiuFSnqGCxwmn2
l4Nk+dXNpQ4c5cMfeefMYTTpyyHGJ3vXRs27wlElYisRwjaUTnU0te+flDgcjM+7qULoiiPuq1Dz
pX0Gabcoyn2fZBDRvKQKm+TP6X4eqV0rPLRiReqcfVkyhjo4gQQZFeNG6iMxXPsnzIzRRHRtdjWW
SBmTX2ajZUlYJAypPi1zaxOh04NDbPA6UMR+6f/TOGqbgaAVEmLo21PU8YYr0BZR1am24O/UfFHZ
bkF6Yzk4JQQr/OMWDvAwqF/+/9DlgWL2kR37b/t1u/TK4j72lOw2VeHVud0omO4M9ZrPchC5AXe0
bdxOPA9Qlv5WTue6q7J4Lc6BPEQDTBDBmuplPWjZD5XD1NlnT9moXglmI4VlCOzviCdVVveUgHNV
c7pkKgrSqxZqt1XIKwWqO0sM4zOSKlz0eKml9/thyNSPlKFRxFk85yBi1AgTUZPf1rOGWZpztmeQ
AUiXlJucYZq58L3zZSJEYAZcOmb6ysiBQfMMxGKlwQ0AvLVBDv+MMzDS/IsnLjvPEY/nJxbu0Q0q
mO9mtYTCtmYthwNSp9dNMefMUtTZxC9n+v+tBAhZiG2jCyVXhn+8JFMCiwYfj0HL/OXkCzV+m1Z+
5IQWiouIuB4H0fKrjX7fo0Yfylc55qboZ823esYdPNqCQyeAJtFq6XOEnmGaATnbC6okHxYXZjkC
5vyxI1tiPtvqg5DchZt1nTVVeoOpdLvJWz/LQOm9lQD+FowEIJk3uFPmmZ171CAyYWdfYGa4Hyco
g6NlBmBwPDFXjH/bKJO0laxJoz+Dm2t/2Q3Az5jQsWoooKPbRIIdgswwEX11u2XQBS9jkPZlzWe7
vl3XpCMjAXGPfQkT4jNX8c3CXHon7TDM9qAEC01Qj5z0fbSUTpBQNXvThI1YAhs2iWo/jcdtTVK2
3f98eML+8s0wBNn0BPlpwj/RrSs+LROfxVgRCWWgxSrO5HSrWFUhoUVJelVbEWWXAddzW0CqIsnS
WIFRx0q9AcHvsW8624fLilQBSDg+fL1QB/HSUmfL968Gc+ehfhc8/pDm9Jw7TBjEBcNbvTRUAP12
7qt6xZ8gUS14SeYJiyf0P6Pt715G+/kxBBfcB3eS4NMTVz3WXgWyLrPgRslPdRUZzjrJcGq9EoO0
7OrO+vzm9udgEwi+vltlcNaJY4a3qYmeOeLk7VdY3nQAGCMF+7lZ3tJNGEtjSiCFZIZNw5qclEG9
mbI0lXv+/o9UDN0uAlxrettNkGwDWE8hFfIO/17H0LeQ/h0MQ2/4Ci2Fjh0TTxodW2QmQE7pMIhS
hMCFh0JJY9BK9M7jm9cI2EWu3JnBAewfb7bjgqkdJEdnpx3lgqNjhw3rQ9St5jL0VKSCmshhlZe6
sZSgYm7Th5jAkjqRstksvpn7kxnVyqHadBSZZ1W0qsErgVkAdkaAP+Pe4CpJUBjRf14XKXHacjuC
BREysiV165A66YWuUZ7RVulMMBcNu9oSnOKMJDTE8U/SoopdN9RPgg7BQCFxlJnFCkbUH9jOaS+c
LmOa1dGxFVi6VwrEYKj5lJwrj+fVXiFIVHtYBQAR7vy83ct2lVrFD2lQ7cEKesqCuIrkRXXe3Vm5
1h6aaxmUgmVc5NxIp1fT4Y6lG+cK7DBBke9AWU8iyDviKaxC0nva2enykBkeEoWXAUkFReUQ4dvN
p3PV953gqnk6TT97pSc3YRR+OWKY791whTl6ye+xLkoXlwnhmu82Wyp8qsme5vxfShJaF3+Y22sT
to1Qo9s5+6/YUu9n2ixp4JiOjxigM7CjdmzwXGxoFd/bGG7Lb0Fpn3Q8hayx1p7ypZlylQmpm3+w
abhnf0SswwbsjpD1xPc7cVXnOGu/40Z6rorlO0pHCTrt4E/zgeE0IwfOaql+HbeLy6L2y9s82wLq
5qJOwLnVS6M/HoAiiQPwHGLT6tV3OYnOQ90e3AHV7uOF/Fjfpzb1fx/1jD0dCY89Y4JI1oU0tcnL
hSAuL5jGALeREeyykLC7sVkjuBszy69WUVqogvcfv6EcARHgbj/pvB9Z1SXbtQgldmUoy2h6Gj3a
ANFdTUDlSh0HuZG6+K74ngB3WtBDEyDnDTW2xLoUCPjCTQ1pXtaqhNysiF9QKBe4Ula42vlUYu9t
++zeKQeF9TrQH/pzXE/Hd0ukm69IbwA5PI9v+Y+wd6HMEqzeyD1Kjh0Zf3DvBaiaNyo02l4avJkE
gQLbV89JxTqIpaml7KLJtfVouFcLlnnztBZlQFKbPgi9dBHOAy5Y71kdbmu+J7f5ttKJ8WeRLHkE
XEd/n/lcTn0G1EquQVr4nHW3tZg42h8Ds4iRpaiSjeaObZMYlPrLAiIzkIunlTVVyVWm0QV5d0QB
pJButLL8VWhMRo6gLEGKGy7temriZ46ZMmmK45useixCAA0CeHyX3x67QtWvRvvcRDqGKoGuPBH3
ui0wjehbqqqnBg1GZ1X4CdO/sbdN7fEEX3M8+ihv5PfRYNeXWni1U+HEwWTs67YJkI2RZ3NNoFvv
3jm6FP8rIUcv6FqA1uNPW58bMk7Dtm7r6FOKF1o+zIHx0jnEgXjuOkCpbkLKtcq/cC3w5xsK8ctl
r/wkVqS5nkKQ/XpG7ZrBCzVVaqLP4N9oJdhxFrlzDfhtR9mBwMJjcYPVf1Paf6LxAhqQfYa8k1Te
phJ49U22M3gNrOQKB/diTIXopVTmKIgZi3i5OmxihhdJ02AME+GBWQvBg0Iiov70PtIDTSFxSS8m
mArWdamdiyH1xchkqZEyoATy78RNRXY558rqfnoiezJz94x1GcBlnyuhjcycdQeRClQ/EnLXK5fb
gVQtbJ6zBlOPzP6FJksiG5RRHJa84D/6olCc08J4eHk6ajMZplooYfpElm80djqxBvNh9gmXkTrw
YsPDt93Cwfef8voFtKLs0Oo06iD7B54yAQG2apMWWzwhzUlwquHBzjPfb4Xmk10Qv+Pr594xnk1B
IKhFkrSK4BFlBpS/MuWcxANFvjydtszIpVNLuajdb5eU73r8EZyfNCuptypwJFDEnzXIBhE13rEM
i11icCaT/I9AGFTT7ZqkQGShU9yCNqceyFc5VXiBdSfbyuvrsEoDyww/s0LZ1XxgLh7XrltoTq1v
8qY9aSe77yQWIJO4Ss2eWJvr1kYCIXrtXHSnGMgG+TAbBTNDeHx1VpJ5MlNntc+0CT+v6MOdrZ9+
vPXZC67UBQ3FNYHKvbH8rneZzsGCRSXSNg/Qys3S8dY6QL44iPlzOb/ASiA/EaGwMn3MmzDGXrBx
ThXVqHk5U4ej4Wp4IUOCRbYFJsE53TOYAH1iPTD+1a+1rwD7j8794TNyvlkFzihAuYv7h/3Yzp3y
rD2U7T6EIa3lfv3ma05Wt0Av9TuVtyJ3L1AZkgFf/OtPClKBdM5Mcg7J0bKVI39zsACRBF7XXTZE
GzJyNuLUxtaWhRpgi0B7RpaReSUi7WJLTFJdSdr5hSt4w4IoQjMjgksxu87wpzgM5WoaUhYV7tow
9JB1o1gdRhN8YDC9v53fU68JrYetnMOzEY4m2Im1KFCZTZwHiBJOo1MnMHfozitphEtqb1fjlmnM
R9uEp6pe11ENiGQF7SwHT/OdWgj0baFDb9U8OOneHE2JsEBHfk9BIiVyAcnYW1ug1fFUHVnZwNFJ
ok7jds/LyZg89t7TqiH2kP+5/jLmAGivU24QCun9qxyoZwj6sSUsYtd/yi4J6OctcEcOm3FdMKvZ
Jhs3w1FyaRRYl0RC4Pup45jbMgrPMg6+aep47ppg9bB8lW1eTKfhSAlO1v6U2fMcO912OQ2+SYH2
SSfo8MduTbNy+5Ty448QpbPkgos8zF8WnV1+4VBTrOqayZ5f/TOLqx0rgTUvkwI9JPC5pkEqvykr
eAHmjMChRPwnuCqhK2LXRFKOkC74x9fUr4HsMWoGpf9X27gJGg9/Qts6HLOWCOO9svok31nS4u0Z
8tWKoUegJ3SHlRUPsKPuZGA5daxrFtP40SmaBwybXvnY6AJKUxFvPf85jA1R6NBPqfB2G6WX4GYe
GFB3Xu4Of4FR8nyvauCEWGg0J1dTbgnIgMslJhkwDnZato2gcm1o+Cmq9V7CjphO0Oi7vAlX3x9q
9XEHiTZNoRVAWtHiCIyDca/ydGiEOH8MhRqvYnaQibOvqcWeP9WnQ66DBL1Z4knt4DTlEsz2TT4k
VglbAxsZ18qYG2yfXYARofs+oYvOAj5/E4AIkf45CqRQ6cf/WCRzboFCRnTkxhhJL8L8qXX95Y18
zTQth04L4CfVhBm6F9ZIfp2xDHGXrlY/QOih5avI4f6E7qlEK069vQ4kI9b587gdUvPoK6qT0M0N
HbK9D9L1wZRh5EyO3Y5cXDPGIgXJLhr6CC/d8Zu2TvC5RNonzHoeDTt/xd3ub0/BMWz8D9jYNfqL
L0U0OOFb4hIOCx9MlhIy/PhLJpXRPMVaShVhseH+N+75CA3DAX9hNhlxIUuccmbRJXaUgGwYeGSc
mpWn9mtZ1uETQQtzXmzTwGrk5PCgc35F6JZ5Up+PG0uQK+Hk9ZhzefK8df5SXTYdhG4U/xzB3nw6
5g1vWMbvwf/OfgIdNGV5ysQyNt6rYaO7PI8r9f2L2hfOheZLzhzA1fLEfuEjFov9hyaMGfKWvN2W
m6NQvY12zSB1BZ9v3nmfURJa7SX7ckkb8sydsSW6nRiejmoZxqLxXFjbqN+FEhkyVEM0SFoM0vMl
bJ9y2mBg7VJw55DGeUNoveQWUdMS2vd6iR/aqb/7yT5HwKn7+0r1DMrvLY62XyVJo+wAl1hO/+/B
1pD4fPF5sEnPVO4zTFs6Nh28cMleNfQcX2YvsVpZhFUqUA88KcCOLtuljcRI9IHAoJWNB3dK1WcS
cVte50R9i+4uJc0Zz87VWxHDfhExHw2J4+z6BwCqTXffcEFe5hUFbWsa3raFueGOKiHnTI3GEH0U
OkdVAd2C/2hm26Xv05C32groB0sZuC2ZJiUAJSydZXmsDWNMJx5s3ViSN4AecPzxAi2M1e9wjb42
Yn5wfrV9+TZIfdD4F2+ovBynT0dbxquc8dsakC6SF0QgWJXG/wmsWr+Hs/jesU/JdMOadf8nju03
/xcJRwdo1HsbZft6ruuYpqEN6kU/aZ3M1nM87ov4qrp9Ee4VT5aRhsVOqh8hPXort7QpTGSFkSsb
MddjGp6i9+OsB80C2xfYck4INYfcOX85kogBL2+YYnuBmdxM1g0GcRvHHRnjsP6jHYWtulCpYEYR
nYDq42KL/MBkPDhGQbg2+r3qMbr7uqkSykqejVfrvjezssCSfeKy8QeQ2hDUxM32s0gz/VNnvLiO
CBx0UCFnBY211NZYjMaukjSWC9VANtCC/MYgw8BV3qkniuSfi+TCxTmmhQIlGSbU2wEjFSPrm/wi
gegGfqaMisIqgRH+aRPdp15SJuAJVwm5hv8PzTBJexwl69nxjevg3EyqVowyMnwZuzAHqiaa+keX
i97a3iUVRfhuA8CxPZrGhnQYKBwC5zxO8idHzXN8g4xeueYNE+BuVAVz1QwxvdN1iCzokNJcAtXI
higfUAKjw+Z0YuPNQ5z4ARxoOh+G6Nx2+AKuQJi9ZoqCYwEWQx5xqCvy+Ag4NkVaf27F/lJQpKON
xYVgBnyQtbOAGvn1PF0r3aqwKoOYwVofpj7humGh3tOoNJo/6yGkk271k+hmldwU17lHVJqbeb11
mFnU865i8KDTgThJlsThaziREYVZgj8iUMDHMLSsQI8TFYi1x8m/F+ArP0dAT+00oeh/RmZBcPqJ
P4+YEPPUyshWKEW5N1UetktQ+v+MQs0rsEJohqFuKlQRJlDD0MVTUQJwkYG2bzb9pGIfXBbJx1SC
8kpIJgopSXvg9GNwGbYPRWDbHxAYjGByCxdHvppbTayOmP5wn83coimCN27ir45fk2GLb0YpdOYf
UnfNUt2tmnRziqOuzZ514YAG7VjzVQcapqoWiJPEyXuIoLTrfzv2eX8qSWoNNvoeWBJ5c0XteQq9
DzfUCiYZYlM6wGtAMGme1IlSscZWQxy5n/TqZ/vm7oXHGhTzzd2a/LNXnTR4flv1AabxoJ9ccFiK
bOblCC7lSIZ7Ylerf2xoGm+qy6iDZUEtLITNADlteEDXzCIJ5z0UkAZxXvfguDxMw+ws9W9ghBzM
vQK533C81HPCvcwU1ULOYhkp+3bCtX3MPWaPHeSucZ+lwHaxMJ12x8DjhyfgzDwL8x4BlOBtJukR
nHZN4sOhM8GuDubcmDf3dHmx6eQPd2wteap0JSxEyNBzOlqMIvbFBOxPzLSiFcimB8so+PlpIn+a
jBtPy7+i3spOnWVVpSPTXEL2IJ6GJJtXOiV65uTBENtcLR34lo4AH8SL9TtltxYnuC9UafIJRIFo
ZHd5iDKugywTedFYGXl79LI2Ob+D/e2eiWPuQzezU2+BT0xJCNzyCTTBkJoJDRDntJ+6UJ0K+QV2
D0zsOrLCGdvihymUh2BtzyyDglNUkyqfFLV39MP6s82I0KKngXnh20eXGtJIsABeK/qVmVF/me3u
UF3nVXgzAvxeu5m0fQqqYJbjhjnvXSfuRlVWNQOiDGH4j3k4GMOnZ6T6nHA4K0GTS4KnRBPaXgIt
Y4kGlkOiws33pRmYM+ibAwnaPP4UidmPqKxW19kS+TjFdnmJf6vxWWRa2ZQYq6KP460TXqIc9GBH
ymxVg5xh+t11ixAbuf9v8RaDoZIOUU1jRRhGgUR2bG7hBSnCZf2DcS+SOznbRShfG0kQJvW8MaQ1
WImkMcPryZNFtCMBct1E7DCv2N4/Oc+WRA8GBF0iGJ6AO+aSQQSvlWn0g0qvn0v5qv1EsNlkCSWr
PXFfOlhedrUvi6OMt9FtUye4AUCJVUCH/fUFOgcVHDgTFiGLKUaggRP+HlYk0XBKNzVgy+8Vxc4R
ms4OE3Iv+Qt2uS+nhCJqHFpLD01eORY8g5HtSmHCZh64WZ7dQOx/BeorO6LFxAdVrI7uICmoo+1i
nmPMrSDm0QDlHD89Ftur1D+HyhOwljbSN6QG2fUz9P0GINjUEBax53EIUUn3RZctppXYAsLUyEvH
2kX+cC1nxK4gpipo4TZ8MZrgFF+C1xfjXwB7qRqaBJvt5A0uW7i0PXGzJdIY7bND9sW2c+PWNnuJ
UuA1w+eA5lxCp5Swbzsz8iye2dtT5/oIT0shnTNuAGpa40LILIo3uHh8yvN1JK94m2OU6krSMEOE
FvcwSeveTAPCaIp/dnlC8DfLbGj2z4uF+0GCn6Rue1CA+mMAHHGfe85NWkM+JTLyMzzQPzs3pAFf
SA0bXK4ONHSZzPKf77z5JLzMDnmGxEVz2fQLcHRQhAuz8HYswpCyeGoZIQLaaX7IbfBDTO3f90gx
3nrdXABzAMD8z3hqSMb1uXXZp3PIYB7p49H6X/p9xw1M+wICM6mcCURjhb/278L87wgE9VXVHINT
5XzfaQbHIMdwXFFVkJh/kicto49A3LIemoBknmXN8Hm1HFonrBrbo6I+eJQXTcNVVcd+eoFbD56m
n5bR1xwn/FJUANEm78qiBuhwDaGGiExw9K/g9XQI4+zjiSn/7A6zi5A3YPuROQRkITUhd9pB+nJr
CPRqR3LuAbCe9PjLIKsQIAj1Oy2NKqqmH6KkbSojRT/fnZ8e2pSsiWXv/nK9sIZ4Qh2fKsyebV6x
HdSVFpM0iP1bursmfhgSxmGgZc4C2dKMgiyNNn83ROZ3Qzj+2S0CQN5z7EovDEtPZ02tdPcw9EB5
R4IuRlqJzNeBRIr/mz4pL9qqKKUwiasXUmhxKAp4+oa9+EfZP3DCmZ4eKcX/BHGIFnwKAcS26bMZ
auEUuuJDWtnpuGYOLoqLTWkf0hpr/GLSbcm4NUDoxJEEaEohMZjN1DsR/sViHaIKhNeu5Pm/gb93
cws8gI+CmkihoIVY+sfsvSr0TJ4s+wXUXiJeYJxdyqN7DDg20oLvjxhrQoXpZzkx1+kiKu/yTQ+d
KDrcoP9BLKVrSNqzQgRgl1RxSY7lZF0oqNy7FWHq2RC/Up4lbJ2PbxbbF4N8Z1KsCmKyEetET4tl
KvRbJrCCSJOIvBlXEgnBWF+4t5fQg+mno4LymM+GO//8pzZlvh5MUERgm61n0k1Idv/SnMgsHetH
hzlIlyQxfH3O7chbITbReF+erUWzPkFb9NCK/wujbWPjNE3PK6ZtBciQlarAFQ7Fcoeoj+j+8weR
QhSXxS7oWedZFZioiUzdK5+Eg9HJvdiMQKldWuUwhZA1a2PmgoKnJu9y387IeCqSAxwqxAdNIr/l
mUaVEJ+z0I2UapLNsrXnSDD+e7T0m/38WgwqE211GNL80HZfbY2thJ2JWLcxpj/HSUmJM74SKjJE
RqsV3zGVvfFXIRx4liIzxgmDDPN2DkRK1Pk7Iv6om7SRf+Kr0vajUyGiyR9V6ooTp/gEHMuNlNRW
agZ8+mByM7dbesk3q0td+a60QOPUmXNuWVrxK2DuFKRn3dGxEB68GOan3d1MwZPpRodpCbaDm9WJ
+vU54A3GcOF/lhhU8qyoRAyHzlGRf9MoSc3quMf4KBLd/GNZ0hBOz59L2bZvsUfHhe0+5UzTPceP
0qIvw/iSXHoHzBLx4Ja1Z6BRxQTBPJMPE8H6SR3uPQQhiDB/dsiH2FCuGYr6R3ZeFbDJ6vQ+IFgf
15GnmoqaAeAKf7FfFMX8cYbMRWo8vneqyfpC6ffipIHgHfyrMeKKdw9XgWDH9eQ6+083c662qpaD
BYaEawqD3EeiIRj2WB3SGq8uthaR+NLFT8/+UAxwhH9LBDL8JFBs99z5rcbYfsLbI5FzSZTHK/WT
qZ8LM2a4wTjPGsoLysJoGGHkqFjADAJETUSkLRByrrLWJYMggr+VM05WDNEXXDb7sU7R+8thg3C7
jh/1jgWlDXAQXOKeJzvJSNLizqFGDqTVpHVgmIbCpZTZFO5xaeL/yGOAqiro+2er0AWxMJ0cHMsK
2RLaWc96qlZpyYPE0kyRXLBK+vsw4EtkPGAvDFCPKxqEZ4i4nuf++yLL93dAUsLM2jewP+Xb4sgd
a77W+ux2LaXJOYidkJV5LP7QyLBSGEb4StWqF+u4Bqqns8diOQ4MwVuvBLfle5ZahbcS+wYQNbFX
ynhbwIS+5MEFGWONmhedHOMlvCEFsEYX/n7Am1JBpvTGRwG6hUdj1wFoUik+DDiRTaHr4sPUYyds
pPYRT5Kq4iKTeSrto7UH+4MIkb5KEEcN94r2TXse/n8A0D1A/AlK0aZI7JzocrCben03MMux/dej
/Q0Ep0vd0t+WVgyJSMGfN9LodBKD1yFAO5lpVrqsTFztoRTGMFAxmdWW/eVNvKIuDaj6K3PuInnx
gragn+VvFLWPp/Cqat3DH9xDhobVNRWwnUYsrNVAKJI1zU+hsixA+jJk+c1g8FI9iCIrjhqrIi64
QPJqKLntgqSDEwYjwb3mgtefEA65AasMqICupKeSSi5Qammis2VEld3rCgcVk5Za+6TMkgcH1wRU
8dues2BoMAW7IjfyiO8Yx2cJj7/C+xg6Dp+DUxlaDSC4VjTsOBcDbc0HFcVgJh7/mTJOlo8nKhp1
Dkj/JyHl6hn8irmA6L5sY3mdGgHREW8NM3dK0/bOWyAXZXK48CwTFJI3/GMW2L+FPpe22TVu5loH
nfILfurXyjEXvqqqN6iDRjgCaTSO2xopfA6W3xU30RaSs51ohUGU43W51EcwrY6aw1LUrbu0UmNi
DZRxqjcALYRq9jFe5TwqJWqwpXPxBmJR8zvhK+S1N9tunTmw7e/BpXu6ndF80eLdxvjtwcAWean6
+4uo+eSGx5OhK8LbFj517tklqvtB/P3WPnH22g4HtlHKYY9Q+3OiXjVIoYcg2dhsMaUHEqbR/1as
1sN5bhhVkAwgAVvxf6VeXaC3/gxIHdDDa6bu2ra4pcXaZu/kruu8AoePVI27DAY0XEkXc+c4Y2Sr
uqBczds/t6EQTkBHOp9TTG4ivH74XMjy1NgdS35BYgnlPcGdDWGCo1eawTE/L8XUMWNYXRse9EMy
QddAzbGnqETTK1VAzsnNw8io4ia8kZWOJnQQh7TztpRpkGfztTLmcHs2WC93vTPeoPoYBL5By6x+
BQQJUXYYMIfY8FslxOe76RfAP008hU8yQXzC5CukdTWs6uuFGyZ/BqJzMsVrdGoaj/MC7NpMY1+w
LdXkMLgYudjBNqIwpbXuS3cMbgtdyJsoBgPDfAzbLhZts06oBxYBFizT33W2NM4YIlInbSXiwPUw
cS6uUxYxht5oJ7TMRGG/pWJJdhGu6ZLlkgFSYRso50gRfPG2piZZsmtleZ2TVkyf722iW87mPGJc
OZzhyd3iFYA2c/eeKMDkFP117O6yH/NYRFJhp7g7TkjnJyXjXriNVpFDqIJl7zvMuvZl+YB2IACS
pjIKr5FtgqwsrO8v3Jvzcj+lEZk4JnWxyEdi8L+TFm34G49x8jUZqcWwrJLXlswvFk+D/CBHRlrK
JABST3bhpJ0Gpx5JsaYEP0aiB+dPvM60Z/ywsMbDjO3LqVGTtNOGEv1ucCbpHjVjTaQ4z43+BvrH
gR4r2wrlmRdTS139GAD183pZcAJ79v/xcLHMuUYn1VdNBXNgYiK31WRU6dYM7NNYH4mjpZzuHVy0
1GQJufHPpqfYRLCuX9hxblFtoXa/kYpNsf5BqdmSuVYfnCh/oEUel9G3jXSYn/1Fcevwc3LyQd47
Zub5RKDfS0sQwAKAHYadeFfZ6i3+44vItr0eN1IcNuCMezS4ywG0wgGlBkhlgyL8nuzNwtrIaP+f
Xh6nouc7wnvEPUQpWl/ZeLLKcY3o5qHFumt9+6b3bKub0wo4AoAwEVmq5mR6pxs3nlU2m8fFu165
6bh7XSl7OY1uVcB1q6KPzG/PR772HG+4UGAUPeSNVeQy/9wNUBpPNQ4YReoTy5oN+brT8A9xX5rM
s+67XQ1ty4NQE1neN3DuYbseh1hWpUde4uiU04u++BKZtf3KRIry9Feth7+KhfbuUABCoyC+A2hR
j5eaGrLoUPqFsfLhB8isUQuG+/fUMHAAS5W4o3B7NBtmxpXWAU3wyMc+GEZVPAoZj27l9AppQ7uA
C+o5qOYI81IUQQvOADa2QC8aCsBfU9rGjKwSbBCWTFOWZGS4Z77rYymSX3laCkhkU7h5HNVMya8y
qhi80QIpokGb1OmQlhumnbB0Q8QS6Yl7dmKpjP9QQgdAVAnmMoB8U1iA1fNvdzwQbpF+mEgHK/fW
W0/qJncq+DeM9Iq4hSQA5KvKufVEYf5GmCP0lFE6E8Nr2R6tavD2huBTUgxK9qqdzJZQJhhzrfft
Uadz8alozCdP30L9MELZ2jqUAjUrWJaOmQvpcVQmkAVS9U9VMliT9+8jRDhxb7v1vIeYQeRJ6pQ1
eEl7IBqRrX+j372a+zBm769KvsOCs3cRHJWgd2SFAHAbeq4rJKR9bXx5Xd1R86zMJWu53Sjk2ooA
FGH2VyWQzPRda+4WseXnpZlxjRfmGrRI0kyx8evP3GLg9krH646X8qFs0D3mpNWYBPeBBIJcvHdz
jmdqUc4FeBx3x4XcUBNO98P1d8g274lf3eptxolmvXdHsJgwDSoWGkqxlfMgVuBiKyxcM1704aMI
WrGyq1WRiqC4v4TZ9o/N/oBbvbBT9E08jJESiMpNyj2dzcLY7PFt65Cj24PXVnylohyIdNLWRat3
XlWTrowkL9OaIqf1P3nCvwdzMXe/wtBH/zX+sAbXc/pvugtmCXQMi3AfdSqrZFl3IJcEyCMjilld
bLfHM3ULUgdUaly3VFa46WZebw7sx1HbGibSfMsjRudWPWr5p32A+uRzezJzuwdIyHPUyterXjAw
iiXMpkeQHrZ5mfeZI2/rzMt/5tcstxsIUP7CU7pK+eMS4VdMazrqoIoERSuJzIb7YDWLzL3kzY4K
vX6OCNcsxWXLIgBZvJRnlI4L6SkluYTVK8CFr10BUzRAeSCXt2av9LVZ85+/hlVg7uobnQ3+lqCQ
jkOmLx77OP+7r7S+AVJjvGXOBf2uSE5VPcjirdqiCdUbeFYqcB7F2V8zuFHJQubTycq/bkdLBybW
9sWO2ch1+/CmZxpRP2DWvN65xRU65pstruU13vsFRjpq5cXfvKYvLMJENw2jUF1KINwbI2Ugf+ye
t7qaqN5z7QBS3417GiAgm+OoPXnVUZapeCPKHywOoeDL4papovwLDzROH5MOI5pivM+uSluC3Rwr
8sgxtO9O89r4JrvaOBEjsc8NUaNkUK6Nk5MVLxLSIiAk5EQIkkm2EBBVr73zXVR8LEu7UxKb+8sG
G1euITWOk97A6Y+wWbifOm10qx5nuAAYNPNn2UdYphUz/St3qB3wNTsNCkDOtXqSVRvf2hve9xcu
qp+IeV1K+7X9nBi0HJUKNhfsUsPCT4gOQw1mRUsmv+IdKd7gpmCrdQz08BsgC2gHDx4Y4ZUDuacI
sFvBj+0crRCzfxAzECFAHrGhdjZ6RVWTX1vcsNhTf/i9QkXImNHidHggE4ua4gYvy/hX3zxA4VsU
/KteWG+EhaA9r/1ZUA+gmX6MUB9cj7h3DTgenIKkqUqUxcFnwyQBZODfwh4VCupZLScPLqqTCjrY
v2NoETfyMgpon1ZGhzlHG7RYv8gCMUGonOTnJAvUpbNB+TTdmwDoWVyLKjhfrpBowgka3fT7Whca
I+Gf9cTtpnE4E2gXBUn8jT4QXeXiphO0AlhnSBuRxtA4JVO6433bKGH/BYf4EfJGNoJSFqzfrYM5
zikUF81Gak7g2A367I3LkvlPZD46umI2q8df4vYm0Xr+b99zRQ1QjqUUp0hOTZV3DnWV4BlGb7oK
EHT8j/K/FoeBZLiC0qJOfkjp4qs9CkHSBTf2sARuaB3qx4R4tv3pJi92YFgPD/PIlAH1WmCTtbwA
UjgrVXF3u5XOcV8pCHXjQ/FgFAKNlE43Y4JbRub0oC1xlTl8lS5YUR7xNX6pEyvUR/4Gn4h7bzMK
TbsyP054qYN+xl4DUmwdMGlI+n8aLurpFikkRsloSkwc4ZDu8gWOUopWGCyLnlxe5ov8IAPHwyjI
Dh15Z/C0DlUK9DSs1vvH8qvuPdH5rFRwYG8r3+DC6rXmEVjdJyF2kScRRZo4bCwu4t/Re0YhT2Mm
iHUYOpxabS6YdMNz56paV+jAQe6ag2n2UpbQO53sn+lWcYcDjWks0Cz6tQhRm6rX7bkbjGRsWJ9i
VBQZum3mjGJfd66GbxUMYuK8SCoWHi+hPNuWIRKGNKVnqRBZMu1Rog0yEnxz3MbvjB3CShcqsO8N
KwZKkONpguYcmeruqqdRVWiadR9VFyie8urFUDpRbBlu0BjoUsiaN4YJPairLQqfftq2B+DLM2X3
YtRQsC36J6xaDckmD+F8e1ErIAxscdvhTMx+hfl+r0EU33AZDCsxx1pKIJqbrTDqHW7Ct9RxUK8T
s0wXXdCW88fIK0SJQKOu5TcaAIDpvINQcMdQ72+CcltFNUq7X4YCDEK3dWn/ah0Y89+vsyhYlOSd
EjFJs966QJ+kdUavmQ1EZAapEC0saRL0pauxINQXotaNXxGB//8f9pbRQ3YYWf3XOH/ZKynmcanD
nXVDT+8T1KMNWcKFm3LQCmkOjYye/8KFwQxirQ6mqmtvsdoc1H+o0TUVOi25wASgzRt0dUYTdjXo
TJbgiyYyY12Emwqq+HdCoxw7liNyeCD4Wfi+iPPGxwkjtJ9Kp2NisRBG/3CB8MPJx7zF7eB7Vl9d
25EvbeWGAz5BqbsVOA6jL5UUQ3pTLq/CRcGXasO0g/dpN0cf7b6l7atOprB/AZRBBAmNq+3NrilB
IbwO0pnJWSO0/GZQ465F73Vlgt1+P/JOXA8eRvaXlGi1wadmpQ8gm+gtqa0Ssp0TVNZyQP8UVxEW
X63b4U8aDH+GGGQH1kVwdovRCAwvlUjtr7bVPhWcQyBpaQrYE5QQV+RFngIXfixvh6JpTYL/HlUY
QMs8c4uaJTm2bAS9AWG+L5YIRO+s1SWPBPpJS9KqpbdxhRaAT/2VzurKJLK02nK7CDxdsVIWPbR2
yMMHInjJf87blOk76P019IL17co812iH3YIFi0jRkdibYWGKhYLtypals48+kA2mqSQeYDrcKZ8c
EI/WgwBkfCzUUXOn8BaED1u3IsB8vY0pRQSkk3qnZtGdTge1OZL9etSV8bgVpgixLidBQR7NIftr
LnpR2yZ/BbBujAyJ93YG+/XZU/Yj/epnnXd7nLi6kIMH3FkBtxJU7P70Mld48834+WPORFojXGge
GhHBvQyBoKYJehYSnEqP2ysFfdGRdhk0xZVwot3bWeeLV+LT/H95mKuplMK+RkNOk4wjV1hE/fOy
ZBb4O30xlcY1wJHvFGqHuYgyKA3ILNOaDFjvRBsKOGcqR7cwHWKcL2B86gjSusombEjwN8EUbs71
R2fpiFLL8j8JKdlIpMjg8jysXy5a8iAuznK/QVk/oriCYKUWc5QPNiNWX4KbA9f8DhGuor1WdoKq
SnHHRs85258HPGCTfa6IqG4af3I7JaNOuXoqxp+L33Rcn0tmtRY6FPZFXu/D3T9Urb1L2A8woN7z
GPHXmyXh2Q9exCTyMdG2hOhCn4dNFZwF3AJQRpxAUw2HJNoD8dNw/jlf06A1cDV1QTgEeHTurvss
9ZILAjuopGEqiuxf1iaYTdd5J8dQ020e5ndDuEkaDN8/OVJYE3U//CQ/c9WoqsbMBxFpnPC2pb4V
9MOL6G+K2jAxfHupQyeScuRBb9qFCbg7e/vpqt0+EUpSAYWYYdmdXA9+fFOtUn5FP8v3jYTnWY4F
vC/Jg8M4MeozNs1xbS7aAQM3+N/QkCdNHF9ZtCAsZ2to3T94eikUTDNXlCslsx5rH/LSgUpNvGU/
ZJc9XLb54GichQAcXBZDQlGxAloVRT4eNdGP3fYSRxikqheq3j2qDch0xaDEPvPxquwIHLFZqOkj
PS/pCUwEjVfI7NfNriyevN2xqG4FdQJXT4vIA+IwWN9ITbRAA9zwVDp2F4/jbohN/+k7iqY7Dia8
woe9K1/RT0mkZlxdRHx6HeMOQYbN+uoZQupB0DKP4ssB6sGiAJWrg9+DuhUNlobZvTf4LyrNsGUU
iCeSiPCMny+vYxu7a2qQ8kTFP9f9pb4gzB4GIH/v6HupybKlWSICW+UWL5AdLGhgJMDCAA3SpV5w
XK64HRvaVKU0fe/zLJ1S++pDCx57H/QviI8Lz6izgaOQjyicaixnHeCGbY4ExZoMg/Vua2Wl7C/I
dkQxtfJdhSeQ812CaTU7kfrinsuwxIBS066iYBavyOhWmjs/6rU1ZJD+/mAJ+pT3bi5R66a7VRa9
N3lFltzmT7OnVKnxYBV1J5lROcLNceDhNYFIFeUBLp8zRQH4Z5ScYCXa1YxADA/WEIEfBfFRN82G
9p6nt6Ri27TMf3fayKRFJ0RdLfarY8cJ1MR71CIT33bqPiezBw6ODRC0T8ZJYg8KlRTb7mzH4dYK
O5in6FUSqRDqBCSrH0NdyuuM4Pm5cMT3SwzHihJwTUxid0kgNSMyQZwG2V0CLfgbmwsoPlsEviha
JOa+CUwKqYKEoudCGwWzU55pBwbBI6XiR9yGotiBQuFIa8t6ifOz68kmCcKNzjUf591I4zvS0oeu
KLWxcXqtyxKPOlWJsaPZcP4mdp/s9GEol87lyOZ9+kYam4xL6q6K5oLHWIiExdqFCfALQRZR0/It
hsKChGjOjQjSg3NZUH/nojq31e1nc1QNeL7OLhGJxEYeEQghVBj1HZoJv/4676o12XpqGeZ+titQ
h4QzNdC19V/2133hni5D/++1eUCo9gcqId0CYKr4s5zQNMOO1MtEEDMVsI4O+Px7obg/Lj6MXTQU
39AvSpB1N//yXLoPU46IwID+yFSjKt2pzL3Ywuj5iu2wilBnTXyOC7KaY2JNQMSFPPhQsayH+VAQ
N0FhJHRx7/UxW+e2Wl0yAcGxDCDeOH6bdMfDgWvnbsAgn7WrmWY+chpH0bLDV93+bRY7mWJQUWqz
p6EzcJshVRzCnCT5u7H8VKPhnL1S6J+wYstFD40g9uEzIRu5nj1FW+30at48ZnYOV3GGmyf+Og+S
PVjTZUXoH1pq2TF6K7G7mCAf8DEWcDpPHXEgtL+wvTJhooD7hsd9Yb0vFb6mDuprmb2g+pV0LEca
w4Rrw/g2dpWL3lNYmTI9xHgTbaigAowHNk107nq5MytpwUMeOsmXMrFq/weV+Zx9JU+N1t0Z8Jt4
42Np1QAdh6Qr2GYhir4pbKxmw+uQL7z2tDuP+p5/JoNwflBVFpwcdxBEpEYwLdj0JJsPdWiG/cvS
G8IkXD+Zh8EQXPyCzQEqP/UImgAPhh3A51Vk/gHnasMUfxGCux8VLYLIJMzJ55bVYsB++yxMxD+A
kcubfNbPwE3xhdFkKsUNzPpI+iTJsU0xHRJGOjx3c6dlrAQElhr0GJLxXCb35hi9U8PvmIpmbRpk
Mq8JVUShQPDfkCgqNV7EpeC5Sl9t7DlUMYtvWRkPm2m82Qf653AkqI1o0UeJLv7XIlkArCyMx/gl
8PUv2h9FjJMQjjtt8I5mTJyfERtbRIuykKJTfJ3V8dpm34WCvrSfefSevH8rIsaNS45Z0Itc4QEi
kZiHetr+TLaUw+y/vK54SPPLz1l9sBEvCidkTDph+aQJuKpbfxakuf95hNKq7SkcQsskcK8V4PJe
WcH0NgvTLj5wZnyVW92VCia7E09uhuXx++9wWKNSHM/LRGffQZ/BY55Ra5pRahLFDgZNlsNJdT5G
SRliDms0IvWbMwLYRt38X1n4eAVSmkx90Y4zC+xPShOkPcjmkXR4d9dLe3kmMiCNngKEOsgwT19V
5Unv6rfQmUPulaUcqVXs9ikIPukQ+2rt2nlhWk8JUzg1U58/LBP8YCeLzB5g1DHIBAiNnlXJoCz1
PKiAAZ1TdoxCyLbQDVGK8kQ/xqqls9NzovvQci8QjsNRNUx7RFz40iF3xUfXHBVW7ZoWaz2ji+DY
1wvqXR5mU5WtVcBXSrMfMAgkJw2QRsg5AqpoVmQ1pUG00LBS8EsG0Djr9WhAOoF3zSTCd+fy8F2d
dSDkDxkvVXL5GPmkCnlcn3YdwLjVinDk81mW2QlQCZDg666iZJ5bQzgE27F8E2IesBE/meewngGP
wdpiJUMY8XzvHqZkXBiJlGbV3odDw/snYtNA6x9dDS1pPj/0VzKH0s8M1sT6uZMlycBbdKSpywj5
01RgPu4UQZ/n8GoTpKrsKVnTL70rF9IWEIXcuI6pmxFsCDddy8U35lb+yRvFu1qEmpoN+1ITn+Jy
peKJyLEeUg7hKv4H5shse51jTD3GLFWtNmM6MZTE+PBvT+gZwGArxlx3J178kW4ve+eaK/863oLw
6UH8qA/AefG98eL3hyyvDjE0gw4k900mvWnHsu9eEmNr19KREvutm6jBJfHwCxE+5/NU5UyBGoCo
24GXEdhDC6ooEfW+8KMQU3irTV8S8wzqsz1ip/sLwhEgrmMacpnvurfcpK5AarmDb6Xp3M3G48jz
ONt1S435rqCMK1Ml9spq1cZ/CoQAQtCeaBRmKVIW+MwLwTxDS4Di5iW8EX7arYzZS13Kri6/GYyb
6Qiv+AX3POxyINxShzY9F3dApgWzvPpDzpI0F+WR+yk9+dYDmwNAJR2BJiOBa3294/766CIe4688
WZ6FuYuIN60Fjs/pv4UBJDgkqMYJ7BmRO6HmohZH/Jrbyh07kmkAXFc0lq/BhJCCQ3aK/3h2sYMF
g9OnMLZUYcDRxWnL0K1JURG1UpyXTMp14BYVHJqUImebKS9CfBsdGozSpyB6pt20buU+i+0Ie+Vk
///nmEoH/ZXigSsko7kp5vQAI+V9nTF7wtCXgkusDAtuIjWE7vRQJB6AiRyVssqeVu5d0T0CQcIq
/ToNeIiAU0ulJHI8GMF1tNJSB7fB1ocQFj3uaTYfUL1O/1oSIhTy2Df/r0mZpaicel5RD2iUDF5k
D+8vWHuggMh8nIe7xLqGhA+zvklrXcyUASjKiHPan1P/HEJx8ZGPw2Ya4aj4Mty74oJ3aAhpYJCy
pianUYgDJdBFCn+YnL1KUoXS7ed403ygjRooCBc5SOmB9SZ6C4IEc3l2wnWByhddos0ycmLMe0z+
oBg4pgGfKrDPFvUDVMmGcP8uMDTKBnVzZ/HEf9mNb53D45OxSqF9m7FzfNZsft5Pd/jGTz8Hz4MX
fu3W4EkZX16XtzOxALKLb9Xa9y1ljZNjc94qfbAzOSCGhV3schbBgM5hyfR8M0mSpnF8xLM2TtN7
d0uviM5kSlWcCDEfdVHkuO3ELsNoPoV8OFR1ML70qf9V6F2vZ1c/xpkwI31xafdbLRTO9sQyQNvp
5EQCkXDpVW4sC41KrOQ9NrDdw3iToYbHKiR9xAmOXP47E7Ch5fHDIwZinEDtPgDmY02j3SoNA4RM
eiEyIFToy2oM2K2tZuVi9cfnRFVep6Q7k9V+mwvQu/LZaLSRDGgS8aI/w3FlzQJNS3Sy/cB8SWLM
TzIXCRvkEPhurepLqjomdIaDw58VxQdeYkdJmPwssZyiExly9nsDiNsqBHbRaaYZCryd0XupqXeA
nkbfwL1Rl7e70OgdtUN3o/YQO2vwsRXiHJrUrLSQ+n7F5KHLRAbjGc4yrHOuq1a6knChnnhodWG5
UybGovSxYGe2AVa0gzTjQTnECuftuq+0fytBnDPp/nzA5JymC6golQMpni19LolfmzRz/P/fzl8I
x73nXv0sznWPUcA5rWil+Xn+eF4EkFAfCsDdcrrd3nh9qxIwdesr+TDz8JToUH1xousZ7MmxrNxn
rfNlPnZklHtOlc1ZIUs/dNSi0js9q1s3dvctBaANXkJiApycklauKlvsLiRj6moykMApo72ea6Ux
++Ue6e+ziQpWPvbavrw8ZyeYcx0saLCNzXMI0eDnYaybEQlEqdpHS66jukqttBglN8jE+VrTFsXv
iJcCKKA8QMhAucKLqzwQha1GNVFo0vxOsA3zrmkwl7C0rQ/Uh85+vCBDSow8vMrGUqWD4mtxUwT3
QnLd6+F7KDIQ7vPcKAPzy7UdzJCqoz59jQY1uQB/ozeUclRQq22NTZArco1ZbxeKkhQrn2falW38
ooHyN3DjR10o6HWT1tFm3vz8009KdoGSKR+C29X6hKr1ak6KP3bVl3MFH0eH6xHmRjR8FQITFd6t
TUG7IjpZz/0kTUY/VSQ/z3mZi0lpxAO0IE97KlAIaQY/ymSGmwRSCVVO8sGEsOmNjKWSFshTd1TJ
frKqJwueCUlKf0+zyYdRHWU76sVexIZ5azOY4tZPPPx4M733di/5oSvGW2vTTjEK0PAYk1Q22exZ
I+DfAijRER//LU/KWnOlGpHbC3FHbscJ/7jmQUTuABvhXWfMcZgwlJZNZeRcCDHR8Efqz360oaVq
fbxxJqZhlPzjuJxa2GTRM4EB0TQerQeOlOTOnq5zktrpdjyEVq+KZ4yhbC27PYCn5h55ty3oAZoW
i/jIkoCwkgM0ww1ruCFbgTe9kM4CRHcd9gnwIc+JpYZd6fgleXreHHLtwq46/exHyl9JfVtzepcO
FPyxf2nJY/+zSSFEK9XDtHrBjHBClEbBWBi1zsZfNWnsp0w8MmrMwczmU200Cz2H7gwYoxhdIxOv
yzDVYTRSlsBckeFz7/H1yq3w0zdXggEMJYztUf3+g6aFSfGV0XZm8ZaldZFM96R+CHP1e16za6CR
XUQlbJanbWpg5b1CjU/rEo7GtjdknB+m/4twNO5A8ME11Fuo3JngCjs2xGClGc+jI1gpw17FPj1M
B+ONr7/MpI4vulh5jVj9xTkCywXLD3msPl2qItlstdhECByF9Jh0Ts8JPvAF0gruKRHTheTlDiT0
M5fn7/otd30FLj38QSvabsnavnS9ghL6PF0qqU4d4W2ypblTt8emHkaA0Fypa2I3oe+iImjIeJzm
jm9990qf//orfDotOcD+2C4cSjZ5+unn7FXapwvkb61At09XRtwNs+jBf+n1ucyCzSCx/HdJ87AK
CTBmx7YQiroGBsuSOJZP+DJ1NxtPFT83mWSt9wPP8QXzAk16Go4jK6Qc+5InbtQpuhgueoD64tST
MG1D/pYabjqlxi+ASncGFicWsDQVDGdYPFqszbBq0Osj8QbJmKCYK/MYBmqORjPiidwzFkGYOynp
A+WiHtnJ061qI6Jc/VHXMz7Bsgb8Dhkkn+zeWBpETBDon09awoSub+jhK2KpkEhpTMAtxnYR5+//
U/6WnbIf+hDURxGx+TjLbbgHnPXMo6Wud+AIRUMJdblFkRyPhU6neH4WxknMidVIdKVH7fOQbwCd
Q16QDu2TdWm6+MzRaBFVs+aeVcwacqCONtjS2o1zjzDQEniL5NIQlG17okUPd/RZKnShs+x7TKTS
O7Rtp2z7BxWTcGX/Nm1IY3I0onHIXa//7lgpOOfcVblK73DGQdD5ms9hQN2L5gwcAOXSZ0eqbxKW
S4UDok6F/lMU2fpDOSG/FHsMb2M6JNmCyyG+/083UT9ZlD1V/R1faMEpVWqyDWvOr9jp4FDFoK0t
Db64rxJFH6u/bjrvvcUU807q6x1VgNNdycfLdPKKkLKbtOeGyqIq56GZlOTiLR71xOukJ+mJmRej
azVyFgSuKUMjPanwxBFq0TTdZ3JWiLYxIIZ7Zl716wQg/trFY2JeVvaU++q2sWt/d3Px/GYpUijx
HI7QQjxTI0X/uvky+/FC6vzoYdQtDl2MtuPGQxoNZdfeZOPWwj2/vUXZZXJWfM9Y8JVeOxaApNA7
FCegqt8Po/pn1v9JjD+aylQ0/1cUdf216FbWgQPFOt552QohgOP8LD+6ww2qkgKQ9Gz3VXktU6g9
hXQVy9v0YzPl/psKSGDkIyOrgYM84ZWDSwoEeYyhD0AQAiEUovtD3VFswwJbRdfP++s/WgMjVn1w
O2NUv+Uoheczy8o61NlPlAg/i/BrDsCvV78NqMmEZYii/aDT2GN+p0zbmhG0rppFPjtz9f5+g9hQ
sYlgq95oEOdvhx2U/cUicHZEdOpJYTqub80PlBEgACmqKGNUFyJOfNa9PmAvyMuj/HUAbH2Xq/JI
rGjz0jmkoQtkcp8CAhZy5QRue2KKuwmTc6Sa7Fwas557FmKm3J6dZb/skvhEclSjFH3bQ7aZ4dZ1
u2xRzlm/bCtuLHGuriutx/3g6UgSwjgCN2HfCBTiMdbuQOvz5VSoenbHEbRixX8fW/Jem5I/2EL3
ftHNWgqjeH7C2oUg+Ce0sfaKMuH8ImSMa8oEj9zX2Mtoc1yyLxBshlGK1P8jKtOSkX0u+2+gOA1W
OC2F/p16AMblnMbgDrod3ttphgqxIu48O0+ZX5c+QBluS0CUtX0Q8jAh4rStDUV3y6JH69kQ/ZQF
8EFbir344YfWlMnpPILVRT+iVv4hNpBRRpUcLmHiETceKo1hUyPEy0Kf7FWiLX3PIrk3i3L3sgjX
4zp/tcPvSF9BoUdA+XYZoDV8HLveaKtoKckaWLBGsf1CT2z8D5blYs9ZUfT3IQEYdiSIyPAGGsVF
iIMzQ6xo+ucSZ9so63JHO0kzp0cULTM4K+gTuS4E1zPellRqoE0U/02/ljzLeRPGy3Wp6E8o9mW5
wEAkfjm8ATqn8n144Gewbyc3HfY54wX/fy3F0mkoFO7xURU0ZrMaicAVVZonGiA2zd/W2fgYKyh+
A9b7L3ksR0ZMJYNMy5zgJHiKGyJZmj2SCkZW841p7Jn1iRr1qAznhqfaB+nUZG7wki17WF/WsB0+
O2EYAjn+T8RNyfragsYypQXu+VQLHy6W1D7RluMdJ2Y+pT3RFSrg0ajmag/B7sR1fqaBBeYHijhZ
LsOKaOp/WJ3CGoUK0bfliYW7xuvUWi5Uu6Jztlvos4ZWGzWHkuBVucXt9cvEZv4JQoPxk3Hd0B2t
mswxGATXhX6YsOilwQN5EHt3ssVHK2H9GCvuKzI9nBAFaTo2B/+Xkpn0q5QxRAsq8eRWer0myfK3
9+RFKTfvQzGsjZJBdcFG/yZKRXOeP2nfsOo2E8p8e05B4PlaVOnPV/LQG5dGL0RZPEVqKx79ErOR
gQqejEZzGoxJqhKtus721FhcpCFiFD5C4hrRHTMbFioNnsutjOrNYhVt60Uq5gf7+/mHGG2rXz8Z
6UciAvzEbO/HtBYn2N2HDgbVhdrv1fLVnHhes3cwQzCzTLS6E8977a1jPkTVbwlTd4axDHt5JiY9
tY+Lrqb1MBwGVUfKfbkSQsKYv10BvDWlpcyBXDuC+i3d161GE4VGjwsZ5HCqD+gnQShlLc2yhmb9
WJhZQgZAGyeMwgOfcl0eZXZz479zcJOqd78k2TzTurSeycbiObeJ5hncFV7W5YzIa3XEc+j0klcU
Na9i0zSz77beihnuaq1eLw3Jdvl+2nTu9uvKPfXv1JlRsoBavK8dLkw4YGzMNgPXD5iVUI0dYFnb
xuAoERFX2vtPBUteJclTU/CTpiN/RW0oxuwV7D/dHckJDZ11eMhifdmiLGgBmB9ydyliWAN5roNs
n0+jxlb53WfykKHcIZewDluCVG2Tvg666uOLwEDT/R18iJR1oe2FUsdn9CBcYeK7Dd58SCf2br8M
PYaTWH0N3x9XkZdltyzdui27BW5SviGQKn7KAVoybOiqSEYAFsgK4ow2FcnGrRYPTqbUAJIqfWux
H2dNdIiwCip5gAOoy3V6OyVKYb2GYUJ3A0zl2ms2wEXjjiVqSCp4icE0QHwSdCTT1sRdDU9WosCF
COrKTWd9u1rc4qjiihMG0v/tq27RwYTxudjKXFBir6F2Ogv40UitY8jzKpy2XBi66zbITVSZrs3B
UeQOo5g3/n7EqCTxxx0fXgqFGH1uujxH8PblMud9PDcLgCbKuYDVdOEK1n+4eSqZBw8f21rCKoWv
dhZkLr3H5FGNqDcwcdmkWG7VLjwfqlRzNFckBEcJxnD+LgEF+xc7i00SmpEtuxz4qU8WcB/eZtfx
EfRb8A8G3VPX4TP6N/LplbJJ1Sdseo8foBNCr5mx13ZvNbxHE8wfFxMTcs+YzTMAQRBVydQmHrt6
0mCjORe6gDoE/lGGoHKBx0rWo8a7C+Ix3F+d/Hc3RVj0azfGURM3VzUo6nUSUfNz2JYj2DzYfiOQ
s/5Wl0LUINGZEr9BcNfNJNJBvC6nfej5qancvY5rN2gt0bp1zFVx62glfOIepuf213hRQffgQCil
qbinAUT7ZFSWaIXnvlyULg2hTO/h2Ox5vyyK4ddxCOvaKHMFQvMRewXQwSiqccmLbrQZ7XnAHF5/
o3xshvTyQtkVgotLOASN58geEdw9xEdbBcgO6oL62totonENp+LsKRS2KqNNvliZoe5jEPc6Pjq2
xMUACY4e5Dr+Z40M51FU6uu5Pcz9YrrcyJOP4u7FE+G9+XpCMZ44/tTAl90rDBAN/rv59FnIMFbe
MmGdN9q9Mw6H5+/rpM+eRjHWcuXM4IAoIwhGDY+U9VLkqNDU5bnEQ0tQdr4Lf9TYj1W8KS83HMKG
84vqhoq9OtBNRDTE8VlaGOk8G3xidUYaOvkrZ9d9AT9Nbrmhf7kpnz6moj9O2nu/dgjpPoR1SyIU
1FUR41rB16aNvs8YUfF0XxLeNanEfJs18aSt/xz2s8lQvvUF4qq4VcSfI6EuE08O3KGUXNh69/WA
cm4EajWyp4QUKJQvsZd7szncHtRAopOnxhCY+oflI/kZFmvRnsq7ygrhSJqzQTQiu8AQYq5wFMn/
CJfc9nKx/nPX5SCt49RQWm/LRSjssQg+1TwqGZnheFIBCG08o++i49btW21k+WdiaM6nX5M/w6vu
1s0eZHK1wehuBZqgV4wWvJX7ONJOlevN3V+3ONqF64gPBPO/jfYu1hgDIywQocNF6mk7i6I7aapt
qJOFO+QSZ+1RPBNvdTz02gYtobe2RSpCtzimgpmnKRwRCEvBS/YPNkYobOLlpvx94SX3Oc9zjnOP
D0yksyVTlXKYU1zWxKVUePblik0Mu1jOtbpp5RifmInVNEMVNb+cMhxEc1/zo0emBh4I6fYtQkrr
YaEgUxFYH4kQsIIlfpIlKdb3mTgPgcitFMiSZSq4jvi5pcynUJ+4thQGiwdL7QVSxT3U0GWyzS+A
7KlTiW4HcgwQou9031GFIyF8e8yahls5yHy69UveA+LwxqwUUCaS5GByW/gc8hxXpePRCLc2PN1i
4cAT8gAThcro9i9rDbJufQ3OVtKIMmdyIEXGdysfVKtzY9t8U1du8ujyKSs43mJxPJZfXA9KwDVx
3VW8DD6Nj/k4EahEzfypx1z/kglP1hfhHnO9dUAz9XcoMyUZ3ZkV7zTtlYkOoF61Up40nPPKu4nZ
VzZ8Unrtm7uuxwJTF4GSpqsFpSiZ8UMEO3GJ8AYiCyTyH0gYkkfey/pwWsIQPJRxB5Zlyb96Ngqe
WGDxnkO4WUgC3gtdX9X8C4RzScW3wMd+gimcejW2EqhZNT8hz5Dc+ZaR6tdOfSx23Nf2CrbUGuck
VvKx/JCzlntWb6cRUO3S0fOtNfaRvbaxXfDITC+urgdI1ILzf+xtbuIVhRyuSCCdrDTazfPxb108
VHa+B9PfgCv3ESC/l19xhhWBFxZTu9NPjD7e+CF6CMduZ6LYiQB12MkvCrOADlC8Usb1Ohp9jQIS
bdOEpgYgaLjGm2lH0V4sHVz6nVgOL3Bpq1NZJ38ZaWlX1PGJhUf9X78eYSDErhGU9wyNw2Jb+cXf
6zvTgIa9eXwrII//J4fIpTkfaj11J61T1J62zthgKqU2BGVyjPaDZJ9piuYdFmoztfoM8JN4aTiL
s+wkvjOCB9efqhfZ2jIXpRuwwKkeDB/AJbCvM9Y1y9muRpFqP5N8jE5wwZTsTpEnOqoDfMnIl1yG
ub7x98SyG1JGuPUJ5xj+lOLXz2tu8fNDTapIYu3wqrvXYnW6E4e4mG0rLFqqvWbe5qlyX2CTSBuH
eAfs+QFpnchfnVlin8FIX/yr6hL+jqb0gU5cy9pgtNDmXpLad5/+TEhk/xNZdOYGJwpD1JSkW+qk
gvQVtnEIU7z2XYHP8dqI+w/hyZ15nLICCDjiEWv+3CIFTDCvyiTIHPkfpmLnPZmTZtAILT2O11fY
tHMnC3C0F1BktsgkKRDFev9eG0recmyxuPfodXKOrwRg5MNsEKDI//1jh4hsi0eeBl6Q46jrCLLb
XhuHKbxqojktby5/BJhUrLL1L/z2w1DwrfaruQsrScjy7UiFK7w05Cc2MJaIHXbD2WoFHyT42Bkj
lDVvhIW5L9m+Y+aX6XmIs0Tu1R3oXe7wH8uSQ3MD2q8rE+8kRKmtoOTHml9AF4PEFePY9peHlnJ5
kpIM9ERXNZ53zm6zu/xA2cptNqsYVMqFZnVBlELwgTvsSt23B9kJ8KGvANzryy5G+687gfjlfI8R
I7lY03sqZoaWIoWdNJc7yS0Zm+tpVawy9Py4xPNDNvAjH4DdxG8YgcGWqb+U3+M5bNT/OM5HcJWL
pIBOjxaWjREMk5OObTn2F0NMNZ9lXj9+q5ICFLJzva9bUy8Mevnh8lAYaCLtytHYqH5Svz/JamJK
0IlpU5Js46GOmHfke1KLKscTlzupJqlL56Bt85SYrV5zS7BQ7Q7T5cM57JtXukETQYBJgxG/oksd
HxBJWcFWrMxB9G1GcaRjVio6g2zsn4V8M7wptLqyzuYew2+eTyC7dTvFQLTb8uBHEHFP+CYL1WWW
jVW7IdbktqcmGYhBcbf2nccnYbRs62RMGHf4blPxGvV6hbAV2l4Y4UbocP3oxz8YAxdMWQ12zGms
IEHjp3lxstsvGrZORZ7ZKKP/OgChYTC1CU2GP+JIzrw91heqLOsyXmG/t9Z5Pl/yNtfozm8i7H4X
n0CY6Ctg0Q8dICXr/PX+ZgGksvpNKGTf4YHM6x+PjrIRrH+x8acEX8zSPXLaEyOXaH58uiaC//zD
DwRl24RUjd8ahSjuR/AAOrgmV9WmslRrl/VkX96uWdAcGJkpLfeOywDBTWPnf+X7CFeIw9FXLksE
0q8O7SN4555mJa/ahJpkHyJ20BdOFkiB7bn8YnEwCcgLk3AeO6+UQFGYPf7UnlCCo5j28bgIQy/w
xjto5Ra2eY/4ayczkCPVuIDEd7KIi7wZ/ovi4wNC07InvauC2cAxShim+Cci5Tww2N/TZu/lDgXY
CaBVZ7Wr5yRAa0VD43eNSPmicUrQpM/oBSfuzx7IUAvO/SBBBgIw8IJGLrbmg5qo/42y83K4hQ1m
uphjtDNpHHBSQMAHgLffXC8cCOYYPkXTmIkF8dHEMKI1E0S3eN/Gq6vkXh9cpLWVjE/mV/ePHwD4
46bGzRHEUMv8QPexZAw4Pkrcxa5pUBO7VnMB7uP/XWjlvWOPiDZj+42KtTtXX8uBx05DBiP7NIQb
mmqZs/Y594nJK5PmHRJ6+zchjXisOSpSAF9dWcS8+NpurADyKE9Ku/wuMXX4O7I6QBQnoRReWmn/
/g5WFROijbw29m+GuyTprWxBNr2+0pyCZ19YIQ4v7iF9aL/MOQAGdL8laScuLNUDDUH10PGb0air
kt3eF9ngw6nJ1YODK1BfIHhqZD8dqIRX+0ye9hLwO6xUi+0JyqVRZXX6TEJlnGm+A8UpL+7s8HSx
YU06ml4Jv+iI/y9aRJrfOwnXSTNzQdxWFYQOzfR3hbY3zu5SxQ8uV2pcTgMz4bIqRV7/DJoW6qif
syT/MEe1YtsAmjYswhBgoJ8ozZLiDmyVOj2XKvvjH4/nn1QEJ1FXUKFjIYaBPOGgWF0qbPuWgp35
sgI1I2YxM+yfb1xZr5yb6XbD3mCNhssdCmm3BoozPlLTfYg543OqyhJE+oow0Rk6VbNTbFqevw6u
F4EvWtN1DVgTKi/UKKIOaHbLaWhOdKlxtjIZhW85m5Z0eQm9Va3APZDS0nHf5MJE0XK8LU4VmE+v
ctRYGun2rI89OaC9mSJW0yAQ+NQaRizhK+vwkU3TsVtzcJQdZV9DFzn1XXcwPoAnyTvBjaOI2urx
oKEhFSe6sbP9h+AuzyQF8YYl0forr6siN0PtBCFOKjN01EoWIL1ci0z7+NN+UrT4qJIHIpYe0ynd
CHJTnye8XhNY1/Ofi2FL6WZKzsy+olmufL8I3gTI449l37XfC4e3mjVaOdevSiOpvL4vxuY8zzcU
Rn1SmcfWspLRnFASTl4ERzFh0VYIiS0coNSCgEETWd1e0gUB1DhYK2R8EmKE341BTvltZTyxTxbK
vd7ueRuAN4eKlVLnTrJ/WfZ3MPB+QKkBY3BL0rL86h0aqCDZPAp4I8Avym+QuMdybFaD1PH5wj1d
nzNUwqmuJMR/W+vSjz1/X0XRX7kq3HZpobHdicp+eER/IOUICj9gNU5pqSKjVie2aNeklmZYgDZm
ZBNvpK9B7CIKIIuN2jYgxDa7yAnJ9BEGYrUS9j/CpvGbZs5DcTIiN1Sf6geWEpkgo5qz5757+417
nmHqEUqohJSxAIAsk7tEKiXZdOO4p3+3N0TyEv/SV4USjDjfYt1OQ6iBEvsjwXy4IiCeamDfX85u
ZWGfdbfpMD4Fr9ElneZprB/Xd64AkJ3ZeNi1JZzzATBvCtY1p8Zxv3ZKDCyotHP6t/wNvZbMtnOr
GTUZT2iuCYlE8lEYZmNkfZJ8WPspT9HEqpR9OF8gCxVxVocF8I8ep9UiG2hu6Hdk6IjhBloSDIGt
CLkev9sNsgVmvvG1rNvn1SbSz1F1lkR8hwaZsv546jYw+CEWgbHQttXeOBZHrqj4DDV83AATLvGB
U7h0rpgtd+SnGQ0nhMI9ywZ2LwnP9/lxFQGqMqYDqpUWBF2w0pA/3tkLKERaczI/DrABPMi+qquY
FlFG5BbjgyJ6iwdikflWDmFeUVyiIRWN9+ApeMfOapNfewGYVtzWSpDN4ieUex+Tz1/jNg3AOYei
2HZpA6mgPIDjWDt+1lcf5hArVoYe0ehSgkV+8L5rH7Ho7FSzkG4Mhxjbfk3E38+sJP6z38lrrNTe
YRbWy7lLrxQ3tUgg/wkugb7MCksjN8Mojp8PE0GP+HoqDaLkUbS2YSEOipnh6qpEMi0Exsv6L17e
F5uZSNoBuY0TnpMOspd2XwBemhkgsNRA9mZht+4yoPSW9Yz9IYxARPzKztUbgW42lLwtdDnTg5v5
xHVB3f3gLk+Ux0gRrdFaO1Rsy2Ys5Ev5kMNrUbvesadNjTKhsfab2GCJdySTABjqbVIs4epoQJD4
VbpmI4mqiWe0r0mVf3llB3uYoJMPxDcZm5U4oxnjYDFx1WbJlU6Ax+DADCqiaxoLbwjI9dU/sYD+
86cbkfYkbut/QD3uNfJYukfjX6cuvQ5FkNXTQk6nnsTBzeBbKMD/7IpstFQbwHJKPV55WrskXSl3
TbUexKkBKobnlMJtBp1EZojYDuod3/uenLH770nWjpj7fxmI6VRHkG5k30Xnq/0oD5xxBGlReUWI
7eLpv3a0xc2Q/2PMe74/sXumqWU5r6rJ0VCFEW/mfp+fm8oXr8q/W7S+/2QRaWquC+FxOBg7xHaC
3er7HqQwVe54qbi25gD1UWLu4wpWohrFxVrQ1J1tDJh02c6IgtBVHTOuhMTEEXkTINhrF50hlcgC
oWgvg9CGnmvZd4+HvzuYKITf9IkBzVxeiTsT/CV4ZxzWcrCUM/KS3e7MqM3oiZ2qe5xb+LeRzT9J
aPHMiXcAqLzPcr8FupTxQkQV3+biU3DyO+ZTA+TdZONRG8QJPEIb7szogaNeH3YNsJ/FLR6oEG52
wMgZCfobKjO5jI1pY/6H9rUUT4FaTUbijdhW4ef6BLoOAkYW+xmq5Sb4CHxV8vBBG0kRxgKWVp8D
funEl2v4rfzytlIpXG0Dxan+EHNqs+5XRse8KdLKo/YWrusrGJcN1GmucEuYQxUuqfGSIsVrgeKR
qHfz+RIL4AnYFvuEDTxxpioInHR6TueBw56lSnPtAFtY9K2/iVomWJ+ZH2r5do97HOIz9D66oJj5
eh/BRJXft72puNo87EPRK61jRFk663J0o/eamv8QFdBBkyVHFfQe3CIu4PbxWtBatC0v8Zd7B/gE
tUYodQJI1Nkv1sDQYICYgu3Tub/edBnrOeuB0VFjPVtRvDQsXf4WSsX2iiDXQcBXu4uk2xu1S8mh
ygA2yrLPhv+du15N2wTi0KbPjojA4/QQEtp4kudGwYbGDDE+J/tImZYYYFtl3iWTRfltzz8K1Ubo
P3Cms8l+RBNe3tLvYM9C0Zn3LrTjk+8GD0PrL++pCxlMfsjzqyEo8DwHAFt0i608ERnzX+DbAimv
/YESRmd3Xq0lDShve1KyTJzueSbjT1uI65tfoEX30t7Y5cLIoH/4Upw5WA+Qq+eGFCfRymfgKjEf
347AbT5WQ+xtVp7ipSZVjfXgjfLXbEDreuCnDZd/QSFOicSwHfOo1QpZGbMqRltzBQrqhcCnppJ2
3o7G0XQ2NXgL6CMKHXDypc0pVxFNMMU7ebqSZXcBoRE/ASKH050tO+enq+1vGERXgz7hB4fDLD3e
rdp0fvRgZT1ltsPmHoNNYwFYrmRyvL32fhAU8zIaAF+PUORMFadKVKHBBP+Imsdl37tEKEJ2HM0w
zRg0PEZsNIv1wLYP1N8r8b5oWvnZv2bAk49bxIvGt5L5fZjb6dzDysjTI80cKSbr2qW/DWbvke8m
7+7BY6u3x6U7CYFQIhJRgw2NkNgeP3SHApI0aG8Cg0aT5NCQ6y8z6FiL8EZhJlDdZTApHcuYtn03
xwiPrsAqMgm7D31xTE+zOp/Ok0Hmn9/KpJpNTZJdsKaYFtx7eo5VlkKgSna1Wb6kEv+p2OJ3PYzm
waCmPni74ZYgfLRPnHQryXIezmAZEExKzxqgUB2Ebe6mgsCfD+jS9V5rexzKfad3JKk/xJ4kniA7
UK2HYas/JqVBggFd+DS4LQ1y1T3Dy3SUPpcmR4NgrYp8EyzwwQA35IQzbV9+YIayNSdhSFIJ5Qxp
6cpgkDiZQlCeZhMyUqrWXZoCzE7uKj5C96OXFjR9Wy4aGiYKkXERqbzjCX1XXYyaKKJnPKjpN1jv
BIJTB491r25x9C3ejssihZOa7y8UODltcjF+UZKgOMMlnObkBVsWXdGtdjxfr7m7Wgzu5GvKF6KZ
pdizORtQfGgcrjS2h3oG3qGoceBf4HD7PdHA3GFOg2hFQ//8UjOC26TNWtZaq8zR33Il+vISEb3Y
9S5ZvU/xCnPAuQnXxdgDPQjHgNtdpl3SHratuIUhJg3NN5qh4Obynjh8zkGYL9FLOH0DVUBuMsGw
pgeigxLr5FOGJ9h8xhKLJDgFXHHnWLFn2jT3pMEbjKqqynv2naDZsoI3gOm45zqHfv71oBJRUXOt
B+zUyGm/3RkcJLhBWk8QQcCZ2YMvoZyvF18Oq8Tyf+2O8MpfYuOPE2jYgBB8N5sRuVn/I8dgDRS0
pKGsa1EASIe9fb5RC8tsXTvQQOrHkRKbVCbxVW6EWjM86hdOR2ETb5b/zWCH+jguL4ennCUggH8B
xqx4jFJSrOlqsvWfoiF9ufnh1DIussJwWWDSym5C7NMNiwePIv8yAKkGjcfioPg/Keyr+Hk1d89n
hW1FHtHZXMiQPDPEcXIZqOYleez5Lc59odSKOjT83Xx9yEkRfFEbAjkeSel3cKk3kt8OO0ccKVJJ
63J2s/ITkPHC3Wy6P9rXT6D4ye6DEMNSTAGYkt/maivdTr/z1NDxgBeXLqqZPpumQoRQ+hExjlmx
QQKgPujJlC84Pg2/bVm9ZepB2zVaMMJzzfFpj+Dlm4WshAuAwD2LKeVI9K2KK8D8uXHwDrQXwE+q
DaPcofZYlFIUUq/VDMLGHnegWp4XSYJdmJXGh++ksbz4uQu2c68BEN5V/g8kiMafS9/YqSXj0TCg
H74CAUIHajhsf5XJOpiIIJAH6+MOQbncANmzOJRp1nonz/FIReVggZIpgWZRqUlfuX3weKTOgORo
GCBWVP10alc/zZaPT+4DR38EjqcK2AJIsOVjVPgRpgWNPb8TNfUKH6J5JyQA0ETHlUEKV5O3rwp1
MlPzdxaBKPlZeG3ctJ9oD2QjJoubYR+oaBRWOW3hBPNEH8HzgGMGjiN5fruT/zVaAfasakpqWIUS
bT5FcG+YDojaPSteyvNCPxmDX73unRfPCGQsAt0BAuGSNqWS8ef4ranMmTV6Bpd/a9YT9ELzvege
BVKWjf14UBqpOpEvLPIJzJKE6Gr+xbRKAHaerB73BbpQ6cCplM6xgdeDze79QicS3rh0NcYtdZzp
YMj9YIRBcdmK2Fg6uzpboKOq8LYNfQk+34i+1vuMJ4ZC4nYM8wH0Fzm22c33oOH1O0FRz0JYaE5W
NoahGWLhCywB6RurFI2Rf0ncPEQJknysmRKjPXP3hQeSxUoKJa33Bu9g5G6cPteyOOyNVROweAOr
4AQBhIxXgglmMNZFsr4DFHjIvw02t/kda5X1e4hYxI2Tn50KUJGHYCUMbRDqtlyCD2zQ0UgruCIn
ucMNyOqMyp0/Si3VOP6cT6MEabLfxRuqT4mby3cWpOA1a4JPty1YnU0L2Si1Dbc6xTv9Q2w/97kj
xdGyX8gqyNkkmKbP2VoqMmbNs+ZNxeWRlFdj83VSWB8b1QaWpjTC2pTes4H/NQOXqy7yhjDxH19W
MdHgWlYRcYzsTDP+dV/LSywbZl7jUqEVvXkwex+29+rOW+vdQVPbbigmOze/ZDJ6tZ/VtKk/agh8
NzMMWTY8zKqeDBpiG/q6ue6VZIXKJ0n4g8ISUyRLbqlSsiuVeRDlw8a9IGeOZfp1WbZh+B3yxKuB
NbLNx4O6FVzyxB15wD5D+/TP+cTaPUMZnNNrXmiJtft8QERlz0R7nntPeg+Sm0pswc0YTCUUwVpi
bxGj9dIe6ComWQIbEzmo+8QUl2yTT6f3LlccjHjNKjRhXEOiFX3cx5Pevy72/ZYHhzTffUtu9HMY
/y5qUVMSnNOcs9SzJsMhTNun1aAPNDn/uZ2/WVBujf7WQadsnaCb5GI+l8pT2NBAWL/T9Um+6sH2
TZ8Om0IrksO/JUn66z8jv2eAgMhzoli+yX0kpLLlRoUS5LM/kyL6Bvo/lvnvLF2mIJ+bfRn772II
T2RscTwo1/EFH+8UhAZgJAR04T7n8rEz2LzcgqudJ5e68S2pXc4rI5iAJV+9KfQNH2YFa7K0E3Au
U65QlguxknZJdVF6wP6+4LVxPfqbRn87dW02ctOD2JOqqJkPTxt+2n1LqRIPl2kNWc/htqyDXRKC
lZr4nyFPNSkF6b5ZRuYUZ0Vt65xDz3TgAGYAEwAAQcmZ6IuOL7UyY+tfLwGstZG1RRnZOibaX2gB
f8znTUNQCpLfLPBj9L4YiO/gbsQYM0zqhNFCCo9VVFOFOzOl1C8JKP0lhXXn4JKItV/jMYBmQqD5
LHJG5d528OmnS47x23gGFWfN1/NgoJt61qC9WmsFapEBevvwQcl0tQ0pDRAIiWljZLy7s3BaT9O/
mFyFVvaCelG93aXTLTL3J1wkfxcewKbbmcBoIib6ZajYH0fViHjVfupMDu/yFC/4WeA5Temwqy9l
JHGk/qNtCQdl9qsNkZd659g0bGcrMchxQqCE+tzEi0AerAXWBJi2SDKy9NcBcZOVJrYWZL+sLwCJ
+QO1qWVDQHK+XHa/+LlDUDbzYIsfBfBpBfsUq0lBw9qG3hr9QdKDaMZomLhZIRc9i5j3Sz1Hqpqt
BGm/q6xpL44o49tNSQaM86LdEQlv9vgSavSatfs5REUnqb0uPAoYKcjDNqUDpIS+O9KI/Em6+l4/
vleDFGRAq4CWGaV60dGEn93Bw2Pz02cRm0lrIIJjkmvu9mOEBJoTqrKo4TY6DxnNI9iY30DxItww
nJpB3mT1OHqemDrLTIbSG/wisqVm61ogiPSEYH2SHj1y950GaaU2nTF7sGjxcbVbiCiHQZ+v+Bxl
HniqbHc7JsEvJRh4yjY43WRAP40mD1BP7vIIOLudn4RFfhl3GSSUriRKdnRJ6W0fWcITwV0Aegch
aGsxfGHmZLe5z8MBci+pc0OJ+lYfMcoC6a6MNSV4VbJg8E+6rLezgCgFSQDRCYeK7eqY5szQyFVm
MhZCwL2L2Sbeq8YXf673vc09Of50/iRag08SH5xZiLEF3gKehJZRd6YDHfir1kNjmtUgu+NcQ4uX
PS1vIndjbzmRnBGUWBEdVSKq/aSG1l4beZ7D2WrOgFZGvnvbKH6hX71ec6lyF7eXcBNF90Xaky1F
chUhpVZV646zKwsiA5tyiVQ7i4J164Y3AYLcqPVcw7kDWmquNDTV1Isp/hda8f+qiuVzl2d1boc5
xtz5CM67QLdUFAjdD6+zImGQrdUMkdQrxQY8z3+DJYkLwgDgeRKqDnmRcK40ZAvdC5gLJWmj6Jsi
otKJm+tXwtsEnhLP8iQw99EguXna+GHUAlB9nxEDJ+CH9vSQrhJu7flnwK/NYAQ4fLyv1tC0datT
8+lx4NkYnN+ankUU3xn4IsTJDmPmCh/aglHBTdvyyTmebyLkMRj0K2q4NoqYEuQsvDfmHT1PJ6zO
Aei2dZzwi2veiqQm5+qpOMgdphhqkoskHSmRo48f7i3QDZzNyqqoB3NAO/4CpCjhzdqh4B0ZCndl
LVlKsKA7//gII85GCuheS6+5wXeto2WlQTIVBSNd8uIcXdzqu51NQxKTEHy8EFrhOBQuTeXgbUY9
CVH2zLKWs79uQB+zwYcepzgt08gesc/Gq2ePpX0dHTCKm7Fh2qcECSDx40cUkCj/LddMr6oOybLn
tFc3q/ToJlcs+SqncLONVQ4JafIhrUK1Hgu54chbWvWw0Hakir0Ba7sdyP1MZF9ABfd1bQXM0cKP
XoTnjJ2+hg0cFwPPQu/yq73Fpyfl6ljadtpsbgnuOeWhaHlYZRn/wrVjANdRxFwxk792/R96ByKB
3+ptG2zAFG8X0CiTqmPwzxPOiUVwCrzB13aKPVJTP4yQvwi/uf73sdrxL0hEtzM/+ws6IFDyJZCe
ej3wPHQj5dprSKh4U9T1HwHBh4aaA/TsmnvSZAVwExSiw+NEdbOYR9B/C34q/sf+pfVUCzKA2ELo
qI4lpu/wjBsVjYC3fQaQYxbw3lys1UvRHy7eCh5hLCAaV+GzH/TwdpoQTFQEtsMVS3OXM+wyYk3j
upnaCy0tFDbr4jH0tCGwJRLtj2zICRMDgsgOkA4IKFln2k395LwSjE2bk6dnqS89N7wFjbyDc1yq
fd6NfCXqgqR435r5lY1C1OCzQmzsbWNOAXpFO8h3gYzmxTFZOy2hK0Mau7GEOG0SsRGRO+JUgIU1
IL+BVOmY57tynzYwdsTZRdPTifWv6TXGhvjh6xZLxBN720RUdbSpL6NnkOBdIU91z9lOHYLEpH/X
sNZ3XovTrBu3Wl4WXybJD5op5beA1DKfl1eXy0RdY8UsRsGqkaAy8N5+NkxkIvALjmdf5KpFECoN
dxzt6pfMYn/lSyYuPmYwRX6yQgfttrZ8tLCLZFNPXWGVL9HnAFmGm127W+/BbWl5Xtaqr7scmzCB
jqBtMK0jcM69TPReSE7+LyHjmX2iDTzGhxZK5M75arXmNxzOximxd3dwu2yB+noOp+cqnQ3G80v6
hKPeXMjcpXJV6m4kK4bB5enRZBzWrFI0fGcrkDZPBJ6RETZwzGIPTzeVbNeDZJPUpuKXu6wzYRKN
NSof9QiHkg25G/1F8yM7OguwdxWY3vCfbzbTqcWeLzXG/0w6yJ5qFKdoitdkeot1I6uJnzwGjBHP
/53+mGRJxxbctfZsFR2EQ7U/wZwYCEMy7vJvBxghoJKdL2BzI8rSuG3yuYM6LMi3LAdTXXJ/INDE
fp3V+1GgsxejBgw18GYWXir7f8C25YM9UlVAh88jscJheZOcIR+THZtPCpAjVBe90ZC0GtkN3yDn
Lsy2/hXF2FUheog7pZZPFajbPTxsfO7SPD8eYptg48IsxzBaTS/8RaFvuQR+KFZUg4b76gMssB4C
4gIOzlxi3NngSG6ms9wXmFilmE7S1Bi+n6IUE6b5s9d47OEEoO2X9QS4GZzUyYSAe9IsH8hGeN5c
058trPUl7X8WqfbukKukSaRLySxzj+q09OPU3CmdP+GwI0NxC1gLbZeYLg8bqWvOrdqSQ8aJNIq0
70harm6ERe3H85bVmYnzdxpyXwy6wr7rtgBLAyQjQ/4IBNW6ZtAu3+mA/D3igjKgLeS2cadHSOPY
Z4lVqdZipwH7bKvA+UorMsV6PsyhKKwOkFuQGp2Z6QIcC69lhjKWG3ZWoDeuSOtY5+IJFpz0pHXZ
LN7BQP8lgEM9ncIvJDnsoTvkefgzJCnE2NDINy/fqTMmOMHuF7TQ9mx9qLwngGG5yBoj9oq9jlzA
1vmK+KoQpF98cVWBXhXXYo5/PItE6o/YdCN5TvMxj/76zBRGqypl4btjt6hEVWlH8VJF3gx0Aneq
c4sGzGUI6YGyPEB8bGhlOQNUMYKrBo1jpOnVkZxAPZ9t+IaYqeBpO/TaWYEtjwzHON8dP9jMBjrd
7ZMOw04kMXSfuDwAPN5p6Sz12vr5YgO/IZD+APLFuRr5Rz8KQhtXbXr8kLQSItavUFZFI8WmR1E3
9ildw3TCWa9EMHR98eXvhZwRRIio6VC/cuQbh7Zz3flYHMWtOqIUwWSdr13UpUOwxggcRioUoGg4
cXyxVppexxMxGlttdaFWxZq1f/ezRDYUm/2fjmFxFzkpvCK5+YMbkAUmt6pp0v1Jm5Sczn67u3tz
7Vo7yH2AsBXs5qStr/LudS2PYHk9Qhc+belIEDGBVGXsLJ0N38a5TgrPUJpkLB7EzuKNQEiLQ3dN
F7K+EwTVk/QsKdzxyrtQ8g0KxbarpZyqF7Mng6aJcf1OZqitxNgrZFrD5ubO+mo4PGsHA+LpJ8ay
po7/HVyS2a8cI8g9DzGlOw3eH9nweVwzLsp+ChjnDYjZVY2ctAOWU1enBaunEVvJD27RA0xjXYbh
bS3yIpPVT8NeoJGavUGZMC+AvJGtHYyb93T0JxRz3Ev1E4VLuZU+wsswgWVBWIaLJAp1u8cWko60
xWhpH4f1l4igws75LM0a8zMbUTWkjchZG3LfZU+3JqN7gS+fOF9NLSDLXjol6SFDgMn17M5BCXRt
caZTZB97P4wuAPWXe4MeEwdanZcfP+67OA5ifgQS9O5GmUjuRrCAsQFiDtiSwa2KvXIhE2AMD0qb
oqlR92niNFN9Y2Xw2dSApSygK4oNx9AI9xvhEWJd44KoPF7FozMWFnU4xlVpMEMLsABD/J3r2gUV
hrX2ZIB1zCoPIMQ5fYmfjrBZ16R4yjTbU65ql0MBvpbRAukV2BN7LSNOFa6+T5EhcGIuDm3UKR3l
8JD3JV3/IMzrN4HfvXYoHT1A7Qs9PzDO6L3CzO70GPqn7CXLHg0xXdTa8yvED5By2efyJxlzXOvw
aGl2YZc8oIOoHVaxhfPO2rz2857l/1117zt39TyhWzP96N7aJ9lQmq5lBMsmGfV7shx0dohUAOPg
NCNfmGMevWvKRRaib82/0oLysdJNhwGwC7QqRz7Ses790bCQZQhHFCh5Hcsh4Ns4jBLfwNJzl7uU
grv/Vu00pb4hiPZJK8T+OeGmHoCR7zDIZnvH5UjNyUjh9EQClfbvfGWDJ/2m7LROV2SC+bTUMtJ3
OoZLiYD3b28ZR2mE/wAfyDwLRtLgwoMCjxpa/XrswWTsFecdAtlGbVxPHcVZbMkJ7QcJuw5Jantc
K8bor/Z89lusIKhGP1RWfkLmF5/mOqEmUu5QPiepgVK+hBnDU5/A0rlUiwEswQPB4Pg2mzYsTG+H
tBWHlqS2Qym22aDEiTPL0yzdbCmx0xjGXlHn55aeQglvpAWsgBxyBR0CFsEK2R3mcXMJT3f+sRXd
lbqDzPmJXQF0ZalRgmYROanVWbjfpawPts7UA6jyCdppg+4R5/FVlt2jpVrKUhFKAF2LxZVDgLqx
Zppq5e0MbeCCGqqiCHOjmKVwB/hsxXY5a69Kdr+kW5tZFTI16QAiYiOt9Ap9GSph/GSeTlp5N8lE
p1DQD5xhNof4PeK4wK/P76RDZsO7TcXA05d5eUjjjl2877KkStc+VvxZBtKkTjgQHbru383SoylU
SU6yEqZeY23u0UphKivikE9lQBPx/yatuCNj9823pj6mUK52gmGVoMg/rLk+HHuteMUMbP6XqIsa
mivEbEkQhYLJYmZzEXZ57cB4c4oj8+0gSszF7CLkSTm4BtBp7Tl5xh0/ZRgVJ490ZoVSksEtmx7N
U2f9wLxPZCXE1qMpLNIG3PPXTaLwXuTiElYjeGlYM2D3IZFUDx27Lxj1hXadRMYMQYAcmy/UUb4f
4QDRzjVEsfgBYdgmcMHJtxvNDtkbrcUG4og201Ws2Q+WphhiZ+9INHKNlTDEaQXkhcC+ENdopS1B
2CmlFqOlH66xD3kv9TTR5yNyaVI1p9EqTASQ8VtK0COImtAKGPJEeAixvFO9G7IGmN3uRe/81C2K
wA/4zLoxKB30YXoX9Fywv0pIYaJl3c8NrxnyjbjXRR8DUuHdtCDPoDqfQPYjc2NxGlRLcoX0QYeh
D7vgZZCqYXCrREJksgRz4fBKod2pCx92Vy/0rWvPbInNHzk2txqzVVDOWEJYeEl2BJg92ZtAME2T
rAVi/X5XyQ0UxCq3pNvjpxmlywNseOs0NjyTXKEquizMWLjGNcvVDB1KuCJfTTq25qmFg5BdieYi
+o/lQI9gTzG6BIG3ch0RwFPcjnIZmjWo+oPkr8n3QTxhHyp9KjoLY457heMrqT6BXJm7i1JdgIOW
uslJeYtxLiMV1+/VoP+LC6Cr7v/VSTWFLRHcaB3pnpBy2vs8VQB+wFyt13Zxal6eluJpKuE6dsoR
C7YjmD3J3oZXXOYl7mWIshg786hW/qI807AAh9o+wyZg94tjseC8jVZzTS2l5tpAzwbBBcYPs0Fb
D65udLrvP/46huHMf4slV3j94WG0UynxnpF36OApN+XrtK54SH27ED+c9oAv7etFeG99RMELVOfZ
LSn7UzsI2bCWw9oip1wSmxrZ37wmHEY/uGiMtXTos6nbBSkVdnXobcKg0eLJ4O46dQyxF4Z4sO8m
GA4IqPK/73BZuNZOnHoyFs4ZnxQNTMY/yjcUNeMllgP119jskN3AqqIFySpHrZI+TxhU62SvQ8nb
YgYXHKB0YfeB0nNJNwFBP17j3StbIIjepOCrGMSj0kRbIKGQcAP0i/QwHWyxGBbV7flL06q9WcG2
Bk2MxezGvv6rRQ1j89BrVbUhOUHhfAMF09ZgfoPJKdZOJoF3tMfVpmbHfsMijtjzT/UqrEjtIYXO
aRdgzrx43ZPw1wcWy1lFg0gE2VqTUU5djDoSML7QBDTMZVWTja7OAYBkT5cupRGMZxGsC5n2ItFl
ZJSGjxyrZB5MajyGd4bUbAvbj2I+0dbMUenlWWRSDMeSMnAk49AsV/XDKhvl29pKvXB0Oxm+sKeH
o+KH4UEBJlls4DZhbhKiCDkBgjY+Vlb45GfupDsdzQUiizczPQ+ZgR7FxEDZdsXU9XIuGvdnVvIq
b1WfBrQ8zeq42uqt4EnIAMJ6RN0TDcUdXj04fEMQEWDPfIUJZtY39cehbF8m9lspNezk+TwfeGks
6ufV5tcFWeLgT0PEupxn4YLuiAvQW8gYexPc3afRJqMRFZxyX4Da3zj67aclcMH9Esz0nuLUJWWz
U4qBHUH009NXHCzKlK99Fd2zvCOt2cTAX6Md+aEOawZ7T7fbC5zzFDQi+ZtxftmkxzMwugC3S//F
1r3Gly62yIMbycu1ufVbKLR/N1yKJZ5/eiWl0G9VPcpXOdaqkBM1s6c12NrfiD/6JIfbWdh+2YLg
uLTk7rWfLDAXx8rnjycyhr5zhjnAMs3Ewa5yOqoUQP+sWuDuxkPo/CMe45POgtePC7YwcIZCn3MN
aFAEbrneFUUJ5KJIgRcZGqjNsNah0ifAHvFC0z/KtwwVnK+RVIgHn9lYduLTwHCeAvhiAyr9QNGt
Lz7ySfNlkTUmvTRYAZ0H5D9O1y8Jc0yLGlALz62Zec42PazujeyZ1T7PrBuXv2VQsK6XEQ1Woma1
MpkPUXP4aclHaKF/yBfEpR7g9oqlBgmYjbKyZo8XhbUbsRTjRwpK0bS2FuDeyf/B25ly0aLPOLIw
8ziDlp3eBbDTQof81k4ngrckIr8GTUrdXobMQ75J/qV5XNQ9YL8CJzYHRSMQmm3TBPB7UY8B4qoJ
I63fKvtGw49x1P9ZTE6gXx8EZ4xag/s34eE0hCenIrNPRHhConxY35OD+idmCMF6dgQeHE9tetrM
k6b+aDqPqOVV711Q2WNLnShXAiG+aHIVAph7vvT2nVx/6cioYBDxBJ/Vryc0sWIFEIM0hDnxK+Nt
Limd6Jgfnwh8YGnAG8BLbiQ0ikV7mJ/k0XbBGb/9ClNg3uK3jChdouFXH7Tt3+xbLOk4fFd9qlJo
vR+Xr9/v0bsz646AEqd91ELt+HMIXa8120xfUGUAp3831Rnd4gB1LMZ7tXtGmJsv+nOTE8cAaqEG
ijnm8z11iKddKlH/hQJJXZzbABC2FK7iWuSqvVTPyI+J5+3ZqqSgVJcVOHwca8mzHaN4HGop3jYx
DgTA8tSSJA8/Hv0JmylrzDS3Ca+BNsB5+RyR4g0MLKHAdlV6w/eiMKnUA+MRqXRq8j3JdtBPIKvW
qeYCm/YgrRVViRjIMGzAP7L+BhHu6sj7XRPsJ80gH4VXflrolBKJeNQMVAZE+7nX5jYFb6w22zqj
djsj2owbsh5d90YsdHG0sb9qNf45/6DDOxunvSzFmrz2p0Zojt5Z37UD7Imqkvz4rh1ezXiW6w+g
Ge3pDy9Wqmz9F/UoE02L/7jW+Rh04n2r2FZfKk9aaj2oOpiiy/hNO/2pmqQ2wkEQxpF9JBcZI6bx
QfLvRzAfHUKkYzYF/DYs/fxHLq1duiwyJ8TObVqngt/JZaUY6qgnSwxpz9i73D4aBzE2MXEy8h+N
zGYsKPbW2mE75T07y/B9vAQ70YWbmHcqPgW5EiFiga3VvAKmKAGixSEy7FwhAuD52YKcP8vWBTT1
MQnj4z7r8zTpMsD8h+EAB/k/qc6idbAcWn4lePNUugC1qOl43ylRA3XZAEkCnmz4HFVjzoE2TTgr
7Pe8WGY9q4xqtrHYyZYPsBGnmx+q9CbXSTu/NIuPOVshkR9nnN5k4G0t7CN2ox23KXrtA9F4Zg5Q
dk7tHAhvX7HE4tYQ8vS/DJsX9TMitQtepuWWMb5sRYUheUvBGT+6eYuPaDQy6uIP8AFClAtKN0va
eBK8aKWBl9T973IzJM03RUXcfFI8Rpy03LP3PQlnzBaN4cN8ru3apyWTSW1rw/dp0he867rJbqBO
Y9rB30gdZxtak0/ohwxK7MFriTBk4+8XYt1HbUSjvVeqhZHZBAGKnquGeB7/LdPE+5tRV2eiDdf1
29iz1HcGMfzXqq0cpsGlAbaqVXVYAaQA+u7MsoSbN2p/MSETrZP5svcIa54ogVzICbk4UkMSl81J
zhGiPXrosJqk8R2Q4I+k04ET5gctdPORF/+LW4P7NHIHGdGVIl1hxpHvoFAHs0xnrLlTTEaYcj8w
pFJ/U7et9A3Iq1KNdDXkHNlAPYx2bwHGKuSSOJ5CxM74zWQBUL3DQjY7UhoA39Pe1tfl7g92XG1Q
YNCMzOmwf+YxvSmVpOj1Vaw0MMA3WwVlSkRGNfZSmstHf7IfCvvAbZ3FG09TH7xaqKhNx2klEdjZ
IF8hw1x/8QPApj90EY0CE6ZSzO9IbbnK1H1mGNAqsrYhU7ZnfjDqPKgLXBJpwZzZNGqW54V1nPqR
bbVkGgxYySc+AzltSQMX3fJRk8h19foP7SVp3WmPjSP/nuyes1pJY/zYm89du+ZG3uWuLUPKE64v
saYYPCt0n/yAZ8Pg6YXBMa8BTG+N+gsFABmH2PvSYMf7vJPQvtVKRKPY0wtUAPAd/hv1yyC+7p0m
YuFi+TDfo9jbdlHj0nWJFoF+YcKuOJXbC3S+5u/2c+Wqy9OyjkLzqFLQKgUAvgBePrxGM1kGVns+
jcoV/4sDoZ2LWGW5zClFPXyC6JGcFcP5e0MBx8MJMs6YfEVb/Z+9TezqQO7pt8I+oJ0oq6kz0aV1
so2qOubY6ihnaAMotpoRQrU5xjapiJ3TQN22aZc5NtcZHMgP/cAJmT1XLjN9goLq0HvZiBlmJXZJ
/+usyJPIS8R5FKsaRS/vbK6J39vMqGLKsqaKQezLym9kjsmy4KLS/bP/oSPOZLn4Wheu/iEqfAfl
61/nCscxmhF9LL+0sjLU+lQX2v+Kd9okRfeBct/7GgIjAcvA5+X08D6PROIQ+SORmHvAR1qbh5Y9
l2Cnz9+RLZPGlToWbX9rXYCghdFRcD2yebWZqQSrIydV1dx6hOjXEVHXi9yy68wi6gw0sGEMlEoT
iIDSSo2og0/1ViSIWMqXQfZD8d4H+SAumBoWaVRw9olUga2V3wZkO4zTtQeOcCIVKwS74xFExxnC
id8YVRtEntk+CzqMy+dMwV7RLhc4edJTBdmTuI8rgKeAIj/59YLNo1jtkOoAEzM22z6aiYOifvh0
TlbuPpMbWvkUBAQ9Q24i50dqBhqkdqrQeWSc4yZQQUyFJ0wiZ3yCN8wig0dVm/SJWmlt/PrLyimu
QRHovwMGOuCUWvs8Y8dogvy4nxBCbeGrvTLAAGUTiaCvkD4PK57Z3MLBlm6EmYw7+QNtcapVwr30
LLI1d5lKXFao2/K9NLPkCdh98kRK+KRyZyh1CEdnLh/Msf8rZkp/IxvrzCpwLyVfSJyUauJIIY4p
K2qtejj+OpdKowprnhY8enYl0PAgiAvqabd9H3GFgSwWj75ujguhgDQyzXWEa5UlWbKpAtdy7azZ
FCkrkkP+plJ3qd44zqyus9VV0sXaE4yFBvLa8o2riMErshpwSJlYHj5RXux4nw4tYi1EKplrVi2t
iQSUPSkm3JKiIA05zpmy3CY12+YErIWZyHJLoExIvnxKX9BWDSjgncD9Ux4cwbM4nHA9927fD95G
AQ79qvzEA48MH08GPx9WfMTrqazVvKn44Ycup3M9imHDQCdTp6U2FaZKrOqD6buji4yu9cBtursn
NrFwLQ+qxrl2Wz6LaZKCfnSbQZjeuCvW9cntbh77FYQQUioTVrZFP5oWmQrHV0HmyO9PMfALzWUT
zFibCMsHAiaSGE1YupJHIwjwOtlHwb3CKndYHFGJssPDQSL2ipfJKA9JGiZx8jkS0FyHURuH4gp4
ZovW7geLS5Nn1zuDTWGFZgETFTXl86ZeRfAzzlpqQr/pTkCxaa7UQcFTID0gTYRFjBW9zLfSRSap
F7F0DatJA/9g9o8BUmwEc+u3g9d+gmzwp/4pePtMPODGgzJOI+AFxkKREFYkFkahGAlsosN7twBM
GPuiTWqQUmmr4fqkIJBiMbh/p9o4Njs2IEfUlG7Zk7B9a/eLvn9e9FihcMxsNCCzR2oM0ACyTMjq
PAFnCeI5PjX70Rk8l7yPEC22f78kpNi02SrYK66/2ceFnzTB0hdf//3VQxGM+5fA5ZWnRcLg1A8I
UbckmegaBlgOY8JIr1eM0fX6K3NlPthifBrnzt1VaG7OG8YoN+vo2xr7yb6GjEMrxfYAeH/DLHk6
JE9+JxuQ27wJab1syUmCPNY+Hi4/nGS28TqIG17DFInPgCNpEsd6Hju+urAVNBjBb6gVfVUl6l7Z
vewyThLB55iPxqLWPpQQqTfU2/MlVozenrkYOvqw72MNCBZujbYKsmzjS/VCnhKgKVYcn+yn2dCv
6VER7B9dMAhuyZpM56OaJe1hKGD/3rZuLD9+HOT/KO9RpNO4qn7UNR1DvSYlP+2ni7Bf5TRgJhuy
j7MERipCYJxRkLjb3RcQj7QxksR+0GF/yxh4PB1ZPtLP/z+da7JomDv32bAtOtEHWaIcJ19j3etX
Iu6L1O1jbj9qah/YxAuzLMiXQRJAYPRQe3Kchc9SVBwxcK75y49gHRW3xU/1SjbIdalgnxSLBz5U
UX1woaaX7J1WvOPhfdmeSxv9CEL2T3Ioy4iN6AhXC2cFb+fQr/WWInW2twhKUGaSlu2cdWMAkKmZ
9f3uN1fKvIQP5WAPlfSjf1YNFRBxT/wfd/+jZxwdF0Hmz8a8Zq8s49mBjQm8LwCg6dZKX/H8Gehd
gxtmiWqeKnYpKScBB01qXHPyqu08+6Y2/CB6ubDWXFOYsIZUdcrAhz98xIZseBbpdh3lQfSCWX4e
VpG/Jf/JRDFn8Y+rI4cihY5MxGZO/6HIXtpQvUYRqiyW9FuCGgXBPQoQjdvtCEOjBH7Ak6ZE4tYo
jaO4pTzTfG9iqehRt8c+gS/Z9E1eFYpmsckhrx9x8yLqVVQiGO2zzDWOD63rxcb6QIjU8qflGkQe
NdKJvc3QVV4Piu+8KWl67adYNI5iTP5ctTffndE13ZObXe0ySCXCJ7K0chJrmO/Gm/sNA0CH/5YQ
bKEO3n5+XOlzA0BDxwoAk+So8rkXY8FFnNCI1O8bjGAu6vabYGnxmEgKYKOI96ttq/TV1SaNp9io
TnOL1NGKPx7cxPRuaip4J14CguosmxrEUQzg3t1G8ssdi+Jbmh2eg0rp2R323j8kviWaXw9Fs02u
BS61euLaFuFRprqrJU4ijhUf0UFpPFpS0kACWqMxnWl+E4J/OxXf3TlMOnrpDd2d+ZdEEq+9/3yH
hDgOx0bPuY33vkDKbtncN0YsS02A4wPq2sl3b8jQ6PcbOt2jpvlx2O5f8WB7eRa6mbDOUED70FXf
Ul/9TD4HI9raiFnUH9rejkWVdjNwxzS8vsST/7mzBV26tWBbKt4y3teJ+0OwWHSzIXPAaWBYVqJj
iXA5VxW1n0XLWGCV+jRE5c2ma1CfgWEg3oBxJtQwupRtvdZ4PGRFIZg3mDH3qjg5KtnMLaupDiGG
wZBw764PG8cDIFJUTFvtkOWu2/7RhLaeKiN7P2cgjGWv0jG4kYYDwYaWAco2YZXlbZfab1/rT+vn
gghFVFVhG5O9jD3f1IW/ijPOURQ5WYNzfvW7miVT2JYMPlDMgf+yGR4G0Vh6ynVz+++aHo8WZUwb
tVHiiNZo5CV4AZOr5EsCgrQHrIdqtkCe15NKQgffDQn1iSoPw87bx74hbF92OxmoR+IHHVP82WjW
2KIQjGviSm8Lq1qZu5iLPje5Hri5OT7NwoIEqd7bV3pX/jHoKWomc+FgrQ9LndJF08tEqoSo3CGQ
L7dnkQSMf2ZhDx3FJMoIO7hUdLFngxKKC0M/IglJrsv4BQv7CHooG4jrydG60avqobj40VlSOHLX
L4eO1Es+YEqBAkhKk+ZgzNBl60SsJr0heyQBtyo+TJqJbRYBHHXnz37q4FgGr1pLFFf8N0/WOhcF
bhTcBQ+mCipKSLEG5aNVQqf2gPJyW57yogGjep5JhndTqv8EyUhAMkaWMrVkjZOvlO9Sc/T0mXuw
nXEukztCwdatfYMYGLhF+O//DO8DZIR/wIQMzcrnkw554WBW04uLhmYzFDPaJq5SWDlNNu8Rxhga
xTMZzi8MCxuEnZL5kEsY4yNQMJFhsev5q3/twgWL9idizzZSzAJjcsKnLA+5kSkAjRGrACjqFvcA
UkFJcU+oT0U4RqEOTCnEifFOd7xdKO4WFDDPdW52nTT1TMSgzAQPzJmBkR5owh4bMxziSjL4mhOT
sL3IxG2QrVR0+2ExiZAncQjrWRH0eKmOJksa/DlaaFYLYQ8scRXHoevLGaVo4RgeuQuYoHNs6G1w
9zmcRYZukKkWc/Rz+vqK5eVbOhUbSaZVoR+SOurfhPAneYzZTnUtTAxfTfAXxYcZAe4YorSkIgb1
f0A83wcAFNuktjItf8nnbWJ6CNDiuUTgrMFHrOUuz4bNGT//wN3p9/bWK9lSPN2PVf8MPh8f2qn0
7ows+M0RjukMn+rzYISgXvjfvgvcMBw/hTfTQswemHGmCHMxDeV8jGOs4W1RyDViOVqBBB18zW90
5P87zVxE5bdn7nhlJcEA2lBz+TCWWRq3sdOJzrxK6ojKCjzHUihrwEzV1pdj4v/cCQTCFTnYT/Oe
UY9Cb0IA9Wtn3bvmgStPJUWdrsZzBthbi0EKMvKMW2zr4UWCiFR0uNA8T47Hnj1pSS7L+pTAxvdy
8ksk8vPnCLWswoz1Ci6z+F2V8VLM8YQoobRy1G7UylB67W1COqFr9+zHV9GmMh5Goj6QkL+O9xel
ixvsnQ7s7gc5+4lnpMQSXOZHhnR/IHFyjqdfJFYHZq1v/pmjkq4zLfx0UTS8X+kLYFDk1jWswPdN
/PkRwuu9sI0eB5akI5lQXyazH/gaNqJ7zZawhc1SDpaQUYWjbv2aLAT1Cd5jnWfCFThIBgK4x13b
fD77mkg4sKM/ws9umlBQ2B6ghZOpTmn4yUKekjYyfDCmHl5gzkeVbGig/02NC7RKaTuQ9sAQZ3Fh
ralRSLxEDeCK3SPCwRYnWvKE69xyAIRcsBkV3KfOv0BRMaEkaDjxruE3IRogVfDkDhq3QpbgjvBC
fOnXqME0TG05PpurPsTsjyEP5s+N+g4JvvbwR7OPenykZ40aSaYaqp9ErlYY1CzlAMXUaKcN6LuZ
xPQYbExZFM+Np4jK31TuWJKrLyKxgxcBJerfCXn/HnWSnXsONJf7r6E0dx7hsZs+xSsvpv9ZJy+O
JJAxXj+CETdctV8BaPqY1VInnRq8+KL7ipaSh5b7/ghqz/D/a0OwFW/CR4nwqa5+b/O/qN/sraLj
pxEq9hMXnfRsM5snqhneUloIkV5RJlrf3yO6cDF9OjYLxkSKh6qmoHokkXUxnzrkZSooUClpFoBP
UpqV5shF1F12LsVjc4i2myMg1b6PwV6BEEnm5ZBi2DavaNVRFWJXAPWD8tB85dRbJXW7qQ0fewGF
vxolFVY2T6c5otXMP52Ph1tcJRG/Y2BEx9Qe8DKh9FvixAZfjEadjhWJQN4iyeM8HsmQ/5iCG2kE
44tBpQb5EV5KRf1SksWKGwJ1pxoxdwdbWB/UcvnwMA5hM3gMJ49gvBSnQVqQhqyN4tqqNqjaPSdj
Xhh/Y4gAfaN8dhAtrtJpzs4chU7vVMhNwfLjupYO4WSFx2Lq41hvtz6UNs1cyGsXzxK3I5tCC4j/
H46TJI29iNere5ud/qFVsnN6n4p4rxdc07NHX99AvkNGYwetvaQfn5xdlPqBJa12uEMvcdX1/oBQ
bLRUOo4VYIhykdb8+gBdAwsPOhUPgaXnwDAWfi60jTM7/P/hIxQEz9SV3zTod8T+4+6aHchuzJXW
OPZTxUySnEHEuD3fakQu9XF5E1RhGpjJbbc/17+X8mAUBBpHmdFtRT7JbrG1Fjt+Obd/tfl+tVLi
xzi3wtRnkw5W04+tzOplGjRFFNnH7yrFF36cmBn3WYN2BAZ2tNL9veIaMx6i30r6lDkr+aLwvYs3
VPX8IJvotEyS2FQQxI4YsIwMKddzJ89a5ZzaAzQKZa+mSlXrFhF4Z13YSOu9xRO1UPaa9amsghm9
7zJycG+BVtFMSAYxIDqClJOCjIwB+zUm4kTyq2yhXMAZapibdkkqaqrPAvfOnWDhDz5WonU1LZ1S
D1Pz0VLE0YRqpE/QxTOqHFPp1LEkWWGcbqoSkm63f1zUr7+Ej39DRua0aA0RztKgp3ZFbkhzXD+F
jKOgvF3caUyW0dWd2HA8r1H478Avk45Ai1nuHQXVU1sdTVuOyWmhXGAoDhAQ839Ah8nRDvJHfxtG
woxOl33dK3zizGyzQ1Ckh2k+w1IJadOIX5BJEPeuUdp09L7gI841pTUHF5nZHxia4qNKBDtEFuaq
3q2E/P1gmByvlpGbqRTkRBH+828jr06gqokPNUNl2FVaa7B45BPGCxhaoYsekUMqfvd4eCZhM3Kp
UqH7i1PMYOS3neGr4VH/327CWLCQkYaKA6MqgHT1yUyAcvVGnIGUAcaQlZIt7q3I4MMg9mIzZSxj
gpCsH3DVKF9KGUtmI0Nq6lG3ALJgWEbgU6z8Z2tERwyCUcBTn3GC5/jUNSdqrtinmatV/ikzNSH/
iuZwOayZVHtJWY8xC37yUV6996FZCfbwFy9YSKdZsZnSycNCKbRbMKBY6lKHkVdj34/Lh0B4IMXu
sDGq0LmmxKz33u8w8ySkVxXE0O+sd7Mwvn6NBfdNBdR+Uz54PT11UEbioHALwSRfOTsddW2mE7cN
AzF9VZnh5tBDRdkpKEkLGwlnAHxejg5ppkOcSFvXO7d4lilSN6P1bqkRg/GpUqJjHAQBdQFr7+Ex
iSKL0Z12socee97iYn/DjQ9zRJ33jW0laxfxKk8pimtVHnPAPdn6Wufh5M9+Am2exyfiWDdh4m1Q
HqkiX4PN9us+723dT16i8KOocc/thLT4J+RIeUgbKDJ05RG6K4kg0LYXKKgrrg3esgl4GpHDaB1k
H2uQXFx/8J7MjslWmfZExD1ml2ijF0bG9NILo9wsM1PLTamZvWLXPdMfyoZ2hVsXLL9F6yB/uHUd
DvhQxMZ7tjjeEaJHajbmtoUAc4ctNmOO5jar/mOn7oOjRRSsBniURhpN/9UEQGVGhRLUyfLOW55X
xDJatEyUlb5hVxzgit8/+YJiZbljKjbx+F+0zkdYx2lqIpRtwhK2nZYMtaFaDqoRVK6F8/uyBK3h
AvNADCCHXZKqNGFvZHIfE7qQFyFuMyAS4arTE+sYoa3IzcEWmo4hgR9zJTF/vhO4hL2WiS8YwMRt
dX22F7b8jRA2ADwte83oIGAdEaGYVi/GBS2HHwLIQw9q5HPDwjChK3bu0uLkiD7cU0aRkIfidM9Z
AuVMux0XQdq2WDN8g0slGUyYD2cmVZxRQ7UHbAlgON8pDEzoyHdUmYNGnO7ohWj0z7dne7TCUoGj
NSopMdRgxBpudtuu9oBaPoqYwtnyANG2sSASaI3snGinFjR27EQE3U3WSOmOx9+lFC83CifyiizB
TOgAEEl8Aheenr5mM0InVwB4oQftMKyRGWJrxDNDVM+21B06bmCRki4swN4yah/X0hx5vRxB5QWl
b7wbN0jJFmAIwSA1HdwYDyLfK1fSwU4ahRoQQUStroxX/f64HbKhO13UP4uSPtwdRVg1p5/Dikmf
QZCyTZ7g0u/1e9efiK912raz46evvSnCJv6+vdMWAZ0t5Z3AZBG1M0db3H25zTU0n89gIWW6Yb47
XC+iQ35rjb8Kv2U92WIuhNrauFwDJO/LV5Qwre7WlBx8q7MbEMNq9SOTaq8kO/Q2jopnDGHeSZFZ
FIvYIdLYxKRpmURkDqvHfcbzW8aRDnAPWSXIbZATm91BfM34iapFLLiqBG2RWwz1TaNWv5dvHy7d
MOxsub0GB4G7kxvtlqrGJsGHuH+RHMmMaIzVHqYau6IvMPLbFZL+Uxe8hizJdrUVLSeHnJ6hDLMb
aiHLfj5inFUB6RX4kctCLGJ4PuUzJTl1Ne21Zv+zDp2imZczRvsVX4fQz54CuBwweuYEX3TCR8LM
33x0JR6b3pQ6JcPPilSVlfN+dqsriq+ibHTHQbZUdHMqJns8/Zkn8VI4lV6o4wA9WQf7x06qCVJf
C9Tlu4tD3cGb9ACkh94wlt09L2Ud2Gx5Jf3JA8pI3WG4H//CvtHrXwxfSPxEHESvcLx2/+zlbABs
ThZF3w897Yha2D5xqcVxrHshRX1++GnnJZ0WNv9rjykdOL2bQpb9ngrS8XCG/3sP6EO/vS6CiIZ2
FKvayUwNI5QGLkZW5pmaCURGUhG6/C28XPoVozfqLki2FMyPg/n1xJAe+gERW3ZuWiYzBGcdgYpb
d+TseS8jMst3dz7am168Wl7n82sl7Yi/LkOMrXpekWB87wQeawnRvqQvfRs1fYa7IvCBs8lF19o+
YmUi4uPmBTXYwL9nIWLJw5Xqvx/goEMO2Bzpzg8IBfJXtrdxYhaWJaKsH10GEFrSbvEibn9cC1rG
jWQZAycrD7U5YLf2VXhLx/WUWIxL156G0tLQylxAcssfN7VJjDn/4MZEGfzDaKON08V1WMMYpbr6
oV9vC/6CtgoM0XOOX3dUkaE8b0rxnu6h6dCeAE2WpCPrmOWZIxt9XjAOG23ffIWexn5UdQgf8JNp
BnRGPxp0okOcDFP1+C6PLaghxauL52wXpd3VbLhXt9tHq1QngrWEhCz2hGm34TKl+OTj8ghU7+g8
rJZNxzl4JNDKLa34Hm3YpHOKdPq3jJ9JFmSy8VifFzLFyolVRu9lw/39RVJBYUdj5xZLw5bUxYUq
u9dV6P1RBHXps0fVGS2bIT1fJiwjFJ7SBIv1nGohfo1pUhV0ejEKXCN1hQ9X7OSVXJAcJWaZmr4s
MRryHGEUyQ3laIjbV+Yk9Hy6n68GwBZ6MHFRJnKCKlYAZlZDKOhQTHp2/3Cuk8EXDK+ewr/8A0PA
eDDj+vQESBgVwiDtPigBkPNGjByHm4nEtuu806R0rMYmnHmZ56XbJAR5alXx6SnpcfBrHOKUUzT8
Rtwp/926eBWqIyf40UAaPhw/+JVznWEKa7Nnjgz3SZDNRPx029SqZ/9pq6n7DCJJncfxIC8BBIcj
RiCoIagMdsR5rAHe12GNQcchbVmKlnafXUbcTQKmPh1pqwawLWVLNN5zCt/8zQGVdfHxs9brt0OI
D9uCNk2GYbUDsIilrpKbx4PbNBOq5Y0i6weBuegbWYEeDOEuSRInW00yrimEMfk70VSy0eKhXZUp
auO38ofMGqslv3yt2zmuHHVAz1UjmMQl3f7kAIIAZkq+6zpfRXbqpTwdWBBTrWOzW+7CYmAT3jIr
diFtw2vtrn7P73h1GCxNJkGmPRpRfDRc2vKSPwm4gToga5pcuOplWZ5okZLGrksipnVb3K7Qt0R4
r6X0q2Dfcpq/89KHDA0CIG5FI5oBiyDjO4eHJ9FObeayOFziNjpNNWzHQiBajly84NU5gS3A++el
XsStf25+CqEafAdfqZLCrEbXbCvQz61QSqeUzlcxPHQ2IpmBD2LQYdWbaxI29xQP3CelOYDKidm/
JD1FJJRYkVIPGPcWzpokQCJ7LtTL7rQz4QajNaMbZQjLwtwklxrI9HhmBk6CeuzshCDW1I4bM9U7
zT876n8QLyreA+37IL+TZ90AH6/DRwpVVHi3HxZMzZM7261CZ9XCjqq96SaLD6P/b0JonHRmop5t
YfrrRaEyeIHWw4OGCar/HIZw+wZ4EGEYWg/G6/+tVlchTI2gaAKquiVj3ZIMRvwc9kKFeuN+iCNr
bJIq4dSSo0qE3gItFevLsPaqtE5nIBEQVHtpeyYtdUy9oTbRdiB3uAWHb64y1oUfRaUqZ87b0SEq
xSkl8t2kgibwwPOldp3xe7opy6GzVT/4wyDkJJYyR3syDG6uTMXkE/2+NmH+TVBgHYSSyWlKJEDW
+yLDsxOxx/CIXsqRCXF+IEEaYgJxJmWHsDvpaRJhxBEIdxprrPFnPo7YtRe1jLoEceL1KDik6bl7
ClBTobBetD28IxtvTPXnxkEFQFipoKCj9XyBv8p9vKJbgGXz2VjtTJzf2VgLtFmNLcPCug2RFqZy
y+LS+wk96ScsTM+isw+A256KzLPPDy7pLgEDcatSpVSqoOP3PmZ/UT+idh5WcD4Ved+CyzacZaZm
Yytx53UuKIBzGgTPP6r1K2THdsoFmX6JeG3QFOhX2O9GkbyEGubjQyGNvwmVEMIUAewLJeHfD98P
1a78OocAK+rH4mIZalUHucJPYKBrMBAJDCFU/wYNYyZAr33f922UfgftcjkX5JYq5d7aQQEn7b40
uRBIHQ18QBvLQp9uH6IgthAUqZXMIoQ+cxrhezDpX/4+p/n3G831I8xbl5BvAyH6GzV87YgLovrf
34j8yg4fQVDw2ohgj+oQyYcL3J0TVW30AHlhnXnIoqyjkzrVh6BHDT2Bjxb8o5F3/wtHqM0L4HDs
xi6rqL/QI9I6RQdMbMPgGDl6GUZUycE7vUIGYwBii0uKv9fhnDd66UUc0FHbm84mMouOlMuCSn+n
FXVF8ILSplzOLCYc7Ywn+oJlLAjRKUi8iaCCo4C0vEeaHuAZPFcVt4SmFNhcKdPMvstKCMF0PoKS
ZXCNsLXwlJGRHr4CgdnyDPfxUDNXRctEMAeyxU6Bx4ZVX8eCbsr/MMdRIFPFp3ifl2Nh/Er+HTdJ
kU8/dfohBELpcoGRBey718GBMKH91kPDgn5PibYjZd2eKMS1qU0OXG8IS8seAJkfXkNpD0IVlb9z
faOUyysTg5OJWFAaASF29eZ2KzEfuqZ25JgLqsvNJimkhcwihghr/DIAihDfxERzokFLQjt+Kyc3
COWg2yeJ/OkqZMBYyDm2hSCvKGvsZI8O5his//4Dx7RQIbp7nf9h0nMoADwDETEthmO3Hayv2II8
8yGEp7PCWLuR8FbzT3kkb772HbxPics1Yhgi1mjw15+DtiJeccliO1d0f6eBlAHpjFwpq1O+6b96
lCbQzmZeqt2k0xBEUj9k/qpRDNZx7/xY2XobyChtvyzYmtFya8b5d0MGmKoSfolR54OoO//ILgzE
cmEP0UGnNbJ/jv55boAGVOBMMbMJ2cmT9rKQx95/pcOvgFBJpSyCOMtbPXg0K+SjpWcMAxAntsuE
aiYkZsYy4DmUI5QHh1GjGcdw0UKgynV+3jNfURKQ43lRzA/KgY4FxmzyuhEms0rwdwGUlxVNYk6C
q5tLwFF3ncl8egtig4PLkZ1brX35bOo0/B3+uzaKZosF90Vddr4cUzvYt/faIv0X9E3kZ4ohaQwE
cGkvn0ul4HxPZ5gP01tSKIkXAum3F91hTpPmnfapgbuxZaYIwHP60EbV4X1nEJtovuhLVwhSdMgp
IUinDWOrIaSJf5TiAIAOyoSp3GLgecGRjBAZqsCsvKwpXPHox4C4WuTydicz/niHWeURG9zNZr6u
QiYef4WLJHhl9Pxw9gPCRTmEmMC7MN9OF3o//p/CG6E6nILFAxGj4GL38sQ+FJINozCHCAP8GQ0+
fLhCc9ovQIIfgJUtc5kqbaavJP0Kt0mTdoXBUFISsIRHpRNeBRYMMnd4sal4EGFZjJQdVM8sINwh
+ji036X+kt05OHR/jVvbZOwWBEOXg6+zuaCyDoiQ3vJCF21cuDOHP9A1BPJZdqBhOglL6qeKjjz6
nHFOQjOMYk7u0+M6TvQT4jAt5N4ti2LTAzuw+cZzvGH3ldDp6oggq99YhciR39R2qJS8kC4Ha5CN
MmghujEQlRo94ZMIfc3kcmFXU/kjFkoN3UlQ4Ob0l3tfDSU+FwIpimGWVQh/BI+ieQR2A2yd3jiT
8oacmKqKKO/TPNSm/z/4bdrDhcwjVzCcXsw0wOs0krfwr+Q1M1myAmbrZoNLgNvxuF/Pk72vKk+k
EPr63mfPXCFTVqvD/rDuhHYQmckyUY7lkE5QTeWyHezyRChv7cX/09EIlI6VvcSQ64G0ErLIzsh7
RilnMTic36SQ0Ysxc5yY7XtjdVtLQ4SF1VwpeDD00utsJDAlJfuGiOWQWzVhpU8p3CuA7E6Nqn4n
7wdbOqR8/xVLBzDU0NRC+KNg5Yi3kyN5MPbSFl4o0gOIpemQbQU/c83uY09a0U+uMZGySS5kymZx
F30RLbijlJJNYee3N6Ao4XlTa9cScDGZlBbE2CAHr8LWW+k/XBl7PCqtcGscFlDw7MHL8okj20bH
+VBRDWDMegE96z7YBkCpk0a6h8HgOcQoAOqm39blfyb6PZKh9rKcdyXGgzarE0C422U33jSOpsfS
/lAy9Wzy1XO0TJ3w1ZVhOT+V88qEI2XYoiciMalr9FRcavYOjHnjY+17WmxrgDk7vlqmkBY126Hl
nK9VSISdkvey6KuQdPcagiXo4bAzaAOQ9Ro1hhQSxkc7kTgGqxXsogv1XMDYyPDJKIW8uAVzbLgk
Y06BcZnNwYgzXrsBSM0UsVn03CHZC52+Ex/7I+jpVBdYPxqsogrO2V//5sszbfa4C161FovmhrVC
2NC+2DIbbMZ9p6nlFpAVYQzwZ7N8/CjjjxQIImlcaol79XJdNxknFnmB6bRTGdaErGCbVMVuKMP7
r0Bju8NgZvLnChQRV9MQKkFpk6Pzo9lo0klL2h5z+I1gvyCjv7G66FYBw6QgMGehjjzJhDJDtVNK
xt7wUpogZmD/oyQIYFq0frKDeiooBSXz/RwtLbis3EVk/8zw1i5Ufxd9+4beDnmow2VRgQ0nXXiM
W5luqCrUWujJUPiYD73eo/v9smnbpp2iqZZiDetiyWLCp7CUUj1wKOW+04mMqLkezblN9T1GZOo8
kwg2CsZZOLwsEYY6FQ9Px6wfrD2dOfYXMkNTsCQjeGNZRjdwOdLRghXdkb3M4hs/KfJ9+Zji9BME
gb9brrNxzkai8T8fKKSzxrtGy3+GHJC5oJA3V9Mm7TfWpk4HK4NRVC/bpZPHabH1WQ8TOt1uerWo
6a4ff5wcEz8IB9c3CENlByAYDgjfmwQPW+Zw33+T8iEGYFsaUxQ279VK5DAw+75tU6Dt0ZSaoiXy
UxyCOLAK1hwVzcANEAJZwclUNeECz+vtST2KaPid5WJvdDaqaqE+XuQTEYY70SI//FTVWeFAVV90
edsEDH/c7N2OsDNeSnLdOtdnUPknNHMIk8FcTVF+weqHAZoT4Cedqdxo1BgaPJdSQwlno/6g2kmn
FZezkADQt+nkhTAVlAyRB0fn5B0PJbL/qf3Kb3FU7cRoEjdDxJylyTfPdi8Vw7J3OpMHGBWN7jkg
Ry3aNwlihzeWEo+3mzYNFg4TpXtPyF2rDf4F8Z5GFGaC8n/mKuT1nYbYef/LVaJIcX7b8KeqPsq0
1S7LS9NNndrn1bbncgFsodMyuOzoyl6/4SdBP+ie9QIfs3GufT5rDO5C/eWMunco1yrwLfT0+KeM
on+kGfi5CVBTbii4Im/+LcvkhBRGMIf1/uIghzCIjWx4PUGG3LMI1ttgsXe5KfmKHFz2WBf3mNMZ
5JdPnKyTQBvWC//YEpMXNUnHoAXDCNHWOHFTcK+b2GUWsKDYeqm9AbUAE8G6yuuQy740uv202hSn
JJhQQL8xcxCtZs6r97GrHFjZhSFXtoyow1TDWCtpiceXAq1ld7vvtgiSWbDPKjKhl0WTBWsFMSKJ
QDAoub0esiyeYg5g3BbEcdZwX6LHb5omS5n9KZDBSkmLq1ny1TrYF0WGOB6c56SDcxqFXPU5vxcg
m9pNes76bpujEOv+k2nb2Sx0uSyl/hbPsVJOAUvFw8ZQM9PJ9BQFi6klfDnyOMs+E7t6FCJ171Ac
1AN5lp9pkG09jMMfG/NhpjfeyVptEYwHM6a8SKIPi0ckOtrf7nf0d+TXJXBGAet4zM/UjHtnVrCU
2e55tcjnNprsXoz0MtV5I3AG6KjhGVE8Hnu5dcjBDvPKKo2Dxp8fJuPfx7FWizvJ5vsbjTMrWZjz
0ouyOWGRQUp1BVEkpU0xGL4pa4poZd8LkgXsP962c4k+rp+D8JSI914GSpENIh3Y9rO0jpLWk5Pa
oMaHL2S26W/PvcpK1YfNHCN4KONTkziNJNrW7b3+4VHrxNDhjNLe+mSH4gc3gA6//ifaAfZ5EfeR
DK8zotKNlekc4We6LY/w2CDN43iDVq1Dqy1s4n5j7SWWvk/nrI5THOrr49phjpVPPHgByp2XgSzl
i8uzpobMQ2VIqTahKPoiFRBXr79YCPDmCz+NPtuB7T5fXo0aiJ5ynOeO00xEbol45O1W01i5T8aQ
molwFDuEJH1lRJcKTxRJBECRkkXT7F6OmCTFgm9VLx51d2jxSebNf4L07d25G9fj0PNCt0AXPsqW
lgUHnEZk7wDPTaAAwnXtzkF4xoDMcrAxgJkeU3L/0HaLaSDsDJSgpaTdNMh2l0PFsGhuyu4gFxoP
AdtwUMdqGGmGorJIpvupkoZ5S6tlk13xziGCKsGdcka0jXCFmHEHxQnpBeT9cbz1pzAukfSgs08k
8hjxyeUvpsxnVEXT/CMLWOPyMsA9X4ZIBTZKf3LU3JGsxlvlikdQzD68I2D4OcT4Fx12V2gRX0Va
oaU6vGKKOx0xhpXSVmqZB9dXgDTfTVWW6v6jLTNtwPYfjKcvQcvlK/JUyQlmBdApj7bVlX4Eh4mR
zi9LCvZBjHMIRe62kulBrO5CO3DCu7aMj9vr58WfJVUYVeqSny9VG7IYlFQnZhBPKyZ2j8Kp5N4I
/wyVfifyCGznoeVu2Wl7QRdVCgBqFtra3lV8sQQYx6T2ImYrw9HtOeHqOFrbSG32cSfB4aL2jkgn
KxZRta+ciBmFQALLJD0ow+A+v+Kp3XfFb3eWdtAPTW4rgMPESVyAJeIEXRXK6wHuxj68ALQKX9xJ
lbkafngJTiFCNc+TG4hce4jCvbOHS9z/yLDPl2QFd/v5+k9Nqzan5bL1YuxF8qfChb7qbgX6VWpO
ufV3yeqoCwhJT//3PqcarbpoDBmfGrcu5XssqmRCigKAstTi/7Q044h24SfKtTI1th3//Rr0QypZ
EoB9AUBTGPGnfRXqSsr7D8SDAyI5DIpIIhdfic47SxBAZwRkzKllDPrkTPEsYPYA0SSOUs1BwGAv
OQdLT0nJMsZKY8TFG0W8aXTSCs0doX8HdW524yTu8xLvdpETCbFV08irkfACP6WssGPmG2jNIkcC
FNo8Yt6KiUg/6FxBb6PqAvMJg+42fVtVKYi+qDfUvUo2VGV6osdjLmROTPlUvFra2ZnmdscL5lMA
4ALYBcmKuVyO33qEO/NvZ4esOqEtUZ/kquQ309ATCam5GtHVLNC9t26VTv7jtPPkXp3y9tiAgyn0
IG3Fu94tncLtzI4/ahzAdF8+OGX83k1kaRht5TL2DqTqkXJtHAUAruzd04HgFMzbxZ3w+kGefMVx
LKMC/AslqmDms0P788oCZfpQO2rib4kYDNBoJgE2vZ5He0/P/zEsKeILGeXuME/Y+47QJIgUOEok
Dp1OHp6TUj6b278Wy5zjCM5rDVVfmtLQnXFctYZyZ0jzUaTTsjLAa3ZCRPvN03ooq82V/nhXhg6u
tYszBj8ySNkcLrAgEqtFdf3z8fvbhIi70LpMOsq0Vg5UXecv0kA/lDQmlVgzKVIoxTHxfRbbbe1L
I207KI+H6CauBbJPDHJYp3RuDIZSZJU2JOR2R4mE5qFs0WC9QwD76lrfejdY86EtbNLsd7AnpUOk
wv+J1W9Mwm/CqBnPArYr8CTutp+NTvCCVjH9aEheJU67G+AtlYR64P1NVw5MyAjBQmlT9uxokNx6
+piHBFYbpfStEVQT8IhrS3p/0CRx9IwDppth/azaM760c/14ZGmHTwGoOp8Lw1EAhBZPBj/8oEnX
MGkgc8ht7MJ379Ns2zYdyF323eJRd6cnzggzMgtZIQRx3GDdHhCO65sTyg9cO67fv+gfc1BD7SnR
+jHpdxotwGZ4gP4XWm9jbg8Y3taJ0Ct1wRgxHRoTnGuXQSy9otkf4l3WCAK9QS9FDVALg0as0dVB
O8e6dMFlx8kSjHlGY/spxGkmyBTWOL3fF7oK6gbWZ97b4Wb65SjyPuDxbB5oGob6XnwQjkXnWLPk
SisLctKmSIHRJt8cZuzYdXVcQl692ylqX2RCFZMC52fIzu3R+f3z3QnuSGpZq7fQAUo6VxL5JJrJ
OdCIqg+r6y31C77pWjWUYwaFSbIdp9f3D7mvyROubXhgC0GH7+6DQkD5N5jrWMgYgPr/0XAEtnMl
0cIunCbuUp2fmspL3D1r9M3GxAkeeOM/hjveICXAPdJC5hN7t2qyJqcSB0sA6e7z71owr464Ap1p
fULPd2j6yVRd2/UsT8cKBekI/i7pJn/nlI8fLdFtHrUiue+Kkmk83YAiAYtuC7cTc5oTlMr6Q+6l
jIysxM0bV9dwPYCs52wgb8SenfsmNh1tgT5MHu+iT6GTm4U2VZWYvIssTlWLD2rr6R3cWONZCpTc
7j6Mf3scdFUU5y336SIovMVD0RKgSngBfpOejBpRR6oTpbTUjDAbzinCnJdWDtIXzFeImI+IHomQ
Cs4E2i0U0wbLgbeknpqvmRoyffWZYwJyds6Q6OeQDaBySwecwBwig4caZScCyH6qz2OQMXNchtWy
oDV74j8X4Twyv4bBVkx3RvPxBBCCZD0T7WrOgiPI4eRqUmcMKs4EPj7E1uy1wfJQtn91TnouuU9d
0Z1526aswhMAAeq2ZMfKR9aExlfvUaQUZweh25uH5Sk4WOxvpPoNHN7YF3eMhDs27b9leQhaqWQY
N89kwNKsgjQ5qX5VPOzKPC3033HDQNwyus8qEQkmxVt3KtLwORxQn1mZaOd3hgHCTRHZ1LuHXDMg
tvdFeS2AMmLEzVpstpjbxJRo6oL8dX2hnqmnxHxSORFluoLEZTozDi87gUt6niyFK/klvmQ8iUDv
kDHTqfWzQrSOUv/18WaXRSqr4Jx4TycueAODYJb/DhbYSggNtEQ8e0ohLDvs2hhTCtgtBsuh7H+9
4rzCkMAYXhmhT2TXqpRX644kB+XMEh4gULK+K0AlNC/r0l/xuWl0pGk0nDpk5LYck4DMMLxKLrNl
uu3e4K/sppfVzXAQqP+B5syoNtuOpenmuu9h3nXQBzQVHcFT2mFQ49HlTBAbaLcWn09bHOEO7UV4
SncGD5eDiupfNHftv8H/ktqMdoRINcxQ8+rNyr5+cxcBk6OxgujgREjQnACRGCEWEVKejPSnGSOy
NaFhq1jgbDAoNpuiGLnl0dpJqeGrYX7aJeXQLV4EKb+rfygNHGyU/d1RKNtiW3Syq7gbzZDjjLk3
vvjzEx3A//SQd5E0CC8nEei46wbYZr+mkLYWwbLGqbBex3Cs/6igNd3eKHnLp7eeAIudZ+Yd0wXp
yZ135/BeunPmD+3BQqguzdvdH0e2XUIa+IWW6Q2/ELajiV+DOpQ2f17vvviFc0Rv+v3ptZSBOKXb
BtwDt61vacM3rNxTsLqAe1AhEU7QMwM+gs0WbcZCOXx/hD3VB6cWHP8vUkZn+N79c3fLDm11PSoy
hhzPVszZNc8hJyc/kGf2AioDPgK+7eU2I6LUum/7jc1RNaIAi7x5cIruE3xhYm4nwnStquSA11sc
JcxqJFLRhYCJh0BfM5eWJalFuU8XK+qahbDwz0VRw+CrMPNON9buJf/UXpMC3L/6jETml/Q0rXkC
UN7ONu7/GY4ofnBsjBv4n0mdO6IUL7R4XcqkPW0dL+8EwSmhTzLF2pwGGH0yOJ8qiaMzZrzQ2Gld
Kaspmcn5gs0yYlv0kOasammY/rYRE2uphg3uuWh/mBLA/fcDARO7PY5AwL/bUHJVLB1YvODftUaP
6zEKlcAh4TR0pDwDYl1cHRU/Wf0D1HHOTrurDSLuPl8qjcjUUWSplVxcTgShcXAo31mQ2hwvgMX3
H1zFsTfdXtdwYZLFVLNbNWvx/tBoMdQ0rnYpswFNfBJ0dyiTi+Ttr77RWNczMazKvR3wKji54WSn
qocxBGtS7K1+rx6D9cRgVNRGIXhvCXxTAqdOMsXJMt7RaccG/Mo7yot8Newy9hdRx8E53hjMVL0r
IVlOCZ11ycZFtg3Swf/yfhpJR8OS/9hCEf80KbNMLidRy+M+k9W3F/FS7PpBRDC3MHBMkxCtv6Gr
HbbJfuYf0CtauWBD5o8VraWKZqng2Z78YN3bWZrQI1/5skO/xV2cHeQxN1rn92y25UHAMJboXzD6
hZaOQYpxzwxIKHrDs+gRmjMh+YFMjoxNjHGTA83GgpSeHyrvMon4WS5FndMBs6MZSzcotjyyKjEK
zXSoYExJtGCocsfY+RXtQc6nTSknV8iafUC470vgmWfvWCildFVhk3fiVxTritkjdj49PVtL0z6c
RjBOAGraFwxaZRQUCNtUnNSJsZ3RcU7pRp1KeP0nYGu2FfPWsT9o2alEbcIu2TrkRP7DNdWjaRNR
liOF/ClYPaWn1Ng4meMLIjKTeqP80b9F4PRd4QAgir5XkAybwfx3EjsEhuJxGjsfj1r4TLng3Z+Q
qwSb9GetLMK4ZVAOgtwj7Xteg+NHUTTTqqPr+oixAOJSMppYb/mhneJQwEqo9gvqe9CnlX3HHtip
bmGowSwVYc0ko+9RAB6d0tzrtFh9usQ6B1uIPFgaO/nWTif7yIxkQLmPD53LCEQ04XAF4Tp9uBB9
vT8hOPwmm3vv24i4u398UugloZVAjGEbmpBfegfQmd7j2qvChSUd8fA+cPLDkts25oZXwgrxobjQ
nKg4BC08S3fha9KMF/JcbbrqOH4D/HhpIZ+yLHDPy24/E98AliG3cvuGM02SDZQTgmcHtd1H3oPS
Hs4iujYga5c1UwM58+NsGrVZLta5D2HvKYP9t+4E5ONA4vrKvPTvFUq4WPvAlNC6BJNScHD8Xpr9
llxHbz4DdigIieTT/IRX80v5CH9RU26ios8q3FnQmFrPjCpkR33QADiYQhW1G5OA1pxMUgcdulfs
nUms1xk3byqS8L8L9ouPjvtDjGC+z36E6R/e5QWh1fx9UaF18jvacJD6L/aBpJI2yYiBlcWSlPdS
yGyhkfEKyw9KNoOElDOktSmXHlOVuP4v9e/HMjUyzk4THTK4XrJaWRtZNxZEVqtzigYC5QWDaD6t
iJpiWh1qa8JUdvCwbBgagTDZiLbPYlT1jcY0NPhrus3nyAXNFvGiBlbatZtn45eFphFaw8Mljx9l
gsY/tZ80onnjsVDuhsvIa1Ve2vfCcqE9M1YJOBNTDP2cWgCwctsoa7l5Q3kRMgfBK8FMFRoT8m/3
29pb1FtOt4QeTnduQIiVeTkRXC8Us4KdG5MNvOTWeS7hsEI5N6xp1G79wpo7z8sHTz9FBUZMYHlW
A6egPuzDr5SyyB3bwSX/JRk5lb6Lh3SrEdQ4/mSPuAxmA+c1xwlfQEacPIxd792XM5K/gDvy9B4c
RTmDqHPNWdggFYqPIMqm7x+rgIcO21jpVJ69nG1XenCNDxZO1W25NCVtlbB+3rbGUuF/NsSbz5DL
vkHEd/17v10rj5/8JeKujtuK1v5FdjkcGTDP1cgBL9SVlU9e5ixxi7e0q+EUxZSjxBTebFpYFUyn
sqw89dtpnC9Dr5c5dwUQon8ed0q8t//oTVTAp/vqHmzto7Y5g3Hn42OO4HUbCiJAc7EBDDGIftK+
0hOM8xchuZFnDjWqUMpW++5Yhvzxuy/PkGe2tYhCpRNlJEtXxPYkDr1H5k4hMKemvUGvRpTuMt4t
CA7u3KDTrzenpKTSI62iz4bECuDRyYWqZ9pNR5hvjMrZ+Cuwd4aR2kR9nn/SQ1Kh2GpdyZ42DF2U
oGDcAd/NOHaMJEQmV5gSCY3ht0PsYJ/7igJyCnAQtdOcFY6+tRrsMJ871AGgEayygC7w7CnCp7rC
f+45/fpKyAIoMfGvtt9Z8d5Qs24sbjC2SzRtSk8mzGQ6nBaYAynEj8e8tuUIcgJ9BuS/LTCvs7nt
rS1ZBLrgvMyPjnhGdTfUFV4b3+N8VxnYRN6oD8ElL4H8MHi5Es1m+DF6zufnTWM0Zib+G365FXqC
/l7WLi2Am36VZ2CLucRqaHHCjhCnknW5s07RVC0rr6l8FA6ccYuZGSxQE5OdJ8pGZJQ34S5mtMxZ
FP4/s+83Lh5yLPQZxyN3PK/kTpKXWIASr3xwPe9tKs5JlL8GdljLAhunSVI5Ogoxre7KEZcew1Km
YxMS7aiGaQzNeabEuGF+aUnnWXW0ujF194n58R59MmI4R5ecA3HjDhX+Q0vH8Zmk12/tqtpLBdET
OaeAuyIEb/fkq6XNzgzxG/hWlZCIsCTBNiEHO5We2bxpr0u2qSFO0TRCo3Z/pDtAx5dfGVT/KavZ
lwm+qklLoJH6tdkUmq7xL4RnsvhmBuORMas5+QO4rCnOB171DFZ+POALRpPZTykqHrQhImOlvgCn
tqBbBsWnJabPKJASeh1RqmEfzV/KJ9mRwNpooIgHD8Rufc3yuNaf70vwq2QUgc84pYIdVaTAO0c5
RCu6HWwX5VGBaqfvtR9zg9kszBbnGn4kv+OuslLJtjKbSi7gB7PCtSz16jjIe2vPeuOpaBEBZYzZ
yihLocrJnTW0Dn4H9Gvsu+ej1pHgmikiA7sbepdYnzyyBy9MlunBRh1sA5wsMFasCYBIe3iGiSs/
YH9cKBDLxf1KVsX8ey86AcocApPM2vFo2RnzR//fCjB2Jmy+DUMuGKwPj+rQ6QCMHDzEcHrPdHew
boJqVQ15Wk6Xx9F1TXTKnmjMo9z/m45y9N5rf0sk8xJShV9AM2r/vnVlIx9/2QJXxW3wHv0szUDS
wiGS4qoro3tMPOZcgXkW/gikETEt0HGC9MEb7KXEcL/AhJFnxPB9eK0aomKH7jq5FpUeml6RSmeZ
6FLMkM0bVUCgFsBrRYNfX+hTC1UfsJBH3JIxWHQtTjLmt9k2/fT5Wi2xepufO3GGj95WOgBKptxc
p0brlYoxElOCW3pASrfYRtulBt5vYuYznz0V88ivWzdtCABPwPgMuzD9DToVjz51ErMi4rSEcp98
3ebX1/l96sE2hQlwtjfji3u13qji8FedlZZu7stH3zp4Oq3YMIwJCueSpNWqRKesCOM8XYQgg/zI
hBBr2/HVDaYsoFFS5elpQscah6sc/87Sx3vMXKzmj8uDOSQuwVBUlMcw6CingYyHZXui+jpyDpC1
gqHcHfiyDo366mDOF7p90LgNXODpeMMdhHOcUqMNN9Ia56JkBpGzXvnatA6l8vXtk29ycINxB5Ub
H0Z4JrHr3n7fayaFPOaAkq+xTDv78mjt4kAz+PYpUa8zULP9OGefH6LpwSy4txOy9sG0VZWS0kLa
lyGPDq9Jv4wR2KgQ3CzZOWCl7UfOvHfpP3DdGvkjXZtoW4De+uiaAIcxH4XHHyiw4O3wkLOEgTin
kwJFVHvdk1+jRZyo6G29f43AVEi/O2quBz5xKlKotPFMcX5rcCbQrOPrGmQFJQ/mxGiPXVSvam+I
usEgYE0W7YdPw3SkgKjQooEAep2Cx2LtNC3gpVwYWb5gea3ZYKYCgTzaTGQUPl+2AallretHvzpd
Jpb43VosPOLnORyUe/7TKbicYHdZY5YnHx5KqETujCNn25Tv10ttGEoDeoqJzb3gLAw1dS7KqcHU
rr6o1nSyvoVALSoKqPGN8yWR2ESgTVXHPA+J9uc1WPKH8ZtxVCdsGTypucOsly9XTjfTZDr60CQV
d7smtRmYbIiKRgCfEJAqtdL+NQvQaXQSyEALuAyk2fufs3HThXnsq9Awc0JWyk13/yIisejAFRVq
7bN+PQ4hFMQ0Fi1HI7Dy7DI+to4H9SJSl0dPIJPhUsjeSWITumdtb/Cjbl64v183gKlxZ6kijnJ7
eTLbeIUWQPMI9EbZkEAdDSKMx/gCAYx2WDgv+kEKulZ9XLXEqgRHj277VzjFedQ7qOaTkZ4lu2Br
AV7O0e7+GLxanPAnJPAB49AF/8yO0bDjkWfxQdpKYrD6sNW3Srvd7F/HnmLho9U9d8tP55oohAGD
xAxYxbgOHrXmF+UkuSWemyCBDlDBBp2+gq4vMFkFqL8pKRU/CbaqbZoXi42icikcJXGT0nccQBCt
CZ2IPr78RJE0oUbqf4kuql4VbYr/SrSckmc4726PV7CRRMZe7vzI7KraiIl03UufZKqta2vkbvsV
YueJjUOhFs3pXlX17yoiy2dm/aBlF/lE3bIzLUtRaF7OP9VshM/MJdGL1cr8dw/DLkShtXfUAsr0
2JkE0y5at86PCkGlgfSjKu4USTjovE04utnc2l/mO7CFmO+NUTsZkv5ff3iPcsBaatIVlsJ5fta6
v3rQe0Ta1W98QIqGXXDXtX3D/IXlfSRxprt+qpCQxVFR5kI4z4P3AxgOwNnAjkuBWG/VSFgMvQtd
kdTCfSsskcQ9+oRRfI72gA35YrxfG0sDB8b0U84PhgROBV0FVVL2IHiP80S4NYxqbCGN0rcIux2w
bTD0pgMqtQCxUWnBc1lXE5UKC2nfH2NHIq9r2J7vyKLqEDLSWj8a5DQglrtb7pm9/NxxYeoePrvC
/Eyo6aN0JEf0TNhF8EtKaVAFgqqEVRKdNKahm+1q2UvwpLHxqtiNpEaHKua8cfYqUcF7OPm36iLT
BpuG0DfY3LXCFsmGoWxzvYBKwyjiSHxKfOetJjybtXLNnac8kLk4s611thGZt8WhoYJnV2gAq3C0
uleJvOJy360m5iymzl7jZU2NBSaD1uqhNhdaIgHJCJh4XP6q7j+VrsNvKTDwnbmsU8Jgpx03eeIJ
1l8yBjMJYQKUx4cmF2AIhmPgf05504XiOCe5q3l6dvvc0uEeV7ue9BfuYJzlYBFC0Xiqrnmy70GJ
k9X7h+TpLHwLik9jZZBCNL5PSzyggW4F/qra58ZiMxTRehELZBk51BBz6b+KFUFxEK3ZeTm7LruY
L12GxVoKr7aRYXFqqN2yjYZfXMLuRNAkE8qOiINOMei5bMVOV4qvZUKXh7JH5sS6OOHBpEoQLM/I
8kiz/eZFee68t943wTIKCMoB2YD+NtQiQjF2PblbkFder4gNARi8fjv1m/rgVm6nSA5IRH41CCTW
x7M08BzEPpPIaTG2OnNkOUoGFpzkbo0yHN3yY6kqDZ5DhK8CZ1ppOxQH7tmBEloI3ZyI2O0zD4Jz
+bL/3cAMxBFZxKDy5MUwcxsvl7LX9GVi9hJXJ8NQ5sD6QIdpenK5MsA3p2/Qh2puux+d8IZXaIJG
OPPvOM31/16378LqCeK61QvWxQTTEttCn+IN+oMPKCCKs81Po6Ata1qgj4Ks7ytejWYI6y4SVz0h
o8b4wue64UZv3D6oG6Uq07Ys3H7q3jWcD63yxTss1qn1e0wZgwvOVf5/4EQnRaSAcJ0nZg4yzXwz
FbwjD2tamihrqLWCuQyPDnAz0aa6K9MPlYGgNcvkb/kjYz9YgDNZl+v3ld0vY843jg0cptjdDm1U
ZJP5KJh60s8LhjYFphCGRVZiFusKtCPl0ZUklnp+jZFvLlJIzvXp61+C7in3iDVmFxmVrJOrJ6YT
bTMWvdpvLh+tnKryUA8scwtwaqxrCG0+HsYZ/6ycu2MImFQAZ+ZxJyV6kCi12mQv8hjYQpY3IxYt
IW0TIFUdvcMMtX774FzNT2PMTMra+fRqNPc6mlfVtuQSY9gAgRuwiA+XB8o1jszmLaOxr/PlXDnx
odPTNsvLiZPqQmR/uYt+UJPrLgA4iRJUlyT3a9xtaKgSZHz282etuT0m8MuUFmCaqiZQdz4wbEzb
jN/l3WTrgQ/NHeuHoSOIe2i9bNdJ0mpLcgC/YCBwANf1rSP93Q8780yWPr5O0KgYDjk5Mlerf/Y2
wBBFfb4vwfA9qN8TowdnWUspDwW13fs3bUOidmUenNbcjjl4UivxDfoTGCVWmOEp+3Oo/4aTusL9
fSkJ1U+tXiXTlc2DIgR8NWJtIoHJLCR9iu6LYPIfdPSPtpGEXUyxlsAdKdIl9LjtOgtab77AAIXP
RNm2VyLAylXlqSA2Wiy1vP6jeoftrUyPDJiOflIEoAEGtCnPhFefzjq7owBElyxyiUunBUXaPPHw
1CC3E1EQ7/s3GTiavgP7VFXlx0Q4PdZlVpdrzzWeo3PfT+DObe3OOMpk0qT6x6kgHQMwp06LOTY6
24QgBioxbNxn34MxcT8a5N9032Uru8o2/y4yBhaenQEZSGVBch7sxvnGNybIoIxF+S6lrwDne4bP
IrCdRWXoxydZsNyHIr/6CbcSzUh9bS5YwLmqUmv/nKXln72BuTQsnHB0Da4rBVRfwDT/6HiktSDb
71AsuFk5bwXe5eeFp1gXmcY+sQ4YInjsp1W/zeR1R9zxC/xGeTqGWc50/l207KB3bJFZHO4FCfB9
T8CHXCK+Q4BhAgm8oDpWGGySlzEo3gCafikr0/jxa9Ay4aWUbUsevQ2q1vFZNkGx/DAB1LS3//j2
yI+ooQRCtiTC+sfFLMgpgHG6WLhFwCVzh2mFips5EzhVWX4l/lUllWIp1QNGBLZoVD5Tk7z+W6di
R8juw8O8IPD0qMNZUCeO+puD3amI111X7bwbYNihVLmhUq6oj+QryN3Szpp4suJtLObLKv0FD4wZ
yZHWYU9GYvCzU2/Uqeyhwwo6TL62Ts9eaFySutwKdCvsjGzOrMA+K1RwL7cZtCAvyKLNO6HwWUHe
J+B7jg5jKzRjTv/VISvlGzSNGloDYB9A647KVHK74HXpchedKtAaRrYRgFPYUwo7PVAlLBpEFG+R
LEfHgopW10hROZGAFxOsSyK6XbVletidPyL4OKczwOeP+IXJcb14Sdpf7i5ESbwvShjft5l5oDU3
GY+4CFFhCYziGjttUVHP80W7eGJzdPhnHyYS+wJIJz64BZx5qHd2DvXn6IqnPwgXouvQktxlYOyp
pfhr+sCpdCPLDg4Z5fPiohmU8OW2Di7vy2DRN4fsU2yFSrO0KCwp51f1jsSFHqxNrNFx63qNxEGy
yGm6TVvVxM0JRsguzuuQOmVW/NOGqHs9Z4y49p4xVoDMJ/51JOpN5QAQ2oKVqADJPPGdeM44wqdY
wplItiJvZjiXUWyp+x8FNGTjRORAP01bd6NOJVD27wWNrghcBPcuwCeiQAJbsJb1rJYZH5CySse3
LBYeZzH4f4U/aX8bFC+NoL3HEvi+DyFXbbM6Y58Yz5D+vEvqwMOYmscaAiMYtJq8RYcN43G//pDh
vJudiPIQiHq2+jtBpkpA5Zb0RW1u5/RLFi1/L7nupfndy3th1wkeY2AMdTzYqh5uYNu2uesXlZN7
u1iPVxN5cX+wqKVz46vBvppFSshN7pRzQgXSa7tuprGAso1q98cb/eUp1A8XlGa6OtG7/S0Ku+tv
S7ai2lQUn7t7GNzQ5bt35QWudhMHLdM9RjUaHZJnMlWvG+LBLowvP8g2tvMvBy0k0zIA4M4Qs1Zm
CrxegV5NFlDB1zOmcBpsBboGB6VUWBxHzC+Yt0n1okyYST0pRMMuO5NZm6PPoZP4ngVWPFp+00qh
BmsUtKfN4rCit2yOQom8hkHDfRqzuMMJxPW/rmt+xBf3OkM4F2K1ZSw3tAVzoAkwk34lgBrOPCyt
X6G/hTK6P2PrZ2iduBIro9tsKPRlZHjmZjtTnSKnIrPcX6nllOV8tMdm8EmMOyazjd7TvN9XPq7Z
/PMGgK6NJjeQIjM+kBVswuXrwy6sT+Ekpa/oqgiBNtLf4sviLbb211j5yLlEBU9adw7mdcUQ4j3r
FHCOPFRE7uDbmGPXINRu+NEcC1nNtH10IXsBSDrTU4uXAfyJRYOqMT04Zn/Utt3TSKhobDmO5MYD
c4+liY7CqTdeCL7JLA9QBhWGOKgrkjvvkS3pANmyrt+gp75MMcHnjD48FCrkYMHhkauhjw7jQaDX
b8+sjQ8FPud4KYUbv9EX0K+CAuNAGKf8oX/NEciX+adIxyqEmex7bjmMjQpSJ5vUZFUOiSRyGGhb
Fm1ntGNrooc/CkK14F4fCBvJi+4nV4XSpd9YFcDNsi6XQ2EBju6z/iESsz6h07mJhHn96LtT4GcB
hP0waAcldZnZT/ttr0jqU9ywZVm7wrAh8hmBwyvBxjSm2hSPqLNr5/XMCXgQ3/7ZZbpkXCAG+lxe
D5WrSZTLOiErgHFWDW4Sgd1RJrt/XvwzqBGAP348fSpl14WS7U5RlXE7on2CpV+3XEH6RaYThEnd
Vj0PtX/I7w3jGoONNKK29f2RQrRWOIbquK4FNLPiRYp+7H4Ib6vLTGfSL5C1imBoeybTANhETKih
qWle/gUpKalxZl5sq9H3v9yZ1qD4oSlWU1qFEpKU1ddvt4tAIMZZRH0/bHXG0f80Nz5CNUHw085Y
AHjaSJae9J35YbBICY/AzomfV4X2LuMwg+59oc9NSO7qBBxgn0x2KxbqpKU2ZdUAy/tIC4213aS2
ae3XG8nflsTlJtIjQqPpWU6VkPNDHO2w1j5ZvHTM1d0mUMsCwx7sNU7RYYSU20/Sn4CidNgCyJpM
aOc5YVOoFOZfLjE6gWrys/aJ6scto9f7qrcg5d6pmn4mN28x+ONHC8HL00z3fAGPvYRlf3M0mkt8
o+y+ce/t8BPJPGtX5rWp49DGl1pZ7zRg5iWzaRg1mA+f2w8SJDMn6XKFiryGiqSCqHSu8Q4+nin8
UvOGSxUFYTDIQpTKMHpdHRdzszJj22xoUPdEjxHJB9IVezW1+SbEv7veJn85MTlYKU+f7/NzlpOQ
kXjnVpL1+h4+KBty9zVA8nO+rIhDnUvojmKCA2bNdExu3M1v/zbua9kYxYv7aH686NyKu9IYO8c1
P6dpAX4vkPY38YpteBFKwWxcXowYVUjuPh9wUOilu+JZ3DZ2tBze+QoWaUGJmTqmf8WJdgHVHBOJ
yTBt1YEsPQIOyIBJK2Ih1K59e/NrYMTBwasDGy1Ls6fdKgqFvpu0pM+NiW+p1/WUrk4GDtzIRTKO
L5Tv2rqnUYI4n9F64I+i14LfOCOYggP4TS1bpTaMWvP3TEyK74Iy8l/SjLUQ13e9KfdyikxxVXYb
YlCSDuT0oc/OuxbiAJN4+2itBUS311pl6v1fK7Gx7I8Sb2GEuCnRbqNs7/aTEPNnLxs6gvyNNX4D
w2OFhQpp9Z58WqbulZe1NZgzdIUermyB2FzpA3NuWs8I72SYmK92v74vbBWlUEMYfUtXwulvoZ0s
9SN2LhNxXc9zgncgeKzDqiGjP/y+Uh0ew6OI4vtcdOpWiykPiNQcveQ6jZjmlB6bGbpd0E1wO5t3
8UcVxDE3nptIWPWezx3NvHQGkD7RRileVbniQLxlzrkWOaUimW0C7y4rz49VxOWwCJizAUDGZdI5
1xNHlAuWZom999YdqdejOLJUsk9De2ABaS57dceun5P6kk+K/PIrJO8hPdbDfliJYnpcq8CJ4lDk
xSXCdZ72E8fMLVJ/Uo5rR49NRVuizJ/E21H+tVnykyv4cO5SGKeXGMsNsTjkisx/JTIJ/CLuUMZa
efnuIyaDLNlloaykUrwGZih46/l8/jsIy+jec3A1kMs+2WugCcrxmL6cduEL/v4HEXEQqH75bMmo
QfHLUawrEAXVdpOS2kHq+jbEgHslC44zt1xTIe55nr43IBYYtF6ErA5kCrjuYtbj1TEBMckFdLpX
+xw9+Yz8wmdlR2Ulrp/fA1FVUQk6REX/9DAJC3MQUnoPkktUpcw6l07/E/bJN+QBRTH/Ed80Pdv/
GSV2gzrXTphXB+GMnLHr1XqnUw7lvA/O0lIprsoruMupXCidbCSkaOm+loI2B+TNX+pP7wW0Txyg
inqFgVii82h06uXfQZlkrQ61j30GlFMnNAisd5rBlT8JORsMKyE8q6CDAO/pR59mRzqCWYLP8dMf
i+nFjVI6hHcuYJRj1/xJhg+Gnil6rhIoM6k6LW7Eyy7jOFkLEeeAIB6UmMOn6KJY6US5IOR5/lcs
edt0wHmZnGUZmrC7BwISKkFTrX2lucczrTX3c+RXL8RpWfCqGNbReYvdP8EjK0WF/o0xa+UEhzlC
emxsqb5sfV1433S36mvA7+cSUi0MZMAc6JlPE2xjz5DTZuembJPDlA1BBqZmMw6lh+UwKrqotAjp
0ruo26+gf0H4NLCY6sLUEFqn/c62kk5W68EvezDO/lkQukfhkF7FEyfPZ8DjFqEVEuoSsHPazuMn
K8njZPsVOgvLjf5pq8NRD4x+566/nYZ0QMigW8aPOOxe+2GHy6i41wq+BZoNzo7F/phOdUQHmcnA
wvY2QbH1CEco/MF6PqBpvnN6sj4KobFQ+//m5Xwd+VACKOH3b6ZBRCfJdtPepvypah+jKsVJ18nl
EAOqMcwmoaCjX6rMbmJX5yWEqN81uFXq5Ue5yuhH1dKIpfxRVIkMtdIgKsiAnIsrdb4yjDouhgcH
P1zvgru1QbNuy/uAXgeCy9DY+kqsIjVcQKmmjCexwFj37n9SW31fe9i9x7iyvcRTd/FLVMTKfWfY
JCYgXzT3gbTOGaXtsweJM85EbyfNbgHNH8IjCCtnz/p4qVe/V3rUaXlQQBPuwifyi3MGqJ0qX/p/
yqScTRgnMnST3QcuAiQ7WYsbxcV9Ejp10RVI5zrc3IRaSce2Yk5gMxFavxVQaEwaP4h/5keE2DX+
hs2FbXJjbdb+nl2ZAHrLfRG3HfEGiTFwhxN0Rv51wp6Y91NjrT6ta4bH21R075r4FkZLsOZonJNK
+CtScG63bswPLuC9xckuslZ+kqx1nn5spDJxrb0CCCzHpppYoGEAH5fLCeQaMC1lo3H7+ieZiLHY
B2pvKl2FDoon18XPdQZaxmlXnGVxON5DkCsWG4UeIv4Ryt6xI4xEn1NETSylR5RlU3uhLFQkU0L7
IcUFWVbvsB34Kwhy3V4dynRAPTXzBjwBzwvmusK6dBwE/xIqCHOVUj5E+TUIt3LzpY2ieKyvsyuc
663Nkw81Y4Iy0gTuhU2yJzf5NvfDzBiP1rSmMW+ebQZzGOhWIUqcvssgb5IGnTT5FOEU6pKiphVf
pUJ31qC2QtQ78lPYSiuuePR0bYY0AIKTMIWNcjMmZ1c1gyfcYPKq5Y4ao91j+XfzRtwObGA77Y1E
NyUp2h3FNvj76QOhhInWJbALrmG8ZAaKvMApeQAIieUH+LGmKWPZ/4dsRg5Q44bIMNymfyMjbEO8
dONs4XGyUmkqScm62Z2ir1KJ8ATMi5/oal2346/0517LkxAbR3+6Arju5SEXPeFsqbSvCtmS7DYc
vg3zCZETXxDYAxteG2UyQnZQHYFaVwkQkvzi4HIQ0wNm906geRc+NwpzUR7I45M1lrMMwqcFvMSx
cTmCCCsSQ//pHApVEUbVA5EhGHbJqbVCIGUWT44irry5ItU2qpKBeGRQiwZAMF+gRl+XY6wjfqOv
+/ppefUllPi9BLaMIl61g5Z07k9q7b4OP0NLy2H58m6/KV4UIhidvykOq3IFZBB2HvRHAATijM9C
AStxSChoEkOYNMm07zelMTTWVb/ANUq+7PtONC09LGb30piGBWjpJ8d52UvjJqEOxEpnDnwt4pXw
DBd1uOE0tCwsLuK+7Jq4gxmwPeDDbIAt5/YNfBC2eCa1+YQaO0c3K4+5TSDIIjoBm8U0/7z8TKcO
8VfpmwtfzAJ59ieP2Ac8R65GxffHGdGckv7RJSqlA9LjP1in1KpYVl3g0n+O6Yz4HDP7WTs8drK0
M8nC2eMeBKhNAv66/G9hE2bMm9lEp1QVeb/iXyXaSDjT0WWSDKmXdNCNJIJawiVPn7v4wOXZgWdT
muEhWrbnUBDhaD85EOdeUEVDqBYlIN0oW3X0LFP1GU0v+g5Ymlo6j5c4/jwhoWzL8L0SQHOTKSK/
q3OVvPSvBy4invi8RrBQbO3Xk1MY67R8LRV2gdGqsPrmA8gkk9C2D4bextZ0frV9XDkMuC6XC8aH
rGXMMY7AXMaP9qQE11NH2YEYQ40HHikPxCuHesFRafkQj3sw9e4oM+a+2mla9MURi0xzbnumD2pR
YfnueWDBaS1cAIz7oXekITYVpwcLHbTLvxC0nD3rO6rB8o4nybqNLYInbQMJo/6uN1oM7f7+yG2G
TOcAI+dF+dYQA1lyKXKNVOAz/Aq85UQsFTAvCGPKB7E0tg3qbrib5zw7DfLHxYNPhNvGR/0BOzjI
Zm9uur5SjK10wlgcBwNvQZ5YcZuuT2JFpyHwLU2xE+ZGwEJpQmW538XuipblDgJt8G247um67erJ
3kz2rjj0e9W52GMvc+lEPd7WXbB7D+dgY5hc5ulU3VNa3m7xVX1YA7JcT6d85p+eSgIdYp32pxvP
+57RCyi+65c8ZThehnrlnr2/eOurRHw1G4QWd4/DuIrtmDl8PtsJ10cwSO15AWR0tugyvy7CtSFE
kxJccX8yQVDnE3stWGOlntbfxa7Hlfas4Nu/KDVFtFGawS7ytO5UsM4KsNyUXEHy40n00BMxMMf+
QWmgZJsjk7fKH/Dr3fdtjGqi3VvukNgJUJ+V1c3XxcacItKfUmAa/WWT8bLVGyTD1mops51HRNeJ
3iXYC9qGR252uzHOhc2O070vYTMG2rhzSPs3IRgvdfxMq3pbhryu5Dtf5xlUERfdAny758M2GJXo
C8iq0Ifqu2FEnMre5T0aowrWNE3SnUfz8VOClfkAwJ6WW4ICFTC5wG3r2sSUnv5y4E8lMJb4dbbb
lTkU2/5h2JRUuDq+OiVHX4HcxHNmlUSC2QBbDIsbzgIHpl+zMIV5KjY3XvvTcOHkdCuKKwAih84g
UkkOasmkmeQSyOHqqUjv1EdoRWCir0AqkJ9jSmh/g8Am4hQiLmjZDuZG0y8MIx5FO3SDvOcj6irF
udNIlKVXw9ocNHKdrVl5+kLHh8NXOksYtJAw2WcIN4dP83l5rS0vZVVkJF1LUUatSz0W/Ma/pHWm
lhFnXY4LqY/rWqH5cfbboOqrKskszeB9t+6Lm2RsVpE6KDiHgVLP6RgpIGov2QU3P1UO1zOv1w2P
wp3MYBSTMkfxGUX7qWrj+LjsiezfIpHBQHXzxXtA8v0Lfvrf0+YRUGFHkk32bmHOm6EzPlBifopH
zee7QhaKeDfUoDIOcabbIIvqY3qKiQ9nCyZqyJESGYN2CA2GXRsTG69QZGlCDk65n8/ibipa+rkr
vjfvhXVDkpKMbPxk152E1rzs9uH6bYqXBBFsM83hizgBrdJrNjFtDBSPb+nlbNlY3y4AIjivMVtc
pUeMMJT+wE3IWBReoU1GlaAo57BqV9rXY1KcE3MRrq5HiFWvJBHp8KaqUqcbopr55qO4yqMcjaUy
+otPqy4egsM7BLsEouEGC7qhYWFhuiGhzd09agg/NhhTO3sJZ+0Z6o4qbCTl+vDp4elOClQgPpY+
aA78Kt+aVJhPJ6JJRwIaLzxLKSrqd829Zy0KuutFp/IxuhxUlhu8GUQybscbeeswUA5zF+KHeJmu
trkZ8w9DKuGLRbBOwcDAxdEU/dpTQry93gFj3UWLfm/tc57jP5E7soW3eVSZTQueU5VSvtGoKaeC
4Y29McMfQ9c1QNTzozN2+blmwr8PS4B0QTa6RAw1x0h3MfS3WOsqbvzyYwq7274uiCvjedO5JqH1
UNO+5DjpVIMQzJNhg4ju/tDtr0TTeJUX8AZ5U2W+i0H0gvkji3qiumtKhLG22Gf9PamO5br2A9yI
blOXm7v+ntCGeQhZWne7pAv0DPR+AGX0VfLXSspG609FKwYFDVTu3hu3TRbzCe3vwF+THWABzK43
VDBXZK26AI46C00gMFHN3vbvCMw48FbfzbootsitYdlCwHWJ/UxRalCjsSMdNaTfwzgFxOaOhzXI
G5WXJhreSOBXc15VKGf6JDpfGqRDyKPcANmfv1MP/NDd9X8UPitJ57pdL+zNGLUJPFbuN4HKXwuB
krZCOsair7nhNofBDLChhFcVo3i8iSy56JyQdopXOPWBaYtSuLjrFqCEH7k9OC6Wgz2JdqFKIVLl
/gJulJWH5xd/h5DIG3gUzzS8leGqf56YfkzHyyB63mHbPQEU59S+gLpfsnw24Is+eF5C0vwwav2f
+GRySRdF2lFN4ep+RT+Ypbev3nVAQUGD7BA+YaUj9p/zxAM/XnOv6NpF/juuc3AghZ3o12CaWFcr
l++FwbVE2JGAf2Dx/xIv84/lB3xtj3mrvKp0ucMwGTTVvJlUJym/AMip4vQbEIJbfVgh/VOqielP
INiaBjjP0wzL9Y+ZwpGLJm5ZyKihSBFKPW3vAlC2uIvSB47YC+ZxiP2xmbmADnFqQfaQ6q9IGfyQ
YgeWv06ljBhjYVjNxLufKHo1yiFdBrBN9OhuX06SATb6vn/1nO9BavRjG5+ri94zBI6ZqLqHJzZ+
J5Z2A6eGI60XWxdQSihupA1MvHCkhNFykDIsh9PTOBBWcLRBeSMN4dIncAt02OjHAaa0vvIfI7cV
LbjPU0WrWirKvy1tt96vtWkvFUUfEJPIcw+LJ8N2t7CCQxjG3Fs2Mcy+zX7HATlZWh6VR1yMq8uE
oW/vKtL/eD2t6ncrSuvX5e7A5nlEUsER4ZTcUcDh7r1MlHMC+UtbC/SBK+Bg2bKEQEAnIShi3Ui/
qzYE4vcxNKh/HA2aTnoQyOY3qgDkdAx1F0Z+sJXW9++kvCKJb6lkqXKigLAWxxCZvc5gSe7eEcf0
8wonMo1vhDDeVjP9ae8v2qC0VqkvAnOiEPQzO2mx80SXdtthEHMfIzMq1z3v6HfNAlJq6FffdWRw
m0R0tloqsN9I2MJqxuqHk+hFDXemRwgBWfwYu11wpou/n7eD5MKz1dDLaQckXndraxOKyfh02Oty
wJ85QcOobjdrqTiIsSOItA6GupZ+jQgv3fVbwRDkX/m9FUUOIo1js1Kd3bPtKSsUFpyv4jbzbupx
oobr86Bq778nGtQ8aQ+xA+/g9w62EhxsjoVE8GP2qNkP5DgulSJqUFkgenNG6Wbvhiu2waFDyPDZ
QMwMQmKDjSzZPVv3XVlUkvvjwCE80QVZfn78cOLXmriItY2xxu8nOnI/MvaK7OhGPGFo3Z9a288u
iPyTvwI4xWa4nfUXczcAzK7dIb0cKXykOakdcgeIGODKTCJKgWH/Po6mog1+LrIqBhJQ9U5An6Hx
wVW2wo0IZEqDvVSYWEDr900TrEHnOGY+Ve+KnNStC5eLCq0EHAsqcTVUOgzsb8anne/d0Zt0p5cy
VZ9r3UhYbfVSMMyHqEz9y6zxTkoEzk//ZscLH24rymrYLz5pZZ/gf8HSh0lCivhYxywZ61e1yk5M
OxDLP4PXUcXLUFDCP7Uaq6A7wwdQ/sqqLNBnZbsFJSa1KtOxKh+RP6VNlzRQPLqZyU55INvGnlJw
wZ24wBz9lScse4dQMrjI5b7UFm8x2uw/4XAlUg2nVARqIWUOJSb63hvY1X8k2XDr0423lQxu/F5G
+uvP5MBMoJ0PBIe4gyozHv9CNDFeh/pHgwdQsmmm+POtGa4a8hLuxzObUisffAWp+tVjUiqsC6OB
y9+NNjLTaC4yN81Zk+ncQqXemoiUyOrRpgn7jIcrHeRV94h1AQ6AZRu9AHLkx4jDf2n62Sd7Kryq
81/k+E81G9TuGX9SQkUzFebQRswdv7Lt52tpyHZqIaaRHCjEmnXll1Vr3tR5uQ/3QxX8s9/lcJsQ
wyh1fk5fQWGl7CsvnsvvXkKeWimKi3NPIbd4NbTGnm9RKQig2CxXvQYT34KBT+F+vjeOzLnbFcTr
rgyoitASNdjHIt1jUaDJJEZYfM95pAAkZAIAPCpDRS2kvJHC86KO6KoU6ZweBxO5kt9K6VNlWTTT
ZLDwcqAEkkCxGr3kUwH8NqUPuKX8U/Wncy1eoMNmEMFoxKVPZFmvIlW5Wy8sE7uBtk+S/MOaFw39
aLnNVXZKTSXeyTg+DRKedVjwiyHEj0mThEdQFnHr16XwGC1idKxpPH5/aZLsFGWiqd5TwMA2fNR3
1P1NB1I3hV/sS9cpcyxAEAOChN7yGscjjUSeU+IMuCvmNij5oudpewor4dygUMOePcPObKe9b+KW
8csr91fmgSSbAerWw+wA1LHWjSjw2/QxLYJqQx9jDSzxfLMuiGFrSpHq/Nzug6uxJfYIv6FL6Q0X
mhrzL/ZURuw0KKxErKsEq7Xeik/Ffl07PbeDcnGIXtCljvjru5x2pfNR/0R13Psc+bcnyCC+XDio
xjs6Ui5JzIkaZrB2glSvp/T7XUBAkkJBXUf6vmI34KlEsh1Ugc3iQKgUs4Pb6fkHVRbMB9BVlHZB
jjk25+QSG6i2u+iNTR7rcQgRIFfDEGoIb0kUaV/S/NwHb+a+OiVHTGeUuou6ayucTwODztFeH8fa
1rZcVmGvdIvDr91Q8wTTy/x9GP1wiC5YDXB6c2zQgk+nPFzG2rc/yhi8Lf+NAmU5ViRokcMLPRkQ
fZkHmz0IagXGwSj2CWFRgRPA+g4UKNh2aiNgK4uriYqo1Bg0llcNkSk04LgDfcLIhOvU72MQuF7S
HWc/Sc5FSP1TL12w/DVPQopJXURT+v+G9xVtilaXWL8H8HOhd5c0j8b5bmT86Qw8u/YbXDX51H1g
jXq4a4BqsgJVe8AdLGoVgzmmuJhPvuRbqIL1pawIXZhlLNXz6r/OcbUu9oQJRMIGx2RRQgyOeYfu
B/1eXpFZ8P/q4OH4OEBKGZlnigw7PzBrnAGbH7w/ZtTuu6ftsdrXWY54RtDUrduUMq7aH1d7aeNH
dhb+r13PnKaTeKF6wTBGWCI/1VsiY9EljwSZ9Mtecxi/14P7WUV5omqv6YIi7eSpafZItoeZjbut
xoG2F3tyPwQrl+EBD18xjWptGcKLHMR8eyOHpenXzniaJqmN1qOnhm79FnIB6A0kPlAAWJpavMFR
aKCv54zCCb6GsqZDaBygb9YJ3WxoRTEB/SfZXIJ39v5IXgHd7PvrryBzBr8EZ9ccKDT3jBsy2gKj
YIs0MXgIbqDM6VtU9JE8wAC9pI46HfZG4E/0r4ySVhlip3hEejehMP9BdwVG0sOnwh+bSG1qXixQ
hZOQd88WcpxYgGKM8lpB1Z6MDclU+pTHnhtE/NCwAYFumuIUslIzB9JfK2Qgu9TzRQdtHEqHcJZf
sN88cmL2IRLV+rfpYQ30cZeItuvkwXoBguZFWBIcu5t29C/C4RrsPngZMAE3fp2gmjvH7kFHzkXn
jKhhikcnURfvoY3/phcSEGQSdmenOG7ZcH8GU9jfQra9q8Vq4gbJFNrjm5wehpb6T6wtdeoKTSaA
00mokM713bG1TQ5t9SnOuFPqUuFXi61zYBWTIge9zh/aywXc9wALZPfX567691aLTyZIvsMlGTIm
PTt5ZbNTG4sCulwe/p7batCbmobvIRJyLq/QHj4hhu946l0w91FqMKOwjtNcOvoYZYI1yWCcE3I9
CcNnIFLi1C73hnloSThhD8nG/Q0yYEvbv+XgfTq3Yxw0nGWR3WmnGxkroqAENRcx/hdRO9ZJD888
XJ3qAQTHNQSOKA194qyk2+l/q4uoX8fqrdcM+gvMExGHV4p12LAXlDo/qbC3/qBkmCJ15VTVNuvY
sK26gklPYdRkupLZARTVnqUMvPkA9J4zha0Ri5EYeYsIO4Yf5hMJ6/UQtsiiOjgEIlV1nYe8kqdk
x9NTX2qIEifcZfE4vqvWSS6zyOIx9zqYBay/3/bq3DIVnX4zDrBEJ421tkuN1KJdIChl3NmV7uMQ
cVJztofltX75SAx0sABlDmvpZgqZSgNKhaeThy+3ZYInCaRTGuAEu9181EImDFtT8Ku3342H5qPx
9Oaw2OrpIhtKJ2KHjtGq8wMaL/vVMYHgyVAv2xvrX8rvkBLUeg02IobTGTsmzaCZYnZyRWt0n1kL
0GQzVWl64cAWlXfBwfkQ4tjTPwZvEOTjEa3OfcFQF/NTLFK2rnDfeTFqE+Havpj2DQoB7wXEbDwn
ci8JeBiSTvVfsDvild7/4grKXDRa5edbl6zqg4mswSISh7M3H4ZWSsqs5PpvjOlQO4k/m0bMSWfS
t1uy0c9PuAIKoXNZEl1TeoJdY3DjbKSTU4iLlCyIeUPiRB92DEC+bHmu1HKW0X6Ahs/8Tt+nfCFv
CbiIlMNV9Wy9iOm4fDDv7awyLdZTNHAheXKn+PU/a9Y5jSh/xvU8lU5qHVUoa/SLdWMZJn+qT8q1
BYmSDyZuaQSvSDklF+m00ibTDNPzUhGXwi+5QWAJgFg+u5oF3FquPpasPWgC4CYz1S5HZiQEQ+zN
2j3mHSIhygIaLXJjWJ4KfYZLOu1vKOrYWya18TAzGfrtG4knhkz7rQ8MsYaaizCsAH1kAJsLCpwk
5ry+pMuWqWALST6BYvTHk7Lscs0PGQUHLTTqvDIesfHJ3lFRkdJLPi/ieXuU3tdrVgm5yTIbGtFw
xoB4pyikA7UEXiRD6/JK4EHyK8naRSgeK7RhmQLP+yEmjcj6yno5zE4SptwWsb162SBqCTFRiCJ1
saBJg+sQm9ZDagVe0uEuKKZ7bX9hcu+o8hX4v1wwLpOuMCu7RxOzZTFYqXxisc2zb2FPAZCpX2T6
97zAyL/2MPyFXjkgW6+LAydM+Hesm4aCYqXjoBJZQ+17L3xNNXL4eAtofKLelUmdgk7o/leElQa+
Muuw3v6AABivf/KUbB1Oh4xrAfWpBh8P/6PQBiwnWdBcBe8pxBx40hmjaWl+Ae42aJy4VDYFDC06
krHWU12ZXyVqzeo1Q1oHF2NA9HTtts4Sz62UA/hoGNjzCJt8OK6ZP6c/slxTRL40N6W9fZtpU/9z
c1p+T7cP5b7AcbvlfNa9xX+8Sg08BCvALdi3h+QOXlUG4zuPQYJHE4uhmsjh2FvPMGYzQ5beuqtf
ZQFQbrppZv8g5hcmPAWgr3E0f0aZyvS1zc8fUba+sBoAzK0zj0RvxHhTOtYzA0EgX6cktqr/yPvd
iCtzkKXz27c/XW2VBrmsPr4liEZPKUMu1UuvXlmJwmBMAJRXr04Mhraqqp26GsJpTKKWEGOOl0RC
mBmfNc1YEyJJgHHnYD2nem/nTyqhQs8+F3cMt/NGnjgXJKxyww+Zib7j1XvziV912v+bhAvKa1mG
vcj3UzJcdxCt5O5ekgVrpQ0jFK8ZtqzwfA2jj+9R/P17kD2ZB6bNKLtu0JWwOmHmxDK9IakXqRu2
FHs5O3H2U4pDJyq8DWxJeKwi4RSMYj51L/bwv4UBDX06ufYZH6p5JlrIZs5AYLObSib30Ij/bFes
DsfQDDTuIprojn0lQRq2l1Wb8wqZkEkKBQpISWMVm6/pUPPjSOu110CcDba2TWcynRcAevst0fRG
Pj0eHVlR4ixksF5miB7KP8iZtQW0+YR8LRZPoOPbwCm9rUBVHrUUaqz/USWentPTuiJ1hQH9Uw2z
hGULOx+YHfwGQrKy3zqdI+v6ZfAZYmae2vxIBpsvNoHGET4rOY/X5NZukzkHXGPNtDAHgwIVbMl/
cuYSrBYFqKDGiYyq4V08BL9ySBrIe6+2OmYGZ93Egou/P8u5zoGEq+hPAmlOaQE450s/KCZaL3XZ
op6m4BgMFPlQne/F6wiI6ASSwRHbIXSnTmIfWXBn/7sUcvf0VRYuZycNL5sc8KbkhUiI8oXA6YTN
B6z6AKnNeX80AxniVO0ORDsRsXm2q1P9b/76YYew4FS4WDq0SrV+I96ytPm6/RXpB5OeM6Fp5f9B
9Nhp34CNY2mkaNc7dhtJx/m8crzwn459BLs0L+Mq/peXggdXGhZOHOmsPxEv7Izlgqg4p7bPlCks
2awDmJUjEaLxJppvoNN9RrMsbqdmv4Q/tfDLtiNA8DKgc8QovA+OeNUmNaHGauWG7Vl+8mvTxgC1
QHXQvg10/Ag2nYSv+6EY8HVB6L9kGXKpxIcX8BQW5dFvIUTni1TWJ5cEAYYlhCPMf2CYGsJ4Z38x
zE2b2HD5ET8ErCdStje2Xr5S4c18dwZtCupjiFgmEwRcrYiNEICc0ZO+v5uSp+ES8MDZWUZi5Vop
/XxgqBEX6dPx/YTlrG03hHVsa2UmINYcIMvhJW4BN6IK62zS3RMqk1NiNQmh87RIhWzdfiEPTMVc
S3aQ/mUO7iLnZLc2kp/SsNqga38S5ASR4JnCa2m4shkQkQ8h9Sc8bqYbE8m37pMajBcTNYGqH+zx
e4Bo0fqBEHjc5PvFlSGJqw2mxG+xzfaK9CUSimaiqOML5w0bI7r20negfwVI6pVFGDZrBwH4kZpt
6qbYXESoMNNk2c6tFs5RtAB/q4ZD1g+BVWdre/iRJdhs0a+wsWvPOG2v09zQT8QStdo5IlJOPpyF
gBVaoal6Oqhof8nY7/J09d8PVTxqamALjs4KMWO9Fb+7zINXTDOgjqgkgwdq0A+0/1uvBs6j7IGe
H5WgTJXn2UWCMR94AgtuL4vBtoHHLQ6SO0O0isTdAk+kkD+2G7jsep64UVI3QSyvMKFdh2oKtJKC
6GM5g/k5S7zXF4aXB2eKxY7yGDAXtfG0KcOaK5VO9NlLtc6zwLd75/t+mjGS7fGDSL1N/VvomXmw
pwTbSxcL1ubIBvZOxxt7YP+QzxwX6wldFywLDz9bQ5NcljAL8YiGMbgQGxqun7z48QTmdvUdxOrN
ry7vDW2q5vb5Qf24W9v/heRFFmcxE2pfZddIxlYBYEjLXTH03IDurm5cqtRy/5NuBCUpjU15n/yo
aJphVxXIJwXgYWuBetHV5itp1Ql35M8wp63ogphqZmrfmDUFBRlThVHJawDGa8DFDOxpawhUn/Rz
8M0dNYlcDtkc/H78Z/RuWJQBEtlnmhvwDYR0cFv27JyFLw2WxWq9WpiPmZFcWI37vAjZcYhRuqvd
X8TKm74VgZefdb1cJxc4IXMcfsr//U+mkhwxsRSxFlr5a1cPHis9LTXsgdrOE3R2eLX9I0BGdRNw
BUy5YavgpVCA86nBCfckPCyLocAMRCoPF9Dwknxqu1lJrOG4iTipS0ToxfAzNeX/RniquCqMxBmC
9Xtjxfdm02b/nqY/uwucwpvoE6xi7MpwYlZGRhUjlcObehG12vEGzgu1Bypb9JYnfwG5wQGrMkOn
fRYAXVkqMMdL3FV/Ptc8nJU8UaeNRFVvlRCtaCXHxY4v3o2iQlAnb0hnoqznho8QsdLsl3ej0Ijc
Pwn9xDOm+lwT3epQ7FMvAhYQyOxceMzlUN5MDtO3kQa9UgFM4Vb3H5t6kP6CfF7OmamBC/9uZSbk
NPE82Hbsne5C+NvEEI4TKyeYK4HCe3XnoB2uhPXe1oHf6tsFzqzSRhfQfv2d5L0jdsPlWw1fB5T6
eYy/K1gFmvhm1J5kbw+gsLGM+xo69uqeUaY4mD9b6tfpSHA7yixn2Qb9ZqObtD69c8FXYOaZIZ9Q
O3wuJKYRhlltCZuce7G3I6gspUR02gAsuAJo+VdbVTeaMnIk3p5fc+mk0YYurcgkh7PyHRMMtDqo
biTYCxhETNi1v1h7egW2tGFszeKucevMvisE3JHaRbQW1G/6fNFoRlR/LrwgClE7ZCxsVqozU+G1
bJJDQpvHn8bxwfdp+2DH+gSbLnw5B4YOrdxZ02ZhsCJ7AyN0/0Shp978ZCBu9tpL62wYGgd8q/jD
kKikyTnJuNQ0SQZbNleABsfmGLflZFV1j7pWMfCEpWmhIqJif0B91Z0XvEFK07QpMU6RGSmx4WMB
lzgnjOFh2wGZ3JBeKdO8e+fh6lpkQHLY9ai3mu7nlF75mKkc/ArKrDZvTeXTK7b7gsPKC1DB6QrF
RmVh4QA844KNsVTVZRDXsy4vfTjVVf67Dc3rt3BVVC92p4u4D5GTmI/3Y2z/Wu5sM+uyX3kfz9r/
2ojPa/LYhexLfNVkH9V0zHzSCRzs1YZfc7mOhGv4vsaK39Dvn4YkbjIsP0MjqvpW0nfGjjr/u/BG
rMyyefHBmohDBaVIbhv7ontxZx0N4HJcgpTvZtuD+rOIaYCO0L9bILZ2AmXIos7gyPupawUeyoKp
lIEUkCA75g8jYNNzwgr7L1OaDwmiFg7ILHjZpOQ/kvDHMQoDyiA0XcSghrn3sC8FIamzoJCc4Mg3
Y110WEDHwKfvSXHaS7kjkNQp5tyu80mjftLFQEPgh33P0ixAj1e7Bh5ARh+9nNZBX/ptEXmnNByA
/Iq1EXwT70OEbRCANQIOt3O1ibbJdGEzHBVGI4YXm0bVk8jBaes7PJcY4HHhfACFW3JTlsKkgXXU
uzDDY+7jfWDxtm9j9p0MJg5fII4A1y7ma1p3JEdho5mRr+fFFM8GVOYnXlC8tWl5fKvYiCCSg893
18oTg2K/ebuEFqh22o3iV8oLTY7TVZ71o+QdOQeHIIG0IpZhcnHbggmyx0aETevFHHEdrBDOvPMY
DqqRfXOvG04xxyWhkY4KfPY2vdcP57YTogpvr8CoqOnwTLZVJJ9xg1rQ5xT0B1+eyz/IaXFWxhnr
FKEyk+Nss843oLXmMdmjWvI+2z/bUV7vIDHKaB8Be4IB7pIqG57pNUSbu+BCG0LHrnijlsVIJKze
OaiMs1Pxe9w4xB0PRxmahmqzzzEDD3VpTeAcgF2f/uZP5Nfwxng5m1MPAaKD7cCdKQGq5cQBeC3o
yDHi90nRPz+QlHDqGwz2apG7HSaVclsISeD0AG6vftQGmcyfqnHPTwY2DXlBH8DH1BFWSsTkWqkZ
7552KRcQOcRsByYgd/rcAFgKFJTMCNaCHg2L0jY0ReFZzcXxQSuMM+FUlHEb1Bwqtqj8jE6U0mbu
FjjZ9WE7v6DQmuooa9Oc1mSumVwAFPIG64hf+8G1JO7Z2hqR6h2BOkxd1HA6Vj+sBuVN+wOKJWWl
lJ/E6IK/LF94cByS8poxFa8zyPSxSCQrk2FtbLYNLHUKF67uqFic29klL6Hat7x0OGesTg2Dawgm
Dsi4CYyBw9vYPDKjPDyrHeyMtPddiOhr7yR5/humO8/wzcgpAC/t+z46u1+ghuxKb9QH6nQiqxdK
l7hJXpXWpJ5WreLnnYHhH4VQ35Or9hw+euj6kScLoJaMD4rjxtJleI3zu6skjwkqYaB31JGhwr9e
7l/g/doDC8cjC+J1xOR5f/wr6VC6TaYw7fWNfgD6Ut3Ae2So7QMKr960h7FoWIRJjs0z2wTvrRdc
gVKs+h0S0mTxz5TunUhUSWw/Mzor4hHu8vLGUmeF9Py6rYijdJnHDBjEfrmrm0wzdFqKgN/SvTjx
sOxwMdxyqaUSlOV1+bKCdc/XguPsnadc/mhzNJ1FamsMB3Q7+qzAEC+QL1utQSoufCas0xPWOtTC
H+e3SZYgUwqGDUcETePJQ5BaeWsNJfNKhYSoGuEhMV1P7TDhH6jt6Gt8swQ8xbGzG5FqTIAhGST9
AcbWXzkqAEPV7RtoO93VlJ07ZmmYKELhxP22Bjkh4bmg0/Db27v12hfjrRb5caxOEGGKQUfyoT7q
65w78iZK4AxMj+qc24ZwCTjp7+hGVM6IeHd3+RAUilrJkNknYxgj4hpixMcP1nyYNLwyiSk6+lnH
AUHPOvjNzzYJp7TyWOOQLCgn/hb6UeCf61uclz2Pl+cZj+HtRKYIogIs3Y9vrRsThHO/hFPMpRkB
Z1DjJVyKUCfQaVoqnrjuYgrS9iuORC2O0+LbxpvscJw70ClJCzm0RoqLQ4ag+uzYd3ztAAT4zPdm
ABEbL+qClR4kOVN0udV9dyjlZvtGkecmn2wiGO90IJFM9jU0+rcseKYaNYDb0lPVqUdXJpxzjFr9
FgNgqCvnuljbXsBul65HiGYeWmjff3WRisBA4bFnUAv95/u+9LYTsWTEfad/zlfLVeB37cbdB5Qc
4zADov1Lg6H3x2PbjeqFswMBodqbwB5i9DvrD/lFFWeG9CxG3YwaL9IRC4wZbnXMPQ2VknbpEv6F
BBaLkMJ4TB5BG3KH7NC8sKEUuCwM9RMYn1RewT1w22y5SvcX+AZc7qGiJwbfxJz4tJyw7/AS3Brx
l6lYptfmFF/MeMgvt1daXZiA9cEch25Zd66mReEN47+6M8Qbv0ioy4QxHFawSlNb1/RVVtQwWfeL
cFNVoQy2zwntAT8sCMNhe3YVX0VpznaOgMCbyJNTk5C0Nvi69TTySKfSKeJ2SNJ3V3irSrIb76hK
dERUk43kBjo07HW2xa+25FZXSyWJuS0zNDH3o9DCZ47vWxzrMZHHci39MF+yHfxaQwKzqfUDAsLn
5CkGrojNGZENWqpIsv7Z9WMa4+KEgG2t1dcnAX+pceyekvuCc8hnLdQxG3hEa4Co3EluzGhWOqxc
oBgSudzBvuOM73q6apHG2dMpKJao+OdPhS1sG3s1fhrLR/0lVmKRi46zH4plQ7l74aoMtUP4nukM
SBblOk8woI43sBYL1bUtw8c8F9guF3LegNKqsB6Xyxcokpq6hRC8Oud13VThGpO7k20Dc/fsinsr
TXZf4mv1jluQveO7Aj7mExtAiXLhr/srwUpYXkBRSck6H4+PPopp06dBzqvSS8vhb+NCJgux2ymu
Y0kKFuA2NvCaqY4RB29KSKRinYqlF4lhV8T+EnP4BhnGRb0aGBJdqHOkCCkKaVIsUXXZ/gF2yPxU
UFStgFTOT3nDLrCj58ywpL6f8egi4g6WlahrhmlTbxr7nTwgp2/QQN07Tp5+CW2TMbJwRADfTI0l
G7yl4lPu1Bp2BtPn2XI1QJLZtVf3ViKiejcJRSBgZ+jxz/Vhs+PmtP3vJMKI4xR/xOFqkjfVZoC9
mUHQ4ZaBv7mcyCpQiSP4bEe0vay64mCL4/ybNsRzhh2TtOS1NopoGW4iQLnZqHaLHmLelWJeo8xl
CporrE/HdtYSdzQaXO5WvC5bHde0q8EYVQ7vWUWUa2BrIoxrZEbjvgLaoOKTWwKYXfA8H3nsIO0M
mxTogXnM/yCZKkAY/P+BqtiZTKl0/WerwyGu/RSjpUJLvOY+yqHVwuzr5BqYOO2OWVe+mX29/f67
3Dk1H3gYuhId0miCb4Z4ofiXJf4bggqsm2PDyJeUcPYOhXJCTKrH08FvXSNUx1cmDtRxDaKCPHkz
cmA9CSq6xckAVZFqGpzcxVV69awW8iXfk8WMP+33d2YIHta8Z0HdAsfRO969QjRZ9WLhnK4B5glZ
ZiJOeRCMdF6liB+bfgstnvwDME/PFVodHD1tYrlimQ9onTnZeBUnKRytuaRiFddsqGYPWsLquE88
/if290DwLjKw3oTJA+y4tZF1XQhY5XFzWgwUB+FL5wTSoBERKfQXR7iDTz7mPqXSqeOKiXdfZiu5
SpGHEBASdo/xob8BFyPtJ59YeGkBv3jEkv+fVrgLmn2RqOjK16FSGMaaYGitB8rhTZIjeHtJtxI1
7N41KwNnKOIcT3NQXxMZjkSsiNG2h5fX1a6+jAC32LoCIwCt2WAkBSlb+5+eGdmuhBRpz3CW+TjP
Dg230FWPG+rsqpX2UzduXqVgVxE8NojMesVYvl0YsNXUSy+gqNOYi8txNoSig2NSwTB1rByUAnnI
ORoem62W1pq6p3xKoQBPLVIHVW0WUbcaLO8z9LRKG1om1kp37MWykLb4fLL+VDGc15qZdChwagkO
m3YAq0mlBLQ1NZcBi72lVrI/yu9yRD15v3Twxncl0d/mhss+2jjL6kON6AenFbdYt37be8j9vHPY
3oKG0EKnviYeKdPcNLOgUVN0Fik2ipVO85hn486TBvNohWSvGNk0//FxKaIqh4J8kfGOqqJX/+Wi
u37zQNsxYXjYNgzzojEVRqLR7CvVdjiS6+CCioXtHQzHyaTiUfaEOCTnNXGkOUmEQ+25HWdeyhTq
xHyzmrOBRCp1Uol5Qnen/I9ucYGs/nqSqyY6IHvaQzqVy5l7SULd513A+MfvBF+iTsEvDx4vFYfV
45ehwt+P5kl0+6KTm7DaVgXzIXh3Fgzbs3qy2GmQfRzAIDEkKDMJdfrRwc0BEbjzt66rt21e8ij7
P5u6TyMK7DMfYF41/6lNo57Pw2o5A1xXwhLNHrZk7Fa/A2kjbyIGxlDewvUTY27npR1IXGX3Tj3s
Onooqgb2vbKZw7OP7UyT6qnWvshnmFyK4FCQDjoYfG5WWEdApHP3zySY7UJjwbuAwGdsyeQutLD8
JRjz6YLh8wxyLTVSv653VJvujNkqZl3polSe6EJGJ8mvCArmfqnMby6LSjMH4If4Mg60EprE4aEY
allP91drN+WVJfF36KIKPmrI1yXkk1SA8C+SmPUtCzkmkmOoonqnjPKpoOO4sA++ghpKoHQ4AC5+
46j2lk5mw+mIk/UDR05gfN68M89HudY5G9qHhofDzMrXcBOy6MaJxB33L8fZ53jkahCvhT2HNtoz
spwVGlq6BLKpge+cWX57Ssrx2ref6xA7lXbdhIDqAd883h225JMWXCjoIij7PMA9ffE/G4Z329HC
PuNyMAAdOkkzQXWfwk7KMPE3ODqs0FlFgE7TBVmycra3tW1QmzCdOfHpRDSk2HXm/YycbkL+16Al
VebDooDdtrEImvh/JrlI5X6UFAvrL6vmPVa0eJEsVOKsyCZ9BT+eGU2x1qUK/VcsWic8DxJ/f3zR
8W90LjZcwtYHwBsiSO10kfEiMHfCDG+v0XH9+EznKQfxbfNUohby2qd8WCgl+64dLR/tY4oeT5hZ
yyT/aJ9tWG8IFTB+zetxZeWbtoBVILJpD0TV4I5JzE1g9G3XXeGqrBA2hdnO/aca8IKp/j/5vDef
fmuUgraJyqQ875YQDaE7AO60yJ0Kcgq+brNHkoW14d24DTXdnRzni8iTnKL5A5SxcKpInD+a6oGf
KKgzQSLDt1pZrEatRvh7mU2P/ogdZxmL1OlbXLpw47ayWF98TbkehXl5maSQOpBxiA3w9JjnnoB7
cpsmLn52VH0m8xV/HPIaHslAE7OHaa9naGaajagbYVmIrbWhYS0advxuCsBEjM7gMmUXjfHsgZd4
nE0J+Mti9xm1Ahe7S/+lzeblBdMWzHunPCkLDx2Nu4/k4uqHcaYkioEFsiyEMM/3W9CELo6jLwgy
oDj49i7ZNK9/zw1UAOJVoqcL2nyIJ6C3qXKExR+y3FT7GceQiBkoEzgav4W7zeZnbQrTaqPZ89k8
XyeX/vYuDDRvs9prUapqLaouaurnxPADyjU+MHNf8QbMbfjo4F+lw+YkjfvkCsrMJig8ieOs9QwI
jGSaQO/rVP1yOUGCNvCilJ7tq2HnprMtcSTCXaXfTDHKw3xI3FA2MwB1GdTT6Qb1h4EPjkLGev8I
yefzbw+D3/RaiXoyvyQgNuykRhv53FLvLP4gJwT9eELh0uzPAreh8gPHGlUmIZqEmmu3a203Td/Q
SE/NcZO6SFtvMv27yzQsxi5C0Iy5faQeB4Rdy681xMCQPShFSjs1IkEl/nDJ39cMu8M1NZucBjX7
TD4HA8N+ipQJH+SOKktTcr22vED6xGOPK54/CMlRZKFfiwkJ2Rq0bF2L7vezxCB8s8Jh7d+DoJRO
z2lLIJKHfvkyjB1M9pY4bpHIjE3sDOo2XTaIChS3KannjpaYexxXouIBnLcBLApaSL/dRuPMXKE6
G6rJc6bZ/3BTcde7/L0ZK8EsnvjPbNHRD58uLVq5+nPSsEAFnx6WnOoGL8zESk7ooA4qTMUwhZBk
IMTnZfKuq70fbqtFanLvmtDHXpHTEYnbcFEhf04cZeOGWg8jlkhxT81KMBr5eVkZpHMWywY44IG8
4MqvRWZx3DoOxpRDpUlsuR2R3HY70N89ubNCHpq96UBmW32yLoUPez3f37PNM4ut6rI+BrsaoI5i
2qSVnbiwZUmkreoN1pTRNjpga+vgm8iVoj4tVlUcwtWNuxe+dg08wnVqhneIaCPmdx37IytLDx5L
hXQ1kNesirwFQC8pFfrGqbAGTiGxp9m0d0IhtdC9zlIQCF2AF0MTpr44B4Li/CoT2VY84ZLRH0Qz
HkJCN/EDRQFC0IqD52qvdT6hlqYgN5f4AlTVxalITZk4a5Rqp1bwJ4giCvZwi/FxqVkbpCN6A9Ha
/daaIfRU29wt6X3YyK/LiiuuTBQyjnoK1lD7U5QWL5oTAiIkNyIUDWZUaGMD//SjpHbeyCq+qKBc
tKVmPCSxhcdAcl+dg6MBqr8Xs1iRlDxW/8xBKh30jErjNwNDO1SLDyefQhL8JGS9E3+4h4XORniH
UdeuccvkOnFlmyi1pPVKMZYhw5wXlfnMH0iftbwURx0sE/Ni99CIKP1lb6Fw8afpOQ9Vh9rtk5yT
skzdKTdWUybWxBF6JZbFAehyYp1qd+wOhSc18nZT82Q6tMGiYvEigel0g1nMXwZ6s4KKaEYzgkvI
g4VDlI8jDwm1V4YVN6IqsVuN9SrbD7KMLwHTh7hOkewPPGO1eVAniY1UpUDF1uYft6p0k4mSFWmn
mjaBRFZ94Dub75J1//mC8BSF5nS0vQaQ96VtmnF+rVM298yjBWW971hdHwDtnMmozKBdALVii2rE
fN314lOeiWZ0IS7FUOdc+v0VwTH995msyLm1Km4fEsdsPUDBXOxpDHBAW7NC4Rt/JK3u2qg+te+E
E7kcXZsls4abNPfPGkkU8x0ZMECeaZGUP2wBkPCR3D9LeeZlxc4E5wANKjCiTASWtgJSrpriBttu
hlUSUex1aMADxoQdL2Gdv5oZpyB2DDIhTYFfhQwVAHwYcbgf3WCvzTtjXcGEk5eswa1EW6j2Qf/n
2KAJFFWi3S35P36o7+LKeFrplGKiJZ/uSwVQeaCW9DlVz2CTN9q8iKePEBTei0m+uPOwJYem48KU
Rr/tOFQ2D+OtrtwkeIEo3Q38jZM3r3y6LOIa8bjloiSSWHlTO+saBc1+NF9pQmv/ICYrWKYkyhUE
FIdmv3nK0CfBjmfxH8rXxW0IhMyggbw98kdDysM9JADlyKMKNQuAfHSQE1R2SrrZwkmo2L0JvPtY
JGgH3Y1yX6f9zZ1Sc3TmmD8FKgVDv3usCLbLJYNpqRVr4/sWAHGwQ1yLcul7bcOPgOeQrN2B5wOa
5q6ZO123FtPzndtlOJ25gFLxuYjcc5/3l1YEIDY41lSjxcw7OcbwmUOWKkIZMoyG79AX9fvozjhM
+6yyjcRXlNsul3iGbgfDHxPjBVp6SseXy9dSRXts1dEyUlTN5egduLzsAzHRnZH/s6H9oMA02iB1
T9QAc61sBVOaP2oG7idCG+jeUwf7KXY1Hdg6dNCIwsE39vbrXKDjQITAnmRWGiR+kZkDk/IrCPh8
4eQncNcPvFxZTOtxDYGsoqx9H1DVGbxzPk+aYR0yh7Xr3Mmoi25yN00pCRoemg64nwApD37AVM4o
UOx6qghWXqHtXFuKlCnVxtMVaD0N6wirv3zqsO2jU5H0oB728OQbWKxT9LL2KuN4UbESjRzaXwG4
MZRuq2WzkuvQdqUWU3fnIQGqj7NLNckU4PYVNrBhBgArCKZZfy6jox64kj8FBHXf80u0HyhurZXC
omrO95upmiFO2evFb6quX/UPphBveGBk2T+bCG+lcMJiNNG9x/SD27NrLn1ZgrYU1yCbZKtW4Xng
Vi8ayJoAMiCsl3RIipj2E7W89CEc1wV4wAc5PBiHWCxdCPJ5U5xluUUcTII8Mumu4EuxztSe7prj
IKRdbKNABhLDDoYa9xt8g/knfmnzU9ergLfePUPKI4U23iJsMczqAExdokjv81OMkHS89HTQDXg6
1uLHrLgd2/qJ7ogmGUP9wlvV6q/p8RpVl/mWy44T8D2c6xDuuIsrdzbnzpDxwn77u3WJsD+ZrFIE
FCEZYeRpQzm1nYM7rrOKjZBxp55jOIRd/okFqgrg+1+YINdiDeL8V02kQST30eRIazeB4/wZgl8b
rFw+WwOgXthQNM9nexPUVc9g2R6NbzjzimN/JA9dgo52N86g/FZNde2Lh5lBGMerssdAYSSvewkv
hIJ6fvpv5MhG2JHSMRUEigu5DBR+u/WDEGgKd6zNbL+uYUjfVZ5TDmTTN/+UFMAnEn0EkDO77gzL
pYSOi8+OVVOV3yDqxB0RbnU69Q3kIJimrvIdlBYw5nRHRaiz+Sgvict9vkv2a+/L7BfhGdtwdsaB
Gm53lwgt6mzaNWx2hMEEBO1nh6Us+yWOnpHxEdvfdWUe38FMTVe94QFu/Uyozvowb2T1UoaH2HiZ
zH0kwziZubHURs5tgA/S91Q10RGfU6gL+iDTn/MaZug3Ku1rUYl4oA5xkHCRb5DdQH4u3ygJ4RXV
/txZzw9g7vLsD1YCT3IZ4FTKY9xGacDKTI9Cr49KlFNwMrkIPTRtaO+wnnVYY+Oj/DqRXE4zYkzC
9OCwfhmnTNSTRk4D/PNJ1OZs9ZOGMwfTuGkorubBZ4b3O9mgnFPNDl+/1xEDoGfeL1+WTCf96VJU
59E4XBSV7fsnYGU3MPDstUxIsMaxphxUJfxpLw6iSNTSbqSEmv47zzvmpQsRPuNO7gPLpPh4bIly
Wg4hy/dqe3mIdptdstChM/1SuDTwIvqUvDSZ/vlrY/7nsFqljeCUTSMopV8jJC04e45bSFupq+CG
FOLUaZhfbxFkDsYc9Y5e24Hvhtxfyk5sgJn2iwAWgu+6FvXAcoNszCSl2z3yRZTGUkCyvGCl4oaO
2S3VHb2Hg+SJyqzGlT9BcL8dv8lGbS2RUIlVChiI9MTtZq40S8cvrQe7dkAx5qcQTHQ8oqS/Ob3a
Ucyqg6k5PVozi5F0EMfe2Ri14egos1ZMy1LPZ/B0b1hWA1J5t4zCYmKWBQGFEKSg3i8OKfSz661C
wjT/NOyXMVScyTGPc3Z8ZSewFp0gSlPcKAxYJ2hrIxYcSRbE8yQZnzHvDsGay1bvQHafLIPqzzDL
ukhXB01MIbLnpFnAbScn9c3diPCsQGUAv+nmocIkDw4MLMaUfwk7xrxRnM+5bC1l9nZI3dXLWwcM
WBa00otpql2KeiAOAUsaFxaF6AH/L/2SRcNwqnGY8o6oCdnuiYQLxM8CNpas01AG51mLVtdqP3cM
nTG7Q3EtCRbssTUazJ48wpzVttijs8ToVIytmy/3Lxaazagv5bb6qRhH53jignGm2csCtYmD9hmc
P/LZ9sfGQUSCgAOtBp5ydIX8rm3Wdh32r29j0apdKQzo8d190alnjmwprDTt5eQh+laeKC1GxFNg
qYf1DACfAKuV4v3rgO4IjiuUsB4+ci+GyZMizRmsHrUhiVRh0oMedr+3DFAHNwfTG1SJRTWQgrMB
Rltg9IMklNUl/fapmcPiysVwIJdF82PExXeFYIBYAEDlgPahsmowIRYZoCj83tE/8I8NXJwsFge4
ZzmUh1vHtOEQp/5y1eqL+pdmKo5BgWb51Ly7mi5dSUvUQvHvSnczvkSGoqcRt+15dcnLs0p1B4MA
3kB+itlPxNgBsEUosmGn9aTRBjpdGHF2qXiCc5Nhn0M3AM+ldg95cLBTWS8mR9Gxq41lDbhyBPzz
pxT6T+lbh8w0JFebdAGuCD3z4hYZCAtLmalwiCRmbSwc5D/QygttftGa7YadJnq945Jksji/s73R
OBeNhKt2Q0ZmJCghAEDfnPZRqDnuiuNMeceL19THt7Sm+BZnc8ouoI1f6HEMrFEfZwtYaFG5zQLL
nl+Jt2dcLiyb+ltayarKKnbPrRmBfeireYy1n5N404JIy46N33BIIyzDr1k9RprsJxeEAU9TX3lI
lUHPMdtI+pJCk90Sk6raL8LrpUCjGhEA1btiSELCgT4WZUS4hQGySIJD4CrZHLeJhltOqg+mUeOa
umOKF3zOTbhwXDYIlex8HAn83V/TjtEY3C4Kj0rB/tZcIT/YQTN90lRB0CLPVZsCe8YcC2IGSqLG
I2f49q+TvXsazmNNLv8BHITTNj3y4xKd0Bh4BNhSoWb/sQvhQOsC4mo2MLzvMXh98wv4eN1RQSgL
5h9HMWib63sS7WorerQ1XT8j3ZnKJkSXbOkUx07GNDjJEjnpEaNac6iaTGz2K5t6HgJVPHI4fN/W
/6hes/amCnq4bB4v04ikCeN44WVzfqtDrwsnAFxSi1EBc0sBrF5Lh+aji9KGFp2NlB51YRYpzkYZ
0cnNp3O50p4Z4gjtQJttAHxLf9Asl8VQoJB13bDj24zup3FRxjF1aWBlP216KrH9C8mQ9ZJjR7hU
4jCQ1hArhqIL3Avbox34q7eZb8LH1OtRmxZ1X7zEUHd9Wx+2PG+GDNcjByqWxxlLXLRO6/SESkLZ
aj6qT+R6y5Bg1McV09wHr5a327e5BzMmeme7L5pL0q+aUj9D5aBbZ/d9RySqYNFmDGsekmyGPNr2
dANps7RJSYzagufv4LZl1gWh+yKrr/88LcAZNd3foGiCb5sfQ/PERXevxc0NtsnietUckNx2LEhz
a6ajlQpd+YaAUX20ycCmuTHoennDKtNAB0xz9UnYDNq9BhmXX3MHpxMcUPZRqt4C72MLQGK1Sfp6
X9Lrtdk01ttuwcpjAjNPqEdLDbFm6W7kKgv+TnANXODus73KPLgcKo4Nf+BvW1mBWO7dHNH3L0q9
uyaCO4Z+npDoqUV/NpEOTSVJhC2vmmtDgjE9Ts1RpdwxpcdMs/aEwWYyFiEc5nmntUl05sWUJb7F
Jb/ngyMAILVsYaB6WptH+D9I9e2kVZVG9P4eTj5MEa9XqFHJQv+qllHIz1FwCmAOyqfd9TFgTtPr
MpslYeaqH2V+lKuj8YFyuFHpSaWCKNfqLZO03IDnJ4M/3qpZDSLtWdmd3JLbQPyvOpofWzy5qrOr
RBFbslf5RqJVSqZiQHKqKTpiThY14qoXqOV3TdEyHPMQ42JRXNdTCn9/P1e5dSwH8KlcWSwyGrA+
sZuVGoyIEuChQOJF8Ryome8fCmO4YaRLXU9YicAMpJOoi5ZQ4kS79Qi6LiBIwCocELRM1XrkdIi9
si/TF4rKDe0clFX6vxZDXAdeyEGp/UzltJzgHhxUCVjaZjCwB2HjmC3X9iqt6hVW5bUmNx+4aRxK
arLUkxizBz3lDk7dHdSVuj/jdXRAKYorl7Cm690YvecuPbSsSvQaJuaxEpQ+jztMxikQjNZ4qg7X
Q4zPrHj1cWqaZaZatC+UpZCYsluPufYK0TxwgLqIGuq9REeNs5BPc/qYqfelPOeedHWCjBFcOzx/
+eTxF7VRd/FM+u3Qp8Jrmwn5Oz+3aUUqwytg5XWv05u3BTCd8oi0ySd7LRIAyZgHo5QChCaBIipw
SLy5HffPtj3KZRIYjgKADxo1fP0dLJ6YqBUthYbRXO3tp1Ykf4yyMSLTV5/lO04cP+aGwKv4iQ+4
cyOmRRKOb3Brhk5kcoTJ67tB9ZGzCFb0HcK+UOIJPW7yIGoMBZncTtQxV3vZBQunFMREXWu2vYhP
4qCUwxEMbtrPYVLobWhVRDyzZ4WINQ0T3EsLim5g9tgfbCmrLUZAHTPT0NeEjAsvrNvtsWsdQcxJ
9mIuSqUzwouF15AycCcBu95tWrWR8xwtq3xylOKTgI8oqMqWixWtaED5veId6kzzCNEzkWVQVplK
GrIu6k6BOCKZtteFmpPOSN3foOmxgF4Jc8e0YOfaM3SDxhIXeRyUMy0enhy4Nim5YBnMu+LlRXdw
RMbVTTiuvLEcLpHlKrodyeIcEEyftepPwnXmj6yjPNtKiabMk9Eo/XB+OJ4vVbquletfWtsLAZB+
Ax007r9fnQPq7SV8AMDgrhXT9h+bu+eCbLAUqZ7pPvUy2C1+D2bvudSzwKnLuNCiYSqGoPS7THPw
+Vtbqq3sUHknRcytrn4/Rw5rm4vr3YbZi+Mmq2hvbpWQU5BdvZbv4D/nw+KQ6HqYlBVve0vfjie/
OhwVTVfWKKiPhqo6CZ1fDURDM/TCJq6RWtpm6Ht+SDsP2AyE220JGwv2LSS2OtON5M4WrX8DOKtN
vf1iP1ttTWNKMdRjaFW30PiZPCibDrCn5vrdZXPI8Oad6y/yk4iRGL+ZbvabQRtmwlPMJBrt1HUI
yUIRwaqjKdYRYJgjY0pDTxzeMcEIRzdKSJgvCXm8xDeYTAwdx84ASEf4obHj+Loz09Aa5QPJjVne
WBdxRdJvILyYtLy9ZwkUXYiKDlBhQu9DvcZyl2PfzjN+8rrRkEkk1zkshzI8CgsTwQjhkjzjM9dn
SgRD2Ks8qpq9ERPopeTIVjnyuM6emqEUHofOXf2ktEwYUbiM9QX+Dgl1ib6JgDsDp/JuZUarw4n2
jWdHJ1rvq/6nEvgZ6sOhXbLQvdPVlNgc/cTNVZjA0Y8uwQ0GLQSayeOw07/f/d4MthjedwTX8mqt
1Ou0KY5wGQJ3oqj1oBP9VP6IXxc97zh/gRpZdHgfJI8CP9GS6uyUtQCAe8UkLyaJvK6JfeNE2ejI
cmaAIFagqh7Ckc6gbWS+YhOj6bmPsysiU/zdyM+8ox+N4excdn888zEQfnqqNLS3G0ccyl0DrpCe
UYZAEe1H3IsoG2alSG7eIYfZ4StmbHWOKp62Llno/cnOZAljWyaaq3UOLcISvvAFax6mLGjctF7R
hugMBr8BA6Ynj1343/9+bKB6cfXIZxacsl7sZKtIQMAodeua9s8FEvttRqYTNuqm8xQC3rH70NEZ
FPjInk4hQEPS62SHSMrIa3aChZXk+10p0Ke23peg3D3WlR3LPCsB/sekLDW+VeXn4+EgPnu9m7Ay
0IFzzODRJoGAhEHfit6itkHplWNulIt2AtlCKUrODBVNQoOcLF+E4P7XGXv40vvJy+TKO53Nk/xf
l1mcDSNSRAnR05qJkglw5nkRAebQknLUMiJUrZ/pUFgamDi9mFI76Nka5ZlQCFLUzB7nFGa2CBrW
PF4vURi/bgiziD2MTs6jecQ67W0sz+JWdKNjCNT30OlPvwbhTMXYW3x0wdIpz97BT5cMwr/1QxEc
SzogYumbSHzH+Ug6rsOpS1HrrWYEX3wJILvZ+Sej6tQAyYeTN6OJNfToR4PDXTlPspcRojJ/RJor
I8OcJvGFlwijAOFgjbYx+Ge1E93Ombym1rbWiMNZHda3CuImc1jvzmzrpb5Kq1rJ4VHgNr3RK9DE
hJvk9g0xHft6EGk4p3pZkmOWTFcs91lfK+XtXSennknM0R5ojwTQeNdmXBp61rH54dQW/lg1b2JW
s/AIgAKFmGgL4JTHltvyqsOyUa4g4LNiJrwXmm0ZorrABQRocghWLxCnLwpH0kffomIbDQUX/FSr
GaMv4FNhAQrhWWemhNrdVXJ+RnG3+oZXn+3uYhs1H10Eccuy51Dxl4Ym0ygrcf5xCWxHmdPtnDv7
mDH4QXdpc2t8ggvrIqOCzQpeE4tBLX5UES/MC3D2FGDqvl4kStXGiJ2bhaR2kP/7BcvNACNVrmCr
dBifMqXuwSOOVSFlH7/R50OzEd3T/UjU4XauHooguF/pF1UpmvSzzZOPaefPqWNRskpsykCU4MWG
PfcZlfcjss/5Q9V2UsVsAZ7P7htjSoNhsVzKdQxdIUkqsCRwPFG2pE7dvMS1aPC7vflzr2PaVBuc
iN42W1GXADjL0F6XJVbgqnh6gpgKSwJIEdCF8nHiyvgt2XxbobHTgsbgm7NReLVKjyoolhKmnG9r
hM3DrQzy/z4GBIjEJqEejBJCcwOr/8fdbY0S/VYIWadRtnPCE/N0egEGiHtefsfZ6YlcioZDnFRq
JZpVcRe8LfO1kjyGJmH+/D+P+hQhQAF9m9cSTgIRIkq0tWcmFEaAanupsYn1jUHpvppCzxU1d2PE
H+qZKUGj3Re7xbwbaoQH/DlJ9+lYmJaCclzY4ph3aF85NfIjvHlYuKL+uNyuDEy1JKsW4RP/2A4T
QmTkT0ZAuP/zKwOz1Eldvw52phj0I4jWbz9ufNqfB5AOJD8ELHryvj4U5ffrT9fYdJQjWK9bra4b
j337X2HoIhnToMyew14GxY+O07ofbUgK0ACE49Cgct2aITxofXUmlf2YKbFnvyfAPWMdhg80WUP1
jxFg4Tl24ckW/MN/Nkbtp+HGtMENAxHdbP92qii3+PAkk+ibplwxwGtJ2W1Q8NZ/S5QpAbjvCEap
aWGwaDDOHus0pZL1lV412WwsQBy3xhED/+ShQ0z3aKb9Eq6GdzI8OYNe34p6LM8/EOE2Ty0mCAu/
Qc7aWfWzcjEJrnGXPT7uVh5+iZG+UXPXxLEyCxMJdUiRd/qLqp9Sc137ODgpuzCtUpAiDGEseo85
CJ9RxlT5C7Jvtjbl5ui0GAHfKd62aUl5VQDmoQhJn1SXRpFY7Nop1A9qveZAN3hCQbdt9SQqWzUB
AGIksEjGA2CJ5JI/vqdOp8arlG+yeHHnU1isepuAPHI6VPDxsPYzEvECMfTvTI2Bc9y01DeYJjtU
6KfMN5LeIIXe6uQ6qsU60foeWGaG9qxFAr5Zt1EIpeM+JPaEpb4UUrxF5ehuQ5uCohPY8kKGRYwT
JCfrgX1WcR/nSrGvx/koIGd4lwJShDlZc9Xy4Pe+mzooXLZoF5HDb4KrzqjdfO74WFh3NfYcSo/Q
3PG18QfhXyv8xskETrWZ31Ueau5HM0FOeyIKhMZoJjkE+s9DQtj9KsPNpN45Gn3fASSkbZLSSsRl
kVd6Msc4ZPD8Ebk38gbRpvaDkUGIDehV7A3QC6Lod4hvqbrfm7Qa2sdTeXqUFLePkwxjcPSr5OoX
lNulIUDUdojs3QWQRMsFOVCsJWFt1KPqXM7JO4iK9V4UwVWXp53NJgblUyI8bcyadwDJf2fAtP7M
l/WMCQ88sYTJD1Q44Oq8RRoffM+qv4m8qaS6SMxgVflvp2H3bAuPRgA6eISjwGVZGwnNvpwrRH0z
om1WCv9nJywG46R5sJnTPVbHzVwrkko/7reSTRanMsNnqGHxoVsuumL+rzNDkS9pi0+s+YoSeE7b
tw3bIx6NuSuJJtMoI7A8KRHo77vtQz0idj4y1ldEZ8t2pUQ823uq/haKHoA9cMmRYSIKU08bNjVB
AbxW+lJpOupOJhR0/+RFXfLJrnCgIoWs0GRhPD45I5PsP97Op7IFsglMtmbwuKuHUnbk2wwwtC44
0MNrjTdz8wGr+Q118Kf0DWVe1GoZMb8Iehc9rD3cFkWjfFt1MMpQUCEn0FQF7BaRDd+BxAYvV8rk
Nw3CLrdUPJLPGk2KrogbsyL0h4Z4vkWgbnSx9jQkx8JternEsyLYdrogXTvFSToS5I9BagbHGHAy
+p7tUOublHTPkqGmckEHMpZQzsMxyTtGKowfiqq7wFByuMwg1MMsSdgmntXQlJVH2fa+mxUP25iO
IG0wDTcgMgNsdJQwglguHxmFHHm9YC1+dEwDJf97wfibXXGWFxVP5+XlitX+rZfrNoCGUrGR6u+k
e5ho/ZrKBt+Qb0zz1nYvI6Nq1BhbWnGOGX8OvUe7glFIUwAIwFBIU4959mxBpypwy/rsgrtrnWES
0AvGU/J+zmewb2gzhMLFODda5rjv+97RkI4gA31w6Zl2jiiu5MBy6VqJWQtpLjqvE2cY2vcKmYC9
BFkwkESnlP4pDhrs1bHs2blzB1MmKUnC5lwsys6zo0WAsjIInK5NWY1LRqJXt7iirPja9l58BqMq
SUyVQqxO3G4zAal7ea9KJxDxwr8Tqt8dG9r9Ek7Qx15ZNmx/nvYut2cD7ANmEDPSZ63MyTqDeZF0
gWlV1z96BWqJU590+uLYGseQfmbuyZ4YOisM/zgCSso+GbspiuH2IpPGxk4D6chdJ9GVz1dtcQZx
VLJ8rM22DwQmz4lysV3AUopbbYXnE+Cm1j38gkXX08eHEvqtl0XAAuGO1qK6fzGI46SlHb+cOY8s
f3ix3J0L1k9Qw4kvjmYtLXrkM3/aNtXJ6GkLXB88BTkVM8/euas3y6zsN4qeeJKqdM4c1BvVUGkV
gP2JaATrYdebAGPTHcn1lYKxpIJJQP7Nq0unYWsOJ/qOoEmrPUXRnl+OqxvFtb9LqDbYPeQiuImz
XesUhCkEKgjJTHMEHUZ5Z8uQC7/fpd5b/PDAQFcKJdXoT0rkh0R2wZhcWxB/5KuXggMPzyWwSKbu
C0RhkBXOdx9ix71syjbSeCUc1Sr9AGBHwLPyrxNkL5eIeO3EP4p6cYBv8iMA3qWYqGyNu8E9NM2c
rC3WL2CFN9+yFNgQ6zzAKJVBkpztFR1gwPjW5Iz8DTjOKABaBFDjvPA/3zN7IzXpwpUjXG7R+MAV
PaRUhxuAG9ar9j5iEdKoAIKAwcunFd2uIkz0eKjY3aMNFhUiDZqRKchkmuZOrYQo6x+50Cnx3ifN
s/fm3fYT3B9SyR7I3t4vo4LOYQRQ5Odg/FUjA2NsnqXV69L62nY+vYofju3HR9tGb7uc+2MI0vMF
yuEmdqh0hNU24pRLYpVIE2vGZXmZZXHO5UuHL/chral3xWHtxVsi9LlI3vB9lJLMhSokoMpLRA9g
Qccn3svru6gJB9XBrQtr0N8UhEBIv4ixlpuaPOkjzSiwg0LFWI6THGRgI0KNmgCH+fQ1nY88eyh1
GWaCXb2xnmCoMc+zgVXMgUAnMYc72LjqlH5QDW5TI4qfdOAhb1Yk9ia6PViLHJHxtB3amnLFCrDx
sV2Pm2oirCPE/puP/6MKGpH9wBA3aRLfL7YrCu83loOwFK2N1cDeEWvtNnSBqlOIvWKPkcGmoCCI
ET9J5cRICco1xY6wERvRSmCKiQqDHz/+ZbFOnFHVchjJrSkf2QlJ6cNwfDiK8u+KmM8D5h335K6l
Fg/G0Ry8ww6/Al/vd/gZlMUTjX2nFzj7nWlvYL51Br4sXsHhEZ0OeKUCF57tOYwVHAUl6u9yXOlM
hSkttMYFTTSKYpbk3xmQv6ceTPaeambwuJwRBqkAvm3BtxxNmL6vY0MLbcDJGAYhIi8kmYTHlqqX
zmKhlmDq8D4N0xtdhiZmB84kFoLKqb2mQxbRixVhmU78DwYilidn+hALuF1D2+VdNenRMO1bV2Qt
m7O2HcE4yxwN+bTk2ckr+qttfWt7cY4OgVnYZK5mA2Nv7R4R/Y/i9qN4lUZJqrOI2HlHrFxVT16K
vbryoAK2D4pSFnJB2WbKHs7Yp6Sq4YJwcoFWBI28etz+4XGWfVyxjKlTj6ZRL1WWvcpwRrX6VuXC
TwWtKZEn/tc13Ng+RBF3HpZRxq/BAM4gyl/5C2QD34ChszJT/rmVfIc7v20QeWOHx1dds4fPz1hE
hpGvlUPM/zZT92B2IKgqNC8bcB56o+l2eCpAkwnL6+fBxmZ3CeIz+Leir9WySQnmoyaz7J7ghUUl
YYgd+9jM/oVIx35yvuHJaLKLc24SwlknnfC0iL4qE9ux0qdNRKXg9j7W/lWDB1Xjk3lOEYS0jBk5
uaGqSsAXfI5QWWahVAg4Wo2XAx9lVqJnt3zpLwjqt9zFl6FSad1OaQ229wXYTZGwZJwzWNoQl/4j
RujUrVRlKhhxUe14+jndqWb5QAEdQs5A0qCIU9ze0kIh56JhXuiIl43AmNsmrpnvlyHiVZMrbyNL
hyLjbehzIo72hhfnTfLVf4/PyRK52GSJtEfgUu2RZhyipWiHrD34jQ5whQF4yQKl7DkJZvoolB3S
CgEWB6JsBVUgfytdom9dwETFxW6p85CqjpufgNHs8MPKGKnujVWOJSbNtoNM1V8qFrxpkHOcS8FZ
MgFfJv3Uj7tmUSv0l4WEgEF6C3QujEJ7o00vda0RtsLd2ep8gtjGCcJkQU6mzk3zTicp2e9gpFyj
qVjrGmHh4KGzFLOFUp2HusbfHM+Gn7TEM4el55SgMnYDVD32rKIaaSMirfFtJdA1cwDtDi1oOKU2
DaHTYlu8wNXjxLJwXwCdrFURMqyTZ/L6LftT+kEFw4Yqm0Hym4+oi1K9U2GcHMUah35Ydyd2dvk0
vUuE17pSDZF6oPA1U4C8T7Y35sU/yH/Si5MEeu+Gtg6lWywskQP8WVpVzsSbT3omjW955mmVWzDE
q2s5Cf9jFLLiWVpwoIkbyJTEM60EAUNtSNdYBskNESV4D1/nOJKEs5BxoRt9miWNrZjYqs2F5kaO
/+0nR5VsdNENtvDVkUlgKtkJ5/oookni0F+QZd81Q1yrN4cDjFc8uidgSSDi9ZMxfG2c/tKPoJQd
50LyDPyBrZxCdzFXxObjvKU2rxcEMJ1yuwpF6cMwNfaV309ilXkB0sT4uugbY4QYMn6ITJGVFNZB
PH5e0OyNCwo7GQQFvZWTmyBDELIn61DjRPUeEr1HUdGeXc77NhQLKRZOeweCmGnFJItRy36ES/xD
773Ny6doADxMWLC7sX8NN4MTmN0xRNLNLZZX9S+xhkgE/ze78Ft4MWH403Dx2SNCa+2OeP0elSod
Nx292FTmrZ3Y8mKhy+foTuKIJl+ZRoy1B7GI/MVyJR6ekBsjPR285aVmtvDMPukz4XF1hZxTiKWF
5YbUsATn4qIV7thtEHwp7AhOGOXCZ72xJSn7qw5VshD5FY4GM41DOUEPyeEkDqsZMlvt25xaHMSu
aubuD1e3eBZRb6KUE0TqlTEB8LOacnwcwr6tXNW70f8c1kZ7Wl5VmpbTE3601AwCRlIWWM5kqu5Q
dQuQpnQeGJZUChDfrT6d+c6SsGGV32zm66w2prIATaTw0XRBVIk8IoWia8Yaue4LsDrhAJP4q1j2
/1M4+F00T6iuxkMCQrEnnGBliIEi9HZNF0+21WKWymtgsuqOtlgvxaCDKA9qlPItkPLHJ5FA4ezg
WlkRcsk1JQyh6tZYfdxo7Oixg67uIPr8AWLSMVnuCel9fECnD0EGtZnQ4P6WM9QWdzxtg5y+DE74
QhaPUR0dWgX4vhQb3pL1Ut5FXdLUoGTmGOQFFsM50+yd7IRHy+YXkl4LP69GlQN+xGjZyWXcZMaU
XrQwOGEf/BhGLCX0mMqsYMHd5CjuvBeezKwuEwUXL6fNWBOulTgSqWQC7qq9eOqFl9HO3IlSR+t1
ZMMg18obkzw3J+KD8sGpBnsMhVDgeA3BBJnjcbKo3cumoGLj8PDI51zOMhsuUS/i6X5T6HGp5D8i
nOGcE0GXbw25iNR/qNzdQTYj2EQb8wxMnCj5sT4FCqRhyFGD5YkmkdpUm3s/jIELgtA1O6/SbTe9
ne/3j6Hi12DcAaWoDrK05z2lCj24b+DxUHXFimiOg1CYFDjqXtdsOwydoi0O202l2X9mAPu01K8m
Lyhgix5DM2fXspJ4HFUvS0g4qW1kHsHJqMhuCHBx1upg0NdOlRHaZNrnBGAO656Avc2OGV8WbLRq
5T1h853xU81o9bcV5OPjyODQD/tXhMXr+bsh3xnWHw2u7+CKUXAmip2J9FclYxyLHVGy6KLITOUB
CX5zCo0xe19Apdgj+7tnI5FafYSOXlQuFlyLrA6u203n7/nuwjlH20HTiIK36/omQ/DizODxigUX
HVR/Zi4Xr8vnh1XAN6P4dSr6cy7sd3FDl3Xpvi/rv8U9Rl/RqZhpsnq1xtkNSmg7jFyYGagBv73P
cDK6G6IaEcO5qNWP5FKXCTLsHnmqbDNLwCZfKVexeQzgpZFo2AbKFhXapir7GWuylRMdRuZh7bo+
btfTOgzti+vWK3e1FdsjkbPvD8BGhfNNVU4koud7A8tBAO5hqmd9ZjN/Y9qAe9W4zHhvVBRmvozk
cC3btBui61YVjTLR3jzQZnCW+AhNypw7bFOUISK5kt9UqfjPFtb2ITXQKrGibet7HeA8OvahlVug
DUdRZ2Osg7GmD40MI6W044WU+D+iySDLKYdAUka4WOHllz3kopW+DvEdeVa8NE2F1NeMesKllfLt
lHxGPNlY0Nh4Ip5S2Bc6fTigRXus30tQupZu6Mza9FSR7hW8O+ESMfMhK2WTq6yvtBHNDI05XEGh
o81LuLWtjLjiiq40Nqx7lWwwziJ1wCXH+AUKaS6SRhbfpgElXL6oPTLPhjen3zyyF00LICGM+/7A
oiPf4/dJXNG9PF+0575FdYjPxOcKtljH9xnV+Okc0+PluodfZHkAczqJsVrMV7HiuvtsSS5wB4PC
n3pxgyuwgAsMpneLOoVIfhUqDWBVjfXeE1XT9Mj0203BBEMxSKqNap3HvFD7Jd+xpdmA+HuZukNs
i/8qdwxKIONOa5dz8h+xhxQbhbEFimU+Q+E2NpJEUqqpF8pgkfg8JZEqs06/gJPK1BC4Cfs+On4v
9YZ0ULawn/337kXHSG3yAgzdeoTVBm/NuLsiB96P3e0YyNZeIxa/0rOL70Xuw1OCnyEFXwdUtf+7
cMybLmwnFv+qlzKtAwD0/E75TD4lLuNAwTWPYvIOkFxgFO9Jwb6Djck0kcmGdnZWuW/bvYkx9tyS
5Tz56QfjvORUPdY+On4JjYW0IrCH/CtyDVXR93F4xw26Pwc01hGXx+Ji+X9nD1/Lm3jb73dFWFH0
Nn3CwdtgSGdhmBKdg0kmZZhdO4FUPm98twAzM30yO4ZA76MLRLzZTNW16jYl8AoOVbCIhMqlxhoD
Y55fXROe59g7+ssXV7iF/LmwxeowvqXe+RunuGU2xlL/e+aJO1qWLhNcI693hPfc9nSPXNTtntXl
xUNQAD2h9N7qgjdrEPrC1QtvqL+nyJ9z8hUZwQ7LBFTnYBiBWb+z1lQPbJbTARFw7eSFcP3FZAd1
JRiQlln0g4KnogZX5wf/yUY2OSvKX4v17VYeyyoBOkcIL+f6OVS3UYc1INoMA608E8jdMOIQT0bX
P0Cv6Tf2QYBabUrRRgYwF/EImJmb684lWm1j3VHxgGf9T6jU7SvVdZHBCTe8pVi9WcuEEVzEFKtD
jVXRHEVg5aHSPap+U8uhur2lB5p1gYZAINaastX2u97JWlG1rKsR4zKW8jZiblurzXBoZBuq3Rez
N+R0cbZNjpXMTR97qX6EokSTRzsYb5Vl2Oj8QBcNP5IHyEKqlHaTfI4eezcQKcHwq3Q1xVsHgurx
Nu1JWzqLwUEA+i3vqqacAo8F4eC+eT7SLPa4Fj/NlDBKo17DkZddd+57vKCMTZmaoTGZN6CvceqV
acDzy0mk4mwAizjniou6FV/EdKICbDUtS7LQwZouHZJ0Aih4D27+ptKbu1gS5AkGm7NGETN2AL/Y
FvKkVmSDEvR9CooiwioKjQgVvdkdopIyrPtm+jMbDKIguhhhEWBaTNCm67Pq8+3Ncv8oUMpiv6ny
q6aYPjgtkFJsb7KLBJsuoozX7f4RER0BnhDZh/L8Vfe2z2mRPgrFmt05Zc908JJK6FYZJHpsDlF6
cJ1XFjvmxSFIAvtS8htfIjqQt6Xh6LfUPz8mExg0aaTFUzzCOzealqoS5ZQMhj5jGtM8R5zRfrky
Xbi/VS+FSPiSKnqHAUhCtLXOr4h3Ht430eWDNjHiRlq+keGHvclrqsY+sXj6LmEo02bG7MQ6lL2q
LpFKxB7quImmHaIPHsTXdqBZ90guGsFVaC4noXap944UjPrXqhCKftOPN5iUk1AbhTVOGZV4mf9K
AboJbij36f8mOM8ashtXIMr8YSYflH2EoW2EZaNDXDnkCALQw/RXn9R9xyzyrlpChZdP5o5+uoHl
Ik5BPHGIaA05vw4v2vjsPoAqSdVFRpzo4kuq6c13CZ5eeh60zDUwsyjZ1qJAQPbMA8gXQITuP6K6
XuXVlOdPfnuCfjYwSg3P9xoEERk76pMU011Edlz1RyY3K8IUBYiPhrDw8E5Iz0rH+E1DfO1dMwGp
8O5t4y7X1Gn/Kf35fWfQmcDH6pqf4l26Nn94aaTxszSkIKTaLfUYgtAwC/jHLoZPo8vy6irhGHuM
9IGgl9kWAzVCPpvepz3qUMEn5Nmpw50lMEG+Vz9tsZ0uG/ESwv4VJO+PfMNvkVvJ1ogNaR9wCT84
bi/b38iewpmLWUzO23gOSsWUyuNNj3CqdEtdF7fJNbFSDOiAqghihB53aOJi/7HHBPKv1mQb7zEm
WoYad9Gmgl76tZMCzwDyQusRCaxK/1M54g0tz0DLWfOEg70c1lLEykp7zARqCgCmELhVvfuEojxO
Osw+z4yIKQp506LT1D8IE1iRTiG0iU3l98tZtkJjIJEzTxEKSIEVbSUF4hs44wgMRFi9c/QL+Im6
sq5rYcmC5a0Ewom2cFndgHXiIDw+x4TzOsuzZiyftnQ3UuDgDZ3eO3YwLw6igKCFUCydUbBCuMdj
o55eyv3kx/tFLwoSqCFCvONrLUxAphIMOkV1ZhWBgwD8NqnFle5NMmssDTNvOByTBD6d9veX5Oye
4Hbzmq49Rc9iNPfK4xloiMaSEq8PXWXRb9CxtMfTeSDvHDyuxRucfKpGXcAvvvFhEx1BBboV3YFr
aYcHPk+1t85PFZHPdnKnzBekzb4HyZ6bGxfvJTs9InlEcst72xxe3tELiuJI/yq5OgutEKFlfJEs
u1iysdARfFOTjk+l+OXSl40L1/Rq94WpH9GCAKY6sebA0khfm5B1FBscurwq2AR6s4MOjBDK8oLE
dyetD01azvhXRzJtTu4uUUyhDHI0+YRL7p1SjvMALFyd5R0FarxG72xod/BAM31uQFX75jvzJ9bW
ChZ9DOFedcKc2FZoPBif2qDDst8pJQ1Sk7mWgN1ShICqaJjYXiRUdf6PfFl/YW555eLt+K3/HLZg
ENKordgDy6Fvztz6yp+2orCCOybYahWp2nS+asCjrT92T9wXVMDVMgWUHL4yxveqXZjzCZ4kdYa9
baup8oG2KBSHO5f3Sm1OBX0PAN4bagwmD7JFVTuR2NlmIdRb4TgfwWT/HQv1y7ijGqFnRps4daY6
o27yjClcXvg9wH6QhKcTfCma8YCPkBgjQ2k0jzfopMYCmLkiXdCBZTJ4ZGzU9w2bHSVoakUBF/0I
cTAdGpNJFP2VYQQNX7RAgF2HRgGMdWsO4Q7+tDbxE9gsAjkKggFULwzdyulcXDSbki1pKsT4mHLU
7oTB0WKp7PNFllOMkZZzG26nTv6G4zSoIuc5tTEAqH1it/VQcj4AZxAbiVC0vdFTRn1mNpO+Ema4
UNeQWw9QjrurwiQ5Hk6UTNXVWKVR+YOCqkjyh6fWpSHgmzuZ/C4howRjF08xfShqroNMgXB3UyBS
WPw9Lbf1WioeUvAGomD+Nxiy+AC/quvRcZKNsEZqCUzZMbWbZQV9Yj5cfA+TVh9/jD42Ckq03cY+
hCcnh4I+8q02Nr4+soOypFAklJXaGphRuFVoou+lGCwPj1UYzs1x+tWBDhgMoKZRKZFExw7fQW4S
6IPAV06+mutamNB4jLb4p5+2CWSeJbJmSOLi+JyE2p+bWTHFgAXh8cFuRaDKSfLz0MJa2hTv8kMw
vmhRTwnRhau7V4kSbBfYmicb8Z5ztZ11nVEbWEMyfMMngxwngCZTHHaAP2qzGNsCPh0D/QqPEJi1
PqwbOvvY9k18dIFiv4Y/hyutYgVCAymuXFG7l/f89m97Nz4N3cySnZr3qRWmoV6deVL4V8Z12UjE
1MuA0P7kFQZzamQrTfQEFpBPZsMu4rxW8p4vwlOMFcPQ05JaY+RfrMDoXLQ5FGLIchNKBSRYsCn0
L5mWLoCpKlr0zSP+1LpRkQJCtVbonW/yb3dxhwbSG2c1XWnZ8lMnDlQIgpWDkTGJtM5FfzteF5g7
GgVS/+V1wBFts5LAhzWEPXL8lLEj7JGoZQjsdANYvRa7viwdbr/hDN3+l1fgeHpnvbtEXOYA/Xjy
ER7g8vnZ8OfU0AnJkJJvMAYbPKgGUpRNbwc0tKggqSADPIohvoCBdifzjjM5849bpHXmBcz8nJiI
Ki8phQK4xWUUNywP0yNSITgnhLl218c8bxruV/R3K7B3JwokWGVhStFE0FU7iZqYqFEqJRHhOwVB
Kp6F8/qIo4EaktYtUCqFacfIIlb7ssewRVhP+I5DUT2PaWZlvomHsEfUDsCow/remcSChORtLdOE
faLXBmcbkMdzlsdiWGDZyIkMy7VMmfE6LNvfY2i5ujwIh1w6uSLOOY4mv9Ull42PMrFIj3NkG7Cx
DjwZmJVmU7GqQa2WkyNbimkyvUf0VcshRRgxJZD3+GFdiLCzesnChP5gPnaiku4CYuQJzevho7Eq
/6YfUPvpo6RK3RAnE26LZAvXVSItwPqwKYBu20dcY8Onb6L5JofGhDUsZlXjJdNhBZaMu0sL3kPE
kMDg8Bk4M7QwhLQpICGIVVV8IBM/jg9WGBvGYJclbRJt5K9f0ndFV7DvNwa9dlbH4cpw0d/dRQLg
8ywNrMWmj9gnOJuXqGBRDEJbTdyBvjV+r/qCjxOyR/p9ZszWnd/V8z3h5UdAUNjdpCNZMfQHdezp
88Gwi87oaSI9+wwMSSSExpKPfiI4l2nPYTwbMEadrVDNfd54XtOs1dIuEd2xA5dklpqgXhshd1IF
aKqMYnwpnm6YftP8Y2mjjOBra+sppnHN3ByZXjLaUxuQmzJMLCiUTno44LW8hRyOkGf42wY9SNlh
o7P9U6VRT+ieKbuKuw2LAQu+fY2+fTJnY+aMBB9eyeiGiodK+mPw5Lp+wH1Kkf7Vo+kgH2lqMGv/
xz+8mZQcKmnww8o93NehlHLSZzB8oXP1TKx0PZV/PL+i8Eq1/4z1j4ZzRaqR0bHLvGAjWaV2n81+
RXwflWcQNv3/jBe0WVxDgdpjUq79rlQquDQu87cik12FM1mPpM6yy6jNHfFJDRCW4lJ6swZ0jziq
wjjKefN2cWpkKypjdFw0wGNoGdQ6Eu0c/vrf9Xx98JvHRZdJ4LUfD5gKWTUvfODJ1fDY220KOFaY
ugxcrQgtNTNhm1V7OUHPApLDbNBNpiHmC6DP1mwmLSM7ME25AorDXXGheGX8uTX2tf55AhDfrUbN
8qEvHMZqjSi3i6bi9FBSqkqMhX7XzOM+XfNxIsaGfSvwZTbz50jdeS+6fFo3xGuhqZSbvV+Z2wbp
9+lHJYPlQCq1W/IrMAK5A+GtAKJ0XRd915DzgFH2VtVXeLvZYHHxotm5FjlBUs+2HwDrfhoSBgJy
QdE1gVF9qC+ji05kKcMvB4mIbjjKpwq1eTV1fE68TIUSAalhW+iD2bW521aoZoEiPhGZs6uQ8Yy3
H/0R8g5RVUmUJ/gINrmDX/a0uxEADxvNS6TW0XhO0vyuHK66wCVl2ZHYDSXCLAjaHMi3+PDUz2tL
CWdcHJSuaqCcjcSCDUYMlJUUMeiBkNete/mbrkY0YaGLqS+/3ZcMk+SfgpVuSl4b6u4glisA5C+x
FfFk7TfGEZzojRkRrDDu+lLIl3h2Fqy0LCY4oYmMJt+xxZi2p32OwTvj4yewUTJ0jAaiYrGRYkdN
vyW5nqX6lzxD1MS0MnAnmk4mkiCZt1Uv7II56RoePO9TkTMmqYgO5/21calXm/yazFB/FqveZL8S
vM5fiHSbJrD/y2F2L4GTtlkaflrufRxE5v/YXPhslwBVvMgPfM5o3Rjfgjdam4d1G7m7ktAoWbK1
tWebat83PQa5I4kaae6ohCbWkiFbV7ADzBkfUqjxoSSErhhwYirTEwklYnqsQGbEra8AwEQonMwv
xnH3hy1hGhsLejRK35GQVM1iiBK+R3Sr0FIoZEhdILlDCJrnG3Qoi0g8ptp7PU2ras6R5A2QBKZ2
T2UlsrfvDDqRkLpMO8QlovXkVhY1VhVZG6wg2nU88rwgwswBlesp0KN+FJSdZB94lJElQvpkae48
DAEpksOx6GqG4dZDcnoPFeeG6HV3bi+o228MiNd4NsEn+I3VO/lTQy9J9GWwICBHEhI7mpowOYYV
eRNEIODB3jaQVYNlPiR165Oa9rhyblCiPstGiKygx7EpxGS2Zl/RiT9u395dBjg3xkn9uhueqP3S
xkf4QV/a2KlrfgOCUYaOf39fxq4b+Y7Sw0Za9gQpyxoL4AZHUEtDTOK6RhlfBHnllDpzH+Oq2o7w
bdnAoyArz1FKGguN3tPkh6xSL7F6PD9zTZFeP5SZaJHf9EnrE+iyagdUt7zv4FJTzPvuR3sFwVTV
tmsBKOxp0C3VNRygscdhZW8gJlXOxyRW9rohjxjYSJJPzD94oDE+/G4/WOUHSyQxExZ9FbTcwjp+
0rD+/XfzNMw+BdFyecjNsIOoEu4ogMl98sZh76Sa0UyOHIn+1cJl1eLvnfXiXKLVjBZSd2AxTgAM
tjZlzB/I0M+xe392XkbScBKURGVSS4FcfVxx6XPaW7jZSbodtOdsbkmpQioMi3PVCRAVOWuRZttu
np5JSEsHeCNvstxeyBChXybzLhAvmsahbxQM8ddAEB0+uL4maQV8b2GKQGyO9GSxv5tlfaoB3XAG
cxg+DepIWMukBNDJudpqpUXx1sVA+Z4tCuTTUGog18uaFEIVFLdSHMd8qPyrIzNX78xknvSLfnTS
1Jg+88xSEAopqcoqiii1uQDdbPjcwqYp0caNXX0Vmw5ousSxjAQ4jD9xfa3aDeBivi9mjx7zrbdr
QREYqFGT/KbX4Lhgtw+p5pDxAHPZvqA2MBM8ERcQydCXWQhs+XuP/jAgEpgU+TuP4i7jRovYa/gR
ASoCnN5oOcrfOz40bv8PGqFKOu2ymQoa/t1VLNw6BOrjtmli44VChEvf2Me+EU7wP6vcroxSoj4V
L73t5fYaBxEDxv1MdOeQApNicmsdbKAXOLKSIsd7Scbh0s2hivCa854UP6q+e+syV15/FKppi8SU
R32Jl2SszQI5QNa3XNRWTTosGhiTScXGjrBMz4pueoYiNFFQ9q8nc1w5QPdKOtE9xn+er0DFISd+
zy7YY0XFrQous9DNjJkeBtYTFrQcsDo81Gz3ohDYJ5F89RxuhvMmKp70eEhJTWJJ6tpS2K+1ezQW
jzchj81wnFKeVcYqmW6RXAoQrVqwQM6xnllUtUGHhAtyCAlCjrqWveH4GhiksctkgifqZbBJQ6NN
Gr5a0G/SiNopsv8gNjlXgwgrMbDzDt7vt6OqW3j7oRlcwepqC5Crnii/nES35VV6b2RulLBAYwlL
UG3dbPv97TCHB+9idMPoZAT6WvsdIzgVzKlYq+DRNqzTx3WHv8X86Af8+1FwhniuREKyGRb8wavT
gvzLsmGqG4NgAqj3vSsCthEo+psjglSW9Lc3i89O/dkou7kb/Ewp/brMOFNL2eObaSHsgkmtpEH/
rkcE+45CoVrIN5kZQpp3n6tJaogJ1xniXskkZkfn4kVnOtYSgt73h+NEWCby6rTWEzUXVbQSVpFR
cJO0KrcHSf9pkFljWoZdsSM2PGSkON15LdoXkmz8UWj66iZx5BGzLY4NbNrg8MfN/6paDiG62WQr
vZ3XdjjElRV92qWeQNZlJqGfIYqegS6GtZXSCB4vQwLnuryL3mpo1z5FlXBgT6nDrVGgC9zKfVCh
MBeCQO/tmx+WCPU/7X8q87e8SEn81d4sj2BpRoHpj/1MAjWO2BhDfQjH9vNNXp+TWnn56Qt4QWN7
FYzYaQpjKSaf/Qqn08OPAeoVYGW7vXU5o4spAYiA/a9Fd70eWCCrqMF0IUqYMy4TWOAsmRrlVAAT
0pBUfHL/P7N7QII9jlrTk6+lvzZ+QEUyMHrA5je1yD25SqNPg9WKckM5ALoZIESawJROKb0XUJ6J
xd6ZqcDsS8BWiXuFF9ywer1aGNqCZw4hViwOwvspJg4I7qb7pa331gldWsZ+sQvLLLbPi2viKuza
0EW1AyYcuxSE2X3Z2o1ISOI2BP+pGjKwvQZHAhJKNbLb5mSs1E4bBKTLSoXhrAB4putQVlu9Yt6k
c4ehwITBLeqaoSdE5biAZKA7YMJY6HAx1vzflSTIrXds6jC6weRDmC14rL//qyXMyuJM8VNGyYS+
XOId9F4BtQ4Zw08mXlJFuPcxXGGSBgPcVh44VHo9hQUrlV1JEZSWLhZJIghNqWF1Ex6i55OcPbQD
8m7QkcNWULHMijHytcr9ZQUHXPLwIX8lOwLNhUgO8je2Dkp+YqAhdMWAEPz5EuNcndrMWffwk/wM
QezE0SZiF4cCMuoSvivOSn8nR/NCMw33RqjtPUqg2MnprL2oe7GgTNhbpRMhiju4Ou8HhlUygqj9
1h0gV58K2UHrH7R0N20w5GBPtg2WnXIYS+30AfkFjCWRGPnAyJjArmpVK5ahY8L7CBNYkMHC6UAs
Vm737bvfX2WmtbsZcGG9H7dYD2eiJ7cHOsKp1uTHuiuxeXLaUKJQa4Fcvb0bZDMP0TLARy+5RsFt
IqaipS3fHX3FPAqJ1Kiz36d1At6/dbUcYoOsL0jDLKBchdzldLm4xgYOW2F7tFk7bO/R5g2MRjaN
G8YO3vZlwghA2PfJ4eBIcpPCLBKxKqZc8nb0VyvH/Lhf8YoO3MmsgPa1PA+m7Mv2hKKiZn2qTkWS
1LKGE2uKiP1aKH603C0nxHvDq25H4hFOYD1p3UpSSFpAuUs7OtxZ5S3eFdRrD3oxQl79k7WyoZVg
4a3InSywSRvohtefDjIEl3nhXognjs+73qFbMfypYM0buvPiCLXlUyLYVaQO/a1inF+rIk7FXkkn
Wo0aB+tbMBUO3VBd3VNPWKfpSxX8ta6V4GHqKm3TWD3HCT/xHdV2e3tFc63D6ASHKEM02JBF3VXg
YERh4eBBLEvRnfvuCWuu71geL0QGBIM2AHUnCrr3l1U5dpnOJhZovPvAWxcdSqxAJ2LZGeWebi2h
w52WvQ4Ha1LMt8YCT1InCoSW5xbQl0Css319icyrVdx2L445xXNYQkqKXtkZcaTnTIxea93+w+eP
yNBUxhkiw9nyd3S7ix5odCmMsBouemv9zgdFyjK09nH+9Pm3ZnhfvaSo/9MszWLZmJPJglvwiOVj
XNPo26YegWvyHpyBQ7l8C5iTqkzaEeoz8nxnclvZHk+IDQdkuDEU6taZ6fP/ifqOcpRgzYT4PS2O
YbC19lKqVMqaZSCXEsCQ+wGja2G+k1uPCEXKREW3O7NWYF4QTcFF6kc5PoVnkBjoK7cww1m1fijG
SWLID8OG40M+6GkjEfGLAhwC7cSvsUiuGyvziV0lBfcvgB9US7UngGIRkGfbX4Drw01qsvJVBe7p
j+GLL2f+P3TngUqiC6ffuC8ih0l+sizxg5ajTtiQ4wYskmYjzFKN++R2CUJAlIy39LFm05Mgd0lK
4YWEn2qRywgwCS8DuldjElLWCubN2Qo0yqOQLo9gY7h/+4rhmQ8DXctEqv5OIiTxuLCFgp86OHe9
TXl44Mht6rT5Cl94ifLYh4Mfxx0qScpbPRGjRM1UV6CQc2U3cB+aotN641k7oZysuWqOdyceeqJa
ebvHsuvaQoQEEkowqNf2ZLHZMfogFMnyToyccGtQLlYHqfF7Vs/WjBPJWTrFrulav8PfiUJeWLyK
Y8nECVHqiaSneQB3xkCsVMkIUixoQuaWMVaTKRYe6AHyh7zOKc9Gzk1tTjDpqLg4SipemBGNgYHq
R3VwtRnzGl0fLjRV5h9N2iylWRmu4N0GhjNFSUm0TpB8J9DxcBjtXuJmDNSyMj9ZkI7aKDl9oL3Z
6HR2KFGxm8fwZ+V7nvs7HP+vYE3nUluDgQbcIsgZoLRgrtFD4LaKgwjMDIN+N0ZjXK+FEQ0tWBhR
TolkMN5onsefxFPLTB89F7om/zXCRBZg3q3DwCYAMc+Va53+awAEj60UT5cL2b9drMoMWkCOWyT7
30hsWOCxS3Ri2O08nbKsbhZUnhKPCiPhnksO4OKRimfy3Wbd9CLDbA1ISeZEbolo0w3GDgs3SNk2
4gYhTCt66SaMBBMj1Y+UFJCKsL/f8ExMQIhL+gPOZJii+e/uXlqBuuPtuPc98yzGY21RBJF3WejJ
F+U9qoxPugbjMiAmxz14FbAW70mNOIZvm4uN992fnzFmwuOftJkS2my2vdRaI3lS6LTzK5ntQlNu
Q62w9Tw6/0yuRxnui1/yx/q9Hwc/N5uVTu3nSjVEh73z6oHgDQG54TgrIwS+f4MLZpjkdUEOxnuA
f985iPXeaT8EOq3+MB7gqDVl0UMkcmI5lXX3GQ3+V0H30PE/v9jAzm2Bzm4TdzHPdTDXn6z1MzyZ
8Ix2gir3Mg/7/+W8yuiA80tN9nglSKPN70YC2FfeKSJm7jNb8aKbvv/OEuPd0KHqxXUHKEDfiPAX
vHYISVE2hTEtMikERorq5aGT791GnRO37t42ehy6kQblrEmatgL0xKx5jfsoMLp0G54k2b3eyGQ9
pqIoDX1k7Ynmr/V6ryBOz2U4I11D5Fbs1qnnWVtDUySioDI5qeGCOo6iopGIMx7tP7VQQcXt7MKk
x79Kc27ycTcnjKrw2vLehtG15+394w1A8HNw8ixviLW+bdwuPaS3C1g2Twd+TXEkEbz6ktHbUYjV
9wC01SoKDI0dnlnoeGLPveHpoY6EaaV97M4mMPhaOi1QX5AuEkuU8rmG7fyHAqZUWSGPWa3bRn8h
dkC9yiLNbnPnIKB6McwwbYELyLpwVHXvihTS9S+VvGAZwP0trvxdQ3OuR+iCpwi80zMScuMu98ZS
4QOzhrYIzbQPXIxI9YU7DvQR7tMQBxegiF4uAGV7Nm+BB+hMcieZNDT9b+mo+/RNlbr9qTK7P6fZ
H0ljRlhmU1M0cCmb6bqkuyuQ9s+XCrsLtGIj9v1kZTDfK2TjkbbOOUVZrHAlWY3hrXkQdOTH1hHJ
6LqpZ9LNZdvmT2DAIe74/mJCQ1vTBiNMBQNoleYeJrOHCtaKy3kNLKDhdDUPasXlJofW4veAJnH9
nS0GonS3g4lp1SFz4zsX4sBk690TDk2GurECyFmV2EUny2Gb0bEweqCW/X5ftEr7aFsiFSnULl+c
TS0SDmbYPK08cvpmBM7ArSs8tJJhBwsA+vyysQ1bqmgUoqz+SHipQLLXlU4sjCAGtEBgyUb0YDQ0
QsqUL3B5Jf8DtVs0q4qyLUuVrrSKcgYOXkOTt4tbpaFiCHyTmVpr/9Let2cOsKAIvu1jWecTbU8l
u9KbHQ+sEWf2dnsZxKJuTcNZ6nK3O/TgwYykrehdfZamVjaTpkiDif6mF8I2bXID2W8bCFTQdw7u
LmAT7a98ocSqJh14sat0NS5SdX0B9QD5LwBmoKWuxg7Yh/nYj82nhXXmHNtemkLgJRJTBzjXYjD/
rJYjm/oO7dEZuwAzPhoFh8D7I4UKeWLonFkmz9aAZg+kXnEU2rRBxlYeyI934zVLWfVBGpL9yaER
tkMTlbieFlVOmgO50nFwUqNXmtaRSweBkGe30CfmLzkBguFtl/OTH8KAB3uA1JouPGnugOzLEktd
UBtQLnqdjG0XgKKNa9AJfQ1Ke54ktlCEhqCd3XWCnelU04HIvCKI2foKc0EPdMGBq5p3BekuFvhR
c6eYyjdFBiN3/POIFJJA8cwYoMM/AYstkm2epyPOC+YF+MD/XNI74Idw0uhNN1XhlumYUVKkVcYc
IitZAvxLqs4mQUUW1aOr6uOhzG3ZtRHibDS7wfx78lUQImM+cxA/m9y2J/bQ2qD9znSYsmBTMNWc
njIK7JOuI6fCdoINwjE97szDMzV0XZGhwziXjHM6EXcv99wwVh1Zj4igkQa5wbpCfoszA0l8tHF8
0QnqlhqXACN7tiqIOMUe3eiP566Npm69qaLOSwqO9LwzSVE760ZfX+67wSOg+aKIa1ZXMR8mn3L4
Zy2xnE3CKKrtjBkzQjmrHY7TexA8hdcg0tJku8BwxHTNE2geAsJ+X/KfhJ6NvEqB5Xdp19uGhAmF
jEmqX7uhk6kKMJtF9jiMrpMovA7oekwKZ1T1z5fCUL4Q1r0tDssIvNDrVy/kyGEjmQj8gjCDKCqD
aXa+vGgxQN4XXDFzxHzt1Uk+niWmSB1T+GfX+hmsF1QOSCupJALO6pIlJ1Pf5z4F8aucDfIyLkSu
u255O6DsAfJjFAbRTznvLIPrEBnYrqQ3jGpHyozDJookzxsTx4QtrMTOxDXo1hiizJ+jN06NFKSd
oGiKV+pHtKxBVACmMYOfGXFjQ5YkW/e09E9FhcfLn4qhwabn3J17AR5VtpEKaJ1Vn+9vzn3xdDo5
+68aI6TfzQPKMR7FJ1EOK0kbd1rHjjpIPtwhIDy5pWjawCppZyaNvbCVxB25bJhGUo0UO+fO3QHy
hL0f5RK/sDIv3TafQ9btBnVlTcw2ApyOquV/4Qz9EeTIujQkKuaZtAQlnvfh7ZutAvKwHO6veUh2
QGwv8+ddfeoGSZGfXNqK5Xx0yMVE6kwU+upsNrGYLypVzGrgRjeQcWA0qPSYzQ9fzan5kafHbQ4p
EoBt5p1I/1MVjF/MAPIhC5Rw8DtObQpTdkycITTWbJNbW2uYoHrBhi0T/1g4zrPQGusTuOQJbeGX
1C2fdtoUCW8yvB+xZpZcignIe08VoE2e9CNRunBDDYBERJL0xsz9lwmUdis2W+bLToPFXA7v3R2y
M/Vv6iqOz0r2L2vlwfOv6JIRBMBS3k7E/CTA2JqxNe5wql+1LH310tEHmtjcUa7Z95CTXD2ctVoc
EtZOxjM/Ia+75nw5m96b3SHsE+CYotJLVn/SEXoEJ4j4zezlT55JmKpPPcYd7D7ozN1Bt4F+Q6YI
KLYyo3b6ql4royRjTgposdPBPKP0UrtGBlwq5IUXfUYu5q4E9zINIUgR7uNUYKuNH+lOOXvPoXuT
M41d+m+EMDRFmWysUnpeqR9ZKSPpyXRtqf2offdJQqviT3DnSCLDCSndbFTe3dPc2IV/gf+DLx50
FVfMfTx4H+Lz8nych9TXU4sZcgEb7T83KWYrTglCjTlYkdXZv8s7Se2vMFLjyJkdqqBeuiiGpmw+
X+omRaubsC+EGO5oClHMnkAQkSq8f0ODDDYy2BEJBTo2BGy0Y7NrSTLjicYgo6DzZGU/8FBw8JRT
gIPVo1r1XR3i/nS5LH2C3fXgpYMRoBLz6HnUpWDPkHKJs9qX/sdR1+GU3AyLyaTVyN726clkxjUh
QakMNQLfJY/HJnPPjdoY0dWY6kV/83aEEnhpuJLELZQiqO2HagXLSzSdaaQ2f/B2GMffQPqwrbM4
dluLLgQlqbFV2siaCdrvjtC+PwKi/jMPhdijxYPSmT1BFL5vqy1uBS2jnhW/H09YRXrXB6/XT+QF
5bBIkdve9nvlGzo6ato+tK4kpn0O6LHAR5q3rz6zhameJsuEyEoj4Jj1SV0JZkljTgvshZinQLud
bEcrJxZLPVFeqmHA34AIIH0uJ1B/8UiCPoqIIJ33OtzaTavgQL2P6zyrQmWZQk3i02Rd9BNkk3hn
S57Uw8t4kooelJO0Ol81fgmqjrgRRVbErgqTWRtjQWSrZ5EnyB+gYRFVHJ9w3/yrcZWGo/oozzLc
1LQ0PHlHGI7jI1FdnofpStN5c00Yxu6CnEKFn5jwFroXY72DRfDfz2PEiLN6NMTLGAhM5NV5/fCm
hiOVPAhbWA+YPyUI+iLWzAstohjgnxKAIkf0rUMR5shooUmDVmBqR942VDx6osDLYze86rSFwAG2
djcAB+KYdyrGIr/KzeJ8oK38BQ1IRCP/ck8RkFjc91TQNvvVq6124PVTMGn4ga/4rTyMJhw+kVLH
Nkf/I5FcOAL+synJyzpeP8W1Rg3P8sKdsf755vvX6rR3QKg6RjSYWhDN90Wc7g2pg9zfpV1AZIgr
YBA25zNymj+tvL2YKjjvf28dG/HQDhWpxol5W/mds3I/WFx4gi/TLa8PWfEvSBSXnpFDF60j+2h2
fyWtvMb8RTPPrO/etEba3R/vRCMnApNuDC3Q8T6HVDlm5gP1jh8Jh+lIx5OMc3cz7NYp/ss9JCz7
ztvbstTa80Kr4ayljcefll14yJZurQTfgTyR6O14C9cDpeW7C0vc50bqJF3c9+Wk5anqjkgnSAS+
bNgJZ2Znpf+iPPwNeeTnW8Thvtr8JwGIgmpky24pZKm4xX7LFNjHaI2DioAivKLQWnQwVV9rlEyu
zRBaxSndoklEZ9AcRd+z+YfgGQ0sRmVgqi3rOYO+c2G6VuuQqk5IUfOTmIa1IDtuHG3F8Kvyih7E
F5UdS2nWJ87Syjl3+JdUfYsIRaiZCLFmeGzNWrH21ksACHdkWwRZE0/Y9x5rDqRQDZ6AxVtIpkhN
bLR29+aA8thstbnGyKEm2tchMhXylwJr1DxzkjhqG7h1ZTbtenhd0r6unZIsgboOdpGs7IpiT6si
JTfvhtXyvHx4CZT0sghmRxteRKv0GGl32bYGG4rX1gbmhfcxAtSJmmPPi4qjWOsapXjLjrEhuSeW
nXRDZHJ0LLvkKjCQDQOV/FY+I1YbPfallzVhsnL7Obn/m0/N/gIFUylPIvBipnGzERzMYTc5/hGy
AgcoKL82u7Ao3VbPzLJfAwDo8igUDN/Sjc5GsF3Dcbuet7k+F0kKSyAqq/8B++9MyyFcIG4NtADI
7vYiWRUxkVSIDJaTjcsLM8ncFULDVBleaFadDsTNx8T3zNcBTG5HGYJuSqpk0wU1k6yYT4Ja0PU+
6HOqqbiE4ZBIrbfqZMJpbPysvrWIGm/lZl4foV2ggh5oDxOPZWfwtG4VP1ukDz8E5XPcSox2D3AT
w8Nh4kdIJT/qVhEAjT15Nfvv2skWcEBWTHCTMI7x4dHmfc0CI0y7u/kBWm5P3e2j1rrj+FLr4I3X
laSXxKE9SjJGwOt9xgRo3XdE6Ln2S9c/aBjKnjfJh5Fe0QryE+tNoGxe+CSLVjqby3cEIiguS2dw
L9qBvFRfLXxqWLyMYCqcGg5Ozt954vcEiFqibSHJV3EAUAwanDt5sMShkpsr+fGtRrHih0Tbquct
vsa+/5I6Y8bq3Lh2IzycATgYtFMKf4KNKNcPSbRj/Eu6FhbbRC6urXthRC5v/sBJKT9wfvLRmV2H
K1PZpW1zejL5wEZYG3S059wCQAX+O7CcFa2Y71T5phgrSJjTj0bhvY+MoUONPgNCO/5OQuTyjy24
j4F8lb7zf2KqBCQG12RvkSUawpvqrZGIS2iK7Uw3NE/kCA4PyHVdjfZIAQdpN1sn8vQWHcTAohiC
2XR+FRdZuPakwYBcv7lFR9yvc2FUxbVpVaXXjHMNdSdkVtTLIzEni2+fKEo6muvAHB/w5BGD3X87
VQVYJAsGjUePXHl4B0HDWcjBYVtuycS2Y7shdrjMVbZYPohUPcl6QafdTaHQWJb41VVUZqN/U/F+
GpsMeFId332vCez5znyCIvRDNm7RHAwE0wG5+EcCNzETlWoQrUHBaw0xUjbTB4NTnwkt+rkTWC3p
ThCFhUq+CVzMMYJxLWvf9G1MYiEw0UhPHWj0PLj7ojndZU7II/9TXJdd6fpxfgCAR/FzN4EmkqW3
BUN4j8roonD3Ij7a7iMIERXXXVdBCcBRQd8O1gu2hHjSgs8vPKnQSmWZp7aBRmfFyLgs2FaA3I5f
1C7ZF7e/86GJKBO8NsaWvbki4EXoFwIuKFCQqIBfB7oib5JCbNy1JaughYpXSunx+0b8JaKon7oe
LLqpNjSpuR+1zIGcWoKWHYlJBLzXHU8za0XFdKQtJtHwFUTimH6MsM30Vhyr/wZqjonIS1PSfTwp
goEMEq1sP4Z8QVgSiKSrC8uqDQg2Kkn3r0kPsJZ8qrSQyM1E1nBYvoyQbWlmIpYM9CzhWsfe6bX7
6lC3R/F0mhDq7oGxqlg4iE0anFAYLrI/656glYSDuEnmfFLoo9Mw/jj4ZX5G+a7rQ8mrQnFQ3XWT
cgR5gsUyMdlm+bH/PGMuy1Z70VE/TFTs5AwNKwJKySz9fB2e1mytmPO5mYeH/8eAB7gpAd7Two/b
o893KOVD4u+LWryMpVYZ5kvcTIUPd1mYQd85FLTjBz8Dc2FSJpUV4F5BRFrtCInjZHityshIK5so
Iq0F9eO7jQ1l/r6sHPfUpyooNSVbDAHv7MaiESV3CA0EIwEPZCsfD+4v0N4Hdzkrlb6oxWR+R5XK
NfYHZuH6913Etv1DMGt7s9ZTso5rMT70eHfzVJ+BkHihbpcCVi3QGu1Gem4h3hRstnRwzCpGYgj3
S5ZxkLtpHm+P/viWuW/cD+WEdHQqgJIm7Zjr/WAkwvQeHMrRoAXdvX1Mef75fUQlCkL08pq+q9Us
3HZIBM39VRVd7DcCqXGKc+O0nPszk9yMxwq6VqRDKi4Yt74uVW2gKNmUg82l4QqSgmiWb9qpNjek
Pslolj1iTc6YrY5LZAoZgZ5siPuXNqOQu+wVMwnKOHzj8g3PDihYfPRD4M7RVaMDKNHPvrYkuuoN
9TFIOo4yWWDs/njJ8ZkDFhaCRxf2b8DIQk9r1ArTNgNDISjT1IWY200IK+9KtchjiQzgX+9SojYr
lPj0Y9Yp89OUxl4QCbEb520I9G1nQ7i2vZ9DzhmMtY6VyGHnBEb32AGn8qTjcoK3Lg6kdjxwiAUd
F69QbWZJAb/v1a80cBvwb2AcrXuWdTXMBSqn3ANpOxyWlbKOuBpL7ixEh0s+1wBVGLhsGZrVUhjD
b3M1z0MWvtvCvpiNG7pHL+8nNf3JN1C56DxtcB5PEU0km0U3hDJG7NCcOEcM8HImLe8sX9HwRhfN
+YduPkGqO/409yFTn94ZcWEtB/7rIhWlsGUA7QmEZnYlgpejI1G2VYNX8MuY0z204x030OePs4xj
6jNKTChfwZUaRS2WLcHPUgrXuWEG5hoD0BP3ELyjSW/2FeCEfbiKXVZbK9ZeHME30ZQ5VGamsePS
asqfIFRJkzPl1TOwlvlKlxsoZQOGWu7fZ/4aLKhqxx3B+5V+Fkf1SQJvB9MlY/lssjbsYAi+pLNO
xlLX+lBTjy2x7fdoiWEyXcLJ3FVu8oINCb6X52e2FYmrUxVPL/wHlISXrFTHqL05gleXCq7gnSST
3cYcJjFDCSOG5P/SaKL7Il36U92d3+iYLSEQfCp03bYYdYz0LywpSJnf3nBR81WkWK+H9iAya8xc
OIzvxhhQOcGqifc7Fbljpj/WTu7wTdPd976QUlqeOemImIXBJYOSp+itR2TT16RRccKWIShO1FZ0
3viD+ErVLcHyisasrC1ebtjWo1v43v8paIMpmTGPbQEEYe+TXO2KTEus/zqr6toi2i/2U4vQqPVy
EnRxxIyoBJO70hJBjQOmj4M3KsE8jJybVUTGRdWtbULKxQZOtw0vbUjFa6RyeO+HgyAhHz/ZeCIx
oKDroUwewCKBGgL7RVtKneKCaWgdN10DjB40BJLcmmOavuxV7UcixI2bMtxkcbKxSE2NDnvnck75
uCdEjTmnUeyjT468KjdiqUhZVtdwwBVVMY2opJ+fqZu18OJVMvU+GJhdufffa+TTrZQMNK9MNnKz
/XA7AJa6khIXr4Kw3i/lzAjSWhr2mvf3Kx0tAnDqiJp51zdyJ9cPjqH8LaDPr1MZHq45HCtfar98
SqBvvB76uvgutXaNua5sooETm5qU+nQp7yv7kJgyTdZxdYGII8ouE+5ZEHhgyXYyneiD9Kgn02mh
xM1OYckFfm242H7rr6Ge7ufuDP/I1Taj0c45IIolx/Wss6aO2Nf9GY7jQsj3B8J3abbDiLCvcqEI
LZcYRE4ylpezdwQ5hWAon/Rz7qJzHBQAM4msuX436dzRuAcnhK8eSzBlrBUYkm7h7ckb/ljRDozl
Buu+mcxnJW8LqJlVOwkWxLuPp3dE7+e+PqjDl/6Vd+XTz5XEu3EPD6qpVQj7KNh2yYE+auQzpe0M
CjeCaxw9xtwTO3HtCGgDvZiVJmfnZadpYVC2eheAxtsy8246PyzBIDdA0uYkV8W8QQXQ8BxHIzNb
yDz31ku1AqUxj6owlkIt/MTzhwDrWpcnQvP8aaKrVZyDeQTYn9D0VFfuQea5h7J6bica+DXaw9UL
X+aHPn1fH223Tp2x/jFUWt7OlMztkXVXjVNfF7j73x+/2z8UYYoU8ijj2yzwC2OjK4RYHGJTz706
HOflASMIMaG7I8pHQPCdWs8ItTG/rVWP9vJiA6KmcZ7QX3rSVMrN0GllbfCShQAYUPf/DH09DBBy
YanEg8O0Imt2Jro5cd6PbomanpM0ruKZRvoR9HM6K41X5U+JkQG3ROI+OnC4cZc63PVCKxNZwPGW
Qtnk/y83WafiC/aE0AriTLAOlUYDmL+OmpOLMp5dH1auzRmNpN1Ij9Nhxqt2Wd4XcunPaGdVFYz9
boDBgYS44VS18uDeOU5B8iMXU0O3iXrNyauO6yITY8zUgf/t613IRf2KXusqvwHyjRs5ebSaKhS4
Ga4HLgydkmG+nVaCtmyycW779MIHuz/HPqrJ/kAbIWt6ZgpUOosHsOx9Ni0pxukw0oYZ2zbXNm9T
qN18IsDeHySay9Ap7q8JIe30E0nqVft/N85W68Fcgl4TDZpXsxVDU6n5tgDZta2xJIDD8WVPsWMq
/S0uZj1iYVvuk7G35oupOMN6e8N1K9VRuucfjZMVh5Ojf0ONdT1OkBZGXlbzlHFN7ZNTlSQeUvCt
UiGGDJk0qgBBliwzkRMBnP1L+EYRpIfPGRN+4XoF65o2liFfCEz5Y3Mq1kfcBqXrt0Ti2O3fzXgG
3XKMI/eHaopHJCa2IHPfnHYPrYUR5lW/oJyua98JqNKZTfZuq+2ARaO9AuOCqtyOhnOQNtDmeiWr
fQbgxgbYfL4AdcgmGYRK9uQmWgBXyZdZT+UL67SIRSEEQ3zhKtP3YxRMwqa+XjBJy+cqul1moyvX
da6D6mjuoxVZyl+2gOEdJ/lwODLSyryBMovK0XMIVMKev93u9kgiqWGc/mo7EAS05BH2XAPHti/A
l2tYmcp9XDfXkT3JBxwfEWg2pBNmNNVbMK4cdJk1k3ZzdkUKJOOsFUtgUsFPT02vA2V2KV70Tbrv
v7hD4EuWMgj8eAnHHLmgFTAAYlX2oYlm9PHrYAJqtdSJrZ6taTcgkM8tEn/FUbk5e8nqgtKR/DlE
ulgXEihaN/T37oA/lbkegvDDq2qlYasdquokdxOdPFnjjymqMGyMIYy5oH1EVoEe/LPvNylosc9a
KibljCJQku8sjw80EQk/k6ziFRU4LSfDku8IEyWZR28uZN6ToYry947uBIsDFaz/SOBemFMuQojR
JgndLoNI/gHlFtZer60LQIbtHtz0GLgdO5OZVdCT16ujKzI5ZnNhHIJ3Qlw3Hip9bpLvBIcmu+3n
8g8t7819OKJpYLXgvQsBj3sttT/aPvBYpj7yrDLoPQ1rJ/iGyOKKzpI5DN9g0BnADf609eVPih//
u+UXdNxYtrZAxcqUJv4EfIcihzlYEe3HoBm+U0j7HErvTHMfZOcMJqUTg0kgtU87+Vaif8PNYfjM
cJiz57vIY4OtZZUCIhXhmDXqhsHihobE4xqAw96D7Gm6LktImBQZ060NJCBacgKsX4s2g1kbB6yk
06yo9X6dQKBUC5n4BXUoCF7CKS4+S7s9p6jetaUcsm8MDZfbGVMBBxOZ3A4ECzoO/PaT0wdRxsb3
t19CUfRPNFpjx6UODJ2RZ2Qf6odbZTkq7n+sxvwXfebpKpmhYsywFPgihAWS7491RGgcXCFwERy1
WJiN9OPXA+qIa9Scbcld1zE3wGYtx5gy05H8sChxjgnX5IqJokmlxOYJ8gxyqpQ1KhtYeCpar4s2
SL15ObWSfoQZvYfNT9C4ky/XcKIu9+8Zg38QPpya4cm/duXUoTafl1xDN782nV/fS9ghrCKHpbtD
RNx8Hhz8WxV8EZn6p18TxH2ablbcu45ahVSinXP0Ejc6xvskPQ/bFv2gQ/EeAyheIMEv+pH5TZnB
8lgxlX3vm8pK9FWCRja6pc+ayCMMpLsbeBM86FLFA4FkP34loH7lVuDD7RLQuHbSqsXHaV/BAWUw
rTJ9zYbCMYxHta+HR0J0yrVCKxjs5zUKJ9P3SVpqbEP2rxAa9JAvflJg6UoUKwMEEZWjXU0Sa+E2
B/lKFkBO4Qszrxvm4kjVf1wUvkMUhE++uN3xIduyb0PTwdavXRXESfSfxWvSP0TlBMb5Sf/Y9rdI
HG5OSkXqumheLP96ZKUCebA2vIELVFgkwkY3gOYt0B5raznJCFwa0IQCuT/XtCRVqL5TY5q6/MEy
YcTrDVquyPtpgNc+EIf/LWU3e2EBXFhOI1FWmyT7iRZ4SBaud9OZ0vLB6tvYHdmhLUSrkd8mqTLk
J5qQqtMn8jCy3UlWtNmjPP4Qt1E1oEs2Cxwnt+LWaNuxLpeotbvXAkMT8wwZhTHZZqP8ankqqt62
Wgzle/gS3+U4/ZpKe00942/yBWaxXwiaCVPp3rn4xLk95re0v6yDrUdbfL3w43/lxwzcoJ91BVNw
kgH8iySVBqwD1633xHSfpGBkHzjFhY9t3EiIi8kK0rG1Li6ZmJQqZTnLc+pJvSdVhbF9XChHo2R5
2md0QnxuvlUwjq2XZPU5f97YrjYANTS1V5TTexE/kfX+Y0gCOiVbvILUObu8raOl+w5jmushdBUs
H7chycMLfj4mqGHjQt3YRJezgWed0G4MIKpO9UA9b8Irv8MSyUPBWVE0N/RKtckNwfSZka+mfcZv
MeAsdgYE/S52SoqCHBbpYkbn/Mn6mxwE9pWIVZXxb5/e9VoiZVp2VBydIhQuzAg7ai7E0X8Zw7Kn
k8kUi7UPAz4GyuyqMKi3OX+tDk+VQMN50D9uyh+YW7UoRH568f/ixc0rpejT9JUKw7bLpKZ9PMtQ
3ByHyzzJddY0C4E6OTUhcaRp1U7UIjKBJTcCGAESg/nbUqUHrzCL9dNRjXbZqAilGWpcXqC+2XKg
da9sqo6cNirIaTuLDDbqs3nL64FR1PugLf2Fe/ntGUmPdm8THtEhcxqOQCVnCU+GuncmbAn0FYXh
MSnX9dOIsveYMi2Y4LUjF7hUrJ4OT/U3TdgV+rbJwQgNCk+er55PHaOI3ewGje6JpJ6vSb8PgkwH
RraZZEV2c1h+PzuKU5kl7XQMwOy8OYFPNQF5Zl1Wz5Hvl/noceobeUMcPlKV3d10dc4ZesemKvHp
B/nI14A3Aqne6z5jPWP3okhY3N8xHhgAOh+S2o3AAwoV4c8XuKzc+DzloDIkKN0z1alPBk9Z+nQH
kY6J7gXG+arlBaQOswAz06Nby92F+oLeCtYroArB6j0/STfZLwKNhitI1mwPEmErzh/h9bwPa7wo
YXlOxYav1/lwe9z5BSQ+fh59nNH7HmqdDgT8Ig17+OXNYupc5WcDzlZNldGqjgrZmu58NP/92V+e
ac925oDOtxL0Q0xrj7+6JMAB/oNSv9SJ6dxmuV7aAN5hCvIE/aZU3UvRX8RRTD1TuEqhrcg1+fwg
KajerPXfq7+Id4WpdriSN/TH0AUb1nqO4aEWVs/W6h+Er7eDKYJqC44pIhuLbA6yURRABUBYKDyo
tWmWodYZBR6lZpCfbVA/j/lNFNx4UbjjhRO2oSHrJBpJmE/wFGesoXIV4F40oVwSJmls6vT7Ofyu
Uf12PjueeYMB/SrDScQyeLm8qf9LW20HVaFG03cLGRT9v97c5HR0B6/4fDMBP2RwCP6lTzxUwCJ5
SFggFvQ9n5GemlbT7eMHLd2nz/wm/dYZWVmUi4Ff/1CXgMaIqSSFm5Zz/CHT2t6r6HxtjhryBdw3
bXSDVMlEd1VPNwmbOuUb2OYUNHy0Nan6DI5WhpS1qxEOjfMjMISCld4J8EQEgkbZEUXuj0/dE/69
jvaCzFm+LEVK0A4MaTJ56dA3FbnpZg0v6UPulHcHjEdY7Z3mX35n+VeYdYcOpLCxIbBBakdn/IJo
jGivlTlf518HVpJB88T1igCmtB3dREVckdmdBTJ5+dxjETNw0elbt9hnxcS0qAen8TjK78orxE6T
qS22ZwoDL9qY4t1ovMey5BhFuVuBqNTzEOPAVbDITRubt66zr5sFcxa8JrssGxQ8I6cSWRnJv1Rr
a4mOcZOWoZsrEu2OzU9NM+NQcSvFkVprZ8MZpR5tjbZ0BsVxvW1aYwk6HWoESG1AL/GWU69fOKlY
JISdBDD0FIGeFb12Qq/7OEchFPJUeiDbQY6BpjJJduQHvjwJgOrEsWymrCKE9+s38e1FuV8nlgU1
6R86EiYH3qw1Tm9E+r/oPBkbyNrxkmdx6khwiqWOytMex8qeZHnh4m6D9X2HINUfrBamj/AQvCsD
IU3tgWjrF6kpc7Yw+L0bOGcNhrwgCxVE16FE2XqnMOBctLr7lKMG3uQ2K1llHnxMSGomxscCU+Dn
lzxUDu/R4RyvIVSqNsm5hAOwG2NuyTf8MQR+2CTy1SsWOa6suBuIfp5jlFFLOlnOa6M8jb+EzMYu
/qaqKagneBebzptLFA3ooiHGsGu8T9eIzJZ4zPW73ccypTKkW1HXRsEpxli9aS3mUY2j/ArEV7Wc
8Yjpb4FvPEXTOuUbEToK6pk0ihdXKwbHhr807OB7b8/VJefI1oui9z4prAKPIJcRYCAn1cSX/VMj
NTjpfsgYm9chPdxFOPZ4/ERW0c/qKly+/Xc08JsarF2eD2UxUoqS/TyuFqotlmHEXlw5VusADbfI
ZJysjYMS/1+3JuamaxaHyqCIyRgV8VFn4QnfEep1QjmcFv0HJPMfbb6xp/uh7CSq6DWQCfm54eng
d0zgwz8bR+qKEkSuc+TqDUN6sv4Y5FUge/FWLjGJVrRV7oEerFKwU9xFaam/D6+DlWffB72KwO/D
/YrWD+PQjaiXEz4wTooE/7YSQl5o+ceUUlDbRUeYU2YxFJrk5pbVCZGHloe0ocGu7exglu011Kj0
6WwxRo96iQ4oPvGuuJlHIY0iqDjednxKqRswmksmaUKSNwx3ajjT0F7IanNIhORonRKv9GaH5+jH
157MKiIU+MQyRkOH0zCogL3x7Xos2mC/IUAEbKfV9QDHEzzcFFuQqxXyOSVs/xijmip3zu2BYogZ
LW2HlyWOiEwnJlI3cnFcBi9szlVb8sIJhEhpiKHrBbpaqOS1Y2KkuiaVyfjiRViOSC+94c+x4GFk
xdVdUl0/NHWubtYeuSLWOxLHaJDffJC1gFqTHuwaEkAEH+hvLefGJ0mNGhG0ChfjfO9cLv77Jz0g
6Ar2iEcou4hYECHIaavhtsDzsoMzt5g20G5GYcvLhXmxopjQitbjKFxyCh+k7Tm5O4EQyNevNivu
pIZI5i0O9U4AsEb6q2QyrBYZiAoQphVjTfvKpGbCxF76HqpzOFUBkAI3jA4RTnX2VLIFb06Z1L/r
bbazkM5ohtP0zUoq4w4dE7Q6nfkvUnDYA8kFn/rE5B8a5t4hnXuYc5+5xFGeR5Q7Jm/NO8n6ApOB
bxdsQTR9xud97KHvBvVuj5TOoaOCmmTczIK8/T+OKWDQJf8e4sZlhNOVnYFiDOUuHIbuyuqF+jCF
WYBc/J3RzLQG6Nb/99Lt5jvtC2zc2wzQidR7Px0D4xy7fcxnJf958e7kq6RjCnlDAtKSsq6Z5R6N
e3WfFlg9gQWK/0PlLUtIBB1NJZ3nxOJFGNddfLynwjEGlfPj/GDZYGAJBINt15V96t0zCpOUK+dl
dtrTaN4X2WrY1Jj36LCXLwbyims45VEUt2Ik6jINEmXlTDDwF+Zg08cqoxgGSBneprdx9/xJhbFA
y3lLrEcOKXAjCK+s5chbksVI2VgF6qN5ZyPp/+/qYmCDu7lnqGFXb4xCLBT4/RW2Ds/k7o/bKWV3
eD4e3Xb4JzjqmkMtFwrHjpLoo67UCG5h2FyA2S7xywx8whLw+hxkrJ73mPZ1x+yeF8rPvb9wnQNl
Qui5T1Ym4p7q6bq/h7BwaNmAkMd+KfuPuVc4kvGqk6wUSltYTIbgbzkfPovbaUrlMBxjZmKy04Jm
O424msxK5g+NZPv/kPicixQnFgwzSGtLj8S2s8nRJGdGeMEnQOJDlpT2L9dQaFdd0llkQFL2VihL
7WDs9RnKvyhNsyWPQGmWUb2oME8Pj5VbMVuefOyNM0OhXDWIzj90b00AHltErpocMBmtieV7WwEr
CJIUTuN158SWDQxxI35aPcsHIt33uiB7KRAfNEBsoHNraxYI4VMEj49Kjo1JRs+4w6CYkux/Eugs
o9jgd37sDeI61D13OYlQmWJQYJkUBmgGZ4Twrzr78U44zk5V3BzhHCDf+J97jhFRxc6A08fwgEuV
dzXq92Tfe4wv30xi64LoT4MdpbLmE17jpoagq2AVTz4NzbbI3q8qM2YJlK8zdIYusb6FhkO5X31A
kAt+56N5r9ZXjQIfoHHj69BFMGtvZ6j+rdRu1dSwedHs6G3+NPYmcG6SA/WnMqyfjxYoEy5w9W+C
tE7nwSmIpUHL1nsjKQrSDIzdGUF7HO1Uz5SnM4Xr4Wcm7nVwRHD0e5DG/Ha5iPmRfg80dYPyV32h
hkE+YFJA/1IpqcjeysqUFL+E13xZ1C4Vh5UmHAWAi58CYAfrzDoVEpA5bem/T9e6boxH3ZUHInMk
CWy9kN0bpfDR90BMgUTRVh4USjeP4eLNVoIO7YJ1+TYlsm1FQqrrTSSMg3FaRpvypdq31YcioHey
d/p0stmS1R/X1XUvBrdA5NRNhujd41hAlfu+zyGi44LV/AQrh15KG10/R2Rax4ktBThtnbPGwq8E
PjuJYrfgYt42RVpzy4eALKhi2vl17zbu8yMyddxuQa9S3Z5j2jd4/trnH5jJSGLvhBjkLk7YxO/8
O9KwkbTsKGUQEgjaMahE0rcrlWqYrs5ux1tEPj5oVba9It6BtOnwd84H7fktcXrpLfrwivok3Utn
HoTDEBUAkrrU6uHlRMiICbPKclkoA3TZ0ZAvp5c8vcxIgGFgcLOJKx+y4ah8VDTa9HYLhkkMVhHy
GFxWF6DXG6OoblwvsOEfBuKwB31qMwwITu3iCeNaJTn6d8N4a3mxUL0AnXYOCE3yXvd/M/RL7INS
ptFpxxvqHWgytCCwQUBarDMlbSlg2aIgF8SyEzzF8QkFq3i5D6EjEJL2lMrx7887EmjaMj3XRwz8
4x5xJotyT8kGfh0xFrbz83QHcFimAmF+4mzqqgbdX+16XYl4jB21sjPp/P5Dbnthqt2oxBc3fdJs
JxR0BX0DdpBchKYjcDHKymDDUqF+E0+ENgHqwqrSFY8z/FvuTRN2Ax6HzaI9ts9vjgZ4+LVUn6PV
0UfbHS6HDuR9KqaOKTu+22KwkiUCLz24IuVFoujljibNxl7GSYJCtFTgKpg3UwMfV6JhBPY2bfyb
zGSAEl23KG7i2BwoGtg0sO47fk1hgh7dlitdlY8DokTp5dNO/4N1BJouANGyI5nxyfAc9Ld4rBCi
HeKwoX/8bIqHDBW/VJLBkMYM03iJiLy87b7YSX34nhY9hwk5MR1GmG64HVo5kxqy7QIIHRQCQALW
dZ4cHav61xiD5enVNvMe3g8X4VNs+0cFU5pjGR9V8kjyvUfF8eoaaBOVw1BkgzsnvltKPovQveSb
jQMe0Z5g47K+o+3GPzpsGJa/0ZxY5VSB5Zao5iigOPUpho0k9UzcXt0aP8a0LJGix2OjmZLbqL+t
W4/9zbfTQ+5sh4sA3x9914smfz0UXpUienXfl0dCixUoCU5C2YVybdP9wsul+Zofi1b1bd3LKAYE
8WVJFSdcx/v6IyPYfrYh/hiNXI8N4CuYTdtRfFtkRaMUrqkKQJveIYLDG5iCQ/mfZCNB+biD19w8
9nVDxPn7/MfDfG/5i5W6+P0qqxqf/p5UymyiRDyaVk0Mxw9ToX33bnxE2um+9S6Xh53OIdb9bPmT
uBT14wB/Lpai26C4fKVWCCS/hOez9Kx2EaDeuIdnPHWoQmzR+LEX8SOh2UmYcz3notuIfc9BtUio
aSqo+1hxh2VGvGxu+cxmHbmUVU5OKwzalmdfWF/LusLQHEID5ar1VtcOcCtEqoBGgAHFUlZjcwiE
lTHGV1u14aBXYX6Hl8pYiaLNl0VqRIcLqrbE5y7fwh3NeZaNnNoiH6BcZ2U25ja/UwlqWimAJ66W
lICpNOwWUqTkfjNPEWOYB4Z/3ti5fK4STKr1LHs1tiF7LsErqgCmhBoSoHZRzHm+Tc5rXRDnenQd
F1zheOurqBtiK8nmm70vFe5O08859LWbb7TL1u3PrGF4aODhPjFlYeWsT3mW8svP4jn6md1424TH
3XkSe93LRTpJq5OjRn9qb40UuGBYLu4tG5DgCvZujxKCOJgRwgpsOnujawYlkmpVQhlbHK2gOtO7
4v2Y6LCWMJGwXV9RVqLb/OJoKR0uHI8pd/wQal3jRQ5uDMOKfue3TYeiTcVpuIO6SZdKZCqhmrmt
iDhyi0WhP64Uoe8N+tmM9TfFyZLByG2XpQluP+8yfYmWWAtDoi6YT+4QswLdCOPEYleYmDbJNIqA
H/yFYf/iXZaoFcsUk8iWkapo+Ub9NEQP4iMOv21EY2PpkQzsGQBMPq7vMcaQtl6UzO4uTAz1gjHL
z9JpvTol5xaycph/VNx1TuHAI3yU8yKLtp1kRYYbWwZmWx9ewAirZACRMgbXsOWp4TnotCE/l9Op
WbuXWIUwboOXK2XXSsByCVtnnYLwYOW1f05i0hIVEFWk4YpkNfLaLVxrHHZZ6DQKCVa/Gkm9bXZe
n5Ih/NZHLRD6pfOQ6IkQieBT04JIDF9mkS6QHiF47Bl2clfp+ZgohKFdH7Sm4kNfUV12gh5PEZ7J
Gv8xurh+A3QRBdLaaPyQ/RTgqF6mWbOeWF4wvNqTE+Zq4yjPYJXiKmmA64pilKjpk6pV7wQRIDlN
Oavme8WVCxiWxVypO9qR4ByFqzKazkZf1lDOxco05G5Mc9PSpc2F3QX/0GFNgHsv8MDkpdL8425F
l0HZ7OFzfv/oX4/+NECRbV05bfxBM+7NoxivNVOqpe4sv9OsP2GviTnZHkb2HU+8mYFTLiKTqUb4
CTwhgVpsuLfa5BjFo9m26UYVf7m37ZKdQ+y+XVjEGUzGfvt9welXfqKhxEs/YOtz9DUT3iXkY0ng
3oJHcZiFN8MFiFXkPnkmLor5to4CCDXYumRl7T2htbB0xe+10vN9pTol5Jz98ofp7UsubxUQHKrr
5r591IqN/Ib2jaoo4Oyx3CTe9AP1vL06uCJouNIVKY3FznY9yOTnkJ6ewda3t8ZKAsE9+qPiMWp9
Ru5yauikt+U0B4C3QanhaiLrzmKlrDxh7ya7dYQ9bMYGt+oJ3WrbGLSmQhnG9Txdi53pBhBkNXWK
CrUX9ioCOWfpV7g5lnPH2p5vyFINFrWhtCwo8kGcVvf/fYIJay+UQP1lZBRQBEtwiPu1E0NqubVH
zMbtsD/5kilHGvYMPs5/xnRZB9egcE7Gu9WNIoA/MINpUohUViAqVODtXVdqVAI+cOCLN3sd7wRv
6PIFcponn21yCJy9NZQIrgiyUzR+hRIEK325Ve3FkrXI+ZiCMGHY1zV52h79HPaSHIkbUXi4bb2f
foMc1Q9IiGEJyqIUp1N/wmnrjd6+GapE6gG04RNQm78K7KkNJnUwoTG4evPTMc4Np6Xd3ry0ibkz
uwzvTpkUuA87q9Sj6q9n4IxQb99Tj2vFH536FMfDhIW3iD+lSeFvG5n5abN2ACy0GWGx18EPJHT0
a6yuLqw9l3b7J9rjiDP0Rm9CIlxYstoavw/bwGyQqkUE22YI9jBGALbtEJp3SEIUlzZ4OvE819UO
toSfpFS0eeCuah335KrKe+5Cwrgbhhxp2fBP3/U6w2+hlNUxhaXV7LbuCrjZqyrvVtH/WFY9QrqK
bNlb0XeHGqVEytqb0OzNJumuf0RwerhmKZSiVz0SDfB4+IoS4rFsF22EfDTHz5sgyWkLZpbsKnrr
/+pE72x9oZZd1KwJrqzQ7PF3ia3/POfINx5LcAs9aII5tmW7I2HbdsyzULk3vWNYoOURjPYjSmBP
RNISdA0KCKbpP+rzHEYveztdL2I8xkwDfOUWFpDAxSWkHgROA4obzoSP/OU6tThRoK1PMy0ycEGf
KTdoMBe027HmvZZRQXZizzGFnEsMp2pMsW+CCrAMvyk8+XDrSc7Bua5JueKZRuOkfkO0DfolIwMg
0HOM/jItXQ2EWSIR+sM/f/fLfhuJZexZOyRXmNfgBPfWmauZKIdZZgX8DR+G/YOWJSGATuUs5UnJ
ZEfPkPyMx0l4Vo7WaJO2fPKvUOJWu18l7/ea9Jp09wYdh1IGHl5pHDZ4N8aaDCCtD7s0gAqmzG74
BHLkUpv9AXAKeCv007ILXynLV+P5zm3ZvthTYnP9jU1ie8HkB79AcIqugiWjUOKSGibFIHUMfWWx
ZDsF38qjPLCx6e5n786rLQ9/veI+MHY28tEZqfCfXnJWJuzYVFvRLoY7JogASIqSbJZL5adyi8yi
4593KRDfwN2DkQWpt5HHn4KPJsF/nu/fRq7IswZ17TAhKFxif4/ESRGnq1/6mAs3YjM0MjB413qt
p4RjA9qMPqVdjJstqev403u2CdrhnTuRMrabyj+wVu5716+P88yzU8y+3XBiZNB6p2Qm6dN7TWfN
p/SvwZLzoPhnoospq8Gfd6tC3tj6GGR6bkp0I15bWXeC/CtHAb5ePqmG5c6cLdcTYebMyt/XP4ys
9XMUDljb+bgMpVbvvCsBA/KZfnM+3L7f6hzfTIfyPbtYp5aNdYWJmwglC0mkC+ZCKWXggXKwb4gt
tLZeM06JaDevo4C0ADkhCpy0fTn7AC8G2jWA2Bt9NszB6o/NMClJYY5b94Y0K6wKN0NYo7dLpSjK
msm7VnkKM7O5+lBSd8s5XRAJNYpawl870HjH63PhoRo14BgN92yIHkAoL7zVJRYVp6X0dj2spcAH
7WZS+qHyBnj/PIuGz3/OwgdKk/ZxgmewonswgxX3gQ1gs6YITPB0byvCfAiiZAGLGEKCfuWfDn8W
Jz7P9C6wpX1Y2EiAy78m0bVwfmIHpBd/RKNoN26nHxKj2nEeRouCti2vimyY1Y7FNs91z9M3bej3
aQs8Fd9zivX70FZXsgSH4w5k+PyF6kgM1rZgXTbhrH8sWgDivHFVXyBSO2hCFfGfrsA2iuzp2F3T
RDmLj2oGrEIEPOEhVn3JFRSt65rqknKetY7l/t03WUuDSyIu7s2nMD9vxLTtCw38NFZNgzzdFSvE
Idk1ySyw07zSACH2F4ZiAmXdco6pj4kefHgDFlcKUEsj2gbaOCi7GyLqescyeVgDkBwYuZgLYu5L
G2A1ya061/gfiXnJUn2aUdpC3c383eTasfQO3IcSDBcnYwjOqavYe6rQMpD7RidpRcRYh6WVIwL5
GUzOyzHPWxvdjG5gmPqZ+aHcsSCwJ6bDPKX9YMr3LZNVqxY6wOvTC3hbMeOJWOdLCuwlM86EXddC
kXfnuEnefJcSdrf9vXaqlQEycqkHWaeEstSAX4w6hiUbpzJnaooUA/B/7SgRm0alXUFG4RMLi4do
oFTJJPzyBEAjGqomeLzvOh7lFOaYkTvHsHK0kJgcZg36M8Iy6TH8UhJESYlTumS6i2y0jO5Iuroi
oOpEnLd+kFyYeHDVC3JHIYujkTIIr7b6AANBOgFfNZqCyuJMgDyjPXpI8zlm2x68rI3wo5MAW1tP
u0x/zywC/6x4xFdDBT8OlYLH98MFSutI+jCEhsG269BomzEThhdvuP5/IkrelhY8NuxpzyzGZ/aQ
5CA5P8Jlv8ffU8/68mY2z77hrPgOMeh2l9r5gOVszMYWxxWdb2L1HCWwBBOBqEeKIub+RJxBzyDP
/deN7/9UNcPb2cPMI7NZ5+IlT0AIT4Kwps0zbkAsIHYTwJ2qQ/jOn3wq9hZki1k4gWwAXvcWSriA
B6k7fu4BMmXjURi62k3V0uHnHr9tPv1f4TtMQDVsHbld+Yx5c1k6GpYQ41vjKCJZen4T2BUPsWUQ
WIjGdRHdeEPfUPcBDJswVc8mo2cPZbKAMungbkXP0/z9WjS+blptNTe14qD5cakfCck7zOjPwtEc
yESmTFZRw34M4SZND8syx9SgvVKYoonQAfDH7F2W0HKJ4Lwj+bvAdOM4rk9BOL1+vAcmUex1jq4W
WlyoDq73ocpplPcJ8f6k8yTa/7g+5qettQ9twvaPwALp4c81c455vBtd3ibNVbxCOJ5H+BAGVNrC
KJV1pkajCIQr7j9ZK0SvyvsyRVTWhJyY7Wcv5javLZAbuT7qRFYrdIT50rssnYM8QX3ADIEW7xdC
Xkdr+5Rrll3S8caNsU1FBwxoiciJ0xIjSRdFxzfextRFS3UgJ/b8JBNvqhxBK5HOOH+7Io4p330+
xPlaRNKd7aGom+JW1DjPc9bmbygPIfnGZXpE8jwRcNhAYo7ikVsNjbaCvKXkE8uCxa0E9c08sz69
4k3HXq35+obLjoFO3kPuMwWnAYMkZ4n6VTn9slSkiD1DQ5bzvkfLy/j92NSFwXWJBpxdGgyoGlgz
bGRhVEqO9SUret4wLeNlWBpeJpS9OGtgCcxCgEsH9O1GAAmgvHQtCh9piw8A8Y4Ip+t14MXVSnVu
rkVessxn1N+jSAiObSxgBK0egG9y6PjuSTzikTyJzT/mF5YGwEQgcCYYAIRTXFrlcJmaOVXKmlM1
xtyU8qd6xE/3bhbSqfG83jVDM4UmuSl546TAv/8aLWd0oG46Tmylr+tBxgSVgx/JAj8ZcgyA+oDd
TVefcscbUspSMKNdiDg158nb7BkRCP0MaFap5cffyMPp72kREHzvrCiv2zJLLFGVT2rcTRi77Xcu
T5YSfx05n/+swNT+x3TJMulo/uYJ0EiAtzoTR4pRQazxbQJGgBHgy1ReK+1g9npYRAd1Ms/3/+om
Q8DX2dbSfuxS0l0tej+1zdZgv/4l6p6wyTFoAz92LbSAFdd+QkEDtgj6xnm3xAx3jIhmHSyMozxg
nvxl/vjs5ReAMmUqECsjPaJ05Xk5pxKTiQ93QK8NzQR/Rpn3VhM1loNq1wSdicQ6eZ7cRxFJuIfh
Tv3SCWrTt7wjz6I05kSm6gbRC68zhMghquTcsTpL8unuLJH0YyXC5GIoQrmjfyqcevOGkSbYheXg
GGobmbrQWzSF5fWRfZoWrlkEjDDE20rc7xiUknaPbf9HWvfpv0QDrk/lxCPcfxzVYvffcn4FiTdJ
ebzhJLGgtqHukJ7hkb3gh38CFL/XUwRQLDdQcpIRsvjeqq9ZvGrmbXaaRuyV0Ar5q4UltjJIBBz3
iborgZAcZ9q8gL1K5UJzqrx+PB30smGtj7MeV+N2vnrIWArr8mEUdInHlQhnLV+K22nN+oa+e1+B
nQv25wIqM5ugj9xz9fe39CFV0Ny6c7pkZFK0cp9zKYPMywqHkqGcoy0LaZGI9jUjIpA4qwGU8i77
H8w7/cvQsRYhxXbsNl3i0rG2Bo7Ux50vH2cNABrMEz4uEJOJoTwqFX1YLpU5dp/QeGh0IAco+IU9
JbiM2GvCPYOtzNQSHgEjAq5R0Frb8GWoOnmXhsb04CS0qCit5QNZQ1eSf5zaiT58SGyhIHKpsK1v
YeR7ZdgWQkm76ucVp+sbk3yPz9XvxA/IcdcOCzbCD6YVG7gwwbnGXVWK4WSkHo4XcoPuDW7OtBf9
5LqZ1bF5zAVcD5exILyCbrroSGkferKOe14NRKWpW0Y/B1uiCFin5z7kg5kRMLMwSWc9dau+VBEd
fylZzHaYeR6F3K+lgHLqEOo7f+orOjk8AUZhVeWT24YuwiFP8yqNaf8C5GssGW3fV/YEeD8fxkxR
Tu3gT49tLBHEJt+U+IgEXe6y9wefyTQZvkW2RvWlkhzZGsmuvxIBSb0q9s6wcHrCvHfp8Pn9E2JX
iCmiiJeIE3A9FyPyorRCyschyhimessuPftzAi76oMWxy/KBSsF3je8x/asbweMHsDZc8kzTruk8
8rOnFDpx5cfUlmCPsEJGbMBfMv+ZBtc4S5sLb4J1C26b1MJrk1cP8/7pFyNQgMrR2GXNtkI0qzNB
P74a1JjfuQEaUw5r6MeZDhvIUUBb0epLvzW3wFq7827mHVm68Wyk0h1U3CXaEeUKZ6tAFLfBEFs7
2Yx7C3QZNFTIlWSInCSYqWlzatd1LsgruUgJqZEmozSc272kGVQqHpNRPsfp5s/Q2zG3XJ4h0LOR
O3DyZZuQW61aIJqaXwFRiRsfV3lliM8zTn/0srFKYLF17BKAQOjgWQpNXEt4e3K6HteRhK9YVIk7
Evh4zjpwyRXtFpl1rwFiAsquPS3bf2+WDeJtsymrVTiqxviDSLJ6bbxWkPdCqdO93Nbe7G6WyqYY
1+MkztT7aAgB2KwiYcJXnZfeegPlCfbs4Oc02LG0Tr9UuX5naqM7s7BdLlzYBKN8jQp5WHoqIbfM
H2acMzOHaoS7ThDjy4Sta7gs3RqbmPTEhZJN7RXrkeeVXvPGyghghTqArh5S9kgDSvt4x0uPi5Kr
lav+5Vrge8mBKV+dChPU5mAQffC/puEptyWCEuZnhadUGQFKNMsyVZHw39GcKyFqkRnB5zLIAZMA
cp035NElYwnoXdYM+LJIF5T28bdYzXGdIk/ZSU12XRjqdxv720OtXWiF/bsSZdQOlK75hFuib+US
itnjO1pcijLwUSw2Zn7XcOssb5PtJfUbWljaUsjdRtq8efpK/rjYFXzXYpyqi+iZGDGfT64SMorv
N7LFkpVTpxCgjhEilsyREp0Hf8FcgYyYdGGaev1otDage1SCHHp+KScLUKTs5aop2I2vrqxtCsHp
PGS4o8AAyQ3T5h4u081j9T7cUeCEDsKMDygOWoE8BjYCUHY5Ek9BzxN7/CAR+auw/kRPqz4qTCXU
rDR5yhVcVvlGCXf83+L46yLMED1VZANpGzofH86/RG0TMi+IcB5qgS41zBM0Qk71ROy0itInjVN6
ywrGmjs1cvoNdHzr/GzRGphXsW0AFnMmiHv0EpkXvzNo/L9ZLtqaLjZKZudoejsDxhwGwwPM9nBJ
7kwXZhYeQDD0w95br2vZyT1sk+1WGrh5lV+6URGpKJT1h9g+3aHWiPpg6lO+J0ErbPursUR1Jv0i
shGfk/7Dof26rBIPte5AnVYjlHLmo5h1ZFhRDlDXsQrKoLIAtwY5hvO1u3HVkTt9ohpeX8pvgy7a
i+ABlfSUE6sOjpu2MfkN/xW2CLGFS8J7iy42C+AcxZkYoMqakUNX/FZEDPxjHO2yiI7szVfQSC/6
PIxaE8IFEsQP0Qgnl2LcuVT03MN5dzR/Dzgt9KIuczo9Dz/sVBJnlEjt+2xQ4oqJQnYKPLcOVuvS
z7l8jinVzDyozn+e1IRbrW3it2AMxrVWKxSU5A0IH7wKDo8dpbRKcalgVr+6f0dgNtIeZ7+AG2+8
3qwNmnTUFg9kO8TqLCWe9iy7Ful9sbrVfMNr3x0o03p8BODvJeU6tkEhQE+fi7z7aXByOE72CFOu
BW684SNhc0r6ertF7c1QakmvT2qGnZCNsreln11ukhZB+K/adSEw7D3v2b0/seRMzd1B5cvMTVVh
NAgzXdcfPiVOxvzIN6u1MVZ4hVoFialfQjdyjGSKXLC4RbU2RMwvIKPqSolP+gWOX1HqfHH8VY3A
UdcQcd/92dE9Pkr8pglfVVuqrMr39O+zwxtdSv+qIsr5Jw9rIsbcR15s6A/KZMEgjc/7xuEWYgZU
V9/awKHuXBQ/ASSyT7iCQWj4KdtiU0sbR1SGlPUw++Yyjx+5bNbwCLve75fWETiEdkX6WiY8+jgf
vFxQamhhNIpkORGoAuJflcwCy8kwMsYwERVcogPWo00YINBJJsmB/hhWNPDFvw+ruZp85vxLsV0e
5jWC0r9N3vFXzs6s9Hje/2g7+V/JFdxGTmAZLw6xSzaU3Pf5L7TGj4t3edA5HdpK1qPpgVCJuv7r
HWQYrlj8T1jL0ES0AjyHig+v0uUbtxm8rd38cmFGXwGGlE4JAKMAMzWjfCUPQ4kpYlNCgkgk+jT3
zAjBlihw/UoY4Mb2vd7HPuCyR8bvn02tkyjW4B06QLdQjPEZ0xaK834VrxSwjjP0xWpmW1ZxRwQV
uKczb2hpBgfyRCfMxP3EYD/3M37wrm8XJCbJViD2qQEjt2PDGy9hL2baS2G++Me0/eaMfHJqYDbZ
fHUKrWNYViSXEpYQGLUZudKuPSxpytfFDqdRnW9AIaUECifsK2Flm9pM8w+4NRtDDQZwp/cEOmhC
8OcOkKpWV9mvkp1hazGPkZIIDUrpoYWN3/+OnkyPeKJxpbB7/XERYP75pulRtSjGILfan29tXjUz
wUHoHAJSkpZVRq3+FuGw57C+7lpn/olpnvdrHA/zGad6MDjQSJF/feJ6oz477Lazq5c5TqGcwgOE
61+pl4WygRLn0eXpneeWpIGSBZRKVwNqxhpRN2tJEiZnsSNu9nJS5nNVbFeCOIiPaxLCMAFz+wJO
NjTTFnG3KKOO1exOZPCoqkfCXVZyt3NGcV2Poh/ci8iodD0b+9oTaSR+DEsPJFhYY4Fdvo1L3ht1
F9ifCFpJFvouZSl0JNJPRmbMfizNbExmGcSM/s9m3V1fWs+a0Lbyeo4npJUHS3qTjyUztqON4Opu
ndNm7h0g41928yVTrJwc0LmqCxNcer3xteLCTsHG4G9iM6Th9XsWbGSQaRo7qd6kwQ7wyapOi+yT
/Fcd0ElAyR+aM0qKtrevZf1jKi7xlnls+Ta5mdV7pwPBTdBtaqIhHpz9+lyTqAJkvzXDUnOXiitT
6mqBRtsWEJqcOnBVGtyzY4mY+Jqdra3fRMLqWOlIoBKkoXwFw283eFHWMpLia2P7cdhW8gAutdaa
WBH3rS7cOATApVUL56DJGMnaucMY5ngOQoYwEu6hE3BDTrog65JBAgvHFbGzaOS7feHh9BNH+JJR
VB+WyAHYYfBoiSYc8fEHIzE9z8sZIhVpIdeze/Ggbl8ia0MdKSfgIAl2r4/61Eil3b6h/OzaZhJm
7LGTRoOD8kQGqpyn5ypOJnvfYGKliLPpiVWZw7dQEauLzLhCmux8jWWJjiMOcvd/Y96OTx1+NykW
OnKMs+absCbcuUz+7cmK1nrHfWpN5Zjv4BBxDISyDpmKSlWS8fS8cJ5VosLyXKo3Hy7bkvskQ33X
IxlcffIQ4CBGpEp+eKhzjchVRTlV523llTNHNhyZ8lRS8hAmENXPk/6/M56bqVSrwT2TYqU8kK8e
z00Xh1MbcTo5JUKy7l0SKvjd0BP2kCTg2m4+ICbIxh5Ur/3xESEOAHVkekaZeUZ7HGmhz1TnxT+/
391IasgrY2zj1Gxwn+qsyyvUTSmZhBTsZ2XC12xNddr0dol9qNc+J7wFttg77h51AEyyZbvozvd7
jxuwKu9M92ddQAz2ygY0cbQwIjVHfR2X4sMKxOZi3bHTPMCXs8IAzKS4ojWE6qCCBvaG5Pk0BScw
r3d/K+FKLu3W5q7ylZA1AuqqX82onisqDBk/mw3eG7Y53/WCqnqAHGWnVTqVQsRIA1870ABJFUen
uw+0Mty/034Y7jn73x2MKf/Lqp8y5bUvem6opdSUoBXdtpUty6qLQ8jwIgquEaqs3GnwY2APpyDQ
CbgJwNl2pFDlaDr3eFBJJ5oaTIENZOzGfpG11ZvbitH/8WXH1cxCmihWyF4ZzHwcpf8IUTw96Rn7
gcaM4OSt9vocd1s8F0zg/wuItZU4CP+we7xwKZyrwWHDFusw1GVQ8ebRg+cE6ADyapbZtxLjoHOs
CoJc1vhEUkJBNRdUW+bAou1P1UqtHcgE6n7oXNSQTmOrlrT49IYq1erZtJxp4jKNbWzdwgymPyqf
sXCJvqMMCJSBNIvvaC3Gd2J2sDMrzjL+K6Cebsra9+//XSZ9i/ncw7XdczGzGyQvbDV/kzlT5OOB
r1sPYLEAl7Akpf4GwkKPI9TBdqvCL2p4wwcF9Y1xHy443U2ihUWHTJiEcqCAbSRkKYTjSlGkY3/y
rQkwc1q0JjNXm0xe8EuRz2JuOJra8YqvD35L1yum6VfbCaZFAiYZwfHhL3xDsnvP2NjOmiNTlZxa
R4J+TM8YVFZ61KNMOvS8ME7LeXHk7s8hNQO9Tazk2h1h37WuAktwOEUGTEOKFlyUhaSbM5qj+ov4
Ztwm2alxGxABibQnU1Cdt9EVlcjh+Otl2AGQCUA5sRJl6aETIMkb4KSPFBJMt9f6nRw0lVsaO1cU
y/yH84rbS0Vcs4eWaMk45PFGSgDVDpLTvnILyK9AvZsPoawkpTw8YwbrRUEYu0g5FZ3Nqzjo5P2G
0QRVW7Sp5476A0DRIcn9e0JWFYrAPo8TrzMoiqPWv7UgG7v2d34QayvcjuCUnqRy3V3Ffi9bQ80r
RUrbsdgCEflhJSDFINuvbU/t+L36lEyvFIbJkpbLzavRz2J8Kd/K3oCpmUFROKOsqpy08/btKyVy
CdK5ykwnUGafEchD2cFlPXT2W0rxmBHa2n8Q5UCVGnXMwKroKSXOyYAQT+pO4S0XEVUBywWZ8C0s
gDWMts2/Ax5MbBhis9F/HHTYoE2If9Ic2rRc4Zx+RfkinNtAQW8eslHqHJ+7n/1uiNUXZ1oRQrfR
qpRVBFukzo43mc8DV499l7s6YPyuLG1KPN5gv8mtFcsdjrqPNoOWOH5KKr23Uei96luOOgXSWqmQ
rgReTsjrV4ZBQquqmzACLhYaXpgLupdWUc82atKUuShUJ+cnQoRVtTrmDkQ5k0rY6HZlP9wvQBGb
Ej7PH4/9I1RiqahjFQTQWQvZmAz1zGh4aF0X8USnAoHlwtqvgAZtWn2c8OMFEBf+hB26kuozfHp8
l513I/R3+t82F3E5RW/Z3vImwNQwO0tPdulLITHbtvqArrSTdkrLiobSKGzEBCX2SFpd3a6isfNA
4M3u9JdGRJueedQPH8IaHXaSR8uMplIUnI3LiM+mOuNPcuSpuzJiMJmrw/7HYqjsciszd7U2O7Yj
YL/yeWcn5z/lIwerZ4PUrQY9Aln3RAeWqMX6xfQwgCNRRW/kSbgOS8+ws6lL4s5EiFBe/00bo6RC
tub5pMCgFVHHNI2QjdtuojOhOQcawowuPXbGoRv581f21vxLX1OXoPI8uWdLywY2rakcZIixhoDB
Gshn5SJ60xOwh2u5amJ+fgX12bcwypVxHD4NV50+zfs13VpPQEko7SEubkVZS/diJ/O2oI6l02uH
f0Jx31Qh+OrBr+u7NOrutUk067v2FvYkAJLM7uEq6hup+i5yJKQnSGlULkWH6sMd6klAql0XwRHP
p55HY9op0Sd4SaDkUd6pbDlIugicjDRfuIgR0DeCNaUEYN6Ys6ib8dABLw6+0sGoTtr8y3LdZp4D
U7os9f1SXGM7wbalAwA8jqleGFKEiAKa3eZEsrZfVDPtGtjgKgIAR1vjK7KFSFVULH+a3/OhBEW6
zbcxIy00AA9f87ZwgIVUcjwICVbwmV+Q6Bkr7UHBfnZXjBAl0aC6/0Rmd9FdbFozDkgjBsWGSMXe
ShBmSXn3MkQZPLFdiF105NEQpOvx6yk+/yR6vrfJBEnoWMhWGCJu+7pcnSTbcjXk/88d7GPKQ8I1
cPyGecfaWtRmcygc6OHVkV8tApx/aL0Zj053SkgcHz1XEwZ7hGue45jqPN7qB1NKxCt0+HKMCpyb
Wh1J6Gk3ugFbUH3Wu/jygIixgTMRVFQNzYCSqyZwJBdXyzpJ4TaY+oDERimXpQ46HL+VYHfAsr5e
zam+NshbyGPSwFpbK0rGNDp+unU9IpsgQfaoqYuTpSELt4FxbvGUPh1RB0TDBrhverXrWXqIcuxL
mU+RNs9eF1KP6iQCTwVw7nYNoG8B4HOB/fImJe6OZlTzL3hPa3RYr1GgBhEsMENTf5vckaJlNzLf
3qMcdGAEFmKSVXy1KDKQ8MZHuSHx6FRkwFPsp0XM+Eqa3f6O67iVk9dr/9RgtucJTJi82XeViict
Pr2rVekUfAFAqip+E6tFItUGjet+9N38a7cN/aQUj10WDpx6k0xy/MjoWa70PcLGS0+eQVNAp+ji
KGeyXXRSKzClQbzqRDs482T7tTrawZQI+QAqCSTheQnZSXWvB2pAqBCSYcLpBd6WWsZQy2n35ohv
/ZtiT0TqJlQoU2IC1Zvk0RmYxkjQF8y51CikBI0qPpeKETmVDm+2HqRw9Tj1AEWgFlq18jiy9899
56/lpXPNV3XoMab7G1PSllAU4KDBJ0OKl3G/NcPLQd//rwqw8H3NCqx+VyyWlBg58ce2w0mpAmG9
AY7gTxrD0wAkecZ54pJFl3yd4M9lAd75aQl3iEtRuk4TaDZJTpZh6dtyuKtjR3s7z/mOAlrvEkr7
JyB1GUU6Fjcog2j+SW6Am27Y0TUagdAYkG3q/MvJpyRcznrfAM63BxCyirkIXkhbiaf8iR7TEzN8
259+5ZTzc1V6Lnl6lDB+NLqjzu1AaVMWM8e7LANgC3U5JOBTZv48Qc4Yb4E+tTCHe4CcmVsZZy+V
7KheudKTrbJuUcuEI8doi+UMMrMFY4Ep5rp2stbh2qSN8Lg8nT4SDN5ZdAB7m3LkNj1LAt49+xy6
mBIsi57tWhvAZtkXqNlOMvxD5AMxxEX6QlIdc0n3e4As4UZWTwsqr2VUEeZktXFdoYb8PViWYiX7
Iqb1xWze7wLtqVu71Apr7DZLPg44gyZIGkE6oVrlmwHe/F4PiY99zsIy3BBWBJuNy8LBsxerEqa8
DLFAAqrD0kmLCb0QeMe+XP27tyaT/RynGOUWoxfguxkgXOsuV/1DuuuP3rWx2jHpn8eJoc/s4BRB
ASzW2EWVKMP3EdtkupGmEv5dM3WrxGVAoNqTgIR4xxGgzoyiECMtahEKwfdz9U5eV6aU3vQMPSlO
vB0sYmKaFcNPzjjsBQw/eZCRp9d0GGm5fztLPSyuz5iOIZ1EQDWzXf8xymUpyeZj9HHP7txclzVf
k1VRDprfUQyKPYwYP5C7ibNzM0gGhsrPBNkHnds4sjtlllDTKzKjEkgj5xsOC4KrkYpEeiX0TCPl
uHjyhpRnGrzTk8zTzGbuvJUq+Hv+KlJERbl9mf6XupBo9C6KvEhGpE6dEJHwvAEPvZVJdDWi9t/F
O9xOl1aGI30JVsOiEqGvYIcz3KxOkTtN9PWAj8MKUao9DGX6IoHYEsS2FNipqhzn7sJPhsFdkq8i
0ECChtVavLdZeHlla7Hq3MCSVJjPvehFCkXJ+e7qLzubWDoHiwJSJA9TvSlE0GTt5lxD7Ohb4o4A
QkD1/DxtfPqTBigMCltJf849LsXWcowrzfPgW14agrZtQfLu4XhjCDkhro9x2UemRJZ+29209q2v
p06QvM+Q9PgkW7LQyy0DW++3dsigQJKgTAZxOsW+J/L9wDTeonAYXI4t4Na23LOgLWdbKy6e2qdQ
VJKzZlsTo2fM1BkjILvATYyS4xjPxcua9zBd5MWNTB2ye0gZcQuEoAbBUZN5I868y2npCkcZE6ie
JFRM7oH3+NoUAz+ZpqFyp7DLN+lfP9rkW2NecX5GYi9y8TxmVLlwWgncfTGU1uNhbafp/E2kEfbn
KeVyCeeYz6MJd6oC4lP6iYbPvHnjRkFcdLZmIRrM0MgNNxk70o9W5H/AH3ahe6YIIcRhj6I8Ltmt
FrW54mwmOgvbNbB3hjUiwPCW0g2ePDmUf2LJO8cByct5Eh1RgfH/xq/XCjbGhhJtDyAi6qCfbxhK
mXFekEp8SDtmwnJvdekPwwprqkCJ+YpmjpUBoy0X8y/vfnOXPePETKdpqHtSwUQMMKGf0yIpqkJq
uFKVFdN9rPiAK2+VagIMaSxMH3LrI5CQ+5Oa1/Zyc3OSn5DPj3PA6SFerMRI3gWpj3xT8f9m94vu
Y2blhsLpB5YcsD+g8WRgJPw6B+PTPPt8dXX8ElXV62s3Qiapp/hcyDJ5/FKymawHIyXFO6aaamKc
bUBXZfoOU/Ijwu20QlG1duwQJtCCYUZFoa/PBc1rFb0L1Y1MR/tvmaHJzDkaGSnKO/DHXIqntaTY
knWuwWuLIdf3ZpgPW6g7HOuZy3ZmoWtX4S6y9whWwG5wSe99r5OvdZni+Vz7RXeN1Ju/SgdOJRRT
2xvwonKEiuhPdEhZ8fwZY1+UfNei2+VlWyGdF/GPRGv323zPlIFKD+J8FbiT7NrWF03du67JgNAi
RLlJ3PNk4zh6NVSFzXcu2UPaIC85N/8zN/l1ktMIttH2jq3P3p09F7bi8ZkiwmzClmkDvQR+X/Ic
LrxYfn0hXGJRJD6CW3M0VERf8BUGul2tziZ9Xatt8p3tGBJNQNjhgLmZ0sGHZMQHVG0HBE0Xa1im
hxC4bIS7RBGfghHiAY+5w7mS0ZwB5MUQ9TvpxUrZztR7QIwfnj/dFlloOC5Lii2NyTRNnwTP27id
FWBuUu7rbgz+cYRdlWzq46e7EPDv16sEe9jwzyxHOocTV8xVzX3uTvAqKAM4Ga1YKTu2oRHClWjg
q2mN7oY33pX1IoyvGN/yLD2L3G85+Wd98WZX2VgEYSF0I5gaIYQnFXReY62ZUx1tdTXk19A40E+R
2MXjKCtuIAVAqwiXA0UPMczT5bMxILj3R/hJKiOaTED7bZaPs4Fz7icD1UC1Q0xb0J37xI5bEiQw
g3rVwZ5A0l2hrXdJOdcTChdYBbUw7ptAm2ejpqNK8aXR+HMkMZUE9cc4q8F0i8UQ1+kWZPdzP1Bj
w4xqJjx/3YycN+9vY8E0JOodBK/KACCzUvACrr2uE45RILa0//y4AU9VhE7lcEmi1BoBIeaYXTkU
mV58LHY0SfiW2FO0yGj6T/ty6SOFwZZtcH/Um0uEDO7h7vowqWAtVhHcYi+1N4Qtbk4sZvjviSQa
UHg84VBMeW0zz+6zyGTT6VC09BWE4x2E7lWG2uJ49OdhBcILqo6IStlwObxjD+2Y+b0HS/Af/ttg
d1ZsPFZjGNd891IKm7yhKAcgYzTH3ME2brvrUkLac5SCDqJUMkcq21Vm3pp9DCw7mSFoA0O+ngeR
OeAPZ0VlfnBWlGX+r10d4h97U9q63RjricC8owmsbzIhEDcHhKiu8oJzTa09dpvz2/zRP/b2pokI
jz5idzXR3QlJt6Fb6pvgaPsNzrFgnislL9ELHr7oJ9OctVl2sDBM/uhEW0l08rfgC1fNwBz6vP1F
l3GjLLwJnisVl5Yo7lhfTUv//LHqFId8Owt41lvXqvIDJg+0Ubnaza9e0uPCL5gD/GVd9teP9dof
iaJ5SKJSBMqEHhKWDKFehPwzmDV5LwWMXJFghwtflI4Vah7CcJL3yqaFkSlrXdzyx6HhJq1nbjDM
ZbZpFh4jAo0mjvwUjWHpmQTea1O1ICkm5R9gwG9AzDp0xUxdnycgIQKRxBRGPsG2TXHNu2XfVwRP
iJsr8SFHwTaK7AXMTioS+2VfRbCnoHDSdjjZ1CDBf/23pPVZDOcbh66rJy/6F/dSqIXkO80q/7Ty
Fu6HMGrVa+qQI2eZCcUsxhkawSKTARLGM/CpmYTpA7d8BXT5UBjU0eID8pu5i6yW6meUJvJy2D0Q
zjNCPz3Peptvcd+jojX1UhwIB/88YAWmz6W3X3bBsHTxW+0Z3stGVw5xJpLNZVpV+edzvJjIAcEz
blU4rnmFG2pY7PkyVMnp6Uu5pEO2jrE4j+xU2rrpQvDz1JkZ9oSQskDGPbMHI/i5dX4h0afhCtSY
Y/o8YgNPBGzm+TbgI52hHe7x40JYN7KsxFyQkuECYYx8gVPbaomTbJZpjhL622N04ZbsMC3ehXdW
D9DnaYZOd0EF3e4CscNhI4k3t1z1dZ8YpaVcJpIvcnSGrq6dM+222QFSqwAflwq5Yn+vrUKuXEsV
uZkX7XywpZLwY/zPvq0YaDN/zZXtveAMAtdP2o8BPxrb8CWh2xclGcUHPTq94mo7Z99O2vmgdrIx
bu8N2t7tV2FM4JkISuzjve8B3S/0o3B31e98w2KFPWtn88o243gDRewrGJoH+bCj3rAbvGF9Vm1c
9omSLUSr7LC8bNEQ9pHKuOpbIh23bbKDUWCO1qjOTetuywBeNAyyvuVoVtqQbsUQduYZlARN7BpS
dXVrVcYcOFGpUve9cZ62kow6I5wiG8qNYbTO4MwUcTtfrwojJfkhLjyn4snFMvQModAOIBg7V5y6
qv5/gnQBI8e+romlfiWZPXV6Lw9nDPFPnHoC5FLLIeMenKFKLqo8oiOh/4mqd+xchkr2d9HytnDB
8Y0jT0yIaRSkAlortEQEx4gXPYE17gk6Hj7YU9RTLqJEcjwaaHXxtIyZDJ8FF7+hZV6Dtfd5xST1
2PeD8XVzzd6KqKSEYO9N00Ndi10vHP+5Ko0JxKq2yAy39wcPGKcbOlBPqHTAmcfVrSTToJqHWpCJ
zdkpQMiugjKgAXOO7XCgjg+sL3emewDseU1icYnxkDCAf5Mx6dkx8g382R60k4XFrx6FC0lByUlu
0xgBb89/q/j3mrRSrpCkRlwghgA1xHizsarQOha0O54nBIFvUPdED5PtDIuOVErdoCFEJ5KvgSYT
m81VSlgQPmXzSpGWMgxWF4K0mWogstw/YK5M2ktIKXi+emdvUC+bMw9nC/0+KbOB8IXw7444Aphh
yNPure4zsISnz9BPsMFAkJyMhOZlZxyUZT3thnOjMMEkEAnI2Ftu/xXudvwXHSa/EI2W6TSjzKms
PTxicx5YqBPmwdfyZA9i78tnsrg+4uZwA5Q3L75ED82FT4tZn5MFz0MXIYdU+Itz2FRRzG7yu6zt
IFTvzqxJJUYEMg4w21RYn6h+KwjZ+zb0iJweUqIfpBV84TnW7F0x+B/qVBwvTJoccFZE3TDnHLiv
rQI2uyypv4cVrnwWhpMu9DORbCCvBP3imBxdyuPB+Jv0cyqsSIjEalr+868/jIkPWGc35TdwNqez
OE3qCJrc4AH1riuXgXn9FG6Cu/R72o9DKN/D3KFNKW4R2Jjqxw59suxlsATm3I5N79oKb5iLUSiT
8JZXAvS3oOIGuUH7KKR0j9xsIzg+UC9veD+Npw+2aFeIW4ssH2W8jKU67ANlUzblnjYO6+kV//ZQ
7ZeyXj5lghH6JRkfvQgW0r69rxyQqMlmbgzD+Zra/a7Vog4n0C09RF6bXFu5HDXBExrRtzSWttn7
P0xfxC/TFhoqMdYDWMsVBasQKInBIDG2kRamxYpGZzrd1wZ4qnyAmz0I/aG+GPCQQNON7cirg1j9
pwxqK5YxwlMXnTIQ7HPZ6ru9dZ1XNFYpf3XsXuhY1l8k8Cm+jQgkVxevlYTzW4itizeLAvuWOfQf
7rN+9Wn9q6ChCJv2pUDIJs111AdFfHibcTYPo1PHl5BZcP84JlChMwqBfygrAWZv1QhUFFJTmjez
ylKwmlziEWbVswXFIrwQXmsvlpI61ceQwNedRSVW3VtHeFI+v+L/RjYnL7u3+aAodJKxEIVoaeXG
FUa+xMKQsQZtBrvyy8dOq4WQIfSOnBfQD1SP0pZcelEKW4OU543zm19RZXsutdy7fCXfeFrxj2ZD
5hZt4NzYDmZ3K5qKJcp7JzXG4Lhei8HMtopbpQzjMx9LzLHR7mWHSVpdiiN3/FUbLTWt+30Gy3Uk
QbJpKgET6zq4NsTRHTiQn2uRrwXEhcPYDDYGTB+/DxN9OZgRKr8/LrCb9S50ZRB0GUe916dCywlu
TmtB7flbUVYmlNjZuOZwJQj1tgqYzBtf+A8Q0OpWfLthh4dkjD6RZGOVnsC4J1nTwBYI/kaXXWGo
62yfSgOVDmaqAdNgzZ91PIVbWsN8iGsz+JGbDr44o7l6/n+YJXCb2wBh3bEN2nvMI1owid54N3ws
FpKcLwj+pvY7995v1eYW+kLdkvdT1khX+RoGSCLFGRi/jitMI2fdaqhiA0JgqatuSDeF7PPtMMED
HiXOVcG/UbauqyOFG5kkaxUiK6HEs9KaDPGWlULW8G3Tq6xxdl8XH/B1xP8HABXjoQ3D3J4czMsu
Ivkv1QOdaZu/O/kQK9QjhkgzocM/eXcC+n/66VaYT6PPDXTLwQNY5uOf6aHDe+ALZQa4On4q5eaS
Gnn6y1sR7E6dljnupUVfTHhOEuOwiAYkjMwP6zXcoey6R1cgikMIEyn4RUul63GPVQWj1JQpdVU2
+RDoNyqUdNDUFIHIMRUsAsojMCxtg1u91SoTERtrfvnqOLinz+IDwcvj1K+Tsyr2cnqlQlhPb7m8
ftIyNGV0D1g3nBGJaviEivxcTfT9LF9qiFqILFG3+tvP1whc43bTMWdGSfWW9rOGxb1jbGArSuvC
oi+tEV0veTUuAPmGNBqmwqitbVBwkiz9oIwHp26fSjZ/2/ap3dm5usWK7CiqBrAUUpDqKsvexcaR
ybZu0gKBc55g/NOUXT0Y1C+hslOuOHqedWd9OhN5HWvCr9PPyfxbngs/YGJ8MVlRnP3SDiPt5UYi
0xH7qWzTqkVkdUbxz2T0JDCqI1hMrbklxhRoZDObgh4+RUW1qAwo9UH+l2ScC/MOiHMTnL2gHNdU
GYrfCsaEbArxhHK7cncTmZpDEufc6MpWXMFbNss1wyWkYDT6cpDmlUC3NrBGQunIIeYKgiXxOmzF
/T+FOioj6MjtoRzX5H6lsVt1nAN82UiGrQ6eBex37EaQz6OVtCUbWSIymClT/wPez9r7Y14s5rsj
CU6zYzlIcO6wxoB8ohjap3+9uRjGnQals9HN5Kfgl+Vwur1k4uGvJRX2b5FMkl6Bor5Qff1Q8wAD
ItNN2o+Oxu03hBlT67ihExH1KI35eRlgG4Xq/Ln3VYJj/2d/Xs29DkTJceWani2469wMIZ6buram
HKlrxbRHzs1rVxyTZeqWuTC1xiQZ4Wtjz/lRPNFFD38oiYS9DRj/77XwaU9sazZjVai+jm39aFTm
Basi3nAGWcx/eDMGCGXbm4Fbo1ezwzV8zesGzXiDdSIUWjsXg0hHhJi3HWuHyHfRkY7jaKJnLk8T
cu7xRooychcEDN1Gge+TzPdY+BZe9hLvYNHpiYNCQh1SwGKkV7xVG8hFUNrQg6PLcu4sqgfBimob
z0mxpIpwSeVtlYbqkdKW9m23kDV/0j7NlccvyeBDNjFRN+0RC68oKJpOAcnRZhYDmn9PJ3SO9QRm
V1zf0G1OkKqpKi6KXiktYmmdPa6d0wcZaOKubyU+zj9O8Hs3tAyAjwizEkypcJqRQ6WRfnpUkuI3
f9/froxztsOdYM6Ibz6MMIEJlsQg2ybjs1ajyL+/T+9+dp0YM9SY+nQThNNt5T8J9x2MBwgFIQNr
clGmkfBNQWzdedcDrhTXnhFhyG4WwHVZMLWwvvxYEXI1IjTiXUHWm0c6TawX8vI1jthZ6fu7kbnC
B3NqQVrSkjUfmByeMaUC33mn7psEfezbJ1hPib+IheLPQv47WA1ADiS6A+iaTX/Zh9WJNNZxkdBy
hKOjwxs9L/n36L0Q9B+Rp5RkPn3cl6YvrIlndgLN+e5Qu3PK2ec/ilhMsIthOnSFKAmnShP6inCM
jb9g2/1AIT/IYSy4g0gUr6R9B4J32mp1OAfQIA1QCy0YufU/fYwCvRwZKeop2Buv1n0UN4rtawxE
ZjRiXGYe8WeZWoTpSmKuqGW+kHc8BmnP+3RF0uzdCZHgaFpRIzS+Hm5IdK++rQrutPhVqqLmCbnu
PPatinH4mlH1JpYrlATDLCyyi+FBLxygVmQy1GHM/7VEiTOjIlgoVG0Vsd2FkD2d3MSoe61iaJ1X
MsGS1n2EOsxL3yqUl6RKoUZ7kl3okYRCf6JgMR0a1L+Ur1wsB3/PaGhWcCDI38Aaz/WLZPpLoaoK
8vQbfMymCln5g3VqxtM8sgmv78LBNLLHeqlqNM9Xk0PkF4uIjy15fWyUcA18dG2zDdJIauc+Ktgg
DXI23iDscjAtmNNBo+wlS9UyuVHOVzMwRnaQLwMzCFTXILPeX2uPzhQsNbyJkgM29DewgYjSU/yL
O7UsqR3zaqc3FJMMU8c25KdqjZIIdYjFchppWAZoT9F3cS4rqeuJCO3Q0amI65tp6TcitEX56jMH
sVkNJs0zo0OgFLwkJZGuPDE4ivLJWUXyR0EwjbzZkGZATsIZX2Odjn+Rh8csav6hjfKVv6NSurjW
Y87JC9g9MsP198DiVdRYmJ3O4E/VxB+mLWuzVLcFE9FvPn93pJbZ6aahvQvw5ccWdPMUEd+Ue8Ck
CcNzmue6wzPoe1wQg6XVFz7popH8tKnJfVRz4glNsjlnddGOrIJi63UwK/nK5Xk3bJaVIVXCEXML
m1BO6YLVLn3ZknZMuCuC463Fvsbtny1TFX0mki1NSSuOf801jwHXsEJ6oRIuKvEYFH5dwlBwU2Bw
GHru6OxAFvVDMlBrw0764xcrT0m2NAgGd0G7WOz9HkxRUts0TBbonymlKK9UH5/cpqFa5hNT99vT
cJ2g+V7R+r3H1Plg3KWFP4Ymzre4xZ7gk83bgz/9ceNN0WobopuLAtAiyoVR+X7Sd/rpCbyHr7rJ
iPsIE3XH3C4nXQWImfn1jJW+7VikL7k+pwPazv/oLFnDQzX4BaFmWPKZDsJ4WIBdpAFkEfcLdl9n
X9yMJmqP4e+ck4OkwvI3Ua6/7O5ZhaUFS4BHA2SB2lHz1MEI6LsUGxYkR+Ud0iQD1rhaq3V6WCRk
OrzdZaz+ZDtlcsaEYZUYdJDA7of0VuRZnt030RmeIT1C6AuX84p8QX1tgYXsi9o62rfXcvIWVesN
Sw2aYe/aF8h0ueYBtose8L7POCPnstXaF6jC44jELuy4YvfeyRWdnIpdLvU547/RfXlcthoMucnh
Pd+1DbWU5XIkXTQO8xt+/gmDcEWP2RCqtq10raTXX5HNFSRdo0GsCn+PuO7c8B7edtb63uTYyZhF
oXXUS4nPDafe9ymCDOTHCGrbuaWsdg86UYeChWDNvzGE5ceLCC86ED5r8f5UyE5eqE2oG5zkzrqu
G8iLsNK3cmzLqxBl8dWGuJo1fMjmiY5+gcu2Wp3cyNqnqFhILdwmGOKCcQOJxXemuEE6zpybNMtt
01Sks9Y12M+1eht4BoGykXu2C9f+F7Np5o6eAJWfo/B0lO8vu8w6dpCgvspFr4lHxNRFY/52fAqg
PHEezKWAO8OQhGpTWto2PmC8MyUUU0Hrqq89l6hDyT02SWyQSlgxzRku/x+O5PKuxpQPVmVLvhdf
rzEqgARK9e/7zjMtyCBaZb1D9s0QYVh3RZ/Cy0+wsAjAboWBsMbbnOY9JE3k7alppOVln3Qyd8au
2FzabtwlhXsfYyxjtE8Pe8yugETdq5fdxd86vaNkIzYmnOTSum1zIXj9GniqFkAngi6883Pk+HGu
0c0IqR6ceryCv7SK9GPE2lvkRppCn7rjH0ixOit3w9Jp8eTYT6LXheHApmRv4fxZGUOXlvWSLNc4
8m9VJOAQq4T6vUOL3VgJhKo9SF/QeZA39mvUtFOQikroet5160y/he4aMppMi+yYaqfzIHKxlyDE
oMGJ7OeL0DAYSag4jc3b1xVnovJc4zpel6ROPonEvaq9AKVXLi9ad2ZFq0U+6SOMC9NIZV6Nuv3I
EARjbtgUE03F6BpQvgZWezQnzBLFKWXPOhldLTrZLTzzvfVREnzN1sCIONC4vUYGyF95ywtevhWA
nJwRsph9QZNqdQgC1IoRbQ24pvNYFAJjcRQNwX+0QnzUY+ZPVyqc44Yi2mxU3SDH+zrQ/iU9zAlZ
UouWsHRRZSWJCFsH0CxVvf65e/zqi1r1TgGfLQtP1KOdQzkqJmZFfZdn2DAMLVfDkU6/BWHlLCC1
Covfv3qo1fahcqTxT9/VDKUxSKO4Fc3ICjs6cmfTcNZOxsRoPjFyLFu2DznMr6CQpeKUHBuwKvKk
QPPEu4kPL76TG3/3Bo3X2bHFOfYpySIuCoP9bilYSt3qUz65rbpKTNhvfv2CGz6J7MNglY8yTk3v
bVQwjYLLkYS9mTgPHL9PZbgEtq3ZNJH/Vx9NKD68rEe/UG7goxZKkssJq0C181U1zlkOZ1ML7uLg
8TzDMWltEwiibimfFOnTuOyER2fRYT30bFznkOZYGmYzMY3OtU8m8tAgVtVGsYYdn8AmblYx5MDw
2apknSldCieXize2zqdIy97XPkOUg87JzA++Tx8vXeCFbTv4iM/Hr6amkSq+0ckGJmIHq2k1RQ8C
YrdUx3GrKASWSyOvacYWX5z6YalolAzPSRWql046VWlbuc8cMwYCSu06MVrgxD+xZk64zhDRvtPQ
RCs19+8g4ZQHkETVj2oYjiorEtliAupxPSpD1y4Ssxa2/cpbAgkcBCFYBzaXLABvqn2RhbWB4eYt
EdKRo0krPKtlLS1Iu4DqyTIW5CObpvpnpTBlIQJDuhbld26Dux6VS6nQCZoxR4GefnFBvcNGHOvP
TZoOMv3jkXMLhaK3NDKCW8zx3akqqWsTxQxqSOY5isYKrRu/zKois7OHK2QahXFJTRdX3gRhZ3DJ
HbfWx/0nGFBqYVURvVADsxsfSp57TdB1b9N+dnZ/VPiZqNjfD1p5Eic3L5WUXQDVxoI0km5nk1ub
GrNuZ4zBc8a4s6x5N5vgEA9IZFqw1zWjoh3j/Vhnw16QeeljTIINVC0B1pXDTezdCEKh7Zfy3kJj
M8KYgxZJ1AGEAWRAhOrtFuhcxsbodqSvsoefBPiuXQdkdxd0q1RviUDK0g1uiMsSiO89rkmpC8Di
c+WROWU26BjkmTnXObrUS6/9vkP+3cFInNSuV/2Aqm+NneguqmEJqf71rEd3Lqi39CGq1FEbjwrY
mHwrdC0hSn1FOQA+ieu4Qk56UnIMXH+cKJU9RduZERZBhCKpCXv0HiqIXdRWOtnZtCxnlxPfH6Od
AHIQVXcwumtDlZZ8PAPtPOCmccAEF7hDlyd2KOFa7CiH+YsiNGiOPCo6ev1osm9S+VBu8icSKxDR
P5Q2+ngKp9Kge5Hpm1oC1iZAklBrmOql58tue1SA0j+uuQn7/43Ya84MFa1xHXVYkfTx81WFKhMf
HtPB3L4QHUlfzNeTPbezSWIiNch9azPvtTZISa6C1ipfagGkTs6vd92iqez58SrQZQr0lPkQyUzU
ZhSh0qDkcvhnOif2eTDdT4QPFsJvuq3vARTPPCcvfE2G6E74qZXh1yrXNMXb0CAb8Fyd3ClPsfDP
rRuD9ccrYQGZSIBZx4SaKDblt8ZmHFHB27YUoEEQ02Lj6dvri1T2s8BC0o7MAnPxnqNg7qc6x6bx
eOj3n7fDV5Lgq2Oa8pmZQatXljMaJw4oNzhNrXqXvd3QealqTuRUajIsSE8pK1OikLYfCTUVwBO6
MfdXeJpg0enTBV+39Px6UdTyG/tfETztHLsfYbVoDEIxiqsd3nn1JwULj2CAI53H2BEVo8+r1ujO
RSh7rjDZEYMhwbidsqkY2h9vrlOmo7M/uZmvNaIrlM14kWmZO21jWUoTrPJ78OJl/ZWrGwJz8mxk
R/YuOtw7b94kWl4YETldOA3nKGbAaU3ZU4+uBxKSUhsmZJJcwXWw3wEmt1m2AsV+FSVDMOqcZy5y
zHdnviW00txSufk4a7Q/Y01bC2SzT59m64eShbXAyi+zq7ulQrDaw0DoOQ6bWHdswWc++GkCrldj
s1c1WL3+vZ3b7zP10ycRIgCbXCKEAGXBun6ZqgLAaCtVuKlUl/zAV2Y58QL+VXE8qqTk2ZKPZYzD
v0BC/VRnLcYKOM9UHYI6mE1DQYY6rEFKvBE6wLTdkph1r60/nw7ufVmhoSv8EBV0FGqOcy8wt5KX
p4E4rqC/qVrCB7bumNmjp9Iw7nIyP3t/tkkgt7OuxzUis8KN8+T0SiCkzEePPfZvogGpdxDbKYnV
T64z+7e8RbPL0ROZ+ScCkBygPug2BQKLF52ay8Rj/Rgky9Bo1g0Frk+GbVnlKB95X9j48QgASk3e
+6o+O9PWa30GT6wflyNUId349Rv9vYG3VisNnjGAVcnyltSA4lajIRpZBCbJ1aE7SAT1x4Ky2jnb
A9t9bSakvBNzl4GVWlMCtj2hFjnBuZCOoAGx2tU+buZOMXRyFjcZtK7gSV9ROChjfcJGAx2N7g3l
7qJ+fZntwklZQBfhhLYq6CeJ8iYX06jWqGG1K0/XysCu9tLzJZ90cu2nHXBhmx37inEsegYrLSwf
cRmPX95lmmdCBYJNPU4SMV173XBuludgeL/kBUwrIGfSsHhGuFfA4xBTPD5uC4lR6w/u6+4ldYlS
38qaDzEwXb+XYSq4g7EHtcrPwo7y4t6YleVPROvDaRWLcm8LvOGGPOLKptky2D294o2VT4w6UkX2
B+wnrLy/IsMb/VZSw2blMEemoRXfjDNoLHAPYU6/uU29WXEzLuex1i4xwBXqgFaF1YZKFzssnE5k
AerPYQ/SfgbQfzUc3Sms5cClXp6OhMPd/mhpVrUR+E1DcZktpaRLAJVL3DnwT/Xfh1GjZMSxlQ5A
HVbOldxwypAXGAD/DYtfiHG+qIZYuNf1YBkrO8BWPwPn99vjpVji92iVqE4MxnxTumBxXGAznH0K
4z7C82XKi5nGBKh9BH8OvLlswXvUGWhvVnfSdWT+vyGe1oyjwuenWhXrsbsztvNGjNS3hEZCSHdn
w7Flk5DnIGJ+UkoC0W8Yy11zLrmuGSdQeU8pGvEjkD6b5eicb97loWH8ZafhhrhxF4fnLZwAnmss
Wlw51e6p3ny3P9leMG6W2M4ZPTN5g3XjnTYycjfTsfWuF2M/d1booOwXNIM0M+EoIa19PtxLeSdI
BBGoZbQLfdsr8o6d8am2PW1Qjmklc5npQP7QVDKZxgDZ5O5Lk8lxbjJN2MiEv4Lu4pxjmrfrEcLV
q+t70BxnKXZAzyNOLzJPPkuJVD/naG6/p8kIKOLd2pm2SzvxAgYVT9xR/fjSzFRpu3mgS54gntVT
ZrO70zAab7wo2w7x91tdlOAUph1+VrFW+nN7JaWaJTtjB+v+06oxF3ytF1zTwbJzslMxBplCn1Qd
/EEz8cSnUIsgwYQnUxjBBRHIQGsxPZ25TMkg3vZ8AFyns4sXtILZvqTwV4l5AfC7fSPLULKJRZ+S
CN6Ac7Wby0efJeIUwcjcQ/jKoYgEA/ErpnlyI/3QfWu5WSNsnstq52DQLeeTmw/kUG98jbBm2oc2
kLTf3edyU3ClZMZrjM0yiGIRPq6jQxzc9tpkKNOtk7lQKw7sHW8ledsJcLPmjMRvP/yOL58XOM0C
WFGPN2XCMFd+PT7T9JhNQju88yC/gj/IfghyDZXCFdwamRw3NNfZDjW5z5PEUi1Vm+M30lGsI+BO
b1Uxy7EvSaWJNrGRmzAWLkZ/h+X83/veqmdC7xPtiVilNGODkjeNMndBhVINvgnckEZqHXFtLx3p
dW086r4HR2Vsv1yIAbSMjJbBzOvw5YqwugxfzSUhbSGUF38o7amvpZAush0Q/Vsfokv1SVZjY8Xz
z8tTFhf8dggH/G/A6u7m8s1fYODpvx0nkAphfqgDMO56P+PJpEIJBWUa4fXR62AQAvXNBE8usMn3
u5/Ln9IrVfDSNcpe0b0+CojbGcy2yoFREnYk/E1v7ShfTvVTWCDSYuvv/AgwxiXv8FeFnel7EacZ
dSuhnQJv5NwCOJHpcKKc+MRYiy4PVFvUyIciFQXmdPG5nY52O0WJ/T3ZCVptRC1LzkZYQi+p5hZ9
mK5Qhm/kHE9eMnEMFS4EoSsNwyMo+Cfl/ScpEZx/r3ZObipsgromoH2DO9XgO9mLhmawXZRF83UR
MhaO2X/kJrT+vmIIRdiiW9++7nild1pSHKza0hqpJppmldtLUXf3qPHiVvmQreaFA8V/qDfvoNBM
AFQNHScBXZPUMltsbrMaax9MfwLqHUwINxJIySaqszKQR1iKC+didPmuEKUKDB7r0XSvvXMXyRKq
Qws1IeMnIyVRxRFcwVcUFYBV+kSsII3kugZY8xyLUVb+SekCCwik4FRg5DYXCG8cScuh31aTyLSU
5GMy+p7zR4hmy0gF2W33B9HHwaaxaHhSFhkbeK3Yz3dBBELVgULoY/wqSenjbgEOozWKy0bndRI3
MbUyo7NZ+eZgan4cJaB+fKknAZwisaGh/wvyVi0+0P9S++WmKtH2gfeziLagXjHh+GRUk/9Joaqa
JaZa3O0G7g09lKv/mLGRAoPVuPHjEoK3GRUH7SK6tMo9QHy0nMvhQKDohJAjQ/X/H440dTZPbXIW
PY1YghP5Cu3C3Sgnyj/XICLUdrjrc6b/rbHjjwnzV1ba4dc1iKlm30u5g0er3kXrGrAmWASBOxZX
UWKHAQbUy3qwTU87Vq4L88NHCGo7jIgKVJkt7kY+aAN6g7UGNBFtg69OApaMvziR9AQGU0jIEXi8
n/rkoUSUtezXNMDjR/oAjbObtFXkUaISUDveqJP1+zhdZbS4qbZ4xaV/tq42MFovux/bgfFolOY5
NGcu6CcRfvXg/Kl/M3J9vKZaNEuswTABQzgItZ2YSvq6yBvdPMuTD4qwx2PD+VQ/hqAMWJ8PADaN
ERn/ua3j4XBejJFeoBI24xfHgiMtl7gJqk7qsbz2gTsWpTENH5Ori7qhPhISGpYKjbfXhNrdmSi4
uOBngN7DsK1uDFZWYsJJXaVU0KZk9tgZ6bQJ/wAC6MPhBzw4vp/R00c4Q8kcmunn3PBk7sewpZxf
cbo7d35q7ou8y5VgXX4HMVmjXJcdTbpGNxYCakvouE0MRSFuobZUAOWFgeTn1T5X26dsC3vwkT5w
VFT3xjBkcftqcpAtz5JNU5L4vUiZf/tqJ0yw9zYR3BNXNQ1ie63ArkC78c4xW5xb3N68V8+7RvpZ
75ekUE8CjcwrgAh/EbhuILRbdkQIUz65Q74xGSi4PPj9WF2lQsIK+mYUXPPUwOgBVZmFO6HNKrMx
+DJpRGQqL329sChfWkV2oFgGx5iEn6UrzsgXJVEpyY8MFXQth1/mORIEd0DyUvyQTW6foAziraMx
561wzW4ZY0FqDu69Hcwz3SsUJZT7a4XdHQ/rnIvdg6QT8dCqtOG57OUxYVxLjcLSxEVMP4S0k39D
RdN63BLKLLJrQgXMJRIcmorW5WMfo5Kw+qn2KSrq0Q9mXRGa3KDjudVn57wWYbwfYmYi7TwoEEpx
R4dixurEE8DvNkHcNL68A9yi5kr/saIAHM9G5pNM2KroCSPUHr+p0kMzYED8r2Gh/JaU7Q0cD1o+
QvUZIlj7CnuZ9iRCXOuuotC5JwZyrqFTH1Xjpng+yWs1OKcL3sUtazzKXkpn5ASUqZoXcPPkt3xl
yJ+BEdOZuYY4+j/6EuvNr8Ja4UZ/QlWa8XHTyCqDLn3ITOF9l2UabF0K06aXz+jkGG7WHJ8yYui6
GflrkVvmESThE//hSsx+EbfR1Q2lfsDKtj8MlOrDtKSTmnCcMIQAXu7mAWEMGR38nJmUnqHIklzh
QyorYw78IouYhFkGYyZRzCfhj4bsSskF38W1iAljn+Wzaz75TuqM07gsnhYTF311k2WxfboLAEfY
nmzKbAP6It86nO+mQYEsvpYLwNY88csfA5uMadBIdEKij33B2GD5hBT8UnxspFu4egsj8E9Jdk7e
4S4ALBN/T7DDBoNeEg06Y9aDJsLVOVltuFWAQbdPDzM8y8j2A5wfaa8jL5XGpmdIOWifONuGbfMu
z8mo55H79Ad0kmAyid0LMDIn3jV8kUTv5d1PjOe28WKjNtL0zMeZ3mai0IBC0ttNybxq4h91+QbP
1iTbBjWL8398cE0dRCvKUSs7MrCyUtnyCzEmoEt/DzVzoP+E6DD24Kb9YfmVFX/xh6VyL1yW8y2Z
mQWgD5WB3KlGH66AcgBGdxs6AtANA1iEX6MPzR90PFnYBhRVSsZAt3x5BC/sLZghTXBVypr02e8X
LoDTXmGqRMrFPjALgoHHYQHirt436htAEHhYIWoqnvDkHGt0CZK+uEliVYPXLP/UMnJcT+deb4K9
nUUyygVBuGnq98pXjYuDGOY28q0m0L3GugeQW5MdnEZ6JdYy/XFIqQFWVTvZO+1QTvsfyeulRXxR
pxB5VrLea7tiEuiSMutKHfOtwpIjZkzsBhHxijnOxz/SPFhZU0WKptKH9F6I4qel/nXMOPDgpo39
Bf6VsibuBK59Q8gntIUvN0evVRksp90Z95Qr+dM497apPR5BmG7KFREuevFnRoCJJ5oFbTu0TdjE
KOiyy6gzpWoHeM1LmLBmhOqFdrHu3umy0bxfX7F8M4BSdSLmWeCpzEiter0tmiWPPcxACtf41BU9
pCCBvL37PBaYI6yq297rPtLCbFsvJuJIwilS7PTqvALQ6iPF2wQzr32Mc9iP//N2Kcrj3Uoxoqvu
FJqII91GVLjY2IAaMqU9Tn6Zmqaw1c7Y9m3qiGRPmYq45nR0d18xVQgWJH4xbUNTeN/Tj2IyssEj
3zEEGdPKXjgx+svKE38izN5zJ0G2n8t6qWtwxcZxFjT/iOBv8uMRq2SkaHW5fzwqnK5CPfthgqIl
5PzMdnsYmVKDjUlEyKp5vQTmtexBFUKNh3DwQjfjC5y1YTC00z6NlPRJNt4d/cJehLyIIMEjV43O
OmgNpX6pnfnTQcCs7oYNuMQJ6adEfG/nf5AIQQBDJug2TKRGEO/W2JIxLh8SHyBD+cn2MvZETDag
5GMqOgE3JTLQ1DFrMo5r7pdmDHaoYEogP+jpMZb8YmlgTflqmtp6Fyp7YFemaV0SwWzpJKklmDxG
I3QKp0xlFjJnwVezru+F2ZHVjUbrRKX1zvDry6KiCl96cJ1k3ahZ0CDts7TU9aADfShtUx9onJ6X
LP1c13evC2c4/lcYXnn6tDgr2dYfvnent//6YR7FPAwVG4so+QGS3ZFuJc+vYHZiFjIjLnNXr2xz
DMjxIYdUr/vKObsY+VVZ0t2d7oHJ0+Sekz7Ub1Oo111hHAcS7qZYml1v0RlgMlkjItaVTd5NosA7
oiwyQuRrbGIHMOa9/TwAQwGYHxWktMJT6pr++VOlwMmisIR00YLUnuAxax5Ic3+yqESpMcHvFtLY
m9yrsMpPbcXCcL9qLHgozOeK5+qb3jq/hGto8XkRfa/EmUUYxB8EQJUvB6e32oUuvEDiy7+nzJLz
rIu8PVaLoGuKIlUhoGUjmuuuY5EPlWUngKzo02Zot3QJ5m26Ok9Y2RIAWVuuqGpRPm2JhgbxJ5KK
8w42PcPiFamdHVBd8zNw50zY5+FoxYgX1T1RYbiDxntTYvIZsIZ0tOEpJIodVnmTdX7z8XQOJHRG
twG08Kp5PR5UJPbUVdRMOcZK2Ao0Bfm6idjhc4oIfaowGW/uF2Lxb79BXC2Fk3IgtVGSPKIIWHPb
bzWt9mcBcbZGnyif/uUQNWJOduYQheKMXU47eEiAOgPK3qd/sI0dbge3xXi6j0HOSViR++q6cL5U
TKNAkAFj431biSen1LUFnH4O8nUaYGPhOSx/yGeJFShRaE0bszZZSx4VSaOJpy9jbho7u10WLUUu
AE1FXh7Hlc5l/U8PBSYpQCYYwXCZNq6OsCkTWUDSKnW4KsY8zA3a91WW+pqVFNxvbVVNETSGxtMr
OE4e0SCEyKRIgGyVwe5rnbUgGmFNdUW0U/pywGDn1XWM09BjjZMwAlZGZOMr8t2RjcUkBs6xmlmc
iY0a8THlW6CVcj7mJBszgTygMpm6hQlNzV19Sq3uHhdYJ9RvG1BSSXmuZ4eWPJJXHi8rWYzFcgnN
82Aep3pfInXtPii8l5Cd3MsB+A/c158PFS+9KCTNQmJPpc+NJrFjfVysOM+aFr3rbPIpR8W6GLQG
UEqSOdPWsez4cncdT6WRvGd5oJ0xv8e40sS+xfobXvq3pE1meuB9kkVYCHsukJsCv1ynTxpFBKU7
KfBNtAhetIWNgcRdjT8ggllLE7VP9tEowa2DR2cVlhMUbImQ40NXQso2JxDA+rnEj+23M+7plU27
N7dbWcSdm1OkfAyZY7uBsFm85SJVIX/99yzbqtG+qDpLByKKr7DVDTc83XZX2VoSgbuDkVc7X3ci
6KtsXuxQb+k7u/9z9uQOtvwRklHO4TY8a7CZCqxrKsmCo6bSmMwuT/DFKuW7fxf5NBKecFZ07RA0
6d87/rSIO0dnikjKw0Yh6v5hqPIwbEmZR8X8HqgiIAG57UmgLwYwMw7b4VQPW04JMIJUN0v2nPQF
rwfX2tqcZ0mDkfTQCQCX9+9TzhfkRqM/XRLcPpgZYDk6Uqr9pVAY+hJTEJuLXTtHKynWtbAlYMGH
b/rNf1jBpLZGfru9rIvgVjGRhcchcndSkuVcaCMDan8S5iCOikk1H0U+Rv4/cQmm/1azK0AF/lAz
xXuY8Mo4QeQ1Nyr7kGNKcSaP27cvavSc4A3L6MWOds0typo8AwIRFqtTqIF+E1Yc2jftGSfIZrO/
F5M/LLFAKKIle9LeFYyxKdmYZ+kctq0FjSMMD7X7tJOP+L/ByWILdrcqlh3/gUVXqaO/Xo2YiZu/
3lqTsK8DXfKOJ0SIPt1EOfBuMToQzLZg6ibmrezhM301I4EyMHgRZP+JA8xTQYD8Cqk2pyrxiq5V
F4ETpOh3+F85s4egzIxwgkST4dEU4a/Yefn01WvChiS2IynTdsNmiROAH37z0FCQyH2Fi+7Y/rJ7
uKaZEukAv4a5WGuvrNJGsgWVYTtV1sc51LpLubXIV3KuPmcSqY2QAU6M2b5g5UjGGbkvx/O+9Tgq
B6+rDf+iGd9VE9BJVyBxtaMNd/d4iQgYZp7tqaBuLqQP3iO85n4wDkHsa4rDhTllzCBzoSDiyJtt
W0RMEqgEL4uVgO4sQoAr5weu3z0A2yhfxWla2lOXrl1jBOX0wSJTJTjKRGLcr+S8nuTHRdqAwuUL
uqzG5PQVFMUB79ixpqOsvFZ0gRdpd0kRl5PnZZSc013uLbtD/x7erKF3lF6wLaEtbG1ra4/P3RN5
r1s/zMUmNjafZg2i+kbz+AJUsXI+hgH8E99LuVzzUBwBX2A0+FP2wQWaPxJkKrJWDvfyxcsegOGs
nq+K2qtx4+zy1XlsB6fYucUeRbZk/GXV02eBsdog+dqyTCxib9fvSO7NLDOc01aL8O9cMXlqChIP
ElnAA/h1tEbHGX/3MWhuvQ5gqmRZY7bOiNRvL0l0aRIxCe3EusoESorK2SDWqtDzti0p2zUecZR6
Xwpqjflva1X58K2lzzAkhZI4egqqZqAh2wWssrep7xRQT8MTOYkft+Ipw5bImdtd+J81XFp2kCP2
k8IyWTHglA+hx2ZsJEmoMOmF3ur6p5dIX+UVmWh43i2et3dhZg0UrMan95bC+XiFo5BOQajLW/1i
3UlT5tNgmG8mk77karHIgorSM2bqddQcf5U6BnMGCS+r554qNg1sohKc3GO+LlpKUg5StenUNZ4l
fqAtS6Ii31TEUGhholJjhg7tJ75SOc7qYREBDqYK9I3C5w+Xtp7yaPgQF4YAKlcooPjW7XqROtiE
POJFV9dn8E1f02rWwmbz7OhjAJgD87mjxtXQHz0vxqdv/do7nW0zgzkr56OYBT0Oy8S8lvZPjYbQ
Gu76fyY5bHrS9onN6GApnYd57YnqHxZz0/0nvyybTbXFPA87kxiiXGXuLbXVcFoJQ13qRimDGqN0
gKhaYlTXPqCqTa7IyKai3wJu5SqQN8BOXANcTwVDOaoGiP67UGGtvktkqzcfLf7d3ekNocxW1n1W
eyMcsgzgdnqq4F/72lTFkNDsq5HC6j/x0E+Ag2laUgsmz2gGGfb6RjkA9oJy8iwIz4Wm/ZAiwTre
JNp8xSeVm2SIDPAmR7rO9KPhsiQTbOSWUSfXpDZSbDjn+covhevlRp+4D9nfdt6NJyp5Nr8RZBGq
1mTIAaJKDTWrPif3N7zewVYJjAyAn9jYzgO4N4OjKDsfLEMxpI3eioho97I/IKuc7BSQggnLMnuH
pbHcKHMjv6UsXJGuS8ZqUv6Vbm7wsH4e/cqk+8R792pVXQLGOHiNtwo98Ekl8bkREHe6PBghX6LF
05kNZyN0D5g/HAf7uSBL/xwrXPDo2IfwQqw80sWZIUirqy8MydMYzA1kl4tC81BEl0HntD+dCFWR
CNHQW9RCmZTRdcJ1Doemj3T7p6edCGJpYBAYu/3nPVKd9cEcCdzMc9u9lAEWflqqcwVMV1aQuesB
CDy6MvgkdJx9HySKaQrVt9MACImUN4ywFuw4Nu+UvfJTqkQnzZ/sRMCoHHIGoWUre75CuPJJmGOE
GXubaw7XkUBs/FsiAd35YskyoGtHG3ltksgSd/jgQO8XaQuirFwFjIjQnpQ8DrzXZ1udchXCnmbX
ahltA8pBQWzd31Z9mJ6fZS077qWB7BiRRPfiqq+4LteL/mwAD4kurw8tSrX3OHNmOoiZAW1q/ULX
uFaEqdCImOIcIX1p/jsxnGbHdGuCD1mW+7ASdsGjlO0cQsB+/70aKPLnXphVawvLNbSqQBNvTH+6
7e3lvbdhcZGNjqZMbqYVvgEEEgZ14L6WnF6DR526wDntg8lwk3rbMYFUhzKGerpNvf+/sONmCRYK
umgoKFo+hLjwf3L8QRBsIb6qc88KAM1u0x/aRRcBCk+Aivg59QvdjeD0YtsIgX9Jgg078fNPYnVl
eTpwcKzE+lS0ro3bZwzSFzyts+4MoMZQw0+5R8CW6yQ4lpUrVi9fZC3HHP//nq98/WN3G0e4LNi9
2ECZQPruMWAqO3RIu3HWNCu3r/+rtOlntd2N2HtmidojrjHl/hH8xC3IHb6YKm1gCxjbzLBxFuGK
BFZ1eURC4z2Yefoa4x30YwaBlg3FZlj4rxSSIGPJswb9swUB8RRvgoXYqlRJeZMOvfdhz7yTFqxo
3XYVihnoYR+gydVxNWcAMGTk6JNACSBNyrcbUtQsYiLnw723CZqtLqWfArO1Bpn8O3QmrYuPZc4U
NalEuPSqE5pYHTfWOf/51R1jJjhXaoSH4wJxjpMb+ZYL2sGJai7tanwJpYl3Bem2cuQ3//BO9RdB
1UZHnoXnkXP+P1cSBNMSoZOAxFPPZzZIhN5UBntNfAIaFTl1l/8+NJ8PfMlY+o9viGfIPuGDR7GB
JF09u6WZWUbX5YjIqZfI1j1b0BGUJAqwOoPSY8nqBqH8ZEmaPPnmsO0whikvjC44SR+T+ikEe49v
0+bhVcxEGxEA7vI2rFN+zObXY4ojP2fhpVRsG5rJsqR+IUJ57RI8l29uxCJ6ENGIaYU+vk574wIT
YuGQzAM86ndShf8DBar3yNcj7sEuegjOL4oIFPfL1rE9Xl0021l3kBswglqtBllRYC58swwB/9zh
1B5WiFXnfPxtbhpPCvwUvA1pCV6lwmqGjdq4ugTBLT0LRCPHxuRvL/om4LMYEFc/6J/a3j2qwXHZ
E21bCgPEgIkAWQrE8F6VuusuKkoy07LZZAhbTX0uuo/qrEpXgu4Da658f7dKH1UT/lYJTLAwZgaM
f6FWfKQbVDr0QERSTBgEEjM1F5f/XVtXoCR2eVsIiYeiJKGxWana75iXOnjKjRPCTsx3U4ZdEeZ5
KQMFbr/ZvyD3b52Vg9BofzMVKFIWfsnVWkS2CE2Y5XWZW8hqBwh7wLlsYjk2xhXMYPPqYBikcD2A
vJsYzmIpGapnSDLUm95POC5iJS3qp+C7aew6tKA0eXaA3XSnAFotfhXMVAVtUxOncdQD9WIVSJL8
GAyQRqkn2EBhDmLJlRQ3zJgZWC8OOT809xS1x7vlggcEOmqafJ7xLpsYSc+RxZDtM7Xq3jDTcg+s
5n31BsNgc7PCjnO8P73JQGTJj5WRZflG8xlpv18s+lpWoUy8cDwv6ERhP6x0+RohoZ2+QFJy6NoN
tCVGTbV5PDwDE+DmlEmexX1QGmFC4r0hpiJEwuRbmVyVcCFZFeUlGR8CQT/iPiXQXLaLry8jw4Rf
xw3T2CgM+mHgETwFEd8KKHVhzo+7EiH93+p1SHn0LX4t9EorPQp5ld9qnH6uGO3qAKXjTniOCGDS
Npb5AHKtLDT5xOBP9j/ICYgmGH9L5EEkbyoAYBFlsgjirzxmm0DGuh09qzPzsh1wHe0mvc+IKr90
Vv0eWTbzrqUnb5vxV/q7lnLSesxFhAxOWVl0d8Vb/QvXcwaHWWREv7WJIID9HCPdCXvE9c76/Rim
U+0jr+tVIKIZvVDvQVt2/s8c9nz5vh9t9SSwPgz+eMrwBNe63fUHZZv8wiQvqwZrWh/wv+on9tDD
GClcBJOIELob+ArlXvwpAqzPSyX0KlRAPO2SJXniSHB4qAcVZWRtvfNfYXH4kqBYkBRLl/x99LwT
O8vU9QDHBIKo85iSbozZjTMOC9hCfjHTawT3aBTIQp98k1fd75cDda4bbRtQfDOB768bbLJKdaEz
RSKXQ11q6FgjiePakCuYcI4xPIKFqknsk/EPSG70cL56z/8mjNqy/7mOLrH4Fc+DAwWRq8InlhYg
iKxa1jFOvdvJOAEicDgCOoNEF4DUgoKez7Lompp6Mk/K55C9/k8LYosE0LKJtJc3cAjxylRkk3u6
Tt2TfzYP4DuEUwOrI5A/0zYGR8S/9oaWabVmyFj8+L4YKCcq/2oQCGa3Lhz4xVl7Tlv63ENB4xHg
Uyicn1ZvwWMlluGfzq8K06ebqqBHBuEPIukCQBblRIc17qBdz0OYZZyAyGVVwgwCGjC+TJKc/hkY
3FMv9Xq+3Bl5hT1Qlxf+TA691K7K1cLJwAm4QtdpBkH53DChxveTQFlqBcczapJwnEUXcl8ePZ+q
1JruIrhebFVPsGJeQa7QWLAsmZexKYK9fpEl+GnGl1mDfoy6nI56+PjqMoLp5zi8mIBMwIeUflq/
rGCsVe7AoIil9GjhCkniIA86wZTx+iuYWKfCBPEykO3FPsVSV+NmqFFgqV+v/IybQLVbBjb/J6jp
OHebLPEcdKRgwQwxTicvoI0CUAE+PaDY2SbO5vUeyE7Hf4wlUrtWi2RV/YUMaUiKLRq3oHMOrpCh
jUh1BJ94t48SZbuheziK0FuGqRxrSYlzgf3+oj0vsPkUEu9Q4aYShYVdhhJ282e9ab+WOpuEROB4
F+lD7IoFL5ZK2XHRY2/8sF5tyuKeGjiLObQF1TnqdWOxsoAMNF8CwaSl9h411IWrvobTIdSBtCcr
O50EyQVC/QT/MJ1g73sg05ZL7VwXs7CC4VmYjLxD9c5uCajCRdzNwNBB48J49Y5Zl+Vz8D4zHO6/
hWNihWl+18GHvbHRpch/lWcAdOPUEIOl4QSAUj29mUhzkXITZXq4+At0MnLR8JUWW0zCr/CQ9Osy
cXRXNzZ8yLxnHtfX3IPBRMYcjV4yCYT0zSUS9hGhPpdQlHGxG0tNJxNYIRehFHChnlqjF9HAigqT
x2ZBV6Va5EyeP6TneoxjRDpcE3Z44MKZPl/OUQtxiKq4QZfKBXEfCAEGNgL6siM/+RaXbDZSfMUG
voAbsyC4lEcMufmIZEU9uxx3o0mTJYvBWCszn3AxJ/KRZN/0vQmX6XnA/0oQ1CoQnb+wLDD7ju5B
rf1puHWyOsbwzURGjD1Ewx3wRrump+N9UuCxErKUogyVVnRpQTPYlI1yRrmgM+4Fbubac3auDS98
Xo4X6dZSBZm/hYZG5KgBYoQ6BhY+Bc2LeH3HgG7R6B4fe0XcekuQ0UXs03xuQbDjhCsBJQQZdJeG
Syni2hf64bYoTb4S5tTdVM0jGZQyNPaOfIbd3tMhRffSMcndzAzwAGoViZb7/zbSE++xjjzkHk8w
8SbyQHezYGaIujTEo4KoZql58r6Rx+LuiG2L7UbLYC2QWM78hIWYConOKJpvzgzctjMV9Y7mtoXj
Se6sGsugsgz1KvA0IP6JDOaV3GCmM/wxXuPOyg//j4yFOXwrNXpyU+fDLRpdkP+213/E73MgBoJT
b5paF0jOEPHKuQ/9N9yAG4VAx2HPtPF4gEoMg+jb6W2/s//+tcu1DuadFphiUCP/MdgaSJmdczkf
3Z0PTgU1QQ41S2ei4upcJH6OHuaMk/IluA2dCkyBgnRfXqQP8ZMsWJx4OutJJk6mXmmjoesTAKO2
NwJdycWvQd9qOx45+aPGYHmxy/TSJZ9DtbhfuTpDjQYMic99lapQavXdQZAFZPgutDlOZPIHo0p2
7wL4Oj9HJ4Xc1kW3tYlgFSznfZ6CmOpZuy6VeATSVsnYIwG/PZv7AzFwtZNdlOhXKsFW6RbZq/Sv
gAPN7H3QImDYOxpGBfwRhBlyCDJRenSslirKtx+n2r5YXkNZacf0KXm9ZxOvxf/mjAtJqIvz5ghn
9FkavfUaTg1Ok3ivKCr7yw7N4iw//w8y75HYZsAZ3fifpt/CG2iolErrBg3suH8LjTANCRiQXsvf
mQwEqQGnEQ2J1xyoRhTg5Df2lasYKL0a+twJ2liBBPmHHX9ilYd5/ey0AlYSX5LydSLfEuXP/HXm
DgAkjwBT8qnVN8E+z7+5ESzFHMs0pS24DFvgzasVXY5EVp9x5J5CPfFvsyFom744THLqqnTdRO8M
4Hotr0L23YOkhb3W0CXQXUgHGm0szLbNfV5grLZOpdlCJmqnBL2suZnr2Eckov67COdpNI995SoG
xVY13YkhL9mfN5/3eTqVrSgCbUx4rHS+JcUhdA4uIYv/I6j2V3RByDC0Nose7niDXCmqd8u0CjDO
psMhsFBtX7ngFFf8DETlORTGTH/k5Ki1NNKvJAbEjWMSLTzjixdfnBt6SKyu1Yl2VoxBS+AQyRB5
dvts7xZRedwJqaJ6h3I+j4CHlsdHI+0nYZZuJ5Pr8LNpfmi7nca+28yFAbRrqORA7Q+FcAKPQxiB
DzbJewxn/7lri76wzPiB8MLZf+LExKrl9BRhKK+XtupYyYbGmkmy8iwO736wtpXti7Q/hmJS3Loh
MEtNWjJVqBMLktZM81J0LI+QKWPu/D2Vrdix52K/5xG6emC1f2Vuzu7sAqa0hom9gBO1wgf/Vr70
OxfK+n+nLTMsNuUkGM4kPIs2ucRPykbCJm8k8DbofbbiP8OLD0ti1Le0zwPMdljVY4BMhs4/gbru
4BTOB4Vm8uqxgCm+f0TkHJnpdmvT9fhLFGxvspKqBlzMBMz8YBHkdp57s2MvRmRbXu2ukBF5sLMA
XawptcTGkA4nHf1HH71sYEKYfDGKBLKcyGuKidODdtncbkVurRuUkC811XgogSf5ycups0769X/Y
Z7eRsxKxhiBCWJCjOfIdKdPclqLEfgMhcf/MoCUZP4ADjj7jh5Tt66spDGdPVhn/r04mdyWoQVfb
7b4MDDywIaxcPkhJmM5PwiBNxyJx24P+ZlqAycXN16tLXQ25qLBn31HLr9kQ+PyYztm1ZJ7Jdyj2
G0GdgIUbww8JH7FtlomIFxC2Hm5KoGdnu/L+fpM2pIePSQ2E3wnJodmr93VXpNbmw+/VveRBQWig
UPzyE9zc0du2Zw841hBMp9BUwpFaNydESi1lQUoUdEG0lgmxyW9yKeMAlLJF1/K1XLBfstQV6gFQ
dy5vStPnzL0nF23GMfcEQ4pFF7snEi/1785yXiPDKJKimz03hlQ9F2xwwGID600wgGjXM0r5vqZL
voP3iOCfmMTHW9b9YEVhum0cirqx3hvXsHg+NOt4FrQ3mzYihCycv6fyTfZ31PlDGO+9Kn81JOSS
WlSPRT3A4Q8Ej/JUpprdpgheYUcXv+Z4eLl2i+AklgB/Oi3gN1BfIBgMpEKoPT6DIIOEoE1QVV8v
H3Y+xpJwQTlJ+4e9as02yg9I+eWjUaWyW0cFhu8NcnjVr+6S4YaBHJLb9YvaPiJlIJzrpvAZZU1c
pXpb1aWfW188zurl1yTHhN4hAICNSI7SPogYfEBeqZtxi8OdNBowp6gPn/oUT4fdoW1eIG60+q9u
kTwIyQ00XkJflHtwuOa2uBO5yCAspnkwJJRMo36LpQpKuvNduKs6865LRQDi4jxbPEdV4MrnaZtc
Kdk4y1WEV0mKaa+Ur/pv1s+UYJO3ujnrL/0tGl5scHXoffGnr35dDv9JNhhmFgLAablTYv+hM7wG
8SFBN6JenPhmLwQf5KTsSGiovFre9ku0eR5iIrMWRG6PsyY6vrSzgcQlYLMMBAu7h76vdjXXldzC
aiSNbW1PonYL03lbIC19JgCqXHOQcVN4tudaNrosEy0HZjXQHP1TA1ZKMy/Dd5sUw7U+FEV8Ai89
9l+qKFNVasoGFgke/7hTvyDbRwAU3V5+q9Kr0zGz04ERz9AbLOZM/3qZ65UQPfGPG6e3KoLPsOja
NF6bEXe0n14b+uu/sfd2zOe0dqylPqfn5YLfCaL/HoNtY2MeWll5HJJhRvNYKZzANRuExvj7L70K
cnxpG5jGHI0fiierJFxaWvbsMVt+5cqJ0XaAimk//6CC1QlBdt5ee5GTcfWsHm16IGzNv6cljj7k
g5uWAgkwPD9k2YyTu+xDJVudOzjMAadHBFNR6jc3xi0DOkUS1pcqx7UootX5JxfrmTPJGPPJoEa8
bmLqP+R5/sGz2QDi05bTvKy6+SMOwWvIIeFgg+X8N9LF70OnAOhq/eOTVq6wU0ByqHNF0pS1B+Tt
0oy137SO4VPotvv+wFh5r/VbmtIutW5T6fPXitn+BgARBPf+LgE610DHQX6wTQA8TibP2+03ych5
toErPrUI6lPvhCOsSbyWusES76VIMXOaSTDA25vkxa355GROhD6sRHsTmvAXYnVTjikfaIb6XkS0
xFVzz8E1Er/3lpZ8F2NbvyQokVZm2fkjwtyIm7r5ygSk68YMyJ+Y7UEs+TfrEa8DNolg9qQJoTX5
WOrTzeSZDLcdQaf+hj6tIUeXxmAmbnSb2kSG0osaCQwDYeK0VbdhZnFKFlxCngE7rQdtypDYdzjW
Rk7Vt6Mhl3aJymgT5j6cIfOF/IyJk9wMIaOLIoeQSEz8VDwzpqGMlZmX2K3FLHb1hzu4w66qorb8
0abkZZCiQiUyoDusoPdG5xRUPPMpbu4TQQzhVZgN2oi4SJNyr347knJWetL2WNStmuFbFUGe35/u
vp3gEyBjDazep3KtObmegl1c7FCCG1M3Gog2N8f3u8LWb82hbFFSN5PGO+9a3yjyE+C3ZFfB/VBx
ZPWhjzC/XV0TAiQnqBaNiR8Cv7XVkG92Lg4gIgYaOjc77Fijm59YqT6jm5YzpOMF0CqTgH5einar
V2+tWoUma6mak49vVCrb+C5K3LPgNLjpUvTh8o3gk5ZRoF+An2KHUxs6sS7gl1Xrt9xsfpG1KQc0
GGMveJCYdQiytihWTcw4VMFBmQp3cE67H+GRr1dcE8uvfw50a9M44meBdW7aLHbdbYhMc6N1zd8y
ZLRmNG2TqPs4Ao7FXa/mGJEvWxPm9OgkG9TXpDJmXQO8FCcb0vgE/8XjzNqX/iXmyp3XB0GUK1E2
hOpBayStt/Gp8RtSEOqe8Yjvhv43YCnNGg9E0DNkG9lXYNbybKDlziS2Te2DVb1sErzwr29RUtA5
qgtR9S/6vYzmGuZq9RYB3EFMNfO8Qz8ApnFGiRkfqR2inHsnlrr+fxQZ+Onnrr+KkJcgK9o3EhCN
sF8EgF8vWeuNoOBsYlTR2P0QHqewrcX0orzD84phb2HIsrec//boaVuFwb5t4wASF9jA5WY5UwR3
UfH/Agr50JXpRU9Un8Od8q+SxZfFA9dNFjZ6Tqw4a36nAJEjnwq20EJj27nogJy/zTAxpjYXVjy1
xNll8nGroCRIm+NFSSE8i+1wjnulTIwtSjQbpDA+cRT03atLAlDkD2O7G5vqvPHOCASuaghxRwhk
BblV7eGSkMLiYXpKRO8YpI0n+y8fz2VbWKrVDGpzKC84BVVGB4Sx1ST7pCP4bANaU66YmhqVe9zp
23JgiZxhfnE6tY0jjBwjJpvPYEFxSnvly8g3OhU6wbdnl1mUHtAUgZ296OMxt1Wb3ov/IirwPGFT
eKZB2u41EKINvOatBwH4Slppko8eR9vwcTmXsUjJvm1HC4Qeg55EaVoKSUHw85kzlVkgFubeBPlu
Uz/B1QPP+3wMluK3+DCZvyBV2zfPvcoUDOiSAuosDH2V0Y2LfeKfUWshPxOcP4yKw15mmKbJHGmz
5Xa36iNvdsGhbo5zm0Qe1VaSkKfjV4D74HTQq2dzGAfVqi0wNTI3yRCI+rvC29ak3y389b/qd+kb
ZrV/CjNlKTA4h/jCX8C1eS9sR+HuBxoNGVZep0MtPS4X/xJ/QPI8QjKILMRhgxu5K4DwLcOmY/Yd
5GOnJAe9ZFUd7/PdCAHYZ0szc2v+18VptmFW0a8zHZP90PQJuPisRmoAYcNBNC/vFC3VO1bkiQ8K
AjGOty+ErPxGKoEYphCY1L75ef7m8pQjf0hoaJP6s8N8wx6hDPz2wXBoXSTL6OGDfXaoXRxn6L9I
1e29O0oFXEqY80OQMkT26buJcdKhiptZFY1ojnJDB8BoosKsI+3HU98RFq89aGkEu2IFI+W7/UP3
iwjjemk3F7COAibdRO38ndtegT/Gq49Fvubh9IvSAFXt3dNlOHcc9/7tDwbuo3YJkG2ZBuybw/0D
rR9COxw7tIEsBZU/mS+c9WkN6LY8XpLpWt37d+Q/XmzZ/wb4larnfBFCvPwuuCogWFtj5E96CYl2
AO5fCteYVHufbCeztSqIbUPDvoRBjn9Im4xe+rZCAkjO1tJ6XH1EMF7UO0gVkWT0A/91gRAZlxEc
P/j5X3+uuDNItbl2F/RyjbrWJPhS8kB+PE8KH9ioDcuZlYU1J8XncZsmoAJGu0mFCBwm8Q0hi83e
F3xbmWljy6S7Y7h/k6iTypVn6xm+MdZwXHJGClzMoB1i5wCV2s5GSlFtYARF3fCd9z1LY1S/gOIG
oOaLUDH8/OPPnidID3YUBu62FQ12GIfjUg3wTqWRBpBqSAKpFASt13gwifa3dwlciVVen0iwZKGY
Zfw3lpGF1yJ6BNiiuZuX061qrsROpkyZJAJh4aXSMycJ9ZQLuws8ce4JKkRhS1qPCHdsXrFLjCE1
CJXlQeOD0rEzkyC5rCfgI/93zC7BGsAC+UdILE7NRy+3s5quieElyKAt0qIiAuJqdf6GsNExaOc+
Ct7mvXr/ZZx0bimEW0dHfYu2+tVsEHDCoEciHg7rKJltY7SZXcnhfMmR7w0QBlcQqJj6o87q0Kbg
WUEoi/r7ZlHoZzp12A4rdVIT+3byJPphE7k1cbSDzKnTeZqjyWlI32hxQ9oW4PdHdxhNklBmSY6p
Aq2wtD6OSdlnw10uPmGMV355rjEpBSfGLjCf5buGj/urMAorA+GvU8tINZ3DMDmrvlzZB+y6XZg4
t0co8v+c71cpgaC5UGavdGlfXwXJcJplcwBEAkRiUOLT4ueBbRKRd1+M+6shKbsL2eLT3KFnVoIo
/rdoi6M6eHmNQmrUL3VRlQqLZvEP+OVt0mxXUO8Js35jEpoGRxA4OG6ncSE/ic+OlwJ5ynHoYedI
DLqSI2PZTBgbXxrFKUpiefJ4j2nAh8hCtOrNA4Fldvv2mvCtCoeWNGkTVoDcKLlbfc6lLplnKItq
Qz1DgGntWkipkREGYiHYtIURZBDXuqIZcPH0o+XcxoiLw26ZVkrG+YCf5RFS8IBq51rG2D8MUmEA
VWh4CRcMb/z3U65a95mwB7n9jtZrVQwJG4PS3X344ET0uHPwFeZk/aUEfoxStApv9gFSkxjKGyLy
s25nIyLweQjdehOgRV9huDRJVMTyfCvwDDo5psOLvozWFvY8TE2SCH/Q4bZ4KBYuGN4v9wrGhmzQ
JidlPlhCZEh8Y5pyD9xMLhdPxLuXkFkaqG8qaeLa3ZoAel5pxde1ijIKCMn0QMf/khgURCj7Q6I1
s/K8vIJ42yOyblAE5EysRmf32gG9xsR5dUeSC3cX5m6B+dsE68SMoq4W1SXbENPlaIV3qyXTZuHE
eq1XdbnPlGbFzSwxKWrcQR+WYNfTs5kdXatnqlgmlWRIzXzaOEE2ZalywoCYCJtFVYawwRMBfxAb
r38WK7AX5qVpIBiE7Entwclz0ECeFfUDZE3yTu5IroExa7BW3cFKoYgubNMfwXsCKw63wZOxdXsC
T6o93LTLc5/nM3/xFkfPeD76DelvE/bnLCbDBPNK61rPM8P28HYNbcXMk1ZpEkbJLU/Q7BhR0DPi
eoUv7FH6sydawXgnvDEtFBp1EmoFrFy+VNqR/vex21+lhJ0uyjOYy+nDylpdq78C51DHcuFQjC5L
xR3LZEc4jZtH7vs2Qt9Foom+Oa/lduTaAQ0gzDwVXFrb5eX+iWCXfBLg+ykVVEEAkLFFbe1mUwvE
tOS08rAmoH9rB/VvSLSXo66AlztaoxswtSVa6nUar/R3ojEhnSa1V830YOqnskNOs86UKfdHljeS
GbHki9yl0jX8quTnkB1RLXhRjTNkBI8EG9mU7GTNYDPbnffTt3oSv8J43OD8ZxF/UVYMi2Njq84Z
5do0NkdOsFx67B0eli76j2lTZJT+MUOzjxP/ar8h40NEC0FcAGzmkcJecTTxZIO8HPhGXIGmELsV
GxOhdDCyEgGmiySezt9Xr5MvoLzhvs/kb0p2UkYBi5jVvZOGKkUuA//JNvOdQOxLAXk3i+hnyB2p
ktnuXL6aRsWgfLvv7Nu31tg1fV/xYxpEoNV8Fq1qSziYjDOao7dt5UyovGyZwtuDkp2elUqnGOtl
Cq68Yxs9EdtenrMnFB0IFmhdR3Qmd4vSREx1Y4vNFs8TYf3BRsHlhfBUmuZi/NurnjjnxDkyBM5v
uGUHfQEoTiO9TXlM8Z3Wtg0iQGmlGzpSHw0IcBy89x/jHRyvXd3GjrP5An4J9LUJW2Ed+QiKzXXv
hA8ukphmKkUgEoutf7be/8qYbgxSL5Mhar1RDbYLTGoCSeJH5541o81JgI5ZKItnZGIa/ddRMEBC
XKUX67BbKXpjVwn7LpxjXGgx1u7QXxcDgXmi/H/h0DBtmYdxXEbVzuUdL165ezDH+AL30QcWI1HG
RTdoNxRAQWUspXNOKbyCzlo8KP88A2SQ7qrM+7lyg0t2V84w+bgsJM5dh7vZusQsIEETx8g8Kfmx
65tm5QU4t+kB9xlGNE6rwEmQsOnK0V7p7RfPsf9amMzAx2Ho8+/nlqYF23Os5Ljbv/FTqcRFqqwG
Z5vn+gzJL7xrSGYMBKXpzNFMRsGUrKXcQy8z8fW4Whshasq+xxe+iLwwT3LIRMRoY/SZEoYR7tFK
ZfDOcxndm6BHrfwj/Lk4qnyjh9rmxb2r5e2LVxDAMSy6aF/zz0GmRFHdt32vL54jTnZZBbItEhQv
EM0IvP/HYYOvbfATs1834RYuQAVanVoX7ST+nKxC6S5/0Rg12pCZOJGQgZNitIb0nFsMLnjfL4es
iCOZPbon35lrwsM4MJ5QPj0upV1JV13rW0ZrFWB35hZ3+2P7kyrgDM+iBf0lrRtS3CWhTtpsU3XQ
K5aeUxVLs2VemULfBrn8tdHkorV9rBiXyr2dZXUwjUfbPvbVagFyssr+T661R5MSaTuWtVBBboGQ
0AgA+pZfNVTykkW0bRt+1bpvFaXI7nyc9yxwIfsRrwUHRA1KARC5Y5w1rl3RzQStTj6oMa3UeCzr
LFXfySTREaJyJ73E3fiv6umXgr48L3fziFQw+WkeZyF4hUodCp3eMwvH5qXy+FWf71ve35Wc4FO7
zXli1DBNNBpwJoaLcEdfLSLTF2fIH1nzNkdyDisRLizvzenZehOByAsyHoe8D525lTC1S50nNloI
3Im2TqN1Fpg4BHbNEdUTMvVUu4dv2rbrskBHs1Pw73hL8/iGpVjSYv4JELph6uuV/z84WHYMZ/gk
ver+Erwk4MP/kz6aDcXY9sKJiWUCNsMjtVs1OBp8F68qF1EqeOCnDLkyKd/E30iqOGg32q20TCz3
hj7lKUQIdxGIPoSCGsG8YBOSw44K+/SiYVIAOjP8XAbqHbjHMHZ4XxlFORSFSbk4U+inPaV2vaj6
89IIyAwLZmv95lKxx7Gv1PVC6IlVKvN6ojs7m49JAL4unyckRXymPKe4WHBunavrxOP9lcxVWSlV
3vf4LB/9bH0vU4dMyoUD2KzKJORcBE5xAwooUHsbsXsnbkJv24xuqkbnBRsNR2lv70z+IBAAm32W
alJ/+RyiyvQg2ZCqQgUORGWGtSAjUgZwWKzV03KofTdys2XrfnSYd+gA1YntAYsKGWACQNXUJFkr
YmEmRvl6sotEQw5y28XKNA2FggVhV4gawt3rIYIaM1iXV3BsHWQLo2SSOQsrfqqSUZVFyc9F+K0F
E3XDFMhg0kZmkG8B9EQ7r4Mzfmowux8aowtB+ksySL3Buob4A8mD0frNOc49CfJKo74LZbGtmlrQ
5xkOnqdGZvjdsYqG2NdGsd7Gx3QFd9j/hyweQ7c6T56M69EjB5q0v8pBZt7IFwY648DGsU4mMz8I
5TntsoGG4BN+ph2B4YMPExT5aCFEYhY186Qcd9HfnwUFVNPkRJi0QiNgr7Z+IVzlsot/SRfARFi6
iYppyMGQaBxPx1wJ3Y+uJvVfHtglbyvxX+zh7wAkZser4pJlDTQeNQVIQRgiUE3eYPSwZxoBcLuy
OuNVyy/C42WpeE7s2IqSC//mTqplm9KOTA41NtoRveQemryOgO3iOimw/RDsOdxtFj3RNEZD3sw1
1E3VDKBiCBsVMQi87QdjhC5qKNuj9fX2lE86F0+q7FuRPvChfNwPqwgTJC0yODU0aBu5u0PNv56p
2bDXlkI1vHuXnfwOD91CXQfwUJgppwVDpyERilWqRTMukUYGm1/dR7x7jaoey2zo3lUDItBPnpYL
9YifLN2QRm05CHqVIERvwnvLptT6d8dOoaVwg+ca0S9ieVEDhaG8ITUYWzEDvxFIbLkR+4ZyqTOs
jnxB2z9C/3/hfEcuZ9z5m9StIn/7gU4s6cTx5b4TFHRoBtSwJUXI1+y6Geq1WeEIbs82vsAd+DNI
ilpqH6/rDsNtmXZ71O1ebZ6f9/WETIVUXbvgpdHLrRToubUkAIrSg6OBCDjpACEbUPE1/8OoZslj
pvZuJ0DNfRM2o9nbFrJPBrDLN96uZVQWF1LQLaDNrtLAaV4T7sYr9z82NK6pMvkzXrUTdSZ1PSH6
FNT57+xJu+7TR6lP5ewbj3ziC/HxXGxYc6TfKJNmWyEE5zIn6g+rrarr7lPdOAcppyHGo9JQCj6f
69SQMHZwEAX9rHCO9OWb40HzeB0Qw6WBWtN3Nud7g3LpXc7/KNGddh8jIymFy5aglWzgdHu7nTTi
mIHA9j3fBzo/aWuaflwY4LA+MVG2gH0OR31AVKOiNTZq1e8EvqWp3cn4yQ8A32ZieDgaMNFVvtgP
3sdiW5c9zCSVTOtzCE/6a1MSYFEPKmqqNusj975hVbM0uS4ehH+9RDT+/+Ir/hpHRMmJ21wspWAI
VFEWKHVJXRQ1YHtgyP9gH6kdPy+N+VjEGLPSusDyAl6+1OmhPY4ZOWFn/NJWEZ0g9OArTcAA9EJ0
nurjeXGNYR4wNdsRaR5ZrBhSCJgsSm1iDPLUDRagczZ980rlWh2U3b9vonCuc7ZqDIOqkSasuvrq
1W/Dra1QeplB/Lgu7ORcP/RNzIqSrfK4ZNzydP+uzYDUpKDy0Fvpk+Sq17pBNoEircyJG+/qZJXt
cLkhna8vLz4IuOGAIYpuZXY0/VWey13XT32oEpZt29aaY0Gh49yl0w3R3lnakxWmSOcSr+jhePcZ
1t2fmYH1F6WRzH203gacTLhKjBjvgPboDsJLLx0+p9s+PiWf9YodXmNjJg/GHEAb1GQbqvxuAGex
3HhE40KYbYNAcI404LIuQMmdzHkRW9egi8d9V4xwJmWlg7XxqiadGGrtgTaRRl4VATzRzu0E7tK4
ESMsuDxjBbQvCXmBwhN+afEzm+px7GPo8coEbdbKZfsoQfqxvZ4uOAHkqAwCVNTC63BqCu0qAn9V
Ht897iuYmYujtRWJn7ZHn/FiJUg07PbPQ3ZG3ImCEqpi4sNLazE+H1TriWtTo5dmSvYvsi/YN6AU
kzmlLTfiHcEKjc0vmZg7oyhze+iL9HP28GCBykYgTcRIuOp3/PFhEucxLUQ0RLeVZy1TgC35gIUt
Io7stNnZg3PbaPz8jGGkZmy6jFv2KO/LUfeKBBhtMObAHXb8eIhqaKD8EOt6ghh43SGdP0LIgqrJ
sRCEQUkrCa+r9u1eeEwgLUL4b/NwONIzAKb5bXtY8F9r0y5kbBAfrnAuHsJ0t8p7ZAmg+35e7VJC
e8bTXVgPraoyuerVENhKt644+dIGv2mIUitpoybJQ2jLRV4xZlmnOT+iy6jzIMDopeQw5DgsP+0A
tINT6oM47QOt/pdmWOmApHL253lzXQxP4qWaKB7Aaukk/b2mTGPEHcVfcQ+ETCFluuT0DP+RL/Ha
0tCYqj7KFT+mVDIMd7zciCxjIDqJW5C05DUuH8EyaQAsOLr/Y1yIl1nJt9QJyqah8zFg9Xa5VK0X
yQ6mC2lcGhJJt6RkRpA2E+odCIV3ngpw3eb8yWzm5qCQOiu+Jy9TDFUsqJBJjsBILy0OGgOY5VJM
B+sW2XjoBcK2gbgIrZ2iRz4cEHT2YMu14YYEYY5x5prhZjMRqdB8L7ZO1F5G6Sj4XHorq5SF8EZ+
SUUJKHugvqGYP4p1Sfh0T0RRzvEzyoVep66t/SLuK6105chuBd/+wiHmW7hOEFyHJOSJHtpaQ2Ll
MBF6iwNtAn/4I3xY+7CqZGriN2PVQIE7R4U7L5ze6h2eeerBpXii2vpK2+YbITyRkzwQ0cE7+2jk
MGTuGyfABTX73/7GkSpdleVC6pjDThYye6chsFzarKPAdMm7+1QhXCZRryETX6nSUkKP3v/Lzm8w
g2h6+LiLg6iqEAw735UdqmpfpHsY3vQt2aldrlrgAvyfqemmblIZCAjthAm7v0n7yWmeqBWza7c2
HKaWT+0H2NUiZUYbX4q/nLDX6OLGuxndQ21I1RhOpBAMbj2xGCGh6ACcQS/O/rvczlXFoA27C4bG
9qFVVfuRE0xL+1JCrCESeAh28hVhCG7HZfaHdofNQsAOwRhmol3mOaw3PHBVtlMbv9W8l8TbVE9P
PwSrij5m083wnb1r/4L7fICS4ahtXyMlhe5CQpmbKCDzjEemuvgfiw5VecF6SkmeCYhLas9rEgTn
LGozoEVIjDhJwuMggZ1mACzblFxPrzLkms2GIXE3m1BbBjErwmbOQ11WYT24feAGvzQe1AaXwcsI
wdFFhZNjv1BURGawrHpYf5HlJgLT0UEaW552jRwGLG+vKiqz0QSg30QnuCzuSETPWNGSidgYFT38
K9KHaIsDX+z7u0USGhVu7ELwWlB3KzuLMghWWlPO1kVPCnvIDrObarzmmYZmmWsv/Dv6E9BVRXcq
5keifozzFE9AcelQLJh/gADU0oiNknSIwdN4N8u1IHh7DNWpr5S8jj4xvoaCVs1yPBd1Epb07/L6
S9Do2QI2Zppq/2Gj5xZDqGyVlWItCF/HMlqCXAIjW02InJXVN5vERoxplhxgRTkuj15qKatuVGPW
XWa+rckNicglSG3E33EDRGdIOZbZQJPz4Vg6s2vgg5ZKijLrvPD4NStrCk7vPM25AseEIu2AOW3M
s7qN2zdvuaMiPsIrRhWQM2YI0Q2Ol8FhJGi5GK9QWRX1EZQY6AuL9w+Z5iPeF/YkoDHwV+OMDb+O
nm12mKPWSCZSewyGz/mjiKyY5oEeAVcsC7qd9p45cr55KKEYzAyZLEU1inKOxz7qtHKc1nYZYq5t
oNs4ZQXNztH1duXk6wI9gHzlTO2EQypTprnMComNRYmcopzPLQmOpcruvzjE2gErbgHCXNXPttSf
Y/ipxwFHmfnowrdHRqoWSzJc2r/aEKL8VFxO9ITZzDWkch4mFVK8rooLxqpuYk/xEWa5yeeqMaUo
BCZIskHOF3H3B/2kvI291f0Q/YsH2nMkTA+lJ5gtEIhzA7+qID90S/SN12hhivpjdv9Kz1shOzRo
bRloYP22eToCvJ+GU5f+2kvcrLFc0MVUe3GmycaHOTQGt3ytauHZ+ouKtT7YWyYYprxUCpHsw5wV
l3ywFyaLl/OvM/3YcCkOjD+3vSThK34p8jsBtavYRI6P09FqTUmnkCzjHy6Fq7Ylj5InVSk2fMW7
Ku0KxrQKasvZ6cKJnFRrtB+tm0F4jFxFr5r1zZLGPa74h+/n9e7kjVtk8FG0n/jls14F6BNkA/d2
n8wwi6DWOF8twEG+CatNoASE+cX0/l6MtZlqfnzwYdaSYw6T58LLurwvt8OeC65hsGR+tc8AlnLZ
/VoOr8QO6w9XYqhxDMryF8Obo2PCTF7zF3puhy2W5yTKKWp8A54utRGX85ifP3QQxKHesiEnw9im
1ExNiP3045jZwAVenrCRs7hKzsJ1icB3u+jc2Ybi/pYLRCj8XaYAt+owAzqFjgvDmiFS5kYOTp0f
nfM+Luq8jFty9cfY401K7DH5SdqhvInFG9i3git/PSr4/nMBQmK/lqcX4vn69W8BGTA6Lu/wZvOO
hkim1ioADE7agCKtIRAgrsUQ6vlvDeM2CHiinWssSX0BL/3jn7to+m5j89GqUp/sQ3CtBeMtWiHX
hcYqeXSznXNi3f6jzXSP74y5Wsx7Z7SAEyiIu+tISa7jCS9nGSMcR3ixVcohZ5PTrwdbh1ESw+t/
c1MMYEEwMx/jn8mgvrI5uMyqzFPu8uSx8ur5xCITwmOzlnQxC83gT6fMM9k7a/geBEqz07sRHh7d
KajbPOoO0qQYiad8e22ne++M7sie992HSc+j5NgsLgab/1zdYuCFrbyJrrR7wrbz4T1UWJ8J5bbO
VBLKCZ92Gjs3mjhvBDQzS6ec1yEnaE1g2j/jGGlfZdzwe1nbp8KX11L2amZykNVwyPiRG7PiXyJ0
eMLRVa+pO6WzTgN0oDlUqvSzdZgR5iEjVPeGR3WHwrvJe9QXWwbyiilM4jXeV2dcrY5nuUyAvIP4
vU7dMIuCkzwT0oNImkOyFMc7Hyv44vKdicMv4idTNzhxvaE34df2/U+RO8lVMccpI7+7MEP1JcU4
Ga2WGJeifF0ipbiJ3rYCzQL83MzTZIak/EnpkvYhMAr2N1BnihqHlT0LjYlBKxMCX8TMv7hgBmEc
ZuGtsHaopDwT5nLvFaDQDKhWyvb19Sq3e7PBpx9liANSi2/J21kk+whZD7qd7WK1IeOaj0ARFxs1
uCDIqYcQu+6lPovShoNiFwj2gkI6Dw2UbdNlL2NZmOCRJ/ByD+RRVJQS3ZTWP6b81GjRv88BJy/C
yOZdrwLqJHMfKijgunE3yJMzNgt7VlMv1rp/wVelpi1giPmYLW8MiovpicpnDwT7RNd3xP+Kk0RL
SWq0NxRvnncpq8Fy4DJpCcrRybjhsS0Yp7QXocbkmi3T8kyoYp9/KTdx/cWzOSMskCTEkGKLIqgu
G5uPwUhZiI/a+4wRo+PRy/KS/aZFLYiDG8bRwdoaxcTpDm5eEAP6yvULiwpKIZoZyuVfLXrTEBOW
F/By2xMQJcXOJhxUXcGZbdCWOij1sFqxb4i2yTZZVFsqrRT615dTLWoh773NkgCtPa/3zZUvGu+t
SFRtKpj+R/sh7e5Zv9ezuPa/hO+r2rBsVegbddC1/0LZKclREidxjQwr0kl5pufE/39W0rvFPQn4
PDYEvmdq+HI5GV1Q0QM77FNgpvaHho2XqsM1/rXx2xboaM/iIBz9iUEkQxsbiORiCeDWGl5pRqVo
r20RpqjBf9Ygkvt/Fk240ou82Fd04MANXujwaD2R7Mi4/q/S30kIqPgRbq1kYoFgde7H0KmP1zb/
OjPw3Sv8dGgrJ7lrS8Bj45EoXl6lnXmSpNtXGtgax4MbZdRndvNzBCCxp/yHGNgDNsM++4yWdoox
WC+t9P8emKZ7GXHmif09RNY6m1Ty/nzM/uJFqLGJaUG6lRfeJJ0odki3/gKa/FH1q6nvGVWLbD3j
4UpEU7RRXo5xiWfhxOef2EuF04rMZSC1iNhrslOPjSAcjaB5flSfnLG/358wU8Ks2awT4ntAQ9Gr
MxWS7a/D2E5BJivWxQJstdIuuOeQlRxo8nOdHpLO6Ok86YI6/staGnJ2ebZwJc3c95zRNug5+9zi
ut0YYerRRhFJYsA9rnP77RlkrWqRg1V8XVxs8V3axViaXozafRw4/eE9tOU/H7p0K0czoSoFo9aO
PkVtItEZ5g+itYBOeLhTKexoVTdgerAbWhq9jnKkp1mJ4aV7s4FeRzczXC4H6IH/apetfYH0rpgG
oM56A1+ye8YBRfiwOiGanU696TBtFN67uAe12GBkOPOSrPILCmGucFBsWXHXr9ezM4LFHhiYSN+x
d50/TnNQipHm1kbsugPxGYuG7RUb4L8R5HTMplry7+FK6e3nbxlaIhbkMponEJ9Wdxdve2/PQX/4
LMxwhFX1BuxQWfFeQqHWFUe9FVYku08szp6ieR7yqIk1bDM3BG/g2daDXleQDTa/gip8J9ZeZG/S
xnl7Id624RBDpbYPnIMYbJHuGUQLF5Aefah6T3ar94V3YMFGj5eh3BC0wXaBpuLPBH/2KEpt7XX3
QAgW4YNYhJ/1dXoRKGHbXfyzISOYDDfGVvCpKTypf2K2WLO2Qn0CV0Amyq+KOFyAlk+xZSfa2KYT
PPi/f/xbSea8gFnIYxfVbVqeForgSrtPavQSehyHZ4u0sP/7lvz3+4fFZ32ee+jIgH0EmVBZS4Gg
OtMK+KpVM4qwhgs60nU7sKuqSdU1yTsMSzldBoH/GSgfdkWz7YU/tPUoJUdrv9o5aXaxETVspURo
VmCRrPn6EO7JWGvg+AGoIyvdGG22hbqPviUWvfEdYfA89wPWw+LQyp5NM2odw+OnReWw6ZWe6OMo
LQcz3Sf4QbHOtu9B+ZQr4U5M/gu8Bo5nCKUSLj1j496ymlcxrgEcWNc6hUmapVSs0hBPfjxK1DNk
Au2qC0830gVfdrZSQJ2C22ssQlK9ohcHmnRmSVUK3fBoNHXShJ0mgX3NwpqXhWj2IZuhHxZ/SM3P
CxLTYG2jaXbtHcD/+62BTwIIxf0MtjIEsZ5IPQL/5AdnejEmzFsxi5nVkOdxXn8yqi6GSIbj4iDJ
2bLKsq5kIawlZcTGGHYWd/OD4eU+R49ish8NZm4TPkmBBWkSRbBXfjQeuvAO9nNrg80Cg3pMokok
Jl5HMYzqt4XrAjCNxEsOLkY0+/n+Hbsdz300oQPxtL44xASiORPI0Hb/EdxBUupyBT2N7WDOsAnt
rEUiElcdNdkd61C6++WrPi6GTdniGEmCAl5NR9A2G0mk41qY339Te1kl8Y7sGWPgCnyHJfXu6Sv2
85tH3FQ2UWkjZ9sPlB1pFXKcVCdRP/dZXIef/+DNLG7zffGPCzH4DD6xhPY5eAL1D16johYk8QUj
wvasG+nlX5dcVbJ2N1xmYnE5+9YR2wLMGeTrp9AjINa6s4esr2Jje39JVrdK3LrBPtJpMq2FlcJS
jJ5HiLaeGKBwDs3hJHQCd3rX7YUc6h0HL3leAIQcTHBoIYBlDqsJil4r11lw/9TDg1vJbj2EnAU1
c26sAIVQ2bhXTZAE21i93/G/tU6G8KL047dm8ib1MdnUiu5qzeJGTE4dm/7OH2tMbsZZ8eVfnD8V
pXDaFfKQFZZ9/Jd9VR5+2R/nUhhslgcbaT4tWmhGypSMa8mBc4BarCTB69xW1xprulR6VkIUtXww
OqhLnlkIDcUuNRMsRYpKhAAGQ5c2rTCinXlcBBvp5HOD2AtMQZ3a9JVL18XTjiaGdqjI75bxGRkT
7OLGvPYLisc9OndTuGe9ziDPsxT10ZkzxrZNpYIZM8R5wk0GG3M+vOUi13WgcW+o4kG21L418Olu
DhN52q05WmxAvtn5rmW9NnupwAl6tlBvKJntdzCRBFzkofRjozsnF3C1cEONLyiF1yLpIl0nfRig
fNwuofB/mWayiMsfKNjADqVhcpx5jfJmbasFDbVzenAjhmo9pEkFelf+nboKPLOOdFTEBtQaUzWw
+qSyjX0A92ztVoEg7MhZX0jBFAJrVq2pCZa5fcg5F2gKFvUiMDQjZ+TFJ2c0r5di/w6k2Hy1x7xZ
DRZPOrmGAHYdJBpX/txPDCOAMnzlJRiEGJBMSyhFDLzUrlCp3EPbdM26rUcuI/JxoISlHXOvN2k7
gh90K7Uc7nUH8Aj/YP/9WOIjzYTP3kDauX5bDzAyyuiJ+TkMz1/tmxygtSB3bNawg+F+9eHb2MlD
RYKzrhKnH8ATW5TVtOYqncGBrtbLDeAX6yfdYNLMQMdyxN1yqVJLgHD7mPB6Rhk40EYNdiQO6bmA
zPpHlgV6i+cr1VIC2XJBG76qNb/A6I+MK8PAWhKLC4FQE036bEZT0wXdPEgs5JoZlmD5V8GqXGhB
SZwisnIqWurMKYLwOixI10BcjSpEHF173LBLUyfsd4uB0lkSBGt82KPGFVrtbGa83h7Y4SA45ln8
PGJWg+3VaE3BFgER5YLky25CaWIyKyOZTpbl95QE3ezfZmGUCdGNxROIm62LkRJRrM/5Ye20JKPG
YrgIigiNcvoCbnltCanVInAFHfz/B25MHnjBK+/bxhhV8HZEQATA8Im2CV0LvMG1ZmnMS2DcnD66
QIXNBgK03HbQS0dVsMLzTJvsFMc1Vn2ZXnbM4tCox60RpdDBP8epGojMqsZuMsPZ0twOBQpSB2CO
rNZ45rOC2FvwjJ3+HVtqN8m7cpKjA2+WOlMdgOerr8kime9g/73jQih2+cpMGsKWSLvDU25SW3Vu
vNkElQuA7mdZYBT5Z63kE/MDUrHx2lg189kz/0ufCjw2/WrOHqQAf4oTxO1ltkmybbpuTt6qvwqr
iumkUzsUL2tGXUjSJa7/bG5DE7CC+PMwJpC49XwWYO29IQif6jWWBMvHjss5QAwjVfGQVrNB/nXB
foY0Qpbd4zReoJSp0ILATWhR/sZw4/wXv76WfRz3O3wF3bjJSPNi5I4u4B/wnUIEX6IzSC5nFgfV
cBiXIcdcp+MPLzeCBgfiqdPVtGhGXhLyiWB2gpkWpkWFt8jAaI9xVN3D1nd0NJ+D0niIXjth3eJf
a5O2O6Pr/x8nW+RpdPLg/GcnOoQzid+hNzpB/JVFGhUbvpqOxcPypVUA20MO49C/AH8T3pBYeaen
hxgH9CbcoZBz3rL964Dzv1gQK+AEcnrLcbV8vqhlXOIevtFQYqYIPOuimOHRufxMw0XwD3vb7c55
8FJYpWM3sFCjXHXlPJd8fudp6FzFAJJD4zmsCIaRd5WIyLkKOtMAMb1r08vlNQhaoJylrsZMv39d
+WWOQn60m/sPd7cLUKZxir3BONXlscjJ2oNZrQkAPf1St+S+efVu9SpevTEF7Mhs4g3hetZISsO/
WCKq4yC93fim/itaHkRrSV0BoL1JkO1BZotJ7zM87NTOpRq6BEgGLdfX9aTyklObMaCr97nM7GLZ
joHcyZiF3eZX/AOb+pK0KoOctzM7unI6vdLktHn8Oub4qmRtY9DozoYq2V97k7vk26ZWnxonH4eN
evwPUu7VFmJqI1H2k3v00Sakqi09KZF+736KRgmXlG+CD8n9cYQoaFHCdbkV71I5vC5E0CHWkT7T
4qUogh/N46OakbD1OgpyoinUUaHOjVR7n4KQqPajjccSUuvD4csu0+gtACFBjIc0JAf69rIfXqHr
sft2RmQqzpNJ+u3G/ZtXRzUC/9BdEIcbxLQdt+SREYwlXXUqdNYIv5ezdEUSo/DvFsL9sFwJOa3l
C1AkGNgoloaDqC8iqcrLjNPpfcVhP3mt96EY/QAPQTw6J5ZD2XqZXnG2TypltXcbLYzcPbyzdBLd
wZOnXjv3wxG8JBjND5dyS6FD2v2mU2Nq84Pwk98S4IZq+7RN/WPd4vjc2OR8qn8VqHA5ehB56ay/
j7TFHAxWHr5YExU4wifeoJUbFnKSVLVaMslhNdZkavPyuclUl84upLoh2aM4EoY45C1U6pw5q7Kz
xFtATE1V+7c4iR4o7aXmwVSHHRKHgzmFa/OkjlZntdHphOINqCOtc5Q/mK7nBunI8bjI1lmQ4P+J
9jTIjnmtKJ0QVXz577eUkjD0B8infJ2lCH0JmBW7htPSB6z2r81BYGeEIFJUH0db7dYL7dnDSero
ZPeXapyI7LNSWr4LR/mUpElf8eVmH/bPDrZ4pSiaNDvV5sLB0BAIrCctIvig5tO45+AzL8qlqWap
8tKojpJSECLzB31i+v2mRS2/7ZLLJypQAOP5kz5TBJ1DdGd+H+7udLRvNXMbocuTKPAiyKXJ/c6c
Lb4oxqXDHNDokn9u389jhtH8n/nWUjP//ce6rH+kh2IaD5EYqSj6UGOsRCIh9Wl/uCwHn3NyN3bq
d/j77owzNm2ficF8DytWkWwYR2iz6wVFwbf9vq1dIkf8IQMBWBtPUHo1ug1ADIex3CJJ/3nv/fo8
XYXMN/6kJuB27vNbtJqmOxl5wr6uqUD+oNIm2C+FSnHqxEvadAD6P46qRRxSNJEJeFJwitc13PkR
O1MJL4mpnhEotF8itg8rgtzDtml3GrfgMDzxd9B/n3STH7REAIpwYi31EDyqnTazWmkYeV3qybqe
DDmnWBSS7RrF19Gm9xxVs2PHL9DBDBivStg/o/jAcJOs1k3tA1JT6Fju4CYnnqA6Q8V5QVTiiiE+
FleaF6f8FDHOogEGQsqWoNC8ChxF60aLMh+hcWBbRyzcvEIpu9fEfHhERbKQmFDlMympbIwG+OJB
eZAD3fYHyU2JulPXrZ9J1O6oG+v5xICZKQ8iyzSs0QQyLkq7l7Sfc2nnMWA7DkhgPrEaiRyEZVWU
RnCIa5pimCGGbdrGbfsIZ16/j4UmlCzT3J+ESZJ0d/YwzmCizF6iauGafxnfcKti1moa2WxT/zx4
FzLAwLucqziC352nkeAOX5Bk+gWMwPyHo1YF4+lNQgaN5Z85v/X6bFLTVIJmrXDP7vMyVpTuYPNH
yXMs+Isflvz1vkH4qwRPWRY4nHUjpU+b5me9YmcDixunzpnQ99U1ROeCVUPHaXfXWQq90q07vfxM
j04FPJXdAfRRhbayhAwj2/4zXHD5GN9JnEggFq+BMk3wxXvSw9fcFYoqf1HV2pbf5+3jtQicT89E
iMhnUuVnFEqlTc0O8ilI9YxCN7z2+Tddgbok291A4y3ddStDgJ2XlCqcVDlQ8pf6fnp4+CQMYad6
PWp9MBywe/jwexJEsslnK7/CSFXri+m/efuadL4B96FoJsmp7JvzCOoNB+yqA5U3i7SKc8a5ex5z
ZWHsEzC19Z13U12s4jGgbwVnNEM5JKPmSBDwdnjGCAer0tl6kT6LEZp47+DYQTCLCBpMEmJ3dZ8j
xEsQKG7am1Foksl28UldnYJ3YfiNZL3dRzCF2v25fp31I5jD/L02wfSSZlmtDtHCmf6oQjyCU52f
iPpvgQb1QSRUUzC75tvI1a2Y+25v9Qi8IEINsMPGaUOfbixY12VjHQfQiQyhHdaxnpJPivsaLk4a
otXBsmfWI0Fo05LFP1dCNJJJVfEeVlKZU66qCVJDTDJpVL6yU+R0wif37RA3yznGtX6ToTrQG5Zq
ju+0TT7h3h717kpnogGixMO4ZdcUmE2rkbh9HRVHjQneYd+9n9TkX0YHVzRcxXz6NvvjIOAzVgNG
ATWLmQZ8jwJBCXz6tODf/BGwXcfZkz//NKgchJMqhsuvdaOkjsDDYFa08TmiSGzzLnzuP+LAgIzE
ox1OSw+DPmdK6acz1j8mFtI1SZTuRYNalabu7Qwik/i5Y0o7+femMWPBDlpnbdq54Inm2LD0YebO
6l4OsHlp21YIvGnTYLeDJSVMPBPoGYKjWGY/0folMGEBSJdvkfajzhHsGN1SrXFWfl62iJpPBZAf
xu7QKqmzb1VIc/5RKJZLRkSKmsGCPhOgl15S5tJFCVbHVTl9Djmc7q674VhGD/twaa8S8fEZpEcB
enRrH7HJsSRh2IOtGTcRjI43XMu3gE/zYm1GD16iJjCqdkc5pkfVTYhnndnVbjOAtDgvRxtAWA1J
Jj737RkI9d3TJ6v4hP846W2tXrfWvlWtyWIwosJfxLQk6BY0EBrYK+Wc3uKRVqrSvzu+JCmSUejk
l9h26RPw3QliloBSn1OYssO6rKZT+v6vqmGLLqNkzkfXGSz/NWu41tUSd+HYt10gTW3GqfSoeMYO
BkfzdQ42tLp92A3ecLNGJwQELtUEQuYpDhq7cq3KZtTZQ4lKJYRnLJgUVJYZOsK7m7BkRnj/MQ97
L9Wha5C1lFaUCeY2LkhiZCrChTNGmXVbU8L964wc3883M0dmcwpa6mSBU2/FPOvLPfbg29AV5HCj
7wOfvljT1IV5ifCGV/pIiRVdPBZUvSGGtTsVdusROQfIvBIsaF4TJLdrLK7nB1yWLYOw74O1V7Y6
VFsOClQXMEhYhBIwMGHVfbCosN4JMds1kRC7zLM4bxQQJ3+518/QQIxY4Put1hGAKlnCh19iQEj3
0CWmmAtS9uVjbjaNsCceHr2X0Ed2xtS8bybIzm8l9u7fWYt3p5xQZMwz3LhUGFpAF3pG5zxV1QO+
RaS1Trzr77BxmYMBeYFMpfwymcZlZiXtpWF+rxCRJ7n8441f+hnkQge9q3qVXs3gPeR6eCDWcO0j
enOxyrSrgZ1lhC9z38K8RYnRfw/lkaK0XpOLYwZVaWOv5/RJln5LjbbOsE18ounHBi3Zdh7yzkuz
8HPhKmbcDliZakt9DjvkkBkTBOAKk8XJOQBLF7Eqm7y4qFtmedGb+mqrb4iZVoCsa1AGEiF++LcP
PDi1PPhBlkwY7YxBP69wJCBp8zTQEJHDgD7Uk9sCSkedHAIwUDIUXXXEUWoWUnpD4+b2efjO9Rxq
XPqvmSl2/mSMubdM6e/QjsTPXCL111JmhpPe+TJHC5u+kfOKP7Y87/4xciK0X9AD+qVm+Q9jjcbP
yjFrEk6MprE1/TkCQTkUltiUY/pZwCtqrVH1JvRj9QZjvNgFJooh6JUmeBQepuXKPFzCUNHDDJIa
rn3bhtnh13wXidUsqlVBkwczaFmjyTV98LnhjY2qZmzGNfFeqtpfsOwBCGP0H1J4ZfmajefNnK6I
F5AB5jZyD6OIxVpnyHwkevYlrPn92pz/Q/KRLbWaky38eLsgV9Ov8t1yd1MkmGCTGm7tW5l2oojj
dQc/F6LRpzCXTPQmPuEiB79hnWil5k3sWm7X5ihLRL2HmqSDyFNK8qDI2xqlroRfqmiE4/4AGG96
z8stHgUFezhQlR83zemxbtKqQGvZLFGnaUdFSw9QtdmH1iTERQT9fVGWj41u4AJhOW3ELL5+PFpt
uK2WBwNkrOdiqMf8yI8tJM1d/cMSf0+a+lVEYjUblEpH/5ASeVfxZlhOZ3VeRJNUhZUbDReFBTxn
x2ncIeLD45p5H1uuI6t2LzypIpTbmspJh1jiv/XcxwO02veCysr9EzKvTflMd0Vz7UkD+K0kdAi4
EFjpKNxnIxeeoNthGFF0WMLd9K8VQY4QwW7iD5195X/3Ny0v+r19rY+XUk/Wufuj4NxcJvCu8gIL
FL8jAEYQ2NzsObsCuQCpdqow64AIU3BPx4bYxInyOVzh35RG/tmj6C4QTLSv0l30o9AgO+SSlBg5
mM/5+mx5G2ZRt3y8f97myolA4lGR0SO48G62yCGuv/zbjTWhsPHAPAVMCARkMQ1/MlAFQoeE8/Tq
BVZ0j+AKW5CvpkwvrZtPArz7kwwYoMOgMSoeo8k4DIrNnN5eNYvce1aDpuRPhNDMlOOmzy70F2AQ
1EmIb9KDK6OnKQQ/Jr+lLUg8vp1iDiuU4AdoX5ea5IuXu1qP+kV0cBVoLQIDet6lAMmXpWUdyWmZ
G+ViGdf9cxx95KlUlDyFxhfJ0ONrXhIuiAPoOKQuKRMlTFkvgPKCSG5twwkd9WBsggjoHcXy5oQA
HN9zi170IGVcJw2QF45Qu9lqnjy7X66Vbo/NmpzGxlzRx3Dlvw1LwRtOTSQOyxwkQHK7oHbkPEiY
auw9A25UXbSvZV2MFNYaEFutilADC1wNr4sRmNYm4eD4J4pay9XQWzycK0FZGNc+ljvmEZefFlwk
Xe+4EwS22gXir0beGvYmeruCS7fS6wV+NDvpjvDdNZ9D7oiMHS2m+tBRlFvQG+3g+dmfwyATGMsN
Ab66dlziXcgYZEMiiqkea790NoVYjdvWDo1bWd+WHsGXMKtFqVaXtwPI1r/Q1HTx264BgScvFUiP
fBJ9UxtEsl77ZneVNSvRjyy0oad/Xvo294Y36gM0QIR6GLA8XIyuKeW0zXY2u7+hDhVcQV0ttjbb
d+aBQ5KZHH/MWrSQJ0lHJ7nDU2FO8KT3rE5Q2T5pWZMgN0h8qpIe7ykbg82+9m2zKWuLzJrOfJ18
JWq7PXtthL6yej3n9GTRKFb+cxCVW8R1Q+HmEDfIC2jshPV+1edFstrldK94ss9hrbSe+a3MNV3Z
fmOEduOVVeQyvRKF3ToboCpMk7OabY4uria5FhOwW0CsHmXU7rIPcyQ/QmZS09nE8iBTL0sILgM9
VimMZWNXKlZorB3syuaq01IjunWOFwB8ZROZlB2hAvJKZKHEZNeDxjUnP/M9T4UmbVZlxuhOf5Ep
3kywQ63BPquSLO6kO5J2xEfYZ843TTtj4bBQkm4uz0ZRE1oab2klDDE0EB2imcgXo+giG2PBQ2XN
/oXa32u32cieSXQYlacQSnikYleGmK0JSFSrPL0YMq5L3P3zNekzuCa1ZByax6R+bhsPEiCsX+gI
r5q1BUXGIpL3XQ/2zIjzMsAbXIb8m7g8Ne+NektlXYw8S551PmRFfMlC4lUfX8BEQvSPg82LEExg
6pyfoVOqxIEc5kpNChy5vmBGtbcpOuWMc7JzI0oD4eeRpGTMrntRNrXHd3gWdQXO29XRx8gfVL5e
D0qt8JJsKi04/WtaeJYp/eFhbqKPhpB2YCjrvju8fbq7nMmq8l2zqhUW8lvgQXb6iUVoS1eA8qFm
zbfQXX1U/ljt5pfHArCja7pjybSziSTuF7t/e2KFUOcSUXlReQtkEetFBvFdPidRd2AaoJQzlLLZ
RMECWvMixrxBJkTfFAMceHM5IQdPMUhAewo+DpvkFkOlKdcZSQ4nECFsU68oPN7dW8skw9omKx46
Kp1sCacEvVgXTHq4fWWzdfaNlPY4HZnjdFIayv6gfiDxQxPHLmG5E6DiA7P2pfoqH6sSMXHfgYOT
tmamZoRV+77NTe0DUs19uq18bPjqrn5d3y7mTnbAvUOZK6N/dwjlOtvfpLyYYkt/fnz8/pdTvsWg
i8ufUQmVqGFXjmLv3oDR6M5Uqn2rv7EtnXnMlGWdH9jeOm6D0MW9D8L+PQ6agTfg5xo9P0j6iUUH
pDQx1D7MVowwqTj5GAlXBXRB56d7Y8HBqo5SV6Oiur1GED/Cne9zk16mRV8GNOqkV+OT/+RiQ1AE
GP+3usFkUjctrmORDUarnyEGLTfBt/poSpgT6rs2pMm3w4uUaJPjBXK3dpmNJ9LZ2Fk69XZtx/F2
lsPpkQ6yShjwT+aiOXHMRLLzdvLLgil/IGgv+zDP13S94TR3zhIi4czm8yUzTmSma8LgHB5A6s1g
gV9EJcgsRXLBhoNl/mXKYh9iYr8diDD/G8oShfa4GS+S+aA8By5IP9Ag54/MVLm0kkiOoS4Ged/u
9okMAN3WBdSHLpaO8hMsVzmiWZt/FAV6Gfcobvw9ewYSYeNF5Y4yX8d0FaY5Rpym0cjzIm6yQ1Wa
Hm30gUhbgjziRduJ8TkuxP/TqkMMyGS6hKy5b0strev39qPzqmTLZkl7vWDk0yZirwasoXDT/t/d
V0vJHW8WqZ7cgKFT6THWUWFHcSsiMg0Xi4MTvwW8X3ATt+P59DnOgNoP0Pvl1QYx6zK/i/h+viuU
nT+tsb6ZU2yW2v71mut1SQA9AqegwqUbvocxObKbdhZIRTxPgxRp1kzmKPfoBGLlShBQPzw/HHAo
5rottbqoRseC+G4/vuC5xIlAwfFLy9TNkI5wZqD7xa+ECn9svUr5BzhLwRgI9j+V/5uUuLJeDRVR
LVTLZ2TIw5ECL5X2dh2o1ykrfnJhYwxKBZ4zuncADBE2S2gG+ptHe3xgSgs4/cuDQipCP3OySv25
mILBEx6bqDWbV8TYfCRhDeEF/iQKldsf58Buse8wOWIf4fCG/+3MRfkbqJpfmi45tP4M+eNB5skM
wjeBNgEZv9HMq5QJRgBxCRIgMTSDVSkqtdOjIlec8znlm8NV1l6hs+3MufztMzlQ947UkJjoxhd1
grKHxcvA2WUCWpJPAaBicFaDhK/dpkMXDqgeYPT8yCD1SsY4RBiqbdx13fcQf96DacanclgmnIFA
PchofbxZtH3iCllxEbgps9mJgdSGvscuuN14aOS3E7vetqy5xSg1CdGWX+blhCIzheknefXGIm5U
n68H13CP4sK6SoT5z3MMcusNtk0m4Q15eRzX6TzU+Zc+hUjrK7ZuIn4NZQxNdonFHT6bq6+wA10S
rClfEGae1aHnL41az2NVswkGYtrce4LlmzeNiiRRH6NU1bEdf0Bv+NGnc6ooz6NNSv4UfuwiX4TI
N7iR1ej/WhcxICndl8m0/Qfs0SjzPFBz/QvaJt/IdM5Ywzz7XSZksJn+bF5u5/4+1uXEn4liM1VO
dsBG6gz0bCaQCeAHhs+l4WjRgi6xtxpEVTOpsVW6kLLjdh6R6TtF1Ds26YpvX8nrhE+DCXlOQUR+
GbQ6Q03eKh0fKkZKQ/a0EuN9nFTCWoQUZMgZFV18F9lAGhIFaT37xkJM44UPabmXU4vxvdpIXoS0
+UB+9dQ2lqZ84AsQIsC6wyorgjjsgaCrIMPBGfWDtvCaOAZzJ9hLuNoNgFBJXmv25zUhjiGNeb3h
MNb82VAKhDa456GsLgfRfQzaXups7qWBnhqoWJDX0VqKPJyXz7Ykq5ZSOlotMEHB168CUdEXBAqS
BWqiErtoMtw+5RJUANs4ubvnZgYbrZ+pCCM+I/sck8mguD5BM2y6PQqmamDpVQ9XQ1VbEbYN+NBy
8TvjHv0HT/32iJBIKahkWCQzu7HVbbMGL8CGbgWDyJM3L5v+Fm/BSt9TgBkBMg7rh/LqGviDTrYv
MNPX9uxxotMlvCCqtQghoEqpEuo5R9VhX/rIbBo/xL9eH6lojqvfaRb9zxBkl9xBRdxHGeliriUV
A5A7yKv0QhZ8cMZQ7wfZOLAv/jZe2yVscrw9YpSQhaTToVIqt5Jd1pJ+JG2dpcD0EtUx8XmARPVT
gRDlRrKW4u9egxkDgGSMr6iaFBlfXsThK3fSNha7UVNZ2wvk6plgl2KcyT1dZu8MJ36E9uzEeron
bsjQpv4dKWuy4/KVGOlKh3MHXm/5p8QQ9X+npCdZ94btFygXHyWAEHFZ/YpWnR83U63De6auMvdL
ja9fk3Y/ErwZnL2GuTVc3v3rYuN+IIfG9w6w/KlFy1mDY00B/lGusgpg/KPFeRb/KMR4QF+we+PL
SepPa70PL6garMAPRuri6fqmhyBVgzXdRl0r9HCUAGbbDLJeLipT5kHr/12xZxK4XkhNEZDXBXyE
ykSgslrGzaIIaWTQJbGGFtroSyBcxpVhEaRSfNTNdw4EWn9SeGY78/hmdSy/aTHLHMUF1bUvL5JX
sk3P2K2f8mvBY6qQXZk78w8QhNI5Lm8B2lHFUcc5lO/X6TmzChmcJT0hCUlSkBjVvnUpyBlAtc4z
olx4yDtF2zbVhe6VCqQ6gwtwgxqItnSHOdXApdop4q2sFvfGSupnBycbfWDtgZykhue3OzZACv4y
NXybMDaYXifjeGU8lr60OPR5EdSR/ag/zdgLgTkTjRWji922u4LbAy0k9PjMBoRQ6+clhNaMsDSk
6R0/Qeyga/KdgD19qyQVI+yZA8WfVtU0sAMfKaTVjz4OkyiOkgVn8qu8pffMrWDAD9BUB2/b/BkI
lYKzN1oyrIoMmyJukRklXBEerIIMEYnGBclBXgQyGYmswTss8A5lOKsZmJ1tZTL4voRz+/Ye7I7+
IGSX0cCA5ERkkO2ytorTWbPspDg1j0jyVUX4XwP9fzmzwiQAnvSzQYap25KcerqYcHkvQvnelItQ
XLKbCWVaQQTWLl/8kr58TFCyymelg10qS8F8/jj5uqV0Y2oDd9ZE3CKV93ZCSO059NfU7olgJiHb
MOXGAiB7Nw9CpUdjbtpCNqv/OUTL/LDzlrZs3zyG5xciHFdWcSvPwcJ5g4wVk2AFYHjMelrekeuE
TGNs9FlZo/GPOOvwnTgfZFaNe+Ec9F0k4pmh22gDj+j9faU6/qJegRYdN29cVh2KDN03jaB2J+N0
idjl4YXISpgrS2oW7n8NMhZMK8dchaQp7pSmB0W0gCB59+XO6ex03C/KRHVeGg3Xr4MP+HoXaeeA
S++h5oyszJa+o3caAhMqeCVIkMYFVhBaHuelY8h409OIsr8gEZanndPYhN6rBKjaVOIXtNqvWKkk
LV15YbMCQjhfFxcNmdwrAa8kyXQv1EB/4wXrYHdfGAn6ctUDSxHkNkig04kxJU/D1EtXnO/C77wj
6LKbC3NyDTG7z2waqIOhlzhOI5/38uBVENgtY7PUOh3pruJQEbSC3QBNUPlfm7qfh0kNOxBUPEeA
NXQqMegMTklWzcNnP/+G7jd7e1hMCO/2mdIIDZjuwQb/01E6emxXNeLC48NRQFinQjRFDlw0uVse
K5c8AgYIGT16J92wQ8isgwVoUxOpmlqgoFv1GoEz+lwhYMC9cCdODc8fdIeAh+tixOwSwUs9ukXI
tmDhYpH3B5S+xh5IL9XDLOLA+LasM8xa4WP6X1u1CJuVMjoG0ePNeHbBh5gefhQRyslVvugpSOuq
U4iy93SCjuVqfYoAodyhvwzHt9trE/1Wo0Id6wWhpCBmEp258spqubhpqwWZORDJM8DbyCRG0SH0
iZWg1N01wjpmVWmyTH/Q5KGZUnOYSkiVnw3GPMsm5io1RmSklGD1QKymREgjlDjhPm/2ytD18Psa
QRFYLhSYUzRKPhyDfICAqR7J6k7Hc8Bg3UqWE1LutzlkMqfT+xwdBcSXUue4Wrmbz1MwrvPQ+j8/
Vo6CUeF9OTUDsRYgxE4nEbJsu+Ta18FiXLVl91uizOe7QmcoWkyHiLe0TAH8RFkGv5A4SMSgzXZB
2XnAQqSS7ujv9WC4TqTqWJCltNtjq1ywppU8OoUoqc5c4noqqhkDE5IZpMYLe3S8W1HjNSvoQUlw
6uGJ5iR9LR4zEH+kcJFLHV/hOa/OGZzJx006Rj2nqTk0dwCt8e23qHJjIcVByiwArXLTODP0oX6O
9wnvyD8aRNfF7kBJVCiU/c8aarxCI4Pt8+qKCnQbsE+6Rjv7j3DGcqwBHWpkQ71heftYVri/a/5h
tWUgdxFszwu6Yjy07Cv3Rjg9+NqC4e52TINZqJ8eQPKuO7P7bM0eFWwi1kaNI8dLihw6rveBrmGW
HlbgWLOOZR3A4YGFs0PbYaQ0ePvZ6Qjnpgs8jaYmdKX1rAXcyPnL71fM226BghBH081pMpJrdQnL
S8U+pb5ZunuTGOC5vuHaRD9xCOxY8POX/gL1/lCY1S5C88micut5XgMVvwre9pXW1lZYhySoOQMx
zmBwZPkFjTZn36iy0CQvv8LkDoN4sGjLyZrs3IdK4P6oFKqDWTUKbF0hpQbVUITKaJxzpXc1ktdr
zmWK/SzuqdmWi+kFuRqoe8ccIvLuabO4y13hwHMcsUEsjnfMDWDjEreRf1U1gOXR1ozM1ZhOYp8Y
rZtJ2I72TQb3/r4LlV8X5zwAknxVyq5fMUgQG5Z9f8gRt/f1r3ql5ET/mZgBvG9fwKOMAdNbdVu2
YGJe3aas4uvD0PH0ZRrEJZhWjlhPRa0fp7XLkUlBoldhi4nXVblIN/qUoHvCvwQy0lQIsr8ktTlp
UdGx4MtBxWKOLHbx6u1J67RnQwA5khtavbGY092/me1boXf+IShcezAUzD5IxTK3lFbJPsgU006O
Eh8YMT8pFfydozv1cx192QgTbPOp2UYdH5DkC2TMs2NlUpll9EgnPR30cO2yt5hWpUNrOhsIXIEO
PVnn3jsJaHlN8HyNV7zqZbkGtEWsAUOo3lkYxC2cG0Pj49twcxbUmmNe5b8H9amU8JSFcKG2+tkc
Q6mgfmlzurN9jLn3WKF0LXIbI1LWGlrpcCUaGQHFyIIxnOqApJT+nEu3G/PwjvIOj6R7v2KnYDy3
LOzafku/qSpY1wqJvNCXg6aHHmxYn+gHsKVDckp3y15mNVJBajObUL4TFw0lD0YWotkYw+SuSeyc
niOQn3LRbjhJCyC8FIjo9QO9zZ0tcDMObZl+R5+LM2ycobji0V7Sic4rsOOMfTMDg/gsDBgysLRS
lcqzfuEtP/4Hepqop5Jy1CUeSKUn5IjQCrGUypjGD1MtrQV04yrI0M3iy7bQqZRRT+d/pC53E8ww
p6zZ+eeXMLjVhGwbiWnzkdWslermHhhCwFqSJJmJLw3Sn45HTdPvySGUwl3pgz/R8mbYJv2O/yuu
1Vg0MzrrG5c/cCnUo/VEHAR2JMnBHwsc9Awaxk9fJziBT8nbL8Z+r+k0nENb6lDwigNHO1o3WCGt
2GfuPQN7RKANGcLw+JQ+rk/fz2txUov8It90oXUh05apSq6bjPia2w53k+NDWaCo06sL0sYSCIs5
8tvwajXwN7nX0/9dFp+20BJlQ7gktbXhDfoW5dCYDHzw1NcEesBJONCSoqAO1xuqC/Ukfj6TbcfB
pP71y9e1ol1IHIc8VntSSSmYp/APKoDTcqHq+CZCYdzPfPGfoM1Gf6wDbbSmLFuclI/hNSDdWeCW
9Om2IJSNi+8aNsNRFLpXRUl6S+qRT51lCnvAVaq63AYbUPrwLhWei+3QN5oJ7hC6b9b5pYfcoT+X
uQuYUrOYe2PuLTq2QgiHDqS31eA8yDXfKF1TXwWSXyEuxzR/cp98TBjMq/7XhMfzbBDUO5UEDadb
fwGrJfmcqve368Ajs8aTAySZb59qwIyPw8eebEcgWFC50XUHOPZRsBCcqAEMAd5iIs25Rd9l2fee
YBDdxvddRFroth0+dtVVbWZpbke++6vSDb2z2UpkY90BtpxxOsb5rZTjf+hWm3PistH4qwGQBEEM
PfTUS9YlitVD4/GuAVOE4EgaSd9edEPwLr5y4xpHMjqmX6+wUvFoRrCOHSFEff5L7yeo1wmX4iDH
iQOrarTRYthdcMthXVyXiUQYgwMcshA8NxWI6I2gzsy/BpaS/ffhevf/cD7SM60g2oCmLB9k9OKp
Vf4+9WDKr75PMpqqw0fEBAeFrhPNWY04y4DCd9/txdOcVopLT+olMlQ2rO4vF0b0/sOKUIFvngBD
8hej4fO9agQni9WVPfAlit52BbxtrLwz6dInpA6sy4uxm7zYbSr/7nO6GRwLDL+xe8IMRPEWz9eC
e2ubWBmXCnzEKPlLFpHnFLOH/ynGCN/feyXvkPopCaQIHdFaPz/rMfsjvdMtJYlhIJdWeXUn//yi
PgBCH0u/QzKpS7vGGBWbrcbLhFm/xHkC6lUtZZZvKDdMmFEz4rrZM8W6x3BqqFq1JdAZy5gaxFa+
JYawUnhl699d/f5KbcQA1FM6UrTlgVCtkoml1SK+apjc+ZOvEhBKhM8wFJkKaKAwJ01XIOD07onk
aZn9GPqlMySoDAXdaOgR5R5GCVJ59qheirxAMdI7ll9LH/4IvYROo2tct9YTSIMgagMnYKEUj+ns
Zx2YxEtccZ7il2vGohJRjAl5g523LqjQNzzIKK0S7a1qI+QafZ9qX7sWM1AEbAQPyv4z0EJdij2J
gTbhMuS1BoNBnqtdr64PHCcErLnLBlCkECxUtUkwZKtiE+koeDVdvTdgr/Zl2KAUX/LPaxqrZc2f
vnIPvKr83xOFRE0FqCNl6/vTMuanYjgWsxRV5t5q375jEN6rynqANd4wYmkqblMlA2fQ2bzzK9F0
PDuDeMQ8VJC/Tzdx6ytu122sBC1iLMH5KU/CRPzy2dWDJgV5abIH/Ypw4gmG2/S1dEGvBHA6nVLS
A0ie966j37NX9vl8nwuaqy6gC25G3iNB5w6LzkmE0MQ42rnJuZhoCrZPjAPHX2ryZXoiivluxECS
OEhZXnjUkYHd9Q8iH2dAjWYbHdUxWb92q6zvq4CQllqdmJMGFr0mlF+TfHmFo86fOJPUqzi/yL9w
rIvHUuQVor3XLKKnX5j/lVYclk0PTAxVfehwv5ModaR6zTFcPK1FPgGPUk/Xojh623lUFYEFVLLb
FnE6Y3WfbYX+0gE2YWDJtj4wMxsZheaf5IrkMUfNXR+c+udm0ovP6PU9SAzACB4VUmRuNK2wozZs
LuwLy/YB1PlbReV1paHB0R1ln6UYtYQyNdU9aajkMcuGx0IBFwUC0VAj9jI/j7T09WGyUSZgKlZd
9dWgZsBOL4t/bjmD5zcUxXWpKNNcHnudp/WI9wmVtpZkRrI9wofZBYu23B8dlr3DvpDEKJFbc98Z
s8FmIXIByFpPisi6QEq9blX0WjlqFPRFrBHLqx0PajFoySeK7Cfvj9Ng7BrIdO6OyS6lAyhl/u1G
vfLlukOxdZ9XLF6NJtT/Om5j71niJIX701bpnySsfqzKXbNSDOk3/Yi8t/lvS1TBL8i0CkFqB7PT
2RthmTa3aTTtfNxhmZLbcrSt4cKkNxLOK99hFK6l6wybx2qPTNwLikfUA81egNBnhlvIJFj2patP
PAh6BvhEs+E0VeRv237IvhxgQhqXWgDwIitUIOTCnethwuDcFCkcMO1XoL4IYPXm4nfcTjOBAvI8
1hylVNMFKT1w41zmV3nIkzQb5Mdm2efWYaakRheSlnPtpD8gSeCQvxj+vRDNP/h84kCJ96n1+SQu
ry0H2xzGgUOmbcGsMxKJBQAAsMsx7fX3mQ6XJ2lshX9PbFziOhNbHTVTtwtTjjDZn665cIA+iQaM
SMZZuQ6Ep0khYpjgtIqxeD4xU+kNuJ+EdlxTTatk7cOot11JIFrOCK1lpFSPSjI82tiWfXeuke4X
AWat9nSqTUGp00fJkvXUmVe69kbHEm1MhwsTI0Un7okmWPi1rns4bkt12R/KKfesbEdLOK9y7IHt
WkeXtkvf908vo2vWiMnB1h+KpiqGoHBgzYv72+eiHTM1MGPRVeSR2TKqBXHecZ8Fze1SE7/G2b1J
h+KJOOPr7/eX+LVADlwFuuHsuFcVYYjKJ2u5a7yo7opJ4MTSNpYG/UFVM5vczNhrL8K/45exoaIw
YL7lYLYSlxtQNbOEjisDspzkdJ7AK17ppH+2lk5hy/VfHakIvYcq5/p1zpwyeEKoDh4VXJBEWE4X
7roxv4NZZe3t2HAPPd6yUftUaKt79/LKstAkouMlUEdpvpAXK4+7J31jzwK9rFTrVu4W+QcLzm1k
IU6nxsMxofuuGyy/aqOsrzcalF5OUjN95AI4gCxwiW/LC3bQvbamUDXMvPm25xcfN70BB1jNfFs6
OqSf4Fl6KAVs3wUiz4BseASc8rKYWiN3GP58Efb55jSb2KvaTyQhtZUAVlne0nklOSbo+g5AbVCO
nZpempKXrDuxjuzsOTqsHpQgSBQahqT3pWhyR1TkSS9/6skH8okhOfuOYaXQokfk3nb84foWh8EK
YZoCsgOSnFN+ekr+zIyla+S7umzwfK3HMUPCbHrTnBDq8rL3rh8rNvd7xlhoqDx4y99vcPuH+K+u
mymeGvyOpJYMQjaLkym0oSbBXgHr1zLLkaUERX/soUDWFaa7C1J8BrmB0a6+KaRMxZ9B4NCxtefj
cXYDaGAEDS6/OFYbmbWxFfMhPh1noUk5pJoIKO7zo79Ha10E1bUaRZYRZCnR7eLR67Gob11TkcBR
M0uZsIXLdVt3N8ip/nxtULYVOG6eRPZzd5/1rnPwLEl6WHRO+XSb0ABLGI2PNw0kOd7zjmdY5vBG
4DQeTqwCoQ1SIHy2wU4uvih8pBqWvLEm7ttJOYwlUvLWzvG/wzMfr0EGnGJ4SFeqO2CTGNYLKDBy
r1BGogJuP6z8irJ4kQTGJc5AfV7TjgAY0IKJu3NSUs7GvgYevUCMdO6GgQ347VzMDK7++tSTpz3E
MTUiRFkbLsy8YQuJmgLLLw9toGV+60EZj6OfZuVAmeczTReVxdcgCq83AAffMurdH1coOh7pI5tq
C2oj3dEK5ub4Kqfgu4QzFTV6NL/QgV1nAA3Mo1loUrlQllJF4SsuX7UnZ77AiC+pBfCbi5Paecv1
Tq/pKGhR6ZMhkQG9jiBrt/SHHdgDGz26FdFa7XPBCUegBjdccjj57lJ8xnAD/5sf8LWq7LiiWOCl
0aaUSHHU9IHHprBdhpe1zBsEeR+20Jn4nnl0tSDlzH3/mjBOyVPAqXojSrVw4IZvHDZKfj1n0qcg
K456iFgsKW1cnrbdqXFD2D7uU/jSsgRvFcChNjY4lgjsRdZORL9kuLoI+aTNYRY0Ra7wvrnNB0cW
6vZSvrw2LuaTczXizQUsodQCJVlXmhd3+pShtX30/Oawve9QM7KWX3tS3RKj52B29Ncw4UCJGIHb
92VYbqY+dqhUa/TXt9wS0WZ7RDjdtBLpoLl94bQ0jOwKeUBe0G8ru8AeYmUxOv1neXhrNvSiYSYD
mpSfi+S07o6bwp3GG34YROlB+O9W6j2KrrCbTnIz/IPNTnL5LCQ+HZ9/zRj7WGy4j5DJvLrxI3qT
AokX6zKQNpMkSrMyTCHuSXnIeLhIGCEfNQxh681edAzMRG3m8LMR3S7deCrRCl1e/fgzT0nwGVaR
t8KD2IoRwNt+oqyD72CMJ+9YtY3XfLgBanMTGN4/4PM1sRIUKV3LWuqdYSm28a34ArgS1EnPV2PS
mnP9yUEbFo1NoWSoUeq7XNKRInJa2ZJmzAqFZZXLmp0PE98ahINFiim5YRcG9QTIM9EJtqGDn65d
V1y6B7L/62/4G0GM/gid7E0yr8MxA8R2mMYnvNg0xyk2KJXzfllxMWWvecIoYFOFtTZ6O4LA6G1k
Dz6b5/xumdGREH+NkTdC5t6tGtxnaCAe6+sjp4efDyoMuMqXNT5D5r+D9NDYN8/ajqovrm7Iay5f
n9KfynDZFVlIm0MBJEN12gkgJOboWXO5PKLHBlxCa16ITsV7F7ETqdkIbGpMwL1WWzaEm5Ek0cdf
e6Hkj7Aj3VVBi2eU2s9h9ZlEq6vHWUVDUE8w3NKOjHmEGBFAaYiB4s0p138OXZQJYBmsPxl2iLi0
rPix/hNK6Sz358WL/c08GW2iw1pZOZ3ZK07g/21Y7abDuqp+br0X0L7r9vnSbEBRbp+QSmwg3l7c
1pALseMF8dlSIT4/1APPPimtctVwCxO4DmY/7rr0kPYYwZQh281v+ejfgs5zQpHQrEmkOILWZ8xY
WjD5fZgh6taHtGTb+uS8mJfeBKYdoqUKGJq7LfWWFjmCfFDya3qwdXklo7hFKn6+1bWVXEZ9PeLH
u7ecHsznyoD7jAlk7sYy6aB/408oHSzwKetmUA/qkH2OFXeaLda4zxCmvF5E3RPNP/9wN+hybr/S
1dIcYvTTg0SV+qPnNF5RQBl+wQ7xbzcLypfcaSkx/tdkx1Kb44xiHyV/ckCR7lG01c5TbJnKMLci
nNbcg/v6Af4H07roLrLR+wVqvxZ/DYZq9rLsrAsfHei2N/nAm6PxRWXc2z8XbgKCWTR53ZLD2yEL
CR3EyEnRHxC+6Fgzp02mKbAo4v6+v9DA2P+G9gMmMxOql2JahbDjm9PaT8oLS2zPWDYo2w3CRMuc
uF0Uth/sxdXdOIXqpeTl62UJsFEbYXPxhvqFWsmQ3zB1hKu5mBqRojydxZ4tJ2ZKRYOlJZRx9+A+
8mgMi9/ljXpVwP5VV09hpnsg4tFoZNWFGrOvK6z+8yjeBfi1Mwl6Pp+ZnQk3eSdVzJwJKiNBRob7
YzYen+GYF8XT68L3Yds55Y9AAF7EDaJiXkfmkWpguI5pe0cP29iVt14B64zjJAbciaMXAeTx2uOx
U4Yb6Kke2sYr/QyFv/mFyWEN/XVMpcV+b/CWeMXZDZxm5s6RsPPBbK0KQJIEUtZqfFdf5H8Wj4C6
eyRaNcC7ZXLmAcHhAkfho7xj9FvPx4H/geVvBSdPh543rdduU3NGvuKQ+G0G58VsDGn2g/IzZtDu
SMrX0ugc6gin3bp3FLlAj2PcWsn/em0wvO+sA+cpvM3QsYooxgleFxrF+NLGEt9oOhcEPahyLoqx
OjEvAU3BmFs4nvi7mup+d6IL7dbc5xND1y88cjniCgpzcb4gCRkuMRHTXeDB7E7UTT1asTQ1FMla
+TeVSGqViO6whTs7CPjvT+n3IPFwCijru1sgNN8ddKgI9Lxc32qSI3UITe7nrAABuvZxJdvX41Jf
hX+W1M7lK8rbRgb3C5UE/kzFOG8stewkXKXvXC7Qfq//Bo262h+qUG33DfarcEGgtA64s0bk/FN1
E0LtmFCrbPw9rsTzHNtK3Mjo8l0Uj9XMvk1Pvfk8DIiRIDaeI+9+mxTHsApA+jGkISeK0AUcM04L
GY1G9FokdNyoccIL0RRhbko5eCiAA/4UW/Bxx7YFFrFL13uAVpFsoG5zHOIiJD/SInYn2y+ROakj
262qrEWfuut2YVhVq1LjvR1l4QVS1Oi7t9LTMwOYEMTiYt95uILerXli5aRlzJOyXggbjyxn/2vq
DPEm2gU0Rwuk1faGOiQMHfqAhlPMDYNB6F9l5sGSYMdQeJTaFhobdWLGPxNwGdDesjSj7Y/MstQc
idebZoz1NCPqkNo+CvqhEHlVp74K32oB+mhwB+1zbOJ0DW3GkUzs5eVO1dpDvJ7XS8N0J4xRYh4O
YKStCkWo5l41tStlLSomz07r/LAwD1AlikMoVJ6cjPodemyJvV7SLbfrkgS6eCKtAeUhfMLJing9
l5gONj3oZKayQJowaekc5SZWJFssmDIknY+wt6LhhtRQklzFBLzVHkgdUc1I1QeW+AVZfqnnRvri
4o/oybb6zGaaX80egtg6u9WWBMhMBd6H8kp4pnet/yMXGkIBCGgF/PaX2Ka11uJtKF4nVBeZYMPN
ZUmAF0kphllTbLMA85P9kZT28FP3VvstI8AlrTnSdtT1MxZ4UsctOQgsfExiIO/14LakUpGH+hDn
Mvwf1dyCpK0FJYnnVEvT+R3iGN0JvJvogRjtRwlnjw7Hh9MP+EZINxtrjq3smYbdHuC49DwM+yM/
njoOt+moe/CphC3NK/Xj23RPZFFWweywMnysNpT+E1m/Rt7lERu2WYjAZc/XWAv5Yj5Rsw5K97dj
dQiPUtuqXnUZVI4BoUi5B2xWDXomdfi2vI2hvXhn99mzA80hYh+hUbxo150bEoZ4xuy8wlmh8c0E
9Naz3YtOjKxULNnTEZWI/ce8HNVt0dzrQnQd95+gxrHHKBTfkQ53CVIB5WYsx8V3wU4E1emdcS0l
+zUfOedcGPEQgMKIFIOKGGZea1pHi6rvV9VdDBRv2EUDJqEoId3FWfTrEs8YYPsWCLELu3de3WjC
3krlPulMSlSu0UMNg7X6YslTGnQJEBJ7Uu6qfrHcqkDmaPyh1P1ERTZZ83XV+20huCiHtoZW4WDX
y3WGiOk3KN9T5XSHJTQ0deyiKAJPH/6q9TKrrMYaKmwHCly1OSWq3DOmSxChK0RIQ2VDXtwQgjPD
kOHeDc3FK3FVfZJxg7oP2CBqRBwY2vQhXEWOZCkx1gz4bX/vTeFapeTA1hpTpKp0U+ufREDKiQP3
PQ8Fv6b7uaFhzAdT4OP+uM/zaCuQHoLNqgXS1gRkMxc2zg8ZGNA11hInFpcW68KJ659231UGqzOS
YO/OnoHvC8cQUK8n9uamAP2v56KLxURaUB0OjEWfV4kWq9LagROlrDgn4tudsav1PR+BCgndDHw7
4nSmrrx7kQ30y1bT/EiPQlS0GkXnlUNMAQ70Luw8/CB5fEXXUPNO3Tk/9tDENOChwe1Lf2hU1UIN
wiwroAfjYXM6mjeh5xqzyW6M16s2EX7HOlGwRl26zjwrvUQXDKsPz+TUSF3NCX7H0xy59FMGf/bW
bk3CG+wE473rXK6O+tAJmxkGME0RPvwlBlXPPFIHLbuYkYcDBtilBw+D28euS7HMbrbwlX2zqqOr
A7MrSY+bfv2gSeD9cRrpVo0yLSbmKVv5tACvtBH+YXoJ49FaFMB1SiiFrQ82TLrTCuKQ0lZqpWYF
C5rbC76NfwIls2irxrr5TiauLqBtO3kxuMlS9PoBMH5L42EMTDus96SPTCj2Xv7R1cbQk2Li745u
VH0FzJu1PBV3G8h+hWUpw/VvmP1PgFlyxei1NMR9iWBn6ofFoF2c8KgveqnXQPSAwnSMl9IIKu+B
7vZpCdjDpgumsLf2sbsVLdOdKMPdecCBMgO2iqmwRWmYTW1dCBrg/1Lj17wXFGyNaFedJGKwJv7S
pxWqdIiMYblk3gD/6NNOVzYMNcUXI/SCIFyofB2ImTp/x3KFuQuRNbHCVTxrAamZtogxXWQagguO
QlIiIZKUKIkcbnZVg1+J8EzC+iC8CL/LOMO787U4gp9jz1x+d9+z2CmMPhHhfGgB7rfdWOjCdLjc
ZqQAiMU3lW+VENzJ/DF0s8f4meGoQwqPL8FlhiHJScpOMgYu7NkMHW2Zn6BxeyzosiQ4FVymldEs
5ss+02s9meB40YAYjj3GED2/blnhQ7Y3HVaoH/N1/cMG6Y1YWVuzkf85soWm8dVn9DM+R6RfE7fy
ygzYuqKdYc6Y+uhdj3TNac1VdtH+M7nk3q4GqhkmFEKRMm0ocuYJCcrGcI6wE6gbi8cELiSAKhA2
WA0XOYgvbZ96MqY4rLkaTtc+isIXSRQKt3/0ZL7qQOGnpexpSLVQDpCCzUnbf3smEBocvGA0BQmx
sdS/OkWYuOBTnPxnxmbFjde4X959QTBOM7if/V86v5ccYLVOxvXRngiEYR3zWeXWhu6JyxbLC7tQ
xXVIVur6/2J2fqL/7mJI98qBg3KNnSpTj5HvzGzi4OLi4gt8Tj5tutsg37SlLPIcVS+LyWo4jrvw
XqUVCAjrAw963vNgm3xhz3pcGxKFzeDC3pKeaW+Y+0DQVIrteoEVhplfInswcAZensRaqwjm3Fl8
7guU0TkT8/cp/S2RG+8H5gZwux1S2/V7AtEQTCU/9Er6Gjdj3vJp7Ovw0+TA3YJs3XKEdl9p0x10
qa0Ld3F1vDYtteROHuI3cAiGh9TSK6SV28OaEhs0yUYZ0lVyFg/zhSVvqDkNvoghlm7+8H0tWZyt
1xObCTMx49PDWx+zwsKNppwQdWerhgXT0lDnRaPq+pwTlFctG1kAHeO7BnORZMaEF15p9GMC9o94
1lL0TsRpCoOYnNnkM9CiDfyr/tvaE31C6GAzCK8yK1lUr3f5/aORSuM9PXtZNHOcjmZcd992kjbn
+nBWBoP7Bxyv7CR0UfoV5leI+0Rc7J/f1vwTixl2TyfX4q89KIeGFsLH6duYxZ/DYMiyER+DHj2X
4TOM5Y63XuDftyBWq/SN+u30rm1poe2ap/EsIkj468klXuy28sNoLN+XExRR5XGSoCmqwpHW78fu
0wFOLr5WMJebQ6DNp20Li3yzr7JUzkreyVANJLCK2d8eGpBtKKwuKl0Y02E1tvIkMtewfmi4svXf
Dup8w+X4Vdx0p9riS91Wb2JRLNr7rtiu5L3XyN/96MDfzlrf4t7Q7N4V91/A6oX4N103NYkJKdaf
VqIRKGS5KW6toYjRS9Jce0wudr8bQIowY9BdMYLnrINcPSuZT4xM1XPh64cfJ1rFMDMIUqmiGHRl
RVkC7YdxWWTr+DydsbwrrEQGUKyXrEIXumnPHa7fBb9Yl4IY0b7VoIr4w8ptgxhh2s5z+45ty01Y
n/4O6uwHlK+4qCa8a2FC6jhvnxPHSgqEeIL5wshOJ+eviDl+6HTikA/r2dxOqypbEbH6vQnFSLUq
Ed27y3q7m9NzsKSRh7GKXAXrIbiBU+UI/aAnZnh/z0g470aJ3nVt5D3NrPFnb+uLonZ1UPRA5aXd
3KMZCdaJ/84fmYABJ3DmKru1kS4j52iS6rrl/XyfjvTivAQKFGFrSc3evlihepTXC8/J9F7y1vGz
XE3h+/2LLTV+gtgPag6PsdRaT3AJm5hcL9gzjmBkeG6FYn/ylxb1ygHdqHA+JzmXe7VB3irCNa8F
+BCcmLsaEpVWvtbRELMazqMkMisiUEzk3AXVsnY8iaqZ3o3+QTaDxl9dB0+Sk7Q1pKTjBFqwWk7g
c81HwFug3bLEomgiw4WQvfN8VTi9k86LmEK0eYnwfv73u50z+DUS9e5mgeWpaTr0ibfvfGKPuKlp
khJk4S0TlHmN8dizrJk9+M4pBfQ/xgassxNXs8wfKK5HimiCVLvVCGSei4LnjFKFO2rBqP0oBIcb
gwtXhYkohn4FrNS/wvIq0qQhGAJo/8QmvzhD2zLTwROT5KdgLkfr4tiBu65NkqyL9wEh3+OzclJy
fg3vQ1N+PhBJMaCwxb27Vj02eKFpt0dxMMlO/4qny+2bRN6TlqZFXvywH4Z7ab1qVKljiFELHoDf
+gAjL1Eb32MTTY500HLUmgjyzZvZXw8Bz3hbugt/vzK3edq+km6xegZgyhIWiiR6DMOAu8NkqcTQ
VgDuAPfeSj9qiREAtlN9mqr9h3jJOfr9XV1OpTmHsqZplrsRE76Rh1e5ARuaoAQJvB83ZgkOjNyo
OFGDw4Rl2O1LgSz+Jp7ToDHs0o3kfrLFuSkhdNdNVvhbQ7RygUgyBncAz7TJaObzKk9uR/o8eAde
zCSXrEZaTDCoff6mjHGh/ocTIKUHsV8Xuvz7IElGIzxUxenTVwlAkX/9egDG7fsWiDa+ro22HsHk
sVDrxEYXGbFPQ8Qxue2tUXfbhHQ03tqxg26N+cQDgNmIH3RTd/thkRmOrpspdBWY7RReCalQt8vp
/JRM7yyEw/yTLe8m7ESkpp8ZAaU5PZoOgPYD+Axv/5dsoNpab7lvqxTr7gJp5VvlyB+AbS/Sd417
KBGTeg3RPJjddrjeKrnqqa4XfOPqG1YCBRHRQS6Ivkk22zJjmGmZLWoXNzuDBNxWfSxXZqGuvanx
Yn+LmgNg0uCvKkpTNEBJ6xReC87hG98/Xh5g7Y0Xym2QuhTm4N2ZocP7bbb4QEROZvfv4bGpl+Dz
jmkVDthb3x7KcXJp+XJvQBVH1Sd9JjEyPD//B01cSehT20Pc02SmvfHZXf3yXSWJebek4NmDJ04n
Lnkdms+cSXGkfG1tDbvwv8MuDyfLf2gyHbuzvsRhogsOwtPMyrTZNTvefLuR2S6U64GfqY8OcAsl
AImM77GSdacQiIntYaZbcIZOTr6CEKNapsIEKbi0618WbOLmgmSdZ99eE32H97b3DyogXqdN1VwW
bThWgUoYgCuUVkorGj8uG+GlCxOi2V0zi8Roq+WO4NqW+o+hrUal9aEkCfUcewJ83UDK3aCrWD9p
Bl2gAkURxpQmLdbjvG3xhMrzSHCHNEDL56aTzi/CsR/WfszHwNE5sK47OCPdSutojHGEzsmjQroc
b3YyzZHK2fdpMXgsWQMVTANfWFmm11V5X/JPhxIEIM8CmWSlw890idYFjVjimdji01sYj16EtGft
524CQoSzH4tlFDIkJOm2T4q3s9fWS3E6AA8oWY4pjUkVypgwVvN41iY6FNB+u/y1BCcnyJuqgL8L
PCLDYbmlvat1/U71iLHM/mIDbRQna0g20I/OfbZsJwyNMU+zATXbrRX0Qn8Yu2vCEZj/72yDixcd
BQ8yNtS/QB+vELqrngVpKCGzNP3JkJWMURdRcq+gMLQPsXjABTE6wYaLW0SvF+PST3oiOgpRWN7x
39Z7tKjRRScyvfXZNvnzFqWVlaLOZK3VxcjM6pS9P4X0dU5sBk+BxMQk39C5cIoaAJN0Zpa/OsqL
iSrUqHDNVGAGVh/8FVjE6glgaAtRag0XDkedFBVRntHMUnDYEmIZmZdRTKQ2qAHEph34iJ3MEOGR
/SJRJZqhxJcTMiDYi3ziUK77vomoAOS8lJXDgBZq0kHysXEZOkPHRnt7kLr/0mQiah6S00YdyUfV
IhFLQqBxVjpQOLquWzxShpL96rA9Vx6Vynyt3uQgpo+9j3qLufQHJ5Q+K0DNknPn2cO275N9Qzde
TREXwKcfb6JAo3j/MgnOQPbkMoEwYEpd5QRbdPNN/lj4Fqn5Yyxt171JVlrv2p9kEWLOFZd7A1vP
Aghdzrh618oYV2lW6XPmUvpE2rsHJSV+qvlYUva/rU3DE39Fwwy+s+1fH5K2xMf3QfduR91nVC+i
D0orSNM1w8L447J1eEuYCcbxdOvXjb2Up3itrboFruL/WfQhwG7ozy7kIFsGvh64otBHR6bBPpc2
i9o/ewZ7JI6avFOiUHhFL54ndv0LlOu5j70ZsiJnOu4qHTtAEReRpIn3wNxBtEog+iT6quzCxbEG
BMvfNNiFqkvRARs8VrIGmswqvrIXqnNozP/QZ7toh7duGH3shQ5a8zOVvx2Unzk/o78OVXoeMBeB
gbFUDtted9KiKHnivupOSCtD/NGIIP//piJhR7ejNV6iJAxFa3HflvWm6x/FYNcvC3DHFRXFq/iK
XF6zds4tK0LtZs/CkWimc6cAyynPGs1yZLlpW+ZDLZQgNv9BCbmf8G/u/EHf2mNDoO20KMCIdYmL
Z3iSyc8yQVa6YB2BKCXVh7r8Dng4mUMriJD/9wcSGiV4Kv0DbbM0uu2VDGPYojfP0Iy1QethpynK
v3Puw24ZbMf/RkY0RVv316GPgy/GhgoUH1M18IRDtPE48i977T76lFvrh4mJR9gCpliyoEvVGdcW
eZVgo45OwOzCGO8cnwEpOSJuF1j+j0+slUSzkdYVgX94L2LIT8tOqAUySc8yWnT0zDGp8Udza5Pq
FNV6epS8ifPxtUiyjPVrEL+k6aTm1Nrw+a+FCuIIbKUPtfhNhItNmK4xmwpz7M8DFfvlOkZlRlJF
9hK6fUQPnB5AMALvhwRXRl1WlGzvEaq+2/UZFc8Fwb5Su/NiO6+eHwAHVyBu1my/adIM3wjX9Nno
xOpO/06syftDOc6SpkyMAxL0sL8qor8mwtAOG5l4/F31/n1K8VH9HvS4/XQnIhOCHFLU+2ar2qlC
Nfw1N02JCsNuAqbHP4IXjb2JUHUfqA85sBPCf7xEj0ueYzinJjCaLMWDH0PE/bd0WklU4Am3zGKv
/WKC1r9Zgjlranx4uyKNxoHaiXgvYFypFIKMYNPtUDWi8uSwBVdBBjNNGhGBPxGKjRyGJioRWVuY
mG9/rwYCJy+NJ9BzzmRp1qf4algAfnO0gL3oYCHI9OqJn9UdX7oalKju/P++xDcBY+FMU7+ZchZK
fHjf72bNdqZF0OJBTJlH0AymI77XE6SHhoO0sFwfFGx9IHbVxf5zBoVWCvhosvE1ASzMPq1aPhb3
PrMf6a3/pZ0HXTOkvRbDuzUG0+BN7vytoVvZI46wpX3dvMYlSwcLDt8Tk6L6t08AMSRNUed86yBv
3ByZZwf/SUj3dlzAjtKfRCazoGD1M2gqNxPRL5pOTLPrhIzqVn2wtwygDplpdeQJJFHEImRfPFc8
0Joz7nEeFwEEnEY8nBMyxmzV2SChgK75V2aexQwV3n/VM5/aBWC0xkbPv4smp5dMHZBD8RxktSMi
7QidhZoJKkIH5a1M6nPnDownoMPL/vWucoRLe49AKDs/RRmY4IsQuA2S9jhlwrQUWLspiyVDal8/
3gEYzhKMU9TKTESVuSPXGoC96pNSSn+ZHKiIX2/xuzxvnXxzK37zUFpp/DzgRVCEaHyF8DE4o9n7
MD4R3OZQvNHilwX4ln+F3ClvBKdgFaQHBrYfsK/iBjZq2SEcl+cgUcgkTNjB+H3Quuj1zc6Kln76
LGzEQaTnd/YxOr6TonLbkk6nCEKR3XhP53tF3Jx0fPBZRrjMe1TvhoxRZW9gy7lVuEzexyePguVU
nQVvEtmkhcgY+aMfrnRPBkJkjMFFxJaOtwld0d9+9rkZZKO8YrNKp9VieCtMCdPJr25JFSzUdeoM
PJ7/+SWNwiCJjnHtqiexrgmxMc1eGoeAmLsLWFtGklZEDHubD8Ke9ekTxlxPyuInZ3k3HlNk/zQV
FBhSRKMLgY3znJ3P5DYqeujU0zB8Cqf9R1dfSGeeI65cT1SVtZoV9aqUxOe3D3vQHNOcgK876Jjm
UZ2f51FgwjHk7MJnTcvEPPwNuVR1Z+tQkH7e2hFNw0CpfFus+HH6U47+Cp3ICnFJpbUi6ly/aVPb
TW18sRWaKA62M2vHIyrmmi7XfC8VZi/uuHOnn5PGu9gvRp36z/3BqE5GYB7Gk4GaVWek49lqm1Po
+79fdbFJ3RPmKUkopM1QRO1FSn95OftDzIEQokA8zJQDkonYja/44HzI3CwZFIsbDQ4AzEf/6KS3
eQ99qWRXlZmbT9SFUTHlLK+TtTw7DD8cbmJhQkONwWHcXLq9rJh2n8wN1LRzLkdmXYZGsySG0sp/
xpcqwQEDkwvwhaAWBaU+qG6Qke7zIZ0+wOXyfpbfDfQ66oxfsnZRoxnBfA063QocLfIMJlRXDFZz
9V/dVPNagdKOF1VZIyx1M2Aj9h/9ClZnnE7KRyGXbFgxFNc03efnnXf/Tu7DDOe785A2IJ6322nf
cywm+KHNg2OeBfg2UPNM4MuV9vkhZzmJX1KOXOrL35t8foR38uN81fr5eD0o+51csJRaj0yZ+IVM
yEahBmasP6ycd2MP5I8YiuQ8VUCar9DDXXL1BU6bdN2S8duRCqSHQK8NTsnQamDLOogAOJ+5/9x0
SB6mSF0oI7R7CSfO6Zphkc4X7bGpHqHyNzkbQIPpSUQzbbJXDgcFQTjF7PoW2d9o3O/VkugFhMM+
Tdt5WvXmh75sJJgdSsQqbaeMBlhQsN9bWq6pMZY7w7XZgswtKRY7+o2vKKKiw+xeNWoSyYczxQMj
ExKl0nqGpwntRvh9KgZt3hsTI/RqoRNGjD2nCU0ySOEfKVq/J9S1MZ0Q7gyKKT5XiTXM6sW0Zt1E
iFxoIOVSArRWgKMhC0SBxQhaAvOyUIfGxDgSHBJM44QG8HI9Z1WzFCDdS1CSRFXVEO0XZjRnRXjI
tMf2kksZxLX/Wn4utpCppNmLFRSShd+pQt5c2vhVitQK7Ss3GdpDY/0Ks5HVxM8HnK0Xrefuw2u3
brOaZVBAtipjqGmubihEwwSnVvZU6ad03RyLArtBdKIKvQ5d7a5+YP077WXf5A0qtqhSwFG3BwaL
xj41Q2006TWBzvbFsQD827YF2+O7/jN4K9zLo2z5DsFDkrXl20+acpH9492MxPEPiW8Pz1v0+u4a
9ej/DoPEnqDHxgOeUQbze3tQXZgpvDuQgkDx19kVfsFMtdEU9jICdT0kC+9UeNvMWH+wgFElFgqp
rTqUTV1VPfhyCTWS12qZmNjdvxOcwgOe6JSbMq80bT8fAqN8If4bGi/rsqB+j58rUavI4k+vWVcn
GEIpDp4HghFl7/AZluPp8IglOhGCEzT4azNikaqxgF1waAiwjVIgsoVl1MKfd6+Xt+3NPbAjJKJ0
qpI38ZxLHVD0pjwd3QbgwbO+S7i8p0tgeSDHNYLnyNcqRCNSl7jHVMLAQzn3UnZ1RNr9179ksxya
7eQUy9/ztpy7uaL8FwdUMXs/w2LlGyTcTpAbZr0CXl4bZHuArTCr4xFV/ufzvFCi6Xvf8SiqnWRg
Lze/OVk6SvooNPbczma89OqKBxRgAg6RIOOWcIS45r7jaXCf9z2uCLNXiX9IA2X4MOZB7y8A98cQ
rqjbZGMZCBOtqIgjgz5vg2AdKRL9KP2Jon/uXx8p26MEFo3i1GdTZkFna2HKNES21hPZ746yRb8B
ClX0fhJMvdPyIuevFSPNHWKUOpSDhALR7oN+Znz0YAWhKw5X5gj+IpdCSYuarb7inFs+Cdw559OS
qSWhtFaOnjRcPd7AlRu+L8JlCNalfryDEiu71oz7xexASAH/t8HUmjVpd6KDREyhaBOT0F8UwKMQ
YWkpObRvKYni7N+dFo+9Qv37oRLl+uI8CBhHVD6IMzF2QdzhTPilulzxxvkkfecfrJEldIWSrrci
pxbPiwHSWTPi7NL/ENNWe/MWqQYWzYEGQhBx32X8f8sfmpyqgPxEkePZe79NvAmZrl+bRIiREgsr
RoXbpVqoGKQchZJqaCDuLMl+MnDCY1xBCkK5zSHLiSgRuoJr4uuTCMrjsB4+6DdIvp2pwUQI+Ffn
oCyYZ1hrTXF2u57SD2DpSL7WgLeYxxDRbwS7eNriOvUj/TYncen+ZD1+B8SJnfTkEi7KCU1Ui4Ru
q02K0DxxozAv2SWmQy4TAZ9TRMCrn7gVD7j1TPEDNFFag8e4BWBq8hayZT5p0yULZ2VCvupED9nv
T0y5dX1Mw5CZPucF3C9oULSW+VniV+uX83+e5oo3y5rLjSQj8JbYEcYeOaQVAHHSBDGXd8Z6bEe/
Ah5VKZ5XUmaq5jwX4atG5VHhGd247kLKW1XrM6v4Dv+LX1kzSlyco+yRZIPXtuUvTPU7nSghJF4h
rgX5jY3BzU/EQwE8gv+SNOQgXfet77PjljACwQxPbENYg13q0f74V+Q0NdHY4OqRr0QCP3kcetk6
7btOS0fL3OzzgxPobQ8fw3ddhmAy4uPVgZOWVLIhwQE72Ywk0P40mS/zGczFcVYnB5GHWL+xKx+l
E2docntRqkYhYnUrcfHKWpCyju298du4NolO+TMIsD/O2eS+9TupTXWcOuw/ZebV5waHnGQ4qrCu
LugPkeOkHGUvPKo5Oy4DHcGOZfSTpGKK30zZQnq3r/jRZE+0FAsbm9BBOxmEo3vH6C9v+SP+JGP0
+kjkuDbJZeqAPFjCZf9AJnEp+39dn80F9cFmPeyfvac7HNaYDFvLohCDGhb0yQBtIJnfC0DNne8i
uSDiFLSNckb3rEEOI5DQGaba1O0aBvOIJlym9bL1Bws4KnDXCVXnh4c7nxSoaixblS9dXqRDGxAX
rGwa/UUi8EItbbOdw6Tqctv842YWQzuRB52mOPAh3112iWYlht198myw+Ph0XqUtFgfReK0Cq1cy
j8Cae4SLIhZ2wo3u8vnWWaSXee2uoQZLWIO1hMlEx1oLS14VCLs0ZFpMVkzBfKS0WwFUTljmCiaC
uOTVbT35qO3taRXXy7zqjpTg/ESyB5xTTUkf5VdH/pSa8v4reQo59maY8tMuPCJhjYrJy14Ilg9j
mJVfJE2tKYQ/V5tUBFiDCGTEt10Hm1bdeA6A2o5h/b6Q+rZc/k8wLwv6QQ6ZBodRS/1TIiRAlZ1x
Pn6TD3mqtvEX3BdiAWINrwcQ/VgLwyKDJGnYOcljM0jkhZQzxRIYUtyjORtNP20jq5F0wdgofCR1
vwwPY7n8fMD1jyp7zcXIJtN19hjcSshPF0t8TthWgoACfIfMrXNRbeH8plVp/0JbKVbxvHrvGy2l
mt/L2IwRMSvW/lxauGMlBkS87c+fSc2Pxeufkd9SdVpG/b00fYMrzeIN+2wwvnAeyanY3JHPTGfy
82L+2uTU/KMNJhwskr3mZr+tgU7wVYfFpIpgtIH6Nx4S8UT9z6hBkFYibxkvC6tTKGkYFsv2elqV
FqgPLhTyDaNjEeseWCuOfxLALoSgb9+snnFxMlVtFhK/RDyR6NW2WYdxsCIFoxwt9bDAqnP8K54g
eZiFY3hqB2yb5gq0hOFeLWLY3DSKS7EiLD5Z0IiSQnQcKtC57yNTQWj0/QpHb1QH6gZFCJMwBXNq
2cNUJFXau3E04Y7CEVC3veZ2Pbimj5aqto1GZ811oyVvu9w+srLtQaO6eAQRQdG1H/NNuA65/qrs
s7ibnR3rBKkO10cGen9CtUWmvHuqIrPBvCL33OoMh3oWkNUVqmdMbSxS7mzpGPnY1XQ4/rcL1FuB
4J8coQfaT/SaH+y3UJekvPF6sBYDU3U+CcGlJyxU20efUPOEbYbgnb7iBzh9nUOhpvSIfSp1OA+B
uvgc7TwAKTidSnV2k9JF0W0ma6OMs6uYRm2S8gzuZM5aSZv5xYk/dySumXP8gUo+jbcdr24lqqye
Y/x556u4t3Rz3IvHbqRyTPauIVnKUkv+0Lb/QhBC5YU8mSHKXct3hWhFjGI1UIQhPy17kmIZPMNH
twUyYHW0SljBne9MZqtgsfApYX7eGVdDCB88CQa408at2HTh3ZUGaWSvEI0RGAecdYXI/n23y55L
W8Bw3Vv4wq75SDZvpk3mQl6LNzIhQkbBdMbOcsQSC9do5phP+i62JsUMfq0Y2lJdm+hmVb4ecy1b
/8GlRiBekAOPX6uslvA+ZGW27kkAtor2RozoJHuLT2JvI2fKQYmnhaYYdsG7rIkH0EpSo+xrQj39
OWv2dCKucJ29FvMfSBYCCB+Lc53MIESu5qeKYjgBp+9D0LyAEjSiKghW2APdlFGjDtnteRnaTIv3
+d0fHwK9voUIt8yzDgmefM2V0QYW0w+IC9t8T14gANW4fg9Iz/U8Pvf7ETSA8IfZEtTKBOFCPBOG
RXdPrJg2yw3pvy27Kj2Jbs2EPcWIB391sej5WAHp7EM6aTK2dcPVH3+nW5y3g1dJk1gRm4qamnsK
eBrj6wjCwjTJNlXa+dHcS2rR+YmwWAC7UDrDS6MRXrWOAusjvwcYigFO0i1whWGMa6h0D36kM43a
JUPXSl0X9pAH4JVP1utS3eVwg7hFGLAi9GjDyYh0yn1sLqyHWR2QrNpdONU+0USTUYEHg48VEYI6
SyjwkiQCAuFNkZthCHrQyfLptQK2Jr6eZ9C4zmAlAj87yjwxo0ZhyUU9SyixLgJLV+8JXubTPq8H
FZJIZSy8/WegbtozkTt3Ol9EgXDsdIgtOev0pO3xVTZilSG8XT5L4DJuD1buCLY1USQgqCfOWnCY
dDqiWCuwqALKeBJMN91tN1syCcxlXK6pamozBDxT43Mzk6UgfRlX5bV+ITdPyCjae6y0EYpt4nDc
v5De7/Fz7z8Y5vctIFJ+tiPYW5stbMGeZQk2Fu2l4B95nX6Lj31kKJDLMLOlGVGUl1Z3YWsU9SkI
Rpuf5SbMWb0zQWQ/5KkvEc48q2o6wDON+5D0iffn0NuZmfdxn76hLqqb5M+vgD9ZOP1mQenpnPSH
ygs/YT0esLJwV9/7H1hMQsioVtqSLCygDkd3jtt+/ZOler7yj1awvz72o8MyEXxvkCtf7H5KM9MA
Q8pwWQK9N+0V+I+/2rbAYPTDSzcO2kRsuwOqhwoub22QhC0DMhU0ZS2IZ4qvh01k9V0a1Y1hiHJg
Gdfz8q0tyXkER0zMKy3/SSmfGlqeOgRDZEziXYsjKj28cYXxjO6/jJ7Q4HxRxiM7ePbmFLi7xCV9
0RrZs0HQEr9Fwe4sXS6QV+fBGN16Z4VbtkdRjcMuCK+ppUiNyQGyMh2xATvUl+soPhLnM7isePK+
qWrRTa91dVYhb7OFGHqbZkvS+4J806JFO1gWLEhayx7oAu4n1N1Ezb+Au4OIUK1P3TeTmlXJeqo6
ZqE38zguXXW7jY5UfWoqvfZd0ca8brZnlFOmbIoTw8XD8+JZ5CpHAEL6BtHNZ1Up3krp0iyKPwqV
FDDSPM/a7pjxP2C5kGY/pBvEF4UknzBqwqN99pCliOl4CCeWfNxTC5xapRjcyFAhzxVxoq/O7m7R
7xOiSQK2gHx6X/MBpqfBh2L6aI1sk5FmtweFKffXWk9uLZvZArwt5eIHaY/ZO7ZlIJ/wbNgmTIYA
Sq92V886ENKeae66jMSbV2EUW8dbO+RoVbKQBp4AE9T1ZhOly+mW/oRNqDkgsAzUCNA4YWigzeid
RQDDdKDARzeUxcZD1REQKHhkfuSFLUbpePtDrxd2++MlyBem49jZAT1EQXGYO5/oyaKeuibs2rGz
D5sTDcB59g1rV9e3drTDqokhBQ6MU7JhF60UteO0j+Jdvo+1jEznd5m9Wk3S5AML0guWVPeN7if7
J7usnO7S0QMZGP7hvAtI3IZvyu4VN/uLHyGJv8pTVItRMvBFSD/wYNOLmyUiqAQXx8AoMdqlEYvn
u7YRv4VzhySkoQFXCCsyNAAJQyJqAtdwz7+IyrCyht6mA5GmQVz8b6T+UTl6WDlbv63M1ZEeTz+o
KHFXarsjUilfRggFEG9wHamZih7at9Ux26LrF7nFuvsmZr3zYAyuxv2MqUYxd8r8W4VnPhcrqltY
PgRgsDCc/3v/faWJ43VbLuMmn1b2gt4Piafsg0YWwCbI1qHQgmLB86WQI83WiUuIRiP00nw4MMt9
ab3UdSGEwp/g/USdHc3h2w07CQIv7mL50JerXtavN4lqchPdqt2utOkHIE9F7Bh4pBMKTflCQPmw
LscWuCo4Y0zm1O0T2BWHCoIthA3dAga6u1ilRabLdp/oiWNaX4kciHeMEZCnSfI+OesJtdws3rAL
9K1R4j/tLv/DawcjBbbIAVuX1jCimrS8sGQrCymnkm8UtXF0E+aJR8uILMJ1t6XrCCEztvtqXYww
GDbtCGV9/+tAUfGe0eXtqO+PfNUah5l2e8d2y5mto5wXatqsbnoawbQQpz7BUVh/gzRkMS+t+rSy
3IBgK3Jtw3ca3V6I60OzbRdA8g032BQ14DajlwJFGr3EZUecUyvr3YWY2oxpbDZOrFTojFLZ3t7c
4bIUlW2pc+Sg0AeajSANHnBbfritWiMZ4Mv294QjxHLbtDH9UKNpvgGeTLogTn9T3Srr8nUXMdgt
s3Eb/ElaS8+z0KadFfkzzM+XgVr+9RmTPEeIwF9lXyDrotRJhxgDva4pjGrH2dDbiW2aoHzUwtff
Jr+bRnFoercF6qYfbXoBELhjN3clFjiNqb1CduDG+PQSFaIMcnguoSUNi0CRhjHxbIj/pFtSUK8D
9jip/NMj5eKpc8/fIRyHEV52sqIoobnlyUrJXCzTHBrJbYLycB4eBNMbKiJHXCXyYM+7VAJKc/cF
hanqWkata6+Cpp2SWj/DAYFRjM3QlkctfCKbzf/LKhUwBDOEKp4Sl5n1JihCKTVwZsRX88NoDz58
I8QGbYBDW/H1t08FZwi0N0FYL2cWvkJbdbotw4P0aNDKkyyiqzOcoyGHwyAyMKRyBf7lLarFf6pI
wTXc1tQ5B7gdNjACmzPOeviyEyEjBfStwx319FKaPholndDtPRHThz9K2Fiu/DGDuFGdffMEzCae
URY5izV0JZNTKC5kWuV+yOSpKTFvBMx04SNMXcLPEcfJTqlO3IhQVLWJwyvTafDfYwKh31Yms+NP
NimghJnJEdArpTFFpWVCbkKYsCwW+L2aJC73ltwLv6Henfw4iSdv8wj8QZ2hn04BzglwBLIT3UwY
P7/mlksIAia+w7hbQC1TSy/cDH04bAKSZ1LtEBOuiM7GHtxsvAR0tVeOvVU6BuEksnekSOZ1aG2G
Go272ZMMk0azm1+P/hPEQmNXnX20Cdb/U/B4BZUm8hx7QRJSaH1Vqdg6AukxUrzKdhkK/H/ASi4c
fl1M/7X0wj6hh/IgwzbUUL8ciduENpuRlPLpSrT7ewl0rUsXsZWJ5BbCEmdG2e22K7IVWlJTgDZM
IBagm8cY/v0JgIhmZpqWijqIa1ZDUbotCPL5jQko0KvyTKaW8TzwrUCw0atwsj2wgugrKYavrBZY
RVaEvZ8sbfmPAz0347nTksGvxTHXtdB0LEVOzmW21yGS4X91XxFnVF6zAHk3IQ/+dJIS0WF4JJWc
DQSqjB1hxLM9zS7ZJLo7NBewZcEctjo+O90dLou1IQfCObPjBbYUMEd1bZ9RYzoVESV+I1ibSKs0
wyNKgzOs7pVgJGoYLj5/i3c0AcdD+g5U0W5FZHfILEOMPuHE+A34DmfxBjQrM1p2qzQ+Pd455iAj
clQ6EYyRc0WdIi+KEdvtKx7cbgXq1Ixy+B1xmvMCJpmhDISLdUVHYClYvsJxhKqzBJjf8YIdYhU1
zaZLsN0BaLI4yedZuRZ1T5BHZPya6F2vxbQ4AZ19SJ3fHtdbBEfU+s8enDWsWMk32tzPVokvL8yj
239LkMXFeQzMb9TeX4/LQB+zK6Y4me8qQxiR0EasNZH1ZBj4yNoG3M1WPUCtiAmRb9HbEw0hbL59
bPbJ7Nj2HsL3U7iplOLMuiVcLSvprAHdIvc1Vy939IerCRFBg+Zu/nppVnANrroPE4M7jdxYnXE0
M16oRKPayxq69q1gMVcmq6Pt3nyge5phdGL6Cp2zeNWXMcsGbKxwhY6bvIDNhIDzP1hPMprJhzBB
CMcuDC7/6DNGMAMMl5a+Xc4dGzFFuzQK9sD4vaUUCGkmSTf2B5HuS0H+FrQjpRFQn+pS6ffiPAL9
i9L+80JRj6oIul8CcdCTXc+9sp2miShFELQLHgx6VDOJOcNIvW1aVjd9yamT6uZO+UfEMQxPID7g
t6w6MdR1GZoV6B9X/6/XD1JNxcsgntvkn4q8KyawMm79MSm7rthY7Sc6Hph2JmQMZKj+41hBcCbk
ZjLoNl0vi2Zb3uiFblExCeBc5Q0cLmBgHUPzHg5ZCBXa1Af+A0axC2/slxQzThP9jwXeoAi+oiNM
G1kRYsuJorfwSD9JLOzlFxKk/DuBsmqBYzpVYrxIdyKawiWkGwA8obVBRCHkh9CvBwkQlq8xdH3t
0qITlsXexRgGUS3NGIaE24CbWN2afZwM5tU6oo/8vCB2cQUloH+n4dQBKCSkkEyjgPRYSd6H5urT
vUn3llAdX4kTm0Omd50eHrrqaOnkS+Fp7Kfx/RbDXAlX3SkhcAvfpWz3YZLSBEQ2SoemFwbtmlQq
uCKyByLZsdAC187pe3SEmS9eMrMGGUI+p33T1cbz8ZF2R03kOfB6ln+eQ1VPPBPJChHcmvtlWHRJ
4ytgbwDalZTlnApq/T/aLY9z0NNiHZ8HG9s6fujgprOK2ZtRYnebeeKS3aQHEH8kNLZiK+b1KDq0
+2UF4yjb9u9fHVYOmaF/1nLA3jvGaDzYnOR2yQs35tAFts5ZwmsOQ6mtmGieS6n9jHsNx15sEMDG
YWKXsib/bMrCl4gjMHYrfA6FI6mdhbT5pXQSMM5F4QgSycPPmOsdfTEb6n6KSuhlKWni21F9/sEy
2zz5ptpKPiAGMVStQyYUZFZsxBTTuFiFGFWQWKBkQlvss5cwzXT++s3rUaRnuad/HoW9iNXU8tP2
2hn/Dlz9NgcrhiypNJOuoCjhQDG7OGF2h/KqcSiXNOWJM8VNwSI2Nnf+6Ryax0CUp6VaoDG1kYcj
dMSwg5fxSqLGzMiRCV13Z5nyzcmWCA/isxnBxBHTngOn6SViUNS7Yrz5OKg2nk9U5cdH0/9lOgYG
J5mjy8k13wTah5h9s76oR02OfWGLCbU2q6y6PL4M9b5N80VH7qdEC0KZi/YleZXk0wnb4HMVIp8M
wzIQ6hd2HypKhe4YOia1Xi+dhZ7JB+X6nyyQyLHEy3CJHD7pGzwmSCy2wubk8IAdvsXwoAschKDA
Vf/yUB+M0hI43vhAUHihT8/416jcILo6OcofZXECbx8R5MIUXiIHX9LxPvvYHpKfW79qz5rVFpU5
0BsIegwGowPFPaEZHoIXnX/6LvfbH28hgLn90Eqo1y2pbS5nLu+17LYdR19vx8eMFtII3qSWhT66
WkQVaSlZtdesOTkI2UYMBAba+RvxcMJz7tqlnxltC2886en9v2H6GEofZ4q7llG7vKcW+JRaj5lE
6qO8rGYy1alO8YZt/vhI27fPg5PJjf5pKycdOKv/T3yC2/MY3PPADMEwoylGy8k/C3Mdf/DB5gk7
Aw1UtB6+4s7gecwbAuaFyMSwbYWuwo2bVgwLfCHIfovicl8O2CKMIurxgymvEpRYQh7AyBLDyFGs
f/wUbLJr1pTcyfwoXbTf1qo1bCC2ZC+HIEm9Lq0PgsrbXkd6IQh9i9Xt1AtHg+D5kIPlx3NYS3Lp
Z+q2gaPwggUpYjN1n2zhgeALc5F8Y3y/to9QKXDHEjGwA2o2GLfYyMbxBh9pO7pzFMg9QRF02W/8
3+ef7K7si7SnkYILimoJCuBzaR5pMkov4HpZ0XhZti7WWtnOgww5MMk0csgHuLYZ9HcZOg3HBCZN
Y/pxBAbjcuy6tbVuzIhv1Ofk5w9fEB0g0MVA4x6rKTrgO4bY12/0u0ANKaWWVrKB6NYyH9I/+fuE
CjIj4djwVXF1A/F3n5uHC/2tN+Y7NiXy3Pz9TsAXRGSAGI+8zUT+U8HvVFkzBk0gMyC4Mst6JdrD
0SCsTna1/2lyYe9Mgp8ITyVOnIqPMzE1C3TrXUCtwG3O5JfyxX8/RxJyvpx9qMm9qwWzqgf7s2F4
/j72iYXRqihP0A7GCPRp2bWiVvXes65+4kcnQh0+BSfGH8rAQqBwXbR0oJCZxUBKOobRmLYsaJ1p
GwUQHDyxsJM58LkxTugPIb5kHy0k5/bWVfC2zhxTbPeQcvrRxktBlBGbEENbQC8fgOIh3ZZwvGws
IhiZh83i8DpAGQY9dLIplPTnBdWrbqzk0yeyVIRHJL9lbt1kd5H/cxOKxbapee6hCPq/EU6tqnMk
AKUFlW9PuKGHGS8jbe6R8Bpmb18h/iGicpPlTw/LIJHH/6MjE2CXJpozEbot8Vy4oywOLsfz3A/X
PQhx9cTqE8G0d79W05DSMxAoAJTDlopH4kSfHkGAuSUS5PdWEfr/SFNuKoqnEGGBeMtYchMYRhPC
yAsYPOO0VZ+PKmv7FJtxguEK5Xvfp7tKq/02a+fY3KVgrP2OcVmRxD1YQ1LNlSyGNe1S9glD7SAO
mOO1oyvY52Jc1o/ERJAXEXwJZPB3NqIRyXluE5QImRsGS5330Ma1/azuq/86ALJPjDb4lPIt48RV
vy//h6RdMSOFkWrEuyYrKIh7DC0iQjfRwu5mKaU9NzAyP3nmHhpazpzviBx8IFiDo/z0+Ai45zV9
XSKBZjzrpa0lfX/GJJb8dKTIISuDx2dT/j1gZ3XDEaQxjILpYDRZkjXsbtXu5mjwzcVH1hmdiavw
GWc1eyNTp8JmAXsBwrrFKy2/AcXxqdag5MlQIoxhYPR8Jo+lBguawtdXbV+p3qT1PNrlXEaU/kAV
hXPSBlYgYRpBuW1nPlbCCLKzFDn2ztvDc9HX2BX9J+uh20DeaqCIksdKz54nZGE6pHb/yUZxXdaS
i/MM/bLpT2LDLBG0WQbpc7SzpR4beHK3hF5FKVoty8B262utbaNCCg91nIVtwSUE1QW/MiPgs1b4
xnR/iZkD4X04EAiaXfoltZV9S85VFt+No5avquYtvBVttfxWHNNZ/8Lzn7evDa1pyDO9/PJX2uyO
gvoumzw9zSvUW3S0/jKOFq8Z6tDaLSuiKMrRPg/F43+EoUrIEybjs7McYB0kvdXqfkX8KL55/LNP
0vNzec6y4jjlI0yqZKCW9HZYp6YQ442nS0sKJLEyPmsjqXEjReqjp8oc0H0DRSAvP7EsuD1hsrDd
pjo+rCahNgSl8EOq3F6RdfLZra3nqdcJlFG0C3dPz8WTUQP2mcUXTYvPwZ5NHw3pu7OXn0jwxIFA
CX4bVgkPaU03ptAJ0UATmd5kFAeS0HlOhKINFfO/xXvS2YM2y8a2u1u89O6n65RLzr02phl3PtOg
wHRPktuWGq8JdmXViROd2BrWD5b0pc6dEjBwmMqI3Et26s424GRP+Y0BJDY/OkdbKoQcWhkbZOJx
QzotsxSHgQc8HrdeB2BCt7uozrfkNOGX2d+6k4BQInOeWOtfPXjUoQhj9frQwkbasrYaJWdQuuTk
v1+GSejTVgOmcRmzienh0jaEgG1EIvChaoEjCZHHNt6+qmRA8QqEjQ7gR5zb1Lw/bWls/sWlWcVC
ZL2M1jQFr9ozbzM7bKwwVdYocLeM1N2WvLMzll1kMUe0rVaN5LcnOS1sJcy/hcgTxUxGeQcl0CUJ
iaLqo9XVpIhED4FQlW69pck3LIlHJ6E0AFDOhQ72zt84O+HqNwjtw4R3hbo0ooZp7G65BGWRzEPV
JxkXxUqVb4sZn1O5NakKhPKb9fTIDVpNA43LiAnlP1jSRN2DGmgw3v/JWWrwTXuGKg8an2hrZ1jl
9T67kNowBGdTaTz3xA6pXth8jv3f69jAfifTZsR+EQzZp16i2PzgPAd/8eTW5B/cmTRdpsPohn+9
dY/x4xJSz8KxC3+cnCUqtJzbh6T1WWjT4r531QAhktne3cSIgad8cpPtmTQqkeUKDReYlI1bwHCz
kzEzrF7LI8chfsGh99+QXWTuAkRkthwRc85XxN25g6msn0FTlYqVm84M/CevU3GY23INfmXXskZb
QVWgx+W/x4I4G3aIPCXA4CdNcdOuvZfgx66uK62QQplPyhGoLunDvU8oNOwxc4lwh8WiI/NK2QcV
TNsPX8jL0NBESVvECfbT1Nn5D5bobq9v8Ws2lCeOunwoxSdRH4MCZJ9y35QoZq5NnoHpnSCvUL3p
6CT6mpwH4JK46YVOAyK36csj1yOaHD8pqQoHPGwjZU7cyoHFoxJpCoOiGBJPDxJknteMCWf8E/to
9AgFKWcK0WbuWjC1B/emo5vaYku5Ov98SX1lj3cqhRHTF6W5SkxK+zq+gEScIYajWQv6bTvTXZ/3
Jdps+Jet+9SjimumQgcRAq8C9EfJ2mxoscsJlP3D3g2iFV9WZ7v5sVpF/JijLnnvg8zE88kAVXaa
1IckSoG48uxEJUzXiYxx2KwNfPhrle0YjjP0v4GaN1N9UYsKr5QTNM6JNJLdj0iuDXj+OY3EDrjH
ZMVEThJCVeoC12bArXJ2sZgM3zNTKng0EJZs04VtFYvI3RdFwf1TQCPpRgGoNISmOu6RmO4DwGTc
h14LGqYOSrdRhcqMLFaUny2vDIvT8yk+gkEMXp2RBLgxYzy7VanwDM/uECpuigB7N7pX+Eq5CuNX
ClKtORQI7mJEqxAIBExJtGuiAdV7wMse8DskSyGJBGmaV4DABz9YtYzZCEViXC3uxRqyWLfJNQPG
sXOPfJbtPgT4wuO5ILPHujIIHRF3VMGHXMTCfONx8AtO+kneiRkzZiMbnV/INo43UkAUUlKxqWn4
rsaTd/Yp0HDFPNPmRjsNDIaNkYFSmwJW1TpLaurw5kk0g8j+VSw90tLvlga+o+Z8Z1xfjeCyHu6c
mdqvrvc1+sVJjw+R46l95eGjd3Y1Fz8PJgZKC4JcZ+kckkpsXdZ04NJbW4MEaPJ+kYKRrgoSIoIj
/s2d2tt+dwaW89Yn/miPgDBTw5U2pldBmtYuuFrZyDf1lXZ+oppua90nDbSsbWGZ3lD6NdTpj2Fq
hBVEW6eyt0iHHn62GiZ33TaSshDsnMzld+gklwAb3d7AqZ1uuGKZ+AsTHAc9fqe65SWKQJSqEE3T
Q3IK6uV0lqZtlz9b/DHefCT353KSfGACgHwxeK6mJpeVkUV1glSsY9e+yw2rM1CTy5K4yueLsQ4T
Cqt2LQLIlPv047Xeede0bL0tCo4atckXaFNDD4GbaCf2kBG5TP8/UvB2pEIchVlb8yhK6UvMahai
/h0RtlBRM3nspn4AdPJN0nM8f2Xf100KM0pdCbWbyn3SrqxSy39qIpW3zP3D6U7jbTY6n2T1tV00
KDpyQZsmDFlISzup8Rwu3yHxJ7sBILDrhZ3YJuaVrZbGRWzpbUj++uZxOVYaWJaJMdy/tHCGTksA
/Aoys+zr8C+WHf+HnlM2UI8q/ng5cS0tQDiJEw5sl8T/QJor0D3+ng4M6dSuQY3hDuZV42Fvt/fk
Dku+isQ/5X0490NYqBF4LmybZrM1QHqPUMBPFgOMUsHhiqoSPzEoR9aH7/PX7grckFPbeOfLBo5d
leg+bqnrTdoc91Hj8XijM+CdzlLwcxo4HQsiXrcjF8s5sv7zUiAKT8rBW/xIRBVh/mAFur4VY3/v
sQfIGnv3o8lAhmdAV+kf+svAh4k3SoIpdwFWGOIKEPT33ZM90CTXSf63OgE1Rcoqhk3PkZ3Hmtws
wucaTnHyL2pUNciqkYJfoiZOL6FPrVFlnpzopBYKJg+qME64OYhnAgXTh3P4EmrjTtIPZWoy3DnK
EhwFVSXyN1yNkxXCHJmX09vC+cm01mTeIt9CnjfhrOS/STnmZZ0B8yfElbtiknarfQNIAJ2Azcpp
jxNxP3dYcHV/2vmUs5yxDPBe+07eT/80ouRHP39jr5wUi9llhhNd1fpb+kj52nHnjeoJGLstEewv
M6GMGMUmauXbSWtSB7Odu3C3V2HZyPWSJAeAbai3R5rr/CpyXJrd3e/7WoK9XijCwowWygV41Dr5
TvMpTl5hRcelA9Wr02UvslbuSAwRfu/j/SnnL2nS7ypDbYrwqedTbt3h69pY3l/kPy7pXceXFUfb
QEsxuMYSt5/fPPvFZDs6eCOm4nOHcCnMtibheRejyZD3tR7OL4MZf0BKHxWdvD6GA5k66yTPQdfe
ISub2VsyVlrDx8Gq1VbOKp/poO66b5NqpC4h7uNA7b0jsUcNvO1cmoypBKGLIW8ibgySosGmp17W
4EpPGYUPY3v0jCI986AKiNc/YJJeyANsvRFn6fsE12sHXXIDplGc2XuYSHaK4qys/urWn8zhtRbJ
fwTahIqx1IkD+mWWvexGcHDM43KGMCw2BQvSUTKw7uBOHBPKZX3u4Uy9CZvfATq90O14O0YN5puJ
xGXN752g05w33w7M4t8RoexJkWymieJupt4nO3lnDLHe23UZM7UtjDHskLzn/u8Es6VIa/6mNh4l
53RBTcWUg5vF/TQNoPid6T2eMkoj0YkBMWepibC6ExHAiQEnWJnIrJNbw3/RZi/4WSaYaVYDvGHC
jQBe1UIem3QgAL5dIO6ERGkXHxV1WBBmhFq/flu8zSOAyly4lnEKlhS+bq+Vvtqe5INFKHcpvN03
GSx8mScpJwDiOG3Lspz/+BNAkxnqu+b+73zrZenMM/HOKfmLl0JJc0h2TlIh4U0pzwQ2+NyuoQww
cWHavHrvPEbJA1IeSzHaZ4WTC+TC289CHQt9xhWhQ7lubB1O2VVmsNaWIOFhGvwIoPQUB1rLDbUr
hrFmn4MFm3XaYIGQ+grigDpo9832z5QBJDJ56lxS5DCLeGvvnGM6dFfnvLY9vIzIBIfy5/FOWF2c
meDe4bxh1U3YM7/WZRRoCfKxVHDhcR7bySamhua8L6vE74m1rx3SelXgFUE3EyGPXYaJ/6Y/ETnq
2Gh2gm2X6LUB8U4JBWScyehHM+Wt1JnAT7nFBxaQvBY8nkRYFASzAAxdtHAi/Wg8P0DhhOHQH855
rZb4607FmeJxIHGwIgeeu1KX2ttjDo7f855quhCFPLgJSIGShVuC+8O9C576Z6+zy2Yfkyy7bdrw
nKysbjDkOYPzZUHdqj3pI/f7/JqJo11BEacbb/zInlUjjkRa7KA3nI9gbrlZ1hddSAvfvZv61XZA
5TBICd8xICPC/W6yMgbfuDSXKY6BEUH3Y/Mr0dJycakKLO9jEqO+CwrlnG6a7RAl0fOtxt2Hy1kq
CuI7sA0BjhHZk6KEGK4WEtB51iOzDtfbBtUikkbI6U2XBFzDZZRCR35IJC4P89+EjPp/gZVog6S4
ezrr1xNjuRUt+GzJI4Xxk+u/8UJsSFEb5T3sl6FjvHGAcs08O2jtFLsX8BwC//LKooyRbc7aJwt0
QS+sXCm2IMPs2+H/C1gRWIwFFx/TDoPLtuuXA/TBA65tyfoBSybE3vyM73iAHZakDnDPfeXShgpS
JV2XXUOsy6wP++5r84Cg+eFifXmTo7VHWwV33y6o0id93nS35JZWpDqDGb16i22yScxAUOfWCymE
a+MKlXgljiHs6HURQcsfQMWbVX0y0lyNOvMILYgJoBZpaTQracjAchxn/5bylLmWobOvlizVfSPZ
ye5XlkLFh6crSKPZKOfJfQ2GMBOowq41CfNUnLpBBaXnAaC8iVmztCsJGv92w+d2Dyl5hYjx+C0x
pLUT2ZzoodwHgdSNyo9lQdj6zsha7izknJ4BiOeU/5iMK3fT+F97eudujk+MT4zDeJhcEaImpAAp
WvaonJKZsJaL+NZiOAa3K3d35AUF5uI2ndSLlrSON/+SAW1KFYnwNxyNlyyu1NemQcucqJN/99IZ
LQMpHwkK8m2MU+/OUkJTR3blXQ06zOqvg6QtD3M7YcoK4AcAiwipSNLyEHDQUh4O4BOAl5n44B6k
BJT74b8r4HlEXGmeZZCmpUiajr/M8ktpsQiDiOsDSDqav+hYaiAFoBhTkkCUMYTQIsD6kJbNMuHJ
FApwLbSiAkRAw9WTf34nrAwaK5WtHnSyDRxjuMlqsYNWTO/hydyaPqTBxY0wXFNSte+LhKr4+Nzt
ZfSoQOOYfFyC6PBmYCde5x4LQXKxwbk4yeF/Ag2EPLgzmeMLXzMr8Yn/Fp0TnYKsYrdAg6yDPzlo
GuMxg+H06jhJs0zj7STGzAvlsFLnhy0Qm1ju0xFQgKp6r2pWpGLy9ES10lh9F3XvrZvD73Xt/e7X
56TPRkw+/lmrvzRyMAoem0v4jqpZKDtQZYsK8O/h1RkeHTfYknmQy6fsaeYhPcMqhTTqMtiQ85mW
4zhUuwUoiG2UZQ1ha1jsCoou5bs8THDeVMGERQ2z/mJdKxaXLoLxLz+EVXkVsI0XJcEUa21ov/i8
pyUWgfNtZkOb6TfzFfGMev4lF2OI7higJdFAUM5UeY7y9ZN4XLRzPRW8DryBU0fEv+qZiCyjc98/
qAWoRrmncckUyhYY7kLKc6KH+H5fZHxaYTCyCbYd7NN7a/vTrMohTZhsZi5mKGS0fg4MXEKFpBQm
EBgNmx0h+UppzvHiFtxLKNTHNwO1Jzr818d4tnC5HgSy/qbzNH/aLUFP2+Ys/7KSF0p66SnljQ+Y
KTmYFiihDQ0JzAH1jsBbvsiErM8ga98ch9p1L3sSBsRERlY4xQvCTFkhiGeY+3v6NMvZTGPRJ++l
o2J78zUBMa4YSpdtPuFfWcOYvbBRcbGNwf4M9uEiRcmt6Tk3EKkxU/ZXqL/9YID6WYGNJ/YPkWPa
NVbEVikscxXmd8BRbZAOMWl9J+xxYSWvvFQPmS3a6AmpmX+BUCYq1OHzmdtnlwfX3BUapux97KHo
KR3JSwE96sZ0wnAG8Zoj8Ym74yN+ZjNf/0HXkr7icsR4FakLWBJxGz68/bMIkIxmsYM6VigXfRdl
DrwMTPdeQ9tCzfMFPXykdeeXMqUC9qo5AfxBzUEFqpKx6CW0MC/Hz5TGgs4IuZBJpXKx3fPzfhBW
jMIMAA0b97Uk6P/5+HwzXQDxgGL+06xL7+rEIoK2+L3Ruo51H/BlGVtgUK+sv5Opj6v7Zxxp0yoF
QDZ5ZiGVThXotHDRu4gbrP5dxEHixo6ZTCvao0k2/zo0YTpMkcONybkxD7g/2efZeSO9mmV47ytO
I3C5j412s9/ByvYjjTe97K+dRE/exsVsMsfTCjhCSZ3m0XMjt3+0mHKM9QLTHU3oPqFMRTy7UzzL
cjMtegYRQLVqIHfpuOLCung6d/BGGD9Wor/f74tf3/TZTpoCi2B6AHjvt7La+j4seuBtgPjPU9hc
uhMEkht2rGj73chBqklX+zLEjy5zIo2ZVHHltZRPw0GGUVWsb7Av2K/b2LDrQfJp4UFDS2639aAc
7alvzttrMDLrW82g4d+dQFvDC0+1XLAvKTFt3Ib7JKPK/Y5CRqmJn6uNQWNsu5AfeyG+LNmts9+h
EHXaAHsOxu3VyCPMCbljZjcUMqSx0rFHZLIF24wyB8ixMfCYlAmDEj/91IPWfu25GEIRSJGgpphJ
spHtStOufA/iS9wdRFolnUmhhpo4nFhcVt84yuf78uilyMNiOwTjip3+IKnW2+dk3hZ5gKZkRkHl
TB21xOeKW+ucby+8e5Cq39PbbD0F8g4YOG/b+93gXiUQLWqewmyngZ5UopqtDq9x+C1aSTKnLCa7
YVnOvM+wQ8Rm4pGlAlLKThEYQoEScqVXEyUE2lYO8qFunx5IywpdxXZ2+rWtaghU9OBggF85YaGV
KutOtzHbheRqZQAGlAP4NmUiOyXbg13l4/B1VV9W+eAemshM9Lj6JnIYndN4rOIQYfmbFyHY826y
J9Bgi+VwtWYOSx8+ddrvUyf3P0q1qN50hDfSB/s9LIKWJ3NAo/F38sQnsAUNwI9rIhCcdZkTsosc
Ojg6twKG9Q8/Q6zTL3sgTn8M3KDJWXxK45NVx5nY4LWsf2SrsDe6oQCrIeDw+5ALvelLMCFOXIDP
51ZuK6uiVEA7oLmOLkRLp3kIw1MyEvzWDvOlUPIJ0hhpl+u7CE/Bha9QeJ4duU26nJhBZcERPxGL
zERPounCPHt6cc47vFNmot68FSZjFKDm3HSEgwSbIWqvmEBSfdXr+mT7Xw7ZJh8XNcA/4xDeZpRk
3f+ifx0I6S7xXA0jOXmPs1aASf4so+o9WL8q2wY6wrF0l6gqtS1NyThmV3iGllcoToFGKBXgZVbS
RfqwjmFNNzetYRHf5tH3rF5j202GWREHRx90Gk68EhY9Ey9GyoLoR/ZeUhnGPtdGFX/Ty1Iq9M+A
x9r5Fn3T4o54wRsEH0ET/jPKS74b02wZwNGZN4LAUWFFcFXwNpWKYGC+Q36jpytQOriQc+SnHops
bECxCsp8+nnCrjEJm7LN0Zrnk0fqegO5uF1cnb7s170WNKCXIhv2ql4zFcbAOU5AGL7Y+E5I58B/
Q7LTvV6tbTzhNHZubHAtsuq1C6xqryiop7aCoflSF78eEhEMoZ5ef6OyEXY+wqHv4CTjvnduDkse
d9QRpxy4XRFFsVCnlnOqdMu08rDluuAqwXNXb21kxJEfy9+Yo5zIYARPcmMZT0fb3nEb5o77oof9
7Kcn9qZN3HNx/ArsB/HgIvojB7wWwCmVNxNtA/7Fev5oWoTGsKgcQw61HwoLSPHXVagEwbvuG2oM
88nhcGNIG+wfyl3LRvcsmHho7KHOHMa5hdPUCq6at6BFRCebhCSo/BW8Go5P+H91KJ1Hrp3/XIGv
2pIwIO5i9vuEoFq1rM5chTBNMlxTGtRIzz8rZSzcYh6lefwiaQvefVYSOop9jDLN5msVNPxqD66F
fYlzvhBwySHNbzrLkADeUiXsswalDjQ39azC+9st/4Zi1w+eOl8EIQQWDkvTHWDZNI9QzNs6kabm
3PkUhTD+7pVZIbBQxrfaM3rQPLIOD1BZDsP5Nx+6gN8DPPKScVblxIS81awfFZDo7QpUVO2t/Xiw
Pycf2BANAJNyNrj1Az/80gmY6jBhLtpTqXPyhyvELThdIggJGo5CFMvCd17RcLtqk+1WHdsVO5Le
d5wtL9BBBVnYnONNMS/73EkbV0XdPnCXaA2nh0CwrLfvDc9boeV8gb4mvQR/QsWwFhaW0abjJbvZ
/SYzl+hm66O1KFrn9MIKSPATS59MrEiPg6kahany8CSxHV7eYi9aOswMQ8ycdD4pEAYlmD0kh0Vm
GKZHypYhDKNDrcXaMlDCE/6R29RuI0pmCXLDHFJN4wZCOdLb2bhXEamKSmjdASgwQLBVCBO2+ylD
DaxSSgSzqwlJHnCEPEm/EkjNiS4S1yAtwqk80J63VjA1JotaUpvjOoHg45HiC4GAl/s9OsxcXHix
CrnwKa6K9Ets9mtopR3k3VTEJBoitPDW/xCuBWLDkbkzGVWGe71t0+BGHir1w78MHHE9VgvYcgMb
eleB5UFuZzSq2vqTSiHZra/u1uYFOrVHaXapxRlBZarMYROPpyNEfWW9MS+1Fpq2Cl6v6riLdCqC
cCmAQLlV+BQB7ipolaIwk0q7t7BWGK0pMwvFesfhyF7XmcPru2xWwazyV/GilD+6J57878Jsox6e
UgceRstgQfuVwL/Tw8tZ6V6TivfJe33kWr5wUe6ZKSVtcorvyJ5WmXTQ1mLuS33Zbr3XWvipRjEu
kZmpY/kCMjvbLrfBa/UTmpYeeidp21O+p0l2UsN4qxgz+Xsl46VngJCQ1+xwNx/Ot88xVbFl5Fdi
L44/SiO4tpBdRzWSFpurx0EwjKB8KDFo6Z0u9D/ElLi44y8EQG1GQ0TZNcEZIjgHCkeetEjFz96/
LSPe0tSoZQg6yjlkmzLeI9YxgcyrbLueQDDWKZkwyvW4PgFm3zxOqzS8a2jnAie5PqI1FvKvT/ni
00atUDRJk32xIOzXBug+pc1Vsbgrzj9rQAsyQlg0ZspyMpl5RKnEwY/DZkTu58KPi52M6TSYnoVE
eKpW4KFv2PTT4/tZ1/pBq6fGeYOIm+flBaAA9A1I94aYPstvqwjvfYrRciCKYTXFNTcF33jEJOgg
2LDQjnx/VN/M/rEmyv7hs70bbwn/tnZYd0d5jwPQSvnESljajbuKaTx3D1AeSBbGDv6kLJtji5lY
3KSL0oO/5z0GLYFK34J2E7g0v+iXekUm8Bj52J56QJ6jO+g1coyjkxpNpayhzi1iz9CkLL68VYRN
Nnhz5jI7cbcbS2rkwoYRvr32g/EF/PqSoov42kHelhGCIy7yQ6KoW4QC/oeQ78oSMTof2pxIdIGL
vwUWAjQ5nLOOMC2SiSD5B4Eiak7mAWQdZc19LnqTG+BRlYu0yFG6nAfyYzy1zwOpxoWwvgxVFr5A
/KyBp1NU6kbUx3NXxAyIsz/BirURpg6wUy/JEO2xoBMC9MZj1gPGruCXx5w2SLY3iqmWkcxzrbGV
3j8ElxHDK6rF9FnxJyNN7q4axWz+6cO3bxyodW1ZzidPvrb32j56zYfYNckXpzifpmwc7SQecDbD
J+yE9Ji5pVx4Mxkg9BGwlfQJZ/zG3lJtJSIYOl9CTJnjsjfgSLUb2Zq7EGQAGaRHMlb6xxAglIKK
TjsFfLPNeKKJk4WI82WHsA14bDCxDPVb7BDY7rFPOHLL9rMf2/7j8tsis/ETlTKv1Dmg0Fo6CT6v
ZCvlaj5smb9SbPtd8FR3uDQkPSF9IiGl1yAVJhJTYo2UD84eA53ZZP2MPQ0xV/K1St/aBHJJ+mdc
IzJFk8crqseFT5zHiCD14RYf432Zmwglag2WU+Wx66QybGXdZ+keq0ByercTcQr12VZDfdLMtqH+
2tU5Zl6Vc6JEsREzwSzv69MklhL2IFgX4khE2+d99QK3QQGb3cfu0yaWyG6/Lv3kX6PEHeL/Zria
IVxXbNUzVQ0Tz4eE98zDAXEVeS9A7QKC39IWm36Nr+IR+R1+OkxFZxYiC/U22X72VkCgab8MNGqK
nrwR0XP798dBnPbOgRkEsQiTCFYxNwJCGgFwofysJaKjDkCnXk0rOf51L2Ch3g7/U1rp12u2Ymk4
rQch+F5CZMyQdu+fLx4w2/OR+8Cg/n3up9wPV/cxZGi9RuUr7uu/sGUwzB7g+0zkoaI5mBXd4j62
olQ8dJTcxZ1cRJZlvVVi9NwJAbQBqlB0Ai2e/+cOkh5dVbaFgqI85fKM9shJQEF3mA4qb42Q1MOq
+zwtUEiKWa9k7SNwtOhiLnAHlwgCOUMQRuffcZhXZP+KIabdCyS7gix2JbhDTIF+Bxyq4BVt4SaR
+EKoGHUvlxEVcrRC+AhrFaZJmRPCpMnPRpB6BTsSl4brdevV91XpFgwXy3u8PvtrWDaOHAiq4Uj8
aEvMmrc9489fClmRf9Poqi4nG5JrgAg964NeJ7SpxVDJqEpyCS8Lif4tEhhs7yVnayGQB0II6c+J
qXnn/pun/BO9hwi2x6fScWuHrKufNLaxUYkZRINbthIJxObuqDG0MOp5KG57vDxMe27+2LfvpHjM
XZbkK3ZFEzPdPSnd+3bhbnV63pgt5DrVxcRXEr05gvCM1x1cW55F4prgEV08FQAtdWGjc2pxgvQF
LWcKRGq9HOPFk5KdyIFkyypQ9s6spi87m2cOHfG/FLFKuEr+QZMobyT5Alq/vCuhlalRrI+OjdYf
4FUH3VF8tU6lY3Xk7GAsivLinhU7pwj+6B9gwCLxv1D7O7OYIoWt1vTft09sW9jxwSux4A9gSg4l
unOwOPiH0iAjhja/8DnGX/M6tlBF0SBlCY+teXSmUtgFQiuseul1zosPeq2P9Lgo6mBPnuUyfO0H
zjEUq5hd7Wc5QaCxcAIj+pxbUgdWXH6ycTOU3i9xLjray0DuoTRHKqIW4v6JlyoJ43oUlmhGepUU
gLdf6/sTeRP3oH2/5I9+7jpSKZGgpkSmTD65yyDFU6sZ5p7CRpgGd9cdn9ai6qJ6l3hrhgkVGeEk
af+Vlu/NYc2VEIYM+5FZDoGWaBdlAutlpuQzGYR01eK6qWPx0NMfxXa1CNrZNVaiSrjJBF3LzWQd
o3z4Q42a726xkLF8cMH7Lw0G7MsqEKXrdC2jGBB+ZtCoSgkQ+kH4WSP+WJNhXEgdv1KMqAfOd9md
/Q0s1m0tUqev5Scbp/6h7/XeTneRiBMdkRhqn76Ttokujm4QX0c6LH5DMM/L2wWs1xuBw9Etv06x
UNqoIk/wRfKkmXrp5SZDTkqWTZQamNfAY3WeH7TIKESVb7gknvWmWg9UKPm05ZrvhP12YpLAoRos
frF712l7ZQGy6aTP/84DwB2iC13vQmCSURjbt8XcUhVfsdlfMGLL/0V90F+OxUYzbINYiIdTuMUa
lKU2nvmHhgx8PIpEqy0g0jy/O9XuG8t2MOi8oA018mXitfs8YUXKpgIiAkkWnXuOCHFuVwZeAHoG
A27s/ER4C2iILk9N9MTYtKF5kKhN/Dz+rx+SVrx4wR3seyK/KXeuu9cFHT1hsK8i8OWCi9TvzxSM
HmiwKYjkChWCvjJDZLkVXocdgAZU2MMCEcrxWV/OC7P3nXFVRucDxyi4kCB3mLXI9mwtMkX4uv97
02468i1UHJuh7gA/xYI6NqaGX7OM6y9Qu2sY2qsVwsJ8MDh+9WYtsRd1xArvgn7UFg2SfctNv0fi
xcSEgJOHTZAoxRnMFtiqYR308q8rFZxFhv+GDv9y4RzH4QeyHkGy6ToHIPd/Pbz3keH48oeyw3T8
3LcCYnJnmKtmQfFQA7Dh0nUuZ5WJJvrNuDyT4eM/JMmF8v5jgV43Z13JXsqH3PCx8n+jrGSIgsXb
07kqJznFEekEz1xraN/xsmiNzIlWpZx8GnQwd4Zh0y4YvS5WZ2ofVTUXDJ8sl0T/Nu4+MogcKUF4
opbr8smeTtVey+lbC8IJ4b0faAs096kwFdobt+HrWaVHXhkOTzyG1xvVOOxm1/TJwssRRBUqcQAB
ADUGtFs/QhwuPAx9HwrX9UAYSacy3pgK/1Ur/oDaioCyvZsZHUCUL/DYe4PrIaCZP2qUMOBZSMuo
GFT3tTBtrzCia6poo/K7wYzif469uOuHm2QedF8HlbU1Yarqjx2xKuQU/WErqbVl9NRhBxtXzvyV
B6siWAqtlaR+9d7Tbp9j9VPy4kCryeqZIzKXCECQjqJLn8lDApT18yRJ10iVsI7QkvAiVh/T/d4V
6RXz+X+xHRYxCjIgkGDfnvJEKtAzxTE/ZC6LA7l08c0Zrl42PerQvO9YDc0aAdsMkJw9PJyF6D9b
JIMa5esUoINx+mF0EoKLYDp9hV0GPnWBUQPYmtaDHlKSKccp4F1PEswVnBZvlvq4wKMeIliSxwbd
gvYFBB5ygd5mVFwC0QrvTGinb/KJS8A78Pv29YMHPFW/HuW8fQBxpOCBI5bXk6aRMOf7mW78Jz4z
j5uzyw8dq22HftieSETxQ5cR41w/80Jggo1owHJ7N8dWvisJXXSKfDCAOdtk71/+OkxARmNRyCau
4JaChZHLHd88f1xKUc3SYtAHD4Yo3x0VbsIHRAq00COm3FGeY2Uj4e9LWLAB/ZZuNqejPAfg6I+6
KEUnzcccfhijSa4fOGswuWiMVmHNA4aYsPcCLipKdyPtzkFA6b+goOmSjOxIEondB40DEIvY3QS1
9rUEM7ETY0weK+KfLHj+KSARKOFjuQj9zbk+DN4MQpZeUEnpmjQt7FITbJM/dTXHEUHVzXcnt/Pe
4ePjUXAhodiUHgJUTrdlcqHoAZdalDaZyCNNcZZ3ADkgXA4Dz3SaBHIxKYop/eKTN42En6xtxuad
5fP319TaGWkd5pHI3zlgbch2KPdw4BBL7tlc+KqOCydEzOId3eVNYbUAeeT0Le7iRsAmMfSwcI5u
t57wSdhmg+Zb+ZZwtS3DBsMbeGsaWjDqyPMBnRq+XfalOxpBormEyLaVXaA7rSwBzzhZMKIzoIds
QxcBgqPuPzmALZMxa+7TFW+2RvI+ilQYpt2ZY8zSHsQhxj73Bt9IZquKyxRBsSj9jgJp15eZhMeo
3XN6p1JRBgVLQN3KZtucgLZzdtJyxWZPAfe/7hqSE7a9R21bQGb9fUTAY7zRVmE4+tZrxCXhsxe/
TwTk3RwwpUI3MOueNj01ZuDnxhI23vGvaKI4HhSs8K6ZrwN+ydRnWurnOtJhef9gsDdrCRHP7+VV
mBMIsWL2c49S1HAOPajVgEIBtBiLaooKUmkgCLXsgA9c8A+aEfTbuYMCxzpRYxF+qSSh1HeKrQio
Y7JoMCnYa9Rg/H7G9kwip9SoBK4HzbQPn8YAiKGnPfBrbKQLprb5bqVMWDBRN/dsWINob67RGhyf
b/oOB9PgZhlt2I3sBiQ8oVyzsQ5YjLwzDIY4H2MmCV91va9Y3s3biwdqa/MrzZrEPxV6WswiKyGG
+tqXjGc6JJ2bJpeWnHXWkQEAx9PzYNAKiN/zQt3HjrVAo2GQB1D7hCFMrs+1Cg/8bKGVNS+41qPH
oyNL+W/UR3Qx1/ce4u+oo7pu+kJSC4G1NHNFLA3b3wbmHILvjaBUGxwz1Auj6G/u6WrTKmWQJM7N
QK5Ugi3GmoZuU57MQqTg00a213XOxrMyNtbFMFzlu/kaylRHfevL+2cfdRoPQvQ6u3zQ52QU4y/f
iqtPhvZBrRtTfpZkDSTt1a0+5knmRbtIpDygG/MOInDnUsaM7LWPfek5N6qNK26NtngqZK38D1rm
wx+qzdriaV+lufD8mxbbolil2UITsQF8nSIawWEjP1LrgQ62GqDiSYmbAMU0j4iKB3RiYtOECo3M
KR99LN2nwCrNbFlOEboNs1tr/0zNnoNffChYo7TkgWEvn4+uLpuuavK5kNTYe18g7R6h/OFavNjv
kSeJdARQI8VKFRdhwpxOjAne+pn4WBDSTHx1QPtctY6r/EOd5MQzod+XzgwWwFCTFS2yDQSsshIO
MgD+CMd6s5xYuu0qdJA6X++ec2MSRdz2orVdQ+p6NbOtQ+oO8RAdggz4g64JoFVtqLRQ89mvBr3u
++Kj+mBxIH23+0C5eSEgcpP8RVeafNxz4qmlkXt0rMr7ol59NTyhEgTbuFiaBCpCdcUVL7mrC42m
haGBiamD9j4WJh0SaJ4444tYuvAkzN1L44lBLVk59YNxnvQXHKmSl6nB2Kdl30vTmZH84OcUHjAE
fIy/uODFLyJBhRxiBJfaWcrbBezf4KyNuXW2UdPD8Y2BpTBAG34Dc2MXOGAe+DP9qLir3UmjYT/i
u5LrUL+Ihi8b9InKeO29ZS2RwuS7e//HPifArJpht01+IdGONkbOhYW9V8zukHcT1WFFuOU5cZEv
a0RlOXTKO0F2mxbHmuf8ehRlNl80sOB4iKMg7d09Qai0byr4PZFmrJr9/yoOQSyd+OcKvUjnsCWa
IZ4f1jFRBVSlm+cKA3uedgiWbVLxVxLPrWX63OnABfT9wq5ztdOMy9GpL++32AjKFufOJb7V5qWr
wH/btDAiPZN3dN87W2tl2fxdXaF5pmsa1z/XE4ASMjklbv+nMS8MSN7BKebjgsDPB/d3HaP9YTP1
+xOy1rCfKFUobZPfhHr7Hbl/1Z16XQk1vBGtUMqY4JjgTkSzqlW6Z1n8D4NwmYNviX2ebsue+KRQ
xc9KtwgHv3r3t+jihW6jNk8maOa9D0T1NQAIa0/bNgiHg/eczA6pRSzsxtwywhTYC9G1K3f4z8HD
b+IYYyGtqTA41d1/kw4sCkpAOvwFVfczq95iK68ADhtq9SNiruKBprBw/8d8tlZAHD8OmFHS3ij7
FLfQDcQ5yJrhdHaSf2D1AoONnm2fyBvCBQNrayZFcGa5Sjuvet0LkJ4Hw68KKntVQZ/JzwbZ1Rhu
Sk2rtxunp5s5lBw1a37C5aL65/nxxL0xDl2lPP++cnJuI/PnvCOXdyLWUU1zMjdnPZesX21ASAEX
CO5nwaolMA51NvSgLx/x4ofAv1NQnL8qWeOQ7dP5l3XZ/rBkKG6nDjZtwjvtbIwtnU+y2Jf0nNOA
IrzkdhG7vUTk58h0QtNj/g/R2dDOMRwm2pAhR4VLdjeSVsbWICsJKqlo0ebnq0CAo3CoVOKsO9Jk
FGPTpAbxkBYOOLeT1v30zxc62au/lbrLZnW17Eg03+6WhNzifaAZ6QyKi1uuTfByO1MbBCVDmFvt
npHV7u/N9zDA6BlnhmxUehGaHJO5GUrCsK45Wz3iGZGymqR16IvGpv2gBaPK1vmN56vgyg8Smfxk
k5gPzhUhO1LkaQHr8hlozA/6SzUGqaXSbg9XfWiCMQYIy7sd/8dbN6SO+4tli8sTBVpFuVDXj1Gl
+/IEIaOs6QkE9gHTh1zUwsYG4JhxUnLWwnujju//cV0exaYz978/L3Jan7i7RlSCCFuwrSL+ZAhL
SmNFz4CPtkqRobqngWVKCorjsrLwuDfl97C8q1Pxp6h8Id4VzjHu2ZT9N8Jhb3U1VN+lM1iKUZBc
Qp9AeWQ0PzfQ8Vh+QXMsHyYX5GGTEq0vDdYjvwzwn8LWj9UXq/IvI5TixU3nA5+/NomsR3JnuOj4
LmCxFqJor+RroMm10IHkAetVcQP8ncJ+Y/7t7A1ahe0+hGS23T3P3MXgaHAKUpWW76sds60BVhij
zliddHkEDX9oqMIxHKP+09hyvA2fETsYFg/sFdQtj/0k/Osaa1PY5NbQOSdgEaUPr4zvQ6kqvR1M
ZIqivniZcLEFXqj+ls+6hrSyO4XzfGCuFsPI/gm9dobPExcQ+EWVh/DRtccRXgopS3Jd/fGhGVvi
juemvVFCIH5fBgLTQ4ZP0vXlcHo2i2YJJNCiMQyCEZyJni+unJ/t8AwmWX4cUketphvVlCiKTSUH
/SJvcTHK40JJwP8uLRFtGJrPAet6XVfJClvQuEJkr5A4HLN8dcc2w2Os4H+PVyDTLZFMnkj2apzm
EL3WpmiBGb2An76t8gAN1G4BIpm9FhEfZzW8ykZ27ywkdxSIVpBjVLkIeSos9j9o3enTasOCAdiG
hBfi//w3tevdufd82xUjj/uDy2ZX7LDPlaTOqwPDRiG4E8fnBxTPvJ34zJl9MRbERny3c6rcEm7L
IjUdXsfCXOXn+sbalCKlnX/PGtqhAJi6Nmj2bc7RRumQqpngNd80Bn8dKxQxoQAc1F+hkpii+wHd
VNntb3KSg7TcZQb2CO4vuhbMvml5JdZoc32nDz9gjXv82e2rbQBGkDrPK3LRmnvZee1M2MC+80CS
fMgkaGPGeGVey8Ui+SGWl+JoO/98ixuRaiFTuzNlkEDrQ0DHR8saO2Np7QS9Gcv9o44RH7kLiBmH
c838mwttEVDT9qm3dIpiLDnoj/Gqkgk2272dTxeIA0xvVXan6T2P3qzdO83H1NgMPTrK3iFKqc2t
pJPO7QjzfimvhXNxrz6Y+iorxRlpt57tWaih20lcPFcQmId7Kiw7A57VwUfg/f8v7HY232wMtxPA
DH1IbH+2GTtQp6Kxas+7ALcVTr2AnwXrS9/Fu3ubO0GqkBlvM/xw4ShVW5a0Bf5L1tuApj7Ift+S
xD09hupPR/gSGQPeJGD2Z/cu9mMxxwLI7rxgra2B4dLbq10JF0JAeLLdXNXZjVzzsXGfmU24JNAv
G71mtp6e7jgwlSE6zCT2iLh6X1pTTbi9IlyqwY0fuY9mpBxLPZ9hpZNc78zlECksT03X+he6ZZl+
JfJ9bibvGvzeAoLp+KcNwX8SfJTSmkHBv1g2BRUEmZd9dZ7fvkGwCoyxg4D/Ap/fBYGiuVA85/4t
W30GmKghsL1HaG3UIhlCY5et5/xesqmEnn35o6LZjG7BlW/XBSXrR5jio7Kyu8eYaDNSgQ2IUt6Y
ghLTwL6Xgn4U1fZrgIQzeqE4Y0XggM+odUzkzU1K2gyv42TkCxlyc+clhHLXSyTQEtbOy7t8ZvYH
/Np8bkCHQnjhnLu9C5FdZAlsuj5HneorjQ0O7XNUyrNvZp/2H1MpPwUsA+j4EnaBHSjaJJwLnd1O
aFcVUa0tM72F/zszdva4GbnUnhXsM+LztwIfIuwz/k8IUdLId2JeNvUKplsjEJ2iGxKz4t55EW0N
FcQVc0H1D0K/Oi29dDYhrh7Ns3K8iv2kBaMxoHngHWMPox6BvHH/cpmiHuVWJQUcAx2YVZ4hMMq9
XXDvlPlX/MeRcg1zDxQkaQ+awWRpDedb5SG6Qmt5hsd7SMomY7vYt59V7EO3nvKswCHtnOqukJXV
I0DUOIQF9wCoWKoyYXqOeQoRNNJ4YhC/umxLVCiApUwA+AoMyO1JU5kbtxNXQnSLKs0/HoBkQQ07
jjlbQJiADG2iXoOWv+0kiAjh0BK7/WcZsTSOE/i5PjO/wcIDr5Lb447bOzqQmDIii+CwX/S0Gh/U
kG5QiMn6Kicq3Fg8i7nsGHOslYXYukwEby/QUiozlV17euRUs3rNYtfX9QS56bnDmgfH7kYPvYzc
SzBs4yn93gB7EDfON/gQZEpBl2Pz8c7657IAlmg6i2Fd2eNNJsBqdrwFeMa1CX0m5WW4LMdtl7Vs
twcMs+2DYL3RA+3e86EvrhcdEVZyVxYf77QkDn9vx/mqiSSq2q1ZQpHVLMgUOpB4mTuiqYiuNYse
dMaTCa2ghaMZPJ9YtN6SMWADhX6zEjDzh4f6g1F3zuCEY4OHgLj1SJ4PVQACSNmsWuZtcP73CJhM
NWz1LEmQlyRJkMIxUJAyt9mfJs0Q39pAhIEwo8PYueCnK+giIdxQFrzoG/A0MPvGT52squzwjV03
T2caMVXgRgzoLZ55RuiASIfFN25N0TD445+uVYca9V/LS/sS5w1CpaaulRD+YDj74GYmWFgh/R/t
JxjmVtyVt6H7xCxGjsu35fMtT4gxSRwkkRAxbgVIT0WGSXZWAAG1huJGt6V22USTkMCUIoDzmx8O
usKaoOJ4Q9mtFeMuIEXE1d2sEhCpwwPdSHZhZXoi1Y/2giQoN/2AgDYBNN532YBGGjRBp8H3sbgj
C0pl+Ra58njJL3VBi0g7JABfkC64722nPvrFvIKgRFCG0bmGBAqnu3q0Ilmhtk+/Tw8XDBXug36R
K1+cNBDQQWXTf/HNEn60bO76vRRkZDt4ZOy47DJVOxYaFyoL2mvt2VFpiwyfxxRr1tAvMizU71BB
uqnm7P91Aykr4eeo5yDItuIQnIOjl2eCuFLQb3Evl5K2QWVReSKzWAmKBpMOu4o8lrBAqerJRHJ+
EKfvU/8jopk75MH5bDlRD9wOgkVVfIQy768ou3TezUGoePH1oQzUiIwI1sQ/ys6zHHbqVpd9BVqV
mS3Hc+K2waGr+/hnHsj5k21tF74O2REzIVtIcMQNtB4O9ASQ5NOLQT5TpIzhjjuFlC6Dpy8/HA+9
A6xQaW04Vw/JBwOEmCcD67twP5M7OXNSWIo3bapdpjsbwvJP+sJbHndTeOecjch6kfdvB9iYSHso
MStnnEQDU7tRgrjqr5jdIKQu+PS0G36vugy/DrHfVXeCKuLZNfqc1KYVJwyCxKgB4l7t1wBUvhoB
y2gOIAk1CMIcj100TeS4CeezYb/CJWKcEuVuMGk1T14DpQFUM6Tet47CWRcDyyS5QnoMDZbKbl3s
pXE29pdif8UypZicfpgS2m1l3HmJHaRLA3rySpGSjBMOUrUfhutykZS+P5QaqbMm5yM5bJGbGfrP
G+YSYKCuEIZ9S+4U85i6dguuscaSpkeLE1q7E0bGbRZp8R4qH0sd0VETK5ibrds32Yvax1M6Uy4c
KsG78/OuQ4Ey/W8NsruViAfviBO8Xe7YhnXqkWO9+FMm6htl4MayCACW7TEb7hsQPsPZ5oz2rKln
aps0E8K4V9bZo0zNknf41xGeNpNKIBiVVyTPBUVojIItoNeitjawS24nE5ONwTnb/0UaBGk5H6SY
Ditszq4SMFXqBlCIFOQusj8E5aYd5dtCnv4vKSbLr/7G/GjdLE4BYa2fTcABwNywG7lvcFOh3+m3
Bp9bMsVCZAJb6sU5ADbptbinBIWfdNeKaKI9UByVmypserGWiDt78dInxVTaD7ILgmSapkOdCmbN
9iiqUAeqDFWaHMAiiyEez/ZHNnIKb7IhZrf2cdk1DMoCwpRs8PDNxJTtQRKCEEZwE98vwcAPwAV/
Ey7wzoknn5IH/+RyUokYy+mubGG6chJwOO3WQvzszze///6FPvgVq5s1gLzCkzNlpIaHDRc+ioBR
2zcxvvo50Yi66DKqtAb81ryYjNS3qmT3uDQTkYpfWTqTi1oyJX2chcEFHBBeC08ERV2ziDq04S4F
kvjnefoR1V4llwlrhJFWwnzf4404tNO3Y8b3AvyljnsMG1gGvrR3wE3HkMrVP2QC68lF9QnvatMN
cn4WLZUeCcK9LrsfJDcOVc6FNh0blcfR9LHauvEugROJyRZCszigJh0Hj8Kfiychrsnc97Nw4r4U
ADQVhJLdleoYElbanvgO82tnm0nLk4nindlMqynVYCOg4HPvr8ow1J2eVy4GIxFhFyXfzQ/YAFff
NOg8/AEc/vwT7kjWT4jA9ktoewmTsKE1p6VGulGQQLJr+IWHebIZ7XtUhKI11Ktkw4K/cPysxaXF
ir+Z3YUvm5Ggys9tq2fadApJYUAGUCbvEO5h6no6Ri2SwvvpxNDApB1EX69cOGOpI5sJ7cLzS+jc
rPTAKZgh1XtOvL1fH9uMmZFuLAnLS4qB8yuctRZ7sTgD5OBPI9fwQ5gGmDkmUPaPA1Th+CTsK27v
VLExitGDa9p25zynlCLBo+61sYQ1s8wng0K3Fv1Ao6FYnpL2nw1ynOA1CKFS4/VqylMid6HOIjAZ
xY0eGTLm4EH33j6oTNpB/wIcCCRzg8uz0wZXP9QfjiPC2e5TjeqiIPEm+5KOtMnEpzgBFlMS5HlS
nf5NC/DBfd5Gj8rDuJuOCwGXgqJJhLQihAsFq4hYXSFa1sXVAdZ5XimIpln3j2xS4UXrMXIV937j
ReKToH1z8n6I1i+NTlJ98exmBLRHflJo37KpaY5O5VN5vYKCXxJRqOqclVi/aywNOyfVSfLjQR3Z
5T7KDigIUGy8gkkFOmQOZHAA62YSsXlZoEroqzXO2Mbanz4Iz84cj/32ka5eBV/lZJ9Pm+s5b2cp
IABsIiRlzR8X+1pThjctfPpZqc3zh9kYPWeKBxuCiK2wE6yF1vcOiqdm+iED2zwwVyZsErPGGtbP
y3x4j4pr/jbZlIXDucEjSdoC3fzL6RcyJWKrMZn2D2UPCkfavrg88TIro/2bDcL4FfP7zHYWg1H6
sAuevsyY8iHJAlWIWCmmAH/qbSFLPMAZ7iYW3QdRXH8xo8rIT3Qho8DLuEE/l0OPNg+1WGLJGxSS
ZMTF/yyf9gEt9JZWjMzuNF3rf1TDgcHq2OZTp+aHA2auKsNTbSTn/JveXHDgArIWG66kHfN6XSPu
hLzuzd3IgA3OEOaIjX3+43aDMu3+nijuoeIpC7CgMYSGKhjQk1lRCi3xX30n/00WNCYalcZ2ZA8C
ZFSUPZ6oGtZd6A0V3rE3r53iENsi32E/qImHNaHBCgTAv8fFtjuMk/eoKLdahfspN89mhFqdyC0n
ecZxkG1WH4IN9yI+nhsY3fkoIgW8Nbth1LwmzrKYq16wnhHkZEzgVrGesE2Zhc03O86+VuRjJs9V
fqg941ypEKSDWc6WtHPL2y74Z25eRxwOtFbPtQHByWGw8GLbyUNwOG6QRtczZwnbi2xyf+uSjEkX
677tKjt7tJzwy6YtN39JAWRMjTIguf8ERRNTcyOPOv2UArCY+ThKkxKU/JpbK6u5In8/hCWZOe9r
442imO1sLwnlIHNMeUdbmXRJVF0UzlxNt8jMLy0O1rakHtDxJvy/6U+UU0+qLJlo7Jl8qyjOM+Dg
QTf/x3v5w8fNxofQuMczRDP/QcFekMKJm543pMWebBgc0h6niAKkPWaYZwlNkkT53ePAs1L6dCJU
iEjsHFKsDMfhAxqQ/a3tl2YvWNgGQnl7QLhSSr6Kp3kFU4VVQ39EfWC4ntGDkqJPTTWYwmAHDck1
1MAJVbUr3Lw2BsGUP+2TFHnKyNeq66I55FQTe3BEiwWz1/7V/ebWsKIWxpk7+9FMdueKeqs8kdbs
j9Mzg02Gdx+o0YZ4J1jayCwkzPWAjfvOzv5C1XsjfToyqSVae8rIPixZmKKp4QXgycvvdeDJr54k
/FWCb3gwj6LeBAnwknjxNU9DtOuxndaeSsdJFFLDF+DMwmX+qwyD0u0mKih8wRF1gZcnjpv5/UUb
5UKx5GOzKAeLBCsJWF+HIHrF1dLd4JO6R3Ou/aLEus3T2+OOhX94ADl9bmywu+ujF9gA8c6yvncR
EkUFhusE8nEa4U2Ee0tztpfif0kMt9xqbvqScSCSbi9/xLuZ2K0PDj4+vHanZy3W4vHnrsQvmXSF
i0Qw6dmUHvvYIehdyg0xf6jdONycOZ7BgljF1PpRFSxEKc1ZcKiZEpGYoHhI992vB9nyg+2J5VjS
z6Wu6x3jdsfL+GDO8Q5Fr7K/rESUwePiZKea7a+9TxwAcmYpcpk3bzEZ5AtM1hDs9YF/MDmA1JiI
SjUKvm5h2iW1JD0uLj5sDUB4jxJ5rvux0OnypZQiI4tfuBU2Qyo4tlOpBA1QUBnc5buXL9uD+U1a
rLMKEgkv74HHRu/Kv6cf288fwFZG0fPfWNjRNi35d3tt3+qa8HPbro0z5FAtFMzGHFlsgdt1e3an
bnkE3YzQwS2trGQGv7AO3oW2qZMFYVDQEssxBWrEFUG/JQVaf8j305po0e7DtBB5at91McA+PUrk
6hmVXNk5fRTa7Ot+XhgzIy5B5pTKEAYfQYFkWm0Js3KzVaJsva9vE2T8OEt+O59fk6JJAY7Kz5Ah
jGyFlKqYvPh51DhQXzj+PUwkrSgfb55ZOPv8SsJDfbhIucfxYt/XQEcZ4xSYixvU7befuNk5K6dk
QfCEjEAXCmtToDPGnkkKdnV12g0SQx0DrnmbpZji7W8W74jWmHNWV4G2JDvb5KA+PB5UvWqqdU/D
C8+g97aTCTiP6tIEYjeC3CChQk9KeGUSYsVNLthZKYD19SFYlcuuZ3QNYqiwCDsLmbwkBAjYca3I
0zNO4nBwHAuQU4o106VF3QGlMY1nl+m7LPwljJ4/feTlBE0q/WgEOIUs4FLonpL1ubxhXd/61QFm
99B235J0XksVOOp8P3fyaSeGoijjut9xUu1du1JAZIiQUXxehlnpkbZJKDkMSgTGlwV4Sj0USfeO
qsCjXTb984+MPwFh/65WvhlSM76/Y/xgA2Zj9s3ZzInvWg801CeGyMIbkZRwBc1wevVKM+nt+rxt
GHoWc8dmbmChQETw8uvOsHalrLcj3hr2hG1tsB2Q6c1ZCvZlOXT+XUufzZ+iYdsoAb0gGC809HaI
JroGYJQ79Xo1XBGH3f5M9onthnJvK4OtO656E+zbodJuI68n39Y2XyieLlVnSNy+FeqYcQTJl7wY
QGwHGe+lo0uy9CRKViiVNt/1bTW0z3yyQRG/tSMW5qNYlbh21JKu5euqqUSRUvbMyWU9eaWBvRnq
0qOdesTT+cjpXa/uWAyJDHAsLzsbz0Me2eQWWAmcd1TCGsrffl/7gpvXo+JhN1gsFmn7mWbV/IFA
PDK9EpnXIbddI0F+zv6l4gzWSjzRa88Dv/SXTG5EVgt4kIpFpr1BSflxLxuzyKo6fNkq6uRJgD+0
oEv2guFYM6yvSC8aj5gp9SmDFBF7saGi6RZx58lt8Wnp/ggL1DVlqBQHB/jKEXtXKKYsPGnuD14L
GoQCSO0B7lULXORYmg3H+ZQcsaS3fvUPWxgE9n/wiizsSgDAKwktUiNYMtSuO5AFX9/3xcaiy2dU
PVKJIBzbTmimvF343AHZYggkyrjCMzgGCyne0T+soSdp0mQBurZxoX4EDvyFnpTptIImrYLEZftJ
PG6gTnt8z8jGscU1n4NYskKT89oSt5CR/bk4tPXcecmH22nYDXmFFdgDJkobq2c6XKRXxYYvYf3F
VzWqMsH5li2C1/KWoO5X5HonqoQa8QRL6QSDCoSUGBKAdXftOzEamFmAjiqfd0Lc5VNFxA9OL4R+
FRvFudRWB7xP6TBBjZhbjM7OZW2EhDehn6lp0b9F99YbQK8oLWk3NOMFNDDhvSQtW80fESF0tSAz
w8+9CM447cyikFOgeyVFsDJNljsupgg5uAeIRpzxt/CylPozGn2N8yT3XfFtPKM30eHfprdTtosK
64d79+Njo2hUzmnfs2Y3qVt4tgNZHPstTJBA2uSGeTRlS/b5kqXY6FCq7HHGF45eubLfxRxYzMJC
qCWUcieEPF044oa7SdxzfP1j9B+92qXEw6J0WoUFXoCxw7vJ/bDy6K9Qgn/1XcdzTFfCvMbWB8rl
OvMqdvBC/562voIzEid1COyMYjyNQnZedhbt6x8gBSbDSXJ9OsyxOcFt1Recn/6HS9VYCqp9mgjc
YUPIDluli5X7mW/8LebcI5NL1s6Cd+qoKZnCLjjW4iE0r+rX9OefAbfeO55p0dLmXqmxHyA84578
6MVjB2AAV9aLS4Z+pwywZAuM/Ercu/d9arCQvhYFtayx1igtwUBWORHkOyxCN+/xaFKg+FlH6gnP
hCiYmZ1ej5mEeMM5+aGVSBHaMrignPL25X6F4W+mWrpKM6AOcZiomLct/qp/TuNcw8hknC5p+qgp
oa3e5/KTl5/V07pW3Y4I4dpa2fPgOKSqdOFGeiuq+leOpnj9HJzdVbeNLriMJtk4TGuveFfmQKLT
xtEuEMOV0umQJXSOCZp0NUwjXXBTagxYvWPre2tX9abX3DFcf9pGp4OsIMJYtUdvJAmXkKIEZXTR
0DLO/6B+/uJQi2UXRVesomQnnq10jSVPR0MlnqSYGTeqzFJXtJqnym1Sr+ThXIhR8quc35ghPEwu
XBIq2LKhVQpvII0t/cF9je6qHqFJpi7JKo0HbOkW0vL1BLJLUz9sgcAGu0hmlHw6f10VoCcoVPaR
I2qvPv4dGt15vb/aJXKYVyO3UI11AGgE26POAjfEh4H74L+bsxDGYuCUN11WEUFQjPQgQiSHaZB9
tfD5brePt1yaDxbS29ZIhJ8169h//1mryvy0q+cGDVc/d/VGKe4GPY0M6jdEdiCgbtN1f9qj3PkG
6dudazUpul1tYBkiRj0JQJ6Qz6e01DpYzgcyyuFWqHb3tx+TTV9YnWqVvRaQB6zc4uuh0/4hP+p9
oR8pJ95iiIztnSB60LqXD0sfiI6n9p+ch+1q5kYk62TfsNiMRICgY42MnCsDSTM31GHSxhVaDPPk
T7R4ve+bniUzcTH9JjutHDh1KxuP20g/ZgxcMFzl0+q2ExVs9wCIKPwZ4TeVXLeif6jOy4JczQRL
VKhbeOOQcxuDFxaSF4zX5e/1m61KHQJ/N2290uOuGaVUQ1AuxDmjg2mjLee6RqBf168LduycGnfS
nh3hb0wOp+42zzy4yyucO9nTW6VmyVgcEmq58fUMaNzlX4WTWzhQWoDr3YE1heJ4/MAPp5mPW4gR
hOaQTnbOfc48vAetvjE5aH6KZBPRU584JTXgDbaLD/CYaBizlvFQWUz7cTyBTdVL89n7p3JnODq2
T3ciOWnVG+dLdocqInD3gRvhKzH5zAK3NI0EOh6J3kZWxmEq87YXmxgRxv6TT19S13DKnKI46/KX
ftMNx1mTUg1hf0jk37HMzKAEJK8hFzUMLt0WHy6sIc/xmWs7TC+NAXyTbEEEmjVSlw4tSh5zcskx
e17YAgjAnx7m9uSKcIUQpz/5mTRHRhQwieyPHADcZx+Yh7O2M1RZgG92zQ9jZMlPK+lphvAY4Xh7
XzXoxmvfvGKjI7XygY7ezzgsfqcvzzR0rFg8ukJQao0OmDWCuSsK2Nqd41/7WXQITJcBPHpeO1Re
MMtGQ/hrdGxGC517K2J8caoEyVc/DaeZYNfUV11FQ/BqQf4Zvk/buE7dDTXsPPlRGU2Y/x6i9+QH
rpG/VfiIoHU680NfKR8rMdBM6YsXaxR94deE2aS9VlYx7sDGajb13MFns4hiHBinCpd7TRi/bt1W
m0rOeSapdzqjn8V4wGX+MIOCIccDOioju9MQhyT8w6PupT8mdshmJXJZPuXK73Yh5ZIsCRpK8e1K
MIcqtlBjiDg9KshM7pwAGW7D75lqwVg2PGnZXIhPxVF6gNVE4PIlqB2SIAvzdoo4oLzl8GA0umXc
+beljVQp0lbhZzgfKQPU9sNoQbeF6o27zSGWWCm/jKMvJHihS3Q2cDkmK98GIOMweSGSPq/VtVlL
xxVQL8RtMHI3Zzgw/U9K377j4wpDGWELOY4SpgxJf2G0vbD96yBjcw+dA8tZbxF26/2l6YHz3NkB
c2DgSCIqObYzapqZeoBBlxIrbbcSUU4DbYS3eIWWk+X1hicKPJea03qsWIGme2KKWdom4+b2Qs+D
ijF9d34PfZwIt1oY3G/elVu+1OjNK0wpW88gfGglSrlOuokWl5TqNVdsLcL5PBZgbNXZv2MoyUzB
nLsNGLm181rWOnz9HEpdGMYQfhcllDwZf9uGmn9ATT6TNh2GBE8SdWuWpofMG3hP0tb/iFijp2+h
8QrWESnXRR/WoEqqTDiwk3h7TR1nd/xnui0r0XHNdyZC4JPFCIXXGsLfe0vcRwyWOn/ySbM2HLka
LXwlzvsIxLLGIDkmC+zq0yCZo1vURhmlrPLjrQjDxDgYrmtHbguA23N0JgaFbRq7XLLzFw+vD+cc
QDsAp5f4KNcKKqBLlQA7WDTr+z/PA7kobqTCyawvlvrj0B4B8NegGtU9e6RLLXFvYt+2v6GzWfKS
Oy+YTxnEBHTjvKMnU8JGaGl3S9kImzbrk6VIONi5zXI98D1vMUICEkdLp6EMp9wj9zPqNe+GpCkw
98rRwVc4lVetpJvnU9/IhFWjlmKmA3x8F79M0VchlEQt+USkgfqrWuoqmkk70K4v2lhrH64gPKhm
mn18peQq1A4wFLFgsoytWqllMTy4ySVXyw2pcAYMA2JZxr+USFpkjX5ZwkD4J0+lX+nJjZNkWjWc
sB/duC5jsDPp4gAo22XbtFexLHQw/CwY77z5+Rzx5r4r25jX1iLs2SwTGd8YihiCDUI3yKmjyKCS
lZhylYr3kItdtpQj8kEDBBLOpHblRymYgwvRLTDG2S7F2trVYKOIDcBP0fb7u4lCxygXRBJ0LQa2
D88gm5HM1CK8u5Fh+cyW248Wyp70kLNvJF/6V3KV/byIaGHYqyNW/sz8lshPlEW9YoFjjeLct+PT
420kiV0NwCTdlw4malC968wwPUWtIsfRESWYKmw1Mb8tyT0niFso3PevfSGzyrqNeLhz4L9pcFvm
mKrwNjPx9kyQgNJ6e/55x2iY/lRQLtVoDc+OBcrM3oLd/0ixFjhQw0SgbOlwV8aUD5FCcY6A8MZh
3Vpo017pUSVgK4cYciEd3H0/EN74NcIWtITUuAkB7LJ5zc+VCRxPdyY39zCr5c0gC303hMZmgcg3
6RdeGcIYI1T+dDw/nhMUNqI12sZcMUdZGmB4k5RBluwYovHT92boKLt2hoZ5CQyBSLsLUrOk4Xyc
C79pC8gdeW0+sGDPqkqEVUOCMXYR0gInH0TD179yqqnK7uNYcoNYP4MzEdSwu4+DyDr1i264ACWE
/W1ruiwd4onI4f4ZF4sROJ+5PUxMZZnAs1xScuxHf334GGa136sHcVaieW5Q6S+XVEXxGtUh/goO
+OgNckdL2/YBlM8emvHBG6YmQiOny2FrolkMRXEPD9VTDY39Yq0i3ckjm/ecrmOi64gKHPIoJejt
B2H0WWrQ+5U118rHShuOdOf8zDNxkmnhLmbIThwqybwZu4uTE9mb2mCnIIyCxf48XiIBK16HKruT
Wsmcb/lRluvrCAu2BFrC4WuJFBa4KHUN3VNOP05ZpUdXgvh+ZnEqO5GLX4S3Hv8OW+OKfB3j/tCH
cWtJlqeOqgEY1pd8lS10/bJ3x9LDYmtT3rX1+q0qr3FXcu4AY0hUCmI3Pzjbd16Zm5/fyhkZPmzG
nDsXXsgjs8v7zz4NB5WeYwg9fwDFxiE73zsnl+XKH3yj3UOZ1YyEO8qMJI/BBq1J0Fyh+H2FeKLB
ejgvGK8S2FmvsPJym+DYTvQu2Vm9kq+bTqINoQhlP2fZk8zXYlKx60Jk3k6gy/LSfCmhwi3hCXFW
bP4dJsBD32hIoDRCnMBgzyOYaFtIfnc2tl+Kr3uZOPGTMJzeiUL78NDlLTE/V7it6awuq3kf7vxH
PGmn7Ylx70m0LDpEru8529IZ+tqX5EfRL+UKphddrSCdFcDlHopIQBE1UHQTOe3v2Dn8q/e5CcDo
/GS7gX5B57nsvjvTaLV3DgPZoCP1rm9ufbNFq6YC8TUe/YO2Qrv49r3FnPvBdrbTdgeSn8N4HntX
O9l7e3iRie6UwYtNpbM+/49KEvXslNjUKd519eGyZKGgy41K1+WMQE923tTw6PyzCVXCMMreWudE
t3esQn7XvjtHkx3ZWj4GzjWYFojkTC6HITsGLv6/Y+PQl7IMoWmtSOly8QUgsIv9OsFPmhziBqPv
AXfA8KluLaiZ/mI8TveBfntkx9G3MZ0vBwokLIi89YVo5SYaQIUnLS4F+NCORCarNXd4FZrCSzDL
VQVw6hBMkD68zJhvAO8TMNgpj1L01VHBjAWELFbbLCRmqQDaP8apZrNHmDpUvGqUKulhm57tQDoj
2saQvxs0POP6wRz5lifn2iWX2EsCLiaB03N0x58JLpt8pEZCESBcJADkLlOdM9iEg9A+1xo4J/A5
gZBaFaNrjTtCJmx9UCMy6kGbyNfpCFKatZeB0oa+WEIYm7l0MN4spK5AwzW0QT75vNqvbM9S3IEd
0m0zO5jrj44rT7DvfVMxenkNWpITqpsQq7dqqMeXiB2CHycaw4WrHfUegdnd4OEwyfjny9JNGleV
7IIChKgffn4sjNvGO7Hl7QUHREp9nW6WoriGGQB0XjYrohdggXXUB0NZoxYK+ma+dn/7N88N07v9
NccQeIGnyLHyKEZhClmCqjszqCvzps23Hkw+vETsr6kWOXL6D31gIKIWbxbrm12ciddiq9tPvEtw
PkyrHVAMss891I2QvNXQAzU8qrCwRo9WyVCNkFGhWuRec1b0vc+GPvxinAhaafsVEsszAoHsgrcE
7mw3UpaSR859m6o7ALMzvCVTHBCPK3ub59lMbaaz6etcxAAcw0fVShsyBz4JGAxd5YiWtPQ+SxI3
1o+vPk6A3B/5UQbe9eK+sftDXql6W+FEhb+k1hiwoBgWe+fJzqgzFlixItfoaiLVR6S3qTDJCRUV
dZFRDnEqattYobdCV2+tsx6SR9pwbY7f6+b3KQtpj87c0bMnF3cxYhnAX4lCg6AN8Q7OzhZuei+b
lGin0Lk0DE8tYPV4pqAE6tOgUAxJY03BxMfkNdXVi+sJftz3A5FSByJ9c543b2dj6F+uChGZSyqH
GweDIIPdfN2FqahlP81azzz+QcDKhV4JmKbJC+6XTkf/Mc3WXz3ikgyhl7JYZ9lsIJRgMsCT/HmI
yrpdTtRrV9w9L8dYCREEdvB7oRatSbpiwc6o9UddYLqN1pMoQ2vvM8d2Jkyb+k5O8DP2Hrd5U+7E
NBwulqlTDSB9T8LRdcgDZT8g2dhLzCUsnoS41XhwwBZDljTR1gKfQOADg81MtuTiD3T3Kd6OtRH6
Bkwd5QzEkDJOxQNQmSOCMg6q7Ot3igCwom+qT4EVBEBbOSOwEn6fqhiTGzmF+Ak5EWJW7RIt6dtA
81lafAK25yoykOnGBfKz6xb+gLKPpo8xlNjUcuk7DaT5vzeHSZcjmNuHGco6cTvuBDHB9Lf8qbf8
SawJ47+F4KTXpv/rh9dyyMUXJeISUMwEnhlIrfgIgqmQjx++o5LdYhXAJlJVEl3T9aSo+iJxt2bq
mYo3DuSWsdDBrOqWrtBwOuJOL5WdoAtzF7KSJcr/nO/37xlprM/ahy3m5PU2Y3rnDUChJ5px/iTm
bcnVf437h8Ce4GdevMhMUtH7L8rmV3T+22G0nQhMa5UOQ4YF7rcdNVtfsQrMxJFEVopgtE8BiS5t
wuxugHDkCYQ778xtWgGOh3aC90KF7w6U6evOEni7B0hNlklCi/AnZfXZvesGQObVcxQhXQ0maBG7
z0zunx9WGyc4aGqoJ2EIu9rTfhMLWv8PBrgD/hj7uAhT3bbjol2TSIZMZtZIjDeaPF9rD4QJH+WC
ceGx1068/is/XnXhw7L2OWZHeK6FeeV3orb2XhMRFnZN4Wsrki0wIl6Z+8MdoEV3hD+i7rbBIInH
Wy4kAA06Haf1OPY2UXUVg5E9MkulCS455j3NMy0zS77h+Tdsv/ulBXBA5/XcQGnpk2TakUSBF0Ag
v1B/oJJcqJMUpfVeaU/kOGsgKHjF9+UCPQ5HT/QpiDcygPION+4cG5VjOc50QokTfZdvR3VJveQ5
GOLMNGWbLfvV5g89ojhJ24mzVJoH4DfqAKh/2shLr34S9uCMMF9ALQqF7z0QISx0Zfdr4SPRpgGQ
22WWGp6pt5yZp8BjMJcmTDkH8Z/ronijrACk5Q+lpsX9imf4QhTw01pFSDk0xpOxNjpxM9X9VD4f
y54JwcteD0PcM3Sbyvwr3VleJ2t3tn/Gv4Ret6vyYmuK9CvWvbMd9wSB7upgz8s7AMBBPDFsOA/e
3nxaURdsKgks0DTIkEy7SrtVFMU0BAjBaTkmJGhg11U2ynWDUQSrGoU4hnRgBtG38V8uyHHBKOFf
XzQsipixNx+sowMXVWmRkYewRzr+s2elJFNm5UMagqjZ/fDkN6XoH8Jmr+zrwe5lgV+eBVVMHVGV
9D2j5MJbQkIhlrAvH/sA01NxP//a9DtJtYH4t7ZzAYW8lk1Gsb37q7c73CC0XualkLzqCWyInHgw
7g2R/xFivS7+Cbsk3y8NysTuXjC+ChWMBAufa1Vwix7U2dCLKiKCTYajtuNkEBFxkPDsXjwnN3aR
V7ofdd7tF3r958R8f/JMP7a0yIF6N+FW9bOD3I8d6lR8JZ9FAOBWB1G29f5a/tZYXnkNgHlT1hgU
ObIEtqhUu+3hiXDsR1ahk5Hd0RHA4AAlS/fLs/AGDM8xH6auxy2P85zhvymtzx1vxdFTMUxk25wA
Im9wO6NPImFp8M+FUO0gEC5H/8JqeUWtofn5iLexvOVh0ulomJrVWCBa28PrBmjbcVk8iu5QamyT
dTM2N3Q9x78oq0VpW3SCPOpl0hAwyCmpft4SKT9oVcPC0S8XvisjvkjZnxlTZKYZS6NfcN266QKO
omSRU+vsIY+I8oEXfIgXnfphDsnvaEK7k9wuz0QowqOnPMntinXuI10kvAr8Gpe5ZPNU+6CchoAy
hgbBXMwW8xLCXcSD6XQWYM5DmAMnrfmdZz+OeRBvS1dcZ1PWijDda89eGjQzOQAJg1wrrzP/tFGa
nnxA5pa9fC5EEVYnyxw0JNiFdS4gC5QjiN+mjQDda0Z0/ckdO2idjNi+F33FoljOnisKFt3nTnRh
f8HJOgseIZQGKhq0whTdtbZSWWs0cZQjicuhf5B7KQxri1DT/PgD9i7XOpczHsrHBwlEKtGxmBd5
k8JYCMO3NDl8XCuE/SpiZMyKp3s+I03Q0d7FOmrR3jK4NOAOrbSKRCp/OqhCdPRzkM9ErECPGG5q
es416RRRlT3B1L8dmaU2Yh/+htCWE0Wel4Z1hSV1ZWZwc/5S5G3JTY2OV1b9BWzkUdwtQP5/OM6W
BroYBB7FOE194KByrsNwbbCxlVLh1O1kqwkUDPWgO3p2LTkvLQwYwzhbgrgAJ0cA9NYHw178gxNp
xnoezJbVUdBbOmpAw/6iRk10nv9KEsoG324EbMidfe53ZPiwhgIJ+QyvUUP2A1P/g3ssgB0mtKOf
6lq5VKua3YqUrR0Ac3jq0mt/k+Na7k/QB+r0PyEdVKZvGmxzcTZA8F3bxo0MgmRe67G4LxxrRgoi
/fpUE89uMIq7kvdVbHW+1eHF7uBarRcWvubwVlzneTfVA+mwFnC+WFL5a28FXTgsSnYPRa86WeLN
r30IT5rB+q2VOsIwOlNMr8lOefhO2U9QiNiVOprAg0y8Gq8TXcdvXUpspqqCsQysiQvY/5B8vvBl
72jIy0zntDp7RX9XPUB9r1EkN5xSMWOf5Tuh/lLWHCMMoZqrQ9zkNb/CywR4K0n12cUs1MU+ct/D
lpm8XrTb3+W9Xm99Sxp7tCuvJdznZXjc9g+qXISx4tekqWDpEKj+2muwjKwpVO5upUlP5MT7t6ub
8ng7pYhjJCXzA47Lnf1P+vuI27nIWBHNdlEbPbOrp3+lXNXYwl98mA/xmItZf/B0bWsY4G7MBN9d
wK0Ye1syivDXrNI/VyoAXBFtewhGSBEo/ohNlcDU4Vw/vOXqOAauUANIRD5U6OyzGsY3Cfwk51Be
jiOOCL3TJG+akZIyDrBErkV39x4UCuVhr8/T1JX3naVxEojyXmZ6Oc41vRPR9NLJLQfwo8qLnkQ4
k4cIfbu64Vt6bjYBbbFUJsx66xtpFy5FPo4NFX3lCXKW5Ov6E7i0QXO7CDqA43ekKyYXTod9Qnbp
Yn68msRIga2oLHnpT7i2hy/fgCAwaSGu8loDi/X1VkfKuW7sr6oR1ekrMvZAXIyntLpGBkWPeOX5
kz/woQAKA0QKWge2JItlh5S9VHvIRABe3o0Jf0EjrCKbg8YkvuVjoaun0iQmsG15LU3aCqmQI7fC
LEA+IffESy4/YsZjgJS0RxsoBLPLLjvzbKx1zsjKqkJUMTwLcR6QSPeIAc7xy1A0Gnaht1rDC0Up
hSNVbLACa2QLK4BAJeC7CB8bNaRldejeJoOTGeM5UcgY9ED0PUhWeaBhrGpNZegwu9QiSTs3jw/f
zQlXViB8hxIgDKfQYpLINRwcIXJp2xQ+oUR9AKvs0LEacAEaW32bHS6ufYaIGSiNxZdnt7uuTZua
T1fZo3QL61/aS0LrIaCrWVpcZaw2WipTkBbaz31WTDBd3+baSW4lXUgicYEYm/PNQngZx76+WOxl
rjN8T1wNZkKZ2AHQNKjNrlLZ1AtSfLBT8ANsJib7qmnbTnkC3ucMq701O1FE5v6NL88NrihMmYcs
Evvz/viyRgKkHJicmiKrKfoKHmrqT3Swyhu6FjOnH4wsdpu72iZOIppePZxDEoOnPduq0PFVjdQQ
KmtrWJCaM9UzRCnbu+5AvrGZBUbReUw5FsTv45oZR39mAhHuYfKYqQRbOR8+IFhCvTu7xfplLo96
wNTL3wknaR6qVEOjP8pfAl5QPOo9k9i/n6Y4JgKchH1dIbvMgmaZ8K3QQl7mX8qh8PL+pqE4fm+m
Q3m4OB+zoguMc8bdo+bHvZqWqO7Jl3FQDWtOFm3lsk9SuGXv87dAl/EGzon/W8gvh748YRq/qvrv
bg/U+CbyPf1KESlZiPrm/qc+myTzqKmz3OxJQXjX4Gl7H20cbF3pazdCNPOAYtM6vx+eAYoEMU6N
mgit4hWrj5vXSAQCEfqxG2+xqSguk6t7OFJ3nysXaqQzfL6c8Vj6q5gY/I3IZPnvkicEpZ2eiR+p
/8koe3ar2ckiiiyyPP2y/o9Wrd7JY+El+Wt9kBTEnmyZ+tmnV3jS/qtCn60YT/VRWgdObWPbC0wU
1Yzy5chRT73mr2C2H2uo+AqR7m7ADxbNZxAhA/NZzjP5OtJ2ig3Vz5W/Ezc00qGOaanMLEdCb2nZ
2YbNYLt1PIC9CDSzeoS/SPOdbbShNsiqBctryEx21irSPsq0OANtuic4kyynzlbIWOQXWwzBJAA2
z8Ug/pJ4DuexTCTrsKMEs6koXf/9qCr2i8fulbkXlaVoto0plKPKWgNbdoKwnI6s1gCPeP1fSVGU
TESYpYgKK5S39wQ0IQDHbaPfozUVWHbDbl2WbZZf0MdMpMbkPENojjAWsc5TmmEccuAqsjz7uS9a
sW3SHcvdia8UAPNpw8iXPkMjk/h+zCiUmAO9JqjOmo8I0N5mf50rsxe6Zd0oO01oCb+nRDchkXq+
/IOm5uEPKmHTVS8xbuT7sLwkaYAtvNA72NEPqhq9bV5bxHB8Cx8F7R90RRE0uPDNk/9BZQibe/Dj
ygEHkE2QMyvUyyPac9KsoDX6j0/pkhqy5cyPCFespycr+QYE2VRwSjLKIyLz4NjFbu4sx1bEuyqM
NWIdzhtADnRZqWsucXhmiMcM1CPWK//blq6HOJboFbp3aWEbwWYkPnjdlMGrmnk3tZFsuTOepgJR
llE3StMjxVE7dTF1rwrMFa7jFHmEbpV5hsXOFW8DJ24koTtgHqeuBlBQl7Idi1GnQyivVyLPaHeG
iT2DRaureq6UPA15/qzO/59LjFBfOB4nHAIJwY+pmBb8ZvlMfbP+X2W+Osgeu4WReZF4n31nTQ3s
EjxWaNo0ZOUP+aBy3PzvFxspbJlIrPLzZjpVRmz7zUXFTUwYamo59rSEyMUxlhN+W6wxEC0wn7SV
wALGcXa9UqYpGFcfFukQMhZpNW8v8sVOhtzP0yGyusAWP8AF2C8a7NyrodXclLna3iAf8Lp3rT2F
uKCuCIcwBWw131Wt+GrTO2G+V8GAGVvJVLbTXYcBxbqXgPjRoA04WARpoNFDivfGYS9Y7bQOi6XB
9J/vb3rt8OOP0SMs1i7hitUEdNao/vMpzd+BRUAZveFpJUWar40eapUYUwLeFJzJZCFbGvzT67qR
XIS/k54ys4LHz5P09dNGjACzrFSulkpqMwgHXNeVN0ZmreKaYCnC6iUeQWCm6k4rKVI4+wV4w+Bx
p+Whk9XZTU9/fHcI+hakSLJXEO6dsxsUUnPv1uaf9xEs2S58auXjvquBegUBGxsJ3fP/fD/hyc3D
7iDplS8njgIL8CeYqd13IiYK+zfUvOB4QqTAwr7OapvDeQktzjo52SX/dtxURo/LTF80fUDZI1Tn
v71GbmhGyCriY4XvdrQFmXvai1cLNB9SIvT3xFNG0cDjciB8L9L0FJPWUmd92UvK00KiSSK9TyjP
r5C8KcXs4SPK0igRCiyynSDWiX7ykNnUnUdznjlk7214HOzUxzgnpeMapLeK4m0uReqJfvqIRF7U
tkFZub6Hyl0btQEg05z8iFqS1meL6jRZPnDd57In/qbvr1BsyDh/+tB00ObP1dSP/r4jcHQ6rAgJ
P9EJdRvhZcKVMtGw9CsMfAvujWkEg93YGE5zQqvJVKiFWZ+EwfeRKIzCtA7uHnQTD8NhHxojyGSI
UGfC2xMY7zPBIM+mHlsOmsj7lFJpVHKurtr3oviSWLW9A1eG7f+vfJ6bVAVqmESDKsADGHA+LN7X
W9oNOQAzvltqpEmHBHTI344kiuCKnbdlzCzfXMzg510Vnk8NHjkNnD5KDc4aGma0Ae8qC2MbcqeS
HGK1VeH+ejTMym6qKYtdE74aYLXz0+T6Fo0dQxIRp0aV5Pibkfhqt2PlSQZyk676cSZ9XVgaPGur
ZJ+xKMqI7T2jtVnlyrqjMhWXVGFmxKn6fuZBmbTqMKneXjuUjnv2OpkEmGWowEqFJCvfJhBRJ4ff
mdXHG79JjMea8B32EPeFSzERXzoHnik1/12XyiMSxXZXOaeMVWBUPImPzQotz+C2rwaZrT4W+M2b
7XlovhcZPBv/OC43UnRLyO7VZDnizIWDTXylYQ+VP3K9ig/4V+bXnGmw3ZndglcR8prNQk5nnXyE
JfjWHbTZr4K9bfuPDTk/xA0TTzLdVo5onIU18R29+smRFOp+ON2UvLYrW7zefajjf2r/0b7yKwLB
e4Bh0RfcpXaYs7Y6sU+LcHbj8NoHfbSTkd5o118NfbVy7ZAAsALgUCKfk+xue3uxa7XYG4m5UcTr
hFWrXjSD02NeFog7a9AeDx/7W/a5XyGcaEMTjy8rwFYMZLYvuY2rhqkK82/2NnP9lsZKvyBjdYvR
/aQDfIES0bAFxqC/wy8dKLZ+oXTXh9zTCHuODdFtaroHepX9Fz/RhYI374XYpPv8AyTKb+KQiWnV
mUel89Qqt/Q8pbwBoPrzZSrejoP1zoxGxD8/yvmJDqGGL0Vsv3WImuTdYlsJKTLzghe9f2YaUISF
I7hWIzlu2SBpLTaobkHJPeWLxFotCnNGigd5zHykTVeP6B5xVtDoRxwkbJNNL14HZLKjzohGSaBt
1LRnjKIpv44XFpwd2UbvRvba0QRO+i6mn3rwAGhJobq8Stu9F9GLBKs0hAdlRYjGwSdUQixRq6ex
iefldGMpdEiOwXWGfGufYnOif8gnu7qDFl0doPUHg7UelOqVtjE24qbobyjrAWxv9LFZngRZLszd
bNeAzfXbW8uROajbh4M9WgABE2zV7fmpUUrlkNaWnVxnU3n5yZqQkGuc6cJ3Dun9lyfGGaypadPS
iNGuP1PFFWOIV6JoVqtnwTqd7WM/vS47N38a6s3tHbBGWD3dLyKf3TqaGjnNvUAlqa/HdLO6226G
JjE+0m790rt5CI+8EvrhYMaTHyT6fb6z9yjjLhf9NMlgKwEnJM3lJcQWCskBMVe08GE4MFVz6yWI
zPq0GWJOnFYm8Z2074oRfqcnuhl38wdMNKOIzjRtCgBmQ5w6qxKNX4E9q4xVI9JncOElHYtQ5e1/
cnq7Ju7R8+vGRJY1Wyo+HskXmFJpm9J/oMs7Oweh8mHX78C+wbWX8dM/syZ8COOCOGZL7hSkzF8Y
W6x6LVaVPLX+KI1ZubtiielQ2qBdckpMomH8QRBzvca3akcHQikNpq4kbs8f3IuUn0JJa2IvexFp
YFAs/zNL+rJe4IdD/nGJz91mZcLP4D9C9s06um+XglLuQSEJ+eaL7AD0SfgL6gDSwpI9l2y4AMAc
CgxALhu/aTNhwrfOwpd4AlQCOKtNgVlgy/Sl3l4PZtcezzTZdBtXsiI4Odq8I2JFEJJSrYphhg95
yEGZqvk9U3ArzIPjs8TFpHj6nSz8XvRzsFliK1hCC5x0psyWpSfLhshk01wSTxwc1uS339pOcTlB
jxK/c+1chC5IGHzPvwVUcpaNArZjhFqIGYf9nLZFVhopvYSWiPssDJ+54gR6UiZ+x0fscQ/k8Dip
bYc3Pm3yOYNnDpjosEn08yzyciJNkJYIrbjSLqQkaQcoNvw1sJVihvdnD6JuWegmQ3bCN680kQdn
lwcbNifMUi3s+2lvcsfCh5uRhSqKd5N9Yl8dNbXH5pciBibKIzZM3ntsWudwtbPaEDTlKBGJUNTx
E22DzXM2v6/u1yZkld/X2KlcRWK6pcfZyksVEQJiaa0eHw8Dm+NP1EhptUHI8Ce6ybqgiToc+CwK
fyXpDI7iHNUSbdpbblCrOfRrB0Z8XtybYh66n3JgYTpn+kchE4PYmFUvh7z3R1lpgjWptzAOOcLp
hCAjmXIHwSYKPpF/K1i6nqwVcpt8+5T58kfudyfmOVPTlbX3EXoSFIDwaxCWoc0dIwsniOnaH8rN
uX8E5s7lwE+cJCj8CC7CZI717YxqobAUl3T0dE2aBPLqWaOa+SIyZEGqE6j2DOIJjWTn1nw0GV1w
8AvyJb9RExI7nkgzjGPbKKZESwyrSxK44tTSPNod70UvC3qlW+5DL4Cord3mLsS8l5GP4FkE84EH
+cYou4sf47mo9cMFVEZgcpULNSvVf6frP925GuW8dbpq5jO5nfX11oR5YTriZ2fAx/Rv5wT/ey9o
vApZaEonQzpRM95GuqsWLmVqJ9oO+JDHXik3vAdNO8Yxmpg7S3jFMUPZ2I6CyxyeYlQuEcrMs8Ib
RxEZ6xthY1IUPz30/wkEso07ql/EPpKECKY+kY8MfcOnm4swt1l/uCAJuzIsEJUPFeZhSr1xy+vL
N1/aZIQfluK9addSU/yszK84rCh+v/FGVy33LnWujbqEvMoCXghholfdun8JqBUWqEDArFr1YxSg
53hsvyWfK8iBb3RL+OQuvPFyhvQ2PMPZO7hOSy638/8Y3BmNCuVkP3rWbQkSqJL5F56SdWf1gLQc
Fi1+l5ppEnUk9fAP8FHweFvGtNGCM2gPI81p5bBXmq3ESulWuqpUznXHeiXRBnBsrw7cV2nNPe32
5u8et2fiWhizdYl5L2VaTyDydDTww1XfkbcbhS3rbC4xQB8aaRtiHT+V/ZW+xQSyk9FupIkm1rtM
VzK5Ugs2f987bd60vBQ3estmkg1SDHC7vyq9/KwrW6AUlQH/4bhht2pXtiSZV8blJjkScA9pfr99
Lzd2QDqaB/yPg4ZEaGhBdotWB9YmqS+rFZ20KvXkIU5rP1j+zol6Hxe8F2ANlyXXxc9nadAgMtKF
cAfVmd3AXIeOuwc4cdVmJWSx4rSk+Lh85ZJrEbtJoplGxS2yBWE7aTZw7NVq3rr9tPGPkfqLWAvs
kMTkKdRBA5gMKgJCgUmU/rPGN2zUfeCIIR5FzDDavLTTqcH1POR5Dy0iWP8kaEZf6nB5eo0uL2WA
bOX4CGH/llLM8hnsx1wJp4LGGPEwTd50OPlIpRVclPklW7BckbtDWAHoaX9iM6Lplg9DlVgvClvx
MgP5RXlAzribAJo/wP7fh4XjY2K++cVVv6zbqfofpS9DOqZOLDV2lgvJusn4j/uLvxBOIvuK1yRT
uWPetg3cLyjfsAC24SExDPHWNU4POIja8t/wWEG1RVsqOW+21caSqdfSBmvyQHL6cGZCEQ1yWAVG
ua7QB7p9evcuovgfet0zZ+iTSYrjYMl3TOeLq/kx9Pc9KgfPVbRSBgpMjTkNrCDoJc3wm2gQmSV/
Ml56b8XAfcjBJxiF1C2EkLyhawv24760JsQkh/2b+Jt7qOmUTvRuWBKUls/v60c1fEB6qmwgc/Lm
uQskCbvo6J3LuLGJOj2O1cYC8q/wXvi9FWzwPKtW+edwENjMvkQmOy92UGC1s/U/FkG1NLE7Fq6t
kU17YHME1DB9oE19aAvx1lZVpl1unFXW+wuqxgdILKCyv6J8JTyqejF9BCP3t/rV6oFaD8PNGphe
NP+IvAR8uKB6rVCUbutXmPlpZbPnC82Xqa1SvprPmlCCnuAKqn3A2Ye8tKaHa5e4k152hYDPhWMJ
PtFBoOw0NH4to8aDAP7hG7gWTbKrpjby29E9jSEYuQMZLaERKaSL+jD0i46+SWSRxkJqr9Fpwfkh
W42KhzUPDfrzHCVioBdxbYC8GcmcEnRSLFIHdgR4LjRYmwTdIo6NI/TDCX6qNoV3YhoPQXRmXPq7
QifwcmnmbZng4Kd6VtZo4kf9C/1o2NrFIbbNcBZggks520IQ++BOePFnn/Uf5uaPpDAztpKg9X/4
xwYp3QsNQSgfNL+ca7ryJagQpjCNR/9nJCvpAP5pRRQARcih7nxEJd3z1V7ZVJAiviMvIxswJLZv
hEfgQiG/GVQ7s22vm0Np466eOWNUl5mEi6Zr2urXzB51+IpBRsOOzuHNWaFMCtyLewDhu7zInsJF
n8b8q9XFIyJ6YZ7kiGrxR2H8p6xsCLmEYv3FXuhWo/PXH0GlNapVVZrnQvr2nVsP+8Mgrgf/fyzo
LDJDCm+O/Mqu3uiWPEB+6HpBs9HztjJj5PB8BR9U/bI8/uz/v9RV0BoT/yV0kZDFMZ3l0yT3jJaj
jkKcu48wXkkCA3vyvo4sr/DHQFHIRPC6/BTS7p4OGZDhD2K2pXhNVZ0IpUw6Zey2P6m8E34g2jIf
ExN6FGG4I0aQdQJ6+R1nVzsA+7Ks1GLQk9K0HEoAAFUluRe6OXYHe2G9MGt9ytrbpMHRhzsrCVuR
s6NsZlvEiOghjgL6FRCOmmpgkfMi6RekVIuywluRt71EpAeI7BOXopifL18iSKGC3+y6jSRIbh92
CIxsiqpSnzHYH86qz4BtKGhBDJNsHveO5esY4oPAM1OxquFIzUQpTSNP8Qa1ymJ/L1uhMjiKYzjT
lVS4L1ElFgxkV4ukDn8AwEneZ7/Mh7lj37nPYAJE3MFLn3YL8joXePUNKXns9gGDQId+aZEtQRhk
Q00hipPdJMvDcdCLnaH3IClQ2YNQKl4RNpfvus/CWL2NWiU6VFEBz25tAcRwpLvhQP05mbFeS+tw
QTPghSPRgqheSg6MWB7iZiBHNTpFTwJp6puYUIrmctYIdcUNG2TYGdW7eePDK1+4M/IpyDWI8Tap
yE9kskhVhAkyHL1y7/PLWhQczNwDYdjVZ2rjgmtNy6DkQixhkWmm2tM2QiijsmRVu0+Ls5rTlnu+
wG1/m223D3oiF79zkBWHMa7CdJ/cbclPimtNG0bEKsGQxuzlWhv6wYDDumAdGDekFV1hyRutxJyo
0EOR1kBVkydeYQx82qtu4ORifWj8YTVcKhtT2/CDNK/LB+RQ8a9LIVZu2akRsM1rXK/zfGw7UGHD
7fbA/OXqQbog95QXRkUJGa8sVIzl0C37EMDwyUKCf5LnvJHAl978Kn0frnhZtb4ClIB4MGlLYyLQ
ao68wuOlYAuckWPuBHeUZzIsuDpJiefZg4mxaLmC2V/oI6NhuflVr6NgqxJ+fVyIJ9HHF6DsHAFJ
c0Jw0gRpM0hYaFm5XQpf5Lv0DB/YFwi9kwD89LGd+5DkA28wz0mCHNlOWGbP27Pq5dNXHN/jjI30
//SXAQpPH8iJpuZM0T63DGvU39dDihEHkgTvB9MnXjUxMJKz/BbGSp3fQSdHJdDPXmr820qk6vjV
dY1y2TDyUlqEcn1TVFm4nb2Vi0wdpLHvql/O3K87B7zxXTo74ISpJDI1O/1Uci5Bn0o7U3y3y8V8
/w2H8MAV2s9QIcD5VSJQTV2X/SQq7cIq14zhNyn2q24wWuV2GEGIhScG302P307opl/APVmEJi5o
7jfdDkSIbNB0vRzcplX4OamHUqgEXk3qio9HgtdnZCK2+ecDGZk09N5GPwFGSG45a/j+WR/+YNvs
YhAa3I66DWWRrEK6rWr9ZbOdMpsAN4Z1uwYH6dXlwqCdGecigRda5wdAdyyO4DT44YegCdOoPAsB
m/DO9Lr0zTvL1Lr4oSWlLfnePre4Dnm7KM1qBu2MCxUJMtxhThJHkPtXgArfkcZkX3m60FF1eEhy
pcmhO67hQU+7rq27/Ui38gPpc8LmIiWtvYjzFotmPFmfFaxqWfSeM/8/mgRNrUbFEBaOoJUaeq7Q
DwFt2UlJ9RcJwFKEVKPxRJt2nK88I9OWhW99JlVPWV3jIfzfX70UqnDZfesNgQKZqXP56o3Jo+k6
YF8l/bJR3AjANIxtmF4lGQO5eYuosY7qlKmUeyQnX4ekYivPgZkmixne3sMSsNE0uNvEwQ5p9BIo
o8hDfpEWWP0WkL86KgaRXRSjETxlvClLf4dLyjgtfQAJVcVLhWcTtiEEKaD1Gw8+KWeqaPIDr7mn
Me8BA8K4j37teFKJawYTYcPRnqeVAmyGuQq6EhP8zAs/NBNj2GV1x0Pskaxe30VcYvrftEhKl+P8
LGf8nfsItWpNJhHKTAPh8LhxdJXdEle5jNKq0Ttv7AVTxs3K4uZt+/mmhfG8fSkGLRcNb6q+Pa3D
+QF9yZ/7rRHYpWu/YTZ2F3UaON5bQ0c5D49iznEx62y+wsxSSHyDaqz6HajPktPJ9FePiVOpcpB0
Bgxrg8nrCH3/S93LocA5Durioq9IzB1GS8WakefRTWtYjlPEeTZaDExDTneKex73DYmtCZTAObt0
mytLm1KmdwLKVKFeaMoq730oaIlvluujq/YDC+nulCR1B1MZPxanQdNZumra6nrZihXaMTeU3Loz
Zo7fxTtNP0dP5kv2BkNAOhT9aK9KP4Vy+SC08QIrnwUlzs4chNRyaX4u3QqAqRolGr8MykVoTclt
t+LLRSQZFm08Ke3kN+N1OEzU8c44wNbbh1PY4kRcLzYOyP62EcgV7L/PpDzUAx6NJ5POUIQlSBHI
imS65nejiCchmcJeLBDZPspHK8JL3fj6QHn8Evttz6B76e3YVENTvHqcvcBfoxSR51NaHrgwD/qM
b+BqrBsXFGMvY9vVKIFXpdOs8cZqVtTBwAkbTXaxMNeYtb2tJqBP8VMEnJkRTrLWpFi67gOVnrrb
x8XVJuFcGff7VzNjV6YbVFDgD+iFnxyburEHuKSQoHPojLbORWbmxW6SgRypvcLUXw/G/2dGheEh
QSvwUu4j5aaDTwxj/BRcmU4ecDlCpBzj+DfkvlxFmHr4jqqk75kNYPcXOIynTn5wUxEBbLakAzG+
Z6rBrFqWLhY7Mz+RMt3quVg+btO5ZrYb13j2R05VuvcM5L03+z+VSeql22RttLCfR+VjTuFg5K8y
3n0VVrOt6ZDYsL1o/zoUiCffV6bonjFFaJOsG/++BmLYLPqoY2cNi1twhB+ZUU06X1pD/e/ZrKvo
cme6TWV9FbJFxRWxlLrHt3+SJ7RGrmjtvXF9nFvi1/UyrjUWKZ+htVLnJOV/Q0azzgUliw8hWko8
q4vCyRpjItd6mP9byyEddJAPOAS5MsrWgEmjUZ7YCNnsehfnG/q0iMmxeWOa98qD9f0wJDghcLH8
Qu2LJzikw6bq0FOGGffVpyK+mhDsK2wvc8FISuubnfRqgPLSWbXtBnRvRvzS3zRVcwsfDLWGjPgS
TMutR3d/FRjsdl5rox8nAjVwaiE8DXlo51/B4iA2vTJALndCaq1zBIgZ/wPSC8Z5kB0AiZyBbIRO
UflJj+WWU2r7HjCqhlft2/iWO8xfOu9FS0q+/KoqFd0w8nHGEUQQQ36/73CF1G9EU84+5Kf8hJSy
Kl8HNUEl8zFf+4RaT3jT+NtW89SzvD5wMJDbZMLaTD/vG53xvgEya4p/18J5ZKpWP3xFNRMEsywJ
vtwdRaTMiH21iTpwMh6kEaQFIG0+XNpFGN5WEjAiBY2AvLsBTmqhrXaPfu17YYwgYsVddUAinKI4
0mcmjTKCkFlZarCxv5OyR2Fd4GokvvsHxU8wDnilXjdqFJLYUm7T/p9kjLQp4JSxF/YOZ9/SL0XB
z+A/zfwbxNx9A7LnDDXy7pcnJVUekhBQs2yEx8xy8UUgtX7xhjfLb/762gt6AjLmKBNuuimiCfar
uJ/o5H3ms8SNGs4EVaPkA8Etygbfnf/omgNcYMB/bqcsgpShvmxHWUqZFZ7BtacPGxUdxFlQyTh2
6RwpUCTwzdcsH1xKJtw9QaHVK4nyDONe3gb6xnvydUJjUHYbkT8LaaAY/bWK0WihrpmGFwiDVvoQ
49ZOGVtlo+ovX5jYgXZ9awZ8K1I+cKJd6z7v+pyCMGsx0Ddu6YCO7NggwsWZZ3CievPsyA8cnIpA
D5Ycy1wMsdu2Zj/m8L8uZb2ZEITC0Z/neovRR2S23V4UO/CB/ECJHT0Vi/Lsj3UT4VIKu3styqV9
Z6iG9GocP14vzxr2rliEKEC6kkKc+R7mYA9Y33ruJkcesVsinsYK2LFGMkdIORa3G8B74j+7xm4q
sY5W0ahsbqY9nSVF2slL5L2gojihywrfvf32lj7XdVeNH6uftmv05HFTW/gnEM/fQj+Js9RBvHVH
yV22UaQFPuTgbbcROk3qYVwhKF5lXHSPwluBPgmv38Itqo3jAnSTUZMJTptxqRjP9B/Iaib5xWoe
KU7q3/GDJovvzfJ2lS29ZbR5cxVZW1nCpCQCX5n4nmOud3cIJxUYkUVVN7o7o3MBZuhFQmF388X8
5I3ztQdaYMghyT7TlBO/Qcz1flLCLXvj1cGUP1lCJjKVZL2aQ6ABdUBD34YnbU8Rgvu1kxhIZuV7
efc6BRY99THm0nAb5OJoG6XsE9OTsXbLOXYf8XF3PFGFmPqad5ICt0ghTv/utOzk5yF6xetJisbV
En+Beits06jJNhAqi3EereoVk7lsCMK3++XcPX80G9evL5RhtZbILy9EP0k4QxZyXncupHdGp57g
/05oVwOc5AxoqY6hjPHjhy5zHmwsRCDjZCjR1X9ubkX5Les78pXK90JAjrTcGp4cAkHdBkgG+BO0
gBEDZFEe0WyJVr1ZFrhnol4yVKp52OgmD0jq1ZPxpRU3+T/f5Ge0VmukYUsxoFpBaKtTeCMMwu0s
EgZVBREilPj90a1qocveVoS+KNDPFVBkDEER/dT+GAvo6fa5QWlQNw/3ceRx09bHdhwY/5xurIQf
l5s4yO1b1f5gnOhrUgUzChGpiCOFiBmQMLS/tb1AHiqbDjPVM6KiKVmyhxDQsb0m28gww2+9xOqP
XDc2+k3xKQfktso11JSSRHkAC2tQkz2V5hi6Re8MfnVYU6Jysb6Qpng3NTcNA/U82SVh/hltRcpk
Iw9kfpMPfkelCJ3T04pdIYFDCjlN/s8dxQ0+3hOfeOIlJfyNR/OKFtQIXXWuFt2zXqCXWri62sxn
2eCGexKzLiGjFEn7dznh3RDm+U5iOL0Cj4OJIQeq5Ob6yyrgdKTEQw0zeXH98JkgjrHxpGuPxkk8
8fw+uy3G+kvirrNsCFW5gSbiS6RJPTxyNh7ZXO89e1FLPx5UWZQTuzIBgsNALyDykgkLL/t4dBBV
xhghEce1UuGVRNxH6D8kaF0ekFi9yqM5qbZnSobU8JmM6NPqDaoHJrwvQpngMFiK89itg8nwB7pi
zQsijORp8VPwJRizLT4ck09voZj16foqGE5aowzeXzgL7jQdmX46xagqzxxZuw6Sf5S4Pr5fYHqz
21/XfFJy1WMg6zF4BrvbCqVy5XrdPdxqb92lMPTZcuzUL9Wp1eB7qYCklYkzjSBWQFO7jb+x0Trh
iDT4m4gmJ0886jmYeTRNTX+ZsPuipB6d8YWEgEv1XMOl0Z0p/Vnchkirw4mgnVcMcf/rGm2LpK7i
aVh9JRJWpLtNi+qLAxFkW8DVdzhIbRgo7oqrWn3OS3E82uhkNrtjrLET4JKcQUNC3LBhQOeYWNvd
QkAsIfzMeRko9JO7z1g9gwCW6YW/YrdoxlqNhiNIaFALINB1JRVDcWH66Na6REybrn/ltuzamJ7O
jSmii+QuW9QQvv9oVlrYpraDc/chvNl9fPmLV3zf0D6uvmLM7u0du8aM3hx78rMtHXFpnwLRNHkn
/V01gh7YIXEIUiX0K7Au8F1tGe0EHenQDyVM13/xQVTOB1tJOjhWVwGkqDJrXzAsGYb+iGrhWAtC
MwGKW7882lugRzF2+Gsc+u4LcfcCqD53xvhU9FxaZQ8Yiq8Z8a82n4PxKfX8DYyCn4tADgjtYIhF
z77O1hh82xnfjMwEOUrQWdkjhiyG6RJCZCn4nVA5Iwk/NDN0Cr0PcyDrPLoYZMXyvEgs1GgZnI7v
dCq14cpx6MoBI+jz3g4+HhFoUyeHxROooMKt/nq0nOC3r9ZcxgH8EOprVEJTjhZ3WyKfPCtpajXe
zLUIWPYcPMsIAvYsYUUXQrT/wINYF76SeR3ZwZwhC760OMEm/8HqISG/mxLJ2n9cMfe76HauyfpK
utYY9EtxXmQ7LhlcG3ooMSDnEfanEd4ZZglWxicXxZtMG1++IclHWkdFkaz1Vn0QPcC8cUt/KRix
uqJger/6G7VX48Mcpc73q1wV5/Nsn+SzGSwEqVc4vlh2/vutF5FEQ0/EQ06s7jiMJq2/9/5FpoRp
LZU4iJyDcg2SxsrxIBdCC0NSJafxfoF0bAlQNUTilLDUNtGm+E35uWZxK5CzsleDLcZSg68II5J8
QYH0b42xGxFMKpFd8KvODEwDmscpZn2K8HBTM0K+A3sNMTr1rONkPXSD5VNKSbW6i7hTi1+f4mej
eeDvhVjLqMaILlBaMEplSxjje+3TF0zt6ESHVMoIfj9pjJVlaqWFTOI5od+GzsmtiaSygvw2oTKm
sKJxUk6amaHJfcfjp5DvJspKOgp4t+BS2vW73qUzTC20QnyhjzA3fPQM5vgTvPYX0eoTxlC3POHL
3y3mJC1B511EfpGCF6mIcsmZxa0a7Loc8ki0i1SOLg+DjrmeaaE9L2J8MqraAnPgPFCEXJx40LBm
cWsl9V+n5CFuoZ87e9RzG16fdTCx1PSwYSVPS7UlLuPI7r/XH6iaA2M93E/dTMsb4RiFrsVXsgOn
jy7Jb669My7oXO4GDRkK5Ghwc+2OOmGrxomItlzN//dz2iCIBG+w+da1BqnOY1V/gPYob6L0i+Gh
L9tDjJyGsBwPH5qDvlZJSPwfetElozcaG0CD5+Rr3cHYliCspD4QcMh35bkBqtprfIMpfGAS3m7A
iVkPylgmtP8rzxpHvVf1Uih1BFunFq1mM/Ek8xlJl0QOMuCj0rXtQDhblXRxTccPrOYq0NLTB1yl
DtH4WmgkuruEvAgAQ+19rHanSBkxT3+uKYzPzQGN2QBSvZDDVppC1/JkA8w1mbQKdXId+bg8tIZ5
b1BgiXs6Moc3aF0VQzNDz3gVPjLoptjjW2NzjWjOaJxC3IV3xYFsO/bg5vXbq78KhNnzBnwkeusH
77sEJW88Szkrqpi0lxIkCyF2Rvz2Tw+5MW2ygAkdpFmsG9LYPuQqEavsKH7Sqq8C21t4sN2mzOPn
QXdVMADJzEtVRZYLtR+TrtB+PnFPpXVVV4gM+iZjbnAK+/oq8DlvjC7UJejQ8plB8alI5W+PK2xD
Z69ZFH95Kj/G6HxfZf5yLQk8IOw20EV7FuCUSZ0Hm9seyUO+QKYbC9m4hNjAxcgxksF5vLV6hFWS
7Zc5lfEqFwVBWzF+brcWzHm8xBr+Wvi1i36IqVVRvR8rbtNCzWIpEYlCO41RWMSJKbl7eOJnSdJ5
cqPLs4C+dKoaoCx+Mu/dCAZAWKNRJM66tw3y49af7oWnstAwcXm/bawEmZ7S9mbAy3H2Oy7c/dW6
hXHbD8QtNZJDatvDvpLr+lIP884cmO9+r61yrmWq+PihVh0qiHMhAEr52nqW/hhE9zNslaF31yV9
DtrNxMsrZ/Tma1WlFKSmbDCWLPG++Wr+Y7jOWT6e7UyTpye3J8Lc6uDYnNG2McEcS3bEnielO+l6
a6tb6ja23hcz0cMhuWYcSXA6aMR4WOwF5xhGJkFJQuKzKlSLjtNlyCO3u0ja54PjRUTiMQqQY9fq
w19l2aHEStqJulaS4PyiGGW1ROcHZixyBdb2x5kVWdbWqB5Ep9E8o71rFGAxb/Qi0Sjkrl6GQlmz
lPOgL5oEaHCr16GuOQp4kouwvwkZTYJByN39aTRDr+p/WptGbdVBqdoaXY0zFh2idQIo75J2ht3b
FCZR4YHwqYl/rttoWhW/jE0gN4EVHd4sy5+PDbIGIRlbBXN1j6OY76ms/KjJTQ5kzDFC3zAlAqaP
sqicLEEBhjXD4LXAx2vEbbE4tiB0K/1v5KM3l2rCcXfce+nPDvCXAFeolXK1DCIympIo15nCNe8E
eMD7pK5uNZGxr1TriZyo2CzFVX20MFZ7zuKLEWEtJ797ibK5uiJ4B4VgBwek8Aie47lQnNwU4ebk
PbBQiHx20wQvLOEkxoPMv/ehRfZOlzH3YuQQ2LuvixG2bLSMNfxltiXo0486FjdoRnS7CN6sZmsX
G1qzPRDa+hPXm1MjKVQzn4nJNtFmw94ULUI9ACEM8dGLDvgFlaDO40f5bU3qR3CyZQqhiHx43qtk
rvefosxKWxS04/C1HRN97m7duP6gMYgCgenp334g50Hp0AtKA2M8a+XOfqjThYux/8SW9k9IDZBR
HtjTJYRbNm+nQdHUZcL5KH6sGlCQpvw2B5TaeWE8JiBASaBOangzjgWNva49tPG0Ehf8ZxoqD6dr
Qxd+PvxksNs4U9QMQnu7y3/57XptySb//fdC+I0I8FZpeaYRbMJqY4B9Orw7sdOFkVbgIXpyBS37
fXiYEysvLVrCKoo9V56kssZEIPhPijCcl8WylSloKYACwQnqkASw7wfpeXa69+k3DS+hYAAi6Vgs
dOR7ZT4TlI6mmVjnieTI6RqJSVMKTa2KF7rs2OZNOlqwOC7s5zTrGVLqAYfobfLCNMs876YFVv5+
oRWNMFOv+U3VCerKmrfGKenRcdIl28g8zDylVNbTR6HnNQ02lFW8qcCtP5JQzh48gAZ12F79w5PJ
oOgt51+WT3oYdfFnbwtkUAefQ3juy6ckzNTsFVyOGvsUbDBQ+j9gRcZcYuIDGsI57PZ22xZBrC5C
b7S+DUnQJ2OQNXy+ZbO63qNXOavtrDSi3Ng8Lpn9IT2p1ND6UCcQQKKjWGOv4zG0rJuwk6CHQEbh
bajp8BcB2tp39TEsbRsJ4m2LGRlj6ZIJTp5oWTq9yBh1wi5R8d5re54POhEMfCAU3/KwLB5TUo79
uZlWYwlFe7DlaWZT43ZKmn+0nCERCwxSXZrTGjrSgZ41DXw7Ne120O1WJ2rXMo6Wtlve+dLHojnV
jUA8xf/KsHYBAy5lx6rOVYathF5+6b852lpWPfN35WGbw0h/7cDC0F6CPOCoTqoMIokpJu0GUP8I
RnkD8KZF7dcO1VMGDiF5ozZViA0AGbUkYGncwo28+qjgN8N4Fgiq1lnRlkprMP9SgqlmFTk5Zz+j
O/pm3mvWzCvgep3sjlP6hC2jhPLN4b5Ezk/VL2X67684UR3i67RlGNcwVziQhgsG38s21yrUjde6
atahL6zJtUC7pRI76qSIsZbthvddwdO2V0leAimyHmQzfuY4Z9CjQtsIilgChnvPytBLrhPhBAzY
2L8SXbhBbvboG0Ki3wJ0IyFmGo/hmJXvjoFRBEMJMULRBHP0cQtVC7QZuLZnZATrffXMrsphLT3V
Lgb5tHXAEiwzT5bIPeBlY1e/y6N5RCMoU9MoOBvUHxd8twdMT4o1upM5Ir03jzjJoHmgwuePHI2G
HC2zmEyb/9FTeXcZcK4ai2qNWmi6YHdT1A/kDba357jMiwBGx2lMMr6FjKJyTUS9b2fQAGZON81R
NSVOuHWH0cIuZA3UgB45oUr3jJmvxFlQ62j1xJC+5uvH4QsRUrjQbph55BF9gi1UDA4FH2c/l3Ra
zJh9okmeRGT5eaeAsArEPWyIQmFfSI1lc5W86m/Z8DfPpPggqm39aWRqQDiFDp+SNXNLlhHLCHct
pCzQXoDHHuCVe/rnf78qodXasAlaWoN4HOLrqkz+rkFASXxPhnOHUbE9EvSNjDw13HptCLAdeqB4
RHIi8yZdNn1df3X+xOPYnTQmAQW7h6u8r4xZQHaMotJ+J2WhfrKaZvV5WHU33Kh3BgS7fWi184up
2DUTBmkZ1X+PhmJOBBtb4Vp3RBwKw4Ozg+J/FGBcqLjdUjMCchbaSecdItETK7sV3zA8MQi1capc
9D2XP3jgnBdiYvToCyZfvAIZnPpqzmqOJUsNMPe32rz2hr34hZ/qhMBReQ8WdNk7i9AFsYMF7jfN
4TMARlonzl47hIoUclZWW7PgKIWBKn8jC6dDrk/e0RVfq3gkHYcDaegtWz0iyskQAqRy011jJS18
5uNDy/GE6495rD/PCzhHswMTfNv+kD3O6EAC+Qi54G1aBsZwpGS2/8VNxV+ceqVUFc0PepM4Kwo1
yvM9HXstiQScsiOn7nx97lGMB0U4sab28FgsroojD66TEdZvD+9BysU9v2rxOH4yOM1sHoVbYqUA
SYU6HtlrCvhqjSuE+djUSdVqx7heFi+cxwnuhxN5sSw7I8poDZS2sJRAHs1DwYLdDH7vLn6Gxear
br+Rr2Ko4oMBsFHkl62axHh00rWRWabfYXLTz2K2L6aSspuMGgtCy5qgftLxmSnB4mipAjjqIgsV
W7elFr9yeX7hGKF972hJkqaN0r2obm6d19o9jflOq4y8IJUTGaJRd/bs24jtv5VgVa8zZSzoqnV1
c2W4eebRQh0CpnZWL8FiMxMQmz+Hj/JFO0vP88EefvxfcgM0ND0iUSEiLOoXmZORxv31rBkT4pxQ
K2Tu4EHbDHRjMOJS7skQhaSVDew2wsxhh7u/qCFsiGT8+3ikLC3WAUV5/GopeaS+E8N5sWQjsabB
hyxKYfRE5HecmPEbtEeg5XzsDvExZqXq7hsbacB41nvWdVNWCQMk9TPc005TC+TyhV0nj+6hK7Zj
CElhG3kyrZMAe5S6l4WqaBWvtgAIiVCvLeBs9QUiNo6LVzZJsq71Ou+nO72Zjj7Ae8XQWIG+LYrY
AmekyodZQinE6joPv48rR1uG42crrn1OMJI1RVo+IrMEX5LxwYo/PhZifMdsPZoPQb57bEnmSYhr
rr6rKBaMmoh0a1vB+MCFytPLd7tmjhUR+kz6hO8CznI9WwpVEqcOPn8gIlSVA4BRFaN1nW8pCiAs
/ytOkObdiWg7Ft/4VlfA4Gu3p0jsdgRZBANpOOV2UWyR73za8k+526ti7Mk00i8dfWeH7YH7L0PK
dEAko+xQ64QMO9zN6sPBRb/X7TqZXxDPZ/SjkZr9p+Cro7c0Y1rL9+cd3tFaNJraV8328WAUi3cR
j/004qhM7sQUnip2bI8yZcjgWnINe8UwrTkXsoreaOx9yHeLVZrujARm3Jycx6A1j4lPjzei7p1Q
3lxQIPvZDVEtNhq4PECGWZOv+/E05RrW1nBSZ3OSLh1qfj/6k3HGNoufaeUXL++oxkg045mYhdW5
NjYc3XMoXQR3WhC1g3D5I7E6IcuoYf/WASnqWvmrR7Ghl538MTf2uYU54usJL1zMmBQj9f2QNHS6
thnIBTtx4y6csJ/OD3OkvbfTheM8JWaK2yyq8zCIvuZ0xq36HrWwDeyjwtGY7y1Pd7LyYZDHVIHk
UVXlWau4DkDvb0zs4JttVTAPBmp4fGbW41inpcPrIwa70aH7MJQRu/zdO7j0uSkPlM6yZsJ09kLS
176p/6jFQdhHvO+fKBy+KtA4ChkMjE2q3+1ge7gXaJw5wJgnBTzQNSmlutuxRA8cFEjrnN5sGQPv
m99062LT0L6lj36F9rLyPjRVnCITBT4nqWlZolgd1r6VKBNFGKydxHVly7qgDXf9n4Jc1rKOB8Ah
NdhvHSLn2H8w5nejsB872Y2D266XPX6YPiIcAr5x/cLONWQnmNtsA4ze2CaZ6LC+iYcddXWah4n9
CJnNHS0C+fu5VbsxVD1w+GuLwwy6JcXG/m1t50l2+WimISHAl8GzOARV42J6IVguvkIzzlDyClzE
MafzF+NBslBZ/h+1VbxPl2vcVHqMMRHoPEVuWjyIR3oC86WVZocQrnS5guyci1efRoCUPYIWGLmA
0+BSV62ATqBweidjvusO4Q382xqPL0jGJEI6DOzttGV6biaTDt2w5XRBnSp15M80EgCkytfO3zSV
0dmFvx7huGbT3syXPtJNT2p0QyomcLPdDEUpvqjdmRWTqb0EB2txMEzm8rg8uTWxmhWi2a7CQJ3T
YJ8n5Sgf5I3nmtRjVGu6GVIQDtyC5T9jha+ak5g4NN/d658qgSSv77Xlh3jQrrStorUBj1wwUDHz
TDzjLyFsa4lPFEJAc4ldZbR+EkSLFGJUCq0BH5Ky3hqr3TGjo/sdc2K6hoBSNJ9cmR3glx3olQUj
uPdjOlnp3poUf876BnSTNKF5vB6wkM5sE4zrK5Y4Cxj8hi1dfNBgaR7I+BGlpPpko03PykeJVItW
vNKZOR4GFqsyUFv3cgMclZAi28aXvv8HRarriX7LtZ2N0xQ6tXhkmrcPyhinpvAN6S+iLJx6Z4NN
Ngt5DGhEjAT7pJJeL71duQDAFG7h6n/i8Ijdyjg7D1b4TOBccR5wNSDHwzrgqbt3ZzFDKoaZ70uJ
Rc6Nr3aI4iUN9WwvJ/LSVfvH6kAu73fGEZKxms6WHJaXnjp26/5AO+prWyooz/CsLUS29olAY3km
prcymvNK7kSQKNNP7/lECML912nEW/7xfmnUeeMypu/7sAL4T4Iu4cm4PksFrUZQk59pOp3lea37
kDEa/40vckEa+gYOQewRFZhcws7h6kIhP5cYwmCFOrMc2UZgfWcSyoKyaHrXkcUwdmvYe0iIDmCI
OC5QSaQY96OuItlgg/WuQsggb4uZozWq0SURmtvbjaAP/pB3vHUbbisInYPKzGL+Cg9HdlUTRGyT
L5sqKz9medVJOsMYVh++CaWOGXfrXR6sgS1JMLPTojtdFnN8mEgoloTXs5EZBnbrwGpQ0+qDEXuE
OTDxz/MvJXr0BLadweDhqenoccts5b22z3MlRe4goDv46jm4wrYNdnAIbTBA3v/tiIfxs/2icAQb
fczPPlLFlRHP7VMMQEVWELYzna+9hd50PTmd0O/D+D02lKvs00QS9PzN2d+paMeUrPfKiq0Jp33X
DAA3w3DE7Dq1sl7DP87//uE1svxqXK9vNjR0L0jN/2t/4ew3P7ddOXYElG6sVyhPN9X6U1Rfjcvy
2DGQz0tqCsBUXVr/rhabiHjehn0SSU4SMe/R+29OC7vAtzQLemzoY9iqbgUCs2ZWgwNB0JYpJ79c
6rdodTQdouCk10X5qO7tnHcnV8MEZO9uNCdDJw2E+1xIZ6dwnkNcXDNdA7ZYpkRVNIuFRtw3K9cY
q3vwbvdUwJxLYRSIj7nSXw6523bwb7UN0qOVc4hXNCJH8OSFJ01Qclp5ZZIuzH38K7IRhUOnXh7W
qY8u7zFyqCXnKFF+app704//nfeELV4tuLmYU21iHP3r94rfg96xcYrfFE8wxxOS8Lx4NFlQrOX9
T4H3pBKigVrIAozoECeslzOy5mqLTeulr87dEoVTPsVmbPwGlhS74nRleu06MyOXVxF+trjIipGr
5tkbxXS4XR38E5YROqCHFIOd9/tELRhSVgnMTXsqxWwKO0LUmD+drB4iz3L2QiWGhg5KPeTXBD2f
gLAUHdu0ZE1nXcFdzfvssAAo60B0Spnepev/KWZqbA7aOe/ppsNGI2TdSRk1j8AJH3o/CGRWqf0R
a1iiaD5jOvgGwzl6T3ZQ3qolR9MpjtgFaovCjzmXT08EmlU/IDm+0NSFQGM5NcMyEnnY4pb8eIu9
RgA9ceTiy/w0ssVQx1keQzXHIp/LpAPvfTftCSCmWGqI8J5SA9nOSirMsvu4Ox2S75q7h1CsutSc
nuqguJb/p63MoBgxIySumbZEx6AAiEUceWbKdSITU7hwk07NF4N0GgneoXVoR6kyFTmFYJ6xZDcx
hvQXbrWm0WXB8IkuHvVywF12ascMTRo6eWk2duGdI4pCpTpL+dVZEKLRdIuxRDYRgRLjMg+Pf5Ah
GbIeN1bjMYrKsxBoVL5KHMaH/1e1WIOaryNkakC71lHQJWZfVf01U4YTFWvBhET29U89JTmrtmQ5
8Fcq+vdbpFUqMF66dq/Nrm5zg/egXfy+b0sKiPY7e2XYJN6nrRCqs3XFmOcWkd25gB5K18jNvJRo
+SeoEKaimypuoU5bzoscWQ4g5bCzclYuE3qAbKN5Fs6+yYK+J2aUVJ7J8WSaqlBMugydgvDU2JaZ
3RKBhuihHnIghpOkVjrhraBaKKPvXEV/YzJQjTPuEeBemXEsr2ghqI5Kjd38EGYJgAK3DdZa37bf
BojtQOxHvE5UMlCbh2mVTENGrXu9BYTcSRKt6uLwfTQj+QiDeEpgIfRuZrdmsX9s6xgF0WkTi3Dx
JwSPWhqadGmrofRNu4UfVagUXSTOaQoO0udPxREKMOjkb7EqLqZbFDs9MtkenzcGKgjDBoXl5s2u
pj0kse3AGKMNbeb2iq7zXCRu3bd7sTWkbS7M7Yw9+WEZny1/4yM/fVtkedCF6zxlWCLEdGyxrH0w
sZ9GNE1Xxqzvy9PnixBqkZQ+4ZXorowXwIvSZNvQa3x7wcUJxi4PGnxydWHqlKGT/q9vEdT3+HSk
bWz/IdEtwR/Cg6tlcXEth65yCbJmWLe0Lw+WLH2N7yz3lrDdMRWk5eu27ad5cya7Wz0mxyEXLxGX
d8DjytBW0vfq+RaRWXLcl1blmc0VsAY67f1rkuAYUwt7zNRFRyoT/8FUz//57H8JXcHxZuT/bGRh
MstOFzwjb0XMkgRfzX34Eqrt+CF7j0q/FupW6N4b3pnPC9CY78xVeDA03RBCke3pivJt5tcdh6kg
tigB8J9F1z7gAOwahZ4EanE6VRa/sWat2baKY7BpnBwKpDpYfsjEkVdwWMVDUJ9FMEptOMX4gwxY
yjE6dz1JMJ8M8KlaTFbV99JCxpoKEsUTHpY9i78mzkPCrKwT81kFsX1jbvAsntfHsKqlraFVy8W4
/v9YFWpskxkc+d/spFXxeZbcZalB5DLg0WHWOl5Sq5tSb9U51ngGhEgL9A21pT+iJj7+LIKrIuVW
7pRzgB25ocJVuytLb/L7Z0/EzfoDefiL7hO4bV05+IRaYTMTnmz3JQlxu3yQmvXiXGJbLq+OX7FH
7Uoyx9idMaU/L3SX4aM0YGfVuU3BZUS3SFCL60pKeJl5LSfar/v89TXRIAboq4ESMewuMEm+YR7g
pv/C4A5TDZekulGj/PPJkNyCivxapM8OwTUohXl7pRWvQC+oIjN0Hguc3aMIKzrIhFuvgKF2AEl3
QAFyMfLcMFCzJOCLmZm1TF0VWc2oL5dAT9xtIuuCWoT4lBnqB4W4PHdb/HR9SkyPqOdfI/JlxGWk
LnWkdZ2FBCSJEIt7zBT+cRvA2EPtU3biJQzp4mg6YWaxvlzCW1SdRp0YyxDHbu0eXVzTiUFnlFdw
e6bRZORp75auUly5FDKnKxU2sfhbzNYJgZKo9KM+eBID/QTKEPfJm5gO1Oa/wCTvZaJbtrTRZaPY
wWKHn2VeO+4G0ePrwoFDEFa1Q0jvC5jd7zPj53IMlaN1xZKNG6LEkpJRJQDccBh6OUPC1/Wr4784
GBXEzPbcwneyBUg0o3RvrNv5Jpz/URkE8gAAD2ujWw/DoH4VgNUwGKOvNuy3fHN7f8ewfanhCKT8
635EXlxMDazWat+9YnSHkGfXw1kaWAZhcBIuSiFgjcwQiH/ks6Rz/UBHatYFhnkMHHDnWeO3nfDP
BvheqMUWnNWx4PIItfGT/Je5jTXNJH0gtVCRlnQTd+MAWG5bn25ylhKf9Kn7HYBVMQwiElB6HEqp
PeoQJKzEONSumF7+ryG16DVpoa1k09l9007VRJ/9+yFJsftE1vZkP0sztUgUO0x9IiSc8OjWyE/2
Jk3E3I4R+GSBaYtEx9HYeJ0+jiTGb2EbOgYQ0ezaP1m0ICXlSrjJ/UIybILaTK9N6ykQsTmRIbxg
k5urThHt0EE/wulX30PmLBSk+PyR+G8faVDRyGotgZcUgJEfT6Ff+HRmH7+0GXYTt/MlwVfHGvK2
RWgmgEr3G+Bonvni/LjL7H2hLSKRB3vAi1NJfbNd3InHdX/H5Q92k/qPxmDRp3vqutQI0tggS0Fq
8IxnsgmsV0xQ/LBTPVIdBEevcPRn5OipPkD5LU/LxUSWgknaQD07b1FgXGZ5JfA974Lnm+fZmY77
p07foCwTI31tq4+QyV9k0P9U98xcPuFkDPSDMVnDBJ8IXTmxNWNo6s8eL4aaYH/Oqg/7Tfyokcn4
1VIuFw66QbRHQpNpEoefQthcB/pv4J9ugxZei45pdwSp9ZwpsIHL9DJLn7YLLb8EfVVLFd/NgE/3
A7ZCX7UWh9XHUd9eY2esjwpgTmJpMfhgcDpUkN47svwtLWCpf7ofmLwd9MvUMqwIKOQk7V7zCFCp
+cij75F16+6n/BCDFcOWOA03qEaHM77ovzgh9p0awleoxy3dUGMFU1zGhfkPS/jVGgcN1Gl21+SR
G83+f6NFo+PFMiBy/1oNWADUED84/hGbXm7WMYsG4ogpGjEI3/wvvA7PP+LiC1VTLXbWRkefmSST
+ZxiHr/H7vueKxsPZxGWCq/Az4pxzw2dzPEC+gf18oi6MJj59UZCFWXykf9bvmsv6V7Rc6dr28pw
ewBB2zZ00cZLEuIJ9BdyfyADrvTbJeZ0RPi1zc9Xx7OYT4sDlPZfp47MFndOnZLNT+t5H/D5WHFX
fdlTMWveyx70rpGVKO31QoVF39MM1vmIYHQWsJ4YHktXBv2JMTpfXP6ol5Ko/kBM3iTbqIWqCKWt
GLjzwnVR6EDlvqO031iYa6mq2DtrIfIDXq3AvsHXcaSzGewtGVHPRXcF1CtCZ2wWaj84TFqc5xdB
KewKXzU72NjrJ5+tUZfBqlBStvt7NdK+Byaa9a5ChBqaHz/C8dmMvOfb8baBe7ob2uLmZNGm7aTL
cV/zp6G04XSdzunL8aJOjD0c9UVPioonpXkHPyfyryw4m3T2ZjmYvXEaMoPcu8KEDd9zAeEQWF58
BSJ4OWrfjZq3TxMO9lz8KDq9FifU8pTGMCEip2EdlRVmEDfMZHkyQIprpYYiz0xwecnHWXBN6YH/
dZgqu3yNJIVmfzJouYgbuybf5QLI9LYyHSfd4GOzK6TLMucfEAY6lLGTdQcDsH66Fg+bt7fBdhfu
fRCHOK20MJxs9jBYXm4GVOrOOowvkg34/PqT4or2XvJ04lnMUH4Ny+lCbv8E0w5RlFOy9w7BGmkn
KDa/3hacvKy+LmrnWNdrpAFtvlxppBqd1yddNyc/DWEe8fiBb62Y/Kp5adX+fT9+gwVyL3kvgYas
RuugvBtBV1X2+bFJURArX4Pd13tfd1LR26yO/I/VSvtR1LvbLEn443lVZ6VlaWs69P0kq9CZHip2
zW180NCsT/Ya3hRZf3Ag6kAmfMPdeStUNXeo4GOHHgd+KSzrshNLNPcl7Sn5ewZJGyhth6K5Ae2e
Npa5YlJ0AUWYulro2enuzEwdqZ9z224IQrZbQaug55kfbDPInXz3MqES3+Lx2zA6ztB37PSBMw2O
16xaZfT/ed+7ygCTIX8kmvI7AyNATnGEDrU+c+hO3abBcHhrtD0QS9EqYT6pRw0cIW4MF3CjO7kP
5SCkBdVldxN7n7dEKnbivA3gGoDPao70D7moBnuprDS9nyAa381AouMwLbhdjLp4xxrR/LP5evrk
P8CWEuCb7Vpea+QdjL3VjC7TwLBoMOQ9gblTajRbjJ1+qCuik2AxUQPx9akQkStJZIfh1KMYus7S
yUcSaM3cKUjWa0zOYbHXMdIeQlOhCvNgjAt19LIPOjPCr7bPUSfWR6I5IACHZt0pXiOg60oXYTAB
T4gtuuXc2HEbKJu7aRYcqeKySyMLmCjXwadwjzPOqFn132CaknxcCca2ugq/mFBjB0z7M6Cag0+P
rcTPBiQILgXYGwMHPVhN6xcmU4PD+MP7Qrbk79xPxLEi/mIQb8DXKNjIfbqQ6g0yjpx9Cl3QX/3D
TzhfEOU2f10IPdNX9VvPGACSllj4dgEw5AmK8wmXKgag4//AFMeKrJqkyjmPvn6u+Wq5cLnMFseX
vzrvHFxs181mj8vk8RS+IqLoJSNxKtSvOckqIUqbH+IuvgBbX4Rb1h63us+qYe9zhzqGJJLrcFsO
/n0jBbHnqEnU5sFRw8j0Z5v0Shy06M2gx5lQ1jpKGj2Jk6z6k/CNYViSO58Go1zSKUoMUhetwdeT
dOjx0VTiNvFn1Y80y8j8HnTCecqOnTmzJLCKLbTMJqd9MZW2aAqdMM/u17w67HmnS6e0k9b7Vyko
/lW/MwthbeoHnyxKxQuCuB2C+lK/Q7eW0he9O5LaK4ICd3z5EqUNTEyTzvEBO5cdx3x4BsLH7xD2
Sp5XrhzFjkX+vzRE4WMNgU3TKrIMy7smFilSuJdDPAVSQnCdjSmAWCt5kpeCS5jn/3xMj2jrI9kt
J12McgHa6wTbCAdGJPk9cic4OkXWtpxiShGkR75qbw7aamuWqfCVbXj7jDP/qU1mH0EdzFxXWpwc
0kbdowx0EYPAzg6EUB5svjFxCyoKUDFH9Uqn6QrrS9Ldll55/81TJLI3iKtx1odkIS+amk2gd7F0
Akrhqb9q8GZV+/Qxb01EOVu9FG/bXsFAVSGxwdCX3lJcj7w28Fz3K/XqpWVf5vLHeQoKKg3BybUa
E7u5Hbo6FBQvFQk0NyxVimM7WZOOZitx+jm54UvbjueRmkFTnCCjfm9RLaQBkpVwmyEadU3rDV7i
IfjnKgps3g9TtGkQC3S6tb5sYsewrS4TpPgknJaQO0TiQxS4lRLFIzPXwrJDlhWV0Duge2HVQxf1
7orOcrpujDe+9h216poYo+X3vQH4EwReJKImDRDvasb2GdQ5riTR9DQhCoWhGza6qhBvVBKypySC
SXSAjoxky8fwgNsVnSyHxTdVDPhAfy4zBWUMeza5LYy3KkjVowUswBNg4X1ZfVh1wEWD1RHQ0lrZ
Tf47ibZMblT0UsvF+xgJ0ihwKeqoq9t1lMIRhFdPtivR+oejRwVBl2uRRF++MhaDr9PNKQF+p+0m
/xJB5j31CVMDfolksKMBLWw474OHBgkQml5YSbBRfybap7hsxFvKuczsSFkm42mpBpPLwVpYXgkY
j/ENPfTaFQE8n0Qsiv+FpAKG5AqOIilLe6W/5hOZlcmrAK/9jBM09OHO65CtFvg/OI55j6/FAa3J
W25uzeJPHj3jvCQPRmZMv0RQNYTU++vAdJtS5WFPZgmJXk1oD1RoeXRs5d5ngsbkBeQVLbIx1hLe
zajunusc9QMOEW9vtcNk3foMcOBLisGBJmL8QV7oYHXTZsFaTDzZAj/len9FAT/LHUPQPNJTc6MR
z+DxfpQzo0rM4Iw3bvanh3wqg+xWVwA/GK20jG4e6lOng/fV00+Vf7bM4xqAXgA6l4xkTJyIDgZM
ZY+eHjPNjFDw3fUwqFTEdxfodvSJzolBxzsVvSuO6+wF00oifkcrXJqwFju5z95Hc98Tb27fpnH6
scr0jU79vFik6orFruTd9xdAqRRi8TwWVUpeQWkzgf7VyT2HiJHvag3GUAFh5XeZSgEWaTUrEUbA
UNk2R3goPkCrBr/eJ8tS7BZXkcboph0emDjn8wZi0KisjxIzCpwWLNVFOaKkLEHzYOSJmCuH1eE5
78ajSAFIRqkHZiayEv7Oly03to5PHdsYYAxasuR6FtOax/WNWYa8/84AxkoRvdpKsOozfDXPmAQR
XNOWjaHBJrUl0rBZcarxRV62FIkSdzEwyyIa7480AvG6G+/Rpx7j8qlOYo3lsFcPrnR+3DElJEdY
A8IZ49tYA7sSyQINGVDgGPTwbYinCntLGnSiNoT7yQ62tCfgX04xUYE3f63T447Tjp0bn0LQSy6G
8tn5UchaRKZmx9mvG25X7fS7jEkNQ+VYGefAYzdIivQSnuz43kTMsyJiQ0z8r7J92ZyGkTC9OC1M
XWEjUIoViHvgt8H571dAQCXKImhNdvNpPXFiN549VQiRfutl5x1hsKc6iSVn9MFO3WHheaqbaKbT
skNpA2y0jTT/hxOavhV9VHJ7HaLgp1J8c9vcZQH3B+Totnbgaqr6bGV0nQpNDxeMR7Fj0eWrOwBO
H9o7BQn1UKYkKIJpbZ1FHoBQloJcyEf437xUPnOCPi1Qg73gsOXhz1lZZ8lRWWl597jKld2GlkTD
H8iNFgnDq47c0M4hB5eGrbfPAFx36DJoHW7c0lhLc4zsnc9OERCeAPx+tfL/iCzB2r1ox4ELYMoi
Al/c3ENiSOnTVyr9Yy0LlsSFYJ1LT4SVFNeYoJQlA3Is0H7FZQAoiWwhJRqiLwAKa1XMvGAIYxrk
QswhY0xe9dSJSuZhOShROJPCVqHeGIcDSqt73GizNKE6sHrlLcm6GZ0ih3Qa+CE9ayq6fheTTwzK
6BiFYLblJcDPHLtyM/du/DQY4W8UItslVfM8tkpWRnPPj4Aa6zFCf104T9uIP5ZEaftnRoCuT/oy
5XWWXZSMPCUfG/XCOx7pU5ure54xnYzaZ9Xc+dixCd+6vvrF6HQp10TDdKMcH4B90TiBCQ7stGE0
9ekmvvtYKEX4vxrNBOVJ1VXiD1zXVVcisY0AsSorHa3kvsVoB0v9sJk0npYg92nKpqrgOekla4gB
WnoLJU5oImskMMl32U2y4aivffO8B1wkNbMEio93IT5uc6Gc4ihpvQzO6yzjeAXxEV1ikEYuu5Jg
JCY3kNvwaoGC4jzuKcCMxmoI8B1hSukPZIN7n0OHLFm0B37KXBirrMre1PozFsNPkphY1q6h5fK8
A/gRIUaxlB0OFSAeMXeY6+iGJHD4dbf/ONWdvghrlYQd51S9/NMIDQrpk3cX+g3bPsYLqG02An6m
5gjTSfYpEPQqxSET1TgjuvLPNJ4VNupO8nGjn/964+OoL4hEUq9Yr3nrzram1a7lmMD3hZnrpvMi
AktFpqOgkeILHeJnIcHGSk+07EH9E5ax7881iLFDFF92EOCixl9vyklcNhUT5sqNtsyGz+EOSvyz
PIEMBNUpP3csJdATF4aPRZTa/ieydv6opK8RN83DX/xAOnLl+O9Z42R/3YSKBbIbBVZOSMAkFYOY
T+xyq8nOdlVAmV/xu8bOag0a557IysyO7EYoXMfzYSIiP9EAY4JJAOC/AJPIWeTXNCDyzWHpvA1E
2xrHpYEXlkJhC8P7Ddd+R8t2BaZso+UeakvIMdK8gSaz2JcRFV1BmIIBy5FoJxdIOpmhFUjnA8WE
2340tyvfpgKMUIzrCmy4x06ncRJdHAoLeQCu7Sh2ykrDz2WZcqMtbfXqZWJFb0FHrjfKvFUsrC8L
4Vzq/h7MG9x+ob33sqZDkPZXSIDr0/BZdd3PLgo8muG9a0iiLk6osB/HQUX7L4Va5qjHbnac1QgG
iQKKZYyfw6wYXWhxPDHSfgEcAJXqcXIDF4AyL67q+1qGtSYmBvEvCKblCD1Cq8w1/IKBcP8bvKy1
WVOHNGRnQLuv+yA0+A7rQ4koew4IMJmQAtGq+5fa7wxaRBvIGDz8NEvH0LTqudIbjcMfxnOISfVu
iniiWk8zFXB7/HEkAzNlyrjuD+5gbonpYlE88Wd7UvrLTNyu6RbNpz9ArXnMhlbbIj0toE/f+eI4
qmCKfIkOWmn4nVr2Z19wbdkizOwUqdnFg24HgPHDtWpzG1gddjZIyESsrHb12aFOlD6qnqhT2nRL
zLx9RDzcbAejcCAUcEaOwAzw0g13f60dCbC3Q5EbILv92ziCf2WZ+J2DUfMagzbQUOGiR9SR1NfS
EPmXT/WK0UFlEC448kwHc70l9T3etiZ14I6SlJ1XnbVg42/hLK8ZfGVuAZ/ePdvIDg7s9SFJWKr+
g+h3TslQpuZ/jF36bC5XvboRH4tT6G2mCH3ZDQgNuthKQ0BeOzw870G6knnpddVIu3eaAQb/gT9B
UPZtIiozNCOXmoxz2GrC3/R4EbJb4xfnq2egymMuxbMCmRouGNf0zHqw+om/JDoKm9qqvbhGC3B1
Q93EnsL7A1MVv3o/KAjsrK4rBXbDSWk9cU2LDWIjz/JdRNeQzVgAeCeI7uNmBA46gHsV/mqzepV7
/QlFgwwJc7O7EMmM4Pscv74UhWmomY59xqo+gbK7bce73XxaDklDvUdkNc2FVzgVwAvwonbWC9zl
MDyvYxVZ1RiNZFg3Akiq/bTTsNW8fn328P8zI4txL30KmlimN+umUFOkuZfCDz8FFvbLDGecLS/1
6KNoVisiel7smDxMlLkK96kW6uPbgkQfG74yov613iYr34ziAZ8q+jhdbSkgDOWqdGxgoZSPjgMp
4dAjjYbpDg20Je8RE/4brDbFDHn9ERTjQzmWrmSv4S90bkqUNxaUx8OP907TkOA+3ooYfqCAkzWe
FzzfxiNLSOgAwSqpXWSuuKeHhdBg7l5Wsj1eKDoypweT40pLtEPVbrjThlvJQPR49hunwRrLFYjz
7Zz8sWNbBFn7DyK06Ps+T0GkL4IwOftKCSt/zb4ryZ27zQiBEjlGnnd25Fdk70DGvf1ab/72WLOG
L6x1gV/5UwF6//W0Ud3XuX0VAhrbovO0pKpKSwSWuF5rKuVWj699qf23nauSC1gbGeQt8UjZN9/h
hHyKYnr4YQR8LCcEKu1HozfulhBOalNlv63fOZfNm8Rvc/nusgBvVNFVqtHnMl5Fs+XFuLEcTqnB
llEAYwurrMxCrsZ/VimWd59xzHP/hE3aBbeM8mYNQgcD4NQW+nUoBVWl6M6tpnJlsdKYR1K2KLSh
59k9Fs8dPSD+y34vIheSXZ+N4Bm2VS1ahkD9RXxKYc+k/wjGxHGxxYa+EVmExkfjSKQT3qr4hOhd
6EJvUKvOwVvdENt6bGVq5pUXPGNAkrNUqOO4q/8i2HVox03qHdyd6Ybr8lg7akOyHns2kzCcggt1
WSeXnS8nvn/+LZ57GBPDNlws768cmrDn3kqExWvCa5fQPG9cc7myOToxAHCxuO6BcQNKk8FvuA9x
DrJYN/d8fh2ED9hfn2eu3X8k+2nu40bgzLULOpedkeqRwZskYX4MQ/vTldGKegkc+gSP3tid7S0e
ZjpmGo+wUZ2pSyyHkCVeO0QZ4pw0hIHo7Gvkt5aZTdj7ZXXLYQxeJZWtx1Icp5VOsNndbsbgVXzs
nLz6YYqqR4QFAcOibo3oeiucZ4HnPYNavbZAb8vqcbLWmZg/gtgJUJlMb5cnGLFNj/5i4m0s4k8O
E1OK8GMh1YwAXDwdV0L90KCfmn02sLkHMFleQbuiv37q+UlOHkTZaFLmMGUkRgwV02FIOSHDq4kA
FW0CjFxd0zLGvQR1YYyGkJsJ/1FXvLjDFbpz0wirPV6cd2eMLZYrplVwSWuGay/JVnutzQawT/re
0LeZmrk7ZxrkHGh2dBeDdMxS1ZkvLoheHtBxJZqT58LXHmQhL7Or4V2D0tZd62+hwG2HCbNAygXQ
S26kcKzagmMh9d8KaN0+8b9uDOv1U5p45RlopbdcxVa3j78DLjBflVjfjw2RSkL+0LMdpeeb8/Gt
plKKLyWJIxPcJ0fFCCFd+smnSHlmhqw7Y3wajCBMTE3EkJ+bXXTK7gvWQCEHCIR4eYHOJ0Q06o8b
72e/mXfEhuojHLYnhs/BwaOF0tD+q2daR+qloM0+Cei97KtolZ7ydvNKsvcYg7VmxsaLZ4TDphW5
9Sq9l+yyqEN9S/7bHiZpqubVtOEsSc7GhMAJTIg5KZFjFa3REATED84H9eSMYACdXCgRzOQrWedR
BH/Wu7XlZAg24RuQYqACEz6+4k0kKtclF51sxhkpoRtJNJ2Q2b87mVj8DW97+gA74qbdGJpss3/H
R9HM3aQ4jcEcW/xP2vG8tyH611mxliWcp5VdpZSFO0JtvQPugmQLZ+w96idPZ1pwpWW85ndSYBGn
fDOHegnjLFldHoRMYb+Fp1D7rZnOLrm/Cgy77rdunG8uN/MxjO0UwIxGQp/6c8TIh/va8TifrSKo
DXbZ6ZM9mxnuwFNabucdC8X0FHlLRlNnqL621UueTP/ZvFYpRRzawygNNfb3CHUvBd88W3lEOqr0
WmGS4wf5m+Qso8LXwQFAQDYM7oImgasyyI40r/t7rBNmJkrj2dN9KKBsLSoB9r+0sH0+8j1W1fQZ
4mk83Ss9CcR6ObHxJEF56r2vPz69Bl0imi1tFCw91tu+H87+/p5rNX2XC9w2twYyWeC+I1SKIXb+
3EVeNbUp7dSlhtsrHzdHSBY2dd4wdyOWbBYG1yiQbnA6tUqWTqd8WjVW1IS4o48h/CTYu6NhbUZU
eRLVfvS45VthiP+GsN5jbz2HtAz1yxxq0ExvEGQRtwKWWddjIsZrJxMUHORFUDYbRn7+bUBfmxa2
9d7Hu02amTvQDeiW4N3YE7arbcOsIqJ0Gnt05hUI7HDWcmmyL/fKw7Vy7rVbM35v30wCcFpE1hfn
mdhzQ3PbF9WmmJUbUT9TnzrT4tVnjwdY55MKUE7rrK3yjWmrMqeYlg+KMA6Ttl77JbHn+Kybq3X1
5CnQfMZafGMcSqna32IeEyzmm19MfzOzKFPi2DJuGi8MO2lHiBzqXhh8OkDZUxL7jff5s8eUvb2r
J1w6eyKE3ReBFwz+980Gmnxc4uEYHtcCsr6fnsX3eJoHTkUeus1NU4nZfNleY13fdstUFImaN55H
vl+ZuUXmnsZsUoJaukC+JNnbIdlF1JcRtvr/4lequvMb4kp+ifZdVBSo9iFEHPmZ6fh/gXWbuh7L
g5jv7gSGiVkmvTLVA7jNoHB0b3iW3YNewr7qGVMyV55uShtvKOczGngx+3/I09hXcicTszCDNRoC
I8KkO6CESwPSJ0TJINdWbyKYnwjGMZJxFBSlKgde+IHFOBGanoce4cEQ5nyY1Pv7zPtD3o20TP3q
lcXLUAh0Ch+1lnurkFKdfKIYpAio2yLmKSs2/3/qCh7BLIFuRMbqQ8DiYTsEiaWk8O80tZPOpEaE
ePi6a/ef2DTk3oGbCdt033F0yZO32GkvTUJ8rAA3XrVCP/bS9bOTx3PJ5B6kDLknl48j5m7Gq6q3
Gsm4r62kfQYAZwohdN8ol9RP3uuZwX363WI91TX3xU88bT3+1SUUnygifVlbBaJ7/QFXUaxgIJPT
g6Rpwx0GaLjk0VPwwsEhWL6OKZXFobmT/6p8edFI3hpoV0QBf1Cc7OLUeVjWth7nlgF0IYylmqTO
WQXirx4y4fI7um93ueYqpOfcv64EYJNuHXkur9RTCLbPu1HcdDNgg721sW69IyTdhCXHS1ilxJzt
vClFIHADS9rvUatyvf3sThrDr/yeRSZqfkebh9PqsCnLXhz8EfajkXESHIlADPVSt8KDJz64KKp/
4NX+SaiirRFixP3sl3FaQZf4SUgkytuYsxMRwKp71z5Sv5Z85smKttl+XM+fdjkFJlrKYQkvIq4p
IKBtBLaLmnrz1C9mCQJnxzNdrJIVKR1UI5f0S0KUXWKuNTEQpDh9Xp471WMwFSJRPGFmXCO98WmC
P+lEYcQRUCZ+QGAvYZDStd9PHRuIhYN0RS2Gb1eXESdA0/YuJ5G+jhHbnptZDI3QW/ssxPNs9L/9
n9tR7jaj8RBJN03nqZf4IZlDiD4LvjFcR5yUXeC5qrnMhttLri68lt+VfTImTICszSJ/eLjDSY9c
OkcXamTezLq5NMEvx2WqjpMwge3m1qwWeUkUeIo0EiRCEYRqvC0xGM4rES0E95ySVDgj01jEKW5H
3hl/EAz5ZmXHX6pMfZ2PW/xw0rOae3CIPqPyw1R+c1XT4PxfG8f5Yy5dvDGtoz4IixtHF6NDOrAY
CNDjl88wFenoBiEQ/ewWeN+DiagZhctrV0d8by0qTVBD1byjcbK7wYIG3R85x59bcxvddQx1Tpom
vnIS0PG2x3r8tnwg5LMq/kKYed31SR5p5FLUCiekdM4rRsCPg8Xi1bSi3bzuW4bftr1Tbm74wTjB
+Fgg9dJJN0QD7Rg6SJzzupgBZlSHPinIDkAVNC5HM7bBBLmG5HrmVXjaLvtsXNi6mSaSkXkKpPCD
hE8lzVjaDX4yc2HDkk4J4/gCmtarjHXdqJZAGcnwSA4WebTBycSyEZmjmJLujZc4gYmK45YXsan8
56n+Zn0z/IxYIfsypaizFyMLgFjER7a7f/LkWTsMNbZ5BHYO5tJBVRMQv2XXL3V0Rh104Z20K0H7
gqhZpVENkEBqE5wuGPGZvyE6NlsBHqLB6dOtO1hJM2Dp3gT0nQMS5LcZ89uFaOwoTtEY4e/+U0bz
du8WwQr9Xnjoo3NLlfuthDaNuQt7vXoyAROSCK+4Xz9T8GCBhRvfCLHboW1Bcw+zFHnR5l/bPwQb
C9UoD1i7VRYABQ5upJxXOYbpSl6MBsIrYbXbdBB9/IonWHlTKPuw9QnsDEdqfxKn4lKQoKdMNP1J
TU5bolACcaN3U2bOS+wyVFnG0q3csUwmjEkPDQf7J+PtAwx4ygVNdnZLrCs9vEEB4/cBBXPn+WAl
+pNt7jdO1AFKunbmuQrAjQvzIJfJKvfLrgCkQZRhbC/YlQAL74U+GmnR6YL0tSXZjG91Bm8eMjZH
eToo0knWhYnk4RUaXN+uS8y5jqxZXaO7BZhfalM4hT97dwDHRhoBZqhm7kW/OdKCK+e7GqTWJpct
TrFls4tbjgv6pEe40+2oJKKuAqgciMkczfcVlfqCRI3i7WP0w/cyIZraCqrAWt/QEd+fQFytT7vy
WOVIqccDZe1AQ7xtPgw+JAhsVPjwtPJbG6fSa7iFHGBuQXxqU2cm1YmBPBYeGa/cD2NchoszbC60
chcqIyAbjGLSgRESWx7lguX5VWA6omYFi9edWxdXezDrcrdwNaQmSrR+6fYlCkhEkmKoyGshZXcI
IW/+NMFu/0PchTx9gAN2P199RRqwZb4p4bmPsS/NCinnluhwNzhZl6cnPGrxDcPJM+bfQyFDlJ0A
9Jf+XaQWahHTqi5CozGyVyGJMF8e2MZ3VfcSKjIAU9U9a3ZadDW3xHKy/6qDGAz99J0ENcoywn2i
Acdh+ejOnQJai4XJoVyDah20R0vj2Veqogsq7xAGRrzwgN/WUnSusE4Lr4TVpVxEWWsUKxvtD8Tn
9Lsjo7bq3Nm3ee82MYhMksq2i+zPvr4OazYPxUnLuymDsRbAGvUFGa5ZV/YX6U10vWb6rZqDZ1P4
BjFIufD7KfbrfjvaVZgeaDZWHaEX0m+RB+YwL7elPRf0TqGTVdgdVF1BDgn6TfTxM8TS+N3qgeN8
IDVSNGx6oIXqriszQEJqzrlwZ+3It9xp8coylReOgNlNHM2MQM5ppjzwC02GAh/PBn1gSA366Tpi
tsSQVhs0Qkt3qbiASyC87rVlNQYsiA6jc8r11Q0aL/qpq8wfEtv2w5ZCjcuOdjd+UFLLtYWcFeR4
EuvEVfSaGos0tGKFLhZLr2hR15hbpGUIeJtgTO9VS+H0o7XiX7huw6KITiDp4F5ziVzRYB5mB0pI
5Ink+STGtPUMHwCU7MdbdCIHz2Cus6is1vwYBlSFkv8fRag36x75Udr+b/ivjT8sQ1IP5ocONU/B
ZC3vknxWxYF+0leWdVIlFSZFOSVNbScgUw2A2tIn/2C2J/dwSb1/LdVGe6Vk2XDJX+MStW6BCS8H
IMy6khzHH3NKe4Y3Pq3wt0/XcQFafe+von7DB7rF1avbjFguEFC5YYgJ38zE79DKp2rn7QiAeaTG
1V9nvN89vWs77lpM3okkqm4cuNNE/BXJ5lJlmx4xs6kgUskpbiUxx68vv1NS81eQzwnaqedcI20H
bjapI8/L0qnn3k3o1FtF8XtZLSnO8LmBYq112OY2qbnKAt1TOxfhDyw920ybz+9Ujr7aCcacJUKA
vlFzsVKx1GhOMlzhwOPI47uMb3jEL6LG4MP+hgsTLGhWszmkvZbnLJwKn7vye+KMoVV7Mp+8XYx+
64QFonsoufHyb3WWagPm1ph3meGlwdU1ahAMbzwk63wvdhdjEVogbwQ82AOR/Mwyq+LE3iDdP9i8
joPtTLX+yIXqSNAzbe1SgY8ZDViZPYhQb1tz09Y6FhlGc9wBK1VcZo4oo+YUDoDRhsuSccwoI8Qz
n6HAwxxW+IhXRqxvJvcqoE6wDpm4c2sXVRQfl4IrzLsGGG3tit6wUPproXsS185SR6ux9un+Bkb1
UVbj67aiaafOTK6XNvjqmvy0dF2pA1DUrJA2OKiWeyCF6NY6AbjvYGDmoz+HdrjY4uW5Y2737i/9
GAHSFe2LfLRO3TlkZeJzclFA+pa/VWcYyU1si0wn88CX1S/gjGtMx3/lbChk9V8yomMDx7NOtoaZ
6kWofwi2JEJyH2jxYeTGn34EDFOJG2yCSWz7WPMYaigiZaxthdAeSaIYX5F9NBFd4ROTbfhY45Se
1+pjifQsuOzMx478+dss/YwIBmDLB26HUCMNYuIy7Pf/VMpmi/filSBizeyp2YFRuSN3kcm8TcSY
lo2WZSS4dw5Y/8W9tBmSNaUQohQYN8o6QbyBmlQZyMFTSv4Y3R6ZWX8wFsd1jhCN0nyhCgmKfQyT
7M9umgCY974lv655iJbWpmhbvGOma+1KCTfOIUOtNSPGq6WUiHj0ZTZozOVxCU6Li7WmV8Mxz1x7
pSWVZmJadnhJt9jHeBQJtJwN3L59pUsKuceXVV73U0MC0HZB+TrFJVxPN+a+DaYY4yPfRr2L+JyY
sCcw/WfQleuxeSGu0mkQ9ydX58WRADnh+G96CeFdTstQI81AvjD8TnVRXmcw8DvQJuaV+PIdPwYN
/aBlMSZZW0Bidt5E+UphUeHJxMngrBE1XCLp4lcOYU4Cg4dYZ+oF8VQqwXA+PlKDmrM2nU4uiPtj
cJZWKs0SqY9qnLZUyjhAQ/l9lV4ItGG6Ebgn0ohs5QwjXjrUv3pZfKzRIacOW2GQt0uH24V41cKh
3/O8QY/k4lRTBM44llaYYa6oqilEiF2dd+0ZHHPiffHTLdBsJ8x+T/H5uqEuYxPkFWeHmnHHur0g
Id26srVqC8By/KL2b/YtSYLv6PMIjFpROTO+asziWradn067yRh49kWrsuT1sOSyzlP05GgOPdYY
YTRFkOEN7G7n9Wu00oH2lznfg9dtBqj8QagpiYeGFTKaRM2eL97bda3dNS26MYBcf+b0zCE4OjuS
8INOZzFMLBBHcpfsGuyPlA7HBY89lptmCr3b0J8y1f/dA0JWmG6nGO5Eq5005omZ3dfy/At9cQ3N
slnUO+Vw/MrDix1y1jcU+btYwLIC4hQa154wllwBt2hM2KZsyO9/Pyn27Cahn1tV1k3/bNcHEHfL
JjCiflnZn4u3f1PRsDeA7WPXnvDmFCqU4wqEZRQ/NOUWBpssPyabhUskhd/4KJgAGQYpC3bA2UYB
14oziKXf7w5pR5wZGyMXkxTA3Zr536FNGxPisPd59UMuR8fVDKCY+fxmb1FVXKUUKPyUOlr7h+Zk
O82Yz5dQO20CEIfKJUnqUIo5efTDnOI8M/afbI8fKuce4N2KwCCKEVUPq8UmiMkel9kZzDYEU/as
kjzOkGHUEkooKAkYAWpjbKd32J1FjysRN/1/1htTge1GXd4Mj5pBtcT09yBWuO5Fp66s0uFIk6KY
ui1p+1dFGMQkuRPE7qwjng18NzjbZK6h4Xkv1hL+kur+hXdgs1lTYJKhOPPVrsUFb7OYH99LfBCB
5JlCdGb8FIH28LyGfgBjwhUwvfc/Jm9mSie9teHkCH3Nyyb1s317K6oYIRtaYkvlN1uq+r7gNT0T
AohdToruZpV78joSJtAPJcAycTefcXJP48O8o4LvJcO3NhA2LutxVV1A7/kylB21PLqGYtBEc6ZG
HjLYgsJXpy7GqkpReTya3LF+qnL+AQLQ//utOyMDIzKBCjCfGZ5zVzefxQ4INT2QRRMwuyzJRq5s
KGx8CYtsfPO72OOj1m6fclF9W5Pb8Z2l+kEHXZPGcItQIRcOEZxqWWL21/x5CrofQXrBnYtZVTAJ
Mp/UYK4LpppqHTvWg8jW2YZ1oKo1iKhS3hL9GPEb5mKOCWS8ww5Z/USYyCVd1DmyszfkdlU7oAv7
qombqE6JISyfoSxZimJ7ARb/KhiF/BZ4xMKtAnuK8MRMPqBT51X03SNhPtEhRNBjXQHrv1KGEy3e
fPQbhEiC3OAkn4WjS4uR+/w4NSPAfmeMPqVUb/2QuQHpsX6woh8cGiyoONrQg+VcRLoi1t26L8d6
fTKbyZ5v+yfMveqxIo+TX9emHSx7g/kTIvmoTL1ZVjScpQsiCTzFxF2IZeCqu0Tf1ktPrv8AL8SR
Cms2gqeNc2L8lw+mx7XlYhFUju4Ybu4hUUadDLfMpn37X9nhw0MCPHRTZiLt6UqtGH84qiYMnoTX
RIkQOQtPVjcsKU8P8GAKP1tYyeezGPWgH2ctxiunATut1fIw3Sw1fsQhybO2+Ilk1xBNVu+T9Z68
HBWp8VZT+4PVgVeonqT/TgecO1fMfIfYDEtpYMgNpjGN+ow5C8YGY++iRpFooJkZRekRAiFwomM9
IggQW9EzbSchKx9kG3LeplLAkTgNNFc8DIyUirJCzJ7KhNNMwviRcOIaXvfEbcExvhVLb5Z93Ict
taGyXuuxOF7WFFqYwLU4DhGE0U8qnm3ooh4ELiJHvDToN8trDS1thsUMGgPyGHd+/Hc/MowwHSJH
qATQMqC73qNmj6UH+plUroQRWTRGo054xaS5nf9zN8iqVdCSjDFyr34aUebyu+mFq9pDcN8n00TO
LvAiXxDPvgs6o0YdffzMYex01c+8FoVj49ds+FVGYWe81Ry11/zThvdJeRvNR0FxHJ5szSpxUmUO
AXRf1Kot7FmYBKPCzjZn3SVGDbmX1leaSGomrffP1Inoojfbnu23eWQejxDW7BAGBupY1ssPPAYc
wKJX7ywrnOirWwcCV/IJ0XQObHE0jCpa40DL9WweQhM5f1GGydwomh6wuuVt8/G+GfCnnzEAyJBZ
Am6ig8V6DREgQDx/8p8bfwRkGhteDKTxIbw2//8mNH12YwlkREw063BvkUhLUmHhDOK1plTElqoI
OnPMcZwWwWMbAofUv1mMiDHELVT8RmFfddsIbYjByomz2sJzIbwT762H9ZMLjtGg80+mw/ZVtm1L
ajOOTGeloJftLujhQb9pKdNtZK19jEGgmMdgb3jqHOVVY/C3fHIxvk2nLB2g/EbrwDcG2xMqoFwX
nk6jvsm8MWVn4sxwt1JNHOCrs3g6IA3X3xxG1+eS+WnAsezE8UrluV1jGo95AagYZ9enGbmsyzDu
l4SOinGcOOmWjDL1/ttx2bfwwFf6TIM/nXd7rlxVojm2BqX9iAOU6aYJLxpdbfsWH6p5Jhtx5LGm
CCdufRsGqaZJOX5w8iUhDtPmIOxKSUhvyayUI5N09/5nezzbvqq2Ma7wITcFQLhzosmPrJgrZus2
yHUu/cNL2XNUXqpz8nKn7t0RU2X8V7sqgrDRUM0kRGXtSXFsM8xhC+x0nT7hoXsq9MS24l0jVu08
btgBp7lq7uljZvuvUL2+9OPqcLbw8HE20jSNvwQqceo53byInQ8uxXJmrJxAg6ywc1ekg2bAeUPK
zXqQkIUVBpmnb9iFfewqX+gAYYVPYNUlkbNQlr51pezlHFS7VyRESpbJgWuh0hCtuyHVv+/lSZik
9d/78b9B9rH+s6+qrXNsvcBRO+nzsnioPta5XN4S6kD6eaOlX9oFMSVj4WTyafnwD0pYx4L+5QKN
mfo3odwGhXFDwio3WqESow9rsx8JsDu23wSqBgpoYBqo+ljRQRvlPFbobI66J5hke+4TPnyHwSqA
kSmoLLzECeXbTvVmY5HrWiEOQvnPdE+471w/AJDa9sdoD8oFQJwP6KVPAOjlJA9KTGbZ4FunMxsp
ueKj/mCegU/WBlP9H6Djbw0LJjULJh6EMe2X6diaRTcpf+RH2BxGtQOSjRL6y8tN9JZpLo2JMPeu
20Y0k9TweYNwUzv4vGeFLwvqOPmKPi76jt0AzVe7NT5Uq16PfHblGZPmoZwEJKP09XEYyMe5s0UC
GeUWLop9qoCCaKm0+5U37J/uGsm60VFrgbwqOhEjza59ZM4lUQ4tAv4bacNS0A+4Pvt49HxaIQV0
r0xptYE30YJVn+n6jFAg4SWduAMfWbv8wZMlt/RHsIgvPc4Z0Xoh8iDugw3qOspA14Z/mLeOlg5r
+TaP1IHM+oln/DdSSfW0SCGSHgcDVsqGPo9etUHTKWg8x9489ZZvnEall6cdFOqLIS4ahx8QEgDb
erc4Lmtwhwiu3l54AM9mNbFt25Ews7t7Dg+ZzzWMf5JzRb8lCvkB95SZOIBl+WaQiFr0sUiSWFAW
e3DwFBByngmJw6hCI4iZ7dRXnmlbMY25RNeMlr3a7iyzU2g2EoQp9bt2IKQOS9pD2iy0nAlevZRK
xRxT6czsPjlCtWWd5JnsAZ8BMG/tTksnVP09U4kEaEj+dYucn3khI23CPehuHID08YftPGyFAVTX
o5HCyLiPn+eRgc7Q0kcJd9L6NjQwuRQnPhc4o+vvh/QOn1X9N4kLcfLXzBLg6Zm9l89GEuKBWSkL
9yeroaEdyvuQVwAhNHKOiiE9KeAdbHPykGe/3Fllyzq4ef/2JHHk/bq50g862ukGgN0tDJsM0rgn
VKuCGnZrJOE6QtEVqobPNggnAO7z8RAGIKQv1ksbz0nhKIQYn/aM7ONaUJIRk0PkXE6liumI0Sf0
7C8d8YbFi98ZIA9CfFKu2T1+o0uJ+lsQ0RJle9Mn16YXXFaimaeel+8C+FDkznBH9eoxH7vUON/H
TwX21jE/s8bo5hwGaQqsa7CnAZKNwnvMeR6wdy2vltHd8w8fQPoBfLsMZWs/DGxYricMM+NxIXRe
DYkhS1sRAyRH1nKK9wStdzptP1ipQvn/hq4OWYOdc455b1XQbKQ19jUZyBhOWJbXsRfGbEqRMoQn
8QsT0LhhGuPF4FyGzR++U9A+S2JQX6S2JrvNWVD9L9EwQTlYJRTT8uvbc9crGc2xSnKuRFd3YYgF
/t8VKLIYgtOKyKz2gVmbHqqCNxudxbq6i8Cakq22r8nEKbV+IvEpCDl3fHebHrtTxnpLjbBBU8Sj
7d1qQ1mHsPwz3Ih+OnunyWF277hoTeK0YnBM/WWVX719QDbr8mE7Y4b9xxYl6QfKNN3WGJXv9tl/
nOp2axGsLRwhNP8rT85sgy3osL5G0ZrE6uJAxtq308dTgodxhtchE4vdMDNeMizD0uebNn8s2GJN
hvfsPjwinTmQFBaqxggJgKSv8ij6jGmtBK9elEdN09PeXLu592E3n6T86tGp3szzEZdBCko3Tgyh
sn8S70slpZnnN1dHhryu4zbyQZ5AgO/WMv+X8N4ZEz1pSKOdRvTdx1Z3DsBBK7aqnqUl80Fsv0Ts
GQCHWjB2kEU6sXyLK61JYY3JnjTHzRlNFB8Eymvi0tVhQ4Z8DnN9XSPnJOVFkM4Eh0q+nVTFPTis
QeX8BFDWRYuX0KHBNubGPzJdcxVkj+L6XL8M2YZJBCCAuhWCTzrBAU4jxP+KIQq+oZ/3m2bi0JBj
jz0ew650iIvgZIOoeFWmBL5qxC51uPU1TillA8eikCLVhu07RfR8gUAlYagMsXOxf1bnlO0RkbR/
1qRl+JX9LIDnz9WBPRcwbMem6OlpR1REn8zIIAdt/y3PIwunrRgv9dy8W1qEsOj1cyH7trllf2Tc
+3fbo+wr3pjpTDgTPWhJToiYzjPZONYe5nVeSmmnEqltPmei6rvjkkSuYp2ooUREx1WqpLhZ5zkQ
5IlUpIqhp4Gd/i5K4cNeC2mb5twEb/xgIWml/1p1Osn0cfu0YEVFjOL+cRuvUnx+0jNVyULamHg+
U6ZcwECkUvFTBR1eYo19cfx70f3uSgkOOJ/KV1tSygiZ1m+Fhv1QworVlFhLU6QEEC1w+GIjVq6p
EHPjZ+8khV3yEGm5Pk47mf929Ljx20MJ13JjO63nTMnr7wl40oemGP/FoQZn9k6i8UOYeDTMPP8W
KCXzTwfZV2eg/FdKt0CqK6RfAnNzVW56JUOsgPqZRA26LGYNxh+rHGxYwCGkw/J4tb1fqHv+NDdb
mhCDI6WDEzX/a2sdma5Jf+eZBdIGFRKa6e8e+k4HxC0JP4WWmhXMJhIqt9bXBOVBmDNsn0mANBCN
aTDYjqb7Z6bUTWhCuYffN+IxuJ6pwY/fz2QW0mwCZQZtCaftROYCnI759tfwlJ/XbPKkjueKtycx
/X9Lnl/Lk1Iur7Rhr0T1Q+OluTEd/fpoTvmx0wncdyb7qcIWDKDn8G+55UM3itDtTHS6OyfZDxx6
Tsd6jkSK8/j5xDp81O4Ss5hTlND+jIv+68fYH8AS5SeqJAipMLvM76F3YC0xqZUhcfVRaQo3fsd5
xVwV+wGR0QNYgTUKoyqarpJcyWqJicWg8Up3t6URFT2Dj4XGIw0LYYDiyOhz9LcZBmqT7EU0zazl
VIqjAh2qCUl9dTEVqtZ1rf7NdvZTuNKsCFMx9Tgu2JZAMytrAe45rRjNQ4EEZ/kDevYK2fIpv3wy
sxsHjaifYpOMzZsU7VpvmTc0Ca/n/QDihl/HLT18oINFUhQHf7lLUfItSdVIhmwHjM2Va12m9BJo
w9pLz6KNGjr/Y3e+EhbgjhSMzMyIK2c2Ci70Z1ixKFtuFfIFfukAt3x8RoadEGE502As6TzRDwIq
Gqk0B5kRoAdhXMTCzpNw/ITYUz2jtvT3hDrqzuWtdGdbj3ce6QqlJChpl/SEpwU/65Q8ao9ZugOi
qvII4yfO83bUrvlVDHeBYNIsPLv8vJM9kA8dFMRPOG5qbz2sEjV3xfnd1LCpiJne5A/KVO01pkdP
Va2NzjdH/MhMIx9pkPXWRNa5H0rAxCqhp6CDqvfHkBwN/m5ve/i8jtixMW3lvgXCCxZb6Ck0qmvc
XYKdcKZ0FhfRXolu0LrzPKw9Gw/X14SEZaHvEk1uGYTs6V35EZsthHf0Mud5fLdv5VNE8giDLngo
XxNTcCPbtoKeMUNToiINZ5SpsYQ2t4juq0t2ixe8Goz2hFkXGtHI7suRJRf1xBOjW1pARfyR1tN7
EWzcbthAxy/gQQrXY9gckRMDrgFT8Tb/6OeJK1qZeeqfeyQtdvd7c+nLt3qe/LMCXbp5ISTRbSS1
cfqiQMH6Pa8s9Symzl8koFTVM+Gw4P3YPD23SQAW2OS8dXPtXm7QxLKJE4Ybcu1vnbZrufCYLHhj
YBXjDnV7a/2R6XKwb/J3BeTDj1OicQ72cZIwQyBgsfdLsKSjst6ea+Pe+wDUJCFwO1LVleDyMMnf
wzz3HC4KOdcMe2dj85Te2gImkprze96q+5X2ygvJM4m60evAuqv5WcHxT6MsBEIzSNhKdOI4QPCt
HlVJvQ+zLhy+aJicfhp6pzTyA1MLiqH5SuM3aUxZ4uNQ0mNh/tRvTrmxXWCFD0AzXK5phW4VRmtD
c7FSv2w+7koXZo+dw0wiufg1I+HNQxFcxYyNJbJvDDg9GfkC9QOfk54QuzMwU9Voe4vIQOuy0wX4
acfVu+fDZ5n6DuMxykZOE1BTcDqKcLwJntuJ0jDQCP/SFgOi4KZ2sp+J6Wox5XS6Tu0eHH938GTd
ZkfsI5dErGpPY51KFsNqkvCxl8OrsiDkbaHO8GNvYXOcx6FSmpZ6pMSVaJ0q1PYi2iM1P5+nuTvh
gS6URVqBiKUhmkFLipT4vH2J7ngliwai7cvL90ycAqzDkFl9Q7mP1s155HnNlofSbsUdtNtlxKp3
h2R+OHuq0CsNnp/SB4I2ubdd+uN1xaReZVuR3mt/Ta/z9k7mZMZgoltUancUc4tMjtrQvelFH8PV
Pv28YiB2ysNX/wOWf3SSB90umD9OuPw0OMGwhuzUUnDcn+IbOAO4+L8sBwOcyC/nm+WtL2+7L1v9
v7YkpjqKrHjq7j9HoB2qcI13x3RfBKUMOTnWRKyg2h5oJDnSLY9dPqgm6nRy13asl7ur4umj9OoL
Ka9Euc55DIqD1bP7V25T05X8nUoP3D6MrpT4/S0dRm3m0uJ44ewKIyF7C5a5L6JRLH3LjIo6AAdi
4fS0WDsykr4FRFkpHWjqFiSrTbr4hBv3Z1IgBTiq2ufEvasI7k1CrzEEbk1B2pkxfeV4AhsJ0jY0
TOHUSC9jKi4KoqbpPVbxKMZ/GhOmZu5DxTj04qid7bYjkAzwcRteTrzIf6B7W9WAu1g8W3fv6QhV
sWafvlK4y/OpSmNUqu4a+NDlI9pkUtendtV9PBwa4hl0tKhLOKZkQFwoVjX/oIVIw7rabQGUj4hB
Zrwp0fmSaUnk2iZlX+Bg7fKqk3IuaQDmQtmPd5zBlhIz43kDfameacs6mFLgpv1T+ZCrnNkHejXr
8FNSAdQcvsO0a5ffmM84eEeZvR7ZySKo5wGSEMVCXdlLPA6MSfb97yNuliSi3fl2xz4s0YJ9x3fa
kghTmRw8BqY6MIGL59D69Vp6p1Bbqn90sRjq2toWYG46vOJmVmZ9T39otAik5WCY4jeCePs+YrXy
7RG73Hzwj6CRYVgt22F26bBEnKiIwCUW6feW1eg1tXDsZcXE31hDJ7W0XDMemzXknathacWXRWjG
BwqmcOM/bvane5NRCFgTqkPK6sJtPylHbzz8ME6r483cW8iXS8CAVhcWnaCjucdyKfbLXrwotIEo
edONq1/vcoBqMmuGTQ1ICbk201myjSTX0va4gM5jxDEyRLx6+Qomor+aJI8pWYpMgymUnkwjhal5
OJtS7UEDNDH2+NakX7Syeb5f2lOnQxlScxKn7/LGu9o/3e1eSvW44KohXzTQLqSdmp/ThuwP/gqB
ekYwYvSZEGiYx3duKkB+AVn3Z37DtlD8Ppopax9xGIqk4RqDhd7bZGsqXicsTXM6PgqVVg3NYn4s
V4A1nkFNpHL+z95pwZAkp1R4YtT6zi2L3yFJnZsV9RGt9MnHKCoSxzHHVxE/Q/MRn22vo3HEo2x3
NMKPlQ3tTyHd3obgMbFzF7XFRaxI6KKu/v/gYXRg5IdX8PNjFWWmYw551aDbFB3mTgKDO+8dPVxU
I8wqqWEdrYqyYuz2NLBcYi5MakmOBJbons3gXIB/nohqNsSA+ZVDcYI7a8Io/ls2qkgX6SLDIuc4
mknqQCzRssAIlQuNnikw5E+63mtZ0aafJnFDvBuorCdSyv151BDePibt3ZqdXl6Dl227JfUVE9DZ
ZgSIdAdCpJo6Bx9w1M9zON178/DfjiRlLIoJqqqVQPQoblEtpZ/8BXuwYixZXfMMIIEviu9LHInx
TgXNY+Mpf43fEHaJlcQ2XN92drzlL0aFusnMAhGKIqyo6W1UTHDnrvZacs87gG3wWLLqFSZE7l/z
W6swnIwGEUSgXTbMJ2NAUONPE15/Khma5Fojs0atJzSq0jKDJR9LPRF/gyMOozoAkDI2atR+lyQT
z1igwIySR1BwcVHf48q6u/BblHdldC+4u8rsksnrGZxZ6aEzz3dKvTf85d9vOG5YLWKpm7qk6KmE
Y37yzgLdzqdTaeRuO5BpySdPGTh6o/xw7yGAjOohC6ABrGr50D7CCaXP1g0AWyFqgDs/5WgXtfNT
Kb48JYaqjsO/Hx9W/+rkzA6pEmY0Kjz2MaUHgCtkv/3pobMzO5NhK+3AFJxnmFqq3cOLCKFvVY2r
fD36+FAWSaU7vnvQxyMfRRM3sP1Wzap76mbh+rPmFhIxts2h8ipteLKMc6PWX+bzGqR7Tte/qrW5
wPY6Iv132almsV+NsL+GLii30pYscYRiT/ctFMR81F0aRV9OxktrnYZFbcb6hZ51U9fkqAvyHTAT
vp53GMTmtrwAJGEwFK7EHe5ZbHeFv6Qs7BDl5lVvYTUi2sn2dMqPYscqAYK+/OJKh748slVOSPWZ
fwSJO7YZeAZxZytLesv4K9r2h64o/1KTsQGglRtJypXLCcv+VlwjEomaNLyQB+cEsap4Ahgv0K1y
Pkg1/6fBi/oCruyFdEepGrRPGQBjWevelyQD3M/ELPSd+PNKYCTbOTRsZSHy9/0x2zXUTyKkgXUc
ycZNNXfMQfCBm+tJiFSYJG6C8DKJQ+yWsz95+gURIugR9DFMbkSlUzd98thCyxOX/upfH2Vnygbq
nQ5VaUCbZOM0Vd8GWxHXDDtSp9W+gBhuum9ifbKOJxvuirPSZYNWAs8WGGb5ZO5wErlZANSajGdE
0Xc9cSoTUVjO57Di3mGroAcV+YYkoxxyatlvO7xkX0bQOgC/TNr9qL0TeYF8VgRnO8ZUvrX/uz3n
xt1KatCvSpEwG8NKqI9JdOxDEfvj44rZVkB8VrlF//GdA2zi7dXU52ZAiu3RbGKMoLxJdY6v23pP
cI1UV2xZo8q594qQHEWENadXLOvcrqv7yZqvSuDfK+fB0iJ1S1hu5+j5QREbeuN9Ylq2rqs2cSoB
R//Tmw2n9iRWeBe+gDgXDefoLhNzkayDWuw8g+kmi+2nsAbNSrqsqNfIXHpnlTzfpqvx6OKIy9D0
ni1OyVnCKqBWrycQn5B9ccYSh2QhXyeyzs87r56i+e5nHpgqfHKhYNHXUWXsWmPwPSFS9EER3If/
41rHT+Qmp9pouWcp+Mc0QZx7rlu4rNpjkNoh+JHOl/j3BO1v/aE7TEGzWZaWiJSvAyzCQeZFqpUc
p9RigUvLIltgfohCAzCEiApFYrOPBbyJpb+PTP7R9UimiYJ/TrgikiFw1thsv2hWI54Ggo9DIhGe
7Umfk+b6g5XQJQMEZROCuHn5xFEAk1gqjLTabPk8zlb8bp8vk5gNO+glljFfMGCpMvJ61ugdagCV
lYYpmOhejaa21oFjZs0CGrk2+e4vgXGlQD2D5UwW8F0EMIHuHRDJPq1mDZjEf+QQmDwbxvnwt5r3
5vJO6jyJDJ3vC139WJGQ1lQRKUaWs6EVoj0fGMU8OpL0Tb8SqVOfM5tlBUYPnaf+fpFwpf1epzWD
PPKOfsGTYvjGaIh84LT9qCVMaWmugJj18Tj0y4cbaTlMqYySnFUexVWhqSMGtWijfXNYqOCF1Xba
No/lQYihuY9DWoXE8l96/oUfMAQLDkjye1KG+KC0Ft0Za1TrsJkvM9zSXoaqzGCqHsSdQUTyRiPt
ozPgtjac4BKzoE8BdFNG4BvTA5RflVE/b3k3q+79rVCM50/H5tHF8oWmKxFWdVwBaG2D6Ar7DksW
pSfPRO4iwQOYbmR6T7ectwrWTw1Pp1FBiCCdEKDbIY8ucizwS9X3IV9ROAxXZpJFSf+QxBhdGYLK
Bzn4AuGcsAVnTo8PMgTDT7nBn5eiKbtRTzOoJaPDC+20k0pCt7ExFR+as+8AaGneT0YvAjGmhaZt
sbsW3OazEGZJlwAsXU1/LVZ638dRrHfOzGYwV3VB2eODqPwZKXO2hLA6yPCSJFtNzPw3bsAcvBRc
N/paRnMEyi9DZ0ylbWwAwtvZTnmo/o8wzY0C5qdBOplNFP+nuw++PJ8uUZg2qbnIpQyJ1Ki2TZIm
Hv5c8juG0b31DW87Jh3wJTySDzRQFFxcWAQQWn3JyLriGV3wYmeFy9gdcrzlAsVwapJyAuyIbML2
b6QW1s6Jqf2CrE1I7sPMFl12fJkabQXl62VWEaadwtzGMB+xmms19QmwAcgXsALmOsBiG+xrxQAb
Ms5PWGUCQ3tuqzaQPTEFCeedGDMmYLdYuvsU69+exd78NACERRX0G+OyHUWVwpzw4heNWo9TRfau
sgzPwarRGr8FgP9w8s95R2RwtwEsmJNwNu//AysXxwuDMfRX4Zx4TzOiO8hZRRQHzr6cAo/NjZdT
i9zdBkjl/Aq6UtMgG/TmkGMbGwJ65YWyI5+2rSA8xgx3LdEwli4aSfRg7aXEb4ZQFgtEL9cW4+Jc
iMY/zNAUXvy4qqID5oE7Ia0dqkSKcdlC4gadhWBGfUPXh0KRZXe878nLaYmZD6dTAih+ILREsKCP
r80n8wp/pAFQ23Oq/DVuPHuBFB1qS4h7nDQSpY4fE4AiYA7I6VM7i7JtPiwLehwJORjmwniFBJFq
ApTvEoldYOOGbRL20M8hhD8O+VT1aXmGcgCcK4A+dMB7fRg1YNqA3UM46Rl9FVGDdRWP7wWkFGui
8K1IaAGgZNOjV8NUHAsmWscoBIK9WPVnx3PAnXTHSLUcU4IAlA6KgYPXKOGgamUhKaGUED2uyCq0
RM1g0tjVTQO6D26fmy0NBLhZ3oWnu3qMA69M9CLHiQWAPpMbhSOG5rhdOjl5/hisDrjKrm3/A8Of
oxEzsR/dtLu/QOcxNjRJkVApnVhUzKG7rApNKyBFPGZpDhYvCVSNjRYzxSrkQFXcMv4IXWWSVRNO
cWMLI9OfP75mw8MWbGijaL+s8D0QCYqBcKp55tC4n/fkQEAHKpZOM+cbT8p+cxFaDw6sFrWiggao
rupZr75P22Y54+sVSFvgKiIOYVZlWOWFsYdpmV7mZkNSu0Qv1dNjsa1JNJjsJWfCmu1aQW2g9bfM
+y0JfU4TozElEQjsmdF5D0Tww8miT5rDhkdE3g0mQXvhJDAc/s+7tjKouFGAKOA+bva0kIC1GI/R
ewxpxQpfbOofo1Wjw5+dHleFVEXgyzPIlK4NC/5eNEoWEfLpEFSHkEqX5CxZT/keTd4Z87CTno/i
D7CXlFZyVV5a3Obg+sX/Ioe2lAX5Nj/PdpQ3Si9TlLL70KuQZrygoF+QM49pYMiIXNqO6lSpwuDe
6fhNFK5+rvKZ4oLNciv04ZsGNe28NwM+tzXZvlB+0TViMZgpnTUgzMwMPqMTrM8mU27oFDfedzaF
QK/c9XJEGL5636TafsOoGiBLkET2zAfTbMS54qcUu1dmeqm3YsFrclhmfoPbXl4gV6QEh6wefg4s
lLAfuvUG0DUw8YclJ9zgUG8vkh487CYwZA16xEZWa33aU5eq9MrtnKJTdQS6dABFfDpZFZzHTzya
k9Aemmh9I96q1bp1pVd8MdxlBcmPWMSkWBo6cP7/FOXgCtSfeTwwjmeY1oXXaAWNgQ35b0TVLMWh
bAJOiMS2uy+JjSNxOu66t3jSuNpHkYdHw9fjgc4DjPEJYgf4BNGn2OaP9ZiRr2oMXymW8QYpmqBq
aZK7ZdGeQM72IzCE+Qb1SuuLlIeAOim1mPNQHqdDDk8mUE18ni88iH+PVC5/+6aGzdH3+zyK+hOC
7MjHyVIGxV/2/JQHQxPMr6Bc8VtKorf1U85inRFrofDpg+BirwPRpJ8FKLe9+ng/PhkJUcsNYfOz
xWqaGLB4uaYQNCoHE3omIr4fmr7We3KS1XEdPbhJjTqeKoqgKeXEEf1HOuUnOE6819uwMfJz4XoX
KZPt4lBsT4akCG1clTmLWaTspvMKL9baj3xlKjizYQCqumpc6jeimaBcB3zBslTuB2DZJoZ5N1oG
VqCaizFBmONfPE4j/e9VCZ6jSPJpF27yl3tjY6n/W7za69J79HFeBeK8O/4jHTO+LzHbr05mvD7Q
/V0nvG1X3IJxwkwqsYcP+PA5kfxls8FjxsFNIAGwELVhKH9dkhMx14VHjx1/bqctQA36IFWRxmzz
ZTorjgVcvpVMFOzzWnjU1l5Y4l/UJV9Kh7yRQ6/bA/jKxt2cbGT+atezOkdZ1OhnSz9e/sPJnllV
W1naiNgypvxCAHeZo/gb2rm/f22VxJA1u+XxmQ0QxsOkMhDicTn2CkaSe10yWqvMLiNAQs1SCDIm
sDnpu0dihQ3Zz4fSXAz9n09yamr8GuosqEB9HrPO4Djsv7AigDGcYOSHOJ0zQW1pHLXo1MJ5Ky7c
80Yjk+Wozu/4t1TOvAf0A/jQaLnS2qFdE++0F+f2GlWu+hOmSJII7VVLvsqHTaTNfg0xVOJOf8qI
8FVlMKIWYLWxzxgxfD1i8uk/ejzMAVPgkobRarXomc2AnEUMxiR91H7xpth3Pybt1xArFYwfE8r0
lSj4B9pzHAn7EqJJAAA+UmtvFoxBm38lb0cij9kuuvCgMeUoZscVOU+qkoT1abtVZvnrlJc3Arci
HnsiEQdq+PEiWkfHenpYuD6dEQqpcAYodfSLr+qyx2xOf3ciSI/ozJPnLocg/qa7O1mcDlk67bTs
l93RcOFtbINS+yiDyoA3EyGNRVsFuTp+RTbyJ7DRf31GvEB09y0e29s8/8SSEUMaTAiJw2Nxoopm
dtEt8n5JimTshVDYJs5K0kvEEJg/5Ej/J9LUQP/vtkCxbDyIX7zE86wOW9EMmJY5cDWnrYWzIVCU
9RSw9TP5ZUfowEYvWY+c26Lok6esNBZBgxcn8kGgrT5FjcIaSsS9ynT3tm7hQfHp8k+DwrvvQdqQ
FZIuO5tkW7t7srdk7Z9tDflVRf7uKJGceJAaNJ/ILaz39XA2/IcQawjiuT6HOeFtDx0lYdjzjzAc
KHy9OdgYXNSqfpCkJcR4G2MyEET8EaamgtFtHTainrYCYSKl2J4rTZOZTSCt7q3Tp0j6GuW7r/wS
TyVj2dFPxQwRqn9i5k5tkHyFfKgxpOisjM86YK+BHoABrq5GxxdyJE9LbmzAtD22Vhre4ecs4SNw
Xn6dzb8nyx7fCshkjMMI86k6H47WNCie4mtMOdupf4qmfJx2Xg5dr5yLTs4d3Euerm3XiXDKewRm
wMxp5oODuTGHmTh3C/zdxV/95AE+qQVBwAgMJzNf5d7T0qDEqbuMpdPcUYTrEnt1zSH8RG+hPLsn
sL/Dd1qJz51yjYlAhBTxYGkS3ZjubsBiAz/gUO2k8XHb03PXHM89jfx1jarD1wjVwFwP+fpoMsA7
JsQoGvtIL2m/7lmtElWvD94NTr7tOVK3xEn3NDl4TDEsPfrg2pRRxV/TLbTR+N0FZWjsT7uoP+Jq
FzdRPd0XtorzY9J5651BJeDCAUxdiyBE4I7bZqFaStVXbeTlanl26OsF+3M4IBcEqT+ZlycBu6f0
8FRVK5gF1PW7TWe4dMKbt6lCdp//IgCrD3ep7TFNV+Pk3xc5v5o/kmvMBef0D0zzIePkDr2uzI5w
ol0Wbi8l7LpHdG8L+cAwgcHWtJOYR2BvpAvBkjhM7aWVHhgu15F+u7wemRnWnNL+u5eBiE+zcIrj
dzZmNk6ub0jABKayedvxcJ5otztBtYDl7p5wROwYze7ZIM2KKjplMAGiDVYfxfKsKifQrTDNsHtb
gr4/f2GT+AkrLHZOt758shCu5AcRfaPLfdwTEqsdtWHgY+7zSIwipkbg7bEXAc/SMfokMxNB8s39
F/0SwTKj92PLyJB0Lnl6irX+we7nzhDmn3GuKkVsxhIanOoYlKFSBzoPaXg5IQvIhC9Ary4PvfL5
QNbg+U0d/KpuazRpZazJBKEAqlEAlUOqIMxHmUq0qnWxXr1jgM55JjLnYhFwDkRYEJoVhAJaeIhy
ZMiYzTJoe+hSEUQDO9Ybv+S3H4rSs4iM8w8pTBSCZLcW1GDGk/6g1Uu7sQgBOxd88/ZWAiHi2/K7
q3UU4MfYnXyJAsJdWfcZyNgdRsLeGHucFVg42QnECcF8K61bQCa01DyBLowPBh/YOJu9TwmxQRYC
ZNVQFGeMLGBO6XjVOnjLozgqjgWD82s+Zenr9QenWbq+28IjMnX/pL5qHym69kSuE7wjBwDfK6RW
bNoe1mu3W+eUAkoXRuukXUELRUdm/TkWnHX1mqLYkW+3pSbWr6hddSb8IL1py6GKLrpXG85NsOwN
NfAdZv4URmchSDRf8r9tkiJC86Kvzyh0jhPfAfPvKKk9mNCXP2WSNnEm4pLiRZu/ZQNIexEpYHDn
+0N02iZAdQHgBv2qvHM+0yfK6WDbY9JlFKUAbiqfrvW8cZi3rbzlU/q1Sa1FXwcwVdbrIMSBwl0L
SkCAb217xK41u+pMwRqHddfLdSKbQZggR5DSkw2x6ewQJHIGp+LihX7y3Pp0KOmpiH+PMIocWDpW
bZqCKpSZq5giK9a/em9QhxcxBQy9qbf+fhV5TOUc391Q9E+HnCfcfRS1mJravL0/HPOhsD1HumCA
0OFDr09BMgOH/4eLV3oBQiJSmtOldOYOnR9RuJyR8YEUuYma5IrOd8ZG/j59cHbkyGhHjH5pK6rL
bnH14ax0WsNXRrsiqfRg4F+ZXjmNbQczqKNkmEMUulKernPtBz944eQFDUMKLFO0MlqPRCPsj3cG
V/wmrx01gzFG+O+vf9nfqIIHX4kCAvQVstD91Q/AaCxTUJ26BNfe3TybyLAR8iLdFv9WD3ZgcYKt
tCteqQprsIOOvWDzC1n8Pa8XmxhQa+b+48EIGa2BpdPOetC5xgQlXdUv3VW0uTfnjv0xt3jmu9or
nCV9UcgbcSg/LVBRUX47d/JyLYoTqMFnwiab6jzXOPMD4ZZ5Gki1oq2DSZDXQ11YXUXYcVXbIZbR
WESSlE1NnKp0C4B8FpRV1D1bK71ocNQTCVJaHkGadvrzUq2wxsUfUufDA8VcBz27BPJ54rDXYggQ
kZPRv0jNWPTi7n6gzIBwXQ8Fum9PZ554GERNrTHYUR+gjchWh8wRtpY/belWyW2I0FR0/2K5ptbw
vDhVWQF50JqahwUuKT+L1ljt4tThgYBUv2WyfLC1Kw6FsJPAIFtuutwj5noWn7Kky5Yo7ZYu11du
gootZXjdqVRLaMPQZEFVljFtcKzcOWD5vv/55idLfq+Pmz2bp+uO9wo2Ur0oiKlCAQEoHVmj34ln
LLZoglg4VOVovY7gvDqItU5ekmZ5HrFyz7axNCLPrMhgdBIqz/og7saHLlNA5XEotWqQAgT6wAAo
rb+6zfIb0+dpbvo67srnY/2gJjOlPNWVES5mqJAae4+lczlTTrvgczST4+I5c9TBNzVbT0lD/TVn
KB6wtMnJpZ3D4wLXam0UHncmjcdIjxJDsPyCZ38IJV9SyoX8HPffju54TV2QvzfX2Aw58sluiFLx
QVKAwF/ppm6JLlvCri7yxZ1Jt0M/xw8YYJnYntoyfUm/EhLumn+G7yIlLOx5PW94OQm4Y6KZwT/k
OBN8N6TV+FJnwbWPG8mSSmldVCEsH9bWiZiC1r+2FNQ1gGuYjiqj8M3xgKYs85c7bvBd4N5srnM0
7u3xeauZ/We/eKreKeVDIa+ClAVwNoWf9wBPgtdBKum9k0zwsia6mTMWpbCdojn8VVmzyIlVYe0V
B6BPQLOQEU48ssy4z6LHmPc/dIJnN+rtNsDQ+UbFOIpQiqsFrKeeziSZrTNGiA6G2bj8liEVzgga
xmO5Hb2jmuhD2+LuonpRH6TpecGvH4ZD2m53OnCIYYP12ZaDPkjU1SOTwyH0wl8bbOrPopT1TXPE
QM0WdXj7yZNdDoUWJSmI6rmzS9RxSPNEYw98tOlQyL9r/z3+x1eB5qocycCCXkAP7aKsmskHfyqZ
EI6exgzMXMzMtYeaR7KN8g0wETK8PRPVsU973JatZM7RbSVtF/WVVqq8I9XUTTgVwBLCZza9E84q
0YIvhSnc5oOIDqsWv6+BzGntVcbe+z3TJw3vsO2JoIbvSNeVhMN/f2Qke6sPG6jd5ROSBobR/r8o
CH4hL04Oe2sFqOzFfAOaevq35PiHP8VyFb6qKd3OhICZ61kT5WI0I68TT3G8XLpV3DWGQUC7teYq
kNNbOcIFGCKxM/2NId7RMHhi5mlqZ1NOMD8Iv367J72fzynHAv0gGzpd3iu8n8BAH/ZwQZWOkumv
j1u2ardV+hM0gJD8M+9BtAMk9OFbliNgyi1pClp9X5oCgcAp2BscEqTZ+Bi0gQO3GPE1G63vW8jo
ihwHLShfg9clYBioRJn9DetwW/nTI792cfK2IWSBElw0hfGjurdiN0LmoYaw0RZ338gK8aV6nA1h
O7/mycROB61LVEHsXynAXoi8yptoOV6S+FfRma1vea4u6TfXjPpA05m+1i3GF2bNP/yTNAW1fEoA
S215RncEu6W2oLBZ2Y1dAYX/wYolJ2J5DALwuaPBn+eO0MJslkv9UFMDLbJiWahyCpBeVnbNFxXw
ua4SX4aGMCKyjepDWNyrPRWDAaguNk9EU+0AzbZAoAr4+veo3zEbPJ4U/wx6mYfaQmDGiQ2jffK4
aT8yNXpHrKl8RDHUegcfsdQ6ZKvCVVPavTzLijTFFUtHt6IaCPXlPGWojWseQ1FwmIZqMS/UI7P0
fkE1kFjuZKv3D3ZMacc00Qf+FZcq5q7coYEhvulr1UwB25KmAB1/KO+bUUpmfDTcN+Y0yxgbBrZg
GrIIktROacuI+/qLaR2ni1dcc/9ilYZEVSbDU3Zk5mcbm2myQ41555K9+lVo4oAD4RpDGwoYDQ12
2iwAf367vNL1eRTG//OyZCT6LKNtfzXWs6/UbtCLwKvWePg8g5/PjIvcUvgdGN4HmfFMo6UuJQ7T
T5o3EbecutocSu8zuTZ2aWWebXvm+eqG8sbk7NpuTxacxYeIeZdKU4R8l1veraxNMnKE6UA7xm0L
Mw4qibBU/Rcv0ML57kfDKMMeTJBg473Ck+UFHbNn8+dlmQWa/viJ206OpwyspDfRr0JecU9lrgFR
GGkWBlNAnmzy4y3v+8maKmHcy2beEiT+GfJU9IStn5P+2AXrvsVma2fTo9LebCYKytiHFH10N2S6
SokIoEBeF3Fu/7I7jgNJNNyYOEk6n+dnvRo9O1UEeCGnq5db/IIAb6xJB6vrVxgEmDCSB6XDL7VK
1eCS5VJc9GkuVguT3sdJi3wp3DTS0WSV6K9XeazWdNqLHS3y/ExkZk6bz0bzVzp27Tp7xAbzYG9Y
H37l+U/qRlc9pVSnx6LwF/NnHnwS3bDdWWDNbfCKfBHA1clALWv4GgtaATIly5eQ46+DRlXNnG2w
Hm9Ri2Tkz7VXBRnlb1EU3lEm5zvbes/PFrkx7NiaykyUPMBm+xEsyYkC/l473HXOH5XUbXiATpiZ
7p2FCnGA9FDsL+iAEirCDZkrSM559MOg+Tr3Q8BcknvpjKZ2H3gt9RVIc9i7T5UEGmxlBtGVRqtA
Ji0GsZqtJ17UWExpLtAyhjksanG7/uzkgy33gIKQzVfwwNlE2S9WkZGBk25jGvvzg9mVtv2xQGtb
nqjgaX7ttiRHwCAi3eh8sAtQlBJEarxZ1rXur7IEG5Q8N9GpS74OWOx+Muj4tFdOXQSMc45xPGCI
0LOJwhpNLiLtYqj3p3SCZMCt3lmiqeplrL0tygomktWKGNk70EztdUtVUNNFg8ybg34gXtYpQzNz
TKBQQHe5rmBkIXe0mSmK+d+gc6AbcGhpKsSBmoGlLBYccS6wS59eu/wv78InZlCOvmiK082ZXXDE
N5+PgFUxo1czub184QR9Czfj17rsxh6HT0gmA9uPd13tpQQ6xLW9vVw0S8Nkc4Ye3Lf1PqKs3FOW
nyQmDSd2Zxs/yd138l8lVMw+cDy2csw+mSrfa4qXNJqKdFNU31VTrlnXRrBbJQtHAez3nUacsm2g
4IerI2aetaryOqPrS7syWHSEzinhscYSwtqQ8vH9m1sFkSi6Ug7I12S1P9dSDxrPFkzpNF9dhr1M
zPoF76CNTK7U3SLfH+zc0luPllIhjA91EY5IIGzYc6uBfbQjfGJ8HjG+hqvsQg9xLhbgOWri9pik
Uf3w/1pAY2XhIJGW8ZK18I7AGbuz2HMMQau3p7WmciP0klHILSRXEG4gJB17ZgDWjevG/5EspvUU
SPNagjzD/RpjCvRqgMpHGatoCXgkwMy65xTFbL2Faw2aoLPYeOpgdYOtmJuLkUcWYh78hd2hmrw2
HDo6WqchDUFzW7tPfhRHwfjZyCEjFiKNkl+IwsJKfMVYuo4EfAeqembLvJ/Qpx/0qI3gUxI/43O8
fU7s6Xo5+F7w32DRvSsoqhFdmlqeQFo+fTrPdH2M0KuUal+/Trh5pP7M4d9ogthSs0FJE+dgmC9l
o/YSU8mAE59CIXJ/Uo98eEojMBmkpd5OvkWf+o92iHE6urEziCyelDGyinJ7pEC/aakRfJgymNOY
7PTBwNe9dZ0o582ipwfi6dBkUpGwRIf3Nf9ijz6AuOS1gpmmFIASERdnyzWAosbL041+KsndOJDq
gZ7EM6Hfm70ht0LuhisccPdCfBHGiLNYJ/OS/qrO20w/xb7oQp+1Ld0qQp8P0vS5jusu5uVLDCtq
2ueR9gBFjbm6+yc6h9c3IlmE93oha2t+As6BwV4cMIuuHT9to/Yz+Gq0YIUpE/lJo4n35wy8bdxC
13d0elynukNOHUZ48BdF9nD/dtdob6tPMI3bDIFNzNPaDnRYa6WedMYa4p7rq4yjI7UYDi6hMC1R
L7g/f0wAZo0+hQN/iYAC8YfTXXam96uN4nfVAIYC97fKtV2fBgSV7vYX/e7v7WZ/WnoFv/fJUkP6
77KTd1luS8Oh5oLGCvJGEAQnYJ0ild8jRc3WN8CytI6Ws3DJ82gQABRsn7vJVxgmS2Kybmsp7KVx
QNRoB6qG62F3yWZLl4SwJRAqweS1ZwO6YwzD8LiGtLdiJmUTB15Q1eoDIHvDCJoyJCwTnByofQRC
iiO391FlnfVB7GOVOvrAUXkA33lhcz1gDXpa8e1w/+ZdVbPH3O5smyWlE2J1uaf+pcBwrm5hBYXb
7Wcy4BTjdkMVDWy0M2MZhmVHofuONzRghG1erUFAkIafusGlwRN7fK0gVAZqVl/8N6qpqaLYyyOz
8KDQxRTaocMzW4SsH7BHtB4OT/RbHxnmRoirEaeVW90/vY3H5rynsppobunqSR0ACXHYLoMCoCvF
CwAJEN/AjD3851uGtmfXFWZZmXvGMqTQjSiL+FXHBJMcR4fY4fj4cMUVAdcxN4OwXFr/LNuw32EH
NjUks2ycG4uxfI695TnMS7nqxWnG/mv8vPzLYk1XeqOgsoCeWyU6XP7ewEs1V5/b+blgEEBogkGR
AdMd5lVbMQY5DcSg/i7atthgvByep+sEkwwnRkIfi2FOKfLboX94J+FIxY925f/MV8B4pGDbTb21
1yhhsjGexBZhs9UPPIAcg8NT9OtgMx3V9hZ5FLzaVLfgYdIwPaWE3zSOIdw4DOCs0GPhtsXuvWmb
sSx/vguDrYtFXKPGIzK9oLZU7JGvYLp5DvZnRCRnL3GydSVxVsHGq1V0PbRhQCKT52F0MZeuNKbs
+rDkr4zR6YBDRfQE+W7Y4cmDnhMG6tKqD9hiywgs7AZDrb58cuI4Jwr9lb9NI5P1zjKzcdFonEYp
pFz5zsFgIulT+3zJPvft7aOUppIXr0BhQq/qPwx9dGqj5BxEYtQ0I5qF5/t57eF3TveQWijLhLAB
KTEHgRS9GG1S/xqvZZA2jZMeqB/au1yRc1QfvcqiR3joipI8KTIt1664E+K2ZTzVOZ747D+6xuLm
yR3mM4JL7CoJ1Iumw+sWmny5Rw1Q/SHncQYHE2BJnwjXPhL8Rl5TfKG1bBe7OLeubkm9IBEU9xsU
DhTJ6cBH/f+wd65jAVTZqkbjPsNNcLZcGE25iw0KOn3dZ9UA5Th7YJU1CifnDm85+y3YM1rPzH7p
THfbkBQkrg0gCrujtRjmRlxQ1YshvlaWtuIUUWzV0gZg7sKiU/FugTRxexxUaNITNlGF3wpS9SEC
dKGXAKzBtsUNKrajWk8GPTjXzR1A7TdRYlkli6bN0NNq1bcmA/q9Mp2UJBWqrKWqr5MFSXBPAuTz
QhnY2c+Tio/L+ExqHQavrgIOIX+wwWCX10jvo1la1jHA4ZFlKe5UCkDZ5tjjLm3sBGm6Kyh+ZJ/M
5ZHJiFxbT3HpTt3QuXXM00yvIOdsjKSiFJf/qT2AmFlK/e24uOodmchcQV54Wo1EqO7uh22V9edg
tFnlhqQ7/7oA5e4ZFqMxKWJGakb0BXSOZqCsWGEn8/W6wl4OPOp7G4YhkcPmj/BvEWoS5pTSYZ90
d9g6dCoVYoAoVHC/CcvbAIfOJuaTDNJaYhTnYpOsHJjoZKcajZMNH3yP2868ZVYtWu9/oTWd+Bd5
NuegQpEOG4ht5eiAtQpjqfrz3HbZI1/6TmMkcsHEAhUWUnF7x7xs52aT4qQzQSwPeI8d9qj4Iqee
O4UzCZy79PvdBxDG4U8BLskx4J4ngRiX3n+EfH62bnfLAAIplyMM02KahASudDvkvmlhUT74xKqn
57ykFQB95P4vpzzbR/7AGEFuVP9EmhR2P7vGzONWkuV1LBsa3VZTR4caOHJM15JDUZhkS9SJr0lA
rQQKohd/81QsP/dLh6FIUvKEI/09sQLe0n0B7ZmSsRTwpf52IZxsgcc0pbqF1HsOlUh0DffbU5Pg
PE4XRRKbq5+aRy9y3Pq0gBSRSd7cbyItuUtFgKOjgZUJp4FKm9Fz9VSVPU/bZqJ48kqTg2K6TYZv
/d/dBA78l/QQQvYRL3OsgojkGXIASbGjpO4rjCUUDoi4OHBaQmmNYMQv8CnqB2Q3pPtm5i0Ptso+
T8Lpn8daZYiUuGqpMC5Y5IRKPOJ2bZVbo99OOSqYbo/voHTJs3emCA1nwme2OLH3LJSHzC47ZZmI
l7XKCDh9GcJFqygQxNXOin51LvwTbfYVra/Ne9QyudMI9fuiJnRoQP9QQkPz9Y7eWAFyWnngqn84
DRpVA67Y9i6Hm8rzhQsRPpxefTn0RwOHPqM4nVvN8YmbHqQD34nA8nq9jcWdsgFfUXVVjnqlXTdt
HWmXQ2MAF3i4xNgcbZUAyR7DY5LT5u1nMdTAs+pPyNeD2Vjpp/84j516Hok9ZfhkXy2VMnU3ZLlY
11F0/x0lwko3UAv5bS+rGnBpb01ui/x1hON0wRlGUwtYWDQ2YlWzRakIqWeyvWnVoycz6xfzOTbM
KXoHVTuuo+2rp5SHo6p9CSoeegCbnsWnCm8xnO6lRsoMnJGDbwaJPTTpd2n8Rz5cupONFJH7ZkYL
hswYrZt+tjoylB6ymGvQbrgUpeGvmafvDRFo7cSUt69+s/17D+JKWLHC4Pma3fgoPIOnTtzmpuwI
mh9kJu0/OAShho9fMgxcGa7m2EfRvqPEhGALBAWZIMrr6YrebUJZwOUB2wCyJC7KfRaZ5WwUiuDO
e3YENDjMgtwSttkM7HCsoED6TeAYJjFxRZ7SYY7nVN8yoe3VMoHqMmxZ2EN4JuJrGTQRvm/HGX6v
RveAzPpVyBj0CCBTNzUow9nbL3ub0JaKT7sdcwsFPEZIZd17IeJoORErZYWIYHnO8k0+W+2zCc1T
tKKqZ86/yeSMUjXfGlhndfkzjTFA+65jmqp1lKbLmFbjOM66ak+oo04ZtCnihI1XqzqsAppE1sw2
fIY/bWAgV/8mchzonfLWMZTmwAfl0f+kCLjTUWh8RQnuaDBf4qouqC3jbxKhY4gzN3cQq6+k3RWZ
O1/EjGdiPuSi3LtMDqVethrxBJY39NdIKfIV5lauddHW/RSZGU6ZeFfSdEIGx+iI7nkDxgHDApJA
JnL5lqlECK08LE9gVHefTts7hssXVX2HVyT7IyU2xcKCrtnNyqRnrdWnDih+J2UrpklDXFuj9FUC
FRaVewtG/vYAchM37ZXKAqtPbfMUVRbUrYXxOBnOlm+WZHBCbXtqDw6v/OnE5P/9gQybLpIs5qrt
obVTghBDb0XGq7B5wAgLtcSZWT0bkAw2ADFshPSNetzIO+t1nubRE5kSHCpgPEWJqT04qaAkxzsV
shZOThAs+phf0jJj8HK2mhZcpar4p4+XXxnpwb+rEpA9Blsru0QdODXBxRlofwFU8tKa+N95WPd1
f1h68v2orh603F8s+azZtIOkQSO+1V8OdGrLaX/QOsGEXOhOWuarOyYu77+yRo5h+oeH2XcJwV45
3LzT9jVWK6vdxIu9Eh98eMOJNO6iJpg3NUHlnKw9zLZXTaJUatu3grGiAZ2stIjofLfm3Z4DyZvc
8MR41U+qHib2nD6CTfarDoum64871wbsocygZ3zurkbvAnVEpFkg4hlZGBKT2z23X3gLnjqqqT63
GTIZ0gx0XoZj8TP7oyOcLFE4Q+3pLTlnh+tOCmKXQuWp1lzOOQTvM0aju+NnhsHU9eh2DGvIfIvG
EMAd03yz6c6ELAlgz5VJIr8lvugos8b91Yt7xyS7dpfZ6C9+cehEHCCzgJdYgvcpqrQCqTh8Q9jp
rXphLOJ0gTm+JyiFUxH8vUMdquNQHATy514izzR5DUH0QapPyzZiSUEgGU9R7it7zF/LGQrBcPIa
dyNkrTQaMWKzZSeeyPCatifOeEcCSQBO2BHVsyxo2PT31V7VB/R8PziTpnJgR3HLp/etMOE8J/1y
lwglup2iskBJxSLRVGqqkMs5vUenmpYJaXRC3QmVfqmLXRkhogIZ9tEsRGp9EV/qAsO3GDyy10yI
fx1lQhl9+hKw8vafhuy1+apgVbdo+DYR23EPuiKw/YA40qS4NJ2QUxU2mVjQn6xJEqjxTyTuQC7W
YQ9avR51oZq4RgIfb1NpcuG91oxUerr5iTyUe6wq0QKsDWL+L2BT45DIR/n6iclb1dFrKySYi8Ro
GacxDUO2TQsZ1Yhj6OuJqwFFQCUUGB9ENiAOfzljM2WC40o1K/Sq/Bgivkj7POIC01ILcMbdCK8c
9d8c14Dxf+/SGEESG10GidBypQvaVm8kYm5k/gvihXSLH+2ctKj9CEopa88ATjnwmVmLDWLCCOfS
CGoB/ylVTEO8qLroulV3L9EwoesKTs1R7csKgHEWUahaHtX5O7PHk6Gleamo6Raf1q+ndveRgQ/o
kNNMCJj28u2IFaUBh/QzfxWN+Dawcp1mFfCaEGTDmOsq77SgPcc8JonGPUIYHuvvDJQYnnPAE8DK
SG5GbALE7o1UUPfQip4RRrOwsO+8s4UU091Us42v0gqoGnbpYzAX9J115uMCiHdI1ydvvwGLgfuV
Wp4ACvzVaemdkPtVALPoH5J5mWavRBhCKqTYlKMGanMWqFhjrWzGlPq/aOvFt+7VXdeXeUqlMxrr
PavHP0xbWYm+xj+5TnNs72W93+iMbb7qrTBU56z1NUmOb/hnDN1mVGnakYB5NH5XPZRUhAFtk4tz
QCC0UBF5wV0V0jyVPOdscs7AECP8lIzaElobOGtFeAvDtM+7XzPfcqKeB6g9EJsm+vAPDNeEn+fs
9WkB48ryG6r1GVBhJjU5iwr/BohWWKSNuTAk8C106SlzJJk/IOZIsSo0DH13QxyTu9Xp1uIgribQ
Jbck5ChZ/GJ3ag/5vaYGO5ptk12jQbzd9r5lcLi1IGIQeXPVHtj5R0f6WjKz3TJoJPXvJ/XJRLdb
dYJ8x8O/c4xVFb09Vk7CuXm/Q3/gS9GZGyO0Xk3YMb/59mVApp1aq8Wpq92q88A4QNY4Erx0GTIQ
CARtWyUraZTQ91IVrOMtark3Bh/c3hqzuk/aYsx5N3fY+mMfYFkRDaHhp3xn6o+5DtwHPhZ3PQ60
ID3K0nkqVuif9sILCeTOJ0IKcZtSQa3dRrTZB5s+5JqkPne0atAA/pOMCL7CzYqWS1UxwA0R6sZh
w8rgiFn7zzfAQZkDKZt4ngDuTwAUnpValAs4GDGvgA8GGJ+yl6Con0mdD4yXCbd25v7cRM+IWzhe
Jz8Er8rL4mPUWsbuB3tL/OFyukNhlqiAPxS+cXZ4owGteq6TmYmdkSZkqbkeVu1VCR6rPeS/HRAY
CcW3kJqlMUFaWMtn+WYF71WwCBzMqpgh32vBxZ2jQkwzh8UAFEy8YnLZlE7p53P0Nyf6EEZionzK
E2sv8L4TKu4vD0tr5AB3E/R+1dIEl9cih9R01YQ7fG9hn3IpLhrT4An4KrPaYFqGWbZcsq+5k6MY
9qgiam5pA3nK3a1tot4J5l+O+i9WNUiNKNtx1XUD7udOymaRtqtSlv4GzH5je0dz29qDq+aW6AtX
SapGdEGuKUvAN9WEN23Bztjdt5UHSB3e6DZu+5womy3l3YZ2a8IOir5TpxUYW9zxuogS54w91xcZ
uX2yOcDzRrCT0yGITKmewUF/RGq2hjBlDm92MkmpesPyeTrKdcrZ2lvabNJzyljyHia8eNkS/OH1
CBNSJDsOcsyvRu8rByHVcV2IOU3qJ8+R+e6FJ5ywQK5fYnkd6Cor73KpwWN+lp588s8ZcCmir5NV
1htQ3cgxG3vnv7gRNNx5B5iycWcf+KpUqTdNJqamerXUlsChrTqd+gQWoiWdYpL36hxw1gEu7ZR4
uu4nr1ftAnaxezhKZWgzMvkfPax3dXDhcuYUmnyffTJnMnjXRp87JLv9030QPTR5pHYT5qa19kg9
uziu20/45PTSutM9q7ZK99g2sWHAHH8m50q3/ODRX3iy8pQul87sUFgW9211YI/kltDJw06o2jXk
hXKzxOG53Cqx1i5WgfDwYxVFeMtN7wRpg/lX8IgyJWWCAcIOsAhG2MrGScdV6uQOPAtjk4zv42Sz
KU4hGGpzL6rsZM0D5jzyyRMcMPx57mqXkqrOJ7BwBzH7aeciZO26dBAs+J3H6XOBAijepk5IXDAc
jDIleYWhBx3aX4yb8rLvI/eFgI2Vi7wfvHeiY/swGZAypRTdRNdDNSZOewOd+VxC4JQd0qf0rK9v
wYwuwSYvFe+UavcUTBoVYhuugd1MbiiR1AEacws3T0q5gRNHs581l5winvwM/7yZcbrRb7/iO6CC
EGDWqIDfwUhyLOoPQRBxndKR6W/pY2H5zBU7kkUxObXpPleJtN5KEZPmgEdov7Zqa5egPhyxYxf4
B0Uv/26ivjxWMYhcSiI9q9/XqeuDOuPQddCGcAUyAPd0UX3jUjM66oKVQBe0iu5Pxy6Sxbw8CTh1
r6Fe5EL//nLkNs3XYLW+KHKDS3Evhj8G/Hk11AY6V0IznNpiO5lWZv+lZKzF283pGvrMmVMUDa68
34wWxLsD1fhDhC4AZA9l2uq6Ee0TU0AO9ruhexMJxnGJDNXjwyjHQur/a99F2P7sK2Zh4MkZrS5q
G1VoZEKr3pZIU5xLHc/QlweOQr6eK07PDQa0g/zvwRdc1CSBttxAwP/lpDqofyH4Vhg9H4DW9ys8
3VicojmY8ZNPPhH+pTb423v8K+GCGFKeu6hDLEf6DEBUfsEURL1odr0ZCWPSxXIFUWa8CXLjTeMB
DvAQcWRNa8Xk4VHfOdpo5dEWR35xyXHqohk6tUHkesYMyOG/IH2A3aOsfd7z5ktDzktVQWQQuleN
ys7IyIqA33h49YX2jbuHjzpQob4PS99dfUOkW9KJLaveAwCWUcOV+F0qsuH73ZU0spjXzeDO3/Sq
FI21kpC9OYwRH05bO/51/eptQu/4ewXet4I//su4d8el2vl9g0HQQ+Nk/pjG/lQtRt+CXsUX4Von
n2AS7iQmjYnGUt1TgofDVaBASFuLRjyzzfZzzWeMbHAgLn5NI66jXpga9pV4XAI50qh6dlTDsRpp
bjfi11ci9IJX0Rp2Z18RYE49JTeRItheoz9SKFdd+xURxtTiQhGroXU6VlgBbnQ57IxCsAf05NW1
66EV9XkCQn2DHI2tOcHmbRTQp5tXGXLEzX6OFyI6mb1uYldm1VMw0hpWH2Niov3915yaarRtVSIC
GUZ+2Kvp4NDtL3Gez/Cj/ZGlW0Drh45BWYw/r0a8lCwTEMnMzC+02pUGFPj6zNEva2zK1WwiDyVx
ABW14eIJUBhhBPsmu+gUK0viipWROf1b7qfuVhSEvTC/247v06F/hYayAT2+u0eWICti+QWWOEC5
4VIlbXcWqR7mnZcH1iqkFJyxEViQi3PjfAVhZojrcR2EQTSspQQ3o6TtAPGW9srMUiLK/2Df0r+u
bl6ntguJMImIUc0PuiDaiLE2f1UY3+9DVgjkXsOBj+Zq/xU1RykMvjuwhQRFHOxhl9O7M/pTeKha
ccZgTqPRcZYa5uPp//J1UMitPDw4CkxCdD/eYYdaI6Vre4bGa3q28lan1MAiP2QpGyYoc3j1FQvO
WVvKsipymD4uBumpDvpS7L5BpEq8gTC4ML1mc2ZzclAdt3D8SsNFRI9gRZWGWdXcJaPF6IsA4ISf
L8pjM6//f/+Ix9v2r2ejgUp0YupWQtniJXVFGL0N/NE19auqJVDEm9qZPvqB/Aaj1yghPHS28kLL
06ZzA87Tqppl24U8L/obHPIkklLi+TnGuwj9GA2N/2KMJixdLdG1ziQB1ZjdTAFCo9SsNFkjpst6
wXfUPRyZIs4gTmQFZ4z41bdnoeDoPFbUWHbUJw/3NAQyvhuyy8ADS4+zTUlcN2hMRbrOUbmCI5rB
MdOOd9plUZuLWdIScrRpXwXLtZseiHsdQ/a/yAgxcjq6mACorscveUh2eID6U7/9APm41WV267n8
8ryWGbDybS6pN6pQNa5kCMFBmozSe9QCT0Ngnr6NjNgOc4i+ic1BAPklQQu+URzoLnQL81BoPe9h
8ytR+IAPp/n9UQGjndS/1Z/K4G0UjIzykCBTZdfz2aSUFa5fZsB4x5xeGPIWbhxAnrToSQ8BbuaM
PRDLH1Mc7PlFIWvRJCMdITREdpCFo00z+tkcetqvDWdqmEZwa1bQg2Qt5AUm6s0g71FrBnnS7d4f
FzLMrZhqMMwq3WbH3oh4kogGluPKaMoZK3Z64szKeC2WY+F+aieTc3HTwYL4fskb3OCd6KiPigDE
eukA6PMQGXxwWyYAj10MMFPd2Gm2t2TbtX4PCHaJhOOTq9f1o7dx+VYoPl9+A12XYl2IyVZaU9Hz
a0vDwvGnH825cGbzE1wcb5XJzBPKknFoonC6O5HWu5Q7cEC+4cBcEHJLHLc3lwzqmEATlCfYIFgQ
54y461zcpfmeleJ+whiJBgB0rwoPVPsRV/lQG57Oehi36qq5OrakrSXNPoeXr0zIzQ4RsTmhKp6Z
T372m7HfLzGEsoL7eEcmqF80EZC8/5Xt66MGmln/+D3AVAOOswx/dEuJbzT9kzbWdphHOfQod8BA
Vc2Msc26ugY/8gSVCGe3jyLsUHGT9lD4u8Cx16+Mka6z1qQ1kDLblXrZmp1Ab78F8aNn1p7/g01U
kJ4s11GscC9OjfVv/gX7H5gI6yqCGpuXyq0Sk5G8PaznwD3gFECObWaMwBkKDH3UhjBOfBTAmE5z
OLjdevRKFu/5vBRMG/bZqfDWbnSILXGU26xjxwNTC+9zKv/IWoxDFNZCTiiwia7pmiMRNQWC9n6C
RMfCUGsG+1sFemMFbu+OZoDgAw7jCZmASiRVDZ7V6irGbqODPqSQU1F/phqcTSO0/2X959VC32nC
3yb/MECyD+Vsj7jAxygW/xdW3Fvy7H7BazK5Nbb3JNQQhaIIyT+92enrXmnJAN7XCxjEl871qRbQ
N3uNdtIY+DB2B61HEb0DjmSpqJaCHhlVGY31eVP7oUd04nqtGwHnuYOpzqBLe+EVDUEYYoafa5Ve
sTXnQCAYl3X1KuFy3CNWKJCnpIxNfcs5QeWTIoJUOmE9AaZwOj+CRjMMT1/UWDE+couyd7Qpmlrm
KePQwKkp9ZaPYlrHQ6vSrOC1JMMI2fi+3d+rH3iGsrvilGEVdTwwK+mP9xYjSpbC9VNNNzTyrrMK
VJfGI2oAHS/Ua2KO5RrJTX01+fJsueAMXl6WEc7+XXnXY2VlT6FfrcaOL4nUxj2ZIZqHfww76yaN
NqvzHivY5UnOzMNdDmPGgEcoz7fQ25F9mYaoDb0uk0LkZxR/94HEA3DOcpJNZxTkybRtaBXXyRGx
2fANYC8e7Wg62/UtQvAwu6JvPeSID+hIWMlHc6gLrV/3tKoNqmjvhPRvqEvhJXJA/pFyzZndMh0N
eia4C66y9SgvNc2NN8hKT6F3jPE7OVziLRrvecfi7j1v40e/4LJ/nyMBgkZ4tthE57OwN/0YU8/1
UKVSQhqmQ+HXw8xHJkaxGFIkYya3XpW7U2OQeAyeizmLgrIf0nZiijbij4HuLwsz/IH8BDkqYusu
gDG4THaRa7kzlGukHTuqClIluXTdJgQ6sR7JeGlUFD1T1VwGpCYZVWsgOWM9S5KkRldeX5ozG6xR
/ofor1RHcJbTkLoefOJ6+guGWw3W/H0Zt8g8O37CPRG0Ugng1SjzAXWasEQMEMSIdJRRbQm8Wle6
PcDqEsMxPWJ19pyCtE2ppgmIygtdLmLcvUjVdNPKE3Ues4+b0z9JOmimo6zRe61anUeORbfz7fSx
o3wJ186Zy1PzMnwCAl89dDk9jX+iIIaauPQeafrFmILKX6Ar9ZifR+sUX73OIbl+9T/WqjMfJYsB
UJpF5GfWfaMTVEJtUpap9DQSQWYTvTp2VqsYMq+GWPJKPHKlaUov49JAJk0j75rgB7E1JeTMsimS
Uy+TXRTlHslJqxK6oUN5Ij1lvLGUq2uIkOXRBkZk8mtnqE/ysv50C/TUkoLwlKhN71qAbwbaCqnP
HIcdOPY3OQeGJIlORGZcytV+XcCJermfoEm6FcvlKL2qsPE4Xvc2UlVJiWxzU7a8xMfcNX7irk78
lHKT0cEJuy1LRDXbldSMfg++b+7m6lO9S++jo1/TyzGpZRKiBzOYkwUydRP+AaDVQJl6Oj1E1969
SoDLRUT9vGYCO15iUAPs0XcCsYjpM43e0DIjvw7NUGlFeFJmB/uzhUQKFz25LoF5Xp6suxqfGBJk
tej40WprsKgsf4iI6PPL3/P27sh7Bi8KzfjZK7fUOxvuvC82jCDfpuOkwokfDLDRM4yxeD8fnely
1GRU7OfTnqa8GKyo3P3Hk2qd1TLnBRloqHjzXvh3o0Ln8Y4e0Ai3VqzdcTFCqcNJaQ9NFgSlCX1a
46oTGnSAoMeQCugu5BJqu55u1ptxaTo76/iC01Nz2VuLbuXxahJUwrnSoVvejRi2M7Uh63GYyRVn
oTViJzTRgI8aGcLyXZQgDVwgPWrxMCFa8NALmuCZ8xxXkkKKwXEfNaqRabl9cys0AYFrBGO77yVq
Ur7YUU6V1jdDu59egQOcDp46sIOuzMfP9At20wTiUZDp2+CWGn843GfT4MMNYxiYy93c4WjzXwSb
kYuZszmkXQDgVGNnIT6B9oAeYhpSmAX5XO2+Y58RAHrsoICS69xNSnNQOrCJcSDk4sHmLINEvYB9
Wmz/PpsEyl6k92ky0Mi8IWqgc1rBI7qz1GnhYXatjW3lFdQyj2O0eMPEuV1p25KmGl8gwsnikQXL
k+IzFMuE/xk4BmXFunQPmYo/NmjqYZRHmDLwEM4yvQ1LLuQDA6a7RFqy9uJWB1JuruCdD7cQOkpl
Zz9wWO1d0dIN558hC1FhZ3wUThplYg0PYWbF2sJgntLJX0gK5gCRTB1KqKhtlk7n7I3uQW5MEeDc
3w35AyH3ymwgxytSYw/MrVWOfHmU9tOLrRAr+Dg5Dytgxp2jzvAsaQ/DaX6PD7nlGDSeDAxs5v8m
19XFY08SaAob/iS2yF5A937O1oSLnypLJSi6rImaFngSmAGZkigcItj2V7ZSVh1tul412sBeMPj9
jsXC1Oi4NNUeZg79J/bsZVNjNi5ClpSPYiFtPvbLwbqZEYT15acP7gkDC9gi/jMHRgj4A8WpVysn
FNO53pUB5yEMNn13ytWLm8AbkXCViOnueUgKtXidQ1356BeMQrmNNGbOXTtNK07tmeOtwYEVpPgp
boVqFv9LJVfkuXa9L6F0PIN1L7yDbFgPDG2kfbye9T0CYF0QDOVJ+YUc6wKwgjtbB7dy2gFxTvBO
s0jWYpPaF00vWUWFU44n4j0xWcQRJOdFk5rpY0sMM2l9jMNH+skQDXPy+cZ24tVUpCw5lVbVPKlx
Aa9WB7mpllTUg+SIOQkg/Q+hViYPIf6NSAeJq+FRi35eGWTvlULVgVnW1o7oCBhTstjYNMjx/ddn
c9znaC1nSGELr901imu5l76M60Elp6xxYB0q0UYKpRaQS3VFbSRs7OYnmywNtAPomqgRwvEJdlOy
LxLWZUMNPuGperLuWf0hZdDsqzubwEdWemNWnaVx7sUmdmZOlqJRyp4iaVi8i4uGJZodvP+xdbGj
zjQijQVLg1vJrmBY7gsCECZxADkA9dE01Ij03yregJJe2RA1/dadXUzfTaqN3F2RTiIfe2y9UP1h
Eb4sVaMf3HN6zHepxR0P5sFWMA4LSaO7jk9d4W41CDivflGQn4zt91AkA44yAep/lurvnGQd0v0j
RNeOdxfW8YBv9laC8DH1lg7XeL8/F+WWddlls3LNpcaoNdYldi5OMNvc5PUWFxfxa5D2d/HSqJRP
zNOy9kvaUR9e0WX8NlR00aizdpFz49YiXFzksqzeQsa+4uwG0Jyz//0wc9Wd8OoI3cN9hEnjX1Tm
x2UPDnIohGTAJQaA9Bi+B/CF3eqdZZFlYNWr0ltqfVQy7GHA6tRJu/Lud+BYe7MsL2FbrTFwvQ6t
+ObJWEhEppTFb7MgZbuKhIa345kPlw62QnMw/ODMJd+bw+v2VSSVLjzw7GIh5s6DlpuzOHtpYFfI
vLNuOuplLHXcUUCVWokUXnodfkyLJGoL1BCouPjfJHV14/RNFp16iWu7gtkljHWPLmb4bwCz2jIQ
l5mte8jGcX+h6bCRQ0r9mC6Q4bfP1j7uRL703Ni42p6LYVOg8cokoxX1t2SuyvHL7yHwqQxPV2RZ
eToOcMEBsjYcpwFsyTp/YhJKxWJfV2CCQYtzMKWTa7SUdGcauc9FoE6JY2giQAr+PkAxpAJjSfge
K4nMwMSOB4RPXmXXskeJCRvHkPr5zNwovMrOhbqXAztXQGJ675vPPWxAJmnYH3pJ5faUC6sjBjg6
MpCOqTqMNatH0l1B2iZHihbu0HZM0tRxrYTRm1vkb//0MAb0/fuzJHDiUP+JIbUFyYUMp9yKqo7c
unmEs0ImFssXymZteD4DDOzh9bPJrVqlVS+G88awM5L+eN1Lj9zHUhx+vtSh1+Uf37MeTnELP76u
eW/3JeanJWeqKd3CfVSgA4h0D1CdIwOVlX5upOrJN1Hkggz3wKlMpIO1HFb2z1MVnTgXHGIb7rmI
p/lEb+NsYjdJtHQLc3/FYVf2T8SU6CXsHsPy1IG+mlqsh1i+ZMHbs953jszyvycN5oRJ7nNnZkCM
zYyPLqwiu4yvSSMeTmYOstMS7wGTO/g762Jh3JO2vxQoKrdsUu0N9sl/mKGxrGacKIDll0rEvJ39
Mb2JrhmDNEXCrqfHYMMfvk7FVtLzv3z7EaAPGuLzBpvZb/wrYiUZy7P+jo267O3tyvKj4pOq7W17
vGcJ8sxYtqS0kQIzu4gcVs2E2bE5KC9xnEedmBYy008NE3O4PDqlhQJTZcjcbx9E51SihTOieCYY
junxdNaA6ob54TyzPgGNGviyJd4yJnikpLIJhxZ11XLdrx8kk7XeEOHsw+TXJdy5wX7D5/ghGN1p
IsG0H2/C0+OVZH+ZA0HPDSxu4kCTUcZLRlnVr6ROVe/f756dXAHbpLfOcPG2SoPrAy9jtOnt9To9
ps+oO89T7P11qp5gDxLjKGj45oL2ZKwahd4nwDu+N9eVak7qyg6XOBELrU4P/ABlmIhoVnvmXTUG
r4UeGO1s9l4tRsYAT0WPdy8Z6iQQRNdTLnQB3WUEalRw6aiwcHCzUZfz4ZwP0/zDKNJXwEzg09Us
kjiBb6wnAAJbju0Ao/Xi3ZzLTFUKhLPLjq5p+OjxsRtgrDhsCBIdtZv3XENeNB/s67+Sx7Tnf34y
f/PJiIulgN7ETQPpB1Quaxjp22K7okkuJcTMrSmIseurLwYREvpSG4bXysm6OBzrQu4Vtwb2SdXE
mmKY+RoEiLer/y5xXT4zX5PrauTE+2FbRUfs4NJeoaWzykjsRl/nggQVRqjmiAwsQgxuJSTehuhF
z+ZtF3mhfNKoJkfkFsxBmCx9kVDjEFpo9uLDmwxkci+RsDMXY0RxpT+X8h19AUymtiu8Y7xzl15r
W5bj0vq5UKKViSk83GV0MfI+f0HElgiQbz/bLwmvrG6A3u4pnhLr2nBlLN3nR/x/+x6zWrlJCH3W
9Y+Fiy1CGNRA6OxOAP77MfhSdvIriNl3ufXeK8D0s4Tw/Kg86gTYJ7+fC/DK/+zriyzOUCoBlFyE
KlYAsxRhQYcXsHgKyKvEpeGZ/iuq3LCipO6PAyazQBInj1aGB8VIBsRMb4qTo0OonhVK3dmw/WAV
zg/NDPkiG8hPbdQSlIHgrb4prh4rpMChqjpddNJRh6+q2mfniapAFFlKVKgEnTheVFvb+zxKhkEv
ER2OCHwPYa3elN6ggS9U/0yQfeZAR85Jrod42UG/JEVM1Hqn+TP+ml0t8oT9SGVh5iknL0SfpNQx
h38v/iTWAQTBapfUIRe4Z3nO9IHgKCsoDrlAxLLIk2b0dFWLfALYfrWTjWp3/OsJgt0emcCTIRe8
QhpejqjEf5JwMkUD2ptenoL2ssKeW6cmwsvsk2mcBX2g+XV3e2eidAFea8Bbqbonl41aTZDS9kq0
iJRjTxabRuHyDDLvX3wpK3UbWwQKe0ETFzrb/QOVTf+8bbsMyDSYO3yedI2fEb9a+JrDBNKjvPLO
7ZZ7cJxkVre8PCqIGkw2XSGdBKq+V9MGK8PnfgC8h7pzYoIeOrHB4PLFuJoKUCVWIuOjAtAgWqmX
CGlsV2QCy1SMiLLkCMElNEdSNzbanhO3RMwzv8MNneGr/bNWLE41aIlL/kP50sX4A7p4NPjqxYXf
mSTys3TM1jlz7Cgc9EmzCQ6uo0haCOZP63Q1N12141zPOAuprP+kXEHOwB/o8D0Y3nmSeorPyV4+
O4M36QugxHKUYu5uYZ62FtxkCoIHqxyM+1J9KDsqi7xdmvinmCQqL+3DhoFRUYrJree02hQvkw+n
gi9tbt1pD4XMucREzUSE2bhh5Uotezrs8WdXrfAndbvB5Whx1EXa7PB6G8aXVkgP6qL92krXlaaD
Qo5L73XhZ+r80qErQVACIbsg5YkHKXf3IDrZoxDu05a8C3akBUd4VGR1cYjXdfSrjUrsgih+61JT
301nEV7to2xYXIcm++706fT/3+v/qpL8Ls36bayR2XGVmAzqY4iu1Ya7CCNihmhbzPlSItLCTP8c
LBjOu3K7VMCBSQZN6LhKJSn3q9w/BZgKvPG7/phWn6t4POd//N+F28p2KO54TlqILRe5jCwjVO7c
AUdlWLeuDaM9Q+fahIU2QmuR+RMeR0qkxIjpbJZe2h4R2ZfIqcSG+J7ikx0eSL51Bjl4+0qjzQ4M
ikJG1K0ZRZgiFamixP0uaPk/En+XJDMwiy04ZA8OLgG+vSDKb0f5t8CSomgttO1wX7VrTnjsIZ6c
lfq20ImGNlC+mK6iAhP7A9zerwAw6ZD91VFgx936fZ1cqVN/Etu9zTWYcfcc+mMFCWOGjivsUX+N
O6acAFcuVxq68s9BHFCrS8+0tbRI9Z6LQbAbpu6vcqDDd1UhpRD2iYBvnNgz5TiK6+gqRoNz+/bc
+Go3WCwV4XHtT8FqXbcpbG86jhnEYZrjXlNNlKdIYZ5LPscKUncAjpgZlyreaQ1rvAB6Qoequ416
nWyj1a9iJMVS9y87Apx/hAjP6UnrxcW+QhrLrZ0Y/H1sW8/tdFhg95ayFzLnZSEP/ryFvECC9/2B
AK7m917oka/vWPp6U58pkjVePjg+Je5kWpX7515N2Tyb/Za9yBPtn4iJGlELb/ED3MkkWn16JKus
UPNz8bvPxCJ0TjNBuQOawnkU/TpHPs3fP7NGEgbdwaYo6+VCExxfCCquT81IRbmngtkukMMLS7EC
Q2inzpQtTBk+hzizHV2x3xrBJI8ol8TXHjJpK9dkKBLVHpKypnu9wlLjQZHwyfBhCJpFuO1cONwA
ps3gb3CeTYGUqLkuAfbHm/JkJibXv9TNti5DgXtNB420klvGWqLoyTAPGMilPgoMLkTC1ZCVVCBe
Jz6Gimov8Sf/GhLiQWkwopzK4IMNaqCxMGpn23TgwGnTHQfx9zkhsQi5x1XT22mBo/+zi1zlqfhn
bli1wxa3j32uX8n4Rp/CLugyLzBpe3FYahqfTvo6ZoZfiOGc7XzaMxLyLaZepx7Oi9dwNEYvwaHJ
Sd+9kGW/9kx0lCs++LaH1U3XFLx4R1izLDrwOBghTHEUP8b9alpBRifdW7iDwtM1y/p405hlkUi0
u6jauuEB9aL1QSlZfcI9pw8tX//797gYkqt6/BIWThbRAndmzhDyC47x99QT2boVgsrCTgYIw6eE
8Cl6/jkJyFi3aq/rW5lpCXitisLwAw39KyFCSCWdBfP8YnpHoytiTAfXfD6AajXJjH4tOCcjjGSO
huArHr/hv9OY0r3ERpfd4gxjS1qOwsmhPQZkp6MeoafbNi+TnnVQSLSq/MDWA75zWMVDZOOsf9rg
iQm/2EE4t8QuyDUxzbK+IB378qOcWi+PRCy5EWZCFGF0E2u3w2GYiPBLOCz6m25+D/4K+TIRhhlf
NN+3wuJ2RJicc4fp+ZP2MHHe+vKXAZ3QxfDvib5/SOB9CmV336bG/A+2F+tV3r7Rv4ej6TRV0WX/
ZMziCDFODF3nHPm3hqofJ8xGesLnq6OPAEWO/xRjBi+GwYLkZFfD0S5QfPjYlQNynwO3z0T0ycDk
ssHXLTE1eRyZfNfqdKtLrBiyHHxVlO4SCnkdNL9NQscze2GM/6geLhCAoZz7cTWGePVNbyG0akDa
ZKm8GnvA2cBWeL26RumeN/TVk/JMLaO9gbpY0jt367JPTGjM9x6c3MHUqaIVFrXtexAIS31VSKoy
Ru0PELhd11IYPWnWAKdbsrZePNpzR3JwbKYkJIFk5KST44wyNd7TuzSvPaoeqU7zu4VtJA1bOZOy
FiH6OHV2sLimD3AOe4c276c65T53UorAp9UCzBnGvGv0WjO2cEJaprNVC1akI0hsO9c5sIGzZQ1C
3tZXt35y7lcYrzRPKy7ZZ+gyvtFhQFLolR7R0GCuuhlk5GOAJBt27T0gsQILSIqG78DLQ0pvWyNS
ZfXk8C9uUj6EITcnFb4bSeD5Q7BnDgdZDXUDs0iey5j3hfsDuDSJryvQjnIscAzeiQMuW5rEFMr0
KqRoMJy66zMz/n7QYJGoiJvdmXbmhoezt8SfXhSjCUm0wxX0uF80aLdrN+HfDBB9yrUWrmqMB9y0
7yYawtUovmgOsLreGgNXRnQ2dZMpUWRRODAl0xxB6nBgj95isnLUd0ODvdWha1lsVfHoytVxbJUW
DCjDHPAGt+vgwFYvchHDpyDLQfMLYpW3pEk4lLORNKatYnUJxFuDMJnlcr40bUaC62DpLp5/5sfT
8gVnQtLMfKV6i8ge8gQvlwmhrf5cVtk8SxFCC5BM4rXF3jt+NQXwOsnC2gdTf1SFqeO6zEXVclQk
nun9YaymBYkz7pPg4DmNI+0nJIgXljmYUjEQu6CmjnN7oHaVANcnNBjzIUA0nMoEr/7hka+XdHyQ
I6i+ajsNRUsJ56IL+gOrTuHtZ3Kz18SoEjGyHUNByexo5MUtk5tqkdy7+niiCEDgMEEaHTxoua1Q
6IR002wDtR3MYr1Vm8Nme8uRqYJPmpx8oKFxy/z5D++AhAosq18GJigbzPIv3cVHNVj68OcS/gqr
nyHz7C1OcW53BHS8Y3513iesmGFAohiWZNnOM62jl4mNBTqOU2PmoKhAVf9IL4pdiVwIzl4mjovS
8CimjocuEwrUAEpy5KkEgGBTtY2eGNH+jIYr4a94qKPX+4XBEkJicdc6DvF8+u4VIQrMNudGU7Wn
z3+5BmKM5o85j4qkzHCsM7SQmqpfznCpW50Ur045e38l1oJyqEa0EWfjJO80z78Egfuu3E0Eq8fm
Fkp92kMMyfHnfdTdSfq0TrmNPqm6l+A0Kz4ch68T8xOmf2HA/q96pzlNUoQrmsaDY/G3gL9N/kW4
Eqp4TcpGySK4z5IftywazynpUQosdwLwBVmTbjKDi5iulwTKNea8jwFP6uYMujMNC4fvuzd2PpcH
wIhV6sq1i2m21Ac9Dy3TtebLBQDFjUaHbVOx9D8auvIkDCgsCFzzLrOhMImHCn0tsrVkk4o7BRF7
tyFKgZaFde9spHv/4Q+q8NispEruyy4kYLCN7pZXuv0lvOogxRnPkD3jzneDzp1CKBQbr+RoCLdl
AOlrNjnsd8Ni7d+CHOHNA1tQD5BrBr97L6QHlriEdjmLWDNL5ytybNjH+6Ve1HSBtOQWB1eQO9GU
mJd3pYNyQ1NWyFONjm/g72Hybg1PIe8Rr0maxGM23Y6uTVlxuBX4Q4guv+ttksk/rSCpUWDpRoMv
3KCUDTl1ZB+XiJSiMHQJ4TkBuK9oNA5Qb8o0uT1FmzWVw1xegYSRfGd4fVKDHaxC1fMP6sYw3EaD
o8nJ/IuXApJChN2y2GTl4qvL1sfcSPhSUFGUZRoZ+wtJ4F1F22pqDjP6XglrnEzOZWH+ZPyClQy+
umRS/xFUgz5N8uSPe6T+XtockQuguBfMs1r5In0Xoi+fLT0OdB4UZ7B5P36tIIFPvUM6uBEiX+2Z
ECPtEP2B5/sqNj/oOuIsveO1gkrgFWHEC5SlTJkOO5SSrZFSSMxXz/tFTK5qajPYgKyEMk3kjF86
5AGIFJu2w+HN8uXveJwpPcf/ob4G4MkwuwULDBJr+HWaAUJU0UGve9ifIhOcoIJB6nvqrxWV4rLk
3w+fusTeZdSxRfE2UYsp+LU6Rcjj/J2FEUTZdTQtfQMRtxfrfbI1sLfxEoJFB+1Pm4THpQ3dvaRI
44eEIm5V/gKJSO8IN3W9WyNQiqHmKvz0AcZiDNod+W47pvgVmBSOfj+4JVOri6cZCIcriCfGxloo
hgiWksv77Uv6ID5blum6zCGhrkLUeykmaG1oHlKoir2xryhnBKo3LNWl5Y1e6S1NTLPMTa6hqxjl
DHN6TFteOqFSpjUxiA5Q+QjmNmVPR7YgSTMGSOX8l1MOntLifwWv7D/PX8PJHO882U4AUbHR4Gdr
UdeL9ibtV5sYq7CLzkZobzOO1Wu3TPB/qnovKyZqYOfMZznnNcjDs8eRzKcT6xyQ/ncSDrafxZ+f
gFXcE0PvxAj/oAlsoSo1w/FvynK1QJHPUa8om+scxEPYjM3o8O4cofbOyyGJobbranbr2rK1TkXy
ELUpyoa4eMMxlLBct0VzLezBB6hKHM1rxW8dYJGZj32ELVdCGrRYUpDRXCX/0g3wtR0eH/i3VVL5
M4TtEWTJVq4dOxFpb2lubYEU65c6fISJKGymCdz8VXsxtn9wa6nYy/e7lx3UXwT+WJu2wLOzjghZ
lX60kjxQYsSWr224TvxS2HPMU1my0jj5G7CMThDDzlTcoSTRJ0J0rnG8qrPxo9rcJj54w5FK4jg1
+TzwGJBBYhWjSyUgOh/U6Raij5TcH+yhOM5D41dJ7+MxwJqcYQllXXuMIpwQ6W0D/HAYNYQj3EpF
7LLbU5YfdWh6R0qAxVzg7VKourfLIT8nEaMlA6X0OyCg/l0PVP3LsZ/rtgjOUENjkbgc5OT9lLpS
qWVcy2K5I8iSbQWj8H8XDzviqHX0KN56ftuoCi9gPR8Zw74wChxcKwcWjzwfzRF6Q5oP8bGxdwXX
U5H3QnOANnttX6wvfybECkiOZQKkJ2Siq7/QdfqGOX1BBzAfjhacfbVQlxMxcn1mrXod8shYofuZ
ETz2itraJwipfuhDyk50PJngb/M1UylaAKHPjZvyx8G2EZ6QrU+OUlcYO7/Uw9XtMmytsZHzSXYD
1Wpbwz5Fxxy6Qbjy7oHH/lyqH8qELa48UrGu6hdoyzsO7iu6qrhZKe+4vVeduNedk6WLtIWSfpVf
fgp7gpY89zBv/E7U8J29EYdCaw2mj8pb3+sqMl8Cd8niaQO0A8VCxmiEYJuSGIVLB9Apa0sD0LpD
VRwWqp9KSH4nWJ/zwtcB+ssWwqmdItmZaHnT8GkfT8uOUdFVK9+Xmd8lEcfB6p8hSHvppLULC3wf
N28IUq8xT+rXvL7cGeBNwfXLfNekejA4bOse5YP6c7tgg7BDBPUij/PwGqkHRnUEflgt2QloM50g
z8QOTMlSxqZJeG81LXW4tHvOhW1rWjhPJoq4LywzvylB168la84827d764ZQjQKRhq1jw4VNWVO0
c9n6bUpf8jt58/V7oRkk7DeS0wZCmx/DspmRtlqPemU6TFqMT1uOyBJhahqsD7d4g/nA0eGucevS
G9fWAUoRxxK9G1C4bRkx/EviZ1kgaMTbVkVOLcdpWwNJ72lmveXamem/JqDHnM1+VAkwZ48q9Jpg
ilU2GX4JnRrg+aHS2Gumo7iZp7rM6CW4BAPW2hHT8/2FY8pM2FhzboEx9WHGd152weZ58I08y9mw
W351CN/XWZLNhISOtxD7pvS5wn7+QXNSx+aVsr17bIM6zDFpLzwCjXJyAqKTjgI6T2uRwdV51zhG
psUXNjIXehWF/JblK69v793IPV0ya9mN3ybKihw1acaXlr9O24omNgzzCEw8BzMe7fnlQjDR0L9a
zePAvCux05UpswyMPgMbXhXF+3HQFcUnJRM+tF/e+dV4PhdpW/CpghNjR4cXlzzRDUFMOB00dELQ
blyJGCNNQAlKkaS4S78y5lwcM5X+3CzMrWYNAaCRdPcJi1kN9K6i55HPzbn6fhoa2IXfNVUuf8sC
Kfju+MWSubnIGwUAG+4mVGJZU80+EDHOKmIjV7lWStLxVxFy83M5Ll0fpmhVHNQK/+SQOYfS7Vd/
rnRWohOVhcDmq5PJzVd0safX+ynCCpG57gWOUjsVe8pOEa09HBNhBWbbQJcQgxkei18smxUAE3jR
2b6AEgeydRHMZKK+GYuSjlaWa4IK9rdiPI43491aup/aBCw6dqHcY6D3xbm0bWuKWuIhGu0HedpT
6Y0FzsdVs5WcDFgujfJJQbW6it3IPZImqD3KTpeZ+edSSQjMHNmF2zYBxDddhqFSvkLNoN58g5Nd
P0jEn4c9Cb66osG0I7mgaa5YsRJSbmpJKek3DvU3mf6LsxeV2XMjJA7ITt0rpIfp+aT22HDDccG5
W6Oa+44mM1RYHuZvHyouImh2rDzh+RVQ0k6upuTWA4DRmMOlc7qaa1Y6imP9XfbIG/ByKZK8ScSI
sLTR3kzYpB1veGbpW/Ga9J0AcitOwOKG0GBT/mYpbTXVJeTsISks5mtnK9uXYD3G4RganwdnhgxG
mBsliFS5Vv1XnHbsNlZvEdAlTSV4AtdMXkzHvfCd37iMa+UkHAYuOKWUcgm7fZM6/xbBtgt+QfDE
2nPgWZrVA8czjpB2/vtODQcJHrt0wM+an/bbt6L8XJCy9QWS2651UtL1UPMhMc5NvI60HyJwAtOu
xyCb1fXehOjqSGu3mY3ojOO79aZ1hxNMvyVGQ6QdhrMLz9sTsWjRnPVaVGypJq/Ybwx09xyrXSD+
bpF3g+dbuIt+30wIyq2X1JekT+CWY9MfTzS88GWIQW+YRj/E2U9fwPBV/gQzD3aZlVHLKer6MFVb
O5AcD6Et6SFUFvrl/L8GqmwUrcOJn34R5LvdooL/emCvBy+Gb8h3cFsq8UC0DlMBmTrCJ5NxYNtp
4dTlw/4nsv42bnlBizRu3eHs4+H6591jcsnPWuByeUCcOxUYttC+ESruZY33DkXfyeFhMDuMHrwV
5+cZkiZNmxIKGosdDryp445f7TWR25iBM5CiDcbFgPgY05SZzzwq1JAnNJFL4r7Y1O9dMVkxyJ1z
wGALfq3crQur9eTEAJkbYoH+7LDNOL1aJ1zJUEuDcULAIYT1ExXIgb2a0OcWqlT5NTCjz99iUybw
+7lhEn5Lfc5O1aP9n5+ypaf1vgL2SAaQuDiV57acC3J7pvFRw62nta6xsCC/H8XXorRLPuLkkqTa
PqVnd/+lalnWvb50yJeIf3puj0JmH6TV+4f/Fh1a21o1mXPLr7mc2iWVv6ZV5W53iBB4fwh+e8V1
FRx6WQX+f9hawIWjCl+bqK44fmjvsblw3G232oHz7wxYqzWZrk+mjMoxsjlIdYxJOIpIrpP2K/wm
+hvNzQ1xMhHHPa8ifoYEKonNGsXwEMk7ZcqbB9C9fFBtP3tkgFOtt5mWiRF5ddxmSyAlqu+Zg224
41SiKy9wV5IomMbHYeUCXVxgoKJS37Wk987MS20jyvf29fq3u6C1YT+s/tuYJZDT/RK5ENF136V1
1jFLdKfTiIBJhh9H3OAqebxV+AUONliysYu7Uq7+PgGAMbKjvro0Ud1bMXEnPc5pMFH5b2q/bryy
I0TF1h0Y5+EDrRKQflWgDpw4y56N4jBok7EHuZMahqdMeW7PMu46iKgrhtmjM9uzlRqLuxq7OXxi
/Np+Iln32ZkJgBWPjYm1FrFhi4K/qbqc3rnnIinjkPw1CMOHvQWCnAkgBTAcXO4idoiLYy0wqMlD
dSLCLhsiBVaVqy1QXQIgcGkCwmDTYV4SJN+T9GnFJQe8hPv11NumBaZCzQX6CHze6rJYc0gzjyxg
PvfIPp5XyZ7iTRZkDa8UIZp/XK0KntLmlW01xRfVGISBf9C4JfMokLrguM1BJUAD9GpIWi2EMjMO
so/pBb/BaquMV9qtnqslqtlBLvvHHuIU53+zm2E0U57KahhUccO44UaIqDPRv+/1Ow1Be+TddDwO
+rZV0fgu2O7hwcgahN7MnP3qC5N8ZSyiE8BVWlxUi8VVohyhw36+BIp1VSs7cAOpPjK2Ub+B9Zka
F+XAl4Ng0I27kMDtOhvld4T8dzEG3K1kxuqXqyvUOB3faGZGkSQpUiHego+94u9UlER2u/xIYgvx
vOvw7DJGZ7zfGN/on9XgYlvPSWh8/y5H8bi6rz75znty+fBDxTRxyD0LthKFUIojUThNkWUDZRMH
cZCGbBKxKrHKh+FYP5v9AYIb08n88hfOacaZBkPTkSYYi3mk4cVzwP48hxSnRREZd8HDYQGXw5zt
9zuGB6xkrDiA4Gk6WdpSDsgaBXbqPn7zd0xBLRMxLOliD3DmoXN8Ao/w/ArUJf4i+8apJ+vvN7wo
wZYrgcIZpR9kqZhgAL3CDPFx3By4V7fsXHfoIVyFsRWuDV0X/SF16bCcLouxEIdbdw+hZG9eenpF
AO8Z4pyc1AnMx0c3UFSSrKRFDONOi/uu9QRm606suhuAeUEEibUW6BMJszQ+CJ5GG5nAvc1es2g0
bXg0CB5WpWZpl2b4Zz4TDQ8DdnvXiX2g7ALClS0NaaVxM5Qw6tAadCJd2P4d5F00gsBKvx0q52RP
gTSUhx0Uu4KE7cjxbPqsjNr0f/CWbpOFKarLpCNBH7xA1u113g/exS38fVjOZ/ruGJ2AoHtjLtd4
eQk1Jks6iRAkS7nd2Xqjxz+5nqer4wlHchS6rmeUoxwF4W7nh6jJw9BsCbYxeJ3pDa12GhlQ77yD
byVuao/21fHXWpYjfXdraSuleLKk83ltugylMGnmwAbd6GbKkRbvXnhCPGcOaHLgRI4o2KVytDqX
wVFFgB2DEmOoHYbb/+4ofKiAK7AixBCEsq2sS/DZF40MzDvy2DInSBjwVrH8R4tYIdR66ndBUYt9
h2YCxEE9TzVHpqherPAbtS2Xb3uJlfYwFabZ69QeW7dRhT0RuJi7S47PoxawRZbJcj4ErQGvF6jO
gbkc/aQfcccYmsrvv5JE7OK/ywjJzMMbMUgiLWbKV1LSLnB76BXrWDCtNuSbV1gXx5HkKebq4Z07
OmCs1W+RTeAzfFQrbvvY1S0EmEuINofPNM4oeyUKdDvQfNugRUGgQvKvfeo2NWxJMabFRegg2oO8
QHYocDfh+2+Yj6Ex7JymMZzSnjN99Dv5zvLOO4inGhfwONwf5n9qdNfzbTrLjMYsOEAD4oANNdbl
9duVmdBxPJWa+aIm9DWnWv12JEXkr3Gn8cII+80qG4ulXPXfDZwS6ysXCx4xwpP/4f7ujymt7Oz7
aibvmQsDdi/iEL8MpyFZTFh8W6bD939BnY9qfSF44qQJhdRBh2mgPoZtNK3K2fE2sP/P+IZ7LCbv
STapwqvawx3Hh93gWetBBDOol33+8QK0RIVVi+mscKukIi3A71qBHY/yFbt9jHoAMPVRIXLJIJcI
kImTNBhxXy7HLembl/eFeujc10AmQAANe/QSVFsX8PB8bT9XbeYF8BQTc+LrdqNK8X/UhLJ5eAPt
6YZR9ASiAeoTbiNc1gfcuft3gn31m/IpSDPBs9aYz+kgq7yAfUC5kNgoBxcacwy61tGcSva8OaNY
XzCCuazJnKQGHeQg9bKhCZocerCbhl4mICldHelK2Z5yeVX2S5JFIRzQuZW5AUEgIW6L4bBgfCtm
Qecr+xO4U4l7o7vyN/F7zL+rOup2wIl3C/mqGqzQxKQd2OrmXYQXOwQeo3p37b4T2MDdvwRlwuMk
O93VeBC5nCPRFk/PhQnHBt/4eFDR2YzPaf2KouH2+5t4ES0PyV68pAYo5x+U5O6VrVSf7ZOZWZvu
wu9QV9F3fSKsWR36prGmZHZjfgC/EOfPttr9viddmVCX20ATN/2z9H6pPZZRqb9FbxSR1OWVRIyV
BY5m1BHRSnwMld+PJyandCXInSSupv6crvUvlWcdEv/b3WMdcvHQM4bus/8FjJMrsSE+3ACjH+Q3
fF9q9WP30MI30yOQnyU5wRYy1+eOQWxvGBQSXDzjcxkIS7W3jGHI82wB7cisxsMnDzLU5Tj+ExKq
IG/OiY6Px+3LmPBMLHbx/O/EyQmvKCh8tTvyawoNmRDoQJDSTx6g2vqbePG1VbfOrugN1NeaLuVx
Pf6vYzGm/Y0NrIZoM6evtchzrXwdEgjym1Ill5Ow3wo9BvdM3iN36ZcsvyrezdwcjYdmKJkBwEiZ
6YnIqQH0kbkafXvqPpnIzkq0U3vvjNuCV/Jb0hBWJtJwugmJM7wSB/qe4YttLY1UY8zfGVJmGiSY
RAaRc51S6EvE3yJHJLTteA9jaLgzqsr0DaPFiUvuudLwzZphV/lQVgSCBG4EDwOmyAgnykWG5euW
9NIf0Ii0JGYoG+GNmR+GuG8IpeeUq+VeFlCls/VKnxGB9N2qBFZULydPA6zoDANR6L78lvaVE1fr
aHVCUe/pBp5IfGt8WfLV/xv8NQPvpVFrs6tdIbSEwOFKnmPkWgsrgtuLzpOgetFt4C/56y1O1IUl
3euX/iq7ZcGFz+9aIgoc+jXfKXCj7cUEBkEPNkFVkL5BIHBNoSZUIfJg35AjCNxHc/lUG59xPAY3
sSDysm56hsFGut+FRWToy+qbY8xhu1S+5hPQOfG2jWTWZo9IOI2HDfjK2rPO7x8UBxKO3DO6jhKY
SEGKpxbRTSZT1OPQS7HOV9b+NZYswf1D1mXy4+3b1chRaHCePnZZ+o7h9zo/GnDdnXT6M5/rB8YP
9gFMMqB9U3/0odGfrv57XGlWolBtFz4xi5mqfUbBjngHAkD+VXSaSSnTv//k2UygzbIUhx47xAgx
QsuYZmZoSZI2nXPD397pDe+C1vFisuZ4mlFt22xoAYUBq1XOAxqPuNzE+IPnigsH/YyEfzg5apPU
VZIVf3j+04Ja1AbvmQ6Yg9xA5sOChRGJ//yC7esuOFjjVnb8c719m/KWvwqefTydQfJgTHiIEdPj
WHXKW6nUMNHukXhGdVrs8JsAqzvH3LB+NWq0mjrkkvHmcuc8Yzybh8R+SAvx18FMYRcUEUW6mHsv
Ii2Z3o10nnXcwWjI46aKNYvz4tRtadlY9+OXl/133etPZib3tLks9OhswRzGhfdgiyG5Lo55CqSb
/6WD8B/yFxSzgAeefLVnvEHNmN+/nnuqZ+tCXFwG/qGS2KDFXY2Dj47O3M+DT/dl6tDlnoCYQdut
3vc/SJhOfz5zR4YwPZPAvGLR5JBB4CmgACfiDFgdW8sqWX6u2oX3Bc1qSf+a7huABhePAoq2I1N4
xJX/QFFlET2aximDetjhBE8UOomxOX2kH45O6ALK8zkhHul4kdxmgS5qr0VzEwDskJcrX5Ym7nXz
fto0Ciqf64nlv/eFKj3Uk8OPFV2Nk6qBYYC+Ht91CLB5vFANCJL5iaH8om89Cfj7BI1woRWGjCog
5wv5xi9Blt1DxqgQp/dPw9ZzYbVK1zzGquFjsNDK/jsJh0DYYjYFd5YeYzDgblZyTT9bikfdmyJm
Dc2XrVeFaZpsBVEUY0gCrrGuwk7fzSrDLyJ17u/01JQZ7pG9B0uQYnOGJ/U0b9eBsnHBeEP1s9pW
5Ip6RS8bVYTWAekOGQr1aH6RN4dlZjGNOhTC8aZN7RjFz4l29fhlnP51rXetPO5poEjGzykuljnL
Tn+q2ejXSRi1zqJbVlHm1CcILmHBSURy7q6tYoShMVoljP9SU5On5exQKDSdeClnidjaQc7bW7qS
zgXO1poJB7oMK3vgf30RU+phgMuMKXy+pUnHcnQaCpr524DJAmh//scWJQfoPFI+b0Wxq/93yRZL
1jZ5yftoQALt5w1fMJZ5Mtyv64DBR5Wm0ztznW2tGSeEolMTR0DfPqzAc7u0zyxL+HM+J80XaQjf
kacZjWxzyCcypLkN4mrSdzKGzaXHBiwYJTIDTMUbDR5q3GrT2PlxaZY1rJCW7nsnhJ0zzKZ9prqg
BVw0Il6XLXtoR1JhrVLEQE98Nxh2Wa9JxzOJZHEnCX3/+CpJb4oXvj9sIVli3dxKrMZJ6JdYdauk
s9zpyh/N49Y3jP25SDeQzPRAaEfV9zoI4VGim8DFs/xz9UCJuI3+PE7RpgE30lqFlrdVYaAqcVzI
O26sKZvgxp0H6La7nzfl++MepLBxCSUeXgyuWcSGV2nN0PAgUc5A58X7ZT1wgyq0avJlDKVWYH+O
fDpWFro6dr4MeI+E11vyBHZP1LxK84U4B7fCvY9kI4wM9PpWK/3dDRyp+JQPcRCUHOrt4tkVMVow
7YO+3gvFbutVPq3kI5leINBOdDR46fhuig1G4cEXkH8PfcJFL1l17Rdu86Oha2xND0QFX13wtTne
Ow3NK/D+oE3kGP/ZMVBe0IrdKW+kEAblUNNnuIjzegQzFwz6cT4SbdnvdGSoBoG0rhg8VpEh8tut
nDbqwyJHCgV1Hp3ml0hPvqSEMzAARYdQ+F2EIBgez+eCLnyo6XWfF1Z79hHTy0m6Nu855rDWEwI5
xkuBitiF+gsJBDczrYvowcsE5kedTFtv1VQhzYIzqujFJrzoDl86LA1zZyVJocKIAbVbzrvBjvT3
0QSSTkFuxw2hWr0rAJone78Je7Me7X4WHuKNzgHUUWTpszF61dSRG2zml7SzQbLhfwguekz9KApU
8h+0h2P0zgI8w2g7HsyXZKkpI7RRDxW4IM+k1aaBHDE12alY6VemdoOZoM5QhyqEouv6K+jF8RLx
kPBCuzigAk2Qr5TJh8ZD1Caeh0Qtd2E+epaYG3Gd/QTqnxpCNAGFITWB5cE+8uvgvNOJ8izxXR55
B8DPmqQoIEAHV036K5+orTZq4GtFKUIU15HTXbJ/0b/g4BkcmwT8TdYlTmPUS8RGlvm/gdL6oq6M
qPdRlQu0VLJUQUCCnb0dKKBYXXYzu8hw0J0hkwH6to7DDehlogrx2H9zUjSi4qZ1Ct5dl0bJMXtX
2eS74bOlM1VY8xi1zoYtYxieN9IZNy1/AP+gJtgia1AU686/1uhLDq5iH9bPVfi89v1x3pySjkSO
w4fGJIg2RhUhNDrAi4cgtTDGvuyjU8R2Oa8VYjOjdDOw55TeGmGqIW79n8JRY1dXBtshRT/sckIV
aOGT5J4+3TIDgBFs+UObO4cTwll2ewjBipT9DsaOpZzRE07g4xIev5Ug1P3kpsiCDU15xCgurhDX
sy4qcpgiBxNYU6CeWsDMfgoF7HiIaII+YcW9riDnid22yCXAi/p/BpBMYDOGfS7oXtOEhIjKdJCM
Y6g4pLA2SVKAviDOSWiZAR2oV/8vbAua26hWeCcwysdkrIeGOsdoW/0d1BOh55nCHSXF+fvrTYR9
BQFJgriDsOSAVmprpZy+Z0eh59z/lPRRi3BxwR9yoK4Sij6cejpQgG7hAcd12ARKagjlY8wQ3Vkw
dwsd+oSKBhATbg8XhtGOI6eiyDoVrN9dvpmRRlZzn+WKnET51xle47o0dAsx+Aysjh35M/kjtWV8
2HDE/a3+AbQZyX+HaWvbCJssjoGObU9YU0czkruo/AspwjnQ0f2sxfV7SkDaNlesRctCGy5Ddhkk
jrdoSw/hgDu3ccDsTHWYjn2BL1C3BBH2NV6eJqzGzY2C3Z/XZFTeoIcvX68wf580B37cl0uPWvNH
4ulRU6b+qqCQS46y7sLDpVi0nZOLh57cxTcmZqAj5xY3lH5HNN9togdl5hGkvk4hsSw/omZH3neU
Zkk8/qp9oqCgDXb7BdBopxJmaMu/NKkuI+RC4J0j1ViY5N22rQEbQToLDABHd5og0X8os1QanKXD
QUW3hQgDXm0ujXLIgUE3KCNLZ3KMXpbX3Ke1t3Y74ztYtspKET//DEZIjFYORLIV0u7HcBdQLa6j
AX0bvMcY8Fqlppny2m8pEv7+ZVBmAkeKcQSGf7lROQd+FddNdwrd9eUwHQmuJIMx+QuXCntGVeSo
7dvTBGyZh/cMOclNztHlqQag6y6bb7nNj7ek7bRWWkAmeJKojjLdtYgLucFpDT4kAW4tX2Ekcfiw
+qdKz2qPGVsrRpV3j8G0w5/BHNl4TJm+qu4Bx+TzV04kGM0W4my8anXteBdq8XlgkqAc2Epr1SoA
T823u01obqjseURKjuAyoIP7LTkDfbJZaHvNXlo6DOORtDOVKIfVOFXHqAxs5r8Aeo0CFTO3kQTt
QpbPGHv2QGMji/SUjFEC9TcQjxrtrvH3GyRILVxLDeGvn7KGGAOr9kvaaN5L/hvz7k02ELx8uuQv
CbL/ryqQT1NjUhu2nV0Ba+IxGok7ilnmx5ERQspXXazA43LowEY3wTyU3Y6Sp2PBprA1oRQwEGoK
deJcr3G6MdfA/q070WCzllGgtmQZ+mHnmIf73Bq+PMJx5kyej/M7ARa20DbJE+olUpq1qHPAOscJ
2gm9QZ7UKWmfa75V6UktJZkLdXW9PdlbiYkYppKPIA/geNWCfafOC/V0YAyAsk3nrA3XaZzzxJGK
VTO9Tmt1phOIJjYSMTYdEamWNuld8u8fLw7ts9eYNREpAcuIjT3Y2FKx+ljKv8Z9cm7eJl1JwNsx
OTROgbD4m3uj53DA4cXoyVVyzHJfKIcaiIbHGpbMwDKHkkvkJaM9eCla0jju+/Ebq8qRJLabMRDl
RSDxyNJonxgi6zE96OWiUon7ayKoDEQ3A0ywW4hUgqYAOhPXzKWxc2xomITKx20wGxs7Uf6akOdS
VICTePtl9x7vm9rBQhTxJgNKMeuZ/Z/XJ/oKg5P+mRBnLqy0QlKdkxGpRshpV6XHzhvgF22HgrjF
7D9ExjTXZNsdb5tVpejHZFsjcTOJYf/B//RO4ZdFs0nVrC32v8FZ2IFqlayi+XXSNMETw2i9n8Rk
aqU5YT8i4TRyPtYwZKg6kSFeQTCB7vY6RZKKfhts7KsLVRXDmanWHA3G1YYcr6+5SIdFir2hJNk3
ZwHrnE6Z3v4+a7dgqmlvWwqZii7HJ4FfCIAQWw3WEhqu+kMyp0XEw7UJ8J9SZ8OhZRqSzl4/spVD
i8Deuc2OUMhVOtBzDb/mmLMRsJdq+7FdOhiv5ELknSPaNaZe0WX1u61maiYvH6z2etAUZ9vQ/nqo
OUHcNkBU5EWEVqajySEfR8BX99qxDf3mzI3BC+hLfGsk4y37lJkBJECS+UniVY/kc7mLQ+zkPg3s
fozftyuahzdlqT6gw3iMPW45TMaSm8NXYe7bJn6IVVD6URwYX+qPOs0E0qhaAy/Q1D1jR84DVHFM
NBTvB8mY9L9O18nRFeKQCGm2BmNh3u7w73OEwY/uKwU45iTVAtwh6J39VuUh1JMGcQ5Di16M68eo
Q3O+2zSOlsW214PBePlDQxekpxczeKqIBXNs/zH9yoncF+KlXPGN5+s2R0GcA4OjJj4chK1nhzXC
lWWvfHB6KGNBdv5RF+Qv3XRRsa0g+d/QOLlWdmVoEn2CbQ7Eidswdj6JG8OLof1O8LcMtoybdZBV
EjzbHn+q0xJX6w4oTqsaDWLdo6GMgj4BylTyr/v7WW5GRJ2LZpSLGu8OxFDLeBJ6NQMw26FVRoIb
PQSAId3FED0qLBUBrKoCqvxaKaX/GknqfFuGD39GZtDVJXLdbWIXE1qTi1sxbmuCdSVegGbpHP26
/M7TW2My2hNPAHB8RryJz2xH3QQSF1ErjCn2jF/iYGGs3eGPR46cacKVdyQHSSkL/dBV42iUksCl
RfU6XM5jr/tr+fQb/wxY1cfOEE9veX3XS7X6HRER0JNMX1f0s2Pnjy9Yh28Fqr0HI4NAqn12B/1+
zUggjmnpDqRmYkExtcGwcQHqeyilEbJdm6bGtiTXhDJiPIAnjUC68+OMXddLoqYT6KBgpE7GA5Fn
TMqq68plSUOtKJefWnUDcZM+CeKeVdFq2aQLrNQ4B2EFsQ6Sz+yv6TbYxssiHkyxNPQpaBxW14Qa
aOB7lxuUhNSklXcVHLY17iIzp3nqMaKcEPP1fOUYP8qkwjfv7WPWg/Ok8FdZfjwp1t6Au9XiBhyL
nTADenQBJPLQC35OWqk6hwFxbjp9aJJYKapW6yBjR+14D8+eNdabDoaJIXvzcdMnW1Kllb51KDBs
TSvU0sQYjLH9/fd+ccrexX/yo4tOm783cZWImCm9soGjFzrUjBDmMpTIfiE5EwTg3Wkg6lJf06Wx
wPLak63jpIUy5jeezowfL05o8XoFPccJKvGUR9DPeWo0KKZsoq3WCpmtNOQt09OldcQFHrEM2syC
BBRifbw8go0VfScDmXK3INCaZObNkwG9frNB+5MIyBYvo/qXQ/q0pmdZDSMFpzD52HpVgDLwjgS7
q+iIwhdA1ekTaxAwJKWh1TkrLnHNuoBlCVwxR/NmztKp6JttOKBhmloBzM7c4fyiswuqF+XwKwV3
14Tto+at3Uol0h/uvsZUHGcjxPgpn/2T0ZlYlPNYThwAv6flCnmhB6LCv/4eOQyVhGzZtFXDgMH1
rpU6TpfcIKvIIaXCkn6oQonutbZ0MXL02w0pVfWbQms2pt3SAWKoIJOhYxczQoDKuQXtyUWWRdsq
zlW7uCvXbptoFRw7KsrKejIKXBqvZyW1K/XKO6EZMJrz0w8IU/RQIh3vibMDD82h5kUZ4KjD3Q+Q
UdoI9fgZyTt/K1qyeoV4BPXMubvaGZbfn75beu3GxTGheGCaVkOOexbrotg0aOQwGgH/UCnHbx5U
5yLokQMQbuXdNFkhzMv6iPX2FJq6hNSVC/ejEW1MoSsl58lkxMzWZyqhwkG2SHh8zC53um1RopfJ
2Px7BgcMHx4dVPCSwP6yrjWnm403jUuZ53I6e3EOBk6TRWG4W/j+TO3lbLkjHn9GPNCB+6uLRCwC
iFE/X/EaWy9J4rpnq9FlCzanZslZkLkT4I0/TeVealqDYuOjQKUN/mQL6xP73wzTLB3Z10A3PRXH
6HJdDz1q3PFq8bFiPRchGjH26idhu7VMfHPD1OqEecq2VL03ZyF4SCkC0SRBogz/pBWtp4iCZO10
SOq/OQuiSIcyHFFOqeEATgw9DhgZ+pccCGn/minscKNhBrmwf99MD150n/e9UtZ9k12jUVy+5euT
1x+wyqf5vEZX+hyzTsWWa1djv12w2Qj5e5tg7RV7hRrJA6xkcCqQxKZ8ZUAMsOYLZLNq97BIFRD1
skNrYvWolAKGYnMOtp+z+JiupOhNsBA8kYmesgVtV2bgxF3aqItV11et8d81x+BMg9QSrJPFNGUt
XDQ5NGHF6zxSDHItre6zpOxwUdvjZbUkZNLJkJ233yxbAlqWLAHYqONu1Xjb+KtJjFMxbNe/JDd5
5lkWm6uMVxNKOVckjoDG5F4yWE86QGZ+koi/tg2ymsgcmcr0KSPPx3DOpW/QA+urANLE/rp5mMVI
W/H2N8snAFQ6pHjG0J6Cp7GP3xBDpZolIo6MD9l4ngcY7bhFUaC2yYgujbms+udR/ndzeGnI1qax
p+AZYNpRtNqevaXNorU92ehev+Df8E68iinkFAb9pFSiz8qWr+N7Yk0IC14YhZyGA75ujy01oB0W
RXcJkhgFh9xhlUzO6Fgwh/ekqcnClHU+ONLaR3Drd0GBj7kMPOvmwW/j5hvcQyUososPFZ/0kpPj
C8mWmd3095Q2QWkfKid8VC7egMAtMVb1ldU1nUNW9UAibkf1KXoi+p0X2GiF3aRFA2rojc7233K1
ohBvbxmIoshfWk9OdzOmTC+sHe3mSilepB25YqzEAEP/qd4CN4YELQ1DFSrjdDE47bswCbIjC/8M
RcTqTyJm32/sa4jfciRBiCdopRQDjxk18pLibDibY9hWpRzPeKSD0RmqdQL4NeeKp797T1E8xFXf
D3I+BDA+G/sJyxVwNx4oMCwhGZQO4BUX6dZowmksFu69ajyMnvSwA14jsMVT7e3ScR3EYUoVmYKO
h6OkMzPOjRj6o5CclGwFTFpLdSu4hRM7tyED10cGy93LSj+ALj9KzWIuCdl0vf6cgpfQDAwWTk+t
TVoi6OJPyc7Hs51dBD2ZVW+UoItfCarrPKsvtFpxqwSNVM4HbCh8BSd7SCjoSrSX3fnSI3Ipm35T
aO/5nQWruwufiIU0egBRWSkqONyuu2feW4nsqBGyFa25w8PQndaGmzEGNLXV+eiuCyUD7XxQ34T3
y/Sk5lsQHtlXaZap1bGOvh8KLXnHhluZb9KapyFDZG3PX6gzoIteIoeICdrBXGRY02et1cFimpbd
fKLKjc+II2wFAHWCeiv9mDChiy8diBEkUg1Wbh/1SlYf6BLox4WGxnoviJvSAwwEmYK1KdMgzMJi
iBUPd2qgpAKhvE/pAf0NOSFrCYpjZGYRNyW54UQqCZ1HqhhGMih+kmtdfDmTIZ5zX8dSy/rCYnAr
LNMapLxo/eZxycxYB9UkRR0CyReWgoNQ2x8qUB83e0/xE/y1oDvM63BxNrYsdX7hds0/f0HwfA/7
GKyfyoZsc5djOlOp92e7ptPmRe/pI1nw8MfHA21Ty6UudA3vhtyVdQHLTuLmXonbYGskHo3Fce7Q
DAdgYOZabpAg6ZZNuTDlDIWchXsbQ6JHcAOGcqSGLfH0yhU/salDgZHNfbODqiJ3SP2cPSr3N5kH
5VKOPjrJrqnMKS88BChdyhm2IyUlZUC0PXXBk6G37yUN06qWOVw6Tu+PSWNImhbvoG/VkIFY97N5
sbtXSM2hwkrHSG0UJgMdqapf9zyy/bR143rxT2c6TFKliJWvfqPmI65c/PlWWSNSBY/zjUXdxFDk
nQDEshm9yU4akM+z1buF/HsME5G6A8SsmaBVY0zVReqkhgaDENCDrtlIrlPW1pAGjny2vnJuQBIF
mDVQvS2Vap/2q/N34z/cOzuWJ3pb4TQ3p5CBoLdQXCBfP68C4GnjubQ31LYmxlEIWzJD0KKm61yv
FO+vKZLKSf5m9/hsXFtXElNHIcwDv2J4NTVeHPgX6qt9OhmqrSUuYjYN/x5QMNiLg/5FDLw7FnXH
cU2zC9qo7OcU/hCrgVPKDLAQ+Qc/F94uGgWlGg7hmXicWKWyJwKm8DCXE7as4satlwVygpWM2s9R
zD4hOkWKQNTDQw2LmFUSVYRG26FYKoNGClgKq4DtWUzu+mZkS7NcgVWdtLOk+eWvorG+OGV/tNsI
qUZjO/+uA3S8L6hVn8umSfcVQQPaZm+00l8B0GUNV8PLPWmu1Elv2wDz7BxtrB4WcbT4ma7P2+9o
fLZjlTiFYebX0B0NtOxoySlSWAiuSreuRlNU0UdxEOAcTgPMuPGOaSLn6Zqivd4JJAAhkyxKNFy0
hjv+d9sIC2D1kB7HJMXtNnfIRujZ+f5VlEH3N8zsp+dZZcyXx0J5B1q855xuOjYm1rH8MjYPckyf
C7hD+a99WqTXKQ5J7v6eOFvRJIqRAHC0HecZpUg9e1M9Sie/sS4x21iGBw0ikUg9Szi8Z3rrfUAE
JKNP6d7pYPYHwBHYNl+9GjQwGV6+hvhuBcP7SZPbZ84t4htkKSgFYul1+n0xRBzAhu2OEND/80/0
5wxsl1dIk1ATl6ksoFxjvbG5EqElt/5bJarje2arbrXTwPh1cTxg/oHUHD/eGXrh0sL/85mP7Asr
tx76GaMTJEXEqwpSAnGX40Q5dnzXNjS031zMI+Cgdu9oP1Yqmv7cyh5y1+fA4Cpum0dCvsnJU+iU
kfpY0VXq9zV9CTvEbdO3XMz2zMCNbg8VAcmJEzlVzyyayT+qfR0ky1FsSWlCCV7LHBYKbxoF03Kc
g2hoTKyYOQAWxDCi+XlOJD0tXmJtTyuOlFztpgH6VtkNUNYkpcumlIvdovTecp2BC1sUtAzzBHy0
PmWnW1XsEOSQbGOeJfjWy5fYzIPqznzGOJ7LpOoCuNGfLfUQeO+3nah/PzznbP/Y3QbTqOMGxLRz
Rkl9ga/293UpqjLhSBnXyH9JLUkKoSOAk0XspBuIR2OSkRcylQRSfbiXPzp0Tzw2tySzUbkUOIsz
Aj/QseZIb4XWHnd1Eqptbbc9sCmAidMNDmyYcGPeWuScZl3K3GDbFq3VcmqyciCWYgsMccEyodn4
XvEf9WwWlNNbTZ2c3k4MN6aIBfuhKPQvGYx7o7y276DZqy7lI22gqJgnDoVCbxtGVThIzz1leKim
03M4q/qhjULI8SP1zq5hNqNRLLHZYXDjiazMfCpBmrjLAkd3vJWznavNGIurZtldqdWdvsjE/4pb
dhEVC0AnDONo0Q9K/a1fJWanV9J4r50zCktm70OJaZ0Kg2ZwWO2aUicMuZca9MMMG/rkFpAyHzsv
7aZKtyG+AJhrHhc6b4rvjPxbusbeYcg19uwLiiafI3o8Y2lPO3KMgY9aUt4M7wlUMgJiiDtPRewj
hfFFkm+byWdzg93lCCv5Z7gC6JIClZScbRHIQWMz+uXTyh0qhwDRw8OFly69tLzOl2odIaWT3VPf
+9H7Wc3l1WUp8cvNy1YVSy9toVaXvXWR1+XbDeGeC3Mz2lY8XpTD4VIe+oiNtAFwhdfpnbu+2Xvd
CCqL0vOKH9qchIqqYZWi8C+Z6YvjhySygcgyG5oUUik6QPMq7ggEjSUBmALMt+WLFgqwfNjOkjfm
LCqF9XSL+cP1My5a0kUnSL7lEQFgFaOJr6F9ABfiq21TSXC8BiBX6RWlg7yBMVxq5OIxBY9+SXLz
nUMUeDxgj34x8h9xja6a6v8C9KYQYlqBbkx76dwAteJ8wLE9+812CjptzFMngixrZV6H96igoMZT
D3Lk27+4NtzRe6uQxuhorA9JJMCQ0C+jbLtstJyo9JcK83TJQR3nniTOApmZpTTxu8Imgq3pWGql
he9OicQuX5EDhx/7DRv7ZUlhZz1dt+kqedodLMQcs3fhJLI7a2dDlDbpkUUgj8wjfRn5eYqqqtYL
EfG0N+eIk434BmhkoYHxR+uuP820EZMI/th/3oABBiKGPXAqoyjMctfZzJ4RzYlleg6CMMkPWx2H
HGHbc24jHsWpdMnDL1Ob/acS0ds3q5M1AGmZgAdf6l3l1HVVEFkMVtKmBTvO4geubmDlQ1OkyOZ8
iwZ/iL9DpoD11UiJk2WWzr7S7Vs3mtI4gOeHQloe2SRhkdvzfa9Fe+yo74delPMOP8LQKIfeT6hU
7+wZA6mTXnHP6xgxzBjoZOvQDvtU/NRVU0QZJgUCf8La0nAFqeEkFxWgAz4WDYOWDzpNbZ84wuFT
XebeWMiVf3dPnYnUGNfj5IdH0y4N6HOsbATEWkVSvk6ecKML3M9gPcc2UwG06rMUIkolxjG5pnaP
+W1lBmKFVA9KY2atFT0P97Nfe+CBd1MBkzGCrdTRjVsM0flipl7YUaFxqPyejkQyhbLPyz+W2/we
Kp9RPNbxdKK8CeNH9+q5rh/K+SY3Zoq131tyJaCoeaXOCJaHVGXcSYt1BXVRGmU7q5sCUo+F7sVX
XszE6Z5y4rYw32FW2QSivgNOHsikSeKDn6oLTMBK+ztsTOXoye2Cv1d7w2tvli6HX/d3MAyCAmdv
K93sGuPAhHrMGTArgAItYvzTM9xy2pImcj8vOs8uzrsTu7isCKL7ZnpQVPOI2bMG1fGO2HutGFqN
uVZMegy0066k9Qmqn6nYIy/lUgZkgyk/vcyZOmkgdS+SpDL66kIvh0K6A4MgFhVFbth/nidYHnnK
HUy8oNp8vPESvfOFDCIPWckxShOqagVHpDwYCIbRq8MskKVO5Ua0Xd5gooCvS+PSc5CvhbnpGwUW
YyQPId0aJa4YCvQ4OkkGen21NKWjbcaq1G/SSMUDFVUAubnQ70PlgwFaFx0nEz/6RB7oTsbmMkIw
GFC/hMFpWMZWs7wpFFha1ni5SGKwSJSdj6EGTU7yk1OQlK5ksHGMkBr/KE68U0RW6r79+Om8iKPX
IzSnv2u6FsIYTeLBtY5aLb2scxX6iBmQkqLLcEkqUxjYzfOcZKPWLdJWpiy1ar3Uu2U1FaW5Xgd9
KW4uyVEn/6iotAo2Xc+69uNfxm5S33G3XHmxKd2NAWNOEuHCI2Q3xHCCEgn266RgiZ58JPQ2hhMV
cb1yntOBlnxGwsbP+bF5CuvUeDQg+0S5saiTmOnMWpOyBfevA7hNDLXO/AeqwpYaOJS7XJ4xyrpD
3eijvR2gVeVIax8jSmLFvJit/rebGnvnuQL+Dewc2U4+eDT662Mw5ORh6M7WGqhsKX/nOXq07Kg7
AYdwohoulpIvVuWNtsQ3TtIAAiduBXv9TgjSguXSiv5CauhjBz1kkIka95igc6xiNxIJERT3OM+u
t6K5p/EbH2lMFSD9t29tVnYDQ3i9vCQAr6StdpkmtRaTb7+E/tAOllV830o7wXiD5oDGC6rH2V/4
tVfS0qIfXMVDnktCOi/wLTnzUWcILxIWaBnXPf9oq+g3wB8oHQuIa+ZPKWCBwz8ICLt+4ypwiZqj
QaV9XiqhADFxF9jg84m+/hSv9mtkB2HYRWZI94MPxB/FMO2ZmGlCE4iPUzIf+43HCnwxN4LMn5WA
2Ey8uNURxDNm0/MVszayG3Cs2n07mRn2ue0IZJHge3uECn+wfkeP95IQI1OiyO6xb+YWQMeBkX8R
pm3vjdmHYkLkq58X1vD2hQ9uOamF5g/4ry0cxuRzWgXlH3nK4gg+a1vzOGYZU0DE1r2YphEJnP6F
88XnpNGyGh8xFKTUm0Q4GjrA8dFgDu5JguxGkAHgtWdVK+fTFt3H3XwVOhzHOYjAQqbe9zKkC+iT
doKOeYidPrMJ4CoWiDptext0I443doi5T4yUyDlJpJvh5uguB7YlnuKsIlOWMmF7fj+szrQFQ2Ej
p2ZrYR5+ziciT56KfQrUAtKF2CQ7BLzW9rsIlJDia/YTVa6oYTlnZTFuEoF8/X758EaN8w/2Uo68
kBRF76LQakSY7F+mn8f7nTDAz7ad7KBRz9F2q52N5+3aZayqRz0LhKAD971H+ApPoWviAbdi7aGR
L+erBIDT8zwUjwoHwkpIZF5KvJ8wnK0wB5/YfHVwTfky+AsW2d9Jg70trCoqAfJVnQzluOMSDUHy
yr2L81qWtdeBgL25v2p0nZb5Ebw30Q7FJlsHAEjVm5qNd9G9uC1FKpin5/3VHILCeX/9zFfu7UFS
tZ7qejLPnPtv8qwjMrbPlaNVHOefcUTq6nZ3QhuZHr+wWw/14BqCUX0or8+2SBQsO7xU+C1mcdjo
hrNFzjnpASqqLwUU9v2vTsxXxZTCs8B1ZdGS1JajGDIXPWxBt/tmPRernXG53CGTLfRsmfWooatP
oriNF0jABtk9amdLy1yyBLuGlPYm7N1rr2fb24h/KMCuQAjQo0OOXRHNL2HY8070aZeL1jirDDQc
QKn0GYpYvbhuqXsGIhDUYqDM6AxFA+W/c9+Uh68Ybax1l+DQCzRLH5pnKXFZigVV84ukBrLdeNFv
WsWZ0DvZ1SRO+n7pLEAqHGOHi1ECQMixD7ftteGM9DWYRnhlsCdmDLzmzn/X43BI/+fwh90J72bZ
7kMfux3liRpy+1ErI6Fz7D0UQVBnVChxLlJyObDux1+M4TnqcJAPA9bEeSwYen1LlJWPOCkrAS91
q7BlP7DWiQWtQjbcpsRuoamkcs7/8oUiuSWlaiQ5NvalBq3REbxsmICUs6E5yBTT0NflVMleugBc
13FNEpb7PTNMPaPjqWF0kp32Qe0o6jH+wSsi8NBHBfUAuCqCmWlypfCXTOKbnAdGQizIlU8juGZs
Dee78E2QaH5xkzKwV1J8lZM8a/1rbxf32eoYVzatm1oMVdXV+q+OzmTfLDiuHyn/Ar8bCNjClPow
nfGQqEdue9hO8QdVZlE8xfrECrz9V2ZbMcAtseLG5H42KD63CwGpISwCcmvonCVOOGU5r6oSMcU/
IefKcGnL6OJyqKe8IIHNXxUTVP3hsU3aHTJ67wUSvZUVSQjI3f+ls1uPME+2ulWyyZW1s1rcy63/
NOtSELCXhZEYAzAuvN8n7D5Oga+/C6aEshNbaq6mL34pYR2w0feHhPBo9F/0OM9H4UBpc33yYGFC
iLGn7AMJdzdI0hpj3PiLf5SZdmyj+N91Nkm1JonvjFMFewDWt0jA1aYf4vT+1nIKZoLtezDvZGba
VRAdY2OvHVRTl23vi12yCw+1B/MsPFUElFeZBU0BjZ2Ki+nZe5I3FGJ0UZ4+HVXNRjc3pwGlskIy
rj41QFtIJ+tSzthrVFHBmBhmEp2YRZSQ7UODL6UVSmRkaJ3l+huJsLBeY3LBsDmtJFjgGLDA+A1T
c0LwhToOaR88ciwtnEDUxpj/T7WYiIhApWQfPHgV5vC2UVD03SoBoqU/wbUKJ/i9opupGKOgGqoW
kOy/QDGOFkyttUcmcUQb+n2MRel18OuzSM4/oVBHm6YfzK+EKTuBFdDKBLcOzUiLbchmLtXaYphY
NsdK2/9Y+Lnul7S/SIY6FL3OYCoDWuza2p7KXAQF+QHCYU30xLsIp2MS8gpK8lNJe9M1WogLBVk4
KdtCptXTWXfPmr02DVxtDH/f4Eu4jGoci6y+yqv/FlHAcRGXoITzMza+VLFK7jv272ZYbepVDBvn
lqq2ZzhJMmaE2KXf2VESS7s4q6yCEsrXmUvJDy3OnCKEQvjXcEPGoLoOkNpIrQ0UiJZvz94/4vDW
XqGLec9ueyNo3QNkVpYjAXseHVqrMU6PhBVWcmMQ6ux1+pvZ07in0gpwSi278VBCkjwPryUxCMOY
GCJbk9KQbXOD/EFBpWeOFtSkEonKs4KLPP5O8GE9zJYZK/rEjZHY1l+fx7cIQwKvHiQX8mCGbMiO
6vyx0z2mCG1xFYADnVMfghNqeD97SKwjJZUZ5O1CfJ14VUckqjIHfBz4ytxlYJRV8bB+t84aSMD1
aICN1zPIHkU76zi87OTdPY3zk8kH18IDy3zBP/sb/Vkz4J6R51up7R7wTuiuvFkoliSxOZf3R5bg
Alx0tbOcEFSKvfoYwLkydsjZdbQDSZrjSdwG5PHyR2Z4T7ilMOic3AuD4S76EuZN29L9+F+Q5RSM
/EdMgoZNaHCmAPnebtn4LVX6s/gL1cA9nqhfHvEEgb3GzbTNloRNSe48EkBoWqu28Ixhj7z05xDH
6MOvVmhMEU9xM933XnqOUxm8smj9W8dFVy/fcSX5sGqVuu0FDlmSflu7EFxEzvR3M3WqX+noCsGw
It053COI7ai7sqMznCKOoHP0k/Qw1pJefWdaJcvn0o//qW5JqxCgdu8nI9HV7Wi6HidMs3El6Ktv
fChIWNPnHmoiW1dhcTMzBdg3OgO7+yMdIrF3+pn1Hk5xmAIzPXLbR5YImTOXBDFlVL2xU6V+VWL8
xTht/MQJVPNkRcbmpbebGAPeeCMNwKmBu1oK+rOi7id1K96WgenY7A/qs6Arb+3HFA31BpPsoH84
YvTuxkpVJwTmP/RpIg9rbytGoWde6jU1aisKF2sfZCrANnjPwhDDEAckcWMcI+NPAAj2/Yqoihmx
cSyZC2nQ/uTodE9uHwthtUi217glVTfvrnbI3FXJnC31dScfXvOvGbfdTJ+PEKrWRzUdUCap0R3C
ZAEvQedFSP+xIBSAydV5Yd6oh529X03uljt0f8oG6cn32tc6Bryibl5KtTG0TCe+dTNV6eLXSeD7
BOSHB/F8jVQgWkGAwY6cZfenzwepwp4FuEQTsDCO2Qm76AC/QPD2UjOJhzK/ZOcnInjqzbvCfzcj
9ckNkQhkgVCaOa4OhiHSkhBNHF3ZhYQ2wc+3VZ5LcOSaV+HhdjF2OF0UawFr/nI0GR+COU1EqIMF
4KstOs6WAy2tMu/Q03ZXItT2UmeyaYnUfdCDNK5OP6Fl/x8dOtJBWnyz90/oQ6Z+gAPEAAIV8fSd
9nit4dqY5RXxDOYDAPBpZ8Eo3ve700d4LCNJaO0P+u6gPVw8Pl0EAEe5IoQWro73x0gf2xNUreBA
QVwr3JBxEPpFagypfp8ffX8Y/IXxLSwBGIHTIFb7mym/rT3hP+q7osbaLgFWeo/gqkQX/MNBfU1x
Z5RXbbbMpnAz5DkY3XHQPHk4H2v6ICGCbnXGmdjN6vLGK6UjB46vY92dGOqnokmY6BYgr5Ws9HAf
M5mq5hB1xcW9qdvJhL3Qi1fDR+QmFVIkDgkWYrvl1IIh1puad+Dp7IbhlARDksdz6yVW1RGTA95v
DRVMTsOxWp0GJDP44ISxoXT5TWY/Mm2mtm6xE7K/vdGe6Dtq1fcX86MG61IOW3NCXzz3/i8tpBBj
ArP/RCKygtKOump2Zo7LHQEsOwU3pBcRaLU0qYIcaZv8JBi12rGmUGJ+umGZl8wZ+MbGucsoTff8
xhVSI6QtJFjJlvruARJqUt4bIfX8xiASHZaCBUMOP/SPvDdTXqeXWaUaTFpTUfdWk9A5qwZ6j19/
0JuvvOsbVGyqaKN+raiOewveB/ajrPze8/vRHaU7BPOuFxFIh+hmVeSTOC5UgZRspf3UBdK6zOAC
y8husch4dJoQ1nmML9xP/9eALcjmCr5M/nHQ+4NUh6+RA58sSvoZBcSkN6SZuFwzXAeP0/7GyN0n
Qprh1qPIUMvdsYm6ar40d35iJpzHO/huDUw/PT3zw0d7MXsuIIUeN8HbSGyT4QAAzYpKXQ0sT48D
xYfEZ+6+MMF/yOv9+TPRy8twhXcXXSXXdk326Rq6FTCoaVKfJKdz3unjLeIiUU03IUX2eK1ns/av
8JC9tGmx0EbJTtZ10KqhUFESqVE0r+rptXoN9+bnv//9vjcFNwXrrtNnB7ywGsLMX+N997afnBRO
8MHw6+c8cRshjZETxG3MOAalPG4HMjLawaGkzBjHvlxjiVPQOozaKKkOp/3DyJkVORiJPvch31FS
tH1TKENIiErzHbKc8foVby5ptiliKToEfAlz/PxpN9lNSW/kgDidL1tpYT8yOyiIHBrKjnShDIyV
F/SWEFjIpKbBhJ2U/uzdVCr0zeCaAf98rJg2ZQ9UuFXc3VYyZo5vZlkfiuu6YWPgyB1hIwSsPacN
/rCQJhh1Gr0smvrOug+wFWDDF6yW6EN7iaSo07saETHtFOffawZ12jhFICXe4YqP9EotmyjDFaP+
zYdW4icydZAAAf/K9BiSNDZnX1JFz/J9RZEJy53bICbjTPAZvLNRqZCGbAyTTo1ipOJQYignei4L
lERL/2YU7p7vfENafp2uMU+M3wou0h5hVOMnXEKa3h3muJXIGQngfmrq2aKD1LMN5TDMZK9bJwjc
tpm0NRhUqr1xE1CLPLfxzasifXAZYh/c3utEAFpa/hI8KCOK7g8mnYNUJRNK2fAb4wKD05lCvJH/
ipQGwXHZGTrYQJvm69/EI2KFaEhhjYVa4Kcx3L8tUFLlHHmROdjt14xFkM37IQz2Qq05njJk+Zk9
hrwmN2dQMifYu5HGt1tvKA00RPrmG1fqy7NqjhbvcuZ//Tg9OYEVvumDqoME9E0e1aUWa9LyhT2z
dj0AQYxrk3UnhuY95ug3ewSc6jXg2vWxKmmmNlcXHeluBf+748hQqanWlbppZ9jRwCY6lQSPjPZh
hxxtz63xwPlaN7yP4ULzBGcqnvEux80r3eAWY9C9SoOkKUoA5pyTwhGmt8lhWXOkkMH9bSO4BxcU
MXrYM1X+WzxwSvoczHpaTe17R2MxfCtrLfeUyeYC75rgNfojbEKWI5cudjPY4lVA6j6LqrKxXqye
FAHllfRuFUnt33rac1u1ohv8/+KIeLwPxIZs0ZtzYkLB/NlfKdC5M9LwGrm2eBVWTcE1Z5DhPtvT
X3w2tb5oCPThkkpUAQanrT7GJo8lV6gugt5Uc/tJfHEZO9BYqpHbvWhSbpqkB+7NlvN5sGEazPBJ
RS8sw0JHDy1yBdh7os5cUI7t8FhvPN8O43EzWS8lJl8sJXItSDl3sWgjWBSRJpV9Yt6IoevRROOO
cNrhes9zx0DozUZroeEROBoBGu3j/h0ZdDeOqvqauIvT+usDfnCTx+9J7zpHOy88z/7pLhx6X5Zq
H1O326s8c7V2jXQWYt8h6YJLrmcP3xiOms4d2N6WV1CT+8hFMNjaMJCtjeBit5o2sW9tle4YmHlb
QZVnEPeRHOShR3SOkKh12CWSC2VK52PRDoveDhpVqEIVQC1AqKGjXtmefLeW89R5W1bqZJitA6EZ
YZglrxIZ2/ej+s0BIc5PIvKpu03WimxuxPAuAY21TR0G++ygQTE4JVrq2hm7mSQVzkalR+Zqssvq
AgawDxC3lehReFEQKdYvL03lLkO8pTluxhNhgJPQ2lnJVcs8aUWOTOTXm0cstAAF8NRs674qLild
YE0EnztenB+JYfnnfSRiFEviu/bAlIGaYFIQXA/lJbpEFVun3aoIwKBZ1TPTCACm21DfRyZJaMV6
Y1vPbguwXdAzfo0FRaDkJJBiVAe4P51bacue8/IFtsuC0Q+zrMpAtpVCMKpNnS93+WmhsX0wUVl5
EOSmDdhdMWlECcbd5S7JzPoSKAAy7BJBxQ6e6BubwB/IjCj1aloCezjzfgsmehmiAJftz3B7Gs7N
3EwHo+SGXy5QeEJUpdGUl4n1KX+dVXT1Qg92PALibVLpORY9qsbGoJf2arnLFFtlSj4MiAjutjrb
94IK5M2gt8d4TnN77c6pvUAN9BGxTfmc+QpLaDwQPs9xuI2zj3+JyWLge/wy4FwobExIrp/1Mjr8
gC72mtdA4ioHX6hDi/O8cm3AQFnTS2pQuml+zzzS3cXuvGbHp6AqtikeNkxhlxfaods416AxdvTC
rith292MhonuVpb49M7sLaEMQtjH05hMIzsvLs+m5c9938PmqJZ57ZYgDH1ybJBJ241nCYpBBlV2
sbaPQb2GNKOWLPlgilMJ0aNmaZiGWZx/Uj3kiosbG/z0nJ2DjoqbZtvGJ7gkr2GBkQzNrbWQvE/S
QK41/WukoAwRssOIE+u6oXmtUX+kA/z+1wn/TfBk6xZgi6MvNep+VMOt1UYry85PTHjo/ymUa/Bf
3oaZbjzjpMG6LXoKo2/98PTNYPVzSbVsRk/cz7XMwO4wQtyMVxa++BWI+XbmGEraUueFJEBg0HSP
ttajbag5Ie3gYOBgPoNL37np3m1KfFksZoZ7BcZbeT9flXhKTGIi0MZHEvztorVcpi921/3ur+Mc
qnYOylbjTmBGSnTTNKc+wd8mv2g+Z+RvWA+w3BFIVeYQdFOq3kDUhlo4kRrPJKa6K1THsVsgTZR1
8Z9xvVUWncjqLh37G2vU7K0CXkozuP0aFgoqq3kjj3WNSXYjhaXF9iki4auhfbsJN3o0ieivJflV
aAw+U7cDmX/M/reUA5oIImJvA5QTsqD9kKM9xhkLRpQgfVR/eqdvD1YocxGL5AhVqYzcmI6aTt/h
QTzG2mlUpiUnMVfOx4tWka4twlMm/pYlVGDnfE3JD/ymPlV/I4w3By0PUVDTcEBgRs2GqtLWRw90
m5ycFQlgrJ1Z4wBOqFFsQM3yY3a4/eeGu60MQCGSKQfBQP1IDB5dt2e7VSJt3h5pjvkK9zGMcV1c
yZZ3Dp0rNHdvqdCcAKw/ROHS8ggHOMwYfmnYOyPyjJtdMpUsTuSmOEUTWDPYxtDh9v50gjnc1Yi0
olUhveuGx1XEg17yfwhfazfiEQOeCODksbPDwDDIk01hZU07/oFEt1HiSfJLpUYL2FS723RXVqJE
h7uCyUGild5EM100VvyiKPQULQYghfEDjGggOenbSCdi7fW7jxSmilQ+k4cF9bpG1VbkcBtHiauc
Ar98M8jWAIun5A3rS15GsyHgHQ9gnNys8dpLOEyL8yOksdg6oT9gVLF7pi0rSa4X4dI0bkQo3FwS
w6FrqdlDO6u1tD92LawvEj6glIRHJ71CC8prCKZkZNl9CjQgD+aX5U4eonYNY8dHVrDXxZl6t62L
6Walnt/uGtJKSg2mzPcpvwNwI/1Y/3xXgyGXwn3OEoRYbMTQ4szGYyJEUYGWOw9AU1dd7hRBo1/J
6N4T+k1iSlhT93XdI7qZd055j27+emQy32th3P79UU/OyAchADFTS0EJUvJ/b13c7p3bmRRn/hL2
44Bpu26uZsyWHpUftUZO0YYkHUcsEWH0K178lL8rUjuMBjbNmiiditvi7zXYUIzHpTtVJR4JhIa6
UaZutb6HGGk0K5rFVR/0BTzHNq5AOSLae8xWs0wp9M/1ag/sWypa4dJK5bwq0LOJrwI4K7XDQctF
n7HymSHjOpcNZA/YjlB+X7JHbAt6Up4sNSiNHkZ/1ePaqfwG6b6gc56dLF7ofXoEWUsMP4kUOMAh
BZ3SYP0XWrVmUXRADHJwk4liQi2NFJOTdU72RQAoY2f5VuMG3xzjtgZmDjzmjSiscvCXWRHpFAkj
4vrPpAghkopB/RIbDE425dA6uooAT5VREyftRJVmE8SVL2/gXA5XPtosm3liqM2DcDmEIoEJKjA7
MvHlaOjDYZfrKVKaF1/UwV6SVfaqUW62etDC6VbHgiiOAvvTqREDQpinX1nVMb9kEWuxroyjn+B0
Mt4Y7nKjz+lTjHjjnif1d/bTvNn0f/MQKBFZqNlCK6RgxIkzj+6IuuoYh3SBo8iCEQf+1hm4tird
D5qJVKP1WLKkt0bL4fDcPiB6FX8QZVojRzoAV5d7RX9xGbt5aP3XEvzXnC7RfMXW3AvD0yKL1VF+
HSD3LrvFB+pHFs9/3857C3h2iS056uptyLjOYI8kEXl0+Z/X8zgoZS7UvAFOyRA4Nff3A9BUtZpX
hk2WQn+PP2da9TiKxjK0r0LcfNPObyWjjU35V1AFIXarE93C55GDetynNMTwtEe6TdSXxxaWHzDU
8PNk5CgbcN+l4Kwit21X9gdgjM/zn1WTV9Dh3DvP2GzNz6KBlNi/f+5uZyka1oKt7bggPNzT8FJF
sqvFrI5RnU0fmF5E5cLRV6t8tz1vI2TMyIMfIP5lI0CVYYQ/AIou7iHpumsaTvgK4alZ56BsY6I9
Ev8cQzSdTPdcQcKKIhIU63Lnu7RRaDiiqi81ROKSqqOmjO07XI9XzqHHMNhzv5iqage3PHzAnTaI
z2XUg3TP6bBB/9ShJxKWCYZp3114gx35GZzUxLyjH+10E1FSu4pAx4Y5m04FFurr4AfBgPi+97NB
CdMBpue6LPaRnkGeBm7WOdH6AzkGX1JZqYKqr/H1eCfqkiDnfj2Re3O3lQBPZvuTOpCEURMujUC0
YlaxlLuNYUqz0L4+4Gi3jNkHuFAlw+eqG8aDLurkdXUfssTVSNUTSL+BuKpKm9pb1AKUMlpnO2Pg
zhEsagWIFbO2M1cXv14IiBRbJC3zL3HyVQENHCIfzlmZz0v/DHuzEU1isa8zllS3PsZ67dmPRvk4
2jsUlwMwgYFfViAvC1D7hQCM3U2d76xHV2YJhdaA7c/Yep32mMdAyPfJwBUZNs+BPdJ7UNvdW6UZ
5Ybb2qnxVEaYkDpEupIe+gXFmnJkV0bRUOYz607iPxabSRazkYyZcRUXVeBQTxjfCtRH82aIaEcs
uZVrdECq5sYX8Jn4Ot3RPL/2ukNGHi2dCgHrfbVTiKUeQ/RAmS85Fix0yBPnFg9Cro558Nn67g8P
Pf0lQ6UL27Ystv8oahTtGhTXuH2ucX0u9OK0L7kFJZI22DorpDepxqlM5rQmucMsIs0dhexm4pHR
2y+bKyznxGuFuJLC1i+7pEJC2uZ+oBRd6qQKkVrfIg5d8qQ6rqhhXXcCUJirxfu0ZKM5eHT0iCll
QOyJsn8Sroa0mMsS9rZx5dXDxpDqydir7rT+O+9u7j8uJP4EN/K11zD2CqR3Wynbsz1z1WH2labO
7lIyyEosqxWsCR1hLg0uYn+QFX0q1JZ++2iB762Kx6or9NA3JxBCBl+gyXajQaWCzV572N6+aRea
dvU1PtviZSyTf61ALCHWPXyioVLxOVNgPTVnhMSHeZ30pp71bFbn9YDHTsZwiIoXi2o0yUWKh9IY
AGsma1nHUnj5x8fSOGUpAKSuTxGoVXXgjrdPHyXgcOAxHG0bgQYzgADEjd7Rdmz41CiryfEmJUOe
saxXJWm01cV6Yf2gumDnyaKX6TC7dJCYiaIS6w6DDZbca7mcPCP0Md0JV4dqNhGzaa6YfDMAbzvZ
/qI6A6hjeGylR06roQgnJRFFZOcv+2Imzrs07vAlIxDIVm27ms9MqLtXUsaSPYibrdqq+KZg4T/K
wgQ+HisZZMOrna0EfdJsCglOfg+W5qWxTS7PgPKEVuUq2MwNxGsv8MBQpTQOJRG7yvIOI9vzQq5T
af8xXbSPgEeBm0gquZMFPkZS1FF7MOZRid6WLRkQMvOA3duOq+2Yz0PM+Q6T6atP35Q/82fSKuRc
xRko04qJpyzzkp20wxQEd8PwqLdI2c7As16DmPqVQ6DBFhjuby0ckLF+RfFjN5+x3Qyo5Us7JmUl
nLoqsNEnUf1lCyK/VZw6YCBcv/bWpoG/W59MQK/VTLAQaekvYezmtsGijnFYLP3ZJGHM9LDtJzlL
nZibrmW5rPGNW0j/uDmHV1uvW8aw6FCnZHwHwmCYi3AT7FNX1N4odMDMX024my+9A3wEpyhU7Nv9
dnGDo1ynJxvpmfPP3ZRx4Wngb4sLPm36PB61esdysP+45eHkceY4zqA6rIAqDruFAcLsKXV5GDCR
4/ODDZ4ZTHNO6Cc512IpN+x7KjW/BNynrA7hZhLx7DH/yB4uuKJdRsmZegTSi9Sgm+/sySgrzo66
sLRY0N5OAHIN0wvRt/Ei5wsMo/0H7c6Grp9BA2bEZpRyD8G+dOvRoYLseb7TYBxIOpnM9hywgBQP
jCUgmEfHcqDGiYDQas4wO2A+MK84PKoQZs+iEQ3N3rPJJd5+jgT3aQuhzZWsztxOJuypIzUfDvYq
1M7xIptu8Wcxp6kBHaO619ZtNg0s+MgHUqScvM7CnFCkv/It/OO9eifD47MtA/zI4iwhkECpabww
sg80SoB3pgARMhObZJyI+e+gzmO/JAC/oUMmMy3ysgbMkN69rxRaxltn+YTq3FCCUFxnZalw9Tgz
Wcz1OU9yzD0GJe4dMeYoyCBk30bRAD+2wD5lpEO4enGuatL5SVQd871HvLgRSeLZjP+u7WnWVluY
P+OIdjnNi10LS1zCr+wtZ4uOM3XJlfZh769xF8XhwXC/DlSxgdEciJA/Yl8blAUl3nh+dzxQ5yNC
5NguekMFxSp656iH/Q7iE0hsFQZOTvnHTC+zgacKlFp30a3Axb7UTh7ccPT4EZ5rtRixGtvjjn6Z
iJCXPjUanz4/xnZjDyLYQTVhz/eQwMnlV23vhEUEWjVmahVxe1ytlXywQBwa5MD66Yong0lt9QBe
WBFiGavtxeoA956/LTpFVXaDD5B5UCc4Xb5jaoZOYcmp4y3oRRHQEESvoAgI9Y/cmp3eZH6D3B1r
mET7iVMdCfGFf3+TT3OctTbWwpXv/+uh7MTUKgYomvIMvSpY0bfsfj+Hs1vG7I7C/myHHb6raXzF
hjJsAryZ9FPsbKAnoPtLT1HVnukRsNrDMXAez4tGK/EWTxG3AXIk3xeFx7BoeArfhNU0sUH9qOfl
V4TBeh/ZgcWyyZol5lobkY04ReBhU8B9gcq3uSJgyF2CeOpP1xRoHIsYEZAhCbDnVCKlxEoohblr
GwltJOpGnN7WWAR13/+XuuzzfqBf6zq4U2g9XuXreed8RDTZ+sZlpNKYlZzklIMyY65D0D7YO6aK
reL+dKjvSlmFNSfiuD/ShjvyFupPrXQUij0zcnCXCCl1Hu3ep9ysDHLkWXBAkmt3JxsL2yCdsfqx
LLkHDkDAegH8BE8W0l9gcaqZ6Lw850UaC2rXFFrG6Lo5MbWbFvsK2xn6LsH0GL8gX1P2rOa5EAV5
NFGU6NBs6LG+wtlZz/B0fGvhkx99+tSNDK4YcYOhmUi0vEv9BWrx0rgVKW20sY4ydDpaStipF0je
IxMnONnaB99cqhVDvvESDxlN37OTyS8cq7egFvs0aYMs5oBehsm5+pikflQA6o+CLCPtifZSMIwu
5ads0EM03hjdZjqnQcwULxISzKNxnnpcIPRsh9eOj9xUMaNctOENQgRkwFSGNVHFSKEZCIA+5ODJ
qDmL4QtZF7N1n9cFUcfr4q8CvIctk5Ldurdp6pn4zNDFB3kv0pn8+QR6zPelBtLn0Vyj8oKKvUIZ
nuyzfW0yJolMX5DzYqXHWrvz7soCbSZJ2fSByAB0drjVwfS4lbPJouGKkr6bLppVj7F1hQBmiRmB
Xys+w3YwpzakcRpEpyKFUN+K+/Ec0x6PgwOf5grnLeEOD91nisbl1tDaywe7mzsne2K67U77VC4Q
zwpG7uWlEgiJYiUf2/GjA+0FUbMs6N31WaMNMY49VKQOJhq4HepS0sOWV7znSNdyrtlndZsy3Cre
paRuES73Os6COgbvg9v372Ew9WiUu4RKMaCZLuSwVv5q7beqinpqeWGSFYKGAXcOjrk2v5ZOEFlw
DP9cWuIwc9BKjxOykrPpxCKgwnom3ayenE4qQ6Y89wS42ey4mwX+xpfc0icse+/4uj3TiQH7x4c4
Oaxbc95Whkk6ZC7a1LFkzWld/Esp4f+9lOW56tP9bfTbm8SYVYBZsjK4XalwE+haeuSwfV/aRfsg
KYvBBEXjmAB8LosjpP0uXIBW2y1h3eBQVoRv9dEGPceoxMnsZsNtjt6qs2jqRqgd16d3FUZoslAB
H75eXsfqA8UIFmiiqcGuhRzfHxnr7p3aM/LDylxYH3/osre9Nsk+HGmHIPzpO1ZDpj4VtlvnvurA
xqb+36HPsxxCgpoojguK5Auk7b8i3ENFUNHwQlQIQq7+vuuYciPRsh7KRbUBKomEuyftoSvz+eFM
fH5Ueil3548wt2l+GPsKzh0Qo/HEZZrkGeUc7N/uCx2kntkKMUA6EyB+MLm8jAwWzBcKqfAtiANh
zh5QaL242JeMv0o2GJmJL/lGBcqjywf2RheI3KIckq+d+t7/9P9ue90xVKfVtvufM4AUmLrZSHEC
xaDXgRYT0SydUQNxzAzXp74kSgsUFxrzYK7tigqU/tLLmo7m6Fl8lu1LIjHMeerTr7CVcSKu9n1P
/MHkKzY1/91z9b7EVHemfwYJVta6oe9Pbb6BVhAQnUMfP4OsPggAWy6KwXYznbDZL3jCZo75OwjW
vTVNfQ1UJCDYGqFym1G4fI8wDssSpv5CrXoI9QhaNN/jeUMNpYqpSf9086DXjqmXe4IMA1RhIRSp
VXP3t60nxTdMECxexzwAiD2nQMQMjzXaVNwqekpCARcO/tUrydLha5K86xh7BpB3U+K8OmwXCuGp
j5rzrmEoE1AXaCErFP2yA3M9Tic7Uiu0KzY/fOk5bCBDnLEe1lCrGxA6bq+hIv+iKtgUd+a4gBdo
o23Te+AtuRhm+gM/umpUoWIWFa0Ud9Sv1hRo78TmtrrWVghduGvdgXyWI5JwG/G9iMmIsl0KsHyt
FuXL1M05K/g627btKBTV8Sl0CMWkw9vy42GbLck3IFowDgiPUOHa1p8b/AAGRcJtR/yv1Z6aT7Uc
a8FDYOLs4BK9EaZ0NnfKiLgUW3y9LyT6HtT4CtvxT8Jd3Stzz/mCGphRDEV+YoozDl9bjhgrAUKb
gZDAXEDI/GMOQuvaHq/U6i70Hov0TrGCNyyzp/ZBlDIsUgnjnX8Udt/2llFmzzAazqxCnmtKASBX
0sXBx2NAZmh6aPTgsWxPrlobRiFiydsAHx5GhOeviFTOcUYNV8RYam6EMBc9riwr5UF7gRHQ3jgF
9ma2b5qEl2bCIP3KHeKtgK5ZhUfo0XBQxo62fXfwqMKL1tJN0TfPsstM/xhmc/hyBbUUFuWyVFOZ
l7r3UsER0ZN1QPxkMHSpoO28n0HiUs4uCnUXpk3d5ljBdfu+XYe6PUX5BmKlCYbf3ueQolJK1eMc
ywotodKFyzzR2jWsmMygtvjOYww04fM9Lqz7TGatpeshU+pM6ZW2zjggM3cHZPBjQuAsCpaorfW2
mC1WiEVaM4fLgdfo5mVvjhtp9MZIFUY7+Ex/7XIGLCd/59ADUr+Z2wJ5zHxV7R9dqSIZPwiWKoGu
1ZA48wGkHi+mkzBn4RSpVmzZF+/D4GLH1vglVdmhejQvFQ333MJlH+6Am8ctsV8/A934xnu4i6xl
FISzOy94whdrsu7pFci5zOJw37+/BtRiO6eEWKMv12bJ4M9kMLYJQogAKKG4k0Rb6gZihcFKWDHi
vjNBWAStYsYo4RW92Q0WlJz/8gB85Ml4gbypfrIMPNUNrGn/Gd6gwINEGQ7iKl47Y+5XJNTmAJah
ILWB/Oqt+npG1K7r3muqW9ORtVvlNLlKESPp34T995yeX+DhJVIv7QlICKVagzxgWTnavGgxquaQ
Ba8m29vD3cOMKJoLkhnSX6kYU3d22/OTufd0wKcAqAhZdc2pG/H7IITWap870GifKoXdrhWrAb+f
6v0Vf7NQYc3RtDE4mhZBz/lEI6eQO3+G0f25CEFw0Fcymxh2hZXSFhYcKTRwaqTpOamMh+lCpFeH
rBbox1q58PDsQ4q05SGgsHAOHtUXHborv09kQnmSqXZ3m4+pt/Rbmp6Ljfw2NUD/FbxyGiqx+WaW
A+mK2FhM+OrbUoRIvsJhVLaO6AqUOCswz5o/8fwDhUY6K0l0/o1SzWuU0Xy8bsTmPD91g8yRi+Br
dlxBVrTg3xw+/vorWwmSufBzPvYyg07GMmpoTO7eDzF/VTktJwbPwBGvOouXPKwF3v/AMqqt8Uj8
JES//h93QUMsXvLykmyLsuGoOZErbnnG0EjCangCo5KoqBf4p+EQ9lF6iZPAmxABhZfIXdMLPntq
GtQ5mQubJArkaO7LS1TueO3/K/RMGOtZ3DzSw0yXavK57Cu049fmS/E1XDvHC6QcALLvqnsVqUOO
PGiryl4+v04gq0FMr9Ifl8hnF3WMKaLJTlE1x7TCvzcPn7qBi9uH8iaLfO731xmN5CovzTRsM2WE
yOBda28umdPeH54iAP3ZbugI+3Czo/WIGMKeuGIf194lBYoLf937b/ima9f6v+HbGv8EFEWms2Ri
3STWWHOc/ExITDOMCzkDxK/bh1H38/JdIsyjkWxAS0defMNLFj/YWlxK0PVhC/rYwtyzuK4krtpg
jKJw14IBPtSjPQjmB4Z9NIZtiFp5jmVP+ns4KgDorNdv49Us0w6kgEA1rmEm8HEID9eaEnA0EU5u
o27oL8vqzirrUntLqyjcp8mtvDCaMbyRVPRd30OsrkanTX3WrNMCdilsEk7O81ZnfS9SyGh8WTFv
i7DOZB7g0jk2i6FmBfLXS9R71f0fYCnXSvq2cHiV9fLTcTnIY7b3UWyR3XYQh5AwAKlBWc6P4YlG
jjUMUWSGvAMkU5NVw5wvudKzYaqXBOakwxjnF8qEt4ebnggcU+S8nYp+U+cjQ7WV0za73mkAkszR
FckHlAJwkfgjVKVRsCM4b3CAsNcEKabcMAlnFYxbGCqEEixp2aq0iqya97kRuMbdxaU1wjqyzcI8
+ueCJoaUFU8PX56LZUrPGQ8TFC2S0AFqez0+X61J1t+3jfyMh9Eb7ff6JOxDVjucbxYZWe7y3oQv
cuQoqE/9CVP77QSMzEkGoxgGQxu0O0oZS7c6Kbvv09d0U/7Lt9VJLkON2MlMZewD/QnalX48Gh/m
WnnDPBhxsCBw2eIqDEdKMD1YJXIPbD/VApqQfzDRgrtjITNN6hhu4uc8TOVtWN4Gohu/FceDfQVv
ydVNC47Dqh5i5GknHe2Yore8hn7Hd2M/aaNuryI7g3sMgvdofIFbISC7Yi4qocSJtQtcB17Z77Ga
MVHtCYoCrgQW1XC55HAU7X4gbLSS/quqpDZBQk2i8Btp/1PzRAa0m9Qx1R2pZ92jF12VnA0av4yV
rZxnSRip5LUi6V0A+l74uxxtIVSMUF4c8Rv0CQtGn8ixSYrn5kPof4FQp3iG3rDVomraBnvsW9Df
p9Y3lZ2h8TPhoMEqS9LAsV82ZgSALX7KQ68kmymDIeo2Ivm13AHt5bJ1wN2jWUpOIXF/KUgbkqN1
jPAcoUW8QXNEeH2cFusd5PaeuyTiHYk3fu9fHSCWWD+HPtRAvci/x0fkkW5D01Qb1jlbcm53nPfU
Rva9rYD3WcP3QMi+RB7H8LfNL7AUumWKnEhyPgLM+8byoPeLoDsqExdfiEWz1vuqjMaWzU4+cvAj
BfTvWlmO9ZxEzwN9AgVslgGMTaGGUuteoHPMuONV/pSFrFQTdaJt/6OMNa0ejB4Tv0VBuRJQ04EY
icjQgG7iOBZpoygPew73s89P9nIT3Dz0eVgmhuMz5p9inwkI+kp4bu6bdjEDmA8nglX1PultfXUt
+dV5vI1TB8zP0Z+0TXsNcPAaE846d8T8wtjkgfVxGSAWwVNl/5h9CW5kHqM2ZQLo3r+6IsKP6zch
CM+6h7ZwEis240ZNXq3XDtdMiefHn7B/vtUUsxox29wF5sXTuJf3v+ybxk2ZNreP/WogtZpzMig8
2C5fhc6ePVx+wfzvKokNuxpo35qoZxKl0H10hU77PnZxzTw7tpOAEsTv4H/AcRA3uwVcsZiYW/dS
9GLTalLwpS1oqcxVJzJYZ7IqcMkaudjlAJ/eVUVxLIs2etdjbicvv5sUc0jr3PrWBQYn+r5Q7gdt
eke+q8UeR/ft3vSsGUn20rZZqxMBy0RmeWt6ZXOAh79RJImdQeHq8TpQa170blFEWJWWglPm0u/q
YJd48zSKcxEil9srxDNvC5a0/VEitDCB+EQTIogKD9j7L7KgoHo+1hvGjS0BnZ+wW1ddS8niRNwi
Uw7WLGJ7zvDPhV/H/c9rxFzLJgZWYR/k9pRqgox3i3/XoJxt1jO8ryAPMkm4DpXQURrlMFA6p0oX
JmrkybCXYCCt0DFy/QfCBIaXbQG8b6EOrOMRKbE4dXNQeq0//vUrvzp2T1c8BtXpJ5BZY7zBDT08
5jZz+CsMZjqI2aW5wkvNjLvNvuND3gkZyjG7W5YBV8UE417cJZVhyprDIe+56rHO02qdniA4hTCw
C/03RN7Ve0gdJrDeyPXkXYcD8HEsqArCu3GQQmwvyOmJ1ohQqD7uAZTz+I2YoD6zLSHVG+IfCBwz
Q7dA0aDc9+5fTCEUUEYzkrhVjuD9efxOsTD+dlJ2dd6QHOXdlfNRRg2kJCeouiuJzmhpy/WXNwlQ
w0fI7632MLT/JPKX8XmF8fZ8NfrYmnjceT5xqaJwU26AF0iyeQMYdYWb6lBo8uEpNwl52wy8xMat
EDaLcj5ThmDszkd+qtJJOMjxJU6ScdE8Wsq7uPb2iP3NsPeKG0vp9eSip5hP/VAk+GrZ16qhblV0
PhVlW7f+8kPIPmSiQ3KBBDLmf1lqWzpjuKWKSamehIOT5HSDcgWa3vfhwKZMLXOQfLzN0EvESA+A
MHE6PJ38QFWK+3/++6IOOdiurNEl/Krn283blNl6h4ij4dFJJLONVizDoxofbe4MhPbLlj6BhsGX
0XNMMy8DI4NH348xk6Fh0RB0np9/1bhg6+qfhuZOk5UAHmqLzFtXb6SzXcxUh87Xt4uaOosZsr70
AOnEhnqQfGOtl/PT7zKH9WSBcTFnYN4PLbqZoBeQAjYYEqNE891D+CVfohsTsWf1HVVp9vPFJbcw
3eSKAOeD1SpJS4bPCCosQ8HgdrZJcyVHf9n5tDX6FroTiCbaI/v28X+wOoMF7xEnl1985VkjrJ2B
4TcJMrP/mtSop3S/uRuXS2AB2qf7fF/Qs+OH37AlPwKT5egLh+EbOLZJ2Dz0RCyIBzl37rotx4Zf
1RqZqGpeFdHbOv6QXlKqn9TT9XGs4q7Vp0tFjGduQt8SnTY0F76MqUKvqD5klFB0X61XiATrOBIJ
egJG7TCPwl+tQOjemHcjLbutI3+eOf3RhnOSvby9+oBwBKCAvmNnuuQ8lIF2T9t4SsThPChVNn5G
95evKyaQdSUilTcQs1Du5avTmIV5MKydww4JWH8+JEhXOfv0TZ/8468Z2eZeN5FYmXJtIkt2VbHT
8ugoKkqb6USpMka2rLsTIYNtspQQps9ZXaAiMpFHU+R4uCGPLyJJd1dsuEGRsozirmeplRdf+Q4U
p7gMbyPKiQelNTRTZrWIMpuTRqmsB64aYoGzNLVmRdgsipOmQshxJ7PQP6xA+gj1QF66mVXz+H5g
xoKy4P4CftK9pDbIx5epD/u8LOzW0OzCWtW246BKe1fRfLOcpdfo8DVhlWMnDfn4W00nLlgpfLSK
dI5uvXEKH997DaHzpJVGYlKdRWja5NEn351NionXtjuj6dkKQoieUxlMfFlLcZnHdxU2NphcwynV
FHDHLHPts1ShvEL9+HIx8d9eQew2UM/Scz9yxyRNSzYn6k+ejd/IqFWDgYpKxhpd0gq1DxqwZDm6
YatMa6iRRUCQZfvXse6dUH+E4xN6ywCS+uodk6qtc2xRiJCKrNy5mIqd9iuZDOSEyWOgg7p+RtIo
7xYYuGyV+paaoBnEt7rp8bOtWH2em0OVLp0IHDHXt8X+6xAMYi5YWiYd+Vykh3vKowD3Ybyxpd8i
Z/GVtA0036nsj6Ye+xEonwZZmDtCQSlyGDvaWWWOVC/UzYHnB8x+9Nm+1ti3PE0jXECQadP4FVcr
k0soUhHoNeeZLR6fDeOr4gVz0dE6Z49YZ0vFFb+4BgAm+cMumWFbVFx7DH/Mof8wa3K0iXmqBj7M
35AzX6wdwFpwa3SiZ5lx6UEHdvbozCJ9CA9XEG0HjMiiIicl7wXVgpvFKwtKPMYMF5xbZ7R0vgO/
MZAWwgcb/QhhagNaIR0JYkcQPUROtR40RHmpV6EfuxJFn3O1xEgXIY4r1qbKkt1C+1LUPcKompTh
GS0omF8Dge/XT9NzrdMnAljCrAdXMDhg/ZvcMxFgp9MAdquTp8mIQq5v7zqcqBxT6Rgx2+Nws+W3
JXUCEtfy+MKIzhTGovXHzE2qUeZP1DgNbePtJzdCIEWNNZ7mF5HbWzWIdVbH04CbpxCbCa5xxlXs
YynkCY0tShmWhFMeyYA2O1G4457hiqmEnwQ+he65jvNOfRqNHww6PjsUvZYOK+R93XXXHQMAC6WR
i2amlBcgIkVYgpgmBN+aAQoWVBtDBB1W11xu1rL2a6OPB20vlYiFBwEcymLs1USlEEZt90+GrS7d
gg8BbrbEf8tme9AfNOGkO5SBMyBitdpJCwOkT9CaO+RFl3R9pH99pan4dGk76FlLX+pzszYvmBx1
FiGbOfdjqIPT3EdnJ07fUq3aHAJh5/+2KQiXk2R0gcV/QHoaNBepmxqKf6xd4QppW+FwQ2xOaFPX
A+0wamt4r8Cr6rWubgltOcAp3UYZEPbliu9sjrg51gaXe45cZLdcFxmqfHEAnto5WOeZ3ODzMV84
Z/nIyyLaLNmmW5iMSYnMRiXjJuvwSY18/+ApWWsxf7/L0y9yrrebNIsun4bdtBlbRypHGu72CSUq
Xo/hP4uPXuX3b9ZyhLh9GY34xdue2aE479EKP8VHukdqGw/vMCoFkke2o4c15nEED2PTyjNkwtaz
sE8uXGmPk0SKxMtCDef41EnNyuV8QmJGXYuKBaJbBjIWNTQPOy18mexgBBeO8mxVxECYDDqaf2UZ
PMz/w3WjeDPkJyYF7pqFjqdPaTEF43SevPDz2KKiwDPXgfpvDSHBc92JjgvPwalD9qSBxUxqEQXB
vo+r2yuHdTIkOqaa2CAOfrnQCagZHRDL529VYS+fIBVAK3wNP7SA+mLB+mYULhCXoj2myB+JQwWa
JtLvCFswHmGzfyB13zZBKJCiGNtFMjLJGzjPV+3XB/U8ZedQTh1dNCFCXaHLt4G+cr3wgFEf/sVD
LSc5zEWDCbOtcmpvWu2888NgnLpYeZ/winE6Ae2UWT9zAYyRmPmo8jOpO7HBO1YwHxk8xrQ8SIyS
zGW1gjLPqhKWv7otR9ZGoBvlhQ/lZtlEnPmWVqvT5Pt2CoNjwA8Zo7U83go1Wxt9m86nTKFJqo3U
/A0HwY3Ufd/2URrgHt/ny+9DmPNrb88SFub2nCiqZxfhzpCe8SVZG2duO2Z4eUyKnNxxZKspWvLd
qO10uaIQu1FWA7WnlQUT7cULaZkIj9vQrIdAr79R32rMBGjK8eczAfQAkxgL7nrM17ufX6EWfpa9
PqDpUt3+8Dz63AdrsIzUWUPxfHK/miPbp7ERDt7DRwC5Fc7tdM2d262mw3dK8R0kLgSBcQ2pajpT
xvPEtpUxNJJPOpfZFmfs0qJf4go3FsaY2XFtbxXmq7yCUEhJ0u2cnlaYt/SUWSulLfezQ8K5dOK5
qYqfBzRWoILs4q+MMLcOzxugH48CRNhZxykqwPs5uGf/zaREai7/1ZjH3CRwwSSV/2mmwawYySp3
mGBv6g556zhyBpqORrMxM4sMxynwJqNEfTui1zwmqV73nz81A7cDK48uWJ6R/ylECPHcr7Pa1l/r
haqTsSLl2MQuNdm5pHrveJ70Wr5DGUQGyIG9msKCBtWLr3aB348i3CyQpp7DQQVbW/B4Y4mwPUk/
8jAKT/RBrg1nbrk7zXGEiy+6Du4Vn4/1e8UOasg+pEikqyBc76LCq4cHI9zsKwG/YwhnmOKiMst6
675SlOjGSz+zRkSMONBHXqZS1TcTA8vgbQ25PABl+x7BplcSJfyoS9EhAlTvlNfe/vA4KzL9FtPA
yapjQfEalJ/0/S0Z2egMKn+QlmRCiFMXNmt6rw0pFqHyyIGtsDFki7ln/Sp8EI5KseLBEjyWnzvU
YuM4p2fkOo8xtqf4JpXKdFIid+toFDPHCJvCKoPf1gvitqkIJY5y11XmyTVNno0D0/0R3NVbi4UI
WHkPYtPc8svbG34bJ9POH6ahijci7Q3V0DJ682jBq28YGs++BOdRacj4DzSxtdc2JieTs1tIB787
M7dnjA94NNsaT69OC3NvyLAYE1VsJEjz7Dtz60Dq8sAyKqAK5KvmkRJUkbL2BqNbMsiPxY+5zav9
n05dSxKP5B5+IkJFJrRjYR4H5/yQcXpxtpI3oUKypoKRoIVmWhDRjhCaMphiDgU6XYZNFRzaNe0V
UPiUpO1MUKyR2A4dFrKk0jNzB+Y3MaePNSF+GfjBfHTQXXCb6iHCd3xxqibtL0uh1xQPqBorEzRf
P/pHvElCf1mGoEwtweZ7Hken9WvszKWDFsRkFXfNgpXQCflun/hHXUC/741zmDqdLR1tp4wEq3BD
fUkxYOFlh2d1ytWZTsO9P8x6Xq7/JuZ186bkttUo1oYTytuaGW6WQqcy3jZnO4rwpURSu5p1Wge6
fusSMyoe8ChaMeAKfywwp2+RFfZUkb/xfrWWMTzMUJEb/u0FjrLUaKCei2I5GJnrGkHmlyKN3Yev
tEivIfOZyJv4QYLtiu/lsNgdjt+D/K18rX2SA9MlhdEb3hdpvIgthyNV3wDazGs/Q91g5YkH6Nk1
205CoUoGwPgxA8Z7JI19LrLSW6PFoTq2zg/GhWOHiWlJszRxX1cq2NgZTZlvISAPXMzIG1VzDZlq
O9ZNIoHbkzDNNKuUh3gOK12atXomPGTlx58FrifJNTCO3/emGmyvK6K5FKdA58CAPkYz+quawBpW
cJ/r/67ObOEtPy47aoHC8v2OP82BrA/kaP3ssFllPDGyEcUQ9rb0LPSvoPntwLJAJQf6xEssa583
XvkCoiBWCDp5LO/cu6quJ/UbimWIiD+o6O8gGWQR7P7UXE1Sn2c/BhCBNhO9tKUZ4HaKg9jsdbp4
KNr6ZyzGtdXuO+1OnWTgDLI631UTqcvCxt2jZL6wy7DzgqGh3xfN7AuD/W8YFGEqsrJ9s+0O3gYw
jjyfyFIBIOat36meEwh+aHt158MKo34CQTRIjkpGGcRDAqGqYzfEZo68PXYLDBYEUJNfE7ruBTqU
bsHtt0TWLoUwMkHD+CrWThnz2/+jKFfAva4B/0Zu1GerHdmEvvHt+v7GX9TBfQh/tRQ+zUEJzkME
IZREEN1q0FRUWeU3MkpNQ8tgsX1rpkP+v3PM8fGh9RKAV65GsJvco/+im8oTUALgkiVcqKHL5u0j
iXw3QVuqcsDS4Eawsr7nDsj3bR/3Q6U8SYqne8ehgCpko+NlJUBInBooeror8JlwnF6vgdw5IY2w
hO8UWv4Febxoku5nAYLQvTmcFpO2eWNwYzAvRkk1EMQhIu3tjROdUNvcS6CZcoFUvpCoawU10rxe
ykVUg/pQzsO5HpRPUUXM8Wpn9iKv5vSXQ0pAwv6R/i56uw7UotoD0Igs24eE/OeoM7GRdWuWhn0i
LnrDxDdbf7KiDGVQLFJeyi6dkm3Mi+KxdzwchWspZwV6yTo6zwC+Qgeiy/yOh2ptsGPSKXQxcVJZ
5bsGkvF7D4M5/l9Gsd8ND9CAWU8orhmaCp60gFhXlkveNjWOWmBnWsgvdCERHZLSLfdI6PqaFIDG
c0jqDOvwZAC5T8ks7KRSGa8MNxJI02IkOqm2x6tt10HmnucI1tl6DxzMraQSYpoFFjotGbQIIDrp
9uv1Psf8w1L9YrV4wwwvY/M6BCmHoWB0/L5VbwVcLyS6wNqhmxVHCuzTS78HAiw6ZOdIva9vcphA
riFjiEqeV4UNgt3OKEG1RUP7gB1qjfg9q3cKXZnExqRAplyZtxNZ2UQxHVgHg2d7bGvK8CrFvZer
+6yEnPHQ2O0UUIp1BRnLvaOdjs6viPR/vMTNUh7KadmMiLBjYlZEL9ysMcmiRQDmZ0ct9+Y8OJfb
qt8VfGMXRFsYXtJmcCuY4wBeGKq0AQEubOt+nd3XJJO/GjNpknqVbV479CQ9rUV4Si9tGjoBwkdH
0gcKD2ouNu06ZjD9wLPHpDALGyhm0Myb4RnVtWiI90Xez5dGPBWCyfAVzuslEGVrF4vhR9RWwiLb
i7ii1jMPLGE6pHFcMbyOy1Ym6dGZjBnaVQUn9vajqWjNCZHeZHNbXC3uL1YHD8d9g1thHWaninWM
yW7ywRODQ7Snlxhzj2juIhMWnO6/SwGg7f+rdJwl833jM6M4T1ZtNvP2B2NW3ZErfDEmkw6TngZf
xuVLIZoiOy4xu4xJkWM1fGY14SM+OR7iL4g4JWffE60Z5jNj3yqaI4fAke2tmhYPHNaurH/UwG5x
jxzY317wWAaEGPG4r1daJHT+4TaXuK2EpYHR4OIhsBHuHQCJcAkda69EWt/Y9vsIZliMCT9hpLap
MkPFsWmRPnIbWQzk/5JuEL6sSn8ytwkWNC1BRtxBKMUVcrgdRjRJ9ttvXxcKCkYSf6PWGtFqZMMu
ReQLzsh/rInIuT0/nJi7kmyupKXtdKTIVf66XElbxf4vj/ZqHyYmUXOmY1o77Sq4FfhhNpKhMB5e
GYsKyq8x2yyYzA7D/TrcxfOpZvGQq0jX9MncKUCVJ+EK3rGU4QXYqEDSGXcGDoIgiVBuhS4193Zn
t/P++EC/zusR7uMBnT6m5PU/HQdvz4eS1LVng7yIUPOmr+TbHesN5fKYcbaxXdqNahP1MMXwzpTA
9KaXCuPHhwHKmZIMMQV0SADtc7ILEv8Pg42sTCRG8C5vPiQj/5cgVv2KB4WXTD578yG/A9V+zEOI
Eh8Cf9s8S2fMK4LRnyhnQw8jCRCQR+dbLFfUCj92nCItBvXXowb5b01lwxhozaupXVHrzo/5Jp98
m5oJNMXQvJ2PzMz5O6Lt6DBBdvooaHf9f9B3P5GBhhWIHFVMZi3PvGNBbda/aDtRvlVhq4DKZ2sx
Eo6wVje9FeiS8hAit6jbw56xLdRm2nisYYx/vB9ZD5TnBxVnFL/T/CCwfF0SMKjtn+91qb32mONh
zFkzwzpTv0gkHsmbh4r2tAP7iveZSWKN2mfuABC8RXYlTuBhUh8lsedbpf5Pl3a3bCnbyPz+qO5e
I3J7gijtbomDxO3op56T5NP/XAQ3/uVDP3ADwHov65EwIAsGt7ETjMKMIGN3uGWhfTEqWB8YtJZE
zPYCgmx+488G8O6pK3TZ0w4kPSdAH7CiwwpwVMkcZjO6JtOwP845j0JHu9XgRFzY87688a3UkMlW
AqRZbzEiSITM/t9KXfFRRKXg9iEtRDI+OtSbwDqZsEesxU9Yo4tLs4mWDJABZqURhcwA0Xv9XSbp
iMwuf7CmmEiFEdrmfXIXfYOHjXDpL82kFVxqefXJ3HvJ03jtiA6A+GCRcr5Ic4zcEhtd+3Uqp3b/
MFYzk1ejiExB5GqWlwO1W4RbsrHTJ647Z9Ms9dr8UQ/zwUMIcrzH/IeUd5wDBt3bI5erLXOFHdgN
FG7wnsJ7yy+NEFRL0EUJGLETzeVyrpEHR4VdhvEPz5N8oUwUEgPaUfLZus4vfpRS3vSABam01Iva
2KzaKvOmdQtn/W7Fk8OB1vqQO1Ik6SVxCBoII9pw91ZCS0viHivoCQ4q07LN500zkGTLezz4QWq8
zQ2UcFxe1++eGNLYj74HiNIdFWGliY80s6H5NZkeb/CJw8vc+vCnWUWJtdMm3c3EWAnrDUaKReiO
4f0uV0E/WglTUGr9L/RPCqGAUxjFjEC2XoyQvcNSC8+7U7DgEqcRlgam2TLPFPzqjCInr8X8IL5O
OAcM+4AuGsj9qo11GZgs1lsDVgwMs7N3DrCDHMiwfponfcmEGm1qXJDh4aGWXtuoUYJSuS/rRwkh
HuE+z0Hy6EwbDNuLBR96jOp+Lfey1r/FeDoI9V6r01AmAZz7f6ep1WnctETmsEoa03n0MeHOnxhk
rVa7aBNGuYuNBtVYHEn2Ei8LuWdOkwi+5W9DjNgHiKaqVl5/M9QuDH09XerJYWmh3EYz5QID3xwU
1uIVB29oICEzMP0JO7dWAMmw26nsYfOc0XLY0MGNb2Tl2KtwD3KsluPiBV8nSbFYDJAQZd3uDAd7
NqKVUJARJ9qYQ/YjNO4uLMx7XN/dwVsajAWqRXVDUMsyYoYYo/Zd2XxKd919cFt9u6R9Nh7W+aoV
mSJkz5GsNMoo2Psf/iZDmsgdFmE5R9VDqde78ITNK9BDlIw5FDcseJIYelvTwz8+WHKmdIZfSDS5
ARGj0o2eGhRYhCmUGkGI7fbv9MJliUmacss87cb8PAtfLwZfK3KsfdgXITU5G65Om5aH7g+VF/Ex
/ZvKqbBbcgP5baccYHmsqw37FzPv7Nx7WgcBu4aehT/pHtkvP5kSWmnH3HYdU71uWvBsRvFDNpVC
X6JyyTUz9nv+uy0D+x3x1hYdpfUFlWrAFimar3qwXOy2yB5B527C8auVY/QNUvr2buEcTffKKs90
q3wvmVyf4qmQHGtB+y5EnXFZbwtBAKs5PVYJIhbV6K50coxoV76YaJJqfeV+wMysXx+VQkt0sS79
42MT6ZmAfHb94BoeVnkjKtWSFT1VgPb86NQI+MAzCeyVzQAYtevWHWiPWMJfxMdx2KrDPrDnbsmP
LMUnFOnXWxeo7xbL/7vb1x7yjS9PVVrYw8PiP7bYIf1f2kLRADEBN3c6t+ab98mhMmR+kYbYb2WB
pfMs4nMbZiPJmwQdnrwtcWzImoRqUWWqfHwx8opfB6CXrgRe0Arh/GyECv0+hHLMSVzk6uGMdiJA
FJLQEUcjwTh8i+n35M0gq98NbvUxB3LoTATMSfRIw+F+ik4xoZUOJF3LJVfIzHtIf5Gmp4vPJuHv
u3BqtkjKE32bjTdlUIkPDdyoOnVfNwTetlO0P+Vs5+TOSffR9iHoWNFIB4BBY8szyWnbTS3TnjTb
yT/j14gdi6LKBS3i4dLJiIZMLyz21r6cLHdwP+VWkQSE1gD7ILSJQUGYhpQVDiTiGcUVCM66+zld
5UIeRawil8//cHXtrF0Krym1kKmSDPt8swrlxT/OdrqbboiVMjbDo1lM5r/ZHWJIZahKbTD4e8QS
nWp7e3nRf51e3FfeeIADspjhWmhEjn/tUz+V2jF6ZbXWg+3raO28vW1h/W9PPMG3u4xJAnFnYkQT
fHXs5e0vwboM/JUTLL/oDnk37HoO2nwFe1CGA5BnLA6MMaUGDQl3M4aqltC84BEyZSTNx3BzLcXk
odlmKf57LQo7HMmPv2nXg+P51BXeFkp/MHScBMj81d85EIEPB7spXLU3odqs9Ine/5FvoMV2/Zuo
D/u7xaZ/ZGN+jrbG5DXWYAPyvQyArOeC9zVVx/AfOCxl1o0xEwgozoAraSwJCTVrGatb4dB44OMy
T/q5X94fzDW0vpEmcoGvdgVJiRxNCDb0wSReFnQh18r8vpAg5J75fAcyKAeVhGqgydjb451ra6Jf
sNv5AqH2Q3BSsexPA76G1/hvMjwhgQgfdrPLl/tfIa4SxQiXdkjUNp4dgoGzN+3edsECayI6VD9C
whAhlJHzVLf8lLGAFT3yRMBEUBErOZYVjbltbr7aAhYGKhKr/WVqx3bAZhN9WukqC9AD0Gv3mi83
/F0uBz7i8u9Bi3Q9v5mo1JnSk21wW8IiKKRAYY/DT3jfMP3kCG3kCVofKsnN+AYMQjAYrdrq1jEn
bATNuayWjKc5oT7N2UfN61EthwVSHPtDN5xDppUyO1DxWzT93Yb6bsIV89c1uiQbDiyqhPNBgnmY
Y1REJRx/uSdh5pjHAEiK5e5qMX/yZ4bJMR5ei4DvNesHodpLY4SJBjxGFh5B50o2pgsY8JvOzCFo
zUfMqBijjUXFm2t1m5twc4HuXvXVBWofsFs3cwiKyPmKgkw7Ksae+95qQIZdcEMJlf1tnHw/UWs3
OnqaSeCyHoWhvutPaMwNPbL0FeXRATHgdcFgEuynWGVeuyhjrUXY90N9HxKxWkJMoxrUHGTSZV7D
JqBZe0xEuSFOrAHuUhueNkKDW0fTtt+CdVCoGuR/4N2Pwbv4/iTTPN/MgobR32pV495kX3uyHdQQ
7GuSnk0GXPDfnVEWjpE6GzY37k7ZHBMxb726uCpepD6c3x7OajlGcLpfqr90H5p7blZ9t0BMouEj
5bgiWhVUSYMs/eQP9wgBVUc/CtiDXD/Xhl0aUxfJbwp4tfGwrXwSyRpxyK1SHMy9KckAsxjzl2DC
iHUd0wgkorLknC+L67GBgao+/CtFs+916p1VEXgy77T2H90ZKGaDvzdWw6kRMQrK0KaLihwoEdC9
T1suVYNEVIGSgiyYQTzQ/Y7uMy+/LJ4d/IELdz3HxWZuwfoKFv4Xuxirlv2RVrCaskwCvkrZjkCV
Ps7hdLCtg1keB9Ih7IADjyKScMiAEvLf12Lk9mxe7g66f0n6bI2KRPTrz63UH0n9ULMc97SEmhnY
YwIrhlDb/HgJ4m5flqunFfxgYSHtmoc9ZArUIJnGvvhttVT9hdQwUZJzeCjx6luFr6GSKIDEX/xp
ufHWmWSNnOhr9B4Q/0k23LMN+f+xX2FzhablTaHt8U1GHK7OL3ZOBvuS0DvuDdi4L0zKmj4b20Ej
HgMrn6Bk7w+IITu7LUU8PAYCav9pRktxVfe80jrTZbG6DgRQOtUjEggWzKxsUFNv2kC/ep3RRV9N
FOgof2bqCD6UokmnvGyZwXiXTr1A1f88hVHHmYT8RjjNIUYZjgT7saO/dTqgp5HSo9RuqCkEASfk
PUjvy51TsohgAH78MnufRcPQOe4U1aZPDBGGqmdfTLtPgpps94Lfk8W2S5OwoSKTcgiMP3drZ07W
sMdDYisIv+jMO7d9UP+PrMnMfgJTEZb0hYrfE57s8Rt4hKwfmvOKG84F8AA5BqsVCJkulBVD0D13
HISwvilsfntLfIPTCnH5FCm8pgQSuv/UeL+/ELJ2xCejbPHs8yIn8OWLdXqc2e/Bp44NIdOpVXb0
wl049JdbDTQk4LjJJV0XRIXe3M1FKxxjA6cxL4iwh84dYhJtxVG1sSIaxcGGvHPcuFxoZi33W097
EP6QRhPkGuQ6htNl8x0DV39N2rFfczZk8QrFvV61ruY8+r+c4d77C3qY2o6SoE1ht+2KOxNOYQ55
rqOpoMeNnDOTv1kUGKEjOKR+85QnKdOoakTWRP/iAJfzVEiZSxwjPweJ190x4rdq1eYsRGRphJxu
ea7LhI9tx3CHrX3eqhOuDbcuo9g0m33hzBTWIQ1eP8gdDBtUoBu4lay6e/BHdxctw78tNg2A2/aW
ugPOmu7LSE2sq5LSvqkagXOvXO5/9WspEaDBKfbBrgwZbm+AgYS1tXf3RUmGXZxFw3jzN3V+5yiQ
+UiPfzX/61IZmsdVRU9EMdIN0epr+vBYtvZiHjgnsigzy9E3+g8VWJnpaKk4llxqo1bubx9ndnCT
yEJgW66fBgQANHQiRw4lyEquGei8iLarlf6bQ2kfvrBmroYjL0SG2lZAfEMySbeEsObA4FtDxc0w
rJKdTf1WZw/SB/CZcC7o6o53vNAhoAtOPBxltrKs/N1787lIC4rXyBBIvMp5M1D0HTfq29dxrbZe
TjE+u6i1VQvNJujAwoq2FAA0PE8p+aPZcQ7RkMrlD/tku6o1EWSt9WWIgMBDwgcaWgO1Uw4bJ8dC
flbculdChKNxlWcmpgQRU/GoTBfHvWXp9LxWcYiZXC6cOLfXPmcWiU66Wb+lB6sSepT4BsvI8kHC
gxHM/V73SaqJx877tVkqY7qQ/Gj/p30JnPO2jJZakzwiTnoFjCL7BXLtri7qONd1oA5kk6iPuMyi
pSU7KY47YYhZkJYPbpNjGhW/28yCjmo7P8z278T4tdXwfdzMjcmg6r6Tf3kFHNwBe5qC4nbTkmqb
HD0upiYgnZPL4ciN3puFqpFKXvons5E7GT5lO8u6GDm1geOdNEQAnLricODpV4lp6nJt7sDSA1Gi
CfcMD4WPf/ztIJzym2jx/CvJWYP/qpELZvar6b2xhIoRgxtwOna2WtGZthREe9wsK3SgWJ7wD82S
hVcfkvmoJ8ygmJ+r9xqlVQSooeEQcavEdMXoXhG/IbRtbClpBNw7iFWyez+KgJX8g4P3tRgMfVxh
EDx4cEN425qYmax6mOwO2iKtvLXjjMk68Lj6FUde/oJfRcVlJkGx0OXSkH/EJ+dgn1ZdYNW4vOIp
xraeqaGDqypoYBtkZGg66YrUy7xzHTeKnYsH1cA5l5+xrRd6jJPbBomOzXppV5OK8dA6tZzzyzz3
LuQ3NnnVduBYBZ9YiiOsYmZVkQ3AykXEgzGjc4A6n1YuwaDSYCGQCbyMMQQxufnIxhg5WJrLRd30
wscOdYLBOTABhA/IV+F0VOgi0ipeAEMrMDAlEJVknLu+mJ7d/KsrXRsza6lzA+Du7sUoAG6I4l4t
yFIfxL5aGUJ5jMRaxZ5B0NlrzYTL27dw8ff0fptmqOKrzkr1yjfi8VHaC+202G5yDlKIvxndZ0C1
palkkQ/BGl9Wxp0dEmtci55op92OxAjg/G0x8YoL54AMSuprGP8Ty3z+F7dJ5x89wTd5r34S80Ij
3KPMBKO65EkavphM8TqIjJiG7bfYrW+ZLe7KwPnnBumEiIJZDH/PDInv1BDA4siabQAwLBxrvZ8i
MM+VchNjx6fK2HLZhbilL6ViLvqkFJo94sgMasNrrIoYaq6jBZQCb6YLn3mNYddJkXeUUMy42nM7
68y4MWFhCkr1nXY7dBPhiEZ01dGJpLLbniUy11N2624sp7msZOeqv0pNSU3cJ7KWz6zNgXuAnqvq
v+oKY4TrDJFVTJlBK2JvXIZOka+W9Cx0pFl6eJDSGQg/3aLK4EmZgNPS1KIH0mVP7BOZMEnj/LfR
zhKUf5n4tN7OHMKnsLi7X7/sVPzW/JIfWvhXr+yxUAeDzQB0Z3bsMzbsJh2y+BC5qhbNuWkSkWS/
lq/3pFI586UQzVEY3jTN51xXSyyr5HDHTeCf7IpGBYGZiBMnuJnnfRWT/1Gr2/Pp1qiwA1r+Z+Gp
cSxoPYImA99PRWxoVbzheMOu044GeQd/4Dvf4CV+oWtBVPHnrWl/wlecp7Kq3KHthl4m7ANkmAuc
t8FvQG9fzL+DRi7LTPLBrRgPS0/dX7gMMMyyZdX9aLuXlRXl5IwDMQPqvd+3nQlQZ80Qc/8rBX7A
hbUAK+xy4H7d1p6buFMPfM4PXDLYFplPbTYd9OI15p3TMeTFtIBpdq/R6hz+qQHjjghk/eK0M6j4
A5LW0O4AYm069vLn2VM4iFqOIJwYqx1oK81v3nRqpDjol3ARCHPVbIph9IkOeGp0PqGNiBE1c5q+
m16M8hr+aacVkMw/X2fl1DhKsnxNklWEj8y2oGyDDRINRTaOFsO04TDqtQIbgmPByLvcyT6TrR3P
xR07S2DkcJP9o12elGar2GGtTMgeQM8FCPeB4eZK0x3z3MiV5c/aOSUtrj6eEcz1mDOcij2tWioK
72OmHQTc/pZFtTWYxpkTXPaxsMSP9QPIej5rpbbrlIsz8YlLWV5a27t6AibKA59SCOqdJZQCvICw
Vqf9tkGO7VAqPfpmXTl8yVFTDTW0eRRPwSUM75jgUZvjdzN6pzC/2sMgtgNE4j5Y33liylXQuYVc
36N2Be35qOwtg6BbjmYIevOg7jWvw4rytYugUElg6CZI8rZu0lSnQRdUOIX8w6wbLbQCJV89XwEE
vKkZB/WKuHA2RYLtHHsDlabMLJYqf3LhFNXk9Ka9Zmjj8/2ZxHA+n141wh76BKt83I8eWWNDOK40
3/CIsErR0RQYO9AGmmj+pltWzjQOPDNzCmXL7ma/oOhKUGWtDg5S03iz465hMH2WqzNPrfc44NZ9
4IDKVg/mtfmHKvu1N3/EuU1peTR6e5vVVq0RhzJhMVyTmevkadM28MnopXQpTr61igPVhTK1pExK
fMysmrIRYGvS5P19lnUfs3KhmLA31lya0Z9o+X+IryPERUJjoYMRl3v8wVHey9xF876FbkvLUAj6
Bb1UC2snq6bRTl/0mxYLPG8Il752h/ukJqJHxUunmGsmn/7UNCQeZZAaSQBp3JdzqJf8J0O7+sJk
q5ObhfHYvET60gtpxdEn2jpDr9e58znxzfqdCWYoOrp2brF9S/LHHTDhsS+GgW4yVEM0ENWw5Fkf
u7bs7oC3ZTrCieSwPsXTzlJPiL+voO+v+vyEORMBtxjGUXQsE5dE/Yo2AUvrWOjPfzayr6W0FijJ
Rz35J6opmAPds3ENOX5xgPvMmSmyK+vU8fJcQ+yelIPVL6Mam8eZDMswB8w77n4h6vdgmcFyNNrS
cWyZKFC0kYMUjW8MOOY14Wavyx22dUTDTI9o7VwTqrpwnWxAkpo3zFrKhf9ptlDbDDc2jJIb970/
O8LTesZaOxTcviMNNqCV7r84iwIWnMA4DQBnJJgTgRw2o5lgXaDfK+WgUYfw+/5xFMto2o8d4NXH
nyM7T5Uhf1VOapNJsBkBjl4WyYozjjpSnTVYKqoFcW3vaFHofZ3/3tTmluh0RBY/AzSLMlTrbbo8
cf7uNhghaZazYt/V60NhbxET6FXA375j1FFLY+Sve5SUk49lyh8Cg+ZmKHYUuqiBtrc2KZKDvmLA
oRFUjsQLeBxY7hOqXbIbG4cSgyKOLyUJVPRjWnTLznA1mzPNJIv1y4k2hyI8YoLS/+ey1iD+KA3Y
TRExnEdr7wRxjHD4RdiTj2r3UW2x9HvofQgnydmw7exECCcleqrYAsIQ9g4zKlidl+YcpIffoPew
o4V68ueJB//DFhTjivOvlJ7HMXga8E/ofeYOWEp08luxikuqLraRWAeQi2RyBzsO2H5FngVp3gRB
2mc8m0Hsx82fHT+3MZz349VLmfqZx8NWgJXrwddDRyZPwg7eDhEqyB5zKNVDB8RmInCKvO/WY6oF
bz52eX8GJcCljncn2g/WQbt14On+OKYxoEc+UCP5GqBuB+HSNFtq48Fe2Z6D+NraiQvdby2bNoaz
uJu9sZDNcshUwJzC/xWzBGDwI9hboU2qkch2v6bIOy0uWKXW6YLxttDVOQ2kDm3lJMzZw/6HdkBR
1M+6CF4lqxcJUzjxsRozOMUJXlDeUzZyuLGP/RrNGhDOR5KPtXG5oC3JVByGJp6pr5DkAx2O01Cc
Mfu5LP2Kkf0dqyMLl1cW6bg8ldBuySSvqvGqy7VGiQ7xVAlx7SWZhpRVq99MptemaioU34Lz64fF
SY/G1EPLaVfPcQ1UA/zwjBSCcVGs4QFKnQTUonRuqcs5rMAzhKDFU+ezVPdsW40/HCj1x7kornL5
fFjY69riX9naaioiG2t7X9mw5Iz3/KV/wcT1Z4cro4vf1Z14VupFsA0H6zedqiAPpiKKEYj+v8Kb
0Ymy2nK83gTI2Ax/4MYNnGeqpaIq1KSzMIM66EDVuWnNdiyhc5M9wzJeQYf52wd6Ekaee03OZiAZ
Twxt6Z2vCBc7zgZUJGuYoG6BE1tCZLLz5GlqbufYrw0dTLF4kQym8ss0R75wPrTe26CRPm7GmHT2
QySiPcaWCgpRQDEyZkQEnHDksDCWhPGADSxIqDZM1n1h+2JsDZ4+Z8BGu2YYZy23WscdcEE6L0E6
qjK3XLGT6Hhniak3RE9KPnEJ10WVNnikL61LIeaLldcwNzn2wcO7AOnOW+aryW0rkmGfET6WM2aS
jOjgTgt/eJ4mnKYsZPDsewYLK8plK19/g6A/mbNXERnpkKwZrYuh/dusYglYh9ce6yMwFuyrJ2X4
XwSA37HoNd4sKWKYDt1NCK1QeC/y8NjJAtJOt2f3LsbZU8KR6OlE/1LiKDVLqlf/r7chRDktKgqF
lXWGhU2PImZRQ7tJUor9KCswW1quyagNaIlztNwTc6j/zQhzd2lWJefb1dv2y4dwNuhR9abm5Kcs
FO53g4K9X8ugixMcGPXyZR4IhSN9s03ZEPzxxjUFlC9pDZvPpSX3WfdRYtJx8vEHTLBVnU4cF75X
nvEC/0sjlxmkkuY7eZtgdBb5N5RuQErFxZiEa9SpHA5CwTKHpnuQEII0iTpuZrycYQ86dIAL3aCF
7M1n6P1TJp6iigm+9Pd+nAyJBAnQ9Q86zO3K65JCxOdXjyfFnscjrWPSVYG1qSu3w5MkmbsTlzjt
orEWQP5LXUSytJ1jIJVmuI3W/5aRLp8UMFYCdqzmb/EfJU4PptnboVYcpE7z0LTjMm1lwS5sYnGd
JbochL1b6otAUI2jZdcRlHEscaCqtCsM2udpZBTp4O2eSIn0FqJ+TriZ8OhqPpx+r3TiMQHhqWtE
NLoWhhbmOaANohL7V2CUnFY42QHUxLUEgaHyP4hjC2LMYTLAihodQpzeSSYXi57Huj92bbI4Kf+j
OLf035x63tWQI3N6YNaRA3wR03CQmW7wLZRu70XfXZHBd1HboRhZhzR5kFbGHKDsjJEBkIrqc4iI
Arleamm79Gh1ePOUOcJEgOGnYShlfzXgZmAi3ygJD1oM36t5yQKHX2SKigg7VlVhEnn8luMLPpMG
u4bhB/2lkIVO52bdE3mvjQpvsL/1UoKy7W2Xi7LsJmIyn18Lv8jDZelwLFL7jlKP/YYRYEOo+sIL
rEThM3etuKbdvLzPT9KpNQLuvRHKCg2LyPg4+7sNAKz9fb++lOPUtBKxBsatm2keuI8JZsLokVQY
joHDmvqy3T1AwB7rxVkkaB+gVrJ/3TP0SLyXBeNv21GFKg2TRbodvUWotFlNBVpZBu9Mt7KDb9XG
3+FLrzie+1EnQkxZLRJhbxvmbKHMO6Nv5qUflfsK+bhdMlRYpIfNF3jl2TVAb+P09k3xO3b/Q9uQ
YFhySSVkefp6vSJaIhkWXncfLkSNfoDzDG1d6HLN8Ba+IIGxsiT3ghTvcGTrGPr4aej8GYIujXqq
SvN+SU6kzZjus2REbL3xNXnTBOIS99hyAxMdbgAfPzfz/98qPyLaVre+zmi08dS3m/j0MxbJjRhK
NCK9jspTM4kYnkefehzrj+rR85fD+JSqJOuLU4igIIWttip7NXUXNcD+oNUQevuY7zJewWN73bKf
2W8l14/0FJUc1dpfDi/7DKbLd8suAZKI3GbbKeb7eXzrmyPo2lwogbOX11z1RETKCqtCsu2tWMX9
1H5eVMSsG4urlJZgHhm5pnCDJOjJt8GiDqgfagHEei+oF00xm3IOx19zk+fJkWwjGQUD4m/YcDKJ
Z1pXLWMCCfH6Vai5M7u1Pg3H+5cH1nVm0qiV3HS9DTZUa4QrxKp7x+HpkkaMm0/UEaQ8GUFx01ga
7ZfRLsmojrFiWgOqAzJDTgdK521Ik7HJU/GYFtthDAmzz64ze3KbfaTO5AwcFlEzv9OKUdTVZf2i
zhyRSEvOKkM4xO0eXT9Y03MKk6PG7Hug2k76LL5wR5/blLFhvnjWiIJnRQD+E/IcNhaaoNic6xSc
oYB4EXMQJv9pyDu9hQxX8u7RbTVkUO+yLjSguOXVl5sbPuaj5oCipfttLGXvfeCWiA+ONm0EcOU4
w1qPffiO8jNsJR0FIa4OuqdrrO/yfwqZ9tOHcTS6rhMM4v5PNkxl7KglOhCXTgNq/N4pc9B3ya8H
GxhUwImxKp0XM97WhR5qNq+DXj5KOtyXi5d67Bqee2wNUZpSaAfbkNiNw18qdhVDcje3zgRWtyLQ
194E8C69qX+gvs+gBvkRaeipWgQJGtO8ln2mRGImoF1EdYwlm4ldXkQ1Y2EtkTIuuebuFZVylzI3
gie6fMZY0D7IAbfGnX9GKdSa4M+cMq8zxyVBFiQztR4EnI2aUv1GV0XqwVMWLPXGzGfiaSasW6DB
KedO5IhjTKFMhXInbkFBkLd5TstDQvqmSXfDMG+xbmJQGtsPgPp/J5kfx87S2ye/EeAzVKDj/NKF
gqacIOjOwf0DwjJo64g6bcjwFulUjlhlETSnnhGOoWJMs4wjSunbhCA4ScAXfgoxDBx2WKb+T7I7
dWo/caTNSmjWRMCBYTVo5ara2BbTQB/8S/883+cqer1rxVUe+CcCoRf8jwnUkiMhX41s0yYbSarE
aSrzSiyQLR/aOw1Dwyol5hu3IABjyTt9OHnM8wPTx9ZcNBwC6guf3YwLhzQ8TY0dXwe+nlOh6Nji
2e/5Dg8wwV7weYE1nTScSvPf5bq+PH4XGeBA6aruaGBAsv60xyB0wPGKAJcGI/1GZVIbqRl6bXU3
z1ArIyQ1AR6XKOEy87G85je4dOFp6Gf32C/lRzlLg1P4W0s3OL1bsjCHdEGo5RrhwQIrGN7imcPY
KAb9xeogWiN0UriyBgwB/uT1BWV7qCOY8DZB1Jn+L4Xd4cP4f8BvmhRNN9rdIx5DPk4Ql/CcqOCR
H1AlfhYOZjK+DpTaY5vVw+ib+RLFvIHSRODEOdVWKYat0TeYJ1HF0osOmbaW79POTUmELLlS+iOq
cIOkDziaqkQ7ju1A9NIjoyg6nyjeqX7UEkt+Gkii6qFaELVgYLEPiK8Ww9YAKBNljGrTzR3aLlYH
8jPa9I6DcEv43UvQ4pm/Teciy1Fr9PsOcckAKj/3HkitJg8zHxUqRAilpj7x0GTwae7DZ+WOVyta
BjTLltPG9/RWw0yk3XQSfZwbQpNAQ2xi4Qtcg2AowXfLSDWWNRnXsEg8kV4bkt2e2L3PtxZI69FR
tlX76XpaMI2k4CLgLPStC9wd0MC1n8GcOFFwbJbm3L4gIInlDaAoKQsXAwCByAUmw8Fx7sbRHaqn
TlhCxV8M4UsXmxgWg7HiUmHgBEIDfE6rSXB7DVzLD0/bE+8e31/28caaFZ4vVa8qmsCaohoPgBag
K4XdEUxKqbWNtRbqWLa4eMEk6xC71qt72EgobyCc8RsltAGiGfjABSiqbyKYW1n2BFSSYqWtC8lF
PQq1uBOoJD/OZosHPqM0Ie/Mq/c9yW//WRISjAclSUlc8QOHLbOOtKrtViQhd/xJ5DLKsefdfy/t
mC4bLxsd5Rxp33MolF2r7hjJZFjRiI4PFo1KVUwm5CTS+grmvjWnYl7kAKYvSwYcXeQzYLLuye+N
gh4+JIU3pHulWbzaQmhpTu+xHXdR8uzfIoVEaLPvpm0VtM3WwA4q1a//M/BgwHtC3PID6z6lJI/n
y4hM6bdOEknWWDwxVIsiLHxpqZ23HxBiGzP1cSqpmRI5WdjXHNQfgC1oNyzazGgEBgwbGepp+OP4
p9LP8EZbMUW5WXNgW3wepZzqi62A1PJ4pioaoKdOMaL/I0ZqKOkH22VWf9x0nZhIrWpkhkzwSigG
bPCjjp/1Ef+uT9D2kqbXk6wOtoXla6CYNQWvBF/oOqQJMocnn3AuzGO8TnSfmmLXTjQuNzdRU0sD
fogJBnnA/gm18vc6fdMLjuZzpZLSK628c2JXwH8I3QIKfwQYlfST0+qbsMo+pZRonysdA/Xf0a58
QxrRUdRr6ZmLnkZXDJbsVUM9nHNgmP/yeDl2nnSq/opOLbCKwuPyEG2ZIlseeEYyqCRMXdFU589w
mmNB1NaMvn9H9h1q7BO6CSc4D6nD1+2UTDSVuIue+gMKoVfpWRYi5Vo3NVM8ig9KozyQmmrdXNd6
iMowCN6hXY6MD2JMEw+INueIbDkjv6p0oMyccXhtVGaAx+pyO6KrLyaIqSCDnYbDFHTMorrI3fKN
r4aufZgGBfEWFrechlp/4Y6Gd3psWgJsVqtlJ9zqr/1Ky9T/sys+7EZ+ol13M/qwcNxSYXP7Pklo
rgC0n+lhQSxRM0ExGYNjeUZyubuAc/NM2c/ufoM9oif3TnjjdPk9HBDSjIIElJss2AyajsxKpRjO
FHYXXQ/0DCOgXTL3vwGqIxmzOAFHwwcOQuG0fpOMoAWyj8DWDepS7eUPeMXsF9phTsYHcFdI3VBU
9jDsqLcIlW70Uwc+MMnZNyTvLlJdZb9ChWcvZNkXMKu9XggpatazT3lHDVTrlGE86RYWToduUmLb
WJr3Tny7oPAIFBSrXU4/GwIkB+5FfvcdK+catVMprUs55JQzYS5o1UwSvncExobpwKgfSF0q3vZ1
g8UfzhsHIUeBoh7AVpU8NTNpOqZxtQsE+fFKeuW4S38lMLw3pOpPvolVdy1/yS/Z8q1Dvizsfk5G
nVQPiZvP7K5nN5BbVZtNhilQXwNo4moh9YAwtcZR/hlUD4uZfZ3g4XMDVbO2pShErGeLMbFdiHRr
LUnnkczQVbMws2BAPgJ8b9PhxPwUN7fXRkgKzLgfLpxniY3GXAhcWShGNkz6SYv1nGMq5HUXor3V
7ymGWiTY7I/Iyj7yTc4iZ7Ln+K9NIm3WNPdO1E8Hhr/vT8WdlldK3cAUJz9dPcMj1maLID/LMQab
LNTegleZAf0PAUi6cXCWFvFGTzp/T65VGIDLhqEtQ1lnHXOF+4ZP9wKOTHW/v42ZwmWEVn5anEDF
+6fjIG7uGU+sMBwpCTKYmjOsC4ZsEkGpV4samvM4F51mVxdQzJwgpPKJugROYtg0mANsUm4LxtFv
rg9mMUPBBysTrjep7r2A/tKVkFrJXeOF86NIb0fD+7QGygUMlxMYlyrefhX0JeWeB7Up0C45llCa
XJFhFSvNZDggmMTST31HFbLvGXUXH/b5tuSn1JLdzImuiG0J885f7sdlQE0Poszwavaxj5QoHKYv
Im9ZmDWH6vJ/oRqCf1fwewrEPaleV8l9VtoQV1hzLmv1nGh1ht6i/17tVt743nkop3Iqos2GivAq
N/plS8FDM41vqiXnYp0oOuMY7v/AbIBYuAs+aIQj5mos6w1BG97RwpX1Q/xBC/JxpLuJ7jJ32MPB
ObbTEbyibANc+UU7SXQENtrMZoayi1RF7ruVmvlrjBqHQTGc3kAohF28io/TEPOKBLYpdpsDFOq0
8XtIwXw7mLhOuYcG0aLoywy639K2mm9KB7ye4ITIaEDnYTWWH3emupGTbssxSbuScIXDohT4KHka
88CZuETqnaLd3aA06obkC3DTrQU0n070txA1YFbLxfdPUv0JqGpSfEu0A2kBYtJ8KSETobXFbm0y
TXnouLKCcYQ4h3Hsxc1FQ1DB9C8vuAxo8s/1enU+zYJv0+d1gScjafsq2dxUIZPDf2z4mhQZTYY5
+tYuNTdXUXwCxH+zACIye7rjgNUQCzE/m54pmZFle+u/AiAkFlJH61walSBARV+pSgWs15LdtKJ7
+j6CPRAi+m6BrHhWr3RrBeIMnvi7kMnNh7/tm98evvgbzKtrMXQTxkBui1P4uMu2mx4fCzEho1U8
F7FAMEllBZtCZUwhxqYfHoi18MeI7FkYtB0+W9lr5cybZrTsLxXi6Cx8SZ5hOo+dSzGnLGw2oTUR
WbBe3PHaufdog2wsfRfJBQpr2c0WrQqHV5xe/47sjC6fUMIyt9BVIfELWsBYoGK0QI/fitniiCSA
ZJJcA3kW1d42AY0bR3rrl3/9G0l2gnrjeV86kSdSBKDLTCahjGK2svJPwCDXb90DK6XfteRfcyUp
MQC6ieLn050YoIw/7BH//rl+OOwrWUrrdJRCEPmfoT7upeoo9Xf2TTwEFHdaGkZFS5wLZCCZ4+Ir
G6yniQ7tjPUGK9Ts0OhNXlHyio1qKkjgkserklRW6NhNh1rZ0Xz/tcX5+ZvBk0GHxan9xcLuW//c
gHJtDdPONcC/CaQovpROW9+R6maHFXas24mv1JNgsrhICTXvEJfoVrWKLM8Qja6QGXwlXIXwKvtx
rrFOfgF3EwO+2e76sJYdCGGeR+oNmWHft2jxm+vFXc08/O28dm7l0lwLxSbXr0dVZiyhPIN/izUy
rmG4jFaowstctXVwDTdzx2inummrrjWvrbKVPS2hFuqsNpDImyBaNpyL+Hqz0A9pKM4GfIgFDASW
8ssWUKTIMYY+/wnUmE5D0fcyShscj0cUjn70yoKtL+2v254qed6+Pv41RScPfXwlFXOMChVayAsa
5/GTNC0E4ko+KIpQPuAX3ERbb5yVmlYWcWz/CDpABEP4ZZcjStXkcEYDBXXhBpUOXOWi85h89qou
TrKQXifjm4620BXDSsp2zwA8VJx92Z6EHGJtVTSPZrZRTGAtD+xnRj+v3EElBt7PvSy81eOOhDbR
pTP1JFIrHww7rsoQ/I/P+RnYJGtLWg5kAVZMWZ9JSpWu7OWYqQdrrUZfBHkyNYYSU64ZdLgOe/wB
K8cLSQe1TEXU6uSpKZFutSi6ChvzWEv/XKdMq69T49nrKVwIC/E0NRKlvok8U9Vy0IHbwML9a2Mu
DVtxiJAg0tjWe4F0BO+5aY8XNL8Hdo+O1RSxqnhiOoOBJiDwJdovYTN7JHDE8EwJW28p82EefOJB
QIC/xdLzPCtjCMlvTdGrTk/Ob1DQ02Xpb3SO5g8afbGeAHT8o6tbLMQT7Vk0wfbc4ZpFNHAj5QQO
vzeR2FP8o4qiuWMlk865xnM95sqIy/pJyV5f/Ate/1seV3hzZ+BBiQxOaGA7vWTo+iNAbxZOfl9X
IQbi/Raviy/iloMp8DW0istJC+EOm2ZQiCVDgqU0QNGkRRlATShexHSH8/W5EEaisohS7IEaaaGg
vLOf9echrb2L+pTO5gK2gs/2+iL4w9/modrcdamy42xi6wYjWrmII96ArVcianwMT48gDhX0uqkX
qb9VMOxNCrgJNOfk7VnHGnJWyAJFonOgGgt/dkqM8uEaNVZRDj2pA40V791xhzfAqYfWHa9D+7yi
NFezY1hVA8R9E3YF6HjyHlR/oGnJDjiPf3NCt6sQQf8hAtL4CqJnIpwWUiTr9OzjbWIrIDWmoRe3
I6KNA5nJ++N8RgXvhApcmTV3LtqVsLtA8O81Mwz96V6X/K0vT1Hlz5xnS59Q37Xy/Qte6GfEcJpf
nueROTTaGAv93p+ZK7f+UPppwn5tLD/svtzofjZXdYWmiBgR4FasgD0xty0FXdgOxgGHopXtzEcS
CMUw5z9SLWu5h/HPB2s3GRb85endcgnTwQaNiUqVg8Ko9u/aiEiGCMovIrZQ5PlykBc1Dj6xxwyj
VmOajWGuVqzcVnebQGSf9x/A8ruULOPMy+HpGBGLoPNX3VHTjofDC2OlOS2wRDdgGFYibXzPIV5h
jDwtxIm5a/G1lV8kyzZdGgLdX5NChK3iOary9WzfzTa82/dT2Hh+BGLjlq7WiV5bPpca78d6FCX5
lPUYrxyBtABc7CQB3duQVR1f7etY6AQGwTnwFA/MDcZO8M7Mk/E/6/ollZdtv3fY2Gzu6kRAMaW1
gDCucF9RTI6dZX42H4zD1sjJ1ue6HxmHGUvOIQs7R5E3ekcwcwOcsD8U79qAEpEr58WUgdifpqQH
JmZ3VOTGCHORcfuiA1zkxp3ZpkuN/izhvxcr6oBbVbIk2FcARJpRNQNeIgAGKB1ahpEa/xBESKRS
SDjmtJCWobK/npyp1zXHEJ60Vle6bWXAcsi5klA3kgfXf0LeVL4H4ajddPSRazlVu+Q9fGt8y8iZ
IsnStUe0QI8M5g76bFKNAAGG5ZT9wZhG86BkbYonpTNqjvTuZa4IahDeQ+zqEg/xxvY4JDiyKO0/
bqD7GVxaX3pvl75MQT1i6uZCmpUB+Fd9fKJ7KGPzYt3C8g1RONIw6LtHmg2ZlfTSTTllGa6x1F+L
iudmesr6QfPdPR0sIVPY3qBobMVdhgiNADI+OnX8oSqJF1EXjpOPENS2maJW/N4N4ojMiieu/129
+oE4K8WKabLiB+sWk4Csr9dSEQ0bVxtukz6WMpnPUQGTDFWeZNR6vM/AY8MlUdI+NwDG1jkhX7hd
PluAKB35pGAwlCjo+DJRzKTBTdTgYUwWfv097VhTD1QN5H2PxYCa5Y0fru62u4orgyILf35m+z9v
XyPe/oniXAYAGIZ5QOtH0LR+Seo7sVyTPG02vPwujQb6EOQZgvqeVO+LRFcQhLlECgly4JnaEnme
EVFctgNiWYgXVpQX/UeFGnAXr0aUKK8E2xNYVhkCfxpBpjmxosrg8jb44Vz9Wy7IF2tv2AWx6Rax
rXf+ENeA3U7rrF0KNdcsKxqvEmCojcz60ND6ZDIw8Jz5OWptBDaZVG3NQjYgjaCxm0RmeIaPzmUb
lwYuTvMRsw6FbKq2TUqNtQncnJZ1W95E2btBlFCuolWGVliMITiWqp+gGAzG18bTlwqJpRAtjvrw
OMVOAxY62zAlTcP1iQiVfSj4F+EwsT2HhJWk5ymyh1DO24Kz9nSqES1ruFTbkmfaYnK3tC1t8qIu
um7V/nf2KELTYaHFcIBbIzbWeuNLmn6AOe6FPycvghkSRBQ+jCrP3rAaq5cvVm+Z6cdGzIpS/9Z6
oe0L4tdYPAcWFdEhpjEefsreHW0u56JcPwb2sXMB4S/HqAt3P8zDsOIcx+wIr5BjU9axJNBWcy+8
zqigvnQZtYgVZKAzMqg2pkb2ZcImXHBxg+F1fTBDbY51PkLWU0/fmKoW/wUNT+aIFGbJEwXQrpvE
dqz2YtGaqVaC6QMMX4SVd10EpPSaLx6URTB2VhzkcpOioXR8jY0gpXqKtgs9ed2aSr0xctOx6KSb
kXl3uNuTjsQR+NG1+6Tk8OUarEDMeMw7nH38hKnNjL+w+aA2SyGhwWST/tgJejgRVVOcJ5iXka05
Zht5hYtwMm863rm5J/t3+SexwFQzqisbd22AvE/WT3RlSpGdvb/C5VU6n69NMEj5bR5a7GC3oAxe
0nnZnpEW8B/OTdKlFySUe0ggwFhjTEpp+gy1NsvHJs3oC6Pv1o3Kwe58qPoJHiNQb4lwtwg0lF/j
P+nZMk2W9xZSyG8o2LToDAYDN4OPdtu14jY6YipWNHUHuwVAQsc6crdtvzXQ+XdJgxCnqQS5CuzY
L5s02MkzRWolEs3kBIEymMySBZ5oj/LrzDn+0DI5D4yy5+oZf8DkZKx4eyECjKcbVZ7z146m13nx
QQ+ivjZr3tgyOV1RvfTY/RUzqvuqSEM0kNtaYvsCluMzLkOSg2XZ/5tF7zoX8CiL/fWAOj9Ql+P7
IuaUGY+muaa2P+G2eD80SeuoK2AOw9Z7aWTtIo3kBjYTzOO/TM3Hi4slS3ZTbz777q26uGvz+IeH
x/npkHspE/8cKobhp29NgCBi5G47ryf+MGkV4OXwYoovwxnPa5oDcHb2iGe4RwerEJti0+F3yboK
ChWfrbXMnpI8r2gWGFtbh0alqgGqO9AFG8aR+r2Ss9WLruSSuxRdKF4VnG6SOYifS0cIt+HSaEKR
aHSeOaNMBtC+1UP61hzUqQRr31kPI95BMF7uKq9ZHvpJKbsyunfYNSRxZ+Tbc3EUvtck0/FiqFWm
xYBqvLNpfRpeNR+7sfzn4bV/yhXtD7zLA0F6maXUbC5od40zbIjFs74lO/z33WfZng9S82a+AkX9
HZ/NKLJZyfzOvB2XJdU9ATd3FCbBXTrh4fbWELzHzkEcr0Ka9ydid95yaT99t6NJ7DSpId0Tdpj6
CurDlaXYGuMF2cbKo6pwVlhe3amCmmxfY3it77z/51alOza6hw0iFI/mNSvlG9r+gVR1mrLAT3wx
F1IFm9Bws2njXhiHABN6GYIMKC8Ny4/2kmyJfRpq59P9tdeuWCpKc9mrQRqDY953ap7b8yhfnO9r
9oQIXF+aCFApaeHx/bapAIkOCcEffawvfge8jQfFq+85iozlHD7UGN9Zrm8HnQwTjUnRBvrN19F+
QwWHWdNbhQ6j8FhkmjcQzxjnyuPyfJ4if3ldE80t6QGpdZlZBASLm4kbMqtb9fguRkygOlP2gPfB
iQWuCSu2Bj7TT3sbMUrXSDw5zZNuuLHaVgnsooVNCBVHkGxQxgpmsPIdqcg7GRcpGPiaSUeMcs+3
5t3d3RbV1x8eshfppLdEHIrXrfRgaTMrpv0OCwUgeYCHeNgyL6Gnm+Hh5gMPg4fpqgy2FhzXV6Ds
em6+RaHMwDnK9SRX6OlSO8wnYpZ7a4UCbWQ+KZE6T7fd3iuSPX8e5KRSoCMC7gOGZwWyazuK7tqX
z97dHaOskV/vgu7IAY96CJb8VwBrImleX/B1u151RforRMR29HD9wACjxncv1RNAG2wooWqHlGNN
JNfhFFLMYpK3sEyl2sc5YVTPE0LaUHAjdcunTnlxncPZ6WsioTju+tJR4GUKZsBUsJikGD8P93Dk
3928FSTMmz68ckeaPqHDU1fysCGq6TnRPbZ9YKtnZlSAXor1u9pd1NpR+MO01XaDLZSUY6ywCgGh
CakmL7cFmpqKSU+f7lrNxABqSki4wJIqPzmzenMDjvAjSB2QoXMtAN8gz3F5XhdTCzoduPmUQv/M
vbiV5pQ+p9mEhILD80QLJ1IJ04F4looveUl8uIPmX8BYxc6s4u57nxtWNL0iYih8XYEewhXoBUdW
QJAltI9Kg3J2ym+GUfNv03Zaztzz89A/e6dworC1CisNoW1CBhi+UpK4qyECErVegQiAekbEa3D6
vnEwH1XOPVENX8luZYa6gSXDkrpireRWaizsmu0vG30jqsEmatNRDDH4C3av+ir/Vo7WLhIVwVMZ
rcivPya3xcWJAtgAHLXvpbJUEV7KK7f7sVTP8EzJVEs9LmqcH7mzFPiMQZMF5PN1PLhJQWb+Nct8
rGt45THLciw7jmMchoPVhRdOylNv61Tdl9UzgD9bLXlnGrvPevSlVnTvSiRyom6+08R774CAuTgk
fEg821YwmG5+Ao/WJNfSzcBRNCFSFH6bNg5+sELcL+K1H5c8hoxa96xWWZLD/YlRupygU0MUex24
21tMCu6g52CSSPhUZrk/XTM03bFiPuX13SQrEP+AzLiP56BBSc0erm83KUSaI0P4oTCEh+J7LgzU
1kKv/rft/JNE3Jo7MoM7R+3qM47IJdlluRsp7beAfruUnU1asdclmcsD4iXOD52JU8QaxydTGUNb
E5VpmJeZGhPyrn0gK6lPgJcsf2u37nFn0dxrz73jXDvaYohCgUeaTVB4ryz9Kr5aHajEzAPFjFX7
tw/UfNVvjHLLBjmNrtG8rxhG4AX6lUJrtwecUi2AcozojsAEx4Pj9xcyYwOYp8WTLusFFx0vjeLu
MFjT9XIf4yn/XAxMo6EZ9X5uxnVSqN0iwcH+Cmyf5/Yx0COZ3gxKtH/yPeQYcx9P7LZ45+7A6jXa
4xvCldbo1JdoefCPaiRzPYZS6Gab7aGkUIxEi0AcHuKUvz4a4H4Hc4/B/kxEg1j8TyOdG84jo6tH
pavPZ1m3ttNRKe5n10UUeiQc537S+bvswHby6Un+p64woG0tRR6gd2uH17Wv6wZShH32d5+DaKUP
LKwxgUIFEhEaAnPr/uMGNmI34RAveTJBkKCLhcNfod0aCWTyUxkcDH2JhqA2HVwTFvQ5JzJd7MHK
xoDruRiMRbOQlXl95NK83rAFzo5CPHyiqNpzwrLV9rWZir17SEgJFvh3CbWNxB/3e9UzvFU3X3bh
hVcmMAdeHVtgycHRE2yZujhUrtF475tya4kJKIdfoA61ySySCdF9NgfHEole/l6+zjnhQMdcOGtJ
FMCcYGPkysEkUFL/acX9yVzsp/AHme/Jdr7Y+8woJH1gCGGJHrceLfVY1ptlVb6TQpkVXu0edReT
D8QAf+b4nij/zS0pn4Oip6+x9DqqmkM8eLwHx16UVd+LumAFkeib5ssN5yqObBP8Jq+V+D+ra1+q
zHT8/CmWUtFbyfg9DVbNREVkCjKSa42jUnF5ucdwqr9fo4rlio0yR0GJ6MpNH9A695ZZsI1ZiTlN
SoKypQde+M3vLTM/SvIm49yow35yPQiPocJEk40ws+DGhQMkYhMbI9Z9H6gKQQzH6pbvog2xBScc
VFTB5KxD9uQ7J6xCmsvgamXqn5kuN+C0FSinTmP55fweV5RzZ/+AGEfjvxwYNGJcjaOdGx/Nahr0
XZruI+BRlPQla34hFxnJ6m0AiQfhw+yAVGZqQixxSGtyFbocFu/Q3/R2DiS/Hm0go/vZchjlJjH2
0hi04vynsVKS2BRk6x9FlBwe1KtHRefhKOn6+jGZFF9l9G9Ue/3+WU/Ea061QV8vscuNR2uGqbyS
492fseXH8tmhZ6AG9xA83hQSEX1ALvK2qMbouwzfbQsOUFPCQb7aqIArbMEU0dvs9xeODbVyz05z
rCDYcXF9sP8VUOolVEcGpoQtp5MmqayhRhA/68cQzf+YZXYAVfg/Y4tnsyZad5AErLa4W1IqVQdg
tlOgJ02fD2uDyEoA0ExvoDZkDFO6cGi2/D9FQ3dopNmAATX8XnmOj2zJsvPF4e81UMjQKFtOzug9
e24JdjfQskc1BdqBvYrlsXBlWSwYjOwe1ObatFPscabGplbugpVz1GqrwCPTOR+nLWdjybPyBWnQ
E+SqRrVQIWhXcZWAVpBm4zsriVi2gbMxuGFV8KBstv8fLUSlUiL+B1R1FxC+/bYZobCs5N5glcHX
/Z3RVoHWOM7Xy0cI80IYcINyF8Z6gAWMrxynfAxQwR7n/mm5x/5TEddhnojA31zNRvna/rnLQWiR
LHosnMv/uiSFfgKIFJrTCOJGsv1Cr7xjy60tPUYYyRLD04NZddMaV+ohevHfiQZbuCaSW6a3JvWs
UIVls8UiPKWL2DWrC/s5J9oTvHTxms1EXl67P2a4OBRrfvNYbu1PMPt2eUQNbvHt/0QaD30C1gUR
NRV8KjKw4aELeFK5x+x42fbcG4DyVi5w9eMIBeRFbwp4cml0M2SgpZlGPQrKkrMZWazcvAeAhRen
lhrzz6Fj61iW9m8jNJ88nOj+LOi/RBxSEMEaE0Y7AoLaUDLcMuIOLCsmTHZEmzTmduPCsXOeVcdR
G9OsJZDieG3kk5RvQLOfsWa2u+Rpia7+3JXvCdID9pBO7WPtdULIuyC5DkgfSt8rxEBT48yxQlH3
imZ3gwPBB+s10RVGZk8oUSgxsT2q7pV4FuE7eJ12Uc3ez3ubAVneBn33jPF7bI1sPFbTOFTSKLhw
Ntwqzzs4PQwEp5lbfEVKr86KzgGKZDM9w5OEiu/4+zhSvTdMI5mDVf2LBf2ieyaf+3rv13auEjs4
Me5l9dcEaGq0RqPYwVh8UU7fYtqE3/U7WEH3M3hvswAbu9d9ORUY5eqkX6BAYrgZnbfgeWlKCEF/
sd5dCNAASN5WK8gWJM50hb0MRJ9jW+DeHkt5gtYiwVxKTjy+cr+tj4z6RXHEHNajZ9PVDmPWVB60
t2gCVuub6uxnUAJ/MHvNPBE9UsLY8JE0AFASlntJqxQbObDgPSt1ctt/Es6X0/Y+av5aKgAg7L1o
0bHY/t+wyNB1m67JX55eY3vq7TFAhA7AjhPZGbRXziHcpl23SQeEIYmg5f8hl+NiwIt//Y6hLRmq
wxbJZ6thuCaeKz5lmKkQUwOd00mCzNtsNU899pFvhLWfkdDg7YdXmTMruFUOu5NEGT4XKQG5momv
hsyUXI+iECKkgoZKZjwOi0uV/w3LyQKCQapJ4NtvowP1kiEhlv4W8vnubQnaBhg9eLXCl1ll9FPW
HGEOENSrQI9NH6z6qSUgVNXlz7REf64hJOXtabbv0IZoIJUKMrdjdpnFvfctxxBEv7l8vyJbkIHN
eEk3WTDQdKmEPduVlNOdDSEHCY9OOX/5bDrljk+mV7c95clDMaU9BWKI9PUwyXLP5MDcphj5MjT+
o9u0+rGdhZ0O/wiGdK6vtodzZgUm3c7Mo0qB4g+fLEABZFScOCBlHM73SdsNUGmzAQLcfideee0+
g2M9RMpsQuz1dYLWa2us1dVL4G9fpbR7xLkISLgGHeRnAXAMq/JqStmluaWRazpDDMNO5FSG/SUI
9HPpQZyQspPR/I9W27XEY4BgCpPEM5RIlEJ/Zh6AuVKAt03WP5JCY3GuC03BrPpIhDIEAdLpNKp9
u1SdYYaKlDrMMf8D15JC+HZEtyDSYuZykSi4lP+cORC+OQrYlPvuqjqRPROO7Uj/uXvPPIjnwx+5
naievDKiLSIzNfDiFMPiCFN0xqYV16HaA38ZKccu0t1+PXr4nM0RD2MhJfKuYN6z5A94MN4KKlZa
V9/3qPzqlG/HovtZWOqtgT8w+NWblMMcuSmZ3UGWhPwWyb0h8tWX8qhnLR4in7Jv08fB1gUGlIHT
hWj4hzO3ya6VOl3RE1iBByUsr/7rm0J8htaoDg+JVbJ3J7Da+u4gjrftFdbcFCrj4k4VA26NTtMV
Fs7rpFZnoeH2telFBQhJyUPTc/QgLAX8qeUB7WiduOeDbczubHZwagGjK8K4G9KVmdEyAhB2jBo6
OmHbHdAnR+dXg5KIaNOjqfMaJ2dESWJpmbdm/jcXCsY5fUOoqNIXUY5mPC76RbnOr4mR5VCYR5qv
1HML/w30WVI0MnDFnhlJ8vD1GtdG53QqBTrIr50sK8qP86iiLfOC7hr1J7fH0jeS1nyBu0TENbnK
kWer4XUq6Cid7WyCIz32yhmVTOWRLCYnOSlNHdVQ+eZSbCeBiq21gC+nkWSfbbdfUvKrGZY8cOOU
DAcVfWcBfBuGgQhkQIe4Bybmus5fDA34VviSN8lB2dlFmWVp0A+fkdhHQy691j69+GbGqfidWMID
0Eqzqvf9GZTNLSCEtQWONLiFJc+9mNN/MQPcwTaXTN61LL8TWRLILrEdph5/LX3M8rUyyMn10Ljs
E/kRjwNi7knZaAUfROLLKuTJ5Pk/rmN8gEIeqrNIC1LQBhDT2Ow6zu3tgnIYT6HZZR6PvfFuAu/o
sp+V0k2lnUloAdgJ+7REXN4STY1j1VfCpb9w45hz/iNqrGB82KsCr2cvjPcekG8L9rOLNF6F5KJ/
DAcfUcdhSgY0OLObzYGvfJKhgXImDC+FNXVFbpZKgLidmZN6igD7dBFNu90HhamL6TdNMdsrX9bj
KEHtkANaEx7rb1t4hjZrjyMhosbpdVJaNsM7GuLcWWF9CLsuOGXQl7fXyNwXRWWyaH8zRUfeVYAA
cOrYCZ1Is9vSCpn1B1wn7D9dn2QFULRe9j69Lbc0P9U9iJ6LDyZXDB5XDRk2zW0a3/+GKPctTflL
wiwFtkAFSn/1N7gb5ak5ogwY3pN9kXG273mbBM2jE39hEcCydcLg9fnljzU+elxtc/38xOE0uyZ3
xlhy7I5m60QzaFTUudQSEv8hA+ujH9Rgi9e5H7jo0GnV0Vi4hhRPl9BC7gW+CyGjeP1N3jdOY6Pz
LqOdi9PXTPYA9zB7aZfcA57AKn9TtmhF1b42OiX58HG6bcITSYUTiryefd7bb2w2MAoEbrdACEsT
aoXaHKVLg/Ryg2HKS3nOQW7UUSDh+5RMnYaAWy6u/OnOZLq7GUiMM2oe8rQwHL7EIP12e4X+kbvt
+BskOh+/JYa0QaM99YBvvmVhd3+SRAjyBZQNr7RqdgXeo2UDjX9ObIrLCBVhtb3TCPS5RLih9Us6
l1xQ6ysZU1d9e6XprtM/H7aUx67popheimfLugGZYsSmrOg2m/Pceb8jA0amTfa4pl26TKMiKk+k
Z2e2c21EsFwt34nN7OYr6LrsVoh7oLm5uJGZw3CBjYnQ0ugmO7gkUldija6tClAoeXZK6FLC06Tk
mtelPInF0qvPaRDeEI5fMJbvPLLuEBbgTN80xMQDGK2A3cIHsTsEvAgUZWHVnCqkq8xd0GYY2G7Y
PmjRSBLNdQuyNqS0lzWP+S4xwSgBjS7d5phwT/Ck0rhUqQj09Y9KCp1O4c9Ry4TFfvdGeSS0zOqI
hR6vGmU3VY8CMuMEP0WQfe0S+RROqgG88vWjA/9jLxmOEoGQt1OI+MBgHUUxFQcEZQX7rjWmKuu4
5Vrr4bPpBuWiKiSziw7/ly4SvkIosTKb6OYC3yaOzyvot2Mker4kNTyJWL/80ZXRzdvSNrUnzBIQ
85COEClQ4np5UkFCSjyRF86oYu0vItMxctc+zkAbjbY12+1mLctCqFmEouDdMuj8gflCvbx5PBv9
Qf0pbmXc3Y27rkSTJIickhRTgdalZP9fQMEzxltIKdbop3YdXV+Hu0YgyOb4smjudRybe52FkLi9
6YBC30Cj7WPsQIf15qDaOLrbHCOkWiem8K0oIEIt/HWVjNDrwJNzZPEPXYwg7+c03nAmXDlsPCWk
JIlk/9gFtqFvzzxU7sFp6fqij1ImBa5jEHvlCtOCPAzi/153KXf5Gk/3MkS+KBtrtEW5D6zv8GGH
sdylGpDEE9H6Wf1eprvz5YT562dKS8o4lNRZYUDQ5IoSYLlDnBZpkD9taGjRIccJFGVpV/SfDhfM
sHATvyR1+VxOUDjLfpW84m9LkUqRTOSKBkL1NTOmAUtY/2F3NBsDF4oSEqiV3BSHf7Ge++T/Y87R
UCeZNsLwMWs1wQPt2E7JDZtUxPTCptcQx6twBSk1uULq1kY/PecxHbnu8DhqNqNVFtwCxJAR59kN
CfiYuJI7kqAJOuoGAITuV387ahFEgaWFGvYNw/rA9vNb6zAJrePQavkqzntBLjAwNPIIx5UQjJv5
kquOIfT6KADVHEBj7GK2dk/tnKx0pxy0U/3qy8qrAzLb3HUsTfSsNZsz2c/rVMZPXrB0QgTH6n/W
ASFxHDbUjpaRMwJhSWe3jEzB3fkjKw007n0NkewfN3nC0IQ+NIVVqt6EVcx3GAxFxPS/qWSxY4V7
XkJmZ/ufTtgUnNdyU++g23eyz5xR7GrSqqwvl3xZ1oBNOUIK30unzzlrV4Es/rAopY7FWOiUUC1J
/R201SiQVqrKsdfy6vqSVvvQnvJnakZIcEUwYZUA2CA2ct7jSiLrdEMYC+ub4v955AtHAk/xGQsr
TKSeYyQBXcyrVPITBqhLZHni+ngJoaGSicEqFNQR1vvq5bEwitTFskYFGPDcubNgNv5AfdfxUl3f
GDbOWH0IP3y/QUPKB+XJUlwFdRK4IdooKNgeLi+NR9zhrtMLoh2zRVuFK2PD6wdgDz24v9hcBk9X
6SNUuN+FVIP2ZC8gY7w9Wzu1AvsLFFGu12VHvClPz/bjB1NWj3Ua/UgFhMn6hfoQTR1irH4XYrzA
CQJCyGiiEowe4KBNSa4ZO+T3WnO3bF00IF+djw8Ay6T6CWq3o5P/8ZcSXiUGVZUOjXGy2zzTLnIL
g5uYnYy5S33wHyyAZr5UVsHlKqRYtXhWMaUt0IsnBXuTFYQ7rgdHHQE2pqgg+LyNo8ZhvX28vQ73
KbYfIAQ8vD3BMvORGx6qJT0nUQI9MhGm/DB1bJndb67gkrDwhSd6yMYpKuczrADh/60R3Et4zfNo
UUBhiSo2SvqPhwA0dibl3UjfTti4SjGoDn9S0E0m4UAO4RSWiWWyQgEFTqpfojkC3dcCh6DRlzZg
71X3tkizAj+opDo1uvrPdvPtFTcBaafTHS46mREmKv8CJqjosm8Bbx5gdhBZy0F2/HBn3HXe32s+
ws2eaNtNqFwGrQfSeo5YdSaeS1pWi3Qdj5rEseDWHgiJLCJ7lFa89JVIpb2IosDOfUnp153J7gMl
+Wr1HMvEmqo1lu9k2wHF/BvR6efwOdoj44AqROJ/RfW4/jDxX3fFoaFg79mO/+uxjnmKzphR0VNh
qt3SbSr5uGokoyAR07GsayTsXdoXJi1kxNe0vmvflMQrymg72MLCr6CyXtXjjk+Kf9pHoNdVE4J5
dWF/QOOUxaMR9l0s+uEADaKStW0pzpFn5O2bJyEV9TDA1t2ueSI7HuY99KlC0Yrq+2taRqChfuIe
pm1XrNOhuQCRGRUymYLavABUVsV1OGaW6UNQaOkoCw4qBs34OhnU8sCgXtA5CoDBAPJDZWapuVn9
2K5eYf1CCTqAEKJvpa67hu4QYT5ufT/x7oxwWeIJoaNtjZrr1lC/UbYa6Icb4U2nnXJyrg4ZvraY
/sSOGVKwXS8++MVmVJ0o0Si0mNN6lRCmi3fHzyI2vhpXoyL2D0GIk2EdzQvEGCeRxCtiFszpGVPp
Re6yHNtrdPNjnoPqX3bsQn//q2e0gsO+dqbKt5eiVa3UwvpbMnoB0ZYPVMoIwEnd2QmJA2Euj8u2
fx8NRjYGVeTwgURcWieyVscRYHIl1IsY2dDqBjOVBRZborUl3dARgA73yPpHHkUOejNllfA0m2Dr
K3oFkBh5S47kumwPYuZWrQfj92EwYHlwKEo9fbcPynf95ytDkpC8YqTxPkg8akgBXLkh5gXNDLGz
cjfz3FXu+zTo2rNLnJqyIq7A9l6RCmE8Pc0cxD3P+KVgs85w0Vx0JSb1aE+BFsMtEzBCMnwmIqNW
7/GhepDtfQTgDGSrJdacjgvVUdGS6yVqt1u6ItLs8lFQ/DJS4Q89oNyRiqKBzoeMn6rOOWIQsEoP
8awkcoHCSwLZngnyvO1QzKuUuepu4AhfTK6zikYsW+fdeuhgaD1Jft7pAejRjdMwSp1jpgllveO4
yOBg9x769yPHvmmBaCokGwkmhwLKzrwj90NDUPtA8iKnpq81ksNjMyDPZkqh1iq7ciCrXyYJBCP7
Bj/7p+3XpQz4UrA6UA8r6IkryC6c/uXr47pqPGsANszhqCP51kXOBk0YhqRqqkAnxa9M6Csy+xZn
ou9V8G0uoKSB6j+9XFnkN8XMSq8AaqnaAvlif+ES4xahHp72tiE3YT4ooOE0iueSJEy8HUWIfG46
oRdFenD4U6jS88+o4L7zD/hPmcgFaucipQXkq+ldtdZ4CmkKnKKtMxOsdr/KNNrCbRVlA9VvrP0S
kvd/lo16VfZSKTCo52mVBgQ1qgDB5onZHP/00lWa4rKz7fJDuECcE99JPdKyGEW0pwwM/QTXXU3r
km3Pded6cyPsSxwjNcVn6ZeoSIgeFAyB0jgZCrWfqeXWigfO/0mFHzCaS0LHMilsw0WDzdA6JCe4
iV7wDr9CTecKFRAr/O6HmbxqNML7yRX+N/rBEUEipcNjkIwHA6ZI11oPrn2c/XCsQsXLCn+DFvBe
IfdlmqqDe/6T1Kfs8w7H8ue+vdZWTghAxwvNcANlbFGuXg9ILIHDGnRto1BDNI9+VVEohQtq9FgQ
egilpQkRN+cdl2a6AT6a+rvCWozcPhNSnMJLv8aHg0R4IHypovcbZT44+exxd6q2VFlxx0stLJoy
f1yuserkrQlG6oyqGZMJSEyq4pxUviyeBbN9cFgA2Bw1/snLzzPXDxsxoDZ6pdmCrN/KRbPZnAeC
OI9r5bSRWAVwCM8vyCgheCDnyHiYY9o36V5ADUK5DZ7DkM/UE0oKFnXDQWHBQg/tRm8y8/GsOuYK
6++9OTeMarPEDOAVxb0uo9NtmBas5mbGWF9M8Kc1xBk+EZ+hu5GVFjfqzlRNmcSoKyulGzpLCazI
3ZHa99C0aKi9uPelFS3O8ebkza5s/RcGWFv2z2NlhXUKHl/U1L6szXrRoBVhZaBWMO+Xl9KZ3K0F
Q41yq+VpUP3urPWHeO+Jr6apsGk7XnJx+RMbKAU8hwq0f2F9lYig/xCQXu36EaBQDEjhd1RBlDgB
QLBMi6aiJoZ2h8gcndw2v+4b4ekMHe+EBtvL+DtrGIjj2ETdugBXG2tgv/HcqG6Tm8iV62p0uZhh
/8u2TIs73mWTIoeDuqCvTdb+5ylagXL+b3rBhChBhWXfBeUCI5MDeSSZrRjr04PvVWCq9Korg4IY
eCuIOmssx52CEqfUHFpZukvZscfs4WL4mZGjJ9MUDpVMg4Dmj7Wwmsq4BydP2+d0mAqwReh7/EQ8
/+Xmclp73H2rtRjBA6uSffQw0dVWqksHSBlSnpU9e2TBt25GP8cYpykJTFgwWnthETzXRJJYXbwc
MiXGPYtDfsgHXhkW49ZGUEHZZix4bJiKzforcpNPilKkpgE8e72/PWV6u77Ra2qBY1N4vVREx7q6
gNZKBOoScjK6q6h9A5b8m3XKoRx/YME/RcUGNwjDdiQhdgnbOQB2Nmdix7dqfJdnsrwEGbZ0zxl2
oOGdpM4YSB6EOMFgA7/60kco9Q+oDsznZRrdLKbDOQmYz3x7OrgJdrRohw1wNKl38T7+IbacuRqL
Y9Vk+FwcsGMXOW06Q4KJ//VljO6E3TS+qB8zO43h4D7SjH+98QoIdXBW/HwdBemqmll/VA/oFYZ8
ijuBicwc9s8cVV/e1Dy69EDP5mshId3r0QfdG4hy4w8H1BTqI+eJI6JwEKO1yDgF/jBNN64nK678
5HrHgVzZH82sHqwcBklk9uWmrli+y+H3KbGdfRlmNnpFtDnTM1aF3NNCRPXd+iXDd2Uxgxl2y1Xz
9WEnDRQyhibqL0its/+vX3Ha9bMVRIB9sannaUN4eQtMu/bfMwuaQt2bYnuXwfaJCSNBNTHvztKh
8uokTqz936QCn903nzgGs2quWSHwJpaP0JtKxjOvpVETOqSwvfmuy+mAgJCIAsKKE6PmStAUU06j
jJts/yfmRnK2KYMwD42XY+9hIY3uumnC93EgC/GXUOa9n7YEs0LFA+vP5rJAlCc9iM+mh3C6Xy3h
3hi4YX+yZcVpVYF3xhDGFds6CUk3qRM72/n2elnhuPYJVLCbgTSSRAhQaxGXILIwB/3duzzd+32H
XA8R8dGtQFgYNlny9n5KjRwvGQA1Vw4F3JsBJHijoPn0LfDLxiXlclp54/n/s7CsyXUxnPoun2eI
L4kqmlBfLXWw2AZjLOf6Uhkfj2xkCX3M4LaO1MlfXkHGmFtMZQkdl/Sns+Tsi+DOXkRZlrifulGc
2yJNI6KypSJZjPBqY5Re4H9/WYYwNjGBoK77rXe1L2CLZdPh8KqnGbU5apKCxIRkKugMVsxUDLW8
qVt+eIURdp7+WOMENVB7c6J2GVYie1OThaDF0o8gTM3A4fBOLbEPjRamRAX8oVkyZTWjwcrEhZoN
yvKJpE6bCLqEjfxL8gH10nN5Tj0umbjuwLy1GiIPJumCBamrGOkv6jEASeomxIURW8B0Z+Z88Pup
/E5kgtrij4eSy7lc2+47IBGa+doaKNghCDYpy6VlKtFzSeUtuvXIdYYXMM0pm1iY2u4VWh9kPiPz
FaFMWEh4pUOosEMX/yeLZaWDik7ASKdBQeyrIsy1tAnO5/5ZooV88HFfZH/+ycKCaJ17F08PNUyL
kokcZw5cO+TzXdIVh3aXv1wydlHQZ6aKBGgu/3UOlmJd+or5MTcrK/3nRmk4LQT2DOJH91ojKfSW
AvYbHTQqJ3VCxiZdxcLy6UOctExLtN9TzJ2I4VXw4Ntiwh2SM8uYG2im6q8ZzfSj074B3NxE3RJm
hHJON1SJLW8cJYTuFzWFUTO4lyS9BnXY210DsI3UEucBRzrN/oV6Gb6l+9xsj6/t1r6QMtPDql8U
MniP59oaQfBOVecxZxlovLIeVBpv5D3+S9B4RwfzBemdLAQyPh+C337lsxDGKdPL6qqMNj57p45H
jmM5xbNUHTtuHbM8rNnylcbYKXJQd6AKj1vi4KbcPmKUQkdUa3vCTmL3paBslYAVAluqRhlqfIPs
ZlZeqrqnlnfMPjoHLr6p1kom2AMfAGuURvT4AQJykFc28jUbyZH8a98Cm23eZacPBrdiKp2xKCGH
5z6uPfFKAot9T8VEi3K5VLT7ZKPKXzk4sCGxx8vgdnbYlifR1RtLWX1T1O3/l/T6uEncPz5hFkqa
hIEZkOswmXft9wYcG+602WYxaGLK81RLtY3rs4870heq175me0iVjzPI4wiAmOnSSh9k8iLRLLrr
09fkXdQX/Yhda8O9A2YWNOU8MGbNzZNMdrSkhgMqzQonidkM5LjPRqY8xIAKc5MJFByr7JMOhc3p
kMPvv78Wr6an4Tpw0BeC+Z7fP1RUX8dEkY151EpdHr5FcOGdsWP0l8RYD1S/x4hGCgVMuBpiySef
x38ILV2r6CVb8I/xIRmV8gETpikX+opHX0OwNtQCL0A3KFhHCNDlp/agNJ12Wa1WUiTASTcTLwhD
2oTmkUh5rPcxBKgrrMrb72RkTT9aQLmnpW5nPFq0XI346T8KGTNdO/qqTLNzDCuElko2UlPN3uOg
wuCkieA85yQsGQSBU/TJlki9IMzPXRCm2cnTG/TUIX45pQfyjZYRAdgSt+OUBnKgQDdOFXP9dtMt
4rXEj2aaTaBTYciYoGalip8gldX9CEv852PxxnL9X1KPwwZRWkxTqJ787DV6o/dC3y1vJI+aixY+
SAODkgRUXanYV1ZC0W6nupdcuVpcAp2jV5x2iQwOsieogVxQA0lh0Pm9gpTNrJ0lX+fmr7MBrTaD
DF+bdyWitpEhyNf8zfuCme62UFlG3XjGeKuvRI0u1hl+KQXeHwuASrP6x4Tgz77+bN2Wu/PvTgJA
B6j47Yb89/ymux6pLaTIX9qiCDbiyjEDkdSn9fsSBfZC9C/bD8DVp1NJVhSezSK9Hhi9TL6WhvHf
mz5EQVAl+IMl2+5qgBAW5s6xS16wrqsn6zXDyxnnkgmEYwQoloQeGTKmTm90/xDmcj8foG+Cxyyn
tQDXkhkjVek8qmiQLkZ13A2+wmT9vuBKmD9sDXGGkTYaiEUghHhuuVBXJiHJkXNsfqw2hCR+TYLK
U163dbr0Tgv/q8h6ZnoMmRCWxV6i9becqA676zSu3+0aBgCQ43G/3WfWyvQnF9H2vzlfbEWwCZ75
spy7y78j7GTjbAtAopaPmOXZurJ/So0P68yq0Q38JbknC7NhBlThk3/BXGtI9ayMIzpBn7s7nm7s
WUd86owNdemr6V0WyS6fTJcx0BXfa0uZxUC5BE0rvzUSsUesLIeXdqn7+64urfMt+I0XWfWJ8jEi
tztjV+dVuIQV2kiTbAzZFSB5ZOewEww6pkKZVIL/aIX/44qNt0XFxzSy/OgPcA/LZPtL4R42awJO
zt+qswrsiMuN0TWMWBA3iw7K/wGD3rUDhHX4wMP0du+MC4weAv47uwxW7OyuojQxxtx39EthGF1w
6bayqxtaCk1/MfwTuFzjHdJr0LRbJaViosFh77tjK6Giue5L/2C/gRKiiBW0cPJU9hC2ECpxQ4Q0
ZiPbduFhfpZV0K5taDgQPAXEQiBIptzwiFG2s3+dKAKHMOuBwgO61k/p1o+w9nRhwkBC2MUf1J5a
ZMaYtBgJmKxxPqQt2CKAkEH3EjEMyIzJk7EUgCYHYNr6Htc0EdhwGXBXW16xJzZcQNQWWPV+fl8Z
OKWkG8T5j56zZ86jNCU3eNrebsrHsCe4TqCHm6GhnwwGBvxR4CVISBeI/L2KDIyqL1LwowWNZswe
/fshiwNBtxIVwiEBbTpb/byOU5OBSsRkNVBY+YnSIe2y0xc+L30FI5Nk5XS7psQ8zBN/ZrjObdEy
hhuyAT6yAy5lkIYGB95rydaOLK7L7NEaiJpi/hT0CgMlDgNiTBF7RcfV2yEzghgLxZy1yjWIDVxx
bJczoO0tyz0QRKQ872vmOgytJDjGXxa9Cb4IYuFOj5AZVqZmRFMa2dh4f6K+ASWhwBV0cmApTqdz
k+TiJnwmflafcdWJ8X99UN5bM4TYQnEGqlxFZQ2oO/4iYVIFVUhlvq/DavYoIHNcig9cSfMXznro
8dtLg6h2qwHw0SmOpq3Bf4nrAMC78U7FtO7A8fDHSGdAEs7wPGAik66UVpQIW+UX3DHphsa67+9D
b779OKmj8FlBd89w6yezNIgkVFUEDN5Bav9xUypteg7oz4GVDeFHs2DY36jIASs5dR1eRSKZalBR
Ja6pXKHTuL09epBZvZVVHxUr81QY932pTIeAMP95QaYZdE5gbEIIURddWIzO8zFIc9Unk48g+NJu
KsFbdJQ7NlULoRiFc5ivcPZG7rjY5nsy5TwkzwHfGHq13loC0QyRdkMRgRC+R6c3A2IYfnO6xS/K
pKvI4sK7eVToJ43ZnGlyGfKvlV5FHYJvNYtPM6+E9klPvTsFa2W1mRvQwMc532ZCq4XYwCFHrFHO
/r0+99lWuNDsDnL5IUOlx5KFbpnsCNxGMojuKW53IBsQox859tDi6WHxs7lCm8MXeySQEQwJ8e/2
SL2JMx1FtNbnsVu3tutJ1EkmAV6EFBCWd5bzNvPP5Iooauu0Z6XKfAQNWmUnqBCfh2RZrAn0r4AG
ZMcITzBQIn7drJdKujUX4aYfNlWum0+RCr7IVbz2BfPPFfbMrirOOlXgBq/d2n9zlgJkLQsHuEM1
hDmyuvGKguS03fbFauyk5qg/PFeca7javDfhVbpIF7wlghujd9eMBzfs0Gz0z93q4gfBFHv+otSg
omb7UlBHqoS3alzMTLP4Sh2RqxI+xAVoh06WcevRJLOWc3m1HWiA2hfBCYfvME7uyj43HO8Adzrn
Aroia0I6lnSdK8XKGnaB+4abUH4BZnQlFcXjiF7Gw77pxwHHosCJhGEDkrgPAQyfbIIMDYMjNEcc
PEGr6FztbZ25sVuop2b1loYk/Xvt5OmWKehDQ6I+bfu0WUtBqNcodVCfKSxIFNru8EmpC7/2S5sf
YaW57O8Z7VIx1djOKXIKtYHQA5kVy4/TG51o8JwcZjt6F2+4Rezb6DmlOz8zkhwC9KNs0PKlI2Jh
ngDInidQEDlSGsbgJsqSGlJeIUBr6I4wQ/7U9ZpBkIkNLry1laNEsoI6qp1xnbU+btt8IxZQRQWi
mBln501A72r64bHYQTitlMVNbfBzjdwwlIF3DLXNWlx0BWY2va+eRHNf0P8TYb7+9gUwCVGKbIfH
JT2rPoYdrc6t5Bcs0+u2lj+W55ZeRukahLb57nYCQQhYiaSnHBkseiB3hTy18Y+dJoPTCGf1H4zT
OWgl4xx9Vj+/b6RLWLR5Bep0edM4mEYFKEhPEf0ljXmZ//yigS7dxear6LWz40ZOSNl+GUryiyyp
bMUFuxuDdy0hjtWlnDsh2aax1qM8DzRdSu5ycrnvZZGcIPjiLc7CAFaNRgha5aXPtjQze0TpUUrZ
/WYDQ70/VkD3ZRza9CYQbf5ycz+a9z0NRGo3YZCT3SZbDQ78vLQpSOfifFfhvRZBAS4RzbeuoiQc
MNG1YDiCFPed/bssVRx4O0OJAp92yzN9O/zW0O8eiLTPSyXps056yTcNWslEsjiiyvuMUtrAt91/
YxSCmp8BCfiazaGMlivu33NQW6olf0nLCgFfbx+i0D1EDiHga5mg/SpxiFAgEEq83+DjsA4FYmhu
+ICar8TccPrEtykHihbz6Xivmy8PXDjFAluk/f8friPnr0uXalH9mN6uezNL+9IALgBfobs7fAD0
u4YjJX50D3qaJiZTxswGIm9MRrBmuBSch3PsEAEWrAfpb5JeJWzncmroY5UNMEojHyFpgpZSFgUh
B0CFdB/FrMqbtF2ayLAelDhvQG15VHYzpheon3QQ0GA8deffiIAHZJ/7lJemphzPWA2ZO/SNEK1h
GrJxfT+5gwyJGKfk2P2Ig3IOTAIbiWbs06esnZJQ7XlIFe8KkoLz/O4/tXoAhwQeMhX4j4tp1JH0
bcVoZDi67atxYAEwqbcFTkHFAF+K2P58ha4ZvyUl7wT7EO6Is6zCrbRoJIJGPpEgGlkgwQ7Igz5n
z7jw/nDn6Wjb8iJMfyKk5pM6kDT2Wdrqid3ZTv9XvyyRZ5yGL+IXdXmWv0hKuWbMckbMoIOz6JF8
Q4LzGubW+D2Q/PAJrTQ9gdqvhEE/xrrIATV0OlDTyron6kdb6nEGxIHgR4y8fSeKknI4o+UNiGbJ
5lW6mEo3iMoOcAykc2JvPZZX+DM0xuXlXHNN2dm3Gs814xK2AQuR2cBhE5Cd9IfKKD0RR+AtEGT+
ouaVkat3MBbAVfAiedZReCA6sjwxiUMzdo/uf6IhR9l8sBkK050LHRHXGj5ahM81Z8DWCRSY9G/c
hBJForvbXJ/LiXbuLqM94yJmPuOMV1iwyT1JnOCE04k7IBS60HZHkbNAEcXzYs58iF7rNMzwRSLd
Hlc/FCmpVxXnakHvqbWyaLOatRT8/HvKOWFSEgjZVhIgK91mz8RWDYxSKnWH9/ECM44Gel17Znll
GN/+PfrNki4PqJtHyW8o3VsPBPxlXEI0Iqb+EpSM1/RstDsqPoAn7u3BxbVfvcafrjOQFjNQOi7q
B96td/ymOZvuxZoRru5ATkFiSJiqlLzChnEhfO4Z8yyTT0+x8QgtgUUxOS8ESX6SA3kUXckiXWg3
LIteYJEp4leIFiUTZUhDgd7mneI5bAu8EIcWWXcNxddXqa2qaPt7LdUICnbhUhBVCO9rWDsPVw+Z
yuufcozu/h8vkerWS52ppC1zHbF6hKNo+rF6dET9AIqzL5ZPHsmMDKa6QnHY1sreVLiPp+wCfg/X
TApQV0l0gp0CZn4STys3iuVFdhtpwPrXVB+T+nSVmh/cje/ttR87h63NuIIhsBdZRXhwoQyZ+AEw
P5PQveUaHfLbmVgRTWVcoRqEOu+eGL/RgORRtUxrJvGG6l1eW3r2gJdnhpq+uad4QJ569OOZ4H+X
YnWNutgVI+HQAfs6PbnklPd2Oz6ZP2RmfbetpFRBv6dTi5fK0M9um/zmOfQBWggKbftVWC9bcR/w
k9SDKI9Q9YFhtkfpP795Og1UHhm+U4BxNzCyKQwIYJJRjpJJ02kz/E5ly2oFmSeJSMPfBmnfF+uO
6tTAPxajMIl68OO4/7rV/XypRFTGSpjibpOhJbiE9AlC3TfKVZZDExhlVaSahch8P5houUfUzENE
CWt5oM4YYE5ttNyMZVUUqntM0avNET16psFoAmj1x0ek6+UHkpAg1w69p66fJqAfOQUndTBJQmxC
txiY+OvqFpQd59TAMn2bTrGygiMopLLEORX7kdFMJwhsVvvDmCX1JAZiCF93lBc9BE7uY+mSO7al
fJPuTMExPjKBPvdm1o+R5f8Q4/2RROpGK7VcfB3KgDnLRDyiKPsbifOGpQg0KqA0JuhekBoXNhIU
a9GefASU3h/qOsz4nL+h5UF5RaG1CzWKZ8YDtvXRNz+Sy00ZHLEWl5VN3zwFj/p0AUm6WH7FJxpY
dAahgz5EFxF6m+V0sAzA+qbE7wZd5MoG4KcTS5/2ep9eU+KJisqVl9CXtZxNp6ZWzq1z+sH6AFDW
BNZQ7MSv7HEw3y5pym6V1842oi+hAjGsC8iyvE52E7Z90ts+iFGILFUrT0HUeCuiQ01O+N7ql3Lf
ASxQfyotB8g9C9X0cAoUSdwwnuFJwJO02dLDgyF4z7cDXZnvHYu7gV3rMHaNUW/p6F7ZfJpM4jZ6
ZtLGYEZNTHUPGtb6/d70fEQ/q1McD9ivYPj8vTQa/JZxdPo5yL0dMHpwqcyGokBOtidSED6rM9nJ
Kc6B6mdeLXF8eXL58oOFav04jljm68K0XhdS6Qz/9m5g6O0as8IpysDNpX+e7XP3RPB+yrj3NknN
/uQkYK7MGfKGiZdlnzy0S35lXIPdh5YWhanYvx7fKyRBthfC71QCXmmOvN3P5SrgZcF2pkGI7y5i
1SBJ7mOnr5Kzyr1NCin69Kq24AlLThEFkI2xR3pKP7I/k1HBPIeBdVQ5pouI1pnGNJLidCA9jr3S
zw8QGd8ax7rlasU/1pG+clg3+OnH7Kg1W1Oi9//b35BuHOqBpm60ZHKIuSyuyy/3fMp0whVckyCZ
wJAf/8IZzRApUrrT7F6PQArcqE5S6SM4Wn1AFgOw5Q282fxHdRFA3gDivLR+w1yYKmd3E3yia6Aj
gBx2mf3qwc4c/Pokifu+VI97JVTrM6Syr9Y5ZNccjrOqwtzResrK/0fh9Y+AYQ/mP6L5df46aiQU
5dKjcdMPsm4r5yNEHXETUmXNRCjbzeLkduPU8jNeZqkRym6szK/5Fgu6r+e6N4hxxV+8erETRAIj
61vVNLqzF/DlJY3MtbV/yQlRkUcefNs6OXEp5R303xk3eif2iF0XvCkndFI/LwxB9P5Vy+CgIfFE
nd6Nf9PVXfrGq//jVw3w/ZJXdLM6HuTjDcjgD5Lpm8Wvk0+nSQ0dONde24Xs3l5MfWzM2kK9d+7d
jfVklFGjaaaGCFjeJFF37z5Q5hyW8T9qgViptM6hENBx9DPHUP87PoeCCJ6xCYH4TU02N3eIeuP2
d7ugX4dkz0Se/iwpnva9BzBbM+dgUkGOsAJJ/dunsnTM8Y2yvc3tz6yudaH/ad7LIJhNUYq2hjvX
MiX/hFmN1XlKt6reIvYE/kvCPk52VlapRdjt1vHBuTODUjOxnwmtqVbX+nkMXNSgQ2+c8cJwi7/i
FBuCsAl5iDaiew6agbGyKH1VRiwDyONu6gpYL4qyj6q3qJoW/rCPg2g9FZIBissfZePU1PAbquzK
pLD2fGfk4pdeWTA6FStVs19LAUMXSIvy3wNWr6DDHBLiFV71IvXlFIqY5k+MVnBXtnVJHVO+VVoy
3ZXTSvx5cLyZB8juiQ6nApfzgAsq7eK7qz/55A3V2gvQEYAv6scWDmQbW+DZeiXIqbvJVR6LEesI
h0TYzh2rBhD4cjAnYoVxMmORXr9GiGnAe0oHGIyVIZAslTNKNWHGqCS2HM9Q2TmEcfj2ZFNWYBg9
ZAR/G5hNHo5KMP5bzDZdr0AS8lNGHJsvJm8DFPKy3bDED/DChTEPlACC4HlRTh4YZr6E4sQK/K1v
yCcD1FMbOLkrvIxzULQL1wIFOSjCZ8wCk4RNRYMzu/vqqXapwK8cIXv+94WKGpTdkFh07ANGKYF1
7zanO64XQS0t6nzCofMo8H/hclw20rIxYeW5OoUtWTiAcuMeG7OThZnERXd9PGCGFan0EJPt/Azd
BHb3WGWbhYdnV5qoJQg/+JS4cWW3IYA7KqaKj7Ga6PhSnnN0dz/S1OiHls4Ym32U15y8rlXYarES
w2O9qrOUgOELiosN6JZMEgY7BNu8FSZt6tajh89EAqJcZv2BIl6qKWRYR6cCUxd0q7pKE7DOKVPr
dWRP3T+e86RRNnU0RjuCRB2V9Y6vFMMdiRaB/YHZXA3DFEf3jLb2qMnckWdcgD/TjgxkoieCql+L
UaWUCIGNp4qhDjW6zLZM9HvZPOgUGpBuQ3i2A03Qwut9F4unqfdPAM+CK9yQ15Zjd0WZHQrLMR3x
9Zg81PYWqQVm4kcOX490UwZ27p8JXJvX/3EcVnI5+qRuVSdnpk1AVOXB00HNzTnhOJICLCVqBb9U
uLsj8Fef+tNAuiHTJAmyvHQsZKEX+2QBtEEeaK5tNQ1ISAMexPfizoLoiBnKe4scKVLhp/CRbC4F
+YxT00AbhqwPRGw7wN6z/ff7rDoE5licRGu/jKFETGhE1dEOpCJ6ElCTRsvrfuyAHPW3xelcDwl0
XDa89vT/Wd9tPThkwjjaOP8rlK6XdQx3n+EaCvHgzPepI/3iJktPmDDeX15FEhmU3bYvhOy7Gs4n
gcV/LKFXZ2cpwSJNXDR1ftNSf10G3e7LLX0gpUoIemgnkSmPKk9TrL/+4T1ohYSuYrTjcR3r1lqv
G6Qa4mTBBbY/9ZfNFHVGF3khxl/KTH+NRyYi6JgHydIAoHQHiG66PDUC1L+zDEuzBNRgEgJJGmRo
ZaWWsTS/Co2dszMgZaAqUk55TxRLGultQpatYc6VAu7v7KyhFkP5l2vtQhY/ZNiezqJTqGzr6OuD
YDVJDSOVj2GlspZPLg5HGCNM6b1vFwOVfmZlMb8PRZHe7YpY2Dhwaz6b29SL/Bdm8E3ib0vCkmb8
C3R2AaAO//4ikzgalbkMK04u6iKDCwr2kToKupo06FokGz/gYUtqMGZ9rCjIljv3bg09iQT4+bNA
pt1aFt1RGOVieqgxmmE+CVNN4bMuF+Far6XT4UwScyffE4d+ABjk1GNDVLykExSkoKi+M/yrz5gA
CZmSexl5d5Q2ArCpk7w+QvH84AjAvxfB1QFOF3T56Ple2lEUWGcmMw1LBBWwjH1rzEiGGE+fAvPu
A8CQAWTSAtltVr44yCOYtGDfsz3HU4MUmqbDfnOyKF2KRIMqA/qBy8wB+1zAA6vtbLvgT7Tsm08N
hsHygBoWbVxbE4O3P25mB/9hNeubvPiioM7oliHFR9ilznR9fm6qHTo1u4dv3nxI1KFdsyOf+SNk
ZTpuD2EXQvxvj+RCPUGZEA1mJfqHO8dohaU7stwHFPplZbDchN3YirDG2ncIhRnHUhY+31SmlnZO
sTuLK0eZnYZ2mSSJyUr86skYIveIK1OygGNzU2NCD61xLHbJPBmNP3hKTXtfSSdaWpVFhyd0kUJg
w1gVpQnswHQdN5tOBo3SeBHv9BcVmNaJT3N1ANyBZ2r8IipJJgmU+PYDDn0Rm9SaFVp33W2cmwPD
IJ85mf1x8rK6zbb+XW/C877KxgWClFg7eFPaPxPMv4S7VUfLGMeXzvA7beqUfc6bjqcsi4aXsCk2
4Etau/HvnSSkakMN+knuMZEEpCKn8cjSRA7pldB3SgRWQlKx3E5uqdrE+97W7/o21MHn88dmzYXa
apn7DeR+aFX68N/jiSHcZjwzUdPJdVgt3zHdSGy59+3iTBhoqt8VLbGzyH1jCQA+WN3J2zhHKbVd
0z6LeDm+Mol97ODiQCVRgFo8blaoaEpWvNA1tX5aWBK1gsfQ2D6itrjn2Fd654aUsa7WH+Dd6yDB
kmNtTDarwxKJUkexCkQNa3L4sXMIs7HdWzrqgNap+o28Ykrq9+h1bR51e7WIVsXMMcSpiPcf0Ilh
mVXD+bAEoEaYU6sxf9gz47Rqr1/WZWKcrf5e2vIabhGdV5oAl/2zQ9R7fJjp1uilqaIxQXoQoVjt
p0yUJ8kmbG9atzdxVL1nWs7Avk5tM8pb+eRVLnKs2r/GN5JROXTkCZ8u2S3/a74zdTMU5XBpVOgZ
0JXDf40s87kr83pY1HoN3LGf/7Ict1d1iSEajPFRl3l+gpRlq52+8y26AiSdKDvKFTchBvoKjP/J
GdbNbsm1ifduovCA5XLmhgk6ZAjRc5SGhtgGwBS9RwakDptIZd/nU5fPmYKxTyWjned18lxa10sf
iWLkeNCQcB9acmB6pISxnJn2q0oamJ08y7N+4LrFHrKezJ3mZgYcUilErxQDcbO07viZCFLDulQo
yUcoZCKkXMJDSS25XE7Jvo9cpwOGmqF7nhNzlwEZP+h0AIL9iQtMl8K48abEPOR8vTmO0mXFGlt4
I/GbKg1cnWLZjpeot0xxQXNSvfdN6a+uimh17Uj2/VbTD1SKmsRIa2C89rUj4MeQbDPFH83Y8w5p
ls/FljJYwDLAZsdfxrybNRM2kfr4aw6sEsccTGFVKj7FZIm1lO+MJuY/1Jh8HuPRjxPTWoWmfSLX
GgzzG+e39qXCwTJZcS+U0bE+h+lUZLX0OCzsSQj8pKgN61W4rfmBGzsErW/Gm90UkhVtr7tbNRwU
TtUNHjXkf4cynCmJSlujTxx7aHwuxGIZVbcGNvzbLCzsVmdufno02O9o7LLrSWQz9XZG26QaO10c
83ZxlO116upD9OTzO43HD3leDOmno5l9G7JtSRMdzpyoc32jLnjcBHxp0wDCemCC+kWutYgCbelJ
qs33AaurzoLd99TgFxj4KjDlxUcybTUZ+i+8uD47m8Zd2FOLrPEMl/RCE6RURuBIvJNt5ACAfrCd
tUOmSMT7okhvA/guYsQwON5sxA3tHFEs/Z8EnOwjVKUfkW8IAy0Q1LyKCfvUuT4tQjLL5a80ADZ7
jvaZ6UEF8HxbxWZiMVTHL4rSgby2SEFVuZFsoUcqqpfnkhPZWoDm0ljW2QyPqBr2e5DmHraTSIY0
hEk+GGf5WuczUq5CPlqp5LAQSrteEV6MIr/LK4TkSFjzP6pOMionM2uALgMBixES0F+bIrtOLou1
xzlA6ED/GmgDgJQ7xcgEcVc0oRgdINQElv4HamqXWgzcq5quh+6PFqu9Hiu0oOAa/LCUuE08fLW6
bKDvxA8Ow95g3OeXK9BNNlTHE+B0ujhSiCN0zoPUM/aR2H1VDr8U4cmlHWUkNVAXdBrplZEitla+
8Fi29Fbw1reCxgWOOGQYlxrBj4DthjHyrFrZCaAoLZZzSwB0oJ8AkMThiznHqWtLITpJxKJmKWdd
3vy6LRpLdbQg3GJ8OkKDNW140ONZazarghZAjVmpuAtHhaNsdpylnAmXkhRCTQtSiUcMGZIiyZtb
xWO+4eciRYRA/vQ4vn5QMB81tCHuVjmTRd3bxEnZvbSOneVNERPD+UySfT7iGQd4Eo7bV/W/3uA9
ANocCXRJKMZZQkVPm0LkBGDczOSuzPdaEgEyuF8C0Qj12lLlrgCGEcOPREN9HNf98TiwCyrH0Dqz
/yEKIN/T/r0DEmyK3w5rIYCxNgUC/UUDaF+9R9OTO/ou8BpdZwji0Eg2sEJBUcPA3pCX7x72K1GQ
ckT2PKn8DQpeBp5avShBFwhk7DIvoip4ddzxy0pVHLBk3+kr87tSC7FZ+a02cLIFS4TuIYO0Ra2M
X5rty9w9avq+gWqWU8XuohEdKeJ+r2hYs+QhqMA7tmtagrejhAudvs8dIkMOevPvEkg1LQ7kEdNa
bXPk8GJgBNDeaQvsyf1+mSjpkoK3QzjBFBwDEirfryi413OJJ/TVChjLRcbF2Po3oMcRHIrje4cS
5OAOFioH4InMk8QvNz+0RxNT2NrdA3Ls+83bwtPOp1WBMU0OQ7XV1q7Ax2FFCqgFlUpT2H0b+mL2
lWGp0iVuuO21PGTJuYNXr9xf4IOdRjAr7NPphM76Ebh2f2HROMZ3s/QhEmw/genjgdcvjTI/qtAW
bgeQrENdES4SCBmVSCkYGfLn9EmgUqcz1D5Qx4BfKYMICwz4Ledq/iG0kG5bhGa2fW8GLtvuLkZ4
5JxMIFfp1v+BH3WHNoNB4Ca0FodnDOKSYCJ0o/DgM+KcwOGQ2Q0MD7nIbNwx9l6an1kAhznl0UFR
j+buU6K0kWaHdB//vALlOtnvacTd7clugg+/34ubhQ2atkx8TViztuR12w5MreDRxYJ0wE18WM4T
yBERO7vz/1XeLPrN0ZENQ7+VBG/sxx0F2M8A5Bb3EaK4nu+oU2EKBUEJDEsYksVD5b0qhbUDiI9f
KkNcBs8ffOtgOpz/HHfNkf3VxKIhq1hFth0KiBwtKVZF8kM851wdpWhllbCu51SqsJF/qnvhio6N
0L8bINSpasJr2EC2/Wx2t2HYzEg6nGvvymJ/keh5dfcsAuIvsOvZJ7FC3xCrghzXjZ4QwPMt75e5
rfLxYNGGwLPECOnkEQteDDVkM/+R4vhPPEnRfj+/rbyuWYoaTA/FDq+zdsyOAcmSHi+5L3IDGTRg
+dYbzJsG9mKZNnZltyVAayRpkrzzUDnEpSWz2Snws3Y7Mgo+dW8k5TseFQYKF4Crp1QRWTaXGZBn
jwbtMvsw5OX/4zkgCArsPKH8ldVEP53Q/XKBkthpBtaEiXQIU9bn07QMoTWHZQHwlXWntGALxbh7
iZ4GH5MWKZMe012KAjyz76RlC1FBtjsvVSvqlt054QSUMl2eEbne+FhpuivEDbo+nEDh6RCB4TF2
DKbRadqu/qlaMKGl7kmk8KYHIVhJO4ApGZc2Z7hYEYk8QN0wBUrx+O/JIXPydV6jIjBlUPssa8dn
wujVFORecs99nLntJfY5ftEMRhJ1MPlYfwPat7Mh3iISkPIannnc/ahaeF70kQMWwsE75uIe1J9c
ScKK6L49KAwtNWyv2/GDGdgXUZlQnZR4Wj5JVu4NQzjZbBxYkMjH2MnHLI3sRnhxFZm9/GQz+MSO
7+YDeYrFZFYkha60XvBhKuCaIC+Y1ZfAKBXp8jxjzqpk3jrhMYLSafOxg6eYGzWHtMEAtX3pVP8G
FiQbab8efpQ9DTwF7fLb6gCvqlTvYpcZNpMJv2gxW8BjSj0j3afuQFnv+12a81G21XDO65oqdR6l
/PFQqJjE5uQ8eTh9mwoDXe2H4dGGSxcbJvf2Y3grSXBNu9cb1cpY9lgRusrrFy5dF2kUhtZ9iQFG
tcsgM9IfS2zBZzKj055xykYxB7YRqoGHEGppN7U7sFUQ4NpT81WcQg/Mr+TqCxL4ujrJTNqDbpDe
/ottCmnLSKE7ZKYQ1qaeM+BxPfcvxGvoKjzvZ7g4EM39lV52jI0lqAX2gyHIZEIbSRZ7+wLJsRHu
zHrnHFOeTKMZ2+DI4LJxvqm4pPJni/qof5/1W3miRmkFrbkItIc/a6UJZGHD6e/8vWn+86tR5fQL
73P+xu0/peMNgV1cDAjyj2CGAMux9dI/qbBU/Ic0oluiWPMo2GwuFej3N+RtzBPw0eC4ku6J4pdD
m1o1WakFopw37nQLAhb4Yw2P+8tTliIftYK74yj5Vg8fvvx8L1M3y7IJLEcb9SmdxgBqHiVIv5RE
mozi3HHK9NrqKHUJwAazPL/+qmE/1w/2l4PDLFse9urrAZvMBvNvoYeKiaVJMVUOpf9thjuGKOKM
2eAKjXNGTblhdCR9/dZbvD+RDjp2YDipjJA5AQ0RPifI8QIqLANhLmtV0sa151DFlsi2nYm/KC11
GvXFqlbbyK0hDeb2GCn1c4Zk1sSwn3e5oFWtL6eT2XewXxmLzdipO91j6YnICp4j3Sb+BvT3s7K0
xtYbz2+szYd4sQ70NPrxxFH7J81kUu8tiw9NwIVRG4chc8AN+glX/4Jms8tdDhSkd/3p6fmT/zWC
dpMMdHRCks7WAB9e+PIIH/gfqITq7D0pPgOHt4P310p6bvsD0uFbur+PhSC4kx3u9pb7QfBBFhqr
ItS8wCjEE4OaWJhnAOY7y0YZR1kC6q8lFJsWuqkRgHREos4mVbD+Cc3ZfP0FOjBXRMAzJRVkeSId
D9FOEUSaBu+oC46MaDiRcIhT1uoBiiheADDjPuTm9neSlH2Eu/jxhCNVyuG4zIgSygVmyw7ySQu4
ETdmU27GfGcuaja3D9hubo1HFY+PzkEBvO3VLjoSNCoGfDc23uLFZBMIswNZsHaIy50x9M66b2oQ
WKfuiP3hiTPr4BLx8tp5bb4INCmxqHbnlvTQAGtSDYkuqrbEaQoF0mQ4JS7BP/9Rz5Nhcj3yW44h
Awnq27wbI6GtnqkNdTU6JRDrr4jQPFy0Y3yCsAO7+SUyhs1r1/g8xyDzI+kty4p31GJ6m9mL1dso
MVQYztOYH8jutO1qCe2jUCGhb38B+omIRKKWM5/t6VIetI3EDE8cMs+I+DXGqbG56vhPb29EDh1L
Cph0fqnnNfnEG9wN0dzWX5TgDSDiUoD7ZcSaKqe4J0HnPjSEQMmuZAkinmB+JI6EnxDWSGxM5GVe
Ki+z6U4KAP2CrDKNxT7XTrR0M6EpRyDrJ46mx0sY+g5Vv1eymwN/Bd2hMRFY7rvsB7ehcOWfR/VW
tIU01Ywc3iwgj3KyunZJpkOYdo/3CBkzS1ytLIOFzx2oa+tlKt1fTdg1lIoK73EIqrYlhr9SZ2aV
8PIAAMEBgvdaVFmXfilvE8IZWNzmK0T20FlvSpTpVnCEqiqglFRV9qLGxy5f6i5yiKLfxnd9EAW9
DgcYefZFUEle91nSVh32pW8En4msSV6+0RzYjPtGgxqfGe7xBd4g4pHGDfl4kk2yX3HLOTCYfuhu
1a13Lt+0cLOw4Y9P+a95T8/tlrzk5FjKXu/8vs+L7bRgZJEAEl4RflV6fDYTge4YwdJFvdkt7EDA
NwLtBI+XO+rniMsQzjZsFFCs2D1o/RNa/IoGlr+iO207jRuMiCX0zq5rOgxGlI7fOgcCErgh+pAy
efpRwc+njf+XTK2uKw+3W/94C3dc00JYMSexyxyuX0LVoROWm6QS+rJmL3Pa8H9QEtBCCw9Ia+Kq
qwj6OomaJAv/Bsf4E7IQdU1sTvcFe1Syggl7hZsYjEDq0yv+M6sEGO5PPW4YARTPF2ZuBSFzqUDX
c7HaEuPbTI9bmyqiof2zFQC2HObQMdzEpFCr04TJj+CJM27EL4fo2qws2kBuaawt7X933HoKA8AW
50eJOLE8TjKYIwIW69ndaYJyVANiV8+NAwMB45pGzatxagKpAihI8Yhcxp0t3c0n/LkVc6Wgi2O3
5vrjF9JMxKJyCdfhPkigK00tCadKx92gQKrJRub9wYItEcoRDv15jXqIVP8m8pidSvWX+n+20bNT
Lv+W/AbMB3lr6T1juFca/+Wu6BQ0jhtoliKuwxsoESp3179Yb9UzH8CeRM6YHjxOWxm2Ym6tc/Qe
wIw7hbsQtKN1GfYIFA2RYzRY3dhEibaALGind85DCirHlxmtuj24eCTlbQeJ+9APkufNnlBqaCdP
3ba4vJGwLgR9zazxdzf9jU4ws5K+rO/ng41dpVgbKUqbBQs1ndtxtKgT7v+W7CAueMsxxEp6iQlc
NFLSKHDuRZ+Q93WpA1wcLWZtsZiHauET7W3p5jyNfMqsZBdIk2jv8POBTueEiSzKeeC6IUdOQP/K
QzS8JEzHHFRbMSQzZBGHOvGL97uKdj6xy3VXc09M51INuAhlRmdR0iTxozYFm5Zp7domt3PFMzIg
woNuvEXFm0kjrucCqvrX7mhQkAm5fTuTu+GVI1WGdR/StmR2xO/SkfYlJ7WDE9pC23E5mAvrc2TC
vzGGftGiol50aGwuGWoqegBz7pHvzZNxjLlindBgBMPEZI1E+S5f+E8uD2bdq5zfE3Gxpj56q4ou
EfqTM0poajQxcxPR8mddC+mpFqhA/Q9FRgTWLgf4vKK5r3y1KMHCPWIKTxsH6IOW1Nov0r3HAI5i
hSSrzLkbHWln1kSdarkyw3r2OjtBDm3psvnls4oVlJ1WiniKCeZyT3+e4znADqp4PX5cs0TyhnyK
7FcHRiywk97AuHoxVYVfwxed7Ml1qv1igxT9yqoxy1C/xUWvFfjFNkRNdzESduK2/YahAFyEbYd9
AUm5KH3AFUhic0baCb0TDp5EURhH+9KKtBtJXrOm2Hi6mms3z5VhrtIVL8OfBTw1DBBPmVwl5Ifv
A02E1+hYBchpkFbm/CEXpD+P1Gb14XE2Gm1LQ6pOw9dS1FAs5RQcC+QNHqYHdRKNHF3/G13RRlpX
PxwpEh7nqb6h34/nHjzBBg6cKRnJQwQkGpvnXJb93Yx8iI6ETPRZuTQGyKIJ7l63pkWPAHF7uWvi
oYmfHWH6oYAbp2kdEERWJUSz1mi6GBNN0D7hJhWQetBYwfAeDYKlX1W22G+bSmKnzZ1q1J7v3+so
veiR7n4NFOVkYwZgBIhesvMcTzn4+5k3haDbJSNsqcVZ0motC3TD0JieVfOAn0z0tE13Kt+O4pRV
5lmdEBbiUAg5wK59dJX+TIG49baTqd4AdYiURZtYcqg6Kj/juAzUTjUvRN3Kz3ct9VW7OCLHwEje
bdS4FNzelF5f2JXBUAcuaBc86+WTdJX7N4bO7D9TTa2dE6VIlACUE2zH7nn3D7QOKY4jY/oV7s/s
ss7Ru2my+B/1rFdcw9oThFt/JMtLcg6DxW2FKJ6d6gziKGCE6IkMedNUAATyQ7xnMAtsmlMsPpvn
AOrVC/536v9kA7591o+FtQnCCQ6nNF9I/mjEPl3uaqX3lO6hG9nP48DSY4MIqnoN6oGWtI9niuTx
414Qoloe1tVCMvhnN6ELwV0LZ6q6D90N9I8m9oJ2VoiMUooOn9JGSZKYxPLYmQsCCTtlog+Ut4rb
gv7d5FwV2B2QtU7f41CJN7j/AiH3xuHIRIbiBLWhopde4VSqWFFAqiVuCRP6pjGIqcRWkCMYaj0T
Aw9WzGxXR2Eq4DsZycV/fu+o65yg7Oc+2cQMgdksuq7jM0aNMWC9d+kfJePaDTttYsmr6A5d7FHo
3F4qBEloiLn61cgUej6qxx5l//XqJ0WfoMRPdrVbXoBWCTFqlxcyBRbp9w/6Et3lJ1FPlRyQjHsT
jiSN20s1+g94xZLk2XZIBLQJ9FSTzSmo+fzLp5qTigmo2M7Tb+L4Ji6ZKE/HF/J+i+/5QJVPTz6R
XLRElksYoowSxwZvS/GroPiChfRLHV6GvefNRQt5+CuaIIuGKdSSKiR4UlrykpIT1z8lOgk7RoIY
/u1c/dUxPkyPTkb7bYHQf3LCATe5GrVwdph3s6xrufas1h+fskM+7eypstkBL8r3zNMjSimQd+02
mzQKEVk5BXnLslxbBXnk8A7X/tee9MN0Y1Axu7e485O1CR64o0733dtFyfbnR19M2ZtXFQtHY+M5
JBKevAzH6xhtVGNTEPZYd460KiWmJejyYe/Y5jUeyh+NK9pIMjCQjUVODff2fMZCV1tC0qbOtRTp
uRZkpGmcp7WzB112M0JVrTFmtyg8509KJ+UkcgnpeL3zdbF7kJ+oVV9wBGyNPb+qmhgVlTLH8OSL
93O996P7UjJbNjQKX5L+k/lb4/YFjguUmW3PUWlLEjUGi9FFZ8utWgrx5/wBoBjaR+X50lBe5Zz/
u/ofX0kjaoJn8mc/lk58++YP3jUTnu+2335T/RE4rShKOjjYHb3nY1JMUCdIj9AKMAlfI+J0aiJX
Awx2rgDL7BRfs7qRPDNGgAofx6x4jWfuBnEUJhe8Rc8E+Y5bQaXk1GdZPBuHWyW383YySnDnSM2d
xU/yEAFCSdLiHdAACjaLggO4sfECxZEujIwY06y+ne9YfSmlVhygFUYH+UtkW0rRJcmcq/yTL6FG
S9fyvE0noVi8sYDSYSoAkqk7lF+2ZO4uLaNCUSBErtAGzLjXM1/T7XfzmF229Kl5lOD7CQanFKsz
owzHppQBZoo6DU2d7qMke9Vp2YYLP40DHNGHh78FBpx4FHT8p+0DMb0UAMvwCVHofF/4nUrt4Ho7
cnCoSCKRePXHtIHyf12YhIW50nwT4thpqLsoSn6j9WnvZxYBkbLrIEgx+WbTmGz24A6DyQXCu49+
8kgWUvGlhaemAT6mv3GX/xNX+ZV4m+Wn5yoGbgAEx4nArO9Isy6pcgtqcpWYs0otVU4ngwBkqC9E
uDJPB+453opWZpQWbZdQRH68pfokfICWXIuMjVD7+hqPFYfGiYqM5dk84JeOJrEefA3HJ/ul56YW
1wgeWb/JI2p0fFMbJJxzNT5ffhjj1dlMmfOBrpjd45hw8SZViMFUQZl0JQ0GpfmI9ffNjZpJzN9m
3BytygmkA3pVQ3KyUBO+kw6VhuCzhwjOHOXgLJ7ONTSccc8NxkPoiG5dddBvGW0elIDgFyX3J4hu
aSha4iIYrZ/UiIYF5LSPEV8dFpVFx4VZ0EXgg4/VWqEjWN9Xe7awb3/hT9O8TFVhjVpMK1WoA6sg
mA+9lJ8xx1a2f+dDQR8zza/qTxgTry38Q9Klnx3TYox3cz2mGIHc3CMlyvHPBwtsOMg9sVvDRsFF
GgAaMrd76V83PZbcy0cuYyaQyxu9VwSBSb+oNXL5QsIU6FYrxgfAYNueCmuvRMmuSOWUDEgw9fw2
7hth2u32Glyte9/JWIn8n09tnDcBo0pIkyDP8byJZMz/jW/gXjP0JhK0DPo8uGB8TCt5TvlO/Kl0
YqH45j/8R58I3ONpAtfWfKIhcHdH8FdaTZIuaaDipT5aE2K2jhLDhW0730CC8yy3bIwuvQIEIc4g
JvWnVoCAcsCZeCo2/dINGnS3ZIJV9LO2r50o+OuBDg04lcJ1L5nwXcftYKT8JGdH8aQ/dVjy6dQ4
wKhJ1yK5lgkCbWG8CMn5XJvs5LBAX4cIFa4gUDWq/PESMthZT43XgGXNPtHvK5sXwSxWQKEpd+iH
m8JvTQAYIViFsL6BnMfuDsuNi2fiyWVrvGqr0aZASHG9B29/0mp7bslV+f+d+cTB/H3qFP1nJg2H
22Tbr4mCTB+GnTo953uAFhI431NRra+4Y0hHWu49ciXZm1iu+uH12oJrzEtAaCvUtoZMtFZCofE0
w2vZB69zwfcWu1HAjJ6LJmzl8RNw4ONfQcgKGeFkTmEklR2P3rq/AvvaPipBPxNXPVBpItcBpiAX
KEuEeHWUCaPkqcyeZpkUoclWX+zrZ/Cm8DUiO0Y4578c7o2ndrDFQH0YjWNef8RE5ysNWXS0XLf6
hjYCN79U354TR30nwlihPMkCbnnZ0YQ9s9Aq518lcJwxk6NGAihsgIOb84ninXDXs+RU0dPOHjkW
LwQDc85+H6Noc475iKkTSmIRPs3Y5YC5MOv79wZel4JnrovXuG9pqMuSZgqBxsttIBNhG177VXKn
eOWvtU45P0QopYBluDL++pwrKWKkvkpp7OExZIqwxih8hwyzJDHti81K2ojxnxUSSlpWJIoAEuYn
AmRzsoPqVSSqiPWZeb0lqcBdeaErvPj3tT7gK2RZrtBBHlFUi2DRAlB5VrKbpS3AvBVgIWFMcJMi
8L8D8VSTnRFAKHZgDOoGXbpLAGDddqQG3YR+4XhPnffw89dRD/FoTBBC3FcfEhpN5SOWmecLPQT9
A88hqm/+bdLNwlj6md1cfroZ8hrSkMuJzxg+oVUUK7Tj9Q9yEcPMsdPHTGE2NcIREOD5z7z2CRYG
mTcjEBEOUFCIplQojwblTuzy7jhB2gRbgBjudqCJjQL5rax0fhlYbPc164XJjecmOfIcgCSSC5w1
Aa5jUXBB7jxfU3phU3Gp4majJNRmGJKs/TWgkfNmk0dpIWUFNpB5o45Bec1xFjkicD/P/o7ubSx+
3P5cTX2vQrDCRfQ1cBirRWxmyg2OSjn/4+AXAN/+bvDqi4ihvBveYS2oSKn+FKtWcuSAFaPLRwHz
tZdHgIkzgo9l5b4zbSUPd/3BFKwk2GQUyAL9WFzU4CesbgK0TeO0RGcUV8SFAmQjCIj58zmNG6s1
G2CoFbH39tRPQTqJQdEVn/WPdZwIcptGnu5gz0Dae6D2H8Ln+VNaH+m5bAA+7oq/r8QGPma2xV72
uh5/HrNeqkBa91LltVzQ8aYSzhqOygVDEIsEE02Pg7PQJhwPZm0VKn7672/kjq/yttkLxnB6CD50
2L4+w4bZQk6qrffw2+ktYd9OzByWFfNiorZXDHAz86zhvZ/+ic7P+DN6Sgr98xbequxF0QnVBIwN
gCpaB2QEYwJSdOsD3PXpnRrdvbLhirwUuIH9jUJK6GBbrSKMjAFBbp0sbYiavqrMES6KGBLOJrSa
kJ8E3EuDSQnSPOdamvECCLJa458C9JDmL17rZcfqT3qM/EqU7SNu4kyaMtzK4gS86Huoe5vL8eZL
h63U+0wNnr9eZ+kRJ5vOUhuT8TDOiyGPo8B42ed0HbCwKWUQdTJp0LVndBkK15SGO85zEQqlmxjI
uJN+B5La/KQpMsJPyD1YMwpzwVrpG3sOnrkRWMIr11XQb+cbuDrOHdDQHnDEcKpPsFiA9NxeXLnq
qjw24RacdBhxhq8FDSgvQRyLQV7T+DvJFa+BOCMHNPUjy1iVxJTYp0TzA48mJLDEbVPFjFAjFeOs
JcioDpCLLvMSo/ETVCkdb8f/KN6kxbKh/SztUQOw/jqH9ULhuQCymb36Ki7GgMljuh4IY+s3AmZF
QehRtkk5fcoUWENGN8VYWWqrsqJ15yiUjkd8N3wj86yhSY+nIwe07bGkZUfD6lO6G3XPGe9avBbX
uxMTyIwGH6hoqB+6B6gFAuIpz3e2K1NogmMPAFI6BsQpeh0c2jWYb7SpmfZCtvZ/u+KMSchc0XjS
GI4aGe7B1u69/Ov/WXPRwdFQVPBAkjKfi5jd+W2XoaodZKq11zYBMx9pPXd3JiF3dvGfG4wUentX
5PjoFbcbKSM/WK7Wiwx0IbuwtVTCBXKzEWXuEWdYun+JrDQLFi6Z5FXpNjLYsExAQ9EJHcOaIy6X
xq3K8D8i9Hp+9IgWnmFq42LzFmioviQQV0X49+QMcj14TQ5stOlyQ697qOCXMQQ2ci3hI81mYNHf
AIHcKYRMNtOQzCogEI+OR/B++iQlZy84Q0Z1d7hzG3j5yHwUbpMoTAsYU4vpiVcHP9XOp+UdyePl
c/uhqicZ9PE1O+NlNJy4DBeIzc7TvLTP6ZRnqTUOwz7UL14WpUVg7ticjO3iB8SCmSAYlZwWtOo0
AwsBbYiZ5eJQwyVSkeifAHdy+s1SKHv3+rO9Zx08haxPX9ZKGkqPuGaxS+C7ssWFXlE5ctmNGZ1L
nqHRXSO4tKYnvWFs9lmYzNqe6wMw594pl+v7lI138gkqiyPr2fHnCSKKGISJ7Cm3NuLQlZBeq0jL
Mvt1t8U80Xtm0NEi4jYcr4rTq5njymYrhSL1FmkQVxgcvNio6+WK6/l7Ihx0NJXEiEf4c0d6vM8J
/krMXiMEVTDLznR4spJU2nA+ptMypC3ZjETrj1LREBl/EbabdWWKsSRqC2IvvgoMZMAKCwBYZ+3p
XIzF1JUHyo03raQE2lpuEyWp8Bq4AkK16YE7KmpF2bUjffg8VMTOMu4y3xAQRcIhGteZbdmQayYp
GhCoD/qyLtvyTrUiLKbVv1b9Q9kp5xBvzb6Q0xZdLqSwLPhlu19gkEbSUeqx4x9aIiD89N/S28/h
w2TRs8agIu3zqoZtClPKPa4u7/pgIFwJ/hc3f6/qYvW4qPJU02Zzn+KQQ5u+p219cWhKqnxKLPLy
xx/22+RH6DPSNHvPjeeAbeNCNj4fb65CC//YWmhCyWu4MYW164iGS2j2JI9u6AG4qb8/1XM1RGPX
VIiHdgsY4ikfP21zz64loD2nCsLMBo/QMnS1QVFJ2L6ysxpxqbYsb3RkAM6XYS8EU1yejAU0aZZa
9JYhvEBa4w97U2TfZLLT6zipK1Mv22Q2WLHr7roVu5sL8pPAA5wK3oWqw9e+qDD/RYHAnOfR+bU1
cfPvEYwx2oczOQHyktRs2oT3hdzcOVCOHp5FyxDYlha8+r61dewYGB0lonkUtiHRxnbBatyRngTU
qI20PEmdsVvH1eoU4TDuKdaqrw7u8Z6V/gGXGEVuaFG/0fRNdvMq4AA+auhW7qqxBzqmCbWZxRIU
1I9V9lZWcgyxQ1876ePTeg1egGRGQRaWtjuqt94VCjiKJbs0K5jwuoQq0T0mp9m1i2J/gXimbxLv
m8v2LiLg0XXOqSfWdkttsxaVmJJTR4iIR7h8jHL7ZlfFR6enamvkY+lXQsZ0YpYLhKOYM6rjUrHR
T9Ql1GF1NdswjgMe2ELGd/KVFwNidAwmlrI8AvXnCLjG6O65IKmFNRFAmPVVboiSdyBO/cnirCcR
NeZwKw0ankBsfLkzC4QeW36w60WtbYsqxswap6T7gq5gt5FtDT6SVXPTPRaAdmNVVtX7qTPR8Hmu
hSoReErWH0mxuTsSHIlr3XzPVQhWxgr9aPDflYHfOMqzQWfUpQbCzSjc7BjJ4K2IK0Ji7NNQX5j8
j8WRFst3p9Av35r37RntwJk05bXnNZeIbOA4HmFl+8pjGV/wcgmZZh6SI4JuPwtK8nsXhXjlDUkt
LnQq04LLEjwMkx6ghWQM61vit/XCIEjFEoOWUpQvQPOABY0JtsdZfS+ONqVmJ5c9arqFhsA0NsRU
ozfNJSEfpnG5qRRdhuT07KmEmcK+pXTOil4WCpa25j2o3ysX9kkS81rG789cEA50z9Mvg34jgcIb
WCOhYU7DKbmfzT93O9+v5tuS6Mt46mp9do/8RqAGEwmx54wYhige6yo16Vj2eUrsKfs6sTVTd5Uw
2c7HvrA8wFT6ONj8UQWAcBSyX3Q/wFzrizRWndCHez1L0TV9PsDmg2V/Bkk8REMZVAyh9oGL6SbN
CMx7wUNeke1mhqCDqb1OMCCmvTgS9ZTfPJX0rOAYdbdbaOCa/qXl1PFV0JWD98kWozhUzZ5oiMgq
1YjY9mPuBQ6S3bC64nZ9vbI3LTxXs5v2z4pXpxB851mPIGtU4wz2vFDL+TexOT0jHwymkpee9S7b
hX0FomF8aC3kmKtphVc6B0SnUfTZfr3qaFKeaEygv59+E7C0C4BVHuwBrIuXN+1VLWO3Y9Nl0Bf0
0bLepKG5P2OUSQsOlpXmwA+fMMTIk5oEtGK9PH8ejPtlx9TKBtY4OLpwahcmW2D2jpnWYOZOznOP
z8YAW3otur/TR2EUD5HyoQqwXyi1LpXjy36fL8oQ+NY+EbmVuxOlpk/a/SlA2+6xWc36A9fXL1H/
LacNcShQ+vY1A8gMfg2jsuPhaRnEc4ZlEKXgPaceeGUyGFfw8d6Ow0wIrbdg43x2VtLcaKpGafjY
jl4x++fUodrMXpH5EhMA5L/XngIF3SDb1bt9V78WAYpYm5WfMeswYl+Z8lAd0BphkD6R5AvIrN/+
L/PihGSP0tcBXJXixpLup7yn4ONKzjpO23riKMYnFpQtALz4F3VogUInfAjPQEhsAZuZHzW62f3c
oKBr6t1lg6TFIxXH0vL79xI18ZId8Fu7BMddjwBt6RV0Nx07XssWkVcFwsTYuFfBMU++HltInHNZ
kqKkkDm0HU89sctKWY/FUUjoZ7x+4Bjpkxia6Jq/WGdm40F1tn4a2mHMnDmfsZhPccxhoNpMKCMT
uMZ5/EAe9znLDySucKKFGGadcDXIFwHiPwl/fFDE+9ITVPpOEiSL8IzGlzsNPQdWNA7uQkmqIt+F
N6VCI6E8O9NDntoJZKmqO3uhjgkAoeu9mwkkF4cCTy8sc0cv3lrGxJX/i8Ux/lYI9RIh2AKx2PLw
HturL9tvT/1R2seIA+Sob9AUhyAAOO2DC+DG5pzCnFy7Iqr3qdJuU5II67Jy7nCYnJLdcnpq/E+z
IvUwmBF0sJBE6OUGVq8uiKQfSLjDXTHNmwoJ9QuxG3Q3IHW9pQBDrAGiXvaU8fxNXwLu5z4/JnB4
V50/ATcSsyR3/OQFMZ4r8Ew2t0taSMgPOk/iTCVxfbvXuiNeWx06xoBJdBqMdpux07FbcZXGXZRr
5JFxmVqg+RqW2G3avjZccc0F8xBXc7tK/rQlqukY3GfWpyepwMX1xwBiK+gUoNpJ6pdzXUToIM/q
4s7VEtKIrbnRjLKw3rMHn5gCCvBkzwCLqe/ic08vWQSIKYfKZGY7kgskU/NjxeINr/NfuLOnbm+N
8IvQWnr5FbFL/Odthac1CTN8yHn4DSK4qqsxNKH4ALWRda2ktV3qogCkX0ANpkXHEb6Mf65ODcUd
/3qFJfuie/fyaoNybZYgNTBxR54lXSbJaexFf1WWpwlj5CI76YEVU9Jpr9y1seqrLU9gXwaBfuqF
3+JyQA1C6bRAGJdPaUsM/hEglIg/cMmfZQoIVZZYio41H5mdHubyng8zsu+rEBSd6lIJARyNNO+k
hqlA+PacVaJZ7WbMdM8vos4nOhvrA3a3OEvY4rL6gdqN2d7vI0WoFDXjxjs5T4fH9gS8XNv4OxTE
udf26zFV0SSmb6NDlOzZTf7J4mpI6n1KvICZvpQfTggKUHtuSAtFZWrih/lv5GgNAUJ85n+lzhT7
m2UNnFyb9EdpxkbZd6uEjiBY24wRNs8sueFO0aXCxX5WdRjFWuFu0mwnEI9CUHYUHAPlTtjfNUzk
QJqlDrc2/drQ3co7UBkzEROgj58zUUK0yjPj8DLTc9Fl5RocF4l15hFOU2MDspRC1GyyuIOsKLyj
E5GO7LVsVTku53r0yIfgEiLm7ntQ/G4zyiNmH1NrBEU59Di7BEUH0HxBpVvJVtKww6Hub2bsJDqE
94OCkNmlgy/PDRa7RmHm5y3zTbU/AtL6XtfZfY6d+jdYGHNqYtmpEvP+vswjdrc+ZisUBVSrPuLr
kQI3vZEq75fLsaQevIUkuZogONX12wMKdRWTj2hnNAIl6Fp01Q4jPKJko1W/k8TY+k26x73tyv4H
NBhYKLGrGCTQwsCi9AgcaINJ0/dIegEgf2LsgwTHxiGGHWN1jKGtzRqbmojbeGU9MifEaJaktaiE
sZ/WnqtLa20MssUerI+SNKASgWiu2mVhqziDvk7OLd4gYSdvTGpET/YJRKJvDoMW/dpRck55KriT
8D2INFwqhYAv3zsl4xemmx6TPQ5D7Mxl1DzHro6cFD/tyCXNuGnen3+j8ut9IJyjzkrBsrFxAj7G
AMPWmGHL1i0SyCwnvOsAqI7Y+pigaKW1VcFMrc5r+m+esJK+VZq2dePs9wPygsDLn5q28+ZdZ4iA
vbSXzQHCA6alpg+ZLRQi2urn8gGIwuX789dnGpJD5VJDhcJ5fKVRsVL18tsSHKOf7g1i2USKUP8I
oAeSt9RyZOzMdThwM6Dx0hzcOsLYXs2u1n5avHYatgTpFuS6o7RiJ1/UTQKwTpLISotT6lTp4S3R
0RoNm1YX3BAkF8apaim/Y7ARjO+gcRjNQe8c5FCiVkfRijgrGWwkRgvlB1yKMrfCrKncF93oHHoR
EjaezoEKvWDWjQiz309woPz2BVmYfRIBn9Kd9fEk/fTZea/vtNI5MSeO9d/FWPNDXWoxW8OO2r1r
e0nWYZ1VL6XCiIWi41949P0etNfDUzs2eQVhLmrKoxDdl+5eGTe/eQ+OPv3KphVQczZyalwrRhM6
qcnyJD+NK/6qjO+IN6porRzgfKykRus/iaRmnRMeiGo+TIT+Or/i6UjJhVE1OmkjJZT0sWkDgZc1
OGKyk9vAsHOoLl/rzyuI7eEsW3PCTVD11W3+gAlbDK0ucdhSb04i15vZ89Q1nCeVY93Hsrggvmsd
jlqnDIezcO5PVOwleTtLGWw17REe6+8Dlxo1Wdw8Grb5xq3sdSUKCMqMHtq0CI6zeWv8DdORnsiC
sRAB6tcGDK0ylE+Ej1lI0mBsaYeVLrNG16AKBxM88RQb4wviR27eRjlm6kXKdxoNMsrX7k3OiNiM
elWSyqTp22Ht+PwH6O/0kMraR1QAORDb5KJSHb2UmvUAtmA1hPGKfXZqFB8X9+sz5ky0pfyQBckI
5IYjGnrJQfGVO7lk6lo4KlQQS1a5BthNYibQHVi10AW1YaiBSABUSsLfA72ss9WxpV2wKfuR8K1N
3+Pa1UTZwGvJzLrUWwZ4bcNR7OQJjnrM/VajfRf3y8NqKx7rhc6Py+YckecRbreJUdUyXJQoeScX
5Utfij2EVvcHLTHyBeSXXTbDX3NyikT2IFUFgKQOYk1NPcVzg+O2HnYA+iAzt8Paa9xFayP/vQ+9
QHItavU61564c+C1u/FWDE1lIkyRYsjcnCcsltMqYbo7fB5VMZ8Piyu0TbRw9CXHhkO9zCNiuRo5
qjizxN5ctLCSGI8jR0o/4xEnvan9aKT/BI2bB0HsTdLl3Q36TW47UdUt/FV6ejr4bkCMBWE+Jrmk
npHpbZ0oHfm6ARxYAEZSDjrYIylQSmJZm7CSYn1r3v2E4gn3MywaOX7Jw2r6gPfaIQq/IBYKxSol
VlpaVvqPI0AKlvUVyX5dI6oVBm7g4H++xPS6MxuyYARvqQ30HPA5FT+orneIWulEloyUgw/MKHND
/cYGou3zZYGLqhudgdhuRLxe3DK/bGlFc03+K/9tmEGGZsxOiVxf5F+k83ChnvA4Vx7/GJxtB3Z+
67Fvbh69JUWwPWXUI8XGNpCpOU4576AAdNXW6riuF/LSoI/W1fFzHZ7NC/S6uw7sejpJcwOBNGDU
tk1tANtvVaodXyFric45+aiGN2AT9QDeCR3w3z7JYCqeoNiJdQ5Ru7mBa4VyQjMbGC+TfNcINsuL
DnfjjsH0vxq1wXibALJO748/JfmOMaP9JdGdN3Wca2spbQKGPerTfP9owUUPFaocxsJGx3txz2MI
g20c/2VzLhqvztEbEjYFtaljmefygBOb9cKf+ORCTRwHBielQm83v2xMG2+cYp1aJJqMRY5RuPSM
QMlTnNpJDIPSz/NIbruEjZaUpWmH/1XqTa9Y4fQ8vbZL9zaeRyau4zzWk7LC1Yh/D5lYrlK3zm8P
B9sX0ZkxEEjrco+5jzi7VtVktsHkjTOGlsYjx+CHA5PEhlD4lR2/3b2lwflQHUiNJy4cvOQhC2dj
o0zMUWMfGen5MXzakak0WaSof+AbBMAlIjc30dAx1rtC3sCEgxPDWlgjWx3pZjDAFKcSE9DK8kmT
VOsE+TWE4wNOD4feiYxOFyowlQgelwKK+53f+G6MeC75d2dYjjIs2FsywcD9zCsKNg2pdrcz2viC
kFoV94JlTAouM+Gc9Df+9SIMOY60ERzQ84vmsgph0P31zr5AlX4BqIStIfAeagXg19WRC0ZndGqk
JwyNF+Ye6kNQpjL371r6fXGGUfHAUVFd2U2iAIAujAHLMLEStrxJDs5gwhP/mS08smtBW/Ehg7tj
j1ft/amgQmDrF0EYTTXwpFLE49/Z670DpAsnU40Cw3qOwfzU94w9fbcjsARRLV7slmfQ9qmf1KnY
LyAzdYK4B9IAjJjlT6DrPv7Smg2X5/ENX0KgVh2KnZ3jLB4FfvOKHxxjWcVU0Tt2DsnyRxefuz7F
Re9PowutMPgK0sXDkX1PEuCIayA5uDTL+ryqRPqKqqExt06wjzpJ/V76p7wKKey5ol83v5pahRc5
DN4/UVHLBDj9gXGvOYsqeOdQm05/IkRjh7K8GID5E5Rwj7aDH7GiN0z/049wV0eZQJUuJ44lrv6+
HnjyunhuOU2DYvLRbVx0pOS7XmCgdApPCSZl1vvkw68WRaQWBw8ha4wXJ/noryFkBXr16gztHGe6
0m9qhaQAPXEqk10RA4IXJv5VuNcfHIZQT+cpUcT4xHg1OWGFWoZ5d4OaVn9xqT5MGZ+AJJtBs6ms
3GxvT+1SBfx2e7cNgBKvvDsQE6VvtA5mbiF8KcLTR5BMmNHW/fVBaEPAdoRBNFnGXPWIt2Papeag
LFMbHuEhkFXiY0HS6MwuKNHRfM9who3ajaKBAd2z0tyzAnHQlDL/w/y4lAaIBwuyKWV+q/DhJf6z
Q1Kibh01dcBN7mp3BEI89ZDGTqfW+/aLar/WnO6tNMqGRsJrTLKf20XXxljvIXG2y42illPs+Epg
TSz7CTwQuUuZUjnYwJeKBtdvcaJw3cnE+E1tsw0z5HZD3CyRRe/52yGfTXOLC7o+0MJpZ5F+iRp3
kpOGX1eWXQ/ZJtSSBg+0YJ1pzgROMmwza7tOt/ATIOAWcII4W0EL5O0Cq1RULtwCy/Son8Hs8Z02
67ntx9vxWcZqtokiRU2l6PdVpcdlcRMGBmqwIVOfxIb2RPOrmw1yywn6JFbXvKcSsnme5hY+BRwc
uhHGEUyXihTEwVzff9cPArLMdF9hz4lhQ91qvMrVjdxFLAY5UJFc6eOb4qqTlvTtlEs5q09rKJa2
ipNWRl4F+/ueJhkBkyQHxO4iPKxvsmxfuc2lB+JZxITOIZgghvAu1nm8YV3C9MhZ+0Z5UAOdPfoH
4e9KN5JG+vji8/otbo7Uxo3Ud7zu72iAa9Eu/XIV/e6QWXFmh3KIhrkYKA4RcR+ujM+vyLSpUn+Y
Tx0yzumEQ5mar6mR8BJA69DfHkPTPNs/xpWOjvzgdWA3gDdpXlNUjo8cMYn9FtDLkWtBvJT8fQ6l
krXMtHaDwHIeyKqdCXd26XalEkDZa6oGUUJWNs7YAttQdLNPm3mWWhLw1NpWynt1Bk0+OJNQ2waQ
hvGZZffHACi6K3qjNWPM2gF57gqRm890T0SsNk0SI9hAJZUpd3FxWzOX18inLmqLMasN4cRhFn3I
4G/xp1dVaG9+TzriNMfD225UUs9UDdM8AWA9c213GouCtP/uYHPp31ugIOp4fyMnFJAPhupLYAvS
MB9+hh+0lpcvjzxKNeiaZ87dRR7FdDJCF8aCTNUrpRK2GQR2XmhP8QEH2mRUShMN+ASQ3PjCW2hi
cc8y+mf2pnt4+AJMGxIxhvr1GtRwuZPqV3cUIdu5EjNdBGQbjx6qvq7nIolwxINbthZkvz6aFVyH
7sgnYGfOpGs6tmQujY0JwXsXjv8BuJmtcKL3B80VvoyJRcjraYFhWs3TiYQtZadBE4jIQ1wFmazu
bhIW4VUWrma0tABZAVpi6mIiX++uyq6bNqxA2F5W1Zkpet6gZ4ABaD1df6vSg9N7Qy+tvmDWGjkK
nLA1yiHtQLjac9e3P0KCMgfMTA2jTsQVXL5p8C257PntXAxGpfj78Lkh58oprB6zJSDTtHKEJhgP
DBHEcUKxr+hemqJysmEneJm3ptI6QTCxlBZGZU6lodcgnGML1zoxIXyA/KzIXh9kPrwh3fFgbVeo
DZeNUKkuzuQYFuQoDSQsb+BGGOwA7Uf1otwRYHhpmrmZT+T5wS6CM1Yq4TbFRlC9KEnMtCdZxxEO
5ULKBi4LbI968rrqTF10TZJ9VB3+fPBZ68/p4/afMND2kOnqK7HmMpsiHEfMgj5CN/e0797dZtIT
E7lHHnYyPhKNePT8OD5qiXECeP0N8RIA+GEi2u4xCcwGkMIku0EtD3JO4m5vZCg29QI5OxI74I/5
/lBv3o8LXx0ahw5TJIHpZpKavXipypytR8rks5iN1/EQVCQspTCOte8ExvHp6NpOZyOGyfnRTsbE
Qa5M1uHxKioY/55E2PQRQpTE3tsJwXBgIJQamh/RxOxtdf6U+l5PxYCsmlp2wmEQnjZbfZPrTCKx
BCSpxg/iQASUGCZvbTue82jxQ6Bfosk2NcqED7SN2Z9woW0ALeALcmTGqUpb1xmuabkrqpkD7Pb2
TswiFPCQEwnHvxkb4BxEgMrRaTCQ+Q4nIt0amszp/Skqu98/DWkGWym9xP+ywnm+2fLXZgfhFE1F
qVySLw9sz3ieEigfpMfJxQPjCqLGPcB5d5rmtBaT+3siIK/pHB4Bn3niYTSfKTV6U4eA+mTabbtd
IjvLGL/Q6aAAuV5eSsbHKyI0qBu0zq1TmLyWFOv2KW2cr/1N3RrhUsSJ8sqUlIeHnu9SxebDCNwT
ctLpVrEmYTxQCSJEXHGstz75IoBK/kuLzrG51yR14jle+99jJyCpo6DbO79xf1jdZKyIlxOGFA+8
gaNxSSu4Jh33lwpFEzKsBxsz5Z4g8G3n8vy1uTw7ooh2gYwocNG2daxcNf2FE0CSafUAE30lsxZH
PoxiVZ1paf3M+8PZ+CJFGu9t+Mkdtihpx3lGl7Taui2IrsTMUFsCYG9i1bZjtxASWFKTQSjoGoz/
lYJfSqvbT5UGuGPQPqjrKDeXZ3ICt+Uf6RoxK6lRGcOB/ds13XYroahIh4nI+1wMSQukY9zpcvmU
qrlVuQa2m7dASvEf38gTB+apjlmbMNv3ajswy54MW3548qIyRyq6fBRxYyChqldv6GcxNmRp/SgC
Dk3m2+mWyWomvWInGyqFWY28JoU8uFFVM9lZYRXz1ZKf3duCyFTzzhAGwv8ONyTWt1dZZt+QuM+J
WWLaLf4ZHOAPtAcg5F5N9RFgQvRhTk7Z8Ntfb5daglQRZH7T5vPbzzz6AUOXrkLxx8FhTl8kzLbn
8vN8ocpxqjEthzS+YtnRVjZ3xXsMexL4P7PgSQEBIPBj37Dq+4B98yRueIJi9UE3Pi7OST8FaEcw
WS6d4iDpS+GLLn47cSoB7EPxA+enho78R8GFlMmdyD901MMrqkXUdQ132qsF0k7BIZX9HJgPAkLf
K3sFOA2q2cDQ+jpUYOPQXSb8P2D/rLr45k2N35UXBiaJQ2fDarVoyO0p4zS1ByRNI78jO80bxTLZ
Md27wW00fK4JvrIE5Ul/lN+ne7YzS2jwRzpQGAjBzlYnr+lNoOzCLSoNVi58LDW64tClx7kRrQDB
X8HiTSKFCDs+t1Ow/LWAO9ilTK7GDmJbcB2OxAzfvVFj6L0X7FdHINT4K6waEh9PosuYk7l2V7tl
feEMhGW5fp2RAYJxeKQscPils5RhXx7xfjRuPcqoIQRoeIGz5ki4+n3Mj+sFETD6NGQdcB1eadBM
SicMt8FItQ+/MULTOP7BAkBlPVcYdfKf9ozvdGJ2/9Z9y5oMo/6kOb69GG0mY9fkFlvJMflznAVO
/RgcM6lO5N6bJHZLa+abb/hLpmghfOuam+y/YjCAEXpiZGzrCybUr+68lQKUJ4CnaiM1iPR8fNSd
cQB8F79zHvBaMwPnyq9PbYxwYJxUzL+pLBNX095BykrtHDclOc5wu0SIOC6XpBpUSCGcfO3DlWMw
J9RJKwOemcHZfO6j7nJU4OxTdUU4GL9C8WYE8N8L54/sppfLKb/Q+ibJYXpqRegApPVSXB9KDghu
0tMdgzrAds9rOpw2PaWq3nckCyQRNog8dBK1X+Au5zj2c7XgE5nP+qRrRWU1jxdfWrz6GVbaV4Sw
3XcONFNsoS5oFA6vV1u7a8S8OI0yCUX3fGhVOinkEPvhXyMCQzTbNQRj4OFvihPaL/ACOvw5xOTr
OeZMwRoAz7c0iLylhX4al+b8D1m2QXMpqBZkEJHOCeCEeAfRf4eHQVU5sXSJ/aQuhgX5lF7Pob8x
+8B5Iqy0KHpID6ohQuJ2q2RS+Uo5Qhf5Z9sH100hXeWq/nTSH4ENin8K/DF6YRFNAGTJWgU8e9hQ
YzfLYhGX+ohN9sB0YksxK9yOwuBF5UV4pBazmnl7Y+lTK5yKOWnU8AjptH5mCwas5rUTueYVAV01
86u9VBycjasE/bmatZHsFeIGU9htVYrlQuuEhKHba9bo0bpW6kl8Vch4pHD9MtDGAsCU08VuDmRU
T37BBmGlqZFBS9Ma3cW9cVJmzsaNjdvx+VN5rfjUB5cRuz0wE162kxaJCerM2fRNgLvp7CgR+G9Q
TjDO6dr74f+iX5y1M50yJbxbxohL9LlDaMH1I9Xv4ByVB/TUTGNEkNt/JV42sl2U+UqFiADJ4DuN
0liStYPIHro9hKESvRijEVv3qwa/UCquMuEKomzIohZTbJrEn9F00a39igGCjHTUTSukodV5Lxfn
sF4Br/HPRAFOdc3+yN9SrnEC3iPEQdLqDe6+/kht+4Kig8IKTySVW6qOHI7st29Q2YxpkQBSgQRc
ppf51+lg9tkxBmYQ3LTtxck1CQ9G92GKmGmRgwX2G4wwH5uwq6s4ojBoonO4F33VXqs8SrWGA9ZP
xy59X0ggXKGF4qjz0D5b5R/3+OMg3OJmeq9Tnd1CEu1j/Rk/KsSRl0M8XlY097CpQ1rT077/MfjQ
NbCYVsypeYzPeUiavfU6ChJqkqoQIsVXpT1ts5pKaR9/2o33lKq0M6kylFSvtUMeEpnayqegv+QE
+cdi5io31X68UFU9JZ++dq3CxmJdaOUhMdMPtvrsAxE7ppwp9AUibEyXeQJwaqvlabYGn+bx6SNq
m9mQ0OJXz39FrqTxlLuHwF5GYXZcBxpfd5bYXezqKGKicQFihpv9btUA4ZNiUxIGNWPYIlY2wr9E
/j9gSHwK05aDRYCzV0pLIsSatoTgDvmqKwtKMuo6PDBPFNKoN5bM7K2i4JWW2sLdsq/GFHD1JWBC
Y40QsWwtCwOm4TzcD8WkZcbxatwQ7FcSqWsRsdjueJsH5iw6UngAUl8yRsUAs3FzCzM37WaPfOn4
4Gx9LkhgO3u3N1y3O+8/69wUE84HMlq69yMpnjng/68uNyxU7J4GRlk+XOKqBwlRDfHEe6O08iZi
6Pzj2T5b6aNdSWhPjVvZzyS0OTXFtRFHtxPeELPF+zuRVr8kuQCnthL1q73bHUTB81hE+KtyOVK6
31Qsp3BlXgw82suDLZs7agHdInjILszSU7GbwYyteruVb/hhDwcKMlArbY7pTsr5DLJPV+iiONR5
AaSwjModi25k+0gS6YSV+BNe1Q0BaXDMcTc2LAXR+70Wy5s/Sorg2o85fcOyA1TX4zqbkxrqWNxk
G6OAauMJoM3hfCeBAhAgt9HRSlMwyPuuKClhrAZPFYXwicV7KOL3UxqXSQBchacOay2gkn/AcbN2
/IdEchn2ANP2ZJ/G829IuVTfLEn/mzy0yVcQD3SiRU8pSk3Rlhgo4AucBztEC9PtGoJ/5UqI++iM
hLbcP6D61UxWYn8tsNmv9EsTMsM428ifw45iFSSYwmGY6xY/18v3gaalM0mh0CFHFlSDnPqPDc2f
w9EVLVPo6DloDmX3fOTPErLvBn1hU92TL7tBYN9VE1B5XdieYEkyKf2z+xeYtjJwdRuR64KjJZUk
Bwcg2HbX8H6URzjTez2YphZ0KQY1MOrhLmbpXxD+0ssF3x4EO9ReT6h73b+97B93NmdnRB6Bh7cx
ax9TquKUeKnHtKw06/j2YBpIEWijoEYzG47uaD5i+wFX6nJpjbSdtDhIehUzzNa8NRZIXGvnR17F
luyMa6omuo8iRXTb+cDNUIbHkM2KKu4dOWkaeIIRjfIC23NsFWfr2JU4eS6Wyady9g4n8nPYod/g
Ao8nRglShltMNkn2sOu7lMQYqC7h/4J93qt9AKYDtZXEPOmcRA3pu7QT63hJ6I0JZb0BQC8OS/oo
6CdJ2E6/HroF+3YzeJ9y2FIlTddR+/8v29KQppxvlKJ8LHt+1CsMdqvBTAKWwMNuosYr0ADzOTJM
3O3EvSldZrAeSzHFkJh7bxb8kJQp7Rm0sCbe575zqjHfohLs8CmyJpRohPfQvwD7Hr2mPV2kcb4G
h7L4AffwyN2d2Ahs4FrSI4YGF0c354yqLPBtlPMOJg/n/XCt61vpPaV6wXZHNGUnytKprHQyRcPr
1XY3q5ZKXVEI8LDq2qGKN6Nh9lXbOJwUckiBWIVehX510VUlhaBwaheAmZSoE+AO2SoXp2PwUqU1
N+zZaeaFi2CuJnxEmhd29BLw2uMf+VfdAW0vFLbk6+cyqLRpZ4Ox1Z+Wzx+UtA2n5bhipHtkmKhu
Dj4BfamvW1PcDitXnUtxNcnC+aOVS4GRfUH8ixN9tcmJ6dLRkD3a7ezu6wBrBPpkiMzYhRGCAq9q
9eSj7izjB+/3rp3eEFysbt9R8ogQlTjC4Y89wUhB3iQ0/ZiCJYFGphaZumcFkN0Bg6/DiZdYki24
eNkxMQYIphb22yfkqA2qa0NDnyujBIQ4757Lh024v0i37A1lAWQeaA+sFWMTQWEwHh91pE3mTtMb
I8m6U4PeMGiFGcWt5jAanr8Uwo8GYl7Ft+fCswTeTpwDVYje1gJJr4CLFjxmiuXeQ765Nbhr/JZW
DXbAufCADcR1B4z9cu8NQx+zbRROCC7KTuMDnkledgZDP0vgRJdJEd86EZcroVg6fIgP+DOdh2ci
j7pVMB8rRep/Epo1Vlq3UJK0CY+a+VxSaOUGy+A7ZjWMkthMikUum1m9CMnGIFwBVFZZcgr1CDNw
jsWBCgXvLm+Mo+kvhtq1oY+TGuJpDZPGei5OVdbbJkAP14AwjG3vDfRM+3QcpEzNCtDlxqiFSxg7
poCedkbT9KqpONwZSPfnkldcslAI09DZrOC7D+lOhrCeXYjzUw/JsylfFnN/OBjJQW1YuqbPfyp+
ZV8TlrNMDV8+IWBr0sN8K62N0SzmK4x6SZxhiO8NT8m9B2XYRtatf3YJs6xiestWyFZZTNXVKGuo
xiXcHs1YULfEsmawqhu8VNFF0bvxVbRAxR7P+ny/hVGABB+OSnIPTB8mbovSSEDzocLl9WfCdV/r
O31hEMAr2c6BcnlwxuhSIoqkQE92gN7NGL1hDElbtYEq0Oxd7xryCWz6Bhs/rRFVV+ikL2wRx93x
Xz2TU3k5dLtdDYRjvEqCkYxIa+ktqyCXxZ1rAJB9sCRkNyMXWmBnJ8MmbECtQQDNYscb3b4czvNV
X7Iv5NdHTRPm5wv7K6NDAzrH1r1pLZLbD/Wk1ygyku/j12sIkpFe9+c8eC4+vEAoNQMbEZvLA0zV
cOO9jxQWDXjZC5RYqHXGBTajHx4SeU+YbxfBxb+AIfGI7+JMVeDqf3HS2V05dPY46ITO87hOqjOT
NLI04WhuQs3zEICB6QSKz6jIAJUzFcAM197/wwJ5/nbHiKwVbfdQCVYFPNy58KUc+/UoQCra4C55
M8XWr+tKGWhIrTsUsU1L2DOtWVFXJa2bA251GDChs3LcxhTUJwCbfMr5OwXBueVMw+mJeysosnlh
VMEjfb96ifZIy7UEUEIn/KHmfJT9aYPN05/1tYcRPLe3Cl0ZIUPpGbJo3oP+jNJzGvQ6ea+8+3cF
M7otihoOWkxwB4JGxaT/X3D9Kg7DCLgHkWaDUoOmRmKL6FOMkHNyTPa8nhID3XenVgDFpvi2WePo
polHo7DTUzMIhU2cDhRbpCbtXvpIMDefVjdudexWrmmkVSe0wGi5gnDEVC0CBHBfawGK8Z8K/kRc
Fe9w6PMRV9Acg6/6JtdY5dUdjsr+CPnMtY+Yxqv8cDNSZqC2eIbvAwLVIRImrWWlhfxPlV7vRz0n
5JZd4m8s76/gdGLNIjSwGscmK4M5Ev3fGWftz3+Marijrc0FcoZBHXEGSuTi4usiGHRg/DkrkS8y
EZYLtVSqskyqdLhmRKAtN2oQdsIDKlA2Y53ulQKcaTHgaHy1pYlOR+Menepy6lmScGhzXnbp1yWV
uhQW2ELO6fD+aeOdnziOkalGZLV/r0G2zfSisLwJ4ZuAr6nOtC3vb9LtODqGc5OWG80/QtaXuR/f
fV0FNxpPdVGTbiJOV17hqBQZfPA5tHseOmm3rlN6NTTQ2QPpsIcIQroUZznaFO+qV+wTUnHE/+5p
EOUZ2vpqEV7D4NryJEWvu9Xhzl8Ybgqy6Iv5dSbl0W9aDxalDlag6U/+POs3eaoY+0QpFHgx1hWP
kcx3ze9xg/sR1HvuoEkMtkN/0mCgM2YrpTXz+Fc2+Kll5zS4QzEvW0VheTnQJIyzkScEGf1EOAgS
4VTQC/wyIEQoLoLnpZeXyqyQORXPb0dHAITbnwlIsvwp0BcFsBhm16rpsA83JoVhvHz7M/R8h8Vl
brTvRXXm1EI8Mu1Ml231t7C5HSocQGgkgPlPnP1u7rMSHld19YmJ4iAJjPJQCV1Yg1TsVZt4iGk8
D0IDCStWeclc5acfb5MudPp+QvsqBwA7GphjbhN29wx934/Cjop5oiSU+OeOCg8wqA/Un1C+dQ1y
YiSy8hu0VAmdOkSaPiEtfkRHUTKHGj3UJfcfBJ6L8HQOlfdeQywENd9gDt6fk/5jVbmC2/W+d6Pc
B9fhs1CLEXGfnU09GrP3VnOfeZSsMcyELqxmXSrCXRMbrlAmim6R8Tnq7KoMGR6HKWcaNxwX3aSs
h3S+76awLEdE/T59otyQaymsvao0/pn6b7vdOzZ8DZuKU17+wpxumMNTX/qi5Dl+SQPQM+DKKAal
wBu0rRYhX1J7UzrGY+YFH7zyYC61NnWWrOuNx/uh0Lelu1p6KE53zzv4NE07XtuKZ3VCT9Dl1MuZ
EOayzHzi5aRED0aSs6CHWypx7/oQdl2TQa5o0IIjMZGmrUsq2Z8cGD9Q8oWqYQYWOz8XNfy2FK84
aqPPZFFWGXBCo54DQaHzC7+8ECr21UhNLF0dY2mHmBPOymaI3f6mkL0H08MO9T9gwtCwUS26kzcC
Fm5GDnCl3kZg11poBkOO+AbdxJHMXM5akrnZrOU9WHkz/H/zkUsK2pwToGFbw1jfpV5idESHIRfr
7Q71s0U3ErkeobvQafUaFXDaPJZyyP6guMO3m8XJy/yESrHKEFMxpecXF60+JWAvVCiCrSehqGj9
hH3uLHrXRl6IoJsv9H5+tcS4REXE+jARqpPa4+SkKAC9lXKOY1e5TUngvnvXKG4d3V2bD9klkcXX
Uc3z7b2GrmRDrVEzYKvmeiw6BdqL0tro+rHFWqYQv5I4pFstjnucTAxYc9ygexI6ZqilfPsxTpeC
j5m0nyRDA3PntePfuK88s2/dYltmUdJ+yyaSzn+enm7reOMraqbjsat6aFULebdOIpwH5VyDS37t
+nwyW9cVPORaAN2meeeTtq8RqzmyfYv4/KDuB0PD7QyH3TmtbxZd8wecO2LoXSNMDF9aq8ojpgUg
op7BodmJ43lH0jQkMcnLtkmBXKgZKtEjyEvBYRdagYeLyCrTnSOsmP+U1x+gZ1os9VfcjDf59UbB
DxnxOJ6umzQWjIfkQahOxBV3OxXa3Qj1aPh00YvlWhkSse9wIOnRBaV8mr5p18j618gVHvjw7S3u
c5Io0+nB3caMMcHGDcrktQft3NvJryRQHoS8IsUmZHPGn5B/u/Qy96usxTYXqDHCfLYf+foL6S31
M3As9yLXiHjSciLMD8HRBpU5Y0chnI+ZgKRQ8EjrbY9/NLA9jtd5eYIQsoglr/2xljdS8JcfjDqI
D6ETyP2ohAoqRT2xdxrys8eECfaZ/0YqVE2ICjPYkW9Mup1FJ9SLZaUrygCMbuazN/WoWm7I6KFi
gIZMtJNAOtalqu4y8koMiCgX1x6dtjam8LngNfmd/+GVv52tmxkn57yWZ8SYfDVtXmtj5HFREYak
AIyH2/E41w2IIgCzLvQvcYwtK6XIsiXtTUMrdPW5Xldat/JInQUJ3abQFRUqIVWg2iRoOhMkuxmC
6kLEAs82xXqZ7OhxjfhK+cv4JU+MucYVQJe+rOE+v6cNNVHOYZk6EzfE5qECgLkn+Hwd5+kmuVRa
B5Z6pcFOFnWlQ8ezakR4oEX4Bf5/37HpDslZ0GIuXO+CGDq0CCjYebEFkjB8x+KHiNRBLdHHL2Cl
0sEFdB5IDcj84CzRqNUqpjsGbP8jG8qtCJz0nn0Pl1gyumLvxdDKg+Uemq4SS1jzjzuwhVG2l/Ym
Lq0enthDfsD3fj43KecAhaeaP2r9JorNS+iRtmVlHD149IubMjee2KcmA41pZItCvz89o1C5fHah
5qxVXw1WxyBpU2hvkpkbpYnRpfwD/ERYygYQMroTFTy6akr1rzyN7FxEuvRt1XJ90yRar2FiUJe8
LCYs9K3PY1yXTb9jKL3A5t39BXI+Ui/26kYB28c2JptSpqSDoflNqF0TuAgg4ZDFGcV5rtlowcqN
rQb11InrRkxj9BsmQTRk+CyuyInMVH932bFXvH+3nvtkZUSh0azICHCyBIt7sV5dZP6ZlPZQrVIn
AhjK9Tduy+SRp6jkTydaqU/I9cQNdTDUyfa7jZ93aShOSuJ/idXrp8XhZm/HkSZKfyuT/96jp9qP
HYzgheFEitv5G+rDBwCUQ61Qc2fGIRx+PVN+5mktBq8/UceD6Z7NOiesrrmp+anYIyx2PFBzQWrN
NCWBUHIc0EcS05oox0FEM195gUEEQorKMacOAPglNmr1huiXxFDwzegveTuE0agj+CvQL4yDsh5K
D/uupQGljusRbJFhS/oMbwkaaH2b1pZeSqZTayXhudxBOZn/S2oWVbwdf9hbl/l+j9Hzcn7GfxhE
59/hUluX/stVp8ChJhufseauwfqmqPsJ1J4UxHWE1CaakkdDbU5qV828wA7ItQK/0LgjXN2BZgZ7
wlZcfuozDbylY4oCY+phlISH4wbzAaaPPdeSR71nQIFXm4NvAu9Ccj49l5rOkWXwRtiNw1Z8E1kR
vpj5/cAE6q+P6xhQMLmmthO1sT6QBLCiQtZ7ztysVBtzYk5hPjfUTDINwF/h5aESVztrWK/p6nHv
q0SPKXFT3d1lZVDesTklkADfkeezOYVv0MnDPgnm/F4a/ANki6e+9gZMLg5Ge1aa62QYzFLcnSDI
T/VYeIgAb9wp4xIgQ6Elp07L0VbxztfBYj8fq8xtgbiBiwh1RG/ubUBx+FEvj1UnkJJiy3sRrSB7
vFfDaUtrtrm4OKa57o5/UqC+GFFBSLJbgFJr9OK703OszBo5KO+QEuYQqsPDJSwSFis+cA5OGwaQ
oxuzWpFU+ZiB04vBepPwOob5yOz3mEsh82kOrhOmXAH060REfpTE0QmfFw5m7hoqbQlAiiDMUE87
TqMbvU2615WntfEjyxGrwtIcfXBoKc8gvWuMBoMl1EQS5CselB7KscxOqWzpRsMrS2aRuyCotRD0
iIGtOf6vtp7z28suLCXHefiWXd8XTcnHPC1/OSOUmP3AP0mBnnXy0bjycAR4cnofJTTXxbmO4r+u
fbQtAuSvXLtLveZq6GqcFszyWT9ecYK4h+HviN89iq1oNnFZ+5wTo+ky+zIeKQXFIYlTVm/HmKGo
XWHkBF7HUI7haRzOj2LYT+zDCIC+ZVIKfO7DWuGB2Sv3B62ljRz7Io68mHhScEk06rAP2YQBqtOh
BUzhrM7l2adrBAX4UjjD7DPnK4ZCAHtDg/2ma4TxIHtZXW5ZJGsOZd/eOtX/TfsVTBLUiNeRKmzW
e9YWndssI3e22HhdRsyW/pdIrn0KaZhL9WVFSmhDNdmf4NGSgWUZ4Eo+zMe1PI//FpkZN8r8czui
R9hX18rDb7m0QiN5q1ifnJsemNeRUZWoHqYr82BPe7j7hSmQzPQTI1iQ7FqUjruWYG7xTxJCRJAI
BHel/VHHbgVTfvsb3sapGFuXZNE0GjbXgb8YFbRI+1l1dEH1SjRcyoYx0NaOPtcdw1+yTjl7REKv
a96yZ+NPCO98/KxW7NoZllUjIUxqEbMJDUS9Xe4G1+ixartOgqspVfd38n13wAN8DoNxrUC5ZXhk
yqHG+kH/MKZsBEFQWoJ3b/bwmljlgzDbTmLRN7RrQvfXWfk15qhmxXxYVJ5CfkrnkRQ0Rl86xgQA
U3+XD97GZbZ8gnNSY8liYtzaBoXOujytKomZyg2OYm3oTA/Hm3w1PfsUeyoDGIeaXPZKydMx847Q
KbKR3KzR0a6ifWVXukmcPLPQ63eC+VA2Br25t9yOSSJAYmyQ3x9fYvLpPeTGB1b+82VEdceDT7I/
aBuzjPfxGiiyxri7eUJbiTyyuHpYVYJ1iRkpmaJcOi94MKBFrtfGmQaWQaWpVdH75PKPi4LHoUtO
wQbvsoI4eLe0LlyokMk3n4UfVcqKF64C4lpmGwqoX+Ak4GPuQIq5iDBIA/TayvyZMYUHXFNzu2rR
RXbUqyqEr+eULXwoLZLwC+Al5sJ8u2sgp5yaKnAqoDwvXfcGexuS7xOKnW4UGyALOJBKjfCfLpJP
r0Dr16twB5ktR6cvyZjh6CEzsAIsz1lhoruVdciSP6PK1dOKL0XS1A9mQPeJB/S0KQVl0JlVxQB6
gHWBBYPICVnMbfqFxRjGtYa3BwkV+pbqtb9yjgM9TnBTgYqiRn9eQWmbfDsvt+PeWGCq7jufr6tA
r0pAxiZ8/x1EAcopRwrW73T+x9V7SKUmYGCp20oppMZAk6sqYfbk0ECBu+ZY+S/teJKEIjajz/9H
6xh52WgnMOulB8QvtB47e6UoCPSRFK3mCWhl7+agANrlXcP7fqP5r9B+cgf8ryvn+BDTUcVm+Qet
bj9/MG/Z4SDRPQALAfrobGAbUCAgXMI4xbTn8V27jKmGLfYO842KDz6BNHmbPQf8bl/lKayiZ32g
+Ns5ppOfS0cpCzJ7nu/5OsLPk2TVXV7yrAajkax4OGvSp4qUgj2cl3SHlUDjGJi7DNFAExzPL/y7
iyVv3nYBfX6oC1NXPkNfINqCeAjv1Ymg1nUmJVkhHSIWPCtap1ixyCk6+awtpp7zeh5/hLctWOaq
w6AO7iuwXojY4CqdF3Bbnu9K9dWDzm9c8Q/KwgRm45/6GOSqHQqeEqGnGoah3qxmRmfkup+62tGH
nm3kzsruZIPa3Q4PxJ0GSCx3jotqcTjFKiLo4Nufb7QsNdqE80TKaGRH4xX2D4Kjv2sHrHclR+Et
WgxFlh6F65QQFcyTZZiqFOHklmu+ihgNDZRVkIkA8/GIO+Flf4ZY/eOGty74sfFVnt+idGPXdrX4
k9nbolbvVrKNn1LOfanU1smw8uV5i138ktYLXmdsUs4Ih7EaskZtr4Yn54QTVTtON4FIF5TJuBMh
Z8xEP75wOJQIbRAd8aCeLu36N9Wxn7UjeARSLD9CDi0slicbAaAkEXegkeK2Xz+YLgjCz7WV9GCn
cRlys+1F3OP9KNWNSrdaMYn5mg7l7/PgPoQZHDr4drqZIvIOe0SFBxmXUTvbWTxSQaeSQACS/abA
qxNzhmM101Dg5LLPvm33TYKBCYqzNMrICTzAHj/BxtpbWNn9HwKgw9tADU24bp4m9KO+4TJv5Xne
SzSvH4pqmHOJfnt/w/jYL1NRuKs9aXj6fVUvDmQKp+tllFwZCtIjVgNQNCe3CPDux5I8kduAi1ID
VvajFD2WLzhHglf/7UcddEOyb6bD/HMFQNxl/U0q/47u1nhuVtMjB6SgfWot0IYoTyFOCLmgoei+
Bm7hjBGSkRJqH/W51msL5M2tmEVnatygghzENxUnDSFD+m0mWZs9sXWTZ+B01eeiiTfzOjYasFru
45xuTnSMquIaEaPSqgx9D/bADPRFVTfWOu7X051yc9rr7cyNO8Nqq1/1CoSQGqOFfBarPFbr4a73
ewZ47IbgkCJ1Asvvi+62z1j2lgW9pCyMTUjH/1Wqt8CKwcVLZkbfWXhb+TfFavt+EsbgZSUDfbFl
7E1oPMqDcz2SWHRZeuXhR1ieZkJ8Mex8povdkwbGAqtmnZuvk6ugk4xDMrkmKbOsmB8v489H2gyg
xKtGkSSbX0XQ1QSmV/feg1WEq+pdwytfPSRgvHBiXQfKQsXDxECw1Hztzrkwm4cIU6T5Ndk3G7kO
xrdYheE8MBtsyaZL77kDpNp+t1O35NL4hmCOVNT40GOmxvMd+Ajg3c7dBW/y8zx64Gkys/aOm+Wb
aPOhhMFE2rhd90eLpLSnwFzuxCAjuFl3Iu0Rwr2CIs/EruIyXbHf7ZSj3wC9x6GwulGra6MK+WDy
2vubdjWefJR69K0a3xDYCun5kMlGGUCKPu4/xISOYQSnotFqKWoCI6U4R/tfQnna4qWYPOyp6nWn
ADqFNV9OwduzHOxg3li+SJMkepHXPbQ+vXa/a8Sa7chITo18cCq5A4Tgm6JayARw4I4Zyx1/d1MC
sJKABxJNJui+74QTGB/Ut905XQlvIDevs5SvXr1ZW0TiM5AbItLlpQvS5f9kqTBtghu/+L9lUvCT
hSyAk0SqkeniEvxgT06BYF81Kgt/uBwCDmVs13Pg73Zm8QcSUyHlyUKOP+eHaQKm1PP8xHe+gymr
8KMp8YQ5E8+G8Kri4oUnctuUaMGpZpcP4b9bOMg3Euab26/S+wulq/wpBYsxEbjv+mMh738zu0qm
lbyZfPsnaabldZ2lDXbc32pErjKRS1KUROyOgIqp2aB8qUzBbRxsiG2TajpAjWnFeytjFDH6Tcmf
L+LN+S7EylGcGdXut5CdvnRmk+2B2w/734WMF6JigGQSEXUelNc6w9Pm30d24aWIdiCF7YZrmcFG
JtReT5w/8TNF5BEAOlYJDmn7pUJjQvqeDrE7Zm71ZHCf3p9IFYQfNPRslByDiRyicI3sCIA9GWwr
YWP4Dy8s/W5P0t5hTfwCwGH5bfpUhmBR3WHgsTbcPv49Yr+a9iDFOzJDfc+E3klWESIDGdPDtx+Y
m4BuzWIeMXSdMb8dAnZwaoxLM/W5o+oTa07PO3EU5e02Ucjxvshp97mqXRoSmzHBYhbZtB4em4pt
WrY1XbroRJt/JsVZE0lXYIC+JC/NKuJtJPkcKkp1KZzN6jBB2yWPOhOXbiWLmWraaDBU5IoDg+jC
CMYhAhYkXGM3kvBQ+NgBPFB+krJPjUwH8fanTgHnYeDDmqUqjnEXu4cjdUQ3wxOPKqpANhTa+8gI
s9cShS4nrzbhO61DPBI07I5EtzcLrkDUJouhxsZl6UaJ1gx+rs9+AlTGpjZVZRw+KJja0zsJRwlA
KOc67s7/crqGPUz87K68zebTJ/DTyEqqGINSQEX7RxDVaMYgtvIGFzf5Vbx+qT4tbxT0ojT4FhNd
98SPcfArL7rJ8go43oWhrWAGuGvB1sl5XfbdQ7YPgr+Ki0PFTg5s1+zwZypzh4U2NdXVV4nf2woN
jPKRinX1PdL96DvZnSl+2SINqvUILMwaZ7hH11JelAF3HfnK/v2umEXc+tktukHHqqHKNxiiHUw8
tQTd7qeAJYOvcFwnEf1bLjQIUTr2fuQFezMS2WIaiJDTQdQII3Kih22Tu3MC2HkK3eIYHXkj9mJt
rx6PdnAC0unrHXYTWF+5NtD08GdWHumDREdsrWPGtFgI9e8pbY7j164USpHOItorwhNCO+DOHfKn
NzEdVqy07IVwIu++s9L8AA2nxPgA0orpLK7PifzfI8WqqgIu8jyrklernV+EDG7ixwddxTwd2WYz
yoiqSgPmNbu3tnik2rQAqTWVfQ5uPTCLJql1LQpUzT0tUqt9RPrJdU8h+2H2MDDl/0i23eRZseZC
Bx7Md+8Zzs2fMWiTIFYKtY2AmFxtruQOqoonD8gjVY02n+BZPV8yTwO2dS9ToOr1azivnKi1U3kE
T0MPD5Vywr53qp/eSHFVqAf6qboHzCQJVHZ5qUpltY0n7KSi1dOidmtJ2skb0D07Xx1/fVRgdYf6
W/lKMb7SEBYD+AMrQl+z0CUd0RZg+yTgaDtRKpZf6EyFcMRgG56NKWXQxEEiMCOkWINdBgJOy6I7
o2+Xd4369QscUUvm9ssdglBVP3jCRh5K+hXwNhNnf1/8iu/E1LUVu7rwTpclG7aK8wZ9ik8Gjcde
c5D0o08zOc0m0MOOfumC1f7XZPqTVbL1zN00iT4K+eBDZkGhb0vZQEFzCK94zQjr93uzIdRBqgY9
GJLhqjgbubQOiLlIBjYyN8HPFXop/8N8W5WmuXmLIdnW2bjoP8z29NOxZoaX3dOjpIG5prKNQpsH
/qnhLuS1daCncnGtGQciN6A9f9qZ344NLWUXfvIWG1snIk0w3cwRoH8zbNuxfk0CKnV7R/TKOGCB
oshEA65nPXghyM719ucpLmgblVKNnsNBgJCALRaBca4EClpj0dPUZMqyFRG6cU8Qw0PoYqRyIL/E
FpyW+tOirkqspjazdDB/Pu0FWF2Ofmkbc7yP20opBjqLaOry158G4M3Bkp58yfLQ0cjU90Kox7Hj
pd+/bpvWXZVhNte4NW91GR1hY8yZba2QAkffVcLC7PJgvi27xFkC8870uHsNc25baDXaoghPmMtT
dyNxTl0nkjJxdt2CC+PxwIgJsvPtSW1CnFVaFGDI2YKsmEwVSLWdM2bhOejDZF35FMhkwKcH8rVc
4bq3r812JpJqglG4QI5IXehalRIhqcmd9wybr8T6AOFriIcjPD74kctmCUnfLDVjFNHPQTlx4RuE
HIW+k0o6DPzJYlxnoA/dtIMrja9mHoBbjdstAWzER7mwioUTRcnCsZ+4DAN/aDksDnHxKIZebSKy
Y9QRqPw9oCM3+3OIq/iVQgO4uUCXLQeRSIrAM47HoHHkJqN5/4FnPCAkKrDMeXlxp682iH38Lx22
OZ2ekqOyJ4ns5ydpQG/2lIKDauhENaYbUEquG6/aGG6zgyUbPy8JxYRJRQhyg3IK2ziEfI+NzAFn
UDmJiCNK3vTiKykpbjifQPerLzrsqSCI3OxETtzIGw7ofwNNKA1PX3h95hZejvHzbFc/vVNE1Roj
fRGTVKzbzCyuC77BuNrMYVo7MPk73kkYILcicQ3XcvJ/iZVOJ5UHCILEVD68vUyZfh/1N6UQ9JMC
P0xFqKRDsp1gpFG5Q5wuIXOigmguR3JqmfogmZ2jj6bmi4TTLa37n+HZTmFo7JJrubKr68cnoNQF
4hfuiwbcVNmcqPlANJ5UgMBrSfD01piR7wknfZsPPcbyugPot4JxNrHM9COoEXj68ZBsExrV4n9s
Z+N+7wNKDKRd7THq+gEQhjNibRNz8/ir/JgKHXtzGg/92xHQixsVB/Mhj/TJXePIPOCuSxacHSMR
oaEc26eEHqsILScmC+/tfww4qF1j+zNBCvI3DQcCIAya6oTa3D3F8TNpHJNqP+W3fkAmDg/9oWQQ
NjUDvrgbnMsimiDW/Tu+k0+IdKawRBqgrCz0cZVq9TuTR2SfvZXChT2awKNHYF3aJ2Km0gqklzgG
r9W+MNRT19TqiRHQlNAn/7vQfH7G9GBEXrMsRjAvsQ9U6+8gV75MhQVHMp9rOlOD668L8q/fx0Ha
bWl/JpfpXEXlW0wEtFGlGTGeZWBuehCRtj6V+J8AsCz2H6lbj3yAWr4yl0UmNcULvkTJtD7Ky0XY
hFygvt+/v34LLL8UtslD06cQxmWhqoQpDh0Kf0KvUiNhvuNs6kTd+H6Qx1pK7g+Q6v0a+SyT3SiF
Pl7jr1gw42emmGQSITEPykSE/CarGlkuOdRAoGSQeEgz0UjBQvBd7pyXJD+SHHzcn5KrsQcMZijK
vpVcqIRJ6FNtI1a291S2Sv+boeLE7SSzAGAdAH7WrZ6zzzhk18eBN++KZH14ynwnCJGIuL0QKRKz
FKb/hnpvqblNhvatRAtEWtFWi/Xtb2fp/CDoAdUz0vux5gBVoHPA0jvlwWxeYgH8PUmh23pnNVsH
4SeFZ0ePEcHAX9rAm8Zh5LJSdhXU+TCJD/MdeLd/25f/x7YFRB9NRBagychnaGKLHxU3lNV+gtVZ
+XAV+EzrqP6wU4sEs4wt0uvQkTfjT7SMwlmMYNbHDYIa5ZfTOV1BU/SDVbZwN+i8UU1J/+meapBy
DU2TssNegpK4yO4WPLIUsrAtbqQa+2e1k+3ddNoY4UnHHbeW8mti00M29wiOxdqwWwR4lUbr4VUZ
i841Rspf7uUpW/ZThbxHhK0M4a4QU+OXZr1+AECH5NL6rEWF34gllShObUf6YwUWzpOZQYpjrRNE
UmkqEC9enX7eGonqM/Vr3ZiCPMclPwSSzjbh+MhSdD8w7vSdbDVBo8ROpRhbfhXi8QOLbFLtN5d2
5zACiVpQ1TUWaXjZGYv0ttPQL/SZYU8q6xdpKTCEJwm7ZYtQG497gTOaECPx0dD9R+6BuSnkxx75
UvjgAGCbSrattmNeAiLAYSKyekVolKGPtBy1udeSUbwRnJDgjwUXWj6e/p15xj4hJCLh41NQjpdZ
GzzEYp2KRYmPX9H3J3XQIwisOew/k63hiqSzxPVsyD5wf0H/urz9OBa61qCjw1JFjqX1Rw7kzCQS
Ax9qfmOGGvaUJJ0ewAvP05doqH85L/e0gimRuMPfEmi2gDSP7D4bOLJr6JGHQKluQtTOxfNjw56t
euTzpa35MDI5lrTglR3SE5Y+TAUElYae/LxcNflacw0jLbV8D5IdNXgJj32dAq6KSlnjde90bQGy
ULUX+KLA+eoYOYUCTpb9Mz1Sj4mrQrlPw9oy0lJ9VTkzZyLEpiIXMqZyIgiejbghj6WY0f3ig9lq
Hs0QyDpGCzXxe55oi4a/3BJIqb1AB3iE3kT4vpi16UwTWdVSe1+lg8fQJpZsps4sox2lQlqAyN4e
Cx2yCG3DSxoF451ehRySwnG0dfdHjAwvW9hHjaE/05+uRORUkCMKSc80dFni4GhdXdBk10szKnVB
Zz+o5hViPNPq+4WEqaApduxTcWfDypkZUIPpjysdAugMMiO57ySe/qZHTfWhUr4Jc8kpH7sbmT8H
p0ieTZg5/CdzZOFZDnnAUh0B82Mk6+DF5YpRD8ZFuSS9fyaXorATcwRjwhjCXU+4iAcQrg81Kirl
nyv10UKdkll9RZJlZqZKAlVK15LMpErz4TGW4lrc/+h4KF+it/c9JPaOSK2Vz7fyuqhdaKWyR89B
k7o3gY09tTpc3uBIRDlRlErRpWsj41VWMpCURb907SDXccCeL+NiUq6ivjSygXMlQqSz4OcdbKYj
pXnhqxEi+7gpK9EAtyKY8kiRco3jNysRQiZKXeVl1E9wBBpdKQcDsNbMMXfJ8T3zP9YnwilkUALo
ryVKkZW2kXhD3wDT07n5nCcECOMmqNOTPtTf353UC6fMLTaHz3bDIx+yEyZIXOE9c+vWWiNWDt/T
UlV3XqorVYPPgN3FZ20qUeRbwtKO2yTThOe44w4rKVA9okun1xr0PtRkKpGbiedAq3jQlRH5A2ek
c72/ADHYkrdCKy+plnUAMZmCTXTp6owKsK4UKosdPTIVnEgvcGflgCFfEhMt3tGP5Rquhn1feu09
GqB+UwyJu5fqD3zSP+hVzOkDYk+Uu0cD15fylQ+6Tcf/qOFMjVEn9jdGzF6xcRQ1UkaLQcn1cOIs
XbQj1jefxm/OTQRkBLn8OksfBotbd5RA9Fh6Jv2AuvNMhsDugkvzV24uQ6E1L65v40lVWNuhACo0
w6aIwWAX+wGD4b4JQhvDpQsFwH7NudFyqaoQmacvb55njt6fhGUUGhFQWCZmJOYW3hBGoHC+7nFe
3LdXgIu0kVRCKI3RFGOJ80OnAUlbuLkaB5XqI2xskGaGF4D+LNteXWsRDWWIAk9hvWOUSP9soPQD
R00F4Zl9JyKhis0eAwl3KghZfbZPPyk23gHyQCDVYljs72gIgnQSChprMsW63fRvCMaqU7/cApt1
YVv1vGrU+IdyyUcdhrhM+YPG5UtosMk9zk8aICapdAJuwtjM07JLCLa4QYd1omdao9umvwWALUv1
kFkYgt9nPFg7umBz5PbdLBSwWq5qusTeqrT36BJCk5TlCJ2ENUsU4BB5uUcYOifGtjRhQBqsPxqk
x4zD3vWWaXTMqPIY42WEdpiRe70GEZ5VoijLR+B0JpYIPBeYftphzbL10FYR/yGkf62DmuRjwDSv
FKy8h0h1IiUmT3bWOqrAb+OIlsEIkAytmESEFJNzrfD2GIucKoCK/Btr+DpTu87Ou/56EKBle+tR
p3BbZRhyvJOIeOgO+1jUtUHqkwab5IKXS1yGvj2eJM1NvhxhJcIx5zJRIHjOJbMOZBjXeQzfiU8s
08aipgBkZUUj6HHO4+KvM6ApKIfataoMKxHNiNFfVGhk2EBJvggrvo38X7vtYewf8plmc588+Qjt
odqTWybjqePaX1y70LEvoya/D+vJTN3Jd+tXQi8TNFwOW5heistDSH+xOigIxirtlHT5I5jC1nmZ
GvXLNZEuaHJ1rItcP2J5anuW7/tmaqJUHukhpZhCu551yqKLgQeyKW/caZGVkGRXsgT3/ZFIIloV
Z9hu2oFwgny/aY/cAt8K5kgNlKesyzkTSGBRAltFv1zoyqXtpb3vU+dgmKFyNfGFUwqPyB3QtKB2
qnQ35T008U71TJEEYBSvGK9/ENucK7S9yNf7r9TDKGfVJTu/h4sOomBk8J5pBjpAGdltKMI9iHZD
uBq5r5zTLpCO4WVjFmtD2ApYjO5v87xI49KS2VqxO9C4btTdJ9L1hV1IYW1o/OsZmA7kD+ygHt7g
lOvWIPNnPB6QLSi5XLCtNNHPUZGEQ47i2DYa9EovchoTecxOURkRuVowvAFF0Mjgg3Y7baERsk7/
A45yf+0oE5PeEHbMsyMNzCV8VkdvL9X5rCMR7eeerNlvmen/TWDb1TzYETsuRGKBGyanoX0eYTBN
K+DmlLMcRuDo1FTstVmRcCEYdBUx6V/ZU42jahXTiO2kTMXyZ7z5MXnkhxIPb8BBb5BJ99C1Hrdn
pCaQzYVCqDzuoO05XRrYTtz8hWdaMzPIyokgjDamozwbGrUVxv8mBnpZKbDb8zNmXsWBTvAA0++U
bGv4s0TOTYoX/MqJwI5Cow8M1KZ2o9gAgOeDQsrMFpK5xxSv+kUMm5Ax2jFtcDQqz/qnzQCE4UlP
rEBJivBd5K9ZvczJGUJwrbk4z/1+Np1nGVR+BxUu0j1yPJQXZJPw+IZTFcdoe231rLq6ns0PvPF/
KVv2IPNVx/VYN8mlvoIYKvxmSQUS+3ceLR7NDe6Mkui3EhDpLtMYB83bMBjxj7719ODA7Xlct/S6
XOaxjK/a2ZKAufFKUju+yu5JXjjJowqVkCCxxz8hKBNFfmEH16DzIy+d631lsrnJCq2h5b9dl58S
TWBR9dyjHuPh7zg2yxX1cmau7A2WdG5GW+apAFZK7nMo8WLiTGK8vlC1DYjXKzwzhA42n8jnVPWk
PHXmQ7wvQmW+mkt5OSTC94ZLmoXeJqKPlhkpO7iC7BuEABMiArXB43CIctlVJmzawfDJ4MAi+BoI
SyBHU2xpLBzP86TZQCucfNOi+0DdIJaPsMLimr40vZ9DHEUV/+7WPj3U4oN4vx+VHTj2xE4Wozjg
08kW70Lq6YFzKs/tKOyCNxQty9pjjaVGeOT1qItzeIQ9v/Ymmd4sWs0q0bLNGPrzcnkQeiHel20t
6KzcEji+23C/7BuJm0W/HYs8ZwkkEny69pZsdhOZtdxRp2ci4USadF295+5FK2pVQG4nfxcVoyo2
K+jP1FoQbWXXlL7Yhp+gsHceliWT2JYNSCfuiOy0R4wVm8MXoE1oRaHM8FGgeCskI2yYDf6SBmor
ovRyqoLFY4mQdrzp0GgPhVbdonGS9kBkVR748ZwrZhMFK0jqNraQYRShch0U4cy/Nap8qY3xJCBn
zfRHfjT6mqlIDS/Fn0vJhIfZ2Rc+cwN3wtgDPir905oPP/zoSBgZImvnSgVm8oiYH4wwhwWt6m+Y
DUq2LtGOK65mdVJBdS4npU35ex2EsDROVi+v4diDws5lIrvWvVNqDXmA95p47T1Vaug4uxdaLUos
EC0E9embbexSOGzEN/KASdACm4EbLFKU+8brRjzl0vsP0rxagySup2VLfceSIr18eilU31zBkBZZ
SGC5w943T1zPQXr/5w0ggBdKbCb/tqCOZxTq2Ot1HYsrFmJhgS3hTC5TeWVeSyovFQxTgKnP19eu
MtW2F2OUgS6Jze2KNMDp26n9UMkKv5sVq2cuPB2tSFo+YtzwwIhAsiULGZ9GDhXnLAO4FKmVwKtF
MFawcVMD94qRS450lMbnqwjsOjSGtMhQgQ/qLt5499ksSQli3ozSUpvFPFzTfgomkmuJ8d0PFK4Q
n7yXTyrPxswxgvEflcc8QpEQsRi9ToiTs4w/QaPb9eXE0N7+kL48yF3qTHCT7a5oCWY1RtjImyeP
YaRmDduS+YxlE85GaOVwMsbW5UffF9ULe9PKELGTc47+pwfV6Rq7xRasM0+6BfrSu+MPdZO/0KJu
VLJ66D/wltobn7bLIBxUsyJ2LMcKgU3Icnvuza3CGsG2ezvy1jo8SQK/efa0V+eIvJvsw0VN8Gor
Ho26Gf7yJZ0l3rA2HOQdxqk5Oe08m2jmT1odd/Cdu/y7h2o9dHPuBXE4FSPANn3HkFCQK8dbyIm8
7C41wXCRYCcaYGWfKwc9T5hiKG/zgAcrTu2TzxnxluvRYSR+wiuvTQXv85wsPx8iLGCo+2XBSIEG
fA2k06QR+UBmugafTLxuz4l/u1p0Dq9nerQmE40Q5lf1V7XaivmatA58gaoNE/IJDJpbyPtPqhTd
AEHoOXF8oF+m6hYZDO1RhHXVFybViCk+x5d+hf2b7XNxcEVEzCkZfvZX9rcrisoJrAi4vzLY55qG
EszA/Vn/nfSmRRlClsVeHh2RcS/C5YIALzUB4GXuYX1aqvFamo8Ut6jDbAXgmU3+6nr+l/ZYj3HV
YDRSnFdsIo66HDQ3zqCLAajxkZZ8/k7mr3YGk04Ccz0DP9mzb/r5jPhyDe24e90E+ZMfW8xy/Akl
12iW+eViSk1VmfyTmJIr/l0XCqPVYguF6kyVcagdbo5j0fjd/TkkSqnjLScZcIQc3I7l325ZpQ5Z
U/z+aOFpNtdOSRRVBKRTLrIn7f7sr7TkCOKuS9YDVOCzq2alDhn9Z7KpwblKFMT5zClM4/tqTx4a
tTdKBp6Z0Wf1gTagfwb5W0YA96xpzCjdC8yu7Ra0pFlBxTVnY3Rq6ZT3klrBHLNpATjFjUnsYdXo
pTxTXflmIA2SWmhFuZ1vVBxAXkDlCJD9AHA25RCIi6nT0SAIANSwf6x1FfXDu+sKGzIOfIsodAY3
6yufEiHaT6/o5WvPEeofz0aOl3gDRY7h7XfnWz9VfnW2m2lXCcm0txy7UlrNBmDYK9P2qkxf/BTw
FkZ+8cjY39+ZihIixe15vN74wT1UjauuqdUjHG9Yw17Xe6Fg6SOFi6j0hPzgM+tKXucZa2NQN8qJ
vwyd/RuVNCDb0EkFvW4zBAafkezU54Bs65IhSLAPZELa/Cuy5z1QZhaIhyR2ok5zKp9AHvX60GMh
FCu+lEHxmehxA0U8ylkIyx+T08u8ueGGdcwFWfuqcy3HgrsStiM8rgftsCRW7Nckm8rq6ckuDA45
UYjmv1AigYKURPmbtPwcFNqsMNWoTi1wToPADqqc/IYCDrwbhySJU+NiX9vs7LhSLMEpccbL9ZvN
eWto48wleyYqnUqkuf6ZLCDy07qHuA3rhMCH8zf3FppiENnrshp+oaOd6WDByllqMWaJ2ULmy89P
CpVmSSUL4cWeayNMzmUWPbbr3wHdTASmBeE3gCtIdea3/1IWjvW1VdYWUFMRIAb7rgEBDf41Ninp
C+GeVjDGFUmfyx8QZUADyz4NI6JBZA3pLFsDBZtjFDGUuWZq94Wki0Df8qtNS9UFO8+Zb0+z6g32
JofgmDBXrOQKyYHYODW5wsg2wWoNDr8uzTdbflICGBnn+bTDjMKBuCBUEvgMOjXsp2cdcqKgZc54
2LbtSAnUePJZimJxmRh25+Ryvj3KNdW0JnfVBDB9p0pbVZXnyWhQQVobd0Y0nJRhcQh/rW4bHyqv
fS4RY4A5wW1h02jXy49fhJB2JtXhwY/8vATHDRqmOL5PJVcpeEiNW67X1oE7FOwx3De5vkMltzfv
s3LjgXJyOe0GSzxh3qk9HPLs90qbeDX1d8zb5EKG677/dcoa+vzd1xDte3/JvnVve8Wns8aKbMDn
vP20FsPA/wJuXJv46b+X9eGvExMdBu9z30jxalY7w1CMYXjqFJcZ+x0+PXG2LPId/Qykg8rdhjys
pD56YHpakUfCL+Fy+nEgvzyvxIQhgG9CTx9FQppmZZqtXKxJbeIiOfG/Xq6pqJRWmaVmezEwKkB3
MzasvzHI9NrmGEE/gT8MTwe20f7VuGPSuj5Wr9ylRAxy6qxqsk3husj7kFanvVTavXGV6btmZHow
327Ok9ptxHQJ0sYKKdpWR97TIMr2RDvP7aO/Cz2xvujitZmLTYfB4pF4EXbJbL1ZueodawB0Utev
p85c5HozndrCMMpujWm3tynSpi+lqaEqHySeAirBHl5vh7vaVH5mFe7hVNW+cZbxSx8KKK/S5dDr
VyXXsv8+Rx4xvUINFhBEdLxo7NB16rABrdzZ5tiC9813esoScuRvUNVhdheqChbwF+K+08FQ/2dk
sCu4dLDdQIOXg09qJ50GtSNRashS4VthY1kKiQTDLFgdvUWH0o5b0t4foRPZWiVRb3xy0nPFA/dd
W2tddZGADf8/1Xp2SpGXeTSzCfX2uBb8uq4sQWvVJ5AIvTIdWvmtVwpVZm9pvqUatn3y72g5Zm22
jtRia23l9h8HqCpCAamHm0puP+qybPnpcRMB4nbD/L04wk6fZyuJ9+E4UOYSNkzn2W+6/6ce9M1v
15FE9+6WdbDdU8PdvW1qn1yUweZyQg8UOyXV0cChGi/mfDtFB4q7+saGahg6F1GBnnO7x+Y+6J2V
b2so2ospkcwOwBhCX27fjRFD+cTZnNsBqd/vJpIJb0NpnUgDMT6VSJot1C6LLZ0+TQZ/WoXeZ4WD
FDfWznuWflCWpDZpSuzV1jzyiKpGJDB0HcCC5vBQIfMRLRuM92LEMnbi8U5CbMhLsQ6ykjxTdyxt
1rHJ9y17Tc5aDAu89zoVNmiDZoveqSvKENL29tkfSc11f9WyeVsAJa3suCkvP1qX8wGO2zU8vkLc
FglWX0uvh8avKDNfIbGdhskJXHkbVHOY9S4C9/+0lYeFk5MYixL1bjKu74phD/j8z0Y1q25iYXkY
Zt/vB9lWiWny5LYwiMve/UXG7WuNemUvVySBcHQTuWpZl4XEXuL3QtsupVXSXpTIK/dYPBC3gtcL
mPY7CW279yQDW0mEjffF/ekE1qEBXij/MYV67StpgvP0HqtfowG2wUzSQQx1qRU+d3l66K1HmcM2
JzfT8rs8mbXrBz4feq/MjbjYJsiGB3IVuD3QYgCGKx+stMcnpAgdBP0MpzVfBrCzW9hw3Ku6IIh1
bXCBevs/y44ZI+Tb/tTMcL7LjV6Y8oFA4DOBJCv2/+mwGH8tlxA7MWIg1PyvrTWuQN3Cxvwv7Yx9
vPu2V+qPFB6kvd4n/mStwYTxGzVs2FEhpVzWdge2RhjxKjj45b0LCIvAc2cf5Or1TKstv59SqoCi
onrS0pZfbJ+7A/JESA1wrL+vuFVulXF2IDtdiKo/VwlIgTaNtw1jqeTxrP0H8muxfjrTYHEpruRo
zzO2n6YqyZxkS0jHoWVPq6JFkuwYIGOZvbQ0J9aXEGKaDSTM0NY99tPKNUynnY1vEkGH+DtPecaU
VY3rk+3bvns6sVjHmzSxzQwU8i1Wi0dfdhainphrsuchjp8vJhCahuAR9KzQjrVFGmfZ0+RvrsZT
c1X8QmEV8QcUCc39IKPX5VxnR0U1OHA5dUE4rotw05fQcTiATCvdRP4F31NAD9NV4vaWtHCpqZQJ
FJX52wz+ZZ6+DqdC7sUKN4rErvKN3I5NB3sIdJdQfnwx2Pt3F0Dilj8sem9JLtBHePCVkrlb8NpC
862p1Z1KPNy2EzWs7lWEMOOo2HaUhxYPUYhCqV04cZgFfP/QWqSqE56Mjr9u/RbnmGCR3SDa56nR
PsF6Zmf0qXtLUUzNWnJFScQVzhmm28Ab+xuv/UGEfgj3JhyXNe501VRuOsgzuCY0QkHp1ceo3ifw
4R5umPunX15JEuILVFakZP4z24mvaPHF3oQ5m+3Fu/HPXcTOrznhm7xMKnQkFTCADP3kg8sYqPcq
gDDtBfasLO7ZU1NoU/AG4yx7wW816Gj5bEZvUR+S8b2KR8tUtd6AyBIkmSmR9ojuoaLExr5Ng9BU
O2ruEVdDxoe1X3IzAU7hDLqZbMdY2fTzgOz5NcgQDioCVFl/H+sh5i0Q0RZMgxulW5WBxyemHrcc
c7FVO4frogRhDrB5KPznqNo7Ug+APTqH+EzKCJr3M10PDt8qTdQDrg8MdLuwIglu2jphE60oEbYQ
qjwklOKlLBfkCVLVLjBHnNJyYFO21P9SPdNe/UkMDmaRslG/rjWKnn3uM2AyiCwMd7oOH0kZqLk5
yCQtY33+gFKUTXVEHjgIiLFiCtFLVsjz5DZq2I2v/RafKTnVF6mZUdKipv1GzSgPtYmkIfcyHh/v
RWaMhGx8d2uZYmNARkjSm/6teRZZUb11eq2Dni2mbeuV45xpA212NfZgSX81RTf7EfViI2hmi3Up
ARbW4mLxIK6TYtd6Gs04Pxinf7dLMobZ7H1nGMpMsSOElpmIR3V56GJyej8fQ58slp433xuDZQnp
DPN57brp+QIQcoGBqVWkX2i6TlRq/IkFhm7rRShz+Ea0ZVYLY0pbuJKSxH1XJ/X9qj3qbItddfiA
bDq0vgP0ERLKnT7NrMEfyi70VPTs2KBcMWKdJGC5vE54YDB6QXdMgHeksW63WUW0MAZJjVcRXW9v
Ec+ZcXrjNoWbNJRAKz53qB82cGFelPO6roqJjD7l2+lF/iF2iyqzJlzw4V4ca27vGV9wVa0tnrqB
aTXpXfEe/HlDqtrX+f0+7Ax+ODp2hUSDonmxo0iSnIQA/+l0R22AeFq+4ijPNN2mvq7bOLSOsn1a
zepnOZ1hy/boLL1GYYqBM9mT9UE8BWI3je7jCtxslWvEs6MzghZ5VR1C+sJcGZqVOm7pQazi7Zf5
6b7Pbf5MdvnfsAjWitM/zSErby7yAzZlmT9sK5zT0y9HG8UujCOfvBcWnjkdmN6ijcyDV7ccWZpI
EiN0Gw8QFpjlIkMBqfinZ0zu32FHXWmzJlGTunjOkpSDl3iQj8p/I2JvF1I2DqFvRB+M9/VzfbIk
AWRKKdpDkdHpU4FtDzRn/YHwCbru4mfzwQABUbGmkghr7WroI8c2eEYvA4hWbicJdXjPemmZHGBz
AOmbbjaPykVxdeHYRcnhB98gnD7cxYAleq69Ox/uHETI7BYguE6G83T0aBrOzs8Hdu3DVe8ryQjr
Fsotdu/Go6YjGN2V5gpRtYN+fJnzyg1Q6fDBp+HtgdOip1xEPVLcQG9OQ8yV/5bvJO/d5IGCevdP
In1PqDSERgZP0Rd8eWn/D3kAwDkO6VY6rdZGfuWLg4vyO6fO7VJ2a0Rt56AAMjGG/a9/gsg3x6lO
gc+t2/Q6GdUt37HCA1Fr3o0XUPt6CLwo+9wFDw7NmJO3b5bxDu+vFnJsHaJ+mHw579icg1jciHdp
HFSeCWxZOEmDylhCxXNvuVl2cSUqMcdYcpJ0jcSRmfJF3MeOlbk2W9gED54E/w0UU3ZDY0MzjyON
PCsN64pIfEtkIdMxyGrff2rPuSIARq5rKBX5tCN9M4t3BsczBSUjs3uHrJaiXftaM6IqUyAPK8nh
+/1BXind7AmWeapMGSaJBmMdGEz7aomY3Usk6fL55zu6v2ZBgDdISDJtOOaaYdm7bi+lTlS0OW2u
OVmqhTg6sk44yFLuRrwrGh/RzeCzDcmRKhRKOVaCCtPwFtPcZurK1/Y+lZW3922pkfCbmgZXAVtP
52qL6MRPccMoE3QvndAorBmiliGKPDS5za2GAgLlqK8meaRtiGFYFibgIxhkNh0k64WmKIsoYlsw
5mwx22UXuRkltapyi+ef986Kb2ckvzT/pLRkJjNr5lXLsrzl92omBjUbFyImgCdhaKTuI+XaZK+/
FWHMb5gyGe0j8tdIlePHGcjQ0uStCGaOEAPn1p2eY1Q+lslFpgSVZl8EhGI3klmNdDr503OBJkRE
CgwVr+c+dph6PZcu/0KDWR2xtr4rjHJWSkt+EDqEt500mfx1L2J/1RQMaoYRXVzp6MxsZ3pkvzZE
ZTTrm1LxK6BoknZ9Kt09sb1zmYrVtGiE+XvgeljTFEiHQESRR3JguLVynRIPqUu8JaIXq7PMBA8m
VJhr3PsfJVTgTVWFkps5/q0Fzz5t3iDfSFU2tHIaVplzSX3QEprYftbaViBGbQLwHGiYx4eOpHOW
HfgbE6LH75m3byD4e7JKxD0EHz0TTTkVbEwvu1ap44uDZcLiNsW229StNKW3AHh7TXWDa1wcWNDe
W8k2FHysRRRmTza7ZdA/lTMZJVqeB0E5nWEO6WhmOwNgmNyBRci+coycicBiv+dZk2+Zqvh5LDrK
HO4+GKXf6nNyo9YGEzbdyMWwKHFn4+AYGa81us0oIn1nJLYbbv6HbgMzXdwdbhglIu1NviqhYyYR
KzR+sToqtslUVsHsXVxNPe2rCEh5NbMl/24vLKXYzt8LrLAOCZpf+HNHB5vWHy8nTZbxosaZdOTm
DNIfowz8dhUVgG/3UFSI2JCR1Tnmyn//6OXZ2P3Gylirb+lVyyfJlKLmGqYgL/wwEIw6S30v8OvW
6kLp83Cs26naKWczqpXE0MCg7XIlTQCmq43Z9lne+opOFCZU6Zoh6RafxO8VY9wRFPOcns9VPQoj
8du0VHRXWzYWwPkAYnmtDdDoAVXfPw0sGi2rnnembbAC5tVKX6FqdgdEOd0P2msPHvwOoE0NspDD
vCW2HYkuKrxEN6Qi1Xiit8TiX02WwGR/XOHlPrS6Xh0BuM2tIPSi5aTHRss9WE/Wz+RU6dA/ouQR
GQ7KhSXooWnnEoGRpLZuyKaqTmuDGExKGvBN0l63bnG3Tl2+ZF0WE//LXyDBrl1aSKbWO70vt68V
L35UsVAQRcDp0CMiRWw6rKjydxxDqxslQp4dhTo0fNYqWsLK9ZY3FR+aVk9GFxBeCnVeMjUK275T
HA4qFZ31nk9svQp/h6h7yeiAIO3gQLj+YjVhZzFIW4dvVvcPi6q4dLdtpZUsAHV83k3+8lE882ec
9BuqjBJ9IaYVV8D/YO7R3zEYMrRJ82w2mwQUP/c6EyWKH71Latr1Jc6M16CYH835tmLMrRObaghT
nlco+IuN1Tp3Agndn8ep6bcvqMwFImkOZhit7ppwyCXh1eULXes429qgWe05RPLtcgFur/a5yqO+
eQF35hFM8eN2V1xk3PG79hi0z1qFvbxeinMundj5rvaZtuHZUdMcsNc+sPQqqQYurptuVI90PMSb
sL1r8CqRMGCCtBE+opc6Edli1p23o24QsuwYC7rqBg1AyjQGOx6nwSANQjsW84Kwo/WPPhD8Oa8d
lY1XzQLHFjMXivufEq9srkgyVxp9KeP+rL1LmCNQDzquBgNHzll3YOvv7tJvMoh06H0yIGrB4jSd
q01bILPDNmg6kcqR+Mj8sI7ac7yGc/Wc9IWEwgBOdw1sQcTjBq1JAONYjLzzMQjwL+5Rvmv6ZNc7
xjLf9xM0I98NcYz/mCri084mC5braD1/JgL0CYATmf3hrKnentHnWnO1BITx35WTZF9OYh3QYQ3V
chCKgJMGEMIKAFGEYAplAYp8sklJyb5U3DXB3CyISIaAXjEDvFeTR7oXPlHBbMHE/i2H+XevTDJ/
nyoxYrx4PMVIXfy61kU8BH9wXhNRKSM1PfSdI4QLNeqPzmWx8V6zkxhUBN+ROYjiae9X2tZxn4vR
aVVb7xGe5YV8puvJqlGqlFmBHUhVU6DYhq9I1zdmhUIMwMjFuLRL3r43SRZlh66wO7IMkLJH3YFk
ZndR7GD1W1wRJF5Mkhv8BUZcvK04i39oo3vT70Z5f1kBZauJFjBH5pZA09SmCv8xsA57KC1EClMQ
k0cYLVhyJOjjMSZxVw/PnSpPcgcXZUkabT9qKKA5osZemgnSUy5jAeF5fGvIHeJBWF5782XiUu9a
+6IGVDZT9oMhyyOh3P+SYwbnqcwT0kz5OFyaH7GPElPDIrv49Sb6gHbvwO9pErE4zGASHMSmV4ws
yL+BcMm7xNdPRlHzUVF8ohtYBm++GeqntXJuE4CiFS1IJS7xlaijkuXCGGtbnps2DSdL0SzWqy4i
3zQu1spuYKkNwG5EGZcwbuWVg55swfRt1T0HjTDhUc0UG5YGC5ETEvE61XL++lp9J3vOrtvt03fG
ZNbCWkEnPqC47XQV8AukihRtcYJIMDQxfYtIAWUh1tDBFDcXarImszt+KMO0C8uodGdcZ3do6gqx
XDeY0QtFRKIWDHjnaPNdBZNDmYcWEuA9rW+PH3uTTLsO9vKzWlyACGM8RkXSG+CPerBJbphp9KFP
AET5ZXh4gGaMs8ZfdnR583xIxQeFqjjCdtRM0DrLTpTM9ZPgd/iQn2kkaiSmFqbiIBcFuu7q0PdT
f2hFORk99iN006BhqNv3DejvYeww4KtEbnoMJkalA54JByHen8J5TBhARaRzJHX6yXm59CGRsYCB
XGfSg7w1IgNxWPLk8kF7HzpHFZ1pC1HRXOdWJcaOxnWh0NuG84G1JxR/ZfejdsLD8pbYD3ZuKiyF
ZLhn01t6smSoq2N3Q8uSPdrKTX6Jrzxd8G4nEzILtjAUsmH/u4BQUKNtprcmYBEB/kfopso5YGVs
11Ytk+VK3w8xb5Lo39L4DLi31N1vC3dFXgB3JkHFZ+OT8c4NCHgSzRaiunnNRm/1+pe7ZIJz6TAO
CWS3re3gH3AH4x2e8HDhfCwMqFf7QO3gxuqdKYHvi96XAjK2z3BHz3P8tw3DEqMWQczI74Wtl0TR
/h2iHsAZx9Yw0n/fWYuu/BHhZVYTDOft5Xlj3WOjVnXrGWbEkan6KFcK4DCDDCZDAmzOIp1zF4fk
GfV6X0iOuEvPgTs2b/WI7EIRe7oDnKrKSUXeiIdV1AS8PIE7XO/VwrjGNore0APFI0WZDkJvrmbj
JnYFcDfuLHq1AvH25snp6GN3yDq5LVx+J43yC5CAd1CmujiXevMVR/C0x2nq8EpNNJFcFvrkCCgM
GGxcwih9w9VaDLPUIV9475VP+1mDuANL3q1zS96MWO//90Y+cQgR0X7gFOdSs0wYC1WYA0Xjv/Yj
IcILCCYzERbUZxF0qRSmuyGKVG4/zvsRyCdqA6qfKCel4ax9Th0iQurMCtNgnmWtjyXsUlW85yB4
nJjjAC6CgI780flBUGgQ79/jCRd3AyOaYrAs8wi+hMpTOwaLjUYu6543ZoDrNe4pvrFN0I7awT1S
4PBJFt25++89/qdHI6Fz95KvejXJgzrCdXxbVMX5Jwv0dpKzByDvJnxUn0NWs/yDRsRlGpm0Yf3C
/npmcqNpdprF30iLDfOKy32cY6qpKBz313AqG7B1t2wv0qRQrbyHgTChHxhBxII0yZrXdttvCJwv
lYU0oto0CG+81P/WwFhWEXqDbLr3p6Z0ZLb96LoAkwzkJ+6E4GHhIHa1SGIUi4Y/f9bvBu3C+ClV
eYQEe7xEvRWftVboohScO9L+/C/kEwf6fKr+gXJjW47jAx1F/cDYhy3xcPOqJKA4WjVpVhQQFj/I
POEFUlCMR3sf/FvzZNzZ3NiCAeampWDafJYRQID8cYL85PEoVOtp2/P2Rk2rOwdWXAFIzc4+M82d
WV10cLbPkaKvue9LgPwgQOdVmAmb3ZNaDrnALnQHAT32lvcgchpVzD5CeiuGVDU+S7rF3VMEUQEQ
aZ6sA294IWBiyyXonJjnU0b597S7+YAz0t4VgsOAWz4S6IX9rhclwq5U0lKc7IavSHbDVKg3eE2d
efaoJA/nUwrMVzht/ALDQlOWmR7ahSSoM8eEKcNZstuGASqlMvkp5TrgRdUGqeoUp1xGl/jk218m
fptUPD/IB4AWd8go606S0yIX6EjQXZ9qUXZMSZ002ADIJCWcY4J79i5Rno4aCio/GVGUtQLA0hDb
fKIsjolnc4FFms5uvsZNzP3dHpyHqo/V/SYx0Oxpk5OFOK69K+xFlq/nLvbMGCxvmHQAbWbinr90
JcTTcLlZFAEC03y/+2CCulA3oUas7t2vabXiz4Y0pOlyX24t7dFKkxKdOFowccEeAED2nhJ5N9ws
rpROV4VAPfJTJO2PC+gjS60s1nM0+ZWY49GYRHNp5ozHSpC342A/dQkbzBsyE1kceb3ZXQCMuMB9
7+nNyyVxaNHGG+Xmc57PcL3Nta1WApjyHeql/yR2cNVR2zj0+FdYXHIU9iLwKcWS0kV5SkyJSDFb
FOI8CyFL/lIEcEdxvoHpLbxamd4OpGCthFCNgRV5r2NINLftKSgywTmb/Axtb8wRhCFJrCnQeFb5
CMKcC5gCipXUSzVMz0sBgIpjb1ap+l5J1JQrXAhlrU+EdpZFtYhFKFVm+axpVc0SBeIK29B6gunW
jjWFr+WGIpSQTB/0JIdIC2EWYlWGkX2Cza68AYht2lFi0/+b9difUs/Pt926w/6jFTu1KOj7Kblx
QVxU/wLsawo/wl79qTLw4T4aJK+anOlifmPxd7ta7gglD9ncMMTZ++Y8DQm8XXOL2hkko9UVP27h
PLa5WRYYL10Q2poECK9kI4OZ7WTm8q+O3Bxs1j8bAiSeJH1IkAmUw+9o7MJzTODa6D2V3i21RusA
2lWPGySNE28DbEAFjUsnQYaC33KcsSpEbQ3C981cy0koWf/+IHrwykpVeXHTOm6oE3aQNpqIlj0l
Tb9UsMIsROVFRRG6Ur5WT9egza/GisE41axPs78kglC0pC91fiJPhQKWXPl5fpsXPtMAYERWiQzA
vOhNXUXO1KW2XZNkpCwAGPlPmEMm2/3bYdwvwgG33IqZFHFgdwJ9w171o+v7Om5ZARnu8oyRduMx
QwJCR302QJC2Ne161kwyfDf4p5PMV/c21rDrX7GyZJjmF4gPBRQ97e25+RwCeAAuDaaULRzcOKoW
2+QMYaKryeugFs5ysubF0tUesfgedtBb77CRPVt4FBnhbYPPgkniwTjbyktHXaOj0bSR5wXL6cpC
hyKouUmqnN2N5pA9lzJ1oFmv4zjZTgoVM7cw+Cla9FuVBr89IzELAIpfENSZfNcwW0B5OAUvt1w4
XC7xkLRFT89WAbS6WAzQ8Rh162maN71aNrfQLcLBym/4D2D96tA7hZp+Sf1yaaHcqLdKfbmptOaJ
mTU2lJV3JWlO7q/+3oFyeqT+pREnDbV+ey0PrgXgoPZXUGQjRciJ0LxWYDGAcPgLFWwjagVvwtpL
AS0cw44pw/S9lyCEagSPg3JUflLSdN3h4Nn//ARPNlBG06qrIQt9CXO5/gssWDv18+rJOecDeiKM
FrQjZsVlrdunCCwA3k8x1vVu0nHtSKpH/gbRUzTZBHb/sf/4MSUNwJemlTzAg1Y26XSEh499StJn
G83Q2frAlaX+9xhn8AEjFsCKHRK/VTQfuXeJ7TvtI3u0l/aGnrt5Ud5euzJKPdb2JhzB0tdn4aW+
C8yFZMD+r8KeNCsK7TKu4V+YFKsIEdVaEmP6gX+qPGEizmVfOPpYJo4P2JhBIMqpdgegnHCXBYgA
hohnhxsPROdN/NfR6zQTkvktDdnNHBke0F3+rVuWvdx4jnxLjlIbyD3Dnb7CgstQXKfzgy8KaPx7
1ELqPYFxZhUdbR3YLKjsKvruAg6h3XkvSj84OFsAjGfFKdvbzkSBe70k9/K7mN+nLuwOynVoNLuC
8KFul0B6oY5bEf9fztQwzdN9n5TXBMPveLC3vB/poqVzCiq+tNdl4PALW5xZOESJ6WagRxs+LSfE
v7z6ZQdtIHahtDUY/m6kCcjEzXu0W/wUKymfCa+uAyeQd+6SI7EdRT3bVchc/M/u3DKf+sS799md
fw/ZT5dV8SiHCi2aa8yh/jWZuP0Oo1njfu7SqwCSe16xxhuRE4LovmvyKOvPGBFPH38g/qqFNP1s
tNx89oCvQB1iO89W+n4/pZVC/S2U9tZyiOwifRNF17UOAJK9EYRty5bZztg2iIC5mkiKfghjodRU
0KoD3d8zpTQeUN93x2LFz0KwmjeaPVnWKq7PZgrz5+Z3iZjo+GBRu6vA4KYgdLqhEP/BtEvVsdYb
ORgABUV1AEtr+mZghhhnP0y/Fn1yexsafBqrJkasa3rlfM5h8oB0M5nV/d6GDp+OVn3umYTeBWPb
GpIjydPi4xALPvfsBFa8DUNQG1aaV+sqH0FHeiFnp1XMRjvU9SblL6m6VBkMigQ0VO9FqKWAZCBQ
FpGpieYBCFpy846OqfA5FNxkRzb2s13FtB2s158L4peMI5O1+vA3ZIpu3mEcGEihhMutzK66qf0o
6y3A7JuluSdxS6kBbLINJrrDvdR6XaO37zQqXliVpYXpAebn5rOHHJWaebHfViHMXD8uZ8px7MwE
8nbzZullpzlBCcHnD40WoQnm8jL2+gVkvQyFCfCayQy+EPhyz1ZQqFYi1IXFPW+c3cUWTC+EDcMJ
tSNbI/Imwg8OiqLMMybwPL/0xpeB+OFfgGUuclYYVXBw/3n9tVpwPJlxe28KP9kQp79EVV+e0+tt
7PW7cMOrJViZlUGjnBxH6bc6vrFZACK5zJzKlb1jcvW3G38qkrQIXXTtgMww1j++iputdnxIM5QA
Fo8CejsVHi2vB58wPeg/3e9h2KyNDn752QSKWrVp/wVHRb/RzXrJFt/Pos07L/tSvwLv9KARTyJp
Yuek5A+fsa5fDEz7HyBl0kpcbm7ozshLvCWkkNpubCFkZDA/PbrqaXIIPkEEFcPIZ29Gue24wG/8
ytbLU3h8hqnw+KtfM8xEO6jYyAZdu1iOx2/hJFDXnYbpU/G5UwXd2pK6BUVUWn6sL0/H7ulqLAfV
i0/jMw8PPqoRFiRPxrjy40A027cuVhZSrbNNcDaM3WT1cGfmtYyL1LQiyTQsY5NPDh21QtyQTRwl
ugFawRv+gy4KEHZ08ONoGndrmVSfR5Pp7E9BzaaV9IpPOJdw6LT3qBGduuzjDyuLNEP2PBA8WGL+
KSVpj7ziIOxVzghLoZ+qnlXXR5LpWUYhmUrQvKKl+zLbbx/cQXUj/cAjjgdVArVX47M2Bu2iHHVb
Zuz/V6BDVPflL1Lm9aomicl2PKmAy3I2UOgYsyTPiCQfRppH3eZWIiEyhXs85pmaDgwbhK8hGBc6
nxUeQsJkpWpBreb99umdFbtsnLIU+vtO789xppw0Z98szutJgi/wqXTlNTwJ54j6yTazsYz3AOCs
ZtFkn/yDIP1heTpB6VLM27x2hBTEug9Hi/gMCWdB+vNY8RG06D0K+XHduNfKMn8aYXhsMjvqo74U
m+EQLEzEK9jwLyy0KnUCCr/FcIHzGpgkYzxXVMAWXgrciG1Rr3eOf8jmKMGOgrYO/oMDdFTMYDkb
bFX7YlkaX+S+STkLWQCJuAmZfRtZV2hLxOIHrmhULtg/tJ+YEOMycrYOngwp/E2l7xGfDkKyHnkp
MIjne2EUFXNkmB/fy3uLVoE3o6kYj8xKgX5xZOV2ZEZPvYYYdJfrSXVcR0uTisnMtbmjaW05h5PH
YDg74Oq9Tp4GmSnjtjgsKMyLLu/bbEnJXAZkV5MyAgtmH8dDC+v0WcYWdM0GmiyOX2Xl1B6iZDBO
4GchryEvNfEHCXqIk8YYZGvLAJMqGKcXsVOAch12hy6/7K+XAsvtdzQ86Pz/ihghnO0AcI1P+agv
M0ARH+0X0roxbJ3AR0m5Y0yEFNXMWtrQdqG3Y5pEOlkM+A9nC4yzHTLNk8EHkhwbQmludcCAWtQ+
HQj7lnLH0vup22MBZaCjFeFDkZtEsFwplg6csbcQebTmEdHSvXltQHFCGj/4v4Mkel9um/+fBDa1
GGxDVXdVnm79ACvRrEMaUfO+mpfSJYmzATD2UhI3wm4YAAqwhcGmNF+FdtgNDSfpUMAoo3V7QWN2
iBZu7cr4KQfh2jm1ugLQt60SK89nzIsONA619Kwt8DFcJ8qooopxiNVs+51ZSta25+s2oDGtGm66
WWaTeOZrZnw54V6K9NaKAhtxRBe3tA7NfPnPWw897S5KJYitPT4MFqT3hvUotsNWyFIZIa/qYjHc
wwxJ9BmP0BvWmTmMiQRJmtmsKxzC6JfXUwGXdca5az6Z8Jo/gOfVJoy3NHNodYRc+aZ3Tj+Kzr39
AVk7QK8+MbN4WQTvv5f6FvbWsKdo3hldEcFHDFbuX3BpF4IZJM2+2is3tyAPfg66CtXGZyri/Qjk
LhFePLTGgJwLtFUR5ePD+Msgmy+2REukmaSMCX3/UhxE3w5v9rT9q8YWjjLkItqr3W5GSA4CZ5Ni
Z0lJ5MZSfbavSZvo0hQzo0vohhSWe/sMXUVe7YJ5xnspw0aQlS6xFHy6oHPVgEKh9snzkXck/1SG
oT/gwPRDlxuqIEKTneLw+uXhdRlX0J2NP81maMB4dQ0B+3qzetNfp/TnVa7MkzS3l8u10zjTj8hv
bT9QC0RWkfwA7boq324ngOkSRd9fuVE5K63jDnnoasA2Ge9U/5bjeKibDIdyn6FNQSMt2+x2G0tp
Omy/q7qC6W5Ve9Kq+1bS4WMfEsjrMdoL03fCS4doU40hYpf8FvRzR3pErs2uTHS9LTnUK2G3ZQyg
7zKIRSuevIeeea59SKFWuS9txR9BGsZjwco5KBIGUax0NkuyD+aC2kKesn0WvtpmHqtlpNgdqw79
i9M7KW7y6q+5S6T4Ej1RPz3Q1KT227cx7vYvWZ07PkUHISEzQI/Z/+13/Gaj14k5NIWFPA5sYdie
UqwcnBlnqXurhPiZVe5bwfC345Xn6TRT4slfXGMehmi+1xJorW34Xf2yNUvnS0IQY3l+Ra50aVN2
G0KEkVhoGeFgOJQRidcRgOgjh6zScG0SYwcBNXzi87UHTKwORb1fnb3jVU9ilgqWDI/QLGxCR0eZ
qQbwBzYpry6jfydRSBW8v9nnkKwlH7Ve6yunO3ozo7Md0W+zzves1hu1Arx+K4+5nen1rB+deQ+k
Jrpq3c9iTymkv4SAlJm5hevJwueQGSmJ0ScwcBJqyv5AuqolOquVKC6KdhqjVEKYjiK1tpBcAm7i
f/VvDg4UiAKIO7ouT1Im77E2dUOcOMo8JA6tw02pJEUqL/9nx+YOqOMd+rn50SXlYFO3yQuC5EVc
v0H2gHpZcXdd642zfoUBp6OEyEwG5b1ltz1do4FNC9PLHf9Uy6H9Isal2D4twF/XQ5Q5z5JkNH+n
3anVUtAlnc/AJzNli1Ret+5sMb/vgys5KnU7/WsaL+j3iKvLnWAuw8bmylFjlmNfiBtR5S1ZzJW0
cQIbY7sQNeLEMxBJhhlY/r84QU46EWkYxykmasoB3Oajz5vjBYyboT2ino1h0aiTWKJGIgJbCQky
xRJYKMd0dVFfvkxa1m83eb5B2FGU864gdw9JVmWEBqhmyAe3RTcmq5qBctkHX/cEC+tL86MoOrJI
Ituwyfe+f/zjkMv5CL0EHV7i7agzlNjvRVS3Tz/EytYgmOvYyFtbp8lOp4N2bD0BSD6EZMNR9r1g
CTFrphL8jXlT1GvIfm87YjJ3caT3ekpN/3L9g/hoi2YWtYxml42D9RRMbmogcuaYIy5Hn4ZPMygM
4j2kSYQxSxFSKNvdILd/1Fi0tlHF+xKBShBstMmVuG8uP8lMFPUVvxIxfp8ttZPxeTkUhH/QLST3
bFjjiCecEf1epcQqdiThqcw0XFxdVf4Oo4g2gkui2Aj/i+4JUGukSbv6qcrLFv/UOgrsCyGyYyyp
jMJjK374gtkGCFb7h6cf4vixPppE3Xq+AnIdrrABfvT1gPmFJtvd260BJdrm2hllXits7YStjXI5
dc/v2Qe5KyzMusgL5rkp+sIndADUt8n/ZFlGacS7QvbSfSrJSN9zTUszvIo6KZcF7CoTOPTId1vT
TYotesLahTFoM375HdSsBg+DJ5rGd2g7tqTD5QFRQh2gFsoTvsDu++nky3iN0e2l3n+mExUhr8MF
9xQ/JUoEuMXPoLI6a6T+VZq78k5GL5XfVM0fh/71PEbXeqXNKT6j11exrvGWkNBZvYetIQfT0MnB
mvNABgT67A1GsEuxCMYia7UDYXjG1XRYpWvcHUtVhrNmXfuwQqyRqnpwhrTX8Xn8IQEFA4rV3acd
YPTVMtZ9PRbiooanMiRo+KFHqACBXwk7zpEDGchyRyzy95+L/QHdIekviZqvXYRUSd7jcLVSvyFx
Echdy5xz/821vxClxaDj3/ayLnMdCad7arRbOH/l2WWQKeGZETcgI8WL+NUt+uKjGc8gFe/zQdqG
FfhH01o1QZ+TvNY/ZaA6X2Dh2mYb9CTosTh+95PVLJfwFvF/hhTYDa5qxR/xf6ZHLUFIGicy9uu0
3bNHefIQpJfJaHgxT6MtL8dabxLfPP23YgT7is/cRVzShdbZwVvnMUyaa7qSALDWmsFz+UGLiVvA
QADPGCdgXiPQIJJRa1LVbMyPkd2WAhRerwtrKQhqb1BzfwSlga1gTgcTA46dloWNzQo1/yABustg
CO2ZNq5rA46H+jjZ8aAro1ZKdqmjxc2/DI1SOfYpjZcfMT9HcsE4WaTJ/0w+GnT/k9LsF4AM9cMw
H6LUg1xpbJ54p0K4qFgo43sWRjMoA3YSS0o7mHy5NX45NOU3Di20ry10BlVSJ7xPw2a3MEaIyd4o
OEdAAF4loRI5my89drnKuZMk/qDySKWvIwSwyCWEpGs/D/sFuCK+pcMbbL1LqDCMY17sK162ceoY
105/uG2O/wC0i442argLNRC2V7Uh0hDGuTjE1JwDoBPBD7vTVqZ+M2WftfX+UuO0A2yaUQFMcRkJ
J6CEDUrvbWJIKtGeYQ4p3ebmN769hR8ZHafLpr4kBdN0THYWaazilRjpsipYOkxNlf2E6eMoUE3L
p5Grh6R5S7y7cxHJxHFhNEtHfQd1rrLaG+OHMM5l8zRkQljtIz4cO6/ejzndk1xunZEkstoNbsiq
CINasGoUhhhKgZmpLrmRrlwSCWlXRXD1fHo1bIVCt8w4Ji96vdCEyEuCSAb45257SWs2DEYlWBmp
6WxgGwGQzj0HH6WBNyCS8jeC6L7okFeebjezVNV6aBr8Rq4Iye5UgTbsje5UY8GzIFOeu/RALoMu
ScjoXDAJpUsI5aLHpphNNGMVHSSFNAVxgA+/z+nrnr7uxZugXHC19lq8VayirpkUCi8/U1AUHWsN
U3stXKKyXDJ87ug3yTbxV6JvtePlL4aS1xcYDVe6xLcqwgZqear9oibt3aXnYB/4AoQSQ8qy+PkU
Z0C5kLSmLCal1oTQ0RYPFb4tp7cd3hRCjmMXbeELnKr7YDFPxXVYTNQa995/dhq+fKhZW4wriB/E
6CB4AGmbuWheu2o1G5fERAfPtUloTR6XHemXFGqo8TLIH36csujEzUMxICVzOtk8TO5ktyeYmzIM
HkfNL0iS+rK+Hyqc/vsjAyJcJtIcobVQJsCWAT5cPlo3UnYCQ9vRZb2Pcd6xhtgWYtHiEtXA5S8A
ID/QQMK9ui6Y5Nw1miw0x808l2Z+43Zkbsrgu9d0vmFfYbBzLCgulcLhJlDkHcfV80iORxJoKzo0
j902RDcTdj4RXm9kswxn1+PuBo7BLZVe0kg9KXpDTlmybdWJS74zue0QYeuSdpsAiobQcDxXX+TI
RjAojBCXfkv2mFeGiJqheAmG9VfdoU32fdyRN54SqTlaoo20xoOK2w04iPPXL2Eud87HpdpSSABi
ZDucNSbfUFwyCwFA5pGgHMw6cWzS+U/k4nd8wHVZ5pzqBuyUxbi/MrbEaY76Wqa9M001XcyFwIfc
AC1nzWHFaVVItl2yXHdEFfWGwBMAipIQkT1W6b8cLCL7cQTRO1otdYwKAM4EQ8ZMXq6bYiZRb3no
6MkeYEvxwpVikml21Ps0xvflTbFI3asi9iELWzsd2ZARtVq7LlXBt8MRKFoVnAKgXOof2hzvxBnV
xXbcX3xjdkzhHvAr2yE1k1a9L3TPv3Mpdypyt+BmOCgAaaT6yWI7hoR76jaOAvHCUxNSKAKfolyX
b3NxikMqisAFOCnv1BBYYH3cDKdnmbBN9461Wu8CgpF77fpn9DV9XVaqC7PlpDKfjzFd8nDRubXU
QHdK32OXkl3QacAN0GBdm6jU8JweE9yJmPExpnYAlWXQnhrP94R757HbdHze68to4nY2V3E49iLk
X2VmoXoCwmtnboazdfYrLGJMnCoseChflITXW5vXQrQnSVaGHwemjrM7FkYj4pgrbLDB2Bs1rwEy
Rvbm8YZmI2U5Vy0Z4rhdcgLXro4yD1YPlSYNXv2NOBoVbfGdzTWWAuZRKWO2g7jevSW3ac+hT4x4
ofbum4WhHnB1ub0whizYi7Ff7d7MnCzD4M/qeb9hE4hd4FtahICNXS9hiyC931oYwIfZ09yEIK/l
WH6VkNkh54Ck4vJme0trEh5lfCoBCBoHXztWLCUYq8uGCZ8+Mi6vESh+x9dSu118zxRRobo3VI5u
UMOE3GzHZfMuCxiEW7ohZFd49bU0rZjUAIE1bCcaIpbmgqacR10RNN+1EQorM+X5+UC16/hqmOQN
GqCRNo6WQAPy5WNqpAi0IXeKmQbmJ9BBZ1MSl/k0/QWe+RBTbMRqfka4yQc+6R0kbAbEwKA1ODpG
p3jxQbAf7CbC0BLmUZrkXFV3TAc/x02647ZMbcaE2uqGobUFPZRrnJGiMBgO9HRIzwBwh/tzieBX
Iyd+2qXwzXWtr7L7mPubCmPwexbsj89lhxQkOxR4AJH2s8f+AhwX1pARNLD+4cK+hZ5zR5amEcPO
6mNo2P6V81R0DFwUjKiG8Kn+itX3uWDj9DI79XPgh86NfuZtuDG6NJQlUAYUWEgUiASWDadl7brh
5MglIJpZNrT401cz0IVtHWyDrPteVuhLs2XMD088Nt0hVyQhSmR7lPkTEOVcKNJXj+9cWVaV3ABb
YmWap9AyRoiWFYXy2/9kbe9PbSrpQqQlkQBIEeG7/YwXkv3j7mj7/48yKmmGTS3HhQT73EHT/QT9
dZP2clT44Eegx31LI5igsnf5iR7BEbgO/xdshBNseotXfeE/y8eeM1jKtY+QHV+ATz4f/FgRLCQ/
fs8ZbtskVIggIuteg2Fec+ESZSh4p5rraX33xmiZpoP2k37eoqEvp54MIRriLkqOYF9/U/H94GP4
EnKyplIX09o3gjNRWpkUfspW7h8/8nmJIAPQ4E2A/byACH8GWA9nuROnM49497VbO4SHn3q6QlT5
mXir/tdyhTF8lu4/7RgXLIwYbTxgMEqa0SEcF4EM62F/Wt+r2M+Q6j9NegVbUN2cGCZ46EJxpRak
2DfrFPsjyEN3gG40J+MyGmko1X7bA0uNkxwrsk2/ExsffZUwcSE2MAFsHUkw3KhpNxm1AwwsOtkE
1XDIpuEx7mWx/fMTyXVc9NdX6qgAC3Q00u1BOLVHvswVIyTSoLM+XymRhFVlmlQskZqBBHIQ5nO5
smaGjFLz0tCgRiaNWs893zAB/czQ08V27nMA4BSq/r03VkKWITbhvF175IjhHAg0VQOCOBD6QGb1
ARJJ2eWnlM8ZgdzgXNf13qjSqWVGSWlLVnKun+TvK5hKmnoJOOn18hwtQ7KGt9xMeMwH/EI3WVxh
uVt9AFoLI3j4RMP1djD36A767N6fYS2CqoCCMO/F3W9wezgG/4G59XNfc22blFmZSCx//keMDz4W
qIa69CTDvewIcc3fLxDpmO5cASnlVjTb79+KIWetavi/mfbiL8IrQmflAkW10FYmsr1QI6S8mRgo
yq0Cnq3lwXFM8iZCOVbLxl4udCAkOlHK5p+7uMdUgbyh+EdA1xgaAqg7kP47BXiEq1sscjdQIDkH
aTk+35AaBQmWNkwA5EJvgLTTu4Fo5tefrCtRCNFpl7tfbx5y7ZW6ZN+HRbo3osIfIv9zqI3MQpda
UviEb28EhjeJisgXY39lYkM406mcJLGGueizMg8MIxn/oUJH9Tvscmnaa3tOlF4mC14pgHZ1NeTH
fUTpZpOSfouiC4tEHCoXxDlbG3YWp1j1IDF7bmE9PlJaFlL5Ow3gARc1t8URjlpltOUGTBlpXI7x
Npbn3cOFe+Gwe+w0jwLhaQB5nOnqCo+5P/RiBfmUBnH2co928iNiJMw0UywoK+eXRJrxF06c0PLs
9tqR6P09EBYR9mGRD1sZaQ835QXheFV8IXa11Avor7tbt8IPH5ToH6lFehIohSLTmu1k9vAtn5n1
S9utrZIVJZaaQrogZFNwTOj3G0VD43kasmo2+RYqnceOFXoyaVtPHGzJlljqgNELxInX5LYCNBLh
dzQmcv9GbcneMAfNj+N26SGlo+smwd7eEol+1O1Qu01RLhTDMWIO24xnLqy9L+iipBCNQ3M8x8nY
M37etgoGZzBb4g2Inyyyvh6zfvqCq5awx7xo0lUJnTvxtFUYZ4MzpZRCnuI8mf+se3qpsWkTwMP/
ITMCEFddS+rcraktFkh3qi73bd7CqJ//OMihzCWycjOpF/LkAU7c053h42WcrIlu5fGQRIKWxdh9
vkelal7xTLGmfg/mEvHddbUSdH3VRhbv/oRzpuDkT0LZ2WUScrXbjvymNXjGbwViL4bI6JjO5Js1
B+I3WVvqAJcG7PEY1YnnMt5ocL8UeoD+dwhQ0G9+s8K7/XAstEPwdWeP847o7ep0o+51v3pvzKOW
CsdcG2hMCmBZGPtJ/Tk3kbOm8ZYRfwItqLk5jLb5XFFvEWWErFYO7z+PJPedlTz9gRibPNR+5aN+
sEB/SLSTbTsptA7uJUx8C5TS5bIeYx6AhWOueCwhYimc8FO7CNWZ38TUt7o3SAqliTbEyn6uic6S
w0rhytntdUZ7vb05SYqUF2bQiumA/cSm+s+SmnPM1Zyw31LK61iJgew5TxXUnt+q4jYd/Wo4sHbJ
5/Z66wi4FW8aVVCE0veBLQGGkAtfNcmD7e4g7hzeJP6Ih5ZLRgeT/OQKeQJDF08KXEg7VP5oVgqu
DTCYVEoTQhDHoELmqPT9GdV3FrHyfoiL+F1sZF0dQe4pOBV4BymOBPuJtgGBaRB9XbKIYixshXgd
AZS+gnuJqsaXrUEKtEm0uNKflyLV5PYn/SYj8PajrepAIflUJTc3YOnpNsF69LkZwCbXERdDez8C
+5j6MkuWOOezjb/IbC31jZO+zPV1C24VQUPT2qebnGWp6absN1GZSMmeJOep0BNTZMsU8oEtwdhM
Rlf5C5jww92ldqHR3rvHxUeS8o+gO8o8x4H9TRz9mPGOgWQj8RhIZk+XQrRXlh2UIScWsJgC1kkG
5KXz+9SNFK38ucuWPp3s3TZnVONhZCrgJFBT3SoOJEGFgHBWi9h0v8cQgkQ58uMZ5nLJ21g88S3f
37F5GbOHDIvcpvRmvpQh5XiuqoLWhGI9PlbohpjMXBj8W6cxdDV8Dd1KofqtXIpMtxsmatF4oG6+
oq52ZvycpHwVFrcjTpu9itFsXtST5KL4rdniGrSgrTflfonGBE6H/6d9Ubqg9FO7ihM0DY1i37+G
m5yEm8FAcM/4me9LE9I6BuygveOzrhYUIW56Qa+hNbYWuWm5uz5zNaTLmZuyOnWQrjB0Mk5InKF4
xxfUX4BeCH6VF8n7VPRQTzKLNtT5XC8q8C/hPGxftnuHQt44MEf4JRTiWJWgPJwHT/qinhAMgwNV
fb4Br/+K3i/moejGq+1r/RetlTPwx59VdJvKN1+9Cl4YDnBhlud07vIGpVbQjhC+NxxIslhbhH9O
G8r/rpfAL1MfqL+dYRl90YlR+ltUK9d2FzzehJKRn/vQ5zzteJpl9f5zF68TZquhCX+GIwpwFgbw
+eOXLgFVtUOe0b1ONlyMP7ZHvwTJY+gpg/eYxblSekryjihjY5L1nf/Ko5UrbFErdRSZX/gzPQ4U
l1KCH8IZmpuwdvbtG+mD2dAQyqiFtgnRKg+NA0goAzFc8+trkO6j3sbrBdOC0d+0Ussxa3WWq/ex
CfzUHCbq5ItP90fZ2lNeC5ilKaHKigXU1vim4l9iEHbd5ZAhtil7rvVWAE4DhsPLAFo7FujWyleD
nLrL+zfz6dDdVcGVSC/QFHqXtJwUo6XMeExoSL+5kwcfcL0+gFkMAsZJNzEhGV+YQzvheYIDpUbv
WGyAZIK1y3045DCGGa7fOu/lmZ/oCXKgY04Wb0yEWREkZkrxHD+6CUT6eztjPtFotyqeGXb0TNAr
UntRwaRtxabADZFiQX06DGbAZOfxtrQSPZrAS1kqAA5j0p5VwmCm6n4/bEAoiZSjkvGy++T5fkgM
VH0N/H1GTAdkihH+5V3OPh7AJi7WWXgW1MlGwu/z+nk6YbHZyDvjNAmQJ3/C+DANR2pqDcmSzJsc
RteoUwcxoS9MZ/79ad1PhS6ZAdvMAcpLDxDTaHM4PabuU/6CnHMHrC5TZTJyHtZMXLweoW9vRTf1
Vvv4iweelv6TEkYfA7bMSLVljOLhvcJGt+Qou3SxjU6AeOyBGx3+uPQWz/nplDgKSE+l/PnBW9YF
7Tw8p49hkSLQdlMdJb0DsZW6X+DtCUttVKwMbHqXHkVUeqevfyTn0D8b9Hh78SWUNU6Qp8RkuUI0
KmvzHTyz2MWv7xPOv3dMCDp8Fvaf2TQel+RiSWlWKr1V8rbs2o+JcUEafG6Qd7XGT8MscUYfRRxc
oZ6+Gm0gEYye1192i++QfbH7nXAy1tqxGbAzMA0wJV0lnburl2Xs5urEB07yNLO75aQVUltBJQS2
CO768+d2kMzy6ZxrkEJnDHCnSEVU3+/i9+fVECI0nq2G5PyS5bwO+6k8GSlmAvis+k5Sbjd6O0kD
jvf5wezLiwoZBotcUpyeY6mqVxvSze6ti+gONLWDpD8ZNUDlMt1zkdlJFIOQrqMV2i9jjW+bDxFO
ez4n0XIctqotmILnY9SExo21+6l9MN21Bu3YYr4staERX6GJxg/wlPrQAHX1PB5WB2J5fZ6TPeTa
e4DjTwlUnudV10/sfkVnC3x3u5hTm50i51maXSjrg+bEDUcUt4KkFa2loaUtUZNt324yNwjXNXWW
dBZLFoki/WxusDoCiqcLEG1EwJ3b9nSzuM0x7UXXX6mnbmVi+9n7vINwT7cwdMvBOlShwfOKONSa
wEP0I8TSMlKnpuo4PKDpAdjUz7GwudSHDU1YdvtT0aIyDGhG8FHxBF/6AMQY3Ki/zAiqWzL5hw2/
O9coNlDUCXogyhA4U1daOvbFb7OhLRa5xoBuPE7QO+SbS8NxqesrCS+oCPz9VKna4ka+EfbsBjhP
nwMedECvFl8QXRXkZmevwRZyrXWZbyMPaWB+/Mtq3jjWX98D5lSnBHoNDVDOejYY8Lkv6AJnGTwV
OdTMshZrUEa6zuID3HBt94gFAdHZqJbl8NYvCw3Iq7Z+cTRastyeY3+lmxbmDMWym/z5VNvVJSlw
X9d6u7WVhto0+1hRUPlJUZfEpev3Od6CTqRck09O8kZLhF97+rxqQDnlnfmEhyzCdYu9rYFlwwex
2RrsTlrcgDLBLjhoPDq3lVNUXhEKSgtduorydTDUEuEfUtRkELpBB4zOe3aoMu6USv8nYPiZd3aE
A1tvtonkWLw1N2s2xWR+wwqo4jmROUUkiTuz17F9Fz+lPVwK8vM9daQOektlZagkKVV6d4ba5e3V
6jwNEGLHNeCo5Df8DdF2P6KbQgnaVkisdzonsgP88t43XX4dyCcmxHLh1tH65cyqaLLpTpRCyWRj
XH9ZqKA76r9FHEAuiV1Te2CnYne0QBw1ex8GT2J8rLBqs3P1VWw5W8YhvVFGTPVXCdtSOC0D/GKp
ancQgvibLsHgLGBA5N5e1H+MOsrDP12sBzuKrngjPvY02Fla+Y1Z5JnIgIYanVlF06msf79200GR
Brdd908vyE9tsBQDXk8uFuHv4htsmSgRr8Xgswx2zCQ9Bagc7MJ3yr+0Bh/gu29vTyTbkAP4OQBy
fgNLyGXeFI890/pBYeTBgvP28pEChYhRvP/J9t/HDh1JZ8kRMdLsDmnt71AMBlfcuvsTxKuJKeg5
3TC6tFRh+rZY7WjadAOlAyAupwFQFVhagv4cYhWNQt1ig7z0NwPNQ5Sb4OWhnOQi7A5gs560wyct
26HP2Gf8pY6bfP5h8Z+fBnya/LwUvQ6pWwKl7C1bT9OpUJr2WTcLS1lZK1F3Qh04Ys+ZVx9eOx3z
PoZJqyoH8U+v1SbMH/GBNMgZ7l/3i3D+X4WVVJmPWuOBb6PBK8gZ7irMYTJLS5PMBssMo/KDEUgn
+Fd9lVKW7/1TW9e3lDLzfAsZ7tgfIdyjZSBMu8seORXgINJ82rCrkgPq9mDFK6SuFxzp1nFBILVn
0KSKcwJVvopX7ZhrJqSItyUOZEclPq0st02vHzsFAnLZyav2CFqw9Jdvo6GUn6zqQ9FU3UZBoWjy
R63D2psKr6E9Bn2bmFqK1iO0KB6lNInXYwwsj8JiRU8w8IM+OYvYxtR5fcyzuEEgjsI6cQcJD3xx
8Is4qwzME6l8DOgTqQ6WWI6WNbGVLQl1OjF+NFl8YwbrwQc3Q2KZbxYaXRvps6wbvGeUjNogHIqE
9hlVCQc7ZkurqiGCzfZThOPCV3Ku2eVRxRa2uDDuJzuoGG3uRFuNViFc0BLkyoJn8EP+/Mkc2ZnE
XG3y8O39xSUj7FU9jCrhT3GHM5i4nIgcNeXfAKxxhzfSlQp1RXOlaxg+EUoMI9ltpwOPlX8Im4oZ
fHodJTH4eLDwV66UHZIqma0ZLOk/Hw5IHNe/EfYMYYQS4hvWqOaJNYWJutFe8iQXrLv8tgZBQwI9
QBudGMo7LznszojKk/JiT6QWdl8u7RZvG5vDZSNt/nWsoCsT/dMS0J3YHMkkRtI6C40ecjr24yRl
TDG152hdAW4yRP5utZKKX3SPaSUHVu/mPcb5sufjYmPIA8kP4j+BRLDOfKoR80DGVhyTgJ/YbePB
NuMIsqoIfOmEuxsSLSTfbZ1retmwbQ93cz8TwwVGL1b/VixOEzvd5TVdMZLHp5q7GkHjiJ5OBYmH
lHBuiwB2f1zUUzR1ftknxRCor1CmqnMO1+IXcTiJ5Iw6vLmxnDI3IgubmY1Z06eiUT5phuRqwRgu
SqL+7heCcDpCMxvNRII2EuV3BgFUgxhPoJpMrpIPbRU2eIEkrHkZZKXmBD7hZcsnrc5EA77L7MTv
diBZ9HUQBN8ocpS9E/aPNdaMDA5tUImveazvRaPRneo5v2OQY+uTkZr4E3ylfveW0ZLhHQzEcUOE
ZS6wvsZ027Siq2JCeHboz3zryffNwDyU7syVJPqn7jIgVvz/YVxkzIBEmez6vBrF09QzY9RtyG0/
HTdlzQp6xhqZilG861sIROxpaTF4BLlp+2vVUKq9wlK29McB3HwgcEhioxoT6OlUh0U+5o5c8FAI
cXQ7ad/d34/Ru+iyrvfXipEQwQZszJ4NvPow12efXLOYTQPiY4aQraz8Ktr79jIXiEWzouJ9AAHg
HZ6LfTrq4vASb/dVBj9Ntm4s/Xh7jtzIdTSp+XYGypJtwWB7ui5Ilw+H8C0QC0iaGdRTDp3Xy5iR
T1VJQjsiXK6nXNdu4YtUqDj9RFuppAnuSyoNGBffrxKq/GLeZXBrsJTIWxu6aGX0fX+ypUMX6RRC
2ulk7FgGX/tAy7jL9aK16BPyI4GMyhKf6evPdagP2sC2a4gM8AkZ/wTV16PPmegHyTykchmrNkHe
/O7ST6JrlC80XumaMtzVAPZVHjll5WjVwAPxzX2S7mevAlCkRzaCF+X4lI0eS/G/JxO8mLNypdwg
1a1P3koH8swTMFwyGNEQOdDiuEmkkZBAkAkzeBJjK0DdAHT6srhziOuctCUHbC2SVDStltR5vcmE
dSFsLlYt4wukcqIbIMyGYKPYksUOlbf0yqd5wa0Q5YjJXQInOLCzZmZ1rjrqZ/YpGm9mLdw3v0mD
BsWmgu7j2rwAQHg+BGr/noMZUwnj86XvTdIjxlX3bBmVqKO4PeiF7tfpYRkaMIiMOoiltdeDLKoH
7YXS1yEA5M3GchmmWI6PE5ePLKf9rjXGXBOUScVPcUCv9oEdK/jPTOimVSBSCD58EMI3L5Q42alL
G3Qw4vgdGjk1FSPxi2AQh38L7K3uzlXXCW9Pa9JE1dd3K+dabQU1DfYwH4Ecc26LzP1gE4XfxbAz
tiY8vTwtsGK78bR1A1psuK0lU4gLqy6wQhGMZM0q3puzEUGMfRo9bRn65SPvO9DZ99LGwASbZZSk
UM590UsQKVPummEJ9VmNX1AMrc+55Y8Mf8UMRfNs4YNPAuoM+nS8FgwURjojLH/jj6oRvc2rp9df
pueBMC414bWVxTPmRA+LY44VozDyVsfcy9kXICK9N/c09IkbNQ6Vn/ZNo7BQKvR+dd5cOUBVdKLw
qeJg09mvLWorwQajk/gMPLjM1hzuEXw92EMKOlSR26kLH7NHi9fsOtxp4qFSZhSD/NO3bs7thEsP
17pIjXSmoqXrdsjNTYWi6f6IrUQy0wLKqMRXcC93ej4mfobvvWAgjAIczU/Da5+muozw2/oBy1+n
5/m6hqsbjiyMRA49Ji3jijUptxbITrivxikAeROfESHLrXKQ/XlzAGQehSE/lvKA0/HxsHX1893b
9ICo2vDc+HLgtySS9JZREGYzXQmOAn73nf1XM2j9Fv+MFRRjTcKg0qZIsQmksdjpxZg3mhl7hG2y
M6obCoR5Cmurc8st5xgR1avwc0qIb8Q2AgL/laPEciwRYEOPAWc87SGLdjswYFOinFTQXIA5aXru
56OUGOG5gZeNqRyOhEBcSOtGZb2l5XzA3Zw+4JmGOmD0aPt5tP51faT8ahS2v+SaI4X+4Mp0z9FR
3Zu/1dE+E48x2LOWEOc98YBIjX8VSaBrVwYo591P53Qk4o20erkPju5Vi6CIZZmWWUVy95atAz9X
oZKBiSCsE6o0n6gX4ECu7HJq5jsP3V1yH2QObHulVzArNXthN/joENp/QraeieJSGcqiIe/SBm5x
kmFljZMvCSjZElWNcyTDLTGEnUP7CyGA7jGmCyLNcQkjvZz3gWE7p4SuIQy3eh1qPuXU4aA9lViv
UfwZC7YPK98IS1yyv+gYs02rcyMo0mlfUvy9R8aVGHmPbDkG2S39385bORS6Q2aaRAYaQDF9hCdP
drQWhgSHZfrvOXOBnEe01yIT5GpWlEWslP1bSqSvkwsKg0Y90Ppy5eni3I6MX1NEWLDym3lEYwWp
QEXVmuoM9x8xC1mKbxIR+I1TweW1pupOyIR4+jWWmFhGXR3rDWEznNll1LlPjXU1lvRfNjTftvBB
o8ityMGEE6sSe6GSk2HxRNLZVQkn9Rmttzm1LULQO/wtGjOKnzykY2hA7BOraQazMuwYIxX0oXso
gX+9QoUp3s8eWwJACt7myrKFHR2T3WBVmo6zKe6/6ga83S+MTrxas71QNrrStNOdD4yqat+TCVSz
0h30vLXPpTEdF2YMbUpLQdKB2esiNUTxe4N7VGAbCmOD2G+vkdpaeLJ6/1137fYAKNwY0Mq1IG36
CvBW2S61OijoTCKmkWBpwQP1mGRdIGxUtpvTWCnOEMUFRC4pmkskRIu8Mh306ZXaSiihqPKslehy
vleRZNKD6ysaxJ4tHph5/DH3QXYdGLRiS1++nmS84IaIcS3loQpPw+3VJGXthbns7awc+wEVugPJ
JKfR6vai+DMXsKD1+mtPna4Rjuk+01ddogrjQQrfyEQLWHFAZ+QdeLPG9+lzW4hplHp0T1hs8DkN
nAxLTgXyjcUBVmCeLWS8uBd5yl6RrulA8/pRtlxM3cPaL1Hk96jwGplkPv9gSkGm4wcpdnvKur+P
o5F1WqKnF/3CGDunDNbIithv7GP7/VcwYRHF5VQbiQaMdsu87fGRP8EYkKvVukWIvkHuZZlZJ99G
Yn5MunVojhMJ6WcwV2ab4d2EQUpg3s6rVKgprjs6TFf8iZlFBRDl4nrdy5YEieokAJQr0v4Ee6o8
3wtgzaxouX6KfcPVi6kq/jnYuCqBFr8qLHvBgLJad3jsoYhsT4CoEKfdwkB01pJufrRcnt6Ya1Mu
7DOMtImIr0twFOoExsYlC5Yye6eKzribGI11wXiTKSepOaaT0aTNhovX152KzLkp8Zy0B1LPeH2E
+jdXbkcLaEyhTTqt/yNlaHyR4cPe92FOVTEL3iA15zpG4iQooJ7/SOqgnOK2FxKXFXYWXRkoJLf+
MThSHZfwSIouEiZS8TCKfxR04kb/HFFrAQfNte+NB1lrw2MscI7sFUrB9p2q++NreGkURvF9LTUg
dAg8MBEY8+SA2h0HtWDw7qW84z5iKgNanvQ2OryEv96t/mcZhaFqLEEcReo+t+dCHJFfahydOHk+
yJim102s9yTBF8YdQXktXJ+NCAcL8p56goUK9B/+SvH7qYfI9Yk67A3SqjHaKSbroIgdBmR2A62T
L+NqmvjPVL85QgdcVkejwdN1wcdKOEMJD8A2pun3BqEa2y4sH31vaiczSLI6GnK0SvmNhb6q4ZdR
NKC0Ph9OGS4sfsip8A1bB+hJHb4qZ62Wl1h1bYgeGTb0YrXuYlnVOqZc0Tnr5wbmKINh4Ybc64me
msIKdbFY1kly0B/Htzvku1P1N9xnU0hMjcO4oLNpGCtG+m0jAaxvUvgdURDoX7k1j0JI0bdSoaHx
RqGSufNivJLQHhTX9vuIC6wxNO4qe1Bv2RcauG58erWUCp6DWv6qUO1fc/If1n6utDX8UQDhz+Hc
bB+3E6Y9+mYQBu2kgmijEE1SSY8acVf/Clmh15VbxaFF6GCpc7XXdr5LCrOQX91jmh0JHvaMN3c0
SwJXXIywG+OQ1hOMyt91mXc4RGUsQOymICti4STPoBsfBAalohzC9lZ0113W9cgFUVwMOyPUrqpe
2eUW79BRJrzjRuI2e8YCUTdp0NCnsnm5BjxL8GV9Y1kB/oPRiq2eh9h2FtsnxcuDL0uzxAR7dbbT
bS6DeAVNvfCPAUsAUpyKbTHyuOP3LSyhNuLGsKa+aI3AJz3s07ZbeL0gPNYlI20+NmZQfiteiSpL
DjS1BZWwEa1AOW1D81VGgl55J60+wGOILEYn31YDRxzvCQ6gQs89IsspAAEVnwL81MqfIHdVw22A
WlFPe10gwSnqBcW1q4X1SFiBXfffhCk+hoXnc0uObG5ut/nLP7K+sHI8t1XaiXxtkzvpwB6Adw0/
kBZXh68jjXchfnl/8RrjnaMTlnx3eoZhTsZHZ4GlqSDOjtxFciORD3breCv4baJ3dlVG35N1pp1d
jovw2UL/e7PzvB57pxy/CLPT7WNmKa8dpEfYIqndTDwxwaLaXiGetUUy4sURAHDBaXmd8NLRk4W4
I+DwCH7Vi6uLVkOCyMhrmF6iHwiXunYPvx6rRZ5ZHFEhzuioR6vj7q9g5JvxmKt24ul6AzlGYv/5
vW6CJ28u/U6dH/5ypC7mbPeHbyfpjxVimpYYn9AGq0aW+A/TuQn3kH8QoIYys1+y0pYrYgcuyelf
HNfnxptnQWKVr2GAErjlo8bIoBSxrROj7Fa4fEXmqjhFDyuGpx2q+d/q+hvI+K/3CNyC+Td6H8c/
4oY9KOTVaDtiBGkwaTiXHLNzzeDltRAMQJZqyv4eiyRAbc2l41UECZKhIZJBubZHLSEghaiSWilc
oogIzsAgONSWqPDj5V/zuSvsrsyxEAxlwrGBgmO9RveGcVUJQ0EGdX7TxYUO7NWFWYZcgeJkHvNe
XGEiQiTCKvn71/x8Zl+nhnuwsw+i31Zxdu/qrFFYKahTOjFA4rUqKbhiG1BZPBNTFIYVeEYLoPhQ
0FuV1aNlhaoUBM9IErIFK6FX82YypMGXd8gP6PANEbWxlfMrsvBNdWugtKt8DcF1cIjz3/oBJtHk
n6ZPr9NZLgfQ2ykoHTZCjibPip4Q6+js5/tUV9Xgjr/VjYjsDDwsnm1qvvkBf5oC0LG1vLMPruOh
KBjNCjOA9rTB38T78f4OrZ1/FUw2y0/bPL2PGekY/35jBTmHPHr/cyio71KL7TXaJ/EEWLasXhxW
oUhqH1MftTTV8cHZgmLv/gf6XuKY24ZJlV6o0J9h9LsEbA3hnLN4x9h/LVlfAtcQ4yB1SLCl89n0
JQ7iFy98THcy3OoL/e+cH+KDYY7BvCWUIEyN0GzoJR7fkwP9UIqhczO2Tgk26DrJbp3PoASsjHqY
8XSxX8T6908++vE+6MRdM4m0mfi1C+Gf+h5s40dw5wiqJobWK3BQ9NiOwO6NbO7PA7Zit/s/8w/6
x9KFBbx3JmsUSWWzCFiBDFFFQGJMsKaUsiGfsTrkpeHdM9XRYhqOJAmzP5CgORU8woJWyX+/fpq+
iB3zjp1Khz5ai1xBAd/gKWIiU8xC0cROfBPFW+tWQDnGPri6NRUxyBr8N6faGQ1GpA53/1EeZu2z
wYGdtyg932tyiFy8BeoHVGm7+JWyut7JfXe38Tx1T8J66Ickc+yu7IZEfbRRLqUP8HuoArIkXqna
yVE3Yccy7QgvJ2Yu8zEQeCpHUV0CEnY7KTQPS2AADFgOb3YGq4BDttk2mddkI1ygdbKJiQydgaZI
EefM/48+rhHyTKfet/mWKFZJNwiaIQBphfV5OFjid6JnZrKabAkUhz5jfYkCIptlZj3x6K3fJBQa
+0gWzwVkob5pIKGaOBF7U15YPCvhoNJyqY+0sC0JdQuMhFi8aiDra95IUdzXD/m1SX7P4V04GDUp
vHuIlK8v5Dl0lBzU7GHfvuL15GqxxaZId2tKCh0IbUPZpGLw6fGCQB+UVl+ijuMhmi16ztOQ1T7X
4RhyPD50eBL/mW0cY4xhxWRN+pYNt3Cyo41+XVLOrDPiedgOW0y6TSxdBYAHq1GD/xumHNKJGsAW
Z/C2N/1U19tySeC7W2zFHMqaAVzPTPJJ8zWXE1lHkc/BgBr/3/LXFvuN/Gxnu+C8pP2nNx9qXYxi
osbv9uOh8uFBW9T6iyUHKr2Drvn93ilyD7yoR1/0GMB0i8lwFRrHMSLogxdgdefR0oISWQBer1d2
4LWlY7HOnLhHYIkSdHiXBI04RRUfj9sG9Ce5eGELGgH9D6n/s498O2NXDf7Ai2whHCO1SHf8HG9m
XuPIhRDrUOYQhuCsoYdtUxON0HGMNs2oO2MU7uSvT9RQRmbEbZCVWgtbFiXTP5f45OYe6aez2L/W
0LRA8w7h/9480/VsO7FE6QYxuYM529h9KsJOeKKnu3AOrjmJlLna1fHscS0t44Rmu0LsPwoEQrze
i/zVNhWnQ770s1qMDgQAPdHugOeLNaAa2O/kLbiW8AkC3iz2I7yMMfD+LuGoeU/BIAfg2qpJzKEx
RLXOm8rbj50z9o8BkNqoZ2j/YCW/n//1OOW/oh0Vi1+65pAWNu2fO6EsK0weqiwhe2DaPZY/LuBI
DCmvOCsmhJJyBdpZn77apZ+TcGtFZWMTGgJXJC6q0QtYbx0q2oeXhATUsDKlIGmSq5AYAq6E7hNV
M9DVvXSkVNa1HSLRCHcKrkSrSS7ZtU/TaaiEbNIcEya08WlB09IZ0ZDEK/j3yPXB2wDP7w0DH+cJ
FrvBrYezi7C7X6EEaQlZ5XtOD7VkYz5C+SY5/Qn7uJLgvOhwpz2B2tMlnAVs4RP5zKMT31qkea9q
6IqOgxQlMuGcGhn1PuqjbVms60XgBEB3cKtTq3IpY2SISXFfdf263PaFDSTMzFo+t1F/bk/hMBnn
1gs7ej7m4vvmP/L9qzhmnYVZ0gI8gdNSVdElslIbQvLLR5IBjU8SBX9ukmTGB6VqJ8eOH0S9DOMf
EawJw0rQtdCDgPSYs9muEdxAXSdmoj76foLoHp10dseVzrcyJsOZ1yqCpCBjfbv+NbJi4z/QkiVx
bMOKy1XhftAR45QXGupoSlR04tM4t+DyFPUV9eui2DOb3ovV2VMfitmsDMmRi0/3UP1gTuehdYkL
vNeXGq5kCXZYFPeq86uIJJBsKfaXr/XNwbKPm388Eg6KBrm9KeW2BQwBz89GUBzL3fZY10xFh9VH
X+vX3FsbUBhX7UK+iwkiMLrMOz+T2mvuDPp9IHHUAkD2VlM1HXAeH/lHsXw7cRBF3cQkQIGwkf6v
X9HbJgguMCKhcfG3In+xxyTwEDwB1t0CV/HoAwr0GODTA+j7+NODiqGo58S2txOFSoDM6QVe2kBG
43jN2PFXSf9g60OJD4k6EMgX+B6MEghfiTF9WJtsl+1hzZKDASNrSU3Bp23nKqP7hZRPjS3p3fcx
yKBha/MQGG1fC275IR8TP80v9ez/IFU16/Ld7yLBAt1hCYq+nMXTRDlBHT73PDQ3Za9WdyRb9PK2
3f4Py2B/G9CV4CkTXbxiXfVNELYj28HVwTK9P8LFGHTaSDQjVUBZqC/MRh5uv/4U5Q12rtDuFyZe
Ev2O91Auz6ZOiyuGp+/9YDT1bG32s50/uGZ5D1Zy3YpuI36mg2bWjMmYQC4yQATojPQooVbiaOjt
AV1OC2z36nr1+K/qImJsF8Hxyzf+DR9UOUgY0VqqcxgT6wFUP1Sdw4FSf91w31Y0PJBGC+IEyFUp
Eb8JvLb8NbjsNCDI1hFsV2j6Xt6hBhe3aepeCvQsN7MH24Oj/11/K++D/BzB8PlGbrw01DYhFgjN
bT4IO/vmtti7Glc3iI+ofJ/qPRjqqiuC9BNEY74Vw47M/NDSYIFQ0OkVxdZMWm6antu92JDNS9An
Jt6hwzTVZQmT4d5gsjeqCNvsHAtMDSzIh596Q4VPWXaAGBUzlXscwGjQp4PTe7EvMCm5YaefPIwP
yOkJ4eLlT0qzcBKJ+ZdAQ1iHT64zf2sDqTd1F8mHcKWLMYsN4UETo065LoZ8hQ2SaewC+C0tFYm9
yi+dZWYNFTxfonMHTKdxUVAVbq0tzoI6rGQI5Jln6kQB2K0P8W+BCxSM+PU3IpsImTZyZtXDbgLs
z69YlTV/10689A6cTnoIzwBryH7XCXm+36jJSkWgZQQiwYdpJa9IQPDOvlCvgHbcmsB8jkZ0SIId
o9ovh94VA+mI8aiXo0Yg4ly89QwAs1l03W+QLw4H19PsAP5I8lUcnO3+LkOzZSTeFfzPqDgyK5zj
bqLkRO0r45gFm18PMjLfVLXP6ChpKCnpIyHxh2EFjflrSJDd4l9TsANAq/vRlFnAZ2KAdfJKZ8cm
Jle8xSOtaz66g5f1AIpNVBFGMug/+jn0U9ROOpnZ4EOTPj8KfIGlfD89hUC48xGHk5jFJfYp0gnO
ZesPqu9QIv74yDJnXaY/Tbs1mSttabAyjmefmsabQ2ryc8IPcVpCjRqaVz5e4WAyVhZAqf7sjlz4
621cbotMGgeMXR0u9xBa2z230tE7LoOBi9vjWtP2nmXUsgHlMHmkxvXbkXC2FSuAzvWsQSLPtl0j
lpASSOdqyNOMfKgjLKm8ASHSIXbBuAq2bY2OUyNUAhnk/APombCO0EDRrwO3dF4OwCpyMBr0h+0T
NsHekWFHK8/2V012yHpNp2AZKuPMOFHJU71jIYFnINsFJzAAf8zXQ6qiBmzGejy+mdbfLoMA0RfL
snIH0uJd3u8smdKnKSYbzuTIOfMJNFLGr8xk/aO2zhtf0et9rKniVOU+UjFVrtkGpayGh0Y2Z/RM
HWQMuH7sRwMD8rtrWYTGLovOjEw9+FemeA6zCD4Vil5IdxGVouyoxwfX2lR/f9K/wl69Xv9DoHIm
GuALofwo4NzVUzmWpu3C9vPhusCJSMal8pOLabZPvhoJpyL5QhWcGLNYfixeeUnK3MvSb3oGketB
cO6WVHbKI4GWt7+H8EzkFhS0NLnxPZD751kHlXPI/ML8dLxRFLhknIggPSfPfyjTy81/AQYCQufR
4zVc/F+zfYBVoz1I1XtiethJCWqJMi2SawBfSYMkyA+KRte8cUwkaiN/vuhicenvV1/Yi725pPnC
j1fm17SdvRUz1vqqfDHzXoKYOQg7yzALZxhSPPHU2tu7billWHgxMWnKJZIU0PMowSmNglc8i6o5
2C6k3hqieGfzPdKoOIr2EbxLQV8UuJ1t5sHERiOLV6rd0APKxPnQOc/6nBXz2kxEmfnHKASsJHbT
f4gqEKHXgE8ahCd7DquHheqKU4KedPeVXRr9lxlsfeHO7vK12m8T67Tq7qJKDWWAY7gSPrUbmaUZ
L5qIJWh7ILg3kkLCBIr+iggRxlxyFTXYVuCROgF4mGvhYHl5ezgKvMEkfAkmH7Sjs6m5DAERytQn
STbDA03san0RCGDkJyb4H+E2u4420O+ER/Ti3lDMOOVj4aDK0eG0ONms4PkzJ/qQaCpKozMKgFKU
sZsAX30VA8pE+7ZYplVIPtL7W/nd76XHOIbPfzy6RwqpT8qrQL09HDWK8WFTEdJchwmXvYVYq9Mc
U7F9obGyAeArEHiAIETeZ7Anp3mCehHbIXwdI1vjaQ/rfVWRg7kMauStPi3sjVWb/I4Xft7lFK6C
sIU6+q0TzIo6iScVpZtUMg2majJ/QD8KloVJe1wVzUirGmOSFhVjRQhxdQfOPJ/qzPBl+9JFgwo4
7zTQUvvKSK9ddP8yAuaMvFr6oJskmMvQfOqFjEttp+qrmGL80WNZK788aei8o0jMzfurZ9li4zsy
8+TNNa/m1Eckvxr+e/GRSkevDRZc3kkjPMVUvQaclWhpvD9/7PhfevUhyPXK3tKkTUYpI8aZI1Hj
gOZSknDAnzT0+sOzxUcCvFsQJp4W3fM1/vZmbXg/BQTgjfpZNnvdmG8jOj7EpSBhcQHj8yR6LSPG
+RCy1URsJNPxdood6Czk0HLEmSBzZfSb0NJWtK+41UtY6h0xSlgZ7AYb+mmQI7Icr+hK9WAoO7yC
HQ/uEij7kPlBP+VALOet3aVG81PwBa5A7XQv13Z13cSIBKQlkjlt092u55TNzD5nYhX3oPRE/no4
/Vb34/GSxKjeIcXMlnRrHFCoy2zQanlS/1YeVCa2fRcDgoEQOuWpFG5mRghZgEgtahGWr3Pi8Okb
oR3A8abi/p0xCwaAG5QYHHSMj9aZrnNXBUGTVWqYKmyMoYMsy/Q7K3PVPnIWnA/cHWcA+32xMkEp
7TBKH/rCIe+s+sFaIsAQa6xXbUuIyAKhZGWp4nPy0ljHCn2V54WKeVz+HJLSU8G1cAOxhlgjGBmh
B4iWj5rNXSpAy/89r+jFtprR0G1gvYwLKm5z/AA4YPs4EZQWxl1y2outIwK3ZrdMk/vmo0FO7tj7
DcjXCTCmCHhNJ2jyse2PdGcL5sKj4CKiVtSajU5gK+9DPMM5ghPYANF5b9CsJ6kv8JJeRmdkZ4HB
ppZkw/rI2qx4G8m2DRwsiy7EHUnnUhDiE0YM/NVpt0YJPm3K1QPx4sAHXY5czr4fUdCkhxXbaMkG
msN8juQdNJFjMhHgzzo94XP1K20BiF5Q0Ajr9AAG3nM/EodgLFSi2fZR9mchFkdyBvyK1XGjtJWm
x9o/wTYZXUfm/hgaM2Gq1md3UDM1ZmvLRuwIaJuN1GnPmiLSXJd7khtOeozFcVJErQ9OhhmhVrmu
yaSPXQ5iNn6TejS9AL4Z2DW/x43LqcsNZdlnyc4FhZPx/2vNNOoghVF3U+I09MsImlNpEP27NNRd
/S5VdVs5exC8eLf2Yr3xbLI2FB0R7tpK/6ewbalJanjTXj4ORqTkuJgGva7hi0TDMawG+QWOrpmO
aG5WOXqKanLM8G39XtMT9zFQFqIVUwE2LGbwaZvdDpAPipF9Rp9gVp0XXrcVPX1suT/w3D/jX4RB
y/0KAkbCLy/mZNiPidXHtzGKgHgfT7/9M0D1kkJB8vrqoAI/R0lK93e9mOLBMfmzd/DPKYQbYMmS
ZwtDsb+OxBQ1c68b1UVT/Lb4OZylXoA2FXWW8TcdY/jbA1WK8Wd90lw8bTtWL9ED4gsppjCLmy5c
92KUt9038gqPGF2qDpIp6zXBBBOmRKeAihOm77qK9UmEB7sg6uKBtxqF/JWOBiRuJn1ZuAZIFg9c
7J5hY4kWbtF1KQrsuWNPJUakSdsfTgSkGwQoIxRZGpo7nQAnhpth8SdriQXbvoL3ClpNhcsbi1LI
7jk3LRYwIWLdRkUjy3J1VaKFx+vI1jh46F0NXhiJsKuvVHkQs7oqTmDTGSp6Ujo32Vfy7bG3RXA1
nM6X0ZiTiIUxiAI0jzQB90Ch8iwj6D3OPMu+s09OzmZ1YI7d7IHFZ2+c0e0az6iUSONOfcjXkBae
cYz43Xv8O0h1/OdDn8AggXM7N8VvjtVA+knxB/qv3ayIltZySKuQXkNukv0lxROicQLg2wULJln1
/1aQak0qOB+TpPxkWgSx9ikjvjieYc5nLU9Q8C2rOljr3Qr4o0e7iLDI7nkeVOH8sV8sXyBhG1Io
Gc0GdLwMSiyoXaSjT6kVFPN8EMdOqmubaPZbi5eYcN5XyGcJSHqNL2Rb+TlMZ+qG2oa/SigzDFh/
90zBUKjakpyjM32t/jN2XQMTrf11JuhNv6LJZRSaeCuwmlZOHt1CbG+O3vO7Zf0qZl+oJoYHeTkh
Ai+eWfjRoIK37oCSI6L8rxTDtPmMLY7MtQ/uUrJm4fipcfoyKtbUF6xvazPUGCzpfw8aVaxpLscn
HNrS8ylH6saAzyZyLTztZ6cKiCOgzBmc3ObEDzcckgPj/WhF64HT/CZRKfIXHQf0M93hwp/KEzvJ
0UHxtXqfXx2rjzXkVxKYXnk/X+rU8HfkYFp7BKytD3SiD/74SNcSQpym3EHGmlSDWeN0tih88MVG
gKj4dEJMO6ku9Qv26iDL3FdIMxrwRWxijzaRCwxkkih+Uy3X0q16wZafrP0eseflcp8ZduIAgqVW
bxev8Dh32IYPUNOW0tyM4FMKxV/R43Tx15Ni3MvJ59YsLTOuB00HfX5Uy95mc+mQISv/KvB60EdE
LNcjM0CBTD7ceSI/MWO2MZncOCP06HXQ6/zl3vSJpeX3aGlmNWzXb4CZrW8h01rBhn5AZPSPHY2U
etvEovTcQ095Ujm2d4/tgPixODseEA410LYO521c0OGU1S6Bq878KGtGIx1rtkSS+qarpw8wXe5K
BIoCUJB19eeclHIUn9EQ2Of5xfztYQRhHAntXXj8V2KzTldEBrRgeXP/cN/oGpp5q36VMQmKml+3
DxY96DKOKpOxrKqdpnnSfRJgkR6q/SO/OuM25pYht9K22/pnfQCRjRpWsrmDbY6/AP0Y2vzjOICR
M6hj3RAjLOaOi55UxjBVGNLHPUlHOXR8FcZ6Ab3VV5sRv3DvPk7lg5+lCQyP1yvWZRA+HWKhom29
0vn3evSgtkOwqE5gixDsUTcP3DyxZLcI59wDnznp8TS5/GexugZuZPU4DBKdo4hDCDLUy5Of1V1x
htnJY5qyQDZJzt9NpQwKb+4dpSfMAK0WoKrc6ChkkhPVlceJXXK+f4iUV6Vxza9tmoyojIx87BPc
b5T5aBbeeOZwIx7EszFjsE74/tTgvIHv2iOIJMKpFyKxAkhq0pY93ibB6Y8ITQrDt2IaJraLZyAV
lhIsqi5i53uSwxc31C5u89Y0q092PC1bG9KV+21Yp7YoCcZoWTx+W6yrkeRyaat4/tljsJ1MOEL/
eUtmC/+C3dp2gLk3IQMWFyhvW45zyRShoVwpIKFA0VQ2/TgPEqIV9RQiuhYcIx+MApddI1N17aSy
oku4rSs3zV6+AN/yjlyjA2OA5V1v/VwlhyvrkuTBaD8/GVBau3f1moV4dcEKMKu3baWgo3pGzunw
9uHp8yBYu6knvEfX+53dmmxqUP5O2OwJH1RNZu5wBtxFPgR/zrJpesUkHgX6ljEbGO1J4yUXr0x8
vN6gROsoAdh7VQ5vTJbL6YAWOWKAJ9oZEV41FGYLW2km/OalbskewoGP9JPOsisycXlkAZZQIbGZ
+lbM65fMcjwjb7BwhWJWTM1au0yw2S50CkQhiYzvo1sMbYxAnhSf+nUycM8ny46uX/gkCNPpoNEh
7ojLev72Ps7nulNRybo9GTuflu/DtYUlMZtF4RtmvWshEE5BcSaCvHFmTq1ZZBGt7VBQdNafEYCK
PqQZWRRU2alIA2Ss1v9ja796Es+nwfZQVqmr8T+e5dGlLAioCnCFMTnpyn1HDrExZtbh6+k1IOoX
jTTTn6QO/Lsd4GiUvVSiZ8Enb6rgAM//EKS0uqStFjbeVKKY5DFFhlZN7pfo8J7yBA4L1lFj2o2y
09miUUpHO+q6R2fZlDeH9dISHGWl+dFjp0eGCDxVWSnK9dMIFAH5d+NFz+ceQH67HGGlH7GNd/0q
0CVHw6AnFhUzRyoZ1vAJXHGXTGDFqsY9sDKqkdcMuo8i9uTpLPCGasVaLEHhzy/YA5vsJ4xWHlf/
YG7PtUlOQyJGi12LqlXKqrJvFsaqSBDD4dfUEd0PNRNCTHMftlku57fdEVkWITdyOefCIzgqGBzT
CIKncApUKw4WVirhnRfA0BmFfMPpwsR+hFro1aHITYcqWFRMMQZddNd9bkUwtGsoA0PyoL/ph+x8
JGmg26+bznPlnHY6zt87Hxh75Yaumac7/BkA7WA7S4ir944OaLriNKkenqe3XUyQzhaf9bKkC2R2
ks0BwOQBtYKUZNC2f4f0zT+9o2/PQyDF3Raai05bQzRtDt3Vt+qo0qwivN2oy1GK6QYJPNQXihr1
fV6s/dpuims3hULKe6R6SOMJKov6jvFNYSoLoGtKPigPyQu4FqCR/nB2YVKxB7D2YWgsR4+xBVwu
La1ujOt6d5+/P7VgHVCZ+ivTqieUmMNosRcQW/+ELHyr1fqGXABjIat6vF/R7KZtAN8psx6lvP7S
cuvBy6j16HLdHcq840Imzft532u1zzm1qdXzlim808B2rSb7dOLGAzRZqHJvZfOMzGHMhjHCjwBU
KzGcoQZMoP+MTawyfhNnIM7AqskmCesmvmuIEvYLlFpzITG7ECSsD3o/kaLCxkG3fXzsfcJRma6H
5wAYYzWmTAMCln3w+IZIBmrspFm1Dn1rFbznmt1UjG1j/ZsC3dO4dGBIfBqYJS9aPlQ5pEuqu9Lm
7VIAWzAKULSjWYRcsK9g/b5iQg2ult1fjHACZYATL6+2EcN+jzk5b5DEH4B/dqM8pzczi9i+PTxS
T2OizWxzrQlLutWj791XqLbKsv9cAlxeyQSFWL0leymIckKdmygmEiocoFbjl/K/dGr/mfitrZhz
n5hkDfZmE4iBpa1zcZKWFEsE5/6kE+JMX9PJ4aryV9GxHzfaSSW30eyewPHxn12ivDaFmkVJ6ICD
Bb+/VT3wTADR+1O3JyMfcA3l11e2uuyikxVyyLQPa+ARcRs4rn+mHZRkLyVsmb+FMiCR0dqm6GMX
5T39SqGR8qVDpyb1I5Jv5GyVef4AXFIgWPBLx8L2N+GzJwejMLyR7HIAQgfvHRfM6Ly/eSE8ko1m
D99HIzOQHisFYQLPzjyvRCvLo7C4X+VdYTnuvtaDVArat5ATavvs4Y290B19HyF9fQZ52hP9cJi7
b1COCkQq/kWfKKdhYaLm5kI55AypU+COofAT4ru8uwkIBKmTODpvDS+cGnY9TvZRu5WiZSf4UDBi
rpz5/dOyBOBh1is38maJyR8C8wAUIiMDolc68OUonjfcMDO+4TOV+Rq5gB6/KfUWzkzF17WmArRb
W1qKYa25JVrkoc9tu7HdU7LOwwxqICORK7ZSXSdutaTGHy2v1Wt4FmL9Ts3uAMTv4Yr4uwEZMb6J
YE2IraScnE84hqnnlsXJKtSxpPxrL0ylwt4wJ8DTPUovZRW0tuuo650SzhbCrZ6nby3s2+6MCr4F
SdaALxbBMrrlNKlwEWVwDNPKxe06SGyajM4Q187XeldFiQd++QwcSd1RuXGBXzHwthlaGQ5yN2mi
oiCjynzzKF7ehGVIBOzSSzIi2dVafMgT+YpzK81N7m9OPF4Pl82Iam6iD5PHbtg9ySc/rQgrdWr9
vN4ZZG2qchDJmSHHadgOJN5hDvtYXbMMbSnAJyq3197tUiHED3H//8L5YQvh0tawyfm6PPppfn4x
XOMYzxs3wkDoaaN9gvP3RE0p2UTEMbuB+j8MFXIFqQC4jnCGYsLY5wVw2bk1xKEMs71RdFefaGsb
RrlQVVIEUiLzWDyDdP/VgfR5drA8TOFDZPKcQKa9O4ZYR4UrtEXnm7Zz4KQSgFQ+NG9RNxiFCOc4
d/YHX4OlrqeuQ4nloWS4g7vIwnjrEJnwC2JOlAXwVZDGtq3wztnxMySXMERurpfz1OkJ7f5sEOT6
GvdfXaHOBE4mrc9ci/nRkitVc61WuJaDSeKHeCuYdlnLeN3OByCuwgNRWcmZkhyXxXvSq3KftJiz
t4OGJVBozpPD2w6iWRGm8iYXDpDVPAcKKhftxNHtc/WHrJ97L6/bF07jfNj1X2xZVOSlhXftYfll
4JK9f+O3mkJii0hPW6s8iAJf3WyPO1mU0BAasztSGbKHfVnyHyXLomEOBvz1hwlLJY9ve7WsbXUZ
JMtC7EQy0aC2vHBgE40iNo+BDcQF/Sly87NbRKHGcp7XR/FepGPPkT872jqloLmIxRINlTU6GBnq
dCv8y49Y/xvGkv5JccVpxw3Mxm33x94vDIN4f60TS8YQ80BrnG0SBEHCSBcIoA172g6jYDe68n+k
kxjhZnvvSXIy8SrH26Jb3vq6hKVXcwB22ms89EzA2rSez9wtzDZWur6dxfLdL2l0Ux2zldu373pb
3emPm12M8m/O75qbZ7SCVjqsxNdMgZ/yO9cJKQtKeN2EXlNYHBICVfGpIjDIJnVHmRj6FzElaqAk
T0c3vEfrSTT4ngu2ZzS8zQ1ta4rvOogwx36QBv/OFfj67f3XKeKBqZNT+QrP1mU0mK+wLqCZMCDi
pGsPErWiuBc4Ti94oqMbtV5kuzv9mafODNZHx/XMvSv9/mnUPNW2ukhNCRrwLonHBoLbQSYuk1YM
BqT+XEv3M2C3FifY1TPnMyY2NbBCSmNi0UpckFVLPdBjY9eaeS3fp/4QRazvXzcGLnWBEqZwYhgz
RrGO9JfwfShe1klrcQpc1bQbUa6KkxsH49uJfjv024WpB9WtRdXx7e2TNWITcY1tGESEjmbA6RJp
smHNItds+kAQhwLZeYE+zh9D95E02qVsoiZVKefHntBnv+dmv5Vjmrz3nOwLGDoZVsAaUrK+VKXk
qfgt4HutAx0y5esagoPJOopFFGG6q0FsbtemJ0+K7WPXy+wuzFErX7ax24V0c7x4QyVgmZUq1ltB
RUGj/L+bloXrhRJoWFLLJ8qlrNS8sJZQdNxzSR3RSwE5pCyYzNYvohK0vsbyKvaspllt69m2MmH2
qw1szjW9RRDyyh2iYZGZm3Xxb3WfQrvuFg/HI1OofGZx8Vm18ejlKzoRrva+w9xX/4bW4BTMfCK2
kQyBVnFwPoRxFbBlH3a/GT1AzVTs7apy+Lip7EfVK5635Y6sf5AUzliqpRg0RT1k8CVaY9vno+vr
LrvmgbuZpR7eQAShxnBX29uXNEZXhCUrMDb4DBXixbZZdYb7N8VVqxnWYVDCTqAkBjfv03wpZ7Xb
Rs/lbaW+hsksqUvpxkV9K3/9RezTg3kXPN9GFYaajoruIgOpiVhw8C+Cbz+DuPMtNrS1eXmP782D
d7Bs2o5D6Vf3mFsjP2X/Q1ciKiA4S43Lg7t/1o+6rlkwgtbmar6khtnPGi+U2M7/YK4iwFIwmcXU
GloLjFrSwf44p9+BzjHDoRl/4beex0CD8SlLQrdgMN10GGx4qVhpPCl8Hav3qaKsIAVoXeaF/F2M
joQ+nL+Ebke6A0SWdzSPC+Vv3rNWKAs66n94rf1/Dn1ysUpzbNJ/QhOV4KIwIjEsccBwBDpM7+nH
Yzh/J1e9UsWCjpHyzrjh7ZT0H/H/ikCTDswX8vesRiHTQGKFLS2wRB6pZfS6EDbefru7/Q7I2X+N
JYZ4Uk4yTxscjxPtyCU9j7EQukKaVfkBkyXeE7R9DfdmmDstuaPLDojJKAu+fH4fH2cF31TxUhRW
+pREBEza2gsLozrzU4kAcVDD6brkY2V3130MYzOt/H/iFe++7cm+T5JeBzjnEq6BbOzL7EB5aSmg
aoetZhpz2mkydqrMY3sRp2Wgn5njBxZFgANccUNbdmbGbSnPOLNc+mlsaNSHnR/u84Jxt+3MmDog
zLc341bXF7UszMCKGbQ9ph7mE+QCUFLXcVErnwAurGes5YIIQvX3TgDnkSDtQA3mlKNqGi9xxNHE
3TKeozd1wJIScFDKNbt2s6YpLMJQgqh9u/3U1s8ZXM5ya/W50Tgn49wl37nPh3tzaabS8H3l2yep
520SydO0PRhAEhivHyWeZCr3ZKpj82vkS/fAaRbKrO1skJO+qsGdvu2NikPqGXqLk2l/P3xtoBG+
TzaEfdRDyHXHZZ2xgFJ3Gr5aUqTkqiQWmLgEu+bHoUSEsfK3wpP7ez0rnGQtvaOEA7isYWwahNAY
sZlGm6gFQem8uHusKqSjQJiBDjT9VLBSU8iUv71n7bBTaax4aw+DOG181WVpEPy/AYoDDBB+j5tt
DNEf+hEBGB9DyurOE76AH9K9Rl/QqSrXSZQzwQJdEiATnyjRbY8mNFPoEkNNeOovHJHUz141Hv48
AeqAEokr08y4NkW25p/LEu2FTkncOSJw6Q15A/cUvcoa5QiHTgxou71cLS6YmSgfKkJ4ddj2J+ps
vkeHqDN2ybO7XzJmYaYVeQleoJSta+ss12ZTO42ow18BAlhNfZddA4R2pcJyhp22T1j4rYjGa5DC
5g8eDcciQWdGSZCArrnExBViHJ/zMoveDRTmkWgG3TrXKz2MkGzEfiIqSH8TeRCWVxykfZViA1F0
VWkryPQYOd5genxQTFeTHeg+m63V9GHhJouelWxLFkOlwbSrdGYiJldEqz75mGT1HXbdErSHK3wZ
C78s4uVZZvbCfsvAkkeqChPvSwMW6Sh03FKp9GQkSNET7koMliaorKrbo8u0giz9RzS765RAcJx0
O3u1QTozwp11KiRYLge8v9oyVuCjXjFKNdyXGllAMqtObrpaNiPa8GS37SO+zHvdtmIbEA538vcD
s9KUtSSpm8iQhdcl+LWjH8ujKtK5uWZuNGA/pKfCQBPm72yUoVNHou7xxuZs1SHz1vgGp9fiti9U
zTCIM/hiuzT4w1rZp83fV9kWHKou+eWGxUnKYI3RfuqE47LS03Bhymt1y8mHBPNH6L3QR056MMRw
HDhAdmd6N4xhOccv3QgWI3+KY0GBwDbgh3Tv2Xj99+2nleGIcYqsspLFlyXTq2wWmTkOC3Rrv9mx
DC7+P35ALCoOo+Y7XTVviqvBQN2210rvIrOpJ52xnuTpOOESCJ4qrhhBGFF6T6IxiPTZskbxxLCV
s9AZ6RRB/BEGynGJRmfuhnXI+UkZoqEU54G+vDnTtgt74AxG6CMou6JXG0Pj/ai+SzF8IpqObT8b
L7eA20hjSILEaG3JP2gL61ONgx7Myy/b/RJXcBeWFdo+WTnBTBHxteWDxfy4MWJm5vIRrJQwLKq+
5nScaHHvjT1AcZ4dCxC4HivIk+IETTmqU/95SNnyjJZFWBtcNpLpSCukf/jyc9g1FN0tFGICAFLI
Ub1Hwgg+b39bnkv2K6Nez4VtEGQ4Xy0GgvkcBbgDyjOFEyiodGo7EvHqiVzk9dBMpVAEwGwj+g5H
Wq2OpMagErNVpXOc9iTIDcLXsL/Qaz+GctAYJZPm84KgjRVDHdqvmBSwY1WJ6gfqZY1lNleiDhVY
jV4mZijAA5UKT3m0tEMqfhTnQ0t9O8PPz4fOSf19TNdseqoLOIRtSevGOD0lW7Ilxz91r+VC1Vsn
TBa6vvlqZyDvYfcAhGjT+NJLWPAyKMrXs/wGC7ywO19sFWLMC757fLtvDaVOUkDfvfKnu77Hr9yh
+4fK4q+hBuubI9bJNqeHfdooHXT8lIbNNWWYDvZ1mNoxtEjnUY7CxMaQ43ZB/ZD06OCiPvmil2a2
LgLI+dEeQfX8cPISJIGvISEOskUjWNL7rSkaoD27UKGac36nIZcmir2Nz0ZEkEBMMZ181xjGq/Ro
DOEVN7FGSsuZwW2JTO8h9QNsXqxyRQCQnnznT2/4TNS0qyLd345Cz9zGqY8fWxTYICzFrMLqQu7p
X1znfnDqWPu4AOOutnLO9JBUo/5W2L1SVV3tVPy2Kq8Zlvb0HetezJNRMc1u9YV0xB6l23GTCPlc
bAjLQ5Aapuq6GMuK47RkSHu21am3nuCc9S/P/dmrXlpXUHaYiZw+KaXltt4K/CTd/hrzFCtjeCAP
SMJ+YIPmuwt0NxIiS/V8zVTU1pQNegPnPFFIAJfP1nI91rE2lZOpCJuB+bqGHV5dV9nej4XprbOo
A7adT+6raCIsYDTswi4AYCsCF48BigWA/v3SWoT/o3JbSZOzi1ce/UATKP47dfjert0HAiCrPbMa
yqLdrEIlY+9InOomtYImb4tzQ7qU+4Ugjkz2Di1OAtcpITRE/NqX0nMLnwpbp8Fn5xcjfa4AOQia
vQ7BkTuIKted0uFDkqYqOBpWLEXuQFShLx8oSf3c8GVukEHlJp7DSFFUqAzQLzapPXZLI7ml6khn
8zqWImBVlild9CHv79oMfhXMiCTc5M3mbWGqJVZ2rmy09EDmCVTVljxgJaYJlaHOVs1hma0TZxQS
DrizL8tWn7Yu7vIwKUixSwen7Foa7dRycJxMqj6pqFDN/Jx3b1tqn9aJp80ePIugZN3BeMGRUtel
Z9q23kGplc3Ey6M/jCuE2eK99C/NoyHb7vFeSSgFfS1YmtOpZhnOB/rMqZt5a3iSBM1CPX/qfKnA
nIjchjZAHX0WdovQuYsOoR7Mx7vn4LqS2FLWM5s3lqsqxGAfOCzhTGfyPsYU9TJQRy+2Qq7UcNp1
W0kgk6fmIoOXtlVqDNEr0s5mR7mQvr3h1zq3GrMbwAICIlZrH5zjhAk/TswUk01rCscRakBWAD5u
5fgHkVWheSElNg+gBjTZT8+Fp/ZrhoCBWr6k/IqDtn7P8AAQ6VYsfWvMQ9A+xL4j5kAdtCBPjnwJ
JAMT6fcbq6TfI116QoPcS4laQ/a/fo4oFzM6/EX9bwaWHIJMeaze7pdu96o16JnRfPzuyb4AjZAd
xAinD3VBDD8Bo3sys3NA0ocn/wHfPq90HOgd3neVXWan+haCU21r4n1ykwjojRpUT6A+dDq3fC3o
KbpBbFTPAJ/Wn6c+LOUaooKtM9hOX2i/8KIW0GJf+WOBoCYs8nLttLqRwqSkJKOAjgKtqu97FYbB
jA5ewYsdAIb+u7cI1htdnMYK9SQig/Fuad+QFNZMdDCIV4HkmTqnoFgmUC5YOLLMFMtec8s44r9N
yMgOKFH7ue9vlvgLOVH9u2XCjlmJXWye0h+gKJTMm7RWVlHRoCmnSAJlxKqY5Q3wJuYnS6worC6C
kUetchG2bql5Ac+N6FggtAVxXt55eVeFUGv+zcYPox4VG+ppXEKpX7RZzD0L6I74V1hrLKmd+sED
tUFQUSeSoUWumDsIVt4wbODlpqxg0+TZQuscrk6Rbxh7h5ZHCBZ78jsMpoAkVjxpWrA+qnzkUZRz
VPaXIVO3rSeVugOsPsqHkZ5tigR085JJ9GFDBaTbrzGE7hQRPg7NfoLODALc/gAwJv27J/FpzM7L
gQJ6Fg2P4wX3tINGu1BR577+QDu1DK1zSw0wxyERr4Hp1mAlvWntlr0+sWdKyyw0b6p/n0avPvYy
N+suWhyHW2D5x1djgplVhdom3KEGU1cbXKHZC98KdQ5gX3PMZeDbpgfTlS+ZwiludLTqTFAsC3Vn
IZXyLHfT777LetBfyF0kphaMsX9X0/WBw0Cbx3CGQU7iV4L8UXH7MU8i5wm4FDz7uwrOYwwPmWH/
TFK77mfTo9f9PeSA2zcC/pYf1XO/tIzcGKnFwNkDgJ4B5kjwMbzXhtqajTYKY/luDY9ZJjBNs1OF
16kjaB2YR/wFiUIWAqVg6PWSGFKn97xSg5xWKLYRtoK724v39EiuvTzVJOcB4FFdM0O041FZNZCN
Q8C5DXOJxlAE19q5tJMXczjfXNVgO0fwKn56C+h8SS/nL/vlWbYdLhvGWwbVJk+aJ6ICENsPBr5K
WjMXNrijDXHjOscL5Ge3R6XCTl7FB5+ta+jyxqaYe1P5bx+fxVmCaAGxZEyNAMxGj6HRSlXDYMsD
wiATieKf6ijM9GussQqyo5hjWsKT+iun8dicsq3jHqb08AgNnUMKDWrXg0AdpML/OiLW1/4oA3rm
DEr7V0UDCeOsV37fwz/O4bP3nS0FA+bgNIkgxTJxjg8xt5/MhZ8jgLqGWeUkVtVZ55w1sLu8nhoL
6aNosIRd+n02h5GNBwLR1A8e6VM+oZ25EYYU5fv9rz6hsYXMcHqIg+oGlIsMxZvo2rNTj3TwyCGc
fxgXNiJ/Dp5/2kMhpfqZ4JrIc0fCA/TunHgZRyQDlVOKZ9tl8QQ1Jz9uVuCR9/vVkyslUc2x94P9
Q1oOL8LWdjYpOrLGXykV8pTVybRq2Zn+TomXHikXWdIABeQLMUWkAQsmsTzPcjeZOnXdhh3ZwhBR
QMEX3X88eDGdfhf+kMCWvgBb35yAa8Rh3uD9zefbbYgeeIK3osD1qmsavOOfPnweIRlNi6ij5pp7
EM+VLT9kQRAkpJyRB6Mepnhdr0ksY05gRA10QLa40R+UOZOfJJ4oDHpEsBLbmU6GN+tVcRnB2c13
944kYXMGGbGXQQFI5o2pfDZtIoI6K2lj8fAhwcDXYL6nwZKpC1jtXKgYxzYsyjJXddapcXizjAQf
GMtV09jAWXhkz+mfPpubdf3rJqWkF3uIXhHgKHHm5UTMutRA3fjIQpt/afS5jVGap8u7tmH+OYn3
CquIlefX3IEyd5dL7ilF7EfAyyBgUFHBnw9MpilrQBdIHVkgs4Ugxs1LG4juWtVyyzChV0De4L/H
dXPNegVYrgB5OKroRvCYI7fEiYmyjVqUuhq3mZ6ghoiic+Z3rwO9RO7DszO+G/mIsPqdxpQ/GYPF
LOXo4CUvRdfKdsUDPbHrWRLUX8Fn0GQQHrcPyQqHqmCNdxRmnRDuON6srjaA2cMoEheywi7Kavs/
+UaXhMFz1ItYW8FvL522Kh+ZRMH5SU7CL7SnVRcZ/VJQpdcqVk45XbZIKHn+9u4sVhrm4cxOECDn
W9ALdOL5m0OQvpg4cyZjZyvoomI0iYPYh5sQxk3qG60pFXvUxZ8Fgzx8ARzpFCL0Gu0Nx/3CY1bJ
fGSe0USCTLREx3bbsUk3MkzAl20prmXGtFntR95DxpqNoG+ZgBTsrN4UJDH9lYRWGYJ6Ugh2TewE
qPNaU6bK5z/okpznCa9gQodbs5sWRXZ2DMTgqUoGHCaE9vZGa6vButRy1Ne/j+mP+act3Dgb/42Q
xD1XHfVnPx2IZSOmLpWlyQSsEh0hzAQgTg7pNlig9lSOTNMl8YFkFDCBlrXLSLIp/3xj2BkXEciv
YMMFtaec8jauCLIf3NzF6Rx25Z4parNUwmfv42LSBrSy+VHUSh0GWXfCOUyU2AkvC9JLpIbC3e5l
LKmoFsCKY6K4hWm0aDo5lsxoxn4CopMQMb4J/qyjRPj2ZnEXkI68uCkeSuiF6xh1ZxisS0po0ovT
zN1fACovq6VAMBwovcRRamAvbgkQ+rDjujVFpE/dY8OGU9vyKJ1JGjhWR5/lLrqJSO8a49Evh6z8
Uf9FFpIcWm3q3qYG1v5Tk1wlO9UiUJ1yfDPeg6binEOdV8uR4mkOdw6ORRVrmle8JbP78gfC711/
5h1LH0L/SvZh6qRDnFuIS9+J243dSExCykZAndPdqaNSI0jWtrho9Lxt3EnsDlX519dIr+rB84/A
/k7HvZOhmibzTCvG7qCXwfwxGBbpz/x7icz3azdSe1RfCWnaJr6RRfrPkwvADBGcqI1FvopSIxUw
w60brLOw3y91LDiuQgdKoAQbUN0smoWX3cY2G86kXGtCA/1I8bK1xxnsv2xo/Ui889VH7ePCe/7N
3X/GJNCXDuQwhIj5edw2LYTSpjkSS1XpSvQq6H1QgwgOrjzeVcTmSZ5hhuK0crtqbC/lYl5/8wo1
v5uZDBWgyURhudZjwLcvhmFuNVgHoyIZ7uDeO/7NGkcT/4IppNKIrFNBxaIJIw75kep1X4Hnr+A+
eagsh4tgVHwNPNkeZUTazRBIZ7P8I8ESY/LNcITqYaaRWzO4fkTT3RUxanmhZrCqN+nBBdGfY1iz
bldRLRV4uz6cliU0TdM5kbny1NxLsq1447UuRptHz1jkPxBjPnOME+27Pt7nj4cGHu7R+/DxiO7G
V6I42l/55GxEJDrrZDXm8bjlasPMtnTGSix2Lfmskn4pokN+7lTxhUEm4R/GvATgOvXryHeLtqED
+Z3A1oAVB5uAiRtlfsd7d6tTMUAlW2Ewi3TDr3FBW3cDSP9vi2bWD9RGXSfHEZ6q3OD4XLdK2eGf
mC4psrUebL+pgSQbLeizLYIe0DiWnZvaEXfvDHm8izy78Ziq40Ufkhc3azvtlL3h7goJ9FVkyGSr
6xPnEwHCouwk5j4jbTojxIS1n5huOOl7ZzfGkG6H3OE8Zd5Rsta/dO6jOgKnINaURpE//DW4FoY0
L7bt0xGqea1a2Vw0z/um557cdH9j7700YBFG+WGqPFy4ev0XMyIRtGiTHNUfvnEtKC8nUJDZ6ZKG
u7BK71B6333wpt0Rd4EWcFibgLhbupq+npdet6r7i+sQLle9UDcGn71wiHXzLgZq+YD1hbc9jDXJ
PouuVrqlqG44JIpbLFE3N/TzcUSYbY70U3DtAoiUuRHn8z5RFGV59gh7W862EI/EWNP8nTbcHVIU
+iNL0twkwcASTFT6q9PR111Yd14DtYZcsH7gQdZkTiVShKXbG/LRVT0OT6hN0FXgO8NpULq8n3pN
/aS7/CRrBYHFUoP1r2VNNRujbZTwFzTyGGrUT+4DFxBkT2h+2KC9DfI7L3JeoMycVe73eyzP/I2a
XekeFa88irc+3u1E383/4x6uCXTcn1WQ5qvD60e12Bq57BYBcLG4Xx7zRdFRuSPIK/ad2vxR4ZTx
+0cMHL13Y84ZfwNMq55KcffDRljwy0H+SVqrPR3H5ch/iHXR6JV09QXeIIiGElyN7PDB/Hp3taHQ
F+NNxFRlo0EcJf0L988DVLID4aIN8vM+8rLOg4SrkGOadJdJP48l81Z1xkLt7LO6UmODmH1exeP+
j09X1B/HBebYWemPMIZaS0trkn1i8yGyJjMRugrt8BRfvlzcZno3JqF29QRpynVd8COkjp2pXWS9
mwkrSl1ikLcPZrRjKVNg/cId34/fmIb7vwuON0yvJC8pr+u2r17EJqMoLOEtCpuZEjxvH9p3OA7i
ugH2OmxyfeXT/uebnsiVq93DaDNqB/brz8iAsDHvyK463mrjCL3+6/WXbZfLCin5USBYMj2uGPXz
5/I+etiDhzZ7v11mQVSJzpaQmdIV4gCmyvbAI07Hs1RLc2LqowfH0trtPfGSTTs9gdM4fDuGNA8D
6AmGtD4kqcg7vEPWXcoGmPRGCDE7MD631HCO2zRI1pxeVkmzKvqiE9HTlSlHzdk7ZH5flR18TqH0
yfXRCxJ5tvKc2QecOOihMzKbuDvksfkIIV5sj67UmT4lSEVhYBf1NkueWIGdIHqZ3w1+uxivgWWC
HeacishR6Z5CtogxHjUYqjtxJjmUO7WeQk/Qo9ngCTMexODyxW91DlwyZsdkqqrpfZbapTkfysaL
Sgyw0EuHBcqN9OZSh/nArdBhvGzExzsyiHi7Hhmp4dFiQ/S/J1BeqcCjHJm7mUwXCFVeyaz8+WRz
NmKPZmW74fkkp3HMKXxMyF6xXSRzrxmGQ2I3eDR3+MIGEZHaF1ZugWz9v2lcek7BqRHMgRcDJ6/p
iE6LvOLTFFr+Jd34R77KUD/3AvD3ek7b0kvCGv+rp7w51coSIo0TMJ9/xIyQj6PaYofsn4uNXBeX
GGh89UzMOjNB0BpkIbDcm6Y1mWv1OIKW/8/uz6fWp3FzT//hKsbeJiLJc50wJ2IF7WCRhNZidKVs
pGzPb0kIaPHBomoVF+cR42G+GFmH5DVhH2pxoMN4omzlAOX8TNbDn9RdhNGEwqymSvpFyfmmr16v
XysPwrdGHwbZeZccoh6rBP5dI4fQSDt8Ugb0gSbERR1nPdA6m8cJj599L0FEiW6xf32evJP74Lxk
6pUYLRxvY5NUmwDCVZFAB9wLZ2LrFhPD6KMIgMgVaZKC710/jVXzuv73w0G+lQDQlR92veTNRq8p
lGVucsrry7gtM/+n82t4xyzJ8/vocVTosM5QyUsCaYxniivvI4djjX0BbMHtDcUEIP3hz1du6lt6
s/HhY8XDa9vsZeV4bfElwrF0dynvyVRQZvC6mcOGrXGCEXzO+Vqttjb7s+oFhHjt+Acj346nn/iP
Ecux7r07FKe09W9KQ+BQAcrhn6vaXLA3cjVbODu4z0SBdF+ToZ3+URj2LKQf4RbsfZLHaHztxFmW
zCH9j3Jl+cXgG7q+QScotDFU5n0mCiDJYzCCE+ccZsq5Vn59TCIvD346dpRtSCn20uzE0iFlODnJ
gtWUj2nekHYYMFXZiL4iiOlI3R9wXQrif5Kvvdux/Su+9hLdyD9Qrejowxk7Zy+m5meQhYCj0S7F
SmeqUm88VUQPrqkptpBzY2Q0s1vDRj3FjQQ4OMR6ewR69BulCnkpDQKWzD2xGC+PBRaXcwZglBqG
WTm1ccxXucNKEUgzC4cJo3hMbIxs1cA8UaIhG1xasskt8QelP5deCkdDYXLyEZh1F9LJ024qv69J
Y7HKDWcpCrDo1pTPddslGzqybGZaalGVt9E99c5f1na5e505yKHJmayIWIQS0GfFL9moB8UpvZiv
kox89tPfg8AqPWhHeoAUWPZmw3GWMCcrNL/u24PMVv/KOFa0rW9TDtunPCcF3c6mM0T9z1+0TFQj
50uf0EVhzKKDUEeo7GTEm4mAdqU16kG32D1MuwvOFAxu3hD3fxoH/bUXNsxmyRCjVSW+bKLZUj7T
wpnr74T6gyavkPMcq01aYH10xs3aEb9ybMH+sweXPcA9Wh2QYTb+TmlH7dpHujdGC1NmiQXXmObI
Sf4C56YAAg5rwz9EfArOdWpUHpFVE7Dek3a5pIAQp1j+iYqQCMw8FIEbz3P2NJeLYgLWEsdJ+mez
feNz15wGw+wMPo0LNwIdQ6Hn4bqA2DFuoZnHEnOxvMfVFoaK289wI7JN5BwH89C9wHLAEOxwz2Cu
HJkTPhjbY2gqVB0jkF4jCTMd+DS7kxc2wCCuhrGuIDCCXWIZmd5Cpk3+Lv+xKihoeiyPkLl81RrX
kmkBy1rp++ljhTlWnFUI4Ma/gbH8fxk4+D1AN67uCwQo1tQwk3oX0oEZXWPne4p2c4T6SavlwGpj
9JBYX+mHSnn/QwEq0mWk/AmZ7KBDmogZKpNWPSfMiUdLHvJIO6D4v4KgYCiU5OfbU+/fjWwO/6/B
fD10wUzBFtUTEhmA+r4sJuzNMsDR8Ptqrev/cccv+2sQGHunRiHgq79nfvEcPWyoYM5nemvsofIH
jq2kynR3DGmvuQ83ggvuEHFkXri4u2gnT63GpCK3XhkI+twlN6N3HKMGN9L5NuexvQQtnUJCNnTH
F6ynHwcyqQclzJifeRbxShsZ9lsgYlJRHVPjLa2WHTwEJc+aVMt1b6e4ZE5CvC0Iwv4axwuILptn
wbT5XchRn+0PLk+nJIw19N7tjQLB/f+nmIg6NQcs4tYTzIBXe8/mZNR+DU+31u6v9w5cfw500KTH
PWakYytfQZlg7PFX0I8cUSt8qiKiYtVg9DscEgB902ZWRwSz25SrjeG2Pt+2mCkryYPERfCWlaf3
ZrSMkC/+SVGTp6ipPkHXAuT84Q4G1l53oBCBQMXuIr1vhZcvMxT4C7dSm0cx5+CUOHW5xjb39GiV
La/k10TXAERnN7WJukXMyV4WWeqWH9cT9xdicgp63AcPPG2TOVKqm/15Dz2110BRltF2rjcx2hz/
pq7SlXLRdx5b9TAvbY0dYZQoIzKvVFTBO2c4Vr6SA4IrQEKlP1qV23lGVYvLq3EiMDZqgT9BHabs
vkzpquwdH/juyTNeCkwItdKGuf/tuzjmFRxyolMJJd4xD3Am17z21eN+n39f/BgjRZARs/fBs3hp
OHMfUGk9gKfhSpDoINeX0l8cbrA/rC/jJJYEolhGjt7kdjJPvoEa966HBzrjo7eXHGPZWAmGxk5U
slKUzvi73+Jn8A+OP6LnvEUUcmX09gKHtlrfBF4clJi5hKDfmM6044xqZdl+m4ejoU1N5Hc7CEhK
IXpkKJY28LObZCFLLhEq69Yks3AuBth7/ZfayNbBZmhMzEQGDHa9Vl+s7xNFSQ81ki70RCrFRN1T
uEYV9VGwvZQx2xNhv2p4rWyx27DqEs8X7Kj0O7QrvUxDr29+rjGbTu2FCCjAT+/sV12WJVS+gdgB
vy7N94yhhjQbkKfUVp2QsxYxZGAupOtAf1gf7sLss+18OmqFKcE0mPVrgYjD06VIbPczqmQo3JX7
Xuw/deXisCQVC61k2zcnrsJPxwpU/99RyH7bMD4MZ7lHuznX8XkavBCEUVujVqUeHqoJVmQ7hSGB
q31bUY58tB7RKBlbxuNJE+dogSJrMdOOZC2dXDddhBDAoITaWsml1yY19qJJE/b/jV2f8mQpH7hq
OJG0yzBc39HeP9u+rzRvyYBOl8If3dNMUDswUzP40Nw1HE0o4m11/IfaMdWYJK0JF8d5eyhtDkpp
dIT02F4/S7mM2/h1VRlvIXca6t/N188tIJCFwRCUdvN8kMIETxPwx0U/wDcpLMearlKV/9QkNyc7
UeUkOWMeks7ruXg5oQCZNVMhujZylQukQslJi2fenR8dARBaJnBXXvUo0uQLc4S5HzPr9lnfMZhL
Pzf6qRXpe7KfzHvIGYYtHFjNVzS44kXMEhZ33JJDotMcsPrMsRL8LKWiFoXiMHlcMXVDMYSWCFDD
b+nuF01egSDekS9ZQO7l9iZu/9npqJSt91jA9QujoNhMTxGFU1ZAWfZ8OQi4aP7WTTOfcvrKhBih
RxRHLYNnrUqkVWt03vrl4pFq3zXik/bP7LZyB64wOuKneDZKbHiLMBls3IBBToAqrsPqBgwPILQ2
G1VbHUs2TApevB3dUNVenCJNt1i74uhCustNiNpMfI4Ab3NpgD4Ff4mqgr27JtQ/RwQSzRKuP+u8
FTZfDp2Km74/2nkyvr/XbG3xfHvN573w15xgJ6j7x3AZQU6Rghdp0X/Wuu0wBNBQsnUkGP48+BEz
hEDNHWY+CzRwggb/b7LzzcbEK5zbsXaBARhJKHDD93MMGc2fBk7BpQHGWya4swk63zPvCDwcsPtR
fd2o7PPVqcPuEXx40MdtmLvTJiChYrEOFgBrmkoNwv12UjhHaKykMzXEmP288gHkDmlxDrLaYoAY
QkJ+jy6SkftXy8bulchSZANLikLbdSBuevJjCT075wwVQussHM8sYC0wdjbxTSY7T1dPdiDe6l7F
15dswUfu4jvuab6B4QUJrAmj83hNiNrVTIaI5TLZOR3Y2144zmmZL1u8L0iOiCu/ffhMQIWq4ryA
fTzxWS3B1hbWyHkE8g1SVBoUvn9NExvx7XfvHAdGzy4QDAxHQbfzWSxNUnZofLFzC9m//rkEUD+j
7J+M/1ItLFzy2NlS0q+zJD7m5NO989oe90Xq2gmyxcJb8OGqasXhyAYEY2D6H6xxSh6Ut9MlH0OJ
Tef2YjoRrPEs516jF+6JZwRdFSHemBE5/mrEhCMpOGNUoe6S3AKyG2SGjdU0D9f5RYFkh2oxYL9y
kyJevXplTGilBBC/cSNwh78PCi0U5g7Sh+h6SW7/aRmQHk/TEeiPWbntBv6c8qzm9ZDMeB4g9sck
CKBJfgccNUjPkWKTCSKO0cqFCn75dxw0sMIvQ5ZZXug8BrqCWnJyt6rg4x27DPjSeVxF6sZeQM6b
ZzTWPmnMcZ40iAs01kqEwiCLWWYGknVW1Li8prnMur+jGnGpi0UwV7yhzuiml/f5dW36czCEJ+vI
YEdhWEoo8Rok1K5jm4m9rWNwBfxZr5o4zTAtUNTSDFbumt9bGpR5grN7LnnEA5uVrmpIAnlAhljX
ommEjgTM3zAIfSDcEs1tyrSVywhPs1KfhvijhTr1ODB9cTIqHwSLfiC84uEAelPSREF1woYR2Bb4
MmMzS/f1ZWF9XlbR+TwAd3ARKUgjmM456ksIc+krXW04WpmMoME/5dOJheFFT5imBshIQWPfBc7s
hr/4iVuf43zUvYbO5DBADIUS62rzoBscw+G8uRi2sYtHSbb/sMwMC0zeADNa6WQop0y9ExvF4231
FpBgSiUPAxQXz6vvODnSiegnVJHGhp2ZgLLUaNkzQsmRZAEvVki/Fkk4/qPKiSu2o906QxwZJ44D
OkhIzmsFdr5PeSQ+ThYa2FMe2iD6wEDM3eyPGTQdVzReX80+KnbSO8FeMUnbKR6+AI05Dksk8+76
81xSu+j5gvbDal+mNgIH3tZ6Vt1JPHkc0z7ME39Z8XEOc3feVxH61xTmhF5zbHNQC0ILsudjXOsY
zKhmQOm2ov5aFu4voshECQqdMwKl0oiD1Iqoskz58ka72WjSO+NcfoIEDiv42JftwZRXxp2wvhw8
DxvZcfqY8NoKsHI7hzILFjm8+NfOsI3NKOXtDsoNBI+nyBVGUKZonn8eW1+82F/9Ay/jCn0mQ9Ls
N886C90k3OEQYaNCdkE2J3UbnVXuQ2Lp5r10mdaL4HoOvM7Isgr7QWVvzwr4JT/YW5/06oatg0mx
DEK2OQ2If1N5Yle80TzyqnIYM5n0n6sFrJFGkfaod8iXtGr000MqnQXma/E7O2cfHvwTwO3vCWDf
yivpTNJqz847MmLlb4DYoysnyckZtHN1qe9lia+uIJwzwYKl4IbIHSAALzqa362sYydTpHnwRaMT
ViYjOQDdp0Xq399kO4kL6fxX8ni97EdIr5zN3lnadMtCqju7f3DkLoGINhjFdTjsfX13dwbm3TEK
1RaRwPDij3/ibSX87uEnaqO5F9T3yVqsDmlC7/8LNFi43PrRRfS+HyQmgKnJOLh2bRfi7h31t4zy
0iDnzmNgeiXTAzo/2KJCfcEkMhua7u21Og/tSa3EP3FJ2fQT5uYRQN3iG7oKSs1L/LRc6Jxk1gad
VeoX4gCnRTrbBIRwz8a12wyTqjZpQZGGWRSuxrzGvg7tMoUTmP9U9XH0omPj1hxzAaINmx8zcfY9
YY0hcyXZmpa6UslufZ/90VMqr1jUCC5RsSeZRPO6TXub9bxCp7+1KxKJ7vmyQpphyu52nK68DN7a
N10kHgJoQD9f5nyqEVouyPAcBoLd9TxBx+IW6ZjpuSt4Myz5SKkQBIQHix73NgfEgnjYSmlWTCDo
binKcnK9CPX2PbbI3+BSCfrtLZ/I1vLkxKwh+Ihmqv9rIkA1mmVOsy5oiQ1VR4Geynse4B3VLPM2
K066rbXwEfcvf5eWG80dw8p9c675LGUkZaLi3BY+sOLF2bs/EfJ/IFQ/HBK4KEFMrqBF3x6NRvQz
Yr8w8YUduz7NjkvsX9T6T4YrnwJT4JCK1VGQ6PeKXRzXbJ3fybG9Tb0DGRQzXJV1eW5n4/4YEB6X
zFDDl883Uwu0KtiOKATlZzJjdteG4A0N8IoqaJAiC99+XnhHGtdqWOLijCZLgm/+7ofQdJrnsA9W
sXAh9rRlTyhas+SkqubY1lVsUIc/E0wT83VYW5jhr+zUrT2a0QDsWO7xnpikC2m4UQa23UkHQ8iE
+y6pxSI7nnvGSB0OzmD6vhXP3C+lul3lKHK+kiSOeos1NHVXmdqSUOuCAh1hLuRJ9ZIlQpkhdtRt
48cw9HVYyVAvSBG3aD7QLsaJEDb40stYu6slm9wyk7eSDlwOfNPRfenZNduPvIgwDS2UUkhROSES
e2YeAoZmrqMk5EuUGTEcsLTXJxCyc8FXVWKq6B00jHp6N1rQdcL5nHuLH4NB9gxrZEdaIs4T+q2h
1170urVbAooNb8MFq/FSoJ12/1+Unlru0VACAQ0MJEiqxvPKo10lvcl8OLrjfhE2R/9itucEACyn
63rWCZmPo/RkT03BdUXCNaHLR5mAG6kMA8yRUsUvUyxpwkJTXHJ1ER3aOs87gLtat/4bmnnLpdzX
SoZ6avNslqXiH5CZiVVby9Zt7qFod0IQ72cpFXWRRL5QC/1WLulyHhiNItTRfi14U8nKfnUaVtPr
RKd1V0t4M0oAeFdTRVICpce09dK4YdeWzDCr9mk6jtT1+IrFJQLqYL/17t6tUDFG3hQtT8NFfOZi
O2Khvvpr0jEKkmsq01m9uYn/fczHUDRvyjHXhRw0CuYKDnIj0yPJQj5nH1cvxQPew4tb2khXkbD2
UNEAMQITqofdZoujcNL+zP47LGg4x9fN9wNy6Sv5VSZegAuP2GNGCba5ktuVRKWccXtFDANEBsMc
UJcUJaHEdMWo5RXlU10TaEMX9u6YiVm8bnjPtoJslZmXc0+DlOXY3L+AauZ1UQLYPn2mKHVbPEQE
qrGZceD+Pcm1INrBlM36koBxnw6hk9cy3VL8+k/KvPPZNRANL+w4zQHYugGALA+8iXu+08ppHNgg
pi8Oq06b80iQeL8u2kchZ6JH81qfxYJjcmd4p4gVeyDxwrqadlsgcYKSJJRJyP2v7Y4EIMZIJu/1
zg48zLxl90+u9iiFq6R9YxJArGf0V1Jhy/w437B6Yy9kpp5otGA4WohB06FJKJ3VtWuTwHtVQM6H
yU4EG5c0ZDNWhXAqoKhcVko0Vx29P315uc1Pfwq9i1zeOa7yshfMXbQjVfk9o9HPZpHpc6UotGC8
nB+z4uh2rhLIeHeX/xgLMKDhkL9JStkdk57ehAyLLNg6fPYoGBFHXMZoUob4moRlzp0DqFDPWZyC
BI2Hcf3yBYDmgSUeMsRtLiYumPscKlUEI5U6NtK/d80LZzrLxGS9TLIEMCk6HB7HXN7MgVcFiPOC
LNoBvQ1UwjzfjiVgVNImSqRx6TGdH//+RHYhIGJP9M4Hd9Xk3HZ3LgLT6JW1+197WXC34YB7fLzM
oaWIVisCFm7aN001NDNOWunbtLIHV3mQmS0X+6ojOC0tPUbyaHgVMknJQioYfZxPz6wWRYf/JZgy
eVUK04Kpmo4Uh4eKAHXFkmufJSyYJwr8S57bdDi+SjiiaXTQHFmKSqryPZJGgP8OnueF5erQ26Kb
J5Cn0d8iLhDwdxBzE5GLrsNj+0bVnd8/4g6tpw1pENi3XWOSCY3N9htBx1Umb/Aqffy7S4J9Svqj
fsNqm9kEWwTUq46Zb0Cb2p+ZCMr9yOU5OvQCIuWm33Sc/YYHkHGn6u8TMItgpHyYlxvtoeMm1ObR
VJHajsk30QCp9+w+wmkMN03INCeMeRgvs2jJ5E/FOVnY7EQ5oveVOoZx0uusSamcGVGSEqFTZjDI
KC118RlxpWiI8RjFlEjfS+Dx+KKQnG1yf3dyTp6atSuoaHF14SSMqWhXGTOPnNvlq8eMaMHqqHgJ
MDsFw9hXoRqZIVhG4lSjNvZ7THvmiqyuMCZhlYHQzMoLlz0+orc74dwaj1sD+akCH2n0OOGZVlZ4
ttUOXIWZFwNuViTZseKYIcvWprV8ThsxKOsKU2rY7EJt83VB62o5xzTEHJTyOuHkjfh6pSPmRVEm
K482+Se5I7T5HihdoYNiZTJCm9t1d4MHn8ft4Lw8+VUvYKG0QhWguvqwxKrUgcbA9ZG8EClS1WrI
ekpVP44yBesyu/c4++3g7pes76sbtV7D6EzR+Ib2UJ7VUnSeH48RAofB7ZH7UPstBTOyF3msA57i
k9AStR5dd1wVGwMsuYV6HreItJsUHry/YEmJyNDokyR1g3LOLwbF7O/FM2ILLIrojn93afZHjEIV
QOYlNS83sfB0Tfy5kuiEqAp2BfajR00L7g9OMhqDwod3dUpQBFOLee7oOdUO0CwKkr8Kysx2gNd+
y6UMURVozKkJ9GGs9Pkt7xK3kcWKlSfMQ3Xu9W1q3VWIJJUc7aWVcplLRr8i1waktrXfGDJ+M5Kd
y2T4gwNzYzaVlEw11pr9zGKHzdeWHxbcPIdZNH6bKrk+rIFJV8xpOwHsWki1fesdgxcARSkfC63H
Pf/PTB+DHrDQElkqbBJQ7kx2o8kxTFbUfLust29n50KnZKIVRRQmNAlWnb8ZmYt82q5ykOyQs7oI
VR9JXrqFaufdgT5dB6XQcEFWLUngbkWCpPquY+CxFUzWIvOKpX1Y4vpzfrVc5zPTTpMTHLD7Kvr1
6AdjqgmFuh2S9ND1/LjBa+EKRpdY1aa5Xujxxvy08qweqXgI9MYcLu7pg0uN+08irzQ2filc4vIQ
MH6Y2D6UzFo+18mzZa/cQo+KDJxp97+yHEQaUxzOhDr0H6rzLzh+x9xaHt0hrtCWLzT8/en1QD8j
ioC0Z8pX6lab3jscxOxXsA8LK178HnTSpRydCK/fJZh26cswibTnP2NBGqABk5nyGddB6ppHjJhE
b1nfILne2cY3aYlvrOoLUeh4y56IAcXTHwfQnzAewcOILMuokUFdAznC6IG6r08CqN+dtuZIvY6y
SutxJUfU22A43rIfwS7VPopQQPOCGZaurWsoJMvghGlb61JnR8M8c58hR9o4oAEMVqCE9/GlV/0Y
nZthRj5sKFyFqu7tq9vHImyVMtNtPmT/UUuLSEhm38fWFw5pmQsbAZtkbKRRohBjs7QopqbaiNGH
VtcpgZnryoEN9vo384/RUaN2pybHapZaCTLJ7+nJ9Xq6k4i9JtEiNbkOJO9FUMQgFYWpakz1taVO
cx1cNueRIe/weARQSqJJStvaU8s7bAE4bnob+dpIB1JBaDWC1fQSWBYu4qnmuw0WAnp2sLSkXpWH
R4dTuLionPK5cmeHSLUj7QQIRfvu1B3rM3vGYi1jCXazYERrr08z5asM8eKpvEdQi7+X0H7taqf1
nTkXN062N1rqO/yiiTlfQHvobfo1+Slao7Y//F5JP6a3nGdFJer+P3lb6VWo/i5eruvvsfJSsZu/
OrFZLhxS3Xd52ImcTGEB9yEleMfyMGFhgp6TJ3aE5Tf5QOfwRbU8RiXPBo9sicBzP5VOwbo5CBSz
C/FOetvFwrf24F60NDWoycW2HdlrvsvQSR1iYa4wjofUXKR2Ri3mnx6xbHQ8RWjBF/ZPXZxWybSf
RycGd7qJQoUDrOMd9YyZci113WeU2L32Yn/WnZVhkn/e7jwME5KfKwmFUKkvcW7KFuSp5BkR9BeL
OykFFEWJasC1GpM+t4yNNt0jLgY/BMUGOF7idLyWPMS4fNBuJlq7Hg9sWKX/Cqzzg7Q8Y4Go+hC8
X6KKFFphtO7WB6ppqxfAxCBFGRvHgLEv4+JYe+8AddlytZ3anwSXcds+bWvj9d2vZTvKL3cX2xkw
ZGVy5+phix0JXZ6HoCzsfpuurv1HA7eMOO/Bm4fjfKzA1jlSVpF2TRrqQCQjX7+8u//0cyOpuYPg
lxzi99uDCW8jclKmvDVUByXLTFhx/WK4prjhyCdJiyhG24pDD4SOv7XhiXjEC0H4yhVO2fuSKzFI
8wf68ArELfBQefFW1hNwPMdUfs3SKwmQtp3dfhtBG+0fpIpBjcnP5QTLDjzT9fvqbvnQS8EYv/kW
6l4luR9vHbBEEEcJAEe3bE22Pznm9QgcmYABBILmIq84Z4aDCLudVo4fHgDr4HoVyfniG7aavvlE
p4TUg3JxNEafmv5pykldW3bdcK3ZM+rzxZtVACSdlrZGLk8S8xhD44XJIy+SLTEkv/bLpG4fZX4x
jWCxJIA2HiKE9c9rl0vxKWNbxJYn4NUHPw9SCIRbyk9lvyQcsIr67aW+zf/8qnajLE4qL9lfBS9q
u+ZLsDXZtb75+YPmA1XHpgUa0fU3YKAKpYce3yNK+ZefXTtfjOLkTG41r7EfiW38g37nHSkC+/kn
MsbBSt1wrKiDm1iZY3fW16Y1KLGxhpOBrb7zWfqPT4nugzJQXZwHfb4TfoAR1CvGcNKN7za1TpEV
vo58dJBeRpTY2FCcHoiUWczsiOgXEtJvL3FJSNA4tH9tNy2BAXukq3sTj48uQIE0xaIP11nWNf9O
QPMNCT6ZwffaktN01MI2YJfQdtkA8MzHDG2L3YRz0/IcyKrLZG4EZmpi7vzo/sx71aEt7+ipUt4e
rGFh/CZda6QIEaG9byiP+xeJMhKR0SGzjGgILoaJyYyADMfYVEZD2382T8SjyuVmLBBRg4UlzVia
Y/8ygtmc4mlCkNE6LtKB3TmYCw+rJBr8LeFo46NaM6uX+mStOcdXIJ88K6iZS07BJ1PdaPX2g5Uo
5vioIiZiyck1nhyUa4tsR9olROzMZw/lCrJZPdN8LxXQ1fj6jskEr5RZIaT009ykMZBVpqWO2bZl
hV3bpFB+nybGbT72FaW7wU44hKEhjd1RBfL9ryIy6AAYegUjQZsJWZFfNUpO4ArLuBZL9o45U1it
yFoUgSkwRzKKJpZrTAURu2SecK3RHhzqGRnvFFm1teTsBA3XrbANBMTYrHtl58QMCNcZszBzl6hF
WQ1p7ZU+BPOVyC0yH5kiWIuMNWyliE86G0ijeGoToqLD8b51tzrjMv7txKQRCTKEUKZu5UY19sEA
4dnDEzDt2kLRn8aA4JELFWq9wAL0YGY/vzzbB0/ondS3sJEQqdnIYgN+tsNRuZFSX+gDnXXTR450
gM75bFscyguKPyCOJcdbhxwGv+DUPt0cGnkmAkSJGyQIJdnroUZcG7t+2bwKMoegKUMYez7aDj1m
69dYgAl7tIqy2O6jHte/5i/XZU0APVBexVSoCE3sZdMaJ5WO3vL16VtuG9wjBr4X87MDFK3xI41b
4F5g1uFu89FePFxV1bb/C1VApL7CeENVqvEkVyxTLyzomIAyWMvox6d+AfB+Jntb3rrHXZwwzFy5
MSsU+GcZ44Un9NF5OYnM9oiUwJjkvN1uG/Tb+Nf9XaqDi+6lijMGz5A8BBa8DWhbLQ2xxkNB16Bd
sKD4BtROdGBdVa60TEgKkp1K+ZcWfPHgld9eGdRU6CbEYoAbdRvmc8/L+xCMXarb9/xFq5QdiCWa
BJ/VR1wwQOWACArVW1EoOXjrjnXAkA8rFi/O63KWEvU4/EbBZ08Srxf34I8GMGl8KbgjLyhjhILP
hOe+tmtw2bS6cmbP7pvB8s5BIKEB/qaFWfUZXGMK2CuVk2mYq89GnnprMcjtx2MUw887O+oGSCwZ
Zg2WtJzpzvSVoMa4j+Uta89EJ/5yAABMbMZeykMQOxYNHElYTCU1h6IXYF/ESK87UPBTmo8cdJAH
fFEpNSJbHTtX+ty1oCNlLOIceZk4lWV/OFI9Cgjio6DEqSPyVWLCLBt6J8vr95OjWA6y28EnYpmL
YE1dl6vbTSd6b0tjK3ipfVAQDSZLfrTtTtd9TUGgkcvtvH/vB1QgNe3DbXg3VTwcu875sFpE1mV3
Xa+72AhA8If7OyLoNlSU36UjzaJFEl/yDNhurFwwY5owqwh5F9s/2JT3+TkxXjBenVd00UrlYAot
yW+RiT1fEKIxg+91T6nddf2gtX/K/Oh5UeT99DO/dsnuwYLxlnzApGxtIXjyZkT9t8Kbs2LEwwTw
Mgav+oytg3yqtiMKKqC0NLvY3FDYAvGzQm0uADsiFT06yCfjrR/ZjhjZ8KdsmqhBwUbdugN7b+Ls
DIzH8SAfqPGBg+6kY+n79yZ2P6ByjEBycmdJE7OMcnhRCK3VkRfkd3vjsJphSAVfhmphwNU0UmfO
GDAOpDAl542vPhhi+6Y8SVZV4tqAKaYSkOuCvu1oA/Qdh/g8E5rCtBuaDm8P7adl+Af+7H+/L8N9
kjJ0CV5QlmwUQsCkusjeLVap0XMTeFajw6sz2f0k6h2NEKNe6ZSy4eh/7EwM40CN+4r5a87wLFYZ
FhcnH7gGmrBxPAR8qCOnL38H1oYWTiY4GZ6O9m/u1FxHqixzubeFhn2xyHGy/Ss5jdb6Jt2F1fGD
YpOYzjnc4AMqAPmlncpaJXu/L1f3YqzIhP2iLmguXzwLF08/f88WemgHOqL/ftNYZOVKI/unztqR
fDgRtLJtzxkqB0QXnbyO2lTWyFcqz9k2yl9xO1OGK1tA9BPbEcXMGxu+LPzmudsYco2TVAL6n5Rs
NiXj1drZkaaKROHOHX+jjcPvCy3P9sCe+k3p8X5c84caqIxbyu8DGcda/FBkYCJE8jEzskOmbxVk
EVtx47Ep5ednoSpcz7QGIuKq8/k08jDldrXXZ9hR4jpFN38cadrGIK5IaS2ufJ+Khfvx82mJP4N2
6O0HDfr5H06PHYPWMw3shXyMjBGxYGUTZ2Lf9+a/QJiZi28wywtWT3dfEB3ebnNRURTIQVgs5nv3
7Yfd/wTABBXu+1828on3i8xVGSTJzUMCnEi9/6yO3CkMj5a80jH67DLIpLsix3UIQaXjPOew8kfq
+qa3IftG1bMFKzU6WwKkNsc+MICMSRdR76lPFUDX/FGUaVb1d8XDWkRJW0LeKGUMADy9g3hkeJvd
wu0eoFtRvSk217VfLtjENdpqv3R5EnIwsx7zsQYm8ZQGaNKBnCI1VYU2aNaa5sQZJSCLEDKozjG+
ceMjic5eYIdj+j+i8eaYFSqvHleCvtEYVt6GXKxVYB+J7ReKlsFEbt7rQgJn6jJJzgLICbbjdK1P
Fe8+97VJ/QC74PteqwsOLxDXKpTbk89w82I34WKNcId7njhQ57qQXaHyjKmODZDNRjckpztM7kwl
JLsvhlclSoShtD9IV/vi7hQj92MRwenC3+SZ58YeaGjjJ2cxmsG7O5A5NjVMaJK5TdxGeeE6MhQO
8LFrreI+z4WMCqtcpF17X4WEWJyf4S0hOgkrEjua+glQPF2ckM7HW5krL4qQFGs05f7BKz5/bZnh
RofP7+T4hp3ZIVM3l6JCbzhLddzWyaXf27XVa0mGkep/XuapzfU2nRtXIeTanOdBs9yzs2DDmDc7
E+3ZHc0NGcZtINxw4DJBHJMieZYyhIcmombdSIffwRAXIRFnFwEY75ZHkPxSRlZiJcbZ/76HSZec
H8rVraG8F4dcR1prUjMeGBXoQCQ1b+1v7srjRUKy8RbXkJb+PI6lHu+wEDVoErrVs2k1jpMauAk3
iY/fmtMnDfeLi0ke+tesnP4IVXHTkpFo6RHzaKoiFfdSx0034k5zJiD6IZ38Q20u4wjQHRnYyPFe
ycKiT26Zs9M694zFYdZ8h33ZdB9+oFJ/hm1dTZwURde4n541WAZXFAAfCcg23I5eKNzf/GNKrYEM
FCJJP6dI8iDuNAIJxpxAl5PXunLg/846OZ4yqA6wAVeemNO3EiTRq4YRJMW5cj3bFasBtnWm8UDn
CvJ94oaHGlIPA7qi7+9mfB/1l0PmkqS6d4RiQLOCKqhEQAFLpidRLUz8Hmea5BviO7j+zbaGsQXa
SvAtGn85iV4bHT46At+4W6pHfUOPJg9sFe8ij2eMSeAivNtz8t175p9V4wdYKJrBjMTe3gsZUxiI
SeFc3fQCUaSc8eWPN6JUod6GRDAhXsb3IKGS7IPfNL5Na4A0MY50L9vDl2onRWFeZ453dzhfLe4A
YrVRQVPNVg0Lj12yUx+34sRXcXwqsBzJBuocQy67MerZ+aMKnMuSC6ABdnRzSpOqawcuVpHe4thC
fzUTpNbikroOJhaFKTpg/ijj3OcYBG/w69KPVyKbmQwGZY3yfEal93b6zFpcnYx7sKgLVfZped3c
IdbYmDAkuuTkAbSTQ0qknZaS9Cg2VWuYlLKxpFcFuhMLYfAvKH+uzOZpQ2klS0rhUenucUINTNoN
EDjR+DcXhsrCY5NierPh9iN15HVMzvogfXa34ervSNmSm+FMhZlAh4/dc3P4tXeyiGUKj5Hb0l4g
ZLS9a4z3VWWCshNGCrWLFE+KErx+7l+B09UyDiGEXInJNAEGuatYOHtQsAa077f1tN8TI2LTmhw7
eh4mqYYHVtHQctgNi1I6mvB0P6jDx21JRTPrYNeesOuNJW3YOUsIlDV4zodSZUlpEhTsxnNCuvnx
J+OPUfqtOeGhVqBMH9eJlVprr4AscoYdD1/lHtXfSJH4E2QqRfyz4aH512VwjFVdXKVo5abj0h6H
V+bUIv1g+BQBVJKf6ZZlRoUKC6jaqF84Ita2hNoeF4IlbryF+EaLIU6IivTQxYA8JMYYC0Dw8XXG
2JVCM7bmAST0L/S1/6PHL5cuwGiyduWoLFKcWhsHS+TlhBJ1X0ttpoycUol7mW1BT2RM8+Y/9+1A
/lkZu8XDu2KQc0en0zRnrWr8c+NpY5ybOKTvkwB+pFhzUExhRRXyt6nYXiqHLB7/F5KTgGb+FJjG
e6pkS4jzbZZ89zn/YX27BD9AsGXWAr90NvPvk+JlbsSuQXJiohqa0POQUhmBFTNvTkr5o0V1m+8j
A5dmxer+E8YLHdvacBdnNEwsBw3+3SjHraqer8wFrr6SGy55VdZWdjClHF9Uu+iKFb5DXsjJdoWv
OV45uUE6m7A4UtmhnjTI3tB/1+wUbkJJjCxIcLM191F19NQg19Sg/BZJwVqHacwQINY5kPtjm4lO
dyxlyYSk8BgnfSQuBK9JY+YAxsutDD/92D+FPQF6zGNPKCDXg2p/VSDsV5it2x7GlRWksLvCClod
WOK7KrpWYe3m81/rlQIghSSxiLOSzn+4ihm0Bgd+SLBHL5UDlJjLE+HaQmfQNE6Rn63GTjp2IeFs
ZFwcTIFU9e7iMCOzeD8BJpT/4aQDHue1yCKUY67lfTLWIv65/rDyYtSpSv+1yFWWeR2I4HJww1oa
1DXvApw7NLN756zCV6TTMDeqavwOJq9YCP/CoW6q71/Yjht0iWhHEvC6YPNRy/xvqCXRrfzrwFvW
dbomsQb1NnwTRcrdim9Ivlf/Zhg+8WIAp0IwIlL8Eb6JONqZU42yp0AgT1UFIKaIiiHNuY8wKmt+
d9brGbmTkpsDDFSJ7C6voRZ1NxqF52Y9QmCobf2oalKTTPZPcxfZYMZgYvHyTjqIBKEl6bHkqPM6
v5/s3+A1C/XYn9RPq2WbOEIr+4lVMp/ZYHFnKrcQizauT2zEQPUOv8aSptSDFWnoflK/BKHqd7QT
TLf+qzfmIAke0M81lNuTGo1GIaSXz1rV1NDXhARBLTF+rorNYLLGIbTnZ6IPLByNkN5VsThHSnA3
6sbmNCa32SPW6KNJX0590tpWbkRmdcF/pLq1FZ4PdmM/8vCz8i/MWe4PFN9gEbjYEUZc36saRW3L
YtTvAnXrwsP6iDgXG/9loBtIlSvrGfMRe5L69oJGQVTHoCF7LdvhETurQENB08ILep1JJJapyw+h
Xei/WgrnfDoVHhkDS21+A+YIX/93ZQp6LC54+a0eKNHPrsFQmxgDQNEvueWmDmJgDqEgJq5kfBmo
YF1PDE4grPcv5szUJ6GQmlKQEdYpGKdYQJFAi2i0lJ2s4Xfj39P5w4/BEOPaJS6nQa78BPs125ps
uBhi+6H7OxdfVGMjO9qzSLX0pTIQnN2SDOdygCcANRkg7ak5iFQez3mieL9uN6dMi6QNLVnSMyIi
Ag7RVVzTQI/SWSdDiob4itT6g+E4opT0b9mq9j8f0+YP2eC6H4SiTki4doZh65fsQKxGcV59iMRf
YSlph9Egw6aVxMG55gEzZMLwz/DNeNC9Ir8pwsueps+O+EqTq4yqxsM4glTt2tH1POpohKsSZoBw
dz/Nhhd5DcyoT7YNbeirL4ypQtWNZKPhajx0iTVlCB8Rbcfa/XEeRHX0ryQpsxaAcEW9XCyUlLtD
TW13fPpXF4bfaxabyh2vRz5nyJVpPcVV0540rv3v2DF3kYCBAekVipyfwSMDZRqMQZHxKKvmOOeI
gQfeGr6NzxuSSFOCgf8cXsqR4gIV1oknBPRxZlIZZRGCSwvykuwLMciKF67X3r043p6070lLblTb
gd40PI/3wfG3CVjgtMop7dcQBlvinnTRw6HW+V6OXk0+RHvXanrywUMRxx4jDQRBghSNyLH89qSJ
U+T84f8VjF7vrOZ/BEo0xkDtuhLubZZUXcH51+rHgDcmWzARvJ86cZUrDR8FRkaQoXiXQfG907qr
YnXqaM+jDBEBvfqk/ZJnlCLFaDYETHAwxD1gbDjpC4bhaDAM6FwANt9HT34AFoI40wQknDV+Coa8
c17GUYogUR0ezx0p/mapODqcVtOV4fVTgwwP2yLCPSLfPYsswBFLE7tR/EeC56NTXilwxmCFq+xq
cq7v+4PC/NfJQgzGTCCO6IcTl5NCPCF8DIziQYbhwR7vHBCt+LDdwpTyx6N8HN/hhrH7k/hMdggs
kUx6hatARSvM9y6w//W+BUtAx99IInKpN/2dFNLj/xtQUSebfOBI8naot9MPJVFfYXX1eIw/kxFN
BQfm6R4396uKAYg7BKyHsGnQ7TFuolqqt5q6PNe/kOkq+lM1jsXQJdMfwdajxdlcvQZCOcm81d/N
4SMRXb0jS3mbJTUCETuw1QStgbEWtzSLtuXwA5upfFVd4tlu4RIjmjPTeu4sS8EZN4nv3CRnd3Xj
lID6jTvhqU0IDQX+FHBuzMDz6vREzEX2ZXKkDeUozsPnzOStD4hTU+n/4Ur4xGVbqoBYCAI5iF3O
A2FVFQLDw3os3o+/0MdHvaVzFlP9FAAqlPtnCH/FaB+cUbnqfwvct4vg3xUOjLIqJR/NSzbwxqTj
4HdZ1IeIcMV6KTeiATz+yozVhO2T6aQFbIiacYDTEfyAkBbwHRTm260lo6JhA2r+jOHZCmecUyFP
rPH+hMVAkn9FGjl2dT8QqbO3WkBD1513AAtVA7BaTk24ji5zvD5xZz8ERUO29rKHPCTsJ/AqexaG
i4bPRXVzQfrfcNU/3zX2ZtUBYORukFC01i0jG5hOyy8faLf+qfSrThr1IBnLXT5aE0gZrDWA5K0p
9Zqc+sOPqrZ8YT/qYhd5FQEPWIhAlXqnTDxB9SD6JBlhstqSlQkAtSLrYg49T3knqdCu7HMFNAbL
aTwZDkwah5IIGlNhPEtn+/6ArDPUlPgc3F3WB4eXcFiekJF6sgIasos0GdWJk4veG7pd5vKq9WSA
oeE97lW3kT6ZzSpta3X8+4jIjDKx7injhvOlDT5XTCcOmx8ZP/bIGsnxwjYQ32jUkQWTkxpSJJTX
Sg+Xso5k0MNntJbDT0WVr1dmoRJhkQyBoqEyjoG41/kFJXBUwxhltsbIcLa1RrQ8aXRkK8aREq2M
r8yg7dxG6ESHtayVogo26vOVK/xv5mKi/pM05TFlornNoapgQ1WF6ET1cud9OPH/ZKx6grDGEskz
yeWff4DVd0Y/nnz1+H2lzjCfoYBp05RAnjh+R8gDEx0RZpYRIi5LqZeSBh9MpP9UzMx8m6Ux8lQg
mfLKSrKcWmJ4xgT4eakLqdDgAoPdoF38/eDavyR0LLVitAe/XKmTi5e9jGOea5ee2jRCO8LTawp+
eNinyWh38NA0jeDOnIh8+SYqlkLWQYy3n3WKtUkLE6USNCEqFeXoGbeRA8twMmShsiHToOup+olS
VQ8XZOzvf2kEP15R3FlOlTVn8c5H1y9jndPx/GNGZXGnYWHGQhLqX5bfaljJAeZ0S1+dJ8xWP3Fa
y7Rcrop81RfStZyZnZgUjEmDFE8Sb8a1rNcFnmtq44uiyExWI/Fvbvmw8CMk/6mQZmaiGHj6HFd9
KcYZrY0DL5Gx6dnRlvFN/eG6eE5lruVO1nI/D4pE1WcUIiYy11xy3wELfVLziVcU8KllfnlGxCMK
rLApgig8uiDYIXJ1sQ4q+bDWsLVWT/u8xZSGpAD+GR7jqvlaLRWiBO5/liZ50h3tzhBz4GwwUAZF
0hfFHBf7VG+7y9k9ZbDIqcqJ8+48CSrzn4O4X7wzR93No8MaKgixyv84M5LTSttPNoTBfKTGIzff
pWYum3z1AJgPAMe1eSceaF+xdwfjAy1uLYLQeD4WwTAHtBOeB1JSVD+ilNXNMw1MEHMW/A+vDh2F
BT4hbQjHLt8YT4XRWq2bd8r0j+kMEjm+yODk2A8TLtOkrL32wkJ/cLLO+Z8f/P6mdpHPwnIn7eky
IaSuLmXVyaVdxGv2WkFj5Jxe8LjtztI9ODv2xgTm8jf1M4mKmawngNu03rkIscPajSpPlc3b/nvS
GJ7SzJB5/fBsGDA0KfuNP4ZadleE8WBbc8bjNk3vrymqXYDAteCx3weji9zI6tXqzy/g2U/PRC4l
LZr0qH12ZB9WFtTNXCvp2JhDGOZFs+Ph+1UPyNDJZMr8+JhcekVD+1g+jqAt4tmRVvl8RFHUO+8l
c7EOAfQ7epaynCyAOOp/qOdwgKLlJB7iWDov3N2Ad96dcRe9XfudoIwMXjEXLB5Upd540XIH0ULi
66NXO8nx7ZE2hYOfafiYWhut4+096COfhmympWtRjztxi2K8VbayjgkQKj3+A6ixAKJDQHdtiB/R
qqzHXvSw0+4OfWzDY2fh+UPiHmk1kSUOK8n2VpwUta4oQ3zSrtjAfZRvPpZZaGJN+mbZUwmvKko0
FGtHNJdJGaj8lCkUmSZ6vJwS4O2P+AxwZjdOUvjSYXnaBZkSqJ7cIQLsKKLZwP2DPUkBP/h2GSl/
F+/C7BrTSRMa+MwSFVedm1AO86mXTK6tS06s0Zg9i02BV9E163sO1vo2pZ2/O2FMDLcIqnvxkU/N
KDIRJeoZVyOLf3yxDI48RKWkdHLowR1GJkRbzQAIgSP+g08V/YFKo4fHlXnDgvc2IVfpU8VfxDlm
o9FIkHx/oHu1Fyi1+viV2FV5UtZTyr9/5qFEvYB+U0mj8p7T1anpegmB79mhrvadYjF3/R8QA2FK
+ztKDJpD+JJk+UL3bMpKazVSKVgZXwmgSaLIT/1wHY4SCvL6IhCjC5PyZI9B45lnFDnw1EKMKAeF
JGr5CzmJJgACn9gs7uTLlCd1W/oxEBktdT824OZz1rdhWEEotMThr6zmefEEB6ohljvvlwenv81a
K+73ZjvUnXCZVBTXSh1e8ryc7j1FrhlEmAA2fzExa0fp/JD16J0A/b70Z7keefCWas0bKnj5ljFY
ktfDjBeAj1UjkNJdE8P26V/1c44/z6DhqsiGxj7An3Hsvq4mY7G/HtOoehIriF2u1NmTNrxB/j4P
NjaUaroP8yKLI0cWDbmfk4cieTUqO1tLgZYa1k4clxDkKaEm0/jzSE5W7o1sBXtRg6UUoHZ0hiBT
UkdSOIeEv2a5cfKR/a08jvMMGlHTocN3PrZg7i2g+t30zd+KwH+kpQ2P3yCku2En7tB+1yUMQj2+
+HWOB1qWjhFOVs+6Xk1ASgDrbrD3HYZ7f7bh+QEk68jJfckOW5KVb/JzJ8Hpn45Mlv1up0ELBMXP
NddfBLmcl9ANKKq4NsqYE1fsnNOSjqK4m/RngAgRuYeUnneN3IBpY27qeYPGRRVeIaC00kH4kV5K
cII58wAeu3oyhEwMINUohnykEAEhnckbY2jAwPjYtd1TQLbrPhhmbHmKS9uoZYEqGpBfXXQke5N1
OcbJik/sCVFs3rKkhjU5A93l2eLr4aJGhJueVJZgeqnM9Q40UBKHxtw8qUfGyyf+apcKT4jDHfpL
DVZF+MtdDsOlRwTh8peK3fvrtqiJqZCwH6apSRRynLn/emz/dySTjCRCJvyl9wbCKxSKGHhkXxlc
uyBlipsxrnDhkWyMFqzo4BC/mUpphG/MDoRRRzPmc3TIT49Wayq/I4LP2G6k4DycyaZ8Cxc3YluC
JcqeO7e42ZCBwegA2IV95vAjOI5vJIouwv0b1XF2uAlnDmogTa6N+Zv9gEqt67brCImA1PFpMfHi
v9W7LLQ+pYwzMXhA9W53CqFjjPZtcncle6eIxrqw40cOZaUaF6Wqc4ShPZXoqw9mFKpy832UCK5J
NGJ7q7LP2dhVWr9kt8zfDsb7BJIC3VNYQvG6VRrytr0IVuYFoXvi1aVbRWQGp901i1fROvOBJVNB
m6GN3uIWqwHgbqNlcwBrf6KuwaKm+QbBkj3XwuRfmZHSH6nK8nBccMtuhPQxLjfAXcMhaS+dBd9e
wlH2o3qt/xVQYL8BvRuXj5HRNApbqxNP5EUPucaKgdYtuRuU2ScL33qHuDO/mIp9+cLPOBx78a9N
a51iownwSG+5o2RyzU67nBl7YmYsPk/vTKqjfEJVa82nVLp3IHXXC+nw31N6Q3N3BJZeiNZg4zln
vXEiXv6URJ7sZEDp1Vsa6kOk1gpwMDL5TbMZPstUEMF2aX7L3/WMWXJ7miwZgUCf4QpTH0I+3nq3
b2ZI4QSFheCGnZp62bYyUD9NnleHs6geyDpG08x0KbFyEKzCrImKRdRLFukZxHvkUmwe5d2p1+FX
q27mHYPVTFRuBVAKCFOvEn1OxpJdpOM3bRz2eDY2+wKsuTSMlcABCBtdSiZsZXaRngBKJQHUBd/2
SLBEVG0TkxLqr28WG3RfwTbEjZt2Qf6WXBCxvovrgswdlfXGGdouMDHUbOjWMDMPVrEiCnhL7pUC
4V/6b7VtyPo49YFykNzhb2jWe4RwyXSf+2DsrFzGio/BCXl3Wk4mTlbUzh4Pfxk5BALAVODpXXZJ
T1OoZLHiYLQ+juiJBuAOAtP+iDoklIEe9uyZSnVJ8Hmf1yfuyX70XIX0DQtlAZMOtrXWB9//vnCE
wiVQ7Gq0NbNpyDKAgl9XUZun9pWlZ4IBKd49loYDuLkMOqlSvVvdKDEPKgItPJTyEENXvU9hyekc
1tZ3ghKqtt5lAK4ek5VOPMaIwIUKexn9dYhRUGRf9Buw9TJnGJ+2NMQ+Y9XoonVUjWhbgguwkQQB
p3m0uQjpBjAeMqISLdkYXxGf5KHNMxKheN7e0Suj6R6lGDuvdg6n5uioC/O72AkeFLNfB00MCv2A
FeRGH0doIXRNi+FVR8RrvGKjNkol5ETqCX5Wjt1SsGGuhP0eI2MpwSOjB6MW8pJvOZASHsGgUu2C
zYjbs07d+L9NE4JuB4BTdZ8VryGJd/oE0mQV9CDImCwG1wgY5odgsvh8qPvsO4rzO1m3pJO084kS
pqwfbcVJcNqWPk/MCus/ODpAdzA0QbytTssNl7nYW91k4Zz/q8vRjI1bf093GLEILyqVLuQSBwgB
aTyPZUxqI7+PVsjI8kFAIFiqLAZPXTSgZKdM+WsJUQ5Hy6Sn+eHbqv1/1pZTngMJSOf5Nxunaiek
LWP+llIie5gh2L7nP0iPZBr0/yb7fGLLSkzhNQKisyp4d+ZrII4PCJ9UBpiQZmCn40BsrdsZRE+/
vDj0BJ6+S2eKUhr13CWwE/31wvmhVnjj+eDwjjw3iVSDf98RAgKWCv2l6R35PjnSZ4UPtjWiYXpC
uhXjgYn8Z9fC37dNQfn0+vMvVG3Dayrh6AXSZU2GzxO5Zs1J9wpF5xQdmP5UCzM1KD9fj8IT6gKN
MHcjw6z8pi6NEPCzTzqriasEu/gzcPgqpep2F5usXM2D6g7DhY6UE3gmUW4nn3P8wc5bVzaaHWdt
xt5IbyPg075xlmgiJ6xG2wLzz5thpA1o9qdYGH4acdl6s+/7viIutJrJdNJrx6kt2GF8rGQSFuEa
9IAFKmtWNMLpahO3aijaOtdem5XcxsWbzzJV6qYyqPcPDHHjiOn2KuOA/n7rEFKnAZOD5lwn8lPX
wzVdC0Dd3ltpLiovMkGkXxGAAT2YxLAnavlJaaKtYWuZndw77kG2qELvZiHv2RcmuaHDPLItWAq0
sxIEc8Zya8VOBdTcgAAGxrqcwd/7vL2N1FerTVmzjJgqqn6fObKcNJRX73x+oDAXOtPPZjp04EBk
vrrX0Yt5+cn/D26GWquncLCHPxSERpTWwR7DadDYX6fLflpFbALo7C6Un+jonYHc6nHIUm/0i90f
VKhIWb/wjFs21wCcz7K6G1yXRvsfmKgUj0ye3k/244TfJLBeBvYnr6GP/BVkXkCTOkyus/GGxLsj
FVEtCokwXqagPRMr8Hp5OkQxo+H1yKLfy3AeaKrLGeKcA1+8s1ZhtHx30r4mx2/FeH55/8EzYAaL
0KmdwMo0RilH/1sQ07o2pzawVC+3uGLZh6sqwuKrZ/pxGJwExoKoIuIWTT//WxNVxx1tOJEtsWME
gxtVoBRWylAowszYLywkk8M/F1jmZ+BSmMMxJLC7YNYVa5S0LnBTlYyU1XJmwwLUEU969ehBSz3X
ZbojGTaH+5yY/1nFSPn8Wu5jq9HBp3Dp0iKmk73ugeyy3rIy02OYp27fvEzyuMmPhN7IMsE1dPrD
D5jmvMkJX07j7DW666oLOa2Tthm5E7rPMjeDMl/+29ftilmxlcKzVoPl2caOXpp18gYgIBCdKN/o
XLvCQZpZxLav2i9dwZJ5+bqOTPEE0+uB+4SA/4v7y+8win4eruo6V/0a+kzNy036RTcA1sV+Ocy1
G/KoOXqDl5HUDZHNcNjItYnTcGAr/JQzCRAyfYiT//nN1fKxmoJzSwfqTUej4Oa8v1XTwj/ZVnmE
5AWIcV1QGA1P9RrfgCbh0zOpLhf8qnZqDVS+JMNiFQDDy69LYwuYYc8aHbHbJj8/lld5qNprSfwr
1Xo93ZlzsUURbopvZNgyy/ygVslPI4RC7RPE5Tgjn2ECfaiWf4IS0Kyo7cZK4WGjVGF+D+ik8zvZ
qk8N1jlMKr3KkeIih1Zp9IDRHiV3BoA78BkpMvysHhK5a/WK+7HVgWUkZMi6eVDXVY5lkXrVPI6A
Kh7rIgy0RfrkPm9z4YHqX7dD6DCBHI6vWEr9QknLjv0GpnWI1pq0YVBPUwtZrCskOfygMHvkrgf7
WOJPf+i5Ka40gaSxhf6XRnjWz7dXFwZN0nGg6kBu5UgQd994Cre99pGpEFj+FfMnnCu8R8tVjRbc
f2Bi3DSvNu2xuDQi/XtfwZRgk08QVyxZYrYTSs2n1BeT9m+hMMaXozegxQleOdIBZlW8MuDQMBYD
iplTkeJxC8Vd0xc/AfEPiO97KmdbxQHsHDmiT+wmGWyVcG6YBlL1lmyUcoUEDtdCJdPdN+qhUddL
wSJaW8jVOj4xnkUALTe75K5ZXM95u5MULgxM9DEG5KDI2slMw8g7Niqit5KQ7Wkpcceeas5XiM6J
9kUh3b1nmqoe0Ik/CUpzZSyfQcozbKQ8F9BG1wpKV1XTUp1AXrQCBQcrZnzUENLLythkbyzHHZck
B3Qe7OZ5PGg1v3rg6Uxwf8/cfTbDJ9vGG8jxHj4ScMYv/vcMaDw48fBYqHHtU6rngv3BxXlolQfB
dqHi32CEZlHJe7egwqo72yEcoyXT5Pm/qqAHapeqQ8XxyC4poZFdCQGqVhXjXxv0kBfPrMA2qCuT
1h4TDaV26L34mjfdspjlyCHdqcGBgkQilU8NZ4CBuoDO9YChh/LVtVvvrJo7aorR1kX4np6kHz0v
zuyb3gR8uoNdiCX5mncS4EI/U01YmQsqOWK+xU/Q6CAUGbm2ojoFtPJeOxTj/iLkpMPgE9MxpFIJ
jRt3ANWaL5y8ae7q2+L+8zsqJlkx4FpUNjk3sCCVl+iTahGt94AWfL5rSDfk0m2pa4RxjLOztohm
uTESir5sL2ngHnhj8DKNyHXhak4/lqw34O3oFwUzoJWZQjFevA3d9m9Sqg5egSKRDGjl7peWxrSx
ubkd236SS7kZkIw9SeGaGZqrJj35+xxOe3rE8tzXYu0ZkyDfIUcgFNgZRhVnNLwIrToM0UM7zsXU
jxf7mXcDD0drMoFm3LUz70lKeGQzBQTispbJQM0oZGiBc+f4US7gToJQ6RoQHps9Zalf+daUVlbR
dHPCc/5ocm0AF1bYSuLWuISTNlG6TJTdmX3c5CwITyLzEUAEt+5kQ+sLnfPTQTUWUREXu1fSqTeo
tYQWKPpAnEMdo5vHWtQ+cVoRB6w/ep55D093O9fjTh31pEoMCeLAGKhRHhHFiZQgFn1faPyyjA+c
ohssGRx/dv/tzdXhf9e4/R6F0mwWHqavt0xEvgQRtmgN6u0Q4YzZ39vXWp+C+za9siwYZssIKl1w
m2F3t7yL1M8hvvLDhXN0DEghRuFmehYyaqBtcHZCh7tTvTfzbQz3Oc/QE34bhBRe4o8DA1SYUf/w
i+YIOSLzYtE2DnWl11bDkzlYOcFMw6CX3Wia0HY5c8oV0bi4ZxNtDiR/WiKi51qc44OziC5dq7um
EkrKMYpmam5oTERm7X/JtFPgwOEyXt50mVYEhCG+41HFr54zoGlN5BKFjS/lXH3EpeyCeF81fBud
2XWWoBvHSP0uQXFj2O0WN0O2bwUUdHePL+FkgEG3DfQm/7lNa91u9DPYDzC231N1vA64Eg6NF/QQ
B2vUTdtngoq/KOGrT0We7DDiVb8omeEYCMz8Ka93sk5GNi1IvtryaxjqyD5pjFS0V/Oel7l70aTE
EAeLzKox0JS5kGNUdo5beikgZBv4+4bCZh0KzS3QaQ7jE9CmUyQTcspU9JLTuJ+j8yRsO9ZhUvVb
EgQ0BDcq0SWsC6EiNz6kDYr/YtStp5/6rqo8KGnBb1+et9Z7h8LqoH6Oxm8DUZTB33qbgMxn/NdZ
d8hAuGiN6BLW3vVQBOwf38lvnzgIrefdVt2eKm2brabihDZ8Ptn9FlpGoBFSWhPT7KthZgqyi6Cf
UfS1xY0i58jTBFl4nBWpQ9lRik2aEcPmInofw7d1c2Pak5AnO+15gpSYKAGkpm6Kkd9aJxGb5bZK
JX9V3AnQc2cdITpld50XTHqu/LGBZmpJuhKtD6gJPN+/mjfwJ4xa2fun/MmNq5821UY/TItoLOsZ
fmnVbRGe70Y9sH+4p++seuDIk+qXYxst6+O67YsGgasvL54X+qPwX95girxleUNpr8xtJ6Dh21HZ
RsEfTGdOlQR6sPr6JzNIBRbhSQ5Vs6H5BUQlQJ7EDLQtl9Vir3xfG3GxR3w82pkTKF6v6orRK8nn
0dhiM/PfcTQxqWa0eav/I/WIGHcXd2nF69pFa6G2pEZt8idx1tFulCI+xOYPTk9suN8OYNjJsEPk
1CS6dTLV2Tu9DFgX/Qn5sPgiU6BqFKtEk+XTvX7OOfBFZtclqEDfo0oeIkQPZpBJCWsBATf0q6AT
gqHIYjd6k+zihpJQjkafe6piHqc1O2wxu8bLUOw/CTAqByTOnNfkpzKkXB39IFp6qW6EWLjXYJYA
50F0JvJTtyg9aFVLMrLvwSgQ3seQ7QfGAWqR+kv540K+aZ+F/QNxHx7lxZunE6oUVaEj11J8iuIi
73O9tU8vAiDXc9evvgCXqRd9LBRy0QQYX7ubOyOfZV0JsJJ1iL9qVoS8kPdIEIgSJrXRo3pKRQ1N
ey4iDA2En7PgojhMRVuVSO0pevX7hCjTaVKUgebQzOmrf3E2KwObCJ194EbuklQnr0XSU3KfsItj
S0isTXSAw1RA8LC1uK6ZSIxUsfITCKbzTK3JRJTvtqTV/DNgoi15XaTaBLZ4NiJT+MmQt58Oxk4+
jktS3KOnleQd+gWrIH7oywuI9bDJTbhi24QWgwV8P0S/IK0jzu8FF4AlFG99Nv0sKNNKzEm72mME
cZb8iaPX2+Oj3HIv8j8zLAwSS9/EEPknbEHKBoFiIumMAG6hGM9OJZwQafxLxzkRV0VpmtPKWRpr
dv+fXWrLfNuoyQEBLjlp7wAKkfZ9twOHoIbufSsG8MWlfjZFrD/b/G9XmkQEL6OnHFQEHXOUIVHQ
sNIGaYH/U5EyUAh79nnXN+B0Hcdgd7vQDuWHtpGrovK60MVNnX4a7aNUNtqPqdKKEU4R7IozP4RX
qHKQz0hScx0LtavhEODC55QT8NfjE3b8Opd2WGBmG8hZEFftk90iheexdrPPSVKAFu8XyvuPr9BF
eE7z4CjGZL/+X1iO0HjWKMZnNFy5qZnUufzNSBctKqbSIuJKmYqzgeAn7zuKqbYLOrdyErZI/LA3
GU2yOBP5znNDe1yApg87PMDtdYA206xFX+UAp5uFlqQhhGhNywsv2etBgbEM95tKhPOqsVlFjezq
bXQ0eklgYBf02HLMdE5zJARSE9q1BsKzMkrO/e/t9TNBouiV5TPQWm+zo/tz+wAQB1hYrzH4d/sS
OD/IJrdHpjBQ7utYtjuiVNbvr9sWfUlxiUB1/xzDrcMpvROruIWfzYb7SsGw8q4vn05JKwHEaKMt
xwhesqSCe8u6r0j4wl/9+Co19J/RWK7XYVEfDS1H/mwphVzsnFVIYBd8ZcWpP58Qyw0yoNPaxvis
P+mxVbKjEASgac49L6E+IvyIA2j7BQTXp3INkg+pfOcUvQjj9o5iz1uohbvAECjy5yxAJtaKx/7N
QGdFQxqvD9BJXU4ISPyrV7Mu0xwNyDyfGZk1KsTfAiSE/HLYgZl+ezlMxYDU2PU3sNZIo9GmWA6l
bv3uoMiJ9iqSZR3GN/pYG9P0JU2dGX+w16ATL0c6lwdY96KGT64HOT1zkwi+uqu2dZYqIhfkDomS
kL9ah15zjCWpXGBK0RDaryKn4e4RQ9hgDa8jF/V4rKYKQaGOuC16Jx0kOSEuLHJB3XayCyRWepig
iaqwUnui9VEzCBoUrs0r4Iv8HFwBJQ6Q3d+EZANUoDaaM7Qr8tG0lpvCohHQxQmlv0TlszSDAZGY
SP3Gk8FcBQ6jHiQXIyPN6x/JO57unYNUjCgHeuhUGEeNpOZk2zha+oWwndTqjtcY5WfLLCgt1+jF
0jxkUvFmCBh78FbdG7MbOjdffk3G/wjFYhL0zHZlRJHkjVsNC5aMInao4Wf+85L8N4HYK7rY6uSX
COUxg3Lz3PVv96gbAy4PzsKZmt+FIAWKaWp7QcV3sc7Wm/H5SY/Gqhqkbea3/dRoYNzG7mykZJ2O
UWBTPcsrD+fP8vZvQfCbLXaNW+YxnGJzaNANFxfuXq0w4A/vbi3fDJ1jFPsvkzJJvg+xZZJ5WANn
1Vbhvr5y9z7s7JD0wNFZ2Z0dMhG+xJU856OahO1yTA52OAPs3i853iQ9OTSHRc9BFkD+RQWNzFUi
FPw40VfrF5AmrzQh9ZK4M+KO4J6HlKwyuPbFIsxREfJznoiPl5zLs+srKX/dij0Rz/stFACbZFlY
k+wPSiKz9zJlVNwt+fO6GqbYjbn4A3JfhrqqMhc++cx5Ak3edgWYGudoYr7/u74rxb1YRI7x8UVL
JeLoFSxxtU822JeCbsRjzYIYTiXiqMdlpyag4gEdYJTW1vW33+AVYn1yjQRWLydKjCTDWb+4U6uV
rU9Poeb7tuNFSOhzDH4MHdAfHp2wqo3+ENXSdc0BJ3ef7EHNcLGXatTn8bkTmw4/AeaMAW4mQ2Bq
QZD+uLR3g7iDuw44etQ2VUe9SA0OCw0pyVr5lqu/W/t3Hv4KdeO0PM63IK/10y148Uw1pEiaZrG5
wDX67r+dkg/wquzUkk9NAswtp3rM9MFH+M2uaE8toTGlQI0jHDghOFQMW4G18/gwGIeC7TJMT5k3
W6hCeR/9fsmMA03nK1sxoDCH3sUUd4IvsrBPln0zMiRI6UfzxTn1hqOALRELFaADM86pVBCD7a0G
iIc3BpbycM2EtlD6m8k45r+g5s240udRnZ2KZoqAU0BPLw1xqfnA7cXI2sR7BSO+hgg0WJeL5FcM
gXwq7N+2c7V2o9Bn/XJZLVb0E5Ewx3Y8hxfYIG/fWeEjRSpcrQLDvzqOpZq+UplK3cm/pLxdRpff
VWz0cAYfX9ui/XBSQQhFSp2+bS9Dh+R0qdDEuJlAc0NWZKEkjjiXH2SzPNnpcuKZq31ZkUvGyp4i
swT+iZOVuIfYQUALFpBsqR/ogB7dVEexgMJ9idB8s1ICG4exUq9tMNqSfVSPGUnoYfkdGj7mxhUP
G94u5mxFd1CAfYTfR06mXxd5Vl/CYLmNbUzYOZOtw7nd+KivxVWb9Jq4hgjuhQw+QXR/1Vn1KzFH
ipuiDd2a3zuhJami035n4N0Fey/yjzDkqb6df01B04SVx3NxtCHBlA2DQF5OlRqxnZ+r3cWUgZvk
OkXDdhJG0eJLshflgSICxHEnahA0ZIyda0bcf8qzzGjhdUuE2xAXw2R4+SCCFn83fZZ/qZP+sadS
vj1KjVQh2b2b+ttRzeVemhAktSxef2bj7W+EInQSm+2G3T49H7fpqSK3n+biW82M9nqmPNZ6w9Ob
T2L13MhYsaB3YA3Ay49ok/o9L6sf7BuT6wA1qLrTonicLNr20z16xNE8AzJWNGBsb5Sy0xGjxyCI
uu+9hGH27f9hghlfjLAddZpGwmP7jT4r3QQvKpaVLFpAvReJ+jnNO2Q0A6RyCaqE3TlAyaAu7E73
rwguKV1NRSttJ20XL6HLH3vcWg/ChW0loKn+xk6ig/mdXdbHsJ4OhVW9E2pqg6g4aHzWxjzYe3wQ
PuHdsMTxtg1Z0J3sCAiYH+k7rAUD7qAdyOvo/+0arSBwfmGIJZfCMFY9sL44tTuZtT1i1eoJ8HmE
EV79FCCzsogg5puVb1R9D3Gs0dlUWUhCgyiOzRiS1ztTCWuJHcfbuGnpJoibYuhWkzvHsCXptNNb
fNpK/p4O7ccwMbco1WX88Oge/36N2BsZDf/ekz9rqSfLp042LeU/84g89FBI88krR/CE2YNWeAan
vSG9U86AtpN16MzYLNAWxalPikk49gWFfQ4Uf4GgIbYwXBSXh69SraUuaeUph0O4i7C2Q8MLp6yK
/ZC39XGp11dUpcmp3a+GmYWUUbzvqBJgGV6OsK4bdm7XpCxfnskVRRF0WlmotchCwIlbuSpf7qDl
T7sy/Tue4faYEC7dg02LhQ77ZT5IE1RfjcK//79BNlIkqoUj0y5S8+36ejE0yxGb8Iac+RsqlU4G
GNBUEztDVKU0qmh4d6cIk0JghIBUfFygpi98eohcsOtm9DCG4aU4MyCgR0AgwKySSWtHoaFZCGFn
yXWAbDXWUDCFckXvIeGYpFm5LoWCn5srLhVzC0TKCfpTjjoVOziH0lk9kF/I02lzo9ppuCyRiO6O
wX1qzKmWK8UHymmD5QofvMHmdghjsOv0hL7V8e41/EWYACBbhsOH+wSaqsa0Gq+VQZ12bHNaR5Br
JcmfQjRaQX7ECbnTUgHhOL92Znt9gbMoAcwHi8fjaxPr+a68uEmoAv/7f2+nHZSZ2irTGpe3oI6+
Ay1kaxE6nqZbcBEWHEo+FqY3G1tWMnFYz60sWTJCLcWvgfLplL67jDy74MWO/iz0qEcpiUbT3gqn
nhd0fJDJXgJ4ag11oUa8leW5b0CywFvmX7IV5PHWdUWckzOq3a/I7CCvKFxX8swFFZ8d21y8fMZl
m491D6MjiDPzTc7a3TWJ99KaUrMD8CvWE7gePHbld/eqWafXtYh/RMNdIbXkIWPn7me4xKzdEA+j
d6ENs+9u6vwfg4K9u5EPhvdTeF/+0E9FiLmQhaBTDYyFOJkHbQWCVHOqAECI1BkxWqAQEBG9fGdz
jSYpChAwSXZhYTCS0Z7/RDu41MuG4671xmxA3G7A9XCclHWeFQLhASWEwQNDGvlm/OSDMs5CoRnl
ObZ9J7usi3kmW9KvqSIKDLLEzJnHW4lSbZ3U/6EVFzE+3izt3QmenlvHRyBdEXCuXGZjl63cvr+X
KsIYHbCQuspLLQkxCW+9fo5AS01NepwBmDgcgFUrLq1x5/QEo+AxZ66qr/XLO4O17M7mFh8d4Ou+
vtvjz/7/ZgRiWci83uK9eEULlYZ3VGmp+fLkwt7Q/eE/WeK14bBtxSYVzumRguwBMzZmaDSdTOm/
+FNBckOjELZ7dYeo07M30jB3sqVF1xHAG7QMUVkAHA5IAN+3UiJWEZZpuDp+gtzaSCxmfFDp+eic
cwvhNHTpEGyHmkY2MRZ8Pysbgvpv7BpO35KO4p+hQQyNkSqcJVCzu/HJcJY/paM2sNtfIxJolOWz
ZPOesvl/eE5d8WDSxG1hYZLEtS6sdAe9QJU6EvrzcxHqkgk0hTWXabBmgxSZTChQsAIIZMRhQe2T
2K3TmP0U2Uu7PzdzBOMUIpORyOuhQa3pElpLGv9UHk+HuI3TqROOroJ4vfdwWuJUaBRt+tjI38Ym
e0mN/Gu63E7Hk1bNVnuaFIZB0V8MJGDAXFBr1PFxd+1VfKetvtOmMyg3zfNhNMktSwGxtEb5PH0K
PLQlY6kNQldAwlOYECp9SsMxpHbSNoZFp4vAk8mVxkBaNrDzKLDanUE7qRp++s+8nOtqg5nyESVi
Wol0PYOZQtaXkUTzCreGYtEmh0ipT3lT2cTEtrankIPuuJZXekjK0+qUZKAsExxnCBxlpCB7B2kW
S/oXnkz8yljZFEvhyQcf8aXkAfTAc3bh/QKaP1eF2RIX7i/c3GfMl3R+sFVO4uv9v2Q5+mY8//65
086OdkRk8OVOvC98G2jrzDv0sEN1sG4yf/eUzQXC4bp6rHvuz8hsHjnuClQTMZcSyIwB1gsZf5zS
SsNg45hFpxO/MSVnuowiauH0YzqcrsaidAW6RjHLD5L8HdBD7xZ87vjS2bpWwoZeJzRn9E1I8kXp
F6mXSLi7B7BPiL4WXKsiRQ20eQdV7Dj/Yz44eJOEsSKQShsimaWM9k7gBZBsN0cZM/hNAqsLPE9t
i/1jx8x3QZVqAr+BJL/PV1qo2FimVDiqIYNSrN/qhNUE9f6iHLAVJNdND0NoJdHv5S2C4WmTIn7X
njvOTm4HOQWs6VO4O4tdljCp0QaN2v8L+fzhgaHwi9rnmbbZUWFdAW8LtMj3vXFooqu7jeqf0vbQ
ljC8H0mfnVDiUE29Rdw1fVcil5/X/YV+ZGbAHy2rnhFcVKOaJo7oxlxUyJl+k0eJ33evS/YoocQg
Jfp373Al46HY6aVI5mDO6U1Au6kMC4ZF4sPcCGHUVTbuAScoB0AXE0bc2/WF9PbTaTeOKMCf+uOn
yd0DUDklHhewNbh1UMAILBy7K8ty7iA9J/mWxySpUYdtLTIUUnARm5gvciIlihaF/HwtP5LaC+6r
nuZoLEIiu8jxGSsE9q/FZwLqdErQrLF55dIz1lbxfECh5ecbOO+lXUeWsF9STT6agSZDkefUGfRk
/f0itFc97X2VEO2ADHNKumUz/N5wrDi832xCm7X9O0wP53OMd9j3A4alcSRlbZovjTZCdyl+4kGm
dbo+QrSWz6ssRaOKxDuj8iLQyOe6se1ZQ7NYMUDIiy4hZ0zQsuHbyZJRT1AEEe5zgKIXeiOwnykD
ULKJtB27mRyagT3AqNc4NKnmeCmEAcdMDPRB1U9MOuwB2yWU1tfeJNJH2e63uptaYFj5ResNjc0e
Y6aCIyZh3w16ams6UMyJP7PJ8YrafrdXPlSLFg1GcwiAop3f1uwNYJJ7eGmQx7xkHb2ZYQnvRjXq
w18rC+iapf6DTohaQXwGbl6ci/EdCc1K5A5jWb0d7eyndr9Dpa+TG/ap+Px/Qtgxzn71EJuDf6Ys
b0zaCLtUXfzQcd6ib+OcdauUc4IDo1grbBo0nnTWQ5HCaoQ40Q9pb1Ah9Ko9m5PTc6AiX5/wnHf4
cQ4ccSfYRIoKLKcZEo6ZvBiwLkZ6wH4Ya5dMAwZ3Y6MThxSran0l4hkkaWiAnlbY0EVftbyagojo
LWI0mHwW/mJSg33sgqDt3BItAKpyAkZe4P8yoAx4Q0uQet/8JWozpWp/kAJOw+fknIxnN/f7D6Cz
G+DwKSt0p8vJB0bS9z5TONv2qtkOBrNK8NHOae+qAV3YiBwJR8Isp+wnz5GHaeUo1LHhgb8EBfvf
Vs2jgkMtEqlovHSAiXgiGtv7AjCJXH6nMduI9eUQXwSp3s5TYJftffJZEcA+KdvZ8GSAtUfgITyP
fqDzJqSQGOnGG2Dwc2q8d3KUJhNRMvioFHqhvIn3vnJw8rStdZ0/wQOMztnWgkKXNAjFikLcvWaU
74Eruizlwwe72G6g2pSi4oce6pmP+tj5otdygQnPTOHQLHYjxohe3WJluvh92i+AXpQbfV1TdCtr
KtEPvOaJqctCWLMFd8pnIy15yBNqF8hbAvOhLVzLWDggz1ttAGjv6y2f6QSDMag3xftAowlOAZtd
wXplwhUaR6wkRC41Q8NGeWBJZhtyikWOjv32VbffKd0txsFWZWCmyW+lwcmxIHLbsntAtR6+MjjF
fXDMTmBTdGZkv7bpPit9GZ/2MBs0BTik8SNfAdeCH3UtoDesgU18tWoqOZBjPSWgi1rHAHaSmOpR
2pTnsw8ydmbtzEFYKChrhk4vzayzrHHsaAiaT+fc6IW4cE8M7HiJ0Jc+MQavkROLmdbBNDI6E4ct
J2opigDlsjyHGBFdYX233EpPNMzn00TGInc4/stAWKGIAOIul8YlWJ0q7Hvp0N3fqyqNtrFt/cet
jTZeNGo3fhyEAku92J1Swy39QcvK/xfr8n1e7s0rUosil4Nyzb7SG6FB2A4FkuFu1N9p7KIm/XOL
acFxGc5MEeTtQ7p+yBLqE/6twMUmIXMQl5xDgPhQpVmbeijpzmgUmGN0JBISzWZUju+Qc8lp40Th
RyOAza5mlPOZi0Izt4HLmxObooH2W9YgeiicCsIgl33Qcy81djFvZYqMcI0ns87i2PCIEGz9WT+m
63xmk6KEIMGmm5CS+zo9+wD9weIBryO1L8UKIDZSGHQ/W1W4Pa0BDkz4SK1xbFP3bCAZU0KKr/0o
wIrxmvlHiopyKUEP+5kzdT9Ptrd0q3mh9p7jGMLiMnWwuD36AE12eNqu5oRCZ6pNkwJ7C6IFGuq5
phM65XIUBOjm9W85VkBPkKPwC1DCHIvSL6oZxFJpvLoaaPc68dWX931+AaC/MALTHuE0AelTYqWh
Dfux+TlAMqwzjO+VWM5qizRwTrTC/HHPnV6rocr6G6LYjMGLOPI7PORB/RqNK0sxsa55X/ubE+sP
QkJm/O9KeMM63SQQXSA0yIXBRqRo1dgWxoAUhnmFhXjubMcmat1VjSlUy63abY1vMBYqxDiHY67K
wA6AFbUlODZEEM2dCXQWPzfkEeZhyVsfi5Dqkt+3CK0H0lZx6+8XKZdXyQZ0yuvsb8ZTjSBHyc60
Yzvn6DcAsVSpgkNaMoLNqJ/fNTMTxSYXm9leshq0tSy5U3xRWQy++DA/i6M4AbcPmHi5nyMj17AH
ZF1S5Lp8sZCXjUE2bt9NvZd5OGdulBj0ZIhMY75G1L6hgdRtzNZ9ll4TrlcEjD2wU19TMaDn5x8y
wWOvY0M4ai8zXTF37J+99modcL33/QqiIF4VEKcXuRFC8cN2tmczq7v1bVe/XmDuIoD8j8jC81wV
I/kydNVhQxRP9lkzF6rJDm+qBIuyy95veLIN/vBYLez1YgJ4o9/kVud8QgGv1itCidRTzm7uETuF
Lic6cTM9JSQH084Iht9/u1DJPmVdhFZc+RGdHnNoSBzK/A1P7F37FnSuKOXMwZXGHJQIRKXVP6cp
Ga4gwAXrZp/dxgQuggePjmDqh0+BamUchtJ9Y0gSe3nkg4jAmi1TVpuKVzI4H5BRyWIAHym8X4C0
S7PgVFFglxlZ8DMqv705+4SFGzjAFec818Y3MmyAvX6XozlKur4N+ZQXes8zI3wGmbcR0YIhD89f
NamDhyqg0d0aNWDQVJ6GxK5SqRJ0f1TbcoeFpkdXXJk3MUj5/HL+OVB4GtmXwoEtwrpGAyl+tPok
ETDzgJGv22antx3ABnutO/VFMP7K0T3mtUEPf6W2fNBZ38XJQKBpw0XZ+Vskf/8Aab7Yc36HO3o8
Rc+4k9/swEm0HauBoyGHtgDBepnjj7OxEdRyhLeswwi7oN3aGGz6boVTTKdYLx4zrYqsCyS+ri/Z
WV5ce0XDdVahT8RQRwGr+iZpOJYRQyB/KIiiJLn64nua3AP+NAeg7e/El5mOEGdk2pWCYc8/ROf/
Mw/9f9jwWVDwK2D4/hJ3gc0Na7ChIue5RFUTS4YqSzAmVeg0n+8mtDPmjl/6oEPPdGxsJWaEve2z
hdCEe0svgAGh53/YGBIMHGqg+9OLdh3iY4/2goD4kdT4wsJlxEXQMv4iGtNNAD1VNVVt9mWBGFwN
q6X2lciXToVq9PtcbeIhkItOWSBNUMVmNa0B8GqLf8HOMwOl+IyfbAr6Suv2SbXk69AkZD8dOCeK
1UK0amuQqPgnIJGNBw+dRmLLq95T5iknSxBrBomtwr121lQpm9AB7674uZ2kUWDpcf+T9d5WaAmV
j5ADDbjeIvHtsZyhjJCItB09iEtFP2pXEUPHixGkUfCWjtgaEY6X5FOrqw7Vlk2OYs1Gs+IoiXJ9
/yOtt+YH3prEn2vYeI9mMhfHRVj3ZomvStrcgoEhIhQ4sSrJoKLnGQZoSHbQXepyF3UrfihlnheL
zHrNDK4+M3Cv3VTDGLgvhIFMgRW9G2D0HuT2clT4b6btnkOsIMXRIfTIuLXQWtCJC2MjsXpAqFlP
E6uozxcze72YL8AO7lgK0KZaQV2y4TEyhY4WhN+fYPu58TYdrZ1lms0sCpvxwFYEtO4MEyu/H/5Y
beMotR9zy5OCU2SI0XkmW6SBTlOFVyKMRHoVK2WhMB29PiZSj6kdomi9l54WbpAdLXk+Hk/9vERQ
5ia/kpIWWymGgftmCFbp3M4+r1TG62Y63iFzH6VVCPFgmFq6OSB3wSF5qNvAGu45IZjrQcjCqpgR
QGXJITVWjUx19U8JLBj6YrYA16bpK/zfJolYfRfjaywyhBdXQLP9H3VHm4bhmqxLRBbfxTwt3KAi
i7RQgB2X77F6EnmigTGpJjcmIG6OU0yEnkHFZm2TOqS6d1ynaQHbBOr9HTZoV+vGA4o+ijDxkXGi
rJGAPpCkOTDJIoyzog4dTCaNg3wYX8cgUlfAqh10vqQe0bwp0IoF/8qxudPELieUwiFh7wOYSbeq
4mCs0mAj/AaBWZpwl+Wdqk78Rbbe8HuIp5uvCbVRQGYECNonqinxLylh4Q/OHKcIOW8BD293gCKC
D/MSgeiJDYfLCdwAW03cPhSBSbF2ltOLzUrqOpWyICDvBRPMOgEA22U5btr+zrzgVpIQ+4C6UR3Z
xzk7DJfukqXw+ieQtB3p6jULgVzsiMaOsLFITSC86QFnqihKijcSyThDpHhkKwmk8u1riGr9yt/6
Q1SvzS775zkHlIphTl00SxTr6oLTDc0rgwQVCZ4RHaUN5OIRWxHb6qlE42q/X9U3eR1FiVVyD4co
erzeLaAOQgIQf0U2n1zHrOuL+5wYK9Rc+y932q4/uJUpkaAe4soN9hjMwnXGyp2NgPXXY/4tvVD5
RNw+tt3izfJcwxCm7RKhSdHahltskLL9xM7moyp9yM1k9ld4Dnhl4HxOUVHUhrqGv21PvQupLkTR
1fdt/4Zg7AMCExX0068R064eAwSjVkk36znnlzlsKBkgZQQN7kh85Ns+hs2CbzffW8ivtnFmDuaf
hcRnxO+mS9XJ4Rawo55KssGbU7eBuT0nn/FxjiROvwIv8j1wgAB7hhuhTlS7vCTfM46B+yCofdja
CvNRNWxUlti8vv9gfbMe2R5MA+1HJr+wQS4bQMbYpXzZfVRLz58OSkE63TkZJVXUqR8Sa/leYeDX
PLpwzThGSROv8HHAUTRiMft6oxLzk1P+TzlnePBVcq1MzXm22scOvBTeKN+ThnCNjg43CuRW1o4z
p+ET0YP4sJ0hHs5z7zwG3NGXwajOuWEAj12+o+YB7jxp1t1jpTZcIJpdRiNry+k8d8NtHPUCIwF4
n8DLqU957/cyq8+mfoLOqVowEqxxe5c26mTmKRIGFaEi0hkS3PksCRxFFY1oQAzf/k1g2DkmuRFj
uOtTNlsBckkU55vR6YZ6pdBjiIyuhcyme2ks3EuUH6UmnQFDfFyYxsG5iW9ps7dRLnoWqkQcgsrA
1T0LUp63JgoUhVSdry/yxo3mMtDB+oN2yFhhxlVLIwY1M2rFiQpuSK17G2cwRB0Sfv64Bwk2iqTO
FmQlKHIR8iys3DPU/8Ih81ig6bUkF1RCsooJippT+7hAYwPwIZg8ESpzA9xxqvkgIc8WuVBFXcs0
Gsgg5HFC2jguqaViN6CIbrunCI56C6vfKDtHKdJQMySWomDfah3EAKeDtpHxISNTKxxCWrTWrcs2
XCFCz8EDz4Z0Se8H/Vc2+I7qML8x82sRPOtDjPhCwbnPQb1/hvJbV3XLE1aYiPrrCiyNtJpcvlRK
IKtbehSfYbkCyLOn40RLPp/BIgB4220HsyhTnOtNWC1eI9yi7+oRAFMrqUeMzTu8HV5vqOIPrI/P
p+kXyO3zbc/XdXO0NgFTGyMu/PB2vuuJdZDSPdyQfxVAoyawU88vfNEH4yRLp2FkpGzyvAXauJdO
9rcOhensM49AMu+u9Dn18aeclitef+qF74Sp2WofVrYcGe8f2CQUcvgERLzrYPbeVz0CoojZPWLG
g2FXwnb/17o/fPetIsLlU74HeLWZXh6BdXuPSBvcgIdDPHX4MQd9vQjrk+nbjnmEb8DIwUglHIpd
rx2nSJSC5h47DyI11pIaabS4tMvocEdyC2yFwPNyq/SAe4tTxC48gIGTvkyhDj2Lbxv5anfnXbcE
JHzSbYErUT3tQ18Y2PtE9nXKrMGqkljHLaFlCu9W/jXEDuEurim8Xsn5sJzvmZBf3Ki0YJ9+a7f9
aazQXB0yea08VwaO+XAsp1YtFUUbE+lHBxQkUcdCrwUXmwMHL21d4/knCErqQlwXi4loit61AOWd
4VZK86ng9Av5MszuBUOaqiXyt4e4FOTPGnKXU42XtjI6GvPpBcKtbjYap2aToRshiiIwFy9krKEo
CF98wlGWOeM3QXAJZH1pHHCmEgaSBOkRRDR0OFG30bVuftL/GVH1gBk8W2Wtsq5U5Nq/Ly0c6F1K
Sw8PLLC0kfMtWxSTis/locgNQa2XWxHS5HVH604Xwzc7Z5cF9gI5/EvIXSd/oWllz446Yntl2QJz
itLaY7V+khbXZN4JDuQza/efFKgb+2+YpCInOivLTIB7MHVIMGy8FUduf5HHc5FGZGkVHRPzfWoj
yNQ4i/un3O8kgnC+WF2X3mnAQ06P+DtOu1Z3F/r8mqRgoHDXtScJDtViNwyxAqaNoaFCuGB2iSdj
5zMGkDO4vBrw5x10rZyWRKuLTF4GiFSN7kak2Bh/5WXvwlejYw8g50VhDMgB7R9TevgHQYEfQwQj
Efbm/DNWtv3PtFLyVeoQdRqEQG4qbECDlv/SMWMfq+nz9domWmdEIlSVswpE3Uiy3s5iV1dZFCn/
fqp0PXMpzTPTvWy81qPkVQIPg4PRypUknyoCdiYRVzmDar+i/fPA01dqwDYTOfDmVQAIQ2eBXYPd
XuX0gdTFeyaPtuKieKeHxGlizm43Lc4hOV9EpMLw1OM5XKi61rtPP3cf53bpaKIQFYYSR5sYVerT
xndh/MqsFv3dF5UNKvhfcP7M8WmF1gLRX9oBYDidpOrZRfyVK5CpSXj2H4koGxExCrC12hlb+P2s
tzlBMTS5STzOW2hAZpzI/D1pxc1sJUjneqEi1CxK0Uo3YxCOzjDFl7uB11yN6A8kIAxubHxaI8rO
d8lXy3nYU0Wfgj5KNum1hz4+4gb0LG709HycUb1NVsnfkCDkFAUPSjfR3WAv4F7vYQbiU/yA/b/z
hZ2esrM+aspwFx6SkUx795jsKMRmk9MunnKcegp+9MxVn/gBj31pjRLNaXszhvv21iDPG7fOQbGi
aY4JLGHkrgiw4VMkB0ZlO/r9YyEzyu1bYr1T331uPTfVYhs4iLehMXJgEmXpyiQuqzLWp/++BPgl
Zwq4fhQZCQfB4lKptdk3J8+ui1VgZK6GOm2Lu6vPsQFcd4MeAgdmX/ifIgsqZ56f22jp4FKNG9Ye
FsvD3B/EGFHKRGN0ZvDfOKiG5+NbYQC82IPgMuYvBek1GI4thelin/Hk30m8P9o91VoKvT/CpIq9
WdlTutbKKZ2jtKLx+a08iioZ4ERUjaZIdycCFwhF1qzFUdgn47hviqPiYPafqTulLGaW5EhL6qSc
xU1GmQZh2JvnWSNOIuTHo9OJeA/IdXNrsi2WZduDuxJfsus5pj5CL2zXJGH1V2+1cp1aKME5jGcP
V8dou7+ya8aGS/VuxL0f4rnh8lgtStlf6wHh+ARzrlgybNdJ0qCNRZFNm+ZFsA7ZLZHXIHJ/0J/l
VRmOkJnw9I6uSmMimbmuF6nLy1Y3dWkKBK3jbYh2klfEgXFcwUUr7Hjfd8aBGQHorici5Eswor0B
KgqloDOh+520AYDVBu3ucOz+ZdfVkjOY00RnK7W/LLXZ2pGNSx+wn+EVDt7/lTyixJMoUxvNlEFl
qO1NazKveKOj1EeUQQGJ9w+jj7JTmcjd7iJXrpDa3IAHsxTg01EdE6fpQQ9ap7++/B7q2KNSyfzU
0OXzuLj3nx3q3xTYIvE7JIz2lH1Yxc/DCnXhpIQcoY4yGYQfWL6k550TgCSknMARJ4z0FTXLAiQJ
kKwbvwquwFepCvf67fQizSJ5RYD/V3/XDvr/6wpRdzbIBjSgw8F7KwUmYdL98Pf6pT8MRByqYG27
gIDh5ezocPJg0xSAGFevOIONnmQ4rTOTduFc6bHkHSLdOW2RizPAcBRRCV6AvMA/cekriLzcarN0
g26ILGkrx4WFwaWswC+9TtaGChwXiH41hQb/zkUy1zfy/udEa7/Kk+n5ojqhdNPsatrTPGuya4du
29xApCWdTwV+Ty7ILguhcn+PxdOr8MOXy+iqAndFT+Qpiay+pHe6GvYZmQfNYw1KKAngMLV9ELpp
vRz9u8PPYDcQFuNB1kMbhhz35W86Vu4O/GOGBfcSveWIQRPohMa5KqflYVrTOlzGaKq3u8/lVzke
8HW95bieAz2vISW/rXhBn9dPyR1rZx37APf7Y1iGNMjL6pPXO6wzhcn4DWaN+zLTMsrgnTCvfJRB
bDkKXBCY+W8A7JC3X1aeJYa3nPZ99he7N1lfjwZUbwM8yKHBU1uQC/oYC3s9dN33O/b+FpCBSup1
4COj6joWtXWFTqMSy9cIMqgygfG2f8J5yfUwWPOJos2Eb4Gf9LzNQujCzRRxoazoI2HtGbnTdZ+7
w5XkK3T2RQW0psUfKrZmTdHNtZ/AYtw0bk9WilQ4xaGB5qLSwqPewzwpyv0A50wl2ehCKO8fH9pa
cm2CCVXVzrpUiNPHl1sHuDJGeMavjor+Z493cXeroTQ2XITcGox31e/1CPvVe0lJJrjNg8CHFZXt
ouAwOCMGEQf3iuds+mV+K8sHfUktwdqFq1ZM9W1Iqg9rz+1iP6BUQm9yVkb43a7TnfREVZaVWzem
FKQ1pZJe+lDAQwtrdfhQykeAfnadUrusHnGWIx4OiAW6Az47vnvzw0IfRWnOHjdeEJX4n2oOTwHM
+8qY5VV2WYpao65em/OYnglRbE68ANWcV4MWZG2hW+vLWYqe9mcshOUvcpceZjZDIJAUtKGIfXIF
ZeJATaqjhM/NBADwjBPtBvSZ1BonCyEHhSWyZ2RijKpubhnfhoS8BUmhtqyCEoXDkbeNml43qmb5
lqta+AxkxTJfedILDLWnjitZIkkVoGfaSRrqPNNy/3QI1IT8ZOybSmt7/AFSx0VDE1rCOHm6OmZX
j732qiYR6E7BQ2TbIAb6B7aVikL1rJAHLOj4sZB6qBsfljbnMioVnX0CnF2XG/2IA/nswLGZbG6t
zWJVGkr8DtAjN4Qwozm0W4hWGzXyMxdGx1kobrADFOpZgU9iK1BQnKuYBw1pyEPO8k8V8aUwLQRC
YTcWhueq4+80DT5J2qzhGqB1exE/Uz458MEbOM2cldVcDumP15KUzDHMYv0NS1NXX6Vizz0TTwCE
usdaMTsK1whx22dHPbN3kWbmTCnlXHKmShoxVymJZdyr6GrxbRVhPwoZq0Wa8jXTxqo6ENpxlHKg
OWAqAS2xDzVypJYRkiTBbDHhJNMKUEHk+84nLSxX/VF2d1huJwTkflQ0pTuL1Dgd8cpugPxFcTRy
ZdQfDIDe4bD/wYpJNyEzuDNqKvQnWJzFk1XkChRC744tP8ZyYukbdaHARFzKQ1MAZ2GwEAYwRhar
jU4poaKEEVXjzRvEVrSASbGtaQiKsCWtU5xfgE2Hm/jUQ0As/IEG43gtsPGuUQIXPcLPbBWG+ggK
2ty4eEbAKEq1/9Y2E0VW1PmsmiUGbPzYaMlnAmBj2vR32zW89fQQbLzGF1aRxTrRRJgP0vdIJWbJ
fEqF+sAB0S+e1RhMhsYAyaVukW8AVGRztsUgE34ogZHB38Eh8K1Amf2jXGEYd0oKUMM6KLPTwlA3
Cqc5BIyQa7UBSAbCxYqHlgyk2wBcHKB3XXOadg50IZh3Kifwh69wCqBHiA4KdtuoepW+Qf0ClZND
XG62kP20YkhWJFTNzlnLi8vdU1wkLpGY/nN0CrrhBfNIVGfkuW/P3BL+tLI9g5OHfAmji4htnwog
UWVuTsc0Yg15ILG18g4txpuNNjEH/0OyHGLTXJdLv6rJ9KZ/zaK+boT6VqR4Y5u5dHO++eCmtb4/
fzqGSBTbpAlK3uG8GCfWaPunebklriL3S0dlAaeBDj7FBlnZcKf1PXMcvNmOD9FneYud4vHu8gSS
C1V+DjSjxQ4iRpQoNd+cgap9q5TFQDwwjSePnc75EiFzKbiN9y2/ZYeGZYh6R+adv0oa61zb/zqi
6UMFcU2n7wbLNztDRalKXLX/4s332Yia5mi0p8QP777bIeUSLLiJ2VL9Z3MU3TDf/LhXE0GwP9IK
pUN/JfkDzYAfo0457hqRDIb2S8YKqAD/mdOlDnzNSxH/UmlmwP8sKwpGhhaNu3c0dGPv/WkYa9UT
35a1ilHt8kmIO2XKVy3IicPKXLfeH1CbQ6fkbevT0QDK1q++mOYUEY+Vz/tmmI8AG66eY27vaQIx
kTs8tO346bjyEgTbL0SCS+OehAE/mCq4hli0lerfTjgm3/2rnsojDFtGuKrxA3ag93Jh+ltgvD97
k8BEls2LtjeNutjz1LUK3m+uNdaI1usTAhiC0rTj0rP81wSy0dyCkK+iqsO1gE3kMz+XVjtcuFvo
6ea+05gOjJJw6pNbWdOjhcapU+FTQ9YFNtt/DqgjP1LfZNthdAsP5sbtMQFEuY91S62Up0Vx47/4
g6fG0W0wvrMS/1J68nLtqTw2EId10pw4TSKKW5iRMgOJoNhZXF4RFt4vDyss5KzCYGMPE6zJpIz6
NfhTn3Ioa9uWiP7dx1mfRg9ehkN38qLhSOJC0hqgB9VmmLmzelYq9fgZTl3pYekbaTyKJzFmA87m
uslchG2vKwv4caetvuR/ol9+EsPMW0fklHOPqf6pYW99rLUPJ736fe6FepHAbcD/SwYHQOOMo8IP
X58xhusoIvKPryILhLuR+A5G1AjYb8nZWLgfpyJiw7Av6YyPTmraR/8Pb2AAuBlWBpfN0Ecs1WUR
6F33a0afT34/HQCz9LI7miSHUzL5YD8XVTp/2VoG0zfo5bPatTSks7UDVNUXKiAtaaZEdCMCAqqL
PDAHeoKhJvBURYwThio5ynF5vPZntewxAo7SKQmRRM5LFXPjPrYphRXYD8fN5jGV3lPUrGzoixHK
+B75nllVf8lbKPOzgsyfhCWaz0JxfgVbBc+F+VadlbZLVABGBYcAZIFoFXW0fQ+K51NDNIqkcpgi
dVeeJ1GQZILLwWZAgMYTf+eF++l1QU7xgKNRO9NZD59gjnb4UZnHcpMMoQkrN7T+C+hs5v9EpfUs
fq81xM2kczxN36SzMRYJo5mkU/kb9y1lxGR5u0lQwUCV5HHDccqoRXYTETiK/WvLUj7+7YTWLw2H
09NCHWAHRwCegDsXN0UpEIFbGzZcNm6OFjbgJffwXZmopkR5/94dTJ1t0bp8soHZ7pTnQ2YEPek6
JS6d5+Vh29s+uThthTB5+0M+mrls0D1BHUAT4/lF8DRTLs6155cQi64cy3TIVpJfp630Tvt0ORcS
ZaFa+VNW2MnI0fZZMR1n5AwsE58ydQns6vJvj3D0VvLDlXgAgA+gilJSMacUiDcsypQkZWsP1lIQ
ZXrfvBPGBdS4XH24P7t4Mw29NmE37Ew9re2jGOAnT+qWhiVm3JEH5/sSBxqVO9DM2N3rOsR+v7J4
BHU97MERO0vp4qUoO6TkyJjrQw/RG9JH5w90olAvsp5oxtPNHGSieuNgZMoFdqXCXLXGNmDhEHOZ
SH8yzOgbEsiIHRfsOhZz7HaHX+ws0dT4XIL3R4lJltkdId66iunCCh3JDovwI8WwMr20jYwqM4LB
uwJsy+oPBLdrcEgJk40R4C8iRP8YHpEQalNquEK2904JZjqxcI0nTb8/4ky4latUy4CvKo1QySbE
w3zNGBgYp7B73lZq04keJM5AoaVcqiE/yz52zGu8JzBfPYAFSpMAfqm+smgfrVorAz/kHPa1BXJk
86X+kVCrTHHPCIOBtevCuAS6YYOF7Xiw1MRTiZfQ5deoYSCuA0EXl5V56C/OrLQZvQCNLarcoHw6
xACYT0sQ0NP0h8WGJfyCDQQaCXaboubKu4ucFP/+JuFjS24rs9EWl/8ZdxFWldue1zVmNj/bVYG0
80eQXGT4LCUnQKDJC1GMDEE2eaYifSjRSGNXZej2xhKZ9D14pepnSTaVLQDyuhvGfbPEaE/cbAlp
eXRq9dxIMQ8qJYmSclvL7hb8KWQBpf1hLO5pEMrkQf5mD/5PiWE8afEIAiNtU4ibzcemn6tmU35d
vXynhlsz0zKXxvw+qD5iXs604aTVShTfHm+ttdyVjoK9W5qSuMZoMeSKOHcbM+hwxC3FbZrMu2Dh
sdkZTdfc46w+v9INOCnJuGSZISP4bVQHZ0qqScF9eGpjs9Q0XkV3pH/BoPNpfae/ta2MtyiVah93
WqVM/i77FdUf+m3S6mdB4FHexd47cRR+GWsBnd9RCH+rH+OZsm/OpTb+S1gqynIN9Erz7F0Qduws
jx/v847c51BQPnsUzJfYxkIPQoni8T5tZRonBecvNXL1MhcFVEdV+gqmmCCw4WMQJY5pOeEfPWVa
uQzW851e8HIOh5hzRMpVtfj9ptdnFXmEA+lWZGDqn9OYQw3CVf0Pn9CLuZIkUGiBNDW1BpHDJkgx
/mBpSZXZb26RkM+0FK4sRUvWKKFGeSepIeqO/1oG4Ixrp1iyh2D2F4V2OGOeYTMLWxBB2kKiUTQx
GD1sgUrHCCTQyMBDUIV9BvynfZpyBmnZoVZUR5jcyCkWIvDHa3MA+FYWtNzUCGjEcqKYsBPKZMmA
a09C+ELUnXqNcF3sNzWCK4zyFkWuU0RrRkznIL4shwMhktBCwsVIRPirlQd850pPsK5NpZzZprUi
feUV/vgYBJT4yoQ/IbOKJwBWfa8EsInlFo1aEsE7pD/dGeoFk9TXz3xxADnzySJBsFqAKHFNBlxp
I3P+K+xAx4o6qy9vVzg0JFcUMtnHsOUBNc0uUrfvUsYfxXEel7jThJEzNIvzTSUeL+Zs//8Ing8p
Bx56Umc9Uyr/JLaRDz74f2jw9jOw+K0fLl3puqJf7VG5L2kLjR7HfKJ9zm9MyAg2cOovVsQgrE3a
A1GwONcui/UmdL7z48p1z7GT/TKpGGgsOKDCvFh2sjkRwdSYos7mmO5FF5l499ThI5ZX1CkC3xrX
2D7j+xkVL5qm8sSU2a/eNIa60D2XXqTFPJPDBCUBVx8bJNYaxg6QoiPDTSrV6NdBuIeGtd3KrXTL
pSapC76RYm6Y0RENK2ltjawcfavLvWq83iCOyOHdRnz2+Ki86he17b/Q7tuq32mqsKXUbB0UQ4iF
Yxf/6/2yH9EOekOBe+a2R/Vw6uUgImgNMh/lOfBRCBxaSW6y7Pg1+dEGB3rVrBNsz7nXNg2YYbQ2
XqSlBHhbvwH+7e4Fre3hdODdadZuS7JNnDo5w+cwEso5Jc7Ddco9/NsQocrye4oOEUe5PaqojtOw
o2vd5AG53ND81g394LuAHE8lWiGSaGefn8Jh6f0mHypQ/KwqW9xXBHfzT8w7TAQ5GCPzkHJNTd+K
b2k4UYkTGn8SIgRN/cN/ERffVSzTOD0LDTLEwHJv8hMlEIPsO4tKuBZCT2p3YZzj+aBnwi4JsCxQ
KJrUsCYwNEqqMOa5/YUB2UH6UcmsR2HujjMC6agPrYFt5luSAocamq4qkpaTjDFnH7u6Hu0dbiN4
6pCCO4XRufDWyJl7AMQjhDP6tDoJQ48rLyU1UAzl6MNgJcbbwoQOIgYES2JJTmdHWDC0nrzcoNxi
hjr4ZcjtLt2/LQnqyheJl/7LvhnbqU5U/ZeebqhRD/+RC6WrX9XxoA3c5eyrNANTyzLnafy95gMF
irXV4CrfD2EyRatg33JeD/BSHlXSbEVpXOMx0q4sE3sSciUT7NfsAPMxepaNyfT9kzTa3OTTtlsV
HkiHC5v/gw13WeAS9pTyMMU38exTa8lILO5V1USBQbnJ8dE6GXMVWywgar23j/JvoPX8QIZqlYQN
jpUkGzgOVVG7NgkZXbh5O2ZX+ixQd270+9VOA4DRkA0fTNSHFl0gQ4iNqCW/IPqU2J/jfkn9czhj
oUNV1OMyz8gVWHRlVx0oeEeNIRoqDMSUg3BF/4lY8yrztzosgRZoyxmCfYCII9KHyZEDGEUUsM/v
YyvJVR30Gsd9dc2olNav1Tk1wub/cvb4AEVRpU+2GQD9YT83HAAT566OpT17pzXy1t3N/hKWLqGc
hUo79yRCjAvoYTQyNE6zJyAdsFAEuP0Jpujc5sW1Lj7qsuENWQ/Ul1Qd5yQOgNsIA4bJAT121pjx
QWUTjLquq9FdFUdBFQcIb/8UY/1C0UKCbCxOUkuDYn754AOsLjIWq7Zx2D0rhecht1nRdpVNDlw+
ItTygAU7+cECmZ6aBqqOemTMPI1EXAtjSrcwKJOyPxPYeQF5hZ7e7a45hnQKGx37wJBF9SjcBEpW
yzgRunFOKATxUdLjHlIATKyQYT+vDbIuLHVbTuSh+D+4c0WWpNez8be14Q25FjFCsm/VaIwYAsgv
JHWW6UZ5aoFW8QC67fdAvk6W+jjtaZ4Fb6ctnJPa14KZQQZngQpcN9b5zqI7XfDMQxKEI1AXobN9
72UWICM+6Nd+U5l1LBKZApI+YCPk1YpmJCsIoo4FtBAtJ0xqZ6D8bBTiHKG7WdIhdqlUU5VFS1Y0
FDyMtKydr9lb0u+I881TX62q9/StHNa5pifqTfnOmbcU68eC7HHuh12uDQov57DojGbT3wbQ2XS4
vElrOt5lm0kVmxnd0yX92dJgBYYco9FpD0umqc+w2HCRBBWXMbfFtSlRfyDILJAg+l8bMkVf2PTA
zySWjPjspcLe6D8QEtzh6EvDRyfoZbcPe3sZ0Qsy/I1azFv3DN+87ANNQ1RMbnf3/JNz2YSwEcNe
mXRy+tIy1pC1d5IgTu12N2YAbmXaI20bk37626e9v2C8swgBoVm2hu0PGghcgYSZl0WRfw4kjEms
WdBW1yQhWih9Ylvv8kuhhap3uBLGyVotK3ZTY/f3gozjdkLj9bkTxtFjJwg8CIkSryP6pbTB6Nnd
PQ7SGGJdwIr1AnP459A/Icr/On3xIAksw0n1/DEQFifEJRD27KinqT+33qa1NJOQ51H8hYTPtNXh
QCmqqNwZgomlqrh4HsrJ296oxH17dRzLmR+390XGXAb8wtbHgACREFAXIgkdW/s32zzcAhVyVlGL
U/rLq3mI4dc6FRVPuITUfAPuRdiNGLCMGZR3lg+zGtrgXb+QVKPTBJVv4uXN8eXqSpLSv7DMZ+QR
Z5lngjMJdftqE0d8iNYFJwz/PRKqM3HU/zTcfsZuZ5KKosVVkGfpLFJkMi0zglFypS7SqOsDevgv
3b4igQ5YahsvNhNz9icsQpJP9cqGZ4e/CPi0L92JzQi6G92b5y3jw0iZ834/STNPVaf1lLZnh83Z
80s1dJ+b82uFKKrSeUgVttMOwuE0U7RqrvuJDGH4yIfT4cgiSjOSvXwBx6+xQg1aOWzjXdVDXDyu
KHQN34Xk0+aPffxTCrt9+VwUWyBzOB60q3QLJ2cZDzDb6dtqNyRO2GtOiG/+u4sdJw/kAtbnlzgi
4Kq5Mq0JcP9j1HpFFNytGZ+gFCSxx+ZqmLGidIm4s9cjm/rsLfR+cb7SwvIRzpYYlHbXyQDH2nd9
8+Zo3/J4dHLJKJjHaR/1EMFWFz2PfrhQwMDDLjXuYQHhU/i4YlYMXOPzfzCQIRr40bOkqcJt7JSq
N4o0OsXsTLb2t3N+LJET38AOOYMjnYygdlU7/HWyeXVVy/fFHuE6xpcbpgyoH898zwOoePuE4YAt
pPfZ1PVaCW3CHPot/Y2Aix4dstkAzERpUO35zXgnNsjcUX85xjNTqMmVSsSrWDdP+ow78HQaEfTm
jVBjs7UQ8Tx/VkCxaSFNzDrZPxH3xU4ZNq+LM9dKxFd4yHWcYxdCZkxBPMHZKYHGmZKbNcyfvSwL
3GzY1FjPxI5v/i0IlXry/4CneRkqLDlfl9JvxLnz169Mx6faXgZ7T7nvsaO3CbG68HgXBCMzn2Ad
/u0PXKuynAf6LTCi7J77WJiU+/tAOFcESrt8v2xQeG0eeEM90OETrvQU0XdLroNoxAkslSaU4l+y
9R3GpbiMgzUtCsq+6QaK++yE8hVlrksTB73MNDWVFd+fVjf26a+GfddzSdCvA8H/BbN0M++uNzXG
y9TapfCYE/xLYaN8jDMWnoS9GMLH+q2Y3d7LagHNaCQrC09KkJWADK4XAl6PPH4sh4ERkWONeTt0
+9N6qUGEMHU6R0h/Jt0jtdT/bKefvDRb0rfeZtNBwjQoiNh+Bh/BN/UzA2L5do4JIMWx0rZuLmgp
HN3b2nyFNmD8nute/rRggH4ODSKltAsfTzp16Ps7KH97RMszKum7nJeMaTS8fJqBGhoqkEZuyzmP
+GGwhJGkmAC31yUGpkUFX4tBV9kVlxO7EEb9ml0+aR1yiZkpVbH6YESXWsiqqJsiZlqymK6Dmeyy
U94vwEaACXnepMoIroONQxiUS/3QHbu7d1JN0b4cVZF8vmpKpocwK5t5MWjMWl6PGkjjRAzE5N/c
bLbiQYzKhLsBeUGRHqvwH9poZoG4qPTgwOWvLu3SUfWCxzAqljAdlHyv4f3JsS6vsnFrBFQ12K1S
ZZ0/c6JlnSioVKCaH8/yxvY5tTVDM3MWQfe/31rbjBbwx1Fgt8jDrMJYUhZiUioO8JQXuLFdT/08
tv/YYGcI7eVSFaoonJTSTweOpVqIyLWU3WMt8VcT7iZuji6Hb6JmnGL+0OsKzei7XwtuAuJN37se
5PPD+PTqWOoGiQGynIxop8r/K9xZAB1CAaSd+2tlLJjWgBQryH60HsABrxzh8d3ogm9WfS7LPC9+
kstMcBD04Y1yC1hsg5tIox3EbNILOkPqL9fW2Ep9grtUNhtt683To2E01JJR4YlNeSiXRac+IYX6
mhsMe4unqjEn6ml/9XGVwXMisR1Z9dEXWZHVQW9yq/khI0wInQdaE+sSqck/ECXEIkhNQoo4sDMH
HJE2e+FeSc3ooh78K6BshFAO39m90uJMMfh6FoRT4z5u3U4VvgHjga1pMvkwu1Sc4Kg3Us86zSDS
ZCzX6kWo3m88tDeb/RJNClC/6xPQNVnInhq8BjJQAxgYBGK6UIs+m/N6xmOotiHKR0fjOEZ4aFtz
6KVtGm4PNRnR14gLsqesU/+1AAi63ZSir1PeNPnaonJDEeZk8ja+b4pNZT1QWccItFUxROCBfhFI
x7yYEyAVilptqt9Gz6S5xwNVMEh9VTbyh3wcVTwcWn/n5dqd6rD7u7JW31J6OhPktz57tw5C5Vzc
7OP0/ozZG4QoYYaYFxFLb+o/A2A9bzkEWMFy3qJpJCs9HG7QgExiT6sk3yc20mEarB7Gh9EPph+r
3yUtRZ2gr1CJJqhmXJRsm0V3mh9+roM0WYjEMrMzEBdaoMJVuywNWfl2NLHzy/v0Q5XwowDhd7Di
sGeb28ITCqMc4VbhibZK6HsK/X3l3kmaU914ShiD7RbWRR3lewOdZJ4jP40psJa+cEFQOFcjk/Ti
jWXMCGBoxrJT1VYmzow/Vl/KyCwvXb11bgBeqEfcjWsyToczdnaHp8hRfiwq03QxJKUtGt6HVCkY
tJug7A9kN9RILdcOwYWnnplZjhNZAP+rJbC/X5FiIprQFL/Oa/I7G464hVOXvAeowmbIYUMR021g
F14kahDDe7J6iLRuyVLFI01ONS0iY9flNbqS52R7fl3jewdOlIySg2kSW0NTdTRwdvMmY4BxJPej
ucBkN9iM3vZ6Hq0fc0ux88G0jtkH2BvLRe8bIYmIlirdN5S6Jgn9d8rxkPx0ToIHU/1RN7GEcLb7
fL4pTSFpYigM9esNlNu3taj2Ufr9pzaq5fHWR/PKcDqjMLsr8Lfsb91bqzK0nHU98Yp3Z125GNdU
nxBb4Mu/H0MVrsDIi82KrmL2N7lQm7AX55qbyyrNjG9oZGU7La9SkFeBN0Mr/obpW0+NMjoqggtX
jG95Jku9UsSi3xpCyHqz1N7ciIxlTsJ/eSS0Yi78Sd9I5ebMQ9YpQMM42rn/L24f4TPwmMEuMjMW
Vtc5kBsEilL8jBLzgneqd1ib6l5GqihMLbLXeNb9UsClM8187oRjt9wLrHx7BqF75RA/OFvkpzGY
75IweBB6sRChLoG5kqhl8nFQSvFLvm04EVqvxMFaXBjKrcUpbHwuW8AXwbt+0RYI1Eb6qjRx92Su
ForGrjMOkomJ14ZxyVamqWHuemNF6sLtkhH+CIcY3fwSLFRIPBlCU+BeQUISb0LpYL8IW7LmWJZc
cJ8lP4ykx3CnPcAlaWKl7ShhfSdz7gmJYc36k9mRS4rkg3+NKkIBp3bUOKbM8/YNGAnv+43EiM3h
/VRw7PlBYG4aDFOKOOQr0KtDeigG0dUA+EVYQFMNIeC+rn6WNwa4EXPqYwisFDFKZTN/uN0lVc8J
FveDjzG2iq4bg2911B3WAGg+DKSAU2laLZoolTvCz0qkiJw3p01wDplm06dVGRNENgpM7EiPu6+v
Xiy8KVCKad4JcsYutymbxW+U2X3fco0eoWV4K9q4dzzjiC/5ED3rYjldP8hQN1aRrXmT2VxrMXTX
X5knY93Ygh381u6ayiXdLChiifulrqUVFe2dTtpxb1V+aVaZLD/G2q/oEbzHVPWHwXLCLbERoegI
AFTrq99Lz7gJy5XkNQ16aaCRhRIgtJdA0e/Ti2NCHwin+O2zXv3WVCkWiRtl6JXwQFDNG/J00dsJ
M7fEcIjpQl7RYOUPI/bGRXDcYzaKTQ+91dLS7yavWq5gNbQhBJzeUscXQRpLfgAq5s9WRi9g/Q01
bA4lRA7ctqdxqcs8BPxt1ZbA7idQP2O4rQV6UK28BgJHfwBrZAxH+qKNGCpKTM3X3xqJAjIDbRtZ
M8E6Q9GHzm9mJxSjUgEsmWE0+qiS+FZg2bFf4RLAZ5AghTAVEbV82cjCiZ3IEiz9L5XHQ28qoRG7
dyz4oHkHPETDcN1Wig+k+egGJoelZFnTjLVlF2ctGQRkx8DLP4IV16cvagxyYDg+ZW3jA8d9vvp/
uCiOdiqKGUpNcHz+fmx4xsovG6O/zF59hrX83TH6PzFkQyKlANo3x7M+jqU2s+/4Uo6ViykJfm7I
zc3ZaGmAPHfwMqEDATparAf2byV8yiqx5S1wN1eWdoy4pptVxI149cSBj+xUVINl6WvmxYYTc+uR
OLh6fSMHeQ7M/Og2cNsoPEYl1ACfFw7MZqi4hc2g6QhmdVRw5dLYhDoyklqns2uV+7Lpa+Zoq6NX
ZV+G/ZTJoYbVrOM8XMLvLC4gA9+rXihGoYuh7iTwl9Qvy9f8Ao6mRgZ4epdRi/RWahklVx6vCO4q
PU4i0P4MBtfdTpEFOqsvmf1VKrCEPJY/daZl4JUdEokfqX96+nu2jdRvSu8fpUn65Vjb/PMUtu6x
H4GwPeqv+t35pG8DfBj+G+AsqZh2egS8awH/F9e2kKF+7DfNtWuPltEMjNsjgRmxUPAyIQte9jlQ
/SOdZFizmLDoKja2nOUrhZd1yiduixEoMe48AfzPx02wYifgIuIkgromjeTOPAMNYEs/Hswi3cgG
Xc3w3wu1QOF7iKZ9risHnJQDxYkv1r9CdYRTcAiIrIQ/8DLN6RmZOS15zTouBLnitAePTlXbh+V4
nWtCmRBScCodWX+rYlDP9ezrNEOqxb/CHGyqSmbf/sOorlwR/EZrrS5M38y4BN3jhlEFBTKe5+iZ
RJyDfDIJwYYg0WLDCJIsINzO1JX8MJc5SNxIglc3+wfblbJxG4xOKhexqE4ATebZHVNAt17ywwVd
l3a4/R23Fs9SMz0OzoyC2WCfAC/rONLcou68pJuIy9UMgmfo5VOEabNDNGvTW62uy8U+FLLml5Bh
lI9+yfsCjM3MBAvfHusUktyU4PAIh4Y0L1YmfhTQYb17lMtwKvRJqdBNPs0aRoMdzIP7wsU3L5SI
3IoPW3bB5YxJ63lhF8gvxXO6aNty9sbDfmDuMbj3YrR1wcTDWqLvV/M+4lpBo7QugY2WBDm1eGlI
JDCGjABJjTtbDeOhts/7/j/1lSRiMD3vRX63Q6eoYkORxjcfaWZ96CUoCqeCwVX06nTONu8DgyIs
uy2CaWztWquJ8+rXGD/9a+zPM4e3nNtnKdr0NKFHwZLdGBfDa5Iz3m26FWe62qo8UJm8CL7sRkIz
6TUAj92FhfYp5SkFQh8xlnXqx5EufQo/OTs1ECKeS7rn1Gq9BXimll0dZV3RQDx0Sy3twnyCR/Mq
T5mfykeVWqjgXCsUhxfmgHMqau58Jh+92Fm8yAJ8EEnXxeNGu+XiSj2gouapiRwc58YUzGaiQyb7
VQnrKFkP+VPdpZianQNyXW2WGhFTlWgFIM6qt4uZP8zuyKLT3h+/oICbXu8OG/EWWhha8TGkMTij
1VIEYXwC97EmLTGnj/zHo/Y/+irjo9Wd9F4wMFX5xHifQ1sBYp0BrRNujax18AAcYD8KSkzz1d7o
l2aTlZkvSs+M5A6LNgzw5ognflQnieCo64nFcZTJHeeivhtvmK3F4qmZaSMr/RF2/voUI4tDve+b
DvWn0nddKtUfHsTCSjWGH4dGjaF7lNhrOB8kD1h7BCIe82t5jFTPVuIn6aHUaaC9BujHJWQtIcao
OrV/+8evY0gRUdiGEjhsNfIbMXSYLB0fqU8XjVQxRpAo3MV/gfLZZUH2STRMMgT6NGS08bTtK/BF
bHBkO87XQeFyD2fi9PPdLSJX4QqLVi7h1Sph4vFTzMrr7zB6essQqqp9Lj9Kvvxq7jDBu8/x/5JF
EOSBeTyeyINAGKObXTRB6FVS8frHQUKlrjiuHEqv/4VjtrhAKJyksbogWANbcWp8Hl+QrBoQuB97
eAm1J1zuSlElgJ25Y5XHnxAw3Eh1PS90421shZTYCgmp+vcB2sXQU0L4+iPlKQJbaT3SjkEPgJi8
gwsytXh5nev/5nx8BwZhUwpzyARVLhmnxgaD/v6n07Q/EMOJFhO5yRl7ZYkyZxTdf0GDRmA+gEuP
nJTIVcLjsf9pgt2pgwS3WoA02fzxjDQ2/d4JJGujf1Ig5G5x0cu0BwDf55qUv+bcyyK9/NMYmmem
iZXjcdnRHKcZdzLTQ1S3MAldqVj+0vVHa8YytFCLCfM/4jArqSoyqRkSXAGHguEukuEen+Zy8Kc2
8Y6QLZuxdl/BHvlvKap+ABEmw6GxNNvyWOXjIh2vDe4shGY7PZNffsw2gAQpmNU9VHuX5sNhmkGg
NIZ34guuYa9dKnKsZNyNR5yrzZOz4GiQAxg1I665HgT0nAszzrXfHiDZUVpd5Z1nAV/iwMNoh3zV
KMHt7O5VOI6PotBl6ICev1NH42gr4zy58G/nyz6kHd1MkwOy+1c0o+WuLHAP/VPHP/k09EjwqfQ3
bHewGVBJGMprGsmA4HUfEi07s5q7GgWdhvD818uNlb5i8phd89FPuBRHy5MJoHfj0XAmplVm6vSz
pghFKNDOTaox2ntVqbKeeDyAqPndL4CLs4akIUvCt0SnXDQBXmAbxrENSpOKEjtbJieYk6cPwPQf
zbpa6ELZMb8eYBlR1OaSzqyWTkF0pEjJELNYlvLkoatAwa6ExuLZ0d/COgQ+feOafbGHhK9+vJ35
o/yX0eOYu7AMbK883Ou8HRvhnYC7hK5k9EzusTiXwi/Xp1Azihs3pKE86wUzB0pzv7/S/iEf3ozj
L0HSTzydGzfV+umPiuh4hp3tn/VNYWspS4XkjEr4vkyfLQ4OLlHoHoVz2ugGq+uK/nr988DoLFXd
8hSe72cfUB50/J8dicGJFVdSI0HWxqQgtYW5ZmDZmv4ntzmPEZL78mOrvc6wMn3AwuooRPBXToae
c3wuVpdkd0PafajhnXAmNy8SNXpY2/MNEVnSiwAERE0sB8N9zMZIgRYGtxAQLYa2ExMO8IJQfaud
aMMjlL1EVXb67Vj7v81djDUoPmFzZOm0ElsuDoOoql9OGBcwd6n2qil3rWabgMK0BRHmQ+2OnJPX
0u+3BScdPILAz8gn7KTtAhS5BaXKhQujoiG+6Z7gdNDUAisIWdAbX0W21acP1fTUw6Jw96ZIL/ea
ocPDdSq6Y2MmkeWElfTKqypzNu9vdB9/HTmwsvdyJ64ZTn0O43y5vbh0S0+/b9OIsmhbJzwU1aP9
Bn7Eop0i3B7DPOUtXlC6Ku93ImtC1VnZ+Pwtgc4ITvvNiOPO0NClzoVm5BU14FfwYAtRM9LDDCzO
ZYGMZ8PbxcFKoGnE3UWCFfNJvUM1U+sQOrS+bg+h9kXvJ8jHgyGaxtNvpnIjN6tq+rL6DAPfvjjn
NDf4V1dE9tsFjvgTx9gI51bQLuQgNLbxFJi4HE9lXaIezJzl/LsTui0SITuIS+IGEDI7TyAsXMGK
TT0uZTW8xX07c6uCq5L3MMPt30EEGGhH14Jz9kmMyBkBGnEmqcSWYvgIpYOgdwWsKXf/GeD/vBBX
+zoy+xmoaQi0w3L3du5736sdJ3lgjFChVz9N7tw+pwcy33sOhqmqj6MgKvS/DN2+0T6ehs40iQSe
duMujOensYNNZToV5YrpSPpoDCgy0JR0C/oi82I8gSAkhzjR587cRIRaNlR56MBtCcD9LH5ZqVlc
GLPxRDjC5IVnbixdtLaZXKboCbvhfG+vm2zSO+RBVhyzBfUFLPnpfrTb8ygi+l9gOZzna3M0OvId
KY7b5cCM+xTeZ6ri3HJPuO3L5WASnDs7FDSgs2meCOVKjqRiGwGHpM/VR6OLMnAjfE7DDyy2Uu55
1EdqQibL/dwT87jM1n5/BjUdkjs3IGrqK+wrQYjimeMiQHLrtT95HMhkR5exn607H1O2WelzZzav
pz8tLkcPu8plBBuJH1yeK+lfJTpZgzSO5bPrD2/6u0FucUMiQb/Tkt7tono9bHGGKWq1w68peTCq
on/4ydrguPCZydjx8rT4Jjn236//irT8LVT185H9H3CqPao82WyaL+FTfz4dF5TYCjieDPSPcuuy
catm8XLs6sH1CtJofRlwbXOJgZtXVyJsayo2QoFg0vb+9+nZ6qAwTLQWM09/dFXjf+vQcWXr6OYO
XNWcupcui4dVS395IuoYXyCK5WTdZgdplVqdLn6y/UjiFoxdUVSXTvghLn7DkUTjtQL0gZyQSQC/
rjJfrrdCIvYZeVRDsZ7O25G2gLSNKlEy0+Nzny86LkvZSqHGwSzBt973ZowEiWf1fhkbjrwkKkUt
Ew0K8/2Zh68qO3R553Acbc5oq11AJiNIv3Akpzqthk3SvD65vzMHGKnLq/X7bOqeOhV09KiM07KX
gQNdnRGNyIbL3mBLgKOev2uPqPa0EIHPitmyoTZNcjHuuwZc+psQMOGm4UxVjlUFXW45B4v7LMig
oWIm/qCLYnY0YMZ/y8WDDmNxcNfyfzyKKUGtNz5oYIWI8Qs2o4aQAYAhy7Rz4HMgHr3sSgaVpX8B
kFDxfcnhEGxy4J39B4yarVQAtvMbuemBWYa3Qxn6MG3yDZnzFDjtEp79ra4vchLSQ4/1tqcw97TP
bjgqv3PQYywjsbNu9/msQUq0z/SvWa+8WGJckdBE1QlliMYPCQGa62VuijXJ0R22F2jVan+xGvYY
nbxcWwByKMhptgk323aqYcJYfiIbj8iUupaQ8QjM6sdrIKPi5KA1pThZ911VNTxUBQtbLm3UTeh4
tGaERM+Vo5C9JI65BFv448mKvsvfLXbNsnC3GCGRgA0T9MT2zeiDwrF19I0a9T2aSDBd6J3vGA0G
97irqJPsnO7j4Q/BVdvkmkmKvpQhrI00EFJPJumRlXJRin5831q/tscIhGMfax5OkDX5nem60atn
bn4kRVEnSAcoxixCAqFArKV5mMfUmP2IKChGj1CpsEZW4H8TJkzAgC1+jkWByqMGK+TXApl90sRO
33lnqk1Com+KLonKd++XiWpi4KfRWIzahxKzxY5MyMj8CZmu+qK6IccCNFhigfRjldcQS3gkdAs5
FZhjM3Grtpvl2iQRy1X5bCFIMwhe4nhsMgsElGQ8WOBL7ixQMZdpl//bNrkHDwXCbDzYDgmZo1ua
fX2H+zf6YPgK2AvBoOCMLPYV5auL6UCOPc3HXxQwm1Xmu0YWVTKfVkI+wOqXVVAG2THgj43as8sg
kM+9C1Y++0exhI9Tu8ysgXnIOiSxiIjrWKQ611KHR4yy85OA30cjyUohmRgUhYbAva7bYxjYIn33
9x4HHmedWoJpddCVda/fPnNU6FPzNYzTKOidOb5zYa0Mw9XQZcGOPJAezBsZVOrMFvusEr5NVWIA
vd5xEyquumvuWL5D0plEZj2RX7MpACUp24xgBxbJtTSpQ/iF7H5VpwCtiHgM8fEEU2M2ZVV2qeXK
vcmvsm3SbjQ/pliMmIqXOEq6BNrzN1eXjqL+8/ddXwG9cCs/UhLzfVV+9DB4F4iWjsJNq8Tfqeys
KIsVTYU50IoulPE9pe2iQmDvoAU9egVNe6CeBoVQmjOWGhBlhfij/WLLbNgYh+HYjVvgH0Fo9U85
j4YQ2ECPbo7RPzFpO9ljOkcC1fbLTNSUeK9ZhcHC33L9JyUN9PJuuhC+2reYBCR5j87ws/0fLaeo
6a2hpPMZEVB+4wMgqNs22gSouecoq5DiFHMYac+VNgr1sTIp4uuyWffJIkqyuUMfqDb+WL4vKipg
Gj+l/8Di5/iYt0H3LMRcpmRhWBrafUHuNv0byS31ZxL9uGhCg7p4+EYUsbF9Dcjn9enKRvjAGIVP
cvtVcA2EIn7NAToYi+cZob0LPAT2VIT9/y+fvO5f2ahrQweRK7xfUQcZRSnpqLlGl35fLsWL35IS
oWL0XqOKuayFQTR5YJ72qCg4/Lvbo4qhW96RASVSXh6LIRdsG3WKMwwaT/8cyiZNWT1WrHcHKd7y
1y4HVyfKiIyMqj+kxk5UH2UTenasDc5qvzvP8u9AvlRCixdYiMmyZr1rStjDLAtKeRbNMXTdkvwr
QKImPTx0FYt2CLfMo2rLiREBnUPQCkVyqCJ87qxcYcFcmnuqXEOMZbn7nyTI7p3NB5P5ZSqZ41g5
8ZZmf3UzeN+BzycbqqRkqB4uAEtJW44r5Vd91ENHz3gzxy5rBwzC1NU9RDPr5Ndk9sfRpISOmTU8
lbP+mMe0NniCWR/0vX/JGx6m5DRFHufKAvwcP1rF7HabBYsHdfziktlwITcSfRLEQYWue1DLgEUN
LleYezq0BqMz2dhltOZvNEKhZuaeNGp2d6BuzYtLOLJo3eCxdJlJs/GUU8o8feRvJWFQWA+3JwqB
l5/Sa6mX6TSB48dna2r5NI2QIbHGPfoSJFp9rYP2323AVdUAHE4/ei/KVUNm60eB4VmmwsQaccC1
PQnGjrHtQUvkLcPzcrFfYpxegdzZW/e7Y/VizxvEdJnGRiKeqN2/Kz5K3IRAjDRLd9cWB1kgkU3o
539NmR8sMtIzAT41JsLfaEZOVXkE6U81ALVQlzgR5auAp8MYqcO6MF0ZDTB127z+MxTo+lXY2kBI
kTFYaUX6g1Q1FBJCnvx+XeJoO5JiduvihNcqozY8hM3lbAKPIE5Sz8jouOI2VHk9LoFZ8gSDlyuJ
rxCg2R45wVhp12fgyPBuXPAc8rpqHm5x19teXNb0ucqFdk6ANiuDhGiiinksyfuq5H3Dv4CPkmQr
J5BJS3IkzNtxU0Ayeq52orm8acIGQrAkFH90bhZ1NEvtmhBwV7Vvmrk/7CSVBUL9Hx81nfl6/lJf
zdRsSXPkS/Hr+0PqFpPifchpNHLmTI6vriOJa5m6DaKUJ0SK/5Xw/W4r2nHVACGx0YyeuPIxz1RX
e+U4YJHYF9ZkkRm3A8LOf0a+K6nDRMpqhxrUlkKuODRfv1OdPgQnlc4w3ZBXxzbdq16TJSpCSRf+
oiVl/n+ndPgMdj/kzIEXlLyO3AC64Uh3qqYjEv2XNKHgdBoKwjfNaskxjFBpPEtvC91dHWWHGkr9
MqU7UsJJ6FiYBnmPrkG+uz0Fws5d83w0IvBcfF4IrdQ2dzoAkZGgAXvtZtF+RIv7VKZuKp16lIMj
VqCX5D4m5jfUNINBpJDywL+wfx459TyjUtcA6LhLwhyqu5iPly9HHgbYfBEZmpKeo2BUhMXzNdFS
zbq8UQywlcbyURWOloWWk29eV6kuXXNUjcBYl5hmP6QnHTb0IVegcClSn05bYxc+eyYwAnLYHKYS
ZL89tTXoOXcrOW1N03AVIYfH55WN5JbxPtR5bjxctsT98Ote10aoq8c+hhFtWUOInmA9c4sh0Sp3
lvYF1Q7dk8U+ipmkCCxyqhuPx7VqGJEPbKtEsGSAexZF8wCzF0UIEnc6nkYvOl3GpDeolgvV1XMT
LbbFt9N3OVHYCtaDNE3ER4l1RRXvX6TpZM8E/yZTdlawoF15gcglaKeeZERme6weikAMt/lKCkoO
V7DXr3yeCtVwMmHP/8qIyKboGtlDUEEZyMOmlCo4ecXX+yli3aNR2RGem/omnWrOyF3q1O8CZvLg
0Zn2Ey9BT2TtBlXFLrRmfB3N9kYWPtBLOgLw6zm6AKXs43rl0yfLS29xvyzRntPNdJzGV8RJWECk
/hbWCQMytX1sxsdhWOKvPBFyNctkyhhxMwpky9+/JsXAHySkTjRhEddO9C4ph2xI59OI9c/zCtA6
+tV9Bxfq4fFA8fxmo2d5CvzG2G7WhZfQLLxYB4gC+WcGeX0qz1seLXQjS2L5xHvL262uNU7Niczx
KbHp2UUYsx/10jLHHv2egVZwsb2BEe/MmJ4qZkqETcYImSDP+GBjC7KRs/OVx/rYsjxpJ1clor9J
74cRLKamWdRUBYC5NLt96OZsFm45AOr4uP5aOgigely+teMJTc49j/YBnEh8nm2TzYoHiFfiD+xJ
DCGk04PtKGFEcKg3nO8POGyajqV53yQwZVSgIq4IlZCjiyqxoJyatHjoxyUYVzzTKN0SEJAraOwI
IuXR5zazsuNEbmf9W/W8DShzyDVkjpIKy8Qh4jy+dNz5Owb2J72Y4wryHsY+2Lx636rTq0mgrM2L
sLsn9e+gjys8ZXkV3I1VA3J/tjreFg0Ak5lTta4gDt81/8X/6qc1FPsDceh6gNS74qSZGWs2ari0
UEbuZkiFXvqhD68djvaxsnH8D2yRsVIvt5BjV8xBeRpxj0NxRCifRGZ1CypqueKAUiY6xPZj6dHe
RKKy/mzxnwqpj3ZvZ9rOrVAR4SOhfXQuy36iy0N/SyBbKrtMFkGbLdGqqJX3hRpDt66N/VW2ZuWA
1183/Dh17xUr5HvApV/+K75sBtcUJ+LbZcBVpjAi7r3hY02maAZOYu9N+1YxLZHZS8MCcTwjcQmx
qQUd6JkXYRFjUSwHyBo9F9gJuzwNX0f+WGRT9yQih7vunIUuRIuTQMQJbizPWyVnMd0j3XrRZ9oC
Al8uLnjGy1ztSwOHtBxwqfZa/CJtoog7sv1AeIX91Rsj901lcMTKq5Ap+nvmlsn62HSN7bEYSnnC
NIhD9Sop4ESKsnGAV5jupEarsgrcJnlOnHIGbtJf3a1cuiSMWPqon4/IiiPVnUEYh+QsrUBsnSyx
ipjbvsrirgeiHD9fczFZUO9Mfe0tGRgU2c80tpVo/tNWr6M7d0No2Le6Yc4sAv3jVLoFTUYaeMMN
G8GL2P5iAJNIeAclWEuCb8lF0CGSDW84yPnWMgSelGbWltWFRPpRN5xixjyNc399Kaydk1+XL/cw
QbOBMbnJ3YfBEUoZi8GT3B1SBPh+NDkM8cezHt5JISzyUkgE4IsQUD6Pa3VOpJsTS2vxx5Aw9ExZ
nr9tYR999ocY4NacaTNRi3LIlW9BZdSjhUh4KwjYBe2m83cUn8illcylpda6SIhaqp3yCU06WotU
1pRgn+LeQut2TRAXfNCkZkxetCtLgGrupNZmB2d9eYxntIJhF9lqOM1c6r7pAFCzJwDJm5W2Pwas
OGhqGsfS0avlNGRWx/9EVnA3sMQbdKIqE9kD33G5dXt5qvXcLr3sOzr9PN29K+rwcNh4KOYQPB44
B+7TfGuDpn+0wEIuA4pIFA3i0amf9ndRBetUVgqhnw+dJD/sxJ6QK69cR32MJaawekSSJX4u+Avo
oF4gmCluhY9xCLVbTcoWPGVRzyz4xx6627VNVhQv9tJJj61Ng5sxxOcHNQcjQz3ooc2CeEmoCrrY
kuFKQ9Cv23I5se6lb4/4r7IRROzYtuSrl2itJ/QU+h7iHj17pkpTz8QT2740puAmKRShRAO4EYXT
Soufm83QoXl7nscwhf3ezLQtWtxEV3lJh7XTy+a5yZrJw4/fgTkzFNCWSEi4pbmGtrxXVo68uMJV
nZVhoWn2aQBzRsDTEPDUWZMdUiydnRcPehS+4SLpAApS+TN7Icq1v9S9vMjWhit19tS0n2nMV8JO
3HYixhbDUwuDh1cv2YyMpNsUHZwUnuI7iwj5ZrhCXB4QVohrgoICq4aMJPBl3GKVUc0PoCptoqf6
CA+OOOpyj/0Ilte/iZWIDCMv6ZpJQnaerxVAjGbFOZi79I1nHVOLjHIz2CdiHH29fVFpCco8v1N+
vuhlsuJMZfuvI+VQBxgplsIIZ4zHJRHa8Zl4XmzuSc0kJMLy1mywSt/YgILvUHJJinALnz55GWUm
jj/zJVT0Qzp3RHoZaUuJpvvz6xdPOhvX01sJngLBkrJbJ4EhY5FHqy/x14zchlTfz3LiqLaq73dR
k7Z95W1wUxV/OhHvGCENVinnMOFLyDOz4OFbaF5WczrBd8/MdUV9NJuzLrfOg0RYt19dni4KWGB+
oBYa6LasB5CJ8yy5H/q9gIqdpDy5YhJ8ey4lqLvrpNScV5BwRA14jam6GXFkVYKNz4lsRBRQ18Kw
QGGhaXzSxpgMphhc7FUQREtch03kXlwI9oulf0saGnMHJMI1GfNJKctoA3s3v3RXvtPBOY3mWPHf
ayFnQfSaSqqiXKpeZGIazBKUkXE3kMJ5MYzI+lDvGoBN2tq/3vTVvHFwrQMy4ixURSfVLogn88oL
iGCuP53upUTLT6RcUetDKqyXCfC3/HikwGwH4Fgc1IFqoPvoUAOmPMDyeHJzjGLQbeu6w4//SHaB
FUSY47cdUTqs/saN1o68xKzQmgGDjliqTGbuDdwrNAxcQKURS70te8aH5U0xZa221amiQV4KaWCC
u+zJPpS/6gkm/nff1zqBIp5A+RnASPVdBFTL1GRQkPKTNwaTr0rff6Tp50eldoXZRr1IbdzQ4duq
DT7GP6woOPAko19PArkEqgxsjofF/zaX238sQ4b+gMQoI43L8EOsvb6CKRa+kbBrdJvwKKUNZST2
tD/TXmarcmMEMwUx3nooiX45lbtCR1Ot04SlkmKkH2wCqxJwhsg0Dcb3tSxlkuqQlRFZNXbOmpud
O/Ply5DmdP7QlnU9FxlEVLbS06dSaO2H4UN58+Bd5LEzm5rIPMJtDho12GKZeHK8tNBPqta49lwL
WCJ4JoVsQXKcJpwegMRJPVjBmwB3JnNEUfjTg7bG/qqFLeeqX8uI569j3EhjYgbdnsxBgDTKUA6o
81jAZtb+345KatMeCgcJ6cBKdAw+qws4AKrJbqpsQaCv3M59Udez7dYieF7rvlV98aVDWuybI7IM
QNKcucribw9jIArL4M5Iys/5COZC/8vzDKrvCNFz3lXUM0/5Hi4rZXIXBBTlz4DhKWoxH1Cm2feA
uM0v1fcLYaiKmoakkV529C5KiaVg/o5rKX0f37faIKqdkK70fUSQt2hFS+wriShd7FfdzwvMmyJ0
oe9VTHBj/wCLcVuvnplvHCuXFDYJc8h/PYlXYER9XttoxTDg3HEL620lPf1kZ/Z4BbHQqI59md3t
kvyHzbbJHjyza3eMYM3nXZpmSiT4iJom7BCpJ2OyyEAj6/2i2cbE2jGR+J6iTp8uVOFx3XTsTngo
s+4zZKmC3WA3hjUtCpn8iyuMNy2YpUOdtO7talvuE537MqIvEJZ8lk68CZTljyjKLaufyE0RfNBo
C0Yl/A587/J6tcUiXovsAXOOfJKG9qH42qNcKXitEilYo9WNaUXvs5ZxpuoVRn38mWZzEUJqiYTS
QEtxM8q/8W4OS7yPyYVDCtbiW1wANXeN0ZDyVrYyvtIzUvKjZkzPAhOZseMxDtVJt5wd6zsvdEVl
XUupFtOJlSoQF+RYv5k2tem46UYmdHaNtFh5xPK3iBjSBjdkR9bW/FL7hyZ5b9lIlrZTzXM0Fr1A
KnFmF3D4MIeys6dP0P4JTdAla7HiEpkH00x6UkfR9DqawTFtUVEs9zz3LpMbQ0veLnerVBLF8aYO
qJy2QFwmcdQqS0hpoarybFaP9Be2jy2zfifrmNgujF2458iqY2mQyQfbyVaA3oNz0JV+sqhceau5
lW5jOULNJ5x13T9dmmBvFVd7kGLu9hoGoLizwWmuXgEeT4g8XPW0qLcMPtfV9NdXkc9Pr5r8Wkpp
hT+kbUQEumVnRb67FVrvjauOp1EHB6ex7rn1J4sJCfGFRvp59xj4uepnYgcPN7fSlyiV+rPrduEU
Y+R5L5YPQMXsE9pXvE8SJJJ0AiiDUpZGMqhikRdGls/TskKMGOquuiws8nh/IYqvZitsLr7iThD7
QZwgUqJjWq+sbAXZ033a5FyEMY/DVK+NFGFphk/vRWhyvprg5ZHR45Oqh0WNkYjUW+5MeA8qp0IU
Lddl0uxQ1wBBEdyc9psL0d3EmhQhDbKKcAfXAwW3xGiVTUOBwkzY2zeIMo4mUOIEkMYkcJU8tpGg
IG85W0vW5TpSgr4Zbk8ipBKnHR6FS8+Hsls6njwLnbXOGXYEpojZCoz7fQenkLKwDb1U+xJgWRBq
jj+TbzJ4UQ/NBIi+diaKYSR0JdigVfxVjouNAJRhfEq1Eoq2d/sjy0XwcAgOHLFimpp5jiiJsc04
E9vpSLSmao7KgvRnWmBIyLVFKvbYWgEFJxi7dL16pdh8N7YL3eiiwM5sS3rfG4/0VrQl7EIw6724
nNMWmJacuJAWEiNyAbSxvW6xsh/QZBHniszOTkUHGCYB/9Ry0//1d0mPM7QYfZ9AI1CO03bJiF5W
UvxCwaW5JbZwPh7QEmoNuVKgT1Y7W6j9ot8ryD80stxsyYdfh1E43+nM0ygWLY8ldgZu1znTDG9c
a90vpnYq3kPqfUiqAk+wPynHPSLiMXA08/kbJ3GOTXcfvJmt+CJh87WmzTUZF6knKr3pi7ma7bEA
iVpUkysMJ1VN6/1sPIibotPolh2TBGlsQYFlAnD17TWX1jhr4IGQFgrPGDwdOYOa6Zm5oDhloexw
oAzJG1Kwhler/YiO7i2hRgck+gT8+CEnlT2b+R8iSZbZmjovsbS0nKm5F4nJwPjP2zj5SDPQpp5x
aW3du4R32HOH6NeEshLIRiOrQwhykLD3ZySMhdwe1bSSt/OfxO+x72AKpudqrBx213vsRZ32UnmT
/mYadxUneQnp2enRitq1lUXkZ7YCM1J5vH2+QYub0r6iHwR00MPzhlkzjwTsln9EhcN0GyL4E2h1
8ArMQ1IWGpgd4vYzDM0E0x9LAGqeUBZyjcUeqNdyVEK6ty9dBlFP2RvU7JyV4HuWOKOMHzWvKYSu
/+jZukABjY1OXHMz7fbQCSBJ8Ljj/CX/1aJLKUcyWk04spiq21sBCCCt4SwW2vHOhj3dvPavg7/w
8XxuBrF6QpDvSUQ3NGJb4GqSLEye+gWiV7UbWy1UGogIRZdz90KT+NaGmkE4WH0/mk5Qywbhxw2P
J+UMT9FEFodC8ReohQjnkSO6wSN7p1zJylDVWka/en8uU9YW94pz5vPDx8gCxCPoeBrbaB0nHQNX
CvRgT2H5Ca+EvHnpwfYAE2ykDdLW6CH5dykLbU4EHJ8wXKA4BsqsGuoHvj7S/uyhPeSHOisJC/2P
97f3+2Cd/MKmTI0oVHz/JXoBbAdDtxUj2+mAumfYmgwV7nCJqboc5WOc5g6y8/ZIiRKeoaPKSXMi
NYAFMC7+FD7cSCdy1f+KpHDFHb7CvKnISQ7KdQDBHRdHypZEHC7/GW+Nd9oE6dTstu19URWx1M+v
iH4rd6K7CRfAUmsD6s9gQ0cw7GcQNUOfve+fyMFOg4U/0MMp8UGnfN/r93mG/YL5/wYthd5wLLzc
ExeKXGFoHoQnr8RAHb/AiIMzumr5AFyRfOSn6rAjURmSw0lP29mpj45EShUSBU/Qqa6o350Y9iHl
DVON6bF3FSU2Iqk5jVUspsP4QuFLfiYv+2KlaD10WdtAEC4cq5Y/V6f8LwJ1DF+KQ1Zf3ZkYhYo2
AxmcJbE3jdidCW6rNh8T/lgQ/Yh6jkv+0icxjNwAqe8hNTunLYAufjlbuTVvZimgV+qEnmr6P3kN
ixL5NTYUhPW2cVAc9VNwAJrFQvQ1pHX8KxwJo+WrQeMeF1jmVZtORdgK/w26UT5xSBFPJeUSHkQr
L+fcI4dqOTd7yF8EAELkfL9yJ5pPVUNLyCmWa7Hbii5k4c+m0t8SgLe9zjE3g7AV89lroEB5CjRp
g707pc0sDF4dcvodNpp6l4O1/Ioq5ht/MOSHLYzFley5LIckqjDAw340+Rb9D6Dirwzhvubnmr9C
XbQTv7ER0ik67rzwm+8zlwudBPtFLDuGnNtsrvCCe13YPwobCvhqENaQs9tBm9slquvDFbTjVc8R
+dviUeIn7RbEFJFGx72bLGNRI6zvkCDxLv57EtTNQ+OUEGi+bC7ERM9QCzwlpqJqe12Ko5vHQn+J
Tcs9brezm9wxKMsqgHNQbpw/x9U7B1W8x55d091lw40caF0cw5uRzp5k2KHqyam0oOUOvtxdYzB9
Uqy5j8+IUH142Yikt/I6NmssdsLjNe1LEHhgOwVr1OpQE70ggq/hFi5/yFjx74Ex+YJ5q1mnz/fa
fUQ75GNiOhOsOHnwZLkNlhgPKzABcLOzpwAIJs7Ask2DnK2KwJi3rIwIb6x/z9yrS5ZV1Oo9xzHf
uvXNj6MMLuG6KeHUULzbrwfbyxT+K0Aa07GyATsB9TFPMBZCXUmuGaIBv4PttgXJnTABuPdhi79N
R68JCszGz2sFPi23fMNTyJB+K574SiiFb/nxFgA4IawgvG4vS8hxVaLnP6BM+l8Gng4rdBkQKgBh
X1I3cx4HtcnKToMITc5Veu4OIvYC0X39ynrN1+cQnHd98CUKx4zmy79M8umSX6o+FCXPHLG0aNv1
pN3LyUxu/1YmOBka4CQTSaaLBRNb/tafsv5pU0iYbPaBmjMPWG0Hmd4gRrIeWIKlq4DmXkWJIGw6
r0QgQKrWw/ro4MsKMa7ZFet85g1Jzs/FN3oJiMoDzGSvGImECtt3Wnmw7D56qdL8EgrIrje6SfkH
JuoEHELVDyF3Z26NsxMnikLnicAEHGGgBVlSg0rsR+yn5HGvlljgQT1oK4uh08k1GKSJgNQOgPZx
my/RsdiiQ48dMkYClKt46Sm325zcRCApczR+MLkZ8gHf4UBHQ3RTzh/QdEDS6cIfGb4csGq8BZ+H
MJMgy13TWvpphsMAR4hBCJLsWf8YiRCq1FgAZydfrnOF/MoItVk0GMnQHZk0619xmYk7v+ZtmV4+
8WsoNBpAt0TafaWrezEpnikXv4sVe7rgKinujS98fv13kEm/ONggv+rlvG5E25AfmDTTTxXecU+4
5A2YTeOHewxxMpR/rjOrVaXHe0PGPRZ/kQtGLOKp+2l0CYwMrs7Jc2YI4CBi1uiotVxRKh4Q3mO6
jvT8/4tTHiEO5riD8veO02137JVHm6Pu/g7MFwGhF7KTwUuUB9T4vXWfq3/c1UN/4tFJEfMV0BJb
18OOf8w9r1HIqGRaHDM9pfCmsODPpWJeBOlGP0AIRWbMV7e5PPul8IO0tcwCbqPNZlpOHInWMdur
YlGWyaAhjc/tKye5LB312jiBlE0N+FzB50nAYt8qabozcjsnaTOoX3RcSWpwCZqI+hWUCo+IkQ4+
aEoSVyovIB4iRz+m3lN6uDEOPLmURN7KaZ7X3+Kfsy0Ik3MoAHMJ0oI6YxGAUEx26pQoAQbxJvbV
/6YOGQTIEKA+gZKTCt45H4hklxDTjkgOVN56GnvtKLx+7/ZcXg2HL33uqNq6O66KH0Tpv5Tiv0e5
8TNAeYre1z2Cx+fEXxrvIMtcXT09IBMa+ph0cmla4KxYPGc/pT2GP35YbnatV00r39p+OZET00Jz
E49VoCOURFeJshASOjnjPKTux+z8xD+mzCmbc6o6ovuHEwN3MbpAOb6pgozgKNWcZH/9bV5+O69y
jVQ0revmvjpGwFE5/hNuz36TD8SDlpwCLIYxqtppdChMRIS5TH/91NOevqX5KNKsqhr7ym9wtYUM
OrfCk0Nw8J7LOhZfj72HUUCGGOnM4fD630b+LfW663BNJ1aGNbH1fiYy7lqKwVZTEdoMjq/fB/Mo
juKkFnt67+XKIFv1Z4Q8FxSCoUXBf+pz+Ypfpw7odqfPJgpwfMqA1KXnPwKGuk6QedjDd4zlXOHU
KvdMrrM3U52aD4xEWetSouk6Cbe5RB26o5ZztBQ6K68jBtXWiAXyvwGYEcFi0J3C77XRLDneJ3PH
7KxKWdYrfIqyd+8CHumBQcZW5852QtScLAmPt3I6ng5K4+j/amZACFNDR4OcxAJbzyRNs0CuRmJn
tTcGFfvI6cJrMsEDDE5UGzy0zsmFKstOraMuL4yol5stJz1yxBIbKSFXaDzfDz3d9N0Ys+181V4F
Mo39JLNxU9usAoeaWkRCcjwcve1wSmt2J9eHHwM6/KICmJr3nzL2PqLGtTR72w+FGubFCIxJsKVa
lfchwwu/OXHh2WWLbJoJxs0AXKVAYF9SJgPJAZ+lTV1kVm7j/q12yM54SQm5Yu9/xuaXnWdofOxs
ZwMcWogIUOJQdfxAmSk6nDVLgWsNfV6Gx6odRQM31XxrULIWkwyGlvrORgoPHWlq7Hr6a5W6Eqsz
e0yepjOpwmMycTrp3Gv7mhrZD11eb/xYIWPDYrL3aCpYCSOqNqyV36oZqMjUufhXAo+e/YgHjeIs
Q2ZuumIZHcssDQjNoTexitH2ZHgwd21mRIAlx62ogNLMzya0BxjGCOIOKqaJ426nzMvthR/TxjiG
kWLTd2funJc9d3XQIl4rihRinZEW+PXaluaqvm0UpD68u1eSAVPlCM16nUNKijCwcRnEYm9jsnVD
442pKapLo3+C8Ulo+Z+H/pKQsDyIhOpB14fVLYxwVHA1nn/vBeq8iPv6mNpqFlfzyrShUqz5Rgcu
fw/V4pEL/1fRnVbjNHCwhnDS2u0fSzb0k7o0IjUu4gq9nPKm8HwBTv9uVzMy9ZHSUOaajcCjGSn9
4zGOI+mxD328+azEkk9vWVgJnXljAaYW1aaK6JwGyxDEKRDPpUBLwbcAT8js5NB4cTq7GuP4fFfp
NiI6ajWwVyycOfVy235VTMvkXMeRlpm4PNkzyHB7VABfrE6tcJf9XN6cqYDUYoMa5i5vG1C3jQSo
6mWOaFZw2HgsYxX/YI8jd6uruyoluUHJqwnQUWtLH9if284N8wKfLZ4PhVR435zfqFOKoaRgS9SI
O7dYX+cJODbcxvdnRBi/bZBfP4OeP+vV8djSyohPQwnelZdxrrbH0LGEPpTHtuMiAFZa5vJdKto2
Avw13TYD4VPXB81G7E1zffJmO5IpQmsXIJiBLURnpWfE39merHmpXC9P/5RsiaDVnnrL7LTnF0Se
V56I6qQDjktk6qbCsptrJtCm5blHi+fhCwaUvbowycNdMZ05PVo2btpNWiCOYVI9aRRbweFgLu02
1/5uIg+gEmZA04+djNRgCZVw267l+7uI5u+BJFcwnJ1epgWvBVt6dj0+iCWltUil03QpJ8vSO8eT
9c3y69CkITC3qqt3wxhzVK6eculUNz1efYL3TE3ZVVxGM8r5cRZFDK/b6aom7MXgzE3laVxJqALt
31W9jbx3yaDYn0LX6bNJVLDkjksn0Aitic/xomP3MUYQuElT8MYSabGq/1VZZwyj8k8iwZFR2Szg
H5r23FKkj6te4Jprshquc8gvXn+UNdJO42w1oOXs9I/E50MWwcZkVjZLl2zh/Vc79ihvvYsZNpxU
peaXMs4MG4ujSbo73v76cJq4GWc22yv0L77ewEPu4Feak8YyuJ409WRgNB91kJzX48rGlo3EX9ea
4iKKlpgtyPibURdasFmlLKZVmjwfz1KDmzDJDsGL4vUf2SaM/tGdgWyd9d4udr9/u6aQ5cs+TX95
pUXi6osA8iHn7mNfuvcwIiG/rUb0YntRY+FjVSuIUJrZiAGbZBQf8P6vBy2FExrwDSkEoTh/Ebv3
Qnocno4i/JJxQMbLMRDwHKtpJXRI5WZlZjzIeEFFo0w6KkHgIUfHXXnhej0ffKDXSrdLq+UkNJL3
WvXVbAdhiqTsoX8YVl1FoxOAFU05DpGbcr/OhFVqngwvkM3HaMNi5TnTXWlJrArXrdec/G12SDqU
t9+SmCTq3d+w0fznjuyC/obn0Yi97EtIKEYmFWtcfcRBBcuZFt6KoEdhDG8ZVWo6YCVgram8cV+8
xGlZpwotjYAA46r9veTD8Bf+Ur2Cg3TXoaMZCdra3gu6VzBcLh6FdNAtKr3IpXVCr+XQau4T9p8j
j3+6V5vvoT58qbP2DdhasXwOc88HMTKYseCtI1MSeJMousGGAJlMQnUnJlSGWhYxDJHzBmiajN+P
pQ/+ogL661yLw0AZb2KzyGdNS8TDM2NpFolNhjpcEyVI1+6JHbOvS+2OX6m4rog+dedw3I9NjVQP
z1eBVLK6PqSFKX854rrcsPiyKwV9bPjUISlShnKUTM0rFZq/99bgFMEZnVmMuwUxn1KP0CIZFaFV
ehpWvZlR/rkk755Q356czN1LSVYgveQFgbXlKyWkmI9QDAeVzZqaEg4coYzABneYxNq5L7Iu5USC
eAI3tmv9PquEiQQoKl5TWZl5HgCJAubyMC5swNZvHmllZoOZ3LIpimklcIN8iZ/8MWMmETIAS74h
mIguN2hmmybwpR6V18cJ3eKIGUrtcpdAIGvcjLlkZOBD/ASJToHE2dyCo46C5P5PEwMiSyiSDKTl
l+9ZrCnzWScyQF39NiuB2dHFwpWzpF5lSTIXI1JZxEtG+O2b7PlsdMzXkqBPCV0Q7gU7Cdh/Jwhm
FjYReW8xO0/gP6SJFHMTUA8QzfvK/Fxdn2X4zrVB0ooG6aL9Xqnu9R22peIfU4y/DOga/hvI+mkx
iFp8TDCfQrhRqOgmzwSrt1W7CmslNLh45Jrtuo1G91OeDzOx9fElxcARYH+f7VHCRMaIqJmP1nMa
OQbpVkg9PG+Kvos7FxbmIX3NVu/hdO8sUHNCFrq0h0xX7Jc94QwM+o5XrQlPx5EjX4hK87m5tGwm
38F8jWgB5HENf9DI+w7Xa+PJRC+iLIbXabXMynDejM7sdlWAoHpxo1ZuR+m+AhUfUbbiKqyRSlNC
5k5jN2iwb1fdYhBP3PMytZepGVo662wJQyyc+Mb2tSuz8PPST00IX+yQlYAunDY2apGfZs90qj1Q
RK/eB3GY0fbHh0VEu535Uq+lsKoRWWLuydi4yODjeWDRfuPfb1j/tplpQbS5h3fwXoT89w9JWUCQ
5EIR8qsZiNA2/xV3zcO9S04WAAvusvGvHTpfXJsA+8pFIgizLH+PYt+RSLFll7AZ0WVwFaCQ3Qc5
SHvLUubOglQWExY82+ejkqvs0VMDi5fZUett6zGbtrohfLnFAo7XvrmUwWciKeTIR928djFmTqyS
doWzVU8IAbYokn5zLlrFS6a1aX1viemhYMOlsWLIi80DEu+c2D53fffzORLhHxSTXUXJiGGIprC0
uI4SIiPYAQzeY66Or7wnQVUM+bhTaEZbPnCqyMY7H93v8zk9tUYeqdgsZw7xU1vLCfH405x1r+ro
9O56pfZqi2VZc6UxCogqgWMzam5EvmwtqHCFJHcOPCiGoEu/qKDOBanhALZc/drYZ1EXX2P3Kg9M
GB/j8alIg8dhRIuwgGnD4GHAsYXZIegHSWav24CJTq9k9iE5HQWnIWa835sSlv28oU6Y453dABKf
bTl4Ds6uONpX4pjDWFwVAKXSsYAq2YhYSS6rNbSK7s+aXCOOd4OHwz0wYIFPio6kdU5L9wye1oG7
sAGKa/Gp2FTbnQeormLXnOfODbI04+sV1SulqdY3zMsUoEmxk/itLKdvhxOtgBa96hwPxvJ3zx+4
BobRccN9SNkCm5Jihambl29V1gSDPRVZnqoas3gtzl/yJ0TzNt9A5VrYWwc5A8ysydoEpumQ6sVx
g8S1JTNZG7whmaajlnKvzTsIEwvw6OB8ykt14o0zILfBSo7L5SjRuK2orPfGbJ0e8a16ohE6EfiU
S5YQP6VwCYYbs43k4NmjgBcIGWsKaBCYzOc84GJ8WCvGcY5oxzOtt9KD5TeSJnI4db1BTcrtcEG1
OIrZSx54WpoRs42vkQC+GOibq7RFSfRPvALt9HQqYG7qButybzvbh/DYOjTzc3dlj6Its0tr5Uex
Q/KvAi0niFMfMajvmf+IHcKIIWF8BLl9evkPPBsdCiuzKSm6AsdlPNL+wYff40M+m4RrDAgod2tI
cr+SHh0RJfQnOdlFS0bW0xM5p/c6lEmGhO2RHppYkSoqOaKW6lS05zWME9mH/yjFelJffQmttcH8
T4ft9NQakuUitJ3yqTTvHxu4ds/+MI02YWZtVhG36a48nGjHl3XseC0Zg8mghBbgpU1sWmsR2bbh
m7ch+CXxd6542hQ2Uelwbaanz6tJnbU9WkzU3wLa8ITBIEEFrZlxLFqhIL7sr01HBwpG/ZZVUhVA
/i0s3hrxbznrmKDB2INq58XMqCEM/J37B8Eq20dGwiQfxek0l5O97MwEwLWAtuWJQYU8uzudvIbo
GTFz/9a39TUvMPe+gJnQ8Her0WW7zeqPN4v0Z+4ABLMg54Yo2Q9P4hn61/1R3zZulZ+J51gM1VQj
xw6u7mUTZlpfQH5qkFrNSHjorWjtjwdQqqSMs+WY/C0Px/yShgpkTK5zwP5aA23cDSj+Hy0NnHom
GCjB112YoGvBmDrau4U0ZxEs5g0nm8yjfPwfXUmCY1ejkKRq2oeng+GITTqKRZ8Eo3XVvmavT42o
7BvG8hblKXMqmW/ac9vLXcT0CYeg+bbJj+5fNbcTd6v11DTslqGE0nHU2O3EqD34UtKVfazrwOWi
xl49ImKwo8SzjHXn+FSEO68BPnKiqC9YTKfhQNLdKhhBle8nHvedHAMRkcO4FybEKH1X+JNYwKc9
U9icahhHZKQSV4FX1brETVn74JdZ1+S1vv2Upr797RVRvR/HwfQOmOnTpuXOMMppbCozvRhE/x8+
IP9NrlPi3L2O9RP0RZaoWIglXei5JFdDSv1n0wa+KfgRz5ltz5q+YjJdyJ680jK//hkaUDZEIlW6
Gl/HdS9AK8uI4Ia5DNuceaoC80vhjrYIKWKu7X9utUkItSbhcfsoPwBgOTXmmFSI6hKFVmBQMZ63
yvuZefvH5oBpOsDrfbjbhVP8Am4wZQ/yBHgb74zVLMt+eJ6TQMNBIpKOPWnRoXvEwYmy3hFcPO/C
uv26tpNmOU6HfCbdjXg0/bIeYJnvTtAXbYplyl1JeFHCRkhQUoopWzas51RIi8OvXAqEjcSC/n8A
lv4TvHceN8x/YDaWlk8pCVt40eRJDqD1fPDKslFksxlxMSy/lktg0vGPWghgRXNwIbW/edPttI6L
ZxrWMh4TIRsRPDPXgT/96tY9qgWsnD1dkwTeY6p+a5QPER6LbbUDDXimd/yyhuk3L8ka7cubFjJl
G9kntfS+rTHfsUD8ByNh7yDt4G51rGvwNDtCifjIWhUVEkTBOASVpyJTJaDluR8q3G4fI1v+G1v4
o4o8PVXXtT+aLynUejAKR84sB32E64tmkiORejI4etIuJR7NugcGBLmugBJp6hyCHLOM83cCXrsa
WD8+7SauXE+g+7FwiMHUfmgMsLyrIwj3M61MqcvP44LnKwBxkJ8JJBP/FYyTKBdpq8p/TF7+apy7
01c5VhIRXH5LTcr6IJpdQHtcX3exhLhFcaAEWtRF696ZUi6dWZKuibt6fy7LmqKVlGtlUCkKhjp9
LVYgavqPcY2nhaxITKu6eEvtiNVVeVTMtgx89/0Mp6QlSE++SJA7b46uVjwTWM+hIZfSQisblua5
XN+FanBdnvEhqqBKjGP//dERqxS5ek9qauJA1RdQB63wFVqMTHefI3P5LGSVlRwRviqsPqHNl7+3
R1UyVXGMWin3QZfnBAJmI26rAMmF/5+LMGA5yr2J1xaVu7uaUonokZ8eS/FdK1aNviZeksHRfc9s
JU8rQaG6HZdPbznumAwlEILLXwNgRHQP90UI7dK67QIoJ8vGTa0F6jDLe9NNvaCmUR5Hu/Nt2xks
DUKVa/h3BjQnpXs42HU0XeAkNfGY76/7uGV5rmXoBc8QmvcbCAchY4E00SvU3yVr8PkO9ubUn2di
7IlQ+Mqyfflb8uc3Y+lMr0bVkd3cqQ7EHWkCvnHZ0rYZCwRzL3ok+pjxrlpFsfh4KkC6+tvyfoND
6kGSAAE13NCrUDjjTRj4yarznsxGgP8MgLYAImmT1/N0oXA5ZCgMNXdh42HsCYcQUbeL0+J2LvJ2
7ONZ3+i0kOSUov+QzzMuK/rRN1u64MuZvBOpbYRT5kcYNbengaXDgQzQ7Iz+vKvvDu1f6pOESKbE
8fZzxuFN7WF3TQpAGMonbtF+bg36/VlVp5aGVwalcz+uIQ6lppc8kbqu985iesTKayLRMz+8CvGC
vlKWwCMqyQ4K1365+3dQaEZ2nY1MR83OWHXwbXEZwXi9U7bSeS6B0579zX0yEZp0jrVKLdGohmHW
f0K175WXaMkGk4GTp9NTgcs99c7u4EpOdExkjoCUL+m1nB/d8nP6vXKHC3oedNHAF8e6Ao0LFKVk
DaP291biwA1FJiYUNFOKXITwqG+93ac2MoiR3s1XR0RbWO9VZBEBdlvvVg+r7J3BKud2QRJAPbBx
oryI9pncxj+q5Ma2rkCI23zjUEzZsXa554CcAQloJBCuwbK5HesIPiYmtdxEa5HUoZLtlcLg9gP1
CWhq+CpckiOzvoouG7IANaerX/YBtZvUT45SPQepDwyBtH3mdzgWBQeqBtW0v74x2hnXIGF7DbGt
W5wbGOX/uTWr0zyK3gMohbKVGPdEGqO55kUpfqt7dLR77IYLKQnAX+982A25GcDJGGJXe1ZlAT5D
w5xuy0wfq7qWLRmUyJxZSNqKbCri/GiDHW6dQ0mdfFjxftidYLFz3DvTVwmh7pxQdSA55GP/QCJO
R7WDOHQciU2IEME7jLoIfyWOdUqhP20s1CVPJwg7qHlyfP2DwbmU2g5L2b+Ac/l+n59lq2jCJ3m/
qo6JUILq6BWZ71WbDOIU9WBl4lZHHvfy0aJ7I0sgsXjqMG28LDU17o5dWHqW9KW4xaRisqYtGRNI
9+g5upYrib+6j3Kgw5ZM5xToxwRZV2ZA+wNHU+xCxwG8btqsOOfhj5j7DK909mRQgxGhkDEt3Ka7
PLN/w6Axxze9H/ifQjF2MYJCxVrqoHRt/h2cZsaxbzdpAhef8Xr31LiuDcBz03W47b47DbME1hun
1auRxx7UvC8TRGVWqWjTpCsgi7SknDn+bCQT3UyYlQrT+Uq/SdrO5jeNEYxt0ZkTM/IHW1G6pR7J
7bg9YaMVnwlOeFc7eG9ddl8cVQwjg41GDZ3pQx2mbHjM1v3cNPniN6yMHxT6YTNOyDuarnTWsnoe
FzUFPfADv4TpoLCgLXhlO8JE8CzUzEBHi07DEP3jFFao/TBwgkWW7u9r185F7U63udLHWDe6uMoH
QMyVSBL4bObgV/fxaM9qEc9gWZJsbIs3OQ4wIllxvap+yVjadjtcjUc+bOzXEhP3K2yfv/V2kdKv
2u1gjfqQGXU6A/woixzQs1EK5k7TuNcXXSAIJZfAfC19GDX4iJ2Wf7h9x5MNEk8wkkjRS2f7FNy4
mZK0Y3lFX/U7esykRHA4T76C1wsQcQrdoEusbV/uG/mxL8m+KvvVkGarOMnbwkCjj9UAOD/4pmwV
jTlfeuUHbHNGqD+8Gdo+1fnl0cvczHUzOv29DxsAR9B/a6LzpDwg7g2Gj3v6nNAR2wY/C7AA3qcp
i1Riu1L+1Cgmm4LAgZ7m65zEMszgBh0mBwx8h0vTaWYeILQRhpYoHeJj2D7ddF4WX93EZJ/s9Kp4
u3XVS73/vfthp/lI8Ex8qUbFItiTH259/nc4bhQHyuJNsZVLVzDzteKmvvO9m2IRHT3Dj+DKaiwM
he2JOi6gLVFsOCHIDLUTERyzS7/E0oFdURCdrsZg1ciSG7upWOspbwLpHrlvju78+Ec8ilPJQVYP
5nSViqd72PO73Zj8KDyGchgEuwx4bv4KQ5L9iqzk9mdBjbuOJYDGqirsGBpuO1BZGd+yWSr7NRSc
t0WxrM3260MCG+JSlR4feqyuZGNLZPTQh7lFEuGzORdgkp+vVrLC6gZodgtg/BNAuouzWpz7bqom
SjXWiK7R0R6QxbANFmAMy4nAhClgjXvyilYimSxPZEdehid9aiRTzPy8lXgQVo9u5+0qSslUy5Fr
KNGsqftgiR7Hd6NsFQ0lUAmmL16DTWpsrg0e4w8xqf222Wn6eyWHZWYHHBeo9Ct0FXZDG4ptt7qQ
W8JUhyL7jBs1XghHYTfMCBnPOFfDS028iryEVepq6Hr+6VYR0QDwAOLlr7DwpeoCIliEHsF6OfvT
E4+WNrpC0dzpPUNzCgCY6lUP4oaJu7c/bh2akVQXsQji9CDFOqFCjvrvsWAzuSpkMGKKItyg9F4h
NN5tYtl1I8S7DHUeo3P7P3tgB4FLiqHIRjiM5674dCFXJubWpXUjHpUrlRQ1R7xkH2djUfZp+GiM
Wqh7Z/ecfE4H03QnYjUWcEEtAbs0HmrWuzERtb6bTaq3usF60vYNwqyXI8TROuOvpulHL0KeOLwl
CgysNnWlbS7FTb1wD8u54uiMR7adW5tEvbPTcQAKnYBqSqigRQXrb1oAGJlRM93Mulxo8B4CHKXX
GAMLZnfhmuOJe4FcSqpbwg3NK7bEaY9XUXeyDT5FyBurVVJ1z6XqQvW8F2M5MPnSAvQkZEIb+nUm
gHZGd1rAeYsf7FgyaVs0119guPS3s/Y15iEL892kSB2VaXyCtJC1lEZIqpnjDux59spu+LKqxz4B
YE1wtGshZHlJaVhbQwRVUCPX1PsTd1BjTZux6pRTbIEySE7ooBl4tZRlF3M03m59GkrioAr4BEzF
1eX3izpWogIRnI1/Vm2jkW9BQ8mTJQybVYReM4OgR1pmiRr4c3cdLX554p5GlU0s4izS+4RzturO
QPkv6bPUQMkN/aMXac37eOa/yG1MJGUTTlWsXSFvkVg24ohVDRcIgFc/6LPwyFOUPR2X/5GQzbqV
tMjszpnI7Zr8tav1MHegCpKIJAEO78yeZtE8BP3tNbCMtht6Lua4qCRiAEXf5xX2P/VGdHpD9Lwx
NMPX3HpSAZBQFbjWVOd9yLeliZOrRHODIlStr9LGQUgBlTalQvOtS/6q51Y9NybbhBiLCkfa1pzZ
26W1edfsvWmDh3FCu6S00iWEuC3VkBj8BuJ01M7eod0ZaFmqIk6yuSRHGKW7899A4WUb4iXRb801
YyvmlZD2OchHBZibB5MlefWiq6AwOG+AnfSaSmrPdvEb3qKkIsLpA0aweejLPnTHNazFLrr59Ei5
iCdtY5Mxn+NI06hDJy+7IpO3gBSLWjfwaUntmPmVySuHgQTUn7wPIk/kEN7F85/1E9e39QcHPOqP
z0Cj0xJAUHaZVX3lUda1FLsFoKx87cniqO91ztFHibNnzIsSCBuM4YecmZyyljQ80QrYDlhzYncM
MrNpvOCHcYxuNnWTNd+K1azb0wk/grrBare17+la9jOmIPGmqCUFpMbjURjZTjDCqiE676G/arXN
h98BhgxK6P1s8lvv7oX2/iQrBD6PdwxhmQKuVYhs7AUjtFsRh4RqsoR1CnylisjLZARBK3QH+IAu
j0CM0zxpXkT8w3JNvo0l7fLO5K6eJOqIAidXqAkms/DSslWCuwDANJoiaibqKHVeFmLhxOA2kyf6
to3f7iKSsieSsE9EMGnrqW1XeAL74M1Yw6nnKBoNULWBngkbiMu2KYPld2ulvGUlZaomeMvjdDdv
60QKg6B9Fw6HiVuAHZ24r3a8gUlSYmLDYb9S3r80kM8AACoQHqCoQzSnY4p7ptk6tkQ/lBHH8mBg
MttBzSVVKjuTaq+p8u8BQwporGlRzYlr8fVu4b7gur3sgJiJj3e2fToSd2ThA5sfOmjwNUX0sHzN
MK5dJQHWmmuRLnN3X4b8+TmfStLa/is6vYzW20jaoVZT0t/f431xagW/8vRCyYidwBqoZIm6Y1Qd
Zi20TOA8903xQfZvuo0FRD/4uklrI4+kVTu7IvAKM8yUWSIahrIg9UPr9e7uGRpWtV4xp1gQEZUE
dVT/a7/aqILBZz+m0UUYnktCNzJPwfKgC+GhwwixKJTse9km2YvVj5AyHWU/N4ykBu4pR5CU9aIc
aFa4uMMz7rNVqaznW43smTxY4x8CI8iG7fbKEMbhgf9e8IlW8dq/8XpmfggwvbO84yiLXBa3zUAm
Emr6jQtxGjRSR4bU2hbAvK14kB5hTflkRYXMxQ8fS+zu9D5h1DMWp22LyLn0x9MnUoMqf1nx+vQy
Y930cdqUXL+SD3sYnsGFiQcYGeqP+eMZXpit/ErRAxE7DkuesLUsjBrHitJ7ZAh9uhmKtcizTQhW
JGQ8thOwAAOyw25CegFaxML7WRRO66rdBZs1HQLK3GZ7qmMvZI+yTSe2XtXBZpCsRIaVavqkemuC
Yj+YxSmyQ04v0P9y7vPunpCOZEwEy0D8TyVTHfsjpe8mw9JodyPLwKPqi7o5xBE5M6GOY5r/15yv
ZtER1P0e1rCKOu+4SJpIOmvf3bJ7uUKKIU8POudOR5h6yuHGz6hZ+w+ElBr0b3m7lbkLJh8Ghnet
1EE5wzhVI91HOLTGAwWLDv0tdmld5pDhg9Vcj+gJzP7/uLJEHsT4IjyYWt4/4bRkfBOITP5hTRv8
OA1HejO4VWquT7OK/I4HORgp31QdSlO8sOR7zDKXADKjNEta6F5Tb3CN1KVQPiSHYT6Tgn2OOLyU
xYfxk0FGQ/MdDZ1cpDm4loe66aHcj1P83NCRc5P4A9jsxRYp0aeYhg0qH7dkAJTKQK9uMBfAkka1
k9clW1alO7IYBAO7pu8PKoEX7FB9TFGhR/FLsie2A9irEbo+on+aet4AzenKQe/BeEmixaOXfQyg
waXzA8NxKIn03Y/ZQvzSLBPMko4g2UkQt2NipzvPRdgy7uygClgjNn6pGLjhC8Wydq71AIOYU01F
3eaQ7FmiQQdALFBrjZRl3hJnacjPIYqNOnjGP9TMRwAHnq9htG4cgjBRBWjDHnlE+yxzNOLVddpn
IKGwvyt2UbfBhMFq4qEfJO6ZIBE7zHCb+e/gpBBR14b0uB54HxZlHPumS+86NZn/xSvOYf+lXuDM
GnyAY4alrbkuj3uWvOWzM37ZXWmIuXcq0sfSXlISSuWrPJ/SgqhxVkzdWB3JvoibaxVB83MPIaN/
M0NEnXL+2zp6LC4khPiVBiH0Wh4CKqwzicr50T9JYAXGbJH3EtGxZS+mQ4hzuNncblgIt5kyMzla
96Ex+VhEAZLqzZNlEnLO9ISkt93vA/N3Mwtif8kRpHzxc5+xouc7tHcIHFCLQTIhgntkURAMR+5v
Oe4klF2zV3rPYO/Q2n7tAylBEUHS7imCgEdyavrC66TcoZ7+5fPTp0UDRyRVbh4Sk8jNHVUqguvG
fwaIQsCjmlripJmtBAZ1+aTefkYLMMG6llEVAce4l/GyAHNecfX1FGGX+obATMyUXvrtvjAKulwY
IXnta7he/3gMsA25BVKrPVuCGvcDDKUP678JAGvwOOx49t3GLfJaBywhCw55ecDOocAJSS+3qr6u
4cQm2xRD2bjxdUXXVGol28aFsD6+TwOJx2gMIVloA7jUu9/UB8vtr1HRIRwxChoU4a5aSMOLluXx
4EUCnsxPZbqEJ1sMi0eUsfQZ1wBu1NoetM+21zNuV8rojiokEaw7KUIedkpzaUo4UIMMSW8BIUJL
CmNiq5zC2bYqdEJu3o+Q4L7LMRz8MEyyFzCOQWSYv0SaTASbAVSNv4e+eNNLwBmgpVFW4STIV0g1
i4+0kWVNZ+oR3Fo10zfU+EATqln/00OPS8ciLoRXVsogQiH6DR8XhpFmGidcvmSDRgVL8xwyEsfY
NEaJsXuhUlF8UKGQ6uh3v46QnMfHhL5GZRMQkD6WdstKBM7SHlfmDQTkFWdH30LK5x1zSQm4xKh/
oGi/A8NUuPDddWQhCoxeNkg45XPkdruxiJVrH5mJCjf1aeD63mWFDNOLXQOTCUmXbeLJFoe/oQfN
qMjLYlkWW1K/YwQkqwtCzc7z7scHDrJS3CcHCCQJg+s5UNh8YRwTwCfDQ5wnnwJPVSX+afUhd98E
DoW2WMHUoDK79JYOjK8FIae+V/urtg/ZDaJdpY+wFag6Of/1Gq3rmpjFHjQGTijelulIUE2fXURQ
G0amkpeZ7oN/K1LbEqs8JqC1yedjAO1HfXbZhwkPtn0NfvbvxzvwKlzT6mhFM6Hf2mwvFlm0iu4M
0B+kXQp7vtOJ2ICR8gG2ifPHgJ5BD0+z6uWv+RxLkvntwe9vZrXKLPbpE3E9ApZfrhWIgjJHJIfq
gXWsKETJJdEXtD/ww+TY+n78UMiSp9/ifi2VB2nVLHlQm1AoT5QZQhMY05lwt2Euls8Aq/Gz0gfu
xPXM4aabAL51R1axzcVe5o2WbrEtul1mOGq9cvFZyReLI2tNhIyc6uiUzTbOn554jwidcYljEwj9
de0wnpXdfFzjj3wza4eQUH/31TKamWEB52iItzdnogap9u0QpRa6AD8/PQ2Ju48xudZO8OoZWC3Y
EsA78/o3BUjZe6XypBKi9pg9rekKEUbmdNn+URtG3/6j/toVSLakzs9aXB3RrwMKWj0al5A4JLCB
PPoueBgJWnxhGra/+2oZXtCd3xRbQkJFZK5qHl20UeCOHsu3WhlyQqRQsY/ublgU0RlpvxMKbv49
3tDB08WVeefm0bSFrzhsOrdAUlXgck1+1q8xA7Np8sn2ANsicPi9vUu3S4+TX9UqTSls/Dgs1+c3
j8ldqVD8oUi51Es2tKnU3CcIZQJsILvwqG1aXAIFshpTkq0s4S3f9E6AarIIMOb4Zp2nqKK4aD9A
0QHCrgnxYeSC0FR0zIOh2N8cD2XP8kXP0v0T2YkgWVCxUukd51Qtq3aFLUPlE9wqPNLWKslGcabX
1WhMd2I0lOON6Ek1LIlrsCmGEI36RU6c6t+815pkgA2kP3n0Ske9SjkAMamgGTFP4Tlt6axf4f3g
6Okoft38JZwXG07ZHOiT8SnfoXwzFqnlcj6nrAkRUvisfwKZtyB+ONfiJYiEdovcIJr7HTpPReWT
UsLikZdBoNbSOcmBz/Up3iEe47DDhP2v8xskGUXnjU7CMajoQdFkd7WH3cSvyW5ZekIZ8ryPaZ1D
sTypU1EdKi7ZTz+yyRzaKl8AuX9Or2ZTcvVjzTw95ChW/QL9LZh5BLrDeuJ5k7sVpMc/8koOz8g3
1H39itBannsV3oHSB9TIrnl130wZdp1YSPtwPejES9KjwQJSc1UEK3CQmasMXP/8wQIuBUB4wCOq
4Qda99X+XhNsaNXNCzG9ScLKfi89NqkfRn3tTm+blOsvr0UBIGM9n/SeV0HJtVJ1mv9/a6k32h51
axvQdBW+gNdNrr9hNytmfiucapYQwW3k17iAqQ8lkUZ4AGND3wOTcjaeEY4BhMqibxKLBEF3yc4U
g3pkET7Vbw6I0D9u9cBks2wsRxTXM8etlfr3lb063m5BiE/wIGqC5OsrB9R4OjiQtyoD1phkIr/I
VVRTO3BBKJainvwBPw2Mor8f385W9q7bn+ScRfI83I9XlK/j2uFB2i/5MQSsAV0mJdmQQp1r/rNu
VFz1btMM5xbHu0xGgwLqN5L+6g/poRuK9pSiFZjCWEbTWFCutLLWJBhEo+l2M5NRc7s52HPiYgDs
/O0HNIsvo2PTHYtwNDygWpY8ccX4Wzn5A7yxpyJcUshhaRFVx3G3YXjKFZxa2OdOX8M1AlLr5uqb
NJWeTFIhgfOr6yk688GCHHFtlv2oJNF+CfRBzQJRmJ19d+JOvEzbpOmnnHFHOI4dr39UPQTMwKZ0
DZ7FMHPu3Q0LSVVvRi3T+Hsk3+HHCK3fQC7HkYJ0mhGvSUS4gZm3rm/Kx9LkgcnZ73CwRcIhAXrs
lIY52RZKjcS5daBYLiQocvqj229AyL7Kqnsne4mssq6+i/ys8X3GEOEQ1/Q155dMFQDFrpkJ8Pu8
z6WcC+97VcrLhcZoUnMRyb1pdbu2LwT3JpjEKS9Ip3M05gdaDWn6J3eoiglh4qmdkD1mR+7R5nfp
Td4lOcnOp+pN2sZxmTOoTBEHNvt2BsYXzMqYbp5vhNFeo3NouS2xCx2KKbj4ZBdUwaER2fY62fa1
m5pSF2s64yNa8+zoDVry+/rfAmN0TyJQcnquJnhJfwQniDX+ncyhUnFQ3BsQO70AruOcj/xrO0xT
y/xdkmHwZQCFEB4EPXRmFj2HsfFhOJvcdUTgA2K4gYbl9DPTC3xflnq/EcIMFmrNbx1dZRTf5rCJ
AbZw9c8xhFI+LW8ybD9jkhKRjfYT5b8k0wrMIC0rlMqSQ5K9cNixFcEO59twldj5dPpgb/NFgEYS
fFGtNReuEtdw+pP24jwSXePZQ1xZT24hqBk2FAufYSDGRHW5pgLB7DBYsyebV6TNBJ3OR6gXtL3x
+S94f6VSgjL4qgyH9dPesF5zJ3OYGjvYigc6d2TQy7lUbd4Be36opNlMg+KH+ga4odoyFpN0PTN9
7MjT/B41bqDUyyc+gwNDN6tGh4ip8/o2RePIiur3Gm0DiwgFcPZNvCGPkicYSljcV+Ddd5iMKiU5
X6goLbTrzBBW3R+Ts/LKVvMiUsJSgVul+S1pDZwBU9rES+R/EBbvg8rBSjcEwfjdJd4zuKZSA2uT
z0xTBt68tQlxpc0Ft5pbZQdsr4d4NZQDc1Wy2cNqjJRiym6vxe0Q9VIRTjrCeo5OF/baWh+AU7Es
RQZAYI6TLxEXo16/22/p30tpC572FnDGhJjjuq8fY2RJtCRjRpnA7v5L3ZrUnU+2Fqo+d1CKaXvP
ej+q6vW0rNjFBkXGletqLoenCjxmU22qIVia2cANahVTxUyyfkrLZiA3SZ5rpPd2dx7l31qv3T3K
FVHz1Ge5PWPM5L7lOG3PM/DgvLVjYe46xhlIPh2dQ3AHaXlzXg/7xjd+7czABLUsMZ6lSwVQIVsO
YpVSbiC2BsS9r4qu3i2/fW3gDjatxOP6q6TLOznN9/92INietaDH7pTPAKnrLLwceeQsSrgLmmef
oDO/atTuTJka8rt5w54Z24JcR9u8VihIiggimcA/XB7uZQypdi3EUpqfpOcKphKEIkdbJjLUU91/
+089UpL6SBoZWBaMAI/0WUCWVS3nH3HjroAp5fpktvR/eQXFgXAx+yVnZuueY/Ac0RAGPRgilRlV
gMaMxn+FIZ+O/8kppunI2n0x2kLb9b+QYPiQKqFNIEFt327rpCaTvVW+v3xn4VocJRT8DI4ANkZM
Np9isaffSYPvpdNgj6c1y99Q+bBezvkSOY7u/yuVBxm0mL9CpDU4SQXGRaLABkiYel1wNZzMKLby
o2wr1qetPS7aK+evDnYr9Y/N7N2LMKg4MW0VW4PhsX8rUJRvDOIJOh7QV3cCAFB2x9alpX+ZPmSJ
daonUZVIbowSvouRQK/1a32ucGBIYKiNTS0wVl6oyAhPyWYrNiFYyHb+V24lI7rCvsdzchsfpUS3
VBvJzlZdveB88f7J0UZSozWQNEln9D3RyvsClSpg+2gXT26nlen+f1xdHHyfNnGrmkBe1yutaG+v
axiTr0k9bLIULJU2HoP71Njrq1QyOXQsaruZ5V0XVH+gC/RY4cVDzB+aI1M4+IdAwoHbK88CjXGz
nBqwY034Iy4J49aNEoDKcyT9tZu5fwDZPPx2xo7drqEejDQu1n2ZGa/QYXREsyo+2KjrjEbsoD2/
XGYLGa6FKNOKjHHhkumMCeSL0I1LZU/Fensv7JRi4TL4bl80ak04kBy/JAyq1K90pFSCgmayREd0
dT5MrrB0slcI4yFtjbPAa4os0AWJczW9nGJ4zx8hHAG6Lx/cDEAjBGc+6zsJpguk5xDiAJQmIi1c
34jqs+tHb/JtlHCYU7Y9+C+xlP1H0TjWVlWkZB89345XdJl3zu9MuyDHY8VcMAKkniExmI1lb4kH
ia5xDlkTVFQuzWPZQMlMtz6kdFFHhsCatxurt96N2cNjzHW8f5/amhN5X2NlEQZExXx7Na0QIOMU
geNk8wFGE0UgWw2nlBqDqmUoeOkY4NPUcjPaqIGT7KGdwHsQzblQn5xJKRKx8UnueKNwXuh5rREU
wY0JgDL2XszI3BKusvxgKabFwlZoOMJ/jItyGebF8otRKh0R5f9wjW91TmLQULuy/cF+471ib5r1
gEogkrSNr4BesSKpM93zI+xrytwK3kj7kR9FtdO8tp8rOThKVQ8MWpElaTB/ep7foFIEidxuoXll
TkKQTjMVwBA4p8/bRxDLM6Q8s5sNSpOYTdFfuX+uQwRtk3VFMighsehWAiAPDf3IYRyw+t2eU8NS
ThoK90Cs5YAriEVa5Dg9yzVCAPtZm0KF1P9pT+lvxnanSGTs2Y8zlRxRUJMkOU4BRUdWVeF45tbv
FQv4w2c6cl71ExBapghFwT3WZUEtlzJQq6+kI/+FiojxPG50aNuZAuScu0w2+DOIAgji2Iv6ivQ3
FuL9ih9Hfg4cBX3fjuus6Gz1Ip0eE1J8cJjn4tOzOyXSopSlsmN+FyjMafh+MkYHy/mLDRYU7rCG
mXz2kxdrHatJYbE4HqwW9jCh6fP7nFbwY4+eTtPWQo8zMgpVP3iceMYsIdSa53d7GNaPuR6csV0i
hUP9cySWESonLIrZKSMPfT3f0VZQjX7DAzKCC/GpQOO1iUkIb9eEdzzIIiEUc7+6e4zNdJUv/M+f
bmM01Qn80dVoBDYyj169k15EaTl5F88fPrjKPVFFQsyERpdNKiUP6KubZRtiPd1MoeRVOJ4MZYm7
isfMmyVBBfocyq0cuA+2B7G9MgWPh6Ir3mCvak+pz9DmsVPHMbeeVaO8CCpcrT+oOFJCNLL4K49i
QoszmHlXbPxIvq8W7wiI9DD2yqRx1uleIctN9sq0BwGsifp4i7XdK1R2nte07FDLae4zZJWuuFMA
SvpXQSMrY8n9nnDGQT7Y9At7SeYi90/LqcLrwebCT+WNj2Lv+m7vkH/uxKQu89fNnmMXljsfJgP7
fKbeeS9qkZZ98aEna5jBP1edn7VAOcRwKKLunxob3ZilT1/uBwfeJBdeE12iZd50WCwjJcnH9wbI
rdY87U62u/Yww+Dl1fVsXRgsmcMELcGUNFxQBX1aa09dJlT8xrHC3dWSdkytjs9TejcfeHSUEnmR
gjNprr8SyV3EH3c/Z/UUmejZ9E/nvUZAg7NgKghj11SWCynRKmj0Q5RqaLHvP43knVkKOkFtLUAb
4TvrTNh/mkmbi9kfDitv4D2OBQGdfCMLx/1Nkn/JnIW9etLMGNliVB4ynuo1Wwq/dJP2zXoYLbIu
GQKpjjGx7XZxnz4Lcym2j6fBZy6xx+UYiOr2WZjVZD9s/48Zl4/q2RE7yKcEjX57dfOdOJCLwILg
kbCwVXZ/GVZInps5fppTTBAhr5k3cLDrQtFlRrWe07oVkvS/VcfmjxOcSo1HuLh94nzYG/MT/qGe
710A7gi3Kh8Tl8kiMobLWVh/d3A8jE9Tj7VoxLWvnKH/lDt/qRkqkb3Wg57SSpNmeyFIJYkneRWx
DwYfGdzNmaaOmixR4s1N9nt/II3FJAxjK4OtgFeEAoRBSPTgyC4ZKHBQc97cPNPHhtH5IjrYvs/Z
43wrSmxYEdUOIsrYyqbmojY3o1VT2smJcrhxvZxXLFfQKlp7JsXzv/KeNvlhK6OL/AfpDhUw5Zfa
JcNSyP0E7T9oC6DrMcTWq8k9tv7XRStoT0PpgN5ycYj9MG2rqZ7BGv4d38hmsf5/v8fnr+6nFMx5
XNmTVyN337bmwEODhQuFk0t++KaeQuifgHpHAgNS2slUxHANrg2HDuOXcyNCOFSRYN5uznZ4Y5mh
aJwm6dxbBEL+zKgnv7+KoH0aLoEOtT/07AdNt9Ko7B0499QYOnHAoKPLglBnOwUaXDGntMHB+emU
Jd+tPrfK8dE4RD3GXFx40rhPGfMbL3GWexrlY/5hKL+KGClKawTs2bPxkF27FmSZ8WaR5WKm8LH9
ZvupkxHmTpaNNAIuFwTa5RhLZrPHnAGl5sc4OxQG8PFp4ENRKIhf0zwUOJL/nTu1+dYaOEWQQmiN
hx3SeLFFn1SDV8PiGKb0TrKrIXReFatSRFhNwMLK5XHkbRUh0bdAsDeU7BMtms8e9Ko/FKclb0pF
0ncxdF7+As58kj/sJgceewP1OYAbO6vfbsSGeEdgvW194Z/Z0zj6+AMsI1hfhIcGBnX7iXZKmGDU
zjYlyN/OAq2luwFoVtqlHb569Y1gORISenbAjoPgrUT7QKp1kPwPs1nQ3s3lT/eezfp4FSVuBCzo
KlZ+WxBwiC5Qkalj1Y5P0O65tjJzM94Qbr4MKhsnPctVa0VTbpxuL6v1Kczl4IOR2rmgwqEs7Awr
13JnvDGKeVh6gG+ISpFpyG9akwHilukkUrTZzgKJkHqnxb+DefNJnOIKnIzJSChChhDsZ7Z1vM4y
VayghFybm5uFriyJxhEQSqaFTjUCqHZH4QvonqWnsoZ4kIgq+05/W5hp3NMCXv2Fxg2YiXCBJ66d
VWJXMZDU4NEFFAsKX+lefZ3IsBeuUQxQ5T6RgeIrDHKe978lEBSBle3HfH5/ozHWHaYYOKK9jKQn
2O2f3NQ9l9v5my6sXDEMuod3YMm9IlkMCU5vyMsn9W5gkdmLlhPdwQcX08JpLEPuM1tmcEeAoEBr
TyZbAIgc4rwY6WBi8CVK98lkDmwrfL7jLgir8s5WG0urPY5OkRe0vOWf6qL2A2OyYJaSPkeKzpmi
HpFVHAzWqtBixNf69nPXKt03Bd+JccvqzrZOraJpzGCkjK29yCm8lCUe9U6EADiXkBkZ3lY3Jxl1
CQsSw5jIOf50wY4WjBKe8rH2vcrYLKK6dC4+Uc2MxQcP7c4IKrs/G6SHLkPC1mQtdC/gzR4aZ09T
ryknBaujRAseRnB/IuRrbJZdvG5ivfqYP0igYxexgYROZqCom1f72U4ZRgbHkpfI1LNfYB8qMpsc
fJY8iGBa/J3v1XmTlwkMAQZ+pWEAGD+fSg3Xs45LwtHVfqFBYGm7Ug6nQFaUIf2s6NQffDExpSej
EGlrQT5jBA9JjgNYkGDQ7rV0v0hOUsZxmgTokL5xDEAXxmNx108MLHKVRlYjeFs6V2CoaLcYisBQ
yO7RXRYd6xZTlE6YePQLW2CqrMDXdKRwBgsW/jZE3SbBHxUiMGMV0c8aiUjpqs2X147qHnF1dbSf
fscjzju5AbNI/pe/UHZOI0e2fY9ZgU99Wmb41S2Al0OlzRbOOzIbrP5IB5LqlDqldMOZKLA5D6wS
JAUukNGLdDY6TzkftK2O0qGrK3JCAOFKsZ9wOgwthQcQK32Lijec4bwgfO4Sxd7hdxVsqFFbOQtR
+dWeeFngLK8gFBk1HcZEmZ09U71EedwTq9mt0j3zu9qSwHQKsJ1hc+oeO891FNDTKHuDUaZ/qoVw
Twox6CogrehTlAJfiMHbKojD52lXRfVH8GIzlG+Q97ka/1YBZZ34sGh2viHKdFiC5G/4PoA7Ohsm
eHl3SclBPpHUZ28u1g0YS1IJQ8LQ8A3j95J3VNQlTJjgvcHp7UfxoeVgY6DUTiXZdy6GmquBQIi8
4kXJHGN8zrTghGFRW6DgfOmnhqwAFFUm+Lhgv6Ntg11dLH5wdz+p5kgZlCuVABBGVxwyRtTEjHOC
g1AR+lRL0BbXU7QtIYBg+LlmkqUtP7BE7TiTmhAcecpKMcm1FUS5Bw8u/C9Zh+6Jqscj+3F56bgN
WPvHeJIxRvkqRc+7p3XasgB9sZuuQvYI6r2KWybMV1bgl3d7OqdRsed/fFmNaCySJ1SPY90GyCyL
cAHLOEf/HzMEN576vsnEd5jZ0FyUcdb74ODqMTvh13eEgJZEnSk10v1V3fG9tqQBrp1AuNNRrnZx
JaEyevZrqroIFEOl9is6dHlGwOXyb9szQ8Cyc+CthLZUzamwwjJTWZkGEsZVq+9QjkIQ2ZOK1kyN
PFjt6EDzf53+jLwA5MOaSlcG+a+XUXRWfovoHa9TmGfyVMUyKFCYEGlL8es2eZGgs6n70uqd6zji
BgaXBdAZGUrLWxE58JPqrxauBD/Ohqb+TFy0gnzSABE/7mudha++5EzTMFy1kr7pjB2bQFHIB+p3
CrIb91g0iUEF4oFRA3xjPr7ipgxctoBFvBtp4R4wk9IKcePX560ro/4gdfyZZtHR8zOhDS0AhU7i
t+y8psCH3rK8MwksrAx9TSR7hdnfcGZoazyWzH2Auwy/lDuI8lae0WNaPqGgGfRzwzxoiyeSYHhf
9wXrEnRNVmmfKbbvWN9B7JPsQxygfBKviCBGmPRgDMEHTy2qxmaCRcrXHNCEpXK00e/RyzQFwM6F
NS6l5CFR5OUN2S2Kt7k1TzZJU7w9rFSh4zY8WbpsqLB3SkRzjUHF8jkmM6bnbYadaXBHZ/luZ9Du
t5GCtA9ymQ4zsyjAfYriqnLGrhY3LD+cJOntX81cCqzaZvBns64bSIso6bVO2oPAivMktuZwynJs
pNf3HFjeun6fIPKED8OxvWIAGuniY/0YaUzOtqP2QkhPzi1jpPMb9zrzRfiJgXMSa1oqW+sZjei9
YUEJW1uENVsAI4cllVQJsy1n/WURQEGZmuH2A6cPZTwNrSlYb3h3XAwoT4wk0AlxZb6TXBzH/0Im
aMeFi3crBgLqZHbyXDDZGID6VFQJNAmNlfBHrtqtXTO9cyITOyAVHIlBz2PBiwC4PaGQQR8Cfku2
vwER79m9N1pZfcPNKac3iJCLBUEY6bSXCZOa9cY33mTm3bezAlDx9N5jpjC+esh0M6ztK4jkCG5V
83ToEXnM/p8njG4jKoMr0VQlCsZYVZEYtveU+hvdJtps5xd2Mf2K1pyqFg/rzQ/3LnkAAIT7i4Rk
0lYvBuH0IJLUiMRtrCm+lnj3QW19Iifdd8WKYBFOHcnoM7zfROj5qW3XoeMWzbXuATSSeovkljV5
+7PE6JZ7xJTmKRJ5lYJFQcI0OGmtKWeG5LDFK0sazAL6Cv/ADuvsRV/ZhMboLkEeuR0I2E0v9Jnz
+1MhmWaVRDIsFIXOIZ01RhLycgG/oJKfiCgAETLuPM2KQCWFMwTvIE5bsopFQKE2gs4YdlcXJT7j
WgJ9doPRLjMLM+PfPwWPCcH2cFaTIfzDMHV4uE92p6YjwS0o0qODlm5obvsqLfo8T3oiS5h3FhR+
7pWqDzA1HW2Ja2wKR2Ea8xlqIAWgiiMiCGjCyhUh4gXOa0hf2vxwR51/Xpze4ecLwwkclAYZzkCX
0vHxN4fecdieby5UwNnIaelmXTfA99sjN0Dx3OuXtXgBWb/8WWiEZNm6xW6/aLxXZCFFbIjeSdvM
FqIo4/patlt8vpIi0S8viiOt+Wmnmj+2qx1O+nV8/QclFjrfK+kuSIG/CU/kl5LnpDd4371uJ4pr
jKzb1VOQjBOCmB+TnH39/tvft5U0OtTY3vcHqLQzm/F3A7sc8aTbQCywatm7TbJfXkoBNOHLxrmx
ilbxXESE19BZ+8fzcsu1/j0OA8jMH39bRMAi9c0ge+5ks042eamtc4F9qWiih4DS/1m0pEI6LxEI
KkExorlTAkeIJinToFUoqb7W2NFxREIk4VgfPG4NO7RVQhkthTvg31w6HYUzU9VUJ4Hf7RiiU/e6
FQf5JdohADL+pRYsoPkUD9XiHl0vXp+TlsKATFZ+8wea012oVa3rq6KB8GXcRiVdS1QuUGG8q4y4
9ci5mbRy/Z/lN9oWwNHp1rqp85pcj4o358hP/nXeefjiIhUKUXx4Jc2G7Ud53kZ1ldGCjtigiZ2i
8hVogYZsqQ3tcO6rEXnP16berAo/5AQA3AYqzKVybPHsl4SxMGdlBlNS+/KpEa73NMoqp8gLnkwA
URvqSDtLhqyJXt8z78SPxwOn/ScNKqypZkHt/J1QGgrPfhspivwUnEfQZtw+4ZDm6TkirW+Lc0rX
FmrijOlsgXIg48Vwp6rpCslk1WAHp86d9pCeek9LI6DurDgDqS7E0Wr1ZAreGI8UdZtY2tx+knfs
ejJb0gBmcfZ0/6Rq2nPWPC1aGoD/j16KeGDDWcZueTkd5uQj2x07Du3Z4WGKD2WqDnVD+JhaEnIz
hvuZEmI7otz8KtrNdE5hu9V9WMDMtQ3ezMC717NbTtO0Lx36s14NWuX/mMdPE+sjEtA/bKoV2ed9
UU7mNvj7EZ8fdH5HuddAU/CNeKcWNY7XHqWQed26LaklwwRBuNxwkn5lePSBxe7GIHtpLCnL9U4H
Xx/jhtub11fLAz2q/Ckz4h60AwRcSKOtaZfzL9UawylI6u7IhGBSaRE+SHfDoGrc0CR0VVQ0MFXS
//Rl/5hyjucavXQvbGYCXb5iphcDqJ5q8vn+84cLHSwKL9ll5xdjToH+9i9urdnVBmN/nJP6pTrM
tBF7gZjxLJmvOIbc7F3AeLF5Uq0GfUWPDGGKGqZBiFoR3u7t7yJeEkG6ej6e1TRH98mQvX32tz/F
3c/wacI4wnDu0PVae4ku6JD21ylennabD2LncCgnIqqylMUfi9XY2x/lF0oyLaaz8S41bF9KS0xw
CW88qPzb1oqnjVADva4/M3HW427BJH0/7sXNpsIr2HCfWT7A8KpEb5PopPjwVMEowrG42jpLmv9x
C8J92+GEV0bXKaovinB3TWSa66mVprM/VHjEushFbq6ToSmLEjouvU2fIWg5KyOVQBbUF05of2Zo
rWmWLnFClsU/E5Mn7phVYj8O3chLobP6LntJBapk6IoUqfOGNG+b6GKgZUVRGSxofy2NQRsgbBAM
dg3RZf8DZT4K+seYw+r6pX2HdQWPCl4Xp541n57ZRD7sMgq8fQjja0+fdkj0ECj5hVrjqKvCC+rb
tH5VijkSdkkK6u869ySOhMxjoKB1Z0LCKb0SmsnlO4kbwQ8ank0kmOvMiCaNLyMOQ7sWgo7DvY3F
Av//Jj30sSzt4lUsxYc7zYIETYmLBK//w4tWSQvv3uGfyKXKs/X7xdNqBMbOCLz+Pas2zZJ9aCPR
5LDq+eqbmgidnZPS1/rygiQnGqdg6AITw8x9TKcO5Oy+qVz0TZCxATJbCnDU0nKneaao/5PlJymc
SD8n5m3or08QXvmlE8Uecj+Tv0b6NxhmXDs5TrtdIojtzhSf83SU4v7wBwpcb5dPvAyoJ++WoFf1
bEhNvtt92SNkeyOSzoqJ3edEkY9HSJAFXxLdJByJTiIWmIfgUzL+L1BVBtA2yZlqw+Kme8pZIdg2
C1GCTiwPwqAB3VMrdce+3cUDNaFNNeqVhf9zr5z3WNvts2hUszpsjKWin9W4DtMakUNDCVbZtwWL
hieyNN4YzAyTubdyC/AbSrQk0eA8+X/LbDewtvTbB56LuvS1tJJfI58eOQZfN1Ol8WEo/QDML/WT
KIEbt6cN2Tyk3F2uCj2Hi3R7uKorKSRsCe+jBSqKMDiYNdlaA7Dhuv9SDi53FozjFzhlJjUwEMqi
sXrsS1Sdxxp2L+zQVSNPejdnJscO5m2eP+eZ/hieWqSr7CQlHpq4ykJ7Ogz1cLTJu4m3hwlfcg2X
kZ9Bl6GZGijQfIxi5ymFRrCeSvPo0lju4Kl9LpMQF22fwUganA8MZNtSRENHao/cHnFhqMpmJ9hP
vvsJkcZrc9ZKKZLOSTJsIIOWG6ltmZYfqzWYw9/trVJmgCcu5pvc1LvF3nVAfauOwvTYyuX4peUO
PudrcBwGlrlP0JKYrCmTXHj/cwYQKASpVdNr8sJ3/CKs+aPRDMSA0eQM7hGDGdMTIH56gcXeYBFy
IYg+k+NwB1ghrOBGVvy1bextOmj4vHKL6Scj5pxpts73Kz5XjFKGWOGQjJmQ/yyNaDexUYXtidJw
Cl2+J+w7Gp2jBIZDHQ8xa1m/y/xJTlMYoREZFSrlf1lpk4cYsQs3dG5Uo1cbbtqKl0RFvuZaTz/t
zxQA+JB8OGo3eC9KrPVjD1wJEOvz/AjJj2/EN8x0LJROpwP9W9BRnMxZAwFqdXTBya/iogxZ2N45
kK6inWRyPodvneVZtFtAKFpV7DyfLQHtSn/HBF7t6/uv6XgJWpw31fbPPRyqBSOHigixZrhk/2fQ
OZ8E4mstLsE75Zp50wAKSdG5p0A3sCN6TkfiyC3jepPzgpChdsAlQETDdi1gWDgp+XwJbRIotqCs
EJfotNdU62moC9AWqhyBG3U3GnhHSkl9vBqRtxgDjynuD4dAr0JUbOT9siTarOJeyCkC6QjxudSX
s83eDzA3j2eaXJJgh3jELHmt2M2M0yEz5FjyzIH6BQqgsuy0GCQPn5Kb9526RD33+lP1NqKKeBh0
aROYlU6ZMalPyLgUELrwb0TXZSzfjRBQe+ZV7rM1V7rtdq/HonP+M8m3QITdWdAONdtvVmBDI5rM
eRzyQIxERPZKlsdZgmiwsDoVMjlNm7uYR4rk3LjvlXgpWg6r3hHiA8QKr+oNMgY2j+OCIFEqTVCp
nuyMgvtvSGcD/3mv8CD2KAEcjaKO3Z5O9UtS1JoHgVnwP6lWgBonYPd+CObiRwlF8KeaE3cIPfBG
NTuzCBS3Ahql3fzu9Snmulw+ZR2iuK8s2HPOmNB5DInZ3bN9xrkZap8dwavunjGnDuuMHTKsIH/q
R8kTgnZbPsme0d0j4IBnJU+5qs6F+EBhMxOZBSP1UCLFnXv4lenPYmrRr9D1n3iI5SaWMj+orZ99
u6yqIs0pgp7KUJJKHnm+Jr1fEzC1jt05YzTs46eRRT5qHcHiFWJb8YJ7SuyYwr3ml9pdKoU3QMqd
AywQgDPfq/7t2EbXRPOdQf5c4ZktmemIBL6x/NhBcyxGmvtYU1bEJiUpj1wLe3RC5YIj7Q0QhiX8
0laxHB27cUyP1UxiRa2rO2KcUdRbc4ctEDFe/rYKIs6rbr0MatuWF7yn8QhP3kzGxMF9mJH3U6Kp
RLzEkLLBGTzE6+YGFPUCD1nEGa0DEecJ34LE433oqyhBjxgm3OwAEsFWAIbd86G4X5Nudf/P+4Cu
BqTF2LYkFRXlPu/L+gfCHqGHgKaAmztFmbcFTfEBnC4serKmsZnZ6sxOdghvhooU/QqGBvqed+ZN
GbU6G2OVbqhVNLp9OLT1Qg38oAMEiRrQura5mGxRyUM0VDkeU7T02bbAROZSGWoVRJFiYK3pe/f8
oZz2QukwhtqIeHsvCfIZ3BrzwnJZAK75eSKa7xJTkDI0OSs6Xleum8kW9pUBuUk5i4KqH8NuK/IS
8aSHHQgwyx75wvhYCbT1UR6bQqSYNa32hJoBk3kuJ17wikVhIq58GFUvqXcurtXijnbUTo1yImPr
Z1F8t3WEQzaPawyhQkG7kjF7RNbqbacnvqkySRLNEKgYF9LU0MDHaMwdX1119XEPLp7NRID3ryoa
dyjzCw9Ufi/z5AiLaNt9MvJf68ONkY+lN8JJmQZNpGS5xx0sqIXXBHQWIQqCseX7CV0IarjAoePt
8FfKq7ASeeriCvvLH/kjmyZys9hZb8obhfe8iAK0gQbWtUYch7VVaDA0896uBxzQsmTG4CvrUmFu
ZmoTtg50VeOTMB0ygHsI0WRvOuFaSDQcJxHRqh1SV3IhsEdnnjqUkuyrSaZSXvkQOWcQZ/TIu4Cv
vvFaIRxktTETtzFtRsPvAznkFNbgIzn+X8HmXvheZm7dgngDJcK0oR1Yg5BfQBeQg6zy9mg4r3DH
Znp130S7MHXjDpOANapDdPJvXao8rUOgAi8mY43Fg8+jtGpjuhTwcXsU5B1+7xS9CI/JPnTC0PAV
WELqBip8Sh+zEjnQz7PBFbewxylsW6Df0CnjpqMHXrfAujZQPghzfurQQbzOHbc0dDpQstxiLFD1
RHu9wRi2Li8xvjyS/xyX9bg9OJNd2spGHZX69OI0VEcMPBpe/nVtDIQtMcHioc4xCjNwV1o2Ph8C
3XxgYHFqUoMMFlb36+jybDC2p8lF6+hziDQGnG6lC3SwuP7N73Ogg+fGsqTPXSPoR1w4DcalDIwB
PqAHYbYH/IkDBuuLMHcngSBscszGvzvb6iZyKmBY84lOKnc0yRke1bantMumkyVluBdTQ8ETnUoe
6PNFHeN6GFrVAt3+rxtNKunr43Z9psiKa3PHbz5qZgemN2HjWkNQ6EVTW5UCpQCBpuGwo1hnO+rK
qQm/DgcRSX/Wr13PhVGXlW25k7U+twWHROHExZqnKOIGmmdFgCyyJbLZoB/R+/Xh4Cm7HJZvoxqS
MJU8mquxv0GtnDp0xMrUKn3xSBjBM3dY/Frb2sBl/IEpCtiEAFIEFYOL5NUFtW13yZWtgBVcnlfm
IJuR/ypmsS2wcDhKMZqvhwjKeZVpXMUjUeEXx2rnSN6KDebF137TGdWCgMYnFZH9dtVvj+SLK5Pb
wvSUdIupsX9Q9P12qGnYA5zpHMTlFbBD95jIox/I5QeslYE9KfagcZNcezCFR3Ie1FvudNxHuGuB
kX1I28wgRqtwKRqJKYtuMK4Gu89hvyGolsnXqfj6oAz3ldM2YZDu9py4TyIb7I+2oLuKHjT9ehpt
N4fHPEuWh7EOVRSsIgV0bVNn7ix8eVNCtcUwVNEK6171eOARkkkeLAZunXyitHRVslxMNBfUIG/c
SUG6MeEfLAjHy4FnyPkUwc7++JuPqcZH8lmk/OCy7ljoOHJelLKVvXJTFG4KyhtV+uvfv/FICPu3
WUKhDPIv9Z3/9L86LdXk5KWF9/Jn6sczWMZAVqisbOntbHSKQKCJQ7n+mfvnJdBQ1MmW4XWgHIvm
KE4vRx6oOW5ykFIiltISP9hS7uNalp/fCGThCBG0gNIyGk7+/y0dCYhZ7bvHEu+z4FfbrQzcj5Fj
n8bt9FhTytoFQFp8l6eD9Py1g6sVsFKyzGx1Fnm5kemPwdAHLMH5vnJKBNbzvi7VxCcZ1E2MYiHV
3h04ZnFkpyjDzqKfDqy6lO3IwtXAJ4qzFV/5WumQ6UXb1p/uLMCOC7MxrvGQOEtpLbyd+pp+FpgU
MbAxF6g8+hvtRyqFFwRQy8ripMhwFBdjLx7VNVH3m2VxRBQ50PSiCNgy5TK5AsdgrPOmqCvN3xSA
xWxs/4UnW0eMc4iFFHN7O6JbiOGJ9n5YcIA2SQ+M/ynKKzZD2X9Skna4uFgkzckVE11dGmQnks4d
GDlc/IJqOyYZ8dh+1PzuU7Zqj12Im8goYhFSeUpka2VdwVAqe6QiEhxryyP3U/ZL1QzF5r8b1Rvm
WjxqaMoGCX5LMmBUfy2lJNxc9i50sA6mUTPMzJ34WURPofe3JMT1VF+9zBwZ/BVPhSBLjgpNuNBj
JEPZXXhj6eN0ROhszfYvaQy7jbp+y9klhSkzPbXEry5NwSVhw6FKb6F4Sp4YZTrXiijD6OD+QFKf
FxpjfVNtCBFu6AQCYpMJsDfUpwOVoeOm+nT6wvEav1qYswBeKQZ+ihwvnxuIGk5SWmTSiZRMMiF9
Lg2v6uCxhgLUIlxRUsWK+tyDWb+J0kz29Tmi8wODpugR+4ghwUA87ypt0xwQ8XV1N1U+XD3alHrW
xjfe6JolNsXhLBTUFuXWBui75XtpC467xqYwZNtgye8ZzqHyb/U/FENjvVugbDvkobmyARyIpR0i
2rKNd8bUq+Q3jTENCg8QHyLeyyXKvI7d9XtgghDVYLodCFsqXCV4s849y0WB2OZ6AEfFjzaSosYo
RSSTgrZ/X8q4JrJQK1VRw7RNkZL/61Nh2GQgFSIg+tcR1ab8fsP5DOjI+AEzENomCwyGm7Byf6mJ
VjQppeM1k0CDwnzT+84dQZtd8YOHvxEDUMoohpenQ2fE+jCUxAG+zawLB5Tkjp920BhUEqL0tk9f
+g1s8qzJT4PCgVkhPZEWOANZYKAKJVQM5Dk6MlP/8qVnGz370e1qP+AZqQ1uJIG13O4ibDKztesX
MPZtUE9qNX4re58r1xcZpr9sesvjCgjJ+G298mBjZ6B1+sIzsm6QmiZhCIPqYleIP3CtMKFzx4Rp
XJ26QInFQ9MJO64gpk98BLImhEwL1I9Yv4j3UnNuFJgvUDhaK1Hpbp89AiOF1yewX6hAc9kMIgoT
rCJeT51o9xDHo75eNh0bH7mwN1sCMHhBajg8YprfpGeeKq226I0Je1sOsmLBQ6O1rbH/Lb70z7am
IecIqej+NP5T+Oj5smc+lNzd7fSH9v4NrxhGvU/JHZEUNxDw9JzdZ3N3Hj5GpF4TY9Hu4q7ULqYR
XzUADB+mx6MpkJUF6BInPZ1dOyf5UjQ/u1UmObErSPixPKxL8p6+dRG/t57hXpN6mbkSDv/TUWTO
NaAhW0X/9vcytw+efsJZXq+s0Qcsm3gEavBhHcjDiNIfqWogKMKUtvDlUfNXJIn3eM5/Hcl5W7Au
d860AqdvcUMND1XhdvID+uPrEMvTroWp50Y+DVNLozXFRPzOKPSjl5xVeyOwW/4JYrEnPw213O6H
mYll2kAWM/WICioD3RFnH90ed9ov1VvxJdV0bOFRZq4dEmFbSY6UkEKIC8M4mqKkvLKfAtAW/Hmw
+EZNWshOM3tgS7YUQ3ZFfzQgrUkoBj2FyYg8gtukKRcLWHF6Aki9FLYBRZLIX9O9x1L8UsBqiHkW
nsruCm70JmdxMdqHQ/e6YQqLRq3oVFPy4wgqsOCaej0dvXA+kO6vD8r/GLp6H3XbEWvuienVDxxj
dSpOnVjqB+su7jkb3YiScf1VY4G8SYHxb6plnuIFaD2pFkv4nN2oIU6DimjsCFZJ3Bs2hS+H2ZRt
lRR/MEE4wH4F2nj8Xe2hyqFJ/zOMm2PE5ZN3xoPDhD3uo+DODOsoRfasZUAXy2fKR1gwbrWuJoaR
7AkGp7T662r4zRWoI44u8NSW0xffYlDBTWbIMx5u7xaY1g6sDPjX7JQjY+qiD47Z4Dq6YFd9JK5F
pnia1aoE9R53j6MTGvihA9bdKXWRW4GvbbmnpxGwr7R+j+Vos3fAqxIuqLfJMcxj6LEmUAAZhRcr
Cfu2khQJkd36eR92/DooEKhwRov8OWCpE5WVqVSc9ORX38n4LcdHMFMxsP8FpeyYRJtATPE8ro6h
iTVJlD95cbEoDWTtNfP8BhsiR6XoVQG6QHbH6ua3MdW3KczuZ7iYPVmey+yNT8kO572hrPmY4zYy
foKqbi2JkaOlQIqTRYS3earwpFCn4qPiMXHLqPISI7eQfZSAXC8zj+HabSqQ8ZHC5j9d3FWpo1TN
gTI+2LnIeHK7WO3rN1XfeAKGF/Agq/Z92bIuEFmcKvBCcRJaciLtkc7L7unDBmFeh5TukbW/eHWu
y4qjouEseX+LnNbRZ8B2875wq9UHSoSHyV6xo2As2UNcKWWezn8Ie139YwUrT+qLRwbXUI/C5H5d
ewLBVS9tV0VI7WvImfBA8LN68JpXrNbv0/qLeOLkcx+wd5qzYukYRm5//S3hGZ5tEjkGC1aFKtu3
O9YvbDsp3On2azuDSOPjj728X5g0kHDdm6TVvArwFJy9r+2RMjgOot4dgVHApzCoAKQDNvzTzzga
7Qc/rRS7bZiEcF1sXYn7IzdNWlcC4hLjEW/A1bhXfqeGGlRIU3KdKJj8Pu7Bytz7R93bC9RmqLDZ
DNotbL2Gfyg6u4TEO3IYiX4ArweHju0oXcVr+ZgfY7JdZM0/PUfYlqwwGE/ZJdc2ahjB6P7MC8zn
OPOBfdlFcJIXvH234TacBhKPP8hGbDY0y9Xr7ffAe/4y5owAfbH08mH5GxfuV/X0IgcwiPV1jAfm
MvhEiR579lQJgUQzTcRNM0EKySu6IupADl1u2G9njjxNObbLYMZPHuOB9TsipN1zz8GzYow7tcl9
XbLMHcL6Spqy/C6Qtcaev2JQXx00p34pbsxlo2a8h17NfLPzAwcNy32NOi/RLpdAWNGRTdql5MIM
0fEOCTNUPrBFcBExFYXdvMBPoKcHpL6CP5DE06zcZK8Q21RJNNeDCihDtwNJ09Nr/jQO+AUtTFMz
UuwaqF0H5UeHVpNUuOqbnfEWEQ13pYAseXr+nTXgYOmfy54/qED0AfD/zwV7IQdlDBmK27EWe8jC
EpfsIeF3kdSvQ2N0z4cw2iRsmnNP9o1JWkKBVdk2O4dfICPe/IvC0e2jXluuG80c8lUXRzxVHuqi
X7X6w6+9FwvF6dfW+A1z6q6p5KpGE1eb+Mdzu4iMGb/0QNaodyC3uElhsvkjkj2e5Q0COKIlb/Vv
nyvCJKB1z3/X/4KCM+aSPF5WFdsQPRnMucyReWloVWj8zNfo/ZWCT2b46UZ5GthxgFSQNW4/Yzs+
RW5bMe6ZzuRfdtl/n6G1Hyp7zCy1IWc1d1Gk0Mf9XVj6ePK4sZFtiuQ7dqXvgsb/01ffmAfmitqa
F/7taExCGnwdGOs9BYurrw1urLo6sFsn4ruGIJItDQYjGr548rWXdH6qYHoNJUc9bMBUntwqMdhf
j45aJ2TlNaIPVmwLQ60AINUZZtGfzyOSicD5ckQxX45F6dlNi1sOXUlocF7nNEO5w75FXkcOp65v
sajaq9Vscea9PnSfn9zm4/4sqBI8SLcy17onDxREdkMPs/OnZfbmBzA5TfEC8raZ6YjHWZ4Qcbgh
ZF+AqEty8xjMixtHgfH3okohyVpKPR31TnQvv1CrirxPal8oSBQYAXbbzzkOTfhTqStU/7j4wOuY
DyVwusDrtfepvaMxNevH4SaYfR3CcPIzrf8ZiFMRJkTuHT+IrZ/BLoq63z2KVDAKBPC/5ZAMlh7X
AVqYDYGpjtFPc2sA0mup3lhgRL+AJRvXGkLnYkv3F/b+4c+4/Bjk+XwhRKH2PLfY+DFy/E9GrpDP
7Aecgph+Q4f7vxNvZd0Ymw+00vE9/atfq2rpC/BoaZ6/ty5CS9g43zOrPXnrEOpxTOM6WCEe5MDA
4U6opuTPDebTMlOQ5E9xNX7T+PsXxiBcGUN6Gc77Cqj3XsfEv4KT1viRJytnlK1yKKbtXc5jzt1M
8nQkyXhGw/Tfv/xpAeeRvVihINn0eEtdVjJ0stNwL3pEQbA5La7FpWmrlUNU4HsAKYIPATVIduNP
Khh8Z0KPSq+skYO3e25wZAP6RJQ/0mEYyCpYztRs3eS6Hh3SPDgmkC5zJtDd7TJqpfmVHvG4809O
8n4Is4guaIQZTnJN2ms/ynfe6z2mYsH7JvBuRJlyGOBzoL2AmM/cMzbRvX5qoAhE1xg0wtvc3Xoz
emI7O8y1XwjZ8XPNFRmkCFRXNbc0gFbFI2QjwdgTtN/uXjQ7UFUXXKcpOjRAAc/CRfBO82Bl/sm7
aitBJVFL/8YX+zLoIaagXS5Sf9C8LbY8cBAw/q4lnqRi5avQP5fCEApqinHV9+17ssaar/83UY9g
ws/DCcDR/iclh+Fqc4y7ATk3iVBXbwfnvgJUlNGKdBI3ZxkK3Ta7a7ZCqaJrOR+Z7LOQqtF4QeVv
V2kS6xrCuSxDjwuCoSJ8WEXFxkottxOPQlC/e6MjS2LsvSS46orbxRC/ZeqWWoaKstkJfzO6UdcH
RXCr4WlVKGap3n3HzHLwDdje7t83GtyYdekE4zTk5mrasS9bkuLkwXvHuChL46lvhlwIZgg6wYCu
v48MW0JqCt6g76YhKgR0lvUztE/NNl5rzX3f8FL7v1ZJzJ9uHyRbmfr9wClkm/xUhYMEsb5Kifdn
Q2tvRmRT9utsjQwVhuqcUYPA2/7YUJZ/pfefGwD9jFbxrTCeMAt4vdynfcjWDvcy4Z0oSvUER6Yg
Vml4Qi39GWsD3q8VCAXMrl2+Y1KIaRZQaX8tRy6DCqlJYvQ6sKfEIGaaL8x9IYZtvpEs7Pt/9EgW
aSFWxzjSYTWf6zEYQRqreP1DLoURFtgQr0b6V8wOr2itS0EhY4ywE30UlSqzPxn19pw4Sqmbosg+
B3vmAz8LSn5afwyTuErO4Pbp3byHgW7Afkd/7AUxZY0GGxq+/sBP8GjagHEXcJVvtoFHATrUfsqH
HaMqXTIpzUiajNSqz+tZQIr3mdTABmmfXqJ1j1IrVlxuiOso5g5uWmOfkrKN+UhcsY8VdD5lBm9z
BYjvE4OsJuw+o8zDzh4AZ4Y0txTbq7FBb6o+dmneCP/y6d8VSzCmzly7HRh6l1mY1/bs9UIKKraA
gOiEydIaivT13TVTO6r/sTQ1+QxZQRvSePEKZXyy2bzwBZ09cX2ucfq38bMpqnEWCEC19jcomS1I
bKbv0Op0VMIApr8PCf8/0IR4sf6yfdZty1AxACFGKK75d849O4KHRXrCmfabmonb/0Q8D2FHkzNW
zpnQF+I3l28PCaTdjzBeCf/3BfVP2djofn8idVwbvR0SylR/adBT+kwtn8inpyYK9+bRC1Fjsd9d
kUXxc1C3Z9c/Z6n+r7SUzg7S0FFz9C6IewBmS7s54/ZXZLu06glRtIG+IX2HzaEu6lF4LlHzre7I
plredMSlfedf4sWLQ5FbGJ/hC9EUAasPMmNE6JqwBIuuTOi4kBFTLIGbP5yzNRpRWumS+LzRLpvQ
oAmBQ3i6emrcUG6I/Pjq0ao7ySA6JGrQqDkzFO8DwnDI5dI3dhSk759KGzkwqCsBTUQHNMCSx7UL
+gQ2Wok4DAGdVDOqOfJ3jWHRoys2+Q2APdTCXpGWj8jfMBw9kbwKkotsjJEeRQKIpxqVebE+X/6K
nlBeUxjm4JsgKRLdH53mBmPsCEVQAdxry5v0xNblw87kraeek8+aeLR6N3n2xfCdUrErg0MlpLGt
D0rpa9mgbk0lAFleaNXEEi7mlfmy7ccSXP8ige91rGZaX1b8PXyLVt+EduV+RDtwmXUmhlp+oJ/n
RRzG8GcivY9wha4Le05+zsAomAlnf39KtdF+wMkl4ALR2S92YhQ10IdTqPU7wrfDLnc3xErOdjr2
vvR7s9zWLhfwTda2K2RsJJyEQuuqWevnJuLTvY8Nldcr+R2c7d3jlAmvzErR6G4Ym6w357JiIwfN
bIc/I51zNEAsPjdhzIESNVpbx/yfhHR6MLtdLBHQnR+2p0tw4SxlSx+mBxdkUgdsFGTv1XWn+Xov
2h553L8ATl1gYAwq1L5t8whLJhsdmH+IBOf6zmV9tdjat8UwWEByVjOGtNubo/2WA3ZY2mlc2vyt
GxquujdO5JxmXIuwAUAElim8rVPstyyBDO2slO1scsjCClzvcApubFmFcBHiYgb1ajx97Ihibpnj
eQLzVlwfmmgcMpZxfD61NoZEsRPUTdwsibLfR7yoaRhpo1CaP8Wt2O6rEDwGQVL2CFlifL4RpqW9
f4Wtb9NpxX5PWL1C3S2CrUKjygSjxLcBPAxdsZrLAtMFLQWne44n48Y1PUbnjNVWtQ1QfII3uyd+
oMiFYZmoquL0mWb5tqbHM988QlynRiCxX8fvM/3sMld+869Vem67Nbm8pGFMfUK5FgKuEGKmsJco
1yVvmXKkeJqYTsILTBnVcZvHJdL72bN3mwBzKPVkiUCoQV7ytie4MQKt1LdyUCIycHwfRKK+7k5f
AeHuoX41DbAxp4aobk9T3aik4k07NBaCdDfl3wl21XdXdsQiBPnPNiVKKQEzYmfULslVsfBocWhG
TWkCUOC8SVaHhEEk+A8t9Tz6DG4L1W0IR57BqV9cuh8UMBfwslQ1yJBFQnA8jiLJLnXNWjb9uE+Y
US52FA1kvoKWrVNAokbzZoOq1K40cryEtOrbb27TRZSBrvca+V2VrIIgdHYNP23wyPlw7HllgzDa
aFxAg0w9baafKFWA7aSXzXEdLVdB+UPvCXCBTXW7NXzrOIC8HKU2C4BMAc3PfJm7Hfe7DXM7nXpb
U84H0f77xyxoGaQ7/S7UrqZ1EUPl/DNQLKtxlO3q8R8BJTs0JRW8EzJW8zLSgHg7TgleomWBq5fC
L03GmPUXO3gIWiYqmftUF4c9/Ja/YUP1greZx6Kag4eO1R1xjbNyKsRhRss/PXEv6FbZm6cwRudb
eEHQasc5u+SkkYPi5VYAqH1pBDgQg4UqsmvqZ2TcwWmn5vWmRMhHML8updfzcYRQl26EzUj9qJIo
3h2yrvecEMCOFt3TAbaXh44E/AwezMhvz9LYeLBhzEbVXp4zFFLdkpI8mTglEJ4lTKE9bisvya7K
h38iTCqJsYAIcr5CXnIdWxTpnGbCAm74o8d4ZZA/OJIjKSHHCZQrKXBAxZxj9xXYsD/QkKJhB+Jb
jf3lYPxaFIlGJfhAgx1hvqLamr4wRVd3vlZUN4PpNe3NU5DAfMh5hUElgWqvgCgxonjTZxfRw0H2
M1mdasu0PXkhG0CUwJnmAvIcK66VJWGZtn7yfNEHn6lJndmj6kU5qMMvB27sSVbNJsBAYsPlM7PQ
dVgvPVdjr8AinKMew+RgE8bgXWPH5PX2er8EaOwr5gBZgKYyparbOC3P20/JkPsuqwZol28WKlrY
5EnpKRcwMF9RlzCKxyspESuDNwlbfpXE6Vk6jGGLsYlCIkTW5R2D0SvhzdQLQ+CYKcftFh7TzfUV
sqwvejK+h6KnA9c+9hfzGSHrV8wlHEWZL9RflM3a3cZhn4uJlHIzDa2wpWPY3eHSusGekgkq039F
dzOCgi3WfQeXUWJnqx6KcQQ7VcPafFgKSCudSWeuOMNy3nVmVILQGayp8LfeKnNDbLgCjIlSmHE2
BjOl3kaz3zIKTkDsqAfoaPAEg8B5BSqgOPiSkx0nqqiZZsJH4BI5Hj5AJTRp0/XMU6wUHEkvzLTB
AjNvdc6x2Cx1HwgR+y0NOvQry8KdSJjBKnskcHPV3NY9JX1xZvW9kATZtnqEzMgiHeS+rNTRmy6a
AdANaJkNc2ExdsOfvZ/JcYKVaRgCxmTGK//3QbEOBsRWHskwd+zhg/ybUD/j/UUawq8p0bVRDTDf
eoz3Br9PLoz7XZ3VMYPLUDxDuGnxDOJ+IdFn1mPQzAFG3hGOHd2buVCmemA1aQpmvgtutIIBZ3Ct
+49ltnxLjdX7QyEWJwoJrNobjmSGjsJ33gnTjC1mS2/IDrtY7YvKz0aiLfLX4x6kcjXk3FPg7Tp+
a7B6qWlit+V0E5p81iUiSefD+b0j4M6F6Cp1UcmXqFvHlAahRCq5qyD+E2lCi+MdO/gy2lmeNeLM
Gou1DmLdd7RBBLP5ewljycB0ElIJaIZuGQgBfpEVK8s+fZAe1n+855iwRTcDjl4eBfDgR2u44eEB
M4UPcCeGQ0XkYqqjK3SpqDvucmHb3lo3xh4TUsKrKXPKQwQROfOJX2dF+iKrA8ri3vPdFm1sttoO
1TkbaA2p0ay9s3N3UANOyhPEzrNpZe1dgakuKs3M1QsIkKGQj/bQ8ecQjxurGlxoXckv8I1lCKdE
b0CwYu+UpJgiJQyI6Chg/n5Rb370gUk9UktjlqCMlUoigUyQw3vjoQ67jTnliZcJjDdVc6RPAnaG
hbeh0avXn7YCeRlYQJRdCLhQBMv2eusficHJtStAdmIWvrSzKYcjmdvdRHFgwGuAfqz9l08j72zO
RJ02QcZ2sXLT+2RKc3nrPNd0BMtrCrVkqAwrzYR0puDcwj8gGt2RaqH9mJCa4+uo4iCx0L7rxAan
/DxQ2tnxBZHGt3J5jDQ2B49V8Q0pX0dIn2qIM5lWFchkJhQBwExo08Dl429CPDOLaqWf9Xf+adT+
12yTWisWTvKIbjroX6/u4eQQk/RMbyPfc6PBG7+V6QHX88CAWnfHgqq30HBhHKxcGbWBEBNUugg/
LDHYSOkS1i1pCfx3Lrabq2FNJ/ehVb/XTHf4ovGH9x7phAR6LmqCKT2ns+/DLlf68+ryRCz+E9yt
iA5cMznvq7QPgT+HzEqIoR4IYUBiACWmkzAVb1N5/hdXSROfAHLjAPGWKMPiVyfrqdMURnjp1RQQ
D7yYb9WRv4dMrBRFoxsAlyovxMp7LaLI8fnNovRHZEzp+6Pxfy6c+duxLgjxLxv5VjnE076IYcOy
kHzweYfmoPrfZkMZAQ6b/ZBtS3X27qy9uoPwlyuNMDd6lVW4tcUXQPOdmPMvAMLoYpsQAp0IQfYD
ZWmr9M0vqYH1Vm3Z2WE7HLfQK+qT8P1eJ4GgmykqCMgMPn1kfgZZtUHhkHk4Fre+AS7D9+KQiUnY
miU/yAn3C4acYJ92bQAgyA0OP4I4U+vkacvfT9IERkt2fOGfZs4Xw1Mb+ix9h3AU18+iSxN+JIP2
6+0MjLiL5xDUceueqIaFl11kmxNzyMuoisNgBhZUPJOkQcVQodog1GJ+WKbLaCC8xJxqI+m+G1n5
azZ9UMTBdn814qDzAnMpu8aSJ1j57dPZx5qsaBLVVad3zEgUwp0Ak91XwDA7EaZ6pFjpqdWDGzHC
YYsyrhpuOexbytmyduKWQLMCrhG6NOK5VFp1AWRBuActhj+s7GRR3tXQoXFsmubBD8hdzQOr88Mb
DjkWWYYX8BS6AJ2f21kJMqxgG6MEb8/7YI06gDA7oq/ZEy+v4P52cw8Qqg03LHN1WolRR646xOAt
IHLWfCrPNv9UsAGFcEKpTWlO/O6lVil6BGo0+rIRR96WjQeuD4PbIbH5RINKqYPwEKtMiWv9pMUe
M8zPZjYOzzkH4FI/s37LdsHL3U6sJUGIQCsB6RfVZ1PtKv7iREyl5Gw/WDIcXGUEmrWqii7zGPjG
ZeGswnay+54QgqfSAHEQ9ep0zuzZjO+i+Fg3Sei/zOVzd9P2RZGLAfzRpjbkZBGNevJOI0F0W0Pb
WgwVZiFUlZimi3NjFV4H8ptoYM6WNJCLo71klVg7Xg0yNlNf8cqfPO2r7bcNdb0zFe/jPkUD6OkI
26MdvBE5dPlY66cFrsS+YCgmo8fpykaXMIsnJqx0xOCnT1RR9uYtAEUrY0QaE+c1jfaOQhosZ1iM
RJ8Nj3NHFxRk3fRjPLzSWl4/WHm7UNnnSQcmcuMwA91vlQ5paZUeSakiowcCFvxgE4BSg40pJSZj
4SCSEpIYcGT1bWNZa41vJ8e1/OXFdVv++ERNRls2ciESkIQCW4vZ+xvBojRLGIxxhtBUOr8QF6Bu
JjWqpmx3EEW7MksxJRF6V0Zz0mZiodEDMHh3qiYAPEu+epEhumSYyH/+Yb+y5jQtBKMCtGfnQGPa
b/Q4rWpWAOxptgkqnvODUAv428qi3cITQsEkZcSFpIXfn6u5PiNQv++eERnrGUBuv375dcRa9EAv
mVP3jTcCCICWbNH2drXoc/Y1RgwlmoCTEOXvAkll/EmaOQUq8GWgGm245KiCcHW/SXPYSBwtoX5l
hpCg+snrHDu1lNsbmLG2uDo6t+dD+s76HEjlxmN0molPN7e3wdFbhbRYsqQi0kkYIWLqB41syzgt
0yDQb/SaHkELVo+4oRm4W74HCuVulWaWVEs6JfJHjKdQe9YkosKBrx5gdnvd4oZ2hg81rzohV3NW
dUHtUCUyLKcagxcJvta79h8Q6ZLhe6x5IGsO/ShdINnf/Q9Lq4qkPaJ8oA3QkKIL5uLEf0sdMXb7
Lnjl3ZABIPNK8Usach3miBlkzzf2oiT/muR72PWAySII10ynv3NsVLl4bN2CtPsivx/3jU8nbCYY
zOdl267kYI/lgm1g2VeuP0HzHQCjroLKVBAkF9S8oaXZc2v/LpRLlVNsBltjcJ9Xz5VxiWEM4aFW
zF/nha1tMFJpRQXmepK5yDnNy7cVtB71H7pXJZTCuecSqRuT3cJkDr1qtcz6vo9EiE8cKuw4MExJ
Bk4Ia9heXTYbzDPb+RBNqTxYkGYsOHHan4NzCQp5oavZJWzikPJP/HH97gaXxR5UmFHXRNY4toT/
S3l4pVJJJK2GvKh9gXYjnF/odIaeif/sjeVwjybiUPvJXsnH+yjNYUMQRuysWeS6nIDFlGgTpoex
3qzUiPF85mLqtybjELTMPU4ukk+19N+G8fMJRoYXqq9KwlmmC6q8+gBZUGIqIy/i11P8eVwWp44z
DeiQmEmrGxLuaJuuwPSrJ8CCeZChipTSG0/IQm9hEQs4BMbgod6LAf0+W8s9snwYqpWz+4EpJc07
3sWxdFmFlZE8L56qP5RQcAu5JEhCMYKiVx8IbFqHu8vZXk/3nqKc77FxwFGsg75qnHg59HBJeBQL
AS5jfYc5CoEOLZTuUyDpg47vYHLRuIlmTU2JY3gU9W4RYFvwfBhmZccoLEKSaflPMTehwxmrh8qq
fJ8Z4MsrKR7AnG/5zQLRUaWGr1ErsSAWlnTK34stTB+STKZWCUQyf9EWGZJ698IBWyoEtnfJbhMa
IKhBpv1UDvn/JPSxlG9dOSsw/GrjwcX4i5VPLJFbel9zOkEyEkHibs4L3NlUv2Yk+MT4CQg8HITB
KeGe+a3dvVqbg3MMY7i52IWB1DT1RVNF4K6HUN0D/aghe9B8pEIeM6+IHzqI+AtJ0qsvoaxKZ+mz
RFz9ECbju/zpmMGe3wJ+lf9EFxIPBPM1UXxfu2aMUi1gJHNNK/EzFTnrE/hOlc62ayldENus7Tn5
2n7iGqaRlzksXuOtkj0cK6ZVVL52Od3g+og/eOvXzBjGWY22xEwesJS1d2c1xRYnHZhZQbSl55F1
mq+gdvf2b/8LqSSMkyl6SAFjXngvNopIVGM33kTbQyT6XDCKsBPWlIAlXywn9VdjKJP8r2jDhcnL
XAiRB0IZD3IN0VYTQyX6uPByibRjL8juO/sXTJ7o4drv8JIkxVkt05kVWMAkBOsOnT+huvpyx6ao
0VTNyvVSSpRF189xVTuD2Pu66VZnlV4EozAWRS4Haen9s99Oe7lW9l7vKdKJH7I5ZElCrsqgyHUq
lcgVXdnc27ntBU9FdO0Xl8jMZFNOLXGYfy0zpteNGwnkpcXjOsyZwAQtxV0fsgNFGoHFx0VH9Ll+
1t5MI/YWcT9e3pL6h+nQlw/DsNZbSYCHPCEY6+ayDpoZGN1Uz78FzdY2uLGAlxfzGYLJ5pUxuc8o
TSF5HkWIEvD2WK6/qzqbGSAqJ8zd/QGtBFCKFQNfnTmy/c27PqTs4leos6IAq02Y8cTPwQxXSPfn
HFUSlFmPbl1tBgkYVWWFa3DWjPIYhVQDQiPL78KLnH7NQfaHbzsR74fKKJs9k363uNWZJItP9LYV
fPyyJW2Sz589uo0FOk1TTgn3/9ktsnjURpdm1tovDxF7hp4UhD2ruFhNkL7vjfXTbs02QeQj3BcA
LQUZoWoj9LjSXwLvuCZhMCI5BKPGQO3Q1awRh+c4BJZxcrR4X0q3dVRtdUi0WZXqF9IM+50hXKCB
+4qreZ833UVfTa0k8g210ORZMpXMt41nR7Fbq9fsc/A9agCUhsK4SeVXdLsza2NEqXoQDySw7tyN
2NYD+ueNP/jDU9BCBFIyepM652Hu4dUDIAE5Vc14n3VOLrafCmxmm4tm4XYdqRrWA4eRFnBOmCh7
R01ag3HqQMmJj4nurvDauzr4yYgMEODOlwsLH4PthGW0xiUph8v4Ff/vhmcJbkKQhPee//LJpEEq
xUBSupO+mplS6GsNWDAu7xU33GcbcxbMWe/6Z5KvWn0tWf4z4QcNLHDdI8l3yyQMwiJOgmCZHNc0
GH47vx/25WN+GP6MTTuv0BtAoOwRSOglZ+kQmJ4NP/9DTavr1U0095UEpe0IUqvCxi4wqmrrYkAA
5GGGKpsluir7XBRYky+7ZGjHMLEHz4N1yTWJ7vqK24KSZV5Y8YJGv5g04eMQVCI0MCmewm7IGkmD
KMZW+rM1WFNjsqePd+yPm7697o6M2E7vRsGkAT/alxGgqRFVzEzgFcHI4o98wztCeguVCtWAQuZ1
46+/VvmSIHNwx92S8hfFr1nOx6k/TF8BgJwL8cL1B8gN6UJXXyb9lpMEqB724TxJKQfTpViOcBBD
x0lPAoLaYqlAqk6SfeFFUQZHrObvYWMKCNSzNcyKFdervzKqp+Cy5ftj7o4jyecJUv4w0pt1Lktg
MkG7N+k0JOyLpo8VurKPAWg54nzLdspOyzU8sU9It1jr+IzGImRGqEBW5N4CwkmaKtZ1Qgwdfj4G
WffKyCzE0a3A0RxrW3SOcTNFtFUTTz0eKCp97rcenpqXvavyXDGrUBu66DgsQJuuJJJSpvS5Qnhn
mrG9Y+ZnkV0+imx/p3jqmdciAy/Af3PHXGGAknY1Zrz2IJ2GwLPhP1zU7sJYa2pVAlDhvFX3Utr6
MEr4AepUa0I5ZqA44l4bRu9RRNstZaEbZYbjeQpqArMBHVh9FiDRL+e5jTD+fM+N+slAdroRjPQB
OeHsiHMpB+F2ywLRPJGP+15RTn8j39ERjMFMx0U12mdHd95n896WfHlFCXwPXRTloaWPJrxd7CXh
4ZNnfWk+rXc9nWBO8vbkEaqz9RrSqCd+VBHKb6XXf+ljP2u5TVq6O2Ff1fhZuk0tXmnizyKfnA/A
+Aq/q0zLgxpzsX5XVZE5Rpg7vNF0ZBORFvIuXnTdKo6muPY20YdcQvLakKxeE+m8QBiuQq/3I6qt
OQWWQlwIIKIqN+FDYOjZIkFsUGzZQciBow6S9hK0lHFlKuWPNpQ3t1FAgyaebxst8DUtMxGXhapI
Sue5PyTfoKSSphMl8IEl2ZzTKrZcnV+kzDYLziSbknIjrspT4PMJvkCp3Dq35ligA1zRX57LXPEj
yPObfTzZK9SUGwL+ApPT3Cyi6d/X8QshxsN67BbyvVTgJ6X/Q4+1Tz/m3HB9kwrMPOK2p/ESWZxy
WK1Qukz0VwNcvO5LUO9mKJ5RIOhxMEEsXs5w7nBCQctylI+OQt8kvXcaUYFZbg3+MDL6ETxqi9Jy
rjslFhrwX1bl0uV5pQLwgTFsAfgIHVnbO7C1Opv3Ef+Pv1RAapwZohyQDZZ97GPTli/xjZ35CLIP
zOc+UK5loQ91AykeeLulkOXcxyh4ywee9POkSP25EJhZrI/zp3hggz141PtvfuhN1mUEG5OHgrwN
8WMbPN2+NcLPTiloa1fDZrzxrrNSmUM/AETqDNQq1XHLX8D39qUglNx7mgR3aad9G3Ade85f3B8s
Jib5eZ1mzSEDIZdndc9LXWhfg5l+WyT1eQBz6ApCzHa2h7cOLID3ZWyW7BQfRivI+N3JJ0sHRwHy
nJWMS3FBALUmfSy9lEF3NYLfzXsfHGTPHF0gp9TX+reuP6dHhehIHO3YyCtvxUD0urdMDS75yPXF
kAtcj8pYB1EbYZGunwLlsGWkXVHI9s13PeBsviMZ7ITN9jft0cTkBJdGUHwoC1iSYPkHjdbTgmGj
t/0/kLNfL3m/WYorHxgcE5OC+YMFUEanjcUtMpaQ+I4ySf+gwbHNUYQpDIAg1HM73/w2tJz2ugag
+c2cZppAUXvv+9OuLe3Eymbx9srnIhBzEI/B/YMUlXLk+Nn3RApPQESv7AhNQECHOgfdOF75Dp72
V+4gRsyVMR2A6sK4yNSleXYbJvtw084a7vzDXQfb5TT+PMjhGimB37VHzxW31Xrc6yRQFCKVdmWG
VakVE3iliNA+74/0hzIxocpse7PBzirz3kM+cvyP5+zcA/RaN0EaiIPdvRlfXqN+yO8Q/mVXBVKt
bzBTEFN8TV2+FQSKJ0KTbouY8wMbQzWFdMpabJyJb1TGFARL1X1khDdVr2N4hxaJzU99u1wJABZB
BZ6ig8Eqfb++M5X2RjokEULhUv1u8Aet98pGjEhLzeCbtn4hDetY4eZbrFESl18YswUIS3I4SfLr
9XVRmJxP9JQEwyJACjK61Y8PWzlgtAyeWadLMTvwCEPnKvcEa3qwUUiT2G5M61v/d00vOuclAwvw
vM8eZTXGWIHxB0q1xB2UiAgmnZEqdlQkFfhq0NWv6rUCtJPDskQcyeaNYpDtUh51PjRrWH7DIl3d
2+BPkeG6kkedXxQ2p5mnpCNxMk6xxBuQ992LaP9wDuNDpgk7Hy+l0cPIT9JyMsCSjM4/DROaO2YY
gF+5v5j0lrz1/NDRU96/1OPfv4x6UxwmtOzYhqtwBlYSnXTZSMi2OGpUxvYAM2hHqocDBQXt7/Z5
c7VAL4GLo0HbL7GbPw0WbycOaXxP6dl9RUhGpyrjUDhB+Mwk8j2F7Nfi+UMdfWwj5Ul5fUx4yXuY
2ZZCq07xxo1LtbkQGpSg1/8GxrgzM9MJTCAphQxFSKh3Jik+5SpuA2eFoDVDMlKZBeA+kjCMvgMp
4ekqr92F7vXKDOvDsPnDrJwIkRF1Llc99dP5hqKIl/ka6D4AGPS2qqRK6TNQfMVBEM+f80H3dBz5
qP9Hmm9Hs8IbWVLsCQ0E2I/6qA0ti7ZKtTMELruSaoj1sMC1T5R0nnTwyCu96iY5i3rVOmk+MyNe
JAw90cXFbUjqH16iCN/ePo5Ko18+fAJA4TiCwGu77r04TFKCFArWHeb7h134NYS3A9E4KPKw0xhP
OUaRy72oljKtuf8+O4OYMBcKn3Sg5F3f23p+zw8DQCHZ/Qvxy0/du2WP4OaOnANxTbLwgiG+Gf9l
jHDz86fiA3QKOSj1JsFtDK7CrEUyZztyd0RKbLvI1+OSLFSntKXUVR2Nmf+CRmsYAgryTdc9gzVW
MrQFG1eBGyP1uAU4oFyPsYnN4DfdUKSSoxjW1M8FwWpVwnjJmDh+06gPtFSWIbxKN/yaGSUYNciN
PfIQJ/nck0CThsP6oCAwB0hG2X1uK0rCxo3YPZVEVueMOf1KR/8U3hqEdkbRDSWiIbNdXX5WqEjK
zGnK8oY/tDX2WSSUsQuxZTWEuAnqKil6b2cmsFbLzrMnLRLi0sHy75B1ys0Ki7eaGspWKF0SgQxL
J/hA7XHDGuA11jEKvF3fe2hlyPa//CrWErPio6fkRNWDUwjNF5js/22o7U2HxytozwNb1uN6+rzW
f81XNguBiBFEU7fFYZr6b+Dl0GX6kJuIcKBoiV4sCmFz3JO8Y8UC5MmjWMwT7kE515zYXU2A8nAz
n7mSdNHk+RVE7KE/7mR60HXGrLGAZPFZhVQu1O/Ac9op0IALT6dV9EEQlK2FGXvlVdc1jlMobO2R
WGUjQ0zMokcgGgs5cfTcUJEHpm5qU/y4Nbpc3UaQqChh1iEgyt+jp3oZr2TTH5VDsTFt99icVBIt
zC6/17+bXL1KHx8F8qYNdknVtJkW8DBTz5cwLWZJCoFiNLZhKZkFdPQZEK66asjlaNsyHonHY6j/
12V6jEHKqYwg6mJR9oVg5pWVGI96wHDoZoQIVKLBqAVPA1SqoDU+blbl+k7rw8YUEHpVYWib63I8
SC/zIrKNP6b/R9Qpdkl0DQ6InFiFqUHz/WiUvA3tzGPr80uwDDQ8w0LVD11Y8aaSurCGwXiDTJMA
X4sIeEd6qJLcjaqZAhLQ+xjff1ewPp3wszLObF/Fc1PFn53BTSqoRhiMKwXq1w0Qi+2ZzK1QdzeA
h6D4iZBL6+zKRZkThrAbW3xeLYj/GR2rmHT6PqL44AITVmJWliBD14WzIUAG5hrYWexYXmgtZGS/
jDsa7Vmj3G1a+4zVcKSKCByqZxiPRgBogXACZHIqGTYw4S3Lk0t2mhpn8C+OcLd0JShE8ZPAA/Z3
OqNOTrIui6Lyd0JKskp3sB+btx0e5vInKOKYpnlng9KaCy5brDlpazjitPlc/Kj9QUGLpnINXnQc
9mYab1k4jdfvUV0ZMYDqMxuKE28sGwSNt//GND10IqWYMStbqp6gwOp2+xLbs2l1W4dbD4hyleNK
v22nL0DQnFEQer29lQs/j4bv/JYaK6mK2YPh6tfu37THvU7oGcvOf0YAKIKZL9Qla/fEPJIt0I4U
kaSAO9kwSVFBXJ/mlNi9aZny5wX6S5CfhcR479VEKb04jsifPJ8z4X13mwnD0AioRO8jV2r8u5rF
4GW0qC1+OSsK54wYesNYJg7s5B5gY86dMzrEpP1Zz99Ulpe+HLSH3q37piLNzxuhu+Lz/mtqtzGI
HEvZ3H91dB1n5KCPrswwTZBzuvJ3ZXhpSC1srUDh2dOa6NI2tcfnlg0LELifELFcceSsYtd2Fos4
l94bDEOt7Lp2AFITaVnMYUunqfZRL3BI5l/Xbu025HXadH8nOEZukSWQqWXy2LG5k6Y8PKzjtfnv
3lhVrmDuev98+Q9UG0aR8XEbxh2xhhf5KSAfIS7JWbFZnL+GG2oocpuDIls05ISANgceWV0FvPoF
29MwlQ30Q63j+vxTp53EXCJAzQFzCST89zdebN/CZFmZiIaSCEc1aWqYpsIpgVy05HLh4emk52WW
2YwTBzWakNBl8U8wug/x+mwUZrqOlsA/ZCS22b6TatdAwVqQo6regRe3ZCkvM3y+pp8YriaqFRYR
cXX8z5T7LVY6ULIQlQeEX+tztams4Qb9Y0X4tBAbDUDrc4g/58IO4GFsPu+6PplwvYKqEhMmSoS7
zkSm1D48zHPK5liQK8LQnn/MhOcg9P6CXAzxJnxAS28iw/0NWQXe48kkxsMlODixOs/qT8SBsKDC
8zhGaWVciNhLkNT72qzzY1ydervZTWMwS1IJgK8GHtPvX4vSm20wZeNxBr4Xt8pnse1O/Pqlg7k/
WqYAZN3dSz4s9jw3RqqV3VhFfLxt/T7R7TwugoV8JJnjjiiE6wlIHLEnMQek6F2bd3S2Ekp1MxwA
wk5MZwMcRiHSzX4YPZpio4u2w8ix8pVh0nL2lSrb0pEbiuLTZJ6oR7a5Fyznw5obb9vTRJ8JjffG
MrbLSobJy4aR+xvk1mNYVMr8SnMfStgXv2JAFKnwg27qN7cNEwlBAhTg4WY+PkKxNKFCRdgg50Ta
FNDVXJU6zsSsuJWI9UqCD/rN0imENnBRCoNLVFck5mKUmX91uV0IcNQNX256GrrJuXZpgk3wdI0z
omIOROHQvu3/E/g1H2Fa6m/7z60hQ3owRNC4iwE5F1jUVzfre6U9qcGVch5BvrqTCjcjPj87okBt
swd00PA0sRgjGnlEDaqcK8tHdi7bMn62zl0CHhheruj54jwOn+lPlVLyhaeZcpvSuL3evgGkrwER
Wk9VhMk8vNKTnRY50PSiyE8z3RA6tfFD7CZiH2c8MwGQ9GMv89KgsvNQIqigmLR15HoFTxJUUije
cXs4sAlzCQjzap2kHDcyG6C/b88fsu2vKdnX0+z+fbiH3eWnLfTxdPryeszzQOZnpFKF+nJWWtmW
YK71+O9idDKmEbhN7dihA96mxZn9mYlaXaXxilRvq9X09OVuw/7RYWJNfwm1GPaadnZA1LzVg/zO
mdN5Z9HRdLSYPrGbS0Ihr8GAuUepmSuycQaBNhK6rgMb1UQPpUATA3+vKxwzdMBK6xE7lyFuDVKA
mwdSGse9reOa2IwR1HXXT52ZLf92m1VwkbzDDxsXPmu556d66IaHO8i0kkn5K2loNC7VcQYTRmSC
JqGHk7wdst1HjqXm9g26aDRY6VIul6S6rA2fUIrS0VwzcvmvrbSPI9bbYx51u6yxY4Y7t7YD8x1M
MMnL2HAgfjrsxmOHQyp4rErxzXgzLMsFmeKWLHzYRcpEiHHkaElLBKrahqFvwJX/fpMueDzdMGi7
Ha2Yksw46idyZ5QzZJVWnDT1gxjQKrH9HYo849Sk2z6et54ytWXszD50cycKGsnawyYChETt9izI
PEbp8gL3zB1/Z7Rfj8rVnT2H4LwpHUJD3SyuJ+lCexfjmiGs7HKmTH1S/h/x/Bv/dTlJYxHKkR6U
/0k+8BFCXKwu1hjnQSPv8H3rmUA5K4eoErCr0MFispeY/O251Q3Gr/UPrjj6q03mU/FyISbDRwn6
FQVAhrf6khfyEaITZzA+VVa0be3ZE9tFLgS2WpJYHslC9Fzzli/4jnIvUAGthKdFdjowfb3C6K2/
Si05BM5BMKiMsiu8SErtvsk93fx/UL0DlxDGUPKVnsHn1/t0dhRbDdPaUxne8CIDRodJcCkPDZUV
uPmKtDdtVuvqzarebhevy9eVWaGxmGO7l/8mreepw4pT57NgPMAwQSteTofqLKt226S1HbD7tyWd
NPCmHrGY9jydL4G2MwOP9zSaXN6lZHp2fiwDRbi0pekg67Ka8rduyLw5Ky9SS25o0f3y8w58M29T
iYNk5HfdAMgygSUGQuboQIh3i6dhP7wp2QqaWsmdVEpCCvzLcJKwcTMQvGMUzdUL2UYB1DtKMNYe
+iY1bleIGM7fnEOrFToyTt9yGqsFJoGlnk9c63SMJAEtUcEskHQYbSTKDCwHgGhIUw8vzqSaeuIp
a7I1clTuqda6PEssQzmEnGlBml/5xit8bpkA/qtwXXP7l7+HlzP2gyQZ4XLpoT+MtmauqiAkR8kT
mmGtfy/MwSvDWfLIUmPl2qOFl+9WJZnD+KumrxdgWPOWuJQQqmJbiIxzcf8uksIkEtHnDfrSGMk5
iicQiqd3yyNW2M/FV2YBK+kDeAZ71r1ojEh3l8H4fvBQU2UEiHbAD+b7be/aqjf5rIkPVIYdgnNv
5lgAfNq0Cd5MB8czt0Wk7lymCbrMpj6/RxWl6ruQ+Z8mOiHO8DadDsvWBNwpily1ZNeKFFBEx+oO
Go4Y4NpYwLCkpR8HXLmZkw0GBM9aLGWBMlnd1DuegXxFildQhQOTRsg4S8O5thpfXw77+p9P0xtc
ye794lxXWD9VzR63OxVaxkApx9orySNQCb5M/r1VM8B/OmzB7/mtRqmcRMnD1gsFx3o3BY/vwCLK
lnKEI1hWXBL7WS9O3HRggkKvBFIw6/OVeq3WQZ/V0FegSBsZyX/wgb7GjNJ2vxo/30KEf6oZmIav
QJLoGUB82/VLLAtGy95utJYgA1auJZKLbX56WmwQUaKyJu0Hpo7KOyfEhfAiifPGMCMDYwXEWFh3
Bp1gN2BCSyBD23zpaCKjxzyRqNp0yjLBnal0MCbVNhmQLhZgKvh71MTKxa9zlS6RRZBMBDez9gWJ
UMccSihqC8uTxE5w/5PFzyuhzI/nXGx3ImFMNskebmjuW6uNAKxl4TMjIx9i2haMb8X07Mi0Z+I4
7IDWbUdq8vFSnhE9gYBa9sKsQNRTN2KTzSMIcVvqHh3CVvbVZDdlut05EUcRCncR0HsxToM80D+4
UxDETxkP/EtoIjzT7nH9BqPb7Rzto3bCgWVJmUQbcDMdXnGfJipYXioORSqlYIi/jSaitwfIfQJc
hwG84Gp+O1PdwAtMv4CjBMdU2wZ7OQ07EI2JKbTQMT/oMkilLJ5JU23dATLkC44rMGtXKYNAJGoX
EcM5T1ghKc7nhhqVFlobRC7f7EgXFW/VXmjTizrroygInynngdMgmT74ou4QqW9bVoFcOzogbWJd
dzK/BEfHHmYdUuCL/+jsEDZb5TJVPFGzw8pI46N8LBs7+xelRWspiDmlNgZvYw3scuVBbcPoPVC+
jhJrRh7NafAU3A0UtbZL/V7Ph/zbh8WVUk6wMsdyQcK0szjwfz9fQdO+cMEYzKLrTRgUw04JGSys
1dsoI76mSNqGGdRmnibmm7MgjrXnxZYr0VTLzuLBmZVu9MqRKJ5q1eND2Bjm9AleBTaAMJan9V6y
6m34J7e1ziErgxFP3orzNRlzLw3ofLAas+RbrNYpjzGq1hymdyLKnfrlGETBD9heNbjU25fvb8yD
wL2CTAMMAXi/xAy4b6zCb//lDjLGkOxGKblPj3y803nxMDrnE5pKayS/FBe3Fwr9oKvB2u8/Rl0I
6j/LZAWWy2ZtI40GOqCMSVH3Wy9Pt+/+KWgPLSIKWfvaD0sZ33qR5Nw2NbZBMVbDOdQ6EOAxGvh5
iykUbOI/5PEgtdvJ9GpPJCxPKBNKgfihgXrK3EQEcAfH58mhnkXVtSw6U9kohNqA84rB5wPjKEIH
Fz2cWIuYfhyy52W9SNv6nu5X6kCuSOXQuVlDMzOObrxTISGeB8SGpb0PMqLPVE76huNQIO2HxqNl
uiA1b5y37q4I5tw2lu8o9JN9Z+AmrhHW6UDtEPGCbrgMCRmAp8Kt/QkRlDwK6/QgOD61OJj1mP1U
CUBhdxSTSsideUPNKU17l/838fL7hKCdY4dL017Oh8K6kdzzfsI/vJzZmwVVC7GSwN0blRKZYknU
fF41m/Oeq0n1XdA29GGzaYuz47KO9Dodhfdk5geBbecChbY0/WkQLUWFvJw4aVJK30KPCngxxAVf
nTpqGnWpGyBP5U4jw5pNX7mTwEPqMh9vdTerU5p3saMYaiCv53xnrjj07ogp3/rShS8d0ZNqTZJO
sbrRODlpwpHe6A/GvVt+cjRZCLXKYgQ4fz7j/zgjELpWhK00+5QAJfeMXLDZlCe7R2ENpztE2xsl
OPAzj9pI5zduRI9t6daT9ta/T6cBQBOEF8qrZN02qLcqxIv12PFBd0AWmoooaC8TzYjNSTiSidFh
vQSo+B63eJ2snVat4YNYwnWpQTLBcKbZKREBFq1KI42GITSkBQKcB9RMJy9xpXShV7jxwHbrbyTi
rYATkI7pB/5CYlZ4OZYobvxLGJ4LzgfQ+Ykk96xxibUfNtOeXNOtdy7jxEwM/oYhEBTs9E3RBhXM
S7Tp/1rukQ+8DwLpfrZ5vwsaTfO1mn8r314nPEutKIx1uUoYcT706uVSSK6GXlr02VuMVoiPu0iV
rui0ikJr9mchQ0bstPF6WkvG/XrmMiALAOp3ee10ppN49eWXu3JaIA3tg1/TpV30OJSExuZfXfyf
3NadB5VBtgiboqre/A2CZuLzV1SRS1YX95nIE3eG6r3p4EVTT0Mw8jAbqxZSrbPOQY63H9VbIRcH
pOk6YzbdihAbdmowIpF5wzYMEPG7HKI5l0zWJqaIUNCUnJ0s5hJYOS/VdJoqrPqMIca+dAJNYOil
lS5l/xj0KanbsVtMJlkXPIiHGlOnqyvrbzbqiUcPGrBZ4YSKbLdN1erzieTGqp4n0pbJGDWXN07u
IH15X79vF8PxpbT9uROuRsYCvSh9wtCqDvMqEqZ79Et56kXEms6hDanx2+/VVtK7mwP/lQaceBzU
c25kCPs473IN6QtU23SL7vI0EvU9wpnagtDiaCAKAgOtMU6OHAVKi1JB5Vb7LHeNp9Ih4CsoEPJK
rB6nGW6DVxYQ8jIwOISiBen/DyYKBlDvodkPQ2hRAXZ7xB7DMTpi/BOyCckiBRuSrxmBeRubwlcn
5ovfVsnLHQcsabJ4eOx/oSzKttEIWbBaZgVp9Wt9g4pdd9A1tLp+cdZOqMdY2xsaOYyK0utSqcI3
T/yKwZecIVnMP+1J+D6XUyQQ7FPlVjQfNj9D0AuvDNrijEQ5jbzzW1+lkD/mp0g5eA/uAh601vqO
qXMU7eDK936mxeGeMmHrpAD4eHarvxl47vSron9S5gDDZJvLSBEBeCUXJxn3z8HCJMiA2Ijbp6Az
daIVCuI7WnoJ/RxCPI7isdGYnHeo8erNTNPMs5aMbl+d7fMPJqnqWNed5n3XiWl7430wAMt0XU1M
B7jGrr+/2gFkolDGKr7zAkU23jOXQ51RZUXym2Oic4TFEn9kfkpMpmmTvcDDH/i5afJKHkabER7b
JBbi/ojwSQ9WeMeYhuOKNnhv7PMJAIvLGAgZLFTagsVp738mqPMFWC2awany3pjHnXwNBf2swPl3
SIGYRfIrD3C8MUjpSPrIoq/z0Fr28nnizZHrweECquUblwUuoHemiGXJSrKNHPI6cZU78oZJqnp4
0ysOufOvLXmktjpeFF4E6t2e8gz4SkYSmfUKFJCtRwTsiqbOy7f+oGXQfAPdXNo3R3sC34viJE1c
uffttdFOTVwTKvZA5jf6tA4HzpoHU+L+acI3td+7HMVho8zTnDk/NOJkKHrXwdKrW6K0LnHmyDEd
vumrP3LWGyLF+xG1eRxiZBSAZQfTQFwKJBkLnh3ofq9Cb6dusG5ZLUvnq8WOK1Z2vU/7P8+YNpUb
/MTGPXdJ+LT2nrP9/w08kWuLIsAvYmPDDz60YtCWreDRKfVuN5cXVC1kFaRsg7QgpVsUs1S5029o
qctKwVzsP9ulffhVOfTfGcVf2CTXh+ZCOBhndP5QxtfdrmuRZhrM12U5U+KIaQelbaWxoVpBBAeS
HT/icE1HHmAK4LGvY+HOWDdu9QizY6narQN/ksUwM6s1wMzKT7lm6eifQ3VF2Amfe6fugloXZuZO
3kzqrK6n5sbU/dBybCwGJ6sxHnfOJ8gFmyv/yKInH/Hb6n56SIYfs8SLIGtTL3AFtaSGQSHSf6IX
LYercOESSGZkY9ZUr+FvQazsphkTHfuxgesJ/Ug6hhg7MMq2cYafFmZR88Swe9xpKW7DHzAPIgbr
0B36qgGBreTOZwNZATwwdn7HagfTTw5Wd6FWJf0DSlr1agxXXZVfRzOIHGCjH5NPIPwWKWM6hkpd
4X6N7q3JhSwj/LGHg6u7nx3xo38RZWoRsDGlyqrsLzYrNdyv9JqlYbjONOi7OtyOlRs2mZ9K9aU4
APn/9h6JRHJsAZ9WFox7kBK4ZAnPwdRr1zj3GbpaL2o04+awtAiWTFlJa0sz83pCkBwHBzq/983W
uZw2tKyhJxTc/BYoWFCakG4G4867sc5Pq9s/Y951iMaVro2J4cn28OjiaLSBDp/inam1cTYTlHUF
XTntVmfJ8pu8lrBVAIQfGrOVmCpjGd9NJekydktzWjfL8H1envikhMYC+rxf9Ug/xHn7LFk1TlHN
CCIJBhx4dA/+S+W32HIcX5T1TaJcVdDkW7xBgjnTvcYGHmQA5BP2UTJzAyLICFhj77lE/jswfLaA
tO88lrRHMPkImudTjkm0c6slkfZPlmtF5Ic4uf90B6GqfaXF11bw+xSKY71Dd567MpPyhveCNBqS
t/X6I+DIlsmVyCzETmuwXqGiSNiOHWoZJ+GypAUsvibHOvSp/sWQAu2R8GzK1nhv4xDa2QbMRm4v
nxW8fz08hiBvfwUMCq+apzoZ+wgFV7BYylvXefFVwo2H0984H/JPH8J1W4Zl1sgF0v1dBtgh5Wlp
avw8TitMVF0t6r4iCnhZ6M3uEWlCTWNn5i5CdXIUun3iun8nc2ezgiD2t08DRkJ193ngyPCTH4wp
klAtpFYY3Da8oBzGBAKgDnZmCaihMc9nD297JTaeBzKRdFbslFOdk5xvB8a7gf11j9l3BWiTIdVR
YsWwubp53FA6MKAb/gQ4e0/mS8PgHitQPYFOT99BZNkUmWUCk+aiyDStejY/MR8PDl4QKMNMzi/V
/vlHwFQPnBLWWzQV+RkWe1d7jdhuoXltHIuO1fF+4O5LnXQ2/5YHo1HOk0XxC/H0pCaYQYeY9p+E
5FKAlTPI8kgBPiLt+3N6C6Lxpx20oQmzFyrEq1UQzj9nQEeD2kPjfk3ppVN+hR/lZFa2IOF78Pj3
tKW473l/iS+qoR7qFQsjAyvgStEi3apscWjgz2n/DrhCeVwdZ8e8CKXK/ni6U+eKbHGhZ7kgS/Wm
G2YlWCQOOajwP67xfbVRjkii2DY39dXwB9HtYmTXOmcQ30vRFwCrfzv9Op9D6zAACO43wCST5YkX
E0YzuK4+HfNDUpFhjHrgkEW3KSipDV/krfFCeDBJJpcwgEJ+xyx6RIv3S/FWKkcniCfo3iHAGjX6
vBedx5IfAHT+YZjuwF4D0YX5uP3802RKpUmyAgMLd3OXrnkF+R3YJ5M4QEc6A7LDJkFY6gsiSgV+
QYVltiuKpKKjXqQvuEDbfsGMRzDK9LxsSCcecsJVKE0AMMo+8W1wHvquwTJ4CpMajzskcDwYyevW
IdpSEb3urKocSMgZulC7u+nHo8Qu7FB/c5wifSV9B4OQ1Layc2Ya4/byZ+nDkTRYPj0c/Af0efOA
vtuonpdXFPscGh6eQOZ32PtyEfJp64kcNWOvxVEbwl9dYpCS+rmdhmq7kCxgBNZU8acenrSHoHKV
uMNoXMMuGbabUXb3bXCadWOpT/cc2VYuLUDrywRqUicGzVBSz2jIwmOrgdRp0GlAmnvBVhCrXp0t
u6CU7XofRBoZ439r53XEEsvhjmkYGwuF9Cmuw7vPnYST6loqoN3xqnClByNJVRstdlaKB4CHZlbC
lIF03iCa6gcDHhIqvk2q0Oq3H/+vfQMruoDjs1dbPiUFrKYbQTKGn6ltcCFPowv23o5krNf5pn5L
IzED60gx9Vx0EtVKuxe2ToqZRTgnL8NiSagMJsWxMzMMm3JI7XU+eTr7D3WthfpwYVOn3FHPdaYX
CBLcGkj+VkpthzCDOP3MqvuMqzzKnBsUXD7l+hS2FK386jOL8/ZeroRQy5iOmPj4VAWlLNrSSlq3
pHzuIQofTmj7F0qEqBSm0w40P+/h/CxtSq6CF7qxnKTe+08uBcA3rEUPxAS1NJraEmWhKPAdANE7
lzatI03dHUUWKMX+RouJQDPrfKRZtxi66dp7T0p3HP1hAehCNQ+nX5BJHFW5C/cwEK7MCIxXHO19
gWinRZbwx0g2z7cLeoXm1amAYS0mGC+lhea/hN1wA3pV7xGG8Yx0lMG1rMU0Zj0kQ92oQleYzctI
dJgjeyMiSItYtuqiPKaDuuMgTL2PVOtghCAwuVjZXaPnWURB26dm+LHhQO/SNtwbiWvFZt9a1x4e
/uQlmp1MnN5GqbA75M11Opy2ZShUGlT8H09uyYCLY4ewgqydvUaouxNJlkygk6BHcLKL0DozjuM0
3kHOGIkro758+uEF5Jm+zghg7dlP59Dv2EEoA3qwGNo8x+wSHM/03oAFnRcXIhBNho1QC9lKaULH
DpwVY6xrRKTQcLnrsoi7RRAvGHB8PXs/Jjov8fNjfwctAqp72Z0dRmSzUePHSrefF/gV6GZ4PioP
SoKlQ5bnkT6GjXIs8R+EFGsA5KvBYvuQGn/gsK0NdAxXseCI0bV8fis+BtoERImvo43t7vkCAggm
15c0Y+p22fjXe/eOd107BZkIDPHNlxQ2+h7nL2VZTY9lqKBHqK5XrGt2g4+N6AQtleA6ryV0cw9D
vYlUuWKB7iFkZPeWsSmudFxtL/N4qo/9vHE1XStALrji1MeNOzpY0JJ0+kvINYJEc2OlRYRR3Cqn
4ZRyFrXV0OiLrZez70vFfinhIA0+LHsUKiFZubdnVR/rBemzaLSgpv/iQJ4fUo1cILjg5+N0ZEGN
A7jWVuBTJs4jOdfCNjPk5fPub3Y1LYcfrx4oSH5j5oz/lWMgM1XE/hVD3XV7gBoFOKEBS+r40gHc
uRVBnpiTs4vCPfWWBxQbIlwOFFNWO6yKpcPgoOpPcZaC3I25dzJBqTM+n/XUJXsuQb7DFCSWLvI8
3xoEKyTI07L/uvr1VwK5t9kwbaazcsFQQ+NVTeOYiusZ64ryE3cusungGBo6Uk/zDWIQ4hQxMaVO
R7aqEUwcURem0nYWAb4fRsLHKhE0a973E1J9SgzjzfBkNnVnCvemlfJv11iPzTwFrlwcOnBCsbsg
/pI/W4elU1SKUHrQQNAV56ivkPNTLLlKJqusvpGYsZfetURlJiBVTa4cW9KqEHzekF8PpuDAGMCw
x8OsjUQNg7Vqd8lE1EbJtAkA6GHE5y2VUSxOyxrreokhpye7N/kBVILNqhTbqsnr2W5s9KW6kyuD
nxtzj9+e3+Q03iJ4XBSALaDo613iDSlDo4oJLl0sqi2waoevjRimUaqc9rcyLH4j6fQyln5Muic8
/ElVWpEBH+EsZ/HQKzS3Wx35yugyvsDxqTBU7jAjc7sgSwSyqo4JKE2o52IGg0Am0CCog5UvQwxP
OxOju690Om8Rly4WbaO7+jquw+NZRXbtnH2IO6anSJH4dxB7yG5z1X4dGukZ8MnFzLGBGXCEc5AT
a4qilFtx0eflDS2zT7PQP/y4dWSpTYy25hvb5aF8jYGcDuPhVYbB1+ojW0DmeD+m3ipLzFD6ozL6
39XtZ6W3koR3Umft4ZAFLVkVnnHmnQ48R/xHXMjkAuZ+j2QXek0qNT7mVRX7r8NWGoPSVGctinMy
6mU6UK7HOIuJU1qDXoIyCiZSkizFeSQh7SKFNzQRREXck5jBhRHoN6hjkrurqVufDtjJn+yUoYkM
xpVJj5sXfV9hCAYmAFNPn/llLTwan5jU3phTSdP30lMztbw+9L/HVfFWtc9XMrZSVurUvawWo/zn
XdiroQBtaPjur39wz3uMbu6lagWXf2KhfM18m0JTPpEZ6xy90Y4/xbiWY7C+0reLLQPxjDGji9si
YotZyYGNmUQ7iWfu6Em235PLiwLrA0u1ZJnEhWGu3yt1WUvWnz7V+FL5j87L9HBdf3lAlO0eCfYK
2G9fUcThFfcDxQKRd5YEOQUVpC13L2HSml3UaME/zjoixzqs4o+yiAD/lDSL8wKvADAypazQ5i0i
+cXfj8SbdTj6QU4mgMPuchtX2Ll1tt2smL/iojGUSkFigQ2OiLjJ7RHxTc050JUWvBZFqbmV6QqW
6buWuxpgRKd2QywUdGs+fr8DxDwtshVgnD73QUjVcD21Wd5oZk4Grk6hiQOo4FE28+R7FOXtVV+Q
jrKE+aSkO2Jwey8B0OGrhkSRXFErMTyxHxBDnOmnRydXBrjDEZiwxse2thXTFIVw4G6j4N5AEjA2
rwpB2zHNyIoz1RTZ5TOQwdrynWRTu2RX0XwjNpAQkeVHCcmuKfzIk6XfEUbsxUxAd6lkxG0F/9Yn
fSQtZlXVknCVymJIeCu70IHI+/e24+2mW5icriZ8CnZ39E9569qFcXMFdhcbiunVcBR4gGL6vu9B
CZSl8nhePJKuJJYGggWjQr9gI2tG4E26REDXbigw5muhjB8KM1ZE2f9+enZ2W5vhzvjBkNMTR+6O
woh0HFDifLWRfjfZAzv6U5n6QtC62ou3kDxt/MSq4JPc8HZj7ngnfx4235/q2U1i87Jt9ha1KO2Y
g1HXJDMlBhx32pd5eQzjTwlu+vJwv58Ru5PH7w/vxT0HHnePaN+ubD2f/akr6iWHDiBFwJqdVl9M
5S0C5dBg1QuYeZsBRxQh1BUTZuqdFPEHUZ0vfC7OmLgljlA4+yR+rXDFYj+ot7VxxuoTTXk3brOQ
MOovA3SRxxc5Xs7mJtxspt/ZfxqdqTcixjCRc2ZSJTK/vKadHRndLjrSeocFekSg9IAJkVhNFux9
6wGtQlnlstgHrKc5exfVM2+rNBcS3374yDtooLgIEKGaxiwRJeoEh+QeT2lYKr2bBEqBFWkUFX/t
r6VyvFRVsI8l8FWrQH+XTW8QXjH0S7bJL6B/mKwic5/CWizUbeTjbQR+rXho/dqvjovpr1Gf492+
smefnRtDl6y8gmxbnANdpKY3+sP72WuqVIAtKKhHmeP6VBKJAK04AqR0xMfyEXT56qO+X7NVUHDz
ZG0tbTpvDH56+Nh/inP1b+sIqbupCj+XV358CdcG4v/R2nwvwDph5Z2Ni7a+M+B2X/DA5HaqX8N/
oQa6mmPHLqYSJyZbT9f7Bhqwf384f2NgPZvHVCT2ZR9yvtGusZGx0L9HorGhGDUbwP0LAMELZdqQ
MQCiBvM/uxw3PcjEJ70whevhKUHDRFi6Mtxo8c736HDM0naW22CK9lUoTJC4LX34bJ4Kh0C8W0lO
/wGqo7XhMwt9Hx3RWqNuYeJrHGLlwcGllkjfDGyF1GK5H+5q14LezI7bYPvk3KMv1n0OCiMc88B8
elINDgnY8nEYsAjzi+Nv2s1RWFTaBwdRWj5I692GprKaw0bWjXtPphtSTFHVByINDQeA9/x9Ia1b
iiAmhG9a/o2j6rRQiCLQA0T5o7d2kxXvcnS62l1sFVxS4BKQtZo269O4qyQt25Rru6H1cQligR6W
FPC91dMi9lc2JSc/7N11DfVVNYrTpzaPNL6G8EY/7winRA+TcSyBCPDg1qN+DFqutoj4oAitY9ur
AHTlz8K8LDz9rjwA5jIDg9uw9NNL9Ntf0c/ImlamLCNfIZ1RYL4f8E59yGv2FGZnZWKWwksv317E
Lwp72YUvSbLv9q31eb48HI5R5ZKGr75BLktzyF31jBJghDII8pMEdSap6c4myl7wIEyZpnG3WFAU
38UQLDuo50QQKAI0lD0cmHtNDyNaBpylmcxqU5P7bKq42Z9uVFllWYP/RrI09Bq2uEHTlCuODVbf
EnFBWYTKYFretbX5XyWHtjSCUAYWaApdnK9rFtYAGKmSJJU/3wcC6KOiK2dveXLzOUhPSYWtEuqU
07+4AqD0MH2PaoNpDuukfpDTRg/N4PFEFYfkn9iGVJOgY2G80dlsjsusdd9e+9mmYL7VqdAoM8V8
yV9fTlm+hLQUFWrIpGz7DkzB1LMWIs3rN9jjgvhm434uPl+DpWXE1x/QD8aPQxyLbZFma8Lhvlke
HvyYu8N5QYGpeN2/xx8Cm7+RD3wg8Ai9JQVhGGUuYHwFSFfnjfJxbY5rGrgeTZpyrJKGm7JwXEtB
Kpv6eTW1lFVKbyAUot3TnSf+oCQM2ZctLlpMI0FVnIdF37+FJSPmySrQUFBDX8cNsuinDZV6x0jm
wkH1XO0HJXW8jZCBgtUoNaZ9sdY7v/PBbsjcV1bq35BAY6rEi9Cs2jfjQPPqD6M3hfFD+iqA1zwr
GgENKBlpK8gQrSsNnO8XJKjapKzutQuFvNu85fLUDyA+RUKp5dOL1NZCv7ND8llrDiplp7JPq/ki
hTRD5H5r2vpxVjVS6QBej6HKSDnGCfASo79fbHPmH4SZthF1dscAzHStmzTFo5a1F7uBjN/+RuL/
XADt5J1PsmFJAk9fEwr3qmR7gNdWJv6oVvR2kWiyY0amh1eeBr9Hhs22woh/U8dnzCGVuqhh8IO5
Mo93haghdacrR4+FUiJfyHadH8XYmTbvqZk03Gtxh8MAnTZLKiFRJKHVDdRqgiQXCofaPDdzRDP4
bP9na/osHZvAbqDcg9mpAm7pfxwI02T2vEq07AJoiXrmqLYijs3GMRZ64rW2fjnmQ95ciX93WcYf
+X9bmaYn8LtmREc45WlZjfy6DBiDH7VYcIk+vNRBd/SuaPlG7yNRK/f6j8sYCVarctCT8JFFLcmQ
5RT2aSF9U7PSvA8Mw4Tq+Oh/c+ExPYtASE4VfzNcEglMIpDaRA2UOCZ3o5jBoAxp/XihkREFux4N
M6RERU7Z02autQnQ6kF3pYavDfRNJkRsVC9kixdi1wgOToRJoMQFj6WI1hUI11VKUP2ZX0BdV/E1
p/mS9K0f/DdJQjm+vL9Tt/jm3nzYjevZNxR/nJz8cgsVo5gFDyZ+ADD+IZESv1GDULwp81YQFYMr
6XBsrcsnJDF5LNpvXD11qVkImAUOPqO0cL7wwAuCIHIRbDJjQnZRPZFBZVj2dNMP4aP6qcSyp8Hr
QWnRhZBRp7pXB3qgXRxR9RrmcZILsW43oRWhbPn78f2C9iIIRBZatb2PsDJJvSz45thagXPTTYC6
C22e6EQJ5QuBonRJQlJNynBHdeyMjXYbYotO4zkJCfi3DUiS+TZ3AIqeuA98dFmRPFE7TxrB57h9
mob/jHViByAH8FPemcFaGXQ/sijhGS0MGYxdfmKLeVgsRFeQcytouOZzMBUX4pv8+FdgJY0bnzak
pEbnsAPzh9jXUpSbJXkd7kM03NQboRnUqDbnj4OXX6+muwQFxZ29/GAdhC1/tiEdn/i9HYxqdpQA
EG+vVaD9nEAcUxVExu+nbOzWxMfm/GIxah4k8kGgjwn98WAoZTGCfkQPQYsgvkvCXxtnj2c71fgy
xGmMSx/4OfybJ9dlj5DqIbJ4zgjtZ0Z9gdKjlNzU0e9lEMfSpt9CJ6qIMJ97Y6Dwprw+/GMMNh2q
2FM3IfvfHhCw1H+Y4k+FyowD4H3pGEEhJ2yepMBYUq47ySAkRPGVMFJQziv/fyISW1e+YK6nnSNW
UiMmLSD7gl10Gu6EcrYRYo75Gkv7AnRYTp/W3uwUP1EQEDi6hLOD8azgMZ2ezxGmQlO5vr+Z3q2h
tXbdtdSkHbIYPV1TSzjvTFqX0w+2p/F8zSZiKTE6OluMQvirAsWO3kMNBuAXX0VY06kFzXjTtzmb
pOsvp3pHA7K0jlEX7dfmiB8fuJ6Pcf2mOaMIjipWDGx+VYGTIjVEV+LJM5hi08coq61qmlj7ebNF
tSrRHqE0NBs+/1e0J5XdJCvFL2JEVOUroQzoxnPJ+Gs9zp4R2VmTVCvZzVTKWIlW2VYqhq8wpRyr
KXVfAKrzvctt1DeElTv4RCdGryBMp4Lmq5X2KWhwfUYClGD+2EjRbzoSDvj+ob9y6BfcKlQf1opX
ouL8SE/D9levkGedENg56qVUzRsR1VCFTV1sKE8kWemH34UtMakV1fQ2WPYGmwE+cary4pwLUJJc
9OWy1hYWnel51iE1ByADYO5Xe+oF4wcuftgAj2QzAQdQlTdBJPJPxghOOcJNoRImkHjooafMGF+g
hGV5msn/mfYQfKr6uKq7ch0uu+egbM3lvtE6DKLDUNuuKI1ZWdtx87ccAHIx9M+3b91Cb7q8q808
bGOVYnzJYNu/JJxCZstVOjka/WB9SE+awfoIyM4HOqpow7JedyRM6XGfCosNKzB7xvVbVKX7fN9r
gKZIITDM/qNoW/j3O9phE4004laqhWJKE96+qMUgNdJiPf0tkIJMHblArIi5M4G46tyFXDBAmFaj
zC2ilbRZhRvQMgDGuC6XohP17acRd2LfNX2ksvWateO3/F+h7d3O2N8BKxf4/nU1lLPOb/WPa0V3
+v8kObiS8b2zB8arJPsn+nw4FBvtrzpAPfNSIBiLf+mjrxQG7EsQpIQL86h0MV3IaBEC/tVqbDsa
dmR2z/wwCSkB2kJYvAD7AXzFChEza7IOnd65poBnU2mb3wm1AtC3RxR7aYsBUh7g5U2qFmHxtOZ8
D8xhPNspeZpm/Xcfd0qrrK6wXQ4kvQluTRJPpXkL3czXFP44UL7bTSJZCcRaBW6q0YHzlIpLShbz
z9DL4M2ji9AjuIbsvAnQHl/soVh2chYEyfhhU4VZmrCxkdX0EodzDYuKGNab0OuuyMgPSpUlaKOp
mfLYrMvPp1X213CvU1nsOwDVuX4XCHa9VFXYNugBkd/6YyeI4DAcGb6g87WDDgieGhj5KsqisyCp
FcHQX7dEdJQpg6zN44tWPph+5lfe89pELxN6lxpxBf9dS8e8UWybkJt6sna92lSi+8BG6CvhUf8e
12ZgyZQKkVtlRG6OV65MoOdJLs1OlKSbcVZwaFFp6rTTp+YC1trYdJIYKiCiKLg0CuVgp4ARAlHt
bpwImNg8CEkDT+plrJZl/saABTvGl5DeQBI4jkQbjMragH/dEcoCIGhwgM0tiZkWaKzF1Mr4ALdh
Ms7kz9Qcb7GTVLpqrzG/kp5p8PAQDZsomRj4tVPKHm/JU3FpKmFNwNrA5Fbf0wL1WnzTd65diDJc
B96//UMDJRawxbxk7C041vZ/yQwz6sEXPtQxJi6fYzT3reWrPBVI4PvF21Vdm6X0GHU8pa9bzOqC
zMsSiRr8R2yGxIauA4IhisocT37DARp/qKyMwURHFIfm6swhuyQcALtF5JcwEIPpb7GbvMEISP9y
XQORPZ99QP6pth6ul7Y8k3Lko2vN0S9swz//M8DQbnhtEbpC0pkylcBe2rb3ESyxm85HQdIOzNwt
wPQFjRiJu+kor5ryXqUzAZ8gtCnChrboUpY4cr86ByN/cQvNwXPVUHEihnzLRsKI49oZDZtaa9ai
HiWwek+HACHCVBOzyAF7QYIW7fat30n/ORvuRfPkmybuhWmWeDsNv0W3pcpkJVO6G2ARQ8E9sN8X
Bwsh26ABPq0WoDeS1DclpBfPjnhO5ccgH8nFPU+hpSLWCdn5vl+tXxMVxfpno9cWFVCDA8Kk5VxE
0lXBjT9wvaoLGY9w0q/1O9q73BV1mLGILVb0e9zn90mxnTA1uphuRhIk4BmgEbrkcRzf9sm4yJlj
2xJhzzh7EQSHW0cIiVlCaJXefMw1PZq8CIffyyELv1cYJnTKz7F77sopJJPojlZKR5IjY7w+rqT8
Vu/4zt9ycnFMUOQfXl3YEg8xcIJpmTIfc+PTBqXCTQN5fQUrlNsvGT7rvwAnW1rtEBpzmU/BUjnm
EHT0exf+1XNr3tz/M5Fd7BJLPhZqZNf+gwdEzAcnLfCCJ6ZvPZQfu9zKkMfniKzO2F9+33/PKOgW
GlO5mK5c2I7FI9ZkQD8rW6X1iqF4/YQTZXmF6I06Hgi3zK6Je8sMdOFFSqNf4zkO5lfVIXcstFtD
sVTX3Crimfr8mNMThAb/z6MK4Mnh9uQ+b83tGk6xQ06psCuongC3uHyhiXSAm24UTorsfw0JB+sr
BSHz6udFvsmExquZvho607tmLf0s3asF3wSZiMJWXCwNxvKM+p6lTV22DCEVwuVlFbiYFRgBzjoU
pjkwS7jFuZrxhIdh3XKzaBpj2e8VuWUFC3ifquDjndJBBuzh/0NZ+FuC3/fNJLZIpnF1VuUWf4EQ
frFc5uwAYrbz9O/RguhaGr0Q8wyyCyLsS6asKivt8U2t01SnhpIVzNNst7alZJpdlH477clkkcSK
5eygXAXTZWcOoOs/XoIQIhtSKu575HItp+TFLMxaEVckyP/Qm9gWP4HYq6mw8YACnSqHpwjzqs9Z
r5tB5jPC5fTze00JLvJWfGv5MX1xZfBqMaUc92YKp2gbqrNRj/D9nQ2B9pElisTRoUHjO9dswntY
3JSy0kudZFya3Q1T04vowkyDOtJT905Bg2Jlos+jxNbEMSFX/C9Sf8DCQoElHBshXnvD9RR/WCiG
1vf93Q599Ox+Q0XxKQlrx4ccFXnagg+uqRSmQVmU8j2c46GNSa5hIpsXN8q9WV4HS/AKmL/i4e+v
BzKQItqxt716ZPWcr37i8P0w7ofhW+uJI5PJjJrRGMlaFqpsne77ecoUBBrNhfaPIyfjw4T8PsSH
TYPjQVA9i3GO0d4QXHt1yci0LK4oaFGv78oPOG/rqbJiep2R095E/FlaJL8R73TlmFRnzJrEYtBy
fblGWvmVPfh0NDmxmncZcB6+l1tf+x18wO1F4U/zUgRm+KA97xGnP6oVfbzw1v/e10zBSLYbYBRN
be0Hdk093DPAQEwoHd9ap0Nk3SLYY8k9GxsVLfX7qtzmD7YEfxE2csYcUcAOnnsWg3tsR2HkCOW4
xeEJNFFpbdfI7vLxG5uNogetEEI5A5IdUjlH3mJDP1AIlCKcFoBw2nOE3n4VuvdJt+q+ikWK6RxE
7fqcEjT8PG+C5BU99G9OO73XEDFGHO6LHpck2jy6Xn/PJbsuVAzATP11Oed1QJ8rqtPXWGF5+aAS
FJ1YLdT2iFrQp9UWE9EWCHAXnvpri1jpJ1njCy7YYDAKkTcFy8QxT50MaCNHvO8nhYuLAat+ulwW
9YLH2hzCam5dNY7geYe4oK6/OnqqdWM5ZwXx8QtB6sVjEROgBwinXhLIwTnTmvl6ZTdTd2/DXGLi
9ZWU4SwyCVT+RpcIXrdlOTqN6yM7mOUEjqrZHy6JnnLw3QwZQYXv8u6RionCfQCpYBBUqLe3WKct
Xx1UcLyRb7o9tPrUxiTQO+WDcPm76RDGv+PRrAyuBJphFUj4XAjwhwvkzdFvOjxMP1T5KARd8YMY
N5ZTSsAWWE4di90PvosMn78ELA6bZ5NkMy41HRtTdyHppX4g6GcxaCXnzT+kx1g6AKwxDxDgE0SJ
aoxSoc2IO3UCPXnJJPmLxS5S18+UXBaUXQxzlNsBsV5GxXU9woSOyoWgblQr0yVcCNX0s06QcEvj
cvBxCsxyAyoJldQcCa+oFWMfQJmAxnPWqmwD8vhndU/WgybGFtzYS2UO0T0TikAgOnrC9HjC9CiT
jyK0C+L0HcUXRPOdwQ9AHIlnmYucEZbITKjUiYVw1OiAX9al0M0nPLHH+k7qsJzM52kw1rxVUsWr
4lCNwy7t4aFGhRHb92ZHyeJ+bO4y4UM85gpMv+o3Ps5u/JtEFeZPQmEDqXkOl7cRo/6+0Nb7HK5b
bTN3dnyl11eqmM7iHuFyqfJHax5cJlshbpUmRhUUhtD0HIinRRpFGkmWDZsW5iKBZr0ug2qrljKZ
XlzIUcnlUsSPCtdKWL5JaSn8JJ2dIqT5WXaJfEtHyxSPy0m09V0QOn2KrKLSOR1vJdBlQ16nvsLC
uHH9ayqsM1kIjNf/VfFSTcDKzFB/erIQX+hZD1X+AY9R25wwVleuikUBSTXThOckS1GNZHp1Tgw2
oEIOuNwNpaG9/FHmvmxiahtrmHkPcLqZzjBiDn7ywGANA/GzbPKR1FVUucCkqrZ0wHME8g3bREF6
f2yaD5UxXvSIUou86mb/2IwD5E4/ki8nOrhppC5NPMLuKigE53l9RjamPGzfDcd6ya2y2WwdYm64
JyvQUD1wgl5wg+BPMaSagDUG+CIuNnR7dTUdRGjBUMOvJGm7Aj+VdNYaDQByrZLYxgKdzG9IndsK
GJKT3AM7ifG/jyEpYqY7QhGwISOHWPnTaGPifOv6DCN/il/cVR36XDd7Y3dmESUzX+NMCAon+PJ/
p47wRf9kJI0rgYdDybfxpfpZjuavxbuXv94apRp779c5iYcGXMs/u5s2lHPUHUQ8jL9wr8393LWH
POALKW173cZV1CPIzmpO4tGUkGCroOHmAovcZQTB+RWk0N6MC38QZxMyCtY3BqOXDEw5XNYM/xlI
eBvS5TPhJScjAIOaRzsw+WDQcczmVq+98o39ReW99t8VOqLTlIvw2siGgLfNbiuEZcfLYTn6jyKz
oJGVPp+MGcSkfb98AYYU5jtKPGo/aX6/k7WxH4ArHbuTd8k6Vn4HD1B3wT6gl8qaVSTSTyEb9UZl
0E5cGvPCbLNVbKoQU4pGupA+YSXrPQQRVSWNnZF43y2yI5/GFDtvVyl9MctVkaoJWIvgZh2bu87X
XOJxQT+ezgDxa/bSoBtmKchouTlHqlujR7UNVd1JZDe3QyAKv7PQmH+uI2mdjuxHMhhMyzKNUITx
iAmEm8wMy1xO9URt9GbfUBEAa9dsrrHNl9UufqC9USRRpSce8SvtXBXlUepf9JB/6hcRPPQ+ci5n
qNtO6rA9JLHzqFaWTSLt9YMH63J61at/iLRpubkbE3pdAZDGy0SuVhzv0DTm/JRNYdeXn6r6lH2V
NuP4HengaAV7/J0IaXIQw/2e8/Ut8QKVOAF8Fj1ktcjaeXEoyQoJXPn/EbsXYzpAZU9ba64xS4U3
cKRx9bU+phLZvt9Z4r22qlzoCfKmLd67Ir7ffCZtSU8W3PHbatsF+mpXceUeePndGvvr/AlNKcz3
O3vvWh0uBo4ikQmNHPVu69mwJR4dmKW6c3W7/UfrP1O6IX5V1xsvq7E+PDAIEP3kju2Dk9YP1zl8
WRAx9HzF/rdgBpMQTyx5SIaBQYOro7dl1K9ohdH9ck3g5ElroE5LIFUTAwXxTa0yzf4tDhMqfRUP
zBgYYcjjGkSzkoRjJ+4BsAMGF3Kn/M8xLPUaWatrUuuTIpX5nh3cb3NJ+YthqCYbFv+VOpQ7J599
TxuCqKTPnAMROY0JSL5kmg4SMvi5uyc40u20vtFPevWepQjDZlGQy1EaRn7EwW0Kplk6e3Hwuonq
XZmRF7NmkgRGNQw00Q91TjAjKiU7XS+3Dh9CR/ausLjGId7eMJ50OoJkouFi+z7Pox47UkwAB54T
WmxapGzVf5ecrmBBkZS6QcKLn8hOVvf8QhcVJtiGU7pmFv5f5+lGr929Rj9TjPk8TeX+FPbu3qVS
wJKrxpt/gMBnUhCfhI9gldf4w6UryznONg0IqZKdgAlR5OE08hWAPj4MsqxPGQ7DacWOZuc9/jBL
7oZXW3ozDikCQ7WyHntfVKFcul9y09Mbt+aZqvxQ0gM3xbSCmJBXVvAYVR3y13a2r3hpgZYpjFKO
uiHLozC9KDC2amP+GfnOgyMUQ14rR538cvXHB3RAA4BsLIRYEDkywoWIt8LYn+9+pGSQ0VlmRvGe
vQJX+OXWWpRajcyIMYzp7nODD50PU2lJLvQNgBpx836ttrhSMsTXMF6fBj/dCY976umMmfAMKaZ/
MNCai7Qv096Xl7rItJeCqUMZBwdZKbaaoVbtzZsXQKIOjxpIqStHntQJbtrDgFftEJqYaf440QsN
kNKv6jtmrlLKL083RycftzDCAe8utoARMeZ60YN5knseEN1XcIjFf494l7GBYnow/vtPTbhpavF+
RZ5BeqawY06ccNnna7EJO/3t+G6KIg8WkbY4eu32NVhTWNOIwd7/Kby/Wre9a+ktlevyLPtaHWE3
DErqjpo0iFXXiWbTBK2AkNsd/sDa2Pw0EAj4i01MrBAE4oClxdz8gHhg9wBTSbDwR+wN4RCPnAWm
S4GkF3vyZYoU8MB01gyCPHbHJ4rQ191Iemqk7WzTqER7qKCiYU65eKH8ukJLNIGVju9h1egvHo9E
JngJndG/dyViGy6A7MHGRp7IYmO7++0w4MOnp3G6VwzG5G6OzuO/8Mciu+Se6Fe2DrC5UtCgQtn8
6HJiHhQ8zDpfHMFbnRpe08fHckRigC7cd/bOzv/iQqkim03NT5CU5r/bprr161wiMLZ/xJ28DFtc
fwv12VcqVJYResSczJzXa7fkKK6F/ZOwYJHyXCbY4aZLQPJxU89/6kY1rqO3KlSkg3VjgueApcLa
RM2G8KiAffccWsGKNieZZEoIOZsEIP/LLd/IM1+r0BhLVDyrXJ4YJMjbqsAHJWx5cZ8u26QzsYv0
IbIAKCr3uWZzDlijnru+vgMoXgVamCK6o0/rIMo7B54jlCSKqNQyLvIqA5jfAYv8WSTWqMzIzh99
3CF0rmhM9WdUFfEziMdR2Nf+oMPEDAzNbFx7dw4aCF/eBuCtcCo7UQXhSd2XARMR3yhBEdmUq4q/
UesM1GoHeMCguAspo6g7CyqWPg0olI791PSoYjs571YVSa07UQ5449jsKc2fjC1kNE5qvbPdNgr0
lpXzAX+tydNPCMHBcVS8dNrt8P1u/mi8Tlv4+sfc7uH/pWD/ACqW46152RYRUbXSy05AWaaktzys
xzthALearH73A+xre/+zXHWbNuc+bUY/SoaL6qgn9I3/g4q1Kxm4dIRqQdcRQH0Zfl5ev1bcnv/n
XS/eB7ps79rAxUHx3nQLpLtSwKcLeH7AXmADnBOEWelv8Qm4grQ9ZWnZnumLJ20YRBXXxptbOUHN
05oezmx652fnN5c/pT0Du0ft9rlXkKBly1dIlDuOhZKVHEey4iTyJUJlyc0wYBxZ+9py2vpu+8pd
prgiIYf6W4GmmI9CsrbfnMsrj+XxluV6SbI5IMPUGZGjtDo6WhHs5gc6AJOBjDPji7AbILH3TUwH
7yjQCkDb8m2yrWz2q5lFuqa6SOEsrHHRLDy6GdnseBm2yJus2xahxTVppXKyDuwQlYCLJ9PnovHv
WGkVdEFRgqHpHtMu96TUklnkWfjyc/5Sqqu77YO60Bjtf6LqlEI8wkcqiNsJkCdfds0yVim1vi6O
IiE8Vl/La8eNdyzPBVTgGt6sgcUbc62Ta0LimB8GRir/oW7yFAcecPxjZPotq3JYi8VqwPTkzN+s
Ri/Yliln+qICTvyQU+yGtTEjEoFxAiiSCBU0Q2AG7A77sbsc3kZi1iXVXfNYsNPA/3092AEurlhc
cYA64HMCaSweARRKD/MytGGc9W2h0AlffsvqHHsV22K9HG6rpimWRZ9XuDJhw1/XfHYNrM0wYecx
V/GAVwGBqJQbfIu3vtotM3X2styc5hBM9hP8KX1fXQqP5hwBzELbSD+M9zsm1wY71zDVHhXrAwOr
j3sfEBBUByo+FHAhLb73wOlzm3XlneCgaNgOmpcXKsAe6RPQzgXPieSU8enZmpAWeJp1qcdA3ZiJ
v2vWU1dvUAAI062eiCq+TdHjLt2lRzJ7CH5HlMjxlu5yWTk4VkjB+zqcpd/bwHtfV/QBIwhXvmC2
UD45qZGpz3ExfAbGSVWf3ZfJfPqe6ZL97rDu/Q+XlBENj6QfQnJpqzQdGOwVJ/AwQljntEDHpvdC
hEjuvAwE4pg+MfynjucZe7zGNHIqgwF/P6+ZrljQilrsBrXiBAX+xs6r2UQKySjRNaZgSnEQXOLX
GuRRz+DFleR++OU1Z1hGFiun//XkqIRyd7iGmjjJcDxmbx275Tv5bauH7/cRA5yUhMR93IgFwI6s
TX1V7vbl8w9HHw/r6YTi6BlJBkhq8RBolaanFRmFYeJLVHOCFn58HhlSljyhej1nW/OkeiscnOGs
brrFzwRuXVuOFwnrIjD50vVvhSJTKGBkpZ76+B0aK2MGmXLZRNRHR6R5U0F/2DGvV6kT5bKCxTV1
nNcGMenfQJFx7erkfUD1zjPBvw15IwT61EfGZB+m3EsDoOyJIBZZ5734KS4NI26TvGQ30gBexPu+
+Zap1thjEbJNhyZ2ypag/d6iIPQnkBYZhAZDV115Cc6rYkIhVDkedQdg8x4g1rrzz/NYX3QtErI1
gViC9mT+BS+JZk2PVRcHh2d9+tNvyyBANSX86LVze0uigZnBEPczirLHaPQlmXq+TG/PncLeKUOD
ygLmzh7O7rMVHMIaJPp0nFUaYPaLlGZH1jPDgUjRZMPcZOse8LgrK/aNf3+3Wn8N206Tnw6tDyJq
7GlsQElB/zM6oONIzqDs9nL/MFHPQARTKcalEVviQ0Bs9nP6CDcPaCQtzQBI/Mgw3P0LMrRPp506
AMAWMtwtjUM69Zyqme37wwrv5Zff405X2y4FmSarKz6xN4xTZC5TYyaKSv/kwwZEEszcFUpq25xG
4zfGoxbyKnEbbB8P5fmelDDy8GktQx+e8d00JvXxCWV4vcvtY9QuPbVLjM+qW6fgPCadWC2nSYW+
ThcPdufrLghWctnQoyh3r2wYgAtFC9GULDrfvL3Gi+yXn0eOIJsNCgUYJXkMncFz1qDWVziMVUV6
E+vxt31ykQK2w02O02eNu/AxyXaigVEPEueBNwijV+rwR9zVVgdJTjS6lXpsvX28LRR3nN7Whhym
DvRsD4RVC2QyVFO1680QLqVYlePf/b0bMQ3H/6DzVKOkVfY96bAqiIXMzzRbnMtHSb3iVm4dhXcD
DnUTaUtigreR7bKVVmZaaEWkCjyaI8fpdK/beaM0E8ftb9sX2mbMBaCVu1ESLqJBVaYNU9TcvWKx
pAuB9G9PZPq7tM3ZL5WKhCWADJL/Gx2amEcbShn6ysJAJmFyuZakSHoPrJ3zPafOwDqPiSMvMQL9
vDwE3V8PyEtrUo0bOir823Xif7Z+j/Xd9lS9DWVlvIupZf8H6Ui9yXEYFbRsXLZdiyo6XUSCl30A
VgQKQ+yeP7tyIm4DaNbbVUzvlWBjj8F+0kXXT7SVi3YDU76G/WAFwDejLqU9AXvgKz9hNEiG2v/2
ljbabbr1Jo3VX/hlHkvCpGOdZCBckbBzIenPq84GBQgCzUSDIiFD8FQ2AfEcojVuBV20DA+UnZ3Q
ZVj/z2hnHXS5B8/JCo8HWzuxaOGlONyp+gsdX21Iac02kv9zAhccddQYi1b3PrAA/YvMULAGXltP
lhf0ccGOKZmO6RXKgH7vNv+cyy0Qg0ki4LBJeP6v5TZt4dIv8EitMizMsJHbQRORHjZkMR53+sxi
lySFTjKm5ESB0G/bL8WuECcdI1maXjgHNNXewX+wHmbjMh3nVDpfMjFII6mBqQ2SmARKspSg8Xw8
CphUNZIw2omVhq4M4uiVf+zHCvCGHtPSR4Cc6jsHmQPWI7UrGJh5tXNqZAwWpy+rGUTSZVr7FBSK
0NSQpTLA34cAKSw/wO/XpMQuwQ+V2rP73m+CzwDeGjDDMmG4Bq1r6EBLCYg9yeIodUzWIOBQHJCK
WuLbF5wHvJgEwHAe9hXE8obpqpZ/O2UnT3vBd69mBSzeowe8/NzQgVx1Av/2BYonVrU2Y7+Q/VMx
1xmh7BmRXfW3AiAucABKyTBTu8ZEU4OQdav/qJRQw4TQyDEy4t2u7g91exWQyr0ypxXhDX0Nbfm8
5mZ8rNEOzULih1UuPEVrSdCrnhEYbgyICcDZihur6uWac0HVC6ypIFCS9rMI+KANBqe5eVzPpH6o
3J0wEfYAjklp5TE6wIYSe84e2mcIkzj7SBem2rCIE3Q8a6LqZzQN08u1uAoRWREeLhVx4hdMZ3jR
9t2M/EBt7sBVSdYMuBX+RVhOMBgvcCel+U5FzFjjpb6kqzT48OeIxkNIUanPA97veIepS+Ch84AJ
Vb1i1Sp/tAR3s4f1qZgDz06mrAnjS5bmhgjEyh7NQlrvNYncOG09m9PgBfiaOc5DT35daVHcPCgX
2XJQhvzeBgBkXV7tGmbrsca4QQgmx5oKpfg9OP+BPz0LOaUQa2Jws/ayFBu0U1LNwqA0qWtxSzQ1
+oZtvv7lQjMxcy/RW0Huf62+iS4VPdovVm+COSIeicaeKo1ei3uKurw9j5m7C3vWrbpyGDUPImEd
ydqfxBA3twfDE2Z4IH5lXOclrxpyIz9ZSp8iYiMNW8EPBRUH3dSj4jGHJbjnCXAYFZPonDnC+Mtd
4UasAjGDdEe3WA/FgD7uu/vPe9UaDFa74eTYybzEmBgGQjOUH7e4L/GgWvqUaJL9ZbvVvEVE85tX
krrPojjXl531EiYHWIWyln8ixC7aL3JwxHU6wQZcmFztB4gFMvVqUb8kkS6I/u+xJQTx8ogEoqqm
Vzp+1Ux335MgMvqgnVNPxW/j8Xv2IFA0PfFq1NazFo95nQ+Hhy3rXGCLWIRiAVKjzwe5UIx/YKVb
zXJhOd7n9AeXhe4Gso+MbDWxCagHitKA/WYeTTXxRSDY09gR3EF4hgbs79MZwbcERpQLBt1vrNz7
Ub2YGep//BB0OP7AvE9yFzzSqtlurTMLjJcio3ierXtfSNfaUGV0z57q4X17N22dJyHdOtTxQdcd
lj06Ss9GzPPiKvSR8hvWf0iUFqCxy+Ayy1qFGlZvd5jPIgvZCbrOeht142TsI87WYFJ8y4MeqVeh
IUrjzv2ATEGk/ZyLjqVRvtOB4K0AOVMXcT1c0TnRFr1zx74LT9cK6OTcgV1PpG7/47D37CXVq0ct
8JhZvT0S5hQIP3obO6dKR/Do/MqXi+/d6EIZhGXFYFdJ+Qd89NwXxsYfMmemVLS85vMAAp2HNNx/
hgsHnbFr183uOFWHxQ81Z0JrkcgOm57Wwzt2rrTSydFdYSbozLUNCcSGEmHTgYfg0il0LqhzQRnJ
PU68ORztHeZ62PnKLgY9k+RsSJMxhOTQKH2LCxmBZK2eWeh/f0IIngIENv3glz2b9n5oyqongKX7
h4KbTp0pNtnbcaYAPubXWqPXTHEdVVhayOaf4Ym6Lk8rWw1qGyXGP1EqS6bY/Pd0UJ7HZaiBnkxn
sFDFyRToVdamJhU2NX9Y5785T6CpxL5MhTe5pjO6qx3pUlyESxAytTLxei/KiAOYrQ84FRXK9GTV
j0Fhxfve3sZ60Oj/kPl6ytrWHC70lsAEcJPhBpZbpPN9Im9HfOUhoFbmWvy48y0/kPYNgesqp/jg
6BQIa2BMutaDpruONI+X2tdjQ/c3+JbQpBO/OicjPDebwZ9ielqh9YnoS5t425BQeSwt+W22qO38
Kp6R2xhAyEPyAIikLIBQk2sLlqLsUaAXDbbFEejlA14ePicji9NqfyymMj4NjQkttl1Y4Ba8B/1J
AUXFNtAzRtif01VY/MuGEtaAUIaYmKsv8Y5xBmh1abtdieAk1ge3Ww7bDnPxwTIDDoE26XKDHhCO
7I8nfHJsW4051Whm/0MWBGrBdD1cBZUvSNjV0qxPA/Ss3gJ5FGTH4G4DjrAHkWvEjOpWnM3fgftR
qFiRCcQHx9GA76PsDMkySsmLzceqkyV8PxRX5d35frgXhU19sfE8uoYVYLb3PpqyIIVc41+utXr8
wUpu61kOC9NOniNl2GhqDopVAvXSqdn6wu/Oq6P/Cisz7ayy2N+qF0D/NsTR1B/BYuWzsCplp8Nb
i7SImj20VFlBWzh7fNHwhDU8RxG+e2PFfYsRtb8j8xNY1PY3MyhRtqmmQD3wT61cmXwA4ZfnqoQT
BgH7+nfsFv1SjsXwsPpXeocVLGq2sxICq5xCybxNmfPxeyRVmi/M05zdXfYh8EWUYD5E61IMTkRI
0CxB+8goapqPJebhJUtdUtyzg1ykHoSiFj5CBY+1+o0/2tGOX3KFxiOwnlzFIs2Ebvxf1PjGJIg1
PsXEAqwokmgM4NFdKbnArFl8DOOlvNWKt8Dj8+ULB2DnkUhun+1IqLoEKtowJA3p7dI8etgCX6/K
IzvhYH4VMAp7epJX+vmj5EjikJ8/VzxDLR7gqDwokDjqaLU4VocW2119nddIt7GjhBaTFxgnA6w2
zqiBU1suu5WdhsIbRzhLTJN6dSy+qbiBs+0cAnrFNeWPrY7h5B5um0mOVJUByMfAhYhxXnqvuw4Q
7SszNrWGTEBinYXub0MLqgw63jpl5XCC0XTzmkb07V8OwSkGeyqgGC4MMIoGk7aHNin+nphWIjRh
AockZn2RGRWr+rhF/67hxcRuh9qqlc4ZlzjlqA5dR7SWX/+9Wfy5BSgT8PB+80mrW3QrHd+n5XMZ
CcbBZZXehvUwlrAY30tb/3nfzslQtl2amle1/IcZC6T33odTN26f6LZeGAgEE9yTVM25RWvcxV0e
RG3ci6jzq5WV0ih8f/5dCsXoMNfXPp6qVKkDjtqnD5m3DwiBTDdEal6/zPEF+e+iZocJrXG4YOTa
AP0p9DKtAzJQm/uDgt2UOz4G8kb8bcXCy6mLvoauaa6bZB0H1oRdQ/YUVxo1TvlsFK9xH6BFVx4F
Pr0EFivpQLLUu+Y9q0C+RPFvzZmWtQ+y/QNCz7RmJ6dhTsqBUg4LL+UlLul8oSIQtMkEKvj1W0tO
DTTrJV55X9K+1b+t2hlVO5+UqwEb/FsUyeZMLa3XTx52O3jz06LlCBTVbNReZnGTM3iy0qr/S4mf
hgvnJGJTmgvpUVz1aanEs1g7NahrxOu4b9Z+QSlVe+79jPqikuw8IeDmduhrmmYxDULp7ten67Hk
zBgoHJpNhcUhjeTnjVPo/rdgh5I4D6i4EhkSGYa040LTQ42pvrekI1CIe4cwz/czIuAOokfHtVXq
op6Uut41htdT3ZSMJNCk5LKcotuJGtnq0vPuA6P6GGtxUgXtQnfRFDTexY9jaf0BRHWCwUVzfaAg
F+eA8ficCvE5zETAVs5kD+JJU+IPYIlc15sr6+L0Wyl3JFqNTPsjAIlQFW2OrquwEHf8O253sUgv
pTuFoWvCj8RdXKTXBKutbCzjBPzqGzpEmy3voS1btwzVejFY8ZeYLNx8N0Z4CM4FSVrd0r5U2fKb
ZFWmNEP1+iO47K8HwxckpnHiXUYziCp3TD6uUBq0HQ3Ui57HoboYMCalz2paG3GIhdMkiL4s9Jnr
DeGSC/ZOCWz2ARrpZJEKgwEzwViq2DoX66I04t5GFyKZ6IiLOhRAqAdiY6yXNFaRCAf2UAONR+Bf
nUz/+0seeUVswWLNkRPeomK4saLfk2O9jpdc01leB8W0S1TaOnHIb6gpaZ/KY2+KWiBLQYM/bsdi
rqkz0yS1BGKdzcmae895QVRtN1SDIP652e8YFw8yWQN5ImbFO30Mr9n6JubVmyxT3afvMfJrShq/
joYW+qZ4t5XvSu5sSH1iHRtlm3k2Dczb+HaJpFdELb6slO+TfAZVi1oKXXetE2J+0vcV2v2d3cja
xx8Re8GKmsyrjWCBSFbOUqqNJlI7FZGx02gLpCBwpy3B0ffASeFcBnoc1fU+qwI76pQFQifd+d6B
CaOYb8qXLuZ23zd+eJANjVYztqfHE/Dlyaj8OAGY5Jj00YJAAkyRtLibn6IvaTmFG2Th/ItxBmBe
G29LU4oCqF6bDrdXt1JKxEt4s1SuZCIjEcvRx3j2NgPv9/dcwH88pSieBGDjTGqab9ogDMirkwsu
uHMl7BewpLCenXp1J1Svpd1lnE84EW71sSk7IgiSYsPVJnHI3DdIfDboikcMOllQquVcT5Grgrt1
AVMZtLCutj+AXSCuEL6RGJza3zcCXASiVpLaGZpdZa+IBALBUTt8Vwm+3JboAXgPE+WWxWR1LUmZ
vP7CCU3DRV+9OupDYiEaQsSpbkiKcnBYDJWLnQVy6kNBZQfRzad9QYXB1nOuQ13jT9dXiQSlYuOR
p8xmJ2mBZ925XCQLFbGXiUhKVtFVIcU/+nx/1/T7X+tNxCxoHEnA3Yb+Jl1jyyiY5C6sVr8C0s/Q
6VlSwIKs2SjB2hFZYlsNLySH2aujELSZCXJwv6CAHbaLWT9R8T6noQIv6kXsZARx2y3iqdU+U+Df
AkejahqL93tS0W882a07NMwGkwg3XfU1B9pyTDR7PMOjmVRwvcs+Oqmi7LwVWDqvgQva3YLUmjFG
jakrM2sm6yUC99MiT9XCMLo7nyKXw3sPs6O6I9fPSyG7LKBRdSZavBmyHHiasIHq2V0mXk7DKWRm
50/CbfmHmFt5r7gxGpUD+hV/hR35SkHsFIDnAg04MA6uK5nIyKIZMaHh987mvXLjhTtf/d0o/Ie3
WeoyMbxb9cnm4LZzvw3plN3rzUoXGq/qZyQ1oyLqd05R2UHni+FsGY85l0C1DFPftogF0+VZj3f4
MPfJZro7ijcVbLBnjgaVNzURXJ+wTtacIAlREZN5gF3tuHKItwTBnvSenCldAzVRghfK6sCT7UKw
SXlqMBvaTqA7gk8QZ/1m0S0JarV/A+/o+3hRvf7Ntxow+1R9tVquxKXoFf9Vf1NI3N9GCR9spjcr
IgT7Cx+X0mD9KKguCMI9eFx/ilFZol87ygcaHElI/5m+LhXAAocKlXJPK5zYQjBFEK1DdWSDnb7x
iHGF5VlzU7JCjVHLdkMHJhAk5YKFTqzaQsUSHmEv9XeegPqZsJTXcM26K1lHoZAfA9Xcs3KWq7sJ
X3SWCOwvhixjXSq336KorMz51ZSarZBFnG/+lrJ6sf8lYLElEDdoJFF0gRaxzOD4+UCCilcQWVAX
zM1Ybp4V/uY08ORYNd5tkF15J8jIRWaLANnXfy9tQpeWmL+7l85qi/HKL3UOoSx+qZ6jUCfX28g0
31wXu5Lwo3RR5g+VdEfhVmevR5iCECMgM/FeRxEwPVoDbSy6S0MA5OsWoULGx9YwKOVlllLIYGQd
qQgNCFo+8zZ4xrgcM+A46+MnqiRr0ePA0OX4SEzQORmL1Knz0CrsDEsrJ45cwEyrJAkkhz9PwiE2
Q3kqKPYrbuttfCoKG0eKlKgmx1T0/kzp1mHIjUDqLvz8yD+wG6E9eRtCPLeMCaullci7FPjX8Jbk
sIZvMa3mzj9Xl5k2v3tk/zRa4Nv8e6v8TAUxUuwl1dm2FquaRzwZ1AB5K/C/qpm0fsICnyJtLMYW
dyywEfAfiOz80pZZiPYmQqhUH79Aknkkep979icxyq9G8xMx2VMm/E9W2uYZ/VGZr9+tibrW1o1z
ZKgQvodGUhfNmB5cmt0BeLLKJeNtkejLNHlU20MlzICyyyDcXyFwSECiAqxvVUK95JX57sDLAClv
VKO7aW2ReUojihtvkJT3Y2f8o8QFtBlmU6802J5LfSkAD94Kmhih6VD49mlfgGHb0gbWM4RuqZdU
pdJexizres59Y4hJUkbQ5ImIP37Lq3pYv5pgsJKL3bOADkMs2ohL/XYEHSkYLjg+f0JY1HHrZNLA
m9fJJhpWEM4W/SLuEGfq9EDiR6kESSiP3j4cD+pfpZqaTEtUv/gcgLopiRLX5aEjwGb60gxsmIX7
/AiUFWIJ1CGQcJUI5vs7FHgDNpky6JQbW/FH8Jk0bqoW7j4tx5fBxEuHDD3/oK6s0xxO+4GFT2xY
I3Ci3XsXBPaRVThNWbelRzrp/nUfZtkAEh7mqgLwCShDqxlY+g+d8g4fHQR4em273Aka4DbEYf1+
E0yfS+DTlTDhnfAuiDi/FhyHCwe+73MDkjsHulkZYgTLggdMQ9kWS0WLl8I/35IZZI01HE7GfX98
zPiR2EgNxUSNa5lZHSd9SqDDDuFLCzJdayYY8d37Lq0kk+PJHAZty9U4/flWCQHVUdD7s0mgQ+Vy
0MuMGJNnnfDvGTPhb6VSXuZXBefUR1Vfc48r9k0Co2i9y2g9CB+xO85mJ7ZLuJGD5gop1Qf7Asf1
YUllv5of5iu6Xokaxo0mirlX89GW3SDvCCzo5Iql/SHztOwnR9himhz9f9ju2ZXieeKS3v/pO0SW
RpTD3P8N9TtY26pVZI6/eOTfCsK0k3To5VtuNKrIto7cZy9tRsnFPylcXGxu8KmIKGJrKYKq25GL
QzXhn8uQTJvXCVKRT5OfsEZYSMjJaePZIU9PM/XYYWdtmfN9wVYA0RtRQxKIuN1yekSvn3PTzOIK
PEeJvcnfMk0FHeBJ4/DDm8P5u7kV5idsOC8Yon1dZq/Au/25kB46jGSBnE8YmaECJVz2M9wSf25X
n+xjLn3vs7baiSG38KFIFccix+kXXXvVbo6p4eMvrijvRE5GI0XgyE0Be3OHKHjmg5+JBFxxYLeK
0XOX3LPRVEUT51BQ+7ZIfrEZ6H3EHlzGqWp7s7i32JxlD5tm/3OD81pR+C3EsQruQlaaKkdrGAYJ
yjcZfz5DueHYfHjAW5bakwAcOFPo6RnETeHYrpXmIFJU3QCyWazozpK8FJu6fyBBP8q+4AMHYcFz
IgSWxmL+55878rSMqDFev4eNIjjITlcs22ENwz31F6jsbENV8oUPATUMW6zRrZBv1U3cYKklfiAP
Fo6B0/JClgArUeiaC69osxzE2VcTljRmmbXIb6uqcc8o3HkwhOeOPk8pmwCw+/LOpovFqWABexBT
VuW+K3MijJNjisQcS0idMIEg57rkZlitWVwA1uRnOUKtedlYu1Lb8L+7qkdSiCre40aMo3EAZc9t
dZjJcpXVLw3hmU8drk3zZfduukEES8S3qEmH25V3mRTblwzNx0iaGhBbAo8atx28xdpVpWpCb5QZ
Mg0gQif3Pp6M2E3LUNs38IgNgfbF+0UQEiVXj4RG/IS6lhVGl8CwSwog4aNOXgjlFrv5YBXKdpST
5aU/YRE7uHnpXXzneMw6ZxqjCcCRQrJAjNACpk+OiGQZzC8l5bnAQMwse8oQzHCQGhmDVTn82NxM
IMA+eVjo9kwJFOLoj5OQqRaY46dr4SrpCh+jxDzMX/SGi6G1U4h3DU72TZTyuaHrIfiwWCJ9FYYu
kcQVeqaSyWe3WsLPuj8MAx8PzZj1fPo8cCh2LAbmzZ6nWT0zFsBmG70BBOLdb7+anz7akpkitB/S
MscAl+sfp/DqPwVZGRk7UdwmGceFMM5TlUqdP5gJCx2NnkB7AYMPTZJYOimSmcg+hy6krqjusWdv
43tjYtoG/ih+s05l/VBfZf2nORrxn0M3g761bHl9gj+EZV8xRbbNAyJ2fDFdxApP05R+RaXPOnzx
TUmGLZqTCIj+n1S39f9j2il5haUtNBtAqVsbyBMugFPahqMPCBMf7cDS6penMxP4/tVvxaQ/SjlK
fVHpGFtJjxH79BvN0hUf5bk3x4n9VzNhtkj09JMTjX+2NzzC6dnFmmZI7ob5CbF40eMMiSEXz0Rk
EGHBsm442NFT3qUPmvH6A9l3oZnFMsfdpgxEy0a0ZcybSV6ux0Pb4AJ8uG/nMwJ4OWfxpMlAn3cI
42FXyL1RVf3FT4DsKN1JhnJvL3sxXCLjycICNE8Mt0yTs0IKEAe0mAEzZBPVRaOVLkDbNyuP0ZOV
6al/5bRzNk6KthuZj9lVrrGfEPmzuhY51uOc3vjAj1a5nDdXZzmZ/36wShgPW+CHetjU1gFEyzgZ
oV7Fncrx58vKl0SY4CN8sajrpuuDjQqUNIvRmUIwJ/5mllPO0YNprBuHsbBQKm8PfnfHCU81IkIk
+7skzpOQjILOBhKZEj85pRNibsbXGEbl0mrUVKqU+xAt5ODUSerwLfxbQ2Ouw1QbJaYGmAnyAt2v
wYMsK+r/A81BgJqiAXox3DCYe/MTLMc25DfWedEGf4sVicruYbpRoLFFFa/HWcbfg57xAc4/reQk
/VQ6CxidXIIdNZqzxw/UgLz53qTRYUvRJsKrUWtBHJuw1V22LZrED8WEHO3XjzapeFE/UOmzeesJ
jtkEVTx9LDlWd1oq4Tz+Rl7IUxFaa5QRl2T7dFq0alZz7rRKKFNftIdI6any8JSUR91lyxzbvnge
CDiPDR3XyhXw/AKK8CbbSSGnO+8L35nTIz8Jmd44lXp327yL/PPZIkWordrkvDiNQ0iiP13XJjCJ
D0LHGG//4TWoMRsDfrRq75Mh/9VwFqLvCsDYaZ9Ptm6iXdfUOhzrTvKyjXwZAa2LSo3noggomZmP
p1l7Aye8rQl72BK0iLliKITkt9oMWLoJht50IZcWg8n2F6t/Tav5zctaA660mSD2vL0ZEswbqrmS
rjoOnjH8v47yjTN5iPtXXwL+H/DMSsUF7uzyft7S+uxnXlEOsbMH+SLKW9ghpzJjIw2Zn/cDXWXg
uS3608WUDwom+Q0TOdgutlJtiYACbmH8t5pagX491S1hANxeLhrA5clhoa//ZCLBnvkUtY8kO/Gg
JpRhq+FJgjVvP9zO7FyS3wIseEeIFQfyOi4wc5AJM/qsjWTCADXTg+BQG/oEx6GBguM5EFchAExt
T4xap/UkeRAaU6pwow97XhC4XWsPnaZ4kqApjG7rkJ5jg9x0Zqi5o0IiaepK5/srQniJYWEfBYfs
6+dGVCgkwVW+yTf1Am+KJ1/ZpZPnouyfhZOb0JX736asIpEiyGXpMVzb4C/lN0JaLQeorQDZF0Nj
38H8com/pjjvupZY40Ci+wCaYvulnZQxzIt0X5aYgn4cziUOOuGc7qaTUwQdSEL6Afjyc+gavrbE
hBuN8ItTW2RrTtKrx+T2nFbX1Sxui3VNtkPA26QuOzFBfE21IEbgBx0+76fDa0tdWQDD/Z9o5qDm
VSb8Ul6dCOThzR4FKczVf02Nt3ovMbuye/YncMLbL6Jp/IldRNta0bxFDm1T4yUYI1hUpigCegAK
V1a+sFaKnK7wiTNQenWj7WKO/Bcwa6CUAuj7L7QdJvm9rGcVjl6y9C0iyykbPgBeZvbSWI4O4HSE
2RMIWKmQRjqzqkz1khE0LkeTMCPffw5xLnDfNcAPRwT1osDFCBP8hn5Wsjq0PzVUzw0cBrt7myDW
w3aPHofRVUDilswrlHEFh99O7bS4SxJ+wf4uIH5Ybd9t/Q10819+26oCy0OxoMwluabtV4OvXk8W
ewlE3p0tf7YD8nFqB1puKyfM9geb+6CapG6TeAh6C+SKWmxb6dghLPu8ynJZv471f8Fw/t0VppJ1
opfMpMH1CpsPCMevNF7yy0iXGnyhubT0ubb5cunzLkNwrYa4uZfgzm/uKV6BYqD560zfoJZ3Fl9v
THz3WV4TLpgaRTl8R4D+5zzcAkx0IJJqx7AqvQ56Snn3fx9T/7f1m9285GU+snZ/QAUE0LurNjFG
2IVb+7RPSeaOkydiLB6tJ1eTMZl7UifWlpiMIkIe4RnMWIKL7t3uzXdebgEBK2yaHgYjkFW/K90Z
DKKgs+u/NaDBnKA15C6tHdeP2f4QyYHBjB9VF65cZ2cXOvr2uR2pLQtIIeRPPrv/VZgCyxH11QG3
NMMyob19snbMp7kQl4uhXPrB0kPPe39QUU3IsVVNsV0vOCfdl4sostTlPbyryZMLZKd6P/dqVXA6
pixYAOjBD1LXOnRhEGqFKYxQZ9PsRaIaAODKn55r4e1wp0Do6DUy6L2K/cfebCxVLPtyDOJn9bLG
rdeg8ZVrEvpuKDU+cAYV2CGND65flMAz25VTD0L7R1fTA6gkt1Fa0cD010QxDxAFBvAu5WDxJoqv
nBrbVWFQJR4VFMqQSil4EJRCTDXU8u3fPmePMfAa6Su+fx+kyGrZ5ETr5XG2gXmyncA4cV+Qu3qf
wKxlJjT06T5sDD+5cNa1JMKibDr12MD6b7YA895zVEGMxzOYxC0z51a73DLq+492sb7UznkrIc22
GXX66D4k1LkOgmJNKHTF/bDUCQBxs9VRoUdkJCOEAePS9JQHWm6PynatRd+5DSZk7ADHvjnYGwUf
QGJu4bFXdu0oEH+jLgw3kjo79ni5+3LmeJ4csDjy1KeSANWPwQZQtKZzWy0mYqhJF2JzXODJwJ4a
zCQZ9cenv9rCFXw+iUiimMgd5Z33cGtK5FGAn4rACHxvrbQq2p+niySAzbtPInWolYvXkXwxLwr9
TovxuLWvswWN14Hkq5aN7h686NcpmsIw6egx+zRVvHcWz+9gbqQSbhc/ujvjCly/krDPb4I9iR51
WX6ZynlUNF3UdZ90Zl9ytbxlbjsA/0cnh2eT1g5q9IOK7sDU49hWzVEf9kzasLZaGfN3Yo8el+L8
WNLoCVkdjKLfqgYdxworwVHspOs5mOH6/sE6tEvqaM9dyg1KJvPSjApQ+0EQke5nshKFMCYJj2+N
b2oyqNL4RKQKr/KNfZesObZOtrRCiDMdCpiG3QgTJVmsrqBpSNV1d8Ukxi7J0iFYkZ25uOQ6U66D
8bbKyLpbt4VsdO8DgJpm1GiwjzsGGFB11jnOkf+b0HMcBZwq7Db32ISDvghYnzwi+jHyKuQtdnxl
UpcR9T8pcTAY9uJhV7MEsDcxj+sN/20/NBSNUYbLAC3an0ij2BhrTnADdulIut5M+u2BytFlrQ/+
VSO55ngy1aGwLaRb1GbYZybX0Aley9YXjRhajfIQ4ehGl9ZJ/tIoMyCZLjtWpArjIVPQyHoDGnLc
zlScWG+lXwSg6mKdFse6QYlYYA6HPlnnN5zsfvmXL+xQYuRlc0wfBT7uxvQzh3iHXhwvVZbK6YeL
J6e955o+Fq+Ukbnf05r/+k6cy9/lv/nJ/jl5M/OlJ/3sdZ4e+ba6g44f1/aH0f0ctvuoM/s3ik3A
G3VTQ705tb0y90NRLmOBeV0gg6+IAGm3EQT+TphlCogvl9byTDbAslqWGgH/uD7C5iBZsy/LsHzx
Z3RWGNDry8d+2A/hKBS7kALuDJ+2K7fIg8W2h7V+wM1HzOYjj8i04N87/yhJrfx9ObeK7C3XNHQ4
Z1G3DaUJvhuVhxPVtmYzTLdZIeErVoQ1Py46gLadq7GjOOnJ4E2R8msKOukeceMcJLyrZAPfeEym
C1CXUV/l/3P6Evt0SGBVXx3uAzxcjhxugU+7Oh8VXwfwGbsdTce02WXH3LH1mgVmVJJa9/pbMQF8
6eums2qC1T3G8FDISwlmahkLtV8xh4ZZlCZsuH/Hb1hRDlA6iBtQZQbMOXoIYhoSy7dbe++1ApOu
DEqlX8kKSc/X6pKIN0U63ygt7/IUTnJCOgojle/3sBupO/2ZsmHLoWkuhapQS4noibDvS1xlL3Gc
ONWqrX7MgBsgZZOYCClNW1n+NuI1G9PO2A7PvvPSkOuLENQH5bTvrcjSw7DCmWNQxY2Q/lBfrRtv
rCIQu4bMuXnVbDV+qAqnN5lb+zbxbvcMrLY5ES5kpa0FKJj0d5aB1dmwfMoIXHgGZEcMpHbh6OoU
YJ+j/prrnzrnJPrbfgSOZOe5D7uopUPpYH3gqV137al2+JsnOMo2xaRbi4IOKa9A8vyjVQbZxiO3
Zh+Jd58OuZeYnvUHsYgOafS8XvK+0/32vGt2RAWIm1qV1julvAZKp1fRvo6NumgGTaWbNcKfRgQ5
p6B7jKd52Ok9n0/srgp9GveY3fOYOBaUui2cKjSpXqT2pE3iBaxPMnd3HU8XVaxUpHXhs2+8BfyS
MMhce1c301LYaydUBNGFKImbdt53k6kThSzidXeYOncd32lndwDTJG5dxPpLlPAhKxDYNsEOA3WR
rdDOMTTOM4fBFI8D5Z1gvfEsDpX69WRJ4VWgiq6Bwt7K9k/Bn+NTVBR6o/NPzxCAKDhLNKwU6v01
eYqr12geMQX+DgMv6EB3UNY8NQD3jt+rxlQRqOHo76BWwXJYyicVqvZ6an0Nfco371KeIz9eXZ2e
xeG4uWrs8KIrcK5Qta0YlGHcdjGTpd9THwxwFIVovKD40/lJfrKmefYkRBaYNMH2xX1NBCY+anAR
cUXDjOXl0lpRH+GXB8q4b4O4GLkCYXISBKkuaRqc1FruEc66CTf1rTljrFmcS/gomOz/+IW9GEwn
dqJ3Kcb1EBZTojj5oML4DYSgb0eBQguD0pFpd+wXNIaKaj8ph7UHcTeL0BHAaA2kF4hjWI06ygaG
ujARH7RvIkqiamWDaJQyiKAPCz0yKcTL9BzadaKa2eFIwp+fLjeAq8LYfdTXCsDYChNIf1K4WNLf
KUHdNVs62inT1MiHuHS8e4UWKg/HH6RVNE9nVhJfYLEBe3jpOKoRgnDiKjhWcrCJ/myQX99Nyuen
oXj8bSlbJgXA7Q8sFGiNqHe/r9PIvwdtBcnR5LqjZjuHvCF+s4+0UZyk5YuZ7E/is3rCSyHjTqab
852NIyNYDJ6SuIT+gliDwVvQkQjI6aSxX0UMYvfCwOA45pUnFbfYjnKwP9Akqrjd1Sh2LednmGBM
75ZGyHGXr/poizsrg8ACKRww15SQo209jMHrzPQJqeC8v6kMVMZ4YaN9/4GQVl0XEkB0Fq8iK4Np
ZqDy+2z1WhiLgIefJuUAqO3sNJP2H4AfaCnl/FCZ9/2Y6NIutIDH4nbeKv1MxiFLusgMZCQKDtxT
pPpmaj0n0REM4NE32Q7igSaCWz/5phhgIg3ZNTKxOZ8J1yp7PGrIa3cMJ3A3emowLDvEAg6jjkIs
99MDBfXLj5Rwxg+aykDMiRsHJ27bcyp4lYyNOcmAfV6KCB9yVusacmEzdp3fVtvWyB2dpi5Ncm43
xVuXvecSR1JogG511T4/OhuFq+GBdCaFOYFeM1OzpHTCzaiuifyGsCQ21uzacS33ItbyjdQsBqp/
PsUyirKLKGq25IzvZKHsCMN8Et5dj3miGuJ+KxGaW4IeMaqEQyrGaltX8ngfbCuuJR24OfDCJuGt
xbz9+6ibWfqK2RY+C9nX5/VlZZqkjmz5Dx9RJPw+KpV5b/fY30/wx9rhBVwihFNvfMcrp1q1VU9l
NZLRHdvNSqsjPU9lzivLDJciUeBOUvBkcdVIu3IRg9nu2t9Gfcobka/KhCK8L896k8obIGuMcBto
7xJ+rfvUrZqsH4eyqmGHmwco4ms5bhsF2oHNoz55UahH8tuoOWxvqd9SHwPhn1e3/bTd7RFLRr9N
57u3GJA1v2gr/ulZgPmfNolT/PdZOeQ6fbL3Cdhz3bPxD/IAhPpIVGhUrHR+tRV2Zvvb+DIjElCn
6trgoQojyeqT6bGt9/OzQhLvtixErTHI1Ijtm7kHaIqucs7cGTWwJiJAd4bhnhFYtcVf7g6EiL0Y
PT/XtnF6NFPqPFEOpdGm4/SV3OJ3Gt+H9BYJloRmnJ37eqvOIKnFlxnJAEkDyqnL9obc/PaqmwZd
fFHR4FNKXbdPWVFwJb7LxR8kNhqweE2E212KmAK0g18XHsbv2khHMltT/QuMAIh/epltNyul2FVi
cUVMYznt3dwu0Us3acnY5HdZsAkOqh++SZmHgvYOhiqG5lm0TRv1XAVrRAc1r+FnCdzlCOMhLUWH
5g6Np9fJbd1O2srIn61aw3L/J1pQBG/Utto4IM2mU9n2niRGaK78BSoWnOw+hkv1p0mG7bDVqfQ3
jkHPwYxAjl8LgTT9zP5FgMBv8tpJfuhNsdUBXHhtPV8u3OmNmc8RQOLLU/k2D0970sO0K3/aBvmq
/MiRkntOK30UnAS3GIa18HfSaj39d5w6/c5fmt+sBLDOgLjoCfNWyvg7x1h1Opj43A02pdIHAWWw
dcteC5zMrhqvAk50nJ39n3iA/tnQylZ4hNLCVwyET62FwVi2Yxkt6zq7EyXAAXmqvkvjTRz1z7XN
K5YKCcvVCMAhAvDCg2/j3BVXiifI5ALlao6MnqpWOY9sIPrVaPrsJzHAyrnN8nRn+s4GNMEFlRtN
lD2JufltwyackT9Z562cetzLfxLdZI0vC2O9ymhFYoO2eDnbUJ/MwOzY5cSPvB6hlFprxx31mynV
IyLF+Ic8D2Oe2ipCqndcoMMtsrpNzFYWZaRy0MuRdj0WplWuYbAM6yfBD6RUhqJcVFHj7mWzqPuf
g7X9n3ljvj+jRy7NeWRNfuG9bfL8P8Vmq6zZ/eMTP541YuEywo4x5kBGSEkt1jMfM2GWw2PaXrlE
FK2XwpWP6AH07dlpCo580t/gVxz8jvDZ2zUyqe9wyyLCWN8HhjC9J2DTzP4dawhV2HxuTy0AaBVF
4yBhn1APGmGvfI6K3U6VSDyeQy+i/TMeiC1rMV7w7L+267DeEhodKsCNLJXbvfut/h/c+2y8JC/7
Jz3kQuF6uiyNMi5MAFsQUK+XgDr0SAKJaNm0barU5Wgsi9jdQ//eejSHAaRc6656o272TxWghhcj
p4Ng2w9xY26z9k8f4V8AlKGEDoj+/36/G5mGHgcZS5/SZbzU1B9dFBSREkuCV9Hr4u+vhTXpDXBm
D/jqZ9Hwfi9uwj+GNu5sVSAsiIQwgYttRy5cejkzSV1+EiABTowDbcMeVUpFUPBqhYaS4ayr6Nse
VgzmrBMCpcKKF8/qwQ9SIKZqdqzmhJ0TfjoRTIkrYlnEJNCVMwvQ1TtJNwhE7votk5RHVGrlM5pp
GxOM3pHfdeNv1BFz8gvBVh8SZJtZjGLdT/r4LuD39eFklnuF2wMPtscx5zizA8lhotmKOvUQPsx7
fTMXnTXU7IpscIBXf5qUSdjNlxMthVHAQRfXEa4iv5X0XaknxYBvO4peMAE94EpQGZnLnmSsTU2d
NV7ouD1CVNlXj/pyrB2hgq6Osq34RrxG6f3HFTQJgtRvKQk+j6BKLvV0cI6+F/h2duIVIj0sHdU1
3ZVJvhVXkTArZ4HycHbQLPRtHoevg/uhFC6SXorP0X5WthU6Fn+9SOiVK/xcd3nrNx5+DuNBubzc
30h1xVbDM4D9utBFbG40uASqENxP7R71nCTH/YRUSF0rLAYYaBAVmNWPwIQNEIh8zqUztN2NZOhH
naZ8pIybOO6f0Bfdpo1DE17o5V7Qu/jx2CqKjBYOoK17wI508hZquBh8GFwDqg8kZ27LLUz1AySw
Uuqo1+J0kzHTPRdMLN8jxwKigbJXiyROz+EK7E3upsN36vHXJswWTpweN7E/kpFLLtnBMKR8uMUy
nZmGc0yjmwp7EN1Hgxrt7ruYYkRW4fsqzdMKGS7d3wLNMVbM/P9vX7QRDMAtuxgYQ74Ozs9WlV6Z
v8deBD9CXb6TNOXWJ1mdnlgSDP6ShJZzgEZuzmwj/tyOWnXKNWFUh3LE4R0HETnD7i798OA/FY4Z
BFCIS8e23hmJm1JK8umiX12T3JTUWEaqcRdqAKoyOudDh7wgZ4Nf7kq0jav8MizlxlKa4g2T68IB
kPHUjfAGJr7Ne+ABD1/0qJk2EyBu7mPbzUGWE7GP4DZzRlPYHOlaY1F0Peprgv5LiulqhOm4DozR
+PJWSAhf+wjfOj7Px710FUOJYqBzScRpX2eUfQGNxJ5/eguqtxfoM4w0AakcOOEPDBoaGdj2y/li
V5e9MKtSE+j7wysU0dj2UXBdb+/S1nHlo7DmnSFNHQTfuB79FgSPwWDNwrTJoOEwFUnRNAeF++Ve
EmzqcrpJIl8y+paPzQAKY3GZiSAvqNAFwiU2raW8D7HuFuLOJsfi3BRqSsD8dcoQ2Mffp/pn+2Yi
YH+TNYmmrUKZ7r5SCyhEsE53jWXdFA+xBOranb5nZeRqpwkDuSyZ+PQ+ALOr5tJI+mfx1Enboydr
EuO1vR9j/7WmbuK7ReDxTs43FOyjl6f/R1qULR7XnPcwZDcr66Yl1EW61o3ToPnJDT0UYGk2s+OV
xL4gcXgDa8uLTtzo/ZfjcckZgsJm8//VgapEOrmMufHg+LpzTn9si4EHvSlGcpSSr7jPF/bSlTeN
gNyhCuMq3Q+xBIL3xOiEc7YFlz4xFBsLFY4Od2Ek7gspGoaXbXufyZpZc3qwBihThzqOEWB20dIA
xh1YE/ivJXcOKkOEiRKNJR0rxWgv1bcOYbdbVMfimST2d5fZRFyPQIKlhbhRLXfby+w8gEaRx/Ej
fTQujzf2spwt36XNTTCUp1G6q3Dr6k0AwmIIAOlELEa9n2FI/OCfR8HT76F8OO9XNv6dJ306aEiH
Xge4CLVeuPVou0GqcDHQyo+JrRYHtm79exVHwTK1HBXjwfV7bGxDKqrGbFbhbVAt1Kqz8CR2DlRL
Ml5XcMkXo7NdCw2jTWOYVqD16MD0fA8Jt/HZpgnIp5Ic5cJTlIAdmoPhz9YpfsUfSaWAYDmWwy9x
UIWj0if+L8AIB1vGUO18bPGaNFt6+sg4kLVV/2Yzbz8/gqhH3W9jN6VX3jn3EuKuIaJq2tWF3Jpi
/+mGagvJJn/wuMKnOuGvSYrkVw716/zcTcEM1BtIaQljirgpc8ZMY8qcQnbOfRJLRtyO1KeHD1xo
kEw4BsEDXDAggHx27Nbq8UavEvk+/lVxQAdp1AggOw3doNjH9QVlU6qGj/bOlkLDrI2CHlhiyCud
UNomUGAeiGJH7F+rFwp9FnVhId1EHE1b2Y7zY4DOh+fmv8dG8tFjF2ES2PHUPzHFc/ph0QvouerQ
sD1NdDHn+2hTkDaNXL9KhAr0hqnHxnUPXShoPZ++69ZMhGNZ8nUI6gTtOLNzqKucvM8NBouKiN0h
0Ah0RrStLoN8U/zy1qoJzv+/k2YBcYF7ZdqDQVQqE+noBOskvAG96iGKGgjlSFyqThZ/rhMng7x6
RRqtiZWaJVWXeKNZ5xoycjlAySAQDexmpFh5cYxVklM52aubp/YW93C43UmuYsWhp7Fu1IH0Nbl3
8rfufSsPx7WAH2hQCnharBwtFHcguoLtpENwlKqnic9eVxxecOJ7SF8CYHnNfO9rO8BN8uSzZ+gF
41mkAO1Zn5wJ39YEBQzpV3KjjildIHBEDl+qN0TmAc3xZJk6fsEyE1sTOMy1zwppn8Y5nAkGDBnd
KDJLWP7APdTDLo9VideuAS4pJinGNveStjoyCjkBJUqgFL48+aAB7kY6mjsiMDOgRw0JDVZT/aHI
8jj68uGJz6+de/87rs/Ahxsnji+XEvIKVWtR4Dwie9X6ulzHsXHzIMf71CJoCtnOi58ndO7DGj4b
Woh2+ixO372bvrY/1VCsqqWVR/UjRzCrO44K5vz8BAyuj1RrNx23kL2i+b6dK2Go8RwFw/KUITun
WuUmI0fS9tx1G+4INfe9JtdI1H3J9F948lGnHDELLO3M0Q4VqkB8grIHJRcPrpkIZjnF+VbjaWnh
YmchCYkWRsd+eQN/4JZq4cWMJ3mM3Z24tQEWs4AAtBX/DtqG2ZfgLQCXAAdT116zUdojsteQg3Rd
s0vmZoEG7rcEPYtMSzxytxdQOYqaXrBDPih2XR2M8nnEtuj+LU7lScEpcsEKeqB+eSrqmnfYKC5j
r/eSQCWYcq3Igpj/5uniJ9MRSgI3VxI3J9/Qnf/PCln+b9uA52xLkKIfqplIY26uOEnKpeuFSstA
5OzIpfUNk+ypSbuk6HMutZdLtgWznKfjPpk7EYq26PSewtqtgBNJ0WCRhb4oF8p1dj3IF3U+nwsF
XOA3TY3GgaMEDQSUjOyphTzWQM9zezoD813dqs4U5XBtoVd9mIb8A87+Som39Zf0wZc5JB6YZXNo
JcN4wpsLk91Nn1u5RLZcGn3mxAtq636q6EPXsHF6wZWK8zRM1MA8XXbkzkGDtnksmveYoMIi1Rjh
VWStwFfkOCqf/b8iPzJSIc11ytBkSYe4vnG2sHnphGguSkjMkEevJdR+GJZ/MWDyhiZ0Qx7CAaFA
G/PCzVRl+ZcQ9mFr8jugSB6i1H4nQo56emViLjcjR+IC/08hWdTZuZmRpeYcoTWDuQeIP6Vll2El
ywu7SFZFxCzBBbV+ft/apeurqvijUluYy+S5ZFC5foeo/IMTsYYwcXYT04pBo9AtHfeaxFo+1pZe
HezC0ucJD0ucCkmjpis7eehZ6PsN7lXkJJV2cnfg7jqHotlMBRAXfXLYJP4k+TJvPqTei75Iwb4L
+jhQ1mBlxgOoKOIC4q9jkOWElaC9Gj2IiP9s0ebqP5e9dHCxy5/WKNIL0HJX7RUD7DtveBguYo+u
+2s2j+yXNxr33uJzxx9hAfVTirtAcGqGy0cYEA6aIeLh3P80NRf3Gdb7E6Edt6TKks1TFdgHzy1m
TEAL4iIYRAgC+98lJDL61Gf7lYn8pIPvne9OPvqZ+bblbx/bZsuNfX58tt2d50Ed4tsy/t4bEkCE
xzJL5Z+xD01fjrcHswRG5V35N+4Sb1GNgtRr6TpuPzaDWME9bowWuv+SX8llOvunAZ2dTXAVxSlb
hhGwYsE8Qjm6XvyD4FUHxIpyDzujW4v5QKqqELxnie4mi3Yj5bm5hw7OCOnzMnRkVozq1BoTQVmJ
jkmfzkLnJ6w651LzC/lKDFLe/gndAdZq6RXrAJZlE2uqF/WDPJf6A1OQakH40hKpUtOWLES2O9t9
QDyFHqVZ+jJVIxDm5LgzeyqyuQL1ptkXIrQyiuoFF1raxnWfZhmhlsS0APuLjUg6PcMgedvy8BLu
GO26rGsOGhDY3EcvG2f4GsXaJMZjSHAXJGEzitu2azvwnPrKCSfnqywRviU2VXrPSX4zU5+Ox14M
tdOLWNhBxGzArXNn9HgF2zIz1v3CjOer2b5qimyBqDutJZNtIENcZqNlo7Ml9SiJ6O7HlGagWbwj
is9xdTNMwH2RTm4sq6YZo/HITKSLg9zJIwhtPAIsDUxKOV3WiPmm6ppsMGJJ78v2Erks93MN+DZj
bxEp36UGQYXSkMnvHUnL/SVWLs2oLTU+ABP5Pjwx2A5vhVxxIgAXt5cMF3yqVyXBaDpXud+gXw8g
nxTaMdFcjROVD2LHbYq/eL9shvQ+PnpdtaAEVASJ7ts+x9EKCrZKks2m6SV099SzBSbtckI31qUl
vNeNFNTHzc4lgr50eCXYZkzgq82S9zzkqqkwtYm/U3q3e3/58Nw9+UZbRM0Akk1DFKZPwdOI1b9n
4DSlmrOqG6CpBr/iSQRZ7EhtCVzDXG7jVonwwTrbxJ7M+qIifva1ay+axMPbSoeTqkKTHLUTFn64
cmOq1EEW5bt+6gPxx1lgTYUoyhdi/de5C4f992B8rpXwsekKx9pdKHMc8Hxt+nd2q44RhD9PzeT/
05R7q8ceN0LeM8WW/ld38Yi4Lk1RwwsIK/mkAk3sse+uHZ44VIUqlpSXy6Pz/TBygM8GEC/c80Lr
pme3BrCojc1kCYVs64Dp3AkiyeeZmq3h8OgT4UkbLQYmV8pzLxHFo+FHNnIhsNeEB+JuVOZXAlUJ
/SECE81p16dozuQ1z9smlBJ4NFDDFoE7wh7Q6fmYTmkDyf5j20nWt5z/EVqM12ib+emhoT/mZUiG
p8OngACwdfa6NZq9eM6/J968b7l3zb6jpchXKxzK8npa0NI/pzP0OiKCTXv3fwy/bbuT303bF43l
c9UYQGIRLhmT6OvHP+9rKRNHcO/jxksBBp4aeMF+m/E0agygkapsb/1XTSSWLwNK+zQSgXMcJwkd
SqUXr4QvhMZcsXx+5tigODl6rE5A2joT/jX/xw5EGz3sJ/TFX2w03UdWy+KYr3SzoRq5Ldz2TT/z
f/PTOysmDXnfXeRVIhJu1H7PS95UgyBdEiZ0UeffbjHEJCl3yyav3xvRf7rGUP2sZAWvAJcc3JJW
VZjYUmvFYqFNZ7v9+q6cB8w0jpvEr5ucptVe33jtOEt+mhhRxAToW9y/BFGITM+l7FnSdW49dbrt
wk7kGDZlbzgQbqz8Al7rKq6CaESiJAhlFaQxML1pXWD4O8fTXs6gpBrj/OssII2IIjTzB5EL59oz
1+mhshj1B2LtskiwsznZu8Rb+5Cv58XtLlMJIHqa8uZMqIJEUMZfQTXaV8uSAAkkeg8GUJvC2sh4
CTqYb8M0tbatyw9AjmKOmtyYrBd/IFH9ND0NiwjydIggUuQe91dEunsjCh/bhfgdk/Ta71/Z/tB/
3L7d0haVu3xwHNQSrOX1Kh2y/ahQ7Cl+LlyGvgMnSPmitc5Ut/+MQZ5Zf2UAbH4pZJJ6UNW7LL2r
XGlfHhrYdNoCfazYXCp77Sbc1N5YlsfzxCyMIg+IyWsjUJsMzPD/nYda7Z12R1wNvo8mMoZlieH/
40YzGMnYnR+DOkP2SZpDfxfSs3VedJfJk9zwIzts096LvVzN02aq3JsDh4TfOYpL9b6Bz/oixjb/
uNAxRGHs9EfEhlLfosM1q1YM6zBL1sP+vyGxHy7Gh9fzfPOdqPCIn7bo5TXfJbgIwJ6Ho0Er6136
azySgdKUrb/rZa51MyS33m781AK62vIgi7mfz6fz+z3PgKyVF929YAVZNJQjiBvl7CiqEschnWvx
qCe4vxv9BTpiLMnHyuacbY5gM51NRM+91k8OQ7c5uORlX2SBHq9S+ls6N4XFj6b7yzs3LI1XU2Ed
ZBGzikxDicW3uYb+CocKVUW7cMsbWa5Xj7iZlZSyb31dha2yCB5CI7FawfTKlgAt95DCSfEiEA2b
5lwR6flEZUK4X3OE7sUgnbpNTPjGUeKZ+wObZ/CKtFOJMIyfsllcBUNQSJvJgKdpfAc1wvbsxbgk
DhSyzUILfWhdCkVN7QFJ2gzcSnQwHr/qne04O3x4ETvJI5Lu7c83HVFktbgFPys5HUWlk4x+rxta
oLj+WhTGa0ympNan4vQqJX+h1OPAbXPdrndVdeqT+H0H4vC9qJK8FkgI6kKMdZNCLH1N73QUHGFy
B+rSGS2nENpMgeDQVROR6BK8AEYtLpzyuHtwTex0UkcCmYeJkAu1/VSXkfwTooafDugs1sY8qwYW
+KSOwmJoFW0oiLer6mStA5EP94g4Bz61RXyVjK8yhUG944oJ4hNiL2pBCn642zfP49bA8WoI6Att
49BzKv98Exrk5xkoUrIurY2E6Tv/EgKJGj3YAtIKpHybN+nOIaj+H3HAKWxIZLCKzVAm2Fu5z9kS
WjcWrKoke1/wDEk2JmipzfltV+X0s69ri0yxldNLYTHX/MCqYxQpv10ENEp5DQa6R0922wkbGzrh
Pu0bzdprk45oyew34Dk2s5W7mlyi3Nl9ONIOXs0yq6isPvWhSxTRbvaSUXDrcEh4rNatq5FpIdti
jet3WgqBYDZBcQ9ox/E/xDFDvWEc42BQf3vRibIrknHZ6QORAPtWDUkwHaV+ZvuFBna8XU/9sVIV
2//rgJKSfhHpj5gC/56Mf3HNCY68ObDp6AI6x/8GvAnbrOdQgYIhHEDVL1FMZXRYnJh9CDutcBsJ
LwE+ew/CctOq7JsAo1eDhvCB7U8KYfxmq8Oz18zbmTA+afVIx6dnuYITGmxmFTuDnZczGmKHQR3/
zF/r4NAgKDCaT4Ax5NexWMnitprVzooW1NXLoNzS8ajwjWR3E9c1eBO61ucwr+y214nv3rqIyfWV
GxzceBktWDTeQnww0jL2/uibh1/0iRUsF3llK6JDuVc9QuGT5QztBmJmWiRlp3pBxbnIQe+pdtCM
mbPHDUViAQR/u16IilZvy+3DM5W/1xyUK7WIJv8boHxx+r/ILd1+HbhJLFkV8BRx1fdfKvP//hQ8
Rf5v1iy47HHyeUnLBKVPkXM9H5DEQDujaK/t9ID/Pq6EWKFph9MgsyN20jcXZPOCrakZv5gdmfg6
UejTYIxL/knMAODkXvlKZmmGgosdWV6qXGmn45dnSnlPHMNTUHCE4tbcxDwKhflhr2lvQmbEQXl9
01SjJ96qLilIZ746VdzQaNSOblVvFxoEa4I/o0gLlN7TSFPyBLBShiNtnAkT3sRbAxAJb61Pc7/3
bswJlxDRng53EpDZcbSZakf7QtSdCVK3UJuqtPvNeF2IpPGYKJH8Z1vHOTzZkO4vAdpAMmwwe2Sy
iMG7iO4S/bMbH6Onc84dEj3pL9lnPe1p7ZqEZCXACYCKtBT2/ATVRt2m3WNOGHYM3vOsM0WXtnuG
CqYFh+b54ijBeTFuSdUkjniYplACCwHEqYgd2KDeUU6htpwPvFawSpT29I5ugqZIFmHcPUVBWk+7
NgfLdecXxDh6rii9TPnx8HSg37AGW++VQ5wt4wBLJznINUB7aL7o5TjGu2ZbEaVOl7DTJUE69zAo
V+YX9wyCgAWu0zJO2GKPSMFsh6EN2eo/0h3p75K8MRSCZ4GIYmHxGoQJkBkmLk1y6on9IohpUsPf
EqvSK3kw5yVA/4caGovjvEp5s3sXSGCl3ASf1ivNL7vM6RC5hMQrBdvgZwNMC62g/27QpkCRRDc9
VsqT85PnNf1MdUJ2ibQKDHP4SzXMwh71V1Pu3k6MkBRVWOtq1UKp7EQgdSRbsZp2pWz6Pybz0i8X
ZrAxJkIvnHS+u2jDD+4h+Y97gghBOU8xlvz9nLEXZg+yQvMKJVd/JCg4MGvyqJW/DMaIGm58RZ4l
6FkEbh2T1PjuKce+zKrMJveV0T7T9zB0wDV18BSp0/vouMR7/CaSpEvdLI37XEzH5CeqTcYjUORK
Bo2iwA667RY8SI2aiO8AlA1y5cthSUS2S+jN2cqe7gZmja7TkZnMosV/U7X+xjkhytF3xRzoDMuC
EpHEv/fAW0NqbO6zqxVl7dS5ny9GI1VHW0Yg2vC43edhBgXrFiJOIAiHFqA6EiZ9WE3NBKNQtNG+
XHztE21tFxGJaeQFIrSbOaZxhd7032MsTYQ61I/AxsyaZ+EDEdR+gFJjUjc/SrkFzBwNTy2zg6at
ZHYWY5GmmtzQZ6TX4jnbzPMxF8QC9Q+OhQFqLol1z1+qB5LwwUN10KKtd8BAttl8v77IavrUuvq2
N2BU3rReQY9jxR3M3VuE79gTFvynFhmfWigHK3hBtPNozqQrSeQew+a/lap7mCkWQ+mMZu3KadoH
aIwdSSuKG4D9XbUsOyNWHndkOrTSPKSjNlUBayS6b0rehPOFOGbUCqe2wOYTAuzYR78e8yvQIfHY
XvIetVLlETWU45FXsjJs7mZqxn3Is+FYop60r3jL1ml6sqKpHgxh7hBLmshlWjjoxcMIwXwNlgfD
oT4AsYDeikbF16BPL84LnNedbQoL4aENXwDSf6SF6q6Bve5pNuw4b1+Iga+y8FP/OFQrr1xaaWDf
Tf0LXgUi7Q7FNLvLyTZrJjtAbAOValdlmz/Bpgt28DZG1CXDJNpiFWEYmtiKezas7I/eD+DR2mZF
O+hmBCDJliPBG03CywffDAG+vSSg1yIAvL9XKYnY0acCGwM4Nf/C7zsTTZqySp5MaX73Fy5AJFd+
iW7F2xsr0ihiLljrq5zoTNNaAeQ/LQ9++7Pua4XvrCWRwDkMd2SvuYwnHatiBytBsVfL7Wym9JfZ
nbLxrfMrA7MxQMZ4BpGoAk3cHrQ3faPuWXLP5aNanHC8QttjmlDcVJqEZ8eAFx3X8PYjMx/TsAho
fmuYumLq9jgOORgXTU0QC5YIsAab8DgPiVUvvftCk+uMyIcw/2g5ZmNZDlocN1XlF7/nemWqWmlk
cN+zEJ+6bXRYr2b1IGA3C/YWLbYA6xPOeLnT8kxwbDOPmxUaMRp9kc1lDIrwkEkg5ZvGX4e15a6y
R8qg+hP5MwDjxBOYLxiV6tSGNaQiGNTnfZrJAqfYx3mifpo97ngPTHPoTt+ZjxrbAoI+oGWeixXO
pR/i1cZwIqretaQBUlZA+zXoAgDNHzICt1FG2Xrx0+lUyO8DtXvCQUm+I7A8tYnmImJunWMtJ4RL
hCjboyROMHBKBbHa9SHc61A5jfM6tE6tVnHkaI8dN9wRasqhV4uiQhLW2sbxuqIH1PDXva7xCwFs
Bxj14ROPwVJ2MuUKlvJfm+71yyOumnQUrBrFsjDqGtuIsoccZ+1y01P7rlzSB85ovwtJLvNcdFTL
iqkWgRWKj/bsz2yl6tG8niXGrQLNmQv1rs0nXYHi/B38S98CpLNlINEaMO95Jab2myFnQUEcdMBU
TlXJUUmFfecXj0brLS4BScL+CQsDe7480Jdka0vq2wIz2ikB7ekXDV/VZ5eQmEt25CCWTaXlrdoU
GBcqZ23c2ZngJsKinzEkytvqbuQhIdD6MTdKNRFIf6cEOT+9gEDYsc7jCuRfbTgiPsuTmfHuaYuT
qSJVNADCGWDegb4hZSYHRdchExmYzB9reG1xY9HrMtPFZAHdOL6DVLwOsBo+WGEZ2QRcGn1ir2ht
I4v4B16HwUSjOr0hAoRJ0R7WIx6xnqNPdb7F9xdl7Gx0PTbxYL87XucI3b0xJ+dCKd8Gi6z4cH8Z
dki53IU6oVdfDJc2Qsl3M558uSOhn8PhMPUCP0SZXYeLY1XeydBax2c36V3LnYCRM2WkfEJYhmLP
9aOHOSrcAMG+ru5yP0h9teuqDDhnmDFeKoZxTZAzl2+OJCIZQzUkicbsdRJz6fHtYv0tqmWkYWA1
Ha43Jj+QIdTev3D+tMmuxyG3iRqCAbNhAVhWvq1N0S3/l1r5KsaCwwe31StFM0Y+9br6SBKmseUl
rO8Zcf9MkKOXzc3UuNVTh19tVxX4P23ogCa/BP7dtnqdbDsp7JuVbi++5R3+tHoaBD+a8xoAz1V0
HM88BQjXA2gnVuQ9BYYJKQi8yY3ZCgoMZNh353ORekvfTual+STqIap99ckydvYDgb6gRwq/wa9w
s2Iw1YAjqj2D3wrsaayQUu8PDqbugd1Wa/ovHRLg/pGlm4MB2ElfOT8joKnjSQNQYt4LuWN8Z8tv
q78ueIGYgfF8ymjSU0/1DLZm0MG5nDq6JrRnY/L4H1fhelo44J5a+0PBnxHZNfXD4H7ZNGTLxWo5
WwrzrGBQ86gmH2zqH3UqaDwbL/HyRs6oLUl36NiVEm4MnRkzyckXjw74rGiUwmta03f4M7tS6Wdy
2vMiqPPd+kkHDBIsWivCrEJr4kzGbKBB4rf1oYkT68GbzniTpEsaggTMi6QChXWhg8Ru4+E1dIYv
1afC9QCuRsigDiiTupWLbsnU96yf92qgHz+NcwAktv/CQxLQYGoUTdsZUsZgP2x71Y3JAy8Kd4zD
P16JSGs3e6bMKx5H9N/RQc0RctfwFTSMAdUZ3uQMaLmVKoOkRRH7JKbgTzsslBoVZETTV4l5xHuz
VkJUNUSUZluzGPV7Yz0vpnhXtlT9beh0jjDH28UPtUrgJFIyt3CB3+jSS0LhGtGxun3Twp89cD/f
8tducah5ARzuRHa8A1EJltNK0Om6CaOLLlwB1GTe5tBH7cuxTzCo4YE7Y28WEHjRTaLTucJkzYG/
hl79h9OB4lkIscSsc/NIZAgTPC08cpQxHUzgSq9IYUzvNNLX5Cor37j/pGZKAdpzvGrDj8U24ASB
q0eeKmFtlzuCQ508c8/3Plddpaq9byrVSNwFk1Ta3gzstN/9FbPMvGbBsVN0/cM/WXzvnpeSrG8t
iBWcetvFbeOJALDWguRN84wRImpqZCltWkzfKzepGOqGLyMgcw/n1oz6hd2ujA7lOAwa9Qy2yO8Q
fxIsGhjJfDq8sCBxkuSRkbfualzwoPPGX+x2MWguWmlxanZYGaZib9FFcqEiSOykX04AkbEhOWbl
k3gA3bSp6Z+tQqcUiSTj1aU2M2pmoftqEVMN/MQVgf2cHrXiQhHdPowOG46j3ukEk3+l2Np/cs3c
BzYnkfaJz8MQ3TFW3mJ0Imluk/JRSOCigiRiyh8ARiIQsoI1TTFnPEgrxdXnogkzsnXLZpZrzHVo
O/qMDOhCeUVM+gL/IA6EKUpUnCvfAEXMJb6PRN8bvk7RL4XDOGmdv3Eio1WE6KG8K94+orzxYz/5
R39ZFOrU1qmDKXpzWJSOuUWj0MQtp4EmkpqZef7zNxEhJIKJPEMmpk1h4HFETUWHX4uUJuYYB8Dm
xVKaaqIYrcDnrK8IhGxb+mzYZ41vAGrxah5ZS6HozwOaD+D5gSVMLIVeOAlZsOL5VZi7XRlBYgMK
x1hPcOakcOO8djWNshZbFsd9hbFFydPyHcjI9GgalLNrhRqPRaDi6hpXRbVIatdo/6ThjDGAopJ9
UvSYbkWko1E/yL0Ww8yJnKts9fCjck1VvL0vru79YN+IwiaCas05SGWA7E/pd7fN/qCNkPqDb5cV
bUBo9x5bTaMto0K1rvXeU7YObthFGPt8X4ZBwSNodfEYWZLr5BEeWTgzmqNUKquXr/Rsj6Rf1fOa
bEFMxcJjHchOwLCgHJGdJZWbUH9w5gr1xbQogYnQhc5UMCkIV9NFNo3DtpZAXSA3st1SEI0c+Z37
idMg6bdK+Im+nXg0Dq7Y0Qd3oRWIwx1ovjDbMfaRapRtcS9wT+1YXLDhd/wDDO9GD1C+CuS1WcXx
4xDktUHgzhWDgbBZxhbeB5puxqypq2zkRUTIS67FAvsyjOSsUhxsQhQNDZ9TaFJJyjUQt6ONLcIu
FvMYJjVLoeKoyWb1cl/bbgVJhVOg+Htqb7Oum9wxgzbQANgpFRB2Ct2rumE1LWEMCgj+P4kEHt6C
3455GgWpXcxjgQMrG/j/bFwr9LwqQfrmCAT3sS9Fy6a1y2CNHvNI5MdgeOm8eCk9bn5NUXTnMBlH
B6zZXL1crQYFGaEw4TJV/tgSIc1UzHDaPch0iHKvVsfQSSY3vaf60DJoNYve7lAxSvhg2Sc88UyG
PCWgx69N/F8aeHbybCAJjDe3mGAVagRWh48U1LEQ6PXI5ncbQ0STJRnygh1hESps9KrGydZXMeca
mzRT9zjnutehIst6GsNkok/rmWA53oNuGOmrTQ9M6LxQri2bslMRrhvXfM9GBllORJhxzHuqdcWV
tIgNZQ6ZvfCjd6z5pply5o3DGuJLq3nu1wy7ysOzaL8q1JoLmURYaDaQ5XEaTVzKbhsZ2yjpqY3v
tR2Ve1BjDVTUIE6/aeYpB0+tmxIxNI+2Lxvjt1dXnqK9XR40eA6dHnNuX5Z/FcKwFysl8uUAyeOy
qOh0RvcDauhIldluXnVPY0WUvkOqDqr0Iaz6ht4xa00cV+tJOEajQAirAGcUH/zJKbnUQOm3x0uu
KjmQHaqW58xkTTdg6JbrqcdzS+xXogcPMNFL26ozwhQ0d15JOcr8Ek+/YCrfnQQ3LXq3XTGp22YT
HaWhaybY7Cd8x4gwuSPR7Lna9Ldh/m55onp1zA/RIYVFkhNjHaKtccx/oMQ1WUbSOAKvUWRMbJ/N
dXVGArvuht65Zx3itEurPESCktoEaXVPe2ocyEBlijmFQsv2TVj4FVbQN/DBboN6CBLOnAfFaR/9
rNfvLbcjjVQqLpV9UaectcNVH3MT0P1No0MAnj8V1rWlYsw4bFBf091l92aCXCedSI6RNrDkLTEM
boWMMRW6ft/qsPWlX4iCFkaNt5Jtm5CvwVM56b+WWbbz6cjP/u4w/Uvv+wsCUPuy3rjvX0FM92L6
uEGHaInVALWwYaZp6QArM4Q0w4xs48VyWRwNhesbSY+6QoDoJqwpCUPYO4KzAYLh6gftncLav2Ai
wCcgL6n+qOOIXc9qEfP2OdEY2TxI9XlAHwTWKcM5+HG+HhUa+mQMqNxCWShZexxtAAynxPvX675E
aQbV9S4h2a/GPR4CEBu45EECEPuaOGqV8k7jsphrZxPlZWK/xDlybfdt90NDDHaTdF5Pjq2ueAdT
cMZkta2ngLVE7Cxh9C+tfKcgHPssin3cQD+Q/8qMRTRy+vw7qBtd7206PBqEQU91uGFyFZEK9Tbx
E0jjPm/FEVBEo1AFPJ3u3p6FFZiUX7XHxzTpXX7zocDKZki0Wdc0fRjmfVFk6+BK1w4qfLSAgR6B
GDAn851X4e0SlREJUGEnvz7Yh7EqkKwbnMYPnuhKtEXbY46UINJe43UxS0WLiY9y+vdlD49/DDKg
anqxbOtmfTaOF7TIb4/V4Bw5LR3mK3tN7W+TBPhLe+S6nMVCN9JJ5olGutmFRIVkPeG6/A24wO25
XlUOvQqCsSUyol9i1EVCy1ne9ID+XqN+/6nLmiBMJz61af5anRFl4wahED39h/EDQMLHk6dTAevb
bd6zFZjoLgpcQPBbTrIAIXpXGFE5UDjqjGXvz8Saf6VMG8/6lbndGBZiI3CWeHZo+Z6F561DsixL
Nk7eiE/PQn2m/9l4L8iPH787HYB5LYS1Rknj3ugz0BE2s3sdWqxyFKClw0qr6bUaElWrcZwaW8+m
MHVEmXfCAQ9WoG7O/l7VbnkCvbP5lWtL0V142QKj/qjfYrZFkVTK+roYcJDZbbffNPCfhwq+gQGH
Xt6QNylZIFPoAn/JvC+v7+XxH67pPekb0rT1zASh3NuY4ZBITUzKwRYxXq0yq6v6oS6tXYe9kcpv
BVjJqt3ssum0BOttRRnPTStX3Aw9Wa9EADmfOJ9ymntILkvcABapp862VSsqzpbnFWQ7xJfj91fv
DNcM1fTryEB7yU0R72Rw+ZgO/Z7ZWdLF7BI31sw5NsoBIlxTe0qXC/KqczUZI8DBztUL8XzP8lvt
StUdEyxWs4SRxJwoWcriNmXJs7dSni+AwhQvGpfEmcty8K9e1HCa3okgI5I7qmusXSf5dZnfJMF5
aKcpAy8DF4l6rIrRGdZtip6idG1wIYHNw8IrWHuOS4TeyLLFZoA2BT/+pwkZp7RYAYhZr+mBlNQk
juFEVX55yQrxrYvSDf6/7zGt+Q0EicmtAUcclilGfDYxQmlEZEcIw6NPE+vHT8MfwB4ubfOysCCO
A8vAm6ZMiVhOB/ylbHqRnq6U6tYik2FWLd3kcbKh7tG5Xv76T87v4WGou3clT8zJ/n2rS1cF3xyW
nOZ3Kfy9+FcFYpepGLQaSlu83zN7gN4SUX2M58KwigJGUHIwgxivRZMUlCJSkKCaK/j9zdv0wmB3
ZKE8HTw8sLejCBwCqdjmOgaFEqx4l/sJg9GOvrlshVGcFRssYAP7n3EcZuS4UzR62m/yXiSuBwxZ
eTlwRLPj8YmoMa1/X5aJJBuJO/AJUcdelVG+3SAlgwLq/kH0VLAxUlzzMe5V56Bb9XjlNm5NVHy/
oCXhVVWp/b/AxSGBSNBFvk8TwAXOy3OWlaAMFt3zwi5HkoZkh1Ow5nCSuo+GypPfsHr9MjQTUTfi
YexDzGJeu1BTWU4fNV6QLt2VWEfZ65Amv9D+YrVLned3vr+CCDM+FOQtNPzQjAgpblxAJpR7NcV5
YvNa6mHJYC8ESQXPKHqnxD7NeGhHTdhmZIKShRFeLFyFAbJ4Yuur8WHCwSrYCiqyEaBmYmYJ6rEs
eiw7RKUvNF0hH3/3TeAtArH5ixXQD+DQvw8pqfeF68iOB/RabYYzL0dvuY642pojDfQHosUGvbsU
hCS9SKmdXOwuJCWCb8YyHLT2XRSN+bqatB2IyKh7Pnh68wj1+pfxR4SKb9Ap1VUMSlVUw+KKWrGT
ByR8peXBshwH9I3m4s1rUmzwZkwhCJGiMvt3oDoNTQAo8ti9klE2qXHz/up4seBlM58PWV2sYQdh
35htI3piMceGT35pds4D3+WG8aYm7XFox+MG9y42XfPtIGDTb36015mNmheDqO7TcF1CRQEMoZWV
m/lWIlUJ9HKCkCjQGUk6IySEtR1zot9+vUdaMS3+OLFJeA4KU5KqRGYGB8yTjLc6Yx1uu7M80YoG
+A7r85hYw5DwY31wXTeDhMyvWuJWg6lg0hbb57zfZ/VvOs3VgTnbof2uVXmJfjl/lUF0JDZIKtIj
rZgou2VvJTrIRFP1z7gdbnVZx/OfJDQ/TiUiv5mnjw2E34ELsFbB+oS+E9DryTSuJprbZM7Ntx6K
8HynCJKwKxcbzE6ZtqDiIo2dGR+glvwfGQPuRJ3nu/cFNOZwlihGuf/8XYaihzsQEL9T8mrKtzRj
Oct0bXg9Wn2GnkVLOvZ07X430uigRuOeADLQaZpmvPL6Ll/7PbX3/gkb3rTOljl4cprqT7sCuw1K
JxVEuE9g8l39qlXf55YPaRtfT4sM6lDk+ZehA4mNiC5K/uR5WKGvNd+ROpN2QhRCJTuVVTmujOUy
FOUOLo1EqZyLEM1DQ8xuobAJbZGf+ymn8OQ/jnVS8Djsq7wsxLow17yg/A0x8W9zYSrFeDQVpcvi
dnwHQkw3zzRtf9UWYlKne/11Xv8kLP+Q9oqmg7NNWoun+RfynI2y6XIe7QBFb2soB/Niyx1aOsRa
Irh4VRC/uqbpbqp3AQN8Cf4xE/iQpNdFRGlg5kb0i6Wsy9I+LNMgfaIJUR70qkF6b2ioA7hk+h7o
BWRcOcpkn4JunYthTFXFQSBMBC1czbC/e9pv6CQzSjfqiKoG/seOX+ppIHmTcU0g3nhmmctijj1n
ja6A5oldUZHe/MH+3x9zc82cvHvuPML4UCJjuRE3LZ6MEHsJVoceJ8KWX0MsmordjcqNz/npediC
eg2bmqGgkAu12ooSvHyUhT1V49jrAax3wP/YRBhOSJ4Ni4vcnEdZ8g4ft3Pe961bssOnIPwpypdF
5Z8aZuGUqZe5cWdC/syX57QouE6PeuHBBvtRviq9yhTw/i8l7gSxCJhVI08VPgTVYARuYaJr1jf3
bvEiOdh/DQEmnpR9gducpPMZtiUdTWpau9yW2Rg09kx52L1u3KXJstezvcYiBHLmdiN+tKd+lNXO
B7CIyRdb6HMUqf5y+J+pUFLRsO0HktkO12khWpMWDi5Yy8DN5wy9enuYZn1k5dmnR8Ro7D4Q3cG7
V1FocmnHbOmMFM6ADYTTrnn6JOY1/4uJjQn61RJWT+/1blKsYssmxUL9ypbc56kB+xjPM7HI9YNz
JIvKNV2rvL1ZuqYY1bCwTh6u19uVEiZNjhieV7XhL36Bmu92vGlnMMrhns6RmJd7ki1pUZ/q7ms7
7tQSsYFYafQbNUUMteeIaU6gnFup7cvAnFgfO58Gil4Ndll9dJDPHDAhfu+O4IdAV+6/EoCyuBqO
UaBwEHsBw4qeCa25jfGlTDuYPr4kafFQIDXsVTMJ0NdHdz/tN5OFq447rZWmJH0/5/9uCBgefK5t
tg9KwylkGNIWwHKBrDwMpnE5uZw01J0OE3t+3H0ZvVu/YtKMcdQPgpgZwLQb6MzZN/FrWusB3rIw
nf929X8Q9+uv0QYfcixYcyDmp1Dm0sYLgLt1Li9duDkcQgPcVke4DiQc7cDiMXBy+A4Sev3FFyCf
Bf+FuO1mmWUjL28o7BL6K20z/bL7J8n42iYZ6shArCPbD3wxD6+VKjAoRVpMXoEwklqEKdbbxiOh
HtWZNNf+EpOjqnt2rD9I3LCdT9WUyDW4D4lM0ViGu7CgBZLQknznNT4VOKXgP0DXPL2s+HAQKKfY
CNTR7Z85hL3py0pOe93LHQ1NTe409NcxuBBvZxY3iVqxFcHuWlZcNzc/8heSg2qws+ACDikRsmEf
9eUFKv2BQe32gfiM/V7eCbpbqmK+RCOg9aGa2dw/CPMUCwTh9mW10cfTkBtalP4LQWxzNLOddc++
Ll9plt3/hYEUgJPfYwa9TgCoh4bX1cItQ7fRbToWCQk8fG88OTOYJX5IhCMBc8hqX8InPiH+NPOR
AktLebelapuf4uEhb1fQ+CNdGzkwE968J6tw25Jv2FM81u15iLgIjNPuc7VWccK6RHtnLQTZlnxM
BBUKw4goMG6+c3P0Y+vDxiDDAAihrziSftwc5p/X7m8K9ivvHZRK19J/9Od7kkr0jugVebdT931Y
s5tvgFZPcoUj9N1ZxQ10gtI6OrH+WqXTVSxq3earemSmIo3l4bdcNkAsYV056qm0TmJ84a39A6VA
bhQtKFZ6jkpto4jfXTyebfVgURzl2bsbPtIKvuWveeOX1YL44Z2Y5znqdGxRh7pitOEJRGYQv1IC
O/Wr9H1FIavflF+7tkMqtqL41gzQXOsLQBVGteeC3gbQjO+BU4QKQXGFmi0xSvyRUVkrNwAqzJ1K
esiQxZ5irallD2I+FLVLMftuF6w91oO+arjGh1Q6+D2MnWXi6naDyHl6a4qGnUMv3nPCs9ZDh+hs
moYLVWdHcgxP+7Be/f6zl/TWotG2fP/06bVGO1F5qaTTuiEkeZncWNq24xQK+CKzWlQXjjRHGaNy
7RpF+9HuDyo8g+psSa/ODQuk+a+yDnHssXFcfsysc4J1Yq0jJB8lckoGteY/jozd3UGfzo+jjGj9
xnWIWqoWGJMh3m7yF7pcsmbjpnsxj20+vuSV8uQ4vkJuml/FHMjHgN5RJ8M2zPcDxbb5pc5ElMNA
cbzCtgMPUI2/gx/C53DGc79DNC/Mj1W6tW50lx4tYg/0vLdOfm1vU3nbWESeyRfFEL95TPHRLQWn
J6DP4nToEuVgcXazJiZrYQnw4bfpkvUOgBlCxPE9dY1L9k+2/ejA4Yw2kih2qbt11qGdu2m/ZZ1a
mK0n5bb/K4Gaa7WLqd1YvoytdH3pejWTtZBC21fPiZTeN75KoYdFIA+YZjohW4+pEmLs7IGMyEyf
FfelHOb469GST1AgQxZlGTFf4ab0/dhu8YXYqLE8a7/SVnwPosvgli8djFgxK8grH4TcUPSrSq33
8vcK3ORQvvB/rtmMSJRfMFyc+Ixg2LFSFnU0LTT+eBd8zCqdVYzU75GgFMYicNv1x2/g+3ClWbbx
3CHIJxq4Vj3xxFQrmXLtdlRqxek5yRhZ9f2INiTtTFlWu3rrv/xqYMscQ3M31r+LVsLD9BqfoP0J
rtmQBKYSiJjzD2sXKksT4ytooNHWN7MKawfaF63+19+1MnRcDZTroxxTHgAX7tPDqG7DjjOg6RGp
r/MGJ46pp+wEiVKjHMag0F6CjK6J8h4SiUPqBNXJv+O+ripuNMBhg+Ccp6dEhvI8m19Sb+Icrris
uBu6utCGWR0d57PDm0bKg3MdSROGhS9oUQXK2fMgn3i1j27TLc9yGfTJbLt4jIW1VWm9CG58W7MV
mDLkl51rBG1r3rTr59rIiWH6ZIWwOrFubzKi+Y9+x1kcL2WLE7k9OL64LSxryUMUHL03wDrAcLL8
6bErP5a8YMWAQvbR2uO4GgmXmcJr08ntgI1Di5CMZ4E2uFkV4afA+vh61yz9lCeDlR3RY7o2mq4d
D1pD0j1GwgPyFWaimEB6FdDmTn5NdsxOYPkhAXaxs2KYx8APiwBGTzZKDjmOmhXsnUuzR730AW5A
bbOF7cDV35LBfv11SCGoJty/g+A2V3d0wa1V9iQHq3hAlyOojkWsu87arwkDQgquOAxjGXsWn09q
SImoZf5dOaHxstlETT7I2bTnOmpTftx+gbTgkIVX1MiJyd3n4MWslw+1nzwDDtJNH3KnrGK/HIfu
YhfvICuyl7YXCC4ducN7Od6Y0X7tjKsC0EE46/3unHseSNZmnb+8Iz+M22WZNP5a4r68uXFRwksd
2jQhQX2bm++3fwbPWT18SvqlglRcUwwy+6lhBBzypHfP8Nh2bmPodcCUvaaMnEa2q1hugV/tJJzs
zGQ2m/nZNtLAqls6uYqM37UN2B2ZHAH9opnHcLL6BH4AWa8ZpjeRxeAAHGMH4zoyiOUOhmezJfCL
tq0t0i16+5rNJCwaLgobPdauMR+wLV/kZML7cOuxUmjcH74gPmDGE0ViaAc3ycXncmXz10SFKF5I
SLWQwUzDfp2oYrmozSdV2Askrhzo1knHEiUnWgYLBme2ME5nnxJs1P3rAXuWS4AjfAQzSOS1LjA1
FytxW7qzu548RlSoAtYr26uIcQmX4agmUyj8YGlFfDlldSpyTkdXcajqpJZIQLOjIz86CK60iziu
9XIyvIQB9I12siuSk2d8D4D25DhT8VFnPJW0qxaiHNvEsFpO4IgeEz74vH2mH+x/2tmo0Uu7pJYk
jgtt0CC0G5uVQrtZpHaFyGb++Q+AnVdcRjMb9e2R9k1uHxWOgsKYrlcSkTUHnjljCudvlEV6ffXo
lkEpJD/9Wswt2oHNr8YuAWhnFv8QW3KHd4Z9hzRA71lEOWJMfu+Dqvjzu9eNC4c8C589VmgmPIbb
Ut7pMdcmH1PqLFO6ois9G5HpY2eGl4hRP/nIe5Dlxp3ncBtT7TXQhf97zry2DEpq4GJsRDTi1mQA
gwPDLTypx5KLlVJIiCJw+AGGC4Pa+xNtcwZhzD4yXAFYUJtU94Ew6f+/AQ+G4Wa93bieMxkLq1Gy
FOC0eUq8IzWKv6v6gv7m99IkJ/SHT3hTEZZVAdDXemZ+fvD+mgZol5DLntbR5MOMqYF7vX4QF9+r
Vhy2DrsoTNDx9bG50HLMyryk5eryTO9Q2hYIVvlnpxmxqZ9AWTWAxkT18ZJYXyiuf1rFxGTFwoNR
hxqTIf3k88fAMvB5ILzyZPqMLAqvqL4l5pbzpdHuF62JmChUZgY/Lsrq6p4kguyRuS40kemaPZ5I
Mh8VId1G9UBTo9SYdnWdkMATg+peU9qdEx+9/aZoUK90fAqOq+gGCsSWNYGsfMFyQkQ+KA0udkqU
M2GuNlTYwL0q5i7w3y1BIR21Z58SwU46918NPFTHEfG7ufqeJd1g0U0qyidJ/H5Br916sgZtbxra
jJ1khbw4/cJEaIuCXnUUMzWazXd61jygDVG8fFpXSOAqXcR1A7Ql0G4dGKp7jx+M/TDZbK9+Crxy
+B3rbpxBHNePcnZ0orJ1hXaTX2pryWP0tFewSRas50VaTYcvCJTyq4fiSf7xVv4IizNAlKS8zvWk
NvhJ2WMPsI7Or++xky3OmAoAhoF17Wf4bpv0RRvjBSCJX5oS8NAmzJdIxYkiRoQ0+n/LY1wDK7yh
Al4Fl8Cznrgl/ekWG6bRxjNG1k+oQHmAD38qN2L1ER06r83aC58f8Ciq9SphhK7ZEo63pj/aFWRM
q/OTjitsSu7Hh8K0ivH0STYNv2VsbLAYvTAprCLlqmIeMbMLP8jWP9n8SRovnHoclOODaXkCprdy
sW9NLnHeWTXEJWXqVwcqvxU9mgi1XWCY+dQp505ZQ6VMIzAlQlQQSn0Cgi5SU5HmoK30Y8mUiXEq
WtikGiiFwcNiQF4wDCP9FwzbRacGo5N3PW5Ms9YwY8w1pgOfY9Wi4pH96wz3Kqv43sVtIff9C8FC
mPRRGjeC+LRcxE0yKwYxjiAp+zxa6lwUSChOuN+LsZbxiWlCtNH6Vzd+wU25GiQ33ZV02egDGmb4
RKiIGY3XIy3DYbeRLg+QSDK731x5Dt/Ur0SwFvCrASNmdPteABDPlP0voCVm0m48Ut0992x6xNKi
9JdeOwNLefyAO64J66jJSVcUNuCmGWymYTxOYdxG5VGw9r9J3wfVsCszTmhlRBMi//6OM7JOIzP+
Tcw01cwZJgFqIV9UdtXr/bzVT/SlHPibwVqj22dyOfXiWHoCVZfAiUv/xOwIIwRArhqzrNJPyD+F
JoIly1p7rzuhAsSub0rAqV2RMOmqEWu3svxrWNJefU8ZxzA5pRcY+jETzU3eq2tWDE2x2kw7xSMV
QQEdDr2s37OrCpy3UF6F3anaFa3sHpf4fJ8odvfKosWZgbrG+2LLw1WxjzOxggAAVKbN497SsUtz
WrjJ+p9DCMsNXg2mqK3A8e5X8gXQIf9QuVv5f6yVdUXMxTHjSdytdpYzrrDzPneVPxY14f/a60XQ
4WVNMTgkZRFu4N+VPQjfee1+nAb4NMaMft5m9IHW3GQ06P/Bxfuw4dcLx8ILUPQUJF92cNRI9Ieu
SwogR3gpzFr6MLc/PPlAic3bkrF0dcd9l90AegxjPjQ1UEB9GqC6BV7SUp2OSNcOPQOpTRva24Zf
t/cs0Y5XFtMBvsO+FGVnKQBkH7D+qvkZOE+Q3oECGNjt4cn9KaY3DvfhyQa+ACPSRapmhLrtStqA
pYroGxSJ6eKJfDKft3ROAyqYokPOlcr23zjkK36evc3/w4mhFDkj/jfwQxerWqRkrGDWe58qbDDP
GkCqxiSU/PGr8FR8B4GTmCRoG+zKOrkJS0xr40rgEPofcoC4OZvN+RiB2Ru3S+Xbvx7s9FukFN1L
ud4/DR5KIs7OlRqasrwdN6mKZIK3gUw6lC+0rkmKz0L0Xv+QXZmNbFrkzSHET/hfdZtRbwlSBX3Z
jeBav3aDR6xDOZZLl4Fex3kqBZC1a/bvJMHxn2kx8XDLdgrrvP1HBp91UTT35SjLaaikLt3eVl9g
sR+i9rBj2cCQzLMGJd+YVdW2ahm9n/wOCIR2hihZUqRYTI3tBWyuoJ9/LaTgt/aWGmclBEqUM9Fy
HtTgN9iVQmAfpAFTJ5r4wifUzxHX+ZF2+Kb+8hOry0fSpMmnuj/CpzI/9VCj1kWsN1OSDrhAJj6O
a12pL5zzwryE3eVKyQblNh9kTqsTpRhX5WxsQnUb1KiQpHtU5hWbtfQwoOv0+Jo7iH8hk1YbHoMl
RKdubEmcht3dbromjknrrUY6v4/xbudo4fN6aPZbbIXgEPldkXSKWIdwtcW+STwDTPqR+BjISG2d
RkbDbTpf/NikuGKDAyK4E0RJkp8q4iv4mVxf8tPpvMLOl48BDECARXbiZPqhMkXo+iJMOJA550el
zcr52cZxxqvmdHxaFTA9Nafx/Y3S416pwwn/BBFTIdOKHv1inYrOZbFoc9wxpxTT9XT36Etu02Ma
7dTUBjMf6cKZURKYECpA0tNxQI58gjzPcCsAICduEQhP9UroFtWITYmk2hyLAERTZpkwnV7CxLoh
vHWYUylYJEzgSmxmTUIVoeqptUzYn45y+LphfGWTtn4a78jHsx16fiSX8zxojlvt1fdJrZLSOmLN
qxn3rZ8AOB4l0ROvAvpR7ZoAb4E3u2/yE7hBkCq0mzXU5bMqLZVjwiR5KtcJxPRrJbQr5XeGKnOq
VyzY0wNeqFb+nSU1nYQon+pQpec2wCRY6ugfUbcgiYO1Dr0xynxw3KceBRzGe/q69I0z/ex7/oiw
x5rMlkHZnzvo1PLGAiWXgKOwcvoZF2y5RX8zlmmoYu8QtREYbRsrtRkOrUspqzzMh+9dEAWDYrZR
2eAznZYSkMsbgjziTXrFaE5ayKZ09+l/2Hw66OqZ3FoYP3ONS9ImdJ8EXbnCOWzKDb/bUXdmFBUD
U1tcFywLQ6OggER1B3W+NBr5YAHED3NBA74UcjAdlwxC/n0WyvmYsTIQ1NS7z01ca2vQR/LJYRw4
7f1rIPdHLz23QseS7c3v+npIlkjvbCVvly1I3AmF7nYYc1emXtRjLf0tHxKIs8/qgDju58RTQxSa
J+MYALJPPAfoc1lbL8W/1/JU0wssdUPH+mLmmYPNasb8ODOa3w2qXuk1WckDehk0Kfh4Tiy3TO2u
9us8ucSqYOkKIoHvpBWkc1+/KaMk8Llc8ZDgh4Q5bHE40cM1QLak5b7jk3REuKRch5UDbEtdWhf3
gFj/fqtAFd6c7SybHAdFCCLHqPeKIOlrWriyPqTvwZhvd5eAXMV31dgYS27wJOm5jqV5RzLdHFFl
vqklaXZyoEL97T7+bahSmIRkpPuFL8l5G7tSm0eqxUV6hCQMl/5pSVCi3BV+3tzyHdd/hEdtlghD
tRvrS0yOz4N7IUzw51X2tgAshC3LJf9wUzcdRo7HLWFULiyC6zkGIELX5dYmvaM9R/lfvNWpumnU
3EzDxyhiHYar8Z4isgtmz7zQ1irdXbAR2IX476rMGNGTPjSpgcmfLGgH0qVmeTut48ljzkBzJTBR
tQzHV+vtB5V5iGTX/R2W8ZVlSj8LNFO36c4yRL6f6rOwZizh7t/Wz5CiaroYzw6ora//+34RAsGL
PxHkYmCKBjXH+ruezFnK9LadMjUzO0Go9vudTe0sCaBUZFiGw1D/3OZw1X8Bk61+4SK9ETBGcLUz
obsEi9iP0nCS2qZhoKgvLSbrlUT0UjjvgOzfgQbGJRgB/SHdeFDeR9DqxtmzvnUGHylTPCp311O7
vjthYslmh+Zg4C63hazTpEJSmRpCN1LuTzbwYArsHPXVvvAfoKj55pvox92ufMP3iruJFKP410Co
BQfswGwdC6Fc46CzSI4gLdxgn3SQoQ9o129xZMegzUQivXW+pn+Gpwqq/vIfdkoAAgeR/Ac8waYi
w8PLEPv/jCzpR4cuXbRWiGFHI5DnYxyljOKmZy6EH5TkwcamSjhENhgs7hM6+YSDy3SZvLZJNKs6
ZCjX7NVlTclxCsiYB8W7jSlthy0mgskmKfCoM3eZKwiLY/b2K3zNgKbql4ymQuHvdJvxNGtRCU9w
oHNFRnU3WPKg5dFyB9lAuOA0woA3/o/R/j6N2HXFLIcGJe0eSlH2Snag6N7fDHNldkcmerT7w6iV
qJCnuqbqKG9R18NA3xuWEhLwN/Kk0ZygkM5zNHIDuWm/RXjhysZJZ17376aoiXgdmxufpqH/12dK
yOl6Q8+2Fawt08uBapefjSh/ND0hN2I3XOQbP7phGvMVpg65qYAbmxlT1J0ckRq0GUr6tI53/MRu
O+y6Wpddta9l50UGH3proOsje/CCQz52yXt3AsNrFGOJY4muLnThzzfh2rz2X08q7F3p+U7BGMFl
zVJLAGzImx0CORdjwwbAop/BHAoJ5RVqHVGnyTjtWMb0+2rw+gFeGoh0i9haDZeG/2pLqwl7QS1g
eWwBiToDOy7yvEKwCAlNDj2Sa5RZ6IAk0X9w/bUYG571q2Etnc/grTuVlQO8vwlhbm15q/L8h3ao
81jLfmhUXocRpOikD+JUrKus8RDpceU56P09e+mSUGEHTp12UzAqluGnC8ycsnpNYlzgStJTi5eR
aasn+E4Tz2KWCK/9NoB9Gnn4necFhdTDILwPIxm0fpSbJ88YIg1CBk6mmvQvFIMm13Usdjq3AtKO
RXv2XVgGhFRRFosZP31BpnXekVvmHWALtOArBSVnhpbPw6MpNbha6GKi+ecu3oEAUCiemNafkOuH
tatLg2Zv9Fdo9owfbsod4wI0TZwSXj4RSbU/O5W4XyVMhevfA2oNTlOL3ayqn0ykscklU9MQnAGu
4RCYEo5B/931u+ca8TTf95l3sdp0eGteO37AZUzCXh/8WkrPEYpUgFhm2Jtqi20coNCOt3keSnl8
JUwLK7Sop4vKFAWCq1NRW6LgJaueLDl99tgTISP9BxrgFwhgHXSlktYPCLk/9a7+eLGRpuER1FxY
J7gfemW2uv7ivMPlR2uZFYCza4xe/2Kp+EFDLMP4LFTTkMbMB+rhNShmnlh9EMtTyzHcjF762JDq
6v/dX7F8WEXITxKUFXOBSF8K3SZuLrtgpfAMNapyUDgjtDam+/JiDHHVgUuD9rYJVz5mtO4jsyGa
G27wEoWHz3pJK9qxTX+ihcB/DIpc65EnR3sI48CRmiF2/DTogRDdxG3FRCpcY7mJYbHARDzzG6LV
7ZVtxEPYILfjJasfX5wFn+QlAokAHxpUpB7zlIkWGAU2Se6A8GBIcj1PdG7KkvmG6tA5WKoZLOi6
Ov4psIQPlVDIJXUVHAxn2hw1Xq01g+VvmUMUf9vA0GTX+ksaHaoP1/uOndVu7WWjSd385VsxE8mm
ulqRTof7wMrA6Y0XAozL900RuYL5jOPOZlnhjpuP7b8QYlGUgxise6GKyvYsWVjp3X1k35GwUvoO
nD4bkWHnEklArjmOmelsck8eYzuLhGWnZw7NH8EusuNINRtanLAr++Tq/UMKOK+KsYZ/uwp3lrEC
VdpY5zF2irO1J9O7WcMzfIzScb7nJ85TW/UhfTii+bNV2N+CHwHzh8jiiHxzEQ49uclrXeAwRdNC
GM5qyleL9D9dbqq9aNQb7dmpoMXFs5Zy3qI0k18MIOfaOQZxTqNhoph9hN5puZ+dfs3PokIMJY8A
ophDwGmTvgJK2ssk6IvuO5fKiCsfbbqzJeyH14KVYPhF4RdVj2IHG9OA3hDRciyNIa82UKtd+2j6
RDePFnpJB2HD7LH04tNyM0EsgP3Pt8cO2V+cfiWhSFP7SrZkOyfleyYkc6LCvY73AqQYCErZwXya
Rt/VqMb8G0VdZK33+mhF7EPl+l13tp6lNZ6RdndSq6AKngyQkpmePc5J+n7FAzqJrSC4Pf353ivH
LKAvmXuUn/NiutXjtABvdf62fgBPOPuEqJz4Qm/j2ZVqZzdVTP27E2ySisXkB2qEfffhszpWhtzu
E8X1R2DZ9/ui32iK7UvWRnPF6DiSCuaZblvVWg97mFbfgxR2Z0wBl3kv/YBw8yuN7UR8aJfyCop5
j24b3B35uv93cs+PVClipZxNb6uFrKeQZt3LCq4ckw2T7Upq7qJ22zqsiIMXbE9z1mfWjHClOAjt
nw073ADGAwYXUOxEUIae465l0BeMbf7mFLLjA1/iqeYuh7MC8CYjYLLlsvxrciZ9ns7YogOImxI6
gZ87PMxWnzYHujmVcjyRe49RuNC/ThqJ/Xo4/RgA6XHd6YoXpzw+iuSSbS+KGa8FXhULXtwdZA9R
Lp2fRuObo0DXL89JUtZyWQtdzzYtzR9cYMA4B2vtcIZAqx5HgW395/u7XfzR43es4pTJftHQLFeL
ZrLfjhk0kdfbSYJAjODZ3QlIzqSFWOwvCu71W9gwuoAc5bn8ct9MxR1kuaqqwSHuhZ3dhiEO5A5P
FwkaYp71K+v96qaOozE0KfwfSLcH/U6tNQLUDCeWef6A+/F0PTPberlyn8DKd/30eAXy57V2T8il
82gzvkJwZKAZy+g8Lhg94hZskqDSUIEJUHTtew+fTZiXXWC9WC5nG0Rm7HlLAc133Cv9It2Cg3U1
0JUPJAvMv0ZAC41nBrJvXVKR5C67SzZGqHuo/YUxLp1T+rAlKdf3EpPOxz/q5V2zhCZ6IDxsIMOw
5Oj/UCwUaRlAR+i+nIOpqiIE3vAJfENJWb6szE8daCUbJh1h7SRyRpN+id/VDa6z/KHqnHoJ5n8G
Gl4iC/38JuCbGCn3h3p+1rlpqKRxRYqRe8RZ5XxgTms1hh+0J8dbrHEAc3FyJlyIu9yytMBAzfpE
aF2jNCh80ujuYM97mG/udM+zRAkGm5qb/dTGjbfJ+0cCFyoSNyZAQooukV6d5QRw2FZXLBH/7X2Q
TI/63I54yaTVqqpSULsAdYV59yCGobpUpvtN8hzF1+XCWBXkCPGL8nsPvaT8PRIaihqUcbLeG3kQ
6pIIMXwIyHX0CJCP/TyaQZFhw+ho8HKHsHAto1mwMTZmQelfMZvc3dXpqrJqJlca/SF3cNp3G+gD
f2xljgF1Jbo8OWB+M+yWtsXL3rtozPUVgAI6dl0Op51lqPXeuQeBKIP/ctEcaqD5cZp2xfTEGXVk
OwEBRzIHsSj+cObLFHi2UaX167opFhd90xitKf5qOgfPQetNyVIvuOzVF0xk9Ch492R+giox5iAl
exA8u6/iWvXTg01HvH9bWStz8xePu70B2Heahe+Pwb2pyjxQg71DFSJD2avWH4Ctk2GQRGhKBzfL
jMLGP8CKZjKabjqbSHZt32ZNZpzSZMTt+7EuO5jIPTh2Kd/FA7hREFCUmra7bLLG9RRtf8/WdL2s
etAr7O/K/45S5lWYfXAGZzGRRLojRQzlXj5owdAmQS+wzFPR36QLAKhFo7zVy/o1EaBwEaOdNt+F
YHXqwyTL2kx4jrjvUqp3Xi8nXVR+PYyjj+2Ee6aKYnVwn0pK9dP93bQi0aNCGWCWKs1O2Eiba9mz
NeNS+4V2el2Kzfy29Z/anwMS0FTNXnnMGsy/05p3lzOBfSMbfemTDP9/Az0PDGJoOZYtg/4lOIOY
r3lBWOxm1LKajwTKFsiQprNAgoQI8neROFT7L48jPMxlOh2Gzrld9iZ5xoISM7S2UcdS33GCSzKm
+CDOUtP3Z2SSDfEtZk2KHos27R8PgeTnRjNLBSFv5yY+KGcB7u8HqKAkbJykxalr2SvzDtfgmHtX
dK0wNYOxMB6ITzHEgcywXDPaOA8QLTDuIhb+/+qZRoBAm3bsyaFczvXQJK0cjo+b3gOfIU3hYKsk
1pTz9OamNfBC7SY8on78YX96QX8bA71QUK3F+8vviK52wRk+6ydRYFFZsJGfI50hwpzl4d7NyoGc
n59BKLr6sawOukEdTPuYIi/bJjqvCRvd0o12PzxRsef/kIkeClWYz0mPOIt05wc/vkrVfl/DaMW9
0QNzPxK5eMsw9XN0TRJy1cRHtLoRx8EI40zQ3ZdUp6sL/Vaa/J31ibYbt2eSIstTjgJ24zuUNBiT
TWzR4Kn99Srs5HWtigBTAmZ6CYyvVAeOXZhzf/NJaCh1zksPrMkZPx8jgOXevmjsj+yjGkNjofeh
tS/41jNelZnAZ66omtM2WFVdFud16ChQPr8mFLVGNBWXnMwU3IYCmXbpGdluqCadoPwele94eBTc
zpzNnKxQu/qYqohY7MdniYgDmXK+hXOfhC+kNMo5zQWp4U2KpJcvj2VV0BEEV6aUqylV2PnrCYMX
zp55ejWiInPmdxK8a5uzeR5UBELiDq+c4kz4RMLEHnayB1/k8HhModewlkdquuAJSQ0CiWF9MjC8
v/5n0o2LplhuNLODJcvzDSQAF7xOwpHZ3k0up+Qh2DnSOY5c8prIrBO3TpW/LSA5k16jfL0nnNuq
fDANfZfcYm9yP6Xmkgf3+D/w7u3e/DlndHd1wATO1d7wm1abjItBWnVERLsjGLwgtjfxw4ytEZdT
cz+5hbVa8cRrZsRV1ALJyPIsXo4qTtzAhaUCo70yO3hbwybdC+3ryuA2sC6w1AwSFYkxzSdSLUa6
TVVomJHdjBV215HnJkON20yS6/YUmHXk0poyw7X79xHAm+rgeDHCiBs/GWD125VLqbpVnPwJtfd/
+jT2j2GDmnQ9jAKSAixCCzS+I8Z2rOrH1NSX57FUV2rsJ+VERacMsZQeOQ9+2ARn5djUSqC6uuDP
wGXLPFjfGfUV6hAyaYmN7gEsZwARJ8Ag8Do+1kUeh/eXFyDb8Cn5HYcdJ6eK84BtGSB3LSuZ/Kah
fIoMUtmW3KHNJSzNyOnZwzWSrtvFQ0saFrFu6UOgeV/MMwljUolZ/6b0cOf8MktBRV54vsOLtP/S
jLe3hDLr5+HIbRq1Uw5asFN+tdI2iJu5VSutlecmDGFotb92ciGWsDhMq7PL5RkdQywspOhhXcgZ
UDfnj+DXnyqqw3crdxp0JNGj7G+rCr6+TlJuoZccumJS7z6Gik7K0y6Xrwy/wjtV7QAfMpgJiI5l
12YZhNInaz6cf/aNZRAiCkOdHRc35T/kFraMpty5MWt1uzG81LQCQQFxdc2ZrJlvWOaqIADWPZRw
77ZYe8YkGjlpZ7CJGTQYV7JCdn7a3T+guK8fbZ7wB4ow3LoFvQWnCbkhpS3F/UyaR7sA31pfanXK
JJS1gK7i+Q4AlHYT/8mnw672w7v2ELFS/093j5+u0hZBhlgY3eYvl27xGFrbm+2wAp+PQfzGRG2f
f7YA2VkhXt4AHpVbdDJqbXTa7bl76Sj4JQ1xuGYnn7ziYEDFDsFPD0zZy6zqeXTvaWftrZgrHre5
fuEcmIfukmKQrWEpovZSuzRXf9aNgHl916LMWx0F0LOjbE1442oXpMBDCH4GtUvmdT3bhooeEN8U
HqrbnD2v+weMG46JGP7tStfrmJRdwOcGHP8vHdU8yhvdvsNaOx6W0jeae9llJOBhtDID3ohATvz8
G65MsUoKEaJVdksmp8gBhUdKc/gmZcz2OZAjqQ1fQ/5/w7bqhD7vVD6oJXb9k8hjanVe3yXbq2Va
M8Irr9RQ/4BWJrePAZyM50nl0k8mBqRTfXT2OmU9BB8IVcLmxn/s2n1lRDVGDp3J8+OXtFYha4Ik
IVsHrVIO9IDt7BeVA/MHjSsL9ldZGxwQkl5I3K3BUV2+hIGtZahNygSXCk8qsWLeCHHCzJBCjjJm
OGloc/PJ/LhtEHJf3iq5P6zPtHGcoLDfP+tJBd0PSnNpvlWra3UrmegIluPTZCvaariJB6UioTrc
NboKtqCDmN0DrwzkE/L67srN6zxyxSVkMdSB9CBANYIjJYm+aMNtpT6/c6mOySUJA1URJWNPd9cV
jZbtlfvXbYWrdPwzZAgvOyby40V6STMKlY2xEhIUISVS8i3fVnEWt7Q2wFEPvKxoBJHeXtDX+VF2
iW87MdzZqUzr0YQ8Q7AcC0VT5aL/fDp7I4Z1o7D6HvMdvYB64hKrQzDsnAQDdO1uFbPZXPCnWZki
N2v4HYPrNJfULKMGu8ufaghM9Rit67CAfVvGTvd1yxsAhjF9YSYMUnIHfJKBrmggqNstgslfKlG5
wdgJOZaE3vwdayPJCHjduWGBh2kSS15N9hkWdOocyrX6Xiul8hWAJSKq9QlTbm0QbEEJPdf+oxDQ
X93k2nf1piDYpLuhpUSlkuCJXIBiP9RPPXX+h+oEeqPvJrG9bkHFyToF7axL04oSlLx7I2Z7AQdA
l1hTtSx9mxn05aZLWQhrZ43Qcq8uSmkkmfHYpUFWrsQ6J4rYQfIuE1tsB2kkLcLuM37iUZxSgpjL
KlJS7zmSNjuUZIWpZFj7GFO9452/3fMjEKMcVMpVDSkIwfrS0Vnxwkeng5XJdCeuCiRr5AhRlH71
Ni12sdbhVMkIMClg7yV52aVz07biRUfxQO0oiq/GR3BHFS6fKsdVKqygCvCT0lH5KX0O3fKI5nQT
LPo8MIIZRI32c1SC2+TfQAyPCUcbrho06EhPoF326YHC42q5irWKEVShTm8x61zgsNLoy/KUXF61
5ZmBPzRwGvUrxR3qYhDmGwzvsaiMfu2R9WWaUZPCWMNqPx/jlBhj+befQTpH8zsBCeA8Yi+oJnEI
ZX9sLXQEUjVuWhCbOYHrKtMjQ9Qp+anlNti8dhn5OQS7PVJxr6+JMOp+AiSgoGm/nGSY5OOp0myw
hh5iIVkKiNLyX81iGRqRiHeUcL67vbOoFy0cUOasHLG2jqn5R1YqlfV4Hd0ixuImbS9b74bYXsfy
t89viP0CywH30+U6/yr3ioOLmNyAlyuvaUU7nc2KRsr+U6PZgotP+8oPWLcLxQN3bnIo/UkjGc2N
k8FOH3A6LXo2cge4S+9JkT2N9DqwcJbYxXkqtCkCKLUkBJSkiBbWAYu+SJgZZnfsxAF2fJaU7lga
UP/70I5YgzsZnPiPRT46VhDLm32ReerLkIuboSRs6rCI2O5DzvjUiRea98rwoJgzDi3+D/V/hwte
csSiYhHnr/X5l+mmskAhRJl0Hj+x9jE/jlF6uVAKB7pX08P5vuMm/U9cci+kNqGiVZ1kV3Nd7+ez
/JT/X+AoYtVK2aKnXEAfPhDEGuJS3ICAJNZS2bTaIx4MkdprZMnMrYVrG3qM97lgmNdy0rBkJr20
lqFBYpn+wwM90P6GqjQv/sjD5YhBvMOVNzvaLKOdike9NwlAa5uxccKblueFQcrzCPZ0BboaW4eQ
Yh7jJx4UYf287yHT2C+OsEwoTtmApTlWp4Gu9B2HsBMDtYSXU8VfCGoLNan+VHR8opSfMBNZx/Bp
64ZaH/TYW+8iMmwSaKf2M9kNCA4rGLPZu3Hv+cKcKk5BNQJaPXyUegkE7+zczaFr+53WN8UzsV+o
mylW4Eoa0tfRnTQno9Zwsm0f2X2A4zmYL3NxbfrLrIFEauznV0kOl1w7eor7j06IRF92lgyP0PhB
40PP3Or8nJkeudNQI/pnmXVCNxeXt/ixs8Oi5RVvNTbikUKc+tMjmC04N1a2huzmFFWhTCR7KFrM
LsbVJqTafOuuiB7jr2iKSLQ4EX5EkQqAXP6p9a2dcwTxeNiG/kZm5DpCvI24fEHzNaPVC+YCAD9y
SETmvcIZZlpCJxZuW2+zwUyOguM8mlv4ly0zN2BTpW4LbVjyv1sBbvsLRdrn9RA4fI1/WWVDpRNJ
i+pZe1+PhpsGC+y7VylYTz6c4bVJktK/CY63lD69N+ApW7GIHdUz9k0XhRyR+wM+PWS542QT1yPJ
IRVEqIdpQJGpYQ9KCNN1RIc4+4tg7Ap0ZIEuYoqeuBfXdKR7GCdWYhgpEBpHRYZGI4zkVI3rsNiw
4gictEy+s+kytuDpi7xJjXGxzx7KzlYx3KC1RwEEqVjz0iKDvBWUcwW0WCE3ddC4l57u0iL6t/N3
WoPw/Je03COIclLPDlOcBeAIFodeCWGQoSW84cRcscheMNS0f5BgLRtoQYk1k14YLz/EHPwvIWHT
1fzs1twk9fuuhDMYPxCSTM6bmdSN2U8nOocxqweV/qRM9W59f5CXtB0opHOlZntKAmi5mnhjXp/d
vx204B+lUCVylIl+8Pl4q14OTvSKrbFzIzsF8zmjYcvJcdf642cZfr6CljRDqlc6IArm/6CZWpZy
mdtjAxJFv4oDzDoUgnPsbV1QYz+8fAVgJHc/jyq4D8dC2KXd5fVCJlIpyGdU1gqQzO0ZIqBq2TAl
QovZ0pUXDuBFlkucEjWKMiOLPPwBuQQ2AaY2Np03gHR17GEoIQ9alhEYwIXQE8EdTYSo2kLd1MYz
rUE5RP63VKlGrzBmC/IQ2zLW+f1iW7mQFKXoUn/wLhauV2AAg4vDFsAqwePvbKq4QXnEA5GWrRrE
WFkaaj2gD/w0ckO0Ah2IWm7c7RVsH/b0bCH9ll/Exc2co+uwLFWQmK2pc9XPOTDaa52palCbE6RC
QhtD9/I/rgZG7YRnwLWEx1DQ/5WPl7qm+qCbcvNQZsXv9QDJjfeTtL5Rs/EAv4h88m9M1ZNoT52w
KsE9nRH06TnnIlR8CSY+7aoBclGMNQIT1buFlKcugmo9WdmIfVNZbF7yWT5rcJmes9CTQJAzYI2C
x1hpS1DJrVTPSHEoM5GtKgvLmiX9G3nSx30Lab5gtiyJ5dI0gLVdGG5Abe7MHI67x5Px9zURWHUD
KAoBGcebf4sBfXcFc7uyOex32rpnCeopzD1l60s6B8DybKN+OhXl7uA9HPfHnQXOSdmZJ7vM1ABK
6Ux9iQz64FMRBKhBLNWEWR2OKVXPNh06FD0Jz8gFiwcSpVQLVGl2JvBr2rSx49sIoPGTYkeFc7PW
8aM9r+O3yi0OESVEYLL5SS/25PlR/8Qqt8s6By+RiolKScXJKStS6HuOnGwEddB6PT0hZ0TVeEsG
53k4psbC77bV8ihToMtW9k59uwdfnno13qvraMEDaJM+WWFE28MEMQTl0HUzz1o3b4RNj78gWXAi
mxlKUs5BL0Vba6yuGekHACis7Umn1UWSRZlsf5VcHneSrUQPnXEUPKgzoDA+XSkGbMACRoSAjelG
KQ6HWai2SiRWn3xcYSQ9ub9QBaTBl0jJhZBr/tbsXuoPCmZPOEcIreUaVAkAj5qAIlaReGG0UaVa
YvXHDGbHufBMpXzbZX2xdkGDo4l96s4p+Oip99LZm+bGTW8q/xjvIOP9nyqNbXPSIuXmKbz0IWBU
hzzCQ0FqSPSpCcGCfFcnIhVExd02/N3EfrYZE4b6Ynk1bZ86x50BU2MgHPN3wmJF0LiiL0jYatZL
Umm8FweX13NOwf4ww79Ea8u3dMF+ftXscyCCuuQRMwi4bFDj6p4w6D/aczmwPf56AWn219Ug0zsh
Pev3iccY4sslPeShjsSxwmk6I8VtuAGxjkCQetmRy14GiNUQq0zOZmiQcu+MsQOeGiBFXjNqzi1T
AjKbDky/pf12yrCu4cXI5GfyIgJH+vRtQp0IVtNfT8aIV+rgTqtaGkIErFjTwd2a14Jm/GKJKWj+
QGAPHaNhC1DXcJoNzpvpEVhq4Rpant7UXawwxlJkB/o49+4PiEOZR/hjA4aHyaT9B7h8yfbaurfi
Yfre9yxMbdAmp7rjs00HkxXB0GaJ9RFd2S46P49cuSifc9oBIR6BlM9tgXGbVMb/yADs4xbJwFUQ
rxH1ZyIIOqZoKyTso56pALikYsQhoNkN5W6yiuNNx2Ski48Uk35G5hfR5v0y2QhkP6RZluh/rtvb
z9KySS24JaFZVnLf9NtZqW/WXjrhRzAnyXZvW+fOrgJUQB4xy/suKE/BYAfMWatELmzZx1BAMzc2
smu0966jUCrSIe++xPtm/xrWA13Z/L+B8puttVB1AwSgtkbFBoVVJsgHDjx+VwKr/UTEU2lW+ozy
wDw/ak3zCZ4soVmRPdhg8fqaj/2K2DGg7BGXBiEr2te8739/toW2pJ/ZeCL4hptqOw9uuwerLc17
nU9oMNrT8KGF18eLV7o8Tx9Zay50i45/dXcHNev5EJF1QsFQnqCuyi2cEL+QGiNJvSahoQ4CnH8+
6fN5cLLYUmrb9FS63NB8drMspCvsdF3dCEnPw1x0rNTyLgYiv7ZuWpYQIcOU0HfCZfAi5OLLghBJ
S3Flz1iTdtAC32ds7tqcOlepjibPp/PETU3eB6WZTLoGwKhTgoMSfrQ4cwVjzGdUaB8/cDham4n/
vv5WNwlfC1m4FuljNbvp8pVwJFA8KaH3H94dbp8Gmp6uiEDSA9kWULkHmufL9A1vYlsVqQiFIrjF
VxSaXed6IOKT8FoOtxLw8/063NTpnjFh6x4aT0fxvs4Y+AEyoen2mGrHjFv4BcLYYtmaC0S1Hvbd
uvWlPMH5pYJ6Rbyobt2hIVBcHD6jQTUcZc/X/3ZmRFx1z8OmUPG86KYBjKdMuk6td5pv7TWRBnK2
QavwN5FJjrTe/Ft3nArvMhYixrX1RfU5MZUcMpKSxE+/K3oMN7j7BH/jjhwi8REFOkWyP9HL5TLb
GwMg7AE85pDaSaZS+wWHl/txRKY6eTwZUGr6fAZClzH6F33pKYL8nzU0vPPabTCqn3oUkXLUsqls
A4te+jjgd3DFCZRIuLKT2+wW8c7h6PskT6T+3mS0Wx74Hm9pVose1ibHBY7awsZ/IoygcHrLW2wF
CFt8vHXTuWahQl3ozoKWsaak7ETarAiG8jd0p+k852vUHNQTgCJH+Um8Y2PXZ8fQlN/BPZqKHHzB
IrJHifougejhUL8O0lQ0wGqRoUIAWkLZTD8mpGSTab4NKza8TIj2zZ2m6CmR0IJTgdW2SU3P94JG
15sHXzBw4PuoN6DnE81ePEBFMSRc4NSF2CULxkYqEQ/Q/qM+stoQ4qjHantXwGf5+oMc1YlvbIdj
1IoSz9ZWWRRNrBNdPT30B5p4rqXL0NEIVHbXzTqDek6mBXbDqGasxdzAZDIdkz5Xftt5C3Yh8CKJ
WpEzCMAmQbj/RGTSlzaLR5TxkMpCJmSKk6nNuvtYXzuM55y5OA/KPeRc3rlZIV9DNr2JprwT+HXu
n8fHG7jT1tTUtyfxNCxfu8GjyOAQCK/jXi5OjwLKI1vP+3ERVkULGAoIHxv+DRNXFMHsjvTLJjJM
hjmGYJ3iy+Q4ZBnWkDaO+2Qf0n9s+IZ6BX2dv8f9XZjKNoZuwQQYIgcU2ttDcpT/iOGwSXdRGQNh
0leqJSpXuDowMt9mqpe9JbZgqV5B1GQofhOMWgrwjZ3Uut9BKy8UpJxoqkkjlbKgT9apf65TiAgF
MEUjHSeBCvCtijrvi39vqecktAi2ED1OvL5Od4JUhbcL6occ9bxBVlPsng7cf4y/e/WpDrxC87i8
wu6bClRd5p3wL4cXweXK+MWrKBmYOUBMKoOoSGQfguugLTB50EaTfUtwUUuwwLuuUiHCQ1CHSWf+
kwgiY2qqBBhmp5N3Nk7vibp/4zCwxkbof+1Yzj9fDS+vwFH6d9ud5cdbGcsiaS/qA2ZFvZYk6erG
a5x+rlBVCg2vCzK8Xet1eEv/sfqf33rnKCaIEexSf2AytXDzJooI3/jWqjT0XL43Tx6Gly25UdAK
PEHJRlwGiFMI21NZYW2boEJvOMplulN86Y8scTsyZF7FIE+Eu1BqO9bUr1JfwlvuB2c1iWHMxlGK
8VjbERWzzGEeLdVfA4gRM31rakBeCFs/0V3FL6pGUS3keIke6LV3UGl6xyT6irH8Hc47n7KKwBGR
Qfz9qw24Y3dHiD28Euyr9tedVo9vEmeiyJLcmZ3ESoFH5oe2LnVesktYYtVReE81B5WKtM1CVoOF
h7OisPDHQ2cSCMCN+1cwdUrIzuoXrUwidapTH3rbjNo4m0+bW5PI2ExyzSt29Y0GtxUShtkvzNF3
CMUt0Vl069vXBDhexdJPHVR5Mhf4pa9I0sc2rOT8aQvk4ETvA7AGIbt+XB40oXQaij25XY5VNC7g
E8CZDV7/DKyLO+SgWZO7CjtUjJyyNPGPjDevwbDjDpFLhEbio0ARNAveMUrouQpQWIh6whJej2yH
M3SBj/fXlqG3CSQ3EHtwnhwF5qz3wK/SZrRNwt+mc2Uj2YRquPLOQYjwvXHvRxFUwdt0xdJvBVLi
0BzdVNaZOJVGw06aoOglQ8C1D7Q8bdhMUvTyxQsuQoq1HwjW2BlApPxXYrhm6EUhTMZcb+U3c5sJ
DXmoJTZKRSXxvruESP+84L7V5C2owH/8OYCKG8LkBCqz0sMNTlyeFL/t6v98VswDITUEkqCtvS6n
B4bu3j2VMQrt3rII0MBoiovR6WVGFgZSszS1dWxkW7xUf7eBG+7zj0zgHH+/MwVU0QpvMz7frzZe
9EiTlwzHlZgNNqW3e6DsDfK6BMnqW/YYf4rzqSJogUhCtRhB3VI370/J3cMQwj3H0Uzo3OUAm6Or
JQaJfnhTavRYjs5O1s8mlqiDjXf4xJSAt0L8+pRuucbkW7ZrcgvNcijPxWJnMsozhyLrZncwyR+5
FqGDBVbrErvBQOMcWJVwo9CTEUs5nSwfNJo762/pwETVf0ZQBTcBkL4Vd0vPvLSlEm4vSDqLWeCu
YhWPyTGzx0BIZzPnncdF3mADYHPsCZPQ4biTWzKRG0HVcwxy4k2uYJVRoGFc9Sy8w0JsE04cQeQE
JFHMamR6+axetYoMtpR+EMO8RB4fp/jQyV7kOpmYvmev+xtdSsrMjCB7WCiSe2tLocM2Tc63iTLH
krEC1WJolovZiW5XdL++HqTzeB5X3T3CvA8VvJYckTG1ABiWuSUVFEs9p9GQ/l4d/t5eMOlDEj8E
l6e6HXYsnnNJw5eanEP4GQVRaT2vYahspyttQsc/i5cyW1cJnhzhG407kE34yNZ6NnOqOfa34Imm
G7veP8jqjAP4rhWTHWnvwQGlF30Eh2NfVpfLuLNj/cIGSViCiuO6rDjZ1nbuszMbyVv/gZ4p+1oG
ixGqtY6+sTl9zrmvFsn5vjypUX96UAiigLSoLPimKDZYd5xF0m5DCjH/bCyQChAdoDOVNZ2OIJXV
XfOAgPaG6SIPNEVDr8JrTm/I5LZRBYhxMP1CM/xIC8yPpun2A+EnGu0C/NMFF0OOl5l1YEGoFuMw
Iz8QO91E+zwDAeBwt+g6UMWNtWrL2/ik3Le1abo71G/guijLePIqwITQNUM8c2IdKA0fsg5fMFTL
jBv05uVftY1MQs8plivdRErlB1CCNwxd2MD2Y+GJQHfBXmyDOHN3+y9T3cny9Fe5N/SuxsgvIMh/
WTBdSRqkPtIBFvpgu7jtYZlXgtlaHDmhTet1c2I6Q8zq6SUnLHK53/tpvIsEMvSShZK1Esm/59gP
gma2qlSXMThqRv/nI687FtPZlVPnmrINJ/qtHx/fWHiZ19S2oUiq5I7Wj2FsqSOT1ZbpeX41BLD8
B3lzsppoqZgsUKtDR9kk8rbgfx7/ow9wlm0KmLy3yr3c5iyvtrSP6qM2fG8I4VRnRRu8tGt1z5VY
Fo/6cbqXommcco5I9PGzz0RfbLaZKLCMmScXN0A7wXjcZ18oDBQ1ZJOslbxIricBMlCxUe20magi
UQAi8CHQH4jpNuxH5IR0Hz3SuF4TP7OOylqRQ1K0HToxM3HOVqbB7L/dOaoJyvHau3aQdkaLsOG/
85TVOL+dIOha7erIJ3TSaQ53e1JGZxYULwRjYEk0xPQq+6Nj6S1p5YeUVx/j9/H5ijiilwpbnN2m
C/LHZQ9V535N6Cat1HF1X2UNcH3efzYg9jSJRQkoqAWf0MKACtTsyuSxZbOsr7BJFLsd6yNIBusB
h3bihxWDFT1hydpdtgnJme3FfAI29B/HiAZAFHlIT5VgdPfMfuCj5FK38o6OOfTGQGkr6bwSOUvI
zMYIlIRSPYmv3UqQVeRQrnd460jdFh3LRHSqc6Y0rxj9fxTheWcGV+hp7sS5EsutdIyz7m82n5zT
XFz2H+mV8ADHFvyCpueMLGPx+lKrxeQ9bGHUFBjDeDqe6lxqhvJM/K3G+qdJDiIGaaR+IMAbaz5u
AW4XYxmytMMjvECslbMNi75rG/tetydIOlTCMPYqYdborLGK6SAOh9dSjRxw+itbPo9Jsxi21LLx
te5lv9YpH/d6ujErhpNGwu0mCtNSuwWdIkUDuyyzYZiLlDkb8ecouw2QXceRcp+W4cR1LaGvTId8
d8JxJSZalwfc2Auv7ILU1z5WVFu2QBc+SmrIUY9YVRiNDlPPtxbJinARcfAetvSXiMwPM5Itio6r
5vJfYGgYgJmA/5BZlITEL8CG1JOe0Eu5r2tFle7PEQEuB7jecpmuVQwRG2PjCy2+E+nM1IlFTQgp
Jjm6OVNyj17OQY171ygLyjjDcFKAHlH7QxgfP3h3IARf5OwdpYCXkYspYuHaQvCqiQonEaL7qs2+
4x9/GKT+7Gt7CR6R5dq+wTEXuOzFV3YK6S1uiBeZps5qQ8vxYBH7oVTtznaMeuK0obD6IRI+/s7K
Utr1m19d4haT1tQQrBtvXmJ/6O2DkArDJ9oH8HthVZCsvulzI6MDMw055FWe/2H5C7I9Qc3Pl0Gc
CYi1BN502/gnEeIiesfINJucZ4BKo2qPt1hh4ffwJKE6CH42hmRS1JW0aD0+AHBiiifXSEgr6EUd
7HM0jLJxJ3cDli2VKudjNN47N6nqzYK6XDSheqikhRVk4wRmG+Ap4CD/8XsvsdRSXEYhA7zWGETO
hvChLuXPbcRtL5rRFq4K8nDKfblsXbkkNFMpumijPAxnTaaenVZ7do8//a0MaYfVqC59/aUj/Qst
wYhuN5w8az8KTh7thlZI+bwFfbczNIrTLNDVqTpCkN/RKUzeJN5Hk5fiD6nUml9CBjfd+cxOcbl3
uEb8cxRgFwXgufqse9jX23p87WbW+OBEARpwf85gZ2j65ftLDf+YC96pXaHp8s8fRYZOCVvnUh2D
57LPEt1o4m0VaSkulDwK1BtjnEfYAlBKYv1PiVq1pxI3jY76CA9wGoBGbtXCk7/+tTxrkmV8CfvF
ripmoC0SacxasoIaKffmxPNrUGdSMGqkAoaV4/ZzTUUFNUzWG2oJU7k/UfOYgm1m6Lw4E5xyJMid
s2yDdkbDKpdpkXQWFmGN0rYsFPjfVAjCMPHEMhAgxIVOSwArasipjMdAf7Cl6FBoLfc4xHKBgqVM
/KKwlVMRP5GWEeChXIEKUNdQPaB6ux4rrUVmEG61+lZCofcwLfCjywKVkCCANRi5Tflru2YZPJnk
VQKAq3IeyreTDZqT9NSMyUiOsZia5xi6cMkqRb0AasnYpsfN+E35+xOzbolZUIMHfYZZQYe4tj9o
nBbmusHX1UdLf8E1RXs3BGRLPvPWu22/6N5Ade7qjAlkaBv/ItCgaeRUkbl+Rme5lFF3sae0ruj3
wrnYbTIxxdonEi5XisusCcRai0O+GX5VZjRxW2lpZLyH37vZxJYQnYBT3mOs7gVyE1knK5IPgy1V
Gu4Mn+MNUBcAClsOvo3+/31dGqBgnNHytbavVLyS/wvu+f/iAWQedD/5EEadgvodMSgxtjFOWlFz
GcTMnkbGpswxQUFzoMmy1tiREMZ4OFiNOK1cfrBLMB+/aS4/OO4LZSS1gDLC4mZBh2Odt8lmkOZP
n03yZ/7fGBZhqMXJpkg9/yEDCUQEEj7AcJmEC7/dnJGFSiNaQT9Iu5jWWZ9SjtSzBEBiW+2/Qy2F
6xeY4oegPiAMBhn5DhkKpZArai27GI4jJH69vulOTycbN34dh6LdqwIvKIWAU7/e+6/GMtAnRk4S
C9jF9wzHu4d24B6EGUsmULM057jc0FtQ9hi4+vc9wUUN8zxqQ3iiP77usVuMZy4/qkNLmhvBAPYU
Ik+g+NSgQTxpXY0gdn523QymR2T65Lms0vZHHTQKh3/6l2DhNHPfL6jzZUXccipWvY74W1UqkQz2
ntplMq1GzeaUJzsyT24SjsD1vi6MTHrELgd/wfxABDmXOuwmhQ8IcJ+ONaqrBZSGor3TxSnKgQfz
PQ18ghaeyx6670T/x7baKYwJTKHRnEyxtGy5npbjd8h7jacoQEXomqvYBj04C4tGltUdrqenw4at
bZIs4oDHo9nAW/XBsHEDb2sH4FeCL7wXMq1W4It0f4R2DwNSLoHcQ6uHHCzhVbxrz385fPfUdJxS
FLUVP9VybznsfCBHTeNYYnGyIe2Vp1IEByZrjS3en9aT0NhZtnAmO/RSI9K0V5Qzl7N677M1rL0a
bV06WoAhT9JkTcQNNibu5mBJfYseiQ8zvXlvodSEtSBg4RgEEVujUR8IZEQtBsvU14DVwD1RGpbq
wyHwygxmjirxOQC271bEWcpz4FNfZbHPGiFj4IAbsL9PEh9AJTS8wZkoXmJHlTG8eN9BJIm4Ahvj
LwHeTG8BfxR4XwDpLkrwBN/2yPlJp/+vDaLxzI5rg4skxZC+mRGNWsglKNn+DyzOZpuB6y0/ZzYM
QTckW3WFDFqxXChGyDTUoAQLH9zLPaIQt3YNDOytBIuSnJsXZE81lah4+VKogd76imoG7+yrZV2n
9bZOYkq01+VPKKXv94I5Gdrn7yYA/ltSmmJjk1RIiOZj+xPlCEVUBmwRzuNUZIRZ+L5Ehhz8T3HR
lYYaOZY9UMh9BvUEW8PaWdp+j1uVb1cAifk4CAOqJP+YovKPvW9sZjNwo6WA2vd7B8m3es3kCCOX
4/nNGHp/VTavfNkjISG38KTXG8GcStKsIk2wC8bwkTnQ9pNP37rqFkp3DKZDhXU6cmWIVK++2lo2
Qubr5nj4ZWw9cpdzcWU72vNWaltfpw3t80MFFVyrNa+tOwkJkNc3fD1ftxjvE5GL03Wl1r7tUpYa
hZfBMcHRNJk9Dh6ymsHNPGRkaPgpQ/a/Etp95tYzqzj7gQVaGmHjn3eOo9rHCrlzlBwEVBEsM6EX
DSToPgi1gFwWpVgmm3qlokdbW+qv0E5lEC9uGEw9bVeAdYElyAQbLb0I3N8+KznQIbU/rKbTTerG
U5tO6Ust5kBiU5LB4TUaISlsxeVGAq+1xNtOwzuaof58V6hYmQy/jJRdFabN3xs/cFzOtjjJJBFN
ZhmJyw1kjzDW9+bXRI7v4UhR7rmErQV/xwLqiQNeOmqnmGp7TPwr2dVDNuGO1SFQZD3ZFvGgf0DJ
/2cuGxIs86oWVHoVZWtaowoyRGOQHgo6S7f2obCDdSfDTmwwS203I00vFOe6Dk1KYRGR4KaTdGrZ
11nKOWJ+XfYfJFbOyGugyzz41jplxJluDzukwqGxszukmQvfBLeK4jGEm4PLl4xPS65GC8A49yJ+
sJeBJw1bZ88HMOTeIF761sNnuD0Li1JkJeO0Lk2ugSrVeixPzxQULx2JG4NR9HRpbWb2ze2mrjkK
4pQyUQRLiMxYXgsrIaBP46aSNtUXmD/VdOvWVNiSfLEGuC75UcnLhNJC55W0MxwaQZW8SgYf5BLO
ZPzYXjN2BsWdVDp65cPArldrfWiAhdhmgPnzYAu2BDQQJhWtjM1KxR2EOdbeJYmSdzb1gQ+pUc2W
wG+wBcLOKwpppaHNg+IO7kmf7T/Ou9wABdXkE61YX91AmAYxrM4Ra5MJWICLMlYtTT/C2qDQr9r2
MvQ3KlkEkjJyXV11w/EMb79SzMkMOyNBeGTE83dHRIngjKwc2jmAJa9651yZrCl7m0hk3d2qFMpn
KlnUlgZS6qH2cYvoY7DD1qEe7yfAETi99FCsIdHUmI0qJ3RL4fbdZXP4NCdLttefGMDGq1UHWU9o
Fdu9uzGJPGCr4EShirLHNwoG4RiksH/Vxb0gcgAfbV8WVarqu2TtP3/JS54LwX6CU6rRJB/0kXf2
y9F7BCedBWVkniKo5KQ5im9Mw6E91FNgaEslmpXgl7vPKeSUtXzUGd7mlaTpTJ3hGLeF3u1DU+mI
tPJ6fciibLZcU/sXFLhGzlIy93D7a1wDYlZ7ADVv4gqFIVG8udyY16OmmE3tio5RKu3fkhBJZHrm
O+ijbxIjjerVQ/llvXKqoSkOrcpjHZE/AYypEMTH7yxEdaRyZcVmJ2kzQHkUx/jjhYdbD2PbwDZS
qm8NIyZ7Y3n46XKtrx0OFFb15rrKD6dTzPpqI9/4f+GtoOGTEvgMVxR830/p3++qGv7dSaEUvgp+
+yT8UVn1+OrZW2qHWrSpOVtJ57j/h0xav2vTVL+3I4JvL7ASRYJUqi/iX3ehvY7caVynnssiaFXq
RwT05AFZftJRTAahlGao/t8V1NW/tjretv9p7YlIYq8lrgpG1OozHbUkZcsqaYo7Ez79r3+n2h/4
0x/xShdcSwGFg+iNYZvM+eBnT5uKSZPy0sy0XtQwSwDr9SWLpeQHNXDBzMCst1vQssNU1Z+XoJ5G
NsM+IdTqkxlKYKBOeHn6R6j75woV15rkXJMbgb187a957detroZDV7KDqDSdQbiCvLV6YAFwbUc4
ZPjKgd4oXTmnzPhpj/XaVf0WuFo5obuNcE0MSLuYgbvmPFO2X9q4HccBlkm4xbN0m+EkGuzdWyb+
jDJLbEqdw0kM35t4ByYGk1EJuywrLmyNtt2PDCL9RW0FeK/Xsek3TnfcB2f+sEZRMZ2y8tD2EzeD
nRmHUctrEhbONKxk9Atu5AdxP7GJOuEftIt1G3MpS4r0MD9dAByui5EU16lAkn4uvaDXCboT/CZL
1keH5MR6yXYsjk5qOMVLvS7Uo/EeXgsyd30mEfM5k7hMKq13tLU1HySjkzuqvEhqudx1gVcoawDw
omUWuyRqvFItwT9gt5VMfWbXuRAh2gP6PSAh0y6CExSBnyM+C08Sfcmx2KFOLO4NCbylRzakewIe
2u/3HkAZJXbmI2ZlyVFHx7gLBPxovof/j8QIXU2I7Tvwf5+rLQwx6+osFcV4morhd4fgeGPwS/n1
lxtHFb77krF5cYKiYi1ip91nJITV/WoINNsjOwX2zHH33on3nzvQiTnLCnAS309wRw5WwMf9LyMq
c7AKU0NxnFNWdwlBvsoceVg73HGl9mS3QdDOL748WoZi9Inx+vbUHNw0v9T0qAGshqimJsWPGP1O
4nVe6VWhvY3V1HkWMBG9KDdDiw4sFSpibSXTfpgeAeeJgGYqYGAo/IehhIx7mgkQj3I6t4Q++NQK
8xaWRYacTgbzjkpG+0CngIws9JBFQqcfKh6/Fwz1rwSynHsVodutLbwcvpcYY+5UgawFQMp3NHCw
pmu1s8GQiXncB28SolRCNnU6UOWkQoGB3Ii8vl6eefJR5i6i9dBapbdVBrUuDbA9zHdoEz0iETPC
b4nEu6mhAaC0iYFWRx86FANHT7icQvuVUZi2gCNLKY/ndIIKZqlIn5JsvdTVgpJ85VHciahnblKP
IGg5te8C4Vf+Jw4xrWGVEejyhBYfA4n77kpXkaJEXy5uUlokiu5B/TJF41TSotVNTUTOJUTgLG7F
0jhEVLv0tszMIr9RTiLkfKzp3Bri3vF/giUJCw+lOFGR8VXgaIdUEU4SN1CT6FGNsnDlrYxYaMAv
C0amKOfm1UQzt0UNL/YR4qZHE2zjuU/LMA174upKibUd5xmMrW1cDJGIi+A5FymaPxtWNElPDg3a
xtHvLLL13JUlXF59BI01jEdeNgWIwS3seuCOBrkLC/NVvScrOKZZ2GnEILQHM4WrkbPtMUvbk0Dx
ici5K26w3meEnhtdnaLMbl2z+d4d/7eOpWMljiM6Cmj9phfYXYK7knP+qcqhKXXAJwReBqakN6lR
iokWpF19H7yEgli9Cu8GFKx5FZ5cO18pYstxdntZtd7SvYmFb7GZTTmNnqE9Vi61Rqit61YwtW2j
Xpcr+vCui22FsVZjCI4B37POIf/TEi2Is5PsC+WNmzBgXxZhE1xjouXbWF+Ud+p+lKgVsxH6Lcu4
vupUkqbzrVErgTq/SQCPJcDLYpFKH4K/ABrVDx4sZQCGTNJ6pB8R0bJ3oJvupsy3HLDP34K2Ifoe
IZlmZEvr/haNHw4XgrrP51dnqWx7fMGb7UCX9FLsu4uql/hD/chuHeyuJUV6RMK1sM081+FlHuiK
yhcW40SwGnbw8lBvykrNKiPuA/fuBD+LFS6ZfQF6bPI5FZo3qs/HJwrlQYahVydFZyxrHocI+c+z
Ss/4qyFW1gKvS9VCvlATn6yxzx4xm7w2NI5AwEOTWMz+7VF2n0GIedl3DAquHwxjBzwIYQ7+8CHe
nN2J+62JRi4rvcERwWtseoo+ltomYU84hib52XfWDtwGx4Be6sLRlsc2DiYYw/SEoQsId06MHgur
GDwFpP9mL1Vji6ZbKZyQ9o10glL+h0rYppnyJPcmt51BMeZAAh2GG6WQxrw7JPLwzDCLQS+8fael
yrKCQAaTrFJRLeoaHyCPb5MeQyKAlIuC056OHDiW7Nbi0UaXmGJsfJgs+cuI6Z/lMfIWoNH6tHi+
DS5MXo5qjpxSiXvk3yrwjfGFs5zQtSZYSWrnqleKiwlJaqCGVf7blD0a3eo95DhSTvR02XOXvN4D
ceuG/P60MAycfGvGIy8G1kJKsSOGXMIY6HeqQniseFTyVAAvEDuXpaIhAB+L2Nxj2gb8fYIprOHa
ITIxzsL1m3p9Ebo67jcgjjCjse7sN/zRBBrmUwtSY6TdZOzgr5zOk/Q+OUai+kxqn/rNM+mp/gEZ
mb1UiLl840BrTtcfSFqQx8oLyq5LXfqagPs2UHpWZ+FrUaMVD92j7xhcnb1I6gfrqEy3rhmA3jfN
e1s9EBNQ4qQv3jeFRv/p2U8xYtVzO4YagkQxx9tWK24FOSOqhPR/RFTuPXOzKzTFFh6VdRWBjUK+
pea5gu5I8aIQbgYKGIsfmZ2y95SXIeh4yqVPOJ5LmAvp0oEiDy44qMqwGWloCc4MXhZtLRiEKH4I
d3zV2l/xZKHtF6DlSvMJVtwCTh/hY1Z0el71vr7SjIl8OvakvGrrtZd8NyZT7u1+KvyMizNzCl3P
kLhXHoLrFYct/1p13Q6QJ1aS8qQH9NgNVaqmHYrWIKsH0vAIYbLifl1aZ0c7tzcpRCvHwG4yXjs1
VBdw7IFOrCUC4NoQVz2Suz2Qw9Igxhi06lX9uBYRolaazeStvWJEuZRJqhwDbAvoS4wix42xgsTj
c28PGQkgZA59VC/KhXGWSy4v3G0Tp1Sj5LeHgHLmnlbgzqUIIaopi3AeapYh6kZM4l5kvamo37L9
L92rujpmJDO/4WtBPehFk9LGl4pFYIIdreC7zERYzBaccgqrfyMFdpgjoYI8l8NX3+MBBToZed8h
0qP/mnbeHtE8gu6473keODGIEbvqpVni4ViaV/fJdoADilMcYvkdqvYHofpOq6Wz1diWXxW9Thu9
+PPmYFu+0xbakXa0dwpLNgU2dP6UlQUvOmBOVLmoFFrg+A87HpX6P+OLtCz2n/Xvb58B2sVZH2FS
pJgH7chNabZwNXTE/crc4Ff7qI3Wkq4tXgnPeg1RDNkEO/Sa+FBuoBmuOtfwHQv6Vz5Mqq3wRAsy
heujQ55z/YPwjdNDlksjbWlanJaqLX2yV3SLaQheynlqd9s1gt7pnzBZFPCM5GGD67ffXU8F64id
iV4agJ6BDZqOiqaPrEocIQtDFA6M5pgAv9tpxKGiRcn3cGVt00Vb6sR2+PhdNvMxkZSciirXTDa+
VQOdFVU3GdpeOy5bw8lwHrTC2JiSxeZ6t2sFJZ9ETu61tPFq8KsXjJ/KtlX8kI+yNFbtEgKsKQPR
YolAGD26iE++f6oaHk9KkHKpp2jf+Dk0cZJgdA9MhQbPsvMaRH/5YyaZuTYEyb04jbhK1B8gxq8z
QL2/GsNZH8fm6DSwEkjEXkV4PwC9YHmNENamLI26OxQY7NgB/jPggYdgHnDuFtZql5orh/E6tuhA
OvTmAiUNeZ4xHO/KrxBkARI/K6XxLKt+TTjDUikorQUk1pIVXtAZUNwytXDc5lg3k8mfh76Mqc2u
m0g/h5Sjf9lY4hrHSqYZGzrdJpz4jEhrBQV/U4I9e5kYjOF9HePZR17IXYFvOf+xEIHNIFZ+ODSM
KX5qnX4jGsvz0Uhuy/K/+/DDK6qKzHru8GrIeeaTNDkoNUSMKB3xzcNNGCzGUV36Yr+g4K1kysPV
2c8zYG4fbrwrgXciHiVsKpN91cBMncKcFWSBBylet1B9KwwsowkCxfNDubk1WE2vPENivZhwZ12/
YQdK61dew9ysJEjL4skHuIJx0AaG7OqsKsF7DzsNeDk/0kyH5UIBQIjFof6eN11WwkRGJ02rn7ro
tD11CKzyhk2mZrfnaM+n9a8yhF6j1dYsBUSaCYa4uDkPj5pEOzbqnCu1cSgxui71V3AOmu3FZdFE
e4GbpS3l7sijx+IuLUuEBKHx2XkZgRl2UMQvHHRV7YnSVLW7WMEozlPpGAqWvTffuCQMtHvw9jnP
mXBBsb8sN1Q+5DmUN5j8BF9Nou7Pwz3ewGZf1woYh/C9JRwXPiuHrRFXl5FBE3Eqn1tloKiNamKb
W9VxCKHvEKqlI1qISf7FG55AkmqmX0Osx2CeAcfa2S1XN06XwIJpwVuBqmQgdwlTh9ybYgK/6ZR4
vo7RNhsjtM65FFTussUqgoxukYdi0LRrzeYnRMKwMncE444XSg/eD+JeKBmnyIixy9Fzz2CP2UEG
yY1QehFtb0bm7iDJn11pDK13UX7aDWh583oDtoLeauO8zccxWCX1R8GQZR7HwPWVOjpczzuLo93n
npfVy4obyXyV+o7Q/Ar9MJHo3YsRkHKGP+GSXolo3Zi76vbaUgnkdkxtsittMt6TUqTjBOxNrhmz
S6YhJlwbM4WdyRHiVoACe388ypzcayjLWOQ7n3XcmooMtN8D7FDt1gmsNS3PTpLKvJspae14UWZZ
/n5TgUI4kkO982dmXP5rdBweRp/vTs6FCO1d980IFx2dmm5mG1oHKX6YSN6P1u+d9B+Zfl7msn+R
035l6tIB3bv1xtA/WLUxx/raeIRUvv34jRtn16tuU3v6r/JrWNGkt8ZHOhzwiqCKwsRj1MX/dLQI
fSbbl487Dkw+HIiAAds1NHK1duEjdLtS7Dno2RsJtDNB4jkaGKLI2Jw/Tty4C/Vg5jHZlXAozTOy
9744vHfIxGt2hNcYy0df5lPPDXeZKFVyZE4xholexOu0xjztBLG6P6z20IqY13MNv0xqAbHhi93v
wX+X2KvfAfAU18hGyfpjmDNROsAmdY2x6mORv5oy1mG9kgTXUScbNNl0IYBhaHTwURPKgNsBnc78
dO/d0oW+14tTy+W7q0bz8pLTHDn5qFEIuj1UiV4NnSBC1etB99PZd3LCtSBgPKEXmNCS5ut4K1l0
mvOBvvbQ9n4gu0sFv9LjTC0/L7ppRDWGJFsVBeELWQAENHRUr1ZxyivtpI5fUekqBHejRVWVMJZR
JOEbo9bc6+BYjloM6iLaiGOioIV2/luxmiPjEIZ4KRjssHoN3lzHhzqhKAAqwqOIOBtyrDK2F3+8
Tbu2tyZ411k8EANijYf7bvhoOASvvvnVM0dUjmU/OPF3abDsmi064oGfEOX0ozUn8EA6hsqPEuq3
ElY0UsqLZRdAVQ16ephIJjZ878VisbmS79cFM1vYM/1bqFaMBvY1X/N0hbL9R8S5uk48VDe19Cso
ipT2VbZl7ZcaLJBjfOyUCogRLPyoXtJhDHfFYM9BVq10JE16tQTnGcBs89hEQxILSF9dnkMXeaRd
+GAunmIJAE5c1zmavYLytdNZ9e9xCp5pxMu8C6MlZHGiyRAZgVp3uqiefXH2fMLppWLqAMVYnpbG
/SlpHJQITcw1lrf8JpMb0Mf4EFHk0E1BU7D5RP3VsVcsVKwDGS7Wci+JDc2+wYaJcvhi7pPuisue
deep8LwtAFd0t+18tjN8nSduZO2+6sMQYRj+NNXSDf9dEKeTGkVpGWV6Ab/B9WefhYGTjXStPtPN
SCTUaoeHhhRR+qM8/ibwrlZg5Ated2a47FzmsrDBui+K6XSJyLSO6HjbP1N4B9Xafv02W2SOEw23
0vJnf5JYeTb7wkWzx4ZX0nH9VAF2zsIgBrswo/QkctOq+rKAkX+A9KAnWQC0ytoJrZDadtakncNy
mtdglE1SdbIY9d042OBd6WFUNJTbKW0IIWyDqfkNaJ2tHmAHhm9bjpZxPLWpmHrnbsr/myYfsKqZ
ZbsC0hXDkRWHZLUbqXtODfN5WRpujVjX1JqLSSVNhXgqKX+c+wKesIlrZJ2NPJygxRnKST/CL2lx
NrGmNV3+FSd6NN0Xtk6dn2h72RRG6o9t+dmbdvNaVF+yqnXwZrmARnx56Ui/v52szKVIia/rTiFh
PU054LfGSwjgZ4zOKr6JJa+/Wh21TEipVGG7rNc8Mjjsjx4NREm16YuoloUrN+MrZkWGTgULiwdf
rdY0N7+pPvbmM0f7aOXH+v8VSh3x2kulKWXKNa/GqP7zpFGGCkt0RP9CgZW7OghrpEedWZU+1bBz
+zcuqsphgA0om0DmDCxu44gr3NiacyBlyMtr0v77AuNbpYQnm15yKAaKumviFEO2ZzPufBCPHScw
t6+9Q966UuOkp1O7AAzwdplYBb6ceIlmciPKjruRHc+LVlypHeogGMnprG+nTblV3xsxLKCCdaH7
0cx1zMwFr4IKD0u7DL2xU8gMlp946AsAr10f6yK7XBAKZysDym6mZDVF69fKSbiitWGw/weAeXme
Fe6eruskcdiwAqcak2aKAhvp/brueUyUgptmzcyMIPsW29FuHKaIyYOi7HY4rvL5Zfn4N6cQoOan
5HFpV/dka8Wb3N670BLmsf9Kbo3Lx4zKXlF6AaGg5d2te5kcfVEu3wo09/rX2Qed+2JG9eJvRCwJ
uv4azFe20ixBE7Q3B2QhrIFvrwhUQi/bDL+6sn1WLndUdo3bjebFfM24XlsJ/xHhHjJb65Rw0e/1
ThM/sPFYuF2VXhlIwo+ik2+56nvnA/2xBQVKfe17vhWXYTFWoFl5T2rh5Yt+B/lBDv7R/PV2HrXj
yVb1eb/2VicFEgxDC8vXYQRfaPkRKgahMc4e81rb0JDmiV9ggt/jxOxqOCFDXtjCXlYb2kQv5QE4
dzCg/kMKhwtO3c1TCNpHNkNwil+NGSaWRF0zmHReO5sDJyRwfQVvxiZX9mFMy1mCIJyGu9d5284m
nGWjZGW1fXCqRiYA7JSu5gPYK1I0okCupNiwr+tWQltEV1qaevh6abBwRR66l6GYaAlzg1EAJncF
Vuyq05wvVsUGDZDB2rrsaeb3f/1Ks7ANnTZKQMy+qGbFNtrKkE85Jjxvbn/KzT7hQ6jjsQjLN77I
8oQUnN1l591llm+Kg3bojrnL572frhBbjECVYB+9u7D/nMZdg5hThVd1KH47pSZk+LYzIcxhI1pg
bUMRGHLonnUI3fDZPT5BWS2cwIJppSpSej0lihGByAPUga9Z+6+8s0g5CohVClMX3ndeeaVbENyI
Jb9p1UvCCYOLjS575Q9fzLo4Ljbe3xq/PVzwbhIrpF7ck0LB1Nq2KyrVPk+S/2epB0dWDnG7Mkro
PPXK7Xi9kLVsRV2QWM46U0ek+dT5mzDPJa1P8TVgfNZevP1UaD7NitANRwego+6otxkf6L4JujRy
GTcPZhPplahsFRvWMQM4o+gZp7o5h2/QpnK1/bSGW06uZNAbbfZUmzgi2M06RpD4P3/nPD2OonKK
1dN498/a2RNNiWXKbYvDvGO1KxoeCasLc3Z5/cDoUpM6yqsqHc7BxgPYcQUOeZtCIwDpYqVDLQdt
5owgXpsRk7iUJZLbaNKjSpMl3PhZgO8t8EzXEP7RJWzgLKTrFpO48ULzQ9ZouvGIHtmkhijokR12
92tXoC+QgbhZFiiqDIZO2FrCSnmesBZsQPkmKLR/9dbwgOt73WsPwRJGuD21Ld6S9jv7pbc8EJ3/
w11OjUU7RbDsIg0RnCIJj5JKNeVfbzxxRFvXnzYbKiJ334rHVj9jy6y6eriwdANTdducTHArJpbN
40kRRL33BcOhHFK3SnMwt+CFkEY+6K0vzDR73AN9P3fQq5km5qOkFMJuSyVvb9EstCpbblyVcbVH
JXqxT3h4QVOthLW9W4S2A8ijiv8TlH1roIpZLYMIfd3MfujOZdZV9HHQskaJNPQY1KVfTR/wTFOQ
WElIHPgBjp5d5AUp7XUkF8QNrv5S3R0CoLHUqHcQf1ufcmF9qfeqhTpEU60+yQxJsJ9Z0Waa5g/U
sjrDyHBOJGRFZQt2dTJIGYUougenruzcOC/ciaMOQkVjBzzWEHMriPBoBSdRXAk7LAQ+x+mvayro
zMAieuCCHgjhEceyVVFn2tWZjWH2B5yKjvjwYHVru1HOd+5LTrPTUmE14nJbwVMwbyQTHzpo65/2
8Ii30GGrBpbokOpta7z3FGdKKWN/vCe4cQR3CntKZ5LmxGKij6qeUFq7mrtnOZ0/bHNo+s9inYOJ
YSaNDZ25p/vXS31dQy0pACZOLNqLRszzD8rakg9S0jL35oGggPQUNCokPCdkMF6VumfZV0mdWt5L
MD7NRdJ6DizkRJZctrVobkREtob1G5w8DJ43kA0q7sxppDK0F87Q+P7jMgygZzemoKaIFO0adFWV
3XX41Jh2c16ONAfgiega/P/BjepUYxpoQQ5CYczh9Eg8qUqoOVLS6ZMmGVxQx4Vfsc0DwW80MqrA
Of+StIFUbQHuMwgmYaeZG5eEyT4nyya+o+fljB7S9m9BEJr8joI6UzKmDyQjxeZIY4JgsrevDf/s
QA1GEIC430iP7zodoPCTxKgK0nplvKykcUtbACK0AtsQJc9xc07StZlexx8ZHuv09VTYUHsSh3hk
UUtqzjVQbILHvXukWZhZxHcso2zMLlupMPVcxZ6RbJvnsbAR1tkGTxOIwTm0xq/NYFiQXHvjSrwC
39oELBe9wuvmoES0ILXsTvGFVtOw1TKbBP9dQ8jN2Eu5GmSygNnHyXGGqtj35Z/I9R/5/AckOBoM
RSP/Xe6FzFkBaOnBYrzKsmSFvXFVZLOTrObNpqqtDs6W0tpfEy1cKEScvaJoqFNjQMGujlOcIUbJ
tGgx2DtMBybdgaFVxT28On9nK4sS0NKrIQjIwjYgo7Ui8nTU7Z9R7O9rjD5LfkHMlkt8hJcOmbjS
ObjHcgrNqwyHLiOeM07LXsnUGqvj7Mg7A0/BSXebH6bIoIjoncE0JYPDt8Fb0KI09Y5ThBnG42EI
h0QQPWy3hE1ohCWANrSVamMxxbEvYqrJ4PnFnTwmg4QDpkKkOgSIW6DkLPK4TQiEq76Jthha+i3z
CeALAG2XeBFYvVWYaLTj9vxsS4nTFgbec6M1okoK8tLD+PXQiimIQHqQUpEeEDHLg9h4Vk74RIfY
Ahv6Eo0pDhT5nHrjd3GAvLk4lHwRl3n3SuNs/N/EmUNIcExeIqpshi+LfmxxmYKJUsxfiHpHeIeG
Hmf305znCsvOKx3PQExO9sOb7jiibRGB/rZv/HUROjuNFTk4A0NjveQ7l+cY6SbYimq59hHIg+oG
R7xrpwrPRxyeKy69bRIJGc/30IqSMwv6riGBkDoTXtmEGYHLSyuge09mmLBDD1UHqIRfSZ8NxWFK
Ff7LU7zJeRAaf/d8YJdLC/spQP7mYa13lqIm75qitihC6oduYqpx7gcqU44Oc2kUUVhVW0eTN+Se
53jtGPgWl0AwP7LPcp+F42t38d1As7UECYvmfvPZKY85ZmjdC/YEVNOoKC7i0YB+XpaAKRLVP9gk
qCCUYnbMpLi4E5mpmxRE2M5D5uu1nMjYN+WxkM09Nu6kdI0ZpkAA6Tkm+WvvaavL5cXVlIFdcsWk
VJIyDcUmVSvIdyLR30I+1TY0hjjeiZea50vDrFUoRIMGqYmjvxdq0xLnKTpv0SN6AsD4KPAiXmCY
8oi2Xh0Gt85F5yBrKpJb+uGuYrCYECR52xyNQMQBuNEjBdQGNuO7ga0wQ3isc/e9pg6euavF53k+
fn4UgJmGeLwOueTBOaj3/Y0Nr1P6HIqy2dScv+QBldcxI3VSCRGgaxfxj59xU5/U5Ld5LD/KNiJf
ZccKcNBIWnn1zmDkLK3YBxvQBGi3BECM90uqyYVPbmx19/Ux0NwFMeP7TW54JGsjXv6uo+xCDwsP
/kYprQqqbZ+y1ltae/Qb99OBB0cg7sBBMtNOMf1Y3ZZ+h7rqDmavA7VXtQ0Km93lP7J/S5ozKjmq
LjNTS4YuGaw0l0HKEIUO5L6YS/Hc19E5K/8olJFbSZtTmovwzurs+4Z1AjLriWr1l/B59+gtnAAk
7IlIFQiFdS/sOAWUdpSUGa2tXEu2UNztQXQw0e/B1FLRUrj7tzhapv2J5i10oYyfWOogj26quw+Z
KNf5bqLWhNFtHi0y9why8PCoP5k2+orWbsuUaSpqSj91YHwOUS2sHJKP8nuOhKNO4PpbrJS12xo3
r+NpxpoAf+6qXBu4AYZCtU2fTereRAL2PRMR1NtnhhFnoeGTL2qjGQ2J6lJhXf+DREqvQx59Pjcr
BBc90qKvDhWQNwSU4t1epki255VmDq11mDjt7x9oAJHlp8YxXtWwi2bW1qFeWmyt6DSGbGCu1y1Z
CgEc1fDE9q9nM7oMi7wFMz6WlvEbXYiablIgRzWuVYhoLhcb4Yh3vZl+yvf4NrcEWKbxSPCARacW
UUCCb46iClOFHbLxsRudpAE5+Oi9Fmu6cJZ3j7j2gpkSLTwPQ1CxvaH+JUYmqAKLksbv/adU4sXB
udomqXzyLtQG4A5ibAKUsqOyKcNsUVPMfxJyt184R+xVhDbrD//bgnuy+Cq2UU6zjrT8iDW4+3jS
93ZdfCytv14gv/ctYtvxDtyYmwChsl5EOOX5WJqlDStJagwPA3rg1cE5rdBhJE3p0XfboSH+uaz4
DQ/bdk49hiTACGReY0GQ1EmpekJDmG1R2PRIVY5iIopWlYkDpICkld0UqGDVQ3KWLRL7q34SmKha
V76/BvNGDd/c2ugLiG06orQS9gMzAAGrubcoxJiNQy9Ikffp8ZKmMlW0kj4y6oTHGL3hfVEpApZV
9lnJXKQhGcXKxgrBcW0oh978gyUIuignxLNj2Ux9LQuLoG8vQXHNZ1CUYRAAm1DAFuZ7BanweOZr
q9L+EeIOm76Zmd3WB+jLGnJZfBIUNglsVeZILPctcWuywf8acclhdeoL/8Buow8v7Id6u0KERjoM
0RhofA7MCW/Sl+KSwqMnTYkKKJFz3xtdy8I8ixib9BVYKfc0siauD99sovt1OQ5zUQdL+RyZqcab
0X/l+gmFWpbPum5McIzekpxbwLxqCCGWHETVOvjtd7703ZGP05RRzj+pP7xna5PTCG9r21SEa0Xy
ZSygUa0WOoadxkb4jQqylAjm5Oej+np0artGToxMW+0wZ8HsP5Y+IEOhEcKyey3WIumqywHZHgyi
8VIw66WXUb9idfx5MEyKnWEb+nvSj9N36J0Sf6FSJ+9gvlBsOAWxM/ZitQ9+Av8IviT0RHtuOXUt
hs3c2B65R4eOPckae2BQnMNqfMIxyoZqSrcpJwt2GnGA0qbzE3wIfTivuV7njQVEVc2BatSsnTAL
CSraNWz1n1AyI1hDl6tdrQ8RpLwDdMss4sb0pGkOqN1NlKiFCW9IdyHJk8H3zVoDVxM9rZIOZ09v
njD5lwW9kcvhIjOXL0Qd1hbfftF0hQlMhmU7lJiLGFoWvc5zK9xM5c1OQdYrn7M8ZhqRQZpolUF0
ckoSHdLuPnSFHDac39kw08XNPiHe+0KkJQXpdXWW6yBYlDabdqocTIw2ukNvsvXkC4PBJkjlBSB5
PHslgXPphFNHL8ne7apNtUCloLy9Gx8ZGvfF+SOHPWjCFOP2C68EIVA6u2SW4WS8IXajylgu4OPy
Xl4Id48BJgqmGvoayse+fjNIMFqburehqzl0OKZ3ZX/JdWIWrlxdlw0SF3VaMAHxKPSyzSvX21Du
RsOv4b+FrVPc9cvaM4myh2eMVtngqShUscpzUbDt5wFJAZD2vkOifjf22RDq34+nonHqYHt6DQbv
Q2TzKL+l99DnGQuVZxdVu3xBhj7dfhwXX+kRLqaFX65SC3h9IUB4RiZ4HLZaFVop6NetQkMbqH6l
SRVluh8D9XI5m/uEHUH/Rz1KzrRZ+jlEOAy98dPXnXRCszkz3g+mvS6/1qCKEH0qqI4lLEVQmkwM
SCNdoRiavUXuKoItpiWFJrHCArkhVwef+7raeuErKu8SvlzbvGyR6BVMFarK3ZZmlAgtHnJxZzei
OojQ09OQT8ZJsPHrfNJeqw6m1J60ms4HI+ngKr5DVbpaFNHfrxSpgLj8jYmTSOkBpbuWAZukD4BI
UU7TYPHzgTMVQLGCZ8IG6Pls+OtQbN6pNOBQZUZIVLreSiM42ByxpZTTdtRX82yDTcYj7hmGPnKr
PfNzpUejMnA2mOlWTqvTAtYHt3ScBbFfdsDKSAdb2EG1Ks5Zpg3/AKRd2QXIJ8Er2H+r74R9DpId
w9SQ4pRumIRNZ9b5rMecJ30RlP/8isD0jsLaR41zV0Z6YcymYCwZXFqdM4w7cdIi+4/pSDy1FA4t
dBwerj40k6vG9++esRgexvs0+180N84/WWuOu1rb/T78stSP4d8O6kVeEOwy9ulIy3x0pwXMh9ml
AYeXKpm2OIodZWJdlKbX1p4mzbNTZwFXsTVlb0Xlug/frYk0ErHrwY4VHqLv1Kgt2b3i7K2v7+OE
v6lCWAeVrLdQkU4hTklpRXN4IV8Y9VF9/JYFudXYvtdGthPwdJq4gvNjTktILDibwbHk+T9wcS9p
o2NqPAmO5jv0Uc67qJYA5L4vajYtSgyv3PgwCEtCVI0h41zDumzvfzAJt+Hk39ZElJ4gdGM7HNv/
e9SlkAEowfxbPxABJO/vqtB+k/BjIh6VlvF/dhIPzys5ncyyNpSw5hNlcpnh/5X1krwyt6Rn/6HJ
qmn3WnY5v/ZlLy1FWaRx/hV+qGHj3xOLxrVw9gvEQ4dC4ODf13DCO+64d5AWKQcP3c4XKx9UNGkb
0x9V3V4WpfIuI5feO5IcN42Jr3sJlU81NLfvh9VQi8KiJ5bkzXOpki1p4ynJ5/Wa1t2cjaYX4+St
8Fqi5sTdAqTK/y/oPEL796/Nw9enF+f9VUVtPHRfrfY6MF29cd1UUsjsXqHG0bcmnVqsLYIp0LGf
E3DrJyiwewMEk1iSjpCncujvpqL5WZsZZumd2jLQvS38XTwOrJN+7D7OlJybSAnwvdFpZnFtI5OB
Xq3R6Tax6RlrXu2bCxLqoSvh4OYIwUkrTEfEPce+yIpI/fT9z51+ylvj4quM8/8lRn80MSeWYvhA
a0toOtssfkJl7L37VSHM5YB8Z8Z6fP/7JAsLlz3I4Aj9pricLNOSnyJXyKfKkymDv5JYG/RHUkct
cuNJ2epki/vKtTLmbagwF8AodhrrzjBwTrbbh0fd6JBLfMpG9IOST1WS5mDS37DN+IHJwwRIoTdF
MiNSej5b4KlRaizAC81hgrKtE0WAz5gitArg7JXJeVpRdGtbF+Bwi9lHre1OZBxeJK1mjip3uuGF
mwQq+lMQSndfBIuM0QQwYal8R9vn/BOQe/u2yYR7x7aJHCZFbZMe6/bj0+ZFzzTTaZ0YQzCL7bUp
h7Ck8Nood1KhoU3ZaxLqpSmvetcDxHOTJ1crORnDsHLkGnv5o1a2vuGCGEHUKqkYHjdmWj8wxZX8
5y0qaeUgDq58MZLWuH9Uo2rIJc7hUKQ0aDNywK04rV3vIXgXZNXDo3q9e+P2U5PEJ+gBbt4Xt4dW
cFjdGjHcPKvrlGZG94EB8fOPFs+5h5uhJvrth207z8VnSn0O/F9LYptjdM4Vm7J7IAq3Ka972ed4
XacLiFCpQQGveteyAEnub7cwn+Jm1eyF24AW454xCN2PUGQ/LyzoawqCiWV3L/whMAlW/ndMY+kd
FJyBr0TfOPux1bPLzeQax+vaip2BnppmbmqYMahEtdRa8tSjzPbi8xrzmdyLZ8LMhN5pD1GfPmHm
fD1GN1Jooi/i09WkEWeoJZ1ypl7hMfpSfEbd6FSODnFIZkJ4pPUE/nHKXCglj3agoLhzisdOFOzT
S+Pp4EC0gFlkUbvjB2J648l2KgPwH746JdG3XBdN8hYZb11n+LhirK0NUE26P7wSAZxqzsNMOZVj
TH1Kyi5jVviXNgrhLVDuB42tU7NzpKMLYRfiS4OS+im/GbaXTNRpgH8Y9xgNIyvxluasOO7aiICk
O5CvsQCzjvU+ourIgXN3luCIG7lKpYGn4Bw9O7B850tRNrB1lgQYc91m8b228Jg9bpZtyvWai2jZ
XXsuMOD82qA5ZoSWHhaRHfm7mrKx6dwyNtRoyM5e8DUyhiO3GqZbt9eoEn/lFRaHck3bnOexHuVg
7svJ/TDPXiXZPYlkeEDAogTHoofJa+dafblu9NrxDe3vX4eCHaVVSDD+9OS7vzsrFycRMrYws6Ld
Vi8CCOAJ76IPCJ2JYWvlxcHWCeKUH/UhOv8T+h1/0I+BpXxU2MhoMI6vPvK94/dVYJBI72SpDVCS
HMUAsfnQdmTfFXtRSbUbeyRQlod/2AWOHs8awXN3XD+heqkIYdd9gIde+b/zIMImYgfaCRlbvS13
6U5I7SRmDEa1rmK7hjqhb/t2MFsz0dvq9HM/PT/QZZRSigYWHHDhvnQdbi5/i41U1S32UyZ9G4WF
I6Ey6yeifXADvaFs4AgWu9kANED8MFcFpEBCwxTmPGHdV9yMUA/D6TJ3pe+FP1WBtXkIPqTOo/14
GyiTzxLyC80gecmLMaek9pcTvWRMSHR9HhKyKTKC7xN1fBwDOXH8a+QQGqAiTG/X5+TDc7Hu8k4j
eaejyW6tsh3R/tl1uvwnPqxA5eCHmh6qPKvOe4S0O0OqN1jq+FqtxittFo95rIIeDauITZs93dHN
49qO2Os6rhNbZzEKnN5tu+5NdTVsoLGemGEEoOBCT4ZiV9TwkRdJURdkqJ7iNgm8XRR/hCwi/4Xh
CbenaFq1NUl6QaG+DLyslHP47sHV1YiSRLqZ1l7tizW60v0gYSFzC/YDAbXS+PtvOdKDLp5aewiF
t8r/6WJL/naBbmpt7+Zr8xJpWBuSUwDGoXllDr0Xv9cDzt+kofb7/JlOxkGNol9rXdSoCQII8eEi
oSrhPwqa/VL509j5ktmB9DrZnpL93LLV4phSlw2P4nWJrfkke9FxCmWG870s+uBODIo4TVsRKP+4
U61V68IAsCyPLoyd3QwyhWBIeek3wsQpPYmVcrcgN3+2TO9prAwG0+SyelVykoXT3IYsezZlBJIM
ir9pbW5hDa9tLr5+bsemsaObHgBHJ7NSVvTNi34XHRWHy9iVSLF2TWcqWlLQcuqivmaiYlZ4m54x
DYnbkZHFdUcN77ZvhXYTHN3klM0YogO8ie02kpYf11ezvVFwTw1xn/aCk+4k2LfmUWj8ZPZQgALr
REiIl6F5qUyfC0mkxBW925kyt0acHGF3pIlpJ5W5MNkyxo9gP5uexcb/N1hhWlAZWAkckjD8HlSE
PUgaCJLhcHsnM6eThQPoGfOacrKcftTOiSCz1C4a/Po1hAecTvrbOxWl5VAyNMkc/IDhf9az4XNR
X+gUeuKrOXCJaQVjgyquzK3PIW2eNfklJ8bQqLN+bQ1AeN7KYmQ9zfw4/QoVk2EF0CXATlWQ6s27
gBKxLB290FTVIAX2iJKWzNc6x4yIihVMpUIhY/NXp2A0C8q6KbdyN6fXvj4R8Tnw7tj16o7sH+QY
UvYDqJ+Dq/hLLNhylnWlIbvhN+equL41L0cRaZHP6u2Weq46Oy0KcqC1DChLIKRX5zEv1rBpOnbd
atLRblTyRVUgy80sbEvPfNFcdCOlDXY6nUVjivgJ9/d3W19GABNZCQkyuwIPCioA/h9ecasAc56K
kqXUukK9x+o3t03znFh3ejat/Hm9IK1Ay1QW9Ti2maApaaNroTjPykLKL7hjEBq0GGUbDDwDg/e+
PJC+hL0T1qnvfwCvg7F7WFa+mD4A8jZ9GULLbL6UaqBWr948z728hH+LQbRDtd4QHgJl/0QFOJ01
Nka5mzn+DySC3EKB68zrAFiD/e7yfkWOqdLGCBF7U6+LQyBl7t4idjrXOSHDGFoMkWryARybtVZt
/90ai0Q8lj6H3UkwX+qh3Nebm2tT7ZigCwAA2KS5xNsW2Uk3NO6uy9Nf2MVEWQ5u8T9FwD+15npk
/n9EZTwLE12cHZUZXf8hP4BPKhGzsIFz5pcGEV+1r7LwlShqFPbvnJZ12Mi9ygK2REkSvkI/QgqY
HxYa2rFvScKWouhJf8RkJB8PyABv0v20cTMegk5IlKTE1ZpFkKGUk8x0aVXi7uQjHo2QvOeF/VOI
RM0PpCIN4RKUfY1iP3jqdfOAgcz8vDRkdhD0KbwBsr1L1UMW4aAYRPo7jet1fcYWradz5Tzsud1C
/a2EiFr1P8q6UH+Pf/QM1qHiEw8Em8HaKv124/VU0wgeUaO2inpEPzbK53ObyRWmYIWykhS/xdc/
ikxikSwtfLnydvFAFxtG1sVXBQhIjmkBp9hwoSMwH49yq24VHVQpP/uoKpltHDr7bd0/CuPl92Lv
3Lrmpy6trNObQCOhBN6sk7k592cZNnAxo8DeCskrR7VvpDyzJW/X9KS7Z+me+FeOvbK2KE8MdZHG
2k6krs3lfGNkGM5S5iKQ52b2ZbYlx5vTszdMxwxsGUrqo8ZtkJZ7QgYyvzYj6DzaOpJ3afjRlB4x
VV4orEpqwDfBP36nrwn/o5iVWmjJzuX5f8NSWy0gjy9lXP4obOv00ZMQo76pEqulM1ljCeHrUkSl
QtsnYbzu2l2CASQ9SMH8kgCv5+1DBkqderx96wUL40+Jne+6cHt+3GVmPmzWvqscDEGxNQNfbU5k
lfYXIYbX/MJ49CpS8VW+gEzOyC18s2VIcRQCcLSQG0El2HgYTvn/v85EAfGoSuBTlOMmIUw/1oRP
IwDIpeacIODbKUgEZVsddlGeW7v2/cMe2osAOI2RxPHhutShlhND4kVGBcocaudY0kKdsxGL+4Tz
ptYjNzEZ3i0gFykoeqtw7R0dQ3Xn0E0kwU3NQm5N5L3+OK2oyunl/MZpUDaDCz1r0deofgwV0gAI
/KEqFgb6wRzJkapr1pKr3e+KGYyed28PgL7kdnrro8VsN5L4rNLPNAFnJsNv0UP4sURZCENAJ4DN
fbapg3hOGEiG0m/pou0LbTD1PgRR+dqWkJWvKZSyVMjrA0i/YVClHTKOAwrgZpHCr/vFbatBZAS8
cJJAx6oYJbeTg7iqZJ3kHeAMzfMwr+3DDi+8nSufBTLmikvEbsvKabYiyzd6XGmnyEm17VgWsUDk
OPn4j+0L1bpSiZ7At5CZ6qgh/i/zv5jfGheenY8BlDB9ECfMZj8KkJBzSyt2HbBUNvN/c58zAiE5
r40AZnvEULkETm1wgAtAdJVETg65VXUAbI1iIxOlDvAdF6ca/8fOQRVz65HmtMEUPxLexhNvH6gd
QL+iSv2ep3sjkhJYfeXvnUHqMVQs4VMbBB28Hlvwk4XfAxFAlA/UGqON1fgan5O1Bd/uDXChYne5
lvc5L+g7vce69szHHqgor6SDq0lyM0ZOF9hdmGzvzXUh6p1YUzfpOxxRPwKr074fFHbY55zud148
dciTA0Q/r6WtG5D5Ktdh9olOOA074IfoIjCKIQFlrgyCFBLJ1+ozkbSpag8XO8tBAfScYsupXHRK
+R6yJXzlZI3PBJDEiNUmBrySoBHwKdPqIT1wMIqcyGPN1mqSscIbVUvO+/k4qWdumvGUIvBzOfwM
EuEjqwwv4Go4hLNlE7wHiBhmfWa9XdjgMsBLGRK8V3DZumwswFl3geOhDStsqm08tHj87nifEdKS
JNa+8GaMbPLOaTp4d1Fik2+DHr08b1qpRVZPVZUR1Pi5mRRgAckd8vPwIeEr0cVI3xKowRESW/uD
oBE1xrZ/P5JhAaCYKt5SFDJFnJAxKp5n7RsgTO1DQC2qFtGYnpuY/aoBeGqVL1L30OKf8UsM+Shh
7AIUjjbNtj8w3xzu2NE+qVNLbdOW0m34meBargQZFMC3fCyDpyJa87hgQkuuA8C8JUH/GRZHDgUD
zsiHNIHzryenves80OpGgM+UqdjNUQSlzYOWUxZWXl+uCGUkC8BihR4bp7uDpckcWl0yBCUU14zr
pp/l5yruB6eiKs9tcj8gbxP4mfiWrJ1Ao3LWNGrxRWvV9yAfNAw5+ShqyH785RbQB/ElUjN8fq2Q
pU1vCqMtKrxBHoI3s3bW8hzmPmOkuKnqHzUpF9llPpQ42tuYquHTRJPSLppmxPOyfifVXlQRpWNF
K7/ItveMLG9n5sBbIpr0LS9SoPDzUnH+1JgEqiEk9DAbaR35UoKnwXCcIVkzawSUSZRPXj6hTJsC
R7idxW7ebC05dtM0uO+bd55ZfxgTQXXNJI2EFd8Kw5Uf1LdKGcIRHrTzCX9w9K+U2a3Ruov+17GK
Hnc4XoYDXs/+OZTT8MKlHqrlPeTF9LwmZBGaB9HNOEnNOPJ0ieUIgyFnsK8WPFFgbZ5gVW25Melw
N6ZON+yyLM5fuyQtbL+75WUCJ21kcVJKVcbD11CjG9MPldCa/YbjqlZSLfRz3kc8XCoQJoaKdqzI
gFDEDwx2zuFCG+tgRknrStw48/f8XrusLQuqubq0KBQ1X5gOlnOFNNCQdVInYuwey8YCvaEZp4rb
6plxRD5ASbIAYjJjVuzrct5l0T7xM/XpdfksA2WGz80lkX1A+75lCyyz67Slbjyem9saCddzORbj
FDa2tcM1Zk5hEZh6GfOOqukmHSznyT0n9h3hdyWiOLyow/XdynfNQaM0WPSUIvPB7OV3iulOFKgH
MtB9XLI3bpTH03VIWhKXyagPPtqmd4pbNrSQgas1UNe+oMdwOi55yHVSb4ZJlWXfOJDGWVVeW4LW
p20HQtwmDGBmc4d45G53gD9We8+snvUOCGY93kgNuhhrXCblD/rEi/mtxWrzCURcmzY9q/zwBg+K
7hzY4K+P1DS6pEnnvv4b/jni3VFlEedKP0mjTjRD7oc390XSJoFM99StjoAT/YhPMUasaiReSan3
lnMYmqLDbhTewovRdAYX9gtvHFaljsvDabxmSfe2Fi1TefInIUmvGDfQBFxAw/OUFs5Rgc/cC5Ac
/bo5ujBcye85eu+xhpxRADR89CscRHmbSgACg9xSs9TaiByEHi1hQdpnjSd9tO2zjXrSfmSb8fyq
lghLxXeXrF2xsDuKYM/anJNKNMvdhfmTN78Hpqi38LvHSudRTPdzYnOxvvKj5kLmh3ivT06fJFnv
KOBvv0Y6EjLY3yK7t9HahSCfKWSTBPDcsbYmK8Q87In68O7seZRdgV5vwT0Jjy+sCv3GImhCgiS0
7spX2re7SfyLQvShuinxsYmbXrT6Gk30ZVvYolWq7kngGRxP1QsvuCUG4ZB4d7HS6M2y+Wbiocut
agTAGEXGRk/aNbnrMOhcibPmmTSjTY4mffQ6cubSydcUxt/8sBb/VTEHzkf+2wiXr53ExlL9KHJ3
PgZ1TXhPjgH1FTIZnsrqQ3abZVdkjIlj2CAOEJwf+uak0UKQvZ5cBegWljKSCxFUbooL1fcTOm9W
WPa1qE+43rrHmV9qF3/kqIbFyjyzjIrKYGamrML2A/PlNtXqasjp3TaKK0GXqszHJFd+w+1diW83
Bbtk5wR9GOQ1PTCQW08oB/nAw7zN+2EvKxTC6eXpG6K/mLyNpIpAoNsXSnU0tgme+ZgXStT15AWX
LHi3nLY+eF6Q44wLpg/QEYJ8eoIIpYoUtJKvn4HdF5+GgXCqqV6ONVmJ8Vk926pn/yYAEm4W5Gh4
YVyBVgj/ykd0vjQu1fkkxV8PfQ+9wOHDxgEXKxBcaUS7EfnjyI8V8up2ZYgKlxRG5t79/eWuRfzC
yt/ZBk1MlWn6G/X3OTliKImq3nThbJFgdXj/CcvM6vzO9NB8eE5xEFjUJqxUOspV4/TaDx0ntv/r
CSozRg42qgUVC4F90Lm7+CKBByQC7vmQF91Kz08eShk9FLMIj77cg+sIFxo6el5nNO4Ule4iNJZr
TgO1duZMTftndvmKGczLeWEeZvr1wibtWtPQquEkhndcpzLB4gFWQKdiZTcvcHcJmWijtiFuXcWL
rBYCmTKTyzXv9Ppc5R7U8qKiB1WPBgltEgl78KrJ69TR+MiAZEBaeL+gOy9zcxQ/tVtN8aKUgfrC
Ks5BrxqcM3rFcS+DGDR/kwvh5xTAtZ4V6erw3DRUguNGo3wAizw+O5GNyNnhkd8GVvKMxyhC5BbL
OHYOOc3HExSeiqxvm19+Q1UgPXH0JHCw/nawT6vglxFbrySfK7pIA8y/HpiUuiDbavacvm2yMUFe
E3TjPQIC03h/A3EgAnlkp5Tz+Jp//Z1IB2E/WGkzHNNl8QVMpUJiPPe6NZTALw3goMxEZ0lMYJxD
ZKcfuIcbMG5jrQ1upEructamspbtY589agJzUIERBJd+bIn4RgWPSD/RcRpLwOX3LqCigCaAk95G
EAl5c+r/h7tFC6wYqog6OsVskcTex25pUFealZtc1nrh5dw5C0NUbj203wHKjyeLtaV8FV4or2VA
auqTIuf1H9yN3pr2lNjjmy1QQZmUeBIY6bFhckGMMVoLKPNmwGG0zE47hHXEiS2Kxv4VdGZ2UlWQ
pBSA3fZpSoKp+KQT6ICcUH0Ie+xzY8q7wzfUG8uhORt/eMwLgVug3ai0+Nf0Flea9l/bpsR7yDa5
8JwlZiNApOxXU0g7Iz3yN8hmtJr4GMpnshdxFHOPtkVti+1Os2CxIV6KegYyuzuggrzWbgR0QuX3
4OI3jemdHzbFSLdBickyeT8VO2k0zFjixW3fQ/WWSlLfa8lKqFYkZHAAbkbpNd6slchHh/RhirjR
vZnT03MuqNrpqbFhnemGXCdbArDY57MnaQnXgiV+3sarCBfP93gM3oCvhUSyD/vxm3hxNINtart9
y4C63/HTLAhDCg7Zy4+/Hd8Wc+vhHmqueLGIddNnSIjKSyuAfEZcScE5ab6lVSWf1PJ6BRNe4KNz
O2chGMAyEWejYzP/mZMpfYOv6sZAZk/o60Ay8esVCC2tyoqrTVMJhIdaT9PvlzyTPZbqiTef9dIH
nHIsvYJ3BZ98fBNJY/9PTk9DIYgqqJ7iGBfvE8GMyVjaU8g7JYTgE5VnO4HTHdK9z8luTlJo8EMD
gm8tTheqjEdHOMVN6IEQkaeSp7YAUpKYuli/iFmLq8pllPFWEKvGOuziCzJrYkOLz2JWcemg9bW5
uaQ5jRpsWeBo9vJ/ykrCSYGlxAMgPq8YUcIzLEd3fDvOoqUn+KYY9uM6AD/Xs0mSsBM2coXA8lmL
T4aRcx0hjCT8OZSMoMcwfF+yw/s1kJHn3CjhKCIQ7zHkWLwSyRshu/0jAsqQnul9rMI/uLnwqmYe
qrWR+Rccf9CrD2UCoKR9TdVvc0Vs69jCXSmyGPC3lTo5PpMbXVNpTGEIZLDcplC6WHjYTz4n8CNi
ECL58TMuq5+S9GGLJpfsuGasmzAiJCCVqdVxkU4JLYHw31hzQc9aCdpEGXWdpCbhGkFlrCJJq4po
w9ai9Z624H3G3e14EQJWeLeTDQL5/YnKuHsdiFbyS0ZwNSgdYl6ichzYmnsPUbVFQc7TGM1IMYKY
hlK4obt0tQ5WNk/fiNsYN3udkXCX2P0Jh+E99EThipnYmk+ksQDkQ8Na+Bh4K35L9RIJUq4u0usd
SQyA/Wh/LXM+zdQeN7zx5scbQZMoXXNDyn/i468sXBMNRr5b060GppTvPJnF7a/mosQRVRmZxAkz
oPyQnzkdvO3aDhM6TEDelUAGjQQqzenkD+9DTZjeD/8PGSIWqkDLmhTUQL1fwjthQfk/hsUCzRtS
sA9QYl6W4/ebCrUbvRtMS75F2PjoCEgf6dhuI9mgI6UMpjNT9vcJLqB11vA9ehvaFqcD81jlrV9O
KA+E8K++vBiH+6DNoYgwZbkzzmORn75lKQYsmwZX47vIkMpYfBcsFLw37TMgpmaijKp93Cbk+hzn
xFdIMPziiFdaG9EDu+8SIpYY530bOcuzIZvsAG7lWuJIQNOp2cFnzw3Bel5h1a1BcOm3jouTy+FS
LqETPZ59FyXDXb/QRStYT87YPOKeQiTibRlLYDJbL5Ael1XtDDoJuUnnXzwqD6nDvoJIZeWYEOvO
VYlrGmw4YzbrPM4wPUR5Hb1eCiCIOVaSzozvYp2gtOdKl88yVfey56G7RARZQJLMYb/d1UT1fcvK
5pIHOomS9RFGzhdZfik38v8CAzVc5P52ZQiNCyQByh/lyQHz8mlH7Sk2frUWAWZT3f0+TbKk/wnj
VPCt4T2hTQEBsP9KFlnAnCgixI59TnmDXJH/Kr2d1EAn88eVHmosC4mAbs8lQml6pGdjX/KCm8qR
e0PWC3fTgDTKW+E0K2wYuzGgOmoX3X0OYvk8oO/VLidmPsgf4x/pKhxTRwo0yA0YUV7Ek7aG2cFH
tKG2WyjLuhYbwqJYXToXkvPmDByBLyRd/W8SXJkvK2G/ujSUO2bnAbUMida21jGGBRnZpXg1Jxj8
/XUsuuaYX0qtFBWRMeoM3FIGZiLuVsieNj0hgLoe6HySBs6bWnlpox2tM+X3wpUPhMwkmVIJR2/F
LBhA7jJqpK0zmqPnS51+wB4lpBTaBegYVw8SPmlwKZKjSpXZwiPp8FdJV0f8k+Rfvl51sjnt0OLg
Lkg4a139Ml9KacC+mJvuYeEhVoMz6YHe0NrYphYQx0VoH6kV3rLptyC1TqBIxtINBKRwzIq42hXm
rTC0c0ubo1Su3T+RQHNYs+ov/aIKHpDUBfRt/tR16eTZWDOzgIvo9dM86LG7iqNfgiYrvtpR9A4V
HEvn9nN81GLRXEMAz20WM8axbZNRSHSZbXMOThSwer7f80fy+lT0TlxNbmxClRsEME0/5ZVQ5gb9
76WIG+1bp3qW8IQuHy7/S0g1DOHw9M5JIo9jObDfrMj4QEEFV6lRrGJEEQTkRMDHyQ0NA/i+o+EF
1oZmwno36vPfTM/hgUAPLR3SF8fPCAzH5ct53sq+jHZLxI1LzRqKg79byKuKZVD8ae2qNTBmSFyy
jv3jqccOsQFxUfn6EYwuiWXMu09EJMR9LHdZrIUa6z0No1hrIa9bu3Diw5dog4PHRnznjELGeH6E
85tAaq7YY1+otG/rZzINafaJXVMdvbCklx/DAMhilSNwPTOlJVOjlhjFPY8qxh3sQqcB2t/82IF9
eUdRlpRoK24NmqnXSre38Uu+DSGdIBrXN1GBNSVKE5747h9ICgF+BSKdUQITDMm6QArBGuQN2Dy9
KLf5nZzeZhzRH05dYspq37NL415odMjd7kc69hYW+9EVSfw7p/2aAd0kd1hRJUA2OEheq++hIkKh
pdKeTi4JLWfIKkcAzUiMHo5gzEjkFiFwXO9n0hwdRh0iSuPTSlxiFAB5M8Uoz1XqjofQoAwCHRPH
9iWuf96eLdtSXZcU2BgOkW2Pn4iILGouVvI/7G5Epa4JOg+kYKvl77SoJrKs8aiImb91g9diUBhc
WNL5z+ODJzNlC5Gx322oYEuPSfZ///p8A4RuJQqs3qngSQEd0LLndAtz1lzKxwV835XuBBYv/A8r
4sXhq9wH3zWuIxNCxX4YH88rxxoCom9TY4FFZESLMuLS5fQ+UJkuEm1uzCnkZi6KA+WzjffcpN69
yVy0t9ZYbyqNOoh2cwDC6iAsp2ms3yGhWXfzrscsWGe7SeYoq6L0OuOZhULicYSWwhmKUuIEupsJ
dstmkNn4PH6hMGVagk0H1wSDGCDVrUArub3upRKSrPnfPiD7cjP5HPuaYhi1Qc5WBK3UmBB+h2eD
9FIED5WuZvyWO7pTrqUIvUQhZIqmHbOsTmj7vl4F1DQIBdA0OtWlFDASsuWEL0kwhJrKUCQCf/2t
ZjtEyk0dQ8N4qGPD7zT7Zia20n6Ue+UD0eonpAR4g0/2+KKesuHp7FD7mzrTmWcFGWGllnQEHUVe
uAUUBMfzBFyQdob3LNXSKKLFBCC+nB4Zvvt7sUJaoxtJW/jP+XU8DC4EeRetN/H0KoVSBP9ITty/
WpkKfyp2QHuu7o+t/yzfuFitECVqfwlc2/k6UEe8swsQXhaPV6g7EGx7mrrOLovcD0IbeMrbTL04
jQBdm2iZYNSG6pYG6zWy529HgC0UAGEVUfTyK4ANvb1/o57ID88e2KYJRmAjjU401SsbzbQlWjrh
chFameVLmedimzbePcjllp5CsSqwom8qwiLbfRV8+I1iCG6WilXc2x6xUYELHDee0fdJdkEej3AE
mTETjo9Xw6lKzHac7RUP2kqTIIMrRfcShB6louGT7aPnL3XgnGLDeA4TZCC1ItyDXWlIqM1kvYo+
OY0qwMDkMQzNpMfno8RQH+vYEjpQKudtaMD0d8beKvjRHNYlQX2zduOK4t3qTCxYFNorbQcduBEb
4gu9o0znQjd6MUJK1Q87LJTCrVkXQ3dnVRP7TKwv1BkUq2GZPsLUpYHLeHX34VoDQTss8X/w+/bX
GsVUWQa9aHnDLnMGUe5Nl/05p70iR8gP7q5ELGhlvZejBj8Mw2RmLxSns+NUzKX+h+AqiCfyCVD2
Eo1My4YYE3Unrt8xFJL6vRnJ68j39dVD2HJpE0JwKb6rJxyJkVhqafAnQDSJiqpXKAFUuiSAqmYw
mq7zf/RMpHEYfIKkJR7pevlM3YGqv5onUIzz5Xrv0kmGy+h6KWTDqTc+ANP5G78rx0Uw03Tzzly3
feMjnD44Tb//yZ/OXfQTc03p4zu3AD/cAVGwdyFtMa1mTaJSqM1nT0vBdBAzupQ8sjH+ZEmXZ+zO
PkbMwHXF6Xm+pTmsZNwtRurdn+UWr2CZmDJ6M5jGXk87zm/lRNOseLdW+o8HL/3eaWBEYNSfluSE
ei7LQ+zCmXvB0j3abQ+bcHx0wgkD3KbW/hkmZduLy8StPCtq5QeaPK2peuQx8G4bjW9Q0Gbg9Qm/
dzdtJbEf7zXGgkP6KLkLHSQL7g+coKSU7Xo/rCOlIOIPaSwcjx/NhoYEbAzhuNHq4FBAbvRCOA4R
U0Onxzbn7r25u1c6h26BQaNkYTxjAdzjh2sXEF4RVVPxpypkEdxequJBY6VinA8qqKZo8f4igaS9
4ZIfJ6cU+nSfsu1zjEyY45DxrX0IhTDuXlckv7edzPdzkbMTGQl30E9Gu/gDftmZ7q251kQuBbFd
Jv5Mn5znI2tuJpzGR9BdqVZ5KF3g7fYJH+2bqHxH7dv8Xv8foMv81r0IQFGea3Ei0D0rk26xiRrr
X4lfJOE2r45D6laYW9Z8PHezF1nVkSrwFRywZrWKhdZEYlA/OwxVzh5zJVDLHsfAzepqiaVltzgv
tGBvHnKpmSnTdAtkw3GgdbL4/XCVwg99skB6bnHvUYMxN91w0YC8+ugqTiD4krvnaILhAFqPUCQq
U5F3yOqnsijJbxnJ9BrczFnqTDu5Zusx3vChrXdfx/jmImjMTyGw0aecS3JMOQyjwhgOdz43b0nA
Gp9TReWGwpGIAHC5xraQzC1sCNmozaD+ZODHkmWMtiNKuSFW9+IZsiBL/OlqS3H6EgB2TdRxktzl
cW4VKCe+jGMc2DT3AxrJ91/IkpVdWRX46jIgdOnHUngZDt92QCQUYjIspGOojAcRnzLjBOkmrkD6
HmnBkQdQA/W/h9EcmSN3m+9R9G3OkZ2NA2V0s/v4LI+dJiWnGT0r5hgMyKBE+JFidVagIlEo3L+n
uClNBvEMUkprucfA5NGVBfe7RMt4ywz59Q1cOsTBzpGHkE+XdgTeALILzbkJl5hZIbxwGmcSzhIa
zuI1FQ7wuiLXxLs1w4tfudyBsiLcofRYA4SDXYZLGTTdnehURRPMb/ynEOLpPwbUcyqWysOPHTnG
jM/JMRN+VajfcD/4hyiTkzykyv24dIvH7J7uxVAEuZRtQtVVNLbBMXl2XDwb5Eh+FO1RmfDE3ooU
sYy9FpXqzYuuieSa+lj4ikO1//FI2BDg0KvNtW9gv+UefbJAGneZjqvNra2R+x19igPDP9oMLz2Z
hKRPOjfVSZpoNIODQRuKrY3FFMoMEtbezzLPR+W3UaGB4gV1Y2Qyn2BCVj49GvOKK4MGOPrC19r8
+9PuKJHzylCYHHuaTC5vqxRKfSmp9qahv4D+Gk/4vLIMZpNXVaBAcbt8AEkGwtGkqn6JKx4jvVBa
MskaSLTW6RSstr3AAoPPBCoiS1vKGXQsjTkCOejlitZsBo0rlBpAunIOcAz0MrFhrtH+EXKiFOY1
JP0C7iMl5HjPeeUmnvA367r6zyeau9/YSv/VS1uXDp1A8dJJz2LnO95YTEp5c7jWruD9SJk1ekRh
PS1UvXBLFSOZ3kHQ0qscYYk4wnsbUwmE0Yn2hILlRO7Knqf4yITsSVQJ4d2LCrRcT9h+EvdIAKSo
RqzEWtyN54JLkpMEYfURKgAl1bvXzjWXzjlycQzjb7op53TvyZKAkWKBoHyOpTSMu7lst3baFeCm
e/kO6+2z3Sduy+jPZt3e0kFV9Wqm0KNh0dHgPRwX+jjJiSHCpWbzrf65sXNbCSC2Y0+hbdNWnpqb
fV4uDnRSv5QkVD0Q3Ld8cPHBbIJDM2UBEB9de8z8Fyf3RAYUJbIayKZfpThPP+cTS8VqjFut6dIp
p+9La/ieiwZtbZZgFYdZ+51R+lHelgkIsiEBy7RyOfFXbD9NFW5DO2G4EW07JXudfKD3qlhyw7ja
g6zp3USXKFP3BrrVN+C6CyfNYINNlMCyfldFwFHABvMTYChwyRTG48jHL7MrRoKQajrMfQUvF1G9
+OtTxWkh4smXy8cz+u4n5YQUHmloRVR/e5knZhQVtrweiYObya4kNT20IbdUvLt/DaWSB9/p5dFy
1tKY0wkF0ingFpScjXzPqbspfrEq1SUtOt/j7S+vtsVzO341/ESqHT5t0ZSUxuNMvELutK6MNrCb
1Bjt8so5fJpXZvVgBxbe0j/XS8+mGMB0yv5Tmv/84yAUpFkApaCIZ3JfYMJvQeYyEO4+AmuTqhDc
xn4edwYaNJytSYzhLVKk7wLDZNSvcW4J/Jvm7W73Gup1ka3y7MclOqkEmTRENNoA253NEOCOHb2r
Z4S0xHWnIQr3FXuZwk2nENZRHAcZyG6kxZkUPvSrnksES/6ibFr4ae87gVmvY/ZLYRzermP5u/7y
9byOlCzVi+XjEn/xW9v1tDNlx9skT3MMlHjtPGFS82vfl78mGfpLIVbfW8YOpJjacheDPISLiKq/
gsRITrQmizQU09mult/L2QYXXlza3WZJMoCDpNauk3FVbDjQ9YVZeqyLODXBv37+4v+90+5ZzFKw
yc4WOLi7xT6vpgj+SB2VRZmnqJ8ypulH2PLRK6eRJ3fVFajJJnAbSDy5mBzQ7CHZFqG6A4wWQN1Q
kqIVxZw/uN2lakUOPtrW/FWimM0NJY7UG5aar6ZUhON7SHLdt/2KqdLtc1Evl5q9h6AdIzX0OQHa
zI1PB9590Oknx5hahdM5LPU2XelEA1ioKJ9U49SFI9AEh5iqCgqLo8ralQylGNRhuPPnALc/9ORN
INXHzBWp5X4tHgGNsOuSF6YH4isnMYAhFcoGl6DoIPwo9O57GCBrHiNEADMAdP3bnEp3EW0cPgtf
lVSd9xB5+DItF7gXUbSoiG078iNU21V0/7eWwFWCqvmo0rWQFBMT2+5iXgCnxzfvBgXFb1nR+1zo
TgWb3gf/tz7li/qhkyBYhGY7eSQWT08H6V4moO4H20pZbgGW216sAN6G7lvuD3LWtHgJzVNs83xK
tuYVws9yOrVCsPbMe9PrlKl++DDF+N53/7jbxTX6+KOwzpqk8//5qQD2sue6qA1d67msEzF3Z0ST
8FpgKl9Xm+MeC+ElIExlMfHb7GWl57FfvxJskGyDqcB15JkfQQ8GFD4vBxSfR5JleaNar7WFDx+V
YKsetj8eOCaIc7SDrGRfPe1Xb/X38qgxFeL90mVpQhouLEe4VWSKFZdj2C/AxCB+02gDiyj2uBnX
BjG129jJmAAokiPckgVVFqVuFSni3bPJsGwdVgq5CQmf6QgmRZBbiEMA75lUCH9tYaKHTeBO+C79
BRSX1FaenQzzO9I57we7e3l65EI7UbroJikOURj+sXBHKz5ODzZHCQUgAoUd7NB3pjak24B/0Oxu
KTgqVpqgUndzejYCqaM0VgNigcWTl70No+J7SmoKIMTJPyTeF4WBMT0aw3RH4zFmp6QdwATl/xbK
+4G6Igprdvc6HLvhVD0TImUDez6R+lrqHy+XXEZMPTumopecR9Pbe+iLL48PjkvQD/OzrKhrSI7s
Bkm5mmrCDG6ESWqcGGvXH+wzaDRc/AZ8QiY1r+n2hf2ikhzOLDF9PcvtjQZG37lgOF7WP317rCl1
cGZNrOT6PM35/zZiaZ9whihRjxV50kYWRYcFyJemyEMesYELQ95ttG2GVVWiz0LCVBK5qc7GyxH8
Ag+UuBz/MTA4Db/blES16Je3gcfvJVSED8U2C9TaqQIlPrMeZMVVd67HvAcKX1lxDvgnJ2lAsNKX
SV/NIZl1VgAeOHkRijXFOucHx1tTBRQsZjWZiZyhw5odsHJ3UKjSb+40YpvXKPKCpZ+AvcM5zagS
a/Dd6kJ/ZIfQb3fq9LtCIetmFFmiW26lU97aMJAFs6XSwVWzxwYodGV24E6t70iQcKbB7WnyjP5c
q5vHoiIkFDPoFRltCzK7t/xM0sKumJR0CdnfWIIqIvCPi/yq/mv0anQYrmqqlzzFw2xvz7v4/ShJ
OA7xHysOvWKqHN2pPBh7Lt8N/0apeaseD8pqmm6tZjbst/vQ0IHTKhy1q1gjG6K45W5ZQVrxDZ4y
EVODyF5t3oakL6Dht1XdPElcLcKTatPAzGPiaP3xDWs0vibZWhKQz0uxCvRcTLI7Wj9nvjLDQi7C
9ATQzQNUQZSizB0WHCVGlSV4rVznTeuvRykI10s9d8p3AC338DsZKukHtPtp5+66NezFAkJqCpGR
exkWQX8jtpFhw/JzXB3/IKo8T8/KLSC7VF4sw/l/xKekxxuu7XA3XCVvuLHWcwQTbgp8mPIBSrGG
mxv/AXWUxw7DbAvSB2GU8vHUS/IusYdPuHlTQk/8yRpq1s0WVYuEeU8kMDwlNy0oZnYmux+RNIjb
wJXhh8nHKF6ghb5SPH16hdz61JkRNFMa29in1va6ZlAZJcumzvWNIiI0UeXI0cOv1vRyXmPGUyWs
N+Fho155N2y2f/DBwPi4dvDbTAzIsoBp/YjPHHMwVxFuigXA3Rflq1Gne7rxDHvD+43lSE3FW4V5
FJ58URITkreGIBJFGxhzVq6MJjW0QioCzT2H/sUX/Tv1tjnyylDzWAnefRWQQNthh8DKiSBEcL6t
1JGNG8r/e64mYmrWqq2qhDdAA9Ndaqb/TuGS3tdgMCpzmIR9H9iXVsgPAsV+63LkDF1muP4EdGJW
v4P7Fx6vK/b/9f3EZ1jS6XupylgWXStFLmJMQu8PiQ56Nn6a3ioSYg3S84d9YudWHwD4yBhLvWWk
W7Zx4O0kFK/zIAeRvpZ6w3lsTGDxva7+hPtKAtqfX5/P+QJlHmOYsz0hzLJ6+O3YBDa0XB30q1Cp
6pX4HtGsSjncQZTTBML8Ofvjat8EHfYuF2y30SX6s+udBZu1e4Uqi8N2Jui2XHxZB48luVL1R3J0
ZOkadzwUf4fauqrrzeyrUux2NgK7z4Ltf18BZMgqqSgy5xhmHhoapwZuyWx1VHIsUIc8xUr/z/eC
bePaVQH/cZ+D849de4IG3pwyXwd1re7EvTkwcAARqYa6kUdTzcb6Fd+tZGyen6TwGgdD7hUz3loK
pHwzdvJb9b5uG8rj5KgQYH7oxgl+rAkApOPJqf79aGwLd2/YlbmUzOXV7keTrcy3/ERXYcnX3i6B
zgNpmRr8pYDoeNTqUDzxOwj/q5vgwlTn8xaKeePmavHleH/kYZZ2PJxQEJLOW7MhIeLjOzzttENn
CvlpQehmx+XmROFlh1qbE8NBIAO/Xu7nEHMF6sbzL97BDisSVdnX/W0yB1pkMeM2ufbqq0nF0P/Q
i3dAGzWgdgzzyzuFys0ZOPMw3IZXaQ5KPH/T4Y3AAV6AwDljdrgHJKFzwU3zg/ediIKBuX1D4f20
ndPHXENr4TzlMsLugcOefy2Zq4mQxHkhkMIDchQE1SyDybq/ZLcyak9i5haJS1+kaWHiFwHtrAxg
7Bzd+3/KcfgSpuevBB7J61NkGipdKVXDEzLx/jdK7ALykoQX+viDna+Um1FDk1+47PE6M7ItbKbL
VsdCauHABEkkSRB28gxORgL7BQpTjeu3NcxE2ol3fPXjORRozEGJ8QlrkvTcNVdG2IImdgxqRtIn
ILzacYVVjfvfaYqg34+yvoS1LC3SCgyCVEN/o9rOHMRx4ocfdOkaaqx9b9Q30hvI6KeLw1krz8pE
5606VrSWeikkXPj96cCZ1bhahvavm9LFedMba6mGsfxEyTuL5ZJAFNooySeU9WRr21Az+F2ZvHMn
7b44FAwpho8FvADoqD4UfM0AS/YGT6vO/tym2ehqRviN/V3qh3pqqPOXLRr0HG6z5gft0LORQjR5
FTivLHAHu6fJSMc+ht0KtyRuw8k5S+xIHPRyZIEkZQ9S1olMN2zJRURlZHGXtu9musw8kY7lUfFJ
aZXBjlCWHgNceUHpoAwLQ1N0Mq0+Sep00wfcDnUFYbwOG5L1ZrThQvrjK9kqqHOdJXJdD9ZXdZGn
dElpBE0EWtqhwFtJUx4Qq2IMw8ghp7I3u1utVd41yfnP+1h3DkvR95CsrUsV7BsgzliNpKK7Jzhx
3B70mBC2M+34PR5Djpb97WYfuFQ/g1nzmT5ga7xdNkwCZTlKDaWawpemi06R8HlAD/gUjeiTIejj
oGkhdlmCZMxy8yTSm4zOjCo2OwhMLurW6mj2AGYALiCgWNkX9J2sdkfJpCqzBfJZmNAWeakyecGQ
68aYOtn28Mu4tAsajt9MDnn9tALmFtvG2VXtVT9Bz9HFdGhfozYRv9mU/1iAqjN/mHpn+ryvfHNg
EjeXi/Odh77tbDpqwIFo24R9L3op7V7sHkeak0II9kr6fybWpgrxAaDtlBGmV8E19dXGpcD3rvld
YuraTlQzYD6zxMxrn9tGKAHVpWY+8NRL6AjR2WUbj4qCboYeD2DCYM1kbQrQirheKVAQH9Z0f/dF
nesQ1MIet/d+i8rBOOUFYoCZUIg+EWAON0TyF/zv/eQXZGHW4SrYdqHLHSIM4jUyzW5yDAFMbXBV
h/RRxgRbEVxb1TDq+i10dUcikaAXNp0PzSVda4k5fVIULcEdRqgb7tJO1eYdSC/ilD7e23oxtWje
WtGjfqqt7T19mVuuoO33EqCYjFAInW+FMbBLO+wsCIL+h+tY1bwP3ydDcijJq+wrEIMgJ4VtqO8i
eY5ckqoLFykAHOgdcdO7ZphNgOXDSxr9vB7QLgE+cbYUcyoDC4HoixaQigjEOayKR/9Otj3qFvdO
qLsNr73JuPYAeavM9jqdUbJtb60vs3Geo5pnYH4OmZ551kAF2Jup8xAZPOzwE0p4kIBXbhN1NlTm
g6H0TbZX35MWfEmNrrt7ygE6kTrNENlRUUcXK5ssJtud+eqQ07UXXuh5sHBX2xBDb0kRvOOLG4CF
jgrQ4ozlO1Gpu5BwFHS65rCQTQ9XucffSBwCHqG6EWc+5uT+LclX49uT+Zq2aicj0+XDaM3w02jj
6jDFdoXv4zByHj6ScyUSkF4qT0PPRjuosBzLRPS+9Tf/1C7/8RtgMq8fRMLvPp2Qe063WYEIZf10
qNnapmxDodDOarFUniHN2GieZM7Nx331Cs4wZT8YomKxwZFfN4xeGP7RG9N0KKPDWUbcOwWsgRXK
qfOU0S599xNC2PQSmMQRsjtO3JXMllT7vrMQYek4lnhchRVhUyrYXz5xJgzVAjvQ3LMgdxL2aTIJ
uVp5oOa+EwpbgYGCdYETjlM5IPZ6VPX74xlkWUvIcs+FA5m94vmGQFT8X0km8zufzmikbPzjSzeO
xI9ZSzmn91lrIJwCaLM9MCewlJ7bov89oMDm/wcejxiP26YQ3BRuT5NDePL6P3NwmIJpzn47/8wJ
PI+eIvzDuucOgdsDtkyVovIGqvVERLLiBoQstr/7U8ci/mMRGDMWj9WJEQqORccFsC+GyM7Juk1E
uV+2DuGW0pLhw8rZ1vA1fkaUg2EY2NQjxQaqXNBkw7cLIhvZHIBB7Jkg8CRtQWA4PcTFS2SsH52+
YoL9OHWwQpqJCFGYoISauTxQ2yLbZ1+xtUH2ZE8spyS1DxkOcA0kBOaH6vkNlhuyB0t6ULAWHXq+
2WqEySKWSCkxTQOZkdMJFAV1AEumxeg6LKyURXzRlDV+TyxjVNJIXTTp1dk6+bEA0PyqW3RxyaJt
0SklKCOvTs7RaEhEEcj21uUfWokP7xdrI82LO8fWDTf0yojE1S/wUgfYVeAJsJDpDViqPETct4/x
vgdg/jw1i124z4Et+lbHH8vRU3jCufi4Seh6H6GLFo6Clp+5t98FBBv36dn7IHJ7ld0cii/GpTtT
2xh2WkM/tJgCmNtMOpyU/6CjQDeGyUz0C85PQuz93hXwbvkj6tmIZekNQ434qOOkck+8wHhbTYZJ
GgRCDooEAy3eH4kt2ccLdUHSqSD+WMuff4wIYBokax+s6syfW1MFO5lNod1Zasu1Urj6eZohhAip
D5DRX2eMJnXiv0URfWlscjKw1d01E71Rq/83q/f8Vkn0EYqijz8T0pxRCQlWe4su6BMBZLS6lSPV
CCYFAD93N30oqGAdeJhZe2dy9wRS+yG84BGXRWb+t9GGvbOmImsuwz+CMtTqGKaj+sgHtDb5Dqib
RtA5/5qeDb7H0oPEw5NFIRWpzO3pa3bqVYB6RjDgDX0f7BjZNvfxB7P9fIlh/pv0yslrI86+HtYU
+akKrLd73dhKbI6WgU2jriyyLAIquu3xE9TylWMFayRocl9g11dN/Ih4o8e3Fvn2LMWAKUTrAb40
EuqnYYoarZOccOJZQ6uTlZkVNc0t4aV/4KNXEpUFy9+axX0XKPYWxgvle6In11K0Mz2Wp4EkcM/O
8UIFBwegTAIwKAawVY1UQQPR5BfDzmUybAmrT7UVqLpcRm9n/gej+XvzY+rHiN7EE0lioLIPcc3S
UA3yGwIkioEwe3CClFc+pxivQ/336HQH80cM3D/PWBwHuQRmiJxPVhaEiiYqYUxkBhGJ94FxVXZt
eUsBjQmMUh2/JQdV9HZ6J6p3fLxqFw5Iz3/OonUDdHw0zexzFNNLmN1aXhxI2ZK4lxsTuEYHydzh
oFLC2YQVDv79JlZzFRqqbNh5QYiGsNrHA5s/oZL2JlEnoJrU50qwYCMIjh1XqHlV/+v7jBax3Qgm
sSaXAikOugvDxqOfn2txOxKY0H84KPiLy89S6578AUss43eNaaBOQvshgIaGquQsYtdS5IvI7tiX
/ueuBScFzfsnYo/Ia7bj2KprStziEDMgetQCKi2m70vRGc389rUemFvvQmIfo2XgLksZeP3YzBNS
yHUZChtepgT9wW704O2riiRxit0k46/FoVtrxiUcZ1Rj385+u2d63aXfYs4XYcEFhM2g4o9893MO
B0Rfa9jqEIgaalbCvmJRkf3YLxUe+l7X/YwYCumIH8W0RXYiuIjvUv4lj6zi6X2pLEza2WMWFQat
BeUsH3spxacAF/kf+la9E9JvrtQwg1Px20WYlZVLEK7Dcmwmo1NSPW5GGGBjaEtT/XzJW8LsoghK
74xrM38aGKPQwUtG5DeK7OnoeLkoQBvPwkGra0nXp/g+l4Qxb2rv3lzKEahFq1RwhdZsqlNlV2u0
jCDm9lSGHsXrSax4ib26omWdiEfO6Cb5ZHDU9aOPRZgB58gwXXaroqgsvBVmOAKaARl+j7GeJdvJ
Go+wJf45SxiQOlu+6MQfi7ilH6Bq+zmQ523QaC+UQubey5m4on5FKcCbkFYynlZegnStftcQ8i0Q
JG2f+wJDQZGJ+f6r2lLHPzK4i8+oXI+9qTRJBYWJ0lz/55wmx3vPoh1znia0tdfAGlK3OmiBjPfB
MYInvhxo8rR77n9aGinBTa22bPb7Le8LVhVXWZlL4V2Q1CDKdFlytt74jAdsbejivMYMXunkzxNf
0xt7nVe/uPJM45mFvGTjaQBTaioAYyfbcTLNT5kXlh+hW3x40vC7xAiTJHn8dxhlgpGKR2XyRw4h
Cst/N9jJIz9DvFpWx3JZ9Oo+/R0pDpSSYmCFWWuiM3sg5kTn9Xj7AbYdouAxRtG7jFCpVyR1EmdA
C9Ziu0VnQfHXY0Mo1GU2sfhT32xdD7Bj/zap4CzfqmFwk0TVi9fC7Dkz/8RzPMqlOTw1kLmt48cg
1bp14oxD4OBWSXVK/u6DSyODGDUn5I7o5+hTLWxz02QonnPtngYUxyl7173XsIywm57ldniDvPvr
8fDUwVQf/J/o335vMvhKIx+/nfkjuy2mW3RObB0VYsHlcDaXE8vkDqM6E3WmqB2VhHjqfa3r8qtX
8YDThF2GhyMV6vUSMwEBLYyriaF5Om1K9j0Z0/IieXk4mfeId6JAFjNDgknFzYbQG9Gr+V7gyrnV
rMaVZuKDiXZr3F3n+2WUhYz+hnPomLiunxnfOKAA1YSqcLCzH7aaPFd64Cc0euuAgIy6rW6dfLgE
WdH3jlx9b1o2RqXI7+lS9VJhnMH5fsmzDCUDHIzFE018MvDuAwT+5yoXFqOYNCMxl3chbAH3IXWS
OClg1sIn6DEz+OoK6tHWZ22o1Ok3kElTx8HPetlopDjPuT7s+dthcdqxm0FglKdp+TRsRCNapbGg
LspDZ7fTGa4Z7FLIFG60S7diW1R+itRGR3lLC0I3pxE/YkcRe4T0D7IWdQknwH3K6txp79ae2X9y
pdoKWgupK6rMhIloP2zjkyPjXzT6ZyMtNwnUVeGX4zwsonHIt59uyqvLl4DrBaGQpVUpdF5g1oBR
wAFk3NA4Iqga8nUCCFFbCe3zSXGD70MnfiNZ6U40YxrdPDPlPzBQeAYhloZ0TbZHgcOZafZ0+KJY
jNDgCxxt9OA+9M5nkZjwXe0qiiEncA9NTTaS/LL1Q2/aX4LAFD+DyrABcQQBuuQA+Pp7lLm8NAhG
MjNKxdwQH458JamydnD5t+CajRlXYuFDtMocv3VnKz7jkh4rd5UQikOqq76WmhwTFOMWB/OtZD34
EAuGCx1t3g3lanWTHhAd9ks4qoMMf31M/0h6CM8InCkEdhQMmY1qDejxBx8LJC1aiP9fuggXDmx/
qt9P1t3g6XWn+leaU6BMCeHtmtQokQhZeZzvsrYGrPtlqMR7ar8d/UWZu5FKgxESP7DVnNRDcxnB
ZXEYElI3FeQgbLnSjBQwyZbWwW9R6hy4C7Jqi077UgLtiWqdJuTNl82ryAlj/mA7vsI1vglAQFoD
AcS2ID+7mutag+D0zCGEZcKpt3WtI1i5YombVupqxyTi4f9aqyOrrQuF/6xqlpsKiwdXaG3Cnmmu
lfGEOMtpZP1//Mm3XzrtcnMvWeLufgx5waVN5dQIHEGFyWwUSECNXIqjcAeXRnyvs+A3WNtpFKUU
/UCaapUzW73ZsJTuzZxARyeT71MWRzVPpmfDxx7Ucah/QgcbcBaL6PUVs/QKj67OSpW5DGpZyqHV
7HD6n0TcHh0mX2ahT7d6h4WOAv1ahkqZqgTTxMOum3+sa7Pguzptcf4jplc6u3f31SbUKHnliGRd
GwK8U6IYx4Hpi5+myNXxLJ0XRvo6vBp81QP0J9fnfWMm99feHjxwBDUWiXF/rU7R0h5aTFt6W03I
cDCbOPuNJP3P7iYmkfIBJTnnq8r+OpvO31AqSbUhOwajb/V1bb+TwKf3meBLLOMqlgpV+nLx3251
5y5SqrvQVK6e0JNDX4J/jccRlW/9ptibtjf8+jWCY9gyonezayPQ6ZHZuADkW2Yvgab9m1HSp/zZ
ZW8SGA2UlZJFyN0JFaINLSt9K9ebz6mrhoYRR9HWWws9ITgSMY/tlweizVovt+y13h8hpM2ZLKAq
P6uPic+A+OQ7Hoc785THc2Ao7McDkB+ySk1/LxbVew7ovKaXYLxsQH2MindGj302fhmi/cs/KLoV
ICM+6fx+TVhBKxTrpYAf93ghA0wnnVZAP+85RN76fTC7tQrxGtj26A8MpBc/UX6k/ndzrwI73TG3
qFWADznx4H7r4izcr+LgmZj07xwWd0cXQJVs0nkbbhrB8idcdbaOPOsobmz+1nrcqT2zBk9oz797
2tLKI171j/W5tDpfG1/XO+86nEceUwsIJinoSCmxOyh5JAAxb7/O2ryEXy7toU90ki6CyVkUYCh7
ef+4p1GpVjj8Dpz61Pb7/ju/U314UKTjZibHQ9XMLcN0gmfTgF4LPsjNLfJ3ODoRGMNA6gJ6hwdS
GyA48zWpv2KNP+HyiHGm2LMx8Rpf1l2yCmpkNOUhjzelzN3wrvZjhmxMhQvbc8SW6ROhQ2P+8Co/
TzML3zxKDqynX8mSkOT+NUNsyrmpoVgqq6TBrCD1RogRogqx+2pEDZj1c4H4wGKtWG9q7FlR3loC
QpD++YGu/am4pvcRBs5jWG6eKJT7MZlvGXejaTSCLyAEBb2AJa5XoIGpz61BzGao5dKEraWZKa09
Ye/QZlcZRBv56q3cwKonWfylmAM/vseB+cFekKeXWmCYQJKT/ba+pVYU8dCh0IYX8+cSCkEtmj+d
BoK2DWhnfUguLwDahwpbo5+qLqvVSa6lDB0TRYoYJt8PG2ikHNMHk/Iqijj8/5xzJXwc6xSp61C1
HMKYL57rPFl6wbolmWbvrSPKLVCyCjg3I/mScKJNZedHan8yV2TW3405cBItXWy1yD1BdkdX8vDV
ajHsSWRkJS+lgrNWXNRV9fwS3uMr5grdpodTFpLfG6B6kdox+nFq43NIeN1iCDBDg9CdRJHhk0dP
hrZJ8WoAUcFKCUTjiszltdKhkXZhUovRrefNj7rC6+N/uufCDps7mcOra8/fM//7+Y/oZu6pw3KN
oQ+goLpR2FI3mtSuiXAEv8JZV0T+UtGvklpSpUBQi0UM+JYQL7NO25NoGPYFTosnTyKzpMjNhrhp
d29E7brVraUwNGfUtAg1+kK5vrpn9KxbezxwyDoPWMkW0sRIH/oQH6lsRbivC3+ekIM3/eQgLZ7u
qFsSVlqXMOMt28iWAioI2jK8mkN8ikLIaSGutvcNr/Br+MgbctH4icHYCNmcF3Ez1hkNOb4V2CD7
UcePr8dqMJtOr9VcpFFhJDJIlRP8THCtfkvTrnY2KB5ZgmoAdYtMxEGLX+IfDIZGZxELxCoxuj0u
0JXYJ3LNVOY8E0dJEuoyVuJVqfR0q9YTT67tOydTqMQa28gIc4wGNjVBnV9GDBCwNdkP++kbEvTj
EMEC8c2VdxjL6FlbmMk85MK5n8yrTA65gviwL3u5OOTroIOMkP682JzId9ogBm67qhGohnrITS/d
Ylr6xZL3tjkduDed+SisfJEL28yY2XGKSm97VuRVXVOezvbCKU4visfgkh4IT1dh88gEfFJRTo7U
vpd6AOysbfu2OEDbH6C+gj0d4vB51iBL+klCtw2Mi4Nv2PwQEtyfMLHizvJixFiIiaTRb4YsK9Ly
K0rj+FTctyES733/8SSo4I85AVt7lcevXsbXzyegRN+XDxHvXN7+8AioDQCozC7l7GOGbs9PvlQu
imJJITbe0d0WbzH/ABbClxPA6DvwM+otA1z7idf0Ho/cPlNNnFRQ4hCxAop5rqM6Q2e3+q6Jpgiz
s46ELm/oppZpovy9X8sqdjqzinddBVWDpoHl0tPeN/x414IIfiXfx9CRB/EYv5SHpZ7QfEM/rZa6
w05ARTvhu3ddfxgqTPeYUea9WErwYG53Cxz4eH03LBShSatTFyAyC63e/CjUhXShWAa6hSVvRcw5
youWQZeqXutem2LSeSdHvkgKoyArdydRIHyjy2ONhT9MC4fRzCa2tG2K7Acnl96XovpRh8b7bZMT
cYnJFCeYU/KTK7Papk3Txm0xekcrfWBpyzeTFXH+VeLub8Ix//9T8PA22qQPAjkjpvWnrzgLMnre
iouCffzoQEQsFWr7jadoozA066fWr0fD5oPU7uS3gFbXEyaNLUBdwbZpEBw7uoeaeLALcnVlU1dJ
qz+i3FT5i4E/969Ur4bMoAF1SHIKDqb42OeZqDJ/WEhTxjYCPbjsLV3srageJhR77pGThxzNPKyK
QkveJFNGYi7JP+Pu5PPHswNNzal9DGF0Xqg9iiXfDvmCyP8NnvWVUzvhe+XOlOJDVFQUzXZ5JlpA
sJzlRUKJsjzpR1SlDZfI1XZj4bUUjGiLZPUYncPZvYsr82BaVRc4o2iCegwafw+sGLi7QZc/bMLR
Q6WNJWMd4XW6iqFMwiBHOE5nLz0omKT5rPxYfaL8mN9aqS2JqqEU/+p2B7mEjOGBz9qdTrv5n/gt
JgzBi1aDeM1lCE/p63Yhlucq3QISVuQ3gyzBRAKfMOpko/tj00xNoqMuUdO18nJx+RNld/b2Uf7Z
81MMXHEMOXjXqdmNM62a6jEulbipE9w2EPmIDegJ3usUNP1AyAlhGd+k1Ja9mgbTahuaWDUAyRmu
utrIaCo8KEJsAftUqSNXlAymrEdGWZ8QDYKV16CybqTY8GkQXcM0GEdzaZtU4I+BiuuWrYmJzaL8
q45jvF3dRBy8O0UjauENWzAg8S9KU5JWyo+QJ4DcTInGa+6fXzpFwhcILj1dF2nblAXtuuPUS49F
FIAJHelPN/+YaVC/F5tkSEwxo/1o5zKNdH4Jz3146X/wwMJNbMbsQfJi8ayZSeZD5FT4aoq9LPY9
QKkUwunRBAmfXdLpWeHo+SvlGiLENVmkd5hLGkWg7eCy+O4mVQO+fobGoy5CxCFDCgh+t0GeleVM
W/mtXI3gYiC0/9ohZDtpCuS7O/wuzHbVjQVUcPsjT+Q4PhiQZuujqx6dY7mHcW10h7doVgvvDTE/
uHFkB6cwTYnxe/mcFb5HeYpEsoCuboxd0rEQIyXrGwMxRyu0iFNFmp8i
`pragma protect end_protected

// 
