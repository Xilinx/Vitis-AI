/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2jbWIUIXDEsnmdLD9wX5v83D3sPkbRozDD7dvmQsubFTSc9y3sKunp6f
cgut1djkCAYEInchbGM3sTaVYeDFOFMNxsVG+q3JT3tGsRHDS/HZYBFq1h3mzl4cocQ16rmfI1Kt
wiEGXVJzoVkJ8Xj20WURJbSRs6IW+lW6nDd1d0pJZrAV/5TQALrjbR54FX8NYUz4CkVtoylygIx4
nM98wh4+egZHyknHCoNxkF6A5cmd0pqoIBQ7uPns8j4Pd2z35970KmWObupJlWwODeKN3OZWmcc7
iTPBBZ4oPuRymWqjqQfPo4pPiYxRFQWwLWJ3UO0L9nrb1DQuoOw6Tuole7eGBL0MqK+YJZ6os+ud
yZcv9OMCseymSV5PzBMJduFovs6QP8xwKMJC7TPhKwonb5DupNIKEeNhirg80B6Tv+yWmauZLTHR
p6b5S3MYI/Ghl0d3YGi0kSowYS5TXl7v6KrEXGt1iqgI7XmUL3hiVqt3LU4tcqznTA2nrR4EHqU7
p9FHbZFBCmYcMTJBhAbK3Qw34lzKCQO61wo7t1KFuyScnjOlIJXT2PbklX6Leqg7ABlR9G+nE8Sw
xBZHw6jaYzM1jild4Iy4rSDiNRj+GkgQsEaXNDFH/DyRV503L1TEjnPwBEV56ogix2KM3e4Csbef
zyr0rAAlWp+FKxuuwyOfTL1gBHIXsHnK07hQuACNYbnuPCLvvtyglz0I5t447ikjArGlV8Fds70W
DYnBnuVDz7d3YNEyXROk2EcHtpnsTPa/Rn2UvWSYne+HggaMVp/kBmOZ1tbEctMLVwkmkExki725
OoaWcLDM1SZbI3zR4FcFnOyymEusOqAIB8rqVejcr5bufyBbwGvom9gQJl91f+An0/Ru4NSwCuDA
SemTSMus9cDbKK4GDAtviu5JG8XFlJERYbo46Q/V7AtUNumQiSmd+fFBNxQtBrumcZtKZmEf583t
U58iD/H4lfKVTwzv2MUypsDugMgWrScvLPBXhb5uPzEv3oPAeRmh6X8kSdo4Ijm/Gc5yT5ET20jS
BQaettkGdS23ZuDHDo8+BAqmCf6Xbc+5R+OEDyJnAuXabn5KlQaVpcPDNuQOEXTKs4GNSeXwFeik
SruHXQc+ky0mQRzG3GLC1qqUKqMd/CZKYTP+8jiy1Y13WTtXyFVa3Ogy91qe0WWW7LFgOMUsVTGy
RnuPZezaZY/WZcpc6mM3+FlMIbZmbgVCPF1PnoC+eEiQ2jvGlOWjc/DRwqajFna4tIKmrrgo6FWf
kN8OyWU1YN3+xRENdorGC1WUokOZx7ugK07J7YVhlz3pMAOh+vduWaXhgOMa6pI9FzzPsWKSYObu
Es3QvRUp+kFirE+5f6NNug2aCGti9XQQ16/CWogx+ybPPUWwepRBqODEKzH4N8uqlLJx19sZWNhg
L/dPOOOlUVgoAaSLwgcaYHbvpCfa4GVNN/mv46ETCXcPdz4D/Zd93X2bEUkQ4vt527ARM5UTkN/L
UIHTYeZ2WBsMIWUmaxl3De7KXX8OpIQgeKo9Dhxw6V90dhpgNdR+38u+kPI+Wg1xQs17NVob23pO
q4Pz33sTVhVKyQQeyMOeREBPXughlOccncz6ntHTExEtUu49EjEkxQBYlPa/JLffhfo/FXD/SYDg
w6Lwo8ioDtdqtOH9poXqLsZoqNvU/1NKzsbvcXThDrjJloInfwxkK2dExd+uu9vwvkrq1kiNyroV
k8+OrYF3yKmzkZi+sMY8sAJmH0BZJAqEY8kyRFnqpPqmtgzKhSVyghYDBMw9MgP/z0msjJPbDGaG
2CimEQ2HPUscZFpKHeEnEAdmZ1O4fTTjR+ulf5eCZ1JwZsmuTY6zfLKVeQxkET2l0lUBzmcLMqvW
Qe2YXYGeW3b5SijgWSz8UjVt8GsYhCCxyGkbSwHBBxFnw7rgrCXsqaYcxIvwXQV3WfY7JXHBb3xV
ok0676bSgLP6rh8FB515rmx65l2/MiGpH6noAolx5tymA5j7tNTQi5FqI67N9ZiEFW6UBfE+eCkE
dyJH1znBzZtYr3XKDdGsF14qh18jKLzpbezjcYXBxGrng83Hc6+4MzVwEPjxRrwTLWeUqrjuNNdQ
xhMpftfYk2WzEW2a1B2iFEBHkd3lfcVyeZzWtuB8jXq2yQX67HtWY38wAu/3str0Flnuz3rpEFix
8Cxn6dkaD2T1ldVgm390HGhKaaShb/0PB60fuIiTwPxtvZIYEflkfHsmq3RGgCn5uSUEnxnRGzTM
DTvoaxsyy5D5n2ABo7lo7PN1PBS3qpHoCGzSTasqW0mvor0Ap8M7tiBwaBGhGMfbhIhN6iIU3JUl
EFiM79w20DvxX2ObreuYSsiOS+0K8t6XNXyWCIuSXvg7ctndq8sQiS/FgT6oaLPR8MswjD4K6+KY
KkGGIrDTM2s/kiUXqsULJRvxURvMdniU9pIhuuEEP82X8XfquqDtqcvcRAN5awewbDz9RNFIs2NR
awglKrTqytPb2nQ5RZFd1xo9/KDUyCLDq2xXvKo4yDqD0SRB0rtl2VRAAYgH9Hmxbm374ooZMg03
5Z8JyXWbgPHzk5bQspNmTmvctVXyIJKSmuknpXtouI5HvXM2cPNXEu5lwGLwV3grwlScXM89KLoO
kSPTHKpmC2xnmfSmL6DdHmpOJHBah/qxE4wAfbWevRNWh+R8CtRPnKmO4LYKS6Lw+ZF+EIkR71KJ
WXjxQhEXThrtBck9W9/baSw5xrqb6d2WXqb6cGG9kkwvYkWTQy7tirsFHLMUF9lnAttY0X4D+v8P
ZFtG/3cDly6UXTT3YqWjUgYEIJb1MWvHl7rg5QHbrtIBZ1VsjtftXbLENybyAKwjD6413F7A7ybo
0mGrClF7AVl26TqQTDW5CZAQ6FfUwKtPzpDFodU34PnWseLfCgZMtEFpH4lRbg6TeYmNXrGdziiz
V6sbO7+SrWdNQkzT3z49lBOwa2wVSnkAw5FG5xWYx67iVHJG9wLWuqDhnB9sa9pW7XGye4eACZNg
PlTRDE6n6FxHQ0zH15UGFrw94VLVCtPjSw/wn1XSSfrooO08YBAGboLCD0CXnFvZkiPfwiuWvLS3
/WJgexS0O5rQT4MbpOgCMZWFrlwzhka1Wb4osP5aVdmDL80nXFJ7nIUV/A3dZOuCeEGYJ3h/8GpP
blL9njvGeK92NM/vkVh6KDguNnXSRjHIfRZJGclfVqF9X3xKpm03ODYRnvWDjX6h9CksmdoIfmjF
LNiDCOjOVCzSGZkkb6m2wLd92moB5M6cuMT3x729eUXSxBG9oK3+s8Q0ANU2PNwobAYrHfL+1KPK
crV4L9RC/xAhugy16wRw6mWE6m1FZk08Zta6vxKnuPnR7Y6mx5agayGaBhwpPbywDpWEoa5g3tLc
FnNFM6lZNSLRG6/yhX8VGKreC43uzDLG02mYqio914sGMjVKpgPWRCuaoRXysEXPp1NlTFLPmyIn
7vLcSaxS/6Uw1GdkPFn9NkAXMrAah8mRS67+5fkKz4+MlC2ky3Ai4gYIL7lgqdaEw9pqiiwXgryU
yTvYaT7+Po5+uCCGBI9xH0ytMdhLLUQbAkGoumh3AigFrg5lP5tI6SbKgQtjk9Q/PGf6+tOh+YS0
2CiwwVlwNYwwD/Xrg7aq+Ki4J9NNp/VRl8gfYAzvFwwBRWgWbnXfalKNRPEpTdpEmWpfjQ/+TzRT
uP8GLFcc9w2gGOI1T2xVWQlRuFr3RcVYhGMQVyNc4+aGZOx4p+0jlYo3bBDpZJoYooQhYePhMaoM
ZEnkTt+k0rGOxFyuGjp1B1Io4JRT8j8+GIBCS97CjlmPNMjP0XuJt15Kkciuh3RlLS2LoUpegIeJ
ivFJcE3ywp1I6WcDxKZaMi12Y/x8ksim8SD2cuCdCORFqIsVhw2UEdnGxF/GwUR1dLEYXFR98CqE
V8beYLp5qEWLTh5SRBiSw83hq25U1wsNQMbhGwYcDeUzytXgWcHqnk/QMVwydoyJNHkESwXa3gFy
yTQk86MS8K33VFKk2rLbuSTVopvnwE79/uwk898NP6NeAlJQdXyalMYudd4/KAQKhkPy6kLDBvY6
OlH+L9ywoP6lnmcwJi010PYks5VdiSJuGmqvhMuoQGuxY3YQTSbTPlkODqA105HYaVsEclX5iGFB
k9v8cqth4NXWQfht2R+8uV+phhXcN5xZjWqSkyhvhymb9KSbEtn7oPz/xWM06cM/x9Rm9hy5K1Rp
DwLkHAm5QaxPImi9AP/0SLuGcfDMPxRP9MZxPaAMbP3gQ8pcE4aHmAl92V0GGFE/PPbEj2tqJ707
L8alxeSJb4a25PQe95HM8nxHM1ApNV0LKVNMRnbO9ikE3Aesdr7DnuZwqAq5yYrVaAXBeRep3r7+
S0EzjeGiryxw9apuj/SuIUtU1MzoR9IUQT5lARdGJi23+zKLMnAUetEcftE7TQNpR+EhL5XovDCg
EAgkhr3s32ZH4rUYdszOB8aq71vjabcXGO9yT2hG4zU4ZW7CRvTYL+gS7vHdJKrV0f0jhL+ahTl8
luP4oY/eLbISHbmars03i/+hJLxsqQOtksZBtY4BEujr8rjxk8+6JduIf+T3AjnSIChSH9BFF3bJ
A/8ItI2vXe5j7uGEDGqPKvh9hWdR/6akbFc5WfFfeTs7PrMFjKhIXnXcOJ4jqVQo4b+gJ1h34vve
tcjuVpwseglmFKiW2KOpkGLTqjEcZDJI1QIrcU+chcxi/xU0B7Jhw43UiFdHlsZZY5vipU6q7yAy
AEchHeQHLYrjOGVvDKTZW/NL72Qk/rvtYz6NcvLWseh86ZTKa+8Z8qs7abTqpuM/UPhsWDhN0uCd
jRYLLIcoXX+IuYFiol4kR4BxG4QldpzFZ+KY+N2zXqcH94VjhjFxCCKOc9r9cVCi+QT81+JBEkKM
RQ3oUdC5a3MVkenxLtNtoHaNDaWKgDJqot6AiuyGsAO5BDeRD/6Yc57HUleOY4JTPHfRfwJcdnTn
YAHNaYJJ+wTcLL2KSn38592whmAG/35ZAGm1+8rJ5e3mMvNz3JpTYofVh/KGTEAtiJj/JeuJFbX5
jp8UUypiufiRDZfkTF7jNSkPq67BG5IN0kp8VU6qyYeUfiNEJ6V+doQAbmZx7QHv1WDizPep7vtU
gHdaAT+dp+XarkU7Unzm5WsW4O5UnhpjU+1SThxeLLcvNqyV5+sGmQAgtki7vmte508+gdbFiTCc
LOf9WmQhlCJ+2fEM0IUytn/9+eOSu/aNXE0MFokhqLYsDcWJ6vyKu73Lkmp2fPXzcYFBhYfDkK37
ve2iPUOdO+V+Mpd0mm0NhuS1bK83SQMoPvXd/PkAruuWMOR78NzfJ7XFhf05MWGGZSan4BVNSnVv
DyuFI41GMXOYNx1Ute3ekP9I+yRx0mncj0aFtj8FDJK+OhVWV5KdNLX7rC2SMsFldwNNTh9wyynb
P72ewJRpX+e/q0IUGf+QMeXHU+poP/Jt28ZdQYzLgax4Lwh34EZGOTSFGssJrsl5/OihzHMhp7Bn
cSnh6/QiZ1FIJSb0694mUGRvBkbW4GvoTFIHkEp1TGs7p4fsxKg9RlNLmqai9cLCGpq2/Nh5nBEI
QlP9/+YRLrsujMTr3NccJ169B4TiIDMvb6mPTtMMJVmQepa6ymeoUSHIfoAxz+BMcMQUrnIm9NMR
9SH82da7B8o5AXAT0kNk4a8v3HevNQTfUg6dQznY6HYx+t48V5j9suiVOGhu9mWsoYp0X7Yw6s4W
vV6T3VM9l+PD0ENMmb/Ke1qyCiuCjPQXW3wZb+BNLU68LpHATUGj9lLAZ2vB5ZUv+vW+SQ0FTcH7
AGAtM02V1fKsKGRCagnKmFI2Jb5IbcKVQKOWjneB0Qp3TlAkF7OcGl2t1zk+AiHo9/+XjedRmRB0
82fn7FqF9uSVS8zNVmXWhZu6te0qT07fBT3s4fbmAJepfmBlZJvrUKl7O887/RB5sObZbnjGx0X0
pEg4Yp9x8EAxwwOHPwbV+f/IR8YRfeNT4sDw2uHY/3SIO0GN5KC0A6UyX5PBSGNzGTDTQ5+oQd59
BWv6VLN83r7uOUhG0P3O+RIt4uAYFrvDTGVB5+be+edBolprESJYwzOEsoTeSaAqSbUSH6OvCR3T
84gEHcwYTeKqRfTlP5w5HyTT+sTB8bdca26BSmGQQcqIF/YpDKS+sQurAFajKlgENdjT3IClyQgE
qcR6T7xkwpO5Qw0++lpV9uznXPxeQuwZrZdjLhLBaJmkoWmF9dh+rNoIOBT0r33Z77i6Sw1Uk/Hd
5r+s6LxUyXz+oQMpdl0Dy/fyXD1QDDKNOsfOdLr/vDhzgbVt+viOAshBeyz8lH0BHw2lpqF7aJzj
HeP+BGru460vSBpl4TWl1OkgMJUQHzrbZmq9WmQ49gfvpRuVwuPPL8rjRpEmc62uPz796GNqvn1W
ORa3buT+RTA7zYt40Ezro9xfHfV4Q2RuAzqglqls/79BLW7FHC209+N/QPgCBxpctmHXcDDm6bRA
cGnCOgchbsrf/lV4jrmKyEmim1yc1k0qi1GeF6h22Qv/BJ5ycPNJjP94IL0lDK0xEvYX27L5zj47
Zd2TzUs3J+T7rS2orspSd2lxIUN1HrMYTZYIml07R0mKeRpU6aqsqj3Tf4wmx3ddyzhtuJjB4m7w
qyt77rXsYeJa0ReskBEGw3VPgnCPiwtQDH6eGX/SbLVpVhaw5VDNbRq0JkQOntG3cYRGq6O2ftjz
rC/PRgY79/oq3U6K6Ed/beq4fQwlY48jlZg5vKylRncFUnPX23shRJAsytH22wj1T8MVqHvk98qj
S3YO+ZiEtA7abEx7g8OnPv7du5aSH6hharZ+a92nWvta6Z4Me3tbD2KTSLWN1j9n8TJe6IG8FWwp
jwWcL/QKgWqysbJNCz4ywEUOgpzkgb81y2reE1D0D5qDDmadSm5jwzWtv+JQ0qmaHl8Lorv3c6ev
3ouht8BZY//9P98Mrz/T32cjxrzhEDYAEu2aezXG/4XEx3t2gaY4rKcy0zgbUgrnbmrUxw444Ykm
vPpF/URAOEb8hLmkBZr9SMpfEbW/4HbUNfS3PHBvOPh3pyyShJi3GU8gVG4uvwbrgVPPxjUpSWro
qrsbFXN3fwCNGOp+uw7HF1jOA6A5zY2glKfTclvvSxusosqILjc9vqt3OlyG4gqNXAEJ/8RmRDVj
1PfH16OPQez0tGVLOAx6YqoLZuTOlcpXN0DmxRyj1e/4t0OKbRuu8RLzfY0GWy4b8eL8xIUrFhkV
LwfXtQc1MEhcr3FEKoNC/DSz3Ze/Xez+3Hykgx+eOPDI+KmuV4L59ZGNGzaFJ3nlOSlRk+QWPBPD
qHFlQyiZZItKH5VSdccKbcmeO6V1k0HxMBDuHLh7KOXxmbOJW8UHtCifO++2V5g6pDvfDSVAHw/v
F12PoxCwGinasCoNhgNJNaL6sddQBEMoy4uRc4t3mZipZUUgxm5qyvx5F+AeJEltgsw9cwiTlOj+
adapVDVgaaBNy5sdQlHHUNvUKeYZnHBYf8SYZYqhn177bI+eKnW+ypMW5uFc5Cki/4YabKVJzb6B
xH83cCy9JJDdPXBCmooNjYhU8igW1+2e8RsJocSUqpiGM5QZjKIGNWIQXmjGDnhrVKowT8CYyb43
aR0o9zz6DLSfrt7Gtq1CmPsqtZsrJ67sjntDrG6JESTSH2aDkLhxJsMfEVIWKKevrEK2Ggbc1zeY
1LFXmQ5Lhp6H+67q9XtOpqi6VgGg19Z2zZhB17iKwCFOpWVHH4N6RR85GDz8AGetdHe72kwkkW4+
Fip8SLsais0muQaqrt2xABs30ykPH9uudKNKgzOsP8O2pFgMG4Qeuz+m3vESswgIeCpkCU1lZk9r
ycw+xoKWXQsAf0ErX/clqztHIQ4LRMfYAaSR4n6GFx/nCRTalUXNzyxOQNClCWmjaDwqLoJqgc2n
w6/7TPIFTODY1SvLJ23Hk/hjhgK4kloq6Ys8wE7IQBUcbbHvsKEeQInZxXFUsmVnU49L0/+fTeSx
aoQyWy4FhTFIBsjJhcbk1+r8GdQQFgmObHALMXL6zk1VQE8cKKQthbn0ouZ1ehtKWUTq/DzNxdcZ
J0QgLITX8RolLSH9RV3RmWz8Gm14PrfGA8AQmFLQa7BKMoWK5GKC66bqN/UFj7wyEHD6eFTqTiXI
v/W0PL7muOeUN7dZPzxXZG89EHi4L0jX5Ah2S2sysv4MTiERflgUp1dyEnHTHZ7AGNKfmJpRsU1k
ePuqTuKTCtNu3jW8MbvNF+RroQtxlD+9Oklgldyj/TDU0AOlDXvneIqDQST4bVL3hhTC/OmHOen4
8Bz1m/SxOevbJ1uetSGfgY4T7/y+l5KRNSRqPLHOkl+uJh7wm39V6VDDXJOBzgrtt1tNbtYh7POS
fB2gppTQLfv7hLmyZq/b7aQDIXy4CaMQtEtrjtFcIUyVEzlgsf6Fdq0x7nS9GHf1JOcbA9PELKtO
D5kq7np9kDWSLuxNuAAJnI7DG+2HZ6dpi9DI1FNJoifttLhMiuZVpYWQBvqhkbIc1i7/P6Ij8Y8M
wBh8t7NmFdQy5nlFNCABZ5ZUAzHtWaWMxyD66KCQHlKpM3aYE9E3b2J1uAEVhDb+o3iJdP3646aZ
VrygFszu/dbNFNMmqR6wXXNS+d8mYMVxCIX1R85rJh9LyHChkf4CLrgSYF2Bn7c7naihqU8E+N1H
Px6OmO3DLSVyh09o2QCKzhnqP9AzlDgU1FRg22yKt2KKDBP32bBM6xM7NAnaF0tyWBiFPfxrhkYk
ELzuobQVXXfVPqOzcsinsTbSWYlVhXdewIIqqXcWm8ijzIKDuCOOd0vjMLYX6oeM53J5QVs9P5DI
I394bouHA8D7z0H4j3Opjt6EdhmTZGGcPXcX81oCi6dsBlg6ze+hgbhaN1COa2PKn7AWOC0Ma3UJ
6Xp+dT9jtjKhh3nDB4cxQVV6TqyyQ9REmC/B6uTqgksrqSd3dTxk7XfTZ0ZZRkFo0p/c4jBOWJcs
q6Y00lhNvvyyki9sLKJjwuhB5ermll2FC6A7KkspDGrJaXUD81lAt/p5kNU3icwmqHPW+Fc5pz/U
2OAo9iL6Rz0X/R9rO3cL0cIxtpan9N72sstwcjQ57+CsbmT9bAPQDvYs/Z/gdHsd3/LSHlTxVD1g
XfWl5LGD7NAwikJ2sOwb1yIHoBgy9aCGohu4d9wIzIUYnP8gdu2tb8FmWMMm/ctYIJJBfn/IybXY
7Q6Q7Z3Ej5/kB2BDA60bzWR0uqAJ/IysMD1SPuGaknKZgmBRwDM7fHF+C6m+9d930uHgOv3/AZdi
DD+ZHLjikiQs/6lqvG/rtaqESOoDBV7ro4IZdsBsntte+yZ7s2hdZTisDUMkaUv7GLdNrYggmj1v
ELyAOJWFYqjQXA2qo79VBLsEU12dYGfApULs1dDVEHZ27Sf6eee4PWv0QKwRcIh6/hd/5CrmerW2
hdB+5acMFyyOkQgPL5qQQxZSDABm9xtkVeX6pZlis6EnSAU41H1v4CGC7U9/S9lDOqkYuz33l5V0
75A2o/IcXf4PXhYEPmvHwz1fTYC7GZB0wQPOExBRhPioXtY71Gnrek5cDOXTO6CRjuqrHOunY8z1
Js8uVYx3J1/8D1331wOGmq+9hlnfOoI6/L4cwgT+0Hs8ccL2P+Ge0eZhtCkIMfPD5Zvlt5LChY9c
riI2UsqPr53pO58tK9NY7/PHNR/U0gXz3GM0NVXmHkGgk4serqCebHbEuvyB9sh3a8aeJ9pBQHcp
3dJhe2QmlY3rW+AQ06zZWzGTY5bYSHxJ43MeoW2KH7zjvjBu+7xfQL7scdoUxawTAI/69u8GEN2l
OSAPbC/EhIfyaV+HwhLaJM9Wa9GAp7p7BcJSR4jM1M+bKa2hW7y9wJ5IzD7JRxS2T4644mdrWMjQ
+8Uf8IlNX+YCE3C5sAYPLmgPSqOntFhbV6F+5WsK/1HbCtTtAuOXAPTBII3TjayuWH5c3tWcohxm
6xPdIWriNFWLOIzFB/U0TRnNYAWX1v/Iv9tfrPaH6zX4X2rTvqyGiCqboxBPXeokLn4l4MqZrkQW
3ZLZW47T9MBZ2vdYBeAzaKjPD8aer12j+I7YjqNYyjvYXlp5FexPXalQRdC/aJeM2fEzSq80AK2o
e3ca3KEEJlFFi62QrOIosdTuHSoET272EO7BIowm+sdRyHbwnmbUvODxujrnMV+2RKdcCKbjjZ1I
+4CRKN4Lj6kPzkDTE7zUgZszV+b1zoYw3ynvObyAKoFWrZyhblPtw20t8T6BaRZZc3K+AN7GO/Hq
5CLz6b8viIu030a9MsqS8kj0uYAuKD2IZZQkJoHZ48Aw4CMoa5M3SBwbUHq25zfR59QzVnVZrjnv
hqIxe5Yxwrmn+u7bB4rSVsdaTdvz1IB+EznaD8G/VjcakXptg8smN5Z4smH/G9jn9ONRzVwEiCK/
poKaojTOgtdNrdc5m7TcHWkUhGbNLYdvU4PEOPiYH6kSdJMVVcDjIpY5fCAe3Vzcl82seN9ZcKsO
16aRn8lK7+gWCmP2pl+G29dUQDXok/b1QK9FrPqpd6rmCx7qCUWcHTbdBjcfbhjn9Gr+yxZbHClo
hurezCVvE1PVSZ/4MO7sgCQfJB2TTsMPuujkXBFYCO4h7niVsD7QkwXG/BzcgoBdaHSMDWGoAw5L
R6i3UnLbEHTHKiRJKaoujPGAHp+OohAD9pfizFMBdPbZAqulmsjAogJSz/QItH+Uw1n9+cql50yQ
JQRQZB9SwIhC+PWNN720JUiWjSSxB4PAtnp+fdZUa2HbsicSRBl0kfCZ8dPIpmBfZMPp4BZZULEN
GF65FtO+HwhZm799BvXLkWRXc8alzlY5SWmpnlgKU5IfnvN9yCR39RaiHFfsSumfCr1Azf7DqBwy
/tRTjmjqcdfbnmxsrf3YGvttzmHh6gqjZ/er3hNgwbaPLGDS7UxHVtdjNXplXEoeAbbV1t+brHPU
+1R4xaIAY+UTELEoWCaAhQHSiaNk8t2wMhFkHGrY2goBNRO3TiX2tmzZ7D2sJFHjtE0+iz+a2sw1
F8ZYDhiVAOrRx8KKEC4Z/dy0uiTOc8Q7HO8lm++IB4RjoIVTiNhaGJBuq8g2fOncFHAwcpnQpXhH
3BwnlJBE6YN51JCWmk5e63OhoFp8Bd6jUkIX1X808C9P2JBVij1QPusawzM8gFJ7Yz3lk+aLYlEo
NT4i6WnC9QUXf4gin6Rr+pp4se5jANMMVR4szTkf3K9cv8PCTzSaw+X/kSPwtd2ZIT3blA/ziZYS
4nDVUBAwwIg8d+9ysjUPTHFL2ict8ib0HlUdnHxHgq6AktXNYseXmUea69j4G3j8MOSjZ9zuJyAU
ac0J+Jv4yMdExeQT8d0mlW3RqO1apiweJ1M50IUpAjMvIURyvf6IziWgG1z+L2bXuES5+HSS47Pa
/6iEZy4aKY+C6DBuVXmcnaWa+C5JO2JugZtpI5hx2OrPEwqciduC2KyG7xQKln5z9GmIM868ghJw
guAukA5WhF1JctvMB+P9ilKfm5I+foUxLL2KGzXmGGg3D0ZOS0NlazVtsTEWAHKEFNIsSXFjUgCE
DkmxOz2zr3qnzQFhF+w45MYo3C+/lcKMWEOzeKMH3SlWMTYXCArhQVTrNME395+A/uQLYfrRxtPS
s/W67QhAQvNwz0F50ezzEJujeeQhNKmmtmcPBtJxfEpVAjU3NdiRLkRSwdXeJgz9oI0hJLC2SdO4
XdG/+191CXmSfq/vGpvhEbvqBGp/4OGgYdV6gxUT9+x5hytzlcPla1TTzi3h10Nst629FgOXKXnl
jpWGSa42thEoyKR7QU6lFIL0ZtB1Gk1IdAtWs6hy4BemPQFCg17NxbxNPy/tGfyA3LksvwIaouYy
aC28aCQvuOIjxm9kgqoFutIqaZ9t1tFU7pR9MH/V2VqYZ481h8naS3HA9XCcIrNOnvjdnGUenfyB
d3icYKmwjRSPLZKRR26RDBzffpzS4m2nc6cYFFqr8pNFYsujVtW2X/QgTr6BiHYI7SrbH3j0zPLS
h/AfumBmkE556i60jzyLV6JlnBz7RnAwKwvM6qQVSI0TsUNqKgk/uM1o/5QOw7O/1D0DgTcy825+
I9nUc1aW016JvdfKZ0KHoBuww+rXjqbrEAXd8rrGoKSr2pF+AUNJHpLVOFMXXxILKcvCEIRaHSUM
5YjPwluq9a5I4XPapB9ILyML2NfeOZO7/xyqLBr8eoGU3MnflR8MzXuiP3kN1Jv8n7Qp7Yi44rud
Pp459E2BcAoEX2/iU16fzu57Os0j46Hq3XB6dGrO9PV5tDMkAU8MsUnJ7IqsDrvwID/WktVaN7tU
ootrZ1uJ63FY93hxB/A9/M04E3TMAubRvYaNDWHhndQhi5QYHdaLsVvg56bGzWDgihjmvbw+1P3h
879rs8RJ3MJhBAOvejoMqfrJqTHoEr0aXWWfOzdLr79z6qPbIsp9rCy5QpuAYbQfYVhY2Ea0m2zb
4oEMaTjv2syE0Auhfu3hXpC6j7B6YXCXo1p27nl+xbPFPAZOqKUtK0s/33TIFl43td/vEQfghmYm
IVmWTBQtkukPXHeWL4tRzePQOVNfykdfG2BaXjT/pWLVuLsE/cUQJ1SKZMbzumV842+TAl1RBpyd
leid/tHnicMOnjPhJQz6pFSv3ivh+D4tg2A73KkuoPwNRS3xBJUi4tSjAertfCdIq17SUbLPGDH7
uLGRZ6pVrKBLD8vjk+xXPpFzNt+HkIhgo61tGMWXMOOtr0Y3UVrqgN87f/jRPzD+1Ae8Nst8C4IJ
1yckLiJuXxGcUNeTLnpLtsZd2LILo/p0j0BGh+L54L0uZ2Rjn819abpi5M0tf5uqzp4h1HuFpvfH
Te1RkUXksvMrqCgBR/bm17jyEFNrNQDS17GYbdb175zY65ULyjGKTzuWES7PDtt9XowIUgpkAjOw
XGnoT+DOl2srd4VoHG9m9MTHp1YaBXEWeYwhp+e27cSpsxfnh3Ql7jImu+IGIgynDE2Hg2Tt8ofH
muC1xvh6JnrcaSH76omtIUdVV0+Z0Xahah5QDBj6w7jFCRuADxNujCtE9qy47PafFknIqVBI+PZa
NlR8GBa7nl02nyjQcJrH8Q0qyZOPRz0kR0Vifab7G+6LJT6qiTLkklIzrG5k5v6N6aQKIYJMaJL9
a5Nk3NieqP2fBKcaMIcTkeFg3Djt4GIysjh2ETapwdRdHpQmJsrgPksTyGx9mxj7NqVoOESyvJ2o
O2F3VuuhGXnboFAAQSvl+Wm6Csjm1glIULWbCw6P5yJReOOhgLmQGrnU34MswXPzlHe9o49IfSjw
1MybWLOw3/Kc3erV7m87usFjD7+nwLr9w9vltUk/SIEdV/4rcsheoXHqmXOSfYDZA0y4okNNS60p
d2Ll7sWWuZNIaWJnUHtjDjHm2XwzXJI1vS36VbAo/DfdS6nc4DIxVFWVVNz5EHoEtcTU0SV9t1/5
glLQlKnzsXJ4KyL4a5Sfq/mqSgNRDv718bbaMIcpuzAOTskukpvUaQ90Vv2zB5KJzFbi5t8Tf8Mi
IxilO7vnQXe3cVLTAvk5/fXeC9BFGNoAdQ4e5gHL/oJVeN9/6cgfSbt+ctX2q6gFALWi4fc4yvqo
hxbZ4EIPHD9xSnDUwEWN7frZPXzJ0tc6AKi3sE2bqWNBABajxn5qGDTVuYX1+sm3HFrjowZNQoP+
wu6youX7JJXZhDhBGPLK8IQ3QZFm/RGNTknt8WP4yC72o1TMt3VjWCLJR9t0TB4Ymk9EAGQx+n/9
qa+kJSDNk7iaIfDpr1lW8R0gIHZpq9mzxE4B4+NwCu3NCy8XpfNr0sYLQsIylidHa/2IIvWTJUeW
ILlfTqPJzculnXwitpSHlHRMs3DfJW4N0aO3KI0cD7wrayVvUgdf4jofk2YtxWdq5YSlLD9q15gt
42jmXEkgS8g+pSpeCo9PCtzBHr0Yr9s5jrKXC0IDY9sX+kFkqTOqmXyaoyGi71VdG9w3infua+58
k4uY3O3pT5eVInUiOgWRgOzfGyLrKYeL8Y6X4/Y6BonL38jkf2lfaG8f4MFvwsg9jkuIDU2jmkkM
9sQPR08tJcwBBVuVPYRLevO9Hpq8it2Ko4f7IPnrjfehr0DaphfaDhLDnGCc6vDhPvCn0l5fDoog
gCmsLtxh8O6YJbNoR0Xd7SLRv4+4Cuzyt12EXC56sMVsw7C46ZEtTYui1AxTS0qgbXbjh+u3wxN5
cnC2Xt9Yt87qzxFh0m/2tea5SvrKgMJtnelg0XfN5ghBs07usQjlIZXLp8GSo2lqAC0wQv/0ycIB
dfD/Jmr8Fdwz6KwMTu/9llu0CRlrEkNYuF46bo8wECLBNHJhYvVt05cYJllIQ7lKRFl5fT/YqoeZ
uK8QvWGj5fcBRFbf7uEOBiX9+fjVKdsKL92/FX12+hnZM65HPBqm5GUQsz8PLYBdTwexOWimkv+j
ax1VSDDEib5AiaJOZH2EGb4AscywUZU1NmI0Tw7KgvbCzGevBO/4q8E6mAjDK50NYfmjLmoEl0kO
L5EXj3Yi9YQJ3HP8nxnO9MsVHHffjb8bNwXlDvOtgKqMQ1zfSfri/lleBhfQGf56Y3YxAnhF5Y2H
EGfaVxMhBHt4E0XTBzqtxqMDGFvMkao3bQwX6z7ICteTk1+0VLOcK7hKdQDrFsovK3LR5oFOtB45
/8MJMJsDQ5cxzFV3VKoK5I+66S4z9UuZuHcgCk1BqIdgvrLpdNZ+39s3Pe8C6uf1t+43KPDZ2gW0
9CZJnlHF+C1cfUJ8v18ZPNox6vJ0YpIOB0qataLgzFX/2LeK9dXSWuwAoYnQFXMgouQskkmEFlQj
yzZTiCxDQEo8yjIQdYRv5JJB90ZRzmVafwDAPVHev4DXlas4m6VzXCExsoD7qw14T8CNwPkVKOv7
/tL5jASTGpnCcDN9UqNNYtUvBfQUITdtgQhTt6WK9hfYgxYOcb4V9v7jVhvq2p6WDG889xSHaFkb
o03JjNxjWb4WmQH9iBaUhk5r84EKo4TWcPsA1DNlyDcIaWUrCndh1KLa7uXw6zKNzkJM1KfnVPli
ihl5tqXjoPR20qQqZVZTLW1Hg89JStRWc8KwKXpYFbae17kJs4YD7zUOQatJJP49BE3hT/kh+Vyk
lPOqf3bfy3TChwaC1Onl3TiHX3UC2tHvifMX19lHXkJ8hkrC8Q6HoyezZ8jn/ckwJFFNDvQB8YwL
h9U8d9uqbWpcRC9/RiUbzfj13qqKlmkLUJKF1ViNRcj2RVwsws2jkr89JldEpbel0St6p5mtuTkN
d4DSCQwt9bFybUU4jigqeT2x2PsNUSqiFhsRckw8ReQjpMagXhclb8dMHDdCLWE4ljrYLeV/mVbU
3aH3d9hV8Sn0fJz6YgPUcBuvgS/0spS3A3PSggYvcdalfyqDyRJrr/0Yex53fgPs0pj4c1EnenlT
UMWW8Mh+2ltFnGc4URnKidNfY5mA5SZ1S9YoavafKq+iDJ1a1ptwwwH9wG7HYQ05aNU162i2WGcp
LvbAa7fkwdfVUW1jBm8PdhxP9T2FbHDe3pFI+hMH09iigxS25njBRKW1q4BOeqSRIfKqFEtvg4jv
5T100/M4ROGn331GA8GzIVLp/SsazLEHooCMrksLHKPB7Dy7TS46bzyemZyRTv3SgxtJ4Y7hDybO
XlVejN7mAAX9Mbt6zanTb2iYd+1eVpXGOxIuJGNEGRVG870TvoBLs4chO3ZuZhxMX8MDCaA2yiRj
veCkS83cm0gVBHrp9FHG+l/R92irIaNyF4FXANG65UPtxf6VBvv0nc4XixTQIgJi36F/pt1xb/vb
qAMr5Uvr2DGN+4lLsZ++VB+Qgz4o6rP6XTbfMX+MCg2sUBx7eqvlJrKbwCpIMvmCjHtn2Lr293XA
DlgH/mNhzIhxUdI2gGMDhHa+fHCGvdQq4nODKXfBy+e7UAmsCaowF9Ry8cu4MAcjLWNiLdUXfmqr
YOPiYZSqWkW6dAix6TrVmfJKg1WToGkEE932X8GMgVGd+C1/QLMUmQKqRUC3+d+ndU+WZ1cUC/pM
qHz4WZtZHphcHyfKObwk2GJlZRoEcVvEr4Bh/Uigji3OYK609MnLkZd1gJyg6R602jkvTd4j5Sbm
oKM3vZKo70YfSb4WRE4XzKGPOyhfOUM/Fq+T5XxmrezKWdbear3tI3LrdcsS435Ju1aw5VR/p7jh
7AcXdvZDIsOem1XZLnixrGKqkGQrD9JvaUTvPJxSDCriu+v+c3Dg3PMNuBwdv0XN9DkDAFCJHn7Q
vfQrb3N9LlbSRyehWMAWPLCsCZjAPx5+05u7m/IWbfcd4L3tx7yAIqYHeMx6AXVwb2KyVIYimy/n
d7qd22cKKK3ntMPFePNZq3NJGhXh6PYPiVk7Zok729xmxVIk39N5PAMHiSwgp5wdrh15NS3ovUoM
7A1Z1POyn3j5hdN9go/H/RaAdWVCR+8z0ttGdhbbzBsMkwYn+phgWtPmre958giqjitFYfgmFpQy
CGhzRGhCUrDEhq02pwXAGiuMFwwdTvIUXBeoWamsvD91CbCZ32k6E6uIDPYeHlQPQJkYGIf70t9T
GyN1Ued95uQ3KJ7NICqDDbRlxNYWDgLe9W9EHjBIQOn0gbWerec5lBj0wKIzAjalshzkDi4cv3vF
2IaYjVxxA65Gqtg51i/VOPlHBWdY5ZKnRnMYygqE6s/hafBZrZQUk5BwJRu/SrP1Ph23xaPU00B0
J3LEhGPc3bv4/vr5lArvMS/xCl5/0nIrmr8hNWsUwjwAxAfEPgpW6lZknRdTvNj4qJtcVCuV+dKk
7v6DxbrUuWpFAxR/dPH1WFK7bT1xCY0Rq4ZuLiE9Ai5aHCZmu30JtcZI2l70xj05FYd9s6cQhyFk
vWjQVa3WkeWfKA6zAnpRi8bqcLTfUUe25BMOLVCDAMZhLWmzdMfsKKvA9lcKBoIGcHQQAz0SeuDG
Dx76AWk/ivODSqO9HsM6H+UYML6lHrn7dGB4yuxnSqglXYc9gRprXG6POEhrXh4ChMkomAF340EV
7h+jPfGXcOyuypJmGctDSjcH8P8jhi29KWeEy5up3kN7MG2TDgnvKzKvbOeZuCTb2b2mPTYiCOE+
kkM4MP4o+yuveGVOZMBTFi+w6MZjKiup6HH5e1l1YT7CKhyfU/JLuEPLMCq2DopBq82dvs+rezhy
HPiJsJWJj1rybc4wdqJhN0A5ll1EJ58n2AgBcKaVviCnmuWHTEcxfHpF2AE/u1L4ST1U6PCaJvyw
ANKIz8zr0n8EY9TU4/RS/S9QTSMqpxIiu/mnnDQiSkZgRrwxQb0bxUcDU+k+Z/zPHb4TrNvX/TIq
kBsbLVSwk8nVPJls9/rAUt0pKCXCDl7S7c/ISGPrKbEQvZPz1/3mkWrqMeblU+GbV/g94g03MGmt
nEEDi4UqTsl7zE1/+QM7gZbVN2xqiyfM5c3anIOVOFCAP4WRgQC0Jv8GT+7jOFtk2sdvWzi43YUp
fEEYZA7y0PWxI/FfbBxDqzOT234mycNOrYU2bO2rIDQtvPGI6WySecOeyKQBLfcVCUIugx36VqsR
Y95/IbmfjB5vHLHy9pO0CDkaDrOWbOzS9G3qI7GxE/9aYSxaiTggcvKX831PN725yVbhw2g8m7zC
0Gdj4Piakzds1bf5fYBWtB0ZLA3X2PHVQ3l3n/nbo/hdLEnPiSayeDPQI3JAyReq4/JxPFvNpDFh
m4twBVKTWKwjFxwAvPM/UfufNZJoZb6D+3Qou37N1Gv4Gr7eQFAjJ1mD0vbQrq0jNwatk7iVXiLV
xWPn4I0lPgeZ+zPZLTi4M7M64zpne69aRxPMedJJoI06GBmBpCKWqDGDhNMLnB/F5qyrBuLI0Zd8
oi6VxDOUTd/zCVlEgfbiVqQqjBD89FOrlJxbRnbz8R6/cHwu176UEaEgVBC4NqzSxfBOmndBMv0e
KTjkaTPzdwLmGZqq6ThN0j8M77MXqQk7STfxwLvXmdGLRDvU+S5Wr1AW96+KvjQ9+Iwj+tpP4Rjw
GvzKC+tp/iJB7QLILqCbYOt9m5MgeFhKKtfvvPargDsabZr9yaBxzaoXo95djZjr+g3Us9IfuF1S
3gwLqHoZy6Mm3xDq4rgvMhlG/Q/ZDPT+KFX8exM+7R8dUHMWSXdK7htye9l1XDqr2H8IBUSToNRX
2txhmggTFgm273lm14YjTJqalqV7KHfq0Fxybcw1I2jmT6fbLomsnL31tQZI+d/14UQwg89b3CbT
jKm1b+zJvYbg2seDPPwrOxUWFSgoZwbhZMbJ7tZ6wWwR7as5PZkGm3D7jKz+JCoRLd8xQ7AaYml7
ZnCeFhwLfsE25PuWkjvgm8+/aAJIT5dmx/dLGXg16m+pJNT6+UOR5U6YXGyQgaEZfouTFaH5uKLu
Drue5nFgadog6FCcB3N8aj9JefbHNOu901mPZUkZcmTK7QOiqu/8Or179AcpxWe3Yv3tf7ZOtc8L
dkzVrXlcNG5s20fmxCCVuOSGHXioflpWb/tNMwDND0OXTaxaQG1aepti/WigXBbLRbiNi4yKBOa4
KUBVs+cHpkotoF9AY7Tnreu21l0MhxzG2H0rhnCT2Dr3YqnseUe9WZ7T/ETh58r2eoHGu1yom2a1
XVEi/7jQxzMeqTOcapDLuy0OyPVXLGHPRXWAw0n8T/nk90dSIuoar9U/tS27c9wWNmm7jVUom7mx
40CS1U++WnTmUm73QefHJKqAotE9KM45ZHtoqJ9fLxXmF9CJ34+tykNer6FAQuYUSuYQT0D1RB7+
2UYu97h7Uk1QyKyVswc1fANYJ/rPWT3KDHH556QCdIFRGVRhWpC7v9zMWlEGyx6jj1lrNQW/u4Im
5LgZgo841CkOUGFcz2UHUwakWalPtsW0ryQZ3y1gHxD+qcBdk9KhzSF1RfA63r0qHAy/cLoPKSYQ
2vRj4pyNADZiPcTy10M8qmHJMsQJpUekXAUKStZGRAiY6+UUKQ6PEXOjKAwfsU37b+7gKR5LIOOC
sihs4tyIE5zwCS43RSlT1QQZoCOgYo7Z+bCvRcqaOohNtAUW0xlJERF33W38jSV/chMKVIppNSWo
fPGu/wKqxRHLPkW7lDXij0yqRccoxvACPCzMLUp0ktNIxTxIfF58FH/H8+0fb4uzajEWKxxDVmGt
JzomNcPoyaGuej7TSESWK/88Q6lqmVy5UdFmyJrXK7Z5HqD4RHLs7ipArgCxOdPwiQBkJAhyMKlj
CdInpylKriICZvIfF2HuZa34eDr2kgs3Dqbu+Oo5gNrl4uoyRKPmp0rzygCDYzO8Uq+WLD3E/45O
AuO/n0l/5BoBTadzedu7gLbg3GC2CfhDUUQZSGWJgdwjASwrPWiW0gU05EMgS6GBdD+wTn9tDu9/
jS/30XL+zpqPkkYzMY7Ep58E0+u61Vwsd4zVtUjX9o+hR4rWL0mJyxoFq1YziKGBC3UiodEwqWPl
5+zFVwYAYzpnnwgJxAy3R5xr+3co7pEFmWypwg4wUEtGlwjED9WcuV1bN+95SnVxGAUJ4th0za0Y
LaY2HmiE+pCKR2754QnkjjP9rrXvCsWt+3SHD0pc8681KbrCFxt0gaVwuOH22Q+AOFbatYpxyICP
wn5pKRApyEhG8CGwVEDxurNznGTDwjpkvdOgsYdRNdThHGuCl5dF6+pH6cWD4uWjDE0wOWdSROE5
IiQ+WeLpk3pf8RJZ1DakunYoX5NrRtKLvrsw+I6L0AN6nzJQeOojTh19y4munGXFkTPIPCnRLiw6
RC/eCTD/QbrB4FUVMAuTmd1OxQN+ljbGwYlWAiT5cKLXYbkfvPomPyu2TB46z05uWJ3WSILI2kxI
RL4wSdDT81CIZpau9J/c84OzL+UgrXId6Sc1OxgS599WJJtflDnaMFcX+kHoBvnNTVoJO+8XE5/V
/ITUFs0kHbeff+rTopj/nNN85X72PfjNQul3qXBt2Q0vbX67jZPakwTTMgoY/+AQG4bvFZolRSUE
EUrrMbTYZWvnku9UrYzURflQn5Cqjxpx7hYzVNNrf6LeqxJzyvd8QB5HT6WhyoXdt7HK05s6Lvy/
DkvYKayZ7kox7R4QPE2ZALp2j6S69rfAHONDm9lb1gv3QmvSJZtBtqzQm+VTuJ/s77JQq4b5c+fC
ymVzOs3mYUs0WrJm0bTa7QuJLOCa2czgDmAse01Xdnkxnw77hieguf3OrR98C4iYYNcR7enp9t/h
fh1eh/a+E7zSJpSkBxaSuegajdA8VRxti+swoQQW+ZcRdNEebULHTloRxVal49y3C1oJbFlFC5i5
BCUCsJ/sJXq0CPrLIvQ6fSt8TNK3ZayUskterA4KkjQMp0Yxmv+FCtKejDGig2kqzzUkvwfgr+eW
I/FWQt59WVI/gnkWJ0KCA0leTVkRzYKttMla7hxo9e/MxrtWGQ0UuTwrVptL/IVi6KRdAYjiJSMD
IV8Ri2g4OA+u2cnDZWoO/3hT2Q9D1Qwn8h8R1sxGf28d4JjlCIzLnzNFAfcpiGM3DCBasEYVPpKU
l2YX+TopNsjFbAOSjlsx0SiQ2b8tFqTLiKelbfT5yYJTVuP0Knb6JBSTJdSfy5IcvVu92BwgFav8
Lec5tyMDyC7qk68Wt3B+Rctc4Y1tGgVQ7efqHMyMTJOIKiv8f0s4okLw+4xR9FPlLAfhvnYIFqpj
S7w1w7SH978dEvfb78RBCr5b9oZevxpvGxB35jQORGUDTQY/Kq0wMHQir1Pk33oW0XFZs1OzLbgV
BEneDdooyN/baBsFXYL5FESiqPLuElcq3IQ+mVvB+Fnx7N3JzvsEXF7rY9oshp8mAZ3G/mTVmTQZ
wvvesj8CV7MVst07TjR3uwnv6el36JUy7cyUI3OUXdk//Ivn1GkmvUkm5cuAF7Kl1R/Ueojt88Zz
UNaq1rGTkuWxOM0JSsOXRD7FkAXSa8K7pWzdhybUAWxdvZxWucOperChwWTomGYdFchy1MxxKR18
3yGvPnonjrAKu4Seqb86+au4W1x9JaEa+bxzn+kMGtAPxkh+Sx3Vw00AIhgNWv3Y2LTKXQ/bSW2C
cK5kyVlXd8cjiEOVk0FZ/v9Q2PkHP7uQfzrMG16/TFccBIetzH8eCNnAfwa8/RehvgX8KlfwaKTL
8SlX9yrU/tTzbRneLYZlwjZdmxD5jlxWgc5gqeMbYTxoqWP+Bu5Au3tNNfMFun50kZikaWgJMeyo
Vw+h2tddgCbOVqMeSC+/cngG83vKNSO4vrz3bf37ZlSm3T52zJzUcb1ddXLlmEtyMJkZBqoPWbIM
ReVEzC9FktikdWkXaU9lae0R09tr30CeYI4INayY547y+1jVdgLK0wM7fDeEcHg+qkO1pAjA2M73
XfwBdTtIucQYZkJCh1bfllyXBJaBNqN5xmYEl0M/jgdYQFQUq/yesGb8wujRYNaosiyR4PUk84yr
48wY0bacWehhgCGmrQ0DTB5BI56ba1fHpjZoVbYlETJnkaW3llqm5pUqlbbvowyPngBq34T18MhZ
pv3sDOZb1FFKWfdCm+QQqMznyDVx9crCydpCqEpfbHcwpwhQw6LT4HF3ObcMX0ubf9Flz8OheAtq
PBfKnM6rdgBozuZ6N+U5IgfqWqeQvdM0KwKRorQc6N5hWZk/ix3eRAPFjtTUGwSt3QzhCXYLjk+5
R4za0dnyWCSYKSFjzVdUK8UVlkCWmdZrPPi9tCL85PO+VLOw/FmiPbpV5YVEhm0rezB5Nffj6a2P
Kx26tn2gDz5hhJa4bLfrKQleIvPsv1xS63IRLNIEgvMliAR7dA606gCYegW0KlmEavE2Pd91DrAY
EY1B4sL7/A3vS4BVhUSjem6CrTUZspWghhMEpxJ8RU2feEHMBELETfLkuHQMX7hb4H13rcun7Ehm
4TwzCy3mhs2Qz9dcCOEe7lqpa9eNyBBv6dgTeRChZPjn1+nS6w8t2icn3oCqv9W+y8BK7SxB1zvi
FaYxCElvMHj0vRX15a/ZVeut6ii4ynTaBoutZKLj2nZJtnpPV5dKXWhqv6+xKG/ExhshhN1SilIV
Cm1cXJaHvdN9yBLtdXBzqcVOgVtA1/zfUyjKme+eVec8aSYzEhUGtBysvG7lyFlN8L/NabcbKHR9
hl2twwX6kta4Au8OuG2gtUAlsuM92TE2fvYV0V3pYcmxPjWC4QZs+FB/eZtyKanW5L/uQSCVV5bA
WYZySiBqgN9ZWROn//3WhI1Ns8SEnSeY317sGgl3WAKw65/YHgpU11cW0fDpQUCwxg3aEPLiFzmS
YESo+Wk4ankXXlAQmvwIUd7e8oPULiSgcNePTw9QzFu40YnK915kDmJYycsw1iVEO3bJZvMqUie7
dvrYhE5aMZ/QCEUgmHBxzBxozJdMuZ4WWmsJJZNfgh9BXy23qS9cH/x0/tBkrdPLhAd+a2QhtphY
fPRWWNLP0t06eoWZ4wTpaoqCzG+ja2GtgnJVS9YKuhkDf2GSz96ouvC1VzmzhBRF4FQH+obcWejv
yUihKNe19CHmBF0l81PbI6B9BOIC3dF+Z8J8bAgDPhAK177Ceqn4TQuxqoYfpIed1/hLo/Ph205o
YAB87gIEs4KSFWF65OxSyPTH7uWsasxr+PdAJgVCuDI7g6jn/fjW3FhxYE2aJc4cuFG/j9Vvj7Sx
kyGqjaHjfilXoY/5shtYxbnBZAJQ0jVMygrq1vjA7DvHsN6qPUsGUY8RRj8IQPXBb7HHj7rOkZws
gqIP971ItrxHCbkcv9D5JuCyjH5C3vYNZFlg2XSOJ7FPHVPoRiW0Uya17AylJW4cZ2MiHpobgmiA
tHjAJd5d15sD4BNjQjftU0Sdu8+mLrJftwLh2q7dTUH//An+3UmM8DS7nOJySFq6zdWerUd7TH04
R7cjkySZoqThbx4Elxf0Thv1wlo3cg0Q9J9xTlR4n2ZXNwocG4ESlg4gT+gMdo4Pa3Lcjw1hDZ0s
zMorUX0pgUdf9iQ7xfPWTqngyn/1LftAK0SKFun9/98Zr/5yKYRVklkj1z+xKBJVXtd0/RDDOv1T
0/VOPaZvOXWDuGxStafMppbaS6ogLCzS67ICQn5rJY8qqa+h5dtCzsp06mJOk7x+a2VPGon+5Gx/
NwqJqbryMYDuU6OI7szQhnXlVE9UOadbWTM62Y9gB8baKiol9aQ1ZiHxLo/MY2z9Xub24C0bxgOW
QtUlnAUgN6c9I8IaDTp6j8JqnGIAa6EIr5g+nHQNJttRIxFS7ORzQlfmPpKVCDcTU626bsNHOruG
4bNJW/KrrksVaNlvXVdDWFRlwDvBLYZjfHFIEhTALRU3kj7y0AwaAnj8lz0EKNAhYPrVDIwjwC5Z
C4my1FP/kbqHEy2975gKE5Plpf4YHNiCVi5fjV7MPfjHDA4MzpKFJdK9WRVLgtJRej9wwaGG8Fwl
T7XtaA1teRlAUpCF6gSEbmHLA+3p3fL9FeJWhGEVUDpdGcwHHPkPXmid7Vae0mMdJVf8vv0xgHHR
ASvCdLIq2B/nmS4yNpEznG75HvhXkSeZKXAZXCZ9Hl3s4BWJLIEliYcsAqjfXSPpQWLYgDmFHBGd
gJ3gvXwzQWjwzpJaW20Yiu5Z1z48DPdGCWnMWJXgZh/CLAAZuKEdFHzGUDQdaHElpxzOpqHAn2H8
erq2YHWSLucu7CnMO9DbcrBs5gAh/Ffc7YbpCuA8KTqqV+p2Y83tgLwAgY0cTRBpzd5MuZdDMnY6
ic1eRPoCQimabMw2iNlN4IkZjVDCU1uC4zR5CzQrAVwwHBhK4nJnveEIFOHNYKUe5wkDNzraT6Rq
R93x1JiteWcc0+G892EkWDyhRR9NhjyFAuJ4ejMDxwF/cH4PIP4umg6Kp1j7dh+NbcXFSg7bmJjW
qdinHhoQeh+XyxBiFHPBcelnh4MEsJ7CeCPOY7ToQY1OmASUslZFHJ8/fOv6asF7uNMTMs15CDeS
bZfCmWLMUwttwFgbrIbQN+w6FA5PrOgjMenW2GdicGMuQuOCJDYhaYR2ONMn6bO1F29DYPeOZSxM
jDLMqYCGJW5nOQ6RVt4YHr4mJodBT7qoQqgI8FwGwobCeAPdisMk1R0VtPaso4DFMucOqThUoUNJ
Wn85Gg/IEZcHdSRvHwrRSEpx4A1/vgl2I82K11LaZHyOLQRBI3QZyhXwJxXsug8agg7Vx8/Sc2Md
6rtTrFH32Oglb1bKlzd595As156dcEAw8t3FWZ1lO7jukSy9/PL1cE1sZxX4b2PzxVJnNx7Jn3IU
pho5jmlg9Y/CwUGWgrEFbnA338W2A6uBcvnGtAV71Mymv4E4S66oeFzYMfSPnVgXD3FQT70Q+v1e
lKSVn+yJdYuLLkbsTYa1R0NWhPreufMAm6/xF2Lj3edPQFpVZkOs3Um8IQlwvqjUuz/1y5k1xL9G
OGIcbnhOUMvviVCfkWcCb24Y9U4Xj90Yz7LUJCsscrlO2ltsJhCmBTTrBv02T5GaWC+/ImTiTITt
uNTPJyfbPlGSWRDDGV2yZDWw+G1rs/yCiR7XaLDlsRWtlfvNFFh6koZN8GDis9SJ2VDpI6fr8Cxe
lKO+Gkc7RI+fvVMNOnisA/je/pvQ8OsCsKnp2tMClY/yElVV95NKZh2wzwUaqWnWkVgvy1NygQp4
oMXH1pIlCEU6lTi3NVfGCZzEQRIae7P6py3ToH9Ho+x/KeyKoe/sBZ1vshB9tghn+MSf+rGPqiy0
vAsuQv667nQixvIooxdaShgRXeMX9PN5ASuD+3bJ2+Dh2VjgMSdROw1w0Mgsjv6gZJYSQZpbwpvi
N0XNkF/k8pcykdC34XFLlukh+AOFyhjsk+aUFu0YUfVHfazwUmSpwZcjtGM1kR1GkuOpViEA3E/g
tBNGBdKLarnqgL9rCOrdwJc88dn37inT5KwwdPD0uVyyjpnRH32v69P9DJe+vo4M06SbXpRYykNt
nHIPfzzhvozv9mIhjfQO9cRQ0P2gYCTcd0KDQXt25/FSH2EEvjRuRb8wKEhBjxknnYFu66CIePyF
dtCAW2cZuhWU3EnBcLxfjdQ+TGfQmsEZtDTSXRkjBO7pBHBgim14TF23hjEjHMoaovmptT/SKJlm
RR6ACMsyRV8ZfJpaZRoPWQUevt3UO2N4xOpQLPI5+5IQOFLJWgf4IHIyjPNP6WSB/eTbsyoDDnaO
BYnnwO0ij48YzkwvFjWXJYkfJQ8sNzd5X5YeKhXRMtXp54B3zD7lLgqhbw9Q+p90VcrdmzF6sArT
JDXNaif4w469wNy22l8pm7UVFYdXYswnlMhXCt7GShqtKljwbR/2AnHX1sCAqKwODy8tGYfRWTAP
R3FXNcJzpob0corYfsU/LsdswqDUe499QOxjyvDTnBw90SJOqcsi0qWddcPrgwamkvZLaY9uowre
4nUynFhWcaWSas9fdBHI1D0Z4W7cF/jwKazdvZjN+TIY3b7Mue05chvkhJ+/UWLQSCDy76GXFo+l
Vns2qCVXinigvdslU60kO7R+BCygK6gT4rnRNyvApeteNUK7shmli8pxjfjNpg4OETb0fRO6zWn7
EpcOk7UTEdgNuN3F4OVbGXmwzxsdJ5EZVgQWx1TgraLP4vvpJ6uL49pHDQeRBKCp5Gs/Eb3aRgsT
/D3LqJt7T/2OyIGE55u975tDaHd9MxIAuHZb31ad1+E+sQ5chyJgXBehr4LkDuyP+ANYRoPB8ey+
8pxAleZcQQevVlEJuaogbqqFMUhm0AMSbQkMDSbieqUHpVm7rS5E43/VdoGT4DDEei+liXvPRKPk
CfweYMHOOLeKO559GvJ6I6/z6A9qEKRMJ0bhYAu2gawMrMe+aTU+LQIXsh90WnfQWlmpPnR/3xGn
AcmbtmB2hYqeKMqs5hZeXr0u5verILivlRmVReXMz9PX6Kh0tRxULkr8VxYXMqMFgQ3zTMq96Mw3
fMvxA8vhCXr3S+ZEVXNQDjOLMl1RyKP+iJq4z7ma2c0Abd+tyXNjR0vOxsiyjGrY3FA2CQfiE5eO
9jZrQVL6cvPyYqip6YxnwhT4uuXfOWjSEMDHtRKSQ3OBaINyUH2+JN3LyHUvqAFJ2WVoS+NZZg1w
3DZvE2e4p6O/q9tsv2hKIAYEa5u5kcbnjTlNJvXjBgzSNQB7wJQFR9TNrRowsjgSeGJ4Rmh803y/
if+mmkiFzl3bCg4wppXqL5JUkG1A2v1F4vM6j0WsdxphsrUsC/bWF3Pfmp5C2pqw595+c6I2eyJJ
YKEpP7rXpUcZ8T6JKrVFHzpdfQotD5SvVnLQVCOnFc5P4GftGHeegrChtzIulPND/v9nAFvfegAn
R9xL/a/ZLrCWibKGVTYbOcjvRJ1jJGPLmWMwlNb26tTJT84MYMEpAvA1KjsssH0ZdJIOQnF31wtk
KCsMNW9wzxoGD/05NsdT7yF3a8cuCqGc2bDxFdwQQ2RswH458G7bjWiIOVemGbHX8+jHTNoPGmnq
8aRdirjVr/r6nXbRvrDqjljJ9qQdgs3c98GVKC+xcSyg6h+qNf3XY+y0zhbXWoogPtsaqPKq+vdr
KblOMnYhAZn7zh6Dfq0ZpjFUX+ZCZ86nwq+2GRfeN3xeBliKB0GAP9glLExe+k8emteJ19P5yliN
GJLuUN7oVurBNVrIjro8rzteRJ2rOEHZVm6cplVligw46ChIV/mwk+MBEpFnVhbZh17N36LbbSHE
T9WR/6A3/W7xnHjsafGfrkvmqT2MwRFoBpE9+1bDUfSTPNJTHAk+N9zz1yK+zQTSNlWTwrHNNn3W
9nD03gnnu2aTQnJcxKn66bKFtqsAPTbU4HAQVSpvaoHI5MpMzuTyWYsgGkbRXGB/Mc8i9mGoE/Ps
3QxJQJhl2aBQcQA83/XtIVik6I9KLqnNi6fze699JWvyCTnk1n8/R8XTyNrLSECIJSflpT5qwdjD
Kp2bKVJYZ5tQL4HJFfokFV0DYeNHQ5FmsnEEzE0K8MCNK+qr9RyNSLCRsxpskkIqYoJyfD6BlUPr
N69mSBDOTrYF1SeF+sKJfBU4WM3oXpncqvn86MFSueESjBLdH/VlOyQ27KdN7Mpdef3CaWwF2IjQ
Z6sJLc5hsQ1ero1aYNkr4evb6BBNuIiM+XaXhU2behlc3E0FpepOLnRLOikZwHxFApCgri6ttjj6
qiQOEC6AX0xfhBAiifq9URIJJFyo5ij2XpFPNPm2vChuscl11MQVRam3zIt36K5i9FN5V+a1Cqst
xCTRzDUz/3SnBjl7mOFwkMXUGdA43Bi8SLWe+FUSOyHmymKa8wFDpPMZ9q2S6XPQgvU4OKdmYomX
15pKaTxqIjyynO3zSsCVNBphVbuAEnZ8HFjrWTfIUU8Apxq8R4ICSmFOyhEXH+LwuZkNGZn5Pg3q
C8p34XFOs8MEDi9nfRVBB9Qc8nHS1PPRjlNJ0lZ2bFcB8OiqHp+JcUULGieZrDzscivJRHCnNoXn
p+V1vt7amDAs+YXK40bQqaQ4SvIxkdRBnjPPXNo3l+n2gkBa9WmFGhFexLlGOXADWhyG7uoxRWzP
4FQ8uSN97736GRpO7019b0ANnxYW9PmV8iL4eIrltNQrN07qYDjgPMT6FPMA6xz7ACoWsXZ3SKlD
qTam+84DLrXzLt8dSO41YRInmtb9YY4x+PX/advhT54eEnW44/aBxfawH/485gHdzVU8C3cAKNzH
RdfagDlQZ5v0Nz7ll3VsCmy5SWOKtM8qbs62isZszGUXD0AceT6930R3piMUtuAfCUU3/LB6EXtm
39y4kB0gVPnYbVUuIxx+Ok3YaFgDSyALRL8QVmvs+fgBUofDAXrCdIqQa2lr5Ear2flh8hE2gye6
UlaZ+8jhY8UgBozbT4yFY6FAviMN7A1r1KWAsN/Qe+FmPbTRbWdKCV5pUvJpuE23/vHgIirnrXB/
bgY4L8/FbDWHBoampgx94WXNaSJWO57U+k/Lt5afTscDnbePRsp5g1sZOCtmUH8arYAlSAVhMP7t
h1e2mxLC1/ROkQ0gghHnuYmXMJJlAgjVt6cB4hwmUXzuHI+GpWPEfufCxE+xEIqPRmZCNS3Mkv2D
5r5IGalWEcaSwDkvkS2WnEHdKgzF9hIrfCp8N9J0PMpGiOOzm+6dEo88sIx2bIZFdLsSRrYV0j7A
5fuImOmvF9ag9oyxvAfz28ce90P6svl/IdcQbxC3/RFo81pVxST9enJoXAAEMwKdKmERITAXNzgc
V7E+M63Ot0Ktk7tBa69ktrh/5YFZh7m0yshHqoAVF628Pa4u4LcBhmZy8jqM9KFeDbCKA1nWEXtR
oDVmrTD6V/gxvVCRtOR0Q3XsChJtQVofOHXu5Eb8mnxvb0ezMFdr43g1cTIqxuirlVHHojLNWxYf
tpPW+p5DarPFi7U4NO+gq0wEKPFNRa9sGNmbYqSI0M4G0rfiJ7loiUkxz4fG9vLOoKiQoR7fiLHy
w5NzJd7FNtYu8rHfwO2MVOVYtTHGQl/QAAgV41gk4SDjlBgBT7U8vA88KNa2WpQKr2HdeDf5zCCk
A+rEnj8MBnSSO2Vt3109iswqfi56NHbtLbZUj6YEbPz6Y7YeUPAWzPhdWUt+vsFYmWiru1rBku4r
x276Nmk8ND2+MoKNSVsyojREsyLiWz8ePPURAqqycC11LD4dy0SBdQELQyUcD8M7fZ4A56p6Mt3O
jSe6y5isPL/5fN8oOiuKGCBbr1XAHH3HKmTBnK4uOfTy/hGwPTRmpvjJuv8Wwk5ikSs5NTs/ViPE
TkWnBVms1svBH5TOB46aPbxEpmZ+Q2KbDl0S2mDrv7fQV4oTH1WlUwH4ThSf4A7ub6f2oui8x8I3
LCEFwfAcrMnR1AmWxyoDsFpvMUkFnWNcsMUAnRjYXJX8KQI6WOma9e3LeBS0XmYysKBgHQYCsTsN
WUy5XnuiQbQU6bxAxgLTwheSxBfiEQa2yePmV5T4BJ/oj8Kn814I9GQI8UPo0MYfSFPyqXE6pHAn
PrUFLUnDRTQySCcHWenEZv3conH3Uu02zuH8/5i5jGUv2v4nBN33+MazsjQ3f3tWwcVDsWUPsno9
jQDj54QE/fkkqI2/wA/r1/CKDg9DqRNxHcbaxx6B+bRcwGItJhXEKfa8ghmg7SwyznQvk7IoB5mB
NLh76nmOLxbFwivRUCdqPwfzbmw29Q+fH0v87eosRiZNQOk7POcjDzMtvtt+KodUCp111MUfiaAt
joSfV/XjgrgPKQPc385McfrsD2jp9wcM/tHmqmYD0Okdm5xtjW7+XORbHCLpqAT8wmqLYRvv6mR1
ZnMUdqZEvdUzlbwgL5pvJ3rivU686XumuQgkJKV1aAbgtMIVV9NQziQCDahZP9bPf7pWfWT2uejk
x8xKwYSSnf9rjjZOxV2HPexifvt118oLBjYQ3+P/Rq2L9LVWklhvd3RcjYI2pBTGt2BQ63w12j9i
WByCwvnlgq2etFLTJZkwkexxuNsSib/meoyAUOUuWZAF8fLTmB9LBO0U2I/GqictJkuHYnn52Wda
xHqVEN/pbIucnt04NEjHAAdWRyPasxoobsJJs8+SzMWf8Pp2Rh+SOrMGf9iA4Gar6ndJ8u3Xo/WQ
2tMWVEhDu1P0VPQDJKvVPvRY2SNNPeamsPtSy4qs0QNiatR7dBD7Gqz/knkFE4tgoF6cyYqa4ydc
kuzaZQjYbsws4iLfzfKK5ms3UawHN+xCo6BvnYdfAwMhgl6WkVjVbwHYHBZ9zVyyV5echmwvuyFQ
FdD7tx2ZviGP7KE1MLTbqM6GpeSGnE+qFrZ+wEELqe+1/79B5/XyUTJVf+Vo877ckpryXHNAYpZo
Bv1+Hr4EIixDKPMl0EHDM+fMPzOmMmLeyuOVrLzylAfc5pAGkZmOObquhByZm8/ul2gWIstfw/C9
zJlVaFYSHbiDbk9ilIcC6HscHBzFpSJDFcNfGAIEEfRt5OvJVdrvwRkzzikP9kIiZ0uMyaonCoBA
nR51+TqQJnI9cr3jJmxhEpJQXrpnG6XJFQqbuepxUGJDpLeEUthPsl2zNIWebeAbld4ZWkCB0ELa
0iVh1Ktz+r+eeijrCxExnCBe8Y7RIyEu4cmjv7hCFsDMZrBZiIf1qJ0maTt7BkPttquU25Zf/1rM
1AS6gKx5FGbH+alZ5ruZsWgupp6LIPYckpTQ3Tlz/4OHth7zRdjoT1irD6q5wP+Q3Jghz4WAU2Dg
B15lKbXDy+XUFlfyNtaiLvQW3nEnNe7ZnOIr6UG6mKzIllGdbfbj1okcYdhOtdhpkTs+uYR2v5kl
oSKUK37k9+02n47+B1qcD3Z9Girl4JMnw9tXzDnCw3CPa2bGgspY/uNmVjFl3XzOao9V6zbgk5oN
LQUgSNtUUCUCh4kJC1fr/XMS+uGZ0C68rnaNIJjZ0heYW4Exkx7uV35hevaIfnmFOkj1rbjtOcuT
7UezK6eIGkE5e0Z4p2nXn85Rc63JNjimlBO6wktmRZEPqpYvIi1JYdXSObl1/nDB7IKKIw3vHrHW
KikOI153TqotWdM5yMlEZAp1W+jeemjs5ioFUDMQVGUFkinmx3J2LJTChwhNB5zOkyuXAw6W3eHG
vRf07Fxh3Dg7atW5WulIuzBUAkGHPAS5F6Js2giZcrXr7vdE5Uf/Y/l9Oeh5OuxeYWgsxVtcxxSJ
gDYLK/J6HTymo9DuJRtmnuJ0GhubKzvH0YPp3CCK2uEcNAHbUDoJl/WXnG6ImCj6+lYckZwm4DxN
cTGx9+JRmdShuF1CwIG7lizRa8+VtnzLu8U+xaUV9qHhDCxVLTpm7TGSF8cjU8mfi38Y9KVCZqiY
oVT3DXuH3uafhzjHUuy6ZlICIfOTdy122AysIh9GxeXnvgiB50rSoGB8Trd+z7swoT7SfvUeNr5x
5xjvKvFqpLdldf/7UZUKMwKmOlfGICQMB7N/7MNqRx200LxKdORUszPuP3Ddf44dva6sWCKQyZ19
rNSVPenJcssx9SRS5VKWTS+ETnNUImArFjO+xByG2bV4rHSEEekCguzmenwaBxpRYn0qAIN+DnUT
ApmeH2WBdxy67aCjQ0FX5T0VW/hV18HFbxJnP54/N3FzMGLfBHMJ9B6mDIY9HBTMQLlV9RS0vdJn
2qFtw9QeXeMOU/NpOjpkIBKA01FNm8jQbqpp3Pp7Vyr848Svk0ohcZJv3lQli07Jlo1EpgrYIipl
d+dY6AufFltXGBCu/rFMCn8+HFP5KuA83KpdLRGYdfMSAjGdcTlsf48ALQrH7OLxPb2/G3z2rL5l
10fjGcMR2A7JpDjCMtX1KhGFXPgRFSNN/OLURcZT2O5g0JHU/UgvUWsYctxKLSttcnWgZLnG7h+s
43UCJqTFcpnj6inVRrLpttUrnTV2GE7LAVmtF0MT92NgNhJtsxWj6E+dKYYK5M/AA2VLwqe3b/ti
Rkq/Ma4dpaCy9AMcIPdikJJ8FYXB3E/Xma9pWvzPShOVSjcKFtgFTIK3IyxlWM4wwZilCIdaVcoQ
PWIK0MxcwpHbFmzGku8IQpD8bloKUCWUn6hWwQYkn09pApaVvfhiCRWyS81l2wZnNkHM9+xT96Gs
w99hALOGKFp3QK5GCJ2j7WxfgHUMJ7pHQfE9TVFGD7mCwYLUb4ShVOHT9+W1LT4rT8ckj9qtBBUo
WwwT86L6lFgg1IVlGWlyPDBw4grg+2r0TcCwLirIJJ4W78wIJC9JRHlWDRJ+5eYrUyJAKR4u86Ib
8hlTxhgRXMLXGDGwxFBe4T2YcHfm1k7u6cku8fLauDumq/M7Nru8nmtkfCbW2XCcRQ3fWZHApO2m
OFKqQXUv0JtF3kmEBJRqekBHJfp0hQlo2+5cUhunB1GOIypgHdDe6aaAEmgzCZc7OWm2Ksm+JFCi
f5lkOcnvUdzaY2QGnG9S6xUszCAjpCEmu7SogK8nVkDU5WrvNy0kPuKTivzrl5M2DBHbrMCqPMRJ
2V9tRy9n7Gh0pkDd265XiEv4A5A5AcaE97dujVEpbHgM7U8KO3Gy1ZUIY/rIvr10cC+kgtkzhk7N
IkYRMI6cKJ5cICALLBHQyvy+UMCmDmvD72AUeeu0md3GtxDMBAKgnY62pqRgAO9X5fNNAkpMIMx8
RTsUWfJ1R/8foAr93i9IhpoiaN6CXTLdNkE6vvDrWTdEKaNv1Zvq1wh4Ag+AX+K/dt0dMAnzLBCA
4o5nMaQoLJQigU9tCHJsPIUg1vLhnZ0vbsVmoejv33Zwk1OLLZIhhyQpe7znruhJWWtCtw+a9rUP
meOoFqMqGvzLDQMB6/crrOzsqHx+hg8BLk8JQFPTETiQB3YqNIHtKkf66Ic+kVYNOr9nNwBLpMc/
R9qM5ZBqDOfuBdBmJridMoMt+MFnBbLAqtnPucjmCf6Qlx0hx+C68daMwZkEOXUWMuk3/IqZ803e
ox4+JZPt9jKC5pzLHLHHBIpDL7tqOEOqlNHmZ7WHK3TBkwn+MFGcc9y/mTNbajpG3vn0rpmoGKcy
JlW6WtjyiGvCaTAKWpyfmDzOSH6wgdBg0vOSP6PR31MkO13bPtq7iNLSu/+uwrU2rc9+Dil7mAd7
F+o8smRWnPM+XPPSiToVK1atfPuDmeGmz8nL0udsMJFnfjcM9/w1IivdHvEbiFQxbNYI2jD+2JKu
R8YtAfx0JP1xC0KScfvkkjCpQBGpw/wvgWYzDfQH9r211CbSLoTGAYYixjDFI63A2YHCRrfYX0FA
QkTF2ECGH1RDwjMPXmB74gz6fYnzgo6kNGRtK02r72CsZvrB5zxcQ/+nyyIyClGD4KLJkbS4QSrg
kVB6HRb65//vZ1LhKGkpdQN9xVEUi49uU44wAUpFoXSplbKHpDgrSGVC8HtkwtL5ubZg/FDNP14r
kYv2n5GSrr6kOYie6hK+W3aSAbB9uk0/P6PYKQMAOlQzt/0TF3Xop+cJpzxh+QSAL88MP1E7Ax29
en3XzSWZRMWWpCC8ZFg4yBJ9D/ojGA+cJoYnubDLfrjuUHHeG5imnGsaqBD91qe0TLYxugVsFkVH
hUUKdTIQoxt+Pn4OpRIn7TgR49hHbnZ/OQQ4HQsmkvVi7JNvl69eokZfBN0TMRxvFNBUIIrqzx4E
ka1OIJKXNj+JPdfc+H9IRmHA2OMeJeNI1zdqigRhc5ixagSi1+G3FvDaXOKQu+NQeiPvmgaF7HyW
mIpkaauRIG5FKP+LO6M4xDex5kK6g7dIEsUTWBTsMO+q9ssvCcrjnm13fMMhHEu4A13bW+XT4Jre
Grepw2kiDtcRGD6FmYzaZZHF5WNtLlCUso1qxzWx+qCBfy+JulzfokWhWdQnEqv0eJwHUJoyNJee
N9RaWVl9iGfNhyCdDGFzuoUMW/zWJse4aFyNKYb81r4PkPEhGco1YmalIbc7FLOiYR3SBxA+3oWg
5mK1VtH1p7bbinMeHU9eLpnox939xMbHToVevdCymJ55kd02EKZ6RHS5OgsB5YY0bnTgTD3wVcHX
O/tnA0hbyG+sonO60SmLVcSxmPylgLGSTOcN78U6WRGUeeKUu/5jwFardsP2LbLjrXJNi2CCjU4k
mhBqpDTuehdXhVDJHf6MND3WGpJjVKTG0PbZIBHQ+OAiIxi0LVAu1DlnhO3mNgH0qykbIJ9+vdjX
ItlKRYl/9uRSKCfgBRaZ6809ZhuCbEUjApbfbLsnifbp2cKcGShnxcSui2TDF3JRN3l2tOTfz4OS
2yuINYRUZSVVLSfzPu1mHCfkOI9zSMmfMWr/l/6PJwTgfomPQds8Lb13hqddx4sEDNeitSY4NmoL
K6b9xM/yJSC61nDIrblRuK9aB5CrdTYZEwF4mWJvy0z878UqT4cmh5/D+iK9xZesf/iuSsbLr7gD
ayOI9yoHGBO+If4u1Wpl1Ym+Q4FKJibXSFV/Huwt3rckDT99D3n27Fspyz3G8I3v25C9urcIgEjR
JWxDW4nrLVykXos2PBzBLCn1i+EMnEtmrBRUjNoZpjZGwnItY7cjbEwOVm8ierGvg+YPZ7dDZfFi
h0IPiDJTR5TL8trzJ/lnTWIG3jMc9MeV51E70OVt0+BWbiUGOT8BI5ADav0US+aYQPwqkqaBcsQm
kuOcdx02u33LkWok0GcwEgoo6qL1SRzuverH96J1PugVafE9ZV6Wmhlx7lgrVeRD37RsTborkT4a
FlUhu/9Isx+VfhLVEyMw5/SMkGRFfOhK/Vm/wu02Hxb2Q8jKUlonxKX4ZjcpSfGvQPBTPS2iBFrb
y/CmrX8z9ggQIs/Afu6rY4BMeeLPnYXXWkkzHKe8r8P4tW9EQdcZ7XBRCsnTZaMW7sLza6dJmYGh
Zv2t5uS15//D7li6V6GbNPvG2G5p4ar/3exkFimMQKttl7UoKVrTkSEHCKY6QhO7F3O7Q1yppoX/
6Qd6VZioeeBxbcSIWdaJUT4X45YPFaPv5jJwL9v6eHQO9CuQCujEHADvT3MOtCEJHsvAeVCZiYEX
Zbo/6WVU0xxSLMO3tIwJ8/5fMSRdmctpqFB3qESsZ+s47esCeap8GwJCvHvnfjOzgT5vHJubr5Ba
ynPbgTd3tevkt/5hv+vin21Af+9KJgKZHW86XRuyyYJmWLy7yi6tCsk2iRbXf13PO48kaCuXxwtY
bhi4MTHVdt7kyeuyboE9fvY703Xq6Qx8DoL9QjkxozysOiREk3GdBfGJ/3lWIvTpI6cF5D3FALQe
mjma4PcDL+w4wkIU6xIwHFZCxgD5Dwq5HdaLrS8uEEkGr0WXpWCZhLtdimog8kTjbMm2pjqWJlbQ
//PElZ+5fVlDt5a+PxBmHUiTdG2VGr5+aL/qzxt13m8NgAci4nXOegxDbLkUoFX94Tqm85tp6rp7
3L3p4royHCdfN/6i4YRpHqjXj2ysalEpEeHIVhow8y8vdqpDF5KuZSku8vZcAbhx/Xug9JUgY27l
uMlERtkAfkh7mOxh8Cv9oVi82NiosNXZ9i1VBO8e+4WxOUUe4ZX656lI1scRSImi2pbDf2bQu5UK
s3jBAVOlDs7hAMiQvq5RN1KZcWjnWfB5D1YTLz+/a+uSs15+VIeV4WvQZv0ZtiGxPlUscgmgg3go
9LElG+IFVP6n/nARj6NWeGM2HBjOB0+lfp7XfSANLdo21n/P1egO8Y4VWTPVhf4gRda7rJdZS++J
2pglvaS35e6D6LgC3CMn7pnkJcWZwCb6Q8hqJX8UfyzrgETmFBNvYLuLqZVsdScT0mJenhLTQE1v
C0ePC9vZand0CKQPpCR28wynPuZ0Bjvu8V7+Zz4M0pekJncDxaBTAIDMhibaPhUFSNPJ2hKLqNQK
n4mtY/b0LnCeD4UQ/F5Na4OK727TxtW7XZbeDWbZ2TKeRiUbfTrLhBn0S3BGjn1AIsi906YvX4pR
PYevHzEIsiJdmeOOKvrOaxaLWBXw1NVlowAiQSlO5sspfKaK4bMuHLyUWJM2zcry7olpoLjCJ2UH
NzlyNuf2SbcM2nEDqX4EWICvpTj1NaiNjpcAjJcs5wi5MJBH14829Ejx2QlCNzeUiA2RJpHOq81b
WUHg9iZkg5/Gc0U4ObMQBx8QPwMD5KXw3MMdWaSq7bKkn6Q/V9QJVqapAgaI8hWtv9GFW2XFGUFZ
IOLcQGdHYKGZPjxJtMXhA3DR1PHCUjHAs3vZHA331Ztb2ShSk8RcvmskM4Ie67Cx7TZfjiZfSclW
9uSi0TqJyGt0BUov/3yBUfHK8x9Juv+gVgzxlmdXH59tzsCnU3H+dOg2P8HwSvfLKpkpyz1zfix9
7bLETLkYESYKRYRcemFEk+VaRJwAEICXfuJ641QD72HSt5fCOMcMy7bWR5nL1Y636EFj6NnR3i4U
mo9m56tIWsHZ01shHvLkOb4ZF2mdFcxmKwQYAs4hss44bWKKk356z3znRwHTnppvNidZAeT5SI4P
jjd0EIMWsRaXOZbax5vyDeUMlDJAWojlEi2Ubl0L9ijez/EDT/rM+fW04S674JuBWHWIDWTsF3Hs
wSNTJVjPab9VLOyDWcQXlFBYtZneBbKdndIdTAYYbxnnFA5wy2u7oa0s1DbALrxlI7tsHUtVj8cm
yGHLxhwbjw3zbex38UuWmRmiKQth3VgW42CphQYA8kAqf9siQkGrYsSR+2nWYpblLvA8QhhK/QQL
pulC6oh3CjxDssXXH7yFdorDp9uCFl3PjZNvgMGPbCl3Cs5yjsCeA+CQYxq7Z+vryjxPhlCQZkRo
dpuDJ+osqlo2iE0XTD7cKxf679Gi8XlvdaRWxm7ob7U0c4sovKMvVdIy+HP6XRThlJuUH687HczG
n8lqdvyw0WX3v39jpXwXs8FOW7VgHbiwl6O3iAxQWY3UfZdQ16os1Ij/Ryg+Si7agjRBXU9X8bDZ
D+y2LCKjffFtqjxi+SmEiiCtAozd4K70r7nA+Izm4WXAynbq+uEZHIwnz8fL+bPjjiiy+6EVc2Dd
8EiKctTK4SQP/e6+Do4+duqbxZr8pXvqrrcXOzBk6da2YViV/K5Im8JL3ApYqb4XU+2GBbItiE1I
UotS37y4Emu2jGVEtW6fdD4o7LfJPwe4GCBWAmbvOygn4/QqjJRgqsF0FYOt2gpXshw+FKDplKmW
244GC0Un9wBqM2Y2yImifWRexaD0Kl1GpCJMC1LD09Xw/4YUBZACUdzlNbtR+acRrNYA9P/RmGsr
UGV2vIyCfAX3edbv8o54AMg6eRhz0mv6OS4pke9CtgQRj9lW0Z//dDLVjxHhEQJBmAxiLMQT8Yeu
GoYotGpMSRlQ8rDNLLGyTXMy5yP+jEz1ok59XippEi1S33OagsfpZZMKNh6k7TvLIaEydAJNSVYL
bYunIUzsmuzy1zGoLiJsFDAeVmASAJ1FFqCC6ilmNo+gyiSgJJTk8G6s+AaT5RkuQla78BcruSTk
X9Am4r6HoJmYN+l+Qzbgfr6vQ2isXav6TWptSeLBrKEN33JzKV4jq8YK0Gv8bqyMebbOTCbp4ZHC
EA0uMbH/CldJE4TYoAI/00Zma8qyetSZu84E4r60xy4yOLOAPScgyhZe4v+i9iLi+XFVQMr8/A+C
BVzhLrMZk9PmMOxtzLRryJFvCfQirY0qVQZjEP7CUXJo9/XN8jEh/I8Y/KkOgOaEZcABbxpWeUzX
9IvCLlUQ+v6daE64FjzwRWYRPWrI4N2WGW7UmxIeqk76UbW/xMSBS1vlPDCRCxHMZTCNWm/dTpNU
2e7WgQ+JV1DT+ZmJrK/f6H6giRwraqnTbc2APy05x9WU5jXg3vne17ONWifZA4In6tLHGCT/yvLS
x9LHWsks1e2aC3gOSwpJAbYgJ66M9A5H6PUdfrN3IzikvkkRm6u2+fCT8qoO3iWH0d2rxd72p4vm
mvcvCqY0Wm1av1R7b94BAZ0m5Zu3ITdtsMgfzlNqTLmhhazkUt2atLpIYNw2E4PMbPtjh7pxcoMI
5j5BHx5B8qKjj7WlYhA7Ik8Rp9Ehz/tatXp4yrLF08CidRlquTtXVNDNr4Sc7YTvOI/JXNvu1e19
0bKslWz1W9qiKF8sUc1HlNnvj8rdjfLe1Dw3Q3nJr6mofSHQ0dsPu4a2Z+TorsUygh/0yO5ekDG/
LYSKACaoL2QpXQYaOPsUJAyZOUIhBIilTZh7pJlhWAfAv3PVOgy5ktDPwOPjFpVfo8ZDckZTy5uu
h4w4nbLjGJ2svu/4o1PgXYzq3nbJlTGWonP59O50CpoiEeZhHZwFz3cZwtdBd0ezrWnRI8lSiChX
CsyPlzpEWJnj7sUgt3IWOw73sX8peRogzVWoXZGTTWIkky3tSpNR+K7b33nk/GHN8rtlqfMglwVj
NOxBM0CZWP2+KqoB0/gDGoGDXAGzrCVyXsshIm1ey08z4NNFY2IUzL71UEfAh7C91ZHpnfTY/+9+
12iHtyL8jfDiDvhoibg1UdPbHOIDhAqxfyL+6dXID93GUWx7t1nNg7k0akTrObpliXxHE9DNvxVx
65vy8wV3OwKEQsm1GCjrwdev368pQhLSeKrQHXdh5IG4XMhuTs9yrp8BwoYMwwcPLhSEmlFVpgRE
t31J7cjaT9iGLEuQjyxeKVdwIZ9hk6SxWYfEtRwgKvnTF2NMd7mf3zz+zvy/GKhBeLSvQlhXOWG3
cbxwgpTOUD5uR4rsSPEYOm6u6b1yyqJzZvyekrTrHBYi0GWHKWJ5dFT0BAcQqK/lPyOeWkr+YvAf
+L51kUthIyM8yg4nc/fFYSBvRx2yLiJhqXxA4Kw+78ot/QunS+1epuzlIQOkp9G/fhBcC5/V/xrT
TVkNpyR1dSyxyAcfo5pSsoPM9dxlvE5EYreRssPCKbKbaP5ulO+r7obrgKTwUPwE6ZHzkxG9xZpe
iEPY1dTb89ZVgD6+OnY1otjfTS+fFWmSxeQbxVVPMCFcDADVZacWRPbFYOsawqMX3aw2U6eNj8bn
p/Apf7U+mVorCkIuVjyY8lYuFlHxe0fVoy86884lME3gt45AN99p9HSmFcbyBhOblIOqVuDoPwRY
tqZ3z1zUChhih0jUgqUhHQhkmozq3SOpNGEWhuD/QhvYXaoutDpZM29vTOByVx0+oZYXeUwFfK+l
Hww39b8MGEMyRlGvUDJwFDyDeYn8f+hrXZF2+iKaz/BiHOnqdfTonVVS6qYkC2S+hZM3aurP+cbx
kY4WD2fKYrpISuSxvY0AFe4aD16YlgZ33tx+qgQ2iphCX95/6R6OhxOm3ct66Zm7PWBra37okpdZ
NoAAKJc2RF167TorocOiTDSHBs8DCuEmcZOj705PoJ2xLY8h0essgOu5X/RXhMzHG2BtNSBhXp0a
6SEXuVfO2okp/fLF4JZ5ygSdCqqVSvD2FibY2fpMLkql1JEwPxSTPMxsxjw5Z3UkGfqEpd/oJgN7
nwXasJPHfjQLQNOARneFoy1aaREkkInfTMW4QpPkNCXrsGrM9YXrXenm1GaU1Rvb6Sc596C/T8YR
hVO6RxQDSgMLYoznLaNbZEK+db7y8NmG3QdtGSaABBCsGVapG7EnNmbpghpu072tnEVV+q2HcAhB
G/Em2lvDg6r+7kuwq2pCF0ZmvlwTd500px5W6C4/4HkndBYQOlcA/xzlzjtSK2vriIycJqr+dEDD
zTn1iXb35+IC491mAFYOMo8LOAX3FCA2WP5ScfJ/RCJ1LNqTfUZ8XZ5J1IiSWN78s+D0A92nmAuU
9vXDizuhJkwyM5D+CDDWg5NNhkRBugW/CK1psl22jEqfqhHzEmV6mK/psDRnjgXuog0iAWXUJr3l
1KnR15mpYoMOAJPaH81SUHoBG1D2IGZU0vOqvOWNByNk+ri8Px2tyhBfgSIRd0xxiE31SKRfKpRh
4H+zcreylj2W7ATJlaXrODjrEds+7ca/T9jzko0U+bZRlr9/dfEK6033FlQpSdfvwi/TSG6YDqKs
Fug7mZX/niFDS8ddnlWDBsYJnY8iSRllVUJcxrCLZ4Y6pQ8ogorh6L2qKFD0ZHWMTZiE5ePenvPH
tu200P0nOPuYbenyTMHK9kdXolTTRl2KT2Tl64eUHB056+K5SAKcQnmgK4HuuAj2LTfqh1ZEq9ES
kiIgQsM/m69zIrzm7Exj/R9vw4cn5TUXdJSxImFwHPL2SW21+t24PYCdjsjll1UTHQq/6wViiXaF
fCuJ+6d+490o1zzrDMglHXnlkxXxL1CFCDb1Lcf8sbiq6zQBi/VYpq828EFndrVK9BL5a5/G92JK
Z8DZ3wJUuhBtukcBhKxZeLX+ngegTXIShLXc9eDaJ6gqDHibrBxiYAPL9HLJR37NigQvSYVeoI/z
CC58K23p1ORDa2xICCx7oZQavA4UPzrzglUwz+leyDuZirba7akgEUL4iU2HT0JORbJEBbQUMsqM
14zz8G4BwF7sZwCLv6adhgo/OJOR7DzhYotiki1J+/Uo5Cf5Zv/m+8j9WGiFHWxzQivS83HLbqsG
cF1d2vX6UhR8JNKjvFYon2OJc3DBQe06MbEqgByGmBTPp5TUKd0VsnWpEvG9AY7qmdWRCsxKQQ9B
lNANEhvO/aJaK4kOLLhuDJV2ayHoCrY9PWkvluoxWFZCNvKo7RTvo0Zf5ShoAvPKjG8MJYfTt6ON
PZBTCYsbNer7TGBf7FH39+j+acfSm4czbDKs5mRMI70cGHeZkbDMm+CwKV/XPoldZk+cvpvSXED3
8rUTpBx0UV3Ya5DxfEQTlpcbSrob+XsKkKrAZplI77IdHsYxA4CbWR/c4sl98e4uW43t+0hJPurk
tsnWGvnnH7Hk9o/+5BFQdQTPUDK6WsRgSIEpIVQ4OFkeFS8kntgAs+W2Lr5GjZ2u5YH3fE/ES0of
awO3QqdtV+GDtMBt/ZRehm+s46sBTex2iIXIbEWkX4idQjf7g+1I4XtKf8RC43J1fArACQuFCbZH
HIRp05K2hLvRmkBQKjVJVJNUJLyIKoBm8EME4x5Ie3HmFlrNr7fKxpoJJB49b6w5AnxqcdJhFmcX
7uHaPiOKoGMsW/77KDiW8XDpwr4x3KG3CTNaAlGJinMyXCOhT1FqfxVXzqpXTL60j+EL/YNTG6Nt
HzU4oUGSXGVLXOX/KldvhNOpBPgdP39e92nQCgyvp958K0OK2dgwGB1S5H7jzTMoEPTQ3w8hnEb/
EbL8ZOE3CGmFMsFfsFbdYZk//B6vMkEBtuZ7TAKbNZZCgF2JOAwqLE2zLT0q9njJJMId3Tdx6b/b
6PYVmTAbdqCxQJIE3XZpoDKkmOlqj1a+8hGbaZgtsO8mxAr18mnxMv1U89714FJUtS6uZgB7CIGr
0dDhXvQ6kklO8JJYj8IG4YBtFHmlqcF9Ln69NzBdEUqF/tDLLrUoyUYkX5XmXXaIJKEa4kfvX0Sc
637Sf/QU3iIyww0O+TVIAEwo8zdbjY1AO7bYxY/9kRSLb+MN14LNPUN8XJ+jB7v9zeKix4cvJBCS
kyFQjmhQfdAo6vpLI9YJUnXI7uUrP3RLlunoyCOFjcBMgwzE63C5nGIpvzUvVGGQvgqwCsCHs2wz
PoxIrZy6XZGVVyxAnzso09dLZRXs/CbSK73mWh4HfAQxk06ReJWkRq7tAomwqin5oJEnJqzLy3qL
0nTiWpwtQUopWqYf+3VkO/O5VcdkrpU4N9/nGBlnWTUylQfmNrDsXzAdYkqCd3RALRJEFllYpcpy
v/KDgWLnt8Gpq3DQdzsAYnMXkLqV9sdlT8LwxKgU6liZm5q2QWzRcFTEgHRVB/ISUUAIu+RYkZpL
K0oxlE9saycsn8Wn+UlDUpSKbLp1cL+NKJ33NAfuS3iq+HPL4T46T0PeC5snPb/YFvvXV4vIOH4p
iogIc9CJtKsMGTw6lvOD+82SI6V6x6o2v634tASha29DcLmlCeyhqb8oJRNCL83KXkdj9NGasBwx
/EO6HEc3IC3fF0r/Ukaegr42VwUASE+0ZQn+chFWCBh8DO1nBtUr8zzTwCBLoCMFc4e9PR3Ccai0
QJippkS21xyEXZjFlPMcpLZzsqFpcyq/4Q+yAeExAiHov3nc+ECeTDfdF25w5AqJvFUCyfJJm4s8
zyXMBRrmcsNDDOLnYU3LMXCIzNURqwmPwt8m2I8Ds9wyy/IAXnP5j2g0x39ydIW9FtP1YkTNiaQU
5/mi437W4o7z6KC25EE2YrEwuQkYLT8k+nTx+xwvLnEVHt+3TnhrmsTgbWTFemZ7MNvFHy4pmqGd
P0r61TAGE2avx5W1qZVMiHirr+8Tk1MkQ2RXB4Wsf8Xv5fhn0JpBOU70ec2YUelrAxt/NoFAmafo
XLVzZ3tEOLuVzGfIj6FAz8VXn/NOyQJmxCi+yhOGXPVB/fPnLsph4VCsYd6b0EJUtzh4cEgXL9vM
PE0rZUb0JQq6G9LlyNcdGJgfbbFyn0NwIqEelxL8FWGmu+S95flMPAMUfv5yZp3fRypSKXRsgbev
uY62smlzcyZs1LoSjhkkEJa7yArcQWrYBZu8cMjinrJIJV04fv/4SUKRzrvWEuzLD0nyP8smfygu
vB1Ft2/+2ESM7lwHXrL8wa1E5qXQaCQ7P/7c+AhExJ0WTv8KV3nt1zHZ66q5DIjodD9c5PvtfvZ1
+y2lnUG0VV0E79H2r8zF1GvkrBJRqEJ5oU+21zSiihF7qtSmd9ejYHALjKqxfXgWM5rbil8uAvF5
6n/lSs7mlD8ZjheMAKBgidgFjEYw6xewxfDig9X/VxcBZTH/fpgkhtIOdCilYn5194enHGD/CXx3
GrOM6npvvUtwetAAuEui/2uoWWij785L9Ok55bX6qPpNozxi5ZOp+/IV4DPWCMx2eB/QWzpKBh/f
jurtDvOEeGqT8WfqlpIET4LobgVRZ8apg3R/S49nLmjiqISNeFxF7ySsA10oeHSqeXCAIlWNZY3z
jxB4WQ4enyl157LM2SDdCyMsggcEyyx6YVE+FSwJefv3veiQ6FVf241/6q0PMtJ7dujUwDxvolRn
46+TZVWGVe9UDlCSlV5sDpof/l48kGuGm6Uye0UKs5V9TwyW+zv1Z7kMhFTJt5PpgSbMW8MVsWZm
JXbTLTQlXxFHtE4/p9/JfXVQhYh6f8jqO5uqfiE3Mk5Mgbo1AInN3Y1oIpgpij5w3tOrSNsjzQU7
2/QeX4kVWjlrdNl7M3rYiS39lCaPin91IAWH+ZktpTyzVsQWUuHoCdZW9lYbOKbh7CD7fG91tSpj
TQmbP1BwuxR+fBimEu4K/UkwoghjVkCSwwgFL/dmXD/RpRnMiNAzMGryleIspdaj0w+H04FOkS/G
oadT5MvZGYwlYFtpxfcJu4Fm3TI8KfuoTwLmnAFyE83eszVvifpb5b9xWmdE6ncn3Jffjp6PJ52I
hL/CwyhQ2+v5RuSeJb07C4lBHCS2QrjB9mmEaq9xaGwg/NyC3OkS09AxbuBWXSvj8ZgRmI2/FgFW
bqc34eFpdBE/+6ClTA5XMsxxpQVxxXq7Lu5mvHmiOVJShZyys0Y0Qs6vD86ZtdvkpmFaVfEn84+3
83db3Nykyqz9jFs2MhUr89OfRai7P6m3MoljzpWt4KHGYcT+ciqhW5//DHqFjIV3tvlaZfiIhFXS
gnB02gB8R09LTJWWL3C80fg0iM30Ape/z89CpIkE6w4r4WUFai9rmIEXRbzkWzzTi0WrlU52n3F4
rio7HQ6Y+Nojq9gkU6KyhB3+NfeXJHBlIzOGfON0vTtjTRaplDai+Cr72clyt3JA2AEc4e+qF19K
Lmj2Kzg9UHpcgnqrBaQtuaRJwyh9EzAqGX6UMLdYwmZfueKX3jPOdkKgGfVe6q0zbHqQ7vQIEE2H
FjlCqw9NXTbDXQqO+agu7v1dh3jS02a0Njl/wjKDbtuk7t1PnYB3Syk72Ll3NYwYnOuY2pknqbWg
uF6ur7oheqW98z45zIXsBia53/32aXxK0Zww8wQn8UiXR5Grv8E0u7WH8GWI7WlqudTFkVjpOjw5
bnnqSOHA9MkweORoOLt9sL/6K4WdDwcQC8FUe4/MWHT9ofApFVbEHmIQtSXxYiVgf4ItsM8AoYk3
8zzu0m3dd4rTSDW7GeripZanczaiufNVoze/L0V4uJBWM+RyKIF+57RUJtZEyg5Rwk8GGATHM7SG
DTF0Vc30eGtpwnk6TK8Qsyjnxg/A7XU65XBWVAwz5IvmArI7mqZ443nB01mOEGWS7ajP845GqM9b
bw/RS1rGaSxmCUPX8r++NnbKB+tLByutUBIzJxnqXfYgBSnzekswHycZWyidsctbE2vAdeNxInO/
c5VL826BRjy2+hs9y3FD91gWAkE50lWtRE4LBar2SrMA9a7ouTtYpqwTTDqkT/q99I5P/EUWUyHK
gHNzzylGKELunMKnr6Qm8DRmo1rtaJBRIvnENF7EQ8e2TCu144br8qq/wikw5mWw/dJ+gqoYObxl
ncgTw6GvnPJheSD4+47Xxq3iR14i59MnuDyzT7goEJwCtU4Bs4J2yvtYx5ne6CXogowKq1nof0sU
nfQrXU7ApT2PY62KHXF9AOxITV+l8tRIqKvIAuUzXFN8JKy+CggHaaGwNKeiwoDf3dDNw3aJncdi
JFfhjKqGQ/kEgmMJWPb5eOgULmnL9Fie3ea6sANbDxis2+6kMtAJlfazu1lWjErZp+a9ZinWZmyp
/wvh7VEStEleCQDxvPZWsJZDWa/HS4PeZ+E8OMTnWqQCXuCxuYISs4PuBpzCnq1cheg/UFnsv3EH
tOwL9N8Adv2a8XF22swOREkbTsibnrUbQGZGG0YzTwlEZIaApm3qIgyH3J/YrcjG/IvV+0vTIt11
FFniKPJ1WSMcZKdGz8LckoKWRloLy7NquTI6sYl3iSm/SHRg2Bcw5gyE6zbjn54aUUjBy3IY1gYN
idVZgzzJsxKiDXE84z6dkeTi4on5pqx6Yp3u6GxJiK9qOyEpe7B75k76vql6rojpUCoQu5XzdmAM
xanRn4e1qFpP+9QRWuO00/N2K6EZtKuj+JLCqr+T/GyJIwUU+jT8P8MyLeXetqTWGfFQzIH/r8BW
d1pnYzYJWLUs8HDxrZyxs9ff4q7TbXg1vkoIZ7dilLOpBg3eF85c3P9YmUBTlBNPkwibZktSt7S6
dXnG/GDeP7IA2diY3lDy1iqxJ5ozsQYYCZxcSKZSMD3kBgqkThoiKK2XEW4bzeh140dZCOoCSWVI
kVhMKAOlvbG95bz3u3eGemmd3Vc9HHuc+mn8QeYSjcyautEva5sPZF7eg0M4TTosYjQjP+Rev6jq
Q4n5iUgmtxytEcMKLLjLlij3MN1dxrh/RmPESxw+zX6MnrWRBU+IZfBK71aGiYnQkY3DGFwH7tm3
sT6XSgR1fgpn/kOeJRTy14bzyEuzmb516RuyQBDTdp6WxXdwYAZ6jadrUShRd+t3FG9xYSodtBC+
AbS/ZN79oMfbt8/Xy5c7loWkfZvxz2s3S8zxc6AWkzpJfHkTlfm1M/PoDeiQo+QWmTNJpk9b4Cue
XcsfLb1ei116pjf5phHOtXnRojvelqtIbvVuo6Gn/LLhEnEjdYwH2uMFb+QohDxLbdiVmQM0Th9T
tx5yDEwpcphAda/7q3IKSMU+ueTQvdur+7qzvXZz87bVoUktmIfJIj4jLo7ZsNUybRxNtJxL7s2k
IcEvPch5X7mQoi2hfKjt9Extvt3rywnNjtvtvrjbFddJr0WLN8wsx56/6nBFSxo51foF5l9PCKBC
EBZLoSpit3C1g07CBJ9I2nUfZzqRrrwMY72Pq7YlXfDFfBsuUWUXEAdyNz5FzP6cwEqC0pbaXVIa
tyx2/qr4xxcU2kSjywAQxDcB/Y/e3b95PfxAOEs1dLQm4gRIxOEAiuPyme/fJ03CaYD/101VUSCo
5s+sSXrkNlrK9rU9wBAwe3YT8+YfaSYEilVuIdOEgXeQfraqtOgoHcieZmjJ3DNlFwdmemPJ2VNx
PDLmhG50KGi6rzgFNfQEL3Y6ipXdbkDosNISkuthNKoxZ4cGGeYBPPZM8ZjaPItV6s/LqUrD/FRB
SPndy43YVYB55nkZMyBN9fBMr1q9IgGdV8s6197cp1HTIYbaDSuKi0ZFdBtz8cuURoVsvEH9uWbv
ny8oO0d/jOVWJDUyKlE/nh2dVOWjKtyZU0oDR8kL8aSChu3Yd+F7mIIe7SKhOqhkGx2wdKApustX
d+kz/wz959PRfcGZuO+uhviPdZh2VpuHkMeSf4NeflVfHawzOw7aD/JRd6neTXPQiPsLIEpokwz2
ex6DqKxV3diTB/eqSc7I+1MbkXjIHOx5DaOjRFGHNAfu3H4WG8P+45ejm4MKHzYcJWn5nwc/87oz
sitoSRi84ePf3/+zle63JQDq/VCgKGKQE3KeOs0QKcYmtrCcwDaS40UccFqaWkNq3YO1BJvl0ThV
KE/tmyUGXgi3NYd9eOOg/5Vi138uOgfRPqUMXzodq3zLlnd2e5k6g3x78j3VNs4Er6EKq2KpO7JR
UOAllglQywrPVCEGhFyq1SXEzCiGROKEYpwmoHKIAA42m+SWvNslQd3y2Zr0CZJr6kBWbD3Gdk1H
8IvKtA/6jf9jmjQkWILhKmQsovNB+voc8iOiOC0KlOJxSfB13TKlOHGFlCPkqrQaCk0h/T9PqwwH
I/LAoDPg4ek7zg8RAVVV9L8I1Kr8K6Ab07FDqgTzMaTiThawRia3UkR3fRom5t+CfbX3v0ASpBpM
RBJLPW7lsxEmTTxFUx7ZOCPpJRYoc60bPb7ulmM3Y84qOfoOMSg2lGMg3KjZDmKzAc2lfwPHy/sy
eLiBt0+JJKq/6pX5diCJxOk54B93sMK3TyJY8FSHSqHbyVI0xBUIWotKTADqLxo2yCBoXTmbnEFS
KTdbnJixQS9J6VqX2l2jJyd9WjPaNH3Vrmts1iHdjWISf4pTikyfaAe63aERLKpTosMLJyheAoki
u1W3jOPwCs+arEV9kkTo9tj0TELYsbZ20JtsGvcZDz0JIBhanqOTrg2L4h9+BOeoDiMQ029N1smf
wmn3bUQl3vG8KGbG+wow+k4WIqcSYxdeFirSC36qgqTmnPHxBNWLsfBuBQeaynff3LqPZcbByGc5
0j6659OXMO75TRtbhWMuRZFAxjUtg9QmgD0HPjrDneig77yLHSw7RrWGnw2XH/yqwzUFPtsuG5Rt
DKAPBBU1UAH+UIMeuZXS9ddHepqiSPY6qDeg84eiMxvJptIel9wvufX41kZ8LOe82rJggdyTIWfK
7MHhxMCm1MJClOEh92DUrByP7XW0zb9VS9mYjPEYa9DDTi2wft7HvEE+0F+t3BzzeV8TfXNtEcE/
qAssK0BTw02UjvjBzJyQ56zzzLXmL57sG1Z2zGXLlxCd4TiY8x3b6x+j9tWVSXJvsJA+7pmHdd9h
Zo1gJ8FrFHg6rPgJBppvQK08fzr1gNpkLHmxjzzS+1GuB/MGrPv6iZIB1T5yUmT6E3k5Pf/DY3Y6
Vo2YMvQDA5HlxidGScY5FCWbw4JDPVvFtXTBdh1aBHeqDpZq3ZzACB6sXgi2q3Q68xno/05HKryf
eNqB3sNZFjyxCqTzZqtIupDbeU8A2Na+fd41gUOCJNAqiNS4auBEh8LAev0lJA6jSrPC9eQ714W1
QmP4W/Vy8bnsQyiTA2GFY3Rnn4RCzI8NLv0E4bqG4wwnDPI3q/ZAd+y0kg4RB8QURrI61Sj3DWEr
lpb64TXRY1Oabf3N1J/6Ao6yai/o9QNzSA4HUUaBxEWiNoidkeZe14M1Byd9UUD/0OwAbVS3sPGy
Iz4xqRr0hLsTcjlGrPkCjwd4QATS9YaVufvBPd0DNoZxTyM3c4OAUVubLVXTnu4uGuj7WHkC2Gkl
1A3wIStqmjeISQcnw4fUPpOWcHHSCCatEKePMXsa5InlJiuDRcBXaC4lDl3ZjL5KZOiQi7qMrYK5
ajN5kLl/gqP4+QbPX7Eju/vjBOhUkdbaOBZ9rf2WDRe/SD/ImZFU0W9VSPrcPXO4Xu9eg1wCJOxI
QvJI85Ul4Sol28Ij9zug1kpMuJ4p6QAC9XZ6zOP9O3viMV6xxIMmVsgzcJMaBQt1G8oi/VeTzmAu
knNJpDSNM5yDnur3LlOkY0++eqNHiSuez9GMsirYTuVyp56g3WhJH030mHrHZOsCDrvj2NQ8bT1Y
iZkD8MhbrZNIMDBmUHlFYerMr+fYe82d2q+p5MUhzL7icz0nliXD9dTlmhifBVVq0pNyRJhrFq0y
r+fkHzOdz89YWYCTL0SNOFEAhmn9MilFZfBhJqkJlpXBrZb0WPGG5smiJXH8zqBq0aJn/JP+xGGj
qSpCLVGwlZpJ3vcmEIwyRWxiMxwdVc4YHyjVj+zThidCop9PrOdTXvl5dq2J2WcRCNsbXAkOfYh9
Ay+YXNLxptvvRrcINAg21NyEIQG7EAnhBADUsXk0/lJ15e3Y3Q2IjJ+gu5VeCpbd20IkBsz+xLoy
vrpnK9fXOIcB3+ScfAkbLKRMsOIMyiuynNc0zxsGBRkSV/PM9PqyMwfAG5O89TWey7oTZBU1FmT0
fFYWDVKZUGRA1rbJjnErEN8TBUF9jvQIsbsgWqC7sRDKl2b3SLVXNBu5OYy1yJzjTlRf4+qYipfi
bHcWWXHigsq0yeUh/kHqmWpT2CbEr8yBD/kBbZQdFcImefAAQY/53NAKjrqGlWggwfvySMv0WLyQ
NnUj6jUuaWzr1mEnoTSpP2YvQK1ha86eLhD3lPWHM49ZFz1DgXb+loT5FM1a4WpFBKkBq1yuCzmI
Ks10FMH1UbVQIpXORSBllI3gUQh1H9sZbc5uMMCVCQ4ktcqXgIrmMhX+1MbUe7lSVI2QrX2JpSWL
UEE/K6gYtUIBks7ytoSr8mFwLI59eUORRblhGV67x2QGONY03Dxvv68PcEnCSCp1AK8rrffHXPgV
pQ0kbsIZ5mUVMStR+jGLXE5hQFd4xubAV0G1QfBhbPxihiBf2iTUDQGaHX9kE/CB3dHz2kuvTlDC
v0k/vJTtzjFI76JUVswoHyzWBwXCvqro/rz4ALlMlk6SKuxCj2Ufj086sudI70YHs8ombPsyIYds
tHMzpbwar4tsHf+PslVWl7y3nhr7SdfP8LSiTTRrBXK4wrIJgFl8oRD0LcUKBBx2VweQN5JYQw9i
xLu7QfUhgs9+EwWRNGqtq05vFmDPj23eMcHC+QMbgE7j5Jp82Xz9m+lERUBt+zLFz/rTs5pzQhMT
kznLtEI4nPOlrNhtEoR3cUeKQtHs9V80L5im+igPjbqJXGWlJp6FhR0zUAmUvLQyDH9XrjjvzTdC
VIsVx07X9Cwe3fZaqIRAm9sObmVb8GkiCnpbfJnwEnkZW4/gf4yS3KxzJwsqSGpuv6aF2fOeKtQY
S+lFy31GdWz2mCzmv2mkUvvgk/FT9JIH5EKSoQIcMRwbJq3WOYEzTsUttoF9gW9nYJe09eiuJ4Yl
Qk+81EGEUkqvCK4FKIaER8qD6j9y/DGrVrT1Hn3Fi3rWYYPbRX4xaA000H0P1kxCEczlkHbKrWXA
u1d3imgLes7RslDX6Sc5Ih1WDnNFXR8SbLIVYFt7VuYNKhakd/2/k8UbQ73lJZsNF5WUFRWKpbEh
adelAi6/E5WqSY01e3Fk/SmWWIvx2ik4z+HpdyuJkCoIKZYt2AEF5ibKMeig7l7jXEBanaW/FI4S
RFusQNMtSDZSmuZcClG/QDaIMGUjfhVHAoeCPT8SpVoAzmUpnQ5PASqWbabne8x3qx1z+WL/Jzrs
aQ9BZquiU21vuJE86BnIejn5CyIezGSAbQVIe5zp1Sb7R3C4w6D2bHQoUz9bNMd8CmP0Sr0pPyWW
lWbJNv3bBKjxmLMdTMR5FD2DXTiOgGMNS+E0diEmG2LO3hyldJ80AG/Rmsu5wpCu5O525bOzkG42
GFyE0LbZvlq8gS9uoktzvLP03xysv5L3CV7X6y/eKpvz3k2svSubVdBcVL1T3q+2UoVCBDPGKH+z
weK2d5kLC1OBY7eGxvXhIBZNyc5eXWPTS0M7U2zZNul/XHRT1TLAPPhknxk55QYNnbCRYD1IeKjY
2GYqT+MgwokEm+IlhGDEknBQ4cf/KwbzOySvjnXk+R15JXeV7SmpUkkh4/LuYJzGCI6uQ0GACBKi
7L8TTqwA1GmG2Ic2Iq4tnYGFCWBsjETTYKvNjwkXMffMTUXX5km25lyX7JbeU9H8ou249yG+FNVA
lwkbpVXOXg9iGoIME4QWyxHsLlKRSBWfPjxfmBNbVNSxDeOzHWsxcIm63yqPxJRoe8/0hpBfdkj4
RotNLeXN6pEIWQqdfU2V0gcnSXQismT7R5ryNubYaxhLccPMPJHYMx+XLv+8ky/7/CYK9OX4i8o6
NlihkCXvVCc5hto9+/vgCP8CNLKTY1yF9FwKkKyQXSVcmwmTQazIsbTZ/yi2XMACM8WLjcjWadUR
3CSOBTLT2ElsJJ5KIiN7Yk2hz3eiKwp7qCXI5UpTycuHM9cpjk3+XUfq4Y/IEhkKnpVZldQ2Ow59
LDffgajS180xeu6TRZpw4D+tohlArzbSvHPctoxu1LJMAruCCaPYJ1gnNNL6lx6QPUnv2EoEumu8
YkIpRU6OCwQ5OVflsidZcCzwNUqWI79nAVeVdOtFaoC++FrByhJFjnTh9m51eA/s5nOu/SESbWTT
L+PkWvoVQgy/mp674eynlfmiXNmKXxGT9/h8sKpkNFsHdTWWIhklmDDeZ0CnNzXsL2hhCGnme9cd
U9CPazSMxynjpvDmeRxshKt0IcJzOtt6/Higrhn+nEXouZQ3NTZE+rP7WZlYNbLZXYiE5mFwHdpk
TJUuDCZk8znAoPbZMFUd6GZa5W+duntV/fkyXqLRDQsne/1+VLGZDv2F1IaRwqEGzsHUigUOl8D9
r8LD7cLbfwoemNDn9h+R3VonrO6u8yoet7Fn6croaZ9y5QYM6uOIbKJ/qB+z0fqYzQFJ+kuF7PiP
7bBsEbMqOZiIXE+gXwuriXSM1xsihGMsUXRdc1sZgAkPtd/U57xp5d0JSNeLaOxds+MezIfkrkT3
6LorDLXFV9ti1+KNBWSDjbZ+QvJFDTSLmcE/8d9ebE++2aNjaNehfq77YmSaOLV3/4qGz8U+ZTM3
p1+OadaW/rww4iIz7s7QqezoAeUEE3oOvjHWr0LfegwZYiO99BgSvFB97H1clNt4UMl9xpxvqcEt
8PT28YkximPPJMO/Blb8BcnO65iEtAIPxQedCeWV2QD84N+svVankhjXGD1xLElFF3BFhgOhqTR/
bcWeBxM27FzlZ+9rsD0Rvnc1mp47z/9s3Gjvj9YRm9WwfcO/8eQRHygcJgyEpgnxan8QPMFvbutG
BCjpLxRVcD3373hXpVPGoXumSlZBcP+48Q4wHXSA6YeWAiG9qfY+dcsMbigyOk0EsesxvED8jhRO
JdK20UN1yJImsfDtrLf86ELknL5toxFNr4hkJZKkczzXfl1aPJnG7CPPf0KbJUatIhziNcfEokxj
f9sM+lzaDuLt9roDkBXTOWHXtubEimNW5QISxqgU/3WnMlZPXLVw7PkNQruBcfCMAxP+ZvM/drT0
bOXk+1RKhyMy8nmQnb335jUtnaprsDFw40mr/N0WTsfk+ktl61isQx6ZZsRliWB3YscavM8YdZq1
1a6wRzx+LduwGFf/pDu5zkwRmX51boYUOWbp/CE3U1sK5QkjsfVD15pz+dp6dDunn0AhAEji8XGd
htaTRLQDlc4/56miTv0hlU82hCVMuq34HSD8gxeM52YFPJomJwYFQpv0YH2xqMEyZtUOTDzUhY/2
Ss11hXxxnphoNQoHfnoXNqNKWY3QhhfRt6zh5P3BtVzNgxI+57Q7+K7mduLNK+eND6a4Oy2HH0wU
UgZUZw+Fcy30j+uO9ly1Fv8C2ms8Iy0Ig3+Jwwin69hPl3DO5sQNWqa5J7oBf37c9DXEBQgXOM9I
gktrY9TAQUAj0Zr8w/6SfJAiMJnbro2Z5IN3hq6unqpyAsTQ9RAWyfIfu1q5lCwPTdn7Zuu1JgFX
XpVV2vxs2mZ7ij/3tbrGzb4Nz7wbFgwcUPiGixjtjdxTxzueebLo/NEdxrxXIxj0jsrwIVjKsvE4
PJZLN8PD8kW75sAorwf+/IbXFnfkwIZfrUGlcwJ8Lkb1VaMuCVod9lJqAhqQ8ihmM316yQlXFGH3
hSZmV/DPLEbLc7O5IQMVRmF47ruY/FAqa4NtwHa9gXHkhdiZb0pwBYtRGOdL81+VAFgjRE3QT5MT
pMV1MUQC9NAdEwLk1XpHiIqB/ihrDi2SE1hsmhB4rivq/RECeNOkL8Rc1TC8oh08Q2EblyJzRZC5
tzN1PXRNLvi13D7sBQYTYkl2EJEJVIO7/Qbs+4HolQyrdv59IWo8bKH0a5DwCDIR03MtiixLVKB2
e8l1cx7Fa2ZCitY8yccKNf0UfrQjPeF7V/hDPdDnqAexf+LgSEqBc0jH5BIFyz3ZdYrfAu4UWM99
rd+nVkblbwOqV4BT2Lrtde8dGSpRePO0KASeK9LjyI1h+QZ8ew9gOka4z3BLspODBKQRyVB+7mei
Ai635/Oc4ZwlJBl3+3pVz1ApBusCpGCJl+rdC+tFVxZHsXYVhdQWoATJlVRvgG3kaTmv/FbNSPjs
r6ap1w/JhVv1EE29Gm9z7nAN1cHOHN3+TO2VxZhm9gzst3OAEWUmhwswCxTILo+sm8v87p4Xgh8Z
QlJqtzd4Xd40XqoOYD+vmmBGFssgr2ChAT1UVVj68tQFwf8mk3MJg3Cx1b8RLM2ZIbe02EqLAoaI
ZcUJrYFLzVlUVb/CmSvQfKnLAIuT6axYQUBps8sJkbPRdnJPWOWAsLchxGJbInMkdcv0c/+MTQ4V
WkNRhpV3n2WOpCSOrpNnCOrvUE/glFLsjPdjzK5YGMdjoV51SWIoeTOCr6DfHEdnqfXPUCHONskG
k0Uo+M4yQWXhZeAsrKyd6BhjSxJCVvCl5dXbNeWIk8I7iSOsWw0WgZbZdlj5sL6DhK9z5mzVjfdL
8Z+a2Pxib+CrHL1bgtpvPXzgv8xzRpMo6hXPX/oHKWoubKlBQEAtDQKUVmsUwIBVq6OLZ5h7PR5u
mimr4KosbImZh2x0U0Huy/g/IAin1VYMfgylHZWZGVnjzhO/opOvTMzmy8M08k3X8m4xR1U7F0x7
tD+vzr8rkLdr/1VG/WHFT5WMc9Q6LGBleeDHYH2qU89oMnCq7C3DAsLq5dZTGkhUGwz7F7yAJoxc
0EKlr2hh6hQLar/NWx00x2NHU0TmOi+v5BrW6edMUjr9wZIRVa2TMiuSXgkRxEhz0ilo0j6i22Z9
K+vAjKe4SKLv5RI5iUhVcc3Dj6tX+rFRBovteA3OtsyX0KGhwil+mj/AlkKITfgMjQp0EY8XTkJm
h6lGO4eoHz13/KqP4Lp8E3N31jJ//tXzqwzEO3Nu+YH9BFKLbp1WvM5RttPgZKrGwrVa4VlDWWqa
ocwyy/5pzrTk9gf5jaCfE9MaQg4SQAit4SJlaTy/HilXh9Sw2vfNyC3QZ2KXpUbqXLi8n//keTkb
FNEqILGzWTiZMEyFCDeKuwfJg8mwdl28xDLm/6Nm/cJ6h65damdDhsSrpugvBzCazwDfXA2GvYFs
gEnLgREoiCER+iuKOWMlN8voDmnptivOaaN5bAQLJKQknaVdBF5ZQvlr2cEi1TeQm6UkQ+9kQJ8V
MbifCY0hPwA81rl3BqGaeiXHn1Ta/K400YoNuQcA6oKVNsabPVwBTrENB1tc/4cNUN/plP6qik3T
nxDekwvdLsJXW6FZDsriXlSiK2PTwBXJcbJzuOcDDuKJs6f1bhnKNQw087Ww1m8wyYec/Ut+Qp2e
RS+djraKlpgiVAuU2HUymVdJjxiJj0G3a6UjdPS4SCDFZtVlhZPpO8e2NbTJWhpOx+auyNe1KOta
ds/w1R3F6rrY/XaxWaF/27nDig8WA/JNzeNjpAAc18ibCe4VFvTu/siOmYGyz0NCEe9yxDrHhrZo
f29UQAW6oFltL6GhZtnwCW6YMaSSdUm/mUoBwh84v76N85n0/KIpf83ItGP8YIox7CicgS0L6Wmo
SklBbN2clexgs+Zas8slsrzMhKheu1aEPjSw65DVMXxg9LG7f4KykIPR561yazvsbWmPpdngTepL
Zevjzm8AlbGYwjh4OpE9lRDxxOs0z5SR3PH8IoUYttE73AAc1nlc+Oy32VVhgjr7Ezzz8f7NNovr
rUxLAdWBAE508oHb0iHcaBbM2UJLjdUmsRhvpa2j1Ysoer41AqYKqSLV+oaE1a36w9K/XrDNUYvi
8gVdYVFtxM/BuyNbmMv+k5SSknEOvQAkjdJE+O0gc3xMh1ks8e6uec8ECXM98ewY79CU33dONcTK
dnMJ4145dn2nuaUhM02SQYbP+sY0nP+tG9tqFd64YzEbzWgKLR/Iltl+Cl/HRK80KTNySJZIowg4
53M5QPWlbQn2AdniH6/KR4JAhZOPI86DaVGztUPyRA2romRj/M8Jyhv661IwUYRt/SfAQloNHeEN
ysar0Ec/22owQVGST7oT9qkJCBJaCtpQNQ+is9VtRWTsPOKpw3+3imze/VJxUgbwjlViMhALmJN4
x8a0QaWn4VwLjm+ona+sZAPjZ/XP4mbGzBIlHOsZcV4MnacPDAN7QPMaui6bM/d2+A9B0w0GhCnJ
M2++7XiJRfHds04lTBMeax675luZavkss+nru+d//Nua31XNg8FMfPsBu33MAKvYKKls8dwONyY5
4fvbxgZxDOv62buE7UpUNs0rQOOJdUeSBeLgdrucxIJcyZaRYEKuPhpYr2AX+iYeolmRAVJ7AAO5
URLTDkke1fU+JrfM9R5A9WC345zAmThWv7ng36qDvhXX7Hh2vQ3r64sefqbqqCEda/BtXKmvz9Ws
uL9UR8rtsLCf26sdfMirxE1f7aAyanDOqZsiR7JCK/sYN26QLcZPUlyWrIYoP6yUIRubYq/GvR4/
EA5jwn4uIeYceJEB88tjaEHpiQDZj9bW/7zN7EjkqzoadqUPs2bNHo9ZmGmJAseCKPWIPvLLASWf
/8GPHdzKL4YpuPTleONKl6+HWtbkOwB4PxaNK73fIZoMdLtRsyyMgXFPn1cQu/Lz8O0fSagj0B+z
icCvVfO6m5fgZxqN7D4fibfiymroKrgtkc88A9iHD7xvn+SZj4riil/OZ0LeKBD4QSNY4nQAxwQK
8DuMDz1xPMS/v19+bJOY6N564DTskgYxHkAXASAug8CdeNg2/NZSsQIDwNNarSuUybwB7Vi4UKJl
Muy7IDm1KObTckHh98bOOeLxGnqMwcPwzE3abiU2uDU6pBcWkYomabezK6gnc9q1DsXARkvW4HHs
Pnp1M84ZNV+YJmByUqbZHsyFK3tFfEwRRiops0+im8pYCAnSyORWfuwMvxj1ehiJ5PVJnFYicyg1
/ehjBVS7CMuNEBFIIoTy2nZgmp9J3W8WsYngBRclnX7DJ2NmPxwhxfyeC7/L6N+WIakyiX5aBLNK
o/1lbQzb9f4MkJyb8J8kQGixJgsDZKIhew5NTDBbxQqnsBCiE9SwSewTEfPF0Qt0i01Mobev2kSU
zXTcD//pxux7YNnlACqJRuPX8c5UNRugxY55l7nC99qrb536twJ2LLokGU3o/rAeTbXRKopiHHJ4
a0jw1817mJmw/rrDN4oPdrKbz8ZDI2xOZs466DWUMh0UXWGqu6DIdyDjHCNI439zdUMQzWPKWodY
e52JX7tbmIPH6RhewvJizN9/FKeAxQq1QwkIr95RZGXfNFZ6a0Kk2UFa4QyB9ekUR990IzauT2X2
Dnshb5dkmBohzGXXyhOJiF4yMR9YZCYdxSRecyHOrO3tn0Vb79vEdt4zmIno1iS3yw8hnBICuLsO
2L3Ph43wGCsAENBTKt4rE/i2Ev/SnVj9HMFyEU2+y4BGpQmKU/w9qu9EVf9SyKIb7MqH+cF78Zup
fkVY1FEOHkjQrEx9UDpemHZxGysevabJvxt+c0k67OQW6mm0OLyOzWX7uI7lV93O5KYb+m+ieMTu
9oUSHOAq0n46i/WlcLt7wRCF1JhAc2ECErYY4ANtoopR0VHyRhlalP3gznJa9J0GK1qbxm96oem/
Gonkc2DFcQlrg/Oq/h4chiTv02x9xy35p/GxTgLXYWV1kUm2W23SrKnFxq4hfbMMgxDo28YruAHQ
j0irdYy1sswDRHviQrbbwVroPHIenMFOM+iPbp54Og8tq3nJLVGwFKzj41NBv33PsnXlcZCn6Iu+
JdaTyyp6Nrg7oHyT8wo6vlIsHOeTE7uWqe8KuPUDuytnMAMIFTNNQkQqbiZ68hdy8E/t8liDk3Ge
dkf37OumEWJJ8/MhXXU1CraZ75j++VKijkNE0hvNetClgK6kywVn4+QAN+JJ+IDfqC5ruAyeyDhn
j0Z7/gnD62G9KD9jQyMHrYrFJZN7+C+8kqZBUTN9XIvoQz75nh9e3RwIJVN99PlVbciR1PT3ELQ3
Do4FXaBVyY/x1H4YBQVkhM+hcmrT6nxfhV0Dp1yxZHSM1GlRTmo12+LuHfY8Z8BkluyRvWg5COP/
VeG9cuSIOH0XKUDI5U38nq1l27UJosAeaeIQIGkF6a7kkuMzkrM4S8YcqwX2z16a1RDh1G/HN5n/
NcPP2kZ/1iFIvNH//0lZq55sPhss8R7MUhSKuaFck4d39nFdovYmRPbUGxs9Bb3ElQHSfOIhzgeP
JIHY1oR94nn8ZE+RIG+AAh8ytJUsuucUGs3nrfsnL9Xj3F9/AOXVoGbpsiFUd7lkfh5N8ZGpunIC
7RS0AkoCQiW4RtlxaoNR+Udb7ABkrjvsw2KSoL//Cz7m+xH298yioBaqimUWiBl7LQqGJkvDkT/Y
2dXiUDmC1hisTpbQDeGRTZHv2n+FcJf9Y2PXvngixOA3WtVQfQBFvVyjYTrF/BPYNi5XL4wtPC2l
KlDoqfRy5L4BZLBXyMPmd3ZhUbMrioQ02rn5PA16pz9VCKsOGFNzbgVPVaomY014Az+zJkzAs0AH
b4NCK5pSb0LRlO2HWEUeUoV4MVCZZhIzL5bkPaE24P0d4ULLR5TNIcRC+t7t/uD+wHdJeczK/LnO
DQP7fg9Y9VcJKjlh29O4G01YwNzXLFetcj5gGdX/3W8tzMlXv8pEmnY9vRJGA5854uQjyFJJTSRV
9RIHjuDA1kbk/8Cj0UGfAliGnk6IU6jAKT9fsBt8M3HqpbfbVvv3zJIfzMgfK/qOISNJztOD6JV8
ALDjRsHSs1w0wti2YTuPR+5LbwJliCt0+KWBU0qI8aDflEL9ZNd4M6B8xKEuiEl1XtS76Sr/9nDw
SIvsP8SfIeNhLkM9vVIEVYSXLzUCNnSQzXAiNJDjp4/EeyOOtHW11GNondv2NxoaXVM2m/Vl6XjJ
fSxbcdVz1DVTKEaDMyVL1Sg2zdR1UXKOoORqAwcLQGKm/CJMPGYs8ViqzcjlW6xxswkXY6h+Mu5Z
dDjqda17Gq2stK/GwMjJPc05fFKg1beYbbbh0lbb5MEM7KiBoQCrIm/C5Zvx19B4WjG93KpZmGJo
eJGZpjKtw0X01cjbDEYPsYa2zB4VLmqiFnhY3mlq1PcSBZhpcWDdBugq6gYFQq+VMXQhKF+ufREe
+BFNuDSOhC/rvOGH7lyOsFLErYNGRUaSkEakm2iE7mi8NaEqhuHIFTNkBFmWrZybvlpiSsJ+92Mq
7E44zJsYPjTPQEX8rzq+9A7t405GWLtRLhI0HvDpCqT55J6vi17LBFr+T6+gdDOTfQ7HFuzIuuCC
K9Krg3QgNrkfQmFZnGLZ3wgy2xCbsW687tmxkBbIs+HL7iMez34jh63fn77NNYOXfbb0z1A64g3Q
GFbyVRkjANwj5BZA9RYC4Ijar8VdQeRa1T7bTamZnIUnJ4hxtN90njuIENlzUvhvZ0loDT1DzrLY
qC3NOR5WqEdsPJ1Psph3TA4o9dgeJ0MoRW06eckd8TIq7suRgQiP0E+sSO3ROeFZvPFCwNrq/Ona
fHBXyCwT7u/5qTnbLqSp96c3aWpWQ/GHbhiGUeWG2UH5ULilSo37kZGfZpnWH4VpQhzjBqQY4hQ8
XESKIP3P/ii1stzb3Zz2zY9qch0Jhk0wilEnKAtmY/VTFlrGvTlTZ9rJiSDpqvAsKKFG+xXW3ohj
HmEeF7XDPS+OAEEJ9Vol3EOAYgSqVRTieCo3lTZQCQECqasTOURvxbotjkXaJCBffrGerpr5CIvM
rGgB1q6YnAafTkrGDzypFuGp72OLxnhYkcVASgNa22Aw3W4V/HOIifFeXtegO7cK1R73LvgFF/Qq
K4Mip73qhkVkVcWayENLKn9RColx1BGjowYckHRP0PRsXLu8YbefA5BlhPBVjMIrBd6LC+pzcmul
KKupnUwfbtR0hifpxd5MWvbtbND42VTgQuVEZm8ow8+sQ9w2Z5s2eKHArNLmreoGibg8CFIwzWYv
xuOOK5aUWeUJ431lY7Xw7b0k+iIVXbduZ1yikIWONjkNJX6XRQ1jgMiTJfw2NqtQ+NXz2TWRCL2h
0QC7qd9NOBJroZTDJdtgcPqMm84sNSm+51StRhjYsa2oSAcP8y0hIr2U7mnH6ghwEqRpa4Az9x3R
ehHS9GZS9C4XTj3E19EnwStr9s3cISJP+uyyYwNsQK/ybIPgmDpOAr7TM7LTz5cXhkk9mNWibg4x
gcuq08J3ElyAqwY52HBmJVa/x1G2NX048kcQe0EH3Ocga1ukbrz3of89Pz5Be1fH3/eeTlwPMC+1
GGwYZCb8vyozVTa/3uV99gFoBSA8JnY1H0ZL7u6UsyEP9o/MW+Nt+baYDyHZe8zjBk3Xfdts5RZn
lHN+L/O0ZZ04/J8mCvX1jXAn2W/mKKoXgJcLAzTNHdJIUi/0WiOgWLiwk9aCPIeCfa5wcxzSQfuA
mHjLUvKDyw6fv9Xzebg8ftcrqZMpzKc26zv7OzkknwsQycUS1XOHdvBeSRvfW9GWL9Gdo9216GlY
w81S2/yQWTKmTXIXpfnFLbLH+KEe+W5BTUiz2oEyKJ0bxPubjVJ1mrF+ihGxL3Qc6pPtGsgiNoEq
hu4O2xgwrPeo0JtDHPTsVpsM+LhQqS/KviI21jvdCKTXTR4Jdpecf2wX3GTHYgBNZjINMa0fA+Zo
bhVGQp6AZ86z0/3OblWsJQvz/zxX+d7zGsjhP0PrNgULouQlt31/Qt7cnTcwRBJNmGhtt+jkjEOm
d8e6iHU+giLw9i5z5gwRBu1b+GQni4sXMfHVlV31QkJlZURNd3eAOgYNxdy++mTfdShoY1J/1spW
ocRKcAY89ZHTgvszklJXqyjiO4P40eVxNgpcTczvoQUZnoSRYONY9rTDb/T2waz8QcEXIzzhvAkU
eG0HqB3bzkCv7oz0cl536C80P1/1Ko6Cw5ne/wjEakj10hWPqCWTfNliEd6TBaEwMyYV1HB8xm5E
XIAHNtfzm86DZN06xOK3vopLCRGCuXOQKlH2R8n7ovoSJc9P0osglyuFaWOs9fJe1MzP8mko1k0I
cZpl/c+lmf0iU5YoKbHY3rIoJmyN6NbQ2G3kx/trqOCFDPEJj0qFwVyoY7bklucein24+0t3hcKs
S3z/F69a9nueNt5bsD1vPl9QAeqlcoErfiugyr3zrjNLbGJH3FQlQjqgMxmekiUi5b7CaluwjO4i
NdfQc/ige74iQzVTh/9HW0hJ+5SLOrfAFmZ/1daGTxHTO/B5unzOTzHJDKl0gxM+LTLA1GFLr4Q0
opKZUNaNmGE4qeKtz6wkxKBjDmiyW7l6J9m/QEoTjJJ2TgfCVZadrNxy6slj+Ia0AMEpyt+vLu9H
Cyi9hiK+hyqTVTZaEcEdVEm5pQh6EoxyrbEVijYtw7/Qle6+hCFdf9kJttQPijzzDDX4TC2/Zd+L
XdoCadL2woUIcPQA+O5j0xOo1dD3jYVd1O85GfP6UyBs7/k2DDLg5cNHoO1BpsjLDneI34SS0BX6
ECXIZJHwBy4pYZy8cib6oUH1V9j7A+dworjrIM5U5eRZp58YigUV85bQqoE4O5X1Ev/il9t98W3d
fSi+Rb1w1GWB0VFbgk4cu+GQnYxGgrqc7m+db37M9GxQHzuFK3NqZMJvzfzCuR1Y8cUE6t6eECS2
EZzMePKq+P8gTsijk8ujpnaef++1uhjCXNhVWHlz09wRA/imuMggNrtDNPBijtwmr+cEoPXYrnrC
bqLfvt76Fry3oJhXQlO3ZnJhI5AcWSQnrX4p9AAtDCK37aQuRAxwM1srnwoV7TdT+0afFz3+Pf1g
q2/vpGROVqw9cLts1Q4eR8/4CIUdJy8zhFfdd6nQtm+bHDi6dIIupqEqdDgBraO4Ztr3Sadz8Zyw
L4ll2sXz1SyXI4m/F0KgrZ2quUBEn7+Ykjfyoo9738Pdk0wvQTSVjH4Xvig+fASb0hrr3XC28YoX
8Ch2LtiIRco3oPNqmJ9zGFp1Hbq6isCyA4TS9VTrJbWchiM/0r8fhpaeLeyMfn4daGlz1msI8mDo
8jKfRUP9olLHCFUiwfeztOufTBOQvkyjgUyUpjd6bOYT/36E62jiuWM9hYJZP6QNsk23Sivq8hgu
vOmVSuwqLFbOqwf4+4e9iqPyV38QHzoThYSREtR6MTFDoFl9UfawFdWgQ3ax1VxLvs5bQ2+fb55W
RkTuXwqWhVf7xT62lgdTHfLWiGoVPi6SDPoxxcxp+hy8S807MPPHRjh4jEbLZkOZm+DrJqNYIJcn
7i3IYKPfuC1cHGSjAEL+0DG83lCJWCLqj0PPyGtL/lr6AoKZ2OK2K6YPpEHv7Nk3HYlnxOA64Kbt
MqIDq7T/NSqMXfjbbR8mYNG7gsRqiYJjhrM8wNbM7d8sIIUJBW69j1fiodNbApFMT9CMEqM9qBlb
drpiu9GOcRW+St9D/0yWKElDNU74xpNVzPUi/aVBs106H2lPrUzZOx1h7bIDgI7XPOXHt2RNurdQ
1C8FIzz92Ajxi6dwPZvbA1GVPnvd/2xorCrGcT/YEZOY2Uk9sVebQqgwZ08qf1Qny1hzSeGYVW46
rOePaQEPJf+OYaPwX+Wl/gzHQUrnBBUxtbrqwOv5DlYEAzGc8CB1g+46NTD499pKEgfGDRQWGmxs
124KtlTWdR+bKpORWfOpQLVPJIT2AI3QRM8ZgV9HOzaNuyLChvNj9nMPw/p5lspFAgk3pBN0gL3O
NsrlZLV1vE/2/PGzMevfRfqrNkwJF0x4sFB0zqzRQ2/dLl1stLGtFV2Z3G8AtL3tjhqidZzoRXoh
Y9Dw5nTG/eEDDsL+RoiP5sPoWjLKO4k5FXVPLx2zox575Q3LuI5q0TY35aD7UAuOGn49MVMfHLEG
zT9Z09/XHfccHXIDgPqzVjFeSmQotIU3ShpZ1ZZbsXqls9A/lwzl4FSUKu6tg5S6mCDlpbsZCaVY
8O+ikav5FnII8aJuFZle1PKcC4ohVwfA0YWCzPiUE46oqLaN1r76tzFU/SA9SSqeOiTVzHawk5sh
WUPnzHbA9qNFATq6dAr+6/iHhlP//vojkKIjavFwOcsCWVLMbyMYFxtmuKtJq6fBwNJKZ9bhcKfZ
36NcC/R5xbdk9vR4MlFcmIWPvibDq8jYCNr+o/t8/Z9IIbWNuPqczeLGwEwd5R5v7WYW5oCUDiVu
9kP6cupzWSVljTkjPcJ7CnxVV7ikwqtbxKoETUGxW2uZI3xfCiW9WDBwaNeNCTA3wGVC9kdlfN9L
mEJMCso4JbR5xOyVXDDriUPj1PDUMGtXfHeSGSlTXu2wkRYeeTglRTvv1RmiP9QMLzIfQXmQRy50
XLDtQJPYHUDa277T1caQDFHvvEt4W+HkZbWo2bpCpRX/1MqrZ5ss7zTx6owQGP+vo+ejP2LSxV2o
SIJWbQ9cp1C0d0FTsVZLRNYd3+81mmwRwCw8H+ByhICcO+2P/bDWVianU3iK/WiEY6mweJE/RYSF
ehckyPiHXjZnWeU4Lqnk/kTAy+QuZ3Rz5lVW/i20WVyJlUhza4WvhmVD6o/2ZhFgp99ulGOr6znN
vHiCKxw/ydQSUujDG5VD01NxvAv0tqYTk70EDCNwrDpAwZm017BpL64U9CFAGYarASG5wR1uYIir
Lo2uJ/z88MdeDhQAcSQm3m9Zwyd9tU3MuZqSjBv+M9/mpKv/3mD6jFfDf2nMhXXyIHLcjsgzwQPd
o+DixRif6fcKybw9oQv6lDzooZQL58XC8/VP8nFAC03FZIopNF3zrD395wZOPZhk9H0mByd4EVib
ZsSn2F4zJ2cFnOWxXgNLocH6boN0agvXGDZjVD1C+uOH4N0HNmIjOFhKIY+cTvYclJnu6Ik9vmh4
Pf7oYKG10g8NOvODjg+1sF8kcx1SEUW9fl/AOTIQIxryzmPcl4lHl7FW7LaxwWJRo7UDMVZKkESU
SkgEPetXwj0XOtGrWXMAUOUts4LkTIy4RU6mdI30UoMDmVK0nqklT5urslb2giFHggLEmIVhcgRd
Ozb+ilVteYrL3YHBswcJT11wNGiQXjko4HvCkAGT5BX/h8RWvqbM9H6LnDzL5TVDn86wrMtKG+KR
+dVhc5M/jk1d0iKeNwO82xaPIvfTmrG3nuxfvEHK3awJXAgAEZr6ueaoVB/jsrVicLuMASFnB4qR
5GZ/LWcEU6/6lw1igpipprdpURnHrPMP46O+5aVfPIX+Ct4OY3+4hdKJU0aNpiudV5P1GCRELglB
PoxYUmX6fJvBQ05jg7NaQGuDVmqIw544PGr6HxwxLFq2tsaHHZBCl4u9jgYk+Qhrz12yqqepe3OZ
Gvk9xCNsjwqzL74HAKMvzW1UgAbXzIONO/V6aVJf3bHOck4N+DiPf5ym1uqLWSlBNcwlONp6RIjy
GdzuLoGGHoBR3aTQ2IvTjR9gbMINtdtG7wvH8HUZdvtUqCK+lO1prqWv+lh7CC7hiUIid9Ibq9US
Tq/K5Pe1es7hJQs9Rmk98A+pNhvQ207d89MKuG/SPw1MwhJoLjzYp45mo9TEJ2kGdffBrxpPP4Yg
S2PoCnPlJHxtB1MKlJQQOgIPKCyhB978d1+8uwhHczmbWRcscH/uAx27fcmkfurYOY9zj6jiPOlE
S3xT58ZceE/gg+eT0u+JAYmmSQnKWFbHUWwpr5hV8FKYuQZ/2EQR7Zk68XNCoUhdr5fENDwn/mBf
eHYNdXTSgLyPyA9mEwcPDNQpjowkZayVSno4IcXtSsjSOAo7FxbVZEMnUUrJJ/T5R64Vp9j0gaLh
rD1znpsNID+13ZXg0IxN4YL15VERKJ2wOwwM2ubXIKH6eYbTL4YE6brxrK6QYTUBSZryFzVALWLc
jH95mISxtSJ+xaymL/Ng6C63IsHqTionEU8LTvyOvOMldxELQJBuJEWpefFQXra4l2LWqpHhBUIS
UPnB8qAScHJjDgNVjF91tIkl0rvmbwxMlDjVv/Eu+8aCBFMe6PuTSckHFcy/xtzK3fA3GJnQ/NSl
eHtJbbvvdGGZsXYq4DTqKlN7mDwxPsZgCg7Di7ebySgHT7xiBE+BS0P06UZnM7fLOcpMm1rSfHum
v2IEWHGzb6PHON1pu+OPQOkbDPgrAclSdrO093gvjNoGFu4LfZIIoGkohlDdIMnKdCNCzVf+AaMc
5z1hXZwB4DpOiDWSBjJI/5J6vs6NJGeW9p5/rW4Kuz6V0CrD0lqb3R3PpgGc4ErQrLqdoryxvUKq
usoWjhkDYZ6U0m3SAfHJ6HsPcAtmERF2jDYCNRSSO6YVmgINuq2tISfdH/3PBAYrL+DdYZqKrhKF
c4sMhU305VUpwUE+BFUIw8VsGEvv1heRYYBw5vHifA8VbT9sasD+iHyFiREz7UEFh3b5IwnXfmlj
yiZ70OzZKdoHhTVj3Dti8/Tc82LorymX27FIEhzPbF+JINnRv7qRAwJ+inm0lyyLLF/7nS8QIFkl
9YPljmhDyI750t1vAems/xD8QGchLncR8prwVDLmnnETTaHMz8tLQsnObNPM36gD27vyHQXou3ur
eUrxcGis3zAQAK7TN22XfbNMv5FC2ldTBxEOCb4MN1zN4gF224Djw9k3kNmWNr5eFSluX0tPvyZd
iMsmsV2B9HouVGNb0OytmszeGA9KYRlvXaeG0rXdxBEuVGdfs3jChJwhnDtrHvi91k1X/Goka45L
EouQPe78ByI9tUiuov1bgW5u6YPlGbDffdrucsoAR7fvMuY0Y8RlNt/Rca9077VWumCLZDbIer66
ERgyJH7Sn276JnXvIokvJjBVbyCkVeA0P2yqSzRlyfB0UCSDTvvpEI6L6HF2ovQs73coJEjhmz5i
2VYJb8zUtco2Mwmp8blj22Jli6YH1lV1Hm6nr9y51dD/tnwkY/CLsPx7//Rx3clf8VVTSvK8OrM/
NPdLEYuthlvFHqNAh6wSEyOEFLJylte5O9t9ulb+dTc2Av6jTeRqOPPw6LVd4Fy2HG8vc9YPbwW4
nYMjadrJm++f1poNevH1sZIlAZYrF4jj8V2nJJQZ9rl+KhlN1P+qm0iJcOvcppOfov1fjarH3iNG
3Nz1OTnQCxicI8N3Ch5XugBEZwmYCR4JjHi4YgQsVKDiBeBk74ALkv/iaJekShh8pYpXoPNge/1j
pmqaQ4q6XhthsLV5z75M7NJ1qte1XfjoahKhJlwQFCjtlHUPFiknY8UOxFFLn1dH7fehPLjlkO+E
DyIRe6JwaL3/Ni2AS+Xh/N1AN8EZf2pe5mGXnIIZRaAViq685hkgY10mfE0hr9L6d1xcCxkniPSs
+LBLLrGKVnQ32PSV3zwOUq8tru16Z90XZevvlpNO9PSA0UsSSBGwLH3yVLtZi3Dvp8+CUCykT7Mu
nvpgdbzMyRFswGJfl+gNaUsWMF+mB8K2zTT+jo9/GPB0kul/hUk7ergSh2GsWmUASVL6RJaWQpvm
z8Ye6icdSMKE4ZsyPJThZDivv2ShlHs8GHs9xin3myakxCxd7azJQfj3OzWZoRlPKRP3GNvpb2aj
7ipCIeNM84ioLqnlaqOoTafS+BYLouzFDISaQnAb+dLKVehLu4m7nUINe2h5+YYwo7yWaN8MeZAL
u8HN+8mSu/Y0RGDkSVhHCIf8DfNQbNmrchYcIiCV65Z0hpqFVUIkuUoLmye4p+NWP1OxUNLiInfh
sgXOyWdBLy5qD768iYTp8I+d3w9JZKpDYcPkgIb83WV/CDX/fb4KlhYmDeAz4p+z4zOpA6Vf2OXI
bvu8C9Hx0h78IIzLBn0oMyNlO/EAdBFgfOo1221kMTJon8YylrMNSmYETHhiJ+WvubF4hqd+UwiD
ShlXrzT3xKNqp3zMlakGdsKKiSJ7RDWYf5NWJHjWxBEq0+/CyvfhgqzsMvTpWmsOSEbSAmXJYH+V
ZOcde8s1WgcEsSOtJiZwcpWO08NETzfn2JjLZnYtEW9exOv/ZzfzTpSqSwUiHlxw8TrBVCRozBNj
lKW1tiEGoQCOr6F/19gSkIiTYMD207KrqUnV/vUuseXrJbqrQcgBgv64w9JFFWycAgbH6ATmABda
JmYZwU+ybJyrCw7hAVlNm4DYZSxe2PcI1nq7q0lW6mw6GlCQb8iRQ/JInSe4Ct+UP1AWirLaouuH
8+R60Dkyp4r6UnzaYklIScIAurcqged3UAA2YAA4UY0gnITmg6T3ux/AX68ppYscza2zoqut8tjJ
66Em/euLXV06N1v2OEiTm3FoKTydiq+vU09a+KCRJF3/sT0H2trwNdEAsh6ctIo0J7qv/0zEBIgg
+W1Y4pSTQ47g/tfgXDKveYB8ngL9zKDMzpVhoaaXQskZennOgOYQ0W2U85OibDcUKw/tbjQfWJQy
ZofqtOuW+E+pUVAxsJLanF8auN8InKRyZABICNqmjlla73r0g7gcvI07Vn1artFsrmXRCMp/GjaJ
Cf8Y1CzYh+3kXBNy5udquWNPriwm8LuK8kVgVSG21qNQXL3AlvLvuzHlaGkr7CnNXWXEIM9Q70Jc
7x4+ixix8W9CBuv/uCmcvftOejRrN0L5eVHIueH4cDMmR3FH6qCK7in9zx1UV+mNdNz2Gtf6+sXZ
e011U5H5n6Nj8W8II5VXeTrHfwqLy/Z/FRaJajbwMB7fkCDI/yz/tQuF+zCdNQm0rC7eN8N/21KY
0QyY0R0rzkicMi4nb7HuNlJ5kL5HlgdZxAjgEgK1uaVABsISZwAMBQ41khRcaqUxF6C2GbKypw3z
qPfQAPKxKC56nty3OJszYt9jiVgYOd7HRcK1EU5pRXcoGTRIbQo4FkzsXI637WE0yKrfF9xRHYsR
VF+KCn7vwhEwKessu21Bg9y5u4H5pUcBhiDWdH2CTCXu5lzQtoruzMus+hnkpmAGrmRcALI2Gxon
c+eXoLGIApt34oDFsSjv48RRKoJfqQhnkDOpBomlZgs/ytDYyL1gAm62v2vK8hcTYjEpUP7saGrp
tpFpqfZKUsNsZj8T75DyL0luwabFR/gjA5H4pLLUl7WAeJ5Fa8XiN0l6yHkNMhtVR5xw4DasSe2W
Atc0tTnKJ70cIEISuUv1/xsplF4qOV2INbs0lBGfr4zVixOQ5Whq/n1SlMj3PZJE1SBZG3pwTqrJ
0GGsWjKWapMV2/+gpgeEpqWtJ/0hEapjspB9BlDlBTXJxjmJ77/XgkKrCcc18bqf6OPypG7N8573
GIZ8dTEjvXeHKwPoG/QBCwO7hrFOR9jxtIhk7nkZOeVsGsLryIelyuisPnKS9vodMncqGQp+sFV9
ho2wMWbIWVMSGCcJC8BC+zaSRAKI05S0wMSXRrwgsi2eYFe2Dk/5YFqAVSoNH6zshyl3/h1vsUfb
jKtfP+cb58SvI55ghbojrKq+vUIgd//0p3tjMIlzj8aPgryqNS9oT6kAkYAyjGPQNt47TlOY6NIT
6PBkAd13JKcYyCAHelBTukWs1D9Tn7h4uqhyPgv0tX2WQggZbuhl/2HlE7oClaNLdQyYYPdAbNQv
3zLITdxqVh2nfW03xWY7Wef27M3dwpPBUZEYecWAVA1JNAoyt1/ygDEdlClncYs3yykKKcS5JOw9
zrospz+TMrXLmrC86ryndUCzZG1gX9TdboP8BN+D9k1VNpmLuzZfj4icfD4LqDggTpPBET3QAnEF
DKC0fqr0hOW3Pn1oQxLaoA1wwyFzbmW6ATabs0jF8ul/DnQiFZbofvk0ljhAbJ7IWrs+tYxEgHpC
OQJm7eNdU1heGgrLxDp1H7rc7APfKWYjvdNZFws8d1lghp82wRAuvvR99Pf21ZFUieW4aZ734pnX
qE8yHMZ81sATAHxoy5dWw950lE5lpOlhjXmjFdWS8xlj07Pr3mNWkB382sX87RIFDq5XUa1/X4ql
mAVegoRGlCYn5gktdYpP57fJ7IBqka1ODvIkgbTpd3YMhEvfuXHCf2sWTXJfgDXEncJzQ/7jQSlX
Lu4qe4cGnkqcD6tc+MdTY/Qdj0cJXbLAF8EqOaNdUJ4ZhgS8A8QnP6doWt4VhyK2bXuaVW8Li1Wq
jTCJAn0r0B/mwW+XR/XeOl+rk0e0Wgh6Tl7VabSb84XDTNXxCQLTqMWImQPg9tU8pwng+ilk3j/F
agn73fUP0AYinNq67XhIW+N+GFV3lH/67IN8WWn6DG2EAosEE/S22aRa/WunIju4sVeoxTcceeBD
wKf8SVoOtFj31HL/M3iOkvXaEOxnlGrF3bfe94Xj8Hc2zTd0ljH1Otzmont8ZL//byZx0KdH5FoB
yCmUg5s5fkQiJXstGGCTzWXsCpmbI1G0/zSEmqFBiwY8ye1qrLcb4A6tVltNPERTIC+kQaC9Bn7L
8X2ZjPHOw9VGlWPN7NsZ71nBx4O7EiffKtffUkzBnnWGnQIo1oHjJybcbK9z3OvhWJwRKbf5ObMT
n2RkjA8HfO9Mn/MmPr/0WQoj8c6nwNZ4NXJyC9YKpAJ4Oqbc6pM48+Bq7WG6FinazzX3W2jIqHtz
uL7t+uLF1nYnXA940eGoCHls9OVGWryKrSJnOxkVKSCrLFzK4sfdit9KPzkQWciFle3Umyr12XrF
pTEDPESAX/9K7cX3ui+fsNS+p8i5GWqKt6SYbmrA6RM0WmeDA0Hbe2V3feisRHSsZsFCkFdXLuLU
KiGysLkN3vM/D3nXybzvRf55wTs1+hauN30ReBD/gi5FUaGZj6Bk94rRY25BWBJFaFGbmfpBtgrH
zhbxvsKMPK9kORS7cSF5ub7Pvs5IgMe9rpxZlo6l6YklzXUn8HRNHb8ncf6bmIdlXDP2VW/VBvnk
2Dm01GvT7uHAIXxnhLecYT5Qw+wf9zRHH4HxX2hNUppdkfb9vjDnxWG7lM0sG+f7VRetVGbyLdLj
XR7x6ffzgXqYiLS4UnpKunEq+nJEuNTP9Qh9vZnvmjKRfUPJ4a5zBvuZhWCoIBhX2q13jZCnEkrL
g7emLpZfohqhCMJ4g+POKxrLPz/p1k5H9kmuBG1DO6tAz2DEHenEInbuiBESYp334PVXVPvPzHcY
iZR1d+at9+WIDO2Zz9HlUPkxSeIcpc5MBjTJ6xdXGuanDYhOW+gCc71nuRqBNvdvoh9ux7siLQwZ
y74gkHYrWEzGP5bQjzAlYlqAH7MXbciVvo9FU/ArTfZ77MW8OvlVvdrStTksoeKIUiXmuTwl6aSl
swICNYSGskEZVKksy2jUo3V//1n/SeB9537f8IiPM4uRHMMYjg2HoN2w1LwiffjtoBQouZftGtcH
7ehzy7ptac3xsKZUONKuhIYvAxMHcpN2wOzwGSnjj5v2JMWeh39Kiq/8cRoyFT2hNFT/IcTBhA1G
aUVgaT2S9fjQjl9ePPPyIKzznxLylYlWNjgPjrtQiAxAmPUVHl0himVt3yUZcSebgsxhObUqhWLQ
kpFWpxHdo94SnJ2eLPO2vL4eZGYVUNxlVUUpHHQnYwEAS4w4ggCedW3Vk9So0lIPQWGc50SbNql3
jW1MoF05EHSkPJHIhOynq7kwi8F7YbNBtQChYMxkVyMgHnC0NwRnS4RnmOknL3bWW8FhwcVNiyVw
cQXc1OKWTtBfVlb0VhU2UArMkp/HfyQynmEEufS1DonBi+hXUxEH5ILUF9jDH1VZ4sR0FUCk1UjG
72gwPUHF9lQoLy+3s6GRZhd/e8J5yruriOK/hfuEsSZ6taU0PZ9dcrS7okTt3XsWMy0WtHov8fq3
zVnfzMmuS17++UllwIKNMWhDIRqE4oBuXO0euQxKExLTGeNHk5j5df1E0JxSR8PWeFEda8xHnnUg
fHiJg/eCWBvJYpaaCsoAYXc3lpFjjSRCYbtatbD0Vr0DDTkNwGnNG82WtIkqcrWk1HvLo/hfhKPY
3BMgdxoSSLF59j9LQiqzeWxx6JEXGG2a8gEWAblLlohfCe8QYRe/R6bqEbFRMrssx4ePbW/m9stn
Ov2PU1fdNjFkzjRhDDBEkKE0azrh6TyrLiVF6pHgNC6VupsG/UYhm15gPK4R92smbniBcPSS1Cvq
5o6cOJ5S96R8BrLG3NhbWCGzLoGFBddlpdpw27uVYYhWs/sJnR3cdKxo1FWhlNPI2Ymo7ow0A01H
/HWG/sLIvRyq+OEvV81waowAnr3uxdSnDnUX8y2f/tvltH8LvMugsDLuXevtHh8hVdAgu46oJiWm
gXA1chZ81nECWqNnzLwrEOiuxk/FM6DQhXB3lD6zG7ayWWEFqjSrwW8dfqHBlEMhoVfDTo8pAfyQ
uNVP7im2f6JySTEGJES+QUyc4K5vM/NM7P/6vO3ztPslg07Sxx6CSadX8t+BkxAwYXwdm6wXD6wr
C9+MDXDcSNLnna7YPlk1JgydPisyepxHNY+lB0tN3bwFsUzwW5YCIa4XwobyjFOyXBBsnK2RH1Ek
KEku4g64xi/RFkA4KyVN0+KcBonxyz3obxJ+5EhKU4M4rTsWYEqObkQeq+vGZrUfr3K3tajyrRLc
8dJd2C7rBBJTxZ5aH22AcPDXXbroS1ERS4YtEbH7882ucEOjSjhAKq57ovQUvLY2WNk0tWP83Nvj
txeksjox0/yw5yuOOPUjxnqOVAQrVp70oqX4D005MP3zR3t8xw4Q0LMQfzauDS/jCFh1Qche5tLj
LNAwazv+kr4Fd6MdPZfHKm5NzgO1MUeMK4cJGXHWyOSSK2eWvDoMIUxHotPTebYfGWBY9qysADOb
mxwYivnz1yalsONs3VHoPQWPMoAldS0fuKbtoAJeHFm9c13/BVCiW8wkD1twh5nXWFmNlBgxRiQq
fQXgRAMiJxNjSLvcHzYPYddUQ3T+xbk9fiAgJ75N0pHhEniOPShMf2CGp+U4uLGGjrBaefafWnK0
IJywIvSOK+1di99uil+hChEHdM0q5mC6XIVtkP/96/Rs/ooaOxY8YWX9EyccDkcvwUBL69bZsmIG
tfSt1ZPj/S6M/h8lufw0NAptldl2fJ/fRr3PeBKEGay58axQ4c4D9B0/dmOqfTcjZtH2gA0nWyQI
GU0mk5nL2a5G0D+kpn+PGbRKs+YXecprbNKQFBf0BuMNlLuFvEApZwDPvRoicB+l3nAdMJn409q/
nsJ3DK25MFSa1BTjOJ91u2AvPq7sZBU0dIQYhvPMdso6QbsmOGjmPxg1BdobQ/iT4nPMBQrRzua1
2ru4Jx9CWMTVXxBLAL5qViPFU0s1yccJxypfIXLCO1oYjoSR1Rebt0Y/Pj3bV90q3VjRx0NaX45p
2alwFr3W0o1QTGsF/gJ5cxlQbR1AP2cuPNwJ6vfGH4aWc8Afs79oTZFcHfIXAg1H+Un1u+dzmzyA
8Ye1sQG3WvJ/clU75lYYCNT547tusLzB01sCUhJNg9nk+pZ0koe1tYTvHpj3rLU+ykQ3bpyitoci
z9kKAF3FBhs6W6FqXKLlx6CsBgiv/XXfYxLYVEiJ0er5ivLc5PPooh4iJhAWFnv+mLZ1xvYWMwpI
Vd27H9LybOrHfIauB6dS/GLgRgWOTed2Ui9ZU5XvgbMbsDSfcrZCRBSAdDuhw2mPZ2tH5r9oNRP8
godfnxIIwnMApiTZpSya8hQyPRE+fPlvpPJut8aN+bSYSSR8dbiDM1+pk9lTXgIu1hA0ake0Eo7f
qP1TeTlmvnZT0jtlrA3QNN8nUVcbh9ZDVKoAgLoL6EgnJ+P8tTnjSSWSYcSfbf8mc0nm2CK0Xv6z
H/3F+kk1VwDeTQofo8NMv/D1fnAkMcI1V2MkRe/s9cB4XfwDihNiljMmuKD0r0IbrsMl9iD1Jguk
2P0lmg5T7n3QexFrz1EiFExzxMtpo5QyRha9SnDTGQsBd//e1Bcv8Vhzo6rdkjWLN3tcg0cfxlrb
5QwkVGGWok60GBuWMLl0xMK1YlvBjnz8RrBEJKEY7YFAo0Nn9mTaFOEUplVoE4uRsn0hS1usWcdq
Ylq6sLJ8PBCT2gDP7QrxMYiQGvsLYGM+GrDFgjzVf2i6wdUjnnly4bca708oB4sc1C/zEqJhreY3
3Wp3vsyCU7lBe1bpma5P7XGgEaCokt4F165RACKiAugCmzA/j6J3Rjorw9YYmeME1/POI0sSKkjs
PYBzCz9dVtolTJVc26fjUbT+N7hvUC/VBdnyHKVIC+s4TzUjpKpf5BY8YEEy4ddvxOOQglHc3siD
6DCMjBdKJOX0gkHb/wJtANjT2NyA4eF+0v72yKuiXiNzrodQ/O4RN/fF+w5nTdCZinhthSSAcfRJ
iPHGqkQJjz6IHr1KoYtnJ622Xs888A6qicf+NQHemT/IgPWbBggHgiFgjVLhgwAUWbMLBcawlqJH
Nvi+gqRZ4lIhpdWZXrIQ7lJN4BFGXVdEQ6KAEPJ/lOyHHlVglnGC+GAu3ZWz9l/67Ob1q5ZBac8t
r7G34T5x/Zh1/2LgdhZ+uzStyXWGMfTlp+t2ELFScj2GyG1La5azlRY90NWY5Td+X8EBkJZAhqx7
gT5PbpFqpTBa+XTNqL89OfnQTXkVOgzchucZJCD2nu3MgPGdWdmlZntzYLs72L1miwLOdRHideEr
zUusQ3TVG69OQu9e0YEu+Rod/ZXtHnkLn9ovF4sAmnG75xP2DxKWfXe1SmegQtgxYsBZJmqEGWAv
ysoHWnRkQju13ZHCAvQVYilEfXO2gv9PeNzOrJprCeJ5B1v+JxFYhLvocb9psZyrWxOVGr2hKLPo
5U291e6RBMI7RZx8aByREyTtF7ZE6x0t0QcZpl0asLgYBDL17Y1yIuDlc8pvHiSUewkbki34pKJk
SOs2nJ+xsCO8DVUip5CPCNbullNWxjpafF2CYTljz2hkwvA2g7cDs3xM/FzDpcU0sXjOj2bSjZ9c
HpDXGG2IRITcUSZvseEIoCRciCD5m1SNgNIsX8RPMGzuhjnDgPVcGLB7oGWIHEqJkD9s03AnWorc
3mLtbpRRG08MDkWOPylHsyHHUeSIQBFneJ0X14K22q5IDRWjfsrvAtF9xfoEGTydEAqCsjtN371D
bJcpLPp/bJZ9q6FtQbZq4Bb63r65pHo+luN5QiZUZat3v7WezZzAbM5AeNnhN3dEs0SJZPy09wLK
3qkeTB1ypvr5Y47HKwp84DJVJRfpnt9XJwLEdUZO66h8sHxz0RWZLkoSFxntAKglDL6Tr0y1nD+m
aIvY5O6mAncZST3f1nnlbzWdItR5gZyz+ungg7SWX8kLmRhO1nDbH4zmPRm3BKPu/DxSfVE4BVeL
Mv7YiaNT8mBhy6dIrGvgC3HWveMmLb40r1RqjMXMRLQ8MqaVBmQPAlU14CXu4xDRln4wwK7odJ5J
7+nIUmzbzFbS36/MiZQ8yeCP081Xt5ElN4pg+Hm5HaV9zITOiRU+t6JRxRKLdL8x53+cMLxe1OOa
QPMjUivZ0+RGQ1ZLWTfdETOf6siAQu+g435+2I3Rv4v0cICm3Gy6DhusvA4fHAvohvfj6rulynqf
MAxKwAumm13XgnDAnwgq/rOpQ2Gx1lVPNu+Cw7r7wicQb6j1F+NgmEh3u2nF/2QifR9ZQs2pysn+
RDhMClK83Lrf4+hn85UBe38XZGkrJamQ3NuZItVqcgTp0Vh3RacSHnEh8zuOFsnLMVYftN86clXo
Hu9yb2ttY8z9P+undJ6oTMARNIeLK/9m8/gIpiLXjg0XxM9EI4MZqUOZw9at/lYq+3ndP59/W6wG
ALyCu0iNCEUiMtFCh2cEIhkm/ZoGAWuhE/xeEIcNhqXzQYdX/YK++n1AdoAHvTpYLbqan1E2g0cZ
X2mO/dc+WXFzlhL+tjb+ocD9DxGa7hos9UdZa07Q8fyyQXTFSZucV1jnB7QM6x047FHeQzLLxwJa
dqRj4AJx+OCZbFtuONBa3L9HGkh17jtVd5kG7apvzgl8uYzS0s1KeehHbojakx2g+ye5iplOVJkg
t529sPkU0YXl6BoC/ZKi2R6kaEbHArPuHKcPKKfF3ftnz4d3WqdNzatbO6q5hoVF+cW4sTJZ82D1
vLAvaueU0mq9b5VZQ97GNoRzEXEeqOtCLOxw4bSGUDf+rFeEnUoUm2AIzzXsQIMHt8Qq3amVw1cS
e3ldk2rtiFeigpzuiLHRHeG/QWAaU+kLWge0Hgt4TNtz22mEIwkv9mqfLCAsa9FgS8KvdyDiLGNQ
3tMrab3fvO7QbdlO1bVBrMDxgxPTItXkp1U+geVxePZGRrtsNsTTrNtkWer0YBiZUqD1aaHvOqiT
U4NZWpZxT6jWjJbg1Fh/0fdJnZnnK1O/c/YjsJ+Ic/MH7PmbjNZABdshv/rIdAvBZ2pt7JVrmPiE
FThytUtOUUN2rHN5m+ccjqDHJUFt67ax7E7934n3mg96/UlEdNL6jdH70ZZjXH+HWBNw+4ax8Lbs
WEQLPHjS+3Ev0THQMJCE/tJcttwCRw0zTQFmaW2eamKeVy+/5HjY37Koda7dJAamMk0w02+tgrRp
g6rAlagq8/a9tKgZnCTmmlGeN6pferb9Ov5YISn6FE3Pe8UXmKo6nhCqCeHFRtGUQ0U+6xdrzeh6
ynbhVOweRoV5dZ4HugBTutvED4nD+9yf0E/bcMmcLA/d1BPnCJWk8EUQbKPX/uZPRiKv4zGZUl56
Jzi/2OXq9C+9tzN6j8OgIUq1LAO1+idfnFoJNkrBzFycd+b1dkNszEifEvtK5G8Mbs8LhWpHq/Tn
XPp7E6m0TpYPsXazmjGCWWg82CC34CcAavuqMn6MytbWphtK0ywEDyHWofbkDVyYhOzK9rXlt4AM
QNt6vYrxdXNUNAcgwXUCMbRWVEGmSgZYbqbVMtHxGIVwsSsL0sX8Dx1no4mFovHZnYo97zWUp19s
1g34qewf5aM0nYRbzbYgfJ5qggtc4F71A5BuvNwvWI6klgEgXwsREy+PuOBf+2ARWyo/uKFoERgP
a/tGuSx40A0r0miR34InHgPzcMKnUjqJ9qcOoHnl77r8swC8PjmQec0IUjUJSgfemm0B86AaiW5U
sOUhP/me9N+HG5lcmWWQqvxKxmvY0pTb7HhqIfP8e+HttN+5nwrIWuXgQAUxqS0mqw8jyILPppRR
abVKnD1vVsnhLpSfQ/zVSGlNrfpnQUFTa1OJbx+6ObIKTx7053tlXK2vWo6WsQOMdNO1yNta0Oad
MDNdSX4nEML2oYao6EXJeYounc3EYooNOb8/nMInuo0pOimDiYnkz4/qsgdM5+1dy+hjRSkJXruR
aQABIblU63/x6VO4l5W+iqVWX9DbAmaXnsj9zRl3W1wk22GImlJeHA60hBMBfe/+2JE0JvwjzPEZ
o31MCwUV64bl5rhBPV9LG9ePvDbU1VGn9Mgmr4jKEWVSUBvkb4NpgbTdjDko9Apy8BccPhzCyqbw
WDmBspQaSs6356L+Hqsm/NRI5Qd+zLroSxMagFHb4YtNiLwjbQJKs3NMuJVjIpSWniVsNexEgrfr
gTno1a8t2QpEW5p+UOX90hu87qXdc4M6Pf+V/fX3tJN985nixSvYoQxGh4p4t+WtDhCc3mBpcqK4
ynzxgWUcAbs/MQEeA3yykPWl8CLmo0IleX2BAz7UfzH659VbUpteVjYgZYmHrOlk7/JJs2nwwmER
bB+Lja4IqT2KqdBKobEJFAai+POW2LOan78P3J7bgWrn9DNArXQ47I7B17OXVXRpbtETev6PYscI
MvrxHoVcm4WlMzjGK1RVYaiKDL9JaXZOBvwga16vzxKWJQAUsQK5DW4+wG6Rn8XLtrfs+iW9B+gm
A18fSeHSU5l1UUyQyJv4132tpJFiACiW5gxNEAxW99WXUEPehxH2YRqdugg8igTbwX2ttAGPYawu
QEqrBygTTdM1EqFKRQ+pE8Ve+jZIZ8+wPeolbeJvCG+AoaxAzXnAZSuWt5LodVab38mC98qmd3Ua
19qQvLC4dpjJWA11AcaGpimWwyDHlPoGZH0OrYW/BI9PFGg8/pSxUsKOgErRfl5R5F1EqV17NyAy
w1WrcVvKt+gCqwJvyAhdSpdWg1L/1iDicXpzZeo9eLmMGWOjYMbPgx9EWzx+uVlz2t96gNpEk6XH
5+yG2GkToq6PQrrPSFMUa5PJ+666Mrot7IxpFFsl40LdHijikk4DZStiW2Sa1SUpyKyGPMi0o6Qr
DkrietfecbrXP4M7/13WMsEC7tXvvpKylz4wuFoAf1+raO/pseu1F4mU6NebQiTxSLq47n/weNzg
Vye/QYRg4WuqRmwNgJs2Es1160E/gKa5gFLar59FYwrkzsYQJJ6rSg+sutx0KQFmTianakgrQs/q
XZ4DGvdWlD4g7ESVtSBr4VELlVx4AbWvNDkg5ASIIeHj8qMDnpW6vQYWWVxIyb6QuRVGg0dYlAoL
JgUmSK7mC1UAacsDhLZIiCAADfmXVCD+UA2PSeAZxmDWakEJOd5zWzOMxcgdY/PbVgNOeIIgyUqg
NlPpmKSUDiu56A+ji2GYNkhc5vnnRhaABXfAx49NFueZgJ7so1jNSZY1aVtIOCqRVxzBggSPv/Sa
7KGlBzzonX5+BayJlg2yQ34zfGDTe9dvYkdyaBq++62pKLF9x/mSXw2N3sjy4LeXT8alTn6/+ko/
C+WKEYN8cMFhADN8Ku/ZXCroLcrFrkpNuzVeNHM0sNjez7ffr72emekbxjbJzwyXxv26YTavRMJ+
3WP3ERsTDNRlbprIe+Ob8mhwZ50cpbA7Bc0mQnFcdFGMOkV6Uhfb5izcttK3dc3KVg3BBjf6XWbG
3psygJzzExiDFEWIa+A77+pWTrGeF7j5TP5nkuPkgMtNug3bd84wZqJhZMXts4vnb6cS1x/AzzID
cAP5ggPPZt7jUJ2CwNk6LA5OmUoRmG92IWFbPbFkeXkjdTm5ju83yOWtsa/KqYntfXmW+CIC8AtI
XcquVXOH/Ci/7Z0SUFof44jECS0Q5EkogUW/wLGaujKVCxeD7aaw8Ulpwu6GWCBNuElvg/ZXlFbV
EvebMipY1/COBRU0Wav0G6M=
`pragma protect end_protected

// 
