`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24096)
`pragma protect data_block
giGA109OWTgnmloyaK8oOFehFym+J0nzNKpNUFWadvEVWaUh0BW4J360T6wMibZ9gIbukwiTum6R
ac4q7RgtfuAxI5a4YpB+OIQ0xGwqGM9FNou1NWDRwhLYRrMx/Ru0mq2FTRbD1dkAyQFfwJSRuMrO
dG3tuuVKe1VmFXum7lJr1WNANxcqdfUMp9DwfKYxPZ7lkEhkLLUorY96jkPJhV1ftBcPmn+jv6Tx
dpljfEYaXoZ5TL4/MOhqtCOEbyfgIIxjboQ1A+kt5yZ7J1HdrTbFF8AYaxpzS66SX1+pPbFPSFlh
U7lVzmv+TYiCll+ZqugOj7/evws5KKc0siF/fMfU0oSe6oisj2BccYq/0luj/jAysmBq2zg2HrST
zCW9JvdeA/HkYUQv7Fsy/10MBprXi/ImmkDpSKkn8r5uuzeHy7QbdxzlIhnui0Fe05ELGHmkdSOi
quytY70YR8J+QMydirNC+4iENw3szXQmnfaTbRD+xRA2SVJoLt3QUEN5fiSDzbeb7q42Cnbo87cx
onqqNgEV0drT9bE/VzWprW23JsDrmHurC7zboGYGlkJYVhD0XbMf3xXb5/RUrex0QG4GIWaUuChM
p+e+TPOFa452zR6XlkDsYkiDh7B7R/UOuxxFZyrM3F09TIb6DyggnOsKf9DzMrJE8iPHJkh/gTYN
NXpjou6kES217vVCLzKmsno0TGqo9Hh3IOADCLc7p8fgaD4rllJiZOr9Fpjlqi85vwAu9MZnAw10
9dlTR2uZ4fkQwFv+Tg4ze9E3MVPkA6VccXh3X2dncDxxTu3SpfD0xzWo9S35q3BHt4fVdoP4vJz+
dOzXXUULSp3i5FvnmFyrv1pf4Gt74GDiFz5YY7A4aS12QDM/BR91B5y69qhCQZiR7FayvrGsb+8l
MoQz2gzHNMMon80IsdfwrS67ZPu0t8t48Op25Bo1F+zx2B6UMCa6Rhph5NiVpduJsl2gmr7vut5K
q55rFv1UJ+bYVbj3f8nr8PYY4LXbqf6mgl7lTSc8kuuTRFilvcW+93hlqj2cnCoiklqc14w8M6m9
RuuQsc1gAxP7lCo9hfePgUMaXK/neKc+NNRPapz9SkhLzt8zmw1n6/ODe3TkLYzIfKJkd/l7rerU
L48Uhs0OU3UBvR3PiSv7FvD5+E7JM6tjtNH+6kWvjSSX81ukGuYAZWXM4oq0y0pcYjVPCKZnFxux
uyrNMWO486yxn84SFYC6Vcqq3FKIBWYbYef3mskSvAhl6LQSfApNKp7ODsb7cZci9Pt2hDE5ZmiW
Uy1CpVqX73DEQrTrQOeB+jcpi8N4iRiUydmyhl8bS6yhLknUpKaipsZgCMAKNkb4LnDRYUTEu2UT
B2AfAj1TOMyVDgg4xFIHat0DLD2RPjS30vo9rLwuqyV3za5zZIgX8cU9RR2+TdG6cCw7w3heihMI
OrzDnV168fohtG2FN+4TvGPKl0pN7QAZ/ycWsUae/hmKPoQ6XAdW36JTQjCKzFyBD08V/EzkMGCp
dhsrNn1zbr/DXNeGCUcxrsuTO4Q3j2JCcgNvgnT9jOanUWMx32N+soj+qw9OZWUXWKioAHO+881B
z2XGRT+MESiWPAs7oZO3PNv1ykfGhga+ChPI4jt93qB13oKdjT+Y13kWSfHrtfhIxMgkEA2Xrie0
Mx3JvhLpY2xIfBTvoZypQDPl4O6mm/Us6nfPkIwf4EqXyrbjlSAL0vofpVgwqF3pXjfxZamwKyd1
yn+HAJ7BwZPMpGDUENRV3xH+e0qnUmg5ESaqWqKiG9WY5yGs+M2z8Mc/iV2+da11sf3b0ffl/q8p
kFky59LmoCtXgu+3T1eAGrG2qMpFgCg8R0tqQ9nLEGcNGTLmo5XRnjyUdCSsruNuvSXv0mGX32Dg
830CmhWe+0NIgCa+Fm3pIoTHwVOFnpEOZOViuFIXc83PQWduzTnqqoJINuvDL8xxZHfhbLQAndKI
WGi/LdnmcxNZFwgTJDXLT5GJlpCtHeRYDMx664R1O5oRyc5+DuxfdDridj+hMHSAB5QdX8vY5qe5
a+5hh1CdMpUaqXc+d9tZezfKyNAU2K6sMuCkpljDLbHDaAL0kd10bmQDuxv08j48y6iQPBHu7HQz
SKpi39/UUabRJCms7jAAYcEx5Z02pEpXjy6yEmmjMLHR1M9Od31HXCsgdiVkfaDKYjQ6MMB3wC1Y
01pnv3F2gHNoIHmymakwNyR2vT78wYXXsetld0wuD0YP0gy2Ia+2Vy9DXDmIvU1fIHNmVaRPB9me
vmfInudtjiGxISflFtOLRGJS6Pb2lkPzkRkB8ozycET0DJYccm+7Qza2k6WaT9opRdPAMis3Ft0q
EdhhuPBiK+AIdZ+Z1iW8RALlWTs9AJ9/lj9djneYbdsstauKuVwJlBuN6IBOtoRmhBO+aZMjbf8Z
o5httc298fCVT7yUA0Nq55XWcnVeZSmrdpvS+HzC7A9Sk3N/yYq/W3S9Dkx48hhNftBQa+scHMFl
ANM7o/JRXExuBlwjreErWN4PSUmMPytv1ICdde9Ul3huG/hA6yprTm7Ka6kDHGn9uCQE72p0fBc5
JjPQAGzDbbcg8OMJIjhUYENK9bnPqYSdwZklLLypv06ijI93twb44BozrwUa1nNFJnKX4MelDa/4
z/VmULyYY6UCX0/hoaiFXFrlVxkvoxW784HEw2HzPGUYBzC9Vmlgl2pbrU72t1SgO18rZBz1fuID
vrsx2IQBbfQfIiyV96HvBiWz95oK3GwzHvKJOr2s/yCtgaShI8Jd6UPDl5QBkAxdXyaubqwEnhtp
9WTGb6JIDFkigvmD4nKu/5RqKV16e/2LhrBWoaculGFohjf/EhkBzRUWDVPmuudCSXbLzdbwNvqE
z5h1XkyNsUynrNJqGV8IHFWuXCOPd80OIcXsV/iwTRxg/0C5A01xy4EpNyarJTbVi6whsIROzHgB
Cjn62XeIS3B3ZdM6WsV6JQvX5pM74BdKlOK49fN1PRJI750Y8RuGQ7t5GGYWw0fXPriW/T9ZHZ0J
LrTylTMpcjcDLqkxzW4grsLl1gVi09IHTam8x+WG+L+jrrVDMnp5ifns/8YzDqnxCNxIYyuEe+Dy
0VzuGm8tYXBLdYvM0fNtVe+hfv53ym4DtGm48IQdfxg9IYit2aLUaaIMgiI2z1AlKD3NTHfInE1g
+TKkbitDNZddPwoCG0dZQq8Co89YcnJOIAsgM+h5oH7cPuggr6N5aZ7pLpY5gQzyrq5zoeiJZc/4
l+Ht/Uu2bbDXP/j0Q3wQaTTL1ysr5AnqOzV3wf4nm+AI5BX+tw0F8IOg7SJe68ptA0r7s3LErDH3
+3iuebS/4IjRVamONsHJaZB4wbVl902Mp8K5EiKC/PbDVvDLHNNFk/kHLtxDZ2WDKPLKUBBDWiYB
urriNZXdI1xA44il4CE02JQRJKF77v207TPlvLmIU6LENwx2UfqXB4xR06O5QGDh4qrZIodex5Wh
0UNKtiwtilUkTS/kfUDFDIeC719DmutFqR7ymQAVboTQ2VQvl/tpFnHjr5JeDJuNfk4J+RWpSBGA
yb+zlxUzHoR6fM3uQNfIJeVhCuzn0bQLCM8erPtEVwlhpv2z4/XBkewB8gvARgNF1m7mRPLoO45h
anScE9ibIwV2FWMRAmXETLQ/diMFTrQeXOaFFHu7aMMxmIWmxhYlF07Y+M+rVm3g4q57RuygZXS9
w0kS67cipzNGnzFe8YcAg/MRAi6m0sQUr1riOd3v7itULSwlnORq5UzBq4M9NzQvqyTjZcWUX73/
wOn2UuVmLVhXEJ+O3G/TPnkvcwuHu5VO2zdiRxhFJj8/eRVs2JdPBnPEJKN585/tiyrWTmavT2j+
x5jxlGJMlSz31eKl2GnA8uDcApi30e/bbg+CzKogwiF9Fm5Va7+uqP6DP+8O++XOSniJb0F18EXU
u4x6wey/U5svH4oac15jdczglXc2QTSAz88blq7xrP1bzj8BTod5rdPcoAyXNcPN70GRO77AD1aR
8tV+++aWcYCsvY5H2c5N7+pYKcEF1uCBjh2lzlRZSeD4/x+cnLJMZdjUGfHe0hsKh2MhTgXWgd7e
axX5M57fFr4UrCzKqy0hltar6d5C/GLqwJwRg9Uyepr8z6p/96ULZOaodFz5vZPDYZmFRRPG6tKP
IMI0maPCG5od3MKTbUhwfy6lwJ7k3sm6lj0wLp75m1Yz3uAQgQJlwmVMBDplHMnw/XZGM4y2Q9LH
8rdp6Ozwr+F8rTiJL5JhUPoG2dBbDm94auZXUidrw1DnLIvhnmMNBP65lZ57+F8vtev+MFJv/R48
sSWpFTcLmTCKeo99s97TL1R3DU+96xnSQUcaK6xaKzUaFT36OP1W7OcgePOpU9eaH4iWdyoODVgv
c3JDpPdMvRwJXWth1VVE9joQ1yDo0RCe8b7QLAdBKu3f69DtVEmLJO3mqwkZ1mng/Jri+nLmbXqS
gBqaaxlNY2bwDZB7+nnwNRM+AHjKLXdWhlcgFLCp7EMd96Qsl992R82VKnu9d8/4Ev6RTjOxU99j
u5F63Og82UjmzavgAqqMhaaWCQdIcrdv55Y+zx/5Wp1Zh22qDeFuxxg8DYYFw10Ap33GIgnQ/waa
RXH86R+CIw1sZzMKS1r22Zt153ZvlnIBVT7dVG7KAd+8IqwLPr3QP+VEOgJTA4P6yWdvqes9GpWd
uCZqihz170oQvUJHuPGDjzlwQgKRFSX77P72hkZDf4oPSmiijzxGMyAHyc1Hg5rKtH/yZmmr7wVJ
zlgdOPXDIPJa6HObaem5tvBB3rvjNXq8odnFdojmA8KCAjsnQRadaBk6IT2sRXS5FS3IETH47xH+
wqfUU2EZp+hjk7Iqe0HjaNDGEYxfl0LNBQuhml0UbnuyWDExTb25susU60cM54zjQzBdTrjUR3Cq
6ZV5i0bIUT+yeLfChM74R+U+HlEa5RNGQAoa3Vol5wPF1tuzMjo4QBtPxMr3gYyahDcOlI5NwjTU
rUO3LDJQeas46KYXwgk7XbZ6sMd+1XPc3zL00oXqOpwu3G+1oRdiJtKls4wNdDZgK/63RTDt3Hnt
KY1rikxRZjxjkVhkkNR82PNCm4X7ytx2A5R1EXSd+QlOTqMlU482OQmSOXVb/GKNhxLQuVwl8y/V
uCyEIKqRhJsBn9J3HuY2LGlu+dU7/+XLrdrg5sgM/f90TONzYqklcsO6wFOkAk8LtbbNuA221WQj
TZYyZrMpWQmXYeWxbhoaJmk5kn/7pUu2WfSJjUeoshGEz8TMuI46UKyhZ6BsK1vNnIt7bnyLDRB0
Arx/e6R7ks3RSOAHuUkyGMtViJVHJDmPepdwPgJG+BjGy0JblIvPQNn/O08s/iNWDLpokVQ4id/K
db0xOsgxcu3Rnsbh3Swd2V4u4NwgqjmasLUArEJdY91NgcLNcUIEF/+fb8vQwdlSII9/L3SVC9Ee
0GYwmJjSHZgaPPc9GxndF/eNC/alH9up+qyX+Bflftfi9WitJSO0IBmlKkCvhhyOTJ1qrip4xXTQ
kD6ihbXa2icY9n55PN1yoCsdaU76gxkwTE7eT/Kny2WX8goFXO2Po1ZNn7KFOfCSV5bYvLJ7AP72
IXZCdz7jKSgN+0jFwNxbP/Yqt3MMaPeCjBs1QC4nAwRphVacCyz2bc8FUS4NF2MbNwHCTWzpeVOF
IQstDrEF85rL9XxdGb/31bJ0Y7p3KKuuEs2ZPW/gxCv3bx1MFXpfye6racqqP9f5fwXbpuAMbXHb
NL06Cyu7s+drmljpoWvLkhdGhD25qmjUnD9YwWSUnr6yLOreVCSpjBEBhbOKT2ejboqnnSMvHvZn
3OkmtaC39e2xtB/YO3X4KEXPaXvpfEX5wLxQlMBljc34AFr+bCvCtXkvf+Cj2Ck53dDlHVS2MrqE
GaCwND5r7HjJ0cDWYxga7IWVvJ1QlVZIMum6Kjw+TZi1e4OdCeyr+zQFtsosgZbuo2HPv0BN2J9T
Jar4dJ22QzL1JkBqgIarC6DmQyMvPxjkcmiBY95qx+iT6QIXESdFvCvP/EDcHKO01HmQdEjWsWQk
4Tbc71wQYKzCOvKRQf0cWbRMoehgbzpy0DmS/XUx5WHS6kdapVSBg8JdaD3oWpD4ZNgBS7UZ/tgK
BNmlJ/AEDptf6X3Q3WtjZkFukYoNiWtF6pkUTfIJsVrtaNJZcU8QvEhgn0zvTmMjP/V6QWZM9Vdq
JT7Vow/b5hmzNbIDNr8uyfmaHxyzgYYrLJTe7be8ea9htT1hsGX2Qnx3NpPO1WCmjGptC613+HLF
qBCEQRbI3+hkpH6PSkzgIaLDfkJZkr2H2vSRzfKBHIbgOQXTSvjieUqa1RWd/6y1B0SJzycIu4qi
SIieRXwokJwxxqbvdyCpBbcPKuU3jXvlpqn1aKCc17VK91eFnu+PhMkatCO34FatiOj+w2Fgc/Ye
6j9Ua0jmyXPIs9gQ/FQg+uGutVyAGYJJhx+kjbrnWsQFMhGpstFSfiPeH0wdUaLEVaYjcjhCNP+r
749Uay6s0TG7cFp6f1wospNSoixcGZtzbRexw6dA2I4veLrpuksIdhRMtBkWXDLwQ5ZQSQZu1xeN
HO5uyekL2R2+eVhWI+NiRspOS4dWNskyw/had9ZTe8C9r0Q2AQfrkh/lxgsR7YiFyDYMIYrJXX7G
R1LPn03QMvhWWZr/GZ8z50owVuz5dVyXcCaqpusj99nZzq5k0zuh7xYKymQVWaRsr9ifrkBd9qvu
OV1dwkffOa5AWfaeiTznCyuvzSPM64CmcdonlQMBHRP4fNhKeNAa2n/SSpgA6WoNDYJiLMBzG7Na
Z/6lNpRE9CTbBHz3WrCn4vViTCBLDv3OpMkYNARNCdGSdbAx+8a/Xecso7teE3ps6b6vabxPxPqi
bKLipZ9YWKVHYDpTMmaf8P5FnYGYAwuSBy2KXGH+OhUjCWfnz9DNQ7OV9SGFeTX2/OPRUhIkGNzN
I13XvsAANgSF7RZUAf8biypeo025vNbm8SQqWfa269RMgbL2a8ORuQcckEsFVSe0zfvbxCKCq2iq
XgvaB4qdTDm+ejxtItgS21KxfY3PHQ1Xu5ncLiJ08+M89XadBvnHS6uotTwvcvfN43y550ArzcD8
RsB4KOQNxQfrc8Top62xI8Z9iEwvUarwHpE37cA2h2n9ixZhGXSSJWVdVENl62UTC9CidWZzVrdZ
u9WtvHKFV+BLzesx0r0DSUzh9yOLuIarRmXhxd5ZC2ybl8LMlAFuOnTxQrl0RY7nVVUw/SMfSDBJ
pbVYxB7yOP7XnXOPSqVUuCOfoipCLTmV9Vagyrq+HY0eJXd+XG5G52KUHlhtyiemjsT6mT8FiK9L
XR40RkcNGu0+lG0YvXaTLw+UGAmQzJNwROPsnluFwmUv0kzCiUkqViyi6BfNOekT36Ur/WSj7NYG
euoogxbgfdSD+zfTcv4ggHZb1QRLiTsXH1u6UkCylX6q2PU88sNUHzVzzM4flmfg6zGC9D+vhW3Y
gQbapDPrfC4DnwWCuPu16QMe0uBJKB6Q9+N17Z8G/64wtmP5lrKiYk5JPtG9LZEe+1URRW3nL5wE
iArAwy1k0hzGbrliwBdKYXleynjhOKaLzT+YZqZS6Ap02DzdhmeHYdaYcyXDS5TwheMPzDWT6yEX
kLeThg58/eP4g/jQ6KGgyb174E3PdCk7lV0A8TP/PMPzGhOrPAfCP+Yj85hSfMX1wsSD37Sz1iTL
onui0sozAfbHKaUkkDO2JyXICubcvcfnQI81txJJQ+0LPmkyd8JMHJymbfGbTxcPnDE1HAi18pFq
hDUZ9UKMl6JoWhFHVy7luXhOMqEkrqoZkxK8srzBd6HZP97zM7YtkMlRkxu+9i7albIwGvzj7/1Y
f+BpHnYuj/q7wjhc5IwCEKP/S7Rl/qHLoteTAVSXiRS0/Hks9oExUFP/iQot1iWLxo+n1ViUw08w
2tA/KPmNd5Lmo3N2U9ItTysSiSqapxLWg+G3xkDc+CVgH+XDWRDflMnS1mGpGqLADm4aMzUaLvPH
LbwqgsqFhikzBpCmZGBdPDVMi1PT35GldAahP+6hTWu/EkAt+TF/ape1Eg9yCA1l1PyMFfGx5viC
t2/JJmQwgyrmGWGMI9UdpiZ5ycwDRnwky4gfQ150uIrvrKWCvT4WwG7syf1MnbX5/N0BLVDViLEx
5mYj/hh3/Oj/vqUj9BviQWng71SLjCP0Xa60Lm9JhOwcwAO8m3CqKGeLWqf7qMYUoyJtiqwtYyEv
W7VgQKvWCMTtIq9WbwpwjXgARHSJCtRzNZpTPn+BRZGZUzODf9J+UhmJuegjCElxWvcmwYMTSOVu
Y9UA2hMQzeqeZJ/z22iGiGjlgqpHDbuY6sEoC2neax75SLJi2/Wup2qE29g4L7OVZ5XUk5Ir2bNx
eQBwpdZd9OIbt8UPbx3yiKtzeSQryS6U5FGAZDVib04x5cOb20Bh68BOEGRskGgKm+PWDfEhE8dS
lNO2JslprSeTrWIDvmisJ0Ltdr69w1oV8uxzlVJnv0himYE57V+1MzSNPbYZRbLsH1FnW6VM8OTB
dfDoNo0sm1XhqvaDgLiPcCWiXIzL8dmNZrJ6bkXhIH7LwzAfiK/+MZQSrz4vbTOUNbfvlm+oz6rK
g5t93qjNmQdwO0xnnivBmy4JXancLU9Ma8dBt3zOZJNfmr7Tz4dWyxEEWdTM8fk0ekWn3MfH/mi5
7DmKl4sMhq0jUbgnlqU0fH6VkLTtJgvmTlpnnl/XvntaeU71znvhTC3jkLp1+eA+KujolWbK19pS
RZhUTmSLMT+kfz3PKgCoMJY1Q6psGZfV5Y1IDvUkwmils5s3zGTCFMSaX/As098hyQPUaLxFnnsN
xGozWDCkHW/8Lyhvht9iWqs58bGyMJ00j810Io23CiHvk27IJhklgkhurx5dFsIs00PYgqAc9VSi
WKpEm00aFsmZ5w7scNsSyB9Jrj+GMe2HcFbSc35BKc5/iuGO9wiTNBmi++UwXF2S4VdUIYgCl6no
sO8pslEpvOmFE/Qe4r/NbCScuPC7iBZdQ6v8+MuqIpwa61zzY++lM6Dlyw5/H6vrnHJICaDwiEru
RhFTB6r1UGlNfxIcZpi7fWYv6wLKMjeMOChJWva8pRxmoJsR12qJcPAC5wBZHUrOzMFlzQa0hZrU
0AsYZDHcKDHRl4CnOKYdmV7uFq9VGgOSKJGzY/wyqvQclSd7A9tYs4LUOK/NZjPCVuusNiv6i9ff
UzJGRG5vyE1ZwsqtAo86fVY8x88uosjJ+mtxGuVNBfRnQRpnhMEYCAz6i25YVboA2biX7gNUEF9F
DRP3+edVX0ml4lDReELRy+NwW0nRPzbaUWbwQph/L5+VOO6xv5kRYjtfeAmf3EzEWL1H216UyuZ9
nk4X7C1ElxRkepfaVS8mQW8qgVZeuaYoTIatVGPuGMJ74TpccKCEDhuBko6vTSYBCmjYYAvPLtmf
WEPiExdyrz0G3WUhpjO+WfPbi69WKfX7d/5Qss9PT5AIjcVxKIo6m9wlfyhLh6KCE69WgRXPN3dm
SrbEEXnTtKZzm+1mubYW4BY2Yd7kdGA2PAvY14H2IJk2E9ZrDnRwo8lt/cEmyTWoCX9/GMFlRF8p
6DLVr7EjGp1TMCFAEz6zpnjysdBONuBrkVbX7YtdC9lzjtVSOqCnK3I/fv+OEIcoWc5nPUfSi76U
x4p1o+Ehk5R8qMjWjyfkoTDvFTJKQ2MVVElTPwWYIXu5oMRyJv5ddSwlAwqskaxOa0ds/sgRF5jb
F/aqkWkXor+FbsO70cf6MpuV0UkBQ0yLZMWLuaGgTDkP36wgMzf3ht31HCGIyEm2isWAI8dZ8S1L
HJgyH/gT06fpUr2l5wSmVcM+FVj3F4S0babdOtirvWIQChOKbaL9BKZxY4r7WIUOkZYPv3uRFYOi
09ka/M0TOpC3ra9pu9qGsL2EqGbeUqjSMyeolUIZPNnPZEdQRBYy+xsBAShFHAQ2kfoBuneE0Bc6
WM5E5iHisWojrpIz+VfonqprMpJLbgyBbR7RvjAlTVVJUAUNTEOCDoo9zrC2Le7hHjqVoGUOU4w+
959Wt3Eh6t61+my2h17ZeWE79qQK3IgfoU5N7TbJ5/R2ipLiKkkUYCANBcxOmTc0uXLk4HYpimD3
uT1i5U7QuWhrktXNfsMdyjgKU3HkTicZVbFLBASnQOWuiqRpcr0deCQwv+zpldhjhoArOwIxCL9w
MMSdA0MQex1Sn31GUjwaO8ByEZFFUa3gMfNUnqzIUhuPqhgEPfzJgpBSIdqddqX1oMyLOcOlYh6m
2kQfu4nqkph3aFrpE6c+b5UEe38e33xTHQEOfqKwnmTsup0mitZpVLZDR4jkLknOmIZ+hn+xhg0s
1SqiPUeL3bjseHtjTb2L2iLnBsdoAu+HXkl+SWRavztTDbEZZciTyo/rAgYZlnegefitjA2L9zwI
ivqvUWd2gkVz6MaeyxOqv4cldpei9WDX5gqDffDYqHe5SojJ0xV0NUa8mDi9PJ+LP1NuNUHMdT1b
JJT0vxQx1UfmIRfDWJ6snxcTZ4A+F1d6RDutTbT07ULaSKsEzJxhyWRyd7+P9nxxivSLiWfy6nN7
Thw5zzmSJrxIglyJbs2fNGXUAW7rW23JWYWD1PnMwoYpNagfxsMP8oEtVJx56+ugXj3eiYAi+NA+
+VVpCLh9uPwlHHtKX4O80fUk6cS1EKfDAb29wN/IHFLnb+VGMqckaB6dGndVf2zzj1ThlsX9aZ5v
89aQwED39EPck60G8xgAcj1PbyqQSicdWVka+EWim8xO3x3mU579oxey0e1eAfj9YJu7zQr8+t6f
GXydSfx2qi/whiAeHEp8iBMNS9P8zwWTR0wXcFbIcZLLgodjpxcPnhR+3VHx3TgcDkK6JH3Xbqgx
yaklcgU5Qa7ags5X9PEdFNI46JUeIdyXdPgsYi1PxNpQgkyQ06RbKMS5ApQ/PdsvKfB+YXclx+zx
tCV9OG5D1j79I4YL0pmZYbZ3V9EG5g46FM6RLlfBc8AE3g6FzLsqkL2ziwjVR1SIaaRno3P+vAm8
dXLMqQrUGnx/Jur9QgliiHylNfhC4UHvPgDa21F+mFdijf7o27losSmlDaL1cMmMwHdzsa2BPhG2
IQqnEEwTrqyHdAPAge2v+wFhLHDNH7dzZiDXi0/xQfu/UyS+IBMyxLiwxEetiuCxz7Xv4DJSymwg
yIHPy02iRAJ6qX6vuZ3OWWZrveh/QmC9vePY7Gf4m5Cb19Jqnc6x/+DNr3KR56tbUkhXqxpJTSnU
K3aA1qeJkhQRVjv51YWIit0tTpBhu/RK8Ppm+oHqkQ0WlB2XcNIQSk0+rRq8ehap4np4f36POAR6
eYUSfm3Z8KdQgunBsS1AYkwu4v+CSSE5tPCFjT7lY1B+uV20aFMOu38nG/oKXrRWutDdVaOlxc/x
MQX7aaveiurH20aWFay+zrqpI5vx0OYMqVUNfLhPPm9eHSi9bb83B1yF/JEbtO1Zl+ZtMQa11tCJ
tyMV8ZQzpBtMFXB/NLhl1P+OTo0jtS9TXveEntxHk055vuLqBzZV+OTL9QHTowUvhQ5nVkiLI+qb
4VW9LydeRUqKobn+/rr1VAutQrn2TZQcOGIqIMKPzRhmrVBvk73JMUUsu9psCTEkxpFFiYCF54Vr
+jdjCeVmnsFhNme744jnJyFiaW+qcy532+69xeyqx6y9waO6i6h59Rx/oUAxyN0p/9nebZ97uIKC
roHbAP58x8p3kooAHIwouTf2zARwm3ZRYdGsAE0FE0sUPa32alvtoZFQUajICdy3ZhLQcIQ0VwxV
Q/hmz9UP9S3YEc0Ah53NeFHxon7AP4Vd5i/zkRML+R3BfmJl7ioDqAY88iMExd9JIqGhCZ9R+Mnc
zU/710ER+38yJxKHwhFzcbWyys6r06B2p86Oo0hIZz4uFLcnoOY9/GIQiL0MGF8o7cNCkIUbS7UZ
HHaF91SYcHaIze0EqVmd3TyN06b/JeABUpgeTpoLylf6GfMfp2BzqZOhfBdzU43Qr/iTGPWlbCrp
8+bsOBZhpXhTX/gEelwOGz/5Kzld9vcBYMv6O60BfVIVpgMGBRG82snwpRbsAKxPf1OT5bTW76Oa
84vpSHSP94rR1BpBBL5HkPEUqelHe0kJbcKRAwpLcEvWLMxvuhBE+1snpzUlqS7BXzqnUbvl0ySn
eG0yAz89g0wbqdi2CV+b3e9/os36Aquhg+/qFRF7DtG8D6jV3w+a5HV27i3VHia1D6NBHX3wcY3/
pZcIrBzKKcI1NKXBlfR+p7KUA6qq+M81Te/+7qi0vxjSebmcpkj8qSyN/CRFrIJZkb7sGpEv/Aqn
gO5/zGaYQya9puhQlPg2AXtKM1Atj93bmMI6F8/WoyxcXxbx6YdkruvLXEfJObuuEE/6+0v/zoeB
asKBVR3u82CqWI1sOJFRsAwI8rxa8eRBkTqOFQA/YWMjcJLyMj3Vy8J/eR7E/fYDnAtBOOy8RFk9
uB3XyU/dCAAultzixBUk0y/QRGzlFeUk7IEWlU+xhjU7Kcfw2lI9bZxR79QKL5SJZq1bZxRxfjDB
bCaDp7bUs5YlNu0UrGniVCwzua81HXucdkDfQqZjjZf2RNENjT3U4xRIKjU8phhZad2kWsxPvh5p
Te9K2/G/NXeFobB5Uo400o73CJoI+JuiRqe+R6EVJOANII2HPD8gexdKEDvcDve8LITjp/I6Trmo
JJ1I52o6DonT4EwfObV9OiN+VpJ4cRPeUtAfBLV+dRDH+A9e2k/zgjSiG1eNgHD2n0C9Fa0KnDzQ
HJoDfi4+7nG9dyy0NUPp1hUsljgCZmpSbrl0MnQqvYbjQF6CTZtEe0QLilcHQ6w51VW83mDK1dV0
GA/ZOnHw5tRoB43wmmLhQVvtt8cu8BBVnkSYxJCJIQ6/Ga5zpzKp7YFcVOfYNi1BqCT/ZH3hIZbU
xr1kzaq0vJEMwqL/h1+5xDcheWf5tEE+zdwFO0Xx8u/99oaOBECgZH2tU5Poe4DjXmVMhhpIIwf/
N/zvQk72WGEUfqCVtx4LHZjpE4izDfTy5apWxLHhekr900CsyMc+YlpdAyNfxMOHzrO0l4jOp5z0
PNGbxsshA1aDH+6HAFEa4Ko+8xvm0n8Ma5JLIlKsV/0RcHNAmtZpH5+RggnSpzbM8+DG9m0aRwuL
6HfaAlsTADtZc1IW3WXWgYkS4yY/BBy2i9lTAKLPgoJnKsTFux/B/JTzbwKotNZ/7Nxbbi7uAVsT
n4n5RXOgqfFJKe33n+M2qRff+gQ9IepSIhfECAL38yt5vEkWUGP0WEkVsQw3hMmfXFcI08pFp9B8
riVoAlJIz7ZZ6oeatpfrDrDUFKlbU4M2m0sSzpFoS9K251kVh9PI1lZMf2gvnTdJeVlw0/pT6hYs
Zi0v6mJmRk8sl4gZ47zUVRBEjoLIJVg1HQ/xKMUKDzfuJQl4y3/achPrVIh7v1kLaaJ34bZhu2ip
EnQUfeUGYSH9E1njxdjP23uLT5nrHqHNRFS9VooFdmopm6+v1R0zXloDinMXsZalwb6m1Mrchp7e
tphD0JY0KNIl9myXdozMa9QznfqcomtjdJpRqFR1lNq/ZvpM9Xd1bbY1RmRTITsPPcomXia5MiYJ
Zwl8npVioTCv+1DetGcN0lIYnSX0vqIP1bSOtlJR7GKxfrIdfZ0llFQUNg/xxapdH78tka9xzLlh
mmQ7xvUgsZBLPxoaQXrF3T48BMxqIVneUNaTJVoju6zXgiVunbrTd77gEqG0p9NZQNQZTdGpMYHq
/YH0iYQdUx+V+JjOM4NvGBwB5Bg1GGPC6laACm3Do4WAaUcv5/EU5UytTf15cQAfQQHOgBq8vLkN
OB60XZ0ov5s+iJR1+xF9J8ugC+ZvR74CA6itO95M5kQrLp+kvFsQ4QkhKi1ReRH3f6dyFFo7sN4P
kXhz5+KPHRd3inZPIq42CMFFrUJMvLp9Io0zd3xhc65SezJl3UaKnAX21fFx1jD31Kq7ECehzIba
SsebjV354X9IawLKoLNOADS+v0UWkpBfr0Q9dALKtDLYnP+uVKZcjNWPv2q+n2jFPpcJ4JwKuKPL
nJLgPNdwcev9tPg4LT4CxPEWrXwfg3RNMV28YEwLUS6sHA6K5UVYRH9plc83OzWmgMqxvokkG0pz
Z0BNDvrck8LfbbdV3FX2tYCPT4EKFHmrf254MLl8kegckpMU8sAsWZAlPcMNYd8VYPV72DnEKT/l
q/0zeSa3s/RhxW0WsVLwefvafCJnhpICIR0s1dFZBKgZpcIOwu9Idg0nU1eAGERL8sq2XUZiBj6j
P/4AUiOyFVe0JayNBAp7ZbUCl1tKWiTjI3S6kNPIdyBOk+m8xmo04rjFDAnSibYbhE9ZWcTjdkiz
GIFFr8FLGWrLUEF3lxZsnTnI/6E8OeugJpdtymyeihZyDYK7nix2S++RKGpsgVWM4Ah4Jo/EV/Bb
Ug6ioCBKVnXHXevSlYJat8OwvdDQ4ygssZbOiweONs//zzVKO5DQY1Gih5lRN79ij6tQsuql8NXm
mzWMvYJVBkuQmG2R+/rHWKMFKz6k1gocVjRjPxrNGeGPrxg7/sp+NVgs+dqW8x4ylWF/wG6CTOix
gqxNUuraIEmdtCU11skVG+UeX6Bw0BBCC3gXXvI6PeQU8aQ1ioIUdAqJq8wY1dK5anTJP+u5vjOl
9vj9SaORR72W3VSUKZmj+r+UUDCmwGaHyBfoaiExl7hcskycFDAKzcEYGvoo5CVwQ8y4OIXOIEm5
/vURr2aXDhCO206hiKvZ3FQWr9D+eDmK4uumHujiUEWiZTuhp9cXs9fZIRQfayL/pxIS684louF7
FQUy56eYdh5iey5KWXVQ0kelptpP+nyGhP3n//Xubrx5SlJ6jxWdjYWjCWkBMDRKNmox2fz5YzKS
LcgFeOR9p+bHA3YVwx9kvjFkOxgimH3pujqSsV7/MBu/hx6HqbIhIblI/wYCSDz0jDf6eg4AJZDC
QMyPVpzOXzEtHOZo7IaxDeLyApmWZ5qiHJcEwg0J820lOabsnSwXtAfrwSlufvJyqjOlhXBWLVnK
HrOuHKAlj/wotwsEzKfUOZQOnaWjanu5ZUo2mduBOEkIDqgOWRLvTECzlQFbLeVOwx/DtKBZiyxE
WR9JzHIV30UinR0lTjE6xpkaD2kjQs6SmABjjU78TrKwJpLDiWufRqaN8fZMwB19Whq2qqwMe350
ZaLo8hsHdVuxxUAoXXTmin7kIIbRITAGY5QjijD7GPTnkD0E2WA+R11PYp9mCiXwk5gRmHbMTp9u
oxCOFsd8P3O5GdC4d2Z8rQSGXOPaoPyBnBBYfL1tTy7RGoeVCJZhfxb3rbiS+V5N87xakEc53a8t
094sMWLJGJbS9OiZ/60zMtB6W8mOI6SJfIfQKTFqB72ymOQmF8NCAHcbeTIIZH1FPEPvWbuwAH9/
0aw1kuEf9ufVpIj0C941NgeQVKiXuH2PCjgRteiRMz8nCfnwx6Q+iB1uAkjDNKVlgNJAFdz/Su08
SHOdCbynC0IcKO/vbCI29bMH7qZxtrKTV1mIzJpNcLhExi94bYCqDEWGFFgnf8iYxWRpqCT4107w
OKdOUsJw3YFz4w6vbIOZuvI2gIYetqwFTR8xJ/eKC1zdKPzEwn+BpiJDHOeK0Og48AWaJiMlNFUG
CQ5YRULxVEw3sw0mXUUOb7xdzjTACWt+Z1jtv1StADL0bp4fBfcs+soKGj6h2DVGozvrtKig7SrA
QuBW33mpIQpVSCZ9YEiSIgw1vIiMmO9Qdn8AavqLeAFeNyI0GndZUXhGfGQNyxctfgWHPGV9j1oP
y5+NJCql7lday2Ayp2N120B94R8Bt+6RpCcSVzKotxYUFZIQS7NhHNtA3bHYVNWBukqL1GqT9hiG
tjD07QinQcryQXKHO176+ajAVTpU6Ah0SLpZLzeT0Y06ZNkM+kvsuQsI2ciKP3qIETifq00pgNhE
urcNrYEsF1WNN+WlTeoT33+qPxMclAn6vNSqwEYegaBWqB52lwu5dtBza1SuJRDPuIVTm3fbvpZU
dSpDJ5SgfGhtoHn/oZQEYkTDa+N9kx61C0o7oRwa2lylFJ0QMrmSUsLCHByGIYwnw/fBfzMMOz5r
yhZBb2GYcyQx1dSV237Y3N5LyDCQkvhLG4NfYfbEj3LHkZaodveMu5uoYDOAkThUFS5HxMvHKcDG
xxFNh3hgUVSSTqNOeWInVTIUy9kg6dW6R98cZB6HKlmtfMxGm6gJWXJ1kayXZKyDDVkYIi8IrHuT
l3oTOmcuTTj4wYICjGbgh1zgucpvIeE0mOPxuSfTMfvoPEYRUcRNZq2MHU2T23F0TTY0HqckdppG
ztvoq6FCMWBZZkQzj3c4xoyAyGo02m2UdyYPJr52vrt7ErLsMBYYlhz+wIUsI4z9TfWGM7s88w/k
2KV+GpWGM3cdewRV6T0H8SrjfDuGJlGBAhvfqfiRMVKU+/xK3Ow30KbOtbz+6ZbmGh8nOaheWREX
n1cSdrUfywm4GxoUefcYx1+YvgGIOXLVND/8G3+5Bmy3d8aB6J3ZdJlOPKN7cUhrflhNLbG6IL5I
ig0y6yLRgUoER7VvvyL8ReVqtI0AiKyAbSzFkmJJD1HJQ3pJn5mv7MuO5n9PRwqb5LUvr4kgkbNE
TRj2S89oiAd5pajlZyYdJtIf9ADwsrGAAle0XprXaMat/sOW59qv9CPmztUGCPc6AfaoqIFw4wAa
2zPg4//JnOCGBQM+UG1p9wtbjiNvk4zywscJpneRSw4rDY9+QTvDAyHzOhb9mKQgWet3yxXRARdd
FDlGD+dBVyodLPKHD/1BKwHX1r+d3jJPB7rbT2ZwG3K7vCHWnvjNynZiGxXpvdNhVB6JtuyAGt/5
itl7HaR0W9aXKMAnksTU8NZhC/kOLrXEPacsOGvHbqUNtSqGEFVjKZ7mqIFbrk5hbG4AkPS/7E2e
eQn6i/XZqU1mr1fW2H/AQ7+CF75deCm6rqlamuKoG7vB/wfNDvz9WI/Am2m9AioSmUjgbLcA9tNZ
PCDppxk418YBJfzrJxV02HKT6/kCwjqN6nvvpVzb1+MvhyPg/Jc/UbI9q8Or4oNkeSAXVo4MQyCu
tYj5yqsRZ6bJjaG5PTJgVN7sL9DcVXEvYGEIaU0+zAJu+KmN+4pO99A4tWXfAMb7r04UwTVMde/5
xSnl6QfphevpgMXbn30QB1BX10CVnyMC9zbVfh6yzNkDwjF4OxUip+pODDOcTHXjMhPNnGjsWILw
gXK8qE2BzcmKuIhZToMuhW1DYkUI6uDU4eB+pkxtwvW8Geocxxjgs9Am3oWJZs4rLtGSUxXrs6C9
LFlo4VtIHMd+d9nRCvif69C1/l50682qEVMyuKjujX0OGbF3q9zO8KDjquq6IijgXXHdqzdimeFT
J3zYLOW81BRddx2iwVKdEVJNy6lCx124fiIHEklwKdXxzJ2+rPUFM83gpc5MBVAzZXM1ctYyZXRd
8qxapo7SSAG/OMp72A64zPiFR+MLot5jGjM3M4vRnVslksBBRDAHzj4Eyw25EHiN1BVrKPo/+OK6
jEUd720iGUgkLZrgflvdCMWp8qDBu/byrTGbtcj/qBOWu0zzg/h5RIjXp7y2hGE6f6wCzRd8MiDX
x0mE5M2fbEGa23cGoPcwFBDyuv3aMzb7DlZFt578VIz3Q1LKEN1hhGVyYgUi5JslbMzHwopv3PwF
bh40ajlX2ws1r4YXGSJ4FSxU5JZpOpxoKeB27L/fvGHyYkJu6FAitXvTpEZ2qW0d9U0HT9pCWDQQ
uC3xMpnxoUJKfPbwERRUpN6TImhcLSNKPNVKD7roSWBwe8kIZTqxsAAv0XHMSmK/pexzuMZtCr1i
Y7EOujdjXeNhE+cwAMUVw2sJfd2EwQ2gwSYXJsLU/bioSVY2cItU9r9+teZUYpNnHZpdjVjLlUX1
eFeCCBuSOFE2CY+aJpPAZh47GRt8A0oqqsS4y7CGRqykpGc3N5pG1E9FD56pb9ow8jANBE6efLuW
033BpXegj+VhHWFOReaedDAOdhVm8ZYmSVFwJvvHFN4GxQM8wH8mqewOr5qZQNIwueR14HCOlck8
COSx8JVRsNCRc79gfEDRSqaGeD9waNDSbb5oabKwFq7naY2PINps1vk6qAMo19k4v6yNL+bE0lLC
7Jee9g5VmrHXswWvky89OFXn+RaNoJr8xTaCl6AhV5RNmLE8U2gpZJOPzelsrRh0VWlz0DH7L4UI
1P1Pn6+zEUxvQOVDb7yyRPf1otk65VyHRzcOjtbzk8rriEd8fiitG0tsiWKut5oXLOUL5d80DXsD
GSJ3Tjxl8xcpOgK/gWE/x+LoRtdeKRylg+xnUNzNWPEuNXsXdCmULlUnp2x4ykGXWgoTAIUOyBPW
0wwCk+/YnwFx25FjZh8ArigTbCbctZSYTAqTusyh635QFRSKDdf1iQJoFluWa+3sS0wx8cjh2rh8
MetZscnboPSzW9DgWjwerfWxon8EVNC+yoxhHmxbTy/0KBmGQOoVfCkfpJZN7JLB5+UB3yXbVzOF
Pp0A3ee1O9Gsvp9w5E2bztnqw/d1k07x8jSirx59aFgkMNpwRqbnv4bWlF0nTZ0nRDLLIk4PmOMi
RcU1T+xFeUk70JOXWzVBqDRPwzqHHX7gisju3eXMnMyekB/fQHQrF/blc9sxP9+E6gHjX6XB/xVQ
InW43dOluKX2Jb58BJGigHeCvVX/+aEpfj3aGbT5XQ/c8Xt9/xmPfyUMZp3d6CPioEqHfhbxph7X
mcFJAhG9E/96AVeDEoY+UTRUAo9wSu9/my9IvIapAyluh+sZqYsNtoOXONIqJWZ6WiTgRuKK2lU/
UVTCHaHxTdf/AubEuOY8qhl2d6xJj72cLvhbxfOMDQTUj5pU/uyq7I//RSMpxbjoRf/sQidfeuYp
lMwMXB33fajOTfWiSBX0sUj75OLMUDIvLP6M3s/4c+SUR/2F0hKuG8x96kOJz/2SriUw07efv2eq
9z2C6vxJ4Y0MDb+IhXjFkQmRB6G7lCNxie3hTQ/H7y+FwttAM33VNxv+6wrcy6kVi5BKn2Qdlspi
lSMaMjbX6DJEmvIKCmKgeoPqBYsen8VownHtlzFba4bWMB8dpYTVClL1foB+g8JCIvQzBoq/IplV
M9UtBetm12EHlKpTn/e51N8Bcqsz9u4uqxjLfMK1rvvsJCCGz6uZcrBjcsqFvKRVC6jP9rjN0/iD
XsqpZt2inCSB7ZGMZCgqn2CURoEPGNJqAUkSKq1qB93jHh7rLd3QIWg34MnfbQ9wcXcZ30NYYs+j
VlQB6MzlAPnw2Mi/iyCdkbV8FPXpVAvV0EigNEF4WWystYF2tKVVp9LGwEkOy1QxXYxZ3PeRFg0t
Aoah+k2FDww0VFzKKlWBSI4eAp/I1Yec2y2BvhzQr93qpTXt460eRlFLPVzX70Gt0/WnvM12DGNy
5S2/gO73rbhEQ5SE0IWYg1xrIcof8p/llknfbTsvUrvowLSeg4BOMIC1/TR4vw6t1fuDwooJeWTw
lq3AoT3xlN1j1S0ukhoGDj/z0znCEWnfQ3bgDYdidyPsi2ghvxljazIKA5W3bhuvi42J3Z+LDXov
9IZh7kPSoXxWHxSCUSfS4r4sGOW2jk/GWHB5z5lOfyy1jamaZ/G2uz2Mxwzq7j/caLxZdahSh/B/
fIqq157pVx4XNhE875kZVwhFeU8F7GExiFRlfnKFpWDHCvEl94SlUx4+OqoFXgIVZdVLKRF49tnR
VVFU2ZB1F4OUH/zYoTMLfxFPT8y0GrX6/NRWE/jBy1uT35i/nVbu+x8cPLTf6D/HYWJekz6DyDCA
WNilSn0mS14u7h7eCwmcNxGWvdh3j4/wvMWmckYC5PUsLCmi9vuNFFz/bv7t9EDi7MSbJQP5gf7l
CAG3dT138IgLkIuWLbEZDaC9F9LQqgyiQqEQjmVULDf5FHpErFX1Ste/UAxJj4KDsqPcCDtcx6mq
X+1i3AXEZg3rYDRR4fOi5TyRYXuzJCwFD47vbDg4OYtOIfe/JIDXPoww6PsexPbjeugW2FN+bVvK
blG419hF2KEDU6aIFAsmVa6xFgQjdhC+vAhA80jvtF8JjfHkADDeVZWgfrkJ8D9xGiruR6l0ZDoW
GtS7PaWL7DRgP+D6a2Ry8vWh6zAfJ3mvIyFLO1aDp/vpK/W52XSpIdOVKUsTUbTQvPAeip6ChJKv
yuLVSXBd5S3+lRx2+0S3IEm+4Crr54KUkblAIdVc/z3CkOX3ypH5O2obC7Xr/k5To2XprqHam7KP
TBrMRYejyNCTfxsZTJ+s//nRuXeV+UmOf7AxbonfR4pCulRhX0hbIBtCDNn0Hv5I+NPl/QgF1bpY
ABcJ6bRFeffxmExPlIFJco9FnXlsp2F3ZDWKSaNDXIzZ3XyZ+HZhZHdzLj3qX94me6kNrjLs0O7n
Md4Dr2XnOlzmZOe96NiddAJHuqIrj351njDruwyczYBEoRvGIncStV50ONhLoCeqthoA3BN8IJcx
uGAULAtVo0Kw88I/9SOuDROhWGEtky7QRg66CHsXjbRTs/JDWUQ3rmHR6IVdC/g/QjWbJDTosh3m
/zD/PR3rOS7mClTQ4mWVxgNjqgH7ACL5g9pnihVVJ+zltUwnihHrpcGeJoMw3pZU5Xkmw13vuaIw
3712mOxUp+D2zekEh7j7BVKFrEqErr0FrYrM6OvVF3x4CgNTgPu3sMXerGw98bFhglkEa7jGUUZ/
T2AvyEV6GKP1vXqIJeakhLyn5gIhKfGqrFxyBVSE2DEGYvv6dBrJIwC7BN3e4+6Xl4QfDGTeVT66
Cb6CJSg/ymLIkPCzgcORLQLG9AA1PJxRSRjz8FSjBqWJHTqQAWXS6d6SW2LI4/NKdder02Vyadqs
GvnNfDoNIDFdLCDCiv6ePcXMAngQA6jfDGyl/Qu4h+14Tj9w+oJGS1egFUdR1XDQ7TaCbyNdaoQc
3gA+8elPmNWLxMOUSDY4qlxO2k4ulPMPaDO1VPX89rxgutVKPSd7Gq4QenY5paETYWS6qNoOVDNc
nrT7jLsklrdmGWBT2FK1ObIoXqUWK6rpZiJGF6e6t+5O8sOy5z+CRDsFrzNqjMnBqhvua+lZmjy4
nFcAC8KIvTGl3sFfPnblAKk/FNcePgRO2M8ceGAKOgzIvzRGFtSRsdZbIcjyvO3/kmt+MUF82/IB
dgFdRJcuDeYvckudqArs2euv41OHs+jslqq8Wsib4cAph8h3Q3ukzxbrYhT54CbrZGJnZxMFfEOf
Qgxenr61jM5xF9kcyxRC/HDnRnzxSQNjueDd7zqu56HWyysPVOYSyns1liXf79DhIMzY3lgfl88u
hoQkH/+zWEt81VTl7LtfHnG5PGU5BgdCzbYoplxaL5X3rlxVOoJj+HTX0Uy04swsaVWByAkFexRP
qLzx0ORzkTdYieUfJlGb3aJNAHIUyzqHGP1c30EnCYsSfh2rfD0KpiB/bDEwQUaVVfILQGQAQXso
2MqWwOKvX9U9Js4Qhq9Zx17rObuGXsO2wWTtkZ+YjuoAiMEDY1TJ2Ks2nCWRdEr27HseEU0/Ch37
Tg7WgBMf2R5Zn7vt4QuTwhU7oHsoxrgTo7816AbwyZ1Hga7Fgb/P3VQ5cMbxEkQ1xjxU1Bfot49J
I2StrQ6X8AiUJvcbkpfu9yuskWtmzSrt44wCbiKyR0CqUFzVcLmjOWP8jCUiUYxyQJvAqIK9ziCd
yah5dREPF2vy1TPPv8iTod71XrJBIuH7PBnvMAu2VbUsYHE336h0X3P75vNe/0eiXYz3uHyg+a/U
nOP99kdzLZatPJaEwN5WFJKNSHZVVCR9yjwsf9We0uaG/tJVg8XpDjsn8fbIDR9AdMNbouEcnS/H
o1nnVzN+fiW+EfHjYm6ECHSjjhIHyR22ivIwyIw/tgO7qu1ALK2FH+5ENVQ2GnrnpVMewIDVkjNl
QMvCm6toQTFHRJPZxhQS8NjobejvBZNKx6SbmdflX+qcHcMf/yrDGEQoIYO3nXcdYGTluFplChZ9
lvRQ7QM0e96oW2YisArL+FzjVQg2Gx7VUjaRz+fqHiJ04ZAiNfwA6Oxz3gFQ43+3nNz60JQaZx20
wD67I0Ee8XFJp1cfbvUOVxeiviU1qw0ECBQhWvJdm2A38FV+9t3DP2eZvmS4ojOeyZsrFfKwSKeH
Ppbp9C1iFkraO082BTdLfDhtDuDviBcTDH9rGHFpcMB7AEDQEm7gDxjj8lxxDNlOVJ3UlE5/FVsR
MJILH2Q52L0IKnRzlXquko26DryVZGK9qHaVou6P1fmznf8SyD1LPpEIjZi1uoY4zxQTvWqshBXr
z4BOq+fxc+QEAXQKSiVvBvZL5fyvvQbRGvCWRx6XaEwIux7MQa90JaMfAtvweAobeYEF+z/un8qp
kfKMzn2N5JclG/lJ5krbvB0qvGjtyEYxRGjf6/9axMbV0930AI1noyu/LmGMX/bvDT5KkRZIdfPE
ohdRsct0AHmuDAHNI7V89lgENTwLb678H/8OV0QxAxAn3p27cZs1PqqXPxD7gz+rzvkuqTsoYswS
7MC4aHsD4oMLoWGanIxuWdOq+PHUzfdO5/Oq9Q4wTQLKjEF42dkckWbplccwy8POS3jYzpjUPRwJ
zK8FVb67+tyHcL/inFpXUZhEuTfHXKZESY6EttKTtHgqy/EX9LeBc4dowMFufBPXPyx+0VRAe6dA
kAOX6305kMftr4v4ABtirvMT7spk6Y+qJhYDRsWJMl1JbwPPsAwmuR1dvTRrpRo/72JRAUMRVCmY
am8tCXSRgxGnEzvCR7tAmjX4obezEXAOrD0fvSJnG0skfwsR3hu3AWfcC2ogwR7O6gmytCupQ8Jf
QMUbZS5OGlUTEYpr4bCPjwbgtR998N5vKo19wFaJ3MteuaVFyaUQewgXVljXZIoOOvpN5/564+SO
0PaGXSQp7Cq6wr3SIgIQZ5OJNtFCzXUCPNWp8Lvojv7ESQrOJWzXjKhkjFpCifA4Y53p59mT3DvY
ILkO5DJjnxuBSbH1BBEgI7A8iwYjDNnPS3UKlA6g3Us0C2s35aYDRNhYyNpRKB6NvJ43ChJrY5Yo
YuQH9Yvrk6jM7/nubUENdy9921U7kHgNsfkl2bYrRr+Q3soy41mEk3dTcfSGvAHAZvOh3VWMvbOD
CHdNEGVYVDo5RtuStqtaMgC/kDQpHtaZXcXq+iilOaSTKBc8e0bR/nCzANern9M36nqnG1v6QMQe
uEAh8bxV2dv/wJR5nGNxdCFS5/W8TtWICwQdzn+zxo6mVJ9wP2+wC2RL2J1qppv6ikPavlkw1ICm
sex4wHZSLpqR+K4ibNm1daGEmtlL5DpVDmNbgAcy5l/LiXsXT8qvwkvZ6HCdIJPxbqjMScJRbuK0
ofLeGolfALMsHbIQnvBe4uKisPmm17knjVynbjpbbH3VyuAXq6m2VjpMeRIDZxdBSl2zfxaMl0xX
aDxprElJgGCYq7VNnHLfofzCyufnEnes3l7WXfq5Tfl+xW9iOXw9botKfOvXefSwGIvS2RkC1lfP
7FpHRLMA9ckyZcFJLr/VMemurj9AjG2bpAFgDkH4pXNB8bs0bPn9sYRgtkRwqnkmZBtlNkXAqBjJ
z72uycutisTo/PM9jf9EqAaN4f0zh/CMRnGfrd0qoVd1iTxG33EQ64p08gyPrJS5fSiE7e/iVG6y
ZKTXJX7TVQuydYzSjVfGkMSmv0O1XXY26i+BKd1/bAeNQobpMaHCORNM8peEd3xNi23/N9u0JPla
ZF5iC4/O4hvm6Az8X7U0fWVMoyqoqPw038xKuQu2Quj4TTKL+JHGAFoiCyaMFbfuOLXK9TsH9H84
zDeGLXm4O7W05Ph6YN+0LnOdJYM1h+sxqBCJ6fhHE2VQDkUzi6Eq4aZD+dJgryUDbh/MrnbFLU3S
Hu1Qh1SLdyhq/NdKI1RsXd90icJqwDh8NWIBMuijUe/PUSACaIWjeOwjZWKazXcX4fHBW75fXdxW
bAaDNugj9IskS+gzAeWI/bApNOfxeCbSkOcemiyY1ELbVmDTRFOnu/h5lpsqhfStyG6xDu8bRt74
a0mrl6tku2DGz5rShIcyBAIUffIMn7rf6QrhRRQYB8gmAxz/PGQOs9Z8vnkghxxstiWg/l9cNMaT
v8YMM8UigfoCCkaaJT2wwd5a7066Dd1muQMkBZwPJ6r/Ks2JfrjIbII8rEOX839l+/86M28epvOb
nlaRNTQFykP5Rsj5L4f4dS0ggZp4OEj6uSRDwDa6jIL+mUm0StQ8EpUBJoe7h9DRFGHQm9b+GPCA
RaWXqTRcHsFwm+ca2pUQboci+O6u/py3j19FWFIpXFGxfLyPXjygo6QNKrtt+djS8kIgbclwVxWS
VRmHj+MOiUr6N7QP3lYuRsb8yRM8KSVQ9OucS7g+DE5Gq2MKQ2F98nw7WUwoqi7LgGYoFodiymE1
tSYdTW2C0zzRrsNjlJaCZRJHkDoAr5r+WpTD/Z3v90xpkTsQK7IXEu6o3xWnOQx1swSNR5+H2i7O
W/+GeKFjYTWBWO39TIuZRIumtJuktNq6LNIRxrCLUpxrV2ZWy0J87SsyKC4qCqBlrhfQERglJlS8
bgj3zVw9qNM4g/iO7hqFF/8PIj8HqVEIpPF1mhzBG9aY//wFQMolrA2CkAThCqAsaN6xBbhTwGQw
WTJ5OtiAJQXEI3oDu2PQrKzkqsyFX5IKnh0Mi1FlO0JFBOe1cj6WFqINBMkvEkUiFXgfSt7m8Ecd
cDyPL4RaG1Vu8nJwlVsvhT1OU3vuGkKwJrObQFsutkmfzlqMNeA/Px+6UUcJ0TG+6Zw4RxxteHiQ
Ekg2D9UeoFnDMw5H1KKelvIGPelfSUah65d2S8+WoEvekKn2hjFpeTwvmWiOKLCYPhqfTVLAUv80
n0FM/BKVbf5GW4yBS7h2b00rJfwdL2+jF34TvQyTEAuYMez0g04lVcsmaSCMww7kdhInzzWlYoJL
LrvamrWx5y1g9tmuNdcl49QkjlwTU8aBDbgNj9mPrL7NinX/4Wp6l0YgKhAR1QCA1FGomJ4q8yyx
NBkrktijj+6Hjd/KsvqE0FJCxOy9X7cs2isUcR/zx1Lnz1AnxlDmF0jqVKxEepG3bOVs8E/AdYov
8QrgzNPEBdKp3nFkXnXlTyaA20TFcbXuaIF6lpdOR3oiT8ZhHjqmrcNvu1mqmkwewx43p2E3y+Hv
j9WLVUO5Y+0i89bQJD0xKND8KytmMFAM68vJFE43Tke2zWSIGzihTYLLqebUPxQmdeSmKu0EbfVA
D5t/ah5oUjZi3INr9nHJBxh5Af6lE8PfX1qGeagLYcw1p3AYNLD6WGcSvlakQa7cR7I2sF3773nR
FU5Uq/MB0bWik9Q1XzLy+yJaFc/veMnQ9ZYlYuAdULLZN9CZ+1w03zl7yjidoCLLHYbbDipgCFpM
hs7KpVwikg2j1eomBn0SXLdvVKlw5lvZzi8e4mRk6tmMApNNTzo6zqcowMtkfaExNLzj3AqWtDDE
7PPbSi6sugyp037UMOnvgTPB68h2MVHRuyDNwrKnN9CdVfDFf/N9kWghJSXookH5LOULMer0tk78
HsadNUpcfff0iFRUi5JnMqL2ZOo3g/FljJR0YE978OeS1uIzgAIEbA31ZgxJ2LCRD8SiH2Q7j/tM
UVi1pasPXRpdT4BGuzFNmyCzPFCQvXBp1X1ut7v0+wT6L2LdxnYp113zIP+Pdhac7X1btnWG/Tny
oqwSH7mscOeHGLTHDYAviKyNYNSlaCcSpBS6MHpyaPrfsZXz2M4Rw99SaeUZrZ3+CSP2lxhfuiXx
i6Y376H4I09NvjXs3Kcnf3O25Zp2qSJmoLqqx0sI/KKsfEPUlkD9phKXYTKAcidyCir0bbuFaejt
j5iw9ulvodt0+jCQ3mgTCHn1ZeOMOD/gBcxXvoqCs9aqY0zWwxLoEk39pgdLL2CXRlNgSRw3Iv5P
LKHbqg8w7l0JBytJ1jsP9Cd/Y+VVkg8GhveH7rgpdXZLGAcNY2RsAx+3Um2lBe24X/3/e7vwvQaa
hOtLCFDvrwMkSpaIlt4Pd2BuZmLzEqUxH1y8t2rW2A8Yave1U6tbrJ2dU5nfQOD9iaXq1+PbJuet
BUS3Fy8J/j99bNE0HBGzuvBqMJ1Xzf04f2W9/se9MIrAcKN3mQ9/0tm6UoveAZVx3Wmykd/1DWWd
j+MjfiHXg2FsKL6zmXmiT6y2xWCXK/vlAllK1heS6jRB4I75Tus6UYw2CaAMAxFh5h2WN60AvmLt
6GCpui/9wYomExPzIVf1pLtYx7B/YnCHb7+DT0DtbDzrzAFRZ7Vqkdp02G2rIfWKgsJY9KqWHk0s
Br/DeuuOMe+ltthbSzXvkp4rbTbR5a1VszC/nBLyFdfhebueobpXIpq8tkRF6nxAZ1XZL/4N5d90
c++hGWJ982IQMt9dJWMKqVMKH6MEzagn8YCtDIebu09Gq41d/EkHqxwF3juBRDx72N/E1PnmiYUL
YCM+/NjSAsbJSEgvq2NGu7Sd1H5AsjnWsmjLccLBn87ZuXUc4tISPUuItWSp3GLH1LXvuxq5OezZ
558PGkGFixCfLh9w7Iq0OW8BimGG4OgtLW8ZVLSs0l3gJOCNN0nTCQl73TKUdDATfZ+CHBKMfzag
4oJKCg1sL5OLSZSZDh9dY+s9lNiXLlFEYX2xlxo91+++FGbgjNjKx1mjbueJTr07MVTuA/kGDUPD
wUzvJMyCukoDejv8/TCsFYZsAX0vgRZJyalOz2edG/V2PtFptMzYQoYSKS5gc1l6QRHqhBeyUhgm
qABOFEIqpFBB22Ix/ztx9g3KIvTBX+aGqkvZ6Eavq8Z2iw6iJoGnfWdj3YRL1a3TxB4VQaxXB5f1
QX3ZWjpixt0VhMgFpRRUrt72KScNaQMnj3EhCLQhOY6pVNvM5PGMAaUt6a/2lSne2WaEkbduLuFS
AdoE9LXX1EJgcsJGKPbeKCTtqiwNI5igO2tOzkZdu5xdeUCUEtTAG4b0z9vWPGdmrozmX+wWvf7N
Toms1fbkxaC74Za18TL4wXxvidE8FJoB5PFPYZUuqNgmrKjJM755uSFBT3+wi1whCM8qfSHtsUWo
5jdfUwHf/9Fyv3iU9YxzbS4pjyqmNAn7OganL9rqzYEjjkh86NYYsuahij+LjggEe/r733rMKBxN
3S/kL25Se8uqLgImRUP9JgdrSfGlSjk81XpjPAVAwUwJg1ZsPbZi6uIoknLTddwbEVcIOk0rg7gF
iJNXN+iOapyaiEFISFC5f/2oYQt44qwdhMa2k79S8Jcyta0E4/WII+04MsfltWzF8WKIta/B41Xb
FvIfGtlOJjSuYkhbTtGfNOGKKKePj0lb2JFNfDqbKtj1zHyZgLczlICHI6dyk8m3qvjaFrcMv3KX
aOt+lUEbMBLl7WARwSQ2I4pm/WT47F9vNjRKM9YYvlNvxq8kf7+Rr2fOJru5nTky/J/NSw1xs325
jK6KjjivQ+D20M/qh3Jw3GwdpDbc3wDJ43ZjXtzJ0W1qO8G0OKsN+nvXOn17DExQBvTxnFy9rrwH
7spd4sC8UMthj0RE8Xgpam3o308jKZYjEf0Ssz8NaBcwpK2TRIyD8sHFxU89r3HsoXaD8XYWj7q6
2m4efypzZmN666OsRczrBOsH/zmuRyoOHOFOhsiA4WPlXzGsVMCJtMXheZ247NCQ7VvuxPS4Hvce
IT6g4umoaF0m1dMGQdmh3jahLDVuT/a74/o7CQtZgZ8IkR79S0QXAq+neMRNzosnp+BbWbYX09z7
joZek7STOHrdH0F6+SeelruYXUmFUL2Er2ZEduyFcadZil+1fUiJpkqPX2Hpow0s3Fl6uw7TGhHK
bVnXUlLLRaQJlc7Fb8im5xyNXb0/OSqdhRk5SoAAl0JKCPMaKwiXQor5dNMVScEWqXPH9kXYFyHW
Q1dBFy1Sn0h6wWofhc8CnHl1FbM4bUubGDRBPjv0sLQWPD67rb7QcTEQlDUNbUl9MGnA8j7QjgvO
/O3rMhuMfWwqzpX5XuMAuIW0nDUYmvFHi+i0LCe5PCdZrhrKWHGMKb6UtJDfJW5gV46lO2ZJ4RK9
3CJMkPpjwRyRzrzh0L0rqd8noq0iSBVg/FNldDUqOUzCR8w2aOIJt1q5J44SPfAZuI0+N3KK86LV
RLiBD5mdOXI4/CUxxn6GbwxIN7lTN3Zs5R1sQPbUMTZRBplxrTPGGfodA/IqBLiksNfkTQJkYXBd
gRbdV+csjs6JpebQgJ9feTpWctUeePd1yIx1CEeX/Doa33vvHYlmlvAUjF4ti77XDdVvf4IGDH6l
/2Kw9VGDjnYPgSGZv+LLzw4XMI6u313dHuCkMCExytQWCLDEnb6bswo4Y7MrQHyq0xFlM/fiXA/1
k7Av6Qhvl3wGrdzJDPcEu7gf2taDdmPVzLVYHlAiRmi3Oi0jYjtUzOLaPtoC96fKqn9TFbfI9yVg
Q7WsGynBpFJ0/dwGqiXEJaRfcYCWRmY03tIb2yDDHz6EypoyiQ5I27RuWxahAljGbYv8aiTFmubV
d1bDVsBPTA3RbodikrufAdzbHcKJ8/wT5N58AGVLhc3Uox8HgI/++uL1pYo3PVKdeURXIxcwMKnC
LeCDkx9AGzf5WMKQvaW80EMnN+XThSLi6xgDEb54pr2fw5Pfn0y6ohYyL5eFlPPJR1Ciy8MwgaNQ
6X6gaIrxFFA35XtOLwGhOd0SIlrzn5qn6wAkCpfZO2GIZ2GSZj215BISXjNki3rzyWgkcmI2qn0Z
M6LSkk59b51MB8SEr2ekrSqTL/tcOeAffKUAuTs3LreujQcvax5MvZLvDZ3ANOujt6fg79GlbG0Q
UVJqbg7NGXJBD1ar/Rprj3BHglV8Pktf3HMvHGwXaqXfaSIGcE7/CtE2rMcd9WNBRi35JqmTpdRj
Xkv32qjYGwH/OtY0E6sRmwqc/Z1rJ/f8987dpDX43z3zQmPNpPbbYZzKgtltigdgbAXarM6irGmG
kuupyzbM2EjvvpAMkTONFs+d6xyxajWHIwDamK+gOg9ZtBT2TAG2kJByAV23kD8DiAjytIpypt6e
3B/aSl8z7wiCRhWbL9ZzifkzDAT4FOC67dsmpD6tOAgYpQMTPwYNrI0joLCgt6klXgnZYItXt5tH
I+fSXrwnsex4jv7jqAA3P5D6Qf/oTlPtoGHwjh4UzKzsJPNEYqeq1Wj7N/tSzU0y1i5DHBN9lZ5s
bjGgWbEWgFT1l0eC3arJkBZTPl2eDhCt5NTllgweIXRHrE4KkBFmGE7J0V5M1Lpd7q2Pt83Sl64Q
wRAqCmuTuAh44LXrwImCwglhzhW6yqHRsl+zUKQ0g+ISBwSIdeeTP+dbx5RVxlp44rhQ9wk5+I4x
9Jg5/pyCYrg2vSrcCvQrHZikLIhmb7+NTO2GZTu8dKXOx30NZj4lUFfvs/b88QEIEztFQ/+CLXlt
2TDkWEvPu3+yucUVcyToGNJNxoLOdks3oKjjWR8JWx9zlk310ZnmxfoWpueNgMOw6fhSlhfDGJkZ
/GDw8eDwSae+abPh2L+kBW7qTekSqSEG4JXo26ETgxwRGkW4DqZ/wGJvrDsoglhowAxXzsT23cdZ
mQ0ZYXIH+42Kcu4tLNoQpxjrIRxugjulQ4YFsKXjHOajV2HGou+n9QyZ5SNWhfp0b3fqYMzSKwO9
2pMHF3jga13HI9ZTnKp5GTxEuVTE+wAEY5EkaHch3OtqVze2LTDOyHvxegeyrVqm5zLXrOzgtgFr
9drXLOudF9tQysb93hRPhLgMsfbXXxnsVWw+VEOC6+4/C5VrnuhrImjG4bCr1TWleno5hZBcSR5E
g+CV351HPcVMjLHjEaS+CkCQ2/or7O0N6Qk4w2kDdstylOYlaurwgw5Pu1cbvT+Uza2E7O8UNK9l
ljuhMUJ1URaa0xZ7KajxDzLGjTCWyKFk/4jZQHf7oe7AketMUawNpzr+VvRa45BzrVvjBnpHIKV1
uyr8Eo4JikcE2TdWY1kc9I33Qpi33hmI0kWa9xDE9RARL+akRTyh5IPyNtaWyvxhuLF9a0tWeu44
cS0H+ozHrAlogQy8r4BRgu4jjaKgy/0LwM1i0e0QSvW+fZY+3KifVTXTTtYwsvIJp2eB9sRM9uBY
6oItJhYKdD2vPnrtaoJIFomQonAcEELjrcs/AHqEwViYpmgWxmcxCdj1JXqzPQxcL9S/uxSNoYAG
61bWtqg2zkCEmkxr7+9nmrCKzGFnfAUzRxbCGoZlhGvP5Xs+FO82R7Q87O3NYnf8EjOzPQcWMRTe
s3umT3KTImHbNIMuLRXmd0y4dHaIOgVfh3MqMaoUXdXCkDdbDiL4Uuv/q09J6NxRwYon5lq8FnvB
/dHzjNbDb5boEKbWF4AibzE9B6zpeuoKbtd9zP7I2z4FZu7U1IkoHk/+EASC9KoZ/436CpGyDfxB
DoT35k0Nc5UB72a06lqFwOY1i6I2TGNNXiwPwaKOHiK1uErZtjUYGaLfnU4UsFvwenY0xgRo4UP0
Bweqfm3f4fjs3Q9CDIMpZ8zw6rxs6wl6Lvw2Z6mawfH4DQKlnjr6pufyu855EAUgV9Y1iWDvK6NJ
cOdy7VDFtj3y4q31ClKe++fVJ7FBo3aCPttI6aVzFLlFlsrEkGhFng5Y0H6hs87QbGipFN9SGl0+
Uxq15CBEGmF57HPf9Toy/TObiWZQWldFPrXUNvYvGx0oquLys8DwTZhKf3UHat4Q2mmIxfQIQK7n
PhbdhiMA2pdMt7yBmw990QSFDaRcjEePGHyw6Mgjx3fNQ0XA9yB6WwOyoZREBv9NfAoBc4qoKXFb
P0QoeVly9QPj9+1HH5bLHsoGTV53BJorOKjt63zFj7eXlA9dIa4oDLUW8OfsWaVze4KBRiBbhfe/
7CauzeQ0AfmoGibfiXAz62B3+pzz9tbtkYJQkyjxTFJmsWhTl86enOQvXiWA6dzdJiLVPTyDEGvW
HBMF6b3GFNpXBi3+lfPN/ukjkz+yGct++v3KLa4/fiSvZRCy86IXNUdrNndGVhYLdfLX9InofHN2
XXg2ta/gmMQKa4WNqGBnFI7XJ4YmvvoUwCTTJgCUntfWTkLgdBLSojUzjL/rgPA3wN4JpYxuZrPI
wkPH8DGBax+pjjRT7x+7RCxqIDAB8xrkGHda+OAlS31E+HWQOfFqjkSvjVilRgxW/er/dkLTjGru
RHsNfk5CYxYkOPhI6Ori0S6eXu0u40jc8ut63u2DGMOFIob5FhNemNT/dk+IrHS+NdXB36znTVeE
xIUEI/I7sk1D3jq591z7aHdczzuYCOR21KHZzJXDVgt32U9SWs2CCQH1Wz2H9Gcw/uX9x8rlIzxf
sIRS1SLC5LtnylNSAcAoq1S9SNEMtExhxQ4kD4TWIw1X+/4qhue98l46djGvxqbMtXQGFy6tSYns
RoCcpPJzqv4lhpV+ofuIs9J8UWn1ea0hdEVh6U81AjTbg/OK0/W1j/STMy5LJ9bZCJDQheAC7uzw
fAG1C+zlMfI68TsdYU9NIm/el6k8qfPQWHG6rtZWoHr4r5PJkIgCf21hrUVUroZrTQh3iXPOubPb
xgh0d7P8PUNv3z2nAkv2hw+ieKksIlcORcErIRW4txUOpnfff48t0mi4Db1vFccOr7XxByyIcFMn
zVKco/A41/DGxi9xTgdbYwS90AluzbT22EXhFSvSDGueVIBKqaCQODuNJqfoxKeb4tuu5Kn9ePRa
5udcRNooYnYtMr5ccfmN0n/QrfZnWRpCzHdaV0BATEulpmG8v4Z6SpV4VWxcUxATcwkI+v+Ooxfj
kZyrOXkw9H5gfqEuyCZw7Pvngzj6Zw6A2exHFGXf9cp3YWNyGRjC1pm/veFeKIKyr9Rzlc8tH9wR
xBZ0veusY1rirDOpGxzW7jKo0Uq/Zqd7GxA88cRatjpjBaiN/7P/xcghrqi58peL1nTUKKM2PAV6
Lg/G9kCZdjwbHhq34M+tI2cZIXQ8o67RfkEcg6BSo2aLz6vb8FNrsl7+
`pragma protect end_protected
