/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 848)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2qUfzJbnzIBt8T1cLLlpTbEJChoxpvkyvQ3kG8Z8QfBB+plqHeaf99ZS
UQ1Cvmy9/hz84UMFlitbGwBU+0JKIvyx5lmmYKFa0+5w1RRly3acuV4G935lFWMtec5oqG8aKlRi
ZKKiI45ioo3j1TrivvsGs2fKF3BlVQDKByV8AS8jqYM+31Y3FDj5TG2IfZuMGbKOplYytC/knd/K
j7v1Yc3Tpw4RDe/UwO56J8qWFGG8mSGbS8cxSHI4fuF5VlcULjEC3+6pJqeSBgPCAhFD0FSD6ogR
bFoV3zZvy26LuG+LBJe/KFKHgAgais3ZPDzcP6dec5KpQbqLWAgiTbZRm6xegBTdL7E/jkdKiCob
GZ6+/J4PGMwQDnj1fCPxoxETpBQod324Vz+aFyvPqPRWS0dBEtgTqPAd2dhODT17WohJhEM4/o+t
X6Axrz9geR3K5VWsEj0tne8cH9yHEZsUIbnnFfTYl06vzTgjBnGPATcqfwpV1BR8w5+2WUAh1wrP
ZUYwTxCu+Iy4PN4WbizMHYOEBr6SAFoNlA/4bcjEAgBjyfynFbu6044sv7TGK3TTqMjQ6BO9GBkm
H8fNgOrwucQS30jffva065uL6YkJceSB0aFuit5lh36c/FMv4Hp0cRpvdvt3NS2ZjvNyk1KIdOXC
B9wA1f7uSswqnWMBdUVMiteKkawuOBq8LuB/NGTWZhwA4KqC/7SCFxyjmW8lOdcMQOSi0i7ftj1/
PF+LLWtMXUdutk6bQCXZOx/kVwTKEnWsF1M2BpjTxGt+x6U1+lKgmR4lgpyWrRtfmsLLCWmHb2es
jZUQgBdnG5DQEgITLeU6dNalHOuuUouP4FgLuNUF1RlOswxCAy2gzvvm4Ul/EMo+l8w0NsiH0367
nDRzW2q6IRrmMeXiKfxhUsDrmysMzUbgPvmLT/9uMZBcW+we2nI2eRU2xJQM2adI50ct3YI/wdBB
L9NbsbuB+4Fn1hzW/EgZC9M+GbVBQIRt4odyT835meeoqT+DoEJ+lRcEODyA4hIeW5MWlqL2/zgb
AGQOSn115lB4bqfwAQ5hic0trHDa5kCrOUdniwN3BvDlg5LL0RNOKMKFkMmprib3t8M=
`pragma protect end_protected

// 
