`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43936)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPalmpDX7c/wz9lvXVan4mBmkObIYbC+57pMXxCA/FMtQqIy7Itc3olDExshcha3hHClTrHoS
NvCC7mLypDaG4xLS/lAsBWbvqJASsEXlPgfA/uZtkN9v3pXVIzWSz022W15nGqKIqdF1YdJfehTT
T9/B3OyJXQZ7gtq06S5mu2ul+xrBCpQg1E3OW6p5YUlduYxgS5KUy9oDEFb4ZyvmdsThEqAZdBjb
hFyQ/ITabHjzvH5zNQNYRCEjbzrsO8ruS07JVCReUYIBoX4EHpu4LyR1NBO3PltQM6G5dPbIqWna
oB782Vry76ixYYvzHhkf/zmrw3fbx7lGqyNbVaS+gB3kvIxdhzVw/xO/5Mcwn1mGTGTOJn9djLxF
KuNrhzZsL7sOntOe8dXNaTY2IiEcDbP9ideZw2TPZj235SXBTkZ4IMIlTSQSaa4G8Slb1CMWe/aO
Ue+0l1x5QMLrr3OmCo0hdmDkdlo1PddEeJ1eEz2qUw/mnUO+yfh1RsSQL/ou/xLjsyCdNX6snfRZ
y1L20Kq0IdaU1FxhDBxrkJZ35XuqGNXSqWaiYZeO5yw+4XmqbOqCjtsSSfprd/xdkaEluNC6+qqV
bTAwvcXtGqdbOUrgNxZAULywha2z3owaicuskuaVRMkxymjePftAhwxGVNWK0iYD+hi7VlzjaEdz
Gm49zdfklRQ992rbI9VOM+FO/avys28hMIPEhN5S+8IUTF1hmby6GfjyumkmzpUYJVK9KO77YaAT
em0ojMdN793TYkG+r8Ys7HCUS9SDb6KIOrggqNFd+Vz5oegLCZq1FMVd2L8CqDNB2dDDURr91jyK
Kf/CiXYCZnSvYHIt2U7iL2DSjSw/y5CZpg4yEiNoizKjvoM0/H7aaoIfEF6MpjJCGlCofUaD7Wcr
Rwo3rvr9eXSyn70g0QeLXO8N8rY1Jmt6XKRjpbsuxzZr042CQUPXzJ3qCbFiVPd7e6RrsOwdEjTx
avMNDaX00RRusTeWDSP/jsCg8Oa0NELdoKmTCaCr6z1B/HzvmS5xfkAAdTDE9qAj/sif51OYExPJ
lFcsAbpGcGw93LoEEeBiDGQKY19/O4vcPu/DQ9w8IwUYZq4aQwydRpyY9M+iyqSgBdM0mdmU3vtM
5YAtwbuZD36PPiaMd4zxfcVzZ+7fbLRsOg5HgAQwNkQlhMl1bQ0oYq6b7Qtes6BLQ73QVTtSMNwZ
T7rr9XFNfBUZ/jNQfmYn46hgcGKUDDOiLVJ3TO9WY1jXT2Fl7+Sw4u2Caqnyo1CqDMDs5bkPexCG
avpGpwBckUKdGYMUmM0D1agLLO3UkX7a4pGDSKsixBsNLagG0/crtH5PmQxZcyBRJC/iHj3Fl/PU
LA1kunSvuJXqNTZb6/pkNvskEvuaQVwC2NHp9M5c3/XBcxE6edn1CAmHr4wpJJHPyG5ufA41fe4U
OfHeBf2jZbQttLpReBDWL9UBqfuzdJI4HUsHj99BJ992SAsNvGS6z5TIPJoy8HgI/+XsIXKuznGz
dmgj9pUr5syk9OCxwebEPCJ5OQdP7bYcK1EcV5ovUZVNS0CPHOhRrPww4qiNBzeLyo6O3xzZ28jj
8U6vAnb3JKcWwxg5XewRtwsaHlnfrdYFZ8W3IiACbE/AssOdvezAQhmICZBtwJY0/UllYSGHxm/F
C3oQlJr2WGKDon5sqIC3WH4bx8AuQoBpMwoSFxaS5eu+xaxyz+a9fu1Iknq+YHT4RofLdRNAAYo8
GtqfwWW/8AO6eLsOVLnAj2EHQ74N7ltjJyAzMXozTYvG9BYF5WmKBpT8HaLSwo96In+U8SRi65Dm
xMRYoCAP4g3IY7G5whnBoMCUFl6N7i4tn00h/CUeZtmGAAb+PnYzS1gxnWog3rx05WpyKgCXv+tq
hRsgB3RodmFGCLCeE3XIXRGgPGRWXJvWXfPdT01rpqzSI+lxI5F+gNr27kzMW/DjPNWBb1bQprem
ZAtt1l4dNMFuwvz5oY1Vm7wqkzW21cid1L+JWKWcZJgTAI7R9+hhMvvW6Ej0PVPskfhFmX6yiPQd
TfL/ltqM4zFonUiwUGzvVSbVFb7w8jLmm1DNUq0HAQzSWqguJJjS0xUuUYte46NIWmMHdpmY9cZN
WNITSx4gSjR5Y+orp7CvwRukC5MS/wt6wRanfvvuteCiFiDo94h+C1G3G5Nkkhj22YnrQfd3rxNj
XANzhuiF6BBst5bBUxh5PUIGQqfl5EqSXgBFR8wV9UVKeuNMb6MCI4nWDL0oj0Qk0t1iQ6Z7RppJ
/U2LYw151hMRnnVW38MDLA3SfQKdCzf/pZ4QILfCIxJN7rm8WPcDfC/xajqtefoVHMBkB27nsKDN
UABkGhhFe6M1chVbbDvPzBIwY+hiAOKP6xX370JvI2FEbkUXSBi9IPQ+VOq3Vuu2gjOnMkpSvehP
YzKrkaqdtUfpdczEDBADJ3+UQvpgnTpUUifz56qiVZxvFEvnvbjRC4kGrPv1u9cb+cMigM24CwPM
1nK9cKIr3n257Eqyy4oKKNlAHpSYUUKjT9V1a7NmkSgbNw3XZJOtTeSO/lZdF/0yQhxNkSs8Wx8v
fjQKYMQo4rDVU7S0DXqEUJlFU+7nHywQiAoJr6YgWIksiTybJg1sfTerETvD3nR8yf7DlgxlHmG5
iPnAdyWVPSVY7I20a/hkrVcExdGWDTkAsaaT7PkPGmSzk0ZWqJg0iYc7FS1Zkrev+G+p/C2sNRnf
TBBNpKkT5zdTETtL8irYKZuYYnlkOlv2XsUO+w+mH80NSi7Up6fqw8BYeNmKQjvIi/tLd0CKi4rE
h+CkUvMzHxvlqwtbj0iC5z/snMz708ttcRqLmDPbSccJtvVmlhnTI1yfFaYvgcm0q+ikUCzDLjY2
ocGxcrY5t62Sf6BkLSs6Zm9TZKogQZVsBYINCAo8qoScrAVJkRBl8V3jRMtIMz0bkjVVhbXiKc04
oRpJ51hquUG2D3Sz12Z/hH6+xWNOs7vPbcDLs5iK+AxbK8M38Efh7cyEAUguQJoaBXba1fDKxwg1
0uGe4X5ydlJXXPuzityR0bkGgDIx9OmS9cBdIo1HCPBG8fzWpCUMSV8+6Pf3y7X7XMwcF6x0544J
VH1UbggAPSVn5O1JPPgtwN10sGgqGFZdF0EebsVBStb7WYXVmfAXWNhh4VDRyOfWv8C+AQX9jfBA
AyIItpwPnDd+WfpP4XjWZfcf7ikY7C0maG33ga0w3Ff/ih1d39jerz0xX1Oei7R9jPWQyBREdXNo
50zQ/gZ706qeF5VJrtqyhHOWH6JNl2YCd6wTu5KyFpj89DzsYw2nB+a6ahGQbItp4N2mR34RmtW1
PmeTsI5dchZyZ7/ech+aKVnux4ed4taPr5ZfRLTCqTvLPKrVOESrCvzD44f6hX5bO/LM0dHKnVXf
yIQBTpxNDmItq86vWjIWNn5a/O/gXfJ8V59d4cnsq1wIouOv+uYoumsS+mPFI4T8YkLegO+8kH+U
oOS/w42rxWZeFSKUGJ/3IRgDneSjoNaTednJFJr4J0EsrBKlqaJZze99NEXSE0M63UqWLNfw9AJ7
AyJBvcpognmIyfHsXZspGzieTHSTFnL7cRIjtn+SfBOxpFzGs3vdjV5hJbpNLJcIe0U9HGIOzjGc
ZW5P+YkX8fMIqqT5KcBySpVbripVYILPqY6LE0KUQ+vjXiNUoxipVPdJnnDY2wPGTKKhyFFknpjL
1DHZBDi3qdDE2U0TSFMZAMb7m31L2WRjEmXVjCD6jwFc4gey59GASp8/p6OE43+0PFhPOYBBve0K
zBPwJCXevn+jK/shZG1jI0b2CgnFtlRzzsL49QWlc9pGQSLZ9TzcMBRhS1RFmpp3NJpem/xSOElC
rfDsmU5DIFstAeZuFBe1XXNYWWRiQwYukovw2bqOI7HVMmfEbUzxFO6lOVhVh1DG+ksqmQnVZhNt
Vk/wmLNhhprbdzrN3OuQ4M52s0hbVmaRhBbh7ud7s6nMbQ1rFsyNy3D0vZQZxU1fYmDN4pqo5Sct
xwc+jRZDU64WS875122IfXecYwKuAgj5FwezAWD00qJULxDRA8ONWjABFnPwQ97JFOdsselfJjdd
PYgWQvF678ZHITvucOKr/9HtT1knXSfAlxHuenq7lNY2obLblbarEAyKyY2248YbpNjkx7pv7ApE
70ezQVZNGKb2/NrGN+tJgL0oIt//c57U2cPBhXrenqxzPYy/rSqJPEhIiOMcafxZERh2e9RvF4KG
ljBKgrHKkoDNH7jVHlWIhAdVQdoG2/D9L7SQ/qNCRLg8oyFU2TWxhrTyI2GNnsfxSNC87vGfh5XQ
5uJ4C9PPjnOgIn5RLLu8ajKogNotK6i9gA9hdEIIfmUvbrp0UgcjH4p+usvGlj2NclyehrFh3jyg
cJjuIS/pd2GwCpu8BclZxBUE0UuzFDKzp8IlusJr6mUcEEQrzq3U8Ff25tUedqODe0BND2NyNKtJ
i88YcqdwNb5pOypHQoFchjvJiLBaHCztDnI5TVRyw7Ih02hPixEtqs9fhI8OEW0eWh+tiLoSVPOh
WCijIHfzkakDa2ZCo0c2KCWyfinrauN4Ymo6N/er00MonH6jqmm0quwV9NXmgt+giqw1IVwtxcJd
L7vgbaKFegyz44elTwARG9zRQIlifceQjaMEEUsnR4kxyLvvt76XIyNrypnUPqe0HaIB0BgGyDd5
DDDxr1acGsO07z0i0CYarf+07RZpOXUFx0X3pFZE5c6TSVmtU4Th0Jg7vadUM2j0ZvUEgktNcNxK
J3yJWtgjkjxSscfWvAtVX6Wjlo+1IDRPWjcCbBLPvo1+S9yR5gu3pXqR5zlGbJVp+rjOZkDDg7/y
BnEXMclI/XKx1OWvR3yGiHz5vNCiIRy/5UozpvN+YKSD2nbls2q9w43OQLOr0bB9M/anhvpY1rUQ
sh8xi59Wzg2x3jCCffLoYUbKu+iGSkdMS2ib+Zaa909KIk83tt+osnNpWK9vdqj+70eWpTko95JT
soy9IjdbbIzUgobdiFmOIx+RVbSTvgBTADS4QzhGyKkENa/56z8SuXb+ohvEI5K+orqptjDfN3MD
QQ4rFJLZ7KcI2PWechbeJlRpAEXxsgKXNg/kJ2aCCKqWAFavHvNLBBcrbHmU3kfqXnBDxjYWdni8
1WQ8gDRO0XAHMftUV+OE2gSSVuDqdCovigFAHOB6CdZ15wWaasL/RGi/FCQk0+HbHwehj6Uxf1t/
mZrD0m1VfLsWlAWiPIiHxxFb8KrKGf4e5e5hA4PDeHprRg3hszJdzBe6szPZontY1ajA0MQE4OK3
F21Ute5fC6ahDjWzp1fDpyyMuN2Lzl2uij8b5TIL6c1G4GMxUta6r1bBp5Ze7mQiskENAc1iu+VT
VIhd8uA6Bt7e0Owp1D6iMJPPZf2TggyOw9Y5Z35ZcmqqqUchHodzGC0VwuG0pYIOYxz+srz9lmiA
RLr6UcxZ/AAP3lwMn6+pJrbOqBMejS1TDCYJdYf3PvqOQZ1hLdHuLe1O7gyvZGaK+6KghXljZPFb
IkpdchTaC/2GM7rYk/5KpG8t3skkc2XC5U7srY5iZTb8DGY/E/FASl7f5ZE7i+n/4bYkbPF/YceR
p8P2TkwG3or8FLboQAFTBDTG90AUpLqw73aW2mJOKn/Cqc0SFUrlz2mO7r0pnAtpioAPYkd0U3DR
2G1KI2WhUyGIR8ptWj/xmRQMJ4WqaJaSCKd7RaJZDRiQA0ewsQ3h1Sq7JiGEjIMv9xtlE52cszPu
qMrNBLrSCXDd9ZfaBKNKMnWie3ZHnSO+03GfhAgmvwbZCvDPtSTWvshfhuBb9pfqjZoC6lzunq8g
RwCQsgcgF3LGnjymSJb//N6q/coLOLMnW4oPuVhRoWFKd6kf4KnPE1YGWeBs3exPElpynDXCFUOq
JO2U/Qu2wP8lAFTF1aWWV+T/MbfrQ/CJVFW7ra9+LXRrrxu6cZgzVN/2+sk/kE/RZY+FSI4NSduL
eF9epDitd7tQ0DwBFmAQGKp3m/p4niuCGV/QUUmOwPNgpK1hJxxse3WRf7QSER40/FHwmU1A7hfJ
irxkGI0cQlxXRe4u04ttXoMgkZ7w2qnx6Ww6VqfcFRimi1ME3mdypaeKStK0qK7qBAp7RMKqy8dA
cOko1cITWZjJGYhZGexs9yvia9BeuA6/R1WOQUGKXj/obn29UB20ZHup4iJvopIPAnXkR1aMbOQg
Um2h6xFlfAIBRoU9V+6htCsLFovricR3O9NR3AusskUUg3l5n51Xf/T5FSx3FVpsjl+QNO7KFghk
W6+TNDoTPAnEXcRcvXUNGzfgntpT+pKeydXKhAeGMjVhGq9I+qBDo7MbJjtQEof3fkjfHdnHjYOK
uqFQq1L53QvHLf5vbGC304q11P0+VXrICB5nOMgNZhuXHN7VU8b6ez8TuvEcIANgruwjBxIvyETo
T/lrs+fyDk54iDGjci1z2r9M3dLZNp+xffUdQXGZOmxVeVinz/oYrcovD9bvtkgkNFr9UhaqZv/i
N2nNmSgo30rSfAvjceIJ6tRLY/y4DF8+97LUFPJ0In7+vBX3PQ5Z9fivp1msIKbDkYrVuFcyVm/U
82K0ZKuQGJ5QtyOVPPAjDOoXuDUqZa3ngnnnDWPfrbD+JnDC8EHNZ///wMJ3+hbg20Lke+GIxyYb
mwzbsXQoHLzla137FbQN0cVOSzJMB9AtTjjlf4xhrBhgbg6GAoX5BafNEzJGd6XJX5Y5qfy6x+Dh
z7uZYTRyaLTZlf3/vD64DyLL9LqnCQM4KdOeKm7wwfmWolSQ8aOdEILqgv0VboTH8gVV2ccueN4q
pPFV228hJLVYv9jSm1pMivon6c789iMI8zOBxDrUmu2li8eaUWOmrRymgu/9bzj+GMGlR9g+xkvV
FiyfjhcbaC7VECA/wp8/hmQwIC9nkhu5Jhjga4y1Sy2jOHB3Z4L35cOMSzdLcoBZsl2X0a0WxGgW
oAT4n8OltmnD8dzOKU5J2CtOwE9RpxEcyKaHOA+YA2o+qv9tX33wVfJAij4RlmF9j4oqyFup89qR
J58OXXzasJcqQ9XckDkgPWBZrhOocIb0iEX5BJlzgmjWPyxVbUGXOwEdasWO586EO2kYXM+U+TOR
gp+rEBnmL79L+51RP93pJUqXBLgarBkCpmHWo4TmpUrDf+bKMLoqYZ9wj7k3pDWeG6qGiE3bQaS5
Qo14shTt4K/OybNjDRZzPmU0kecoCrjooQkLJoQ/4HG9WuEM+NMb2t+73ndoIsXZjQoUp/vjjt0O
clZR81NSLKTutEjBOT4Em5aDxTBmyaV3BlUCzHWYJdFBLrVdkfFdpMx9uGIbpiUfo6dU2WcWMMgd
MtzYtzkmqT1B0sQXbLpsk7J/oI0SZ2LZFw1fPqsUDFZPAextccBxOUawXw7LTbqOf9zXn5wpItqO
LXb9u7OrbUItme6mVObjNGr3O3sPsTI9MKDaOG5/zJQf+w+xW10NwyYFo3H39af+VNf7oEmOZDWs
SQJB3GB1Za37nNpJhMJadF17WT+UCkFyUAFT9TVB003y9A6ubWKG5j0viWs6THKevgO1CJYJEl3i
iPnafPAldzyohhKc/W8vet/bkMvXG0k9zIclrV27+rUkF0XqhNP95rsNdii3PbtQg4k6ze2EAQW7
H+KZHLrH3OGUQt4DmJokUq9dQwjojUG66xsj9Drgz2i+QBCqZ5ZXTCRaMQX6200HDnR4N5lhIgz9
MfFH0kA6c9mqYYeTdlncL5Xf4JcJF+D0hYr+2KYMkZkxjcyD3A6ijLgIFgd7oY+olUSLGGUC2lgU
tLK9M8SxnkAEjtHunq1C34hUOkvShv1wmrDAyG7uk+sMIj3HkRluXcTdrX5uNZaTnLGvJ+8u5HEe
ROlsk2i9+qp3FpAeoUevpJP3gSQT8Qg8ZNFLK0daF4sPbfvkZijKOZpkKk5aAuUWrNXSqE9UEGTk
AOsUVk31lp3y8VDjLnTugzLTElw4nTAQc//8Nk6M1u54CqelMBdCFuj2XcBssv0AVto3nVMW933d
pefLlyaPh4prNACRikr6O2nnHRqKLtuLhJ2HRGYit3u3hzGyu1WBoOlBnOKUqRY91sVgIFPkHgn6
xrRs44W7xgEBKI7ELRSYVDP5MupInoCrYXgQ45qpF2GDx8JpcYHQXJLSDWYPrI28E/sS+6qHKQa6
KCl+EE4ICWlkJwy1fKLn8lOOhXH28V4OjiXORz50jro9CatFurHOwtc4xRQi50xiInRSwjpcWMAR
ld7gL+KO3ZPjRyu43sUa2Fzb2PpKUwLruW+KocL+1qh5HLQqlbayAivKt87EMLRRchR4xwm3ShFP
Gt+lw68aGmFoNKs1hFitwL6Y8xgLsFqNzNcUhIWr7Na1W14Sc53Xx7mWJIccG7wP8NHVP8jiUZrq
wfQBGUUOu/pc1PyNqHJMGZhTcLEYGUQO6eaFQTpiz6Pd5v5MYSuP57ji1LQO01jHtk9N4NREzDCP
mtRJ6UVxYBdL3Av3He07x8STAlWEUaqUlLw9caY+a7HTXTR3aLvZIid/IaQeCA2ACTE7908lf0Ge
x0bOhIK/m3SYkg2PMrDccxqvw+p33rGbW3VqWqips80eh8XiVShQzzQ1UukQIaWH76WfsQ7S4rwS
/ocMjZ/kes+1okFSX7xdH+0bNlDSB/Bh2mnJqONZjYjYrWdAfGNBCLpJv0Idki6nZzM+GYK/rPNk
qcfuINOG9OSh7SaheT91fJkNYCpcZ90UQBGRWeJj6lPh/Zz5kXYBQV+XBuS+FmqvYu3VbXpcyBAU
KEihKN8ZLDniwAYCf+wTKA+obL5rBAeuK8xj7XgJcqf1MX48rvDFam+EHGq2aQfxSkEnYw2fkL9o
T/D5joUJgd0tPEXYwgnJmoi7GM6wC0b6fYXKbVJL9/glZglJ171ruFtDkshlTH7JZpmDWHUee+fS
UOaWpu6s3bBIpBT5U32ZriRPImCZs3LiotgxbNu+X6CuW8EavbWe+dY+W89LktnwGlNkvTOLhm11
XuufAe1KPgDYKJL00x+Z/aPxAiZlysg+Pu3ktg/wxh6hAV56CR8RMC2C9DSaVASQb7JwsyADIbKs
CW+Qc4AoMVV46/T4XLYag1DgMZpiqlJJ/sCQVIbQ3z9A5mRPyTDjkmmBxq2CX4HVGfsPUWx62EC5
zHT2/l6rAhFnv4egsLPupGFY/JtTcPJ+8p6Yw95WewXoJV+8ZERdSfOiMD3uLeUEFgwOe4Q8RLDK
dp2+hVImO6kzsXHJNF3JI7f03LCqnCG8wnoK67ONlTq2StBdsl9DcSQWO5POp5nQ6cUm/WaZTU+B
RYijxtHFQtRxv3hL9IRK2DUet3vGRWCQTVk67AJYfrRVrGCgS8/dzvXtwY2UjiHmD9ADkwSLFkVO
O3zES5OU6DUOGSczGP3WxM6vzCqeSTacPFRiBfXbZ0R50w8VcHDwp1FsyIdyNRfRx1v452jwY9AN
A4sDdXTWPkr9RoRPjtIE6nW/NljDunQtLz8DVl55c5cZyuvEI+P5RvATb/V8YaApoc7YPLJJdK6N
5DJR/4J/EFvXw98356wywS+id5DdpCRk2mAw5VxcKnIJaKuQDGewPYDdm2h1AV6qQ1PnooAnVqnE
PZFrnkTRnbfMesx4ZHE//bVuMu8QkO5XoEq/nlFe5Ly/jfTQ2ENGzaRpBatWKGqZsELMnn1egtTR
bEsLXpxj5+weI3cH1bMG+YYFrbJ7JBOXL7uUEESO5uDXBcn4hgQB6pnLxTidnHsqUEYI2+j+h6M6
C4Jak+IpMFJdhbrStvnSzKaRqCjLIH8vMWXxIdbqT9eOskFXYU0uzv6yavcATgUr9as0UENpmkCF
1epQKEc18PyObfigWzTy3t+w7Fo0aNV3DGlO0g/lXV6pnkojSiCUgvs2uDKx17vTmVkLsWWVp+sU
d1Mo8zouCGR0FCkTrx4k1ZC35NemrL4Q8soN3EcJ9BNVE96gK1X1R6iEvS8saD6leG/NtCI/Rbyy
2iyWLlR5lndNY6iHWhb4t9ubtsPnFyanx5Cvad1lGkHkUalfL34sAEUbuEMQwAxjLo/egARpfTDh
50I33Ck5OlMuOPEjCZKbwHNbSSuDYdkasFBb/z06yygs5eY+Z5M2Uka9HpoolP+93+vxeaopC9mC
r0P33cxMJC86nL8KvTzXB28rIfr5mJc2yDY1Xq0xqOrQbUsRNuH7HxgvVTkb6PT6QLXdTzzaSGsw
6t/MP5ROEUEAnzFnIeCHuhP6J+gARhYRrn2JnAznRbY2nnnUO2yc4mQsv+PM6ZtViC4cmBn+FoQr
NnYk+K/TWKOBf1OF6NSZXimIpz5DRmx0uZBX8pHaJKdUN1bEB3vX8zfn5DPy6N8/R/ls1/BWmesy
zjef7fkE+SkntU4wvW3q22GFxCwsYJbUbMLMIEdLrcxBzT3ZpZzc1yS8zBgKWcT75faDlKwqyoqM
0TJDJZ+TfHvRPtoRbfUFkmXl3RG0xjh6bmemrQopsPK1U/9HQ86pA3GYtzCqWMybxnnzurCfH41o
CN8QaVYJaCKALbHk4ynnRhwj+qB3MhuAgm9hJvo+tIKLS1mZTPnN5NoBcC7UhTyb/02LoPt7+nc5
K5nSCxMHpnwHYIozDDX2oB5XkoRFADIEyA1qD57PwpYcW3Gc+DYmItJnShridSyyjQxc14wVAter
Z9X9sWdnwicCRAGomlQ6RLYVZbhovv0D/mD02NjAy6KQyaCXLhaSuiLyY39TLSW8plLzc/9GSp8/
0Bt8HuRet9AszarO8T9sGjdpiOrYmgS39xV0ENCjnpE+tn307eNnJvcdsUqwI7E+EAAFwjqVLnZ8
EXZZehR1AECraFDfUEgk7HVY/PjE9Y2Kh8Lxgi2jVzqVFh5q9gJ5womdUOih19W5/umGrfcXCeoW
N6m+AUCLmmmaJXatWUUnqKwPOYAq+mL/zCV2/nHF28vPprgYk7um+EED+Kkul3kEbfUtkcM4w6n2
jyzALrT5kATWBHaj7ie+saW/6l6o7pd0vG9pzruJYc7fPtu+ZXgf2FQgqJ1HpTwyLQOEANcyE8df
32c07mmL5ox6N5baElU2Y5+tPWn3ZmwYfODUVYYxn021opWzJyT6eIxxB9T6fZ12vp7H1qfYDMSW
Rdep8JClUq+sTySFXmbBlBNRn6qNM2laFrQdv9YtHtGVXRoW1PbcH4ROHbS77tjwvW9jJMpkvb+H
J8twZftTpzqhZcq9y4xkt/1YzxO11WYrtB6Hs9I1z2wVAWNJQ9ZaLuNg4aJjpdixWkHPKPY8riEz
WYya6rMuqCOf/3emqcdta5+/lU2nfNK93UCNalJZ8yUfCKtrKLkyMyP3n5xKHzl+wmoF3iIPSnDd
t+fxXqPuFSDFxXmL8Ba9EPg8F0um7es7oOWzC5135F3wRPhTltbh+XknaXLNai5dUvRLKs1sHJEB
k1QLcm6UOmsVrD33L0AWaWapL05HZu2OcfZr/YbzVec2rio9/uSlrTwEEES9z1QcYRmfQkAu7Y3o
/swFKdDk11/f8Nt7ILt5kpwwmHSA6a/NNuqCUCsUuHCc7jvMk6Bs74GupLHWeNc5YU2P11/+xW5a
5sG6XAPaEL22rtuDvV4sOOQVqpXLV0rIQ7iXxCsAiP+ONdkjDAtFyoC6ARXMp2U2UO2omc3LdKt3
ksMD7mIEOGSjc2rv3rtcEuO4nT1t7X5bU11B2GH5Sjxdx9GXTqRDt6aQXwW0ztRogHzwJYXEXgqP
TmDIPJ27V1qonRQEO6h5qW64WdKOSpN4sUAgOzmOH7kTIhwv4rYe3xGa6skhHmQdvYztvh5w7LEP
lN1LvoGm5Q2IJfvuUZALeuzpG+LMpiepRfIAmr71K7LxmzDnPqX6Ojo/eRYWXyX8HVTgImGrd0dg
8ODoS4JW1/TEkAkxL95EwF57mwPgYpviB4pHuVLtlBIPAp/qoAq011ZEzEuX/tDP63zmYKCpevKg
s6/+cPajjyzn8RBjuNqTn3Tbedo8JCR+Xzh2AvEiJ+TErFaQ7Qt4AcxamDa0RlKdrxRBxBwdJJo3
0M3wTcLhaRAKWaw9whKQHXXQ59tbM4Z372Ft3/MoHbx432oPNSGWzDVrUBk8UM5aOcDsN0r4jifs
raR2E8kGh1f/A7KK6QjI8nZ0jz1RMLp1nCfL16QIvc3jqysaitneKC2+du1G0DiYNMO1eiRTHumX
+3cOid+uzYzUH9P0xllN6QhSZR4MpfUlmddtmN6sWltNdTElH1bbnn9npkNYrzhiKdfBId9QKa7U
BsxV8hJPCm5kwRZ8OgZK7As1F0IdFSdU19TH1+NXsg5CEJsQprlHGugAvZPWrSWAZDlFaZPjG92u
o2YkvXSp41TjvSO1+/czczY7BjgwPraH0O8RW5Gmury1Vh+LQnb5KR5kPQ9iM4ZaZFjpYnB8MzZk
C/6yejZH4XZ1p49S6zIwlHXDP1+WW47Txxp79r/IAdTJb0FRbSsiwO63nzmuMsBSkrczHWnfdBAr
/edqustyaj+kdYolpNi+i7xcuvdU3dQTKkzoR764nkSa0pL9GraMqD90bOgACRfTia3mCZmSMivC
t2hqf9CEUkuldhH1Q/ba4Heb258XjVjNMCsV36uE7laR020mvRSOgmBL4p0HjFfvqGCz3sAUSaoX
a0iimaR6E3kA/MB3tG81xb3UfGbl3P6m9V24WmLSww0ncecrkfxe1/+ZdWgkWPg8MEBLukH1HR8w
e/fct2Ss+dKd0xs+xVfDKF5gNGsX3HEIde6TcNGO1vISqIc/7wOMwqUyM7XRZiFeOIodBHMwsha9
97mcdnElxv3Dpg0d6OuxqocQxEzBAmpGgeLZ53QJD9w6HXhuU5lqE3GzFcef7vha7N4DwV+Njq9T
FcotxGKZbyKyrLWBi5bGotB+HgVx20Yph9xoORew7A2v5XfRjFSm7pmefvZbCXaltGrGa7gKLxEV
mDUoKjITcKylSeFIftRF4weAmYRnyflGNWMJGoGPVGFchZ25n90eQnTPZMX+6moWxHKrYgwueeLr
m+gJQdBVAmTGGkbAuelWlfJqFOWP+EwMMmzRIl8Eg3sl0SlKFbYxvoyq3FiaAnTvoQQSCQlWDdbh
EIAV10bv85XaJMsmLjudA0d43YyG8s0eQ6yvyi9a6eo/AlJ6Afz3JA8k72tENdVedCb1WEp7MYVE
XPw/M4lJfDncZy7AzOmtXQsQ5LudESJEyhJMZLEunvRpzqAodYu7YaVK9EwIhjOavA+2RIOuNX0+
ZP0ePcoS1NA/3G1VKyzehlPpCxFjax6Sm85uUJmgPFvapJtBnAotqY1XB8+LKwZTgi3zUUDXiaaV
aMwc4l1+89HS6iJTIR9yPWG3JhGoyT6FalNF4uplQlmg6TPnkDi4kkBhkwvUV1uMCe4RGq0GWcHq
VEt/6FHEqfyCi5Oc2hPGlptVhUH20X/1OhWJHZmzBWiqONCH189A1p+CgFdPBw3fuaH6Ax9828gO
ElLyy6uCke8UTk+Ec17yPXGqV++keCfdA7xHVdHzP5LXrwlMG1OCq0Nudni5hqH5kC8viLDtN3Zt
TwP5S8cHfJtYnnsNArWbeqSk4AG6dAI8+ixRv7puNvtvhOpQBbZDfwa1x4IV908+WscXIm1Ik9i/
aYgo9K+UshXqg6DiJYuDf6N0sBSd2MiFRUtBcXqMTSM6YCuc84MCYo5Xwq5PGTfbflTUtqK3kIzI
wXNthSQdsZUylCGwJ/ZDn06zlEBohDghiCwuGKNLJ2KiJGA1jNOh/gj1CSwlnRv8gKHQntLXXjeq
9/VOJSwUusg4dCeJU87vqJ/ayvDSz2xyPYYLQ8IRjVIRKStUb1KWccWDBs322nDqFyl4zPEM3yhb
VV1ePqn4qMIHz+bJGT7PXAy4xok81e4Ghwxyy/hYWSTsq+v7Ebj5kTxYnknFpkxjdR0/xNwWNtdY
YSPl8ga+oB2btBbJoSt14WYDnfp3GAl9ocHtTUeECKB3+bvPInRuEgg+eWdC6rtp+Ytqy7hUSrd4
e+gj/rNWrzJIkoo1gfuCNTfCYHp3YDuh1XmdUJc0l0cm7RaBcKiPhYKiWLrtR0W7xV0ZniYyCnlC
1dLKNSE6/4yEVKwp/lf0v9we2CvuqWL5HEKwFsBAF4j540BnchNAX5dY33hi/WPjGPBsQxNnS3qw
8hJ6Xefv9M1WhLwnKcec3ztO5OOdYu6GCzOtZHfzuSbGnP1u2MjsAfezctdYskewtiSN7La7YOST
0XryaDfLLmfupH+L4IwHhDDVfiHsqr9mhF2/+M9W7GGNSeR6+72X90wehy7xZjaDjXihK95LfwfC
kKZXu70dC6uagKhjG+PRy/4vPONYrYuSJ92U8ImD6BQo8h3PRmcG1V/9KOsnYZ9EaKJQRkEnmDx+
suHvRMpkV6oRmeyrODtvJma7hUJcps5cutiEn6+IQQvU4askTiRb1J2ckeM27ymNDAM816GEC2VH
Hwd22FuyK9xt/OqdgzkmVzJ763qlHWYmvou68OH6iOok6o51Gi9ApGurMVbUTzj4x71VhM2c/qbv
MyAw8fllDO6bjRLsDmuTWMKwwqCkCkFrrVUTyKCpR5PFAlQ3Bla2dn5sPLlEuV9p94szETGeIhAl
UoFlOar/gP+pIFYINuQuKiEd2XwRsCr93I8+MuKJ5UAKS5/aPqLHNcD3KwWSOXb001+nt/0uAzyE
FDz/CahsYH/XXYe0QY4Y0P40uANdD8theec/TLeJNShCeoOT2ZCWXIAfDXLkW87StWM2a8r4PtEB
57QN5vPvIXbx5Ih6pzl2citm5I3uZBGm7+qrc71NBD1JaLeDKPqTxoQmu0ikVPZ2Khexc/XjYJYF
NTkzmx44Jz1+bpKfik63fv8bIT5ze7BeYsDZ1WEBQVAA5Q3TgEhsaw9Oii9r5sEuifB21snMLnnJ
INrG3xCqgGN+C5qEfqxnbXaPwJ5PzwZQbThSMqQRIbRsTHSVmt9K/goy2ilNwZHhWHObyN3/bcpf
FW/AA+QDvPCrcO/Au2OR6RqzsgFPPPlnsMAQAXlnnTUNnW1dBpNcOw462hyK7aG3G33G5Yk+tYTN
IdXj7nlcnI2KfTNQiM05A+AthZyQWU1q2luKyggLzvQZkyOJPdLSkcRi0w6JywrEvejaQWnAmQC0
ETEe8KFIUzTm1Q2qcloAMPnLVlUhhZSBZD4eBWu20V2j4lUx6JnQ3bNGdLkP4UmGIRkuDnmxDyea
7hcCohObDv19CbAuPFBFRb8uxX7Drj2xBjbnT8B9QQZdKZT1efqYPxqhmbsNYqLh205ruDqg1pps
tkj7qqLxs4tq/h0E1GEqLylU97+irTPVYaokCKOKx6n3XspDQVKan4HwDaBel7iC0TdIXJOVGSxu
fDD7ZkNQliKXns/Y3dSnRMGY7S6ESu2UFt4LRFTCVOvzkA716Tuikc8EmYcvjlDHh1OFqDbDBcl2
cCLCN019Na+AOMQPz56f4MOeuKqUDytMQKexhGO/1AFM43V5jAQBgIM/7w1DJNmLCi84dUvjq+8W
q0C0jx0Ke3IaFQAqSQXRWdP37ZiRLtqx1kbfhM7rXh9redQJvwiujKXpmJJpMqhW0z9SsqRmQQxs
iaqwypA1v3fdz60D/tG14fyRI8KgM+i2UruL9lgG/F1vaK3IW8wBxRcozO/eH9+0hrMfQOwjG9HV
//rm1Vhm+3CPpOic5KH5MhUjcqsN5I526CMTu2NW8DXQpvMX9LBmT3+Bx8KMXe7SNBojmwykJPe4
iXQImlacQIr8CcgJAKTihdY6inDnGoyYGGDWQU7PabJquiqYT4aA8Qb44+N2Kcg96O8tIVsa+NBZ
UupUCkhTIOhGEXnrmNlINZVFCgpSkjs1UZmo0ZT1gB+37SvpWSAGqBC44a86BTaHY8DUDPjdNxNF
evWsITKwwl6QRY2PABSEl38XHAWWzVENWd26wEIznn6OLx9dxRP4szwiQSZb6OSDjUL6Bj97KUHk
NDuGhqzLNrl1P5w+FvxjDMfB8GJlR3/xJcV1F5WIHve0v891/JEyeqi2iZKvxyEiteyM2M/6XLsq
emkgqiW68iPj2SqgQauKLksV9yRotu2rzMBpGSxA1wqF6MY9RWthYluuEEYZNh7lC65JnaPWk0CG
N7wXKNFmfqQzQzzvCgtraVOtA7k8CzeEe4Lk/l7HEIIsdLR60RgQ+jWDyL0Yux+h5aepu2ZjiVst
g8iLuUL05Ef7fswJhxfA1JdP8cPpMuQq2beiASoc90ZCAGK8E2salIhr3xvCuiOQRNGUff+VoDv9
663OcO0liZpqDf1tVJipTl+F5mmuCuQHqc317nGU+0BUNAQV7GIkX8KHjJQ3huR3TolkisGKK4qF
PR2/jOliuiYOnz8F0habQQSiH+9o4mEwHz5n+pSG0QTO02pihrqyYeq7acmzLc8v1T/XPZO/XXKl
UhRPPZvzmJuRXwbUxdrXwsLQTQlsvLM3Dhk/2zbTpZEmxR0M4dpp4MIWyroz9nzMZpg/Mvz9PHPL
pI868tINX/GYXTn/iCbOte9yI7wmFEMUR1zPIf9SMf/V7H3TEikIN6ob3VDudqhL7sOZuDimX/85
UHdaJBx/oSUIg+4/+3Ypksv7Uef4VsVkhLJhRVTVxeDASOs3esLLrTOkInxYIaRWw/HOQeNdZm0K
A+vN8c/fxPpMcGpcxAz3gIWJRuW+KjNqjvqeZoIpUNvCjQ54Nd+PnDTbGnCJIoKz/a7fXQfhb7e7
rcNSa0lMqZLDvQ6u+Z4r9u+WijdetjHvs/sfLCaJ5xrdt8+5FzbG/SX0oBzd3E5o2LGUEzGl3/QL
yhegrhZu2XETcdutYcq9fs1FlcNJdNRXU2DEDmOPBlbTq2AjO+mPa9XEFoFq7eC/GGhb6Eb6ym5N
lJ9g158PReRIUhrG9UMq8ZXy5kQkL8v0HA6+kcy9b0wOvlsDfETw9lDMvUAx554TtKgL2c9yNwX7
iR0oKVrQK7mAhfyMBb8lmKByvLjtztaaQ9ZLcdwSWIWTIEgS2ppg1WJYofcwjVWZecDW+THS59Du
Z0f1yTadcYjJCUvBNe91lx04EUg5tzSJs73pyqXhloDL/5oaOZ8VC+ymFcuk+MP7C+KLIIJxF5q8
mqlkvGOs02a1K4ShjdhRb1rnL92rnNxiGLgr+qgaKkWODppbsHCPJOhsbVjB/8YoyY+p7EtddrX+
wvLiKDPIUu9/ANCV1E7ReKGqwqWWgp4uKkQIYRPAsEYGCl5RHhq+lTNxfB3obdqBPqjzudTYwn2v
jeE+/oVR8S+B3yd36Qy98wWZopGgITpa4THH3epdaWiqqdQ5w4gQLcM9dwHsP9AXHq9G2EiUG8G6
kdV9M0GBMW/5GNu/h2dhqkEJvSZhp9QmbxGi1esXjal6Fz/8cbyCWCa0nGul3HcDI2V+RXGYWpWt
1jPG6n034QdYqxOzeGzm7EJbyKdTDUjtmGnw7+ZaWZxJUJoJcU41xTjXo1GN4bcSW6eWtvGUqFLd
9rtZyKiGL5WBl+FOfCOuzYvciMj1fktQWe570vDgbUv5yCg1lLADfiJLFO7MOB33QSpFUhhuBnLW
06QtjE56PIfiBqev37SXsawFNqgim1dxAZb9yrRLpJp9LMjwW0zCn2hcTPVzo6YNIrR5D016Qb4x
rGlFPQkps0vNmiN+OSv4lJqpgZAs3P7oCeo5c/M6f5L6lRNgfzhF8BXd7ICrrf2cWWV/H4oton8o
UZItOhztfS6z9VJ1I9loqUP8v3PhJv13yW7Gvfj3Mh6m7mbfUkq8j5BhvLEpSnhwemJOLtfyQife
b4n6qqJt3iMsc9+2nTFK2BJIs4iL4Yb9WS1eOz7394pqCG5CWlq2HQGoXDN8uenh4pH1014Ig+I3
iF0V6hKuc/6YHRpysAvbLhWmr6+Y6K883vQJKaeA7/rWmC7cWDNf8orSZFlNfsmaQl2wtK+bY15J
qYqCUYTB+nZGWcMvVLCLh7H5apaWRCiICjqMurj7d7RTcX02xtqup3PDJwgj91eYqo9KleaRAk4v
rGgbNC/pXQLZbcc1h59fmtypsn1WDxI0gjScHqiz7jFTUheSQ5mkQ7GsNnfBWM5rk7ROeHlDwEAf
zaGBKrTyPpyBqUHSdEPsxw2PlmkNyrH6MlnYq7WaIqeBPW2qTsLfvwB/MAhCMJPDpxd1cgf+tYzt
1v6KQmhUMRLkxaUc56HDF2v2x2R09tG0v93+fwG7Z78D3OxhgQFrOjpMMKrtql+4kJfJjsgarTxC
eDcUnQlOueUGxnUnpQ6Ipvi80iEH+oVBxVFv9H780vt+0Kifkn2d8BIQ6p+jmf+NX/bfoMaHe23Q
ytHg5JD3YJROMel/8kakOtAlfCbavF1DU9/8cY0/HtKEQ8ArLjkBmDU4BWs99kA++5wUM2cvcU0m
ReGzyoWe10IQHkhySHBEqoB9gSFXSeUJNuxhi5Yl+cdr0YH68G/HFLm2TLJAKgv5RLN4+h8RanVO
X22EHx9P74GgnfJMOdL5MvcPjC2RWDzqypvAGLrxY8Kq8zFqA2mhJM4mKlhYcxo7sHQXp6+fVtC4
FEE6gsNWSNCzb2OonuFI8b5pxX9PsaS3YPV3K0IXmHyEkSbMSer9cl+zQAHIS3uq4gXEt/jy1/2i
BRDt+tY1cgkKWIg/QKVwNmN+dTGGIRloWc4eQOdZVqnlKdhaa/7J2QDjxoZtOKhgjIN04QW9HDF5
DfiPKDw65eK9BtxsdyfimlZopXKB07zJfnmfzS5YJFqqM3Oph/h/4QUu1fkgSJeJtHC+F57dgQFq
Oe/7S/pFXPm+oIdX9s5brnHThqhN4s6LHzrFvTKxrMgDPqgazZfr1UtvQcbEn3nG4LI9l/t+cnqF
mXnmNELZuX6eA1inRKl1gk14Umu1elqVXNuebOdHW06cAin6YCW0G8aUBywmGw/WQURDQLPkfNAS
iLY7hsskLwyw3nxm3asaVWIspcOn7vqBn70Zfy9mNr0cW3pR7CBeZLH5o6vNB/4ZkEWvlRPSNLj3
iFljWB6LNDaMTRQYvot6ohrqpPQMAOuaQ7pFDr2Xm/auf8F3CeUm2YgvCa5rOq2KYyA8YcDqxOT/
dsOvmjUadIAuhqh1965A6+wfeuRxzCJJDR6wZJ1OLmnMUjttl/NAq+eWaNF1jt159+lef/SCASqz
1MVuJY/WxUKJexiqBRqDtYTBMfZ1841bKHhX8imGwF/hTFaEZzOVVDV8c9N60xyOCtLwd1OqYEtH
ttW+JIMIkm8Adf4MTmuYfksigZQkOC7joMVUrRS3ke0EKm58R2HbYlZJ8q5EQTrv0+BUrVB0gRrQ
KT0OZJaD4sEb4lvUbdpvYy5zTFuFpQ+ZPKKLsmOh/G1WTfE9tL4nH6ccWaA48SrVo80KbZuHdQQg
UjedS/+MN9pFkOL/p1ektOme7q0iWn+ndGOF+t6Qv2c7PIes7oHja4Waai1mVtIq3QR3/M1mOE/h
c07SjY1YVLKvP4U1l2Fx17v4VAXcAcNXKECcQI0qaA6UNZ2Vxu5RL3W12PwosRfVDeIrmnCATwrc
XHBfnjSZsTfIRuAorTjQHy6Zw7abDxjEmCluJ99HVvcP28yg4rdBexPbZrwH8hbHKbDTCwPGgptl
aJUyC0cmw+XvB+OwK5oRl7WP5OnVuF/xk26S0o7V6Im/+XqMF84EPxp6QNSZcbGs9P1nyECLfXC9
8PJIVWT1/gVNmRGroA+xPtonIRW+WQWRZQQQ2etjSXLqXalLselrgRlffntXrMjqHDRNZsTWQrsE
m27Fbj9bliUSScH2OEBqz9DC24f4ljMD7IEfnTIF7dYAhzJuQBjjoZ+JXLgtXzyjdR+AH2dsXoi+
WVhNYoloswCZIy4whAlDeAohvq1xEQY++ylJfo5drMVIFr06bSyyqGWIDx9lT1XFh3IygP2lhpsh
wTR72jrXDxEEkvU7xatCrUnZTQxhfIhTXdFT5IxTYVSYUgOtuyO+l6mCwyQbCWApenVyh54VhvKH
sYRmZ/8VS+hPoROOphuK+noHYCinY25SJgcu6pgYarUsFYjHresimb9qAVUfA465Z1EPzoiSuu89
sWkhpisLgBkoxNgSengO94WUXXj/oJKHZ2Z2KZIgVUHeCOflEGDNvkIGJiH0K8R28XBC/hnW37Jr
fUdcg6EaQ2Gp2Xlrk6KdXzhFy1GI02oHfBIdxiBHFKb9AlTCEP+UQkgyndGjiLynboJJEt024Rfx
L7wUMaEwBCKvWiBUuMVt1Z5cCzfoLm5XVsFldXqgWIBNZ0bI+o4ZH13zNMV1tLGxU5vIIc1tzqMT
4NIgRmZK+YPb2Arvr/K/r9SnwXa3VO/l656YyjT9RLZFQr+SDOltC5YvIlQV02ligoDFiB7DVUo2
anQhwPBWwOE8y4Ars60s0xqjE46feoFS2ffcUwS6JXhXLleUnpYixUe2x8EAQkvLuAziE/UYfPmT
tJ0pilKV4kq5/25BH3E1pAXY/pqvgtCXCvS+b30J5/TfK18agksjEqM4FkzZUTcOTVrxKvBRpM6r
wSN+mLUOKptbTPPuRRytE180XdPZAkmMCM/gq0rZQWLhsoOxrbnmaz+KYY1sIiQr8SzR+eYRz3qC
2uW8w4w/9YV0jLUTu/ec8chSrDr4GTEKyFFK6hLDEgf+7Kd7wQOPZuY38w8Y4o1SRwY3v4pDA6YT
O2DmQa7XQFCh9ah457xxeqEmsifoY6DM5qMWl7IEZWvBtMGDLP7YcdZGqFZr//h+qQkUO056xjpN
zR1zrnqKqnwf/lioNB/I14pd/vWjM03PgEU+g0O+fUzSt83/+kz2RxvDvk8xJzYvBs1tkVLBVJ9j
mPptLNlMDOJuMF28Mt1LG8XnBGrfm3u9N5yz25YE7xat/9BritbZnCv5oATZEqlR6s68EZ6sC+WP
E6vrpqSd+4PcmNaQbJraYiz+VBEitKhLcIVXwRzMYHLHaiGSHdshjwrotMyEwUlaeGnU71c0pw9p
QE/5XYms142XY+8P+FVA3N5mGasIad4oqHIniyQd6HB4xCKXWqaZ36fHMZUph+coD/4i5Cygqrmv
95R8PAVQhQ/ZD4Nu750A0K4beURPREwaTW02QPx/wYqyqHcU8HXboUgXzYiq/oesuxokz+TOTVog
Y+pDw1R1zDyAS5uKoxqF8eVjRpLmOtJfOyYUIXMsoGJo6PNFksFpLUMLQGc+HxNjf3DhY7z+aaHl
kqaPOZSeigHSh7Sl1JHKqS8ZfSkmxb2xTBDstcB++OpZmlT6GcqdOocNxftyEVggdlgGdU1cLKFQ
m2Mr9MrN6CREjffS2VO4AmzGDbnOb5T3mZXyVeKHzVnoCrTxoZcNZko+IhxmRZdtfbxexlqP9VYr
+plM3dLkwojD4nBm+8I4MdP65imMzS3fvk/8bgi5OsPyKnpsXNGOu9alLQj11L6uuJJc2tfxZf5u
jsVp0c4lIwUKznIgn+l70WGAtxLV+NPiQwCHpSMTVJWLXle4f2lBsN59/JdOs9DrqfFtWK7qYvN9
yODVgpl5cFfGISm07Vn/8+lIjQ2phnIelLoEt0X9OK8v1+ezBP+MLav4Ex42NINwzaMPv48DRL3J
46BLPIo2y57mJwYATghLj1mo4Dczd5pBRVTfLvFcVaCnvROOlC4PMmnoZ/B29Tnjhp6gySbVnKUs
+FD619jLqQ5+QBs9cWV0xGvYnHAuzQbgPGpI5BpnY679pGxKGVnTsx3Dv2K9poerwd+lICj1hqyA
eIbg4cqGIgxZIsCvMTKtnk1sTpMP44GMml6dMdatNYvGrb9CAl5oHRKSCUJEV4CjR0H8K0qx+U0h
VOU/6SLEzhVm2Q0mowPQypXepA74HyGjvHIGdGomy/MWWUvM7tmAyoeceI49yZCLo6kDk/3WJELQ
2foqXtj24JIrcWQOmiZZm16AvHXemLFt9ddL45bmUElN20w4prGSWzduAIa9DCHm0f2ZUj+EIHxo
YEhmGPJZijvepI9U0Xv4gL17GSfuVhb1AzCJusTXBg9p0FSKhnerg5BxDJ8jwWzi040K0l3MZ2j5
GMYqslGZOJ+Wmsi07xhaVEowG+C5owfV9Fy4CGYoWiQRQ9bqhalMA3l3Ia09JAb4XLBo9mwrbj5R
/k74PsLd1+GjsEgGYkych2IG+r3Cjo5UFIA9R+t3L95pIe2YI8axGEELRbj0EY0f41e3ydvVLVLF
JUaBNfYaSYO6vWWTMgtEWzNiwkLRxl/nmmRQIEAdZ2BDHEA4wNfrUfI3IzabiuNdL6e4XNJ7u3z9
tvi9RYShsu1FxK9//Xj9eAfCuCY/BKl2XHr/1/BVAd6bpRjs2lG/RO0IasfXhoIuDzLfvm1H36xZ
DYnU72CS36mR31pQD1+ot/4LhbuZQntWqNJ9rVg7sJp8ubdj1p4lhK2wQt3pUAcBx7XHi89jyClW
YvlPjcD9nyYsrL7VE/V3iM6CS/bygt8tAuFh//PFNZmWzfz3VSJMvU3JVQo8fiZsk47BKS9AzrhL
qG3a41rd/GPmMVkb643x7/nCTRib1iE+vfGDGulRf1awJBjafusHvazFQ4SmTKwB0nfP366RLKY8
tlofgtCHX/UqKtP9t98fpSndc5HbrSSTNNV3gYenmXDbAlxMQLmVjmN6IyffGx2fXJLi0hrb5Ydi
Uj+tm77qQOoZw7q14njXNjZjn7mj/uUd3TOAgmjoG3AmZUyAOzuTX8kVFYlC6J5rx6V6L9nXvDRQ
6Mk4JQQi0/ArubzvAqRPqePi+xjNyNLmF2rUDMzQDJm8uZdt0SUN1IIw6+3N770LWLU/vGJllg8b
pXxpONSg7Iz34MLbyfJGiMwosegPcc+8yXBENgb82R/QHKOmR+N1hHDEfpi/xfu+qv6QgpMuXadU
KwS5AT3X9GVszj0gn1XMvpYYcMxhh3tDy6XEc3IZpWwU8uh2l+STl6O4i/sIbhEkq9sdJpPEfkLE
npQvwXyDdo/KJIZ74P4ZOtTgaFxbyiFCRf/cxcegnGzH6FSkoBKsG8W4b77BPV/mJdNEz5VZXrAA
Gmcuidf53KPOFoJD+pdISFVFDsAe7DBJXZ6zPjJSAcgPQAHYFSVRWgRHlvXg2c6h1d6eumME7cFV
PBgbCWWnjYwFaCl34yUMc+BrFFaDfQVO+UoND5cNbYRd9lw1PivmDtqNIiWgHR8JPhwONT3YYMA2
FTjPZ7vvTENaqRafgJvc3jsdtY/GkOGOd2k6+NcuxCvy5dN5saaUOW93TUc40swLxVOl1TltMjwK
wNWDRfqRUnCguIGqC0hLX5kUp2/rs8aYIAoWMdPBawBK6wddmtKQnbAr1fxmVRaznQV9LtVnrnrk
e8XLw6Vw/u1o7v3wxXuu2CRrlnBxm3TV8phJzt5y+iVxutGe/hyR7dTOLikWiC5pwPobict1RAYY
8PryRHTO0PDZJr+OaASTQOkxFP1Dxvi6gIbQl5C8/wFpqiRMLU8OllykFFch5oV80jQ+NjGfSyI7
xsbWfW/WR6jb5K0I4PHaObCXF8XMobz3WxeSR2f6akTeDuhJ0IvbQh4KzWbE61CMA7WtDX8wfZie
UTUsV0oIKp4Hr4fLPD4FFAvo/OpDBlauBtxJ3jWFn94kG4jgSCjDSBS2egAJ+azxDlzACQ53NyYx
Shu91jF2g2Tle1ngEXsT2QaH1QPojt2jYC/p9psTysg/NXkUUMVSE6pooEVOEdYCa599N99to+RG
RFi3mWlvuiV98dFXG59i6996/Z27XAV5hrMKJbGaI7ytklAGAH5UxMd6Fomskt2HQBZYbehU9XA8
Rt0YbR3IwoIXeHGkNNYAb0Uk9/GSdRAbD1RVkjDBrfEfPnGpIA0UnuxYev6lLcQEGxP+ZcVqyP73
WfW3zBXkFEkXazpfRzBysxwCY7n4pjxFGT4DEwR2klBAJ7RpOrBdZLzjAAfx4Fs1DeOMYPTgDdGG
njzaC8wGNQfQunVcBcv7MtDHt5iQGJbSYHk/8a0MQkFXZuwotpCfKcYHeXJ7Wax+ZWcg8rJ8Hu2Z
+Dj7iFFsubKFGXKG3bJVjMeEol2sjK4cmNTQp9EYokMdcPI86zN12rFZmPVyJyAJ86jUfEIFXBlK
q1n16kno0VyT79o2f5Fouf+doKvMZv+pnIXi2U3ewkKSzQmCtA06ouVB5wjWqDcLrmC+gQtBwPaW
pizqqRbA6dIeUf7q/aUuC5HJopYNt81i/gNdu1sfEPIt6JKgFU8+JqAonsMBUxZjGmgN3VOPUcE1
tXh430TrSndXVdEjWSq+q2nue2E/QqYkq+J3qSodTgqOgQOYRXGU0Hg8/ft+cncGYj3Z7lrwifgy
e0j0qxAKwgixoZpPbZ6iSOIghhX7NbwN3/CpIRxtqK/H0fW5dQfZbqgUr7XZj+yYexUZ2OehJ83i
wqVG58B1pC8ZgZyejqvFuq1jZm3JRBEtGuUjGkBQXE4cl93olTfmxhvriRMphaRWyzu3ETQJ/cgQ
w1ADSbsYANXkh6jnZL10+i3iy/8kC3yyYKew3w11nWFgaoWfCGlGBo59S/6L5K2JYk+gj8aBCTWM
tuyJ7li+WBI3Q45gXtBhrOo7xx3UzKLB7X12e4X+4TZ/EkM0vGMdU+5ExylCi/ruAxFLvwwf4jdm
fPL/OFiaF5ajZlGo0CVSWapy17YOEieZLNXwc9pmloagO9DbcsTJPkkhM+L3q6mZRWBZ4iTyWqIt
3eEcppD+XDtSbhsBU0IlUExcnyVD7IALjMopqPayLreafyfNRt2O6nodSTeEGvKBcPfXpHrj1jWq
aGQ+Say3UI/fDvdwKEldNFAPoT3a7WAgfxuCngF5Vx+KnaNU2vCIrK952EDFT0KIK2IA4eROTssX
Vxb59SMSZKYZ8cV7b2JAxStFewUI7n71vyAlqv1ahRJCy5z46iDHU8xq/DDEcnHj/SRZFdCHVYEu
68fgnwPTqF9M47aSk6B92G26Hn+EyqWpKoCAa2U7iuRebGMBh9MGeBCDS1sFJVJjwnSbnhPOnt6Z
mOSg/Y8xNRc5rHzy16VoLThv8IpCbG7v45j2KR70lNEAcx/UX7+Ct7FyXqqyU/P4PSk32WloJcZL
w3CvT+ffiyuV16RBzwPGuzKLZOUacJjO52ac3+rPEYh0jpDus+AkYWf6xdnM6Mo5UJszqI1bGyOE
PSTC3qFMffZfNcO7l5hMleR88+DOANiKjzyMw89OY3svra5A6VoXcGNXyx1zsFRDoiLRcsNRNtBk
8EByWOs4vaiyWGr1hPbfUJyT6A6nZe0uCzUyZNpwtGPcGpfQohYVUm49nYgJ6MKfls/QOFcQkfUu
TsbaO5ACFww2hu0XbqR0WRQsF33ugtJ8iGKc1xlmFB88lSmTWsl+cpF/Ca4+HHmmkh4DMAisPo3c
tb1Xe0GNL2nZml0+6vhfKWb6svq38TNyN3Ll22gVsVAeaLaevhdpUy1fs8is3cz6LWdG6wJMn+Um
FNaCvTEHnEfEiQOcTRHPaRtaS81KSZIHVCFPskYslrpfBxKlRLTY1wjXYYef+7S3knyp9SxkpA3d
DSUyQS5ffIOvr14/IH0ZmIaRL3cEq/xTl1lYy0OX7qCjRDt0bqMlXj3d5PeBPlxzSWZBwg3sDqkw
J0UgBBht13zqHeAY3rOC5jiHowGvehHF7Yntb0Djivb/PxmLAp3n5SNsUO0ioTWu9AaDsXZjLQA3
2kWTP2vtVO6JcwiOGO//hDOTnlvsMUw/NtCEzTqd17DumGwRV2QuyrOANBuXoK9ZAhziQ/HFop8P
aSbOVvqdsrDn/bVacExykkwlkE/8KZHeUUzxHqEjBeUmdiOl2MiFuiyxX8bfY7K2bUL5u80fmH4S
Rs+pO/QukE34u0iAyj91MmY1KTEKXiAKWUNDvFpfj43fXdYwJZFdoSXQxNBR/LQjXHZWTkdd7fuR
OKiz2hIJuKVPyUclOWFAixqYZ9r+sR76ftFlXjQXtJEzsnxjpiIvYB09BdSCxQ+9ASdfB/PlDWSd
Wk6pvRJxSFztS6+7ARfTEtkWJQVrr4njdTYmP45fuICMPb2aQ3MtnoaFzZDM2lBIvSMgyuTkc6iS
/56BOemD5bDh/X8PAnbhPTlH/hpCfFGMQCBKZFt6WfmexsP2Kgwh+9zD2pB+/zhd+5VpTm7dAEGy
/MybidO9pXNI9mPR/frRKUv2jvsy2bgT1TrvWuEglpf1OKVIxD9NcnSpn7nU7j1ewJIJua5sPBpo
FWPF0e6UUoLEp5284iOfnBVGUKldErv+wvYZ4f5ORrzPN7a4XoOfzZT5IadYuRMYyNlFtqIQmtSJ
m7aJGECIaUgEE9qbCZOrBNbAYxyYg/WTNdFsN82SHXwK5GPeqeO0P4i4J3/9xzIiyR2zYND/5QR4
sUULALh6e2e9+jUQ+K4zsFPvym3ci9vFr8MK/U/MQYjsh8hWRLBxy6hTImeqxTURnrKDc77MFeod
oTI9vK0oeLJk762SpMaPXahsugJmYBUbYQ/uuowuTBX4nhaM/EHrPP7BTnTU9H+j7/CVUoLB25w4
YvEeLYRvpAbDDz+3Pd/O7hf8PyXKQ2VFCslkNnp9BEIBXJZP7gTcRyCLsUGGGhY7aC0IPWYertmJ
n0SMb7CDKPFKhtWY9SteTdVQ2vkT9A3N4gZiDsdRJTkwTVcIx36vLyUBr80LRQnOjOEUlzMFmG73
lsOgc4qafMwVawUPNIQvm1tpg7zgw8qZn/tN3NY+D0e36+v14Sv4xTMN14DAJSYddxFdFPrtB3To
nMjcweTEFxBrDgOiZ9wCF5ipU3q7aLmA8mJwAezMqSpJH46bXU+pZEGNJNZIqB8yNsrnh8AxTk5E
Sj0/XJEXMNSRSW9PTT3RPV0AMRCNgy8x/htCtcXV9hvslqwArgEB1wTHZVa0QWRkI4+3xgdieixL
/XwOuUWmeS9eHayekJpCabXsmagIYLEjffBaEVXIUmf0lyj+n9NMbyxEAkUTMRhcGtzIKICjTRKu
ztHMgKSkNTXS7voc2PuJzcLVpIG8R2Lw2Rf9MNqpGLYFWvRQyUybA8vdvAd49ryV40xrXHWAeInF
iS3h79SBaO8ikLDCRd5dCx4FoB3AFlQ5owkY1241EoSadSIgulngPQfu50ky/BfAqR97iGt/+1jD
MGIvyxTTG9WMOACFZcT6zu4drNMumt1uUe1jccXLqM8CCogW7ohpo4cAgw2Z4DcBZ1SIMjbsC91V
a5VRYz0J0mjSIJaV+Xoe1eoPeKKbVlLswO+wSP2Jj63cEtIiIpjmTFQNUrQVvduEHv1ujuoLszYK
4m5fWY33954VsVH0tesQtWTXfuusxx5dAmLQzbEa1o63sWFj2rTDTzuxROUItjJzbZyinaQpAHag
AuvG9x+zxdBRiSgoQPiHhlzpTt/ONYg+EwSRU968qDc5s3Yfe1YJooweKWChs6cMwB/HY/Sn9RAS
e9yMsvPwopu1qbNKYkyyMGuURtipdJgyWPLrhIKXVWSpEKi0Pyq76TPIlPS0+5RoIghEfBsaUBW3
OVYx0Ui+zee5bLiq/evtUvL2fcg9K/ts11x6+dgjzWM7YBWDbNqNwPj4MU0BjtDzQ6VaySo/DJKH
42Jcs3gOC0sOpx1pfD5mjUneAmJa09AjuOI4vGaSZFgRaeA0T0/7di5RxUoqB8rP/VbEBmvFksD0
Ly1NMxKy12D6Mc1x/AUNnkUL8TTkvFlvbQWMJkXpBf8n2mzTH+4k/geJXaAztdYblWa6FDZGbRqu
GgWV4KHZTyxXFe0Elwas+lt5b5uwvVf2osQEpFkcINiQIf1XCaSTw8T2XQQwlCZnQYX9kfdOnDpf
7Zwjf+J02l8q3watU9yCU+1TDR1zjcaddAqIYDsVMS0jveMPfqgm959X47xNYUi9NeDRZaYfHv+D
UEA9gUnfteeMMvgN1po1xAsg8Qs6zoKkbXCiJu1kmXwwuiYqZA7NycOBkW2qSj0CloMTEBdbw4zr
I2/K/nZYLgectUKooZBbLvDyBg65TD7rlGFJef3RbWi2ZWGNCQvisZbiaD+adQ7Sd2nt3A23G+LE
AaFeLyVALpIzpYxQ3tm01VUr3bPzbT6E5tFHvkAgOwUlaOOe2Sg8z2IPWttr7qmFupZ39t0gBw1M
zMP7ZqSmQxaGimneW1qRbWF2d6oRdVyjT9X+GZyq2Acznet8CXKxNkrCdp/N7qiJ5YlGaoSa2qBO
HJVRDphpkMsucwfTTXHMpMZSVLXaWM1sB6lSZ4zjwpj/kas7KhPyDyLdr7ZrJNMSHXmFoTRwr0rh
HkmjXFn5w7tpqZTs5z7CGcLEgyqHlpLb7HAoi9JiOMM99KDJn6ou/W6Yt0Ciceeb3tszrb2LdyQk
o+wv37jzdXLO95r08NDZeMHnirhPBog+1VcMur1jGomJsLyl3Azj99iDo3yGjtBK4rcUXHxol1yo
pxaAfLRooYJhKQZ8nIIVyHt+kuUnkJBMiaA6XirvcMkooFhqiVsxPGV8uWU6OD9yxrMdTUc8SfDn
RXbKzxf1AFZ6p+jdxNIZPerhgVuMD/qEJLZS+B4Oe/3DCKjVESaKlkisHlSwNvfxDiikgqyoda/C
pM0b95cF9gHJHg3Bw/RWHtd3iSx34UTwm/xi6TNmocY72UStROsXMe1QXm4mrHsPNeV0WCY9o10F
yDUUKXFv1jVgvakgi6OeJEdCD5GduC1P45I3lVUMKYh+aietcQ+w0USYqR5roTWyN3h0o9cIBYxR
sxbaeJg2PE8BZ5k4riNLcy/qG8wkbW0QADDQ7QDC5eE4+aVazVI9eNczQvFF630UyQe7bUM47Xzm
+ykx7Zmx6zgaWkM9hNOE5gZK3E4HwJSLk1LznPkyqGmplHKZ8G8mFOw6+MSVC11M+e2Q0syNLcHV
Kqs0xd0lUsA/oXtkyA9x9kxTbMSytY0MvYnpdQPXmABdeRTuta2LpLimR/Ruq8zlQ/5E9IEHDLtn
zUpfTe/1euI6CbiPTkyjfEnXFTe82/+Hair+eXbPPiTlI+zmE1PvOrNZQnkRg5iLpyQhhSxjH5XH
x8nhDvyF/pkOZzJ8S7r9R5SNFFr3MHElaQY7EiXudYc8Z8IQxpIn80L4jcq/mw2RtG8nKGs/C4ph
vRQkyGwVEuWiNcQVHnG5M1AnmPfvtm+UvdmpNFvurGeSEU+jngwNyPWRTfQtI0awKVYqFfO9g3Ef
f1C7FrXc43j8m80EIgIX/JFLllf2BO4wWPdEUO9LJZHoFw1USS1D8T/EmybHc0iwVUe+ZHknWOuT
12IyKJ1cA+IvdO4ePMbg3POvnqfpYWFj9EPJDO0goEf3Q7dmvar0bNfKzkvCYjTElTP2zPQDBmcS
svrt74n6jL0fo1h8wRuk1sHHGmYAN+eHaE95NZ/eX1m95qzI0imb1uobpnoeAaL0DEV106utgJxc
/CIdigPU5ygaaOss22N7kKvrRTremsqvH5+FrkLzk6bBud0P/zEzT/Q5y/mmbBR6b+5MDYNK/MOC
fd0KeLqKrPrG0/Yj+SYgR68PggrCm/qT9wSfRcf4EkMBY/+l1D5/3V8G7eNBbsdhdtAPiJ4xaj2R
5yVrKO3YSSiJNThhIr96A8Fi/AOBjsl6ncEe1apXMzJ63FSUxkjURr4w6S7bfm4B2Jzt7nXnWPGY
q9pr1YtxPCNZA9GItwVNqq3CnnNIHbTLNu7Hb3RNZ3IltqQwrVTRaAHgnhIJMI/iHlEQOLL6/Nft
GonJ1/X6/yqEgRJjD7z9oMGTh0LtHxmkVLxLEUhCaBtVaeYxYrHNJDoCpknJCLL+9SRDuc2FnvoI
v98/oaXMGoZwVfGT6/xELdPKofECvp9QH8hbz1imz2JKDu5t/fSMNMxTXayOwsUzvL1c1jBMjiJh
8thn6tv58LMLnok3XaodV733TTJsr1+sawkMncQsNkhssap+fapCO7RyNibuOf9kBbr4g+rZPmrB
UG1Sahp1hHCeBId14OvTJhuklPC0z8g2nDwEEeN128O1hzL+yHWNt70fKJfQ4gyVj91/jxzewKD3
HzGWGycbdi7QTo4XzNw8etHh6LXniy7VYfGrAfJdhGgjEu8LROVUuscWbIivxuv33sgWFPzm7H56
pm51PfqGAYyYnDU7Tc/XkVe4klDd2IT5MXP0GNXHohfjoH1Th0MzRTyu80+euNCJjS8INQl6wvJ7
kpBhrzigb4GrVB3Rcg73g2MdREwZ/pGftj2H/S1SUsxLFictOdYCRi/sd04ZSnGvJAilhAipqK6O
BR2xjYjGB3SZHN4SRVLpGVM7MAeyd0qTTUgnPFBirsJYnSRyxJN7LewU1VFzitQJzTyaIITasVAQ
iKet7YTujLx/T4xTOSRP9whR2bKqAdmx6VhZ8n63pjSwNLTRG6mZiXH3w0oUkaNHKGAGqr1eRR04
W00J5Ej8vNDQlTZf8ZYQNBETJoHO4j9gACBq/qtBAyfvM4z2UrZnh7sDmhtGQ/4bH5veYwnr9/m0
ko4crRftIkZr9dITm9UYd2eE2CekGRvWd4dAFDEgsN1jekzCH5r/cKlWQByL8QsX2yC6wVmP99wC
kLPvur5z6LD5wB2502y7gU0ZKslL8VcwmjqpK/dqQdPOFtV7aXQhKDij6KJo6svO+lUKivjFG8SS
oDlHdvHaqB70Y0JOPfBJSSnd0swg7Xzp0REvyvyfxwQSMzqB7rU83ItLv4Ct/ecsKHq3MQxnzP82
XNXcT5yA02zGm6UFXA0g1bsF2ogcvcjcqg5qUQ5eAB/BaW+KtuqVgNj/iyPmbCgzN7ROA/T0sST4
YFssVTtTEGCroTC7opGxV+PMHR72ao6jX6DYhDOj4Q5+M4kULjQ99l7Q7iS/rolRyvopUreRzF4X
4pLYvw19ks3OCHQJ7Kkubi41WVqG5dLWlgE1iCAX9SLi+/oCBIQQtFOCeVIpfqXZbFZ+Opp3Ks8o
eHr1gQ1iaZ1M9XfsSR90v/2QzRGYj9hG9BXzqXg4xW44A4+xO4dn7KzcRjESPEhrk7EZgnMG7zPj
qIrTPVvFdfAkeCaOhcGr6hu29FLv1Z0aP+xvdrrLpKELm1pR1X5PlL+fJKezEVzWoygITIbmbLLf
85WO1gTpFKES+fS1wksO0ztHpZY9AI5x7n819D6YUSfIVNsZ1H8yovckJefM8RAp8OBVn1oFmIY2
MA07zEW4PR1Vw5CcNZ2VUMQEzSmCghe1PmNiHM9sDJrySOzRD6got2Vvb/k3RKkXwu0bKO9CaQu8
WXc1qZV5NpCDgNvlgUVvG/l4udnY0rsO+blJlWDP6wNE8xUzhJj2kt5lgzILzRjI4HtPi3K7ivrr
pYMt5G6sKruSNybM9oT7H1tZTB77t0K5Jr0apy9GuIZA7S/J5/GaVX4f9ugrGJ1l07PZ1hHxQUPS
7rMbTlKmjXzC/F8j27DrGarE0Z8MfuJhc/W4ikmvs3lcbhmB+DPPBY8Fh2Sp68IMIu2NBYvbxwLf
H5Rxl87aiNIPAKias1u5MFt81vLUFQwRB8ZGi8bXc/VjP7foN2AjOIZwsHymL6lC8FjOrFgnQ/VF
ElWnfjqTkAxFNrhAnv+GGMApR8lmJlshkNDVt0MSFRxXqIdHc7AOXI6cWykXycn12TUXOdgNeKVT
56+rP9KRuHAlZfYWXrKhMl3RoyaZlqhLDE6GEjagXx6AL2Rek+vA1l393qZxNEol2MLOKzZ8XqUr
L0RmVueLrepXMU6VQ1s1CFdC5PZgBUDDN+26d4Qsthkc6TgruOu7k+rJAAP94uk58jurl8tQzKtu
NMjNvALa5KExILsgQnFgNmM+IrbZKGZ1nDcfHKiCgcg1EOAwouiZ7/tMHEFVhaLsgNOmoOBPQTg2
9NsOxXO8quedY6G1a7ubL9FlGsu9xTCH1a5kE6Ok93Cpw5sSXjVOLwSsc43vRsM9zHQvScMsbscS
y3DXt/J7BgvXl89lzW/WbXs1VXkGmYQp1OGZe2vRUTbUXCXVmJV37wAXJWGuW1wd9JgQErc1Rcra
dIdd/G1PbFAEq3gxN+GsWPVXeVoAqNMC8+lHZCL1ZwzKzxbix21jQ/zb0k2Dn+RCozCY3FacTWvn
V5AckwI5ntUDOYiGKDY65yf4pBSP4FZKPLubyXecRn85sCQIXHSvqNMytTURsfEZ+6jh0+8ORJiU
61YriKUJCnApg0AbtBe1ilEqsRUNmWJcU4cFv3KhKO5TqbSbWenDPlUO9pp924rM1AWHyZrgOFyI
Rlp7wjrytyAOIHVr8Rbq0iegrgcb/nW36r6wTB2Emfz3JfLqfNip+ZL764TABCXtrn1vq2I1xsiN
bHH+9bWkaauWfKu7P6H5P3Kg2NBlm2Yv53YSxQ+BZ+t1n5tSEN6AlyUIH2wkwaeYQ6U4agfEGfx4
vXCXMbXOxTfJbRLFCz8tsIWLIyRr/fs7P0jsnjknXbqf3pOUT2sNOJH7Ykv48aRYZ7i+uFxVKAAG
h+mADB0DcDtyEnmh1uKKkelcK037SWkV5vjfeu3q06cmG9aXLdAw+zPX3W+mabsMP2uce6vFPPdi
vuCeNbZfn6ycQbgh8sjuCUItflmXuwen7Q7S6qYyR0pgcHlIZTwe1SQbaKAENN/YJO6HWjZZWDLS
hB+Se1BfcldfBQ93LLXwaQ45lEuG69wve0B+UexfNpbXi8VzqtE+uegJBBJxQZ7PlXwjNJ1CJprz
m9TrlGz+b+uDEXzTpm48E7NfXjYGcca9hFv+ebwSsozQ/A22UMq/WHgga7dwzMxdvz21Jtt7vn8G
Nfc6c1EfDnMRzXHMNZUE3Oh/zcGAZWGA+6CehTX04+BFMeg6oq4gaOcYofFBgUCb+Or+bkGVG00r
YoupyPiC+QAJQWCuHDX1kHJ4faZW/jo/xPbjAugXiWnVhvdbpzYXmnCif1z954l+5JNUVGKqO2AJ
cI4lpAKnvZA68334fhApWIoaMlHRLb3t8e4RJTmuOBH1B9fGIX0ZyEu1kJQG0tRQAgt6vxqsr7sl
c5ZrtXY4EhFYo/sxoFzeSSs9oORrD3APNcoHlJokrgJqm9R2SZmUFOhtRqjFROyYJ42S4A8uIUtS
Et7inubCmMQKWNVjTYRjc2snRMEZre4QaQWgbkuFuMqs8aD26TljwR1cyeoMk75L5uTOVPx4OffH
fyOBbU8Os3en4unDmhFM71K89PJs97HfXoW07APWf7cvWy4qlV3YvpDxaqYfMwEynRUgJq29+Tc+
NDrXAIhm2l7XWOpv5uXrMPNaRP0Uty90+nUhOEsjdL2PpalX2WvpIMglOkUGuzq+FRe1sEg0PPLl
2Vo1dEd0f7MlFD6VfRq/NY8L+EiUhKmhWHAJKh5mQ8lKbXFTMM2xscxr1loTb537r3kIq6/jeraX
Plx6+J3S2IDDLoD9f0NiTGL1IG9APC6uiWQcrS4CFuLNq+f90FlrpNN+IN0F0QLqUhoB5YxGB6rk
Ru8ufLYDgmSShB+76EvhgkEB0YrzGzxH/y0U9bEbjcyTyswq7l6AFd2liAeLSvy1zr0RGuHfJSWC
F6oYkSVV1mOHoQlTC/bw0lw7mZgJiycBSQ1+yIw0lvza+q2b/rjQBsSxD+VYrmNFyp/Py0aSLdYI
HFDhZ5EVcB0kjeYgyOnwzvfFq1E/mf2PQbFi4mMNTdJfwqTgNmGK/AtGViePXSxn8QXCbrw4F0yL
9/U7TfRoUkzn/1ds7VJzc47TwsE6bYMLLRUOCWWrD7etOjwEyPwcMTefjd+yLxR5iPDQ3Uja5sys
koht85a+/mtgVgtJmaZbq4/pctHggTb5bISClR24jQGvAS4gE6htrKhgtY+XkLuvrRKljOoITQhM
TVpMp2oZ7YxJSydeCCkpM8sDOXX5b/EXVC2rmWG2w9K4OL5jVML/PM7z+W7p5AzIM4V4WrP1b8OQ
exoCiBalw+iQaa+8F+d2qkQrXnmorAuHlARUNnb4LqrTU4SC325SVHvNKPQxngN5H8Tdfb82uzmZ
37JDy73JTYZzoKlRTHORbvexXlVQIMv1lDzJOooiNwA7nbmTIfGDlaNqnVaZMrmRJ0SwydMQs6hm
npJKJHtpIB0kIPOHX9pvQpnXpH6Q//o7yeXTVWy8eGgj2dGhC+PFpCgENHcbixacOqnLV1YKJ/WU
B1nWNfXXLAmmEsVeaAd377pMUQW6pqxQcuAwwcqMBvHhUxMk4wf2/TXPEYp2+o58+Y/36kusahr5
ciP40qI6+QsfWi3VkO9YzGMFfg0w1u8mqGnpwIS8uIoAB+MRJPYfOX0X3QbJg3ddGpatJFgJ+Kp9
b6rwuF8+5U5Hyb5vR24nQs2SollB30vn3HONWp/JZ7IBZbT3ThCyl4zcKUGSmI4RHks3PAx1jm6x
8mGL6hGhxEHuC4aO982CiuHOjLoCiBZUg1G2w0seepTVbXjsVDp9kmQnrxOZjPFR8W2+1v6hpu9Z
XI6N+lh6+E+zg2qtNi2g7jRiTtX8xrSbhbcwwmHqvidSuVQYRBbEykxGDe+suHY0Nxb2fFJm06Wu
9C7fd4ltIgyCi5uqUxgLqZEMKouRpUSgN1zL6kLJEPVHYSblGzhESNp1+QDCBp4RN/VWJN7MJapz
Ly7YFXJHUaX3ddXa5VN6wB0aKn5yAE9GZzoJVgiJX20+UVd66sWfbjFjZRyFDA5Hp38UdEcCkfeW
GIBauoGIrx14jDPz5Kr1bM6RXmGy8BcUiaPCeIMvya7Q+uiMD0WHo0ZvsHxbDlY7FNd5+uIZ4etJ
HsqdxQAolN2HsGZDW9ru4KkWm9p/fsPsIaVlNXBBo0kFfhMC8BjlQePMRCeWe4JN6rMubzcnxN7w
tG4Odn1yrUoG1nMGhA3Hgdl6ct4WCCf9lC5aVWcthse5h3G3c7TO2Ua7kkx7//QrNDrrkbqgqase
6Td060OxETAeODIKz92d6md7n40NDhkrGPuGeddiphL1zo0/rglXZZ+Y0KrtoP6/kducnYvuLM8b
GbvhQ8hJKcA0hFFLixb0PW5/nI9F3TBWJdvTlxpyIehWzmFRzOe4tBffthW+Qtw+yWz4hP6+gT/W
75uB7l5XZrDc6geva8w8pfgZidUDSpZ23eP0o+/rskfRb+2eWZ3Z5i6iyvd5NAv/ST30JW3Jf0UV
rG2tu9dp6b4cx4+TNjCXlm9OJiave9kL6+Khz7EP35A0eEKq4pCwyaTOJmQRYU9rZLJXfIA2zoM4
lrf7Q/EEnkfcLGWd0La9m7EIzKoVzahirg771e7PtsdOa8cw40ENpBh0hxfo31/Ul51/+5wXZNP/
SmwRA+uO8YPzBz37uz1DeO4F+Qj+9tUY1YTbWLzd4/qDHIIcpqpvSsXkmV6ko4PdHZsL7GhZe1pr
EFW5IbhG0ANehX9myHLpqOGPVEnawfgjifrYEle8rs0aAC5LxJ8vbMIDPJiXALMAbMUfaWC+hiDD
s4S0D5f8y2zSpGphL0H55FbDDJvLBOtDrnuJwjyqmy3Ctk7CLDDgpdRiedROKAn9Utpyt+AKFkh9
XAcyNNny1wj7TSmw9YAoA5xoilKx4h1XfFjC1YisVWPNxxh4zT8q3XbduHFsCZd9BqJPvFrAqgbo
lRGVkbH/zxCQ1lp0oYWSsNrEdfMLJk62U6mM+wfx9eOAwcjzcYufGcJCo/1HtoXBZtk/xJIXgBau
B9YAIQ3l8p9zxzS4AFBNp2166w1w4xv2X8SPlDROYINnHTHnqEwerY4fwEBrUTakX1Gxy2UvJ8F9
Irt5hbnjRv2J6IQBJOWskqaoMlf/RB/imKP9vYDKU7MzGN3LOivaSjs8shaLAo4RIIfkesuNhK+O
nCZUSEywhRMH2wsvO83ZjYBm1mrLser02F05VjEz/uOUmKS/Df2I1IcrFDCwCk0aHjHHadJt2H4M
4Qn5122CUu3x78RAZPpMDbK6uGV3547jIBoOU/NQKBt6QeRfgv6J2SuW29kFkjmezTUtIhKx0/u6
zj8gE1CxtmmZ+ZXlf6dQeUcnWiDCyx6B1EQQR3WIiYN6uPU4WL00Apv3XP1LftLCT95c5V/FH8Z7
yqOT+/8LbtIW7Fk0JgJLdHAQLIc72NDCTdSAYmz5PQ/ezYHhZVtRIdV4FUvpHKnXdMsj1LpJ43DL
m7a2kILlpCwFk1Y7tvptdapdZCxeg2RgljAazSN69P/QCV3KukvofLBwAnWJqXZpF3+uuvKTNf+6
TozcN/tZuydXaAz3vzz93KhD48DGgwKHogIKA4f3LJIjb5Su4onD7fGYFeatxL3pzUikvepDN4Jg
8cun6ChkVlYVZlMW0JOrThLvyEumsPMMMJtSg3NgIBKU50FXn3JqTMt7XxU36FvwP8H/KVSrzAks
2Dmze64LYbsjP53B6vdda3t9bSsofPocVrOOcSb6C7qlRFjoymn6xfWxqR/AX962C+2Yy+UHIn5k
O8DxhUBU+3FaYNdGJ79NCVfhbSIz5WyyPkm9b105GhNlDFhvmvWlLM5QqETQNa2MsconJthWgmrk
H27zUGa6VTcEQFoCEFRzl687up3L/0njcYkoJHgJ8n004jOACqNoIq8zFggEjr5V+W9t/yk1vMvJ
qAcO4wlnCW1ldwhfeacq8xtuj0wlQUq26eVI0vPqSXMC4lLJZBWv1MOsrKRG4V8hIJI2irJpdH4c
fw4W3UtTjfadLblQHAld2e8YJF3id1Kmef5OURn+4L2sIVQfhdFZg0OQPzWFlqyadnsM7aPycOF4
Cb+YsL4Mr5yeH0RqtmWP9i4plS1i5uC6pkIyvhSiEZZonNdyFJYCobOKFZliKZaVZgwE5yAMeoJo
2dsJS6G0j2VUZhXEdJZzBi9K3T8WrsvAJjGHbZZj4JZAz8ni7nUZs9R/2KvK45xugp4bFEmsS1Ms
V715Iw3WqiQ6cVW8NzazEm/kywJvgIDo+/IQkQmMpuWoptV6nsWourToRgdM3TJbDHlizkzW/dmN
oqEGu9JKOcH5VIKIZEX3tLLOMGHUGGqHamCYoPxi3voxpH/UR66v/x/SLwrSx+jAsSzAC/cvMgOZ
rYYYTHEwrrd/3lIZHCUaxYhghZxyn/0YucZX3phti9xNbm7Wk8dI35BIe3QOU8jxLNbmabus7zVb
9ccpHZAglYA6p2VoVE+jZDZ7OgBCPfqgm5ougxprj6v8gWHGJNBNSS5YZCLDyaqcsv7p7+QkHm/8
sez17nC/Qyy7OM/hCZ/b675c6j7rNX66P/E9hkAI40C5/FQIlSV6ECPiPQj09lzghP3r+RXqaTpA
wf6DOG7hhnPclkcAKN/MRnA0nGJ23Fbw73BALj5iAKKUJuqv6deEY58rgIZjGwoT3/XKdX+1vDKJ
Nsgb9V15tzqEDt5FxoHf1vtVIzdB/Qfty7zMRxPV0nt2jv08gUVeHqhteIV6X5vWnnZXTCNn+UNf
sChUr5vBCt8lym5LtGQI8CH15ieLTg1tNckJXcWfe5e5Rt+BKyJivkS06eQ+Np/V9YK31nh9zn9r
pfWuwXQQx1mQfKbASds2LH1FV2NHG5hPr0tWvHypRMBccdC3qRNZTtE1I/eIZPK5rZDQLaJyKaPg
/fx/+M9A+BPOpURryNImVTJwRaFRsadXwN56esfceG69U7vZ08WNzNSA/rcHydE3A4Uw/gjFkh9E
7t6mHy5i6CuSbHe8Pmagiav1EAaMCa2zx9bU8Cqu7HziyEkHtzAbu2UohZs23fpp2Snd/JAIor84
ku8kAd63bbFr+L4oTne3jdD9q+7Kk2/8zLmM9yRyypX9wLopghBEOw9gigQl+GTGxByLxEPB8uPd
X+seDLMTOXmHUB1UwOoqVAZ9gjp/GH0IHZRfCUtcbbZs1ZjivENYdS4D08tXOd1b2LRxYjHBfzc1
qks19zV9ciiMPGDxPl+5MrKxirLCYcVejePaR0AHYTv/ixTIQZNtS9d0kjuesElGhFGu82WxhS7E
yB/ufdQ3zH+gD7L6n8y0RpHutW5yWTKCM9sB4k/OH0b77+JfufhWTTwU/jOUGAeneRGOTKz+ZhIS
HWc0pKJmMwTruCJ410JsR5j2yLc/TutfzxeXfFQCMUBe9lEZY7+SYAC+1x/9f92i0UfBOAhP0vI6
7+QjNTKerRXVVuxgvAvYn1fUBoQhiQd/qd/3s2DK6lqxo1Bl4vasJbi00hEVSxxDDw342riPXpcm
UQ7Db43TWmUQqozM+kGWpN8de4KdW7XhPf9YSBf86mQAMkjmc+QfmZKltOHIbY9ucCc0BMbG99wm
jsiRRvJ1GVodxT1lF+shvJwSStD0ZBRQLBcGzchms8IePY0TXV4M4FT5FjxIh9jyj+VZLLVAgL25
fOPRjGxp4D2p6a7HSLGp1vIvNaH54LpZgamTCa+OEbs3nIWCsyAViMobhGCWtqVDl2C/7B5XYFWV
R60k95XaqqOjji2J0BJUPUdD3EiBx7Qkp8LqYRMdp/9IInBglE7YByyxdhipDs1z9k6Gve5ectwN
0DVD4K+qGL0ek4xk2H+ivRLQAZRtnkZBpklsquBEjl77VYOjwAE6k3LeXQbXQifwlQLjiJzqOeIi
VE/nplH5k/APwIF9EkOCLE2XgfzenbVVsi074fPyL9oItaYvvh2eAJAbw6SbKXV39qPoaHBVRTts
i2osed9irpHcL/jCExqDPfBrkYHiQRSVfYXZRQ0NQM3aDMXf77GUhGb7p8o2Yp2Y7GOsstqRHYmA
fUYcfYwwGQ4j2UxPwtGlr4MvX/XtFB8DMDQq2O9edn/I63yqBjpzuRmNE9Ro0CjO+NUgXVFOEPdW
59v9GlZGX017TTWIbvQFlsGwmqyYA3/Kc18Cvqi3G6AUkTlAuXa9lMmJEzq/QWPAnoXRw9bD4w5U
zFLK/P1i2kd+pfNMEy9ajjPc7LnrlSkOpe2HsdpmZakxZtfzfHvN07WFH9H4GKsRlI0Ox711VJ9r
9KEJMwtWnGuEYCs99HViEtz8Q6yqrqUHtSzw44ijX/2SHi9GzvtVlRqhfR6QCSwxzPQ8HoIFD2rF
FrVRwgkgx4m2zYh0KadIC37c0FVvuM9kRjo6uVJaWla0Gm9D5hpoG6SGiTh0XpEQfv1K6g0gVjvF
AzaphmeuqdG4TElycNM5GtsFeR9mK3MMqpglFhTTGnGcG33rUF3CrbkIlDCU8suy3poyk292lAk1
NvKLJesuG6ztSUQjNFNnraXd2T/Ky77drZrJHT5Ex6vcmiPBy9Yck0SAeGSOBAEN/fl4Z4TZbX44
3cP/RJ4bIgMqubpF4Fzt5uiKkmxGqadxK8jlou97J9LGGcxYg6X+Tnfd6ec0hw2a9ioEdH9DDKY/
t19PhyIHUHJEeBI3FBddSaIisQqXniTXI/3Mu0sZOcG5MvueV1lYz4Ek/P28uaASUU6ZKMOWWn/k
lRcC4ebuJL42pXtZihJS1V+rJlko21ufUtqK4rBPPT5ZSXRNMWLo3pLK36Mx6Zh4WcKj1MjEcoH6
soK3tBWA7H5AVE7XAfqFtbdfzNod2POXFcf3Qd/TMVaVet8nOQO98qOPfyMzUvwP14odEpRFpB51
DK0FYc+Az8p+HPf9YoW4ZanxXW5Bna54mRPVDDW9IURfL2xN7cosDzrMwkqwqGGw5jFc+UguS6TW
FUDst5gqfrBE0OhAiPs7+HuALtU9ysy3uI7kNwatVxKBufWT6lShIj8OrCsrs23oSUSFoxc0Vd2A
IE/AZ5i1xkEcfHEKtVcF97jI0M240D3YJR+SgwdR1OwgNJol8XxLG6AYtK7CEeag1BGonqHALxX3
KYW9TbwyVc+5zdUabAV3o/EM1+xtFAThNXIoLbOuBRX3U4ICfWSm3gRLHlhGxNfL7toXZ2GmhdMn
77JMWCbMSK7vJytSk33AHw8VTEXRnP3tk7U/XpOsm4AUSvc6mLqEfY+3Xm3ihiQT5WV2XMCtRcBZ
ECxM4i5Diw2txCgbK6fYbt/JM987PUTj81CcGfklZB43QXOIzT9BlFsu19LR6qDzqBg4vYiQpqh5
V3gKUD0THSoahMFlobw+jp3V21JGOaAP0+yATIgYG+SM24zC/GQeuL8Qu+6UytHrEhhBKETvl+aH
s46L5BiiY2bbRHaQSZ6+hUIKcXRdv32threM8qaIs4+6MXSUNEKhxvhols+AmkbTB9mP1on1aFfz
VHChVNcMaSD8ixGzf8ipmpfNiOlslv22fpeNJ/66a46jKPWcsPM15JP9dv7Uvvi+fBVpmTRX0NRw
/k/mf+UP1S8U5EfT4eUSqHGp6KHanb1sYJ/8rbx95inRh6FleQJh2NcLq9MOk2CyqVjrOYzgBJLJ
nM68QvP/CYdBbzMwfQWtj6IvGK2hveCsUbuHaqdsnzWPWBr6tlImwvJTaMAks78/ZG8Dl3b4nTcV
AaH/eA2VDneKKX1cZ/QV4BWcuVTTqg0ivBtfGAMcFZFsmVhNYv+jJyFwRdWWAv6mZhqQDVUWJ6Sj
J1B87Td6NHrQh1sJeu+yk/ZgeMG9tEvaT3iTo/G7XcnKG+7p4a4uybvKrUFlrXDtUQ1I6z51+0NI
arPRf+QwITPnflEPsyMdOigzFM3mRRoJoxkl/iVYkgfMfmuG2Bg+jkfilJC0EPkly87tz3vadLom
Iy6BcU9HWWiTdkez6KV2CpJrXT1ZGGr1CY4+VzErQo9DPpN0xAYsCqIaX+ibCg86JH2VP1de+A/F
mrPWzFVNNowbnmwTjY+JaDRfgWx5aNEyn8IXM0SBgPM3jySCyXDxZRxYxm39y22yHImyBJ4NYNAN
TBZR9JVYLUiVJZ3x3etabsj34YBEYuP3FNZYHEFcIjeRnbhFCTQFBBRmX62fdvRgB1Bf81lW79X6
B0fJUEwfsbjvbnDsYwANzX66MbvLmg7z0cp/OlQNg+E+3kFPBUna6EGRHANAXpDcnT4hKmvIJ/iI
4gACdJ2rMhbS/GuI5KAVtVJ05gjbRCdEJwXx53A7F1/CkOGpH6X0mci2s0sOTzh7zA1eNaiFiUt6
Eofw2gXuRdJT8DSvpRvjJ/4GHzc0bqbH+CK8aXHIdJ5FDKtE2cmflF9EiguX+gpDXy1uetPmr8XN
AVJVPCCUAwgB6Z7swtZsUBA7ySg7CUky7nMXHoIFAbr2RUhVpSO1RK60FBmkDDiVZYCJ1vaD8QRF
yGoia+8FGfOrR1y7Sr3lkfUeVUPkQDd+cwkkV43LMSEJtQTz6eoOV8MjHZinuDBamD6ySUCh9a/N
o/XFpY6NXgfWEe/0FJewZmPtWREFksa/ABdAbfw8Q7G9mgaYrAGxcYcZzO06HHUOiFSvNCXSCgfR
MQkvDx9mSCSTN0jTsr2sI8G74pbHocDqgfgi5Xrk8c/J7TJlQQOftFuC9AqRq5oMjgmmHk/3VkL/
rX0lkYqTvr6X3eKDUAgQL2TSeWbPl4Qe2KTHUimMxIzHmfmgaOyQhBPk3ljk4FlbsPK9Xoh957N6
n+CQ1WSB12wqM/n9AWtvtzKiDAKK3KOUEjJXjiX+dDOyj04hK6J1X7tKY7Oda1KnhoEPURxTj0c1
3XbBBOJ9i/GiJ7VWDaMchLxeM0WIdA/ruM9uOfch6njT/NpRssGCM4QxFkdxaZsiUcPpvlycK72W
V98puTXTG9tADVNn+xsqxhbFtrxAdAGMDFc/N4A0X3qaJg3Yi3m+S8tQujXGymGhA7/VOr/qWLGZ
c1AjfK3m3jdEAOACOIVgj8RFsedvmpcI4/M9J5TBnWAQ+gb4GKzaLPpPUek7zD0agoRFmTKSJ/Pr
zMLx8TxBU+NZ5GdUvRIiv4fhlfZWvWq/Xeg6a8QOjAO+Dt7h/XtBydRgDPcmCR1wxfOjWip4N4Hq
qdwWQZ/McHnHtWd/TV+AuPfe0rUOAqC2ZpOGpKZ26HRrNzyJs+J7vSY/aiVQaKqWwxttx3yvGxt3
eNRqulV0oK5pioqYBm6jscJkUBVUX165MTbpHHCx+lPGnhNEm8Im5IRTpTpoB/b/fd/pFGspYfNx
BEYM39Fbjh0hw8U1TBTBqWvJKBV8jqn9e/jZWlydSXt2UU3auGNdVcW0Z2chpzVnJOdh9xU/E++g
TaPpXQn3UinfwlvnSc/rt/6Cs45nOwR5ph1bDiLuABYSJgFXEapGoekt43nSw7E+7s+/d8SKXPb/
VROkPuxcag9ManpA4ChLYQGoSLC87WroWDxGAz9MyJ8tVQ5/RK1E+qvdF53yBBUOb5ZfZ9ooJ4UW
VP43IPJ2lRb63QUx38+7p/2b0sZHHfUFvg0hi62B3eUz9pykExTKNr26/tvNBBgSBL3ayQS0wG+1
Zjnd3Ofduqs6dH4h8X3C+y7RJFlB0UZghQaueME/G/cLUL2UJY/xSCgzzmAFSU6vo9iYxY1b0Xf4
aTwF7AryHvPccH5kamZtrdLJhJjv6mHcKLA+ns5CfOlL98yMxCS6/tZOW15C4yYjmNNNlsgEBwxf
NBOy1T4WyWKQqHqy0KlITuKqOav3mllRoE9J7lnHCxVvfHzcD9aIE90Vnt1vzf0A74rclukFfH8G
eHpGbt+ooum5xqbK3ICWEMEpkJl693me0gs+9t9sP5UPG0cMZS4V4ejohshTgeluCvc5TqoZ9XkF
TNpxIQCg955oXT1x89hWidh5KjsXj5Q6MbWbEt+qzM6dw99vIDKbO4ruRdRyw62/SyWBip4fFd93
TVsbuR3YO5SKuJ78exLntgG7wxrbaNtcnkrXj0EL+SHxATSdrVZKhz5Tjhmdh4ApLhTsxuhIV4cc
0zRkNmpMPJOLer1H1p0a6KmNChvJ6OJ4cL9+pIa/p5ym9ygM1u7pwvPqIv4KKhh2AIkMO9uOzBMx
KgxclwWqH4jXXLdXTtnVYB0+ClVxXuSL8AeKABD3ooTZYgyp9yIW8sB0apRJ2OTSEQ63oLvNB+nM
F//Zpwj8pVtlMaAZnFh14tmzn7gp3Am6NlsOPrb0V12zHe6IpMhiY/hEuEOAbwSIcimjKRB48ue5
STp9VBcVAVefsLcUTYYmXTXRgDVeLcs+cQqML8UEmqpy6Hn1oXgGbLN/v6THIzLOFrBGwl28THUq
s5d84zk4wRrhq1Oi9v/lrfqEC4D8yIkpMFFjZKxHwwU4S73CIwCqPyd0x+2AhMyEcMOiNoaGjVdu
6tD9lA1IzULdhDCJxDLezH1d2VPDst/O3BQZ1MOdjI55PZ5shGrtQ8XSJGFkl5bf4WF6Q8PiJyWu
tvJ25zaruJkkAV8OyuxVTQxDltVRxAi3EB+d9hGfVf1Mx8J1W2Io3Y5Z9Y6QfY15Iayn9lqvahdg
4o5qqki6CTjDlA4TprC6OG0sPXmWAc9kIOKMPcfpbMffHLdBBV0njr5LQshc7sPwFdhxJBT5C/m0
1ccKOWf6OvYYlT/KEsk7a5XW5+mStnqV/JHrwWeYTBfJ4bvlClOLad9dQf+BUfgFq68fVC8pecqR
YvHYY5rrr/vkaUU9Opt3grvvkdBX01yJx4TMabWvWamDZ4adoVf7bLGO2ivMWnOs3onfctfVH45j
5Z8ANgGj+eBIP00fyMwMoQ3cchIWLGZki/7lznVoxN1qohHI67uF36oEK7E24wiK3/h81MKSotgH
Mmg5parpoLyAEiC340wnVcW/tmLkeH+xBXIaFfDYA4Y7mEUZMacCRx//ARgwlX8Pt5X4DDriZohH
vEEbN6GqKCLBonA6hihOeyV/u2VTkxgU55y302KCDkkLnr5dzoLrWbMkR5c7dNhLoA7E3JL0eziu
V1SakHhSngQVh024G4IYVzAuCECc7RMGZz+kLRrKViFoRBfGRXefwA6lO5WN8/HpJpBmQgJZ4dks
jqyTTi9Bsy2Hk1vs0uy8vxuvIF2Ll38GQkVIxQbWwxaw7ZGTKoi5QAMcJmdX2Jcurqt6nRkOerAN
O7lctPQs3aiYiOnaMNdFNHHKoMmHbiqC7dn9HsaxwEduiVNnCfm30CmPhAodv+aWlaAi+QlNgUCD
TC2mnFPkqIgUolX9hqKckWE19ffGw13bPF85AB+GivWyJmb2n7saQfZUxPr66tzp7QxxN8BYlrOK
C3P890VGVI5nwWMoDrWjlmhjuk9WXkegoZCFlMe7T0wIKexKkmzYbEoXAVu/JEShbUwQFP8v9B8E
O1+bWKPCzOTO/aPvZx8GoeSmzatle0QC/AGSHt4gkQWOcSt0I+FH52o8Kgt5V0ayQVqjeYrwAfpt
+U8uSJGMeOEOwhfSGKlkEv3UdHTFCUyQOW3LlyrVsyTyHA9qd4dX8VpXZ8xkkPD8GFg2T70fmzvw
oLuLo+1+Yoain/GFoY4KHiwbk9FtGxiRUMv/ZBPl5I1bWkluv96Ep363PjDxWg1iGBpKGjpWukum
pY6VPZeeVUirDRxiuFb1NnRgEAe5KugZbgumulN1gAzFLxgx1dVLufcaGvJUSm2U7+h+fGgU9li6
BJiCgXHrpOM4yV1yg5aAWHH2ZO5Dbt2YTV6K8AQ+XWKbq8qrkT5zxjbNH7fntgNs9maIdZsu4sxl
LyRgZQdXeAxs5ogveJIlTBB/aqsfYmnGOI76i+riy6o2eEbLYhwdP8XLQMi7yheZoUwu69Kegd0S
vGoM4hmFCv1rmijvDDqn5yq72nbGg4mBKjLxUhKrp9YfbK1vfgSKGeCut8KC+HZ+ZVCLetgPwQ7i
uo79fYNJi+LT2LFROE5GQKc3D7xJBzpA44p9FCEOJxmmySINzcehtN7mYWQyE9RWpbI4GgIJT33H
DCea6+Urp2bLw6phhlgw9OrQNWXMTL/AQ7CpH395AWvQ9ZKyGaAc3d9oMBDlDVbPz8MamBQVPDKL
0YlgEW4Aj9iBZHv7PdQSMPU08dOSh4RJfJCXtWjVWekE5sQkwVrJd0RvhOucXIUyPVzJ2nVhsLF5
bDN3gk7bSxSu0wUukwS/P5UkyOOzHgJOvTVa6UKnarARcaPR52QFnddIHI02vB9Oizok38QXJX8I
N7EARR63sQ8xGnMYm2FoAigFKwb0CdBg1wzxCV8bjbTc4HfAYbM29LekSyPWxvzVhp0oXC640Ajt
2N9P18anQMxi+pttFsGSML+JDSFqD/Evc66BtdkDmy6nkyVOqxXPzzXLwOIXiU3ea/KnyVd9PFYn
yDAY0QXp3DCCPTkw+seuLuTh7eHEDSZkK25eKOEj9zwkH+nj2KYUSt4s/brJADPkWvy6YTZ/klp0
qxMMUlAP90D5Ryqtjuhg65P1PJkchcr2E+InujlLptnqyayQuwLveDsc7vFH0n1/xHBj2k94+Ksv
OjyclOkXOOvwS95JHjWv1mzRKtrs2CtVNFK/lWSFU+0vj2S/OfU8zwNH1N5JOVOctxYynH/N7baA
PbeWhXH5pzEny6XI76/k4w0J9dLA7+MIBd97GyUNnSiWvIjtb+3v3XlS9bSK6gX3/1VwvV/nOUIE
eHBWQFz97ry+jgg1driOTadZw9QfC56YREccaWrvpiGBJ79Ggo5wrbzmaZPkg9JLjnJI8XFdOqiV
x98eAfbRIFyScpf5q9qctPNb1E7rBhwbTWEF18krepGlJvyYs+9T6qRMp8GLnfoq5QFF/qmg6Gtg
D/ifjCcPkUl0tKjMNtmCfPJU4UZn5kshg6/cmFb/lwfZkXf3TvW2FrGHVP0VFuptV7rYtXppB/ua
1dDOTT9ydts62hCWQbBaOlAFx+UNlTN++gqxUjE0Y9fzEdtLivMSmX3CiH/yEJsxMBzfsL67f4yb
ooZqTsbDh7pdSmA88GlGj0iI8qRrrd14nxNDTnBT9IeKW+VDBMGVW54dVG3idyCVQpcRiwqvntv4
IBih7Emm0iza3aanNqWd31yXYC4YMtGUf7xb8znGEnFLGcXSSlPTTO08gCJFGu9g0ezuvYIQCfNk
tzRqhttfmalpeogQntsa7KeiYfecxZ2gMxWzX5QjVMsqjNZu/AWuzpzHbgRknGnFbhdwGY6uP5MK
ACEIyOeTdvqdi8VQ7yjOmXZFe8dTAxavTG98sUf/CWQdOnUu15R1+1ttJ9ge3Oly82uRqUvZLY9f
ueMBc7R8ppZWkjPnz0JYMYHGokvbKPX8+cki+GB4FyIQi+icXA3D7VNPOCsXFKRYH5YDdN/r5lUG
2KMl1iyDR2Xk3qKWCU1QnfG9wjhi7ejPa5JqMnrfIQukKdar+vdQCWQZo4tyoS4cCqpgD+TFNyxY
jxU4vHl2RF7T+zwTX5DfG2d5iUd/WeAjkVr8hIQVp4EKu26cdl6zJNGXqL6RBX6ahv7pchDihFHF
5AxiRzxdAeQJU7inwgc13FibgaS/lb4ABRmwDQXgovPZCMSdkYhE1Ofiv6VRfkjA73Lqug6GXXpT
efHTfGjvIQXvbm3OcjQQJBbSGZk2OtNg7jNb7RDW9T88bqr0BDrM39or+pji8jo/VVeLUTmXiWIu
rQkZ5gsb4/gM/QNQ7OhwTO1GmQ5dbjpDkqDYlP8PsglJ3c7inNRNlBPg/ziaL0DihobP6eHUbZSy
XFxunlgPs0lm0CgBJP53bkK5tx62Yo5QiwNyuUBdby9PmfYiY7LxGG7bFKU+4FVqo5eh1kfCJprl
2hCFOYjDcFNXsjMhEbW8tsXpS+HsHHF4YHP7pNlRgNasPCktF9I9gAo152OVrRR6R/jRcJ9KTz+N
CQFWuRuYci50e76X/n2lE+0eF3VrrbEGp2JJb/4xNeS64Kq7flYbW9sUP/GIUG6fPJk8gm6EGCTJ
OB7sOKEz5fBnJPydR2Hnieqyqtbu766tbQbuf6qz7B8jmCqeyTHelF+TF34pMF5ZGOx76NwbfkHt
2OB+8951EOqZgCQsWICPTBVCXUM14n0jH6rHURmoSBSoGOcPjwxLUm1Ieykjq1Q4NG/LxC9rLjYO
F3xzHb5+/FVjfeC4MsJ0KYMjkBhjPHGLW2YhRfUEbPb+pGNTB8TObaOV5Urd6yfuEKsDkwU+RsND
nJ7YhsfIU5VpJgfK8RQUDMIroMF/MixrI036KvhoM5cqcnl8uoBmize97a2yDDn+0Y4LVyIB9OTU
yjH8glu7bZWorUPd76bC/9z3TfNIEBPnESBbQIKokubsi2YQ1zsolSo4eT29B3IydAAkE/iZc1nJ
JuP/he/OFy/DpZhxTqgkmsDB3aUCU3VSqOlRonwgrTWvtS5yZRdyVIrI+HP5EL1l0DTyQAaHwS8L
8XdYBVEt6e8Bu+27tmkc9U5+FI4wbKC9xdKvb40PXOXExJPqbVddR5Zukbyb8lrpW4Cncyr0Cx8f
5DOy/CL2qYEaUb1ZRP7OsKJs8+qRnjgQS42HM7MrfsevNnYbN5+xc0Ej3t6GTdY34k2EOX65UDTu
zrURbYw4lPAfE1U2DycmMM3WB3hLbc1hFNz9jCxsWKCx6tNLjd5Z2uEqf/SXjbypKsqrEQtCdhVU
50dxrb4RSM0HWvmZcV/3UhZIDoM0mWFs5EXBYRkSp6id8JJeIc+DSQVmJfSrqZqSbsmYwRwXiWXq
qj3frEenGANm0OMMcBT5eJVaueoKoiPi+m5MWh3vMCfgt5xPZsSB1SG4EME4OB1aw8jvK9jsOllp
EitKKWvnDQ46IrX3CJNb4m0q67wNBPQvwn6KtOIsgJjPd95bk8qKAslIJsjPR7HZV5K/k/UuqihL
wFDqCrK4UlMyfvU9I0hFW3mlI78uUZFyhF8mO3TLGSqPB3FtXfUIrNsscO2PfvxVHOhUHvBrMQQE
Hm9i6o1zqjBtIZnKbuV0ITY4PR9jfKO7bBldu/EllokD7VtOJ6dNsWr0rL+lXoAKGqcVABUK4qUU
a42c9R31sEYG8Ip1oPaeDa1wA5Ce6Ja0qcY3+IrwQaEg821GcC2WEbD9Ne0Qlyk+LwvqfbLjSoQq
QjxrP9kQvEerOyxULImO/j6Ddx1ZLxLPy9lio9BkFBU4dI3OfWYog+9y6QXW/TpRh9Pcb9WiTT0H
Rcaowk2QPbcJ8CGTx683S2VLVs1VZm+Rrm1Xz6tcJMlyF/JD2gWKdxrxhI4Lo87j/ypsRuM/tXla
8viWuP37f+lkvcPzRl9zOFsA/qrkrd/NvK8ph4SKUZZnnXLjCNllvMYdhfK9gg7Uj+eV0+6IGmdq
OO2zy4HQyxEZ5VchxM7ZaYcymeI1okB1Mcvjud8y2lFP1n+DXFVlUhs/9N6kH/qi06xICVZrnUYb
tOA1ihF/zo5Hzj22bynR/IdB9sFD0LzG0fQs/CM6u0vGe/17zuzXouKpHjxeZJF97JN6g0xmhJct
V5Uv2oOzJNiWLWCfFhg6d4yb9JPyy2RUjembztWWR2UX2GRN5yscG3RMVn2NqcMnx7KZeWbZgZBR
Hq4ZdwIredigblbQZk4ZsBO7IrNToCGhE7cF/xnx0WRRkYGl1jKLaINh+hbPuvNN1r0AlXOE91lj
DRqz6RHVDFfuzgm8c/16TqTjQs7lx1eXQx6Zb81yXrl2ZAd/DUggqMpBQo82GO2RWHJbRPpR4yzN
bC0mjsEAZ2W50ojw0F534tzxk6SNmqfov9He0PWGlwBKppjJ9hIYcUwIRqRK7z8S/pgR9YGC2dBh
Wu4QaWOWeSb0+vwoBw7CRtEsUPd4DyQNBQo9zmVeo4/3Q+vIGqXsJSFKBdvHs5cUEyReJ6XTqi34
1SpMD5ZXY53Z1yjAhpK+rzFSiiHs3SPk7am6ejJZxI7NIGyN1hKsyD++NkkI3H2giPeDdeWO9TEg
k/eaesJpnzNGXNoCzUhvpTx1YHVPYWcEzoJCvsDSzdR13oPPpl5DBhDi3yjBD5GukXF31mHEGTNH
KSchmdHoKqP3cVn3aPAsqlk09XBXbqrm33nn/wy7fFCbViczXGRzYWck+EAuTTB6KxytaljREB6l
s992LZSM7UUap6AQ111gaDXHJFkfcRClrLl0TCiKTHpq2qVn3sTYD53vMSAQsqshiZsMmTFfCbRc
b+ZIGMgaf2hX+QY50GbIHrhsXavwcau9vnn61hbvjZTYr6GFMbNNvoZGuJabigkHH/ooGDrAL141
vs3T0DLI4Laa97CnGybD+ISD0pdqeIo29iIkZRgQXjyy/j1Fhs4wXVZspWHhpUp0s0x3h0K8MjAc
aU+ODjCWRjtDHESBp7nBuRRpFFD/D+qfgMPKAsCJ5iOdfBWK32luvf/xpEUrLC3l0aRcKLzUbLph
qID/TaE05VU/WFU/+Cs5YBAUGb6unjaYGugeBjJrHy3H8bGTnoTjKLh3YC1i21qsj5ILi7Fk2sJI
0kUTZfXGEO6jddFO26AI+jcshG6TFVqYr+gOlZhMFdIBZnXwnWBPb1iZoyOSh4kbZnhPrPnMwdCX
Q7TI7NEDr7nM2WzVU4QmjGOMTcdCcryrW3HqyD53Pr9ENDFZCYQrGrGj78topChg0jbKIh7s40ET
3gjwH7pVG4teu8xYhRbBp54Co5j8ypPArGKa4bTNjQRRjL1rCaIi2Aa7X8UrsTgztaefzzeKNgRZ
2uzJGYkmjzwNQAQn0mdBLLUGYVlKM1CJ08Ip7Ixqktt0B9/52539Ae07/CVrTQ2yIKPos4VMxodV
xPLaYStRJy0J6aIFXe0fqZnmLdH2l9Ms58MUFVESFCNh9Y2OVmkiaV3yWGYAuOtxJM4YuJ0J2/JB
y/WzHky2G4QF/3WwChMlJlFjc2uwNU8LPBjtphqAvF5VC32nk2oNvIaU+jDtKNpvLWhWoKQ4AgPy
oyard7bSr2ho/FUbM6Y4ZEyHBOKdRVy5h/4AlxLiTlVC5urP76NT6R625t3HtP5hCbmadp1BZ0jd
7s8SVeZgnf84Xe9H98vw620rsdff7Q6QgvsgcL94m+VUIvWU64Sbpp306PeJx7Bg1Xv9rkskVjJk
xbFIc8lwuJMeLYIyBl57b7grFQy7a7FwF8f8GA1ld/mb19LJcONfaRKLhX4aBq/iiCrbICj1nhxa
WuAdQ/BDJTMljmYt//1oSyW1u+CHYJKQIbiMS7KfsXdO/2OMovhlOyvoOdd+ptQw/oVJoWyPQBEd
Ux+m1RVsQMBsu2a3CwEpINJ1EnH2c9LKYaSQgui6C3dX9RT6CBFwFe8DLGMSFtVn6u5WEqZlJfdU
NvtD3pCI6PwSuSL3qOUkBPG2rXiX0jfO7jO1/W4KD/oUAD4Oaix2RDt2c2wS1/9tv7hkVXQ6XRfS
xSezwvA0BybZmMuWFG4MunVFL4pJKyjtv/3FriXJ5UFdKsxfz53IfWezkn2pgyRdhatzPSXbev+y
l1H+gQQ0vj752v9lE//0v9XjYDPNUvEooGOEyX8jb77D7Oi6Sf1BvaRI4cqBEl60Zv0p4Y813xwU
WdXjMNC42mN4DQBWWUnlMg7Bjktx+xeRF5Y4JTRW8QqXx4bo74RgmIH2E8TB5IImqm4RL1SCUgpD
hvecFn2ka6anaILBOKBcHpIThhJCyqDfoca8mTWvMbO1YREIgJ5pABfyU+11wLLBYVKFDSZmT0He
uLrPaQdQ7lXHLnj/VoyQNg5woY/c5EoS8o2LVLwfFN8STNTnSqzsDWC2ZNTJnaOKqCWgzcTzvTon
qMC167HwTHETj7FzlRVhWHnRm3t+9q1xa4IHjd82JdovI7r5vB5B2YHsQ2u+Cz49ZePyZ6VCcLVL
48v//STXOgVD9uovzHuOpud4p6YijBrHMnbhY18DlbyYwlaw43APr+RwaPcxvKz1WIm7PlXiJgBK
XHG1wPVm/RgnYTUqRET3P1O29eQbFpydaj/Feyrb2nthbzODRR8EJNB/MpvobfccpQXRfQPJKH/x
mQZIN2nls6ozNsYnYkioq2F5Zj4R4NzQGh52wINzORo3wzPoxV0jDRFCzh+zUwwjdohUUXzz/t0l
QJNXHHAxwZgvKU+SNxlmDAlTTdUC7HBUL5AotF/w8PUjcTxfziWvO3ZtBWsdVoG4BO5Q9mwlNJcV
W+I9M7BoPPj10kL4Sv6oPvU1+LdKU6HzpUyG98uRNNVO54ownyKf+DiSFuvLgiITckGlSYVQ9RKr
OLjMXAuPsgs8Wae16NWd/tz5dIoSJ/0drjG3LgZ9ftBveZWZM4JwxEpsigthAwnuMe9eQEFTPBXA
A16uSyuGKD6adLOJIn0W9PvCLce/oBUphIvRRj6QDNbyYXkbsMeJ2bv2LYja9i/+SuAlMpFxT6hM
aJfAegh3ql7bHMgwoLWRU/sUGReVFbkW0HQk+Uu7IApz//OYeHGFpENkJknQIedO+SWPCFvuNtM3
928bTpNzEVD3F21JIJmFopFyT7ivdA19Gr1kXei05yBLbrP5BmD8/O85JP3o6CXgeMDsNsX4gRKt
rctkWB31dAcFO5+20WeHfxd61+juaDYr1E2PEQ/65QkJf4qcsNyNIHoJu1lhwB7r9KWTBLH79xYp
JmONDj/p0Y20bdh7w8QZddEx8lGMXxle+Zz5MUmHRoGzkid/x1D2KDbl6npbwyX1vfUVlSFv7Jii
IDkiK+xjTFTb1tz17l/Ht4igKn6KMK/l58AerbLqxF/IRSdWlK85i4GfBxXnWAkM1foAOg0UFVvg
G9qgtRNS+25vAxzUfl45mGkENJJ/kPetenXG8qYo3TzgbbAjUt9L08junGhfIY/z4zr3ICoANAYx
ZDGvoRFp5qYXq6IHmQMSLnkemG5gI6vERMBV/xbnudontJK/hlc9hbOz8IM4qNINO9BHTLzcexOF
jYw/Ms3c6EPKDMlOp9EXKR4eHQbowvIr8wP7aDA2E4m+AtmZc9Ik9tyeWjb9n/NOafT7e/GuL27f
1esyuTQiHUVdv/QYBOBFXWB2tZGkj0D1ahutQUswvzkMsEVVFmSjklwhTBxBPh3r0eaEAYYHZV4C
Dj1OnSPlSaeTuje6gQvzci3PM6pFCzzpUlwgtohqAqwYz3l6DgNKh0vcs/FELWoKWvt/lDtu8cbk
tP4TGwXIiCBMcbMBgIf5asVq6OYZGp2rpYo1hZ4KQwW+bLjGyqCkuXphqY0glRzr54Fifuo/NrSH
NCtsc380s8de815Tas3EjpapcCvCH2SSt6SMf0qWvJJE98LuVU3mOjuogEOJ+rEX/bzTKPLjAXhb
ElH76X6ylPECYrKpVQ0ra+L82F3wpn0HOyWS5lsNFEY7FdL9Tgudsj29yOhC1X11z2occrXj7u22
jpUj8CFGzEaxZ3QZGHSvcjs1tp7CH4zyzKHSB9ZryV9hWLVanJ+QLUxhLe8eEptCmqVtsFQ3k75C
4OC0YA0DP0FEqEM05qseFhV3V5/fPvZ2uKVuGjZOqhIuQAJZ8rf0/5aFZdEu7A/lHe8wFtRwtTzd
coZnbr6FwXgf11TK3NPOEg7oeLtXvKmf621Ytuct8d3BzPHwD7n4O8HPP+f19Kt6p/tYz4GGCsfF
v0EfMPBELcyDjr8wNlvj0YpMO/C4VyfvlzpqByuxRHM1poYsABLxHDZmB6lokEFvMsrDDOY6xFnD
5+StgrwMDg/hVKp8xrBhnJ1WdTFokqZr6P1M7riprJdYR/mLAidgtXhqrDSb+MfHvXFYiRkyZaDt
VN31AnH87nz6lEHgPijp/FNEK+Xs3YGfc7Dq08DScr0np5kWubtE+IKOD0bNAxXoFs0GeLhyhgOk
ITRyCSUFC/VSyGRrEaR4p4iAe/A27LAdIpBcosPB2NFJTLTnBTdClmdgNMPkNxI39bJ8/hVnpZE6
j55+KoJTX0UOpSP7royLdF8KtaUTPdG46YaVN4BZdIK6lfmqChDImFD5/qWYpbEeHj3+QTEG8Rtx
ICLYuhOxPtsQX3nEZs6HBN14ujnFFFzT1VEBdDjzkUcDdPjr3M8Z+gkJ5zEKFJ8yTHSiRLWLcRbC
VTGomtS3dQp4tX2I38ijGp/bBAISggTZJR0qzxJ816iG2CK2fPNRc9GbkoBZ21omBiQzkO2iwvV/
PY9+nL6CwoBsrhX5oK5GoZXUhYJ3K9Hf2NVqrZPoICJ12XEZWUKMWjpJpBrQYnuOIGxWbaao1Ty2
U9t+x2eEQoO9kxx5U+Obe4RcO9zv8GMGKjh0jtzxQazuw1y6sZm2R4kvDev/I5MWIkAi5nkkpuJ+
gq1iMLICH9PXcewUq/F3uHkHmFNKl3fI2fUnE0SvwY2J7pAx7mlZpksr2LncLKHV9lrFef9nvjHe
OBxiDpLr56OKkqISOLFodvxpud+wcE0V/Xc2ZrSuIvEtvYnD1aOBEWZxiFviHsn+PGS49oxs92Yg
7Mxhx6ItKn9qFNoeYvfLyOOiJqDtjdC3L46TqzCDTLr9kG7IE6/K2iVH1ykvPrPcHUbyaKi1nUu8
M5t9evNlIcuw1zjOWpL4Q2LiobwEk8GL089FeTaaZm3YIboVYcincp++rsQ9BzjgzQAvIsB5pTJ+
LkKMue4JtAWs6n32VUrx2YaPgzCDpkjRHAxPMTCXRQAXaNZk2BrJ1SBNaSWDPLEBx38hZk+dT37X
qIBaE0DnMoQwxPY35cVyf499glqjxTzjTUBqRyRlorZEVqBzGWbqU1VOdT75SZqlgVqsSWyoiKSS
cp5VWMzhZXchtsBpYINVmYx28hIrOvtKXg9+ylbN+b2OVMDQpMrsFUrPV7xD0RhCR5mIBfIoIBtz
p/iapSHquAgvFRVIJ8/PL4NMzUsG3iafkpJps8l2L0xAVBFhtcRrrj07PBEnJOyvDVk/btFXychw
Mib4LQHl+SecElPXNBonNvPA6WtYarLg9KL+EZB+Y107oi3lBnFcK9tgm3KTLQo1JyQ8uIvVED3S
uuG2mrjrlr+LEwfW0zK5cbKUAeb2Xf4SwNu3VnmEbN6TedRJlqKb2cslPsQDHpCxAM/A6aKzI/5/
JHYCcgP9M1kbD6n6UmFy1payIVyAGrl9WtABxx+o83yj6pUr8EUlvX9CaqPvrVtZ20qHj4cYAiYI
g4U9MZbvngp7Fv1tehFb4xPsdeH+sOBPHPoZYTJTwKhBcr3Cv3e3z6jmG8XN7KJhhX3HcEf/sDv+
zaPoYedpywDIDavufXJAE7zRgeY6vRJzsOW7bZEiNSmJU8VaemZvArME378bR6YoM6mj7abKi00N
OOEPvCPUrhyfIss1CiquDtN5Z/rEbD+0xcScTPRL7uLJckVOLhlcj3KijEURuaKIGQhVWStqTwpZ
+i4pwVrz7IJgdGx4xeqSiVTa9MoKpaWxk8cVDm1TiDGuDltLjMcpvok6Rgz3qSeUkr+ufq08Bmd3
4N54S1YcXk6wDCMiCH5lXm+EX2D/M9oCEeWIT3mfmQTxfikBFsHPDjTqe7QDmcyzx/+GNLAGvMl1
aWAMfMBnv+hvMdI/o+fnHuvTMD//1FFHsCOy2EWflUFo2vETDCJZ6pgAXW77O9pD8nqTgQmGzGRk
orDqqmSO9Jdp8gfA/TCQZfvANZoKWFBa/gzNzUNtSSdpeF9kWwcOefuNcQPAJ11Rq+tcfWN7wqUT
ZTpLoUJoXkjPNGzqaSBWw28PeoX2daw9BMUbDksuwqShSXXhlceIfFV9WyWQZs/4C5x3afKdoPRF
o5QYNeXrERsTLF17fd7Yi7djkFWHWoUzlP7LfDl9yemKWC5llMFvLHoJM76RruzOXM3IxTAuwIf2
sjISR8SdsyAzWN8gHIlSUfopVmhNnvkGegR8ryEBlCB7bAinIJMNLTXnZM4bR/wB//S7EDqMIgK+
ioUCXKTwBfs0sGqnMnZBckvz7PrtQz8tnU4tFuCJw0evwJfCvkM+JMNSaV0Oxr5WV9iWZvyHjJvN
h8fE5GLQ3FfB4i0G1TQo0Y8q+LZD27wOFm5EZjUn1oBq9aNRc73qu4jxHihdyKGcsNv7v5hfl5st
6TUExOF/WDo0kBiMO35mkMMjciigzIB0NQWcpQDe4oRrnyfy3ytXikUcJK05DzugYUU1On6V/kGc
+Cq/YripVFGN31gkVCcm8HazeO1h+ybepM+gY9MI6o325MBnt+pihfcDYg4p7jzndAR7Gjwb2uE7
wGdZwa8FMlnkPHOeYoE/SDrNl7/oUr1LyiG0axFpTSHqs7IfrfRNfaFuNFDXmpNRAsj7lj7QY6YH
X4s2BqfeCubqr0qMvyYIOf3j/Vf7CY6Jjqmcot6swbcUFPQnhZNe2kpN1aTa/jBJ3Za/Nt491ne0
q6JN26E7M6RtFa/AZ8nw+8Vp4LHFNxiHGdHrmOrWC7DJsxTqzrSi/WXQ/RTyuz437caw5UL7Ct4z
cdQGy4OUiRzcb1XeZm/g3JMOLTlKhm1Lp71mt4m9Xlak07ynu6xY4dDfIuBsho5KOmnYGkhQJZIK
K5YsWOu7qyHIN85ZFURbImRq1VJmLXtPPNfo2LFRaJFpGNEACNZBc6eyLcXPsdFFmwzmsSkHopEw
hTgs/AXfvm0OhIZUYhOMyS8csgwAiHWl9teEv+EEVSV4Ymy9xqMHpnpLOYIuE91mLnkRgnywG8np
PA6rTRVfIyyVngYloHu59M0AI+yIc3Ma/ihUVE0RMOMnmEzXPwNC+yH6P2u16+W8HtqhzfDHIazJ
7DP7BdBAUmEVqCNZQbrqyQDkwFdN5QnF9KZOKub5EBuKoK2T1SGydXU91YXYrJUkilgdmP6FKnqM
jpT71UzjZnhbvsZ+bj3FKGE5WjKWZ3x+l1AteiAOU/oQD9qxx7K7/pHtgzg69M0RnCmz/e5RKPYF
Le/wPPDmlJZPICl5NKMOy3z3N144+I4ehzjxfBNnl+AZ6NV7VEUzZu4gfK4SifBaRzpOCZRr9hGC
IHqbiRcMKam3MBOem++8a7JDazMMyaGgipTBhmgpSL58yS/b9SiAJ3CRowJ45RWk1P3Njdjb51Jp
1fqHujWlsO2XyyqogGCW/2sD1+Xkx9SH+Ouq5iU6ZTmF+CBGzm0Urwu+eezWSedaiCkrnhNsMFRg
vdXJUqsrC4U0WSjWUeFKjTRCyLQbVY1WvoXf/xdti25Nd0RJRYf5I4A18gU0ZUFs3vu7uQzPvPMq
+Nqlg8+aJqUk73N+4g75W3IzrtTm28URHNqrJOIeQK2AdIRjgv6/zckeecwJLxMZ6eDtQbbMthBt
hOmDR5MG+dDiZIalOGlVPXXAiIET1lDnydgi4IPvwvtKXD6UWsmjEcm1W8EaV3bcKR5myGOeKSTD
IRtZzcUNbQnwoxUmWj/yYIPLaIooTZMizCjjjS0Ielygdl74ktS8K5z+UmS804Ap0LYXaDHO83Vn
RL9mYBmix5LOjGDBmcvYQevjkVYkTgWg096/2jOPhzCnigtlvLdG8sw4gvbr2IHYIE/EGxyM0jvm
yBxZgwXIXfGQb6isDrGhGQrLiywl4KXigtcAqZ/TdRrptf3u2zZQz8uRrZIpazL9WN4s3cqkYDEz
3fFopVUaf25h5BiRCYBW3qdZrQ9P1940/M46FiZQx67SGxM3sFsMzGZCoWMfuqUKLm99wR+OKMuC
4q/vqMNnuG76HSuEGFLjWmd+3CM/RGlxt7qw9cfHaNnzRjrOSIBAEH1ko4s4zvh0989cc/yIMohd
lPkHPX8bw8RrIZttG+S9p2+e0HrLGga0DxnrzVgHg/yZUW9tb7YOP8pTt+UcWbAi5WWUY3FPRwOj
mwicwLGYvwCl1haB+Zb8BL49RMX6oro08biq2dIz4BjpmUj7+0b4PUSoWOIAXrXoXlmtcgbY0Lq6
88Pi/oGbVknbSUUt57vHNCReT2x5S04vKvb+9NbbPW8Chc3I246G75dw+dhSc9geIhr2VB3iTVG3
rQTq1WPMUK3t+cmp9sVgLKvPI0z+posM5kGViyOhPRjBOozCJzPJD9o1BFNqimCzCXf8rYQxIVY9
zy9sjBC39NGPTwxUMe01wRMio79a6D2wmdrM3Brqv6pDHdB6T7kRFVpGZybIyLemHue9/ZwXrACd
RNMq0gUfczbrGKdHieJfrUcCtyCufPBie2tnZ2eY2TxnGfjOXq+/mSpSx6SpUD+LaQKDVmRniB8J
lyKDhR61ranFafK1YAglV2H4N4bpx8xnVlyEzugNMyMSann8+WT2q+O60JKKttvoUksv4C7PzYu+
sThVWVHJh0PSYQ9TE58cs2jSYfYSJnLPsNW1G70ogL7z6RSUCLh9oXtQ02tGm4yVti8NMuExavfH
0M7oRYMI86qrU2JJMgscXUDGZ4NP5Cmw4uo9Slhn2Lp30P0SxMWKTjWpShZf4yObITjNk7u8JZsD
ZjiZL/1g14yK7l9vfimWbydgVl7yPTuovOXeyrkt/TdjiGoJArDzz1uU/oMhStvxdp/O9wJ1dAUH
ZKDWiARXr712A4XxxOl8CweLLvAOygT3TfELkRItIt7cW7FZQJagTMJH3TmXpdRUNrVCiMNyrUmR
Fe9KCCwmKDhFLxzftd68P1OTWPziad/rib7w8bgkzMwFI01bi4BRPBkTMLZpZdKCoVfbuYqw7OVY
QmNLQibE46oR54pF75//QdGkTUSCK+HJBgLuX1LEdIbbu4Ypk66+NbrTOI42iHYjt/OzK8xKHOzF
0Q/yFdpBvjqK2AMHvsQHFCf49ApMWW+XOL2p28ozTjJzto+CrehC7APAqKtpFUxZIs1ML0QP7BNr
967UiIf7sf2/kaAG6BJzgE2HymmxYrHZVrGAcoBEOP5dDXtHvWCwSwPudUUt8SOpDJLNag9hjKJj
EvZbcTqWfillK4+NGJ4Eiq43SMFAaGorRi01VjdofrVxiSuDWxzoSiQYjs3DKI47+cL0drIQh8tm
3rvT9ML7TmW56EYf4+x2Tk7krinJdvAphTMmc5WZDxipxyGWZVqW0xxXi1TuAZYCgEBz3bgeccW1
UONvy9v2x3cRtCmlbo2wLjASHaxQ4aCNNrFdI8zxMRkqs7bjOTyZZ6H67Kg0+Z2OGNclgsbpA3gU
hRjmKo4mdN2j4kw/qHbS2XIlRoAfLoe1u6KKsAecdob/AD+sIUn/Zj2/XG9jMyMFTWdmlYuq9nJ/
aMhyTDvtfgfS7cZv+V7FUVFn4OYFp8sjz7qkBnJxlBV7pOaj+kbQ1Hx6/67B9N2vki1KbFhVFE27
tFs7YExBeCoUq8le5W7/nTuQaHbd4ekPcobQfljjAyvNbmXv8DsC22+bMBmJ4rBspnqvU7e6jTfP
bjHXVoiGnxVTq/BHrnf4Zgb6IcsHkQhRYWHtZbhLjsjL6NFo8Au5pKoMupgWL8SSpNUCNgNdR26a
CxUqLhXbo7ICumgte+05heGQoCehJzKqmML5bpn3FKVlNh/lDZJ/t/KH+K5gMlyCYy6V/eGX7/XO
94HYY8ULiA22PXu9C9rIBAcSmpXejuRBiwdSTKifVUnYrd6ISxOOfkRbIpFepbtbCMAP+unXG944
6zs/0cTbp6ivHAcPcMNlYLPr1qVxhPLCjKUnl1fR4V6CRFOWgcsEzUH8KTEG5g==
`pragma protect end_protected
