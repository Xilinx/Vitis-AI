`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40064)
`pragma protect data_block
giGA109OWTgnmloyaK8oODsiRC9RZVQFcgf9mR/obyjke8kkfwHUD0rFD2w6Qg5sKJtvAY8b/b0q
V+Sa+ZX24LFU4BuS1vxLWFGohu1WaQVSB9HQcsOWHML849yQr1UuXHS1H7VUn17v0E61+/PqUzk1
X19/pJmyYW1BM5ZHOhJulHdCd99vhdUA5znwgIeL+qkiU0sf11eCHljau90FYmDoD5m6woWzKvoP
6gHK4sf+uEu6z5A+3PvW9Z9m55mkt2a/UNoD0i4Gx2DEeOPjprF3CHknU6QtTGQAHTnbS1uZPoNw
J0Sju40A6smmy7thIuddNnRhbf0CPzWagreerMnokI3NggFGrDin/n8LvbeWVkG36mWUjreg0ac7
GQW2KXC2e+k4aWwFs6cRP1nROgciyC/wmOPKGIBjPhZ4eQAYBOQjgvvUCCe9ExMj7qR7U8om+fLi
ZPzU0ZCaSJljLQDuWYZX4crwPg1njFRO8wiotrO3OWLo4luY6iGT5gwbIkairUM4kjp0FfO1TYkL
b6EDQVKhOSgjlXLJhVyZkXrnVMoBfvh7WNXKfvZ9VsEBskncFc1mwkxB4G5qRQm40gZiGU9EE5EH
NIsi7o01zo+HY+28rQRaBi5O9jkXEt9d4067b7T0jDdWk+uuhguBpzor5DnMjb5IyfWyFpiOcmUX
KbcsajQwN1MhDbe1GNktQaaHxvDf+WeA4wXwiXydQtAy2/pJHpjhk9LvdAWvB4mxCFNRInsqpzfs
9tWUuZr6GJbabDU0gD06Z8fn1ihxI7FIsKZ7oL3pgRbV9TLH3EYxBep8eUbi993YoWN33O2szo2f
2vEGM9GuGGJGlHGrpq+TdWJ8W0oQ5hJDEC/O83Qm+Gtftd3i18qWdjV48xr/IFqCGRa0GEyzE+/i
tRbohzEQn2LqwNQ8BDIsIdkEh2aK06HiEHESdT0JhYxFzkRXf+0SbOJMYx66eumsPHgSzg5/NvEO
7gHVd5Ww4Re1OMv5KVqkzkfAZzeeUMFDN61DPk6k0f8RrlMT0tRMKi5qsuuIFZlMtQDpsIQjB9ba
34QvKFInwOM7w+RWqqr7nmYLx9wYeSzLCoZHZoYkYq6CbXVUgw/4EX5W3dk4hqUfUVZ5VdEHw9Ah
xTprFbTJkKZQzUSw6mm7GxHU8P/MaHXH1Fp9WZIMJOYfhiS07kIrHKDQWhjfhwmyX6+lva09lCMD
imF/mhut38fMAca5s632zb/UXRWMAqMz90QPej8vB+BWzp41fMyPXTzv+byl8H+qgMLHNb67tdrX
eHN8goqNgsqkWb+qR0VmA9uq5r6b4TxsPDljPq0qNP0gf5eBViNH7Fr25ycYG+xiR7d8pf4nlVFZ
Kq/G71qop7K7gmLs1tcaC08Ou0f9IXYUplmf3beJGCPbaIu5HbFCg1MIEX9xQuD0l7g4e2ZK8d/v
wT8S2IMeWLjt2MQKDCfXAH7Sv6zvuvxlBGYayMdK7W57elFyAnz0Z96Z1oK6lL+FVE/DO9KSodvv
QsaursPfPP3W0WEUJlV1cKRQrJGQ9otKf/CR+G6SZMHBePLhbxxO/JjYAxEbw9hxnd15EEwZyD0Y
Tr28enpDIh/C4PZBlT8EKRgrR34msWny5Cc7VeKbw4iNnqACT/ic71ZjMU86umxaAYsXjjDxU/2m
DHpwdrrCae8UviscxwFtLJ3Ix9tVr7ABV3F1xZJTPQ46ngA/OiO6Ub2dQQAIhUD6MIqC2gQ/9mS3
ecVw1qGuUGI1sg0NAEQiNOl5OideLL26bBR5JujC4Veuezk6d0jSA3W/5BSGtaWwo6SRowdZ2n1+
OkqtWJkN2zD/yccoxgznDLFu48MeLYEU1kuMXRy17HTdTNGdd4SXev4gDEyvu5vjSh1T8kftdLk1
dTZ6oRobtS73Jc24fEE/P3PNFLcekN/H8xElpsHJNb++Py+mYIYfhVJAMqxbzHJAt5BpC0aGt+GE
qDrH6hxlNXrJvcKTLDN4BlJlq7ZNyEcryuUD8lHuusP73qVJ7ErtraEZB2+LuCyVkow0bGc/Qo+s
9mKqSg6W3RGUAJ/4lpXKSD6h38JWtEsheKOo13Fv9h6ixHbqLZrfhjroxEswnwkOIzmzh35SGgU0
QuISrvnBF0LHC5mzij3JgX/lXnHk+IEENYk8ByYCiln6e3lcXTPwzuMa+OvV/KR4XYcV5mrcG8pM
EO6LZo/+WF7peb0NkCFcSrwGqI5lDF/f3KpkOtieQmJpNTI8/oRrbcgBAt+bgoCRo1MY7Ls5R/Ul
SOqev2eSRfD7gFHPJ1SBeuHmlZmDFr4O4k9trVNRiPwKAZw6QOrx6uPZ1FGnNBl9u6qiFLsr18rv
JwqDdAHZaSOzHNnKHOTjTp9R8Pa6rWN/mYd37V0HghQvVp8s+UVx+BH/mBODuPwv7MY+wSQo7VlE
0O7rmTYlI0ECFvl00JPbRtHTRBias7PXDAHSDIfLGzLIIGGgPD0jE6xpu/+VHsDY7/FUKuhlSP7K
QL36dAwIiXyp8RK/0fAFFKnNAG2NKYf+RSPgNAyM8c/UOXxdlHV8BGEKnOZmwDRj5ft8kPcYAmQT
FPMACLjwHVDHw3udp/dPV68oKo4zWqqGd9pMx1CweQVL2hC1CFDoUejqmyxEDCB8bJKHcDaw4LH6
o+IwUBNpNIJS4H8C1dip+wlRDY78wjyepGLk8qKGnK4IqmknceqLF3UCJIHzqbF5a9fvcJYajfZN
9tpk0R2JkGKboLDxi/wEynF6iGuLTmgxlfRjViPxExJ2sq9xXw1HfRYiW225pLoryca7l8ICHXBg
HIRVoMELu1RXBKF+80GxLJOOruiGjZjbawwCCV857bxeKvl4hAF2oRZxvH/Q/kO7b0dm4j9vdrq9
I6AZfx9Ns1JEeoM2u4qnVCaGaRl5kmCqFS35ycmd/Zj8VUT5ktHsBdKs25N9dY5+azOFmWraZIw/
aLMvveRWuH3CzMNqUMjIWnUG8GzXGkeo4UUe3J0TL6khBgpbFyFXHYwF5qHLR+ZdGCGwmfVbA8L7
Pm9RF1hvbrucvuJhiYzntFeqJ9rKuJ6Fb98E0ijMjQqVKpk+S4I2SHqEkeIzV+NYTpgTaAlhuAIW
f/kbY75SQsGGsVU9TViXBq9iJXU4p2AidnrkDmwrbZjnogDZkd7qPSQhzjvV/7TnIQ3U7e5PSmt8
P50BzqEY3a+hG3WFqMoyu2bfuLTysrUH+BFklWUZwH1DbsSpQVobbBu9J9RgfiPlol4rZgjHfxGA
Mqpg9NiTSnSmDpZOGI/F7UaBHpFtUMdP9Hv6iHgBR7bTJRMSzSqcZXoCGkXh9yVK4pJbdh3hI8dv
DvNTE2qTzYrdH786hHA8eHtmkPyhz3ZgzYO3v91QSEEVtcccO06+IDxKHCqY5EJlL2JLgbg7TrQI
dPW6tyCxpLkEGMXtOvnaR1Mdpa1vG2qjO6QpcKmOOpbn25Yq2Nb1lg9bf7E6f2hijiGlKAVDYwOx
/Y1IofbZttA7nphk0mZnyhUxCGQcS9ylWEqWMK+1JKP4WVsdbIwsmeOShYxBD1FlhkJPXW1KnsKE
d99vz+PxBkQdqNPZwl4LMNUuD67q272+zTc8/mR5xY7Zs+wy1RyCxuel+fBYaUhYNNQgmJgfvxSO
xseHVCtkbtgr00vUlCDuA4NPMo9FgN90VhVSYeBVi+LmiLe+3lBGqrhFSut45xJ7pZaxwAV5DLRg
YL/jYCdFk/Dyfhe567CLWBDT5JdvbKXlYv28VOnyf1iHiKKoL6pSPyKNK8W1+cOd8//zvLHAH88Q
VwFW2E5UoX+g2BxyZKoOqM0sr8g2EYpuaphP6S3t3f1SVglzYgyC6EoWGfRNN3lFWVRtRxH3OqbH
LCGcyEQVrMKjrebfn5MgN+IvIuZoepbD9IBI+lfcaRWD7N/2Gb1cpUgS2/abuaBfyWwAdIDFf1lV
l0vJ46qiNjcpebGaefjfzcOui4Kfij0DooeHrAYRmP8YGQsxcywmp+vrVlBajjb7lz1gVk5qV+E8
h0csyoCBSJStmCAGgJhqxoo2xkHuZ8SV5MH5pIN6Zb96uQ975cn3dOvAX3g1j9wh8aF0PlyQwtrt
N5hltV6mx4qNb3DECZrz1qoc4mMzXqrDk6wXgp+PhWHfAVqZH9am7RWp2cP+omE3oxuOed/TuoV6
iIcpNjDyXTpw+BI16Q2JdEtvXo6q/lgtxtgUZ+aBB/kIq4Nv5lKiKTeqKvE2X1MBHNGhmTlgjB88
gthiq4qw7H5Y6OyZU6WYyDaAgFzAbjhg4MG1dQNJcT6YwZmP6J77JJSIcZ16eh4pTS6mOSanXrY2
P+4FE244YNlkQoqq/pc+OWju0EtItPbBEE0PSxWnoNe3YfBsW3py3NzyjywSvMe97i5p1LVGLElU
jxiO1+eRz86HU4nAPz8LtnNbAXdQdyTiqRjapregNd7KcvBd+wojbuCGC8W/Y5Ilxp2r4vWS12LJ
V18bH9b9L7P6YN57zgnG5ySqzBJ00aTilu/niDwPboKtI4itWTYaac9iQgbLz2DRJm5LHDh2J0vD
eNdRKIaerFDZMIb08OX6j9MG24Tow+WEafDsck9fz4S4RS2qZaVedOzPnDoopA/zBbM0CvKWoDUb
Ph04BapP5rkdQfA3IjWTxwrOyibfQAs1dUaQ1UifyTI2AlsvVJIeYQHCpILg+L7aZ5jcDwIQ812w
f1J9JX6gKZZyJvMhWEX65KAKw+eq8m2XkVDK3zw4+PouK8vPXzBxawBu8t7BlszJXtYGETeRpn5o
514VwPtDDVQ+rv21P10Xxa79ELaKjhj06kXcSWy5zc+eCkyi1Q6vkRAr4VHPVd30rcz5ZpuSov0y
rjS9alm3ALNVjPIZR22VQWCeP48DfMUYagfU7zTm/OwXoEOML8nJnJqqV3OD10DqT1AhzMrSKCBM
/0XbvNhtPIBNRPDKh4t3jAt8RgiS00QOdoExMOuh94Y7hkFUOmfR+AlC9Gpj6WCHpk9aS++O0t9l
uguuy34ahfmqf/r9XPLKZ4pNluhdnMeut9fICccWzR1pXok0mo47LZD/3OwQUOL3yDH3HCWMQJcb
FJaiIqg7PuBp59GO272F8hORFAdRCyDfDrW2WOkk/LQdUF8FF1WwrihqVFClSG8sgoduseBZxYXE
gftqy+oY4Yrf9kVWWXrAjlqTngMwx5ycpXETwvufv9VnbFZc7MYQFn+wSjIQVKS8mhb41Yq+xRu0
58kfO7IwBXz3PnU4d0urpNTBP7uqlP8gRvhHKPk+VhA4mo/MjnKRu0KV6QpS1O20NamHolD1xTJx
lNbcSi02JJ+UrWdZ0aEPseIYDM96zAJRrJaG3O+WLnjS0/vMQsp3l4wQobL3ToAWDv8hbxBuqljw
gn0/DB1t3Am8zpsNSDkmPSgmfgw8jDHwjXRHYRcCb4ZuPdhUBrddYAffI2GJ5gscVN7pAJXBZNoh
FI5XCtXMgpUD2mvKvd57qA6GY0Fhd8nO6atWK2QQhE5H3eR0qu/mSPl1PiaXO8U6ycH4E00UlJcR
Vs3q17EmjAxnUAee4hwuNZOIe7+2p1rF82a74UNckzft2SUb5Xt8zwDXrPQ+ZV49Gld9HlZLszDC
OCPpGSyfwG1JjdtjX2LpFcNLojBv9R1cmTo8h2Vs/POYQqHgrMxJa1CnRtkPho+VjMJw7K8Y0XKN
gE6pmrG0QeMjR8hXi8N21/exiHK2g4qxaqvy0H+4jUkvfmLXVRIVPmuJoL99tNQP7mTpGoJJYYgi
R2Xtx4YZnRv0hXXFjgbmFeofNn+ieAAyQSc8tNT+7rIcnhRUvg9nWlwI+8h/FPPpz/tWOsF1GYiC
Qu1ALcnQcCd4+P2qVNxptMSuQAnudm80Qt4R8UuOCSgIzzuHJsI6UasjVcWhKWTC08iz7bHiGYZv
ZV7l+5F4pmsUFRJgf2a9wJnLbH1ceIo9xuWeykw1cIdwTfPIjXZOYwz5jJbWFUBO8nWX+VwCdtpI
uIUoY5phqE6883GSmJlhGWspKssPysq82YQgI5VRxAz4KUn2v4Vkkh6eYpFrNS1yl2IjQB40aw01
EWpVuaQbWWNTtBorjq/w66Nrihewm/cKWSFCD3SXSGIbONUSQw5qygL5jmngpAxNrwU5JvW+QCh5
Cly2lfa5sZIeRV3kNcukq+0wpClgGTCsQBuCoLT6XeIXGPK3s/C0oJzX2sy/hqNNXYbXDLH5lTJV
EJDdGGtG9yi+rvDrSMNkiI5LgkWJfDR7roBGoUeX277Sdi07bs7wlwRjTwMPkwWu+ePcGLF6AUH1
OetjowWVQ7hrJgNxFeJ+57vUhj9bX21qbDm11j6sf//jPxToYoctGdX5Yz4zYxiVWZ+suhJYRjiC
INkjvEuAjgjr0W0h9xpOFCuNUdnGlDi5B7/PD6PbCV0um36LN2mbuw6jBGpOdeL3Rrg+CpdjtxO7
ANZ/W0jNVi197yVN7uzHpzNCFmHqM5oCsisFI6rVjkW2zb1pPoEPJCjXYeKcdIYVtrfHPzBTUY4d
UkFvwPEzCNbT4BtzPP+h2qAR4d85IJ7fX1QRHAOQNh3UWncW8KglvLHU1cI29a5eROHQaUEek5Je
YsZzWE3wTpL9C1mtN8R005V87CP+Z0HKm57Y7OAjKzHJJqjpu536HRQXmYkCoJ7R/v7loiH9jm0B
aSMhlW+Xcyca80TPC1v8n6HJZjIj/Xx2OfHRxchRUJbVlaqaySHp4FCXHKyNEGFtYOfZ3tHzlDC1
/1mfyEWhSNBE+WmUEmuQutWc/ocmxLK3C3hXNTdUGzXjPMJuw7Ams1tZwVkjh7LC7m4SPGP6H+D2
vSeX80P/WHjcdjnUDBQebAltVQCAgr2HNKJpv2Hmubq/mj+jyACQI1a+x6diaBJYVoRV96e8BY2E
kY15dheJxdQlXauCpDnwX4JiFTirsow1a8hZz84vN9YvWNPc4SCjDya4spUNyIql9zylL+2ORPFa
y1TD1C8pFsg1g7zS2z4JiECiGVxTHEyHI0kySdV1teLgUG/vX3e4Qc2SCP/BdbSQSuUjhYSSkOhu
5ASpLyLe+sr839r2JkZgXGYuMEoMs611z6on0NVE4kbLkPlfsOII+KyJF8s9BbiGiW89Ne95E4fW
K+YqqFmFrKDXoKuHLcxBod5h5Rw9tKTSk0zQfw7wvcxESDECGJYB3D0i2ZmX8nY/qt2c/w9BWmma
F8M3cnVCbUBlQke5nskor4tUX6yGCahih5bW5XJkIJnt4hzz+syOWDZtEdLUlHAWR/+OkqVmj+LQ
I5Hie5r1679to0y0dlxcYADg654wAVgJgIYzTPsYfYXBs93dA+/Vq+or9B5AErADZTi8zx0RFHrx
iaDlmZGt7EDaRymgQN4wK8czRAT/tmeXiVneSTpRMfF2ddgy9aXGBznw6xMutNlECGtmm4p6rTab
TFkE+vRR1kpAeaEOoy+6OMDboFibHaB6aP/kOsoAWBgToBqcpLSyZKaCJK2OYw8c4pkvm3YGl8ek
k3keIcbs4HmVK3xCeXQ3ntStGpudoX0X5y7JcgB+bzXVyEwCvc2O2qp3j2APNSwMplB0FIijUEpo
59LBame3utmQ73bactpBoh9Km91YX+u9QT/foko64PV4DOJkDO+eKGXeOQukrGAp1AXaLUx/nyQj
MOue9Enc5hL0hnvQ3R/xkCfTPkaeTtqU5kB0FaG2yxJ4iqqXIE1PVt0eRBUpm44/6DrxzJRCwZIi
iH5wtiz87Ou+x354MZ1JrBxOG0HMN9BPxbtEicwR6Jpcti/Fc+wZmqxHxrPXurm8DlDMXK0MXZiN
JqJV2WEv1osdbu1VM9XWiU/y2zw2Tj0c3TNLdT0AE/7yXmtqjC9sxCcMD7ER/MiSSi5vGpB7RpD/
8aNUtDydFMnIghlKdNfxfxEw5NG62Falg1WKHTTJdY6Rn6iXjutnMr3lALvZKFg7gvuQMpQTV820
yiYvcIVE7AUnykGfUwHZBnGru76HK8taEe8MLk9ko9uVHTcN8r+vsNxpp04+IfmD1I1cCs2m1cd/
2FAgQ0wehPFb6JxJGyS0UXGdVAGLUr8GeDKUEzxu7WstybI0Ec7VX6CTCE3o55socAbLVyN1ZVa0
Brbi+oB31JZfBccHmED2GNSOtgirXLW6+Ar0Y3q7tmJm/I/TvrxZZ654re1Rx/9dtMXicA31kgqd
gPmEN7KpC626BIO6PkFbuiu6C5yX3LlngtvdJ0KrjAg1vjIt/FMDbCvqDGgzbkBpCtQ+rZjmERDp
e7FVDhSmmsQYbSpWxilFLcQ6+zyxSU7W9749jVmyMCtTpRXOUG8EAcngOV52dtpiLx/j2rMuZIao
RJxV4xI2bsPDkcLZRiCHdko4d7Zg4rV6AtnZrOZ3xKF9UpzVlX62Wb/ZRW0knoqvVC51GMhXf9de
r5qHKv0CrKwl7341kmY8fhvrBx/a/sVER4D+uPtv9iZXyXeitiTRkcgT3YwneR89Q4rXa8D9xoAy
jZ0lAbiemPyW/P9zUXe26fRFqKmD+FNtg1dS9b1l9dATMnkk3NZYnXAa80YcUTwCFmpnTZ7oa/OY
ebb0/14Y5DJTgvv5v/P2jiNiXz5NPvdBdwUhPL3LIGHXNAa3XdlfmMaE80LIY6M21BD+jd47xjxN
dXvpsgw0EGZzrtKjifvIJ5PBFiIK2j+OF45ak3FpD5ej4Ak1oFYisLOp4J3LWMFa/HJ8bDJ0im+f
po3TzapKlY/5YNe8yfK6kUMokSLMSze22C/VThFfbTDNOGwJG4rKzerRL0jgMAijuU3BFBpETYFN
005n5sHqzAe626JyCqCIk2It9btosoTqIbwNrzc7JbZKFRZYG/KaSDpdPwum5uio2nJKQ4JCXwop
60QGIkHrIQDCsDduS0IFwLqJbjcTXEw2PAUD6QappU0sxuhE5DX07vkP/JS0w/NQGUF7iiXuKrY+
ItJN22F7CgC9BnD46ehB2dFq2N88AiSMyvjlBtg19gAHXcO4MEaRohkeIkrGRGA/lB++JyTgFHV7
DfmN4ZWCAgFlWer3F2rmkYPqB/d5YHuh5FfUfosz75dEr/5ltSRVs5eaXsICcDHiQ9A2m85t2Kov
eyi55wDVr3NCWSJQTlaROrVYTmPzPuZD6AwUMteSG0bNFzpcO8DL7IsSJB/n0hvlKsK9ufb7yA4N
qaYPyUZ4jLfCpiDMX8xlL1pwABjcOzVQRl5amxsRMVu41tUxKph3NxeWs/oSHU28YPv/z/Nae6tT
FX+BjLDeBMEII0ZjOQaXKOebLB++boluoGRi5glot+h2uhrFK/KWT1fsI8++CRzFyLcFzxrzlCqL
QptieN0LDyQFzFNULOGb2FQYVspchspV89FgnDoJjY8jxucVX9RsvHNaP7o7z9whg5rk+PIAB67X
VmSF1vSb6uNOdVAvvi3TA0lVQqYGx8mqGV7CIFVzGxJ5jXxcBTj8SSimzUzECtC6HaG522+vRys8
ftey+5Z6uZRqD3YEnb4LLExJHU14UQ9IRi4YwjjvDmHEbMXCwUiQzVKjO/mP0rc2hLZTNOKvzy9G
JrXZhU/xboAB9WoCCnqVfqyOCXJCGul/GaYJhmfYXtgmDDQ5fbxbT4pQuC3wPo4q+h7jBVaH03qC
nVh3k25Ldz1HcHKhiE56gfR1z3sABSF8HgheMXWXhMd/eLC90XqkccOfzlMhOfpNppnA6WzcTh55
j1EmtJasrwIK8LsZrudqV6uRub3HKv13oXefUu6r+dXIf67tRTZqYWt1BB0IxAMOzRTYgb2A6+pG
oLOVBnFgCbgaL/1Rgssm8A5bpaDbe8rQiF8ClIOL104C46Cdb06Eh7okE1zJTZRsfigIHRWV/xa2
F3TAzd5I5jBsLp+abpMTaRl/VXqVkE2ejJEOk9M55tgro2Ku6a64d8gNzhTaKaXoNAqW3V/AHBn9
SFaMENpoTJ3KBkTpv74r6pBhUlUy73idevyVPbo7Z39wH+Kdz+psPSfAVAHLPEpTgJQKhAQwRKHq
7874S93fc1JAQAHGuL3CD4WCufGW8YHm1CgckOicQbKftrjSWM16d3QjdqmNqEckbbe/Ur2y6gwX
jzOE0QroA8UKCyC+Azvj9AjkM7xrLiiWkFa+mBQXBqvxHrEByM6+obMPVfCmouoZC4AGnFrCM1l0
BerLZctjXi/btYbxDCXfeVAAMAOiq2aBsEoz+BDdkpZtNvrCOqcoFuijEy7FTmqYRcdQtoG0XUp8
USE/yestNxY/atlZV61eL+DBDXJDmsNyPxZscyywm7Kgfhu1VNZAu9JO0HORgkLCmXO/s0He9tE3
UZpCqucdapv3PgeW3f+RlAUetp3H6mdf1J8y10JIMsrAEkAHi0BP+4BbxXMOU9HwbOWf3sxNuU/J
g3HZWSJjk3tRr56e2dm4y5ccFeA9dAeC87tqS495kvD6hd9hn+qCZm0C+EOz3C1zkho7HNfpWahB
owisL55LUNi6hFblRMdCOEsOIDPtq2eEwMTuav5Woa0613khDpr9uuFaZeZ8m7+MWXlWuo23TIQo
cJKvXdSQ3+vxaGaDtirQSg2B9ahTtdNmqfg01SQang266vWC1qiZxkWG61rsZDl9Y2Mt9C8zEr2Y
gLVlz4aaV22xxUZaTlwa7vGet5StxvohDc+rJ6RaWwPgOR3FfMiQnHb0Y/rsWZDVsbI8KQAWlKxh
cDCFZlf5goMu8eK2Hl8a4/aUzxF1ATOxFrTNvBfqdh2pu5i0X5WnoDgEjUzw72m6Oy7FAjmd/UDg
6gdqKqPRBBgT1KtqJqEqeApqR+qH/tj42b6NKwHvuk1L9qloLXmI+dFP717nc8yCcqQasBCGiuF2
TJgHwOI1oFesj4W8MI1y4mNcoHZxHeM4SRPHJmqe2Nus563MIh8h3mASvgVOeDNLpgkx7gDfVh1n
utIQiTu4ZNvoPRu9zRR10Kg6fzgrzrfOcITdZl6eiYAEozosXSwDk6F1/Ts2CayyFGpmZpZw63OI
uxYrJrEv0RaOAbF1g3P+w20VZQS4Fg44rWxnHoZ6G0l41q8tqaJ8+MUNJIaVagA7v+nUwJ9/azzK
YIys38ftZcfF64bXN4tEX8a2voLw5rTVd4UEE3dhNSCN2IpgFPXoGVbVxLoxMFFJ9NXf+Aj/db+l
9yA3HlvD0RW1eWIAG+mKd85PPFRc7AgG+VoqtJz0w7SUxFYVARZoJu34Vx6lpwiBmOoPt2sI8bjj
St2xyj4PSM47SFmvixcOI03APaHOP0D4XaBJQ5U0z6HO0OZjxcMFkNz6szyuj+m0xlQkbEKHNvkA
CHCJIHozvflciBUqi95Cq9Vvw5YtSCgzDXPSdeT+tyANXHNtuhdeVXsp/2nnjHKjMaKT0yCAaYre
uxxCBihLztRSBsTNtLFSvIGxNK1u1GTqhF8Ks69b0IXcnOGCtQ5119rhwRuXTvDKGpIqgin2D0gl
ze3QFdHj7Rq1Hqj6C7k1rSOP2hRs4jEEBf4oXMXdLn2s+nGeoZd3s0VGt2yEHE4z7bDYuOkHIfBh
ZsZC6jUHqQXfaHbFrybyfqCVlAjG9LSJkgtoZVgzVHKspedRfGjTnhUckpC3H82NPIyV2BAWUL8T
C3haaFplLpS1bP2tgsrdlc9F2CakUsD524sG/P+SoGF1krJL4ovJG4MhmTd7uaqwPWJGctIpskby
BzHeejIyO0d7YF2HJQ7zZltzKz/MhH/VQNsxnbBLBU6jmB3qpIxAnL39h6Vnz+h9NW3e/w3QmIm6
fSnDwXTRL66Rml5P0Qx/6sylSzxqptdr5KMkt002pWlALSSij61LV3Adhor/v7HxxE4yUSwlQnuY
bKNe/IKH3zObIku8n6D9GI9XHcLtsVWwuOzo4jIP58Mucx4iiFaC++tl2rRSrvHA4Sg3vjRW2Nev
qQOzrf0GM6bMjsQSZUk1DK1Y3zO39bdiHe9S0nEsTIBaOMlbqtGU/xow1tN1+45af0fzrzqbGle/
UTXd9Yg8CBqqSFdNuY3xENk/IVtLIjnAmXl+LjfcrtuhSDy7o44bg2ZCC6bE7iV7h8OfV4IfwraF
AmPo3LSJNjS/hSlPvbl5cLH8sGyHtKdmzYRMfgeS7Ya32nf0Dl/S0EZvY3PVaQywvxxrsIoxUFqL
+qsZilC7NxEdIgEPHNog1Y/haN32nyw3ZsSMYkCa5VbGb4NH3DnL/X2TcOgZA0ciqhUOtt+tmU93
qEMunOkru5ijkdO+/UlTtZWNd/qpy7/qPMZQ+w6po0rWmN0A/+97CnzghfElS2FKxjDW2+NyVQta
X8XajxlXjrvcUPksNnEcdA9FWFz6ICnf9V/xhFvtUzHNZDtuIonwgZPvlyLplx+YYXPvS7uXfMfn
fRS6CHT/MuOgPj12CtUNWuTEmJK8DqcgIVjbTlUrOqW+tQeGLMR4e7K5E2ns0gpJmY11jJiokxYv
0RsCrSYETbEw+c5o/ITPLO+z8sRBohVvPPfObQNmYBR7el7bsrC54gmyhtnkkVUUhl5M0gsEv/qM
bgjhnQBwBNC2s4uMhWpgraAeIRmwf7ab7dVNVSH/hIx9L2FNoS3AxpxBPLetppepBtBwLncW0ZVS
qb/L7gyRMj3d3D/uhzFMbcHfh9IdGr4OxtJdhohaNzQly+yFeVXaz9FedQdpvLIHVarN/pdPY4bn
AheFdoj7K/pgji5bhLd9Jxw4kZmShq9sGnvstizEZQ0i3eZkjfkHl5xe9doQN+CORnZDE6kk3Ybf
FDsAB9nkevLe8vakKzTiU+jVe/7CFSmQBuZ4t7uL6khF84cFGKaUShirRny8KWb2NzF3IajnVOsf
RnNJGjChdstT801uYOHbD799vLPYU9AAVvNpHRb5OV8Dt6Dn9cKvqab1Kkbr3+sle1+cBgILejei
gT71agsQ2A+Tp9z6Tkh5oDCVsFNkTtpY40pKF9hwabUmzXbglIYWKuGf+TkBclQ/tqX3ej6LZXJw
5MAE0JGK8Xt39ohs5lB3KAjohYSdlj6qnMMgEagarRR+0RiZ/Jr98AKnY5hnfCDbndnmoTW7iD9i
fh5RFkm+iIEI0iawXajnMVHs/l8E+rr5QA0bn0w3OwwPd4nfoTYmd9FCD0zXTEQ32SwuxktW6VCq
62q5UuzPoJWim3mESkbrx0ZIvrd9+BmGwX9tuLZ+zshNmobgbnJcm314GZm0fyVuLlGUCblZtfUE
I38Ie+OqH8w/u4OXvJtOseu+KOWIUwT52ENVfS8D/5WslYzL+T6d6IGr7Oa4GsHZi0uO/lOUftnw
d1tWdOuc0ZRNKPchbWzJ6eIhEaHcDx9PxATlYQWNER5nj9428MzDLe094NVGsBSp60E9VBtvbjSl
PRA9XJVomnpr/kW0CD672KuCh6+aVbHWJLqmCAzovGBwU4OXRanGcPzl1wzdGSw7sjQT/v+cllZI
scOaCYzNTbGpU31uQCHpQG4rWFlsZxskyMmJfmegobHaLXrA0Nq6qNc/zwx6SV57MjhtKA5gMrzL
Df/SLkubmM17M1Y5NCCh2SI2Eq/F+tG47MMZ8EZIaPk/DsO0sBim2SRVX7qvhfxYW+ReYJg1psJG
iRhfjeR52pQkysuW+8Ate0NLzWeuwnGQ+xvMQKklEXBuHz1f/pozotsM2HXnIXWAqTeomB+3aFtX
mcLz7ljI6Te56DcrXZQMDEO+LTnf04Dv0vcTIHa6GF3Pqvv8glVfNrL3dhQO6X4WvdMI9N/SwGct
nAU40InJbTVucriqxmOmgPuJ9XEgbDNFX/t0YJw2s9hDG6/fBfjQxlR88W8ctd07ZOZfs6J2L4Tu
RuynXnkt56FRWHzsneD4Lx07k4/anT1ACFeHwbYkHEVNv9AfRGH3ykjMZGrK48xXwSeCOLK3yX6v
rEr1UKPg3H7OVIU+P2BPq4mdI9K9lhCYv0Ls5PH9X3HUTI3GBT6SkyGoTOfb48O27PqvCWx1fDrA
OKLJFCoK4OH9C/5psLBqkyZ7NcJah5yxsz0cdZhBgWO2BC1H10LHCVTr+Mfv71hBEEnHYHeiPHav
bjovbEXnX9DNb+JQPi3IH0iFHw4/o1MdKynPdffb5YEKyGqGV3prJTjRau1pPkv1E0MMnsjM2rL/
4sP2bPXC3WDT2ScuFunQBJzbAvt65Yb6nI2vpJvULHagaRthz/UWj+gbc1ZuMeMfhbohopnWywPm
3AqWKuZcaCDKdciqMneG9B52wsgPd96gLrcwzc0pByU148+FEcUCSwnFgcCBtFnnbs5w4XoCKCTS
cQ6McIlV9a2czF4G05M2EDAokGL9ZZ/ksbR4l9AoeVJNU8OMS7TRvhyXnbwkq4xnH695qvKaBgPp
Kcz74vkuLcwr6SN7HwPiIuZOZctdqCGYWbKCUtYtbBItvQ+skmmvsTreCAZMfFwBto22G5eJik5C
ESmIpSsHavP1ByuHdo8hWX4H6kztOw9lmSnF6zTMoHs2uXHnLalcvUHSaofSkJdE2ofIgkYDtwnK
pL7yZFvaDkOJBYmre3/Zy3dGNueuMtqwEsPIhJcRMex3P+gI2xAEVx63Z36A1YnVDos7YiXfBm3W
Q8iXz4vU7z2i1+DkNLwOAzoQUuJNnCuIwcLddYQvzN+rHiinrVcAgkB1ObwPYvvrsO6xK15o1lNH
QSwrslL0FVFE7jLXCxQRxrq9w2MYaojnDm2aj8S5jJOIDx5stUKA+dOo6whvcccXLYSqc4jGOl7t
a5yDWzeb1IcbtxF7rEg2xXAJPPKtIj+X4f72POn6vd6DbVvC8DOg21uryxRJrGQcdMjz0bMgPpfb
nXA3ZMdqa5R4FrvLbj8IDF2DilqhkaoLSbLs4Yil7nXBlBkI2mw9yP9S7iaKI8OhMhRSF6+/6at+
S3JP2PpTPhF+u8kVxqDUWnd3llBkDlCzNmgnkPPu+NwWysKAubdtAWG5F0aYpfTZg6OWw/Z95m/Z
EIcni09/pnHr5kmWhfzuCFBjnsezfAV6SHR9GSuoMI9cbqAC7B1hdNT6NYNot10E23zm1JTfz0aX
OQcoL3H+yhrhnf4qsZXa1g4bddm9TrW3DbY68OINQNGkR3HMXw+jW6nubxjFRFdowm+cwnwjX2ff
wZJ/TIyCjejHuAItrzkwxu6vt+WZVtTC0UjV2L1yY/6mwRTfItGLoW+qZTtimCY6ZV5EYpXzRFWn
2Lt0pMufrvf7AbYEKTkwa+p92xLjIPmGhdg31HBs6g1sGUZDzeiyE2+0T8R5U682eNeEALdHGkrH
KdCpPCSgomsCOr0jfuXUe2vCeh10vz19kIhgHeyT7Uf2pW3QUbWYvvtaKuDKpn5JaQPF912kluz1
/ld5ZrKsAFJId3qInUROlJ6gTGhfyO3R1ut+iR4/GL8FDl0IcI9QAYPCkiBHM8RYf0gpqIoVcpnj
gDn1xv2wak8tVQd0kMsFh2uEGDlyiBDrSP+paspRH7HpzZ2GvB69MaYQ96rgUr/6mK2lQsUiBROb
1l2yx8aOnzpg4MNZWyvU8MNn9PwZ3Qo7nIpwrNx5nwzZK2Q3Nr4BG+CetWEUvzmXzfJR+hsucA7e
G28gATzRhl3JdFlMlIQj14UTMQxBeWLlYaQhlBwdpCxOjgLqN5Li74+VkCGlqsFxjekMp08Mm/VW
/ISXRQu33Mk2v9ZzSb8cgfRtwjCKDtD5ZR3yEKoqQqHMK7PTiDOsT2Pb5U8ljAsa8sg1lYUlIyny
w3oYOhBAlg+wWnX7ow120tU81z74SfdSxrAtGN+CpRgKYph3H3VTCIulooKWZ0ufMsplijZQCgag
8vtV1NqJI3z667x3l0klbpASee3oPeGBBLYBUC4gv28vMYuNM7Wcij0Qia70Kaieu0Et0jrNUSSJ
8nAZteS4rHxMDN0YVsmxDpk/pz+0H/NWg4BGzZ5komNHPKVs1bCI1aO+HXiixvCstjq6jmc07tbL
lfAglsYUnGakimzUCPpiADIglgpv7jZ38E6fszYf9/fhBBrZLUliNOAz2mhL0nd/YS8gd2SX807c
mwBpZL//ff6yVPurbMfNjGSYZGeq7SFyYk+jqs3OuJpfQXGaP/O/FttW86+k7dZCNm2RoIjuISna
AEQbdhog+ENJHOCTKv+JMTLqS7yqYgu/vB7QNkl3ylR+7DjIbIFdUcp6AvcUuIk/bqdGmxMeaAlf
C6E13n76MECFCMhUh2KvAq16eRaMo1UeYx+kqMHvGT3lNYKj+wSdVIXwW1/Ce6titzGKeF3v401F
Ocxl+agROFZkKjyK477l+M7OHblKi5BRAK7UUWsFn1eCgJOWQE4siic+MBWt3smcGEiXvSdQcOQF
MiMkJumcgkCs78S0niftQ1FM6mE0z4BXrNnR9T3ycwDL+eN5b0jmSh4mc+n4auzf28tG10eUsKcY
zyFbgATFSOEBE/VniA3Yk41AY0A+K/pnrJ7GMjI/kbnx5axeSi6KFPAOvJeFisdYzaFy0+OPcNpf
pu+DMfDhmbscP42pT50/IhJ8eHgZzDTOjdw5C+68lfyiguBgWh3Nk2jI4oELU9a8P9RIVxS20MaB
MVm2+p7qiH9ZQ9H/lD3FXi8tuxDairy+k8O+2yhRyOzRd8ixn05jG5tcaehxRKWMVfjtydmL+xZ7
N4WpC0zRRxKWyKsXUmIt+llADZstLwyB9g52HLP6qkaWeHeMcm8H5/0j4LoA4LCdxjW/rrMd6q1N
XMt0JFVxwoUGHXO3Cqg2AZ+9h5mxW2PU8f94VY23alpoNoIXE8l0AZIIgvXbxrXC3p0RxolKUqor
PL2HXKUXGYQjA4JnQrTjg93cYwwcVpYBDFBvlxvfHaD8BBDuNzBq/Z3uPm2HqEWs8F2PtMsqPf75
wCjW1zDAa/v6ny3GSnZMsx8UEBRySwVa5tI/4qYMyD5X0S4+XYexlOWA5Y9sJJE3UxDM9L9AdpZd
ukv8m+15ar3zoIotSf+prDmxrjPacXrMqAogg1bSJNCxvgSJFc9lJyah/sErEP3CBXrJK2bojdqh
fBZ/FQpnQbhvLHgcQDTTWprVF2hmGtJ5XYxK3srHuwYluq6B8KW4XKsvyo5ootS7vzwy5CMOuqoN
W4JnMI7FRd3edmmBRHzwE+HmHwdMGt64erwUzCsj6oUrlWv5zyHLcyrLEFroePNBv+aeugP1uBE0
tGjF2DqDsVJ1DmSceDofyU+eGnQZF+Z5Uqa5whBDQm8LRsBuhrwAasqE9BrhFLn1jDgX7iWx4+Sf
ADhusd6QaPmj1gPJqDWkZdpUV28Hfe4PgFzkfnM7iJ6FOnLwAFRvZTjzHBxxTW61sNIDYUbEqz6+
enfsvaH53TvR4EBFY8d7Uthyzg1CBE23iFYl0n21WTOH2KuvsomZ34vzuWLu8LPg1ySLpUycoiGx
MPwLnBsaCVSY0LO6w097V7qrdURNQ9EzjxdUEChayrNZtDb3jPTI/8Prdt3roa/nH01kTBm/NTav
bw+E2lh0w8kShxIqdbWYux2D1blTStzgqz9yhFscSahuuSfwdzUiqT2UHI41EM+pFztdgRaOmv1n
tmq2ihMaCIy37xBVbiMbOWFlBgIsNjPjCnJLgm0f3pQ0MhSjtyWEt8HANLJVQ9kaXIm/YkNCaM0p
CJLivLVyGs2+sWXbN4gshZXi7wC80s3EAvR9SQGx1iYXwA1xVuyIzaXDEZWNOXCbXidFRxBUW1WI
AWrr4V8L79wkgp+ahK7KjaBYTTVnrZrfmNMO2kQNRLjRLm/wbrr09SbE87hVDBGTG/x6Ud6whMb3
l5dP63n956s1mGg0P87VdYD92OcuBgsOxACWlrrfNfQ0tCz7Nt2hdnSeLdIMAqpORcuxSAIhUqW1
laTSGiWr9C412ZHZVNhuOSrKflcRNlfUJ3fC3cHSTYRK77pZhSlC+DPIMBrnaGC/kflr4Frf8AB6
5r3/QBPaCK/jZ0PySBMnG4IicSJUwCM4rbCqgI6tdthPokW3/JbfOGHOLEOs0n0t8hcbVlOUfA6T
mMX5lynM+aKObb9jfWWLJ5muRUgFiXAiZNCap9xJA+/l98a/F0bZRq3OC+CA+5FXtTff6BBX13bp
7lkCLBZJVt2IMkH0E336hn+AvEGWgFljJUX7KF8ktRfJRmCeORZCHNOiLtr/qqlWSL+ejW4DZrQI
2b9lERlNgMqbgDBuX1j0/uXvd+pAQvaQ+A6JrVz8KFyhrKrOGumGQp7Ez81fjM1NcKkHT2VI7oJ+
RepmAljzOXDVbuf3f2dDSsfYYDBTzn3XzJAJLQex6G4eEkHPKL63gfy9BNEX/cReMieGxRZGdDMd
FVLLY8SuibEpsM2dI5xqudnxuFyyr/1huo3SaKkJqZZTaHcKt2aMfDY1PR6x5KHxLbKnbF5Bx3Sg
FTpsvH7T49ksreCqNmZezN0qc4zHMG3+1WcD6iWF3W3dF6W+5TdqDxzF9xlg5rDd2/rP20CHr4MR
xO0A6DXzsClzXaKq2wRZleIiXERLK4HeczFhZEtzrcddGQaVF8zh13pOYE66eVtD3u2hD9XiC/Wj
tzD3OhMlDUUY2C5MlV/ZL4tL2faLzyeGCADIlUptLLA1qIIvBReqE0yGnLiyXZufcJnbT5aVn1GX
K/aRpwT3H0OPsW+3dUvPT4C8pai9O4dd4p1pNjc6/qsXOewvoVb6XeqRBpp9eDa0LLLfYAHWoM/L
1O78JKGW9lJWvSOAy2m/qR2j9VCOOQXefSUfbSNqKTUbEMpTB+p7Zu0SHCaKg+jurigArtJy0DRX
U6wLXLvnc+JYhxlDfYJHq6fWeIiAZBIj2iBCasoGbQ/D4DwUSfm4rDToX0CcHBoDTRtQKmOl8glt
BxoKFPrzouziSpwIp7uzMPumUTMbfNneLAFNIrqfDLVKT1t5W91zycq88fYuvW6BfQsaMhunCJe5
Vd/2FWQzVeNXDeR6cVcPIi+bzI0aITpaqtAW2foqIUCjQmLHgMHYaPGcOwtnFo4+RN3xr3YcZgjh
eN5FgnY0sag4oi8RLnL+7fIPxoE1Z2PJcwxfoq9EGOMwEW6aahYuybR6dMucuBJ3fr+mh3lcNNlE
Pr36+OcGT1AAx266f7+eeJF1ECdIA0A62fmBZE8G2Km48nqR+c0SANueBGn5ubGKk/qpIB85FG8K
y4pz4d4+lvNcY01Tye9xpNZ3u0Y+EQLcz4st8cLJ6JX/EzqM4hlAoaAXWI35yR/hmKgwOcu1BWKN
YEw984E0J+yaFLWSplZLrv5BrTEcq2BDJiiaVwHJ/izlE4lyAPkOPKGReRHpuVOcQZydBjkNthlX
SWS6OKz6S3rEVkNmNCzNeoMcX4YmRMytx1/hH4F7n3bN8R5eSUbXoxmBUQ+6DKHErJQA459/h+c7
khqGxtkerm0NkjvxUbYMCyn8VQ9lIGs+ri8CM7OKyBV1J+Rqz9vdylqC0HlHijHj7kUHJcdRLfCe
+DKHaJLDXxqx3l3AFjtvJaNu4wQtFvMkCf+zPjX6mVcmKtik4MhQr1a7fs7hE3BEvPHfdnK9Ec9p
S7seVnXXtCs/Rz5Nm5m6sZcst16yRHo2Xg+i2j0AE7tnzsKobM1NRiGheHZ0pzJovfbzYYC4U+FJ
8wicsOCMW+xjkbBhNRX9INjJ0kkqkyQ5Yr/j1TGWE7TSxIG+LrG+ixTlUiDbF9eFRzde4Bw9SMHJ
Bv5ofb53H502dmNcQa5BjoFP9Im/NcTHoTvYHuEBN2V1cNdCGppNRHHU+QVc9X4LeZ6gcT0lR1PF
h9Ne2yKwp5FJauN97WNhSPpvnNUhhZy2K/RO4FexlNWkmjuaGTt5bbnP0PK+oiPEaZdj4wE8d6bs
f19TFseSkfnbMl0bqTz0yBHMoAnXid1SoVhZ7DEM6UDpzSIcB4Ghwlq2yng4qw+qolctidD8xI5m
ntG+nwi/S1YzwrQSMB/IFv60eURvFlEGzIqMQueDVZ6qWJQiv5ieQ1tCQz1O3+kc4sWKflllRv9B
o6MPgJTuS0G9fgp8epKjyM4/7rVVZq86m8QM/UG8Vcg4dT8AjvB4RsRQEPa8bcwSUFJS/UaVY210
qxGrQ/BzmLqHROR0lYvx1P1CpwIOF16p3yVf0P1ngC/L+cighe6eaDciCEe1Chttu1hEL36wSsHB
eoT5E+Wd0Iua+giuY4+ZwUwB/DF3ZL6Wk3WsqgBOPHoNf+cCRNuBnnWqb+R71xmbK5lZtGe/iTPa
FKla51pEpks//K8QoUZYpmwexPKHxI28wnR2U11yZD5q+xuJoeQOcHydn5E9ssjn6j8TcjLb2G50
dEgXFZHAxagGGB6RK7WJ9SM6tA4lnCenr2+1p/xHrK4eOCiPCePqNx0oNu9TnPiPgye3P91vMoAU
XMwkOYJ5thVmKa8HrEWxJ/PD6FIx5k8pSGdEnzUZ2ARPDtVRMY4QsARjPOReWgNh0g5Tz7RsPxZC
pbzM+9+Nf4y72oDS7WJ+f2u9IK6X9OfxT881DHP76l5O60f0UjN7oTSD3dsUxj/9HeelT+LDZeYG
gdDCkoJxWPz+UoUu0GPDAPiXIVqMlSUAu8YiKRtJDkmxANMLMbbm080DfhqigqwoxN4sFkOPjRgW
rPbmBMMkfD3ATvOgvC3ATdLDKhXrcxLUXuKP0Vs1OASaAzrlySAX1kgx7wwAEYxLPN2EsAtHVl+8
Gv2bTQQq780wH/kzWT4UvsqEE3b15HzqD7mXDADjSyCIgeP/8xqGok1p9noYc3KLVlsID55YT0f8
spRZC0816VdBEj4B4z924/WjAVLu51ZP0KTkKMqJVwWDPXx3E0/OkDwd7wOXalZ1QqMx7A1BlNXn
T+xxHJOq4hTuuknWDl3H/o8LxITztELcipuLRW8H1EBZIej/tvWfOwnaS8N2sVYB4du/X+9UsdUT
R8bxG00gJm42PMAwcgC9mcCOfyHKiYzRxMxOG4h6/YLyrgQPEostioKd+X8/7/ZvDRFnnimGGbjq
dkUnJkFuPTKbF0kb31+uEi0zjOYXyJn80U8UHiYQ/VnZHZIqTJYnKVoRCT75BL5KuO2Z+CwWlBOi
gDynhmFutiyKqFwVLc6ZYruF7G5ql2u9QFkOC0nMEPL0QpEuxO3/EmXLI/JGfvxEo9SDtrXmFCed
nG31E6GwSTltHd5n+TTqIfu3LRpP3qvyCRwhcBVXW2Wy+6OIHqwVRE1izqOTrfYhBUVd9z7oev33
A8LPtRvg9HsMNSB+2Y4ADRAg9vcExcYDJ8Rk2Q1WEkcv9bdlGTXCgKYswk8gLbI24BHjBC3PnMPm
3I7XggjG8XjLR8h1D3WnogfUgBbPrW61AU1a2VpA+pO8LenEKL2SObNni/WfPs6kXNYzpDyInIuq
urea1P3BQuDZ/tbrXWuC7k9TvMN4h6kfRjPN8l6LpxuWdZnOrx/PavtYEl44bZKExXN1Et5xLlzW
Ur4KtDisxEvtDc0d8Et88ufQNi2MdyMWjUrA9kVVeuLGw12PEGSDPUmDVJmOCI43Xf1abm7U+/Sn
h8XnCJr3Ulzy6BMXzS3BGI0my5SquxhM6uWKWD9PNnUmSl36nyms65WGWE+0LKmaSVjVaeB7sXLo
M5GpYOfYwGIUGYYzSMqTl+6LnmjxMjaCDPv7fEdkfq7aatPHL7mSYwxXrtY7su/ZhuD/IhK+Efcq
vFkZmzFOYuVc/j38w2G8QfmNzClu/0z9YyYOxCpmFXhTlJZi9jFkV28V6Dv21n4jev8cG6WAeS6N
IPX0Ftfqa6itTW24kbJXvprf+r0JFa4EsIxnagpGX1jVtlMZHGYc0ZSxA+2SFw6UHIMOzrbMp6Nb
eGcvhQN7hK2JhRRrWP3MeM0s5XWqby063nQHE2MKEIolNc38eCTrxcEsZGseFjHvjJHK1X1QBowY
bKOnp+SQBNn2P+J83nTYnkzDdaRoR/kuuN1PP+ckbcNOA19ZhulFuQZAxuvsxMpF5vKbVPvgzgrj
FCPAhbjc1WBC6g4SqIqZP/ZeAIzUSUo/DnOBWyOlR61vXBD+40k7YxRPO8fuKbU0cJpnGuIPl33t
0plMcIVIfqD41eKBK5XjttlT4OCjIdKlhzX+6JIBv+e0VuKjhDekXGTkPpxpJv2At0jzKlaOJJ8D
Od3F6mPE8BcD1Dg5/no2AZF4Sm4Ftxk0UkkO1YrH+Wnjs1GCRYAt5YCmKTmLCOTtAI76vdWEjgjj
E2w1c8kNAmXlS7uMmiKnJ8+MHjzxaRIcla5W43f/JUjySJz3bPp6nolECg9ZjWDnvQlEsMxUiyKN
TOiS0daRkrXKFk2378OwGSChYg7JC20BIENikPhbCF0IZEUt2+xJXj6zoX2UtUsgJQ44pt2JacyA
W1SqYkeEmjVbLtWxgYWdpg8/q8KP5stOnidmW/uHJskhFKm0WqDcqDCBLqeEU9QZSAagtHhIO9vh
GdTerYN6Hlw2WgqlevM/6iH2CWe5CCbReb53zbrm61A2zAp8jesbZ//qT+eYkraHotmRE/K7npZg
QNFdW+bTAncuXLoOU1X/xO6FOQwi//OLblwf9TsRjLW1K94ifz0HHX+dLCb9LS/W1VeeYsHW4ATZ
h5VI0L0oOyZeKZjRWSAkGEUp9JvZFPfjnAoOrO3VVqv3dSSNl+4AJAR9wJGva2qhYmBR0HZtdIgQ
V4CpyX3nlLxl7Vhvv15gVUN5eNeAjQV+SGP+6n2wm3wxZgGFleMwF057lnRMfQhSjsViT/NT9gEp
Ea/9b/NiD1hAADP9I2CUE8ED3S1p43X7S30fRNDquy44ssvPpOG0ZrvcgZPb9oCYUxoGtBKAFGO2
VXrCbMRyolSxBBT8B6z8oTYsYI9dIOsIKPC8FIEJfAScCLKPY/sWO1UX6X8XnKBfkO5ucQM9tCwB
0PZ4kkH1EPXuvDs+miTjfy58TX0rMrj+WqLGOC7YRPTkaWdjZ0f8vEbWMnmFHSs4AWfhj+dMAbmT
qqgzrDQ/7kBUTp0m3UG9zhH7nP9MZ9sUTuQu6H6wp+0Ue+TJaQ2gxQNWzACJnz738s+7YIFJU41a
0wwAWxNSMGrpClU3iUxy2A3ULiSoP5PNH9uGJBnwXUJKYv77MYnGgbqEvyV1hJsnISfENTYs4LuU
XYFmpR43Kx6WcS1QzFgk9+u6Bn9I8gbnFawI643coXZxtGCNPavVf2cXxoW2R59hW0wrJ/efY784
PqQ8ntMM5ShBP4j/J4GLgmt+HTBIfh8BbXisuOqIlIYEISr9HfhiCqRPvyGhlDyOgJlGnff6LXXa
j3XbTMt3iVxQfsck0gZDceudeia53Cr3MEAX3g107OAts3oI8XNj2IDT9MryMUR8jH2Ee0VaUrkq
ZXivRL+Ply674YUYV4i8Wr3J58fEkSiU2MIbKLLdIS3pMwlTogDbZ3XnQa4qsLBIfF7VA1MgczOI
QOD02twdu7MaWniAvcNE7aEx2cssgpom2P3AFR49bIdNrrAKbrFk3YZ1x4UoFzsZ83C0Cu4ywZP/
ic+plFkaBMv7s1LoIbLc4MKHvQyLipUfYIDLW/Q+jH5p0GgHqvb8Fkdym/SnekKnf1STGsW/AWAz
juLO15Wfhm6khUBMMkBPekwPcfjfos4pD8hhd4WhDmBY4XXprzqASpVMNazkwOK51LAD146BujwQ
L4grVG/UQw6TNI1KnJ3tmhfv6y57rK/CubBEPIbIDax9Q+YTc/ziJiqOWa+HcXtwu1kEj4/ikfPm
lTOSu50D6KAZH4qckmliC4/5BCn4Ht6zL9XywGSb83C2fdszP/vuweO7+Tr4NrAvMypr/SLD4S0M
1kS/nnPbi5Fw9S3UFzgKQ22/qOSn6exEFhEW71BZpYe2H1ToRodBOBk6mvBFUftG1p88LI2uKf1w
2WGJvbKdO6G6cLYciNjTOzWXztf8UWOSBw3k+aqEQrVFmEm3AYj+bhKAUmVzd+g5CJGTO2lPZQu+
sUcO/Pv0ldyxcDI5rdr+XJX9dPZSLZlygKfSu6nPzd18FYPfG90vtmEqvYdZtvAIQ6Xfm5k6RKBF
FUQgOgDcWNyPOjGcdyLJw+VWLA0XcPxsPFifRcOdfl1cvSEj6V+PU400825yPJnqyUurI4Gz1fr0
9jUb6IAFSyzzN/EU7sw8+KVmNhOpt53qeI8cKmbtZBWEWcGrfGLbu8syCSIXQIT7FopRVJoydM/R
dvh7TqEZuUhua+BNViRVplm+a8zlx15HRpoTVq6Nwj4WZpuiiHV1fNrYmGJZ4EEBwZbVA/8I7e10
eCkHY7GyOrLF9fL5WVKTM6loJ6+44UT+1rxMfmRl0PWdpW4+Mxg6mhUVThIpNJJhnMA2UEBIJb8p
b0QRWW0Bd7CxXWzBqylfFGm6UYABeq/dRxQW/IIeWp183eJ5znQGVH1dVZJ12kmTiOczOk/EsgaM
vonPrYzMrR6hsOk6XlQMaPzXROsXETFZyRnU2ett/7lrqIe9WCVTWbCMj0IzRFMiEqVY0C1/IYUF
ZdXom+VeJ7M8ApF/zm4aBWP1yXVg8y14kIOdh+GIzVderICPDaCmRrNlvjyvZ6YpZqwiU0iQ7QJv
kLnNgpEhpudwbOFdwCqJR1cl9Pp+P9+R9stQmXc7JTKWRAFL6DxeVlUUZxmxI8yU/tlLVLgEqZX0
g5c9fdqnz0BkzX6gt3wj17n8LaZxwuwDddizexrB48zQwY6Jnsw3JER86T92X+Km/7u9Bv5/b+UH
gdWvRtHPhSRXqCnuGh+c5XaE8oZDYQnPEZ0rVUdJ9rTcD/q7f8FeMcRJFWS644M/bT8u8jAEtyOi
4GWmYhv/vmd40v6+kDSwTY+OjUhPYR9v659rP5csX+ya11xxoV+49r/VxBuZtW/D0mxI8lmf0qMw
p1anOvUk9E8wCslTeYX88Nu/oDh7hMF65NTsQTHakEpx4weLlNr3gRVjENhGmwjCgF+fOCc8W1xF
XRANzLMmJj98EteLg+NrjhWCObEWag5dduRf+KerhW+r7LadbyAmgoo7mrhAP8HCwPAh2185clVn
MJQQC9a7KRI01/1/Eo04nOF5v5Y8l9pCTLGBoHAHmVxS7VHjfTRpSSuUBQo2DsCZqv+5zvyylRUl
BaFVGLh21Xe8glh6Ese7pOcNcLEtWsuXJljCste0jE+whPXKyAy/4vGaQ+C/TAZD2zgtO5zrLmsw
UeOZH7sdRp7ObVLKmPq7CH4sOsSwqYTId8z4oahfuDEn0TwIgrbu4QHoBKvArYpq+KwiK+8O6olx
KzrRYw0iKhXtWZmdPpKaG3VUZgn82XaHZzEzoJ8VL/mWQyGYPBQl4ThEUWe/5t4QLCQZmyQMZiRL
omllbZVHFgAL1EgbP1WVVahX5tAe4eAef058LL92tOC+8oPjNnYYPbugDEIuR5pTn84INaAiAYuv
dsp9DIHlwhAsutIJUzqhT3UpuM7NYtE16NxYaqNyCVAiEQPCWCON3TELcN3sIpraUftYlv6L7dCQ
vqlnpBleAUE9f4vxuCUaziO7VQgRkUeQopWfScS8f5hdC9WfYuFnRD+JAiY68aeKvulj6HVHfiqE
39ZKwJTf0Esru+ahVh+h69xV1x48HjquG9WI7EtmC+5VwTNIeBx/bb6NwpFrsKrvlCfNGFtw5AW0
LyUnCDYVmCN4fnNstDUaLZUC8iVK5qmjiik+WzKjpxjdOcrv4P+8TbKxZvy0cSjVSzff5xmljyjb
IAB62/wPRFc0S03c43QNmDtbBZaYtFtmMRXLM85QoqCROlCYSP6Sd4hSPd4DkHgQlAiZ6Ce0hggq
+Zgu1CMTnTqNjUuguAWvfVakYJedp1dBUQhJvPbEBeP7usq4bGqEFsRz7byCm9J7UILb4I4NqJzW
kijUhF5cbZnpkT8iFvF6e301z+0ZCwpX07+UPRxC3STriFPr1/rFBz0oZjKP41klg2Ci9nv+vBfX
vyYUFQEY5XsfSyvWP24wGDV/85DU/T0weoq3acEVza37oLnR7XWIvxF7LmWucmakQKCjVU6IiEUZ
WkDNz2hGUv1+TsrfHdC1q+0rdsMw9MW95mbvQJ+eFdZzdu0IVTLQ/Y1Y2yobsWVSKI9ODay3iHXR
xVexe68AXrd4+78vpUwCpOIUi2JnpVzowebNylfuPIsrV3w5LNi+GepEraUP/FTOigY4c/YX1XIr
n1lo/mAXaRJcWz3PMWVQjmYQlTOUOt0fhJS5HxYSZb0cZYVowZNiMcZfWfD+ABI/tLdrdYmNXI4Q
Ki0VU6buUSNOd612wYwINTW1lpILusfJD2qOkDwmqM6lZxiz+mW7gCl9qwvB4AeSHqqmEA7X+9a8
guqIboEMQoukqxqiGgHO4LbPHpSb7vh++ZkjRhcrYzhXoMhOFmVOu4TTPfp429lT/pyhQECqlPBE
IGL0ctqK31szjH/UmXjnVSTIsKVa5ki/SWfTYDpZY6e82gRwzUD/ACJnleflTzCqtOsWq/C+/iyS
UOSkDGO4ewRm4ySDZs8QZfOxesKlLUFcvbWVL5V2rIXgBl0tR5OsyQwW+DhrbkqLGdWpreLAdMIT
ldfTELfaBR88n0Su5jOsMR3fW1tf80noedwv4mFQk6dlshxuPELcRgoM6GfuzUx3daDPKtvXMFiE
Lkd4Z6DWaojLva9VX8VJKOy8msJFRScSHmpsrw+3Z6UJ/BaAv4yN6NtkGg0QZxByTegYvgcblVOd
zU5B54h3oNqMp7X5VTw8hcXISfyiD9YR4mreomt2Us/TTnSryTi9Hw4J9tzR1n/7eaSMolA3ZIer
Kn5s9OqPmc2yvyTXg8QcAKTXxx1/IC54eQHp5iZSPVG4XNKKY+ijfrTwqz2bNh9h6z7/59deA28T
pz9L7kpeaeGVpPataer31nPrzkG1QceLRn5D6M5822M1rdzoAUuO5UCuEyMJfQsIqzpO1dGoeQAF
3y0a0/2tueB5RDAvubywrXZ1P4S4/n6kpuu1njxZLYPZnW+uwQilbNM3sF5OKWe55c98VjZcFmvJ
5+KgpXYsSsCH4PIDx03zUwUmYJK0JVLQRYyNShcT6Br3t0Lv5B6kAVUIvWcTjpEsgGWNXYnU14LM
WKTjNBNIrYZSTmsGpWPhp5H4zvsRdBAfjbcHzTyoC9dMqqcj1FTJUruBKoQwQAbY7kHWrV9DSYbF
N/7V2PT/l+Gmh/kTu61EieIg47sFOYTsg8ejiFjNFMvlUoEsSRrcO1eFH14MWwHF3pNSzQ2KNDGz
grYDg35rsILMpMgPdKgeTZXc1QHkYp46BYHP856gyzCo6ZgcK+ChzB0JUnxHfL6CXGej49AWGrb+
w2z4Aq9nlXGOSFbZifko4dnbdbeLIcTI2KQg4JB+f4Xl29i4KuvBNCGdoQc4IRxMXUuw6A9zyYMQ
Q8T3A5aVidCmSD7iTB3eF2il1+0+Ri9Pggys5/566gYbn+OcP8p1LYh2eIh95GCiGgO7CCJo0Ott
B2QXGAlfdm7UdzPhy/svLkG1DfOEAdsGJShGe9CJsqapv2nhuoSE2tZVR10sNcyeJ7x9ssq+8Dcy
KqZ79nuIqgfq/dOrBZ5E1hZ2uxdI0x3FifiS0t75sgCDOpDs+ZyCctr3szA3NQtzDwFOkoUBO03h
xCz9P44qmEDcfJnwO0PjS6/QJNhYdPtesV3r2MT4/wVYDL66T9gOpst11WWCjoSSH3Dnu6pwTIaE
MlQTr5yF3GvN7sqCg/Q+H6FqFrjufrctbXu7c60XcN8+m6XVC0PczXHAAv/Vt8OE2nQITXWhCVio
aU1Rl/84jkEraiCZLuGqFUQMr5/UmD/eRCnhmchALJxsqUue0g68pLPNGyEa84CF6ecaUPJfXBRF
v/3VPrDomgB+vCITyXh86dMkGxtgvuiBU0KI1A3z/6Rbz46a76O4gwwVg18PLhub7p/Mo5PRetLi
EfJI7RgF500CNBx/53HgeUSCfzWtDDgBkE01kixnEw5NQBxERVBKPzFXt5pN4bNjMWeDeIACbnZT
svDgRbvV+/FgU5RKrt9NLeXF0gZbuSvuT+C6MxRRzmPxaMaT1dLXuZL7BKArVzfWwtWJnEyRog8G
X+Wf0OTyvwcXLhvfqqjtDOOxIJgjDoQpjgErg77B3oWrR6qMe0E3t1eEHCohrTr9qOgWvXZghGKo
sgNrPr244ggTQP7hIg8hJ0QtCKgt20WEXZGgou0ofHIZTMgoLXsLnuCRYYBj/glMSXIL2Iq3o0Q1
i4R7L9ZR+RsCyEisNmOwL++oISmk8ky3aclfZnhAB73WsQZ0KwMNmYB6tQdhLDqXkuXCrlsGhKoV
O1Hg2ahOsq7oMf94Ch/xFcyDv2c7HPvMiz57+RKCGvhevlavC+vxjkMXca1hT9nO7ifhC5s3BpmB
xJVnR8tBNuqwVONkZVKusXOTA579n3zB+k+OnT+/bn4F3LcpP1oTenJUwG8/wwsjTqgy/8L6Ru7O
dsOUlOKbvPGGBrJKMTEo6L1tCwrud1YF8L58Dm5BnJlwtceMpZ4Ikpo08o5YZo9ZZ+FEGBMRQLOg
z7eAr8QftqbiB5IwFcl9QHkSHrnfU8LGQN6ZP3w2VHiEcx2wwEoDPyE/mN1fGyJe7skNd9LbrKH4
ZBk0fVmGatxhgAOz7kwYTdD94oKl7YrumHY7jretLsVHSpInynLaQ47nVFtIukpqYtK+aiWoYv61
L/60KtT22AoDsaDZCOJ3ruAigyDTQry+XUkyv2WCHNTOIFfOp2qWBBQMJ0RrpdwhKxluE97h6XrJ
305COOMjxKmxq4fcbZP0lkgx2ZtfvuzL5Gh2N+Ls5XcK2VOkiEkEW4inkhVxxsNH39ftC9mKxOPm
FcxBqkzKk5kQFN3UWIQYxLiAEL2zKgK1Bm4dpdG9Vq9ugOAbvH/FNBP8j+jHcdRB0QTD1NEFT3Yp
htcK+KTOECOoACWaNZG+OThH7aE43FSlbFbBtGrEIHrEthr7mLNiO/LkxJnLH65WW9RHlTTMSSkx
qOxz8Pr8YxHTiUYZw61FMk31yhU7DyQJOIhYgjUBvhrmSizZpUZPB6qZqEiMuGEId0HydNpHSM5I
zYWgpz9oe40VdIfLanOVmc4Ts6kKotrebHtCE03WhT3jLgJzbPemA//Axlx8AZyUcleZllSXQfim
faBpXPHm62mQ+eMA42NAY4CRVWGIAa7C5kZlpxqiP60U9PKhavvIMoa6VZEivVTP39VmPxHo0pcg
Mlbaypcob6arLW0ET13yiLh6zJXa1eaE9fbQg1bQ9vKk8ZZm/rCNIuVDuC3w+kaZVppBRCJewEIr
/Daj8H4G0vB1NhH/vpB8PZix6D4EIIngslVKoWvWK41bCyUwZy2UtHH554bLxzN36dpnGUYMBYtc
Kjbo3/jVHwXfrJt0e8jx6lfn+JvK0jrxrTz2LQJsws1H/Ls9An3oCd+D2lChQfAlOlxWlxvnklzl
wOLS0DMeR1V1PrgXISTI01RUGAYbQCZ+bJ05HaxngCy5XO2ALTu3OvCVy/0f/FUC+JUa/ma0cQ7d
K68Rb9hy/JZVn2GvFYWvozANCgzwbeIok/eXvIHAsCl9VUrB/KHB1P/EC1ow+AIqYBDUu6cigTCM
2dAL7bcMT3Audbd6Wk0KMnZ0xw+ZNewcoiobrYs3E+z5+2K/veD94hRhJjO7mhhdT3txodkr6wZa
xFBoRnzRedQYuAs/nAlCtfSglhyxRxRb+aIoUeC1h9iJ8N4EpSRaGFN9QCEYXnEFQ8HCfqNtRBhq
ZcYcy+13wwlzG8BmSnkeWi4BCimj4zYOnglkF8n2sV8Bj+qfZQBCAXSKHXSB82k+6ReB5uqMAAma
Vq/5RTJLTXY0q29DrH82p6GOzbGHjuiSUVP65MhUs0jC1BSWcLwzlcSSUuRdBNEXYhcE/rwlrSE4
wwuEMC3b0T1bneOIwCyl25R0q1KKVgwJhof7+wlkEc4786XxXqldz2D1zNLcpbszZhGdt8yH28Ps
ve+kU+RprHY2IEk2SyuHjEV1UXV5nXLKGDg57wHJ6pbgdP0GAoNa4spiaKka7/ag8dC4CC+bQCwa
Wm5vOmo9RO9QuJOBpB9Ls4gdvGWmVpGhHf7R+1kSS0zKMaLjuPI4ZS5xc7+UGg9CJSuW26gQ3oxK
qT/XH/+EsfPqa8B8GamPJkI4d4oNJD2URJ9KE32zaDG6xK9JblS/2OlsOz5Z0fPeFx2lyFkuTRsz
w/eoV7ugL4SIKWY7FQOTbaCWpCka4+YM6IuOjXfBt49JDkfcDDtdTekWLPUBirLGEgvqHsbij9CQ
0CjAjs0NqPug3eKJQ6ycPbre7Xm20Y199SQfxzbkrQgLtXj/EoQ2AK9lAzQpV3QU5kgQs+rnLkNo
+Mqtdv05yrqfXI2B1CmKLwd663VxNOGjAU1O4jPIfHaiUtnAnFDf1/Fj6uIP02yF6x2gRUljwLBy
e7WAEiaLC37KK6AOidPlyW6TMDivSC2TldYWSSYmyDcPcoqxGOiAX11upBeTixtoZ1zaKFPkx1IR
ioUopGktRuP9+ZBoaM/ZtlpY7PQyZaWG1z4pxp1di++37YoRlqCG6IZl4rm0jZlQOMwkWPX9ptjP
ENMq+rxQgU6bgKnO4EN+hqbmW5JaAA2oQJHk7RaihyF/smMmPvt+0J6aje9Oim91/V8KlWfvgT5N
VompwwNgJP0Bd4iqgjVpaLGMm1ZOW/Vlu3S7E5p/B4m4VSmJdB4EP+LinbNbxfB3LBQzHyg9Fbnm
NvSLO+ixZa7DCJXtCwIuv43UoLYVIu8wzOqL1DXNgpD4GmWt5VYQscFFBEK51EG+3H21RvECj/HO
3fXVjXBcqoNDnD5MUUlLk6HKOOaqXbbe6ES10Td912P1VAEVF1BNbqTDChzty3AZ1SDL6R2RD9cM
dZf8Ai5Cs53ndzr4Omh4TDBFv7OXK4kHJL0TI+Xmfd1S7jkt1FxiWDKdMFFt+jKKMJQG5WNqIM9v
WMl69PnXuR4gOEgBRQxTHA+7XCO2M7unoDvOJTJBIMLFOy0fzW3SKdZ3XTZFQHd0G9MDQe2kvruE
uhwIrkAdCnsvH3E7dzJuz48q3NZ5nSfnMkeAnFJ4p88wnVO1yjqM38IbyHG1OXIwhFctTEdjG0Gd
DH1xNdFCxyCLAaMZvFhAGnL7wU/SPNbvgQiWoHb7xA0z7eyNWS7ihutxzuLDBKvzOeYQDl6iUWBi
xILQWt4F9AXnpOK+MJwn0qqXfBtde9RWpOlNulwIzJB0R50i6XszTe2A6wcypn/X6IQFBZuingwc
+ewdg6v8T63tzyiTQGxxP1cYPd/J3CXlVqMpaLtdQKk7Qr+QumkRzqChFltQYeR4pNJmbkQgc6or
m1RliSDEjD5fgdMPwgWBI02BozLNXCLrMrxfn5gOZCyB8pXe18s83G5xjYfKQ8Hpk/rKag5q0ywl
KlYT4t81mMSBZ9oloIxghkPPha63yjxU8JTwt0Wm0SbiqQGtv07o1TqBRbSuTwawfCpJXH6ZXRD7
j38Aw6KAnUfG9jWFAKIw0Y/18nnA8dL7SnuN4x1QZraUSWINpZaYy+cDYrk0PYqdd21MsSPCdLmc
SgE8/0MYMBJgEzOHBk08N8RrYmnc3rFhiTwgLFdI39juIsFa+x8J6+lIXQTY+s3KWwuXT+O0Dfr+
cfCScXUGWucVUJLkM3WumZjjB8FqUAVzdFmO74KLmyA2b1Da4t64HkEeCxRKOrpC3pVe+o1SyEs9
9A9DijYzEn3snGINTMCnk+K25S4h2IX/R4+yzjy3hNMgqo57ZhXuNicCEu+H2fvt7rEOIo8Er/GG
lhDkeDQGkCFTazwPenvgTjEZPn1z0Rw226dwIu0kdV55JUTUyGeV2wFKIlr0vrQSA9qCrOi1ylbB
eM/ANkDHLNks0uN+zTXi6DP754Hn7z74sv80UQoYml1cYziQdScGdCG9hJnM8zpbV1a99DvfQifD
/YpkQL1mmsCwxA+6ZztRM444KoJRJL8/0wOYHR/nrAw02lNmJbjlsYcrt7STbo9b55wuUhGV6dEk
5+QTL7wGw675a+sPGs67F4U4E5jJMfcKra4yWV9A9aj5JYIXJPwWMlPWP5CZjuoyDB/khETp2uyR
pi2GkMv/Dryw9TYaYEgw3bIdF+DQDSnp4REUEOiCD7HxNRufHVDZ9xmpMjEDVsZhNAZDSgr2dBPA
j0tSq9TBNJorGHXUAACA/yLcbs/t8e5ULnPeWVa7F02IfpGA6aIwl0ULTp3cwFka5NMlibkyvxK4
dXTrT/salyJtuP5uKcwp/RJd79+cH4PK4pd16OYJFrLTi+fiI34bjgUSR9NTpDYq5o8MSTXAkAgR
Oc4XjPtFbqz++cU9QCW1ZzV/Lia2S2bKrU4ZODF2NcSHcIstXbvwX5FhVqrtt2qjXyDOaDRd/RFq
U9C1U7OaWMx4ht1Jxa+qb6V1ZrVkuhCPfJc8uPW8RNScqDT7hpElHqLkRdwM2RDm7pX0ECYVAkL3
q+xnbMIRcWg86YQorOLloN8jRQzOw6MvNfgOJMd5OaKvhxtl2UhjOBSpnP28R3pK9L2cEFUBZ4od
YT9hwjb6lrNuEXE8YNRHb3A0jvO4K5tKEa+3Us8bDSKec+IaDsChllTrIqLzc+LHjrxj9NnaPbKK
+yDfXK0WS8aFCJ0fL5sTOlwMl/hyfPhdnp6GjL5t2V+DjXF48oi7zhhb8uoiEGE8h1GM4lV8Tx5a
5Rl/WLyWUHq1iggtvklOjDXiGqcYH05yPydWHhmYra1fQCvBJsY5hDtIjQiFgTvfYv2LTrJ0MM9s
IUp+qsihQWPM9phasMZJRpQp/4nJ4zKuoRrIg5T45BErJOM+vuav6/C0OFsUk/E0tW/+C8qEzrVJ
yiO5U0oxsFBSvONnd51ptJgOCTIqX3FBRly1DVYU3nj3EhmizUknaeAmGdClVNNmjkA+pu9yss8o
j8B1eDUBk7mMvUHyyzFNYNEWtqWrs15pEQmPghkxGmZ4F9TPTYYYxafmBFF1xOA2JmmLH6wAt2Td
wfdhsAnC126jXNUCcQ+J3v+1S4+oJ/hPFxMXxZctfbdycrz75hZ6tExOqMoEr+3WGGm9Lu0hi1xb
8CE7QxSiIYi3LrqfZGbzY8npPwK7vQvIquFffnSEfr4UUQG9waLsgFRQ6v4i/26sRH8K2TQ7gt74
2V3tMphXvyJBvgACq73jMt2ke7rjb5znlz4JeFB/219RbM6lFplTCjayjnfuamOYF2gu3V5epHn/
yo+ELoZI8TvReMh5V/i9lcGzedPKZwJsfkBt9PzMwzh72ggYz2ybp5ZYGG3TeKoBGgVFHQ924eAn
P3csaG4JT28tkEKRdQaDv/Z6YttLomROlSmM4sN4PxXHDYtJ3aV/FIDcjwxvfbtimfLERxO/N5eR
avME/PdCaGpKhaZhIQwkNYow4Y6P8U0CJiF98bWPXjQrzQT3qQhoLpKvab1Gkty9eVa6zwZLbM3k
5EYm1ay+6Q4ofnpIP8uwVwNuZESivM0aQFD7T/GVm4Z9htY7d/pvzXZNYzkPsbqVdxWr/M/0nN5L
45PTcPhmH8l7SY19adSPS7d+WXbx13+0dxhdTObb1Cnf67XXA/iYyXQGQGtpGY1f56LyNGc81F4G
H784ks2RYUAMn85ZzwAZNg0M3fe2o/mXh2uM3HVi6gQ/r2Vd0do007CdUX4vghhctTmRAZeBRYBT
Is2vp6Ri+e3vr3TYDCJlQNZwUHLoXIZ34Xy1wZUcS7vVWiG6utzlxl1ROoSgTLP1RMeXIV8h2EIG
ggmYVLdXHhkxAFSIkWhZ/X3/cSdeuBiNlM3VXzB3yiv7aJQ9vxaR0lpyu4ouB0rdYy4x/shpIGKr
dPXBp5W25zzNgBjPcpV+yVBtf+l8VnPj3Ov/N8mWvE+7Sgz/gsLPku/80WqOIwyQrTrKleHwMIKZ
fm2Z/DBjXCOdKSPglLKrfRJ4C8VyC5lHMmVM9zve/abZa125yh4Xu1QClr++vue0ViYtXGokzrY7
jO13/kdgx1YoiSZXpfLtTldIXH63J2fcTROFAThm6cmhPdcMLKYq6cATj4H7R/DiVlpBkfHY2wTq
EcakgMzmcAm0ztwDRiB3CTWsWSpqaTi5N66+xSi25wLtM2tgFnZgl6zj3O1/pROO84+CBMIIt7rZ
gmZE9n71xDpVCdibgCBuPIjGVRMsdYsIcFXAixlaAV9nBjot7E/Ek8WFMyhkliXo+cyJc1nE5iXT
Ujxli+FtMi/mWKjU6xLKhDDONqvVvh3aw/dI9YlY0UkdWEXsRVL+2YcMBSq4P6jfNAJ6gdOk/UX5
3T+InxTRxTgVqCzkwXS/yRK0DGCjJ9+Spc9t/28Zeob1rbL8SSgwnldcgXCD4wYG508/9DKHi7N5
PxCh2sQNfKHeEn14pqulZzA5e6tjoBsNMxVMW1f0A/z+wQUzqDoxLoE+SozM+B8A36zXgPy7dj+L
HHl6gL95BjU+f3vm5wAxjldrTQ7/Ssv/ZnFCCxyfI0/b8jm7cVVUvdAGAmRfTpkOo+PptHC97s2f
QpXb+lEM3PMWMQeGos1dbQMTsz8AKNWWAvnO2Ppxtz77eLRz1hzjXXYypXs+BKrJ+hgt8li9egxP
VQfbJLNxnWWLOtXXqlFH3Zio262S6TrWdVOKSm9QeQ10zOAjmMNu3kijotUCsrHRG7PZczDTRHi0
N5RyyQLlfK4/X7KfqVSzulxFcs6J3zPhEqDDzZ6O/dfrqP7lp9JTrq272ZEn/KFMcJxTgHBCnK+X
UDLKYFlSgcLJUAphvLlmn6FLVbI1HDdjVV3uN6+sd6UvsUGf8C1yz5vwlwnp5TYoi4ASS8ISwytS
2u/EbO7bWDOb5XXlkCnPO0C14xufgzHA5Kq4X+4A5GRcHjCOzJs714Leu4QiSOlvHDQO+Q06Yy5H
6lMLiDCpfMDwz0tYOvArPWDJv+IBn1z5bHw+MXeGMU9Ez8hzJ/cBi/ho1KFJzSVW7Gdn0F+yp3E8
S7OqxvaOq/J4HCO8nEbJNktBLxA3Vj/fqYQ80vJn+msSz09peEOcBuhCP8MngEqSs1Kgji8J7VAA
xNuAl8cfpK+5ZREBsaZN5rNARbfpkxCpgHvcAMlTl64gWdYy0A4YqKHrmI9UmZJUduQo8MftALW4
0pAlQ5vy6HlbdZjbXVLjDiTLnQgl8mq+cvE72jEtZ2MVwDxb5ccC656ps5eWAfIq1/lsenDwXkl8
TW8+lByGx3zqxonOPZywSNVBX80ZteVOhdNCSIaESs2A7CZx+B/VL2v2H1XqABKpytJWoom2zqXV
dQzNx0HmdoMOk0rFz61vlPt49FgEy4irvVMNticLvZ9TKuvLP3Z9ly/RF3OEiE9kIuaclW8YGaql
MnekjLcxG35gtl1f5ToJRHctJaFeyuLDrJQSTJIwn60H7wirkpK4s+b4TDJWdGaGR1k7vlZVs3lT
ch5aoeHcm07o3zn4m4X7ZJdqnuVFpwQOoWUbpgKGJWJwxQdS17XpI6zs09429ZK2E3x9FlCfkGph
NZoGmX1y7gK0PHvVxxEQk0D/1CNgdDt3DDdcXDf73Gxq8wj3WAmRWW58XO6+EONysvW0p92dJXUi
IBO5lVTnFIdq/sAMkmzg7oFL2oRJ2GtOZ7O8rasqxj7Vpwntz/dvZ5rq7sI0VdMu01Nu3rjyuDKm
NN2LruO6w0hTZVt0g6bLxP0Oy1PGn4iuLvFjG7quzs6FJgYKaRb+z5lmRD98d+i6QgPfvNFB1gU+
/780tl0F83hw5bg7Vj8dA99giM2jDwgQZOUaygsEu3YqQKB276/ocpm/jPsj0/6T8nzGZfrx2I5P
J6BkMYw+/x7VDefuhVziScHaULkS3WF6oa/ogzUzdgQhGASxtSwkNtGifmrLbHaahISkfxJCbdF/
QY/sIZQV5eVoh0b7Rf54ng2gcqA6tJg1iBc1E5Elv5nDrGxTtONMa4E+GPCzmz5EU1qK8nvd4yUJ
B38voyLpeAHTubz36c16f5sodf8A3xRQhfKvo3xrRndAeuaMaLDwMnDjkjM5ratJISxZO4/JzMXR
tvYER1wPVN+hhEn7B+dHvHrBMxDSwCj7f+YBH73PQaQmljyXT680Wxxx/uRCANpu1ANLX7dw2O2G
Bjdc69o02jwv4b79u+EjVznNnEsvgChnEN1dHDpD3kh2WhyEiAfz/unj/6RiOlEru9OOZQQYA2Wn
AuPY2o0m/oV34HLTfnryo/xrsvXyZ/eqZLOnImTdFR9b/mhOY/mWSuS7RqvM/A2WZYCsUQGcx5w0
e0F7r0aDRcbqpsOoFL1B3Krwv1qpB8cQHP8mPPTT6uCWRcAI6LqYskiwHOPxD5u8Du4QTVqg6Ps5
GgF/Lda7TyMTnVi9hPKWRzn4WlcmzV7HUD9kMheZw7qdB9rNqxKEpKNmpF2/pKrSji/3gRdgV/Zd
QSF2GGpNCyNPRkiDZBmo7XpSj+toOJI7TZWx9Mvj/IQBkQH6PBgZc8sJf6oU9zhNMNtD/J6dVQFs
xO/Oro2wfv6qkYPjFpq4IYJVV7fqQqfVXojiLNWnsGy1cDz20gYoXhtEq6qNgxerZLNOlUxY9D2g
QLdiMAP/sLFEJE87vBTNtzcjju7dphuc2GU9UEUNR+4RWXpu9KfjxYIyN59dKz7YgGaoVg6qvHUs
iAHy+/mgSoJ237Wmk0QVJzV8Surcrj4fzBy4sXG569y990GnEpI5RgIiphVht/XWtSTI2uNXDSj2
ad/oP+F/iLBZEBj+Sif43/2w/yv8NUYNslS0HJqehgZ8b8/ZBv8Vw5y+IgPdQJzfkUc9qWuKU/p+
cxnEjGQimpI2dQZR2BRrVPOqbO5kE/UfBf3xqbuFpMo6LaILAafINcdElFBlzeIpX3oVVBxHY0sX
+QXQiZd1Q9pJQDhwUmQHOMZsVjWi1mOLJtpIzf4348hP5yD791ckyO8ah7cJ58or+VxdFJx/5DdJ
SwS/419drrPdn1vdOXX+DYWhHrF/m8knpqjtnrw0vmyWj1tlSzAZE0j+DaIYo8+6nT4e3z2ECiJk
DOCnnNpg3A9GXq87xScwXh2ZgMIAUNGJqdAsZ6k6WwlSTtVGVl4JrwoCRBTVQsAI3IQaYuANM+Zx
yBjgwI+Yhgx8/Z4ybII8hsWFjvObx2TlzvrlxgyWgXXubYzy90+2D+VhRaAqd8VNlWn8I3y0yMtt
L1K5ulXaVO/7pXKNBUQLaad3C/zaDcs9+NFgF5lhiOaaI7Nlr8vDeN7hvLMS5bywBGg5BwzZoxjH
g0eeY79s25hypJj2RyDpSGLIHmxyrTtQFmG4J2npB1by1ToQ50+8WppKV4kyZzimNMUnV87w9X2T
DHPPTpvFf6GyUOc5ltPeEDTnTNwnDjTag970a7cSqEJ7nmaLDtjwbN+lNiGILz0hoJfyfzz2bv3Q
KB8yFUufbD0y6NcgniL43DWTAD+1oXORvtOuU12n02P6TGhaYP7BgaJSdgq8AjsD2BQDHdGD+9lJ
MrLRach7HOW2KoXWVag5QXD4gZ5JobK6l/YMGVQr9mfl/LG9+jlMcS8LeBdlvL+4ky990eYP24DB
Vnjr3qK4GR/Ub94aJU7/NfGe4G0VJk0RvoJac3ZfDOe125nD/eLo2bfs7k7kPTqM/SjPeyxYiWE9
eB9UznN9sG5nwb3fLCh9AIVV0Kw7DaVroIknWz42L0fD9aX9n2KAewZJoHzGMUGe62aRwxHF7CjP
2v/Hkv2pzsdHlit423MwObXEhsBldOQFXE5jnM/G8Ev8mgaWT7rHNvA64h0fi+nA7o3SCBW90EX9
84wHawJDfhPaFNvDPOVb/Ru1T3hVXwT1+/55gyRyLNnz/VTPTzxd529ZEXhdkn1paqZ78GxmAqUT
ixlF2pzhDuaov3YttzHcF45PG70BwSocBpM+Yv1E7iXayGq+XWXd0agWXKekXxdI2QvISWfvYhBY
hAz5XLXNXZWV7l9k+m9VurqJGxjtc34M1dUjfIJObzy8H8Lp5hadyx2OlvUJzEwVLkFLS4Nlvep8
gZaZMgBIHgqQvRqQhk6eHg371hRgO3d6utzdA/u9lOq3UvK6jV9nlykxzBi4EwbHIJruAGdIMbJA
v6BfVQHotlJUYPmBl0PZJ4tEXb3920vP77CPzLbrM0M3NESXe7eZF3q3lmlme+xOHnzNl+fEzCfG
alD91Ky5/AvHEYYvHgbtCx6i7EraQWHB6Te9mt7YjjS5nPDSXTR6/3iWXlMbADJTMKFZdLRazIPd
MQwr+tcZdIbuB1m9qeaRCOhr8YM7GgpGf6+GqvBzJPrAWPbKoyl553Pr/m3AMjZDmW82HApLRlHD
vI5vFbmR90JFPcezOsoQCxZJUF3eSPCFAVxXPI/hbIw4yEgHuthAPzvVZhV4JbRjSX59Mbm0uf8T
glzlvwRUy36CAU/V00dZ3/p8WCVb5Pr3hVWFzRMgVAljJ/euJYMNo3wYIqzi/ikbYbiKocB1bJad
0WMH/l/G0UGbMQMGa8YzeR5TCfkt+wBLM4+UXx0ns6phDX2JHd9mJoYqmQiMWppavQyf148RuSwz
uPO3I0/tLv4/p0gevGJKzFJd933rq/EPKPcR/PptcgkRWMSZ3fqraXUGSNKr6DSO1FnASiyHTnBW
EY1EAMcgscWDdT5Q+hmv12FNQAurQ0Nno0/7mVKCVeUUqOiez0Tw42Ktqyi8FPP+82SFMe+B/jPx
IJFkwn9oqFl5IzLqUw2UlKVccCkLnnhgGNNeduCREJ2wfjGVGIH+vmI8RbCrtDxGsKXGCgVmbUqz
NwmlxIPSZtYlGrUZH7k2/OZfDk45bdsK8eeferCOsrGz+nKZm7eILUp8S4Q32zIhtSoYXvKf+IWn
wCVHHCa6YZvUHZ84OT0y2xxaEU7LReXD/SMR8qLfoefIcjlempJQW5R4pLWDzSf7uUlkRNbvSBUE
nFJIL/nO7ZWPlWj4SNlEaHJ2ggkpvHFa+IBQPMjPoFSqamwQ0vOUSSN8LcIp1WjKfx/bLmnpgftT
Ezq2v16a6AupGuxTiuKjI2KJsyqBIvn7LnJfjOTkfuydfuf+A2YzMG0+H6LZDumjJo9/1c1+m+Bl
WiwHBoY0ovQQTIVuBN7D8z8zOOJHg7AE2HyPx6bnl8HxkqjQzwGK2GBmGQsPLyD1eu/rYxZRWBy1
+zkiBrUZrIZCLduQIzw/Le8uiUfQZ39unqPPJdPKKfSdpyCXk5j3TbPeuCB7ul9xfL1bZ0jVDI2m
wtEgTltdnH4Wz+S+616JgXaAuLQ8rVMNs6J2ZrLOOBzuRQUBhLf/Feuh4Xd0ZEae0f8vsvdCSnri
dPgIAcqRC+KDmp9LAElidaHHCKhW0G7UONxYbhS7Nw+8/RDAR1Mc8JWzZgGXG085+RvvrBUC02oj
y8YKkcyydWOE0lpLIjwbCdkUglx3Y53bUJB6Z2iVFoeyeEyq7p7VUYbgApkJCukAeHlYmFQdGHiz
680XCE6LsisgE/svYKUVcxwWlC6AnpNZitSXqMHnsS99iVxl2Kb6bwx3FxPuAPJWr2y7U1WbEATO
QHWxYFGlsh4q2UdrF7H+YwkPCfKv2ustLzv0OFzFCby5oozc3I2aR9ty+7CgKyx9h1sRrAxosalr
UdzyKub6HGKKPcVLtt96MTK6o1xSerjjtG17ZWDnF3iu3XdF3dvCHwFB0lqHUfsUpWp/j/Fc/jGk
A37PW0ekkSsFvLglxfrQTUMNTDppgi1gNI/q3cyzXD0ZYmA5CVD725S2kzkn48NvMbgBWYsTicp0
Bs8YcXqJJY1c8AcuTs2Xq+OFneepkpLnh8dvEz/wTX3qc64Tvi+6ky9FlIOXTJ6D2jMiBrLzwR7H
Jo6XN4Ntn2HPodHJyPiJrH3F4MLqtCsijakMrj5Axpt4VBejIBtM/WA/pTS2blbQsJS7Y2rreAMg
z3oJKUj5OmRJ8LQ3QsPyBDbM/kR9elx4qiv4tQHguw4MxFaSropJFk0xcimHTZkvvojIhbsWTx1V
W1rGYJwymjcq9xiRm+4RGn/oLzfueMM2spDjGHkpPUPBqYsWzNvQ4DrIkJQohh9xYbUnU/gyAOy6
uNUeM5Ig7Vp0D+VqSkHpkViGdM0iuxAocPJmJr1Jh6Ln7vWtRcaaQmVUXFrHNsgdaYTz8m+rmAEG
z72wO3BXpltln2hBPaMHpRdiwpBzDYFEB5kBhULNETBQy018eu/onq6v/kh3XIDvhg4sQ/JWORNJ
brwaNiEDbGNENZBkCopYmXNFq0X+uvU5FhH1ag1SLtSslb2D3Q2q3MCydGJyDM9LwURYvnb6FTnW
SnbPFvtigCEUOPA5acLwJUXjALMmdEnHdgwSkq2TOtXsZNFqSHUpkxdglmnmzcYHIua2h9ZaBTyh
WP7A641kCKZjhoi76spH7exFMD+EKDHWR2Z5cd+5Lwl6zMfF5Rfbwuuvw2EQSiw6CfIT96Icky2t
BClB1eSomsXPZxb4NdjBipoM7HfcBkAvByVpTmLlITgYffL9OQxDHGt5YjvC92aHnBB2hxdYtd+d
fNGGiHb2sfonc4CysXEbWP180yOek8heXCO8T2GzwkgyFBGW77aAXDeAvSZmnMlgUIaXytIJll2G
ywKrBXsPU/HAp9B1Kges//OQM28pG3nXk1rpbIiBM/Qsapuxv/fckStc7ZMZkLV+I89+yDiSOxLm
4vZWIfzv9p8oviPj/Q8CXQAOTW8740z9jOV12R1FpsAoZ7hPkU0nOQNhGkfEGDfaGmRc4hgXy9/b
aQkvqZtdrFs8JcrBeNA0cM2xob/J7lHnHx7NUizjwVvqpNhpUp4ylRbObi0lW+h90wXOsKo9r0zF
S4yfbDGFF+7/X3SheS452Tf6jM023pJEEOgkNkB/aMINTpUYq49t5qoDLMWzOVO+ZndYKHqBXCy0
Yht4KTZvIyt2T5o3mml3YMaD2ZpMWSGJB84HmzSpSsl6FtFW5W6ClI8IxqSjQkTesS96Vy+4enWK
C9Az16/c1dtxytXIjzM2qSQrliQYlo/TRUqX0q9lAJCyz7D/LrUcgBbzLG2cEjgnI0YWnE2EwlyS
nbnIuSASPkZlAhLdijBz9Vn32DSZW14oRc9jgI6O0zoX0XwHYMUhuRNLUx//Yqy5ZdZ4HL6vXxnI
FfacjEE5deFVlEX0QaLGLPEB7SZhnrAx/Iw+l+jUMilXZKexXck469Ex1Bq2+Vi3zoaPniNvSB08
n2ZTg6fV/6U4ZDFYchsIDF1LhuqVOAChCMAENxruYKW/PDkp5u0bg1xF7X5oymvJ2UwAgxHszp8C
yZt7wwJ9AVTqa378imYcA3Bzjn1d4132iX5Jrz/swzY6npq8sV8CZ6dXiO8GS+sn9I3PADY25/O4
DJFhe7InmNBJMv4qKvYkIV03UAL7lQxhaJ6/QEt2QiqRKowUca3rzdtG3gPbg1KPeNsvnlYOEpWP
C2QPe+780iwkg0TjYRMGIYmImzSOqcNecpi80of4BA81E6e+5budzxIc2Pcs8VWRCxuvOCOFdOhm
cJIf4x7xpreQ7kQcpJIwM1l4am9hajR/6P4LDJgIdZJ2E4L1Rkylex9kY9LIH3Y2SvRQ7cAfU9CR
160Wlikl+42etIhvHr9u5uhzKQXbPA++dxD2WTTROdJ6M4KT/0LPIBKlFo3zNSfx/cMl0oKe4/t9
EYrJMwn8zOxxA+2xFAUJpBuLYuwqzd9/HMwch8jUMkH5OTIuUHNbHtLcbB8HanYCRsiAHZ7AyRtp
yYuugwcpZSIb9eNqekaJmPGTnr5ik1NnONot9c6uXnwQgGHyqhlqtOuTexNOzgb5eqHY8fAxTPix
GhxBnHWvKV9hkT4WWqQ2R1Vc6BKWT5/tlOYJGoE1O1vivvG0m9+BNNnMf8qBGfr/aLogzor3+8Ex
3WSjFGXSt9qg7y39ixzsxJl64x8XGv36x8beIt0Mx2KbffP6ffj24nkrwL5rC1JSWXlj4v9N37Zp
hwzMwgOLM1oWgduWFvOHc7y7JvM3K9OzK3pdYHuyUWjAXOtB4OtkUzYHAnq2Ou150exObUFnRD/u
uXxZqxwn/MLkZ75IMYgZ0PnPMnpS2zKgBFfwbtpBTCOR/ASsnCF9V9IIulQbYXtzkLPkTWCA+YK9
cuFOlLEJA+aURFtvTGJl5DwIR394jBULjkNrlNOqcZkFP0kl2BIsDrh3dYp2cnsmQPeYUzWaHmqS
gJ+snEo4H9elJfPjr6WQ689g0UvfhvxQcGro4EUZQGysd1gYdyQ4JsAZmAd4PiT8G2mm081SszbX
CbfbDO1wH5kR+PcaFIllYodDl8t5rwYL7APWNX2/iLz+I06d8DRGUhsy3LAg6E6UH0Ls0DYp66/F
oZ6L+38SXbwG9+Ts+amK4cxJoV401HHWnzV/xyeih/wI0A+yhft+NX4VpyMdHSNIGKKrMXUuCjz2
kLpYDb71Gpth/+kDI8Eb/hie7tEnIMDoguFr1l9BJ/4fZR8BFT+/uJLaeEFCAIiCvMa7h6WOuOdG
Ym02I1I8GZc4+TQxbEowtWpBznxO3AK8sGPu2+2IsainYNwPsOrZPz8CSj9Y1HeqivJpM8S9Blyn
7SHOWq2kSCG8CnDDDKBSB9zZIWiEpysILJ5mL3i/cJsnH1QZx4RO6Aaq/NOHsiiJDbWSwC+UYyQf
xWuDpwJ9EYo1dCN5NckPGEcpqwzJYEMjCKC9i9G3GlAny0EUziIQ3pM7mwloXAHucZNBGBUhZ6f0
wqjSbMEs+rcvCJ1EMtF1NZRsobP/fwffMlqkLMcgJHTS1n/GdHuRAf7br0vpMSjrmdEotux1V3Eg
vE4vPgJcbfyN8k4qASg4B6hcMqrOGxqP7aBnpP9zBC0KxQdANVOWUPBmt6GR3tNv4Qahs/EUciLx
jN0a3ojYAyuuf2gK+3s2S2gIX3rTcq7XDnlQ/XXJ2uYKub4zksJft/Yhq8YZCbwdejXduEgdE9Ts
2be8ot+/OxEc/wi/1cpXNXSeCWqkYhEsb3JSYMRfIa6Lg7Hs57vm32hSlh0Js6x+37uIpys9BtCM
QUGfCqfb4bkLW6HJ0oFWMPUNNpcTHJuaegkJZx4B32a07J2yJYAZ48y2N4Iz0AxVoFCG37SyLug0
fksFuW0pDn6tOciXZy7TCHdnkcbBA/QUTChDaT81WexHwjQx2kxz5XSifNNlMaoWbW0cunqtZ9b1
JeC9wfNoe3niuQi+BCrrz6nooiRRqmmr0Ez5tawLTxtBVtUqtZSQZVp98gHoLfG3G3ZNXxc3IXRb
2ZRXroM+sXljLaW7TiHI3Jrm7GRIGt2TrAQcE7k6i0f4KGdb14XRu03FYTq7lJ5ADqmWW1TPnwB5
ahSXaml6COETEjWChWfginhUO0wQIu6BizAggWp+XuqTG8czJIoWKOmT8pzPv9Z22on/bXRN2g6/
tHRgePmpBzfESbIXRMTLTw4M1BHPv+Cn0Aiji4NIW9uq8OJCUOi6KYT2+vXNOTjTV9b0tFDaQejh
1goRerexnQ4aLTViEwKcxFQVeTGcH/26/vzXgjGYgqeEHE+gprxA/6u/KpV5Aak679N6J5BgXvHf
MmX+4RSpA82dIxTztMKPx1bX/PpA1+yVaJEY4vXa4FoynBmxkZ3fU8r+iqTgxsdGcQFfRfU4yWxr
CXsVvC6a3zQ1htz0aRZpqXY0k9WKJi913RUctVaAL4UQYW26FtO6N2LGa3M+EDDYuHVeERflDalu
OH/kb3vj1l6rtaS+sBiy0JM4JN/DnpOUhTlfO0yMO28Y/HfvARBhVd17E5cS9P0pGCRowwjmwBx1
RtxtAWD2L3SiHr73ngForkJtkPkQ842g9KOgmyi3IjNjFJ1qHOAZQYkdRmaLDOoLnHrElWMEh+Pf
hwiYfhJrTmRjPp7cNbS9h4guOPZS9bRyb5RzUCCcEeRncm4CEGTMUmEdo8+YeMbNp/RALHHGmhaC
kLCiO+x4yIVxxaRCkcpHpzco8CF6Hv1TTUR6Sd4VYqgVrKmjFQP50O8x3CckgtXJN9JSvRmu4ubw
79cUGl2QBTv4Jvhv23rsy6KnfuA5e8DLjbrhT/jac5xJfi2Lfc6v0WlPIo/jTqQg4MDw6WGtWm/M
UGRde4TT25rTbael7F0hOToebac8vjazMHf7BGZWsCgry3rcTnvw2tIAq/4nad6kmW3yx6XDGk+J
4AnoTkVOJEZ0qgmdTI3Lw3CZGHfVAbpi+Sgq6Wbw4jT3pQrQq7DD0DcuOqWl4cEmAieabVTwEkdR
aBmFUPz1Dpg4QxQQtQXH2CPjWBFPh+mAPl8rX62BB+gOtEZy1IFSoB5AayQjQ5eQpmie5gMyWU+L
5LzjBlZdM09A0GXh68AyJskOFh6gThCXDSTymZJITdiihYpe/SLqlB5EbcTS1Rob1QK1lsRh8AVs
iD7eFxtwo3Gji2xZPhRyr/ChYSUArW8TJCWx776YTteAFZ/gSWFhnX0cIGdhx3O6z6PwAjEJY0b8
ZMDymiadx4G0BoMEO4GCm23WO35Hc9HiDPKLNLVJbrlJzx3ZEAOTQ90kKKEeMgnmnBwWmZyehZvw
CPEg5MQL4eykrCQMdxc6syefMg14nBoAdC6nW8cQMyApsjUmm/3/JJTDD8M+HtOBSGFKX467d7zd
QFQFad5eWTUL0LPIdQlcpreJ8K64C/1wM3P6EgMlq501+iIrhNFx6XVHsGBwX6usYSJ863VgiVaJ
DCaV0pwzEaYEPtUuZvJJ4ZZqi/0Sq9phtD3Glu+HIwbdxnkw44nExgNlUW/z690Q29kRfGGu5TMI
+6LMSMfxUQhhnBfZpHoRZM3nr6/T+9ZV/qTZao7MJUanl27f2vMLzzFAIqYLHRwszRGa0svlvuxA
QpUbG7Jdktyv3KFpiDQj3Q8NPTLr3woqwlrQgcZlAYOSOKfE416g0URKczbpDXS2iY6OhejrxigL
5G/FBQqYBIVveEPbdADAYevImWMtt2hUkfK5Tr7HGGCXojtgV/b0f/ZVMtd9ARci1HALwx+SoV6Y
BXYqgYgegC9LrWcEzzMWozJwUCna62Z5IHeye6kpuGZ0kzsj4BAvMYTO+8+EQ7ptevUaymv1P1SN
kbmShCa4S3EAUvSH5hqnuADwxtDOGtdH4LX50MHLc0H75vlqaJLUgfkIXQGneBJKa+1+gpPtD4bz
iG4ZoCuL16yhdkyTeaPeqfpMlLqKSOZqc9rp17NS9XKTLeUCM4mKYb938fNmtrZnV2B820AflgbD
KvAX4x/Zbl2Ztl9fYrn0AucDlLKwHrtxFt6ntfu0S6dyhF9jkX95F3W+bSMJbbI65Sq/InS/3FMN
LHw0DItXhKVyCKX4oZb8oROWkoH1Z1iBZCQROchJBj3bl+BrGaiaNoSeZX24P9eERhb2YXKo/hxs
/r6cQOM5D7kute2n5blXjiZXMr7BfmCNUeT/u986R5ybgQZEaLTbUIh4AVMbQYqGhlH+PtEgRGgD
Y9+evNU3VrzWuO87RS4uY4H/wcY0mziJ9ZqK7uEyzZxlGrJXp0dsGnEuyhgpAKRDqxRfJdz8wp55
FdTCeox1Xc3jJm4Psu8401Hsup+0kOCcpAzyfC+3lhPoxDV/ICYHH1yZfGhRLOoKUTN0cy8ZMcPr
gqC5CH6D7iNz11dH/pY76S0ksjFUOKM/f2OJXvzh9a57LIKE+STqEtmzwUPtCVDZRMJYDr9eHKuq
kHMYTXnNvfoFq9KSNA1uT7cdpGU1QFnP5oLi9gTQewI215xcEFeLywWZrh1Nd0fhwDjmtNmL8K9E
4VaZ0QYmYJBFMDTFdidhjI4ntn+BJDEO6p/G3EyvwKjPgbDiNtHlIHfXeYcELV1TIYAg26I5uPnD
qnXG2wYKurG/oKn8YMbt3EHGHtNjOmAINRpNi3lUy+Ojn4aFbuWtWEIHLm/F3a/JvfujkXUg7CYr
RNM7zlv1+eJSqQT9xOpCe4ltHHuoL5TfbdLJFxLNmxzhTStTUeronOglql6FK9LEDSlSvvtQIhf1
8duFCn8zIkrKjX8X5WA/wPVBZWE/kEfSsCfMoR/1DiXrrOxO+KRrUpVXH7u6ZUz0f5zsHNlx7Okg
jWY5ijpaLXaNMvItDMILzp0DW7gzc5fg7R+6/rQt05o39kppN59JHZYzSyzR35m/tcVyOLffCiVs
/4/HPhN9qunY6E3wBi01wLSCZVj9cKQKfH1BA8o1e1piuSoG/PTX6lgHCy3ysZNq98wHCRojGrqj
02FIa09ZtSFAy+1cME23WsNO0qPdXdi8QvgypAyreqK3AVvK22zpBSuoaGq3aSb/AD+qZGlLds5v
LyX8xcosTHegtGUGxlU1rP1xVW6544OExddLFOZTMBMr7iZu0awUaN8KXPTbZOXfDaQLaP5XK5NE
3tLtS+AFoFXDgLQ5p48r34R4Uu8ySpRDbjLyD4pgUz+yoRX/11rZVPaUeUB07nbdFpa2M9rDhQ2w
nwTcNHtr8Z0nCTgcgYt5Qc1064B3Vp2WTzrDOqJhufwZ27IclPuURTfDjy5F6Wc+osArPwI/WdS0
Ih7YnaHY6j/Ne42NQQ7ZtFR6oOikZEYa76lweswFCIkDAHKrfcGWzbTeeipMPXeY6Ax1QuY798ER
n4i1pE3rv/OCeCCpXZmWFgnm2ixP4yqbMv1reY3bOjCEKfYjMZ4+f43/QXJxJjSR5ODovg58HQcv
DYOex9Hzwp8OE+SRSgFER7GNx5ckT+8sS5870jW9x/se0RT2z7UusOPM74EzzZwN+IpssG2J8JKd
a4DQTf9fP/v/W9NWPoLT6bkUklM3AYBr7WR36xJxV9VmdZS81Naqt1EIud/0scuGJlr3AOXcq6EF
8YI7RAFPbUzKy7IeiGcF5LF1/DZ2qDTZzx/CHUgq0TB9cb8M2Qi7YgtWllU/P0iGJs6dnwHuy2Ey
YeXetgpPcC9Qr26OPWLFkYDVYCIE73ORIRVc/7T+N00BexLq1U9+7fKBKpCBfwnDcj5H56Rt+vNK
XUxliKQwQODF1Ewrnogt4KJHWVa5ps77CIOrAIzba+Y8N9re2HrFkTUKh/pK3q1xAntPGxGQ8NZ4
/XA3Bw8fu8N9/ryfzKX4Qdw/Og9a7sE6qk1DZfrz/fSFex30h9gB5vZA+JYFf/z1HLx2JVtuvjnV
PSYcDhSVIbCO8B4J7uZPzHobJp8x8U3KSVGjNGYsMEidbVRi0JKj/jU2S8EY07T2bC9GWvDpksCd
frWsvZ1FzZlG56yBVS4hcDiRRvxWa4SWr2SYw0tfQ4JWLfggmG4vN6Z2pMObr/7Hhu9PnKhkKAeU
pw9QgEQVd245Cvq+ahtoVv94odJTLrH3WsgydHl4X0OtIif1zNNgkAsBvUNszI6yd+t7rbQjCLgF
gEeLkrwpdVYF3ZacbAfD9kykJ81SUr7KLKp6I0d7qj+vsiwslm+QTMb3hHImdujx0EUphhGeKGOs
6Z+XSN5ql8F01KRSRXUJzp7/0E900bcwRLclWj4tqsRFHDmtnjxulgJogYvorjKnPT9A2C/qQKYQ
bGLV1DtvutLJR14RIHaCPNMxAMAQvxS3Xp+NKq1/GUx0jdYuiSfQy1gqfZq4OydpNvIxERPbRrfe
HDXdRiqv3brgO4yt73osJCobZQ3Bzfbrh2fyZ5qiyTJkYMgNhTV5OnMC50pqro2O2hBJrNYehiSt
mVLXg0XTqgOK02d80ro40ae4b4lhPs+PEw6NqRqLxr0cmlnzFPyQwqACLp5OfuaUcLaECd9cMOrG
B7xzTgbDRuQTeS7wXtC7ZygVNQ8bce/UlGpUzryVMBey7wJetfRu0xjOGjt3XtvOcjuAACvq4nvp
Uw/JpRdZ1YvhCBOAeYbvUCC6mHQR1ze7k8ffkByYlu5XSWwUWmzaudRNqorSBC2ew10BDmIXMVQS
0JspWYgpjOMzvLihIlsOEUt6iAO8/q7BWZfzhvoJQPqkAJalpLhdm/CpwAJEQ9WpT+wg5IhvPaxV
nJVWcQTkzlnL5ng391sHSH/R+85NyNIEgh900sBo5TT+1hKQRsbG5ukPGrlPiEkRy6TJUBocjSAd
uks5tTyPNrDTJNvLceFRJeXfkcPUj8cbHi8XQ3UX2Ktf08TCS2TfBxJuy3k5aQepN2IBOcRqJiY1
fGvOPyjUrzW/6m2smRD49F2e5nLpLvxlibAqYSG63KYq9yfNZPPJdC1+Anlq3N2Hg//oWiWJAI8z
rBfdVCutBb7KVIK+ZXdVowhmN9X/04ce3KXOcepSpG5TVZSxfQ2tSJ+468WOMVQiT6sGkKJ06xw2
fC5x6B6c5Yx8ib7IG/gmM+lSngFgw+NHdDG+pufGp929rlNFhQYmFZOTBe1KfdOJG0w65zUq5mYv
O5E4zm6Fb1BeMzVsfGh8bqlQdIR/Rtnr7ijUc2fe0xiKQwbrcbPyg8QKJDrwsYWYg4RzPWJXff97
jNmXm2wBe7E0ZtnX2LVa0rH+2P/q9FTo63XZT8GRV8NVC/8cX1/2HLIYUVrqXEF03xBLMA6tOseT
6dQoT62Yk2AsS3K6AwPVB3ztMdbdGkl+W6tA8rgwP9EcnZH4AnRxKVT7xJB2LIDPhRPRfps9okys
N6QRQGh69G/rZnPNH/poAzlgfq7bjw9pHYLLrcgpxjFLkv30l8udOY+gxwZ0l5L9ZG1BMgOJRJLR
bZYEnkxve/9UpWQMa9tvVTlFfCJst3JS/WbqvBZTE1GYx0rcAjFYcvFYGxoUpj78YzHf38BSYxF4
QZK5bZMXcBY3cMc/OZFa0pSPcLJZDENLKutZ3xkX3nzzibM/2Vg8153zutidkqBMkyhWpdCaTFRH
uMMc2/6Eaf5Hcq5XBZ4NkfAbXaaaqfjecXME9C1jsNo16F/8ezOTSvilMK8DEp3zO/Uh/ULXXjFD
NA5BIZ4Dcw8txfkmbGiisQTCdWT0xG/bjjzh8dahjGYXA8PXA3SPLPTbXhfYvDl9hesWLPNMVOkS
kmjl6lySpfFvPgIu+1H5UyLGzN1RAMPkDs/PH6VQMq9uiv6q3eMMYLFCatNB1lozSMqFcOFUTZoy
kn5449aZdBQ7Tcf8md1c3I7v+gaPiko059LGGsx1p5t1TQHcVt80s/BlSR4aRzd+XLfImgXh/z5t
NlwXYKMjT6KvSFI3or0zet5emE/eF8Oq0cVOQamThp6JBS+hjq5BmYbpxSCcVad/O69tMS7caajk
wHZ7WJ9A9cFPqo2G3RRmNC3iy+c9f0fNgp8wQC6EZOj7/D1cagDRXMKpprqELnqxb7a7r2PtEVCg
fSwNzrrt692IJr6mKCmybw77WKNkIVEpkoikPceFJsopwYrJfrEbT5wEj85N+ztTt8KGrlHrJD8g
4VhCRqwB2Z8CxzCqEiY/LUA60L5R2Q52ryQ7Gj5T5vSVMxYMepjrjeSaRpAG6hgq1To+K1irGJsX
S31bfe2oG070IQCX9F1imjyehgUBDLPSXZOYGQm+vQFwX2T9WZaJVmrPcd60Xc+Sxa4za7wK0kZ/
ccf1kX5n4xU8ebMYKxiQF4nZkYEd7FREWrVuoq5O9p4BQlYvrlRYatx5dKe77vNOjhNl8gImzHwt
+WHjx7xK+n9O/m/SQO6mwB+fHieS0pI/I6Nj2DVy5ccAPKNT7+BiGOC8+zbjdeDmahIjZ75kQHS2
ufv1fTGjsIPs9uGXimE44X6fuArQVR8XKABXRk4pB66wgIlLbL4JBXcqlcwYFuvls2m/PlSjYTk0
dUZ1b5nlVLN6M8nGE4OVe6RvVHu7cRyHmPWJmE/A4+/8jw69/r0fI/e+XOyxGYEomgcfzDa1OP/Z
fr/ca3WgqNigGOABv7MGK4JHHOvWT/4SpJjRq73fkBjJBSqZ5d/oLqA43CXYjL9oKI8cSNFHDNZ9
UFofTOizLOWDkTNHbJiSwBpeEhQ9qGGDBELJr1VOxwM6RJzKfBZ+Y7vteAkh7AZiDxmOKqKtGYtV
UbPjJVmNIFKmdEXiEgZyOud1nyftkVW7008Q5iQu3LoqAbbWJcQMuG/nbiAZdJtXfYD1BQF1lR5k
WLpNjUCsdPCTq/+L7K2MunRj4VDCG2hzErL9CNL1C85Xtx40UVD38AvT2JbJqr0a+pLv3HhxjchP
Lvw7bI+PRmzCYNU14XIZd5cRf7UrEaf1v4GyCAkblH6KSeYwE2xgoC47cJGodBwpWT12s6bkd5uc
b+5EkozaVM86UmbhiUl2NmPY3xiOZHeXnxiwv0FqETJ3ajG9Dy177UrQwqznPHQXsh73HBN9GfpD
3ijMdHkghPIAKaevsgOzZpDTAdW7sSdUs1DVzDalRn24NBkPdUmtxAJOkwY3zB/4Wmm+OvVzN13M
qFM9Q5IjQpNpNq9kyMleI9teWkkBctms5O/R8+fo6OX7DkGwRhcQ1YHM6IgkpIFwWnL40CNjzNmq
CGncXvbxV6ifrW2ljAwaa5gfrm7kTtKUfbDxzdt4NUb2TiSrBetuAaHoEfHB4yW1uGDwTTlt8Aou
/MvSq9ldOQsih3KaZ8mlQVYxGOTkJmPhNBuF303x1YfjWTJo4EPI3roBeAmThRs28LrTWankbgO4
rqi0dERHl1ojO+fEZ7YwXG2BjdyhNb3KdysZu+8JBpyrj7ejMDOL5F9fD9T04bLq/7lvW2lLG1yi
MHvS6bmKBSklzgpsZGsAwYSGlf/RUyT8NUZ2i+SpMdWrDbS8GCTeZm8JwIDvfvpDI5FG4stpq1zb
CSe8NAE19N1zRH+qNVAwlkSfVqOj1D8k7QkajtPpkiwZfcGRnEEIPsBo713Tu9ZfYP2Tsxa4uTDg
JcR4fGUkdN9x0LB0ZcYm28bmhhYHW/qCbylfeYl0TacVdR1CrUCAnMh46wU41seGxUie+Ya0jXoi
qUMCDMMrj6sISxW8ay+uuy48H4WMyUThzAM8EO/z8DN5gS+JfpOT+o9idlZ5Y/QkERxF3D4vWza4
zRwmr9ZrLf7jJ5NpB8X0++dDZSIftRDxWEOjssj2xnEy+xNh19ror0vI7SCDU3cWY0T8LCXXFnaW
+SRec7ti+8/2fTy9NEmGp/bdCx7s8CRyySEkbdHprcmYFKscxfPt9i+9eQhRr9BhdrRQPWhBtoAC
hOJxaBQ8KKmDC2QVNlLjxDM0o5uF+xixV/aCfhkw0Loy3kxBiLL2vw15IfUPJY+yUE5+utV9JCBL
nNyFyEnoQX1JKyv+tvWR3aT3cFTf9v55UKktir9288GKYbjlNn91IybXHXCEPqI8t0SpOwybVyX0
gJebguaaPERlhYhoa9etQGnjGRrCzbg2gyICr3UMbWQbagl/IJRy9XPfwd6OSO1TJHszmtSpMJRk
0weu3W7BnxTMrcVHkX1waMxxpw36ye/SGPy4h057S2n4eyj7fUVlWPwmdGrxzU/zUAQBGEoj9KIl
jrYKCXg09IOssBGac2UguTHoSiavxW8+pJ7aBocUiEesMBzXmJH8dDdXOOiQmr9FZbOjJxIYH7Ar
YiMEJeEgpb4V3jwRIntQnwdhjT4t2PR3g45+ZHx1Fagqgx2TNckjOJgluuhu8ExwQyiqq6d7/M+l
WFu3fzL7+iUi4wNpGb2R4vB4faU2IydQJF9wjsJpqUdenIyRU/uU0A6SeroeAlKNRG7f0Pmwlawo
INXVQ5hjuTEkIXJIrAkXUu05Mgn9EUjwbIg3FIxJtXQ2ZGfIlJvaS2X1Q/Pe9b9EgRrchnEyH784
BN8OjQ074Kvr5CbMcvnYoIW6B2cmN2qp7i99vp5JPfaUEBhqCd1CxPQWlbH9IwNtVvXpB1F3H2i6
AimSfKnc2foqjNjGfcNV1XmQ9WNjF0vnnpzo2zAdw7dG4QQ8m0V0rSAtFpWByFrU8K2DMPBKcqd/
o/a90NmN1/Ioigy4GsN+Kv1Y2laLrnJFf6h0rCbeAgOYIY2XnfBNXUnqdhaYNMzb8G9lmgtETbYc
GRwDgBeU/DkC0GmnpOwNgXl8bC5S0p1L4mRWxIWFSrm/05lU6U9qs67usHnmBmYUu7E3x3S58yYi
yRoz8+okLg9QjLfXLaW+BeBfUfoEeCHncANSP3urKKR3kPV78EQHx0i3mZSlBPlWQK07B+N3jp7G
hfE9D9YwtWT1GexhaMBB0zKHM4YAi/U9xuu4QpEh2eSf3TzA9+FiytrpFfka3sC4VahKg4Kj5nnC
U0xKkUmkT7CWpu6f3w7wHTC2VVq5ZIJ4Sa0whvYa6PZW+k3uMO4p9FuW3DH9YkSpKPKshWZBRnGQ
FDcBKshgVumyy2A55WTuPqSOs/DRDZ/BkTYX0BkhPWwrIqcFv+rRKVpMhJzlvriPlMOVTZJwNw/v
XzP6joghQwhzqQsBW0rDUKcHb0Yvq9k8rti1RN2TOnNdZPK9+pVNTe49YJF6wyFCeQMeb0x2tiRs
nypY/1FnzzqiQDgnCHwxCNRJ9YCe5jALEfvsP+ySvb5iv0rNt6By6SmP8kpD6NWc54ICyWYSpXwA
Sxs8sOsWyJ3eH7PWZyUqvVoTCyMoHFLXqTSFw/YGemtZ+d4LQIfKiDqMHRX0xDne3STLE6IDC4wL
hS36zTUiug9dfioJqTXvV0TeIyP91sBHo5r19KyRVRbkxfbBjrFvZjAFlWidoBLd6azECNDSIFdC
CFlxPCzNxBVuu4zCEM4FhSh1057YxQaHXlNU7IuiHe4lbURLXUjJHQVxgq+1u77eLcfaTHNjEF81
/biHp0SPH6JQUtzXZr8atTJPYo/TVjojKmOEKtRjvB0fgOGQnEFs8T7J0qfvDNSQbH0xd0Rq3BaB
n3JIgk0KTz/erqLei/0m3S2jVyuCE4qEHYLgIi8Ny/RVi+RvU8NjCUw3CaxKLtIQnsMYEvBCrA8y
b8b078Ay/X6GLYUDg0MlDp8iQQmS0SmIinqk75U5sgpetSUB9jk5qiG6fyKWZa2QzcsFaKyVxP4v
tz/G5Rf6f+D3LGytbvyQZIHq5XjkmFSnDqMZ/MWT86Qqr8Y43J+LfOXHCdBJpN3qkYJR6/K7pSDG
Tl+n26bL72PxaU+cQj3j17kHx853zXcJ9C59GVeobPw+tckUytBAvvG5ilBl78b/taeCbbLmgPyk
HQvzZV7+O4K9mURIIfYb4v7vWYUyUkhg7+IMtLKZKOnN54Yo4eWQAOKGGYzW/7s4rLZeQcrqX/j6
3X1fS+WilUn25mQagiNVY/Tgiiy98GXAoHFWd0SZduhTi+EZ6qAY16ti/veE+trR6bvXHvJuLxUC
0Pukd1NRVJWswj1SsUS11hXvZZyiJw2DLeNfBTRKxisbawa1eHgOcSyk8HROAGaz/4mQmQ232ybU
8W2p2Ym6czu+fKT3dCxKLM+rRFxfv0W+0Bu8Q2T3dCDNRy7BeQjUvc8zu9d7jg8QX/5YqQu5V5W6
eV0w5yQ/wnw32+MLQ8tC/amo6lVLEWEKoReonfUpa7lCiEcOACGEmKHso8zunFkXU6c=
`pragma protect end_protected
