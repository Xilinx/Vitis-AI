`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXYEdg7mMCNTHvUAl9VVnYLWXPJbc9wIkZ8nG8PUYbhfddjimIGVDFPOm
/oFGz+h4c6gpVRy2GLt7IRfhDVUXKHT3MM+d2lzIARUuYYorTtqT3Jm/rq7z59T1gOfV7O3ftgfy
HjXX3zJjb5T71ZkDKD1WXYV4P0wqivJz0DgrG5AljGNtVrVGNv9UAU2838pgc68jgTQncwcU6zMo
EngUrvhbU7Qyi8xb8PegaN+rSS/kt/rcFVKWYYWJ09ASDLxcg51DWfAHvN0ZatP1tWF/yb4QFj2l
FyuF1LDxhUFTYRyzwNsNYvbaLYF4jZCWts/NyDRdPZaZfiP+sy4oGjO4bFNYZvOceDUxWg1CQ34i
cUhzlcUj9vcBVc2ArY2jrcUCmvojGl/+KJcjlZ/cQ6ZvDKncvgVgNk40IDfV8oqpOWhFnMqYp70e
ipW+uTgixb02DyFpi3tSpfilO9qVZWCVvYDkWAjxMfGwaajxd+fwwtQ1zYAlbgXQEaARnaICWfUm
RTY+8oNEU/CH9e8szUh+jjS/H1PWh66VGMB7PX3GVEfVjZKMCD5foT+0rMA2sRIqQyjcwCvK/cM/
mwtKjYffHktfDcOIg9AWea0TReiX6klGv3M2DXJAhdgO072gW0b2jaLccGluPGpQhekYzqWdvohd
YoGUbrLfpENiv2b0bHZTi9m2A83RBUeYf+4LaN1EwecwJxWyjZUXgPJ+DYKi1B0clI/bXKmCiGUv
fkcxiqdAW63wU1rwS/NMSpHHZFUSQ0GdBdwTim+itIIxXNQvKwNdUJojgBm0CGfBi+rDwFjuuFb8
o91t9QKUWcTW65+sKH3jcqP5W8lU+wnQFRKrNU61GbdXVGyYSGWI4zFd3bkJBqkKn43G9m0M23qZ
IhPoudpK7NDwZxIR3VJXhhY/bH8lFWrARvdwc0lDLO/1RM0RbzyJR2XhE/ku0eu3cw1sXIrn2vi0
I9oRmC+aOU4GzU9zQXQ46COpyYZF2rxWXtKYxk8QxOrhSwRl5lG9HgowJyAkvDYsiyKDfjHCl4/w
hRMxia89ZCq8NnTJRmAXX/MVmm32tRw6K6sUmKrW/hPqu0aiJ7IKLMABYFJ0CIrZ5hnQjr+GEmD0
Y6hAkghxLkp7QW9CKG3c+u502mY+X/mTFkWJ6r7X05LJrKw8nyApmZTxHlmbGz5032LtClsWyax4
ok1ECl6VEGl4wj7DcbSUKjVFsKR+92auUTqlg3tL8Py347ldIo1wJGj27R35msrJDhRPSWxaF2cF
ilpZTJ7FhWNQQCC1wSMJLV5s9ZhJ3rK7qDGsozXSsVIbCX+JA0syOPW3nvvDl8g0Ndh9DS/cEd5j
8wCo6sK7g5cczRfYX33bjF4DHM4GSzgYAEWgo5mw/qsz8zVKkKtZJ2L4XQcf7R9ynxcMy7+t+fLk
C6PRraAzbwY70JJcgaETAIjz7kM8/rx7yutUHQ2wfDNcVm6M04zN3q+s83le0D9KEGVM3sxwr1W4
tP1wWJPPk2iaA6vBSOAUv0J3dvaCtlgwSprCC4ghT14ZSo/8aitqgA6PwE0knRoQqOX3eqZlw+mF
CoBsOm7Q0Um+qZ/zJt4Mlp5bYNOBb5FS9mhRSAUguRSnFf0n1PhZ2melLYKelEYxsj+Fjnr5AusT
TA/O3y+09E987YYBlvb0gm2Kq25c+YGR6afUp6l2SQ3roawFb9iOgmC259lDpXFj5Nhg9wSdYHP0
SLtoo/TfbRzKqJhNLEGEE5p7p4ZDOw1fX5WImn1LjIpPk7r6gV4SH4d87F/UsJ5cQyGP295/rIeu
P8tR9USFyeZ+4qLpSALoGkvPB15ClA+9B7IEuB1AQ9gSmCt9Z4J4xNg+AMBuKnTA/F563RrUwqSz
qjgFAXh6AQ6ohFvBD0eVCNaopX40gLmtyUZbj1kzIkxyUpkcH3xUx7EZeOEvADx0LgSiBGWPlRvP
o0JHdK86j6bG39bQ+6E4WJC9qVBdSL7jBeUf+yhygd6HF1/zlhi1Ti76hAR+N1DS3ujfdcYCw3oU
n2eO6lfnacnDqNLNBDOVYq/CQJNXzLV2gUcZ+ZxlMZ7f5aAnu60XY7ZCKqP41Irp7JVx1IiK4q9W
o9p1zAAmj83hWtYDKCjzvHBTDnv8n2cDYSW6snWZkeNWqQdmYtXJY/X/LhL7tu6jD1Oc8t3oz1gg
Ig16WEtTqBWOMzlnzSc2Q7q4anbVrgCVm0ebTqK1yqDeAFAo85iXm8kaDy03eZLyuDOF04M2607B
rmIUmMoB6VdLMpQRS5PEFROeMxdpV3mWApAexjIxn+omspYdfQPfEJ3ew/AkZ4IynYiL1NdwCPfL
V4FdVb/odLPMeb+5U+sI/eGYCKXXs6+O+x8W18mhlGfN0SW0QlkDGxl2qaSQhSt7JSGPpnEg1qEV
mYb7yFp/7Ja4ywYbn9ZKyyKcCMQUL3sKwjjn3Z4JwO7SEbzA2DZsQE+r28QNPUyggIFQu0RBMpeu
JQ3E32M81HP0R05rW2cag9mdaqsxUaEjre5g2/O3w0iRzZPvF3LTiOA0vmT7EIk4rx3HoG2Pxg2V
fv7qE9FcAx9b36wsJ1UCdt++EuRJDV6CJnlgZL48rdQ2lwXknn1f8+v/1KhasXsMSS4oBG/bZv0b
FajzBSXri8w8b/noXbNZg7v3R8oCBTesCL/famH9I+wrGHshuRpZQf6Po4TKm6lNezxVEHFSTBwV
/sGXnPaPiWSiJeDBdU/o43iypk8NZtoMR7w0AmsablrBUcNZzaZ1valqWSPn2Ze1X2NfIJ2v6ebl
NTzoMbzoWD8MQo20O1RDCOvviLQrhNQnf4IrPriMmr2swQuZuaUhn+5859jHTUG6A7MqbIUT1gca
Z0VPNx7xAFRegVe3jDp6U01Ws14nlSKHqXaTvFm4c1yVSnVJm3tIaFknv/hpzYSloijeECx/E086
EJraxx8zcV/BcE1FDHjxoohAMhJMLz11kncnHpe8sdeL30dxLZtV5Agti8idS+DvDvDLxM/k72xC
hl9n/tuschlK7/A5mHQbdXMcOxtBxKYlMpIz88I0IEwiuMXvDe2sq/l1WDevRpdsVIpzw6g73hUZ
A3G/i1xG16k/V0lPDwxigKZVj53t7udB5QfUAE/6e1soULOSVNmBorxMEQuZVDYGeg0pnfYyylNS
5l5V6ZFN4RB08wfZrIRIrPPqgk9b/0hTZaM0zAgavGdyNtUYJGALiYM2BLtrtd8/4jPaEShzIsh4
3YOC9Gza6zEi6+HMV7Jz5ORBk2kLTmLor2JZNVGzOUyziIYYCaPauD8XX3lKxdbzHRnhyqBUzB4h
ovTWc3ZHGfWYKZ2qb2RTMzk311BdpT8IdP/KoGqtHnZO7jpVOdHrsgT1T2aI9iEtOXwz2dp7alrO
aDxt1Vcf/NuSzHijlHipyT+fSa/pOkBuKxZLLWfJM0X0J6UYXPbd2ZxGR/bskAZBq2AAu4rN7K2k
k1pUuLo/92+bWBhIWbCeNmRaL531UqYH9JbmlhLI5LiRHwSfhYeTeGMHw60K8PE5/JqlphcHB5xM
0sfL0xCZW8IU9PCi4P3ZkDbnNsPPN/NqPVlgbCs3LznKdmvXhJLwm34auUxr3mp1DrY9Aa7MhtED
wq5ZGYdWZMVGlFDavunVkkgzMR+U88kABlAnBRUlhAMZKrQNoAEOx+aUpbBvFzsISSlm3Q8OYJub
01GVr97ZtjLiDy/0VYu2mcsqYStSrAut7fV5uqGA3FSHA+Bwz0Na6LxDAA2Kf/9NCyzXmJ6PLoRJ
MK84Qe7W6AmBniV9V+HtwWxVAN4PL3CoMyBrD6HUOhDqzJWmD28kVbsd4LyoPdxZZGbLO5nDy9Za
AKNCGWWjPUVG+QX4fntvnk0hexN/i3bwQxQ16zROiHM04aHfdKYAvOlJrGklnimeaPvwAIRsk1PW
65PeVmO+ezKnHjFfTTuWWF9ku3Y+PucYjOHTJzrt0d3YXRCMnXRisoiX2PvxVDP2cfT9j9Nh0yb1
XxEwSp15PRLoY/9ke6BW/+FxbxKzGI6MGSbWkJm0TwTnRzC4EBdJI3oQoz6JOV9Ni5eUF8Ud/Hon
Jblxhv8bcctWq7wbYD9PYvG4ByzmMCZrmQbvbeTS6hXHCABw71jd1o1ut94Jkjejj7FG7PQxFHpN
jWyRkYGJR/UFSc3FOGf2iMcKnkBtJp6b2ihQbRqhXur7KrAmLBpkFZperrGRVWUE4aSrzyrkAsgu
edXknDUDl9HAWDlCLHqOajgCLORBtCMqFDoha2Sb20KTU/ehvHCBrCsRCW70ctuAxDv8c26B53xn
0CyfRzZParEQsBHcct3SPE3MofB91rePaftA04r4jaZlMmpf7n4J5BpOB7LZxozmsDXkOJ4pMHVD
56f2iJZyNEFdGCJPpd+DQp50aqZ8fZoGzbjE2wtfUfXe4mQENrqsxle204i4+mJwrOGv7i9v0lxK
JDnvz+brndF/vgMuvgnVJDljhdh38lgjV0zgF+mEkTyhoeF9iJsb2w6MUoowKm/4jFto1PNHNP2n
Eb+ZE2Qv7jkbpk3HWdVjoVYkTjtQXOVvcHzeockPzm2dKwwzymcsdW4pDEB7zSK2dfcZa9UDXCtU
jTPRHRTZ3+t8vfAwpTNNsmh0gIhZopYqT39wSbj0baxr9m8LmLlvBZ9Zptv9LDvnBGU8+Zi00Gqa
Z+xVbQcYNjQds2yS0rANqeraS/6ZuAO2PxjaQvH1Ug5ca8LL9Wy2hIIn6JNCOhVMomnbpIoifZmB
DR4La6TJV5BlqrN2X/HdFuR4DSt1WcoPoiPbEPvpd+fRxwO4nVmT0KWexVMsg53sraulLRqV3ujN
DtXzbnySUVFTG+5Gql8xW/EtLKYdDTX0SLgGD1QG0eaMrNkY8sYkqKmdVaKdUMigsozz/QnzVlYe
HcHGxvV1uOzZRIApuIxyzMLdHcrDMomUKj7jBJIKqQCHtBb58As/bh8vFU3NgiK+G1qVtvbSRJhu
3uCoDijAhcexGWSkEDobOHpaFzuhOxCG3ZJ+KM6oINqrY4B9sz1zxDu7V2QJkPMPQ3kdvfjt38Vz
/PRkwzo=
`pragma protect end_protected
