`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16704)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT9rrfVTtnv6Z/atBuUOrnyXqzLBAxGGYaY60hwY/ffGQAx4GLVwE5nNzZAdz2oUeP2NIOTM
dRu7Yzz/u9IG7+ardU88KQzL8iJpAAUqRG9WbZ3iK58IZP4WCVIFl8NwTwZa+E4VnKdxd3LndlkI
fa9IYlq7YUCIbeMUgUUSIt6EEuqBE575Mat/nXRHgLPnPYgsPBYXXxA65cC3l8Uwo+gbMSNuHwbS
sk0pUFxTtAqN4Hz52qz1uC/UUuOPmqdbQnZkM1CjXi8MP/IxKiUja8esgYLkfFNjNNnjVXogrcbg
YRPK55oowzQnweeSI6isM8P8yMjsk8ZkgISGS8UUYlgXoWS4UEfAqzPLDRgZ3YzBuOhTl9SxHKBd
ceBTmdFkkoZJDVcD3ObeJgDHiFcUPTOOuIv3MNd/7L8SBE2CGGm1MOh/IASutmTNk75uiETd+bRB
IKJJBfR8RdyWjfsofNDbpZcaNOw1Lhd+LfoGQJ7DVMW+9VPPE8ESGcs2prjMlDESSktFIz71PVaj
bCDaVAfaeERQOdeLAG2ifhPCoyqIreMWwLiKCKQRslfWgxXlK430NNi90giNyT0MAjf8CaS3eSi7
QxJYsICL4tiFXqfCVH88mi7S9Y1V01LEJzZi6NCRF0LlbfnsxshfRIJDesRcFcS75VgWMduFSzP5
wcodbndxUIiDA6eSYK0aG5FOc3khE94l1E8YSr5F9KbA3N/pqBUdnIcQwVF2RjlsO6TscZBlu8E9
l5ikQk6nKLN0Mqa5SSOvqLhniUKftMwyfqRd9s/bE7pB7qaS5kBJ2obFsQir+PenxSSQPQLRZsl3
kNeTClJzEGEJT7hfq9g0GcmYukZUo04SVYJ5FE9h888wrAM//mnyPQI0PGAH/yp9VbVyVwPkG3/Y
m2x4yHYCsWFH+irM8mcrr2qc+L8iyCUN47iNEuooTrhbdp8tHWpCn+IxahokVtGIg7oNmtNInsu0
NoDCS2he3kdgGZV9YbeaFdZANMKiFzw08FspdCSoFaAlela8vnhxVHxrbBYkvoslcfCTnujVWtUr
207FLVxzd2GzJCoLjf9pmIO+IIddnmdIZ7BbARZBWxqubkd3bXdve+sbk8VxZW1SC0hkd1WNg8jC
pQAuoaqRhwfC8beiHqx7batdnPcCTmaPDLDm6cQHJ7tbBaum9WMOTqiObgZkn9q30mVysMKc4Mfh
SgT9Z2r38SxB5KSmVjUCpJPzWLU25xMBl6CpjVPOpRPn4DrP2y1OLjnb8vFAKUk4MePfTcsXz1du
+MHib2vyOhMaay7QCYpN+T+QXzplTr5ZppLzHVvOgFw/2O9WGFQLUOQUTcjb9VIKu+ZaMaxLfgx4
H7Ez7W2dhvQao2i6W7r2XTS6e8kNnKItO0mLdfK13s4K3g+O+ZDirpLJrpat9Yn/qvernjZ89LAz
y6P2HY883pFJKSga2mZNXthqs/MdbsqtP+HZ9WQMV5gDCdvIJP8LjNUen5ph7QSCtD5sn6t76SL1
oqjDtH7ZwBqBNjMB1SvVwA+6d0bn7a8yHYzQhh8Rmt682LqcoeOFXf4f1gdD06ptbvRB7W66LopB
F30kLo860RDOX2cLsYkSaGHFxKDzRa9QFpzUuVzBIP1MfdEL8zJ63+bRawKsuk0WeSXvWgzz75+o
6Ba44VVGdpNXx5cBMcd+S76craVyWsAR5+PZIxrE1aHrbyrKik6KFKGQOpAfyZPZ9Y0jRnV3B++9
P/tu3Gy8h14f8jrGKaHHL8gctbPUuKREDzHBZ/Z26qL/GCUOa3E0jlnPhp9GJ6V9eLWgnG5A9/ze
iHCisaM0Y68OJB9wvmU+NilFKU1e/Ety0WZCzvyh+/GPDKxw+tt6alOuGb91tARG6BXA4bWLCagX
4gJZwi3TXTPXHG4bFheFNSVGQWtFeJOwZFZa0QhrKASpCh2gMuAglQQn9SU18f/QL8/7Rb254QOE
V6W0g8BpIpSCIael++rxySegcz64ncA0MASFBWJhZ1za0gZrXR1WRomRHU2YS+PZ5F/t+xiqVJTG
fyIDwIqGH1khGIiqc4ErOeljtUfGPBQBv7vsOQNQnpUinXpClUzTNJFDyu9GXw+lHmRDmvGRWy8k
Evf1S82lStXKOkcjDacX5k1S1zWWCtDeA9QTT1YxfiNaLjXVJt6oE/sKeXDhb7livqfZJsDfVNKr
IrSTKjCzZqL9QSCfnN76OsQCi9puH3hO7PknQm6Y7t62bp6eyaiTBQeHvEQLKIp8puvhYElVGXGZ
JM+qwsd5nxxnALpxsJsSdq+5HtKJHN+gXXIERdBNw/a89lzAYXn9aMFIXf0gRZAGCR8Rrh9QT3e3
H4KL1dd8+40sHc96dmlggqLWlkp7TpVRPV3XFXdxslEgVLTiNkR9tX3Dryd06prd9M3Tmm9n2KG2
mj9UCUCv8QgtVB0CQaX1dLEU3Z5do+FmSJVdCJ5Lyf2abFqG8KDCHKOw8yBhix0R0bajLQAcwgP2
8V/Gadt40LGjnORb6cl2r5dCrJepODV4LdnskyDcmREg9wNOvkc6a6vVSMtGGzO0eoYjBh+75lcM
VR1hpKkW4vyGomN0uJ8IbvU85MJCe37Kukn00OdhXT98hhPPSwHu5aGIIJUHeg0vNu1MJ+BlTvm5
thsSIRAY79dbaxOOdfuz7QuQ6kg+DcK8mIKUj/CihlXa5/M3jxet3DxmKuoVMY0KaJghRTEsXoYn
6demjk8XnJEoR4iN2hfY9Rr814WTFTzx7WcxwlLaaKhYXPJKWuDLpxYifZrG7kIr8uuQuBZ1KsyR
DWzJN3KCkrPqO3/2CjVWGZIUyh/46WwqxkcDAOS6uKpUMi+aprw8BiTmzAvmHBgEySyLadh3WIXW
SyVhe0UxN9AiBz3ZCWXKMncV+RdUD3TyzquzlWdv+zgBqKuKZquh+8eiZDdYzhYw7Cv7JOdYLsZ5
mOS/lIasEkNDxbi93jKrKaZByD9NfJs4T49HbAG+umfFzy2jFmjYtVc6tU64Vq8BgHlQP8K1kj9q
NP0xfqd/d7dDYf1PLUT5vBgVw/UPxDPBxvo5gAxJDzEi/1XGPZvd38KKuIcejMar02AFux3d+3L8
nCjERlgFke1IH/WCY1CZUk3YCvy0gogqYz2w2Dr1+ZyNtnywy1LlcmQ2hNOl7PQpiz8uWc6ksULb
Nkkot6KsaOqOch4/FszllnQ+8DjVAthGNkqcK2Au/O+uokBHQ6ph978w9pSypaTNMdGsgnIeF7KG
C9Wo7qTXshn/ax67ejeism2V1RX5sTQct6/BAGH3LLx79+ssZTIyKsd2trIUFBRA3uNNxEeeLIyA
7zRzSkTFkbexxxzsKWYzuEWh58IK9EV/iag4k13x0Yml4Fgd3oIa3urKDnB+Zcx6d4CrkUH/S/7h
egDpsym9ArxuO8w1sT6aih8DZg4PqnvAaIWEocvznjME2QWJCsfIBHKQ8P2VTu93FnRfnGP1YHr+
3ri47xnCpCctoPoppMSGKF5JQQPM+nWpimP1Bkn6nYPSrzF0S+iDoIHBxNhkz6E2Fs20nBoakMVC
7qECSlbooOYxHeqAkAk4zUOPsTrLx6rOLrrtjraewrshDztkVa7kqlTxUSM3bc3hQcaHL8QYx8Lo
hPzEySUtAYUNiuRS4pfSwdsPxRUljoWlLpm1ay0PWzUayK5t6gZtPeX1MxMkFF2yx6mqw6/n1RMX
beA0WMOQFu6iNC72JTsPwZnb+edfbF5HUWP/ovHV+d+kPP5UcavQmewTSYl7UM1WoSePLdm2UMJ3
W+/OGZHxTmLvqcvyoXhA0/earrRO/MsFKxwrsLYnTIlQH/BUF5mMV3PkX8k/bgP6xvogXgHOWtxS
LJXz6taG+L0XEL0dGwU1RWxSkrGiryhEmcsmqQmxzQ20JWFmut9M1vDDl98pkjlf3b36L6cQMjSB
0rL/YdMrNS6VD/IMksZisa7uONIDDHxtNWVw/d7KrChjJmS5FrGUBkcFZpIa7eNHZhcHhkXsl7pS
nVZjlyaMUPabHIxg8Uld8FyHJOd3tXnPy0kQudXsMaRnqicgl2iTFP+1vn/gnaYfXN6mtOWAURkc
LYtLf9YDfYS7YCSshwH34H5xRE/WBLF2ZBLeEEp+w8lYrJbO8aDLx9TuvAiv1YUtllYjAP1XNbJN
4YCCzpWdo7K/tKCkh90p3JQNQ3owu/Zq2owIH+n+xIxMxe9vwI1GVthL19LpxoojsA9hhCXtEN0U
9225XPcb64Z/ZTrZ0vkEeU2wLKZzILD58LzhiymddxgeXcYOMDCQcaC9pU4YVwnWQTYYbSHYz4C6
+kSN/33Jn/IMzJeERpAnslU8uV1UqIwCFWlXzcnfb2KZi68sViq5db3uX+dQ5qxhGpTTow4hxlUR
SgBS12JxvyWxX1r2zswFkMKzg8l4nCRAaliRqiaeNqGd190Zsd+EZbSiGISXTF45bGXIAmj+Lf93
aarjsehvX9NQkIK/AgHWCgHlYALXZqKQabTsGvXkqlqNgQFZYZhvT4JeA2Jl6Z2nEC126NeAya/5
INkhn0D2dEpsCdILOugvZ3uPIipIsNCfD16F6a/8O+8+EdIoW5RRwg1xsFem5ECBY1zyugKEDdmp
te1JbYtjz3/x6B59gSp/PXAiHGseMAHkSuabPe/4TA+pyRVitjDT2Yxc9ZKlIuskZKxtLfCbYBK3
ms+1zC29W7QdGX5GMh6FTyrIfIgO43PpVkFncEyXcjR1VfDS1E7TgcqCkzHDmxmV660H1was0lOF
1FWJRPztWSBWzlE0F+g01XvunD25dHg+aXT4bubZfx42TJFotg1RFgiWHOBefoYBPIpBugvXQXBD
6n+SAti0ONwRiUc10Xf0ePpPyJZ0lPuPFTRcE2j/uFkDMkZYHoZtSg2XS1Vmdn3ZD2cWVWs68SC1
cpVuz02dylK+nEIz1S6wYNyxCQ4K1c4dVlDN5D42vtOIt2c2dB04MScR+h/67jp6kyNdxrJd5hgq
Mrub7mB6SqATbM+0e5QUZkeSdPrLHPdNqAmdwdey3J5IQ8URgpQobqbCX5ve6yl2o72R31qgb9tA
tjJJKmodoYd2XJYfn9C2LrpNt8aqMENmHcm0DdUO+LrBZ2hplXcjkM5w2P+6d3tBnWTAD6DNidfp
HbUCf1JIgZ/pvvzl24viQyBsKtu0nlDnzxzmGDxGxeJeae8ruAANbfkPMcahDKykx90Dst/4LtOO
WDfyFwR81r+8pqGWGB7RvrdHfkXHzdjuiQjuZPFbzrR/5z8VS4ugE3gcvQlC7JuMcgmRc+63jJdO
Tkxw+w7QEv2UO4LZUsMQbt4aiSfVWbvpF3YVLa+CaLneCKII4IiV2TTp45I34+MuSq9BjhVgjcz7
L9muegsCUhmYOUCYmSpFBs8cBhLVc4n+77TQkcvjtYARNeR0DDo0fW/e68iNfqokRa7T5s+dv6uW
uuEsfZvRegrgdTq31J9a6dPrMa3abzThZJsbSstEWKnFLVdnQi5Hup10qHfT8OzQoMpPmPhGrKwC
2NN1PsL7A91dp8F22eqMm0QgL54TLjaqEAV7w0MK+6UERfDfn1oleTnvugAAow8CDNpPZJamRdzu
eP+IgU/UV31Y15Nzkmi7FFxZMRyWlYY1W/KErA7rJIL6ywjg9jM/VL6Vw0hgQPQzUdtOoaSWJfRM
3f5yaMeH9HVlNAs3DGfRUDIHxlHiKOevGxcgYe4H/vQVkoKXLDutiG7KfxDSMTVxT2g62hAfmCWP
RXfKIOKSZ+D7rYZ6qttTNWylG2g3Vu+1MvicCI4klMRS+kUinVczez3E95NpwohxWPPVghg2J908
WZbEZJ/jxUuBiWaTaxQKeJsxCLiEz7luUv8cbFf0rsmsBX+IRgx7YHWue0KkdeLZBNQ6zKD5Gbmc
74o40LgbZHv9X36/9tB1a7u8zuqeHY5y0/2GF0hk0JecpzswRbDJ0yskGjljdd+xBY8Tfo4B9MUC
BJb2SVtpYLpGFPZmmKyxc0CRc/s4KRcR5r0JEBSDTMkyTFPPprRQrL+tmVRW/anjPAg8YbsVjtSk
S9lXwfo0S17+8AUgBC5EpmU9Myl6Nkc8YmNQGr4fIhr3uhI3f/fO0YSBCaM22kH7Bt9Gs2nfZcL6
tqGRt/eQ999iDxtrEKIVlAY2MRj87r1q276qi8gy66tJHyD61ECEOlvZTv4DgKczAXT3ZM5bkF/E
szXnNLvqDDMrgCmIT/MBmLbvybRWf3AyfiLS+Z7n2NFfa0bJZaTZuOKxkZIsHfXMydW/Rp47NCsn
sXJ1FzWGKIysbIiJOZP7KwjuEccHaWcmJxMGKGdN8B4XKaJkEcPVRaPuPANGKTuKYvHEPdhS0Hz5
x0Labbh1P1E0xBN7t/wtlO1MMB5/saGa+bMfAHE1Qy+b/j5vPVAfG2vegpdDOQ79gm1w79NGxs5l
GdIsZOsaU0BTkUWHAHxqiMcBE9m7dKOXUDF/bZOkal+FIzfAFifcUJLz1+TB8VQ8e6ypvD6ZQhHs
5Zsn/N1V2L78zuGqgfVBJzrTeA3RhUGzbuY1z7BKj4LVeh2r8Feaw3Iv2wLCskhBXFli3J1/wIdE
yXnOqBFhtqqT9/baisHtSqmvQSCjzqSs5QnUtwtF7BsH/WnBvoRX0xcUhvW9adA3dvNDAlTK/1xp
7TFAjAh8hIVIxHghNjoMJMRuj6uTuhdnZRzGuFaQ321zHNBvNEyYxGXAFjIhagGsjJ1q9tw1G7vW
APrjlWv9d+e4aMqvPsubM7tIv3+wx07AsNhfbvuKZdZZdKVbdGRL0YuRxqtAlaVIx14E2KSy1Xer
S1kNhHf1QuJfWZisi3a68hhyqN6/gCaP7wzR+/lqUcXZ1LIo27Qg2goMna4HN20xyZbyHHhZVAup
2/cRv41yPBFZceeicwnfg9HzpM5alCbipkCZ/bsgfgtS0lEaQdzDCizMNoFEypTlTZRNbOyb8uRC
l8Jv6LKT4N3JZotoHld3pOahDw4sSAoNs49X4AWM5FmLsV5ztkHF1Nq+ZEFE0ua5FxboLR4inPMy
ZrXuca0TcXrn12eDG8gH7NsQn2yRnc6FGGwl/hkRonJdmHXud1lHVoNtWDTbaEV8apwoP+PhE1+j
8NEkoc/lt3PHqEzmvWDl/mHtl3JTBF94SP6pOkZIoArvTMpP00aO5PujG1ueT9bk950ODCfnPkUi
tj0bebKOH9v73ZM2+t8BECSScW/ykn8lPTihpGE7lD9wERg5eOXPnklVT2wumbnoL1m7F82/XA4m
bOMdiLiLlFEa8EFsZcBARd5H2lU0qrpPwpeWztX0yQb4KIqYLNZltX8sGnh2veufiR3rS4qybqgK
c7Z+i7tTo1uX0DRvNZHxlOyfxbgYBwipp80tYAFXqRocg/EutkVEFfMeA/AvpPcn6Y/X754h4yvw
0dY3zldJE3y/2rtvAlux6ymUHDPmO4Dj6IlvW0FUpmMUtiyipgP8UWm09dekYQLkEjioTO8cabgO
1KXTKDDwexTdr4+X8FlTedXTtLy+aI1NXwRSREiM0khVKQJ7Up5akFzp/ENGYmGLgMczUumWCtRX
bYi2D39orNT9E+/HqPAGUPl7nf0ZaFKByrO5l2Omf607TV+vyKZKUxFnjqhO8qvQ82Wq5Jusujtn
U8i2Ll512AnO7fZsec24zzQLEdlmGEt+kBeuJNEGWxECzW6XG0kzxlUlXm3I/XapMSwkNJy7w1l6
ggud7bZoqGwdIwiS3YXlwbTpjZCWR4fXihW3kw5Q/sZHQDdyAu9c035Rkw6nTyYkxUHscHR63qwL
5czCm68ZWxh0CxMaDN3vhaoQNFivaV1AfK9pCpflyPhd8vOmAtow1RaZs0x9d3sg6ZfgA5x0v6qo
forQng0IFcqB4sFjLRkqxFWcq+uKQapIcDC2L30rZPdQaOHWgSnKM4sLAKdsPVFgDPqfsConryw9
XZe+pUNBzMi9/rP2yYbNUbROy6sH/pEZsP/2tnu/qpiScaHmdw0h+o0ANO//peuN2GeU5414jcTF
i5WG6ozf6zkYnCMDFjtmFVGhyky3nqfDMqfk//ymraV3F+3HrW4XedXqktHLQDEFjERobWVni4Ze
m6AfkLpSiJNCDRaMdfJTTPCYcy1b4vcLSo/jKdvQvLNWj6wY8vsKJ0ZEZ2LTz2Zk8f1FB3oMFmeF
hbjqMYt50UQOr7MkYEXD9PfUhw8/MafrQktfLdPWyqgRnTER9Q5xbf+TQjeSjcvSkg8AXNLVtWxH
ckpzAO1L+daiueLlSznPAUabNuY2ivXclm+WyVBq0KViRXRrnJNAaDWxirIPd1kXViyqIRuqbYw1
VC5h52++3gDkF1k68GXMnWPgoM74qdCZIwSTjqDe48ybctGpJDzMemuUsrpriUesLEH4C5fYqQbe
34FYBmMIyjIZQkJRZfqq/pXd5/p0FmqiUpOnsU98gLKbEBoyocnpRMShmjuSb6Zsfcd/rpUW+1qs
UOIWN6+TAur8LM2Kae1v/r17Ks2wWdymFNqxqrh4BJr/onX3fXQIYWgLgwbjUBvkWXvxZgZY/SOW
ZfTh7LJ2YQC72dgf9LdG96D8gTpwuRwr2XwLdXh9K+1lku9FadD4YkKs4xychXnZ+NNLOIhyvstk
yUvQyWtznjXQftMc5Cer2g3aqBHM9zoPOTa62IFtckNGaSrPk8eAQkL2hfaDVf8cX88c2lVBDqOA
XaPjI4c8TJYSg+QuhH6CPx+ri68rwPaWk0jqMhty/MzLPHpGRPs6QWN/pqjWwY6zep03rHg3OF6k
NqREwA/GA0Bq7Va1k4S9VPukXzbUAefX6YhthAOqz5ahrdJwMTitm+H1jhTGploAdK2HSSdVbPv+
/ZnQR72gT2lVlh5YcH7VqkGSwee3c9i1k9LziiN/giBF/8zcEYtxSUcolcuHpYExWCNg3VKTPjMl
Lr873IdXwe/Y/h5meXb6osx9orFv/J2g92QZMYA7X1kBAsEdATWd48GixF2A+Sm0SOYmNWwbIbYL
Za+nF5wMEkzsE+lsNg3TLpiUmOJuR2dppzuRSjt4vxyWrxNNm1pK8yhwcF+DxNisA2cp3SKe5yR+
CJjPhLhMMqsWlBUSu0pdN3FyFr1ziGl5exFGWv778OKZ7Mz4ISGn8R/G32AMNm1mKViSp9KLFKQA
JXZsBEC+s/QD0iwEDb91yd71pHEmFLrap4wwhZE6Vr8OrzUG7zwl8qEfncz9Pa7S2ZttI8LZ/q5L
9C67nfsqDjkZfIzgAtZ9DpcZRpn2PHK4N9JshwCgRwl9zwbDO7QLod99jpq+kt1w0Cfb36bhAQD9
ou07usfOgCFn+lT5JpH81O0XWTK/+Aht3Hq0SNZlbrQ35oXoBc3tR0gKjLDjrNfnUzXXTQbTg0qG
nBxsxjZUevhDSSCJaopFPIwfGO2sngqvS3rKFYQW/Lja1Xp62mVdLSL3blDenxl/cpLcbboDZ++y
JkUkaq4lPY2L7BJEVRQu9YSh/D4U44aZS+EY7JUptIxDu5GTVvd3QWssEgRBeRsQeAnvjpbye8hh
Z1MkplSHA1w6ys8ywQIXPqvKRDCM7Rs12xb9hMAbyG6DNunM7/JNLK0cmsNjC3tSQaroUpFHfpWZ
SUt2Zwl1uHwDoyiT9QRrIMfRP9WdR50GL6hYRcggETdSWDLrVhKcJ3DMDXRZFZM81xoSlRpeVQlE
v+EabLPOeiTOKTFYuktO7FrXns8NUxIWFJTgUnGdDrQlHst32wWp/MO6bnMKRrUyCZPMBmUkEKAg
VrBWaB5pd/tn+BFxSLXRljE1Bs8zM0QFpRCBkRcLU6QxQRyp8di3Zn5rPbwDjwjAR5MaeWTH5509
SrWuSRX+LbtSR6f4KNbM8QSuUpir60EGbPmH8OhoPW8fZMbLW3D0auGE7TVPc9vshuZ9grCNVlcV
0KQ/DlbMB/lxnIgJk6mnSUUANyZEVAxwEknKZ28XDqlNvIxsaIT32zu8m1DYcq7DDoK7mHMWL39q
1xwmaOC1t/nSi3m15UrZUfH1OxW5MaRuKKes5nf4Z0/LMjUAu5PLynmOefTtosFMYytSzxwjh6zb
y+k9B0OxxWkxecJ+6rnD8VOkcQVvXMoejo71QnW+7QPLAFDmq+4c2dMlCTPW17itNSVGX0aFXnS4
GhC7bEmCjWbD9dCSPi11eXXe2wvLsUod5PX0piNg1aJ6NCiuWtC7AECNCt2dphlWchjG7dYAJ5U7
7dDerV01z8ti8XpyDNxZ6KDl01KBsdSAJ2RCSDb5Lzp1hUlFaYNm1Y0uwPBK2CFAtuRTQFsY20TB
Kt9xXwhdkyLqcuEeV/GlFOSC3nCQBevllr2M455/rcq2nU7L4A8gsouiWtoX/8V2nBc8tXEdi993
Afj01bRwMoZOy6ZRkWml78fnzh8ZUOvLjxYgY1TDcfzfysAZg+MAkImCGEzD2QDHV/QeeQ++yLvm
+876KNbAr6J8666R4UZoqmhWhiIjZXsHjFW/OrKJ4bGlPpYjZZU/Y6LD04veIRmNIrzRAXrFFN5S
UVeNqMY6ZfrA+zypM2QZR5xbxxL0Z1Uannu/4wRCyGQ4QUofnxN+rBHVXOP2zVlnjNdkppvyU2ai
rPik0BS3M/tL0cRW+aDWfcFbgYe2HXd2JDfr5IV8MfJdD0+lapoe4MGKSNRurZMbPq5g+xGocifo
Rt6Q1a3u+RfRUyQH7qsAnrkCdmbSxqnLwUEXoQSBfMGEftPBNh9beRWppVCguzdh/9wYUtLcHZEK
WaZFkTADRM35xTLJOIUQeMRyEyn4SjUvAIHMNVGp49bQWPLQSX580CjkjmqlJ5l5kw2/H2pE5jv4
KXNFAEeGelXX42k6+0JI2BFeVHUp0Uv7ikLPsbjrAV003QJtRQ4U/0MbJJ9dYP5RVkC5mfW1t1r5
3wxaEyium3iKVkb98EV4X09dTyPY9yJQKHeklkgg55xmw3N5EJrB8OhSFnB1IBLFSid/TN0LoWoa
1i9SL3OiARucw9ZUmBLGyUyaZsufmzRb1xm4GIFVwXrwTaDUk1ikzVSkbtxTBOypWYM7Cibxo2A0
P3tFkhZt13H+X2z3Wb3GdbGuA/oT0VyiIQULX4WyXK1/pCg/Q9krwKjMHcDkf5ejG4N7uYktZDO0
+95BQKc46Q/J/mg50OUdJld7UcJV6TBg6rg2m+1WZH6BtgfekOKmWC5pbWyLKVIGzb5r+Qp89eqj
r4IZ3n2xojLvff8v5fuDAiuLAuW/J4Q0YhXV1KMTf0OVPpB0FvAsyiLH9L3A7NIwN5e5TEk1JXEQ
81IGtAvnqDQIu/i92b6nNg5B6GftQoz4sddC9Yr0441kKJMoxmTc/9hGh5SIRMio+53c4tDcmyuG
7HWy4jUnO8j0KfOvv6po9SgPrdG+VKtstw97VBnLLJYQEBMxqMnaXR/Cmy07OS3YtbuFtzeR8MlN
VM9COkM+RfV7jLYQMXFJ8442dx3p7R/o/bta979Wv+1hUKdq6E5qTs8r6MduMvU3BviWjsslePM9
BeaxA6bJR/B3myylbELjLxXG5tYF/qEMS37aXuU+tzCqhpQuUOgztm9/hueIxQN1+QKndUwLXOHD
m4Z/k0JNKB8DdUG3m1nBNczrmIhC8PILNFhle8aHmKbDIGpxfwg02aLlTDPHgvAz8i/aqcI6Atza
4LSUc0RJOy+IRB9sNM6JJLxkoU/tdLh/d/j1Fmj+Mj9CDY/7Ta270CPSVaO/te/qDXWVUlkLeh/6
/XzOZ2Ms1pjJ8EsrH+05/cduR3woMV6DKJMw4hujsVA+3U7ETrgW+V0/G0m5O87YJtfpfrbLbJ38
y6NsiRYEpM0/8zjAGvjGGcufLm4IVNg1WBK1NPhN76b6ecQm+RLGf6tkYL5Zv03+qpu/el7VaFoh
/77FTSUQczlZKZtu4338NRB45RQ8fiheJEK/UFNxn89CGClWXvflhRZdanbQPpi4papCD68RizSo
of2bNrlE6oKRj1XUtFWBlKhUEdj1EbiXlKolgBrSsehsIziqWU+bDYhMg+v96b6RxGhDRAZlGCZ3
Bikh6ZcHrbXMvzhEcEYx/v3XwLhXdkOmcl2brPaXGbZG3XmzEq9XFYqaJHJqtb99t6l+aij0Hg3p
BY0UHY0feyB47KMtCs7CIuPSrqWwP4IkpqXNQMqmDhhB+An6ceQCwzYa4ThuOeXKDb3/evtL4CGm
IPqm/3uycYUb7ktvUMrzDolHvKNXttKnI9W1DHgwgKhxMcP4em1MQpq1pxR5s+YzVOLYcZ7M86DO
2qvloLFev4D8qGlD054ZzUbRDDlYy+KwlMO3FjeV+j6pPiE6lDYwU+dZ8GpZP8QxG8RSimd8CIwy
TUWV+Rw9TG14x2NQXTAA4IwDUvOhI9kWNEauPS4GWZ7+S1d8tZDYPdwb2/IkJRv+doTFjTk1LXt8
wx7HxDBDd0Sck6R9mS/w7HlURknP3fKBoUw2d9uT93QuD6IxTHTjxB2pCRCLsR77cRsQYhe60P2G
TvU+LLyZJnFG1eTSS6a6UUhNX1wb3qZQaTIdoV8XqNIt0+CzhSDdSExjZ3shA1UK9ZYE9+bqF+0z
ey70K9weU+czx6gW/A/QHPYmTE+BG3eSe8p7rB12132R0yb5Uo9QVQK2b7VWqgZe6zX00rd4weF6
IzpeVsbl18XythR1lTAE5YA8+PXDMxzjcuApzD5x+FzJGsKAszSAft693HqkkiHXc5ciXgpdaGhx
qsOM1m/45/jvW4T91TcC6qDNLOsYfjoIO9qPipz7eJn9yhCIpRP/SjiDHbgXaORole7ttFkznOME
+wCOl/tu0LuFaha7IdZRMEuXDstyVT4aCa2ITIGqa0L5l6CRJcSDXHIWuiMOqM+A2dDNdGHqz3wY
+5K/yB37HewztnVJ6rsJr4UMpZGOSdYXV/YSx4YTGk33fAGXT5P2H0rLuchlkqj8aRWTmm+18jUL
3nzO/p/gNwLjSRn23AVnb60Ar+mTDvNi93vMkI7m8ALHBdY7ChzqmAcaef1iDyUvNPfVHnvqH38c
CDw+nogRbInWLAig4Pgrv4E+6/OHiZuBleU2yzitnPmWscBkgg3FVOIlTYSRnb7/PHTWwTnG4RAb
lS6SVIp1u/Vv/rjN0FbmE2TaQIJoGsklnpFnXdb6tU+YazinDwwMjWSS0U3EPhK5bhTCEjPyJraq
pvKZvV1l/xY2KRXdT5ZORCfIcsYmTkNfJVjlydgPkAox3Yz9NZeALvY3cvqWBbK6qVGy17HRAPwI
OIqSa0+f01lJyt0ruQmPfvu84wIYaKu9RZ5yZSr1g9rWN73BGXzzPOvuJVunTK8yM9JcZmj0AfoC
mDQtFITzM0ZJ5FXD4DPOoKBDn8KPtoZxdANY/s8Z2xOSEk5kYrEN40DV6mXqSjqVTFMBy0Jha4FN
3hrTV1jQjJJOhzc4aIhFIZpkF87pFA4DAQd9ZixU6/FnKn8fGrwQZCVI0opJkE68ynyzOO+3CDJV
+FDzCKTq9w2EuyThRXgwRbGsg7YsMa1LDNkGe/D2ZcXmCjxHypjQWGkdz95V5cF+uNvZln9IqmWQ
UE0ObcPbRlLHm6MC9v4KO2w8+Yij5Ho2JXh/0Yv1uRPRrFk9ksbDOlGsloY5TRK7Jdo5dd1B6Lnn
mIu51DMcGyBH2lKoa+G0dmuRdGR61HCpK3r5QbCQrlgeMlvBCG4PLKn4RGgcgQuuWwi0LR1rlWce
9SnA5bpXKUaa0Cl+LzU11gjaicW3kBfTQu5UHj4kvqBPo/u4AO0Lr3StutmPc/8No5C9O7JUdXEf
FkLMy4EFukv9TJup/tVbyPa9JtkCLfWI0CpfMUXPo957//2FBdv6C1BcknNx/rM4HgxocH3gimcO
XXn5dzlLQn9pFoCivpK9eF6adpCNEhX5FFRWd1pQTUYyY0q45FPmJXtECESEOSdiZfXCJ4k+x/H/
8oVc90ZUEnYrQ1g9+0bCfbVK/6NsVctT+SH3vbPtIP3hJIG6pe0WhYTBrw2nFcD+gGLxifH9eYRy
4PL105tCyKLTnBMltvJi+7Yd8IBZvlXsiIC0QguPr1WocISmcpV5NTTLu/bZy/1fES5WOiTa2is0
scxyPROACkmTbkkrFgt2Z5BEK5lwo9jem0VpXBjhrNHnja5ObZlBFLBi5BVzfX/S1Et093Vgnf3i
aZ7Jkj5N4OMMl6g6NPKHKKOA188VrFy/kkCBuNOslP1fd03T1wztTZfgP0zutxYxab3eWNyWxThd
pz8qzI5BxsqiBKknL36XphGdXKEvwYoaZofmzvRRNL4xFRXlO/zB54I+/h+752fW8bDJqUYXnFfU
T+/5Ca4rbwTr2uqQapHVsJTuD/4IyP44XqYKxQXwHvPXEqtQ7kMBUtl72Jg4GTbpzWrKLkJoXZMS
lZHhaHuPy3Qh00Fbx7LOSRuAq2FDspwyw6rfK60HN9zAD0DKiduVKCkVY0vx7JzZIaVHEClModkV
G/M7DEKJYYafUqDQLZ09MYprFbrt/hzbYQerhB6toREWpDsZNW5yVbWih0Ilt/yScPMkRGJBBMcz
JYCvBb66EQU6I5M5OfUD9irLfEIbVmPxZd4beMQOcw4q1oiPCWUmJ69NIaT73yOiDJNra0m1K49K
lNnQn4N0bW3Y2Ah5J1829p0cdkDwQYyGHblfdX6nZ+q5hbYSTM8VKkVx457AG2Id92QykGocwf5V
1Xd2xLNGBrlhMrVizqUhjKha8wg9Z7nvOYtI18OZ91C0NkQJt/TT+gZeZG9kSqpmkuxBPWwqB7QK
Cl2IjL9vbFGJ6EmFMVrzaLNxETntzAd7TRqdZK6alFkMxjnv/kF33TZbdp8H/ozj1Oj9zbh3yGKu
pFKcyPWAZYIg6OE715mT2mhLFnBw1EJPe4n92VTYw6uw65RfrEl9nxt4ERVT6wOt0ZXUh0+tE/OS
OiJ0h0kd8CPI0jUGr+2kMKIyJq/JhMU2lDRxLxk1uYs5YnBVlrmqp0meb6xllCVw/ExnOEc6zQyE
qxQ8dS9qwBpsrZjvOx2HOXgy9+3EL2OgMcMm1nO6WKkO6CMDWKuZIV7+vlAZexQKi5buYfh72sL3
one0ExADtEc+noQq3Y6zhJ6b+5NEu/BLIrw4qLb+NQ6EYvKa5x7/CRBAli/aXc6eglPM2dAgD9ey
bmxUU089aWvDlOPNyDb7IFV1cU4BpCD9LlO3WCmIbEsGpKz3jN6znPg42TjgXH+NqRrQ2uKhj8Pr
MHLu9uAeTabkzWH8Bp7LFngIXkLnHhJzMzOTWwIYKKkB1mhxbrv1n1KI+TzsAOXQuM2my/bR7x86
9sJGO+CXdvHkC6zw6o4xnHB2fbiNUw4cnHKwVybhPTo12U2rFGGzpzLR1zX5z9dVpCbQMNDI8cZF
7siV4YrFr2CxgbByDutKHAeXNfMdbkucguRiUAGHBqsoUCb3AEhqB8M0SFO4oK3KDfIIFMjkejh9
lxKwcD9j+8Vgi6Iqs4H++/D3/GFxbcpB0FXXvbUgm1X3B4/jUtDvSrQd9OO+06VBxlVGwh1BVmsv
8tiIG83xyZdTPKgVYmfGHYsgnzIFPWRyvj6f4nZPbOT/JdeaMtTbMhU+lF8XdUvGh+Wr97X/zzqZ
hBHRvuOdyzW7UbLgwpkd8xEpwuZ3YyJjV9aP4fcp04N0MR6212SoQIUowjN6psXZBe709nMw3wsD
029cw/zCtVepyVFkAX6qrezH6czSq/wjdTm4A5L6yaVHcIHQu0roOYzEsPp/gcKIQfBoSx7deMIS
badQP+YF/U9jZ8Ij1v72Jn1GcSOir7kxNMxBUCWp2mIifGCQQ2oIGIAU4cdWVq6J+h246xclLPxW
62kmz7g12B0qmqn+tb9B0UHNsHl3zw6VJzT2GEeZFBi9B5CZyoFWsBfe+rkTGvsL7R0CpXV7q9vg
NA29M2F47AZ18/jTruG3iZCsa59viK52VXiBNu7a5u6LwYEZ/wMcQUqvCuSu+9C39WR7twIAOK2P
JRsVRpZvriWFVBh2oKxVwPO/yYb2zMEIn1X6Hg9DE/pZeb8VbSs42KgcWLvsB3F4REOPwPnGrwC8
XCe6kU6zMqaqWVaBTZ4lAHkvJTWx1akZNZWhGdq1NCppxRyUgrNsGGSJlMna7vhxRXzYqeJPqZGr
S00MNrpn7vZP/HZCFaDjYbHlfUePXwCan2h3/qe812PTUVMEAV6Qzcu1fC1JmCA7U/cJrckCBGc1
Wjud1crqYo7bYApE6T/DtRmYsYcRT6XHoGAXEU92u6MorNqQQdUMKqpy9ylzvgQBCWKbNHJ5ZnDQ
eje3/gIxkyEnGBaB6OXf2nsf8dwgvDYV+SkKW4XzXQNBkj2iBGbtaa23JHgmlFludrTtFQUn2anj
6BykDkbCuB1xOgzos+lK3S9DIepGo4UgfcmAIQS1jNYD7UbNumraGOqQf5GQ7fnvHk0B+hT/ofRH
QHO/4wHojR8XJ+nYU03ibzBZClD4L1ojjIGzT0ILCdkwmxBDJ8coqEQ1DyZh23R58JyF69YhP012
s44CIqcAgDYx5S7Eid2TB+A4f1lb20zgJwu1rXuRz00lO5eoAdh/XvdPKYJX5w61OQas/O6YeKbL
g5GAYQ8RHyACB6003bWK7teJCigFYpiwyxhCf6VkvGTE5ou5vOs0xiG44YXPfv8zIt34MhgiISLR
zyvS5vAsa+7w4a/r5qpxtIS1cLMUK5yj5YU0iFGpHrRMjGKA0Bm9srkQGoV51j83Rz5sP6kSwzpD
ucVydad1kXyf3TRUPCjEUDBvorxOMWNE2JLvwssYDoY4jJECO+iUnkgMk/N387v9q/+wd52qxLDx
rrVe9XHnkxpS2uvry00dzl2f3kPDB7p+XDMPIyxHBiWtdGJEqfqNKzwLOS3RaQeFulP6o8Vsy/3n
YUYO1ALSRRz4yC3pZ0VGcslihl6va0FMt7KwknqfD0w4Z0wD3xxW6TvVcsjRBFR3HRdR8jusMgt+
3FWc3xaW1UqUsYttNRWoa2d5OTdllWDRvv7IkntjHp5YoQo5p7N4peBlrxWuLV8xER1jjr+6uoiN
6yjwCinallEq8IzNC7UdJ8Y9x7E8vRDFtRk4203gW6VpZnDo+kfPykcDCkl1ov0ikmZmkFqrlXy1
6gbAtDDRVJGRFXc56xlgIJQwNelYtAa+A6pCChJ98KCqJl4yd/w2LxwpdMWk63hB9lQjcR96gUek
jB2hgMTjSHcaUPDSOACgNMkXrvbPvyI+lCeaU1C2XKedoDRvTNrikTMk/yS7W8yYsaSNYjmeVTFY
LzSfQDvRI6RQ8jRSnM+8eCZmf5AMeTIo5jvs1lPysS5V+1veQtfB0PAbvbTYHd8VYoU0qIp9QrMJ
UyXrC6JY59g8NYm3I4/VtbDwyJ1JWdn2O094z2NiHFY8FE4GmGlfBsYroV9Y9Xa005QdGsmj9eYc
1BVxBRJLfsMo/3YT9F237HeVULYx4s1Eqlapv+1+hmq2Jgy29AZRAd7TqwkBlgmns6OYrDFyY5VH
5q9rLioA9mHNblDHcJy672y+Vj3fvX7ZMqa7SqKSEt+MxoyQhttPt8YPZNYdy9nS1qWG76KJWiO9
OIypzkEB+xehWuR0GoZoUZ6eGnmYNS4A4askWwCDffk4CPQYVZf6Cmotg4ZrWDXezVTnfP5n85R5
I1WtiblnZHGmdjR7r6NEUW60zdSVEUU7GEmnYio79jRxVAqPo5GdVzk+BxT9UNqxibaJzs4IMVW3
gwfmGVddOywy9M9O44wg3UOWZDNYnagRreIwf0PCueYTsNnvX0xdPvuR3rgrrINRWxmBT/oj5MIs
wXr60XkGMfc+SPgiyYB/Vl9sMrcUEPjhlbVT6MeJpILvTnsDQkl4RY3RoXTnlxXCQr+A+8MmV99c
z+CofmfBBZGDSj2XvYfwCiA6l23MRCelO0gRNz81dOx0SSWdYGl0QR/WwdcDzMnt0bI8tlmiZuya
CKFDVaCiwJKVJPNNkYKkWSMz0k+Y04snk7m7kxlLpjSVqNN89t507YFBRg6IE+dxA6WCoS1/ESdi
DKZuKjurTtwG0e5brnfI0RDI98y+91EzEJPLkcjEhxc3WdV2DL3ncYSFSLSdhuOBRpnsUNFMkhMD
RdFDpCENOhWZn9IvJCkunnpH2k+yRd7a8yTYbahh/LlodKda9ios5tC6RsBeVdYhBxxH6h6emZtN
yEGM7BqFpRP5+cY1Yez5XFMfB/ajYnIlGtjr9DPFWSYLVMli/qEXMEhonvs/XMSE9xg+ggAU/iKZ
5rnioGmBy3dgrmkWuBlHIBe64mAaQbnP7PFTHXraNFubSYNWlXXN44T0sO/i6K/+C2DSfUaFPxaZ
l2zvuwZ73CJxdKYeAeAB0/vUBWRzRA48h+/WdXt/pcY8/YByw7ijLOMth6tl3HBkp3JmQ8vO5X88
OMYO3V4pJqGnvP6aWe7VrwtmBh6T+8HqT1q9y564DeG7yoa0E9oXK5G7sc4NeOUyy8wpY5dnd6S+
xP5ygRkLH32symbFY/aIMdmDoV+ZpKIiNvi3Wg9jlJT6C6MM3YwTaFpvSeh6ljL0qPYgP7f1a8B4
DgxYzbgA/7oFh0fHq+R7+pprxTROGOJLy5tNZ25hhRd3VvPD67hhgKl061a33Ki4c3QRTwWvn2H+
M/k6ejqQSH/UXv/M2+LTrXsygwYU3Afs1/3rvaFDvU+JtytKuwu/yOPUS14kBwjV5ZM8NVgMK7D9
oJ0USONuH0UvwHYC7j+sGUuCDs39N13qZmvOQNOb2cKiPCndhvu7MF+nvksF6CkeyP4zxaDg1USG
qqc7BxAIrU+pUuokpNcBz004yVpvyYDQSmV/TX7kdBaFjowitZKf5A0mHA+QIA7bU/ZdCBiA1hQA
S7gIwtwG0rPi2zZ6Qj/57ecf9zl8eHRwn9QjTvWLlTcbMbtz/lgDEkq26zcwYzEIQbgpr1/xUh25
DWhyNDBLEXixalJ9ExJMN1iDYi1+GrqApMbqLwVO4LOrRBieDyAJB1qze36VsvUlGAwJtls5prEb
i3aYKiZUlVZaSbY4h/l3dGUGdnejXcY1IkxEUw3VJyE8DgVBNUJwYWXHcdiqNUqEgF+GnBVWLEM3
yg2bqm+n1vadXME13Cln4Opq2bhyJX84t6I3OwdXhRLA1mEfpKlZPHJgDMUW+/CU3FuW9Amv89bg
85uKnzKdrL7JAAKx/7g24QxxkCv35+VwkGvdKwlR1mmZ0eFnIkvOo9sr0QC4Rw1GxA2gsZqzTwws
e9dWpSMHsDeM8RskiemTIQBZ51tjFwQEtNZTjiwN/GGdS4j0UAyp+4C2t1qpIW7gGZkkdItNLBtK
B1EmTzFt0eEFp8hbU/rWN5MAgPOFiXbt+pP2E+t6MAiMDl9DfnooCRruN0Z6g7aCTwielG2K1Dz4
jKbe9njtjJVDImr4T2LwY6YEHehoMQN2nh81Ocrn20ve1AmK1mo25cF4iB1JmF9Wi1P2cPmO3ZNY
t5rbpnOkuQBrtezKbgFEs8/CFga9nYCyqUHQZLtu5feHWaLbnonihzLZbKRqWV//nbd1tHr3PSDz
ddAC89qMDXX3oL7xyJcMvcgs6vUt4HTfzd56/mTI3fPXLMPb1zo7fNaBCc/Lfmh3b74wCDTxgIDQ
Qx0PHyPimC7kzaVMtUdGTbKBu2HqqPSddlupXImbnOLUYwnIbFQ35ArTh1QPOeULvktkOp1J4J1N
bu1XzZ368xYhaFIVWpa1uOJLm6yt6QIjmTEULuFUuPKztnUu6uW1BAkNCf0fxNWg8xhyu0g4to07
dFaZtniaSPjpbSdmISPsYxI33scHphv2K8mUYkLji+oe0l8vkw6lSy4JPxcMaVDWqwaR4B+vQf/3
Az0ItfKFvBu7pJDjDdtAcBSYiuEvL2g8bFxFDr6FtUe3/B/4/WTY2LUIyIKsva+JeF1e29Es1dIB
w8MDfDIEXCacOMhbj+/CmedK2NVKnNy8QJiz2nSq5/VVimWjXEG7vQhaEobvmSjlHSGPCUQdFcT/
hctuUSkJuxz6Muunc453C2dNaOtIwyhyUMoyArjPJf9M9HMCu0fUdIdvvtbAyan5Ia1WxIjqNjYL
tebQsTwO54xCnWRqan7gEVoFD8uQ6uj0RXRH/RkrryxCvSZitbp3s0jY98QV30mqaEaStEUFDRVs
wppQLmlFK/Pz3t+xA9hBvgiC07lddxP60xP4qn1WWinkxzQk6n36yC0meNjTEpERLCyWTNmtB8UQ
htb8qLNeols2tgWFriaBtLZ4lfQtbwVfT4evsirnC6xChhv6M7FqGRlZehIkAoGZJTdHfy8/q/UZ
5nrgTUmGLRSCv1UxKSorKHjgqoJl/UvuhQUDxX1LsDWF/c1BFZywJsxWAjX2z9I6pc7DJVUm8i0V
2rwvTtDcq+3oHQZrJ9wmAjT7qS2hnjXquyp+Sqo4ndz62M4cb0Fd6O7DJGdmezfRa8/BYfUPBpGw
pj0Jb3uwmuAYZR7Uw5FHH0BGNHMpxN2K+rStS/+Ug4blPB11CKNMndPkDXKSJ8o+Ud/hzsTMucEt
02YCnNqAkGjaHtSZl4Iy8W/l+65gGBMutwAGom3XBcvFLC4l01H3UtlCsnzqRWO8T6ngo5YZbh4I
TKk/VfQyYJf2N/nqyW7WCTn7KN+cCn/+B9uLUfHUXYfjUfaBunvyiisusHqegM1T5sqNE/IV2q9f
Z2oaQDGlUOGKZ3AAN9nzOakpjjK7kbdyOUy/zkrW1NMCx8dNTCJs8L0TuEndN7pTiSvpIFLTdTxi
6B8w7uzAnjE+QAogfxz7zt8D7DGqHV6U/WZ2Xndf62WNTFC401K4PUuH7ksGjLLxK3sXzRV2MbZ6
HXySLIUKBAnn0oJnIMJ0bv+eBUwMdhMfMRiWBhciQyYAb3FLOSCGClFE0G7O67508OAqHv2S/Ew+
E1cnkdJCDnAZ+yedmLRwOEbbC+kfGan7Rzhn0o3Szj8GzpXVsuZjQq5nV1l9PrBVVzNEA1jA//jf
JQNBxZXTIKB/jEKjB4U1AgIDk/5ek/UPxxLe37O4Gh841rXOm0dPhOzFCoQqO10OpnTs7nRnywkN
XIHNAldScjM4bHJEy1J6avRGs0TCFWtx011Y84QAHs4oSMwkHADvtwnOs+R+d/NNlv8QLH+qJplV
HC26XISQilnzWJX5C+t+QwRxUr9A61gscoSbjlrjmeHZXu6Drs4cJbU7aJ/Jg46AHqkJP/l3m0WG
ptH2YI7r/vu6WuTlY2XkY4LpKrWyHY9DApSsRRx+UpuW4RiezsxcSAeYDRYmlNqKP50UhT9B0lrV
dHJIcZoJgskLN/dxB0mkKsVLyjYP/YANXY4fuRyFhJ9pdnmJYH2FReDh6w7uLo7v/liEBdwaSF8s
bmhZQt+6BR5/SHFYmHMrT8qfcG+7zXSYUDuz40d5DrefdL1kSMu/IpdxxQP1kSePK+WVh5anmrGr
ZWeKFAOOS+jDbYTa3sBQVaJepBXN3omETHUmcnq6GmBngmF4g5WwUkHPyS3P7cm8M75XH7G1oZXn
nEBkC8rENa1MaLF9HChTP8+4T06J96SvWc1EuCnzLyH+oJLlmkcC+or8RbN9nU4J2ZAtiRVr9gs0
y4cHVrz6zQ0wT+vwQfJ3XtGw1Xv42bAUzhZdX0rt91k6+bViLaEsXEa4Xfky5aztexz5WwsHCIhB
nTP7Wi2ofryekkUXrnqnqHzWLeF2oWxupNfJOkb3b9ITI//3DMYMXCSj6jMkONqqWghP9Bs0hf0v
nXXn3EsoO5/g9vV4re03l5QTzoUEXcEAzCQOpGq8x9OxPyHASjNN/mmdflswIP5VxzcdHf2Vmbim
jPvhI6iMpXdD6v9WwzwM9aIvw/XjXGYPrlmpOG9xk3tKviQ9qIqLQusHhcVBSgqTPGrs9so9ARwO
FNr/ym6sMOgpQI7nkINpU/a+ivfeayoZJ9L6bY9+yjWuf4lkzWP9fhWgPC1hGIOJtNegpoJSa/yu
L/80
`pragma protect end_protected
