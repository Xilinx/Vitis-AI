/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1061408)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAC3VlZPl11OkqdZSnZcSmFre7g4Z0fQ9BKjIML+nNvmPdVmeaLYCM656
jFYCND3ffJu/UWxYLUc1LPls+OHCGWMHMifgLT8gBqQjKSGlJSolUdiiXsPn9Dpniym/LWySF5dk
8ta9J1rf8/37TSv1nnGzIVDnldwdH9sPnag0MW/lFcaiXc7G8UpFoE7hhc3KuS6+MAkd699ERym2
5Z2Iq5MQ+X+Fnyi4qezxzvl4AkXwSAQR5TOjWD2BXo7C9pAFTvCGiUVVoo7HSUuHv/KczKegTrMt
9zGi4lHgriMBEe8Hna1AFdtCYjREAeKKW8IU1x9y19p+pM41WkEaDMxf1TS7tTlqX8mP9w1e2uu6
PEp3R3BIjRKNAqOWJOLskNCMqOzUfGvIvJpYriVUc4VTQU5INBacnzGPBvrYlM/Vq8JHiXEhHoSB
RkZwU+4RFwuEWFEKU7gc9TBKeZWNdFA9dbgJ/G1LuI8YixFPfQZn0EkUS88BmKXckpOCWrq0Bn32
4OchkRmzXoRkjj2TTtv08Bu8L0NV9ssZ1iqoCuQRTXD0L3Th28WYPdvy6zMm1+EvhrtPf5usnWD7
efaYzAACHvdxBNvwX1RUnZHf3zavZ/hevg2CPzf36Fk1420AB6qBbTCuE4+PzO2Dqb+w3TvDnRha
8VfNTCxNgEhUaBPGTiZcDm6DXkIG9xRh6AP2sgIpQSdBl850WYHseNHj8MPgl/4HxIAZfaa/awp4
v42PgbAui7sjhEysdxwYW9iiDsSZDIZSDIE5gb9UVe09T2NChscTA0+5ZI8zOvTIz8HOPumnWt6O
55fQI4K61Mh7lHRNgpZh7w/dCgiBBreUolVhDEW1/jyZEIweLi33DnOlkaR1SwM8DyFqmwpqj47R
WV4G/q/sZ0vnkx15lCGmAesRbWJF/76e6JqEFCi72ohBW4yuL+HxPu1iGpxwAlTgamPV54sOxD4o
ArPsVqAyxKrfzWYlX8WtipVVBi6n9lwi8s9o5dTnAl4idZeVrfwSqTVjaImpc/oigJLzJqWko8Ds
mCywWXY+M1y7cYlAfN85b1eK0BTfyaGefK66oBrqXUHWoT7CYG4Nx022CjRVA+dQd7qhHLFRFiuG
3l5zJLqKmnC2YeB7f0nrgTr1hiITY2PLhX0mW68uG8YC8UFwXEqCYPCuvtxGav4NkOiDpvMPgSgr
p1BDO5sLBW677JgQePbaPnUe2HdF4ncLrFI5/Wzq12v+QiY7uPOJP9oDBKERqEWFy84zAtw1na9l
cHSUcGB8ABdZc/LXQgwT6bWsHyKUPsFd/z9+P9CW8oHhDNq8x1Ws3IqIvJCA44I+O05Q9z4uCgfh
d6l4h9Wiw+iV4czfI84/H7xet9P0KzOw35pREwF+FLffqvH4BEpOqa0eJAe4Ki7fr1IXqIzeNQix
WBEnPZ48LfmRSW+TZ7D5nEQD/ZNTU2BNX1FXPLWZqL5GMxT2uq6BVCC0S15s4tFKxhesOnx7qDU8
zL5OICpNXK/UnXQy1Bl8x6bHlcLsZVk5yMgxU4OTo8D0qarjZk/fivDmUXG/Gwhc/NW92DaC+056
1JLoR2szBGsDy2vWKyTQgrzeqxR0o5KJ6F4OaYKXGQwAbfoocDb3HlJmKAg7NunyjgBg6x5aEhl1
tBStugfO399hJNQ3Ro1lDvCXI65zIUwXPxsSMI0rJ0Ad30tkSXDIriGgodWUeNufW1m1yEoNAS02
JrDiIyzEV/GNqGs4j3vVJVXK2vk/l6xjdygz0PlzRMRopz6sG8we6syNXrEzos/nsJhkAYdfWuCs
bDG+PS4YVmoBLxBtPGRyPavUy+a/fMv2tz1wE0r78yzeenizH66+Zn7VzDueaNdNZfEhH6MkeIs9
lODe+AlmRrzD7braCcLKZXAD+XtBfosMSMx0QFa8LoEiXDbKKQsLjtkGSEDJsg00ZWK/2qfjXQS8
wHzn1EMFDjkuUPYf1hQqTMYMBuAR/z19+/bgqcVqGGIe22wiXoF65SKk1xAdkhIWaDlhOQNrTovk
xplQMk8v7GUifWpVM22EPJnsxRpOk0fNQxTo3iGiSexJKvycfQpEDKkx7rUfMGqjZOP52Ew/PghJ
/dhsyuxSjx+pASFYiYhSXLLwpTS/XpXSJdD5az8dPZLEgxyx0VszHTfGCyJZk8ZCeloE66aAFB23
ApONBYnQ03iDZnBoFwqm6wav/VbiAxAuLjtUij7cE2y4w4MXdhVSphiw+/LoOWOS2SZJdysdkOkM
EB5+AB97Fnc92p/BYMF63iBMULYXGbi9getNOHvZyp9om3YxIw7+zxij2nrLxU2FFMj/eyP9FUaB
PYU06Vfb23g6RzobxDs+ko/t5chTKUTWHBKqCpC97dGTu4fAmI+B1yfBLfmz0FFla3NvK5mZmY6B
Y+z09wyu5YmnCnH0X193Pu03W9W7A9HNwReQIVL9c8vFEbRX0kMLS+97Qhfhb6ayhj0ErbtYXlOJ
YYjvVAfcC+/Tnd33FXH3rJdDMT79HDFmI8DelvoEDKldALWF6yKIJNVAHglH3FnHpSLElAX2B18k
lXXQXEnys9BMqqhr12iIQLe689/2AhzXtA/f5zNoIZvIsBal9wvnobJs5fN3/8P5IwdXAfDfnd/C
iOAmDnu30vIX/6IvGOpgtRehu8kt6NeP7z3Z1upP4CBvRSDdg0N3Nl5pvJSYYqBfA50Ha3Frj4fT
jZ1q9i/HHxCl/hppOAkLAWWkUHvFhu72DO3wfpB9wze5LhyjZxLGrjkzgQ75XziENOaiRAtilqPp
O9nE43qhcEGR2uSCFcoxYxR/C9fOgaGArxmURt7YpJdSziUQvo4EQe3q7s1LdagjquonxDMoA37M
SWmSo3pMS73Lr+kXVmiuAEb8jo9mDSWK/3DB+C2X0rbc6YlVW2l+YxZEWtXMnpK4hJs+B6XeFfPG
QbVnHaZkMo5zGSm1jr1WDJdJiC+3RmGoFHwpq50NQUC57VhYe0NfnOa+GUt1Ymcrjt6hfWjFFdA9
t7aQatDA++Op+Ryj533vqBQmUlE1OPXJFuOXAcs0aQNS/fWlCyIdRpL6S5opQpqJY//E8bAODM+b
yhC677punnMA3uCic0VaK7JalYRordVuLq6scwPnc9ujfkXYCVr7iPyIJGGjTq0LaK03V6IgMD/k
p0vlzPZK3CZqHhzOqllHUk5CJ69cLBchU1iYRt4q/AgFvbeZdISZl/CS3ho+YUIYBW0rGoWWZvmW
jOnoLWceqUDFK8DmyhwVZp2DG9sD9CTAU1SabJJH7EMPU6dc47ZASc1kscPwBUrfIY1DnA9iTbhe
uulsZxg/8H9cLFyvewVvsaSkLBQ4kYohEAL+M60TUXmKuu8UnaUwXxTc0DrCoyuTt8+HmTXQdI6F
NQl4j/4iVYoicoRc89+nrLojHwdnczCXG6DJ4c64DBPJaYFOAHhhcHFmOlL4AjbT3l8spfoYZAS7
+5VU92qwcwoyC3j+2cwJinP010EJldJeiXxEREUbxJ+LwaatlYY6/gdx9prpZZBaCUObBuzzXMpT
ToA7jUYLEuRAmg0POFeXPZh5vW9Zp2ffqRD1x0+mSQtJTIvL3WO1bpSG7AReWsVr2aFE/Rlm96m/
VPK0T2N7eRxSi2q6uXOB7XUX8tyGPUVp1sx/HvDSTOv5blIRQAjW0JJ5/i+D5YzkFq044+cbprD9
bQS7/3BxOc5nZGFS0DEPW4OiIgtuZ1wFQPFl10BgxzEoGAtTRAyZUAi+FR1d7z24KXJ7dT3P4/8b
S61E52LmREetbieWz6P/0TqD7PIlKJKK93XWIU+BXYJpnMm8H4B0i+RpuLLRkrtFaEqjmV3Jc8MW
wsfPAsUyV8bAMvdE+fEcWPFc0OL+USFbhz85MMPahA4bgOMjQ59Bq9bh+JVhSg1tZW1S0hneNxCN
kCyffeOQw15LIowp+AJzPevlqNoDLXANfX1Y+U3zNqKgi5QgAObcKnKnBrOIqg+OxKCTLnljXPiF
raqV4qrppNJf33QMogJ7yE57CoAg65mW7i0JjlD6ZcFgiFmtM19uz9ueekaAfVLvp/Pkc2vOlVGu
Rabm+itQhQ3izytunUBpdaNzJ3Z8AQp2w7qDFEV+iq5qwKnLlT4GgXbvrhKGu3ueYVn5//lJHYvU
CI3BOkKDPq5A9BQjEaxBNDOFTiDDWEmeWAAQhVIns8VAzJNCJh4nOmgT2n1vBn4n0MwuiVfi8GIb
d9pxv/nTh8cuShCQM8sBSJ5tB+IfGVh6a/tXxr+yWbjFCT5YQ9tTBV9kJFaeoY1biVIiWyarH4Yl
uxICq8qaorhn1TOElv0RGFbukYRbIJfTKHhGYNst75/C9WaVgK0EBm756CITR+312qv6EKkLtxCw
+4xS1FXJG23rD4jVqL02Jf7/3anMjwNSJJD7/HmzjXjrdtYsz8YuNiWWARwMcuSnO+Cx74OxYHRm
neymf+iMEYoHrzq+BY9wiofhpKDkzD+GFIKQGjz9gDX+ljqHGQRIs4PUoI8PStACOTKRAuu2djuf
J+L/6R/H74iLVYxr8LEzOZAlJMLGvz7WilIMVLGykQ2pMwbwyDRR2TJ0ucPxJO9tCerVp2LWDL63
aWIoD+4Pi4RB7/TycCgT6PklyY1A/nXguHCVNKx+JMXzgeGMMX31GPZiQ22E7IH1vz69EPUEZ67+
Q+znhQRNPNw8oZUhyX+N5Ct2+3QzdpySMJ4DAdlq0zu0YJ6IooOTT4YHtc5SnwtexhvIIuu/31i9
WpmoCjP+RqisSdihlwLxQ/oEdJiejFcIQYMZcGWXv5DUDE+ZHRF38ITGivMz1+2PuT3Fx/hivAoB
0hFOTUNgbRQdOTX+ZbLtG7arYQcMYvf9dOn+mYbYqVl6Op++x8iPHFGfUy8ThV4bZ1V+vWOMq8rp
Ypx/P2ex0L8H0IVfdZzNPPxEhujgJjJ8rvXZ1JJeq1jhZ7M4NnJ3F7RTSIOpsOH20MJXZD5iGR0y
RSd14FrhUZK8xf2VX/07N+XsplbpJNioSU1NeUr93EIJCyUzBYkVUpyI36aJFTKC1nrPCjFWTuqV
8/4GPEgp4itiQu+ZrFmY2+rMHFxxDcd9ZlHQaiA0lsLUJXY6DjhMVHG464f4OYqccI6vXn4fb7xS
CJq6bfLm5rfaphfVxewdVkAnxZ7wXOJ5/F9PVx54Y9KKVSfp8IWwo7W6bQS+ONzH6Ac5kS/5n7Pu
qkj7jCXwjJp2yyHOPS6Oeqpyn+su71gQf0HiB0PRDxM5UnUfbEHhc1KZuZxoW9He5x9BMtrfN980
3cXS0lf/RVnBopmH7zwPb+MXUsy1UXi9MvCdp81jzawBrpHkA5ZKzzfrgW6Mv1EvzZQ+Cn5UF2fn
w2P5gXJIvlqUOpnHQCGx96Eq4E10b2HgR6HrJePkUMJEyWJpkgxmat2VIjswK6iooqun1je5ijII
ggYyr8kTZT4BwomDGBbFZ5AFc9hgqPJGj3jh1/UCVwDBtBOG4kOSJQ91dYBHOjpSGsYnRO4s+ixv
q4/3KXmHTBYEkfNuRtqgAEv9v8XqPxr7qQ7IjGItDhrNbzRjAQe7lHVGTktBClq5K9sBwb1pILHy
q2tYJgExjtD+uAC8YVnlzi4Ass1qH0ldp3kUZLgd572V8AUf06TRbwjonzRcCIt/nxj1HWd989n2
FEF7QM+9xDFkWMQWxrAM2KpsKTNHywPXvmJ+tZzCLLVmbqsrgymw18rcfdsguFH2r2P2Ea1YMQQ+
1e+H7ZGmNxFDmkEAlKsBS/H0NoI5qApHTf8uVz4LiOTmjWJVcACRaY1xnNtyWnQdUCZU0Vb2kdcC
QvueWNVkIOhAPhDjow6TzjbGpfGUtS5C6BI4Y+BERk/Qg0u1lQh3mRd1kgWRzYcudpQhWRuBF+Em
5ZsX3WweuYdjF7jazybGiaE3fFgzDOS1QkG4VKPglmq2M6jPBeyaChX+/0MdPL1DdSL3HctMVQ8r
W3VPjXKpSc8d4FiL9QWJrxIcO4dhiAUwz+IM6L0zluJmlGc36VhKE8wl0EuwZ9Botam4jce3fvX9
DHCmdwcPoUEUaugCCRhPuBpm1op04zdXBM8vH2PbFhiKpaRG7Skd01Q3Qn+5k/3szEU0AzvrRilC
PYWxzNRarOBab9K95RQbLUqgEObVFc4RXrkO+vWnkjbfG8DkYCSi+2kX/jaHKaL8tAqZdO2BV+m7
dkLGC59OdaBAvwXtqqfE01jWSWZvDd0WXq+ClUs5hLkbY0QqxxQAivmYqjYjUwEXUHHXy5meQW4E
ATNy/Kpxz0/+5QZPDCdUdqPhMHqIgG+wJY0V2WHAiBJK7vZjAZ72V27TtUhCgUTlad/OyPKrhaJP
xr3AGN/IKCBYqJgszfxdEe7mtL9zc+NH0mdvHnT4vQcrHDSi8nT6Pji8owsP/9vj8h0wuDIjtndA
XLb8wNBq+So+u35MVbGVu/a+oBvWpsTobfoPKLXQc3ZwE8xj2l9pSOr5A2mDp6t+mnhKSufk3LRw
QOb0PlddHYM/eaoiGATPbv/zAblgObD6JUftqjD9JYaCwkjcqKPlwPIN6oKsDIzx4562UfnkHN4R
nKPIzz8LEUWI5Rbri8t2Dhajap+hJbLp0stnklZ5DvitbwyW+snoV+ivgFAbcCyIFMWn/HB69BYE
tTOP2X4BvSDf0RviAUxxzfgCHHOL+Rx+m6KBwVnKqajrGVXs2nnJy6wBVYIX1gFMCEHbMzyaNvV0
WxJ7nz1HV3fCB+J6G7miJJnPnzzWuzoR/GqbaUycdZm+cUCycthzvkDbdTScS9XSLZjqyZWrjNAw
p/TugQX2eGxhG5q8jXshXz/a0CTjIhG7Jf6TEbsOrfFi/p5f+5oCPr5W38LHnI2Fv+LDcyiy20Te
Q8qIuwaw3KwCaih6ViGEYPxJb+pChC++R9h4V1g9Po7X9a6x1eOoz+mXKhoEP0vVqYujzcuQ92BG
VWgAyCobcJh7R7hL3aPKcrQKb2KHCznqUc/xba6BTDhEaDW4gLMOdW52g1tIofVTu31Q0gTd8My9
H+iUGWEkJ6+D8j7YQBHwUzHWA/QMxeatuTv4w2N5y4+St89GkmH9Vfo6lOAp+ii0XoFLJm86jKqr
8oEP9stApWbTm/Wq4u7uF9eOyQbeOct2jC2/n1RxgNd2V1DP3pBVfO1J6cm6b/ci8XoLkLXg4cSC
XNQMF/CHAyZDZKQ6LPcN7jI4SEtijKsZyJpXGVar8PUdcTSbyf3A01ZjQrKIcaGeksOjS88l5qj3
XA4jK/+aX1a4FoI7Y35MHdIvS+7luwBbKsZ9Ovl58TBAHs7hzP8jJSkqyotXHULPC/WKzwXSm25w
g96HYTdOOEQQd0rsKo3iolTEEgi19EvrCKIpCypVlGndAYmWflss3BkJXFxao0PlN41+SwDaDajW
Y8feAF+tCPri7KZXD9MZToZljnsSSXkZw5fXLbkriOb5gYqKwD+kf53VIpoQuf7grLX+jnYJDP0x
ThxfNA91mPlec5oweyOvbkhubVSWKDDsTotrXO8mCCv07Cee2/Ig5YtaYKZG9FNu7qzmZyvZydBS
7grbND1A2dBFB8qA9ZAYHAB6+K8AiDXlMT/AAeS7qpB4bZNoHWVu9qsM31MWEJsud0n8RtIjC2qa
XV2g7S2mzRVteoM/8V2iKBadSCeP0b/z/dP6GE2QZ8909cVmFEN9P9n4aaFBUpCA68JaSloiMc+h
16TMFBT5AnKCtl4Ru/gByfB5ek3XhFjmyI621Mkr3lGA1J2eo/drNz/c1hWAHTaMrYiZiMPXmAr/
fnNSPKECy/Ahb9spW4xF04jJsAi72rWPPAMvzy8KmKpJ851UqU6iZ/Uvu1iNaRUlukmOi1sWe/8Y
rY6ScESCKP4BWnfo5kfqKAQb13piaIRP1GKoavuYS1c+LNYAm1dy8bYPcCi/OsxBo3lAn/Oj5qcI
qQrmVHhgzdcuzHflbSNN/pg+3ZMPD5tJsHald9UJTVyw4CzKFV+MaZahb481qJT67kReu6lYUdhK
Yni7kKoa7pUPMTriih94gAQSL/DfWS5rM8WAXchpTGKKa9PASk5umP1qcKdvxzjyTtDsKX2rCGTh
6sRseQTU8/pNerc30i6XfJ0KUJZkd1E3Epb1sEcCeleRWZE1xM91z+LaPckwcFfQfdI5pnho8A3P
ILaHKB+QaZSpYXNEYlkf9hMwr1BevKrR6OH9Owior/jiAkse5u+9+irYb9tsdMth1QtvWoXZnSx3
+FVy0Q0hoBb6yjyzVKBTJAcsr/t9kKs3zCRRUP7d0+5w/Bz9IRvJqR1OZMGhCh/IIciqNv5F3AFj
zScbN8GAgGujeg1Bs2M2JLbk2a1r/jcZfyDhRbhJzGGIo8GltnYnBkgX0kUz11V8obitz7QLoA/8
OOmb/hPujPQF8eJfjmxEZaqT7KorRZ4to/Z3j4eeM0zMxqAt3b4tYt/Peqi8Fd83lblLhTp+xtLA
9ZF2wWhUvpgNcFDqwuS23XeAQkISfSlOXrVKgRU9EZjPXgZE5W252lwk9mm0prOtB5EAacyhptiP
h6KmNElwADg1RCv25Ar9HEsIsRbpKl7nqXk1XrNnQhtBK3AcsbM3CTQLcuxTefEXTQQJOVWGcKEG
1MGwM3eyQ7soq9IFiBuRo5Mc6Pfap7DA+uPOneFJ3NHhTzwfZNhQ8AweqMaX4qnv6ZaWsM9aHvfx
9AYFWU8UF9YcBIChbH4h0/zUlXHy7wG/10K3C5+YFEJeXoQStRAhikTl2Po1TWohyOS0l5sgcRly
aDKCpqHMo5M6JTQK/kWf2jEBUabpa/9+sIcLigH3JbWgqKABpeWzz+YBVbyFZMeDAL7U5y57eg8g
GBrANU1gqvk0NLsKvVBjgqHExO9q32sDLAlvtyBGwEM2HOSsbWdjBvY5lyqPX2LapUJM352+8qYU
1xaOz5uGaq9OKQ9eBMHYGGtCqaeRunY35fBEBo74VVtNVPkyhpnJAUH6o4RUzuix1O1mBksklIQ8
ZANNAw/f3DXuujP6tsPWCyq8mZx1AUwudAOACqM7yi8D9vtfHlBIoLp9c3uNauMf0sKdG/ffHFav
OIjX9Qr2IR88w+GjChNaDl+nta0zHvHs7p1jiUOb+T/zU0nhrJvQ/pfIbOloQgHbP3+nLrR25IPr
xn6R4G7sKm2exxtSpANDhCtPcLNAXFm+SlVzdodLNhPtPH3hDga0MtswjHWLHigbG0Y56uSIxo9W
ydOU5apS37jjwnI+mIP1r0qc7rhSKBRb0r9ZD25Osj8asU77AG8M0yhAtPkXpHSVR/buoHxIuyJP
Zf8v5uDWzh+zmK0zeQujIlj6pU8zFVBT5xmQzyJZwd+f7dOqvMJf1codyc/Nn2k+d+4iybVavsBY
ZpUGCn1dOdOGUDs2Xt5yfm4w0bFM6q3O9gW9tpNrzx/f0xcNqcvdFHZ1Q1hBcTNVNCz971BpEdh+
IAnS4AhTW1QI5O4/O9zhaa8JvhzRIqMFrJbfIYiVdk0llbRu7mbhakWTbYN9n4NCYWAwBg0GRnux
HBMZsmkqgBZVeaUllWDMtHdpqg1PdJ4ALq9fZ9VbnUPUorZ0uoQKxbPfyWnHeGksCbmKGrQ78ULP
Jz+J9/dJq7ZvN1+0ylVTvQ67rognlnpap7+eNpGFMpjCVjcy3Ccqt1Tc5sN3aYf2dbg/bUJm3Zks
czxO8PtWAP6Yp1kUozq6dq3vzGhwoLyYYUqdfsC803UehM0NCZQxas5wFFMsJ8BEU3rQaa5Fv8lf
n+vvDvFwlhQpTwHvfrRNH/3NlPsQhem91tAJlNfyAPNyMUskRC/M1WHZ8aXqSbVTyWNAXtb7FzIl
RiThF8B6aBzMuyd6gov0JhXFhq8u/c7pZ7bMIbFo02pznDe6t13twSIKq/wfw2n50BDQh9EtbUuP
kOcEV8nlHH8xTtY0UYZYxg66BoBVQt5WcCx8AHeGI/WOgx5nG8wNZl4oOkpq/DX/PZdIGbpVKXqP
FK+Qtw323dWOjWcL2gl2gceupP64U3A34ER28sd9rR8/D/G3SUltcWQ9DeIPbtIS2No/lJ2BtfyU
L0OgaiLQ7CPna3OkEm9+esXABr0MoOpYelOouZCrBzwrP+FHXlvtmG7Rcrgb8/oVNJhhjpn7e+m4
rFoqhlGNjYzLU9TSPPfM/gO1+veGHXsJuSRTq63hqLjDKb4BUXNin7xpVhS2vNhVN8PDdtC1qAf5
YmwuPb/1qWLShgRNPt25m4I2RSj2niYpA9T/1oa3SNE+rJXTxiMrnDXLwNe5eHaZoJpS2YynH29M
9t5uFFEYPa1wsak187MQ7r3p/Ri1jLositvr41sv0/qhmamr+Gj3ce7wsiaPbZD1IrV6wKDYbIgK
JduZP4NAAdPtOs/JaxaxoS8G/c1BXH00YeQtJ1Oj0CzceuvM0HXmYVlsyoDLGpwEn90w2pBFvXXG
+aguHLfHD71RI/xNA4XrmyL550P3LXHYEWgc/bInAQvY1Wzp3rEgMaJ+ZSqc1+XNUiyZgKfT+vbo
ktPDKgkf1zbscrwavDe/JVNfi/cU6Tagx9V7jM/05nqkWD11fUv2kUQ4kwrEj+tzyaJA1fFSl/TP
sUWP9Dl8y4hupWIKKagQRuamU4T054Nsvih12bg4Lv+551mFLmUEnH0rDeiQpfY+VA8shHOSid9P
9N2xKPfVq+lQ37rYCJIQNAX5oZodsnJNCm+7ny2r9IsdMJTr8ZbN/nSf/gFRKs59k8XI+mrvc/ym
oFx//HEfqKbjCVSqGDkF6yDVhVTWmMElaJtEX2R8mJe+PK2VKcfXPSgzolcKR3q4zhJk87spHbU7
FtxwdhSlfzYUPXkqluCoRifJfa0xBWqoR82CGGvPDIGvxCjqpb+foTBkUagUS/NZIpf15uZLXl6E
QW5LS+/Yc+dP8lJG3NTOPspMw+aR6XVbBWzmOuUmoupH1UPjMtDyOj3990Zo75AVOcgJjvbCRlYP
a6ZlEeLXWNXCmWVaAvxPGk7MbADupAkg0h8i2EeADg6EFRID9bytIb9378jDlhNtIjYG0BYjBthK
EyEqEMJftxP+1nqysMwPGAPEADhbRfjiVF4SKbub6x6jbs5aOSxqVXkoaD9BKo03xrZCPjUBrVpy
H/K86etZMYyTq6unIt6mK9TiNurtxACum54Fun2NX82Qut2CfwHYra7W58Zd2zAfMFcxyiFJeaXE
CeIpvxnIFYwZf5R90mS//3127KB50HFWcjpzQoSLWowD6z2hV99SWQmWQsFI1zDSWoq+baNjZ8mo
zBdn2BXeCj6wjLH9faG+BrrAQ+KSESIQ8Lr7vChAXfGCnNYadI9PaLKRfPZdJ1h0Uazcp+dpoLsL
UMaghQ0qPJhXl+/Rl0v2+pdsUNXkNcN+9lqd665PqgcjfnypHGU3LkH8jw34fm665+GdXOjjJtT3
sKL2wpAUSKeQdZlLpkKXpZlI7M3EM8/uJoPhhnsFvqiFJieQjfjDGATTv+45ck8pO8Kh8J10Ljl/
0CP7TTMShcz5WPUKdCaRSIPjc4zRFaxx4GGTaBa20CHpmZmHYvoRY9ivSH1QzTBxS9TYhUzc3DeV
de1GP+PM01qt5kzbeJWFdqI5+ooTMnKjHuTcBSaPIii1lo7T2Qv2H1f+hftJXv+4QqVSnTUNCC+u
4rkv6f2IllX4jkjAeT3VVxWNEoxibr5e9CTrasEF3r/xqTSV88NSGQNP4Ri2LcJ0isCzxHr2ZzhO
d5DzZZfcGYfqo3jNz7S4RMw1qk2jtb8g3KiyDyvKgmCXdS6bUxYJv0tfYmGeExtCEPcJw4uJvgXi
M/4tmaQ+Y/0dn+YNi57Vp3M7mpaMEs2tlG7Et+J2F5JXDoD8Oxj0Fec928gau99Q3YRhLsGHkyO2
1rK5cb52U04RCjkCIf9yVundtmaHWgHU+FkTqN6lBmWbFd0mBcTQziZ8flpCc8W15Fx7uqswbHSd
Bz8mKoC+BdmK613CVf/28o6n7K1/uYSemccCbSvtj6R9Jz1Wq7Vlm5bHpIPf1y9fWEwXbJ/I1owU
0v6rATsNEYI4BqPF/iMcbsB+xQXVIu2CioQVziEMmshq+l7qUaqaXjYNixAh9WaOEvOjk134vOqR
jckTXdpdZATn6yqxIb0AQz71CLX96WaLl5RBagmMFsoK1RbBl4RMFGlPvCvE+LXbehVGW95oGntQ
IhH+75+2gIS8NsAQmhR2R/U/GN2+8AbhN9bV0NedEh8SQzzx4ayE0lPvUT0a75D6wrXMrmUKIyU/
oOtNiNds5daedi/lf5RrTcDQ7Qb/3oCAT0Dgz9GWzT1iyTbIOtKifpw6WoFz5C1frzf4OxX2MTDa
mKcsTQjmGGx+fF6WX5/ZWEKp1TXGe9WgrGq6TugHaIjNK3oWeoM1IFQTWQVgUDXKfKFJNTFXZWUi
iuxlfYA8OsadlQ6VxuJ2cGh/iIxUsH4rAHpZDCWXI5lXvOC7TTfPvVjMhJ4bKx5hQ1Z0E/VEipVI
Xe7y00Pvn3Dr79FQeAhh9176x5CTIVlLPst9zySPtmSls0ZPZJ/57hp2M1b77UBuGLtgGgu5XUdW
wwfCArM7LT17Y0xAZiufSUdXYlUcZHwlat4bOmz8nBpw7zQK4DyeOi2+Xhl9I5k2a8uVXG/1VRTF
6kOEO58K+re3AWNL0gxhUXZxCAfg+q4boZxqF+2cxnEtqMPmOMXbflNUC4sJEWPFKn2Bg2GfwhRO
xySq1/SdG0k6BTErz7POG5qBIcLI/aXlBX9oiMAeRw/N1+3v5Thbn4iLR+Oh0qpgCiO2+cGbp/qO
zQD0hdVp/mKD8bpNC6Cx1dXJkVql6Skf4hrpfYyxS0DjsUrBTy431BENH3S1GLeDM7GJ7vSCZjrZ
S5CkRhScFTpj7R5nEyP3zj9GrnY32skt0jeBfPEc2rN9ia7/WCV76ORWTJUg0QkyyQwduudG9g5y
0V8PmqY3whay3zjSc6JzAGil12hLuQ5/IuavFp+0UuIuaqe6RCJlF7thXlCvqQQdiWX+9Q4e2k04
8K3rS2pwh8yOPH/dWXOgZy5dPk3Rx6dEaUwTc8u6bvCgXk+wFwq5d4eZKijsFSWuzMu5wdDq7N4G
xP09oK5rTCvE2SVVScx5zJFo734lmu/Nx26IaPOTl2NaJqCS9andyOmtDsBJx0TC147HcI+dTJlX
JKc4Uin4I0xMAmgtZcOHdQBsOtCQVqQZMhLxIRL+5n/DkoSRHXxPKSZ5D5XMcabxgVHC7H3dynbL
0opQa3WyKaMPFX+ivPm008hsm8qaZnSeNw59mwk/3tj5u0EePtjdz5T2qW4Sq4UStGMxyVBcJ6l9
i4I8SDh/9+K3x1Oa65yKQ7IAFViwrI8/blNNqh1bgR+Ch6oEZd1DNXP71cJYEp5MmPJjwDeYOO6e
D5Z6ySo1Vab1+8qzNRgOVkwLrTNUM0NCgv2FnbQR+7j+KzB+64b7PAFBnldLxK9tSxmELzE7JwvM
vfO5jXQD5MZRzluE47ShwOuQihTPctVrf0IkRjBKi+DTTHISvzFuWfVTMLGCmjbsk6+uCXXcHk9J
3/FNxBrjSgDHefKEPCGdFaDhueoPUgE4hOY30I8oNMOETvcFttsKJY0Y+VgoP0Y1cKkKN1MY6rZK
UlTFz8jFmpMiF78/YN+CxFO/Lm3oCzrVmD4Q0vIfAK+kr+C0po4dgI4N11k/T/PBWVxSDokCiKtO
QMHWYULfP7zhc1/F2CzNssKAbPizXuk1546PtV7h4bJLRJ3ZkFL5yZV5QRqf+jVHF0wl8MEY+Oa5
Ll/B7mvBhmDi++Jt5SkKnKECg9AZUkl7Du8bjDz5WO0Vux/aRKqv+JZqLdY2WZaRn/DSl7S4CD7o
FGmSvfEg6yR16i257dkDlcI4tB+1P1USKFXh0DO6R8Zy1vJUDH/2elwN8kra3jLnKpwL6GpYxIu5
dlwSeQx0AbMhQY/C8fkTS39A22UsYkg/MRQc84Gt5+idlwe6stsziTJ1xAMXoSSs9Rqwfs/V4JLs
5T3uEDIeeEsvjh7CAVVRgGxmNGBK1+gVT8RlT2aeAXiyhwdpdWeSF5DbXYNyAYtAx2XtBGrXz9u/
URy7WsIvH/r4li+4jczkDWplbxX7xjsK8naVXvoMaoxFN/HAab8I0e0AfzZRf+hENFAhpRGUtJVK
obBwD1yOW3hjCLHUqg3eBLX/QYWQsRx2QBfxvKesDc4HfhKOXalWC9baS54w+jaPhTpJQG9Ng6sa
71Lq590nse5QpfG3lkUVVk8ylSNuOz15tt/WDlI3AI4iuCx1FXRPUP6MkARJRs4m+bYk2iikQ9EW
5etUXpmzr0lLXkWFD57dHHHOWxDkOnGh60s5AQl8nnp+ydKz/7PvZPQS4rivtdw74DHoDDS8G0OV
pWHWVLVZFgNAz6bjQjQXJ5s/HgMSp3LisI9NpG09Ho7zzfaPgs5XEyla8trUqcJnew+pJ7ziqS+d
5kdsYBhlHd2TyOI+SrYCsp0UJFdOHWoZFJFAb476t5t4LRUlg74u/O6Xq3tY91pK+EvorA/hCJEe
h1dAEuwpML1WA05lztdsWE5gkcMdaXNFuupbg0X56qdU+6+eIdoZvzF4aF4lJytXV076zjPfvifz
0UMF05S9OZrid+ZZiDQsiV5TK7+nJuPQMDrxCb5uHOJnoPp+LX/4MJDKUNNDWQ4kukUHHHqv3h9N
vm6xTKbAQCdFXKUGRrCCeH8okqzo3H4SkxBJ5c+WeLTlb9WKWwiNnNPQ4+P9RupkLQnq6BqKTszS
j3x0ryIfCc6hIkkqvnBFk0kIo8rKZvmH2d2p3gSo2R2GeMeijDozgZup0lPMT5PW75Zvsw6xqNtz
17M1KkB//xx9F7b1ny+6Jj3G7qTAVeUcbqKh3XrtKzw/doo0aUf+ROIYg1WGuA+8zCyE1FXwCiIw
gZTG7ZbGNP5TjOkmaC7VLhGUf8dZJVBW5345p4qAt9e3m16xntAnZmRRjgAh8ZpbOePI4Cvy0oUd
OM2N7sguFg3Y1h2yMixLDUbslUKuct1fvyczP2nmY9OeQlgHPVLGt+ICKKdFikKJXetk7K/WPNpQ
WYvhfLWNGqR1aDLjQp2Ho8mIiPNp10WOnp1bIWI1er0P61vpVOjDGlT19KfmI5BjYHwmcZ6//rHh
umefmkLLnnlMKYRiOTSADE0YMhHQZMs10lq6opd4PLOAXuKB3/CS2kryumaKBwF51/aBml3nWBd3
Vc7g/zxZa3cpYrVtZgKHD+MYhQaUCgxC9B4N922dA1EgFT0EAREsCAet9LpajQ8yiDOga/43uDJj
mZNNBPKXSg6zGojCUwGTBUyPT07fwCkIA4AQAfBjtlCWg5Ogq4di3PUKcjdZIDAzdtTZi/krDPgd
ZIiPLw0NW4oKc1DJmY89dqTaG5CqBOixu6KQVCs6phpRX8oCJL4YVEUTTjTNyxOGJpnWEfLq9VRS
vqOEJ48FWW0ojWKRGjZR3MnfDf076ylgnwToijsEM9ATqUxhb4IbZ51bagfBTVWFT/QqC7WckmmB
Xt8qHCS8mR8XI1Om0SR3JDgwT5Y64UB/e3rpyz4ctyXzbooaYqnxqv/yrf02QsM/tJA1d9vBGhbr
FBk3Q6XtwpPNV62lmQN1J9QnWmwmwdnj0/6U61NR5IzIO8RnU8K4eYC7yZpB7RmSYWKqCLlDxEsV
eTXxMjBGdx/QRZ6KA/mZAwFV7OnIeMkl68SguU6tNEhM7t4eQImHWXdtcTTep5uyXtdOcURXqPKV
ME7d6tLqHoQe4yxywVhRE/z352Kbg+hMfjT2Z823/x3lSEyZn79S1mi+n4zXp2JxZUklu1heiJlx
/GakHSVaSzbRuozGdRU8kAmZ/T5jdGRBSh5t1EAB5DFk9Yrx4cqrVRa3oX5cQ7aJ5xtl058vZr64
p6neaATHVa5aHGUTfebQiZlGYzNU4lIEOXtcgPFBOTYh6mTd2rQV6xqnC2BpsgQfHqnduaVWFDFW
wU+La0ndhDTyEn9is1Qe4DUf8FdFVqmJMLyepNR009xUQUCvAvf/82yprsoVdfhiTIfElPamN8yR
3ahk9pBhZj7nN7Jceg/AQyClGAgIjKEBaQ0WgdLM6+EIKGDA5d4fWRec3Qy4NmJxIZ+Wd6dnVbiz
UTLglY59AKn/An2pxrt0/NlDqusq8m7vHuPhH0RPtwBXXFoPokHrltIBH3qXWDdiQRhQnGSCkyq3
lx7nYEeThXGM0ZUqUVkNuZg0zwNCID1Sf45RigNLJnyE8WWqNHC3+BLGE9psdrtTit1bt7FJI2JO
V/SKRmuq6S2SqA/BJNj8xB9S1fsix8V5dV7R9hDi4veRa2BpEYgvWCI5M+UlSm8IxhbFzDNiMuG5
khD+Y5oyocBHFyoTZcmiIG78E+cvqVUd+++K67jHIZ6XzPTNlfT6DP8jFhZTcN76GdnWMNhh9v1U
CKiPrNPR6iWjRs9dCScH1vXRXeDO2OvADRiwH1Av4/43ZM7CVMkCjM3EK9rMShcXxDZxWpoFiHeh
RCcSLfwknhfjaV09jl3uKlKaVfSBTts6LEje4bzGv70+b9J0rhCI0XO6SOHOkUWosYVw4NmE/MO1
TxdlAnVgDoxmEQHYDH3JN6YcsPYxTBfdbVHwLQMsPcKNMpKivk7tSavCMWmfvSk/DC6R35b/qgpr
9AytvauG9Hsv5FT2UL4PMLIPgaGAO1GEAZkwTd/eInGROwIn/8zoeKrvtrSXMctd/m++OoSHJKG1
rqWhZA5/GMXazr+qAKSpQooqxxARaPIqSZXbVQBaR15TACFUfh5AsdZ8qlZiZRBnZrJsdjQgLVil
7vgo+WYCF6nv9/woDQxjvP4pHTU9UMy/KMyl4jARNd4LP65OZ0ZTkNbGnFEfpWF5z2ABfAHUEsFM
3p87ec4dVkZQXZ/FAMVbiCj/4ig01x6ytnfXFI08YvM0MXV5h3/0s8wAcG2iLx6r+MOjlxDyXja5
b/AknYWHHwXxS3+U+Y5a6SfR31ZR4U4REABcoRd4zlNn9JQLJREIkN4QuCWC73NCunWawqoN6uWE
jQ+O+QXT18Ufb0Q7lBK7zvEMjiCg5JgB2zokeytGMDLHo/Y+m0GlKe3WHYBWDu7G6CMsJ+BQ9K95
23ZS4ukCAm4WyL+ZkX0tGjMvmejN/u23mz46ea0FGODb9S/z6ihX2Am75hix3EzFTpOWPutPnjGP
vqC7VNEcsvJnO0Z+Pg2u2PQk7/ITRsx7VIEQdzxmhp8y5a7mRtA3CDUB1potnlSrSvWzlGY1jl6K
z/FLKmGdmmBA+KM4HIsmXJ4kRZ/Cr/VBYKCCQO4d6NB2rAulYmLM+OW+XA64cEL2A7YLZXo0c8yB
dv31y0H3H6nKki8jxOoN0bOwgLnHU+u+emvpHqHkkTigiPbTwGkQoyIJKfIFK0wSm2vzMMU/Aemb
cZBRZ9aD82UELroMCMbgFgUeyoqUP6Y7ysA0VGIHg2YCb4ij56tMK6Cj3H1hg+clVUfctbkMt2q9
vLZEPShABIHkZFmkmqKREOOGmhqdcGUzxiSF/s7pnUoJdw03yY+OBKFfrHy7ue9r3dGh1kNf7+MZ
TObHQ2VZRaD5GG1XTXSsRdHHW/eXwSvzFub/riyJELEpmvcrnA1QHWotCdVAdKfyLKn5pMfv29f7
409AKHqNBuQIpVcsdFE0derzF5zS6/o6u784btb9Kjt33wG3bjF0cuu8tzFZJ3zmpMECCgcHMb8h
OxBYcscX+ubQxoYsfKXQZ0Q9qE+Ui2C8uU6bg6pO4sjlPsmVtniWE5Ee/X5sdu49w8zclxP/b2mL
aM2uUEVo3Bqcc5+iUzXBRRBHA808yC+fHjZK6P8POAdYcb55/al8x7Elnlr0mZ30NPksOzi56yUw
qB/JuEeSBPquqtPekAkNdWyyZibo/4wFJJatNzi0xjDt8RIJ79lAgemrlFsp4qQPEqGZXIdaHhah
89hb7hv2GNaEubb/VNeYQAymCznON1KI5rgOowNzxnRDqV0B77YKQwpMxZj00rZR9juuflV5WQAZ
IG2wFGJq2W+4+odQyTJl/jQzISht7ZngJ8dgj1Cm1hmNYwO4fbeoSiMluQHJ7j1bGAqhhOv5wtxp
q+wIFmOKktdlKNfy9JqlY5myqynHEXNlyoUhQDcTA2upPqzDjqgxolaRqmfj039YxZWEFfhAkYsp
muCnEIvVu90pt3fT4V3jTHiK+XwmYB9br0ponvZbGOLIFSngMGS2ZH+uqlwrA3M308QN2TAJj3OQ
E1kTGt3HB6iksM0cfWInlNt8l6RbgITtVRmItJ8vbtIsIJSj3eKnoTtHxJ+ZrE9maW9Ozl+HiVrX
/Xr85tujsb48JJ5a74AplX7L2SuqRlQqlB5dqwQeNIaDg3O6rfUaYDgMzNZ68V9qsJ2V4xvIzLYd
eNcBiL2T4gre9MkcD6Qci20UwKCuT+sRttitdRlcz4soU0SfL5GflUJNZPPpq+kG5Zi6X7+MQijL
10dvg+lymCYQTlhfY8CfnW0RMgUbk0nLQiwk/RUYxHbyDXGcn3Zj3fpE6qHU8l0qTOPBdIgCQ05y
U+f4fcyTv/frDmY7Xm8G89kCdBRkgHQHWyOCCydoIj9IIz+mywk9EZ19/sG+2Sd3q8A+7m5ltwhW
qjjCxogwXq1Drg5XQ9W0AR4Nm16RicOprebGdPo3tFAa35DhLmBExU6/rNR1MCn1rwXoXKc/i8WP
xQXVh3Xo/rfoazgDpP2O+Abrbr6W6ZFqL8U8tcM6/NETtG5b59julccjdNUgMtr2Q4/Cgzv4pttv
jaRzWibboTmFpxz4QwtvkkMqjwFtQAEkTr5ws73D3dl/ucT/eQk0BkSmZikaS4hSI44r5xaFA52S
4zWxlY6KkJK4xuybVR1hqgeBdrcDSIo/CRuQuVGrTkSjz1KhgxHoR6YP/FQxISnHUZZgK7nuyUYv
cJJeX/WRKsBIm38kVu8m4P0jyG1oN0hmmDuKZpoSWbIPglMQv/0vK723USIDTMT4bcv713k9JkuP
WbQsPa8VciiZsTj2MbwZ/u9ThY7p9gAEqAYZeACTjaixhJNWBok9H576vWaUBuISWzXmLdcs+cDS
00ihiVBTkqT1K+k2FGWyQ7q7dlTxfo3gtP3TSdQcvGs64vxXQdanOM3U3qRq3byvYIFr2nk27na0
WjwcUeQkf7MOnc8i0GBZYpToabW+6AvmEqMeehdL7ZVlahPGNA730r0mK9tBiUJeRAe43VKQwD8y
yu7scTFzXC8uIxpkcfD5wcmHzrZMC39zE+4QeidKo1s1YhLPyeZMQbcxsAI/nM0bHPgtIyjieYO4
KxEwC+UTPuVtyaBDKgVv5HSOj/cKqiG52yclxr0Sl0JuVzSTJixPNpVExlhcnkc4VQ5XczaMnG16
HZXT14t5AnjvRVyhTKXxuBf1XM1Z+T3/uK6NR7UIjUfiOE9387pgTWdK2QPIV+PgJJPjZRcD8OCs
cPPl8dB8+InZaOzNbo4mmtruiiriKyBF3zBqjPE+QD4r4kAmllWSfzvDOJK67YV2dT0DiLJG4IHq
0gJmTUEwYANNKcZCgcfIAY5DvvZCaQTE1QOxR0os/gc1OYN5YMJRJ0eqhl8Dra3CqLWqWCTHsfsB
seKrU0bsDSAfju0OQJpifA0hMbzpZtKJIoBXDdVHnYwzCu3FCpnNPcBwxHG5U2aX7yK9BgMTmjEH
2xn8Rc4NoAeAzhoaO5BVmtU5cqsprkDB/EXUoqie/2WsntseYOw0maUb+WsOe0ovJjhn7HicPBNq
PsSvSnRFWt+YzrDj/RUJTRHOQYktogqIwPAk3TzcK10ED8sEOGm+8X/puVDUyWl9jM7UhdVlhN5D
SQtaV6KR6OSA7OqJ+sdPJuUfBcoDJZJFXYdg3NK+4jSDXaLgQkiKRkIYlDUf6pckp3Cv+ZlEYyG2
4PRQmSOlok79BvtbfXc+0b1trSmIkjXo5WR069plz945est3kX1YpZ8noRR4D6SgCKC6Sy8na6/E
YZRnguUjxnHlNYvCgWkT+sI96tNURfUE1QmhMKEeK5dnC8I6aJQHOQyCvW4BosDLMn3WXM1s0ivQ
dK3U9of01pTgQ+RQ3RozZzybqT6glAxeBMmE6N8rhJH2auwjnoaG4qh3Vz/tM9Vtwu30e1YtmGTs
NdMYUUW0midk5u/vHeccgMnVklMUl+Pv/yP8qVHj87KdlN/jCpzXgsxOwhnO6KjJ9V+aFVUxQ9vD
FCB6i4SQJWk7zbhniVq32YofQUl+wSxTJTdh+O6THqCys2C+agZjeokPJi9exJFxHrkS2AzVGYaK
TaZN8R9Yr82+oeKPJBZDstFk3UvE5xB4eHpQBd/aWa3CSq035uvxJpaZ9lUVms14oDcm9k87WzP1
KZS3g/cXMFENvFrhMZYaM6jB6n0v6UVHEnGXNCI5u/2UEKelPHVNJKqtKNtgQV8gjB4YiN4Qx7YV
HoCgxNRrNtU+PU4qCYrWek4bILrJpHzf23J/8cMAUrBcpDRiwUiiwMbykMX4xeFgCu1EWV9Z9VEo
65As4lxlPPkndrRDHmCFneOtW8jX1ViRIw3Aciy6EA/QWyt7kkkYpRPKNrku5FDt9Et4i+nF873g
WVcBsf/GEtJr1If9a4YnfvJ+JeqESigzy5St6uWjeuVpsvTqr/+U8nF3oEXfHs6YlFzd+Ozh4OiI
CO3IiORZ74m2QT5IUgFrab5paFTOzcFEjf59ff0dHMVe1XFt4eRj9URzkzr9pQ1DgGp++iAP6Ft3
cMfYr/+/boJPAweCzf2Ps0M4IQb93x0rmnV31C9ES918d2ks6y0H09dJ0MhfuWI/ltXrZz9nH0Fo
uM3ubsLQ9jYCnCqmc0/X5mlJXWwS+sCfmf43BTzqjZojdLvI2g5bkVr8kkjDqCUS+LpY1xU98g1o
MTB+MsBtNCop8LnIMVq6857vhAGhZxVj0Dq5BK0Y7aOcGrBG/ln+75QwyX/SJtuHCWKEHaYqi1z3
9aR9dtk+wtTH4LlY7y/8MSBPnsCl7eY86Cb7k1sLtc0zZ2gu4yQbFWpwWmIRxfeurXTm3v9376Oz
fYYYz+g1EFj5Fhj6IRyupDkxeIYlXiNM8wiHkE3BRVzvqtN4nXXjTMyHH9v1vPPjgF+vXtCzsCPm
6hsOptrKmMGsdr+2HvB86jo/Wy0CbKEmlWPKLK2Oc3VtUvDrZQAzB0yXxR2Sj6zqvj0p7WEQ0F6M
hPT/qrm+eSfgwnGx99tAj9XvcauJ5RyxFd5i1qXFaWCH6c2fsy8GKgAkBVDiu7WiMqhuzgbTGL8K
bWY+Oj+sv6cJF2K+8SLlcfmqr4sDmM7/sXV1RV7OJuK8/aYvekEPRG07wUW7k+0EJekJ5vldCntl
uDxcC3aqsf8jKaAtTCPYfV6PtzfIbuMQwl2EyUSKCIGl0+wHBIoYCUdimvOFO3eCjtC2tIdepdLr
tgm37p5PmICFv9i3c0lVJIs1Xy1WVCivApkl2iW5W7DAaq+YsNPulZa8n8MsM2VJHRXLE9AA47Fj
nR42ZgjJS5wch6yDsvue4BgmGLJi2NwN5KHlbcRdOuyMyS0SX0qbszQi3OdJLGW6WlJqXanMI+7C
jKzFfxBvml4zgdVwUJpwPkjRQt70IDVSgnurrOv5YTchaJlmqQijUaGXwXJHPQ3/oVxLOHJZq0Yz
WB3alpKeymwgrijx2orTZ4Sk1mIPWka1U+Ce8qR7XnlHiZrXFMasSCyjFblH/+RY11nN8W6QCCff
k0ATxgw4mjNT4SvHfbqHBcXpjEcKHAFu5CficuQMrnVWWY9DRL7yvTJPEPQIAzigEYji0Sx7+IbB
WqEbdf/E5wJygDL/EZ+3+sBeHrDaEXDv+BgzB1hq9FECNu0iq9zTIjCHTmrHLVKfjk+xWzf1Dapj
9qsmy03/75YLiYwySg2U6ehpVvu+c8LvWo2yn9To8gc2FWaqus1TOQJSneJ1Nwcjxl6EN/ON665n
/nuCSTmfLzLC0tCapDt4yl9N/o9Umou+rleSl0bH9Z9j6XyuDfbPbyoUZjOURnUB3pqqHv83ZLw4
VEW1w4Xbi/J1LEDduIMn4Kwy01yIdGx/ll/UWTCxoMbwmsdUgWAqbwQnysUcjI3BLMWv19n/i/J1
XUSzur4fMIsnCFLcuyRyOJsgzOc2WoZ5uLylyGQSCtt3LP3qLjEZ5ukGI1plOqP7vdpnNkeyrP8J
o6DBc6BfwaqWoPyDhORO5+r2knw7ql3UruV5jiK16vnQamAqcp7pzqD+RepnL46YvHuyEGHsGx1p
uk04dcA7BrFttUIvJEVudFZjqSt7p/EmOnviBgZzBTZmhGUgZa76oqt3jWN4l/rlHWTAg2YR2+B7
+tOoaYvFwYPhKfdeQwavVeJG1J8bsGOX82sMLeNZQ8et+cjDYVt4AlaTlYK/KvWPq+Djs7YcP3UF
PTsgGRFcA9Q6SOrYrQ+XD28mNNlb2UZQ9/738U1B7XQRK2JlQ58z6OD1LR5kRDrJF/0WUHK17lEl
xyayrie3r1y8Un3HDeW4TtgYvHYqWObTDGt3+ZPu0ncHIb5BDCWjDqtQNrupORlPc8t2a+BhjdzR
y1BKICpZTsiho8hBQo2LZcX6bzfIGnwMjlAdx4rRqYuV1RUudxtPMtFeqTOi9hVBO2PkLQPbTiOV
3lfkTJeRh34M6pSPEtbLThQhs0899QvTVUaA+/VDKyzcFHP7ryML9eqyuSnpfDA3tWhhJRzd2fFG
BdRl4iH6qdzu8U4mH/EH3rVJluV7pK++i3E9fH2WAy/+Ug4kmG9WhKnJnu1D0ls+hKzP5YqFLxeh
ckXgq9TncUiI7wED6WKC7WTqGqilLL9PaBPxQU/zOuBhV1NJl68sHLVNOzWq98nen7uXQWcmBvAZ
GqEDbO05tT+Wy6qQjMgoOkNQqE0D+9/NfNyfXpT0MeuavfUr3ObfIq+hvcKIcOvwf8X/ssMVhVPC
sAAdWlYUAOygbi/xZebSupnClfZKc6VpPSKB9y5+BZqLWUgOhygzxHIBdHagXqajyHYJ1jaOjwFl
GNW05IJUa0kQKB41X+gAUUh06Mc4vQwqwm4IubkNgrqx/h/Xtxv2Idy5f58TtcOCo91D9+ZBw4eh
BQoFsaeYeVad3nV2ahv+xAeYDX2gHx8J42yn2UXL562kb5uAVxxjsuFkGa5XU2kshmLbOupYCxsn
+7Gs4Tjiq46ZbyOoibRcxp+aoOtghgZA9gN26Fz6J1wafkd0GGyF9cIdGU2T/i9vOKSzqP3qYBcQ
MlasqML92K5GvBGu3LoyZdlq3KE055xBsyFkVVqTsr9PNfjEi/+L/VOx5gxC2svqPOyiajM/igKe
DAT8qyTwB/Yk3ObxNklErxUGYsI6JamHDCcuBhLkLD7A/hLs2wb19qS7JK1nsEfDBVfPN5uHZm7C
24+s+9A9WT8agWVL96yiH2A1GIhdrOWYDu4aAKMsD5jg5o4ke/HWOCXy2avui0Db1gPsIson1WRa
PM3+mGGG8Pp+vi13//qTwxLnMHqvIXnBPdp7szMqhd5zi9z/JBvi7gKfW5W4y/1O1Z97G1QvcqJz
Pp/hoWzGc3/vxHMxbYTwpJz/LgV9KwPTXFuNfEXMieQVz6mEigGehmtKNf/j7qtAPDGFhXxyp5La
OaccycBlnzqyWWQPgmIvTOnb6MpOS7K0fjbk89W/NTCeXRvNXnF5zu1Va/2aBEmjCqMN/F8aOw2Y
01QSAUUNcOkzmw9SO6Z4eWOIluSm93QDahY38ZGKr86QOmnbGm67sdyuuwLbx6SosaUNXLESY63i
q9WVmKL2laIiHV6ymLwR5c0M375BOnAIYY6a7cRI0tLJ0Q0zOQ+mvSR2h1AErYhiysZsgRMBVuWr
CHRERMBs7Fm/+oa15YahH5GQ+CWcR06rfmZXHMPRTBW1a3rnkBZlrMuMm2kCZqvZKa7OSx+IdaFH
gH39t0YA5UzrEPheaWdYBahA95EZgQVenUe4q3KgJrdV1LQU+xGBNhEU7r9RgzH1M/MqiUgQEDh1
1vp59enChbEShj8d8uF9vPXnhODwbolwkEo4TNTWW4jHvrWlxD5aWRi/i+G7kbcSazhoOmrhceWN
KIGFuv606yo5Sgw4oZenX+odFGhMEweaA++MU+OVP75Swo9m1S0HsJojo16ctcd5nuFAX2MNzD/3
esW8EOoVyh/EnVbtApfVYrxgPuODVfpC5McumkKElQE9cevIaG+YM/m4MALyC5q+f/e+Fw2/9v37
ejlJm0C/kKvgXKnNwgq94O1ojStvB0nqpculAXp2WRJF6GZbYeYOUbR1PsF0sWkDItloJHirzOG7
MDmK4/RdH1l0XBHRYSHWSWwlubIgCGZVEv71XcRx60vEVOygLAvA6/CW8z53xhkzm++dmuvbt7HK
rlvnmz5wIJwE8mlwqeVcZ7qxrING7bhqBbeMQ3uewkvTZ8j0eYyifigN5m02xh2Cze2UYgPUa9Am
pTpvl3PwFIrWqV7ZLGLLX90Fqg7JLCScwuyyM04YClbk45/10wc7vMNi2ZzrfBSGNFoQ4tauKZC0
zSbtjj0E0HWFRxgPiooEwWRO3CqHMJ3Zhbfqr9/sM76Br7JfxXxwGgFUlUt9XoXygngwUvGfutJH
YZbe4vh3S3MNnye5lIsrmkX1B3cjecx+cDkCOqNDCYqXaqlkC4O99i+X0AVQZ+0qexKlUA039qWm
cX97PvYtamBFPbbcRhCIEoIJxmaVzKXShrKdDQTP1RVOwRm9FB1aONlOW3YlLmqTNpK6DUtGkT8f
D6T9Cr626zu3QWgrn0JmDJhVLUrQ/gjoqOlrU7a+RfpPdUT3012zcpskX36UfMcCb/ucdnQXAw6J
MrzSoaVyAaprHNWNdNrdrNCDbagZ2I26/mskmicKws1hikGbjRhBnlT6XLNRgKhPUBtRT8WayX5P
iMeeNucTGZJ5gN/6rj36JKoVHm9mXbdxZJ267lGuxjnHgDHn8hd/qou4XQSFlDI2Q0SeLCjJjlQ+
ZcaQv+tTa6/MDuy6Vcm0p1JUPP9xWKCn9pRuJbFIfCvTbJg2GLiUulfiaY4K6IQWTUJ2FvgRMWlH
UEs5CUjfXQeLwdSSDxSYtXikZvDwVyXfjzv/DZJ1ucx8AjnAuHvVtgnmgpcLl2ginnZdiD1dqeCB
fm6toLy89xx4tLZdXrCeBr1YqibY7qLtiG+OkB1H2bWyPLZTG4oZ1XpMjYf2/g+nHmoZyyOlL778
1ilL7/cc1ogZAtmChSC1Jg6XQ6VenSrjnt0nt8END3B33METzHRF6K6klMeI62SVFnE/pcwg52aO
AMCf9cJx0lnJcKCoBldn8vu6eMn8afbFYwACQNVZXiDsDNTKocxQDdP8GFXbZe8B5INXnf0n64af
RnRgdYbZQ8aNPAUvIUaO3R7EBEnJ5bzHX7j8qumpjoDXxMjkWngQTF4Ckr6xvcKLHLCXeqeQyA6Y
4RgTOM0V5Fvrz5bPPOusVC484iskI/emVtULaVcANe4U6SWCfB5CPxRqMEhPptr5fzaeXWoN0eXQ
+7nDh8eXFXISnkTLdsrjJec/SDJjvqxmuhfKbQysPAIT26GRX3uY9hTaBKnCLvHkay2QzCiykHZO
MaB7+MMToDqrEyFDBBIpqyac34oBM3PgPirIpMkl4fE8HeA7b4iCXdHK8fCVt3lBqV7iS94KcM56
rQoqPiEny6/OjUHZiwDTfpuWZyGJbk/5bAQF/EQK4m61gIyTelrHQEDgV9c6uEFhZ3y5xYAatYEb
34y44fDQKxsxf3N2EY9s7KuvF0eCGbwy+PwTIH0kU9FAlkbsRwDrQ5r5McbEW6UjExgiPdshTTwW
vGsQNxoufgmz5poyzJ5xJpOldNzHqOr/Ct5b3eendHk0+nyGJjlFp49+Xpkz9bhf32W6gCutZ18j
VcAisA41eCzvLMGV6OD4aaw/XpuF4glInS8T7u1B/vSdtI7i1Q/aROaqMQakO5KAVONhEuIi67J4
9vSSFUDDo88+bs9kmWrPhrEUpI8yjSHyatnDHOLd5vcVdN9X4oSdAs51FLYKWNd0fS/MSHmzp3SD
K8oyLYSW5jl6ibol9G265aneQdwhy4vcsBdxUmXxiDblmlw9j9DdjZNT1kxJ007o7/7+BQNk3Pza
DUKinLQXRCsncyrAz5URQ4+ZLggwai6yHBnK0amPQZHAxv4NH7bYYrnsD2AwRr7ZIRAlPxMHoN29
8D29Eig9mHu2FIZBIswWwE7J+F/UEFCvOlriBjJiTufnljK2mve4xN8QaokZV8Q+gliUis7koezv
r7i1jCF6GKfAjhQOgx7AuFiTmnKkNWqX809/L0kbp0Gh9mPW7KCzAakiSPbMxvmxBUU7ybkp09jQ
sc7EAtzyx8zk13Wv5P8vNU9fVJ1NI6+o5DZbNbeOdcVZLYyxZMS4/UliWOMAZCgTQV5vswe78ama
FTm4YwXNJ5clt67BrinRf2TdLEkuo+7GwYq/AemKX7DvabBw8oMu2PnjE/4KIvcULEZnf1tB8z2s
dvTp6ptcaVbUPqQas6sOOJqTHT/ssr25w7GE8k2ZLkoC2xZsvfBXOOxK1TOsFgxNNXSRE2b2P/aQ
x1dtHZWEOctsIbZNrEjS7JGgTuJh53WmiFojSFzhexRKRqUbW9+qGNRixeaBRzeiZnH/S2oEliSY
ldw2sYfu6w7g0RfEFtE+I4i8ozFqiIupKgZx3FKbunOhHO1lgpD64z48rpDuEDAx0ZsmhSBrQFMJ
ZxZzn6SChblAUoTncIU2/3ZcwDndxnuStjiml+X3+PHDaem8Nu+4v+d6p9nyQHBd5/C5+WWSn8F5
0QpH6EWknsoosvTJST17SdL5fPJr60LSrQvjI1NMCtEejwHcz5ake6nPAlp3kADaRE78+03oaKGX
y9FCw+j80uzoxJjV1nw2KO8BqeDVCHJEbI3O7tJsAX/U2jpjPEXdWiRIqM18r2bj/GVYYZ9PXU74
KN+cp4pBwSbCl9Pw+uZz7dlRJKfK6fjxpkOOkWN/KQQae6LRUdD3XTgsFrpv+z2HZ5hX5P1vE92L
hkAgskdmINBK6TIE9j383G2G3KJ5Twm2zVUHYY4WI1/YqMJFnC0VouDc60NkpUkM9jDHUJ7uUAVf
Ya9xDo0UW3gpjIwb0DnzGoev/UuZFjtIHLE/Wr6FElZuyTyUyN2AcbvYJRlBPZZhv7zHevkgTJG2
KwwHc2VMrqhDOARFurOieACfxkw7Dn/NQQrJUrzP5Xd7LtYBpI3Sc2GUMDqcBQ6hoJelav70WfEJ
UnybEuNG1kw5vUvUHYLyV1d6HqkHSMEec5YrH8ByqSHiS/j05O9EanW76/ymiXSeOWUbRSzSYrVE
diatFJf7TwlvwPkUXD9yu+65UXPY/3+5E4reLVH02JNHIoLhmBvorNbNZkSdGDOP8OEi0YG7fpNZ
AIpGsj2KaqFVBfPwzHYIIdvRHL5VCMvwDeT7Ypn3KXYMTe4DQZ2Qt+bree40YJfnaTPo/aUI8rjc
4GjcOj61tNgssbov8qy6knUeNd5yhUx8oRdBc15H7IQ0pFW33Y1rjJLw9PTSs3gqEe0G5wbLLtTR
8PC2EdNm44s7lxvi3xaKkNzD77c7ZreGCuADDz7fephjpLQm9I0btkr7uXrq31tyVqv6N2fQm8qH
6gBbka6Dj4v7o4o7WIjfqtgPeDuKnCbkUgxXWWL4SSaXcNFG4EU0f/+rQylOnl0n/A1qvNEQFPBu
wTaaT/zySOQ1N8ug2gY/Ey9uIGMaEWFcD6VmWrSQuqRKO25xM/7D4ooPqQ5k5F/ya7qAgQwQC8x9
fvGLFlHmTbQA3fizuOxrcItREs/+jHs1PT/Iry+b2vozO8bBsUCOJzM+q3Zl1piCO2rwAbaK4TFq
pOFEtetJF0noEs1aZSz8HBd2uDIktHZ12iz5qo1B8R+lLFwPx2Ero+dRMBBBXyTkee63x8/J2Rus
JgmPeF6CdGBSyu9mjwxLYABSrcXJNZ1B4ZJZZX8IgkKHp8E4D4+YeCrddr3hJZ0XdEsLfo+XYNw3
tNK+ZJScEj85U02rFv3hBqhAGuLSavfwMIdFbvPdmlbLsRW3gJP/Q2jWOOwWiEW979EqpVJATutY
EtKPKRBg0eza8wJMw9d2aWdBUzOewgo2LQBXO2/I1g+zrPqWilK3VYVnzfjvnnbesXjN/Te/rpIK
GUyPo2UTxJDTzSDpK2fwp4SRYRL9k7wYaa++S849HP0q7DkZsiqmypnUhV17jxdeFmJPlJu5VE18
IHBnxBNQxzYJYcwG0fIHkhub7HiLGW4kdV+P0L055cXhTVR1jbotdZuIy0xCVUVhwFNo1xE30eXL
Y7U27n/d6oBdxsWSUvVygvgQVcfm+f3rSCA5C/U8dmcmrOBvlloW3bhJ+3J/YU0eSF2n0eV8S18L
zM7KNg7yUlRoIaCJsZuk8dnSf5RluZcGhOM+gzwu6is3Oo15QpaJMf9kQP1tG5d0D2RX0uIQ04AF
CMwt/vMFObfRvuwR0HnmmmednSxvJNFTOgMlzAfeofQaB+m47X62dNrthpwNkLoUbCcUTztcuZi6
pQFk6DlG2jOE9+haZi5ed2lh5K5YQkr1PR+1fmiIHuCpLQxwEVuG10/Sr/FXoqAWunOUtdJXqYS2
Xx5oFNjtOUW+KEcAE5YwVrUeq7JBIYNqkJakbgtt6x/Kpei3hPT9XHoN4ZG9nYQK2JjTctcknmKb
gAZ2sSKjJtyoOC23Q3a7zQy8vHsWNTOuYV/eTWYJ5XEHilAJ+kLeOz5Pq3uYaXnEvdnuypChUeGc
x4LPQWWcfv6nuN4MFTe4+ZcdJIUmcpFL70Chwi4Q8uRNXPQyJa8vItZUSIO6ul7Tb4Kxb91VmJ0Q
yirTINkFPTHMheKWu2t7wcgjIRwe/HsryTkc6h5onVj3A+fPhsVajiyDbutV6lNZsXEoTDEchZVX
qmgYUWSzZuUL2Fnt/oXol6SseS/r+Q6VBxBbn2qBMEU8wAz528+cG4oH2PBwZ0lKwwwImWLtmZ3S
GLu8XLX+ElvvbKhQGZHQ0NauQsemVVH0xPegSLjRj5BqdBlZ7lBvydvZyzCynuSIxsVdy7aWfSYv
d9y901NnN0qM2xHrkNV05+mvO/mdWnngh06R6uQ+ki0PYYYnPJAiGimx0hyimOc7G2Rvx9wgfpr8
MXHXY3LW+W2/QWv075RRiYhJyvHirCBLFVHE+uRYgQns/R98Bw1GeK1VtS6QZav2Qtp6Pf2LTGHw
ch4R7mPuK8COEd7Auz6kxAPJufPIlMHnaY427tA/HaZOdgTRRl+Ov+0pVyCV9xtCQjl3M9tx6QCi
HLUmKgH6SbSWLhzYSxk5ZvpO8MvSQxfXTg2fvP30Ou57BwYQiESvVMEMKnx4wsHn0XxISXvf+gLc
8ShyEE4O0Q7ynvtboLaP10eAxEkd46oJ7e4IWqHkPQzcHJF/Qn4IxeL4dUEAy2AB8OxN/rw/eSzy
IWO/G26FGQFMNXfRVAt+yllQVCaQAyiShYuCIWRQYX4K3RQf3rBfBgcJd/X5S5rRo0t1ZRIAmIG8
FSmoIY82EQ/CTO2xzX0FiMRr8KE+FgndAJKicKUQMd+jhl9zAOvxBYQrLMyNfdbxyctbplkD4FLQ
3pPZJW4427/IRPIz74Sd7hT6nsutDBHw6fqunKaA3JkloZgHdBd/TRCrV6PXWLBgDUyQWzYf52+S
ceYlS8keN/ynx0ZGwAgh60bh56Xf7v50KM7HIVCGcwxq4xCFrD9/gNozLfWtAvYdUYkn6ixIHyQL
f6zdV0kJdmfgNScKWJveCyrL+320T4Kk4nOP4UtjhzLrGduGYvBhaKeaEiJ0mLsDMli29HzfGAu5
Xijwe8e6Y68VjgqHqPnh/2nlQVOfDTQ3LFI7nNhveibMbjPhCBEiFLJup4jCn2ZtqX0JMNXp6rlN
JEMbPbryrCQt3sQvi80XSa36smrKTZQkHlepePYp96ySyNw3hixC975N0FQW2+04o4kHMnzAXko9
isV3opVTnNP7/Ud0Mv820s4afkMz/f3npgOIvTJ3BHAFrwUab7DA6yFvwmHN8NCd5s1vnNOfhA1+
C54W0cuLtD2fnEt9hib/1IKjX5+uD8QY8fNvc01gCiFVBGNZqpj++3R53Iu+0TYXzqAPoeRpO8ST
Ulwe7lLoxSAhypL5v3GqM9E3lYVEMqpm1i2n07SZtKWO1O0gPBDfPreS/dDZUHASUjP/HF78h13o
8p1cueWPW8esW6KUmEMPXXQXOrZY4vVcRWI9/8MGh1RlfjfskP517oKPxU93I/KXhnfvC8BoHMMf
DWB/B7ww/U6+Q++kG2GhJ5WKXtbj5ndpQJfZ4FHo7IqslSqdlhz8IhDi9HB7HXbunq2P0L5xQ681
guOKtVjX+qEWW9K/xdv1xZJoBABomlYcfdcVZ9Cj2tLX/QiWJLeM2rvidicezVIUWnydzf4w6J+p
8kHtSgm4ses2qcjQVdYUdfrbOq2vMZO6KXroMwLrSmgYcFFheLQIo7YV0u8Bp06VpdnqY2epZ4ZC
QUqY/35dLquahAFvxyynVzjDihb3pO8RmtdWpg7+M8y9DcdEFNIuSM1bRg+B4rHW/8GPzdTobbHf
GDIm4STjJTRpfH1NQEyL5QUkyai7ivmB+B1ztG/2afVW+PF9FzEGwDthueGJR/vwnl1GmbHYKvpM
NwU4VpEuGN/6A1DrHow4nVkOgrDs6xuHlG35XtvUwVO0quCpVYWpfC5JnNIddGnNVcACpwI3UqWC
Z4R2cvSE3mc1Ex5riJLQM4vkaYlTuj8CY/H4yD/IS/3a6UW7M/57aroIZOKjqaarFwMsAqgINa/U
Kr4ryR22Y3wGhQq0pkFSAOAJtjd/JJVo4zNd8XRHc1Zjc/ivMb+yPXQ6Vzmg920tgBdNpu9MptN7
VS/9NfcO0yqAjoMw0psOjPzj34IhzFLXpHo6g+P6vea/mfMYm9lbHxPKMnx6odulX5NzLxdKfg27
Vd9oABMquSoCqsEzHH9sD6qo6eFhqRAPcIU6MF0XB0s89p2PVRsdNAbmFE//eT43dpjXjPAlTVPd
6wuS3bwvFPaPedk8NUmcsEEERWS2G3QYNAA7EjuofMS6km5rtW+WMjFdS+Aqd/qUWvE0d3KFSu03
w8JHBTPn+68AnKoTmZUcNsNoMoz8cT3HJmzypo+QKd71ZL6jRLsGg86ochyKlsPqOFgs1VX6U8ea
Ns6o9pezYBS6D40uLV1E+KvZwZp36T99ggG69UhCJFxqUDLeX2RScArLLpLq7+aqYU6XhoTtsjcb
utF7GrVhM57ycUE0yuC/jQj7QdQTOVO7l6r1PkQo5BV4bdZ54zqp3ySxBeBaVIiCfGChVK3xSb29
gDuPi7F8t6WgSQ5j4x9tkXg7Jv9beF70xIkg46j3+jjnR/8H87u8ITnjWBerm8IYcfXBAH6VcI87
6fFSXVnwDh7AC2IfYoJf/pDnioMr7OqhNQ8k868bTE3v27LRUt+3GsR0y1Pq9+TmB3fLvWXX/pbG
x+kVbs7JeQQV0wlJCyOlhIPmbMw9XPuWaVxV7kGasgGKmeYUThT7oYWogD6d1rKavK7fPtc0Z36X
YElCKMmUKMsI+JtCl33oQSJ7WYmNYQFRIBqUFTrfeFyIl9qV7yF2UYSC13SOELpsUnPvZQZHtbhZ
HOKSQ6SNsuiyghQjw5Ojp6MQK0Z4Dkcz8oVjeiDUFg1X4DTtonTcbLzPZ/iMnnE7rG3DpbE/k3Db
IodcR0oK3ogvfMX7SCGdumCm4lE3nHvUXuw9iAHVvdNPediKh3WJZcBZ0kN1827faovHQ1+6psBv
a+mTP22zxeKqnhOyQkb30OwXdM2yv6pveuywk3+1+VfG7sjRfjYS7tyaMJFK9VeWN3vAAZm8h+UY
8lWHR+fRipOkPDyiKGjUjzQZsYrl7lyNOgqYtnSeaSB+ckOYYbUY88TNEykFBIJFuLMqJVBhtU92
lTDlNT/jSFrSv93Qy/uYdCndNCROqCWtlohR36V/017ucIVC2d+py2nj80IGn+IhkwShQKaXLKOs
0uw2/HF8j14/Dpyj4Dpo0u0uJECXLN3Sm6ONnkwhzbTos7h9UfV0qbIMYALlX67Tj+zfGA8k7l7U
bm0YC25QtNevr9h6wHZyFvEEyU2Zqx6GCSxtxdULlmQFEzWckoXwuBnYNU4FwV/0lYvWXe8mTsRE
/g5itkSsHX3+efzqUuR+oLaoYncze+TOxFJNgVjrdvYxJvztZveaaPyM6JDNGyaQePk1bL03PlK0
q68aLlnFuz9eKM28ZozP5zS/C7NEd3vKwt3CaUaiHn9aLQdWTd2VS85vkAykhPUPseoFth2/TwW+
hTIGudQdHG7iaENmNGc2BrZt0TQXIPg2EOgDCSgMyK0Qp+4D+wuPlX1f4ysasweRRplu+p3y1Jud
sk52+uEblDGwtjfJRMr8Syi6NN1WAt9luB/fyGjYhImEp7ttyOvvxvx0txeg+SRvxCCEmY+hmckE
xNlx3H8tQCEc+5P8ijZvvhI56hlhIfDU6/KzsnS3kGAaCdgGN2IDQk5BbiE5d4lPdci3iDRQC4Js
OONyqo8nS9zWOj8yte35qdZW6twc5FgE9yjlMJkmlqnvuJl8RJ6JxO/i9QwEG5nCPGrKOunc5tlY
moMyQxphF5GwWRyyQLFWbc8Kdib1pz3jhSPRbJ3Vo4oCoY3xbePed9FU2cHUBfuqHGMbg7PY6nw2
svqyB7g1JVebFPAES1VBKAV89U9p32zwpxEA+VA13vnf4BjHLFTa0v6zjBnUokJ6xK719X9LB2Sx
zdgHNzEi8fvo5bveAZOgfRg6qL4E24ZUw5BwKuCjwqM1Ci9xsH+MeLV4FHmUF9mQxz69MZ6MkbyQ
O41gVnIZgqnC1qyeCp0T8CBbmU3eAkgP+P/evMd8PA8E1vkOgu3X4K2Q3+Gj+QpPzcrTNH6ZEGUg
XSvFjHT6i5eZ98brscBpPYawKsW+U0U1bXbh8FUfp3AxuYv5XNjrXkbGiIPHuV99BRhxaUUjiK5X
uqPj3CfSNuLoM3B9mzgjlg00tGz9DjPR7gp8osmbEwQsZr6T+2qQdht6rT1ErlShCiOlubbf6wzO
Gn3biRxhL+Q/3TsEBNe8YeBr32iPzSqnjVuZd9koVzB9omrwmKRO70+wqFiIpaZrRC87BmWEqWxg
ToT1HcEJMdW4m9N9K1KOrsTzJws2fKM02udqn8T2w+Lvw4eS/VChhA6RfnaQFAC50s/7FYhwv1W5
Y4rYhqxmFA3/i/MYRAbZ3D9wng55ljl1+Zo4tHLP5+4H3t3AyE+W8kjyUUm3Q6K9++MGMkTSuCJ8
XWgdDrhxo5guAMefTiIWoHzLoxRz94F+gYYlkmOZO0qtp1hO6B8D+F+5CjZACp2FS6QCdOajBQ+n
fre6ejul0S9G/fG5oA6SvWFLywEGD0zcB9Ode5fCfs+VhS4lo7KqrcjtpRW6whnaYovQN3tz0DGf
nS08cAaUzjoBGVIaln/z+F6b/rp3Sh8bxiJeal0XEsiJlK8diXnlZL/gFbPjaXVGI+6w3tor8ehk
1cNTGZDK38YKxlkOrSD1B8XdrWfbFjcwYOYxL9tQiWLlcqkY0G8Dx5BTULZf0VmwBEjRqfno7iMC
E8iPTRg3OIapK4UVAs4iebWtOrg2Xq4dCAUo7ELRYcWMnfy30JPf+ew6J8Fbbre2VAdMrBXhbZVt
W64MVQoG+724DzqaXkx3J30gJEGoa1cF7rE7VsfiCPkGzEyOBhcL/gWdmHmMP5/WPW5V1RdM/D1t
hQKoNKoLPu8xd5eUI5Udxr6ggPJWZ6aFhsXZy/t9xOlskluKF9SK+kB3vVAitzO8l7Py7Zvpqqlh
HGrYsRpimziXaAtUE4XmpeWUK8edp16a16CeuMYPwSxqVyUBlXdjC9TsjMGd6CgoBBt9XAJHvjq3
3ewrmevEeqsF/Jh0J9E/2MpQjQKAjGkXNi7L1tKPTBfkkTPK58t+LctRGpX2GRbOS41YvR3vs8WW
VD8615oe1Kz9l/+IjhGtkhzqSs42aTC31Gy2SWketxVq4El77kaY4O5MusNbNqM0eDvfIK0l44WB
XHbTIprTL4AGuRjZdCWffRnVB2+I6xFv1TZtmthbW7CNsJiUBgoPsr7TAfqSHeJ7kcu0HZdfoWsf
g1fjBKe/KgaI7x3QANp8FBaAbOpTnI9LMYQgjbwgod3ybm6hlpfIW0FNNPXn8SrvrgPqX0G0TxPP
B4OnOkwAKcMzA6vBPMeLQMmLd3+35XlOo1wNdQ379ODo9tAfQPoFO9Ruia1uoxZUHm9Dof4aoSUe
k1PdhgWzygMBEL5ruzFUKKfsXtWVLZ/uaGwoGofKJenTPsAq/c1a8mrw0rHNnIBqqA1rvzk5+g41
Djw1rbkA3K8qxeZAJj4qisiwvQ1XYBi/U9p9ChoSNzMMSxXfz4B7+tgWS/QJmB5PC7HKNwgBjrMw
wXSBBiZfSpiDb9sHGDgLxoT5hJxg8kSJbBxGt1GWOKih9vx8TE+s9cUJVyByq6H9+2QxVpoA3SWW
8+cRwD68UeNHSmpTLsWk0XKjq/cYd/EUUYDNuxBfIH4m/Ns29Yl6jOIzGLvnOEXERIFcXDL+dDX8
JFucFf6TVzMxsbRTwKOmKJwbVGtnVhDFlnzFGte76ZOyCSiZT/qmLre9TpRJuKRTMRfD8mHc6xUO
BGQ886s/SPX4VGeuNhZgwLkg8xPN0GR+02QVIMlPGJlinjk25pUt7YfUIIUjNFE8TwAIXuLpUT0i
4mZY5iHlM4gZfLgDyDe9YMvpASJ2usZmamLhaLDlI42gkVQq8h6qaO2p+nXy+IOCUibM5JI5ngTi
c9aFTiY3WUecL3vQMV6mzemXpxyrqj0xYc2KbwNgTObf5knbw1ASvWtI8efz1GDPcZ3Iwx8Pzjf7
GeLBEh+ycm31NbpkWjzgg6uPp77sdymakIuOZlH0a9dekGyZCZUrc6SHN3bxgbgXnHG1ZByPf+Ok
Tvp9dIMO0sUZcheX90S/kKdety/EgdRxIjuGEqTR3Tm/k1N0OuNjpPvPh+gox3jhVEKO3sEuW29k
vFsU+0ekxdpd5iySY96t//bWlThMZW51kZXPYNSf2230+WbtQXy6Xwr29XGHlBHxHuARaMEJYiwQ
SV6i4agHSJ0+KjDgKfsgR0gTYY5luVyiPtwR/WfvoXCM0bUcAC5TP17Q+6qgJy+4zQWbqfRL1e0y
EUaESWgYtyTgPtyKZ9zNlexHFZvmwfOcg6Dp1EXeYxHV+tk6+xA3qNqHj+ISqhS2Nh0A7ZvbmPqT
aTWO4fY58z85SkdMqnMzIJ31SWwjIDjTsdU+6Yk/JDrMaK4e7kFqJNjHCvBey12uNjD96DyNRMVk
yvMJuslr7OBvH7OwvXh5YYeRsFUb96Sq2Z27RFX+WGIXQe2FsefTh1J6kBJiZGC+89lcjy9sQF2M
P9KUUTAWDvrbsqqqtjx36erwdNfGqwDPSckyMpC+b5blTDEyaYVM3fEdT3ta5VwPGZ65pIcrstDK
UkdJMt33BVvwRYRIeIk0RVXkOZ92SLOdB/kEsRlV9J/zyp47k1RjXwDw/A7noRcC1qNC8qcy70MC
Zy30VHhq07IAGwEOudW3PvUlPkdS0eoAqmRmB88rwQzaeKq7FYPDFPMyv5jy9ltzwfIinHE9IXmw
cFbMlkK0HkvaftfsEqKir6aUQEDWw+ho72oyCjKHXsLP0gTZSV4GBI48GKaLYQfYNtBO4APSj5WL
MyqyudnRbuDWGxXEUhfVJj3JldyKq0AzOdAsDTPdYfGUaCSYFe6jfHouK6J0w+dWv1ZdQOIE503P
zYnvz4yXukI4cHzdkAlytFGQ3jLWa12zDBXn+8t4mxwGS4A/xmvbkRswY1KQYHj3L+bvBYt8mQAK
AX3dGeTKJPjezi1JVJzPcZDBkWUXfCfHNYaLnIlQQ9v2eQnmpF97+Ga1iHm7ZM7d0NlEon5sjxoT
iW1VRJatyIXCEPf2UhdIdL9sA7AaiC0B2Lbl5ru3gxVSwbQltJRvGx4l8kZh6B2UFmdpmNXocAvk
VeQliE2rcMe7NtBaiRnjt8QZmfSkMJCoVap4I8n+M5ZMkSbpgHx4vKA9Eu88IJYQCg6cOZEkhj02
5um7nJOfBbtY82JPDaqiq8YtCzgqhvzgAqBI79fagY38r6WdDxI8up0v4Fx2pAZcWYdlctxq7Zaw
rVhMMgMqnC+Vp08aQQsPTiGTlYECB/+IjDMjQQHJQ3RiBYryJrd6QpjnqQwb/GvexyCHiNO9cqsI
Ag/QIPnK4x3SOovv5nlX1wnM9wataN3aYRsurIACat3WSNFj7XmFTabE3izOQfZu1uWGcr80Z6jE
8+KIUKcBiiap/uemLJGakUe2XyJX/T20LP1OJceAsxikhqHOLbn1b1GKjLWFy35km99O8o6AywVW
EIYD/JRlVrsHnAyQ5O2p4Ho0Vd8Nusbav23w96VXOJKDCU7LcR4PnqNl48q/TTHnxtcR+OLJ4btX
vR0V+hz3sXop4H9GraBhF1rSMv5ZfqKAE9Qd6IKbwXqJomz8OLr4UxpX5CVYBHJcNbNhIZyUHDZr
Z0sQfum/aV9Zw/XBamNVt2PREENNmFeqpA9tDQ0XHtID8mnyhiEqbxN1WJtqwWRxHndFKRKyHA+7
Z62up5w/b5/XmjhULF13RIfbgmTLCdpqCmymLthJvH/CNvsmA+oP5YUBvRbTkbxs3Edn/1vYIwMI
Gk5uIlGYwCYaqq6NOytTNzbKkRD5Ek7dYc/2HG0TlG9Yf0Ps3llcpml305bC9nHdfzrsg6Dp2oUo
uFjjE6v63BTAmWMHI+mBMqo2ytqTMIiQFwPD7MJL/fMEmyoBnU5NkyQHAqRo0jIXFzQ7lxfWRM7N
hRh/2QguoQHTDABBnPHA5dj1rYiqX7b3ul3Qffcrxk6SsOWQPNg1rZ326RBtvxfEacSNu0y2uEg6
SZM5lilC84KLrzoEGbrbs8UZ3QnsqU+zB7JGLKYX4Hs/tOMeSAcPDsIXHf54B4C43Bk8XmisrGa2
1529rit+LLIN3jdgqi2Fs+sQ9TDeyORz82dyvM3EW4/L1QjJ4AhBtc2kwKr2uNFA7v8SxwY9mNW6
ze2xazyg5ihRLNp9rXvh/5s0/MfJN197rI2Xa1YNtL10zvFdlHGsaL0S5JaV4mw9eBnx+StS80bd
p1oic9WjukQHp1i7TDJ7D+pSNeZcExqDCGg2pD8VrDe6RfkMIPWfWuOW61fN+FDcOrMUPMwTHQnc
vKlYAMANlQ7g0CGNXyDQnCLqHPOs8hLt0T13tfAAsh+ICf/peOurDOfbLgegTbNsKhiklIZISLJl
GcmJJTgqgClqZb0VizmP4MeD305bsiaCu79/oHCOFAlqffjT1HzIfJw7PTNi2Z45ytrGcDPoyc6b
VHk4sozgFhy27ZIGskfpHLi+2fZsFBGbCAaEUROY/cj78oPcHO5Zxygy1eUSURAtdTRqAD+IITBc
oBKgIqCQSzSDucFCQv7NJU/puIRmxpceVRg+MyjvJr+QA5awebEXj28Bi8UUlFBUWlgoFd/YZXOB
Z3BJtQmwH6ya++xvzBV2LxRJBHMCZDQRialvqimnB0VhXs0rUrtuVeYHMjhrfoAp6k4NAT8HwgTi
p6mgE4wdALAlefQr1ywQ1B6yBns8WRUIrDVK4z/RsutrmV/NUn6GgArjZxTLiq8xWCl9EIw5fJer
yte758J0UK9Hof+EHd3p2UsacbdZ6A45ky4wv+leRO0IKavrRF7ocRH2a7SFD5rBd32OEVKE3gvH
U5cVgrRZ3Ovx+V3ftop/CyyN9acSF+aswTNHgqxzF3MtvwHdNC0eQcuBPQraGbC2Wgw6Nq6qjruw
TwPslDt0I4UlydqQO5HwcqVdtkkg1/Dsntu2CGa9FhZj9ni7iGsF6a8fTj+ujmy0KmC9Wqzr/N2t
UZqCEUG3/wSpoVQfkGyDmzLgBZq3pbSXE8uKDAWIxTPwE/VxjhdTTMazepGQyi5qgCicng/Dz0vn
Z1E2Y9NhOd5G061oWTgHSsDw0y5QenkG1Igim7PEqU/pOqYPM5rAP0m2r/CfFSJ7jA3zgjtax3fZ
/m8jdzfMgkFsuyiWlgBmRHsodHCacLeIwhZBs9WxgZlfQFzvZ+N+0YZpOSDnp6XftHwptfYVLpkj
xZlW4fRK35/HbZYLF6vktJiDBCOrFZg8iiGTTF1MOUvUGB8N7fPCFqomov4J3sdpReOpJM8MpHSD
xbzS8q0AM8iHbKcShl5X5LV4Iaj/b0z0eItkEfYBNJFQMlUUH/rEg3fk2zJBIaRYS+vJmeN6H8W4
6ELXF/7m18ulqhZvs62XfF/WlBrC0wLMpN5CgPFeAnBvgq6CpmV8QYV27v/SR8vEqsyRW10uYRkA
MXXYxPGoeNOOiqgBQ/5GU3LGX2NOE8INPR46crONwm56Rzcs1FnTrr96Tod6GGYAjGUPzgkAdTXK
rhZap+45aFChgzgN7M3Tuc6NrDJai+0Ir5Hu2447bPrvsGTbuCwgiIjpTcKcqAlpiBmHesVwCRtl
2DTyE+NAt3LLSHBEdlTL/v01mH1T6cOokLIlMlGqoiLQuxE2cLcrrCvgcOnEuZB88svAo15Wdnw0
L+5Jk1Szbv1Sr9wibFP6gAAtdJGMZGhrkI2SNvQGWsAMAdqk3z2Jh0Eus9Hn+7e5ctcHRYI5zdA9
BM+eUOZaM8fkPK4WLFpoU7oIc4qg4BkkCMX0T3nBZLmcBhNg82i9NhL5D/zEMvPIG0DcvtNJeLyV
m9euBrMrGGrov7zJk95RRxE0WhMkAi8ueUceZ1SfB8uWlCRu24+Yc1mRIrtk4Uyrl00o9fmh9kH5
YckZQ9f5o8O4KpGrB7Kcjr1wCjx7ImUTMv7GXCOgmdQApNRltuqKD8r2ZhIy4sPoD6sANhOx3vzs
/IHAMyFJE+rq7/dlUkIWktv5npTR7Mq/yfzXhbC4vDVAcjrjbjVdbFQL2ZyH7ZWwBfqcwMYKTKQ3
UrMPl9/9yukLPPWfhiuFjeJ9uIzVjIK//j+39Np/kgX+QhMDf55czBXld6FGPojylDwS89a4yKLI
WD/Alz7J+1toWvjlElJkW+8YNquwE7/VkZAAlm/iSnUfr2PTVMFmF+tVGuNKQK/10NlKj8p+2t+8
9bc8b0xbkV/1Yj6b0/k5GOZIIn5tX/op/ektZCzZ7FgbyQIOUCAdbxHLTGTg9AxzfYQ1TrMiCqsN
36r9Xu4MUBjIw6kYhMBY6yYsIkOhlGnX+zHBbzdzlEmeGxw7mo/mATEzNLM9G7f3eCmsitfYvJmZ
p6MZ1a4FT9vnSyppEqxGkylg1TSErk59zZml3MSsA26mXeFZd5dmmogLsj2LAUrgGoM4BhXZTUpR
eYsZJJ7bzjSiA3CMEDlLh4DZYN8DQc4bey3aoMLYkNR1+FrZ8mb4wrwC/cEBJKE5bf1E+iwpd6Nu
wBe5n5EpX9tdXvwTIjSLWVd2uc25sQtje0pqjSbE550Nf563+ftTXZAHr926K1H9bLATh+ZUQMmj
MDHpkp21zppck4rGEfl0wscIMJavIy7JcoarZFajQcml89ssQTuMDxHpG+0hAlUpuN3k+HWOCb8t
okD50OET/dxI6lM3H/pHavRCl2xtnGeEoWzsxX1hYlNotJAtgQG3cd3KattQkKGKF0QHBAGx38rb
nfVy6SgheAesExapFkVHvkH7XeGqPaKMQl20idqHvyIce8xEjheOO13rpaXfaGfCx2eWq+3M9LXf
f+U5FDV/hE0AN4QQOX9ZllfWBHeNxK3Ts04S/K9ekcPeeKURgFD0xVPfXrY3UyHQpTirmrpfQ5av
6CEKnFMe9A6Ijl0nE+m0p0LGygf4dxwCcaZN3M10eIp9PAwyI9p/KDHG7e01AP4iR1WVH6g7djw1
4oeGzLwU4E6N597GV199+t+BCJWLuDT3uGpTSK6TiymhyVGIzCJC+rDnpDJL3kYtM2Oty57Enudp
SKXPdghWNfQgg/6O0tzd70vy2ndNrHq59wQjuNFeAn3tdI8fQXlKOlPjPETF9UF40KXlrv+BDuE/
1LbmJzSoTRfqBOC9QISjz4AmePzjBDGV1gWbqlexvKtJlsYavUsIBjcX4+TItL2qi/Kou9jjkwpY
mYdsxuJSeEEUU2R5ckUcUX9r+7FpCo8FvvNya1zx2m3q8SSfTIiaSBecLuzFCUDgHoJ0BwlYAoqv
E1JaoaGvXAizTRUSkNyDkv1jSRol46/8SpYvomaJTuE5bOim4ue46LnZ42g80ty1U2t7riSUm+tT
2i0UIJNuH7RQ+66c58jBoThFuZX31IreefsyXIm2yHJPHaNZGKUyJIExSxWS4c4W+xYjnLvGxNSA
tra3zwMXazXk9DgElRdX21K9eQjQhgcj6uTQRoiqL1qJyok2PaOFEWTKow8jaaaMYkGs6JHwhmcb
6cWur+PMeosLFKLQTPv63WSDs8nHtZm68xd0VWS8i6rT7uZtrzgEqJxJfWk3GYG0Qq7tvM2KQU0H
5nTUR/Snvq7ZARTILkKXC8tC9X/Y8oK3X5brlLaWAAqN9rbsMuCCqN9saRH7R20bXrWMhloJPQo9
EvUVqlH0Hd8fn71d7BkO20UDsUBs7Dog5yfsDjvv5PL8zjHtCyxFy/Vm9Okwadci0zz4IRk/TH8t
CkQ4btGvSbpYC4JByPwV4/s42+T6llJhvLVz0/mbxW7cKcmUKRGCIgltvqRLRW27kwqjoWeVTR3/
WY67mIIrwCEz1BEI2lHfNG9+0XQ7JsL4cYkLfKz0cUvqA7DVF1l1A5+9k4y/vG0watBlv8K5+KAI
Ggu07K1sc9RZdZKzpOgfk1DOYsQ+7EvqcHkiO5Y0Yd33Va+u6zUfsQ5SyXhH5V033XrfYXrlDSaz
AbubGJTaf9m3eOwy+dFMTJCwLWWadu3XzrBifK3s5hyiLd55KMJbSIdC34k2MTGujHA/D/llktBN
BFyjF+k0Vgi7bZK2DIhaUoSS+W+7H15uyfakO6gn74bbHWSiK+VOalfXpa1sdGve5WP+QYpAVFqg
LAQjgGMqOHdy9FVyB8Q2Em17qTrYiYfGXpgr1R7/brvpr8+8o6igM1RFLz48LueMAht4e3qdCCWO
Z5j+E3PTJ3+0TrxL2MjeeFBx8Vp1vvDGgGPW+A1oLbEbo/Jc/Jc4W2tdgJjWIPphRpyrwSIXkTM3
AQHbu9tkDH3ACK5pwPTSOFwsFVLAWN4l/lD6caef1OtalfqbSi06iIpEp4eDcwU5Sdeky/2879Q0
BJ5GRMv18n7OSUWvVML7Jb4VSzrpohlFW6MFw4b9qvGvBBxYXCWQbroMHYf5aobdUa8XwGirsZ8m
1gNBArnQv9Cz+tpPaw4sglBMIYFKOcO5JSy+zwzb35YwkmPUu8mIlhnCkp/ylpz1WL0tms0TOOlk
/PNq7SYxOhO2vbglJKgS1df/UdpUMKMKtxWk1gtx7KiHAddlj7/94wHmHbuOpVc1FRjrn6QR3nPe
PudzIoVUFrKuKE8yFSykvZYywRY+LfTLb3JKwA6SdQam1iElZ9gYYZ5ooHrdHyhkdX2xOb8oLw6m
yCEIT6FKubA5rSgWtkzRBIuzebmHTGveosP6OPxj7ekYWt1HsN27Dr+O/GnWq6oU4HIfHrVnRh8j
8flwub6+dA6HCpx1s1Z7SDLNVfGUYZAnxoigddBHy0la6cKa6+7JRBD6Qtn6CQQMpcqNQ7DaBib+
acIjNkv0iG/EGigi5v4t974CVUMLyRwoTVrccvkoagPRHyB+M7VhbZHZ7XvtqfruK3jNC1Z8gA7P
9YTBOEv/RMBGXxMTnUPWx47P6NzkPfZy/uvXq39EsDN49koEnaUq05yWM2qTYv5faLSUHZ8BaN73
zAXDcL0kvRHv4Q4PAwjNiZd/hhtbZbF5VgKDIttvHKfXugTJkoM3ymrgSHTzhCsrFR0Ip+wWWY5/
wwqX8p8f0KwEyMhKgI2t5A0ShNdhwHVX6a5E3bn0S5N2qjXQI8r07DSkKIujPBx/r1RWyefehO1a
ArThWI/VGFbjqvBJixlJWG33I/7N08THL14hPx3u3aNwg0VrhjBQOTC6ax+RzE7Bq8MPBjk9/hyj
W+yoCx67VqUPsurFaskowmRQ2WGVeMCHD3pysEipB0/iau1p9FrLCPhOWFacjAn65Wtx9eJ05JeC
2se0UQKTtdhzfhAscyuH4/YeFdx5a3h/Sjp4WQrvaby4Q6kaLMxwuAbIep/M+vOEcle+hWOQMQ7O
HVbVKMGQwzf5zucrUCjGfc5vfP7tEYOF6GnxWElIV7y8v6p7vle7SnqJqwlg65+rNRQfiRWqJoCo
tE+m31kYZxOHVlV7WDkPwbcHzj06LXQmzqBp5Fspqyb/jGGeaxUkAmSP/3dGoSFpKUNTvAoLcNkb
m8xz+rmC15PHnK4lN7jCRDczkcj50NtKMDEsySDn+qZf1E5oAkq57USNuOr56ZMew2n7ikBEhPzD
BmQGO2uYwSHgpyMt1ofY4Y41Q1ffn0+SrG+m3frB9pBdmH7mDlhbkKRlNIvDK+Sv8RPXfDts3D9H
qnxDQojqeZmkVoh5MWBxWWhb4SI+IvyxnAikPFGQbS4+c6FYWEFH2yiTFz+SmHQhe4wFtlY9Y1wv
BqcDb4i8Usum5+fzEiptAoNRXpbmSKXGZ+pBz5TZuTYrOmz5GO/xuXbhwlShbAEjYVLqabXCjiQy
MSQ4D4+bQHuoslFievwDpHL+xUBbx/ZKPC0mxKH6w6MfVdjSBI8mofD9Wm+czF5sNIA6gdFi9lnk
k40e5mmDwJMEBIsY7HfzW6IDPx1nJHkB5zUsIoA3eh/8cdTfeij3aeVGHG3kcB6zwYk2oOa0pVMh
XLmTbfhbVvVaWqFl4pGeIb70D7XIT71JECWA91GGwzWiLyWn3dWQSaewpyqdvVT3WbuKA61NDrRa
XzS29RcpBx2OjzXTDg2ce36N2gto82xwaCqs5vxaOLsmkY/XpqorlbBPL6o2EgAKUThfxQZ7klNF
DZ3hZhtUEmr2BawW1y56u+ZKAuX5ieZ/QWXiO0Ku93kI+Hh5TuNI3hiZQBMg0qz5SrJ3NP1CC04g
mrsiTgnLkSCv/ac3W6F/3jNVNI6mM5BKrlQ39qgVJxFIXRHdDhZ3r7cX8iEWcOSsA5pYivVjPdUF
R+toga8wWWsoiL/5Aj0l83xFwnG9cB6xuzqQKJPSvfyqPB17IJiUNL+Vd0YHhIW8Ot2gSO9tB1Vq
17gswL25VerV2kgWcF6YGNIXUBb0/f+hpZ8ZwtWBe8hCM3v1qd+wRp5EZw1ZMOW5Sy/zjiDP+l7U
PyL38zHiMpEIeCfxOGFIenm9nKNTZveA29JkBP17TAHbo1t5iZKuSS1Gg9NKEZayf7Dlpoowr61S
p208hSRvbwFnmXgSr1Y5lHcRSnCLuLhLrXjP3ytJfsA5u6t9X0EHN8J80QJABHdvDfnDc+mPi1aC
3U4wr8UIo9y7etptUjm8+ezGxfeW3fXRFluaIqh04ju61tJuEDfpaYETyV3IN2B1HZACvXUGqNN2
cpBlNkaoxnEv/OvtQlOeZaIdYwkgCcHSvG/sb5sTP/KDBACCIeI1ud1+GNylM0cF2oJE8Qjdhmvq
bqRWRhaKQ34q35JiZzBIj5PXMqJvEfOctvJJ/2cWIJr3EYCb5IHHfI5f/xN5i1KqOGkzubifiJNh
+OWbm4YQg+VkwxDpas2rOmgLtmOQc9f6eyIt4qmfee+Zi7+eYmIRBFXegEqa9My2BQ58Fs2+jbMT
4qFEGlJk+yRq8iESItQ2pJwwVKaAc9M9atUB59T1QE4D8bFe2pkKOPNjhxKHruL6NkqFab0yAKWo
CIy0vL4ZL8AXDGUD7th9iQ9R1jNS0NnUsryoiECobzeB+zqvDUNuOzz596Cn1gV27DId4uNRnBFA
XzBnkF0SY26ivpgTZS+9g/dAQCRsCRCPSvmgj7ckZHo29iN4syle8UfeIR2HJp1R3AXGWzv1AXzO
QZKzABucFRZlq4wFMQUUlHpKbsI9C8eJJ/IpCf2rPL4d2QXfARVy2rg+nSqqyzNTVpZUJtxBQS4R
ppB4m+060mskc3sM8UBgHIFxJhiQEjQ6NYN+0s75vxVPLUP9mL4Xjfzvo1V6zHpORcDm9hvWX6WZ
joT0R8GO1pLQjsuk2T7YgxWMpJnVO7Jj2jDu4f1LOJI778AfvgpQRXQL8Q3vnHKO2oLSZV8aVEkh
bxRnooqKrfCKGZwhHbZVnjyWNr4Ij+1FUo43UxpStYOGIIxy8gdAAqzZGjdlW+QE4UVvKVTVJ3MI
gEGMu6Kb+bT9wD/AFY1fbWZ8er+y8hGWRptkHbj0M5XuR7tjb/gD56UT3ifj9GZXU4m5stTOKcFe
yZrUBIHdm0TUTuVnXv8v/S8a8KknuSRKcJz7pox1JL3AQFQVo2hK+oRMhmSRtkwKaMO7eQKmS/az
Me6x0Wc6RraESR1rpo61CAiNdooVBxHjIdwd1FbLAazmrCbwAbAFb31NiQPQVGd+p2TtgLZtdNyE
rfx9DTpTuvKrpYHDekbSLrjZ52mBZEqBaYPeiZFBsxb3UVQKZLZSIz7HV4vzh2hOaVRBHJiyBtT5
PiEQ8yRSby+KRC01ERAXuhthT4Xl1wtCvxhJbIFIUekeDx/HftGW0D0FRLrQwuGuAYN5bqeYbYLv
ubsJU8zf6YGxe1omIZ7nofRcVQbqtHBjExCvGA6wKGN8x+nsLc/FjADrz4isBvgDQHXEhltL6VLb
lp+vuVOcBbxdLZDetoS6BsDJGkYG1jXfVr248WShGwLW7JjnF2KbyVQGP56f6UdAzpPth694KmG8
PUj2EBgfo9dCxnXcDe2ntiiluco5QhiKIq5B4UavNfFFhGHvXEBECNtvm+wjPEBaQlLd6Rx/Zgi0
ATkA5l+AdN9jxCmbBnPrbUuaKAL4AxPkAXm26ev2tqVqLiDq6gtWcq5/MJlP0swQO3VTYRJzlqy/
ptzD0dLVFvViWt8AkdJGFFnMFZ6Dqf1lKzW66rPs7M5V+qUPaDM/tm6bScRG0AmZ/dAK2O9E2cdW
eCxRikNSOSiuHMdtBe36znBtpCgUXeR2aXoWJibKrLqiJOS7CFeSUecRUd4MiYtub/vMG25W0ZHY
FiTW8jat81pc+FqfJhe4aW5hpeKztR0b7R+Mgk7ecw4Q6a+nDSjNIJYFHbc9L3U4A8ioC5u2aXyP
jOCYV6ZlJQRGDKaOQAW/BwpPpTF6Q8HiDVDmOMJRTS5O/2MZpAcPKcEkPP0orJQB5NcllHnqGoCx
oSY3leCp9YsQwZNntqD0JzATlWkryUU+RyYoksa/5/YSM128WmiWwRX4DhpvOo4JJfHhbKl7CbqY
wGC/Rgf/a4EqwhxOhl4dIsMeJ4jR+VYwwse4qXPPCaoujXhjyAg7k/Q8d6aJ+n8ajl8j1+9/xgu6
0RJOOyVib/ugczlMojL75YiqBgFHUlESPdIE6S0P/eI4vaQOe/q95QYYKXoz8CnN7mDvZvnPuxgW
ErBqdGSHhM6dFJvlhDWhsf5iWNjFEarsf9nYPHhd29zUemfivu7wdoAbsG7QFzCO4XbzTPFUZru2
2FturBTZxQWA11LR+qMvi0/5ghL8TxyQcZ2YPwzH8ThMjXZzUpoCyIbbc1FRri6iRDe54/BwSIJV
xCzC9Ez0UrYpazFqdfVK6xlDSxPzL1fzodZilmyg6iHnfdlQFb2+lfTr13cUWKDZBzxTYQOIHk3D
vImBtAuOmy1riEf7YkVtrfppTSYFnPY6E2lWKEl7EGYVGIsqwYouD5kWcZYTLaVjp/TMJHzlObCJ
B1ewRFEmEhplfefMxBNEjCwj5cIx8NDFNHX5N4LPkeAq8v8W3GDZnKuTD+Lp8G/lgRm+YjxEexpQ
2jV5b3PW0GIi7cJVNTaXXg6EH33JY6P2tTa/3xPDqwEarLpjLBuyTEW4qI5XWCw7RiyLpTToTHbE
U62gOKonsfi9ysRy7mPGpEkcqcEUeXERcTdL5ccvEnISAadCni3/+TsE+Ad0X8Y9NgEaonX9pS9q
LsoA3ZPxpj5lPZXiXSs9kOCdJE21jswiyaP4k2O/DAb+QikIAhtlabVdeVAIY5m9UQpT+pq1zal2
9++TqBbdE+Nig69i2yWTIga827xiEZeKVU+hPWKB/nCvHl+NckLRI3vBLXgozdVvt1+QH/fG2/S4
+wpvsiH8kgq/TO6NA64X5LnnIpkzD49OqqQKDp0RRS52SYi83HsZIJZ/2CVOInKAE06a/uJD90Ud
XST3jja7o4jQn3JB7RUpSrmz08JB47/HutXbju69/JqPIOQ9yFKesYhum6/YjG5S8SN0TlPAd7Ez
GPqLuiavww5JKKTutkzo2lVM7+AtiyOwI+1jC1x+4kYS+OuD4apgTC3Da7RwYJHlMUR+qTUQeIm3
KMM5ZOXt611NzhpNW/3e8pb+GMKlktaQJ0DLKVEAHjaMh1XXlMNDPJTE2xEUW37YJZJE+ajnx9OF
UlYl+PN6IC39MGYZ8CJYaHGdKzrt/uT9onTYlH4IF/vZFlw2+1mn8vyUDKTvCllCEqpVs9kchhO3
NhBhAdB8EGpfUsF62fEMDhhXOfB6Icte7yz37RJBgLtXrZW2vGM39SZFGYcN0T1kd14W7NHtngMk
fGPzS2gUzPlTanPij2w7wm82A13fwNMB6ZWP9+D9+mFud+HYWJyIIrjyrrDSxmygzqhGLmdiw2u4
srthrY3csk8S4ROmlsmhi9RXQpVaJOvdr+QSqYE7sT/WqfvoEQ0vaSerw+MQf94AHYnl1RkVzS5a
sRVy42sI7Amj0KV3iQ+JJL7dLS++kUK8qb/AN+hJX1oOyw8leUJ6C8frYuYRMEBxulYavvi/Ot9m
SdwmBF8PXcmVnCsRUJpE6jHtdFmGKeel/FSaebHnSYg2trWpJ4l23gD0Tu7XGyBqcWgbDBQqeH46
g2UQaAKDY+JTCY4aojpw8IIZrDIceoGCaWbcpOrJNA92ULEzy2B0JlVT9qig3Cffbpoa37WWLBOq
99MRK3t8KbM+vDNfR/oCprmUCdbv1d5sZi7syudeel+4I97L6R2xXGJcWfA7KADsWYgQH9h86Z63
5nLQXbLyRp/HnsMA93ilzp3R0pZUhm+L4pd9Q5oucAEkIpx2k5W67ns9nNPJ9mhmOmdwhtIIyLEM
Y0GiYQwgLG2XZRjfMPmO5CX0BiOAGwslH2JfUDAds2XMSJuOE/v0HB7pskcFSqufzL20tcW3LpxD
q/3vF80oFjGlOA0hbIRjlUBRqHXL1t930tyRAhYou8dSfX7UZh3g18DS2884Vk+cCO3DL0Fqdnx/
Iy3Dr1nLd/lFM59pJqMwXTJDMOOcTSjQ3phwnrfcWebcndMUzZ2vD85TsjvRhjwwzTiYOewDo+yf
5QJ1cynbkbcizbCmAOdXOpNI4ZKQLOvtkSc6xMw8upbe1k1h3zxEGo2zz3pzduxnzv41Lq7qj6HQ
bs1C7hEeHf1VFzWbSKS9uNYLF1/wJXNetl9uAOcQrplLI1/zWQNyB4G/Wd9WC8c7C5wSJt+MP0Ti
1PxO8Bl5hoGPeaxcLo5ti1X6dD1vPM5+jiHtc4y1IzW7G7e+0YhsZq55aX/3VUJMbl8/c9xK2S+Z
elysEJhNdyaYUzXNhOCP+a8xccEeZg72PPpDy9y/a0WQwvFPjoahAvwJYZEkLHdqHXEpxGFPubnJ
+GiibJRPSF9w52OZ4pTRAEsie/WSZZnPDYDJ0iiPp6QL8ID/Hjpz+RD80rysDckqUQ1w/9Lv3J0s
uvvWRvFl+EDAkP5rDbk5NJJNNlEJrhSOuj7gFIrc7JQ8nnmpPRif2VsiI4KTcZvGk5TQacQIaNpe
UheO5LL+oqv3snEK9VkusjEA2DRWAYDVjw1g5h8ubq5yuPXDSlKJvATIzZhifPz33/uTG+WPUsl8
GLElswbXpD+Q+nsCmAJugdlsVpSSOpaZzaC4EuIvxvfF73yyNWnMp9O5hTbYeNzw/8g+b0qxpZuh
0LuG26DNsYWkjQm5FitGx2jxjltGruqKE/3AlVYyhf/DVHaa7jeLHT3/PYdBupy0Bo8FcKizIA6X
vCCugdPYV+2/biZvBSKEEoQ4CWfto0ZIHVjYs9UpWAGhv9UCZVi2z+SbYf5tA5TYH1ck+HqodWt5
jcn514l+IUUTWvdupwB6AwGwiWuZXHqXPuD89AhEgcNb9jkORnvavEBla5oXlmqjUayr+sYXuheu
aGIZe8rtYrMgWGysV1TWahqXGrG+tiK3jML4aNgp6Tk3/q9utMN/O5zUXPrv9YDlQFtjL9DGqILC
WyemrgwHaL0AnAktkr4aGMveNw4ILOfLN6Bnx0VvnO93kCc9rZSsnZHQwt2KKEtDdgRnNt+z2fId
RDNkvaN0F28XTH8kJkNRD8My6T3bo8HDyZIKzCQJL6dg1EsfdHTP1dLW9y3af5tx2sFGoX04uD9R
zV0A+kl1qFAT2grOenm8LBMcjiCKI39yBRMvI/1uRZGowt3h0umgfDIexTrQC+lcnNgGrJzWl1oo
rS4aG0Q+WIbC1lsc7D5ULru65m/uwgkxsRoL81FPe3yYGMluddbj4+xU3unl9pLw8O5mStUwlONX
oexsHysOafGLPY8e6Jd2IH5Q1EN8JBbaJVy+9IE+cGg/hcxklEFa4/pRY1yvKZFw2JWrhXJms908
I4stwtiMI8tJZKqGjTQtP2ZFAXOtlTbjKnFpadu+BCA/yKWRorjawOXMBtPmNMfZF7/w1AyGL53a
vM9jIxe40bhw4BhdiBykM+wGo0mUm9XELAotoMhCNhW9TfH0FRAO3CY/F8OhY+r1dB/p64Ql5MQ1
VsZJ3j5/r05QIOlnNNPRb4gw/LKwr6+J/kAODjPt8UzZmd6NLGqu1Vjde1fKr1fFrY0087e8jFVe
WBmebpI6pYvE3GA5K+K1ne8n/QWOjVx+Zh9QtBnnrCEQPxctsWK43dZ2i1umkiQlwErCGtH5gMgY
Y/MKDvT35Piu8kRXlLy2Od0dy/0W7BNwl2LYOHC3PF13B51dYltNTXnk1r1UEHXNTnYdjBZQ5A+l
Y1fvKkvSsxH0PqDCRnzEvl6pjfEdgTkY+Cxfa50h/2DHVGpyvEdOInzxlWyfjgAv7R63bogD91IJ
nJlNcl3qcDSAKvd7YR5Dfbpe9o17n+JRqlBOC1UpQ5b/4uYna1MUYEhHlDEfK66Be7Mk0dEkeRgw
AiaR0OEzk6REQ1iEHoSVph0a0xRNUKC1WftSxP5FzQF7nevehgyD0qI+KCYHq4vSShJC0Vfnka8L
IzgPO7S1lGZkc76zquOkBOCW34wIww3cZCipzVP0hD+SBDfLXNzERpYLdVlgWnTMr6ZbTrMrccMH
x3VN77EdPF1kPWR2VXRvLArApHjkKQgyniodtL+QbPpEtvpjzLrCu1PsK0dIzETLTrJFv5WNah7B
t2/6pExMNT3N+osw47JlfzNX047Z9qLB3AbBCnh6G8Dbfx1ChyAxfb+uH2ZZFqgapIGaQuK8bLpq
C1jmmFBHHvE+UZRWOs7C0WMGIC3hNGkim6Nb8WKrl8y6irJzrNsgu1TgN3sDxYGpZkhJUp3vJdvf
TGTggG27sQuXBhb20GZl3kWu9LkRmf6Gjre50QEsqj4necGQmnTJN6RQESNg1MfiGNRw16vOuHtZ
fUPyOo/gvp4IIPKDKThh7LcDAP5H6G+pi3U20EygpfmEdlW3fnZIiey/IPCMitdrwnZYwH+3UJlf
x2aA3+CDsuiy8Ph/Ho5WE0f1/IJHD66HaKGDD1yPgKSZbegp+fCj/K4PCcwyqwFOyIVjrhyML7bZ
wwPr6RT+to42g14dcWIOog0Tq1ixU3+1nysairvnkfGF915wESZKDOtXyLM8akvtR4wlqKvNkTyr
wTqGKqghFX+nc9t7drpZHoLwjuBfiIgplPXYTNRIEQQGSZ+aCXFt4kIBymw2PORWF6PoBPGEmjwS
CpDen+Bx8Ot7QndLYWd/gg7CCgyU0mGEBjX4wx2JXZbjcV6u1YGQOBZNZXxXvvzDrGkZ40bmdhep
9SgxhSyAmif/YFASVuNjVRAMMO9bN5xLUNkVkMQJYIC5mDBy2PTDRbguG42iykL62DULE339ESUX
yT6SaFbZzL1xtGqq66qZNQtJ52Dh1vp9SIQAp0JjZGbicU9c+xcYHjSjgIdNWFARtNdqeOMM1ekS
CPTQDS3F3XVhfny0hgB+bnSZL0sUMTDdqXeF/fJqfX4TZX5I/TF5UdEa75/hq6irxttwkRxO7cbi
0r/wcfhLtXdIBtT8sjAPY6MYfCqMLka3DJbvceHX3x3Bd4n3RJ0S8BPWyYgBubZ2+a6bIq+fmD2z
dD//j5nsIIlUhA637c5z5isogRBCYkkFnmNcR/ufO+aVhf8mSAZ90WsSBbH+Mc1RF8TfvbS4ZZ8P
Vyyd79kbvwYcIZMpknFmXj/17akhh0lskmU9Uho56fzJ0K4afycE1WUfW2Jumcx+bU6at/rPkyHE
AGlOW7tWC9zl86z9sdwjyxZNSDhkCxbwBj4od+7zV6byx4yqnQMVCJM3hKNm1otRR47nEYOq1XTh
CpHbxsw/bnhkaLHG3LGvxh8fkY5KqAXgoZfrB869L2iOPsC8HrzdIogTZVUpwzMQ7OXjMfKKI74n
J/XgJy3hwX72CAkq0/Zqv5YWeFgxw/TUUkq7YZbzuXHTJk90/NxYsrGOsP0fumOT/IsY7WtaRhfD
7ig06jWenke+HkUaPhWFeE8YG1Ue9G+fbTFLMxWL94H0dQVTqWwIwd139nchYDGkC3vbhQ86lAMc
fH8Y77ON4z0YZo2wPm34clMjKs7cjrhSeQGLdvMIvmkzMXz0Kz/G+eNH9l9h/XgzKLq7iUalKhdL
YDOWwX8A9xxCyNpBSkWG3Qayt+9ckD0SRCVNZhzyUDfcBgqKTtPNQJVJAWYSNzBMrxKHtky36x2X
+cqi5msyE/T3fwAif9yUHZlTVVz0q+buJSHgqU9aSAgCzqs5kRpP2cYGXXZ74PSALefPeCkIhhb+
J3U6ihVd6sN3FAx9U2CDnx8mRi0Jus6GTWwbbXyBdScbn7q9x3XJmjzC9+Zn/3gJooItpRZ+8IzT
d9/uoVbzIfCIGWHDeAiZOsmMG9amgzSUvFKwDV8tc7E/0urH8UAOcCicB2Mro3Kt6ivTlb3Csyhe
4XiohCTxMxpU47wCfD5Z6++aYVCQ0givXxCIapIEgys5VoHcZWTQdX17TBJWiQH8fx4wt3FWWZen
eV7B2ZS0xqclkaIAfVHlP/R+NFEVxIinlQW/ANNGUMDdKJVW1q7WlP9g7CXxTCLvH+mwVIJVmTIW
OYXrMHVZUoRT18NG+mza8vbzAvkUh0KAt1PW/3tF20+fZACttNJZXLdolbemDUMLjxtXdaRy/+kg
q2sKwsTIJ7tH71zw07VZD0MNcAK07RboDxi7s0C2SoKnqrUEktxBx0n+bm8ukhvWO7DUVxhH1BcJ
sl5ZwO+xeTxR1Bns1IRPJ6oe+NtHbFxOFHf2OAJvRRFq2fW+cdBOTu4jhf6hTb/3hRtWhdNQilLc
erHwFGM6I4o/OfyesHqHsBhLNvmwAHBJFkylf9I4LVkds9bMkhUpfUDUL1F+kz8a/1v4og0FCLdo
qPH2pya6S7EnxT0NKTLVE3yFY6QtCs/OyAk8E75lFZOkw67/HLVnCpm9UeqM+9DzTkvRbPy3vEHk
UJF49KJgVxd+KzmjxzCPCX8MXBRHjKO55fW80/x69MQogMyWCKGaopViQrbO0jizfyga72KYpjOw
M7DpnfRxzAXw+7DS+9UaWMGGebYNDwRyXC1oBNqzN1/zecwVaBaQYjej+LhKE3mxMxU3ikd3PJNB
B97Ru7dWMY7Ug83pIgOvOSm99DZu1shb7BhDQRvj52ZppgkGBtznNzaGMnrhu0bwbH8AAy7FwVJH
gxl4ofXjDqXxtaeFIZ2MKELfjN/zAmG0Hi3SO6L4wTUSHOJwxHpG2TbubkLez7l+yoXebcRxrLiG
tnpRwiuOxuxrABS/BR7PT75lchxQ9rJP8cdujL3TPyFgb/BLeh7LWbFkTV4zgxqkUKjZPHZ4s22v
9jgO7SEQivYLd+wI8yeLk6z+FToh8VPQyfowhOIdTTVc/uXTSJ88daqzULduF9I5+O7ES1gwCjrn
8tX+GX+labjBbiiPHxo6APm0rXeuWVFfhQk2pQuxuGhRc5fpsUz21o+cr+BPoCoXyYKWSfPcbNnM
5q9+tC2ZUeaiCT+oWJtA71+Ds7mHSJ+6lGAnsZ2LKzxSEAJtU1BCt1eTvb7CPmhsweTv3eRhLyC1
wD9KbDWfZJq0OWpr2QG7Hv0pENyoL2M/J0sWr8MzXJzTWekTwvwYoXqnz1mEsw2+0SBIaPecJaXb
k1KXxfm77EKLQlMmVFLeDwJG6Vd+hykcRMkYzRJP9JZdMsIERmxuM1XgM/OyWzVoJC6MCB9V3SEH
DIp9I4FgRP6gsVFAegmwpRioZaLFd8gwdM3NYbwayPpjTN8T23yavdsxRPOG7DMW6/TbC/T3UtMI
K+Z+8cYKNoAl5HnoDdIWLLlkhzl7mgRXCN0eG04mtoY5PEwNyygqCROIHV0xVUQkcufcWckWKcz2
/uEOw3rDekW83W51xfuk9NzV0zmKk2jTlRW3f03dL71h/fJ6bL067/qRiqs/l0oq470GFSgKfZ3h
FnPUpRgPPPvsVWGvbkLJFBh1D/5gWjbQA7633wyiduLsb+eWd59xzrgt/cSQCoKndNsbIlH9edsY
+TFsteQvJUkB0XGi+/KLzT+jUjnQ07EhSU0bT06O7qW0JFoZkYiaxm0fye073qewtaVrvLq7oKYE
8wlw1WhVWuOCfmGz4xigD6gswHSg2sdAfV7uOxNfYmQV7+pz5rg5CJcjkJv7xr3zBdtpe8MEPOze
uAkQE8MyOeutzrV2U2DjcQDfCO3cD9nKwuJI+ZIaLyK8B0YHphaH3Q/ZubqPbY5D4cPN3ZQmDMV+
2pDCCRBB3ls6/WI2ig9WZhD1athcnrAMxrQ29kifn7ioOwMs+EZP0fSZIj7osfn5niZTxGOBP/Lw
Gf/uVRcWNc6P7JmVKpM1kTxrkhNHviySgDaC6S+B7oGHucEuY45Sl+pO+HJx7uYkhqyaBESZ2Hyn
xQfL0cMSj2TnrnovNkmuPUt8T2jxAG+pJktbAQMr2Y6euTXNA8Hu+SaUsxdtH/arQKPrg+lN6tub
4dXVMft56mYTCcsiYau+RMDOEboLC/wzz4C3n4s/pICrL4ro52ENKWxCwt9QsgquoEDmPewkTgV1
OPMPE+1uhO7IqwwDOj/HPtAEz+CLNgmPGnQFRyVSydlzx7lL0RXY2T8habG7L5BKltkD/pWbvp17
+30tlWINV6bg9gzvtQVeucGlpL4gApns14dhWHVCJWm1EIBj47Mka8Ok4LjssjP0qwuNQlgdV1Wu
1evIIm9HYxFJq3DVaeKfpO6pSOj0mcHWn9gzIFkCcUW8fiwHzwCKOs5D3b0b2u57E4y/Oq+2Sgc8
60M5/tbIBXUbzn+A2b0dnbU2bdo5wH5FYymMVVy/Yliv+6YKRyuTdpLUeiz6baVkVmaVwVYgOCbT
YLzMboDGcYqrtk5oHEdb3hM+qPFm9VCdrlcTJEjou7Q8DmRUWQDvPOEqgOux05v7Q3RzblvCV9Yz
KVZMG3+dGHMhaZrOjpuVT7sjZQaB8kbxfWiQ8WSHThCRHfqlh9DycNLK7rEsyFH0D56IaL6GWzrv
GdrdoDBjpi8rqu2zMY0yL3+nALV7iRXh8JnUUIltYApgMoxug12ywGa3WV92Ex4s/x0bfrKX19i0
oweYQ6u2vOhmiXSKrou11yjGGmA0cK6+2F6Jk7diENUHd6Dr2VFDTwxrVdb2otxBGIDeeIi46vF8
+QjWrkPoygmeKC2chl4XfP1bYAghFRAPfDVjMo4dCM20f+U3cmtU09lbEdrXa9zPW8jSndfz7rmu
qulLybn983Aq623e3yILmzChsYRc7PZF7IjyXHr/GRbyGGRWzGF6eMdqHqxtb/b5hBgY0gTuEQMN
Kt5EFNaIcpJW+Da+FcRX55lyujz4zjnBU7OPRnl2BUSnlaJYy+gBIScMvp4eHyP/v8i+I5D3HBu2
8iXvN/RdExVNNSUqrU4D8qFG+/k/zNXHJSdLNhI3L4qAYZ9+XXcoKZwoUaU+JK5CPNL6VKY3LuAK
0A8gYex5BPjqwYaTK+Ooj/0TYbw2oDQBIIsLPWDkulv9qdht0t8JalfZfiuT6UXKPPfFSFj7UYNZ
djp8qfotrEF7q3P7jovu4VEPFerFgyrHEzZS4/31/BjTAgjL1710iezXwTZWVUA2cePL8D79wtiA
l4XONEkQTEr3D8ddDkTDeEZM7LZpKNw7eQeDu8qu9TOCJtqf3m6wf+ObU2oTYkyQ0N7acK0PmFmU
473/PBxfgdqP6G3ktCnfcaXtPEnyi3c+VjjOcRXxqbTKJabLUXvdWfm1zK+MVWekWVUZ2juOILE8
4Uqrwd1Jp6AcTNMCbsAaiGssuCb8PcOQqKZITufLX2yW9ucjNtPp7G4Le08I6qnLLzniAHXbbf/Q
Mf0cx/QCEplSqZztACTE8j6KXAKYRmRWK/k/7HIoqdNFNIP7zTUB0buDsixNbKAeM9I4tuVnXKCj
SC7OHHVpaNEXuI58Or5+QLZr4JyvOzuVM1wvSItk+4ONL0uzYrUCguaM+J0sSKKrIQXStQ7Y5LGG
g+sZy6tQAGa6wLvJiatY+Z7In4HM/ev6FSTJNEkYKMUmxRT9pJu+iLIsAS2lAU+5p7dsQyjvZq7a
VwxXn8568Xa6ymJbndmFSyudr7aNaAPP/zVRQpRjjFb99C9sf3OUFolz7B4eWhLS9Ppf0+vQW7oC
pGVsijhJHjISUyZheno+YmRCeq/YsMECgczhvfUJ8GLf4VIDXAZyAnOJjltubJbVUEvtxVk7vUce
MCDFCAUvjT84LbEwCzibAxhxM7c85v1jWXSMDrXkl3jbtbZfxPOgYiqlomvZxfcPH2lKij6qpD7E
sjMq/HxhOaa3Zw0CGcRFInE2RMYQs2L7QfZSSNsSyvJtSzkZyt0FUxQM8kBaF+uJw3vxL6OIyyeh
RB0r6N79BjbvpYijNOoQdMymjioJGa+Cn38XLcOHUDDt/EPq4Ph+7G9GPl4sXEwSNnaWm5szY1Yc
7385fuGOJUpJZKmOYuAtGMjWOAaDrtwgCY79t2Do4tYFybAbBEiXC6XsRmcynqdGEV2CwUOO98Nf
4o4nsuIuV6COkqt/rmNkBj8wSmnBLP5KWj1YSRtHZmaig+7qD6DP9OsgcbtVa/5o9Zi8MT9IE43M
wil3sW7EW8i3lJoW/O26DySErkQCw/fWdKylfzfsayk4flCcaUoEBmCsSOzwGVwrYtdqqfAWUN86
UdeZB4tUwpHERC9NQqCbzgTnsRDFdpDLiDyDtRsdzJNrJFvGSSrIdKNgGP1nNAQgVU2FHBaPUMKZ
6G6erUuS2D1dFSYiEn1SwJgmpNNf+FAdW5nC0UPn/5NYrGTwbUTkyR0nvKF59umq/Mb+acMqCX/b
LjasK3eNOIjVg+09rcWrtajEzELoNawRDS+DNpMQud1YXMo0X8DZL5Xni30lQ4L+Whg5NtUWfrFs
GRkJkIy6MWWoAwukNZl8huq2hWYevX64g/Wkg3fZjFtN45aCdOgX+Ext7wPmufVNsQTVJIBPNg+T
4m+7GR2/bCh4HB1ZVXYAdzyNrKSUePX2wpcCEasRq/RxhuQcnCMEoLrymUriGJRZiPl42WNQ4Hxe
yZbzPCbjFATnffWPJoJUz/EPuVLWeT/y0C7ynwlBQ3ykjXgBK9wPEyWiLNnnV30BbwCuOO+esXSy
n997IAUlS1fj7ToSrTiiV0RDaqrVA2WBNkkBSH+JdpczESFrv2iIqBjBfAB6dF/DJj94ezlQCdI1
gYtc7tSaYonoH4W991buRX02y0ZByF8HpqYQXOQIkm9BkT+c1GavcdC82I/r4aaEBSuFSzXWdUQ/
x8dRSDFdFn/mSyWHJBS5biar+hMhTo/oIxOGFnkh2tvo5AeJTZiYuaLkArNTSBXVwidZyMjofF1u
49ZBX9ZfHax61YSKhKK2qJVwn+v47SXINHQQs79Xtjto1fkZ4TOSCHxn2IilOvxHi1+6eETIEX6v
fP8tjXOHk8RL0NA14EjCxH8SRz4C8ELeeCDsYJsl99UDPcR4Ym/UaR0EPm1M0LATBp1yay2Hazn8
wic8OfsUz8QhOlqfgB3dnkTRSRqpLRcqlFdtPE8y5Q23ORiccB+cnCLsw8Y24pCHAzFbHSMQwVHx
TUQ2on3h4oAfvEmzgS/JyosTxSTnMZ5PJX2A0i9rByd9Mu9QWx9+16gQ9Ln9YRIPR0F5bK3VJBgZ
UVScGCa7TlaMnbNMX0VOduRdX/Pbn/bmmJUhz994vZy5jrFcp0uLOxfeVotlL5J5St5z4SkUoLoB
DhRucWIjT8awa0/GbxGg5ZqKcaE6hRXeMMHf7KP7LhwGedVHUYoCt+D5TuC26GDbqP/u7V7PkrpA
ZMZK3P62RTWn88Gw2EalqrUJOlh/TX+pyczVR1iLkiCc5EobCEtfVuNcKyLNcgt0/EnLAuPBPxOk
fS6Pxp2brhj3Sf0VUBV7d5asm7tYu7rrV8obCUu8PTohrDM9iKz+AFshGz41HuY9k+Z915rhbfx1
cPZAFDTJg/uQKt71Osc6KKs/FH8M5uXv3m18FvwnJumY5b4VQJ3fVGuELS6OGdpNjVSwPFGJS5m6
NqGRIgPBZtI3GgYwQocYSOfk+PWjTvxzLq/72gx/bL6iDNV4ZzPUjmFqQ8s27iDuBXoNwIZqTS4L
dMedLYZjtB1w+uXDuNFN1K8lbMqZInsMPnIGw25PivYKoUdCcRs5igeyVvs2kHW1i1YWCuiWH1+I
to1HiIHDpfhhF11kXIjvcnL/eYPfsapQqYPg7UbKDKwrQ3MUIOO0PbRyrjUrolSWeaEwa2WM5hfZ
DmkBL77dTD4m47B9WnciY9700Q/V7hhxiD/RfdZwedxdvk78OWL+SmYSvdvslqgF2yDCw7ohp29W
hcHmkyRlFHzJi+uQab/bGcIJVx3KB+rI0kzz5oNJoWS92KCsUjn6sPHCKOCX8VpTkm6WG1FSndKW
UFhHaqDGCu8FuwfhS+BX+FXGfxNJktkR0ntQkipni0/p+p6Jxh2WiNswjSSOQqA2fu7oTk5ROWlq
+nNy5hjhS5Ah2qYB891dp3DlfuO1tVhk29K6n+UTMBVex9sejR635M4IMPi3gha/lcHxjJmV/l82
JJBWXMRZXfKMpYdnyxaKwrIbk9ipiViHmviPbWo95JWTFWtoGi0RO7DZu44A5cHejD51QvZ1qj/O
mv594kpMJXQCiN6dadiYp07JNxg7XQuYqZQVskhU+KFWj0mf1rr+rggLo+xQephXl4XKSRgwFNLT
1a11OyxCjNPmtsQ2/73Uxn5aTYI7YeD61fLNCK2fiGrv/wyfLpIOGOTVxJi3FVYgW5aRj6Pe6nkz
CVuhu6vYEskbnk+SI7FuPDs7ckHUums5PcBH8gBBuN74fWWQ93f1ailmVd4C+rJUVmCUgbYgjuJd
grdSqMgEIguBNMlgRunDR2GabJ0pi9CzRcEMsc5YWK/6cSSSWjEOjbJAQi8eH6pXerp988iA5zJt
2yCaa3kHIOfoKHvFxbuvBtAV4qpyD/uh6kV0SVucE3RpDkwHRZ/vrV/TJXK/Rtos9T6Y52PDylrc
E62JDFOZeW+ryUBWOREgBWG4dK9p2VYh5bvSnZ5gq8zIaWoef0ypIKLEX1LB6SFtxVZJ4Wr/3zLd
3s5OBvOG6qe9eH4PCeVYF1J6K2FNQAWZcpgWfjk/DkOqx+dcgwjJEGFFRRfkSDnvERs+BqOws7w6
SB5xbznGB+LQotOVajgPHEW4QoWAEty3XU0NL76biAyoMEXbeNvjd4jWrFpm65VS1v+mZ53lSL+L
oUEne9g3rT0pLCmctNZCdbcUsfET7CW5kN5rp60ksJYGj124+Mv9p/qcVnIh+6zRIwkwI8dWewDB
60fLzLpbsO/5ksM3jU5chAAf+5cfD36BXIkSa5SNGRvZUzlW349fyktpiJCw7jZOP6pqsHOibmMr
g4/00YedyjP/H7r1GG3fXYlnMb8rg0STwruAWmPUkUqw+brIptc0fovJKj6DJdhEzF64/TQS4KA8
DKBkRgwHiuLFPanyL8im3J7qlJZVdBMA2VLzJ0t/J4nH3vEe0AP8XyAV2z132682AYWDXTzkOs3c
/Cg/ttpybadMwbKCf51KRnS7HUpRoXDq8tontSMpQA9Id4qBotUYmo5Rbgwpwo61UnGkJQiBcePw
JZgOdkUy9wusJl7UuFYq6y8FIKL0utBStkoTc8qRDFW4z+0HYUxKw4+FSPF4R89l04M5r6KH0Ose
d/jNTFpQwc53KbWA/8hKDTSbrDsIvfU2g3Q1TX0PO04etM+F6GHum/9xAwruJv9cREOZaz713jWD
Mh4Mvc61P25EIWYIDbqUj2C+ICbZTGKLk3PYhjS6f2IvlB6aByk0SpvS6ABqhhBrTkQ3RWeWj6+Q
m6owZHllzQNYosjIsUBkfMfdmGQFVNsE25rpj21dZgN9FZgissPV5dSm3lCOAajH8OgX79K1f/zy
M6kmXOUKRaPpxcOJMHNishPdVgijxHlyw0AFPCtBrPdKftBGgp8Bng8BvqMY0ColHtBWfPOj7O9q
z2Xxf4+yLvGhSMl2PK3JKQ62fILW1DjaQt9EDD8UNiez7RJLBP42lngzMGNIc3aUnZPDbRoYryhB
iHrf8FKBlR2aJCYsZljqYafCyLJR7rzygSssSbnLWrX3f0fIH4V3lBiXFwAmvF/fy1EaPI06BKLI
J0oWGj39cgR442GsYv/Eew04aQfGWyuVJn9SAGHmEIjiYkLMSvdjsxg84Gk1H4YMQJvHyfm0WOLt
AwCmSnj4aS2gaxLAwh1FT3bRUt6Dqcg1LNFujNru7xHYYTb+m8/5d3THDu8uKnjknzXhPT1uQqYP
YeMl1TvUu0rv9qVdVfFX1l+5esRd14YKqN5IwA81ymgsYg1APevvwd+yf5Jxmxu1bjb/oJXHwCHJ
Bg+uD8LgbuANffrE8QK+h0DP+O/fLsUsiubFawvJNZgEtxev8Mqn7rCcO8j6QygDrkXKGXb1VFxC
EdhnlTQfwZIPaqFW8n0IGj/rjHYrBdbRH0UkZQvMVV/ayKmDaKfhq/9wztkCMN6OlLo+FoMdjfWa
8KcR5J7LBj9hA/zO1S3p7DXunV+C8gQVuo+3cesyKj038sUn+JDU5jkU/J1ZT47nugN3a1z+DxiT
EqWYqF4ISo2TMhClsqk7wLIpm+aWitucuwtfostNUTDkPSMfPabR9mAhvShYYp2BBI7WsUjVYiMG
0Mat0x++a1KSGlxUpxH15F+eONGTAbAvrNwPyaqP8BKQZikVnc3w+gGfdNKu1xl0QmpL8kE0029Z
w1X942PX6rh/sxeB+eYkSkavdW47P7c3UFcLgFV/7GVxgaPlKrjrl89Aems8M+3cha/Tz0Gx03Yr
ekul1WlTWbFKZmOJV2ygc/1KuyV9VDXc3k9FmTlL/KwxRWJY4dBMGBZPH5FMve0n/HBRwi9JwcCo
ZwWAjgFZ1vQ/diZ7PNePWEKmy7vpRiS6GM271Y4qR0nlmO7nYyBL3gzaLl0ps5Wnix4boOND6VLa
amRcqS1V1+mH1HKv+ZY6cfEP7syam1crdbGxVyCmQzXRLp77JpaBKOe4qE35Rp43iEc+6ITvOK7b
ilWofBLmS8s1j3R0jxR32w/pYqSLH+3kbzYC0pM7WVzRH9ZJ2YLHEV9XKuGHDELSx3UctP6jtBoo
jBjXYNntnG0m3EaLbkLNuf6vi+tZiqZsi0OoafmyzZW5A3KyKjgAWVrItBfnHVSeRx5Y7W5Paoa+
nRzhnqIZJVC6JlzVKfsyJSBj8JbEjNmRdWQZe+m1O/jZWcCWxTVDTovbUyFPURYcQ3bYdOmChLEf
acVJzG1tnugMrhSRCGgfKHBQsfqDXN8eSyLR3XUWZ+s0nG2bQFqrjEIgQHc9eGsCY8lnjrIRvLdN
tUIM3OMsrLss+pn1dmNICAxX0US0eGa8mc3UxhNmDp5eXEtdoD1GKsjQ8CqOJCReODYs/kEnC+yq
byd0Aq9PyWhcJv5cWon09UQLVgpY1lBsMuoD8wggaySmHM1cVpJkZMXHqjZ8lA3J3c/h+8Tc55QX
VAr01j7UmnlOB5GGiKxJe9/lyoip/ODo27m5xTREohdncyR6o1sbl7oCyDdZ/1nMrO336Lmcu/oL
k1iOLM9yeGbgfQMubnKPMmGclczk9RQBEZy04XhHjyolofM4btmrCDcqXwcihdaYsF+b/ugA20gB
7CB+mnFkxBGCxjEn64BMRFZRna9fmI/X7IA4na+wImZiOQ6xF9AqBLRc+B9ar8q8rHUSz0TkRa/c
/KWwkCQgmYzbPWga4ZvWjOz0CBRa38Gf0r8HMLh01Z0lcn1/zQlj9/0DahREQMrT4+y0Ii6KMm/c
CFp0rfVeTnDzbMXBy4VioKiPNZmz+Qzma8A2KNbDkHWI91DoMHK2Jdz+mVVvOOOj0ETGb02sOKor
FbA2Cmo65O+mwycgarhNVMdbeXrULR02oyscbrn/UOq0jZop7j/t5cn4TtjDQrFhznUR9Nmm7zS4
ckHNP6BA8z5kD1EdRFBYvVQjm4ASuqEyC7mviKSRnQEftvAIRlRbmMnxbZ9gy+mzOT1JrUh4tUOC
ZbXK7f4cReBdQiE/mtmPb4M2dKDLQ1F6KAisQ2Qa8iYT26LTS8fekizbxgQ2fK8z1Y9eJzVlnf+W
tFtSBH2hIYjltdJ8XIBhyvlsFI8McUL5nUlIMHHACFnRXPhtQwn2zI0dre+ahBT4HYVL5iLUWi20
cv9kvWExr7ENoQtSzukp8eia0TgEPOtrypoySf5o3j83RJaFDO7f53jrWfWh0twGZKTGpICN5PJ3
HPKJ2c2mrpqhyJMCK9FOU8UKQmuJsaznP+QhMqHDjEmV1DXtpqpdgLy2WAbWl4zO5N6BKLbd4rvm
ttspP96ABBk4pw4+J74DHpoVBnpy8/Fb9S3Jd8TN5wwU7TxEpC/hPqzzMI6O23vP4KY8TSzMDIss
s56wHFZoLjShb1RojpZvglbS3JYOU1INFNg2YgXVy0Sn8Wih8u6zWnYn2Vd4qzyRvGrL7SrbxWWE
vzeIzjOlYglKysmbrYXJQD8i6VXW4dNO2dQkcrdlfWHlp22KQOhTGTTCazvxJbpHnYaJj1PjnFzl
XN9kKfJAd4xOH6kVrOJETM4+zRk/6KORXv16Z3/4GS2NwpfO3DmW8mXAnmDWmsZBcGl5MyttNr+n
yrjrpAgDn/wbZkdMcOp742jLfQHnftxsEHq7i/m+Y6A4c335nAVV9xf8Qr8rM06I0RR0LvnMxmqm
htqCmduANY8PBycJm6cgevsQkJJ7ythtaPHnaP3rBTdODN4/RdDC0M99wf2S0f+h05nxHPJG1ri7
0PySUTxckw4RvjS9/HRLg5OKOzgMRGAXzybwGLEpk6Mvom0/ris6BZvcH0o+3j81lMlzuR3PZ03e
NU8has9PBdWbs7HVjxv8ovLY48MKdEPuAzi8D0Z6f622rO37nLHboZb8u2NRcn1qXNnFtmiuGQ8K
PFWKWvfJEArePLBgcadOVSgHRSxNHXnI8I1v+I71qX5QlQ1KEi0o+6FjFOUsJeZkCHEBAUQpc1Jn
9rbK6iCh2GcmZKbmmUCryAmW5GUg5fk57LEiamW3kzBzNAByTpwMxhhPbESdvyelwF2PRE75wAGV
bYI+EpxMnhEoR9BOXecjT3ASbmRVpUkDuuEHxCgTW0IMk95pALqH5L9BFRw6dPaKQAtSHcAci2yH
UcLTClii4rAGmsQy0NStcHhRKtzNN9mRmuBzo/CJzJixfNZqYvXazt790UD6YbonEYdCYo87qXQ3
YDnvwb+0AYqZvXH4gc4ihHaV5jgGlB/LewcCeG2pR3mVMoBFP4urcfH5Zn3JlZ+hOt9csuag3swv
Hn8CLdEU64a+u52U/291+kuvEmgrlK7y0XQBhaKTD9lClltMhnnkS5SBS+uqpoomtFhfy+ZD6NXO
sFvY4nqJseGNj6F3g1vC2kn48hMBYN+r3R4T0xYLS4lcl1HF3aTXNQEwvG5Fj4kFC5t2AbWucnw5
yUdu03GBz1MjHdGAL9YWmgSnf39BEZoHJpf00kQEsYY47Ogkf914V//e7tXFiOer1TxpIYEl5vB5
Y8fRAtFlhl22Yhk1vj5zqU3PN84Psj0Mt1GOwHpD7GWyz+DswCZv0uN6/GGa8X7gtzn1Sqi+WNdd
GKBLF9UNQNh58qCB3L7BqijBzeAT0uFkaiT1cYNZxotmyEMQdtJH8chQ2uIq1MAZgFpClCacLTYP
b4OyqUFQ7n8j4DkcuH9Q0fy5tbTGhwQ20JKOiDuSWGzsJIc82rkqtvXhrKFkYiMubZZTl/dBNKSE
2kWbMhfkoOR8iLVb0bec7jl8xUhryYmgbsc4S7pK4yagZ0ffe3n70+WfeZb6sBK+TrerExsQBMlp
56DY1hHxbp6Bz2zyVwaOezjlTKA9mJ/dffad2TuSa8Du5ocw1K50iD8Wmte0ggG4yt/IFN4UnJQb
7HOaaySTOSZ8MTyIBRqaH8AZOTyttCSf9y/Q7ABpF2V6wQLEz+OJJSuiwLUxPZJiCRVNAztQobVx
r3m4ixa6zVpoPo3HMMnRTj80ZTw8siE85DATUMENLw8DOHYzV6dBos5JVSv3Ky45VqtSLAA3b7wj
5nnKFIlt9BPXHROjgs/48eVA84LCkJefDgTn85MQb/uSwMRucgsd5uuY7/bOlJPKDuKzo514BQb1
b+UO4zEubVKeRFTvHhdxa8Cl6Llv/skhqmG7OoyLNODD7XNw/vPDVRf8QP30RFVbvI+UTCufIx9d
Cs4KKWhHVsqX0NooH6j7t0vZeXk8IC/KrE4cMYyDpoU3mAe5VB6hNNmdPYlQb8xSCIqx9ZnEHuiI
+eFipCJu3FoCrC85QPG38t5Rovk9oKGw80U8O7aty4ue+su6CJGnBK8hGhMhx/Ouzsa31NkxNh0N
c9mrd7EV7A0Gs3RwZRUw6FI5S8srOEYb6BfD2qQDR85NvH487pox4ozPes1cQIqSPj99ylKbtkzc
oaevljbkPeYLtzHjgZH85mQ30e6Oo1UTxLx/lNYThXFBxAAoxTJoDElay5cgf8TJwt/BELhDdvMW
pMmb84uhen4MF8AYpC/mmVBnrM/E14tizvjAn0FxctLvWzfvxLfaNWK+QUsAl57IeqTwunYStWpp
JbJIm8rqdvFYyFnsYvVh0JSA6cZSh93T00iX+Uv3y4O9DbCPdpl5d2+BgGUM31L8ky/R8DGPe2H/
ly5oNevNh5N2wdFJRbzWNGxUfGTE+uyf3VrzUa0yDvG+6cbC9OPza+rR2FG9eOfwjGmsK1B05Hkc
AmwX51HUDv8/M7bV6weS0tRZFhU/Pwu4iOhBQn2+LLrwwNBGwnHcqiB7Lc4MqNpaV0y8QWvvimOZ
oRgTpk253hIl9TvibQMfdcZncGaDq5S9bKFn8zDc7rg1DCEcz534QyfdHjhqaFW19WrpGRFj11Ol
mj4+6f3w0c/5oU+m6XE8KBfZMSbibCtD1bXE0eHVhenuZAoOJW+wtnYBly3opiR+moZTa7NEhy40
Q14Qv+uLuD5BUGmG7p0ngSNKNCAxDtoronK3+PQ9i3KdOoZ4916d46lUoug3yKGtHWYxlAert2b/
l4ICnSRNxBq4XLl/DDU6upRnSGM6UfKOX8PHkRqnZi70L2ezjnuYp22BSOURuPDK67IzpW8hinya
5/VhXNhWQXidIYOWlHq1g+D9xgLD8g+fwNQ2k8L0gi5VAlPjaqixDvZCth03gHGAD8b1q2JEy3RU
AcfPeoz/kXs6UddAX/irtTF+UtqZQH4SOrK7xfxoN+hZhG8hUFeiN1+7R959YXHYD9AITKP/P7L7
D8mZH9VEVSadB0h0cH5KORSd2hOcaWPpMdHqriOtZQ/sLlR5PdS8378T4hZZz0PvTl18zOiYfa8S
oMWjPhMjLSQthJy3905Q+DNG0/PechftBc6gSvlLzfk1wRIJSmewyQU6UQs7t2JpOFzOGjIxEz3u
bpcuJn3Zbd4cbkeIZxDE9oyUreOcIIMepB5uasZKORwVWNXm8gBG1pJt1NRVVFhuVA+2vHcFo3br
hhHx2qNVOV/OWTUmIrqkc7gEFgOXNjfTaMz9XHMaTzhvXNQ1yGlc/0eUOXwNYoRRPcvKeOtqlUFL
ODwDQH7h2D7rLWeTQdTGKQrdKtto1T9Bm2nxTHPwEg15kf6XwCqaHRplf9ycBNyajF3Yr/XWHzqe
tfQ1sz75hkjw/CgPThh86Za5lWmOI+n89B78CjPZsTFM5SOlnN93Tog3LvRwKqjdIdZwWIJJEkmq
SXwrLqL5ZM/+TgCF1nQb/oFMIBO9hkJVS/OD2muI7lfi9FRS9KR5IWEbjIZsaPZz9vp/YlInXTV7
hjRadEADN6l2ZusIIZ3Mji6IoSwmFKtwCqTUZJTGz5bFccK+Yn92IsDDzfvstwuha/aJKSmB2DoV
ylhVVRghsQGKU8pdJtIGeYD6EFAYTAklK7zDRyA3h1QkXP3l4JdDVmV5h8VekGWWbZ1BwQBsEi24
DB88xCZXMX4mRhzIuk5gzwdJIVr9X0UwLTzCOpNvOMtFQMKItMG+ELsCiLlXL/lZhwm8lVnGsUW+
+Vf+HoP9Xov0mZ+g2rbdkN1dYHWaxdlBNXLYzSQrn4FWv7iFUj4nZHS1DSQAv+RZAqOqKyuA+WAo
loB8hfaVai0/tUmMb1P3S3Ec/imjgkgBIZW7TXrQrXoGQBjMXrib3RCizKMlxpDnyAyPttr+hkX6
QRPDQA8kV2mC8xOgvysu9iqi8a/isrOYybE04LhQhZnT+i8vqf82INqJBASAvKXkw8ZAPz6Tuz7Z
8x2RBg/+4QfsjGmxc+DdX+jpCZZC4ywL6mvr9roI4ljTkWUvGoPxlTwgQTEuGSBePoQHxQfW4GAG
EeNNNy5fztmYxljipT7oejNCb8DielDW7cpfqDSkJ5VNt+GMvEpigf0GU5YvYePtfrK/NTQrIclG
Dqu2k017W2Qz6VwnhHauqOEP4e9ram0BAg7vhpgFib5M+61IeM7p3x2yuOYYoP7oeZOzeBBmsAyc
ALg/LO231Iw8eC/bghkIcH6fijNY1KDINhTQbHFRwLnRaeZeWAGn/psTlLJAj4311NSY8rw1Olez
PyMQ4zewPYOo7enlA8clz3495peN+WVKeQyeplrjmrfryIz92nm09kU7DoShQ+0TFbCiIbz4a9cs
C5sJ+kRwDYp/2XuEjoCBFrRTztn/WoRcjD4H1Y25CGiaOh5Elefslo5jIPPwsHELC28OWYtTgXmB
OC9sTWXjuVSQqqNP6DmYu6j2gdFLAurXsXf1QfmL/P5HH7CJdxh4e5u9XHHwIujVTFysZOM17Ly2
wU1ANwIo+bB2a2k7Jn7UREV9DQpc/ejFyIbT9yOh2F3SgOj25Q4FQRYTWP0RqXXtYIkJeLSnuEbG
8SRD6Zw8hqzZu4Bzt1o3MZd6kRZ1Zysdu53E+5xCpQlzEAgnHSirRmmjdRxfheOlUwBpELi05T+D
LJPpNRHTgERi4c78S5PXVtQEIpsKOJ0f/bS8hkITKq2IPi+cLQdTrtesTIHEkMbwGPpgieKBWZn0
Hs5REWZncatm9ir8PqRlKOxTW4ErZuKB7yJ0iUPdoiADh2KtTIPEKMCdZEfpmuM41ifEfUA79+yP
MDIHso6GH/gGI8qkA9HrLHcHN1iQdjF8lahy5QVNWvHBzNi7u7wN46gs9nfUI/qtU4BwXiRyBIta
LJvS0nHPJ5sqyfjUi89JRYmoOt2s+i4NROJ8MxFflhyxwjXP5xa/f7yGg4zz8gz2aJjWR0hQT1Tc
8Jh2rq870Ln1rPXzXH1s259ddOzb+rrRWgyzlDMbk/0dLmlQWQzIvqudq310+hKuW2+duUTM4uRH
26JcMc2ASvCMLRd66TqrRxB5uNZ+htT5mlgoeAr4OfuYEBor1D/uK3obwNcQrhc/qBnTD/tRHU86
K1HHDOd+Kt+vIvNDqZfQDfz3/I6tM3Od2vW3SlLJk5/ZcMgIoI0dQWQVqZLznH1/VWh6nXDNHJbK
P7hdxQMdzaIykHqZMXSlIFTBLauvF9HlzDcBerZHyphljXGeniLxvrXYMZxDNjq5JafB00qNBR/7
qMFnpJ7wV74CDHlzi+9GkKzwqp+F3AX2kAgoEzM4z4tv87/xHxgrNUdFBbN65jwEjk6Hr0kIAU3+
ljbeXRapSfhNRUerZS+pIJdGC30B8nvNSrymJUO0yk8B3h8YwatQtxm8iHXPQRbIFJGCPJC/cfIK
U5u6LkfYLo1j2uE0koV8pI45LJcxkBOskUzveKPfeg/Cvi39CuaTpKgnvG1qtEW1/1FepJoyCrHZ
UBZEBTpn6btv/I/p/SkTof4PLDsroWjehVtBBjgKoW/5P56EYpNaiMKMIE/izZ1tbJ+lDo3ZGFBh
gSpHrHzUz1IX3VU4EH+rRxwo5SeEFJDWONEImRl4isSpt4/xdBt0GOgCsEjT4gWIowLZvxKayaAe
mlLM4RF01c3ADFz0nHQi6bJO7f3eXU97UTj47Tc8ilU4QSjpnlCjHx3m2Q86atZRwTX59Ohk5lXQ
G2JKLk84ZMINfsUI+74cn1lEgOCvz8GlnIy9z1P9VzLc8Bmqy3b/Fdd2YN4JiwVtThhLQK9b7f+w
aOzT/O7UUDmbx0obWyKQBKWh1rQyGsdIaEFP+3jfa/rOrEeh+E7LkxavxD0Wwv+LRf0TE/JFfFLN
iCSDiC9fzOom3PznE0qZRyWLTd6BdnUOWQ6gn9tz37ekiOS3eDJJcdlbVu5Pr6xhN3irsRZbLbld
z8mBkiChNy+ebT17JJngDQ21cihLZh81z1X5rxh4yaf+T0xWF3AP8FB/e0ykwM+JKQIHP7SzynoO
r0EvKM632rPm888cc9T9Ab2gZxY778e7XyWf3RG4GPzPGViu1bJjNbRRaSoXvYsbIYFI4rmWgmjJ
MlWf3GkpofyRrw8/vdA3vO5Lb2aVJvVlz3/nAF6Ry3pnQbJEUPfRoX2UBuJLU07Mv/7b8n1PBEYS
vTovLV94F39rhVffzy79f6pRdTUSpegSyeePMMTb5qkYVDyJXZoYL3nLYFXkmKy69pKLfldMjQkn
CdzoFTr1jlz/20RMZi6+QnzcprJqt/kJjldL/mzoirCHrbziczKVxL+JAJwIco/sbRptSnTTHjGV
sinsglPjb89uNxOIuEbcn1pGd+Bet2zl3GmFxreK+7pENQEk13nMEEes1kwz3VF/vtrKLKQwpUaW
4B9CD/4t+1V3332By8n2Y6TiuiX/Qfc/6qWBsCz+2DjZ0lnl41Imn7CVp36ynQDDiaQkuTOKJtSQ
o8TsgX6yZj+cHGm4Pd3l+YIORlEVN43Hqadae4Tv9VDENN5yBUaHvSZfi+FfpF+G69t7Z98bnK9O
uGCKwKP1/18DMCNivuJWdNHl+LMv7NtSXua35RsLTfaEmXjdqfbOBB4G9PmBoorIVNmf2Tsdf0kc
Fws8i91pDAvIqrTfuh/XZrSAfPzuoDKrIxUOt6n+8moMYomFsbY6RZJtH9d9GWyk/yx5cSS8DDzo
FJJEx+hrNswqQaadh3nZEuDwx58TqHpSugGztFRK4QFiOlvD2/9rA6f2p8XOconYHR+WtBZ/veG1
nO5GhbCTVlzAAZo52es1RYls71QLm/Hew+3JeuRwFYSb05TWFWy1IQX7rsvr1Yb1RUnpuyyWz1ei
kflW2H1uy+AvUtGQ/GUh1i8PcptULCB2ozQuCWV+Y3Tk9x5teUwgCPjo7g+QAhk+f6fgGmLOEei7
DtF9YGaPsKsuxZObpLecHSo2glYBgRQsEOf/2QmSPfy1iAaOd/bU2PIoOhE6res1HtDNKtdQ4YKF
zlNAemBFour2ix/eV1yfOFdIHlUPUfznKo2PQG72DsWfsLvtDAEwUpfI5ogXny2NHcfQXjk8kZOU
HTiR3F44j/gPMSsR8Wo6UaseURFc8R2JOP1ogH3suxWENY2Juto2D/OiStFD8CrryfOJGGrhFg9X
UHETsa+ZkMRWbD88QYaApGZZR5Vnb/A1Lcbpb5xKqs2zBWlnGpadsjUZbdIOjit43n7Lv0cqcxcD
R4ABom/kfAFynzSbNqg+pSdD/4fCDWZD6ruAkz2/ZqpTJ9fD3PBpAwD1QDJccOo42k2y8trKB4aI
ppXhBk4L/aqJraNJqf9a98cnPq7vyQCZyqyJaRSrI72v+3kQK76TL1zJlOv9oElnqHT5kLhgz6d7
SDmQsTqR421r/ZzPRMtgHZs1y3HOCsPqQ81xT5p5yXMPuHcjFbr5ORnMOXWkF8fQf8ZlJodaUw/8
guM28T8XS2YXJOO5WSBkSiwxuUcjP/tCbD8ULMFnVgExOge/ol+BPSlLoJVUaY9bboB+DWzbZhMH
cuYAyvxxMoTRqjvnbHuvVb1fbLEFqOhelf6tzd5pdyeiEB1x7VxsNlumQcCdEQ50VdJT51pU+Sb+
DGB1DbLP/evampg4OsyFXQSQHI+JSg+NumSAMPZj0PWpTJ14WScFIWsUSa2ASKxZbXp1WOFYPHAE
5DbewE+676sZVuBPJoDts8ymz8cSWgRSZrOxngWxGXqlNDnrXcaUU+23SOZ4epkMnWQKK+u2ImLm
BdbbasU3u7J6msG3Tbl/NRdOwmadzgRYtIVque8CoAojRTffE741RRcU2ZgEzjYPcjESIQIYZFLd
lNpgiUtwBHJdrHotCEMg2xkAxkeDD2qqwRhgxVcgWLb4F0mEY2uGJsz8rAZl/4+FqI0TxLO7gtAt
NwxcOiA8PfEftNJRl3kwW99ZoL2IF7XN/Tn3WZAE4yTbvZKZszSZ1wUSnt8peyLFBEgwpIpoO01Z
wOWmfFhgsBoVtmch8xKtRjo+FQb6SDzvPArt2IEPbyHDChDVo7IWa5PapkA+hZB756oZ/ugBaZX1
L3reXpTuABBsoCbVmnUQisSd3CuvP+SCNNwJUJN/VIA3nVPBMYMUoi2h+C3QvScjzDrgwLM/7dVa
vyO4ByGaEbU8/Oxukh5tIFCfI3TNoyyYLglmKcESmhPZF0rUiiv+OXFGYYBmIN9ABs4DUIgyLpdM
JHTScXaSZHHh+jdZPPcJWZx/2+bXNIrC7p9ooJM3tbZ06T+TYQ3ZgFpgazE5z7pOTpwUwbKSsl4B
DOLqnNkPzCrDv6xvDnU63ar/pau6f5DtJglKetGV47LMckAryNfN3JYpyKpr+Nm+DenS1LJNco5C
id+zlDlF/C5KnizCee0ndqQo+Kun6amkt+FzZ/goG0bQVP4CYADxIjynC7J7EJqEegqZIGj/K8rU
RFJIf8m8AiLfPK2pECEwHSTZ+MqjtI6SpSlZgBYOHMnS2uQY9+/4ZTlChzI90Hthyh9TogYxSjvd
CPq19mIqTIWUp9X0USvTcLzH+87IFh/H9W/hUeUbRcERA5/CbiHyRgRiShMbAPmS1tER+QUabRTg
UrzpyDEZxl2Rv6KUEiVnTBwx3jWs/dq16wqXAVWw8dh/qP//+VXfVJFsFWfxdUPXIavhqG1K69TZ
lX2jPF9plZMTn9kcvd55Munk2jSWhnM0Lg1P6kQHpHX9TSWakuTLODOXsqTPgWRga9z74iFunYnV
CYR6IvGjD2K+dxsCAr6Crvv+rbiS0Z+ozTEMTHk3m5ZuVUI5/jUYwHD9z7b1ILTHbHuWMK7DDzJp
pw2rO3fFxOkWENpohE3SUfFkJcBRbW7MrDBjWPTyBymG4gnoX9S6BSO8ajE7DqPb04OCjqHBcbb2
5a4YWTZ+aHrIoCc7MoCrCkKiTpbkeZqKtbvz96HOj+BVqEinxgoXx6kTo8Y7gpG1K4QMICbpBSFU
HetOmA3S1MDTT9l1zeJL/LxnQdpHO6Y8+gR+IHsKx8LpDUggiD7rBl/OYOvFYHvW+/K5c7oPNDeR
4a2CVYn094JaWPmfgWQ4fR+WIz9kUMDSTRNW8r2XeYZdIeHmKeKYHJv8uA0q4AGqtD6V2dUwuIpV
lIo3PwcW1NIwKsi8hE1xD77fSnoH2rOGSUR6aoaw+3xH4FrzayrvW3mGZT+Jc5X7zJavpbMdFar8
0y1p1CvA7fc9EVHJvOYqTw0b/SypxdpOudd9u0revzVvJ7ng0iZi0CfYOw2Y3qw11a9IflwTX2Ov
LbA0GSZQBP/d5sn69PeM+pN4M2mXvlaPVT9qH3b+FhBur4ZB6pcgyWNPCQpfK8YwH0EArooWTFpE
0k8gb4T705iO4LfnYvOv0CRbHhVMUQIjewawlZ2GMSee4Jm29NGEk7XhmUXcIVBnZmCzPW7+abkq
I3q1H8bBsYNbqFzP7q5fP5tJdEBYKV6M5NVycffylFqr6wzb6HrnAjOJPo/b2FwiqvxmkZUOBs6+
QndfHK82SI5BZhPC2+oo+p9f4V1Y9AMR2esYQtDM3LzLk9OQbGyajHNVk1BQRXUMU+NRmkqw6dcQ
rpxd0YyDCXhBJOpBCq6PXI5Fs+izVmYs3+aCVzFG/ZBiV14W8LnkPeeRB4fmlg4thDUm2W7DmF3i
HWiXceAE3GWNReGZyh0i9geo33GEGghN10OBsLB90ooBx4nr6AzhypUC39mRbC/IR91S9+I4QLSC
/dVOwW6B9ttFd/qJruSQTGaC31P+1PcEOS7RXqkba9NerufltuUUgSjVl8uWzM3YSKzBnrmD7hkQ
B180+s+EF6dgjlvdepCRPCLcdPWpjlSfBdFSqFj1IdadoEGDvJa0Wq99K07ebfQkAauJ4wSQHfCo
bGeXzHayOuefx2y0CX97huOEJN5OquV/cJ7Zbazh7JrdW9KDGyGso/ILI0zl9ksNCFvJdAu6O0Lr
+Y9FOAK6KfZBe01GoXpk8lpurD1dq2JbQTzLmuvGIXVTFVlsWny5NKxzVIKZ59T+28EUJnP6tIgT
SCP/PH345YzRw0mpaUQUu0NauOP761IMq+aQr0LIKAxBCfohnFIOrXMiY9c4mCpWnHEyO6XX1KtP
9vUaook/43mZGhT4+xhTuK41vY9I9GpM6THV54kaJHBpVkDYBHM9LIWGJX/xdRpRzZtSIhTcFSva
iPo281ccRwMk/q3B4qW0RscvO7QhltRa7l2T1x9p+lJPP4HGyH4TtKSahSueylWdQWXsfzgDPDKk
L9epn5tqZIi1UWNf+lspBInRFDjVu9o4jb1qzcCjLEYJ2gK3u2UHORCOpMN0eTm1cGC9jo5ty9jn
hE1+3nMB/O7wTdplYR5wu9bRPRqemDscQnNxubidCdt45SwSqOUA+eJkeBfspDISJqyu94Gzq8Lk
kASqV+i4asOELCF8LZtr7teDe5lBYr1y+GEJhYSzuYR5sBKwUp5/JPxkSM+dyKfM/HvxYUsyJYKf
VvWZm3lLgwX9UDe0qhJkxyflR/R9JbmmYm/9HJNoSOsAcMk+pW8+eGlZaiy+NHexitfbt3O3XmHu
U2eEX5dtPdS+MfcUuTlJgy0suDfm1ATj1kDwErm9+wsdvrPy52f3WoPZMFq+C+/4Cw1Tv1kbUTbz
7wskasbet8o62Xp7iMdFvLnRu2QNxzlHts/sc3KuxeDXdW+kxUsr7ka4z2CjtGuZK0nMtaLJXtpI
Wj6871ehk5SEnqmRbgtOk8s8SGLsmpe1a6ukmmLnkPz7dJ8zGFyoXc1dfvZOldUSvzdrfMZT8L9s
7nVKFuG1JyYvV+bkX5/eZiDYj/V8Wug/SAFiXllpub49nR6KMkUrReUSJlbB2oETroF9soTtVveP
H9GcR20X+1pP2b/7ZnodNBH6uZLD8izsyKBRFsXPrXCyWC51kyKuTFXez9qLanXuDut8AdDPcvjm
JuuRz3y1yFTsYmnO3AVx09j5SE2LqdnrOkZdmdy6UBMzJR/zhM2H1G3Fsdi2WSetz5KJVr5VpAMx
r425S8LE5gpclxVCGM19nB1Ip/FCvfUAIQF+4aM5mFZq+3FaXUt2WWxjmHrSqAdhB/rpyTj9FQql
2djt/R9nYioExWpBSo3DCLramP/CUveKuC6FKlm58gsZmuEAiKpKsgYoEYs0wHMrk/5LgqdmQvp8
V4kO3OmGlTDXDlR5tThTSloPyBlHT12sCLPrbWn7CWUNBzQx6DQxTsRcbFoI2aLCI2qMzkQQqmaN
PiPjBnRXBbJ8mkL75Slgj1NnVHWcNs8VsA51mdSwhIg8qDFZvob8CqsJ0ZPmobkX51s2X2k5O2yr
QZ083rJVeIfrR35JVrvGlElK9x4GpsAf6dqLmG5fAHw2UA8/OErnSaXRdDUbavN1LWPM9/k2Z7JK
S9j95p1E8dHdMZCLP/hbbETAVCTD5QV8Awai1bjSQQaplckytqNhTivrsdEUFhoXEL7JpXdPPboy
mGinL9toT7/vWyFskFSFKlUD2Yt79ima2ijNERjd1DFwnB5aD+AM1Zfxi5jHKxZtQ15cDmnuyjio
tW8glX0oSiksQ1R1en49MkfcZC5r/pcEeQ3jU6LVii+dIYtmAPbLii+uLkO9ZkUgiYcr0P6J68GS
83xgIunixHu17xRJM1eifLpJnEBpbOstpUn1Ba/FTlKoT4q/vYQPXlFV+krc7uZqoXRB63ZmSnBq
kCOrkG+nFIUWmA3oY7p/1Qcc8Gn8HTfHYXcxFR8fxcIJNWfdIJ5OYn7R69g2nTaqeeEPziI7wfmc
gHbeDc/Ro9T7dKyEMmtC5vBxCbNOqTf6/efWv5o3MTRmtSKrgie/bYOXDtokIciy/qEPs9o2kYye
5i/8aXWNl/yH6LpPyss0z7Sn6FYsAPRM9/HfYR2l8vbyFneg2cXo2w/1duuqjcrXZSrgxEa5ol4G
KeBq8z4auN7xscj2pYb0XYz9uMjnwGymM5bJmdYlsvYib8FgOnj/Qzx/19nTF9hG49HrfE27BeRU
J/0mGIV9Hdlb0kuy160XdCQeB3ZBbVrNErQlTuiusgv0SeX3GEW03Ij5/XCiTl5qZQRNb6as0OPl
esGOkwF4f7pRjHGILtzN+MeoQfhCOA4Fg+nHWWvCmpTzshvs5MK0SihpqpuXn19WET4M3cjrukfp
dtmQeiBQTVYvHVNtJLg0kQJX1Tu1obGIfFPTGhxJ7mt4I8ssa1VjT9ESkDAAJceh6pOY5XsmSA+n
ixZmiYcC5qGv8gctV8iXTmRt/gMrOMg+KqE4o5VAoOGoerzMyMLi41F2NAEtSAbrR0jAVEvAhd73
+0nWk8uBAwmI8Hjw/KAAQpUQ3fY2JunsGQw7BBrYS0215KqdTdZt4FbB07eUayOb1s+zOsEpw193
Fj7zkdNwQ2HVm8dPYh/ZsGWUPc/nfJWUpCWhuppbix/GnVReav1wiXb0HRvV/+T2Q5fFO9FHTebC
WSTmeFyEAHiRhaFXuVkFv5pCDID+YE9oxtSI+RsHNzYfQcHQGnaaen85m9ikSXGPKvYSpM0PCcTU
700JSWMe9CP/61PNfgw2j1yA/0TiiDKoFbKnQmQJtEP8hLg8+uyXMtN3qO5v7v/A3S0JnMysTr5H
Ec6twI23aWO5IaTF8JAo2a830yVvGy7nQrhKmEbnt9nr/OOZfSBffMIUt4s1OV+rFJhfBRrvtyj7
koaGnmgC7tKhcXiHm0jCJjGbfj3CdEX5+Bw5HoKFepWMLrqCnp9SW3fnZgUolrBPiiAXdiqOxPkQ
etXWWZON0rNIJKhy77yN3vgaGyAINlBt6I5VlU03hHGtoFKakVgWdWr1cc3avZY2fDnv3Ib5Sm/B
4qPZZmc8oBK8aZlDx1+Oa3t1Gkx+OJUSzOYOg7t6eYgPZlwgVedxtRcpFD/RgrtmMuxUhvRRJQAe
AXAw98iPKRdILenqfxXsYnD9ypFZTuv9yedRxNDlSGXVfhVvHFJ7BGxgSV+gzuvz8Z4bj8JzVcp+
8OGizIyTYTet9h0jO8i6m6FxodNUcH6ARPmp6x2Ly/rt4baGpTth7jFrG4HOlspUp7oCi+RR/bPV
N+6H0q5BXwte2fnj7AHIjkHQtn6BDotWkXHesOV+RuP5zzR0wPpq2xyvYU0n6CV2I92To6k/gHRa
j84woy/K+1RiVmnlolDq7YJXRrX5oduywwj+toSwa/N7Nm5XhKgr2zRo4/s0cZNTyt35QG2xrgWY
A44R89E1hqJm2x3uRfvhJDGBVToIn1H3juYAxI+BERRwyml77hWl51rRbyh9m006IPVGtg/UE6E0
Szxzqg+4bxUEHMUcmhmO97VMK+A14qNNVbxQpF2U/Zr83FF0Jl0hLtj4O4IlI8Rx042LixLXtprY
HKF098cMST2TmG+xLvF9uCLhMChK23Da92ZZGAl1Q3E5I4p/eH2cYhL1RALmFCuRi19f2D8RE7zg
4YBJIGvueiiRNp9/Bn+OacjGOAw6G5NPOyFan4t9k1EDLNxa7oJBoBQ1cCr7ffFKMwsik1YvQwwY
UC8AEX48/TVfHaopPiPaGkYJGHM0Nc+AAChBrppA/c0IcIR22iXVzCbqVvQIPjZJztGgi3DvuSJF
nkzj0VLGMtm0r5T7prlhNtRV+LyScUaDvcob+wYapAqCDvC8+bB1Jc/V9Ay4zxGKu31duWgytb+o
E9oiOZGcVdAia5g8OJLiSgwexMiZK+A1nCquh6K6Afigss2exTkprI5424+L4ifdAUZPDnkWec2l
3hcNC9pLgGmGcrJai+jC+RmJZ3A6pLqM8hf/zzE/lUm09OxuajsZbzehiBuW449Czi3unpSsvqr7
/k2VrsqbEyYAVenHrLZZ75V3Dy4TZadd/0HRVd8vDXtSv/Pa+wYSuTwE91SwFUgTddRkI3wjZcG7
Q7uYiO2VucLSN+xeYfeZeyBFppAoOpS9ctqLuxmXFkAOw+Pmpw2CzSOYgTgSd0HcZl82yM32XnQ3
nkmRojwWPWWOMcQNoTXWiCrr/LcRrioMKmSIE3LnEKoDlnb8fFItD7c+TZU3zwfWiUK8mqak9bQl
nMwegWu6s0Kb+v5tV4pdNa5egy5kLx9U0yzLYIVZz3zEtK44PG5Apx564fiBxBOhxaGQWV7C3yd6
JamStOaeUo+5yzt66mQ5mOppdh9bJYRON6KvmYfdPWNtUwUpJ/+QiuWPzQKk9cF0R1dqqV/ZIQNy
MYXguN7kx6FwbVSNjU5rC12Y536dbzWz4N7zka7+F/u0MJwoemxffUJoedhS5Zqh49Ao6K3ggrKI
52HaAKXtMixlAJzKBvLanD0uMasb9sMfQ6uXWcP1rU67puPiJD/6r3690CgK83FHljIatbFkKLg0
XremjwaASOUJRFsxJZTPaIa/RH714FQbGNNybMm1sfst7BqDUpUK/hySEjXnbQXRq5S9O9pAPn7+
YykCO0Ob8/36QsiigNVW60Fyz8o5py884X1Xr4230zECBchOCCU/Scuz5spJfaTxwzyU+kkFd3CX
dXtEO73UgarGUFVR8aQZz9LGP9SsfFlC7Ygf/BLvPQB43gLe2qJX7Kj5eWQNHpEuE5/mXT0EBgBC
1B9T140k2sdzvhOANwg922foGRkjDg7YVFTUiFfylQP/6vvmERZipmoRRHVSUgifPisf9WBEEGf0
1t04KbrqPDY03ORbydw18+hSiJRyuDKXJ+FSFMn+AHmQG3dkkc+jiNI+F2Xx0SDCXsq7hYG5pxgi
OOf4R+nE0i/nNl8Am7OGQlxtTqj8aqyMsbCcct/E/Uo95BflojGVpiUYlHqff44W9UaiaSvW+XzM
sjn2adbz/0cTSyKrwPpdnDF8JoDHeShS/sdawjFLguBtbwE7R/CY1Oup9/+sZCc0HfdrN0Gpp5Bs
D+L+HYEr82380FHANL2GeachS7XOiM8KPIc289WyFevvhKIkMHWe4nH6OfmRyiyYvWRL2apCbw0D
jDj4vRjY5+sqBfu+kjcmix4bKwa/PRmUxIhN8FmIrNBkY39R1y3QGm8T/cZCJLJlXdVDIx9874Ox
gcpwY+YeZYnV9MC0i6/urpjahMxZ5dY2iEPwp28wQbBoUw9pWh84Rssuyp/gGCAmMLu2XUXt85Zf
evcX5myeT2IlYWLp8KLwnB/EvoXSqwmZvWYoBOSFliAZKHOo+19jof3R4A8tQBZE2A5mVIiPaJuZ
Oi9hsliwol2U/7Br7P0eSTiDpwX+lTsnSPgZBPvFRnSlh7ldzhwZ5dQWVeOr/KXcjiaenrdJzozf
K6a+2JXC9QPmWMzu3gNCrELEh7rmyqUoVoNZTMpX8p74QvC0rMxJHEQPq5X5/fq/CFg2Es3f/keK
SEsrMhJes/LzN+ISWjjscrxVNEn4dJeh8oOVGObS4EA1yd8zH8/9E0FQr61A8p61mdqsS/CKRpJQ
5sQBjsXfrCuZPsEzrbCJl+l9mmkIpgBNmLYsPSP+3c0i4yrZyHP6dBWSMH94qqMk+L5FMkasnXiT
1CfZB+r4ZkkkQ9MkJk6rSi+VSUNMySoqXhFn+LNcd7BO5o4MbpK30q350pJioFrpZKu0/xA9v3p2
a3xnsm6FKKa9qgens2BhimgYDaREkZHX6hNholUK3lWYh10haXbbyerT15P4r6LY8ndaeOmMKEzG
XPPQW+s24o5ZzSdfoCnJfUXQj53KUuaXzBb/IPBi3PDFoNcGhzkA/3mC4kp7Dm81c6oBrfpNN+vn
IU/6+66AGiVg9/n2vh3VJNHqS3LXOq2d5K/Fpzap7YK2/dzAddY4ByAvp9W3TCgWgBK4/inthMns
NlNszlheEkBsrfOqP0Kh22qs/7TUMU6DiRQ4IgTKs0B4W/QMsD5DXtqZR78Gk1ihJxDUuxO06IVQ
umcD3HY3/sa+pfHhxHQYsfVsPWagBhBHTwyNNMPw2KNqJqmLfQ+cZXguNsAEgWfmhdIzT2xnFCQ6
wkTG3lT7yREEKDp1aS15YIuQHy9y5oHMXqnbOIn+WoPxP/+nE94kZDY/UdAWedBNbuhT0ceTibsz
3SxWwUp5zhwngBxGdDlaC4t6L59cjvC30xfqlVcOruQGq1faWY6n1RduZFSw1CiDZ9by7cTTjkSM
5pLDmw+/CExGOX1znBy4d8gAC1Lhh/+MABIUYHNr39i9S/CSAUTa7seWHVlHWt/5xrmRfIhK/cAs
1Ea8tFrtfBqdi0c9R7zKNg3PMzA/NPyk9EV6ijTS6OgbZus7STs2xVEtpl1UrGPlKhWqPWQLy53T
BRKPgRL0JlOQQYZY1EhMyfkZGD33A0HiQ7UCO6czhqVsJ6O5QN9dBFLLrzvM9CQgBDJoniQ8dUSw
eJZRn5pb2miUhcrCPP33XizFgCrwBVjlwJMNeTEhVA94TRhhpA9ogV4Lku5O0YDoZfIxb5jSHFd/
p3YqN+xcF81f12c/e7jvxYxkQ0elLLTyVmvK/3nlQHiTmkjOFJqfAqKeh3AdfwMaMpfwozhSUl9U
9IftiVituwjuzyeqpndd3ITnAd54VFsnj1F4bRsoTGbQV9Qi1n07M9u04tXchLZlymJDjJM+/Yae
gpX5MOuppQnUD2BX1lFHBSrocBuubB/zY+7C0Lr+BfBgTeywLpKL74fZq3qaBirvyO4dsuK2vL/z
p7z2aEXbL/qGt3RuNaIQgwTDBAolMLtUf1f6SMaFJaC00eYnE43Ag8PzeY9NhrHEqcTIJAr2uHq1
osd/Rgirg7NJ8Izfkrj2F/eALpWuyTBciFWDQKVzxp0WCy9jVPVXSZpzjHwzSfCAZz9HNjSx5esu
VpnhBt3GuBqkvBGx+1kQsG34pSotKk2ni6GU+CPamnfTXYriOT6Oq3SOYW0FL9SzvqqE19ViUV3M
V7DZC8OGriee7aaIZCWv9iz/GnjqssCV7T77qdxf/lcQ5mZ5GxNzCDzcP5d9Yt6YqkTIbpitR+DZ
bj7AlGeIar0OKTiEPpXwhWs3I+6KTi2U9TSMhVo1qFT+j2cn5/xIuXS1ipW0JUfQRCAMwImoaqc7
YsqLniqOFwfD38L5dN0CLSHw1RAVtdFAUOGD0mnSly7tlHlyWQD64fDl+ge15MRbXO4ib4Cz5KXA
L/EUcmW+c9P7q5C1XxuAl6OoPi8FEii6o/trrbg/scWv4Idlz1BSruOQIys4ScTeqACa+YOLpTjS
BUeWjNYXjY7Td2A/vnfXDAHFtvwV4rqa+7E0ulf6yxuqYjoIQpsuhak3yC4yoUSTMV4Zw2DgcW4i
q4099N9gjxzfI3/r8vWeOB25/hv6LREtOAUD7Xh3xCGsW5xo9psM/yLougR+hCKqe2mj5uS6vX7h
Gml3wSPN1FP5EeAGF+9LP3JmB6VmG8Hm8FzSTho8sVnUq9Rx0gTTLkZfw03qQSuD+xPbEHBCGU2O
EjBWkTQxVt5Htta/HxtDDzOnkK2tEu/At6fOcHd8hnKBSAy7raGFwBfeNze7sEvCNdid3GEhn/Yj
EBHqjEpp61cbbEcwLmhig7Xh2eVQv4nFVfdV4VKEJTVg6tG4Xa6BYMEuWfv7Q8b4DabnFoPpFiUL
wC2b31bZOSdkV77kWngXo58/cyEvjPgbIr4pBwhS3O5ToZFB9/X1C8N2QjRKkGdf1irDi+1C2CZb
pwuhUCtfCZYQ6yb0u9JEsrpTN7s8w227if9RAEaEgDX/EBSDqzfWlORW4rvFO/ziH1f0qA1K0XVk
698kii6M4R8Nvc7qL0If1WRkl/75glqN3Adi/cOdyc+vxJlQTi/umgQvSNLpbMYNb8s4Ff1FSezT
YqoxuID3oxUe6textOVcq4DWpF3IRVp60ezjV9wNP/SDx3TLsyW6NKug/QxeRTTQoTm0XWMjF3wJ
9qGVH5nmeE39a7VWS+QaelApTeGAmoaQVZ6h0gYmsQCRUnG6bExsEv7pP/pRN+yUjCufVSS7CFFW
wJFKCWc2m60l29P7gU4OhFI5oJp6LJNjvGqItWeMrnyXiuvWe8FDGtH1NxERqYegHwvTk8J7rzF9
4ZlDufxohkYuLbCn2hywSqHPRSNOUXzldvJ8JwvDz5oJC2Fd4g3GDw7vLW8SOTAXOeAFGFleazGs
d+VOYf+CeXA9wmZ1u7UiVQrqOysrxqEwsn1bjFgimJa/qqixqW8VvoIqQQ16+oI3FpE8sJLlqUqf
+1bHnwuB3lMaXMLbk+LX1NQLtz7+AdKF7ysAO58KTjPOc69YloLOno+quN6Hqoylks8LRArld62L
PD9OUrl8khm6Jr7gTblP+tQ1g12Su66OPQkUnsYZ4ACr8tWiEPuWIAGQmkQHsOxf7c3O7AJERa0u
XGoB/AJ9rDp6iwzIA9p78JvxOWFGPxz75s9wsIJLn46zrCYD5kObnmnCkIWMhvuHXHPBVCHIxIrl
nszBzWf+vw9IUCQuSRUELvYsg8G88o7bqai1oBP7jsoOsB77szajQ9b8ynzYneVFBwtJG7/WiNFA
BKoYOII2PI7rinxQEDLGcozQN3QiU7tAGYOMqmFIY3RIa8QkbsIY/reqJEdBkBmg4L9vVe6uw+6J
Qws2MM1Y9YWd4Yw3TJNFYnscomUz0kFzy7H3yUKDzMHS9Xl4phF/RZCv8CeRVaGfCtKLQ/U1SV9s
kZgDVvGiAaAOFcfUoomT40V6kd+mx8ZZjbjoCJxS2y2ftQQq2g/ddhhaAPAt/p94tYqobhw9zBKE
GeNYh+QG91a59TeFnbmYEhEC2nHPu9awX/1spK0hylr7jJRovCCjUNfSJxzExe1Lo5sUmtm7l5mb
WNjYaR14S0ckwQTACJ8fAqw0bAy3ZiOBl2HJKiVNCgZAV9MuwSFws7jL7LJx8aEtnLV18NiOrbrL
O93CLbnSMoEz8KtJQcRbLEMGYH5KZlit77Fs7x/T5VUXUhWX+QO30HGe8qkfkwzxa1NdADVikmD7
X4lZct6Ib+EvKmCh0ZcOG/XMhxfz3138UWWBpI+tEQd2k40AdoknW/7ip+ZNRqKogo8wA041aB2W
a7CEpWetHWnG/zR4mek4caqwb6xe94PHhAD35MtZ48swf11uugG6ShiIoXLSTNc7dMSUOmbsL9P6
fo3fstUmN+x2KzGqFWNyUpid8Xl8iC6qLzAWTpfycEiVXRf3P6Oq7O40yPf3llsEWlTddpvguyTo
KXFrNmOPACGWjmsx1+V8Sir71C8aKyuMhZ490D6hwbbyMz+Ez0WYH9WXkbFT5H2CNTuF+hbKQTpb
3A0xduAmXJLfpf5KmX6ln+m+9wBFT0WGC2lSw1EfjW3dziOX3tAhkTY7hdKy0PKPD8HTF9qgnC3I
KV++aBb21r+XPTeCUgo1+vQYPV8ktezHMMF+61spPnoxNlP3ZfMOr9hVellukY2CdP+GTEZizSSW
CnrCZFMi2W1VKr/AMf6qY3N6WXqd6s3/lGxuH4ddnydxNL9XB2WH4lIXaLftESvjWcFKWCqPZq69
FC1nk1xCzNZ8U4qpSvWY48pkePf6ceSJF4aXr0q7Nua+CsSx1MJGSuL/YqGaVCUrkj7JLuH/Vwox
8jtGhhucMCRusfnVAVmQ4qzILT+uUD26XInZeW/3u+0LpDwJVhPP7SGL07UGOilT1HHni9D0igsC
8bF8wVsZOYHtIwOdqi/DOFrvOIcxkhmk+hsGhKJ+tPs51qccRjuX1gezIN6LXPX3YmF42bzZShmB
BNT52fyOxKkvJtnXQkhdBvZWkiv+FMQI1/eoFOElyfaktvz4xFpAKeJAd02aHucpn5Np19gfZ/kn
5mnNxf+TSPO0DpuLgnhY67OzGwh8f0wDaSJYuKZdmiLB000ZXPpJaZHE1X1dnJbhcNu2hN8lpcd1
5af+Ir5gwnki5WXY11I+O385KB17SFoO8tsiIgTbBNuTO+lbz5Wge2EKleR4cu/Oa4HiR+6YVAsE
lpfrywsYpTcVYPrSG0qEsftVl1V836K2WlgdUg15QLMpPz0ifVUusev5znYxp2qXYkxsPwlYaSEM
NwMmPJXyvkRT++hzznHOshRqJ5/BeQjjheMK9zhXNzseKrQGWAbgtFt4oNgHLeEY+yS15zGKnl7E
EqrV96gnWUSjexUaFkpKs8YPX7NGljGHhBif/WmU9whQW/QGw0LNrLVJnPVEc8VG3N9j3YGmZ9Kj
ZGrls8RlI1hR0unX6Y3T98iWkZYiQ6UTmyPsFyOrJ7kZTP6Q35Ftqb+po5AwiCCW1WBhhJrmyrNo
zycXRNKOK5WVOiUGXwGsEhopQ0KfARHkcnccXEJk/ZcqUR3sZdYL44gS/TiGN63av1BJil1WMoqW
HEYmbSylMgrfwGjVBT8rYaTOIdik1SbB6dfpTZRtF/cHHiTaFs7SgNouJCzAoQ7x5cxL6mBIwDFa
1J96K/Fv7gsMvMe54Puxo5sFXKxO0rIm5L1zSM24SSVVJ0v42nS1P6zEHfHPSZlHop3rSF+I1maH
wX0XbUbWnwj7NrhL29gU4uwecpLLNrin0NWorgiDXtaem7nOdYmO+BY+gPEROPJ9WZFLR7sFBAPF
VLph0yDV1vg4uedIq0HR26fjetlWP376ECtLmRxWXJrCXD3J8S6dFNwklV294obIO8lnIZD7fjt3
ze4ilzcSK5F6oJcA/9+9LwAX3EHtHwG+G6MSAPrUsrniyykyQDzd//++loTbX4n9ptzdcPtq29Tj
ViDGqHaFZfHWUroRRXEEPgdU8mEdFli2t5kZ4jkjYQzv98YUT0ETE3ndRXlW6tt0AzV7lt/bpy93
/9rFz2dqmBoiLTca48ATA6Q2XuMCEQ2OS0NhYY3Aup36NHFFLwyOOYK0VvYqBkY2RJTgSyux7u0A
pMVIax43Cc6UuEiqjCy2DyuM2jN+DKFH65CEhQwseEXeHOZE1OBDfmgw75wWXT44mpgXm2WRb8o/
rITv5u3uYIyh2U6QjSR9T5IOIiefK2kG3x42EHcWtyz+ZTYOg3OEMenVqS4relpS5mqCOX48TBZy
NeyylQILzfQ1Ss+uDHB02B/TTOmY2RJT/BrVquRE+2G+oKsf+3VHZX4o4E3l/KzAofrR3L4NB/l6
iIIy0fkj0JV6yqwARZVwKz+B5nK9TNgDgdFr0M9DpWqbcb210zhjoWK4gnWtshmuY5JP8mJJwyT+
X/9SFQTraox97yF0DgP1qvRL9LfwcyTyooLG0H/SsMq6EdrGI8e/e4G2DEQyDjP33NIT6m6pj2w/
78ZpgN1fnNuDTRcuRydLSVKwHChiBVsuW7IvoqmcGm+w99JftadifGjxHSDtiW+xA9q9r9U2/ZDq
3jSI4k/cOM88G0OrpF1j8JiRZraYcP/FVA5dOkfF0a9D0mioe07884z+H+hfgmzW+LshrRKOR3MI
12wThShaNIwEx83PCkHfSzLIIiOo6g16oi6RzmWV9VUgZw8OhA1b9feyJVzCTWk9GGWyS3h6xjh7
eXwsJ53g9/apIn1xG1P9Jkjci+NwE9VsMEl2dGAgJoFT62QxgvnjSggXkJzh7NH91gKb0m2baQpT
NJ2kRPxGBoPetzUBuhC7aH3jFwNnjNTkDe2QZ1tfqF+o6ilXSC5s0Blna6pVuDr4L6vu6LWFLXMa
Vy3ak8TTk7o1j5lTStL406+GkFR7v9fQnVxciXeevT0V/iyx57ueBWKFB6s/xGPvf9cBDFh0rYTq
XLiAVLx17uHMynwbGUf1VewPCxCqimUeApOcoKIJJjlNV3JKFl3UAtPOpopM5qKhzOeeUJ/E3x79
xszJWkgvjRX40yUZAWC6a590mMpoeUjleZHBdSYjubQ+FXFmJJNDAKQpFZfncKAMqB4Yts00sANa
Z6/xIslX0Gk/Y4qwd47HHLBr/VcvOPKX8eZRulh5s1q7yTM5faMFm1r5KeRpDThoP2Xc+LWVRSn9
p5zCfVC20LaWUskSP1I/KC4tYGY44JMn5lx/VQ/g5IgXd5HdqkM6tSUzzkPLSMSVDhk94HKqXxAk
JZBC4QCrcwsAOwUFQVZbwTxq/4M30BzLHxTeG9LgDdRRNZDHvR5nV5GyRfZz2hwJN4vu8yUH3Nv0
hGf1BDdlyWcVyoC/bX91p0WOSrykKEtGbYVM7BxmGY8ebns1USJhSRhwOV0NdUqdGYS0NWHLPoJs
PSdyCew8ScCQ5ZxmEtEjinTvA/rAx6Me+RbEjllhlfOVwzwGw1hEfZVDRC0+rO7XaGopx41X84XH
nGBlXDIBpSNFhgr2YzhMz5Udijqkl8+ejniEhb7p+PBC6DJb4mc9pfKqfFv2wp5zTnKZPaiFBysX
Lzcaq84gntSChwgccp0QUWJgRtxu4LlmuF7i8xd6eqbx9E8L9mmSokHkuR4QZj5ThB5GKluV52IC
Zd45GMOrXPQXyrjWFftSHY25AEu1Ea/9y19/hnPjameSSQ6KIHZbhp8ymNrqMJrHtINkwz3Ctr2c
QTt1hjacO6qYzs2kOl7UWCFPiIkfbYeNlFmz+y8Z7bfzCRF98QNHb/oTMqvf6ckvHutVohI+MKa/
Pzg02gomvstpU0k2bQoBb40PGjDcEpG5RgQVNhbSLi3TGR4Am5eFOktekcGaGNdsiJw5Vu9NIhmF
zGP6g8uO3dyM0DcxhkFhyLLUTOixQzyAiYDZ0CGURJOK2xVFWRozaEpF3EStBpgIKjmg4vDpB8Jt
P2T3X6L9D0IL8QPsW5s4TVFf0102Er7/m8H2mO6yU6xeTrZgtW2tpPb277P6Ih/MIgN6enpUyje7
2gU3fHQxXXSZIE0IpGwOeBD2thbXQ7vNNecWgZcxrL0hn6hysObuhDuozGEnHoytDyqsjfo2ZhoM
jKj4AGrpjWqZpLmFRZto/0pE7Zx/AagsclEay1Nucn/wgzQLR7h94/FtyafPvx+1MgFdyi2pTgSS
V0aI9cYheQZiwHj295TGRdFgtR8ONz3695iwyjHMszPw1kQn3gsK3KcjlQ4aVBJfPqvbR23PkxiM
DOJb4gIK754YKC2rbsk1EjgNr6COBGGG/dyHYY9zmfpAMwGcl+Pa1dgahSnIBJoJbfFkIYHvqWqe
fZ3C+8j1cpZYF8tHR8/xwSEkfSd7Im/ARwOBIB19GRrF16N5qbAA+XA9cFg0SEaOjQZs7E+V3yn4
1fW9bR3HszEhonAKY+ia8vkqc+EB58KxhV+M/emGiLkgpmCLqNw1WnJtSiWHleHNUafOrl65PQvt
ngIsdnZJOviZd/O+9Q+pKxd8/R7SsTgYfELYETM2sCxV4iLkM1ZdIvYB2MNc2E07NSBevKPUa0Ct
+RvA0QpJhlSL7OKXmgU4eZlDJCq+Q1CN31+bA6eXYHKevPIAAs10VRZmxfEVgbs+/Tx9vXCPjshq
ezSunN1CIVanAUWkBentGJC6SfLp23LPe74rsefjieiGmWNE6Ti1z2O28POyD8EAJQdm7rar5FQf
TLwj9qKQr5PCbn7hwn5TADlL1JrkngM2w4nA62O4iAhnLeS3Z3q279jN8O13R30pE16rPjQI0SBv
omwy3Mc4CFw9RNYqaWj09xkKv9YlY+7cd32Lo/lIt3+44ObT3fS0pj080NC8AaaroV+UV7rjbHqw
9i9AQRRpfPQgks5FYcjbvRlqDlSE5pU6o58kyzb+JDTOQ/FvaRHWK4UUlB4wrQP/kbCAo2+AgvjU
YK7r4jv0mMifhxI740UUf7DEmUInnMIpBsrSSrzL64o/cASqXG16ilKrLpDSSTqzVXYL1oTvDtnb
09Koj+obKg5ml9QkllHntqnBfxphFuEWjInO0jOUkzCKUgdsW7oIiZrpwnRf8gd1AsTPZKOVrztq
dqtcN9knn0+nCO7yg+X222v7+muaBrfpl2b4fcd7ZqhRQMwZmSOMGNFDsOxF1cFsF4osuIpfANl+
UQUuVXMbt1283ZyiRsaR4TSg1fYJQwawEXfFaZwjMmFWfpFpk2h7uEwD+CE+prj7DKhjwsFKSe/t
oQ3HGyB/fKX9IJrBqFIvHTVuVFWQ3p2vukXjhqahcXieP4MqX3fyd/6kUm35I8odigUXXnpePUJD
stwPH+uyZ+kZXnavx/TYVQYCkt5AcRreanAkbrunT6JKYhbay7j64+/INV7Twktgcds55raqkOns
pLXPUYLm4753XbQRDu+KUIpFAMIxgJwLgq2dQjRUUtC2RXcjjTGgz3/Ar4UWJyLG/Ac2K/kkdpUf
GnS637x5QoqbBDqFCsDYz6uVJLqLPlRdM1dxO0UB8T8xSbJGJvbsVh9sEbgA1xRymDm/VH7TLYBT
HUoxuewkPXNSEO8cePrsCEdHuAgNLc8NRLOSCfnoymc1O35UFs2co9GhR1Isj7KOfAPOBKek9bXl
XbkSzSIdses2P4xT7k3tJahGE8qZ8cMz374fdzPpROEsiUe8EjjzI9jYeJqt1jAAZ7hKfsFNKSQS
x7XQSdoOdSUjs/+asqxXIB3U+4jdpFVfbAZb14sybkWZPKXUDsaWBY371rhsFN4S1K0zCJEYbgSB
NeVWLQp2T1CApM5u3rMR/2CyDMcNEZ0N3rdFacXZV4fnGWSEvKRoysANuAYWPnTtO770mu3BBFUZ
dYQMLtoE+eXa3S9oUo5gvVi3ewPbCZ706OgGEywONEtW2XjB/JbtluGGaU+1rNxrKM7ktfvWAvwf
oaIudHHcG0tLrA9bzmwBfThwDwDWeox2ITFh6XC/WETVu/dEwEuI1RhROpFz93WezNF5hKUQVEjd
30H+KWb1rU6oPQ9YGF75uRuGZRdwGFKytd+g1kYxEHQX0AjF8E8naMa4NODrijqSrYYxfdbp6/Wk
b2gyuCw23y5uLxNu6qUoRJ5qWCFQfL8wXFoFXU7FSt6d8MzsJPc38whB36F8SX826g3gfKHtAgph
IXrRt9yWTC15djNC5QoXTx+TzDJaDU0dGvHpDZauly3WVzDzkpYoXUyIP5iyOlUj1By0LSU6zHgO
v/G4DNTgXCtMO1h5xTyyXfl0hmr8iL5P2cfnX/iDF/IfPJYD/miv3NscXuhkGuYrjoNGlwXZ8NIq
XDMWxwFmKrLDaQALYTa/WFVzimOUZKWbKUHaR43nIyi3/CJHHnmnXu4nVAyvTVLgWUbMUTZqrrIc
THuPfN0urVa3VzPc/9tAf4YmY5PpJpY0Eivq2RlbbA6o0TTZ8fK1ujy4PoBHaRP11o2mAHp5Apjj
mPOladhIdYR4TPiydTYdpfrGpIM/iWF9LU8j+xRqcESDhu8AVTFT4oXpbndtNGZhFRgOQNhIKw3D
ooABb+KQO8MGvTHJpGJF6k+Wqpah6JQQYToEc6U1D10i4+e6zmQfQD1Wq2Z/xYKHL4ILshM6wgrj
cy6Vx4MhjH6hzLnf0T1gaxbGx9VBL5SqDEA1WXzpEllG+83/IDlqDWMoWwQcgLx/sI5Dtv0VeX7R
ecy8APsxFNpQqpomGJo7tdAOgw0vNkPmWKld26CAGCpIr9fqZf3zVC+Lr3fMFwtjujMbMKepzMAh
n1YJTb7SQ8jsjFuAMTl0vEpg+KN2gEdzaAfeLZwtoGqpLPbPxMaNRojE2IzCU7GQfAZWaoh+t8FS
1g8CdHBj3gpbpoAttwcSFS5BzorqwHJ+TMLfBCQs1HUYTspDa14xMbtUEiBcW9Ja44eLpxxW5Bq5
g5y6VWi8y0yk9augVAgH/37YejaTxA5kQ6cEYLMCEBdnkXE3lGKJ89uMpjeO0KAYUNXwAVe8Jj09
5c9KOw14lskBHHIL/MXNIY9kT0Yzuouq5L1YqW7EnssSdCPGbSZ+WBsQ1js9qINXKnN9kwLT9yIx
vIxw1UZDKGYRElXNqTurJDi2Nh6wWdzq1I1yjIHgdN1AcKFgSkrf0YyYSc/JMxdLsRqghoRg7Lr0
UrLlhJeQBggyj9UiYijGWGsWqKaAdNhj3Dl0BXqgQxKvbF6/7ON3+8xDHc90EAQxdNX0CgLByMfZ
yFJE0U4mQ3Znf5H5w4e7fY141CrW3EQsDKb1K6Yosmos6Fcmpj6Z6FskmXKBKqCrMWzux9jNY0Jd
2hLhRGxNNb/WYfjV/wztiIcwTDVl33Thnfx5UhQv82Dty6QjTteSXCmD/wfv3lQL0VJPG2gDWZza
7ImQ0gdBt4dZhTTs1Ch7l/RQeqej4lpgcR027uNJurBPAUORPMRJCfHmN/NXPDePcc+LU8d8ry+e
nE4cCqz5RCRb5vvNz6fHyRgYyzzhbaa/sZ3vWhhhN76ec51EvXfh+ioCLOFncdR4GdhD1N0/dwWz
NuxBWwnxrjkoToFqGU2YRIdzkIlCG3WMKJ07IRacnKy+e/jkEkJn6R8jKtxW1a2LXxc1kD6j9eGm
ZXtFaOirIpJ773iPc1znDmwuumet528yXoJgG1Sj3dqp56RPNT//nE/os2f0EbOl1/2Yp+s/cDu4
nwWJiUFjOa62ePTEId+6e1CRhgMzT4+eNt73vwjyqvv2BVjrjO9wQIAApr/qcN2CEr8npX61eYcY
zf4i68A6l+6+h3eYYErA5P+HYtkGhVv78f0o9rpc8l7Zd+paCkZEsK15eg5eZPRSrEPedKI5gBNI
DEc06TweHg1XHjWUZOKKPzgcVWEGi1Lwg8OV33de9zbMHdGyE7/Csb2pywQVXVnU2AWWC0xq+ZRR
5tRFe+QylXUmwGsNPYdmx0oomNXUlE2CZ59vrIIp8Bfa9yKOsLQMWtzYzUvc5vtBXEHq+/PwDQY/
WPcDaqCLLNR5pCfBTTCRmXe6UZ26JY+elPCn0ZZrCzane6go+SUByMkIdFUQj66jcjkGijJJBNKv
v4durs4TqS6IjJhDOb/dSFSbm3E3NPKhFwpz2pxNKTA9K+N+0uHHKowYaK0AknsAb6dhJYkvmymL
d9ZkUdp9pIlQJLlnSqKPBhXW/3F3UPigQCtRt0LmUoBcG7S2pBvg6QXAfqdjpiv4XtNMGzBZCI6y
XNuvulICkpIHA1gcN1hxtGsI3hzM7KbMxUPPUEQWaz8ziHiOWPyorQlQJnUIdZVYqxjwMgUW7mcL
HfN9XEmtaJokpmuCA7VJcZGGY8UhdtXJ4nOzVrypbqsA5VCwldYVKctYRNMQSnQ8QcrAivRehpox
LbLmd+y4NU8Y/w6R32/YOec6fsims/eyPZv14gVJOHcjA08ffr+VjyWKmRoujg6HqGXOKv2Tz8VD
PywQtSb/KF0mrX8dE9D/ZheQ4YmeF0Bsig5X0SshDCVxg6/s+EMltNdBtH/h/E8vNV2DB2b0cTZ2
G1hlmHgqpqlXEEQux7yyJ/TmKj3DXUJ6HwNhPVIzZJ50RA37s3PiDie57PWdkcJI1lAQNJwFUx9K
0ih9UI+sB70FGd/TtHEx7c82ao/cW8v6kzzr9LMut6m/U3EKH013coA/H8sNHzUhI5OfxU/9erAv
8LxqyZ3NgWjfjhALWBjZLanCmcrayPKz5PSSdhCCFuFgUJitUb82z4cYRsX4kuBBiRn64geEp4cO
MygK62znSbTm2koNVsE2LZg9t7xKJEZzSYRJr8yC7srmUoY99WGQC2G540U5UHp4mPG2NYGk8l3T
1yYJgE3CmxCs19OMc4WbVIM63yUyUeld70Dgu97DJFtibGVTGUdF2k5E/8NH8lojmIUJB/cD/ecY
Jt5oYtZy6YTMEhbzHN4f7ky3VqmlbfjT3h/y66UE/pa78lyouLrM8DuyKFY7vpZuXQsqWw3IUaQO
VNRImJL3zAJ3XcsAtPCTschAWP8gJvddCq0Ul9xymImscPQDPkCBnrTuvxz+2UxWZM7KDvVxEN7Z
assO+M18QX3VgwIlGpgqebbmWvHKQPTbxHHyCQZBUdhtHHHiIpLSCxNTnV1Tn4juYBVvHv/w0uny
kMz3hlfqTOP0U+z4JYLDaiptsb2bFvOhmgv81Rm1V+ackNp+ASYfuHrZ3MIHZKWZfvCypKwzscud
cAnzRE8ilcpQlgbzpnE2O8alKB6s3F93TdnTduQH5QMqCy5dx0BACGwXqr4nc2WDiNtbQ+fzPGps
ciGy4+nZEU/eBlQI9CGRIg5y9w1KG05NsH3XDjS6QgiF5EiU32qotZacbHcUJIjLHDNwscdvfrtE
MlgJAQEtBS2RxO4vFd232HxBCdUMbaIcPHzVyA3uWCRNJs2xDZ+XBzAVGDCEW9+46XpCRFi+SVT3
f1ch+QIOGz5oyuxb6wrYr8MnAMjWjLeWqL2qLSGovci8lVeKJd9fAeLvWHyIvN3F2kKFjncyTuNz
v64ue006+B0vNRoqs0BchEFAq2jdhbzLphv+7LPtvvSdspeO9MK9BopaQsfzja7niY4W7CfOhvvx
C+9vy3vX0pTf3RilQUfji4ft3+zNH5utoFdh0jC94Z24NFgFwgFR93EWfnsccnFN7KPrJlBb9X+9
BBpJ2WDrv38uZtdqiLQrZYmZiz3bbi0RL0QSDEHEFr/2hpAGUJqAqdyfvaan9C1K87ua9eCVIZjK
JDxkWrK255fPUcqHSNrsqVAXwO2jXy4jJ4ayaFLktfE7SPdQc1hiw4D8J2VgCxjCrXhNXHlyMjHB
b8HMnUAa3YkP7+PRRHqsWB4XdWKjdHeibPpJy14gZekLuyGGrUJm+8B1flfwK8wHwCHyhT6Ue2yE
6et862EUdZzJtzs1QovFL5pEwR9Jp9MdC1IuuslvEy6++hMKzUzAdmrvFIAmWUaKWlvGL/5qdzYV
++FGxbMuKAuI7U4v8Wri0cPg8kLk1xj+Bf00//wqW3vio7CKUyM//h5zcLZfPW7MQkYS2d78viJ2
l9uFNkG8IXJhSQpKPDZM3jcG/QEXE95mRtS6PIdjFhKwWu8+8iQ5Ddtu/vWr6rhDMyHqVismONZM
Hnym7gHio8JSKBIaJIEd+lZWnOgup1HVpKlf9bz04V0bDE0a41Tq5arbZ0GdXpOq5Ku+P3KMl6HX
mJls1Omb4kqcxGPt6kFY2pKNZWGKDpmsXypInUy+0j+xSezwB6CBi/5NoWz8uYfamzVI4fxzYbBX
C306z7Vwpu0oiELx0a/45xyaZfSl4+oBCavyOcsC6xhEGOi/iaqK38RnYJ/CWoQoZU04onp+vL3D
1T0zIz+JecPhJQzkVuk0VWLh2T49vAZ2Vqmb6hmQmDliqK+52wsVwOH11PKvhuGcImTeuZ4kvb4n
D5p9p0q+GEnRRJofAi+/5KzaAJ3o31opPK+nGrruJ1ZFm29YDQUMwrmV+SkZam5rxaqWXFX9EitB
NHTq8coFml2IyJeyEmv/CDaGkuYBonwR1DpAgM6lhUL4hkw+QnT3kC5ZBMTDPmYybcJVvOen6n0Y
dLvGqSDJSZw+AxDp/UZ5U5XkCcGIS/k0wuT8aKhhaKOyta7foROxcBgzDUrUouE8THtyr3Z0B2tF
rVTYQG2MuuRkRc3TyUI2OEXa1II7ErsAPCy23pKh1ySKup9zw2JUaOlupURhzFTVoiM1VhiIkhnH
eiv7271GO9ZykHfQsI6JtM6pvHo7LU8ZM8NMu7YWhLpogekdvf7HtxTeLqRPg4zf1n9hhiNAcC2E
UsD0Y1aPdalksASPfX4hRdbspNlkDY23S1iUzsZy76t8ek6awMR3hoz+SBUoawuuo7jF6MNSjsPD
OKP5dDocMuszuniBnzD6PGD6CO3TGAsMouoCHSFVdUqoGqJBYdvDlp0nyAS+ms1yOkroNa1isgvk
zR+CjqbKpDlhXymg6hLtPpNkaTwet+g+wnMjaI6U3bPMNbvlOCh4m/vMPz67DxOBtkSX7tCsMLQe
SjKHFbvkpf/RpsBrRFwWeLnb8h/CNvaX+b5eTpH+cAXwEvR3hlywS6gXnWm7CWKoxfGlzjCkYFOr
FzAeDm0FIGOAPhxVEWcjhNH24FzQPYNpvCiFITqfiXvEQUtam8S8AD9umg4uXjpCU9QjVLLMi9ew
cpFt/g2kZE+ul3cVxPU+I5rV7nOPvubIKgkZ4IVxZ6eQm82oeRzJoYxJWpTqH1HbBCHrSy0zAoRE
dNp4gTFqj1UGfgtqav2ssK/UNHSnGSH4iQ1prMQtmCsFdAz8lC0dv4o7Y+CH0ThCck/PyDhgN6km
3EZqOT4+TS6azQQlV1t1amFGc8Ws9uDVU3B2mM7ShbnM5S0vswiJAwhaCFr2jbIgjUUkidibOqr1
fdQMZHK2fnBAJW8KxtD9u4cFIqSiFfjSDj2P3eJLQVxj/dAlrHdFzXDg1a3T59A65wge5WrQ4zuR
87cW1k76dhsSUPB/68hF88U9bASRutzPnyM3/oLKnD1n+Saeg6rh8racQfCU2KmzMEna4K5zTbi/
//vsyLKPHpUbI99rhWNxeJJcfLPtvYJxNnhEPa+coyuh+EdkDArdCFfvrCipyMufGEFECvppeV94
ThFcYc2/1XqFXMqOPgLzFokV7xsV7kYywqBDCSIgwcf/TLO8yvzTpmnF2PYhV0mA8JtvuWrJixB4
dAzwGKZTVfUp08HVJw9w1froCJRBbJf/vAW/pzQKjLacm45D9BdQxtlAmEZOBErNTQfy1llisek3
0EwSO4BzIy1jMbcKNsoLwiJj5zZPaCemFq70eUBWLzgIZy8EH1rKTqFKoHHTDSpQ2talboccWMM3
Gky0lQRAtveYze6hNX5Zc00YgiEU/CVau9pGTLftUY7pcDOvSvUtjfhsdwd1LjaktbzpxCxopZU7
ahtTMrFOltzGNaueacDJS6nvY4V/B0YhdcRA057Jx7a0/3dDO2GOUn6FOf4y+oTqOI7DdqBz4WwS
ChCfjtmJT0TRLJVov2LXci4j1WzNWMmn5PzV3ER3QZxqgVDQ07hL6qBP1/ebQa2zaSzLFaPpKTI+
IHzUFOOYm3RfTN4pN1m27eawio92GSdftApliD+N+f7zTD1bUB1qXNKbHeFztIwnuO62z3crpirQ
lDo97JH08fTUrC0QJX15VlKiuGVFo9kvyF62ivPaobhymRZJYn+aVtUnDmpsZ/nf1WV+Jnr2sLS7
qyxMuiTSUke+tnasvBpxLPkyID1dv4kXcYr5FyIatadJ/RSHniaHndlNmb5ADN6PyozCxDB//n9A
76rrCKqw61JIOtHPvPic5VEzER6cX0k+GOC45S6FD9katkIEospKXaV20XrHl/hV0V/T+luS0Igv
jVK5xreNVlcYWpJ0xyFhbRMkrNJqdnNB84LXooM4MKbzS+hpO8l33dHzIr2zP7fJTQs/V4o8zgKI
ZXP85VbExnjJqo023wv9pr+AwJm9Hbowo+2vBRkykEg+pGc2Uw7qFapntCXfYvmxJLSxfrOLm2YP
/DmcFyCL6j1t5DU1nh4RGmw9tm4G8velsokv5y+/zzm74PX2DcaElpq4wiVWhAtybkwGhAwJbK7h
WYeQr9s47fH7E1uSS6lph/iVTErG3z4RMNIiaKmeWkerp4xyCj2ZGvK1tvJeAfA2HJfxI3PIzkfL
Gq7uwRFN/SFG+bnEedMs65k6Afsy8rIQt3VKsAJQV6CHb1t7YpNnWmhfLo/vkcfol1x+SoZB17jg
bk3ABWkZEtoG6L96wa/JBoQuT5efLo3BBTWTwG0/cMv/7TSyFn0ppF/CtyH1JBOMdLHwfvYJGU78
eMbmWCmrfUZzrcUoNjJMKZWWMxL1HXW9DJTp6lbWbT0/UIhZY4aZc6vKy07pmCc3gLugAcueWbRc
kCC3fA0as3okvQO1/7GRCZFEbJ2HlXF3EFgXbSKY8nunaPDHWSjhR8PbPKgX75Tc4Vnhmq7nQ+ga
y/FcFd/bzI2Yw8xlnAgbRnA3lZqEsdfO0FQOSTlwlyyc6kca6oRTs3KRRaWr+Jcwk6ZpVfep/S+O
TuwopPrVhamTHwJaFiqSmgcs7SZgYS6uXU1LSCGgXbiBq6KxmcvEHgUCk4lqDwCOt/tGAv6H7PaR
DVX93YVBp0E+v8uBYZ1fTpvQhDdom7+1v3NsJA5ByBsDorKIfP1nH7F7kS0kKx2OJYd9ArxCb/FR
lDPlGs0Sn7TCW/XcIj24/89bQ5JkCPXl/s7nO7DQ3uAaMa4HBG/+JxK/FKU+P98zgJ9ChcJrjC5E
TFYSFiINIBfCwo+wHcOC46qii3Bt4BvPYACFD9KibQBmaDEznDnRqmkSFoFqp+SIH4Ml1zoEXG9f
8mJSzIbW29zfWBsDkNKITlukXowh4Bj4gTed0JhA1WbC3ST1Glct93Ha2q/iivrCFzdkHqH0dxEJ
i+On+XF0UeMXbkfRqUewnLboz6x8nNbuA09BsT+UKxnVa4wXS39ma5JCOje++p20dXfjupuFKXpg
BI3sl0rxi6ZJLygeVF85tNFnybN0fSCuErwIeOlzVkdTg8vUcbk2RU5jwtI9mokxfEhq2SJl/BN9
YAncCp5HXyGr2feyY1oJqyOHAg8Kcg2tr1QSXAtxedvO+5wcjCwD5fOZyNGL7ECQLn/54TqGoyFP
b/tcLHzxOkuao/DlOThHSKHKR0MtqPkLSHy7bImuWfKH5A4fyXnZRma3IKVSKn1luQg6VJ3WnbGS
/o5Bgf6QSxHdyGDO1EZbahD/d1aQ9nIbpx3tE0CQ/k1+/vMm3Awj9hK9ZOWtuGSLrEomgsSC2Q1A
m7MnbCNUjfKiWJOhKTUAcC8P40j+E1dS0W5F12CKxFZTe+CNH1NmxaEUfUQf6FXfwX6QJKB5CO6L
if7tXoh7DlTaBd2/EtyTDjP9YTw2iPY3qgobZX7dV3A1jZmEy1HYsCbMF0/RGQ43VziCBW7LusEw
VKOpc7ev5F4GyFFtNjbRt7ySNJtHPMlJOmO9CUuXkz4KPj6YPVCxrWpC87psbc8cMs04KBNgmMeP
uVlvXD+b7HzVUZf7dWU4rNVK0sgKrwWlD+6eUqGnFuRqhg5pg9nDsfcop4FIUTL8wCAC++3VtPru
Q7ZUrv439V27X9HRrRDwyfA6hMOREvIvE9yqQPRlKlu4K4eCSesvfKEKwwpvr0R9udbIFcj78NoE
mNhiioVafzl9gRpqV/oaXK3n8DTXBAIqBkWAmkSjLnYKvU2gW0tt0XvRroob8wy/kJZ3IaEPJnE2
thQ6D5RW769RNWucs8uephnT5FXz21e5Jxp/h6Dh8bKHIQenIoJaj52r1eHwg0ovEUEiZvxmNoUw
Bjp4hbxdNN6vcowm4ZhhvsTAnBLub94pGfs6GgXlZe5MYUS9XdrmM1B2eNOPtO75wzQ/wutmTva7
Gd+Faxsn0oOOuwIPUzpT/bz8dAxMHWMagsUKWPbnADeuS+QRdG/14gdeU8ksHJMQk0Qcl08rTr7X
VCxZfh+yGFaoddl9NM9zPA6bpJ+L1DCUHK7AtBPuk/of0PKyAsb5gLJ7su5d0HOS6LMhqKoshVJQ
xr0MkQXwhec5k0rADvf5CKBZqQxV5TXLDRiDIzNFLwFXV8kxLY0CDlCDJwEdTEvPDHzXr32evlbT
GNmtUwqz7TU2zImC5kQ4aRnPtMJiOFdYLMXfF+qmuZ/IDc2plPSfjFDk0P9K38horpolIuAUDzLb
M8ngjbEdZ9GHquOMOYYl0zP1ZsLY5TvtXuatuMKIxW9DzyelLNYIz7PvRy0QQc/NOXp0DkTcfWdO
XV9cH/v67TTEqnMDlva7gfA8wR+X23am+NiKgehvf/gv6eW3rSilNT118Mjc8eboqV2sjC/rJw/M
tZ2XHuqyk4Zm9IDu3otr5q/iOzE2UEHBLxIjDRCBzJo8iycaqMf/TDbSKlQPBbALg8zfH/EPkJfe
6KJmsWJAgHAHY1W8U/ZDRLCPf+zIecH9zDkv3H04MBXenfpPwBHMZNGmoMhmKIVPH6d0r02b9W/b
Oq2U8gA3aYSXxeQm99k0RvDg7CO/CwRRS9gexViueJ7pVpIijnduNoaqL5g+9oo9jzym/pS0l6up
e1qC4ltI7EGWtP68UWq717hhqtnDcCeprHwwPS1JqxG4LDT583MzDyeIvHGrcSdlgqsjaFRFeBO9
1s9+UMAZ2X5KSQQCu8++U2VlRPDlQuKN9eHl5UV2196u98INWkQQrj7jPpuackB+xeZWHor3nCpc
v8CmiBvwhs6uQA77tJIkp6DmKEhJh2XKCeVwfIgPrQjC8HVgwb85x/rH6MuoPKse7c4egFQX69Rx
jmv6dlq8aONXC/4gI171Sd3teNOnKfHiSF/eaezoj36WEp/udHPsjSu+KD0Fu02Uo+bEK6z65R6m
ohGdvC2dyrQXX2IZYWgrV5AnIIZTq2/RYU7N/GkTDZDS6G4PjGXk60/gp7YFtc5LMQAvtmSlcu6R
ckfwY8TIDoquv0PiMAiJa2PxR/fygUky++M8XsX6d0W5yxWtgYp3VmPbZftNxWqQBaspoPHl78b8
1f6QpP4Ttzx5/c3YSLjWfSCZ6R9gBj+nrBmE2WUliDTso/rDmCZwt6JAziWOfDgeAIPcdfGHAFjq
RxfIsNRVjVqIZxNta/Hfzm/42Vnbao+BUrA7vXNmgDPr17ndRhF7nqeF32QN+1j1zaY5Z16uaTQ/
ukaBIi66Zb0bfAYduxU3w6dxzHuUrQb46fXEM8nnS3qM9+jmp8h9P8jQOHigXM7aEyP71Hir+Zi1
FcbuE+et2LYrLf8qGijsKDpreXTnzz1yGar8/5h5JhulRarEcZeUudIGg5irZnaKeUmTXP39cAgc
IJifgpE1oianfx2L0EUxvXRaB8X5z/uZgSaEHQKhWnOH5mJueJ6qP0G8ExGE0VJerosZM51sPWpD
ePLqVKi/hfVGSQk47ucCYu15xgwj+OOVci3R69goTMZCeiZFCj3NdHL5qIpnsr02qGtCwmZXj+j3
9w7Grlk7wEEqtNysgY8twwjbEY7L8JsQ8xthCVCIn7PYovdMuPra49idtv6E6zuPjP9geTpiePgf
NVigrx7kRqokvwKmUuQTLRaj7myb+qmua+NQn1U1fi9fgSAAKlEPKJxRuCoU7InUtQLmz9AilKs6
4RWTv4sF5RTDXQil18x/JFMLEGfcmpcFKZa74W1faKOymI7DM/lTIupypmKftdH3GCbuLQv/hC9e
FbiuSHvabKgu+vqjOEyM/QGstFqIdeuKNVoFr6XoEpeSmNq1+YGP3GMvym5kFabriNweS0smLQDh
Th7HgJjXTMPXw8ouyoczc8FItIndSy5339PAI09o82T5/DEOFMH4beJ/cSc8tje+R5W1f2emm3lk
z8R0pDUZ7HL+9EmfzMBW7q4g3RjPSkUshrvyanKTfvuggTn9OIyGiAvuwvrP8op707grRM7biV7Y
WHQzwroFrCr7N/geXhTLGQ1EU6Pnokg8XAfCFRqAM8jo/Ga7DWZEW1557ImIpwmWRpNF+BBBhgUf
Pux8JV+b2wfGu8LKMVnd4p2Royz5vAQyf+DtslYH1pGVkaVTX1Llp0dalJB0JddyjyXPjSDdUWLh
mqHR+dB8xL+4tQGPj9PL8wqtvmbOEAaQ6MpcXH4qtynap7vv4uNBR1CWIYdVXjIgYo2RwyJo7xjg
5DF/kFwF3zzw5vECWK6XRiQVt0l64Z4WIpqD5+yh+Q8D2LWwMBzZljT4zLNVEz8X/iEZ2tESQpLV
38+S7eC1ajzi76I5/jv+4op+jrN4Mnn+KjP9EjwF5vprdGzjqowvasy6DhJqlMLaXVT/as+xajmm
tv849215ShZXcA5NNmXuTQBZVmSXpnqNAM647jyANa8fdgUR4i0gS/pEftywriI3J4ikmU3wGxLb
a+Iwksc3kjc4FhlQkZvrH3iyjVbzhqorQEV1ACQ2ezjUZdwJcCFJYKBA9VaagHj1rL1BAYKXG2qX
bPUB0UUDL7wtlKCgrJyLUcCWt9w5oAZ9zlZxfqkpb4LhvU/YHbw3ZaxiisZhMTo4EodhSD4SQUpo
ayfU4+3VS9zfbJtATIjwiWskzKCqFQjo8uoIAJZ29OLIVxLYsJ6uunYcgGm6Z1NrlCodyUjLrR9B
0zNvh2XdgcRdnCghMRiaOA8z7m4lVSFSfihF978y+7v4OnSAF9ee2VsTnWUJUBPijoOtOf1cnXjc
1NZBLdvsYAVEqnG60pXDL1SWkurpOXERcifQ01Pk9T6PWQ+QOeR5sIqLNHGLpvztSiarUJlxSzUQ
4NZFthJHe1MWlzvmFu03ntuCg7g2BoeGkwjxs+blr5tYwpIUj5rGp4KTIMqw+/Vss4xeOlH1+V5g
1e4nyl5r2IGAa4K9CaKft3ICKiodxTDfwyIQK4AjD+z2fB6pjy1t9hNZpn0cPwox7Nob72MwmCIi
gJXNNHKKUrEweHlJhx5rfEbGqwDhYH3wa65y0+JUFJJQGt6qgjPx0MuYbQCVXm2Ax8Af/6hnHqRi
jeCFAkKlLo70diU3CoJPGm0Zeld7+x9bUU+euaKtvImMptZeGj70IyiGYgspUPBnGiFsTBqflU30
OUtw/H8vRzAREcnTvQG9WgVq82TQ++F7haLTX6nz/arzqz7vehxDSeafymUp6NQc1eShm3ohIqoD
i0pmbRuW27KFrw0C4KGhyv+8wcoFk25SbBD6hpKvJP0svjhLkQjAn1L7Lz9JZ29jxMXtvOAi7pAA
E41nndFOv7SsppO+6lAOPAx9hPek2OwGObGD0LDQHlVU+aShEqxPlCJSBv2Y1g3iO03lW0bt+UHv
XV/kVzDwmBAHtbsf2gl0cuxHZ2Ci3qvITRSZi+7/k2i4xQ+8VPL9aIVlNZQ/1w3grcKmjjPFUi9Z
Q22jMaNqp+QIATe3/72I7PXWOrV83cuLVxWmamnUYMGO4fCtyjPIV3UhXXl3htUtey3LsHbFNjiz
9aBbq2umyFrUUPwdHpGL+GAA8nMRQwMv07WWnxqH7EWNYWfzurEeJmFdG2JXDRegRt4v6AA3yMAw
9rpKsTylkFDrt9Kngxj/+1VNM2BYgCEKVrJfKAmyjrE1+Cr/BwxziIuJhds6WI8SjruSq75CVLSE
gKMp7opdOZzYaB/k6xn7ZCWSORVVey6ZncZQoikJm29RWI/IK6InkBNYmXxPlh3PWhxbswWt9oou
1JMMMHfunsJmbLPk0KTDji6Y9tPbel2k50zuT6CqnbemoLRED+HbmKG3QjL5x12b3D05J43zbgks
nt+eT3XwM3t1TV/yXnTF+7/OJ6MUwWgghl95bd8MZ2xyX4HGE1fN1PsblZOxUnAMb6R23hfg/O2J
351H0tM8Odfnh6w2Oh8CoOQ2MKJmn7whURvQwmkLS8V8ftzAxKZK+OmwCBwZr/p5BJ/uokVVe4k0
qWQIdXK4aOAogkJXG3v6UdsHbQ+l7XWBbbELuuw1VXM6VaKGHpJQid9h+5r+QZqUBFqXnPDI6qmS
Jt+3cOivR5w06dbxs1766rK7UyKY1XoovR+rfdCcBqH/TwtzOhseUPSKTkhEnVF41X9k9ykg7U66
mWCnYoiX2rb712uoD92x/AOnJaXSDv8WjQrGnTsLV5W2LEXyjJdNZkRMCK0KLubKFNLX8bMA0elP
yFJ+S4jUZC6Mea5FOGbfROLml9uN1Pr/fXGb/Fs49Y/va6gq9qNaFmNw4OYnt0TfikR6tmmSq/uc
lrkzHKpnEEUlrA4JWVN6ESD7h5znFbb6I3bEMCcaF6XLtx8wBiC/f6l5ALW15qLXP2N14S5JUBM0
rX67lFHhEYkzid2hp3Irlv8Kv6FpRSaze3Yj7laaRXbFU3f3lNEXaE4ANa3Q3hozR+aD63a+oEJm
u6cmNf7H5FDa1rY6EUc8BG++vC1gBpJ3nxUzqdkuuxM4aQa0GmWbTxR27eoz8yX1hOS7tlPH424s
ti+Fzj3Q+NqNdk6kKVztcJpX5YQ6OlCvkCEtDbV20SQAO5VkRQxTbWnzursN0Jtj/m4lqfnUObUo
1Yi0zG8ufWqBIJHaUn21OBpK5eBs+4+YdW0afnsJBUDCAJrDbGDdHqG+Wa5viMqh4TPkM1nUADmx
bMb2PkBrGXzFQ2GsCN7M6vrrDLS0NxeQlT4arPY+44E6bumuvaiPjrnQrFkV4vObzzcxHKLq8zv9
gz6oFbT1TXVEr3W+fMlpVllWbhwi+qDBQoflhXG2eUrWFq29/T1Y5TFSXp8sbHAnc/htfxOfIqIZ
GOTh1kuQcpYYRxlETrMRXvHc5eNC+DhcVqsit6Bih6bXFQREopfd9upWswcbeNRfQlvQzIQIJCAy
u4gZldxKhBq9kkwzhaUhqi6lESTchlVLzem3+TDZTmGce+ftcgkbHiZBhnX04XzQOXLY0XMGD9Xq
SiX+aGyKhlUSvCHO1rc0Jh1Td9053fDGwBNx9ZPbJxHN5G7A3hH0GUwqS2MRGgLQ6hjPAO3L6R2G
Pr81MfYnarFnmIbI5px1i5kjgaEPsjnqq91s+WOB4+7mPfCGP+ppSzrEJHjdxt4miQyloXhs9bBa
tWYFW3k56j/ASaqLLtpQB3S/Ratu1xLpCCK5gCBEVAFFNpg5vZA2UWaQFVAOnJ4w7TQPQp9GxHt7
ozStHp5Flf5HcqabO5sGkpr5j2T+a3av6EtvDsPfmGCBcc4YH7POCXz0mbm7WdXNEIjqmvAJzZaa
CMsxQJ90qdFefhUQpkO3x6GZaQjR7Vz7jfpiAzkjnJKf4zXftLdbKirVPaTWMuyjaAdLD79NpcMj
nL8G3BILrrruBftKD3bdFsspcqpdYnSfkifjGqhZFTXeNF19CaM4vnXAMJS+aX/kfyV1VC9gACdk
DxJ2mvSr9EMLEInzsy/fxJ16nN82DtAneRcy7gtFn33ep1FVBbHvBIqEGR/jiKWFzLe9JJ4lKYhB
OuSK1tar/E9JdOoVnHXrT4xx1/F/+XVeUjyo8KjNzGqnAD+uBQAYBndlv1eKde68RD3Yzuy/4BXi
syUlsa7l7YTyDuGE8Qjwmxv6uw8XyXI+srO308O5TizXJPRaAAgL/btbLjgXNgnmkNBhEgkflIe7
HW6xnlncsuT7D0Uv6Mqxdogcy0m6be4E0BRYUfm7Fvfulioi+GbLGuSOixs673UXfI7qN7q1IP1m
r5yUVSvyXUEWwJ39n5tvSVuJ30b3SndXmAEhKqpW3h+eBhh+92V59qzqD7V2WXyeh4iy6lVfFIrL
ZUIOeb8uUIzr0YPKNo/KnQAzYdkkn3iOvSKUsLw8NvQPWiNkSM+tmc01aTi3QfmA8BBEUA0TVGQk
fyMN8P2FnEO1rEmRolI5TXLeu2hSoxdsdblTjJ7NtBS7BBxLj9UhWDnFdWcsp8VyYWz1//b0KbPe
fKEfzZHjNuO1syhSjuQ++kpeO4v/2l44g/JWzSZMvKA8N0jMvGCGkO+OYTs8vvlCFWnK/3BtGfdj
xypHsT2mAnsUD6B2XdMEhnpTF6cekPcdR3UycWLAl6xkrPDfKP4mP+iaW3mZxsMfcs0ewwjTTVNm
hRXNizPEdsOGTIUB+39zXjtfEydDbwblXeffSnvemNKSC6XejQV5QLp2n8XQcDoGUHP/mXRJec8W
4bS8iBSfRjdTNwrg75WD+16UflLLNOhE30uyZI4+rZC8H3lK/LcNp5fAbwVlSecJv8Sp4GTwNTK2
vlDLxx4shO5vVjGF81/3bO1I+f//AnlBNgJRlsxGYzJhpaKbkdHI4G09NIn8jO814PizB/a1uDcg
meCILBs2XE62p31hzHHg0PX7SFde6Gm1X3HNvPyAh3MJTWy8jyUgvLCE0EAAQTiKz/JUUL83Uhqh
qEa5YE2mqwYnL202OM+vvtkBiUtsnVVdpleApzKYRR5WLVGwLP7TzIckbVoXyixp1SjxHgHXKtTx
g68uleNDFSEdxPDMlCXgt41rCAeDIT6z6Wg4/q/pTv+OFGHHeDwZsv+n3nUjNJpnlqIB9bWhVNrj
JDzb/Zwy02+aS+qClwmQgAX4UxSfP/XZ24tzXLq9dNB+EqxzToyQ+XtvvSEjph5+SZiqEEJHqVNT
7F6wQc9SNfU3drHClbmyQ84AQY3Ca2Js9UQKR0hqxJk+zc7sL1H0cPyzeU4+B63F8kCOn4ldjtDg
ylHIoX59gEIvJgKDvbcMm+Gi5rILdliPKhbKu669+xbOWSZ8HteecvT1xFUPEeEnwnyJlXILWOuQ
XYsPjkirPfZV+3aQlrmZkp4qaJYeHSqnQiLdFkD0R06lES5BmYZ/ISIXcUhG5NAt8XBLgwSlg3G+
wtIXcrSDfZ98LddyCgWhHmYFwo6kxhLzDhZ5UJQ4EeYLuDzIu8j9vyamOlXbhqJqjy4FRHfVMtJw
XDyzHsJJLNG9/pixDyN5ID4s0uZ5y1NWz6/NmO0ZgqptsJIDRqBueVPwO1OTlfI4YQ0yBEFcjuwr
XsIJ4wmMEILWNiwU/UxCLtXxujaGROeZnhQ8N27H46KOGJKwtzDaTwuK2TDt/tBrM//fXSOczfs6
P/9sC3B7CGCpNluxV6FPGxVvUxjLOWEMb5L374dEL2tXY12xE704ycXRYELuePnBrmVFyKeUmjjs
lskzmXyh6LLJl0ttRBwedn2sABnhPCp0fFSjm1syS5OUcvZCHPDbnD781iZSYR3GePGnECjj1LDU
gEElt/sClQRfJU2puL55Jn/mluKtFbPmOzvVjmNGx0RuiuuPHNIQOb9+nIFuEzgcTfte6MGhuPa7
T1WyUOQ8GRKViZ8/XjNNSgwHMaeXPKXeNL5YnMqxa5Po55IIPbiVoniIX92Xs87zR1Aoh2VTGnaA
G3tbn5CMSA3GNbGSz4zPWHNqYrnhLQRKOpHHgl19q6nkGDGxdFa1ChBz75uuF9rz6Ub3QfrdwI5a
ECMBpjoCjq5IgFo80R+5vFagrbKl56cuz2Jmm8g0BH9g8umRqrbvegum2S4zEsH+05DpUPi//6ZU
tDpLKPVsWpeNJMjGIX42dwVvMaRKPY7ash1PZoBfdY96Q0HUahXxP4pFDvBYHnhMgm5a3l0WyVUT
1gRKfrD6gEYrqV3jnk4/xzAuBl3d8SPPJGMD5yXe62sBq4QYbsDjijUnRFI8o4zj3Es0k+jeEE1c
zISj8S2MkTkY5z6MlQvMF2YdN/BSlu8WeYk90qGqGYSw4A45f2O0A7WnfQn1RFhdSr0y8QfDgBRs
fOjSTRKWNTJj1wy9rJS4BlCKaTNVEvG/l/G0nphGed0Cl7DdcLanonUuX/c60G7OQ05R+zc7YNM7
KbU+VEC4eJ3J537dsnCMTR/phh9xVSt+aj/EiQeYGF7PNdVx9ORcaw2/y3BKhSZRlbswttY16nPj
JV6mak+/UrGg9vP3CpSYkKub2t4j0dA6ltMuOGS+qZ/P31WytQGAs4vo48XEmUkCcY0TomXARWGX
Sg4G7pgMiCnqVQGPmGFqzH+WGxLfjlhoEYIq+3kRi/zhWJBarP9Un/4hSCFfKTQQzQ/JLGwme65m
X9HYhygTzUHajlmDRdhFk3ZeEd22dx3p8pd19hexpyKDvoCdazNXzOuoI6Eee2ZpuROUJo+OmRoV
K6X+Xqp30+hfvsB5r5k1/Mv99A7zrwFlXlawBgSThjPJu1X4IJiCJ9trVaa3nLFavdTtLL7CsSNV
SOH3j8deEes8JcqsHIWoELg69TVbuVKrlXFmwOtEoeMLwtyNlNDWdxDC84Qsc5m5+Py3q4ZeCXmS
jzAhR5ce5QbzQbm1tObi4dVeBIES4vVU7Dpb08TSfc3VpQwzYXDdUxMjuH2OLoUARWaLwYDc7ftW
oOpUKYKA9GFAhhPExmpj+wKrXWJbdTjTaKnVZ9cHut33MIiFIxfbbmKy5DaAhe0Dx7TCUxFFikRB
Vnm3IaNwUH9SUxLJr3pj6pAkCZsiBaSd843PjfbdpZLmfV8fKkO8WDZLuedOIgWfXbp4DA8MPBbT
/WOk/lTSJitcqNB3CSW7lXqHGE/G3AMPRiqeiqP5UnlNL84y/uvWqbyjNFr/f8O+WxwWRdG4rvsV
n+sSVaT+xjjfLzuUvxI3W7+dgywC+xlt5twninM9wVO98nPi8Xf16aClDjvUvIugpOlqnms5t9cG
XozKkqe6ZZruCjQHVUX5Ut3bo/qFiInhjWvFuxExl5sw5y7aqjnP/seWBpZZjj79tfCK0KpBsw3x
o1xVWInnyxk7gjNpu5ipQVR3/7+LIrBJuw/g6Pm9Ll0vy/KQNx2IhZNQ3b+ZhOPJsdtuZgecH59W
Da7vwHM2Ep4P2pd90zsJ2MOJtqyza5pZt16qRLyGTaWRYaCE23ipsscNC/HmbSK8G1MhWgFhaeWG
ZMFJNEKSW86nzaIsnYZej7QnQ90xqngYdI5bH7AtUeP0f/YOPKySeL9gKgHyQKIErXtKJn1PSTYV
y1XufgEOV7V7oiqaWddTdzBN11ZTd9YoFkD829EexQScS8HCNKzMLBW8EEI11RZ53oYV+v+Kc7MM
sL+thn8pXBd3wPe3rMATwXcNp/LvAzGdXCk3OF+geQfzf+UF1abdeuw95T3ShH5vLG+QeDtf/I7N
M2QP2804tUc1W1vLuMHXGB3zHUABX2+ijJ+DhvywrDB9MVjxD8AfqtXPZ4mgqaky54XnpVUP01vM
pyiAj44AuQcTsj32Dh//pHAFOEWzfW4aTI5kAACmgG4MUrLza7GIjWYZhgZNCs99g1lz/qxehTGQ
NzhlyMCj04ZQiqsJQ+SKUWPjwCWSdR3ywjKYcKnVRp6fHfBPHf3Y8X9p0RC46zV/TkwYGaN0c3oS
ZASYFGUkhKPk8W/Qza5rSJKJ1W16AZ1X5MG7kZJ/GtwA51MBL1G/jnjiONMQk6Fxbp9KM8AOG8vi
u4B6xsxjO96026ZKQ9PmBrArlLzrTTV77PU6n5aTGNiHzBbHqrZz4aEyMNolNuQkgXaAkXGLIITQ
PR7/WzEejZoR9yBUbsrHjsL1/6qIGeEAQzWE9mBgMLXP18/CMJWU+xPXzhO+Frnz/wNhKfOzNpxq
N4cwwlvvcAs/7qGwxaL4RFT19/F3zGCQ8+srhfgQHvFpg9u5OwpCmTTgHY9lDjJVjXGLywSctEg1
QSAwAmIDwRUj8mQRDS0VANV0E9QJjHbndmc9IQLJKu5WOpQIRDnOX4j3zC7H+5RTQ4bSTwzIzjMv
ngKfzN4BrKnp1HSyiYYLQAv9xnREerToBQhz3h/kEu4lH1Byplq4KOkrMVF90fFhhEU0fr9KBoib
tTZrMhLPJK/tem65PRlCG/SrZwMXOzfbUxNmZ7rknj2SD8prBcOMWIhfSpnwV0GKBpmTWUi/goAC
LVT6DAm7x58/KQcQVypkzc33DK1BtviGsLe/GRYW3BLUZxpBPT3mAT9UaMAxUayOY7Ulk6/U5KHb
dSNnaJH0K7O6FiajDPdMTd6FN/XF9Dq35aY3wAuLyCxJ9atVp7VhhwSTp1+0HtpD/NhLyr6nxOYQ
oepbynO8rtiBoxECu7g8F07EypCtx4Ptf0qjGGnqF0kRPTntwgF/0jlo7QbZPCMUq7VveY0rckQc
EmLY7IDLWDjQGQylyosOALsyucTUKQo/72hqJ1glHy9TOa085DA/f8qPejVmgKA5CxuWcO37gOIK
ZG76UaQy8vCOwuFHZqoay8Xs13swk3liZ5cz2ST82aedGiZ4iRk7i8ersaMbTJ/grjSxKqaZytfD
UvrR1YafdKfgxkuA8F5ntWcEXWdeeoG8lCUjuVOK9DRUdJ6rCkrBktvJ/x7q/M1ekovvirHmdp3U
f83JemdKAE9hoT7SIJyb7xBwY8HlfKmnsv98mmr4vZZw7+mhF5lzPXA6t/g//Ps4MX8yJx4gmVtU
PUBMTMycefbun8WOn6yftIeH+ZgZe86q9Q8ZgkBq6aIwl2gAX9bQ2/w/QxcJ5w/KsCzG24COS6Op
NgRoF7OxFleGaCDfUjz2/g+YBjKWCRuDHnmSSfKF4FH8hvhBOWFHs7sMFb3DsP18TTvR04q0woea
/lzNfscM+Rt7Xfy8vfo7etfdN6vWM0kbMuFeowcQ0bfS8ZyD53w+cTxcuLixeU3CdsNhNHBN5xJR
DkL5XaXHwJLq5CmiFdhSgftXHQP01ffpzay6NbCqPc99fhddxRsgcOgzLkW+1jBVJ8hAG+peMJeG
Bpd55i4lW7V4OPWo6ijgwZJPFpjcVRtJsXYxPl1/REGF8/IgH3ZYmN7KVEDJIkMhggQU62hI7ZKZ
bw8IqRIPP2mPhEQBsbtEAJO5GSNITePDjkZDAX8f7GFoK+4gN10IEihM/XEcP+l4JzgOTW6YZvDK
0+i3OM1eHXoQTnP3qJ4yG0Hzwq3OMGohAIkP0thXglCc82bV3n8CaM2b3YoMoktLVIZ1dRT8z7ej
WQRRGntt1C78rhdlckUoiZL+3RXn3oZ9HKBcphTwEbuOvKaoZeniiMt04JzZ5a/0oLRHaCXeGOPm
9WDuG+1TxJ6NbnrTSbwmV79Dx7utlcBocjjjpmijF+YbaBOxzPQKnazf1e4VsKSLCPzB4TpmkSgG
QaYh4zFFgbrBuwi9JZoEqJ+LMMW0sBC6S4f+RqQhs6AkamR0W1CdP1FUO4LHsBXbF/4Ovl8X2Pvx
15YbsnoL8ZUOfXtaJmNlsHKGkP9mrbYTZjUqM/83/UKzEOsM62L0/KKWnn9PnreNwmtUzU5lOPNR
sjDzWZxjmuKZVAslY02Qz2Ej3AtR6wFvlSYS0P7E+q4ftFD8v9ATsgC4ZevJmSCCq0qwFzJbaUbL
YHaQEotm29pSJY1+zYOQWqTRf5V1z9c0bE6BefMseDVrV6OAD4By73YiVg1IEIRTGpA3yNdvqEOP
7DP8rAN16FKmFaVLmHud8h5RtnW6sxOJwr3ojRcFGaTLSjEFNglCoPDxCIFdmEC+WU2PUTdi/MZS
Cj6onLSyS5AdXPyRtUspEsP6YzkoejA1AQ1+B3GvRmoWfYvyyPNWyj7Ik2eGfZAuV2d6QZpUzk12
O6vMOSIVqfHVJdQssqPBDWBSlrE28vO3aYGpMem6HdjGaaf4Y98sacqIgGJU4IyivCo3/nET05CN
25juq2q7HGd85kMC92pYhxLW6WkiFMK5fBDBS+aeDTvOwArNEJVtS+vTBVLboPqdhjnBTm/ALyDi
rOR9Hr/57Kv7+AjUI9D4Eq47zJ04aF8dakQDG673Mi0Ltsv6LhqPlk0+9KXb+j4anfA6rnLn7DNP
H722OBXxae166rOGvOnR51c7LPVwexqkn19tPgo4B2IzlDnJtRw03LPLwRTWZXvfjN+PSo++6T/A
yz1W8NTvOJu+XNJpKpU8FPuR0iaNqEeVOimAW3rQIL/2QKZaMJjYD+9YEjm0uvclj5u2z2xAxZHH
7c9JYD9JgQJmPQt/Qa1FUATV9xyAQSnQiXA7isODAU0oZTZLVwzbcGXb4g2cMJ/KmCJS/wst1hC5
OURHOmwyXIACqQJbwolTGfqbXr1lLEV8uS40YeZnwfX3mmfrInZkpRPg/UfR+4DhJCtHlTRPd67a
UjQIRrjpNMMmnmqMDQdH9iUz8UQI1WXYl9I/DT6K+L5dcJh+TOmPldmu+a/EukSn5WbUkpEXQqzz
v2aqGYe3OfJg6bV1muOSJrqgK5kxdPuUfZ8mIRB6M6iiMA8FkwfU7WtNZGJgTB6qftedprYqqIuY
nGrStUMGf2WR5lpPIgh51gD9HnScKjqyMuP6PgGgh95BcCazAnJ43Hb5RG8f8OSM+AvWqNSBnW/4
59aTm3OZi6gFs502mV31/UZdXBl8olujuf7Ze+54qCeNDQTteYmcPTYftLnOoglpJHdXoH8KezAJ
6S9uBCQihpN/jXUlTTU8qYcHUCjo/f5fQWWPiHA6ypDyVBfpBM7IZC1Cw2uJI+GoxNUpLK9Q2XD/
tkAUCVTOgSg9cnKHrynlklqV4Z13D5y1qzxq5TYIJKz+tK8blL87HgMDHnB7pSLEKqXwScBZI8YK
1l4WPHfxX+qe+x257nkY8L8Z1J+/oF1BTKIgtI0oLNDRVCuhBruh7gYq40bUygw4F0ok8xhADkWs
HIIiypIFrxk+nUy7adXRQajmLo6wLRRhHA+wS4nA1QkduxD9obs4JK2YgIfTo/2TgVBFmZGeN+oI
HdKLomipxOCGTXEJM8MH34HDiU51Qu96aFoK1vjy4mGWxxfyuecvVxdgDRwWtHaCt9r12Z2seD9h
DyQBC6GZBSmaouOPwelNFhBCLqmCA705EjLducn8VpUytIKBxF0/bleXES/U5mPyuFERmA8+qjjG
7ccLCp5sVfH/j4PWXb918XZ8iB0lC3uZTiFb9wT5CakhMdxQ3vrpBwj+DFT44DusUTEahxxInMLN
BD1GNu5Xxn1sHZRAmtro+7qA8DQhsPsOdBGtKDKd4LjGEOVqejLhiwjCj3qH4ZByJ1DvXDSabPhY
lLWy8TiBXeF7oelVBF48dOoCpxU7JBaO8ElFhrJTwkB5HdHmPOMBo4yQUtIjmzCr9GsmOWw9JONV
Da2wq2bkkfUUtchqIWOb5SxW2q5X5ZtHbgpoJbLEsLFhW8WqUge5vk6tblFTLedUAARZlhRtVCRN
GbpjcwzuzaJLCfzA4oaraxW4+CnrFQTtyhMxdsT6eSXv89uqMppDWfp5TV1IcxEWLWfCN3C2ouTo
9Q684JkDUcrkUqrIwbarpIbFwmfq8HcFM6tQEC16Z25BhYFpaaLft6fO7cPXsopoLCBVuUCoeg/i
O4G1RmXJBXhl8u9xwMMoEWmGLrtrJ9b44qx3o2FxNwbzK/xe2mbJFDYsm07oXnanvULIgLbhhxgE
CAO2HWjXXXpFWN/UqsvRs59DSuo5YATq0cpsg32e6ll8YaED6icMXRPwysZkzoIQSsXEFT5Vw8KY
vpWZN3HQPielE8kucGcM8Wsv4oomEjZQwnmbpzSHbFJUJGmRpoMjpSd6ucjFJ7nqdEjLAiLUd3pF
Pj4OxkE+N8ef3pkE5379pMLczChXuNfrQ22QIuZwWXSPcXukm6JDIooZnZRP3RDSfqv2GaL/PUxg
u9owGIJbJbJBZpiV4dElv5sGp1EvhApiXXK2kDK7XacKoqvR/lpudcpKQw70MCoDAPeCE+sPrhFv
m0KrpUb52b5wdWWGUzre+0TBiYvgLgLprVGJZZSxxcdd6H7KR406T6iXx8RFHA19D1X4eLwgew2R
lkxeX6Dj3efUjCzzidoppyl9nuEGJ+lyf71NPSD/4+hm8DPXNDMjvgyuoPEH2lyWfZN/eIwHJPj0
qkM4NuXv8B2IKP+JcPHYEidLl6z1SekZxasPlD34hJ4k0ZyLHRPPt9gxQ28CrmTcsFUCXRxioDmn
/lkEnuLGFL6RmYk+RON+OqeM4jhFfmXiHSfQ4BPugjH+3uRUV4PVtKFAsJ22IXMPqMX5NBxED5qo
LB/MhRM7ZT0Tj8r/NTcEFNzba4EH718I2vp80yQ0EpGuC309iiEkviSzHvOc5EKnJZbwGhCeZTHS
CkH4pzoKMtXCxSBvqe5rLttEnoK2JTXq/d+n4sBE6E26C4tcu6KOjXJKatYBf5O+Rc+vJs2FPxlS
vjKWMvyz5Z48MA41m8Xtb8+vRAv2qeeHjUN7hdbzFDXYnBbKQM5SrvnmS+ovrYUIREqKjjeaaXC5
sERsNt4x5G3pPSKo9DMPdsUVRFFAFZNzPLBxj1Y4P3jYDtXWtGe06UCzxYdH4gzqNbaqbLTxikSu
afsP6uhvXh5SkwJcw5czqGWiH6yZ7GN4SC9rXotWPF+eRWvifX1Znr02W3a/mJw00KS1TL5MaUTj
f34+1qEV3rzD7DxLPK32uKG3jjDwfh51Bfwj/KCu41xnMZ2+0ff2beVK4jWhvxMapmcUGuuKOQz3
CJPu8cMdhU1FkgHkg8L0PFI+eBRQTvo6+WIx/S+HuSrd6qfH1hLV6eA8S/1v5YRJc7l2yukmhzmg
e9OmUv5T6jEsxfYte3THBwUtWy7DSfFi3EuB8u5DgM33cQYQ9dXK07ALvn4ycBCAqQ27+ZGBExDe
tAOInpPKgahnHzws4pZOKz9ubORvrweq+xBBu7NAMJ9Tw8Avcru+GKSZVUDYkTqpokXaJ9SqLS75
xSRkyxTmq+uXXFp2/FiAwq0LMLT6jun/dQ7CCD7BMzqYmQM/yFONUcu3OhQjnIyL8wAzwMccpbxF
DDclLQdKEHClPNqKCZh4j1EjwlrgjuVfnRS3/ZIFv/n0I/VP2DWHHsaReb/GEW13M827WcsoS3/W
34+7kcujRvw2V+Fh66MsXUlh2mCygiZhyEBDkA8BgAugQv3mKFXA8PHTTzoPfrgDl5DX5kT/pNx8
OebFbmQ/Itd2JYPabRBJ/dgG4GW7Q7+r0m+4EMy9mv5shfpqGPVMCs+4krLjAuzWIFPtIAkbBJxU
GasSUus7lCGc/c4ltFTVzumzd0o8xMVxLU9K3y1sx7RUlnFEzj31SAiZxRD98cLJ9wKcu2y+ZziP
SHcdo8bbAK5I5t9RnebZ0zKexzECXF2dBqJWCMMmjoasYYxTjEOomSjj8jlouEbL89OJEqF545rx
bWWOq3kas4giSZ/RzMK6RZJpSPlpYUrDznRLKpzNepA8jD5oOx9iecYnhAIaHdUFIRne17PlBkW5
miv8F0Yu+nvJK/WXRMapwaHpga6QTLiSn/gXqwkCsz+QBnWU89/WT8s+WnaLptxdENFSRmLorlFP
O0omPJtdEB6TYvLH0xafkLGrx1ALD1r34Wiu2dva6M/OujPxpnexScGD1iBS7cybueqoWZ6pfqtw
dkv502wUQgnPTIekU2zTLR6Q/KqVTk7Rj5nu0grl0ZxWb4T3+3JTPqAxKqAM18cjO6hX914v6W+K
Grn6igwM4gAjuThyVy2kUqgoqxnjkoVM1fMhO7OxZo3T+vXujsozM3l8D/ikx1NX26b5QjGcUnbG
bo0cNl4nx9lQK34Dn0Oe5Xe3LsIW1v50zMcWC97Qvejee77s2/C8jVU/yi0SsBM0uCQwqjz+0mQF
IHjGBluXloYHwmnJdaOAhKTzFAU+JalMkKWMnnql/qCyFHjAqMeuSoUe/Q9ioLqys6IC5vge3g1u
jHa0sBRAoJ6opbXkUHnVIyQnNEUi8XH0bBVNfq4cKiRWh334eyCaXuh+iwjGMX/o4+s7jMuHrXxa
Nh8TG8AXhbSV0zJNDRYfeFhu8iMnnFkWR6Q+NHEwpZNcYqzqRTXvDaJyLntEIegDv/mAUPmcGrzF
j++MlosZRDYcCIimaXZLChRR0as7j0BXAMvFERHNbN5xAj4z6287fzEJ/ZE0mxfaIDeJ17i8Rx/J
1sgKbIPAr+Yz6QZ/G1ksU9ivxZmQQQFm7sDevVE1as06f4kfqwfTI0L1fZQD8evuOnO2UZDrsFKo
FuhV3ZkuIIJevwC9UvBcJj8pD/SaecxXo6MVJu0iMBmwPuGKTiizwTKKP7OkSKzPTJsDQ+U99zVc
xebClyzrqrJ6G2jMUcbCKqcEhibjkvcSHuUwapJBY5Kk2b2jAvZJ6VyQW1fKB5Sk5SHjBNM03yVi
2W72L56G63PwRGAcLuu0gqShO/ZWABZSDQnjgoDLwEBZ8jDg3nNjI8C7lulHhrXPGNQ7kiSfihpH
SSUeZIw0iqVloduG4ZIth/eK0iApGiI8o1+zGoPuxJwe9nJclX73JXa1NGtCxA65H9uvjYTfQd4i
0oHUhCroJPRu/ISerIwaOkPpPMiL29eHHjYaFBhpncjtCwVP9+EVY+RuDzU2DpsZA/HkEdsof7hW
7PPRJqNhdZXxXWWah8+sD0pYwXfs3WQT2TAcSrSU7vb0l+SWQOweftMQga68NgPKuvVCZKM9ACW0
Vg9MPV/MUcF0lajntSDdYB7bSpDm9ZvqBYUCYbWh3bEmMVsL11iGSRygn0lcd/vsQbhPHy1HqNSR
zFLSaBtb9+FjVEdFstn6QzM9mqQY9D7VlevyhIii3FY40uJcSRDt45rJa88ppysZOcld2l9przxp
T8DzdPwo0KhuWku9DTuc6PcNeN05KKlRonalHLUD6swj3QtdFHmoi0z9hBZ337CwRJJEZOa0AnjR
TDOeF4VoY+t9gR6+/keoYriJ+niqgqzQRBYSKb2hCA8T9llYPMDrUIH/mnhoqhUCLCG7FmaPKn0m
odHFuCbVFixfxPtoDPTRXoflq2hoKpaO8BBqKL9lAOVXb4zgmazWZsf2J8DiGuHYB0+tOv5D76l1
692vYQ8L88715JQRt2/7Nm+ul6V6zlSYBYXzODC5tGxPfx4GH/Cm5rTnWrxF+V9Vzi98ta5/VULq
LjpRsxUWCRcgPCHmdA/nTZ6QZ2JePYWb11QZec+k7uy6zSteCqFFWdL1PFiCzndh4nmcx57GQ2TI
jfKV9M/mW34PAhnSYcLE+3YKl8ZJegwvjBQ2Qkesj6MBbHSJyEOMRHl56e8dR8e99xnZHjkhMCYF
osBr3sntn30jPUgEvhPENmgB+ub5ey0GpuHBcNgDwsWD6WGHiTRltRuwdjUO+k3bZT9Rx+hoQGSf
iKYmXlb3pJ4PhBvvWC+2dyb3uwBYirpbVTzp0KhyvAp2v+MM+MGBHHPIxuDHhVok9CW+EFc4taZv
h4Ld7XzpSn4mCAu9L/hIm2WTzJhwCfrcS87Sr/3nkV9ZaLKOLdcxObKJUTOZOBWrbZtIOImm/2d2
64hIG3QWicwAteSdgPSIYWEkizsrE2mRVvr9xndpioEf+dgVub3pt2UwWAZt+ELxZS+8b/eb9z2r
MVKOuBx55Eih1p3zC5ZolNGN5uEm0zQM0ZRgrSoLFDYYW9pFMcHWx04zFRwoFYaYSURzmHjHLRSx
soE1iVtGLye6oar0B1cOmzsKEaaH/eFlm2Pw0pURTuPYGEs7W1Zl7f4+J5EGpnAEXzeuIeWx0Qw/
ngaKLFHlh1SRya2KoF8KD+IaCaZKzJmOhGdSqgcRWE1n0vLRx2xmwl6JwPxg1pVPKiVW1WH5QGIC
NUHdDNfOSpYbjFbMxU6W9T1RggzdkciSobBrOEzfalvqVbHQQ7SCzNHAkMK9rQfm2bek/uQLLL8h
V6lqxuGdt+CUJVRQO/+42NimGoyQ79JZqnkXZlXfpRSPR9X0YjdLbsPtdyuW22wlnJ9bFaf7QKvo
1gD62Ar5eABuD9pVvSxCfa7fTQi7UreudLAIV4g8KNJPmEoHe/zXSGzn9TT1CKQdzSjP8+JdnbKv
h2FuFkYTqrrJhIcNbCFc8j+0DzXdXt5OiAlQPbuMP1PSXaGiR84Q4/8WqAuGoRKV1n+1GLCDuMSL
2ZN853d6rxM5NJo27gHCWfqEpRDakZonUwsmbIE2gNxMmlFVNmYUdl34FVE03JSh/GXHmZQPTbdG
P+9Km5495AtcIgRi6PUCTdhIWf2O7hH8UuChzGBav11KiUEwR05FYbRl8SKQ1rVtB1NCNV9rXAGr
KPP7ryklHJ7KiCdMhbc8Y3etlRIyp41hBPnhqBt5I2ijqXbffPc8jA4R5l9MAaZIlqxptrDkmPtf
/XplrleLVCisQrEwc0bXz3UIJIdfJBj46bfTgHpAseoZlVjz0Sd3/Jq3ZerTMQxQYXrLy8IXV24w
Lx+P/KDZsUQgVH9skgOzhnuZM3f4BRBDVx1SY/usPcb2zUoJK6A9D4XUpAmM6IT+/I26UyTkcZLU
eaWuoZSYqXjsF9MEKhWstCQrfo8N1YAGRCfa/wFa6bced/4NT1VQIaff8zpeava6sjOdD+ga7ivO
Xlyim1+OJAqxSamX/LoTjpwh15V0A/dt9dVjN6pIVhAu6nuM51J0qmyV2gds9LXMnGCORgEPWMUd
En9hvQEkXLbvskjltQoeui+BdhGvIdGB4iryf8V4qlp7o1IdYWNxxYurgpcC4+opCMCTp/s0KOrR
5UqWOcTJcQuxgKz1dhgddcL83nfdV5bjgp4hOcHQDG5GU16nnCJQ63m+qpZOt/ZkKPnEjsAfLKfS
mCo7c2oQUBb4EC0kX7PiOkHSKoeVe78/72F5vSaGDLi0imghzo6efO1sOj+MdWOq9u1XTC87cl4a
umZF3bdOSb8BuxlRrVuJsXQeNiYhn2hecjcsxH6r7iTfKdAfrURx/II/oOk2qLJ2483ffpHJJU6Y
+jq5PLUwt5BivliqwyS02SrnDjZmewjHnxSybKGS57rOYwdEqqcH25l66SZTRKuPFIJUkS7QaqOn
yfQRCXf9JJxIglbLimw9eNJVAzJD/qcfDAs41uGGOiiNT2lYwz6tPA1wqfNadumW8DX/vFUVsqr4
QsENO8UrJMklsbv6ETI3W0MOtbry0WTQFI5Tnt9uz0FL2HaQqp9Bsnf4owJBL7rMS5auCvjUQ331
kylg/qySlJjXJ7BUfpppP9n2FKovkJpo/8Sf/1jEq6uSyX45x/Tmc5stpSfANS1e9RsRSENf2fJl
53AxE1P9dhDwJvoCyN8tVld1p04cF5/OlGvWTSbdb8NayTuCYwHNrJz508wwEGc8iyQfmVb0I8U8
NJY7VYa0teONza5cGhlGubRrJdISuUyqKTOC5vaGO/9X5O0ykyyxfwhEQcMiwQ1dFsIOP5bpKJ6G
8mw2ifMQ1veqVY2aUT+RRyTuo1nYlpo5zmh2GwNNGiR+r4g23wF2DISUVcQSTCaCt6F6qyMa2SNR
Z6dH6JzyltQSoWSuXd52hPV1GAgGRzPdyCmTTEt3YQB+BnfbmIzw47CTQvkhqDj7JPkrwJv5m1Rp
AvlGPhM59jIyABBfWRe9UTqhLbJGQFXHH/Ojd+i3ubi9B+k6DCMVunHwEZyN/UXZOKTuKsA35AHD
yJpGmi02JOloa5dabddhW7gTLC6i0AvEwoNvCXeee71TsOxUwCHhSLlFs06FpaTcvP+jyYs/GzcT
ruUCNCfw7BClX8WEOYe/VguK07bQzldIzG1rCUC6OSZKuskWKBwtVGd0JlUubVt5p74QUMjSwwst
uo90I4WbXkJl3v62tSH8Afqk7A8yHQrIE5xToCf70N2DBGMB9BlhSyN1dufAqe3h82MV3zezo7w4
l3s5abpps9bQr4qNMUyzGocae9fRYv3vpLk/mlf9gEP3guUEtYjlvo0udHtB1sh+YM7KrNvmTKJM
vIrGZ+wn8U+xmOeNBek6qJV1LSPMdSNqvcXoxzrzazAXfJsQhsvxCViPbPzOfqCBqBzkAuv+nd3X
IUOhm7d09s9h/gnCUocKoBnJzCQZv/35ZDDNlR7/4g4vnh/VAW+KZm5p6mDX0RPUt28DP/edURa9
pOir5LJ57dcyvoEqxozRk/TdsF4B3In+yTezcG4M8XlXn9tKD0JZ8U/4d27drl974OLXPHUU+ggH
mU14wmow7o9Lvopk1ViUiP+2XVyS947kTo7xfN1VssYdwSHMai8cgeluRDtUSPPq70JlKcAh7DtF
tQWJea4ftENgCi5oliaHmMFysny+iaSfS3mhHUeDkDyytu1tv5lviz9gB7CvqE47pk3G+HYOqHfx
F7Io3mqrGiGpgCDST3XHk9z92Ma36mj0W8wWdS3+p+3Ce5ez/AJNb2J13QuBCtqtzL8PCfbxq4dt
rjwHuwg1405ZUps8NgxbA7b+cKo099O5JhML7HxL56r11IwsZYTqhr90GM8XEMl/UGOeu8cylsAK
+3wbVBvjcZBK0L3e+6HZRrhjUcqmtQ5x/mSAUqm1e9gLqa2qpNI5f3kw6x1810Eem0AU4U5O99JZ
KETar7IG9BUmLH7NgoQ9o+ctmtkgud4Xfno/2HjtZ3i/V67zKtnxweS0omcFRgFgPOEBL8Uzh0f4
/3OEMpd8y1iEWn7zhXuYhUgl7y9g0RP28sJ2uIdCS4jEOWaalx3bY7+XL16Hl5DY4EFozHhoIa4i
2iYc6s85WicuXk4uHWpzQyQfqhZtFkaO9XwvKNQL7BZqc3+u/4epMXf5tNr68zYDtvzhFo9dySYj
Ncy2wWBT2hoChQqpp9nyRS5tyxCtmJbdVEoYYCoci4e8adfRjc9qpDPu0HrtnjZ+BLXQ3PEmD85u
xSUoAOVWe6wRmEYqxIMkvZXIrcTnifwQwOMXm+m/rBtbmycAtogNvKA9sBJe7X4skNiFRO/yta62
3+B36YlaRIWNFThsYeQadgtv2Q6P+y0Yit7b7Jb1d0SPwTr0/OP8OqbdUaSK4m3SYhnNYZGarmz8
9Xs5F3mzmJTh+nMroT2VF8Vwoz0G7DlbAuv7bD9lKDgrgPYspFADg0jxE4Jz9OLiEeJTz8CJyyS8
U5Dvtjfff5+HjGSr180LJCDJk83MZwnWhD6jXIR+S1ufpLHcOfRXVmJMC5fVKfpJtPa8O3ej3Ett
gvGYo2utvTvxEprI8/feTOMkZf2ehP9LCtr4Ai45kzx250/WfbQby/kkP2PnfIsYpvgZpmm71XZg
c3HY0dhzmrJa3VgWriMxZ7fPOnJCExIdIqqJjRxUoTfQmG8WmvUkLovr/dQM0VfNq6fZ/khWcGB0
+2ZuCVFaEnfy1FaiR0fV+l5I5N5KdTTSUTwENG8fFoX5w3yxJ64s90cFT8spCgsMxoUlh76F/SHz
x9KGXc47bbtrTDlqFZM47lKbJgDrUvD00bLA6Zfa8rrLCqvV7Ln5fG7ti6+meqMq/n96MU9Wmfua
9U40aBww1muDGZZV4toxUsvrC4g1WyRCHScPc+p+ttAa6XSlmZSIy3LW0w2aCvqB1C53Vz+PxqOx
66N+w2v+lMj+HuMKq+2Mb+MVdW1kNLH9Thma68YVowEMy9qvaP9yRFfQF8aeIlLdqQFIXIKcPPpi
wuphu7jaCd7aq5A6UkqFFxuZjGKkbiIB3sPTzVV44P61Jo4yZi/FmNtO+9Vfir7YRvHZcXFGvlfi
N7UenLMkLO3zl5uakC4JMKjhy0IU3aEn0MDDpsCfDWZLh+ezxN0nG4VX6yv6gi9GjZFWwGKPjVtY
tgBG93o2gDwUZxjJFlmuhSNjuqBf4EcN2ZQG5M8CFZ3637geRRYPc5Svi64Je8EGY5OXcnrj7Q9b
Ubxe4t7cVFJyKBic3yPBIZrCNVg+brDVEy9UM/aYxcsoaMEOtLag+8NjuyN0IA4hkRCXDw27MMH+
ZVsu8ANBjqt7RMht4Ah0rPj/nVkiWKHBCEu+xCeCMNyKHBylmHvWM/StRXL2+4qUSoKQELwTRN8s
rO6ggUm8f6aCk0fzdD8cpEA2tJcA42BsvUMNAC4u4obRY/NXUeF+3U+pIinhwlnaftJhHh3CelUb
UkuAY+qSQ9XMpTyNmAVzv2zmMMa69vmfzWeZrIcLrLUUF+mKgpipbkGy0pqQlS3V+tBbaO/RKlmd
zCuHsaiMyekmIX/3kGdcG3RMehWDbc7RIwnUw/l1W+7/THsbABazKNtTQmBVs91R5WnYjDVyOGbA
AUeKXaHQwyVrDSEFWCjeswaiF8YWtSHdTqPp3U31kYaNFZx6oVnsV2CVvkJPPb6DD/12FEk8FxeN
bp0uc1D+qaLLm1wIdp/fqC/3wN6gr3cV5nUuYVG+edXHbI83Vx1G2JugCPmJYG7zvcWcjcZWUyLb
oCU3fgoJh0LJh+9Ucu3GLqpIbOqaayYXAf+0aTGDHZktY41VbFazOKsMlWMDMAEbRCBmY98nnwgE
VblJQt//aADXzuq5lxcNG7H3EaDAeMa7cCSQpwcWJ8MKeMNVwALmzNFIAgIoA0WFYHkeIavGrHIE
Rdr2aGxxD4IQTxu8z3GEb/tidT2UBzQkZe4u/ZXEcq1MtzkJL3OUP7qTDaS7JlLNnM4q71zWG/2z
sxtGHbi/bTYK3Auw8s6GEmRiq0z6yYiGHFDyNeGdOfabywBxY8UtGhGV3LXK8hPXJmruKluC4NXw
w8rDwNNtXYJMt4CPdb2tmF3dW5jO85pRELbKuWUIiJQmlHXliw/5+bW4bsCLPS7npfcCsXhU1gh5
TM0bZNXqrA3D9QAmBM/PeWzMdaGbkZFFbb4yVhiJBNHVZ7LKV9GqaMxUSv6TvbxTGSRU/7EjqdrD
VIo26rV08GYdAnghVeXaf5ntieWPETezmOfgjT4LYr8kKAVF8TlUzTa8T3C+cOvt9b6joYMrCbOh
Ax1Bylz2c1ZUR35r+4wzsOYHD/4OSErwSf45AvRgCInO0aJgfTjxUOBDuMkuVgHK1z449Yh8P7cl
lbA8E8zSPai8M81y69de4oMAGrxrpgVmvQKlc1APTqVHP/eHAjQHuoLVaiwnRS5VypMU1padtLiG
bAZUSgR9dTgPN5NTbxbw8fOhrtCAhxgLSu1AihOuSjcquUNF+WXDEX7Vj4nzAGSOx0kInxgk6qLk
fCrhMk7WHetCeZ8TOrgHIWrXVELikivZUwBnP+o5ln1VHOBSG7KsyVC+alshDWlGROfHpSdKQ0QE
Otr8qENK7gsB5jroHvTQeWntPFK95/dtj5FV7FZvQvs96gPxvHk7E7suzYTBNSmi3zCOGxF4Td6m
bknE6C44rNttjgVSTYMDkmv9/oCYx5IgZGzypmNnSHeuslx4MsdHDKKoapDawveTOs4+AY8b4bCz
SdB6EvSZvoGQ2ZycDq44ZDs1XVZE6lTuJcJGWcYdNmiBxsK+jlrh5AqMfW8FNoiLWz8UCxmh9CLY
z6MR6fXsXkCbNUr3aj2wfCLRn885F7h7kZVKoMaD2zgLVTGra34XNvoZn1RlRpF2wsve1tsQkN+O
kdO8Jqgf3KDPO+rwDVpGNT4mJqEr5vSG/ISWP9qUuqmZ2Mvzqq/PlLY0CcCe+lAZhATzoGSsHZue
0ADLl5gvz2oquAfy7nm9M6vkgQyOAUHiOd5f32k5gP0sUHHNOa6YH1F7cXxL6DmU3rlsPeg6MFXm
CsVyvFGMBWxb4CZevFkCaOk1t7UrmS8M8VJQOZuw+PRV8IDrLYKOla5YPeDT807Dtqg5bvB4j+pN
r4JC3htiteCZPep12qm71yKE+Ij+l661b03lAgHqFJPVA1UTTwjCLTNNXuxA652DHwPt/pjdoWlx
rvUVV9dYFmWGozobbPIFviPH9NMkbw0LoLKItxpKZirGQMQULz52Am+BMROogmOnwHMMNxhbbWjT
m86mY9kYDDaBWoWUF+m0pELKr+N2B+cRph3uytWjsOljuQvgwguh4m1SHE3NGEpQxh1BLtokxwLw
zhyjPMphLZf+99k/BABh8G/kn3qPeZjyhzslTWtATYGsrxROxsi9gu5Ftn8xGVZzzfxEH9FLLEpb
EBQukBg1ZD7qZ5nHvxml22GCxJluu3U90dh5AyxCSFN+/4V31THp/XYY9snX0ydfHORZq0tdTHR3
+lE//otsBKhks+9wplGdPixM9+9+FcqfnRUKihiRdTmVftZD0iz6yb2V4HmGS9huFVhSV3AkQL/Z
AwnZSStLJYkvOKAtGHNHec0q+Ce/FPAtBM0OCGol9gDsYctYDWev2loY5kZSR3VzaOoNsr3ctT+Z
yAfFeZopm83p0/aMC4WcgLcdMwQwM8c5rIARXzO0tRYfGnlwlq0ho48sbGfl/LasZlINOOgZUVRs
LnVXxC0KE5fdmB/3zrEnU4aY5rr0GAAc+ajzlapFXvK47uqximskFihKJ3Q09/bhYEsMNFTJX2qm
+KvdR+NhFdBr+Xw25DTbAsj7PDc8w4s8I3vMKdxEp6mRH87YCML8bNwnk3N1WaLGZvUB5o87O59n
i7/yecg9scJR5G4eRMptE8IvgRAJQdmvSb6NFPNiqZslXRZktI7xQIo9DKeM6hbpY7qsWknQYDHM
NimlPq7hbPgLZAGgeTRiLl/kjP0ynLRcv0/eMw0Q62fYiDVasRWtdH/poGvfbPzLlpMqEpF5F3Jo
nA9RY2Q4SN9zioUPYYjIbYazQi4k15Omj7FG6gxmhrjVn8OKPb3uNp/2JJxDwLyeXFZHScI0YcYn
AH3qfx/HMrMpGELthA0yA6Y2fvKzOQfz9TF1LjEmifUreSRHthOqQZutWV95wNdUFej36TJUfk7i
4XadXMnVyjs0C4H49YVnZ5Mdon7o2Y3j5vlrC5f+PYHuLPZ2kxWjXKNFpzT0F6fQXlvtsaDplgLg
4aHlgcalIoWIDhx/ZZDrG9CowYF2Ja0dJE0QjuRTDQk1EG3o+vOdJbIxUe0DlZmnWUZCG63OccDX
8Yg73f0Cmsr+QPCnO1z2ZMauSmDVyu0v98rKk5yShmYBi1OuT+W+IsFBhC9vt6jBpH6wa1C3WjsT
lGW6jKh6s/Gq0M5e4ygvjCplVQWE82V+90UZ+znLE5XqNn6C6V+Hotmr5PUExN79FRpsyfBYHH2Q
vd0Oez2ditJ769Au4wK9dc1C075T3yRS7vIqXq6uPH2nwP0oySIhf1ww3oEc3SjqE0merxe+yJ5n
o2+oADHLy1icgbacQpWKQpz8zJzDzME5XGd+KHEQgbo3kqOB++NjkIppAFmaiKX4X3OkS6jrI0GN
oW0Krbjry1CMhSco61u/h3TZogluNP6b5qNJQObBNH2jZW8+umY7c7qOoPeCu3X1SQ4WqH7DppdK
RhcgudtXmLsBBgkEZGZKLyULOxpudyq2UwW9wOkxb7QSakbwxbvDbVxXGWgQIJ46Rc0uZcXS8+JN
mdSzHD/wYUzyRa6V769uI58D/mtNczvaDIexUDBwAMc5zRV7iU01ZcQXSrJNuv3IY81BcAGIxkYn
5sNcHYKdOBN1KxhctkSF68xit4ZhaaHunbDBLuYUKWf4PFd9zt8OYyxutEhSY6TTgdzWV3YXLGCD
72baaI2NBQgzDNeJzVuldjNxQzb8++WbhRjumUU/APZouo8/EoHYu/QnM5M9TST05hx79Q0vN6x4
v7/rotsHA2Kru+4t3ZmUEt+yNGiHbLa84TdMpNtFNDCPR+Yo4lJZHcQfdzhEjavEZieJn2SecpHD
00F+qXQ2aEhmrLz9yzMRQDTiwSK8kjKg4ppZcv2W5385kjRbbNKtwq4lVPbGCpPXTk8cSmgeSs/s
qmie+yOs3rYBVg7leH5Vz0nvwex7JHlrbLOpY1MGMi09vY61APFj1/RJhO4NdZh0Ae8079Odv7Y8
0rzW4LFT6TUMpSSM2P0golUmWMkvmblSpRqhjjDauppqRWx55bqzcmuGKZ3J4vC5HSbKUx9qHm0M
605s9p74mB8tvRFkMJeqf4nDGKWfwuoeqJskzDqkaHoilcxsNz/E3NHt79CLKhz3OIxsQLjV8DuK
4VPr8liy/fGOMb1l6a5MIIb/awgVBLBJUwSoVKcOtxyT7g4Z7+0pv7f51IxMs2ICqOz/ezxjKjIB
bRKz3mOjKYsQnt8aCP5/NaHtdE1QIncvzbD42jWkqZMdr6JsCct9ogEXnLrIFwMvBjmOWzN8HqD3
yzhorhSRyeDuKFu10iCon6CUBJ35zaWMZCi7iYSWyn2Rd/3QMZZjobcTDQ9PP9Bl4UE+pzf1v7Gb
W+jSiJwKS7tNRsXZE3wK2vCgaop8KI1vwY7RdVc5APTy8e1t+r9uNpzQG+0IK4MTkjIpTABKMscT
fLnqGPCG7C5bRcScjMxMXmLzwM3aT4jcOghrLsIs25jtvU9j4N3P+6Hvs5Hes7f93+pm8lzaTXf2
p1A3LoiWUv9QuzjWf5hxLkWEC7z3U0uoi6SqPvOXH6Ddn27Ini2ICarXbM9GXoCRpmK2CJV7psBb
MxXtWzP9Vumc+EVtAeutDkr/xUIjw+gQg7vuBChsfFb9S5smGp1jHX9P3B7GfedxNxyxNfLKFd5v
/ab++CVcVRUscrySVKi6jlq3nDhDusUbVj2ZJewMXIzdIwOaSvnxdfZhYc3oo+1pm7ZHR399LXBf
0o88Yj/l0TI+uYd9stqVYA3XwvFAKm7RFU9kRYrnl1VBv08gWdCopyap9IoXc3NKtYI+DM4mXFKx
XaLZwXw5Xqeliik6EK11G/jAkm0CYGfB+J7vboEHlPyxuo2rD9MdFghKeM5dur8eNtWRvPLK6X0i
/K/09knkegAV7iKsWAwpHDToRroUneaHls46wIBRSqmhATBrVQ5aTOfzlpDbRsFF3vC2BGidLwjf
Uh8QkASUJEypnDzf+X1FcjPMVNSCK/bg3hbEtwK0vswwtPKq3JqI4Ng/I9oX473iB8rDeXSBUJAT
GT6oIE4xTAOwx3g7e+zTYBqms3U2Ai+ZEJXh1KQa4VZsgYPIgfjB5yHGQiAVNMhTEm5ysszU1FrU
QX+Iv4k8DJpvea3UEj/3IbtsvNQrD3JBoymrzilDzCGk1fPXjzbctP1tSUTcf13x3j8F4lQQTy0U
otzJaG8TjOPP7Evh1sQDNCp5kDAu3g7v9zKtL6B7dtI6hgTfqh2UQ045f/LZovKx1YwuzpkU1Uxu
vkZgc9Ql8ieItZtep5Zk5iTR9+u77Y7HT6MbLaeuRu3tYVUafsey4CcWKJKV+tOB+nIAEIRWjHnz
4YYXK7AN+nAw9m7o8d+3ncyYfQQhWps2Gm/9kckEGi7liFZuTsvuODp3lQx+GDaOLyW2JPHbwYJ2
n3W35kL1c8MmZTn38pHbGwX7Y4kS1YawylZtdFVIZ37/rv8xhoOgn6Hyd915cWyI+xS3c+oYiDwO
qIucCteZcr7YMoHX/qpP27eJxJYNkIq2Dfl6hyezeUly2Eue7HHHWHBR45MRAmUQLIj4evD3oR5N
Pk96dihd6jJ1RLkftwt24WRLPhzGlxPM3lzoudi5frrwMwW3UskFUsITXM24yfN5ekx9LWyBI0Ew
iUqu5+UZy1H59rE2XYbZCTwJcVt7qk6bXHyH6vMZgUOFc9AyOEawSX6KenTkQgibArvWBvbtq1yy
jEHUqmtt/3F3BUo8EV878dl4fFcofTOXsSdBdcDK5M3vNMxLUcCzR/loiz4iY0Jw74SpJ3dDrE9a
NQIh9AE99dfXgn9RzCa4mmzd6UzycjTghFBhoCkEAkvCFogW3yDRAcYNQIn7xeB+Y/Mzzv9gABkx
7hFUtNg58BJpYvn9Pw5ARu887Y+9aSQkOx257uYjf0zW59Bblm2ht4VV3AH5pbPcIJNfOoiso7R9
Xxop78tav1B+6+Mdkzzl+vakvhQJOFPdDVmGMyCceGLrBu/oUGOHdmJimxxoD0XHnPhbHzkUvs90
Zn3G21g4FGHttXlu9kWfCv5qfAB+5tj3y/Dkhcsx4EgGPN3vJIW5G6DOw48Mi9DHZrIJEB+jeDHV
xkROo9pm46kC3TGncH65SI1Z6Tu2R4kAW40p3Xby3uEYN4DCVhAYgXGUsO/gOJGQtvzIYMmK7gJb
5YIqL1JaCrnKmBhilBNYy3hRqphK5YHwaREHOKKaP65JPIsECmE8d1bqq2a01qXWcNfXFiwymwGV
bfFu0hEKJaJqCNeKgRci8nkCuvaLlBdsWIgAvXNQU7IRzpJNb1HrLHA7HJut8TlfA5tk/f2auJJa
jDnxqU4OCJz5F1DNBWcqKSMswdP45WnBEwM/H/wsSlpnbBr6TWxYMRin7iidUreptwrbf+g/xrus
SfnhSYx2I1Q8d7QDMRgkUeYQpjZurCwrAM0JXCAu7hBGHRTFokQrsunosdKLnMwIsgjsUEPGm+3i
C6Ams21olG9/ht0r/izYnhf2EkVDtKgmjFBvUlg9RzGpiL7qdyLY+Ojz0a73+BOU7b+F+ALjZHC3
66Jk6jp8BeoDchVCPmDT1js+WvAprCLBe2F/cWwz04wlrICw6Q4MRslPkuHYXwZPOkVoQy6DLB2F
Eqs2igikTZANzQdKJ68PoU0XFurV6n6ParYi7Dj2BC8FNEnQCs7SLXS4e6F6ZiPnrg+WlXn5Ooyi
YeaKGLlz3QNHEQ/CxeeXrG277WBGSZ6NVA4JgtzDb3Y93TGECdKtaWdgn2IsSyer/fSVKG6hTaUa
BSCjFPLv+uNIdSy1EbK01NiUWw7p6Jru2h4qU6/ZuOx+kE1nm8ZWlEOkXmhdl2VQ8CVa0F3ENhhC
2X65q81bsGbzRamwuWFNflZPEL5Kesq9ePqXDYXUL2OrjC2tERfrhltrFtcw5WoGu1+c55cJRTUB
Fl09fkyzFbARVLW0Jz+SD8AsUfVH8cUAG6D8U6esEp1j/qZJ8vyZSbpnt2UDuoQr++b2BHCc7U/q
oq3B6UINrCkFd74k+QVihsuWAnqU1gCiE67EjJvUFbv8cjzIwcbrUJeOG0sUHY2HsISSY6PehYPt
oVCVj8OZfEnYpgU6r4wAtvAPwc3fzOhcwQCZwybLjf7mORiktoidZfnmmH9FxOl0VrSVPU22sJyO
MzbRsfvrTjtAiEi8H1KYfnmskV9HN/DSMpqm+JNjxiBAcc+d6OfW6udsmiUktuSt9OmauuUoQfpU
jFPnRcG3MwSTF+bXYAzAP7jJhbJ0gzar6ykCte9LX911RWOQ4RBuZvGLof7p3vTwq55eFR8S6+dz
13pn+yHvDc8NW4e3V6Dq5bDS2IgZcsoslq/SPuwmd988GkvP0tDfEMRd5URl+3dy048a9CqWN5QZ
2DWCAj/aAfff1XluzUpEoeQyWM3sN+UgVhNaEwuR+iHUkVuAtuJUjAHrxV2RPxci2ovT/fZEY1AE
jnzmKHs0TgcR99/CZSW98TZZgGXmkIkEKH/q/pF68lH3SFW4nu2Cv3C6OQkZCLypvBym8wY3LoMO
5pehKtIaLG7gn00CnyKlbkLYriShCKw0H2AtgeJaXozNXD+6nvGFhnwwdrXPn2fthO41vHK3+7kA
9EsbILxsuueNZxv6MBpsZjcfLG7bwIzadpexajunIIfK8EtlXxa6yv/i/n6Ne3SKlMWBxefOQ6sE
iiJJtS0sg5kMLPHhw8aUXPPPW6VvYa9Xz6l0+3q6rSOndy0hdvHxkm8FyycEfMTKmK/MSOFLcfEc
R9Qwt7CvZHN/8erNVyAEA52NBjG+5smhjaS2iu5Sbi94QDiv+a+XxxbFAPhealn8UJ05TqjVblwq
vu/RwOJ02dIqTlAuD+8oo+ljvSvU5xf9Cnl9+BwPWQgwdPtqGBN5xLqWavBM83aVCRqSRQYBCQNH
pmYkOfoiJyMoP3OEjvLJLx8fbVIsjyFfpH1rywV/VBnYU8ateGVLcSZaEsnMiJNN97GyNU+FlFru
D5lh+z3q8bnTbVNTQECG2vHOAL5CdW6sE6DfdxemQRQPUEfBzEYAZBC6S6xYcjKFX3PZgYOtyVw4
VZeD+TkZxF6uPw0oc32lY8sRbZLW8B1FU0Z4zZpfm+WpXD2escvLKdyDJB8V4ZFQRBw96NDOcyHV
tXNifqdVPFtfDfDcU1EqFd9teIoeQuwRnGdOFRGtL5RwyIEOXhTXBD/5y1KEiLTMTChLtsJaNwGk
blyZwAGhApKq4U7Hnikv5/rkNBoi1xjVVh6QM+t+JrnwUcuTrg3fyQolTKZ4m4i7NHzxWti2t17F
YuOEABwpDcCsHJe6hdCUNJE2/JkYD+PUXz4LrY+57rBvAMhBDrpfabcdOnHmuKl8cjLBa/3ntxyx
ioswS6c5XblsQwVEYDq9N4IDOQI32BMKJnqJEza1UGEELDcP2d5xGad8VM/jD4Li8fRHDItIy6sG
BizjI8QjNXn1lY0h1aoaaDolTUbhO0jsiJZfO7dSn85NLqyZMEftTfHzEQWRgM94RUt+GJPtxwyx
okQ3AAPzh2LOAmZA8Qd+e2C9dHmLLIOJQOl8viAym51dJ7Wqub8p5sx1HZbZ0VlxiGlVaFGf4PfM
Mp1cSRCuRfT/C7rmM/+XDbtw4pavm9yQbv0MeMOgIluLZGfseMYC+qtD8wkim6zYAYyW27dWnC/7
O33DqpXMzTK+aTFKPNE2IWCQuyTWCLsiu8g8hv8QlGPndKIAULhcu+zfZawIWrTpJx+ayr/OPv1x
v9BWrd1tMmmiJC+1BRYz0KELObm47gPR55Csr0J7dY1FdT+b/HoEhyZ7NBYM0YwQhAGLA+cbamPX
0tmfWgid7c4K9UZlpwKfFh4rvm5LmAMPat60+ZCupXk8uXPVQRCUrfauSmDMs61iQBu66TAMDoFj
D2KKvXsVr7RE8eX6BEjTwUu13tQqju1svT5QvIsAwXuUmNjsYDWAMx7aACsqFkLaY1v2NzLIgz+8
Ve/M1oEpDEAqFdIMqHOGzJTsgEN9lf3dUKBdiNu+0zFiEFH2bYM1SGhDPTvw3RmnJnPEbKYQVXgc
ZbwwstZ8bnDxpzFF3n/fnmZPZs6STJtclW+Bgy2gw6AEpMEUOQewahcsGd4SQraJKTPvOOc5yhhw
KJigdQWGRLQGD2VaAqcVBOCcgv0LfMBD2SAHp5dLrlKnsQF3hOqFBAW5w7iCg72/HiLyHjwxGm9K
9P/ev9PDkOfg5G3K+DKulaCYWov/rTlrt0jZLqFos1534G91R4lxbTk7b47jc7strlWXSDqfhiLx
J1n0rFiy7pVYEIV3QxMgT4uUIxYckfruS/80UT/D6ZwJwJZW94Fg/A7Nxxm3worwJCpNUMgrHApY
kCODICxo5Yl3lXcRFaaBPOUquMbIJKT4GjH/ODM/nKGgZ8lyjzJrOmhigHIpOmvJUSXLPx+zS1rJ
vxfEtHaM9LiJ0vbG8GQTzERYc1v5EOt850XiTjMIvzxtJlmb2d2nGl6DO9TI4dtVSGoPke/zhzXa
RjIhN9Sakx1vM9kdXg2NgICyZC0IRDIiKhMOX1XfaeX5hVH57jgvsVGlOkBK5oNidrozQ+IJzB+7
jxLSOvfZa2XG0m7v6Z/DtD4VeSUCW81ToYlpg8vOkh+HVwrah6paTlrDO6pX2KYUDddlJGyLg+71
Xy57+XsrOu9+4S2gz7/PDpg0D5I25A/59APeBWl27pvYroKYZF2u8uOsyQ+/Z9At7diIm1B2Ds2K
mSFTRsWvxkekRkW9sB/kp7z2j4mO5h72b/8mDK4m/F10VDZwTBCL5qIlCHwkEU+f++Fpg1+Jlo27
5SZkPJPwZlGECtc1Lt1TXz3PLSEgfiJvz7PY/OadDgVH+E0TZReVJMOpCkViZqQGVfE6N4buPdoy
MPmIsFseWgtDXg1COgQBgzkxrrs3UD9rl5ltfuYtTt+UhwdZ3n8Ge5VdUj0XmkVImB1cqyNRutXR
gcd84Vbvsv74GOnGBFyIaUZqQ7Vnt5eN0XeKb/mT3X0hirEZm8sp8OKNZxZ051qJ2bSRww+ID2PI
kFTTwieTK2e9aW+r5ilmPGv6An++CodL9+TiMsz/qRCfd7np6boXFVxRI/53nPhnlyv1nTi5Mm2M
1mgvLhFCFCbupFhJ3p7q4Rnb/3/eup1zpJH7RXJa0OCdCni9wQJG1QZskM7ZW/DLyMaZ08yjEq1R
MHozby1WvmCz1o2CCGEMejBP8M/yHThz6ZAkiCudWcNXolhbZDL/j+QPgUi3+cPy/Sx7z8hC3Api
XftXK/BAn3+WWPXvg7LuBbSnREyNt75k6Ekp40+BfdWMxfk1attsNmuko6YVG1j/qqySn88NsXdU
wSEsFuN2y0gaiZeOO5TD4mHp3eK6HpyurB6p5CHuAZPE4ZHaaWbSC6LBJEj6eEb1JU4JFIepS3br
7NH31L2xopW/ikdKLvThOF+ndO39D2pWhweNU/LzYNo9RPe3nr408PHFMlDOm3EJMqYOrveMJCIX
u8kCa26tqI3Nyz6Mq4gOpvbYjvnYugZ3N49iK672SgWp4CZSDivMbnO2BZzWqWzz7BHHmvPs2nb2
yFtVz3I7PTF2j/N++0KyJWo41rYpsG5W4R0zb1P1uz6hYwOCahW9ULJIoHCJyPzphCaRRyDLer3P
SOSzHwHgYFcPzvfQBDyXNpEPPZ7q7eVJS1vsYeBJJ2eNH5Mxcs2fqZY1fk/LkPNDVjzyGNegZ8kB
I/1Uqb/uBkGFop4V3FqaGfHt/upC40fLNRGlOUFHV3u6GLzruJ1JTJt63qaQ7DcIHuqy1ERIDTTi
BW68LSzxCy8cZ1Tkd8i3K7gQ63yuBYMqHqjuPbeHQdWwrcxK99XlKDo/9t+W+g/zUYAn25DT3iUW
GZe1HduAzQQRbNkgssPZnm/IgTCXjdvnQvEXs8vgbSE1wWfhFoteDAORfJmrm2mn5cU3GW+JZ+A+
vM56uV6opbL+jsA7aKaXCMgys82k+ejv2sfTGEEZJsEb7FzA47OQKNCwjRthuOguVXPhCYAqCylL
L/39nC1brnizozPVK88Ol486RMSKxWV54oO7Z6spt5AE4ObwCu/Ymbq0TZQyO7bk0vhgPFI34jx9
Mit7PSVzaFbMk/+wG8QPP27GgTFoPAQGiNYkRRu26gqaUilyay9Lmb0uvATZ35jQPORa9FXGTSy1
OXf6ZSV8BM7k2rTFOWvTsdZo/VjmUn88iHZAVpRU86BPapo0BK92oqD/Alektbs4oVkRL4APKV14
EvEwXIewE8k1lpS8yUjEbK6Sa4Stu1eLsijbbDGyRnyXOdJtSCwTvQ12J7+0ui7ZnWwtKR/EUXxU
s4up2yN4RZbrY6rtuuYobJaUdZW9hgZ83OY5SUZrbvWL+PX1Im3tE/7NuQHP9HbL+cJoIYoWMOB8
yI0ZfBPtjM0Qi2anPlJEsb1/Ai1BE0HdjduhCXgwGHUEZHdQqtHuPRvtZJ4NmaIVxnDY+V2M4HO5
9qWNZ0MxuKM5GpT+kqhFQeWSRmbiTmyGBhvBEENWc/uT+eIDY6EjkgVK0iZ5G5O026VLWD7SbCZP
OiXzRlcPSZmGXTlKcw6u3bylq9PjRV2r4lg8b4IXL89DPVgdDAUfzeE+drVcP1xLSBNyLnjMD8mc
/S3KelXoWGb5o4xFBYyPYxIe9mFdUR7IH/lkc2JwznFpg/E4iq6iztJDFWP2XmWcRHq644Joi2W1
baNkaN5SYJsupw29kQf0wRQqMvIsM1b+XYweJCV7KdBX/iA86p33l0m+MqzpdCfxWq1xV22Qa0Xj
zh0zXug3LyrCSGIexqawYt7UFo+yx5gmsXMxu7+5l/80bpTrYQZ1ckcJ0sf0ZROjRy/eWNDVM/pU
t5yUGi3MvTxHJPkEaXF5hBQF7rGJ77W6+lZL1yn3Kbf8oIKye65qAhdfifQuZMK+4iGmb1I+ZG9z
WHkP/kHNoxd8q4GSudsLnD/CchAAIGcDyQN6G+mUMDO2LoTy3E9w0vl0Aj+48Vn8htne9Z0rgP4Y
BzD4IFoExtlomgRD4M70jpcHcQ9eToqErVXX7GpBJwvfT1j6Y+wDfdizzVupLGx7KCBE4aOkkX/Z
sQko5WP3rZXLeRR4OQVeA1LYShjCdiVeWi4ugjEnvNc8Z63TqB6mYzGY6Y9zbXYbtFZJSyHgJu4Y
I2NWF4Prrc3BaQgXTdCfwdxDT4nCMyn9p8ik663glLSodv2KIj9lQdp3W8mlKwc2ZQwszmKprOoW
T9zcKcUOolVlSTf8l+iYFwzBhc6BVIijs5Bintb6gFbAB3HbBtooiNXYoQ+i+6n/RfccEj741MPq
y648YGQhvEmJmnsOft9CUBG5/HdJBFOBlSGEeH68B18vezW/kjdm8A+T2Ru3KAI4LyyO3HXUbI0y
hl7/tm1cARZnSRukLxTV9Nw6Jo7fpCaCfRxp875qcMJoTu468cfcpIJ/CUBnvqPSCRxhcpnNB7L8
Lmd9FKC9QNMDpQAvrI9PBgUf+TU01jFEbFM6PUwnuhHR7R6AuDKqb7sdxuNiKzrmpQxyGnpYOgER
WaHIdN2jpH7wK9awCJlPODNf+355yikYuNtIOl8R9PtX5GdlAcQgQnhz4AzDwZvUghMsl6a2cRLb
rr3lQV4XvvCA2SBKhHf4mj887TDWZHbydbb5zdZAPxmYQDWJIzum+1zCEgF+xafOGzqBXUXTaqqe
xnxLQsx5H+EBKOLrqkdrx71TU2eVp67hZfLAumm3jAggaR8MhDQRTLn/PLEqi6kMnUNmKlOcTeYd
swxccki1wXiZh+KHVM++NDT4GwyHb7uynBjIuOEC59OYXvQOZbQjOJe4/TFnEJPfUczNKkK7GnQh
pQwwlgKozL8zvE+YMIIVZmCln9W3wVW0AbcK/6yqw6IX7hhCeiDwiCS47KOjGv96Gz9HYrNl3ufs
5eqNyES5fjHKYu0hNzZkwkXcNgjhv8tFCIMEYQUVC2k5LjgQf0cJBIfxWx5OUlEsEiR+kZ6GFMtv
RG35gEqfnqwcxzPBgJ3HMpkxneIf19pn1EGrpBvci0T+oFVEwNhGGCyWBq0rhDWW8KlcBntM1YJT
qWn589AK+ABnZWiOaVjVLeZjb9wFHFJPb7QXu4BhlXt+qn/w7XURX1ACDeKP4tE1bagAAx1cnXyg
4wBl/RIvql88ILqG2i+KO4ep0U2i/RfA3U+mtxyn3Vsrk2uIkYLDyDTjJssSNTZ18STg3Ni+vhu8
7k12xzX4vsUpUKgwdQ9SaKl5zbNGAE+PfLEMWB4gPKDxXrtXx+rPlu1juPDAvVa45X6lOsFkahwa
u3GVosi3Z4O5ieiS7qx3lu4Sd8FOWshI03dmf63/1zSBE8KPrJ65c+DjJCCBIgB42SjYaiKnZsv9
53EW/5gijfTaHHKeKVIVuLR6ezklgbQeiP0tspV5nJQH3TLF5A5voYNrqoZI6bOIzpyy5sVpdiND
ny1sV1lGESQ7hWMsRipRm94j2sTRlvoWd7FHZOLEDb0rqZ0Egt1hBSNG2q3b0iw1oH1WCehlUxZK
QJzSXJCfj0gA995rocw+gapfkIm9QxhVbAabVW7NSkIvDMWsABeBqQmeRIErV3b4brxOBdTgZkVn
QpCBvGayz5hFWfY3nhEubq78bp9//rXSguhwHCyGvsNpksX55Mpf8kRKRh4d16Xmi/8r5vndExp8
xxBv4YOa1pGG82/lG0SaMXtkbF03JEDsT2lP8pyaaoVj8LoqAyXOYjeTtotlPcWAcX8zpucc/cPj
DTgOAmFU/JQBQA5rx4pZ5dXy0yihvacxxq2vI7D2QpAWVGgygDFvjMUsmL80y9qdtl1yJ4kd/DfE
DJ7TueGusCcTXqTYnY189o4/fl+pVs9r3wfbe5VEQQbvwgZG9xjld39yuNeWKJuGuLx9EtvA1gtf
wHCk2kmHY/bd5GZsjEZSv9qotja7TcevFrBpsLuZrVlkWQ4nePorrQbh1gGkTr9bqcCp38vLKcj6
JzPhMTqY369MKtYJfMScmjBArop0mw+lwQB2T9MhH9WL90SCbPrqf/70K7fxm7u/dZB7EMRC+sx6
qTv7hQPl0tIAN3OseFI6KByMH5JOR3aMr6NVOfdP9EiXkSRGNYNmif38oF/W4pGRPuCU9mq1910w
VNeYHvUCVWImB19sa3ElWbpUrntNGWV+CuUSssLl1Ifc7SsKxp9dOrejuwZHOB3p05xEu4fHqQBP
BG4d+bemQfkEdoxIKmm5VXQHuQZLCvbolbkpvSQwAG6M5DS27FG8e+36vEmQMwDIrjZiEsIaMJ+c
9+V64EX9KCYuw2jUI8nXHU0U4vDeWIMatTifR98CX/ixKptJHM6ZFySsyQgmlB+007RoKMmoc4n7
QnNUOHv+38aSPLzVrwJ/LZv2TnW+ePDjtalD1JlhvdM0CrqiMFVN0FFUQcVROWrgnzfDue37ZZSy
U/D51M5ZYpDrB5zBZFL9bBvJJ786abzw6vFaQGzz+1jHUq6UqnyYGK18HGEarUny/AENAi2FgiJI
tGFs32F8S49kQHdF2UxaJT+x+ZhA/uVGSRtqxcPA5OPVKx6589zR1Uer164nJQg08VGuUbLK/yv5
TF+W5f4+q3oflkpWDg5JJZwrVRwt6AoVs2i2wbwkZL6VaB/qH200eeTZfVmP8psEn9TNg5rlc7Wf
Gfh7vQ2wNLRJIZTIj/i8SIcU89sDE2ZMa8newXdGvPJyD38wBQTQGqMWWsHo/5UwijXNVh3ORKw2
YpdUS39FTyiVhVu8p1Jwyl+5dQLtiHiXN2mX2bewJJDhpcjTDy9a1xLk4QtvhzZs6XYak/Bluu4a
cZxWJ/YBq8df1SkkQMIcAbjB6HjexV9OsihB4xJ/XEL+qYL/RvMKToi/ObM6KSM+S5XQMbcP4iYd
+U9epTbVfcsDHxblAgfghgj5cLdylqgdbEKPrNGM2ItPQ00QIK9aVln8rOBkrVI7SW55ueQUep02
pJ4WyTFs5gcwlgpm+aMn40/kxs+DCpeLn0zFt1visUBH0tSYm/OtIYPCxZILAIUN5NTXWiSNdLwX
a8/tBQCuJ+DlwflsNoSMiA8rg+EetHs+jQopHtPhDrYu5ORfzWOM0alKasXv9TPficX63eIvnDZH
71Lg3gRLttm2GfSXWkJhpthQMzshPbZmAjuPoG+mTIjRZ3l7khQ9yEdcWK3PjkIyskhgUNb8Cvc5
wp6xvDcqCXItLR6yGisK6MoG6mfPLemzIWa2b0jZq/1eGffwT46TNPZKQ7bYTFyAoN4T6flCyPa2
uvI+fVcsW0wF4tCski++B57EyveLRiM3h1oAFiOp1uT0y9QkQdKnIKTGqJqRX3vF2ndCZSgRxZMQ
lzVnVydwh/CTfhHeMA3LTlUMjNWEDx0EVxW27rKtwlSrTJlEvZO3RoqYz8DymfYaIfsSIhoYIRQN
hDpmFl483ElolPdX9xy5oSiyHKJo1c6++UO/utb4m6UHY9V0vnPVJNM/RjBiilEB3GzcP0q+H45X
QDZYP+vDQEWZ2xvLeBJFG1xP9OCaFWfvN0efe2M/W5fh+HQzOIeG2TGXhAkWCSlkH+tXrQkh9ys2
QC7gUrwkE4YhJ0+joxTqPYfOpdUK+Lnbuxd6HNPfYKjfS5bI5n7rqkWV2ceEy+HPojt0fT4DNfFq
cCtiS0QGv/lExqabn38DibyPZnEZpy0/raXMbOT7njc6jqZ9v27fal02hAUz50jBTobUm0VaZCpX
EWDpzAjZXMxYbW/OlRCH3qQdZpm43uessfPXMK0dIr9+vWclB5tuqNo0lxt95DoK8TQXp/z+sF3m
n9z99J2toqswg7z+Y6gayv7RGQIFetZh8iO7o5tEbfBotvlmVEKS7UFZP9Sr5+TEUcg2LIoMCMdO
NE0dNryxZLK6Hu6EkGH+APTxb5BZRl3m7B55ISUS21zGGAoBxjqcj1t4opmUl3T0kXwFKFEYsM3W
9Nj/Yj95zL0AFXycaYWei6cTvZ7ws3UCBu2QrK4xEVrqkwp9dNuKmoXj+AbAwhxwG2HNIKa4ZsdP
QuGHPlGWtzzdwCy6To9+ox7OijIdKP0tLfuVZ5aWmqmTHC2VvsiK1wREojkJNjwBl+gJoRzl3zQj
ReWaJfv+547qQHPgLlvZMM4jcB35dv1ddteDJcru7KfxqT/PayTic9SMLfM1+j2cQKBl4NI/lXru
uU56hDEcw8CH7pCEV300Lwieg5Mk7o0Q+abvpvQRLVBYehpc7ElEBbzgTT2eRmaDrqp5qvqUoQF+
mnaq65EvNKYN1s23fK9KS5U7kS6BnGtPiTjwZEXF/nxyrQmfJapK3S078cPUlADLfr/pmfUn4nGv
UbYm7Z+Cm0UdIHAKotnQ9DE4iTTsCEhu50Lnx20QFRL2UIk7cpxtneqp2FAghO00B6YcHklKL0KZ
0Lvx+D3o/JYTBTK55FWjGukKCVMZmXDB81qdh2R89Z+1h6zlTjW7Ru8z9Qen7Ixc+7MMlXZIO1uw
UJw6GPhAkxHqpTQYbWDQw49mRK41eXySLnQ29yd6Xy1N/NiECJrE27seu4LnpvXkgv8Jdjk8FHHz
IVfEpV/t7zv57mdoAM3yNSKOoj+vfAcLZjXLvnR8olhSYCVadiq9FKXA3iZ0r2oPXOnITI+4/uxH
VNPOZDg4s3RUh6GVKoAwUHTo9wrgwqyMlYH/gYjLsFqlqaVf+IfyoByS1c4lk/uURi4dtKEyodMG
2yySxng8oI33NM/ptVj0s4pGwvtkDPua0+YgZLBHqeBsKt5XNJ1bC6CnKO0/C3pLRCbsTcP6/TDm
bgW00og07LV0k1KIpTm7i3MDFX8X5x2e2l+k2Dhodr4bgd6XMW5oyv876tl1AM/dmPhPqJMhN9OF
5VoVVXenznlFRtINKhHPWUhhxLSrL0SsrnnNrx6bcevM0bhtSIXQx1s19woKYyuUzl2JhLtgkfYd
BOHtPSYrm4edNKWMbsCHIzskn6NojaW8Kr16zCJTGu93t7CW1j1nhxYg7u993aCiVY2zan2wB+Qu
/p+dm+O0/u1wg9v/ZX1HPJfIGY+NhnNuqdPAJxOx3VRpm5c6xkXy4IHhLGak7aklHXTroGjTOZew
gB25Uz0qMkyt20eBbCeH0MXYp8dN0cU5B8JlzHApZT14bM+4GWPs2dHq7otU1UEDgvR8dBjnc4EG
fByCgiAy8NyYiWY/WZuOxCtUb07JaVq2vdqMe1HHMBQK6ZltylD10m1+rOcO8IOmhtmhXav1NDxY
kENJpUUJjwigeemy3WEwhqqLbkUJ/SgRwZRmSZLYkZwkrD4jMuf6cPxQ6HZsGmm0CjGgsyn2T/07
ZhF49lRcMt8BRBh3mCvfZ3mwd4Fk6PiGGJR7M6hBL7WKp7qViZhJlIqKJW6dqhVsTulJAHHLEBe9
3yHw2mAx5/hRZDAVb721UsV18cxePi5Eh1zP9t9NQH5IOy1vdcBLUmUFABoUv/xiybXDraN5Unsy
69s/JQruoXLD/0hy8ktcOdNbtHNQNAMIGZ6HcAlFBuDy80sUIu819KnicHpE8RQZBF0pQEO0tkSk
feHtnlGsMcd2MxhrxdoDSqKBXOUytNZyTyOaEXJiCm+V/G9z2a3/DRHB/iy9H2cUd7o5b44Jt1iZ
gvlJw29kIvLuWMhIQt7IHj4iQfCCmUBj6vd3IWWuPWOk0vhptUZ1pva1GRelMFWhalXEltFRKXHB
Czb0y23PK256uBJ8aY+ePT47YrKDmNp9j7C09zs3n23OfNyCkpDzVl8z+5GOy4Sg7Mikzfzd+toU
st/1P1xtJD/h0pJb0VWj7uhYLRFonn9AaPikKkUX0s9dA9A9/Jwi7CE/TqWc+EI9xlItk/ektkIu
OtF0MdaQUkCJmmMmnu9qfuLSoVmJtXVksCtmtWG6monjwJib5b4x6WS+4MdLKoltYz6nu/nnqXbk
FlZtSUyQCFluvonLeYUVkjnVCEL2I8Q5S7SqpbP0d/Ue7ggrX04aKmizXANQ8s52bQF9SUiEZjMw
9WCwK++ctv32Nz26Y1Lqj4TBgzFZo0LQdFoGamymrTMo4Jhc6ET4zoZaLSOfZPWgWUMMaKJ/tWnG
sKAe86okCvfF2zX2Ow4NJ0FhcQV9eesaPzC23o+C4NSHzPlfX8WQDMH1AZWq9jKOwhd3wLkBPey8
PQ7wJ+Lg3NYr9EP8Qw7S0Ix385g2TTb3jFLvVorW3bSttcw0afux0sotC7AyilF8oZneGnfqo+Lf
DYnmD6Bezx4MIg24GgjDPPMCHNh1r//363+mwz13b1r/dduwU1mcEGp2oSG+eu6TOuWzNXPCUIcB
uXEy7WIdiq9F2yWP2l0vzySj65Vnrsixx8iq4nDoLn+Xsubw4ZgwtI7rER6d7hLtvcWf52B+aSKw
CP+hRWCLw5pnMDSAMXZ1jlwDPvRFS+18ZsqOkMf7K2QC6F6EUlHyGXOaSOpot+2sn6nESjfy4yXx
CP8C12AF7rSXzWwr428esk0pG93YbGb5eUwKHdL1nYweAZ8YmkrgSrIucWQrZ+zA9npcts4AsMdC
czNw51/0KR+C1OX/FWY5Ub3e39hzrjrmXCe60+OJ2juRp+Ltl6+1WR3DOokKqvj/k19atywATgQn
jXe3wtvjYhbaHt/GhzNs8BzA7XxypisytbxkY20tu2v1f6Gx2O+4X4kUcHrH7Ov6yL8QoIUbd2MI
nBCb8zZsGEo2accFgCs/meyPuF6A66IRfInYseAhZ0RsxsL2zY/+HklKWIzsVoDfK0rUUtY1uTUK
i8PQ0DH/GfJilcKAVmgip6AjOKhQhaR6CUvS6SI4i4b1QiMEN8onipVY4A2I8JvgRVnPNz5MrOJp
YwD/HQd+OmHyPy58sjduRbvxfaivCQQ10Uj0gztJQ6Er4r39MdJScjYreh25S+dkRAGDushzjfg9
sOdvoS8sgBUtGKYcFICAT44NFJQKomRUexXgkfTJqDx2nhRb3piA5gHOs0pMj+Bjre5rh4Zi+Ukx
budWkwyS1gIB17WpXt+S23Ykk9Am3hsi+GXzmUK27pcQDLF00m7mLQv0LBaftMtHGPEApir20/Hn
vODm6tunQ4hCii9S83hwKh6OsUpfSdqwGWbwqDUBY6pRCn+UxC+4FGXyRAiwR+F2iVUhIBj/d1tT
u2IoPNDeVeqY0mJplVdzPQ1OlY0KB8Bw9jjcblyq+Vf1rllc0P317SCGAs0qH4wfO6ewtBC555+6
Zru9cGle0/TbuyaHRtO8WbqFDg9kHW+4SVQ5nQcHpp+uWQCouip+X6vIOk6TNnPxQTgWyxuLrnUG
8S8jls4um4xf2GhM+m3isbGscli0Uw9S14bQ9syYFvyvA32oDloI7Ru0zsIY/qki3gmfZn2dm6tW
+enFyU5QyDCx0lRSxhI3T548iic0/Dh5PT32aZFPurtNbzJ6ENGwtny8g7IBMr04lYmHBwMdsQ9S
4273+EC00dxSaOSxdEgak92ITWZEcjQCYnNur6U+ZbBDsWzB3HpC/wqZP1mWs+t7POMjmyabJUYE
nxWr1hY1TFdWjrYkaLYgeAVWGDPzNyrlrMftKtaVNrpGpWbMLn8EDdfmbSR4mvm/kLRiQTFceySJ
3DqX8BEv8TtQUkiiNgj8OTeYzb3IrgIiKWSosqtMfif6/UCGvSgOwcmhZj7ZlPHLTu8Zhq0Z8OrP
V6PGmBMN06pZLKLbzfZDDYp1CK9+7RpOHmh/4h9BvVupWbHW2XLkLoWOa5Gy21Vjt21OkwP6UAOT
0VapVXpmkHKyzedn5adiNhmHxkZE1PwrqNS94nOzY7DqBKl3/7XpnxuX5+goccigmCaBFDELdhtk
w2PMIan3SKTsQl0G0j12mzEI/jJRPSV8H19Ku/ceUGv0Z5YbZazbbCC7klGy7577W8gg7Bx+mgrG
tuYKAQ+HbOlA9+mu/+hSNyvXTRNZenU0JlPWb69ZWdgeOnvor2rYpmoevSFYj0ET2U7TSAjP66ng
R3BYaeqFrAZdjMa+NMkDK9d44FxlQi3a5IMd0x7PK7EEYd5eYS2Qv1N0b7RWGhgsueB047B9fIM5
igYoDGmxdmUDshvtHrdcefZbsd9mfZCLp52KLv0PQq7LQcAtQWxAn/lBg0ieUuVx/VWTukfb7tGR
Zfg0luHtiPRc+6X44KNlUahXvbNg2phW038nyYMHNmZ78PiGL1wfnVvzQFIftthFwyotMvHGxZvS
RODiNCQphIRYreMeF0WchvQh0Ok8ZQQURShFwUUCih30vb4OcO+B/RMR95bzlIOaF6GJoW7f+m53
yVft1pwWwzfAQnhUGKosIrk6Yq2mEU6cMyetTxY0d1R/4/mfGpU8UWE5p3AH3pVG/Rw5q7V5vl/y
peWg13Mee/Cv7aToAof5JLd73oAdCKH4RNKTkbnYYGEwWrrfuOebl3DmkzMOo8/eNgMp58eFtNMc
poiczGOeJT63VmxtfsVV3ozKceP5ysooV57Rv9+qKoRD7YPxyFhaxhouJlGLJaNVapEE8dycwtaR
dB0kmGAVZ7zSpeVz7reuwyNzZ8+08RDRFHyJMNP3KFj+H+qe+I06dDaU4YE/VfKbXZ/NhUKYrYc4
HaiTHzo7xF+qlCs+TbiKVTFYmZhnmBwXInGeYsUWM5jNVPL18l7QFb7ydj6GRTpdgY8iffQw9Sjf
UDGGqhcXxt3ozTm1lX8epqR7dyxgWsEAMWd6N1lNpKgGWfSg13jQMHh1UJ/fRcL2hYPlgP2m4uOp
S/Yj9VNVrGTST64Di+PRRRiUsyvcUsQEnu5/gsiTJB7hNd9bKiOJR/Im9/an7YMM92syuKO7dPFl
jyuyyKxcPkrdTQ2MSc5hqXHtuCzNu5rgD9GnEE5Vxd4HY2Js28D5W5IRXZTXRfpTur9Nrl+qyxhS
PX/fl3ddMiU41zFBVS5eRSQ2lGTWzysAqDlRyRBLOfrkdGFZfATYEQAeG3q3cwdXNvIkOAohor4w
nN+FEwpj+XY7fnnCMPNRpjo6s5UlTnFbv+yNI3XukbeSRCuE/1sPFVyxY45Qq5gV+6oIat+aeAE4
NkOkDH+sLlRJWv8aFR2/NtFJWVw8FCoWfutoHen2c4WViwGrVA8blkgPYJNLF9ITQWs8dOKJ9SbS
TdFeUY77+G0QNV8hFot4JGF4XDp034FVtCbXU9O+PZnqaDXS62g2hpuP0QZftL1vpGJihzsC7+tf
1kkJE/jomWIKAlj6uGWy/YAwGrUJe4CNlJSYmxzwYdAmzN4JS5T7zayZTg79Bo82EsVsVWDBAtGb
kbTd9C0do+LkUwVLcOQvW+9Jbdc5VOYP3j6zOLyo2V0kFLc476JjctM5YSlrRvHPHaCvQ3DiWp/f
U3wAuJadrZa5fZ0FXKcSFWMdj0MHniw2FnwMQmRQjTc5dsPasNcGJw3VENVMs8S/NxVnrMJgfW99
DvcRM+0spxRUPTR8YnwgFylMooMbPyt087xXIiPDEeGBrvX0UbJngILxeJVBmiV01Vw5s9wSi9Hr
j/M4lzvBJvtZyZSHDWWn48uuYqj7M3vajdjbw6ewLu8pvjh87rrNCKpITspUDEZZ/RFEnzk0YJwa
88zPaB9IgP/I5uUCumjXW+tOT6pWc19W/zJDwbhK+GHC+XcehMQb1DBh9ZnDW0ZC6VA0o3J885di
FXJutDscjv4iSOOHbugLKdAS9EtOXGdaZVjTaIrPPj9HXxUFPG0ASelWZDkKKhVqZSX5OKhSc/ke
NTmH3ZUz8tGDmDxx7kVCaD1lHEjjrXuIuHgm4NKtnrXFhDhZTNr5YyqpzwB/Wy28S/J45tDNup2m
WKQJldbspkRadT0xZpzJ5nYYOrUks4fKserwgKvGsvSQ2puCptXuz5+tMfSasRE5BbVHr51XWbAF
jJyFVrbyTw9IzNObFBqsyHBO/4fvZkLr+GUByp4UZRUD7NgeGB9/eZ59qbX362m523ySoUrvNtBh
2bCJOfcNpSqqkGu8kRFtSs/8NCWNypdhX8nEVvl0Fj6vLxc/5k9BfkN69Dot3cHsYFEVu4hJoyB3
UjC4xJzqvbTP63nEEvY9vkIYEvrIPxIshl8E0HaIXCCoaD0uBTkn3D69ZsLd+sBW0vTyfcAkHHZ2
SPVCLyPeQz2IHYOLQp+tD2whYqQrWhQxp0S5t61gnheFqJKB3iqMjFrMMI/0PrkssQguGUvCXjM0
scOkF5TmCoxSDcwGy6ZfQDr8/LqywKX6u2aqAsWpNmjKermKhiwJA6TS2XcO3NP5TZdSrlX1N2/G
11DtKEU2HF/5OcTVJr+69gCgRkw2OuIoNOzST4iV3gPW6NFRz4BGKcatk3fAbSOpamuNe4y4xwA8
N89t1iGKGzHiwDeByJk96BRkD/bkmXIZJNkzgMRnGJ+7F7Dd+PwzrFaesP6rl2OehKiOVvNZBZuU
71cZM5sTSxE3QJHLBLRUUjQ47E1q1WCQ44wE+Y+EWCasfFWsUDoINnSYN/1xvv10grQMqUsUUr+l
9IjLbqKfd8qbO+Kx+emr9OEZkMqPHy6Ak97uGeSGtUNSd0keqlIiPg9ZmGcxLDZUGr+/P086t7+S
x42IwsdYXP5rYMWBFfQCY4sXMVCbIdWb3ivxZdq87o+WLlyBNK/ZBeHEVGnYiE4Gu9xmn315BrF+
PZcez0/MoetbnHQDxaWYAACfhBOAx9NGuv1jaz9QfObx5hJg2BAUhF5NEagy/W+1g3hjYPJuIuBF
Nr+MK4KWgcie41UFMNdYhbBU/xBy9+dDtNwdGuH4f5czp5czbsKJ+Q7pQQyRfmKewl/EyVX+VK0T
JBVdLdzLVY0/3bubAG0c59saWwrMyC4YvPo6W9aiMyODIzeyk0FN8L3Yji3Bg2HcCyoQHSGK15Ir
jOpDv4TE5ermll81agueXrm09ln4JkOuUQiav15Cb2/kahtXp2GDA7f1ho6ASaOFi3rP0vhDorPl
NMsg1CMl8oJVKfliT8Mf7dCLoJLKSDtBUwJkVuJ9atzyMLVqyDDGLsptZRZhR5WFXOQXCyB6EpBX
ta1Y9jNUbBxe7OSQFslTveChBp9qZxO2+6//pA8axqtDWCcYXlJxBAVrrrvVtUwnunTkEVWrxu9m
Lk0tiT/5Bv3xAd+g02U8njq9BLlN1DvW5dMD1Ya/PmkKVVMUxy3K+cirpmHVUQ2+BOMbLqF4JIwH
Z4w2GD2YWfDe04mqHLugszoG65O+fLRQ04amRVuis6DAOeu8SY9uiytbcLXVx5rnpEQk5aYFvdH2
gy6msoxBfoDWOCRWDIN6rZIrSSjvZJMMzKeDrAsEGyo1Rbq+EA9qDIMHm5ubKCl+JbHI9yDLSyn5
jMe9ptMzs60sZvaiWXJS4KUjQD3J5i+pht3Sh+t/ETXcHN8pO8r/TE3vRPmG+R8IlBeELGpYkIyq
/74mZ4yeotvQybLhoOkqvLk8PEHAhak9rRiCWbdOmwbCyr65rnKr/A8HvKyxN5d3wUi3RjmmEPS5
Zf19qV/5+0wMvhutl4n3oyVmY7vmH/yuBvC8/XlT7Qv9HtKZk3KcYg6Sny86d1mxWDNf6dhKCzmr
nqRLT+W2HDF3C2sEH1U4KKAB6fWRPlxYrd+V+kl7AwJfOM7o25bjHVvBFq1eGdCihH5/zlPiLloU
Vp4yD7nbNBPwKZVTnrFRv3sevrXYcm/ZvUgSRYOe9WJ/u5lVMus3ivBxrB0QbKqW2+vp443cfyN+
lgY+W2GiUE/wmzA3/BXZH1kQxGZzIWNL5zXNbkhKE9Euve4kTVfSjfOGIUQuSR+pcCmcMhhhVaLB
figc3TL4jJYxYWHEVc808QdGRpwPgyXTqzkmflnTENqTfrGcNbgBib/l6LHtXePrnRv3XX5pScL+
JvxSO+AnLPFTyESAuVoZTSe/DKJEoeQ3zi7h+QxmWkeeQG62qs+qRLKy+lRQw7RETohkwblB3GRZ
Hl937oN5ucQyYGvbJ3bwhmTgpZ5fKlfVjD1EXPbkiDxaSf3XjhkOI4Bnt47ziW2dLSmaQBLnCTuS
mcUD7JOqcWFqNl9kr/c9/960fJY8eDjYAuETm8aslBq+6S8vSWacxrYEe2/STOff5rRI1KqF62Mg
e1epyQ/TZoSrzbTl+1NUhj2o8cKjhQN4G57b97aMD98Za07AF7CBFX+Aw/3tlxUuu8T/9/oRy6zM
TZlffukHfceGGeFJJuC3T+cBfDIewbM1g0LPAQBA73CSfOdoJsK839kUQSnsEfIF2jPQh486/FDu
5IotiK0yS+aSCT1lJHNUYGPTLEb8uR2okALoa9MNccs9RAI2hCVG4V354r9isNg31VuXBuUabbp8
6GWuQziTwpl83nkuClGdklhKZbD99va/5QZVPt+dWC6HThxAmbE6lhr3f2TfJX4WbG+ktX0XlXjx
Eoc/Tr220iSdpj36GBu3IPe3pGfGlJ7/i2R2vWrdWXAFHSUXysFWcgYLN4MoVbeUZislysDFw2MF
pEB1WXCxiXWh3/fkdw9z8jnMRuZNE5imujCE95t3AEZsavrX5Pi3oGCVcqskmg5EVwFIL/dV+5Kj
gwld2eoYWOs6IIKoZHPIwxwBszE+LCFniDGrcrTajHbjt4GNsSwVlhhquAvv/2SC0uOxLrFDE/I8
r4jrh5Zi+fJn9MAB3XXQ8cLVRxOrQxIJa8BrxX2+lPZtWHEmALmP2h/HRwz1mrR8Y/gNlWAb3dV9
KVc45XjCpdk8Dlp7ufPiT9bXSG1vDL6okQdUZOxsoGshOiDiUqm1AtdEKcfcN188IvoGhNiaGyEp
v5/EoX7Q/TNO+Cuv4QZWTd2Y+orvBwq6kxsxRJKuPms4+JVO6rz4nGedAbWW7IkqdmlLLqfy9B4q
Q2qLDqErlxYLW90vhNSOp5isHdL2gcKvLdLBfVEKd51cab/mBWmhz0dKt/ZEfbuJbCdho4n/zv4v
Il6XolQtVnzMnHG1ZJvrKdOOG1s4/FeAy8gkex7An27E9NSVcA3/CAJ5vSGXmAGsX68msMmeZiZW
JQB4+HzoFbm4XfziMJsqtIZT/ASFcFfnOZZOZacy+cPnuTgaRdsEBVR3+QNDN9BWQEYCb48cmzOf
BeD0OFt3L5uTJ/WxZo3YsQgVavoVDfQY6J1YT2o4BGassT4btKyiSoCj8IlyPCHAxIlMgEQpPWFA
FkKjooTMepZyOFTAlCxV7b0UY4ZerRuy/rWxsFrc9Zn22fk20yZL1W+oh1zjGQLtbrjQnyKohdEV
kkkFUGURJdYzJB7GxLJJkWvjqoID8PZlRLMLQLYTeEWI0zUOcYgv5Aw7EiYaop8E6iRjfXoCVZFi
QOZEnNFcn8pl1kA0Geizht7/uAexzSPrFODBxMDLnYQC1YPS9ZBxxU92vl8cA7dFt3cU8Cgap503
RmXz2U9plNjHzloRiO1R3NaHrdS3IAQamw7WsWyjjtm4oxc1InMNtyuEl4V0nyHT08Ba2xNRPMPl
MeK5ooiSU19Cv4SlLirArlqGKyTI/vgIq3JYRoAQFg4HFuXDnCFHMa8K7iShUuQLxKmzBT3fNuts
O4qiJFbuKuNMKGV8uZPG4BWIrEjJfE2i5KOUx8YVxF9HI+neL3Ep3zrSmOitkunBKpkbZN7Mf45D
YPie7OvcXmrZ/3jBrwMvDMFpdKwuh54euNNhq72c5A5h6uvXdXRYr6gPgBNk56GDJtZmJU16vP8N
jQb7M6L64lN0PfonnSM3OH5M/TW+os2HQa9ThP2kkKG7v9/Wip9qd29woMxv3ehxKEyNMuyY8s6V
mUMZ9lKTBNQr2G91HzHhAt3x3vV0Br2Ng/NWj/EiLKf6/zyHevnpcqrD+qXsEREonOvHiMKUCPoi
MePtUmSgzt6zrdMKQ9DkMSMKK4Q0Cx+Za2Ouno3MfeDCGqxXmpbIAlzFOtrQ0Qdh3kJ7nxqhRuRC
s3YWAg+6uO5fgfQaMHoPuwhrYjSB/2CVofwOKqYIuNhC7QITMD+xWBYoXZPU44KppEbnwFpQGs5j
rsOg6XcnqWGO+43iwdq2MRWHMS3ZuisErESOp5kdEfZAZBUKlfSWkXFBf93rq+2wDEQA9xcVLMDf
kJh25pjXCy4sNhI0MdbzAGwldrqYO2h8urSBHqYyE9yvMh5BwZYt0rcUn3I8D4tgerzwrbzMDRJu
3MnCzP/Yoksjv+TXAh5TuiOns3rTlZL4nlUenydCHc63cMX8nKlcTzdnLCQfUMlWRpofE2Fi4hGg
oLkWMcqeXb0hQLBwRmTzYs3icaUwSzxDyexRL4sBRt4Or9q+p6xbXnXMhk5x7NPFyiVMdr1e7CH/
JqXWbK+GvgaeNL67w5B+D+RJmY4GbPt2pJg0KjuVxc/eOAcw57NdgRJ1yjpvADIEt4Qx4s9H261t
kK3gpi9+MLD6F6bMUm+/CFzNYDCoj7oJpug2JwX9SLyuROnR/rYEWVauUODmv4R3uF/r99/rzs2D
iUe6tP8EZV3bK1iNbTzrNbzl1Vp45AFVhroFJ9WmkOE++Ujw5WM/XoA35Jw0/U7yhguJBJWZnhgM
ZmCVg+utw9palWXq7TKZiiGkxADZyZlu4ZbLIU/WuQANg+txYPgp1ra3u2rUKngr6WjG50H7iVwT
j2JmWE4dO5+E9lulRE2tzK+zy1Ox6bzJOkaOhw/eoP+0r+XbxC6LX0T/gKg3hThcfi6JTSHipcnl
RymxnZJlxuO+VcTohUmPwav31jzf1jL1FLj09jS475LOz7XF6i3kaLz8IU82T/aup1DdM8cbBu4z
X8866p/HuyyVqBc6p05MkDiBbj0zLYXFTg+sW79Is1voQ01S9dhTMm0NmIePjLqbHTizuVUUpiOV
VQUCLsbvvSeDTgQmj83Heo9jIKafmC1boNsTyz6zJnNv1dwJnCXK36qgBq2y/yRMK/HbdT9JtolW
jITRKPGX+JZokDmbNhwzYE8o48ALqazdnWzGLY+3RIcYgVwvj1L9QZdSZ4vVeuVD3xulPeceZlyM
BO7sNnPLq+ioHCYZVFXUvYipOk17AjaxiCn6Hx0XXaI+uxchwQgiaU2nN2XjTWIUsaTUd/QlWamM
kUzn2hG1XXvK81wmo2AhEpOBJN8OsR2lg7WYTs/R2BhWaISxaNC7itCiaFwlWr8GyfFZHqnMwW0n
Wrzdx2SwzB+95Op5oDL7kBqJ/FzGXKyD6vRZMTXTDvd2mODO9laXgMsk3bSsfZ4ees2rG2V/17Bw
HRMtIk40475cbcpPnx1JPJGo/SHZ38tPm/6sVqf1hcCPzwrYr488W9BpQ5apGDxAr3PdD+fRmase
iqi2FPm0hL5IyRT1N+fsA6bgX1YC8CIHFHdj0T7Sn6aCHAJBfLQG/UmxjkPLOvHus+mYGy+3xjzz
lXzR4YRnksTtL+HsI3bxgQzHetlcikYxKTPe8mMD1+g1vzcoNdE8d4MLfJbsb7L3DmQp4cAHtlMW
M/gNKIJ6xly6/5YHJ0f9B9/LRZpBNFgf0487JiT/nBLcpGRDElo1pt/MT5rfSG5J5CLBukrV59/W
ptt8k2VQ46CFYxyRNf0Xs2mdb4j9+tBdZkAUMAmVXIID6MKnuzylcCWlHvCl67pxsre1PpzdeFt8
3yrwvNRKzXl3x+0KWsOAomuQHfzcIEErpnXlZ42ZoX7UhTe3/L5WiELztgqKDJ1+GvaZTIZApZmQ
1yateRvDjNnfqoq21WwBNF34QuFJT2iwB54abjITJ7nHrirPE2732kObnc2NRoIfTkI0wn5H6ewF
WutkjZG1n2SqgU/n4DwCQXvQ+O02lHNDra4okUYNk5k684fPbigffBNzrWlecdPlLtCtA7WYddrG
RKoNVlrSNlLjbxBXgEyB1BJdhYJr4kbyGUyFtdeUhrn/Im43ibRJcRnUBVQuIuZdaZvja4Cw5aMy
tzWiZ+/r5LYIYOFA7VK0A7r13+FSXo5fBqI5JbCV1HbHN2Tdl/MrB4XGm1dJgNO+KKRpy/qMrHxW
qAjqlKdL08gtZlX1nk9sZcuz8nbq8ndKVsuJgglHnW/PGs1DZIB7IPEOAJt9vw+Tf4yuaBqkRlIt
Ejbhg11GDaUbxUPb6On4uPGnnOTeB4GRmZxEZCmGv8R+ODdhPuwt++VY3mAOTDhqoFf44a/zuPzD
FVrB6Sved+SD/IjmS+zWQYIqEZ9fGkFJho/z/qLsS2tUzB3P/QSOX0dLoETWxU9Wc8QUf/u3sD+W
SpAdXWwUoLCgj4WV/A0a6bFaDTOHWiXK61oChFv6zJGbs+J2KSI4572koFTf9NwsY7EucWE3+fnj
76Ehu32wC5ur62nlcEljOmOusimHVqEhdczb0EurCqhEJuMQfO7oNcrDd95D0rSaiH0M+ogNyskw
Q0Xr/0N1KK7lfif/diWb7ADNWnq2WJVUdS3NGe13yAxtPBRVvhPvD6d0sP2GYEjaveHctcA2W570
7xzLyJv+SQH1OdtXwP10GawN0cdtrxQH4Q/edZlCFVM5kBoUsqvd7uA60RLlKG6k3/SluUOZSL+D
XzA6dQDIsnAzwv03GeYSTxLss3tdIDJDJRx4nl28iujLY/3XYihHVct7+9r67RS/98Doe0sevwKN
ogkwPKO08qyKVk6jtn9PaNpi8nRt+250wE1P6ITZaQxV6hy2AOBZsuF0V2z1eocfNjVcgJJzFGY1
5RlWXoSQwUODkDFz3OLuSWZKf6Qv4+L9VLjrxdNuIMd4kkg0yKI1581TWAl4XmNcZii2FqEf6Uar
ODAh9175oVZDQ3XWGleC1I4ibI8ZsmpQ9D6D4vP+iD2fF9GNGHG9oNXUaioawievP00wdS04SNdk
fBbbv0DyfGDjv0kQyrbtyE+YaWTBU/UmIiHgTIjdEFHzcA8QJFVPcxFh9uRkyORJMW1s1rPW8ntf
EWghvqffcX2yYyq0iGoY0A9QduRQTelVvbe8bEBnU3Mia+Gu5prtqHjMU7aoQwKmbCc8YMPJnUXn
B+40Qfh6K8Ps0coIUd1c2qtTYhL3kKaXsZswHZUQ9h2BXOI3PNapQtVWCwzJjd+m4nVN7T6NypJ4
G33ZA0wkysUqNzkcXd1KngKmFDJ6tYpxYzYCQxUGss1xGMAebIkfKO4Qg4NRltmqMDLjFIQjPv68
i3YScdBcDQud9nvibZOtf6aCFqkPikYfo+Sln4YxALSY4UFctGbJrQXIbCUB7DeMWZAa0fvi9hIO
Kf0NdICEoGU8bHkBANn9xiBERCx7Y0XrfYwnGrJWPHVF+ENAcjf2VGS2VwH3M0MVDxRtZuQpoAEt
4WNE8Bws9U+vNeVANfaidcNb0BzBAj3xOX4/wS99J452A5B3pGp83E17nqJvvqRvrUPVdy+ziiKh
uggk2mjNCtQj22jhvW7Y8kVsL72e97yXRb+K50lFdrsIr5gMP58IHTn5QBBahEeLkFbYBp23i2Vv
BUNZ3h6Y5KO8lkEIz4SGG9s55Y3VPG1vO2DmvmcmLXa9Px+HPw6ZGS2fi698DAX9MF+yldP2l1my
wlNibO2Ogz4VJmd2FEtohh5eHB1A9UE48CS8cC8+D3xKoGVyiovpUvRm8eWtG8P3zqVkG74QdbEB
nvM0A2Cxj6JRYENb1+96GGJJC5bGPQLwcu3FovI3rCl8pWG043OeNrrro89+ckv3h7TiYGtz2nci
6O5m77px6UYhS9pBZ/0WwMjZvn2TqwtjqLre1BGcAe1Slas7djpBy05vQXcaDFUIhnZ1NyVCQOWG
d93DWiBXNQ5ElLqQQD5O16VjLB/6KhJkpRSuRytg3esUmaQah93sZ3TAOjAZXQAXcNE5OGWxM6XL
Zt9ljwsbsRuASvgtKshZfWmUWt4Zo1VxzsZa/dT+hE03LUtTGu6DXlcEAh2uQVLYqWtuoupyBEVs
uVX4XKjzQzLw+BvA5dIFLvZhFclYj7Yu7LudpDrbwJkqrLgjGEuJSxu53O97Uh6kXLoq7T4T0ev8
2P8HPKPDlLqJwfANnzBYQyUGmSmqovf6LQ9nx5sS28ZcwVArL3wpR55WWEPeaQhA8pngyjghntCJ
fJPrvMSYFo7Qa1fN+EGxpDZ+U1iqmw5ZdG/Gp3ssfVlJT9rwUTDRGr8mClcMhyJIlHVGcnzsU/qB
GsX9Za7f7UV5T157s9aditsn7illn5SGHgYLXD0IUdVKbs1b4KkTI6++UsEoO68+WQkEUYRRk5HQ
N+ZDrJhTL+0zZOllZ7sITaImS5u/TqSA1RFG6NW3v2ZjvA7ief9yvIXfg0AZjgNZ4hLdGxomS6QP
GvH3yi9syXF3IrDCpJMdkgQWmR0h0/P+W8hTmRvcG3ZX70sE4mYG0lZXe5zuHWH+tIlcUroyInR+
g+LxAd+myBSz55oxU12j1c8lDcTEG+kwssrudQk/cret8+M5TBNr4zibEBUO0mmO3Ef8I88klH3Y
oazeKQq47TS5o2Sds7ehR0OodTSKZrX9eNet5aPOr+wGJvs0xwwh2mpkq6H8+xqzSTBomgitSr7i
TNGeq1VtCEmnaUUriJ7V1kPpF0jq7Z/sbkjgSLFA9LPrCkR8LLQos2WpJv5+o3FAciacwAKVwXw8
pVQTHg9aM4Tb05QlJwJfzRds/f/lEjzr10EIkkVioAXAfl4BSX19y7WG03aSX71sgRc/r8j1ETsx
4+mK2icnvejxYsLwEc4INKwPHpamS0z3eMMmmgipx0HRhelBmDXHp5wLeVzA1c/WHKgvWyohlkcc
0jDfvOiVzv86bvWUEbpkCi1/mK70whZYrHmBwCCbeGVv+GvwN9V6BHzSGDwWWywq6hK5ajVkg5rj
xh7NfNgbuY7/3Fru98lmg0GsOr9SZAF31tIKTIkJPwT9yQCqZCA73wS9/Usg5AUrgway30IP9RTx
+AdJ9T0nbX51GnRijaBBiCeNuj5TAnMQEeZn3OCtaW9jOPOK2g4zQo4yQdESUTjJQLQlzjDGEiy/
2JaNo/CPS+yLL/yALL0HBCa/uBI6ZbYg3NxUTpIbIIUnzjLi/TX3K9pKapUnybpif+8RRiL1rZ6Q
HuXNbUNbA6CChiUNk9QQS7rgalntiWzjIYUBzi3Kor8mOeJZhBoqHmoBy+o74OXSYyKvlC7PpkLD
f9SSxLn4qkCZ7p7Zb9GEtTGh41rm/oU0tC6bq2BMFU/9Np7fw2O5ehW7gvUPZYiabcFmG/DZT57I
xzrd1aFhyJIkYqwgJ60Vy5ug94tElv3CyuL3nltXNKdrR6jdRdUXpxuBHltZtXS3CI3cZApqF7XD
IO/RoCViePJu3W4kd0q8DuBqCx0V8kcAUAVRGCgPcDJBoABnq5aHoln8WFaCmj5VE9vfnd/euGLK
Q/rVFSedC4DMDIr37rdY9+qn72lpbcArL6MnvHLS0btt9EFGMkup8V6ly84GLi+7Q1nRwUK3u7b3
KQW3xOEJJrqhYvfuCqJktkolxcwq6CU8r6LaEev0imt7QTBblU3SreQCIq05dmFGrDJqzCfT6i2h
z0hFeFPqvtZ7JUw/AB0JjzxjTWu3gmVZA/cvCimOLANkAyFto23fKLlCUzcKPU1lA75E6vn7zByd
NpLI8nODqMUf+4bIadiYixcn0pZw76nk9IyCM4lRT7v6aoMbx++nxsQW/wtuLewA41kINNbVxLxC
wmfoZ8/9gUNZ97FCCuIyEPtEzulChdJqQS5rCfNMTg0FGemU5NCU2Qq+2rWaep7BpOQB74/cZXzw
0z/c/Lch38XYyTEgz1X1AGDZKIqOiXb5RaYxoUGWvzR4Pa2Ku2kA4fC/oDz75IU2B+DGZ+iiEvVp
f//r6PlQPDwQ5YqYUERH6a6HVFQzT+gmEdQ/R7UqVnNvH6qR0X25SjxQvTbLsZBrD/CeZwEGgIY3
/VyCvPdWd/8Qq4zQaXwEtmogC+/Ddaghkmb6eRMH2k38U/9pMdEXRBCSxiHNfT9rGf+F+CHemxmD
+oOjFnfzAke01glX+o7HWrO135mn/VEpQT5BWDv6bBAHx/uip9Ljg2rnnLfAlAKyMLlwSeX/HC6v
W2ATtpJsV0YtiLUPieY37SPgweisu+Klgdq+wmJKlyY2ntbrDB/DEx5+NH7z4hDI7kj1dNsfz9Ti
0PR32UCzdmDyKGOIQ8tNHAwaWlStqIhBvbn7YpEuL6/h2ily50OG8y9l56qUVztV5HfzTeaQgfYu
UuQRHCXTkWI1HkXTPuXCUujVn8T4L7r1upVZkDaf4d/9+B3cV9gGzdiI7c3Ezhj6xfVgI8WFV21n
1iBPYPpnQVf/0aICfm4M4btuD/EIbi82bUy08auR/usTiO/+1gI0bLITcb1ZRq44VwkTl5U+b8gY
PEqcsVHGU45KbAFt0FqKr1E9ICQiedIZl5g4JeXiNI5NXSae7Tscfy2+EU79v9rfqmWqujb8IsdL
1YIz7xJQ2lyKZERvMVc50y2GXoXcSWrPcr4qcjFCSJVvBA6MQRXqMtjoM7zAKgNDL+JL1HvFIwQk
xFfRgSKSCzJtB2j0FBWeqwA3KGxcNlrRbLbfOrvPUIn0jTVo6jntUk8TBM/Zuk6znoK+8pOnr+na
YRwMclxLPWLLDr+LY2SseXlOTDZMjpXInScHalnC6+Mrxh9cb2lnQp9Kqc9H6Q3g9qipvl9EJEl3
Y/jd0tMO4ZUMpQnD5q+2WQHT0BpIOjfEZSPZ/9dawGkk82emvgCGjZFHV0n6jr14J5m6hLa+qyUF
dhsGxBzYEHrarofRbrx31My+UUO8UZqAKgtMZrMU61ioTXhEuhhsrsCzEpKem+Mvq2p5hXFbqqVR
iyqxRY3PNJ1FuCQ4Be6MF3EZpYbE43mRepqAJ2OYeDd25KyzJY8GOaF/Gbm9yzYr7psmuSQ9H83z
qUsr1WDPkt090lxJiPbGY+6nTCfLmJPBpd22V8Qbeq+1Ap7S0/XEMF7OkSfICK20Q/zqSiYA0X/q
vJ6TDloFvM8vFo39BxnFKRNjZFc/C6kfIcIkVMkwH4e1F4IUNC0sI8j3J6UMYX3TwEbispDz6yMb
UNaBl8/pbyKpZFZFnIAurxO+dj6HAVB3alZaCBTvxen9BoVbqoiRndsyEQTWvyqYCBgOVyFZNYVQ
1bmZJZArovlWudr7TkjL9ofZNEMMz4t7RC2eCI0Tag+QitciZDFEtT3wIszzspK54+nLHUrxCEU7
ivOYKewqIudt88XHu9u3PkdaYIZK+MGI+2moRYfO/Bd6taODOiVN1tKnLRmZEtGwzhq0XNBkUL+K
sqkABssOcMzsr1dML1cB4IU6qJO3QHVBvAVuXGHJb47x7Q6hRj1h10PZUB3KwwlJhBI+meGp2DJC
Iycxsw3Py/NDtR2F2Ssqm9Yl8dh2YZyXBs8QkW/DYoDDOUpuESDL91pn/RFBMDuyDdLfxX3S+lXG
H6LnG+JqY7I54ADveLJzUde7I3iYn1XBgyNjxoJu06RlgAkz3w3MpOHz6D3PrPbseJ3d/M4Wr44k
8FEpSl76/IFxuNr2UIHsHu4YJ74OogpxOtUtfLPaKaMysDQyDB0toPXYYROCk+EC3dETfiAD+8mP
lXsckvMHXLH9olIJCOOpt6dUIZDA8d2batUc5sarVxzXL/ScyQhD/jETmxU5y5OrMLMEkwCExy+f
OKWMIOdP3UHopoPkp/OxTS766/Ff4VWuxOVZTcVWhkC0YhDrPtNAUUC3HV9USdkGn0KvfYKsP4as
K0VAHEHvDR2eyicsbGyteXcIQpFRcLLD/2mGjf66B264rjgrYkuGoWfqoKNKGWAiKSVS+ALw51qk
pM75X40AWBxx8+FJnZk7R8oMBixgo3BJSEKpdSp/H9lAANz+betcwTs+M7yPfOO8VNQISYtSXl9B
RM56mlacD1CcJvM1W+BJ53LkWT682JqML4tSe/bKaaXmXh3xqo99PQ/M2k43sUNBVYLvZIUNtGIy
aUwI4tsYjlXkFx6LLN988mqXPbZ2NQVGKydi27hi1HLjj+20Iqw2EYWbUH6cGQ75qlDGbaWWHhhL
tSxnqrm+2AUylblAZF2OSX5JthT0xjXtVoCOrsKkHa6SnNBh/T+kQPE3GDw0/4wXaEHm+JD8mCzC
5JsFRjFT0MQtKEz3aqqYwf9s7wM0XEkTfXImJ1e/b8bz+p7ROeyir2xeLIdoYuXkPaMvVeflQ5iT
RIH5QBS3s4En/V1dPdef9qtIPQEPRp8HtD5jvhnbU645LksJbqoJBuD+HNmR0K/IrLqp424Tonrd
zEQkrSq/h3glq1CSQCpj1Jyq/ppR4SC8apqEX3TeESjr0fKr0uT+WOZiEl1r4AO4EwXDuzHEzwYL
WmnDbsFf5o8oID5UWO8l2lIsF6VwgbSVzPWDH+wvc5kmKGb0SlKCdaSgz3BREQ7T5PCIPw5DnqxC
CMQDQn0eYZKZg+t445NEGcEihB58BVvLhQpaZClpU+mJpB8UlAPt8ZAdTSaaGnOB6c65C5WKRa7n
GoqTvcJoUjXHGqjDiMlzSBkvy7hE+hqkbhKJEys2W08ZkhVfLLh8+nuPQXxkTZvBN+lTMaP0ILS+
/aompbf0RlfVj+ZtSpexH7In53atLRp2rEzy1XVJ4LDGKer3Z/7oQOaPGKkfg0LOjXCKLCtWIKaj
ofKw+KWEkyoloo3EJ9xOOxdUKmFPUHChXhze8G1CIdLtT798VN9OhRd29/I53teXEYR8n/lNdiH4
0e5TFgLx35ttoIYBxtpoNeuxscb8RDm+f1XVXA22IlXsYWamEtGOaxQySDhbjm48ALcmT4lr9+9E
4WoSjpguwd37E20362W/JHJgi4U6cEJH259IWt76ViBdeKLfcYajXkntiHwS+CUNK4i1yEjcYtGY
HQrM6sASA3tMZTYetZDGHHIPvP9dLVW0QgjkiaPrN4Pkv4G4dXrWJtxRIYL/SLj0Utg3epd1exhg
WfCWCoF+GnSFXcOYRQ+0Bd7Uck6ONyK+Xi1ZQ9212Z236+9OicuolVcrj8XGGGBWDo7VODma7xAN
Xmd//br+paGp3dpqNdiEZyhdq2XUi9zXFNA4cKN5+vaoTTUenAuFkc96Ksy34xjaBTfa3qRoaEou
Eyy/P08xrhcfEl6upXTlzhV9F0HE4yFadZiROGqExhcSgd6awv1fXVBQyWIMsjcN5egB8JemrH63
6we0OsEnDOcqkEUFVFfCypKblFudpFGy3+BdQ5upHnoOwQLfJLItapnu/LyBt+tYi/+7/yTxBnSw
3jw2e3Ji9safog/pCtj1nXGOcXhvJa+QBLI86KbAhuwlHSV/qQI2OaliUjTHtpBZvAwzCu1ridKS
8y38gRo7ZV5Y7EE/dBwuMrb4CmbivHXc5ZGpJAEzczsh0TR3MlWCj9NDCWMypTt4Q57kA0uJFzGc
5emV7G3YmqHO6BUW51seRDjhYIQqZ1T93TDhe2WC3q76CKO+csY/0ySJO0/AIj9vIm2WOhCImfzb
6AqugZUx5o7OjvURSzwmjCgrwhsU4SbpBewOm+vliJEMhJPCkZzgYkjUpuapz5WcpwxeF+TaUU6C
vOp/VyGUYzRRA5tUUzEtFOJlEzm0zMyj+9B8giFB/uEPyyKpOdYLN7OlVsdUaN58woetl2Y7pF9g
FhyHwJ/DTDdUSCmrdFE79SQA1CsbZqKKS33r1e5kYLznxfBuOQClKIm4L3Ce9cTJgVGvtkzOoTw2
O8VGqmcXmVjBpSM8MvMtFCdmkLvHQD+UEMnINvTVGTrfoVWINEMRwgHaPAINM/BGQY9FB3krMbWw
TJg2MM9uDwqsCg49pYdRY0OE53WEgl7O+5VbIL9ACeFgcgd966Ieh05xo9OYpJ5yjQd/iSAQk1Li
RgKpfF9miSpKLajIOS8o2kYA/RyxkVvSID/qUUAQ7i4LIRouuILb3OG0EQXwOiYohO/jSXjSW6v3
5lZJ07fsxvoqn4UbJRHnlw0MMYT+7weT+2b2pc1u7Eeah7vSkw2oErYbu3rpZm/7hjhqtgvZRQ87
rm6Q9NDLujy8Zvd1elemZp+MhF88qtEjFkw4YHYciby9tKJ8KA5pFqOQytPjcILqyXngk42e3/ak
0yFjgsBpsOioajMyUfDWMIvRqNsEo/jN39gx63Pg0BqwAXrLBIkHv3PxojdMFU0bHoVsEdCg2Zs1
c9aDYFDF0iTHd2g/ghvIAPYvRHJm92a47ttrXbs1j1m/F1BxdgsZ2YgIjGvF0neZ+RxzQN2ts1Re
qytTuK3dsYYzExFUtssQI/Efxb418RkXP3NlpOyyRHEr3wk/iEiSis2LUUpru6tCAVE6cdmTM0AZ
/0/+TAXYjW6xp4r+wlDqVsLbMAcX28v4zCsIbr1RcKFeXCYI/HaKoRKjhRi9BFEyhfT76kZAnC/9
RwD1EEqma+2mlxC4Vt6ZkwlmPolr9/JINUT2mp9S9NmoIA0hdbAC3uhMsx7PgGPSMRHnVjl3Rk46
f1TnG8qY3nYlnnPcjD0BCetzzWJTM53yhKurP3bge52xhaEonishGC7yDXjNdC6qmUUKFxZr7k0c
F5xD8fm46FsZpsfVhTEKebHi8SsmqZALk7R603/cZSlAgFuisIN0l2gkYPuU41YhMzaPpgQUGpyZ
bYtM7fIPH0yZoacl1SOMhelUb68ewsWNjxVUVj53xhGA/p61JbtRvpf6CRAw2LnK8mENSuLTd5Qy
ntHRN4pET5Wtu3f0q1ZFcbIG+Ol+xN4O1fts6ztGk1mjaLl29/uEXlURVX7s4Y2yJ9HcLc/QVGfv
WAAUJ3bcQt0+4PwUnK2/gVcKPl6cbUf1VdoAXsaUEesiCB3UOwspeAwh3Qnb9eqs+KzctxdOATC0
glMnFSePOanWWM3/9y5V6zelpucrODRPJNqMUXdogiuEB78k2qaZdfUOecOL1XApQzFaFRK1LrRt
OeQi9A3kvbLfulVxZx9/dpO3Mvum0XzVmOOMxZewE3+QbJSV4raDBcvioxz99Kn7b0dUhiHxIuoS
5+IbBFUgZoByHZXT5XB1qf0wfikai36Ah6iyibzWli+1vNMVJclKPH66G7Ym4aZfFoLXGfrqDXeb
E/hHQdwIK2oTVjsywp3wYtPowADnqvbXedz8oTXkoIJqrE+vhMnAGQkvu9pz/fGXcfF35Vrg/PMn
mBmWZ+Xs4N+tQ32OJu09D/KcYghhsBaqWUfDcF9mD5bqGswggdFP2PTTVwffvHnTcJjo4cJPIFjZ
yD9XDZky0sl+VDdyGdYxwOrxSJymidlHgAPo35uHQw3EXlXG+Fl7+0SsQ2iSqC+m+ufdhS11Wkrh
qIBpmkdCq4EoQf/e/fDDM8n/DLFH1tipmJEF57NT2T1gH6TY3rihbKreVqBygqnw6dHrIE057Cn/
h1RvBMJSA2Mp2Mqrz0F5O0sVlIQCsMJIfsSkWHvOvkLHlxCYFCAWogMooiB6aPkNcawvpY8+x2TT
OvXLSYM02sDRf61oXEd4nhgwqr0y4wbYtgc7zQejakst6g14ebvnOgbZI5XA6itft0pevSRnLkKm
CfDYA0NRjvR7roHCnrPdBqtJcQtyhsRT1QrZvFqFHhd/fgwRxSnSHU7/cdAimfzAZsK84t6wyDhI
cdcBSYPhlnBzC4xxqaLukpnCKVxX0BrfO8gEGricS5wJ+S9YYTw0r560ZnWabdUFK1XBeQl82X/O
zn9tE8AjCS5QHpbokAB/SDqT1vXf3P5UtgzzPzNns4EZ2nlzZeGFt4qfbwAs/Q8EjPgu/fNuy5mP
ZWGY/YnSz4s44PaUi9U9glZ0s5s38fi8u2OjfoYOWRgZaLG4iqWbottpzqLDkmcHCepLZ323NmpJ
Yjno7thXCEYuUcwRj3s9/Zt9B0z8KWbMxhT789fX+K/JXvTd0+2iGhr+LnWsshO7h2Fp1Kso3fOl
NbQbcwKzwGMXZ+2pntZKQbez4YEAA7NJYrwaiXpWBQy6p3Cw8Xq2IvH2UiS1TxVaPQ08PqgXVLpN
jGONLOuCs4WY7ksJgbUcz28sJ/c6GCML/nnWQ5I/SRAVpJNtBkyIeoB1mEbcN3iyCbUHBgf9KIVX
x9ELNetBmukpZ9HMTNRM0fQtE8svODHOPE+Rmrg09Uh9voF0dIHd/9TtqJ+Yrx6KTEL85LgXVD82
Zm31NkM4BlIyl8N2t/wOo+ctWZfK7534lx/jVLitvrprG40pUttytwX/NtxlvYWF8Iar7CLQAVrA
PXv/tCDOBoTd9NDyu79gJuiSYqaWfpkuiXczfyxOdBLBi7lNRuC7h5qrPBcOkpsjwJj2L+sEKK0v
sTCRGXRfA0Qn/mg3SsNTD5kEj2wAZS+squ41f5MXu49DNEJ7VdQQkJx1SY2dTLX592Ztz5PVYeDD
tWF3EVEQXhycXq5lQMyaJSJ1Ets5IQY4k6E9D7euHYyVA7l2dvPnkonC5JfNdfc0uMT4GXzrd5c7
zUZeFh7RT05EcdLMrljydX0aqYzULfG5uFmxUYrmwTjWuJPu4pUsnXHOQWuvKrCI7+LdcWEkrsN5
uHUMhoiI6drFwiypRgOo4duO9v0XdVQ2xIMVwenRuoy4Ns0UZe937ZAhX4MqfqL6DMJc3uTZdKoq
seyeCffqLZLdQ8bz6AgOLIzCukgKsyzcrrd7KSpZEGT2wYr69uHFXJt1ksNSviz8mcQ46U8083qH
FzBY2aQCPno887HjYDcAGV6lOcMo0EpNHqaf1aTlUmxbJGiQyHVWn2FBLC0V+77vv/88H7HgaZP7
Y10OmcAEjL6GwmM03mwpFe021iNJ98OZSHnl7Sp13Ia7becGx9wdckbPChnBZp5jHx7T9YzUNUxO
pKWs9b2citwacFJopHvgsGQYyS6IMZOvSfMta76GL6+r+c1SGnZWmzXk9JfoKH7/iz3QydwdWGbh
dYHaOwHN1hBo7mfy4VssFcfrep9vEs9ChIKHbGRcWxUe7f+fhZ39x9GnXMDYK0T9VNgKOltVrXMT
RaDsSOe73irHjPvJbU2nb1yh8jX3xKLVBK0GEkQw6IQifn1FAtlGySupTOb2hVTRuMDerRjWMLGS
buMmxdm3qH2uOBXJmXI3tM0ernNIHCd4ISG4RMW/sSblN+2OzHJZtVvg7sEMbyc/I5OUZktzcR3y
iaGTFf/+hup3FrrNclJ1JF0hoFyen0GDyNuwoCH3oXdu1+g5SjxMa4lpdAKWoPy56UgitdoGgZsG
+8cmWMsssdY/NDdtxRTTymThl7PalcDMfOT5dg736wnxcpY6BCHJZMEMxZNcBR3IZDIw0jAfrrw4
F7jrc9z3gGkuI5UdVt5V6aJOekDDhd9sgOxSWO9J6+xuKiL62L0yUicC+MYY7oWwJGNdkc0SCtV/
o2VxP2DYrILZLVzUapYa/Q1zd7uy3e2YsjEoPqAaTjNAmbHkA19S2XM/r83cDbpJZxAqSvzV7DPy
fPIcBJiJp864Je9I3H0n8jDr8BfCDNlxdMUfzBmwbtvjun/y47Zp5FUbm5u9OU7Zl2Dch5IA7o+l
gExByNEJxWTJSHMGiu7xvm7x9ECBtnxPXg6cwIFjxi9uZs8EdvNxK25SSm+9nIgyxv5Nak6IW9Y6
HXulXWlkSrcLtHAbbpeA7C9vSpcCirvg+NSqVXX0tbXXEd42Hm3FRVsIqDQcMELIVLXQksQdfzjK
u78sPO5CLkmghCE+PrsoD3i1p3CXZgVHsVoAiRvGnVW9DLHDZ3ZwfoxvU/H5MJGdHp4ANoVRV9m0
e4sLcFozoBXhTjgwjazcU1eU5/P8HQr/pgKE+hI8Uerm6vFyaOpMemVYWocqO++rumjq6jPbKJ/H
4e1HZmD9UjCCTt6AMzacaMfjt86+2oP8oi5bCyjlCBgUVyT0VOyBBV3dTBrTkRcuiIXNEYV8T6M3
q76LbjHm5DGbLZothv8MzUUVexPMzNN4pxJm3UxKaZJtLQib4o4aaXcdQzN0ibtVZt/jNqA4BrlP
DEJy78h7uQ6WASi865phrP54xL22tffWUfbxrEHI5E6FmnF72ZJmU8mAcgHjVqKSfxa4QydvjUWJ
rexakoVEv/Wo8tFsKShVV2JfHX9bv20UDHp8TPcFE+fqIyBU6y7k08Rr38VVpSVkDxiPPr5YzgEd
d/C92oRli/pQf/c4TBURI95IV7PU3xcP+IVZ5BheVLpY9FcLQEFDzleJ4MPfoPcjOG9ta3Qnj5dv
TeTYPeYWN/BmagyQFGiDTSsZuZEPE8LHHkvcvFWs9RxVbTKqfuSl91LwBjeCqnulNzsnbTq1MSxK
3qYglt4He9yZ/kM37997V6cURE2jhfoOD92u5BSHko+RFl1NVPEFIkhm9wuw4VqNkyCaR6i6mzjm
zEoPnWzkKkGCzEW/8xysSXOsFrWjvBYKvtgpVs2L+ncO0bojeg0DP6Qk+bRBSoIC9OUnnrII+r1l
xa1qgXTBVjvyIt+ymVzs81JrXah16Q+XfDoISAMIvQST5iuEMfb8xI3uBVH45yNFc8NhekVREEuj
5pnfWvyicAbN8J4U7Sl2fV6rqxYmInqMLlJSjTExmV4Hx7T9TUW/0fUdaPNmobULlZGNCLIYjiMq
hCpabR2HTbibzjL/91T00j0kw2QRuH6wVogC5W1rvL6ShJaRLUgmJZO8dxIL1qCco/uw0Mlu66ev
3TAJuroYmCar88tmahrwVp2fWO0D/Bml0YIpVHGo15rhOiWf/VR3ZiDNuD8k09xnSvlxUL6AjN0S
lI+CZuGmGTw471mUf9nSQIpFFhL47I7vqrtjKNhxSXXudE/jyIAALfNL8NznhvROZCBTSEg0Jpf4
qrXFzr8pNEQeJjAQJ3+Ou9VgT4Ll3sf9fNnPn888m/OkrjUsFtgLzRrs/53Yn0Kn6/C4142vFxyA
WXUmL1vVbUWgz1IyhiWaZluyMHNj0zj1FC2lhYprBEZWJbnqjbYQqAmSXGjxFBo/0lpSA+IKjt0P
VVB5ncLawLApM5q1tL1qyCCWlkIzY6//myy6TfS08dgLJQVRlm+6CqhZIhzMkleZSOfDqUKmOuAe
UjP2waEZEgTL4SbyahG0y0r6r2cA1KdaqPsurIr58ZJT5VRiXo8gM4h69MVz1FpPPxBKEXThQOZH
a/PJBru87cCcLzYfj67MiR0jHaL69hR2fJxACzNsj5HghChYwSZLgIRKKf3NKnA0NcqcTny7RgPX
/uKMYcODCamJEjvyRBdXjJgl+aek7DHEoUrqA/SDC5X3h2vPLS5Icp+daBnVlymayi3UH0ttVDBE
NF2enWRLuaknO61oxFI6HEH4KtOoCCqgo2Wo1ceVcn+5/1DiaxQRPhB2kwmAnIoX9ew7MKpxqXbX
OZaRZwEP5PSKRbu3wXJD4/IwB+VJT0bB4Y0DmF1IyFmN9QxL44tDLsHeYKKuK9HUXlTFMDLTESK3
zi03baU62mLbSGRd+ro7moUB0UuVnN1n/JKyH54u/n68WIUJuhqgU3mI0JU75jYwyTBiJXTuhBiq
mWMWpIb3mGFwwR2AmaI3uIrLJuUWxjTezDsJuhtfxX9S3LJ8YqgXWhsgtYqIpRR4Fo13jDZHt5Fg
gB3AzsBk4AgrgZh/eThY4bA5feNDUi2WCjPAXNfP6p+n5LN8uWNxLQl/UGCEjbVkF2LhptuZtZh5
xJjQTVhuaDHnFKABwBwG/eps/2tTPpozaImrctN4j+3A5aMGkKPWf8gFmHv/bcXruqxS04h3shN0
9Uk1nF0a6NS4CVA2aiQj8bSKrQALWNp3m7sLtxJjcU/mdvmGiafDgsTrdrc3wWH81G8sRR4uwJfB
0UpjEm0Dfzgn86LAD77VwIdIDcLPAk0Uro9WK30TzAtZ1doFL6Qgv+NSdBUFIzq+yAfN3gGFkS4m
O+/UPeoOUoyVXXK8/msrTHnZ1i+UW6exJjhUbP2C60ewDipUy59l5zmXNfASDU6zOmA4VefZkgxy
8oocyBP4a3hX7Q59k5e4A20JwEY+r4Zzss5uzP5DKaipBUdl88nHLKkZDYtG1WSmVWrqjkA8YfIa
dRdwSe+wYPx1unll2KQPT3w1TcMVdVI09XmIgGh5uposDy7+YVlpDL6C+92luS+7ZaH5w5l5cfHE
/F1vbkMLRY1gkJKY2UXXRSX6CsK396gPdT/nYizIAfTrw6XDG/gDxOzBEfOfmQUQr1fW9XMfjvch
GyZ7Wlod/1593nkLrr07HZZNr74+LXaAztFU41WAFjCpTqvAaGdC9xfnu7pQGNP5lFXhvAHr8FqT
mNtgHtuGkyCaIkGrVehUQtbYBNr0Ds9eho/D+8DWYevnvFK01GpkobforAoxRsoZUfIgzB2pmJyc
UmtY81YdaMu+n00O57ROckDrA+pWbXoqlZ+LoJDHxPBzq43d+G3sp/3d2HqtK3UrPi+VaLFmwjbb
WtDKvuwbrUbT8bZAUVgWJ2P98U80bCU8iREcFUUfAKofQKYmwZsNY4RYUkASM4WSCNgy2verNC3m
gD2TqezTFdC1AZMEF4PKt/3JOdbOKB5NdZig0qYP04as2WBBDfotXsiMltEKGzNoklmZShnyNfFI
/hGi4mqTt12sZBuGO5p3SgZRxgqsnr5zJSfo+dQoIKItOrYwEkuCpERFOY8hlv0INk7Sq6QXu95m
vJTf4Wvh3u0mVtlx17szujTlSn1ti0Op9/Khado41LytYcGLu4dDIUBsYYShoS7wdq2Zfl47TGHu
EEFl17Qxgm9ttJu5A4/OJSMEfzr2KPk8z4YI4U5p/5qUceRNdKqo69STZqiQzv0rdB7VBXxmYUl/
2Ec/qvSfJ4Q24Y2p+rhpNCqHXA/1YhRoRIRUKq3pHqvvcVe13vezhmAVsGslHOUOUinuhX29R43Q
DJfOfiOSgxmhZGbWyxlVvwkFo+NJ49tUwI/8g6BMUl9zLHg8ndLuG+oSvxx3s6xXCZc0WWhFe5nV
0FyLkBFr/KTnhCVNeZXVgz8i1PREONJdQdKZgtw+J7VxqV9Lq+eo8tGtw6VIGqvCmj/taHqJZZti
tl24HaJpdRJkAynKNTlDyW0Dg/BUZj0jpxkE0gX5oCEC0HXGgUWONCoMI34v1Wve2BTj8xwV7iYn
l+sPNOU5ScMiaet28jBO0ncletEFaPHzfaOKQfyI3i7FKJuDUyyfJSZEvXiPZqXK1BSRKUFdzaUd
hEQWFI0Dl7+HPXt7/nK/8ZvvLfP0gVmFgSTY+HG4tAWfXahUQEFQfCEhzu3Mbb06aPX6mgOnbQgt
Bt1K18rLzW6YLy/QX5Bls7ccnderyn7KvOVz7Y02sEhxXJMBMCJ59u/Lae/MfcCHzjAxwkh9r1Zu
QXNlpTZ5T/5reC61CGQ0eZh5+VbaWf4ZZZClqKi53Q98UkS2w9k5llFFL5A8sxtvco3c1Aaj0gPp
aj6fVtGlydDQOnH0CAJrev0u2q1PcQp0hpSCDrBD1+61r8m72eJsTxgh3BZCwAtcv7vT+y0v0DXJ
vnML8hZqlIK/47rt+w+nIslnq6XODY2vMy0B7LEDlSyj9NIRh+mkaXUHXQhu/G4sNzDg5T8Peu57
cU9lKR63H7bioBGrvK2+tEcuXp2lLklWvjiDJxoETPXJAgaKCXC8fi/d4EfOoFu2euBV5QpLR3hj
6e+JefoWYPbHKqP43kIBz6RaYUilu0Mf460Ih2zEVisbUPihCk+1OJBxkbkyMN5XIb9Sc92YJHgv
wn25pHMfBXfshi+cag7po0QV9UztfjS9Dt8mTiRT+CAXBpJN/pcnca7H7vQTWjkjVE4xkw+Ii+GX
iFjs3krOvuVPeU9CILiwHZfSb3qe9l/EEyxT1li6uBZcsixLAgwgHqv04RR10X85xoP2b7BHIX4n
xYtvWhqaPa7NbdDLZmxH7PdXM/10n9OlECefFMWJm/3q3KtjlmlkMjjKBUd4lsSypVscTRvzzKyO
BgZ5Kqk/2wAQQIld9S5qvXKGbfukFG7hoXrwCmaUTSOpVtN/cCp8CVdRc7uRMWD7c18KuJnBxNlu
V+AwpDsUHMBudDhnManjePmtYebRkiEuQJMEutifG1pkXYXCJTGmilROvPdra+3r9IK2Cx9lSCTG
57ZHltsD24r0afQID2YS16rveDI3QQuH/wjYJKGcMqjtZY7O6XEKswCxqMIqhTRyh3OmQgv3nbN3
X4x0q5u4LlgcWyYEKtyrSkslgLWefplXhlcTX3VKikk3oGGzVbtBGV7bPvaz5+KvXoSZ22nlN8vn
2J4oG+2Va7nOmn9+vvNQz0mHNQZNSp2mfixzk+ruHg80mPBGmNsjAOYQC7ZxEp25plDOBQ577F6V
7tu/nupJmikoH517ttvSiogxAoiNe3WBpGW5zDBA20AMDhmKG7FLaNjiq8PKKBklHCdrIAnz5ZPT
FIqm5z4fsCRLp42R0B+zwVdkxcpM7rF6ps42FueT96RObrh+0ot3YwsrK15KV+ODA4cP9iW/G1lc
TLE/bIfrEKnZLbgq5GHC3U+DB/0/tCgGDoV/y3qDLTi12trR86THsHFbu/1FPF1spV0Y3T2KNoQH
uQdEmsKRsyg80nb3fUuDTRbMirEEax+F5MYrdTxQEpHF7CGgq9zULGuq27gJ0yFETxepGiy5WOXn
rBjNz3vdWVjW6lw4R+ngUi3/8+WJuUX9Nzf/hB0oGqV7CizDOmhSBJTj8oVHwfaXITk3y+Ia9tkd
Bgl1Xe45F2gd3KI78qf67IaGE6NaR3lXSwzJ6L6QHOD377A5UquRakegXLJ9QzVqdOmE+EkfEJyT
4V/iqvrkF88KigH7LjHCClXLnPlqQ8+BuvKuWcyhHZ7U0tkq5/D7uxWy4VlagAPF4fECTgVuE9UU
HrCzszxTr5RIF7KbFRJBmfOn6lLubqKQ3Ou/3P/n+GDdYqPkzsiIHUqrLb3EKJq4vyYExXyyglZt
RiuwvK6MJscwCrcfqtG/+Ongj4u/Pb6UUhDtrEmt7O0utZDLvn9l9XELaQLlJLfPlVexAra+3tr/
7Pl8l14ybepywOmNf3DLVK9oGh8LNRiw+/fMML233/cAhbXfslf5POOH5T69oz7AeOaSWy01OjiA
9Bimid7D20UXwhNXM/kGqsHsjjOfpBtRFiBpFmamfYfuEQNa7YbArkWDiDzAqtJdwJitJnwnxZhq
InS3PaydGIW0Z89Qg9EA/25nBgwr4fg+f6oEOK086GNFGyne11NURCOk9eHbCiLLC2DZVlUZMi7+
EgbjPoyOBjpPB5uMEmKYAQlMEj6DHR/0MKMZzd5FfEzDXvBknVD2V+SovrlkXJT+KrCzTSfkO4kn
E4UW/XeTu/uhfIMGlNuHZ5f6LMpwRotJfN09d4JzYhK0bZBTDxIAsTFBU7tMps23KTlY5dk6Z5W4
+RBeRSqQkBx+7WtFBgFCeqXmrTE+nmIHN4PpSf5P1BZX67z/6ZPEhv/uo+ozzjgBUljosqB1BpK8
EXrDq6Z86w0g/L3DjdGxC/Ev4DI3EkyuKbbftr8W4y+kYGK80wNRiKtlxFrslIqxivSlJcug9sUb
imJQURigxInMUi6LSQiQAIT5eohJjVKgPupYdyoi5i2YtnOCIpu8yZ4XsgIvSYJFDgWWGll4j+U4
7u6tCHlFxi5u/q/itrAvDxDcwj+WyXJ/KETHFIRt0BQnCYn94aCF78Sy+0/dEjQyLlLrn5+rYqih
NtpblyyA6rhfNeMDmPJIRsCsUbXkUQpHszEAM995KSTvx+/n2pr/oFj8eaUtSKHRQCESfMLutP5O
ooMGJzPf+mx4RhyYvWmJCwqgwtetzsaF5cPH1OZ32lt7V0ztp9F4Ra/Czw267BXWOASCLKOP6ARR
+xcA75vCVFgfWotX5KUnh7FkJTJsxIYVMCVbgCNA7lFbBSSn7bf2c/rjSxG5xT1jZIE+4jtMeO5y
eKa9yYD0rWbxJB0SsoSgLAQrWgxjNmiVmJ4H+tb6l+MmEv9Dq3PU58nRXMu6hY4eEwACo8QePZaA
JaB3H3mKPdw8FfWHq16beRnhjB6+3A0AWfrhDNboxw9VHVGguV9PpPMePKW8BDjm1+obTO1MDO58
UGxy091aA+SVNHex4IvcVly5PhFclAXKcbdgOCXmqUxUiY4bCpNatJ8uvXzGyubCCaZPDfKeMmCL
kj9vx87aR1sljPH3R1O2HdKKcPe5SIqRxc3lw8J78sM8MlHbng4FGvXNxDzfYxjP3J0dxTwLar/P
GxFB1Yu00FNkEbJdG30qPdin649JvUJEkaUhx/CYGrivDMI47u/k130pHxl46Ysxh90/oPYpVKg+
EiPDChAz30/w+e+WCJY5zZWX/X+dioRfLKVyor10g9UaldKVAYNMXBz7MLR/12eRAVbziRCFFy9d
8KCp+W+XYxopsIPUryXq3nCgkIVsB2vt6UoBSBC6ltGuyQ72l0+mDfcLFe8aZrP3fhJKDKqYGypi
1WWWyoYAV7/WuynkrbBg23a8ilswF+MtmfEmf/PWE4GrwcELf+cB57GgEwMySe9FAto/BhuhmacZ
tw2ps2z2DqcJ/DJJxOc1wSQlfZSWGjYSWcaQCoTHu0XjBBH9cMD2QWs1qdyS6ortbNzMI04Q57B7
6r2ptJp3QE031npWhloZ80xDvaGrQNnpjTBQTppRQzh9I+p9KJZ9oTm5gUIb8C6qGPol8RMai04k
mTd2uWEHYxf3P59MllZqqgyVaMoUwfy0mbmmz/06I0knCwSc/10UCvd0swr8X0OgW2TT18VXU/cb
WGgfYw9hs36/OgCEVaklGS+7rQQttXJiFoPU5ObDQSqkK0Tk4BvwD6/nXI+LX5rx22YBTgPjmk0I
gIe+w0kFGK2zHcNDIopnIX724TEA+4ww3jODy/tAf4sTWCC/4Qo69jPKcmIE6OY6UQNPWz+J5FgC
/3qSrJDRwc2TD2o5B9WEsLS27//NIh8cbBy8tyIcIaBAooh7oG1Z/3q0Fyf0Zb4mteff31az96L5
k9ocR5ZSlH4XggryOwaGr1agLRMZeqF0ek09hpSw01gVeTkqmbYbiuU5L+yMiQOgBi8s64z8j09z
y/OeHLpZr5KkJ58PqxkJbGp5G070aA8RK85X5M6mFfZv+UOx8yfJjqgbEaQTFhucibhg/S/TgO4s
bQxLG5S5ImMEgbWAK/PZRG/LKiRKBdQ2iWCcTDzj3GGYgoTEKiXQ385d48Mhc1Q/eWgOOld7F7fS
GmbaTqfhY4HfwvPhdPATSAUTeBn1fw80yi90tD5+cJfrpUjRH/uMcMTynvjyuiN3FwGOpH/J+OQ6
DEJt/jbmP1doipcAtCWBCEsjfMC40BqtpAaHErx1sABC+HmPp2idk2VvR10/18TCE9CN6rE1s2KM
IAsY/nNoldQ4/mUWDYqaW7lynw7aetu2sGXJHpc20S/2rJ8r8plKt/bLcFi4TI1HWgs4g9pU6Knh
1pKBZVhx36BYghntrVfV1ZoPMCthEK1RIcqVdhi8Nlddpng8u1pJtaFH6fHujV6873DnmOsD0ggs
K71TMmQVl7Kw0vypB2CMWZnvRN6QzBVYdYERjV8E8fJ0Oy0/VbJuJSb1uI2+OCxM13GUbVxtNTS4
0jQ1/NhJhaqghQJUvcy3DPru2oLF3QtTrB0IZL9rkoQHN+r8NrR2rMjb+nek95kHl/dyYx4bPQdK
hsi2XWdHMQOSe1cydp/rBb3DUxWeb+T9PmJb9MNz5/h5Be7iei2/rZYrHRet9QXFiIc9Qphv4X09
7+PDyIDltjxm+FArp3Pnr0t2uWaB96Dwb2DPXhEzs0+1hFA8Ca69YfgSpjDIiUZ9/iAuuXw59sW8
F7zMc5ChWwCZiLgBfqBq+dJdFeTgcT+4ef9Cz1T7p54uaaNxnR3JCTBlvwYqUT3cS5ZaoFqdtcgu
gF3Skshvx1UMTrcoqNHwao6OduPpr02Dd45MSzVaJll6ROt2ci1XW61g0W+0mDNqHwtrXlog2Kwk
/rC2rdVVIWXXZhgwiNx9mK7l5afM4jwLM58cfESFp/Cts7E2ZRxr8u11F0HXudBH+zJy3v78E2L8
NV7GS8GCga4iLir5OVyc4UUFLFr7eAE2F1mVRjyRyykMVvlEUS5zzje+FxrfqnJjny38GGCphlY4
QRwtQN+3bjymuGE1wOd8ZE8UsSE7sqTGpK0cv6+0uN1YHTTc+XPp47jpW5RkCrayyHSl6dAEjwN4
MYc5ijcZbecDbU4JXkER9OS6HFFy+Ur38EyHRRBsT3ZByJlkxXllXD0UAiZ5xYE/PHMF9F6ZMlXA
j+wvJDG0dLCw7hu16lYWRTqQjAPeV7vQL/yZT/+6ZYn3XLKnygKIFHzUcAfQ09BkblQMiqmdQYuR
QzW2pAOCNE2sY9GB4tTPpBsaUkSriFNLEwwLYbqtX+kYjBpUoLs0MGNLQWXEbys+lm3Y/I0OPypG
ZThcnIDF8CWEHNQ1UNNQ1CyH62ofbgSCg1nY0qXbFkapaN6qdLfRYTt/v8cY6+VgfFzkzNNtuyDH
sYOBcjZd/Ps6Yb4CZtsnbw41zvdqxQfvUxIrtwfkBh9wYTssC4L5hifsl9BQqe5nhngjNVF+zGKY
luP0y7OOW18VzbbwL4LADjUtk3DdG5mF/O536AOnBrhimNzPPatTY6PyNa4kZFjcc7vlZgtd1zPc
uOGRBsyPKlL2nsY+LY4hPngQ2QvW20eFP3jS+rrnmUYwknxE+orUcZNtoJ4xzaobhD6xOPu258Mm
7888YpeVYXtngV1FDPVg2zROsKjOhWtVnMLHcsaPvB8t6uHfsymQI4KeLUYKK9+ZW+G24jrcZ4x4
QIYmgNxQqRjlBKhu6rXhspgtxyuu6GXDnf3qUz3CfszC07NTQHKWrnzxWApA0easSY63yLeZlhn/
45PHw+tXYtsSOtOnaZjYroO/rbbwtJU3r9gEC6qsRpdPvnejjnUVbEnGlxtBP1WRfxleY5hj4qcH
j0Q02Pd/eWNf4PC/1bm1cuyjxnmA5DBU0MYHWSw0A/9oNPcPoTUzpOkrRv8ludGT0+Xy9wGKb+9Q
KWgJUsaN6QF3m4F8LTOt6/dxWb+GHfMS/BRkhuxoltLrxzYi6sAkSf5g1KP2MtfS7kmXV4R3lQXk
EGmdz7NCdon9JXDCUpSFuCWC4fs9Bl/6dGh2rDcyR0kpvs/bTR34mLg4nEzUJ4p3PXyGWzEcrCYy
rjSpD41C7YR4vrhtWBjiq3SzrDyPOdSMj3ApRWmloR+c6eR6PnlbuQXwv9JFbmbjeyH2AqXUPSZP
JHxiEsi1EQrG0tKrBx5rj8PWDCOn8uT6tW5L3U0OuVIcMwq3NgqvxymOWB2+6S8bsT+ivbLTPaTa
cjYcOmCLZi7cw23WAqI+dXg0F0lJ2Mm3lU86dl02VB7DMI6RkPTb7GBdhbfVBTocJbeUYlcxEian
/XUmq6u7hKKQw505S1usOZhkOXAekYJnhIzFZsBqrDhBt+KfWRKhvflMo+ne2TkfQH0UIeun0iuZ
Z92JH8G5i06xO+kBoiQf9XN6s84qd13TaqeUTGWkwZhH2E41m1bkpBZClXd4Io8RzYPXrar/v1OS
Pgi9c50RU0AoholsCTWFzmOeilNDREM2L8Y9ynNNbT+VUQKQM+NNQqe7iGwV7NXeBumyWzRNqUet
u2AYIcrFohpi4kzAc2dYJxuIz9PD5lGQXc8OxwEzl8uiHdZKqmjaqHEUJfMSytSKZWHJwqICBOx3
SiSuMrLWonwVa/LHmOy798WcNhuygjKJuzr2LP0oe8gHRv0D+tBGobiQLv4etrZOS3rk5Vs6eQDx
chz1/bOtKXxKyBaAowL61Dg3rWYdhZCfbYXKvd4gWHsYjhPF4aSDWwCb6KHLbxgeFPVnL2ePK8O/
V9uo8QS+7RMHO/L/VLDP0xBP16XEH3nX4yIdYwiiKh9prsdyDa5qvvKOyGyCqgpSgubjOUMwfFtF
+ReJZwwsXBTAfyGukNtLWHlFExcHw65tnE8GF1DUPVQADL+rt1qPeiitjhE1dr7nQNR0kb9xYfeK
pRJCRxVsv2ZOvbDCe210LDgoaTkcOv+iPvDRXhb7vhgRCGj5tsMiXXk9x8QIgE/5kEYy/4VZ/ylT
nXVIiy1VUZPr7dz9tF38ThpDwfpgOVYfw0xPh0MfiVq/b82MXXvabdUb2gNlzxtmJCqbP1+mHvcf
vdheOrKs8prIVhNHt3aKOHLMGTRoCxk2hFhaQOe5DGNiDUeVdDXd7Zixn9MkCgXDS/LEEAN8vicX
btXRzsS72d8ipq5H01ATYafyn0+v3qg2YtEIHgV+YzQw3PI9mZxMr00WIDebeI4R0Wn0oUf/tuJq
Kk1KbIpCgiBJETzt2iPFFBwkua8OsJ8gLiNsUnvyB3Adimibu4vI/k1+0Ko2jPMVL1igKj8l0xsN
JxkqB3+6nPUXDsTDtAv2u6naWQBNuNxVJwsImB4B9sU7LGq4lJvIjJyJ8vhTx0uPYMctwiusfGp1
+Ni5XAAYygHye9LvJWul08k5xtEK2R0/id5p60H2FwZMroP/jLP37K3lk6/PDC6zlShq83MwgS5p
FOIs9qFuI//d/fIt3jHuQejpF7D3Xa2v1/MaMeRmMPqK5eglWQk0zRdhEIAZ+9x0/0zUhpSdBzPf
TSZZpmuG9EZoMwV60kHfn29tmBNSSArKwhouLER26mVUob3K8damsVRTcBiK2H18azSpiRmvKEzC
vNLiYaxe+GM6Htu1jsdpzeswB/c5Iomy/CEhpBfunCohdxp+TuoLfxdFbV6lLdtjxG9zn2lzrBGM
8kaH+qew4pOkEAeXhReC6eaPETIYnDvqXmk0BFzw65vrzYu4vyRzq8LmA4+v1a1FUzNM2RQcRYe0
uc3E5jflKIPiGaz0vn2L2OUTFle12kyUJxQVV5jRVlDVpSzFDuXtudvUh2HfuqTz7FJCkHIcyjOs
JMSFtz5qgKuC5Yu32pTybuphgqqSaUjwZDOoMDMl3nnigKsCahANxrNI/5ysmb1OOLy6e15lHR2f
FC590yKG5gTu9sM46kdV8P6XwN1vrqoqNRfqhPK7I2ihqpoO5aQjayoX3K4n2x9czn5Ipie2SyYL
qsTjDlAqUgc7QGf51tifXdBxYMFD/9J899uGfEQwD0Kdkedo+iLD0KG0N7qstvIJK9OpU48j4Grn
6+e7O0WDEICw4iEc6hEi63+f+2yT/0m0tBHz5G2md5QxShbqFOPaKkETP+F7E3UiT3uP8S+bOz5H
x//phzAkjveqYTx91QijWWPZZOdEvrDGNlG3DRgWmSOu1R9MVX0KqMbU/CJ4/pMkdpCTIMXC3Jaj
b2FfVmNHg3ZRkLNMyqWgyEBPlOi1IZbt1drfARzDkb3/8yDJzuKnnTgWIQntN2DezKkM6b2JfvRr
UgZCJBns6DrYerTn22UW3vb0IRRPpPMuVkTSURcGKvcQgldqzYjtycAGwGn598alJgjH+dCVi2gl
MG9yW7rJnYrNVQp56kxq7KtVYINtr47/OvrHMR3TUxqKzvCqy09X3+yhZ5PS5PfYc1sNDsLSoMCp
PVySFYks/LlS/wFv6MZGWJkImwxsMjXItev9fJ/bwjoirI3VDrI5A70Rz11Xj8SdnRT7w1qBqEfw
4ckry34u+Xd4b69KjKP2hnYGF4cC+H1ao0ai0+bCHA963fYv/DDBaVy8V7PzCJZD4HZRS3jjbx4K
wRFg7pCrciXpTERzvurq7b0OtT5l0cjXp4Ua62HjNoQrdi3POKiPL1Qts62i7WEHieCVb15cxm5H
ThC7346aRBNrmlseYTt8QBzMinlBSu32CA6CHy+n36eVs43urg4AKx1/NjWaLgAESoG6WTLhWiUr
R/xVj/3qDGLF/0nSiRdoKkWLiGYzoXAi4ptr/TujPOMUxcRl81n/PXFYPT4hvAZ4O5gIla1CHIEU
t/9i/ENWTufCg1b/XvyvNb+8qC9A4BpM7fF32DeoMzpx1Q3oKHmNAsLUOF23YlrC2HynBnC1Qrz0
4m/jYO2ju0XuRY/P/8S0aMPPrytvgU0lw3J00zgh0ogc+GOBW2RsabMCaVW36nSKDGljecJCWHVg
PQ1NI7UVkCDYs9PANw5kKD7PINuRvxdxKqjHk4LZEQ1O4aDTOyVoKzVo0ECwvLcLBv3kvgo4Yj8e
zRGxBF91hgia7zDTotFHaCIFgqhnJxXAwjo3RZ9DLhTeVYROIG+pOxC5oHR2uBLRHtYunk2J0zMt
/YJTmm4HesCOz/NJkDhtKr2ljAii/n+bFpJfcg0CpxifNPyeXBW3pICoezWosP2SFpM1s3uGIFRl
KxaAVBNA8buB+pDe5BjSxh0457WzqTa3v8WoBvKZpWMIYgBlmfcxxBqe5CMuBzffIOiJGK5jIbzd
OKQqOYVDzYkbSHmwvroMQT4KlYWhh093yEzFgoJO9++UTS6Np5gt9eohybiC0GD+zOmlGzxBh8nX
u2LNUPWnRJPOmvikUOrE8JuH81pe6Bo2FfLhR3+zrwWFdOuj+QathsnsLAPRbAGbnA1Vw5uMQYcQ
yJ4PQ2emZKBp/TA9sAgBALUFbSaX3l6l26puL/ePFgKoL6QFXUvXecg5qzU/JBJTfFJ2vyMRt+j6
l3UeFZmHgA8HjAK5diaIXt7DoUisGSBsg/OrD2Ojz+ts9t9zcMUgfGNzLEk46ncRk265tsb3+O0S
4LzprX92+nzgqJ4m7V7RdhYcRRy10LpkjBoltUi7hm3qSsm+F7sSxWaBgM0MfcLNr4mYYC4oQ2Xj
cLSwQEJsOswKVTYU+oO24wBWnFrcqRstvaMljQDf2N7XhcnyWRcxQxULN4gLlSlbJKzm9QTzK13Z
oGFNahgecTiJGr7IjbE/iLs+8+09yGWbjTbp/LI7fwICtpJNGt1eLcw4PH7JtHBm8GSOVr3e24hP
v+i84nQf64fLduZcJu9wkhkw1tk05x2OQNT2wXQPXTzS3w/6mg76+12ngNB0ffq8S7YndH71eLkA
VXSVyRGgmmtNHAYgErX6UAFlISNSV0Z99bVWFIRvOs6zu6m3TPWyTpkVqV++WPhxJnnptsKZ+S2h
QZ1+NHu+v6IVGNI3PF3j8Kr7lCboAvgJaPCT4RRTojvKNOziQx4SRq2T6QkpkrJmh0Kyml+lmrDp
QhO7jYchT5A/EReqrQ3WwXwBtVHTzA5zSnQggR7ABnZs6nkmcxkDZz658M2ghZvk9I1BgUueavAO
2SKnEADHtUSCOTQcSXTd3xTSL6IqlzR4X5Zil9YB18nnGyjDx0bd0dmjXHy0sw2lsiYeFHm94qVF
k+Tmq5iit97jaPsRjHimvHLrWzH+NjDAnPbssoQG3vrkIubUY2yH/Im3Hgpok5eCqZVL0D5AgZk/
7Q9r3oWjqGiRma45zSTqVP417hPEzm7dz3oPzSrwCNlqsAszHpQModrs7p/waRfpuiJnjpaBOceN
GyCofG4NJxYZ6350SE2jDJp6MkYFBX/dqB1Vqvq3KD1mBccvr8tPXf4XfuAHubTpMfrg02uE7WxQ
rV5ZrRYO0DBTpQw5ryAvl1yre+Fm7i9ijgVSuDDOKOeC6l1W5zUrRSv5im9ZOJ7oRHZaSNPqOulw
ZbZH91NmCfboM8LC/eZYxqwq/Rlg0A9oKtd0eUYmy3UCOXP04NXstRfzA3yyPXHDrFFh1BGlFh08
T/1ABkgHWmLh+PeBOKv/BZJiafNQ8HZHCtU0Wl1n7pRJd0p6ZFTHAr3rlS87fxxIse01ROVHi4gy
340VAm005yWTPTun2nJ6qYXy8ZFM1QlCpdXUQOpYb9p3FKthLXY46OuKxVrAMcv0xG8n2uYDHwps
42BfzC1qAKg6bHbHJ/A8Uv7FOGRCKxd6hcG7xtw1rJH2xGs0k0PGToRWL/omuda2HpKkzj1HH58+
QMoxdgtLHIq+6TEZt05C0lJLFZNfrGd68SVmlqvuTFcmCb1f+Ro3A2zQVuutWDaxBpKVEu6rcgqz
+Z+jKv4Q3XXloAMB59fJaNuWmjR0Ha4ef8FIoBTYlyKcT9oVq8pcQsrAjMSfBkeVJAthO+L2p1qb
Sr7Z9rdItD/wpJjd+EvvwFLHf/MF+gOD2JHP2R38xsRSZ4g5rCq7GlHETYP+4CxwZCBtcaM6WMeW
5uTYgYTx5v7B/Luv20ETJjEEiheh3PMJ+yGOk5ZZrxgo1XijTwFONvO3jBbUyBgOC60VK6BkyB5y
Zf6Fb/+VRsMi5/YPhkXV6/dC3NJ4+MIdnBwXurJZE6qaO8Cy8+fN4TrEgDdP3aHSn8Hw5jPF+eSZ
t5ZK02brA5/McaRtvtFKpxfL9CAnMxW4l+w8AfQyz6Yb5eMNw3I51x1GUiBMIkJPWouTPpNZuB2l
o5lsSJ2PxgsAYK2rFheRlUbAnAE/8GkaYtppF7RlX6/fNFCR5u3VPD4oqnVqgFxb3uF3TnVwGn6+
Hzgbe/V+H67d4AeZfPIy/BRO5F0yKtq7aUm8IEEHwQppMtSmCctr/e+BUh4E+QLFZYxWr6W9j8HY
OT8jsX9TdIv+7M7Xa7vIGHf3sPHub/l7iFc3gpIq0IjaqwcQkMrwZ7V8+7ZqnbKsnL+LDg66hk9X
RWePpMDHK1DRNiIs8j023znSozYJ0+VGFhg31UVENMDApY4bbnLH4wDAFWK+icAtUtNROW+PliZV
SfwFRkERuM/fsxUpp0PSs117Afo0Ag6iJrlcGTO5g2TQB9ZgVohozbD5CGfTPQLtokPRT9p1KSeM
4S18vvKbY8ijLTAu6GGX2HLIC6oocLPqlu0hB7G8Ee4xmKtKgnMIYL6fOJbtF6DiaHFIBWqArXoK
uzh4jm+HTDQV6FIGeG25a0RfiHAUC+EN7my5s8526Gfg5fC1t5cpKvJiM+Mr+cNu8xpAtAhD9i7T
ObV27Dne6hJIZRPwkI0XAlMBa2qk4ynRBQ5S+1WF/r46oZ+PiRNIIWOvlCjRsSeuwVj4O+Esu4p9
2wkUXslYGNNHe3diNYO4arIcdeGstmwtJgK+2brAn+X+xEy89BDv1r51CT0AVvo2MCU7pj81pl6S
5JghlV99pfU4O1t8B2QZ5XFiPTBMk4jQqMlRMXwei0Tc2mcGtWhhXFF7oPMaOnqFtHKJFH4FKOdi
MtzNV/59HewQMEccDk5oGCgSenuaAWUsnAE0ZmJEuu9nCO+ceYCQAFVleODpD2zHirrXIdv8Yt34
Au5zAXnOp3iW26BsOCfKR3UYrSEVJbHRHj3ctSrcLVBS4qqCGK2CpCddo0WbLHi3/xuHuRJG1W+J
R7+Akk6rsDOsm0G4JbCTQ+Lq9laW7q6M6bqA/ViAgKh1qbjPZ3Fn8DD7LRIEwn+mc6JStGWDNI2Z
gA0uqEZktEuKDkBiq4veaY6SYFf0+VFAP9nxpLUD+Fd0m6DqdKbNEGRVyho5b3ztDvLxS2oI7I3I
HVosAJA34s1v68nIPGeVx4HRAjnYSCwcA2B02JtvMvasIhM2ZpY/geGeon04r/0yV4NzSVJBQPqU
+zvEcP4cGNc7LP90PBTzGkHxLlBSek+eSN77061d/rsaSuYyQUdCxUEaXuik56n2TNZnxNxzgjS7
U3qkAYsIIWYoj2+R6SNWglOMszX1tBTkAmiGQHQ6ukv44aJyvSN4oin65+bC+qf1RqeGw0CECj8U
CqueIbOsFcszArxjUF1NEvulYa92+2I81vA3BJXnDFTfOevTS0lzjst24hcCvbKqp8vzLhMJ/Uhb
Trlk9f2BSZKcWrXlVEWFj3NDgrLBChffoo0vLWguMDouYJmBL1PRbIBGNXmkiE9MSDHrxGyhMsXF
B6iQGkIh/+yzTKwYO4+jo5QrPFbnDTwBbD55rIMZ8nHfEjsJtFJs1MLi71GkIFTDFtNnL4EeCyid
3A7K8kQhQrmq3+7uli1hGTw8iIsDiQkJIdH4rCf5RC1GkNIM3D/s17njjWJ9FYTvPqHcU1Kqmmft
c6ePOR2PiaKimvuizcGbHqSZGSZ716SeAJ64T6y9GmpT9GdY/kAyrcwTzPMozLmhasOXFSzYX92T
X2brYiezARKZRW3QBnlEJk6vicU3sGaRXg6zUxKt1jMCp9C0H9DQNtXlw3bSkdQ0vBFQ99xWFvSy
ZhXErTQZijxMybaYdD1ydWmo2e1+UGGbEFSuWReznJsYvxO+FTlUiFjiA8Sq8GfT14bofKXa0kuU
CR6J+DkQSaIkMUWTrQ36ytooXq/tuDwWkNJ+bBQDvo+YlZndsQ24zTIIsgfw6uiB9FoCqwLNiJzy
vac1kBhjdH/jeznEXDOXQ7O/ZVFw3i339WoVehkfga2XwDMjiX3ToNvxCYya/Vn9RdfdUGwYNlwO
lmhYXtAz1cj2aq+o73J7LgCsS7cDnnfWrGxUN/lTVIw/1IAV6K7R3JR5uhZHKpaxU8F88TMOZjwp
i5KqxkaRGq0LyKf97UxnQOnMIeSy6bDsjlyTACG8WdHPCmwBeUTM4+p7ut0Fw0Uo5ltlwUxXYZcN
mVAwsdjMmyJVvTD8aOg+HU6KR87Xtz4XVLh4UO8bNoe873Dd79YCtb9fpeWkfr6DwCVQs2iJ01z8
rrEDfBwhqtsF4Xgmiwcr/M2Cu2s9PF2S3sIc/w33TbxEe3BU6TjyQP+uXkjXFqUpKFcCYbhJcOJy
YlPqT6mDXrC+6gcQY2+ZWpjrdCUfuxUOCO63abesUGPxx4OW1BmqJURfzBCgSZ7ZjrL+hdbhgGLy
1YVAIKCZTFn/DwUPZMRB1sDgdJvIxakBkQoWx/twLLfS6Gqai+xgukTSQp8dSi3/eAMHzg0Hs76x
WXPEPUr0ZrStOpQxOnEhv3BOQumrYSQHnt8I2yG+YbHt0KNPiFpw9oJA0UMQ1S3bwMNuM3H4zV5a
S5VfNF53UavsOP6ABrfEze/Wddq6keL0KvubtWdOXuHjaL/M84bLEwxXF/T+mKBqXAyCTFfJ4emj
YZlM59a2kbyqYw8mJcS3t4x88dmV+crHlGEYdAu6crLPoUx1U8Ni2LVDhpvLEv7P928Zm5rjqZDV
aEQ7qG6+TtMuVrnGg+XLpsvM0+WDSqEiQGdn6IjjQoD5qplDJdgysV2yK6aKsnQ4Qw7kGEhrjkgq
o8CCL4c14BhbiYRX8didHY8rf7WvO5iluiAhCZW3/dVbvk9IJum9W6bpkZg07yV6MPWiaw+1gQF8
u9i8NqoeK8eF42OlephtSPzo192SfJWyEbwpToVHAahD8XKb0P5eAWiWSSZ+aBeow6u9VoZhUvmz
1E9S5gH0jaopnT6qnL4r2k0mwIXf6Ngm5hFFyzj/igltmuXuHzol+eYs8YrgPrNVNNcpdHwDGhSx
bf9LSdAXQKrM9v5F1iN8cYN43JwguC7brLXYPxSBf+lQlnY3cIywx3k07qd/P97RI3g6WsOjwdzy
fSb4dvZKo7BS2lxy7V+86o76Wt7W7c0KtrSQ10r4CAdt+Dn244jzijAID2XTHpwnrWY/wcQSKNta
8Z+/6buCowRCTTIL0XP+JHuSdBqjHGxZTL+P1ng97I3q4ZDrjElFv6Zhg7msP/yU/TRf7hWeJqT5
tBlKBbggAF2SnyFezOShZOfw5BcJyymQoB+IX4N+5+ttXx6cxVjmI3/N7Pehj+zJbGSiMJHgbqgZ
OIsCRjsp8uSEYh0WXjkkIDMr2AJnkJrpXXAIz93MIpJZAKZfogxLRAelCzuHSPkOpeykD6BrI5uO
WSeczO8sHVNoQxsOke1x+ydTYEfJIXMn9xx3qH4Woc/ToKcvv8aOo48c8CXqmmxr4dGrzPBPOs1Z
AOR4Rojl6OcsYySh4W6pD0rYdeL7vnGZuHrzaFP3X7zUu/IaOns3SLRNZRMkKMEYsk174zxv+6oB
RMe3KDDac9SoFePz6LDeDUO/uTh9I2eMTgWQYj3E90h4UW6/TYw4yyven/PlpCR5KYaqHXDKL+tb
aFqK5so7pMwG5OC0cB+clNoPpRY5jb/T01yJuN8rSAHk5XDJaZMb1krV/SNG9PCgt5uxtanlYHxm
6EFNDD12LouBOodDnfTrXmBEkZ6m2tf2wcq78PKDiaketdd6nGf2wtOsdDl42JJuhH7FXvNcRceW
iYECpgZmrl0YMUtsAE7Ak6JR7aJb7YCAo+L1GeXsUDEjxt0MnFGRRKZEEOzwojFXLtpJhygfr6Mr
GmgDlcfYdr+mi7z4qLTpFsq1XCcHt7WGUUpNYsq+S7l2y6VrOsqCp1tQ5bL2PRdrOyf7rWs8YR8T
eoIXmTq3KI6ppd7p/iogqgEamUGDFrvLihrFQ8vDLZbkfzWQc5p0yMEcpoHV4QiDPAy93guotjPI
Nv48ePBr0XUHmOf4gB22zdQhMRfHWOfVNYJqReARD/3EIxA5H/enx/vdDmMI7Yo3jv8tuqf99Rxa
MkhLAkORdtzEDjPUgFzmh9P50JFO7yxFhkZ6EzGphFLCd8ZA1PgwpGl4GSRHr3TOe6fsUh7kdAHf
gNNBi+UVjNX26eMVavQZGIlt+tzwZhlZc9ZtGx/kdJfnjkheiBpr2br0HFILbbhfn4UgERU5x7A4
2vFLI3ElpAxshogVgnv5G0xmExqnJ6uomSUAiyCJcF/NPX4fIUKMkXZ0y46XPwL/Tuq4rUOkim0F
g2rZjqFsKPpHQM57KNiIrDKrMc+qDf0mhRxuzaImIPXWiKnIBwFr0mPutXiVlSkgnqw1xuGa5G7p
WHBRSIbh1ZIu9DIKnT4nW4p2jIDTkS7WaRHQxhdDea8PkR9pLF2FVxlQScJELENppvb3y4C6Ln4S
BmVPctwdiia+sXPtBchFr7rPCjRSIjL7pUdGpui6+VDS7R48KMkWzLYiHQCJQ6BEEU/8uDKMfk8t
Zlnky67b90WylrJzVY+7t2kHH3c6M8Z78m6nHI7gTzXfSAZjmp9jj2eFNqv8NiTnhHrXSFJ3G6q3
ZyHoSiHRAu2srs0/85NEVnpz5vUgRkoS1lx8vuL4TURe2/RQJ3d83dwcXCT3VShrrOJFcufd1KXH
fRhZ0gpRGVKtbFYMjoeOfV/BoCUCmkS0Vjjk9995S4tgdiT/+DW2UahQKa/JzzN1BVzcNN97DFMB
TX0WBn1n7EUeFbgrfoxS5rNatOdVvFKmcbLmdXfNsUW8TfWt2cmYgr/kD9kYpBFEfRpht97AZcAm
4mSTtGwzLgi1AY2SUcavLlTFiJS7+8hPtwZilWLD9ZGd2lO2AbXLF2x03BDzGFa8L9aK87iMziVa
bsc2mMdS8JI3cM8lD3M6EP4d6gI0PEDffevnVZV6DCo6qkqjPTzOZt5MLlnrNtqZNBmaXqS7wgtf
QmPP0J6fThu5XJQGwkgLssmenI1QMftwPuTPTrNhh1VGF3kRIqXZnTRsS70C3E4uuqc7ZiYQXvH9
mwZEutsKiQqBP0LD3IrBntxJU+5Z7EYDd19ZGpCQZ4TexJ0RpDW2SFl5Un3hovkWArPM0iCSxWLM
uDqTbSXwSU0z0M2/mDpMwEV0RDpuEF3c7rmA5eULwHUf/t6Uy3CcS9myAwrfgZT2E6vlXH/5N0Ml
Lk0wYhLHxsz67XOqjdiTNbht8As+8R5SbLFmyKM81TiIYBLy/OYkhEmiXMa/txKtZda7IgZgxuVy
/9FTtYio9BUwlo1bwvomSvVYxJwuM7b9fh6aBqzy7YsCWtzJuMG4PYdKYPhTQWUh+q3hu1VbFxcm
mHXkfYt3KY2BXfmblDD3xsUtEjHtg3rGE/H9Ti6ixneoN0P9rDr7pWz7hmZcbPOqSLJpBazibtI0
F7idbvoBuYF8dry/uQfd6RCcUNHCaCbHVy5Kdd3cACxPnLegT0jZGpZeYYi308uhGejD//A/SgnS
u40D6sp1qPVI8UL/3XMdZS1IaU3rmjXoVIVLkiEqDikMGHDD3v3ADKEN1YqJeicipugbTbl9yyeu
UY7HB6t7hTHYgp13P0QwrIhaHJu4RvQcxzo481d3i57aozXtQm+QOYWVjLEWDMcFIbbiPqm5r8i6
FN469xYtED5HfCzEiQa0+1Xb9lNJqmHh0OAGANbmKMr/bJBOPsoldj7Tq2naqeXWFjPQxw46inEp
tMLiq7oPq9YmqRcOlu+9aBwZd2CDeUGlvAQ7L5rbJK5XxJ/TFXYHb291tanlZbrU8q/X8Liu4tZJ
vb/xGkQTUOKyc/WdGYRgM/IWU4jYntSuMnv7NpnMM3/s8X0fEkug8haNQq1zMSdOfC+2qq7omoAv
V/rGTKIidIwdn/IuQnsrzfHmKqcQtCjOCZC6l3BWiWgj5Apc80b5nFWkFgfnfHk6zeDZzmlod2/M
1RfBDrGQdOzcJfXKt09WJA+nP3gGtso7MK6cdDLG4BpqIwEia2vbJulvuSUMYMeq/aEbyyblxaVQ
NWj4ysqE2mM5Fl8rXPBdKaeltr31PscyUm/D2Q9F85tkT0a/iYleS6ZhB0Tsgaunk3s1crZt5JHl
7Cbn1iUvqW1G/UBIbQSmkw+nqLuqOiMHrGq7+RAHkrvivrUmG/uLmHrOOAMFtI610cTTjx3Juhwm
3nzvf946DKk/kcpAIBZhsgl2T7s1QqeGTYLtHO24oMf7Q+sZLXChLxnLWFq9Aa02I1Ghn7WM3O3X
40uisa9QZZz9SIPeAUZFkkgG1wcwdkMZNNTbmq5P7rKMmRxZgc4ZACBeS0qDmNt1BG1AZabAdDyg
VR5f7HO5xnNVxyngd1Jp6R8oyJQRwp73VDBplCiiS12oqIZW5fdsOJ9tzIZaPoOC6ToMOeK7NZCs
/gE+QTuSSnSOK6qxbbwAD8iEzWJnQk7Ov+XOZ9/yO0BsZ7prs0jpV6qT1f4sQ1ezynXadtOpZA9I
KxC6ctAYjWeLi9NBOajXwBiFyqhnRIAgA8wKeQ2WTLMOTQSlKCjyckOeNFIVhOETnMWBRG7WMvjZ
hKU96fHj34IaMxrp6f2ExviFMcSaWTlxjTwjgNBx5BFsOkX2Is0KqFwg3ri84z3VJYi7KU4GEOVG
ZWTO38TfSNKpG+cZb+MYu05OyP/u5w0Iu/jvY55v8jCwYGORjy15Y4OrTQ0i3jolleC+iyxfTKFI
2RzA/nndOK67qOpN2EI6K3juC3dZfdfFmxRS1N+4ceUWB930nsuzHzan0KB72N93s5tKngfa0UsI
qLHcqwE1GLUqA1kJsgGsfR9rl3WA5IIuaLQOdSkBCvDycGC895O3eWY2CBEvNtGn47ExjkUfXg9R
cJIMq00IH5lZjlPIoyPEaealU5l3kuVVHaBCXJseQFSrTZxTahWHgrDLf9QujexKs2l104v9z0XZ
44a0K4bt7eCacSYmiHP3GQSE3H87I8V+DkOBbFJwO2NBtOMWGWyIV0MUCkcaonVF0daiGTzjgDhu
gPwoy9bP7Z77/oAGwIUqJ/+NZO2FdhBjLDSYPWDAloMQHZalmBZhyji6XRJe+cPqr3Ajx2PrNVxr
m9mWF97UjTvEROIQfGa8Noww7ymsRBIkjMefPse9WZyZQMA/8U2AGrUT5Ljoc+8f/6WgjEoqltL5
F8uVU00ugnFShVk675x221ErB2PipXA8GzHM9ZsT0du1doD4NicwjI1s/iI38KPyBLoOL/8PbhpR
feVBZwZqEcZpaZOUajU0t2PY/QVERxjFT/174Bo+6S6Cfrm9YtAuXS38nCq/Wx5oD1cCDPTkwxtI
9zGtyZ9y0B/aBTMM0px6yPBTxpc8LnHNx0qJUNyThUkE/L/pgDQIgebpUVd59aZUWOOceEyBnVJZ
3QX4taKgi47qsrk3/KXRf3tcV9/acOkSE2zCzV8ivtquofeEl+cNKBC1ThyHeIN6b5nu05vEGM2B
IpF3vg1jrYJhCcZtG3wVXpEKDYnb3JEL/S4W3TZoP7m2T7S5WmH+7lJOVq7+YBceYkxotPOvavKy
Tb+R+c0dMjzKmT7xHwshCynwvLlqFIm/lYUwJr21pj04kpCnADmwCEBg0QpE8zlm4IBrqlogIidf
jSZDcUqCjaPaReKq3PEVrmejHs/+0FdBhmS197aHL6ziXeS0yWy7LxSaJOgW1cHJjtGGj4Zlft6K
V8pzQMPr51J1dVVFmhAFvjY7T/Ew4olR+PeKqLseDK6krWCv452hk6pmROuA5IXYqyL9auR+IFSw
xQnb3O3se6fFZr+0v7vxGpEt7fb1iQH/GDCPhU9rrtST604W9rm30SM3+uQOI2QisT432Bze7U2H
po31VHFh8oyvhjWp3q3pOGgEp6PUVM7NjtflR4i+UMG2qHu3htmQ+CgAXF30ycsgfBz8wcb8GiDm
jF8DvYBtMPrL4twxABO4uo7F+RGphCHLBm086sydfCFLlC3II2CAJ8i5tAOR3AKG7YX+RdW3iKp5
zsVQXyFgJbnaAHOl2NTtOnHR2Y6qM22KRpsht2u50mv/c/Y+8U0fHCvfbDfiZuPphQhXcVsyFEgT
8IdxatxJKh2sJHkQv+08zoH+f1WoxBeT63GU1Dy4cnsZ0R6WCLkVSya8fCYoH7iDefNfRaZvTpVg
MjfIApFV+QD1f0VxEZ+iZtrcOLVtGJ71O/r4a2QQshFaCKDIbOOncPl5xhmrdlx9lqkzZni/gZ8A
a398N67OUT2pp0JHHqZrmeHwiaI0et0ZAmt2UsHKzEjDbFEpqC/4uv07hf3Q1W1UWhQynQsJNjiI
n62IuG/6sv2NglxuxtEbSngjs4VGZYFVrS5nNiqd/9iHy7aYfNCS5TbPDfOgeZNYcD0b/9MgxCz8
5eAOzfbn84U2oqy/UTYzZ/iq/MN3vFDAwgBH9l78EMEsVRoQDNMWm4HG7KvZ8pFjFimHC9Y4nest
y6qmogU9i2n2TRGcfS/XquNJ/zrCbqI+8e2NoL6gqvRaYPwVMpOhQzGbLGyQZqnNAnUbGGYaQriC
sTc4Rlj1Rw13fEnCkSCfimECgIv7x1GleY2rYWpenpNulWtK9Hr3mY3nH+tPkMzWp94QjUo0XbCj
uG/mW+GbsypoZQAe1wuC4harAJtLo/r0I1Vn/VhA4uzdIEV4SchA42uVZ/zUqbaUzjXjNsABv7Ab
tFasIxFqFKj138fhbpieymWBrUuD4LRokuAvBpgeRCnIWyH9OdDoAE+AODiktWmlklWNT3yaSu0e
H7+jVb5U5xjXZoTRdSZOC0eCA6T+Z7JGeoajnuVYPruiLndH6IqfGHDEdTLu3+5xmSpp2KRdXSyn
QvEp7LYUdfuqHOgqf6v+E0TPZdA5bIjw1/u5T8GG+2/e5wO9GMg5/MttwkZ4bFH4JuYkRwTCQHNo
XvKwhASn8iqIkX2PfJThUap99vOBvGV04In0stv3IQIQq15U4y1lrw3qxlrJZyGQdaiyJVVRQlUL
+A4my/UtSMB9qV92yXOKDcb9/qpt1J+dRUWiTu5R0MY6c31zuKb+hLzh8vUpYbx1LOkKoifh4fyS
uDdjkDviCo4k3LOn1131ER1uOn3IgbfJVeZsYZzkNzGwJFwaINiXt/g2u3nA6yrQRlUdHhimqIJk
TbjHAM+Dp+j5L8ayNLQkeD6sqPHwB/JeuZ4GMbH5s6ZfxZ5xIKP6gp//R6C3rHOpbnMLsOdMRL9R
CIzY3D0l/ZYTE8jHDB+b+VDytyFDeikvBJQATlf+8fFkQI2mYhdgpwQMOwy05sN6hTcMJH4cVskc
egLyURvIRiaHaCul3QSyyLRY76kLnhfdXDediqJH9TuvT8p4BDq6OIgL21sR1bedD5ok6gBCXADS
oPAOAHG6ihchUUJCKCJYEvOvBwoLhi3rsMMk/523wLqokn3pGZYsIJwn+khWTeJhmTnYeB8Xe3uu
oVgqYy9NKDOmEwcwWOvrA6IXaLEAxwFFF3Exuf+la6gut5lXJSRJrFqPFUc5M9egfV+7J08GECEA
/yRlKi/9fQ1EvtdiP6dzGNrdrBsYnjXb/AYgEkzaoCoFTRBJvxzonvJAB6hCPKOgkmwoPdFd7Zoy
RghviWAmSFZ20W6NZ7qghyDf/pjwQ0Haa2aONYdFXspTBVwgsO4Y7XxS8TjmkWDNWXxEiZBnJowq
IDseZ2L52f8xiigw/VtzLHES1gB404MkULJLL3YLd8jdXB2nKgpwO+PuKCQpC2EZnRUoepdwxagC
uOCCwWIC5xzXZbpwxkRfYmPLFlYJoGEbEXrGCo/ZB7knY+i/eW/kd39VK3NM8rzCn36LpvFEm95E
d5zOk+tdUr8LvR5/iYdWwmCjFaRk1vPus8DSt+aR/QqVTBTs9F3uXIJUYsJkanraIK/AW21ns/1N
l3monoyBPX+I//j9bhIPMMuAR7hSHYO5XBfLUUW/T/1ctmVoTduFnvttYwadzjkKDeLuMKSAUH76
mLIdBfRK6jEtUkImoLi3UvVAD5rNVrGdQC/Gvo/BB70lNVwBOXSCpdQmFRI2o0cQqT0vn92G+gKc
/p/Q08vP9nUpeGs+mqvUDJ+odJOQfhfdCGYKKeXnZHbVM+qSMOrGHCjDEkSXDUmt2PC6FV9sKbdG
rOEFVn1WCaDU9uvhrE7bJViFe0wsojmqserOL0kyPH9+ip+CstG/pbIo7j1PeAejvMdDyKkR9p6S
LUuSnPFFxrS2b7lLOq5TgkZ47XKiB0TU+InqmDB87A5UHalS7RW+jxAHqOlrxWeLTYP8/U84z0N0
Z9pfG0PV3rue3NB1lb6eAiK/g2teL1B2U9oFWkjhNAtQGCYh3SjyeFtt6NxRt/IM3zhCNN+gHjve
UojUNMl3NW+VwgfvC4WqgyhhLbBiohfDduVI40AmZ342EbaJ/kb80bP5jdSQVelXxurOoWwvnXKk
nQYcwfHz8sMCc3MDTmUWIqq2RGshOs65vckddXiZKI61cvWRTQhpq5FRmFHr+6fux+9vV9FrLDd8
cgVmAF/KmMhVUh9MSVqcI5iY1IXbBLZXkqi7+9dUGHsFgdsbo8HZ+bDJsqlpbvGMy9SIVJgHTn1P
IGs7X+dzgv8NXDrlywmpZumz8N0+4kV/0qOdo8hvCpKdV/NVKmR+rMY1UmFaQrjZ27S+LnlpowOU
VYZeGRmsCl/4bK6FbQpoq7ebi2EUs+QkWHgGFBlX2qGKomWCjB8GbYxXMNvLDlfO3mYlpBmc3SaI
JXvFfv07onSDGF4Vx5RTCZR1q6MkuF0KueUH7SlfREs2ALVrpvrchOj7OwvVTBSp+U0qmSaQM/Xu
wILUAvT4mPH0pzQL+7y5WJml3YqezOUlpOwD5/GmqZuvu2pWQNtKK6Ryx57HhPD5/eAb0KxTrsFK
g2Z2STZWafhHZv9MXwxNyE+Kww/aF9tW/NEED8kUjB2HulBO4DQ1G6DbfvUz+SOdEgaPsRmGDAUk
Tojr+KCHyCb2QgCODZWBFs2xN81sncuKbLCgo8hzoWieI1mY/j7yPvuPe9X8+JTg1W55EvsliV3Z
9S3nLj6NLnxaNJGK+/7TgXsUzPl5Xbsa30yxDH40WhUCDtouBNVx09GgcWrXov0lfZTQXHRXIkDC
FUfS1ir7hKMOKTlmve3BA3A8aGGOLzI0rgfDuzJmwu2F3oG2bhWiZj8dYCprrrnxz/YUmRz/usHw
M/LIt9hK0vuh83excY86wBlRqNWkm2fMMaC9gj1XcmRJCaosdZvsNfwBKCuLNzEw7NfauYWnlzKx
TT8z3YyXA5OG81MKnhiQdAP43NObOxwn7W6oehkk4G9d6/tLCPmgJfCfBwaYrbmpdCtlisBac6wK
q095d/4+jNthi1+WznBMiIpaAE1JCT7mYyV0uoszOb/niJd47Z1VWQkG98eU5D2BdpDic9mB2ED5
zckBuQmy8L0ecyn2VPhNbzDclZlZARPZc8HCEJcIJiihOND79P7A9HsFGc+Qd0RexDkwPxJRo7rb
4V2Ne2rmDPPJI3pyG4ZixFhmQGe7cBkIxaVCtStPKv/pgogLYtsvmSt3iwP4DP1HGcDCqIuTjdTB
8hCMUwGaDkUt+6NOB7u/NxTCoAraYZ3p5QdPGN2q9ytLvxnAF/6pMOxI5OX+jwybK8aQ8YwcT7CN
Kq1SPOr5/CJvnz4OZXL6REEuEPUicOoyp+rjy70AvCP0rr1jiwpudNQxUrXfSOIQ6J0gG4rPL1R+
wjhPBKMzu2+ujEWxB9qBPulJe0YOgY5mmGeu5d9zEIbQ1ZDIcwye47vJs1PvAXdz2Cd0NgsCTSWl
WKgYTlpaRHF01GIZDfQ1xokwIGF6xUbwnpb71wMJelsHD9672XQgtIbwyvpOrel9Wjml5hPrGr5G
uFmWsSyi+xhjsz2aQ2czeZENHE2snQMcBGh9ju6yO3J/nsgXwiOEKNmp8W+/Ku9CEJZoWC8Fedcr
nE7Wos+Zhjrsk2oPAugSZoD8BmVAvdi2JO3hggvnBTeYK5bagi+u1/eK3sXl+aETM/LlN6x9dlaW
+8i3OY/Fy51weIuY5Ts2LoA7WUcxHLwO5He+SMGnBj2wmozIv0e2UYCm819GRUApuXvZJw7OcIIQ
cU1dNrogAoZ63VHz7FpnreYjEa7cesSIP5ZcQuw6UWEIipHQt2hXHIEG4DxNZWtFPss9PjXShBhi
NhDfA53hjVqFQzfU2bYbLhvmX2xxlOhYTTTfvKOhJ0k+I4/GvKpz/8a6YR0H7bpZuK8H8BcYXvk5
O+TwAatFUG7pY8qqLT60wKhZlb65UZbV8y9onCbErIlIf2cyoasnNt+psnKC46Lo5Eh0rjM3Bfu/
4lGOl08SNGx8FJoQWKWpP9J8b6SI+TUnn9QgN+YzB1wklsyuqHGpt3vs9ThTq+LE/VoVAQ72dGFR
Chr4LuWZrIKGNTfkosQn7N2CQzT/QFbLcAghFz+QddY7amDaUuxj5TSWiSzcDUMQCpot8/co+Bmt
V+AUcptvkCfg6dhrh8ccq9EfzVJ5gPA5chCAjybsVLPF+90YHHGn+NKhQXSH97TPMx5l2wg08uun
Ogwy8UtRrd+V8h+EfTisLy2D0awHUDJ26GDYROh31OPJcaabhnuyds+RxN8p2qZ1Oqba83ePp/Fq
9kL4BvbpTYDHEAeZ2gW1+mVz076fi2Smr8K9Xo0PeaByUesejO+oiIo1mzXadzfzweG5Ok81WF4B
d1DPZzL+xN9CfrX65szcqX9Srjzu3UXOI8aIzei4w3QjecAN+lKhEC8OM77Iov6TH+LjkfNAA4uQ
86PYuD7i5oxiLnVrA4ZPjxqZDIbSVK2+EBPpSClcg2+v8vb8u5Hy+jI9YGJhG9C3Kf4P9foNK9iL
eeT3K9teFeXbUbvlLw3e+7gRWUqx8IN8pIuBPwkm+pdbDMC/DTbGH9FkR+EaiWLEDVt59HPnKmFo
oufOxFRpB/wL26+nWl7F/uNXp5a5JS0ej31Se2iolmczwSX6427nf1ikBmgSGvau2ABeNihwHq2Y
QI2pau861NG32qN38r3Pq4JKXRFaL0Kllchfk5/uayp53VKwhVgjDtAoF3ySp5/OSAeWajilHiVZ
e9cpJFq2Zt0jUPq7ho78/CAX2MeHnQfQk5YMlJYhzj4kp2nWWpaEg2Bm3pc1zkqAHqurZnr23Vum
mUP0OEM91LQqBU1zbqTzkDJKpPjvrtFhOZX87war5CNOGuUpZQhXSbdCRwAwvUnHebOCL1ZQ9TrG
RTfA27mom6NkotEtjSrnOl1zRJGXLLTk1ZkzsPfVdcG6IMUuWI++MjEle+wgZrk25rxHp+3PhXYW
3ek5fAzbXv+M29/AOV3ufZktky9qVs6pgZWPy2n2RJZi819IYqVHv9gG7Q/cyOEA9bgey1R0ggXr
9dLnAK8pmvypCIC8IwEdukjuwRsJnuadRfN9lKiJJZIBH6wX0UDwBeijTMh6dXqgdMr8xcadhbTr
6Lto7uIOkokBqbOcuQQQ3uEwZKx8byhDvAHlMV6OAXS/rfQ4VWCDIOfi28G4xE7pv5pM7DBykjqB
VSLD1aNPDDo8tv98pqKr17LuFiCTw4Pd1yAFtZ1r2JQ75QSstz02Drv/tMVGuesne8HS9e8PLdpo
QN7qvlbvM8kRGDvLpkBmtoqwnSFAs0rHuEF73qVo9rBlUil3/xB5YG/PeXquyqfAaEB8kXMjz8bX
HIeJBXUJHy1RRILcm47IfiIncBQfxS4lSS9y28NtlH+5/jUO82l0JYqaVkuOunL0im+A7UmuPyyK
61F/Z9cjnSnHWskqbn0KQCO+RwE1KR/80jj8r/s69IiytDrOh9lX65jLyrAG2tvXnm7Qz3W1Kkyu
8kxq34yPu/H/yTubyYWQlmakMGrAzsyPcyqfePIkH8Iz8qshbKxEwc6hkrQAMQ4RttOSU6XKijk1
es21szbeZgJSne7FN7nAGcAT5Q688d8xRMLHpd7YFmflPzvM4A6XIDHNl3mTq9KnRyslhFD9x9Gq
365fqrdg2u1L1+8KUi4qzMjBYvetJ0Dbl6MbZ1PR4s9Fja635A4aNhygsOiy8CTf9itd+8ELRofr
GjkGYsb6Fs9ENrH5XiM6jKF+P26WGhz+nmmzY3owDrBZGmBBA+w69rtFCMp/s5qR5TOkqFDIxEpI
dDz5rsO8owpUhVHpUc94xL//qUjFcNqfSL+kses32cqdIYd30p2OAlts8jbe8NVQjtFsPHXfD7oH
BOaNaB++s5PI/05zV2nnb9tvQ5Rs+kLb+TSlWlX83fsFbxgsJbisPoBEsKXfsnh5vCSCWllG9exh
OGbJ5tkQs+JFMHSCkC8VXauVxnWb0q5r8Ewpx8RId1rH5PXWC9NGb8NLCSsLQFB3gDY+40FRbkwY
XYJqxcXaHcb3zk4egzKMrfqt3uDwF69PfHnf+utkA071lt0NOpwcRiZV+bFCMhAzTiyqHdmUAeKu
CcawjyXNjJfHCXuI/KisJol744Sp5L66Ui4C3y2UCWB7dCDWQnJb4LQ3EihFL0DXH2O8KkGBetb4
5IKxJJKVaGpXdPuNVl9JslGjk1oNjNP+/oqiNt0Cbr5gX3RWPPy/8uxX93FH1LeeT9OTcRz7vZSZ
ubXdz5pTA9E0FqVzZbq0tGgzMiB1XjhTeaQr0Co1Vrzph8jy1xeTmPaR796ABdmzti8OVBRyGYy/
RJOPoaNIkYFSpJ+enXUQK1xf1hLljRB4sFBGRooDDkBdZ7cYX0tSWbREInJMaFdBfJKmM7QibLFC
cHYJG4mHL3WNa30gp19kjMEsJO7g2ZNOwB1ItAV0TNw4aBDbc0u6iM2TL8bzO3uJL7t3seMM8gvz
JexdwdmXwArilBOZiczCng+rOdNZy7d3dM3I59r7hWlsSI5ZPK7T2/QCNDfRysrcztJRo1VAq3+q
1WC87N9JZ10qwkjGNJSL3kf2kbYujjJHgUelKHgM4YZ/sk5IsQw2pH4FSCgnxCvfMWCzHUHOo/fs
FP3Or41zWZQECQztVgRYOI1h0Z7F21Ffmyd+/8io4wcnRH7ND3BGNHJwK159MlaLab0le3PdfSNm
74Wd0GJCI+X/pYXmSuBaoIcarP0oogo3lSLEFV4vGoal2d0GBCCdBZC39PeChjcJUsCJt7r6dsxE
nZyZxrZoxpXWQroqP/Rnn4xkaTICr8bZ0EuI04dT3c3TSOHSs5BKT+duJHByl+pY5fvhxx0dy4d1
0GzA0KktNeTSyL32C2X3Ae4isGhSWdJ7wqAKSAA1zwB4sdDvEAIkPk6IkpxxiU0F8A33j3zlpLR9
o8aP6ecDWVkuWcWSoIIUhH1lQBHDmPcC4VT8uY5D9NaXiu8uEKY+ipVN7TA+gl/wcY+YYezXLa5V
Fjzqb06e1D7byX2QIi8J3avJzhy7FWBkDm/of+6Cz0tLrV2DvlMa+0wj6MAGeyfhh/ByTR+CGdUA
XM4iwdCPemrBOWId0hOUt4k2w6ofPa9B1CZvoCHkQcmPRktsNIe1hdjVhWbpgKi3nwB8cYIuoZRY
QUDiol7Ds3F6AtlnVZKJ4Cqo23VcNNmcyA6DQPckdpZsReE+ce34Dn+seYbQNMsBiryI4rWz59Ai
e2633lieW7us+E0pqDg2EXcMuoGOzarWhlDn/iExRlckaLJR0NdvR3akEFsI6ZNmVDwJEkFKNCqX
sbFSH9dp4J1FPIfoQWw1nmbKy6aGZodo4gnhzAaHrhGpVOLkXo2+AcU/ljOiefKQplZtPTd/foZX
6SDFROX95Iz3TUnDwGsvPNtaiI+NidBij0wJaIrNx2m+CnPTshPtXL1kfXNQOrnG0Iqqe3+9YTHZ
zJF2qoon1QC2bIeV0ieMtvxOST2DYQAeQn5GOq4AgqPQ6XhnrbZN+8bnvEOoOL7YSi90Ll0vyhSv
atO47UYgklVJTtOhccbhNmGgg8MDcIE/Nynbr3i0KOSrzAahpTc3CKE7PvtbDRdvFdaJ9DK1PyHB
bRJKcT2zEUnIDzfcgY6YFwIEuae9p16QNCuhw8FVjmPdFhxUpQ6O7x3f7CKUbemi8rZGgzdn4Ypb
XvqtsFEsA+B8ZjEGhzWN8TPlDJIOOjM+eRi0nKTnzKLkXqoazU6xF+j9sA1DaOoCFPyi/dKFpDPT
8h1nbFUgbeWgx3v6ecC7vTbWGpW+yk3aKzwZTI/ITgV+6zuPAy0XU3/WbvrGudZI/J3EnEEFsCMq
vVEBJ8IHPOOAs1EI3Xj7JY5OY78SI4b7NbagPYiaIx3hxETtqf2kul7hahP6QC5Nlz27EcxyMKnm
m8CBp2Q+s1YCeUknLX4rdFIv6JLwPu378dADKhvvabl7d1yWZS5aVPYd4VF/WZPtMKqWAy8e17lR
/CB27Dnf5QCwsp9zY20nzq0drdJmzCVDRZVMIacnfu8Bcm5jNmQmgrImAdpaA4lj7YiydU5rD/By
rrLPFt4kGrW40eP6FYWZBn5rwf8WLB5J1rYRNRm3lpzDfz0ZiXg5iabfcfWPW8ODmzrbPXizS9lo
xm/60AJDdnbNk46JJS1X4Ng8jELM69jDf/okrKUVbrvKbK6VtZX+wdFcnfa/qGWSBX5YrzzQcsKi
SsjXOZTamOgJYVwfsCodW5ntDnow3hNFX0nhVYMfXvkdQ27WSCuAYJRDtL1Hy+DYudZsIq7V3zpq
1+eLW+CdOB1FHw/N1rtf4M9IiKMNUJfw5/qYGjfJBipUbUhHHbSOS4jBvAoq7VfGx8PjQKVIOSUb
fA/YuGL8sq84CwjZD15PYMWISR0nfwTdBdCBmVV01+W/q07Fr6Id95yblSwX+aKBHpGVpRFfReSH
STp2//ihETr8SqwUYnjImZSBcws1a3AZ6m5ZxbKJbukiayZZloZ4ooL5kptPyWKSN68y3hvR71sk
Xw7rB6owao3jCPusqrJjWVDfu3K2A/2pEXvEMFX3u99QMJg8gEdzGx+a+/2EqEyyQj5efguMkMzn
JAxt6lLRf2j5mrf5LqA1oTXPStHKKfHhrf4O8yipIK0e5hJTF7CtJyyzjTJBX8ClVjuKICvgVQip
mssKR8DA4Ytc+H0nzmdz7xqE/0uzcoUcraF5zrDgmUe/TJk6uYuzb1+zR9mAw5qwL86k6dRZ1Mne
3VDkeUj9nSbzCOtQkp+IfKQBf/RvAJgOLXLN1LIzaCgCQFGY6NWT4Vphcl+ectJA6fP33amYXjY5
2XAJ7IPbDzAnJd4kZVh+OLm7dwIm5PfSdqY8bjsBjHO6sosItpkeV3ejpeIopovsAa7dKYNynavg
XasVmoLhLMczpI5bFmNfoD3L5Tna8FugrpfU48BppL2kI1qizMPop4p0U5X28Q6qMkOua5778NVt
kKC26xqJbn4F7DwzkPZe5E8je63QlH9GjoIpTOV1TUATmTiXMyA8vHi3xcbFFM5VtjLr3OXtnV7g
Mo7KOrflZCy8ctCedfrmys2uhd4QjZrQU2rNhlfLOsY+9SKEN/jUmvkLweq2E1oRViCh1l0mgvBk
sr6Nww5QPcztfmRhyHzJIVn2867lQAcYBYBVXoI37ZbMjiRImaPjyMP5f4eImWx8Jwee7TavsG1g
pMTfK//aXUoH7qDTk+R7ktPkkeXCC7JfOy7BZa8a4Vw79fsXnDSWtIa8I8dKYHOAVh/Jo97j/E96
IOmgdO1jqKQ10Nl7kqGfeC+F8tOClk41nV9eA7Nu88CLUC5/5X71oKVk5AJcrsOdh5kmEfdcfrgI
cRnKigdTnUfVZ+J2GTt24DLJrQeM4S/Xb84YbqaefP+LaqWFGcOOC4bpse+pGhtVeDytkn0v1cmP
2gfcT2ekZ3KMvcGebFSOvLkmN1bKFvXNZKGVObIAq3BYsG9IYWk5ye4+l+1ouCVXBksNbXU9LLAH
f4S2nqOzESXOaNPAE+L+7HtyWw8yTgOg3JMhNrtiZ6AwKnOnTu55ABh44mtNeHdD/2o6+n7Px/B9
fQXEJqa8Cb4jahuBqnqmcSbUZOrdZhy0KmPH4h18WN1/IgH/pFV7UDz/uvhww9YvWmJkh/ngK5iH
cI5Tczru7WN34tfqIiM9qfk6U/OjbPWKPitSLkIV6mKScTb+tyWW1IhW27ibN0IpgmBpNuOy9fHt
jJNUA3laLeC4j0RbFQiXeKaOSP3LNmxjyNDwAn92otZ5hZ+Cd33zFKY9JD3kypNicPMuCJBIwbSf
prWiN78v96P2wWV5qtoR2J3/tleYdAVEQbxPLBaGS1gNXihUSaRL4TTBBAe8rNIbNkXpyEs5QzPb
iCwdrsD5ToJ+dbkeIfRwMw/TWCl911DsgRcgyKDiz2KTA4KVK7UWgF4DLrP1NBZTvg5HHFKiKTIV
4Q/g9q0vggQYbIJl5Nc9kvb6CW8iM+6dFeg8tuxS9pvV7A0TJSYTEzuFh1UIjoDW/yMem0DcUP2u
8OQvwEFTxEsnTmiRa3lVTIa6FP0uTlqFL1kt7ENzlcq87U5Cg3o0UYuH7h7ovU7cPvMaaGCZkBbx
X3L8fWr+5oYgoBxZiMWWVP1uNbqdEGmyZ+3kIc03fs/3FCbM02OcqvO3BUJXkrXwS9coZzp1zTwR
PixmX160/x4NfDghbYoYNqn75Wjoa3fJGbAGGbfBQxjRjapRurgELCsW7EfEIAd9j61xiXw4y8qs
b0hI0CqbEyQll9reh0ZvugElqYigxw+fueA/2e4nQLkZ4w5qaJ9djv17rT82l5I50/6BM0qkZ24q
rDMuTFIMaJKf2fQEVZg1lD/QFqhnzX7QTgxe3UKyTfAfWOsqV6nOWnsOEZ229t0rmZQHYfRw2Z3U
7Lnok3O2SgWFYBy06eV2CiTe+EPOiRhKBuS6ZahcnQxn5ekrHLM8DuIBPrD/t22Vp2Q33nJC1+Ms
lJIf0ET4budGQQUdgZIWIb+TatKum498q5zDCgZGKlr5adNe6yNH3FFTkG8qYaAInFftF6P1DWif
qPgJU8XZvxR56Ca0wt211kRVza3srzki+5U+9d0xT/kLkb4bajGM5N1AYh7pVBMzW6Cip+eZWCi3
N82Yab9T5xn0FKOqLvftxHGMz4h1bvKKhy6FWf4TseIoFMRAZgWXmNWUv/qVWTiEwxr11qL6ag3H
0Ta25pGvVtavtcQ1+07Ze6Kil4xoV6IRFS8tlsjF4YP6dah5mh1MIzgWatqH/phImcSo6wjFmpai
7jIMl3QcepcJrhctwnBpTiJzy2b+zJSR+j5ZxjGL25uFNDZIJG22JTgzfG0/joM9uLlR69UXPSPJ
0Gfl+JpnBrgDjLNmrOneGJGscd7CZ1BoDaW3jAJXsdbqqlbQvUxyw5h7ZY/eHA1Z9L0NFoIGJb63
XijWNibMaHlk/QxYEwhhMNOhGK8HgJcq4CXq3GGP7x+m6skZYK9BHrnKtfbD5i4E6fANK2E2Uydk
fVfiDquMqvNESAHu+4nVleYVc90r6QVC8vx+cAUn9mKS9NdP2IzAPNPDxyVaVeI2r/fLeU0eYE4R
6rz1BeR+NW4T78jdvDhdKxN1SWOxZXQgJv7EeEavJAv8JOE2UfAf+oYnIggkMcBsDT9ECM7zXpaK
p25aYwffSMXEdz4OcnYT6qhWipPPu2iML2dAW/DASecn5eAwvEiEuD/yRwZLRPpzFrlMJP8olYRw
QTOGGY+iFH7he/hyVtkJ+h6aPTa98PZQFx7xRTkYnk2ppGnqudfComozM6UcxuD+yJtlCjTxbtn8
rZGRvAl+Td+vI4hQmtSMvA08rGSpF6IrN+m5l7A369nt3FTs0Lld9bBGZW4LLrlY2b4zcpdJecka
H/gVFF9cKaWpCrNdM6X3DTbVBgrgxI7Wkut/27Z1jqQLURricMv11eqrvYffPXN4G3zXajYkC/Tg
Ilrxm7VF8SkOOgrEPwhKSBko+F66rRPgPidY6omLSU6FUfVBrfUCQSR8zRdr+QAeneq0lp8Jx+eF
OryupJ2q/+64OXLwfw9xrE7pCQ6j972JEz7J5igPcg8Mp7e9I00DXVf8fHbmaSVBdIgfk2drEvOf
qJdVrTFad6ybt5YVAPxJ/S5HqW8pfhe6uB/L0CbeKDncMmeHa3JoAKLESjkpnaCPvOZ36dvSRuoF
rdvxYl57y2DY8QtirZYLqRKz3A08Bd5QuJFpslQq8RKu1mo1lSuXhdbbFXvlkx6wPuKVHXilQxZg
jt1Q0geouLhZZoHl85HkObS/BMReQ+yNp6/9x+jIM4fvmNqLBJZTgrsJ4DVi/+OOUjQid++tCCkl
7EvdJqUkidylPFIHgqWIba+PbdtbsukIGIFz9HwtfPOlweQaB9d4McjIzkkb3Qc5PPKUd2D45Is0
boq41N/g9BAkB4urSM1LHtnFOfVEzNanOh52xWQI4a5kDndAhYH+9omFP8K0Mn+l/kyhRqmofOui
cObShYvtoSvfX2H1RjHyP3pk8TUnMy7hApdq/XwCH/vEaE0g08FaPLlkois0lrmI5ig4x6wWDE/k
jKaMRpaOGJzAuD5Zo6hFNyxz3qqCK8zOgzjcKMao8Zjjrtw8yEB9j6tovksU6gsf1eGANlCfZ3PK
7WxZBWkOhnKSfm1v017xHjAOwtXCxcESF1uut07A+Y/bA5nY/Cf+PlSlP6SAvFkkSbiTlinj4St4
n715lu2l+6Fb4AoGUIvc2hpM0LnZDY29Vr7CO6QJoMoU9tJFqJnGhT4vnWm2bfx3G9s3Fuq3S/SF
GN7nngyuPMN5PuqvGvVy3MCccpKN15eT0WuWar1bELXmj2W+rAXYzFnhyossq+C1MvCw1vYIl2/W
nFQYJFWFx+5jzfUNhE0Ee1vV5YW/wY7j/OvvHIZtULE3RmtF+66Msj31HXKX/eW8PHc6v/IXEvB4
xBKplaV3PofWD3b0Z7zvsnyu8Nm8PqaVQxWBFTPwlYRxcfxxji+E8ksQW2EOmYi344yX3MBMTW8G
iUJSkKIPT8yf76Kpy+nus1oKS++R+mNC0zegZaQYmduE9XiZf8jRueU6O3Ggbs7z/lZkK41UC0q8
U3cNDhgKD7W8vKO8VIRNwuSmCMi6T18+cA5EzdmgRd8rtB8q8hZF77K/ZNv73Q3nmz4L2Y9E7goJ
x7l7wCNeX4rT0jMQVod9SzBl66M2ieCffeR/7l9AP0tgtXMmW/qdvfjGoxy7ByD7jDfneWvJsy5A
PqmLrTBXsVRjWmkRTLQ/YQ1KXPBpMcs6rtVfSfp1wrH8yv4p6ZptfgWSLfQxOK4gI9o5ft2pvHe7
rNYDIoBZnuYnQr97RtKpd+nhxLyWB6loxQ5O1HueadLoJ6/tfq4XRMtEoiiRhrAFXzbVEKmFuSSY
m71k7r5V2ezDNd6j4NrJ5HHdZFtZnh1n4pew+Lz1UoDpDgVEJVopQYScWkfH1lzP7OSHJq1mj7p3
UeguyZH5Hrux+f22lMgYDvQtkP+X5/S9dVwa6KP0dQ1yFGmYaGFo+qqYs4whq0sQXgbvCSo830IN
hfx4vZ3K2PbGBIS3c7VoYlqPxP585J4WiO/qz7qAl1Uy8+vY8aAJCnSeGeIvbZeMwKAJsVE6j3/X
uTPgvqVxXxL58kEb86YL5c/Y1Qn3dHD5UpqGgbzLFJ0y9M02m+ts6tKzQ33evoAQMhBrlA5SC8Ce
4QfpP2eGCsTrKYVn9/vsY/j6RfBvdNbS5bwQq9RRumaldiaD6TbSOVfoKaN/ivGUQTwgajnTrTac
gSIzgjU+rHLjlXo4VNbpTkWf4Z66RuuvJ+xEpqCI+ymzBYFhbmA3H3/Wk7v8F+lhEv1bIK/5T3Ln
2ZQOnG6vunAl0upL6583rfcUaZIhmCO0WhHpiG261ktXnzgUCRENdYucpiMgh1puqTjYPQP3bbrV
DbZR6ak87m2XA6Q+6cpDRgulhtotUChFa15Tj6H7GW0mdD0mZe1Gr9d2T/tmOulNRINi2oYpM6zj
FARqcl46/EgZkWOM+iqcu5dQvRsIFtqmSOWR87abcB89h0z3kW/BU14G25tcXygRSLCwZ7Sr3Jfp
sVPbMZoK0UFfczf/YfBxpn8TkWKyqDkBULaR8aMjC0w3dkuL/veqpiiV9POsDe+D4IAMGH82K+DJ
xOT0nrEAIHg2Pj4IUxRFoZWMUw360n3Spfa6z46Y91123pFvNUsrHOEmwC/SwE/WbDfqKNQQ0lF/
8mrq1sywRN9HUv+JLPGNwvvi60bUwap2M+y8fS33K/IsoE5hLQhmz55fOYu8+mJlxzgEp/llpczD
lD2dAZg4JLFWWkTfBY06GwJqzdqUD6B9GQK0Z8rLEG+jQEM1a4/OqsAp+i6VgEcO5MgmwtcJIJhb
JOHffmoCkaIFR9dt5Uq1XoNF60hjkhKDk7wI0DTjWlWAg6Emm0c6QIrW267+yIfvRtYx/LkiX9Jw
n07dOHj5w/rUWLUOzGHrj99X2SyzZTHob498iueTXmlLI9h1/cZeK1rptLEwX5TvgwCRbzsVmEpj
5InuwTszjrz19nvg0nZKdgaQYCZAd+Q/PYiUYSd882NM10WDqCwRG8eR/TSED/8gVllS9fPxMO+Y
sgbWXoTnWMzcyi9ou6d9ke4yVeAdZAcBrp60x2o2gkU4kYfB/JaRTLWiOuN2kXLi5LVEzD40gFJR
atgi+clB6lIN46ETeSRXrsuDEz+I1ercypnWioLMCsF1huDJCfxePMx2WpQc4yDIDIniGdDt0/gf
AZ9JxF3HY6DJW1oZNU9tpHaM73wfUGKmnqFCUc3VH1facIluQIiAF+88kAcXn66XY4DYwcODh7Ro
dB5qXuZPZtxm2QjsGMfm24ezcJJfruZVjUVL1p+gSJnqQurUAui3Yzd36JVQ8x2fOYwXs0uzFsSE
+Y1Dbz8D8nFrZiamGO/s/m8DbIS2ynJl2oVSCpdTm566f1JN44GKTl8jgbdShGULsS+PBSUY/5DO
/MWDeDxCVpPHnT9Le6vebA6Vks9eAlcIzypF7ibCCz7LTC/NH4fPbgCMbmv6vagFWG4/iSGhg+qm
RKnEyWbMByiiz0PS/7SlZmBhpOzztfj+X/21KgTVjwzl6mMcJ4JmKUnBWohv6nDEuxvjDDytmzXf
cXGpQM6HvHFPImVkXdmJMKazd81zX9gRegJ7GHoiIoF7HHjdeqbHwOTKETDpMAuhOm5Ld1LyGISW
McvNfS8weAlL717yfK8xH5U0uCXtnkBfrerp9YicQ1JTGTc3+zJjQ/2VWY58IHCITOueD45VfoYc
BQlppbeJYmjO4+co4Yb+08i/uMlF78n4QlopWMTgrRkVPaScG5JoF8OI2QKjnjjueToXi03WaPOk
NhSWEhvG9JEM4P0joGCweTPLG8Wt4BPc4h/CSn8ZjqBoXF5o378EwjDcxSOVq03Q/JVV8KUiZm6N
slivBdnc8HOwBP+o66gSBG8M4cJrbq00DSQHx7HLmqsh9mjlcLVG/wH6SXesuTAYiJ+UfGdIJsw9
SnP5wbd8EF9WfOqu+sq+8b5PIiPgNBKHgg62x6q2LTrOSzoX3UOVZsnGqn6/EM5t4cDt5G637Z3l
HTyOppAvtslUv/PwJa1O0cgrtKj/dk4501G2+MxMGHCtiAHp9KzF08IO+Ejcq+UOq9hpL/5amsJJ
BZAh7LBJYBMPRvLOXsun85J22Jg2wo9nMayPen7UevQk+m9NQSIhiAOpTWfMP+VRLMM9n5naU/Mc
n9ApWCcdqjXDT1FgtjhHDY4x961SGwabUY+3U/nDTgOxuEpsl0lq9y+7jXtZtT/X6en/VVQhsPAZ
BY0aS5LwnEx8qYx4msFeTEy7oM8lUCd4e+xCmFA9UlzMAEbTIFp9e7AAOzUjqY6st0N26jMHW3vO
b/gIhWgdrqqeYeC0Nb7Yl+OrNi0QK2Me5Mq4uEFJt9c7O3JV+v+YXVnu9qdDExseeSFdEWW09xQb
LAuoWIpO4vSVOM6lUYYHQ0bdhdCix3WmD9l7FHU+zoTvG4wewrnR3P+Thz7gyycCJyMQhebLDM5x
o7mQmLL8QQKSe9TOPdVBXqIEubVkfuWJsRhVp8Bo57VR8559NLdYLK5y+JybIRRtgcNFo/kdVu9G
6jy5sIs/YZjioIJ2vf7JOJ6lQ+vVyfztJKoX+9V9RfWvMMzgYI9pTaSWMnq3jhNge/I1gYs80Q4i
GmmHQBOnLaFvU5jnFGSMGn7bxL6WEziDMNlkbezRTMnIOI5yt/li1gX+qGw6Kr1SgleF7HfGnaLS
fOpmWJJZbtN2kU0Nsr7S7gsawne6R7lxVIwbMtJHTYY2MStBapnIsviagcc8roAtxwYtWsP5RxNK
KLnG/rNxcbk0QjhvvtWeKa4mVXf9B8EvE49acJn0laSrGqaDRdBDB7/J6mth8+z30S3J+SpWNMX/
Fx3ZKBvK6a7xpcXGhdr/NGbS66UCIG+n9Ril0vqlOvmYW8FYBQAGqG6Q1c9ylAfgWGJxeWluxAoC
k5Oyt5NlFKqCmiaP0l72MWFm0Nq5ctoXsc5jV21K6RWyN+eVQt7+c4FM15JJdMDpe1iWHHEmPq7L
gafPoMBJqrLBy+ha3mnemunLzPesQryC2D9X0mRJv33vV0J768V+s6+0foPhYjGn/J1nk8Oq0Mv4
FE1n3CfmVazwhoJIPsaPVPtiZEE1z4dwM8YYg6ENRbCw3/aem2QvhCT1VgoTu8tXz65pRszC0/un
nOb5FQtkNyanBdby0pRsYKN4Crqbrbhk8qi+Q0Nv5elOOjbN1i0wMBLM2cw4mAwO8zpI9SkNDVZS
wg3unLAyEOjWPG8/CAXOZuXVgRwMxDYoAFHOgQ5iiE7WrbDmYg///ZrYUU/+R+CQil39PzmijxrO
tszXefC5CP2FQbQlCnycExLbULj2jWPAcVQB465WuZx6KiiZumh0B2qJPaUO8q8jXmeC3qskHCWZ
MAsouHd0Bb5BFiOYxWczipquy0pzNwZclkWrcgOXiZp5MGURLcC3OWScvVT1+8I4qzF+3hcqoibV
4JmAo0bYaHJE6Ny1txBUI/r3fCQoDvtSsSL3A3QRVdzMT6Lg1RATmjD8fuHQlQW0SAyqQjCkPPxg
fHzKI/pyshvaAUH6JKfLgJIkDoNapzL9wcPr+wBtTVUe5ZIrHBzfDH7kBDqFeMTH9H8TZFkPplKY
Mt9w19eeR7p3dka9KbZkX+GLjLknXQDuOSzmhFSXjoPs6vhQxJlGgTNLwVeGjBAGOI6n0S5ZWk5d
jxdq0X4J2mcdfmd3f9rDz1Ukxt8UblSuZX96N+cwDbzkZKgwc2422tiSuAzekQORqKh3wH0A5zxH
gd6qgWr8cK+IpIDW5s/xvMYYdFQreFzJX5q8E6FLXEtyoBcNPI/NNFx/R6Oa0G3igLYkxip9NM5H
kjZY8JyZvV/I4LBvSIdcZmB3bOFtApe1UNs9ZVd7KiqA/aRIFwYs3aCBZe+FPynGEfjQfwksXUke
ntWQnzpubrNw/j1rH/JiF5BfBykOUIzz9CU16iWWlSUdse0B0WZTgYfL4Eha+5cxLdppgenM6odP
iBCvgyRCM+xpkK/1Nx0u/wNSvpYIUkwbRXRydzKx8nno6b1pBx8v8REFzZcVbSu64kpUEHECfcBQ
PYXdTi8DO9LKPUc99Vxd/MfZQF+Zh57mS2b988cANc4/Z2rKcAP1mXP8dpBI9u7Fc0/VD/5yn4bq
aRfZddmhpU07Y9QQ6f+/9GCH3fQtkhVz96CMNvy5oV23LA94oep4tBHYAj/GApRSAu9Rc4G0Q4lv
VsR7/+aROXEbDuKatSpSDSIuZgmdmq2bgLEdXkD0YfaYxzb0RDV19juYNZlUxI0cOe42iHJz1lpz
hNoqjcioyp0kOJjc4sHJSoJWnL+egf2+QXpp+U/NKTEQX4nOcKhSWSYZ48dRQILGNrFkffrfPTH6
9kIyIwSy2bdXwU9Fq4ETqK9Y5aZA0TgSkB77wVL0WGQGnbC5zbcviH1DCHp+K7XoZaA4FFExRg+o
WPOfHdrXIGHkf85xoBaeI8kMJE0/qbZnYDSvZbDqI3ojyC4G+HRD+ZOPE75xrglwm+glx0k01+29
PM7uKsE9t00MFdAlb5hMUb6bEoQG2EflQmE/JO0hw+3cj4DHZIghNaqOp9v71mHNMfAjQ7wHOuwf
piK3s7yHItzKgbh/OJQb1jc5klW3kRAUbV/4OV9Kp4NSN+ndmEK1SAnjSUDv/w8kxfsed9xTJUQQ
ut5Hrv/S3jtUfXYziF/f1WuPdjhi2ZqzBn8m3B6b7yhiT1Y2dW4qMScu9GlHr24RWqtODb1lY82V
/uJtO8h7lHfP+lOsFqVUD2uBEIXV3xThkEap5SgfJakZFGKhgEOO33CKkpN2INdU+E7+zW3Dv990
3Y3XqY8BXojjv5lsBH/U5b7RXd+jow35VQ/iXFyIcJ2Ddj1htv5/1qW0iTMWGaNkvdjNW4RbHBi/
94WuMAQjougvyMeIElEe+LfhV0HMRpgMn6vkUDr4TFSNd0Ej5D54Z5bwJz/W/mQQbxCzWZAjmk5K
CXiT3tYSR3kHq7AadS0foK/EhOcfVZTiRk7xp1j4qqzXk0ujL9tho2cV1NFkZlWJXo3h53LKAzJd
Kpp3AfT3zg6GITuOBq9rXxPh9Z1n1ZL8GRu3zf+XdJ1rfR/FSywS5FrO+DAAYXRHcztRlcPhERdy
FVcI+F+RLOPozu9/nDR2eAXijDIvevsUDYPdZzuHMgKfWuq4EeklFL2+chL5q/udhqlPB3Xn6hT6
Ql5s69IEEHUtJiFUQSFMYmWBpdM4MHPB7IR7t5gQqnAehUxLPyCPBbPyk6ePZtcv5OQYpGJbwNMu
b6N9uRlJICrZ5RVGQLV/S5HBHM9IEz8PbJaafK8pTK8tGCfedlkFBslf9+Hl3o6eHHmPFX2DrDWB
3lGuWyTy/VnJhnTPIefxze95FVTE23TzbFRAUW28dI5K1EzS/7Ah0nukhTN/Vb5MkqfP626ikE1s
c2uaGCazUzjuQ8dFzEpXyYoQseq0x7eJBr/JtnQFzj0flQYlWxU7vy97JrJwR8jy9RJUyaEG7kpq
2J1dqk39Qg2zkw7Y0SsHqDbppKeV2hWHmlFpxUDB41quWy/lN9eqN0VJOVtdc9WqPJwrsPE9Lysb
Ap4ebc7OzLYdzamHvcuA1SVFDn7ISW76BJqXEokWDh3kSc08jmO78U8SYLTEAH0HcY8C0qfvOj9r
a2CgUosfCy+GQrOrnFCnebsVf8s2PdbQmvzUNlwFgACmg9iayrR8lupQanxRhsEzRAms/lmL3vam
n4B/lOguOWveJLSPzGJkTDtd5Jx7xHHT0ElGypS7Ea+IHNBvmCE0uZauEvZkTuYd5G/OPEqyG6Rz
+T/Ro3zR9XrMEk0i0Zk4wE48Qe8q/Ub7C1NIsKVsnLzRTFbsQ+IVAk2JBvdF2npLbmdXpBwyunV8
autOSjBnIJKyHbJ04Ny4IZ7YrcL962Lv3ceULfZ38rc88C87akwFUlUMyKEhegHos54PHdqkB2a3
k60UXpgSWp8IhijlQLig3RfuJxhuUpMnUGzJ5R0FT7Ca10MyzMHZaGAyuh7TEPI+Tw2SCEd96aSH
iIJZiZOazPTbgf6/F3zqVCawspB4hY/4s/GOVOB2BzW6CLOGkEKNdoUMcf54smG4QXyEql+YyzD1
K1s4SuxUgs/BV8rO8GSFG6r4K3JNNfkynwTsRqMdrHMzq/nN9Dhrsskia9PZLY1p3wJIZTossdM5
IvgL6d5wGW4yPgRASdE988X/xsSHPKhsLQbR7J4uLMKcRqRaoTuzdSjyBW1sK5EvS+Ewok2b6oF3
2sMMfRaXFtdiAmSR4DN4PwNKkG5sDSBT8RddS5vEJFeUyEovokTmLhVQROJKF2F3S+XjcbuCQHLY
ABOhAe7TYYwFSexvYRtvkYII5NPcN/F21vi++wyiEltRet+J/ilUnkMJGm+O+kqVX6P7UnuFL6we
WbEJPeiS/qjFuqhuMb1Hi6GJG745r+AJjN+NT/5TFpPUHbca36QIYYoQSRPvV2L6ThKxtDaeuF67
5Xj8TXhhgeC5ReQd/JNeL7lticPQ98xEFIsEUxoUA2TtDDZXWORUlqs7elToJ9hXb/U3qYHQz6Sk
IVUSVlgcSpN1ww82oFDTNzoO3G7H48uMLb425tEVsYPEIXbDBjFqrx6kS6BTdqNZW4D3v17T501z
8EeRK48ZtTfxxmamn6z3UGRizNBSUOm1CqjMykmPx9ObYNMWcW/mVYrCDhqNcdcuEhmA336JeqB5
2iLTtCMe3SUl9PZ31i5M/z/GiW6e73XpfTBb/pFrjxHzNmhxeTmzgGHbXjCssFjeW4+cHsV0HT4d
qvt1CYxza3/NpASn8Q5N0WAMzjis/+HEpySAro+Cv6pcrDOto367cB4oe6nBaldLRgcgs9WGzmsF
bZtybqbQjTxwoTnOx6wQWoEJ5Mg7kju4/NnL4V6iW00zlzEBcPudP17baYfWUu+mKopPF/oz48ri
WGGHGOdZMn2Tac6D+IORz0DIm5HrGeoBUEVjOeiTb/xdWB4o9KrO+NJgUeX2U3aAFKuPPGPWQ0C/
SiYxkV9thZN/7qi3tt0K1hR9bbArgUfFb2HJzlBSfMzDhx24DbsznCX9Tf8SWxTJs7Vmz45OGOkS
YCfXfi4e48NurhyN12ajMqRdx+hMCEKOH4bfjFBiJ+Tnq0348TD5TLl5IvTjvdgJmf98fZm74VB0
AZ9OPwy5YXSqvGwEJozy/gNp6xqx2LBrcnFKvF4K3Txnv7PXuPhIY9M6v6qOMtHw+ocj9FcVC1Zp
rXiw4nl0zwxQi3s8AtR3tJ5fegZCXOA4iTA8AWRyQ2/+kk1DEEtzGFZf5cvgI5Pk4pdLeDQfJH6n
s8uCcgu7fq3UjJpmL+z/rYUF8B58Q7DEpFJpF/wiYwqFX3bOK2Q9chSKC4mNUPDTQfjBqElzSmxs
fZlZCwFwcUTI0R+A8N6cIr63dlfgj2X7SAERqyUqrFtsZP7aNGVXh2YMghdYtVuBhdlrurThgeMi
dKtun6cyxGdpAD4SyAOKdF4n2LS3UYSlDcP69fOV3zeJaFIvBdwOZ98bNvedtond8Ym44zIiy/p4
TaHetPNBU7yXuIIniNNNs45bX9AxdAc/FfVRSeGmv6ZnDKMzVKXLggSoPETmQ3VxNz0Fc71q7vvZ
tCtxC1ZTrq+duW6iu2+DO2bdOeeLRHebdFwE+d4y3bWEdM8GhR2W/f9okZ8tvNFu8HRes0302tDx
gOqnN6BXZ9U28Eb8zl9lmclZzMwsPEKuHW8ounoyq+CSx0vhQk/7OLS4iyMmbDlmj2i89W9JiV/p
qvmr0gK0k83mTvgtyo6HBcXfqiLXaSNIUsh/CZJVuvkuMrIH2CzwSGAcmcHvI92IdRUCLZrI/7EX
GF64steiZo9JMfovu+m9c6NH0IgMchj6iP5ExAQ6i/qRQAMczfOC+S1qXhOnX95eatXoCAWChU3x
SHBtZx4Ng3Ljut8v8jWXRTYea0ykF5B9mAG+dzumV4uS8B3/HEvQ9WtHkPcgFu2eS8FgMuycDVPu
6HWX6x0/1oZjaAZtHk7Co5CGk2TAnmXIjUZ4PAJS3fCBBFDSPrv8gNqweZNV3QFKvaPNIFoIBBOE
My4Knx+JOiPseWaixJeWNPQuEnFktFDTdFW6UwbzdTBRjcOu7z5UYulrnHA3C4pWEWQjMsonWm/V
c6oNk8qVkO3R1sDQR/bylbm5tLYY/q/AMXILdXDT+dd59XQpLCXz/h8ujVB4zUJqgV1RRindRTU/
DwCY7fniJfglnb8zmSFKDPLXZWwd9RYzrAIllQ9J4ibh8H3iyUJ0srkT3KcDzewCzP0L+QH7a+9t
tMFbz/GKfo1lSALgdIu/b33vP5vGtVj379II/ZPVZbsrPzsvtH4Nb3kANOdRzmSTqnY9SvVOyp2o
Okp9+Bf44IqwJ74thojQOVVQzyGtugZnDHAsoZxxOUBBQduC5h+QFWjK2lKdDWOWvXe/DKuztkzN
0ahnakLOhtWzEPpNQXLhzxPeXS61GlXxlcY0SdQWBKtAEj/7cSkZ11C2MPuT9y5SDkWrTvcHBIra
LYLjPrhNtA0YERCRHmbjP4Ia8ke5Himw2BcVDs26bv/5VLMcjfXGWjXgabwVStPf3MyOFGaAFg31
1sciJAMGvZYIRFfwCS/9AhdMruHCNbYbw2jvYrva+JUT5msjqIY7cQO3Nj+oY+7bvX5FQ82GVfFZ
uLotIPuZUF/c90PKqguRfxtwhGAfMLMIdaMx5jEeaRQajLZiv/kzA37tiQrC4jq8fdSEVNiGhNjp
xXCyFbhT6WaH5RqZkP49hgkPEVUorLuxv8IXxA+e0bUKWt9xV/uHAdg3h5+89nc+5w4U/mF7pSFT
quvWMgYeLwtR92ABcK+k77W2t17aK1Lvf7zbtSq1Hpy9mCbUcsRhcaPSm46tYzncOvRl+oh6+3Rp
ydOrm9B5J0RVp3uZRxwhpLPOmN6VEiA4hwqu8+gEHkmq0cQ/RXEkopxHhSbv2AeE4R3iKxsjjmyT
oYbET2afo+V01etOv77olo+3wyTb22WZKUIkT2mM9g0dK1nQPEw+z1Jv/tzLVkJda/NrlP1qTb/0
hE8o8sHmEKW6qlqhLmCz8usvZj2YvryFIJl74Kfx8eO0YFgHAMB/R/EcTVUur+2iDvXyZ+CdtPOJ
14Ng3NUfaCnQQBU2FInk71lVyhIfG04AS2AMlc5eq03sCB/cRVUcgD9df0tlpQ8Y7laOpnNygH+6
ixTmh4RX0O9DiGMlBg5iff2OfB7dkHcQbCbb8arYvAPTrR0jTx7NoQgCaWdWygvQB+0Ez8WPSdIz
ghQaFNFju2276ln2yocrPSWki446vZmtMdzT6nrjsWnl2hrCBL8wrvrx7E9WGi2up5oDpY8TPmw9
VhyEIrrNCuDIQfV+NlFInX6PNUijwpgtLNu3H+nJSOWt5wXINoQXxcqQwi8yLoTZDFush1+PAKA5
w+Wxkz+wtU9442l5u28DtOw5V/F1oRo51/H/BLnzpGP9zspKS20sE6bi0ZGJLLzoDXIpmV2RL178
jACzdWjQz1CrAMz4D9xNMMZFjbsVpYleia6jNeOTGhRTRjeXMyqpE6AHQAH/T7/R7zxHC5F7Smw1
fwwJp0H0+RSxJROi+M612KsQ1PWppJx1XX1j4lsawFnNGKI54hknX4aSpZlWZLZ8IBQQitmbmPMx
r9H5jH3Z9XDfAyBp/k6OSrAH/TfP0U2UNESFjY80zdEeR9d2vjYYD3uxO4QZa6PW4o51I6AxLl6V
WpwxkFzNjiln7x0x0k315opLw2Kv7SpfJv3ho1PXdUeNlc1h2cC8IkyhfWDOH/XJ/foKfXNcgPGC
ZqP/ONuOPquNrZYzRmn3Tj6wQR46JDNj/xdqke92/BH/1UIoGcQx9kuVmfKdvMb7+MJs1H2Tw+ID
tWuvWeMVvjZgAjskCny6KQCE1KerY045HIGjv401M6MQ/OrHZmReiP1+4WaJBiyG+bhVOF1uiFUr
cdhNwQMQDzy9ZoBOydH1lZAp1pm38Ghc7dBRHoPU+M+EEfY86wDZ+4X2lWj2TGtoYolPe3WjYlzt
zjj3hDWh4xh86H7hjG6w5peMSyN8/qPvMNH+WJbG5FhDLwJXiXEJHlsyoKrfiGHClNwLC+gZltoP
bllnUfr8UiSK8zjCE3dngwpnQbtxygRcFl3XUkCREngrQyC17j0SaAREJWn2xKYm9O8lrz4FKJQC
lgqXmu5gOnSykw0OCzMz6IZMY+oPQTa0iEJfOpmQrH7jhvtZr6uqXIhRXpzRxeyXfCE+5VqFHakn
PNIbWdTwh04KbIWK/zvwi1R9t3kFjbwjaAgDkJWQDeTwzL/ua3UJVUl7U1qCurwf9c8Xkj3PIBv0
zoUnugbv1x9b8cVjuCHItJGVfdc11pxcoIX/gdyppuuznsqnnhs7ycEPQAJZ17kRdUqo0MVT1lzt
DRoY8+D4ollvtTDZ0ccZtqAB8aLuinRPKWcW0O7Cg3zZCjOR7NClR2QBxkb7EdgDERd9NUd3M35B
kteBv4tQ9eB1xqC7ER9QsLvqt21STuhSs9c+aYLg/yBHFUf0nsbFA9qJVoVmTn5ZMSn4eMhRGENR
b4LqgC450LSwyOarQVaLRZkUiuid3T0rBxBa7oQdKFRTanfhTw1VFV9ii7tCvX9tyb55/aWlhHdE
PJ267Z1GnMZZbc+BZFPLbIzTLJ0yj1Sj/ehnfOYtJfNypv5a1sPnQ4ah9gfVykQCP3dbcP+N4fmU
C8VXYJp8W+eDVcGm0VsrZgcgKiHlccnKfyUkQvcNsfpixsuj7BdhZg/CP4zfeOLcX7QRr4xSL5oj
tO+8/nN1N0U3Bjy7IdQuHAHTsh217oUXTUl9WUECF4RwWdgxFMW78RiEzLjLrvA416jgQeUFgXBd
daPBCgVaRDXA9NV0bqwl0z1PBIi59od9KNWRNES3s0Mvhw4ysElGSdsYgoHIx39/Ggc6KLECg5Rr
iMqrWHIWzgc8BGiksWfBq147/4lnAQCZBZ9t2NWtcYGDvG32DTE2CfQrTrLrSXeiYQrkzUF0EcQh
nF4pfiIs4mlM+Ry4go175ZPwz9jqMZDz/80J0N8LBq7eM+tHNYVyTNMSlHgTG/sT6cvvr73F90Wm
Vtop4L1B83vT2EGsCB5UIEjCrVKHTkQxnBhzCn+GhEVheKT67XATwWkZVO7iVdWM65jgPi9w3xo5
dFxcvaiiVM/3QD/qk1C7GbZqvwRZHVMdQckC/rZE5Ev51unryhBJcZZaIQ5GIwEUj+vpkT0i7PgM
++BUyVYwW+i6MjTo+tGfoZPWUAPIhj/DEjpDlD/xLD7rKMVrxsv/lituk2lxtSgQKK1SYmUzGFnA
dG9+WRyjepvb67VLGZsGao2Zp5XSfPECh9VWr8SLr+g6TtUL2KLl2EVETCOa3wXAWmo7C7YsiOn4
q62QA0SOkMd58NMRf5yBQDqxDnvKadstfmlJj6eJk83zygriFFGQQu6Bek1uKnRw3J/S//B2SsV+
884jpsaH5B6XRdWIn2uMoBzMmpvUZA+qoeJGt4Ko/HlIpTWvDWEm+JSmb6ZIJY0TcwZQqAsFiwvc
JY6nEMhYVItMRvBByWDrAPA0TEoy0wd/+c6pHbJcVlQ8D/JbA+EMYA7AMArGdNpqHamW2rh5rwoV
D1fvMn5OIVS+zyprwTIyqheoLIRRlA5ue4ZDlt+6oSNy2DBzwciTsBUn3qsizDvobQfWlBgSg5RA
iVyG41wQ93IEH88T/FfXNxlLmGWW8EUIKzH5L/NhprxZHnny+MtPkpNEKCn/vl7GCbQNsL6YkN1Q
b2sCbki5dTZVRg/loZ6uMplpPsuvnXBT5V4GEHY70LSU2oRAO46iD512jMynejw+8/EkzPKzhmIR
Zb2NuJcmh6jgReDFc1ZllEo7hForCkYNh62dKJATA4FBmQdE/hXqfqRjtO8T+UmwTDvDPC692A4r
hQF/rFV317m6cBA3b8EGtb1blh799lJl5boppqzZ16xtpx/eFPBAVTrlwPGUee8h5tdkj4VrGo0y
3Np+EbbgolHpA5xQ/5c4dRrB70CB2WU71dTvotZc1bc3YJnl1qxX9eUfu5/XhKvMuM+r1vvhehSi
xy/wSW+w3Wv8U7rwy7JeRn3eg1W25GmK5mZW1rkdusASOA28Aat7UoFFxFys1U1wnYMC/ZRe3Io3
lCbuNpe0OHQQfd6gvHiue1Nl8JMgT4nzrkY7F1M8RQmiE0Kbzf1EU1Ujb8+r7AiW4aZKRmKEYzOn
5227wjmVSPZG0JDxZgHsVJpdotx1dmKqRXAcRPm02kZQVHVWyvRzIjk2IwOQYsxg80khGkaZcBzF
+osBuS8iY5WysgeY50/Phn22ZmxmrqjFybHKzcVpXKRqQpUFDIItuVTq2ZRcR28PJ8GoZRTaRzKZ
zmN0EKy7tLBJf/1nmAziJpcwuHnDVFKQOYWfAzy3ykqqM0U+AtUsT2S2WN4+pfWfkChoemOPmySS
hc/u1/MkL2o7+AM2H8/9xBVRpZcySyshoOMEU7EfVVJ/3BENyHAUvXYjynEjte9b3Xp/L1fqxi12
K2IwteiT9k69L/Xm/UA/K7kYSz0jsz4wJzoMk2N5eK9CS5FpneBCzRqlVCNlFh8+OzjIHX0jm5gf
jgB0Kfo/+jmbla8AzdMiyrah3pZ8OjKojNF/UCmc/vMgYd6p1LivOHvR7W+GChHWveiPVn9MN5eJ
7WsSdFa1weA6cgdtXVhH7q0SCdEbUXkpeWRZ0Ilx6mvs7rTWuigjZws1wYiGF2ESiSFMn3an6IGG
k0EkaTmr3QJesisdFK2y/4C0jgvZYjowvsstbG/Zz8R9STqd76nloeO++mbe0wPGIqju82gOmXEL
W80TIy+P5tJOWiu9uFiYJyTCQCN4fRjtpE4hcLMgeGkjq629j1Yw9IqtBmqDvOQO/fHaW3Cof8FS
xsJ8aTcLqf0uI70aKw+yzekydnFmsz/Tx11m9FUx0c1IhYdt/pwRPo/5huoxQHG6d6nLgFpH3gqx
IvbEPJfaTuVgjRIHF8Vl3YIoFUDkWDeMI+aNTtXltUcEl87rIESOAQxjcLOu9uVgTKK/yxWnddLq
VyKtSk19p6Q/gguHXbRrZoaadmYbiBHyT2G1YQLzs9aK/xsJ+m8YZOqi+xZskk39lncG76rM+C73
5aa+RzM5RPfPscnI2B28qd7HTR7rbhQZni5d8+qhAHnGJYX2coD8H7WPQW1urc83dKVyWX1AlXLY
yuoAbEksylRNiP3DIPeh2JI0KzMMSvHvzreq2M3mgXrns0eYTG0N+rKpLAA9F29w3/wvh0YnzMob
OugcrfdxCh2M3D/VXjMShLmrQnUPuv3NrrRRmAGOnUjFVv/hbZ3CATcHevLnNmHjMJLwg2Lh/uzE
Q2I1JzUpmO99PFOMQFC5J/EtlBxCvt4y/trlcbqn5CQvhrxxiwjOJVmWhUPWeCE7DL6ZkLylvxa7
me9fdFpA2SgtwM0Lk19I9iubqGbvV2gRB+E3RR5jpdH9VzvLeOJbxLF21L9daN2OlUfPMvD85EfK
VFB4c48/JYkV7gub64Touac01WUuTHcnYwH/QV097eGVKlJzELV8b7SMbh4WWWaih7sdAE6Qiw98
ssbVdczD5t3hFZ2lEk9uYylpL22ixdfiahcKCyk941xDcXRdvYQe1pmnUNfg6wzxSLiOWmTukD0B
N5/8HrI4hZHsZq3aOSPCRWhvQnsCUP3lmKIqGWIHHgVcS54X2PLChse8Cfuv1l1BDvO8sQZJ0ZsC
5Dm6ZNeyi5cUhkIVLDTmLwnTBU9e0ckfbl+gcL8yE9k71EQQKRtjhEpVEPJoLkOWo/Mvw+e+Q+yq
6M733Y4/x9ZJwDkwKYDHdz5+X+WSshegWQzFKCcArICJ7yYHc5KQzseKe9AOwc84Jy/iS8Vanpcc
4oW89qN3AYbvftqgXeZoidA6PK2TlZgfLDXpS1prWgQhORQOJ+gCTka5I35GuCxNSca52Wz5xOxa
cL7/vKMFToINhI86p5QmRuFZbKGM4rqlYAixkySGs7E4q5HArKV8TtH2P3npBAfio2nHXz3zNKr7
6WKYguDTC7OsR0FW94zFmW2aUX3HCjzjULk83x0Zn1cA6RdP9/C+37Bv9aRnq5DG0tutpza6IT85
iMEM3J35Vu2TT6G34h+o/fjrfavgleUqsyqTQRziTV7CtX0Ix43Q6VLceq6V2lublqfOQA4RnvTe
txoJjT3zmeVU4jyaBVoYskFjryG8i9O6hxSXDVZXx46QvVLwz/Si/ejUGzpHYNAWZ6e0i71jaWfM
es4Z3uUrs2cgkH/TZhcxaaG+gxeXITDxaQyAfqqlSPN7gFE/8eYc2PWhbUxzRjLwTYaFsuR8+BHI
4wiXx36ovvb9TlDXtiSksUJoQ5ZRDb7qtrqnp36Nnsey2AwxJKUkbBvKIaJCuv6cR4EZP9tQn1Mz
Ww7cYJ/XaN0nurMQN40EzKUjHPunUhKc6RMHrY/uVLCOph47m8pCWoPayDkx9lnknxetWQ3bbEFa
QPtMIRqgvgvAZ9ASdM8Ianfw5OCvPSQmWjxhdg8YACzmpBi7Ewtg1dvPlzJ4L6/5ZWRCEpf78Rm2
6yWTwq1CjFBWbeTgfPzd0pjxd3+FWQ92fbiyA4E+8FlH8LaeH6XnGVJbxv9dgL5aIDn1DHy9uQBm
rOZf78YTpfvTmVHDezE7fVJ1vduilnSVyXf1DD6jKF+PMuqnGlb84LMYxe7QY6amJFkhqG7znGew
izXC37Z6bI5TzgRLUE6Dn8z0mWevdwX6PBq2qaPun7S0w2dGxmkWLqj3qYaZGNCzLOO0dG+tKw+L
qRjrYp3ALNHEeSljaXEeqcSrbYeUrG3ev2KBAlytucrCwRJMxt83Irl+RuBc1At3fO4re1q1oqcZ
876x8NRsXZ+mYrKUBu407I8sdquE/FdQGZuSSybDt3fkuiMPaJAV9X7z++l1VgXC7erj0hc8LZH7
8mN609zWMkzy7x4WEdG+tj/km9/2wSJV6q3OQXs3pNOYRKBKMMO05/4gtlBaA92GJpfWHRP2gMHM
uaoMyqwxMNxSMPE5aguIjSZr40I2d3hUHBG6/CSxEGtmtLFQ5O/AX2pN4zWeqCIC621cwXhizNXh
xJQCBt/hKCaJvFHrKIRJxTamfzO/QjQnfGtO7s/EVpEXmOyldR3DTEpmS+0WAAwFjaC6aFSFS2/l
IjpJnLyv8rVeE2I1khEyvzqA8dFO9+d3zZTThSyAn9iBNHoaHFL1LSKduodOSyH1iFvobTHlpdvS
RUU8xN9Y2PXsCtBBsislvyVySxj8h9DZTRz7MANF4aHjb3oySzaBb2Qgkn6RB6Z6MzVmXxzSpxDt
mMvXiHG3eybGh+xpml8kv8pZIsAlfe0/hrlSwD7xkSZYjeb0Xvq/+syHjiRxuyca1I5CfDHI68Ch
fDH+DIoIvG+d34nACqbLn1ax64ULu7c4Ruk3D5FQ17jmzOYiQ7ccnQ7JCRGFlWWBvXZN1DMQ6QLq
6ufi33mhyFfpGw6Z0ZjN9h4NyJ2ocV+kubJLF4BnJRSwQHd1VV6PzL8woBTOIqjURI4gLF1Y7TWD
l9WrRliRgW/OesgZ7sFZ2qO8KkrcEu8QFj8IRjb+7QyNsVSrJ/SaAAJIrFz2kbQ8Zgzyr0gr31s5
byrjJ8h5YzLNQ3U2Z18gvrYOyikWK+d8367lXn+5VMaIc2QAdOqLHefGHm/3uzdFsTa+2AvloLQk
goAWzRnbMq8TKsstCTD7XTyUE7YZ+r7NEOyGR471va9qGj9QZbycxM4eNij3VylBp2jqc0TFngb0
2QC2pbIsCeRhpF4ikd7OJIJjbQXOtp03E50hzu8ZG8WeZhqr6mzI380rzfQF7dmaSwHbCXrDKtY+
xDJ8ArtqUYm5Yeu3UaltiihoJMxwLQyqAfa6lsXH+R1+1HjG1TB4OWgUffm0jCpedBVgqM6NBIde
fVvJv3/sE4n9lU7FbkKfJ8G+cdKWhqI2KNO/jpZQi0IlsFdTtclKRoZ/fdaIU2vTYpPjWXPVWo+o
TBapo2RTXVNWRaOp3cirdodhJLGGwIAXktDuIVzBjDZSCQqm+png93SDft4uwICva7FEd/z3RorC
1aMfOtUiK/LL4gdxOzcug/sRhRdbG2THln686+UiPVBK1XD1QOiHZyGiLQgfM+oI2vZKmGsR5j1i
Wg36ISNn4uy1gtJUWjl7pgjYIgRoAM5hN8fnxgnpdWB0d36s5fVd0hVJNxNjBNabt0DuIVE9KO/G
cFa3zVfC/DpyVyNetUWYxpGOLTzH/vEZ69CdNcc+Yicn+61fA7tUpVWyvDzEZLBvIeTcAKXw/Kk7
QLb/9kzZBsyv+sW23lGl8pZX8Y4C06kCjwBkrtZ4E5vmCnK4hZ1Dr+PZxiZalTMIkEpmG7seRprj
9nS28ufNaE6qmvx3e+KAzI5KjeTX3+jF3MBVC9bdqD0LKKZACxdrtZ5Uc5BqJFD9T0YFe6yln/GW
GF25A5hM0ucLWmcrZBVYG4OuSpZju0BvtdmzjJEOr+X4OYUawcevE89BM/0Su5GyFiKcwnmfsq27
6uSI5uvUeocXa2umlCt81BGKZ+uLF4IuTezNA5ru2A2rnAlSPHn6uqGbXlz8HxWDdbliGHVFHBmw
9XP3ENOzidQe73c43fzoFaTuJhOCH3JtjcPzAEZNvKf02ilalYvIFKcJdcWCOjm/b7MNT7MXEX/8
cqURtdUviSBDzZHHHovsUCf+SNFC/WR4NfsS8FAdssPr3cyvOo2I3SfqNSr5o1p5dFrdfNnG163n
EPE9OcZfYiDoc94S/kjR6ixnxmL3Ykakrc2i730ktHZHbLEzYL4DW+68C7W8XB/tcONNwYoh89W6
dmDtHOdGwd4Zp4iP20zAwmylzzRCyJI5mCuRsCkd2AnPbL5Pl0Ovow8VmPr6lMdHOB3Vo4Bmfnqi
KQkEMHVWThMiuS/I2f88j9p1fkIrDjdzlJvtossdFuAc/I70R5ccD9DUDG/y0leiCkfssEpKdKvc
nk4xtYu2XfMk1l86UH0wLFN5YezB9BYeWneuI53X6wNIfXc9A1bHetkOVVmUtonoRRff56wgieLV
lneqRFs3/JgVBeoHP/ScVOoRaRpUP6ngRtJjgY8RtdniLd2jjeL3VQrgLCtG3199JdXV54O3z80D
znVyGm1D8SvKAnHolxeW09yWRhhqmIEepwdK+MDLuU5Kedybtf5kqIebWqk7si0I13P2H5zvc5Qx
xmyfxwSkb4Nf0v35jNONqcjY9ZSn4qgyybXj10XvSzY1fD9k9zUiWcw0US2/EOSQykSETa3Ua65q
lhE4NadEn8YJThjW07Kd+79/auZO35j52B3Z4XwoqzYLMrYgPUkAqHsAdeE9+CbgdNgg4pz6Gbci
SZlkdxfPjwNa6L8C+opNpunYO4jG8GFEKvfr8XKxhqUW8oetV0xF47xN73/1E/ZjZHxJKZZYIk0x
vPP4o64nR2D3+yCLYwLY/bCVr+4muOzYWDf8eQ69kqEqRFTVQey5ABuhgEvl3GSfqdaYlD2JrveL
jkVFI0pixcxDoeVkKVtnl7IPKW9fDZZl69MehTSGuftniQ+QwncnSlpLbyzkqN8G8UaleZZFOzVP
QGL6zhu3S9+SVe+sw/Y2UA2uu7m4fO1Yb0k1qLugVLX2NiqCs60oOWK7vJCqVgZY/8tazKWnj4Ds
obG5fFzdx//mDJWPdK0g2OmrgY6R+BVejorsoU99QGs3s3gRaM5dHWVpihXYR5lav8l2TD2B7wRG
nS0d5lXVP/3WXtPXK7x77BEP6aKSD0X0+ymhK8m3anrHZEb/pkmEf6tB2rhW4yyGGaYXiwwTxFo8
VpqRc1WNmpHdt2NbOpOE0gcraVOn800VLgY5UYrV1okjJSFQ8tDhWlQpM8mAUjVELwgMNXicarYW
5iAlf3LEEw6TzyBxAldOTp0V9l6GoBNHVnQ2JlMTfOc+PCsYx7xGpm3QtHhsZwEmj24nurLz2Eif
fUkNp8LAg9OE0GERKpXn7u09XgbImebziOF4yNBBL0LFlfpY5v1DdL+htUgg8QVUyK5RwVmJ5REL
olhym1RSszxQF15vrd+FMXobTLMYRixl+BEWoxNH+2rExYyV2wbRd3S+Dac+VTCJ6HGiqY8RnTJW
bXkpcXOvFXEYlZ8Wu0bedlaZU7UjIyib+pV/OEHLZzyv0mz8B2GPFujMwMVX+63qk15nfZ3ZQjMo
DzcJELrz/s9hfRrlmdKAF3E9VXJb2Gzg+EU46JD8EHCUS9YzlMh7n9cOjQ2ob4486SU30/zmvRA1
/SoDnZgT2ZB/yCQ163ZU1+VAzayAeoB0ZHQg4C6dExFhbo+P9++EAlKZq/ULQua7KO7UI3xbXJiB
MvIZIB+2eolu1f5O+VMj0+mxVwY92Mi8Zb2AdrYXw9xbjaMLbl0kSEaIyo7Cih6BbR6NoDuSCuzc
c295oN+FlwsQjOafFUhuDl8pbRApiqmqoYN99s8ThnZhNRY953/031xnVSschaZFY7Yb5WG3ouZZ
Pwq9oW1FjRlVNwtTKkYz4xY/8sxkUHLbh8JES8eHRi98te0da6Eq9UEUykTuLEYAnkxsHO67DEsv
Tl/MUZ/UdBzBcIzFDqofR6O7ka8ZqfTI8y5+GZJXM+RsQn9/3+fQWx6t5Kh7ti1tNbA65J+p3BoR
k71uEjHtBJ6y5G+y8uPO8Q2zMIx1L2b08y+bTY+YD4mpjr52zYDW3BhDl5aitfKeOUSI/Yqq2s0d
76rpaBSmAXcXsD94WJKXc87rD5faX8lK1Cjjhy5LgyUWHrCAJ4E69RyqQQXu41WyOBK2Df/ynuAZ
s3GLQfAnxy++/UutQxqJVZangN6oRUWrUaCJGPYOZHrZZp6HOyT9vTcAQO2LTliHYupehM+Xi8rT
FLJow8Rx+p6HjH63o8wk4pJ9plmTtTWdTx55zOK469+0y+JyPqmWJyx5GGVTuhzv6qMK/VbCYAr1
3hZbgOZ5akeIUk+akaOU3w4qMcPQDabomr1R3w+4shtki8pBw+NkWmUA5pW/oKns3AHqv8BLVbYK
wyMCrFIE1i5QvbcDN4ZDRfL9VFokAdyXNaMvQikLD+A9OHxwjCMhHqKwvwPWjg2lxFYaHC+yEiu8
ocdIgmZZoy2Q8fyeUB5OcpkmhOmfgRPpMW5M3rc/HnTdapMvCHjIdvzU3zKJbsmMoinkGmlBTn0S
cLKEFKIopVmvZ4oFXUuvuwLqQ3J1IreNLeT3oUx0RxPc6/wsf/sG+cHTO41bxMix9uhpG2oyrqRt
qgoUX6EFYH4P9Ar+0LWiJOPPRPUoTXQV3IlvFtr1LWPpbQ49c5EMmGmzizKIAkmYs0KcgwyMmlJx
4GsGr0d5Ec8G9jo/XkVIDUwB4fN7fTzgJjhDdRwrcbMoWikTGuPiNw7Rgz0i9pOEZVOeSYGGv8VE
ko03ay/3Lip/SyrXtC4fAgkrexl0CRpOztE31+LUIZAUafEwnAOBrjLumlsQrrOXCG8LtNYolPKG
oE/af1nM+XFCNIkN4IuP9Uo3J8Wn5EwSKkqhLjN3UhsYozkbJYLrylDY0YFASckNXGhszOZrcIlM
/+mDLYUbqRpAi4/bpqVkKo3btRSZZ0jpmwnqMNrtPBebLQN81hoqhzdd5UPHSGTVmA86CjR41l8+
QT0TNvQUHYblJ1oyDHobP9WDJgA/q196RFb7nFnMok+WA1sWSCUiDy3psacAF04kHlQv/hMVucT9
t5LL/aGFTakTYR+NJecZD3yu+S2WXYzoO5sytUd+0NmAcxJdCANFKjN3KEaFOHGimFJSQibBL1FC
m3gRfVeB7rTcvGhRSDBKhogZxcAzlS9Owx/fL9DQUIQ0NNuFfiq8U70Dvx/omeB4J+kg4jJlpGyL
oC4Xshrc4+6KE18spWu0GSCbPiQT3QfevGlQ14v+x1AuENjKHxDMIt2Dr2NBeus692qodjAwUyg9
Ri3oWcsUWku4H10e7GMmQ1BdaODUnxn4aPQqeh4EibI1J5ujPtxOYjtQt1QPBMUfk2xmGhRJADao
TBXHWqEoNYPRJLUjABIxBFNXK7aSyPUh4/JH9fTjLGS0Ck7Sgaqq1vrYHnQhnfxoMeEoJXa0nneB
WvsAp2pG+omqSQomPX0NBL3WOy7wGrBxFPTJBHOy3+0OlNpQFRPR0aW5nKsCki4mmnNfekxcvj4P
Uflt/IlMjSsdYMKVmI+YHfpgBepQprngBOHrrBddz8Scn5z6SMqf2WQMcwFbNV6vmavGbYWg5eAp
RB972ZMLOB//v1UYIxlkFp/AZS5gayFFKF+9C0Wn43bljl/CUohx3a1r3QScJlTWTDe720fc0Ghv
wfFHB6dq+KypFgzTnjuyVCCo8fXUY8p5IOLg5fMQAuidzSN+P8hx4xIkZEKSWoItyzUzZSy6an4s
JsBjvVRNh5vnoSBP3i8jcQoB3jXZHT2z1nzcWMrus/XcYmcGf8XLMn7RiOS04wFZM7bco7h4SkHw
i5juUBVphZehpOsRucIzwEZcdIkOrtpTUOdcY8TmMKJ8ye+/DrDd+lNl+DK/Pqm0Vaozvr74KSf9
FSf/RH4kOLkqBI6BwzjoWDihTITLrFmIE+/yhogBbZYaAzrv1vXXlNGabOTtt8KARaZdPRitKRuv
M/1CM3t70vjEZQk/PlIRgkb05wEULoJa4dfuJSNqpVji4Kud7ZMChMkpCpCAT5cm4mFiOtSgN6Lp
zsX4bPJlha1HPhe4dSLDAJf2f4UiSpeLoLU/C2lMEJLiSyAGO6gQlbcyBd/gSYIpQn8l+6YyKpO3
T9X2c7sS614S0yK1780SkIRB8ZyNHBmQv6yRVX0xOjJCNkPS9YF9thJkIZdFNWqK2dYUFi5ZeVW3
s5bOlsQIm+1blwDXQu908czoTt8U9QAqPvn0TksPPfX5lbLbptQdXoLOSt0jfaG1RUPxa8NjHzv6
1/sPxuyxkJDpEwSHIB6mIzz7svsCjKJiNcoF+8vPaBBd+tXC+orm/Y3XyZLJgDSkn2+Y35Ssw6yJ
o4XjFZY5K98f/rfj/1g+m9hFX9oqop3yQj8WU+pVGuI9VAdti7bAuh9IZk9I+MyZ5DNikiUmXGuy
YSU/CJDOtr3CEFjpniQ9V2C7+qo6D6Y06rZMpWXANubOJ/T6pPXps8wefdcBoijK/rHQNiJi4yr+
gieYRvVCht0C4K51Aa+fYWkX4gg625DB1o1cN1UVA7PeAKdawREq4HWvPe7VDkv3omMAoE0GYSxR
+UVMAnjm5DK7Al0Ia78j6WF5ram9KbQXtYdAB+R4bUJwVK5dreUqiZo6rjex4y85fpf8LVkKEys4
1a5xmhWV8gAzGxSIVyCP/uAj6bv87K952gjQvSkMh4UBF3B1y124+5R7R1JC9RRVS/CdljivrwtU
8JIpvWuQHn22Rw/4k2ZAInNy4COe9RrOS//rnLTJFjnpF6GrcFaj48VDhAN4PrDDn0wVCQif9EC5
eslLWJXzTsooZDYsgd26sXe1R/ycC4X2esiVD0r4+7PrUpDVMrCNUV54VXJ/VrlMt4fcfcUHwrqw
CXR3Dol1LeIwX/HsMXRO2UkiR4Bnq6I3sJdCTFkCH3TrsbzgmDYMrNub0AZlTGgP6NY75ND/YJ9H
i2tZabrx05TKclu0mOLQqOn4eleUdAVmzAviKsQ5dEhktv7ldYyscwmqaZAhzkaZ0ZOrxqspUCPR
k6mDPaADIGEtR8mHx6EZ6mvAUW22bkQ7L4WSp+5OFO0TfmKT5kZudVhOjj5173Q73+/hktFf+SvV
gZwAPm8HWgi6xI6IOe3sHlFSEyP6tby2KCU3NC/AGSFC+wYr4AOUdv3wZWA0SXss1HJVNbRT/4up
CgVw9BtZrBprdPOkaUmyfBmuEYhjXAeEbI8Cu5QQsjydJ9qVBNEUcEFVSkz2zcknPBUbR1mvGOFM
a1YOc7i16dIm/DSZttp+ie6M2o4ZEHsYxCR0iETwqCLIlj3iTvR3WDNEpQhhQJAuhccdUPKLDKuA
4sfotOgzIwf/h0rtyx/TqwWYMDZufkD76vV9HrqRT6yaQP2kk+3Ukzwb5CKhuGluRALO+YHTdN1d
G0eFyZQHQbiHjnyHZkj36aPJzt8mhcAPNUb31Eh0A7wvCdRQkfDyC1fVlVLV7d7/zW4avNBzCmNP
4qlWhTQX5w95rXjcKpaWAGXwD8JbgZnXjfUvmcMNwcz3uCnTnf93bKT5+XMy7pTi7EPPGNLYRJ9r
dd9BAc9vv5XDqt73J7Qi5lsuwlW6xBqz98Iphchp4CRioDb3kExzR64g3YOKc5IEuXtH3MtVQErg
rQZtnN8IKya0m/8koYYS+De9MrTXEBDvgibHjSWR44kPo1FRDmh0o1l/rdLM0zRC2IpzFSRaLc3A
dLkaeJiyDj2pLQ+O0tf9HdsEUTTFHVxvVJDVTiapHBR57iiRj45rh07uG25Pbopr6erGH9Tyhhrv
M2yUzmIMWeIJDVMeCI+nRDIHI/r7n1n+WkiBB5IYOAN6jr1qeijaZnau7URCWSVvlFAwcj9HE3mO
yNvNc1MU2U+ci6MPvLCJ+qYD5ptwCxzwCS3ivUbSawA50bzx1riGiIgH9viU1jMdnOmyUcJz6sTg
X1Yd6I3la0GpLC7XlbJLInSA80/O2hYMEnKpyDIdA1qkdXsGUbekh+gs2hXMgMY44Os7qpB6YO6Z
PHYfQBhct9GVrAYWpf8yqV1/gFgIjkETzfqzWdQxQixnAfU55wO5+RyqEOr0hajxuOVHd0WWsfE4
Y7qIrVNoPJOjSimNWydOT5ILg2i0xd8WfGBmp7ZAkgqdrgAsEUmrWwHVBdMEnJC2ldcHgTAFCEGH
OHXz2M2R65q9dZaWim+B2PxLLtfAwkYgkgnok1hnlv+sYvL86xJmkOcxM+GMhH9mgnWqD2RpJxVX
1OQqZzhawU9rKxLtturh6CijBkCrpwH+JvvGU4N7g01LitqvA/80ViL6FIpgUE4iOLvpEeTZAdwH
eWGI6LXK9nzO/cIDlbJcyTkfid2HgLVYo/eDJtlR5Peofv8jwjk1656xZQ9zBcD3tmI424t9R3jk
2Wycxd0wgdFv5Hk9gHuWetGCmzSifX0dacylHe+z937zz5rN0PWhXTBYVWHgcyjH+0EhvcPBP1Rb
ctLhndTR0Ylv3xqs2v7VpuQYVOGgI/OLAFEX6MMJIHAniUjeAb89+d8yZy/0meSmCE0yqC5K6XC/
eVuzLAG41aJFp3382bnlN60erizDx6e1VhKf+/w9DF0ZKQgfaXOnTjz13KIsxtPZ4HCGcNidYWEj
OCb6n1RFw8mSThuQPjY3WvCfRkC7fe60dsyhGUhlJRLV19UtJKkpNBbze4Qq63w0zdElFRp1Uf9H
Urg1Aa3DB0eTRDuKG3wMPJCfah6h3qsriLXf7D0RNblIVg6AvLtWRRQi+k53LWg9SuqOzKUhITRo
05R3Ils2U+28Dj7WHgjaYBIoVo6Cn092BF6x2vIoFlJxTGriQFHOQ1Oe5ab1j1LMzsRiM8kYfz2z
dQs9yGiHsxECAvbDybeBP76YkFvCOyyXjCnSFgPrnCgmOR/AoFbCpN/fYEnrMqbjuYj4n3slZ6CP
qdDzRFTfqnv1ejj/YO7UAuq+m0IJG3IsWMnV17p+wqruyBi4WH7D8XGX6VYJ6gwCZsO0HTo+PKzI
QtT8+0ftXuODreENsm5d/ryG46BeYRVQjhL0rr72Ar3i1hYtjvXspvJ+IbkDj96ITPhr5Z705hv8
DOHkm0SYtRzh2Lz5QCFD0Sahm0DwG80Beesyzw45+Bz5TAJ6AEulzKq4SsJDCVkhwJi7MpnsyIPe
uUE0wk3ZrENZt8rU2H4CetVdLEjPxKi154PL2ypgMWsW+3MZBKC39MKBuqYj6XYF3gKRCgIHtHi9
oH/pI+Y8l2xPfiNvKnaxk/6ncTMe5XNy6VtnZNuOLJEsPnhA+PANuaIsxyNYGoBOveQ25lnwns5q
n+pjP7TxtRfc31/5etuOGuHnLB6ZDJHgRwstjkL6dRZg3hfRdc8rbyUO+BdIRovVIlEczQClFGJ/
6M4dA5BxSs7y4EAMT/yCYxk4VRVUW+7GL+LCF92GLJ8/LojDdMDYNkeJeFOycJL8oh2rgJioRSlr
Bt75U5XN/ZVikXuw+Sju5QrlISah/BeqdC55P+dAl4BymFBhYoRPvh5714kZnceQxVe8YRaomGbj
E/gkh8Ird9rzezeybNCVPfQVkRwjhm6vSmYXSCBqDP8+SB7EqBrxcnxQvM56b1EP+CB7ejplS1QQ
tpb2w7Gzw5dwI4sSGkDYzdxvW91jtStTEzHd9KgnjXau+HsAd1SApnxMyqe/aeau8+NQS3uAVPEw
FjDyOhB4fIe82/D+Ia35TKnDpXkt2rVHCy32PQrgx3aX2iEZvQKBeDLRqVEhjdjHoj9hlfzTctzR
dx7sFqhxG/GGCioRE+1Q+Xgn9JWy+33LdnNZU5Pz+I+0hSiCXp4wj8ARKe5vIHKsoNRdKe0n30r8
tQqZRFiUnyG2/BFfrR8GG2qTXzTTWMXKgXYPNwtcQ2rDBupF8br1qUeaa32e6sn0PMaZRDQwS/OE
ZbGfVMxOmnAVy6YVzt0W6ZxXL1RZknO9IRBpBFvOs7T0e+CrOdKg6NrM+q7fdEhZ7KrT3XyEqwZa
ZvYukc8G5pS1H9YLdKs+h9vI5bv36mvWYLZ4fWu4/G788gabGQD1K2K7gnoDfH1IbZlS1XqSCnO+
Kzn+3TEsZeeNzAR8vEYmKq83cj7kJ79SZjWIha7lx+k/ala1+hrsyugnOPS58GDx0H764ou8go7w
Ilaf1Nk5d5TGIaLs9s6et2yTVpU3isNh8zfYhg7YI6liip539YaeLQ5NENPEDF+IdbyTu5EJ7y6i
X+UlqJeE68TLZ0TyxzC/eFo5iCXFiP80vrghu9F6RkL9S8mSWjF0Jvsuq7kQ6ZVse+xqrD6ovxuW
YZ3NbrmRN6Jy2eSzYBAra8GKpQALPgL7KK6CVvy3DYm7HN5z2k7WOvUOqYaG1ZevfGavkABbkse5
hJx1oYOUWhZhkA13JjCqVGsD04SI+M9ZbhX8TNwJtM/wJ5Do4T7a2Lp4u4E80PKHo+zJ2OJg9Rlw
muc/47oVRtYTSeh5ScDtkTIrqGbn2RtTGWgqkGJq/aM2f4q7OpMrPQ5WaXzkNgySc0yl6GVJmfwe
/gLJNGm1IEDMMz4ggq9alN2vRGIzC/9GBoMOrESIM3y1NuTKBOoP0WSAhRgVzX4J+z5euF88UFyo
qrepXuC3jIb8z9sWyKg3DW8r/RCnAxXyr1BCIBzHjl5bPSkNIn0YNO62La4dkxa2HUvG8ZeOHYjN
QN0Gsx9uuyS4PUZmBouuzaI9qy5E9GzWBrh4EJ9424Wsy57UDa5q78REq2ZPUHC4j2BB4HWZa891
IaUjW092vdbiN3fC+8wOB60UT2LKDuAYFRjbt0zoyR+P5hRjNf2/Hz3VR6OZNHMl5rQtxPTFcGE5
0MKWg56PVvCs3b2q80+cIHNmUmlNRlStdJRSxkIU0j+vuA5fcBN5QoVqsEVFznlyDxZ3bDyp1B1B
lTpJQlab7iuZf7tGY0JhAYFmwnWB9Y028AyleOo3mbe8asqbj/gRn1+Gzclqyx6WhTCsVplBg9Mj
sMAXyO2ztsjzdbGNwF15Tpo1v/sQHtTRhHiXMVBjWDedYytwT5xWtSY5yvLJGgKkk5OtvW4Ijf4m
dfRL3wIChcwOH09PLRZxh9qlgCOzdXCCZI9nlhtQj2FG1QMZBF6IkJB3TeZ7I8XdmaiIXGJ1VCL/
iEaC+y8DFRHbpk/pHXTbcc+04rAptxDbyQHF7/g+ovqBwucE31NR0/3oC/fow5yn30f/FhjKK4wd
GXi5ojWHaC/pRFpVkTDMsPzIQNfXIfM5GnetsavKEON7dRBxSo8Qeo4aS2v4L8BTW+uZRM85yB7J
q0JGGMy2M1jOBSTk5rsuJIZZqe2f1a/juOYi6itP0MeR1KE3ciIIznx+l4+4N9r5L3T17oL05bKB
pBh9YQjoN7nntUobEZon02Ub8DC8CrwRII22p3lMGwouI3jPrLnN+nASp/0TAGCkewAT8F8vhXIy
r40azXZ25pSIjIdOzf3NXltMjyNCzgVss6HGd0GycM7XmnfUgvB+8dHpDuQ+zPEinyNr6Tzj0DND
/qlahdEluoiuM8KEF1urA/TG6ZklhQhNcPptB5REH4LltmrnQD5rCrNFVVs2K3NLJGwt06vqrtdU
vMpwYBO10VbuL6YVlwotgN0Sz3p2XRA6z1t0kowBhdqn1vYzBho0/7/uHDbRyw/WbiDkiRRucGKW
T3/83H0J1B9KFDOAQ5+jsklbKO0hFtgU0rtyH8UBIvRcQgAPkGknxgfWvBXFZjlhjEfjEMOdrRx1
5SpFiXUzQIuavjtghm/SKZRnl8UApuFk0GxVVqisBVnw3qWXWmzf/mGskyadeXqNjiynDKa2JxDK
KefM62vp3qtPOZoj4QdXoSWweOS6yR0Dc6A5gcm2yi7BbZOFleJgufGOop5uyB2iEyCQRRgkmMtx
6i98iIpCmADT0ESEMgRMjcckDxBO1AmTODIMH3PNTt4VU48J22ktZbOGYv1NPAR5jg5FkNopWh8y
WIJzd9rWkmKCeCaAPrRGxjqTI/fJ5Acbgbd2uGmIq/QTw83ohuYolrpsS8NLzfE1Y8yOnaxXzAEf
pkDdKr9ephY65vKFd0rpK9PI23HAaABBm9rJym6V0+znHFqSTLXekGL7tb+0a9pmv2VWtuJcYFBT
b+fYH50wbhm24WEA9REwSmuvPDsw3oRXNfyy31qUDrgGt6oLCSOKi18fDfXUH5aYQ5QikJqF91Ep
5lfAAmXe2DO2rAahVxDPDGTxjKgKK0XOot1WNlpHLb/Z7AuDkPuxmXYDnNDAxzRARVW4LjtcLWqk
Dx7PEBGbyWFIUwPPc4n6MF2sVwEBkLfujxcsBwcBAF6Vj1TCYC6+LYq3H66ffQgJPkvkHkYd/1Lr
SeqtpfDEFrFZQwsuUZs60O07T7NChc45vpJyP3QO891BZvQHzcRAGslcljao0SH6tTRQ2/uVx6nB
3ssT+rYtcE3qLSKAfLUYr8NSjy4kp03qdvpEjWHyu+hh+kL40WoODXS8Sc6/AvQj5BeeXZ4JE0pt
zSo4KC/3rzzKVEQDRizLfCKDRdjrPD6KvrLfYDqybQPAuOUucULjPFnPWvfva/7eM4hDDT+rHlNM
CKqs8FAatPXjf2jVIs8YU5/exp2xaf0EEQprXG2oaP2QijuPWdcyZdCx12/L+zHZY70qHebT0DK5
2ED/UqYeFNzc2JKZ7YoA7mnCb0CZszrN3ovGJIpzitwfiw/mfWmWa/sOeA8FdQzEjfmigQrq5GZa
iJ7HxYhO+/cv39Z0Yzw/jDo3AqyjW1HWJ5NsERzE43UwZhAXa4/8vJfmMtvmreKSFUwZhTi50/5x
5H8OsPxPMmfQf64FdsujceE7k+GwDZzvJ0vZ94VHB9/RyYy1hRW3Rb3bV+juxCHaY7W+nQbOB1cm
7Dii/5ylpOdyF8LINanUy+skFxrAJc2ZvDZymOfb1q2fggfqmj9TVqXYBKbUPKtnryvtVRPbKhdt
4msN3g/tVW/90AOW5K+voZldRndZ/dsPSBb/SZ6py52gsGAp8nhWxlyjE0v7aLvtQL9jMSp6p7AF
uAAADIPqDlM9CbNKeoZ8hX1Eyuvq0FXyn25dT5liUKjIxb/vpgEbZZGMv1v0477hNS4H8KK5zXi0
TCGjwFvodNcGPEUKf8+SMs7DlyGaU+w2a2FAhFpKj/fQqkZiBw3mxC2w/Mak7AoyDigC8vE9N4BR
JLqZF3xLoM3HKrne6t8fDdttwNVNU7BY2N72rulTbaBKCoOQHtP6PecBdq2RKeLJLqy90yyeuDUH
pVQrCWZOcaeAgEfktMHq4fAdqSVNuNYO5XMZh0IHO7VmiLky3b2qpiazcNqX70ba4xAcCO4BTye6
qddcHyf7mNNDCPwrpCum757VDr36Ne83xzVSW9MWIIoSumsqYi19WAsflL4i6+o7gSpuOcyw8kHp
apzsaralZsdEWqgXzjhFhm7gOxa2VsUgShu5v3kjnpgNqoVatl0Vfgt/Db8Kz/jbWZRHRnacYqf4
D73lw7Y2okXa0ndG3vFc0KhFm9gmq8HG8SuVTYBIWLD0iPqdiQm/CSmVGLC/E8TQPBAzDMpnDg4x
56gtoV43Vr3tESdqlcK9UWz8+lvzny4d2wsmt0WZOAjBBTtLJhqDm0RH/a8EDbgNfCnLMRelTlBW
mBRSczP30pqmYBFwPPM0RzyEc/CkCGWnFxN9yBfok/mejWg9rohGDjT39BWu67UR5xokIM+8bFiE
BIUQepAbVoH84JGGm1y4ocjhbI7x6wBOfdV0u9x3vtjB3xNo8zfjZ1DiFot1vpdvZuDNjG1MSBLd
wYhTO2xqmPCJuyCeV8XTSuYKOEetcABVkDsZdMKTVjh7lNy4ZtzStg0940WF4y11qaIlBLpKH8Ha
QMx0frwKQbapbCASdl7bMeBjlWrZjhRWON1BnJ/lk2TcOWpQy9SqgborSdUNqdEVaPxxRKxnQbxY
356AIKlS5FhxqY0zSrmiUTU0uEkJbaXVapUU9hV0tBuEmVw0NImDUMbcYEaliFin22eJCBsIkCdw
xUSbH5mblTeqvMR2mV6aHrfmW00Op5sW7taKS98ifUi4DV5g7sC3iBqWz7fW5NX/qyehcJ69w/2d
iTSLDnA6xtqKB9NK27L8V5maj5ER+yQTK7OV3pNq1VC7EaZum2q6Ou3NVLOTLXAN9kU27uQNJg9N
y8EDxQQI0Xg2Yy5xX5b2F6+T+J16lzRWI601xM4XpLfnj06agiogWplaKKx9mHhhyzHz9jwFN3jS
D2JLsRi/l2nULIhJIjclfupUSgbpgVOB5qPie8dXfMNEhq8uZ7TPA6FpQil6DasTVqcLZMa5gQSJ
Q/db9U4mLKOEiZQtsaNn4BCixXvvvifkbqCaxUv2WHDyTNGx2bN/G8UlOaWqnxURQaLjVyQYrMYy
AwRihmHf9MkGyzWFoiZkNwgfQWuPprmbIxfBoXkvc5Pj5K9hjYOXxiqvn5QNrXeaLH+9WrQ04zTs
6Di0uai6iwLFR4oqMuVVSrZMNKBIh0+mVYXYxBz1IfQMzg5MiKbIoWO7xBWNKhSmNIxbEBfPDuSR
6nhTMb4gI/TcjiesJiZQUjACYlQ9W8EUIhSvd84iLAqp2ThHYqsOjduedK9xeAl/EYOLuw0ITOhP
GsO+Ifnv2Ov9yNkKX5LLR+p/riW2ltWnpDF8DnDO8r1wDjCR9ucyF3Y6uaMuuLKB0YsKjW4kaY48
MQ2VRsv4nNG6V4kgaOEpUKRMNqsmqg+rMTVhhlhiBCGdG2GE3o3HAfR82nru5UWigbD2HCrnz34P
VxKPpuhCI2kuvAHJgH36CuoyJLDwzIxyyLqYCKQ+xu5cHJPlZ70bdGfAMJRCIzmyoiuj+4IGrHyd
LbRBNztPwIOqyBbDxe1Ph4tDd0LUZZrCN4ZEMpxPndzvcOwsOo5Ty+51Ga8KkS+LhaU2nZhPQsLb
oKd18mRa0Wsd32VELuOQXSAUArUpP7zBuLnfdGeful4yvrO1k3Jxj4T/lJoOowK0ApmHwa1JoJy2
YVRZxXQoob1MSjU3A/9ral/s/pSvRPTFynWnDqfoAtBGqAp1QIjYTfO4ZaEwaKpSLHz3QJhkzbVf
JlsyW1CUu2jMu/8SgnAvKYNOpIuhwnu0AMqzF2ngqxctDRbi5dRQVc+n3ZjdT8TR/tuyzztiT4N4
x7IU1nzn/SchbGOFSKdkEnHB7ZHnDy5hn8NaUamp9iamBwH6kX+fNOXqQVTUDcrjRBPa7gsOLbr9
yZaWEpFbcPmyChxH+k7FGPHrY2ArqmnbrYNMUpjIVAvlfdsZVzUv6vfU+L79mTR52LFr+UIrcwA6
62Os33OIMLoiYeyt5tkyBsGmyi+cavnAyn7ItaJ6Mp+ggLxB+g3PxuHNZXX+ooy+1VsVPPDJ6gao
9XHb30woirFrlJeZw3RdXTd2HK94R7arkEguwkIvB5AOlt6thNkhLMUoKcHqapUc/wCLAaTE7y2d
aHa4c2CycS0L+KGK3EkU4OdCLjPSOhGLt1C44qj5yG99rHByENiQ/Hc4EuWKomo6QLQoHPt3WtDq
HcnGzho3uihbGmx3yHJLHzgSNqDVoZn4jfG+rnstGUg+jFmRwq/95tye8RoCvvSxY7XI1sICMErN
7HGv+PBefoQLyn0mfsz6msebkGDnbEiZbbrW1bia8+d/fG2EEr10mHSsnbhgvD7aYL7upXMdj2Tl
NDLAFgQ8Nn9KAnRV6UHV4Wh8TlSI9NUcVvVsSfo98GsojUbBrAMqwlhk+DIMoaXF+fkWe3T3Adzr
97gIV11hRW7lWBS7+SeNDcPBeiaTj7UK7GxghgLZXlw7UTjAw/UYZHOKZYdhwMgNFt67GcuoipOI
G7U3TVJSefhGbAqCudPGGv76F/xbrajv3tzsM4U+IoXEwVs/gVQUs6Ztxg8IQOi/UxzDbqbg4Vch
ANJUlNpZu9zOJ28OxHSISDu+n8wJ5mRgWjnlTHMCuzVg5mB3YoyLiifY4qlJ0tz5rm5bsaBisFq8
ahLtkVel3X8lIimeDyWAAzoeqUQh1C0P4VjeYdAg67qVHPW1sAfHZZ529rOp1tABxOnAPpBkaH0/
paB5C7hgA5Pa9cKvtlNPNLPB2pKhCrCFRQ3FswR3/n9IuAkzfpIKZiJ/1FA1xvtxdcjjxKvuW7kM
Uj17vG6YkWydJm5JLNztt0Uyv74pTw+O3qPl1r/kYUPCCA64/WubjvBYoL8cKokz3iPhRwN0Tld/
pPI6cLrW6/KRXbfwSCA3dem0JPJb+Xr4wNqJdGZHgV9oJxGyKr2vJwWgY7ZhDNTHBcsGMxfXyLum
qD9ZldWLscCbyDZKrM4kFnOD2FdHlLAWD+Rh0hQUoGyxL8Mdj/sqrEitI+NxVyjWYUXUenPVHan3
yhl7fI67fUlSOR0rjjWjw9AW02oLDk81RRXYFUgC0Lbocwnwkt8n5p354Y+db87lBO62p6BK+xc+
j3Yhqw+HG/fBQ2MI31qS0gqzHX9DOFbGGRudI72CV0jejHmxxrDqS/aL21GPlUo+j9fk+rYJk8K7
I4OdXvxCWfqtvQ1Svjw5cIgOvGnAn6LBIhqAdJ/nAGjp/mVKdqRYKYZ2nojOQQ7jDpCzDhtnguwA
XZEydh89TRoxslKXNUxCBgMgE2QykdsQZeYqASW503JTFd+kBXEk8Pe7nb5i8W/0lrvVq4PspwhE
blKOQ2F6VriHiWmacgE9LNLpTU/uPmZQ1fLIiF1BPuSd16BKn5nugwLUdNh7gC7cgLIiNr3cNx+w
OP12c228yRhPABnjjVcKSM7HfKTiLVX/oIoXaYwvmH7Lmrj8FuL9JILcKkr49KBhOKG14e+PD9CG
cP689nc5WhQQsYV+ERkrdzFaH2aZDlNwygErWJrEaiDURoVX85cEWEbIMLpZgNUMqwvE0N2g4as6
GL6MI48tkgd1Jy61APOaotwZVUfzbW8CD5Z9HbWq45SRV2IWihwVUrown6h5Bsf5AkvSLnrbcwz0
FY1XGevGhCdmyOjwcha6s++FDJB5Bpz95V5tuSCcjNGlnlhFix3e2YtmWrQO4qLeYIpbJ+H71tnK
DAjWBUrHoraveXwhYYNSBotuIdupOPRJSl3BxfbBNH3eLIz6KUFI+HyBwSLfK6i90S9U3nVyZRgy
ut5XHIMJ2/WKgO/mCTtXnrN+gR54dD+7qlSHJWTmEkZenJygq9IYcEOrHlFO8RIhc8ZlBJldRKaf
8zNXQrIXsor0o97Lr7REr3ajiSxdwDXYAjdybeenYI+BD5Co09vgOapa9iF9o28z+3dgYn95ISmL
6zUMBnqees6sT4Adg9WpqFD+mGjwzzDWxAsPw3znsgGnCnj8ES8JYyLejgVILj2Q2N3+5VBLiz/Q
EmxqHvDj/eh4JgvVoACx/NrmVU7vmr5YpxWW+ZsnLAL9HPOrRSRGKJ1PouvdWOwcg4TfnIG6gga5
ZA+twMp9DyxpUdaPTKAKwBu/DaTS+6nkamWoLSMD2i+Ah+t/NX3ValCnWpciq9E9JGptjtIRKuDi
HkaXjZr+/0zybUpApADzzWzFjM6baxGubn5J8LWI1FuFQPYfuB+hDw/xIOhkhbvjMXG8qyiZG77r
Y9FjCQEDdGUAiAKmM0sQKUscbE3NBLKsEJTmrARfkwz/L4BC1XaCo5C94edqnsLV0+jY/K9pvMWt
f4T4XCIDLFmoR1WKzfpdgrVM2CQf6QrSgKYF5KSw4fL/WCNrjC5G1DDg1M/+WI4gF7+zve7VTW3x
6MSZkXAMKP3o9vh4LsmLWGA6qry/j1bqHfx1J6b1HzMKQ2/62r+aOmUzf5h//dlkSQuPGox+rIDb
TaPARXUBneToX+vqA4sxNlG7lmC51W/mW/79GVe2f+M+THEufjUQF3y/J/TROj+g9naLxpbOMdeo
dgCsdOa4P8D9egfPLDo1YiSmZGBEpTUymLgo9plyyypz5tQhoPr1TPELTeB/pafBs/lViErnAKom
Gj4aAcWq9ZG+bmqp7jUK6PNPSQ+fEH8w92iI+sfhQ+5ZGRgIjHoaZ2u6s2kNyeswu7CZhC4d1AQi
EBT25k/Cu3QJ40ldEgUsamT47DI+PsBxwQcAs31b3hy2bZ1PXWNYqGQippwestJdc62nfoydKHzq
Psrefsn0i5Eaq6z+k84dbBOEWJh1g1qriUlGty0vkbGBK0MqftvU8FaS6Y210efB0Mwxeq3+kwfL
Df8Pe7I8/ro3wrLcMwWPYS77LE00Aq019mNze5on9AuqPSTqkY9Hi3hfvI0ia0qo557NWNGWwnZk
AtLCWO/tWToBf3611vn9dxEOV7EoJINAeH89IvTGL5gUtQ+ijHYxbMVWG5mIyvXiwj1vDflTIehP
tPAPiu2P338qN5WYmiV9lThx+5d7CeozFZwdEmOiL6KCXn3Dy+qiQMm0QH5r/dKSTNT3bUfBZlme
fX1h4sSXMlecH02QGCITyvjgS+TffeqlMCYfzVeHLL8r5uB2G9d2cIbbls9cLoJHScOBXh/yL/gy
J6jCeHmthkHoI7OOs5prr6xzzdMKbwQ7iiFxIsnIosHD7fEx8dQRMWgqcg0MxWwWrCOhX9CHnG5+
5opfv/gEG2alCLW8GpohtUooiEXkHAPoWPjERpXdAb9hVd+lMDTd85oXOflxcHIL7wqzDK/BLM0V
c0WUabG0uWDlcFs4D35JghhbNiS6UMA8lL7evo3tC2+0U+WPLeVUerJUttqCkjB4gPD7hA6y8T5L
ENxIGBvlmlfMqNy8OBob5tYwLR4DQKmGKaAoLdR/nuzBgiN5QTtjEJIWnV7wgPY4O0bGsTAb72NM
TCAvdsZkFXih4wglS+oHB62EPtW8MmQLEXYwG6e8GyjffZypU9KF62STAE3pccRzHrUX40ZWAHul
pScgXF5kxlA6Yvjf8JDqDAszIF5dxgSZV/ko2AZVlE4N5ufLFSjAVbC47eAE1VSxw1EZnxJ4mxpU
wvg2EZRpMDwpaQf4DZPghbWlyDeHozbqJAOOdl4On9whgp4TYb4zW6JowpVLinY8Bqoekhuc3k8V
jUt9vJ8Apg/DLLKsPP8WBjMV5iXWfqpIJTbCHnQYSbrX50Iw4BJNaEO9etnAgM4Uv7BrMWqnI+oi
Cidnj1rRz7rpY4zsbhWtboKTF6fnF9ja7eVJtfUpVkfPWGlAm8z9s8Sdk0LupZMxJAWYdMwc/kEq
YKeEmvR6OGQhx8962KV1P0qG0MC+aO6F7ys+pUDyVlzG8gZGsXg5ftin+zKZyAg3T1MfOOlRLarr
DZm4Ys+VHHKygzInVYYERrq1JpYQ7clNfJuhRjZvZtIUCcAp82Wng7ePLoBkWnKFSmsscwrYPwrL
Z9l+bO5xT6ryUgDuEua0BFN6be6tOBOngHMwsMd8AdyxRcmxK6zzauBHK6yCTXf/Svq031VzVsp1
2AK/ooXzuNBLSVqWP/ZMXTJjBhvHdBm43g+d+MnuLJgQ39oc7MEw7aMXbcjxcjnQL5oZ53t1q3IQ
E1f1dCCIT8Yv1l/Ulp1Lky8EvQgQhXdDYdTYq2Wvk8PcGqM9JvC7h0wwg5k7rpeqshd4g1wV3RW8
Ezt8DDC45p9AcykSJ8L+hBh3ul4kNDzE5RZbM54LBKKrRdHFx1+jilGSFCu5BN9eYLYT0G8vfvyQ
nDBtadP7Kbb5c7jeygo1aeKvA0Dm2YaTQ+TOaggCxOMvH0jS9G//2OWdRBHQaVkXz8HjQwIOd7mG
52FgagUPqKEqtKWPCQfzVKIEovb1wheIvG4pX0y6wzO4AWgmEeNHqQeCyaGfHcTPtgGA/nsYV/OK
yYwRpkBgVDb5xnbh53c2V1aUlKiHFzbGL2Mr5or/sMvI6fp/1U/PzDDKepv78XD7aW35K84HZedg
n/UZWcpL40nCP+DE/fnUojVs2AI+EuHWv3zuZQ2z+k4NJW7uYm7o8ERo+JzoywHA25Yi983bywnF
yAEx7AyJHBoxN1KqmqsvZdj8y9BQGfYyDSS0E/nF1q+CMTJ9VIF74z10oqxm1vcb8yxCjaf+Mx6l
Yv3evxTfMdPaWB1q4RRmXlLUIb6zvuS1g6ztN+P95VuguXQkGc1hXXyOfu2NsN0sj0woJWgE2zHl
7yNmt95+Uu7GKZAqK1p9ukOTHkMDS0Hy1UPCcYpKhmDMY7tU8/+Omr1CllM8nkoUJJ7YHG5v78Jv
23EyfUfbNvVhWuuj2/EcBDQn8D9HQ/4J9554QdUjd1Gf6VfrdNyKdD7JqnyFnzSWqLAFEXxLIUSa
aOgQKcb2IH0vn4dRaeqqbKEHMrN32AN7EhKEc7sLIOn/RMS9WHykACY9Xu0vH8bh6WbEUtNXLOQw
5l83OBEZ/K5p+N44sIs5qq8sAWgPbMCnYpdRckcZ7rG379YdMSN/aUPHMTfAh50e+bW9HZ/b3jbu
kY9wsAkQG0AjOCMRp9CQyNkygI2MsEnXmvS/4uS6f4l+wRiNZmgpFeQ+aFqIDKWcQTxoIaqqmGb8
5S1apaTUPHWcQWkknYGb9J2+L5iMlpSEa9kmBA/832PFsPEixOqo/xYpd9H4KDI9Hu4iVSRmWidI
qBoN7RtHs5S0rWiwhSqJhXQyEW1FxVLj3e/YMJUHiscENqItMcK3GsVpXd63zflGwPpEinUmNq0B
saWc+3RPXGFA1YOLvajJ4iTuVfW/v7Sz3rKdTgLZzHnk1SqBKjt4GFjbpx9kPXve1piBTVn8WWnl
9TJaHOdd0sIQ+dfQDdIxsXmMO4K9TKnmruYhfxswnDirjWaCuprSAv8F15F7q9Z8U55/cpqYCCJo
y8VjqQS90HzFGnh4YhEhf9nYEMFu4u8f7KZaRdNw9b68zJGT8UbgHSmmSiFlrUytA8GSuvRY3QtI
omcYyqUB8bxvWqoNcYEqOp/2ZY1nnveOzLU3faD/gI88//yXWeqPIcRanVrT73Y7P6kVKeU4ZAfP
TvrRKOnOLGypDO3dVdTYaNj0uEiZDqED1++bV+v87BAyhsRqe5oPGr70Vn9Ns/5GWhM/mNxgafSx
yUiEF8sRXq8MYdoqKKtcR6qPjhUhekfL41FqAZT1trBkCBeqap1lUEi0V+FicScV377x4Ki2W2NT
F7VCCy0GzlWk4uoXs8CBV5g+ySjWJBblqP/Ta92fNcgLOEenFNbTnfrtn1xMhYuhroJX7BJ4Nv9o
ebb4u6P8kZKamQhKh7CZxGZbeqNGqJPy5boZzXH+eu5kHO85DBWnSDo9QhdSX88QYELrEvI1jTgK
XhPWZAchtL+w/1py1RiVRXSGpI/83ywjQiKD3PeZgnpKphUtnG0s18Y4gRYxIkMkCQ0Wqx7jQU56
bb0hHMP+WqMffGtUUXnjoXaiYzAVx8IUuyh6/qjhwrUPmKBFgF7kHJAFhBLRgfRXOiwMWxQfNWCX
vbQoWFE0r1EGHddBfLN76Nt3TkMnS6DcVnPTyp4VsNAUtwEPiuR7UxKmumsBU0E7pTVyH85psOhz
7KlS8KE/6IAa0IfXNZNu4bIBFrlvFkJbcN52sBiwQwpdDIVlkbiKHaO9HsEfZ8hUtC9mMaWdVZEl
Qzz1WhStRYmQrf5aVYbgeE0xygnbviA7J417GN9QRD7lK0odls+qE189qarQ+mIm5g0+gegYggDC
S94GP+Wh46IBCzkp0HT0f8dEEtA4gWJq34GAuhp1PG52GzcJCvc8Sny/fZRNZBvZWg8cl5Bte0uc
RdHET2Ca47sqwCdtWvknevZ+Ii9XwXsOyeAbjGSr730Mp587WRTk/7tq2YoS8+nueLZw/75H8H+V
8NmmeQ55i/NOpg5O2UJsBbYZ1paXlKvz0tf8MJdIwlaZpAie0Gp9ThzhaSeLs/EI8AsoYfARrn+T
h8VPED8xsaZ/2V9wav0B5bvhl/bG/vFEVslwLT4eyasdjKDdoZhkVOVGxmA0S1XoJN5lbtNhJFrb
YsyxacDFtcSE8Kgua5pu62Or4yCTQDPcCrdysMOBpwxSIiarrBWqSl6tQDVLEP8cLxCtf0WLfRI0
yyyLhfvjrVb0ebabwapdH3RYI5m9DlvzGTk6iszJXCP7jm+x6AAhsfGOf4eQu6hu6qJjVGyTsbeh
NFwIX8KqYqqSSSqbAPo0DBAYETA+q5WKVPvo7LRyPdq2p2vmv4hQofKCOpW6fLzPC4RrQKMblLTA
kH5oojEdGlA2KFCX8LWXOF4yGEmYmKpN4LvqVr06w+XANHphsJXJppoGnS5Q3zvsxk48/M14QHsx
OzQJQX5oP9uNi5409RUDw+xw7WP/aC5k6n9M40HlYnk3BtN0Zm2OOaSU2nb9dlz7So6zTsuhuKNW
/n0Edu0rC/BjMAAu5L8eAYwhw/M2TW48v6yn0KmMTTHzzjaLvh+4wSee3uuzbWrPUSUgI0PhsHI5
phEBhaFYu0+sxeWWeAGF7SI7F5Nq7OaPhs25odvqRaMkjjCMZtd85e30T/OtXZF5kqAZiF/8V1sN
VfrazX/QTQRciRKvBSh8B+BokswSNN9zAHFhhsS0ShQxaV1b58dOPBgxBXbI7xcE14P7kRQPfJoE
qQSB6rFqDUJ7l5yXvQnXwv5Ra+dgGEXTHxiXwRsor+Y9Bd91lwQZPCqRSMBU2UBIrG+3n1g3ZIqP
QLWjRf89LGhhaUCTHk0WU5V5GjVfG2xuAGiTzAsmVrarykFEX7PeRGogmnzTf2UsJ1VRFZK7QXdX
lbnPI+oGBrJLSt5i6RuLP+fcNf5V8fw/ysF+mrQzYgdMiHQM6O+oXhaOOOlbRhG055OCnMUc1/uY
WU//ce29qWgA8DgAqAcqHadwCD+rPHMpv/CI428FWnt2F+opwAu7LXQMX3v5xSk4yPnbvP5kDQFP
6/lPOb4eaGb0d5SQhxFEo4YUtIZvRNznvcWnkOgYemKYo6PpqG7AmANBWZGPoUbccQtHElg3qLHa
B54Ot0DtQA69mpECuc54W+XnmLTY0Eg+vz/g4mU5DDdVFg56X9JK/sJheUuYOjL3FZuGnLx6Dcju
5RdW77+nKa7pCaXAczyFQa/3bX2mW2fQoCsbQO3zcjASlgdv0fryjT+w/EG1wFPKpu8mEGaHMF/b
lpxZWl/VxtndhJwWl+6H/3zk+7eoTWs6P63qq8CxCHKAmLucjvIgPcuW6VU0mekYvQhIcpOHxmXL
K3aEdMwdjUvAnRlH8nVXmZhl+0e/Lqlqjd5tUYSvRK05gGUCgPbxkjck5RRo5zpofHkU0leb7Gtj
7v1uf1MBrT3lHod+xAn2InTgkWZIkorDTCpsb0yWIR//VX7ZemFv7SYGA1mqtrv9HIc4CZBal0I6
CSq0yKq7wTqjvCutKNmn97hKBDY1Gsyy7XX3KmDZVewKmu9tjiXsWvp77QHP9XiV9Z5yEbHXD+yu
Bh/jPyTyvm0rKgNLDuS5kWPHOZmEOAoM3loe+QEfVWlwVrGFGDSR1EpqWHqiQ56U+ztIi/wq3rEo
wkL5zA37QVeolBSsmkqBTykAjuAKll/qcbiumCwZ8z2H/PmnyBdVZPADwqk+8rrYQlu9TCXhS6Ti
a+6fIBTsSLlmiSF2Sbb4jlGJln5DMaJnLm99iwOoz0Tfl9xfpM/WRjfkMvieeQAhhd6u7mQHmO2Q
P+LywiT/lwyplDao8WN2UDorvXPLbSsj3TgdUyheOsq8uN2qgiXuiuyCbSuFzR3zqv9BTvQz/lAO
GhJ25xa+aT8pKSCdnKMSlHKsUJl4+ffJ31VBaC7k02iu3MYbEg/+YhWNO4Z9NsNJUQGDOgNUcB0c
+lELfh6kH9gjJBfgVmQSXfWIoz7S3xhR7vzfuXgCwjY0FoOsxjcgwhhyGqCDTbeo64mSce+Sifw3
zaLvLUHv4gFAoLY/RL5I06OO8+bvEXKKLbTpj75k9q+o+vCIoBr6Lk8KF5anV8juvZ6c0nqa32qD
3YJuqJwI2/LNGNngQlofytu8mqUvBWHvqWGm/bOZ+qcpqKPjXwxeEuUMj5nKnBHCzYyeKFBABhqc
VwMJs6u7XF0YJVHMXrwMz8sNHCWbHu/ghKeWEIKX7M0N0TETi8zKscDs3KmlPk7ynU+5R12kMAVl
x9O680N7lEqOCGMOIOvgsqA4jY7cllWv5VnmDE03zu8n/WkUSq8OgM7iTGjxP2arf4O2ed4wGleS
geVwY1EvfkUoR6hJko52iFcWW0SIFbX5Bk+AjEPBS5MlV4CI9N9QmNg3c9n0qGxi+c3+Xz25zZHe
NmzSUihVm7NCktntIc2mBbXJKIa0QbSaUxSHd6jsCWTG7ok6rOWXH5xf+oVmOfyWHDHNtn+RrJ4a
H7JJJtq1mlfCOYVbQ/IQXfUdWtN55My0mYIs6K+E164YeC6F9LO1BibJbmirRfZypPS0UgWOihXs
HY88J2C1M6aWbLhn+gdrJbWuGaOh2slcU21JoDDYpvMyEi1nKyxVXpluxFnq1Z9CxItuQq9W/bM9
DiCBSrZ61GwPXt9IDuPrnoG1KBoYwc99zS0X1tiXqYXYwgJgtTAM6vSMTdheyjod2ZufJK7hGaml
MLKFziwRflDocKsbzp8h+HGr7N+JXC5SxkJkQbRGy4nDgStFvhtrBr3fAjF5N2b017ptEiJf3Ow/
OnOHk2Qq85ZiUeGkqaMgAWpwxwO+G+Hw/oI7Vbs3LrTUhWxMpsM0lAibuAiOq8sNIHsc1x59mJHZ
daozKbH+hTI4x9bCdVCZwUG+ITbFpRH/hOai3Xc90fidGH5Fjx2sg7BwjMpSHs1AXDFViDjDEt4i
oY3ZBe42v0e3IuhmFRkZjCtXVbIgZPRWlg0ITu7UwqdYSFFLxNACnHwmMh6J01+dINJRUBNv7b/z
nJbkA56a8fNiZFRvpHcYFVdc8oQqwT0C8kLB001bqFQTQBqfqa2U5OIp2NVRF6tOQpzI0pwlVd5C
XX3KhcsfwynJNZrY+vXAa6d/AH+rYuTfEJzt0hHRcoauEuIVKiCLwGMgVS0Emq7SSE7Uk5MKQgjs
xDP9OSeRX8wac7U2MayaSNAnwUygHn8ylAWt+J5/sXKb7pM6EtI0tpb3avhsmeXiMlU2vuUBM9s+
1PRItR3oXMXZxYSEh7vZr5DcDo2ILiCVB1klJPXSSkYQQY9xh/ieDBpEEFYA/8K7nOE5PLNbQlj6
e7yQiGFaTi/5In127YsoNlqDOkN2y4tUL6OQadJxcTBV9t9DH7hliMl6K8oin5n6NVSIMuLscdkj
RVp8QQDZHCcutsRkWS2doAnxWJ9ht8NL7kzW8yLYy6oxTP2jtjawic+/LEyRHzbkSZ/3UVQ6Pg8X
sUt4Yyvk/InwIuv1KZzaWT2REpcFdkOwoVg3INIB/V/WWSEODb4zkPMX94gyXZQuyV+1NoFU69fo
Qm+PlBNaDcaVg+UafZuj6ef0pwYxcBiJ1SZ72tS1zBWc0pwYSqHTtVtXeGnwO1tfgyX+9dFSxCzy
yhd2/3qRnRnG5eAIbi6bbrncVBKPYlABTJauWMp2Br7fsU/IwKBONSCy9JpRPBOFCowEy+oyOd51
eVMDg2HDBKvCwoozrFLY7NGYray87VUhQWUxuncUwshNKpHqldwQqCZWK1wILWdl1czQOtYJT9cq
ha8VXKQJsAFuXqX5a0nU2xQchJbtdC50Fr1Hjtjxlu8+kDFc+QNzkfpFu8sbkT0M5SFqyhkNd5a3
BtBuDOvsA2d1DELroOJUxCuaQ5pQCPuxxJZ6Wpd2WvZuIuGvJqwwx46ti0nwvAttQNuex5+BuG70
coyYwsAhKM+pHudosqEeoVj0Wpl8o40HhMUV7Ps+KQa+/RgisIOrO4+5UqwhmfvtFDbEvHPTeRj+
qA0p50kLu2U9CxlnzcKOU6rVO4pDK1pgkOC1nOD6pmumuApX7IQ+vnyg/f/cX1vgIcpWTBBfEdeT
8DHpAXGF3zDKODfUaHeBDLvPNbXssV6Lspxpe90vDfm5QgjZOzxEotiKcjl7It2bo07xTqagx6yh
eaek58wSmXiYgp7CwtT97qqF+sBaDehTlUJEM0F20z8cUpjoRtcvWNIzhqa4mK4SwEeQpRQK/Zz+
dCKo1MmrmbqjQ3/E51HtnGgHYaCG8MCRs9oonSv56dp7ivBiOD93I6NI/q18DRhmnSrAx0rHXvl8
ZR/66wuwuQO2l1UcDhl4QPP2X4SVcy6lDploeGOla+c0pYd42Oh5+tJxUCCnjQFFZTW5TqgP0IFY
I2gzNG1Gku/ZSttGcB66bYLor8RQFjrohm69e0O36dtIo3vSfcBYsrGuJMiHpIUACilYOPTqu/SW
mPryejZzYOWCy+28tJYKivjW3RZjuH6bsVFQbCATR34qMU7dWjbLjcVVoVq8iQ0pWZqXT2eAvA5w
bSab6hOCIQ1I50DSsNzLCAHXkZ3/Z6ubjeNRqXV64kKztdVvKbpZkS+1TL8krZjtpJd6cLvppPC7
f6bywOZ4Zh9gU6i1OnMfwIeHftzmJB1OCQl/fpORwFqlXtZMvaK86tJal9wNpg1YZdo8p+vv+CTD
M3oAsiBDbvQSdGmmWsuxS3xVbKBkwH/r2b447NtzwgRFsYU0NpLV70h9S1pNr/D11+vCfjiYKb3C
SzPmoVIMuYVurBai/MJX8Hj2eixXhYw1LYJMvDg99xirMeLD9jv8FuaTjRljJTXdhjPOdHmuP5/j
GFMZ15EbdJl1z5eK1bBJ5FuzHz93LUI86HetrLL2ghO3oKXElp3nzQm5OAEJvlstcZJSPnePa2I8
9ZgbDTyyvEQZiVdEVsGfzbPTsZ2rnzhFy09AA20twush8j9DtVCgOnkLUVIL0OZQ9rtQisVb/2qx
aKiHANbfc3Usyh4sUKOHwBGMcJOupwdiYNh53BxOU1Ba55jfAXO0BpLUh+v+XCktc5oxyXpxx5tr
j5ed9C5Dm9QguFX43Lx/g4uRiIosAhXGHa47kzjrtwJZmN057d1NCEEAl0lIhs+5K3I4geSRC5Ya
XAIxki3a+nXwlr4EK/0qEsV7w4Sa9CYPMfIZU7O/pgN+z1svXPAiLrzQX/NXIPeKmhAGSpxRV6MG
9l90PwUBnsvlaEScbGULNwX+H1aoC4nz/aPPG9i3G7RytvZsM0MBFCVhsSy27erOmTYkO22y5JAq
gtUwp/c92hvqhK90sUKVwV0brPw13iZ0iaFjkUhBfWhrS4vOK84PVg6CBf57SQ9BHQuIcXulLY+d
VxfHtQo5FtiXvAIETPWxnZiHMT5JCy9g3Gl60vH2BNiU9PxlU2Kp3tCzVjuoT2pNWr/T5EL+B370
oMG42C0VzLoXV0cmT6Vni9z3Q590KCdD8TZx+MNIfmBPUYj04m5OvnIS4MYvspXbVT5Z3WwHlstu
SBGhufDJM4MfiVQVXYqmE9BiKKkuhx4oWh0Pm6qdk/U3VTyWNn55kY7EkFypHLUDfztx8owpyZh0
0/3E5Fs2IkUcM+Y+Y3kXGl4WlZT5Y7vPVnzPK3lzKcO50D1jWld3EdbgQN2No7fjUfR6ZKmHocYT
4p2Y3cfwR0MLWoY683ARzagZQ2RQP+Cw1vA0nQU77CtoWDQTpjHV+KIKKtZA2oRMXsx/t+B42Y58
ailA3eFqjCIoYC7lcg6n0EXlXqgfgNqpcVDinXwE7YTPMVypOS4WrN/mNcm7B63u5ROSlUQIhI85
n2x1ctLWyuM5XG8g9b8tDjssak+QqvMxdqShsuW9w0gpDNroU2gv1HGe2vwTd3XFFWGjHEOPt/Kq
/y1qUw5R+kyNlS1/GaBU32yA52tQdiDbhXa8r2SDWnJQ1Bf8a4sZvkmUGP4hFN2vrNAza0oR/oPy
BRmBcQyMZfc4PsI4vzEvGrfzCB95n90m05ybWZrbwZZVRiSuWZFCK6+j2seSJG4tjz42ZAAh3KON
liT5EjdOWkvd2w2bIVlfP4iSy6OiDOXalT12tqRfGayhCLut4Lu1/XNQmqP5JJUl3v1HvaODTBVS
7sGVKgesEgp2d3Ogmn2De4fmfbhfDtYo03A55xX4GABgHY9hJmMxoBUpcl5wohCfZwqd6geoiwiP
xe4TqGgj/tDenlAPtDB+mvP74jpUaCaXKm0cNFvl3YOztW0+F2sv9olh351cwAmT6fPnt/TDqAgE
oPUXEKh65VNVQQ15n36cE5lh8+Jz/F+2w76qk6Sx/2CXYtA/hIbmQT5pytMEaisQbZ8YJD8ZA8zx
aDWBCZx3UqbHwdQ7PAKTD8N54uIqE9tt7Wbp6QvWlm06Nrw8KselN8OBk2qjC+xi/oS4UqvMNH5E
ImZibhNBssGe1DYveDx3cSKseUgaYu2ol/nEI8/j5p1gw6KbyigfrGelf4w8GznHc+hyCw9ag7/r
tIBGBCUeyMGjW96oM7YM055rUp7a5VSAUb+e2CMA4NH6PdpYW7OSrpOG+NoX2lXk77SzzuDunMY6
gPIzgPPIbIgatlvh1U8FNxsCbkk6QdnIrKM4/AQQhiMVU0mtfsY56xTKLe+iCWiNrFtvvWjouTou
6bCXKeduZkYumwAG7ju703lEjH87uASScolu0pC0cBQ3PO8tE0B/Eop/2yqg/vX4ZE+4500HMftI
AZdqht08qXMF0c8Ua4g4wgGHZJz6fi4htoLGXx2t4buo5k/RK3OH+7rJnpcxAcvw1Rzg+oBXVn9r
XMWoohWDZck345Gl0WpD+Fdpd2Xpsa72PuitJontTtc4H8nJN+NbQ/I7Z4sG6/PNZ8x6AEHTqhla
/SaHxD315Zvex8VHRka0tBZzRnJg7SDmUiHmcNP+QcrrFOiH6sU+0UYdS3s6FwfyCz1uHFuZZsAj
PzAupmQ2VkObm7z6biVR0m6qDvgu7G9XGasE0AJR7JNReUKrj/EKiN7Vz2VvDcA1UbvNddt6OYMm
JN0zf5sHn/4yAp2iLOlqCgwf/SiwriClDd6OtAZxe36eZttKNWJq1B1vAgu1Z91tVnFobFggJ++p
Qyvy6XqCABt9pwmbtLPBMR9z9XSz2RkRN2ZHv/3LwgruUR9j5htdpyS+SESmvWmhFLeVQ5jYFzkl
Bs0Vmv+ZL8hpQS/NroFY1GvXYQ58+UaWGATRXVzbLOLuU/QNk1xI7RJ0Cc2oeZRg7buscwIdxRM8
pGUQgDGhyuNfVahIYfECLJUkh2USRV1j0bVrznH+FfYBcsNldXEYSlnCQRPnxUtRUWV8gIUuLYLn
+fsSc7ZpX282aK6P1Zg2gz8xB7khcsFAbOfzQHotkewbaft+SnPiUf+Kp/g5eA2qGS0C/SvquH61
nWTuZkpwnMCMSbtO97Xoui7NpG71lUVwu2ImuwZu+eEJ22h3cx8Vg3p/RMAzziFC1UK77JGLhCIF
KrNl33dKQO2uRf6xV/yP8e/uY3V2pcDdObmh4I4SR/pS0ssQR8FRdPqezHsTgxv0b3hZm4z5Twnh
zcAbjqsMtt0YusZoX2v4q7XffU3YfFylMRvqKZfDMnHUbD0awjQ9MgPgHVzdCOn2mp3Pk+WRjENA
C+Au+fsS8N/9aom1G6V+O09S+MQYGWhCzFZLE5ut43XdwQ4i7ZAaerfGiC4bnchf1eQqIM74ojmn
2WLZiTzUlcd79dgVuPmUSVoAHVihBV2sWpROh6leBLyXTL19rv1Zn4KcIzzEjyUMswe+DCNdy7Zx
OniODlMtRL7cRcbyILXQqNpW7vLCShpvzFHMij0Wy5icFnUDFn/jDQzBK7J819hJJuon7lgcxJi6
D+ZPi7N2CoMVYJqbouf9y0YB5a/j/cG7Qi/5XZF7RKMXcvR1jsjTIYNNHQbdXvEq91Waq9rzMIlh
cM6POSgZKvH5Cs211qSLe2NMPtxH0j664gcHreXVMqHLOKWvTQM4yAQj/s7L2OUK2Gmp5garsoEG
OEWkwFlU1rRVllKLifdCTaI8CLETkX9YXHwq359u5XHsi4NeYviZBXtrLkaMHe4i2qW72YinfoUO
Q2DZcScad4fcG3VhaEMaA31qy8PU/ngRVCRGA7Af4SayC3a4GjcxbdekL3udO6FmAmOyF5KgW87o
aKnZjMcl4/f0j46THSXjyLpUyOKrx6QhkJx/1YB1KTw/JaMBzhHH0GuvV2h7Ezzcw2G9UR5Ov3iP
2uEA+z9XQDu0wEWnW7BosZA6tGMEPYoZnwvJalxmriYV+M32YkJ1lRN9EwOqKIplXtM+Nt4MueIT
5FxHUsXmtyXrYIMtp9Dnh0obKQMWKFfg/LeuKrrR7mmE3DzZIpRpHvBzWujIU1cAJ/AlZch7o7B/
8Y+3upOJ9CLBJ7ZbUzeOJ06BJx/RxOku1TzwZsu9WNNMgoWptNs/SjkbwjJ6XblMgIIQiRy/kzfT
H+6DPllvRQ+5OLMcmlZWEQFKXcw30lKv/W6jdWfF92qJpL9KsnyqPJ8cqDpUGqprPXdOcsw7WL5D
GgMOZMGnu6+hF+itFQqZ3REJXdCYx7ge4hprIy5xQhmAQeeIOT/AUTzSRpVQ5lHpVXaoUc8bQKiK
JdVKXjz7l8LZ8l/5IdrclpdmlqepIRHWJY4iK4BEzbyg3tK888mOQ2VDhCI2hzHdYy+DiD/jta3o
LcsPVCeSVe3Q/miqmZZWPO6JcyafLAmNwc1hkate+9fyHHNgUbZ//lGX45XUDg5IJv7+lsUbC1kj
k1Awhjh3mKk7Ed1o0tLtdxDOEjPAJcTrouFURtoN1bohgFaU3CHl3dEAKymnU+A3SRVloUBj60dX
lGj277JfGeoJssm4iEBiOh8av+B/pRVnd0NSsqYF5Rxkx/fAa/K92JzqNUXcMHUwcjqomqa6l2s7
3wT0T8pBFULUwOhCLnFuBCUIUIfEVDK0vfhLnF8jhAPsVUlndN/+HPhWfPTJsrbqh3i4U1zsn2j9
TNF6tkeWgW+4m21UD58fRtcEA4Xd5FwVqh3FSxzO5pY6RPJRExMhNq1azoxpLLpXpTfosaiTrrcb
bI2fu1KqwVNB9F5kYn2afrgS25HytrOrlm/kTYusYOiHKgpkxqhsz+zkH+WPBiiVWKxzrP+piYBm
yvg/KT+7z3Cs8uogLuP+ldVF5FE42PvIAtzr7esiAT/t6QkpcpP7t2Is330JrNRxuYXTEv4GZfjn
x7mhNiOj1pwwA9BxOCYXn9cy7rsz0Nm1BhWuIVXyRQtXUoTbLUP3JyU0OAmua77q5GSnvD4XHRkH
Aoe7uLplUUkFSVbZgWcHwyz5BYEgcUJJ0XyRoU41oXTrNvIzU+mQAt/2V9kd2Mvd4e0i27znJpE8
fu4yiG/p4k6BMVlTbhb81wC94AlyC5OJ/X9VR3uDG7IChtbx4BpvAxEhPd2CXhOEsor18Lo3snXQ
6MlZIR3JMsrKMGrYg9pxCBUZZ5Dw0fE04l3+yGEIovNxGAGsKDc9nbRVczXROQ8k4F2+WEYKEy7X
Tg0df1p74uHhGH+SwrV0SWS1XFUwxidT8Pve0t8iXRJbI80Gb3LlXDz6FoTApMIIDd2XREZAb6C5
n8pJEJYxE7l27eb67ZiQoZoespwrwYiF+H3jcVIlkdAOKSzx2ASy+Ek83bhGN/7YS6Bil/yNtsAL
Z6sQvQiMCzgmPUntirnkpZnYXEQcjYi3//yBE9ZRBj3u3zGvfUxNhDCpn4sFY+RFjB07DM6qhrpZ
P6aVA5566eZeh5jwM/7DdLUAQmn/u3El6TXtSMGsMBakNXrX9E8b4JOh8ckjheLzyCxF8gp23bZm
1EjziaWlU+C0iF/SUVg8GCj4Wi0hy2ld+sqna5uTucIu/v03uSdob+GzAx2ncUcIXmIrgABCsKFD
G0VE9IZ9OLG6IaXETKQMRpIOhgARTpTaFeV0SK48hXoxPWw9dPn2p1fr55SoSPJCA2BxSOKt6E3A
27Zn1YkQIMhyWpzDnpFcTkze7Ko6GF2ulTQbiXarcMxiGntb7A8RWiaUPlrSHKAC2Zm5iiNHJ9XD
+s2Abpuc0K72axdWKIds6xQwtLd+MtWSiRXe2fbPBa80AOYcfSrU1j8JQQXS9miq/W0N3gUzGuP2
fa1+qtrLJeCc2p7fKreeuDeMfpiAUayOFQ/pxNJiAH7Y8m05hQGds3cO4HfegggaL7B5Y3bTtYUP
+FZiTgOQBgkFzqorf0hzXpnUxnSyp/gsGgYrXsDhzKjUItIfy6oK0whqhvXNAHicd9qUK1CvheAm
jdAMWWkDIYPY647g0zDETB94tEpPe+J5fJbXu5L7dpLv1bQiJVZqbFbaYxZaFoKSKB7RBLRncDSN
5V1G5dvwryI8gKAuy4ygewRN2utrRA2BSsCsT7JTH1Kro/zvcAH/rXtArwICzAHmPYPLgfLZB7LC
9Uo2mry5yHMBOd3UQ5j9pylX9T/NsgkBcdJ0/K6r8JvDqR4Lfxf88fhQwYHE32i/kH5CADkwMLgJ
yHG6PRtwqUNCW1/efTSir1QHQuZQdiANlnJuoCjZ1XKyeIcmU0RG8LtOea25ta2EiXF6t2NxTeMU
6MTpHUVIm1ZHyqUR2KBDak7pzn7eQUWYgB42QRflwP+Kpt2ktgeLzqBVWVlDYQ6yfiuPFlhTmoyq
AejTQ5ZuOE//zQlD2IUR7PjLqFfqqt/ZEkvcKWslMntvFVf2nO8gf3tGcCN+jNlPPboxrHCP2hbr
wU9i1AakzFUN1e8lcrjOGN7m83VqgGLig2fHASESSFFnORm1WCCypoi5m7VK+OtBlZNkJIk9rwei
lokwaE3bINP3xVYE92tStMOSjUE9dt3hpZORQqNCxOU51mk4Bduj/6J96Q8xX0iqBgdD/VKWGVU0
/LDMcUKA6iDHnc3fBAOgzaqsV1MqEqMiDsi3o+wjjfxLoHBZcC3PCATPZssNPH/0WRvKRQj/tcZ+
G/W3Xtt8pEO4iOb8G51kiGn+pIA2jw6b+UUROq9eUhnQBAtDxqm9Ur+MuBRNo7HKFSBhUUTe0jMu
7VvM/Z6WwEjmTB+lUkQwLRMske/8LDmJEmyaTXKTbEwgymTkKyTv8GSAv6nqj1aS7hlN++yQgWDp
R63V0FvQIKhWvSTxjaD7hAzYUb3b865r2CCW7kIOj/cXSiJuUI6IVSBWUPWab8ngwtsLpcBlK/99
tvWg2aGR796CA/xoWkc83+nScSlNcBLNw/FAQQHdWHFQgHVpqQva7bI2AGf+CIXSOnj7cn9n9Amj
2YNsGz+7kH3ZlirUJEM0MwcTxw6cilBFesHJVI2iattNS5Rn2b78CVRYrzyx4KZXlEA2xPov/eTJ
PT/UgqxXi5WgJYsCWfmEj1pf4pw7iYSr0cyUa+R5nU7ZruM/kR/pwiMehBep4C748hAqQrJ3+H3u
b+WVniCcP//w4ORzD6CZ6Mw7dXUl/ExMSlfcRhqk2BLsxBMlvSZNTUrEkxEPJoBbzXS/p/HD0pdH
EHIobm8cobpy0Yl6Jp4w79grnKwCJnYMm1LwyA6a0jF4x3IphywDM+sViYlLQEpQHR5S6oCyle/e
wXNYNTwTgbZmWiIrhQ/GS+KYsDbl0DI3Eq5ZbiK3BtX8ypN4Ki3zV6eQ9bf6hkePqOGlM/YFFTGX
ZlUWM6tw2+PACK/iRh1s9U201vIVF9HhS/7R+f/Tite2X6Ra7p1m2JCSgNpF8OUB6aLLb74ORdWA
uQ4WW75T5DxezxnRtRFVtRazbUmhfCTgnTE8GNQZJF720nzSflg2RxhpWHBTrS2K9BbEmRcRJEnz
ht3u2vwHlvEANPO4PqDR758b3KYTy7PYHzDxis882t5ZVi7iPjyC4z1B0kp58WaVuC9wraNrTG+5
pjAIcyoR0FV1OPOtNdq1q97y/nYSKPrZqFGurdcp6p2PzA11zywQTyFCjSJ8WrD3nUqueIkdCQLC
V+3NIKLIO+OWwT/SMXdu+hrOItBEm6cP9qinyaKdG6kwTcQ/FwDYRnzIDF9dCGJjxew6i1ECF3/G
yggXzjdhASUcX8Th1iUJaCgZxseRHjoJEIdSRZ1aTq50h1XHkLHAxqQere2ggWDCZdqO/TvLMxIH
ulO1u51+rR3ObTscStMtlCqexjwvmLZSXQD7HiWodQLi8rBOERc7wHWPB2x7r7LKpeKvtbti+nxR
pDnH7Vpz5K8MMx0KyVSeE7YBSH5go4iPrtvfjyoORnfopAKD28dGjBqyYlVDDbB7veJga6F759xw
M22d8tFYqcU+Jpj76lRdV4IiYlJ1WATZZRgezykuEDI+XUfA6xmXi0dJ+HjR4AvBfPuajTr7jUJy
yZEWq1AZDtbdK9mmtn6zeT+MaZ2pSHKFzCMo/SSlSip0HCaOIaB/lCVmzV9iZ3UyiQlDUy8WdQDv
BJbXbkUSD8ZK5xmYW+MepNd+v1umz/b8JCImxbE3u/oel78ocsLjEU9GOTTWLXMHDlwLHVyXTYhT
tR0pyGDUwldS3T++olnWdHaYJTAET6xUDL+xK1cpZGQNytWHzeohrA+kFoiQ4tV03HqhYadeQSFd
xkAkyA3B6Qem3EOLsSCPvgfN0rd4Fu1G+A0Mte+uSoene9g78ljXo37m9pgGvPxbJq1KxZx1ErXN
YwDFI89ZECJwEMd91mfmKWD4J84vlLW+Ug2Bda9SHvs9oAAFQU/sbj6icUwJ3PCk3Dl8i4wwRUDf
zRvjAzQk7Cm7pj0qfO7CXjGbc2GDsNV/fyso51I+mQeya5bsgFzDL6H24a311RjAImwmlx3JBZZB
1MT59FjD+1A6Cs5rZyTCRQyYuHt6PHVgW1EegPw7y2xs3hllcvX+4WsY8ANxUktLmyUJ5B2jw033
cNq7CWElz3amFQwQogz7NbQ5hjwU0BN5bpZtZowyaQEQKSGfwoHODAtSUu4IMx6Q9GW/MMQ85fVD
tIPOFMeiF/acrHnqZ7AdU8mYTN8AOVUB3BXNohxrLWPY9YVjEkFiZqoVf3SKVYiu6qEq5CEoPxtw
9utlddi9nZ1l4KlTVgtLPV11n0zbxHP5SVhlhO6iU/ja6RMUE9LAAPm1bIcI/8LnpxRYmqSAROHY
MLHzilr5vRQ07CRVwy8EBm/a/NA+pLtEXEris43e30oL8ZeALB8gru0qSnfIjVViVdx+IZPIivkj
+RYKiwA1Ds3mAQ7Y5OETLGnm3ccY4oGZ/UUzQyNUMTrR7Zj5UbVwoCSb7NY3aB2Qu+AH02hCpnLU
BvKX8V2bRT+lhILiSWFZj1qNMHpTcZDv5WLauZNFFS4hu+QP5lGO2bLoUBzBGbA4leJ8D1422XaN
L+wpC6KZUK9w7hzAb9HLvSnOgm+PIYS4uZghw24o+C9VY4XG1BQK+TmSk4aPVUqYJAKV57zEM7Oo
HUOxvobt6a25VESkEeVfCZWiNosp6oMrI0lrTwDH2tVXObvR9Enq6L3LfEFyeFS2SiErj8QboESF
o7pjlF5tH5QRL/nygvu3tx2okXS75UOmxUTyKh6Ci7yxxhblchK+UXbCFqP7rpoFvGNfqvBcqUsz
oZpTETwapdSQvD0VBlbeuyC67DrMTU9hMHX23V7typAFv95t/gcMdapx5XTnyX2MRn4bjvuyfCUy
DTci06YQOWqGaTv1UJlM1bOFS7luOmkb4FR01MxJaJbIm0Wb4uSDOF9+/XlKxYH4bQ4cFm9nE1VX
JGSVYW5rkIGBqaA6H6/bxHJx2dfCH5pjZ8DpMI9D+tXSxiYG1sJOuOevRzX5xdhVmok5Z9AgH5GY
zldutLerMBm4A8NJhAVU8cDGhA7/j5RQIQ7fL9fCnR3Hayg2q/PqF18nMF/OvM9xMkKiyVsgNzw5
pZNNHoQBvg8B4W1pZwd5FjmOFk8W5JvxcMYnq2wPhD7aMVuSothm9R9a+YPaDk1f3pILsG6xvb2q
A2IEogsPSOXbnuYMAmz+2sEUOWkw1NvLvW4oLc7BGYo9rYE9CCemH3D4QMBu03dVQtRvHRo9HDcl
YiKve2V1/7PsKUaCho69IzkJjmi/HZUTR+JoWawkIGYkMa0QFPLE1co0corwdRiqQKsQoHbbjNuD
xfJVbFwfliYDZabR0VDG/KM8QRLiQghUdd3LwdXpHObQ/IiB8dKk2XHcaFiA1QkImJ6nmqGQiU1k
GujiqJvItPM4zWqJJ3ppJSy3Ooe+eFX4nbTCuNPkM6eZWrKGw0/p3Ln0ck9MwwtO2K2DQa198TUC
SToTU8tML8iR/jYUn+0mGZIapGN0Z23zWnSkh8aJ6M7DxIeGYtoyuTDFXy7egKQExCN87nfZQGRW
pYDpCN7H5F/dhSvqEUyKg5F6itb4BGHUpbZMpmL/s3zeKH6OUjQJ9yP4Jh9VUdsB8wrlZPqmbCWy
jEBnds/7YMzsTEbrKw8WIdvvHvXqAchUNjnvvYy9jZ7U/bPYvMJwBxcqzBUxq058ywMJva2mC55e
abdpTb8G0/SLkAIG7sAOHJpItG+B2ti+onvJiEtMn/9x9K90Uv82y99WmgMNCqD9pq0HegyWAw9g
aQEXUFIdLE4Su4PvBBaauv0rF4d6ty2L31XWsI4sh2M77Ko0HI0ILH5UTKzWb0am3adO26b7SFZV
mvH6SRaDXRxplKXPCI+ikxqykYOX6FKsDrR7hvHZqcZNdagmVtoYiH+nlJ9H2av94nQiD1ME8/1Q
qQGFS0cY2EJhxE4w9GbCfSYrAowau/xWKZzAwwER9FPd0geick+lQBPK0h+6Zc5JK1HbhLDIkBy5
fOY0o9p/QXTR28YOErFBjzSS0hNPmrWg8OrkZjVNCtIidi3iNJz9wJPaMMZC9R682hV8S7/6aQW0
QzQoi8PZc5ej0uOEQe9KiN7j71zakOe607Nw7gbrgsbN0gqgsmlLu1aZSqAm5rdPH3yn0qtzbcq4
D0fO5NDrR0oRWMIx/Z3la64MqhxCXTFNiYnh/XH1UMOQY9QdicZFy6aOGH0GFuvkzUGWDcZNDvgP
iFVLQsFTkW8PfdiPvgzBW4Nw3WfU76OcvACu0gJDj31H2VD0duf5jqlXYdiLGXHLVknUSK1nLDha
lWpwS1zOtVHcbniiXLG9MB+hf8395MQUZ/eG/+augeDY764AitBxvDdGbR5d6+9JDzm/6mjP72SX
mQSqYu3+U4yvtplL4pywRzDre8IZYWxBjaRJWvZ2R58OkdE+5++GIpvyJTaH2JrFfhNe5+IdynBK
l4OAGepFEcaauCwKRG5afKcECmToB14PjaeQ7dOesC7Ek6pPw0UYGVxyKKCnexkt+VaZZ9j7xkbF
4uIF84wdeRlCQwmtVcQhK/WGTNWeyoQONYWG+N3JvkHPadU0IjSkRfgFyWiWatwG8dQm2ZkauQwx
7pAUVOn3ZOsroU1sTFiffb1BnkNTeF0l5EKsjhybuhF3nBkXPRVSxNZfCspwSaHpKZtgClXAr0JT
GZEsp1/3j6wgcwHSfj9w5tkExaiMN6B+ZY35f6E20UI2svuZqUW1STySqSXXDqkgkkOXzqg7U+09
8B1Ken4zq+FMu42VAu7CnVWq9v0aOVjeJedx4mlqUNxWnLOqCFA/oaDG6FN7pCDE8wXNe3wspoE0
NmxghiV6EERzmbb4Z3SSDE14HUj8WWg0+nRz7xriwrmwGDCyFxAWoF6MxmZg+M7BN3mBAcQq2G6I
U9/Qi10tPnNJCn+NsjejjXU6ZJQFRLk1D7aJe1XZVBQi1+N6gZTGl65H4kor7+TBMiJGHND2viDj
zvB64wvXx/V4Ufr/M2rD/ZG6WzUjiHMVhvU4i45+VHKAb6fO40jQYq4p1UBkRtgvKUBbGk/EC8fj
fy6sYBniu0aKzA/6fAuCK4gwvVKPElfUNLgU9R5dsBG6Et8AtfI3W5YQfFt2Xj7G81LIW0mf08Eo
7ODESpfKxf9TiV/nlEQ7/UgN3ySdeyTBAc7KBuEJM9LKHRe7p1tjlWk+GpiEC6BI017tZH8m9LIL
RFENXLtTVoJslT0qLYlt6Qbfy93u57AfbgnOYHeOkaR/S0iJg4SrEXTzviVT2cUDIqXPMlVMhukf
jXyObLedC2bqt+ZQUSBYaBi0uKZqQM2LMPQSRLSMyAQXNsMxzb+nx0en504GYMGPJqFU6eMoUFl6
f1hhDBheiLKU/NrlkFeN6teShoNhvy0xeNzXRLH8mTbpjKtpu3dZwEcqEsFiTjezalgTGndIS5Cw
kXsUDs8FByfKveShxXP88duTCK4tQQ3P5YgY7lYBEYa+tKSMsoIcl8n3CscdxZnGNXsibloKQXJe
iic+ZN01CCjFA53YFt0OqXtThjBQ4rkcyhsiUHpYY8+b5QHfQL2fxfOM+aq3zmljeI9yrhRdGfKi
zprzG8ylCtbU90XVaDeKGYhSfJZVzQ9E8SsfLP7321EDNfN92O5HrJ6LccHbwty+1AWP9kKpQxHA
nh/U1efwamgZANV3+EF+LZbm6nA1bPUtf6BJUQWYkA82gdG732cNoutd94tmAUezzbkOPfNZwzCN
6lBUGW044nnnOUDmVJW5zL2blPGFFtxirLhW31tdVj+MCgxEjuOJO9xtnn0m2UImMroUeEPFvLro
c6WKnVxAjsPRZegmXL4l7lbTbdCTO00egDbmtYrj/wajZ8QgOGyGazEJ57E/AgER3pUs8jA0YYrU
PvMOID+yI8rFyShQ5ysfxLjltg4373zs/geaP4mtzCM86RGVKjbc5EuAkFx9Ln8lT+r8vKmnwink
XuaM+JaN1WweL9kBKda1+E7DY1IILXJgwcQGkucFJaN/4Eq7WrjfPNGV6Qxl8FWHeo763sWVwwH9
pzOYLYZO/B/pOy6p1RgcptpK1C6eHlSm5sPAwpZiOKGZwFtdVK/I9jD0qNdSy7OXUFVSxeXXJZV6
AX/QPpb3Iv/J2C3T3rnNHjsIlzGLDs965TlIdtkyqQGX/rBH/cL9MSeYAoDWzbJuTHAXNICgDCC+
BVoL+4bNWTMakElhylV44QQn6QHy6X3Hj5egXAi2zdytW+jKAMsnHtgy/BtRYK42gqxQ33PDoovP
PeU4ysDWiU0Ig8NL1xhAc/qsU7kuLQ/gl4tOPrroej2205zn5+fQyRgkidRSbctbRpjwb/MYy1+k
yEIzFTlx4e+vrrb7s8lXZKybwg2waNwn8gqD5GoD3dTAf0t0Ob7EmtdnO9y83+6yFbJ10ceb+zm5
QRIVlF0yfElJMkL1KJqobYK0RSkkIgiExs8ewKc4Fy3xD1yjAlWjdPd1WeQX7j9Tk51rG3XlAzuX
XgeZ1J4tWuBTHkVrZXW4SmKYCjHftS4I+iiXihg2yulFStNOwZSCT59T1QE3CdgZ6lgF1ZnDK0us
HheflUQDxKxtHOviZct2Eo2pw3iVDPm67LZCgzxMz7b9N+yLKrU2VjUXHlpcv22Ki7lVRs1pHjiy
GVPobr0i1LWX9x10SMRwrlKgrF4Veb2lOuL4Gb2y2zVGB5lY9RkFGbbEz0TsyWfqKmUI7+ztM19W
YgkMCi/a8H0GvXzoqokkANiIcdd1G+T6MIlyarUq9mZITRcjkcSafsYkqE7Cs9ec3tGBNcpiVh/0
tC2rB1XGkou8c/eJ7p6GMCKj6Fthi1uwCRo9bTLUpdkeIORtia/sKStn1LdjIedY46B68/pRAixr
jSQ6KhgaiB3yEDMOLO3qLAfyXaCeSapXbHwqpKQbhNHSRalY7i93OM9gXXsO0/YjqrAFaZFVryLH
D84mtKyS4sAjT7RyiwQJazoIJYrxzyx+tFXuxD2dXhlWrk+/c3Cu8+3MYcxuN5ymCRMns655KBC7
FMPGl0Sz2QE81rZyOusHbNX0z6GwcKu4kLrPb9zDaZoJnSF5aJTcBDEjyf/0Y5QmeAhO/2rCELuM
vbXp0E191G0HI7dB7FdEVN/+NNuDfPt4BVno68e6jmkYTyEjAFh8kmaqra6ikVvE9/RkJ+vkde61
46ujRvc0nmQsSp5Ub93RqCXdhn2gc+d46+fQgPBtHZ7xfux1uznkwHoXFi+GhqL62JyyF7THU845
7rHYZx0wzZVpE/97YWNEgdj8CkMIPPLEF42N25T4hbNuvi2QWcFNLF+PgLm5WvOtgNoLZoWUG9aP
BrYD3p/EMBA2JNB5vj7YZS0wMLCTdDYUCUT2gfak8k0MdjyOyvcQuRhucRrqApYhU3CX1zxNNQJk
G5JHBly9werEUVm/BTN1iwH8QpbihnOfLf5FlqfKUt60TAWpfPtdGcsmhiwFaGnZXhkXlz5nRGUV
fDN50xPQ7MdeEtvWUsv+WYXdk2mtF7NFTOgtvOYkR+TH8VEXUVAaoi8YeoIPULOzdGdtC0RDzkLw
qGt6Mi6VeK+UcuF1Iyxj8/2xktFLRsA1JymA4FyXqXAZU10d/bLhJwrpEduihGqFPK4Lsi3Ke+FP
WjErwdcO/Srjd8IbqnVreEKjRAXOOpWF+huNM4ioVUE3v4CHIZfrim5XxvddNho3PS+BA6NYO74Z
SoJcQKaw3dUj9SDvzxHkgr3KCvQGvAcCIrmTT5Fv1S0LDlFHqIUACK6pStbHysiaZgx02TadT8hK
p7YKPD7EN+8tNL8ToCcchqj2ri/O+sbEZNagNgun4aZZDKonHkDmKyZ7v2td9Cli4A/rr6C+YZZ0
LBSXzY8rkZ0c9FCx8H/XebjidbvcAn0R8AZo/nnNL6WFmVDBt6hJOoIFNozpdWqLZtw3WZMgIrZm
zIcgc0UH+Yf9KSi/fjs8qv1ZwaOp9Lf8BkYFvIMTIIFqoaqdKf+r7biTOCRKjsxFeE3oSl5sxpMh
Xc2LDx22VEFnJbpZoPi28o8EY8RXVDCgow7rhxXb0nV6nBw8cGD0cY6Y9lA8T9mSZ9yFkNXV4E18
hUkkI+x+VCro9DSKoBubUXV/jebPixwHDOtYtcmukaE0PZxatgQg3mQeF2aZ0su6hkMURIKBQMZc
hqd3Itd2aH0hKS8PRRTk2QGrzXnlMz3IEbt7vlepo7jvSA1zKJ1Z7yE9CMZ5O35pI/lzuHChhmkT
yYfynTvNvs8xa3QWfq7IpFj25woptKl4CijfcJNS684x+hTZGBChJ5cIE9Ygi9R0M3xJ+brsenR8
JUl6CnkTocrBPyR5t2YJMzH6b/S/31m+yXdMN73mGWWXsB+XLuYORDaMeux7ISjVuwWKBE+znv3k
Ey9vNSw90xeSeW0iZ0LwB63ol/jYIZOBGr+FsccE8ZPO+LbI5NAo/pKrKGSasVFZO7MuQZxRgyQO
xYVU86kLglvvC/Vx91qveZf/CMMWkU4mJo96fVcYmXs8IXY2IfzIMkOHRvxzg4LHEXqSk0UOQJ4N
89vKr/SKN8Q4jJPmOP2OMk5by0yfRL+/jPODLijty6fR2prIeB260dafhfXqtTxZey09tnGfDOnU
Fr4O9J8xcshZhjb0Dpwb9PUtWqVkq3CSo5cmxvytTx4i8xeEscl3HE/HyJq44wm884dS0N41fG4v
pK6vuDAUfbcrTFK1kCHTrA9zWttqg670m3eZKenwMEG4L/XIZc6hFMldFRyvQMDMy+aX+c2n0H5S
bhB9IN3AqxHEVdnk3xitPNQpAi0wyqGJNrImRye6m5nfvbkxnHw6dH8H1zcqn1punyylk6k66mOm
AdNBY6K+P1R0GuQfyL14/mYcg1AsFl2Zz4dkhZqM9LjqwU4cRpDalKdiMXNbIWZYkxCbkYvkMqyv
PmPD+TmfHAqwwrSJFG/2lsQt41QvllFhO14DV+7fL7+DrbidzYfXRE5rxRW3MptcpHl90sZDns2o
52EM9ryFEgJCaMZ3FWMzlIF80ffJDDpWK6GYLS6dd3kGN9g6dL5Fg3GUvTiqAnCgVD4Rq7hAvR13
FRd5V0okeN87CBzjU8C/G+NCAYcySCF+lMjiA76sofIc1xWKVxK9glzUSdORz9xqLwgYBAGoUvo8
GEey3DW+repVzxozzABX2aJp4YQoULAKHacHMXM3LFAX6hA8RQi+xNgFq7++OhYnkLd6v1uJ3x+L
qksznTsb/rlseL+iVOcFT6i5guFsPpAxbPAC9y02p0MFFbPbgmdDNe4xwUOMpq2U+5G2pMvJ5ssV
KfbgEKjvVrxTbHtzFHH5K5sXb+ogeTX332CmIt/e2NsegrVdG8P0HYKOgkXm6T7L5p5DHd8EWVh8
BaUbxwsMvjb59tkw2g1VHbPn73GT4T8tio4Y4jlnlwEuvd/QUHRnrv0OQRe61An5+XgurHJzei6g
1DqBJnpkKi2TdqJcncpBkYPJ/ufHRSBg1B682/H+ffCt5L+TJni+zU8BfGqoNLc/LKrZigvT5Cfl
Nfkv5nhp6CWGAWosD1vCk4CaTI2D/Ww5YW1KyMRUnD6yIDdiSduC9ycdLQSsxu3JWjLRURAijbjp
Gcynh5iKyPhUPaAJnW17AE3KsVjdCCw/93YLgRoGykTJVd6qlSDTT54aEYANIcVVI1L79a8yjpV3
jHa3+tSxR2M8i28oSRaB2flnQNsY9cjhN4j4QIQl1EEigC5GcVHpELyWafuX8oh3JwnMbzCcMK1z
iB5FFaKYTjQy4Fl3F9flBFDQztBrQDUviq+gDY/Gpf3twbPtGsJU0aRuHBuun8ZmKqe7cofyaFUb
2JvPnwWxuQeFXa1OFzoaFFB1wq7pd7jKIMGKujxcK4CaYpd6/pdunFzjW2LCaGJ8wp/y3CZ/OXrU
K+CRnk1I5opoUWlZV5qxxwjrIdmGAwNS5Svm0/t3qnqnGiq9QEQLpJoPGqHwqP12VstSO6LT66Hu
9w7gRmuigDrwPl1FqlNHico2RGnZzGt5KFo8IGSiPo5a2EDcC2y5OWBErVsEXBGTZsmwMT9vRAZA
Co0Nw6/miDKADw/WVt3dHAsT1TLRYAH9Ah3DCfWWWoCeZrG8DU3RFl/ezHelv/VnaP2ESftTp92u
1Uqw1NpjY1/LpndpUsjd5BjE5NypyZJTmlABFnoJPMo7ItjgLsheUOKHEcQCVgCcFjYo/Bx0hVMZ
EZ/olKIozljQiHzGvX3Q+3cD/C1KQ7MN4liSSpsUkBHaWPYE5sWkF7RxAD7LtWExlYfHj7xNmG/9
+vr6ONALa5SSKLsmp38ayX0ZAmFrBKeSDdn1ZlCZQOpCafM2M2ubsXjrXROM02PiJo9zCxrBfQeb
kzgKx979gZAMvXyu/ASUPPnt8t8kNQl+6bxS6Y2Q6qZW1UjP+4oR8zNAmncv5mA9X1R/mq4hdNlS
N1LJtkEoShJKassSfHPzyksJ675lIU4mEVOIDpsC4+bM3xpAwFqWhJrl0uqdopiOauiUAxg79ggM
ojYfTXBRjyvEctyd/H9ewbJWd9KqrBuxUe9iDtpuunnkGC1ersy1Ps8KDDeX5uAoUcYOWW7A3Mmx
h3rkWLQJcEvXMFll/MlKNUzsA0CLW6U2kn/aZjr/7yaJ2IjP785IEqs3uGQubua7NE9m7iQfJP9W
GLVj73CeTJkcQ6pMOZWiPpX0B/oQtGop7/GOuoWYUlINPyYQu9w0CxHvP85xkwO7YoSyl9BrHtOj
ieJGFk7pejNzpLmqxE6eXlRcTw/g7B5WE7qaV7vdqsqVk2eNJ3jCGoJ3lCNczrvbGnp+lOOTis6s
wXqqYi27E3eRVgpoiaKh0XiOg62k/Towhaj/2xtW/Tl4dfGM0KrKe21B7dWj+daFOL2tcwGKykSM
vzJtoVz1FGAjOBeWzJB75BnYI/Y4fuFmGgY5bNEXJ3duwS5mV7WjhWdIAbdrP9LZnDtXN02qUyFY
8LDF9rlcuWZVWzLPMUmYZsB2sZDauB7TSCNFltCWtuj5TBYP1Z7T4ebO4Qj1OnVWt6d1B6FsLVDW
c5poSP9gCn8r7f3BXWVQQ2jxrdY99VGhA5cdKUXgfybl57/ftTfA+Tpj7uF2RrRPgI8yfTC5ox9M
ADID9aE3p5j3jPIExZPy7SHZtvpEF7b3ItaPgMdYXFBGqS9N9ZpQTI7VtlVRqUK/T6wkjUI4jRBg
qikc0BUs37mPQFjls+WguOMAdQ2rikQEI3dp9TPhz+/ZoI9/E0fbzdxKM9V5TWrPrro1SAmocff/
0KagRwbHRXzVyX8tj2QSle8QtWw6o3Q6m5eNIYnxxVHcW1Id7rWQamx2mQBaSnTiE3ZxYs4wqLUY
tq2U8mKk54lsNJ0nefP0tPKnQWxx87niyGXAiPZPFeU3rI53FjvEKm+L/KLspMoDClq2ZlKDCqFp
NeP7xPQmyZrVV1bDDQsV6NTvfbWtysK4bVDWt/8UHp94wAgbvzZxmQHCGO1U+0VQnCpQJzkk9i+R
Dab++yYw+Zz9DVqCw1oU5NQ+3j0HCyZumxntvmhInvn6w/6x2qjQSxpsO/Psm7HyCDmSqUW3wumE
yPYh/OTHzfWTswvfUgdThm7NgvSJQE2Uu/3vs+TaOuh19P7a/nfSJshM/TBZ4sUnjICAWxgr7gDV
NbhrzPGe0zS6pv6U5Um05l1p7fOAW8ia5y9MHHa4HpncVGOuawQG47wfnYnl3l4OjYz1EgCx19Mx
bickyflTHwLI8QqNGw0C+IoUuC9TyEfz4VMU7Ng1TmduYgC96bL8zqiFZOmQlZDCndCwo417/awT
lquV6Zl3kU+1FEXdbbJPR4I5FpzLkv1YxtHsQ80TlkV91LPVYClOpvHeZ0HiNQWlNZ5I3HMHzL5A
AjmENRfFDKd3DdJxz9/Xxf3B9dVLANZRsN8+bE16UkDgqE/36Jj/uGeLmmzHtRoql0UOX41cUgSM
UW0E5v6gHQxbZigfsCx5osmY2fKRkVGT8ENwR+ZIrJ5Jc5NOV5oNUJItc/lCWXYwL1rF2Hje7ZkR
2i13xq1B+rikl+AIAzZLTeVH3UjMDy5JTf7VByPwxSHQ8FAF/qACB2SB3vBqMJXyb/3rt4iL1MNa
0LwO1CqnueeIj377AWjc5KreA8XoQ9tZg6ru9Mq2mDA3giqSFXdKx/L/QVoksgzEkYhzGDPIzHvK
fwKwe8wOH4YMltIMH3k/DWrbuu/d2kGobyXhB9CmiE86s3tjpK4AhHeM2tXqfmmUhFrGmCRasL4B
hQ9mUQlV+7ZEAmwwz91BYJu9ldcXnCo6NMsocQEdn/TboeSesCRB0soIYVC40EIDFTK+n8Gg3o1D
6ih6Re5DJHgMnbhiOstg4nT5V8McfpF4fxAkqaDK8uVbrMArWq2AP1XZDmYsHPK72/eSAfpjZwnr
TYcuNS/jN9qGZBniuj3T7L+Zp7f1ZYtNpIZRsh1ldB9oLf1BjzXYwgoBekI2bgKv3M8c+y7KfMGp
4UiHxMoIYLu46NRPAGURjPefKV2Kd+OUAMTezeuEwlvN1FiaiX8IQvD56wDM3klGvdy912ntCpzN
eKVCGmzoRh0xztXLhMnq33LgyC4NAMgwYdlS7zCdwO6ahP4REamsqR2QxCTgCS8kjQ42AJjWlDZr
uTa+rL+cncohjSpRIPmJWF+DWtxb2waGD2nmcDVsdli680LJ2dw3fri/b+c26sSnhskdLDvu94Rw
3q9thPj3rb0Qj1NQfSuThHWrFknQaRbOBPilXA4O5HEbQjukA9qYSRHCdAwXCLyFEe1q2IfuC+qD
u1xNYXcbfHJYQNYWqTsy9Ql0xR2HXEhNkZJMkvzOAW/VXskaceQa+qN5fbPfsVvl4Ux+s9GMK3Z1
KtI2XYhWAhAJFqbDScgskjmf0129hwSGdWZ8tozLTSCpURvOhVRGd3+JwzEEJCdaJZZY0TaCQU13
1UQ4t4kRyjHUyNsJarwmPj/tVGZELqgk4hygGzcNYlIAz6jzsDhFgn8/tu5so9TSd36dqCqx699P
INH3PM8gsRtjYnbmFlXR9Uzaw3Ued62PnLoAdsZ49iuvoeWgx+tDIPUUUKsiSv6IzQkKZjAdPH6Q
KmUaElbvD4ViBk1ilWXDXjnGbgvTpZrzn7E2z9Jbo32KSPpPZwlB5c3o+WwBlbDY9tRJVgYAMZUY
S7iBUqA3M6ZT8CRDtzVfrUYPtLX111dBE8Xsg1I6+MC89vHXqRFgCFXGMIPKWWmJyE6csLG2rMQ/
bEYDElW+3kDCZ477JQni+sTaI9/BveP7dHf4fewmLovr+xRuRbal0VcAKsv+2J98jE3xnpj7ucAA
Yp2+UflZc6pHaj0EfHkRWsphrx86p9NhesFmG7y7Tv8VaINMh/QieecRyb8Op8QMj1F9FAs1BErq
QgSbk7t9N1yXYqKgZF40AnKtXDWA3PVWmXUASoobsIVZrWAYOYIp1b5qwWuAuMXmp9Ny67HSlBCz
YYVkpGJw+gkZECPU8gYLHqyuVlPsgweNkVJrGN9re42Olm/OK+MIpkCe0eIU5U15ERHfMp6IvybH
T+x4MH7nQW9BkfelZ/s4sh2zlOT772Zm8HDe/5K5I7S+TSkpAHBwvdDsOeJ9CHi7WjqhDXqsikuV
YXWQ0ljkFQv63sCjyzGy34UetLkhgq3EwFjx9I7Wg/ErllaBssFPhiwxmDL0jO3Zpw1dVE7AT0Kg
JUX2Um9LrCW1Ny34qt9QYurCdLluAFdnn89hBFgkMN0fotN42ak+cM2MH4qGXfrIKAQgk9F5hNCr
AcPEOj6/2UfjZ43CKGO1pSLaE6701zzWhaD+QK/EKywPFOW3PA/RxqeaIyzF97z9zZlTLeF8JiIx
Z3/DYmG0hPSSoqy9j567uzER3NUBSLJBclTM5dQCj5rgN02rkZQzOA6avvizs+oiPm3EUqEh4LF2
KjQA5C3qYk6iLl0jgB+NQ6ulNlXQup2oVlSX0iqB5PWw62wfOklGrlQMP1JmRNgTuPJOyzuEIqr7
xglp5YuGrkcTLokSm3W/nOgtJAF8gOoc3SPnnScbbHFwXEIq6owKMPnhREjYcRp7jSSZxqdvI06u
E1a/5leiT1YYdbodhmaozSUJPE8axVoXHQ2kh2m09iISYn0YV4/So+1oZIv9R5Y/catnvBV6ITa/
ZKgV9dnAEzxbai0MBHmqGHcYwfasjxANR/7AvXvcm3z9Vh+pPC45Go1Vh4J8EWm+JoKp8pXAJpKW
SEo9Y0gMZnCaufNW7neGwY4nzhw9v6i5BGAFgTL4UhxV8M2euWK9ofZr64GcwgzTtJ73gpJ4vtxZ
w+cLL1LXj09LFkVbVE3dOUuLJe8nyqm8+LkIRu3BzzVD//DonL50SCbiVrZEXcrovuqB7NN9AjJ0
lDWgQ3qXMM0Y0ai2IlR0knAvEjuV65foGmUfL7dCgZoQ0IyuI/u4QqHXz0/j4F2/rGEm1KC0fXFA
kpzokbDGggWnt8kL5zG261jKH/cE+D2NKHmzBwSaHWLJRK2bu9XDlCMwi/PdgRs7Sdejb2aotkpz
fwa7Amnykm0Uu7eEsLGFPxtqCBvcg6t3HRXvv3La57YuknMZBprtPZRCHsxWMWKX35ADATgrwNoE
oRXyenEr1TKsWFP0BL0rEjhsJxaYjvaON7Xxgbq+7zSOkdjuWIdZTZBOPAkSKZ8OFJ88L0MW8qH8
uA9NnVVYFyiZtJc/t0KOXGM0drDpYam4sCwDxy/7cHV3SKxvc8zy8DR+nm4zfOZXM5hyv8q7wY8/
V/lnNPgwjdTm7ZRlFYtFW+YTrb6qBgx7EUbeUdNJzw2uy2MrqEGrIuVCK5Q6KhOQvI3deOv2PnVW
qvzMVssx8w0GMOzgkclluUDct/6KLf1Od50c33iYgFCkSQ06tvMZ9iGceoG5ggoYIutQ6v4Tsm1g
tDtbPAEB8M2jEjlZrzBZdtdxK3cEnF2M+rk0GKG9hmjSb6maUgS2DTgaLj7tDN+shTA2rgjAcPeB
qLl8OTz5Hf82lxZ8khGGGN+yxNHC1oCbTY7XMF+1ZVBL6BVO4Xu5cZvs5CJYra3nuu3y9S2sX4V+
2ZRySo059w3WxkNJyq+5Qz+3rZSFBJZSYXyvI3SEOf6zrt2XIh6uzSXESx6rpPM9d6Vcti3EH70X
lUOH9l2sLOGoNrZcEZKxmTYpxSp8lM6tb7cKEMkD9ZGGKyumXekqTAVTSlrjYdm8EEliPS/Erzmm
mveTpGZFKh/DEd70dYGwRwe3WinQ88kc2wm7ndC/qfqhQKgVq5+jKvsjEJ2n+YgcWS123g7U7oYF
vMJJucFMyjW1KnLh3fNPdrXu2R002+E29WltVKkYjFirRvlRZGzS3fajfylh6glDTXtgzvfWWYzf
Qv+5EXjh2FCMnvmBldLOlLIipYxl8KryIzBMe1MMARxbiKq5SwLnwqRe7F9kaZYwzB8m03CsVyZg
LBKZcOolV/s2fEJdKBUXkE8W/YNILr+a/Yta2pntBXIb24ufeCjHpqFmprc8ysQAnA7S7/CNKTvx
9ivXyO9FzXQpOR0k4aE9Zek+2dFYoenGiypcg4vDqw0Wq0cLOBRTFXgT8lhpagWmjo4l4y7mP3GG
s50AW9XzKBIwVAPaf+ocqdvWolmsXAofdWEclTnuJMDbsGt8x4GlNcroWammVBuMq2gXD3Sphtg1
JM7BXSsQMLNCReMr0cuKKcT/sD8Tw3mnxqIhpD4lQsiLM3qIlx7hMrAKvOZlgbjwjjRD3R3MvrS9
hh3vadaCwuIe05E2+Fsljs07Z4AdA/ynmCPNDhRPsdFj0BPcAzmAUZoM58c7wRLv25uOUPSUoR8X
nHNIhVYAS6/DXJkEuOC7VWxOUxPtVxaCXv7IyT1XU8jnu8LeYDDh8X29Q2OWn7rqOB18j+w+/eQz
/ygy8nbWzsUXT0tEa7/fs7eQD84QkJSrcUfwAyA4UgJu1Me7phxo63F5ahUpcmfl/eO1UjebA5ah
IPBKLB7nSVkv0Vk/61LLk+OJT9DLgjWMjUj12b7GJXKDhCKj/DV71zPe8NY9gyWjaTOTXXyWINUE
TZSG9b5o3eTIGHqNEXkAVkx7YJTy93zHUSoW8kpQLzZ/WaMlT16BbYXPIpWgZPl3v0TzjmtCQzSB
7jdxulpM9zWHEY8fHF6w+MlLl7Kt8wjOZsisSAPYlVUurppX9pCerqFHqXe+H/WUd2dAUPinyDhK
wDlijq2GrzmYBA0B/om+jFiPgc5/1pCE5OPbJZjqaENkwje6oDQ8C/P5FnVbuVBN+MHY5C6LXLGZ
fhaAaYbSer1JZzZqzwZxusqj7ih/nCCsvk0X7CyGxyMujE9vNz0THKbwlaPTE/G5MUtIj2zq3QL1
+vZCCv6+JuTWMY6g6eYlfELmjUJe9BFlSh0/xNsH8R8AfmIkdYaJiSF9/H58lpziMeS35BUH+BDV
6LH8I/sjHxP8UBH4fUAPNPEWqWwkDyl8W60wDSHEP3h+cF+AbOF677wy4EQ8iKb9SAIIjLKyAwHP
AiUbH4RKgnbxdX1cVi5qDO6j8k+V6zP3QxGCIw7kSdsdgir5NjWG8mNto/asDarXiQbyn+uShAL6
9MBdGa/kFgh9S/tDHweciqJSco5McZxfus+qYPkM7Jmmj7S2xP5IL210o1NZZIi02IHvU+Uf0RU/
i0IKfwprp27JkN1NsEfJ+O7GqGd9LMm4BKRWtW6xpe8wMM0NvikdwSEfkJESi0g0s4VCLe1ACqgN
nSbRRKQs4VuS3VSlnmga7ao6vmNOhojUkEINaw5XbXCk1Yf3iuW+4CTcfio/49dWJ3Ayg95GH1qX
r83r/xHh1iGfJGWWqrMRAiOnA0RxJIwfrG9EViT1XmFgUJx0gBYj39LsXffJn/YKrN3EKbCuNHu5
tFFeZSljap9pcKlmTOcoCg7gWdl8BNrvHCih7mR7SYy9osZGxKtgl8FlHJpS3El4ZGg3bLU/5JrH
bmX9uv7ytxpoE4kjSZj5l8Xxt/QLd6az4v0Pv96uuxM6pt2ElCgaN9Em07eN979BVxTNlSSOATsV
5N3RJH/p/Hnz92vZC3pSeIghjY0kt7VSbUh5I0GeE4bM4UWJIvOMgVdP5Dr6PqbldNA8YLkVhzui
ex3vTJ51rz3j8BAfDdpvRur0qvtFqRjDb0S+VViylcuYesBgNfJMLrqR3+UIgGrQ11j2ch1F4APU
Tiec4MLPrgDZkzWIi1D3sHhPtuikWmXz37dOxZ9B58MSDmysK6YOx1SkVAstjUcbIWGVwGwgJMOz
S3LqPgbDQSrIMhQfOeAUhL2oZMCHcVTZLCyXLqIfHsGDKsB0ZdgJBdnii0WkZ6qdjL4urhD+b7ig
PF+qs2L/lil3YT74hsbND6tk9l1q7WRjog2Q+lp9cRoys1PFZm312ZRAwNAu/5ao92OfKDiZjBPh
FTi5B1Tyyc+SHDnowJUsuyazkpKmtlDlNuwX6zHS7IWDqf1ppP45FE2auwtzj00Z4P+yzoEDmqXT
laZ/mVRAj6RG8uYWIl33YrE4igPUz0upIkN0ehVsb1nLFmucwCd63RRqFyNZ6NeQ70h6WvCRq6Jz
OBF7LPaNlWkSISEnapITEkvjlr49WJSTJ2wTpXDaZsFd8KSnrHnRVbnZWyqQ9be5U38Hn5cK1Ppo
bWJBJToc2HDb9phb9Tjn220zNHE1SoGA6x6JAbl+wGQk3RhIp1ogSZn+8DPesZTtL8sktlebkjI3
OvlAExp1Ynb7hG1ewFz+s6bFab+JByc51/GIADkN4n6nutIPbaswNiKvzWbRyvedptIpDL4S3/Z9
7syo9PA2ytTHx6HB7RrH4H9SKf/kDBsMsuHmAqxEarjreUZKSrkoZuJ//LbnfTwyFUATQscA5HGO
+F03Edzud2IWHcOaV1JdwWTCWscTKEv7itR69vQFcy/I/qezl+nBa9tWrYVSM0IyrwuOY1skaiNd
T2d6rcs6o/6hHz90JJEC52awcJOgWRrkntsLoGI3ivtYQIPEZVfXMEIxeLeGYOmFovdpgnq1+QyM
BdWJ31s0U9TNLXdfe+9sqdlczIuZzGub6sSRn6EAHmNxBbzS3aCnaPx3M6h2j1DejpE3a5Va3wo4
3V1jlW9s+ytzUusITiJZX0aGvcqPdJYJ8AGXR3KvASlDyXpzuSpS37u3QiKAiLTifHWBtwVsdMsu
/4JMH1x7w0pOb5B8BrQw5pSMITrUZnIPVSPFs75qu/vbH1KUqfAVdN7dLHF/mP/u6xtO9XhqmIpM
S5BTAIDC3AFEBv61VlExSxQvo5MoS2ssEusVASWG8qjMmEEhb9JjZ0G8YxACD43xK9JxPFadvRuJ
Szw8q8yshBuwR+qCQnbCOeEG2yAS1fcey4hp1nicKCziEehK54NX2UJCm0l/r46SZ+57o3Fzh6eG
MLV59YHA27KDO6jVs4ove5VuO4cYJMa7jMr0Z4fpxe6Ue3eSnbqrgJ0uFBEFlGjbzmw2DrtEvBmt
8vxj3rSJruxOYt/yGsRKoR3dlPzoB+C+2QNJ0CXmpsU8E2Nc3D2nlgOi5DBuV9ZH0yBH03qfnSgg
irV6CsuGylEBH6O1tf4W+nQmYYXpKvfYWhW+Cn14Lv42l4w9hhPKPsKSjSqzrP/APhDkgLgWN5a/
q9XuckM/1rWy5MVNiLtz23m7vFEwegEDzOYJYHwUj9mvluvS1zGmfGaJKPs7JoyU8nymYwoE4Gj5
WMlxIlhxqvbsrbUhO1ele3xdIHeXmj3N1NdEawEc/4vH1T5T0uQWCgheBKN97/O4x5/TEQATCwY9
stPyiZirtd3Pd/gR0ujalklYolclLWHnNIOBliPlpT6ulv3v386UR0+b0vBhMYuBf3WgKHvbErmz
HQEGLnmbrxhnCRhk4xL9ZuEl8m1j2fipG46F5G5kj2rRLGbnP9W3dtjA5kDFfeiFWsu2rWcGvORG
b71gVIbQCdPhO2j/oR+HbcXVDn5OnUokv8FxHDgusQmhUkVTAZAPJ6yFV1jSp1b5HhHkqSw78Fmj
SX65+5pKneMmpBSLlPRKlf53+HQJNqpPRavb93CGg5CabMvJsFP9bekC3s9k6OEF7Akh+2bPfoLk
Z/CGcamXJL5OMSkwhtm49cCUW/uC02BsveUjjqoMhKGi3BiHRbDTeVwaZTGy1nnQMKyEYwOMHwPQ
kS3jQUatPNprbg5ckIx6UmTZzNtA8dvYjkLoi57WVEqPO02vMECtKDCnxIfnkmoEJHitbAIysSgW
6dkR4LTiHGtlyBayNuePsVC2wDOEr+Ms5umM/psMnArKkNXRsurMfI3KuTqrB5EW/UzuA5yU6R15
zx4CvyFfANl9TEzPaaX7mtBEHuCCGSFTapbW8ahtcaAq+VZINKPsBclrvtsAQyo/Ub1DX6Td3Mh8
Bcj7CNWdRstoKrf0EbCUqSD4wt4kLZvL/QkINzX8F8OZCSD2tE8847ctRWDpewYmRpgp+l+n/yJs
NKeEu7mUgzfHGeM9HGxVGBksrnIKYetQn+eJzP4WpyMbQ5tTnIUhr7T9wcwiINrbwWR4GWW4Nm39
y86cycNapkA1h26kw1s0LiKOwMinldMPUeJ7A+hk3oEyzjXhtsGTSfwr4GJdnroN61WdH0TlP0yo
aUft+OSfmTQ04CcsN3ZiaYYWH8HtxrQw3ViA/BiCT3H5NVnXrLiRZq1ZkA8Cqm7gZ614PW9W4lqV
kgNW9suq7iyAFEtMmkRDO2hP/xa9cYOVKwj0jP+lneG2xiKTpgbjs2xoX6kxJsGqBerHixn/3DC+
0Zzt1MtrFhtO9s6SU8JRYVJJmJMH5zQeY6F8m+ZBLr4d8x/cIlsPCdMMh0HBSIhiWYM92/UFYNXS
hQzHxlt0+R+ZlIAjemN3vvhUgkuwugynSplueq7PA/wVnsVAVdM6OQVCKfERLjH6PAIj1OhKcO+c
dlYIA298Bie9UhzfQC4bll4MvRwhVCiIsxmZ9tGHdYo47u6GquaqHASdYkUgvY/SST8bZPWrJa9p
uCd6DNzLMeuzrs/LzlPyp66VNYmoY05VvZz9xghqcvXEA0LkQ44juZIHG7NTtmeYbVRgCLJSd/h2
+ieMRT0dtQzj9SBKdWwHiG5HACd9op1Ho4+p5BEvRvk4qPyHN6bdiTiB3OkTl7q/qUhdp1ji1s7/
LCW8MvWc+dDpzjPUoIQYjkiuoq6GVjkPkIKPezYfvtpWDTmmRUlzTxSEu6B1/pL82Xvokpj9RnZZ
x7X6oiz8kbmrpME5vjcHCXzDwEcNFbCKpqTr5RA5IRD4TnuHt3awrlKy+CijQitFmL8J7U3exuyL
KvBbjT0NkPl4D/7GcuwcbPSTReZDvU0AaKqSdNkcLrWligzP0t+K959+6dQZe8y82BZlZZc41ssB
3VJiouaRu55BYtLVSTiJDi/D3dkHzF/w31LoEQ8+Ug8lR169bWBykWNAYHCTKxQODxZc70O9/UlE
DLpoJgy3l9QH4wd6dnrtutGyVzZIxAyEwgRW/+s7tRlkw4XaMcCQB5cVxUm5NFmwS3i0nYKETnc+
Ll5H7NywFtpYcxIEPSJvyzqZzAQOOgEkr5RDBzjfT4qQo+Kxg0ltynuhMpepT2BlOUIdO1l2c7yU
0Fzjtsz56uiM0Bf6VoKIKOWxmtR75qvCZOXJcDdNnaMJED0vALWk2CJ55adp5HhqYdiQ2eGUeT6p
xL15C+ywHP5L73lvfzeMk4ky2dRfIo33mG1XFnxRfxtnFVzwFwVSWiTB+F7uQtSEYVMbJXLBlEx/
SZMQb1hz0GtfFyVbRTsPeTUk+/XaiCsri8TU4O1geMZWvsNM5/bD8m8yMPNyeZKpcm3V4hd8+fyZ
VE9KOLj/Eo80Da+/GvLZ1+OvqdaQ5v9BbdGxOP4y2Gei0t/pCI9qRNum95EDqiTaKIC1Yy4YSBYu
2zp5+274dxW3J7saL4xw7GTgmv+L2AMgWW5495L7ypfXP/44PtESz78uWQGISuFg1BDUlylYgvSl
jipjCXh0xjIvDbqJFqveo4Kv5UAYDX/WqqKYm5AxjH4sb/g8YR9ipVzxfSwaQjGRYEKZrjWpVW76
y1Ulfmvc2/yxdAl4hZQm8bIj52nD95LxAolLW/1A8PL5BBpf6bvumKaDo5Ff2l++vm2INU3Sao5W
+53UdaWWSsy2I+krk+emef6SAJbaW7EjA75AqgrTYJGEfbJTIQ/1EgWzRWqom4Ip/A1v3q7sCYKR
qAMU1kvH9otcwUx6Tp8EKaOmcFhxHYuIzzBRI1JkoBCENCXlWzVemqkF1xvjW10bg5xRKJq/Bnvy
V6tvlHPQxiQVskAuD/nUAnCWWMJT0j7eJs84bVY2pXsUaMzVLq/iY84JpAH1B6LYhJrXnKdLJ1rj
tRWrpg/jxeS/9X4Ooi+9g93/c64T/h/oxRDCl1Ck3t3GV+6guTlg6QW+lV+SgULZinIz7NqcpUw1
V1min4sG4X+lEVwzagJdG1J2LywpYVbKnJR9NcBbxleqmz3OgLyw1YQ7V0Ji+1InSQOUMcxMuAc7
m9oByK+zNejCoP0zhPzrEIECg/2muCV4niN9NQisONCJBA36M1BXqKx9Mn42ESNw9HYIk/2jhjdt
sMK1KVowAf+KPUXWIG1mwR6dbb+CQWdHcuwEvdwvCHyiOKkggygq6Eipp6tlguF6vvV0TrPd/VtH
brZW975hGIaliYKGuscIPnVr546RfZW42z00nQpxaNkeqNA+F/AdVUF0WxZIl45g5XNTYTK+CSBe
937GU4KHSWvaaO5SSBA8oUnpVl5F6pyTxs8Xn2Ru4e0d2Y+rsUypE/NZJwqX911i70dS6Hw6BcIN
gHuKiDYo4KHpd2uthdcA+Q7Z/ZBtmeQtr+vIdb71K/Upk3yn/1KEvlc0S7adD25f4ubhyZDhTji8
QPUfzOJxqGyBVTlQdwhFLA/vZ0fCOIvogPcEOZ1RCRlyRSPjBXVw1Focw/lsNCzXxeaPOiwCmM/u
ut7DmfZ2rTDRSqyRG5DfL/wQ7nEcjTAvyTLvaCrhsvTMX5DH5EjfW+pbG+qYbU/9HYJ0QQER69QM
3dMjlap0kTM4mXfMdfXGQPo3eehdPPm5iex2rKQ8QjEvDJinzRCw6Y3evaBkJVyWA/1SDnpOz0Lz
ON2/nsvKOnW3JE36p7KhmMR8UQZYnZtL8roUD7uTU+fs5SlAbxGqr47YYzrnaMEE8FZVRVsE4Pwk
8ibFkJxKsGt7ViEzWiLxIRALgjqx71LwmqQGO84ngKZ/t/UYOJmSf0KzO9ump8/eM4/d1mWUf5GX
oG+nGo3rjdKGbOG7NskYb+dMRBZz1XWYgZSbl55eCpCCJRxFhvnQ82oICKaXYGciexVr2aVxZOvf
vsMl3tSUThH4olVdU1XIaUJYFFZbUHV6BjQUfJuJk2+NglwvLwxuDwo9NnbXYXFKQWNMKdKb2R9g
H7thjRUCGIh/e/GgCRDHY5mU9pAN4pUfB9cttfR5wT05LP8intg4k7ioh2gWtaoGHDmTY6XPy2Ox
IZGZqdzyHKZUEu1lhvn1EBChP19vQa+a4qUP3cI1slvTZfULuNMLtlONEmWVzzl2wwoZK8o/Nmzs
wl/WkDIolWXhdlZrWkU/aOSwl/m7wI2+gcYZMubRE2yp0UH8cRymysYBEOJJjaQgP1KabAuF1gkv
xnC8+FcwejaRY0qO1jOJNQlV3R6dqfMCoBeM0XyT1jc/EIjxb7EtB2syCKJS9YaEHu9y9zK/QxT7
4p2CRg91SdC27xoQGeFWlRldux2wf0VO70Yr40SdXmU0icKSLkknE327HMkXBYXwLLxMg3ii/vuu
tYZ8MXU7xy847SurwP7GPuxzsxaVC2fPTqC17oaw0ZfjVYPMJ+GXJMDc7b95cclSrOCPlbSjWY0e
TlcXIVXCy5Aw88m7hf54xvn21/s7fPefzn8HTukT5Yut2Tg2nfBBBTfVkmGFwSXi7lZJE2wp8NPz
plS7gN4mpRaObK54PuFwv98UddN6cGFRQWrQqgUSvIYSV9UxqdSO1qvhXMjr3avm0rls+a91Xy4M
jZTTDBsPrUc5k7h+34PrZT0/6KPwikp+wTBYKfHQobxQTH5rMCooRz2mF5AY5IKdjMKOq5ixVaCe
JLGDdigR0J8UZF9o/dtsJcD/lu3kMHoqFpPt3V/AvRswLqNIoyN9Z2KvPyFYBGBq+fADEHbS13pT
IdyPHE5wVuEeYYAiD+NKwv8LtmOsIKYh8+Ry+zYQfNAdIlbZ8mEEoWhqYrY4noJqb6MxKPgdJ5vz
8zZXMOgbG+SW9pKPofKHlq7ONretppn18BNkBaaH9XxHcL/wKwRYyOfIi4JPXImw5mf44k5qrkLR
uZZ+b26aLvQzY2IXUgL20Ms4EoHPio9LWzMEX9aUaplF1eH7QXS3/U+5lf5oQ+uBVFyj4kNC5cZ8
0hq2FRQnszs6ofGRd/Lh9O8LOOaSHz81F7FVkLBaf/SXpvgV2jwDKzldrHYQRSIPLdB6vUMswfeO
bX+ROGsdtOP/xvVJgCWDPraqskKO9Ymj8YyIntCKxm+EN78gT0lorT7k3fwXBQo23OTj6Mj/ZFe8
2NF0Y6rmFt0u1XhRwWWXAtuEwQTFisqO417rxI0fe4rT3RwNSh/neDepwqa084xGsGoVUoTM8v/D
zkdypYme3VoGQWOFbCVcMDzPoaXnXxd/BTXdhverCMEmtwpmUyhctrmDg9kj2k7U/icY7pp9hVHz
OOwprh+jQZT7R7S4xjAjS8PEqq3KgFCCYXKiVA3CO+O7L1LmJhNcX4bESOJ7vryzRnlIn1kmVUJV
0r2whD3P+QQVseNuQUKaiamuXBdOGZ+7pDz+DG99rAOStYq2h8umReeY4+EWSvYT39cdlGNnkVQs
0SqHdP5I/zE3TXGQTohXMUm2A0i4uOX4ogdXJMj9WF0tzENoVQLVLn3O66jsurgMLJSSJyPUKWY+
fRDCEaDjomP/gI3ODDAN8TzJv3BrVIz4Jj0zHSO+lWPT4FIeuLv8OFkKhp5SEIPUZS7LZSLrHduW
uQs7uT2QwBOQD4OQu0eQZcqJkeecmm9hWoSjdAhEzimh10gray3qIWxoadPb81nKkPWFHx77MT+j
MT+dBIZq6Lnsy+bZ7MQc0/DVNP2K7YimfH3DXeN1SVYb+9qT+rl8/CGcsZfGt8juqm9J/Kd1XBJ4
Y+VYMwjdGMG9jLUWHCiZbzvFqpC5TXxpuc87C4pgZVhJIztk64RQChVIMxyUqWd2d/dy5S5lr5Wy
oSbWbz4DRJqlPkMnCx+vTZOUr+bpI/Lk9BpzrXnfGaA5RIgb5rBX6+cR1aIK7Y7oBQu5mNfZ+pQy
VoF0S/cnkYovlF/G7h3Bs8QqREkp77Em9UYkOerWt2j0NbSfNpo/dlw8G2IUxTu8YwLHAy6K5uPf
JPCnwNk2UZMimqboMK3Kq4W+tqhw5d+I1uxcXCuugtBRWMnE4vhTG7S0eomTJ6SIpiN+UYxJFc4V
JvrXZ0pgd/IiNZCyCFv5cinT7OfTHmU2BZH7MCD4t/pRW2a3ANqzHDsXhX4pePKymMQF2crjYOJv
EUDeRMDdG7hWcAlAJR25m+MSm0iwCRdYjp+g+fSzXscTo0mhucWAJgUxGJ+PYOWvwSJYfmDCKvxR
8I/UQxAj4gBpRXphGqPIbq7sYKHJELag7VAmlZvGNYiO2dPB8iVXIzV7ZrUfPsMye1Y7Fyit6TuE
Vdshr4LWI9jvejKhEAvH6fLt8n6TIDHUKOoUwFzOXlFVLZDr8pMvAAUvoVkErfE79vvVvF/87p/c
T9u572AmKJUxhkYu3H2Oj6GClqdA24/xOchBQvJJZukoC4v6pao2MyFvuPCI3HTk3FghQLvbTvr7
rwacpDYL+L5IrCa41FFtwlcGtkzrhXhRph94h02/ST3t5WPDL7qmzVo5lNse4Bk2uyHBn0+W1IDn
f0vNl400CeKG0IlTaHMeXh10Fw6yHjZBDtlBN8xTOUALB2f7vwVh5J/AtMRZ5X3ybzd6p0Qk8rSu
KTAfqRD6Xsx9DCx/2sj5AHGegsl3WVQCSU+K7XMBZq7HqS0WuGy6sLdjqsTN3es+0lCrjAH3PVYQ
cDxyHB1hw6CG8jier8IU98ykZVV3d/JWnQhw7O2yeNSWV3axpaacBfbOfHytJinNrRzG7ltF/0qz
090/hB4TDYcQla7zcYPcX5OMiFufVuZFcL3qEsJr1DdtFx64hhi8SPeWkye0+5qOijVKNsM60LE8
24IPGXkDJhnLDaXG2yGQQIXiIG2qzTpK1HvUlDZ1TlEd4VlJIXLUU3S36O7MwCnswPOYoX9FrPn3
4YQ1WnG4Ejjib3KOYEhOJu2DdRqvrfUqBn8phEus0cbrphxBLSqiNp2wMIX6+y+nO8R8JcDv8U0n
b0ItCZ1kf03bjk7h8xt5Xdstz67O9pYtZVIf7vQrHSmOpVP8dL6i8yava1/Yh/yZJk8cesc9xgV1
K+8IusuIDyqV/DzzjEV/qQGa+jDFruGMKEEMLPw6W5QThIgvNu8Kv6APIzEGk/0zbhnw5LWL93ZD
VWUWraZrvrkeIyzjP88405Qe/nNh1QtUvPVrmFg0Z3VtlIEZuSisUxm096VJ3W36DD1Dn+87NqeH
YXdgTR4yHUn4Ts6MfNKMl0lN4k5yMYq886dAbLoaN1BUUEF0zAPmc09oqbgcbEUYap9iZgG9mav3
mTLUj3TJfHpdU5XHlNO2Wx9WziuZxxPjt5w7Vh404ltx+o5GYLcRjdH4y2VnQ3FROFFqYdjlP53O
pru9y/UcTeIHYddpeEi0NnqdeVLEyPxJj0fqg6XhVfMtYVmv5hYQN/UqrbgeqfIei5Fw28N3YwhC
R+78p9iv2gE8Z24cEaYe5BHkr1qQ7qL1vP6P3de46BQqN+0xBG62yVKOEDLm/T1fDhPCeD0NN1yu
v/bl172kfzNn6KaW1veZqi6w5Kr1xbhnuNFa8D42tr+9TzscMz1rKZ/rRJoR4EepqZXN8hnDYzrY
h3cYdDzvViCcjrTDuT2s1Kjt6ii9Mm3W/4a8XDPaPIy+cKlLD9L6Y0R2r0AIcs+5na+dZz2Q22Qh
qSWKLtbRI5r6Wx48RMFoLga1b3/SygNbspN9Ror08jB9SlKsbiurMadGFwpSXd5YQxaNkLbBMup1
TyFKcaKFqX3Gj/zn9V32XeQoVDBU0++oWXwnwHzMV4AKAAyJ8YyGu9VgYsvk48epHYrs46w5isX6
2OpfGr5khomFpSP9eAKEBVF3P49gSXPnjJUQQIdYaz0qozw3a/LAovlm/C34udgGB/DxxkBwnrAF
rlioQdG9qZud2dnosBPnx7gA545TLK2vj6dZC6gDc2r5QWDoCnhzzMxTm2weNUF3UhYGABGCQKba
fdtD3HZeN/G4nmkAtCL0Z9XDyupRIFVlzxuKTEFOwRgAlD1P1srWib5Cu7s9nGwYYctbBThpI6Qg
OhF2EHi0+U31ptSb4O/QtyVVPRTwWK+qRgEcvymBgnhDSVJwc5tw7E703rtw3wEg8T7GajuimVvS
6SVH7eeQqPS3bHPhMjfRSiKu378n79wNGllKecQfNzPrndLeHMjBrw5YIjkFNRn0sYYRxRlKNcUv
00vE+ktXEQM5/HF/FBMKG27tS31YBVn/9CXuUgiq2m1b+HyR16p/PsE8y8ziTvUIyFOMsGxk7GtL
emY5cMH4wthrZQ8tdMBAXomTwsKvRhf6Sr6rE9E7aZHr0hw6JbO4R3rAKfga71SWrespxq8hZ4WC
+QpDxJT0HTdlF3VyCnKc06HcaEa5UTIVD61TCukw7nO0OZErv5rDvsHgbCy/ixNd4qBdJerbf60T
L36//xexAb5RZIihqhuKTJA/UnP+hFmGYUpMn4nQVaBQYRoY6PjNTVIGjTLo6WvY16mp0HqJprz8
671i1LsGiDATvIm0+rAogTkC+kzd6wZzHzfn5ApHdzQiK+jLnq0E7SZ31TiR05rGiB1Ob+h3Zf2Z
Hz8vCjjTiIw9CkCzGHwNSwc4xrrV4cjAPW7OfXff2ZPfHXpf0cKp4aRLJqVGdGGp2YyqW++S9sjv
A/EhA0zjqRq8TI5LWJ9hGR/8bcycVOai5WOvXFihUZnSEEFYEHpXW3RuzGI6ooYWqNKzynCVdt1u
heV4Vtb/S8f61v94r5/TDCBf1+qNsetzgsumevH/ug/H+BATBoyxAgO+EXtkKc1tP5/+r8HD5F6u
mZSwP2TsLAG0+l6UEUD2Mc0DWq2PSPKnjAM+D1YJfajXwB1/PQJNkh772bkPoDNuQRGi57r8wCj3
uQdvnhV8FMRJxvTVrmxkqOeTmo7Pu4JpJL15LIntl11E3x5dTiH97b1SuLKa1tNtH5ZUWnS8Gd4Q
YKYgvaNRZ/6M1UfabAOjSnnOiIMOexzMdORE2EHXOtNc80IocJP4iYD2DOsmz9KPTXD4IXcVgetX
pGV/oUZ9aunNuNLeYU6mHS7+C6qSQs+vw0SDq1+mbPJSR9bmlUHi4QDetsu1JxBy616tkrn2Ck5M
hSDCALEaRfkXVqg4FoVd9SurXWYfTA2GdwIQvYIuZfnPOBAk61mfsXgmehNvx8WeoQ+X8ZB5sYW4
DiB4G/urpCK7bXoMXIk93gKmFF4CeWnGMg1gWs78wQcXpkRFVi6Ts0TBTf5jh9Fw8cCCg0edsaO+
wdWgZwMI5cPwdNAhQmF4b/HbtS2HNl1UKg9jBnRzihGfeGFAer43VowLDuUhCaqvUt6hgNiqlyGb
qdi+ADhP2BwJ7JDXlZSBwJZOufwezLEoQrGKo/xZR/Q7K8ehFpTOkP4b2rDZ0lKSmDEgIOeMSkzH
y1ct3sh8pf81K08OkTP3rZ627zJGXXRzVFxh0Kkng0kQnklBjoojTNOYzTA9+fZyc3z/lAMjVMb1
973GI3w2vKy84aeF0/GUYHKGWz+ghlC3WhldONKeHuqlHFQEltI/7P3hQVGVjs+lnKZ3QV+3peII
IdBan8xQ//VRx7RzO7H5RjXDymwbcx2MQNrugg6T7zfYC+xt7VC+zgQZcr4q4zfZexGXHlBqwFu+
mmxw6dJCs+t7wnnltpggGk2PgXbCwGWLbaxpDeLNiWSBebUXF2OezZ/53QOXKRF21ErG+kK049K+
iV4QfhyZh+4MD3aVvNrSNV2iR5YnZ+n1MC6h0BnRS10mSXwLvhHvkEGZRwl93MLgt1CnGfxwciBy
6hWCEw3scflq6GRvSKfFTl4CTS2XNhY5ZBdb42A9VjKmz4o1Jd40IYzonhoLLIyb79B/9dVSyDh9
t7cRb1B4zA9xoQ/ky3R1J1zcxDt0y7IfC+pv+PqwqvZnBSZ4FU/0+HjCQAM+12/M8aDxA/A4HSeu
nnDC+enLh6a/oz65DAaiz01PdRl0OKfo7A2SLGTZzrUWyB4H6Z3TK7DTIKNuIyWEJurE9cnQUzsl
pNdNWgUOoqvmhSORxzAvQWh7b/G22TavedEC8hdFmkcKe95BHkAOsETdQOO+Gb5fXY53+Ea5/Xkz
gWmxPoK+DxuCmmwLPrbz7AkQlPO/nUvM8w7xGZ995jbwyiFJL7YTl3Om/DokoZeKdqYK4xz8Aaho
1FdFVhLAkE6Fso1nR0ji6iP3/wj1y5k07aVVBhtVWXcIYVe9+2MdvrCYXla3vefOhE3TkrYJq4xd
Xjb//v+WZwyStVV2UbeauAhw3sxEl22KBruwMaFyiGUzmYmwe5g5EgFrGJItrzRFoaR9Jw+TZgoq
DZvVbpHim6t+LRwqtj4cM5JKpwFp8MZ/k2yQNGkxzEccAL99ROz40dihQWzoy2sTo7tuXUMyAyfs
ZqpnK5PMEU+emSV4lEo8yLuYz+kCW5rgFbEkbtaMeOAlCEY523E/IoN7UBnc4DXE24E/rhPynuJ+
HHpSBajj+dxtE87M4K5pUGnRy0G+B2zeD++Absy92aukNd19+auDiRyjk0tX1a+aOlicAvrQbXS0
IW2tdnbHmwd8PTJnDjIU+6ZBTr1kklzG5Pr6W6eu4lJIByo8mxKAs9uXKH6mS4TgeKaPwsgJqEC3
qXQCMO+ABmCUjouGbOz1o7+LunUhc4pBCejHZ9cPXbEInGMWJWa9ywUqyqhtZat8jFjfy9fMXLot
/LQrNgPe9WYOl5VFp9LET6wcZqGVqZKTCs2wrzfULz2zWONdF6bdyv4rq0dBNuN5PuukACGdXJZD
A/MmVdcCMRr4Drqg5SEZ1doWUKJmot7kvrJOlJT9ou4DlvEZjF1OLfX4yF274kC3Y4BAzxdGtv9C
7Gqz6OEoNhQHI7qUjubH27VDP4rUtTEGVheVEJ3YQ4B97Tp4az0LCAeFl8TL/nUUi7HOZTjkXyMb
7aGjjkd3B4pddHsHDZxHZUAtYpWegjuNrkher4bpte7ZtFaxaqkbkvLe/vXb1gaOTZZVY1YoAnlB
xpYU4l1LSIFD2oAf8Nez4Lj4dq2H3uQJM7ivilKAEQoQPV6AzWr3jJG6Fx8iVNCoOc790sHW5QJ4
yeZihHOpkopkfnPgpJAigi1St1a6nmHLoOaNpPQybjMuxyy0b7swdTo21Oi9UGvgc5Tqjy66nOPX
Bl7ks8OVv/cH3m8v2FpcoalOQEyASL+hGsPrMMud6hFp1fQ0+21DkyOKH0JgjwJl3awTBmuA3WmN
+sqkhk5PjjHqZoXvNFVy4tGg5hFZOWFrLBkD4UhxM9DKpn3VbnDF/NHNGosazJ/DAX8tbTXE78ie
qJJSgoJcb4lnN4fUErK3ECgzimmBJOJig2+fqvU7xOmNn/DN0fEYXoENmOsF5i04c7TOPfVckc7U
nXS6d3hYMhMf4omdsKQ3Hs/m/UFccU7oSPk0EOMZa8CjwUkR+Q0MwK02vKJWeG7bMUDWfbQOXVkI
35qEJ8L6wkJ0S56plnI9RvOxPWNr9Dh3qt0VIk/5TA3DrVAFkxVYonj42MFIba6Em1JGZzfD5YXK
UYvDbBwszQdR1wjA5XcnZHLgNMz0qbEoPTO1iNeAmRIhCfG4FlwG/7DjNmKQ7MiXzzGjoygSXx5S
Fne+aK6ID+OmALTvN2Co8UDURoL6i52rcs4OklJe642ybnRuxD5pdOR+id0GvH7iUvL/sR3M23FK
RdFePYrpevg8mh1vMp9nHBPOpg+39/nll7klLyhEs2kweZsmxNW6+11vQqSY3J0UnMCdfDpsyN5f
ymvOAS16nO6mP+/v3HU0lVraFapfXQzYZm/x+I6sIOnBOtgTh/D/5cYpUo1impEAYTrStmzSHlSJ
A+No8GPxudVEWPRz9UbhDUT9655APxOjtVg9KqGDp6txsyw15DY8qtufUbSDhdjxLoSJUxiDpp9w
VnAx6ZRQObv1ZOxtDojvvfamB8/kBvK0GG4nwaznZxu9W3b9K96Pd4BvsHIJCm2eXypqnPma4wtu
DsqsLTbAKNsZc8XZYKkylYmaipJCpq8AguusYyLTzfjAl9lTrO5zWZfCO1IBxgMDBE8HEFmKer7z
nTO1sKACqq+D8jpdR4iCa/S3MN68YGhzbi002er8mbvo4gu9vfr7NLCeuyOA3N3YriwnAI5OYW55
/4RMmdtfsRgnlfd/am96Rz1UHH4TDT8MgOY/wYK1XOwO/YFjR/Qzp8n8gpgY1RI84PIFbj8EAKgv
hpqISdL8VR9AR4xivVCr/Bbge0WUgElxB4MsxHynKRJo9JURzwBuq837D6zQ6sUMlvqbqbO9tAm/
d/jGmxpkCvFhxUWi/kg0lVemxY8GxocdNK5odAhfu1rmI+TYuxM34itRptG1ele2HE9AuzLAiNp/
gWNLM0cd/IH9Mhw+HiAA8wsMvZHiY1VT5KvIBM+1BiIK9ziJlfu8Jiq6Xi+XZWDxwhMt2EFZo6VN
QfQxZEwJ2lkbLfhVgWnqo4hovHFj7Lir0FHmPKZkUjLi25GW/W82wwcpTWm5eFQ5v4hDCNaebgG1
wWbBmxm4aMXCXjpf3F0y1NOObU2hYaKN06WOQ6LReWqwCWHHkd2luJ9amnAnwdUHWXl4CANagNP6
KLN21ruAMrO54MdnwSraKHIBZliqUbBuair1pwWp7P3TlRFEIDiwCR4YE9XSXxsQ0mcTQ+RLmQ1V
Av3yF2F+m6j/A99zS+wBzAQzwFPnigWBHbjIyqoEx0OQWVigiTVhDNMUId0fyaMg5epS6wtq9wDW
wrT0oTw+Ts470TbNX+ETYHRJw5rZyIhzfNyMep/78GksK261ZIJxydCIdTV/jdZqmQwXWEUistHZ
TpTtNtv0oWsNUfKT5CjIz77QXRRs6rvTne680RlA9ElJaY1mWS31NYCo1JmeBlBj6T+lJwpivUic
BmEfzLikpPEDcS9FPokWNaytIaSavdUYZK41RChNJJSgQJEwFMSQSzd69rJZicZ1U0YrFLid17Z7
SS1ggbT+ol+XAVOrnqMEf+gJmiEUeBhtQrfI/TAii649jP2CjH4JxYaEFcUj4eTe+slv0O/pcaDu
jPaSrrdhdhsfxBi+cQd5Uf322wq/gkgKKlAUI/e97syP7YTYUkh8eVfyvzvMMas2Yt5qTdwKwjEG
QOiibsXJIflHv+2qqTuWe0/ZxD0H3kMRgk+oRfehRen+D+ruUbSDgsUaiRWRxe9jcVTsYUFr1vfr
Z8yMhXLF0xoxo48trGbP0+4JQSuLc1Taex4un2GSfYonPsjAvBjL5ag90rU0xrtipVjzpMCgezE1
Aj4UevkQOoi5eBZdhn37DFoHq6MEg4NhuAP0RUwwM2jRIxjkofhRuKUdSkBa6WHzKx8IzA0imY83
6bNUw1T2CnDED1DuZPP/+VI1aTRp4xZrrBFoqjflN1SDLzpzoSqXhDpqBAxXHZeHGYf63q1DW5Ix
fOhsucEgSMHCCH2gOVDfejl62IzIUnUtYjwtYg/bmDvdbD2z9dbA7baBOr+oDDDT3/IM76js+4uG
eNUykk2yw1+gdJ+sBIRDtPteGXrOdNdNa/0kSYzdCVS7YoS/vd23Bdta8S7y3PLPyBAm88YtZKIw
IeA9wg71SBULxD6c73CXy8o6DrR0qFkzYb81ozai7ZZe93upbkCMOfSZzdwwN5a9Ffn20pkJucql
ofORkaetdRzG0jBq1JxGbHh+ZO4In32f801aXJrE5J7utiqtXewLHvv13TyCvMHz5U2EQkoajFzt
052PvQ2uBjUYa/9qy2D3nNkysBusH7DOsuqv6fYE9CAD+1s5a5ZweKT+keSCoSnXpEE+TGEwUwrV
yqpGYotJIq3bN9fECiE9DcncUFw2kr9nzAWjnAt83zkyomdb9I5SP4J4qAKgcrtWpnF2HHeMS7a3
HGGAM97Pt70GbdS2EvVlDiXdEu1GKXDbJ1KxHhVMjY1krzzI65FztazKzBehS7FbnOC7Lb/RVCmp
FrvqheQ3x/sDl2OnmZKrmfzlqODaVF7CUZnCnuEYobAR1jVn6F1r9n7ngDovINJ/dE41Dgs3YBAk
12UtQSoN8PEXmbTjVs6Fuf9PY9SyYxf7X4KKhoEkAAKv9xR/VkGObOLpw//Duz50SNGPqO4wPdqj
8xb03tPBc5HRpH2BJrAjqiYByqosBHG0OhQJs5/HTin0NkXyciRh/wYtoGgPOwUSTwe+ojVPmM88
h4V2jgeT3t9fdnVWVdR5LD7UDwjx7X3BGZi36/8uKeqTGw6b8XvP2GbYStco4IRICkUSuzCtEzXl
sP+qYcanc+mv/lwZU38hNhV3YUgdUfMKg1q621SGRAf7TST6u6kkH6FFlJjodUqW3uPkAw0CjikP
hUgJu/MBpmoiUklV8hodk/rMZiq2MRTmaRD5Xv9uKNGWFphtvQW4PBjaTwmEHHsRQh6ONC6ec0Gg
hcelB6Tfo12N9AS6TNMiUQu15wKvysDB37BVUMbEGqc76xwj9lVyzvnB4uDB1iR0bsY1Bv9ZpbfU
eIR2JXcfgf94ny4DxF1xasMues0G++4WBs43+3+jR1OrIkgEZzHRrm9Zscg8cC7/UhlNM5ItBEP8
g+DrxzJYBDrFf2jg3ycho2lO8SqdjxqWi0gaIEuZYLBAwGKsbl/blZcS+/+HQjXAs1vBuKfrOnTN
Pnbd7sDLgoR35EeH6i8hGxZAUfJTqK+pkLBMfOy0257GRPnLxQO7BBmkg5Q0oCZek6c46U97yTBn
CYzrB5QLpSHmW/10ByOF1MTbX4x+hHrdgEr7fgVA6d6lFc/P81ftWptDS5QMWc4YrKXbEjwkStyX
PUDqWlqypJR1qR5O6BtZ0iAHopxRUi/PQZqkpWxD8FEdy9m45eCyUxGCH9uIjOhcAXTwaIplV77I
vfoSbYnOk/lMd6BQqDR5fXpweoSHpbSYFSdtODhNw4wCfCHDo0hCh1JSVvWHQhJQzm/A/aFvJLkS
HRF6keCLhzAy/LHCitgJyO2UXvlKzE3Th0rYhn2NZRiOR7NFOFWYK33zL/pVc47fPRSrUnasureK
N7FBTOGDZaTFa5Ow0og+4ipt5ICUBA36GpdODfuATSibuRi6Mi43vmWyYWs9u0pfuLMc0l7W0Rvz
g0dsHNjH0XR0YjMGbw3Vjj/+Xw6m06O8H12ITv3nUcJ0e6H1KfzPdLBLHWQjPdJDSP8CaC9iiIv3
PTImH4sXcXh/gGoU1sVV6LaoyurGWQ+2LjIKYvvFqNrUdsi1yXVmCsNf6h8peoIDcYEBZMF2KTeA
TVObAKSFLAjpa0gAeFHqrsYnB4XTpN3sJx98KRDS0E95Zp1qILc+ArDU7LRx4WGKebNye/ioW+Zi
0yaUU90R4GTw4EPo8eQ+yJvAa9lyjNgjXojqH4IJEJCkNN69pCBKvEXp3ChJQqvNnpaTmvzLtwjB
DjxkTSwmTkA8jarYsQ88grEARtGLCevIEXCcW/OsPrNgWgdR95AqT6wUMIW1hsMJR08+56OJ85vw
KZS7CbywC28txgQKsEVwrvaqxFTIpd8zIA7djVhxEkAbgOkyjKARLNDUR1tizm60iV0Z3i5Flkva
2S4ggCrRXMwcWs9BfqZRUYZpZ6xm0kZFEuSc43rOZB6KVjArC2N7suH6N/hfCJuakf1C9DOOm8dV
GZjU1wg7yXXwpAQV6aKVh+oHQO4U2aNJfAuI/mdAyw7TeAqfzL5/GVMg/nCXxzcYptO3IHdTauxV
q6WqT/UVgemk+SCQTIYt3OIkFUQmSvqRtTAdYlzTsT8TN9T5fVB1gyClIvx2UsKnY8wW/C4FWzOt
jHkqg98a1XxW64v2tIeQKAInoxFA4sN1prDNxDBwMSK+j9WxR0wZ3/Iz9T3QOlzgDl0xh91OZQx2
P5JFe+rChKrC3y/VR9oE10TUfF4rxCW9jxxYMwSK3h3Jacb9B4MRfk8WO2m1pSAwKRikWHiVThRU
mWrVGYMsuZhL1elJCGLlR4DMfYJmD//90r2JlWIIxIgsGkYFmcVy4XaRFDhR1Z5umoGbD0b2gr7Q
2E/PQeoMuOaPgmzUoX/NZxhKuMU0yiH5KSPckd+kvZTICRPsv1XUKHwNiKy6nmIUonWFySNXhCEl
vaqqjZK9yHtvIk8DuKQpEFTLjAkfhmQnPE0sujBZ7AX/JAGF4uc3hcbFJoozccCQlLxIJ+GzCRut
CNBw8twutN4Mz5VoJcsGcCb3sgnnz1Z19/tUENmcVGS9f1ahSs/G+FCH3gwytM6xqdL9lSPxkPyx
aSu8T0Sz4dBgkQ8HpqO+CZHMRVt1g5fB8RTLz8QLqFopiuEfZqX8ZZSZPV9Tat86I4jo4i6hhVoi
EMeXx8lUTX35XNBf1TxzxFxCMfTNkIxuVAP5h6lFESLmlHUvFkcOB0NDgspbtoKh72sdJCX/P6cx
iSPDpevWqSv135aBnncGc7BskPvqv5rL72W/vq+Zta1vR2E1TI6RrhUD/pcYkMuvxm7SB2FK2qLd
CtnuZblQ5qYDYOBV3ntJfMIXEP1QCjHrryHV+PfN0bqukDtOid57T0Z0sMbRb8+z8Xb9rSyftAFo
fgCO7AOIcuf5rQouXyyOy1HMV8n94O5zKZSzh+ZYhh2xf+n+1R1kThYCdv6G0LXa3kXE69B5bcIy
lM2IfVJqtn7Cnr0oGMOjyeew1no56VYbU6zUOwqQ17wIVPX7dCjq5qCraDWhMIN0oUJOECvf2Ymn
VxfaLWCENdeGR2cu8Ja8BdpFUVRELoCOrm3+shcWkT+9jZ1KJxJzCviM/HZJANDdYlySSXeppc/t
xt33n/i2LRz/ArG3eidxdrMMdTcg474IVlkbk9vCdfX/Oe4gabCaWLL3CJkgJLw26xtxYA3uPOBP
gMYKWxt0obDIAPb21AkeY2BJ9Ts6Fl1oPCtcJEUXeZro6wF505kavi/mdOGdbAm01C9qCukVuX0R
3jCv90Qjk4orv/34j1NpLma96+3/xZUXNbmZMz8p/c8nqr8spH9GEJ/+zusE1KxGij5g9Zs3qbUL
1vwuLPfe+stc0ghvYwsVNEd4KIT893wGMmWWeHbyZKBrQPnQ1dYjQY99db6TnebOJS4iSnqO6BUC
wP9GhaHtIlBnoZP6KA/NtsqWYloNePmXc0vgXstT7ppSvXEKq2NqePH0R9ydKCnT0d7ZkoAY0uYE
9gqjr7HwOuvc/5G2UzZXjuPX5xYkYEaWvChCmcbBJaHtGiclU4HUxZ2tuFD4acnDtrJXbR3CqL/e
G+BqU8ZfgRAKTav0c1epJ1wZGEKIx/pQoweu3RN8gD1RI0YogC5bgVZBhe5G8t++xomhzZ4UfJKi
XX2CF7Fwp6K3B3c/FOdkMSrgEE0BOgq2Ieebsbvwc+lfWgxAXXwV2ruqvog90eyBWxYHZTkhBofT
T2p15nLtciZlfARYFoNQIM0ZGI5rITqLQtEn5uISmpnz51teeX7sGp6eR53Kz2um/R2mryYKe/Xd
VhwCEwTut5rxIA+iBVdDNJviwzimPfTUcCw4KEDPbJpKnz6r2U7KyZNKaze9CS60iZaC3woLi1Bt
nNYqrRXbX/CJ1omCdW60WFY2CDtXVaLaydHX7ghqljMF/v12310L9JkvghTHpQJroOKv6ftaxkxw
w1nFIl8UWGZtDuegZWuVE4hvwD/4Qa0YbtvnMZdApspt2bXrvcWvjrMXOZMsCmkENht+IY6jWyHk
pik4QnKGAtSlnrNQRy0yekCw62A2+VCJvtaJwHg0s1eUvze/ykMvOq06OVjXsqRIHf1Tz3Ez8bfQ
Ou9r0WKGqxFXl6XfA+P9V/mQEhZiPQKq2S6UELkXVVgpos5jeHMWHHvqVwDLdQozDWuFm/PZUcgA
zCyDNxD7MqCrSBuU7yp4DxeSjSM+Fmvpabg7IjpbostFinluuxOpV1OoXI01dn8rF9GHKiaXSnPL
sq3asog7qKfpP48jME9YPdesWj1jblJXf+rleKIZQMJuuHPT9MeJPKSA+JVRVSQamsa0fWB3lDFB
QcD4MzpYgYYxuU+7PDWj3bCLUHylKOP0txFIjTC1oKd8JTbVx6s3spx0xDdw4kXjhaTY0jgOSJb5
1IUoJ/4HHu98kAfVLLvgL6BJmIRmQ4x0qrfz46u+TPLmQ0SC6PK5E2CUjYNV+734xgLxW8xAG4hQ
5ZqLLNDOEXaguVo0wmzjFHJiNv/1e+bvgW/i5amyDv9le2HEPoz3pMBIEU43fMP23rK6TxjEEj6b
vl+T/cs5Rif1FmW3uVS48EfEeyztvl5ZlbJEygF1sCmSuEE2C9J3h833aZeqCRCRMlYS92u9HqP3
rUNQYjj7ToG2l+Yme2Ihjc1vwS6rAQZAHT6DC8I2HfmET0ZrtDTlcvJz1oPTUOSurcqOGfQ9hA2d
s6z4oYe5XG8BEFapvBJTS8C4Cex8JNYJwULJlbcCEZQCgtt/FaJFDI7CR3D2HcXj5CF/2DNQOuY7
9IyESBlu+NV8CWA0KznndjvP7ocGIhW0Ckfl18hx5MNpqN8xMXH/13pR1/eG4oY7b14XxJqicVLy
5WBReAa3Mfci5lbrTQ2Q8s7DpF3OAy5l6vbChx2TzVAwgp9Nt5qG03qhsBa7kXbEEF51y/hFo1Gd
YuECQFPbWPYcM6Haei6eV1yRAe+rsnc0TK1PH1a9jbG6Z7MeNxmCyBdlkygGWJMSM6OGsABZ3BMu
0UwD1Aqlewodyq+AVvFZvYSZ1HLpOn+deFz6awZmfldkIcH3tPqDm/xyXjVScbSamZId6piKItXM
UOhtGP41H2dJcFqWmUGSdpdgjIF143k+VSAI7aJ8gT3bsApsdwYPbl0DW25fb+tEhDXYcZTAkuls
jLXx4R1NbGB7zgJQM120ckk5Xa4vCLoF/HkatQq0LlOur/PwdqYeq/X+PwpsIXOh2hcYswsUPuQf
djKmAC6Fz4ysmCSosPbspezi3OW8i4uFupQ3LPSdDgxxb6BQfABnXt9JF0a2NjISoG1r+GfXUPEW
JbmSydpeo0B97XhML8BbSLHrJ0Xzkdc3yZCfGqRjCUAL7xzMAGDqVQDrIm4kiYpAmXfamJcgyRBs
ZHZ2STmxc6abSecjdPXcunf5m8AJLuZODGzHi1gMXsKwsKs4i5BAe7lUoqj09PkeCeHmEpDf+HWG
msCfm8DzfDNMcc9KO1hRELi6wZOV3z6a+8E78nVhzQrBGhc4CQ2ZLGsbUv9bIqlzH29UShOwEs5B
MmJWXC/Ef7N9/Sqw37g1Bch2/TOB6qYlJChrtzjCCRHJhlDwddExnDxqI3+meUPIT1kWuqJU1oj9
bi5+vGBgvPjJ8JOmlgBoH0lndNphoobgQ4PDsmZSlKBK+5MYTHhz6k1WaAMaKz9UMfnjuKDLjKao
5/G4UK4cViMN2VaaXW8Bmg7nrs5cLD8SkzO5QmwBXyj9a+0YVIdyeBORApJSFh1efA+ap7D4tNid
CtYjTnQ8Yz8Id9lZkZG+bd7yMpKkAmR8zu1GXVJ7/i+Bem27yEkp087Zrc1CKcOOQiRK5cO2RGlL
gGtWHeObGyKPae49OqirVFlxjwzy3zWYXxZgaoAx5rli9bvrFXBuIYiQZmAKr10K/Yn30BFNXepD
9W0ryishENrJhLjVrvkQbv0IyA6fkoFaZyIQ/fcZh7axC68kAuQMD5bO4ItHDD0YaT1QU85+32nP
ls5CASnlLQ5EnUf/4MKAdzZc+NGBiMJ8avS2WB7fa1LZsuD2GDpy8RtQSB0xAAbdPXynfC/7tizE
qg4Q0HpU+iD30Rsr7Bhg2YjDmNoN8kSmBaxHELQ+iX+oL++9aRQ/DDaL8eGslA+wZKsgcoLz41Dk
4H+8OcycF/VEObVAEJ0BS1W3EFct4V4oD18WM56hZW+p1tv5kSlu/XXju6m4KT2Ee5XywqGcrRkz
fv2B8AoOnfVhP6QMBmV7Qv2o34KB4uzZvVxFnfxDQQVyAT8+1MEL+oXRv/w6kttS//OIF0sLDUkR
6HX9HdfZ28ib10kaYpCJOx6WmtuzS5YoDybSJNsX6YQZ255nqNG8fwRLrrR13PZhrpp55kDUb2Y8
4TxTgj1hK/KuLXzNTxRCptRp2h8QIO8pjIK8iY2bRMjAUQMoHETCiTS9jgCIszQw192SmnEcoDnO
+WjVRNDVFGz56H4HvkVGqs5qp8s4laDvYEVHaO2uMWMrVaL8n2OTMWPUzQ9UHKyxCaw5dVqa0oGN
St3d+msGJaeWkWt38cAzAXBbdhi46p+xd405+YMqAa5H9AWLXnqrdO9eYP9LILB8u56eQ3R/0w7q
Cbw60PgBuQENE0X/QQMUNTqiJHySLcmzOM4UdAdwU6c7NmQzYA6lFK24fSqwJ5i+He7hCAyCwwtU
HxK+AJdyuRG0eeADIw1uH9bhXogTldzUkxMv2jmUVUx48oONtB0+DaVDP+ntzBcoiuEn9pC8yDW5
GACEeB3JSTVlFodPWACMq8toNBsfG2yUB3tpkew9R8fInnwHFLY0eBINLGll3HqTacYWgVzoPAe0
7Yg+UE46hn+kdB3nYDNDsX3m2ckorfgvsSf1qo/3nfNLZ5RWzJdtctcvwZuDDw+P95h5E/1pLn4x
RlVuJASFa0tYZU8eo/+A1EC+f7jO+Qb0z5TntuN1o7PClTJXHns5DbI8HmJPXa1/8jj9Q6sW8YHI
j43A/U1JKZo+TTjWvaFJ9JoF90MJyZI66RynYvrH880tKs4ZCBIlMT0uBx1N4cefPwfhW19tk02w
IiOxn+xpfnGirEmPC74IbDdpytWU/y3aZndukQZ0gCd1a06a2Q0lx2ACQAoRU3j8nxpEy7+9gph8
8slrpoTBvT5WRZjJ/Xe2oGGl/ymJipvB/UfTFKEUohHj6CWffGCHHuMiXONaSGD6FLLgmAQtJWuE
zz8rezh5FuTc8nt6N30OubUyKQfKF7XbJ1b5jdv+r7yuiFv3ZD5//rwlayYnIruxeiY25kMJVkUg
I2gugc1ncJkiGwfZrsuOKY2AeAV/VQdnoLxC/vQbA/QaPuyPlP8BzwrJW5RCwqrn4FpRd1uwonEj
Cg3Cd6B2zJE3zTE4UEdtxVMTdj1yQ55PNKhKqxeX9kyFTzR0/7zc94GQwZe5koMy+chV3t/LUPqo
FDuPXhyjbum8h/H3NHK6O9AqmPUIAzHNaX5Pt4oxHJj9MK2EHE/B2kmWRSuFgzr53+Sib/UenN/U
RE1ux05RaUCGYuSef4UHMvID+fQjxIxiPujgaDmHLJErWt1HEkwHmECminq65gKCvfPvty0f3xxm
or9opnlFTIXnvt324luOJplAk21HvLTwNhLOWYvTB/LRLbxdlhMtIjWf2ERGXP7uZtqJ5Ss9AnNy
fQBf3dC7h/U/01yaPp1BMttxv7dMbR2/+5Sjl7cJcMxO9P7gmqG/bQZmdliz1v4SihameBXF+NWl
JDvQijSMZgn9fu2ExSrKkrypg6Piaga0yJSEViPYp9SMSHnW+2FmSCAvZV6LIW7zssYaBaMnJ+Z3
ONtRiC8I+NgrgtSVCTPbjdw45zzlwvV2vZtEJtF1G65Ge+MnkseZZ1xHs7iLffc6XV08m87yvBDC
9UVdEX8hcZTHtw3GswHVglZVcyUXjMZZpjwWWHcdC46UaxVLWX0mCt9kcQH1GbNj3/BGOk/6Jky3
/wZaskuJw4gAm4LxvJXNzV16KTsMtffEQFCx43TSEsJfENWsUa6+aj8DdqBqMucCmsIlySgvH/29
7k6Qa95WCgGV6hf3Txg83aY5nHKjEZp6VM/gHpJ+Yj5p1xof2lzBy/kcghvQ+04UkiN1XOpFXVnO
ISU8NXpbfpYX1nUy7WZxcoM7S8az1SOTsyGcIuLyBBuxdgyi37X7ZBr7vtipxyj9C61j5dhr4AjK
wthmRKE7Jz1/2h26LuiTecc+VuOx/bNPvOSKkjaXLUmH6HKeTsbbWUn96puvrBPy5U+DXNs3j8JO
Ei75eB8Kd/ixaxV8KWFulZ3Xbm4SF0qs1YWavooSl0UHw4T6ZMejXpEaRO39tV9+gsfWzUPkDDCZ
/8EI0lMxuKX0Bqc3iLrLWlO6G0hCtYCn8kioKuzB7l3ny+htC2Ls7CjCh0j94+t4GliZ3Srnq8Nb
jmqCLf8/jLImq43dYMrpI+gH0maD8n5m/Ru1YicYQ1bMUGzRNTqqPk6ivoTMKNUAsqkwUopAfpmU
cHcz2Eo1e/5mC98cPKrOeUACN7DvxO/7ZM4+OyapHb6N0zeWW2rjwmju1VmPMG1TJcoY/OcPRD0N
powF3yWJnMQ4PCmpWzUtC5z8U7o6Lq34dmX4CQny88OYxeajX4OaOFWyTlBQQWHyBdHpup4Yh30Y
zYlaVcQwLvspyZPJ7HMRF+21cz0HFDhV1XKa2Dd+pKXz4KDZ4GE69Tgnj/NYxSCk2cwvq/M0IX+h
XZp0fdawc8WIVhUeCtT38D5lz7hGZgvPL+foVDqXUuSs0in+Mq5I6ShNrijGS2MNIrLDabW/iNDl
b/GYHqgIz6N1c3Adgn7rucm0G/Qq+O8EvAL0X0jj4Uwdo5CoFdWEqlAbiSGQr/ECz2QnixitTz2B
9DRtHRJpsa1I7lbx+0Z/AspMPC4aa/Uwp3Mq62wU7Tffq3c4ojqv4RaC0TqgL0TsJHc/yJvguXXU
CBSOyZmXwZGlcRhvLWtlBnpYOptC74kqg1n4mtyuyHu0WFJO93WeRYm2HSfxStaSOPlU40bHk9bi
jq/aCJELE0WYYxBGicK8WRvdOLvdpN7nZURoHiQpsrDHkUn20B48xzcpQfrtsPhrP6Lp4QoPl3eF
hi04c2m09KshjDkJmCzZTVbrobo9YbqhnbCUc5ROWVzemMxkq9q5XSIJRZ+QQhQslWbQmOZXHWIT
x8qLnzScWU5xh2MDFUPL0BhHZT2Rcnf8mXrExw0ZP/Ah/aR7ejcMeAKYwBvN2r4fcXG5VcJg9uTE
M4TZO0f683zkpgPkPE1bzOEnJsCsp/2PBq0hp4IR7MtP2ZdKJHrEfn832xzxKo50Lhtvc3y3+2al
dRtj8d83vxdJt6C/Rwq2Q8Ii7BVye9IbpOOf1gm2PERRp0tzwaV1X+pcrngC1KFrMk+c1boBwkNR
r7k1RnC1g8x+qgaleLVqD/n1H86yfflCFxGabH7qm82Uu0C+8qA/Y5OQNtMhhKK/MCMCUsIOPGsV
x3y6jZYMOHshdgrjw0l8lbgE5VQv72FkanPGFIYTmyPyjy5bxpCRXchXsBz5w2SNh0VLjg3KSt3z
4rhM6l2WWnLiIrNpAsYEnp2/N8eQCu0IBnWzleQCNrhg4QFPs4kNnnBxycYyijYWd5UQn4/k6ZZQ
E3MJtPsfBvfcXYxLqtMLOx2mHKmhEw+1anCDQHZ+49u4TVr8I1cCvY+xBhFHa0wcBOLSFO07kUPX
EjjIE5Mmc4Sof5uZ9BuJTHqpzfBtaMSXJkqLfQ22iX4QImQbfUbPcEQQjdo4gZLYFikrqNBV5cAa
RjBJohvbFUCR+auyo24NVXUq7gtZpArYgEhTiMyIvwSbaxYAXqcuvfPCYy6GVztsnQcR9tfOnIXy
c/24PyxyrFOvfuyLY//ThHY+xnSQ9a3rEJcxyCfV+I1Kzafs9z+WFVYZW+IagYduQOHswCzee6yh
+wY/pVupyJ+twFAxtuiV09mouMBdR9sWyAZiFQ4lVzL82VRnZA2JY75q38dfdm7mrW13fnlUjsEY
W+6wQuIofUynZq1uB1t5MLRZJhXCy9bhNFwbThnhF6mvPQSJYSDdRU2tZzz3yOu1OX3WTxIo5TKY
lRP0Z9YaykPZTjP3RKJadqiH0d9QxXeA66iyQaZpVoFDZZtiYT8AmQ65WwqhYhk3TM1Wnu3UZgZR
xvTSfexj6X6o3+z/79DUQKr3JGexjOaEJaJa0gj4TjvlXFpvCIlXj0iMNOgdgwOECCHr/DN2yPxg
yygQ5XFgmEOXY+dlX34mKUnKM+z06j+ULtaDIF76Tp3UJwewfrzE4l4jJmWF/kg0qn7JuuFPzg3r
j9tsTVOnpxMzK+W0EBDRBKwO4bAmOHtIR5h8ophAxMj3y823vzTJQlMqZQv+Dnbe30ccn/5SeX/b
4pEv6LUdDsGHNP3h031F3M7Ke1gShUUr6NiQx8fb6HUKjf5f5X1G7G8DeXC3v6UArVgX2prGhLYe
/rC8Dm3iAtuueQh8kzpZWhNqwMTqiB9P95UvC2VYMr7UoFgsKCeLLuUucOLT4fz66XYQSRgxDCPa
bXW8ioNgfnXFEGHDrl6GlAXp0GxKbDARVAZ6gEHu0EsqPn5Kq/FAJE+VS+v949cubTq3ikX2d8/B
tZG443joDwYj8EGYPb/KsFyK7JopqGccq24PaVPIUbJAuJiEsyds3Ht+Q3IpB/8xvtOV5CpQ1GCs
NAq+OyORUY+Nwxgr277211ppVbCxr2s4GzUPtK9Fl8+OSsREdpPvNNPjxx8htqzNMk/ZScRn/A3t
S4IHdv4o1GyW++khyPrtmYUp353IqX6htrJ/s6fx0skAA3Dd1jddq+Z3vMTVkr9MAzfp1LJRZdca
2BNChTBP8nbWqi7NTlIXcEbzlq1dStKPim0C5ZRaOH3Wyo4mQbAlIjEXNfNbUiMCXEQG+EaArZRQ
VnaF6MDN8WB/xJ82vy0mU+H7tiHrdk/yNK3BtFxqUpmC1DdwBXsnZjocEiGjYuC3T+/rizt7eb7/
tm26Wc0SdQTpNxmswabw/KMB6gjMb2z0IgUcaKQ2zrkABWOcrxFbSlgZpzdbDmX4IKrwr+sKBCvl
bBys46T/K2dPG7/WjRMcHTJ38OqohE7OjeYWeewSwQIroGQyN7L8hhjEOmiqVd++dqwY8486yScN
BywrBKnr0dnRB4ubEzpGeNoI6otAgoyLeRQWC8lLsK3KXPk05RrURIi7H3F4VPVzk58L1pV+3GKD
qE7ZpZYyjTeim+1y4eA0vL7/eSMoqjTDngQzM4V0X1OEkT1cQL9SQIUO2dMXOWItAPzzspwj/N1F
J44TBfQfkUVLFWXqMbUjAXTk8SYlInsAByViQU3LIwz3rGs39uIt/+Q4GkIbkai2g1LYCfOs7/YS
Y8TH+FMRcRC1gapP4i9TLSNWdLSqg8FmekBsnkUV3bc85uOBJMsE0dPipRH37SyqxAXnGw6vcc/S
Ro0BazTVG5qCeoGaaIp/ZXKfP16+NMz1trnobuM9rWBHNhd0ZC7ggq3leybbFJeFR1kbU9FWiJ/F
5MmCWnh9e4K7FZEBskwBmRhLDfyzdRfEgzhOUixRB6WXv0H4QVvA2ePA6s4//ISTmoxx7pYobdp7
PRPJA9WfquKMwQPcU2qYi2jaMoRbxHpZc2bxnT1B5P4ctwzp7S2yIh58xXElqOL5x6Pg1gcHIbmO
OROLsRYG0LEgumlP+39nTQeuNEYZ7ZhMiEP2leWYakz1sWpr3TUI+FzDbjoOoqRAU3fnYmEgA/i8
7x4bZJ3NkEv0epjtAXEtZxBIpRXb3kip60MEE3q05UBrFcJVhQWpla09FzWdm+wb2znEKvEVPml/
Sq7F01S+otTcapIQebUpfaaV35WyjyQhGmCaWXsiRNqWScjZ8P2TRbLDWjtgragh/IxUidIzsDw1
L/7hXgwg4WaVAUnmx/inKqAZBcuMfntfCPe2/PfImDH1hf7XVzUBtlkQYg+gL2gSlONEXw67niEs
VwN91Cyc3o2WFJgdQxbCFxWkclgei9O18BE+lHAZDBiE/tDtNa/ZqJKdVeLkUPDSw5imbs6XQ5uE
JTPIYBgwx4E+WgHQkQTu9WODp0NbwHGGry/uLRat/QSbYsgWHu2ogkYFzhPL/UjpceOgeXSfH2h7
0lMV/s7COsstoCfbuMozriXVJ7xfi6btq3oEtODA6ph6LwJNCnQOTQxwOchXOzhvAeiVEguhebvz
X+gpHW1X/hKSgNKSCZTpBKpCfttWT3LnHGgBgak+m0MYfv08XtqUlNE7ZYnnQbdbXGtaOM7Cx494
v/QRBRAWYfhIA2WRh269inHCdDSmepir8vFhLlgedSni+KRxC5e382KlQk1jQT6WpwTGHzfx8FtH
K6GFiCw5vmBnTVkypMvSFr5a2Ff9GD+6EC5gcjhczuT/cJMxcKhfuSgCeqwma5TkzKzJELRGxW/w
FKFnN3X4G2pl/QOM4WpCHF2MxjfzFEqKwyAeXmaLxSJa4KJm1TmdjVz8lpBMZy9BfMlKtVdf09+z
yN278CuUb0eZJyEV3Ds7Pgs5wGdxvAkG2+YacZTcMTdw7hWvQ2PkQKckUx/GXpn+iJuuy4SrlZW8
0/CETNBtIEs8hyXiATUT/RMSLZ+qNfrHSK7HwyG0Esn996aGWHGg0zGc6s5pEsPUp5OBgwFKOGlD
UzgSaAFt5tadbm2BKqUZUavuODqGmQORV+oOthbIRA/y7jm7f5O6oCa9kpk+SDW++rmq1NjBvYRA
Y09WdlJ/yArDaKJcFV41eyTWd+j250InOiA3cTBZN+NrKNsUk6OYcVYRCNNWnxUXXx14VT8bQSeM
ObyG6PRjIxuZYrQG/k8R66rOR+FEFkUX2xflvPr5+v9u/TA8Nj8N7N3k/uT3epLTpj84Eh93nTTN
5anNRRE/Bpwb2myxUhdQ60ltCjwDKmQjTFdFSTyie+aekVa3dnV5scjRm4pKd0b3gGHgJFkLgUDI
JFbGqq4cKXkPep+pOgANKoGBWmki1KdCh3rqIZWFbChtG5uTiKUeMnj7Tpf1QNAzEIi/4v4SQBnR
jO10JJAvmxdr1If3MCneZIMa4y4PZlFowlGuq05Jq5fXsJVVewQeeoSqs2beMGKJwD6N4EDSqceQ
5h9g5Dq+18Kb1GeTxTO8l3vM5Kv2ymTMwYffXTGtZiqB24wlJv4PcZt67usQbdWaTt+zCiqs49Cp
PZe8qvZyq/5G7rr94WlWQ6IyMrfM5c7Hl6KV1zzCFyaqEjdRWrpCwnTY28V8Mc8SgDW88wNKAWYo
bu/sbOI2wrFLVEC3Gtn+HWq/+WIcv5yDchVxu8lNNfTtx++yoEHWgN2hTa07NuhoVUlcSrrtrdtu
hqx/LgHfxz4Q0fMgSa0xEblNdeHyNoQ2g9qT5DYrzDC0fzHZpVDLoAbHhzQ6NS2ih6IS2kZut6xT
6RjyPKLwEHiTtxKvgbzgoh9LB1gqt+FudxNdmgYVp1CF+RXukTNSVlcZC3nyo9AbMzhELyvC3dyf
tUSGJOdyfckHXNY3c3J7WRN9SOKTpgVb15Uo4e/sHajtgjw0C2zQKvSUQw6VfiIb2CbggZBb8Gkp
EC0w62GPo2qCcLShNojAIy1FcU6gzKst9ppxqRKqPNhBP0lXXxiwG3BkWcy4p0G0x8Y1UA4//65Y
ErcrWpBFp06ju/qRXskE/VvOFZA9AGkn8MC7Zvp85gTBfLHE7v8tHqDUZvdqFqXFr9BDOcGQPP0r
lvFA4Ixyvpf+iQxviccxyd+LZsJZ0VPLqIlBqD2xu+WsZV3rLOv+Pi/aXeIUBir2OJbVQgRKoRbg
FF2aNvKaqXn7903QyVZNBireS1fQc5PW3kb+/VM1mnxAaDkuzc+ha5c5knYO6vPMiJGy56fWkz8O
Beeat0+gJwKdjakMPiAfrr9U5TQaINGIRoWH0obbZVqqsR5FsxnlQac7Qbg0bpFrp2VflKxt1HBC
eh+P+o+GDifAzb8nH7VNq4nFlK2WlyoQIANtwh6YVACYK/IyJeDUMaf5hY44idLpSBemd5TtAzax
dA7j5+rMgGnfm5gFxeV8XXPAwGJk+qAUIN56to8jTwNsmQ5ODt5hr1a+LFRMebwi0Qo7MlgrY4Gd
JGcpI5a7PD2reqmkvbakA0uGO/0cnOyEt+Fviz+9Yi1IFRpdIag7yVTWH+m6CEB5qUUAODtYCezT
UPi7nnvxRfjN6PImzSAU56rmG1CeWIlJkzVT0JdbGg4ReqKVf6MAx7QDVpFgw4WUxKeKPXrLchhO
zJJErg/LraV+3aRYOImh1uNrhTKWh03Uv5yLMgfQ+86BEUuy9YJqTZeGtY7Y5DsKiCrAzvjE8udC
hdbu8Q0lJxGi9d0vLltDMgUSUWyMyu5Dv6tthXtmjCyF8tNpWK3vyzcWKTBdxBQAw7MiljLDY8+T
90J4yyugIx76BHmQ44JqRhqGOPwCoVodvrGKhGuaBlI5cc/DetvvaH+UFeTdmCdCtmZ688q3hHFr
gVCnC2EtK3Cffk2t8XK1MqRYmeLBAonqeNl8qrdvxS/cGRPxNRIWAiIu6/yyVyGeC4EZBPjDsudX
GrmtJGY4/oQO31i6Geb2xtpTCxbbRFEjNKwKaGlzaUaMWijUBbj+TVnILHkV2Tjau8SH3iYqVOXc
CMl1L+xbqA4dGTc8iP9+at2bmlhfA0etxeRMpalQ2zslI3+t6C+am3YWWO74b2oAfSuWfhmwU9Zh
rzFeBgAHpZMwMejyAzY4L6AUJRdxVifpFXH7W97B7LE5jBEUzf2rnO7U3ixSZNiyj2W2EH4CeefR
XDb2ljxBvl3rReL30AGU9ETYXlrNbbdzVZXIizjTvzjiBbSPVn2XYu1mmCoj6ixWgkCSiHNr7Dci
XC2955Qs5ISO2CQZUqjqPMgHZbygpFmuO0kCASwdshpUirjFuO7CMUQ13S9RneahEpA9eSwSFlN1
UjSIV3Kdxn7dhu7JeptnBI/uUqMjOxbUmc5i5/56aXP5inDY5ioq3qlLLsUMHghFOHwjqPN9HppJ
lik8knIRwYv4PwTlVYa6OD/u9h5VbScfFZCxIoU05Q/npVTzkWIgeoc3IctSiRXv7Fa+PQu+Fvr/
T44F5K8qv9wpkbWKRxxaydsoWdQm174AtihOFYxQowad+99jwhPAHmgps/tL1/kSh4t85puCjgms
o1sOVKpWXSjNAVHjie2mcjwcU+w/3FUTEGK5BfLdTKA3zrzLMGtYs7pt+KFZZBFksgoQn97Z/tIy
OOcSBkyOxC/5zzFXGDlI4np3Yb+JYRtMNcg/igWoYXPJLfHIsD5jmDm8u6xrNdzoRe9Ge23VCEFH
m/LQVXL25ICidejSPPbA0AC4nnHLc/9ys/kSFfuAHvB1Z0CKwGIK98USk0YMuN724XHkv/daJ4eX
D4Ax+dlLAHfzBX1+ZZNaQSGeWK83p4BLZEiPoY8z8P+cov0I9cywwyDaJNQXJ++SJtDLWA6z1NVW
jvsOXjMcMN6gPNw/ZNefJRBOw0zx/dZNMx/O8HdjLzHFpLKe5o68PS1qxgfShKxkbrfGCNdy7e/h
Au40H5N3OVhTM5ut+GrN3b2qyRow2au6aEuD2Vy8+LjLKkoWpF2y5p2Pj6aNiSoSOwG0sbjpdqmg
+0jlKuOKWdl8BVOiZl2pZ+4UqN8PUCEC6+Zd/tELAISjUivgRxT+JNuivUduoDmjYlrRQ8Z5Z8qH
0AGkVPoVuSOSSc2cQ+tAtDZ414ubakRrBgxTI4JuQSutostQ4erZJgtMsYzHCYnaUBu9+rFAsjRL
4WwZCBjAqcMLE0tQLzsuARXb6xP+zchwxLwYoMTXX9mp4thsQ62VkQS4N02c2R3dlYswq362+nTI
k14qJx2OQ/YTdlbSKHrTAXp5meyD8H776mFV5Sc0LCieFvhdwJlneM+ulL42zQs+3mpp72RIW7E0
lZE19zPjf/X8d42VxpZXG8MaprOURtU0Rm0MTEUgA9NkHehtvM3hxnfCbkQMgbXg2SsxjmuV2L7q
OtUfjOpTNCp03b54EZkCqK7xlcIP9vptNjG4HldkZCZPJlK031q/IRn8k/L+J1GkjQ7Ke/IrWGgO
+hOjIfvuTr7yKEmUBTW6SAnBn/eqtBzC97AZxK6M7kRJysn45Rp74p0vGHbU5XanMlzxtmEUvCmG
y6zryYjNJMde8dYaFyswjpm9t07CvyXHD3mtWjhXjCFxwiNbcMdWIIo49iDktKOkystQw63MRG4U
N4DNvLlnNPAHjo42oNIPV4KIzwVpQtPvCST9E9Lj//AmxjrftDX+YwYn467WpD671ecMn+nUIjUe
QtVTYGIcQJvoSPciT4/h8SOkkHmKaICvJyOHxHZjkilnrcUfEfdYOILNqPtT90OWAGsXcMQCKJMZ
dsxm/Jn9Xh6PkRchCc+XbcsIlTZAPopfdut06uMspFNw/DEbE6tLoXnhHimjlSFTgb9ncNWJ1w+5
waraTrMer0yX7LKyx95cYpQoHlQOwSjgGQxylL2IYYJpKnOC26+C6DsAAMLOfjHzhli+WhvXro8i
qwCAAAqnFnp750yILPj7QuyMGSDQGTPBZWTjpiCoz9n9NUrp5Efp3J3tZMZ+iQhUtK06T6QZxGfb
/4ulxht6LsPT+Ko1waRWNX8426GJKjd2VMtCRAD1wyNb15h/n8RJbEl9C0y6tB7fOnQyk3VGI/Nd
EZfIl5uRyxtl7LcTDEn4TM4oBKWclnIicSVkWhJkOm6HYxLp+GQt4+rH8rdK4d/2g/1rVZkV9yIw
r2Fz3NYtFClPMOVQqjePMywW5yxz0Sq8DtDs0ZsWkeYyImfDyTolXQw0TLukNxoR1icOYAN57+vq
FJCBuJjHoTQGS18SF3WU4c7CLQgOhk8MkfxCNgHLu5Not0y31rrTB3x4mCx6mPXtLylRl9d3y37k
Pwhz3HJl8pAhCGwgKQTN1paxLJu06q85NaC7hnp4kYcfhcf7cLp/ACuh1T6/Xli0xG8Mqiq7CU+V
tTrTEUHk1pyJifiRD9Y/v51uuhxMsFaHY7li9NY0qEH78f1HYY6Cmi7yEpMDWKZfwTze3Da+S3Wh
FIyaUS0+JatHDExvma7qc7iJuSirP+oIhDgHnXimutuFrAf5TuxiQJbJXy/OoFYKGyaOEYMOcMAJ
vweBbVgzkwF+XFEJV8hmtXbU3GxPOwSlULDf9MxUYb12hMdM/yVMlSPck2HSte5qzVNcanotSA7G
SBXS2hmSRqCkFiDX7qqUni18gH+POCqZsWmprHaY5wvLnRABYsMh+7bi28I8IeEDnuDU+UWb4KJf
0dfkm+0zySLjYgXr0z+0mQp9TqxoOULsm7SWqWeYq9U0qwHPs1sYqAn+n/Disd5hTjDVHCogh7sD
z9nag2CNh+ZLiEUhttZu382mN42Sz23Sh5Dv3EO9ufczmIrIoVjS7uRQZM0no/9BxEGOdYijeHDw
4b0e+DKkATFntSAa1CMzi7pvdgth6lw5chwmdYGqNpjNwtq/mV/8X0xx0/vr5O2bOHUk9RVdjMPf
bhV9R8NTS/NRb7kN1fWzb2+x9qN7v4L80woEHh7NdRXrfKKv/755/PX79AhpYFQoB7ipcd81rDTF
2fhYRejs1e+AWL0X/PhvXAC5DwQCI2C/4hCLBLMUzGqwwXMY/NckZaaBTT6A+YApB6sKSY6AFKAu
9krbCYwTaDdMAByNfqPHAQ08QKGFyeMM3zgXdRw2RjSvlEUl8PFtTXTC3/eoLQ3JUzsIATnhovSH
rleDGhCiuuSJNJxnDNCEiG7aD3Uq9NN4Fworr4SgoSk8grZgHbrA72EShr45952Q8X8D2O71EyLZ
aZozKgRb1/3ezPM5Vh/IicvzULM/mcfPPR0m/tw7+8DZM5eL21j6+7dmi7LyrOyNUQpPtuEobCcX
cFeMiD8F1rfNfTEouPwbl+x1+ldZiGJOc1xjKhhztqM79KotHTvHpL7XopOFZwAjCBmTfSgWJNCv
8tmM3FRTm1MBZPNRMuAmhStuDkLAp1tpLAVXpni/jC/0UQ3E28soAuBRa06GZSXuPDuBIL/oLvF+
tS/jQZE0rRsMM1dfjM1A0sQDb+hdaeRi7T8TiQyv/u2PLJXlLbk8mcHF6wR8irZhL4Pe4Ei3jtf2
JSbsDc0cD0tX+hGmJTWVIxEK6h3sARAIDnVrPh2VVh4NoKvTTtqFRqfbs/X0We1wJWfYCQTgi1Z6
S/NsCF0MYdSxykcKPsre7+8WA9oXE+QokG5VWanBIy4DAAyz74VJXdP1uFnassj/CiHjGPsRUzU3
djytEICbfdwaDv8gTv9O4Gy6LcNfCH4LDt5gBa4zTKdpauT/glaSKlUDh9XsyFf7BqMBcHOBM9OR
n+DW02X2dHhCD4zFbmnMcAWA+C+RzQf+8bj7PZRgWjt7LUv4EeStmRPBPpwnSTboobdsodUkYwD8
UcajW2lZqvkLvdrmukpteqVR85budSTID+/DlnYDdHFTQ2JVUk1xHtXpCsbmInm4GZHnZi5awqxs
yt6y89r4TD9szbkCl/pgYnl7mmXkFpUeN29cy5V+U4zk3KxKlOURZRaPVJbc0ikP7n1c43d+G2bN
1rujDmYJlAY9VsX9CJJ32x5uwhxt4QMUDCS+z4KfJrDSw1t2DR4yHulKzDrfclqM0iKkO3hfc689
2joGKxTzAEg1Q5ZHMsHqJcTtZl7rchKk8ub13c1rfP9KZOfXHohwDXg+o4bVj0sKa3vxRA4bu32J
qCnDjNw2n9thPePwZYq7AuPW0pLFx7efLZa7C9tXhjQTdp+32RU0d65ly/Sla5NyK8DmWoVIrJDk
7Q3Hfjxu+ZRuH4RBYNjtq/gJe+zh8ON7XmLXws0sIX2w7JW1yjZ9Ds2/O/yLzWKm1s/r3TIm5Bki
1BEKl8eOLWbNnjhkDaLrTx/KGliYezMeFJfQVaYWZ7vGogCQ14jTUKSRtmgyEWSfkSCJIsWj31T5
kaD6mv1j/d4AXvm3ZA25lVaKsDw83BORNbrGDe3Ax1PAdt+XyZh5erm+a763JhSLi7ViPo/J8Lc/
IHO+4cK7WEWqDIFsUS7wAzJbN9nMeobUVhJPVBVP+VDO0c3K0udcLmTIE0e6ydf9bdnZyKagjWFz
Bzm5j2OGpCzWfCkAnF3m6VMn2nMFFUgeuEQL1mBGw95jXLbw7LmrIYO/XFNBVEUCY+amGq2ypHdu
Lxf1z6RqzsdSTQGKCNe2jgr7h0Mdxou5TQDdO8SEPRDwG0yQ+BXLhUoHZ0mxKNz7fk5c9RENFdD0
U6Oh04qvXV88BROXuF2d2LjEvCho8JP/EbeTorSRHBELGDhdtyxF/ZG4QPIg1dRzVHanxAlcY48G
ZDXEnrS8+4zk237AY9rfTVVyeqsJAsnLRpn4NPI/ZJn0RsW8OChsuzor7QTRhtfHJLGnalzgvt9j
DMiBBCdSNFmVudEk/8hRyqxwXmClOgSjPyBcDTHrya0GznrQ/4BjZRXULmNllieYqeeQ73XXJgek
HTry8g8mXMGxjiIJBWnSfxOuUvqKjEGodV1+TJmcjjzvWQS19LPPt2EgXqYJ5quBY7J18M0jMdCm
ADrmvR4WNTxQGyO5Kl7U5+UUjBLMzQa+LG72djJRV7Kn0uFTKJ6qAs7Y5bOht4VjTr8qT+XNhiKJ
8uw1OImpGAwt2TexiwOvi5++JnQ3Mqi/vlKs1eIj67tPSeCSs79oRcwz64HbTG5qVXL5nKqhmOb9
9ZvjkwO/uQXzMq4QA60P0vGlKKdxPNN+6OYz/vRFIaJ4FVbROBSZWSau3aeGBtN6PDzEWyMWnMLl
F/QE3ZNzHyIi4CqK8rlncVHLf4p4A9uGNbOH1GRRuG5RONGMR/yaenfECQ3xcwFrnQW/OuCv2Jc7
r7gysqpsKckr8X5DYjj/qvmiwR+bAlvoqDbHfrQ6Ou776aHopEuptvQtl/HIXcNk3huuMqZ2UreN
0e+UOxbSHYAyRWCXImqtIDrgD6ZJbYZi+21ttdK/9IPJVhQ2XOQNd0gJt6xKwsPpmITPmOFK1pm+
sMVzqDWHNtwinpD55+RrQ/sFTVEh9kCmLh2Aty85648AE3edcFVrbIDqegGGWRV5k9gk0iEn8B9K
rVNvPaj8576gIlZJqX0+x+d1HeSBi4IGmE4bezu8dPWkZW2hAGjiPvUfigz7ahPtOiIEnfHi1ZrC
ZqkmwviKVMM39XGyEDRGy3x/9o6geAqAnQiK63qTs5gX1kN1S/A5lpiL2WtwCNmLkhst5lREai+c
4Bu6z99M2eHzLoJ9hPX/gwffCEqP9stmMeimv+YRPyC/X9WGPjeaRXV7BNcxftxyt+24sM6PwttX
FPPl/G6W/SQ9kfO8HzVEub02S+gwrZUgRkILsf/5fPwKLBLEzdBCdgxopk+/S5MTiAwfgL3Wl3af
M/GkJjxkohnRoTQSAnAPqtSkTvTRLEdI/CuL13pUbu3QoygKM5OgGkTCFhNsUxGebl8RKpl505/I
pMagqVF2JbvHJ2B409jBnHwt8XLo1uprG6ie7aXd+lyNNDAn63jkYLYj7x5oAiMwVY7QWdSIy5Sr
A1Gru9j0XbiX/Bho6/NynHW9bvDbB217FQv6gaf5bqVdaLh/5FMrgRFRV90c0AAoRuZ0bYZd7DI+
/Bk9NvSGNaeqnuzfEh0kQDnzBaGRIy/9bZaajKkabujEw91FkLaKGFfci5rs+Op3ktOw/XmSY7F4
Fwbbd3JhM845A7f5lyzzuPfarYP7R0cUcSyo2VMsheI8s83diAXjVYXLgdNrUJeCQFC+ALwc4IBy
pYcISgdOAFbd6Jb2QBPcM7NLTSW/o4zDGGyeGpGz8aSOfIPYG84TAEVVAIvkoecG0T2pyKmuA8HF
a6euUGtGg1sV4Qa58P1Oi6rUjj2vQwtHMa5U30/V+yKMZqG8uKLWWWYMs4Ui0i5p1hmF3oG3pu3e
1Jf2yhwO1n2G8nm1yd/P4vJHdsJzeYRHZw9yVTBSrWQCoSbKgDFBT5oK7QhJwxUb/qYZJWIsnwG5
oysgwjXIRe32peNGEPElEok3C4bGBzYNtbGuP0xywVbVVwQnreUFAL3Yp1q2ZYR1QVTT4FR/bHVP
bsteKcRIjsWzQ71AORIlOOV66PXN7yehj5Pc80hk3eCrVsvJtI+A2h/ucUHJegzuGLxGk9rCDQ1x
IYJFnuzVGhShR26HONtinpy5vNYz3QjiCNUBmOlWFlosplLwGLoC0gXkTMuE6ieY4fC7Ii3nLyZB
vZemKJEJb2iQ3Xm4LZ5l8nu9SFR4QuEFiQUofpVsEC4u0pfFJntfazl0q1afDV6bFmVgpkXEspwd
SYdnuRKEK8m1HhmravsMTvlm2BZNydmOe79vtwtOgLyyuE+g76h/2eM96HmBHfSL1oKlkXwx3j+I
eumF8iWCc7ZXf70ZX/OQT4ec4UxwxlIn2K1AFxrvRsOROzOolHt6A+/BoCI5PBxxobDl8KCWl9BA
Y+CbjYi/KW0e8QSc+WREF1rS3sPibGqkSWo8qfzgnHd3nJPAaDKDOervhq18kE6YrfM0+gzTGCEJ
aQlG/g4o+WPmMb5iDXnXeytTGxV7U2unVMWXbmPRyYZx6B/rhhcbFGgNTgkG/Ffliie/++9lLKyk
JAlXqe2gsiHHuyIKi2HlV35Qa55akvKotd90iVajrG2dS+JHVV0fu3XcOjXg3ewPYUNiDK/dhHK5
AzIDMrgW5JjfSZun9jRBmPvpzuriGKby3WxxFzEOcjKycNXVo4OZo7Hi1aN1t4e/6L94xGdhhZ9L
8kIu7+YAmZ4GKJHFsUGDecUS43E53TqauZjqEc2lEzme5cZFlCLH0C0dOzLJfRWXuwLvQwfI1TgE
Z8YnvO1cNzoODzvdiRTAfGFGoAz4JGhpcsmn3I6chNPmgmii8JqXWRHM5/weEC9kvB5OxBu61c5e
Y0yf44nvTUdqj3t7CJmi785vd6Uj8fNbdTJsImrWImG53+NHOnprA2fKZiD4I5uG/wi+1PnO+mhn
kb0f1LyCpIsACRDhgr/LpyVlJJ6ZnB6KekOPupXv58p603fRRFDDgD42aDQt9t91miVj9KIr29/Q
qyBdn1edbCQQU7OM/1K/d4kFhXsp11tKzqjkFlxzjOqHzE3YuigUMSB3FD+D++Ngn+ionOuIKDH5
o4ykvNmj1hPbzHMA1iWSF8UDHZQudaxk2JDx3Qx8ziuhI3xGLRxeZOEC+aio74gfXoejI+jLwciP
kCKk04ZrNBVWGoh680kvLoZMH3OLJgzWJpZSK4f0oTZ4zmBMmlCSAGH5aoKoH5u2yqtiWa6QuQpV
mkHD/4rqV+GXrY0tgpE/ufgXM2labsELNop/WZQTc04txwe06pgJknCp96aJnmUPzE3EY5DwfD6x
Kfo4WDvebJqagQkCb0QKDelLaGcnMxX4mSUSzGpQgKfHns6K0MieY9VyXAfv0u86Qy1Pm37qx8dS
t7NjceHFl2oorFpaJgDi0lzsZO4s4Hq8+IiBWcddzVqV2UPDZpslJ4PzOkQDukMUYUuEfqS/OXkz
hiaJHUuGQ77l/OxH6XZNr/YNxWZiKfJqPges0Uo5ocLLCarWkk9H8MKQE7DPE0PuDcFlgaGcD1R6
FyTwZtgqg1byQUyfot73l2gICCGDGspeGcV6yApYb/7KfafGWZ8C6CIwV5IgSC1sP3xrVh9DoKd2
GbaXKOD2cMOdzZTOxyEaSdCaxhFdn1OdlnlK/qt3EDgKFYQdvkaalyL3LauRjS6H7+fR5dPQYunx
aOvms6iztPRrYpHxygJYrRkP1rA/suRuJIAUjI+UUmdNhoYVPKQ/lZ95wdfoCqCJvYjO3r+WITB7
tU58SzJN4J1Zi1svzuAJhOe60ZyMqErvDEv6lWUy5BP6ScZogOsuQDITSB8GDT6+H2/FyYcPj0dU
31p8PVwQPsxYHGrtws0vQYRw7IqxJ4k6yZQ1q/qmeTB4hejT1jVao9UfeisUDe3pvw+KoRUrTm3q
SP97dVqDgFGRiySH4ipZ76Vb3QkVyFPDAe1UPBylETT6SZyGAfpvCpWs4r1OUGnPOkb3L/oFQk4u
MdK4bpSptzMUDdfSIcduF8dGMnIRMzVVcxEZ1N8wRXfHUMhyqUeBhS1sUMzYaAC0BdBIOQAaI1Sa
ySZGfwED5FeZYnFN/bzQT1jj3zDFapNpeZiQx6FOn4SkcsKy43ImZjSLaYY4bWs9fP9UePA8qGRh
RdCklNfVFUe73Lmt8RxF+oRipOuQhWSywSMWnuTnSe5IavwRv+hg/qvc7jWY4oJQX7de3s1fFL9Z
gNcdJuCfTm14OtNH3qgfH91faXpXaa3bKPc+KEtLj6kaK7NEZWX+9y88L/ZXhAxxz1UDaITQMWeb
MbhukJH4ZCl5Zelcm7EHTHo/UgzCujcnhcXZ6gcz/rJJp6HVH85a9gA25ORfjOP68zE8eGb1sRja
XZLzyzZKWieyEMOHtbkQeoyPmro7XnEhbuB13t1UNiu99hfLh9stIlgA2eqJJm+mUji/2N+C7pn8
7J5Z9UgTAY5umnlkpvHKILrw52Pu985+9NoKtBS+iNzn/6Y1JycWO0DgIW24a/DF8FvRSs/y3aEK
mYkQiI4SNbmLEUPCNowDE0+rpgRe/1tkOLzH627Hw3YH4JM0wUPQ+BvZz8FhidauIKQSEM0IDYad
nwpQblXXzVD8eZUatDV0XHONV5ibvU7CBQav3ZHJP1cg3pCDrg+OlhZlXvfT+yytdQp8BHkjfxua
3F9Ofpdh7/sZxZV55m70ZP6ZbEGuTOMcpM6wBMjkDxdQeBMURdCpKxGSdPAHCnpXRRer6Cjc+Hhq
tbAoIG790j4v2xA8G/C6SxloLMFfSiPE+cPlzoV+vNivTvHs5YSNzf0i+J+ijttAUIU+8hWiEMf2
t1ZWpLZEZkYbWQ1sPTsmfV5wtfXcvuQnSwhLBmfNo1e5ielfRYrfB/4BLJFYyjn+8GFlXDTGqe2O
WBjoSU8+8Rx4V3irh3yTnTp1FmSZTfDpAsZCeDCdDf6aWrQakZJZUmKsJkwva4iB6/5agIvo3lPn
ln01MxB/v63ieNZSnNlpqp94z+MkhxBeFlW4xogq5IgAHpwTQp9HgoX69BdAcUitir0Pwh0+p9ph
GnQiHhXv9qfNn6/OWqjvSrXIXXJ0hQSnCqqg+wWO304evZtZxwl0rU5SY79kUJrRnqzk6lntt9Wg
1bJT9U5Pb21wX29lj4b4OGYgODew3KKwc/gChDxGgktdjTH7YFe34sK6Qe4NhtLUDjmtbaMiOtQa
qNl/SCQtukWoHTGtFKpZtLEZLm/SjQwys5Jak8hubruI+tGcjRZEt/BxxJDKFeH5cYVMZex2D6de
yZWCEozYVH4x9fmvFHMWDDoHOrcj9nYo1+L3WSTvnNan9V5BWrd1Oe1b9IgW9mXfWQYTfASvh40T
ZNSxQn7dNSuT31WfBxOvesYkcA0SbNKxKXCDDK/ckrNv2efnytnzo6ZxMoZ61HmHmGoq82FSkos3
Pea5JM5BrxkYi4S4uwtlRBSfIE5u7eGIbzWfU9F+CJW45Xxer6P1gyBw4llZQabs8yMq8V7m9HHt
i5OrO+vNkXn7QZoZK+l9uNRr/CscAIyfwk7tgElJ7Eb5CtgA4VW4GK+yy/LRvJWWGjNWVZUp/d+D
f8yFp5BJyFqWpB+lapPqjsciLDaDZ2Nw4qZceaD6d6aOOLNvJaMmVDA8WcQvg2M8e9U4cYlkDTzE
oCMdHh+TVuTTt2uZIhQaTVR90WmztsMNhTqpBa9Z7pBotaWFhxGz4kR2XTHUQFgTfDrjy4Qfqd7S
FenFqBbhzK91OJ+/hNEFMgantdqURjX3fZ8zfusbm3RwHd6kJt6SiVwGezz+uC4IvyN3yt3t3f/a
cFW10a6qX3gATkn/k9jK/CLS5Amu3/0WPd52xFPKYfGN3FTDk0TnirZ23+FuGICXr+2yIAvJcwS6
DHHukDPlHxP6bvLACKulBW/ZGvhxgQ3eDpbC38/Ujik3f9TMshbAoYVD8819NCHUuVqD97lfXbqv
7QC7+oyQ6I8glGSgJzoZxV742rixa66YF+Gj3plJLAh4DFeFeNirxrFtCZRmwKiEX3HGS2qbC9vC
eycqmYrydLBZtxRbLuHdt8hWS2Ok3WJRCvkryw1aGCZBghgPOEpwj6jiQeT9M2fb4m75MCaQAnUq
JFpflcMxhwrvDip82LirRBZLTZmWQuHjtO5OcIlNCXYLa6Vxa1DyP9FJNT0sJfN3wg2rZM2sdXl0
s/0R7G4FP+S2vTrB15xwD/69/vdbbAAjCjiwJlg9BGdjzozG935S8k5G8wn9rVQeWjIeel/d6GXP
cml9foRQrbOOPD3cj6b+xNHQTyG0gZiOfsxJOGcbBZhS52TivCYBOfsymrswVVg+bPrFgzKDrjQC
NwRmtICgbywY4jAD8ToqZDR0BV3waRdXSdkNO9OvHz4yGf7SHAm4jD9gFjPD4uxPYFy0LCgDr/yE
pgZww4FEOPDj1CmnJHaBMN6begjRdvdjWJUAlYMjHpN+acXuQQ5UnKcOneUhe7Oku9F1WIkF2jjY
jTrJnZRy8oF0nA+tcb8a7InrPTSgEeMM5fyP1QPk7UzDPwl8Td+XdbU3rrvnwmDtF8UPRWU5sxl4
QM2D5BoDqK3HxBhZW0SkZIaBQR9o+Btq3H8R2pBiPVBtM6KloZeqzJnNEgp32TvLWg9mF37kjNPd
JyqJShsVVyJFfHt0SOOnB6cBn+SZCCZTrpvGID3D6g3fr5YRUWVqIl39h4lBO3QroL09CEQ8aYwW
xJqse/vRnmLdWjisd2kWSz9uOpnRHswVgDchXQJneSiemQLcqAMoSSI2/ObAssPWUdX7aSdrB/B3
50PrRxydm7wF2RgseBwWfMKFpYeIWnqC7Xxzq7z3v+NROTd6bxtnjJFH/0yvohhF8xmtfYAnG2P7
jQs8xRCjYJsPsWfEJ0fB7Hygl/hGPpUyfoIGga847uKiFtAz52OXpHWjmnX7WDMxwL9hFu7GkPSR
HJi26/BniCQ8kyrHgebF3OUvO8XL79mPn/T+HbA6BfJnrcNRCkNxS3J9I4832P145nzfluJCWWW4
jCTCGrVxlgz8sgDFp1YI0Ja7rYQZjvABW9bVv6MulDafymrJ4dbk0tabpz3az/uGhqRGvxInsjr3
Nd+LEPC4UH1C9omiDVPkWEnWgVXA8+jAQEsuJU3TmW/m95hPuw6mG4r0kJmzc6WyVPP99GtYGY0m
LRtf4RCsnMsYGrWwIfIrbucy6X26EkAe19eHhUgx81qJXU3C5wbXKHmIQDqmP5gYuW3vyFmzEW3S
PNLWEPtATJ/idWN2oZQW/aKgjUJeQYRJLjfx9psxlIsCj6p83ujxCEMn3q0CivQBfynGkAWnLR2z
vDZVMmCGbtEC/LGFdmttAeUW00x6fjNC8EBOr0+tzUdTQDoy65xLK41yHjhMWmWgPV/jrZCGM0EU
F4OqPagH4pKE2VTTqqm/ovmp7KwhCNKNDov33HoBu8gtYziH8TKjnZMdwNefePoDFp+wtBAl+pyM
vQQLBq/69jQmtwajhyYCIquRdA6YaG//l1Bh0l72Ygf2Bs3lkapRswhgYSdJCI3IwMcoVjoplTrs
27bLFyhBaZArz5JypmMXoy46ICJ3vXGcrlvvaJoY6tMg9SvLy9zRuDwiF7edWLS9dP6h9JwOGLzU
OIBc4MtX4uZXBfVqj+EEVGUTyiwqB7kIWN6Phz/W10+PCAfSp+CZqRJUFNVkOqztbFNgmyODkTeS
WbREBTjHJBQKliz58MVxftcFdLkbidYZaraDpeTC9ISCUPVMUgjDiFYvhXt9fymoIPUbOuat7dOW
rIwaNEjMIW9yZB6ljRfqAYEwunWWYGNL5AUCFNm6WO+LFjVRoejKGVMoW46snayTpy3pBxHrUbJ7
Mss7o0pmhA4GXU/ulPn0ifkX2Z7rYG0bPvh7EG3KP6GwIku8QmWhWTv74/1dauNs3y4dAtdNOGD8
Q2xXH6wKCtXFl7lixFszpF49SzYmGaVL1oavHNXyf6ql3BWSdQquJ48UcX4xUa8J1q6ooSykunIB
4ohSsHDdIIkJHdsfqfIflplG2OAmT+W4705Yq8sv/3jLiBR3QkmPGjnyMHM8t+7IT7wTp2XeXT4G
hcQK55RYb9WsmbksMRyW/ljD8CW1dyvLdQ8oGy8DpV9K4Bqdt9P8d0z8lFP+81Sr5VIhKBh3dm2G
To4CZMbrsoXUXg5RDFRUpItoAIbvP8p9lZ2fO342nJ/Moji2u1GD3cSjWHvRbpAs9jAfUQ5NYdeN
buo4PPeG6tsgEWsB4/ArfdBAI7w47CXuztRQ97DHvQjVLt382TLKrQO0Z50v0Mt96ND+XSuCUkq6
CgXxT7lHsj7icJhNXprItdOPvlWIfVG1Iwg7YSEuzayZ2iP2utLV/y+GP9iQrvABN25nXpZtmDkC
DbxMNwBI7MS1XP0HVl1UAohk0EAgBMuV0XPa0h/cY/m6k9ELsJzTMYZNaV2x8xxHppHnus+HtfHb
SjubFxuBLCAkYO63t54GmuL4AebbprT3QyKaPs4uei2w5XDJPXL/yawUBZyZBys5vqijZ9t6ltpp
ZhlRrYhaZtSbj7eMzzbgUKsbVoE/LAdQZQkshRybLzpSC3HsL4e/me/1FO/J5/2TT8bmzocV0imP
3ksuuvLx0fMWqZRAXOKZcgwGeGGBRao079i7Tkeh/lOcN4OXo+OViWt7MeIj4r68vghNjEmqXkd3
mayannO6EQSDNsSatMEasWCC+SBBr3W6G5LVaPQtOztUqYi5qVedb1CCU07yHZ0mZyAlqPe36ZSI
VFVPt9HziOguHd7RNTr1au23wjuK1h7WKwiRXw4SZIBictWK/mfaLurmEUTH4ckbKMNix2QNHQtQ
W4w1h6G5lrGjX/lhlWBNozhSBGPjhU/VHpc8PiZtxCFLRUaRtnWNMtxzDEnxIeBxcjxJIHWVjl5q
EJQnz7lSJeaP8f7dNEjUQpQ0GUdnXwFcjocd/gpogJyWqTD1lXdNfujP3CrVDbi0u93Nh8ao20FG
68HhfbMz0VUSd641nTMXIl7B8vZbtuMpj8OHHcbOGm1OgHa9p8aIyR/6D0sokEyQVUChAuDW7FMm
fM4lssQAh/PEEsIA+Ro5srLADesN//AWB8eVSFWr1rjUIUmpn9fbgXSAvQIlf+YBdyUeCVtTxz3D
nOcpw4jo7l2BmLpHyWDnIOudEJ98ZGjseILcHYVzUVmq52aFOaKLTn5gR2XwgE0BiPNVCVohCTNF
w71iSzY7hJXIUKie4IgExbUaATDCia++FVOyjauTTB/okBh7qgQZ2LVp3wbll96A/dcV+51ARBpZ
KK3+ZYJrBqk3fHYIrszshnb552Ldw8DByf2eiCkjTPdOLxWaAZznm6fFQZzOm6WAEFccpZhzyAOu
33WxaOHeOx7NjOvEz+2mNdtfkGGDvFUl9B4Eh2RINrG5G4MzoQT3NrabDaCQpH8oHF0MUmSR0qRv
I85UACLFdA9wexdsYbJMOVLqGO1o4aKjagKWQhIzZfaFvgEP/NLstMyHVLWqapul2SV7H2x2kfgr
RSyS1MIONPDX7VcKJXNtN4COT1r9x3y1vL49DaTJ7n6CRdqFZHhz8+3d4m9XAM1gOG0X+U7YG70t
ivMYwjpZrsf+PATjgSjw/tVCSeNmIY7kyayD7oXr3BKTQAHUSczIT4csz2Uc83sq3yZ2HAeohezt
8k1rn6pOKzahr/OYJwEevQTV21ZxaU/jWBSVz8IVgHgXfHNOOj81esxi6/81ivqR6XZCT/fVK5PW
Gg7g4p0nFbDeIs1ngvOzx0JUfTZZP+mZlNza9DBQ4/5jwYJZ/o5XNhDL1vWYJzQ1WuA1u3wyaAp/
LgiUWIuvwMcaf2Ln3DrpVBvqsQfn+uevGEnJzCLYvdCkxOcwbsWW6BkSLpAXkteQNpiZZfmuXeMg
VrSbZa/DdIEIgqVVNSrmr4hf+6p9yrWWMnsdpkDJHHnbcrmXw3eLDmOyGFHcLiyVp479PrBm8oJc
dtG2NL6nWgw/OXxdv90j7y5KLKsyTNe8gMGmyV6uc0uKEW0vnJzf0GsJ7GG77Ybbic6tM2/MZs49
EX9XaRejOHKo0X0E7rwY90hah0/DPq/KG0Cb1Ga0xKdIkjy/Jg7JLIFVNGsvsXzJd1hg1sw6+AcV
g1bCx0Jo3iTGL8GD6zzhro3yutbq5k7vjKzoib9IBskPf4tbARFutYjV7dq4dcVsfPY9maO8P7s9
Fj9EKmouLzNiOgglWThtVM74Q5v9RLoLR09TJH6KeR7G6rH+iXnqLfeKjWCwwppnOT5bGahkb7mR
qalK6lHmJ4Pini8fRsX13ElTQ9HEeT6zccMw5HDgPrpuV0dsEdmPGHVfzMnoG1rHVcFc9c8P0ix3
8x7aR2mKoLVBQVG6WxQ+rosHOPWcP3g/xzehLfE679BgU4P844Y3KoIP3NZPEouUSvBxCKcoUUcg
IQDRZSB3WWlTWiEqA36Dfwf8GC23xopx20Lp2H6cm5fiy1ujs9aN8Ag+lqZW4z185XAbBmNR/xrQ
nObSyLjHU7BQswo+2St0eFxR0cgJwQPNEaynFfSPHtnHDtYidio27zEJUNXVbVMe50cq3SQMXTMp
SX2B6xVCwJkiYPu7/ZOieMjhg7ASlWuNPzYWYzlkb8HlzzGjHFvzm6cKxIN7juyRJgQ4Kgirf95k
3MeRlPgKqvF4Fs/bgbHr9+omT8prDsiln5oskt67ZfuZL6Fe1euFBhWcFcb6ZcYRtlpXkEfq6m9I
PxoY2kmW3PIGITk6+5HnkI+11f7XYIRzdAtEyTR74yWRWEChVH922neE58LSFRTQU1hpQ+aqBXfM
iptbSv57p2MT9lp91qXg8GgF8TsK1eLUxlBehBBkse2HuWHwPP6+9pxjng2RMAbGrB+fLa/TR9oh
s9rY5ODWfWandWZuYjkskavABx/D68FfxWg++87+7LhUC6GAt1ziNjuJn5qKhV4D+99N+/yj+MYT
SRHfktNyxyacGlXRIGuHM8g5WWJE7FxKuoNGuaNgImfjY1j+3vz+q54sTzlmfy/3lgt9mwfVf+Go
SayjeLD/dF6Ou7hBsYOGyV1184iyLfF+7lQYbv6pibUI0N5ciO5nFPpVHHkIlOODh9w5j9Lo9Zl+
j8yu6PWUpPOYdfW8sm8RD9xwSkFiFbVcbLipoBNVcn56P82WobojCUypEBilCEPBSlRHyY58n+kn
A0144AhnVivsogP3JE2Nqul1E98EWAXTiGcTZXMNgh6I9MuvQ7lMh5T0BP6Dy9SuyymWfIicHpwy
3lEYoH0yzONvtYEDPE47ykcmyknG0Xi8o2t7mFfuYErvydg2x+sJnBE/FXSLs5JbfU5Qrf0n49Dl
88M/1ScDsJdID/lF0DEOLZjFmcHDY0uVDfMLvdyBX5OUxrvPEZpFpBbIDxQsEsRdyvZQ17CgtEP6
wiGgLJzq+Cib3rmVDiHLma7zSzfctjZDTBqVwrpYd/VILd49rmKS7WfU8863dv5xNzxmbLd3d4xs
lB5J69GW5FdQdyceL44H5zJBHrzQP4LJlA0+kbd00b5LbNLXqmgDjsYBWJxH7jdzq0AXbs7lKKkK
Tsb/UFxzj35bGlHQNlX/NwjXNvEnhSmfT2CYObYp3xb2zbW7o2BjZjn6ywESxVRSrowk120XQGst
zhjy4APkUJD29hJ794yRLo9IvrI5rSsBmiSD2YbB6GpZStCm8PdJTv9bRK6OKKJ8f59SdTKz2Fph
Jyz1xgEGAbBZOl1lFfMrbxdp564rcpaZJK/0/cdLfIU/cx4GqrCX27jHYlvEexLaXsL/E41cedwn
+KNxE79H+ni8eqQXaskYyiy9aU+SsJMy9YswxFPtbESl1LhzSLLs6UYwwZNMAOM2S3CJQTwZWvcn
ywG5ZeeEFmzh90xnyDp4cbv8tx0WTF0WUMwk6L05LiZTDGYIXmfRXmCbR8lKNJGVus1Ay/ELTL4l
V5zj7SJtOs/G8e+hFaRVVbUKGPmAE0xSSMubVwOpPj8CyT7E80boowpV/uNQZwdMQQtN6A+xDtrR
LU/Y0+2hbdFirISjcRA/WVH4avXU846f6Oiuw22nb7a0WpRMcTU5oo01hoqECmMdMNX9lyjT1m9O
bNA672iR0V4w/eqsSmbku2P5rqZFMvu1TPpKDfGIqtkHueD25OlmoUaMbW/ifJ2/bO8pZn9wpbRZ
2QGT0vgszxtB8uDV+itty0zxOrRi0cN01ydCJ82QmyXPOR3o7qNCvxSK/KCfnzC3STatHyVVyA78
xKMBAsOrht5hvbhSYSn+UYPw8xoomJmQBVy4J3heVlZD107H9HpNxNXS5yksUl8bCvhcUUTy6pb3
P5HjWxsBFL7HA7yHFWykxrCYS0WLyk3sfCI1xMv+KCFiaYJKEttmgyJl3OmRJiWJE1z4N3rRXHqH
mtt4fXSXwUbALEH6Ou8VxORIgLuAYYCA6/I3BQCb6zq5rva+AGoWLkJ5lTosw6I6rAVvA9NYkose
mZbyulP4lp+60ow7eJheo3KtH/cHEpwVk/cbJDfxlVxxLfl78pKHsew4oX7UMDdnb0UWQyemeEy8
ePDQ5JmnFxmQCjyg4KX/e7opcEY5zK4HULxyhyiHqY3FlQE8zTx2yEAfOmuVMhHt8GuEP2FjadtK
KviKRZScTIdSledyy+xDcwmn+BeDs1ZcZCq92qAk7yKpwWnCRiPcs+SyfNyxOM4GJKW29kvfzEl3
nUXQ6QYRLaBJ5U/8BxvLZ4j6BKw01TvZQBrXmtJhrT25B0hKGhIgrr3Px/tOdFgUAg+ArfuNpAdh
Pf/NWX1skFHbzqt9qAQEN/YNNJiUI5R4mHq1Etjd/Dfc2VcDrj44+xzP8zYCacz7Y4qwzPq+HctS
AfSM4KTMkeMLvvElKw16nmyoE3jU3+EdjMDuIVEa2FazsL4QpEVXeeALr7PwU0CVj+cuR571GIfq
UmkDpEFmXTrDhrVOorONzW00pvVIWP3yxVlHertu2JyDu5EpQMdlkbcBXAOUl29TwzfhMEpLruC5
AP/4BIZo9FD2/mKjCs9e60T0KZgaGP4D2pzxjTB8zMmmEGveWJ7gfmDk7GvMooRdLU2JfhNGPbY6
3Cg47if5ujeUydokq/HJCDkv4CfzyyIam2Guh1GShDowRgbMjCZG1IF4uswXvFumYx2RwI/kIEUN
z0sEh2MN+rUq4XNNllaAa9PjfUXDdPnXTUEoCZoH4J6ZuiHiiCdRl82xSENM8k+3/fcqLq4sB+vA
woBzcbWc6ycXmCtOdlqAq98+VW7cNj3IP6e8OkLXB1T8XV8nMU7dIIT6X0B7BeHWOdFRvGryWkw2
ggY80U9z2rg1s4GIt8v/7qgNn/9+56k2ylwdOaPz52HS9VihZhzu3kmVeYi0KChJ3xlI1IrQWODU
sx68SMfh3UosZrLNzOexbM25pmnspUlTbEWBiKZBneaqNwrglMMqWEGZdv3QJchNrmAneLgyAAof
uSy8CoNfExmlQAKtO+AKo7zeVq3cxie87cm7QuJRuV9tZdzj6dDhulTG09oKhZg7LSaW3vOVlnF5
AYZAlPENyNqJ5nkg34BpJlsFp+Yd24o+6Wdj+JRVhBzBbgrm0jkqunzq4Y0sMUnlX3TzLyDiIDgj
2pwQJlo+ahZXdSMIysALc3q/c7X7a+UkqrnrMfVii/NT/DUiY5PjKBcN5CpBRyjbJ9ACAeLz+1iz
5uBzCi6F0sKHo/yc4Ft+kaGx4v8dTRThWR548pgsyHUFCP/jSrkSw4w14iJnBqWFqChsxRMb39Ab
zuHI+A4aDIlRLMQlJhMFiJM5CfF/v+FkAco80NBjzbgFFjvb7UNuoXx7EVFZWcQltMMcT2RcoLas
kbtybQOprcxa2cerNbN1x/FEbU8/tDB8X+9h1uCl/w0y4C1b4f+EXDmIQSBtntoPg8PxOldzNt+Q
cKOxp0VIL7+9o+zIBxuvIcNTDNAmHf3mqIC5W582b4g8qRICpfB7xd3u42RT0tCmNKLxnISntSa+
lBD3kAsAaW4A9g9Wxjx532F+G6C1KFrG/GkS0+6MdscdzfBgIn3dv3KiNAf9+sMuVyf4eSY4MTkc
bAKid/1+P3P3mHb3k2dz3/yp4ZzPKb8JowMiK63YoQ8NqlBZY4AcZtV006xk6lHQdtb6plfMewPt
XFpf+gu1AbL9Xo4/EPl8heO5yNpntAQqeQrhvoDML+7hEzpAJfCC1ol6MJzFUXhaYydv4nLNu3zm
6+X0gJZvzDjczGgrGBUPyRqi9Wbb4fLP+duW9g3O+gr37HKSNm5vRl6/IWX/d4+G0J2nZRvZPXIv
sfYtRU7o6ex5CAXwUdv9blCc0LaJss0jLbMXtUKcXYusHi/5fDd2L4c3+u/lQgM0ox6qMidQITIS
P6ykDaAQN9jFDc/UZ0lx8NxF4zLSQ2B8Tzij6/48h7ESzzQUDOfiz9G4lVFTpHK5zws8oyByKOAs
Kre723zc12sx9tYf5ZEXp3nEp7bc9rfBZ6cMhmMEoKftjRINPHlhXG/BwyPFkquBuEgkmsu2kXYA
Q3l/8O3gGzcbSXlVoie7IorFXmaXr/Nywi6FViVDdafoIOHyBVsph1yYR1GHqdmjI6nY9Zi2eqU/
dmI+3UkuYDemrTW6ElWg+IP+L2qyCiybYPQmfApswdWRsoS3+Oa2G62X7XB9rKvsWXD4Yzl9Wa/n
n5x2hGS2/QypaA4c+trFHGVSz7BH1KocHHVenWBeir90rSUKloJqb58dG1wYKW5hgGask7QQnTGG
agHe/n5Cz0W53LizBC0fHtnTy3/Hr5X4E9+sPn8ToTdd3R3YUhmcEAy6EEMRfTpQVYF1PCHxvtZY
kw1dAVr94sCyFdhXAEIFXBKxhhGTGi2UEIofdO0ScOJN9OZ++ucHrcyAdw0sqH9vY4vvMb+rZlRX
Slt67x8Kv4kh01Zf0LhUbn72uv163GcMAVzd4YrZBS5EP12U4Yhs2qUmqW2ZCprqx4jeRGXM6B/s
IvluD3zwAo/D19C3CW6lGOQDv1hyMcZTJwHg41w3B5nPshuJCfzSkQcVdibtuh2sBdnT98DCRfTb
LJHv8T2aiMehk3irxYpwF2MKOHaRM4WDwcfeJvJj/cyZgNE2iDNGxHO8FEk5691C7GKsHeBG2EOp
5sxfttcr1IR8pfSG2pE2vS/zjsCyQzkCNrFY9eRZhPxgfCH5W3WQexb0UrDAs/vR2aJBXYg994eg
BjrO/UzIfOlmvuUcNt1oicadvDvBJaRrMEoG57GfLHipOOEnM6+oQRER+r49OmohzfqF7YuFD6RS
ounkEmY0Jt1HdY7GwV3GKk8M4FgIkSysObZuWNYWuoypOZbVlfXwLVguGnQJMwC7otisqyp27Nc6
JeqxKhzEpYuYDXrSVwDD0S/anJMsGJyz0U/dQeyoleYm8cIUmez6Up2FE22AX/+OFrJp9jmTyCNg
R9nTvLx8ypIng+hrKL0vJ7KZBJWtpD0EdPdHGij2/BHzPLtIBdjCndpfIfve8mnUZ25WlRxKI2JX
zh3WK1UGSlFb2HWsO/REP3EP6Gn8uILK1cVtksWqvle51YHpCQzRgceHyTyAuysNe3Dy7zFDjnqM
GdRB5w3G3CxtwUou4HUxt0/cgEatjmrE//bSs4r8Cvb4xt+yxMf1y0BPt/ckBQZdlsRSyjnE+w/w
/PKnadEi9MG7H2rzmmwKvXMUa1GEk5ZTtKP9taxIRS0xn7o6TJzaD8PFmeNynjQQr/cLyeI7IZv9
mRz4NRcy0DeZgdLbOzPatjWRvI7c+C/W7QeaCQFWKLe1rKoA+OCjPm1hwpyumbeSlKeQYdExA+Pj
Z0WbtL7n7rXG+7SpY2diNQl4Gq1tUvT8oNgrCTwodzu58qd10wX0r3mbQR0FGGPAVwsZ079SNCir
P5d3Wt9poif+gR+3Y/JpuSIPamhYsAfmR8KKz3xx1dhI/ZVNoUc4AIkuE5W8zlOYoAola5wA9aq0
V45OIuotUNwdVr3KtBfPLI7YUCE3E8xSROTJL/kQlzAjuEYOXRWqB3JLzhMtm98qjPvz/kBZBxjj
NdL/VV0ssePeKh6IHs/3qXC7ly010s69CQDdU5ffAX2waxk/6n3Q5GDJIPJMhBV9FU2RkFfetHn9
mPCcuFWqRXr9WzaCLJ8x3MgLOtIlFPDZltYCmxOGzmksp0giHvXYz9MDxqTe/W/GP6GjijOShaZd
N1GyDB9adnxL30/W2g4fdEcpEWfzMHBrF7FnggNVLBE0bSSvymwE+a0kmQzP1om3zSM+oTvAJerI
nUkLPF1hs3wDOO9/aiZ9zDiT9jdgq+HZwfUNGpcdh9+kjG2qQNNHhAk/JiIPMYXQ+Q+QnRViXLJC
3tq2YxPZdC4HXh81NHGf99//k8wc5G1UEpOhphFi5jraLRy5/LcNhQaIHe1mQ2yAVl+4id0XviqH
cRMoCw/ErYq5KEZ1JGvwYg+C9zx67nu6QGhVi0jziplj3xMtP0vhjHlISUzSpSuPV9SfHzEAA0RD
9EPT1KlCRGxa1PbHsNdcsE4qYSXH69cSNboq4JRr93WEvJ2qNH5yz2pVoqgSgxoc5F4ezXrDoL++
nbbjzk7ud8ZNKh8l6DUSqogcPk1hat1ImV23xrgHFBgmbuB9zQB2r0qi1nQmlraVZDJAiHrhyy0+
HSNWpJqXmIYbeLYXBzFdQJ8SpAd74WX3nuLqSiGd8nCKMW811INo/dkD2VlDsQi9aMbckxQTtlPy
2ZxXAD8+hHKJclYYb2zVRVzNuZgTKE6txVqopTWqTi1GT8jEykBH+EKY/l6eKvnVzWj8LWHaZxaM
QbDR0XpvVtr3VJTKrI95algaNG8RZVkhzCxjm2YQMVEUpILQsN10PcbmIEymdLJoL+/DH3ByVf38
gG9D87hWnEQNkQ4vIDZmr9v7/FSb5pqiW8pCuTwyxsks45UAPQnaAx+yzRKvWxYE0kQ34GPdsz5w
Lc4rQPHzEGy3Qyu8HOLnmH2iWTY3Pu4kjjQYZfqQfEp7Fk2VsJ5hB6q2d1TSyu1LxfgXfE6m8CKD
fRSlDDoOLsxY/Qf1y0AASTES/HCKIiz9l2sULpwF2Bs5VsJPkTcSDm7uxft72iPSXfIN+ZtQPQes
nxL30fZjs4B0BHhI3X0drcRkzSIvDJbzRdt27xqCqkiiv/8OC5Ux94IZCTeT3ZPDV9I5XxaMOQhV
tTIohSGiCwrcM5aLwnxLCOyeVYnzLHIvdSVjcz7U1lCeXV4AbWVvSQk/j0EAAaQ4t/Dh7ZbnHDt+
G0GU4dx15XYSoHuodo9dCYzYyUmyhB5SjDJ7HiaCjoq5+b9R6IQplnRve1qMAE5hYSk+4lhgwCqu
Pqe8MxrsphKDpuwksry/qut2PnQ4xbV6hc1/TzfKKu1mIPkSdWrl/LKDx/Q6P9jHyTb4U0guC9kK
caBAMF43C+XtzdTxL+Z5Y4Ys8bVLMRmxUzklAuyiv/d4gcDQuzT8fPDuin5jIOoXfY+OqmotzwR7
M2vWs0oUVpT4OCH+uk2VPcfCvuADDwB34QUxcrmX+lMeFfQbCjwfmk6DmEOIDQ/uyKNi5pfTMStF
ssnQv/hUzwWfKH+zFZW1rdsdHPMCKmJWL6CSoakCfPdnaW74/kqdLPpzR9Hx40V+vL01txfqw1v2
Aw/rGhw1O6MsZ4M08OKPURcE4WgcPqKr5hdVWRNFhmnhXtdZMgt/IP1IHJ8Q+l7THc/stp55Ohd5
0xZmvHKz9JtBdj5Mqh03YM6xE3Igb+ktcQXuDx5MyImL8E+mukpWxXpKGb9juXJsZJuaeYaxilE2
H6Ac0LTXi3m5rUw7CbbMzNXvzoagSjgZq4GHt/W8a2ve8QwOyLFGbcSWIu+MeEjMYrPl6tzzqj8T
P4sggdNmA/K+h2ayTdaOt3H29iT3nmPPPT51Xwaea8LB6p5p99w45uujR6p3XdGbbAZ3PaFYls+a
gDlUEnhSEUMHgjZayvqOscULVWb5GMc11XdDjZxA6MYH0fhfoeptMGO8y2+o6jSJBGNRaqNYzQbN
0/13A7gdMnjUsejSjIekkphp++3sPnq8RitdNALhNPcsKULGPO3WGt5cYxisqbIk2wV39WFWi1zb
mhwDzYMSsY0Bw3hQGrUkGymAusvkR6hH4loAJ9yIL3Z2hypvLJP/PI16fak9GNcCqw8AFGqitl4v
C69rFeqce388bG/YskeFxhTDMjXZ9ePhOB1z8DlpxuOERmDliqyLyiIydzCcCCkHOFnMXL8Mtkel
O1oJwd2BRDS4woJz8ejOOBd4qmnTvd0WeL4c805PLSYtLRoTpK81UdqvuqMTDqI0Qk/A6bx41hw6
cF9Xr9qmFPFYIyGVOnAA0vQPphWeJOuxHRZwZbD26viTHfltAiwqUutcx+gJUwt3n4l7pvEs7fLs
ODA4OJx3T9UcOfNsprAC1hKbX51cD8eQMB+j9rib0JcK6HX6mo8BgDcLV1kjFnq2leg8DNT1hfbx
7i6bd9d1iOpK23ASlYUtqWHZwsglet+DJ6cWDqYHBigrhPD5higE1LbvGD5XIGeGq4Y2eq8LDYzx
YInPEgzu28spAjdQrpIkrkqiJm2G53jWhVOFSPVT5Xu+A/9XFkAwhRyGsnKCNXQz3S6OZMxstbkb
P3/crdKu94THLWRCwAtGsGCE+KMEC4wJXgYtBuc5FVsCQgH02DdjfZQ5COOPWH95FkC5CoRvHWrt
2VIg0nhoW0jq1kInfSl8ThDKqOiYwJK6mdU9Y9up34sdYVg3g/f6KqqQnZFdyxwINPVFbdYQOc6S
KcwsNiRlHu3wss/dMVZ9AAb0wAVRipL53had2pB8pmf4UYV3jMvKNazlYl52MSXrlFgTQXZ32aOA
cjddhPB36DSonvBzZgk/Jxmqw6v75ut5Bryo8k41IdHTNLhUrFWyy28G1Wa8ijNdwX6N4xUJTrwH
kop2FtoXDVBXgi/MKKnXpjGGvA864I3IhN73BzlwP1o424yTITZ0ffNYhGAVRxleB+dyr7DCKg3e
Q56EOVOCQOivIpPBQVUACkzLmnbEip4bPYB45GILi5LM4P9XtWdUbU8l/i7o4rKFie2rfUL375fJ
hLCQU1EnNuXdAImn+ckuuC2zXZbmyPOJX3bikr77OFmGmLd5J1wFZAX6qPj+0CJMnQc6Vb2HTbKJ
ZTRQ77nummf2clV7WytRcVIpQV9yiUGA4RrV0Tm60tMmfz9Gbc3m7NJ5yR9AX12k3r/tmnaiLO0M
hpcHOZIYAw048703KYSomCPTYcwXEUPXne4mTNqvBx2uVuKS1ZSgH8ZEASm1xCZmUuLcUi913jxi
IFeB0L9Oje3NoAmMgWufCCTyLG2pXyHzld6XEsZpCCpi/GBY4d4P6XPuu+T72aCzRMD9q1NadoKb
/1MbLfLl5/+EyvsNZhknfy9kqCl7e8UwOjycBZ1BDyHv7V+CXRdFuqL3SXJBeh15Gbhxb67R29Im
t/0JKC/BXWB7WGGCf9hYZyAJG+uDxOB/jEt2wHvNigqUrlG0zA88mmTki1vREF5ndDu2ca3uSbUb
2CNBXYM1hwcP4EQqdrZL534KyIZrevmGpa0TNJfdtL6HftkgL3kzHqNJjoG0mx0jSt+LmBUUqcr0
/R18KXEeZg81lJDOAhFqzAnWkHzuWKySXYcfbjrObQ1rghWWr0aBAoTTd2gNisEe56DL+QEp/0Or
L+TYpz7D4HeLl2MUpnmNkbl93B8QUFT6lRAH6bJZV0/+9V4AjMEnrqWxNT0G6ke9xzpdpLb/60yO
a5ocM4cRk9NuZ0sg9QK/EgccgrVT1Nhprc63+YGOZ9lLHl3v+7hz6b1jZWBARtb3mQ4sBFRgGSZn
dS6gEzS8u0dSWCXqip40XKi0EZzpjHt53bUIJhWkHlLn6IFd+9r6iT31izyJX7yUNbBHAnLjrErv
BC+vSjeT2Cm9LXiKLN9K0+nybOlWtTNDwR2pz2Mh1vxm9bAouUpXQtl3NjzZjo+4D0Baqu2yCqP/
DLqRrzgfDQUSIwNCuUdNqyC+26whj86Z0WrgOwU3f1A75PHlmN9D/juEJ01kSz12pCg17mSFlt0m
2cJ+px4DZETMJmVLxn6aX1Y0yPv/3vXek9UL7rgdv9QpCT4nqgJfRSQn/p16Ct0Je4puI+EtClfd
SBmLiMn0Pszuo/3KMRBU9OGWEXqrrx+kjYbz+h57vgGcsIJ5QNxUKKC2EupMOZX5T6wEDBNq0vMe
XYgGUY0J7JbXfi0Mqxf0iFoZ9TofEjiH4zQjMnIVX5/vfrd2Epe/vowBxxhjP9Mme434gwyoe0FS
doU4RIvGELFBxuhitvK5dyAaf5kGA0c1wZiWKjfA2LZjGgDA6SfvNSFOZFDYPMTI1N6TYP9amGAg
ZdJV2jREKNEGrwYilFQ2+ZK0rNO+iH17cuRhtAqbmQfNYDUjUEaW5RNTGy9O3gaOy8euMlf6jGC2
DXner4ndvoVt0dotkgP6qAKdePC+lbZZgcrgdJQ1/GMPQMLWhpOSAzSgH2lVscZyd4ELpNMevVHP
MQqo0NwLsnB8FLcpIevYLPK/lZIaJI/vQDULPnvuZsqRT31piTdZJ9626E1HOqFcMGvcwY3Lt1SK
if8kgCRFcF4xg0+mT1G9RVJVZvLtRrwsLxpMaIMy/g/rerngzzIrGWtldQcR9ZDxAG73OL+r7bps
ooH/Mn0ITH3dz9BsSlSU3XdHA4ae6zIXNvCDKRWKNpMiULqxLVvnavL4P/qjuWqWmVNYMCs3U3XQ
wzjTumuSZEj9fZpM6R/r+a0Zh86LSb7c14bh+ApK17iC8cWiPDihmBcngbAJwD7XoGsXLI/GXReg
5qT2AVd9hDWvO0qJNcly0rc4FqOhICfuOCPR4EFj4erDWDOTXKqBsjuzy1B53fd84+8xni5shv4t
wz2pUmO6n9ymDKx5mrtP06S6T7/mnv24LGwbXmM3gd8xfotlz/remvdLMNo5bcwIVFNvhwJbQXUH
O9DWYBZ6JgojW+vSlkI1GDwTDGzxhSTbgR8eTo6OmgatczFEytgU3nEPuQOzvJgxyPTKaFEeZ2fX
d0mwuCw8Y4I3aiCxiL5LhoOLevVNaCu7JBbOyFVJgu14wF0ZsD3A5BK/649iEeB72Oc0oxBXIawK
Sn9q1WVhmYA+kDrr3Wz55ZdC/+wvL06IYoHuNO7+rW0im51DMN3wmxWVRlMj/39txBopVMLpx3+t
1STz+k3r7XcJQDg2w/Tdlos1efULVAT6JyrDDzhWPV5qponCRzks9qX55Wk3Clyhy45EzbrXw4h8
DrNph9d66X70KWbmfVmbFhqnU2f8OHrOribq/YNL9O1yd7B3u73z1kbk3+DUiwR+T7p3cng69BZ3
lKloOrgJFjxIfEey58SCqg+roS/uus56xUUJlZ9/5SDpotnbNSgTSChqljGxf2c+Uli1vFTaSCdy
OfLVjkn7gwvN1bC+cKDdnq4pevm7Fd2GXcjRo9Oow3VePCVDSi1R9NYC0JF4VW2vm4FTFyNNDIP6
xlDStWW+Fl5X0oTvJui0eviWNFQvoToBxzKqs8X0edBdPTrXDhDMA41GfMuBtp4Qy9a35M5ijXns
k8Mlz/hsNNOauhQVCigHmsAHFG4O/mhBC1ceoKkNtW0fl/Uu6R3mtjlCxz7jMsNi/aITlTzPZVUR
4CloQ9a4XJ/kf0emec2uw4HCK/o6iSTd5Bon8hDTmdLfYfbIGCjgOaXUAUg9IrcDhi/SkJpdF6aT
u+Kd6PrGzgVc+ZOESs54OP34Wg4M3OEvn8abWLuNv5Vp0u8MawOBCtXQk6RLpYHvZ63PfKO5mDel
ittPYCH4EAziOs1qpq97R4SDzkGzFall6AUO8UslA86aBnODoyMcKuZsbMcDRFSjehHfjz6pBeBt
nEZ6vtK88/XTwo2Yo0PBbYaaJX1qtnBBCTUTkPrCHqrXz0gDS67mbP1MiyaJtKcaCmL+ba2lNBAY
lB8wtP40aBqrHUR30eDHnyno971U19Pph0m2brp8xLEPNLsrScd45+LjEzPkhksOiHav8/GVODTf
78fzHwCgx9cRur752b3c8qBKWln6ley+DGOVpRCcya5IRKIma6LAFx093Z3B6phQEw7oqzFTDehy
uUSYQroXhE56JZZB8Fmm0HvbRRqiyV5YwjiGFw3hth/4JJCyKkF7vPztkqn+y+P/m9HGGnpUifbr
OMsFVAUMBTl58i3cvAGB+/OdH99ztBfX8JZP1qZpR3CSE7/GLkJ+2H94f0YzsJUawi+gz3+gpwcV
D39ycfOt8zdj8Jql8IBAOLFE9TvRjGgUIsVYxh78uII7njujKe+hjdofmroSZdDbaVR2mIjusy+M
iwpqchzRWxpLrRINhZLbflYiZkCgIHnWiHui6JmHl0hs45JklycechKXt0WkK0Y7f/d22IeysITB
A5jCptRMJC6lz1Wk1S9WLCL4Hi7AHMuWk2DjO8AgsMrgAABgG2UseTFxhcgjaup6MxlIq2LHxXE3
T87+as8h2mBfOXluBFYniVkcwDHkitNbeIS8f//EThF3Lh4THd8ZOLJ9k6n4N+cFVolzdU2IAKTP
vXx2hQWLuBVItIyB606xKn/uvum2BInbXrhXI+ye3+JpnY1a7ZkGhAdP+1brv1CjQoCjyNRGpLqz
8BBTbZmtSo5cAefjoK+ulaahbzlsU+t1n7oseRCtRzd3yWBhZHC8leN9REvM4W8d8DHOc68F7S2/
6+2hJFC7i+OlS/66H6UNaA9vwym/8aZr2UMv39xlMwoGiCZrJedaQLNnjHsFR0pjcLvkChmwI/Mo
LAkt2xO2wjsf5DE8Y4yqkDS/n97pTcvmsCZgNcqFJv6bN/bzmvD5ZL95JY91KCaARIMPi8e3ZmQn
LYlQxeIOlAmOjVj4GnDBFLHqVql1F6m9zDgtYtBFvxmvphVDJzpk5aPtXKd1INPt2HJeoO6up+MO
AOsd0FWSVUYLCfplJJ2rGbUBVR13566iZzWSjBcLjgbas+xZE0ff0OSpIPNvrXAHnLSYPnqlW6t/
BEtKeo/cuD9DcAqDDXyE5R2cxbiWlLUNURl4Se4f5nYnBBtXVTXh7+zNSWnjxWwiuWyNKoNrFxt2
AlfVWULveSiWWpaWhVlskOyN4QlOOaGmSkQX4BAifh/pShQTFwTDsV7I+t4pNg5nwOBjgZhQHWw9
x7BsBOoi0rcZSPn9kfhfL0ydnEebKFZC7GsCVrDfn1XQGmqhj7DhB9hN/WNq0k1I8TAxBFH67lpZ
8M69Qn4gBhRatoN64wT4/tQL851j4mulGjRQmTECeK5mBmFoS3HtQ5+w3fz2U+Deyu9wrHmPEHJh
fNHWM/FZKCEaS4X9Cvw71I7MgLou7pGIvW3XNTGmWhjyRAnEHFc+aDMwqpMhVaLE+fu36A5aLFk7
+bwFt51IWLZtxaTANqEIwxjqQM7X7jZK09NSy1nMNqfKC2dVHNRO2lD3nfOjXrZ4kOrfMm3dzINb
bCpQOD5uI66MBQ6VQfFGzaOg2ZjALAupPbbxLCWNCZceNyCln2VkCr1VrwCiJMNiJAurMcQbb8FO
lpgal0pMCWKk1YQwgeceI+iudzcxNvMYVA25Zm5k0XT7VKGTgmbdSe6BxZvFyqql0lzQitfCaZPU
a3DTrhswH40lbFb7ylGaBJ/CangFMaHnNsT2LNB0WvR03vegdfO58aUreOUDdIAi6B6QAZ81G2/H
c5MMH52MquZ9jZfGK3BqWkJhcBvBmn/IEMXZHwn+IA/k1/QeCOhD09vEl1cVl3WvfdPPomCd9CBQ
tZzzchLOJo3y9VLVEE5yrCNaQ4nIYYSph1ezhY2rGBjzaDXB5O2mvraG5bEtK6PAhCO4V7TPwE/v
Lzf4C1gtWR5uzvzZl6SPgY/E4yC/roAa/NV7nz8POREQ7zpoLQOTa406SJyKjcuZy1gS8Wpz8yFl
j25Cvt5B73YOM33m1Pd6UIElM91sPscQV50oam/blPmezsgUa3lm3FuAscLwFNGzoMNkJsjmhUMh
buPBEfIaaZHWbstvXst6BiMzZ48C8mGEZVni1h4lkYqIwFly17OXtmoICZNu9FbywLVsIBJzmG3u
ct0QFQoYq/IYjws0BVP8ByVWBkVWmjuKsO8xdztDOx8be9LzFJJXG6uCMCLHgF3vb8DUojUoTLTV
3L+ydlWtAsZx0h6G4pDrg49WwEpdj5bvZtSSeagx/yq/iHT1+mL42O+Q+l8IVWJjFNNvMiiHx6D9
nWE9YSWtp/s1PFgtrvT11e+R8QbHB3h1wq1MNfr4Va2MEF+qFsvsoBVrIUvQBnCnUbv332iN7lxT
DOdwUwCBytL4osJpAzq6LtQV06NZUmWUxPlqH366B2asO7Dbd6nxFX7ofWDwzNQBWRKNJdhFRu9d
Mm9CmawNvH7FvX2NVNkhQu0yjgIZsAhCUywpyvHBOVWpXnqPeiMhzGFwP887LKnfTkvJpVS8jG1w
yTeoGoGd/wk6G8joFuNI1RsUoC20fWpBCmDvn8kfMjLahM7x2f6eBcx87tN6xUQJjRwgUarR0stG
jwPUfQgOPm9Y+EkXPexftb4u4nqPIlktlYLEjhk4pNXhEKNj/fbyHh2b9195z40goEOlr6GW4h6D
m7ghD1HapDMIAe2Uxd+kGGDkntEMw4m9HLivUv4HVDwv0q/o1Jwz/TqRp0O7UyyfGQ4m9F73yXZ1
6j5++p4lMlzWNOXdDIH9nGPl7AGeIIYWKOmpBixkzaHyzGD0s6CXGgn2b1moiL5D/33Al4kyfLcy
BV2VzduxC1kjkiuTon2JddNZ88IOpTGAsLwlrmpIdqVNMPTqejOKPCiM6N6FUkVpFrkhCxn4awFu
OfNcU0R4J7Tbj7dYNpjrfExJJtbi6vjwhF5MQqMP45L/Zc3UZcSRMSuDsB0wtsmaUOkGSFU5Xb68
tqw3DQupy6aZoefVIlXGGNC/Nky6+WwzyxUOQjdWt8SgzhMNYK/gbwSVTMivxtfZ+SWN3FIYvAxx
fXHOxV8ESvqKWmTcCn577yQzDepfG1a2rjSyvDtw7ydtwYjgsXlGDIDQAcZAmArVYT2nYTeeVOEr
iUoaVK4Vwaz2puX9vHG/v8pBKbWBV6dmg06FtTiCf0jLk7/6ayjPv9E/tzFPiUleG7uh3r4kph8Y
Tz8CZgtrvVFHZbKpj6cDXrxDjtx/6CdghYh8uSObqv6sHRX424+91h5jCutd8eucisA4VhUTlitZ
SjiL8EI3V5veyuXeYVDWpnAs5oSKBjDxJKfg3BLNY3TvixUrsjiidA09T2AD91++uuBdDKDTvRIA
f0IPyWaSntalHmL3a4TlYDN4UFvbJDaDLFa64RpwqZMbF6ypOLBAze9RUaWz+TkJWXprThfAqFDX
oDu48xYO/+u0n5f/u4/hCOX5SPQwvzQVCu8ypww2WEhiVf4sSVPEq6tbk+VC/O/0gfQTAkBvRroq
+xwpqi3k1KiVtlkXJud+avXexV4ve/jAmt3L/s3jbBw4tw5fNIk0+GwAVuKVYm3yPT60KetanAXP
zndeLVwQiSsOwpiXR4C3PiHMPRmEPGEzIHHTqcZ8wjKb1NujjljXgw5AK4mWDmnq2T/JyLphg3fv
EW2Fs+VWj1hHbRj/PNMugJ0IQb3kVDByTzDXn3Nm/qVRvTHQWAz+HlHmtXyZ3YInG/Ga18MbL0NS
65OL1+Emo023x7cbK4CN34jQaYY3WRgnvMYA6BoiOFNI/F+0OxvwrBtCG73JXkI8h9FSrU00zrPV
L2IQzhMu8y5NnzjLKwDfbkiOtAYUuIRaIwHADBAk/zBwWuUunNz2rRlRrhIcb1Kasx9g1rvDUURS
ZCkvolAh4rw+DyQUmQnHG3qMhEFJRRnmukE7jU2aAcLx3amZVPnHIyGZGkgorUuEP8t8nTYcmJh9
P3SsESKLRaCd6g6QW10oplQrMwZnsfjCnjzc4vetLtG40YX7VmOnFir1JmpDiQNfqlf9/t3eExns
SeFYT2xCCexqMsViH0uJ6cjRkmVUGvc+Cn9Ps3cK4NiyziPthAfpCpnLtJTfRIpeBFRP3x/r01sv
Ivh1BZlHRx5WwPA6n/d7Hojf6ApGprizF1Z1MSwhezZrB9SiARgWejbH1Ul05b9mCiY+Y2h7xlGd
gbzd5gjzDlOmiy7Mov3y8ZsR9g/OnZxE0KVYGqMH1MqWfjokEg1azuZDs60JFt2bGJW0t4+9jDyX
fDe3iqH8kI1+AqImO8qBMcuX1VRC+Ui0Xw9uQmE5JPLs2iHqQsx1JCrdheNvRRr9Gv+KvnS8bEhX
V0iGyHYkbE2cXUZ7COMYV3zNMo8RDIQ0nf/wKJW/z9fVWZ4yXbOl6V4ucEp2naPMV6BollwzmcTz
H38h3uVJlTcu4Q4yZmu21LUTz5Z//Av20Qfkz4rZWlv1jShsBjmGEaX1cyy7tMrDvipez7WamRH5
UeTeM1JZgy6REAUhLWW6jc/a2Mz7NstU3XxbfaxIg2f4u6Ej8ZT/KWB9Bjew0ZNhEVjDnlzBQ4Rp
dGPD4SKeXz53kxtzymv2jGhSsINANBjyOj0JzSR1gVVFfFFZmlCZCK8p8HR134CoEeYnDAQrr2fx
it0ohE9c/9cd6L8g/agtOil4uZzVnfkM+pPVihsjI6arS9PHs670C4uCH2Yhi870kDr31ojkEec6
xNnxY2zIMCJtRUfjs5HccYyBDUiizywvqefmN7H0xvF8RdJ8ZTWgdHKlJlKHbSyPkkcaPgshMjLI
FYAZ8HVDxI1KIRPQDt17kGre5hMc4VP8BpzKw/kXYeNrpPYTIyu5DDGDt+tTgA8szLLDuoPXb1sS
H8AV8+y7qwBb3yDHll7HFx9PaVPeNpK+IM2pKrFdxRMdM6Xe73nlESKZUkKatSIsH4oF7yypzrHS
9P/yqGTkZtQz9nVEMR1eg+By7KOz9Ml4A0jtWUeH3GW7hgKn7MywyofB5Wqm12Kfup/GsZyNrsjq
0Xc8c+rd52Q3z8f4p6bvPgQvg50jFvMT3RMBbMMckQLVto7waodv8ydBSkbdm7mdJytpK1wnlHp+
F0wZv93HIENSYKxiIY1lJq4jyDn84hafPgTcb5sdENaXlCVCTspNB3hSTHccKThyl7Rx8zTcz705
+DFg/MH3OWodSaGTMs5LGCFS1k+HWw07y8/lgErTO1+yE+KUdroijYjfIu5oZbTPF+Pl0+z4nb9i
Xs3dfGmxz/NHARWNYAbD6FhR5/X5F4dxm3FhAZNQt0JYrbJKwwRneA8bz1i9lAHS2xH4OoLlgiDD
XNBARm5KTwH9HO9a0tOjRKj5p8VpqqlvzLBhWahKnCXoaQlEHlABJA1EN1V9utD/lQ6idhs+ReOB
hDpRfTFS78IhP0EwAf6dJBrsbbZfFU0WtW51scM9RnO1kjDZ6iFtLPvOMSgdnCMIdA3dciN/QOKe
DOq0RKQSkiLPEQQqqmqTPu5GYvzsD7nud4efiyCYZP/nJbY0xR86bkGp74nnJHma3J0409aWL87w
cS3tmL3fFPXwxAhc/DtgLXiYG12GGQ6Dwqp3GCrVGgihtYdMNcKwDE1zkm7APcFC7RRhWwrYldhK
FlRm19HeVAPoWTLstng+wOg0vlZa7vjuZULVAcQSqleaP6S4576waIuDsJwn5Zgxwh/m4lpOu4gh
L70B3gXwv1QC9bAryb/dAiLkdBmO78n4P5tGeexRl6L42n5VP0842ppqPqHKIzrK8RF4tWRt3B2e
b6XXGeWfZXmapYQPaWrfjFAm2g0k1ih/dFfj+38RGAIgBFzPLyMOcV6HxSr22bDRIOnQo9udKo9Y
i0EHP4FvmV00IUa8FHB54EeiVBC+FYxslmIbWdlmdTfHBZ4XRQZDK7LXeDTf9FOpNUiY3SDA5oZ/
7e8+gEbEFWvOCZggHsZ0H9/KrTP/QMV8bmSffK1m9jocpAqiPN9rKg8dBoU8tEf7Db/iTzoiQa8j
VEl7tEvC39DC6D9uhODRpMH0RkMtD2zRrBDaDmXQqEsf6M4+7VkmASopa2f7/GRfRl60W8+OnjZL
t5MmGwK0sPk0Te52ymLPH1nyINe3iu0pZq5AM/zLKGSp3K8O9/v9fgrP42xzPBdYzu8qTglTmwNp
yGZ8Xu1j2SiU62bakIkbZz07ue//W02G87D779Ym+CsdHFy/iLvcfLZ7zXGuCHoPw8fLRHV9CbTc
4jeRqBGGe4kmhxy68tdv1jDeeyQ5dREn/ooABhbHW4GPWJ0WVjMCrwecD/3GgFCstEpTTGzwA9rX
QshLZpbdZ44XZRGtMubHhJ3NSFygRAAtaxEJAHbycLzOZhpI5efHXVwdM7muzfikmcyRI5lNEgCN
86nL5l29Oo2HDoadjIsw3RhQA7PcP6tJLKoxvaaFwKnBzS0vqekW5qXH7nZnO31tPaDp43qh5itR
riW3xUeUfxcRX9sluI5mIlN1h1l9WQjx3UiIN/PA1s9EKzG8JxTqZUrlF0PEQKOqBwolk8NJvpH/
FRSzzcCgOCztc5qtV3vo6+lGpozZLjZM3bwI0SH1CPUptFrMYxjOCD2LWTFgKg5kyuuTizhazVRq
KFjp6x8b8/aWtkvS7WGIhS+iNyjKBbyH2DBhuMOcVNDgGvbetMt/hX8Mt0tkFU4DWMdwaXumL6J0
y1E6LId9qW569/HF/bL2Sp5JQY+X26KAtz9Y5AcXwqDuJI/gA7ZT2m++BN7wPEproYApN0nmJCmg
zb1eo6WAhjiRgtFjG6Zu1bXhfLmtkIs0w8WqQ9GUCSJOmKNbcsghQRBR5iGifjquGBLzexkyObtS
+AtU8IfpSY+zDG8ChuyToyZDweRll69/URcnNcAECvD4gUDX1RxFYzxF6LUztgHJrRpQhwFZEnc8
KNtykrnkjZNJ7hsx9bsJke1uUSrdqVjK2UeIvw/Gz7aegQ0XjDxq0/s050hL83lYRBBajtTSiDBj
qWm6eJM5EUCZkejIwpwDnmxNDy9GdEH3eF2jjJpSNpP8XRsgyjR2iqf01IOQWdJ9HuMfRf9hqWYK
xrwTOAY0rEnhsl8W6nlHIJf5jTtnC4Xjx1/LzoU3SV/JWjgZti1GBuBEKmU+zvhoawjuPe0Ii2XK
JeI3BTg9eoc5A4RuA4ZIG+seFTcqr4MVFK2NDXIx7Q0DVjOfHHv/qo2MSJECHcQk5zG3MipFGhFx
5xTa0g25GVlr4MHu8kb5VibhCKAKd6gc57CW5j6cFkEJBc9LMezR7FwSRXT0Tveb/ebcrpK/zITI
y06X1vKj5N8YMy0GEpd74xX2Vc0WDU/HHe6ciaouv3rVp3CNpkRFZdcASeittlXVnZUGtTexio2w
bKt1Vn+tkI4yiVcsjYxImmV34SdBWWYe9asZEU0TZwJIunl9jeAqFyoGah6JOHGEbxsw3PSU+LcF
cFAc8dQxJRQToSHuucakWBCFcSHR0SvREuQS353bKsWf+gAsc5V0FByfdpFopuyx/I6Et7yyOx2Y
9gmKr5e/Qnm1SJyZNlIpmn6GVjx8ORJjsJCSqjk+J8tIF7Ln3NhULzXIjEIyPvEosBcTV5fIEGLK
xMJfdjRBf+FBqyPOWkHUF4YQ6CEJfLDMVL4sCVqXJ19Ya7xvXo2X6TtbDPpYUpMeuXMSQlihJWHa
dDXMisgxXs90a8obyxsCaqBXlWLZFEewV/IJvohhdetXFZYppZvxakYJUFUhBejqqp2HP6Ehx6Rr
Dom8dINk/N49iOKZzQw9C4oZpgFdO5PGHnhq76TQBPmwcB1KxoxzPZLuKklh6PKcolYtXPEQ1vnh
jIYkBRjsaT3AEhYu0a1vll8oWKjRDipPNxGws8rJHnGtfdJI+xprV4Y3/SwL4Pksbd3ELuMXfnYq
LyER90/OFQJwXCXAYg/HVqkeoc6oEpke4weVDs1s5rLvxCSoH93M66Ms+Pmt4iZ8eZ2zyV1fkkSb
/XegNqEd5tvpJncmnoJyj/KlDEw5jfCxVlF07FPQiIsO6h5vlMFLFPz7FGYKcmH2GYXpVQiSSd4H
EYJMq76NSvnr/1cwxL9QOQu8x/PhwjTFfR9Hinftst7AKvhbtJX6TWZM0vqu3Rpk1AjBVHb2OIir
ZeDuQYaaPM67zXv1GN0NpHzDqQHRGV+KMlKKl0fLW6waLiH5+M5DtRIAdiYyNkTbrPXVqr/dxo6W
6xzhomlUHLXcoJt0j7nBVFDVg3s7CS63AdXImsWEeBfFeqqTXmMUyZc2+nZYW+TFSeXEdg+q28q6
WDstt3NUJrkdMWRP4500NnDs3WWfBWO7kYm8Lwk2cAe+jgAgWWVeLsvlp1fYyWidwAkf4QK6Wkl7
H1+Ngp8mYHcsRMhqzhEc2tLBaixhYNrJZWMnueY0lumTExxaVGq4aNdVQnwaAMfm5rZspLuWosJc
Z9vjs9hR9LjAX4/FxWUc5eZlEmhhPBu+uD028his84SggQjk/64Rk4YEruzfU//unik/RO0MEp0a
jNtw9eWo3nFIC10wA083dalsFPwzieCZ/xPylkdO5zpJcax/S5BUF8OZqqylkwnI9xkWLIVxnvYI
B4/n9pcJQhh4TgKM0fkarmAW/ChF8ox03kL1RoVdFH24CgH9VOKp0sk5a6ezeC/edlEc6dQUbjyF
LexBwXfA+JcsMo7X/sxbaBSgxNy8nMLuoht0hxS9ZAurFQINS1JYo+S4CE0GhG/qxNIfg+ROTlcp
smoTlSZfQuqw7KAHLk//RRZ3gVzzQhjbHHlnJecEVuBY/9yLW+gLZtYUe8uSF1scMZH8yVU2R7Th
38688N8pLy8fGjiJdhtE+Dxhgib5IZAUQLL/T6zTXghYDOoUSBWsq24dYbML/xV/ymO8qWigrg6q
6AUuCb1mUtFc7XVcaKU7opNM6WvL2mKikkkOctB88KRoXvyjIGqMGM4YacSd4/oBwmSeJENumPmt
hr9oUEdpH8KDFiyTg2pkILta332WaoExb9882OR0aHL/dYGgfZ1ZyTuX8J+ofyjIuM462VGJtSup
N39rB200gDGZr9/lWaKKuTS5uvlph4Xu4TGM2yizi6GB4UVYHqwQPiMB12+9QXz8P05Wp7UXdliC
brC9INmcqmr/ARsrhWNS5cwFM7q1laQZRzdvm9UEIXD1ueJMmu5jHd1U89VguhYDNhRZj9BTZWfc
2p4lmhVOjD/vEz3TxaIKHg13uHI5xYc1t9mD0nwRE1PIgyprDkMAqIITgXEn9idxIUSxbcbdCj2W
cN+k+BHCwuKau1ofDRS2u20xoLtZbT0SiGmgIcc0aWyW22yrbonGl+9s/igzJn21uV/hvTemhitH
VtY3rziDtvvfnvpG9UtDSarCVYbsyI8jpckTaKvm5B8xI2BlEqx7W9huwBfz19IoQP3o7W0xLHgI
q0nx0abrXr80kjThNy0Dj1kJW47eJ1DlzXX3AtaQqh+JqO1ltdQbZIuYR5toAK78EjL7RLcuXKpR
/8e+op45P/gQhxbX+4Xx89/iNaxm4AOnwTAQvuZnvvMqKpeGWmK7689IqZ3tSawljufJDqWpy3x/
BXvO/qBXnfKJGGFIjroI4m/5mjeaj8OHzL8IRmtmSsOlSzHyHe26Y5VpDKEqU67xolU7yjTs+KTO
0ktQk2JsIYKelsuWfFGIZWrvk+YI9tDDlhH/5EUljMXxXrRclBgkvqkaCPsAhNhHdCvDhZRAMTwt
rWfoYWW3EpCduNYxOIU7aTYS381k/36PV2NMLIRio/q291ZtDTJ5gtZD6tPq2hBZqobn50dTmLC9
sxZt7WoTxrphRpJ56n7pk7bBbHusQmSwLOxQHh9eDGu7Lvsj0xxLTKXpvuWpJvB/zhdx3aWCKoQR
Wt89I1+ZXqic665DF+ovILtULTDoFbQq2ngTMyRtfZYfXaSS1OIMz4DT6dmhkjRjg33ViLJxPH+V
f5GYLG4kN3tl6PFohQkbIVTcXoxI+/JgNV67dPKbOzkHflJLyr6gcgc1uIIWSrY4MUdWJWOhhzan
0a9vFw1x8PShlnNZVAklBml1R8v0mm6+eqk9mfzZfzBYhmd95WJsIGochajRnmVHoUDWEIhd5QMn
gPOqZfIBc1gX1kh9vDgmNaX5+5ay0ozT4jNHsOOSJjtokc3T7XU32cEq5pnRfK91Ro7mnWT14mF0
V803HU049n03oSqPexTpZISzP5XkgNVHUznVhyM24yb8JPWdn3pjlOBkHQpFzAEm10nRRMf/0HD8
9onPgnu9SvqSb4U6zD0ZjOGFosD+BamLKLksEzHfSueK33YFnsli1JRRjW9ALMJqoQeb+1awzFW2
Asu2+kgHnmUScEX5OW2Mb7e+FnvTfzSqppe0DYEaZIPjVjZzXAlxKyAZIu/fPMpUVyIa7L6i7BGk
8ROUVxD2uiGwrf3eQngiPXleh9sQPgcCFknqYxsptzDkt3FY2mD5SAmjhadhAsG1rr8OaZ+LstiN
sTxBnCyp33s4aoHccxJl8y+z4PING6y7vf/df3WGspxtMKySBZ3HwgTzI19lNPImEs1Pp53p9ZiW
qpUy+zHDnsoB0fESqW4DWHlyW6KcAqNVEwNAc4VjhuqyjXBILBhSjaUkRsKjskYywO1Fl5P2hNaN
JNWo0/G28QjxCTpAgn26XVbyjxY7Rs++HOybgYpXg+Q4obEVyVNEZsViRZnYfWYGniP37nvju/q9
EeetKM0TR6QCrhvLCk0c7yMh0+r+wYCOZ1w7nPiJ9YEn7XacxkaIvcs1VeWl08nFfPiBBKky6Lii
lihL1egkQSkRVnPYIfA/6z1eH8cY0qjwAjWi2Gs00NkvYyjbE/pyP3k/aaltz26OE5LINC/fWbsM
0aPqgKPmyZaMfjAlmjTksdLhzXEqLgfESyJcV0q2qQqpHXREVawlME1Gt+PT68B48C7v3KaE2V2g
Ne5SAJdJ2y75Xk80oOBh07X1/1DuI7MLAPqqS3U0Zci27h5zU/PrrLiShRuQETe3yEKnfQ0r5ari
Wj/w5t2TGaStgkNzHicl4xmRI+3MvEb06IUOvHa8HrdmEHQVyaWOmxuhVfEmdtYN8rDre9vB6lSf
18U/TBcx1yXKF8wrUYVX8bNr3Tk8qeopgLvzvQZvmubG7t55gXq8aCd+fV/EhBCWdWqK+rcijKHO
wfM9teVYTSTV4YZQaWdR9UmfQztsg99TGdpsknyt4snT5+vzqZod8SzOFNGGNYD54b/fqEPDA0jR
rKU2zIXmrD1dTuoqI1z1EXPXugLlNL3sIcn1sHC8IuXNAKatIuhc9pYRIKPiEC7pZsm4b4ZdBTiB
nxxJv/ReytjcPBExiPdtLvdxibrC2ycrxfObZ++ajHG4oFYnNiLD+Vv9S4Mnd093vr5qbN3wmk+f
9hRzYul8wLEqf5Cy+5fLr9RV+ibUmjVyRA0WuKDZTzyTRQGdADdh2pfKTPsDz/7Ure1th1UCaLXV
RN3rVkloI8jPbr0RMiC53fjNAWT64eCsjVIZXmcvvptZx7q77L2Ni75l7/a4JvUi7U4Omo+apw5C
6Jb8mMjoWXgpeSc9s3mSTu8qQOFckLq78Ww/9tU2Ad4C8Sci7t9/pNonYdAHRCPNVUuN/x0TWIiV
fpOVrVJtmSSL0EBImc+jdG1T/bsg7HQE/4YBXOeMmj1pvEAuxTUHnUgKgqhlevQ4skYjNhc9m4sX
KXnBLF8zMs/3VT+bNSDX1MjViqzBTKTDq/jhU9oxq251IitWx+uPD6m/BT5vFoRznupQna9CAFjS
hqFE5LW8ZmItqItx8gMiClvLJWrc+t76LK3kEkbgDk8Z8zh07UyTeXEQYQYjkYYGuWzJGY6dgJr3
aJ49dmIFrrhEEL5uEkpsnPMqyKn/SjmvSwNo28Jo9PWKj0qM6fjDjZ6Q93fwlAOkvLauIYP75W9m
nzSYI/tpKhI3/DdBN4yzaoZDHYY/0UV0K8f2gQNNE4IkoUdMjhJoOrVtw0u5EqqgtzgtyTpVBfyk
ndXkvLINL5XzvyQt6gWX4/L4KRK/FT77vlBGGNphHPxB+ePvoHDlw87dBPxSW9pIDMSJkKXi4lt4
Hir3h8CpJDtDLnyBxBP/JpvhhVyyPv6SpCkN350ggxkO5VOAiVU1Q7fnySf/PrLmHyIyc0nFzFab
6mL38Kta9Ai0cKoE+y8I7hz3xPOzRLqe6piIwCYUgoMtPCDiHyFAA5wRSLwtqz71L+OD+KOzt7cb
m3QXHjrcWV36VLSThdrYN9ZdPfAJ1xmZ3QdoibHWftEeqwDPrc7683cd3KtHkDgxnek/TMzCvRb8
+az3J3IN/AiIFP9C3xOfzd0i5u2hG7YbwOP5gOs8EOCOzvHqtabC2/x2ByN9IWLaW5/NwzUal24X
wf+H2z9aJL/xzpZ2ZRQHBlZT6lV6ffjVyAtNT7219haSaIljvbN1kSJXK4T83bGWxfVoCSWeZNZt
FdUXZ3+OA8HGNttdD1E9KSkdmkzAotg27ooWm4Y7a54pFPeKo4uUMXl9CoNg1uEQ/5gBXeX/5MBL
L46/T5sq5y7WBALfaOjWgE4re7bJuyRbQ1h3RARh+U27jYS4SLO16ZXgzNUx99OMFn7SQN4qnp07
9GPbju2CCnPuOAeuh5w2N7AYLm6pPayQXC93PGVha6U+MFdJv+0aPaGVlLFc4lUyJOJ9cTbBWOIk
j78KaxU2VxR6luryXHw0KMVfiZUTUmTuvXQsvPoTDo320nry6nuO4dBURdJnSz51ka/3ieoGGMRe
5x2xB57+xTTvWCuvPmSfOdKwhZXLuueX8FLjJ+9j8MSy2Je7TfuqQr7K0fCpHOAocDE3X4Euz9hn
gRIYMfddxshw6jj2730MOYK3lLsfvcHZq/S6Abi/HCITajN6eX4/EKegK4FKFdRizb6MLJb+niL4
KNYFx0nQy9/PtjuJf4Py8Rg6raI5V65RNwevQFMyetC2ziH2+KPaEffCnBQumHB981AZi3MfBzdR
T0pg6H4Q4kUMSlwvVYSVdBlk+DrVJEQgL0vZNZ7EqbXF28fcVl9Yse/l+0fJJNyGF2DSZ1+b2L09
2H26KqoHKPPmlHZSuzqZfYcF7PxZf7c9uNZn7jNxAgl4hHXefI/9LEVzLwfwWmtIcS2KG7xKn8di
X4Lzrhul1+je7KcPTyU9LKGI7xAKE+j972AoNuu37TFsdTGG9M/aisnK8qtNITpRac6zaKFJWZyA
Phlc06lM316E+0sxhQJ/5iL8PDliPuhQiPPEruwJrN4fPRbJXD54PCYShO5CTRlEBNjjhfedwNt+
iy3urAQ5KctkaGbbsMbiQQhF/ZHe9ov/pyI0SHh/DfHjv94K1M6OVpMT/z9Ono+wsUgjNLyHvIhN
EJW/iFIxCMSUVMyGQglKOsAEBqcrDZR2PzaG+JmIVnNH1jwNhlFQDr5HyA8ox1YCDXrm7CswH4r/
xBA2araouNblNkSqnrmukOfyt+Uc7+RCYVnDhHxILbzIj2yAL/gEA9I2C2pMtNfHJIed3OSLFgc3
1V3WCp3tMrQbExk7f0FxC5nAscqqLyvM7oYOmbKi+WGlvM58ZYItJKpWOwD3+NXB9x/9qjVsYCfV
NDfAA7nnmWGm29peBYWNXB6povv0rmS/U46OPcO9qkKt9ZQKRg739o5TUpsIMudF7MMdBt4aV6Hw
M51IPtDbExH2Ugr9W520QxD6Yhl45/B0dmXtM9ohogj6Pplq+I+D7b2jPmYLDjmdy1THNFior1z8
4rKdTVcarX821D2TbbSF2Kkuszf4qftCXSg+bdk7321/V6asHY5EXiZ9AWK2z7svQ4EbuILPjzA6
//rVAbEQJsBOEcTQoJI8aVMsCeM9Ue192V3b7BSlG4fL6hH9u47QEWzNWA74ji2Q8ANF9O/zVLIL
sR4TNQHm+wD21AWBO/QcD4NhRcHDptrwheRqexiFsTK1Rn2836QmxSnJFT9SQFyCsqYNCYQFsK50
NRfSwhhfOuGsapScYKgANQKZnCbFaASAbCBpp+LllqQJPA4vnl6sfMuZiH6O0Ryhmt59jouKjwAt
Wb1zA+QfRFMGJl868FcgGz5qVSjmsDFn2B8aNO6AwYmNJDuGp7Ajch8zT/EtMg+prJiUZzGSuGZO
p5Zr3frJY6VPVUeHMFWRe2Z5aiaTPaps5EFQsknw6nogEHgS9y/E+jXRWvY1k05F3XvD64tq28VC
r7dGmMDNDEmYwgbeDZiQDdQajFDu92Ut/Zx4c44vPBDiO/uJjjxPyl9YImK7kcH+DLem6Gvn3DnV
4HQ/gX2/bEorSv22BfZZ7W/3YaiMnx+VBG06jNyCsaWw+DlFWPJdNs0UB028hI1etBrZ0QgeQFyP
ZDZM5gk028mP11+FDX3/+lRYf91qYIhvWvxtBcX4aJKWb5GymndFqJmj/XHIha+8EecZqdWXe7Mz
vovBCZxk55FVQYkeOqWgkjHFQrKbW+zexFODtZp/IIEuxzPwoXirJG3WWbwfID1Rx4BN3NCCjH16
jdUc2JHU3ZhGL4LEaLkMyyxEyLITgoVNRJT3DWa+J9/b2nvD0qTjRxU4HR4meicDcOKerWpn43+a
UiKZ0D8CkV8lgF4lBaD3sFaDEqElxnGFePPhIdbZaTDbAXbATPppjkVke3UnNlRKa737YEY1odeg
WidQMu8csi/AYtm+u3dbNtDFBS+G7hO8y8JK0miVjnYHPJBTx6sHfe3yWwbb80kL4CRZ0v3O+VaQ
H0ODVeNKiRIDLT9xe/i6SuszjN9lr60hSP1eKy4WVL3cTvsv9m9dPdrEdwX+1VXbj0Gv7sXMhdVC
MbtQwq13oVNrnz1Ux59QxY0ozigdhziQESiHU4NAOIiN6slhypC4Aa/8p1sZs9m6NA2BkrAgnqGx
+09BKIwyI/eAs7SOhNtV3GpYDDAVDFnnF9cXsc6x/wKXqp9kQMDfifSRKdG2hUsZOih3ERZkwWBB
9qXxQKuC3Zd88IeLtq7zA8kDocDFBXhJXqQBJB927pG44j3AhmiOuGQiyA+Iq77InVI04N/i0uP6
e4E35ipWFd8PUi2r4PSEsViebgaFJJFoSZr65O0fRGDUpPBHTDgVgjS3YXnncmT67la3c2goF2iY
PbPVRjjE449CZ+M7bLlgA7EyzHQsgy/vU3HWBZwEQiHzzJsNI+iBr8wBgEGe1W+I658+S8Quux6/
YRKzbRHHa06vDQLvtU35n+AuaJKxDgWKWs6nCtDxEYY7sb9ISZ8J3rqKshfJPHL1cSAslrOQSr54
VXs4mamP7MLqhnAYnOyLFQCZ6kf9odowxzmozw7CUMXncWC0tWHItRzFWjS78GZVkELvS6WrcJR7
GLc+0SPIui0BcmT4NnhoYDTNjHcskMHjlF+J45k5mjfmhMxMvdzYwIjLlkwBycuppKMmsJa3onVq
ebhdWfbrDXjPq5ON2OTjv9HpxQANb+umKQXKgB74DqV9Zu0kzp1aZaMX7CyoQTsBsoBHQjAvRodw
w3g/wLFsRorfFZkedlsZMm6x8X7MQTo+dhl8ksmZE6NCZSAkrUdj+sd4YRmEU/dw2+Pd7e86NVBe
gn57I0OyQbrlqK+46b0cXE+5PRJOB1FPjtz8JSrzUbzN1H6SfhfFv8GBSiTkF3RtX3l20py8dlaY
ORc/okgLmKgMd9q/4x7GlvGSMpM3q6r7H4bFLI/ROeR6HQ9VYbM9ma/pE89zwLMhMxahCsa3TN1r
NxmLcAzVpIGGGc0tZDMRt5qyyhlJQt2oW9mOgSqE9ivcAlt9ROq63p7lz4ipFvFcJsjGkSNZJHF3
LpHnoxg9gay1VgrsfRlPcvzS04P4b73i3h7sMLkhH7S03+FPbNr4W9aznPQg5snT6Pu/btZuamIX
0W1h+0QphwBhgv8WzElJdzv68sK5jyqI329uihVngI+h6cCluLjZe6Ak20v8a+/TYYdtWptK1D7E
BHkUX3m990odcZp0Sm2wUxeyBN7JF3oNl6An9fYaTUOlmkiD1YrzoixuMC95IsCHEiDMgIbCRhbo
9DFwAXekY6zbAytDtXCioWkhlgl/a9bh9v5jAOWC7BlP7Kc1vKswKct31b1wk2MykpyhZ2Sar4TW
VwwGMf6N/c/35Pr2e7SPQL+fXe1tlUaajDHFBPMMTajRvf/05wfevlOXNQxS+16BM5QV+5r4FJvx
T6VFAgJXxY3NvWilq00QooL9b+JYmFGhplCG/x98231us01wEEmVUhOqWEnFp28/l8bimrMAUPqH
W+26X5aQ3Xdazzsb8t4X2356iqoap/49sLkwU0gVo/9iGXR7uWuh5efE3lU+VHuYbJewtQpBSXlS
ed/EA+ZBWX6tofVfntTIbijbeCqyCQwgY+aRHINLPCgTyG8n7WDZHFuzAaKO+wZ8NxLZ3H7lMj4D
23Da8cS+7uMEzrfT0aCWNPKBtx+GFSGY2EldhNid966BXSwC040wa5Uuu30dhj/YdQnt3VchXdQl
9ybn+twSyw6GrGkzMc2A4/ilTbO8vPf2cdO9qd7lMy86SonayD0M6GlH+IVOYMWyEQjL0tyOgJIJ
RUSNwuO2Hb8+Z4ssB71er2tZ9blLkwbsaN8qMhZoYfSDHCs7gCtJplMEY75xvPc4LEVVyeEYQBnX
ntCm30EXSyXIHoxtUsOIY94x3J7YTKqVoyBC9Yt1hEFDu8V0Bl/2AfvvL+XsL0XCyHCKp5Yfd47y
l+2ros5VNnVPjx6uUx/id7JEIfA2B6+KG8pWw+aZRP69vprlZ1Qji2ZQgGyUEnrWw1SxhqjQt1Cn
xNslxK5MM1/jMvlKA/n+qTGf7LjzIolelqjxqDnyVFpL14uKZy3ykaoBXBzECUx6mtLHEabmQUmx
3q5Idf+z431Dck0pBdop/ln6OtEfcFmXJWPM6ajXauYb3ugx0sQPQU/13mey9hQ3qxaAzdqzcmZa
Gshy0zdkjJN5p5PnBEhNzWDpFVRFZa6Ve/etu4SU1xhqfQmRB9npAM+v0Vpa+PCXg4J9NTIaxL+x
8Fdt/bAqlD8Sz6Ua3bBNJn90ZlfOzeFE0qV1cxIRNmqpS/GxLsYzajSIGf2MY9aTGJMvN0rs045D
IJ8GWsAXHu0H3NBKCuWChZ7mlsSyKrr+k4Mkqgj8AeBSVq6QCQRb2uJO5+pDozU2bELlHP9YJe1S
DB6Q5pacyrAzbJONgadaEhGWniq/uYfZmnpqyp6bs2bet9IGnpKMwGKHmSsdckbZwMsQBMHaRe4T
OjXnd9MZB2RoFhntb2oXNg7TEEmNknRuPaH5SD+qZ6/cchrqE+XuiLHPDSq96HY2XFGiPxeRs1Gd
3iXRRoOZmi9FAwmhrxRj3WaqnevmBDx+pumjwbW4MmLOv8rCHKSFfUvsTbi9CHvTlWs+c6LBwS3p
PerlNJ3PL2Nf2DVnzzZH+hhfOpzQ2OjmC49z+/yaTfDoEHVZFWEYyEqotjPEabGCyMdP69lnK2A5
BDaFf1aGsf4p0bpFR5cZwxTMIOwGxp1IAq1cYCWVBnxCV/rRLhNDDSEGgIbW6oHS0Q2Uzu0r4p1I
atnqDx0rt252q1FLHkk8OK1z22rUgDPiG0dIEeJW0GNGtKkfj7CzeX/2mJ1FtYbAJiC4E3ePHwlR
9VQFt3Xen9T4YmYMEqcWrZeU7nbsYxMma36qmPOmXgJFnsKXvIKTpw52RS0TLJ/Qcf9olITm1B4O
mmlND8AFgLdLbo5+l5rQoX4yHzyeaMBpU6kFyCnsrzU3E68scVbmDsJJOuukapU5lsohRU6BYtMO
Z3lFE4vjpRNRV8ZKScA+KW2tBj1ctzkINNKXHmv9OJPYgOPYN1XNub2SOT6YNVN8QvmxfvZCOZmJ
XEx+qqDH/YWzJPP317N4vEwmJzizYF9fCxphh+qVGn6Oj8KQAnenX5h20LgygKphIIxNkYlgoIJm
8Ii0wHC+8ausi6NnIHM1u+dM3Ttc/tX5qVgwT97AA6OfhsdXXkpSSLwQ03BjvBhanFDgYil3Bp6H
tGMvsRSjSPaYlMRjbYs9hJYXx+E4ZZl/LKeadqtEhlbaVOiUVDNgRrGE255ViEh0kUTF8UL5D2hJ
GcouxMpFzz/5Uo2rQmeI40MeIznWejR2unPeMKVPWlz5rMdUbz2ITBxAJtlNkYcYQeOUcw+fbB5+
8P8qWuStud5Uyi3sD00rMmJgDaT+uqodV9m+ogNFqOvqPEmgRipEeL1qQryI8Prp9/B+zO+slwar
nhc8rWBCTh9mk57o4t6ucRlG35oIhlxC1Q2gsUm3xygi10tqCuie5ZYivLqsQzwIshb2tOTgutBQ
OBV/+JoJ2Bk50t5vtlBIQ0Rr2SELumazn4c2G/yeO9BZ8hMnPYUg10fTAbAzR3eU1a4N5FXNvgta
HiugfFFyx3xGMNmxX5ytC+j+k1VFE4cOTno+FOD/fQAR6TXBmdmjaFgDy9CS59X5s9Z97r3WUzqn
0iNv5V54rlSqdgwEhK01zxieoThD/V3/41hFGKaW8YkI9fyiTATvkm6UbyQqIH4k6kc+iYT40Rl6
pWQwUXiflpaFg1ql7Q+VtKZnECSoK2cA3ageI64ClK9KzewAzzaHkg7HA0hcert2vMdWNhF3iRR8
beTiMTpFawrJ2ATa2TtCeWv29juKdqmBuycqcmjZ9H1FvkxvvZKMWZlVauaIjLdGzmp+LJwxwLhw
rAGp26UVQ6u3gJOaP0Bi+V2m5Qcemuf6Z+2d7rGNSbDtK4PPDjN/hDzVjkYQLpxXdvAxcMOtQbC7
sv/NEtaJI5FplCs0aX3E82Ng7cj7wJCHEISFuNmYfkR0DS2Kv+f+R4a/9x40KyxdaU0yhdEoSGdg
Ci4+4NVFvqq9pE7OYvm0XClvzidG4J1UrYPVG0GLLiQyS3N0geT/ayVbSm2irMrgvTbW9zkCsFw2
oOyX8iTTbQ+FV8Zt+e299CMxIik+rdSKs/42/zNI0q5uDAecGlYpBLHuoppBLW/XTSYeTqDYHuP9
NNZOrB9s8EZYiGwni6iayWiW48iWsMuP11nD+fKKyvHCZFp0gpBgW8wh0MTpM4LA2u5S7VewHIrH
NMhiSHiuobaHpHGQtu4Y76d89g8vm9kSRho7/dVOLUVhcQtBhqOBkaGuO4HIJibwpKp7lpD7sVpc
E/TWt9/LA9Y9N/W1ZD8z5eY+R9vmJfRf+46ehln/1i6mv4yw1FIKw84FzJzBt/0e0LB7jvR3Xnb8
cdSojd/XVjqP2bQJD2FLMNXz0jDyH7TYoVVgCbn0+gBPG/Mg+booChsn/U7WXX/nLIlBwzRKetNi
2T+KW629u8jF+VRkSxVD+icQzx9ivFVscVsg16j5GijkuKT18oVuYKclVdn6OXwJvSfi/foXb1Eh
lD2Iu34Im1xnXofyETK95JI2pppAhRBqBmdwnumIl7LnfFsvc3pXOCy4rETI/MKJcgzwCLrs0nSf
H8hLDTrlCMMWEdIIRoU3PnegyBPZCTnC8o1691F3AVnyYA5mn0Pat8Vx2vlIGVDHZnwUJzpge/Bz
7yFJeuC2KcM9EAKefj1Bc1rtUTEWbHtBatR2gqeqKqxj1Kww3p9okxsPbEcs0/1SCIMHHcNeDnNn
2OpJilGYm+ROmnUal5vkQTLn4ucLnDzATKVP9q9dOpN3/HUJppXMV/+3TQqIY+UIQ1Fsqii2o9mP
X09H2ksH/v5/fZje8uSAq843PVDKTyUtyx8Yk4pXbC1OzfXx11QnVYqZrnCaLucpt/ios7RC2jbN
QF1hO1JMRsk21pROYd/+0Fu/VX96fgXWxl3clTsXa1bAvNGQoOb+SCOhyo+WLK9g+0ppAeXC4G6W
G5HDCxcLxBunjEm2g7k/Mvi88imawIrOeAxGVNOnSFhs8SVkimE9cBp02caswOwq3bFRMzUxVyVT
BgZKM58ffDwBvXf22B9vVMucg/GzZIR/YMkhbxHOr7SvEe7uOqZR6K0a2oh3LUXaAksUo1emQqBo
XLadbVD0vQB3kZXKLh4CkSuM+7J6uW5KiBP/Z13toG/EuXyYerEhzCSTt9XPtLgUY55QNJwVs5Im
mg4HBSr8J32WsM/Op95j8ipyJythrnhW/c5Owqv0ATihlxjO046jWyZDQI2j/nVapR2md7uoOPw9
sx6GGXZq+EjasJfMZiJd5nqGFZBsYnic3/3vu5LRzWCI0TTkuIDnCYRzj3Adp2qVnvfBZh/Wmesu
kIpG08zyaARjQ447kMcDYNgLR21MWcs6h+2BKcksOVBuXAk5aTwrIKwAtwE7VlhPtpqZzIKNlWH+
CILh7n/LMGOOBmTww0TdKsLkgX9STxpN1AiTAPQAahri8IZByi/3aQA8E4wRIrJG6LbPgRR3YvDO
YZyWRzacMlLqtggQibFhfVg0EadFfqh3dc3HsJo6pQoTSDne1VfonNkEgnhphRN2g+EK4bebQFhC
nx2zYVFZCTcuwyOFEoQlAL6zkXCZIKwLCgMXIzyo1wjZ/WsxebXRmNHhR2MN6hiEV40EtPlK03fe
DTuFEsqcNW1dKYRbXoZEw18BPOWMrjCNS+X5DxJiq1DmjcoMOKzjse9iFwJYNYMqWLL3j6uThNms
u4hyaQJ8jIX4s+GrJOMlu0hBrBHDYtk3f8V4rokBX/AOUw9Qxl76QrxPeyOM65V8bi9IkDWPzRkM
AjSz1UIzWHQk2lWlzkFiLzE0za9FJNDY293PDq/9f3ocUEn6NcLnvpyJHRG4MQn/clJ29yBYoHCv
yGfrvnfueFgx/HzJrv6s+sNYASNUXxuVAjfOVfhe8ZQezJafqRSna9wD0YiKcYXsQoHZr5WTG95C
rn2Mm0WDPkILqXtpx68KDt7aVgsaww6pzJnHf+lnOsW0NqSvN3f7KzRnCNnIkmgAvkk1BX6O5d+A
ydEss3sN22URtHVOB7O2F1/Paska7pVxfhfnVaN5gsiE1sc01mYrIZVkF/wmpc+iRyprQFi5Z+uv
gMNJzdVtRtWcEjIAiRzAW6gGrCwhhJY4X/sYkoLLc5z3J+9eX47cPzNarKsU1S+UF3Ytbz6IUrmz
R0XsNNezRjXHHbc9FlS+u5FZRtXFl1VMx+he3tMCqi3Cofa5S5lS52mWK7pYAv5lc6bUvgVtxpda
UwgXghXEjzYC+l70r2SXpoPIdXhnBucpn1WB+wfgd8cqTuEfnCfZwLxNitfYu11qUJH2feIKvaSe
eeCA5xWNWP2QEW+mUkMywO3KVvUb6MMRlc1ysw9yILBBHKTtv2cmJArXY6qimIefGHvrd6vO7mTM
unvAVcYaDjjcvQrjlKqsMDGdZQu2mxLL82PKRDuEdqhwc06b0bddR7AAAByohHAb47Z6/RkWDW+x
+NR51YBLkCxK270EihsWetOMwqCG4NhxxdWBx4qjFA3CRJixBFHNonPxaWecZwUeYxPxeaOX5j2i
mpTQVHZqI8OcIZae+Q0fA19DfEwC5+v2WNuBqF2/8LPmQDKcQ1gqE3jJwM0571sBzrDRxtX+GoMP
ClsIIVyyVejKXg3NBqPc3O4vI1HSVwjI/d8iMtzfipbJ8WoIxYN9oh3KbREd4aTZeQip+g+WJPsx
mncLXLqO/pY8vrbypLyEpi5D05jN1yfBgADJyKEUZnPpKI6rsYIIr/ghKZLSUsD6zKolirYaQRrh
iMSWTTMZ/B/j71X2Ja0i3fpL80QhJWir+lqLahaSSffL3zzKZL96+nwr4z8pxlYM4LFfOcDkqHCh
vwAOvV/JAFIk4IwP3vJw7TClgzyAQ2e0zsKdO3oXIUOT2uNFkgxVXZXszGy5F5+yGFD1uuN1jf1c
izhCmhfP5mATE/QtK9GRRhKglLN5JHeyLc0yaOVd546cCtVf8z835P4TBNhNx7TScz2Q2WfKmK5F
COXQilYb4RGRbKXa3wMnFkqDO5JuxWubVCfFUB0+7IIjKW6aoqS7d6vNIqM0mSVyRLDG/XWRqxz2
JqWOkcPJf0+EdIiW6nX40qtEp1ULyEpK7J4QMMh0QEXx1woO0Ee3xdxTKWX9ZPnKeJLayRIkwyyP
Z0UOHcQl+iwouck4m4U1wWMD9m7ZeXdHsgyxQQABuYXjNZaZCx3cEYvyzsHT0qKFgu8XBI6G9L6j
zzEN82VOCeg12HCaHd/SDio8u3mK6FLVb8n1EJwt20z40aJ7/P+G59uRVxB4pmLg0uoefViRREo4
S0STPdbIeqQGG2yqdJXgysaR5mgNb/ptHqlEtpZZah8kF2JWJXP/olz7nMc8H7XrY5VMroQbhlTy
cMSsP/OFxL9DEEktSgJeVkhXOv4cGHbHCVHpuTXUP0p65EGGwYBKDUTdnfTCUp8ZOMsutJBirL6D
5M4Ae92MerG/px/Dol5vDGio/67nMHxVz8OHu8ljNiuqZeb1+v/5ruOZ2HC5NecnEuXwg5TFOSeb
ou60K7o4fwV3NYnNSMSmhJg+ym13Z+DclcHBY4r6b7Y5Vr/n5fOIy1NlnFDGDSXVh1q7prTOnZkf
KY03HrztdnBRtjEruye7PhL3062iRCImJqGrfgy4YQaqKu6YAdB7UnGFurg5DXWuh9I0F8RKC4jA
bKbTUC/9upg5H6M1FMgq0/FklNAVxeMa/K4MlxMO2tl0afXKr/UrFYtOcjMnRDaPsbwB+rvW3IL5
SRm/A75q86SeOcGwHh0FZckRC4WlWI7TyJFINyHHbTQldRdANSLpyf8poQ0lPsZ2LEKerYJhqTTF
I11pj899Qu3da5ZDJ9si4rFfbzekiANVLTYY7EY8Bpa8N2LfO0y8097C4IdpFuCNwevNrDYvBSw7
ysIApxx79lYhWPHVSPf5mEe+PlEXwWMbsBqPt1c2EBKDgT0osug/56Lirt2ZzcOZzwvhFL+REobG
RyLFJNVVOsOIU0+3cPQk8/UsJPJd8Zs8nY+sOgjEgpl20RO2qDRB2BrOtvjvp4rNGNEh+eBpYsYv
heLBRe5fBCKvO0F/uTyoRxTFn4hRpXD9FBn+vrUxS5Td0YrKyGXjPL6Mm+Exe63AfaF3NdCarD/S
Ml6uue7NAKt+bSRnjG0BGP8mpU/38jLDiel/7TKJLtK9QIIssrJUDNKzSFs6WPT+K2uGcJb3IC5o
z76oMhw0lw9HAZKcdvQQhyn+rikYT7TSVqg4KhuIIY8JYzozDuoj4+Qwub8FQDgEE3BBOWm4P0gB
I2TTdhkaNU3n5ANDoFXF1QUvMlb/cbRPOY/oi3OZ0cZydjuAq40sExcg6hM2wBv52eh15dIL/tyN
mUdFLEzsTA2joh+BsZdLU73n3yZTEZPkQhx7K6TAf32DzR4PRRIRODObZj9JZkRAOHNROaac6Ihi
SfMgZT7pNRWIDSljpNFzqF3nbdodi/E/IJs7XqggvoDjJHtXzl6+f6ZBdJaQqD0EsxsAGpeHD46u
rZVQDLeDxrCUCzA1Yp/2n0WDYpVPGwBXj9krkU5HAq0qhGR4B42Bvrs28syz5BW6lPvnc0xvu3TK
l15oIFXqAX3w9BjmVI2+cTpcvdf1Q4UYkDgxCs2gqk9l7Y5CsGiEdR4nmolRiIIVY4GnJFv3NZUP
S+L4dsaJgb8G826XqfU1yQPwRZtfIgQ5lB303sCOuKzPcVT7oJWJTtRsZBtCtHMFqMKhJsvSFajn
5EGcXBhEXMMmS1XzEhqBC8gBdCJMlLg8l8Q5a/3iS3vg6mbz7r+guY0uNInQBVi+u+ulwNGNYbAp
3LiuK1kC/fyi31FfYGqULp9mZsWhnqe20aqJ3ExFB0fUBRqgGvegF6Gx/xF/pm13s2Xch5utynNl
ePAI9AxvjqX8bSmQW50A4dxcUZ1jwWohG5UhFtaN1+FRsHnoo8v3fB97k2dFYx8NAv7NTclIONx2
aLYk8lPB/koqiHJIW2IBxq9KGsejU49sc0JKDuiuIKkAJ9tx3KdAqfT77LRbz9lwqobErjBwBYQd
CmS7ss+FwT5T/Yf6vbIA1IXZby8u1OtLNe8JeXxq1fXHTFtWyZEWPIn8sDlRY70E7x4HyGrEB9Vn
zhNrpqXhlhPNd+3UPQJBJDkovFhfqb6owtEmkldQwpFubrNkxxud80rorD5rkL0eH1iz59fpGe6o
GwcRk5xlyqJRFgLfuMOYKehwAJbBSkxTlN5VZDG0c2K+AcarbttkXUX3gSQkkC4iIXpJVA7yFUDg
8Q97NkKJtnSPOO0ZCLVkdPPFPzIL74e395XZSch16y5fnctUoGUI2P+eTpNISZukXwdwOY5+XeJs
0jUUXe7yFLtZppydpT69cRJEqtmRW0BpCqI/CSxfJ0vESi34q7FiOw9K1518HrxLLaUks5UAy2d3
FxvnXwWQL9mhW24TYEI+nT6XiYAntL8gbZ+jdxPn0s/9YtmOL+QBJlaKpHtnOj/db2Tj1jorMM5q
ghQ5AoSXyHKik6YJKUMZF22nNaFhQ2/Yk4WP4aBf3dffJoSHd+Q9Lhb1DkPc6sIyjuy+TYepm83U
4h055x8mbjJakpe2bEo9w6bPw9gf1VAlqeEwNbcALt4mbS48hQdVwdW1RSZiyaGmvOvu7smyO53A
6EsyGxDrmAs3G61LQ7JMSLs2d6H+JQQFCzv46trJ7vA75kXRh9pxSrbLlL0/MFiGtBAmpIZiY0hW
4sT0in9n0+EmslOOvYyV4ZA/etNeWVuMkrHTHP49sq9+HrHp3E2Bv5Vw0YfXu+tMibiPFiyhfCmH
yU9ThuDv7+fMy4/8qw/PFevTSwX9QxGhswLTRNBiIniiK8szZq259HiTbaOuWXOP6bpq92X1QiHj
mG8HpvXUs7mkf7o+KtbnQtu82+dChtCeZmRAEmq8JP96D+JeCosy3Gk3AAlx+PWSpYlDKwphfW8g
6Xn8B1jN+MM+7y6DAxgcIcj9Mg/qfNIcKbls/PTbyqd5wwg4CtkjUynpirdSSKXhMM/pOv4x/aUz
GTdqIQGOJFzBg5UFPma6u80nCDE9Yl7bmQ3udMeC0HmHA62gYocnDII3Tck9nK7INODUxfSrtLuk
n6D33RRKHD1C00W2hb5boStMeYBDS/QkrDsKmVXbalrfTy4FmCom+t7EosTBBB5q35qvBoJT522E
o/MQGgrmEVjWQcWZVqoWDv+T+jaVWSNfebkuet1R3pP82twNDTboCmAcwH/B0aG/j7u+GCcpRrBf
/8szuIFRknsqvtTo4ewm1wpXeaSNWxtde1k1vJlTf9HLtkaC4F5+QQ944CWeQIyIht9YBksaZ9x4
Z/6OMlGNeajI66QLj3zmTK2q9uhmkzZV19ruzAEHzQhTPYNDWArN4APRtI4bc0N+04yGOhiYCzvp
a2IUjhQrIFTHqdTA+QELpW7Sq4ooOJi/o3/v3vzPqzZDNetPF1hHH6mUjUS3dzCS4TZGYCNomS5R
AFnXngN4Lrl+D2t8yp48phk41Gu6oG2FqExeZOkkk5g8mMoA/9TwiOdN2ymNyIjpde4fgSaj7krM
cLtL38jqC02MX9VldWPdaJZpaLZgrGR7hy97p1yAAohwsaY5OJhZtvimolw8RmlV5uUN1JFcpBiX
Yl+r3FY4UBm4H4KIPI8krI2lmIABmo+GR2Ua0Dg8Bsx5KGLSCYwcTu22r5k8/v26lIIqQ+WSC9g/
uvaxWPdBpyvJHcpq6a5hP0+XWjDaHfwhs2TvWvDW/X8L6+IDJQORdUkYn1uSJCykS76pUWVVj3I5
9vEZAYatN815Wg/bTGuzJnLugrCGiU5egN+PKi2W4gnHag8i7sza619eOHmZBincZWU+U7uPgXro
LEmDLR0bD+3ktmZxy7zonq+Q1CaIm6JCxyoZVoQ0XXVfy9TL6B3kRkMHx2EYJQ6vFJgPUi9ZKN/l
YAj3SuJ/h2mgLCs942V/s3MjATtWKg4RToSlAQZWov41rA3n86Luxzwrpw7dv5ZOKIRBPCFZr28B
69Cc4RqGYtVFQDItXo1kdJBkVJP/JI5Gwh/15SCVopszv03QYMv/BMGuPVAPT+WiYiq1xt22u7Qi
vjIWvSVsswuYbWKBaGCmplWNKLlM9arFRdsP/HvhuAhn6+M6u/NW5fVHRMJEYdM9SVcDYkXel1x3
eh76d3Fg0+bCLrITyhsYDmESW1bMjHtbC6Sis35C8AxV2NmF4IccJC4WDtjAgJHdZtQhX1fRDCGC
K3mXnheZJQlFA7g/tKBsXv9dzSg29Q9e4zDAT7woYVEO0E1ecRHZbaYHNFCJgrOahEhvqGUT0CwK
Dw9JOQNf4wP+ME1mhGF2O6Vw10ukTwXdwqN2Uc20k1RCUB1mOi+q8gdyF1ZKRLuby306Eef3u1QK
WtU3wrGNiBXdn9CoOsMX1eLrZfvGMZ2CkjtPJ+cezosS0CZwQMedXHy9rIg2+QzmdEhTQ8GaEHo7
O6bN9yqAwCG2opbHf3qbP5uBJUZf+qwlz1KRyJOvcayJ4cPu2bm6tNXtomcK73yxGkfihHd1TadJ
/HNp7SxYk3lZCxu5WvXZyLi3nsQZ4ZIyTOUwIgABtpuW1fLJW7GhXmC2UmdxPfQ1J3kmyXlQe4Qh
9LoEOCMOr1OMNZbbqwPUmKB7TVtMDVPRqA5Pu8t2NiTLnDF0ZKHoGpdZUIXz5Hn7XEoku55b3o1Z
JoYfUnTBjv7D6J7aUAFPgnRxeCJijCizBmFiPYsGSGD4OVBbxgdPlQD47eMZv63TAfBOMVnjJ0jL
M4cD/3soAwmlvETdLO6JSD9MXdbiPFTb/taM1ui9j3j7r7gV2e3ZP9M/cKy7qb4jhdJEzywbsfCe
Ahe0p1WdfPSjhK6PVpIGv25rr1F4pU5yMXtmau3htpJFeP17dmOBfr1kko4CVj3OVsinD1r2kmpU
1pbXGSSxprduib5jjxa9vQmizToyHCuYqpxmq71ceram6x1vt5rtzgq3jbdAYA2RZGcDEdJIM6kt
wW7Iomo1sKX/oZFhTYlEPnVvPGnwx1XjQ/I+9voZUABWdUt0klxMvcNbszL2wutBMwcLDKtFqvfX
QkpmiDE8Fiy3YZ9daPxRTIIUzh40H/y9dsVgTOhzsx/dchswf3jQcSQfRTkF63jJuFryP9aUoNJh
2ovhqS9pG33+6BUIGblFRHK38IsFp/lFoazWyErQXgvgPm2HxS2W2p2QTfk1jG2F3JB0iHnHjaRD
GZRzOeHK20qjZKU7BwEPpP5K5gfLDIIy3VFS6wmLPtZrJuaq5BSFocG90Xwna3w48DYlkoCfGELw
AV4mvGcKANZzAPrImgAnWGLmRH4sIXeKkJbZl/b+zl/Tjy3yQggTCnY69W9v/DHsYS+9WDp4M2Z/
dl/Dv/Q7lLwuolahMIH6XSX+LC+KNJDoWn3HZGySHszjn3AzoBiE+UYcKzknhEcz2/Vav9g1JXW9
VEXSsCKKoEdkj4AugXGiLq1p/XUkVPdJuQA9M6xYtWe5tozApejfSkMDBacRshgdg+QQNAZfYEqp
l/3r6JXSRQCYC3JK3SVoqWeF8ra0siTfrMqrIbpardvqIqRUZ2F+0FSGWa2+n9zJW8sjWKuAMR3X
Ofsf92k4V6f9sqDPM4k89EuzDHTNu95RiXgw5nY7UY2F2JEdDYozc72MnND1V7u6/JIRlmfBhFAS
aoPWUoGlGRUxT2u3k//CbINPkPYvMvQASlHrkMunPdIJGSAgylaKyXMOxn3c3dZ5HxI/yz9d+E25
ZKwOnj70ZHZdsW4U9g3/ekUMeofimNLtsyfAkWVTKQjolK3CgChc+HCXjwT/fwUkqBnfxnjhrnv0
XEnFlEoQKqL2Iyxbj13rSCfAj5EKyI+JvYbFR/NY7BEXY142KFiaZYdDwuxztPfIxsxMw8HYdvYs
R+z/AvmSlefieW5FrJSavq+fTaYUnmBcYX8cLhTFNKZA9rqFDcf7glC8lWaYJxq18Yflw/hZrOGC
Gogyq2phP1Pwf4oiKL7Rw/SukBmmS4FLPvEy+xakEBC5tgjh0wtOdzS7/pZh3CHofR50Xzzq5tSH
Qcxmw6cT1N5m6lx3CUxA7YMyGYLrYGIQo0ALUkRH1I3Hkoqof18YTL6ozE5KBPrnWBrQxqd8ukbd
KrKxgqIiH8gRda64Z/XhfCbTe87Z16hRWulyTpGcfV7/q6pTAcVnc/1t1wcKJzUy6rEcKqegOxgT
9J3MdX8rlX9TWTs8j5wHtGmDNXg4pQ5DHwhAT72Y6LOp5cIBsV/mSh9vsJXIhT3Gc2DuMTJCnAB6
R38CzJ6B/PyBEBjPF0/jHIl8kbZZmpCBej/45jfNBg5slZbC/XX1/UsNPYW9zIW0yQxY6NcUXz1g
grx5OXcpavt+l5V9SdhFrJTWkLXyQqIKulJ9bZ7DFtffA/WQsBBOEUUWoTjOWDAjPOIxm3TI1Zyf
8waDyZN8eM9hCrvhY8JtGiXJA9S5BM0/G1ZanIqRlxZEfPc3MqkWRb25UWx0of0wah2txPUEHCvw
1jMWSok8MmSFF7aYP4drgiq8BF0TGhLL+ejgdOQwkU55eg+mpiKRmiu+mEPA3ZV6S4lkR0TQS8RW
sdpW/76nBnW1B+o7ClyA3LLwZHDgRd48RQBLNohhFQv/jBSjE6IFed4Pt2fPtWi20P0lSaDcDnvZ
YnF6OibhOwd144NufDtDFSxAuFolquTBiysH/90umgjVSgCAbsKRlK5MpWHLJus3niLszTYOm1Jq
ZDFqzF4gBBQAc23MiT9H9jeFEISycXITuFRG9GAjqI0FzU7RwEcWddvrRXJtZRgn5fRI1uwFz0Om
T4pxQf6k2MR2v/Uqz5A8k6gM8Pi2fJfDhm6Nl2T7jKIXl4gZnyBQi6gio79aumuy7uscLFWzS88L
k88+jcMDe53zlXX6H3HySALA7PpccAaW9nMtokpLHd9/HM370IHUmDEX/AYttuxE3obyIEdH6J5N
WQIZmOBR2cVtJ2GUENPcl8PMH+cDZf27aOgg5jL4+S+19zvTj8uXV0q3QVuHLg11M4Ox4Q/G3e98
ZnZaRebsLpoAna7pSWNyWEncSBSReAxgQEwDd5PDLbdWeFnahx9JCxODU8t0tUfQcHflYnToS+gr
Yqb79aLBrbPiDO97z8YjkfQwj15Sqk/fSYI4Z1sN0qnaNTbvUcM1nZj2jg1DehiTboaaMQlY80En
aLd1bIbxvMSkXVtm8/MWSE5vi1hdBVvGkiffi8STEGSYKylBhfjm8wfpYIZH2+mLTfgMUHenxqCL
xkyzpyt2NEPwq7YQsP6TWgIX1O3ILarcHfQW6pQ9Yc9SbQfCe6ajhIIPu3+n+Q4WUFcvfH42vxpZ
idOVr+QLTsNuXlx3fNb66ssa3KbeacuLiwq1iaZjUMu5sCeIxgBoj/xuqOvbRW85TB7xCiMMIWvd
WanvrP5fpcejmKV/Tv2vhBaFgabLZIjdD8K8jsVRlL15ZHuDVne1VMBQird7HhVNcs1n8QkwnSm5
mtftDzjKe1/DwizmR8qqG7RL3AoJILt4ZQ4ltJnlSm3Yrw2sRFTPRBBsGRMIBGutRmUlp8IpJxj8
7F8C6NplLeXeLOAY/JEuHhxZSQMxiZux2Hkb9XilVHsezpLkDciVGP//y1CKlMwNGEVgGg1B/f8d
d6Dc2tKqi/0uLenNZaA7afNWAF/nHcYUKcAvkFyn0Q0VFj4CtSEDc8WIeJNuysvw6Zkhi+fdgTfl
GUTSQUDxoyLB6EirXgo0sheIWJbW5/+iFygy3njP/wwOvD08euGGlCoK7WxOCS10aygUQppjLqkO
LMAP7cA+BbNEOLhYqWvfv46F2iULiXpgaP10+e75c58kG6W67mmCiB+qbwuU5J7voLlmhfwgfVOm
+f/xjqjEtfSGD+uDFsTyCrIHRH3Gb/d0pC1F2Fgj9Xj/VXO2GGVIyy3GJ8s0v6TCkAMAEF8gyUST
QBoZfGIuuKSFh6ME54HxwSSvrSYAckg7TUmAbv8mxwXStYi5MO7tgouOMoE2klz3w6Jdl+F5R4bT
xUdNr5yH6Gyt5j4K7f7PkQTPnm2koUxppgEP3QMC+OdIkn1wZUa9g/USSmSOgf45d+8kfEMfi3Zl
0fPgo/ORZ3EMtOIP0dU37htg2+0GheYQKCfb925DEUWtocpbs54YT9eHjE4L5vb8kW7pyL2z5Hly
bztfk2qL/SZNHp97rUAlp+eZiClPwIQ7SyFPeS7izfiAor368KvcM867G3hiOEgcaG+r1g0yWkVB
uLEyQmPtao5yi4rksPe+SOTr1BWPCwTjMkIx0kAlk7FT8dVixRHFbHT8UNAdWmVPHGSW7fLWnsiN
HE6r48gv8EsZzECspdW44CPY9pn6IpiThnda9Jv0YwVSaF55v+ZQF31/oGgob48VITcqZNRkuXQ9
6Cb7yGvv/SO/t610vs29capiq604fOsqg9cMZH93k0qtYtdNMrnLmaDw0PvkH/GqIP3Ri9D39wWG
lB2uE1iEH9saC2qPnhP55W/qgwLtKFIXwwkxd6n90wYxeyEacePFA+0A4incsoY5a+/5CunCpG+p
keTOWD3jdOT+KUDhXj3brH0m93rKvWlFbcbAiFniig1H8JQ44VF54o6wLpWP/9JwUb18RSgLGH+f
rhO5pOW+/a50hKVQ8HuQFWJJLz7Fu63vLjyjLJrmzKb8IeJkrisC93GQyXVAqZOCAqlRcjt0SHz+
SJH9Me9LI9zvBCuZ7jJF6awYVHn1YAsmB7gVS9VoKZw2fUj4tw1kPNFBLryzJpnXqrnKC+I7PXSh
+E3aaOmQm8owc5v1xVBcTq5HrZvu6rpg+Wq2EcU0Kq/WrF+IfY+mdAddmXG4O+6VdqbIM+Ew5PrE
wOO+rTPzHncGkm4uGYL+wzgbTP1D/mPc3s8peBLBHt5qMpCESbsVocIN7xXVWQADqoEDcn+p/ZGp
JC5xk/ytXMOTkRuYOvLaBcap1VtiwzDR1ppZMr2P4AqbkuGM6pC1nfj6vHSht6HEBFrFzY6Pmnp4
B/av356qFAY99c64ZiXt3g69pD/dyX/8meMp0vbdoIfpDv0FR9W9KACH4b8yDxhluU+RZCCNKms0
I29sFhch8g+F90Q+r89gMk5OXk5WJdZ9mqq2bfH+wspLopM9kMzeY8ryXMAKvUohksSLiSBcI4Q0
ecYMANgLSX+Zdwn82OxvTE/Fy4RQ4ko5wYFCh4VCvn1O0o5ybR8dC6s6zgVCmp6cI6d49xD2V1Rb
N20/Lk6gyRRWyfj3sCKVl9LGSeTDR+OA54NskJ3OS6gIA0TuT7PxsVYWGU7LbXqrx7xK/4LHvcNC
ig1BayeM8jS1tECxdBAcWKufPIvfsrwkv09MRrmDN9F5vxySJK07BCMLB3MZ+dmuzzVg/80/Mfo8
n0H6eLkvqAC8lmHax/QWhxkJsMdD/OokY8mRzSqyDCaXhJxbZw6FxlW5sf0l6+sjLiiPKdiNUuxC
79DFoYN1TZlU+mtPzmbW/6zzewxxa335qBVOZv8862lGfSSd1ov0RPWWk3WtAZSlwPpm30FjfRuT
diRd+mH//D0/H7USzYI23GY6bOIPm8ocAHqguLZxmHH5tZth+p78llz0gq8m9yNwtXvn17UzBVuE
DkgFT/A9MNb805d14ti17oAb8nVfpMkqgV56Dj3t5X82oH2uYw6DouIYjOIvOoDc0bAaIRrZ2Lsv
37bHzzhI9k4+q9pFz1ZlL0Y1tP3KgwJIrP30YdFaPVE0bLNGdbmgyHpqpwxTbjtpEqxH6ugzciqG
3Wn0EFJRqyDadq7lz2l0aKf+HKLRRJQkn5uM92CcaJzzDBKeytTywo1Q5RmOUsATxy1J6EiFQI3u
I4vZZTOORRnW7oDZL+5+hZu5k3VNDEWK5JDv4DXkhbixPwcSuDM2jYUutSvvwquXKm0fxe3Ds1Ns
eq5WJhccsFUDhQ12sWDXiOuokfWHHEW7wUfwnksVq+xbFQv32XbreQwwwX87LK5fBgdpIJf3fqYe
kIUrnkv1ihU3A+YvRQD4DjXWEhhJj2B63P14nJCje7HoFohOvDSzIvUVmwPNMpKC6H72QGte0mff
Skmq3ImRh17C4xh0n1dW0E3w6Tl/kmS81mu0M1TLfFTkEED058mJrTcX3778AGAo6l3Xu3+a2CTn
bNTlRL6lwc4o0tIZWuRLvy8SZZzqdfxQTWC3/lqss/UhXD3+lGu5yjEEBTAIkOUyGzjlM2LWhOHz
+dCUqqhSu5+u9vJAClSfoEZ2aJ0BrFAU3+vdj+ABB4MDO1SMnEGswQHs18iCGaXJqQe/fsrvfADi
hlFJGnDeWSvC+2oL+vpguNtZoCD79ANVPfPDSKgqErvUoxnQDI96qqQ0oC0T/zREBr4l7p6ljlIK
3UihCIxoOle7XiBsGmEUy6cOAl2YmUljqeX+YpeIvFupsEfjXVQ8DSggSZrTIZWUFsztJoVvNnYe
jf8pyb0ZkoDOP1ItHzg8qL4G9d9YxpWnVkVLojVSwHln2sGgOzXHLy1IgFpfx5woNuodqPCU2rJ8
ZqjPHsHMzY2iiuNCYSOziN2KUfl1YTSlhkfSTlcG9LuHLLfI2D2goyM96D//UXFmOG2VciqD1kTl
xP49FC/NoYBN80fRAT1YtnfAdBApOToAu2K2Tn63v4eS4aWREhSRU6/MPO7MMDOSX1IUKc3KlCAP
BFuMFvt4eP2SFy3uVwbDfRYXE36iO/yBdzMN+zu4sZrx3DEVedBxtcFUwk1H2WmOoqNUJr9nu2Xb
BzXOjNP0hkNu9YTet+nH1PMcFz4NQlXNsDD5yfdCoevewXi3iaQrwLUp9Uyu3Aqe9vr3ImsGhy4d
9cT7bzAoDfwzcgCx3bGGgizEIbXjGi80qjxGEVqr8aOJiMMm3OBdXc2hGcNArSpTzcl53Bp4PRbs
PoURk6s+ccS5Go/WCwnJkDKxUrXqZGKYaeFlx8ClIvMJCX+K4j9Z0aOc+8FB8EPu7iiapjoig42g
XVI11w46nT2AEE3RSAWa9M65QfFIi/kmgCR8RYtE99WR8FFLiP6BsrdcKFlaySCC+VPnL4W/kZXH
0sLggvgbe4UFI116wPdQogH2wjAgN/RvzERuzlROUfi70eEAF/zaJvS4u25vdcHRN4hnKNUA6tfh
P7yIDMlQ39j+P1CXnVToJRaq8uRnS8RWyAndKiPlEj1znQIaBkfgyk9Ul1nabUlb4VFq3sRJINFN
YmkpVwgxt8lzh0mdJSBjSQJCUf0DcQPE5aHl9uDMlOKtaG78XSwJL2EdMb0kclxh8GTBFOL6fLxs
QCvHHXBlma6+QUY/yLDGYSITq2GOwzRjYJGrf1AnE5JjTLuoDgzbBOwWlWjzLFKOYrSblguXxMFz
P1ZN4Whvlq6nJl4wwVCr4+V8gSL6m+YJ9UYyRQGN26M/+4THxzPIKhHhjL88nl56szEozfDrnPfV
vS5LOs7gc1xbfcfDBpjyQDmnpeoD14AG4QPtGJVSmbjcQ1cTB9vLWNHW7yLXLiqB7k8ULGE4Dxvk
urcGvj24kDoLpzWSCOF7uKqqLTOE5hVwgk6hXaWCoOBVxP4WHxTyqo8uwGr0H/GntHciFCtDZ1li
uBZ2gjS7XRpRtdv/v0QX9M9eO+VS1a9RkorWXb+p9pqKMGFfETsZYBj1jy2ktE0gyHyQoy83l/Rp
DKGSrKf/R2wne9bZWdVFO84g9UAcU4XsMHvIrZ+wqMfFBVabAri2btaHKejFwyllZ8PRpxoKnWi0
0XckU8udeTgUt7ECdDs7MOhKBaZsfbegylols6dA1WqruVzq0XLm2ttYFtK1jsrBsOg+VdYiwRfB
VWKx+lgvcLElurX/4CCn67TGQqSNmb3nJV6m2FBR6PRjQYUQnwlgl+I7fohZLmnZWlpz+RTmamaE
bGGVulsiuB88VmzX7MPTGS4rt03A5ZeLLXvcvq6aiolgtzQv5ve8UFwlXxU2zcX+TSAlxTVkJfBC
3pI1eL5Wip9I7pUc8IQCp4Jn8FLiCcvU3lTyiIkqhkNdlCFFWlg2NyY0i+EqaznJqCryjxCzZk2y
XqZ7PKacPE19ts65pOB0StUavAY7llVKp+2XFT9OhE3x63FYjHuxCS/enAD84zEATF/a/YNDSCDX
NyTZ6HuMdJ9dSU7wr3ik5dhM55cAGcAUBsJK9ndarKN7qgptcAH7AoCa7osi7hbIdqexO4Rjpr15
X7Rqnb/EuEBrNX+7kYJx7qQ5h0ngsoGfDIwgFZwlwFZanztzvD9yAsS9fpiEWWKGlEBS1DZXkXJB
Ep9UNFLOyclJcnghrbilt5DL9ksuCD2lOAjUvkzV7JR/cYO0m2Uy2RAD8W34d6GYJC8dpX5UFFxL
e3HAm+/xHXYx3t04rBfrjwRcGC93Qvt/pLEifKNq/TTbvjTsINRM+uoD4e5KXS3giKf4HBLgW2wJ
46iP0L84fcot/kphkq7HWEoyNbx9WuqJk8Y5ep9n7iu/pyADf7Cnv6CueAtlPgoVGz+wumqJ4J+Y
IjEpkbD0b62Pj5GzXn2k9stcVcQvS+T55n9VG1kUxDScKXC81MFeDMO1TemznJw0Cqcc2M3V4lX9
hSPWvLF5AuKHWdPW7i8igk4CMJCtFZw6wpyXaaX1l6kanqyEhPa8kkiJPExtHq1DXProHfIs1/u9
20jTs6dRM0lo6+vSGhll88SsBRupERnnXBMxoiw36H4O1uZ1Az9M+VMLEfhPeEXv/k/Bv/BK9i6L
MYbZ1FpabA7qT94amjscqYYHTDXGZ1vpTM4iO6BjjwIpWV7rcIQruFTo1y+Dk8ANNASNunR1LJkH
D17QAAt0rqQox1L5R8VvjQrHpneGrGagkRerzr0HwdyOGSIviXoL9vxlgzM8Xm0fo1tZNGrJxzTB
CpxlpPIV+RjCNacCCGkag2Pn7q04xsSdLyOZOPLhTDeDaK41lztFxld80p9Xrrcnjrv+5yFDP9Fk
5jLAtI4V5gDoeSi4cHvBQxSFhRsPR/jH7a99ZJYi0pxoJbtO9x5XpM3fKQBYa+NIjIxjWGD6ATLy
0DeXhuydftWrkTrc1VgqplT68K/MSFFMVaanZOrrQsC9Kb7PJbNQExNMl1x1XxGb1H6dLAmZzhbR
h/kRK2gSJq1hpJ7BxUZMCvT8mqfFJMsFbCDh2AfBTUpkYy/+SXIW6rT7N6uc595ZR6M322SmF1Zd
vlqteaZ7aRods1jxNkmOJKblaXw6aCGLMMEK5h6htorBjZK31jXO6suSqtocEN/jchnE+fSBYKzA
rFXz2c7uotwY69aEfLZFYsb0cEL8GhygAZlYmzxpo8ZrturER6IlpVemtM5YDMEd6aKoiZ1tIKEm
iQhr+F7RML0bw2VA0VogwUkjeEdaMEg05DiSZqBVjGZ8XwSnFUiLABXQbe+H2L5mWmBaiiDOQPCO
D/AZlkC7InxV7yEcNna+pMgIvJHbEj8fmW4m+T97txMPTdgbhmXwC2bkyV1FonPgr1Z9SyKnUenA
CuV6eXVt9GNUYyD2MGjmYhuc6yQeCDlkVrGItwqZLqqb5LTwohVq5/wPlBwpES0/qFbq4p8T3PLJ
jIBuUWg7CLQ3pzPZ60zUIbsmh0ZTc8Hc2vEfxXWINjMw+7K1DIAlvhKiU2nce1PGqINEPhOPRfLx
qhBlwApoopHXMwobPgm3j+Xrp55l4d57MYsNcXxV6bjjycZCiRzMK92h9c/YBaKtF8TLwG9Cewih
6cvpL5HHX0/TkjvjSlGOZeAQ7nlBOmsjlqtv5ugQ9stmbeftMNNkLhQTu7/kccJKXsywAVhsvf/l
FMHqFISUoWkcxWr61q/nv4FNUJ7BF31fbkl2mr6HXHRmMS3+tTH2Os2qDkJ8N307DDcjB6GdVmvK
sX+w5oIEATRDr67cnvp5yc0n0SbEzj9ju3Egr8dPXS2WdQwlwdn1FZpL6dbjfODj2LYeCv9blwWC
Hi6IrIJqnewlNhBaqrxUqwzbEgiEd/mL8YBebAcjF9kOS1jGhPf10qm7GImhMSTaiNNwPdBcVsJD
Vh4mJw0+zl4zoDHc8bAv1yylW++IeCO1fIuzLrWaKk5kWO78RDQBmT1pQITlufVu/lJfL+S7etc6
3ieBWz+cAtg3Hr9hlg1f9T5wg9sxGi8rsXG5tBr/a+uTR4xmil7aAJiqYBY3mp+2PFF4bgkZ2FR9
w80lkaJd4X+FpxceSjHIsx4jgkYNinVaEYOCquE9Vi6rq88immZXaW+DjDoj1C5sk+K5sdikRH+E
ApfGoPWRYXOereGl/eZ6YYvrcwIg3GKgXsGO+ayPR3+dqJPspaFeaT9BkXvf/91rKdWPd5ZT1Afx
S8m7GuNdZBZLgHTPq/M9jDCh586Dbt3inyuuTyZi1tdCQFzAaVckfoaNxGkGj2MEMyAv0w+EEA/i
Cowe2ZomAND/+1PzzekpOD/Ym68Fea/586j8E5Db9XFwhIxzgNr564cRBZK/AcFmX2n8E8ho30RA
0ixaNLekCL6MPAT/S5PjkWk1PHR8QJMDrXzS4nEyi6cEkDYoicnq1rlAbm/CWGo7FOZ3TRnTtY4S
vcxtqfGF1IYXMCN2Qsp/oFBni1DlJfxy5fGqM1/XGyoM8VTblVHLHRuO00hRqIjxy+AJod4rsm1b
BL508YH7r/JS0KrV32keja1gR6biTGKQwuM2/Tw+I3XfL3hb96nqaliyl6uOFw0n2+vfpthBKp2A
iKtV3LHDmy/cHm1Tsh04nAY9jcUkPVexeKhSxzBUuZuck1bu+6CKBUSsajXNk4AOQOkgdp8Tlt+X
V+Xiu38oi68bBjSvGu79Capee+J6oam1mYm1BwUZnKl3+E8Fi2FJozPiumyYfMM2QbaBefg50Rww
opoJRfAE96FAHewnqRv7jw8HRs6aN4uGkUb+nkI4LNFNb+dUvaSL7ScpFhD+39qS4oGz5mW1MzCY
sWtIkBuTas3HRsxOsHQWB9zfW0VDPK1C9ISL9mdm1gdHval5nsQa899KwOez8YWy/7zNPJVmmKIq
d9YyTtngFx1hJIxBUpvdGhGxZWKAdEonr7V/TY7NDUVpY0RpugVVsoajIMBYio4PCZRCQ3j092GS
DEtkgyadVx1Hbxevs5UojsCBdGyKjVv52nkgyrxM5PrUQL+P0u9rblG95tGJ9wy6KI9QE+oOALZM
TAKWIzZKXUI9CUyPUD0VNCNc/yLvm5kWJHffasdSGuhZWm8qoJztfbqbgUc+dUEtoNaFLrC+pN3S
f+H/3rUfuejuW5JwfrqMYGKmrJbYrd01T62qgGQ4S4WP/1BE+W3LGbqkI+tV8WfLuZhzGVkvoesX
kQkBB0eerUbGGzxI1bb5lzWtvWOM+uiJjEfgYs1Wf9VsotoDK+prcVxB79DhOGmN++3uPtAG3jUR
+cOjH+UScXW2GwD64fbmL7xYLoVbSGfjvDGbCwn/NrBX50FoxJ/0WCFCKxHNNy0NFDJLo73m0aDt
lRIqzjiEyw0mJ8pOrdeqj2/YdniiSgJQ020ixANcnwpDjDbpnCuCD5u3SyZqUt8NVMGMAKM+gRVY
jbeLnIIHsj9KIpbdwydgNYwvbsyukpXxVVQfor04gK1Ag0SSILyAaM0YbGEEMLFtl+WIe37jKGhm
tfprAkpwQ8PaEnGGhmVnXxrIky+p9RgBGWCEMzjUj9pU6joMVNISfCf84NCxEuF9mJxj+9icBeZm
DfDin2pS6eGYu6h8xM4lcIjHUF4eRVkOv1B0vLEu0xxHj4HaWzZ+zrRcWfYed2yJhw46WwPdZXyi
0Ey5cpyyjfck2dyuT7NvF9hbTOlhJkeutS+xOSM9MP0dUl8EBY+KWSDOaIUplA6YpgMJkcNhy7XR
5r5UCIIs1vP4MHe5S3Wv+8ckK907sG1rCj9G05upVJfPS6jfXiLAKRSCEDa3X//Ht3708E4pxOM7
tyqu8N71nFq/BmSxgcsK7v5sKXVre1N/3QOCw2PAAKOoyQgxHocPal0DvAAnpC/r64Y3yMcpZBPI
80ojpA68RjUP5esNzP18SBw08SYENTsJ/GO7kfpxtcsrgjxDmHxETI5eTtEkUPxH7uTM4TqBoMb1
b3mV05gSbujYQ2o8iY1MVZXIAI/b6JQetugxLL4feM3n99wimytSK5jAc2Vpo7feRL6QsXdFuliG
YhEOAvblc0DBDgnEmciIrVcHSHFblbTBJ/cOYBPRUkY06/VAHBTqRGBvy4SSMvF8dbSzmIItY0Cs
BG0P9kgEDJWXZ9/AY+UVQozyuBBC+oC7+caICRei5jx1GFSXr6vkJJvBpPHvRmsxQizb1Qi+KU+5
DVRkrnNZ3dFgmjRSZiTLN9HL6hvYwNfTTbEWrVeVXUtAIp0fEHqDkU0UBMAr13ac4YLFtS4szhcF
PGRUdeLrn5ibbPOjFCVmUJRAtoKPwtBMAZI6R5p7F8UhL8mHZ3yEBE7HuLorp7k9Ts/qw+o4qQ3l
RjLaFWo5wNNvXPKduN+Zyicj4P9KFYeiMdgEc4L7wrXOLomosHa/2l/yg5AW6A4lUjS7EbBxmNbk
HZOVlt8MBGIoeKVOSqYr7p6/D7weiPdyxPgyHH9hN0myjEIj27m28UmGhfrhfoOKaVMb3jXnhRDK
u6q10LAWQS5EKNptny7yVTfdvqnukY7OMmGu7ES+mRCIK0aqAsIoX7AostxXqwKlStqfhtbZRzEU
ZcV/cJMG23oaekxw4+dpV9hSMtH7mAX4UPrVL12FQS/2FZP6cwas2nxmy/Q2JTL7AUpFvxkTXLTf
d5kmWrIwxbXrDgSKKx6ilCpwylmK4rRyiCHkg4VSaaB2M4V4JZHssabDSoGDwPrOV10ksRLhoaDD
jdCpEsFMKBHSEo00fQFRSk1ift1vvwS7BUsa06A3vyAnO7IRbXsP/b73F//HMwYJET1eYqa5dLtY
7sMhViwSGyJF3RZQvTP4bxC6n2gsg0HCoB2Amtl29ifyKkNQOuA4mMgUgBiGLYL0R9GJeXTwSBqB
5lgd6FdUj43sJC2swljnVamhKV4fyN7ZcBuwR5h/FxeOJ8zLSmtiJcVWSd5KvaWoDuErqz+MUYyb
RIrdZ9y/LPY+5c2L/zijrjPDh4rh1Po3Re4oPLy5hkN4/IssYpuP4IxP8rAzJvj5yjX8kXmk8jGI
Ji7MxuF0XmPkYgOnhtXTPv963pGXjfMUFBN3ofSgsL2nmW2uyEOXpCtxpRm61S5hMQU6BCBxoGTG
5k55cuEHArdUQfkY/Z7fuQkPTl5GmY34L9QQonCII5s3PcFm1tn/WdeOpx6qjBXYAgYHwVnrekm1
IkZ9VoZzLqrADaXa8EgduvMSKJQNerKsBHHy7zJc68uR7+eE5CJjpMbY9aPovpKsBWeuquD5XXnm
kuDkDhOgyWUff2azRbRXTyfG/0Pp4DlJomotVh3NodM9Xqy5r7pvFVogTQvkNAYTnbNtzBK+wCD8
GtJye9SqLKwEaaB4JTmQvXhrBCoWiL+Y24KDpzKfAWvscN4+YsDMqHEMt0qsNW3RLB6KF26DeCMm
HLBriisSDVpl8ePO6W+W90ibqVcsFRllsqUVT1dlkb/ho4lC5OYjI8wpWMIeZT19xdHpsWDWIL76
Uy28Jvi5S1giYawsnb7b3woqTktcl2BSYkzBOgrdIheyzfkcCjVlSB8ErzEeTTE2OwiGh+K2HnQE
0Dv+mZUGOkE2CB9WsrKOsxSsVL8TnUJLtIi3wPARytzOQ/+0YnoU51OkmixSpPJfrJuvyJgM39+C
k/QamOy2RqcRy1ytz0mS4T6qyWDx/EllOo0ELV4VOyvOm+2cOu7e3Tg/OBQK7QXW+7sWgXHYPHtU
Qz6iJudaaECkuWWn/fLsvx+Un7L5LepcRi/s9ddoOj4sUiOehsRvdCr8uZqNIc6YkOQPqU/qZkfa
r3Dn7DJiJmJSBviwsLFS1SydU0RjgIWB9lqi90w+YM5IcnFz+pIQ8C2RTB/YxuNWgMR1D+40qhYY
iVrUBwazWv8QVCOlvlTUVQ/vpYgIFhQxonWFp9OOo68BgWru7HN1vsaZU6RZHClAOBcCfZ2VyL5F
GVgR28yEPdCrVSmL15aQ31g5D8oI7W6rWGXjY7Nx7Nd/6hblzC1tCfDE0/5X9aH5WxwMAR5FB1Eq
L99OlqUnUj1qp65ETrYRb8BU68oiB1TPntYJqLa6mt8SQX+4rJoA/HNV3NzWc6kBn3u/9cSCQZh4
AJLndigQUA0E9pSpAOjOTI1QCfujrL+SDvCE9+Y5r70TneMhtti9+nHoQxinOcvdd4tKHhSQhNEl
K4ppCMWENGsP79oHYnkEJUMBQGmi7yTSXp9+4rJGSAOE7p3fZOX5ycs3AZctVbS0ZM0T03zEophs
4evkQrjsQ2F2kaky2P5lGUY73pb2ADs5lGkwN+WYJlg0f1oRV46oJwYKs+VY+/mQ76SLh6ohPrGQ
OUcbBo0mupmzWv1rXG8OK1pWBAATHsXB78LXbcWy1NrTXL/860B1fs3ZR+2Zustg2W7czaneu06b
89MtvIZZyAcLv4kJb1ZL5w94FEd28Kb9XkIeNpU/bZnK04UhfijlXj9p3d6/IR8070+XDJvvpC22
Awu92Zf6ueC0uEb+ho38efmFs99VGOlWKqDys0nH+4nY/4iSYxLNzoZsoHT5Nc04IMQg/6gOivTH
KrbWtmV+wIcEyAsjgCGWKLejpqq4ihyrGkdif+4a4I6gKj6ig9+dYL0NXYWt1qHJrZ0OWmyOMmQa
smcCqFoJK9KfWXO8T841Gom5rcdZZkYigYypY2rZQQsDwGnMU66EudN5sQzI+dws9ejnCTXmIFQC
kSsgVR0fOvbVHl4YVtQLXeJOZqe8zeMe6dkaqDIjOZidJM2m8S7F1ZpySd1jOgTxBV5lcpJBXNQu
enOV/TbsDPPym6bCAmR61UjYN0OpdsqAJd3LEvUcFrBzJj9eW7Q9CtiY34doR6ryt5rWWixGQa6r
q7Bx1iwR/AWeWTRtyTlZVFp7izn1cZSQaH5M1rQ1bxQOsyWi7kzi1NVucKy8pikorIt1nGiGPTUy
E4/LJ3HZV7g0V0dURAyTIDWlPoUA3rCbuZhVoSVLNCaA58yhfIOxxGstXuAwe+aXRTEyyzI2sVvA
/YTMeoS3k1fHGO2NwCJQYLoeUxlry3iiDu/YO1HXZoHo/k10lt7VlBv2yBFuDs3J9436Yp7+huWZ
3JbMwC/KYlOtZfaxBLoC6x4yhHGf1oN02vAJ38oX3bkxNCDuh8nd9OoQ7j3zTpodd2I7VcAVAW1D
W8fYianPZ4KzqYBxy0S3237KUbHYArVJulJuUcNk4MKKVBCKl61rbbALdA+9F0QB7izJ8Av3gQG9
IA+6rj5opTP1nYWRgepW/XOiFDwaUtAfJGl0ahRSfO54RgcwqmpbPsagLzNZhVHDlS+E9Ofwop7n
CoJXTyy/2BRIde9ybktdC2l44S8jLPBqSd919fVXOmQwSuwrcTg997Fzj8fNgnwy1i84tf3u9Y4v
BP0saw+35Xre6NhdoOLwvrpUF0dWbCw1Q/prOoWdAfvATivVe72/GPFsAHtqI/px4bTEsMLPWm8w
Wgvxf4FwI/P8Ud0YF4qXeXnegHTmE5t9GfplgaIWEA5ZjFUreRmgqnW0VLzdCZFIWYUAvFJd4ddQ
TrDxlcriO1jzR1E2dnQgWxHjQ256fh/gAV2euy3UNGr2X+kwH9hDC85otXBviaPc+OZoEeXJHVEs
Sb6rXsY4yM03LYJ2zYpsla3fK8Jr/+eCKCfSuBZXw/wOvFp6xmc93FjDN5ljUIlWaxtx/NS6ETvJ
jmo2GAjnOqJoykfntpH3SpH9yxjs6wTOmQnBJbHVyuhd/sinwA4XMqsEwLOwrE4rBwSxQ3/kX49Q
BC1LcsvEUO4NEWIFn8Of0CH/a4/FYtqGA1udcmrc7xCT0KT+SiA8Lvnw5NvAKmlaUhO21wlalpEe
qGc8h8Wb5wnNP9R4uw3b+7p7gt2BEOqqxG9LpmgjK/KBqLLBQ/Ayo+F9lfDqCPFoVn7SiIP3azzC
FoKhXy54XjNAOvaTu7bmjPAFZMABBVkUP068uhihtY8UtxqAak51dk8tLay5papQh/igdvXUas0L
DQBLfNxAQo4moevKltScJvQq2bNOdb9lWAF97W6p+FrmpCv2RL4klwoCeGLL7OGOM/hcXfQ5yyXH
LsNruxLNnWTxf7sOhvchAv7cFj9/6TpNXQZS6HARb2efhtgcvJZ1EcWznthdWA4DTXa4jkn3rVVq
+YH64uB1nDapGx/DzCt+cGvn8Z7ZZbESSlrPH38DHI6BrccQb5eoRRxfiVf7vn4jO3tK3hNeNbJe
w0Lbw1cWHGUmLtLwYfAaZGKDUl1CfCVR0rnOmsQANSYra9blPlLKkYw3IV6LiEGunELl0KZGWsj2
+SW49cFY4Hw+fMKB1T8uSRHK7ZiTCcjEk0fmLIliiXhNbhS0E8KMNY0a+6c1MYamQHMtzRmd22hg
oyJI9E72iUVKkBNopZAE863lVl0RzzVNtQZLJreCHrMQukm6Ypeh7kGQ2dn+dFlvkRmlWL9L/kV4
bVDtOjVBgvehZokPiArsD69PQPnlD6VWkLtjm5hSnMUQKuv4ZehKkntiJ7fKns7jcHq3GFZEJyVa
7bh0PcDiH6U42B8m+i55e75zGLbXZ/YVD3pnu1+hjHxw+DJiV1Np5ZUot0zKu2rqongJK1hhaLaO
5Q7v4te0ls04iNf0bjmUJIAxEqEF24C8lJevix1wSXvaihTEde8bNnGH4GK0IPNq3Jw9nRgf0Foy
CWqtCfZjB2Mlh0xn3ezdDbthHTy28VsLgKn5GR32xBKEiDFbh2Bd1etQfRlJ5gC4rrw6O3z1vmh1
p4HZIZURfBEKASG1t/z6NOhDF4NOUJa2XkZxtyUzffJ+rDfqf1z5oQUuHUMVmmc9QispKYM/WGVI
FA7P8PT5qBtLYEKclt1TC7fG7YGhAU2AeXKXa6eH6Yc26bis8w9R7a6EIOlEKXhqB652a3qlc2Jy
/whWMcyJ8ot7Nf2t/coH9WWZYhcJm2aHCia4wKnnoscLcJQ2SplWCk6TB3TU3CG4Jun5lOI/YtJy
gkID6etUAQbDm1qANC2ZhPbaZtqMtA6zzw7YLJXqEIOtQkZw6k3zHmDj+/f+X4ijG+wn7OcBWetS
TCxLszfZAQS4bocmEfFnAQ/AhNsaiSzDJqU9SQlwURwxCa/kir3jw8v3EnVzEUDcnhxZltjau6q4
9fmJi7ICcQ36S+/vGEn6T6rl53rICQKbRce+prueNo0NAuSY90riIZkf9hsBLeL8GYrOSBqI6jX/
ZGX/E+hwi7bBQHUudCRAORvZJr3Ut+qg3MaBjttwyHDvspRckmPvgWvmM8pgWQQeE5ejyYdTMLcx
WDh7+vKOJnwq/ZuIrl+59XirYvvzpF92bqxYTdhpyFxjnQ0vSLs+VYZaA2YIt6QicMn8jrAOux0h
Kx7shLVhh/s8raahzHFKFaqpb+A3Mc/4ofoTEX2BxL0ufSWhNrDGHj2XB6uvfFWkKGex0Ubp1Yt5
6cbXC97F0Nwb+PWpvBXclulfcnQyL+htVarD6wfQi4jOO/cwk1SHygGrYmzUNWFbbCTjqjDwpWka
wt0acpkWkek1hT0Tqrk2h/xL7L3Yo68JRpbba1EtlQGx1BPA1NO3BNvb+3FgC1NPRWQJXOG57I0W
jG7dLYMN5KKy7C33ayxTGFcSGOL4X+iSl5Zr9khrYuS+T6V/z37pBE9igc2kY6NIAQsVY99CBdkL
ERUyG+NkL6n5Z4aPEpuSfW7Vi3sRGIK+Rfa4ZM6lW7+pRf6v+X/z2Rjfci0XnpMwlnW3edb0kd0y
GeLY4JreDz2xcsZMN+uhva9ABEFcXV4OfYyIlk41lKjvA41QrW6SlakrNnJiAJtv75biyl8N3E4P
9OwHKO8+K/yvq+PxudZA782bMIIIV+S5wp4OTKVmHLCj82NkEBq2KIiESK10KfI9ZbQCbdlJOgAQ
mIcQHWsDArWWJH511oQKfJGr/uOAf8yBzB9Z32gIB0jJmulkEOfBIFw52L5eHvEEzCqlrRmXRp0G
lroLaaCNP837I/AXjhBd8AVt3bRHXMYQec/DGTOH+ZIt0RJwHhoK6EwWkDKOhINT8OccMRwN8j4o
SKYqQwdWCTSk9ErBQffEvez2ZkovJUkRqWnUjbVOsV3T7aGb4C/B/OY5/kdKw9vMU/qMX8mrJ0Y/
mC/4tIQ4U1stfupms3vW4jGyO/DlyzTQlweqCJZ4UDsqPVziFmG1tOrZsJP7w7BZDoTJcdT9DhBB
tS/MFDWeUMIfpNMCmFPFTiZuh8dE22ADE42Qz+NV7MZv7/+dLrHJIAK/9chwZcvUh1jPxSv3tbaK
ncZ+vbSw4zMiZem2pqFgWBxYipQQO6PsDWqOKXYiQ1xpV4SzTOPQSsEsgDba5gywcYimXNutKZzz
K+wcMoJ+/+6MXVwt5OqaNoP62la0nXxshlAiI1nh3uXj5JjdD2afN698pRCJkZA8qhlvRu9/8dE1
D+S6w4/UIeYvzKiHpkeWJaiSNtgGYuV7+E8YGY4KKd3fkNQHxz93i7/Z8xA9tZWNfAeacTw0LfGg
JDVbSw0DW3/oD1T1CGBnVP8N0RNEiQ/NIH2UrTLz+DBog8kEMRI7pZ6vDsdxh3FZ64FtoECthE86
12aMPdZdUkGFDOZS73iljDAHqSpvugNoYfHWgDMbRdzMx/J+ea1a0xmh3xSHZgDUK97qFNXjA8cg
RbM7XXT10tJ6VJs7dnvREqSLwcRja2cy+vYBrbqG1Ulh6mox4/v9tpOd5GRKq0lGhsIlvQ3DU0kC
UEYElr5/iRmdELgdSXpmOV+umMa0/di/TUJ1qubhlgECQiDbI5MPtceDJUGKkuTj+DDZrq+BPY7r
egI4nKsmeGhOLxO49KYA6nm8s6M3WTp9m5ypOTuc8cyMUSVox01OL92nHGaALYUPSyLn4NAnjHJd
eRUiAUtPNlekZyQ2KtCDguKzu8/0x0283XgzCRjC2Mjxw58sAMtrL67p5OKXntt6MiNpv9aNjyQi
DnS/WRo1BNxr/hsY6Y7lQyIt76vpRizq7UHtMjF9d/Z9rzhSd13B2nHEAYoNf65snr6qJfd7FthJ
mU3I2MqYmjICkUJE3C7EDbM04DM33nqt0fyKdrovmZIWTdt+3POjX458tUbFQ7mBfVxIPe6d8xKr
zj3bgaPYFYxT3IOaQ0dTFnlTS208gWM1oUqzeiMPZNZ0qJ5ub6qfUrMZJcTbnvLy5i/1ZdvDQCL9
p5JiBZzd3iu0w3bc1OIYbW5GiK/VaKA8J+aLEDb/twV90YazxaXV5Y/ZuXJP7SEv1EPpTJsfVuHC
BgjnDSJLi3kgYUh2mWkuDitLh76fe//qj5bliFC7kEpHqMNh/PkbRI/wCgWPfiJN9J11WMaHkZ+w
7pl/MI2x4qxdfkacMj2n4j9aj6CKBdTZQ3Eu/MzJy/9hEyiQpje7QRadmpwiJC4zs77mLkh6yuVz
SdR9971psYKwC1s6q7KyhynNN3DsLXOSWQifl0Hq2HbxpTp6WxouzbDvdUL2rY8oJfPOF23QrtyR
zcJbr3ALniqeOxZJl6a4FghSRg1k4X5WazkXnK2EavNQDnjg4jKDvOoiaID9ak+9zh60cR8s7tx/
tQE2c6MbjBxMAGQ/g2b8x62tQkhO7FJV8ayAIEHT58FYY5k6BYJ8xI0QzDoPGmQQjD6PqIHg1ukG
VRUX9NfWORn+nD/F4jslPmdZCWUmgsYTqRPJ479edwTwFseg8gX6RU305J0Kj1fcxWa4Uvp1zIp4
8Efix5f/vGYHKqmgUF+j+AoxH8Oe3BbfdMbNEuBjArHETFbtkx4I1rUwzlfwrt7umLaryf2hsdJB
i+t5VcAbPomfkDGDKospNuga/Q79dcF69M+SAfk74UYRFYudDMKVm99Y2LZfSFYMdyBoem3jwld+
+wJGtPH1tpH/4Mz6SwlxEozdUHt+FVtuzPkFNuNc5/87N7L/suUMZiuqIjr5cnx76Kil9gyq2N6K
/QdFBx8gegE0zfVBsacvPz4d3pZJ+tQCgTkkNkck3cXB1fzgrschhKUaiTZQ4QnF2/1yukXzbAVP
RRFUgc6dLvNtbri1EfhCopGcs+DLn3GLhKsJZVwjoy9aZJ0jSVTWj/j8FWYRDxwEBi+AQx1b72q6
OQM64squXqcI4pzZfBZJyMST1Dqnt1+UWqhc1eixpxVb5M3VARLM2Uephq29CHoaBsgELLMk9f4B
NdxP6f15sAIxaU1SRM2grEf/8uJkShUVBZFVzoEIaS2npiZmllYULXjZadclJqw7fgHJiyMfXyVZ
7GRORfztv23T7mN7XUWzho7wsZBtQKqEOsMpAmuBMt86GCHd9XGan4UrBYWptP+Cqb9VT4f6+M7j
AHqhho+pIUu2KT44R94OMQDovfL324EClu8YUJenvMB5awGN036Kwe/NfNfEU+FgCd4Q/98D1euk
uObzSI4YleAM6UxyC9tQIDJ0D44Ll9YJO4m3njUBKCzckViJVtqCkoz2J7jsYJcbxWC03EcTGa2B
ukRRcBvaOuSL56WTpcPWvQZcxeci7/CGoK7LJt3e7FEYSsCYi78nVFTS21E4IX41e9g0P6/YiWXa
ns6ukszGhkzsTWEr0aPDMw00TyAqbzHS7E6D/Rdh6WMnczbDOZbfLL+c00rZ2KXrlrXz8CqMLWvA
nr9+pWPVrHUxBIV7hh3UjQhomkSxdqP4gdRYT+OrwQe/2+xxBsAXtT5bK0O4kzJaJumdczoyiQUl
Z+6DqcDrWcPxcO/RjxPxExg8hbepXddB/T63AziOXt9JLYW4WqRNu1pv69cpFuoOuR/IEEkwsmyk
H3XXndIWAt48KDz9HO3CPr3E2cWlyulFdTLVh4LW4h2bk/5m+KBBqQn9FEMbqmlH+Jp0G2mAK15T
3JUrxt2gv+UzAB+0arNbfcjXEOQHxif5WEiOxDYs1tofNbPNmnSKYhd/LkZvwuEvq3/JUDOJHxAj
IKbYYPvXLpPtM2WTxqJNIgxxCZQxhE0B4WmjQmWv7+sDYNf4HAeOju2ib6c5VBceJmAVj9sWPAOp
IVBHCtkzKYer5MJTfUJmrj4RgKDRk2ceAxla3+CfIlt8ckqSeq8lzqTHPYvkIV5UdgsE89MyiCn9
b+XyTr7GCWH1Mw7vzd71zF6hnWZ60rzPpVicA6DMC7pMis/q80SeXACOmvGQCZA+D00jJ/Ro9nml
Y0IyBZ69xsi+xeJu9KZ/5tkaKt8m48RvjkQ0VjBd1PaNV2JJLjs58ZyPNyzvzGIhoEswfZ9n5aP3
4SYFNOPZyewoiFBm5YJmbTuyxZlY0V7/rxeZVEEfVgEojHUIHX6YJ/603NFPHVjVzSTPbwH1HOvj
txSJoBlmn27MX5YBXT2o9omzY03VZm+CywMTwjUPWOF1C90VF5FP2iGLBv+kiID9HKmJbvpkYzU4
ELrgcLAwM95+YAre18q0VQU6jPI/mxSmZK9IPNpKwkp+pbwQrlh6P8UnKRxhKHdxxFDnAIZsgypq
EKIV5vM63OdEkPaznS7kBPO+3PWbMrh92Cr3t88PQSCa1kbikg3OdPYO9QtKeOq5ur/nHdjo9hDa
qLiq/Ij+g4/po8Zvk8t0qShK1rCH8TY+c9RwWPsVAQEdLxT6Rmpm59drTYbQuTV8g4jePfan7RRy
4RFikT3js/NTFXNOEv++PoprDvEWyKOXGuf0jvZ/2n0jw+2urhIYYWu3XliRpEjrM3wfNHBXLaWt
BI6uA5SCbQJXs5eDOZjEBs+f+60C45TG/u4phB0VZUhGA/KV7DWkT1Fym/stfvwfbJmDnxOE8719
OybGVNw6bbrMxIx7J0yjdnZhgYzY2Pyt7iTmrghwy9APIBfl+J82k1oYwr0kOwDyG0o0VmbiZM+B
t/k2WAbIb/PcgbHwCR1b3JrqiucT85nx+0AzLKhB0y5PprOt/8rRXKOSD1oK+tYGnd4xmPhmhWLI
i4EkWs3pDRvOh26gaYrt4u9pt7Vd2yK/hpNIuSibdFm5/BKhdSk5CbkxeuqpxPSRIeWyw3kZOG2C
J6Te+CeMUclRwNPn21f159z4i0RNrDpOrHQWNiNamZ1c5lZpFzvFiZtlJoTb0pQg+S42fbpl0SfA
8g+S1h0NqivNulPXjKmG1/qjo7p1/hMZRTJVIhpjUGsQqpFeHpsH7GG97NMVK8Izc3XoTB3XBBW3
VOe4LCKlmfyKV+eD68+ouORce03Whu+JbCM5rQZdPuLcIbWINm/cBH429faGmfhHzoKxhPjo2x3t
bx10nM3wu3e5jqPGCbd0TZaoJT6GCUS6mkJggKVF/pgoXj+BUkRMIK758lS53Nin8ZLNm+lDjmZX
F/tNB0Lb373I/vqsfOpbxLKg+Jtb23zduY24VkpNo+LDarZK1VLdxC9rvfGGez2sF3bQsQpB1L+y
s7+BgESz3tV9AiSSDPkcUMtMNSczbT2Z4JjniUNRQ/KAxc/bgl+xf10F1cUpj6zYRuAuORBuC95i
EQnPeo4RpwpLC0SfPs3lq/B3FSfbKfgWMm/qBAihqYNJKWw0pOSxiKKsVToNrW8krgCPQr3oYU8b
+kQ8Tn4w5cXmds34hh2siuDJ5WXz5fK899J+LjVzBgXHCukmL6CM91fZLznClH7xSczJGiPjrz9h
uKxHOcDeCTcS2/cI4PUyIaIGisOCgxucxOFoQ3XMoxMbDRZP1oMOSP/e1pr0kSR6JqaEZKwTn6iH
bow+ytP40MKEbl2gCbVhfmYAOsBzizCT9ZDNQ/ckAN95YDvpJBAzDk+++ZqPgp78PsZACFeDs48i
2qe67VwwMvMIC+ZoqFxtEWXCwtwCxD8mZQ5UlNAt19jg+Pv0eTNwUU15G+sC0OHweUHzPJgMVMIR
OJDiXwIF8RmxaacrwrmjSwYblxTIgC2PIiHnUtFRVPcIg/KflZTWGDW2/JHuugyNQAv0SX011nyu
ybYNmyQoMlTVR6GqI/KV5ZG3OZtdaa4f/pXVzbMJ0wBdM7cL0xskpdcBOXciOfDCdZvE+BOKbeHb
tts9WyZnuBO9KMxGygQvvKLkeKoSXcmtnfKE60TAnchChGEET1nIc4nGNgjcHHyWapuSVF3gTudJ
1jQpyYUZDg6iZJ6r0olQiUp+TRG7tuiLe7PNPLA1z5ZURakCyHQvZ5jtPkSbxP3NlT/4OIIgbhtR
xk/RfdbIc1eP6qimGqmDL1gY0mv5oGukx4yj416kyh2qnEqA6YqlANtr45dJW+v/QCP94KihMS/v
mh20bmnDb/LQwbRxa815T3u7s4hEu4nP7uuSOTZSGZy8sRYq3QxIh8JCDz1jKwkIA4/ENXyt6QjZ
oYkUkjRCmZDLnxG7r00PCEclpkqo6n1xQrQByhAEXMqn4htIDG35etvgMvcxWxdPMZiya97fz5nw
A322IOydPWpz4pGru2qXkHITA3rUJl9OTdzds8pG+xZjSt/CJB7YQLoeSvn+k/lsHBQ2ZCsOFCML
LBMOHNmO+jCvYENkFlYOGxsmkD/BXK0y1yPy8Ti0UxQA1hQ0qGghwNdoXeMLXJPQoHmfDlR8i8dx
msY2aEtyA0iER6OWeTI9hYce+5RWRigFviDPQT/bAIItijHn+2gZxpCBKBI//lJ3qp+A55T5K5VA
qUrWXr0uIzeuvawsSCjJDJmz+ARUSD7PY+DNPsHv7XyiN5hsu6nU+ztJ0Tsgqa8+CQ3de6ncA+E1
zZHzPbClCS5+Fy4vDiixIIGEHNfOsg7uc6Y9m9eu/UVrTN2jA3awkeQ0h4VwEcUhVGveHtzr1Zrw
oiK60vxEp3s8jinNZz4BAqCX5DC0nc3iAGsVHR46NLkii16vAnhMr6KUefytWvxpUQBZDTCBprvm
h3X81DI01uzHReiKmyeiCSCZWwS9scS3h/a25+EVSC30kdITcZPGurGiAncC7CfqtF6gkyOGjoVx
hBpfPmNkMfdaG7IOkaZM9MCiztqyGzXLWunch4SVGP6DxTCxeARc4vVlMG0oZVrg8L979hq2XYBE
XQZEusBpsEZ+2aUQrRisN10noDjGlY0RMKsSDPnDWzht70h//gO5bouFdXkm/JNPrNtaXxxsAkTo
J3G74a7NQgEuGeVipy1T9GmY4+Ka1EgGCUAGCfS4rDGiJk+vmz/cYZ5wjoii1J2fciqvJZ7QVvQt
lKP9gdrMg0i+haQU24M5uhXmYaLS3tHVtov76auwyMwlLZDht8d5l5pE8ZqZ6uKcYDOph1i0X6c7
RaheoElsBN+onuDU3cc9Qm5yyzQmSSqJwXm1dSitcpJnFvLnLzD+DG/72iSXuU5M3zssPDAWzSXR
CQx6vsY0KQkGiFfJwj4wdhd+QtXx5PkB7v4J7kGHGlO6xqU0qDXvhtI3XZH91BJG120T2Gi6cGkG
1yZpR8Ekk4kMQdQ/pi/npbFrAUjfT5LjjYgIDzM26Z8ovgClmgbKQURXfvmpan48O9l5ptmiHXYc
IgJh3EhwNJSFpQIcHkhXfssT6wlEZQSXyYNNvFKNKLIiW1FHiT5tHyqmOvrlHdlLD9q/AQQKTcsh
8Bq6qRvFU0L4wiSHyHBJeIPPMQLG+9p51lyO+RqLiOZ/BYJ2BS9/BVvlFTGJ9RUUD3EWYwuAK0F2
m6rN7FgvYuN++RBSQMVKbgJHRR02g2qzD/atMJTsgt12VFaF6v5NfbmyRH9+t2CvDWGJCactKwQJ
bcu3czDgbbgT7mnLam9HQvl1awyTy8Di9pryoBzIrGL/9RP/553aoU+1Lfx+czdtUj/c99cY/j5z
DcgnAW8QXFwMUkRusPGTdep7e07JAc+UpJZxQHdiWtbJHU1F92TU3/jEWtEwN2M6HkKaNGmCxczU
RnmaqYeBzYCzBZe6m/acF4A5gzY4cW/21S7zfHVG/TKsSfnTJ5TNlLz9qIeKiCV/jcYq45/Jhlko
4Hiqo3CUHn8RZ+Z0oQ22Jv14ba7X/TCfv9ZyRVQc4/PSN86nuF/HEkdFH8b54oiEO0HSISW6QQi4
dRMqlvZ/01Nxt5XHjXoms45uMIFdfieLBONTP4Fjvq+PKHjCZTTg99RUKlEqOjfXDeE1Qp7uerqA
AMmWukIFC59flo43VvY6cEwCeULobN2viTOUxMNYmULWCZ/TCAxzNQ37FA8Uhp1kgOBqbJvpE6Dr
s1+q+2WKUKf3e9ftHV29U0RXHi9Cx8Wbk4ll+m515bdvziSk5OOQZGGguqzbQoP2gUGKaX43+Kp0
OtRh2vD83ktPHxxvvqPVC4bP4+t1lJitdTVvoPcZwBxBJUU4BrRQuKJINRDM8+XPlLwNQKYJ7iJQ
X8y3s+GP/Y0ge1bnPHPrbL5U4ywrAlYCQsGP0mMAQqb9CjWkhctT+rYz42F3ynUsh1nArG6k/00e
vTiVX9Q+goomyYh2JxIEkwFWLh4OdB6f9l5k1EeK1K+2uShWZEGeDDnFvcadUFGIFey4ANDYvFIW
i6mmbf94p/WL1XMy0F5haX71xVKq7oXifTwptGwdYMK9N26cy6aTR8WrqOc76b5kw4Oh6nq06ENA
zWIxbE1B0luhhXSrnr5i9qbialbQa3ZBQU0S9ylE8yBupcTYCiy3sKtpcp8wHY4gUGgJAvg+/wvQ
8NoCIx+cPGddn28HOaIzZAX7Cx6OMByIYCSnYJ1eG6QNFdllpMZRXYjA9ZP9LZsL4tgaL1VMdaYu
RV7OLOCyRg2NC4QLG1NSqv14LYv2P5i2iQ1QebRN2pUfnAszAwFHcGRdXNJ/dM1A0kBhac3bz7Bf
80XBCfvGHqnTDeipXZFsfn8+9TiKLos1NBr9v2BLgz1S+sDV4CUNeyK4iK21mXBuiSnPcX0D+Meo
hbh7KpY5hq3+z2LX6Dx82b4uBn5Gs3Pvr0xcZQpa3J7KhINs204PvaY2TclqmE7ggqDdmfz19Sqh
R6p/W0dnbGOUAmYPLH3RfO17vWyHCvLIgNpqDAHfwvnxeo/kqwJ3lztTmfPkKNM7MEhKzENyATIr
KInPG8qrLq+WObfi5S865aX0L9EmofWZA6IC3ytHXqrlKxhTMcDGszG/X6SEvbxMULFcUW5AqN1S
rjtZRacB3iIynsY4WiA9JtaG68U2ohKoUtbXuoH5LMgl365hEagce4eUKhKzjSEFJg9UpcV2EX6F
b9XEfw1oxSdx2xBiSanJ5+XlpG4e5/BQkYmEviPcW0ojjCGBisViUC8BS/91X5wSzgTeXKJxjyS5
1YmA/zA5ks0YeDHv1RhKo17ekl5SgcKhMAj+O/0+662jVelMKcg0cneg0NPAO7H6S3g/qyKV1PqV
vp1D/gihM47z19YSCUeRKjSunDTFjNpBexjl4Tc7P7EVlPrc81tmkz/Hb8mQbBPn4+5kYvc1LXI/
k1UzbDv2GiTDr/01LWetfIODscNm+SJ7xXu+xUOX6J8F6dHEAxvDxjB3/F5krctvDdQgKsQqs3Pe
IdIOo+wY+J/kFPFHgwXMWTNySA+/Y5u0Y+w+6z1qwaytXJZRjWi7KyJh4iyT7QzLJXQ/OgwmIZXc
44XhbO8CSL926vMFl74dc1f4TygI+nh2XsLjWgrEby8On4ZJVxi7LuaY1hEEa4Cc+ey/fvI+LBe6
kZlnbZqGurwkm3GiCb7SjL1qkVFWwQ487I7PFZhDRuau9Wtz1MY0oCsEUDquMi+Fi/623yN2krOU
vhXXJM1OthrXZ1arB++rkJFGtODGgfhBfSz6sCm9xdkBSDl5Qe7lA+88KcoF+WNBczMXtMPTQXRU
NLaGy1vXTum/j9CTetUQ3qvbz2G/04F6qDKQsE0pWdiHFsb08u5A7Q6uT9jpOeJG74JK16HY9cKB
jLKfQwWLYgAe/rt0kKnKbOfQj6FQ16s/Xoqx5DIH5oHYXoGp5AwFB2rzmECxXu0v3LqATdAXdS1l
iZ7SVIIyfD8EHzgqGWLuvCtiPu8Q0VkYDYUXiePSGusBHcEf9BLk5eA4/klu3toACIKEmOw7I3ae
Q3kyjtnQbS81Mq6ttjYhoxhVs9QUkhOYMXWAKb6OCeLtXJfI578G96Emmeaz3TYMTUCuLIEmFbYx
Rz2HBwLlEwhcvk1f1ZoNNQAgVyBLKyaAIiMIWv6lN9ejYFLo/b18I7xx01wcyvBh/WdFPR91d14u
QR2d05l0dyCaE2HOp0magedybHnBNMBtdgTLDrccJFB3mU1aR51MYVdhCQHwbSUPwobCYAA6J7ph
DCwPImwZVQjQ8p1frIIg+uyZHKp6X+fv4x4b3LmhMF+cW6D3UXW2ercZLykV90mpSroPOzw1bsuJ
7omfpFVdGDX6F+Sh2WrjcYqWXK+ps5ZdHSEoEPKfqLW25taDhVF08VhRr/E1AL7Dc2d8HvM79Xut
+xHwtRcBShHiYgyjW+7epOB0Qpe2Alvbf649k2FB0jOjsnePhlLQ3+X50GxHB10K6FhHby55RCZp
KsG0kqjk1MB2BUlogIQAw87hZj2ldCpsoQeBKFiBMCOU6Et/Qw48gz3jAI4gWQ3g3TPZxCcmOE2k
thkDjMyurSQLUnLdGUSkqSfqCNXeFUqgsF0V0kAHxb5sQs3kGyyHgwhJX2BIOsnePFz08FppMsOZ
xaJULTEql1oUizTkoIA9N/rkipij/oz8cRYP13fOLRgpD/q1/u5aP3GKhr6+fWS3dFHvG0a2Iy8l
ci767J8gEAjc25cqbL1/JzeDgB+enPfGKPi9ajhggZyqVbdq+SthwUEaTT30Bp5OwAc2G+3Kozf9
lSfYh2hH+n8EJZkh3LK/9DSM7ZHc/DRjT5DRepsxu5FB2X36TJuJtgunObeIIcyGf+5uditO5hGk
p5c0vgLZPEQsvBaGpATa1h8h3jF/h3xZ+8pePWDMQGuPQxcvCmaGxlYtIc/jqGpfKwBoGqfFP6VV
QuCJAUAlw0JgeIXCWriTH2VSCQ8CicBjLjbV4RYloAUtP6X3wyPn2CewKxPmcAG7tb0KbgGELSug
+ilM7qCZn2fgU0JjcnahRoxxxpfoAndA7X4z4kRJnfodAfZq8UY8zNMfwy+KYB3RtVklyEe+/zqh
tkwLEk35Ro8SkUIssdWNBuSayD8ABaMFsOen5m2F5wBy8XUtDoh1Q9o/TmH9fkm+WcPBJ1IZ40Gv
xHuDkzivbJZZx1CRLcrNVvIqs1S6UPswuEdqv+gY73K/Hpm/uYsXkNdjBxKGaI6fvZ0uW4dxmpG5
9x/FGODfEn6eSI3i/YXrQ6RSYW75KMzMpMaXc8v67y/v6oknglRB730bU5LDfcO2Y7i/EFBfSmou
1OICS/ErlNWDQQWCDFUhHRJHJbVZXA4Ikc+TRtU4Q7BC5mCkTJ3GDfbreZQDN5fbz6qxnonMRrc/
qdlF6uHBp5j45CoxZNShsEx0tSILG25IO1ewCk/47dUbndLRd7zY3YT/MtamNduG7zs9bTe713Do
qycEJCBvz5L23Puu0Nn2hOvTW7qdWZg3sXUQx579u6q3s5RaSh+xxoI+tOz65jy5dgRUjtvBhiCz
w2RaRirhaVpGEDZQ2fPX8baN901F5y4gQKbC6DHnupr2srI4Z2E+QvMyo6oD0FUASInj7nY5fu+V
LRSmqlB28KLW27WGSM3AgEAICiqzB10jeSuOPeAvsuUn+EKXqn6AQIE2tpuSl48gCJNEUVeQS8//
vY83kHgNo9gfcMpWPGOzXnRM4vbBKtN8bhEdiIemMJgs3VdjREuq3HSDB++vPp1Lh8dFJbN0kFsj
RLSXTZGThthLzKb+xUqv9T1BU0TIVecsjBHp5HxAYAgmktvWoH+1nuFgkO3eX/9Lo6fTJg6YRU6u
pMRMsyfc1jYDHDXxKjVShjWADDiL5Ya00A4BbG7vB6kCDPf4qz3eUAdjHwHACC6gy94r9ssteAur
QMxbCpoNcqWeJCBGAsTDTNwavyfuGdXl063yMtgiw4MmrgitloRXsYacWS7Rk/6WmhBrDF+jkf85
5VQyhF7iHuzxSo5ErODVd0HMr0OWnJ993500VJxrF5qvMUNztDshagpPNW01Uxm6CLQ3AEHbrr1G
TXD+O0IcKz+ZPsAGNK28iC+1etLCneWawx+AAn7dAVBiLM9Ls33yGpG4pzU4HQzGKdc4lmdx0fdF
JUN4NtaYtgP9smi2pRJKgTWKs0iAvW+wgxsbMScT2y/yXpGx3/C0il3/17KBDoB3rYH36RX080sy
HyBoimc7JrRNtHbQyQInrt7XH66Ly+YLPy65ZetsCuSeMq/eflfDNOS5vQnganm0uok4S6K4Aupr
GEp6fdjDGsBzCgn2r3HaFRNFPrfybn4yYjlQmnLcpko3uL63Tk+dvpG+Y5dT3UdIZJmxDzwX6/BC
e5u8vedMJU3vHIu7pEidTWe4O2xrL1Eu8FspQdwaHs3CC5FAZzHX18NCwUpA17sWbSY0O6bL9Izi
nd5CaYTbYY/c/zkqxj8uCLJkYpGwU2oF5+XdsZvljSVsiYtqYGXydP6JMHHXMeR5fSAF6R0uNpvc
RZ7Dcd/N4ERIZnZB6aZgS7SG7Rg/QTVhlvTP4OXhWv5FDEqnzVQMgS43qZsg8uQpYA8nJT7d63xE
U6Mo2oGmZtY93U2xtkAdtekTCTqnZyjOffAp99RtRRzElcPTvkIvfGfx97L7VUUuplMcxgFX8BIg
i8zRqfaFmUytWsRyhj5Li6aHGAp5K8aG08+G79EYiGpDc8RZPF2MOkUntpfv+DJzZDr0J1Z6/NRZ
8tRtaez7AfstkqfWgPQsnCckrMsmrjlASyqie1sGDUyUcWjGS2SeO3tAVAp9eou7+wgoMIBH28uX
f8bqKPhED7CGjhSNIEHKU11cnaj/UGuzD9iheumrVSP8JEA9iFI9PurDt0L2AvytS9O49waAnHWJ
4rGjFPhjRN9c2iVxYrlaGPjNn5tS31PqSV/iKLGNbDe+VMLja/oYOjilaRK8rO8L2ski811zIxo6
znUawzFlMf/VWiehhsHGlcdm/pliaa4Pop1rsxdbXXnjf0m7fnqodHipgDSNe4uq8g+N972dRcJP
KvL4EGD21yfuuEiyC+T+f1xztKXS5sN8zXON6Illd1z6Ghs03rELMqkJXQCl39J0FbrojJB8oTM3
DJMUpLsos2a4N9Lx4AjXQzqXcj1ROHEBLxKRJ+hP8G65wAd3dtBI115wkWuk6jGka5q9sMbn+QB3
m43h1geouaw4isV2nBR7mWdsScfqNXlD3ZHaOEfqJKbuZyu4Pr2z+eN+ltNDGmQi2gPUm9OXXEtL
OmcmfLrnmcQbHWzTBqUw0jHk3mFvM3jZ0Z+5etGkzOITmdCHV8IAqcV0+1cx9IwLIb2U3XzGQ8FI
jdzHKvrd5VWg1EmGeYY51/pRKtITQaoAdB7Azbwf5zmiBWAyyyF6uf8gCjD+fVzC7Iq6O39DPwbu
dI4T6iExq+heu2IbbySR+FcZYH8E4dwikiWL4fqFXBxFggGkVBiy3Rz5aIgoLmG4VJPZcTiFwRNf
s9jLvrU6eglyO9xPMPQ4moXSyYrzIdAwpfghh6YnV+uIRWQlytHSe8D2WR88kBeaTOIQ4BWfKwnA
2Ry5rPhACIpJb5mNluv6rLE49nIwPLlQgyFdCi28UHsQ7clc8mdTiIzlogaPH2chmz1SqDbhW/hv
o4R2jWShvSRB2VknyhL7CHv2AHfCzcFDwgvqRQjuTfUvZXB7RQwT/PhwCzzNvk2EPkmDDw11E4BY
ZD+B+5MDNDm3XtZi/OjcGaIxoY8Cf6Jt+JMq06OhR5oNodqhyiFrUBGZHDpxM5DglbHnA6oSg1sV
tVaLjjgYC4yTDyztg5PQzln+Aoox64o+36MiD4KgC3iHjWsa2j6RpN+oRIQ66z0Xfr6YwRvUF0ke
/7aY7Wgo9UfDMmDYiamzgfT02CjkCzxg6RNcUp65lRE1bw99Y7hXja00I8fnE+7sSV6sRjaVYkdF
Iw8aU2J8A7IakKmxiKVMBz4P9XS+ch2hWUSHkKtp+g8MB9SK+3jYzen9RTVLv5lBlSx00apxTbY3
FYVBV6og4nX9BlFRSiUNJ1radXI+BWdMtsoyZXS0eqsh0xInseq/BQbky8hKdudw5dE2eq50FGSa
eWKHVQECbJx2iapBOAnSxg501gllTnAqT0+wsBscYHbjfAp6jsE/TLiOdRniCo9ZloX7glXnHX5P
KoYc+bFAr+SaVpXxUyQ96U4TC4FroaGWetDBUY28tCjGuKL/Z1VuQd00kjLWoLqaoKAI4mBeQPCr
rvfcFu/HWxi0gHK4WSpknijUF4tEzmNZpw4apkuUtHKl3DnxFqxT3aeH6kqY/QloFydnpoRw/zUu
JFHh9wZVWSnYXiOsZAKdN8Uum+fPM9yk+qYpG0X76fPDhOfC4x3a54nqQIAtcJOTuk/8kXvrIf6F
gwJeKrrUdu5+9eSNqZRtPHDcBqZK+9gWzc13HHYPILVS4Y8oM79cXC8sTOIk/B0hsdLEX4qgFGgI
8ZrP1iAPko+ys6xTo8mgZDOh2F+fYPpI7ghIJlxcIdcx7vLr+aB+9ykk+bY1bIUdqfQkN23zT+Sm
cEXcQ6rfWv2vtNp1oqtZb1r1x7FO1DFyhzUrrIU+4oXtHhZTjhBzOBWAHpdSl8VyuKgPo87WEhFL
JnzHX5ELVwovVeWOE8b9ffd/IH5V3ILTtbme2s36CKRJtU8WjCivjBN0YBIwcHhox4CcE0N7NzMY
aY0X/HeIxRL3tq3p0GUJSdNvOQkP4eRaMwGOXDPUK+TI+7NfklPEdtLpfCYxH0IvGi14BPDNJMB6
nbwGKxvIyT620KhjYUl+B7paWGXEupwT8AuKFvGmmaEQnHYmJICaZsQ1K1sz+0xsSlCLW6GMoVHK
ax6o9VqwaSyB6WJm9kJp0F2GiF0NLSDu3be4w0PpNlvgt2zjDhk4Etg6IMPJZcnpPCln9tMdPRbF
Ii6+HuCc159jmleYnzRfaibK5EEmcnETmMUx4LfmIY2xbWbubvLwtvfX3w3FyneJx1mPVsuzh8HU
H6J6q2qcsbVB9b11/KOVO958r0ZZWGllvI/QIpPYCFi4BWXQRjcO/4J3XU5JDpxRQlmMlgXV74uh
VTiyKWkLfl24wxDqUhc/4KQn0DszZtbTXCotUoIwS5Y8rUaaxD9mfUNpvDhJB15Jf3L+X7jgMzl0
k/EaZiTEMu3TLHhKMZf1KT+jYWP1co0kmQmebKk4DAALITxAFaqYqUK3cq4ywYfHDPJudlqmG04a
HJQwUFDt3h0WjiBvu1mxn1yn8EE23ZvJ1pvp/jOkrIK+Ah/pQ05YBrtVqNzx2JdvDPSSDKWbAr3m
AP+xqkloNcRitioDIywGcG4VB0IGsqbnhHtY/8goZupt/xcKdksnVbobE8uuiYncrtGnQWod+eRR
ygMcveBd9aaBc/17yveOQDYo4BDG9Zwp9l/+aJJNBN1UZlMdP3EvmO1YlzA/+7hosuMQes4MJ2jN
h3jH+bcl8FPteqnGMw995R/99YzmqS/qWxyUHvdpgyGvgHKaI9B4bTtV0yU3ZXsm4Ulv54vjwi3p
5M63KZvm/HQ4MlvS9wnNOb0mqOze4dOqARRfU52aBlSZIBs3trdfdDs7vSAucTzzllgQV+9NZ1Db
l1z4mo0LmH3/l46ezCseT522JZSTMi/jIfPeycZx1kmeYR4KIHpu0siYtwTG+LbsbtB8CxpXK40u
NkNRb00b2nUNhSchuoL+cZoT9NtfEhuz1gEQp9guAj2TDVJR0bPfo+ncT3tvkch0SENmfaj5NG8V
x7+q+Ds9KhU6b5G00VW+vMSqilvRsHrWEM6aFANzJ110cmNaNAe2YwN5iV/8zKmHKaAMTtb7m46g
Pbro5j4NPddDM9u8xVkkM9xOIGwsf7ThOgL3EyHQvwd2UjU7cj6Qe6hz6ZOolGAd7Tk29Vr1er6M
j9idZxm0g499xfZ/i0pVt2XhCo54xxgQkbDgV8JQmc+InsqBgS9hZ7HZKFdW3dUCFCkrXXQsv5Km
+VKZlpvxSsD7jjgZ96jK85RVIWfE01DJn1nuKPrbWNmij7zjdcZimXTlYj828afXUOWseaqX0tOa
ca2WNpEFZcic6aUff/FxyW7gDRNdzQ3qtksqGTr+gx9IesrV6NTlvRtEbC8LGTPSbJcmULSw0FPo
fG8yYSHPntQHS8KLu204oZSwsJ/60AeEqqhwPcvnRL4Ig6IdYz3w/FI2AYcBGjDvI9sbk5nSNxjh
GXyJULa6CiFUZuZZFTtpek3gHqYM0gojt015Lr5BdPljQdNwQmS8+2uxjs2ynrVu9uzq7wgGDDTZ
td3bPYX9AnYkVgkVVT+3nco5e56kNqrqRw0UImzW9PPZc0okpmTU0vEon4cmMxoQuhy4bUC5uaJk
mJCU/wEKggO2WFj98/lBnzECfo0PaDZ66PsDcN1cluPjuHHgvGuEIKHD6NYs/HJHnchzt/UDrFmk
aaC146hTYa/IEa14rJ2wjYUVYsHuZIYQLMScNJEBZetnMJaNpQ9KEXJ+1Qu7SlSMZlxdfud3115M
hWOAHpzHy03BpURINv5yqPKM+MUFux1TJ/ifqG8jXBPWppiOcr6C+WPtQvv2umLJbV8IZ1F/aHRU
CPOz4u3kzvtjhH3vlhFeW8fI3YY5XHGJduIhh1HFrbgyOHbeFpNZU1tuL/jdc14GAcLkz11RkmOV
p3F6+wme4tLASEgfWbCevWiOwMTbzsmdamn0MMQ65P2mkyveMUAPj9QTzFQE/tRQul5E4kIfkPYh
vDO+wbQhHSkfOF3vk2jkM9onx9cLIrFBswZa0XOKpKeV9SzZEjlRf6aKsiVZLbTnoc6srhV5JJ2W
MdJtG15TwjeG7ZOxEGbN+8liRZFV+3PGTnWY39eEJ+TTYfsjuoAyAXE67EKLgYVkhFzJdiocfWut
HnK/ZplPMWCmyfDMi2xfZQHVdVFPFi0CJ3K2M+MMo2N2UuHWIt+PTrL9nUBPr6jUoqb9DqZhdde0
yeZspztxE/eggu2Ai4OkP0zMmric6wKEAaFdQC+ib8Bx47jZN8uqnFkBvX1X0+i/CAr2GNFG25qW
ikeG58dKtBlpaS2j+P5xtEE6ho5LqhAj35laicN3HVXOJirmn1xlmfS4RmBvvEbVGetghAWNfxT9
0XSF30+QBRfOwQCU139MF50Ig7ZfRELoQVdQ13ExPhHxwA3aZ2hzSkPk9rk6owwe+pCRrheIektY
NXGI2jAJcfaZcAj4AhTbyuo7hW55zlN0+Ucp9KnXn7gxk/g2LsNN5GgAESSnVZhwLSwtgn37ntPO
lEqOuBLSsdbVKzS4rfZlmIIRfhm9KWcSAfI9eqldFhMJGKZUK4Egzf7hRZcK++3oZGNuEGOpjaLu
IwQjs0vSqrxodJVPzhlVB0dHNnesuedEw9HIRV87OumQ7EKL/q+zaZLfyJLBcmo411DlhnYSJBTU
8qO/lK41yCc1dgAdwvkZ+riicm8KLMFPLVyd5L7T4pXlI3z2mwZInuzjNe1R0fqeQIfjqoKT1ltY
zTj2wA0Ae3X9LdhJxcSzQdru7ENS7YJiC/zAFyMxefQ3dEnO4sdo+0iDd/q0OY+zlfzy0swMzsoG
7AfGzvLHzX1+dp2N9wAOjBawLLM/JEc7JWHO9bFN2ARvCad0eLNUNcxvyY0rLNGE8V+/7zMXMSN7
weuESsBLj+D9L85nkk3qY/qG5D4w+DfxZh4peyXj6Gi9hz+9iXAOKwaQ7qheA8Drqdif3V33Lire
sOMX6/MJ/wi7DR3imDG2WXpYXochZkd3GdwNMkBTfN/6nwf0VWITWEoMaAIkdylvopBXOpYOkRjn
GWQcUkvQlLMFv+6AjKIUdDiVHU5whDHxd9y/5dRuteTP0AdHl0ExXCTbsjuwhWOKUrNxKO6Sa/XW
//rnJKEcuCTzG1wVgkwXj06UHLcvfDMKE4fqxRGuiNt8F+6PHdcTb9FN9ULfcYvVcu1pLliMefV4
nB/avtLXk4ba899Fp2JGJPaSZ7q9bxr2ibl7dyB2Y351y3/JPL0/UGwfhdN67vY3A8UzZZo8Q8WC
5BHf1PkN6+7gfUIJP6iXQ8HJBEjjJSqi0HI527Vr4XP9l8GU/oqWgNTCwDrY9FlEsv6W4CtVcVFO
hOaJfyx7L2m92DZYjn4lHCvgr7YiUuCfWEd0GIMAlc8Oewzog9PFBEnzeJ23V1q+EwPYJEPdXMG3
A5Z52mucfjH03lG53juFpJxumMcpfmUw1ufWx2Kegm8DIdEFbxShOX46RBMMrBt8A5ejKT3hwS4W
FzZYiLApns8Pcch3FTeEqCSo2FyParzWntMJZGkh8y4njKaDQMIRo7UxgKdhND9aYdA0MMHRM2Fj
abrj1hJ15yEnXKk9C5fjyiI7neRS8/bE0FgccWvT24tCpGjVZSd/w3VjuBn42B6cAFFoa8t2hQ7j
Ubd+umODoKfhMy7+ftn9n1xwGgvF46E9QNugcp+z6LqpZKPzEFftBJyC1U3QTV0Ls0W4aEQBZUM8
OzgWyS6hxSCCMoXh/2JbQBcisl3uY6FqZ6f52XrSieRRs7b0LlGDku0ETM5rNqUyiy8F+OqmwEGV
kNvz2VkWWe2+PhS98N9cO26SoGUwFc2zqPQn4T0Lr08Tc9U5NBcHBlnAWBqrSyFyI/LMGl/zRcK0
D7hhh1CV49BO3TIGFWTYFDCkY2eu/ZnfZTrMm216C3v+IQhuM24yzA6KGwmcwSg2hErkiu8Snepq
6m/oFDhoG6n1vAYQc7cdDiXWse+fcUyyerR11rbW+CPj50a57nLNnL5O0FjT9RrHfZoxvzrVTNY6
WSaMuJcxTJbxvPGuW6uriKz+PQtkKcYoe2Cs/PnI8JZ5SwyY2fUhqbPdpAl9ZgeE8zR/7vtcaZMe
qmT5e/5JQuEBMBoKBPEy5CKG9G40x5BQTyckVTf9Ec24roYM+whdFlZZWss4A2x+8N4lD7fB1BPJ
lxooqSSl41BSl2C8IwBUYr3wRFrh0qSWB8oGfTT4OteER4/t/3bFDLpYuJDnIRalwe5QULmmfIQ5
Phtzju+AEmc+3pdR7WZPuEGMk4enCJ1mVnnMUY333wP1cd0sVSUOopNzz8JUFcCNB/FYkgjd4mUm
Nn+AfTuaq3s3axgWbLBZd7WlZO/3TTe7P5mN1F2S45b6nM1F6LuN+0msIuaqtQXShEMW1XAH7oG9
qeFjpvbu7EmwI+SR2XtQ7DRXSiGnSJM78iQMGkaf6DlvgH09k+rFI4ALpyxDavayYcrL0xRGcPEl
GnVd7jaTBHKaR+DJf6rR38zy21+MTkVQElfSG+1sV2HClb5vbdfTQODSsNsSjrgGonVEGYaXlZGn
+ZTBNExRPYylE6c6uA1Ci3cQ3U+I5VbnmxVvZh/6cWQVLBFW34t3XKmF4OQZD3gqb7nG2hyRpJUg
jInszcWtPxfzKHBVN51cey3dXMuXG1agxIamRhWsYvTb2gg+aScntwoRYqmQSHwSz3a0L5lHabZi
JiUy49cWpu0hCBWrJfNItM+nbkTRW2mt/BtFfegc4nxBSSZL3VKhB3OS5DFZalP3xhPU5oKpkRLz
U9zGDKR/UGse5PdpdAwk+j9II9OAG56SmeGudA4/YZs/0zqNCYFkGOuQ7JTuxcpOcMWTWSrsJiGM
cSC5DG0a2HWrGoxcGDMQ3UK6oVSTi4TMhi8o+lwHpRnD/GtQ4wdxKxsRdBtviAlqs73IbSfGuS2L
XbklsxeTUpUDj4vOX9HflaPBTcri1wq8sr+fvIWfgRHV8yqkbjD3qibyAWj1qfZATTKgeMzoHrEI
wwbx+10/M9r9J4xoIj7/88xw1iMPbZVUfs/+mlpBGA2+/aPcC3VMrK8Jt4dYXgHUoZaI3vbWEgvS
15/uQZalEWjGFxQKUFiFFXN7JqSVWgxBjIlhey8RVXR6OiaBdhsLM667sjvar0aMo6x0iXbhK/DA
ixRhjgUOOcRINe5V/g5Y3baxbC1vdDppNHsUrtp1NhM4zp+x+RdPNg8L4RUOXQTaSne05QHA68gH
EgHe/+LGsqlsfYfQEKDv5d2Ins+D98gjgEYMUcy11sjuZ2/QA7qjeuaDoaAVVfiIeuH0gU0w1vXq
XB/xRfC7Cb8gaUFgZ86vPvC5lqlyomMoi/hvJ1iv6uAJdPM3ffj8wqCP09MVH0r5nzif8+cSMmD1
xn/L/neMQNC8UtRvd1SA8mHDQn/Kj6OtNDQ0ASGhHD9+R5AHTL4yUdw6z0Mwi8MQ9133qp7HbA8X
kKC2QuiJoSsGZcJX3wWDUL6QVYoL+9Tc5aCC+1vBDKQ2+y2FZRynsI0v+zroxBVwjHjcYMOUDKiv
VddG3BDgZWV6v31JonwZ4eZi7KEevMrRTQKSSDIBmGKB+DG5SFBuWQ43AE64Dlc8jpepuCrcqPIA
upcmuoY0kQIxnFah1tQJIuDuQqNWTMUT/+AFPPGz2avjjPGHlBBMndS+4IhTOguqElVlACQcJXpV
bOafY5rhJOUuMJm0RtRaSBfDENjrj97vJpCiSpr8AZ4aj3Tx7H4iez76R3NQ+r05g2vuLyhND9Cp
di++rKCKdiqyKZv4HCzJW1klW5xltS41gj154SlTAxJOTDYh90COAC84YktvMTt9a0NXyJs4moFu
ynAqj68WsTMtZib5s4npeEl1an9b/ISz5MXUmlLuHofpgZDYoyPj89jOdJ+BwMIx+YMjIDM/kReE
RKVl4+q9mcaKac3nP1la/5iuAggbSG6vMqefzqNE+YhGIcyxaSc2rsdPfqZykyRugPjRNTqGpsBk
UqCtPe8fe/hbYqBhpCGYPqRB5iKywhALNgQDb7jfJu4pHxjfsjMHGENpFxtZ8oQYH8lpSWPlg5jt
4E4o47s8nlZYewGXDokoaTMw8+XhTEtDDcVCTmDnqG5k3x5APrdHvvHPvOPZNeIdxLqfOYGTBS8j
Q8vtKjFki7D4k5o2ERAaRWn6I68upHWlQ7OiQ7MeEfVwkXA0kjDKYsO/+p3GBAM1aTHcTboeDtbN
pASS6h14XFiBbpndsAadoy9+lEpE+X3KP4IrJZ0Qa1JQRQIshQPn2++Pe3UUkD8/U4lN8+as/mYs
CHzQlIr88AhBDrJVkMf3hxj4CRZoMAOkazAa1tYoeTfVs0hM47VsRPqfE27tl7IsJHJP+1o1uOMU
7VqO43eI1Yf/HUhf+lZK92Y8LedA4X7bsimI/tRwcbjq817FcZ98DbMq4FquuMA/Zk8wNM6Y+OQM
c4j5vVchbclUqHcjCtigeS3xFrJB6onEan3ZMua1Lo2SaoGPXtcQTC3ybzMqYnvfzxv0ZGd2dQUI
qbyrVLOhvhxDBwW7B4x6FPPmXKbVIbqjQEe5g6PAlT5iVRU7Vh1yLBsw2ele9y1g1OY7Fu2OsXrP
6o4bfTpfaO2Mq9OwF6kuSfaE1YQDQniOXXKBMhnh3AP6IrsaH96m8GuAx/pJq0s+ajGjrX/xVCbQ
DGaDSwZlfvbEoge1OQ6TDp8p+xEACy1Q3DG2qpXcWJ9ZMHfdCPpeTNdofH+UlwsdiO8aGgm5Uogl
Oa4t/TewDr0IR5hs1CgZmrKfnsLXClZgEnO9I6iftp3aCtfLX9Xpsjd1cUuMi3MkejoqrUpD2ZkS
lDQ2GdvGPHSuLW0FmxWW/luvuACfV3OqZnnwM6+Y5e5Axx9MSDSUdV3VuG/0yriT+Kc+H99Jlxex
+ayGac5l9e9sA0VDN8MW+hRlkancdTzmtQGupgFIFLsN9pXdu8De4iQ6VgeoPPbkCbz1zzq//vq+
G4BbXWRtQFe8WfJ4VHEG3DKXN1nQ9lFF5fe2fhVLMjvtGUdfruxlqS4d6anYKVdVsczpkh17YlnC
5W8Frd14QJB6lGCLveFppSsN/rq1IVO9UWMvjxXd6C2/BZAQmU7yXlwyaH5wgsqFqlAxtDma9Hid
pQHS8mHBiGU8K9gBDgNfJ/0St3JyE251TzUCoXT/ooUhmw/K17dj6wMA8Rl1W5IC5dH10dHdibXl
3jx4FZzCZSZBiWyB9DS5A3HHdAAiHrvrwaE7FhptGaLoZK/MtYTPNxvkjhOiLO4/t7ucJVqHoV4L
ZLGWLIScCT+wOf5Z7V1K9U38rDnVtfvjxrmZ+pn2F31LbGu3EEi7wrQVe94Dl/wbUDIB0WLmme+A
IPihcLbs2dtoD+5Xkv1gv7/mR+5Jo5Xdqy42tBa0eJv+fCL7vNI/Mim7YKA+HtX9aFeSm1xnglms
2tdu0Yqa9RwDbxXNJHtjQ7ogmCGPRQy1HFgdh6y2AicDu1M9h4m2YAGWB2+fGBXQLJqFcigOCNfQ
bHCeBk8xN7YZJPsasAzjzy0LRTJ72wF8XM45+YHD5dE9Qy0yKGAU/w8p6CX5wXc663yvHf9qPXZ7
IjHWEjRcffU1HQ4xnboPVzjisJRXXeYgskjccRN2Q1eEVWm/3csHlHOQuKroSaPHVPqARNVY/MJI
WC2p0OdbgOunU100/DChOZev+EsTZ41iFd22xDqHWSRweqZyz4/6eL6ktm1hc9h4nFLW9aolFo8E
kvN+WLpjiFL1a7r5OylRT1yu7HO2ur47oQqMb2OijBoLskbvpOoDS9LhTvwTQh1kQ5nE2YUQATF7
kO7MivgJJSRPO6Xh4mQdAw2WgCSNyD0ium7wyJl12PJ6KPqQJMHZtEtDKs87GnRvdbs3GNdAioUd
2L8tcTMUUuAo0UL9PKQBJl50C/zvN69siNtrF6/ucUVtCXdUpNcyd9ZhXTQKOS0e/bIuU99uJU3s
vc6MLhVwlIxtJap7ou/VpLhMQHIkqVUk6vBQX3k1yffHqukRVVf1hSjyJO36qhH35hnpWmjdFNsJ
5+W08DI53AnvPE+IdcySqXVf4TfgRZ8kfDQ0qFULFvzwyMy745dXFntsDttSM4qIN0+iAAhoJe64
Cu1cV5L6KPvb4SCQq5i/nWeCOSxh0rQvnl0UnwCMdnXMn5SHA/N+Q/4SsZBFJBsV6/nh26a134aM
RN8tgJPRp7EKq3K6/goxkD4g3mnahF7+kJd186pwv020e8VyPSwm0okCDwJrd1InHWU27VtImA+R
P7TmUppJCzXmxXaJO2y4+950xF0ku619ALyhyixFttvYUPUcwJKHacRAyOxrbJl12Z/2LbI6IESe
hu6GyMSAUBIz6XxFWGN3xhcSEEyPw0GqHkr/1z6sgE94gN4GK4ZWFWVK3G78k4r9dOcnDB9GCIyX
OshHGdSA8oC3vs0QNkgDqHNGEuNo3p2ws/UaT7sGHMUwJn1eR1ZlzZK+RrWTPYHNGJ8lm98CkxGi
sUv7zp3lZXpiP9As7gMvpotz0GemRCaLVhtBocSkM++9IRTP71NT+S5mv79OXTK/Ps2gDMj/cdF6
YU3rS4tM6NUc9NPRe0dynCMkf3Mrx6JFKGBgPEHmW0C1l6Q4SmDFg+p3TyHqgK7p8oXY7ZwEwka3
94oVN5M7LWb0ZHpICeN+vHUK2gM9hSzAWNg99TPxbugr6RYT3iq3Czeb9BPM2wRZ98KmDsr3Gzmy
Ayc4uVOlvCt9kV4FvoyoEItTCYICKw1eQ05uPvSRemxsiqP/nWLi1urmr/uqbWeu3rSgkpPZDT/9
uV6eW9N4BakE50trbCAH2hwe15aCUWxydDh49kd5nfssucVCxB41wtF8+W7Q1rsAyqN973Hgkl7q
bwL/19FyaojG4yp2bPnahSWw8fypNNgJIEXJEDImxbBou2y26RIHg6dIaKTgXVkWS8MJLPSDpB6C
cqlozgaFCKdsED/NLxDAx/g5mCndE8ExwZPKue9uB8DC1bUCFvlwozc5/hBc2K9qYd5GVZT6JNJO
B6Juhe38ztPJQrJ1dHMHdk6GVj0Ba1bfBUeeq3suYLftFZmJt+CMH2jRGG8/lwSfm0eqoN+SKo1g
qHKQjG9wk8da5xSHMylcx8mfDfGQ06cz94GfN2Fi8XT6t+W96Mge9BIIauGk0q3vYZdOBtimhbaH
GTA7IYuzpS7Ukf3By4Lw+8s/zpeAM3axxctynfQFyEe34ZIAPeyev6Lt4ecrqxBID34l89UiF/1V
a1VrzGR2cp63soJCmcnejv4AdpJZ813TJPmgKJTNg4HDN3el+osZot3j0WnsfqoMcqFB/47MHKXS
k7gm9t/Zv6ZXPHDxNBd4j3bh4ekcjqarHxi1cCbH7MAF/aWebvRamvUhWQFy6o6RdnzxK90m0vdw
+2vuOephhZX5hP9AhygO17v3IFvcoeYaFdYxuP9sMHJWDEENAjbAvXRw+bDopWvIJDdaB0OYvk4G
EegOnXzi6qe5arc+seFJ/4b2QiJNgq6Jz5nIE/cksCnTY5x02+vJDxKmmukE9j3W4hZ4OYKnWwKj
9CLtpZJXxHcCGQtFYmp5rWlenG7GVikv8MxHaEz9YlRztvTedzy4hzoEK9yixGxi1wNqz5dUzB+i
s/Oha1SP3TEe72OHvJs06C/AaAivbPG9619Pt1x54bh350tyJcfMEaEzD+8CrASEXaqpLEVC5hWk
QhQ+/9bkeTdquKvWgB65f8urMQyxpvwO4sGN4BEDDPFG4wRcdWaEjiVRScd6xbJHkrMxDWV/Op3/
gXgDw8OwHBLNXFXypgn+AOdkytvudFTBeCJcjVc3KboEYBDTN3HYTHgwTn7iouncfLLkdtyJzpWw
SUhMLv5ciNA/3HtQtIEajhI7nVZkuzJcE5KamlGb2/oPuM7lEZR49+cOkvR/iV9XE8b5UVZMafBK
NehzV5JRDYMWTdbJJqeU9UT9lG10m2R6xAznej+vO5UHXRe4WOMBOt77qq3EGjza9l0dlSN+uBI/
IyU2COKUQr2tFZOVwUqEpErKFmo+7oCMG0PUAFqi5xXHekBAqrV2jdSxQC3XcrAXg+r6NhKQcsTt
Xw3p1JQBoRm6HSGUsexeWNH7wbeqSUxge2nkR1YbJnaVP0gXRezIK0K3Tp6pm37Ff8VImILW3QSK
0qJdyxTTgqOK+uj82WdWI+YXzB8hJY1cE/h5pHrZ4b/ifMDAnCmBDmz0z3yfQrwfIvkxKDs38Ehl
ORLCsgySBZI+jph8VT2nJ6+0eb97JCF3bFLPzPqpu3RJ5OqlJSOgzOnxGGdv3V53yjdhSmTK7Ptj
yWy0xZXHrdo7zaBS+JcRULvK2Kp9/Ku5BlkZz6mqRH9K+BnEigRn8rFVQBPizGU/dsBO/Gh/o5S7
FmUI/LCHQh3Amw0a/98Kq/vgqbWPsV+oj4SAsVhe34cgmNpknNE2sUOFc+AW4o1UtxEQWnIrKCu8
wq3W/m/IPc620hXZkRk5Y1uUn+obIe1t/pMD/J0qkwyS6/sq8a32MS5vDSRjvzhWdFUznU72ec2W
AF1ewaAmwBx9MIjN3l+mxQUNWdp4qdevJVsY0dOlRv63KdI03oxRUk6UfwlVSB8kqNdqvul9Pq1F
LZUl44L0jpkhY2O2NlBNWzTM0lryYKrP4f0MRVuyQRSI/gyoiKTGWv1q1rqi/3mFHZJg5pnK6HOS
XkhIuaAA9ANLpbDrI+cLqG2rgaliJswJoYpHmEuVWiS/J5lIsyy7/F1WX4m8we5tvCIIRGXGOQVc
RHF7wXx9hL1yOqGRR2V6UI6/SOltrmyf85ChpDuLhqhTr1ofLuXqjdjgcDw9os7D0qUrc7XDGcUM
Hp8Pd1Tpsv9EtNAZdgHlScEiuFC/+Yb/B36dEuZ68ZYLEhscUcxmIwMynECQLDId0+ONInqpy7v/
1V6ffteZiI+jRoRAkdzb2P4OFtMG0BV+fdmFKO3SxspoUhaEG64irT4+dNix3cBPi7IcCcrwfBxz
Cze35dZvsGw9nGgFsttwhYHieIXkP1zKjcmaexleoDDDTFpgiC44GuOARzTHSQ1J15bg31jfE9xV
l4Wl23Ue39CEiDdeyamixdGDAYjYarT5jD8W7bi2rlbSlq9RH7TIscKwsBdmVjXtjODaS3bOVc22
3esdZTan+AzHlUqca2ETPx2RP9sl5NvtoPKRO9GRsoqKQm/bJyFjKhnDJg0P1eVeZjFUfZiKAOnT
LTbyConeCygFdBu6cX/0m2sxsYMWpxM4Jjfshs0RN8KL92BRpKRBvkgFvhEi8CVB/16OyU5IGA0e
9Wlo1U41Ip5xOnQp7kHjnnj3GZtFphCEaUesuWHB7uoVCPHBKeA2F6EG8iguN220nuZckb5J2lQ0
sUgBgdR4sx3QSb9DQ8cX4HQshQHoiYrTAtiveDbgin/61Mu89VYWjyMIlBu6LOllaujnn+v9frkU
+ykdI5rQ8n7mERIKjvJLVPCQmoKNYuV2fZCr6tPsqETc/qg/1Y3cGD807EKYOWT0ir4lemzNk+J/
1QA1w+gO509Tw/9VXsMwHyf1VWLdQsRI3jdplvrWIGDAAGvHW0kT8USO/Gc5zoUojiZKgS2wdmRb
TMg29UKeMVtzB8ozCWIwnzoH3cfd3GRrNitF2LU/kK++aprFYcOjywVVOMHptMwB6RkQDu4pd2fI
IErlj5rDBL6iPeufsv6GJqxhy1d2oTqFegkDqsJQyb4PvR0Hg4tFwfiRr/LPC4CobSduNtZGZgEx
OTum5z+gXJ6pFTFshD8qolJ6A2ClBD47RDgKUS/WvG3FRgqhvZ7XLNVbPdM4LiEzcxUsQt8HV/P0
NZHCeeGc6DUVER61k81jjdrmkvq2v3Yu3yz80X9oB20jCiClx2ooN4wMJTolXhVaFwVwTr6JfwAM
2pQt743Kl14r/BEbUpQFsFxlaDWu5N1tlTVgl283QkkaOse+hFrH4fh6K1n663w6toj5kZkIJcSF
romlG7b4uU4N6TgUBYwWWC/QIh6b1HVVm4zzbinUXx+BUoXOuLldsG8O84ITz5VcRPOzi2OpNdH+
ByVFqvsQ27UtDMMblVaVTK4hjBj0FAS4N+lbseSaz+CyXOMPYObVrc5PuhCppMQqUu/eW5jdpNiu
GuKQOYytgclZ0La9ATt+Cg3qJy/K9xJcyKjDy3TfrFmO2eJa5309FPmxNNYyukmoajd46Lya+nsC
60e7SVodGs9ZVGWi/qULn0qImpjmUXc0omOlndxxxcl98igRAqQgfj58/q1szn2uQ+XG4fPRSDW5
ddfVyimivrgqan6Oj2S3PrVHl4QQ4RX/o07AIAiqB8usCpB9dFK3GyZ3w2thDoDCzfBEp8kB+E/l
4Jm4kmDAAba7L+4Xtuwtc8QiKxxshfOuafvxPRFFpUT30xZN4CzXaC5mLIz+gSLJLf95PG9fYDUu
FSdwDt1uzXO9dJ/+u+8qFH1E0gs/Fz0l7gcDsR+mGUpxEO6STyBoZU3S+Kb+o2SJn4vujz/3AGLg
V37c/kToBpSQoRlj6Wjr/gebQa8E8XbvrQ/ExQ6TZPsBtw4+mi5o5Fj23/owiAF6Y/p2mtBSzGRb
Oub95Fd6LWavA+XY63ZFmjlGMiPwb4wtaCuyKaaxgVXyv5k1rP8FbhUIqG3X66nGA1xvCRD3nISR
iOJNaCoIXSaMKILBV1UNzMHZaiaTv6ADHsEzkn4caO2x/F1LWwl/pdg4PQkWP1IBpnekFj8EqNDA
bCTI39MdMZIpRmEdU1pK6uU1OxcYWxJJeBkWTJswlIE8sfQ6Gnyh8Fy/4q1ychsvPY/cXQ6UDbou
1/RHGv1nA1StBBftTqK8JlefZzn84AsfydB9r7gUgO1x3ZOjYrajngB0C4uylFaiPg09zt+2yEhv
V1a72DmRpki6M9qF2Nym6V2ZGtUbLE3mcL53LjM63PetX7Gpi+RbTMRaEZN+IyWJ15uURxRsJZz9
ZxAv1WHjIgtdDTp4+qR6+f0Q22H9OzanwOvXXAJ9o02wbGRUJwki67C3THJXoiH6gMRjspwFQ0Vv
lX18wIvQdENPaZdFlR/EEo/NUJg+VsAR9qYvd32HE23pmdZJnbH8mfRLhYON/3sqc4wz39fae/cd
nlwuOoaUEBNuhO7KgJToiYFFVPOd1clCtDMpUcZ7jSFIPpw5QJFKLIhiz1AWonxQDfWYPE5ucrF/
ndhWeowiJ3sXD8IIYaB1OZhbSFIxtjN4iUGAR8ZeBq5LsgVnp72aOsbm08LgCHOhN0mbX1Z115aT
OOv5l1oK0vCecdcKfIqJ6xpvg1HC0Jq7ZPzHY5YpyuoTmQRE42IH2vMsg88zvHnZ1FGj/6aPIHPw
I16I9TSZ7HypWrMXVIj53pirRDid6V11/VzGQ6KeWe49AaxihIs6PvQ7ZuhazPHcZSCXgg3duHSJ
eY9o4yH4TVA6suz8Ojq8LiDcP9tzCU6LYlOOPMIha7VJ4VO42Ge9pUyUh6ovDr/IFkDloYElIp0k
ynWjYMYLQXJQa80N/gKfrOBj42Kc/d596+I7stb/UikwKRfkeqsriFSnvP0aTySE5CLaF5J91nec
mO4p/j2pHpTmPRV8UBfJa3cYvM6WhO7LZOx1LtBEis+jbu3Cz8RhO3L0WijnEPFbSPEGiWiqIBHQ
n5MIVvTguQJycTn+f0qngJizDDNw/0sAzunSY+eTLgPcTLhhOWZ5/KzmJEU7BLJinPrt5rijHVEn
eIrK6EQfcjGMZtqKJRvv7lT9bCVePzYW5Vu+q7X7+WlQKGnGT+r7AKX0+HdbazCpAsrTjOHBS7eX
/ZYjpow7Z8xktuirvY7kT/p6pzSHeeWtBy0grGYQ7c5erIHrbXoz3WQUKXKG9JFKx5wXKAEQ64TC
EBr9z3g2ZfqjEOTi83mWUi8SQssAUUrobeJcvxyjBIA3vDZRJvU3CVB9CxXbbS4r4CLDR94sSAYQ
ArE+Y4Ml9WXCuNOs7KM1kSMTPxnjS7dfaVyWlz62+IUhrxBS9uiOMu5Lpx73NHfy1/cbti5T0gd9
wHzTWEhNcJIplMl7/gSQlPKVF/RmiFu5vAax+FyjWOVZItDU0/75dxEA7RsUwb4G3/5tUrb5jeQz
T1laIgNdXGt+Fs9ZtR1+2Baxt2mi0A37dgIS1d7MEAugR44mgJgYGxk4n49muBz4rKvgWG0IXzZ/
6TsQoKOsb+cixHr9v7qsecuSaVo8fl8lovzRv+G/YdmGjqmLNRivToRHoyzECxV+cdNs7A0fxjDy
CyHuPSK3P8W2osRZtP9UPfbFuWCMBsb+eJ1XLBc2V8slNjIwDERABeykrSCpyh6ZHAPLKFvhRL1q
x+uJ2trjt7tNJ1MBhB+pyX9WZ8ju5mGrfdLvWpA7vMe0UIzoLCWw9krGVsxN0/gZ8UPOPDDUng5Y
rUVkjpnrBdIRazpuYzi2OXzZAa9pNbXUxJ9KJWGq7//sbo+7SzNlO2iSIr8+v2Fspoypdnst3D0b
xIIi4dlf+HzcRD3aZsJiSWRbgN6QlQ2Iy9A4vCB0EUrteEjfvzrpnuVWgILNgnp5sT+oiiav2cKK
I5tb9/c6dnsbaWyGzvVZMqLsSYfKvApIMqFQHiKFNwzSNtOVDmaQ2P2GiUYlnPcw207kaoR9HLQR
jRx7tEe1SuRbrMdnzCp+6nzZBX1M+oLpedKGW7Hl+588y5czCHLwwX41gm8VpAJeb0xS4y6e225u
tj10/E0zRJsC6+HK7GNrM4eJxf7O/uGy5CAk04tzNDpZueYTkZ/yUKMIr/s4s+w0WWcwakp02Gng
ytPInhPVBAb9kfH0Z7lVwSzHY4KSXxYvderFvhQzUzmFUmb9lB69L+zzldXBElYDUlbM8kil97U2
rJBNc7OSqU0/OnO2OcdGWZvRD/rk78nP40/oht17QM0W9i4DsALTBa1SLadQqGqEVqCw4Mhge0l+
JxB4Y1Il7u2p+nbF3hTh9k6yjzQFqUfadwEGVApN/5RJur0r2/p0kBrF+Bg6z7Os6+UiVhMCiAO/
6VRd3YlSdexrrMYfz7DvTQk3ReOrYQkapSqFIYHN7ZNaAnz4oWlLmCzrTuur90dLnBgr0gn/zQL1
uiIW0GRT6V9pdZIaJ/gx82i2Q4OOXF27I+xgzJOQAjM7uecqXHR5gZQjyPj9Q3GRHmEP/RrNE7OZ
hQi2umMCBj0DYWoxsSlTDnnNqSkBwCJK/JGTDTCIc7bqr23tSdBHN82J5lxThRECDCLA9VW3pyL1
z/icwDd2p7IxEDOlPDsixtRiCmx4dCYdk1NwiWY4QU0gQyOqyOSMA/Jw98ytZEOSRn+Wr06aPgpt
XgA9E59/3qYIsiOSGtqAcNu20kcT7U0CCxy36eLpfZvUtQv7gYkzJBJUINsNSboVRASL4b5vf1Fx
d8w+Vvo7i6X6lx3QxB3gVyRSb2zLllP/yMeHNaNqc0BGgQUWNwvo4dOB828QafEYMNhkW9+oCh4V
UJpK4nY28WWOidtUA6ScBDVISpn4I0v8AP8q/VVc90IJOG89AJy5r4qvm6PWWtCnwcTExYPB0pUG
hP9q9s25NwSnX179WvNKyMPlDzKu0ifzjWVYJbp+gtDTa+ysNO80xcbWoXtUcBxWZM8GwqjzmoZj
ZDtUZNemMWaq9cShkcdRryA/pk61gwINeaOegOUejYDv/fYeBN2uhNvEPeh9YOo8vDpR1akAaye4
jTctfzKSZGHuy9Kfx07O8E5Vcbc+ZAsghV6js98Gvkx0zjG1Gzxh3+y8TGXqa8VtSKfNGRcW85rR
gNlG8sSiL4RmIYoewFLUy2OlrUv+X+h3SWiA23a299PxufRcn+wiAkMVYOKZSv09k8TMuZfhAm4A
20Al4zuld2zhMgd/B9L//WsPSWkFqhxZgi7+YPfE4mWX9v8z7yQ9ZLXAcdy7J7Cf10AH0jjRwewJ
gbpJ7tt6Xyo/U6cmS9R2uczazk+O2DW42c701FBuf6ycM3ZOgmG6KWsyx4gkCw1jv1Gi0m9tRH8y
R4NzCHmxkX35kLdOLmpkADGkph5xUVxg0lYgdYPSQEQnrRmsQ6YsDSnVJFeU1l6krUuLY5ELSCD1
cCRhxiilsTsstYu1Nq4FDZxjPGd+h3FfByIlNWZwOMOM9sUe+izE080qFQxXz+rN+jOOXFUCPZQl
Y3B7+5zo0vOCskXE4oYanMWUFa43k1AdxCFrVco/ppoGAGofAhbzK7/BKOHBOqpxfPBp3Lgwwhku
9n8mxOPoBHJmBaruOAsf7x9fXLlBE3UInbumznw4F75mD05paStrue6sOK2lJChK/xDVOP+AmBi1
rDeNxBCSfM/rSZRVL71vkpXVWr0a0DvCcHPR0j/o1CraM6yobR9FIp88rNE2L9vYvPwCZvBUKZXA
yim9MQa9yOsUVjAIlZfiHMc+EdJftSp9NLZ4WnaZjmF+SX03LiwKp7mHTFgIh/pP17hkdhYqQ2se
D3XwTRf/zXSKjt71TxXJouYO1wUhKUdHYAhVLBV36ueg2c1xFY0LRJCr7UVKnCOAcwNPyogGOQJq
TqJHt15mqdcEun/ImZaXgw7mnK/VZN8veo2LGooUVnCS2EkaRJRln3l39RmvEuR1fM+l3AaUSkDZ
W4QG9/8RC4W4SXYOf5hrJyUVFUgtl5QtIVaEuCKQJFIKCmTRq5QGZqBJ4o9jjNV0PGcwK3JzHB3H
NEKlH9xn2MiuySAbQrjJYXYoyJ5a1H8b8d9aciSiHHx89IOBMAYrK0Gm64I2W28jBU+LCZX1JnSK
0oQvfDVIYfzzapR6W804DHLV2Lu4r3XWJQFmiGCXgMImiYeU+NwiU/4mgbwycyoKR3nL02cFZNJr
JX9XdWWfzkJFisYAJH4ZAu02Wq6Z2VIbAOrhXKljp1P346/dKpS+W9Fu0x9TOcEtoHsjhGFXOSla
fmTbZLp5qcsPpkmGNoTyii78I81AdnU1go5Ts8okAnVc4By6It3RARR93+uPDlDjMkCQLZmW3PcG
6HChzKXPZG4h8J0LEwlVumBc2g5A+F7VpdbrcsmiuTo2hF0gS/Ae3N/j9MeGYmzj29jl3rGI0QOK
09f6oQIg8xVIUlRx+sLBkksq+W2iKwW77FNASB0fnyNXZTTmIdZYP8RxaYkB66VT2Zx3n4OiyWhI
q76T+iMAc9yJpR0/vJkzGXe4wx2Tcr+l47SKX7A20QEIGu0SwMtIb7rYApKQWI68obpcqte9ea6b
kZslP7RupTqhaVRdmHt9jOwT6V1e9GpmFur1AUpwW2noQ102GfB42dh/3A8ZxwyFS7SoqP+z/JmC
xUBXzN7ls0JEUqTOKqD+cgah5O0VP87IVNQ266QuPnvC6jMF6BMnLI8Fa8X1K7lbpJLuG9cN/8FV
i3idch9q6Wu0clb2aYTkv1SicMReUvUUJYedhGG9uiA7qSgcKhe9wQK2Kq87RQ/x+TCItXbsPHZo
V54RXLKy2d5RXIDEj3cALQTkwhjlvVc/2g+S0ziVfIHcA7e7YHgJcExNvdnBcQf7c790OHOrNA3i
ktNz8TMNATl3uyz5ws4jc3jUzOju6h7FG5xm/U4aeIcp3ZLwHv2usUxNQRT9ZkT4p1FJlqsP05Bt
h3fCvs5mgDTL10AGDqlZCS36AufK5OUyvr8RULaxK4rtCNUjpOrprh40/xmKoZ5RzWU/4vIv9gtD
irUOxmAgz5/kdb2Onzzh3pXaXDhv5Zbna29evoe/pRTcpky8IVPn5MB2UvZOJfTNLZrXkhC++P8s
LzchSk3rCeQnQ3FYnR8Fj8JkvA/1git12cYzd6x9MTEXN+QB2g0fiRuYhENeuYf1rqrhNSbZq38b
pORzLIS0F7m15oMka8qmc93A4jvZEkGTkZ5G3HYwzkWDTADXXYixz4g0K16etsmGGnbLF775//VA
pOKwdgyjf93Id4aUTL1jVVwYPBqtVR7TCx6cYrDKuzj3/IqrJ4oj+ESs9NwRG+TpFNjmkGmt2Z+g
3ZI9H+nFUaq2Gu8sygi4mXNGF229/ifEbnXjuQOKyjPXdnlyNbRhflt80hXP/ORDgk+ciatJctMq
tV78CitGKOufu9ural+HhL9pRaD45hyXUr2CPMUMOgR8ck+Obfqz43kdZv2pfGA7D+1q7G8GY4E2
XCzgJ/t5i4rAeBiYjgcbRnjMg/H3jgefhmNVGJhFRduXYddTfplCJj8E0U0CIGQ6HJW3JeIaIP3T
N6Zq8LVAUzLiMZ3pNvF754YggW2IA2iEj7tH39D9EBBHTEAISndRaa3hnV5qIwA5ckqxyUR5am3t
oKNKUObPm68Ca366uuV4PmMlyuLYG+iYB7tsrp+e/CDJJGuLXuR2AlOviatFRiOIKgwiYpdjoU9R
kNKVVJi+Tcu6LTpMM3sENywrbS+NsJxuq0gIs+zWvwuLOm6XPxeHeQuEOhCLlrY98lXu8MIlRmVC
reJ5IzEuMmksKLHHwFJhuVq/dMhGDCp/XanS8ayxnWTYzuMbwlBLUz30KMsCzMXhTLDAyWEIgV1C
6MqU10GXDKPZaKxixOgWt5zHOo3llD8LGsjUnHT7RL/yl9UN7cB+JrKdqAgaOV8HVN6/jXufTUh1
u3+92q5Rtg5xubci+zt+k8DT/QjkPkyfxpGtcOOVORrGpaXgVl8Uj5J8eL5M/T6s0jasx19QU8P/
sRI+hz/grxkKo0+gDwODFbHvOeuF/xAqw4KD4QF0lF6NEWg7CHq+vRPt+CpGNIaFxIybiDwx7DAT
AiSScrUUZ4y8oQlrF59dZWvSbTBhgmyWVVVu01GuKv2gdKFE+TZ9yrjBT0TZVzX9mUqQGKOs353B
aYe10eplj4waWPWowvpZi1djPHaW+TKOOp3c/H08jEI6RSQVoAuayzkJ/J/qtkbooJB4wMMcSz2g
9FhM3VGYFUiY854GwLtFGQoqNg3R+kZGCC2rflSZ8y713ODLkgZrkjoe3C9JJGh/ssiVGc5fiUzJ
drnuP7pf6CnYE8n+/fMyxzx4aBxfUV7x1PnWn/aDc+vKgn8xiuLIDCweix1TWqG7KOhM6YhQc0fY
A3Rcy/I2n7KhKrn2he69BDWibYInR2DNSrKYdcYbymOwFcVHLpbdPla2edGpcQ3hnKe7XsKRw1Bw
HuCAh7BR3V7RK2ZdzoQ06/cQhL5UmzfsiNERJJblcThACTriXX/1xXPQPz0IWcrhXw6mha7P8Pgi
nJHaJkFN/1iYaTmkKeuImFgnrivEDqL+ivwWSOQiRqBMYMdC1tZPe9sABNQbaV8y1QBKoejBVsiY
GI12BHcOYhWy0LGk/9QKqviAvCcUzxKaNFSuZ1j0kVFHA4+kveYUbKs6D67cObggElOOE8MU2nh8
DMqghm4sEYXM/Fh7FsFPqxTcDy43sAYb7DjCgt3u7F7D3WYmEvo+y7eFk223uMTFtwv1Ik+Yidz/
EcO3nCfuM8LlRev7jQGhLoHtV7fnBsJb3RKemZ7JBbhNBnCNZGWyznx9/c0pHrku5yeF9VmXDAwV
t4f5pW7OUZKjqGqdpY8dcofLiHWS/SMjmvuvIZw2ngGELJRZRuD1VLRPgQb9e4+HcZVrJXAYl9uU
hXHYTmJrStOOq2MCr1fpdzA0a5U+qZi5+g+HjPi8iqwAyVD1XhO+X+3m+t6Jf63Y6gm+/M/bvuw0
w8E1S8BMRxkUnpcwK0qtWsEc6/1lJD0FuayLB0XH87gawFHQdqBFU62fUh8oPfI8B4hpFNOvK7M/
t2zXz37UouBnRQ0lD3MBYcVEd1YLBhQpr/KB2O6QTlVLifX8zcT1aRNyOwKhaZ2WbmchD+Mbjptm
OgV5PgwHXhnYJY3uxOJ3CAud6PoW6OVl9Vau5VjNbKFmgUDp+MuCPJiVsgFeftqxN9Xaocf99UHc
1ak6StGioWwBZHL0AOU/VAmJbyCR6BAKD4FealDJchIQT49H3sTe6pz+FLrnPF66KGuiKbsbJA/f
6l3hrnWpGFFAbycnDjQ7eBSDgDwcl4UpoFPt8xhlmEMWKFVUCwMtbOzTtrIy5wpFI4G1yo1aWATP
AbVUUL1Q6QBslVAqP0miJYb5ZC9xEnu5CpXHSmFGOrtwlZSNIOQjeb5mtEreJ6lZeO3fLgCja6GA
1DUcf2u1y6vIpQ3yosCEwJXdhQ4IiPida4btRLxpGPRBGyP60wzUfEWXz3wEH7qDfqz4D9fIrcTk
8T5vM/pi4cF/T0APlqcGS0We7LiiqIFQaqXWxCsAY/JjhW/rJzOic08TnWvoUejDuFCuQr91jhvl
o5DAt7Ju5pMtA3HHdIsLeXdJCx2B1VJaao/HR7fjXzij9Pi42rsez4fSswGGmiGPrtpgJKq0tJ5a
B8LcFOjCgK9tkp36EqcrwcMXgEX3JbIOVTqmz3uvMoS9YsJWBSfBN5q2ReDv98JUrAZFZ0zKBpoq
3yTwjmVSVAbKrKYuOgn2qIxrrWsuKPrZ1l6lHxKyFwg6YhZdlBMZki7c3nVhxSIPm2SJ0FE8mLjr
Fgd13guOYYbCy1SY1aQMaN+SxLoFFvN2yPnC9y5TsfzXl6x1OBMaALW5b2IsCFmLmRyXRQCy3GQM
aZwk/atDk5mMK43t9w5YLliJoX/zJCxvDl++7ZLSDfaKybg97vV4NAZg68AChaHCDdl5Y28kv4He
RpXaDT0WE3sLUdBFUwpZeAv64nZKSM1WU9qQ1Uo097zlUxK1kfM7vLNTIiyCB/1Hhab0M7L7a4Vf
QQif2u05YvTatjFuKo1miibgA2pIcqKdpM3pe+anhsCTzNpQRNCkIywJ78RcrXTz2jBnJ4cj17ep
ygKkXL1UKG8be1MQioTsDhZsRjK+cI3Xb7Nf/nA4h6k8tUUEQOqSaLsI1of4Qmy+zYJ/cfc69iyp
8vguV1sFwr7+Zg3Lz3IwRHwdLBkGvIxKjRHtzAj4rQFxZGB3cgBG+r7JMFZulTVYmvaxmOEQo52Y
ceaZ3bs06/6EuUWDfdfO98oiM/IlUaxZc9lUYEQFaQtE20k/NEtHytgTmCHRcr3bGRNaoEaW9U9w
nl+Ngm1+aYWzS9cR42aEGygylfg9IPV6+UGjP4rmB0vWDU09FZnoOWVR5F30McgABReUi7tGo7p/
D0WTVEcKJ3eUrSt6qi1s2f7bccCbfua3NAiWvhBlcphnaCKlD/zRjvU9JySFnz1PrMvsyvQ+kIN3
wXKQ1FDafv70HLsUqc8gWxE3c/YE2wzSi4R17GUm4ATOXmSvub4akxopsrmsH+f1inxiuC2ySGxI
uNGplVR2VH4zuRLIk5CBl3Gu1kdljXvmcddXfwNEl7r/PRZl/DksPhsYmAlzcTxU4hcp3BMSqe0c
wEqS5RUdIEG/vSppogV0HUxO4ca/w9E0tgketbu+on5wLzo+kRKIboYNG9j2inLra/KjCYnz2Nz3
/u8WI3+0EpNWzHI+OqmWYrvUNZ5Pp0OmIas+m8PCSAanwSgO24n1XWAv9d3XCvPvY9Wd6LQfvOnq
vNid/i4qG0LsKly5VtYf6OOzDVZG30zuuis6iknM389L2qThXtnv0mDk/6QdbXmWY2PUv0nkoptk
hJYMT5n1CHAI8EZ1CR3YaaTtwb83NuIy4MYfSURlpZl2//bAKMenQpco3DSnkT18VX7HnKZZo6dk
OpmP7MgMTyzH1w6FF97q5jwKIUJJhPHYdgGhYyaJaFi5q8jDYSGUPhXdjDydb/KZ+MJQhV5eLv6b
eEjMtnVxJcSNVEJtK2z2HiKufyQM1aLg+7ZygUiXJGRny/ROemVvu1riAsZ0pZfIH1cbtBrP/5qm
z5/EkLYkJZhbGnwwb2TZxB5/KxXIiNBXrL8qKdVSYUrNxwZRpiwAKXVAg4YwVEr83MwAwXnyPHTm
Qw1+2EwLU3wRO7dJm3Xwr6J6bmWWUY89pX10dVtRS2KpZxfIDIr4VCm4ukvDgThYJeiHEU77/91r
wRjSGj0CWYqkxIeD2nCg1Tsyp7aJOXtaANXdVhdXEE0Ir76khY8KEJ1iM0NPYyRYL/cfmDzlPxK1
ZO5TdTCvPrlB/wVn9Rof8BMRAipd8nCiJ4NsWelfWpMknF3s162yWt5pogNqY1Z1BdsAwIvhz5e0
hxS8C50rxmeAXvZKWg6wG35TMVC1VCSahpaRnDq8rm8N63NgjoKNixABFveg/6nJTAXQ4dyjRQ8h
NMZduLbWUnItr6NSURRkaGJS41OtmgN0hgGHePL0jS6Bf79W/wy/TcVrdWZm6lApCDTMH6jwVBBV
rao3QTDhqzBVI0Zdz9Gxt4usUUm020R7rO87bDhbOj6smk3D6NSDGQw+0/BX4DQeVN6vDG38TEbO
ryUnoKDjINMNYGLidIHCRNojx414hwEixZY2L9UnqfBcp/f/5vWrVgMnmyXFFJzpizIvlsUkbLva
+eAlPBMkUHn8VfzhSsdtUnt2wBkCdWcNlt99FIgjTK6ink9TkHrbSFSbAW3KiUSwLZ2ZqftnwRe7
3PDE889CDVVhiGWKJ3LMPlQZXKC9HQGnzokBcywMp7gHgSCe0LE7xo3sBUaxU7enG4ouv2Cp4I0s
uQyR6AEqPA9RC045sxRnqPXEoh5sOx7Gxtxdje9bGdK57WuQZ7ElcyCgQRKiyjqZc74DHqyGdNlF
M5x5+J2N+32eTupm25yBwNKRjGvVUp5u4lnkYyYoboUWxmc1Vkuo/eJFeWs50iRSuAlVYWkgWmQL
+0B7M8CojU5ULirDW+Xd5Y9KyXdftsbr5N784wocDlq9VIoerkc7w6x2iO0Id8kIqTeiWqUXWRfl
WLPYWUTwNjpfyhSglq01B4rNaGvT4AHhEHWhW25CR2RJz+awGKvPVfxV4a+tgBWPKJATl8Kk9ogx
pq4uD67HB2LCFpUWxDgRF0YYVz2pdhYIfDfbYss/dUCMoFRFvvZ9sQtfl3eIgNHPZBqSILLYdtIq
uxE37Bjz1SAS+Mc1dDiD1cvoXhH6qXRo0xbpz5s6WWEx2Xpg/MkiJp4EuGfkQiwy0akQ8392FN6N
j8wwagfCxKghZIJ0gqwGHDLS9zH+zJw1KN81QM5PvYyC3zvlkbo05qyn/wulyOk/X/Z9Tzny5r1K
Cn5Irt0Si9cmy+UKwhvOiI8oz4RHJi2N36LlEq9uwz+93F2EQazCggyLhZKlroxiSp6mJtiprQUm
xiiW6WQrLbw5Be+tFkWHt1SSmFrXveGucwL5VUmjPcE3aH7iZe4gJrN7xwKFuWOIa+Mjb4QZRbe7
x1wE8F7sdLURDfanTnl2HzkOM6IG8oF0fUzfJ6ldtYh/5LH9N9fkhoOni4T9kmYcEiwSKaYetvV5
TPq7UI1y3LFFhEu0cV9G99cORfMv3q5+rVrQfoY9E6yJEY+DnkCagxCvL6ezrdW/EFbpPoCply1Y
3rK5vMGgq6JQ84cFsSkyfVuJxWKgmdAd6ddKmeIa08L+/Vs5t+Df/kpxtMyenv3XLhuNvzxT4rh7
njSeKqO73anttCukCTiVd2whH16DFg33RWHlH5zyQi1JDLI6bGu8y71RrdLVplIbqems+g5YsD2k
83ErVKEGg21tNOw6zbA3q5az4g2OgZxE1n5+8RucnYldeDm/cgkf8AJvFCt/lOfZpIxkK2IRgVDh
LMQiZGup4QQ6gxonD6GaLKb0GRQVjPg6dGwZ92RuL8RhdHlPuRZurY35AQRbOtW2kKyTsGa1VNqu
TyDsNmUpRikx4NlfyV4PB2Hd0qGEnyZJYKDFcl+WtyO+DI9BeLCfVVOWS2oTOuyViXhMgjD7gGyk
NczSxyDIwlTXSQFpzmRQbmsfwJQ8wxGzspQBgXAqpqRGbwxWXfJw+o4XPD8XaPZ8GOm8ttz9KJJ5
3qz2embNSyglHAvujlS9EsysshIEFfVG3m6+5GmfScFdg8BUWJCtBoGJszLWKqJ3XvbkU6di/cf1
YuJ9iQlzs4S2Q+XXzJUppvlOJpBRKKHbDQPdH7wcTWzuPnqIDZC57kTPbJq8/twEarWynCL2XmFR
s5jNeFH0rVX3EDaFN/Bcdg0MurcCBoLSDdR82HP9I+bvC3KXT53M+cGvXJkMn3azfnN8Kq5H2/t6
rvqELG9xYjyzaH+rYJRLYdMSan3ADmoHr/Ejt64NyfS5w2fzQF5I2+IFSuFUtrEydHNFsNoiXt1I
IQjbNmE5wPhIB3CsClH9paDNj6B0BrXpVyPZS9O/9FWUFEvE6N1ZiPU17Cs1WHLf/3NGhogRyuck
lTE5RTinA68Rxtb8JIs+THNcrwDa8Yyx6H1End8natknI6spaI2W1nUgEskUMfG3Tz7UrtkGW7Pw
6Dxkg2RnN2cHq7mvG46uccLQbvu7Vc1JEaT5+hS5dbSuuq8viBL3Bz+9wkYEQfMg3c4oHvjqb6Dh
u0/bYCzwx4EefB9uuEARrn1qYcieBUIA4qlYnpxqAf3s4LOrhIsAEv5egUORXwLH60MhSFfAhzYj
Xcpa14Z7qopvtcBn+tAasewvX4LJVu1t91cHqkTIQ1sVMTuCDmnhEdD62hcybH+hVYqB8Vl/kBm7
PEeZ7Sgczw4nR0iRc+xd8onIAEId77B9qqqRA4WsiFNkxbYuzDV7VGOExcpSSqFQ/3W4BLSJEUWS
bQYiY4tWZtWJ3MujxLoBhDg+I1HkWWOul5eeC95TRhMlv5OLhIHfOKUtI2Q045aXSUlOAZmt2mEI
G11pAwraUBmiAgg//pHSQmz0NMCwaElfktjgte3JRPkVDijoRd9G21xb9hXJPHpBFcqr6cNEYjDw
3cnF9UvSC0Mf2ojzCM4hRrzW204LqxjiV8r8JdUpB1TL3th1JoXGltmPGjM/NOjYV0iobsa9r38Z
qZsIrV1In7g8+p625BpCArSdkoJAgPbKqsVlGsxTySjdBTUZgUMym3PZladF7UjgGqAqE/UT5pfM
NAZel4VjHo2GX1lJJPZwdo9Q9tOOG2GH+VtmUiCU5ac8AM9KpOxkLaW2LM3TT1vOsVMTbVO0fcG+
wYX75WHtkLkiqdSpKJ+eU/kh8OAOCPF8YzpTMyGoJqocbUmL+SSD/nVoIfsfq3md7ILvu/uUxR+z
LbXNCodSS6479tNgS3g37pchLD5JZ50PWgyHHX5u1uDU0PeXNXgnkz33mYg4IILJ+51ABbv0cC1+
xh8C0CxLmtX3p+hZHdIWVcp4q272YZTAGtE+SmRzAa/S1tIPv5+E4+Bei5mdG44lJLN5fGrBbire
8G/D55HmOptG8H+lIlXiajVu+CSkgClOZHPfaMxPBUB6Hc7b7DMiyU0qjBgCK5P+EtM+bWlgl3ZE
YN4kCxkWGe//rKEM5KApyKdgHJ35L7HDTJQuCASOz0kgsJHBbobtVBNDXMkaV+wr7PNBoY4fbNCH
YS4qyB1WCSEaQ8FUtJZqz+koL/d9k2ZCrKkIuxK1t7NMOgDW2huJgBPMppZk3oMbFnh4eli2k0Xs
fL8jmWhoIpkHj+hCUQLWg28vymK9aBLDY7+JsGhdcKRv5PtXhg1y4sep0crYvoQwAwOiEuWq9m57
Yi6km6dT1H2RMJSljn/8p9tiE/8kgl2h1jRDmoG8abNaZ8lQHXQ02ANSprFSCXNa8d3yyP3ujMZR
C4S90uqf5yeqsgMUdf9z4hjkSdsBtSdP4GVTvX2vsRYE4Lp5volZe8mn4EMt+uEjF602ch/lumDi
coyuLee1vc3yKaB+9sOeL3HV6oVoawKVT/8HLyPcmCXEfp9G7UaTU4AfJHWCGiEhJkkkUEF0d4rB
6sEW11966Y3XI3tS3on1aWoO8mfh6O8W37kT9U3DX2EAEWVlscQsIyetyi/h60WyRtiLMML4oXR8
wP3VrxnoTUWg6k5LM+IgCZfobt5GF+KrvMGv9zg6D63f8QdTlqFwxhhHE6E5ojc7VDzt9dfY2qoD
zvBWUmYFssUvx2yUv/ZP9GSBZ05x55uT15e/S/+AI2QjK+uruh/cPhJzdEESPxdOketwNVrbaIcg
+TuGvYDzosuv9CDplo+IjELenrHOYCaWTkzvQaX+Smn1saxxUIBStdgrysD3C8BhVN5y1JQcqXou
7pXGpVYawQz/N0WNyF2wf4r2hLZr5hvbvzRZEAz8GB9K+rdeU+eDK8ZsFH6OWa2mrSmaey08dqTy
TdUT0iGuHuG8c1+UprYdaQGG0lpjjnzKarWS/bEjE7pRl3U3kr2gg2Gohb37KZP9kbjL2+6oHjDo
M9ToZop4YuXkDQ+DCuRLiFN0xxGc7/sYXa1PSkTnfnIY0g/N98tG/0uYOWXrELPPktQc5011VeG1
9UkwPBZeOWc9ibw3OablWuJxZdAvYPIpW37V3Gy6s6H1lVGte3Gtqu9fZATVAlPb56oDZ7wkqu3x
TindZPLJ3MEs3G7GxKF/Ehg7KAr8jE1AIwVM9fP5bd/DtIos9adgyVrdtop+w+hwzLtPOa3XwSUq
0rWjN5Ca6iuYRo6T8GPl7YwnvkAncuw59UeEoIjuiHBf3eAf15jm2dZvev1XdCgaySG1drqVVAfR
deEZPmvwcUQ8moNRfQ7fp5gbvWI4AxAdE1f+J9ym/NAHpfsI+2Q5wNfYyY86OTvGW0SWMmhqK9af
nrl54T0OwIsfqqneKRvkT1j7OiOK0C3zLdgi9oAZceqEzKA8Rda51GT84FTkgk38v6f+uQw9gCDh
uRtgOyOGW8AWmxiJmMGQ4ShC+5MlheDbKxa+QR2wJ5DZ9ftUaV0QVAW3kEoBHIGo+rOWy70nMWtA
WW4pDiIQMFCSFv6T+yU3U7y31uoWdQM+aGPw55BTqD6+sdFJBx7QGJhrjrmrWnxPImjkEQp8WqJP
3qrBx8GJDHnZQjClje/g3yuTvkjKkaYtS4YuH1LGFxp6ODYpQUOHBiP6bmqlALl1kku8EDg9DRe+
1ToSR1qPU1Gt40aMr242/4Dg+/QU/Xt1KA32mq9lHDVY9f/ioFccbnYC5/KxHfoj0T+WhChc9IqV
Y88h8nzRZDz8rfnnxrdMr/OpMBXSQctyfYONuQN4/F6QwcOSg/+P1PjVBSsS8IkN6HT4STGdLkkl
79fQbzGZui+OqKyZ8pLloTywPUVRts/M1fuXuFyxM3kdeEJP8k/2sAzabqoSlSmjU2CLhrlhtA9m
OeafEypGN05h5QyOe2/hvASxDWQmn+i0sq4YRfDPdoNsUpelqEWHOGrJlJSyCgPsjEWqvCxk9q5N
gl5qprGKTdnw5pRUtfSfgg7Zp5FRQUYdhmTlacF1CzSU/vVTIo0EzDm0n3mDe2riCcaoEqLXQh0k
eLx1e0N210ZWml5h00NStz31z1d56otIIPl0l+gOjVWdRaFDfePK6eojZ8a5/d0s02Q+J65QEQcG
2eEMCzhNgT6tw9KeUrecJ/zl77kWjDPJN43fYosMfHpqqbFhi6rCnNiBwLTvRSLa/7oqtfFZJYFo
MMzWjIyodWHCufnjg78h8cX4Wk2ce39/dmuQ9+ugrsB4HZvdwljPWa5CCywls9H2E19SaboMwBam
mP6IGQuDsvb9f1rbWiyTuD7YmBNb3OPW/cdozTTfGoUMfyA8A9iNseH621L9mFdq1LbBDmd6YxHl
klb/mLadgOHyAd3OoT9VdNCNmvXTUoaVHzO9Bd3y16OUA+Qxz/4ZfMqhciPoMXDVZJjtph1H8GoE
hWNEhjUx8rl62s+dSGjV6SgtOEzaZfyVSHxsX0Y8MQrbJN+8PhWa9wBbzvkAWpxfuZXEtA761seL
KFIjhCVJO1dHoDecyLGKhw7YWObRHZKYoc8027o34b3/7THtGj1GSp2pi9W4njMQ3kcKAF8r6R/l
eR/0rxs0hQmsc5gK+JPB3v8O3RKUH3euDaKJ8imYDGvDWIP1WRpnnqjBiVccqkBKMyTqDf6UmGkE
tmjuXZCblsmlQZo+zYwQ90qFvmzxOJi8rL1TDj+d1LATJ/I20B9gzmq8yfipkx+UscVsjc3xY+Vx
8PmeCMTcXIcSVm+jIdVvxgE3IWkd10S4pgkz2G4slKXlN+4oyBQIGEUqZ+gpwJ5fWLLN6jYBdm3E
lPV4xJWOq8SaiKcMsgjy2Lb7s5m3nNQ1a51i86AoEKT/fXUU4t6nBDK21UWLu7mfV1A55XVWWOrd
vYOsj900TxZHdwLnlq0zxw+iEtxhOXOlh3UtI6YZEn6JFj/X7qNJYm7wsD00x9mzx0+f0Mj2nPVk
Q9Ma10FjmQG1o6KPBMwVNyKxr918AbDPZzB6oxrDXkTq8d598te2M6NVd7tU5AD5pwgeWmA6wg4j
Y25/PIJppSzm7y+FJDZpDztqfHbNVHi7qxnC2edlKOyieYlUQFroh1GGMb8TquwTxczGchzBwuap
3JfvzbvLdTylRtgyAU+MqQBZvXqqfR00MFNIEL0GncUYIGiuso2p1FLipbdLTcPBqvBo8L/bg0j7
N0t47vXflvRpZ12ZJB2uxrdz1jvD9psTa0fKGdv+YOzj0ihafQty3TsnWFQJM+V+sco17yxTAgvo
6w5W0v+89h+n6JnlXvyx5ym9LBXblxXMhij+DucmSP04acVzhuxlLwKI2WcYKMf3+V/ND2HK1ngr
0WZUxAiKPTF2n3yy7inlL5MZVLSp/lzLtdCofGzU1et8yn0S+4upUg+I6VnVSIsVXkpTowPaQQ+F
1b1cf0lWPzGUPk1g7hUkWS2HvfKQEWzJhKvTtsLdaOqdYdA/U7lGHZFEtaEfI4Xb7sj+1HbVfOLm
Sdow6vfPoku6eGHoTucIa4eAS73uIvKFFVIGmy6wTOA06ZwsjwPcvqSrHSfYajCLoatPmu0HPWy6
Z5Gk+DE3j91YSyGAqWPyv7zkFjvlXtVEViLb7cV6OMdWj5hnMS6bSM23cCm98eJs0Fo8l6BiGi/6
jKz5CB2kwvtcuxGgd0nSETBt2sS7G5NAyi/tFNyyMgJrkmFyUyw5sn+NmSZZNZyRyj4wSkcHvbWC
xEVJ7QAFEU70tyFhu9FnS7ziHe4yDPtrDBJs3jWfn3e63AfQRhUR1dqkQRf1d6wNo2UnRE7HYPDJ
Rf4zI/A40rr2jDMIMWSJvk4FkkMr+BurIZghbUcFmdTbDFefTqrJHcNgUUGDHXIH4HGOtHFOh8Hi
G387PrH+wAhb1wkS+jugQYlkhM1sseibZM7O6pn0uck+YjzUDGr5G/UELWgxxlNd7EQtKsr8AISP
RccnhRKnXjtO+cYGiqiDcTPVrTtkxHwSZU5b5FCZkRYOXfqWdLccxIgYHOv1XnAE7xJ8gau1vKhc
EqxAZfDovFgT7jJwPJNtnJSlzfyDgOsUqLZJBf2XJgkP1czTKqog/n2RnvshWrX5neG6a00erKOf
nUYnosBy4yLBc+0XNEXTIY6fv1hUpefUJT4EXWOueARoHakrR7sdSzWp6+9nCmuFjhlsykyCDdH6
3lEqfM+CB7qjF5jUX4lxOrGybVbCItODfzHY9SHO+/Vb/+G4t0JuiFSdDq6+5SkWOz3X6iQdOoSg
Q/8Y/jt4ltZagQcOM1xCQALJyh8lyDggWJ+TYIh0hUjd5XPsgHe4kXhwJvSuRNO74zUapO9wHmwj
dgZn0patRYZNw33b10OABQgHDVZz4RArgERfN2YajCnAmZNfJq6oEDE2VWvfuGjcW0RAAk5TGBHt
VOClIdWHLXrmzlGCPdM+VllV1oYnCbtHoFvfuFez05wVlNmTHESyc628faHyGTfxiR4v7f5kgjzd
gnrp9LXRejYifzhHsmXjFMiN4bW0yAY0CvWDRJbv6EIFXNP05DRocIqeOgmFo6HLEc34WDzZUU5A
J7mWSWYlo5VUU5Uo0+E5FhTEA42QH8AV/9eUCU5RAz6585XdtFKF9KXNBvYgTt5fZZeNuw2AleZv
JJ8cDID7/AZEIQWydzb22l17ZzCVKUE6hVTUYFceN55c51X4mhR6Yiz3QWWSJwVMIwTO2fVTy7zV
IhT9p9L6/3N3YRv1kRodcRyGmCmciKpqxUuH3L1E26M7fRhc7G2oBfbba8K3xDrhTklQlphiQNIX
rTEdWqJ7lIXBQfdOeVDBuE+t8Vzs3heeSqrnghKb6f2tLEjY24ZU328BgVT89tBdcuIf97Yw11aj
6cM8T2XuHrhpe3bG+YVeJbIT2Ed2TmRprWc5xyJqtkLESNxfb1CJYQRrias34U2P+Y56WaSX/+rL
2Y4/3dKieeF76MKSTisy/0bOc/ipRY0WzEy6BAa0FhyBgfk7XNUgiqoXkGzXykGh1eqeyf4nlGNX
znbWBT2q0c3YjnGOgFHOx5nbPDMGRL/0ctMmfjLOYohLKSHhjvEz7hYEH7SAQuk/8Ze7rzzZxFu+
1PtPgNxZ9i6ekyZnH1vF05EYi5CyhFxFBFkTVcg2v9EoJt0PVQcQ3sHIORr8eRnXf4qsmAOVBDKF
jxK/VtARKvkdhBz0kM/G2uha4jZcXAL+zdSasdnKXcE3PuCZpl+bFmjUsSjWrxp15kN+YoQ2PCE5
TBgdMUW6Fvm8f/E416x2de1o7GsKolJfJc9u1fAp5uZQzmebh7NulZdqxk5WNsek4ARrnkcgQjCG
XfXy0No0bgJoNQmBYA7EBeQymTe+YoB22kJM43EFj9j1U+UDeg4Fpd00s6oTCrG3+lol5LGjUl3c
mRUs2g+m9PfC48qoR6UkhAPt7BN0EEJRAAJWIhohBu5cfBZMXy7kRnzgZG/oti9oL6mr8j6b9r2z
jxNjao1gwHFhaR8DdqHCe0PnlR3uSZx4X/j1ATPaAQ6fcmuRNAhVc69Hd9mm+Vk1q+7S4Z/dJCV5
0tw5eYFPzQAgRiN0QdFn9i9LzVv3hDkvZBcF7Rpw8a+NqSrqB3bw7dUIQc8MscaIYaVM/J/4T2Fs
nNuaX7yceMqYCzJf0CUSjDpZ+hhuGfisiRJo0fF3jwPH68Kboik7ai44qa1m0pvgdT8NJs6ehD90
xkNot+rZVorYBN3nSiiRt8gK0W73trGbc0VBm7Sk36M1hVMXnWPkhb8he+wFQmIDx0cYXhCamf5U
1wjRY7b6uf7RuBZzLuyJhaNbvor6GABzU12NaZ3TnHqMMApgxXWQc1rrh0wJygeMaO3btuQR5kM5
S5ygErhpEXqOd5iMVLHX+EKGASc3wrGVpNaYlZ85AXFQmgIHQBQ0G3PUagzqTezeIoDfiqNtWksG
Mjl7N6IHaShoXMiofgye7Gpu+2q4kPNWMYzVeNEV67uiq5X5krPqccACaN5RPdMi3BsCV+tUbML8
sTAZMMTDdMX8UTnGQ5jnZBM1yRMJCBXTXyQuW4q2X7BFj7m5i1IuBYduZpvNp7txGa9iLytEI6W7
4NoIdBacmVDsgeAQFWwa0YalRxrSn6IIx3thS54PnPjY85Emhunpf+IV3QgE6fcP7F5sXLc8Fskp
E8YUaQrhyD0DNrIRc6M4vDRVYnXPzC4c29ZPXqVrXY0xI+YPLgKShWD561Hn7a0ahT/cWwDbivf2
XdUgm5ah/7u7GWO7yq/MNML+fanEQHTOiHVo5TklBF47NRbJyO2+hxxirUGH2zX95nhbkeaihe1C
Pp4fR9oMuFgLdB0oad1LT3Kxim6ykCt4OR3BjIqHevuyLHrPBNHs3Nqz07SCB+rwlfChV656/Ktf
CqXT6BviUzyRZcaXeHP6NwltRdVdgEvyPgdgFJNxJsGXpnnL4+pw//lrxf5HHK8nuUbzvc2Dtw4w
ubQa2VeAEcA18GqcU3+F7k8Q5KGt9UDeoxlRDa424fyeu0jmloJU1fIk37vgmOgmbFoZEo3ix0VA
BE8Esbzt8YC7yh2jm8DS+pdNFMveNE27dfT5DGobdbwjvUu7FW2B5mtA9Mj/3Tq+KuqrA5blUcws
/EdSMY3T5XRD/mssYXMV1G7oqlZAkfRcgejBBdpg5tMkjNbvlTUr9NbVrYtI10GbvKfj9x97gKoN
R8VzAWMQDh/iVO2UWpJZICzbjYXpQPxpOXg1And/o4O1IOP7yqeFFUV2Cuh3ei8erB63l1o/e+vH
7yqXP4Ya1uBc/6ZS+IExjmNyxjefEUli+mn9EnRbisMU/zvf5yRXQeuLHJIZOxwT40n89cfHRRoR
M454F8GAFCO8+b1rVNdCzIMjZB1/2xcjAsB35eqBNbWGYxHy1GUiDUUY7yrxIgZPHQfbV2Uu1pr8
RrhE5ufAGYdUq3Yqi05uaYlzDwzvoXD92pHh+achbTP4y1N20U7Zmz3qwxbhuSJ6TSqw3EGawAcT
2oQblyJx33ZRt0iB/F2OpjmUmVCDHhCsa7Wqh7Zw1oX0zt/HWQ29YS64vUdKwBKq/5O2Q3U357t4
nQ6iwDAwLLSNORqYWEevS4ERz9vOheI7dX7hTvAtD/pIvt8vC9INX2vBuHl//MS6rBtYJkjCJXTx
Epo1N28kkcLjOcxlm52aeCqQGjeKK0wbQLmkogOEuVigAlkVSgoKIoAKkTgkw6lFAOqS/Sfmx6fv
9BOVjKCdaVsKclBcNCM9nql58a2CPnR6l0b4b6dF9y+MFD9amvFn36DbAiLqC9AcYO9tacSVL9a+
HuV0T+K1L02Nya7ugQnLsv/3jrDijBHZYf2UlZpVA1e+OblVkQasikxdWyJxqdoIxvH4YjeNRsnx
m2XEc0E+Xo0GEDsbS/WeFsYQK6dxpjGBunyuIWwfaljy4yWjERTGKUolyOyVMrugJV5OnItBKJNW
Vcd19cnQm8wgjvZer+CQvkO2spT/qaIi5aXaFhYPyDWm0S8eY+yM1gxT/jFsYgLRger8zZRRChjL
Q7xCeELWf8la60CCD9PusMqSBcpYvJHW1h8BRiWpaepNF39b82b2A8qeYToMjukwPPoZ0oDrysyf
5Ra5x+ZfsRm7Tn/8Wykm/k3b4s8JdE/9H5Tu+b4Ad/vvCkE2M8xh+pB7I3rlq/dpmIsFDHSCrbbC
ZKDzRogczFbG/z5QAzl3HQNS+JeQOQXERYyaADPYiYldn6vde9TshTCHs1L7WUgtZtRVvY/73h2x
lOggWCJ6O9bLseI2GRqGkpF8yQfINhxXkc6OtbhOq+8uMq9EgQ9pLHAIezGwIUQbmlubSccL7Of2
DgY8uunmJMAHbbOdcP7ifr4lrAy/vR9A5y7nPMpHPZ0XCLI4ashTaHr+7CdPr867nBHtQBBhci7b
DyqDIdu5kxbhr/2VkMCh25JcxZLjOr2E0D5XCdMZCWXqMDq81iFd+KmUhBqnPyjlYeH0N/RmWbdn
KvBF7A9hGNF2k7nm64+r7iG00RurUm/sFQvIHDsUMkeLGKdDlkH0p+DhcpweXxnHOvVQHKWwAnHb
gWm9gmRExM17vMeWkF8NcV+0qX1dQ+Wh8jPFOadajnY+9TsGq+u2T+HENYp8fadS89vyTeP1m9Dm
OuhzzhHfQ/RW17clBEid3sYGyporvAsRxaT/WCxiwaJ55CcloQp8JcFmCfGtaAYa/p4boAIMmkE1
haCAw2//Pb0iRYHBs142/hc4yhOzF93vAKn3Q3Uds8Pumj0yU1AUSVgooHapZlfigAS9PZCM6R1e
iPYU9Wp0DXtigtXXTOdgMkhf8zJGjfVaw0XzDLfNS2AVa1PTrJgUkGQj5xELZbYSe2Hz2ESKm69F
+6/QZY4KZTjAZTWv0N7uQZqicigvb/8ujfLJjkkjBVAgjlZDljJNgraNboqUzLLzi+y+AsguUxv4
fWsiJolop+fFwgOIeI5yL3p7CnH/VXlFpzfeXrZdjgIt3WywSV7MRHXCOPSahPH1wb/R5wP+rXdR
fDV/L8W2y9sc3N5KEDWKglZvdknexgrvCezDlDtJQLD+ddrlgczVbARXpXVXapBCEmpUaq+8iwyx
WmhtHJAJOqzYqfTPIsZQAEOOmt88pljxwgvTT17oEWVzvdDMMViGAs+oitlGVK2oLON34vV6K3vX
F63Xt+4Klfj22hTxet5SwoNFqdZDOvwEbg8zFPKDIe69uYw7YZWksFIrw3v9BQOYfxk6gFXHUJHz
+esuYOpeeeet/tjOyRjm4FEpyx5UAYGRO11TXk0bcE/ExPdZPNlSEk4ZGNHibj+YpZ+qXVEC6JHd
NEPXPM6n0SkjUc2L19UdNLOFaAlVG6YxYcB4ZtRGea66QtykiZohnoblrybTx8VbNDiFkiRW+pBL
TdcPS/nRxBtZy53dcglZ16xobs87qWeXV98oGVbXAss0CmoVcJNTYwXnK2ogYvltndw72DnNNZUP
nIHF5/RglnGlKjnJmHqLYd6IyoLiDNOTx+WpNj/TwmWxqjvmxeG6AFfOaD9pszyZLDwMj0h//LFx
FoBPF1wgTtAGWbGs/DjJQ7amX1EWHOVeLkIljzaBRyBm1q0m+5uFlL3GMTm0jI2rEr8+k4Cn9OLf
V1F5gi0XI1dfG+HoEctEiSO464EaXug1EB1u0YWrn2buXeVAAg1XUpwXikIMoag0tAsx+rA5094b
ww56rBa9O77bqSHjp0SHF8KnHsuV3+Hn0MfZdq46tatDjDitJTbkPgLdShi7OkK0hLjedulid7gB
1O5/eARTjSa6++8gRhbAD+HAcIl/C7jM95LrTYyJywY8uqSCqHyubYZf6niKsf8RKJ0QbI9ksrHW
XB+gcRa7uhDhBCBvpm449U9gLumE1DLOdx6btiREqmhqXzM8bwrwOahAZiWe50ZSKMW7B+eA2PZH
l8GuG5y8ZjPmh9ZVmx/qaZMnhQ1F6slxZFik/ODjKu1T6ywWFmFXA6Nwon4pUO+EfZ01VkXG/BVw
mbiYWGHZDUw0310fFVjQdmB5pkDFNa3mmgpwLR1rWMRj/JkfCtUaBM9hpyWc2jdf9FieGxCcSJMa
h8f18rxkN/pjMX/msIFFnSs0bSXf2PZ4xU/bbtajWG2q3gqWPdWk650kcRGXIbF7SK2jGchx5Jzq
Z/ZLvbP+VqYoCU+D3Dkhilid+plREyvJM6lCtBA8IOTx1siX3RDpkkczTJODURteIhRE7w6pyJiK
hD395RF+uRQ6mUEdb05qmyU6yI3Tep6wRwhhedgTG34LwZrNM67rGoUPsL4R/PNXKYwpQyq5iqRd
qTM2DbM1vlfv2X+ui8vtgOxXjtC/bxYtYUQmbo52vzeo2wyz5zzMGHied3l2PXWBoAMNzVPj61+s
OEvNtNygdfkbTqwbpUwI1mjpT1c4aMRQiGlEtbnk71v0+g0MB7NCYxo1OprbMMxLFR8aMbagePcV
0JaQPwZxJd7A9ArcnnYL74RSnfRbKviB0eRbD4kqebrMQg6j3ULnl7sJsKZXCPteG+dunYR/21tw
fFtbgO7Th57TpzwtRaX5c8BEPf+/xQynmlY0KZsKNcLfjPDbmp2Imzf+Ng3WcPCU7NV6zIkpboM2
cWG203b2lWNycIXV6w0Fl7exz8JY0y2GkfCcF7jBVqNmN5hF2t1ukBhLj8RyW7PKwoQzBY+lLehA
yCY/Sox2lwy/J9zJp0ncAOWq+UQsDDqrxp2R3C5l/1Y53sGvyRZy2JQ9DEjQq5JLDpmkG0NriF/X
MXmiApeSq3kFG4EGtWgs+UFI12qe6OGs+QUQ2Apo2XOIur/8DjsJDRH46dO3xqCH9j2QP9GfaAKk
q/GXrj3OYG5K40V//tnxH6vzecfdqXofVy1sdROACJTctPn9z2Q/Av6FkX/Q0kDwvP7Lgq3RIuV6
YlBNOnhYQb/gfJ+D2jheNmCe20yOfG6LFQfSHX7SbdYda76gAH6KpLTjT4evJyDdz0gI97eLNp3a
i+hOiU+utFdbiXtJo+N+D55LaXI7X/T40odbDrd88QBXQjdJrat2aJfabKNQkb7SwCa052+MivH5
FTalWnoFiCU2kDUHbcXA1OEI41OBqze+r1+YuqA9j2oj4ay0IHOB8IkhoUT9OiQJcbFJBnSiENMF
FrzRDOioJwGA9LXOq7CvFm/O7c3ZuYw8ZADVNP17op6Zx/g7qPcRyjt5s8XErcZGV9gMLcdc0OoN
LdlCrHHPDpf1cW6PaPvBiyAcq16z28D8WXUcYJ3KqbM/y7wE+FApMomRf5dU/qPx0QFw62m8XRVF
Vw+ZmsHF840SC4nvq4eZ7P0m2EBSi3sW4M2BRcQoWYD/yEysK5yp3ia8wT806DZ5F+JikQ8qRMp9
rKjfjpCTP3U/OYWnI8r+V+mS2mpaTxJ2wHpxDVOSYC/6XvFLZYgmSbWouiWON4U5Hu3OMVTcWrrS
bQ+LvR1P/HbgPJDY+emxoubcGKAd7VH6aySHdrauyF+wVxNN7NfKDF+ywXxEempMuGJ3dL15/uDW
THA050kDW1js86hxra0M2JL3+VsEQ7HonkrlN/uNd/BMjbCK0ACwwDRDhN0fLAvgoUhhREd0PKMm
AXaR/5Ru2rdCkFI206zjMQVLd0IOY9OKxCDHamZSveZuAwWgy8SjbZPBMqj8LoZbS20jc6SxVVDZ
bRa4P3AvIieD95WlGsbtCoGwObnGEbFKjH2BrxN7kZ7JYaMkNHRFpaH9fICA01AGczRZgXWceFQr
c/zGhlW8kBs0z9EozhiVdAhHL4hEUGtBDn6OOdqDXztg5xOQtW10ywwAxs+4CkXnbCA4lOPApc+L
QK64Jex6rz4ADfFpzKPlbchCZs9hqdfs7bvlRQA4NIT67JlCPA140EsRNzmNnQCUA+7OIKYs1ji8
q/quo4vq4WxITeMspLBaab8mKvAHVeg0JyVezBUpCr7T3QdmUYmttbyEK1elsP7zu2xviIHdevK/
yJQHMkeTXgkEeEyvupQI6der/4MAmFYS9V4tZNjQgvACCcjOm9t9d1mwiIN7R1mcq0soRM1ZZciX
KNgVzcjrbTve96mfVe7t7ixn4dJpGWgXacVSJ+h1IcdzlC2blgGCWUgyJLS0dojiABtK977KQPP2
o6NpmLWrXh4aMPDf1WjBzD+O6ldJCvzYmCH2POZ3RvLvy8AEbXpCxPZTflidirHQ5dCJXUjxup01
lqwdrUTKLMfIDn5QL8GqGKP1CIqCB1sXNyVe/Rk7jjEqKmuqEnie+S7Vq7D8A3VTHgiEZHxGwmBO
9k0784VlFOWYTbhJ41XPDqbX6Fv7r44GZjc5ib9krgFpi8jsiM6/fsFBrpf9bmfKrYjHpoIkuSqX
qnRVcbf/vBfeGCL2qRKMH7hCmqud+wUjGe1EmvPJcNfHZbU21IA4y4Xz/wgjVQrdfTJZZxNGKmXK
HHrjJjGSWXCKO7e/FcD1mzb/Md8wntznaNB35sCinGF2eNP5KRfvqCGyJX3PCKX/oNOHctVzuVsn
7z8CgjOu+httffal5znN/cJSmlTSWk4DbHOTh5IFqzsUpQ4NTgr1HGM8J52qFhFVmMxuLj6Q2MUv
0y4D6JHoVZl7Cvz+ME1qTiF595Wn+vG71nxwhVcuXYdvuGDsld6OTUO3WrIWG1gIqiOZ0xR0piyq
1Mm59XapaOKgdJkLjYxsMc9rvvK89G9ZOjtKa4t7+LifwX/r4m12WxtYwsbZmf29e56L+pjuNZ4w
3YKKKUjyDnAgHHHc1uRNInIBTRp+8bN//gdIM7WjkPRk49cXwcyrAd7psXDXYYs/AL6sys9ZbRuM
UvSUgvCpRb7wFiZLTrG56i5otEQhb5DwyqRbKeO2Z+1fuuzJaAWltYBtnd4tZeVa5225VuoWD5io
XqoPn8YD5NLT/oQQ4agaTAsZN/PtyIc64uX5e5fyW402iJvMRXjF7ETZJojJtZKt/pTvo9POOqpg
zvreGLqSl2DU3DmCKJUTQIY6yHOa3GsC04+vBiYfOOYlVHsGEzfvMhBJvrkwAy6EUrdWrz1lYf+z
5ION318clAu/GiFrpae+5rix5rDrHhUljePaJ4wThADLfW8x7j2ptZE0tWeYNKw15fs7f1jH/X5D
fBk8rVc2VOOglE2JWuZawJQgXk7S7ZZrg7H4207P2wc1aEEyCDds4CgeN/qs02xIfrwvyj/2dzlN
J7uXfZU4uoG/FBMmkVODnDnrQ3NeXyCru0FcCOSGzPUGP2S1xA+ASMmX4jzRJre7ixeohp3+DLsq
T44obiequBIcMWayaXF/1IRAuOeM8Ma+qWbatzITdVqVjeLGHbGnXbZVpxTPhrAImiMssbIXhsny
GG5a8h4GGeKX3A3z26gP9yfcOjQWrVktaWjWvFsXgBNoI0TYId0lZVkIW4sgDEqJbHGKWJDXhQKZ
mEcNuCVEwQZ/JptxwY17OXZwGbedX6aNDFiWyF4/tcVNyc66dZudKxNNyu1wdnyxaPAYvQnUsoKJ
yYXku51VOTuAaEZMAZgkYiq6HK5wkpFDvXQphCYHgIh7F9F/d/9xGk3KjAKBMILaMftrnC7l8aGI
CGlvEUSvokaOgLM/qRcu+K44h2c42veVMXrArribsOKSW4+cv13DRpdGWvf3sRDYcNVDB5HHAblB
6oE+Hj04jDr/rMz1h8HvTNd4EcLcX3f8l4DNv14o952L5oxJWne3FxIymVZdTCOwreT1pMh/JToA
7ArUG7rhzF/4uZ1n0EnFkAl5tc0PcKoPd1VNPR/Z5Ten82sBxf8fVUOpHKeRmBNdSZmdPNvuDt7B
m2huhnvPPOyUw9GeYp0x6Rke/yco7HWFygs5CAtvsXXWosriGNKjnSqr0OeqSAOCRP28GkjXghRH
LPEmWNve3bdzb3h+okRn1CAf1mv4IxmDXtUqfI1An/zWztH/Y9pQSzvubB9cFAsKS0X0JKWZjCY3
ufw5Gwzf+00ILdad4db4bi8S4bQPaO4loq4HNuBFBDHpVPbT2HRApfF6vVqy12kQvmgQ3Lfvauze
4g3nRA8YhtUVL+tX0r+zmkHNVGOw0i9CMC4mDvz1OdX//FNQjGnI9KE3DfDs/d3amkJRcmRIUOr8
P6CikzT3MGdufipKMpuHCGqx008N6qAqSP1i7z3XdYKqce5ArRUqnege6xUM4/Ovqzrf37ID5Q+I
8DXmrRhw2BlsYby9YRdiKL7sUYaDpG3jSUvFCiqOIfgo5Qg3Ii2NbTLmQjLAkqDu9za/i/P1fi7g
A5Jbjk+ke7qQE2HNjX0PR8wUQJRFG6+TmDPlfLdCAFmJ5kynjmAITCragpkD2IUQzVwO+IooBLQH
guhbKvi0eS85sTLuBxRqt0Dx+PM6d6OkEKmv8SGb/zn6dJ7kvxjJAeMKxwej+rh09syRcuRPfabe
F20vFieQkVlkl47ZsV1TYFKviCIPMe+LrzlbN6oRDhGtSOavU0/mCHYETr6b79j7y/5atAm1TE20
978zYF8qvzu0U+zzLc/pO5xhj9ojTYQxQjUcWiopAEV6b3w9jPPsnZswkFif/Cl5fehkb7v3xHrl
Pxzklf/11HfHdRt39DV9CcP4W4QuOGfdk4Jc5+GvbfOkvH77Ulwe1fQGU3xysxFi4fdzt9wV8T48
smXhHU5kniLUz4JK85AZvBYeIuzi4qX0nTLHTiU4rFdOhnXy2zNUnZt5RdII4oIkpE9K16pqIVh9
uP0gnbUEZB0a8fwRrWf0Dglc/3RIpFq4ferzh9DTpPJp8S/4t7CyOQsKkp1R18231eAWB+GnLx4F
rZzTdRDJYk+WCZLMHqKaTB+VCVu+/JnnpGnqJki2FC76TiprI3CW7lAisxhkHu0c8MK82Ra8HxHl
VmiqPzRYPogzQKqgwBEafLKxfiib/a/s0y7QiPEQKX5Ucaji1DoUF882VB6BmbNTYYgQ7uPSsK1z
d2gwbkaly82xxV20HcH5oU3BSDrJC7fVB3W0tTdXRZl7BjDGHAygrqK2HgGEqRURelESMVi+sjcz
0ZoOyJQrnmbsy7NVh9Moy5SLhqiDhAMojPH8T+6ic3rqAm6D4PqmuLi9RqvletLr7gEgqtct0mmh
1FpDENZvlvJvZfDue0TEvCqUCBntltU67ZPPxgzb02vUBUjeI8pBwko4SvRboDwlrA8tlf4Jt+qd
tWC2SWJ7I9bpJPFniwfBMHMpkipAAYV75LoRNg903nt14XJDQCX1v7h4OEeYxRMVAnbEMzg+vNSB
n9m1RZnpqric6SaNRy2QIzfcaXA9xd5EAuerBCkHBPJ0zkhAnJK+rTJyg8ztWk2WHBzqXWL8Z0dh
WpkOHAwpdIG/eWettGf7XmF0nhqK3DvsH9OhGYDmo9u2JzGsmXkJuw0OLPrNF4eUx5DuGKp/VT7G
CH5dv6THp7n10rzvFabw9wgqDXP1MFnUhmCsfqMv3uePRzFQyM0wWJJ5cPtF7bHnBoX23IjDE69m
B+qIiQIBGqliiII85HqBkBVFBKOxVRYe8lgUbEXKSyCBFNg3hZQ/0Avi0bGVwC9hmT5VhOWodjyQ
eIsAbD1XDrCbBrx998XYmU8QzlAOExP+j1b2jSEfCFtRyu0ngxm7E2W7NGeqzp2KjqCucG5OXjyZ
1owgBaL2VWTBYR5icAGhwZt5ElTgobpgnXZeSXnyslWDXcM1Nz5Cyb/zQvsLmRY0NR/0qdlBK/Hb
g2OmplHO6+RfbnBmUiX9hqA1autCVNUNOISyLfQ8asy14N0pdMNDOSWG3bM969fveUMA4hJtkNSi
4W83sGOEY+SVVRfakTne1rG+wUOedxDQ+Wii1NCY66NCOSj0zCg7GX1Ev5J6y/PhYBo5AHeQvEJD
MBpzC9IKw+NoxqihJWPA0r21I7Bd4abFfZVfthCVrd3sTEXFoKA1uZy7hJhy7GkditR28hndHK5z
b2x/U0ky7e09j3cWcYJVH+fKKUHH8wCEffCDkx3c1g/OwFbUaTowCHxh3/ASmVC1o3N60NB7q3zy
yD57Idr2Qx7fQGgZydQ76MpSXQhL2MCe+jeX5soeFfkW9pnXZs+WUnMYykBKjfSnuFYBpEtNLmGb
0uQg9R1BImpTovRMs2HlCdAZ3dxi8CK60VJ3bxM5ke5eGRNsKbgoRaAIE6/2/sXQIr/95+vZZFh6
vy3Ab2RmqKHKL77lju/pwBnJ5bRd/ZVp9I0LeWiaA6Sq1D4UXusbgRKHFhYXcxs1atnw4utZMzQ6
m3MxWd7urPQDE1dBtDRUoMZUP/gsSuDY6/4qaQB8JpRh0CckjxielIUCrmzmPMh8iI6rGp3jccF6
q+sgTdgW+xyLuEE30Wrvuph/9omv9QZLP+ZbX66yUyJoXL3uU178JkavQhmEjLLP+kj6H8mMO+vr
AZp4Bdjk0Pzrx+tugGtzsgdvgMUQNjxSp5f2T7xnojfaG+ZWb4poHexuClvFxwYPt1u/p3tbifeC
KvNUlbRbPZIJq1GguxQ7pjKXvJQXSJ2LOYiIVGaq56W4ZrbS4Pej2MwRWqWA3HBvhNDTX2uZTuCX
H0bBT8uBRGrXzgM66TTtw5bOO6hMXNTTKuJE64yzUPVGo4sQXk2xnhrVAtncnTm9HZ6YiO3UrLWc
rGZSqjYh2sOoie8e/Rh5JE8wLP6STix1W79zu9Kd5NeT474h3bhaFNLINU7yNBoX0k46KOdpPvzC
dgt/Q8AstSQ4+eG0MH3lZXPgiWQHhF0AL1sFm3nzvrGxUVUr5nsTi+FkxG/L7vhEIZcFn7HNuknX
Ou4jBg7AhvPXQyq9BZV6owx3A3XNvOI6uLe6KNyiWFPs675eZehj6TXPhnhC0KupamjhxtvcpvF2
TwFVprkpx3J+EezrVL3RLWVjhF3SiY5bxd+hMOkGVe9z6T3NJTo7OGc8H5vo0QqUjtdfIrlZfCfL
XtGmB/bmMyY8ST0INOHYZ/ZaIFC0ST+VDzA69N/EnuKKv3+gEY9DMyd3h9TTwVew+m7jePd9sgcB
g+cvpz96m2tF+lz9mTMBv2Qpr5szpegPKLM1pC0IOLFGThpE3LtLBqklWB0x3a1MplalZQXAEzBw
dGcPElD7gSXXLsX6A/ykdFU76ggHh2xVoZhd4vDgXSPmhySpEQB3m/NUMFMFP4MBnVPAX8TNxBmR
sPgTyRdAcEnIpMvY37rm4C+VqzOY+C87oUxQsp1aPheS5JQbHC1KF/V/J4fa768ihrap4pVvO+TX
VjdmKpqXNtzElF1cSMk5AIfErvJKBP8yVMki9NkktbnoXwEaxB6os0lZyjMa1351vam/MYEyp58i
PMTFREO+9nG0yYcMhMHVluRLJBTJ/oyPbPqjx/haRCFToxKEyjzFlb5pQTzhdbqT19MjQn1KNy+r
EBS6lRYBFPEn+vLe0QnFVsKlMFLmsqJq7YGeDpJu/UNVBCeparcD/KZ2zo1z/EFd6wxYdMZd4px0
/ZnCNtwI++Rf5GRsPvx6FjM0Y7cJYJ3YKbGS2KrrCj7UbR6O699Ii1UzpFR+1mB8MtqdNL+VnNcS
JeozWm0QscphzRRdH6aMYjN3UBQhpn4yhGJ+qKRhmBaWxRUVNr68lIQnW91FZYV6DoKBYiQy8gBh
59osxHmR0Uy3IY6jWC7eqtwVhbcLuqYhq1RJ48oz1WcCQ0LjfZ6uUKwDAJgNsZ9Wf34nHhL5RUHI
ZGwfGIwsIfxlMGSRK+s3KDYpjAheb5nmr0C1kQJd66+PyY7N3jdSO+tChLfhe4l60vOIedQiI7MS
c3iQA1gGSTRh6p/2BosjM8tt7SYG1k1xbiW9LMPzUtb5UGUz+2FMtZ7U3LrcDNSScNupsuD3Io++
w3fcM5pLHV/OePefcur/Kgt8e/eAqGQe5Ro0k2ryPvAR/iKvbhtII+/CE/jMLHuqKMYqMgWI8165
5fJIjQy9DDQJVx5dLZDECORlxwfEU51LOiJ3Y3NbygoDwqS92ks+52nSyeu3DEdv6dgYIitmsxjJ
EtZCjxiPosJHxEL+1m0JQpLcKMva595pIOo+gNrSVl1ZU7SVqc+jyQHDg1SMdJJV+wH308nzWvh1
HjkKVsKXsIMCfIcur/5rpX2Je2brHfodv/KS69dUVRiw1wtQkgdFwYWnxQ51WcYkjOii5PdObDqA
serryra/waS9UE2izUhdWGzq7qTUTAQxwVubd6WBtB2PE3CJGR6flPLq22QQvfoNOmskyK0Uqr4O
K/FrqFCa0gbDRHbLCWeA1QLEw5NYE6cclTUIYyqNtAvfQXvshKK8Hk6Yl1P/VT+qzzYbWEdI1Npw
H0uE5+dtnRbbV2U3d5PYknmzNIgkOkEp8AWz11Y0HNku8CpYQC5F7U66IT+TiLyDG9er9WvCTr3Y
xAu2k+eCl19fECj1u1CNEpet4MnsAKM9tLNspqAfYra2scWqnShD9q3zTtujR15mgcOy0AyKXji3
E0Jt39nfotEmNZSvsoW6U9TR5AmSfTcNEhv2GUHOjVlqnoGhXEeQmUPscPhcfw7kroyodO7FG2Tp
skAFGMjyM/YQAyVM/3wCpwYYp3I0xU8QNsVq6F9Lp3/L+IXhphaN2n93x6uAGZ9Em3K1qfXmCV2B
5LEFmw78uM86iOMFiwTJ6eyp184t3zVozWQa8pPW48Afu5huBv6ZT6wTP5393OZHNTWxn6Q2ym9W
a5KSDbusNTaOetgEqshT/qom+1KzKt3nwaplg/rr7K06FZgC9uOpionOC+wxRM23bunNQyauQKp/
WZ2VfysSPDhIuTZOXbwebcjxQXJ+zudwSFHTBcs+rhmfzsmn0wwTsHQqUxNPHWxDBAGzRP7SPMSb
cs2DCOwfu7tsfTAgR+WVjRS4iauD+iw+p+ZcCza/1kj1+DtRsYhtxZpkNC6Khd2bc+1O9EhxHHev
sAlhobLT2qJt96bMCDwqXps1lEyDGoBC+pU72MODEmguB4rrhsiVmU+ArhtzXwIQaQE0zcIWmqT2
q8ULEkLk8Wjk90AU+kEi0Ilwx+qg6sTUj/nvj7ha9wItuJ0FPwoS5UatKlaTmpOPZU4MJwB0B5bg
T3w7PCeVd7o9vexPuXYV+n6vY9RieXRRPmQi08GfR01uI6xHbeI/wDpQ+C3/en8OUP0as710aEc2
6bPUX9wsnAG3WAJDP9yZB5DWeYy9xfsHr/LyKwGEQbO7wR6HhGlXoBsRoHoVmPgxDWBpVlJjzs12
4h8YE0L+XMNy1nkG0Zz8uy/eMLNpmnB0MuKfqHfLP7zOu/o5cE1mOOk+SHG/ai+WkQPfT9KSH1EM
xcfsUbsaz03tyUKmLtfugkomVjK+u2Ku2nhN2EjlZzcd/T8538nSvxc6a13NtxaL1JL36sarpNT+
tK33flV+sxdUIML6E8D/AxoYfchxDQWXkQWMQAEx9TPL5Y56RR1+VgZiGRMHcwDj/hsNQFWqx3i1
f439Dbr64dssSiv8CjY85pIrH58iLzghdTIFf2wTioG91AhoGrMCvD8N5356Rht3WoKOhzXuK49G
aZf1plZkkrdRD63urrLDtX5rIQBhL7w3ZULkhjekIcekuXawkYLf36m56KTmTJxFF6o7WpC6CwHo
Iro7rWS8hiiyLTbwBNH0EQYhlmqkN1Duecd7V2VFT9PSKrJQlwta2Vz1KCzAA2tmjmcVTU+t7dos
GboJhXJ6JaFGL3XPs8adrvRv0sNFQvqk90yPTiySEDpntvJDzfJ46Q+kKuCssjUMzLaup6bFTZXi
Hx6i17/sudbmUwwOFse/QWg/xIiJsabkBsWnhiXjt8M2/DnwcQ21cPOIIdQv1h4T5V6cjN8CYCjT
iGL77x3gKfMjfj+1LyLsJiZCw0YDgylRrVuBHXtOWR3N+ib39gE6Bio0CZ4Otq1VCe/qVTv2NU8z
XtqKthRKGaJXjIQ9tsNanLun80oWVK9+bwCQQwtbxvXNnRiHpfwB/2SdgWO9IYYKYQgfFw53dKvN
nbOimFqEpbxt1BUKYOA9wtDxUOKPJm4hTj6HJPACRj8aLTCJ2ht7ntaXgYkCiZeFTzH8MBP9uf2B
1MJyWGpa34qRW/1+byoD4d5Y1xPINgZA6cAIPMkGKGJmam2/9Deg4/3PFRnFxoAnXamq8SiopyjX
r8FqzfDvup7qvUyS5H43DRMbnEFGlzMPPBhkrp8nSrHCjoejz2r+aIL0iSgCnax+KOaPlHRiRSBV
A6uE0+/rG5Q6buMO1TGPMmgUiZT3A+dfNUqpbbvhtdLVtfGvjfCbhWtoJiPXy67+IdXzXIfOPDge
5xWCCuf9Uq2wXBhsnjsZ2aMu1kJlk9vQAUYrqpjUERRjVPFV12DVzar2xCydVQTP3WEMByktC2A3
cSQuj6wVtTjvnDDhDPv8Z6792pTkQNJ56nCbQZxpVeWrv2tc03CkDNxbjObj20o3bu2B1KlCwK7n
i27gy47eXHObBqiGmGCxGmtp1GrhKOO4opM1wiIXB5W2A5vcpdqBGuqtfbDZxhtgGPlv6TH3DJF7
iBh9WGqgRzwvbXYna4Vj29+kA0CR+ZQPSpZ9ydqtBZAm6YummWIzm8EWgHQMfa68BmEQninkpYUj
rVsIQQN6sOFUbVewu/sHuw2GToGLIHim/4E1J6KZy8xq7teAD22MigR97HWFr5twhOrNPb0MeRl0
wNEq5aUWQP+nDs1jAj/5a1ny/ndBmVrNUD590//vZCpiTuiM4dcGgBnXfpWeYeaAKgA0KaOZsINI
rMHKqPBBE2XOZywtBj2wtIMQVEAQzLEQqC2rPTijjnwv/MrP4USFPRAtajo/RJwB9n/bxxQa3SDm
FIkwpdC8emkKxwwU4cllP9aYmpmmt9fU/lEhU66JaVGEI3mIjfXx4eOf3pnkSsH6aANx+QyVqL5I
mqsKF/UvK7jTwbkiFouGg/XFgym0/AyhACdtb0gz+lG8BtX1x8xWYQ8O4Uh8cv03BepoA2KRJZKq
OMXO3Z1KrwKq/Fu7Czp6OqaowkGgJQZKXGDM9trhfJT4uEqAUV6xbiT9KQx9ZYdH3ptB+ZIsSVUq
uEET3mTYiMEdHDa1Eo0eP4BiTc+wh0elEj1sOD7E/G7inCvHoIt4fyqlxeffWFG1YmDMpHOi80Vc
9MNv4W4C92CdImoAi3lDl4sejlUQIsWXT4utJcNz7iXhHDCke6GeF5nwsEP2rdwvgJx/Gg+/TBdI
NR+X6KPlL2CS8llVmy8PxkhaqS93oHyUrydU0VRD3QGLP5IugElwHGixA36NNVFeVb4zftoCwZJv
PIT3xYjaxdqM8aBryxalRw7p02r9phFj4OF7BQLttFvAE1emVhctxp9PRuluywep92+NE/+2a03o
NR0mM3WkSdSBQNZruXhqHeEF0w4mpg0LpY3kfyjLEkEigLXuw2f0ZRD0eE5D3S5vckpE8jGk2sN3
FSP5fw97sW4tun74GkV8PxFfeTmIBsTAsDtPppWf+pbEjKJETQzhSY5VzuRb+wBe1xgd76m13zFw
AJxxsBhp8KpcXp9NgCydO4nCOQnM5v17/xniIYxpz65QL5Dl+IJctkmRUECH9sEvmrnHjHEoHXFL
dGcG9CpfCfQ9kTL8DsgCMRwFTgilsytZAKDJtxFyrPF50DPjpWQ7bEUD++I2VmgoYmOCgnsiJFCp
wPw3MFRp9PLhOYdfL+Y6E4Y104N8z5UmFinYABqE537pDEON/XRmJF+MT/izNt6ieC0oU6QBRh6E
g0Kcq1YwxdO1qPvJcaJhxHMpLXW/40CyRk8dprpt4mjya31Kfpu9rXEUoQSib1mjYjoZ3bYnB/gF
ZhXeSXWPnkhVuhb6dcVR8PqQJE6X48TIJviQ77N5i30gV6mAHrQchvkQaJVxbNLIQV8Oz4gUlKzW
EybPos1AfhznWoOehypD2tTkXGcgS+/+wvIz6rsvGxMdcTnhR9DpLQY1QzmfW+CXez8/3OOL+NsO
FBkBLT8uyk900NxrrGB4h3ytAiBS1Yzr7SqyIC2pBqxGVSnKbdTUWhEdfgRwWwb2LMnAz/1dbZcO
KoDd3hYKCLhEXzExZqn/oaVh2dtJWZo7S8IpRJRvTVOfa/hE4ptcU6FfGX10++WCVNOXg2ucQ/KB
j5c4wmt4uEZ/Jk2A5iANB7zPH2xeD5MzELkx77r9T2w+m7FuYpXe49OterZ89/QdzyOD4WlRyZLw
VMrBUJji2xuev4bDH67By3MzeO2suSyPvo51mIJ6Ss2e7pePRBVMrYKB09ZmpSb+qmAheG9j5YOM
V/IyAO7BFhAFm64mZJA94EKGC9aMznqja1hlePrxeLq/q5b5O3yGdGt6DmsgNs5gFUwwTuFmR5EK
gpq2RT2YdEhasw+4ad8HOaKdbTQXhzRPjbHhhprfItk+BG5/OqJ73ZaTdpgjLfMsxi8QKZv+dsmY
GWd9cNdiXArXqDvHp0apI7U8fSgKGEHDN8KlWj64INIOhAMlS0X7lKo4jnmT4Dc6y6ayGetE+mx8
Xnt9yM5PvFq4zePKaBO7iuScyeFWlT1XLpax78Zq6Q6bklfHcxc8FKIig77ggI7qQbW8mGTl+HYe
tlbl4irBzUWwwyFQC6Rb24dfru4mvoZ1sMT5FbpxqqBXR9lwOCEQUOc5gZeMz7cgNhlGyJDcAWPp
9RL+gsz/nHRq5EqRd6abgMKt1hUSpmxl40c6lP5KFPJXNS4R3SSl4CndY86rGYE8AxLM3XHUqOj4
7KWI0g7WNUFpvwT6EjOsMPtkQbwExWc6PdXzyYCKKpikdREQRvFSpRU6viL8r+pH1BcmcXYrNp3r
uN2X7l0UvoAP1NgvOr1RJr2gBYBmzTudMRDcW77I7NZtiHz3PsOLpgyW353msVFgvGN6uP9vajZT
M5mOPVY0rsWsgjKbQ65Bl8WFG7780dGwYoum14juQhhr858vUeiABdPvqFO4QjroQwOwLNK/+idK
N/55eGR9pQ8E98IeMjC5kxAN1ixcPnVvJkVAUqZgxDLzBRvBKXs7rjgMHI0LUKgNWrsq+DCsFoXp
glxqpdVrX7SQF2E5bGI5dmcxeROWoUEO+PbiMG4veya8CmkPs1FElHy+HPhkz1dXG4P+weISssQu
NF3AszcBkDn2s4FultlnWX7WwGXmza4a/XXpyPFm+rdV7zUogpS03HQG90WVzC66A08YQUs8lDmf
PNsjr7ty6O6xERSWrwQuEpL4KNOdR2mCuAPv6gRo4hkgKPmhgTd3928G4sGPXnWhAe+wNsgYqIUc
jAfeBO1KDS94/TIFohi4fHaMse1xLI0AdXrrMLoglk7XCOazfAiSre0ErlYWRZ/Tr5vNR+aMdHuE
4SwpKe1Lq2eb4LbD7PKmofv+FUZgJw38S2dhAYu1qdVo2unx+4VkeaV5tZSo6/KAbE8wVUT6QUpI
YdOcU70Y1Nkiw9X/TUVhwLOYzIydJSaMYwOq2FTbL1Zq7PQkjQ+5kIujdX+pmWrOfOZHtZk00+0S
OB5DolaCU4KC1fsrBtqCWWegc5JW226Nz1jbAYymmFHnFEnatAJSd5tmWIk82iUFwRicXOp2a3rR
PAADLh6YQyKB3qnyb4HZAwG9IJ8dbC2c3pPwBBDFjMqeQ4VsyQ/kDp5MQy4EWcqovBfjuFQAAivm
EI6OOEF8SGXpMiVqsUys7lOQv+BmdCzpZN6esUS6WO69aQ5ZTm6ocM5mqs/YnGdR/h1xmF+vj1BN
r+8ELiMhlMRpvIPpz24ZrV7bOZUuoXZpfaJ9v3QNgTA4iukaTOYXOocMhmWsF8Iqdgt3DGphlWWp
ttMFETrIi9eGdDps4I7/Cu+6K4LP0syXIr26TLg2G7wVGx1udzWW+ZiQDd9ASQ1WH7Zjl+RPRXVh
/HK92fSiYU0UDqPJ4G0PKvFdPm8iCYhwoBmEfr+e0zGjP1HKcq/KTJcCnc0sUmguQu9BruChXCKM
xFohMGb2v3OUZCb8eJ3ldkAYF23AOsoa8F+MorDRwYx5iZ0MhpJvAT6IDVDE0HtFL3iW6opxcKbJ
zWOCLdvjthS9mbNw7HzhpLgXRoeOYh1TEII9GDDP4YVnjvDkPBvbnnO8Sc3CD12F9o84qun5gXFi
uUzXlghuiL5MjXDhvxOGHQSsb0NsAUA413kfB8gRn9ga0sqfBxUfMG9NrEgBWnC1Ol3Q2C6xGJQB
wmcsssFNglSJFodW14CBAp3HNTRy1oQklT/xaAiWZ+4D8APlmMA7m3ianRXnvKZx4ch9OBEddS6x
6fXG5WYYEpIOcsghf0AQ/k170mSQkcyq+DRgZlfrcURrzpxXhDlvznt6s6Y+cxBzGgK2WofhIF4l
Vj1jkwBy/vcCdnp7zN0YuAnErpHxhazRJbiIJ7vcVuatjOuvFcrfUcG2cpuCsBPjZlxBtbSU7ODt
75sCjg2VrOsMbtnk9YJPra6w1sujR34+RN71102M/B2BWXBQKwnnLfSbBP28imT6IS0ZT9kd4LVV
XW8zuzYPP+8WpIgbCAz3nl3K6AbUNnqNWMhkjX5Qg8KVHJXMbL1vRUyh8Q+2YJgagpKFQQ+yJTSi
ybnpd2VwK+9X1dESbwvC4n43Ra2mbJRL/LhA2q4Q1PzyP+ux3hhgAdOQnDk+lvTVkXDyg0GyUEkS
ECH1E8qa0YYUYHCRwtIxZrfe/Ki7gKK4Wek7kB9G3Np/DisnA0fDMuJIHQcxqfw90887O/hKzNEh
EZIdQ1iDPnU5C/U9gb9BrEkIhfCWXmowmljRVvPzpQPCiLETbj5AKZmrASQmDKbQY9WI/EkzgPjv
J1BqQUGnDfh+ChuGLOLoPggzo6yLiF/0kEoMnIlffLJ/QuaSGJBz+M6mQonYN2v6deFnZTq2eQne
8WUqg4suEs2LMOnlQIK9xjsAR63ijyrCGupGM0AUKcUgEHMQ/HdJqGKtay/TxFaNLHWyeLuhiUJk
mcP69xQdQbYo4T78APljX/tZKEOiXRx3zjzXLHQhlK+4AIcccFn4w4LH9k+7MpWQuGw4ySHMFfP8
sCp6qqqLFc669DiZY6KLm8MyGwR7hrQPuy6nW4RgnW6YxGK15mMlx2yUyDPLKuf3ClIHZBnAm2Cs
hsNwc1UlM/GVaeO9dOrcrVUrAwJ8BeTwBu2Zg3mvxJIUFV8nyzuZfVwuVILJyYO43+ouQR+nzOgm
BjRHHwZUxWU4+/vY3km+tXrUjnBmMJ1JM82z0iJPXE8PmzOIcXo01E2uoyFz6C0K93tRrkJy2FBN
WaoHsEAsJON3bC632fy8kDLOJflc/7vG0EoCzNZRwGtGOBMpRyIGMZ7JzzXZJHQz6AmtwTqYKSCX
r/Ejn6HoIWgZxffri9Nlo5sVOtfc+qbm02OxKpe3rXxxeOwrYdvQMqWpw+kOfBtvDF9xbRyKWB6H
Sv+v6Ctip15J2WIue1pd8NkGkEsduqvDGvrdKVxQBf34pPQxA866dav3P4pAjmx2hnZ6mhIXAhrQ
VwiHMPjB3fHCtywn69n7xIsZU/VbEsG2uOwxX0SBOXDhJf6Ke91wgCCG6Xo3C7q8E3c96BWu7ytO
BnSuk30ny0Vvpn4s/Jhwd1Tbszxg1DsOY6Nt5IJy7LNDewOJUCqK83KP5pWtCzxTTYKlaRXFvQaU
T/O2xSBld9x3xQh3XKCXPJ2viW6NHjnnqnUXZmwEsibB62/NDE3q7ukMPkQOLOxCvm4SxyrdAK96
HmZvVf2BRHRyNbZWYimRgu6JQC5SSBc8llFMm/3iDS7DU2hiN7/0szGq35nNsP65s4+2jBS/3a1+
sVZRWtBpWcGUSqCEnpj66YrN6g30Iwi/h42h2QTKJBQV7heUiAdU1UMrMj4nhkXEQgONoa2jFtyA
7imnX7RPE4Jn4CnczjYWq+8HkFy4R5EO3Eb1WuoGq/vjNRbtW2RxHPJm1MfvvmjPKJETGoTdqm8+
8JHsxML7RPZtn1zGH+sPi6S7xWAm7uMV/t0SONy2mmlq1YClk+GhW1NTUMGhbMlkl9nziAhfqLSz
4d8OCvnQ/AmZVIujn8BwHE4zptlhIblzemXpCGOhkg8T6I7K3C/fiiODDtI1rMW54Fql9nr9K69G
362CE5BpELMjbDIPutjNw8g9uwTtv2orAiWX9WAEVe6+7vsRW0d4Fka7RSDNtqqxqz+HhC7o/Nsl
QCbWMSW19OTG9tpSCFDLaBMAyotue247G6HBicxulrtcrcR6BwwRPnGbTn1XjqPVH7eTDmQMtuPD
tNra9DKKLdbDCZ2Hv7y9bkAwfraR34aPxVT5AkrAixeXqP7kl9nPZQWG3fIXPjBO9h8nGPdlVDvA
ddidO8WU5cdTjTQ5czPLyMjgy6Quu2d45kkm4Ja5gjdn8I+Vc179ghfmLmV17pSlKpEStYNVOs6P
4C7m2R4aFvue2G92d0XpOon6FDmJjgVgBFOsEjPV0miT/ZytwWaaE/8dqERtNi01fqoDm9If8ujb
5EJoAn/v/g/fyEyc8gQM0LPpkrWTCtzi+3YdHHG0MllEFv56pN588wGBf4/wsnIqd1X2L8fb3Thq
KmJNV7lMb6NjoxyQ5abTpIicy9kEFXdbq/pWOCLXSZii5sULJjnnhQxSH8p7ai2E2KDQENRKuTq8
siijkdovlgBMqvuLqOpzZFM3majcbFeTsgRRyxSJTv75/4V8SAb+PMCzUN4bOiNOYK31O6UcgqhQ
gm2PfDYNM+zIWNdAKpmK2DeZHrR74OXkJ74ybcpdsOdfUR8rzcDzoQE2HJHPKTvdgtLAV7liPs7v
5U84RCh8M63rO2QMeqeUmHpH4oUnwVkSR1xXth8fsTQ9X1eqUx4xdW5u8oHh4kxTJT/BNBtSHdht
kQu6wVMFTXN4HaYa5PcQVarJn9tbAfRXXtzmOJOXgBlaZQK5t8ScdPAaXfbNp+xLVxdr4IHA2lcl
ScJD4fvJM9r3KDlx/PPMGltBq0LnlPGmzpHS7smYys3RLEDRoyj4HCezt9HV8nt7qzCZzdvhRFIe
x6DVYAxa0wUvzDkW2nCu/pNWaxc2WCgZVKGLQriWr/f6sY4X8Dn7GVLgTV6Ssgl/0fyO8neQo/AF
VV5YNHgcWmdB2wpzBfgOCuvJ5s4YogSvNq46lIi+O2PxOy0Uz9rTnaIs9UBA1+VSDQVkP6DbPnhV
eaPpkl03BgQ3rHvGxYFbvJpgINxzubPm4fH3wdt8Ldc07qSewRSJNqBXy7Vp+hp3PyNj7r4TvGaX
DxdcSGxYhMBIRaMvPzux1qWXb3AGdj8+h7ldDPUFt4bfxwtKTZNIAWIv5r9mCist3Ytlv8/7lUSL
mBcGS+MfjZqTOWclF++0UeOhDer4dsUHpkCt7gbxvTYgnZykI/irVaW3pIjv4O0ukVjfduqGGLqb
w+xzB5GuM0gTbE0RLNR6pgcZISviek6dzOreaPzzZNFvEiI1xtQfxkYR5FtXQy1qAVLF335jtfHn
bqOK0oPkne2ecL0GI4DstCwN8R0WjuayFnHfTzm1KROCSDJJa8qse/CcjdUcrlihzPsoTCBGTApo
Ap70ZZPQJ/LiJsY+APFbImoyvAb+xGiavgG9Di8HaQgr36phfUKFmUMlugo31WpWAbs9nB6G6Fbi
lSX4UhQ3G9Wd/BUjhuvu5/EsL3e2yxJJxwqxH9tpyXtmZcK0JJ/kDB+QVPZQldTKAgHbFDBD3oIK
U7yhcm+0n7XGbd6/YS9UjSttwK4QP/B/D3zYFYgtyDEsILkyxJhyJV/BGrleHuQqZFUkISxzw3MT
yPQLtTfqXxEDyILiLAcDrn8fxXRJmGPtkcycg7Vvi2wEaUVZYKUEcIXOngH88wdT0xAtjhRmso7D
7gAI3r+jdh5egy9BgRW1lTMiAf06WCTY2Q+4zh3f51B0Gzsd9Oc7lEUSzBBxThU6eTHSABwGi7+r
BIeTYLtjHAnuFBEg2aHFicrGw7Ecvusy+5EqRRHoLilOwP5QcwYkDIy6Jk6uPo9bx6IH1Vwoat3/
gyDYSoovgu7IiEDaEN9A+ZxRDZNcJoxwnC5feNpj/3xR/0FuRjFdFFzdzqjOLXl0VvfALIpT8ZfB
wCiAoyq0z3gsW8Z/VEDT+HL10WexGsb7HDYM/lMDLlcRJag2H0UfXy2O6fmNg/ie9EGosgbfAIkU
Vel1arBpAGgbJFVmlGoI3S4seHfXt2jzW4eQO8QEGy+jFWSwlzg79L7sI4M+MXT2KRzi91PHNMgK
570Jn3tf9zMq+l/ntavdQ0shVtFP0xSQYrReLpVYWV/UXn9Pwbt7/DxT0eJPhjmCFJdhHWGc7sWf
2wXMLH9FXVISyw68dKmMO+5m05b5Uqw6Hvw8LQoM4ehkzQeE7y9iVLycKbike+FmH8r0VYgfmiel
r7lu7QQnqSs8XvSbfpThdZgYqQ+KWFA1tVJSVDR3ndTq2YC3SoJXZIaihZlOWo/qLxN5WMjZyZDQ
5qNqlYgqnBklPIxAeQLQCtTIDWu6NP75n+Vo1XNLKDIdV516sc5bcM5YvFtzIL7v1qnAioWbrGj7
K0thj8wpyizx59dDMRoZOGFHdbBa6b3cD2ziWzDth3Z+r5iCJ6XWZF4mI2g2txRy0GUNUk1boo5Z
opP+dwNgEPbvqPGVUoxISz/t553rqiuV+ma2z84EbU2EDZIcQoF4fpJsHlH78+9qlV4gYZvPXZPo
9MsqFx8EIiT/0hy2S5JApdruXfu+AS+Epqbb1ydT/HyPHOdqQD6Z3sCjNvCN75Cn7/vmYQ/cqVXS
R/pwKwHxQV4Dij4B+ig7zUxurwSZ+bC/xUeIPeHxY41pqgbxrfJIN4o4KELoJSjPi8R62fwThhMe
dR5Tv1HxVzi6TdrSF/o4b6SIEVip1JakLUvYMbSgJrLyf4nk7CI1Qd8loaKK1n7JVYf1oV1VWJfT
qaIPLTogsDiKhvAj9xEUij4+ePijLFlPDNzGNiRP9hjZG6Edp/kaPzpFLj9wyA/2Ux+a49Xf411W
h3x4SFyykWXu9+k8zdOv2YuKcuYbckJGt2ZntLNaccJN2tzCQfLsuiU1NFZS4v5FSXnwD48qiP28
YC660u4axWIxZk4mKvSGsoLa0FvHeMkLvmxcCQ5z4uYoisOpkfXT90S3aMD2miljV41v11kM9guw
LEVndVLUL8nsqi/aLTf9ISbZjezJ3+C2Bx+jrs2x0+qyIRzpNhr2jC9t5XHHp4krgnXq/arRd5V+
i1+f8NDX7XWmCZ1GWiRFw7T9/8KUPlOmDi3ehqHhWnBjtCDmCE9mHLpW2cfPTg1PNdtqPZAVjDYv
4TIemb0rVRw/Fvia8muBZr4lJPmKzxxW+52oKDiMAoAqkfa1b82GaAez6prrXb3XNcCXssmEdy+K
4FrONHDHv7eKjAU4O/Et0jYBgVatgXOwiBOrqXfefOh3t8Jx4aYKRjQDif9t7PBbjwJAyygkOklJ
7cUnSlJXOnHJhAfAXBn8gd/5QPoq947dXhAuZyO1J5tn98OUZYRtJXQrB+kGh5EuC+I7lEhlvKZ+
my2PCgo0sz6TPmmu3SyUQSzzy6WFrXs8CJLvu7pRie5GvJL+Koc97B6JPfy0HeGreCljalPLVNuq
I52Pc0S/7dDPmCFYn4gtNFE2I+f0E0EMw1hjqISYgtgoQJUjbHILIKS0c4j8GH+Tcs8iFkV5ABkz
UPsMNmQabwVuD08mWYavdCn/r2SfLAOPPu+Khoh9PjrMbTX2+bkUqBlPiNVOOG5CodACqrJ5YZ6Q
wzFhvW3lBLn2lPX88V2KwX5pvfuyi+7uj7x+0Z2UAtt6VxHLDA39sPsq/41qqbuAznATot5ytx6M
3MVTMLyVfIyS1nwXJQZp8Fm9CDDstW0cxwKPetfba7wUqYQQSsivaiDYEjXqcLR+K19Ads/xVi/G
LwoD+nZYO31s/6+M2xofcoX4Bk5gzTkvui1esdCISfHmOXr3kNcsw+znZjD4e59PBstYrpCywQh6
pJUk+dwRYELlUuaex3DW05kw79sT50uV7SdVy4yhrwqC5voAG6LWj1KSfKp9CQSh2TSI/Q+G0Yo/
zx3+FG2Gt8VDura1eMRbiN92kil/YT649KvrPW/TwXT1VhohhRn3vbEizav6zFPO3QSYbb3CoVTT
Pk1OFCE4epwjNr7macCxmxWEKqNOR3XeL/jEExyoA5/U/xw5GJ1B9zFIeshV/UcAlXwvTqcCNWgT
FBAU2+FzsmwSYBQIZ+B3gUla7ieTym3m+qAfaV8+60qzYsvuZFkeO8Z7fsvZwrW7s5idLX3ASJL5
YqhGHbfa3tVgG9PgxrLr4iZc+xSQKl7iYmG/SXwdZX0M5tBN7wNtaeMeDkiMGgem0fLyP+ha6Uu4
nN0UpMJ8xFWO5ChRW/1QX77yrQiCtYmvDXXfsaFG4lzFFmSc/cby86omUqtrVJnvupuIcpTGaQOS
YsCr/nmsXi5Xe6qGTsm7bMranjnOryKRiq26wzqNvGH8OURBNS++y3lwAxzFVOpQq7+AjpKHVYEn
jnzk82mgQmDogM+dR/RbQmO2Ew8nvHnTE15cEoU74797YqaugPceZE7xh9sVohfCc81LRinsoIzo
nqC58ApdUxJOvzckN0+evInsmXqHAUZg6L3rZVx0SbRqAICzg/M8fl58gVJxmCt8eUPCsWQ++qsS
JJiD2TyHLr10JDoZLtiau4FOtggpDVoyLHMQ3U9qJwOZo0frr6zcwat7sbtZccmbBvFYmvdRaMia
itLkn9FA3ZR2Ar6s3gWhIlcLYpQhwu7+ozBVRSUUiMoqgFROd70OZph204LBly4f9fFYHMbIQ1at
XZopcOTdnu5AO645KUN4EBniTRhUtZzeWfiYoWmyq2KrtriPeQK8tdBvPHLaa4a3nfvMFe4STXmP
+DBbMlL6Kx8G/okYygKV26AEJYaoZYXtahji5hF9I0BB/YZHUPDjcaQrahrMihoryXd3aszRfCUo
FgNmM27g1sDNFvnGMPpE6eOUepYBga46Hsmc1dNEg+CzKbXbPwbcCuZwpq7gqf9rc1vRJTY7Wm9X
ekIROmOo2Aids9jmfMgXkjWiDIIMBKRgYTtwLWZ7roFqI1yFOsh4dSQ057LOTr3guMghF6ZJsAa+
xt1zPOVjbj1aBY9gh1fRFT7IZR0KySSrhYKd+1NB9HpI7A3gKexL5Z/O99CkNylygitThRgGB5ey
+DsMrvrlKapdxZhBtkZZuxjJfBLiZG4RooD53v81rDFEIAtlb6E3LFEANfnznL3YlM0hS1wXD2M4
Hju2jFvMdV9nraRD8BLSYpz2UyhskARzzcU5YkQEnIuH67j+eymDcTxxIlL/VFhsA71LPEOqXeg3
4I0K1lJjc2qZXA5YUFUNP3gE9m0UbxypNbUg84pIXyAzSkNgS+aTCyvqX98DV4Bjbo3LHdrHbaq9
wHSlsezednm2Ec10fr0qFV+tkZ5X6frR+IRtOypP5Dhw2BbOBnrTL/Z0wYqgSuduWYk6n4bKWyDb
6OW5EEfIuGWzai/znO7TNAEu42sqvPzdwXfAbbpAiz4W2tJThVXRq2hVPAKh2NWE/96jv8hS57H/
zk3Zrtzl5XbDUTBfqGG0mc/7FQMZowsURg3mNilEzcWlHBtRR++U+qhXR5dXi8MYqpOwWidCiAPm
yFBv9vr0B+2xeGRYXaNSpQAWCzLzVlyXVRdVE8hkYx7U3UU2/9/OASoGGGt9uC4bCt1h1ynuT/pe
Onsv05Dtw1e8fg1QNDQIatrvIGY8ANlv1tyXPRktXQitnU1R7r6CgCTpV22oX6yNjcFFZBTvVOjU
pqbpUMyl3IF1HQtk8f8ISBEoxTW5dDJeOtwsn97YCgGTd39bNDAF8UryQnpnbfCRLuz+fl2T6AHC
eUBcHYhgYdKfTfJRePMopy6ATc0NdanE1veMP4k+sr8QdeBJODfgD9kwVzFcr/9b9TI3B+MGWOji
zLjhtQI1kF+KQHV1c8K9uSQeHoCrCwpbnqdhWz15YJuYZW5badF+2lg/czPmABv4o6Y/So2dS/wA
QwQO2jk1BRGZ4JKB2iOt0JugolE2bPUHLBsseq/9AR0D4oP+3D83gi3SUG5jn0bZkQmXf47zY6//
Ugay26qmOru2Bzu29kuES6YLV0afwB1oh6u3o1UUfDsMij84XPTAJ7auNoGSNIgjTPXHb1JjcQEw
teCx7zAZ2mXcEclFY+Qp2/leEK/JokKxmGp3Y/fmDuzeX6jdJ02UddPoZkOizfKLNHqVY76NkT5J
jwL5WkrulxGknV/rsMby7vHjvjrSfO5FEms2tZCOw/suJ4VYSSEekK5f/xDpATNkTluskLdLTzAH
EEbmyLaAg9VcbYs1Tc7eVTwB4o5dGjFc1FLU1ENW9U6BCw9QyhRA1g6PjE5FfRBqxbzd0T4gWoms
yoQCn8ZwWDozOuDe1VNmflY2LXjwX+lzB2MjWqBi7rUdJBfMujfgjpsMuGab7fW7Ki6U0xlrdEdd
7y88G2CMf1v4zz8tAesJPyy03IpyX23Dr0aOEMK7JdLpVa16kgVMPdE8ffglFFoaJlovYpzzHhOi
UFwB+8NgJK5ymYSYEnXivbphG0nXSB9KQpz1CTApZPPtgHSa/XIutDLViyZ+z4RZiLKwnYF1s4jE
+QAGgnrMjpmyymH2p/IiZwplKIbSiJtIJSTiLzSBgUjeE/2GBhysC2R2gpLcqPmMVwiXzsrQKAmC
XGU5UKEW3dkCCSXsln8LPeuNqqkt9LMqk4qkfHvJeJoTExrF+aMR0py06KeAXdKUH0EUJOjiP/iC
Xe8uPXiTN6pcTwQRe4+q81Z306ipwuHpexX/Zg37a1bSQpEzUzyOKHbMWOLuSyYWP03T0VDUhUYe
I15xI4tcskrM2ux5WXg7clEuz/drsT5JQ/lGLyK3BxIqGL0pYzupoHvLGp7iL102fdv01C5zaO0H
pAMthFLXhiouUQCtCrAtnMCZZRhy16xfDPeV1iZFIVxE/NW4r9S8GaA/sCjiCTsld1uuRdeBw521
/XEYSpeX4QVSsR1AijkcgUsWGyCmkWCMS1l++nG+S/U3FtAxisUb/a5fwA3n9WvPy86kHgIVhJNN
3PzduaDdwmhaqs9vANOL5j7Yk7ArALJ3lQt8z7J3ZUvFVZlP7EdRlDg8ADnL5VNUQmucYaB+I4OQ
jRrTMpnLtLf5TCj0Co8vd31tatoxyNoMy99TWKwGgZDgFDeGL0BneDd4uaPecUCWaVhSL49/oiVp
iiMk4tlJixXVGTvaJsYQyhvoRD8zrZ2/aaeur/XlHBV6pnOQYIeH7A2AnDh7Pg1FEID/qh2qmFV3
EGJ5mT+Ax+VgCnSrFOekKiitSWFQyfwKRF/pg/3HZRuBIW3A5r7ubhaBNtw7HOFxeN9If5GMkqsK
s0n7EWbqbMVLR1nS/9+0dKL0/o5eqV87Km3Oop/p+y56zqvG7K5LjCeMd1ghzsZPqhtZlKtzz+ax
cx9GlTtJSFESQXlD9dlZAyOKT5/BSYlGDBUzlN5iZoigitxhBA8DXWR0ytyfDMKPQ9/jUkgPHpOj
psVu2CqdINxfBLCoCmm75r+9ErkDyan76XVueT/yAIj5NavlM6SUFrE8jAmUBhzajMcljoJC6vE0
ja73BuaoPUJjFAGCQrnFs7MiHN9immDqHj5sFvNydOdfbRIF6MzMNubcZUAosArdV9OFxFTmFHOQ
zNUXXz/3UlX68n6MUbMCv2v3RGdWtp2KflYGkrzmuiQsvdMoxDVcRpdKLXgXlKRDDQzQMJB2eUZF
5IzoMw5m+fmMEWHKfvvSagMHMMpHcKGSQq1l89u9CYz/4cZIh5D/xsXaYkT69t9MSjxCajDN9U54
vZb/1PTfCTyKd9RYkK3mv0oqv51XIWYwhawXjQTr6QiXMimsEwomiz4Z+VpAO5RVNNqcOmxwEJNS
JuKhKr40znd3bSaQlpr/9caiGj56BB6l23+x91zsW6TjP+GSl5/XdR10jmBRnZXHXdU9KoAqbesZ
9L6Adit6Y+REBMfzUybcUg46U3fcfr+mB15E0wl4Df+iXzNlPBVyvo2uxA3ei/QK9bBk9UhMz5XX
BLRpICj17oUQ44Yzd87r8WYo3MUXXFI3gkao+Pr7WkWsuHUv+oKzVry/feJ0zicsu2gQw7vu9YHd
9YcZ7+dR6S7LvP7R2ZmyGgtcDWXN7u3tGIAcEazuDpccQAuDF38kzKUztwv9XSjPxWqowmNkC1Jd
k0pNLXOl71GrjAyS3JSWWjaN4YbUeM71itLpxqWFol4mk/PV6XfFVq3OG+yTRV5iMVxDagOAN+Fc
uNfEd1dF0/ujZVMtvvpao3GemkxUyUnKEMnKpc9LRpLO+nd0qjP/OsAw0VlXuitJVAOqphHeIUHo
2iAMquCsV3S9ESWNxULwqisoRKyDnI7GCgqtA7n5/1pcnjsAsVt3/8ScF6KdT9bUmOukkM14NKJq
NXWwi8yCvnMJ8jrcRHTlf/0jxPvkcOGuCxzPsZj2rMJOZnV8+CKCuFUuO8IeEVmj7hrxHw0ZF+7t
e/dBq/i0R/sXv2FhossVBfpvigAyKl1Ulv/H6wEufmPKnmTsNV0K8D6nJn9QLAbid8P7Y9nkYcC7
vER5du6GGkVV7N4UHFZwXRojpZuSU7zowRc5B56tchss3t+/qYS+/jGgmb19Ho82IVfdF7/tlrx4
icjY0tGR8Tk1o2ojJLHtSd9xq7IhMrKgl7vdOcjWjT9yEGybGv1jXFI8GDK9weevfQ7cM4s2r2JO
THCVVaKqAa4pcFnF5QzqRYVyIvwfEot2ycN8Ms9rhQhrWq57J6vHXUN+edzni7hv8eOqGCsNPo2h
SWqv47Pc1ILTzc9DgEKzU8f1KNtRIIkX0SVSAb1iTk8w04m1t6EE0GptEXCwlv29AWGU1WrgjXjm
uCC2gU3FCIcT7x22NsSbR1lsXn9A89aN+kA4CY1+Qz5TpQ95HpUqpLVzesu1J9zuvI1K1GtTBq6o
s1GEP73t9FIClwm1e9Z09AxKmbpR8aXexCcWnJeXqqNODxJ4Ewe0lMhpKU7WTLUMwyBz+4Wv5W8z
opT2LvDKjvthAIwPjDOKpcxJbZ9endIBKaOZBOwJS+utm3K2y0sIJZSV4jnpmaxSwjdz4I84SNXJ
97OUpR6yGMhqgxiL5/6pwhux8I8KnvF42lxWob8tjLIWMoHxpfbIehg0uqcvp9sjc1jcGYawRczn
3Un2/dFSOuBP9QcQzb3TYFfl7deJSVjaQTy2deGv74RN1J0SWfhbxtpyBRYLRDMgOpMIFq7aQ1PS
UJfoDoX+v2ctsKhjdvdF1MqUyjlfEpAxsT/nBg8SxeKF4s2uAHXHBib+tvDo3UPforBGfGohMm8V
kUKeHLa4qCFsoxu6Aj/hI2nolyYHV3t79YRimOxPiCNOwr+2hZ9T/2D0pL0Sr4zc8pcA/hjJiDi8
tLvo3TN7WO3wrmdPruH8hsL/IAQLIzUxw5cF7ETPCB4zcaM+GjwgKM9N7fDI/cpIzmLnw++rkxkH
A+B2LyMt916233mPu3h9go5aHl0sxLRGfFSii+faGu14sLHSGcNqr0cp15eCRqm7hL1jdsu4X3ST
RPrdohSBNj+Av6Fk9mTt5VxRXknNdR2Ua7K6zDSgr8SzC5HYBA8QuxGivDG6eKkeVGIRppSEb4m/
Zza3bloKExxkAjLh0XxLGicRNuuWjHorWukFOP9xVrw8tAgndxdluukOrYvv6P6UQnqPzKaA6LKQ
hQoBEYF89/vEjwaKxaEVdd3z8vOPm8VrDqJ/0/Y0DqErxOy2BA9zNjLHw7Zhzzftk++IgYuw8Fy1
DCdSyAPsmgtRgbYMktu13HREdD6pPs0PV4n5S8t3EbkG7kWFNw2x9d1qJWmRh2Brt/mlBFNM9GRB
hKZJ4fvg0PDbKbKxyyOyFTdSEDWIPw1U4f0rITWaPys0uAY9P2eE7/FZg8VdOLbKwSi4wUMsAolj
8YWoY2tV+pcMfcgcKpcs00uFM/8UWc6dL1uBWCSUyOFDYnaEDcrClgqwyftF4VnIRbnAoo/SQXl4
vWpApWEHSGsd6num2sp5V6mYMOxAGa05nDW6eUiDqSPpaHiMS77Dodn8+v2urhttvPqziLm5wKCr
8SdvvGj9FamRDY/t09GlylsSysDPDqcKZsPTP9x2NW3XmYa1WIrII0Le3//PW9x0AZfTL8Aznntt
d1Y6Aws9HqRqNFUIbvGqEidStOOpflgWrJsTkHCf1fQAkmB9cKksYNeTFYQkIXYAR/vHRzcvb9st
YYLCQHs/nxV2i2nV/hepIXGnbyMvAwlTwuDUNY7skIa+t/L3xKmygaTaTw2+9yCkJ8CPIS/Ql4L1
u5CgYah6UT758yAFjZAoJLweUMn1cbtBhExzKK18cUHzkpuTzppZM20WaXWkfE4zy71oxZPtVMOJ
fBfMLnFUPJo65gkmj5KwxuIVW7MLfs5ni1gfglr92MEnuqCotMSSmi+S+NbEX/g1QM1MsNB3JsfS
84sfsSY8kqWCIm8OvJiW5Er+RqjkI/mKGy8mdcH7vxDy+t7b7qbqsiNwARsCqKDS4PLMmN6nqxKc
H75ABoCNOt/CvAR9D3SietScwm0RbbxXm8KmjNINwGsJo/dZ8bV+QH/jAvG11By8EPC5/agJE/B7
0JNE7Vb5Xr7ZIOFCFCdXDPZQdd3pTpdiWhJoa6TZZAPWebO9MUrKifw6QgGZ7vYUbpT35blv6Zeq
LiJQudED4RxD889qnjYigj9QX2YaXTKE9Wkq+xx7fuxbwCz3Dy9jR3LcBE5dBA+Cfb4GDHaYHliD
q4wwOjFUpObiQQ3IN09nukKTb16ybaB5TVbz800gp02xnagkl4/021YB/n4MRVlZLeI1TQ8EBLfm
INCbPXaTuayUvlxUcMT+b96gw8N99WglmUL1aFTxX6NsUEPzaRYSlGFnQRUu1tBDg8NtCI75bPwG
zZlGDV6ppXA+Nd1ZIpg1d4qx6Y9uZkRKSJDkaeu2DM1W00P+TH8JOOe2eHWvTfEUBiu1Or1VkVrf
guSYFI8C9NNlM90BFbN8dKydJBZV0MEISImK7P0Sc8BJinRcvM9gGmQAgoGYvBk90ZPzGfsvJT05
ztIfClnE2MszSXq1vzFz7BUYOWuvlz8gCkuVwNMdMdmuq9Z2Tjxf0SdH/GAJhtgxR/GZNT1+OD9a
83QeDPMduchj0SuJ0+TkY/Vqu+gi6+EsIj9fg8/VIk6ebqq7lvlG+iTWyTW0VIAJQ2GYMbFEkgaM
grsTQ4i6xoHJO9tyGglBarnZ3oVPUrGT1J3mm7NNuibzEpZRetEycsaEtxLeOjCP1U3YQWpIeGrP
Jxfja+uo/pc53qf9ALqRhQFMPyMiGR2f2pLHsDWqSgrY4iaw0E9rir94p2s2gphrunhEED5eBLZk
opsP7Zk9JjYsc+57L/6lf6M8J0Qeku31RNQe5cvExfVKj1T9YfLULSjUD3ALYrNEb6zUlX0PJVZo
B3iLzqebktfpXB6XC9WMAgYzV+S7UYpqvHBqglj4LlFlD49Pd6cFiMaMgKRU1RO/E4rHAZxFrDOw
7BO+hZqMLvXx/b13HAM3pBCdow36dQklfzzAX4h8vyJzfPvm4gzaFBGFtc8D+Ori9ODVzTDl7Mcb
cp3BqLoKWXhirBuYRUReLbtiHBGK88UzG0YByNoi7N3DLMGzL6SjGlfmo+rkZEaEGQB3TGmzsxQ/
IfJpySIzaRzBFHeAK8Vci6KT5Jg+sWhiC7LpWaqG7lKEECI00R5Rlm9yeOgQvyT4lB6jXvSCy2Mw
PAG0pCXApEaPuUgiV33pmJ4mod1S1f7wYIPpFbNo2/gmn7p8SxaEE1pHSNDwzAXaV5Gc+1La7/yH
aEFBEighjJkRvhWbUA1fHlXwRcBqtkZWqxkfHfusHlpVkXM7oIlViZmVDfS4YI+PBvIywJxzNZM0
sRN1JBTaKAxz1aG/8fdhebITxEgkmexSxYuMPs1aQpGzxy7Kd7PDE8OhlwOib3Pnn53cVETlKiuZ
6/hV09N2EBtB83cT16lgff5xp200bE3jxX5f9KEO1t6z3BkKMOzm57SKkV65ocbUzIrw8BrBqngR
xmpljk38HA3UTF+eJNrpmeAO05XSxp2fpZlO/VHKYxIi0jAZuPaksuNugp7Zi0sWx4GyvD7Xc2Z0
LW+pv+WEsFig/eKyoKMG7XFWn7BDpEs1j0Jod8yG/wy1Ng093W53GFjkfOJCwXAzBAVE1hYrKwup
jCkLf7FQo6EBghHglXwQcicicqe8TKxDXE9FvMZU/YZOmQzpZTsYPUVNS8e0cxin91fIHttBv42F
QidNP7sJT2mhzj7dTMyrVEaBNMgjS+x0Ujk9UYTXzHRlEwF8z/5+jJ866181uUdhvPMF1yaHaiRr
MywYnbTZGL6yfcGMd9yfnquSxhfNMKCI9gERVNaLYebz3wzqItV8ggUQRuqk/+nGB8AGGi5inDgf
fyBLCykrvyxikFZAc+76qgK7O+Am7kz1boguSRO4PoSFhrMbNt92rfM59HrzihvGSj2tNKKX3iro
8lgWGnrDN8ERWmZlu9ZvtZzPfjfUBFPRi20UrD+JZbutP4UK/eVHV35/AsTqO+pRWDNH/PphKryc
Xs18gJLnFf75oRc6f6BEGt7tysVfjlkefX+9r3G2TjtPeRakPpfj/45wUyMW+Bl4jzyzyhMhrhKV
iDw0lQQIa3fq9MRrOeR1SDpwZSuaZbwyCjjPB+rfioYLe6Ztbk5Rm3GZSJbEfBRPjjKxtP/+MUQK
/+Zg8CK3b02Gsod/pLyAkioef/i5bf0s5qkVZOW1xAw1lLMJUmWXE+HDDWFqPfRppqez1AOUemzu
u83i3yveMnOstenpkt44SJZ+9xK1r9KmhsOdxjFB5A2kN5zUpHQiJuMPuN35EkhpgtSad32/Dwtn
0LFrVBT+B5jL1+P+zMexC/GJlzBP0YMPojotL0nSPa1x2kGH4sCUAuqmPrFR25PoxDOUMHy73f/s
3dw/xeFUL0vXy6NPdNOkUnEI1s5gyIKkasoNoeKhs811hV0hbhjRrxddcmkm+yYNl70CHDOmLUCE
5iSMtcROyupmyRF8X861iLSgeVEOaCWSpdedXjnkQso8aplsGcYpF0pcaKb40NANnJmnY9zFEwVk
vSEAMsTuPirI47eKBbNh2mog/cd0WXYTR/Fc3WD5d45Y6U/7vlVGma1Vp8G/gToInsMhafYwpnEi
J2rLEHdj+6rs4/hI5f+MYiosNz0miiPoBB9/HN+AJp8b+xcjy2lAqInjjVgZmf+QNaYK4L9W9dok
yaCL2a1RmUExGQZJ/oE+OjqzP4u8UV6C0aOtfRMeOqUVHWRuYJ17w1N49T2f58jxSS5siJ66s9TG
/S5e3OUrsNlX/7bjT53nelv9Coo898fmV8fk0svTQhA8Tcwpi4D1Tboorys3+Xt7qqQY9cnDsyIC
ItU4cqqbISVXUgwSJ2UTQBbRzOnqhh/ZlMb7K7VCdb5cs9Xjp5OMwenp1zo2/mlUK/RckOh80TPG
jV5/torO1lOh0ihUq1wNd+DlNwwIXwx0A63F5vvu0bCAy55WbYracRGJyz7s5o9Iam+75VRa55OM
WWNyHpu2Shd17YpPISdPRW5SjDD+J3v5eEPOZ6rMvOc0jVwhrLGrfwfY+s0NCHmXZKbyfQli7C60
PnPdFj0TlIWuI0GFIJe2ABV1SCZA3JvpY2MMsG5PacqsNGEZkrk+szpoAbNs+SMQs7Su5ZMHk8os
JPH2DoFfXBIuTyZbw+v8SiMhi4bWGDFT7QI6lLT3vRyeqVN4VLl9VVZeyqhXJDC7840W3n1ic1dD
2pR3j5szWe3PU8nCrMMO/sEwj9QTBeKsQyYap14xTb1kFC/33DKcg+3wbu1KXdH73VdRJa0y/okq
f8X1oja3dymdy8im7XaJb0+tsJJi1xgiFOLHS/LKiU9oNDTzLgaJxfrEXEEHr2gihdCgJFa3qXiZ
hcuCVpmij4POw71fr7IhvXLqlA6ioKUPLBCbIRiqEjazVUxEiKm7J/ILYf0sNSPjE1aXQFegn+o4
+ZnFcSjY6s/E6dpAv2OyTSnKc0eGzAyvLuJ58mEwUdqlHjriMvCKkwljqVGryW8Jyl6YhC0rd/uy
+XKKjGGN4EBC4YCopuMP5XhpmbDUlPXedix0AdRTLX93XhpiGukN1RA2uXYrpY8dGflh0ks320xY
J4BEkZWBQjgVSUN08uDeEYwrcN783OgDMQ8/UKG+eo7cu1Fo6CUQU2iu27HOH54vtabEPFOppauK
d6C2oa7x8XFOAkQZPMkIGCufV+yWGtZ4DTwgqhlVUI/ul+8Atltm+RU2TRg4gq/28SItkKT8NQQN
6Azbl4xz98gk/yp/SWIgDnf3FeZMyjBF/oCuQnt5T0XqQjO/xjBxRqEAcSWtcCgTLqbLoRHaeCNM
TRGrVL3NNI4Oq2wHV6Vdtw8Ud3loTEUz0Jr0CD43ifPHOTb/n8dSvTzmi0yw+dKIQ/wk12GEYdif
2FFDyJZdXuza+t1sqUlxMwOOtH99OH6uNey6UhTbiJ4i0fU1/UqN3HVy44BeecnM7WSe9Tbu6oU+
v0sXVUPkveng8NEXGhLe1lAe+LtTcnrC8DZyAA05ZB9591AO8rgmzuCxzH/JQr/k65W6rHDb5v0u
QmyT9YthKnTsHvQg/OrBsP13TgSMR3/F9aMZuA6CcXsdk5bdUqH+K9jrDHQKbeLKTWYpqxyhHZ8A
LhM4O19NAF5E9LTDPyPn3hVrFn50/PCdd3DhpIVW4+pezZ9v2ELiBMdPq/wEdsRlfSjo0G20q+gF
3WtOuyQasZW5HHSmaEN0E1vmTvkmFIKwoUslM/eDSuNdHwc7sZcLwT0FwVTnui1frg48inf3WGkQ
Z+TkFLMMRmL9bHzCzGzzcluaqxmVfbQljfPyfrgX4V6AC8MR7A/qWqw5nZqYuHW8DNYfAvWHfqsV
VNAr9G4hhJVMq18ABOZqGEKV13y/18lAjNdTWGT/KZfJX5npxLTShXWaNzDB3+caV+4v3hNSJMl5
UNJmj8kDDeleD9qjXHq9d7tK4xA9KgjPfa6f/lqX22yLKafqF8/LPfiyGMe9QqZft07PQU9KQ0hZ
V00McqUz7AiL41rAzJ67Cybzh0vnPVWboMKLhbW2a7WJY9JyC1l2Y25c1jXSl5JNRHzd/zwoeZ3x
JgjEl/PAPP/ntMC2pmb1QGwjKSZEJezV0rupQwaghCm1EiI4fKcjPz4iq7imKrHoqbj3ZGuXwOL3
ids520MDtBCh7waONnqNEm3LedlwLWmpzPKC0gxL70JZbSa+ZqeLvni+h7MKN1BstquE+gNfwV39
oIp/fDaiHjyKdBbdJVU9TRvTsez63j9h7QRidIxzCFfOfWkcUN8Vv7z+/0VSjToY4GfacIpTm/PJ
ToNwEugiUdrJkTminRH0j8B5gFM507vuYR7mPIYBbqS6BL5QkkX/+c+JNVM8fyK5Nt3foHL6ZTMO
93gtmYrfs0uy8dGiWRts/OBZkEguh8PwwvVk3zpwL0qxHq8kxbSl05UziswN9S3WLSscLI6ToGin
CwZ1h5W3Jn7wnNhwYi2Z9cGwXkfuHImfg8+mEcJ5oMdAg9lQm65Nd0PJiK6MEdRG5hQ1L9zLH7HW
dYXoOuNKCG+2jBsD7ARkKIsmKWWimMWCeORDkUw0QmAnrtYa5hSXP62Lo46op+t5wFw6G9xi0c6Z
ygmtEQwR+0cu+zpZ4LjjeDiWf4iwGgoKDgtQwLysvEpzf+n9vNVzgESMMuVRx70L6n8NClBZsuK9
tH/icluQvGrfuC8gHPZoLwOoQHnuV4j6wReTiD4beUtupJDxMFgP92ngatSMhxYbU8VtjgMDOVgp
cFIO2C0BDAx4KOgGD+4vH9gFqY1XYo0d2z7xkL9oRZ75JhRnkXaJw3obekovUHH8JeWUT+X+UGyX
/bGAcfytaMaaY9YrXPxLsvHKh+NtfwHxl5jp6KerGbNDqzkRrMtoQMjnhV3AewwOWEjhbPYJbrga
dvmlhAsLBdi7o4AYv/phsGEBRtB78Q8DMCrRImux49W+EmCXuVKHaWd6pgK6EAQBUBkAhf84HqQ+
NIzkJwmYJeFR7pOZxbstGcCQ44qu5xWJwHxqV1m0ElDcET/5wnfKouU3RIMBRGA/IFdwtwgeKn35
FhSCYROT3bSa2+0cTXQpQMDytLuCqjKeFO7eD5hHnCPDDx5Kul2bX7SzEOlcjsJAd8IlBU6t6yZq
R2T3BAOrE8XjpLO1ClfNc25+0tvRUQjlje1RLUYzH3QJsY8LWsF5hRyo+N3jPfD3Vu/UzbI24+C5
i5mqnZW2b3bXfW5eV5mExCsrCCYbCe2JzpmMgRTKBr2GJk749s8dytcn+zEWGIWffnlkO25zUb6w
/shVYfMd/vbGV1lRp7sy7K/7jgyFAx7AqyALxEshFcxjYgeeWvFWn0VPlbUMu5lTuzFoq72ez/QN
UqPSvib/QLOmVxvPseAvBXBipRyKIlzKaJPMVOAJsh+Oo4YdXphF3iZDTDX7s4eIbxPL0mexWIAe
sdbIQSYihGLtQAV7wNwC9EMVXjFhcHpP2pHlFwl5hbTB5RriymsY6bGntlAxBNTYTWhlMFs0zipw
6Xi/hPP1/e1Q7id6ccvfHVxUAs57i1uyL7/9NgEsdI0wNOW0ijSvjntw+2NBEblMxK0rtXi4toxo
tzMaWfDFxTviPl+1HRS4cD18mhK7u+m8xpIgENkqkxbpuSSIkZeCgJ87KDDdN/cf6TLZce7xGHbh
gcOBpiPrReKl6EJtAt4QRf73zObnjbU4nseNlhaeFMIdF7dnPdftsxayYEcmnVGUsBHf2gJUROot
HtK/Zg6Lb+jpTZEPgD4+B6/ETeiN8SjpfpKPezrN6WR3vEym25IabojnZD6zC93/SjfpqOssyPLD
5wmptUfEs9twz162NTFcmpuybbyHZqIC6CKe7yTFLnOLXfoaz35Saorx7um9rMeYYdIdMr3WukBm
oLKQzRAChme/R8I3lZxtnXsqGnrT9wWkUIypBqj+q5xNKMgrZ4PkgjSpoV3EeTNRHP7Mg3fznXdL
X2MdGHsSmW+dAhk4naw0JEtT6WCKYTyrvXZhtfX2Kup5gB/28oQPZvS6ocDx4qNyQS52O09Lx7vt
AkYBHNQv/N94C5w4MjxkEgFddZeN5EiHWU0egfiY2FpBODU2jqOVFPbexZrPPgOUhIu8VIwRRuvw
1N1/AwFUEKMjdqZfVxvZ3X+HWcHDhQ5oJUQHdlWJQ6a0axMgmpkxPpgTHo525RmvN6yNjMxZRYlh
L5AtJ4DcCiB1piPy5qjHzVkspeT7jTaLjRFr2S3VRNOC28amFucsVUDMfwSg3dn9PF2RXfIUzrgz
WKjPOlXQt8MG06Ut8sDl58op7kW7YN6qiBVNftGkSE3A0u2mQUt9RPUey5OHrlWclYjNndRssZat
lrBIqm+qqmhqjUZ9fTI1az7+rP0Y5OFeHFBL6vLT0wNZmTM5Iqpe5hQpHxAnkOByRvuo5dcQgvbE
sN2TAGSf8Od4uvuPCSWmQwnj38UO0XC4j3+Se8A357lAjLQtpHKyMkOnYIrjiQKT4stkCP6ik7nH
11JFCUfe47rgSlx1s27O/SPFsgQbLu0hxyVWJD9PxPP/rL73WOLMd61ub/Pm/vj4muu6KsmDf3NI
xe1Cem7t3GApjoCxbChUeiv4zTIj6rDNh1WvMISDrCy3twpO6HVdDn2RjxjkI2DcSgo0Nt81u14e
mB9H2FEKdj+F8OVO1sphn3tElS39Bdhg0rvTug4GY+Byzyoa2zwpX7YUSmRpN7ZLNFR1+H9UehTO
RA/FEpyfGIUt6EIXZ6QuAWesoPRGq0SlIn86NqF6VItWiDwvfpX8C0r8x/EthpOmsuC8ehLA2bId
xfVvxVPi2nOwUlK8iQqfOtdwUcYxnO7mmehvyewmMJwtD+W+pN8PCP5dOzbEv2O0NKWX0Rwm0maa
XVJm3MPIsR94QEB1AwMll51RUaxoUuETO+1ApyIItESvgk1KjcrT7CU+mwuZ24NqRns7YZ6WKKHo
uKiQwME9UwqRiXVadkNbBOI68dvQjD7rm2sq4x6E9JtLdKYra/Wshdf2fweZ8mcBcM9eLNg3xlJm
rejsOpl2NZTeiPFf/fKoWh1ehz+GefToLyDCYaUABlIwElCZODwc1MxHXb9Z2Y4QvuloO9uSdfpn
MQEk0M1gkArIuxm32zmt7yMnrEX2L8hjInSXH0smhObKGhLXnpyZlQxVL3SnHhZ7boBIOUDCPXuD
ohNnyXMHyv23EnY8xN+vBXKWHZCDMgCTB8VorufHYt0BqOozlms4THH5MFs67qP+vPlSPuFFkK2H
APtW2FrDv7eP29x7kBGm/4HiMPplra4LIzFOt0AmCHdtxl3/6l8CTUHJRdhFqJIxf+Bhdff1ijyq
oJdj5U+vfsZmc/ow5qdjekVVlXr9uBCfG1R2wvsGD8j9/WEwsvz6IW4gI2F6Ir6G5yWQJinELRPT
I0KYMeo8koNQcj6y7hiD2kpsVL+E+/cGXz00UURs77qREkHcYAcrFRSai5soxAq+rmlB0BQgh57B
3lbDn3o+d46F/qUBZ3GZ3LCXhV+/h0hLBxVBwPW6Gm+xRJrXI3iN8SOBg/60qx1j8x7OZrqGaNph
8l6/GHih48mkYHj2uKTfUQNzt709zqZxm/MyL1OjvFrjnWvwXkrc50DYqDUg5kBa8R8UT9nBjwMx
2g9HY7XvW0ChBU01LzTSzUrjE/u6gap0OI2j4Ggs8aqFmxEeQuoKM7oooUBkj4weSQnXo/TSq/RI
07XS8xjrmh0e/soTK/jn3ce3/Klqf6iWhdLQgS6wSQ23/dntMcm5stivwBb5lAZDfgbqc7fVp18O
dQrJwu7iO8DujdPUqHJz7/od3kG8cUXh3ai3BLbtDvNdwMi/XkAXyd3xubN5UCFmC7PXBlxyVfeB
pClkxs7HHCFdSu5HFY0d4o7Yhcq6T56VWM/7z2vhqljaiwlhm6V13MfabEcVl3bR+37CifwBxcgq
5pHkCYrPI0oBa3UPjlADuj1tHhayspRTNVyAsuPaNbTtA4ctBW3LmAEBdcPVxo56TifEfzQi3zB3
DcGRf6bJnlANjkfA0yBHFqJodBk9FQPvy3Imw5EIX17XtFlI2UuGwqZEXhPMld+AhsjHAR/kSLYO
7TIM9KIP7p37cP8jsegObjS2cjLnFqdHm1nmT6vsTJP8s6XOkJQdJx4WUCdF5U6pOzFwEej2tF/A
2fjNfWqjPXq3X8hvfiYkr73U5yB9OX/MhBjZ8UBTaSPY157T30/ceAl3Z2Kskm3NB7B/eBX/zcBN
ZI3XqAaXM22ak0XaD2LBRGcY/4CVgti3254/eORQW0HNbcJew0ngbtWEgfTb2LYvugCYsanMbPZA
Ydu1nuHdWtC/JJemmiywjnrDknuMN4nBdfgdbTsioxC71KloKOuP+T77DFToFxRSwcIae2X1yrV2
A1Ar5yqptnDmaUcbAaFVwfsP8qr208HMbmHou3CFq4LTJHICXmYB2jLijIZcDAK2SdOZYnDmJ6/e
KE1CdZyVQZ7vEL47Gr+SUT17h4VxUc4QpCAR3ie70SmabDy5OmdkFdqqhikbBGMturYL8xgtbc9k
fBh8PRdBKYmjF7M6aaE8vIWgi7gk4ntCuAVqHNg18aSA56/0539bfSgmtF1JH/LTdROjTj/9sovr
nlp09P9WN2ZhcoV3oyqWJGSV3LC36xtlW+dHDPCD4So8lphl02P6lVj4qG6HTGC9nyoaoxbw++FA
zelmUvRGjHfqlGDkPJfZmyk04kFGJLid/6a2z0Pz/IkXju1Wg4Zwm+P4seWS1079FEe1uy+KarzS
9sgJGU2KqOKKzqpl5LwKI/UhcFVzqc7wMYYY4kDJR2GoqMvC3ujqDq9hvw5FVctEc2vo+BBJO8MZ
YpQgDIbkm3PBc9Cqlhg5Wdcs6yBs5l6Ug9kRd4tqPBKmti6zCNxFrolN0K5kYFhasEtfHFRc9Vh5
5AuoxsnJL7h1KIIU5cW1G389vyWyNI+ADu7QVcWPk2Hpw6frPEAqX3mbFKudUnwuUXW5EBSdni0U
axtG0fuShs3tr3lWwitHaCaDRr3OkbHuxjVW11srQ89KYlqyZoZvNeCG7f8uyOfoYgCGxHC37oAv
DtxYfAEXjRZwiOz4w6t/V8ezf4Ru43fVsIzqOxIDSUgwWOiGOCJAWinWWu99fbtDZRea2nSpkOKS
Ylj8kzc3rImBmJX7NhCej/OHwk8ToRzKIxgwWVwJxHirUCdb8ZOS9IPPPtsIpqEGU7p9nG43Wv1j
Gm1cRRTQh9RVe1CIljKS+X1TyaDVtVfEKh/ldQiOwe0dyGWo1G2lH8a0VmRdcX8Sj3W/gkA89U2+
WzgfSdATcvTZuqNs+JD4vGxSaAlyWxJScHE5Dfr1Kq/fBCE8qzbBYoUEN7drW7zjfpi/qe8YEbfF
m3+K6fsqZ7m6ghwaoOE7sxSgr2MQN/vHJtNgPKYOwQQtldEyDc1/ANGXP8lN16vK7DDQ02sCMmuf
9KCq2AqOojEJ2Db7OZjAgI05kZZjv3U8F9PSRylwYqWAwb3LqokXFqsMmfcBCbX41c3AaS/VhX+1
ansOXpI88NKTo0DBplSAQJ6sHexeWJkhlILnLnTk8jJu9Pvdd/EA8FkVv+kuLZ966dxxsvlR5zmM
LYaw2Tg1mGoMLkDkd2QFP9rqdctFPt2gNx7WWeXHyFxv9kwx3vCwK/cEo0Wwsw3HKrecqpL4kKIZ
AYK3MXTGEKtpDbc92O6vr8tpmu9thP7TmVB3ar2flUve/Bl8NeC15FX7lGM6ACHLg6BM0dz3bY28
PS5auZq9Ql8p0XbVRmOq48blm+yvm3Zf+ac1RFeh7rmr8eSo5kI94Jix2BguJGC7VBd5x7ZNCTcK
nYyvE8Owf6sE6u/pP4NAILzzX5dSjQUx6vBvVaM0L0bFvQReZavBHlI3UX7VuDteJw6+qH8Mvzmg
J8hqSai3lTqn23+IsyZSXkNdvRkOhc9YbzZouAdAciP87gO/BG8RQQ4Wet/0VHYsEy2vpulds6pX
M5C2lJuTJqlg9IngTcTV++rRhBfc7Y4vnagbYzjtm1mGLG40xtwCMeecc0/Ss8Y7EgBsJELqkLfP
KT3DqdJ8OCawsgs6Z+4VGvYNtaXi2D3KURBTVKfw2qVP8L0gpRioamnjpq5mfIwyLFO1MHQotxKu
80Vc3wG/BppvDOZCQ/IIPA3Fi0epRBNEWrUbnZ8lZyoKlL9Zdigu6AI8LcPHYAupobP+UlBrY+dl
SLTqNglfsnrZUHa3VhBU+TOp3O5rvT/5chmQ7FkqR5HpAsXu4TecJQRXh+7JiZlh7WJr3WSm5HGI
DuO1BPjMqHsIkxxIaOWN9ohdL7wQ/QB7Z5LN6kRbKyszqZILJCBzyDU74QwlJPAuxteKUMtOQPbi
0+BW/HqGlILaWuFrugd9mSkC+mA6G5DBFC33LjXBHY7F4/KG1SvDeJEU44Eoe0pV3UGPAQ3Gt5+d
FarbSvRt9WWUelB4TanMDwHPmq6zXCWspv5yJctGoGDDxpFW/bHOHXH/7mHoVoa1QdBmW0rQv+Hy
ao6telZc3/0s96S2SJAT7nG2Q64LYpVeM/9s0GjTm2ivpmAPlc7kyH0nsOQTD1AzlCwHO3kO48sB
RwWU1ktlLIObXhZtMTZwhhXcxoyluidbU1T4NGABu76AGqzYsio7XatMayi0SmCbK25nRHQR6NZh
oYtVUTy3MsV+5xu86+RGL/D+qDKFGIBrxG5vQXXkaUNc1KoeCqVfxG30TRGIu2QFF4x984S5BbNO
vUWjOQVFQVSKKkcnjyKbMq9WP3lUBBoYLc6M//5E7nuGiLkCorkJ/o0F7G8g6YP4LZ5H3qr58a/f
IL9vbZ1bt3lR0DO1gWrjGLjdz2u/O2MR+aMKt/JR95sxmSq6h7KsqE7pbz/0YAPgsyp+nkfmGAGR
DUHKjO/MUHMX5ejbSR/tusA/0/JMlSOStytuI6aiba8F6tBb9b4U0G9o2KaDSxppZOHnSzw2dUjB
y5ElYAwX1jyxGFBuC01XJfuJVAgFieSLJj/4nNhuFlazINDEkyb7N4w1Bl9f06zBnjVtzbm+W4rp
GzY/CbUJ3lgUd52nCxjG1jDfuPKISCJBsOrZLdovIjqzfyCaEjB0HkX0JlMo37tmDkdak/DxMnfs
0rN4W93b/jmTEzcaAVuT0LyIVKsJDVYOzHBhfHRN4vVa4V5K4ULMXzsUZrsVPH44CDvzQZBCYCkr
8u6XCesUu5nssJd2sGGxeCBSA2fZCybhN9RJSuHLG7RWvnnvu6efPo2C1XUQwh9lUNhAQnU5M9hp
CVn5yRjqHKKvwWI2/z+Th7vPIlTlogjv4MLom3/Vw+sk+fAZzU9+ZhgkTJ91Xw/9kZ5bLC0ZT/Te
hi8x7bv8MizGCNGOrs9Z+vp0TEiVir0x/0tO+/ewN4bmk+MFwX1j9/R4PQ9Tno9utW3oyumzCOiM
lsFFXBHEIXOA2IcljVrta83JuUKNTJyFN0BZgm2I8VbHGgreF3k+92B1u8m1m1ghP7WFdwz5fRwF
/NtgqFr7EIBjM5CBnlACmhjyGSdlDQNOoACrowq/AAYbPO4G5jKXB8+8aO1kxrzYNyxx2i7Hx3Eh
/P6OvrTrjDUeJGJuD7inV7N6bGQ+1g01d3mQvDNBtChnmEieZK01l1ot4hyCF/CNVHaF2/cDC0vd
oU630cWCiWm3dSLepsQ0HYgQOlOkvRq0dHQb9q/qjWFdkuH4zdr4sAu251mWXO/MSQL3yGnWzdUp
NldEdF3W+CcthEZuHl5R/+NtdVQdJPkQKPxteREa+Qj1XSU9OyDGYIP+1t6k68yZy/sE80lk64ph
Szj/aTsnOBZgUyzcUqR3O7sAaP0gEcesbIDoF6xEsg2nNxgyvRNVuzTfSTTi0p8FREX/Cu9OGURl
0AkuiPtALGUCrAMpzHu7vEvduxiwvMuvZgD6J+zmvgK0597IIAZ+yBfOuSIPxCHc4Ph4dHqMYo6f
/jP+rhE8q2N6dUyNwfOR374UYKuU3mUS765GaSMDU5unoXh8cMPQ9c54yKSGJYvrUdQoLQDkKS2u
koLoAQipZoujXz1xIllFOapoR4egBjWZhOITMgCLkrK6HtP1qwxcgUkflMXtqzU0wdYdq3fX2mue
JRJ/udHedLmIxC44NapOSzO2Any4JNnZ630HE/SSPFhvybpm0OE6kN1fyf4GOSZtpj0Y/CIKdixI
5UER5thYu2mlX2rho7UPttrbK1dnEiLDm/VT9ZbZGPsXe9mLq35RpvF702t0vaE1OZlvLV+eqAkF
OQfU1imYx22vmsgIawwvjvyGGE5sIziAy7nEvve+KiONZgEXburHSyIOU8+YLS3+Rhghlh+UHhYr
AoUKDCFJ/eQez5cIN3ZfBr8wIKV3EI4WJB614XMN4X7uWI29ayVLqd6j+Is6EhObyYOYqpU1neQF
qf08FEvO/vCUXXP4SdnMTz9D6mh+MEnR2KFCzL443TjHPMVzG9ztgFNG30KJpp/qw79IwOcGksoK
4NhxcGb9CEOyDeqdB0uNLN6EDBl9F3vQdmDnsU4AYfTsor38mVXRMfFifE3zksjcueW6BMuMiqQK
BBOprvNljDQuocVJx4P4klGi8yEG6/N4xRtALuBDnLq+oeT+H9PtedCVhA3/8h/B/pn1r3fxkr1k
GLxGvVS7A88vGofFYeNlSe2tfErLHIQ+7pvPY7NA1vboNDYN8TfZiz8Sfkn4KSk6RjV6lrAe+WRw
Y/Ol72TIIvrDx213ksvzg4vBrhBPsGDXe1VbKsMf7thnqK1HKd90BRW9YF1UNn+Pz1psOd+ijH+R
GKqxrkTkKRwu+Q7NglfMsagm3JJUr2B8qhvgwyantwecUbn2+gTtyTrZxqIGAWuB+dT+rPvYD3o3
KfL9MOzqs6kYUKhl7ghBjBXUxvJiWrr0X2ui4/WYHKvPI1o64JaL17/ZA1faFgqJB/jBNvksCnKC
yiuCq+c0TnMhQJtYWoDGpFjgn9bkam88YnyA/lAVCXPdE+bMulSCa8C1IJnUJIC6Q6D/LDpPT4Sy
SGN5HEK6qMkG7A4v36HRjPdxSOehEY6e2t3ZwPdwZe46KcVcM5iKtrWgKwsm2jfIdlfP8wOM0wrd
ZjL5valsODt5uwm+Z4Mf9NMDret1ngh/ZZBlHzqMZNQnlQyuPy75swJw8QG6Eoye6uOKIFXwNsBa
t4+qocrv29yl/lJ0Ffrb6u0VFxD+dvH5N4Sc29hkiisqmx4yCZ+/ozNr3/BcLkftR4NSpAkkF+ih
JECd2AWwiOqMfAA9ahNCXCzfjmjqWwL0BDOn5a8kWWEYTYCjNr4i/mSh/tSC2WntiNJaBvKMlzfM
Q4LmG+kXJ5FPocyR3rF29xCrLEBlNmJvD24Y5e47rUseMTXUe12/cc/DgRnAXQAKNAsCvkTleucO
Pl+N7LkZaY6+W/C9HwaoRl/bg4lQ+McDZbR6rh6uC6hIx8TxKeRBPDjl4hPc30ZqKqN+ThyvTpNi
1b33o0JLkq/BxKU+I8t+aINXFP0l+rPuixYW8nMJxXcD6I00LEByqqlPEfeJEXdqZwf+zEbBMf23
6lX0/CPNg/KgJdl1zfEYbbQjO4ORmuo9iNs9+gAF2S13W760WFr3aw1j9Ky2klpDLNXEBLk0Z08M
8Ts2dSMW0bivWh+VAAfPcv7CmnuK0fy4JH65SFd25anDt4mggRdXnTCaP0cZ4pIqEM35G+KHC0uO
Ib26lF59/doM1bXnjpKiEdaGDgwU4kC5xpDAC8MZchPDdHu1D/q46NKTim3HUQwn7h54Z9kc+37K
G2CsiBLGirzwUHMgAEHCpZceoQGF2eTElfygBPaxLrfJjGZouVqKDQi4U9y/2RpCRIZ6hMzasrT2
6wFh91baU/XkHFWq+HLPwzTVf0f+BIpbsDOI9T8q8tkkdBEARhcgYYevu5n+v/xVJfLYsiFZvuon
nUBwS+pXj7hLFprQCvaQmWEqfA2VzOhcaB30SwSstTlBk/JkUD4zfQm6bRHwaQIeDx9qVXh4XyLs
qQPbZ/eHQja5B7UvEo0Toij+NGyORiEpVfnxsxedO83ppC1wbmlR/2PndMDIblOXG4gWcIgqm35W
ujt+NydNQNTAxrsQV62C9VO1nSoHX5bUDI8rjvy2OXwQ0RDISwcfv7LhImqVFFTi7ed0mvZxIFt0
TKXd7nkzfF7dWlTHT/2I9SjIWg/w9cDUcgCFx8Ffg3QsrLs2A3QGOu6SBHgoFiO4CE8FRHraVpJx
sQt9zbFTJOvk3BiCpbArg81hgYiXt88KW3T0hhEvvkuD23u8QjQu9AiBgVGm2ycHh6jUeOyKmvWM
OxtT+Moosm/jKyvXHFXShHGOR0FYHg+RyVSlj7jvzqbZyhzE0+JZab/zJ3wHUXPukJCvJrBYXbQg
+6sBhwuqs+B8F6TL1loAOLSHXw0tNL7F2gCoOXSorrssy0G+NaqXvaS93XvH76xxyjJ4otdw06CS
g5FllKFLtOPQmwErBPByU/9GhZl1nCoWlxl6gsAmQi8+TB87JSddEQado4a96d3Ruyre+hD6O2zm
WAwzrnhmXWHczXr72en9hfa0YB04T7fUwTyIPpuRZo0aM/qzVpH/Q4Bx7EroN5GLQT/TarCJw7pR
aAfq38sybjT5QuynIh2EMUKSej43ppK3FJJ8lHh/aFnRwOnplOWLk/hmoX1nJuzd8l+2IuYGUd2c
8x6FVAGRzBC4LwSTKru/B7WgoWx71u3eSu5xfXLACjQCejq4mX91LFAtXVzidboDpocvnWOhjyA9
J7eM2/BvfsYC2EuF/bjqzpdIEbQhlov5vasKVO5gmiIZkBrEBKdKKoRfI86ObyADSHlh8F5B7HQ2
WOtqcUoe1kQgsCm53GUPz8S3ZB53TGkAErMWzfuYYFTGYB4LtlJfwZotq+8tsrP0qHyTWzPxWe0D
ZtqzO1SjJsLmmF9o1ejsvoERaPBU7sXJ8iiIFsbbevxP1ygY3bNV22ss0WPv5HL88Vqjh22x7o1a
TXgHwP/EPxlnAZ4sBDoxMsHw1142DhVmNU4o9P9VHRvRa2bKi3zMIj05EG7giKHL2m7yQVXR0GkR
dsdycqr1DGKWBOx7EhFpXA9ihXTheWZJwPx7crwZQhzrNRRDuIEpCAw7qmEpHDh3BqOLrFXn40E9
sQNYvQf/ej9Sx2CxkX4WhS9HcZrrVZ3cawbYUDDCa8rtTqNcLCAxSje+YhNJHUgLfqNQX0EbiG7r
dZ9TgOknb+rp5SXvib6/Msk45O008uUovG2QY5oEaL+yMZFEe1Z5iaYPCWDIjOTQMM8H0yHYk20c
lzHq6j9Cz+Bza2xrRwptqjdQNidExPO6W3CoOX6sI+fNB7ehPgg9iN0HLmsAfZMkpLSJpQEKBsU+
ZrGKrw+V+dzwqZMsAF0BTyKF+vLbi4WrvE2WQxvx1nR8f3YDDtFWzGUvLDYjB0Xm7qHLplNHfok2
U+JBi4daffBjUCTU2bMV8YcqlsdFUBptCNhMYRVetLqk7Je5Q60OxXQEOP9bV9T3vcV993HWQvHS
O7oybXMgSq5hJAdGcy3EuS0+4+jL1M03qRB8d5QUiay5Ega9f1W7W26THl9VfPZ3s++jaF81HtW5
4qcB7ogqNvZrY+ZsBCR+2bFIJkl60YPMsCBghjBXie1uRWRzOv+RhdUeHK21U+TZX6GgAtvOFNai
GPebGuYmeFoX1KAMShcQmUjaQH680WErFJ/aEc5mjLhUOdpTOdLSNR90i/V/vzCdAHOz4WqX88S0
PeUZ7OLB4wg1+GdiFeAQxKaONvkFM5sErqeIMhmQjs6niFpF4DiqwtWS+Ne/FghgM2e3cE2CYZfo
8TGDFmtLqDfDemhr8clTYLh7nQ0g20y94ndb+8bKPeTlZrCKc8tMupICC1zmIOpgrmDfab8fh1gp
mYE6hNegyEUnZwmF3CKAnQ5KF2vbvYi//UfDmj8xmSjs0FTFKt3k3/eDA7zQ3a/9k24jxL8TsvKY
pl4rSjjBaNaw+NMPcmNYQ6e3UjZpNROsQltBo/YIEwfUpYLy9j50PilstUdBgOPVBGjcQbVMhPlY
W2JBb2hF4cw8BTovQSL9zpPM1mJSAE1kxbLMBvbwlgMf2OohhBHWszBUi4/3IfUDb/o5kJHlOEJF
hlLtJyvxiopq0wIZtkZX84NRqcR7EcEkSMN2wBbWOSxkEU1nwnxYWqOvH1tad33cia0TtJNfAiWo
PL17I9SOeCB1+q0T8Y5S6uTl42uBoFFWjwTeYfnJa3d/omHErGDY+MUII0hhFg25wz8s8/93wnTY
xV67+Hj7Zdh7HRuWuN7X4yLRJlReUcMPkndxFGZcTjS4klYmLrrZ0mK3do604xtxWfX2aZHqDgDn
1C4SwWyiu85nGg80UWgV6Oda+Hja6yb59S5ZGh4eu9+MXZR1/MeNd0MjcPsPajvyUfOXZwLidO6Z
29JtfWvHK6Gbr5ETBZ4QiMALBfiJRrqvI7PGoP5qQYflsdqUSdlDeR3RiQMT4SfUFffmczQ6/nLP
y6g69spA6mfswmZk5e3CmniNukctjbawPSclgMXWjmWCM30kzEuysh3kY2tQC/8fVnKOBzmzNLag
jywmPGNeM7bpErdObOxrpG25Z6KZn4YGKixinHhuBx4RsKrVYfXXaZtwJcmCf8QYqQoVHeUp7buD
QTa+pT25HLRsigOgNVJWuSQzHFzl7f20FYYBS27Qt2y4TZiprPwCgWWbB8j54dyi8s/hNul23v2o
QY6kIMpXSNLBkaznpv9O5olYIVHBGC4q7SOIj3Xo99TNF4P1Hm7wRdbm+MQlAeJelkrc5KJK6Eg4
2bwCxysjhwD34a5nN1Eji2fauoBcB5z7y7LCfh2vrOvNDnukHQ4Fe0d+Ohb7/awMTnnndICEJvYE
6BBjWBsVVzotjpNhRJh/yWitW6WbUq0CfJZEVPRABoFn7tqWwVJa3ue5zzK6hm/nk3/2zp5IcAfa
03HikOOSS/Ic12VrdgI56t7hsNMHuDi5WVncpPMqm18tvHJrv6ynGYOMs7swS0CkfZDwb9W0dXIv
Z+L5oY23T1MYdpxaDT7VoRoGfwIHwkJdtnyKNQ76TjqkPp50Bf3ZrzhKkPE5R0NbeP6A15xCgcTr
u3nL2+wuB/SfqvkkW0/yHUZx+NlyGrlXr8z+W7etULpJ1z1xT4z14kMZ02tucn9XolthQznIq9Ww
Di+N0XrRUmkC95A8jQdBUqURVyV/en97I/IPE7oe3PM7FYYf7YlSuy7DIXIVHZDsNA0JJqCVDDKn
A6xKs7AnKGo2sKSwRsVLPRsLNZpRvNzMbn+vQ2W7UI4BxLf6gOsJ86DQx0NU31uSwmhhTui/DPRC
rE4TLm4yWLBZlXcF7LvYEfO6bsj/0heUKZ431GusPrH66vRGRcltgL9Jle4R1BJWjJVV5H5W6MKy
yF6cJALwb3g7/WEwsPtcdU1rrmR6jaMMdNt1MWyC8hbwy8ttaTubmQkQBGa2DCxPakY105Eu/9lw
EhBlKRVmoEus4+y/0m7pcGblSZ1dnzH5KpO1MYFJnHEVEq5TLSSSB6WmTY6pJdV9RMwkddoY1lNC
II4TtAbWITipLEq+1DMj7oZvyc9v3oYz4RWLs/27GgFFqK5k6efoCQmOH/QuDrvlnrbVSYw1fZuk
I6bIsOWXIbV2eiiszLDce2XTdHqL9kLoQvXGnorwRW6mAA8Qte/Efk274o1hY+/uV3UBRdDrg3p6
rCUWzySNVSSBmu6KuRdpr0LQ/S1TsnUUVvdBeZOL/2xn93nNABibDekdEbPZslh0A9MIXlX4hVT4
+8jXmpXHwrWEw9m6l/qIOKNC8XPgkyuWt+osYuggMFVvzpqymw8qrlGnlB8Nfue/F6Ng+g28Kz+F
57yMN8/kw5dAjMjSGl5FtZ5d6LhvxKrKiVg8Y34oAKxiPaTCEulDWQ0e7+Tc/7Up793jl5xy6fbX
bf29vxVLiuxd0/CnHNtk/RzXzEyh6fmKXUegr0XDEAycQ8wBh8CP/3DP3KVF+yuNLLH9SnkA4HKV
hjToJKHGYJZTBX4hOL/49yul8O4kLRniHDpbTpZb2Tu1hL4C4PWuTyxcFD9+mJubn5CYOQS9nQoC
VR9XJBCi57Op9x7vKyQ/NpD0tBw4+A/q/VPJhszURuYwzYKQR6Oa3eCTgNle2Y3qnbklsbYIhctH
eAlki78UqrSlLcg1cufalOuGTc/s4nnC1PopCCyi/ZFw8pm5h6DEvfCs7RsXfNeyouohvoPZD4qF
/BrFHJUsDOhOBH+6LCzEeuLcIJqwZHp9ntiAzqGLGSwhn1g4F0k3PQmx+NKWWD+re0Cy85B/rW19
AWJfSCOiWTR2XAbhvpgCTER1ydAC+M9/HngtvseWS1qNEhj0wn08WN7njdAWbJDcU82vfBfskNHz
6r1XM5y+kg6kiOx+2YSPFRNvuZHR94G9g+RJ9ubGG5ESIKc3OYb3+OHHTWDlTkewe0Rb4sNh+EhN
vCuEt8CeXyKoyw6IgvBJGCXf6LLuA/4/gfO76Q5IW3yd7nJlltSWjbEs4Cz3FWKkJr83HudYkjvu
UrFPxnIdicUDf7shWWdVKHEtMFXoi0e6zSq+izZPlhv9xWw2WVYyupwhsOQX+GjgfWHbQVOiEqCq
dyHOoOOQ1t0S7d6Oib6xwrLjU9mMjtnTk4f0o1tAwgnnw3NbCN2pST7jQyD/DIST8u3a2H3Ws1B+
15lIVq98HT8M+nJGpai3pKdSAuvbS0X4nWpQ3/Sp9LIH2S2rBAUu4umty/oivbE9UG0wZd/AGNLA
rfq1zmqmBsFTXTLIRRajPHNlm9TZmGDcZC0XX60+2+4rgLA9wC8FBtW36EzwGQ50U1kwhlzpJzbV
R3omHHIaOU9+NUo+2R6v4h4xQ9cZTCnxidfVBTH3AoJPyYyL2pRrDnEOrZCLkUgpIs9Bm7TpbtgV
ZQY4w57KRQ/mEsmZg9l0+x6Gv3HSx558hBO0ooosbiB2MBEAdoizm9WZiMlt5CAyw5AAe0k3TeXc
ZIepw8iIgevHPFNsN8josu9vs4qu8G2BdNORiOAgcJGa/QmVxigdnn1K+rNKRYCcbdjdA01IYpzs
SCv+LiG3VL3hnQj8KjihB/LDEGtUZPUZXluMk97GvZn3VSnIAeCdeQDkZ8CUqdG9Hvk6/d0amdeM
ilNlGFUdnm7b7l23v/p942mEhNONcqWscXKgnb8MYxwbdW04w4g9k3f9l5e5CPhlLCJ4JQlj0Zdi
W6FUSlnXD3B+xRS5Bl+D/8P/jTKYSIgHolqjK+8+N/tFRAF+K5euTVxFV6hi0Gg9p2LVeRZifEAq
TwqRpJk+mdyR2udcReh/Zkn1wN43pCFheK9XMS6h4j+9WS7pLUvrt5yISf8h45CtbW2JZyoy+it3
CMIh8/EMJ/gsc8zbv8b/eN5aMnvyggl9Ng6pLn51bI+QMXu2lW6vDFDUJT7t484wsK5W8Z1ineO/
zpRP4CHjXkXQcZ5klp2XmdKegdCtkh5uvXmdzkLktBWxg231LVij/K+Fqke09AQblz1gYFVgMEqS
PawvST437mWql1kwXGPr0ko8mclzMPvWvqeORDmr/Z6O9IssFw7mCzxFyYXtrIoXNfymx0CPhvAr
cJBKBvOQmf9eCrpgTZ5O4hvC/QWzk33ao6Yj9pJ/sZMHUvr25oIuWp4wLRuvSMS17dgGzV0Swf2f
hRFF8XbNftcI72863Au3vBRVFxiApWc5KQmSf8elYKB4iGXYJ0lu/flB1VBup4o7YDpju/H2PD+D
nkpwZChBC4JL+HHCb8xtGI7Tn0ZOjnSNHxXv8IqCUwr/ck1bL9V7ecvRDPqOW0U4VmypjTnxS2jn
ABHrnCw8G9AZhtwtP0p+k+CEmd/wLP5aFHvh5gqqKah0W0Jy8T0TNBKdvSdYYZdiHkR9B4zlqnz3
fBROhQT3p8VPu1/2PlJkfey6cOYBJ8ob4xj+leaJwq3a4lFYsxH2ZysQaL1G/WjWaQNULGChgYsg
gqIbp4HkR0+wyjVkYaFwyYN2xrmX9m3OkcSkL0gaUKZgX8a4KvInQm444ajL3ddOLXLfo+cSKN3v
8KRByZiCKWxJIH3E4iNbF2aF70lp/S5YoDc9DUa6ebhY0cQqPk1TQQCiqZwoOoeRn0TVU0XYY2wh
ZX/vgonTFGSoJmqdyFLVXRX1YXyBktZEqkqiKkdnP/bJR6TYrko5fKl8MEWU9kNioVgSJK+EE/py
NVqCvgdghBOK9JEXOw/u3FVgLxNoN/xDcG/1dKoSDK/ynhMhj2kIHigwfd1EQmndpNvISKYluUMA
ojoh7Qgp+D4vi2zJeLQRMGqhleC9pWlIHW7sNXl26QWw+tOp4akbptAUZAbLhhEirk0WFjpgMjzD
SVV9il6djq0CIaeD8ksSxsq0L+FormvBR/zHqWpVwRcL8LT8QH8jpHsqIHBf0uVAeINHbhfrCUgd
qYu0DxxrjC3i+pk/ASeosWFTICCnSXMwmD3gX3y9ScvGBzJ5HiDDmsWpKpCeNreXFMtgg8TBlsfA
5bb/+hIY19d7sCzXedCg0cdCLj3hjGfiEAvl7SKhdOYLU+ByP3xLPlW9pwqb8gY4dLHSHdKpxtWh
cIvB/9AGVMbeA/2MTgV8BP2iod4nyd1LJsvkPj7nK48DctSXK8xwJzXZi2admWtOP9oA54WMA823
VbC5rmHsxcYiktRonfyNTmRHzOhWjRhPulwf3U2n+rR9TV41Av7LaQEv93NbiFUmzD0zdavOOCjI
nV/zwP63o8ewOhMjigOru8+jF1MsfCVM/oyQUiFuYjHUO641A2O2TQIQuoJFL22YMdgLbt6ktw2B
Ui1NUg9ecf1W2tPKxyJT4CGi2qgTpoDOaik+qPOU3J8RTYWBMhAbKhpR3VNhebyd9QLrTeL6gima
qD96Zq5Tk+Ug0zHBzspoxyU/UpViHAUXu21Q5jXqmIY68Lm6stiXNia/2H2T9i0Od9WuAVI4Prxq
nCK91q3i3J4FkoLU6PeuAd/g3f963WLT1pFB/yWc+kUi3vTbHY0PkUnNkqeiCK9qdKyKPQVF4YqH
fKGC6qgiz7VttOsXNznLUqCZfG+668f7DadGPgyFfR2Zu/MlpDQVy/FUItx2TlmmjrM2wCRHHX2e
7lIgmdDUIt/LDxzcTokI+g7NDSMzmhoQccUD46eYRXdTNi6Tmr4UokhihmK7p9cQDGOraBhz2xCw
txkDjqW8YAa5qjXDmaxxYd0+Aqoaba97Bg0QmUYCMlkPFnl4DrRWZbyAqQLqTn55mhpWSc9EQai7
W0wppuQ5EMx8iOuVRNSiUqidAqjLFhwGjObojKsqL0LM6xvpoLLQS8KqSVHaleC8jQH5hPx9HljG
uLFCrrwA5V2dqbp4P+wxtNxMusPa63NYrUeT6Gf0/vu4R+kc7k7W/hG9D4LXmgxyoj9VQRIUD6Ai
NU2fVtijm+REYxcjFTfX5S8+p7plpvtH+PoyGJ8A8iYxvO3Tz83p52ORtpxqNQ/nU9MI6bQwct2Q
QLI/nzB2HiwxKm2jrjrc+1eFN9tRn1EcfHna2BpnaIUKjTAJh2irKAoJWc+aRVgxyAxRlEqH5GEH
6C3zbQSsaLU6zL8zRfgY+wkFESur8OJfqsR7wqeDCxCyEpYcZgD4lqQmTFk/8iCpMAwZ0ZJJDaiG
6//bg7/IQIXOQWih+E/3nVEFW/RkdtUeB+ejaopxOVvPvvclWv5LtOIvZCOEBxL8R3mmq+dPcKMD
xqmju53egHQAjIQJa8g2T5L5HKQ8vu4YSb5r/9gpxozONeb7cDGI6E0eIaZwmxsCezblZqa+YIDS
ZZIyYwFVNa6ft3bO5jCaq27xUQGvVtcx7he4dz/NhBA6GKkNRR10IH8g+Xe+dZ/FkPzRhkyqjuAB
RGua24fWfPk8QfoFz+AGksSM/u2d49oe82gghJax1sU9emIPXVRoMVddpHfT9TsOH//eqVpXxU9L
ujPD1spUCjfuJ/2MaxQ2YxGMzesTRJrq5u/3hWh6feVc/53Izr/Fhuf44/WTwrfhTTVTHRn/W2mb
qEBk0nrhZkMjUoEhvL+KXYTk3dEerPE2Qx8jGHbztOc6B11+wJ+CvXLiJfT+Ec3FTuFOibQxL+vT
ZwTZounXmu3RoM5hZPqXtwSmtwijC60yDVJ0MDVh+5lJl43hyHIIOCqxI4RI7G3TzZK8wLOkJL03
oiGU+L9/Q40M6lTrMdUHFlrKdsV8zXBtYDhSHoxT3frRbFVgz/G1r2UHEON32GYn0g7pt08+FHxT
GT+szMwBap84UazjTuYRHM/DNjnU8hmX8LvBh+oA0az28a8OKya8XGIO1aGfm7I4UpPtBSakDZ2w
PiRreIwo63UqhEf/lZep1/tqW58piRozepXkii9hOswzsVYNAyMjZ9IMgZB5ab+7EmqVFx03UvxA
pGDH1S4mO1GlX2yQph7LQbboBhpx7EUELXmle3WYtx7D1Oyxmhu6EKH074azTp83S/iVb0jXFgp6
PD/t/r0jbi/BfT9OpTZDunSPMXiuw+ipwBnqDSWyfuxLsrjPpp0l99yd7m3mEHFnEMbJoYBesffX
63gyGHyeQl2LBd4OLBOWjsch3v6TgmBetPXVHdR7vBcXmx5MvivaFWtLP/6rjEuPg432Toq56zB5
1C+SUTYwqEsWdiNJ7ZvgIwDSrKJGNsSSbaM+0NYTl5o9HKKc3VBiVT9yj+wWp7FE2NODONSYYpTA
to68Q6vYl6WO3yCD0nb/MBPoC3hZZvqfj77ZYDUwJUqnVijknMEJD5gchqZCr5ZHKOR3aG9NSD5F
jnSfQAe3984w/BZ8pQb1AAoL8TFP6rMMFrD9JBcFcgvTcACwCsJM8L1MQFo/7XnZ605vCI8kY5jM
LtpTDBDuxDtsLxjE5PwfPApLdrzyhQFkbDOVdVmU7+F0e2/N+F4EhA2l3GlrXpY/kuyQTjH7f7QC
ADJvoX/S1Y6gLZ9hLwgJcD/+c/sCgggs3OwrdGS0p3a4LTdZt1ajGHhOiXblb+kalYGlbsnIHP+p
tFPi4BWNEvcGf4fAO2Xv1euB+OgqU0vWfgAZm7RLu8inadZ1X4TRw13VaiT7jMQeiRa3gE5qh4Yt
4VY5BIVpK/s6KqU58nvIuBQnUKSF575g+7SFGWS+AGE+sNuMApHsPNRF04qfRIaU0lDv0zbwJgph
pP79kWGfRBlcrx2f5ccEgzd26QRPcNpz0Sj+yoWFFnHPIwRpckvsDtuoDaxl2WJXPx8KzMGLGNnI
wuHLi/xtFi3DSyJFWQ17s6b87wzFVpYdYq9xrNpVbzpSNoKrBE1zS9Od/LL7yuJs/e/dqDZhGZPW
kaCNJmseRVjA2svhFObTn9Bvm1d/IuDhXqSLkniPBa2TEl9YOvpIwhso76eXPVcE7GuqNmRfHyOo
mht8q8MqNHB+hsstsce7IpTJpIl7LK91NJCbUvxmA21w3xVLkGrlrQilshgYUn/XRKuF5pAUsw1S
hYrl0Grx0Q5ozLHu3nqeA3D5Ai5xYW7cmKUzib4PQhAbO0C0zS0TZ33RJ0rDM1pa3/POodYkeDJV
Tjxs8RKz9ozFWG/eFfwmhvw4hZUozdBqvs/sIQQoa9kK4djNR+LGyl8mPHH2CEjs81OnkupQKm+r
4lvWyD0RDkcRKgXfREreC/ZayAGyxYdcnNzhFqguMQJ7ZhD5l9iTnLd6qrELu/3e2Af3q2+32mbm
ovYVSMCFAog1GWn05VqT/pTpgFU4E0kmShNUUp7dNwIkwX0dxmqR6E7FlmRH1uH9go2a2Kdo5ejM
B56VAiG2TjC+Y4wTtdsfpmeW+8rZT7Ts9FMsOP0o15eVTpQZZpMKQ26w5VhPGQHm033Tft3rG2Rh
xjFmgyJGqfv9akIj1IMFBOKbVnzul5RnfqZnkgynnZLVaMmKzuarno9pFKRCAAcI4+V7JlS/AWEJ
KKtjotLyrZJFdwhVOUf/hx8wRSjhPtYGRHhqhfgR0cPXNvCkLqtp9nZso6k94PSjmNJw3N3tFJDr
5PZMqfN+wiu5eZzqCQ7Kc43qamBsQSfJVBaiAXFo+qYp1A6ILQcx7heK/vCGnUseu7W9W8JyPrt+
ATBWC6FR35pL+vff9vSBwDH07ZkOuqWtNcLqlM5SpXLQulE6eIskN6AldNCA8+LcRkZIRq3QcP+6
7van87GdYtJb3LVStrMtGDohYJdXz3E9Z9HzHt9tljI7Gc2j76dg1I8aplJcA6Vjs9aKyQta2O/q
Zh+gsKvUW+6ouny0I0qHR9v4rQJ5N+tveWde9tI5UIPaCHZhRWa/EYwXkbWV3BYT1DivaSQjIQ1O
M4Z4LSsQ6LAGVY3ayMGBeY8OnlH51YMXOZWhsGrR5H7iHdB58HGev2kDrNNZkktveewHWl3bWa7S
/DK3ta53cK2FYSh/OBclTGgqJ5UNGQ8rjXDufy4USM+OIuR5E+keDjNUsrfcm1ofi06bCheJjheW
27eEPdfFqP5e/Sq2AgK4aYVW2B9JwrHivy6r0cTaYGAk+Pk2q001se8NFpwNeM3nyuiPxRiAawXc
l1cFd2xWjLbRSAegn+9DIIk3v9+/NDJwDwfBeBosmHwkRTFgCuQAG+67g/W8CW2XEmW+gNNQzzPH
7HMdMmXEtMTvNQC+YcGca4TVxcdRc9WsIXcA6PrHDqotXhDS/4PAoXKs/66QXfkf1uR/KPSj67HF
xzLjRSzboaL0EKGdPnBwihml9+3H/uXy4v022NuFiS0e2OdL/AAuloPFhIibvFRkwidd0VKxMF8y
obEKnAkZC3cfXeQKPL6pBOpp65vBxi4PJ8PpwmJw/LqBT8ocElOBFpvwfpRU9DAg9ofUbEvthK2B
19IRJGF1mv8p+W2eiizgVh/M1coDCL8GG8Nt1JPC6j48pgrp/1dXZ5g+fxAF+pAcEBnPg266Zv4z
pYBasN+ujKCV8aqH6P45CSBYsoti156M+ly44FHzUT0nNq+gOFofzyVs1ZVsIA7Qu0F6eNY3IzBy
nFvZ34zSMpRm3nvf+FPXTzObMrX9A8hwmT+Pv0V7A9D1OIMyW5IrCOZFfb5af0kwc2Lm+JJq5+i/
eCJygm/lEt+VfRMNdTQ8dN43s7faoKtU5zWSPxBmbb9/o849jhyJ+xkEUkU4iWpQlnfqhBBKncHo
2Y2R4dpOlgDfoFY0QkKc5xcIeLEUOt42eHBrk+EpmlpE3vRYaddDvmNxkJ+1rnul6Zmt5F0UcgTl
ivZiKKUZCSYZ+mulwzS0S0rXkDLizuKNQDvtiQY2LUqwKH6kws2VLAhv9uFzPAuzREFBnl46yvBL
GzgmiXFnJ2K7xO6hfCr37vy8wC1qVtaUHqgeFUiK6kq05mP0A1aZmTMjiUG6eAhwi3fYC7ELykQd
p+5Acf3RBFe42BTpc20kTS6mqy9UKSITdqnCL86Y4/x2ZQXEVSqgrayUMkNhU5F6XVi55X6HagUS
+bpei201mfpa9jdChW4lw72yuQVS+iX1NSYfLEOHzg8xkaw6RfFtTPRl41aHOWXQcmnpzBOUx9g4
t1SK48CzJ9e/eNGV/WWwIfuPOSkiJ+AibcCCKGuVNN+BaeMTNWvTK7Cuw258d88ZaEzf1Hto2xRB
TWA9PLbOkqz2jiFKew9V9tkZgBCqJYrkHTPAVDY80u4LkmrVAcSphMPC3mMpUD+zXzxjGEXBFtPB
rFie8ahDVHnd/Lv4EDmby4hX0VPgPCtw33NlHUq67x7FK9bRxc7GUk04mPHV+wUbQOpV7CpYiJH5
Ey2DllDiPiaEyKukwydoCLZ35PgKToF8Q3V6nJ8vVoGyFpCQEzhp1hiVdF1P02oOmoiVE/FVyytF
nXU6MtfGjZpJhZOH+cCejD5XkXE6xbjdSw38XTNaEtfv9RGABIAN66nM4R12xl+pukwemi3XREdG
m64GMuhxI2LiJg+bNnnS/JTh0Oq8vubL9RDvh5s2h2LmRBJJypp/Crv8N4qLpPHiavrsITst5PTN
tggZxVG5dVD5QFpcgRYdMNcpsLzx45Bq0i4poRmFpZC5r1pYfnviOVKGfaFxUzVa2JqrDch529Np
sPwvyBPT7/vHe+6UGksAPi2/g9SGmaRHKAN3zFCmm4GiLeAvYR2hn4wXUu4Tkrl/sLw1Kl31T+/Q
csrUb93ll7yON8AFI5CYDnfnc0ycmen1y6CX3iWKMgZB52/ZwgFNlVEXvbhAJlDs1n9gSDEMQicd
RLPv0Q3E5P/M3wHIjRKKyqmMqbIuPchsYOo/69n9LoZjVF7ccTpeYkIoA2fm0y6w0bWmC6frwEoI
oPFTz7B6l+Md4cXiFWWRUi+vkxY3bSvEPLlH+HP2LCYkbynRppK0rHZla7x1/h2XU1+mjwsxami8
JgJXbaYB2uYqKW4npo6czS70Ck6NTcJFDM2g+Uat2uUNctGOhuYUKBuKh74wWnaRrFujaQCiTRqm
plkc2IY6DnrdXwoVqq7DEuYIA4UBOMFQ8oQcJu+EyPullKtM1RBjehUXPDJ3/xSxlBlYWd/f1beK
L9v2VdTPLqM/AARB6tnB7ehcwPhF61Ovjacz3T+EXeqMj4c7+wzy/AIEm2p+mMEVzwS/NMXGg+CG
k73oQ9f/XiN+HOi2lNN18dZQ5x/HPlHEnWRX5wNenVwdlDhQMrbWPTwdFS/snuIpOWM3aZPSoP2D
CwN2w40Gdb2plLkbvzHQOUPxw7wer5UVGJgDqzg3FmF6xGBXlUvo4O7SCI8SQtFn8HStAOvAW21h
uCxIVt2A7L9y9NJ7L0dbog6ogvlklaTFLUKNWekqDylYJbUHCooDasL6XnKpG3hWUKW4YW7uabqG
wxlpwMTbm90bfyYGNykhssu0+o7XP5x43nJXSQcmPkB2s/2BSOKXbK7tURgKxCGcy1J3+cYz17t7
cnMJmSiWXFPLgHlkRv501CO7z8EW6A2zhJWQI/OYXwST+Q0Lyma5KtEK+dj81wU9Mm5KUyjfdZbi
ELTqROzWhlnkejXhhnWqI/7eDg6EE8Ddg6pVRWAX1n8APf2taUtbXmQrcw1VwcjZUhmWrNIPKH3M
Sxa07u6EtvmXRjEZtK3hOc8YbJzs0K5f2GuhugySiQJkIm1mdGXqxmLqu5sIETaGu9t/lW1nvi3b
6cE7aZirgvyIaQdynMonkCqZOINQvPbamuJ4boP4gJRdhy/R4pRt4CJ0kWMPDsNPYbHZ6TBxsnI1
edRbAj9ASBvMkWb/PgCcTSzpFh3E1Qo/Stl0VHZIwYWJ7T/ZMPG4lcoZSrPQ8+Er2nB7MAPEbDHs
DTDfAPCcAl2BnRI8M6BoKEvmSNN2/JGbodBdXPwtF3Gkr4G9kaRFu/CRCVIW9UoKSRQzcwzjY7v3
xNKKLrDLtqoM+zE/mv7p7ml0TQ58myBMfEKXMNl5843A+ENSjMMomIrsDNLilg975uTf5GePj1Cc
hx5C1zbVOp8/emgHfTdpeRJekUHid5bfcUZhCkHaK7R5r7fo5Xxh4qCf161hc4/DxccfVZhCCPLa
Ww1wxEj8PjrO05n8hiltNOBrfzrNbYoUZLuAsOEuZKV5lRFog7Yw53JV3yNoNpuJk1kQzLcwzXRQ
TPipT413vHOJqGchjf+SFAqav4XtCBxoNDgnXkqjWGR3WiBoznn6gHRZYqMVg4qgJPXLLPc3uKkq
jA1Pka2U0+3H9QM92z4LLo/pRVLj2w68n0dyM2d5+DBNqLxAK04dbmFMX1oIqqcF4l8p0y91b7Jt
0FzWhAd41VGDAxXYoB1W9SMsm1rwRi+sGbhgardL36cih1Ig31axOHpK5FHxiYIdQ6G+aUfm2u9k
QcVoHR/GHoLGtimolqYrJm/jeneHQkjOeglVEbRa7BSP6TFLHfHtGyFxMe//W5vWy68/hsJ/gqem
TiuGjEbN5pCWwhCfjZlPapqPr1XnKSYVbZ+AxUeMV16kMOYPJQAl9HsiPB8HWrzdAfzqgTAwakAv
Obc0iT+hTyyKXcnInSoqslUrEXUVYewqa21YWfF8w0GOs3J6iB66kXD8FY/5cq1F4aL9idXD4A4n
VcSEABV2rapUTQWHvxT9/hwHC/h6Rzbl/MUjU2oF3oG8ESoen0E+MkF4coYUjMSthOBBheTQUoT4
bJQWLpDKyvSpeGILF5D/2AHU2nztl8ULBEhqZ0RVRkxvjtqWGol//y4ZXDX/S5wQJ1WynaWwn9U6
0Ul7fcccUNTpg6+hsgH6O/lhl/fkFjkl0FiX8DSMtU1PGudAGz4JXa7ykCWCFFlN3dlKa09NCieN
IgrgTZ0A+rtG4PdsWJgyGjDzfjMpIjd07yMDwtw7JWNXQX6TB0N7Ccgk8JpBtGKTo+v4liSPjutv
sEbFoU2NBv52hsmzw/Hrc1netm+UEoaYA1x2qu/hA1geHpcsqIIOMH6c689mBbN/neXviifBuxRU
jbs6PrSw3bTFZqi67EWG3Of65p6AAR8pt3zgNoAQe216ghLct0sXRRMggH17bhd5JDbnUVyyP2qW
G7aF7Ng0S+gQBz6c31pcMCB+Zbfzj7OTPCmz3rtGTI79N9O2bQVGBOXs+3y+nY31LT6PXIL9cUTX
7NV2GXETcEUf1BZfI9El+Wfk2bZ6P/+Izb8oHgqRHjhtfm1kudpSK04XqPp8GhWvjaPsszLP6pxi
57RSrmlhhXPI3hlOkP4h38vvQ42owpfNIVX5nQVl470E3kGfn1Ln7VNyu/yzP720JUk+pt0eoIrS
OF8CifukwdqNjThaRwnXtYZ15AWSUxTn3Aa7V8p2E7+ECKypsYdsUX6/W5hGy/DqlmMl0zjh9XBm
7Za27xR0YOBWSHM8UklENMNTDp6d2K+9dwXcTYuEX2EfSDff7IBNviWb2AXQX6HboKyRgvOvrc0S
z9YSC1HZq1PH9QWQ17uzNxsyqqm8uE35UT+rbjhJFrP29LuO3uOaz0NErjKQ/Ru5KsGQRdaFDvEj
FyTozCM6rj3Gk1jorQKFnvsYFRUlp/wO/P4k84DQ2k/DpQbp0t8jfoIJ9wtj+eFkpRV1UZyh3CpQ
WSKA0krgLNELmH8ADKwwHBJcdwdf8HfiE4CqjEqLGKcmG/7a0zg95ymGj0CiQlETm3QW+FonjwTi
/nIfxM/oSeZtWnG4sK6w667oGv5RrtnciqGhQKk+y+A+FJ7Z/P5LRw8aTFCKRpXDipssiwfPE5iF
Rpq7ET7hhh8dD46Q6SJhOGcardCWbCebrrWmqAUffRVFTfJpHTGKK44dxi+e9I1qjfnqq284iqyK
8Ah4OZOiXGN0d6t0uQASx/6xwYXKHRMRNM0/HIHKLu9i82sl139gktdy/uaJ64XUM+luYCqvVx0g
kUhlIjbniL+AcZB2Bg2BBIFkjYZBbysIbeKeh555y2lCPhhmogGTkASE0Y6Cx00Geiwjnb18jzK4
cpQpLJgQ5XaHr3SGqmTQRUG30LheRhA+RRQLWwufnYoCbkh/45eZ6SHIk6z4ycHNviZzi9l0+QOQ
OTKmzQ7atTWynMlFMt7ayxJ42v/5Bl0FX5U2hlwy//n0xduyEVrGP1Tpu5GGFjZLkt1ub8bv1JNf
Sp2ARvJwu6oGizj/7M+RDcPxJHW0lJUrkPb2MdB7x/K27dH92dXbVtGfXAp3kxRGTQ/XF+rV6By3
dvZAo6UVGDxc61H/F033hR9aYSeKTZgbpsQ3Wqt4RyVS7uBxdKUwaDSBOKD6hjEVXnhqy7XpILld
LSHxFTqiCuvmuwZjkOfs+Sv8l7Dds6FJXZDQ2Q7Plb32EvmKDJKA+ZvfLj/l54wLQ8y32lkW/f/1
QAKXdVBSvLlKag4Z9ZCxi8RpkKsrDzlD4saLDYykJln7iociiaIFebTnp1mns09D5pxNhDNvZlLk
LL2fetOciB60f3CAvGuQJhxkMDDFa3RUglWL1+t71lTKkqIb2W5ARuPglahqtcZBxffi5tlRZETH
xqg3hrRnyTSZtOtpZ9oQXBMwb0jSO7ZEuxc4tjMligiT5A0TYVUdyGZ1gUyB4J0Fv69E2wZcDUA/
wyU0rOJnlVxqzCoqly05LH9Ug9nBgowt65kB4roeOaflBnzn78/9EfQmMhlqHtRTvFBZPJv3NhnZ
CGxbEY6/Lz2rJNIcqgrWwvtdy6VrmDYBNBLrgCgILwqr3unSvesCe60J2DR8uhF8LSMUV6ScGW2l
7wva3fKerJRh3BnvVvsURJLtp7/QH7Z7VGVrll1+y3AuJMUZambMieTZ2JDJNWy/DgYuiPx8TRlq
UXHI1pGEqk2uDvJS+21d3ded4yuazhLB13NLt1Ya64j0WcEgI9+Lg/uDByx1sjl0Vl5RvUBeTDjS
g+PxSle8wLnVjQ6t98kr41dZ9HN9YwvUfjJ55C+EJvqteyNJb3mRQM/yTBOUnV20RdJWAYDaahWv
E/iGJs/C8dDkgMlO9qyhd2BmcqmPW9Q5egiZF6B5PJM3IYajQodVZoelEzHJVnvZBhEcchBXraRx
p+6fy4Bz4aNn1RUIaMBJ+3U0F28ry8/hN37kUPgBSRDUGhyxw1lJMlhlpf3WVTTWaGXytRMrae+W
ZQn6OjvloQIhYK1Cr3jXu7daW/Co06Inrzi3UGmdhESbNGIZ7mEB+TNRwz4naB57flPomviXsYXM
05dSCpy6W2wnY8bd+vVEkM1D9TxA5OTQ+jo+dSjQKe4GR7MjjBCu1Id4tFFwiKgYO6DkUD5/M4x7
H/MZKwvRn2B8NqboVlBbbF1RSrl3SZfEjodNELrtx7726D5H01y3oRmzp7Xqgazo17XgcRL7Q42a
EU8TEaaUgF2m2vztmc5Pzgx3YLyjsyfTNoWsoZuqjgezHP+7NNa89+c9Ny1zoU7fLyDbW/T7XqUk
9dWN3XHyT/jmwUAMmAwYDKU+Pm2tLBGce5Kpl0d3T4QWaKDmu+JqSzAVKl2eHmhZFGmIirgmtSWE
L5kfOqbaOqyg8fAJE1KApEXDG3O+W7VAUN31ZMKW2oefJDDR78oXi0ywhz5IBt1aHwAg9v067FdH
Mp4++R+NVVDfSygOCgshK0jzVoU5a2AMK4qCSd6/eRYfP6rLtXQTxjWL9SZgCRTvOjAMxwxoP5Jm
56zWusXvYGJUBbs86hiz3j2U9ZKZ2PX0qM888mptDmIjv9sp1WKpPw8KY8g47SqxTEXj/gmpBz0a
YENcbs+JtfomxHs4qE8P78DPuKPf6wDYhDzzp95JSAV8vrMIO6YnRuAkHKNx1DVHV/LhxhJ39mbm
UOwKa5gCCohddXsiJq9h8BAUGd5N7P/h4wLaN5JqwZcyX8E6x9PO/QRXFCXMyKkh6IiQ+Jr8npyl
KnN1fSaIIaLhOVTp8tMqvvjRgU31CpBTX5Ifn/R1osaflPQ6rGRX9s8dc13CbSp0/DahS2ksekZH
y7omwKnzYDG+zkLWib4xTHUXTWF/0tR/poZp94/xKuenVLGe9uXVcwHwTGoVrzDgTTgzOzWca+8i
JQ8eBIxtqo+MGnZujCm4BBrsJDVLV+MpdqSIiO3nF1l72yP7kCl6DQfELB5O4HVtu3MABXIHDZje
MPk9tblfRwHsDrNMtclTny/mryC6Vi7r1X0L/hFpykk0UjmNHuw0iVG84AfAvZHG3o8rac1/ubJE
LYnNQE0umn5qrJzGvOwqAYZLyVsLQ8ap6187W39HFttddkx/Df4UEd4gfp3PzgCI283tgbn3CB9i
pIMIeP9xAGbaUjb3m31sxuy0Do26AOJtWzjz+3Kzs3jL+RZcQqvpzg68746UdMfIoTGJMdvCXLTF
7HdPm1V3h6PO5SPT+fIcYzwWB9nosBM5apHzpG/l+jsoQl12ljcad0jFQnhV9c7tvXfkyQ5f/9eY
2a3Be4LRNmVtXOYqHMnX/4lmFqAqksI8MiKMfvLPqKFsd/AUwyP2Z9+xHN5JvMMv4+9J6nt2itPs
5obwr9zj47OYMuMy7zl8kXCGEPKxw1iFdOoIdYEQ1L1HSYzKLCn15cbiL3nSjIbC1GaWkql6ZlQE
cr7Un5r0yDaxDU0yCFM3SWEr7fENsaFTmS5UcCtCg8AJAAzkxoT/KtLG40lQIHD0vC3dodTirj7s
Elc1lwjXnooHCbZSLt9w1KVTU6mp+RiPIl0+TgXUM4GRcOQMT8LWIXknsbEc0AvXRf7COG3cQPX8
wsuUhLHTDntap6OpaEODjTmfhnjSJ35rDQ4zN2h/al3wVXvRRBRMaz79nHQYEZu+pxsg75wzbR/F
WBs9VA75NdR6/xb9ZbgL7x4wdV7m3VioLok9r1twxb0sfd1UZK+Grq2LJ7dHfia21gPJIriAfLOs
Rclsi19UMTNbmLMi24kiUc17HORGhRg7S+uSR09ydgLuPeSq6CRVn5IH2+M/r+m43xE0X9diJ5fI
WAFWvWoWxi+LA/tkmWoc0rDr+vVopHcpv8Gf75NEuFVURyt8eU4iUACuLqVNsyBXD17uWShjlA/d
SoQ/TSm/RQ2oYE6e606hjFsDVnrRzHT0zy1T54FC+sK6SNmZeyS5xwvz6/jVMHOA2Dd/q7rclkzx
GHlznMNBCrhXSCzIFPmaOpmMndG/Sk52+RcMb8xcLTR2W9Z4AFTB4xH+WXYav6qKKnjuxxfiKd6N
TejwAbvOE5BQK4OwrVW0zGS3WIbFZwU2OnY+2rZlBvW4QuUqvTYQe0qDSBmOmMtDzL31KW+TiTVD
oCWcM6l2QsfObS463X06RghkBefA/mG9ERAD6BmKoC+to/hrC9qnIp4YaSNrLzV0B5GxLJH0tQ4j
I1Ric8zjZRQxR63vGY38PskKxIUYwHgcvr2BpBI4AMiPA+98LBsidSlU6csBXk/nCB2t9dvwtVCq
RVjO3WH9qbjCKR4mn5O2gFD+K45Ni0GJsGMwPO3Zm2fFnpvnllP+TX6i2ADTnTi3IlyPTUFueSfF
cpirou5r76kZYPjU3ySCxAK7AUia9m0rZKct6GaKoCjLAZIcUG/j4Kem6NgxXRUbUIqeKWpEvDgt
z985UwLBouvpbYJ6RxiYfnGwxvNRsyXNdk+uepzE0JhzaJNvLHh2vFaiKzVBQfqOdmFJ/qc1p53z
62vRzgcproFLdDnEAgqDcCwVMFNR9skp4EWsDB8+kQgLh0a+X3mS7ovtMhg6yPM5fGqL/WayxCpQ
9W+UYMVlaLkZmWbdJ3TonRL+Uac5ig1Op25WkjxPWOiXQXUH5hXHEMLlTNqYJpfHjgMBdi7hNcqP
KMtXlkhlrs3GUMysCNmONs0CeFUD+kRwEH31FZVb4kTz2oB4hnBf4Rmve/Hm46RJSjASX2hnyd2b
Vf54EEdRsqTFAlPOgjMdw+eCToXdd34znSz417LiqnODG+x813xKsyz9hL7G9Jf1sGsOOl5zbQGp
zZt+DLVWsiPHWznh3gmDrObBxdos2mwEg13CVK8GDvxSUEtubyg1ckib3ZmBbqMSpwcldfuZSf1Y
mWzatCgsC46p61tKaEOWtKteLsW4zYkCFxMqYfb7P2fYjgBUDC2dKyF/Epa7Odv4cilOoyRY81ht
QksDu9cpmrsvQ4pLxfHWNXVo428L5RWIVFlEbsViglN5M4OvsdJ3feJ9Igrvp6lOJ1ouc2YlzAG3
ETj5NUM2IB0qsfGYler9VHTp3/7Rt3YOhqUkKz39T7OYu+6n8+N/Nio0iXV/lfD3FrsOs8CB+kdq
nK8HOot6VKpgIthS/ai2LRaNawjvJQQwt/grFXsDy8z1DAw6iWv1GA+pUSmFxiScP97dCPBcf3Mw
BPypstb6f7yNgLepj+cI9vNQLi+23RxP56tSjCylai7HeaUXlYkiFIrTKDOWvzgaP+PiUHaDlYZC
XCpQ/rsI9nheJtB//KtRGhX4D8tXuCJTEFZv97/MuK/AIF6yS72BlnfjnglL3JlEhtwNRvqWliWX
BXgh+mYH6U5O3/LDh0Es1McimaFw9ZNt+eRtY5TLv1YzJTHDZtd7DyX2sraTMzDhflk2Ndvd24aR
hYoDWERJ9iwDo6ZY/fEkI/CgGUZE2oKohf620jMbkjdob1hCq7SBJmu8/3n9EFSuBBpBeZoHpbZK
JtJCjwllUJ+OfxkLY9M62UavtM4MuXIUGKJILT68FlsjxB5nACv6jLwDhUGYOeReyEshWN9+sU2a
9lmOLodf/NFFaIEwonwXLueal8dsVEBnNs6D8uwVjY/EsDOfoI5GZqpZ1NA00IUhJX/mIZ7Shgij
4BFhzC1zzzF7GA9GH6ZVmCdJoFfS/0hDf5qtvByPfp1HaM7iHwrawHVpQqhYn5wlwAACwfO8M0o1
X3JRlCGU9vefPLborIje74Gx4ftuMCvPtpBglEoP+8HKUzuX4TbR5hMDzVoz4A6IXRykCN+HrP2d
RU+r7XGMNqN1WepxaGLrIFQtRQoCZ5m0arrkDb9xOg58qTdt6PgldeH1P9aYdAUpDBATN42Co/lZ
CSRAGPLlFYyt40QVQeANenZIOHOJpk+hkYTZhrmIRfHWV8mJV45wYS6KXBU/70+Z06xsDyOMTUZK
O8RFqTfppE5j+wSpxuF8SOHvpOfvJVQVoBd5v93IrDCsI3miN5/R/9VB0VA7RkYiacdFEidqC6my
Hh3o6Bw1QVfvMHPgS/jqSB8kvp1IEYyNmjXd2GGeTnxfh4R7zAhEUZoFgdCNCapKFYYE8fhy0zIH
EQU5VFAYCecvchep7sqKdIgaXS8+F4Umx54CeTmtwYo1fonKseFhEn0Njckk/QqGdcVVHznBdLAz
yKCp02WhAdTzUrysI3/bciyLDAG9u8h5hENPxSOv21Cj5C318PZ4CtOywfHrzG/tmmrePRbGgaV7
LWwfUG8a+UjF1QYB1jJOpP84spaXk3dkdBEGFWTZq4xo+2eMwSk8n+ZFyYniY13Emi0qEKPEZtR9
jVcEqxLzahmvE6uDvt3o5Ua0P+wMizQakfCFATd/mTRrNOZwWEA7Fr5+E9o0Mz3bp1GmHaW8tjTg
OLMjFWkrvKxdNKKFZ1Z3ZWJKzBI6kwvNuH9HcrBfQDz4LwHnRLaUhPpQ3fjPTiv1FmEVCscqQSSv
0Uu8B9fWqH/V1H/koT0XkPrTFy/HqwRbZQ7/osm0H+z8VN3qbg1T4VKn9qeO/zoXFQoDBBxFi5ls
co+0L53d3QvjsiY7jLLX1kJvL/lV5jkKRhssStC0cOmrhlxmlhI70kIAcBSi1xYtRZLDwIwKu3NT
vzdoEg2G68+dfTcdYbJnP2JJHaGtIefsry3Dz7x1mrN49qGUlDOwyUMQTyNOL92cjKHcoJ1oq5NJ
8eJPHpHPiJVUsKgb92uZBuvLYiFGZ0ZHZpGC52jR+L61kI7KNFeFYJWLUQZ/L44HcwcR1ThwMAnv
2efgpdyVv4IO7tTqk5dgOFsQNU+n4vgiTQE7phHi4ix1usdl5yJhmnzMl18Tqz6AG/drJ/xW55Mt
9issO0TzpSTdR/gdFXEIoD2MMyLE340gjR/Le1j1gkGM+6Y1QCIs6HLsQTU/8+41RkvL+IEj0qr3
/rdgmyQ9/2KDLM4aRoaM5uWwLj6a3di6re14qlETCl1XNFiVBnB/07ZUXDlP3EWYT1RV1xpjOiqe
s8tgZ9Fq8xHRzt5jYumy8UiOaGBdciTt+vJJbZ5M0h4DGWaGbI6tp+MK5HzImHqErG12zcMo/rkb
NL/vGZmDiMpXzZ2rtMZmjKW/wGQQr8te5mGxBYwOq6nUwxTW8qc8XA5SXntsDgNdCmCJSZYVRR0n
wpt1e5vB7HjuxG41ZLVg9i8RJSg1DiI3G9KlR7NHCzbPtunjWQqtsitD+Kw8enxOxdXHFz2mZL4l
rmh+6Go2fsC225tHUV1MUoJqOeABvZszBBevzUlm26TzCqhVcelH3QlgTtsJBU7YEqVSngn35IhO
TDNu+VDTs3SnJPNzbZYEgJHqXp3YV06ReP3Inv5HgI/bkC51M0cGM0b6U79OvHdJCAsZTM1Xz3Ni
Q5q84DkupKydqoXPfnc7X1Hl1oT2rMI4alSPLXCPshsoFS4TjW4FJNHjcm8wRvpNMSQfN2jTbvyb
24iJkFmgwGrSWCKbtVTM5e+7o+gVay9CiXchng47aA30+Jol++WUuZ6OEK3oMVhTvQB5a9Cpa3Ld
iKegTwuSKKuQlmeVyAFCjtU2xgBd5vVMnwwuSioXGCaboH48eW2eJxFpCE34hmJ7HKMHiGOTtcQ+
18F2kROh1BHXCiZWA9TCCXC89YnntbTOS/a6FiqGRx2OwyO/10cgv6k/tdPxDdgyG4roXhq+0Nsf
8sDeV6G0C6ETaqPYOdyk+1M8zF39iIV5dypZ0MwrfkDKOpCLbeYLGn6hriIdaTmK496YeU1tGuCw
E95EksYIi4EWFqJoHh81jx9HDGfpX0+POZKVKkvuHinCGdEwvZ5GVENUVr/r8E7aFZzc2v6rUoaz
LX1YfkJfulywJLWcQPRNxz4NWd5zED5So1c+eh+03eoPwXHxuhqY+4bGE+9IXVZ6ATlHX46VnYpa
givXkkE61cLEWFs5c19SITZzRRXVgbeVucOQrVvxyTEVd83Q5Q88D6y8O+sbG8+tfLXDA8zo3vOp
mpipSAuNaqr/XsncKYG7QNTe3balEQs4Zk8sKLiPwEkMfoPEE/eLWMTuiY61UUKssGhUyU+uR73X
dehvR1qalbrqoBNjvjvDjgtp2TsKAbSTSRIIsBIcu2NcQHN4nkwxWkl+5UHcGWmKVQ+uQDFQU3+g
5miaGkbbCrEl62XncbvyJf6jwgaX6vWKACNzaZ0Rk9i5AdnGv7pxu1kvf/GIgQKtXZoRNShRvvd2
93XZUkH/Q4qv189ejIE44cDUotrNdN+agq/FZ2a50YZDqntBGv4+bSFnqalRFFikQLTS9d29BZuL
s7Q7/zUyWCIZh3stRPsp+1MuYUxPS8Z1oJQ15WwtQ9ToCTEaIxY1DAzvQSw+4zwDsWLFsSJxmtRX
8nBdavDcMYs3iGLbw8i33+/fMyu9dGw5VA1jAzhUu7xjFKZTcH3HPMlCM2bWZmUooVbWPEMzlTqM
IGvvQwRAicp8ePZyg60ukjyXxTy1pbKAT8AUiZEKy4AJkaPQscjU9v2cEAFgEHf42VtRfNHNrX7e
Xjt6yKxRS1ZFY/D/dgHWjAr8UWHWEPTKojCG/VVbXQKPxlM/ewG0hpV7Eayrjbny8C7kR1/8bJrT
Hd4Aj3k0TT/fiY3BbKl+RQO2hBhtd17LyFcsWuJ6XPK87TEPHpmdztzZek+H3Dms3dmadE4mLqp8
wm35kqZ8a3H2RaOf6LH8RJJ9zVEZAY4dqtLJqBYT4eXv7BDgAAB2hyDEaIrWwm5w/J2hw4GoXtJW
/byhpKrKhknDRhSErNnwvoxGC2+pTQ5hnFbYshvaU46KCP9TW5ahLdeI9l61hKmQViZR+X6Ow3RE
15gBUA0Oo7xBZZ08ct/tvL6md23A7FNPUXmNgj+9gpsk4+jgxrHLEofDH08JbCTTlfsqrqaqnpRZ
JKfvrUUSt6zFN2vgiJ1+CC9ITh3+e1AbhmYGaLzt6wwCD5plhy6PLIMFV2dp5Jq2t8F8njhtv2rd
0xTsaXAG3oxrjQBc4i+Mr3aJeuKy4iMTwsdwUo+En4RisnNRrLmUzBa0osiC/X6skHmEKjJtsYbY
tfjpnTWl5VAp9QQOk4ZHnYbb1z/YJhp//gHO0N9Fi1+/3WkeduLgC2bUBvD6Z8uO6gRcDQjCbB2+
OiDFA3UyPOoMIyHWeXI+IMVEsuKE1wKlwYsL5qn4+DbgqZ1J9EqNDWiI4MZS/wnkzthqshze/5Oo
k2e+VmmJie/kTkCpPXkDVSA0Qkc1BSXWpEslUo4lnRIbV1SUGRbsHBu+5oVV7pc5Rynnavq6eOtI
3A+33FRCsXoz3xjAXuFIpA3/vtBB7ruU0tXvTUjK4EnKitKpCKHDlbOtKZTfulQOpH8fT7BJ/dX6
iCNZWvLaKG94ccKQdW/1hJ08In+zERg82bjVjG3gtRmlN3F48mFW+HAI4qclgSCM3BsFWg4MBTaB
U7p4M7P+ygov1Mt2Lf+Nnzt22MYNfTt2pB/XIV1xAkogp8GgromwTxvTSUxaVV4/2vcULN0NdXYJ
TNC5Owum3uHGXeZPV7mX2q2Pu7v/Lah0ZeOkwnhGgbmHgvfGzO9K2g3oR9dsGWyqTF+3ARxnoPMQ
knj+6eDcDIcfqzEBqN4qWeSZTid66wjC0MPqNwC6nAg4nMJlJtdhgj0uACxRbpSHvJbBFi04bigy
fUzjjDdzqigVXD8VQmI5gcwB9bh/ba4vMlgX0U4U0GNA7mjzZlgI8ubDi0OrPhGaJdsPgvOo4UdJ
K7AK554exSyf/TwMFbtjbaKsMlhGJSRDICgpZ46sZ36Edtbqv/vVqId7FKYPQtVLxYWeuivkBDmc
jgxWjkKqNIHsQ6usB2DDgpP6NlX2wc9R1rM+eOWQuSHW3TqTbihKZNRrCyi5oAnp38uce2WhUu8O
1qKSXJIHtq971naCzXcGK3ABoO6hEOVootO0uvb5m0CqHRoXWSDDJM7YLaQ9F9/3R/3ml/vpOvv7
YRjzY15VerpNtNBPfMqgIS5g6J6QuEt1SqN7wATz8dTG5ZKLrXACcYES2FI10yPfk/xwcnem2N5F
N8lKJOqy80bMbJZoQ30wL15lTfaJYAr0NdoWXCWh6lj00mZ50aOJ0VPmV496vGCfbXiGKr1nQ3u4
7foe0KOb/YG/LpPTaNlgxnPueAJcydAVpcyBc6YQmB0c9w7UmQoqL25hW6jV1SCXSp/eub79s6pw
GUJwjix4fM0BQ3f9DQQrPf9xgrZSnD424GyV4aBN9imPEUlX47cShPU21coIoQZKrl4j5PXQKwYg
8SPrddXZc4LaPw+Iwq4JuDdm/dw0+7+vmlAJOX8RytDuZTeZ0pnFtJaHGECap9jtCH+rLhVEgMUF
x2Mwg02mS2qiZb34dB8bF8kaospo6vgbuOrAGSSoAZB5uN19aWlt7f7qo9coRvjv93xP0rsNqwT0
myLBH3mFSt6oEubvBhCMQxNMcaFDbVR8QWQDGyWaPIlIkUw6UnCS/I+VwkXpvq/7sQgGPq3Q3JUl
8WSjEADRbQ83lb6PXM9j/GbunMLWfBlpigKJkXEGCagiNLcgkeMg5af7UTxpmLThNMBJHiYOp2tY
sKDVdku0oQIj52VHdpvGzX3UF4P/eeCHysmTRYzPjnuKMl121xarz437TJjc4Cbq+6KILtF99Dug
4a3dxOy3xNS7JX1hkymQHWsyu0QYHVdJ7XQrIzDajtjSE0kHVO+Z+u6/0D/7M+8OYjp9pcUjycZE
+zNbajkztwlc1vsod40MmL36ARhbMUKKmyDtkOKaDrZ/h9RgXThp9Q4wx3b9fSyAUyKZcrXd/utm
3wq3nYT2t57D+t8fV7vsP8yLCRHC0ZXbhqWiS8of7xRYzfJjs42Jxbax5Q4mK6sfKvBmQ1H5zsH/
kOQY4Firzsz75xiMvf0EASVQM9risFAZeA/tpVFJBF46/URObCnnidzREABrfav5/ZbpuiNEXbx6
EtSXxwZhPInUV+zHUlWz6KuLEinsivu6PbV2xGIMXe2qqyyIgzWI1Ozpp8A4A2gd+RD0+o0W7wpN
N14d8tdl++GSNWCrIxSPQfXc/BMddJlkcVUFCjarX04pKt/eQEpBxraTCavSSxxuGRFZpNyPcNMW
KQ8Px7gz8XPx6CNAQLJJA4sMbLlui+xqyo5vJkYCHaosmmgRtIYTfCueTbq/PvMSwLtZSn/joqKA
+RhSp89YEV45fOnYt5XyFmoyN0DbXIAMllG9vSK/4tIHL3OBF6etPMltDWiqahVF04D1fSORbut1
mDIx1cmqluov/i4Qzeu1Wfl9KplywoRAvVdGb1KGwZzPpaXVGofUdcf7FDbxLxDoETVZtukKHeh6
40U26f0lJkALQdQ/3thT0OPbWvXsgW6hPQRhxwMsZ3OFwgvK+rRc1nl+mDJ3h4Mav7mawp65wJJE
No06iAMV4Ar/qCCh9BJtBnCCKpoQnDkjomy8F065JU2OJ+OUy+wmxH7mVvxAYOA6LsuXUi4diz2E
iwKF+qcSqMcTiR8tk0p3sNO10q9bCcNcRAGarZZH6io5T04zgykm16Ne7OWhIutptgwu0Jd5EuN4
uMy3hkEQRYSX6O6TvQ471uXGdxlVeBAWNpjdYxZNd9PPY0zF1NXJXpcTy11Vet5XM27hPWr3VbtV
incWAH1a7wUd0OJCu9eZ5fAbgVhIuG8s3axGwoKuhURhR9vty/w/ojYD+5iGfiwz5ZYxdh4fNtaz
FJmhY0gjGJIRHN2f8JFyX3ArQI1l3jOa3ReOXKm8w048m17Za8ndCkTJB8CFuJrCqszWnboQzqJ2
DBJLjrM00BNbRyYOwhFdWcDSVQnL5DYUsNXWYaZqqBbnB+sJWzi5yoWN+Hz44vie6n43GmI8ng4D
pgtK+0sbnx2zBXW3Qy3GSeAQpUKmQp5ZUah7D33ZrqtYkaZxkAOmipgJfEzma1T/Xoh855LKv64Q
7eUFdzhhKvdiijucr2LnxcW4HVsNRprTrMxfEATQQTEwjhqln9k9kRt5dV1CBCGXHuqHblkteTtM
v/0+xJYozkivETPHn/MgN2BIUSGCydXDvsVXSFB8Bzv6s1ZNEvac0kpbQdI77c8ZoS/AbBLzeGg2
ARaP2zvddQ1aMoH4SMc1OC6MlTXINTqRk/LU4c6sHnJqwuuwJGv02YfTtLmQ1Ut+oy48rgkUkawc
lW1tQvncM0UPPYINIoQtXE4o22ECMubLXvjHXU3uiQ4X1Q7cUTQujnq2vBMR0dOp74tMfIjZ+gHI
3ETSi5vYQR7NZrheapS4J2rIxjI61DQjK6LkzmiyiNEfAWDfb073fkQYkcb8zyBVuVtvlKGbrUi2
51gzH58N0gXj0I8FnSoDNAJ1BuouTynWpff3NEzD67JJnCwIXkbRRPySaxy+zkmpaRHJ6fnMc5tn
QXUA6bZ2Y0pZvZ5heCfNDImDIUvh07Gc8UFmcfMKUmFBvVNWBx5La6ec3EHXgMf/Cc0cam03LP1i
o9jOBi1jZmxVUnzF73rQBF4idZzsHDp//Tfw7aWIdmfnloV3NG1FqIhnrKPjxUtr8f4fg4LBd1DP
BWOe63HzvsM514Q0VK2nztlE/x59CHg0JqUFuF4eb7w28F2RZOSHzqeGrhq3odyPSQ5bRRyVARwM
55Bfj2aZVhNdpVMbCyHRQibuPWllo5wRlMp3YWzKILjH0XGu3BZOoV5R5jT4BiHZhnmRoJ9MHVVa
ZU5xq2XFkc0bUBRl8dxIvjwknCiAbZjWhTLJzpSs35T4quq0LjInAf61t3exiKLrnXOw+0DnHJFV
Ee9l5KNp9ei2V4XNesMe8Azbuc/haMlEHE8N4Ks3zb0CT0OJd1P5lzCOPzJsCDbSzFlTYL85Rha5
cuxCxZlhM4cSNkA4Q/Au8cyy0oj1NJZyan/SMG9qkTjOzp5cfV3tzWKj9onHpVTAuP8uR4vTGAIF
uZ8u4Jrr3KE4ayPY/DowojS9j/m8ZGfrBJIK8Zu75wuC4zMBTX1LlC2AqNNw3uorUqazBMJ0Fm19
Wggeyfq2oebS1SytQKskUHV9IdVIIBvxEvmbQ4ZY78U87w2fbUhLRsnJsHedC3AA/z4okqsekaCG
0ps+YNsvnCoUiA6hmLSVIBK4XP1g+LmRk51fqGj8sVVwHNl1T+wmKG+vItGx0/4Q/AL+eljnXM1f
4Xh8VB4iaZgyLylDVi8+MIaSSa+u8s3hphXJ9R7tcRP99gbfWw0q54f9K4o9thzUG0I+bo2Zm8fi
2io1P/clnyZk14X0jBWUIaHsig6ddiuLyV3YkhSHUZHr9zYkwTB0NBpKf3cNWK35hsYmNfusYG5a
pd+VlRc8wWKYaDrdvW0qFTurNg1BRBDGDzOHMkXkRF/ol/JDdcYlYAek/1h7mqZYBPBFrFRV+XjZ
aG9eYERPaO+tWvJlO7kOLlJ9ozQZbTvyCid/AxbWl5l1NXAJM3l+lnLYTnQP+hjMob9Wc8ZGBey6
MJ2sTTVhoahqTa+Gh9z2yI4L8yj+KmGRRV7uk6ojNLp3jN5n6YV6UPC/Ipjp4Cuc/DK9LMaanl+9
V/M9FYKp+aUKbLC5USep4j1vXYTGihFzHFqokNkvjapyEqXRs7SH3HpOsSBePaqCofxudlOtrkhA
vEZOwDWd3tkcNxuwEryjgaZKuq5Ujm8wbvyKjRoRjwPx+Pp3Z9r8/AeuL9ZfbYxIqvCFlhSWWs7e
RxHcjqWCcycS1NX0ZVfN6iWNpS/zVHrNKTyUd5QP29ligbT4Tx4P/p+Qrun/Qunmdu42vWjF3vlI
rDt+qIP51CknPwRZcnpYTQ0Vd2pwTbmWRydflUgg6mhLvKFnjyQ//z8btEgXyluki61w6W5SVDYV
HSniWj22zkd0zrtllh7JmUxpqAPuCgXfvZ30FDn/+zLAVLssOlR23MLYVrsG4VS2kT3MEUzXene9
9NjWmYmpaMFBviYfqqPIFyOml59/dtrk1oE+BEP1JYEokLsx0sdmh0zcsHZKoOZvxHFDohzVBaej
9WQkDsA8zjip3xfF+/rmV9Xu2dwbUgEUKMH5CS0P+1lIVG2MmKY96F/Myjoimga/UYSKegxCZdL5
q28+36dZGJo/EQ9IlijJzeTphppvZHpVu/2sAFSdRz8ThA596yF//qOnoi9LT0JvPPc0Z8SIL8TO
dbLGkzz4MY3mfgWBLFBSk0lHa6vivcr+R6IO3Zkbw3JKism/UHeJV0QXLMhXfkZi02k4VJBkVYP4
ga+FVXJPanTJz6fpPwhYZlaocBoh0sqZSgS9ovLq6h1XUyJ/Bwx3ptC9Z7glZyFlYwKsavx1NUZD
w4BQh+j14JurYWdu4Eclft89XUCYLTSydJMlnZNkTiZK5y+czY2nnbb6kfaB2LAMunFYSv28a4mn
dxu1sOWX8LP0rMANUWXZu3E2dfZ8DW9O5rSLae+dpfbRhDlCHliOOdnKs2EpKEGgip4gW/vOsmc1
ZrRxDO69PLjo5uvlTKGzbqMcRd27HOB+uZYubXtpo95aaUK4Yxnl8sgzQf94nWeThj+6VuEtGBZk
z4x3ybFcPE4wRmocVSvgFUekdqh40XCVvsIYj0JGFSbW0ICD1YoY5V7ZGjllSqg+8RYdl1yBfML+
Yh2GOehrrZI+cn+WiK03pBCQXPgyCEV5IqwDwlLzzO93R4KUQ+QeYLq9M6jyY5a0bz6uR9Y+y4wu
3YpMllPbdx4FZ+YZwbpsFtW34z5yJiJSe44AL3Jqi/IIeXfaYT8fhVD6wRwYAbwskQAqbXBiJm/O
2a7PMcIYP/bktswuM18HuNhrt3Pa3ndBDRr5pwR19SSyHP8wsxsFqsZMm5P70K8GdMQK/IAyeOX3
45Vtbqo+FXHrdZXKr1bWblFkp454F3DZBLMptkxnlsuYNDXxcET2yOtBOcxtvw9eyOcr49gdq1Ik
WqRkDrgDZBi57gigMLkOQqIxC6zvARiWgntDU4CRLPYRSkf5h0d2m/cy0aDJLxuAUpZpyotCMpT4
rSvuxJKq3qeLZK1S6L115HhDFP3+oXhfC1CYS+swU40wk75xn7ID0vIpXN6Acu5BAymqyHjhTO9k
Z//tAHSKdEJbJwEwqYUZS10FiW+xqJ/TPpFp4NmdYABdA87RdFMA5VZEo8mSgaIyDUg39kfrhHou
l2lUWESK47qTJt4LVGpcbUwiOnvaaZLBFn0tMcO+r5w4txtpGe0iFQNeojudZMWUXeVkfTC7SVqz
XN7BTeS3/gUvlQiGLJwckZ+ZE8BusGF60rmx4HmThxstUrPvqPYXkTf7g+vKtqWoc70VwClZtiWy
3H0J0yu5HA1UHVUNjE9hqTHcSxJfgEFOTO6afVAy4jvvrQZ3qigG2bRJdNwaKJGXRrZgODjTip+p
JKM8zlQXpB9U8Z3H4x9cOF0LBJ3lWw1z/4rlc8Qp98IGUGImIdwMc8gciqCysYlOXQEW3QzJYjWW
4DTqlvUntXUG0DBWkWuq0q0eDw5Q7EW6tTbJspFv7v3u11dbhp8jlevYRPPhW7iHUxAw/rgJhtcH
HYl8qSMEwkoXCesqa1CVteQ6JRHEPv2UDnrwvPdnVZMzew0QsTrdgbhdky6mtrO49qjOPjzJlczP
LapaW+Ow52GirOQoE3FtEECdU1ZJDmxCt7sCVkm2ODily9WOaCbG2cHec0S2oDYa+pf03Zar6ByY
pNdEniTWotG5soVOrV9qztWqTNzLgyp2rnqWHuSGM84R2hHaVxG6SLOTtWz3IpmADcX8AqYbM52R
cKUR03Ch4Af996l0MVLxXfhsEBaf4o3IgVGEBugFnuZ5UN5JSFiNnDGtSBUCWFB7tBFNHCVUhpzt
6XVbC70L5Cs4JD83DodRd6PSPWD9iqQ9UafAP3gEynHfbgtpAgE6ZNr59pWaw+gxPKBxZfnIxdKi
fLuKnqP1ngoWStVzaTG5d4ItyncS4BchwzQd8AuXpbXlG6fc3K7T2EDRQl1kcUcj5BR6XgB6Gv7b
Sknab9tKdVu4K53L3t/vz7e/v/eiq5V7XXAN/ATfRy2/xFfKxkREtTjMwWGRsxAVJyi6uKtB50gE
6mt8MLUyWGV1QDnC+cr9kOWNx5OPZkOTIbcqS9Je/e3NX0Fp3Fh4cysIZ46JzfMHPWYUwC+khsK0
LEUW85hUI5UtZKyAHjC6MiqaOZsPeaTCV1OrMbRoDUQQsO1H/mNht45j33DGhYaTsy4uhiV6VhAT
5Z9cAraDG1aw/MaEQ6RMrDSzqFUCalxY1wAyoHk1qfLO7F8RRUuNZxVl9c74duS03/bYxJCVSMgT
CIwz7/7BQKHtgL8c1HiAEKX9vuCwArYjUEcE3MJNZQy0OGKP8zrwLEbJS79TqeuyecppmpwFu/SM
jsTtz+0C2v+KSBKWw9bmseeyyus1EdA3pmy54l1RjKHDwZeNxEzZeN6yyGotSlv5r2KUmLzlRQ/x
erp6O7nCYeEISOuU07yMPkYxCOotwYFJYLdG6i0OXiVr3EUontSqkMjulryynyHK+46Qt+xsvqJ5
w3LCsnTs1vMjLnKOkZvTKjJd502B4vHvg5wjH8tyR63xVKlUyHqTJ15qSCYRWDLSSErWlofA+y+l
sF3ZVHjq8QLR/V5q8AU1VV7WWYEFTy93+GkTts3wb0nPNIjhnX9NV5bTN30F2nDqYgaA2XcYNPeN
xJhDOWJSWdElQwzM1EAuU/zepSE1fROkSEFP6X3xEexNczpwd3RoO+M9haPRRVtk8GWvsUgiD1I1
uyHPAxYvBLpKWabfKqu7Nar4JcnCGb71oPuS5dNk+6klvOqvQ4I5ZDW0/PZsiS1vUJ0uxMMtefs5
C/JxILTTIx0Tk6xVs92altld555F6gWanmPidmjQPaO8brwXLVPeq5xyKZo0Ec6cedGhVqYHgjTZ
go1kHRtshJY+e3hzuIBAA8WpxnQ48p8jwgF8v0669gmisupZ+g5pu9Z9sF+HCSosZA3JFhqc05KE
9He8tyZTDCUqMZxfirawbSFhZ/7MVjoi6Tfeksn5eGZYxWhoXUMOKxn1bpUb3ext+TVdh61FEIc9
5/mJ55ptIJE24Nm4FJCFaCtocEM+mY5pz7vMJ8n5dxtlnopFd6AB2WnjXCLO1oU5EOgSJ7gmhxPd
P9OPtYOXmwXj7Uc+iz3xPqX/D7BsCfLOOZXnJwh/3w/WnSq7MRkmLW1kVbm2YH1HkjZn38T+JdTL
a137m23vjRjj+Laya7HZhuz29wbMd9cND8a5bstaTYNTTV4ibcqZ9X2147sfIbK5Q1l0yIoEb+1Q
9Mdn+7oR7p6piosoexdtobB/Cl34IJuXLNZSddv/tCml5/N9GtBz3Nn9GPik5ZjkFeZdWw/griC/
LHeDkqxzgYQVb+xOrUXkatjQW9D3BxnVtbuFxMj2+4oBA+M7nF2ov2yqkPu5EVI8iZUBasBW2Zp2
yPCjjwKiKO12CzKFuy11P8QllgNBKYSJE5J0TAInahTlkFdnfW0WFZHfGMiTvkmGZiGxpX6QPJPG
dqB4bepYjYqUcu4zYI27wmMEORlKA+c8pJz7xr9ibrX0Ie1acmiwiLP0r0xjUKiJkHD8jOWui5t4
uhXfrCHUFSI6pttUbBUibxCAa8LU4cxG7FYtUSgYFhu+Y54uPHXDNMhtb2wnZRCT7RmwQm9c2N8r
bcVjkHMDk74N2FRaYTQHHPwhkT/MS2efPfne9YgATE7sGeGeNFnFqT1SCTS9d4bL4Rr2hKjq6rUU
dgx67FpCa4MSmPyexsCpSkrdIiWC57o/oOJhCvx9/lHGpfAYwSecuhIx9cuvXFmLzMwDA7a99nwc
YXfCb74qE6El6HjL0H9yecwil++AgS/F0ORi7/8JF6YbAbtPNw34F7QR211N+qAj1oxl5o4jyWnh
jAFrDCVPzWAMuPwN8M4UZGPEuo1R4dlH1LnVCg8rQa2tguzqHslMyfsID2+0Q/KkUQtMSqx9bWHW
foocG6vI5+wetbXyWTr24lwYMR25yqV2pkJBDxjiwcqOQ/5Xk90wbDQUJVig+1BpfDYzXLJUt5YR
OlUF2JjaWOcoH4Dtya0e0GkMhupXs6fWUl0ZhnaxNpHmCUTOOW95Ug1VSmVDuDiq58nGOBo5v8/P
lBYSHsItSI9TCASj0wMp1GlNduCjJlFg8irziY9GaTHz6NXQnDbRfY4uRV8cmGcWUKkmcGhDRPbR
WppJGi1ARvfv99KDioI3Y99IQMYk9XOgtF438znWfOA/uigy7XOhvQSCNxwTKwR+T9OaFH5Cx8W7
CXoAULOMdzFHsY3gBeHlg4Fr029zjD92H+sVjHl+OFlNHMEOF4a9ywA+cxPnC0sY7LVY0DLGrE81
I5NAFAQyZzfsZGRFeDJy0tnO6cG8IzcAXVw/o7ogWrfMPQ0avnRvBwOKyDhHB6aNp+ubqzqhy2IR
qR+HQ3+FrDuzdnA23mK9XGg6brC9aEyzn65q/IuCe7QjoXp5x3lJO9F2DVoCTzVdShs45d9xiUYF
AjW6bK9F1gnQqVNwQ64H6khsPs4NhFsqmmLzqtkrPScTg7Mg0oSgibtd2RM4ji9IDCjL2o2LKqbE
nfHiMOio6nxS6jEVlwbcGi6gPr+P1R46EwDnBwGrwbUIl7vP0VRNjBS0rocMXZpkIp5jrjKlGXBR
7sjktTClSgT/aZ882Lyp7HV+akgxiVIS8a6l5SNf/qBv9AAA0DrBu5jv5ibsw2ygxxiivPwa6obH
jB7StJAtZ4EFST0viPdXJ9OskdBqNQTuITLXIG5+5+0H77V0Tao/F2NxJI/DYXP5NZ56tuoZSznA
bGLHyYloTb+DoQATUvCcLFo1sXDx6fDKmEhQSEwnIz4KNbC/ToHjCScInwPirYwozVnZZ/ABqM+7
OK8JvVjUAc+OitvM5zXxM5gmQO9NO5N7oKa77Wr30fV7k/UJURAFsjZo/ihaZ0eMawC/6xzW0sBr
/2R0R9s5wvCi6o7retJK0hIee6fAqWnuf5K4vJKZaEvULDevE2WEvROaVkrQFvbpmRkKi1lIIVpC
CSWPJEaHRm6lWu6FokwilAo1jbwVJ5VlhSsGZW1J3R2YMFt848Cs0hx+phuDiQwdWnZhwn86SfON
djy2d8MoDKSUZkwLato+0dtgoYdizaW4YufLKDRbn0goiHiOG8GohVIEwjgZO+hcb3cusAKF92+I
Lsc9IjXgD5MLUHOgkXp5msJRpPIUnkppttO/a6DaXyHEzw2EHOuRYBnsX2IDOg8WfdZKPSUgmeoQ
18S3uaQxeTM99VJ5N9vwGorLoPm2XtQ3m6lGXo3vwgYmj386FLhHMiN5kqMjnzF9fV7GPjoshYQN
3/piOnID2VtElulLefqbQe6w3266T3HVyKI7VPbrT4LiDPB+hEwPzMr17iAomkHTwOrVHWJUH88e
1wG+DrrxmoAQXBW4ObP1Jximup27IkhnPgMSzTjjpLzBrzJd8DLWL+k41NZCfUML96sP/uUSNSmD
O/NXxg5vl7lmmOQfFC7dev7sUmbrTNgo3SWDaMl5KxfZe2JEteGjJrG+LdQA24XDFlFwrAFpDz6Y
wO8gliDwy6KOTRl/MVnhoW1UR90AggmZx9HLp4G2NPiU5DlYg2NQtzoIpe4N5kLJsxV42W7gEXu6
EWt5NWt1weSNMqWyR0QSdHq2vEwjEzGLugtMl2Xf3WFJmCtg2nTL23M288sLoP6l9Yd0jNy1WHAs
VWpBOaWGD5Zau7zMylUVWWPYxUPbE28uZkIR4bizQFLR/qdQRlLQQsRQovbTe60QbAMVP8TMc8Pm
5INdr+hHCV68f93LgRqxV/SB72Oh9QJ7YpReGcJ0cmBXGeQNns1wL8Qsgrle/eJJznFMJsB2XFwJ
VqUFXAasM6Y5fwXEd9I8JsVo+x2+WQgTbo690RP/2etcKP549EAvUDeoSqV6x4xoP42QDHiv89Te
wGdau7LsS8yzb0/XUcjz9Phq5o3YchRu5YiGPVm1+sFlrkO7n85yBfEPy/GIUvxFFWUZ6CfvxyGK
uTGrn2oD0f9Hsv1WQYJUS/hxAh2u13RZwwMISk8z4sMYjWQ1tJLEEvo4zYIDi4MQRmyMSDgHKTve
fNOP/tKsaSEwqqgjnIChI9n9y7Jy8a6j2Bv1Vf0/qAwB83sOzUGGrIMOnJmIgMyi/aJvUp3EV5LB
KDw6dFvGew5IqVLwWpEQe796lj4fC8iORHQPN/9GqCtPEQhxPDHr9p9GeHEgv/hddAyFOGtLbdAT
De0TitqABQEgbLGcGOEPPYHbwWaJq4GkKw8P/77N32eUgRfzdB1GCbR+ybOPLTXpO4KmPZ4XgD+K
lErcfd4aSATm7yumrphrJi5EaHc+SC7asoDoPLpu/TWrhEbttaT1wQjNgYJ4UdRIWQs5mujEtGcl
5D2EZz9+QTyfXeH1Sn4h+FDWQVjo1HLsRRVvecoIfnNpgQ6gUlmLxIBhQrhvVbFji36fNzAk5kZj
c9+XyJrUv/MdK0xuse4b+mIiVLCaxiyVBFeqAE3S57GlNxAYh4WaUXAJwGt5vXZNzhg7tcet72dd
NAMagNNYwpUYAzOFx8qeJmcU0i5PQQjn5wrY84ol7BnGBDw1AdxuW2pyLnwTyDc6vC2+YYfJfKbA
g9fsHbS5XQ8P3EY+JMbgKqQjQWCRmCtDwuM2KUtX/0jNgWOCye59HK5DyytEKA+TwPyuHirGkduy
f5JBZWQSMX5p51nO/GJeq95rvpPNl+BeHlZg4iltmqkzNXw3vM+ul7qWMbXrgre/rExKvNb87nWl
/SQY0zG/5Ph2i92OtE7USgA+9lXMQPYeLeZMCjtqW6wW8F03TqKUzS6RZR9MZzV0yN+SKw1KncS3
qbQt249tDmCZWrn/IGIpQCaysGeLnks4GFdWhO15tt5prlukIKv51e2K2Z7Y7zRdjrpIof6H7+rc
OfRnI1W+PqhwLoilLipN9UuHkfSe5c+DjftNY6dl2dh43cdC4/fMt/mzdjcaMPVIrVbONSWNI1wz
qUscAAn7LLtf6XbIJXYUlVd6BnqJF5iTK8SOa8rgBctthweVxAR/cmEfKxnYOv71IzepcaanjNL+
yV0v0TwB8dZ8oZQ6EUczxE26tKPpfzdV5A386OnoSkuM04z1S+2wNYMLoV8rWcv0JMaiml3dHZBZ
qQg7mwu85lEtcKa5GkhQPyj9jhUJEnwqF1VflY9sdvj9c6idTKOeLjMPRkIGLatbotWMyEqOoiLO
3coF43e7y6KjIkrF68kzT6FJkLcaxlJI/4yXLPXyaBthyo/lJaWjyGNvB8p8HYxj9Ay6bVin9SDr
7BCjgK6sUoPCwDoAWCSizY0zYFOP7sYOfitanR8KfnYVeGVF4571whv8IVYWdjXAwDazo/r1Yc1+
XozX9NuCiCLWae4gvSi13DFrZ6lnXK5RHrOeFd6z4UYA0iV0aaifhC+wU0blL1uwd9pr7e8D2pOb
q2grDBBnm/JNj+H3nITOUYjFQqtBanJTm/XolMo81yFwxYNs2zEerxHMFWpiSPjJOch3okRHXkdT
q3iNL3YkfFdc+UfEzu70T1BsA767kJzAE94m44YGdor71gxjNjhi+4Utx1+nG4DLgbesYiRtSt3Q
SX7zTzO7BBSqiFxM3mAH7vRg9I2yyVTDnUbEqhlH8ZjFE9Yq2kja7XCvbE80OZ5SWrP3C3pxm/I/
x3omHfZIibbHPLB+yNNJ3JrrgFJL71nrL71JwKb8uy4ol2HXgCyAt0iASdS7j8iPGV5hsejzM2WB
VqPYYZgpdHR7hAta8NOhQqapnUG/NsmRCFtJeIbJD0UeZ1vcIPAVFP5zFXh7A8rk6Q6gx711aKeZ
xeJoJxo9iAXOLiWTdZ+6DdDSRGNqdIEyulg1CmqZhE6T8Ifti5//YPtiMtqjCxkMqaM9ilPSSUyt
SFHRGdCq8xVUbbXt0HHgBYKdk4vry4bD8X4xBV5et8hD0TXYQtVGMgHkTg6GXUI4WBsgCs+IUFul
0Yey7sjICVbHil08qYUlauf46J/pDfVco/UI2jR46Alym1JafQS1wmJ/0g2nc7nGha0zKEEbrgSC
7+KYEuV6KFAySIU5G8LXqlq/IX5xMQwRJi/4U4FRB+rb0G+6a7/tP3mcJ6B8SQbSa1gdMPRWun1d
wM6xfV7+oB5e7fI+c4JGSy2lYTu4Wcqi9LgVTWwQbR3ZcSwnS0nKZo8lr9aBrBcp1VtOyZFuM7FH
zP+ps1azftxX3nLcHSy7ROWwPAB364+xiYEe/LPT1xzPzy1P2lgLByNsf/SY0yKkDLhF5Iezwfzb
zWaC85ebTxKTm+1qBVaYmU7AIVbIfhBaJbnPzUezxXe55JgNAD7T81SrmelMoojPvTBRbT04rPz9
wTJWK+yYR0Nza8GP8PRJuSC9MV23JkBAAElg+GGp70Vvp+VQmYHDFBwcpK0Tvo47wqYtiAWsZ25Q
AhBFx7lqiNbKoJ331qIcfJauC6p0VAtjoObkCtY/x4SvVXz8tjVbXdwl9bwaM+KrYOzsvK+TrGy8
hn5MEJvgAUmadO6fazcZrw3d5qy/Xm9LC58M7ZqFK1MFZX0FTJndq+9Tup4SYBTcLrxcpoys4CBE
22pCH5MXl7PXCruzBLl/suFcRH3YGupP8+ZsgX4rXBY0LEL+mtEwa9TyN7ce+SPrLT754jzekxhE
o1ULBxcBf9F1woBK9+ykstMy58q0r9MdyGz/tydoC+PVKUljeFxNzfsA44yp/0kEcRIetRFlPoNg
vE6526WoDMQZAQt0WUiQRxSEyCi0YmS9UxZRy3S7L408wHKAiyrLWWvl7y2BO/6hKCkJMz8/x/s0
AqC+PcDOdOBnxYfVY6gNshaGn1OF2iJYQaaR6kWqpS6iBi6H+vnLpn2YBrOHO/4b6Ja/s0x6R+g2
Lt5TTgjAhXIjfB2KJaR/HyUpCXDURiDBGij3hah+ki3clPAyTm6fCBP4jGC/KT/SU7GEQgeWnOj1
cMemVx5P4XHGcR49FAQRtLubiGS8ZR5xgfaorSe5hpj2MY2tn2Zd+KzrcJLhdet51mw/1etE+zU9
8fP4teruDDLvD0Or3Sq9w/n9kxQNxaKpHIApsuOgP9Pbcl5w/Yo/5xMLu6+plLK12+Qqf6w/ILqT
3AX3evVcqSb3eD4946e7pZUZjRP7tpKDJzVTJuMT2CmoYiRteqw8bUKln+8+eyvOFufMcafNUPaI
BOOGAnhFryNDJcQ4dHN4JnfIj1643fqbDp2Hzc9UVR5y0GsAS5KgJa9wPTE0P4ie6YnNVGaOXd7b
OCdY3KQzsbevhRu6eMlwIv2HjIW9SmDnCDzXkrDvwaTwTu5CC1hxXTZnTeuaXcyEEoWy/bS21Y8+
35deh96idmdk6/9PlzT3MoerKMbf3LKqn4VkM6ibAfIEMGrJkAGaDZIUSmGSGIejGtcIZjd2Z3BL
Snv7QdP458BEPvNl51HSxgmO1o/AYSbaesAKL3iWV/fy23w/Fs7VcX24lugXtCNPdbl+g4DvSXW1
JtgNqRJ5sN7rBYiK2P4/tT0XZLkDhdpdaQOHt07M+augx9KMQxKrL0RPGGO0QI0rGfhOPSFhFDJ/
pe7Kn6r9jPzGHshGxB8QhFSPYmeOSJ6c9BUiBljo+lYnyzptOre9V722+4CW9BdqDwstHBsVtJtU
vffe9UhdCrCUdNoDhFN8Giyw7RrdaBzdQ0pmaKsc1NIwInN5KG4f+6vuFiOeSlTYh3d7co7AOtfj
pwXmzbvs1KtU7/vdMs1pC09brJSz2QL9Ea8fakLBsJiA0z/6wcv4mhtBsQiXAN8DiguZw8H4Us4f
VV675xRlWun4FK7IGiF2sHLAI5KFcjtmdHjzVf+iole0wR1RCaWKNEj4sSYwiBpS2Qr/6L5dtMT6
wGcmGOHswpfTmKlYcFhsMIv/zMu65QfjS+TkSP3JgA5Z6IZnjKh0blTxhHfgXPIuiBK2mvmWWdgu
eaf109c+G3YKH9Lsl+HlJw/jYqZp7dZQ0N1jgL02/Hdd3cA4FPZu59u/MfjraF78yzkFuONbOMsy
m5RS7Dcb+i1e1iwf2J83TQngqaC1YCtElO1T43wvBbqTij11OdqutKl0yVfO5AYxl+Onf7CrKbzK
d6kCRVvtFDTrRIG9TZEMocAV/wjwt8NPiJfwjURGDDxNEBl1RWPglzG3q77LAidwCgqlGnONBbkV
pf/40RxmES8Y/W3f8mi89aFzLZoD0/XaVPS+HIY7nirtQI7YSu29V4utsfUi+ZzJ6wIZ0mVcHprw
u1rQ6jX8f1nhZUMGNUXKT6TpMKLfenZGfKNPsfq+R5YPM5O77/W+qie0j+DusNcS2XKY6E1KVZIb
g4tpaB6P+VaqNLe22gCtI31aQdjy3YgQiSJa4kAA+q7qLmoVUQbufNfiT40DYR7hT81wnWB8w5nV
x0SqJtiAcZsvHm5WwkFcabmhAuVhjqcT73pW6vANMpXC/obuBa1zgbiwoW6mkSo69ZB3zT709Vv8
PlA/DtlYr3zrc0PWrEvBGtnZfc7dEgmyAMrxTBaIGeOn4B2hpsEb6m8RZMAZDG9KhZmJ9SyWMIIL
TLFW94E8o2acaBJI4Eknqq6WDBL/Kwipj3NLsbiO7rXfUauea38oPDJny38EeomS2jWy8zHmUnng
f5mPeWC48eutnmLrafh/M4z7IVfpwAWUwBeUvgCexdBtTiOQt4kwLQT4w0cgO/ueTRl5iMJ0ik//
fXApiKvJAdopItD9fhoJChsX22qe9Gmikl/KX2XB13ktJzf8U9pWDn/439KREIHAXybgaxnjFF55
I+ZTPfcNZiFX9HRiy0x0iE+XVhaCcjw6qf6s8GsG9cq0z/2zLALh+yqYpkZ4gc6T40YJv9Bv0o9C
qA4n9HLacS8YnP+4vVkeW3GhcclmSgK0hlBeNygf6iqVkUEzsfYtwKVGkinb7k/WvAmAoKcqmdKz
LaZkvEPnwCqOaFeVdfZTuO5aHMQnK8iAtUEVk5mk1DlYA1rcs+YjQ4gKUkaIawFAItolRmNAveRv
YSz8ETXBK2RvXtT+CmW1diDHlGAU0HU5lM0uy+dzFYit3q0zxYGE5likWGuYdlEwTlSbhUx3SMDK
dOhMZIlScwGB265dzEz4bvRW7V0ildhqJ85ZLOSiFvBYF0e5WwPScudn30dqkJp3MSLrKjAFUSJ/
gH3wTHvbWLqy6JA/C3Gz/LEa8hJm2ztKWnxXSjT1vhN2YbtRZFOvZx9eypVjpfYqm6oR6PhMyNf8
2yuseIh7bXzVQceYT2ZwLcliPa2a5U0f2n8++nQA92npVMEHX8GtUhl71oib78WcAh0agDioQSZl
r0vad3VWIrriwOjhlPpvVsHG+/dAcCPjnzqeBq2rolR28ZPaY4HoXOPkzUN8SaRQnsRK8xDm/yXP
pv/Nyvafnx/MdSDSs4JMLOMgM3ylPxytGl3DcYfktRFsHfhUZnDtTMwSKuMMfCEvqsFVAb2IWOWp
YcccAOnNcV3Hlat74DhTE+2vcDIeSK17N+9fI4AuqeCBVYG9ThM68Ivms7LQ72X5IHNHLUBjpRl8
qA7Fcuz47Q7GY60Bb4q50S2JqU0KPIbOpt71NHDBaZLCQDP3PfB0aDXmkvT3QYsbqvfupm2IqB2U
Dvco/llWgfG5MYTx3RBpBS9SyjTmAbbXmpAE+TgKdKX2S35DPud2pHrSmKo9QgSQSJBIZRuP34eb
VC50YWlrvm4AC8Sk6lg6XeqGpX6FinAnYrmzj9hY5nfXUYE//MZIS9n/ULQC8maaKUxcPSPFWZfZ
meeWbw0BwlchiogbdxGWufiBig5TERoGi+ebno+g8leoJDH1AuYPaZEzN1VdEXnAlBokGo8GJYha
Sg7yIGZUH038xQl6g/U5oiG5e2SP8Xfnovzs7eNuKOO/bTaZUDk8Buko6Ll3RdI+XHUVZselzk1Y
zjHG7PaI0NadTT23hIQWJfP2l1VpMqEdohb2DTGYs20nDGrMX7gjyNVvbM3B7gbe0bz2Go201ihI
FColZxX6gSobVQkfR4C7g708uA4sfUXq6Nzb87Xf31fBWol/GwI7cuQx++yM/pMRqIPw6n9OdwgB
pdsV2gN9DYliotyB1ekzKGzN2WqZieeZV/PITOs3Rmq5vfGR6Stug3qSk/ar5MSMUIWbRFXxMdNP
Ul1g4SH2wqbtsqQcHz8V+Ci3En3YsrPKS6jumFtzFevmV1KTchoTlmqmQnVxovrDDewD5wcP0Vvp
1x5egbFDXfFXdXEPWcchAGi3mLbdU8loPyBgcr9l0elR/qFvSYTCbojG2BxXALa/w7eqhhNGC7Fe
X/wYSR/h3v12JPDeZslifcqva23yvhfSAVKOBKa737QiBDxc0fBG21YYbi5+TyJauY6T4ucRuxYP
aBvaw7RXJXFVgFiqMSFC6Zq0LAuqLmP6/r3sIoF+gyA5dJ8tBw+e0fmpH822bxUhlkhzc07npK8I
VwxQViTqM2ZCdahafoqE8d+ZkhfLhjt9vbLL6Gisj6j7u3M9A6SPwP2A6xlqFhS5KZ5br1QQ07QB
M/bmzvmF27E/f6WsC1dHq/STFOgeYz46hUid5ugGwUYC/U8vuJ8q3JHIdhAEix/yeW3oNBsGbuqe
ejTPdrRQDGKACTCC/f0BsNybTRZeJL5IKqHdPqYtGzE0MmXdKyA4kiFH+z6fNri5UeCI6vhxpW5M
VemrxSjludOYVPYNkegGOjLIYDPGVSu+wPOtsewS2xZqpxXiAEKzkNZFLGODjvq9PonkD0ZcxlR7
smsDNM6V7KMvgpWzmvRLbcg7vKXOfnzBpC3/WGAR/MFTe6CCWfD+GIZSKXx37iwukSMPzCFUsUuj
KDMxmuttJTYiOpyH93kqzH+GLvQ4GGD1OVB4PAa9kibVDv/wT2DH8AUlJ6JbvwjBL031AuwZeClP
85MbH4fOsciySwZMlcou1eZL7y81ikuUgWs0j0ulGZOu1jW87JTGjf7EB6ZeeO+mpcM3zkw6Zs7s
t/LBRVrfS4kHSzMOM4t0Zp2j+DwgNApg14owv2x8RmRk1jpG0I6xxUf+TEy7cd47+wbJgFAJ05ga
445W/9SYrdbopUwKcBH8yC4D1EZwiyF5WvVNxwclO8+Qaqn5ESzFmO6CpVObhDCCJeggfdJMvfS5
JQPnd68BWkoUO4YrNuY3hkPtDR/q0j9AUpR/DhKpdKAqci/7mceE0V5rh7mxHOY7rlQXjhMa96Pg
rqGsRevPr2rNpZYvKAsty6i6ptahOj5FH8FjWceo+71WLsvbinQBlX6r9OcevJ4mNzoJo7PgytWd
w2Ky1Fiju/A6S11EH2Uw0dtGBprf6SnvOvKQn8LLKsgpD+i30CPWJlSPFrVaEWQJaP4s7Igd+RQR
tNwiaAr0/UmCJ+AlHk3cwhHIJECUJ1Aw40TIGBWqs8O6+1LNWU0csZy3EWiF35xDsZdxW9fiiZHF
5xYgJ4wcZpHZ90pablLWe1B9DeM0Rrlc3/+D31rrLNa78CZWvQHiQrm1dCU34o2L4Xa27Kg5mM+n
KpsASAGP4qwA9msxH6JidAQMJTTN7E39tiGluDXMCeZmLIx4eAB8EHfu9/aWIMSl+DF9lG2p4Zu5
FYzw1yPWSsIvH6p0YNLMvjxWKXfG6RoovtUsbK5JlJ0o04FzsBz//Q/Q1SrsJyAdgV7+dSReXEh5
RLZ7yvpKQtjOjWE8TPd2Ojqw2ZmSZmuAn6fxTXWYonPMg6jiqGHHhu2uqZfRx5GohfnJ8lyc68V0
OLnwIm50c95qhiYmhrRHOzyv5q/nHjs658rzQbDs/tyDziXrl28tYZy1mi05Tl4QfUQO2CS0SdAN
9MlyHzNvYbAg/QBjsyrLVoKgIARJ8TmSfbWqePyxumDxEsFQeIgxO3fDsSfo8Lr0qy9mqDJprH8y
iSGG8hGc5J+q4pSHnoMpnngKvluYQW7nvjYNSmbcrY2B0AjSf4k56uEc+zrnmktAuUYBVtirFLEE
z41DGwouXzkFbqWq27NUL+t3JT7C6ic9bS4j52MaHrUUYmhcxgpeMQDCpnzio5Qayv8ykFbIXJJ6
5ht2/jjxOPD8aDKVP9T/rm6J5TgLeJT3ffgQDLheCJKGmzh6VwJORjKANRqRpYTtuJg1npS8pQal
PLeN+474jCtHeJblvWFeWdy+XewUZXUqWOwFRfZOi8oOJnweydlRiibqLyj5eH4IpGfo+wVAv3qb
Gl20Hw9fT55FrvC1ViQpGSGANqCcgFH5jpM89zyAxt3WNLDj4rcSVtgwcMRZ1CddVWyg1fYbFssf
oOO47UV4lOs1BTYEInxyUsqkR4iyYqW01Tu2NEjSgkPftyJcl5mamuBKSPnEYh6pNzZdu4VooCTQ
WireVsKmJLsR7nvvF7HerqAQPnRgE6fJ39J4uxVy54LvtObdUYPosmAQR4BZ9HGx27FnvlABmQuc
IM99PxBr3oIpTAJQ5SBSYUA8nSmuOFUBK9wa4UeBxvGckAy+zoNf7rYd38vb9VQYg4HUgjDWacL4
+Nai6zvnczrZBulHS4D5kdIdWfGwPsz6r0McDEF1uJ2GZuZpT+g3ekr1xN0O9kvyzc57BwBu540H
JC825nsXoXDGVShsCHfdKI08ydIESIlu1SgLgVkc2LX2Ho/c+gnWJtO36RkBPy/L65VMT0ioDR3f
ge/BAn6a4aH3e343Olgi1EhrXwd+orf8BweK7Gc4gFQ2hp1uEAR7pCOQwhuhgGYV9UOVbm1VqYXE
fyRJRK7bFwveoYjxkkBxu5gsN9qnSDDVKRGF8g38trO2zpH2923gqAA8rbFrEsx7up/xfAFQB/XX
na/qz2uAN3Gm+dU+DlOR01N8Nt3qTmzLJZttuIEguBNH81rcftTVjFJDTqSx0+n8oGS953J0M10+
7WvWzZn1ahZ1WPefZgVP5Yf4MEfiL5D3/u8G4w3cGFuVusZTwW0kgo+NpjaQX45PoEW+p8oh3O8L
I9r9haK6rQjbeziw0c6LgILRTfMq7aRT/gBIUUeUtjO9/pnzCysSudlxf2j+MgiXhsfVc9yvMFzq
yhc8ouWVjngyIlE9/gLw4mxakz/4g/zEKD9nzCsm4V4rvsPuThCH/jqpSVBEckn5DmGTA2OFmsLX
zU7VSGumaToPA6Wxay2AyP+avVD2weY35YwxsUYPnBG868g1agwLsBfkCRmY7Pvwa7X0l1WU43lI
EfmXZJs3BR23SQNFlIVdGN/DKi7C4l/km+lXnbBrwZhJJAKwslkTLd8T3DmkMPkpXmBjgPyiP+eS
wzjlCXLn0p5mz98wsB0KKYm+sUUNexPf3qwr7dZ2zkQDMoOIedMDW76wr4Z0a8UvcOK8DJ5/m4MW
JUtLuaSoJQ40XL1Dh3CuDNug6i+vlF7mxnzT0LFdpMGnHpGOd5HV/+DO4tr/Ob8oTXcqtxXHBvwq
Ox0aKH/lGZ+a1XtQY8kB4goHQeiZun7RLqdpW82HzvbWL+sjDagvaKlBVh7zeIKsfSjeJTWS1pps
wj0UoQKQEGfx+zQ8/mfU8Rt/goLJXSdr5VVT9NJ8FmBi6azwm24+9WD0z0kHZGI4vNyyYXnLn5NH
HbxiGKqZEn5cAnh3cDVnU8Sxn8vPMKcs4jiFVs8HdZmnsQ7fB22ESvEXa3MhQFx64kRIOOt1Ycf6
oSMITjhZrBWBqPpiEZo37b5ESMo0lnNAeknt5OmUS5ml3i2ecwNz9a6oLRpyKMuJGQKQUVgAynaG
N1/kdCjajg/udALKvWchqHAEz3EdmQ78+sJJBeXz2fJSGvRpJBPI5dEgLUYWFk5vLOtMq3rqtzbS
zLwszlgunY1yLYJer7Xjr0pIB4OxjzvvNmT6Oq7sLPzDbjlXanxKE4Or/iwxcBNoCMxHuUqFHaRm
xkGyw8CATTYZ4bG53DcHxDlmw/NACEPIWxR6KefqOYGcwQOKyVFAfowGICgMYkcWFsqmEvVKBb34
8U75sM4soFpzgmjfqghamBb31DVu5KtzCZZNw9uNcnOIsDsRJJZ7oG35F6JI4hY8vvNYqvBjOxcd
QYklRg9ci5p73AYCtUMzcWXVZk+A22+U/QzQK3vw6+c7gH3ivaMtM3YB1q6h7J6qToOIJO6pDMAd
LG9UTMKVcOKuzTzmxEY3kHI6ii2xz0lPyV3Yw05YWIMOeCMR5V3XlF/bZQMFsjXEMa8aSjaaUt6C
qdTGtOSPunzTJVrDHHKHVsW/uhLs61L2SFxHC6m1vebmvlF8MvJwS/sMj484QordJh6C0Onq4q0O
sCefKyoz7Y10wL6fOW1KKRRxJN4hxIPY1xYFH1H9U/0ZWvZsJOKYQFtkNXKYetjgpAvuD4Yg3OT8
xtJV8YsjTd6/StPLgSmPDJRj+BlBfoVEawRlpCmNUWV2evP1Cob/n7KK0eEEjIdIopfPS111T5rU
Ppm9MO/lBRp9FopmTRbWUWMW9shzILb81Nre/GNDtDRotDC+FvQQCsO9BzfHePIL61v8RJgZMCei
b4XD/b//elBp1kng4bYIHznWjD1wLYpBLKuQm5+Dw97PkKAPFZSBXXsIoNJw68JxJHFHtgdADxc/
n/uHauMKT1PEsPGfSX0ieZhNJZhAh8exxUrsKdVdK79DKslsFiUR7nCwh4Qfq0RezUJe4RPvYrMV
nN+q9nVAHkuvJyyNStV+58L1VlnXSoVW1cKzq65L+nMBB5zhQ6ZrFvCBwLEku7iCiOTk6cqGcQLf
ZJA3x9DI3Csb/tVD+Gg2cZGSTxXOgOxxEbgMNG5om6fW/+xP2xAGwxxotKM21JMw/oSsR67EVnbO
eS8TRImbIhXCABEVlpkKRgnkig6RoavpEfdh2d65boCwIlCXBEkZ1MPkXKaOjn1AUkTG3ExzcdF1
py8nQl6qDQGL1tYoktyN86+MvyTfJ3NhHK1wgkw1xRNbXjOoxCODvTPeNj12XbvOQ1dGLDbXRU66
ZEMbX7JLW98J/yfgWh7niIsNIcmMxX6KJXOYqS5YJuRCAOwTMIKxdxMNJprVbjx5SRluoDzPO4wZ
Lg+PlkYJdw7J8/fBufcihOF+RnI1285G+LCz6UiT8QD+6HfyTQ3sh2c2d8Oq93pJYy6liA1ajoD/
LnRMbA61W+27P0v+0MvE1lZeCB+8oPDnAmNtrC8j0Fi6Ylamolo6tT5Tj52x8oqLH/FTN0H+NpFr
Iy8R/MUKPjKVU+26mrAxXV3KOyLvwbsETBnQ4CDxW69bFxZYy7Lu6+IZBxzMp6c8gF05eUBRF3wy
wMDoh3ECEZHo7jadd4sIufFrxhRMbzbNur3TSEHy3zu9OUL5w2i+grGeOVIPxsHQLZBN91A6MjeC
PnFTpYnU4JqQAoD57AAAi0pJ4QYBLXySq7l7274yJIV8+LDpRN4+nc/WFowZCF1KduYX39stKLFw
RYFgbfJGbhjquYzWfOPVL7NC41f7dAKYz3GcCn/mo9Ge/jEii6Pe1ylmIWyv6Lc0BWTKAWAPb1Nb
MDAztFVLCjU1lVHA4aA8iu1KTHIz6OLyMANkarih/22uVbstQqV/OAIU/EuyIJTfc3vJ9khDcRbr
EgBAbAXzhmIR9uONT3J2kzcNBeQ6el+ehWF0mmrjXIhmJI36HpJA7QgPxwg0LCgN3xtq4YnYlnqk
EABhHC2Mu2zswvMonMew75u2YSSLIDamG0ppm9tiE8CgITT3/buS+Won5GSXZiIhec+a+fcZjrVO
nFf7hmqP/1ecrHsbs9MkjD2vRu1u4U8DGg5ggGcJz7Zb2csepsMok56Yazmk+Fuv3XWKAEMKNTb7
AohtSPSmBHtts6MP5I5n+PqwMg3FUVLI1CQiodo38IVFhPlH1pfwwh2u5L15FmCiFPIPBDH/CTjJ
x5lGtwoJvUJNHFXZ1sBrygKz2jdh0jO0a7YfilT1hfnVlBSal7S239K61ltfTS1eD4ljDOluqL33
/LXp/qauOOy81K/1XcsUfxd5c8ikfa4aLHYUPNDNBKyzfsu9xdZiR9MupJSVi9OtwIi6OvCRBWbT
I2R1tVJ7bClSg2uPkMSMv9V9WrP4/F/9NCLlNQnuwE/AuuskBzrg+E1ehsNAse3BPi4DiqvMUWfG
X7ynemqah6ngWbwSv3RZHIBmP6Stq8aefP1Tt7SF/Foumo/QnJSDAhxyETdwgOKOaldjiLb/ernJ
ULh0K7YmxjfAZW6XyA3pnqX0YGUxJO1Gvy+ZvHutvuE/JpxvPUGUsgDP0itR7Tn0Md/Zrr29f6TD
o+evfRpT3XfqONHIWJx7RMfxTsxcKgXsVJGDwQQrBUPrYQqE08/fTGRk+gWFEzVEs8ZN812ErRKD
aw43qqpAZxPd/ltxi+BLxFQ27GeCXs79dr+DnhuNTVUopQOQKcVEgHuJTOcixfmrvT9lbY2q3Civ
rtIAPchABgHr3IYHVQtubFO1UXDbyR7Zs2fH2JIrU6CLAGO69bZipiJmiwDt0R6eqUkFC7oD1nN8
IshV+3C42POBB+/cvgXNhVb8TQ11zg9KbKqn1wFIUI7m4W9OOP6DbfooFm1kz85Hcr/qWT4ME3NX
QH9aKr9Qr66KajSwM2t75PxonChlPIgJ2AdhayleQiLLxVNGhzEKgQRNAnh1ZkrUeDB/Bs4DruFi
BtcUbcRm0sk1mOPHy1mbBncHPsl/S2HOpLCJtRCEq44OEqVCb3hqjKP0qNnaulQS700MMlIK2/Z4
jf0BtK69tXUl48VyQAhEXsXmV8mn7420+Xg2JjWrNrvkx3nrHIBMwu+Q1rqSYPMCZ6iLJm5eyvFJ
OeOdd1Q1VQOrpS2u6CnRCQfq+bd1bZhAYmkDQty/elcKu3FVerGv4MT+cOczieu6gE7Zl0TN1L0C
nRXEZflUlS2ihl69CaMnRzVFHoyAkgDFyCrqSoJ2ZATB1pwcF8TgmzOfcauNwgYTeaLiy3xN9big
eJ+A8B908HbOU4Q1IHVUyFbeiFBMjKup+C/spGG1+TOdFUgOMQGrSAFdS8zkz6Mg+iSlazGyWRuh
ojwtsjYKtbeE0/SUBS6ERyd8eWsuuK2KWHkJoQXni54ZCAYNDJDvCIVKOdRJ4VaGlbtCa3J+dCJi
5n9VXFzcuNolqvlgto9mj9khr0JCmO4ztCAzt3dCuM2wfWuOsK5zaII2qLU4YCa/ZVqgfM6ZDkRF
UbGqAJSS9z0bKVrQGVCjTc+VQdPWGWSQBrwf9XEhyvZvPry64wAhCz4WBy2055fR19lq2cLeYrmi
DlUSmlfANVAVohQPW7xSh2/QWpCe7KzfKzO9IiMQn6lV33peVr2mk07kDopOqzHZrLfLu1OMlScY
7SOFTKsBx/Eh9jTJ/tgNb5qpGU7hA+R3kYCyjr8oNJndt91hjFqq+Qdjig5AdLMEMoxTRJ84ybFy
nQmNynrjatoukcE7bxvVUwu62O5tkqWmxdX2CDDtCmczlD/GcLQIi/ObYxNKAA+ghtWxc/NMJwU2
eIOOGa6EEU9mgy9YwKDuG5RrSyMME1Pk5bHEJ9L0X31N47r8c0zfjkK0KxrLwgdAHviIitF7n00l
76tp+UG8Zj8KHoWaz/DZJbop+6KyhQymVztnpBn85EZwCZbR1UC2eyKz9kXRZEQv1hfyzVQti6w2
ECRPr6fS2c1bel3QwhdWZ6swsKfjB6pTiYVk8o6LQEWoOy1xlro28sj7jzmmrpOA/LJBrDjuCeBR
O/hsdcr87LdtYgGOb6APW4j45YwErbd8nw/X7KmceunA+ES1JHT6p9KPM+Qt/4kwTwLJAIo6j41z
dot48FiBixLSzV4CEGO4zxI1+FaOrK0n5/DgHWoXrDG9zWgFVA62AnGXAaRjG8pOY4R10iCI/fTb
LG8C1K1mI5NuslZ2VveGOMCAvL3mkP8UAHE5plCUos/KTzWemd2LwazmDqppi5jy+6Cnzab8KdJK
uNp9QdYsvkHkJdBjYwYoL7V66cL0xmadKlV607eYLhe9np4jq353xVt5ygS0/nYikg7aHXK0vQsw
ktjlS5Vo4HVLZ6/5jrYOJWx7bqBaV14Gj3/ws7GqTcmtbv9rKYO+R74Ijd+UaqFIdogWQrLxX/wC
MUy7ea+/oY44JI/RyrAfvEUPFXCpfE+58D1fm4dGHmEy2EP3MH18m1p8bCWWQ8FWdPWh2Qudv7tQ
QvfHFEzvJBNFqTP0YqukrOikkgAXvQYrIqGWh8bmBrAtS3SWSIIjaJZ7442qxS2w3M7z+XrYztOT
pWrcnwGYx//mMEdYcYjjQiFwrJRfKvgep5+FhOwmZE3fz6YXf7K/nJD/oBk0w4pBH+YxpWyGM+Gp
fiZNHlHADKkphQ0C9esJQQ5kjp1TW6M0Nyyc8lAsp93rSmN78/ANSVLUvSPLCC/xWUZOb7WtKZ7P
xpoh0gVaDJhZKtQmwV4jfH4QhTzCVHibzVkay6cKoCNKlEpl41IhgZSSSWZlEyTzFTWw642ObPWD
aNQWeU6Gae2Tt5GW41tdnRedy1oEZTlgEJBSwiGUmw1rE+OaYGaqCEAoPbkG2558I0ssyf/k5DZ0
tdmQ0SNby7k0jjC7EmkAJq8hT2bjuvmmUQIuyyzgOzvhiUFbxiKUXPpnT3B8zvmvhMBl8i+cLiWG
lM897TUkSZUWqwjXEkJ+b03iGqtMrkOdsuPeYTLQP1xKJhS0X2rHYukAYs4Y/82zcYJyEeilH6nk
QilIqHxzZIFxZUiSyFpX1AYfcVjkIR6QyLHxABf5syPVjJPAOdomuUhBHqhf4B9DzA+jyI2irjh6
9Aq694u4S8oOyY/ZgXL1jl2ipZ1zqGeCk+RmybA0oiQGBjOE9bl5LzyoKEcwnf4RMOXvDRou5f08
Olha8claxAvXtB2n4/ghi+8pa1ho68Hcr+0UjDGro6tafGGwRx/adJnsnCiTIhMDQCj3BLkBkDQt
xu4vPVbLFFXlOWHHt6DmTWrH16sHTYlX0COsK+UEVfMS5mVuIuEqxZySYerH0PiYCFrUO2lZ1Lnx
aiQm1BpUzzOwcuwalyu481/OzAgA7oINH9ngsA4FfY+O31pl1mfs+KCx9IxsHc50+SKoSlRwBBGt
bncH6PM+RuUf0CW/ah7Rcx2pV3mxfF5R78K9uw3yUawDY0HLywpxXXfvQnYFR/E9SARYZcmk89wq
9W8EJ9Xs2rOWQF5fe4Mhqe35aSilPsBLeYz2vu3QlwwIiKoiKosUkQBs/UulG1jj4ZEJtHkG3RAM
MvHb4s4QKlCrJhdAe27gLmaZ+NxGBWTA4o784qKRbaeitUGnS2FJ5Rj/+uuhlLZkVWPpD1gsjcfa
Kr93l9fZW1cw8ug1I8DzOe9hvdwdOCPtSFVRoSholfrm2GgbnIBixYLCrKiOU453c16gO4jdfiv2
4mX1g72oPYPTNj8qKQidIeKPQSFJhLD6xsj8ySY5yi4N4cpYJ1TQl6UHZYgiDB12SY+Kr5CgaW4P
ceoh1Y85ihVUqjfoALXrLl/A5r/OdgLQybk8c8b3Yt6ULT0JDjkjf+NeLwKHdGlZOY7hPIWXFEc/
9Rsx1k3y7IgNkBQUNHMmCefQ8yGiK/UU/jGz0m2vJSzvM0d7VGU/kjtTSzBCVBtH/DxHL26XsbEj
IXOkX+UZyNsTp4eVXb44R0ka3K8tFYDZ34HvxqPJzN08bsE9h68fFUdnbBVgs/PuMmFRxouOjPkY
Dk9aAGgJMZKauicY4BkWYmUenNjPA5DYoJaOmd64hGUtIMSe/eK7hvnsTgoLHk/Iv+5nJe4SE2k8
vYS1NhSD24AZTpmYDjdpQeekplg/D1npi0fcl+GAbclM7iWqEJoPX0dOaFSuCCoN91SNrDsUjSdw
8az8rccQc38H8RmpJ5KfOOIC7ohGu6A5U4hIMaExsCuntN4fCNBjc3rYmjIA6Z8KQGyDCdnq2Rmh
XLeb6Jcw1k4PVK6L3M+nDjFVeJciOIp/JqRuof1LVHto0Zc0TuuFsRA2qfgGrLYPrrtZRHdXVL5M
5PrKXpieAGzf+zVwycv0EfIQ0chGpEGJLLAelIyM+rov04e4UXih84C9GBkt+dCyK+L3wO75TVv0
wuCC6HpNe5CO8NFJ1pnjHhU4K0o3P6AOPNturltwqNHL7Ezg+A2Ab5ic2Eye1+4a+VBMiF0TuNkb
wmmzX8c5nYaTSS42slVkmdsRZRJIy1fpNvv4EO0UySLoVA6DA9LCmJdnNkpHleyVY3St5yvuW2sz
Mlwt3K9emWDoeV+1x5+z3Zcj1mhH1AXccHE9pYzfj3jLmL3N8QsRVLgZtqUYaoGx4/hYetH8fUC7
mNLZ91wQeywbAg8Mgikn8sRlfaAKJSnHvtFpn1UtphnuLrz7xhO3v9Ku6uphFXBIDnWZlX++C7wW
5tl/KgvEAXAf9Hb9m46QbuLO4UlJB8nAVcl5QyPLnYtMjK1GYW83JSAi6PddVbMXdxwFRz1n9JkC
U5q664QwwxcSrBxmtUu9QGdHW/NNf4VeU3tZwcQEbP54rgHT++WgeDVIWKLVfeLDEcqDLfxh7aQ3
35bTIpvl4qF56LsDRHE26NXDDe0dqZj/tRikWpRfOmd0/ziyY/paz36cKjnDfJMP4TaG/8sDCQjg
35cw7fZCzTyGVShwfXcwCniNLFftr3f/toeQl7LRjFLv0RFe3YUKHJLG0fLqzYFMX8cAHclen1oI
gg/74P99rXE5JO6Kwt9t9XW51bVDAkQGiMqPDAoEW83r5RH0q7epUR5qxdcSHuL3vQ6H/I9v7A5f
FH+CQJ9MVlNatrhN27zM9IrX1NQJ0e1frRPnsjEtiHf6+2cN1ZUmRbP9fh7NSmUN4ffcUOnw7iiV
JS45cD1nlyrSL95/MEB5T0aT1dPUYaZ/kG65bWwv8+7d9h1mP+LGa8gZACZW9YQ8E6Ebn9QLv9Qt
oZvVncMcuqQ8MO1souW5To4A+EEYxAnLZg/AdcnyDzFEio/8yhmLRQSOKcaKQMaV3lwkhSDkvMS2
Vz9/APdW64fEQEqe8dYg6iXwFUlWzsllfvpZP01DLh19+kR6x8vU0wmZl6RMLzexs/heJ53M1aNV
3xKijdIbq05j7Z1AtIa0jzK+qQfxG/Li+HubELlfenT+4wrAyEnt9SpBwFwcFc6XzPhxa5PZ2v4B
F5dkFgCzD2NwBvq9fNS8zHt3PfssviN++0hSDRj76SsfCMWaRJQO1zijBNnkFE8jmmhddAK949YP
zLNp4UNnNwQ9n9azkaPawldj0+8ZUSI/yw3sa3goYst/Bl65ANyM83CfSI1CESABrNQJqEupyt2f
JU0v4KaoPRzLxGvPcmhdya+UxQJG8cKXb2N1oy9ESo9jQgOYsieYgn68dk1Qy44sHLL0a7Pe/xJq
Ho0QUKs9E3z51AiF6+d54/rlRCptpoNYd9+Tc5Y03dTZLGfWThqq3Yw753cPfEtxSGhhzXdxtPa2
mXE4lx+RCRY3lBqy8lQA5zSblHiTFicWTBULLAwdf1EbWjDc1IoF6mc+sOpYTJLiKQeCE0vc9GIU
3C8GCwiFaTk2Gq7395cDSL/BVzkuJJ85gQd7UUlFtj7hG1F1cPYecPJaiEBhcbffSHE1kno/Lc4j
dj08ck9uIGgY8eK9+qHwsUWBFwt6HFXwrP9F06r8fzh/QiUQOW4p+GWkbShk9AeiP8S/NHg0lLxf
qF8W+WCPeX51zYEKmpG1cDl0YzDookULd5cyBOpEdf8mR2L8NJKyO8DyESVc+grXLDyXXNy0pgAn
Lwdq8ub+WWUWSQEelht2o5Z2t3aqJEjBwPi4Ay41DSRIXrfL6nOJY8g4RpjLl7vrbUALcn6iOb7s
qp4bLcrfyLKP7rAXvlAOfJKHTzehGZBnqL0tC0E4b8KzFQtV3wnPpxe8tqrSt8w8Nf14bZNe5vnc
E496FZhEq4OiMSkxaXnwNvdGWqDui39fig/FE8A9ibmOls41xafKl5lr2rypNCprsGRStCGv9eS0
ITFFnTEg5Vv4nT1lUy9OJYiRD1PLZYwkTI3DgsnaSDRfvP6OnA+RMjEEcScDOmhOIHk+zCeA6ofJ
sf5y+oarJJ6XY0Cbgeue3bdBgLrfIkOl9NAB1jN7G2ekXP207KENZlwaY51aDwKfm2U1wHI9Fv3a
CLklXKACzsi0kMBdQqFMGwmkGBArP9gg26WR8qK0JwMH+Ho6IqXWGFKb6b6KXNC30yjImsL0DsR4
Cz3LDQCGKds5B7+pctz7UoWpKfMLlADCWgPErSSyuEaCW1KA+4sj65NHKSUA7xm51NN+73iwdlDL
6ypSsJGlMD/bRjLGcnbjyNkFPJ637r1Zaaxr3sz6Cfr9PS1TZ56zOFbjBAkWMyGJtHSHjcwdQg03
LSBb/GCFxp4yUM/0KKptAQz25CWtfxGm8vWfr8+8ty/6uGpXal+Tl803Gw2uzjPfU9a5LWUnbw65
9pvEPAZJWak4iVS71fMhyPXQuNW344ZMHGGb6d+qMAhfGrabb9p1XmJyXDOJy2oFT3FBkiTOllBu
Q4ts4N2KZ5oMQDDZ/bDKxutRqxwVvV40B9tKnsT/JCZp2vfb8J9aFwHMPgUNIxjvTK/uMUm6sH3S
m2wci9qEDlEohnnxH7NQ9SWOdv2DQu6O8wn31mur0JfdsxFFlPIcmN+ac5YTKrB9qyNYPpcnEvDK
uDSxS5bC+xPA4qu/zQBMInEHiCrbMatfK0muMY5mD/2zrYvlYY66N1S93jmsAGV5Sov5Qy2z5zk7
drYM9dqtU7GwyPzn9b8C14UwRlQx2//Mfb9V8YiM/3fy+oLaKloMGscIYVL0Vz0bnVmgA7QK4jB5
B95nS69/er2hcYXIcC9+u4m8Jno6fjwzLaahX6eAjGX89UNjV0fxt/J/QQ+eT+Hr3txKtQhi8bqp
ulbhjftP8YJvaWobZysrNjuSfa9NxXeU+YbLg/V5qxfraj4Evmr+Yi+YLkXXtzIiHtd16Qgc7BE0
TyXOLbyW2EiU9QiKuTZ9DA3Hz/FPb3ak3NnTrIFaTVjhYXbqbmJP4HtKa4IG7fFj6Dx0IMWmICw7
6uUyHt3DKNkbmoYYf2Rk4N5+KZ9RrRS9aEEkaHTx2annhoI76Mugn/lfkXwy7zBnK/mP4AsAU80f
wvM44a5yQ6ovaL2FZvJcKiXTC9eK3d7iSejUSLWLXbo4jhFFWcomzRrrLcb5pTWC4fIiowF7snHG
k3DhqdRgLhaj0PR2L6yDV086o30UhPs3TA+wQZrp7ToV16rbDEZg3fgRmu1F6RqzH3CLMHOZU7fJ
GpiRTpfwLaAeHK6PvmxLEPJpNsMAiNcSODX7APX9gUps5AObr8ycECxNRmMciC+GqbAtqvy5RSvD
tUDC1wPYHCK7MMkrT5NwvrGDr1faddpYTn33pkhD3TkHjpURLQIjTMJC5TbnGGnqllUQVph3Awer
oUVQwV20VnBIfREeaMS5wwFUJ8rFryy7oqzZpLttS8yo5PddYOijW0GojZPy1tG+Q0c4fy4iBav/
MGN/grfq6b9Xw/970GANxkwoVOt1PlNqM9n9O02aXiJ/DIdyPN/5yfEbG2NLg3PK7OMlHES/oCw5
AEa8aDZvUy368Sh9rIPCclcFIsNBZ01fK7nFuAO1AZDKGalKzWIIgl12J0qnpYTccf6ksg5Z9fPb
AlZlmr6CJsVEdB8r72aXnqnnIyxeQO0mEFqL7YUoGZziG+JKoksWUSxGrgBK4LpLhp7A8sDNh0TI
CBmLSI+uyEdsSGkV1PfEe+ZOcMFehSrLi6wg93D7EBa6/6kdAy0ozq5Wd6x0Wj/xxxXH+sYClhti
LfhkPR7Z5tVjTk/QcTRCFlbbb0oRff8eaSEvH3yRG3Ln97ojYMo85AKzCF8hkHirsG73mducRQT6
Bd4AA8pYZ3m27C+lhHmRhmkgFLj9ZwkIw4z3dE7yiFOyC/NleUH2Hca9NTf4NqPH4LZit767OA2p
81oytluyJTaoxxxE5+xoCIuogbxdppxXog8ugc8h9nlexBmPU+WGc2ZfHkK65o21vAFk4p+eUcfY
WFg1zjNN/urFHtGHGs4EnrDlD/DecX1I0UeGby27VdCEBEIJ8+9hfRTrrsDcpNP75+pQVJKckslj
K1jDE5W1dXfamuMvvN33uI48GrFnlYqAGMuX7lCpdxk+lPrC5wzn3ipgAyB9eZFgOURXNGI3A/Fm
V+gpFvQbtx1noZOmLV/5r7vtA/Cu1dquWMBYwdlBiDL4bRakR/HyZuX2Uq4SPeMnaWxgY1ngY1Fn
fqKK5oDYecITB1PO1xwTLS9ce0/ddBiBE2/Rm9RUqKnCoX9keT07rN97WOless1QXQfyZBN9bJVM
/9jxlTbjECzyFt3Mg7ga3NW/wvNl3CtsnUjyOB4wMPlPabq8xtf4wI2sKC/vRZeUbCVWDTmckfxO
6QOJrJ3XpIcFJSHZx0n8Lf/ZYR/Hozj6M+X/TtWtkGha0l8wpipbX1/rF2NU7BbiCN0nAzXImQo6
xlAG7o+vNMkPcFbzNx9KPrshdfhQLy/HK5hmgPb+vbqoY8vzKKssTogtafwYLHHTlSgxR1/GbYQm
38fvLs3lvIjHrOcVy8hXW9G8T6KtRm+UruWnVl9Gh6GHGBCISSQSZ6XsjjYz/LZQyOFylStlk1wy
OAKBHxbs9dxkGL0LEitUqehrTk/7OJHMvAia9/fLMcvsKv3Uiud8wb2TgcnhKxOhXZQlB8urcOTk
jkQheWxPMJdrkwhC4qFQeAYTZIanFDYQi23bWmbhWmSE+UUTQIdKIpTvhPmlyy5p7I+00ZNngtoI
x9Wzv3Ve+MtbuLKINd3KWi3wobFDU2uKKH3nvpyUPS/IVqMgSc1QAfC8FlPEQUIGxCmiBWzEs8rp
GNbnfJcPTb8X4i1JIp29vdVVZznGHjm5r6xu5hPXhkTxG1a7GFbZURp6EN/4OaSD6Yt10AA1i40e
H8Y3P1M5GVFW56lfq3jiv9YikOoGMWYrEQW3ZMYOfU/MTlgrIQHTkrt4DpJB00FpkboyinHMOS+u
JGcKPCK9Is1XETCTx+ZoYIiHAeNrHj3+zIdm5NRIEwsF9sXhY83sxCUbG25KRNjILft/YK1AJJzf
LimaZDsDhX932sI61KdSTSVaHAUD1N1V+nvtZXFdVo9/tXO7M2Vm3H7J+JJYjdhILIQTsp2EtSpC
/JmjWy/huH+6NOyLSnr0RV0Yb62D1lmZrgQyIwbC+YAWb/pN+iOQr01ypcykZdG550pBcBS77qKJ
5HqWG8CtJqsgvKGVeXpghsigOboBNu5zNxdIZyHh2R4yOkxNBKE6iSJF3t/QwihHEA1J+Qvh/dPL
UZ2uv0JRxFt86ESevoVVmxCqFqSgU0oc3VmIDOrhkFOzJskl5ytILFlYOMgNBDiIq6Gbjr5Cm8Kv
zNw7EixNxpvQ4leRm5TfQGK1NNm6BeaVCXtOSOPtgOgqhgNl14TX93GPRhLKH2+XXMoYK8GpCZso
TUzBjtgU4KQdQKicnua9ucwIxGp+IN6JV8lq5HtxVAQFEdA1/vH5yDGNQNUSWPxK8UMiw+i61mbB
KBoucRFY/bRD6Wig1/l39maOnFMbNkt1+cKaQVPhXbXLJiIu5tUxpdgmauu13WzxBLfAq44gVHyo
ggl2wEvj86BiEKBgMKsMCldig6GgJ2B0R7NT4g6MNz5TPeSWkvwzYxRg6Xg5cZVKaihyvIouhkWk
Nl5m8NgN+93WQkIBuqoClzQs9iOASln1Dj6CSDqJPTgaxrcqoqPe7oXjpS5Tbz7boimjiarxiPqO
cLIHAYzKeIUhZhkQyPYEsAyn1ee0zvuPe7L8eAod8Wn5pIs3XdL22PGmZ25PNncY1hHLbF8+owHY
jem1dLTGfVC0Y24BKbWW9BAovWg1/ME5lAtiLEfobJ1PJ9Prys4XH/RKSU7Y4N7DTqVpCcufBQiM
OXegJ6mN8P9q67VUkhOS27M1/NpigWdDs8qnY3p+ZlCaXOUiNb7IDblLThWVtkEpnTFqT1Ndvm6t
z66p4N8C5HdRH6usvS54rFNoPfITRL2RUgMeDu0m2/jXEBEDbXM04qLgC58NkZ2PZA7uGyFb2TQI
G6lF4nmIPAfWBzX+J0d42Ox9f08oSk5JEzD2VI7OXtNbVqnwn18HNY/p7ixIrq7uVjCbKaiWmNGI
JFX0ZH+Nkz1rVHG5TviYO9CmtYFodTTzLW8B+Uo202JpdUVE0pB5zDD5qUhJULvFAD0hDM627KQU
YCtoVhF7ObDh+VWJP+xWUX1FuHYfs62TuQtdVU4844Itsd89IsPKRMqzU0Pf0lAy01iI47qd5X3y
/9hND+ga1oB0R+wRWR95x5Z7wj91riF4O5s6cwgNnECmmIePr8t5wos8rK5J2TD1icQ7yC0w9DAx
Z057T1gE9vm+6b4Z6/1PkezlfCPy3q19X16ojn7+BKtbvJCssaBvvj9nEjmXVv3ZH3Us54glhe5X
YKlQvl6bzKbcAp9NZdBRV7niqbWuxBRWBiXdAqb7KDXz1vXlkuEcBKcrNtsV3/0kTkuthuD+LYgg
fXrNR2km79UwEuNxlOf4AH9swhpm16cQ38VoUVU33vrq+ZNHQrF2wR73UgkxKoGXwQJ4LT1l5mcn
9zppM/ZTQHup8zW/eYAL4dCtpQH5lnMEpMJIuTH8hPfgJhgdF9M7P/tDyg71vrMA/nIAMW/qbHFb
PdmrRcXCQnFmbBcYLvx1ybvJ6iUc7s4HY8TDH3HolwiUjhoyb0mpNt1B4mBAFz7m4nHyQe7d6O0M
7A2x/DDJ77T0RGd2tUKLsv/G1sluU0RiaR10x/oWrGGJkKO6yQY9M3JTcGha80P5B/EG08yqy3aH
fgl8EBu3KLrFKGwCc3+2bIG18uMPe7fnH/iKd852iNtkQ1JDz72VgO8SU4I97MxtwEWuRTBMcrR+
gjRvPtpmsagPvoWNE1EyvpyCMkVfC7SxNl3W6jIYdAOTwcUwswNmRLpjv+kQnmWMoB66L5dUqoFT
WWVRzxLKLVK1gPiIJhZRiNoHWSM6FKmWa9EJf5Vtp/b1t6DL0ZEsiMkuH7KZXLYS/j9kV1yHIGBe
I+GbkwcQF97K7/HwiWqgj9+lgAtAxLM70XgV5Lgm/MzOHaGUhOexQJqlxAh15sH8O5tiN+a96sLS
O6hZvFRN2hGSt4W2O9xLRRkkafIVt2PMvtAYkBcSf/ytdjQNrg0KpCOOKLQ8XXVqRRHfauA1Mjp7
PYu01Mrh+Llvb6yz1iu2HidUyx6t1en8YABhhIgiXRMFJHE7vHe1+ixsKNzdtRmorFlQlEiqQXkY
qFf3vpWHwC13Hxztrgiw4Dny4+4SUkjpzft1lyc76KIm2s+hhzWApXUMVlG9Oc4fqLj3lu742XKS
DhgyGvvZ4RhUyUnvf5By0RyJxquO2yic8rIROV2L1iCD1khsnqo34G294u2zgmZlmsPZVanA7Ked
fn9TXnLzYlWkSqGQuVpaGerK1joY1Oq3wcDuQnLdE8BiOrZH9u+jCKxmTdPZiZADrDy6YaAwABXd
HF+gDDGRlTWkOi+iKmSdVAW+WYADhjgDLusbiLvrfMFKjTEmCuuwGm77gA9ppAdCE1OtSvZA9ral
l/tVvY+xhc5XhPREhsPERw5Fuu/ixI/O+ScAklRw2R+Oc8XJyZQHodPme+pkGD8XNyNZuP79aEXo
M6jzIZ1bN3k9G853iKc6M3F08FQQWaI0ptDTuDc1dvnb71nFky3Z3QEyGdKqcemvHUvANFgWjkR0
j1NWcKU2Uq9x9nrs4XyeqFH64OtKA71DCCY9g/QcIvF+FWIBtwLJwIoeR2qotatu4I7mQ2YpgMnZ
/04PWdazS0AxjxZ022U7U0gjV56mMijnTDzO5z8ZDXi+5ETtPsIY91Gku5fiuOborS6zz2MirBGu
tADGeBt+mDhC8p1EfaN0+ZwXXJWBs99cqhg/CrdnZjIrBrWAK41VoS2v7trfLhEgRWoEah6Sw9b1
5M+qci9ZnHUC1D4cW+VIR7aelw2nIOCostvatFPJaKYFsY5vPwXgrByHc+v36dMnoBGN81a+1hbL
ZEVJ9n1dwAva7sIVgllH4vsCXQzDUwZ5XsIbJdT78WqjMKPHNMP3EAvNzyHaVwA0vJUZeFuJ8AXv
MM/AVZ0Bnt2++MljVaeB40jDkFPoo5cXLOji+2FpiEgoUchS+oDSKV36ov8wYJ/QPZJ+oGWwUtNH
iehnjZvsiDs7A3GPf2mXHw+NvUZINc8CcD7KM9k/OKKBVt9kCtjOcT5+6GFcZlhR5qD/YXr1JWzN
QM0las7OYqWbLvnybfe4LBhNVhtfBI9Z65pXLIfJC8rboTMk0A0GRy60dgCxMYgBTI/zzRO6/0Uk
clBKcE3sJFMHte5McelkoXDPNEbt3ex9Q8F0FHKwfkhTuZrxlaE+OtV/jLNxHf/qM4TN29EUmlDt
dxQJHDbkAAomzXcJfTysVU15n9EhnzHVZMsq/PHSkseHwNdPC6mqCvUhy+p2XyyzlqGbw+J3WFEH
7Bj0ibzN/6oYfLJaMH0EWeKMd+nlMgSPlqvZQx6hPxumf4EPJknEGWL8rVUDUwA+/3/cL6u/mBdG
v8w+IxOt41+MP6CFFs9yB65QPFLMN00m1rgA6pRHLNo3dkmOZWfKwpcRJv+2kCgjnGni3b4tbLuv
gz80ybtA1aQN8b5Bh2b4Woa9xVwznuAy6oDYWp4noj8cBeih8hN6cB0An8zVntlE4MwdxyrkO6VE
CqODenwRwGVEDT83yeSU5kJB0b3LiXFUb8nJ2nkL0Bji7Z9XtLtCor7JQOczmP2e87VOD7bojgpN
MO4tnyTCB6wwN2mtUqpLl700AYf2TIpf3D+PEvcEamxmei3QUV/BSyqLO93mvWEbT1PAIClt8jfh
TdAStdk9gxXQI1l7TMVlE77oHqH5CoKfEVAffGf5bMT35l7TQ1skLFx+TZmhdYJB59n1mPNkvJ3N
bUmAeFoTFZLpjHpb7ivk3pm0Zw/ERXumUJ58R6Wdk2SEKDu19eie6rbsE6PTFy81MzauI3AfPEyx
eBzHZ9X0ChQ344T3DOwq1nurZ7E+fxQeQ0kl0Jss9h51/mQFE/GiC1KKBhaZoxO/O+YtPfLU/jgJ
t9pnOjSktagXymbzsL1wDDfPcF1EzXXLFOHWDE0yfP2+qlmjPqDGtVDrk+gmYE8vknXwARdsy57D
qJYGPnl6WWbzyug95pHcjsrkQ9Jwkk9qesQlOnSfujJYZFPUoPXV0UM4Z1Zqiu6vJC0f5Vzh+aFN
f/uEOlPJuwQLreRpQB3eucDbPSIp/E9saixfzEBy5LuN0v1TMGV92kSVJ+xX61fS9nZgOJ7XIiPC
K7e8gFPpMH2aUcB5DG8aXWOVcCYH15n6n+uZUR07GVPMwoTjtIelDN5ADCK9lP9S5Gm4RA7wYgdB
3wUfm4KBMVSwP0LYRMOc4ReuyYkwWzGCKxLOVohrIT7lRdFqoq0fveHSuGf7UDoWoR0/qjWQJwMZ
n9gwjdyf+rADr2Z0SqaRfjcFxwk6P674FMLZ4LXkWIVjYR+n6VDmV2aXeJaTLMdpWWnGdKMTfMgZ
aJBkts9cMst3MUoiKgkuasIUInpCV/Z9mNAzHTmpPa9demDS8I5JSRGwLGJDRyOEvtQjM5CUOi0G
B/bWMPaRkny8mWGofNtpzQSi9hLHBg6B8WhYyMHmNgLAo3844EEvuyQA22/OwlEJGOXWPz06Bdgn
HFGVBWTcPiba8XD+LrTWx/pnd7kA0Tw30ri0NJm0dfdEpBffA/I0sd+JmIvMch58cRDlYWjC17/A
WE2ZgKf/irjQhi0kIKprrlCFaMi/IDbyZZZu6PWEEXHviHJrVN/qWslpIHGPQontYopuABfTC6ye
j/ZpYLl4VauI+r+IbohBVgEnKUzurcUYD24Fyy8BYmq5E8hec3e0eAi3xnvGEw24t4Pmi787+s9h
j5v36Wm1C9UBAH+Gb+18o4k9ZPOcqtqo0+sqPd3XSIl22PiobJ9urYLY4rsF8phI2nLc7ZHtxz8n
HJ75zhu4TvCJhygHHMBBB3IhKau5MofiMvmOqAW/sls1B32Dm6buq1G+YZ8/wagLgQc8c11pZ9QK
gkWh6U2WKvrPnE680I57PD9AGf7zV8idcq7/yu5IajpRWlJL5ha3wBvVQg5XcXoJfhv3sz1s10QL
161sYTQzz0Lxg7EUGCf8i6NR47suriTmwNKMa0s4MYizcOaIMOrKoTRm5+rOYW4dUlCwBD1c/roI
zVZZI0rWv2lNkyG4ARjji1N+4X1HDqe6D/2+VyENIkrMtcyI1M715wbFzL4rzsQ+yBX140zhfJKZ
fn628zZt4LhVlbzzQtfzRCyNYInrzAJpNqOzyYQ4gOpEdvusD2vQx8Y2cDzyH8BwZRMENg+lQE61
xuS4n2F/or9B2XAcTDhD5H7lhqX8mBF9EZxts92XKoeAFJgjV5tPmSoIdJJdIr8lH/LnCfoNLYiM
CcLWo5yP0ViJWx+SwZB5F85FTDHngYcqAGTyiTch0ygzCxVxRAfl91/nreWke/1TLxouPLKeg4x7
PsRgqB0TSxFqnc5hhv0gocRIc1uapbacN9DgDnTr47uFAFM5O2W4r9iRDy6MnaB2dUfJhiKgFZG9
GEwbHwJ92bm0SyqA1Q2YE/O1SVStr8TZ+H7Wcy6KPynCPQp5oX6TywW4jwYKTVJWQf2kihhNVHkd
tks1oBRi5e4sp5M2oUF+zce7A87l3KPBqUsSRUu5BD4os3RI1WGUDBALDNfQiRVtRCg6kMmsv6ao
QHGgZmAT95TyFpUAaMkrHdFT2oy1WFEuYW8C7iI3zo+rWTB1EYCFfCTgmEWIwk45ZGbighng79nr
A6oDhjhlsdaEdr9cZ6fo4AXKT4FL5XSyotgozvkqM22K3nYpjQ/B0BS5ujjBXH8J4U0f6c5iDOVK
7VU2/IHzO7mHRH+jROnp7ZarK7OITXraVnG85UkVX61Jt5L3OHp5Kp2W36+4SNvZsknfg2+SndKF
fMXLVSmw6aN8tQdLeBV2JXif5ValyRoMZHPCbxZv9+Xbbkpav/UB3Ksn61ijgdVusu/4d8cwP327
nHdux+gsTVJpmSsyh7pNlayDwOwyz43j55RpHUjjBnCdDy9/xlIiO/9zI9EoysHWzocq5VhXmzeZ
y6wpANBTINy4n6rob9I7Oz8SCnrXhzoLRia6bz3b3Ub7YEwqZnhjUcSt+Z1qr1hGLQd1a1Tynr5o
Ep4Jd6VOC+L63rWOqCbs4wah4twALSom1EoHvE840XBFAfhqbJYAPOTV/TTQWO4PgzIDz+rICkH7
D+wwULRo/9hfjxsUDeyUWXze9bKzBvTSSJ3hWeibaPkxkCuBgM9n9JocgRRpTdS4D9WrCt6wdGVJ
hzsu4CxLUlXgSvjbrFvbfKcn4keuzcwbcSkgeSljG7xXS2NyEM2WDyzp11OYJjjqbkq+ZmgBJNIB
yr+VxSbNBDNpogYlR9mWQ66Oqx21mNMigb8vFRjM1EOjKyZM5x0w3W+4+tSB67VTzSAgu9jIN2Lp
YccOPUgCQts7r9TUGOO1pNn8vYuv2O8m4W1no8wMGwwyhRkiuU3Zswu+ViyLBxeUv8WOv8jQ0LLh
IcX9JXz/pQPGXDA+Pa/MZw95JxRXMJ1QYMQeLa2SfCdFDZLaAeAxT73OptZUmz3BqH+lLK5BVJIr
356cNfzkIUk1Vl6R93vTjbRQzB2i+6yVEj/WhsHTDf54on5B7duZ1f36EDWDuEOVy3ZhvGQPYQ3q
X+2R+RyL5L4UN/kfQ5HcbJlhbOdE1KsHvzNqXKWClZIgAahbaITV0z92M1txD3CqTs2uMI7tviV7
+jPaBcZibboGPwsmscqeLtwzgDt2xP1+eigY0yHthStHODDg9ggR4JIczUZzkjoHYyprS9x2xf9z
2U7ngNqm/MDuwuDbc5jz0H2DfYN8bcfpaxoP6PFUahAMYaBFEJrF0IfX3iaBAmYJue1THSFTryVh
lpV4WPRvV0Aw/zQdG2AfBjD8tTX967KDBULU/3myVcrBlj46xP+PS0ved/yZqFNsWSP/E1EtlHcU
FWYB3ZlycEqBTGZw+GSdVPc83S1MWd14MySIcTPZs16hOcR0xsm0Q9nfMooFK5P5HAOHJ/yTnfzb
etw0W81Z9oR41fwaniKY+704lso294XYcIeWiLZ5MACzt7IYUl5VJdvXLsTDHjKc66MwG7cSg1cS
p/NGwt1WcCSle/DTpiX9AjsVTKNSl9krc2+6XcTgfUJOCU1d7Mz8Ws+a0y9gVLOXwbC1T3YCon6d
VGFJYDYjSuLQcJCUmnQYd8CRuNN4VMez7ZTkUQH3iWn6hAIPl+hKSeplh4Y+drqLuoTGEBARQsgV
6RgE3k2c30C0T46HfYIEUZ428VKoW+LACrjy5haOX9qzzMHpIBsI9lRh6KUKzpj1fhFoZ4PUljSs
p7O3soYjltJGm8whK85M+35FyvPkx1zX14ApC950bHmagiWrqLBeZQGwct6o2u1EjqeY5OKYT8KQ
dJYmvvoybQyXb20M8IA1IYVP1YC6WCp7wVBir+0A9cQUBdUAGa2YxZX81XChYJKS1dAlEfaWCvpT
w6oqbEI+AbhpTkApNsUOYJ5T4Y0MbRsGjjJ5jGJ/VlKqZ7288Q8EbORA9WUTLtOTAKuGbAFut9/p
QO/gO5IeY1Z4Dfja8Vx+7okI4fWF6osRunZ6ehje5QY008xFZ0DU8IpqFyNHbLDgbXcjEWY0/KB7
COEtuKkU+WfJ1+ghbF3VLzwn6DFyPcb+CwwRF3MvsPJn2qS/yndFGXdphaVSsXK2SsQy3i+7YtbC
dzDeCQxLvCf6Y1PSwuSRH7qOK8e7W7x1KoehKh2vY1cmvuB5kSpLBjh12gvmod1kyMgd/VzF/19y
KlComyqZnaY2qbCTejLdUdxudkMoN85j840q2awt0/q4s7SaEUO43OsvADdPmCk2Wu7ntmXOBkDe
Va1F9cSx5IO0YvTVWMMuyqbJC1Y7lL46IYUWGkRN9RcDEhIxwLjvSQJcGAmT5dUyqBuc6iZzvZ6w
Yec0HgriESyNsSvfaH3W9Ha4t6zO2bu6Yu6ii7D2zTFZm0ti6MbZzXwlxrJVznPzxhVFSbElnJPC
/ztvzyMteRNyb6dtfbqYveJny7D7SNsWNfLMZRye9xdStGIR8z0F1RoVTdO7R3t9UB88TwqExWxf
90Z6kYVqlqPMH/BL8RazO5byrj2kPNIa4BiUtmA5x6OGIR/YJGBiVVv9FqsFMZsYOBm71ISFKO8Z
WwMwHBFKuxiazijKdMJUz8ct4kVAPAIDMZAiV1ypaK3RtnIc0BGivpHezH2ShiPXmywVpeCmQ1tc
38ViQjzBJLbOF9+Hx2xTXCC9yTm8fnFvkM7+Pz+Jjko3onP+JijNwXpxgbnrIQpxJOuR9JWI1Iow
+eycUFKYQpy3B7DUhpKQk6NB3ycVL36IaQNDl0AsM6yROMep4bPaxzmpCTjfFJgsp3PkLUZUbK+9
jI0fulnaEKmNzmp35sU3oWpsUkwUhASKB9Hw6bxHw0+40t1jL/N3pw6K5pLhW67RtvPYmkJAWcxM
x+bgISq5oQKZ4hGuBBij4pd9V+Avo25kOKyB3qJx0+iEyJAvJxtWY9Kn0XjA4JTjKxCzok8BwszT
K/FiTAYOOBuDiHN5a9uNIq82iibcTwtkIk8kz39m9ueFebRx/J+u5R533ktotRvmQDafBTVKAIwd
D4u3bGPLnMIW79EypGVjZrrCY3NAznbQEoiT1ssTWDkwtpSsb2kSAbL0AUKzZqZleUX8IgqyzbZh
/CfqxPYV6mk5rdmKHedJN8tcA2NcJAhmJ0R1kIzJ4580fje98GmKBG5Jxf+yB4iXJJjlzd0G9wa7
aLy6Jt9rBFC34qPEkRI43RPFRMi2ggjZ4X4j1eS8tSNuoWTYpsl9830NaoggQfLvy5U8lFcxhrmK
Zg+/dwlxZ6uNmjEhnzWXPw+/sq/MHRUv6mPliYMJ1bjckvZGl8dExLYqrm3VqpQsKUaiDL+etNN+
8g7UgyRUK7ZMcN2aQK/iQcpyGfFfnjInJYdy/UI+1Gl34a/3uxH650ZuLdN1frJ5spmOpj40NjdD
oXkUw/wNQZ31BnXMRow0taKUNQXo2ZjrGKgnzbQkF6CKTbRGcRhOlHexTXv9KI+otCP0Qz3K0p4J
6UF06BH5vnqDL5sY19yOL8cocJhlvSMCjiER7xWz0K9te+RMkT1guwTeRxQL1CHJArX7UrVPfoZ4
z8MQPK36xhCsxCz40PfVguSTD93QiPo3njsImiJp9Zkj43uh3Rzb8MwSB6mt8pcE+xjvcrOX5kf1
1VFGV2ZR3vGEQQCZEYM1ZXONGQD4wib5gBR/tF81ym8nhEzUvBMwKSfIm+i/3U9HZalO8cLp2HSK
gWTyV/8e1wZWy9ovWGcFTgStl34SObFkQtKJukYq5o0ZdOC84ZvQDMtAunpdxpgyhm3H6RPSIK+Z
gG2CKf2FIubrRaYTPCYfG6FXYxTs9JmNt2ZJVxeLSLRX+S/LsRcWb1+WIZ1T9NAPCkiLzowoW9wO
9tDBh4gZV7QJ8TPYLZH+Akjnyieu9xVn9F1WkajIjYnDeN9lk7q68n02xf4K5g9dkDdxZtnrhwOD
RVoHFwizViOYMxSj4oJRSiKZ1+eqlY1E1SXI0ZOghkur5yQaqpDHfkDVnlRO3S8c87GO7xe9uFKK
r19SY2iI9HfLSUG27NLQvdANOG/EMaR9JulVqjVzam09lxSyB5tH4Y0jnUdTs/xWWn0V8lPmJh7d
zFg21j0Gboq6234QqHkMeeeS2kRF3diUovmnaQ7+j1AbsbAYd4vVX9QHqH15GAY6Q3iJs1+jeQx1
xBBba7ETczQrF8PRB7g8BHWy0gnZVu2l27/WknECWg7eAb9SV+kekubt/gJJcvf86KxcqExXIe1z
4ihWoEMc6bV8Nl5vGqcih4Sw2zHLDikBfZkUNrKgbuCztxEqZ6QCYkc8jQgIdT1pvFfFPgejwJLT
6qLDUJOLel/dVBh71tPZjqw6qqOxXe3OVZTYwH/Jm4e6wdejz66XnJEckHDVufctbZw/5cJzTyH+
x2uFJ/I2a7M4/92YWfTR0CL42oGZai8ohhYpnuv/7zqa+5dD5iiKsf6g68KMfDS/ciMeZ4vxVj0T
TFBc0fCY6KF888RXfk/2FOQg+g/dy13OtG9s4OzurjlEUE6wUx9dTVKrzTEupH0VoR5J7MgvN3eQ
vX5Bzk8Cy8RQu3IsqwuXDp7hgOWqRy07XXohr9z8Hhx7w2P6vLIGX7dBDO+l4zmU9arx79BsiuBg
tcBq7WV1FpSoKYE7lYWqRajOP6cufSrhtSiGJ1bjxvrfxmR0c61Q/AWaHFD5xSgYvQqa3GvT2gj1
kQhbXpVRUTQCzpcSE9H+EA5U+ifoR16mOOK2dNDb8DkcEXpOVUjsBgr1CQeybV1cmZSJ5PVA/k/1
l2VJ4kReU50OHZLKs3nPfO25CkS2pVPPWimke1avRPAFgvpqhHx+MNTq5VCq3mBZqL3RNnujTY/M
EoKNVflhhlSHOKxVupkNqRGwU9a0AKuLN2g52mCsb2gh7f42R+JAmE4M08jBaO4qjtZDFyKfP8wG
BATRp4cjjQxi+mremphfUF9sIaDcjltswq5ZdNaKZMGqphOuguF+ODOEkjgVOLzF/SqaElsg4a+k
hz4bj9jecIbKF+FDyy9p8NqcNOYaZVT1Eaw1xliZOyVTiRWEvSJUoqTvua3Jw/GhZj0juCRHCVyb
g5kbNlgLLMnEzAtk+goZhERnULugUsx1aJV90B0nBpKm1igEBBbBc3OyHRkJGztXuFwpYTDiajLM
osLDKmCTe7aw2C7Gsfeap0qpZiieGdY1Rho8je8aLBeiB7FDIQZa/n/ltwWgsaRbXyEAW/DZYC+c
8Aw1jlB8V2M321otLjdZgfl3xIjr20oa0d0J96yh8RzF4+CqEOy6DyyJsFv0UxX/fXqm+V8cL+RR
zr4jgCP3ZLEVqvGScbfbqqnveDQozVeEeRWEpWu43QP5pLgSFueygEEWFHqar4uoB9c8txMPOqxw
8HoKT+6hb6AHS7f9MqureiqF5dxcwSwtH1DnkBNJDx7WcW08WmTJmIudj7p8IH1VrsIyNmmQcerA
34edbOw3GiYsfFHGfHGxf4EhSAHfGTHZrE1ItodYWSR90pXl6g2TORK5h6YJDS56gyIRQBDT4nds
l33KmR8qIbpJogux1k6Wl3Tc7CfWKBkKEDocQEw/lLqrNiHMdTHEWVUqSugRO+Nz2jSNTq5UCDzi
caquHJEtd0sUFOa43hacFSoHaPb7TKZuoeeaWKOnDixJ77pPlnQlovNX+YIKEmeS4dpSximWQz2i
c8RiWr2zhu4Cnn87RjQb+DIZLH1EjL1fhM2iw3vrDNuRsT7rDMke5+SF1eXrQbDSgKGfkvcWbjou
xXnm41BF0PSPhrT1y+8DrDpkP4Bqn5k0pHXHCToENAbkZ40ZS8XAyPV4WzB7jO4vA3FE11uHx3jN
/Ja1xDofgqUgXVFf/exbbtumJTYK74lYoozuWUAFeomcPVTUwFbSjwHrL7ntgzz661vZyExCr6eY
47iOmYBqpzFGRfuvRxX8Nra7Cpyy4PBGTzlYOMhRakH7Bs75qDlTQKF4mOD42krapP7VMB6F8nY3
Pznfchzp9H13QcmOKqVXVZMKCYDutbd19nM0fjlM5Wcv4c+rUe8wy2OIqeIzddd5YriAzN7zvvVj
INZ6m+AP5+Te5P6IoB5QqryaXBdGHRR4mPe2JoRDnUyiq2sMDvHseyyVtARpyI8aHnhUoRZ62jkJ
/BYM+lDuQnJwQEhY2GpjATJrD3SujwEwdqad+BvTM1q+iJX136sj1VPb4ixWuVQIu5dWVqJTlH4T
iNFyTAubcd0Aqh6bIkfCDuHADwr0s1XdRaIYppWFvoiJzkMs/0XtJf3jotFLc8+sG7KSAChrk9Ae
Il7N4cvcary4khwq2v4Ci+9wcny7VX7ePCMmpG4Dye64b3K4GhgcgrCEL88C4rsSpMkd7vZyBqkt
NjHxzLAZg442WdOmY9eRmu/N5L1u175UJWgZ9rldgYOd3CFH9iPDf3phi79f6w6AXZ/r4z00Izar
XVE2Mzmc2h6ZzonjxiHqi1P/wQJ5VsBgw+rn3R+aayzDw8xHajMIEsQ2Dob/o6Nbb9XHBO6tHraf
ngmf8LFC279gM8GkqKtdi8fPevB/2E6DbkF5afnGOnd1nxKQal5IZjFIevHNFCqTpfT9iSEy50vz
fKffYZY+av4HZkV2GrFFSiBvdlzIA96ANJFeH/K7yFzTCZTeeDnsp4JiggU1+7gJy/geAeM0Adqz
ywiCdE8U61KHXqjmCIJof79kYzo/Ki6fRWaZdO8fOjyN5H0M3cTKSGKyvyk+fta+5sYCkC4boguf
Hb4rfnXwN4LcmJ4KH3GZ4chq8hQWI28BgNzGu+ElIE1Vrvvt6Mpk8uMKEFDrGrNVYmN2NkuohJD0
IyNp22Dq6kLAmCZIfWyql2dzg1Q2M6LVnaZgUbSzh/89mTq8XKqVFiDjyJeKHK41HAHCH18nBAFG
trUDPs4juJTQqkxqGe/GlMVujmwjOdW7bXw4jkucsIr24scuVuGamaKXy/Mx9B24MHfbe6Lu/Rke
4lklP7+80MMlvS4T83zS5+ymuO/2Gj31KoZ8328u+DVyJyPH9wr4bWihnH7ktsEokyFRfQ93CG6a
PqYDFeRdS3FwPDCJVPgouB5opD8+c1EZmPOUmOTER4nla09PVOpHx69DHrWYmc625ejPls9gblvw
Ziy2aSxHJpplDcIScCjOZ47CorERPaIXNEE2wmjgTfWwiuJh0ps4X3/h1p2e61pH0t8POPBHUoYK
I//Alr4Ajtg0G2GzNDRGsfWtLWvWwJLP6TyyfsMFyFunqXiTyQUImBQBSxlORYfZXS79c1oHfi40
AjnMu8VZ3gHe7PSljAjDRElaCn//A5cgNxdltHGxc5MMDhNX1pZ0EqTQv7lXFKb2KmC8XDLZBPDT
8iFpj88vF5luqeA3lddgTxGAP+5F1RWN+KPVzNOPryYP4l74YQ7rzIokd6kVjB+NDUGFW7Zpl7z5
DpBFxWnTUdijh4FLJ2pO4CLiLtb7tpyCJLWERW4J6bKvgNyksO06m3o6ztcwnK41d46Rrc93CDMx
6lXvkhAOR+She/AUnaBeZZP2jzQsImaOZMXhpbhHczfLUmJyKZm0SuMzbgb7iMqvB02BnRFN9Eoa
aZUvY367tR+bRGJAKCPxw4R+cvQNBraj+rhIJnk50DkWca+CzkqR0nUJ9PoobANg8F5raTCirffm
QzmykYBrwaQzd/32Bly43yaockYjWnmRZpA0BGcrbaMvXVUE66/RkwC2FRg2JC5yhSP83lCgenxJ
24VG+Wy0VF5MYPEQprupS9j3qbIZAIHx9EtwireWJcNxXyb/IZFZ5sz2f/MLnAtawS4etMobaLVE
eGn8nAtZ5USBd5hNc1RazB+oZfUdGgVIuK9f9sotFjwpHd1ADnfz64e+GGMqoDRvAvLhQYAe4X0X
ywPn+rdhoZEKLT2fs/MwOdfLb614bGDqVo8bLJSqYa9NZWeLe74pQ1YMzm3ETvGsT84Jm9FjWXc3
3Gzr1AR0yCfr9XuKE2K7isiAOGKra6IbJv8iuSdSF1mDnne1v8onO1mmx6D6iPlX0/nsZB58YihA
R04Uzl2UjcMYJ5E/2NVVMkF1aV+u6Ku0YsrEBbrG5NrWW98FOIj0nioVw3cguHd2PYRjTHQaZnK3
4bATowMNFUqyuoRJPKT4KQFMZwgFbXfuM+l+FoMwAO0afwTkAJvUXKUPyrvoxf5dP3GmWhQzsJRB
62J6CgQPtNM4/ZlAnWKsfAuxcImE4ud4mvVNn8MVPxtHgyHCOGxONHHbRKF0QNViCIbIk80pk8iz
zOpw8y43V29kQph+S+7HcLwIj+rYGnvXwSedaXGb6QDKITTSxMq2QGsqH7kSpucFfx2KcQsBD5wa
bWuoXB1L0KMQKztnrDzvOcgO6TwcKaUoZ4M3UPUPE6vJQQ+0FEN1zRxdNI4RCA6zWAjkh2Ra48lX
t2lLfVuSGEWYUddekxAenQUJfNmTS5fZcgqw7a+k446DpZ3BB4ZDyX70OD+UTA6KprLYtxFXFCT9
2+IW+coLtB3HQJnyPzTsjnrlf8pcCJIERDl+Xolf/XGR0NE04pKwh3uscepS1KTxETfRUZFiGbkH
zG8E8fYQyIlvkDA3DsWYuyl58rs5R1Cq6bwU+qfmZFk9jml9HDIOHH8lqVa4ICtSW/M2+Tvt65Mv
yCdpDlYWp3+VHAWjIAdtBlG9oWmVvsAOR9UyMu3D6Xh7otEC7fge4Ke8tepIpJxXJCMMLfW8xfYX
0MhIvq5PnpkDE2A3uS9Gsf5PNrrNV/A8dPqdwEabuShNcOl71TNoiGCDfF5Sg5vRQ44Su5GlKCkF
PC2vfTLjloUjd/3wteC9YDTHvS6zyEeQUK7HpA6zLAguH4Th+8djuYp86ZgXVzS3Z0q33mOajmFp
+jjrSSpnUUQuD9wqAu+L3fPp/OqfY5NtNjUs4GltzX+v3BT37Xubzfb3648rTM3fr3PqGyVzpwMZ
VMEiBbXD9dCMysdhpCuwxTlyU8LmZM0sx/udJzbdYUZWfEtbhwwBpRit/qITy3v3OZJsfDu0fk0O
qEa6AFLAme9YXJl2dgQkyYAT1IILrgNlaE6ojbnpolQHDx8CdwZm1pAnAWdGI3+ctjpW0qRNjaEb
9/wYg7hxZDQGameA4gqI0Y7g5BuBGxiLpD938avoMluPVcWqiG9n2XAxa5eqWO5bIN7l8qBrSLeJ
xJcBGRPdUnbA2TV2pKTdRxBGaVKJKQ0VLzHnTF6nIxtVmNb2C6xt8DC8wXY8YZ2Smh7gnCiTyhKH
hz+z6j8DDNZpkEbEGF+6oPTR+uW/hEzNV4LpVso2I26w8DKkh5dgKsSSvHYaAz2OKQO2z8L5xddm
94A8Jw7Cj78itTOookJK3ZJY9ztBGOFiaU3/HXOwouerbPzz5HQwVQDX4x+ZHCX4DXilE6C5UgyW
Y0zlIDP8rVMeRRM8S7BHZ+OCkIitZnV0vYbh5YcvWxl2k/em7jeYk9keQIn1lS4UYKb0WSc7J1vZ
Wv70D/tPZB6DvV+wVvDkF685RttN+0Vy7BVKbpZETqwKVBiA0lxqW11XxTVfz8J87kNoDo51rpUI
D83m1Awm/dnNl0qfCaOXSFhresSCFu3enboju7UkAl7EI0kEsAf1WFmKLx5zZnPCQtl9VnpwE7Xn
a7n4I9Egvx0o14xVGuKHfPAdGxEdKz1N+oZlrq3Ui9cGkJ4/N4goQ2Ydv6mVVu69WL57mSnq6HOu
6waxg3G09vOIU6aTfEDr9E6DgOVYaJtdiPghzBeqM7EtYxC84diyichV1J+gRkoaQA/vuMEUcwvh
5r/8RK67jTmYbseyMtjstulkrZEc2e75+9xKfa4nSOUmO60evqE+UTzmF01vjdNJn7DvYsWLOQbv
Wr6tj4j154r66B2+3BeqIsrDCzbsUXIgNMVJbCxc213Ba3YCpCpG+KMVLliugL5uWpHcNb23dVBP
U75LwI0rldxnLtMVfFcGpuiweRKfwAy8jE+GD6Dd5DbRbW2QhSr/uUDs4sN0PXcPgBHZziCYhGK4
pKVJ/AyMYZkbc+gQR/CdChAGBXuO6BlaEU7ztVKFoJfncuY1lWDUgav3dkKNZIri72NaMOtWx9bx
5X14Be21JXex7vEqpa56QXIkuTVEOuK5tP8lFCpZNHiOtguwM+Qql1hdIC6KtbGZxVTENaJwwX+Y
VfEQ6EOTg+RVBlNxkZBKxBecYzYPWyhG4lVVEwccR5PU/KHKrYbphWrFk6PraIgHiFQHEAV7g8FV
T50i5x4BI3SBDdxyuh0gZBZaZNadiwCZuIR98CyY1CAyUHzRXQZMdWo1weGmqM2ayls1b9aNgZVy
pH6IA+THgZkKy2D2IFGtoQY835gONKhQ+Pkud8HT+twUukOpaxeFu1kNo6VT00NjitgW8KEH1m9k
Ut942q5RujwNie1nq9U9YykrRQqCnQE4J9dzlxL3SAnQmD8fqWSrV4+Fr/9Lr7xhQM5mrpgPPD41
RVyvw/kMcnK2jfhU01kNg/xhluPscpusmd/rV/vTf0MrIl/rfpsyHEOGBpqBL8ZUFChB2TkPfdx7
m1eFHKgvzJHx04wJsPrySUSfr26RwHPMfLV/HjU2hvpEeMDXKIezEhy/4+b1bcMEj05OeYSDzJMV
Cz6U5c8yakbFF/3D2pH89OmWBDsjg/M9hKUBcRJjeGSUgcyH8v+AqITDl5pM4cp+bTInGlTnxPW4
NX/rbMDRTGlWf+zmk+wo5slnbZgRobWvnr5sCrHgSswmxXcLm1BNdE4RoIf4YEC8e8xFw7oqjJDi
ZoTD1u/3H1jERCjU6fIqo4b86OXTaU9aR5s71+XQxU64flhXg7eUEzuQ7Exa16b7JZxD4dAzgVMP
J6UBFTCOVulPPraK973tEZJGX0eQ4so3jArY6L6ZdFkAVBhTXIusGmE3uVfUf+b96gVy5wtbN3BO
ypVUJ76D+FdTvJ/caysQiLnT0rCV/Dm7ggp4NGeQZDIYlr4i4jxLynuCD07p4s6MNRcsvlkwOaNu
KurkZFrz0zlejVN3Qa3zKDZ4fu8F4LcN07hofdmgrkKympV8o7e9f8wB2egLyUmAbwJ5hOoSHXAr
Gz//ICZHailA6fJUFM/C8OVA5i8PE3lPSstycvaW2qwS0SxH2lYlGdafq94hWIevZP44Gn9Jt3rN
/c/qARj3prRI0kk3c3c9OvMqlQBOOn+nYqgUncltcr3HiEe4mXo3ERDdsuYpQx1+yLJ+Y58IEmAh
f33HFUq6C4kDyWF3bUWiXR8bCJ7QBrdxkJDikHCWAEN1N9P66CwCzt2EM0Y2shf7GrkygVH70DPG
5KJT8/KyhRwhQbuebbvs0p/jfM/Ansn8NrLEtw4UVZZxrjoVMYEB+ffiAjHHsilneuJ8oJ2rjNvN
yZBEH+zZMhE8N9pehDwkiQfu95wHcljQRyG1tCY9yuqNtcmOM+6HDVq0GFUoYMxa/Myq5L8dPQGo
3CwW+8rIrW1fxlCXBSQ+15ISjmi4T7+Lq004emNZrHvgr/bZlsUZbV2FbcFAE+VzmTBXEuqKxFE3
8q+RzTa7+l3DLevgMzuw8+H2Xv35sUG1SKUoukXC8T0/M8jmuiXYBN+zq0GXyJB7ZUO59+OJ471o
ZVxO7iwJZtF1bzeDZ8wB/yQ9bAOfhWte2NQ7ykukgt5FRI37YvH8eiYyvf5QJqzC3SCGYw0U7Rsh
SuwcpqRJ29lELjnBgsnVMv5ecGsNnkajVPlCH3N3nxEx/3qepg//IhqGzlNf5NMSVd4lVeUrzJgG
hKfUDlcJLEGjZBf4sY8eNEtU6VugyxZDymmKbK4DxGeV5oOLkVIHoQsZtjzqJMSCp9JC0dipHS/b
JO+WbbMygrtBdq9Onfc5Y7BATQAnUGy17lMtCgtrkyzjkwpGlRhc7mvHPJJZZFX4HGXTOgNOA9VR
+xkRS6osH0OK+IkFG2FXBkR3QWb/g6ePTLNO8XZp16zZTQqaxcBOpOW8i15cYL8+NkPKa3nSwEN2
Onm8xRA+d5IGhQwnLXrPiA8V+Sgxd6W1Y5mzPSUYj8oUbf/TjmkqAB0lXfxW3rv6wxGtrblMQHSj
3+zpSsFvvjGbgke7N4BF3utNba1h6YH3jYLNTKrE2byNkQT9cUQSg4KHdvGb2xeXVva86P+VIWmp
B7AO4k4qavMotgTQ2Ua5mPWTli0f7Is5w9mGPjZcxFfAjsvNmj2L9sBxOhy/nH+yvMVjeqarBQKb
bEzoMaz141dEVqJWEiaoO2eqPMoucZRxKq8wMka0g81loRfDSdHTlYkSiaja466llFRbnTk1o542
bbmEHamV4VKMKWPrV05pMo2avR74kArv5iGZelgh7DIpw06yJIjYL72sSQ40cVcTGdn7xTTln0VH
6saQr0jUKwV0QkN1JEVaSVGgXrFU8HLNnHP8dvrgoC7/MqfJ7BwWHhqsnBdGCMO6p2SWVJf3L0MY
uLz/3omovyVTC9L9q5SH4tOE0mSOkR3cLxE2+sqD8n9TbegEjnZXAp9lgnApFucBcgi7KCFMFUCz
fLD1prhxuBE8Z1JpvOCqitlCJt/d6I+2ZD/jF5G+i7rap9UBZ1d/9iVyGF1RTakcPMZIfb2taAmU
EGn+KgP6/17zaGdNVusZCVlGch6KkuxjabYagtyINQPj0kD3QVKeH9KciQ8i8S7H/n6UkljK+P+S
JwOHvm0l3ed4QgzPZd/1XOqsgWWib9lvn2a8QYxAXCjJUyHBq8zkj7R829ZMDE/MBqp9YS104g2P
vMBRDteGR5gYFFRzR6FHBBv5YOj5BVCQT3MJ9nrZah7heV1QVToiv1tf9/k1MWlvKbr5YhFgaG1I
ufdz+NOyFXAdMJdMHsaTPLYHNdGGkdY4+FB/zTSQESRlR1v+GUmWz5K4ryYv+2XCiCV0J0b+1C/u
Kibpw4DhpoFerkHbFrBMEPn6CtKWB/HtgnQyytygUtdXDs7AknMIJmGWln00gEBB1valu8XgvWhx
F3m8oFlYrWyMuGAlhWo1fVt7lqs1DZpIp1vH6KM/IbuRpoSH8uqHdMNxdUBVTvyQQf7llwA67hTz
CjIIpgegWMvXtd8AxrF9S61AAIl+CmXNCe5X7kRwmyaFtMRIKzGjOaZfcnTkDNzFEckZwnUrSDDH
TR//vXrkVxZYYoJF3bInDnBiweHfw9T2/qcDp8qMYK0RBBfrEjG7de4O6mAJDFIawB9Ei00uvx+2
vI4qmd0D51eWPjTw3b9Kup5vLya1mNrElaFqZxaVwL8F6XkZaMbEveWNXXZRhyAS6h9r0hO9hZZB
9xpDZrfPyR+uKrkPdERVA/AyQDjc2eOUr3wVqLqBo0T4ucehbyARPMwEBswQPMo3bW4qZ1Xxnw85
e21Bk7G/A0Ux7aUzEG6aN8jB1Iv+4DP4JBEkHu5WqKqTEvxyE0LqlyXEZkZqnv0LlqIpXwLoIm60
DqBa7KFC6fCVRRjUVbr+V2q6vUzjFZYHR7QfAD7DPrga3uZHZKDdGqdslPeT7K9S2CcyXrDeaMZf
Vt6YcCoraIT3uQItcU3TeIrZ12LrYgSxaDVH0t7cWAqsyo9uxEML6LSkCEjN23Yhm/5qFl9MLG+m
FNWcmbSbVf6J/bnSu4yBTUi/1bxb6L1CCuN1kCeUSL3Z4qFrLBWPu2Qfgsf1vYNcu9ZTFW6BYpMl
DY56tnBQiz0fYw13C9MX4Dm4glN7AL5ftW4QzvSgxZQFileCSktzYrr5h9fZYU0GcD/+Li67eh4U
YBVoO6EsVh4QDjP+M9ftnOmBlybqyexl01+hjUalxHXIhQ7s4dLGPbSIQ1HEsQ6+4x61jOJr74Ct
0Lk/th9nUPgLsI/OcV6n/Z6xUnJytG7kCRBJgXVAjL69PIjRxAghc74I2Tj2jCu+TtEpHEyCCaJc
hbFQRw31SYKUQcTTUvA0zfo2o3YTD9wrdPVYlmJV5aml+9xJXeoJXA1enmiISDsWy8oqcMYgGMCL
uduJOnO0hD/dAG4lcwCN4HOvAjPIdgvsSR7c/iMXkrH4o/Fgc3UAOrryLiDqKnuoCNKvqm4iwrDC
9uqnf2NS88i5Ix5Z2w1+id6pLhYKp7aujH41WP3QhUnzXdk+dlAm7Yc9Xoi7PXXJCBaojz7sL9xq
5gwSZOrXU072QdNu+lYI5QgXBDCW98qRirh5+seEuWFxGVDKuJQu0X6WXLEUnhayvUv9Bj1RZ1Dm
SbsNscPoNGnqh6HoaVoKcg7UOasfuBfQ23P4EnE8lcxIjot7XAk9XclIWXvJhFpEBPr7LdH6oDr0
hibIltSsXG92XL1y1uh/S0eSNy00XQ3AEwoLBuUi9ZBln90DaE/D8ryG9AfxB8ncZuwJu+w9xb/H
Ok4Q0Bhxp/8IxwohwYQhO6sG/gQ6SkrV3j+/FfEqgzvd4kRVkN7JyfgPE86YYl4HvH6uksrbY44l
LgGHJOTULbWAAumxE4DIbMzq3lsePykDWaSn7Wvk7xWJe1bT+DtF7Z2xUSY/+6LEOm0+2wfgAO8f
tLq1NKiYmT5a7mHovnmSGYXDQWp8xynBx1jIx0WrNFOp7vMEegr/Mzio55P1tGDifTaUA5/fIpjd
Vhm7dYWVZ7zfQVYi12C4mQlguRhILRqBpGnMqs3IM35lLNmX0OkdowA/yFk/D7MSpWrT54C+B2OH
IZMK50pgd9yeNhquu9z9jontQIL/pXKdsYolaWD3t/ntDjQoXEAfPCMrJ5Tl4j4Od7bSG36iWYOd
s2oMNwYTYCJcyxmNPAgBoALdHMB995mGuI9JI0aouJl5Rd9TXZvtS5pSGUlbbLF0Li0qx1K3Jo13
OuxaC0O8PPu6zu3lkckEd6umms8pdENRGSlDMXW1rKniRzFgDKMQzb7sqzCdDxXH/AiQwDr1S/Eo
/IAVxQWKmuudoXglz8cd8UspykAALRPrT9nTrxglDCqPHZdWwr0q0iVZOxkbPGQYXOkcmRSjZg7k
825lCmVbIFs53dnEHHx9bG0hFQ/bbEtYkyS/poToKwi8ncSj/VJ91b3qLaLu/Lr2ppMCvHU6oOdg
aowA6m3+6/8A+WHSt9szl60TzT67Z+2RgGMFfC5FT/9tPoNpqXo339Eqysb6H4zr90qV31schMYU
3LGPuxFM+2zFJKFXlL5Z/Yy+fZ8De5dLx+9RKDJYt/50FsvTfcoR2J/8RiQw0fNs2/auvDgI9DN5
Iax5vZUFb0i+uIpgbQRBoXqdzvAZX/ooY5LSgZ2a9tk/NDtbgVTv6f3RxhOGOxIJo3fkNcTULaw5
ADDuUcdqmi/GTrjGkTzjd/d4yfaaLQZsKUD54VS3374kfNZEcjA4I90CAHKDBigIZkW0FdS7MIKo
BF8m5e3zj4ubTg+ymmg9GvBpkJXIMa7spDFtWDMNa9dkQvsOOQzDo1l0p1kIQUD8egRGbl0bY8wH
/vy6xLN6n+iupOTj1haP9kJ3FORS17pVzXX1joTtwGR38wVj7V+xxnDl+FG2wAWuJVLolJ1DBIWR
fg8UkjTxbq8lx7eNt+0hTUX4OWc+KmGrT8Sgnujs5HAdmnRYzDll32TF8ERfT+Bfa0R2hM8i1I0W
NPhls1E6B8f+PD83OrvQ3//CdjPtWCFdR75CsqwBJ4H8TDXFzTI70MGs1PUSwyd6WEM84maZDx6p
LGgEyd5admVJepRJuWFz+7oqPc1BvCSIQlHL5JJ2exy9+n6k7ipKQvEkD8nRYQ8iuHhgFupxqMag
x9yth0YeJF1VvJR4ko0Wl5e/zZ8ZA5DK4KagE3QxWJlH8V9PT2oz6LDyQNpD77gVp6U/ebXsvSw0
E0fNO+3JJdOf6aexBm6W6gcjn0HnmQKCcm074vV9D10eTs6RxwEzlNYHp60Fwt+xz4mxs8VrQm5i
MqbfoLHGZ7jWZBA3CLcMQhFXPppgmYSxlSZ7b91xqvG7V2kDc0sxpdPa4wsD9DOVUPSVahPnVjoL
gD8uaHS+CS6cw0impm8CSjRUVCag3nZgsdCfSBIGNRKcur/7pr/GMhpyeIRdZeU1O6W0z+0J0p10
pbVdFRG2tger7Na+YA0itEDp+cCEH5A6K2DMsRR0ju3/iDIZ7TSnovShdMPY8szfYIKzfjzKqcZM
JBTrHLiHZS6CaPQFB/grs+MRym1tXFKfGb8xt6q0FnporiJGQt5w3+hsLRfFYy6hMVKlhaENWt4w
xTq8u6C4ebnPeJvHMjX6lYflSMNf4ICJOO7eUXVUj4xmb5pVR1ZDRpi08cfwIDi3vLpINF+zrH1f
NX4o7GYkroiyfMxFSRCzh9Nq4A2QmPCmQxupMKMQoPciCwPU/DcJ3n1nl8ouk6Gpsu7+1ZzPM9xM
9VFHNPabdhrUgDlHfzRLiy/g+JcKn+NhiDfliB2g9rlVaeBxTClHgYU1XaViERBhhJ7GBpvfH0Kh
BVyegteVuyDO/fCsiV1T3oxrSgUTjS/iDQxi6ssTC0ekM+saHJWisP6miLhzZX6j7eIwnfipHyRt
iOlk6rJnZVOJw7lrfQdX+T0ZkS626RTkTYfVdXyb8X0yBjfsyX8tve+MQF57fCGP+lyTNhlpQiLq
IKONuQheFHEav5bxqUNGCE+Knm/KxDVQZqw836nxuWCplFNaP5CuEtImQ2N6+yxTMDe9UxLphm+y
TqjzdIfd7LtcyYm/jTy2vShwTIksDoHXkejlKCHjHEN/8YEPEzeJ5fITUUuvU75SFowUqJWz8CgM
pAi/ukMlgDT2spwMEnuvLSXLaQodg1+QDLFNRBIaQKZCknBBz6aadLiev7j8d+cauQMUU0J/P4ja
s/4tNoOtNk/kyxXwLZFK1Kq2pcQfWk9LKJ6Wr5c8dnRDWD3H6byoFKQnSRcF3ovTmFvmwWpkWorM
VtBQwSgJxv/DWRCAtt8eFgzbSsCs406b5MkSOsxDv7/pECL6Q1790iVcMJVAoZT+1KZ/w70PU56N
B0FO09DRXehBYkmoiekUMCA2ElBKgNcRnB/vt/MvnPIesvhvTOiTGlRsS8lbk8dTg3eVYHQjeV+9
zE9oWq8kLPIDq85XcB8OV3Rz3EQp03Jm13X5sbK2jEVSghFvzej7sWrFRyFauEmo7WWqHZ7WPBLu
Vklbhor3RI01YIs/lPGybWHl3VDe1sCmO05n58r9t+xPkgRF7JYUZiX4GkNfFciUsn5TTsFXVsAJ
LyU/mi+h2HgWs7I+wBenxlrXgownU237teWfRInqz0ruvzr5esjXygqe94c+tJ7BgtUlyXo9QOGt
it+qz+AydPD1OkwDsxTwote1nBDULlCCciSgCGnwZh+xqwk5/oSzElEBShv0Q80Au/aOvE9NIDcL
Pb30dsaoDX/4TFkjNxp9a54XLRqzNyqWJPa/xBt4MXDc3m0ZJtoox7V+DELPVjx1ZlYPXKa24Es/
RIzKkxSHjI6nsqSnDCMFAHP3vztzUU5fR+bjOGmDnafNLivhh1JnfZmlVXULeRvrazHZmhOd+vor
bzlVuOQSF8vkN9GRBIQYm/A2PWRKSz4H/tIJ2OiX2kCK8nE4U9JA11brVQ7j+Xbzdw9VSW8u540d
G4b6fYQDKXYDo+3hGtrYOZQ1EiWMSZK1mi3blAsdfVnEC2YXOMCXj+C7Nd/bIULI9qNgMZ//Yymh
pwFpwhdkwbF9QFXf3/8cuJtqUyJ2gdMIMrE9+/B3ZUlrT2qVntBuxU0mR4x8hHuEB6qGgtZB3/6d
ztGwpiiP1ZrpB/2oEFswxg+RBTbGQNkjoOLdhO+QI7TAQgIpJ6cUa2aXMEkRKRXiaiu7mxPoTsub
zO7hCPY+kUI4iC/mXcRtkfizmjhj/5zfW0GJYefwTlwnbCMaWGbGJz/oU3za0p/RmXfUDJtnneTg
4lorqgFKPErjK0qTkfHMphazuLuoCK5MOYSg/Stqb8ns0z6bgA23lnPvuaGd4KV4US6PrhE9e5Zx
ZLcIIXk5yEemCCwQUGRmcZwiaJIoje6XNRkWleUvm8IzKORwcBXO3290jrJKo0SDmIibqcHS1QMI
hVKXD6Bdrc2qZa09FADg2QXrMTi89qUISuRtGV1kYgvFq6JglnrEgp8NCD84jlmRPY5gCIY60Utj
cGOGD6En/Iz+o9NVcftACE7EvAGG5U6lqMvtb8hrSh03poiH4C678rxzO/Qp0m9Tntst2cvSilMT
62P5hYiEQGQckB/KHqCsG1Bc975ulDVVEXNsUaDeI9N7/Xy9syTvm4rNP7yaQmV66H3/lrDPKePO
S87gn2jq2o/6Y8VWCM+x2zxONa+7PmKX/A3fay7sJybqpGpzU7WBram0V2dqxe7R+U3isCm4+dOP
jL51ZAh23ibxoIVeJWFY09eYGWnYFDQKP8xVsckwqWgafOqIBPCZfrhwla7iDMzaAeo57+tsrTW9
61YWUTAFaNNqWo9QWbB+UtGKO5Z464Svwl12cIyjD7kTtVP3xuc1hakubR45nTo6pttfuwog6gMg
Up4Y3oP9kBlR0E4IDzaqGWAMyRwzy33wa4FCcp6/0dWTEm+5dtv2xFlj/DC3XX5/D3uU++bBObk7
H87Sg2rXV8hL7g5NMb565sRzHPTnYumvUcFW3vlUclUPBrbbBpU+Ofs0s4zgb5jm4brdpR/V5ueN
ulRnyy33h9gM42woHKky3xWU+KHEvCvjI6UNY32JtmByY229f5QGL+/JNJDWtz9gVL6AFhFM6mRr
cfr51qY7ofZT3v3gJM7cJqT6FhZi6AEM+VDep5qvj87b0IGqeCNVEBBKXPSua+XAy7nSUB9QW9ZR
Y2Ksp8P5aeoCEOH2IMfokp6aLhTjgPhdpR59m7rIfZax+9tiHSHcVjQ9eMGeM/Nb0CI0qaS1loBF
PED8eySAKUS4VEjJ72yKAyiLcVQUijJ75sYJaDiKAC3SgiSrrCuC4Rqd7thcjeXb5mNNYzjvN3Pe
B6dQlBPVknxPzm5RKGWHE8zBJ71Kj/eHlioLI9PTsBiM/novtc2Ae7xCdIqd6gBMJXRxaErKcKpG
aWYBWrU0TOtVwnAFSX6MEKos56auPfrlPga11DQRfSt6NA3AD0ujUgwcjCZI0cCRHE0e5Jkqws/0
xWsM4NizzEA7cPGrugTMan+6qVXt0girmahjN6/jtAuITL+oMMa7Hqc7ToUX81+IJIz6+PI0alB4
3qKFHb7K+XUbIN+Bz7cJhI25/z6L+WYdmhY9JOEX0TmowzLQaTfjPUK/1vNHpKUe5SpTFSgWu3bn
NE5FOWnhopVLor+D9ZumA6tmIuoRCqA9oDsSW4ceMh4Vb9ggW6HyIKANxVsfXxTDH6VX17yh2UMU
eE20gX0Ji/fp8UlImb8/47jTsICowLNfaSHnJHr66g8U7EoVw68FUnayyhKAnDNqA7QmvFlOUE8C
g5Nmrv6MxeVhxVN62fSiFTnZzseYmnvjDN5kHLgcaA1DV2v9ZOLgP7Sfv6Zi2tdvP+JuGDZtjshW
SsrDZYB1OZvXfyO3PblHQXsnoKkHIq5kj/CgaB4/+i6NCEPxlO9vNb9KqWXk/m5wGH2WwPu9LTIt
aVUAT1E7jtS4k3+yC0LBmrYuOoLs5gV20afZvaZqo1IQZjixssfDPDR1htD+Znlz8RKqp0fcveSl
mrKfejbzL7zfeyzf4M3uqbz3OWkVH9YmnkujFdteS9cGqs9p8q8Qy4mwy3vA1TnJoUjjeRSg7iDB
IOaiOEjMwHr1PXcuaEnwEC1mOG7z2IJkCudO+UZUbpfeHTucwUipD4JY3zKFgsDaSIQEAu7efUgF
ecWNozOVUNQJGYXEEBSlwlC/CvJkej68Vv1F91OrG43KCEX3wgg5NvjmnBBEXH7agkhC0Zkfvkuh
2W4IQiKzYrjy8DKZ8zbGkGrPMLvpvlXs3Gbvm1rppEqy/n0jZcmCweiRjMSM2wwXKmvNjc/kvTcI
CnI0Mc+Af4BkKspNgbiw9ONN+0w5vjZ2/xjomT4NXQ9uEOEBYo3qOF3jDXYIqZTI+dkDSjVG4fAo
WRygbKgINFBG3XHQ6rJABz9kOB9BE5pGEqxo8BFtvKIFtalPWX6HPZBo/cyT9JomZ0nsOhSjdCKE
wsHX6yZMV7a8I2JSpkMpsEHYjR42FPG6Ri5uLovmR+RLtH/BAp1gltV+dO39PLvEKk69s0acMgSl
hVHvBR2wklcbjX4sS9N3IdCauRrace5ZnNs+xVu38IHFAjd99r6OYBu4h0rxk2qfSi711kTEA1UA
B500KI9NPrv0shSkMo91MZwVlHaNlha5KrnxzykwI/wQwuNZGjGZlZLJ410RQVcOwAP8f93CXqQs
mBxqaak37vzHGC6lLZD/vRdFj2g3zfHFn9Qx2EkbwQY12bSubXYK5405NzuEeknQrSfyhhW+QxTY
yBYYJdxTEQLQ1bje8NsJ7fqDOaSWVK3SSrAcVNYuMz0ABdwA+gULXSt12F7pQCcJ7Nu+q4MjBzwh
C+WotOVtMCfWPHYOhK75/dpkcQ3P2OF+kaeuCaXfKSizX+8l19uve+LbK1Jiv/XyTNRjX71giOGe
DHVQb/LuQPFBFgOgz3TlH4RCacAN0exhKZKEoo2LDhOB90ISwNC16cxwmKXSP75U2gTLhi6X+m8J
TkAIH57z5dghk76nj5Jzzvsh8UVWE6NIrrMJmjfDeQQKba6i4amxzvqxuCfdx5dxubAkfeqg+eOU
d7r/Z382wxjrT65x/wZs1UR8D5cJ+26kUWaa8Q7ighBMw/Xs1fH/L0Qyf8bhbZlAJfhlift17m4U
xiHSHAj/bmSqpU0wpe3n+DiWH1sHeDLxV+KMS9uE9Vq+4s8Jaiei3WVw4SeJCoqaIVVeteT/G5JO
wtREiPifwIQgnxJTdOlGTy5IBrqNMdRC5VIy9GnE3mqHrgJk7WPewVOLx1pjMNlHkA8EHbFIFldq
3xW2LZb6GGCNoio3zqnwQHc0GawO45QfS5ERKGMNnJ0MsG2ujZVhokVwn3Wt/d1F7NnnIzbhDspa
0PL6wrFRhrORrVecR63YvaZTo316hxUHbTVk50HaSkRc9Yizv1ZyxDo6i43NOcJFKoCQd6SFNQUJ
285nWvZ8X+4QPU7Kx81tUAV/y8veZg5j8JxyYF3eduvljw4Q74gkSPUmziQwk7aNW3z9TL1gDSUx
XlN/47TWrGKbfsTc2ZNSmcRf1ViGAZlIdDc3zYrx1kL7pnSVuedJKn2KIABXsvEgAUwimO5caFk8
ZftVj5xCwrsFOTDYqrR5dlRlJAsFhiUJFZDXqyO4roTS0uBqtCiuv1fGzkBqx0SMxv+NBIg5tZSt
2U1D/N0/FFAtzZT1d8/YukNLVviYQS6wRUbgReLWf8367kynOp6ejUmf2XQWq/mMQYYz84beIWje
x8M/Sj8y2H1wG8rMdJCnB6YB9l7GyxMTvy+ALHryj2l4WLXr6CTXIjHqxEy98xNfnINzJbumVNf+
ogUw79Mv+zTh3Bvo/Z33VOcA5Vv+R1cB6TgQD20JPcrUtg5GqJQGjQ8hi32PLRH+ZMZHzw+BDS+g
YyONcNPdlgp0AY5C5HxRRLL8nDK8jEQbIxpktggY0fN2n20KT+cS972L9NdzFlTpDCR5F5eDeLcJ
Wj5AIfFds5cMziS4u80kWgYC6X7ukYJctM4rbBph3M8vR37dWlzTfEGABqwEj8SH52JmiLwaOrre
LzhZ+WVsNIufnDena8nEfJpNOM0u52+zR//YvB0ku9bGm2BSCNQGtnXyDq/LLpmhdNu0hXKTDlRk
Kj9TtP28/isFA9Wrs1fQkOgm8Ih1G8pW5sT+bg0inGNJy7UbAcWd1tsdATZEaj8rL+mVUPe0fOtM
BgxPCY8YTnbyTjT1XbbGg0KO+n2YthRt5wmoymCLllFtnXzyGRSeksp9XWG1EjlkZMkWuKyZEIIx
6gvTZCUZYv9oPUJtQWSTOAH4Vb0aaLZImRop03YJJ4q9wq40qaGMRaKFh0dtl9fg/+lK3MovRCiz
rNLGpEAggSNflfkMhj3qMhYBX6cmbfC5eAfBE8ARwrq0KzuetzO6FG2e5vMnlMlvULRsIFl7v+dt
2mMf/O6ws/eaP5uI0dhcTjdCQEWIovL3HT0HonrPGx/ToLkUmDx8nIA+jvfB5Ey/VerLf1CmZdK7
0kq7F/Sartj+vrdxgg6QHQWHNuP6czflxFwdDk6umFRxDFMO/PSUtlqGIILGgjINQoCy408T3WUX
prr5yv71hSg+He22uqhkA8e/fRqrOvCuW0EBTRZ2vOUa6sdV8rxGZAopAoO3sdWrzx8cLBwYSkQV
mrWiPi4pl4LTE0H2Yhhqc4Ks0nQQyoYRqHwNzgJ6xoIK64E1X4zkemVksx2AKGzIoA/sB8gi/7rz
r0sB8opyKWhe8qYu2B9sO+px5s/xH6YR5oW0d8AQ384UpWgEx/hzgeiGL2WdPJ+OMFjTdSsUuxYL
2WPgkoUJ9wYFx4zyGNFAYeL6sJ3rq5gqOYWeQSKXpqTmUMYwNNe1U/4xRRJzX/qKy5Z35xhWnF/A
M7TwOVIAL+4RhEGF4ZBgTQO0ahw371cl+H2e/ZuBrtIlSic3dM3wfawZRE7RMSjjakTboBsc5Ajp
Pj7sXPNPiqwr+wQyMBGpXjWc1pWfdwQZ/VwWXcH7gaQaZ8dn0xW9zWVXJWzA3rg8/0Ypb48MrwJ7
6bIX7J/n1R3Xno0/Wb3QDIXajKkW+rWZuTehgJ8RaprJyXy47rq2RRImve20ocLA4D+JAvJAl3im
/tft/MGEfK56TjCbF7USZHuo65YHiwXX5ATyDWuZ7/BZERZoSAHtjMFMo7/IWUxcYut4YwXqTRIz
44LOyfC4PZN5cvcpHHTyZhv/xmwxm7MfZI4i3vvapiYKLTWSmIlYjJ1ut2fceEjtcnbOxqHKWcAb
/SIBxrWIjyIV369LdBEIwJz5lmZ9a7XNzzL2XJ2zxCMlJM8pDZefv4IR6Z74M/1qrShyjsPFQ45E
8AiwFgzrlagjbNLWyw1ucoiCgdlz+NpCUqaYdywvPN5O+K36Rbe8N4EeiNjDKAC70wgK5LFJdzdJ
Ill+UGrOHEUkJwlLS56Yx1dYGAiCiDL4PfSxPzufHFJYFt9wOivnsa2uFoHP0jbBkQjnduBWRWOQ
XKhS1D+3PfX4mJRJgeeUDwngjLIPn/yOpj4cn77saTvdvov293cIMPu86TqkdCukUretS/Q4SHqq
CbR2AA6qlE2BhzZ7ZNZPgJAVbSacA8tNYTHgh+PNRJ9gy2CA13Y+y/MwcCYhVJZwx/apjrhYhdhA
HT6dn2AmkiVp8wrtkKZ6PIE+0ovCfeKCR56yoEx1iFkEhq8P2PrbGtXw/XQiUD0FipNZJ/T/HXor
gULlXkPebIDXR69gQY1Mg5YbhsbTH1j57Vgwnsdr87lD3+2iJXBc9Cp+x4DefXkyyxC4UP3lW41B
sPw8Zrs5aSOnxvjtGL3uxGKsaEeT1Knq2woFub7alfNKl+ssj644kRK97g47zZzoH+FZh0Jg4VKz
OHjOhFB6ZthA7f2pEwMb6VDFSFQKOZdWYhZH5KN3D/O3kz7y9o2xJioG3BU+vYbdz9swPgJVrz2k
LqtH0OxanE9ZEn5psBENwfdhAgAlAIULCJ3lbr/3JnFtGUqxZsELr3jbPAqaQUj1299yn3KkWZ6s
BQlWYGrVaGUUFKXLRy3EnoND8hpx199CQ3j4sh6gd6radZLmcGCKydRDOMNjPMg3Ae9m4cd3sBw0
VHm61pBKAbMWbQqtKNK9d4zQogaUP7xI9ZpSUZEbfcCdBcL3mgaxK92ZhPnxSZpWoFVv40allBBB
by0c3lcKLwRo/73lejs0Qq70exwMdZRll4Po5eW9HLMTqxXAocrNn2BHwJa32ivk9m9DWWRp+GUz
T0CxzTFD+rCxUkQ3V+vpwxgPaDnicPzax28OW5uYICOhlKj7bcl6Rh74T8CwNMkO4nNHX1LmT0Ob
BHGTKpQoSvQWLg7llWq2HtgBkkAyWXE6pyiHLUiPF2cYXnUl4q55SpqIpVeaQboe4KDccKXGnjiH
AjzTjOec9UQqfHdmt99BrVlIE2wm4QVsUq5G58fU7KFn46QxgbBFdMw4zAC3ysQdbYVgJf3sR2Sc
CdOZOkkQBFRCZ+WXDf/EFsq7XZJKd1swkGqv8VVZ6cOjx6pRYR+6o1v3FP2RtR7q+PjHhJ4IPsw9
GEsutrgS0vir7ztAQQa/7wridxsVOLCpC5IqXoO4igaP54l2M/rFO61SvBAsmEapmJ3epR6zKRJu
mTLEyjVUrQxWDIR1S2v36he+OtWgGC/puuEy4NqpFx8anVG3pDVQv5Jg/wyPGDigN4nAgn4X2WJk
+cdqUwXl/jHSVNJYzcu0SbEAEzTkq+HAKwys39qYri1hedBLBipgcWtfDfik5jljfHNjMYciEwyE
Af2d6YqQndHpgkoSQl3nvvPoijudQcBpQtg35dF86vWcXEq8UGwAqHybMsT78Y8t9XKrdOSjcQyz
kjzAfzqDYeKTFVBKL+Yei7vd1eCu/4AHpCski+bZXgEDNKvpKBa9NtG47NTRnPJYiMqzpsraJSBq
M2hJPg7ZznLKglCxnxJwOa4IsYGiFZKVTbkX4vjaoXbWpgfueHADXeHlvy4n0d1bhOrPH/+9cGln
ojucosbjrNnSBwlcir2ZplxlQRt5ggYzEWIxzOhF+SdsWarM/oLolH3RjSjk2E6hADcNuyPuWG0p
qnQxG9Yl5OYuEEp+TfsRMcYmI1mMROLsx5odNMEbPFrYDJ2y/PBpJqUAQuZY2EKeM5x4NZKjLq62
5yJ9Gcsz11KvzCiqTp5rjnGFMkrzNr0AhGGxyN1DUEBqie5VAeQ2Dd14qCHuPCbUBO7aypjVvG74
RvnbbJgIp8zFMBCZMoschZ8OqVoSaf0rd1DOFlakUYPPMnJlzFzjHHq3KmNMRC9G9tOFblSjdKmR
FWh0jIQb6uxCOM9smRG5OuS3ZbipI/bmNG0XgewBt0MhKUCZf0ZgeEiwLMJHp0u+NFa1aruLqcmy
yDNsITAyDsX/68y/fnxoCjpEmMceSwnYIawEkvqEAx2xz7jsz02uZhOEheXXh1iGwqw2GUrw+gr0
eSwWNFSTw43zyX4sJS8m6qlgPNObcImgLiFo3bqcobZ/PLWre5J9E1qm9Cnr1bNvtDvNKr9MS3TG
eW+2s4xwLaQWDR/K8CPo/+c83x/Nt/65H0TzjUrrhk4bYVMj+RzQzMqZNgAgjHmaZe4VBF3NS1Us
5Fl3YHVdvQmwhS47l/4yUKsjPBRZw9wnJbCcOESwsD16i5cJCEEWjEcTvOveyIlUVKJTCYRHC4J1
pyKvzcsdCaHWQQ2xGA3Xb/qACq5HYnrIcnFmoHzWFWsmoxo3ZCjWdqn95iTOe/ciwta+9yZ6In3x
L4cw9zxTmFBOmXEI68DH+dVe49hgTZbHI5fmNfXu6914oMCfc4MaWrW7g+PSwgNJano1x+W70w+S
CA5T6/T2LhKiw3K923Mnjlx880klHQ7cj8OJfPqQajeorNjpHYTm1slgM96p6G6JalQ4koyL4K/9
DgcRlZayTpt7qGsaaiLaHb8c4aVRLm0jcUlrQ2MlCNGyVyNc10QSjgl5Po2VNmGEmY8srJ9yfZiv
WwZJYS7eZtXIL43Iyvcs9L/JtjjJQX7s9aXih3fyU1AEvU4Ckj/Dr6eFGLWf8mYYnTY93sPcYe4h
iM0bWtqKwOBwLr7D9kylXDziXgHYry2tvS790PM3eV+xXoOcMweqj6UTWWnwST26wVUl48c9xJRL
a4X/oJYDnMiTM++OjngwA2xXXdPmEjr2cky0l7Xh8WEJxe/YJK0yKlrIJSqqnA7BMtVksBru/aB3
ZdKBcBsx3lnXmQmVNP+pLxPvSBEI7q60YCbiwbBe/XsdLe9F6LpLfwl833tqB+rbD6zpwhgFb6ZN
4r4IGQJtM3bbrrUleNifALnCB8CZip4r8wL4v8tn+DGbZFxKp8zw/BI7G9tm23JlEyeztYvsRGA4
hS8G+SgQ5l051BGvcf8q8gHMJKRuJvz8L71jzqbzqD+UVd9zNDaxbdpdwTCgPD/DAjOtUvp/0zwo
xTZsaqySIa9/qEd51jURFmjsHo11A6Tmv/reqbmVRWQBLwaSA1w9fo2Q/dDv0aBdzYHuxp7Ynia9
q2+0s2Fmj9LGQNjGAQEGhKFNe5EiaKQ73eq6EtLydbiUeiQFsXxP0unEUSkdFJCrUU95M5kvq/R4
LRtIKb+Ae+HLKCgR0xQDVyUQJwIdCaU5vX2k68gOSm96eVhT08VXWumwu2TVbZ/MRWnsg3Y6aLhi
LHqszP8psW5GVHcK4WJD2GZbjHhi06Jp3auu/pKghpA0wdjTk+TmbAI/tstQTr6JMTmZfx4UYCVq
RQ47GS1VGpESF4/DQcdtjGKu4IorUcHwPPrbCHTru3+dnwH/8jw05RjwweuV0xZY6bBfYbxcLa69
BsSNRqNAAX9xjgfe/jN6i7xBfMd23uvuvRdAjmbWHrLwDhWA5E8eqD2gBWknMTqxqgTIXLOFB6Fk
x2F7KmGS6t/JAc0pXKJoDAwrJSgNI82hNNpeq9W6TL/qL4Y1kuzJ7VOzVt2jy+k11gXOQU+gfXjv
BySbE3ZQsVDIhE6gLfQ9VTPVaNX1K8v329VV/GNACGh5t+8R+nerx0antaSHJvGyLXFl1rTuSikJ
7ZpmJFPAdidaSQBqL1zSemnuVU8N0KsqLeByd06zFXI31hyt329wB/HqCUEXGKPAJu6MCtE2oe40
6sLWA79hRIJEwKngk8c6E0XmHX86WcGNMAJAO0VGFuILFG/VClL4fIz0dFPU3sJMtG7iMnertGKM
Gpv+V/7sbxZ0IdQme/PJaEzN8lSjJwar6iY/VvaQbAE5xBXCoq3gsQ9AeSWLWZUfXYJHtNpVrJKI
/2o4bXde8ro4I2knUJAk/V4F7AWIIHbte53IygvExLikGIhx1CmqvGnw5XeGlzXCI8aKj4brYteY
wZP0qMK0pgdeIaKG0FMmwM3fLzJ82yW4+pFMJHhiEpOAbLZDJm1MOYeoUtPboMXSF4wZQ2+48Wbt
bPYXwNfoeyw85i0znfR8MKSQnhPPnL3egoWHjqzTdjKaMrjNWsxDkLNCRS8ckhUeVEjTjs3m9F+s
EzMTady6g+jlqwdQ3ksXkhUWD2L64IqmOyRELCX6v3GulS28GMryj4bksW/6782xbYbTUWMR+8Xb
EwRVC0WNTuZ+H9vvLa2Dcs6ZRTRzX7EjGMZfyZz/Uo6YAtun0esS4toRnunrqYdosxYPYvLwT1xD
TMQCIdS/duiHqQXNb8kmy3+42+Il3EkNPrpqhH/7/0CVfQZ9hwLqruniZrf5ugeAtUd4Y0lCufBn
kr5hU6fdPHDqWtApIr9qnQQXFy2zvP2eCxdLXHKlKJ73WzQ6Ho7X1DbHxoy9SGeETxiiw0qYZ1xA
cTGlLNI41iY8n4bJw/Uq21Af/8kPIS15Nb+/KYpos0K1YND9bB0aCrheCTfETDpOelKgvqz2JSHT
F/2zJ5dPbq+IUB1o9EGel9AMx5BhFcBo98pKhtmM3TWWBywg6zAaAWi1vLWcJ75bJEgHJHBlwCJL
2r6YX2DkUWvkLpCbYuhOHZ3bqEEFvaENlZ9uvTOUrksv7jXRY5ermV6B9GbZF165i6Y0raQtXh00
HgkRMjh+cZh4o4otRjAjsZHdj/NdmzGW+wyTTm9waRsfrfhbFHqyKNIZd9PrwZvpFN8ohM1D7CvO
oFSMkyAOTe4Qxf04xQLt0JGr7swo0ymKSfF64JoZQD4k64XRe6m36BmR4b/kMa3TmaCob4WF4fBB
mMDxVxkcqVQD7fmabjDwyoSLH+wxPegTmRi+bTosWnRtTTLkEH7PQPx+wmK8O5DonrA2X4RFTRSu
yRb+CFWULsgGjY9AfWGPQWKVaGVVgzgb4+ksDeY5SATVrVw/bmbL1wvMzMyjc2GRUud2w9j27LT4
Ckb99EAg2yjhjWSn/5hK4foCzuNC8KdwQg/bsuTw3ttQaK0UT31zCkShiiaTXqyzldu0WHu60uG4
pQAPwY0sIzIPhc/AdAqmgzkxl3dpYQ/VamW3Cf9f8mEakfadf2kqYFbo/lrhwuxpBzm/q0LNkFHQ
FrYtch9/+XLZ5rcSm46rX9E7/TeiHkNKak+8PjTj4tQwhjSK8P2HMVdYmPv5kG+AxSULrWaKSZbb
Te/9bNUolXx6lZQITG/PCElYlpYtMArPy90uv+YbfofW/SXDQX29azLMri6W1Ff+KdOyAnYOkhb8
mqGboC8bAkBXhX7M7Rbv4Dw+io/WSkguNLLTsTwaECakj5Nlb23srVS914CoqDc6mSWUMlE4uM29
jPJZw9EKWBKcxrfw+m5EoYLRU9zcyp4DCzx0JibW0PsN0bUQvM82ObUchWYYuRYds3KCed7kjBlh
zkpPTzXjJTsknu+W5SOurE7O+DAcOiGgmGCw3nzdjPsQrjoKS+tFznbQ6Javak7wjywuu+vSAWnU
R7xNUOESg/M/pBvvWLQhZQ7QTvH8+2TvrBpncitbVbiU6bg850e1QUM3wQeh0vNKWywAaFlfQQpi
6ONQ1lealsK/0EuziFbXwMYpFu5QTSrhjmSQk0mlzfXTBpiW3ZjGlzaN3KhZgdOAMZUIHZIfmK1A
flSpAuYtWHODIOJN4t1EmWFFSP4T2o/HJLQAoYnces1mF+blQbcGr+lXEvMm2CX3oRz686ZJsbsX
STYkdj1PRZR7d1Zi2KxmOmiEm/MmKgeZ6RBYQzJF4k1qgWfH2W+FctMu+z4SBx2ffI6FO/M3ICMS
I8Y1wuR3CyfBsAfgMjC08HVp0G4q95+BC1+QxkhmMNaNXdBH1EPhLii/eoILmE42EAuEkOEgB5HD
CcoRn9iwjV/5xN8/91MRCi0IvzI1NbdFl5gaJt/PEqafINKD3O7I+rcAhzKgiYMAPUIiFd8zo2UL
lDj70UZbm4F1C9xE+Q+ANpE00ZMidLhUndL1RA/RJ5kHlIubzCIUUbqpjDSIZD3fODiQ8W/YPQ2T
Z/MVjWuvAkdbFjpoJLOYX7q+3Kjhv4xgrerULLzkP+vI+uxKh1BZG9xtLGl4u07dOVBG2P9bjM0N
SETTK2PLbvJqKSJw0tHFMLhvNXECU16Hgn1uTh7Mcm4ULk53/ODqthjjw4qEjNPDjMdJHK31QYGL
JbLkeb1vSWk7CbVIeOkjC1j4GkRz1CnTwzmWfYej6wcDlCBZi3msu/m9xPI7TIlRNe8dVQ6H01EB
rXaezLhH8plgBCmeekvnYXroVhxML5HZgrEDhJ3D+dwjFxyp+oJe8lrJI1rjTe9s32QxJ2bQhRZk
vQIBK/cpjYu8GKssgYhr07L2M7w7v2emU/OlwSzQQFsDrv8a4zpe491j6+9aEvjjZscanSSwgk61
yl2kYWqUA1YovQiuNngF3kFZLQwbfYMgZmyI8dehjUcdIvegpZykxe59VS84T/UQ1ocG8lTnhvOr
t7/N03RJGYbdWadpBwlfQzuTk3bf91gdC4ETj3izRY3v50c2QdAfJzR7XgS20pHBgavwbQe1aP7B
4oXXJ2evyV1h5y5P970s6/SSskTEUhMTzR6uz91xT2oZAW0fkhu1H+WX952GZz/NRbeiyJDeUD0W
Bm+Ex8gMTp+GYI5EjzxFjHDsztjbahIzVkhgotA2RuxhsX62h1WFKUhUzqrvm9QnKswGDQvEyc0q
XX8fUK8nLhveZzpzbvEt+wvQskg7Ax/r4f31EpKYTpUF4DrD+UnNeZ94B0BK7LfjMrX90vTp9vmX
VKUDvi/T6oNBZNQsCrQ0DT9djtBWObAcjvlTeYtGay6reZ+AxMtkyNk8CvZmtj5N61o+MdHn+/07
jKe1Usf2Q2pdYFOCwSoOMhBPBpiT06GBQk3pvjNovhz9UsPDBE9/W+mpqb9ziaRFHQg/5xuqPMgR
RfTm0mKANPNRq4YJF6dZNJzKtqvccI7lk9ryPXF8oiBUof0KTUsyJLIxU7zl//SNm6OINhld7wOx
SHK1cjNAAGt/qNcoFEZ2PtNh+c47zXw9gsK+SvZQsP0zUGSeA3IXspUqwTXXSbzpIA5WpLxUpgaz
uHsMMd1mAR6TYNPu7Wnd7qrMdrbcx+f0XHL3czo0EYQFMim6mquR15eiGcWT08/+oaHfN5FgQqbg
mwqPiJW9/KR2awpdhHvuuUveOnw1RmmJPENKgGHNuctEVqkpSfOvL+cuU8MoiOYc7OmPVK4bTol8
HViC7dxFSsBOPanfIusL5XCOyKuT+wgWeXIlf6PLesr4BJ84hRhKD2P7xIwyW1MJyb5L8Z8WcJv9
qCZOs/LL21KaqwcVZmcFQzYFLO2TWp/IKrxoo7EeBMtxOqcZl2ueivU8Tv64ZQusWz2aDulQR0rO
PVpXWXskVEOrGiFZ0e5kIuXQBCNhSDsVTlgPp1fvgBNcoEOu2Yq/F9PDQe90x8+KxxHXrI2JznVa
NFsmO1lTB7GPSPBzmpAexVJWBg6CfvuOyKTPkkHty02QSJLZlPCEc34Z/edhfTI0A3TrJA9dNrK7
vjbsXHfQ4PYYUpfpNAFqMefq4x4GF9UYz4B/gaNurJ2zkKcU7qnMjA2tCKF1RSnrffJIQidmzl/G
gPkDhwQurA/qCjv+WL4Lk9ECt7Et5VN77tNVdC/TaBKyM7aughTGmldffaVyOE77QpJlIay1Q/XA
CbickSS3O9DUAdKt3uBSYtdpID2SI/NCzytltsgOL7m8hxLcKVYQloyskGy5yctOnwjyo777gWQW
QkbP5cou+C974XvuLcFoPfsAUsVec6Z1NamPOmXmSiNOEk/8sz54DjrL2Pgio2vNZVKO1V0EQR9Y
znEdeTNfkcUW1tTXK7GDqIWOj1aRvQi/u0RGkEmV13e/jz8l2mrF4U6bV++qktVq2ian1Lcx71vT
uytxgVY6S2+C/gsdXPsumoCMfB6HMxAs7utJ4GXKdtjESjOGP0wR55aILpsTIED6icMTERHhv+4G
Is9AC4ZS/LBepqCLjclvI7VLJ9zAUiDDkgWX9gmJXgnWhQs2mht+GmVIWjhv2COWquSb/2T2zeU0
VlUn1cS/+6W2pVWlcTkjRILvZ2FQJKqbTHVBnpAm7OLeeoN65JJAeXFkFOvn6aFLlDzY+Czp2p1i
seSEJKZIfMncysc2soVgiy/kYTFcOEvEzCbcafFsoy/LvyNhdX15LJeBJCugnxecZYDSqVp3A2yU
za8vj1BnfouaKY9sZMoJVoa/SZAIOyJTgTaPiPd7ldoI2zp4/TqZw0+evK9yS+C/fuvwUHPJ1VZh
hEgjvk93Dx4POTKzE584yFcj3b0XiPaLnC4ubq8ziln7yrMZz6DcLEn4zjGDjTJKrQQVj7UIsBJ4
n3RKZgH8dIUO/WHAxtaLJEdOZtnu0ggo03/F5M1DdhWq0+MkuFS18EDnEJ1oZ47QcW3Ftwf/aYuV
TrdANW5caFR2Pd84EGlc71+FR7wvKRVsPCeofm1qiosi0lnahs3OYWYs+KnvNDTc7xouSEuED7n1
ZWW8trIiiX7ENqBT2XhdiKgxNkEALsdolvOz4lIUzYbBlz61WOz7CIgTQ/n9qx/P/PRf3nXx5i09
elzem0YPjiGD3A6qn5FdGiA7qn6jtCRAelIS5diCD5ZtnWwh1xyY7cK/+5YBkM8bsc5JHI9FBjIC
+kOH+5HTelUHKzptg99ApjyuO+0iJI5edSo3E99lcxPjCUtWrOqbOScvv3FgELEvGvqmdKZxSU/j
bIsNDKZYd0HD1e/zGrlL3ujDw8RGOBOW2LBJqPsOzP1DLAt92zHp2zhhGe3JOrEcnpabqW54AUXO
a/x9FssL+4SLzSyUVR/nLF/8/R3Lndt4m/WVQSmmbOZXJMDmNBWBa+eNWyfPW5klzX6vQJwUcR27
+gJ5JFIuAp3Fz2Wk4HHlVd3yvy9bBJEiNslu9pCqnSKcHLqRSuZGG+fIdJXKOn+AvbjFS4sAKYBI
ArHcJypJ430cCGENEnCGzUO12+7jNFOOIdDoOjl0k3WofKc9k9kSulX8LfReb8wQy9DJHzIY6T66
7/1LazRkWZPk3g1cze49MOt5MVN+hpx5O9nO6CqQTOgsdpkayxt7ed7WG6/hr/S0752awufYdn1j
s7WPzuQm79wnnkI+SN3NOxmfwus0te5ISwOQouUIMNT8DJdW6J7m9jFcpeTghQlFxMJrZTO6aBMY
A/4yMmYJiKX9Cg8tPwnfN+ECBsY00t0iBxSbbAMcITLTsIEnhqPJaeF/Xl/rRiRZrwu4W0upRZPz
2Cv0Ac7BTjJO93SxU2NlYAciuG5+YCrhRWZp3Yhk+8Tpo/2rDvoF+cylVnGZRS3vAc57ZjMc//Px
0zyzGOCNcL4nzbfGa2rRzt33c+DokaYhmrrYzoUBNpMwZo4MMCcPf1w8FZKC5El2UHFtoC11qkFy
hiPubWtXWd8iYYtbG7aQLZbq8PelCan5DUqsM2ON6TmUL+6Nnan8jH0JtnxEGfynqQ9O49Bmc43/
cBWKcNHanHfcOiXqIg2MMreDX1QbUjybexGFFS8C94yBklxcOrKDwTSWDrpLDdR8iYEhtO+DNG7K
RFcALa5N44880I3eLXhT4T58Gr1GY/KSz9jInmmQHH00UzNkQZMXVMI2+nZ4EyCVtO18m/WPfAjv
fcBYfH4QeU1e/eQRVYsJZ3plMq/mntdhYmawggn7muRB47fYDiKmemJep/FPaisOZaCOWjxmOUps
j9itSkcjlTstiJmLJ12cvLvZADbkkwW+tjQ4gH3Ymsnds23fUnDF2BuggG+eqehUNfEQGgQpUaoR
jnyt7CnSi3QkSyJ1WoohMMQRRtRDxC80kRBmCB4SqI9uTJEj0N5k4aQaB75gO13Ya4tX44Aa7iNS
tcz9669vWVSpR817pa6Yo9du3RlYuwoTQlhmt2sKN+dwY2dejW48YrMRGH5QSJgMn793xjOhuup+
Y7lvN+ileBCbngBd7UHU0aOsyg+RGRddK9l4ac1+17eDwS3aDkJeu4PzOsyFMojCfB67lCKip7AY
/+MjDwqLbzt8GClqTOFfnLfMBgm+8X9VdGSTzsr+Oiqxu/cVclNyfiHmpXfhdEIxzVzKOmaP72MH
wZlSWh7TXMtMkr6Xg6hc5BbPVXx+Qb5gRgxORKK/vYg3HTFJcP4Tslnp98zeakzD9diNpvu5BCqm
FvJn/P7WjOiZaDFq26EUODUltkPLgI85XIZYR7m7aQJRFEOdt+UQWBxRJIs+cUxT1AmzKaRfwMwJ
Va85AeG1aV924XxhbosOq/1o0fGgiFBE5TskGhtDDD4i4h+5r7VD6ZJi27wArH0Z5xFuS4E0Zzl/
45sb2oXx/b1AZ1lhVzj/riwvd33Ru4G9znFMSNIc2HZNexehy00ZVDh18RvRn4JhRkWu9g2acCms
EGy4F41f/rIc+fDbqFoak+HQhebRSb58Ceeaemj0MPSC23fGPuW+m3ZJMasXEg/t4JYCWQ6rnrQ+
V8UbVK1KJtso0HDu1rvwr+Q+vZDfUg5cnCUiF8odGUUXMwirB3vMoZd5hAk6qmj4kvhCZi41zi7J
HGCTuPRoP6pZeZmk0w9JMcve3tSrokBENjHdfWETg1Z6XACfLezOLyZJKssrGl1AukHcR+RCUg9B
TFBuOAlI8UAaakQgvDsJ1I5nfl1ZHyyr4aoBd/s3D+URGD7BHFyebZtb9bHTu5Q4V6VTKIXQE4n3
H9/0dP3lBag6rgOHx14pPzwasCPkNjbINa01++7vTomwHJb7V4yv0xCv4xuUt5NS/GNPvP/Uh911
qffir4JS/wQOUTREjbFMHIIjo9vOOP77TQQmCs5uoilzFG7EdhwQO4G9qVzfDXY7xivJcsWWQMo9
t4kwdJNAMAGfzp38mJpuAlJPrnZ7+0P21R26YJ2FsaT8LxGmhH2F1jxcyAIBdEcoPTRISGawlf0y
YGtiScg/NRWBqWEGwSQDa12Pfs/Ek1bV6qjr6wBdAj9FDZ9kjeUdLXiUMQ/HE/sdLwIT5TK0tJ2m
TKxQO37rRKvr1184DJ2Ed9w/1TjwNmLqNJPgRdG28Eg69AZNiLCrhL9hl7wZHcr3Lom/cnykhOYf
7Whg8f7DoRRfx4Knjbfb2yHi5I8eEYJ1of92mrkWXbI3wQ4GtehqbazMCQCZXEiGdqIKivDWkBh7
5Neq8Omu2GYZWAlbVVW5tdJleKPZAerENaZtFOz6VrGnBfwwbHrFnvvUZea4HcCsjwEYqKp6Vsfi
/62/pIFF1vS0M+5a1THAinCSi3crcETSEd0YjWHREWy0bgvJxOFUgYHG3NtfR2oFo3bZFm1URyfm
o3KNnIV6LJbaBA7Ll4tQS9hEN/piN/h0lr65wzQyyb5nJA39QAZXN8c49k7dFAk45ah9WxxAAcG0
OQ6Q5Spz4mE+08B2IfqvAbmqj47IIE49LSCnSc0Z0/VUddTToaazP0fo9COz+Xr8s0TMKcUjWZpd
hhmuUSmVi45iihK2rfVPtuC3vbKGY30vvxu8LyT0zEDhY40DMoy1TSYrhUd3wFvi+XCSNFinYtQN
VqHha0h5O9Woko1No4QeRkgN81ysz2cRNgtEWNG7hOb0AhkcrrXx6fekBRcN6LyP5ZsVDnL9cRCz
nn5Vpz0QXBIkds99+mHXVVixOO1aK6cFvYwx0DCflgtSmthigf4NTbO9wl2470ayOrbUaV0D6Q5B
jRFGbKHDNKmXJWh3+tBAncGMCApPqiFD+kBiEjSQYWQnsBMIlCGRicRaHQAMDYDW+DwyivMoiiHD
KwYDuTGhGcssdGFtqRRwikhURehtz6N6JqFpw/K4GMb2PSCQvVCibzrtbgs02+MLdbC1NaXfzKo3
h9cH5ZOFU2EN2A6t5Uniyy1/MRfClAqCl996SA/M5K0MLS1bujFtXpaFQmyG2pTgJRflACK2lSQT
40lEBLsat/ti+xaX/xCTiP9muscyQjvkG3q8PCaxXIQa0zUQszCm19DQU4WOr3v3aUQaEf5WHCgD
bSKV2ByDMcCXCCypSLwM59VuQW8nsJiPDZic3oWBHQfGTyrcqnA299vZpxHGyxeStuXFunP+07QJ
pshNEujC4SoSiaLXRE+uZOgNyKAfpxgLyN+FP2j20OhLNALus+jVvIBVYr9IUx/eQErCB1SDBOzE
oh7JfOqdKuXnTFN+xi9zYSdf75EVXoZjsDiP4vx4RcFif8S3H1+zXy/l6boY5K0Ff/Al3rtNqj7a
GoybWq9ZrseI4SwgSB0aMTlegMQAhUKggRwG4uM0Olqn+rmWOfoi9dR7KDheWLvKVI/ChHFoL1sE
jv0UI+OQpMtKXQ2bT3Rc88Jsfsj6c/eeqJxrx8k92aZmnvgW5ay4XSc5WLIhgTIIGnFgx8+X/NAY
jGZow58a1PLDz8r3vEl/y2cXJWtWltyZCxJ4k9stIkdnfkSbSXpLMZLDeb7mUH/n8UMc/zrK9w5I
ciFL9cDztfC+8xG6KLnXoMRMwC3Mx6jHpKVGm7f3ztmhMNPPGNZW2EUZ8knt+q7cUPkESPooyw0i
q2DhjFxAiJWWvLsfYIHA/IGSCRNZSsc0Wz2yHrC4IUW1DPOUPYhzuugqQtBWAdRW2+rcHJhAmSdK
xDKLmXxY83O7AIKdN7/FenJC2gKZVY16wyhc0ayaa+5Iz2Fs7mvbVNIxQ9ciYYUrhNW/EWwk6yLL
/Ccf3kRiEkR6yjNDO1lDfAO3EBK4Hcd72JI3YzAoTAw0cpGWNf3S1h+4JDnE8GLfhdrKzBJR29TZ
JbbDh6h6g7QQYpMfnsdOZIOpgQL/Tn2QWSkYnkAzlA/tUMBZoJ2+g3FeNN5ezKK5SGRjLreFRGv2
g6+c++N8nhZ1guKYcOmcp8LGuZqIIcwAyMhp483ikW/qpphjENfClOuMfr1QC6+va8CmLmHsKIPr
iU33Dwb15ekV9OB1LpvzVkVUiQIqj0LyuBt9P3jaIUZ1byZWzZ7YmDXBy0pPslyaFV8Op9mg92Jm
1NnQtc2HiXbUofpnD30lyBKgGHF1PdJ11z1w+85dxoLfrpml/YIJpXT7qRMlRT57BZhYwYJ26dCO
XisTeNBTryCDgkqA1VAlmKH5Nt8/GijDPfgpzoTWmwRB1pCZzzwf4H8L+NawDuvQ1apVOjo/9No6
3fybsSwNxVHu3UUOAudYFssiRLka/QdpEOm/e5XnIstLIa4W2fy3+XvdjU+WWV/Nz0fp1ZRwI2U2
XSeXMNq31cu0fr/OH0g3mw06z3oGDPAGejOFdLWFSj2khNwVvcGvW+a+wr4zzVVCsgSpCDe84Lz7
BvZ8GQnVl7CCRGLCQ5GgreUPQRBRg1rGMdyg2EO8qUk42CAhGv0nO59XNfCrG1RTM42xfskIcXwJ
7ja0BDskXqqjt2DpUy3dUFWoZDBzvnh+qRR6vBXZh2jMAsP80qaVxQoKc94b2gCkSqAuyRkubnB4
AM6Zb4HKnSZ4YPUE/NFIr2Zz0ydQRyD8ICKCewRQpZvcCQSoX74W76sqgeYOKHQbZGrZvQyRSyLP
p8ekQ7aSQ8iyahOHMIVsbFRZHqfpFtkduVdz3mbhJA6y2QyeX/sMINbtAhCskQ4CAdFOVx0+ZsIr
zIwt5zpWT3cnHLQmXi5JJwSTV+pK4ZxxzuKKOyde986VIiLaPSIiwP00M+Ep/amfBBmLhzicAWKH
7HFzyYx6HGS9gfCwDlPhwhPFgZs05dJ/5fUifwFRsqmLfTY2CnRiW+LuZvracKeQohvosbGfR/Td
OKxKJbtlG3IZuvq7RzcBbLUqybDgqYQlhPLDcDtAPLCgVFNP9oUe7eQNT8aYXXT/ocz2IILIQz65
TdJHVPDuSv5dAcGssh6CWNZtw3voSs6C6KI1ASNwVy26z0fxcWbdwmIRQOkwGwwkavgUktMIlyeM
jCuBqC6wLdupbs3lbkdczY/2erdIq/elRPK5Bh5XkMTTWHUSbTlwCO9nD8V4uRTGdrehilYijSig
DppuKCxdGtvWJC7AJbH/eZFq9Kp7R42LxLABmllfExTMXffv4JFHlxUU5BXpnQ585l54D6BjSPdF
0qIGlpviLDL5gQpMsaRllAf+QmQ5Z5IoB+thgnb/NVSm+AiKNWHewTl3scaiAzlH7dvmTrUhyVvw
nsJkVXD+yfu4Rekx3Fx4J0QIFQK9L6xGXhez3sGvKCcqwagZJnZBjPzkWmaTvHuto7K03dcIGZ1D
FOzVdoV1QYVD0IXco/H7/O+nZH8oF7SQIVknrfuafEioF0bsx1dEfarKA6QJ5kNRbbv3F21+tRK3
SqLndww/X7otY9GycppNs0xbHAlYloMPEWuqVgI7Uj2EJUL5cXHJ0uT92lWYlM0l4hXNF1vjB1XE
mmehdpG5lROwT//sTsc2c5jf3khp+mzhbdIYmHjDrRhVDuE2UWaDZ5slSIJSz4vxC2SqbUTqKrS9
kLZxBlfa0YKCCyW60eimzwefni7BrQL5SZOeL0Tmg32RdleHHGGLa3szbz+D8uy4gjBLqC/aUtTd
6azM8GY/XVjhWZ26D0vNfD6AizdjCwbYyEICKzoJAXuAmCvvPgxQzF0JtwBysRRkCUrMYMPYRwy0
ltlGriub7MGbK3DPChEKQI6hizIRMF09v49HojMRIU4weYZkquaUqXnpil+UQ+wVAvhGRfYG5f8b
A1axMpZ84vmBqAeJCvDs9TAiV+ApDmAlmx+8s7ei7MqzRH9MFvmBYQmTGkVDBGD+934DV9+AxKPZ
UIX+450cHcL9rr/yxYbf9Qa5hFptcgYE/gobr2eDD2l565XK2QhcAE6IJy4H/arUw1m0MpC7vXG3
3AN89DLO26UXRgJj1MAObdQ122vpOySSIPWO7cITEZSKlScopIWYPqF4SSGOzqowQaYyF9KABY05
ZuZK6KRr21qq/uVO9EUxTrJD8t5CeSDjqaVEPaPEQV/h/qhQ3GlCUSAJc4SFZHSJ4AVPrxospDY6
YNSu0cn95WWy3qWLg3AwxooMn10ga/8kbmCsGkVwtORH6KqpNa2Hhprc1T6I1tCqSKJoNaEl12x/
5w9orUGAFSq/jEdl6wwjR2voBjB2AnDKu/HjAUWS7kSs7hyFeRqQm9baPY0VkWMlRNFpgkOeH6WK
fYVmWJj0XcRU/eiiXuNDu1Q2gguIoR/qt2Nq80azN7wYLY/AtBRtaRJgqSj9XvdgH/zoZT470My+
SQSq4U7YXx77EhU6uYtB0EkydZiUXJhKF+4RWCboTiCdbI2j7qCeJ+76Yylq1se4gLCoJb58EGta
+6q/EFEhoNPdnCxRT+OVCX7j/BWIobKoUCl24wkG7ryz2MNJEendvPTKo9MbFn+GnfqWgIp3biCY
VxnOKF2gF4eLQ3fHIJc9+I36mLQNGpHmRDGAqw8IOwQb1EK1H5pwe7LZ5ISjdMYPzYMWg/KeJeEn
6gGkq3G6/xFnbbdB1AnP2xINYDnLYLfdiAjXc/zyMwpvmA5RYrjUB4FouIGuGc6moiZJLjIOjcKt
5RhVGSdJx9h2f2dSI0CjAwlr1JXtUAVx6BP4iMvGGDKVYLegYay+keguy1O71lPH2sn7/yGIvY/H
8HxxkGBDeG44Te7rBxxgQQ33lxn2w2j1fn7zOKa9d0nHug4txLmynT2PrEf2udHp8Zm5Gmx/Gl3I
JRR5GmHb8jVCGQpChSPECkMhoP5N/dGEIVxuyxWLfVZds4CBwFonMIYD1zNCRahIZ10EVu69NnRj
ysWsu5UeX/H4a5IzmkxPEfC6ubFBbjvjMHoMygh+W7NmznvTW2pJ1++Qd7R63u2TGJWBsrKpc+vO
uCC42LH5qmCAZC2vsLPXGKKPQXxU7NzzZhbXycX9pEk95eQZYvAIfEN3XwNMlzKzfFOKkDofeumS
8cvpQ0JYGeWzi9GRwlUGj2Apbj2qBv/+6f/z/QFS7Eb9zCot5/5t/AxK/iJrHEltR4wL+K4AY2vg
k9WSBH4mPwWA3vRO0H0/Q0BuNPW8Tj2JFOk4o+U2PtBGnU0M5gl9Z97u8bpXWU4tdwMz354Ed9fv
y8NZFCvA3QHXGSlLrBSwdHeNGHbCRU1MqWiGEl0njd4F8DtyDtRaKaItiPNy52z4x7kDt77m+iLo
9nPNbC+TpR9ePJliJN3El5isBHHehpoIAmnyS6CopmbTaig0UNSHJa6NiqT2AmNdsLCEEBXObLCw
jYBUK1RMEGjwomcX6k90IqW/vKtasu50fG6yNWSfso2sRaUEoDyFqGoMQ7Kyp/VyEHYVod1chYaY
0XVAkMlUSHTIYyWFilNhBMysS6zXYdK55IGnorAqLWAA09tHX+pkVoms65n/6RGZDjbDa40Eo46E
VXiNrxiVFvA0hBHNO5OeYee+yAWXZcsU9AUAaOGstYdecq5BcSjdpA00DT9OYxCX67/QviGYzqIM
8UOQWCn8tqnaDiUy87NB+k115hdukrThl+sKi7vPI16/RqZuZA7KGG4YuS28567gr1dpx7BKWWW3
TsskkkO2UT/NVUB0KMD0MnJ+PPDRvm8Rkr0Gws7CnBv2FcSaPCC9zXy/cIUodnLVEkKHpVC49p93
E+H6eFZm5diCbKgRrrr+CRaiiOJ98QWvtQt0NvRBERzgUJ+wfx8meKOo1Zv9wfj3ER/DmQuuh5pl
nJz5FEA8P7e3Qikts37E7u04k9rwFNx6qnktxkkv9bIXdDfUOJtZuIC7kWxebg+oZHfwEv+1Ewc2
v3db6o5Owfvt5+E5ioD5IeQioZEpT7+8adzaP8e88Nmw6+k0zq/mEuZQPUgEZ2By9+h9HwfOGnNf
0aRnsK97ArhGlTopSlteAzZrH47nAzhwqG7Lh1qVBGMy4KFkqjqGGDjvArKd5cbXG2NphtMg+u5F
RjwvdpRgg0tIa853oFfIEHDPfMCa4FzlVs7lXoqYzzCGbd1kmqfQtGA1MZQywncpB2fiQ7N/V2dJ
jueFUz+JEwSLgm+9x+tHrrC2/Jubqzy0QLDpJunl0c3Q9NTj93GKBFD4x5ITYvQtQF+OkuixYG+2
CiX4zz0psqTJz6HyxrEuqXVkSVbAArCxlgNTxCoq3n5d/V+5uU7aLxrjPLr888a80zmtACq2/Msu
WKoI0CnJz3mKUUFpMUUDOE05ZV3xip79viKH3SJ7xjNHCmrkQGge6vID39Y3kKzpy3R6Mopr7pj/
0lM/5+IXnGxWiq2ih6W8FQH6Nso9w1jvsLt5xLCtoGGfFxsxbMMduqN2R2WekQU0fSHY3JgztzsZ
7Wi6xV7+JN0zzzkL9AaYN4YLfwQcS6/sE8eZ6zFeSl0VnZU4elpRKN4i9Uci5TUq1y+UwRAm7Si5
mgZ9Uoi30XM14V09qPZEzy3gtzKjdZE+0a5Zv1hDTbOKnNlLSRD9Q+Q38ldPG/APEEc7ghNyooew
gmjESi/SdB4alWIgmGM/rb+tQG/53HgqkVDVbm1Eh9TniFkGE5sdWFQH3LZuUX97tCxwX5CNh2aY
fDhoyDqEwsEek55mzbmkEpMVXLnl4//o4QJQt4m4vHytXi9BGDd0wppwGenozYgokAWanojXeR6h
eK+ZmeGAR7vh/w7tnQRQxgonZBGyB2RUZn4UWOxshFjYhAqD/ODK2bawxpH1j3qGr1Z3LqyDLdSG
cXajlY2V0OaLnFWx5L+1u/XEV9Tji1ekFM4lnxPGLyyN4TZEem0+LCf5JmvbhKwIKSuprVKtGKdX
Uk3Cp66uTahmQ2mHQYABpTUQgNWcvQs7Y/vGfl/L0sccPMtzjJyp3YHAD4mwcpPGLcGM3L5UjxLJ
akC2GH+v7IvrctqL2IGQBQpCdrXAE5qaVwwelVTIw/51RyFibE4oRXRjmNOFjFrx0tUVb1zC57ho
08ubltLaIjak9D4PWdgMGjMb+fXuJtXSlDzkvYK9iWcOcBKt9FiSkyoi4q2kZNfjciOu+1/+N5b/
/AU5HEw1ec4vR8RxAYGYhwj8zxMFiOnPHhdoJJM2KabuegFRxiTwoNuWc5deJQjel4QI/G76eFar
pcBxbugEWNfUuMLeMI0KE8YM9PHQnx7uCC/+C2NUxXM3FDn0vB/ZACjT00YX9DK8DQtyPz2ne4wP
Q1gxmT0Lq0ugGnXIomfGK7sggmGxeJIAvVj2dxpw+rpLjsacWxKpePe/5j5Zo1uENVZ4pt4Eo3xm
YXK2JpdsrIb4KtcCOy3E3uTvXCwkrnlQkOymwmx1zFHs5oK0EIB3AV0WGbFahy+H08wdA/gfJpEN
3a1jCejkdnwl8d6FBD8XVMfixO3bYThJbpWLfMcCPKjVke6A0UPKZWI0dd5tKvTJBlhZc+CtL4HM
Myio3Xv4wwjsbK4Oc0Yhz3qIQ3JFVSWvo8ibdxomDqPHLng/H6QPEpSwUZOhhmVFphha9aPvIwQ4
UsSjfpg+1zDm9k/gLEMl2EFlbngRpOAZWTTDy7EiPEqmEVEH69k9zGAsXJ7U7DM3oLUUvFH32O6Y
JTC1IBRZXvXQCpvQaR4l4nY0FUfSLlBMgZNXBI5gI3Pvp/L07oEk9yHeU8OHktRRltaxEvNd+HWC
q4HjK6nt2g73lgda49dgoAwgNwkkJTjj1gEPoOT6ft+0DxpSiWZ7RP/VpoboCzrW7a7JEbgXcCQ1
y6irStuT2pYs/UmOH1JLXWGAxpKB7RymZXiz68FNZ0ehtuhviBzO/7hsBM1cOzMjh5XNBQuiip8k
x4iLtrUghg+AUEUB/wi2ErUkUv2xO/KRc+rgyzQoaZtjaqcIDUaheUqADlQRdskZms4f6ohOTlWK
5EBhqjrKuAZ5aGQK+isvDeJ24+uCfHrVlm5t2/RPx+A7owZbGMc9sMp8VnaghTaIu8rKIFVYz5Oa
Y18LVTKFZNFq6gvlcpc46AoPbaehM1skXh5q8wEhz0YUmhu9YQP6bR+k1DbUK4og37H0BsFWCGd9
3zPYc674+PRYU/4D9GF3WSQ9709+z+iyDDxuqH1j1PGKgpDyKQS7t/IPGOq4JzwsQEvJGeUimjPd
2NtS0eZ2cF9gei4rzWA1DXXxwKMpOxYqS1Z8P8GXOyllFkE+xUBdLCHnCm2Trlv9HWpiGQ/LBnng
BXY6mGEwETffmNQ50xjN74CGVKFw3F3t9bjqmoIqwetTTOKz+IG0GoaY9nrvJoBRPZOM4TGfMBtk
avUIYGszypfaE8PJyoUpWq1zxvPebyEfPqDOgmEksUFkJ+w8mwrF4QNL2Sw6F0t4DH7PyYDCt1vc
KDNfiLwMvccg2F08aIjPy5xZCDGAKRTma3PjUGPmAS+yST9B2P2HvLV19YsGmT/luLZonxHuu5oL
5M9HKvEqg+65Fxb4KJP9+gPl1ftczENGfkO55DaTJ2hbTYbIKYExVUec2nbFWXFtVZ1/GNYSTZjZ
7CslqVVX618KKAQcE6OSsG+3Xkrrll5IXVFPns5pU5z5kZ9O3UGCpv8kQ2pCifv+CqDqm2L1WwKC
cbZiILTFATy9JYWBzSxy+txiqjtJopDNEC9aRfClyC9G3EqDvQlFKQC9IJxa3rjTJ3mUOSGrAX0i
RnxdvotcWrCM4dnWGh2QypDl8hCCSS5KMstmq+wYWGCCUBKb6skHWRkjUTtb9DI/bRjEEKtGf50M
wFmJkEEFeZVObXFo4TuxBck0RB6QWnrS8SL9qIvA7UD62kharCJrIXty5RnmztIFBVOQdLOvTFyO
oHwSXxeqRxCn6IwsNst7kO4FckkKrQ9NjDVhBBVrHOyr86C+jWmEIyJ5mNSSfKRH1hxVZO3OXdhv
p03sFEFJFQ6wgx4xwVZ0/2/mRKI/nJZS8RFgi4w5LG08Bc0ekCCz2OJhz3+6RWoS7wKok5uRiYys
p4b3T+3C9rWp0gFu7WllsZzzqNSiXQndt15ijpIfeGD/FHxT6SrgjXZ8xvJnnkmNkPYZZpkK69Nh
ugi58ymprNQlAUGxiP0hYVqOELp9opI01tE0lu3lW0pPfsNp65ngJzfj/xkv8zGM2R1ouFAa8Rns
JK4ZO7TTR4OhFVys9Up4QZX8SjT7u7eNdlhYviLW5rsnHqR4wrbKY82zgzunP5t8C7kCo2mNfbQg
4EBBXVnW2nVuVsOQn0AHSyjp81tWrYbZcmBLvtGlsxnhpnT1ic6JtIXRITeIkDep0r3gn+cYY0NE
n3oCJdJafPeI2J6T2JgYyALOSB1sgS2PXDXy5hiQo2ni9GFUSt/oe86m/z2giB3eoSAo0/z7kMCH
2kDm78nnyTOIUFOGTKz5vD97c7APm7GUCZR5QUCycNuGhNvsQTPnuEl1p+A19vr1vEnTFCHcXUNr
unUTFXFOwRHF8IubQD383PaBGYUryh3q+zD/Qse4LKc0VyqZR+r2a+juUeC6vC3MrNp8kfzsYlHg
2GU/C1F8K7zCG6dSUBtvvLj9Cwf1K70o98Mjx0xeQ+Abv44z0QbGZ5HBNtBcjgdMrcRWvBMyYVFS
C3i0uXF+s9kut1BEmUrxehNkAW6vZMVoMaw+4GHOGcbntQ+0wi44CKam/lmO5+o8lrFU3hrLUEoj
iU8fw6+xv5MvtLIwFWFzvvpx0B2FXE9RQq19rSXvQIxAox4A9gyFtmGULAS28EYMYRC1Frx0Aegd
opgCq2MItnjsw9J6B0U5l/fEBEzDaMLW9jXts7SZNv2Rt7umkajsSxDSZ5X8b5GCxZD/p3bOueoV
ypEoifAw5yg+ev/pJ5wY34s+2bZUMmdDxeMtufXzyo+SnedqFREt6qZA675m6l5aVQkYX3cqgpGr
9cfbso4TUjuRRvTf23a+oK1w2QvV3hv1o23Bf/GESGxJxBkeFthb/a9Y8U0iHQGyXMdmAXve4+wK
F6ywGt94bBv+5APbBX4zPCl6uTNBiGV84QyHwj2YWwvZeiGi4OeY/UHFwLUhPWgs+UKLiGV2i/fs
EdYjBoCjF4UlUsCFD4Rx89jVw1iq3WbYqCWRoSE6Rxek1WznPhuOq946tzffqk8yxRv7rT+Qmthz
S7CMKhxhJdKS1cuEznXALYYgbABl1HP1Zv8h1nZSA0ndXPZfSglq1cerYf6xy8SgPRS4d4bHkozR
iIu6l4kKry93dO8o89KxFc98nTqZluAa5adc5w+TSHVeN4CL370+/K2MBHSMyhXk1uHGCMsq148A
Wz2LILC+B787yg+fy8WD5ZSCs0XWdt/k3N36n6j7yKtwCVEEJAZ1r+Fm7dHQGj0LPI5yFwWP2UO/
vl7Sf6hI9+PyVrGv7fi56chLnfxfO2CJIdFvCm3im+DEep4tIyebtFD5pUYKA7eiZ8MDq2XNxFU+
Vx7o1ddtlwgxvPaHpvCn5qQci5u/l1DyEEPgwPElark/0rthk81cC+eOiD0gn8t4uM8DrWY1vfD/
+G8mhBCdgeq9BXqM9fOCZKfCQMcnONCFquuMzpVeEUfr8cIAuuQ6JKKPlbcxHq24kBRg21Hy/h6E
WmCHoyqJRqeQkY8cBxa1SaZ0XX5ybre0Y7qxfAtrruax1kAEh6z1tNB2/iy3U/5C5lYNiJinhZiG
6D84wMVQ+CEYX8gpbkgnqjBXKLAvA3Xc5uMrGPfj4fkUeQ+9/QW2PqSGTyIx/xbH5kGlKt/g94q3
k2V7j87dIC7juiBOHZsDKXNRaLE3Mt9M+UZh6RkTPeSwHDivFBpqAAHvRF/NbTPczM/YzCp0+xVS
XyWRpXOm8XrEbD5rVWgzkYTMvovRS43/1D05B1NnqbhLLY7ltyHaN/8iRQDsvzsyr95t1wVZfR1l
zRv+I5mgCm+l19uMzYVguULKQdVN71Yx5gxKQ1iLfXDZsMCfOrKccwy3S6LKiLtLzN1ETlNdDM4i
1GldfzY0BGustVv08K14OfEKgCeo2SJSar9iA7mzl4dXR7tlGnzueAsk9B/ozNSE7V1RPfF5rjdy
EH5bMkF2IqdLtigTdfAepXMQUfUCdHNKgJASysq+oug/kxpCkaO1HzGZXf7lweg91MrlewFknk73
DEVP69eqqE/j3z+QlGe/46fiC+UcbAkRDWxm/ELlrBABOiEbRxhF56YJkr9uHblIjuiVLUUZaeiw
ffpDf/CsQiRUl6VOxzaUwMmI8Uc9Uzft5IBAgFNNsXteoxklMQxvILFx0cqiNT/QB5CODL51xjzo
YTLKw9HDwVeClh/wFBaGfCVN5dEuBgkGn1dzy66fDCi9USIU7pwfsU/YDRb7P+HpOHm8zxVY2Z2D
iONlMhC2CwDnNIrfg9uQj/oxFc4QWq2G6V6ywX8baFBwvE8FlGS4UETxSM96jBF4Ff39iu7ZCmyc
yq0FfFl3zh8G5eIAATRQ4YGnyui3Rx01S505uFPnKAeRp0hQqCT+xRV536ZHyCKUZVEtoJ8RELHr
eXA5Ids8uEVCOJR+DJYyHmim4XUDYNQxg9tjqBpwyuMsKrFn/zWQNWqmR5gQMVWb+S9PgRXfE3xK
iha9wkdFgDrVpeuzmsB7YnLGbe4GVpz625kd0al2p91TrF1qOl/L4/P+IkswbHEclWUZT7vlo02F
6Di31eLZsQjnd9xj4uwYMZ1kOanji25wHRRKcwnndRndpKmNnEG40AYjMLFm0lKhcCNbj5vmZ6Oa
mEN/eANcCbKyucDboOVFFgL5LFErKQXXYqkzJ15BFBFvAmYLRmhVA6UfWF1Fi4LIR6C4hSm1AyoM
7o4veQNfKjh85Pa1xEhHJwrVkZf++ORxYlKuALhWpvUkt5xlHPNgR0wcsCtIg0MryG6ZW3t58/5c
0jQjA2+bSqwTEik2bb4GJ84iyF0SG1M+DLEQ5EPR6/zlptxvGkrz6g03H2foAnlgQOk6wOaqSXWT
3FJIJWXWy2Sm7uhkHxRHTnnFL49TGHsEs8n/J+X1KI4biFq3EFHLv3CYy7VHnShq7xoRL/G7WpCD
LBwzT9mMOANfmxUal231gCxPY72G6eiBmENZ7jCRe5okWmv03G9HxgVs6AvMl6zwX8fGGlrl4uGH
Vrog3i/d3y+Xi9OQ7y6mrHP0eEEkyymTW3DPZNUWmoC2rLB3ttJo+YddXjhCLR2lzyftXdVmqjNf
RuWz935bHfkcnfEmpbz+xBhU5yoMPQ3k6c6B+E5tccjxnEMvUb612gY4YiXlq/Jeeh3AlYCs/7aP
niS4ovtsmvHp3rmn3tixDZpmX8rnj1HHEYB+2V15RTiUp4ImzZP/WmIi4Gm+5euHKBihw7rhxr0Y
X+LIZudqvGpXob4fzQcSn7qw8PTLSPz8mCafw7BNOOPO4fp64BHJYROcTlv7t+9SwW0V3SqQoMWt
kLKA3FHMfUa6RPZxHiRiC/Zs3RGAZ5ckP7icVJMvLehJISu9LuszfGAgzE0mlE26OGhei9XqIQ7H
/QWUXJsCryadoorLZT7uoU84/x2kG6XAf7tsPfrlS85xLlHVlXhqTvqk+sHuXhcD0UGdjbk51kWA
R2pULvIdAKukS3q9bPeOilP/UhrVO3LxZ+rywkb68CAi+Szhi8zEY/Lcpk4OeJFFN8fIA98yvd0A
y3ARLNLV16Uwh4f9/1RJVnr53jeL13J9sprsfbHCiX6XSUP89nCE4YxhZGqiVNZMm/1FSvope++d
ECyvn9sQN85TLo5P6i3TaIldzs3sAAlJnLBIQsBlLvq+eLjulkhg64A1OXqXl/r1NQ8wNSXzBVe2
lCeFHyyw4IvVEFHLwXqK66zB08uXZrR513lJHLUM28cpcEqCadpjvcrvSIahodJLouXL7KXJwyse
LQcOrGwKrPEnK3gBpeW6FYUgo08CQRSc0TpHtkQqbBsL42Qaa86eyPSPbLV74FYhklwOlfdQV2Hy
5aoSO7VSInXxrUnJNcAcPRXgIkZ7A103wU5DpX/8i1pWfq4atbWGjkvKDFmS8vuOFELOMMrfcncN
FIjfv/+t6ykjinuV4l1tsu2iKR2N3b9VZAAwGIXuCBJ+SYmzH9J6YjMiU4xOT4tflaGnBrVBLa/c
RriOMAQ+HPqvp7o7pz0m2y/Z5jXBfHa2MTzSC1RY8a3h1Hoj6DiJgluyFxF1GNoKa1joiejIZ9eJ
gTpaS+84bfx+GRQ0HT45QmzUUdJTudAOTag1s2iGwUFDOPFX7iM3GvJklhHw4DgxvkL3rped6n8w
J3Pz/mPxgIOa0T5nCScV0eME9h/HT6qNMnX8FrW2s1rr/PAhVUrQHR7Egsqu0rPLTfg0sT/Dnvn3
fZ0nIGiZ2u/dMpmED7zrpIgz1O4XYJO/hkJo+07ChupRhwkKRNh3+O0TqkI53Cg7DhIdXSnWPXkH
QG2/dDw5KVQLxgxcYIv3Vd/bEgQiU9eEJS8t2TzsU4RiETlO3BH4N77oaD0V6Zp+V+l8K5BrEJfJ
4qF1ggk/BnS+RGIxjqZLFnnNGJwyNBcqJgQqsqqpjdD/iPSa3zmKp4IC6dWNh6BcYH976afFGgTo
1cvTm97+BT3hPVjgzqiSfE9+l1nKlZWJ9S9gHnb3tU7I9k+OVIxFRAw/8WcGWQ+WoLmNdjCTUlr0
hvthx765ivf10DCH3e3RCcFIGpVRVAGvBSqdmq9HZGK07215MjiKZ6uuUz/3OUsFpdZAPJRg+kaq
+mWSycvgCSfXsP4sjqT9rIso2or2ttX3ltWtj1vHN0RTqMZGOPEhdCgMU9gG/s4U7Eju5q1vlyCl
QTEBP+FJidA678sEJ0illpzuErzPFiN6WwrX2XOltq+oTrJnJ/NWL22pEtM5f1n04P6tQ3x7vMU3
oxh0mpE3gyk83soSS/AOu42T1H/cAXUqyVRP0EZGi4T6lBYBkf8S0tSf68XyR2tvKMJegO0zryIU
/oYbkRMGx7No4DL0ZXNjxRSEh/kh4+jfxfCZREDrvn54+/KwF8hH/TOlqkXegaxIUMcFlctNKTG3
XGOQSudc5tzzZlRXJrqO4lgoMZei5SvzGvLCH4Mw5Z1Hp3w3us+s9w/aeeaz9EQEpvXmCw7ZWTzQ
YCPtG6MNCzQlD40ChKKcRkUKLgrXUD+VYKNalqALC/3dK2pTI20jezxzwOIbj5EVqWytpq9RV6XD
6HGjqOanWDWLyfA/ce3fqA4nFKG6wLOG0+jxbBA6nsBDMnmnrqbxVe7Lp8W2Lq1gzx8ysE/cjFRS
Qsm4TJR8Phug1hPc+cmesYO6nfTe5gX8mLngSQ5bocDgQhok2QptK8E2CEhc4ue6ezaOlN5hp78h
L8/JqdKUgmlD9e8HgD0XygD3WYVEhuvXcIKtTGOLFb2xvLEytgFpWCyusRihiN7aAdnMD2BSLma+
nHBU6YmcrFGGH44VKQkcSbEcRWfcwx9z1uUtq4BabkRABoUjjf89fvsxvAylpZHkbiW9lUdQ29bU
Stp3spM+IjMUwVMB8UFqE0cfEiafya+37OL8O1JNzqS/87WxOCrVSR47bCsacBNGLVDtJPczCyeE
JpXUuUG+o/2ERGTpNDK6c/bA7rNN5Qb3qPnve7gwiHv/DKfiy33IaFQnSTFxOZqz9cjnzZLOxmVP
wOd9yGsE4MFBZby53NhkTT1HYVezHsC+mC3W88+6mfIAFQnChzSqsMab+bujq/Y2nFrDPZQG1g+s
S7KGijTHPzoChpKS/OJ7zz0MNnZtH82TnN6xXdrCqs1Bn+4Gh/phgcTpeYkerdh3P+WaY17Aij/r
tCmKbJI+/f1BB30KGfgyq0VLNXF0+bynEWJB2pulPJQpR9yGfV/f2VAYTGeqJptvsB6JOXCqSzBq
BeVe6B4GyH9ScAwrxciomCToAkT9Me/9lVIwi8XmPvjLWKVybS9Ukyr3hyRhwiygo8g5szmXjBhu
xqn6ad2bIK4LY2+7jC6lC7Om9q8WXnsuA92tOQubq5UiPpIgqWP86o9dWxOtscybdI1+HK2DCfs4
fyJAUc+6U9LzEV0v4tnfWA16tGwnfTWOXOMikvufdWgc0i1odHS2sDW30MQhCyO/NvVTIb8hpa6A
2zmCRNqBPpGM8CSz8aPyCawGPtLR9FL4otmBw/LMJC8O8zf2v8qwIRDVSce7cHDBQtS60NBHPevz
Zxfb7U8IcGUuAWDVELmBrqNO1Je3bweET9F0th+vAlNTGFjsQ4wxjcxNnZ8TeXf03II/Zgsr8u3j
phaMvo7uaprbBs1/ZsshcLZ9opBCsY9GVtOS3KW+4flTWqa1l+Lq2j4jDZIu1fASI4sSg0Mvu0XH
x1JSI6XuswvkfdRfn10dU+/6us98+ZxNLX7Ndhtfta/KR/+GqRe3qr7kMrHHcRANLc0oFU00BBN3
BRtgkDxSGXZ8YkHdnIZmb6IrDqYPdIrFAkiS6QbMKTB5emGFcuf41pCwJiontJQVEi6ew6dnBzno
n3/aOZtqweHUGRgRP65SYEhTMWZIA0gyz6Za/5aDLIHUjtyfttrgqWi7gycgZYdVPSS/BXQj5swp
rbjF0ivto+dLZV0zu3e5PBveop4C0YcQQ5JBlzxtPoVBpdLyY47ephpSHg2g8ylg2eUXDDzEhgi3
qRbqu89tU6fslkbf0gE5PAaRMtviIZt9BjKuhm2+Ax9tpN30TLRir6WlAuwtauMXu3c6C56gG7qq
5hOz0jua/07HSrre0MSQuZWRkQ7uQkexhV3PBHTaHK96XOQSZdyQAYEs9a4+U1N/Qk1qeMz3PKkD
B/scV74HP3AHYAQXarx3P6A/vUjjygARLV+uKhTOXEIplw6mw1YXLKiKN6A6ycWwBh8HUk6CKdCp
J7avnVkCDre2UskS0Nrot92ajj5rtFJfvsprejWOd3t5vv6HV/wrGvBksviGsxcEvTTYYgj4uazs
BTKavkmYzQxWcTqb9+QWezIcZG54hJrNYcgYqJLg6XCI2UR2t1n5Pkm0h1pWWIVy+LfNBVpfVYWo
ls6UGgKvwcQ9aI0GkSDIpZhVDjbiJLRKaMs1r6dqGGuhqKUaKz4vBibQpcKcZiKNXiDvaxI6PUHn
BdcGa0nvqBjNA4ppPlNPNk8ySr8PVDTUTfnxA9NEiSG9+X0kGc//67i2PfkU6+UN0kZBb72ZTsD1
gw5ZnksR6zmrYQk5mkXCaVApgVw7W03BMX5rUToHhVmR6zNf8/DUtSJNv+ILFu64e17v52Ny4Olq
eDTWWXXZ+Oc9de+jc6WUyowmseHr7wmY3dze6seO8vXV1n9W7RdxknULj9Szyrhlh7zYFAIbSGnu
lLqTAUu/EA8DJVXSW2GwSykw/TAnh/2vzzvnpDGLGXF94FUEoSrO9akaAecc7ji1EvFK27Vxd3Se
/2h2JeKZvWQ22Yt6vJOqY3rLaBCon37BUnvMacZvZKBEWYt3R716PXrf+Ks8Hy1NwMVCe63syxUb
hCFPUMoftrkpLm6BBWdTjYUmnWLUqmRyBsdTVaTDU1dnQyjkzxKo4dGZpSfjFY/AP3Qa/TrezJ1g
ock+WacuyZcfSMoO8Q8pDo83JzSRorzfrVI/8vcQNOv2lNpdt3gTrnlzY9m/kJJW5SP51+CvGL3Z
GNn3qZd9w2gLRyWBtbBKJnN5SzYf1zzfFGZgQvMciVCmoTn2WvrGOd4OjgI3PutTxaRX6uK9HYCx
5K5juMMmpJz4EQKaAjKG84a94/fPz/hgohcZ8NgyLq5si2N60zq8huXtSlWpwFy/ag3x9auJquyP
PTlnAfgov/6fkPJBrR+/8TthFd5sroy4bD1GqFXItT3socqkZm/hshf/TFjfIyHuEB7Czo5qg2sj
larmlU/uFLwomUOGd5UW7Iz8x5CUly0IwwNRrie5tOX6Cs8CRb/MmCvLEbBrUSEOUodPgIzG9JUq
vKuPx1zYHvRIqu6/vxDvayMKF5tZaHvm+yHyOS8x9hcNj3PfUwmdHbijcK8co0gPHoJBqwL2RumG
0nWSPUXDVw5FOr8UWdzbpwOe3GhBWUq7G2IIdXVxoLpvoy17df4SY84YphcT6alY2Hqhk2Up3aWE
loJ11T6ESMC7DoeOP/qZ+9SLpGTfZ3/SQLnJbtNv16PcHLtW+esn65XnXkrkNrmIc2ga+WzqnKF5
YaMvWBUdnmaMsNNa9YH6c0BwLD5gzhx9pJiaj3cDDKSrD9GIF3Z1xNuBDkEL7ycHElMG/I6YjhII
gbKP/StaQnMS2RMqgo+dV2I1V1j0AC5XadxqCnwScUUzXEekfk/+7tv4srMeUzKPOp6xjNbv4m5r
f1HM5kETwXleVww62cjhmT0WnVq5NXelIso6DNUhJmtLLI67Toz4Bpdn6+i4bITuEBZMkcVbtg2L
lYPphd4xVLkhBUujYKgS2pSMv5F410EGgHZjNqp/MI7/FYu1CI9lUAENyWULh1Qcws5b0PZtbw+D
e0PUynay7ePzfkelckRinu/geOzhPiJwFyED48xX+8zGVijjdfUcyxeQkVRhUPFBshTVOqCzdnWq
u6l3g+k8JL6ffepHgtFvrngtBJyxAKGmeO5+W5kng/4wHv2tYNdOHZh6JjhYVbGNH2rgksTeyFm4
PVcGPFCioq+dmzxNkWTFt36Z+OSeT+S1FwJgID4d873TTfED4c+xS+MSvSOF9BeIPQ13vd186E0j
uNJP71be1C75BL02XARFDddQVRqnlbFREoZDp6QFrBv36GcbWxlNMUrDkX3a38W0n7fgjjJsUsXG
EyVb1ZeNY7TiGkSdcuMQ8ofUn31GZrD+zdLesRTCQdYMNFTl7I+t5acYDtw7EYO05WMpMsoh49BN
/IcHIlbhi4JmECWjbODbkwM0mk8Y0jSDgFO3pmbBozo8FEBAeYQEP/GszcjPtZqfKeRhYRrgd6xR
D/vE/ejzkkpWVhKA1+YKqhNa8vbsVw2h7lTT92/P5wlxqPK1t206Pp+u72I5FVh0KE/irDQymx/m
mAm8jAgEFyPePfd7fT/U4YNBXUlQJvCkNQToGxLsocIjg81hVftUORM0zRNGkYu5OmKXAqvmaybU
3tE7AxNC05y4KI54xRrHyOIPMRVoXZNzc6qSMunKUPWX0DTCGuceh9jApbMLjZILQexdrNUOvON8
UqojG63eKOGqDqxHG4AYUYVtK54IsIQDVF+xoHFajVATjWKj7tBJGCt4BlUIZvasxK41b2Ytna0v
S6pFwvyyM4JCfkLZ21+BG2Gg95bMkY70TAnWaqMxYgdUrDApaM8Esa6PuzcLcsPIDaW3p3O+stjP
Fd+bwc4OzZZ8TzJ0EbFNJ/LXbPmr8bLbVmkTVWhgap7PGoPqQ2J0GFMU+FDyN9oFPYEj3s0Iv/d4
YzBPVC4zZrj0fAPhYTJZYgYy+UgJU2LwFTJKcWjaDEwO4CM8JPi1ibSD7zUI2SWV4NJxInvAD98+
n8LGHNrdvE/QaqQZncxtVvVlPuDjgAWAMYqrl44ykOhEr9irGBQx+QJMe9OqwOmg/EBerMPH8/zH
92BbXLHFjXRHsf1OQHD7NB9hfQ7pEBU1Xa0kZiSjmiFg42kvTHD/xfZacLDSaHWAkU/eMAX+/X4Y
MMTH0dryKT0VV5z8Ydx5N4qbI7PHWaArRtj6nUSzwj2EPhrPI0oV9iVXDDMRoR04iaV4BgYC9lJE
Tb28p8y6/eDVCznUQlEohNM+9jtP2GFWKMTeQSXr9VdaULXuWce/StFV8haFXljtVgp3ArO+X+ML
Q18PTSCgfU3z3UniFI5eqSzKNxy/dMNZk8q0ZqCqx++KgHgOK7F1xuOpQKXMsGglhrq7ZZtJwr/s
cZyEeLxj8dMN0gkAS7/fTcAxbr0nnM2hvQE8ldEvXP4/2mUa97FZQghk60RhXrLKaL/xsSxC/5wD
ZOpjJG9CTBVmCG03hsvy7kUTtpbMT6h8Kp9H9jLLdAHNYTgiwhwyHxmgjrvSjR5Q8yadnAQsxJXP
9HI4p1/X0SGwpY+bVvCdyHPfoqpem9AJmxo47A9V1S0L3Pq2n4rBbkc9odQ7uACvndIBgMRUlT6h
IfNt1FJqMUjzhEHPdDc8GO9eRVIJIyFo4szxD84vQHOQlpYHKFIFx9y1vrKUhk5/6yTxa4Wr3BCV
67aouWv7DHq9GpgvV7uwmoUjY5QOvxo81O1He5NJlGpGCZNBwax8b97f1M3NbqPtaxGcHC8+XKQz
FuHUAx+q9NKsRZA0x8uulsX+hu+QCv0BrOvsZ1mqHVE+LWyRUBYfO363IEQ0+fwN0ezDR43j36/n
iW45eRHoalb3LMG18XNpKIeWK2hlteqEp8pKOGCDoYbUC3PA6z09syGTMBH99N4vKQRD52eBa7bL
QrFz5TjglbdMiLSsnIrL5tM0O1PJr2Kuu0tqGXXi9QsXfAXU7sMwRoCtvZoPyfpoy6mNIilVV73q
m/gDGXb/+ef86ljLpmhEkWuglWFz6Lt1jvNY7u8+LAeu55tuLLrAcE+82w8DH3LmULH6m4t0HntQ
nS1BCZAbEbXcNwiCIVpgc8TWWCFU3UMZwvb/HPbRJUd3lIbND56K4DdJMnrCeXbY6rTk1T9KfknI
JyrEP3YZzEOu3qNnkaQvuAHIiW+gvW+M7i7NsEP1+SzujoMfUeJBbA3fW5CvcvohQDW4KCK5Kfm2
Kw3QRmI8mLNPxO7y8xqV8mO7Pq8LO9TOcr1tTy0fpqLbMKH0D3LvNCPo/e9J6DLQozDugyL5hdIV
/OQ4V5lf3ftKAQICMNj3Ya8ghhJwNKSz8twGp5A13sbS0L9wB6lKVqg6c3OwKbtAQYSrjwuMVGvs
Vd95COCJUnuoIkDRV8NlkZhKbqeT2vVkG8+KT38oKpMeT3Mz+5ir9DMT5/S6hsRdhTigu3CAgBKX
XD4epzC+kHWexwVEXqtJnqPRDGTRfv9At9jSKYjFBmCoTw8UbF/giddkUyfCsFnw9ORSXe7q2oPK
202HfmRv7Upt4NdDzArzYZ1520LP+p0nYyNjr9kfOTcdWIxNifitcbjPJPmkPoERZNXmkCBKKfR8
YXZsiW4FL8d2g3k5VOqsBMszEkzcAIHwa7+8dh7HDHwZdbIau5iH3dlgTmeakudw/q4InJtmfUQT
qIqLnQzYpvKkdOr8ctmZ+jDqz4OUVymA8BFQE5Mh3XHzMqrD2b06ZdRqa1/2XP2jp/UbssI4o6Be
cLwJnGikSf7hvAiYx+r73sOnOV28YECP5yDBHWHjvnT7ELfkWetXwjl22alMrHLaWrbOx2ZMO8yg
ngMbQPySHs4PH2o3e2ySVSauXfdYvCgbhR28tdfk2qcbYv2RKMEZHiJnjhEowIo/MJ+FHVmxcHaW
4z3EPgdmw6lThbHo5lo4TyD8cjgvF3cB0Lwc/HH3EanvfhsJO7mE8HdQ1ciB7uho5/2q7uONBZiR
unU7yiZ0qSmNLw7E467zSvkKMUcebCqAkxXQ+5Mz8hs/ajEgyVzjzDr1T5WuOU8+2vY1yjctQQ3T
gyM6OSF4Gdi8h01xFOsYNGEiQ3hC8XlOtoV6UDvtgh8MLbqCCMw/Gxopgg/HuRa+rC1YZ+zgpyQl
rTGeiygTDYordsPb98D6+gffOwigpk816pEx78He4Yo9aFwvnL0R5FrIAhPzYM0Yj4sj6iD0eE8k
79LEu5kE1PQQGjanIX0hlb6UR3MkiPPo1QpHHfozuSG/Uu3bdcBCFBVNGqaOX4fhfbkchnkSmcS8
CvSayLE9ZsLvDVQKnFgd1k2n9xuCGxP/UoEE8XtHsXZDJ457DjI2z5BqWUYOLRpNIRw6SdIN8EtH
Zk80AV32FE1v/i+9TeIqV2IvZqFUWd2bHISSgZndeBs9csGwGXPxiBvLPktk/S0queutbqlLE4rn
FqwiHgiQP0ZyHEj5Vnn/wTQwUiiAUcMSYMXgbG+bF2adkthdxol/FzLdRI0+0is9Wbfy7EDYZPcF
8bdA4HpGp3LR5zGkmCSNBsv+bpdrxy0m02uMUd3MVlcqTZZr7UvA4r6qFUbniO4evRUDA95B4c3w
nkXcyKKlFua4pBCiZKi7ByKT112YdUXMUmk5h/eisQ5/pHx1jZbm2JTxQRxxQmeekRjUV+7kfZN3
nnF/k+daAD8LUTsRa9nXtTkbSX4f4CJ6D9T69f6T+OJWpN3fQgLlW+Mmq3WzeOVsZkq2JbKztJtM
ud6EOz65g1jHmXaP6Y6dZju0vzu8Rjrn45AfGNCdPugnu78ZYnA037yXvFXONckhheVxjOVShZJi
7AhDPZyhtKZq1dVXqWngC4YOtR3JRRYBys2ZS8Sd05dJpXALBfYrRreF/Q2QCEACxw7qE35DC8vk
WJrvapYfgD0mMTVojgGM2r/ke1hjsU1GC2AYSAXmC5aRgivaDOLdnY0uRwyziR8GqIMwrF7mg45J
XU1SRA6V4/pR2Qz/IJfVGpf9+kBErjOFwilO0fxElueH+wHs3Ltk9GCYAp3IuD07rPrVVlQ5+Xvd
00a/Q1p9FSMT7xETyYJ0y5H3UOE/M810dF800AZU5BzwBcwgIEp2ChZqLQhb6FP8JrCtQsFnSswf
bdCNcZ3IKUnvn5q2Mm6mFApbkSuS5Xm7K0Xuq1bUj98ghATsWEBUe8fnkIHnnsMHRKlEDFuIt0nT
dJu7p8a6xay4iQqPJ6imOEwV/oyzNFbGixEMudHhOEnaEC3HmGfx0mamliibnyyHsvzUDV2TG3xv
bUWTH6d8qvNf5mEdYxRor3LnWhuLFJqG7lURUTJY5+klaYOSZF6J8SgW5Q83DTjFNQ3DOoCWtwux
Epq6EHryWBwSOYIzjztDFHGzfX4GFRn0inkAFioccZWjbRBFEL11v0aChz/r/1ifynjE9L/GB8tq
LxthxILo7QhDfqB6W4CdM5M73t+xHkwYD6Uz+DEHkZ8x6FkxGGya/gJGj0aTP1Vqv8tEr6i3lBTW
JV+OQLLU+p+PQbMVKt0xrH2k7J+YB8HH3YIeWZrLlrBNaW+I0qLdHxlMIFpwn64cCloKqZVIEo78
J3/xp4QrNjoqjLinxe5mh+jvMyzIo3laPav4mNMrM8TcGQMw0HN7g4Mdcu0qz9wNauXjmeWQVoMa
S0xO84longSAOywUYIZ7AF+DdNOQYa3q/Q04Sj1p6yj1lRihV0q+SkEfw1+pNTOYBeiXM1z64Fsm
nghcA5bfHT6e70t4b/e6Ub1j3KWvDgoMmc+ROBJycr5vNIgHga+SfeExKPHYjj6d5gdKpHXyEoc1
xC4iRGoqoZh4Dyl4dAJF1lp36Gz46n9WlMUIJrPnywIfchmU1T9aAaGmBI98EPvwdUj9Z8LC5BxS
HAaalK4L57rCZQnx6ZuYyem6rIY5tcGYMT3HZLCrFpnXga4R7jAGqnMOCFbkI+VtwM060hUq6FVZ
bbccg9VxuBNi4jTz0IQdfcr6MvpKYSGNiWibsOTx1C7QgHUkAH+olTUC+V2VolsylIcAd8+kQ44o
/kc5Q236jkaLosh7kx/1zvvWFLdVv5ktFlSj6UNI56BGiI6Nn2Mbi0ubxU92CDUDCOIFned8I/MC
7mb8qbr2DUHoC8T+PvXmtsWenUcrTkT0iDssGf2E/fO7c3i/6YphE5HC38RZh/2psCoMRoFehw4B
ZP7SwhCs/R0BWD1W1t1pap24no5nboAZjI/r7v+aXdrn2qf+ikxeOVbJieqCDfRJSLI2E/ZM4HHU
mHFpuX+Cfsn78HpQbMN5m7OXZEa4ewkMSWBmL3Gqbzh+hgZtCOoUDx6BwkyNJbEpiB+divSIFrte
3hbidwXX31cINmf/+DpffhXAsMaB6lFqcrrNrU14zpkjciK4qpcHjeu6K14ywjSpZsU3ClsleXEn
LctFlF4hH0QgD2DgrzG5cdIn+QBUTeQ3ZsYu97xTLsclLw/JBxbgaSe73kkXogyWdBkdyuVcEsvR
xXJaS+AVu/aNwlfh8rNvyAS1jDLHj/y28jtiSVtaFP2cyRMCl3lrXItb9n2+bx98qzZDqzZliE3e
IAGL3dfsI70XyPHbAI7yJAMVZCHFcK1px9OXno3h/iYxUybgM0E00UgnFykN+Jgi0muQv9qhIcI2
WK3kn315nS1IcjLA4RhVbOmt0YQb2Nx85BKI44QO0mHKk5N56kTw1ymc0Nc6T/SJv7doUECtyxAW
x+GVbmxnA8+4cdkEXjCsMPC9OgB75kXiePwCCCDXzlfTO2Mh1MyWvj+T1RC1DfQhM4tUVmXKee34
rnTGjuQ36SjlmYNUmJ2rE1wlcsQXLbs1ErHH7qVXgPAsqHMcmCeqO59v+UCAW5TTFKIxwLE8cLDt
zFa4+iScJABi20CrCuWQm0gAeYij6J084ui2Tla3K02WxuuJBkCZ3pNTmeFQ+6w+NYvdsvFaThAE
Cb1bcYW4DaTy1ZA3ctmXDvLZx55vnUQ/jZD3zEPm0OUuWeMvdEAZyvPk+uHrIULZc7LJKPjqWnRs
YaqrsCwPZIMBnjF8or0sCrJs4RYqdR5yJOLVCNUOCttVng4FmdA/fqcmXiBVuZ4d5ydey3ZKadnT
9sBtMFI6xw45A6ooiW6tBLYKV4k2i+mZ/UUXZraBkpJ3Hfxw7rVBwe6NVhCxnuj76JZEH3zMv5/R
ptGSWV1GCScKWZlJpqrG09YHpUxUtSTRkEKPOTeU8lauKtEH/sxskd1dHRrQKAQ70iK/7CvZceLV
3TqJZJZEnNHTsZn7enzn2TLlcF8q5GKJCA/6RPElrx2pkgz93UZunrdG1Zvdug7PDtBQPvKrdd5G
/3//dcDlHNVY57DDVBtSO3uRs0e7uBm8c/NXdyGIanD0J1PxLwmJRslaXgfPX1BaXYyK+0yvyL8f
XSuwGQY6gaPsKrBgoFLrJggOW/7AhdSflBDkjl+4skSR7NWPXWqfSr85efcB7fPJ4jZ3xEqKNm97
oGCir2ebnbr7XqcNz+dqTE23zU0L+2pxf/cChxi6w3PPvrJLN56/sGTjfd8ab0BEQNgU4Zqszl/7
IX3a4C8Vc8RssATrW9HtA5va33YkUXxxYRXJHrgK5heHni23Z1QEOT4vFkSWMR8DTY/qaRonxRZR
Esx3ssbzLMQXHoOlDHpAfOx/TTnhon3Jn1vai1L5hgk6walG+HAgVGZMMZb5wuSgMr1SfUq8eNDr
QmgVAANEwz8BsxEuFR2Ab2xAIZVbRb95h/IJfa7EZcE9mp8sJCPqsMx4CvUSizfJ9Gl2s/8wM2ae
FYGMkNo794C1KrJivaN4BQVB22p/Hr4amK8/KGiyD2LTyLZX/wZGah43/fQeIMczAJLYxwL3s9EP
8ytkH3f8WASRiSyWZuz/H3B5PoYvKIQVVoVs1qkPxoNvC2V6m4A187++xHzU9vtP716ESBSGRaQ2
i+iMPq5MMf7KptwKNmIeHUs68e7UZ5WK6ujl0dwyL5etd6BJgqEOjJhI8uH7JRVjrFc9kLnnx1Ud
TZfyJRdks8yupQz2Y13BywIo6DTBULPkYOl4GRZAsScofFdDhlbIRxVSVEyVrPBfHXutnIT4q/5A
1JHl+5mLajdkj4P3mkjQvEC45jzhdU/396rDGAJ+/ThFX1CUFGUkcAnhNayJxXBqSS6tCrcpZCk9
9zC1/hhuDjlT+50SENFUMyBqCLOsBPifr9FYLZkS7WrsBZTh2gfmeEi8mZq+euSDka+y1TIyPCoI
Hkmg6GCu9ZJExkvjJJtTtPKJzjBUXlglrKmXlwk8tLlqeLFAStjiQYVymZptAnQOCUU0NDTBBBcS
d6UAhcbGuUnjbYmnEUKq/1R0C/mDgnL4uJ+otRX5nTBlZ80pCSS9GZIgZjpnHBPL3Ch0asNya/zn
Zgj1YoIltGzqNaAPDLGNQkVps3haEJSUpkC7jkSVxS6BxIO3vbuLMdwtmoHL4ZCud5RNCAk5LZy1
jLvbMDChet5RpyX4AYC08bTmYRmUNg1SlDOm/UZHB5pG9BdIMW5dEbnI6qk1H4ncfZLPbE6zjbJf
8lNqhwE0EgULzpz3K8nodzpqgL61lTpjTyKLASCmWkcg0obsXv+4yUdGotWU2R2ZRDMEDfOq8QxX
agqHZoOAEyNCXPMguyHQBS0vLQzYoO9sIwW1pSTAPtEuhHJmbDon3wvgbIe+xEm2oD2pKu8jsYs5
uraiyVFZq1vCYmlPW+FEJNmnyJUgxRnBvrhWLvw7mHGfENUSzic5MsZ70Oby5RBjIibEEiQkzmvr
mwPqaC/9So7dU6o35XORWU7o7S7qPhCByPu0X2Kaym1DRaEsrOSSsMH3i6ksx617YikNEHAmSN3X
kSr3FsQr2w7MXJoNIJTpIb6tR9uPHzifvgcZ89fX9ikS77Nw7zFTUKtdW3RrlTcsc9H5sNUHK0hs
uss3J4ZUPA4Qn0eFnchFhgKqjxEaiLDA51Zu/zHg65ms8yySajtldoTCXp4JEzO3yZOJWx6ccxOR
yepaNHe4MUcLZbCKFJ34mswMo688tSmj9+IQ1dEVp2V71BbmvyMRJ1ka7JzOBUcxqz1Z4jrsCXU5
h/1RWjphK5leypFG+h8eGZ5BHDn5H4AmgESiSuDdLraCesbDr+R1k6U0PTA2tYz+h1WFXghkP9Uo
H0empHtna33uJtMHiKFvEWY45YB/IVaubcgn+fqzxbL5QiYn6FDO9ll6oh5tVij6IjTAx7JFnSe9
HPUCnMMTNYBGKlZRlpO/84xkWM88KetIh+MFULBAPa1zKcYH55MgM/a/Q1fhNF+iJUeRMBzd1Gwj
dQQ8xBa75oqtnwL5HmFql8Lr88ql7IgUVi/UtDJPqrS+IjGyMhCimbymxS2fse2Giu5JU2gQA/bB
nOGx3/mRUMy9NUN7/8B57TyORtVO6I4yZR/1QCt8t/6dyQPwtrEXQ2gSqDxRRpDhDXNX1CGlSmMN
OWGEa2kAwhOIu536IZ6Va4QkC1CS+XsKJPPEfUUkI5ie198VOwKsEfrMwYaj490TuFHw31BzW1eC
g9Eaf/DSRvsgWTLSeimf5+foEL3p5FLKADsUgjyxWTKV8Yvukr4UdGwJ6FpNcJlNoDqunR4UzgJg
YCtJOmz3dU5783K9zIr+OMhWi9TJj/Zk+OaRPtNsiIpGa1ZqJon+G33Wl1XvloXAN+XHx1YhaUEi
KE56AR99m1ZFf+wP/a8cU+scEczH34qf2wEmTWCkWYV7YaHJs+TnR6QZpdtfQ6qMQ90eENP+DdD0
WDFy7ZHCpMdXBFjpUWLxMTzaZWQGHZ/+UH0ODTVvIWS4QrbUW/9WWs/PB0gpVeswfky8to86pgXc
3M+PW0m4zit3svFqCrJZv1dttdwyhlwLkvJd/VM5iBozNxCpR7VyYB+5Ew7EdeoCFz6Oy/19EKe/
bNVfKU5uEyNrQnUyZDZ3HxhtvlADOpbWXSYNt5J85cEqNhWZJ1HO3rYfQgNnF8uA0Z36WxjTDlPR
EGwGVwRIys+WD1tGfX8X9/sBWmIoAqDCJMG/FECIKU/tuOfgJM3nQ/xRf/0I3AXWoM8RBbTTWPIj
IKzm4qrqFpv9Eibhe4eUw/JQBv+bni++WuftuD7wrvOkR9p0QzocCVIgSyIM8XGoYXiA2gQZDA05
RPgWg7evsyt+GBXGKNF3tmdU0rK+e3W5st/7erfGIfIQqR3TuUhZjzV69hyVy7aogcMRouexawGl
xuyDUTpHbWEpIEcCQcVQrqhIrpgR8X6jMmYQAcjzInCP8GKiLDjSUi8ieDQWn4bxVt+OQfT0YGRx
zXbG5TA27yLYOEVhwNKOucTgu/TmoacRDgQQW66UTz1sjKkZLobTlLo4Lzlw9IQKTA9n8Xe6QtVL
ZyAmkyHgt+7h/7qQLUZyZ6GefTjltuh1zhSxuxuoqC5/fo+yE/YvlWdD26AI32w3UqU3JHlHYzEA
J1JYFS6GCIsRzxVn8XCy3AzMxiQ8/rlWC7nuqAQ47qQkMqg6oQmxNLYYfmA/FjgbLg44c2LzoQWH
2GyQxvfhARgq53rhJp/5y8iqI6v77qDtn+D9O+RSUCtQi4TgarAnMt82BLFQCEPAX1KWbsJTf47C
rR/42Zt9sq4BkjbAw33O8JFhL6/N7wAoHMA8lIBIUAtL/lnAK1rlGlmvOYGYwUy5PkEJYqK2acKi
cYOblBv8witi3teAdW3dE4ACpNI75IBSPL8A9nV3pkbFVY+SxEBeV8k0VMFVfD74uPQJkfFi4k6w
nk8JkDKRm7xNUY9EDACi83tn2BNXmMWXWJ52DmII4OzW3pUwQQ7ycISIDKnqo0D/tUoWnUQffvXb
mFDNkIZICONTyaCXeuvB+HGGZzFyP/I1hzec+OpdmWs4Zqo7qKTAlm9j97eZQEhwnvvvXCElWSew
7gFS3o1Ipzvg6zGe44WrJJS1C+Bm0bqnuvC8Qg1dlt+R8R6FRnK7Zcn7QsjFyjXITpDI7YKbwlvz
9rSVcIJeaX7NKasT533VErevDtt3otOTGDFcgULTHvA4BwQHrnsZuZQPviFjacC9h8HLVq4u6J7g
R7xvNvVNCyhdZOnBR95r6uFKm6eYs0E6lcGd1kH+x97sAvtO2eHHnlI17MBDBD3GFbB0S+nzN1vI
V5tvxd1b+kxPHhnbJsRVk2jqDosotfGGw9s7VLqXDzOrgiejvOSdiIMF5qP1VPcRvnAQiexkyhVC
hmPM5jJMFN2HvaSv4qc6SYYtoeEvrP4SGR9WrXXhmGK/1k28XbF7J20q1c06DMxVD+p3AAMuSZUf
Ks6ajlxe0546k9YWd8bLUdYGjPjtjjXDAnDI99AnnCtZpnTXDHMD1q0P3j/cuUZew2jU60Yq8OyE
dfRugzn0c4H9c8eRp439QuyvJUXrPsqio0PEP4TKA7iiyTTY0LTVKFTt01cQgnBx9Sj9fupStHm3
rwiecUPhTibGVnH6ykktWip9rji/o41ds75zzzVcQ56l4cssUk45+KAlAcQTOMitphWB2WRYxnQD
zf6OBiWfJXVt7qalyS5do8FEaTnLO+vdgfpkZMrW7sBPKzUMGBwo2FzlwYH2cJ/TtJe9PxIRT8Ur
2YP771FWefKRJELLgvWFjt58tzGKs9fpHMxU2UyTmw0/4Cc6KyJb513JOB8ykRCGjJXHl3NZUv9w
iInX/nZ+HSlV+efwaLB47YGHYpBrz1Ano3IWYnkQ5lUkTK0Pz1ddIn9V2pVmWzH6tY7SpVyxWXfP
tyUkKCmUIhgOL+kD7px1LULHmveeeN1sLwqweTaqNOk8en6Gx/xMX1Z5V5t+SG6Lp7TLBcI7QNHs
i6qg0kUYpbbyualrd3mYUhr0R73M7mVbden6SXMou9QNL2470c+s7+zmVzQmoFFF50WfJMyrVClg
9cjJmxmFF0Xf4hK696uRGnf5V7P4F+3vhgvPQpUzbSlZFcaOla27fFqvwNLhCV1fuXWWSIqDee4C
/duYj2x0DPULMG134XsvL7FOkA7vi+npww6XQIkg8ZzKbz8e5u4oPaLa9jiZOlultlGPbduE/ZpX
XnyGIVTxsL9fAFlsrecvgkxfSqAuBMPE3kGm2tAd/+hkZm6u9rpkvfc+1heOz1x7hufg0swvbIPH
d/EUqChotYDM6ikDZMqGuuMMoEtvC7isZoSSsIBkK797fXdSyGqnba4bvqL8ihMOWvzoH8dcp3An
lJFpeFpRKcKGZxPYkC9D3/YoKgIWBXh9UmWTHVf0ItdnYpfubNrBfeOVGiLC5vQ71pTsGJxTEHqG
CVtQ50lM/+WEEJ0BEJln/hgmmulrjZK1U6PovBmXTp8yAAr26C4YevI9X6M3X0swpqV82br7CxiI
xEAYK3wG7lcqTa51L5k+FgDW2FjgOfWAlAz19GjfBLe6KGnwoxOWO8e8N8zQ3R+Ow/dbmyeEAGZb
A0ie9vatfH6wBAZBuzL28RadPtcDcPSeMzmOv3QLE4oTgd4MpDMT32w2lOfmmBo1wjkTobUISOnF
rezF3utBsyFSUqOXhNlclOSP75XpJEwS/sGwb01w19ZMx5LKKoVif/YbZeWtmK/wIESDu5AaWAhe
K/3rMgBGFkScezWKMSUBzMXnABef8ja6JQPVQF4UPGSHt4502vSG6j0iv9MmYc6HopTo4NA5uHQu
yw2BcRgISVq3u+9qWe8Ejxw9tk8oI/qRF9UOu/atl/SduMOnYe1JRGBMzWWDWpvKJqdtROX3yxVn
o4znRqwP1vHahzbMTZJRA+ejBt9xScHQHXvTo3r7EnhL86+VlwqYIaoYejGFUnS9cjIfT5vDLxhV
W7P54Ir5zSSFMVdepTGxvK3DdA4Ypxy/kyj1QM8ky3xWzP7KJrRjWcRsNI1TkIjTcSVCAzCm6Ey3
r5t5QY2IcEmWehUKmLbt1QYDKGCIBJaeF/1pxrbpkvwjQxnIV3iQtAzI/+pA2ObMxMlett+E01qh
jCSpFKBPYyyAENH0e/Sdb6gkBI93f16gu0QEOlDygNZhxW77GnChBOHiySats102P/hWAf/7XDiI
PYTtY/hT7l85KjomvdbxlQiFt9HL11uTuCUMd5c0XF1a63jM6Ug4YjpnYVK4VWSjgzLeJ0za6Nj9
9qDtlrR7rq0BLmHH7Yx/+FCIQrcFeWMUpQ32flSoAga3K5X8nB+4Ca3/Jm/XwR+YFKQK4PaM7NX0
JI9YelKCIIDt/dEHnypjOIsbHqi1MQ1QFRJ7sjPHpD9i+SjYRSslkI6pXMTQ8E65U9HMmjgR/1q4
2AHrkkdAus/WB458u7K2jlXqXyJqaB4D+V7hRQ5UEeUMrl+NhzyiO38vO8mqfc/wGGlCBMt6IbET
0ZZFr7J6qa5Q/YfGZutsiYVNvHaaWJU4WwLJ5QoWV2ognhwXsYTokIkiFzamGgoOmnAit+f+uhgU
htuy7Mb3MXAXqYqBYkNZxfjdurXY0BepD/6Gm+wD/VZO4JsNZJGl3Ji0NwUuj8fvYTE0vECBlMk/
a/R1OCB+6m2tSO21BFq4i8bf2tV7mfk6feWiyRmXbnnzsuDV8MpoGJyt7Z/2Lr0LZPJF0Nx3JMbV
FbcRyGFSexoTi7r4T5ZeEf7q69E4x2Tieo8nl4PpyMMkFCzM7x49huhA+p5kp1DsvPHHSfsNcLnv
DequSO5WpbX6cYTm1X2aeL74KKtb+Qb+Vnk/CZQc46yZcm5NCwIhZaPu+q2fJV3UaVSoyAynA56i
JcT1XO4ILSqgo5Ugyu8zn20XxpaCrO5AXixp4wcMiAr4M/UNs8VREFsoxwD6gZmbREXONuoF1Why
PViWxVV0U1xopCE9CtmKKVUWZ6xglSz3LcjZMzcNUdyn7krKmLwFr1exxcZO/PvlJBs+wyGKhiRj
iVb0R2B+Wm5Jj4pug+hPiQWHLls0hDqqywII2PzrLs2EsPDMXbgxkDe+JLLLUvq6ZOeIpXwnF2j/
z3V3NtZqkVRYo9j2zP43nTKNq+6ZUL5gdAfjttKzjeLgabuGDjPy1vR39HZop0XF76U2XsBQ7yYV
O4Y+JteLJxpm+jQNYmMSX5KpZVJCQgqDaW9np7MDTELL11LJEVL6PnBRql5x1wyzP5ljZU3klm3Z
xb/FcIe1IRqPG6zp25exEC1MkG09vkstYKsozfHbFD9yJz49krcw2CXjG5N529pqw/qi3SZa0Mkk
je1jjSJfUtFzmRQt47FyhaC7zzyE56odn4jYpKcB13fm5yyI2mB3wL2WKtP1V9IEHxNhlVp23KVu
ocs7CVABs2uSUkOxLMUZFkCwuwNxbOzVv4JJgVfqkTaZcNL2v8Jdt9HO7ErP5E+kLtShyldWRkmh
bOKPs1QxmiZsZ5DJmAXe6U8JZB7+sz0bNG9XQThXw3JiS0LmyypdqvOTF3Bpt+1sB1Q78zZ7GZ7r
6B/OEBTL9a99WTJk+b89k+7utwFUryGtH6+7Qu9HigpfE57jod+3H3oLasPN6dg7ID8k5pA8yRaG
XzPKxVXqtLx1E5xHpk1b/ZtezrfYwwOv8TO0J806fH0y5xM1QxsPuM/+J57w+eTVhVS5sQbXn5LM
Z9UOkDlHcdJurPU5ZIHe1hSX6/8chIzhZDiJyq14ynyF3wBAUnHAgvSK2NeZOWEf3y3BdnciCqH6
Lh+MQCyRj6ZZKk8VkYdELhg2Ydxc9ZhuSs+Uv/zVBjqlqwTFxSBTDAl9xOQ2Zsp/m1bTXynCa3DV
D4lTnEQ6hJhLsxd2RC4yHrnvpQF+/l+yeL3DQWu2THlZjtw1QjFdmHXHnI5PmuqJG9ZoditUlOyN
Ij+qQixCYPUw31r1eWbPwtWIw9cSirEAKAESn8Dm4EMf8DFUYFlfIVR33YQ+e79NOVUD5/iCvs2d
oQYzdLHWbJfb/KVNv90lXBiiLpWLBjhVjtmbqG6DKlSGO4LlOjJv82n9t/DwsDLh2OFHf7YD5xnR
5KffBnQpCZtI6SK0wr9enK6IOPuGxqsfCpwgg0YC0UD7eolEEegBexJQW08aaz01hEDy7zDWwc3N
/P3SA6wkv6FD79Yey3z3JKWKHWQGe4ndCTx46fC0nsbfxK85xgMhRi+PCzVKUXZJ2OFlvVySWX9C
0kWPhQ1K22NaNLiwkMmRnDm77RZ2XfXpscA0uz1WgpdNkGhDJtp+c3yhEdA2S0ygAdi1+XSZ7S6V
ZqF3Ti/wWMHlYmnkztCap24wilLcyCsRQM0Q1/va3b+w2TZ+xIIKYk2LLJIl7CbpYSv01QVGfzwt
+lmlUIlx1oCqQvv7QMaQcnYZ+TUOTBtpN3C8xeW52VRRdaisGBVJCv199tLL/zavKZ0udag+f1cJ
YhmUgFhAqmEfI3+gaCJ7Dg9PggUetCwpcmKIhkzXIq9mkepQT5y+YAXl2TxoynD2jEN5Qctmut7G
LiY4sVzTPqZTVn+SBDcyfbzsULRhxcaGmLa4n/b48mFra1Bo7qWGPjQhUVC63X8SrGF1OGyoocHN
rowhKmZbZ23vsEu27uoFBvcZjsM5hceTilu94FR3uKfvF0UeRQxpNH4nj0jQ02O1qXsWGdNgWepf
BTfYbVFXqlUS5zmVBBaBVUNZzK62FoQdx/myvecyQ0Zk3jzj/SBGVwhyo8TLyxE1TW+rp4Jzi8Et
oH14Sx94fgtdooGLxdm85biGYU033MMoAGL5hLgOPdFfPN3vWbxB/7DTMUqj0m09qLxwFWxmpW4Q
+qd5qPxqiT7SbLIWFC107kg2nhCj96TKY7ragO94Hgg9pcRMpUCdCeW/mMu5yLCh8V7aYU4bQKhV
H25CERGTp0qWwg54NgfMj6as7R5BR2uWzVUSlCKUUpkSSPa6sXdCHfmy34Y9h4zjXgIIPTopJyAa
mOEwsRSUlS0oe0vPcCITyFmBp87Wr5M6Vi8fupaR9umzZIAizn8hnXet3LN33nySaubrqJG/gcUQ
lBLKb3Oum8GDwY2NQyWg3a3c5I4ZfH9PJqCy3dnQG9+WVWBHODcRjfG7eLXRSTG+/afsgVDgytk1
L5WvNTLXZLoXYg9Od01nEkyS5ne0ONdl3wYu3you+iACTNddmrBIS7Zfiimv8sr7sCWJuj38sIut
0eSuvTPfBXATPb8lJtvZigIv4WmJyBVn3lq/D91JZRhjOaE1pZ37JE7aGnauAgiab1b8/hrzfMtF
ttah3SYViIEcuFizXHYOVDBVnN2aAUwNztOw5VM0ul36eIk07oSWD0GM9CvnXHhaj8R/LO+Tek9d
jeAUPMWF9xtiWacuVQMQGYzQxTcPuD5eCmX45Es94BOz/ZrN4Dwbk4WKhk4GjwbTNvIOePRemBWU
P3iYVqCRO8ZKRgL7FWDqlWIar2q9PXgjWObXnTDGx14dC8GpceRkVlPs6FVTJHIJhXeMUBDZ0oVY
ZUjcM0HK/7zNi69eOUX2lXS4JiamFm1lBdt4XIPs1FDGXFhOpZg4Ht0W6pHYyYQYjI2R28t681TH
uhieKMmsfITh89T71eF4taq4ISAKiveMn9eDPe9BXviJCr9NvQ24AKKcYciaAsebq9eSLuxx50RH
Qccjy9pLNmBca9DwUZ5jzFynjJVtKVGq6UsY+u3+WTjicpG2Lkt8kbz6/HK5GwK5bT5WSafAt9TD
Wpsxon/rXgLeWrVS4MoWkvLAgQ5A9HU4Obb4ICpuo28SnyK3TSLa7FVNmNWoU/eQjFjsbs7+CYDs
HEnxLDf2k6TGO4s5Ay/sOzBJ5/hmrUKm1SCXJFbU56Ugj0/rfsCZ09Ffpll1o4dIuxD9qvMMkVLZ
MkBbyJjaEo29FNsGGr72norqXIp388A1lD5bj2Iti8yzuREF2oCJa5+Gd/R2CA+sepsPVUiJvJTL
bOl+ZS7Nc7W25YjlLUW2iIGn5IhnMW+v7NyhCtrcu2//9/IlG8KON4dxxoL4BCQpWQQFjEBwPLNQ
800c5qZOLt7uroef1oCzYBnmAR4BoLfjpCOkxX74/6MuwhgtPxHxa+wctl7V+j8ZjOdnmzyP+wnx
I8JhTsfE5KMktFb7f0e0FdJrpg4MkRVWiDrxQ1OMgyoafhWqopjpQyMj7oOons9bYFziqzJNFZyb
7yAvqFbwR9ZAVNZoG1FHn2ax6oOMI2vD7EG2l2rOU6TIE5hHLgWh1r5VRYrvfdE9GHp4eMjRB+XV
SOe1fgIwNwITKQBan5bPi2IqHZt11Latr+Ji2gp2Fn0yMVFK7gG5/6W90cW1gyLjNlQalVX7yV5A
C+0ciP0+OLUtiSXqpFiynkXuvMtztyyQHzafOIfehg8sFSfDpHpsg05bR5jsXmTs8yrtmbUYELa6
pn4ExQQVWA22H/zY76Yj9mZ8zhmE0NhQc4F9xVLKSigRfzu6MNbDN+s9c3B4NS2KF321HKFb9Nhr
fjOiyvmAT/2JDsPcWeA2ajesBLHR74F9qMHt9j+O4EyViY/Il3569w7CU1Iu/i1QQsI1tlolTwUK
dmZq6J3Jr+J3OwSYVu9TMua2ZMffB7kbBdeRtveq0878j6SRrz5IV3SkvoHcp8rVUscF+0VpLE5G
CvkEStUD1bfM6utXSL5h+tos/dIX63ZlB5544SYrsCZmRtmmuW75ml2tTQeBPcL/i2dP25whk0Ik
MwB9x/j1ZtIub7PGgSohs9p5T79Y1BoFLNSe+GHhQrdNScR8bd0hDXOViF3zCaKTetvy3aqi9G7n
66JZ6SJvMNofKRuTQJ6wTyqBdXofdbeTN5aFDK1sEw8Td/bAFk+WDx+85AIqWijYtmgbptEiNZeu
RJ4MZJAZBwXREVzJp3a3WmM3WFMyu6k5wYWBn8m6JL2xHs3VQJGr8+jH/aG7AIhqexMi+SFM3QKO
vjdfyZToZSUnjRLzaEfPlI53mlPPJ51AHMi4VeljDSpuq2pEYMrKudY5fxOgJ+yP0ZCoDBmy1ryj
usQ6KFAJCR7kynVEdRM3i5hdVaJPcsUMsKTIWBoTb6ThYUvgi7nTrj1dK/wQF/pUssBZeGbOsDXE
CHiySTCMKwdWHSqyY71tyLTU7BKkYY8z5H7LLSGADdYcYm9ul9gd+bXtOQSBLc1sqCYXsBLaDgkM
UcZVg0/5H4MGOXXTy2/lrnOLOJ/wmgoRPqA8zJdfWjpfTT5+kRqklM9RirRcFFR+/Ha3L8ip0wCY
6Kx2WmI6hErVJPMmvYGodDf0RG7cNSfsLWUGxZawS4vpns8Pmp8qaw+EjylCCUJf+j7/UK6mPaxQ
siCvfusL8WnVuzg8S67IeoA9mkIVKPc6hNz6x4v/nEttzTFfweQZrc65dR3JpiavSSBUZRavB+7O
o9n221Bfi3IPt6Y9/FG3jCOmsIpbwBAk9L12d5tg7Bfjm9PYr537mo1+oHbgUUwNMNSrZRLPloaH
K+OOfANEgaFZbOcli+8Q2D4ewjRROKl32Oe/1tUsLWgeHhmZxmKgInvnDmiO/hH3pAFuh6/4ADhY
+llF0TIOMPDyn1ezByZUZtYFT7whNHaP2eLqFuscCEmPfr9mrvHPBZQTVZrDVO/CskUsTYgqHZB9
6+ls2RKWqgXVnMZZ7vlIFmBR/9Y/ivcdtbRmw6FEX73nN8122A+Els0dffB1JZ4ClnOdWg0C4x0z
CLfHNIdqG25zxfTQP4ebJfkDJEYes5ujh/60fxBFWqrPky9gzVE0TkZAZaDD8uEvqdzxzaN5gstW
I7eynwuyywdNeDiMAMTfUrrDqB2c+1DTMkwJzU+T9phOkMOX374YRZSvhu9W90fOEpmi3Hamxej2
mbSRxWnso5RBdOr9tgSwhqZz7dY4kfm3JdHPX4Iz0zx8JqQ0awXV1Uns+bOPtquw/pvgcq2m9Tb/
3JO+Mhkekj33vTQmCvo0dtXw1FnV2cZgTrCXUqJg2/kmPmoBu+CwuO8Cd2rAQ6XaWeY8eQnaKrij
bHu5Jfc+EmKQQaRFunmX/rdMmfYzzOyh1SlaWCxcnygar1XGb0eh+zBOP7zu7w0MTlIdGxEY2gC3
yL2Qn0qqp3vIJEkRi9kFzvTbqUrT0jJl1nKxSCpx5HwgI+wjojckH0i7IHQKsHKNCy4/pdYwdCtH
HglK2Sy7V14azr7WYF7ETo4YJkUwyBFtOXA5FW8VqP7nHZcGis1QD+yIL6sgtwIv15/m8iCDy3Jx
PZLpfQitU3KfafIAjJA+dES1+PNKICyj1UzhI9SBMvBylUPggaTkLRGWQjNAPw5cAH1Pznb+vxrk
OKRYLc5dEFk33lGGgPKgpo675uB41ijzmXuYFuSoF4ojNrEb/3Kbl5ktFfWuWf89UwS9ijvkuBQZ
U8KL3QxMegv2QDHvlZneMqMaxxJ2rDAYpJ8rTvzbD0x46Oa0omlq6ZaFKGtxHjwSX7lLg24SbzVB
u9FZ7c26R24qlaGdvFBm1dazgdqRb1CTz+ZbN0SvrsWUagV/vs+b5KFJfaMoEbFVNt4jAQlmWhFP
uC4R0a2EGbw/kIAG7tJqwaf5TPAXjAc/X05zVJlhlXukLckxpHtznQoWyYFzaXA259GpxcYHzyNe
jl19oqupymoc7hGZOUWyE0h75Jl/Ls6m6RkSXGYSikWsbxmSMT8v4747nIhgH07WmdyztW//VpCz
BXoN12Ho4kvDvb0BhT6BFkpdaWpKAxIxv7C/Z38b8qZdos4eG5kahkLiznRt7UeX4NoMY8f4cwf6
rNa9jdHYEYBYJ8JsjpHdaioMihb+Jyy288Ke0FdtiB0K2XYNyfLD/VZ5/dRKlhLhicwZfgM/qewc
mUFK7wBedult/VMezLbZDk/1N/Grtd76ola+Uo0CE32Zy6oevil8d9WqbI6Maiw9g2oSTQgdddER
VtNErQfINREyIi34ZP501GIfr8dTu4HYv1RYzPgKJCUXfDHHtshR5XNAJOJR5pkJDNPGjpvEc4wC
5aCAW0kY3x3ijw7Tff6S+UjCHd4gkNsBrdKGvRj6ih+6/Ek33ntFK9oGUcYkeCfdsvKk5uCCgzZo
3fPa+UT7ZvpPqH24NTVClT7KqyS9gy7EtlF9drFwswwCKbiXeLPpW2s3rpw1uV1kRxsZcw9mV5XP
VYISc1BZ0QU69Qw4jOF5wU5gRzy5KZ/d0uEwQhaWhxFYdZqbkFA4Xys2Blf3kEp6IsCcOSn0D93W
zzIy7sdD8v3YmqN9dRzaiNBR5j1Fbioyz8NKFtwURY4sugq9P/xjk5vl/fX0jEL+RrpuUtFWmgAS
dTM04JuZLbo7j91q7S5AsA0JMak99UxbUYF247yIFCkV3ebAsCQAj5F0jjhUfQfOVq7pUt7BD8YV
UrZon4vlBvXdy6FeSyCT7pBmDHGIf1y3uG50pZNNCLAVFNpBFvXz4DVNQ19ZMOI0P4bCzMCmJlmm
z/raZiw60/8tsB3eTt8Kqw9pffB1oVCQggleBVosQMWT4kTsaHh9DzNMH/rLKqcvCGWingyeijc4
VLU7mIWcAGcnIr5Kc5LNFvJyvDcTCqpe7BsrTSkvlo0zwOsg/WH1MBNn6+8qqYl/r8YJvk2F8jcm
NyyuRsSdiezJ6YPUg5ROx1Trl6BPkugFWsw70zULpEqWoOI7ctvUJNT81PuZZPAoy1JYWQpGZFVF
JNaoNDQVyrYIU0H9wJAhw25AMsDhbGrJzZotDSxddbKOcjc/3f4LhKfXVI2w020R8gUs74fsNyXs
YT1HsKs/xFnf3gu6vuYOOp2eqf8SBcOmmByJu7MD8KEAIX/oS3/vqEDyjMWQymajCwjTMGjV+zW9
2alcvmEeGW27KUoScAgWsYjlsKV2VCOdH/kqNDm5bqz2YFMoCmM0NQ1NG1ETq/6M6rITNamJDMt2
zqi4ODUHWXYm0IOmK3RhQwNyAZaDJmK14fY/3WtJC+gwuJ9Xw0foGL4Z0KDbasFeK/y+xUlUv8Ee
nG0bGeHO7SP6N14lWWBMVbd/2XL5SNc+X4L/kc6AN+y2SqSet3gfQVri2wMNrpDC0NUOXmxA8KW8
D0kdOk/OE22CmjCIuZRREsyrMRY0GfGARIB76lkbOXUAAqi05UypTEaQNeiFU/OfZ7t2kwCHJ0df
HnSueqWopMjkgFkWW4RWJoQRjwF3zAeBgvYY6IR1iVxs+haJdBWnaIP3JIrh94uBp58pi0TaB6A6
5hT4Zk0WSr2vxj2aqd0rDzDL4w4zyiQce8ZcHmTR/Z7qV51oEcUxOvMVmcBwwr+bC9EeRMkO9/+v
VwgTJw1uzidImyxJJF+7li85uenoG0JCgXrLKoRUjyILOPZenA4LLqi32qPB+S1u0NxkJRPU4YhX
j/qofgIqXVj46xPkGqGT6Qbp6AB/qFPgny+r1vyfLgxkHIg48kOu6RvdvXV+7pgtIYz/ZwJLMhyH
qFE4l4RSVIAkCEGEA8H3CqfV3DvmdXDgWOdNhBz98Pym4cbDrWUWpMl6rSB55cO3jihqUAAEBzU5
MNiy60WPnzfDqTuNY9yDBXyMzUiSa3XW0dfJ9hMzSG/4cYJY6v6H1apEhMOkSOKs5SXGDnBfijto
M8dvKKYzokYaV9xn+hr0rQr7720+rgHK2mssxIdjI6F4Pb4PnUmRGBahoWdCB3HYnXCaZ0LVGXXv
kg8US4/OQ2U6Wgahb8PabsxX4r3cW53K/Gjwx1g4v4neYM5fQpQH6GiGtsyvKWcjNU4al7PRgNOr
usvCpVjoqTLoGWl5cdF/xsRFZVfawV9fq6/LBAWbwtKMORD1ZCVJqio1dyVehxuf9cd7TUgsWo1f
UdlzCZyJN4lr8d2vKKFrU9hYJwwjOZSpZabTfuZsV5yuZvqeun3hfadw+T9E3dEo1BvjGOutA0x8
xmAzJGNaqDwOMssLUc2ARb4BTBefIwmkIjrCMbDCpcDTF0Q4L9dHKJ5b9kaRsj2cRpDBF1PoCBQy
e9r/lKQMfWXhjb18fpMx9cbg4tkB/69AFdS1OOxnUEBwtxFJVWk7inVJHlS8HEdRUZ7cxHOUkPzG
/zaTXHJB6TgMpqB/pi/lTT6KtON1Q43GqysahNUCrdyXCNMgAiGrTp3fpEs96dK+8UdqnteDwmPh
4eGgu901XOq1AmN17H7XlmwEcmC8di8ciEmE9hPn4XCEDUwHVkDkbuHihkTV9CQegY9hELrYOjc3
bW40AdKNmpj8DOXOTtnkLpKyNm3ZS7UBxN5S12MoPHn6I3p8+s11T/T7oQK1Addm/jZaGqJr3AqB
m6dX2m1d9Dk1Kd0lsBwn3An19HNJPjgfZYfel5NcQ+voBEzJayM7z6Pnp06zJHUgi3TKspbTHMtm
gehEvsGboUp3SuY3zgas7p5CtEX/fX5DycdbjcVYgc/ToNWRFa/yti0W7mZaW7aS4r/txySV77QV
GtVtwjGfAQbCNfJZLMiyWSJWB8oIlkoX97VNMKiiAEOyZKu1ETHwetIXI85WweGy7TVQQ7LmxlGh
Zhu+Yntm+ZBol1S6aDya4EMNAX62ORIq6qgdD6aOfpqBOCF0+wpFjzlDrbfLJis2wmA22LvWgktN
YOEY1CHL/V0Kv9BLadOJZwgQongY4dLy7yUopFZlgeTZ8H87xXy8eSAB/p+xCPXCFZIUgPJjAc4K
FUNo2Sf6wSnGm6VZzaVjbYh9XdonB2pfurLLhVnQDZqzca4+5+ZkVGpnvWKmySzYU7XTxY4le4jB
TJyQ69JpFiekJuY7LVctowThHDQws8juhUSk4Yl5vkILr5Z3lJdDYu99i60QTyP9i0X02ikYhbR/
ygtRXn6DtbcSIVyRP7Ijo2wWdIX+dpyamXrGX9P84F+aovan9UALXjMRdcd2dnJDJKI0ttXlEle9
yGik56excKtPEDKxkFh1t4tt3c9bHQWmMtmvD+qS4bKXl+BQjNxy8jpvF06JAtorp/JEgDXT2yGv
wxExeQ4M0lJfKUw9o2wFDSXJ6Efwu5Y5jMKmOz6TpeDz4mp/sD+EwLJJtGn4pKav1YGzpVj3FTeY
sUx1gQZa0xBovR/CKQhXnwHO00bqU53UfSgf9OWoAfmd0l4bx/nFZpRg3CgiQNok3shAkv682Tv9
sKnmXMS6FgTFSloaZQIGgIr4U2qG6vX3M1D/SAYIkVbFU3V0ezV5p8htyTJw+ccym9MG9TYi4Sqm
qMHWrSAWFpWgsNiyfUFs6RLkFwmP9v4pV9SaUA60wbKv9dj1xCrFer5hXhTaFmzvGRXDggBZdWve
udxi50iuEJVAjIorEf0CaeTlXhmufrr7YxSBsDvlFxNitM4r765+jk3+e48CY+waKIrL+hm2dXCp
30nvjjIaIQGpnUKl6rnuYZVlV0l33wJQqGb+YHvllezBB/Gy4Ryqp3KVo7ltjyZrvf4zBQ5+O2g8
fcjKUyIzznY5WLaVdevGdIR8poaDF+CHXu2TzcWPAWV0Ee3ZPDmCwkjG0aY1vCdQ6slEt9oJTmqe
I1O25Y8S25Zy2U4/WCcXdAdlZtVLPrO6zlZBJizzhZPyMh4YZdUy0hc1tzqU0W7aHypcE2oy3J3J
zwRqLk+BqOi+ZYAJgoTqJWj8hNFDQFUnpScvg52+BnvSxV1hVkZ5C3m0U1AUvsDAVFTP7S2BvYVZ
0SPOupfK+fwt/WgEB84ia2UbJGm1lerV+i70bE42LWPdEgiQhdXxlA0gq5Kp1dgMn2eET5g6BKKt
z1/h6qCRT55w1be4MWBohWdW4cYECvTdzTEgrN6M0CYFn/MTTie3sHCWeOCQBYvg7wHILrpqs+By
tQZ4OEF2NKmB8ot60flHoqGeD5pU5MhhH1PcCuL2VvE5Ghh2O9MLAGbQ5rRzFHiutxN4aUC0hSAI
5NCO7C962JcDQ+DYYDR79ir1GCnPhMEWYhdFLkhpU9kYWc9w4u8u6PNoXmvx7yWjt5JDAZNyPhUI
JFqR3rsRSut10OBvoHbQfakjZkcROEIT+xd/LXvL9YpNAtH+nhLf5fX72mvWHEVzN3WWtUfRVdy1
lk94umithBpdBKreOW1RWtOWW1omPHlg5KA8FycFTzRnyh5lCJu2U6daLSrkfXa7Ykk0zN7TulWf
bq7q/9Pmu7a84rBf0+DH8eUc/fMJuNs32zPb5UT2wwSAxNl+a0ulFenJEnzquYNKj914Eb9KS/u9
pbkX2SHCXi7NiUhY9QmmFknWk7c6Se+2yEoWFpZ8IjprYmnXodpT5yxTzpoBuX4FYfeQmTxnTKTU
RpQCEcL1FEaUQsKF2NAlv4lAlPYwhnV5GNLAfNsjx/IjhDhxaNROHFjughYfhZ9SxU1O8hLgrzXx
5/PShfO2DVnN6b5iWHy04/8px1mb8K/aGiu0ccHc/kS8v3dzi07lOYgOnFDGlDcaF54ehbQpE4/o
ygWpWV+rdILw7kuA0DIh/ZjQFrypZtVY6PD6A6/iaoZDbI1PO+NXd0oH/UyFNgW/VhGDuvs6Kt5r
PidRbqR8FirRHfpKwAGxA4MCJdi9jOrSyjwP4zyP1nJzRYP5o7D0EfICYIWA21lkpDt+HnsrY6kB
8i6z4M42Ntbz/ppueTWZy4itTJk3d/LpgVRBpf+wi87CzQFXBUH/wM1Ha3e6EUqrBojAugwLRt1D
VCt+PpD4TtG0f+d5jUPzx4TtHHFgYN9Bk4rxU+BgMB8I6kd9jKyCekNvvt105LVqShPq5gjea98N
KX+IgLiuJFj/te1gztS97Klm9JeduhTAD04BTLXdyIBJKuyuB/8c/BURGpXDZsP9ocnQwg0oCP3E
hybSLYruQBnld0yBrGaYPIgaFOC0ALf/odAF38ten1DByFLZW2J3885+mtGf+F3DdizAj1MeEikT
eF+N4YZq6nky+stP2txjJ1Ai7JpCz3k+kt0qHpD/L4nNKIeGZD6qzohNGTiHIKPw+GXX3TWWgDKe
LrNsXJH8xo8AaJPSI4NzeBIyTq3Y2+3Oxy3rCN7XR77gselS53tufGd5vdU6AcsNPsgSuz0ShGxk
H3no0C7G5NqxBNAKWnaS+KOlVLQvcvcKO5Y+qEq3zDCU9lmCG6IRBXJ7fY7QeLNiP4na7FUPGx4j
iIRISwxJkHJmjEg+6rlhtFmHVFzFMaTjSg0/yH7+KK9U84FxzcPq6RL6s+i1l7NbVpI/o5Q5aqI/
iIBNJRnU/TdUooMlAFK3D638iD6j6tR8Pomt4qFYdNCqx/O6Kle7l9rQooYeoSdAGI3xZ9htTiVB
fJfGJVjRiC9wxb/At5hivbi7lSjeFJtOQg+KHP5M1x/t6h5QapOavg9JJvNe8/vPHXvymNaQ3WwY
THKnMIbFMCc8zUJj4NL+0i6auSrln/fxqQhlRgMkwvVtRQ/HqGcmYFufqGCDRWNqYxUUHj6LmW7N
NKprk8w82mt/RDJj4A4xPDUokTFlLWtHhsIs/onvaGdRw1VV3loq3ioLGqVKcwSxarBcKG/w2Qtk
u3DZGnXOiAW/gUDigWz/64xuWFTMaJ8Mz42xDGOfbVsHjvhCo4u4KrILL2D149Xikhch+bidzUkL
W+w7qfNCCONDIS3tnZgMDWlSkCmnDJqbzEFCtvg8dUJfxleC2tg49XiqUauz60juzQAmmk2clpru
uBgkb339BUOgJwtj30tfKTP3KWwi+SaGolEwLtPkkZG6ox1ERRvEyOy6NPM8yZ5C9262RZl056iO
ciaErWEPbt5VrPpRxlUowKXizXsBHV/HwMwH68w1upj35WshZepWcM+M8ViF0OQmMMKbI0CKrFr4
RnuUVnxQ49N/dOMm77Q73VJWea4LdICxubOMdPQ2XcRW7yfxsIgR+GEksrsGispKLXcp0eOiVAOs
KiMZTj2NRN4SqB2ioe6bp1o7mEC3OodmsxFQ8ZZpqU4LBW7P7Vzf37jryGw2qUtfuzpystVNsAKQ
f228QBalHtTZiaDvoXaI9oVSwJlOQ5rEAUyTmoHJcq07x7JXCZo9CLa+8ryo0UP+Fd+q79ntjzpM
p10NgvaSwMqnnvqcUWLPnpT2ts0TDqKw1qT25fx0GImHVE9AMaw228wiM5kXTtNNmG/ESWZJ/SR0
9hoizK91dzSZ2XET76Cr2NPppwVLkX9vyOgTCu1cH3G/3I4RGbjD79Xhong+DPDZAOWiGjg6Mx08
TTnUnF5eLIJxbAuf1lH4qy0feUUz7zZJyc2+Gp97/flt7zlfa/bC2yN6yiuQXjQ2dsDes54LeOmd
fXdteJPkl9QiPQk8qx2JejmBh102lsigH618VUtya/ALJVo4WjCKBOYcOLxYrDW3f013+iVJx+xj
aOjuVHBSeaT2f9ZtY1lNGgoW/HYp+ek7716iKg07VZizqEDmVfaB6Y2RBU0MG+FY7QpTNrITwL8s
FfQvXJuRtzszLXd9J9WC61gwtrJd11WofH5WgsjD6TOMpgF9liHDP/8H5gDY/jt3DE2FQ/7kOimn
m1ykIA12XM4GcfUy/gkz2Anb3uL7vqtyiZ0peO17M9V0hPY/RnyK1kwjDXjDj7a2Q7FGO9njTBwg
78eognAfbky7fmNXTEx2B6vI9bKFrq9cZjxKGB/PduThBGVUTET1QXbtlQoPldww2hNW0kvt2Nz3
9hYuFzD3Q4Zo5reZ5en2y63wmeY8lBtkE6aQWw1zKL2G5sDpr4rAyqcR2bKTUgcbqq8UtdG3JETX
YOANkSOqQ42lh2f5l94hbArqCxvA09E2nK/WJYSHIctTkQGMqpZrVZyCzsqJiA4Sv1OT4sH8EdZT
AbNKPYnr/7nAeNDMn8AqukcCG/pGbNkXFTjH4eZw9SkoEeGO39uHR8vBKkn06XWMb87hbRUfRYGu
emdI3zWNbGGLPtvrUkQj6CN5ZIL//vojNMxINI9jwHAMiYU48KrulY3zeBzBFra2G1EzKtZcKjCN
0bZz7MDhzxMeh2FpuWSkVuNvpGIl7l75jiUfjn3g1aS3DFpN9L+e99jiorg6ednOAU6TE7ETAilm
tKBlOy/eWX1AwydKHsdJfkLbV0t4G7pDNpZh8ZuYFbFibpo7+M2aUVsYx58qsv/GJjCy0iyLUq1o
wwS0UoJpcwCL7ptCfXUI1ufPbKwbTRU2lj43m3wpDgLbPo9b5xNsiwYHHD5/tiYXgcnvtjvTeZII
QmCCyIhMdAfHBNpp1P9bL3dBnhDEcmSlohRro+vt7pVpDLfzhsS7PtgSyNQbESBxxHuKv9N7lQ4Q
B1G5pGsfkkqQpg6DORyr1Y4LYyQ63ZNQwm+0V1Fw58Mipyj8mt/c8xGF35wGIObpxUetOy4bYXyS
S35hmUSzUz/vJzoGz2YSM5aa2hM6IuWoZPYqIdRnAVUubK9R4VlMqYkKdVN7ab2tQzkv6BUVX7ei
vydNHl9NZiF8YTc6Vh+Y+JXWiYq7AU+rhgP6r2UemShC8N1XHSisnOVYs+hd2q2sKLdNkhpb5yzE
3vIqrMtqtW7mkipG7dp3t5iVOXyXfAKQ5KB7Jlpa+kbf5DXEKGgfiByue1C+RgjesULePRHEZBHd
ol6hbPX1EjuTR5MFDbc4PXPpq49qmR9iMvITHLEgo2jEArQi9rHs/+3EYUfYMdqvEyIfBDXwAEZJ
y7sZglMUmKzx/rF0t2UI8Emjzoi24nCD8dqiB777vwkacI0d58VzOO4T4cy9P7GBekLMJxSMhzLb
cF/nzxPrmtKCiG4GW8h1VSALNXXiN0RvFooyo8aEgvtvVn8LLBWbPvVsIM76KMDNyJhfaCdNCWvi
DxcTEZdlVTjj3R0GAjga1ZPwa/hbeV0x4+fMAvln9QReDiLCrOjIGYGM+2VhIKvDnJC/DPJl4Cm1
JrOvHvwKEUz4MiSEfiVOgxAuX28fQfwdYoEmsFWqyoPjKgV02vYpkiRFUNN4rAP6srWKpt5Packm
NbAJZAQMoZYGzGhJPc3waCdEEXqrL7Cj2tdPN2zQVDrLRbVCrUqwHZzLTLLrol0f6bNO8k9NH5Fw
4XqP0+7cbAWsr1nkLKDCHw0xLZvhkArZhLqBUMDtY+E6473uzH0DXVJh9JMe0NKakfgG5OojNSdT
V+qgwqvGaqnnW9KkR6+gBdGtqYDiphcmOUPGtZaaUMoHigKzmpIOmKDfpDTJfykXixp9rd+Di7DU
20UpWYNyvxJBUfySc+e/zueck+cGsQM5o1zxVBtWLm5m9fSkG6fvKAqW8ICZnZ/UDcU+JcUf0Q7K
gjDCykpOP8eSboGur7F3SeboVh5lh1GcN/BES3tBX/A3H3hZ+mwvcNScwb8w525uSlic2T0cB515
RckTNJm00aa5RD+/ozGEvIwq1yE1VaIMOvfSbqbwxpY9DyyTfd/rM7007EgQTzONXePlwfhvK15a
+/w2RNKLcFlg7eZ4mChzkyPM3WzMbVDNyvSehsrl3YelzLnlvnssREJNhN62JCPiw9eTe0/coB0K
jG9Uigblp1b8IzEkcC0K7UDiOrlwhYTfiV4w9J4EojoAv8OmjPqMeUAG0PoUMV2l0niODrO+Uk+E
YrwCTg0OFCSlP7AbmV3QQGkAoJl8ihC9Hv9nn482hmOgbCf2XVyG7bXMO+RHVwNeFjQgR+025EmG
GbtqP5icKbb3Vjd4jy0qMPARYqEKdnY5GnunqdPtamHO8nL8SfBBdOOuGmrKEShgLm1Jgw6wz18z
E5SmAcSCDEmqwcdehCI/U2XesmLgVClN9+zwiCInDO0x6IIh1beK9UBbsIp+voLDoSEm+Rf21dAI
8LeJg3IYLxP/LNRInvuO7mnAjyfJqBOQoWlZF8Vh4uqYrTBUnAph/oAKj9pRiaTccqqT8blW035X
I5G20RrIApxiGV6djsEbV49bRpDDOnX+v0Vl5YyzOhYz6c1dnzTs4Bgc2PXxkjILkmZy5eYg3YKJ
0kaXntEUv9bkojmy4eBtVs2HBpNLfS6gZ5nt4gFqi7OBZNN8+r5Lxz9uv3XJddeZWDMWtSRxifAM
QBPP13AmKVc96ERG9ZOE7nQOmdc4NtTi6+A5iaIIhDXa2VXAemE3RrAyBN41ZuP+3mshyrsezwiz
NX23Hga6PK/v0p74TIk8rLbDa9DghViHmuc5UqlYsQIMcGViMNfUu38321RVoL8vX/UK0c5xzot4
dZc8iQ04eFlhhFnShep8GPEW5I8dkPtxWPrN6avy7qJh2XCuyPo+hTGHk4dxy2NyWPAuEwIlY0Ib
oduRYjYtoHdN0ZGaxLPHJTZT+r0hFnImYZYdxZCHuv/V/oZOgY6d+SFQVRgD6+v045VJoaUa0+wV
K9XFCObODKl4lleSEEredgM+Cv11UFgUAvfYgsjp2Lyn5tqc+6i7eLzmXP01rOdunOjyWevvgCUt
+e22i+BAdfKGWX6dDJr0MkeMQzBmdzgfAauf8YWJ7gMMjKCrwsE6rkdXw3UXzXxqLPhKvZ9P3U4Q
/JZTG1IB4UI8Ox7aiQ6RwUa5tjfbXNi+r6VufYAA4BtC1y6fQNW1ogeZqqbXtgdIodAeXy00xmWy
aNqmAn++1XudwDpM+u3LI1sSaRp/Ra6QgHvmAoFA3zu04OQ40DXGRRkawTi3Tmxeio+ZgLYV6JdH
OolRWtVrERskbLGeM3Qk4LNcQTmQ9KuOA/kdm0tu33Ey9CVUhj8Sml2mzdaVpRYL/8T8GrlpIwoi
pBkLIid09dCEUlc0Xpz3YJ5TM45scJZi4gA9qP1W2QHYmq1aYXam1fdpPRxdwdzvUhb4JBa48ypz
yijPxKZvOAcr1oXaCEjxf3OjnnJNe0ZTEINJWbpbhq6cyyjUjQwjkXGRYEJVSo8cfmYwpBnzcqcD
xfYDPfNyeTNpeVyOVGj2vHvoftf43VZuEavMuNevWa4+A6Pf81fpKCtVPLvk+JjSTaS6ULZADSMU
ebbc/UxWIm1yxqWrR2JGcEmBWLikcx/H1H49qPl89Sf1Kq0VwfQ5wH0LpVVM9qYUrX/9iKpWF+dP
SCxxVhoTy9My2ubb4aDrWrUBHyfOwg10hm+pyV7kAc8hao0YcAGUFZsb7iOQBk1mbiw1DZAtO0Ou
g2SNrq1wWHsWwjBVZuxAcC11u7vl0EwQ2bObCBxzNdOGGySFcTYQHvMvValZghNH4+m+wSXpyFKv
G2OlIjgooxIZTEOFkQCNIqI1uc2CZIUmuxx1NNu9GrOCvhSHP1uWj/RHQaFBVawDLB5yt3rG3+Vy
zCXN43jO4QBVY4jpYVeacMMhGls3Ph6iUJKhe5nnfQ2SoWxEWZr2Me5LYJFomim8VzI2q2wGXMxk
2yHKJvEaFMA9SrtQLIy22N2HDsUYdx9O6G7EpRPBDmlWVqU1+v5xNyJOozmzBJLoch3E6zSVle2m
N3swll/o8VnyaZebt+wnfesmuqa1O8p2Kq+8A1v+OmjLvm+z0c0KPgem9Hedy9HS7CM56mwKBJbp
ij+0n9JpqneYajrZXzdXj1tSGC4GvsOFVi3HTMNxk4tKo9QlS/GEPOqZTdCw+S+ZDurMeWTXEHKd
RJAYLWrmCdpNoqc2Toi9Fib9EibPQdNEQ1z/KhUOG8X8wNenzFFjG1sFX7f3Qc6p87VyxxSaSiB/
MCsQ4LaFefYlmmXPY6RX7h+z1X1DWlTOjJlbqc1tHvh2pJLh9W4qXOBctlroZK7HGcgbhBOSbRY/
Xd99dc+/eP00AiSbeSRzWusQO2Pm++N7v5BohznoZU6JO8ImbRF6ry04Zb1OCFLdkH4TY4QtreL+
hYME+zjOX0eJSMbKz7qhSShrTiHrTyXCixhTL5HLeFqFT3Q7las8zHZVASRROLPQZ6ugdGB0IMQx
3HmzABSh8lxa00eJB/Yhptnpa6DPH9OvHJHFZzOWJplgE8BuBOTGaPOOaqysNpODbWf+mQhImOEi
knyq50Oew2VCZz7Y8vr/4EgVzULeNSyyIOdGM4anYZHIJdKz+LpueU4GBEw26wOMuezR1gVDX2w0
3ZEsjM1dBohr7BlXvBFzEe7lZw4vrPajCS9LoVQ+ZvaeHZdzie3hHlu4/X8ZLIxEyAsSSffAxtTL
m1KRcSBKC1DH5d0h1An0PWfJ3xFxHUXFrIeG4oAh+3xHttW+bDw+7Sujz0xM6czGGlCx4bAL5O7C
JzpWxBZF1qi6quY+qkYGJ/PQAyLoZbdLAcRH1P5AR5HnBPmyA8lSeJLS/aa69fR002M9zHPJ7e+4
oR7s4diGy5QFaoxiVFJgb3VnMpKtl2VMVT6OCJq5hPcBpbj1z4FHSJmX5Tf2HxvsHe2kLQaPWPWe
/Ifg6eT3Q8aWOtyezp/c1GlFu11YhBWLKe2rFlhTlaruyfj82N+INvCMGgmusRrDM64hJ/hlP/jX
6zO786Esj0AWXf9UCRjc5PlS2VKmdQcHP9Ys7VbS47UlRiBTfpvcSwXf3ruLSiUFFuUMuc6EtQY7
dxMZClLq/6ijp45qFOZTg3ju1Y9xNkuzuA+5Hg5VQKHzYbnRYqBfweY1Xr7CAL+eiOVshkRN8m9C
yfddj4ZFsVDvTWkbb20j5Zc5dphmSHuXQIW38eyCwvgaY+1/BxsAaIdkrrz+QI0t/eOKHQHv2MwM
Z5YAKggUzWD1wHfokgutioMQT8sJjiRM2Mi1u1o/Yyj6c0PgsdrlOB4AfH3h6pQT1ank7JZn5BZK
AEHklEgIJa1rolAsLH1gM9yRCxPBe5qL7kpQqjju3xwGYUAfwF9IlpgjF5XHzuqoeeJrfT+Vcyl5
j/iWZ79eHTcc9G1iHJPMucXrrVBgm0gxrppOcUppbhd+lfQj+qIm+Ul06tUkRmn9a2kAA8KP9+yS
zjnlv6PvQVnsxTslLSCR5oTrRW6CwGPCoF002PKDqkX9ASpGBgk5cSyAz7XRTtGsiqyr/RMRXphj
zctbr9K3hiPOYxRsQ4aDAKzIjwZM5zUnyZZ2UVRLXDX0ZAxSUxGkClvpZkMy3SyAZ+KrozpuZ3gM
0XPI7CgO0EbIPaTwmchCW/SvZBXqshz6B/QO/1yCxx0y2+l8QNS8p8pmFj4Xz2abNfFioH8EcZ1l
Jmvsp3dLFPpPmfuLv6T9Uq3vFbXmO3Rv5kDLOvBi3Xiy2E43zkSH28xDPg6uiuYMoKAUyv8eQE2R
KAa8zzBymFlMzaaiZWCI7JJdK7EMhQjlMJ/jZPJa8+YaXscD0KF4lxM93/76i1uCj7z9a6RxkKC5
rAXsuFvzEsmGDXvHQPZxtMKRCTlm0t+CiRE2bClYsxPu4LtfTQu6Y+o88fTxt2zlomPR2k/KWke5
MbIvfLXwQTnOJYiovY88fDuOh/UtpPGcjHmN6E8GP0dG8Og5J7G5Awq4NnH55n5OQy2Uz6nFa7Ye
dfKQKyX2NcS3KIP6dFg7/AA+tNjdLaV0DIH5TuDXNkLMcDpspyanNA5pFOYJgaBzbydwQpSbZ+Po
wTZi64/OqOWjVr0d5BGNJwZYt2W6FlbQVxqXsOlcPf0QxCpVLStXc6xXXZerQ7AnqX2O8xA4gSxL
aqsqhZzHm7j6umz5XXzhQ4euwF2B9X3FJmsO33iJuQJsNmgXdWTF25BdWmb6jJjfv1yHcHuBMlLY
hrL0AiuHRsACQvabsrau92SEc8Z0m4fNt6hSgzbRUO+Hh3YG1wvtRyp21bKMfISGRBMrrlFE6vB2
3M6l6ccJBsigZZys1w4usbT3IApJxC1yU2VayhMxrUcEuP9+DqX89txLVje3iHkdjRHPw7akk0cz
mRPaSMaQNUg6LlHB8WMmcnKT/0CUmHAAPTZYfZBzYtnE/RNFGA0nTXN260WvdRS99C2k3If7bFUu
wZRrC4pQSsZkqhcC1DIwxOm9dzpi5IROxvakzttwZZ7uLo34+so1xVjbRv3HbHLwzgYyzuqzawml
EJpz8LHqRS1NZ2QGdvexrHao7nKIW3K0ZAGjjV+3JABCcmgQN/1Dc06MPiYVyyFl7aLcuMxHLDQf
bnwkcs06GEQ7KshV3CeDMwI3NQU6aIs4cXjYXxKeQ4sy7oGX3c2ZxrLiwsmjioZuM3Ob1XQ2zHz7
qMAq7RdA5ldhSjZbvhaaE7VZU7ZGjkizO0S+XfIjqjKwcDBnAp01yaAQjS0lmC7+BsO24mTpGQal
XXVAqSYWZ6oHYdRA25mN9pcix//VZ/v0sbCjgERCwJ7oAQw9spf8xC50hePLIfUkBdt/NDOEiHk/
mk3lbsl9qXrA5n6gk4oHTj1+3cUFIIxS7MzvSQFYIBhGP+ykagxXzGgKWKWmIyATobPFGklgmOHC
6A5Cx7wK/fuHxZz+CCDK0YjQDV3nR3aj5vCarvEZ22KZb+7XWGcAQ+A8VypRbu8U5FOwePcKiWE5
CsSwi+BBaY8G6z8DbUOnQCewa+CQu1+6TpAaNAZKXntThoD6/vnblSyHnVu9qnCs/+Ww2ysNMf5N
WkgjHw5h7tkXRi9YlYoecS55Nu9wpojiSNwUv6EUMlA53KsBqGG6um7qCdg5DwjjtWVJoqWLxiLo
K935DfMqQQSYX9mRfaE0u3gwlYtVBInsRkvy5vEzsnICPMWEZ4s7+toCvhy1JjUFe74GzyFoh/Ih
Dfq8BVupbEYFfDJgP+Orw4pqj05UJfZv6obPhIo8JH+rAbUn/BI1HHfaqVB3XiPXUWAMDNU2oyia
Aot9/DQkqXkj0nK7U2c676/IMM/GlEwaATZQppl5BwdHzisBFCmN+RkECyHQqL8xv0BM3ioYaMBa
zx4qdY217vDBGb/pTB+1L/gtDrfvthQ+vmSiXMRPbVx/iQP798HuepxpXWs3Lx+1IU9T0bWwhNsP
eZY+3d/GcozZZJ2D4q2XIygWAtcwBtZCG7hmIXAyRBpB1+wpAkunascAvEluXqRpVeZjTmFZWN76
Cp/W4gRYRF4OfDiWkUhnZOdE7sWxNILfPG88Z/aPpciZTn8IsZT/bXY82WCeNWKDBxOZfM7kpEI6
fvfsW0PyWkQd3WZq/zCTGtdGk380GgIepH30iBjjUSSVPGdlOTj1CTEkDotbZU0yiEy5yvQmXZ7f
Kf/1Si2Ve/y8OO9LYcDfNgVYmwmgeEzeUJcDkkRP9ZD600URUmx8xKu7UOQn02BFwi1n6CvlEzXI
wlYkXi3LwfnfrprMOk5hYIJm7yWV4QJNRTZGQc59ay5COnCaCUU/LFOgZgAXSy+iIjbmujHf6bkr
4L5Wb85FidqkD4hSMkTGQs3jaZiMGHRmYABOq1x/qPd7w7qPUlXcehnEOtTH66tY4YMnT1LVrgG0
szjDMzTJFr4TSJYJZlcMFQb/JmtCAIg6RAraUaKMNtcJ3MKFMZknEwEm9xHs6PuocuZPwns1oTY7
qdlY9UplAqfdiVCPP/m1LLaJO+AnCtzGseJWdlUmKA1Nn7gAvnw+7m2KlQTGLdmlQg+nsZyoEYqY
bZ/foGtggCmYNElkFfYg/FGsbv96NdYSDiTiH6DAuHS8k8EX2EbriQVV1eDEzKAM9A32H4BXsmo/
sTaxUpv4Wi1FGMCB9Lf6zgbicir/Oa7KfrfTa37pcKY7AHMARjDMq74N27hWUh8CzW7MUHiWzKqo
Omml2PbETln/Y9Ya6vAN9LkJVl2CezMnqjIm4VOZCunuU3fmQyEDd7yq5YxqiU/Qk/ijG9X84U34
mkPOl6j/RqN5DwhF7PMFYxiQf+8LuG/S9kzNRXGBUQjPDs9jNhIU0j4bECrQVd5ipMLGYcoPYIcB
5kxey6tr3nBXrFZfT/53d57XYCn0gSRsR+3JFvyvsbCrsIZT7xa5WoJ4F0S6JicikJeC4thMSpQX
EychBIf5K/Q+8DisBvHseDOH0O+wQXXK8/uEMEq7rBgtTKlQcvR7h2Zc9u8lmnmD6Y5PbeZL/xMr
8fr7vzAssMe5Pvy4L0WymMYneXqBSNWkc3KOHzNhkEYBw+GpHgT1g9UiWwOqVjZkQwTY4MGFpP+a
5pdXJGZyFZbpGgfdqOD0HYbI9/vWK9tqV00KKfX2MT+9kcNgR910lbuN9z+FxsNJFz3fgFd7GuNh
LKTfJ9XPWRSPrOr4ZGJwzdu/39wRhDQ8Iyv1C8uzVoUaCAEyzrqM5Ru8cl2bjMMzbZ8hG+GM/Dt5
BXJGE/vLChNFHAk7ZbsK3SADKwIW+0rUm+lkRCGphkvpjva0cq/lMKs56skHAWTc0Vij8VA1cM7t
6j6Q1q0gGiZaiuSC9TwSR7n9dpjikrO9TuVYN0vB2+byWBz9WZdJum+JBii4A8GXcwYhEkAAYnvW
iCey1heRn40zH4tEG8qjOlMl5yxYLCdR1N/XAw74ee1/GwHWyLGmKSXs0ueBQ1LhsjHQT/Z/l2iu
K499xCW+ulRyLRv2YgvrbQ/d2gHM65n+LxXB/g9r8Al5THpx4U8RJXkoclWDTQshIpH3F6Z6csfa
zDqCJie+KpZJpyBNIiU6BcYVdjsZinJipnF3636uS8U+8qbXdoo4oiX5IxfXsoNGFUYQorvXDH/x
F3SJoFt1NaasyW6lfzkiHjFAtqbRxBRFHQYqZdtuBZzN4vsDhk6rhodIQ0/R41YBNtfTWiThhcpa
MoMimw4sTdqXI/wycFwWAhSf13Ng6GccTdexQba35l5SLyNVkbRitQI0afn3Zh4ZBYQULXHgW3dn
BueX/BNzl67YBfbQxKf6uDDNw30umMJjrqdBLu0DnuY0V373PtbOxkLzsMGH0jsLDAYnVTlORyAH
fRPa2Hj2+kzdYX3dYwYDfbKS8qaF38dn9mFcIoOQX9iYq06PmHjQnHv/Z0YFZL9idUkL2qTdEsdY
Et6C/h9XKmxzGr4N/QNv2i/Xt9ZKsMf3dZW1X66GtdzF4D746lCO30mVdeSFBpsHcP/NUDPvGwty
8jsFnMbfhn42yS73/SaXyWHNzNlEdN+HSyon98dCJjZDHlHY9koevFJY6cYKBF/egL0LtKIa3UgN
Isi+u+D6pfPdt+PyBxdPVZf+Pi8YnZ7NUq4VEXf7La2xWNFOKDkhkfzhc2OB989+gL0l8hgou2xz
fr5nczcORyq5fNTVdO5idpjh/vtF3L7mcrSfxRKVTq5f5ZY0jKMiB2ttNZuL7s+u6oGJPcXlA0BD
dA6fYHUJf18iPt3oqPnVwTHhj2VgvkpcR2ZEvaaYRefYdQVzmkIUGrO3Z8ijxs0RXNNFeu4VLbb2
3VfwJsEeSwcVuiQa79iZAMzZQYuD6zdAND3DITfoZo4v1hffzJpFv8SxYIuEs65jTQyX68ajnnxr
vP3KuXz0J4vUHye+Xt2bIJPQfQk2txmGFw/O5m9/ATvWBGti+In4hJ1Vd5qaM4b3bFYYiyCdRDtX
jmYX2aomoqbJe9ka90cdnT4L1l0r+NdTTaMuNfdj1aVC75NQyM1s9B3f7ZMFKyFGGyMcHyYYoDTR
SWmX3cLTEH7wLElT5EJQ+fqHIGG32hs0U6H8EMsfikKMgz+VfZeNwLvwZQLTkYK0jwedw8UKAddD
U2zROZ326/YcQ6WOwuAGIV7oJJ1YFTw73YHN65CH7nNGNe08fI9YQy+u776caT//K1IElRptjs7N
EmYMh2J8sK1n8OY0oa6HTIaOHJ//EV1YrZCaHgTgWsWt1GZIkF+KeroybzWNr/o7bakwRTbBnSTH
5tbUuapodqLNcD/wIMI2ZGzQ/iNpKfMSMC6JyvshWUxnoExeWJnxztHbMUB6BFDtkXw6kQ9YK0dF
MvJTrw0nypc0WranbnGq5xf0zDfiGEg2pdXkm46cpE78mjAhaaHXLt0QV5JAOP9f7kuXpomk9MlO
ZeHWmN7DCDU0I7TQ2a5+NCLPLW9CM92tHwLrUGGftlCtCgMWJj1SWA5dcgDEhToJrZJp7862F2dD
dX5folo/RUU5guVSOesvPq4HxifezGmvARG0RLBl88j9PdRNyfcfyab5BzBZlj3qwp1q/1BDrpJf
rsQhyXjoo7o4LakU+GOFpE12cE7ctnNDfFbCLOFVX2sYRS7Lxdt+qe/o8Trwi2/fU8voBN+Eu87j
8I8HKmc0h4bWvqLxmbAKTUtn51lwgUCn44APj43naa+xe27f/TdWFjkKJwMzamaxq76wEGSzJXA6
2NfFwVzhm9a6jQI2Aqxmm0R5Ms2wDaTEy0cRnLHH8mcF5RWa1/8dQWEzztud1sdaTQZY53lmUnwy
Z4EHVZ8pZWWqoe7dzYIygdEeZzUaHK8zNiGIdSAem5gVekgMtfeycqDspxT4g0QflK03qWF9V/Zc
JVSJR2CiSH9wxMakWouBys8IgHfBFA7r4WOJfLTiVJY/tib5aARqNmimSexV0HVzjwc2c68X8prM
6lwz+S5khpJCNXyNf4vsHWmFK0XwIvJ1toOH0Ex7RfZaLQddgMMFSTys/SgzzSYfChFqA1QLZFmi
Sj+ak9v3lBI9hSoKJaHDaoa4Tr+lcwvZyKPTMl+KJTW2R+YpAWOj9qJqiytnuu+pE3WqZw97GyD9
u6jKqsTUOk3BFZ+lwdWEYs3hBkOWTEyOPAO1AbGMhTXK1qJT5zPQ4a0SEVpSw7QhUUVm/ac/WvDU
V5rsMYbgR9XPmkHdGSfD8iz8qbq7qrXx1+5c2ex9tu1OXnoj2Z72/u39hYCb9bRfPQ7iFlWQu0/y
9IFXzH448jVpDCFLNx0UP5MS5ZJ6Izm56l9BB/rlxp+g6mPMrn6Qf5ARVmVcjRrkdaoKtCYmFTr8
rNxb5CJ3vH3k6CJWo0ncl3IRj3TZlh3VJ0tEAffrXxJcvAjaFNKFd1QNWX2ks6Mu/mKRAvDU1jBN
Kw8XxQgwZJ/zywcxnu/IeuDzOgV4Z2YWZoyeNHT4RbqYxk2KzcX0tfaA8op3B/NE/FlHE5Db2A21
4w7V1meLVbDj+LUJ+vH29LZCsmkrdkJ2B88JPZ/B9Co4lUqLPEyOyHb/11Wu0sHxZd0t1XCVTXh2
rGK+UPSOVSd5tGqAYYa/Tm9CdcVpcic4Pa3DEUqqpsxzwmxwfzbpQeK56AKXdjJantUAcrubjmUh
UcrbCUjKFdKf0OcQdVWtRxbucc8G25bM63CwGnswUvIpJR2juNrEvrc/1/f0v+SPxj4U6najG83a
Hi+y5wh/9RGJDM0u/JbFSuNC0P+Lly8DYuoOqx2OjEN8USCpELSoq+FiNYFJvobkic5iEQ7S4SSb
I0/SbsgFqf4hoxuSnlDa0oTjtqxFfeVfM4+xhg7iLFJSEJq04H+ejl8YOyKZ2R1/KbVVFDjv6Yp9
+Xy6MUdBZ5Jm+nVygeOSIsJLDHORYqRcZedXnVhNYToCEChO5CBrWAVfmfkzsTMlEy0T3G6/gIA2
J/qPzeFFnfcy5Mrc67j5isJwriRxo4oQWJCTSsAHJOk/ZUuO0wrFI3PJIKwlRDW21Z3O7A1NqNKG
uuw9TXykwTwWaEklvyEf8TQWScqN3ySyYpbk4DgSEuYkClogXnKEqGtbu9cxRNkFuAFgLjI4HDEa
4An3lstI+l7Bdun+0LrVomdEqpxGZ+E2TFJS+CmNgj+M8GuYpSoats6cu9LNgw3C8iRiuiiXkCob
3iFGavbFKuwXjHY1Q2Ev4FE1VbMu5KgjJEU+yo1knAd4fDXAjEwlgQ6mKKP7fPvjHHWNaYs2ulh6
+suGXuaFU9XDEeQAe1YLjbDVv/DgJf/2DVas32umJ9muHVEgOhpra8VYiqdXG6EslgWCzF1F/oiY
I/hnR5k35tTrbIl+dSXGvdAMTi5+sbr20Da16xs7ipdF8wTmFH/6YM4yzwfLAlh4cEONauJo9/2p
0tc46ihMcpoMLnk//wlLQ/geJU+lYXdPHl6ee1bWW/0l32NVnwe0+rGErZjxXlDMfjFY6tZEOjdf
P8qbfj1VplXbkY54+/HWNJv3DiirN4++coJYc/2swwPXUU6rLFlmzSa4wGZIlbcPm7cWMr3oLXyj
/RgNHQcJ2T2R1ZXP+z3Hqva0WgxCQXGRL3RhGizU3Vy6/y7OSdVYaHw7EFNRiL9QUeoKdSfGtyH1
8FhFx5Jyozs24oSIl4anpBV9Dj6FTnb7It/mLzs8ORFVviLx4q9/ohuJ9/NgoIbGxfDBy0A7EHgi
xd3ebCLzfcJq2j5QpIFFmibuQ41vpe1Tjv3IKLZHZb7EVWEbE6l5pFoJ5oef6WAbRnE6Y+teQJt9
0FFlhFklailUvqTCGYLhVUwKUFL5ij9YUjkRoncLJMnGM9bHXdDRGJxxQW0OIgZ2sjPB6dxbpNKt
KW/XwZE9zzY9dtb24x90BlP5I/mFrzIZQkYeISzhpEDoynkYP9yjx2FVT+vphTS7PiwCSQRMgXKv
I1Pml2iqnk4+mFWN4EUL49+Zt0UPJAzfbpHWGVH4O84qfQhvVeOLwDx2UeXmXO0z/D4dcUA0TG42
NyYK9lMMbRvVcxLgqXlcB84Q6oQyhwWiTDfVBvJrNC7XxZZOebPMf0YqsWJB9eeMKgGpoeIueS4v
/2XPQT9LexHhV9WHRjsVheZz8vRkwkdi8QcxwIZE9Pfawe5qUm6OZkLlNx0s5Q36FAtPm13gqry5
6mNwOkAqm5b/EHDadlSPV3sgK/H+c5/2wVZ7RKObMaTAJy5wcdyD7BdX/XKPz/RYy4rjni6WY6kf
KEHvMEj8Dz4xUoeMebHXH3Q5tMLAQk6VjjYH6GPR0Oh6kvB/+LfGAUldBSj1eHkdIsl+OOBRVnxh
o77iwMFTfhXgs8AE687z8B8s33ogX4tnwvQ4/+ulLBHRqsPcShFgUcXiXAWZQn2HwI2jfTlIOIpv
CzjGtW2ePw70LMtXXM5css+eDpDEOyQO03xidCkG8FeDC4g5Pv7AuJYzi5RXEueuqY4EmVksORFb
m0BfsE1gZynCGCZ7zsFDQZC/KBJEN99CNykJAWsztQyJO3Jqp3icMlShWs5skjNklmdo07DESnIG
tLIlwLdvwMzAF3FcCNCHlR+CdKvE0F/rWZioEwqrA8Gui17oAF5vdG5q3ej9OW7hsNWrGXZPYQIx
C5+pyjaRiBHj8G/HBJlLThu33Rm9rJ+PwONXGIUi26B+PdJij7nnS6bKE4LSMhuWqFX+IbBXzyJr
60m7xTBMXFdMPnz9KEoRRcWQfjqw5JwYc/2uvctZfE9Kk1JTVGOq4Xtxfn2l/VUEcoR64zA6hJ7u
LUIPCH2X8ZU1sBHGdtZYHheHtqZKdMcQfO8Ny7UOvh32RxRS4NFSBePOOyuEKnFOcl+Get91yGPp
YVS0nJ/q+1S1Od4p+g9U3GMclIRflZhImFDSQoBDm3MoypaFxUbkv6+WPK08Zt9iAa3bqw/J0PNE
Lyg1OGxdx/CU8thWE/jSmFaiZwcJlLNuDBMjv/WrRiQL+VCOMw3GENwgnNUjzPTnvSGNTrd32gIg
A9Ov8uvr61K3L2QUWExuh8IZKnVFrXWcQx+M8SMWUApEbGAWSkTG1muggcR3gvt5F/fF2njX3E1R
TD6WZ1zMimYNJYATkZPluEpDfhy9uvFceFDxF1pkcxYhn9NlGo3rzeQEf+m21kSLurvJr6wvxtKp
5DBcpKw88P/zVZmqVBINhwB1XhJU2NF4qL0ZG/Yw77QtlKmdhXy4CznHAh+iboxHDPQ2NsGxsT/M
v51GKplBHYDVF32vJCEc/qY92XmNghlWgXxsjHpbQcyoD0Dxuo0tkzarv+rR+SJ8jXDn2qHuiX79
qfPcEHmVl0al3NZSwDZz1nyzqdZwgmo+k0yzhJVJ76JCxd8+PAsSWEM58WlZxSmUhpihmUWo6iTj
gX8Y0q8ZTyslZgUMuaLOCDcJCuLa6H4eQgRYvjMkOLa/V0IHPbrXisanktDks9GDuR8xx0gyIuKD
jezZq3ZK4vEWS5m0MKDCzsVFz0D21ymNlIT7Gschg/7YdSMMSfL8QJCIyeEh4KM09HRiinsptfvL
7ZmC3Oj1GirdwuC7fgmtm7fbH6JSikh2/10cVe354bgKeQU3ks4icJ1rw2Ei1+IdT2nQB01iHLu5
MKtrgML7PzXXneIHLllHz+n8spAsZnXVB/Sj1PBUyRppu4tJP2foFaGURDvr0tlbZztwl+nrHCGs
/Zl6me9ecmaGUBNIWrJ/VS8CQ/j+J48zbqBxjxH8iSuzL19pJcjrt4H5jy9BoxyE/ub4eGZ3NpVA
AvwV/U2FAzEU+tuLQZwMcdcsBz+jiLUpmdTxHK6GWIQBlVYpvdzaXIBBRWT8ZcVwngTr+xFy4oHC
nlFdam7TiTYvfaoEFw3Mm9uwXIT8PBw0P4dZNex7PBz0fjWmBeGV/00AK6eHcvMmBr6ZMUqyQmye
fuMSYWdI1ODDo1emz+Iy+Chh797nwJc2e6w5funkXIkbM+YIARBdP7FqEAb8538AgjagylMWrCdx
smQEJteN4/ASrBkdK/zNBuDDqR6oYC8/4iKbZJijLvglae1gF+BSez/xyehNh6VVVQuOWp7vyHTU
o/Ek5eRZ7AjJsCYV06+a3hPYX4htnBok7miNhoDwZwlhlJrGBK9eTIxM9/+Zi3dMKfNvTrj1ETo7
Io+PUsnBGpREFTIHFeZ6D3Smv4aQ+EpxZ6dLYcamXaOlFA12ifDFCFoCVtm6CuqwOcLinzPXXFwj
jdqt5v0M3RQ8Xs9gJZ2lU3x3Qo2EKXU4h8FqtUMYQPRBoX+iLOokUaqNeJlm97rDp2i30173MCqs
7JZqHkYc6dyc8EOglPnRoU1Q+0SMCjgbx6MNhcr8kkRGyYrRX2k6aDRHFbs6EVNgfPtBNUGbULA0
LzDYthZk5y3Vwo9ANYm0PdzlMCrBnpJEn38WXfZB2oecuuUMry4Oye87CgHhLslzattWDnhH6bux
VETMxq3IAuJ+UuGb4cNUR+peD+bjuIEy42w0nq/eaqGHe8tpyFrQUBiuGwqCr1Ie6D9k0wUjUxrf
A2oRzODd9smKRz6V2guJA6wDSb4nHfSWlmyXP72yEVcEiABtOKzwqp/b3Kdvjr7Ps5HmWSSbSv2p
MGZC96zCTjgqAdcivPtTeqtV0UkBLcM7M4jNP+KnkD3vWqHZ81OU/McYVFDBbm/VB6mBj4ykSEjL
Hj31LwHBcYXYehDLm7rgTI65wi3p8FDlnf7Ie6dORtrHBLjq2GONj0Htd+GShf3J9g4cH5fVnnPC
WcrTS7Zer5MOERjlZbXjFL9gTTer0CUnxmTJxPnv7yk/WJjPTldex1guQ88I/oxQqDZd4fXGIju3
OP8EDZHTfKFvTGTBbjuWMQXEQHjrKlkVpY/oC7CGso1/zIUg5DbAxfjbilL9GyDq1KVwb7Z4AU3/
qqGAklsoZwhlj4xSPqAYTYrJMXGH0M5+jnGIlyENAfiynFccl55Yeg2EeN2ltAJrRPmTBYxtVQeJ
DGHPwLsNMP2Jbf2zU18SvoRRK20I7SVqQyAObZpbHskztW07nNYo9M5LRIMLeP/33yjLVqxh42ss
yi+v7qD3nq1gG/7glAU/TAWDaAPo+An+mMw919nUL0+w8IeMQ2LJ5Hamdl4CCuC5/sg5POaHvS6n
g5PjTv/PnVro5GpwqqempBhDxMQkrjcDF2ottx/eqzuNWVc5UIdvjA+3MjFDlEo5I3iN7oDNB0jf
W3ztqfi0XKQUmiUNeohtIfxuk3JUzNnEAnrs480DboOSNS1KwMKgmohQjOLhujm5WbdcN38hDfmO
CzXLWyJ7Q3WC6DSpkqEzqcfdwk/22e3SrKnn37U27CY9aP40CiXqz0zapq5WX8BYOkuEldFGh/jN
kvhK71dV1mtIrMfod5g1cYLtYEataGEbm+Z6+jxwXRmUR+i7ctfKv5gNurq3ZY+s5V1TKfZTSgAt
nf0oDblQJNZS6lK87JI8Fh8XQXkzQ/f2yTARScsQimU25O3CBaAVVfRUDMA5T18SM0ZZ6aMmPtQV
izUXm3FuN8vBPl3PBrGEvOLq01jMMKEcXGERIS7wmkZCeqzfbb5sWD/UDZ8HReeC95LLwAu6MvqJ
aMzlGqU7naOp4cifEJ1WM3WtXLKHtoejYAZPGYfkDyaHfseBdsKmjEqwlL9u4/2xKIvmj8J37OR0
mChSKsb9OHZJHEACc5lBe7Ai9W8k92W7DQkWfkOlPAAF3fpOxlF1tW0LfQat17Lsr3kEUk1ZtNRD
OJ1ckJCWofz+U3idoas5dWG6bWc49BsIuMHc/4R7q9svxv2RiSzh/720CT9z8ajFBDq6v9+aLyqX
Sej0k7posQhCwx9K5WnrAfAeVMcppRNaoH6TkzepyaVE9NQAi4ciT6kXBFggIF5lOmEQeC5mWstc
++kBvSGeDV6SDFPtxJ10NISoJUwD+aGIShk8jWFDvNiv4Xm3DxXXvxr9KL6i8wGoNSPD9+SevkAE
MSpuTerRwTkuadCkw805aluFZIK8D0OrjwYjrNDinkB4BktNHOOgybp9wjXI980rW9yGnHo9Ywat
VbgEs5Y3A/FVsW8yZJut4k1zls+ERqF5gU0tduhQ5vfmfXqKuqueMft1EsJMwors0ZkowVd6LPAN
GO0Z0Xlwm0o2mbRazV4hNFv+EHULn5/009YsG+lze3HMbxvrkhcv4qpnwBc5JupCJSg/oBCFybrV
Sm2PP2CCf7Qh8Rm7ZC8xpQjrVWe7yXA+AyqrNe1SxNoydPTX/dHjkxcaDJPDUriHwS1C1LMn8BF/
qpKqykJftZ15mV0R/0OdZhIDwDfptad1N/RUxAyC2W7O4Fei068+myd5dEZa+Dex8IZhnRZWlfbW
4pfChZw41Ua2BsKLw3vvzYvQCX/59Borfso6ZSdUT6QPmKoV/y+BMhzyElqOv95PluIIH2danIG5
XroteuTROeMY5v+/Qq1dhwoE8V3ul+JLl+5kH8e0mC58AnYLWZCExxpz0t/sddvJkHWRqiXy9hHx
iJKXfUjEgUPwTKJm0m/6a+Wz723JbGYMy1xZRV9YcPEy5dh44qJ48Oc9Iw6Zx7G49PlGZn+t/1rK
pDn5HapnRAKBNIobRDOhNGU9pdvQUP1JFzP4wqoSCDO3hdNM9t1l4tJFC98MkfT6AbdIfT8W8Wqg
pckCy+eDHo8D3pZ1T5hQJ2IZOW7tAa+RiT+/6CpZVK1Gp5CS6wnwH2tkE1XJvqsH74FB+Qe3NQiN
bQ32hFRgCKaxbeiIFP1emksQU0BDDRkoKwhJLaie5aF8If0cOCDDRdQW6qQGtBOmozk95sXiqtAf
MUYi/rtOIwIVQbAKNWTnJXBmC24h5bh94xU+4pjZ8KX+s5a0hUafXRLDN/nuwFEHf3OTpcnVMxao
cNkcfSiRcwHmlFUV2eCUBVucEObt5Pq2soG60x6yBatOGJI0CRdPtxLqw0SzogrKtWzSpzR01N9k
I/f9zUndJwkaVK6Xom5t/Rt/17EzIhs+VCKnRLy64JgeY0nDIh0OdW6LI6kyQFfSrz6yQHPmLZN0
6YQOUzd6fBnajVQj+wyA/neoPm/aIQyrBuR9Q8HAZKcD1GkOzUqfIlcNAHTjJq0h3aHxsrsnh5Qn
+3X6W4VUqrDq+rCnv4D2W8eYsq2zD1+GTJPvR1xIHxr9XBiCMbINfttJG8m67us/fTEE7gRrOzsL
VoP5Fyv/kIh7/04F7woBnHGmGPNi8g9hE4qAY+KjKuRVEcrf05nErdHNECSskENXLMeyWURP4Hrh
K9JZF//BUMiHSo1mopvXzL1+wJwlKxugITDDk83ZNJokPKBp36KLFoFi8Ci7rifsUqZF00ztm1xm
ivpRfu3OISYECdwP4cvSbrsvqsP6w3/OtywcI4/1WbXIxnOck6S0OV1X2BsB4c+Pgg/1CZv8KioT
aXNiocEbczJHortdNYNN+ZnXrNktG9CV0VjMzdoy8sFfEUIzgSTxBsLKC3zVopEIlGBmW/HcUcKk
p4EzTmrV2W3Wj5mU7Df41C80lD8SOuneGrb5g7zjPEkSYuKtZHUwxkZx9A060P9EnnkW/8GHwZka
xAkmAKtHs2uev+hQJ9IkU5rRpODsXqREtPUUY0HLlb5BL0zOYuyS5uSEE3W4Pxow+6UO1Koy0wod
OJQaU48R8u7f7fVjhv5huctbf6TP7krkFuwu4vMIH8K82va5C5b2KKreQST7Zp2a74rLQFkkZuH3
PbTIbydj7VZqxfLOa+7waDmP0f92QH5kmJJdk+sKmthnSfkzgCXrgQEKVY7HcrywV9G6cqp06qwK
Dp1VM41bVku0Ohc3O0I8VcKvaiY3Ck+0YvcTH8ooj4iSrkRxi1DsRNBssnRu1TMbdCQRIHTvwAqw
CkcRnNa0e8betRZt4Y3/Ohgn8EykTgtOadMZeIh990oZK7sGloMTcBio1OqSDiFbX19+5HvzTaJ9
rGnDtv3QO9vEpPi/b01KGQn3hH0g8snXarvVOuUCPJubLL245M1RLDyNVwQ32xx1aBLuozw49zsc
HEospzpcGTi2AJ3fhw5TazNtLeBC+jea0vzlc/n3buScTPTVzh9w/MqFDlfMX96IHSBEa9KG9cfX
45ELivSkF8rSgLdH2O/DXpSVOYDo3W8nzCOGAtmMKz8/f0tu3hL0bgrXRs9ss+Hi1yDv/sfDpbHc
yAN1lD4Ht9oz15Od9RTBJyMCdTc8cAjpWRxJt09nz0MCjSEXDaoce/HyXV3iU2CQL8ysR9ZDYete
il4IJJzyRCdjzkyHmCSFENiLlnRiGoA870yuA1ElQ71JdX5cvfHjo176MBiIXRccYe7qbqTRwcJx
pKu/05yysxlpHrLWK0rrBhMNIBv8TBXvccaRIaw4BidN+jLYWOPYGTJ2IDxwmgBVDxjopqDLwC5R
9wsiRK5q8woQLU+t3UE7ibzwuIkCXf57SXwZUSBkMWxLbV2HPpyo4UA6nEk2x3iXu7UCxMTxI3WN
YhWmBGwSYdTupOtdr3p/2m7MeIbkwnH5caO6C6rGsx9/aXzuEJdKLc5hV1xMILN4fiybzvn9aoks
sDyAXu2Xc/Z9BXA2Xv6gdOzypsJt8cEUuH7kfFQGvfDgiEJXhkBHZhnX0dLrl+C1USUY53rkX0jC
sEYX0Z/8CqC6HJcHOdfcENkhsPC8tOQ0PBGAgRTmwNMgBxyAvu8o7Z2V2gQEwayRPVJ+fvL5baGl
lrn2iu5fPV20dQ4EHlvEqpt0CIkJLdKzFzVIIUBF5hOkP40MzfToTWqvbTBEpKnDdHpt9vS2nZe6
fOy9OwVo+/Ald/4RmcoUNFNaQcAbmRK9efEUzJpWRi2aPsbL0z7V1bUy4qZmqvmuMGTPJYhxlNzK
zdCJ6E112wg9GR8ALWSvnncS8vHFPBsJZbioh98izA93wv6Bsup7MnzuA7qvwj88ZN79TAp3RiYd
QBNj6DE0OBDKTYC4a2iLUgU7lqcTcXdrdn8pi4tNy4idQqBqzfEmcfOf9UK3j4nYS1gvr8pQ27JL
7YobhkpQu3MK/orDF0hw6lKiZa7FMMrY3R4kBgRGD0NBtkT5Pxg0qX/WnJxUl2/Ol61j5NH/0Emx
m33am2mM6MsCCjZQFBUdZDlSgSWMjRIIqaUTxujpbQtkI8vewHL0KINt9cSXlUsN+QTd8hRNGAuw
oxkmMW/sidGFAGu+jMrWGdsLhLMqTU+4T2Jp+js0MofIyL8ncDS76lgpX4eNud3ZrQ4IQ6bp5yK6
TJmQqBfBkEM24wybSvspWpDdEksDZkX4LCzvSvMfyzVa7WUSxaMMg/w8T91aRdtVDOyfKgTQ69/d
4vJPmsyXQXszWbOWy7JH88xmrrDLsQguC9VLDmJpAS/s6GoSxwcPgNtqa6/MyIsZk5nTs2OKNLRi
HdMW06OnZaJmQBoDVYi/MLmonu+IRYvTq7TIs5VpXdvBENzhLlZO6Qbaim5oaKzrQeG/eEIA9wna
VJvfOkuYZukwEUNyrPvIKY2qCWzH1pIirZkCPEovKrJTUErQyZUbCWhqRnaWfeInXof7JgNPyauS
UhbHtDO7JiG2ed5y/8Yrn8w+qzRgIoxzKDfLqkugIZWSVht9awqaML8PsqcSKGe9Zz1MdjhzNolp
vPCrkraFflim9fc7nY8Hh7rQVBouYIeVoKIHOyAcicQbQEvedBqEqLHYf+Zb8MIW+oKhuqI56kCd
rXtOoLk1nB7E8BJjAHP5+pcaY0fPi80uB/ULhjtthd8lmq/8beIOPj2O05Ykv3uXqFHCVQWKLfdy
yaL3ejhw/9JVssrDcUDzxVep6eHxMaNY048094y0PTgxwktIrKm9vZWU+Tbo+EzoVMtA3qhhHLOn
AteHY+Ue74KsL5Uy6SdgO7O1I/wS4z14DSWYEMu+M0FYsQfwgmHYt13J8u2VDpSOqC9tMa7TOgk/
g96r/v1IAqzZeoha7IYLHPziEGYvhKr5by0ZnvJD159O7CgGnmc3V6u4zYkUbIu4QmpRrKeIG8q6
ldjUS/AwgWqzBUR+doZbOQAM8BGQlJnS8n78jLc16hQpsnefd/FwoNIJVO5jyMPmHkBiTGLvMwTX
yyiRBIs3VCdbMKud+z6p5A+NBOXjRwZGYl/okgFo8mVnkth8n5EHcXbie1TCAurmZ95l+7dLdGxs
MYejVfSHRWmfDvujRihfMmRif2OaEi/94K+l5lHsNiN8i8PB1lI37U21FtuevgXInT/2eLW20GqL
ojCWLtlOyV2Vvbt+ozWt98/rlw4yohwDG7AP5QZ698wx/+5WfRLA1wzaYbZ3crnynLS5znPaPEdJ
6zLFyQdshLeJUCOhib81qkSWenDURWsUxLnHXdOFlgXwypWdZ24VtT3gGzHxzgWm9hQbzpLlGD/c
D1BXPKw0Uet61DhnDpX/OEAqfXHrcuPK/pyplA9NU6RjSUD4HZoLxm1+y9aVzBk/ZXHJPxQKYKP/
kpGUR4WyekkSy9EWihazfzzhU1TDIU7s1QTLPXsicO+s7kbAm0sJ88f6uQ0+kXT/9ylNRsmY3LKF
xGulYi6QAtFrBOeKbH/Isc8M0IQoQaNO4zzbBvYycs3dWKd/GVBwwfk9QbmUSjTeQqzPidzm603N
dpTCgYiUBHJojTbmY92xDYtYG6aecR8p/NHyezkQsVi5Q6kG6lfPORSsYABlvbSMO2lzwh4SxwWl
MMnmHzuBVUHSMlxTXmeAUkJICZBFm8gcYPgj5FrW9SVflQCWSU6HLqw8ickhWxRKwE3yXsx+HLzO
eIWpjsIG0FZdG3YxEqP3v6/2nSDtOhyHspGCCJMDffcwd9UHM9Obp+bW+1dLJ/xvDcGcMKBwfYBK
Q15arbQ+9wWzD4BPWdigZz5mrZG/WKSvvmgQg5d2LqjjVR6DsZm0nWRGMf0P3cpO3Ruqy51yMP5c
vJy577rUzEm0+I0sWHrvYKBivs1crDWb5eRVfZihXiqps6uYExG9ghZXVv9cQkt4PPYnfTyUd4EI
rPT8jJz14O+OGdxCB7VezBVEc0A9GW+V9ytSOSiqOGykoBT36M0kp7vDGW5rDhR0Z9hDhGHHmCh8
e0K2kwVtm6/jycBQQucVeXutVzthWSCsDd/weuoqLwD/NiSaNJvYFrNGE91jmRlfisSQcrutDuoa
q7/tJAanXJSrL3Fw1o5/C2Hl54d+h1z/L8r8N6df0qYVj91lbOSl2uWjBVAxWlTom21GUCQilK9N
BOhcx4mVyQeiF2KV56Ydn0FwQLPcPPQTIDZENogpunASJjfsbKEXfsmkUTh1uH7QPteLOv+ngMU3
dzq3X3qvH+c1JeYtbtNbvBzXws7HP1UWsU59j5hOA2XdCObm/Qkbw0IjouBVdOmMKmj0Gm4F0R3w
P1E14yX0Xj9rHifCCVSI27efZsTGKEqE5wbzE3NoW8fI9qBthJq3jp0SKdc+8/bZ8keBJKg/YlQv
qH6AkuOYWAZWhV0BG2gDMX5o1rxbbtjyn2i8IEyFpo/ccMuL2k5ky310XdpqIuKzUztSFaepdMjp
UlXXNfLwJcZVpuJHcpE2hODG5dFJaO7zFiouT5iQhcE9MX14BpprF0uO3xy8h8xQTmtZzGpDMGrI
CJIOXAEuo0hWOM1AolkN3bIiFHchP2eb8JaMiho4cA6IQxHK7irL5kIjpgUu0vJAbMQJ8AH2xMj7
hVvyewjNuyO8gnZpDOpc1wF4UebnEoX9k2inNUhd7XmFU5/5kXF0KLEqfpmwMTLMbroCxHRwhpWm
0gZ3cabPhy9dqLG/zIpNPAgR5lhQdRlxrrDyWo9Dx8rZQdRNRqxosdDyuD03ne8aMoaadN1lrR8T
/ZokXE5qMvFp+Bu/QgeRj8nBiIpjVjAudMP2b/GWxK0YJxJTPp1NTh9250XsSn6hdOmmmkD++Mv7
wKHs1+W13yQHNKZWKiKWRRX9WhC6b0vzZ9MOrlZ5MRlEZjpaF5WyU+RgD7J5HSyX4wtb7ybxrgQF
PCdmzjaVPu/6zq6eszc/ebBGp1kYPcJrQhqv+DFtLun2iVAakpab5NKZ9g8vVEwSw3jylwJ/lTya
K8L7OeeiP6mPNhA6v1NClNL84q798dQRmrQRtyJmK0UpRh0t274xwkfCJJENPmxUGmhGM9znat0r
0UsW+kH+ZPdWl4ucjJ/EWLJi26+GypnfOQ9tSH7jRs1OMmSknlFWuzPoox5qk9oSo0g++DbcaJj0
lMGCNDMBvonG6Xqu7apEHob7fDweVWxBbaiIky6m6Aexj7Gn0e9hiPAvZ0M/j0bn/IzvDMeyCdsm
hBFevmmuvWf+GqNlqRyHeanmo6bF03mE4j1v6xfumrDzcMyhz8dwFBscY0R7NgAuTVP3CG3CBNZs
mVxJAHxtSz1ulov+CBV3mZshVeyu1zqb+Ns5P2Kc+Iz0tg6KcvNoGlJo8zKQcx7GLgh1bxnexc0E
AqXAYqyz1w/K+DATG4RPQxhEkmHBWDIlpz1ofCjZFP3Q9kZQoM33kSxG84q31kR9iLsIKSd3RElI
TzILfg+Vi84wqgc7lPkxdLoDPWcOy9ad0xUlI8lLoljdQ258APNItWaP2H1nqGztp3TEwVrUWa0K
nypmd/2YzVvdlT7+MstQ9u/G4oyK37AXNGUpbKxUJGcRMpH1a1K+5u3rgCSkIEtE61AFJWApcm7A
g1aA8irm9ePrGk0cNxHYe8Wkt4jcouz17V+TUEEriD1yPa2rHx2ng2FQMJ8LlD6MQBPlQ15Nizre
EXklbgfWgOJNAdUlpO4tdPVDAlCdLmW1LHO81ILJ8Tes++XjpTeM3y0GArxQlAz1WC/W9INYvZiB
kqkWfFQUzhOa98gnGOHgBg5cYgEu6RuvkTH1PdH2h6D6fuFO3EOa7DqAKFSLmZ5jCilo95wWC5K8
0R8NRxAcOqMzYgxYkv/w2ACGWeJQPIEWutvRcpi67BVeHV2Ew6AfkAOqBsKoZUy7oK48GKMRp3bk
tHhvaT+w2bR7UK64rx1NHoaLxp2jo+KvvmEmYHQPSiEZglgbIgdXEAIaYXpZ58CBOZFETDpvSomd
VTO0VqN0BgSA1eHpS6OLiRMrdcjyxqRtKi2WrfjyG/ETQ5Qf/uOmFVGHb8oFJn7BEOPp3CH9H3YM
AUIrlnExqV6k0tKDIEQmgmOOMY9CDq4NC1nzeWmijsrvHkH1uA5+4h942e6/mf4Ej50sgErTUKKd
RSWlI3vOrBR/znA4bbXHiNh7cikN3bEQCzXcq00fzXFm7Fv+KvKtMFGuarJ3puv64mxzqTLbtKri
ugB+WPi146N32w87H9uNXvRmameIYJUBfZZVrc4nCFt6FVhKtQq5H1h/Kvv7NnzTxQgNxG1/pFdb
vBfTa5Q8kuHe7//DMXaao0dLbwO6HDNlBNxZZwPaQ7tgau38cXfeE8UPE28cDBMcK44wspByz6Xv
Zf5itSjigInnuldl2VUXrJHOmv9/IJ//EeQgaZVYq2BKL/kO84/vK6w2VQH6Y6XJApacvYqwIvrV
/BvCE9b9cG8fK0itbRzzoKRHw6TjP4aIsuoFIGEEIXPn4CrKEHM1dDWr4AvgSnUi/lkILvnXp7fr
b+FEzQO9aeZk67prG+dDEMdzwMaFHLgRL8CyOpVoYAUIoAtYyrb2tQXYro5adea03Ichp5xtHrNh
0g3EP50TvEU01PvwyyI5jeILjWxi24hpJO1g5wT5LNaosvoCdB1sk+nUMeAVlCo28KmOvuYlvPC5
W62iGGl8lOXS8d+RGjMizXtBnoE/niU2Ombk3OxBwHt+edv8PU4NEut8dvPV1c+N+Mz/H5tAjDEu
390oiCeCko/LU4KvF4mZTiV3crX8jv70CSh4F4Zw/pxj/Q7VHFos7a5G41cNPMhDxVVZ8HedfqSx
CPK1cLyX8CqGWwwzQDfF+pTJ08CyAM0rOvB81rS/WQMSZZ1GD6tcCFSRGc9blD1cjQhFzW70H7RW
XMJeeXWhzNGObvSWk4GYT8t6BD4HkmXsmA0gYOEMgqpd2hTOiL47rmHV4nFHfWQtAYlIP5UdxvRe
05QhTk+c0k3heJ5JBavPrv/cwv+7MChr3q10mxNGxxgShct2dspUGHBb+IUO8n0pW+5t67oEM6Zj
EoxQZ53mDOCMUklYZ5vW2SdCbty2FHg1zHcN2T7Ihb8qadmw4pQx+sLhIkAmI8lKmh1FXau3etAi
7XmCitsVPuAPHcQm7thSZPW8QW+UDMPes7CfuMQn0olWCdFspH92z/F0dl6r3yIlIliQIO+StXM6
xTS6uvVYcmmLh6VMXwKoqWpx++91YXQRV1cSlUF2xr5nhfV/uVgwZKGcpaCZlGwOBBBmEPjzc86/
CVWJnXdU7px2qTD6eUimCfd2x0hr01h9S3SqaC2m2C1og1V3EzipaFzZ2xVBsxxIpQ4DL3fFMh9R
6tlz3cV4DvCbPsogWfM9SNK+3pD/Z8a4yv1I7j4duXNxjUNQUB9rZk/GkmVCq4YYg6I4cYPTLA0m
MuLDMdOn14YoUH5jOl0oHvz/EwFvESOQkI2uBT+SpLJeV4qI89+y1j9FGFAR1zyaX5pFqnuY1xPj
3dvvDVZ/nxuNJnIIUtQQ4Hjgx9Xg62qHPk0NnOSUNkQFZTSm4AHrZM2ZCZSp4UR7B/d1RV0tXLuI
zHOEpKHr1fn7zdW9DH9LGORYu5Xbykg2rrdxVObEfv6Y/85RCer9x7RO4qLdLg/vm317OajSY2/c
bWNA8dHpNp/7WD9g9W01j4Gi69kyFZsyU7JJ0Y6eb+Kx1jkcZVQrJbTHWhcAuZDQxchXq8x1r6Er
Y/osXRDwhVGZzZMH6IVshsPNB4UBXroqWN42z2l7ZPxd4rU10aJPHbehPrMsqUP8ljfIhEwX5tU4
asVZfsZMrLf/9N2aQS89mrQk2eHM1lkHjz5E+viQUsYwZJ8i2D2J/vfO4toE81LkSWWPxgyOwRcE
4j5MX9hxE/YlzLifTL5BofAWMFMFcZhLOA44S7bJ1SEi4WSLef7lj93pn1I/wzs/P/+BLqoAxFyp
ueDh5YUmNOxtDADDtWC03BPCyxhue5jFmf+ftXqHaWj3y1QR2RV23o0WAkGakK6Ie3vIeXfuhcVv
0GoDo27wa94/LSufKRs1v1LZrMdf0ewPRk7doXsRDJ/RXDmxSDPOL4OQKlUJDzhPv0isGODctftk
IFAdRQmb4e/+J74EavdTrzVGDClNd+nkjJ+Vvp93gkEbX5KFXbmnkn0ORwtdV4L8m5Ar3Ga6BPze
k04oNZhWfQ5MIgB/BMsR+Vyqjj4ic8karssApugKMVudWO7zQhQHK2ye/LwCi3vE9MUE3O83fNjc
Lgy6+pn4Ej6Ppp8iP2dNyrteNOj6bXf8ZX2ywsOm0WGTbNWiJuTAfMM0bL8AEZkKKihx+sBoeaIM
rHzYW091OUMjJd8GoM36MxK+I7Pxn4LWz9lUzSRTh7bcx/zX1bA5qkF24WOexevo/9DEiEeWr2Z4
aHtcQVxJoLC6/SnbUnPaD8u3UmDW/plmUkeN8Yfc7B4RiCglA9ufgDw/TLKVaw4Cmh3fWSFDf87b
B5WbDX1Ah9fpj/CnHNRr3f/iz/qG1rC3X3C1AZuY7tK8vXbY5HsVPmOyhkelkTx3bpKHWt+j5ATJ
xM/cmSMr7M4CMRqeNBpWXS7+xyIQf6DTonLKzsGxXvAaUn8ypdRMv6t9RD1y9Q6LNcE4U69JHqQg
qdSkhS+u0qNB5hI/dlQkJKs20I0LBtSRCKBSPPaOyie9/JqckyZXwfVQnHAkoSJmiPAAT3nougDR
nGvxGdbB1zbQYKLLPOLnhYP9QKVJdP7iMoiKAEtpiGHx5qDHo6Xq5e03Bji07m/w35uU1g6rTJn/
UnlcCtnN4Kvq/8GOWCj0Cpc1r7jjBEWh6meav0IDw+k4SMzHyxmLc7L6OOkZF8hCQ2YUG62lc7nO
Im+KAgYNxy7LwdwtK3Y4feSyfPdz8qq5CZ6JB0Hf5VtsGD6sGd5C70nsDJ8Cuif64cLOBiY1bBPp
tAr3ya/aL/h36ZmB0Ow/k4UGRXFNc++PJCBOSCGx4u/krkQlwft67lR8DTROVt9OgTMrEP/wef/J
MPSfG7f2t9k9xRx+R8q2BLXlUgIu8WIMfjBJm+YByyVUrK6guLHDSA2iuGBV0mRn8Yg3cvVXqjuF
3aEKdpcKzkbP0KsM6Cjg5R3RCMPS+5GJbPv3/OQaKxTCXjsUNGf8sbGXhBlF/PK5C0JbJ+tc/Yzc
G2W6y7hi8GNchMPxwQpc04SuHHZmv9KS/0AQwnl35/eb6RZ0JhTrWD5fQCJZk/H1Qc1RhSpkL2Bv
A8ef2v73Lkug/M7eMy7fJPgJ1Ue/H03wWt9fa5/vg/qB7EpGTJQXrenJNST9GenOSAlzHjtrV04n
/A6i/PPazZZhcraZmJrBJ9cF3YGosZIFb3Qt/Z2g/Fk2Ya9atikPBdSma2w5DH8rLolZ8ki4Xjp0
gW7cssKeDn8Mn0XVcnLtINAMSiB8TkrF97LVcQNElG4UF5rSGunTUb93OG/j5/Nxt3WJi0hU8nWp
bbaj0ExB/K6/gUBvlK/l3TWpMpPrF47r3U5ugQm+cugqigBFY7H0M6LoOPmUNFvG0ivNL6YpjSKN
Ar6UdUfxhV7EEehl2kXiKJGDqvMNTUNY6aufm0eyTFymqzgpIqK054k1KB9Va9fGANKeouOLGB33
B4ezxm7dglx+t2WhfYpO2qN8LdmyQTEtg5kpIa+lMJV9fN6rSrp0sfgbyY+mZzgSmsRh8JWvfMPk
QpWTFMyLHcawtQ4nI4KS7zBXwhFBopB6ZZe2U4CYEdLczUmRenruj3bfIh9UuYXaZEvH1M/yyEPi
jO8L+EgwJf2YGbNFo88TiGO51zwsdbN5rDsQ8CYG9Tq9Thkaewv0XqU/pxuPrcHcD1miu7mv7FqM
6Scyt+NkmYqG05nnRP46b3kf7oCuUzXpAI49JiMcBgmLnzhFMIpFY/R/9VIJFyqfbzUqVfL5ws9Q
e/Mdsqf37flbMLBn8vRl5FYHsXzOr2nYyu0q2zRBokmQa1eCnsNC6wj2SqDUJG+fKzddJ2BvzIlX
K81ov+snrMdDH7qwPQ+Ba/PCeiNTvo+1lf1vHXaDXZ/ejcDl2DMDZb//KL73LnZ94Mb8UCfviuMX
Ns4RydIe5qNbpOcG6tJqE/lcXeNEdio0GpLWuHC6RLE4qye5fJx4wo7kPNupCfGyz2xGM5Y3aoif
vkFDC7a4ehlFP9di+ILbUXaZVPQJW250GtJYJwN4+bfAtSOeDmG00dilaMX+BVncuXmWkEwR4gWT
D7NynMZiLrQ5/TnaEIbQNFKVaxH4Q48kecNiAqBjFFYQ/7Tzbyt1k6e4gXhawr1tM61p0H6hQ3W6
HWzHhtKTfKtd7zPuj7SxtWmqeYy5KeJXAtq4jjok7wm5XFTzdhpcOAq3kvqIEPedEXYcmRMLc4lw
WNleAo4CnZjodAUElt8z1rSHRnpQBZhcvCSam4wovtQ36s695j8slci/jX6QKG52otvguZtf2MCa
OnyNbd4WQY13WDOua+N/hLhYJgBacI3F8mcrkBPezJMh2z3fOKBg82BwiYUyxSKPuxsrjvvk/4op
m+DcplV2SBavS0D7at3h5oVeZV6Bs9CUwoKh/EvTwVMVduYlHZ5axbFcIidHks2PFkAgMhMAA5h6
KDTovBeQXMyZ/PgzIGxOrdDF1pHlmfUPa3aHmJ86TX7sdkjfGGBpD8DuGcNLaKN6dXiHZ1iKXwN7
P5CJVQISvsAscdTpz5vo5J4wVwnmY2USIGn35KK9nPNHZZyUyMkCleKtsprWYVbufBG3Nj0KSkQH
Oy96M1F1qzuYc+tI/DIHBWDBSBb0V6om2L7zbFZxyKPAFPQyg7VAcBMvytaek8NXwlkETbt4Wqru
KMoYmJCMt7WelyxT24OuFGZh55z2G0oSiQTtTw7Oe1a400o/ihpBacb6gVgr4x8yU5Stp+J2NEIP
lCy4u7hqxfOOLetLoWmFC88r/b85JqYxbgdSxuSa/TFo5bUbhicJQyJ7UtYPN3or+NLXcskiY0lX
3K+/TXilaELeojLSodP4c5iHDXSSb/4j1XLBRN92I+X8nSc2d8xO86spC+vqx7aFbL+dkkrSPNyK
wbs5nezSNHtINceQLYTpIa67A8IEeNMrarkQFjqYA2zUXcwX/4XeJH2O/OzIUWcuTBWJX+x+I5M6
9Rbs7TFp5K9VWqpHGQmgzi94u9zQ8QjZ2T4x+y+8QhIwGFCkP1vg+8vDQ1YtiOgXBNF51KJsfznE
d9OdHq2RCFGR0WhENsFhN9tlevRttm+DG5cu1HkDDBsMsDKMxh1VwSqrSnrOqYOpk8Dd5Ct2vaEF
9TJbKkCLGYiI2lWSmccYgUXjidc7ZL0Z6uyghUOIrK7/wESEbbBVLkkBbKdTBOoL7qSWuUN4TPpp
rSjgvXnIy0MUsKElI0CjpkhTw4qF+3STKbiC0Scg2PN43b7m2NUznqIY+KdxkQckivs+dd79f/WX
NVjTrGddfNXfapzxE3GKiqmuBXKQix/Ea1ncb3pJCWnsnTW2Jfg2h/HPwzN3vrkelz+5xOM0cJRV
WoCHh5ug+CdYyFwrssq/LgygltzhtgI09LMUBRP5L/OFYdoswGN0fmFGt5kGY1xDD+1mM54aCu5W
SUN3+qcJ8CK6zVrugxJmfAyk3Iz43z9I7Dk5fb4CI20EySG92/rsdtZNz6dU2gHnja3ecAsZLW0r
8ICuSnW6aJL1Lg3TBDWS+TlMcH/4kYOxgzdG+xYJD27GaPedfvvddTkRvemxMEThByocS/XPCwNZ
LVMDXHBgIGt2gblEHd8Ki3ElMkIMCwOUrytFHxci1souKrfHC9NsEeK7OdFXf2nXcPPJ7Kce23vU
gO2z1LajSwWfbCZT4/J3rkHKs0V3cM60FLz+DF4ymZjiMWM4HIxIyC9NPssT9/N50rBR/V99eE6e
wKZMZUUO1klx/PVeaa3S5O9Tto+o0ITluPhzCzfPoFeV3Yy0lKa1DBgpaw7lp6Fq8UVhdA0RjYuF
5oaebfBihanlgXnsbn4QR4n7q9E9l95l2zKDFagzNTt/8qIGV/7qgBw43TfToxh0qI2NkR0I7X6o
TzAQAQrzRWrDENMIQflSPVsn/2YwOozv5ee5Fj95YG3WP+xABdmSWDX8sXT6Jxc3goFyaVDS+uGj
Og6gORv4cgcscb5okJ3wruwNYP6+cFUuvZwVIoObN+iTybdtOmZ6fr7Xq6q6KMR96JRyDtxvkGS5
GhRugqLYxSnip2TRyma5fprPGyRbFy4zfsKt23+cB1doTB/pWu0F5DPOlAJaRjzXWIOOUozzDCVt
t5uuRt49Norp5K09PhzS6Ue00p3evtmJpTvUuj2RegEfHgUb3wBJOcNpcqfA+xkqykuj/9HUmOxH
qfK7rdt2x1egxlL51x0ETUF8fmA+PirtE5/tu6+iVgU7ZCgjuhBLbjDJYbKiS+nwBXm/yykfoYzZ
LuVPdFzTm1f4VXP8xgiqzTxF8d670O+0gbMBMDpprzFQq46dR44ks7dsVxJuaRBcvv3mZAwqz3fZ
WhOpTohVgchdT15/Qp88pcnQ9c7CN88FFEDWEOu3V28RdUmVaNEI+r64xFBhToObcxFH8KmQIFRE
/+8UTGNTbbR9wJlKF8+PzoYVV1ACTB2zCSInc1dBp/OBYh947vY0pgWEDLVY2a2z3oRrHCcLZut0
biZsNkA7TIzZqIleoDZq3f83zM+zmUnZnQfFQ92VfY7K6p5oKWv3VhEulpF7uBsST5e2lI4PDYfD
9jDKALxO9PYGpP0rf1l7SAL77/JCKWWTVTvAlHAgZm+T3l6P+6C4gRmsUF0Y1z1zRRx/55o1JBn7
ftcQ8zXVZqKxiLqHfz9itKwM5s7AaSRBLh/fFtxRJjtF2ZbPW63zOEjVam2iOuK1oifeLVFAI9Kw
bkLSK7m5nj0gNGtRTL83WvZKwWr/c2g6kC+Oi4GHAIbLpN6XRIq8koDmdHr0qv4BP1vtExtYRvkh
OcztDIsWOQ7AoVNZqIA7Pp0d8cMeXtvPibE9aXqKTQVrH4sN6YDfbpNsbzoYcE4mpv5RQDZIquH0
thaDOv9mho12r3Q+wamUXhQagufjrsB5ijYPsmZpD7nVthRv+ssEOhCEAm2Fwm9dCcrJPWC6LU6T
1OvryhAArlyVyUFICFYwBI82TdbtggCJICfsonoTU1Q9edpbkT7aLTt3layDTGX3kXen0aKDOcUA
8RMIHEy88N7AwBYhR22+/lGLq4R1mi4eU5skqYH/nFo/PlyB33T35OZvq4TYr4Mj9xPj8LUh/bx8
Vkx+UQszj8lKQgsBup4d6Rrvm8PJuy9Hy/NucFw/ZZ4+2dARpzdQgsKX4tZsYttexoeSVhNF2SYM
SgkJUVyQppVVICCOcwRQ57IF57QUTtcQeeVgEqEMkwZlHGyizubTar2TgzTEfQml0H5BrpLZuzCD
mjEPUNJryUfaY14Hj/UzTgZUFlV3NatLBp9PGiLDsdET4UYPWk9h8NA8yT9afixg/Eyl+yYrZY5s
jLCabKhghqYYEpjt3qoAeiEXfpQ6D2UGa+ah2RFrbx+mnDldr00KWutAMqe4wuIWcDtWl6c/LfhJ
LhGOt9orppzJwNyKG27Fu3o+hUkoXgBdy//oJxtPZjfwNvG7+j6LwGr/qjCoD87FmBO6GSCIYcPh
LwaKa86ha2hLZN6JKCP0eRSFi5VvUK+TS2vH462+8z4JoNQ4w03W0eQu0/iDC72qM/NDT3pj9oVX
4X3ptr/tOcFnYramx+prpFrMi7oQ/vTUyer70bFgXIvU5aPJ8L4/KIdSwfc2QU9upH8uPVuDAvT3
vK/x3ccngHW13qlMhUuh2rRv4Hd1g7yUY9ym2XZiSqFbwWCX9y/73QHM8afzmSRHnJ8BpBlsn67V
PdupqNA4gx+SfKUHcvmRAh4YoN6PXcqWHcByWNsIXrAiKf9EufWT9t4vFIHuhxlF4d+9f9CAfA8S
mSmIOet0dDYUKZFRZSpQf3y7xpar1J+chlfyKJAgMlw3zYzy6mtYFde8psF2uSRbixYkcnp4SH8Z
37dWDT5y0jIMaCr3dTEmPCZXXjbw5gZBKam2U2yrCd+0prRTkpEtoMjTeMUQfyVkP3bp/tbc8qWG
+kSTtBA+0du2vwMlDo86SjBULb0plyCllelg0hku48HoB4zR5plq4zvvsTTZ4abP3rz326MMb3DU
6yjbeFnMZnlOKcHq/jjASrYo86Ga28o0PoxVeKM44QeiunJTwPFUz+0Wj6lOInwlAhcFzUKVDu2k
prG263qK87cA1i+tdf+tzawsOhW43gJLimXlXWHsCcaWYgEgg1DuwW2nhJYu3ZOX/ypdxPltbBky
V9Roaaq32Wx6y4wvFfvtlAst8ty/LzD5X7Lr11pXFaQyZPM6PR6SlYP2F3rKanr04ZmzKI9ZDJhK
AkyVW6lPb39UBnhMNTTlDnYC/usP4VC3EPN6vzXLaobmw9NHg5k4xEDI0ckm0cNIthCX5DF6HfDg
gDZYxVLQNk6AS/9XGg59chZ1rRVMxYAU12y5/BZwF6JtqbVzlD5kfBGXLDMvFt1ZhIHQSq+0Vf7K
fQBp9RWh6OwU2mfhx2iE/qaEfYKpXCUzJOonsnp3AGlyIAoiH1CQw2LyrwbsOsAb+DjG5Kl37f6Q
AFy2rkm2L7IanNHOLwPD/hQ5+iZmY3N1kIjA0fEl+zB7MkNBzdiblGHV7FA2pgKNLmYNEs7IqWZu
jEtqKnO80ehKxMYCSp2UGhcbllffuRhDCQN2jkKtNmzgLYSUMMhpPFyyWsRCTERyHLXNhLUrcqgU
SJLeogiJ0otvYXeDfu+cgI2nnKKzu+Br1lhNLbKjPDwfBfeY4Xh/hAMI4nEGDLYUUhPH5yxdZLSd
8dMJU0I5o6BngfCQ4/fpmwKwk5VYgB5AjGwEtBBeZJEZpm7P2veYDfJhmeMPWO8C21iIh0adTIkB
Cr+GUhRD1080arYsSyeI1zFYeiCEVNags42Rl7gkfHAmJAo+8fw9PXy1B19m+6rm9WybEjOMsurm
v0NtWLZaw3j7fw/TY6bsm+TFfRSvAyuqTh69RxtoMMII3rHVs7cV1xRjm66U1kGKJJ5b3MHdGACd
GajiaoTzfiNcLe9GCQXpQFrueLad97D68h/PIhkLaj6Uap2zUxWVHkyvjFrsczS96YKt0eraExx/
rumN9Uor0Jksck6yY0uZV+Dt0s0OW1pfmH32ejRbMMpgkNBISOhNo5SyrblYFmYxb7E8bITe++ql
TIKPNL6MyTffe8ZVHg0DItm0IzHw76eMs2GevbKwYiUZ3+6YwPSyRjjSyePwT1Kd1G8GuamhyfWl
5MTAwEl2RshRKNe3wlP179x3VD12nOIoxIajVWmzL9UpAnqFnCE5yipxD4x/pbYAtg1TkTfY0uKU
tf3MsMAbdhktj2VGC11DzFB1XfrEgCZvmGNZocxBODkibnh7YEtKBvDbJ2k43DZmp6cb0xPoYqGG
HeoSURRdS0xq7tP3Y0QJaifT3h4xl1ZZcTH4cyubvtiKaa84JoSsQtfAxWmQAJrSn5QP2QNQaUIm
Iv0cA774b6mTJg6nY1XZvnaAWam1Hkim3Qrx2MzmP13hPD8tWaZJao4h8XmVWLsV++a9WJ4TQel1
+ehIcHHZpL5tUIdNEuLm+xol3jflbeYfDwgQfKWlXW+BA0HECTXCdWrk9D2V/ZEjAvPYjE/P2+gu
F1zZkuD6EHtUHAofKQ4Mi9SQFh4PugTiQR4S9TA+1lTB8cQTPgi7LenOSNRDZ7NEHMSnzHmIHqvo
z/AM+FA0urPUp+/hbOuu0ID1rhLFb9sLaIrUmBBV2M7r0z9CKp5a8ZfGzR7zutmaXXuQNyQP0Jyj
GGGR/95rG8Kd/cNO9wbpdtkd71L2xl5WxYZwQStQ5COimon8Bvfs35M9E8m+M1cE+ZexpNAmxxKE
Mxwy0AkGJf1R5sRj1uIi3DPJnbaikcerCrKYH1HcXFHHDx+xTngZy6NC5sKFa5uAjrb0xk5Gy0xM
Ua5HvXfpSfLIMbTqVBlxVrTRcX7lYp6+rTyth5B2ERNitSPRtk/Dls3NyZun/IzvJKovh2MbB9Pf
d8ClupKm1KVTuV3sMTph4DaY6dG4UNz+ueDtj+qnQytYxa7TazhLVCCpN2PdgsKU6DIqw++Mb6I5
ffK6xUGcijcLRFT4ojyNQ4EvyHquuo+ku8ooMOYLEbspnoJ1L3AVYThWNjeSUy9aqXeam2tPLw1A
dm0c1w7gB40aMpuZH16dUf8f2yLUjz9sPCN7s3ZjpQf0o0BxiWX5necLP2upWJsmkjRQZTe+kFrl
ACfFVGkYztmNz2NPnyIqsrGTJudsb/oLEhQViKBMGJCN7+2txR3BcWTRrWuYNdm+AqoO6Zt/Uf3w
h7RVZhP4r+F3491C+qLdvkkFbxUJZJZlfk0bYOb7C2sQkjNTvBoR0kF8l43Cx9Z2K4uDdZZk0Uln
+uEFrgml8a4m0OclE1Vwb8ft167TaNhnvenUptwsQD64w2oYEf2o1vb6D0992UwJ4oG0TrEJktJE
5CYxEw4Tm/pwg94zdSPiA9cQRgRCNTerDiBqbIKiL6PlYw/NKxiaGLhhxgoHuqC1Dl1whH1Xf6+e
82jVAAkHBapEqSIT8womX2YYw+5Ewx6KQiLznioHHrVa7wJ6cOE6P7HBOILdjzeCrXpV6wCgKecq
+R6w3sI+it6MMtmvJMw4X+PqwqMQmCaliXMpE7r4RkHn2psc4YUP40DRXuJFUehtZu7WGiu3o1dw
R/MK18O0+zSu8z+qpge3YxNiJ49Jb2U93EQDZgNqnKIFbuXinnHH/iisDHAYzyLPn25t+xQ/IaQR
TVg3Mu+uQj5isJIgFOrdnCQD6ydq7KrqBwk0K1a8J+8RIaH34BIU1gWiHD/6bOL73aBfjD9MzmNK
WgpOFSQG70QF9P5ILconaZ80hzSchbfqDyvgWHX8+UlkbD1b1FWQ1lH/uggdKO5bSVF67KFfkpIK
mCRAuZQGjJWqiSDUi2kHhTDrHw03zV8/OFUDW1nORhvGH8r2coKOamMnG1iaSahTb1JE09g5qyqa
++OhiIJ/tozwzLHhCPrtjIkaWad0154JDvQMGSv0F6sEUXnhuA7hWxzMP32Nygt1C5HwY4T8wPF3
j9OqA8bNPLVUCOmpS7/ydOj895X5LoVfgr6jyNa/7y9/2uk7qQjzxSeoKi5hFQuwPJARYaC/xaNA
CI0x3kgJuDSDoH1AOfmNcb8XplJDjLlm+EFMZbAMm4aAAt96EvItvbeDM/N00d+aLQsnWeRWoOBp
wnBFQCqAbn7kzAAEiXHEWN0M3zFo5wdbPWQKYhdKZ6OfOJtBz0IyaJmrV2Bl+9MYAr3Dys6sHXmK
q8LlqwxJW0IWmwW9HVwlffp+4sNyGPny+r9niF4mu1IJdGryte8B0iwcf583NBHNIVQhW7vEJH2Y
0lGZNVg9UKobQQsPWvPkW0wVqtRXA6vD5Zvo7xqSt78wCI6AP8RtxZPGmbjKP8FLRj4nHTiq502A
DcyIVUvkxKXmWnj4RIJeIKm5uk79LZDhVbphJNwpGFWR/6K6lyNkFOzJPsKrqTrZLH47uSnP6qmT
RvMJudWtmQeTRG9P1hL4+kVHQemxhJYdeIwS6FYne3eNwzWnMRrkYwQLIWBWKaENrP8tuR1r5Sm3
3lQJaJB8KAMICxPJtAGwKt9UaRvmThlyA7vdr7UmnEsp9AzBNvYzD/Kr+LrfhpxlVeQXRbaedbJw
YFj+Pwkate0oczkg5LBiPcnLvnoV/KRKJX2g3aJ6bpUJwKyNkbUQ8hySGwK42D8Z80TdsirjF9Uz
lL397wFqTQpSyhWkyl3hHaIZksgs3dIO91GG/NI6iQZA+03xOt/qII5bNTnGEz0PZI2X50ZHO2aB
0UL1ezQJZU4HNFR0p6CxrVtPjbOetEW5WSFWgQPV/jSlsaqHTi+BC6cWeHKNQAG/AO9Q0tXoIlLH
mzz8csuhDL78nknGwUfDC9WlZvIKuC/X2vX8WGokq9e/o2A+d1yCTTJJA2o/Z0jRTPX271Q7M/cC
DT4+oEyLO7Fh8XpU0XgZqKtSV04MTAMjeSXiZG8xokpY37ogrw5DZiyE7ypkZGzIwzwkYYh7CTR/
eXoqHNnfvRGQMTiPYx5Os+sBV0moSfEoUogfhkZ3oTU7Tpy0Pa5U+VSTJuSS9HsWXSCrhF5mr2Fh
HIwhMZSo/dsLeRK5VjUXQThB5IhloStDlW4TovtCRNcRBcboIC+JDOOQF0S1MZWgy2Ww4VCgJ3zB
qUSSYwz/rRRok5eU6ZtoSQIKhNP/XI5irYkl5JZZsuR1gNhA1R20ZvAIuL3Vq/HDxveRZuQQujSX
RhhX8ao8beoJstQCAsy2KMWPg6Oljggf4WQcBt/fEInJJW4dTbUmahoPkUAxGu4OnKnEnrAZ5nt8
7wCOEzkc+GEk1RCnosqa/DGyyYZrElKGEe9udvcRKEqkaCmnv1W6Cjz3suyAjAxM9ylx1q7tTM7A
XCIzPKf1+J+g9kd3uBauNhyaqYWSGZayhZub5nbjft5ifl+0L0tKuJsRsG6m/2WwaSkkunLJbDAv
j9YuRlCeIKTN9SHqtTv83/DY7v39qUw8GfkTWHIt1U9NU+8/QdnsGGTlxUVOXoIwZf8AW5F6niLH
82kKxWnrXaGmkntn6fGDcDiWo9wt3oPGwQRYAztvtD5AOfqW8j9tMZ5jR6bqYRCZctxJ5ezqigtq
qcDWECV9IVsqitOM6I7oCwXa6Gz3RdX7KHIHo100Q+v1xEa2uERX2XyRdLHLfwi6T0weTxd2cNqR
c4kuMqGpOAfLs+VkDRQyTJ+ue7qcGvjF/JOnnBFcjgcoKTht7Ni9EeIRW8WJ/7Thxf5gZFeR59vv
0CsaTGQe4QCG1tHp792esVWLfp7XxapErnpnSKv09eQwYJ00Hg1PacoaHspWKfle/OmQSsXh37Dn
1AEIutvsMN76LRIXqbbNHwwF+cU1NjowFRMjH77wZHJtG+1PVV1vok6OGsibHgrVlGS8XOvxUTqY
73JB2+sS+ggkYaFVUai+LPAGuL47RxmBnQUV6yh3d0VicO6+nRxUX4HD60LcsSqdiE2cTwbolk23
CqU+O7iaU2rorGGfs+rgr0q4bIXSGyfW5G52eTVIhY9rY6NLPC2SaCeezn3/KxvEPQGyvGuVRd1A
PuF1Sucqt5miKhXFRnvIIe44AzCRO0Fd6xTT22maaouhsBENFENIFhPy1S58HtU4ATaSmf9EDeso
BRb/V+IEQ9kaEHNPHgVv7fYtUn1aIEqbrw6OO8VyD500bciDD7jKxRvfHDVxzBdknt0ze/ZE2pIX
O5ksATlkhrBz2I6IdMzOYbP4pOnUHnZpozOTAVYWG6w4v778YCx7L/Z+HMwXSPkO7cKuLiTTBiTB
X7/TBKIt1hX5q82cVP/78rt5Eh9Gy/LkZM8tQSbK5h0Br22BgPVZInToc5TsbJkbBVouUatgX7EK
Pt2Ud8bZzUU/hZjJLbKoIOGAlMcbogPNaZY4/fYY0wm0JxFfUuu6+hKPHl4vYRQflImJaUiM8hD0
CoAbYqslAPQiuzEVhMO6h3ootBWC4tPXmbn5FboZfXvgaYpIDRJqMK8attkLyniTwt923kOH42hP
wwaM0tjT3H65w49C1wWD7oWtvC3HjxxDvfFKVSbPodxHRmR7mAMHGxUHtBAq+z5tCrCiABgF/Psp
QiKTfzjF5DHum155GeHxS9JOmr+7Aa97jFOjz9HV6+17Q9Jys+FPFFcX+V+t/lYfipcZ+MzfcLgh
rzmCgVDL1EkqVUs6Z8qJ2cWWy7Q2uJifhEr7hgaRPWmDb/s+PlksXO33v15XWRTcY/0QYXv8DL5p
+bOtM2/JREcQdJg4Eb4Nzhusu5E5rVazrym4SiX8ysbmOP1x+s9qUO5L7XPehnViUP4tfEU6/9d8
Bxgk5vdZQWjMyih/h0rT8ThbSSUW7/ojL03HQDekAel38wlO2l/4SrY5ci3kPyTg7ImytTqRMh7I
7e7IYmPbkDBA9ROHmL5TtcM5bb58Hv7kOYnl5g8HzG+jsv7xX8NAsqCxQBB/UzCSiCISl+q4ZpDg
SEN5Hz7z2LIe/nyqoDkVc9IYicErCLP3748fu76rPWSg26n1LqJJIs2+EiUWRrFjSTCTmoErS6DS
zkYbeyINfVbOaeqyU7nXV5K2Fk7nNaAoNuqGcCSbFKzBTcjG3u6zVPZ+TREKfqLN8WZeEGRN6z78
yRN39vi7CRSjOMIGqPGMe/gzXMRou/TO+GOp+VfreSUVXvDc+B4BWKRgQffHmEkJZ5MnjykSAv9v
gayTviLXjFAhwJB0YF1LieuQ3jhrcaT5IsCLxZABHtq3fmvSqK0QiAetMWBK98cLICFRrGyppO+o
uswrlQ2MxNf+WUtMH8KkN5fSqpSM3boI30FsowNdyk0UJcJmIVIww4cCQyBmGg5kQWxilbKPMgr8
JY7pFG7rz1ZrsY2uKsxLqX9ziML1VsawPcfVBhBT0o4V57PVpfS8avDdjmuPXvgpxGkhx0tbScyp
Kr5rQTl/4dFuQcmpeG3vs5DMjgYlkc0/i4S6fk+W2DItIUTmJYAsfXMTUfcNQHLQysIF138GgfGs
DrcYWnQ6cQQr7+PnD5mzTIqTCO+jAnqPCDuuVIEPWsofge1wmsd4MvENctKkwk8VP6emlIjfR6CU
61sv/6/TJohb73FeC5Yv7dn8MXGlBr5e3kkl6ewPUAKZ1Tr58psG5qXNncquyn2rt81E1U659S7X
S07YEz7h9k64DpluHcHvsbHl9kMDQnj35IjeU2ojmiL/FFSmSOQ6unFtCo/dQui7ppILbhUwJAod
MZBbGq2yfCnCimpnbAYtlJNxnbREpeHaJXHdk66tCi+YX44IAPPDO+XQTcAjDgQq6WrLcJPUo9CB
F2fCLHJ3EDzICa+eCnA0utJ8o20X/zj+gJAzrlqLL66cKVsONepCrF3Vp1UuEEKFUggPN8F5mG/U
OgtfgojnyFPd6oKERc+0FXetybz/Udk9fq2kXZzT5Uwclrbt1QpP9Pk0/p/VpkPj/1BVtjcsDLli
BokB/8N50jyxr6Xe4SSjrCzMOg4vLELNvmP1RKZDk8Kbvvf3lwq4cLuHJCfmS9IFvJifeitrFEPN
eT2t643coF167l5GmyUVwQVkDHrvRuDVkGzxOav/9XAvubEYBRaLUpj5e0lXm9KSwtEO7UMl2f73
vqdaWPJB9cN+RbsyQXpY5maYGEgD69AMK3Yv1cUbbguXkTRtNjyxeatAfEO5Nf2ftvCg76bULjlf
9yD8HpCSlr1Ehqbyu6nO90mUNxGpUCRyd9zlRyTXufdzHC3NSpJtckiMwMlCAHu7hyr+IAUfHHEI
34wNDqW7KAjKZ9OH3r+PCTQB7bspLPPeF8ACIWIG56ZoMB6to0AVWj55zR6WZpYc9MDNV4fEknM3
MTQK4+K918iy+PcTB++DPEvkrqkDaoWZsHV8ZThcrUhVqKSGBc1KZcjYinjO2lzR3NR1owLGDp5n
EovlTESX4FfgABGbxxIYRgkoPQYxVPGCJDE5zBNzHGVH92UpxhuJ4W0AMalw5B24l5IEIF/x86e2
4+nBfp7Ic0JuaiZ3cb9koZ8SYfMGqpBpNUCqPCuPelbk4xTf3SyY4egTG11JYTz/XgR6ecCW18/8
JCP5pIrYb3z6zuaeQ679olLtDYpEhjUIPNoNQdQRBa9mVfrgi3rdf8/Dk3goTVRhxOCWMmVh1oRs
i6xDFWsK494m3vRDWMRx+mh7gu+qD2+2ZL176hIr710eFGQBWhY+IPoPR+M/NCYDrj4shRncTtVC
fr8dlp2YheVCBoa60Qo+FwbIVTw4zkEGpYkcGuGfk2g873JLXBX3bJhWKG2Klgr+AepNjrtWAZPn
VConOEi3HcI2Hs8MtwwYkxoFpZg7SO8ZXysnVtjHA6jIPD3yXQRVYpSj9jXInFDrYGW+v1OmbIxl
fGSgHKLX/cyqBC8ur3J63WCAb86ePsHEPUDbmDJlSGawmTpHh09eWv6pTuaQ8dvQOKcrotATX247
8EJIhzcy7BpfnnvGGFNPNw58Kj/UFPkWivDQNmRQcqKtK/eDzcLlLRBwCAEG0kTrpWgEDC1o5pBM
Wc1j+1MTqgf8pS+IJfG4KK8Pdye2aWkEhuBhGjTEEM2P0pJXPq5BmxjEZZz+DT7RKjHSKoYltARN
YP6xDu1OAED24gX+hLril/3Wqng1gNWFqj5y90pcotKUacUJ7Bolz3k42bFL0TRNKmTheS1JSRSF
lhtnL9RSGznOAw+SJWPzvm/SE9WBBGsnkHw9sYlxriz0bcm5yTZOCsi5QBN8rqVXoLcy6XyBabnU
aKoKXN6RAlYw2M1lSYb8PL54seHMoHssDS+g5NRiLuRwDZy+pH82AuUE5ER5Yvehqrk31BNCVSkn
Mdb92c8MnsiA9NSiWiyB1Lcq1ULYWLEH6RV13j/2hUVMpIqB/mWtywNGYCl5au4zIokqWowdThso
o6tcDpvVDHT4F+G1gmExoxeh+NeS55b0qVIUEqOfNCq8tcHFuVWe/BMNv/6wGxSTECeDWgZ9w3Cy
+uj87cZj58qF4OBQ2IdDbNMqME49Ret++AR6b3rF1d0SLK7zzLs/mgFxB1ZNGGqcPZgbD1kkMHKo
oWT3QZ6rQXXbuacJO19pc0ia93O8QKKxdYAu4QKHVS3IwhEUPvgKU17e0mLfsywWHkD1IjPlj8T/
SOu0iykvUtV3Ct2xem0T8Zo1YzkjWIiLjEwJOTTWBz/4Aw6BUipDfhYhegPqv9B+hQL47vi3keHU
57y5Azjjo2w13SvP+YoJ1ggVNvc0fr3oQ06HYBp12nzWnf642OeWVv6Y9/7xHa3DOwSV2llyMQof
CxdbsD4eTdid1UYFmAAUA26aOO2X9T/2p0SJwp5vqW9swjkjsuU0dOSVJTc3MfAQ7Nm0FNxoaGYZ
o5A7lQZI2XfH4ZYHErs1tFYy2f9Z5r1XPKEs/LeicmrxCA0rnarJESHJou1QpYD2GPjGSScX5VF8
4nl6H3TPxYvhzIEGyqB7qjcnDIS470yGGm7cUqWSM/XnQSNL/LYM/112Qa/YWDfaQbJCw6+FG5Yw
TZfz2KjfFItFs7o1aijOZGHrig0bsUnjOsjj+qcfkjCmHmJyTL6Yh3tRH6NnX9MaH2wKLgi5Xkon
GN7Y+N4nEkVFIpEske7QG8HiWGqJztt4w9X3oV25ZoroZgL7P8E6wMrgDM9mMks4lhBQ+ByMZ1OX
RbQxSqLd3p4YIy2Vp0Om177tjkrBsC5pXckzUrFWwUIUiGUIMKxM7mkjP+wy6gVhAFrtWDKXlxo1
pJDgYxR0KV+osxJLA75OCD7/G3811OrNrnU396xjtD48r5O+6S+WeMi3cVXkpBoa1zZ2IRXF+rLR
uKr7BjrUVLi69x5EICYZrVBrRNKlyHonj1xqtjAZu0DuqpBaSBC6eJmmu6BoP4cu78pF1gMet2KJ
ZFmTkZ7uoeOOhCSdflhd1Oyrkuw0GlmEGDSi0UCdsQgG91bEnwUV0R8GxmqEy449rpKQKh76bB31
onnDuGWumdXoDuRp8/fzXiQofGSw/LsVZayOxeiofUJYQ/m2zeC1K92+/4ilLUTR+Z0ZkX7pCec1
PEmvQjNwsgV5UEum8NyRZbq4YK1yzMwipz/nuhb2YGTQtFx4J1t8X9U2O2QvoJFIdlAcgh4QAXon
ysRDAMqGm5lNscjqZZOhdGhjrgR/Iz/l/9aF/a+0Zx5gpN7kT9ULz6nFfJrlN0QxuRdLSij7cUSK
ifPP18pui3bie1e4uhmDhMpv1dUX3Jo84BZMyaNiOQOpbLIp2vUR0uYvfzjoxkFByOf31OGyNWfL
Aql3pn8sUuMyUnVKVw+fRIHDuXjexaaSHVFAana9YkR1k9YDVOG6XA1VWp5tzPD4qyqveIHNyFty
KqFP/YB4XO/VODJ5IW2nACd1i2YaNZLMSU9h481JGHqYEu0V3lEKO/xKuHvkuCo2OnK6KOQ1xttU
llktZSAo410VNlyWsClZlrJ18H1sqtQd+4jFlW5NDeousY6/m9ihCH/tfTl1Ut8sTK0NJtPVOGXD
RCP7xNhyPUBQ9gUnnF7zm6IoakLmAgw016pG7AoDqcl6Tlf6M7+1RpBKV+fdR2tu5RFXNLjnpST4
k0hmnY5g4oXLreaEzNbnMMmXFlR85PXUfgeSvSVaJ1pKwz4qUNHIuHhPfYcFexzmYGQr+N7AN47v
CQ4IoChdC9N6Z2BqZEQw/RVAVZJPMjFxdNMX0UDnpRtgOWtyQWaGUK1Qfzb4FczjABbG830o/y/a
P2oqkjN0WNe1XUTwO2aBdXOgxgs4iACUDbenhUvjsiSTVAgZb/Ttf5UmBVyHoTAQBQfFG3eFwBfY
uggyiY7StggEjsBEPjvTXGIodggflZ02xTN0EcMtzN6SnwvYD+aOjRvbHZAWlpxMorSuR9BFoVku
Kldy6hTWE0LKIIBd9ho8R52bmsCGFk6l7HR2d+ehI2lsyg5en4bouH4gphXG9+/hEE2agZBmfaG/
YdtWHR8GWKMzaj4d30Xeq55q0aJRb11OXTO1dRFBGTW/eYaz3I1EsgkWnlPtuIkIjSdj9gkkYdS2
GUuKgmQjrqlzlbtAQI8ikgiq0m/8nbYTkDAKGaYUQ6UXLYj6Z3w6pd8nXfvLQ2t7IFzffR43ok2q
LcZfSibGp7DSAlIHh8OPDESc+mUNxO7Shg+081S554E5weAJB/2czW0D30Hy3sKIHtBeQZwvAt44
jn1WSYqboX6Et+nKN2X5KYZm5b/xyrdtGGwAEhWd/w9PKrXd+iyQ7UjEcH/L2cz4YCMohW53uAdw
DGxx/puMyrtrB4gkWWZ3J9ZcNDEjT1FuPU5DgI81dwL4xM6G8eW7upMymue/GTmEBXrhhVjdg8d1
YMowT+fvt3hxqwl53tdyfGnk9dqYNy2v4EOh5eUS7jP5GcIsk7crNpJLkni6o3y1avLDChVL9Ahs
NZHJ1W+VlS1KcSxjKwCfelP1N9fZesOVefhHeZP7vow8sq6cDttZlSsrSwUDgdG02Rz2hRVRUnkB
9wbI016QZNiRHhumZW5lje0ZzXWRyTPZyskj090sIgJqLiV0W4euMi5QXXXtTE8yDXLljX3yCVMu
VO/jsHRH9HMSoqIgpbZ4+0TUrsd2lSMHjpPrREDHst7jSqZm6fw3NT2kFKnfmXHk3E0BchWe0Ie6
C+U3dUTuZ9Ele7VkSkVSf9M164g8GzEWqTWl8EC6hRaa3fnk3DVZDWgKNUdfbukwWD4Ay6hq1LSs
RXEWU+b6bkfKDgy4DpqK+ji0m0SStYmxKZ06aJ0YSzJuDaMsmVGJYmpCA3/2Lvh6SPoMQJ6kHYYF
aA/3otHGtsGd9NOx4IOH651ihREMzwcSxbK7h5hJT3SqFHW1RDVvjhk5LIfiom3T/WycPlKWYkO+
kdyWHW2kK2Cw6Zvm92XxwW/wBLdZCZS7jwc8gfxbPj3LyCmhZCHDSKp6BhoAph4b4ciFlgRd/p85
TAdi5ElVqm0lohtwlG9702oMQdZHqjR+FkkPkdzgt+B3+wrHyBcapE6V442kkrzx5LIAQE4crqEe
lVhJQywfrLz8dOXaMifU/7ZfA/axKZjX6J24E2/O7PHu7Eew21r05cBCE8tJG8ihW/7yrHaImpsF
dLG9DC1+xFo/7FT5eKjbEoYwD3aYXkzP41IyIhE0W7dm9TTQ7IjkI0Anq3UfxwANacpVSogycqM5
Edhi+YToBoc3uqkJMfinqE98KLhX4FtHD3Ob0iLn3gcrAXecJo5jsLbu6JcguaA5k8W3c6K/mOEj
jYj8TLgasq4DFvxwaXhRV+CEFkJ7ZArgMjrKIIPx5//OITrFQN5QA9NYBsTR1t158syWBlMlgCqO
j+KDhh7mN39MDvg9sj98JPZyPSDPwBr9N3QX106HKyPgSEN7JG0O5LuUzHHNRoh+ekAFRDalTks0
9ebRfBPaO1ZMMaQ4GRHCOyMEQ+lhRi6u4BCoC9UzujVmhByR3rOh0Adl9OvPx+T4tx2Nb2h5WSqT
6jbrbb4v86qRkG3QaJSiJv6Fx6kgMQvXxPuX98zk4NgNiwL1oQFjljTQu/O7ukn6qjT+OUi2Vc4+
viXQul9qP2sarZJBjqdMPCvSG4tOcSDzMBc0F2dJoQZkYks2U7wa0nIvOPtJhPm03FWwP+tNuoXs
notD8kT7kSadcIV897TIHs6V9Kmg0zNi1iyjZt2BbnZXyYq2TIcMCtwhBwUAq5qNXALtQNGI7IvZ
PVzuXd8mNk36zxamF4puVqICYZUWMmiasknCWpNXA7QFRg9Ehl7iXNGcV/3Dsjk0dAC0Hrj3Xt1a
f8NIAnhYh9X/sY4Bp5t4mxnpG8dZavGG4WGO36KCBKHKmDpwVzxVw/OQbcQY6d71leI5CNrUchWu
h+bs+2vvG2I13gJ3DtzIEcl3bXhGthtN6qQKHJjU0844YA5WJnGZWHvoI/G3qWj+DErUurfDLH3z
l7kCndOo4wC6mOJLTVTrqeOL8BX735JNV1qx7fdHMxjxI4+87AG9ub1EXS+V6T2R+FMcne+SKNh1
tI60+vHBDHKBwyrJuHUy0wtyFACxuuocIGfOWh+a5JbAB9/rsi9+M/JM0/gso0tj2dLnsg6EyNG2
23dYSbkJGJtWHO5zznxYHzaCLhVKi1IfYjoEJwuL+MWbObLtcBih9G5hmwbQsTIoMAB2AjteHudb
6bUeZyRUe7ixiKyAr0Prl+kbGjwiDK85py406XAe7iPvhZ3sdgy360GJtjHlf4IjlhVQMNfEV/Hr
tz+TuRoyJ+1R8Vf/u+l62eOdgVaGUx48zU6mgOPOjo52hsPyI/wUTMRJd7bZrw7mAdV7WHbrxWmh
huXLmByTmHiYprpDZmffcbs/jFm9vDuvdpvtmH0fYk5TFGNrcIAHPZKzi3ZaaaDbNeQR5Hnjl4lU
zsNCzSmPY0oUJ3LnbzsCtyoEa3WvVg8LWWrCvZVp92i1zOaQjAuxzfBRJ+ZPtbjV7iHvMumV71tG
zi4mQWL6PSId2I4MJFg3s9FVNOjQGSPYq/Mcjoxp0qbF7Wmo309UCU6O0pUd3w8aX3Fig7ALIvYL
3aX/UmtCWz+JP+kRpJGnpfAsVLb0mQ2BI3jkJIMHuE5Ycs3xAfpMeEeCIMprU5+7KyiU9pOMCxNS
nT+CAYiVYoTxo3ao1EbDcyu/sVhD3NkIhBdsqFNhyuHU9GeBJbjzX9StmuyWjT1nBKLne53x/rGr
D+EvuNK/tr2K4HxYgZ45b9OCof4qB3eN44YzlOL/Zur0k+bnST6z7E0z35ZqlqhtetjXSAGq0ZP6
ZRBT7EJkprdYobFZan4ytZyNziwiVJCFbe35dm/F8dxvybjEahtqZzTL7pAx54V42z8WCtTxR6cn
ayDKQP0N4bw7OBAc2mDb1SkmBqccGYPoIbG34domV1LYY2a+kWgYBBfSsYCHUS5TAiDsilorzET7
ReEUXQojzMF0PrB2cdQ46ZEfI9Is0ERbcNAoa/a/hkUwGA8HQROaODjTpsUZzrzattOr4IxQWdV0
UOeGnnCFLbw6Tq+o5NjtjfY95ubLRGCQkS2SdVtXtYeMetspbGSSOLJeBVk4SAg96zmRWe/hr593
i+PCEfTWraMBAY+S94ekZLnZJJM5dII0CwrDFYz7J7cZGw+64d9c7qGWk7lYfBcSL1MvZ3zWiYMu
f2f8jUDEkKgVUt89J+byV3yPeN2LVic/U6XGbJH5AyU5OqLBjf/Dcw12W0nr3TDBWgY5qH70crCM
SS56L1kytW2h3vFaS6BM9v2h2KwZ5XfTaqbfDd7pS8kSlHsCZmNCCoBeFrWFDxf3zk7XJKhOPa9s
Xm276Y2Mz1PkZyWb5lPii4ABPatnwOp0bU1qRwQ+S2VAVexiptZ76wLoAlxaHb3Ep0a9wUwV+7cI
FBRDYD4wnY8R0OkpaPkqKlpKUblzsAAi7k6g6oeJVvJQlaawlJyVoVYo6sGODu0KKJxj6aAh2lfg
LJiArQJQrATrdG/xZqx/+yNihrWB+OenspayFU7/VZPgMbn63R2kbHPiS/4cuspiksX80cdrQcdL
cGUC3Dl4ivmU38nNKsaMJ6u7HwkcipHyuf6VgumZ9opQ7wVuLxDT9h82wSm30ekyHQc25TlM+1mS
6+SvfaMwqxuUWajNb8ZHb/643i3X2TDdrYHPbqGwla280wRqRSOKleMCmLA1T0kkb/0TDVLyqyVH
7TpCazoR+tkOzyINAe7pt3l+Qh1BpSAdfeea3WLkqbDmhsRkNUH5HEtrZU48boj3JszZj3Olf9z2
uhuCOoFyxVOn2w68xJtv64ZKurwmET30PqEHeTiR/su5jLt6r19iqCBEZteUsBCMnWO1loDwmuAj
WlpYdQHVGfXtllBcj4TOm9+uP4ElWLptzjyY3v3RJYiDxFQMeMAFcaVFiPLtlYhgKcO40PtoR5j1
nIXsxYp5CEMicZFkPZ4e+O9ouqXur10mMcScER/0JJzk9iKAWiQoCj1C5pqwfqTNv/quTLl2kLw9
FIofkjtVFCP+EF9zfA9AIiG5PTj+AYkYfTe2dGtSlufxom+SwKEgbdYcJW3D8AyGxU3zyuq/wG1o
pyTppJpNaIGsYmS5LwHXaQKul8LTgMxAuA9negd2sKmd6OG5eigIbh/wZyHAmfI2FQvjb8j8vkZK
TgaD+0hFaX31mkjZZ4/G6TCL/fktUYFrDpFZadsM6ERmnE2TauKupjqOcDosOOrZcThsisl+ub1n
3m5Bd1yE+tze8mJhZpi8ziPg9mw+hjh6pGpcNXwtEpuTJExxfItP4vYCsaHeK57IwZbdaesjwv1S
Bge+NxaM033MORSNZcscaPTASVPjXqIP51SeV03F+yqilsHEx+Ca1ZV1HDIL+V3QMZnLyGaji+dj
z1Zj998euWMBG5BzlJiA6NOjf6qNk9uGpvNcJTXrSXDkq/hLulhY5C8gwKGUwLysnLxIKHkW5qAL
I34/ikt0h7j0oT2dyZcOWbnBgn4VEindskhoMNiwzd0x3JKgNK9lPLggBfmQEIzYgf3i5FkFmbV0
+yAtI4jeRBtZ1+yotVuQ+d3tFx8PoTtt/sCcMKC3z57hMP9Amrm3n0nZPxRGnBZQcJHPuZvnrpGu
sl1SLexLEhgbaYIKk5zgk1teKcqa0n4cjKIEWte5V30NL7kixIdHMDmGPrY/74xqQ8CENCML9J21
mhXOsX3tAuZ5iT7agMKy/3QZCFpVn4SS195KkngJs0JvnVczXu31XgyLod9VlwP0HZ9wuWt/4M/v
anicrimf/ORb9mcR4IjwvfEU4BYXHEnJpP2hDy8Rq2S2U6tSF1c6Lsa4IUPTxc5+8mTyyzsf3NJd
HuTqbuwjqS2H70Qv15Xh8C7tzdtn+o5zg8gRPD0pwGxPD95y42TjrACHJeqrU3jjtWV+zW32WRGJ
JoLtlxvgkxohyD+a8OH2St+NlEsMKu/85f2zwZHXU17oZ/QIgEU7dFvjI8/Y9Vf872qEri5+VENo
s401PQdPigEIJ0fo2q5t10dZ3mQl4bti9yes3EwqTZq/g3eQNez48vz7vsLZ67qx7uObcGULJLTB
/Z8WD71KCMqnD3qpoodmpgeDfoX/PBGXPj0FmqokOvQGO2VGUmVKNr3C3bZu2mk3S0o1tj7GyZ9G
dJiqNSN9nHAaRXiENu/KKMG6Rgx78LFXORsr8jCrce4C0hQKnqKX6KDLnbHKK4QB07qGnAin2z3d
qwNAsFf0H19ISURMzScev6IxL0gI0xdoejRDtwtPZ+WD1l7rad4Ssz/jI534e7qPPjELhhCo316R
IgmfcKDBNUwwCQD4Vuq/q98+vF10zzyXcR/vxP30LEfuprhWvlWkcN+7dWKp++uyEQ2HLEwzNEzR
9FknP+lpXZpjCrbAVGfilfCILrdbv61x1qINK+VrinXuF7clnNC/7mdWIO5DrMtlR3l2KC3klziF
N9lUcFzAcxLAF2O0KwgtsNVNsAo4ZaZD4f/mv7Btd5YU5JzJeAcS34S2fJiw8gDTJb199MJYqczq
qN+Ten7IeXrjw+XC/Z4+QTrP4pgx7hf5gWgZw/26qb5KnBaS2SG2SWdMkfLbXIUH4pUOxV+rYfcE
OaNV87ttm6O480tyyzEq+DWx8eCdbXhozPxn5M+RFSbYf/eRQb8MqimAR7YSJg6QYwuDfz0Yl8Ck
HQUBZyNEDEAR0wn4c8cWHZ4QZFSSpohm6eATc8RxqFrpRZNJatzewJWFWaYRXpitquNKLaKEYfmk
VjcqnkxaMuwrQJ1Ymvf6Y5F59TYgxM3pNYtJcXs1AiSdktqyFk7GLdR2KVviJ3qyuVEUQAQbMr0h
n7uCjGf7a5EEWm4dZ+DM12e/DWS9eE556DiGFv135NTyiOx3OjXC9lt14oth4E1/G9Xa9UNCtn4X
MGhDEXCgcKrOg0z5m0YkjvOtCRfnmLvzjzsOaykRvYccBar9xTQi8usv2srDXAoHNMu7Ixi+qRyH
PWIOO2DvJrqqnTrlXZwi5hBrO5pw3u1GNZjL2kXHQ5HwOjPIs9o2KISAMACASuYMvJa1GVK0ElSP
QqbrnHk8XzLa+izkFEFTebKZ2QutrC2IgZculjZ2UgYzluZSivmCuDJzwS9KaNYpaDdtxXEHRVlN
4+r7KuE58DXtnvl9zGuC6ro/dlmgbmBcNNqi2jrgtzEnDKbcboOrUjR2U2r3ejfaE8ewKBC750G3
MbZQLHm6Il+LMyIwacCpjrwrBt75arRIW6EFlR0Xu+Cp4YTfO1E+2oDKiNDhZQDZbSwThFWAQ0rg
Le+VfeWhDyka1HuvABbBGPrAgNzTaGCg6i2+M0OqxbptpfCLrFb9IPRt2d6WVaMGOWY6sgFUi4Z1
UULfCDtF9wcWhjbk1hJPWgnMzyEHluc+u1WqGkgzkHqC/o3HYoIYfqU/u8nsztvkOrp2ZBgEu25O
8Z27kxz4ivSa0CyUdU2mFvDk30w9xxhyKGFx+ghyibMR3sSaZNGRzPLceoCnHe8LwzbOC3DOu/2G
UNM3Qi/OthvCy32mMNsnNXEtfMVR4oBTmpOZcmp+tLb4WVHxQVmk8VdeuIfzTJdp8uSIUvaDaSOU
M1egtGp1IFUwgvlSRtN0YWoim9phAzutxSgmYk2743jilhEGrpyzvmwpg8M8fgeFOEhphajoWLlQ
kkqtvOmryTwCqowwYzYxB3JC8zu4qwUwd+bgzxu02PCd15sc50Iinf43BdsLOg+nOwNbJ56NOFZH
9GcCBztjJr9YvGGDgeSF9itSL0iQjS8/VvPuHXIxraptONHh80rqno5un1tI8aEs7V5J6clkfBud
4Y1f7jpCKeuC6O3bBwnjDohZMkMTOEoGgf2vtbfhAHCte6eRw2LYz9zNkBf6lH5BUuoiU95hmIgr
w763Tjw7fEcweqbKFzpNbv2eN/BTpviBsXkbIPVPgu2QFEqtWf5Keerwr84OndztUZ22ColA0quO
d9W/0ucxGuU5B203i+3XM+skItlUBBRTydnWpKki8tCcNmL1l2mDPdnKs+O6T7ViJjrGBG/QqrAK
s7NVJlqOIPfWnyGoyanwdiEiUvDUx8mCYjNTSBcnUc4fmcXVWD5iAu0YYa1o3CVGu/G7XXXBaPn7
V5dHtVaGHWhOFUfByFpNMzsarUyfAVdvnS29iNiZC2pCl7srIvrzDr399JKfW+X+eicxQVqWNsk8
fTVMHbO0tv5ODu4EsunTfbh1wMHQzRUD5D4ySSbYY6p4n8fAkUrTAkiY//w9C7AQ5qALPxRZM/c+
S11qjfHQULxu144OJ/UDq4NrkuIaPCH0iOuBvm1j3RbglfG9yFkOMoblp7A7mVBHPgMH6svabx9R
iIrWnP2UxGvp2MZO0EGRDg/pIzXBGxTLXTFYVPc+yPl3zSn1q7oWfDeuLXbFMKEw46Ot43isg5kk
3+/AcJFHvgpe1qSIjXQp5ygEzpr5QgfsiromrU2tCs2ydZj2A+8f76aDU+uFMXakiPgWagrbN9NZ
MGSmAYkGPqppov2AWMjxcAr9aH6dgANxVDNGW7Xm1AYrSjZq9i7YKIVgIKAuU7I4FaO2KU/uj7sr
05hj3gi8EK5x+uX+YgcT0tbo4WdBfRFOx1e/547zuCPZsV8Lq4qc6K3Acnov/DYvLk9jayXW6FFb
EYldhqDPdzxdEZeRyp8Zvi5icuxiSgsLRVzEiq6rrtb2vy0k2fkT2HKvjJ9rtdruif8pUY7mio1a
86yGm+vLcFgoyFGUuw83Bw55dTWqxsF6lFq40ZWEzc7S8AuLTi1nUInA1ieh7myG0L1UxKRUGiI1
fpMxpMR1W686bHwh9C8cWIAzoHrbIicqSBIo/sI+n6tP1XuTrdFAehqaisxs0vbq+omExlD7HS1I
MEP9+4QpzuMcevG+aIl0srhdqEdT/DYIJJKSNxXPDgUJAOesl4G3nve8kgPEk7h8vMRhVYm6tvJw
6hBtkEbZqoh3c4HkA2rcwBraHIWnxej+/pIQjKu/fv4/JnauP/+Vf/+in05igDwIwCKHq3YqBmNW
QM7EL59hmjhUZe6OAjBoMLJG7qj4pftmxQwGTs5FMsAXsS9nORhD9G78NdbS5bcCPjRvTmqGPpG2
ouWW0eyAWlV5BeNY8WSOLsb08OGmThqY4gKh2vdRhnUHL4LStUKwalFa6ejB1Hja6Sy22I6Gj/Ss
MTKWXriRsBTcW2c8xapaQIaoV8jV2LY9N3xImqCIIFOSeAa+kPb1bcxzqDMraNtN5wfHKJ6dNKkn
KYbE2UWAxpQuM7wxGst87Gha4DpZGOhqEPisZjJ2EjLNT+cdhCyh4qJ60iSyKofAUnFfsoekIFzn
sGKoLdHNBHIuj/eEfa2kjzic6/lczdmY8gEjyppKTb3VRQRotvWEM/JxBxn3skq5NF4I0A49mJjI
mCFOlutEP3yTXqTWPiku9NHOJrbjMqkxnRCd8Al6YkUr0h9sirWy7DNTyDL5nS5GE/x5nZrtv5A8
cook3Vg3I2QQ4+CJ7NPIkMKiOWqN2vNPQ6l/D3Ut1UVbbSkR9lpr7LPbZuI0gOHGW4xzwvEFF8Y5
kIIY1VZuDGmabTqVlVZIgqtfZCX1uQbGHanGuBDOTpaczfH+SUnd7q+TarEt9/qGuZ2pk0pelwNt
i3zzxJa2aUnAP2FTQo5zWcTQPa33K8A0zreDatOAgyKkqvMI1kcR0g0ISNidpFQMDEGezGvSxqCP
cyQCCIhxgMdeiH3cwsw1AhBtl8tCJwz1G/PJtX+08XfOq0heSCP8QcJtwgJQ1SOPVXzrSi79KtY/
cfHIMwZEvLoHDKlTOpbGtFDwaTwpCw0UTcxoF5UEktoJlyD5mLpehpXCr1SpzgaoEBMoiEZsuV4E
8RJ7NNFEQB1xqcGb35+WFJFmSfA+MVSVCbdP2n6QtHxoXVbkt4QQH+u0BQ3d3CC2C9mtD72vJmyf
VBUv41AhnVM6IuL6Pra7ax3nfyc2XN9xDVxt88wpWmRuDdhVvGdcyiBUlGTKXREr/iaiNEqm10bj
jg9UnNXqldEFzXSvU8w8hmpbEKuUhHM4O5sM2kAlyb0qt4sMnYwi8lGXSkVIK6zTIQcXTsdiOWLz
pZop8Lbaeo5U0VTzb0eVy/MR5d+FtI3eRYnBcfS0BVXthZ0c5c6FRe5FR/8y4oKszluDJ5fKsZJE
KSLD/Pv4Vke4Im0DXcCAc2q1hg3lHXH2lz2sRaNTG0uSYbCfwwuSGRhZxjWPomwCceTK28TpJkN9
thI91/U4ln49deZk4XU3vJqWRkWp6WG2mbAZXXENO0UDpiS4O/rx4SDbjocLpfyGcN9bHa8nP0iz
IDwOc241dnK3r7VF5y2OQ0o/yb0MBYgJEu9w/1K7z9bhqreMLsy5TgMU3vCoRQKtEvYG05eUXDZg
DBvMgV70JPy1IGkFtq141Z3Or1GkHgu0t+VElsiyfkqg3nh/4rcl6bdsve7L0+237ReNRGJEM/i8
QoEgedTIqtUblVyC6Ha0dimuJo+9SJIpcKfyFZin92GwLVTf2tdxtPJqnw7403oEcJcpEA6sX4pX
/C83ySbCo6b6cviwWHsNz42GFGTFH0YmS+YtUN8l93vMtm9dfWr4T6zJRV58vS9baWmuBFhSfGNp
M+N3f5rsr7e3Z9xbAGySNwKIzfnE3uNKFWP8lSmUEvymOjdUDCAd5pf5fSgTuu8r3ICWWZEOzQ1l
nhvVOiWmm4GPi6dKTtW5d0zqqK8vqxSFjMQZ5Jfw7MJZVMtJsp5mqCC8T0mNFTaQ0cXYOBzDdSPd
47RVqc7O+GY4XkFClCs4McMh0iYzlTrnttnqxzYAFk1WRBwV8hFkpoJit0EhJujOVysRE4UcFgMf
6grvsweC7E/yEpORxyiABtt8NGvhD9zVkT0jWqRrBsu5RUJm4F0YKgHCKbtGMQ4BjeEbeb1YCpv1
a5egvB/IJbMxYINJhBpMd11AckaKxsAumzkIRgNCJZdtAM27m/kdlHZOlbz4quUpj6huDZT3os9V
5PmPIZzJB6AoTk2cv594h2PYZOuwxzbES4rGdorfXMmak/bjd1xsUss5HdeKNGPeKgfXGZWTwAfM
EFMluQRFCQujgMjBBshogBPhSGra1s7QTsuH72LpzEN/GwQEFURbK9gvrDwuREVtjrywAm92kGbQ
HLZcfxPQwX0bxqmdyLEA5AmflYmkG5YWMxY6OteEy/kzZEJC5rA14W7/wQ5i8GGOB/8czHlPoxE1
rlfD2v576IoLFeowpRNUxBTZ7Bo2XE4NWzMFGWNtGQZHbYub68vmNsCIxLMgDi28wwqmRj/X4sOJ
PflZORKcoK27VayE+I1Ud2S/J/orPz855O/YTqAGDA9gBGh6pJpQXw20d0ujyp7npA+VWtc8cX6y
7VgDcX+BxmCFfgSRs9MMncuzhti89K0WhS+nu4xeg2G1G0qDHeWlu1z9/lmfheQBKDj+zsQcTiZi
AGOQForWCjNLKJC1Pw7hMWMnvpFGg5mM3PBDxRXGAUF9JcQTHQZSO9rCmB/RC2PWxuPIeXZrMV2m
iLKR1OXcp0xUEbLkxROO1wnm3aBY7nhT7R76wcRX2mgL0ECJhKJLZbGU6iQ+QIWcnfNs/Ohb3/OU
DSNLnxybI0m3Z6M8MwXnQev6SO7pmX3+N9KNvEaxG8hL/BAb9SU8HwjL0G/YFqJe46H+skR8yqnH
uEOb0DRssAMvvKmfkdFkR1OZkgyCeFTkSpsIdfFVpOplJvX6QRSyBMihY/YejsrlFAQYc2iRPu+A
FH+DPdZDMsQonxQmfhWnoENrbKMcKfe/wG4EB7HWvXx/XYnxmmAgdZhpKo3a8vTuev7OsHwwYdar
ScI0t1x/YS2oKJoznEYD8lk5O0nwQ3Cqp01RsZNOjI04xcpjH9s787TiJRub8HTtMsCOzLfz4Mwa
THZoFR1Rw5SzdzOUuWd4J1KEpSnudFtxGXnDA7I7vrZ1Z2g78adgpubtIB43DLNq/tUmB6dXk8UC
TgskNgNr2K4woE4fHhuaIAbeCvlm3C891hn8e+fWGlFDOr0Irpw2vzeVVbkh8P8HovrwP//w0wVQ
TNVVMI+uz7tl6SayWEXy66wwTP+B6KsguUzPzjg7o/xnLcePLrPjwS1/Btiz8ELyvLJ0GZ1boBGX
LKhR5B9vRrerW4T6XxtohRv2vuMlWX6fqFu1klG2l5Wveo8bztvJiCLNx5mnIRPa8oB/6mI0q6Ss
iJmqqDIkusJ0bBLqEZmYBKP3U1guibfjL1gsf5aLUxTDHIEJmEDAJYDbOumF4TM2SLj8xu/Xto71
jTOcrRQyC5lgQEP9X+cHLQUvWz1iWdGrR0q0M7hJPH6RwI74Y2vjRt03cMcizyISw9YRJ0cY+smw
T4vEHM0ZkT6rw2a0AE/pFIA3561KEKENAGqewUGvgNUB1GmFjDPmUMZR1735eBWlaRhdeQWqRwqf
7W4qISIcw93Z056FvOlxorGCOUnHFuk3aEqgOD3Qp16Qp1BPCkaexw87iaDEBN+rliTtbwvNOKX6
YxgHlBb/efG5bilaoviodLhmcmreD4kXuS/w3T2Kz/BwSN6hCTp1afAeU8Agg9BzMSQO4w3YAWuY
I42EmQ0kXyD1yOqWnL3S7D4tS3OcEyDM6c3vfJlPRWI64i7T+rnOsYosrPcagaFCaLqYsqOlK9oH
2m5/cQ6axamX++6kcvI3mHlq3zZF0aHpIayIn96m3wLx7yrptCbENFFTBR/WeKXNPDudDpSrmW0+
Ke/b9s2U8XuyTYG36XgvEa9f/uEwUvc3X1tYDcH9IFO+/3Yqlb0tgd4ICNjLhIM4/x96QZNTOXvp
0SUbKIXS7GVo8rSJ6f9G12HErBvQ0RRkPvxLgZF+oJi5L044eiskZ+b2Jnl7aBPu4Mz1kvmmjn3u
IChW6noFc5oFEfegLbPLtOntZZlIAg9GejeUpruXJktgd0iqmdEIHAuOWokiG/BmZPeyuIOHPZZW
2rJe6vFT4J52fVmZWZ+7RylG90MtQ+IBycIn2j/XhbOy6EfkSs2Rjqbwq42waH8sDyVok4+mBET/
si+Xbmoc8xp8Xt6GSgul00KqTUX+Y21y5O5e3qC+WGc9ua8+thoMmQH7qSDHIH/AYgHsAnUtgMMi
Cu0jZyzDVY5jtN8rSSXpduVdoqkAaUePBHVJhNpge6LXTrnX0SWYQOdkni4fvpieVJbR7KvgmOLy
t35pqCGM9MvOlHYzVfvrVAZoZK7g38kIcRCz4XPJtLfgomGtDiLGAshWK9IqU/AQM8dtXHx2YCWs
wsDqAJZ9ScUrlwS1bj0TUBQy+PB8SUykzx/jfFWhV8v1oqTYQlO+HUwP5wYWpIcPF3P6pZlWA5m7
VAA18EfHoa0VbXtqk/n5Q3cFUHjscrG7c5XYvy6x63z6ICXHe+OXhUHtE3JQy6WYMsj2WigpsJHf
PsUNSFYXKd7ovDBLdxM21/izQZfRkVkmy0+zAxl48liKYImP4DDMqP1pNer6RXE6M2P5SdpcTFpf
xRQ5/BXHVK64u+5AgN5QnOY3cBFDBC3u5VsuB7PFtNI9pRBPnMwPSHrfGQTNMpqFiD2ash+ZociE
aZ+t4e/7eRRH5hwGF3IUgwx2x5rTU/5PaPBIKQY+DCvyf+HNvkwRc/bU2spk8x7+/DjEgXWJSaeB
KLTZzjPhgZ3fN+rly4luvops0vHZXMnW2yEutlqGzx1KgZOyAmvnRtKpHWnW1YxSddG9eCY4Kqw7
yMLqqeit6F++DU8S1vPXWvK/A5s6OlHGsBOsM6E67VdXh/mcDtulpGwSQHyfwMvrI1qTbnq4P4MZ
ERMx+TuBBb1X30s4eDdWArk7kAMRAoA/U2PV/hQJ1BthkwyfbpfSjomCVfnGdd2pKs7crHN+h6Hh
BeNyT74Gb4IFoNYU+3FKAB+BUK23+roOkjfm7PGp7ZeEKkddoKzXIvtbLryyZOa7xaDKcz+72hBV
qXeWwsIMl++kjVw6TJPGn+Tqni+4rJUTsAJKLn4LeoKSkNVHus+3+pIdgODjLi0JRm04GOudlLH+
yToiWWYh5Z2EadNzkOZCXf44Vwk6PuB83/WedE6kY2IGFgNe7fEF12atxm3zQmg79WOcwV2aYkrz
D3J6qeWGkFpGZuPxwiqOLlUoN4Onkf0DxbSeZ4JmaWZAxKLcLfNWVA1oKKEP2hRSaihLPIDLWsw2
kppgXQt1O1NV6+32o/gqB0E24zFLqzj4ihielEUjr6FdAdj4X3KKv26w2dui/ilEJfOxtbk2Q++u
bJ4D3qLp2KnqPwtJKiPioLkmD93MmMP7X1JxnhyihbUwSzX07YrhLym8JDacEk9VZMGAoDFZK4qP
doo39ekR3LH1LwIF+MfvmpOlKp5B5lUODy4sD2EI8jxz754Ei1Md/QqolBVL+0jMnNT7uugrmRmI
5l2/F5XFzfybYlGrSq5V0Nh+j1+tGNRUVLPN37RTcwZfMJqHTLCYAn/YtojOZS274WO/IvdnaVhL
wtXPexiQ5kvWkeyRtHHK626OgWILTCxxzsOQTaPL8uIBop4G/xO1s1zawe5XED2JlSfJAnL7UPyV
VUnllgMm9xtin6nN89QfotNIPR/leBxGel0dVT3U0ea935Y+X6XKNjOfUDVVD74Ain9+tZ/xPrMG
FvZrwFGKHGebvrxhXLLJt1CE7Q3iVsTye2lKClpL1R3DTktP0JPkY5eW0R3qRIUXsnpaZyJwep9o
gnivtbMM75dO39nd40TFelXowfiqqbtRi8CkM0kawEzA/nb06lFzAWbfmRdy/QJzWUkOo0u4mFQ2
hOlzKJ7VWujomkrl8706aOjJpJnr2mExGCFh/cp08oXqfsRl00QV899NzR0fYMd5TCNXOXBVNXE7
MwbzbSu0QXG5j7FtYzoFbb2b2FWsaDJvb254gD/i0CLs0H9qqFuq82C1OrAxaZcDNa2NiYKKmu9G
XDrE+VDIJhTvg84x9EhVFMY8M9DHWMQBQ6rHXNEWjhyhlvmxs5tsW2mm7COR62tY2JQ1L3o5lJIE
63IUDnGfolTOBMOv1kYocQu4OeotvrXfyX+M+gcYKMg1JwUt4xjmFsSjhCp1DOE17MmGLa8ErJWp
1wK8rVXBDgYtqwxJfGEZA2l0bl4QMorRKrldGvrirRBABXgSQDtsdx86z0EfwFWO9vlPPhECuAQF
8maZvBgwAf5aYDGFMUJP0i1YBAwAqBwipEVPUJcY12IlArpX6pEf+Jihik7W9327pFaHRLrPwGPu
PdNaphNVNXpVqSNOcMln1eUpSDP4ZAImHlYOcUnI+4DOAuqQunCr7L+Gk1hTL0DSeOvjJNFHEMQ1
Gb0pgESUrOnMLckR3ZEU2c3pG2D1OS9hxnOXNOaKEF0Tt2LBkvoeinyohhkWpCI4UfSQZQdATzGf
1ePjl6wauMmJGjDBlQXMaZXQnSQlqWFIIEkM0hQ5XwUJw3MzNhezt5NbKDu5g5Is/NCLxVFoEZb/
ono2qorXaN3FDO9FUheLAbd5JAMehnZrD2C53JsL0pZgExBAnRNI8Q5YkApGtf+oWiPy6GC8Bm67
p5sjQlTKemQUwJkbCzmfWe5/St4qJnWfaOfPP7fvuis4thtUclnQMBg/uoxgxiTqih3S277+xpbU
xqRlnU16Gz6x1qM6ZhMinmYDoE5Dnuj2xca3bk2J4aQ3MJio4txXxgL2Ik+TuMRDLSUFec7eoSbd
3ZpLAa4rM0bRI42VjTrYhl1JgZIuIOOK6/khCy5CrMw/T6+dMgZw82566D6GiXHtYNqY1oTTafZ9
8IqMAEotcPzA0C2rkqIxbFxMjmVj4CGRGooVVH53GBrjStITGjn017uU06SVBD+ZadzMlPIWVwHA
L+/VuVdLf3tfxJtukIeDNLUwslRTU0nmJG6wSaq041PhIy+3yBtUoSrtx5TN432Dzs/2R0us2Jgi
HYNP3BMp1Gz1YWeAc9aSXZtbhV2mXw0L87mPEg71Rl13OhVQ6SyDENmHjTPLHuCwL/7nAVS5vIUh
qTRI3i6LJepKPN4zZzfErSFi46y2KIfDSErBEbJ8UIeyW+I9Ge5s2XqQQRUFwR8ggIN8gL7TxwsP
Q1JTF0m18LgB7X4ML5qvbmPeBFGTrVZ9/G58UuJ6S7D/dalTlOWStchHCd15hkrvUA0BaPmgn132
j/OlwgCT76TZEEJU2RnqR8qeu9PVrLCni5J7Ocm9ExCKz4kgxrEbgomyh09zFaZil+h976Z6YJ6T
TUXFXkhbK7ueRI9Wfr5xUvrB0Cm+Mm/wXVoaamqQt4Sn66PfY0cQQ+F7ofQ3rWGcoshQbwzKbGYE
R5LOgdhjmYazu1x1/Lj8tj6FKQ8+lnSGoQ8SHV52zHM24RrzR2n2GoG3MJ5STit5sErGTnN4PfmO
U7RcTqi6VqZ296g9cnvlRTTJJrB0iurkhfMO3DtHHMWpPm2huU2tHtVVTLFBq6v94wsjTFPrPZAZ
dLjJc2WT2yY1uUNyPVuvt5w8S8chN6rqIEfP7unNoS6chzi2dAdMlE6nELLIzkp1Dzn7EHNnaRbC
+Q4kwKcEULNB+d1o2dyrCJdiPVBAD3sIaHZV3bwqbL8G4RzglDw7sLXq4HvvCVbh5+v1GnTBtone
GCtGnw63c7VAhNLpi5oF7SAvGqGIMzyNBx3G+v01CLH/NvucJjovnbyMNO7KWSbuWNnYhVjqfXD9
EJLLvX5FACtMJauYVaeUXSfjvHquGV6L7mIrYiqzjdNa8d2HNOLjM+CYhU4AGUgUnZ1pWusmqjvp
QHFJkRavRzSmTPxDohfscWM+9Ex9zcNV2S8zaHP9uW2ev3TemKv8rxnT98+7U8Q2+AwZ3DW8M0C3
y7OJpLoRuT0+6UIeAcuICuUOpd3EZSgATManV6khBy9wUaOe8TGWTbIgwRr/OiitPRsthd7rVRVL
P1H0+C1sGtY5Xn8FWAIh69sEmyfjHLcu4X2+yqtJ7tzmTQhGLwh7MOGkrZaCkCaghqIU1UU2mpLc
7eA6K2cSnelNBqiUJoucy3SOk34YsQ0llIMqPYMllUh6/MZf1/LdFaseM/Hfi+me8jpBDlEGkd7+
Plgj9m911GvL3isJmdiH4V2G2VdGsvOL3pneBq4BsHKC7v5me7V6tIWhlWwSKAdcg3ZIchspzYQM
GGPvqrLANrAiG+iU+IrzATiCPqznvkHILNbANQFV7psxpMWsBYih1ggmzysX9apfGn7I4jDukr1M
8Q//cfji6vGkJl6/QK/ivvhiVvNEUdbF/jR1zeU+DBzx/vBK0OhInj6oEAaKMSHSSDJXQLZm3fv8
FrTpaOj5Xbp/8p9fzKXUQoUaIVgj7Y0FUortHcLVoqFut8lMWzJvSU0JRN8+5desofi1caPSd4y1
eNyLkvD2uC+EmsrP4SgX+S4noLTWwXfywALHvZplQzRjMZZTtw8YLj1QdjTXhsVWpwzbVLOTxGkz
9vck+L3ytJvLxjKSlyab4G0TjmMm2DwHIG1HAJ+rO/8choRCr0IxLPSbxdOlhGR0gen07WnaIiUj
4AJdbJ3AQ4AnTLLgl0fH8tlRDE8LNt9g+xlBfi3bBHxMiREu2WaeeqQj4Btl5jMvGkxSLCwUxA3y
T0ABmCl9AsqQVtgM2jQjf9p6KJScM+lUW5gd+T8IB61Wyhs9mqAk3Np45qkvYsvasaIYKyYqfUZj
jQON38GDa2xu+0Xxwl6k1cjBWbCFsyHjSefVnj8Igp45xuvfBgQ3A6QC0BEkRRX7rVYwe2E5IUk8
YnrGE0hFMbNkhatmZXmQ+KFs51WDOn73D6VYrtHZ6k1WPT9dR/m7KRLf4wA9Y+TCjylpc3oBHWcO
iszck2Tk7e2Ij1n8AKD1k6/rc1P+Zib7CFZCBc0rSuHVTgpDHYbY+8Rc7BaQDiSujMXS34KYhakG
ZhhJj6izuYBNGPOsHQFbWitjtXCRu9Jk6jKEMiUGRjX4cT5/U1hjFOnRKYnQgKYZIXL1wJwEtUd8
mXmWuGWfP2dlztwloRa5jrXMe4IV8cxp+VGIZYBU88nrX72HUPJsSNfXKkCo4/ftW1CgBVCz5Ban
KopXT4ptlGr2raTP4iHvK4Em/82Uy/yJfvvfJSsGV0uGmuTje1mN4ebYwp7zJX8D5u5OyRN+gS0m
9MiDePdRq/8CrGg67Hle6fUQaEDqpF4eKpwZSlxL3jr+sdZ7fxJDXs/AeWOA+MIb1N5np+wo7qit
ZoDtwhSjjCPTM0MBxjGgToME4FmJ8ZMAFyRf16nQHBIwhL7IJ5MZwSJbuL6rwgjqXKH8a4LFbl2b
DIvH9e3UttvitczdZmE+WDbwExRF8etgue+BWzvp04XWcoXTmYlKRGxic4yCsxZqyqs+sayNwf5D
p8rggFz7WsQmeatKF9fS0CSlH4OFqgFIpJtOUfUxbbNcKrKttkRx8GFbyK1Zn2fxZ9nd7/CqXjyM
eNWd+gSjlPRqcxfez9fjzakIkw6RCFGyyr2Z8mtPjOQ860Fb/FeVTaWqQLssYCRwoxYRZJx1blNc
wM6daczkpR562E3y8zEY13mjp5nAdwnfNZOZXXw5DlDR1n2OUrVuFZ73CMYJoH8HuII6PnkhCK2m
2CgoxYq8M+hZichdL5d1Dme6OTMcZfh1Sa6YePeVGBN+vHEeZWxF+MR/cHkTYbjBIBNT9Fclg3wX
wkdxN6BYLJG7Fjt8C88X1p9I3+GMvekt83/GxDuM6fZLesBYD8jxAsO9ER2DqNcyPVP0RjXpt3J9
sHrfssgAl4LufOmtIvW4PfKNkTMnGfJZ9MjGphP7pe0wVHFB3Hu06CBvCrD8m8a1BU6+wx7uYr/m
JLdLODQMPw6ogz/LYhtJSesLKnwMCGhTmPWdIF7Zf0ebPcqMvecUCK6Ve8BXJgtzCVnwiqTQEsG2
aiv2RPCVFX+9pxiU6vtPPqK+zh+iJVpH7Fc7LyeOvlaRk1SC6xRk2u4eyY0+pqZ0a5QOBx1zJcG1
8iJwBBU2wURcAZspjbpQEGnHrXzstc+mhXBc+dft3AbEz7UimPcpZX62BxEJ8MOA9g/aCd/7uqHH
WrZe6jieguLUm7QwF4LiCgDwAikZoOZAdT3b8DjysAkWg5pgDmYc3XTrjW9bgtl2CML7bwNmORQX
Ro6nh5o6vfUGtaoi2AHgHqkq/GIVpe0wLDbCOB/CXzjJ6f/A9eN6S153T12MtqBU/jUlPyR+rsV3
9FAGVdIK9yJugltaQh1QzhX/DmzHDnOqi2HdHuTf/MoIapsWEOZIcK2cBZybWXDxkiawM5WiKCSY
p5zzaSaYg9t7xCNeXMORd2Hp5/vWXiiE0jG6bJKKRSdqrywuhNzGdr3Vo1f8lDlR6ldPWES7fViR
K/8V7WlYUhw1qurvWUEmD5GhEE9UpGpjs3CP2m4Q2rlLV+1hhV5WBsf1VRtVbRkD9jAS/pCYmOIk
Rj7E0w8Yc1vg90S2XAl1PWpD8368RZTWfJFbjKf9gynNw/tLL1NO2GNuZ5zqjl91SeszVPJVmtuw
wGPnJB2lpuom8FJ0jN47POMwzkX2ud+oDXiP8MaMRY+T9nIHZeSPawnjUR4RnmqMmQW/sfG0E8PA
rR+s2seZ8G7KN6zbZr7Z9B5nlHIa9k6rSI8vZVhxLgjlQ7d0wJb4C5jhXp5YRovOXGP1jnQgh5nS
i+vxYXBMnds47iCOX6GzvXexL/b5Wjmfr1pTYXqzfRKvEKFzqd4N+ED0J3AvPvrdw6yv9xwTfN/M
6dHG09/MZ4pIWikr+MbMTeqXdShrgh8Bc8k6a+kwJ90t9FWtABOkxQ7VIgZefjpd17z9lEtx68te
OFEaeeuUMEz8DHLwvaW0jGPvIMKP+HdhVPrejGMW35YV8X6Xvkj2rwGxFZMtzVqB4VyJKhqkfCLv
r7/KFGNJuJvXLwUs8fVSrdiIQ3asdzFSQ5rGE83Fs27bBn2veHjCcEKGvXhwabPssOShmvUZLCSH
9CbyO/uQOeWH8XC8S3OWiELgppcgBzAIK8Shj6WBpGZzNO3x7VlaVXzOL6GQk3xwq//c9QZS5oXx
LpLc/eL5gEUpB9OgAcmpuukOM0olYY+tSLtsKSqesJVrg67uKLSxA618+/Zq7oWd53M/cUeBG2sJ
+jtvnpuPl9NYHmgktFNrC/uWjKuZCUocVWYqpKHdPkK3bmCL3T2S/NaZXMRSuM+Plq6oO2JikEAb
x/Y7ChXLoEFZEI3mCqTaG9SQXMaq3H8tDBV4kx1ipYbIJc26xo2Z+LN4egdeuzqtRAaxe4cx2A9y
49z8yHPDWxwp8P9gytjoPE9dsuRTgPyAE6+dmVdJXMwV6XQpYaR/LdKAs9jj3MzCsUVQwF86Jkgv
Iy4OutSf83LXrIod7M77HORHlkEZ0a21NGt9o+gscC0d7UbaNf9jh9Kwcj+ERkPqai67KYMHuim1
C7076qSw0vXs8Sgo4m9G0Yfws8LFi1QaiqnROW5iGDodClX9bpXfKI7KQLA77Q9AKvqRfUVlbX1b
zGbxgfhovJWLTqMv6CDxjUJ2ttveDSTti5WangE4CCedyQTGTNTulri/ss4F1f67aE4C6x6uXGO1
Oqn1/nkZtCFS6r6rgL1W6QB7a/bJVB/tDvcCCiYwlpDei11BDU+heoVrb2oF+vW6aMiNpX/wS00n
JXLdGxj1ih1MrXghS0r5M87MkxFad6JntWB/NaKR2JZSBkdgNVIO2h7gvTJAPGbPixffX5PtHG99
ZuejE/RFk+Sa1xvbVC6iX4gzMMJnKKtgBncyTXxKhpSQu4Tubw0fBsPm0yz1fIlH/9wDNwgt5c/E
V5mPgGPLkc0wPJ6KkEuSW2doXKJETuWSBLPv9GUp2R3xkpQ9WkyDN/78st48WUJxG6FoPKrE1gef
PLUrskQql41Sooy2P910CHtLk350uxaTcuO2OXsVYOkTt/Uebda9Y5PVoZWx93cGdwEBnktpe756
ln9vi4vMRbrrn3J+9J9BdVmzBp85vykf444L+oHyIL/uLKFueSm2hBhLF+UHG1p26KC00xcpWQfA
hO5M74asss6rnOv121Hs9Ik1vVONCnMqM42eV+cZROj4VpicBxJnKUbPQC8KKmGLH8gFfGM9K6so
Y1/37HIAmqY/sRiRsqqM9jxeYvus7sH5+cIlUZ3QR/7GXaJYplbBWQSlcpX0OoKNKG4STU3P8BMj
edgDrxYq06Isw/ezyuThJIGXK8gSK2r73xMx6pt3VxnGyKenDXTq7pLLoqfPanfDEYBTX6IK75wk
wRgvNB9oycFh2Vkb/I3o34/dgmT2oP7GrLxlK/JYlFl45DTCD2jBDJL4KBYU41U6jxbRzJuWMyqt
nv1mz3GskRk/OYuag79DseWOIprnInszZFCTzQ30rMYZ9kwbJ4YqLfvxfTJJ0foJqdh3joxaAtWJ
Auyl/k3tsErvjSoNkWLQ/3RbviNWdYmPSnQbo9aWQx+HyWVx9B6Vb61MjRXj4NY4PwVyVUH2p32G
aj8F4YiHc9xYahbH8JZKB2lGrkaxxqG3XgRu49Uy0ZQUIvA2E7zpX4PtaB6vLoNfllSALhmzyp/d
NnspVpl8rmPj2s1AKjcaQ7iq+jYwYUL+jN2yFyfVj89Fmn3EyMMbT2EeCc+PK/7Zxr6grMslOoAU
+6QRQ0F9lLmuz/ecJG36oVsLxuEqsAKPr2aiBsaBsdkJZXAaqUwCDocFh4hX0EhXucQAIle6Clgt
SZLg3Sva36mVxhtZfGVDE2NYIYJx1LZtCRki0+E74R1xLYYRaDY5upqEvZZ+0ZtG46h9u/DAsL0G
ROpizUiKFJQDAJitYQ4ak+H5AMG42WKhPOyXZu2hov4SwkK+aWkA01eCp5i0ZA6TOZ25c/HpueWS
CLg5fRfiucbKfyD2rkJR3KvWox9EdH9WvK0TwwVneoMxIeTXfWf1Vc1A1rfR6zPXMRCGrmZlqJk7
WAFnuvNti60S3iMHX/mcOO0IE6d2fY/dtBvXTz91fuv9EM7YVXOXAi1HpKy/dHxhuEcpOrklU/V+
cErgI2oUH7mIONH7AFumDBC956oFHh7V8XsSjxc8IXaqriaeHC34RKC9IjSP5+gITfQ6ihT0qz5L
EV+DnydvwQTM4Rn4UQAVQIsCm+pTYyZ3k0xn54uM+bnb1GlPr5dSKd+mUK2BVEgrf51Qr+OIoGLY
9oBfmh4hysqStSeb9wEzoJBrskMYO+nEBnznr5tdW8XO1Zes7L2ldYWQBdPV0HHENx3e49mN5Lub
CJ5h08l4/l8oHENUGNKpvWwdt6d51N68UNonVEe0EtiQrLHC5VdxXJ0TdLE1dsHDZZMv6FX9c1qw
b6VUlgE3w1MsBysddd+yWuMrAyyeG1n8cuahJ0CbuvI2dmuP4Sz82Y9XCp8mHKbtBeZ/Qm+kpjQO
rl4Tw4gSA5Au7nuFZdnLtDD3IpdmCBkt0UcmycKq9AFqKmN4+yfOFXSvubwZh4KP/Sfiqc1uKJxe
voR3u+3LkrJeHZDXIhvXIwg1FooxtVOaS7VT3esBeL6EP2aJzko5W9wY/yj0mS5m4/bFrQCNaIX8
u93xBmqPqNlvp/9ek0S0+AF75BurXnsOfjf3J/898qX126xVLk0KaCBfj6TcjAuX54Gw3vkYCfPO
9zq65tz18Ch79Ex7bOWYZdXkt9G0apwJM6VBDu6ZuJGP5E7iooG37g+oYN05LLnNJxUJgV1mAJ9k
bUnurklQQQFXPpLzohOTO4qtbCLIuUDRiFQH9pAsKHnFNat1DdXJtNuq+0ofXnx8QB7KtyLNC7KM
7wPCOZY/j2J2QQbTrAfbttqs8RpYn8+AwIHhKEjcR3xXDBgVN65OvnCEHrmwKv/yXsAbdk/p9tyH
uJPWKOJx0CYosA7IbWbtQbdjJuDjr9KzdBMZZWQMcCb9MF38LNnR+oRljXBELsDqjGenpyZOKZRv
rEp/gcqJXyQgQgCDOo5j9292oq9qR8DQiWb558W4cdTENwYXBMl3E7zOikayBP2Q8LLoLU+cdD2k
HGGGdbjWZZeJ6hG+wcojDy7EgP010jLeIcAaA9GleaZLPrzSyK189BNnHT+5PRnAo7al/A8kW6a1
XxDoJxhaPIntCnzZFWuxXoF265KUUIagQbQI9+GXh6UYxZ7ZnISfVptEz/xfXDmMgydVAvy47VbY
1AMMTjlZt2OPRH8gJdSsr3qr5LvSCw2n4yGjGhgqS1SlM4pTG7mvzET07VG+RG0FJ1n49I3JsfXg
+Pu08UJ2lOxS9zyNPFqloQAqxNHsvqY6oXYD5DJzBm2StHx+wk6UPhVYkC3fpP/mIiXKzUHRNXK5
W82zr5/uZx1a/LQBFrSjIBW8mzkzczLH+lZ33OfawE30aDhMtyuYK+qeNZK5Yh/4wA/UmrVabR5X
DGO4o3z7si3Sij9fEjYcRqtl66N2iCqVVUK05yaerefXNcLUw3pIX5hKFVzYffZdyPQwcK1uIEmO
FX4OkNZs1G8RtMtZRQzXJDx8fr0OWVx1JDyMtO0xYyOVTfDJAgNTihnJmL6Auy5AfpD8S23tf1DQ
HVl6LQe/5M3lQRKtH4YcOIQtwPZgH/gJirOqB9HnHLvYl6dPKPiAJR5y+rB8k+IPzV94lbrlgn4N
K1O74YXCGcWQVLCIA7sAJe5f6Y8UL8Padb3lHJR/jXYoVMoHcREKPPm3bWpxiu9nPkZJHshW7l/Z
2LbkrqLZgDKKXuUcpFBNXv6C9WHJ9YC2w/Cid3DGFjzT6Fbn0I6BEc8kStMHJoirutFtDRzE+BWn
YFDvyS2LDNBtTeneaxyPUgnKuFJjK5o4EQhRLb2p00bsNe3NAgHd8u1uDQiURALV/XfDcys14XNP
xttu0W0WrGv3hcC13EtzEUaws0ZSBOhGp84PkDKf35QMjtlgECrBZBH772ZQSl6ggpKlCg/XN9Yp
KBMUjPp2vJd1Fc/rwYUv2UYouDYaFkz0ABrRGxWuidH1533lapCFNfeZvQE1arB/ZhcKllxfoXwx
oT2GLA1m/hLu5LjO/mHitDyejIkWFnPNerKjIs6Q/+AaABpi0POIrb8bjDcWZKf6n1Bb+eej1FUU
eN0ERKkhJgk2A6vDFy7lLdM3i4QsTTROuE5+Fx5h1uzUa0zlyRYCxEE5EUDQnzx+wH7kj6MnGbAV
uW0LlHQ2cErq7VGV8ZqkDq25TYMWzVhjBbGtbh+MRGz2XWDcxjTacJMzrPlNfqr1FPJzSy4YfEbj
WS155smspeF5om1dFSmLuqrc2xZ43QxKqWs+sZcSUx1dzZJ03H6iZJ7so8yWTE0WZGL93c8Nh+Rg
TMBzh3+0Cfb172T9cjK96HTsYs37fiUbWeGr6/xJa5LqZMrZLdQ2A0JtXa02ayoHaVqmH16IT4XZ
UGnm3BmyTOhDxcMaJJ41vTPtbippgA3WOXKodxltSz/+VMc7MYHftavD5fCHInCJHJaVcwojIngy
llxpSY2Qtb97yhqFoSMrSP2dSO0vdHZi1jrTWpRMniDaCS7tkENHCUwXYrO7+uF+p0MsqMI61BuB
/0YrRj6va5LnUwDeQxyxzlF/0umgnDCaRDm5JKdVgM1BZk/UUKoNi53DGNHFaMP5B1iv1ub4J0Re
IZLLZDzUsxzh6p0FEP+jiTTXMnrJdsLZbwh2Dg+1MD2ZD335f+cDzBmzAwUiIM93GrMdcQbt+cit
kXGBw6G9gCdi06xdFxWNvWIFPa6FJIjqb5AzF8KFg7KOVosPL0uZFQLcck9afsdA9M7UmYBBjKxg
hOqzJaEy1C7Zbiv80AbNE/Ro2/RJikx2CUFZ3NdQJDEEjON7UG+sP22xfqAwkFGlzq/2gZ2BlSLk
eoBJtir/mYsAKUyleU0Kh8/bcadn9KUdN/dl11Bv5oqigOo5I5ISqjBmqrfpIFBCE3FctxCFy8s1
5q58ZKY5R7Yk0x1X0SELXQyiypaZOrnBGfLAh6CAQZcr6+wqNBgw+vPp1GFkqdGUB2Gai0hvn+ZD
lIZzb/x4Lp5MeRi7y6DvH+yUD2ZZQ7h3M/GdBmuIqFzOmVFFRcLIXj/8FWRobCNQEhsaGbbvlG9q
w02g0wEO3YBKJJFryDGMTJYfuokOMgriiHByjKhqFalfYfgc3Ou+d6Vms+0wO2ucFJjhC9H+TVB/
C3fbgalWpcLagsjdiZD4H6z8GrW27Z647Zi4/RMEAiykLdH/VAofKD0OzjDQ3/+t3PlIDR7N4FC9
5ojSw/rcLAP/58qJYnXPWMDzXEfktOFalIG7rPl8CJCt2gjjgJMnn/P4OPeaBqd45G+laLs82Let
cCifW/NAcOcISOxlOy4ndF8WDM8yd83zIl69utJVdQ0pYV+PlZ5JsmRO3aEF8rDTn1IwYO2DhvTX
Zvku/m1HieByCFwiM2V6RaTzQ29FKUnNWccApSPkozjTT4wOstHtvvH2GK1jTqFqmOjW/I4T7Lr1
khS94gu/zXf7R8d3RJRhCn6wO1sX+dyN7s0/xwAtywFetp7bpqt47FdlR7kBjXfl16vpessNoGez
cRLZv8XOycRdlWbcQ8pj22WZR+cyGYAd4Wg8sSY2yxX66nnhty7W2mM11FBhKSslaXow1ipQwDI6
0n4I4xhtHa2gkbNssPFCK+koGr/mV/pWPK9seCj0hn9eyFDHaT75eY3YJjPutKQbdYT89bykF4VJ
kcayfTPQx2RYrPNroX+5WaQAbw2HZYSh8JIVsdlRnmsCIqQIJ8mC/Qh8QEOfRpiqbttxcWcoeSeP
FcD16izgtQdnHvbqRaoM9OLXC4u1NxmAjriKxefr6VZtEZ/Etgz9E4yCXYpw/nlStxBGFnEQbRKW
jWNYoPgSRUdAIo1BivA9oqhQEPM2WLp4BuW6lJRdZH/rb8Dm/BDU841TEw/n+flYHdjKcj1dALjN
IJpZzz7tM9y7yK26HB1ey6dSH4VTq01Rrkm6q0w8ZEVrY79RZgS5eYUV0UaNQ5Bj7X/UJ5/lynb1
ECGnopSbSrVqA1Q7c+J9bo3SKNc1IJ5dJfz50kC0V1GyaTrQUgxg5ZBFjvORssLeB8owAURHYcft
yv8j41T/M87Hkrjzm4z1U4zOX0TdtLXUDUUDFmgx6oAhhIEZAT7KeHdUmGprdeNbzZZqgnWh1+Va
82KTfGATZs1PNqWBnW+sjjzSWOFOXded8ylUNwYivy/9MQ0Hk3B6ZVHE7h5L627Q2dxDD1LtJaOz
tYmhusZ6cZS2cI4yPyJE3XdHX3GdjAAG75ZkKwCSVja2TsrV4MECD4VU4XaXnyj5tHxXKde2yT6d
EEFWdwl4x+3lSLc6GuICIRsXib5GrO1FS9iK7QEOgpLDy2XCZkYfv6sl2Le0HFBE7EzTu1y5n5d7
VCvBro+YsWYTdXLFwWr2PwD3nxeNVXz6B0NKqqc4XNukr9d4Oe1XAvzqvNcF8cxE8bY4VoqTTpZy
q9j+NwOs53g0vBruJmfeeJHhyV3XCSCExYgegrlSdI7Kx4hK4VWRJ8Ip2K81GUGmjCCMlZqw50fD
5wMgsQgAWI0IFBivIScOeLp8zpsYP29KfSb7F+bTGUThC9/Tlw1DjzK/7XE5hoL83zOamQ4ucoZR
TZ5+IZBYQl0PAde2qfYwc1b/kRPLVEeclePCCu1yEY1zayGNPndEZrW4om5vhO1XtUcepH6DrZEn
4DZOE1X2z0Stpm2yMlH1jsCcQD4VX/1OkAn7Fl2VG/kN/3djXuFKG7PDOipiZzA3DcFOxZf1KLWb
qNQvDZrHYEv1xrKrfvN+ExbzK36PzghUy1mvoxkrI8/HfJrKz+vzg4kYDi75/nuLhdJTcPMwSbJd
4G7b6wpeXpqh+ywNiiruEssB9xZhNP7gg7wEDbVwaTu4f41TEjv98Whw/xjh7UV60b9Q2m3htYCB
bHN5r3OZevbKoVCTOSdgRyD+Rwtl9/ItzUeINOsaDTW5XWgdSk+PFYq28QdT7Y1lZcRxs6dvp+xI
JjpAzkzrWelFduV8r9XOTfxV8sFo7a9cepXMNQnEnspZai5jhuAvayEZH0L4rPuUQTUDgoy/1nce
AyAEy5bmFSPphR0XuIyMVCu0xw0X//LlKcU4yQ9FvnHwzZQbQdOjsPoIEBTmTKQDUPDjQOoqVCfE
BZr7oXOF3hAqlM66QK7/NT1b2RXpNU1BHo8kyKuhzN8SWFkxyhV9c/RJmqSLU1dGcF+r9jS8/ZvN
U3YWZpYTHYrw5bgU1/5Py+VgdW88cFwxgTJYO1JKeNVidaKqZd5r+CX1HYpRtAARTrD/8VD5r9Bt
cNlPuLPKYv3ThyENINzDfeHRBftWzuy/vTgJqOGHHZp8L5LDwzKXBTg879ApLH34vPdbCxjfXJhR
agvuj1iIWYF27inZ3psf/cQCiR+UFiZS2RZMw0Z5jwkkzUY0U+qeCbxEyiN9+AWflOVZ3878Jk4d
/maz75RyqQAFuvYQLGqoITsnxQHSg+D9+NFGsBQeFUaYyvwupj+pMiS7+D28aaZXLmTsJ9FW4Elm
6inItjLN2OUKYun9CGaxI0ivqKFuDhBOzJt0wpYwxoqiAoMM/4208BtOD2IWSSBkeN7NTAEA0wDY
qAIO0pjrGdhRn+amM/+HcRdyxJusjih/SMvuIGaeEm3x+SoBALCZhIqRLz/FYVAdohWfwm2RcBEg
7dKDkaUcKSZ9Qj0ydWmZrOqJIJ4qnPW4dUFt622RC85x86mHiigAoRDNbitVr+svyrcHm3CB0wzO
zSvCTVufOW8qSjHAKxQZD31PqhLHr0WvA9MHbLg/o2eqKLr7bGfxsLIJ8ccN3SzEnNyJS7AC4PzG
0mNfKZnbRAjJSm08UTArEjBhP8l+aKrGFDAnTmH2pbH6CBUpc5Aftvni4FYFoLeQEfW0fGTZ58lk
csztQwZr9LzpbTQ4x+b+yprr8reuFcsHgLUuQ2/+gyOqBmbs+twC3d3ijb6Wim+TE9GHeREq2waG
LnO8Lc5MoZE68n+w0WnYLDSVpyJSwvFUjFklChDcv/FBcchVfVaW65nyfhAp8y4ZTq9SnpRLEu8s
A5Vf53YK9GQB9T3lyZEZNbzVjEggi6lKjSR5oajT6jQqmqnOFJXXxyOz9JKuqg4syoOt4wkGz03G
KPElmtCs+N6yyWZDNTmKendMX9HaIBhus6CdNL3zEUCGAJvZHo2PAsR0yjxY2O4U1WXmbGn+3/6Z
0DWK1Oylkl9xnqFBdvi1jxv+DP0+010xCjS5I/C5Ga5IFhpl7h9ZYQpiikj2YSpJm5jouOUCUnbV
XTCXrWd2qSkZs8irA3sxtp92jrIHuxTM8ZYP+WvbRHQJCQE1LfyLZVG25McvEYLB3MJnDgz69QGp
QPuQZn2vXe7Y4+bFJ6x38zC3Gp2zko4ll5aNScAmGBTLWNWoGQcx38y7pmO3lgiivweK2VCvlLGa
wEnBWZ+WfhlVCc6vQQWEGoMgx90+Yg0fuDh94oxGuHNlsv25vjpXRBvkGprztYEbPMUAPu7veMMx
n1L2z3HPVLgZ9eIkxbzDaLy+JtkFkQsBzpAT46SerNCAQeP236flzfpPt7XlP/dwffHE4xAteOTK
bBThdLTbBxQHl1aIzjkK2sh3+a8st1o/c/JJTWXlXgQDXpxZMZGkQ01xL38ABP0Ekwby0GqBc+0x
xY50TK/KMFHabLa3Aikh+a0w59LxDJhsIKmnjtDlBmwaB05uNJY9hfYB5EAsWT3NYC80TRIc+eEn
pO7jvJc40/3wpzjrhtSvlG4Dm7zZHpzqs7n3zetmHQB7h++sbcTyjvydFQDJUhPuyq/I+4b33NhD
4XdJknBG49yRWvjRoUq7+XpZ/ev7jE9EkdH+bcW1evixCRDB442NzwZbWEpbvL49OQRS5fwGyhx4
rECBNjxEigXUlTHX47MxK3k3vQ9yH3Trq5Re6shOByoSJkxNZUBkIRwzgj6eEPb1ELbc1sAF5aGD
5t7vv0fQdrd/381SLUTHIbVfLPtp8xwpaO2p09sChdWPKaEJIePaZXSF6HD3bBpwyPuxxITo45cd
XXrHcuts/Xd25g/t1jmRS7+Es6K/TGCS+SaJ+M5pNVQ+PU4UMaFqOrt9IRHo6RDDy11tnGCpaBsO
paXdaSVT3yluJ5ax/xC/CrSaK+uy5tUAXPr9UasKHSADRmo7ixSBNPU51Wl4ruiUeyEz9+6W89sj
jFDjbFl15RByNXXWjjPWLyKUmY9uvQV1/5b/udo3iC9aQMoGAmCEC/Hl35iK+FYbxH8MCMuduXac
lYYRa1sUBaDJAWtu0f7X6ubz0ucyk7MCxokV7pIVYq/blTtXuKv99Du8Q0cYULuUrEi8dPCc48SG
7a8ZbSCc3y4GLa1t/PZDg7ErZfxy/ezvQTaL64UQupWOEGejq+puHdjVO02hgYhkGRvOnIcMYu/N
Dezjsui3geHC3Zumv6YLx3xGBJnSswkbHdIJVxDMacWILCZ4zXlLOh/rrWdHC8x6RZhx/82d3etK
FWZoLKTzecXt8NUSgIHulHwxG520HUgVtE54ZA6zZOw0wZkdqFzuedTMMysAyPBRfqkTcSURD/iI
nuOm+eCnVzGawLk2X0AMkxwadrT2DG2cId/WwYmz+3MNkP/JBwvw22UCqvWJmMjEVA0Ynt3qrsqm
KHQ7LJoeK3Z/0JRN+UrshNlWEIEdMWvim0uoMSoarkTBIsmFz/VyVsMc8HCm8IQWCg2pzRZ7gYrJ
7bv5SDvSnh7v3GUdM7XmJ8/PTzf5fb/cFEkUM/mKqEcOFhmfg5fsSpd+bunUKXEoJvWU/oKBXSxw
PP5BfG9WDzJHbkVaP7gUvWvLpqzmaMZzBF5f8K/wELlsQ2PiIHjgf1peCmAp2j5YvmBTn+jk5LpD
nOcQvwpV2DodNgQ3Ka8W9j7KqufAA6nr8sU4Awb/Pze4JUWMvJ91Xk1sxzjh2m+50oEWmARHs2gW
IyLfU+DTX39QZvctwy+ZsK0ZPUjGpuWKxacDUkgu4FxbGa7eDjtUR07cmO8Y8kPh+FY3UjpAVu85
kf4BfKuhnY8kp++F65MJObYQdRAoymjqUma5n7OlCQoRSJLsMXMmHfkvHYyRj2ZDQxfMtackApuB
CWYFr94K5JpVdXSFL5Y9NNPichRChYItdulOxiuJ+uLv40Ms1T6fozrX9M6d47Y4+Q726TG2FBTr
lTFuEK1OTLhzshrJZzUwb17msgBA/CHLmKDP4YESf2/MF9NRzMzZwc5wg88u/Cubyf2BgfM7LKzH
+nHCoc/h5j0g2LaT46NtEO83MXDxPr3k2NSk1rZpmnWFyACUGxFXXgsWJvR8kVphk8I0OC6Ul/ah
HX9l0JTwTfHRHwEznO8AAbSkoprFdYEYROGeA2HoahOdUjh15ULUVlI4nLW+ujVLXsk4SMIlgee5
BrQ4bO4CPgMqcUa0hBUwy3jAEhMMOufCZZYA+6blfULXnZ5si+NAzW1vyJxPfdmF/ec28l26c7yA
KAwf60f78wrGGiK0LUAXRway2HUUO+6qqnx2XzJFkcV3H3U8L02VpQAnneC5Cv9yDo7WwCuhdyXm
oRY0f7vnXa68LnwRJgw8wKTO+GD1NS5Cs+kO71MS8tuF9sPKmi9eqTEoq+DNfMjzBb2WjvUJ3VyZ
lQlGKCQCCMSok4TNHtuVvPVNMOimC5YAp758Kog0OOsax5gpRzXTJbwalz8mYoAvJTzNBZTAfmWv
5aBn7vx7da9pv/xiMhn7RAbqdJFx0Q20B++E8I7+nFrXjJOOb+RGkVHSicLZql0rDAPapF/L0gO5
NpyLXNm9jTkL3+F26RDaQ1zLmQSPK4wduTFY2O0ad/iBvZOrzbrRE39cOnNQJiCl57Mx/6G68/Aa
bhwuj917l7rn9pJojLKvlmKzXstUxlrUARvxZMYxrguuGGxjg2Oj4y9NLxrv+H2YjZ+0cZnopxux
GnRfZtwBIFJQgdPfQecpkMbTfJKm0M/lWTyEG7/dP+rd9AZY/bOCs6hjrjfRWsoWUmhXCdEMEW3v
RTdE5wda/SvMyKjvNzMj8u9H4Hkss1lK4Ysgw6mQtgaOVNt1ulV8AOMZQh/rb6QXHr5JJ0KtmiSB
56gJh9fajTYzdyAmZc4fvYAyJEW7cQg/O3rYyO8XgWYyoKFl4webeDfwzz3uwrlN0bFNtKTohhGy
tY7bS5FIvhdmucHe4j2RbquLrYO0Pv05rjrJ1w1DUiLv+70p/DNcfA+PysNj4E7RRLEAOljsfJVZ
pHp2R4boWMfiVzJoNrXYJap2bIIWzNi/uZGBAgSOlYbdNtnnQZ8wMm+2LCsNZvZT5LzrlXqIjUNu
SYnzGp5nWSLqHhZARgcb8DVOZ5B739sJ59qAtQbwGIY+igwU3eDU5g9A4VpgorOIzOztxaalGqYv
tKIkWnj6+a/k/ctmfrSI5YeFA/JrriliT86q9TPWXXst6iBI2tQY5SfU4SXCindqy79mMkBGhesU
pgzr0X/Sax+01Lkrp1UU85aJxZuUxVb5Y7W+7BMrelHr37qir/iPNs0GUglN+BHhtlLyw6WRrcvn
DQVZvZGrVjgAZkHey/yTS4TJC5UGyNUiaMKug171svrHHI6Vj1LM0Oa1OsbTC3pPYc367SrRhxGU
j1JFyFQzUfXsOnO+Z2pJTb1nwWWArF4rT49t24XYOcHsByVNzRz4zQ+uyqxjbW8Axlu0OSceX0aD
ZWywSJd4NG9pYpoGqvy6auy9Gz0ZSvQD9BMN3aT8R+GUnWE6P/vZFsQpkVbCRq3VySQEViH4yVX4
wBXcipF85uBwOic/BSrIDM9vR5f2Wb9lNdnMYVSZQjJIDCX2j1NTGjQxEBT3dCXxn3dgeEz/bw+8
6RqQEuluVYIh3wyRY/Lwdb6jQ9bKQNH5x4KYBYyf1Hx8tYpe4Qw2svL4XEy3s3lKJjvFEBSbBFus
wmkSdjcvTOPDj8/Wx9J7FgzZ8nje9iWJ61NF0YmWWfUkeTcUNugFNifz5XKJ0NF3smk36N5UPMLO
L1DR2uBcXY8/3dgm/iIhZNX4oRh8YXu9HEZUGM7qbO2ZLxG3AqRC87kWMijpK+Nx0ZLOWaLOv19b
io44h9HOLTgi/Lr1pNoy5bmEjri/YzlKqjya9hr024048BbRwMUo2Bg0JbYf1/gZOFRwQLjgqwHx
zMywfx8ilrsDia9gMQEApGZZmpaQmljGxvXO4lw6TLy5oOk6AXppu2oni2zje9Zfhk6qlcv/BtvW
oGIVsrE4+XJ39T8ZVJxGHvE2/rAG/SCQcGfbe2oRz/iRIefK3OeegXd8piLnqaxfuLZccpq5DZCi
K7IXlpVsmzs/hnBUog7Mw3QQTbpZe8190qqz7I+t8dfH7pM6PLRHHrvUPDBJQcof5jKQuSd01KVU
8nkbJ1uciGx1rWshBUQen+iL7OxfK7KJGQmu6nKLEP1gIW+mRva2Z1Uhlcm9ZZwml/Nde0L+qPWk
0ImrVZrIKrYPzwWP+0k9+inw9jZID9rNPgT6WJV3WKAcUrFeyWY+6S3imnb9WhMn7h3/tjboadum
yFLHuyrdTM28+ZQB010y3016u8l9LhdXVhNihBDkHxt5hdPXRrVgDFs8uttiCJqc4HBLaDTES2Fx
u5dA1NaMdjX8sMiBDjVzhOlMRLQuXL2yoIlJSFSepF9sm+1wItL3YxXZdSlbZ9Yy/oDp+PiRgcR0
6Ua2mLS2hxran6eOEtEeVg7pVbAoohAdzrZKkjOht0pMSRKqdNE01f+jLW/YOI2vAZaXunuuqf3h
phSjN7nSq4k8fblU5mPdG93O6N4tiZMHe5KFOdy/pgbjJwV+m6y/YOy3DQ8VMj8w3JaQTyJ8bORO
Ca7xwhQEW2ZQ1byeTCNk+o1C48ot3CD8FByy0wSlviFgxyeliSsVyK1DyTpU/8CvzK7Efntrh5iZ
kY7W/4y9TuKhRFDrv0SHLLxm05EDZeBq0CjADR0iSezAl2pE4mvsHhkQQ+Hy0hM1IkpreJnM811j
hhzIuGKTLtltkqvxyOBXNu+KeNGyIv8/CafI/WPuFJFzPasqfpERGPHFXE3O56DC/zT1id/S9bD4
thOKJudNQEWA+O7Qu6uhe+RMPMdVoW6i8q2c9Z49wmFCxcTLLf8/mhpe6hKV5TQPGa+A+5k1+qGg
hK5TsguF+dn6jB/syZC3jfJZnALmkc5PzlqGizbl6qOVo2ytIwnXrG8l5365oKIZol5e9O3HWsJJ
K3lG5ntkfp1E+CrcmBR67aTLfKxWJT+Bnn2ytYVClSLat89X23lqBjs0hw2mtI2lGZoCBniH6rGK
aeyY/ttrf4PkK9gwp6VhgGVpEpoSxCx5+8M56xGLLQiJICLZhi1yRsqsDZsNljolQaErt7dEkkKM
rp344ss/YLCcj2/nZ39OD5vH7DDtAMq3V2Alhmgn5SqtWiin3kVNaJ5RfiQjvBs2EUkMevD1QAlv
kVul1CswRMgAAx4XjVsM4yqM/JUybRQ69iWq6R6jTKsvC4QMculRAmzE2ngcWu/gVFL8KhvyX5in
Q7rNSaHr5kjAhICC8GND9OKJgG/5VruwHsGrCSpJzZXVs1phj+w2GawKOdATOkT6d42QsDmyH+Pe
SaXusxnUuOhyiT7Wxy+gNvDnYDvv1mw3Qc8TI9NhlT3jfw8n+/h07qyxzdZEZa+kCOjlq5SGhgnN
NxeH2Q6zsj4H/S1LJ2tgr7FNlwgNSSo4AQgtq64b3u+/iQnhJUQ+0HTRZp3OPgqSyOFsTQjl3U15
HmZAMSTHRugKYvgZl835d2/jYgLkqEXPgMqqRG7Zw+kaVxYsaHvfIbx/kLfA89b449xosFsH+HdV
o5l1/JRL9OdIm/74XY815fbRU8gToLRMv2m/iHQYd/sxeG7nnNgRAD7hUJHN8UzswxQ0gQQT4aO1
jReykJ7qxJljRzKKQ6e4qmolRSdlwu4BeMhCmAAg0xERKl88a+DkTaOiucZriCqbnJ4/GCK980Ro
zN4xK6xx+x/vrpHvLQaS1nN7T/q6RcH4Q19yQ55/SfsDx7eBEDHpdQx+jXcNHzzv1UYQFr4k2N04
JNMWro3DRb4Qs7j6pRBMPZPKIyuQycpEtl9Ig+eNWnUuqA85YYAtgJPLftzNfvcLZx1z2bkOBeOU
62PZgqp8fYP54LzUtJ71ttVscqt+f672oajcHAH/ysPv1XcTyhBXRq5TzZxY7klRLACqwiWlKQXp
P3s7IjObMwrt3r3vZRcqaf3bcw5tCPYBRzW9PFIjul58MoCAo3GT/EMupvi7zPMHRIKQtUfYrhwi
6MvxZVK/zNqjF/aZzCdzFnKc/lj8M+rBKLlHYWQmCaPVfumWKDDtxDxjLTFs7GfxtDkdsQzxOc+W
dgmQsBF6J2f0s8SEyfD52HVOJEhNIJcCkmmVJp+oAeUFPy/slTpL2vkIri2d33W8tz5A/UOspxwp
OHND5apFANY+6R0qVKBmSH4rk2de5Obq/PfYwlm53w5U+6defuPVqLCTSLUKlMTHpfHB4kvThsXR
9sARnW0SDmCkgx7jrzHe28Vb52VhQ5GC9W8E0Pf+yYw4DPOXYiABRBtmFPnlRrcWkOBhGx/+lmYJ
z4X64uXppQvvuXT1+nL7LEgV6Kz4UYet3YeRM72AafzsoBlPHGlnkI2pq17k7QG5w9Z4o7p2KXwR
a5oc67mtUUsE84h8Q54YMkUFAbvhoLBeYkLBcBlcBqbTgDnvd39KhGFAv3N4CjXmi+bB5rl++OD2
qrjoIb4cAyVwaEz7shTFUhoL06X1efq7jnAeidY8Krh6aw+Noa1DjXYgRQDb+UZxBt+ej+gf5t9I
o9VDXR9+4gcf+lKhJ5ERXStRagajmleaqpm/tZWM5DvU86wuxqGp1yYpCWYUA3d3MclU0YhtlUcg
lJp7Ax6GWhNENfqcs4+XQS5Dm6KN79SuvgFhr58s4ulHfWV43R0v/rU9BUpCOeV1PwbV0e2mjZto
HDrlqn8JKiKPAL2fBoKbkh4R91yOmEvE4YlqPA+xsF+h6LpdnsORwHqepQngjhuDbptV/xn3ktlp
cRP/Gy6YLSfbhPtRKAk/U/iLUhcRdYCg3kRXAwN+LNXYWNw2VFp0B69+zMp4lRlu1y+aQh+ovIO9
GqC6Ga8R5M3WUW5p+rgRV3fNsD4ZR7LSLghYGL+PilyX8gLj5NGjq5rs3Lb9Zk2JJDVWfswWmGxl
48PTXyeoPSwZPUJLbshueqSZM6Z24p5O7iJRPbVTF+XQSmR3aAT84JvmXUfvnrcUM6eIWOtqAXns
butmPk/ChwLXZYJI34zVho6LSy7wZbxFWu1EbM/rPpd2thFy0LOEDobKDO8aG19o/sBPFsigrwRi
uq4Xk1SKGZEucNibyiILR5d3RkUD0/n23jouBf0RqMam2MVIgx+9lk+GypQGbkdph1QhfRqlhE4i
UmKq4O32wln0hU88yiXTJ2gVoESEkqjgMOzkGRdG+OSRPcb+aNvFFfeY7t1YfnTJuv+o2NQPNOpe
NZ4tAf32y+JOcu8c75+r4d4qXbhhXzYcXhBtdzBKdeSyErNodESJAABe0VoN+IknIixqCn7u6b85
NuXuzad//plTuJuig0NLPKA9z064OVKRMifXtF5gpAOKL8BzZgPRvwaXbstrhXtUsttP6hGaTyHs
veDPw4GGiaFXoH7uHLW72EdF2H9G3dYYMzVYDpUsD2N0joRMLSmBGALila11EbGOhtynuMxknbVP
QAJgayc9RmfpwdwkRLGGSZ8eKGfaBDoAkB6F4SBJZzaHhy/AelWlAUdrFVGyfTCtNm5QwAYr19Ua
UjbwAU1MKm/TLgQUNOkorPrdl+tgEHKf+IS3fLTAec3kOPuMlTSlyiHr1YV5JYJNTqIVq3m3Fa0V
uH8tVgz5K5pVL9qrtJpquzSWG9OPaaQa8oLffLODdm7TF1OcJzH2wW2N4pYqOcpT4nBZOM1xA5WX
Rv5VepIcAszyWV/Wmzln1mJ2gLW6GyzLDBwXGh1lwkLZEo6f9FNGCOW1AF2biKzAe5bDfOS8qAzh
kgS4FAcTwNoiQ6UU1x0NNWIzA1Fc8hceNvYFveQODcJ8PGVKyFV8oiNp0gw7f7N/fUKcnfVzoQDE
oUozW7TzWWx7vf/b7Cre9fFSiPHSrIKbhMFlbVLHpcFjoDN6Ym1fYXe79KkQjGEeTwitlkRQRZWc
0WTm73Qm+szwVk/Xkipl3j1KSmdT/dzzhzdg4uVPPTWkVvyEcGurOq7bbEUpJessrki8T6ffuhwb
1eB6b8Civ9cHWESQBvGhDxVTdKqzrs46EU8MIFnrMdxC461RmYQ8O1ksJhCPYqLEEwGoqYmKikwZ
4OP/OzjIZxnTr1nQU8pyvD19GJzahuCBdU9Wo5cVCEZbPzxvURSuoUUEgEJMzfvtJrVng5f3Sk+D
fPQiiQ6+kRWs/eELr+8kcsDcblcwgKUUQYLvPJw7iruj7FsBeS+4PsX5EwQlp49atmyJiHWPQram
yjKCsZin+fBP2Bemyy3dlrPFRkrrKIN30fhSnul/m+degiy+afJ8NFm+5SWKiRRx0uE7JXCGgbPM
QzSUZ8BqEZPjIEhZR4VYRJIR0PdZNuly/x9ElG9S1OlCe2Dt7g3q5iG+1470Swt9XvkIQENDn6vr
Dc+Idu5+oXA4lheZ7mDkQAAf9bps86wi5pFd/wWDS1qEN3rdLlWooJFvnlDL0qYLnNuLfUMqG+cs
8aAYqEnZsQR4Vf7k9nSK1tYHNy/PJGfG+F2VspArycknBPcHtEzwdGlHtHwS0GqArHKscu3WenY4
VvHMEFSmpkVJXTZvPrRfJ4uxvIC0wZLpjHlkmHSddDg5duMPJIAxo6zQyO53Bw/6b2Z0s21ZJPbt
Vpxw8pzS50YwVqmmXLFrdI8HIrbp8Dw6H/cs9ck+E3x0tSeEOtzew6qacvS0clkHYtD6FWnc31E7
amLlyTngct20FJZfKYHX/RIDVN/wRhfax0F48XGYJC79egnAc8wBmn4M1DkYoL2/BL6r1wvgte9G
x+o03WNP7SUBrFCs//G2pbn5PLUhSm+o71+R01FEpD7gfZVGJK7URghnjxxVRja8WikSTD0nF2wy
6retbOWgoZzkjGeXRYzR4pdS3qAFvloIakm5rYqUqqh5U2hRFaVps4mQE0hebDDpDbJ/lGsiMnZa
//k3e4pWKz9PsTF8II94ZM6R4r6rDIybypYwUuJTQJhAIqsRm6v905Bt2geu/plx67M8ULZ1OdD3
V7etshUzCUhsVzFQwdUTesIaZ00D5h416v6nqZYe6TRhREt/gkrk67YJxroIJf5ZNKANPQ2fLLL1
S4BW9SI/b1TPcEhmdoqvLRYjudFsunUhwUZk7Iyf6SM6Gg4gR76rYACpAVnByIysLlun2f2coav2
qz0u0b8n/lN4orGjdVv5n8jrLEuVqkka7ykvbfAAm4Su1HUwtrzAQRStCGzUi/hGeaYfW4yzygeP
eGwjebMySBxDJroG0IV9MyMlounmTMAHAeM5948ZCOYWMvyxPTrNCXo/McX+B7HDReHSg2Cy3B8n
2hj8dYSayqDq5W6bpknMEUo30JA2E/C0OJIi+ZymkmAkW5TjIHHYWFvLyASULdOE+umzwV75Zi0d
yYlmcqvQMxrqKKjjqh9gnzQVRzcyt09i3xbHORLLNQAcnaQDWslvssQiztEBeUc+HUuf3w9UTVUn
FSWrfrQSs/4bEo/4BPY9/7BW+ySiiPBSXOhCdikzhJ20T5Du5YqEFQoLjupJXELTuvddOuBY1tz7
uL9VE4Bnt0Zi1jqGDRjbEzoB3GGed01tRxfL9lqW3flAxAZryPTkNSk6xKWhCByeHzZ9eaYgIYyz
Uol97yMKZZqsyB8NAqoh6d+di9EZRsskC0i4oYUakv7vliH/PINH1VXIQUtqkZI7O4systfnz+3k
B/UBXFc7JbQ9ubgTmRVV0cSLUUDFIinw1XUtmM4Pe3UsoSiMX3TBcEy0AzLV6PEDdtU1Pc8bZHE4
gmHE7XQO8GimfwkPVHSTktrwCblMTFXFU18lFdWYkHrfOXKqgOtc53Yv9dEiUfedFyEIkxBdK8zL
5qfW1NCP1v8ZqQ9v1A9vbKo0HO9tuBxp8ySPiWt1viLtrx5kPCnjkG2/yIuNbflRv24+7EmbbuqN
rYDzu5l03H7V43UP1pK9LSd7OIPs3SmSbIs2keQXZiUk+XmTMXiY0gMWl2LR3W0VXxI0e0XeSzLG
HrS/e/hIDYqZL9qwGTAwQHo5PN8cid+fEpoEI3+xL/9d+jMftZyCkr1iGzZCtRymb5nOj0dd+M47
XlKrvEjM/pgtBpqGUXrD1Yxmmo3JCvzOiPrHC8Wg/VH67ApBsZ5S+p61VSDlKGA63ax8h8IX1Ir8
iBs1vvzPdstQPBqBIXs3ccmrUYU3evvEY0kxKt983TusjpKo5S6Uxd5qO9lXbiLRz0GtBYWqeKF3
0gsTVnquL5/rH8EAHWe9dL3iOimibKhVOinUNdxxjncCYVzWkmcQPcoLG2sPoupK9u2EnlhdsgCW
pBBem68orP1hsp80jY510amMSSZ3XEJRO1PWHMConZ+bouSVOkyiKKq32+fZPOcpkXoiNhSspFt/
DWCaxcrHB/YrTa8YUO/wQDdHdQ1CHun+zjMmKqUz3FvvPV3+34AM3qqdoDwekYNTIXqqLdjdsu8Z
G7M9zEaDWfYBKiO6jD793iBY/U4fvk+AS/njwn/z58Xvg2sd0D9UVUy2O3tYW+abrN8ulllWql5H
eN/A26acxvhdAaFi+LkDyVnXDBHwBbXaQSWA/lO8yU6wbxwjIhTPVnsIOuK0qCRIy07a5SHLMgzL
A4vK+N6/vI/amjLBhRQn12OzOgidJURPWtnCo80GPmSOdMAFW7qPX0uYwgkG50eYI3AqHvr1X1F4
tcyTmWrukD+CbmYA3aU1y9Xc1f91dyH4tzPb6W5axpv7t5fn9/T2KAVf9w4AyGaERHs7scZp/iWo
eX330i3Oy7h1oYnoMIVTJO0KZqzX1RAn8xaW0wmRRtVQRcuJICozp3U5OC7sPgnR7PxhvuJqyZQI
VwJQ+wIa0dufXJzpy71e1dMlOJCcpJQQH7ABnzViGgciYJ7GbfhzxqZOnacfT/2hOOgKP9pFbZRV
1QD6SDyBxgvAyxYtWlNWE+YGfbXGyF4qf9uR2q5Hx/J8CdBZhZ1rv3L6cYoF+HZfgoXxrrlsCGEq
7ZXeVRD5rl2BZEaX+X6IIGu25VDhv3fDCAKG4bYO4iHAIlGFKddJ2UGkPEFMWak0ECyX1bzUc6ae
vxCzyVyAF6eEVrUrrjajRHlKiOeoHZcs39HnwT7WsOgRg6Z0fmExsZN8Uznu7dLQ1DvRxz5zX2oB
ML75iHv+gr2OVcBRDQ3ZOjPoeXHmz+ByHFg/e6XohGeGbvVlPnRDFhYkz6GFmEfBvYsLfdI/ZzSo
f16JYwQAYnRSOCnSDo0cNBedd4xt1G2XlgAJOB9j5LGy/2HCa4TLZVr5mr6zas+8KYN4abZp9UEA
b/aJvj/e4NyR3hKNCEjK0RZM+I+VkqJ3hCKBo6YXM92wpmde0p1BUjr0OlVYXkHigVnm3s3O7jfA
EuywzZ7e1AutqkQbHlknBL28+z//Js7J+nWV0Toh7pnxogoNl07PWqAzx4vDId3SniHRPgxJJzOr
Dl/Bq2/7WtLIXAXbKrDy66BOHve//7dDjIbx8c8I+qOFVy0Sx2y3/HTk42sDN34IUzkd+dW5KUHo
76Yuc6leUspzlvxrGi49k0Va1cCZnUhppZA2wbS/NZXEP1vHkwrPrHrIVgVOOSvXbl7W2eLJzGM0
3qcQTFMDoOVjqznfDdEib8uoxuiV7Yx3qGEgZAl7sj+3jbbRqgjPWjw0gF3P5mWGXfDdr3C+wxg8
Uq1CS8At4xQzKAW8hRZpxPCqixXfYW7JNwxD0qsox6o0QOIT9DgKqDqiCO5dDKIzS7DIpKjDtYre
mVxoXoX7alE/lrtQY4BIJOq4Uf5g7NZcEcrvLVkUcNUHbCvYhXWLfXVk34zhh3eY6gacwfvmJQVc
Ev3dmasEISa0MGjrjc4Sf3SgeNs1+iv4IEpmdBNUGw6ekSsxnq+bekpSK5d4b4W6e5rl9Gy7u45N
fxr0pMvPsZSxsRW48a0Sg+tFq2aq1KnT17JnbazmtWX1r9Ry9EKB6wWsUPYNnaoTc2X8SXHrkdwf
MhL0zG1aoarBZNzEx/tTUZSCBcgNz0hG3302PhXhEWlqUSMN1LzBmGtd+rCQ8H0o2Be2RK6hHh72
bBCQxLzo8OD52/xucX6tNyQCgG+8b2LWvBReNxKtamU295lq8cLs705zWkHlldWJtIPrLfFCr5Lg
sxT0/qfo72GINCrwIr2EVpPWdmS5cojW5wZXXuKcEri/dUws7JYgs6HgrqSn/wGqyt6jq42y7/EK
ZCsjOb+x2xAIHt15BIMa0l1QHZRCV7LGtBxJ8kFPsnYmhMxVDa8XgTPi9bQhw7VPdSaXdxlN0B1H
oA4LsHA0brnUANDZgsKw9grhqZzgFzgrPOk21aErQIyCRYoGUH94kC+ViYfMauKlEiCXP1EnafkH
+BrZsP27lJQZA+nbH+drtmE4dHsMokbwi5w86e5hCznLB1sFMaoWVCYNa/delYsdV+0P6RWt8R9Y
hS001/gO0xxDMSpPQ++9hRVWQAo6Dz6Qve3Noc+g/4JhJxMyNOsDq+WIHq71pgEzaN/AqAp3UFz+
HB+L+WtI/UetDzbf/OQREHu5Tl6qLUIMxv0Sem1E73k4h1qXJYB2QLqcghchYrU2AUa06T+1C0lj
VjISSTybMqeRbs4vRXQwHXG5LAh7E156w1gDo28Dj3wuU/4GGO5O9dox3eCkeWIZauawB5RqsgY3
MwZH53JIOI6slKPC2/sorH/bxmNwHJudaXAnxRkQdv1wlXXmDAvl6khuzA362okrGA0XOcdtQlw9
Hd9BqYw3v3MKLo0RxnzY0FRpMZlUrg03/y4zDO390xG+Ld66opm54evM1k3qrZTtg/vassLxPl/o
vBdK21vzh8gQqO9WOn4S9psnm/C0ocQ48k2sSH3W90IK/oIei4Sjw8SLUCzfz0LBP2XvhSECH/gK
OoTN6GHD9l7djz0s2Ivj2DYCc9dTXE46AUawc4AzaBDqmhn+Sqe4As/aBnzjruixEWNwuOc+D8dM
OEiKJts52+AKZUpINIvnnCclTN+3u1kolrzeN0jBOEep2C4djhjB8WeAX7IMreuJVM+u4kyfCyNc
yM2r/KeAarijkqf88I5QoxXp7NLh8l+WPTBts6p8AehG+WydHHGT+004RQSZ0eARCNltZbl1h5De
ygJ8J28QMpHTICk9+PSefIM/YSLbfyvi0zdvc2aN0oiDbaWCB9sGnFX8tzUC/nlHd9wwy8zWqhjv
j9JfEJGvonz5SoiQPGBdUDN2aEbZ02KRD3JEga+mw6jULk3qOWM7AY4XTB6jI1ebf3xtVXAFBxvP
XKN/KvDoi5UOiHF44Jzr7aJVLVSwiCEFWfheFysI4gLzu863plYBmWn58rBqa4NqhDcVot0/Khmb
NRN3+F8B4Zuhl9A6gR2dv+FxHth9QXtZKrSUvvW5IOfMn5has7Y0p6+OH+4JQ0mBNiB8tRzNdQR6
5tF59+LeVrGas69YZ+B/5CbauknRfrzbzm1SxgVre1cskHUgUGXvDuETLe7Tey4jUzJ/1FRNtFdB
EZnECM5Brv++Vuh/g8qHjeUs1IUduNP/WkXuKgJVXNDFF7SfhZlflJC6CeYLrEFQu09MJXGvHnvt
/w7gnSDppWJxqvotcoiGmQ4lLEWGkxsCWDcFKBpOXpmgu6R/dLAmx1au4tLSxlXgqQKVlnNwlkLf
VldTU5TBamD5O/meBX554cc3wMdQDo0PQWeRUw3WTru4piZWXVBptv44ojCkt2sw/DdjV0Jt5TaI
tVCRXXDCQBzSW119JXKq5Wlh3xM5XM9qCw7g3FEgVufBiShWYud4UnDS+wz16Hpbz4LB+4VmYDGF
On4VOPLQx5Q36Twdrw8+f9wSXmBEweIOHssdX7cD0XCdZhCVQf7iMN7rsoC1EQ+hALD5nhf39uGl
RcV9EZDkqt6QCrfnwbzUsSmqx+fLnh1BiWeUpGQCNxqTaEal/8voWm/NS3xgC6lVunlxcSkLAkAv
5boH5WYOJDo7vSvskkf4s9EyNUosN04tOjJnQWm0q+XxKjolBDBeH+m4eZkUTpGLBBI0r/JOVW1M
RA7LMCX6whdY4EnfXFX5GbiHHTOM+wRzTOvPXyQJXP4bLy9TdWvF/cbS3iKW3ysaLzv1adOs8ihm
BjSDzbJyZBq7dsiIhqEY3PuTVRe+wUO4u3/8UMfdDBpueX4dGrpOV4yuPqpH3rsaezQ30Ty4yzPI
yKZlSbC2ydv704F/4iIcoIji6dUCmgUvApPz2BVJKq6vn6EJkzqltMa0iBlwdX+9uv3h3cjx3VMs
igyI4wgWCkdiE6omzc4K7eYjMhLImmQ4vmJwxm2Pcp/cGiYQ+s/MrsHvKirz38X9BnsmajnaLjjp
QpsXIEwC+MZwfJo75UYbWW7it649+0rrsVNH6LYlTTgVZjhs1MNoq+tgUkByAK18SvU3J3fwre19
hubl/GZgPz2l//ucN/0NoVLBFK2p+xGW/c8Yl24Nz0EQUM8W2Eu+TRxo3+gEe/t/KX9/vI6y6dGk
r5jnBSADbCLPZzPm0OxePpNSGXVivrdMAm8WIBCMvZFVf78zGoNnsTZaPfUH7mARQ19sUwy+cgP+
kzTHs+2xD1BPc6NBaZ2qlA/TsqtmQVJ8TrmTZHaBz6NHaaQGz9rOKpHunV3G4f1ztgxEuUqpCdI5
v8IHtvSRK461Aqu6aDpSNFP7erUE1+jzLwWsiArgDqkoiD37SuJ3PsxKM67OfZ2xk3VuwE4hJxX1
10OaQpnzCPFXDvbSoNaLrIGm5BjiAV7zqOapMI098iauOo0cfW7MbWz9eEk89DKc2T0Nct/+cXel
Xq1Ily+jReAke/IwNPIrNWzH4GbHkrw5KCI5O+AIJu+tUV+hzOdbwSP5J3dZ/iUCeah70R8MInh6
2/oHXFN2WeHlRF2NQqihOaog6ZEEH0USSOt3vz3Z4T1+8VzLOb41ACN85B1OuLBoX2P5O+PDdTwn
NpH1dnswhTq0fUEZY28m25Y78wM2/RuHmABldE/2+yxfWni27JNP4JGXCSKw8AyJXE42w0DF5Tem
9CRs54JA//i9RaoUIZj6UBPa0dlL8cKS5nnOfbB2/D2wmIY0E4wCCDHVZSNfuhvZCr6T+EMrvjjg
FNDSnnhNK9jyuHA3QZPujX3MDjRdwFjOL3Jb7KXBYGOPE3A8ZBluc6pLSl8b1s1JDt7uus2SmmM8
IR7s/67qEu2erMDIiIP0kBe6hyJgN1hDOjFkUsIFc4nNDvmtimV26TMdO1zNv069JmUV0UqORsBI
GR8slDl65GcICY/pGw+m82onAO+oQDZl3h14WMi8MaZQx9BI35ndokdKEOxP/S85Tud53n3ZuiGK
3/3F3C21NZ9RN/TnkYW8OwQyNnog72NYtWaSEzNMuexgZrWQpPp4OFY/omJA/wVjtyOS7Fk9qvfJ
6ugNomDfOhVFIJGMADDv7qjgVWR8mzioMmisACDHGNJcD1DUIqzQsRsx0ewuyS1adoSDcj9xCsQ8
KM0cSaXxD49B/RabBhxMBDyVrjjJZ3Vdd9qj98StqB3yXzU7sc/61iNvRdbpUzEIQlL+WJFXA5CZ
tVGmEULcy1uUOO+5PxoDuEwlMActYiODrljGhGJa8bSj36uGoLpSTtJnPcwNgBpHCLAB6JaqlfNj
rnJJ0auRn2iuH59rLQsCBa9+RV4L43dUM8Ckb0wlBf86uC+TJAxFYJNC+2x50ZrzxpYieBG6EUA2
7mXZ6Y0+nFI2St4ntn71tahp9SA0Bep4A0BWnemg8QlYigk/lPKU/8TVJkMYivCOLgDBfPbKnR84
xMOWBcG2ksuqc37yxbhChacAQ7xTRBPXC2xNf+hzdAOOP092iYus+OSuFwpQ8LxTsG4tbKsm8pzr
NW73zAjeRf+vuTyd8/M94tAS6zFxXOnETcNpPcSPdajwb/FNtDipVKAj7qj2GZV7hvCUQwbgO5Iv
u5lRE+sMPWO5sxuTkwojX2auXiTXgg1dDPhZB6DVRpHZAlc/UNTKCBnrOWU3yaVPayAp5cMavup+
ICYEn5mYVtoIPUWLO455V59CuW2uB2d8+YhvMehkAE5Rc/qA0x8jiPXxKH8KR0fpKXnvlkH7LQmU
XpWYu2Ss09ZXDXOa39nl6rtrB8bxH0mfDTZhvHHzzpVvJyyKSlrndnNnnfhgtQAYx76nCnY3cW59
Au6w8CnVmQKyBgaLhdZe67QhNKEF8UOhVm7sN38ctvIUwxW+RWudsSInk12ZqWc04R77oBK/FDJK
dXpeqvpWk6PeWW+UJE38opOW3eZwSYhQMiK5gR9mCQiJjIjRHSP0wRJ5A3QpUCboII53QjaWHQuG
ZGvguUUIcPx2PySlRJgN28P7vA6M403aS8RGrf8PL4N2rua5ek336H3L/BL+iGaSPI/w9qZLy4Oe
ziUYtZzznDJErn+W/8Ms5GwD/2vqMoEEfxhEtk4NuyTgH5fxL9Js+DAk7466YSK7WxKffZ8CDVAS
8bQbQEyZuWyMBPtAhrNGuAFXkqUBBF/xH+N0/LOiexbP3ZdWwvVJXJMNswnghCGuCjaMz8UNtX0e
CR8CSsWtQND4JpuJ0i1jUvsR6v9paNhxq+LOHcBRhQpM0CHemve2piE6DFjQsXi3iFE8UExQ+wWM
ymrcKAH1E+tkyHJWh43jLMfBtEb7HT97uIfHOmB5OPnKNIDqKGrv41zdBYQnZ5TmFFBfrRLNhh6F
4H5n7/pQNf9gf8FK534+vIhcaa/gmUF+xfpCoHoAYNK9k2A+T5xGaKUw1m2Zg22jufYaIh1Hfsqn
L1mQI+emOkY9BorG5sBmAfUej/7xTwuLT/vskKe68RorAYe0qWzP5nzy1cf3bq4WzHxX4ECrXt32
6ktWimmVrgRXkPW16Bc5ycflY1pdo07sFzMm1N5XRodl263TAvmA/iSZlIYLaQe+Aj5/IiStvtof
agZWt+1m3yiJBbO/HRCjg5e7hBBsaNu4bW5znH5RyIHvHvE42k3dEwQfKEv5lgk/QeG9tkXIxK/S
6VqytOtp/2QJnIFOz8F4CArEdWItBQLUnHZ5Yy6I/QwAMqAfSoFw6XBAOiubBG/xrhrybqzvoZn7
RCTvQ+A09H19ByXyLsY2Nic5jpRLZLypquN6UKFdWiZc8IZj0x6a+Uvz8/SOBTsuoEWXaR4CpF++
MjYtVgqLN/ZPOEPl3ZQXVJFVhRJiRwXvLh8k3FtwEZB9lr4N/GOTphvyz6Cgd+m0MskCpQTTnltt
4ZJ6vQwYy+Xa9iinMwyQ12sPrNth28efABUiJ0Q0CPjcZsDCvi3QNVYFJ5pTqUbce6x4XPvAF/z7
Rsgjro1srumxUWJWHiK6WDrXaVrYyzYrjURnBJpyl4MnTjPaFuPTcdOOZJ+g7pCP7GHZAdPMGrsp
DUirmAWx5zwOtgVbSnDM1hCILYP9mlprEIfLtBRqr4jPDIv8Zpq4ifeoWi3J4irCA1alWmAOUmqa
DA4QzfaHzioqT9n1enDqmUBSUGE9ZKFEt54VZ/eSzy2EIWtop1RiZouqQAP0IbRTPfeeMDZu0vpY
AgePIddkHytj8W+FUOfti4dVjdwpfC9OKVYKuAZWCd3PGxEbZbm8awzeCu0N9817sOQAdqaT/nLR
sNn0cVedX9Sc2Bef1feFJKMI/lseBvjbD03P7ZKI5BSjSJMcPBs3aWCgYyKsYsXyLOv1ytz6e+lh
R4kSwS0mtM9F0JNJs3fUWDRCeUe7dwobzxAs9Ri3bMLPcF2L9p7ajznk6ZOn+hFHTeKUFqniUEg6
V1/ndvqxpwTQAGuZ6aIzwi0LCJS4/z6o+w7w3iae6aMUBz7qdclp7aGOtCaeltU1KWlloPQNR+lV
7MuA1cenP8aCZqXXoa/HWO7x3tQK938Q5J8q7lVZ3b6er2wXVT9Uyl17aHp/YgCpB0BliVp0RoXD
5fRSGl41CbeRt2Ty51g8rNu2uewIMxGaeFrk1knY6fd9zwQExX0e2bqpnd87ucWVRQPepO17hxax
mIiHFo19ZXzou74eHbIbV4kqobQ3lnANC1Y9NyYpDJ94f1qiVa50ylIddbvhzH00I8SgyIHxBCfs
JUzGngf26TnXsRq9cIU754x9jaYBRyMo9SWcc3Dw1d/EU5kCzM8sNZ7bm2nUwKwRl3dGS5JE/YEX
zu73Uv8RPEJVOTl2ZRCt/MhWhiZwfmIUF1PWUeF9T25y/IFv0q0wP2fgmw5G+UHPS8vpMzu66cyG
VNe/bGq4i2MyGf2oMDAx3pCoSFEiB0gc4NMAkKlGsJjd7Wet4rge5tuyd/r82PoycV4YuyjpoOGy
uZ2Rz4/eKvi/mqvTYgoyO0V/kn0k6oDXfNymgd5PKG+AEL3yC0jZZ1g/61j4cMzB6qR1EdANp+4b
VdMR7NxDJQ+XZJ9AOZcMTbPC+0M55cxmUGxvv0Q/fQsz0E+qM0VHjcynGBTUbo93QRtfdrHS4Y30
9Syz3ULLsLQXHhul3L8G021+kaj23RflrNX6pCBatgL6ypdQ8YCw0bTphwLrbG/iyVcaqCNNHCHT
8FdH77TZZIxABBKdRCoxyejURbrSkAY4C+qVbohhlsRB6GMLDgaIPyQpqWU5Mk0UA4au++sD8tNS
+613nNh2ceGaWTasMX980UTva6qOGknNlcbhyx2SZOq85up1q4IrTnXVkDM7ng63Qs+9KkYYGErU
UWYvLHorpZBVVypMSFjV9r03MixuMpwpfkZWdZ5Zpp4L/GtWhUi4sy0z+M6NXqdeZ0C1XAuRIvtw
2phn1dqQvpBn80bCZEMSHhd9jgGP2HAL+zJ3LPMJkJkUQLoPwVAMBBxLAtbSDH6nN9a1MIr8F97N
3Yu8TQydxxNEY8wvXB8ZrYuXZRreMd7r+DqfvLSJ/jbkNlRiHEKVwMVk+2WtkNRw7FpK+IWgmoU7
ZweXHp+cHCYg0XefE/rnYYhabZWkne3ccSWOte4f4rQ7OzrKM93cFn7uFZ9hnTOzrQN+Yq5n6U2e
6cFLJjcvzsJUasfEzVqnXKGLoQTAaUDQGMcu6L0XAe5Z5N+DIV/k+rlx7fuvDSdarhPfUk/nBLqR
vto4H6DKhva2/lbX9u+FbpMXdWFzSSnktLw2Xxfjy8XqpLKah2LCjL+FsqrBp6gda9N3obFZHd/1
kITCq3/5+FmQ70qDGV8tAekLU8TLxCnxIuOLzx9rtTootm31r9r9ZeMKpvzKPeq1v2J5/WgCHucv
/4ExlGnvof7eYxFfUIoGCRvwIFJN0ddVZ/WXavAYKTCdwN5jpsjvGF+eqC11SeVVfJeP/C8OpBF3
JoFnVHRP4hc++Je8MPMCi/qQJwEvslfPUjHbYygg8zxu4u83sATz4XvJOlVb3CfdCP5kru9oKU/C
FXGStQjJieaj8eKZYYI+rxbHbSzkZM55TC+paB7lgpYmYkI/0mP0iNN406MA8u+jGbcmzvnnoShV
rogP4MDB2EMrG03hCEaxikj7NWZF5MSgn2WiIuSZBX8JVo04P6XTJ5zOsVeBOe/+WoKWrSeuUqHa
I4juUi3vQcZ5Y6TEHo/uHJFu43UN5e8NoQm/gOZ8a2WROfJYpv3KZK9d8jd8MSI34+cB4CqYOhZf
Ve5BUGHcbqXJmTbpetUy4PZxAl7R/J/W/qDDKn2eRmhz8v+3MaEpWfIeDNkjs7XxtVBBVDFpOE4w
mZwvnUvT/TljT5EFgz2EyEgdVaPNYX9IEo3BGYm7mp6U49QZ22JLY2NN9yGUZ3juG7CYkh5anwBj
sm3D05LMOgko5pICLmelhinWxXiTU3NOsnuB2MDXbe7xFgb7UTCD63lVwgYV4JE1wDW1iZAWFqfk
LoWJzPfTLTUgNuZVd/Q0ZEJCzLMPTnvEqkiyTY6OLTKcu0ryHmmnjpi/9z+2AlNz3dzBQgBRFjw8
qkWuhMKcycDuv4x/eryH1pI56ipctMJXzDE36WcvS0T6zTlAQhxi/nYpWJnZ4zs4WR0WyzIIGr0f
rJtB8Y/wiESvmNmzBTOKvoeoqQEAqlB23+oFi/SfjccYwCJzgGkbC9Ekg69UDkXeWIHJh3q5l2th
185aVxGQOfxITK5d3gnnXUs8Af83DIV017xL0W1OlI3ihnaiVjupUWELcAV2zrv1zaAcMHYFPpmf
MszX6IYvsdyK2b4vERmTq5q2WTUHdlQs4F98e0HWnUHPSAYiIdaDHYUUp3nXXiwALiU/OWs/bB35
vp0u6zU8R9L3W4BHv/XWW4SEDcuyiJWXBcs1lz4NltHE1hM9gJkFlq21JiDVM7oX2RGIGFxcTGx9
UvDg8Da4fOiuzZ6N3/vSFYmaDUyk2cLn8PoH6Ez8MBKe9HJlLwQPqa6nu8jV7dqq2SBUPisNbvv6
qtcnC4ucKtfC5Uf2YfQhgtuX5C/oiYW1JPSxgcuKK/PMpjBj4tK3n3ZLwNWEgAgSITzLXhq14q2I
rT7Vluxgi9dRlEv1rXsFZTa66j/kGori1DF4ajjkOoMXtmagmFHMLwDExueLq1e9hDnC6eQ7+vs6
oJLbv7DLYBuhKBaOIiCIvrZk+34GVDwwHw9jlRYwNGMc6QRYtBtYIV8bbJEnh8/f6cZDe2aeWcwm
kKfKjX3NfwZLYn1RjIFN7AHMG2qyn9YqWDwUIUIU8g8JLehMoR4KJS69RyuA7UhlO9utn+08E3j8
lZj6Ln5nRCtSUUp/l0x1lF892e6uKN1Oi7AGg/ZH3zWsjJqs4M/H8ic6L/vnwIlCIGYfeaAS9hZ+
OBui3oCqa1q5bB5MkjS9N72L6XLxdxA2/Phlh8VE9sPSW85bTDg+dYfMnaYIK0UWMvA1KzuLLYnq
OeQO4L6dbx3BlZ92qDltDT9K3ZhbdY9A4RrIqQlFfUhioFEFRiNYltIKAlGzuA0W59WI5zI+w1Tm
ISPR0Hg1Io1waWL3/GYAuw4JSWp4ytjyKK/ctYH7p1X4uv51+ldQicM3gf9Uh4IrPcRA0JXaZiyx
qFgfkLxFo0CMn/KN97BXSvShnbgsJLZlQ+TrTqjblySXyQj75gWqsKGrYLx6u9rBwURWeLaVUw+3
G1XP+iKjrcCJgN5KNFW6BnP2sj5aN0HCPqwu//H7K2N6IiNDybVr3qWOHYJfyEol7CBP6WMrohfr
U1faTEe00T1h1T61tdTI6UCFa6nI98wPRVFowl6cEffQAAarBIV6Kn1X1i3JK1Lhzm2rc1GLJ/u4
uuCmKVO8W5YIFe9L5URxF3NaaPlU7PCCihhik8UvtZhNKkl0BPGUL5cD4CQmhPrOGnX/2idC3RQE
XOqhmwnd4/CQX3e6k+e0NTYqkp9NpWoMCstxVPnS0U5aJ1fQR9/2X71epPkt2QWT6gslwbWjJPQI
U+0kYg+zXuUm8CFRdp5usYhNgknCyILINEiR1nytAlkn8l2J6sRZ/GuAENCQ8wBHxuKAlB6tfvU4
Pslm58UmrEGB0DJcHON6+gWCsa7Dear6cYssFV2odmtnsHsulGjg8xMxGVhGQzivbaA2YsXlBSf0
mPnUBiLdFn86RdOQ2s6mNuSxVxNk/mUglaJfTkS21MMkO7yswq6yiHG4w0M/rL12Ar3bJUxd6KLA
t0UuUkcStTg23xLwiAGuqNoPxyLDpdcQRhB2kYb+SQQMMVyXHqufX7b87If3QZqdO2PJHm8k5tGi
/SU3z/PXyGne7TK0LSkndS0b8kEqscsKwHSxMjeFcPgQb1E8P+TrzGdT5G+T2RmM7+k5Etsr5N4h
9OBfMCPQp3Z2Eqoxe3JlYFseMwJbxSXmyxaAXSvyEPPurVaakmbCMhF6qRuak6oUN0s5NzdFdn2c
Cm/WfKi8TllaDfMf0NtMzQgjNyzP0zYkKDf7E63U0Wm74pi/6fh82IWBQwMZUOFp6OZuTM7Wklkq
R3wd/oiOmAheDRl/wmgqztgvwg7tIFjtgIlDBEQ9sD7hxy8FkUQQl5umePRxDbYZCzkaGnl4flip
FeYnZ4J5z10bqKkM9IWsoTMILEeny//nlYDOLT1iISpGvZgMK5+C8lAsYBq548zM5zVufqqMht5S
ivOFmxvk+4ngkZ9X92uealteeQM7KJfBM6ubJZ7hUS8C5zL9rb8jlq4oXMcG1G5oaGyulc6kxMTw
6nrCjwhFWIdFXbwOplEgK9wiwwcLQkBUCp0flku1b82M93GG/JzuDYqwUvCLdG7/+2qBUujE2cXR
mUPCp8QLJuLlS/ODhqPRJp4yTy1hJOj98X8omKcLg3fgVB8NDZ6e4AX5DAxAwkFtMbu3cfDHAIZe
zD5FgqWMjMQJ7KVCbnXypUQm70uEMplYU81VH8+cei51E7Dg1+N3mpB3JNpjQz8J28fh4sCFFF4u
j8R1C+N6LR6JBzagXsag5HXnkXD/Rn+pHbVlrq1vE1Gt2XkoXMemv9OEKcXC6uHTsBnU6J3FECeN
YCeTgaLoScHNoPXIYW6E+obU8Na/YkChv5PrirdD0AT5M7IEXz4k6tDFPzLQKa2W4wEtgZeB4nZ1
9Fjg2yzOAraoQpIn3haa18DFJ1VzHY46Oqer61eGB7whmGIcddKmPty5aAWrP3OVzpY9BORf/oVj
pJXsrSwoXmi7RU9CzG6Jo1LVfKCb3rRqJ3jW2Vpr2pD8Eka3eDaDD5VOWVfC89dPw0H4Cm5lZUL+
dbawq8ciGBW2sNDDgI2+79C1YqPG/Z0dNbVQC6XmrwNH8mhRXHDSa74esnRKYVBEi+g5val1lLHE
NnfCIpxbqZjzPE16BjwzHHPeQpi37WrEsQk8jVDpu19Y0i74t9u7brlIyLda4PnQhodxj8Z/bhhK
jQLGPXV20RpZiOtK11er9d6ZpbkKJQNemkOsN6Yk/PLuKHgQx6mONn7BDV7HV+J3UPNltIlXRlM/
J8xQQZqmNi7HpaYxnfuhGbNR9fuCzlDZAV8+4EQFa7PLm//v5KEuf134JORmAFHKM1oKEH9KHRop
Ryy5DmdczOKB1FBuUle4CLcZaPiyRqLnaSUj1lUQ5aJz+QVC+RUv2IpCVXK9LmmfZfx4U3VCj82/
PM2DYkAse+BBSeEBjJcrraAu53htSyCVqe76dRYWx8vFZpp/cIeVdHBJptAlcIOnAASZy4DOSrAF
jZPgeNvWzhNnFJK27phrLqJMkB2H0sYMoY8Dt0rG4+twU0ix19RJqzAoEEz/Fe4GhS0fWt4lpLEQ
ZfABiqRAzinwasWMOAzKwarp4jPeVTOm8W8qfUeAsDnY8fUHfHq6wMm/r5WRJYreUr6B1nOSqWLK
DpxSyzZ0pX8JXhcAII2ph+jNltKRWizA30OUvFE5dAIRSV5JziuXmxKQmp2vzjtqAXSpIG8kxBRp
89s+vlNBWiDJ+7RnxwGHjauULVpg6+PyMN1KZsZSlJ8LLYnA5X259IaHGb8RTPOhKbXQoGGn0c8d
LylxaXofLjTbc7ligjZRml4BJm1etbwHZfQPchx5PvxMWQ0TNdR4QeVNC20YVAXsHvENXAGFFl9L
ApfarLsxO+bphhUbPSXoJS0NW6i1hxJbdhxfmnUb1va9O0LyVEiOhFrlF/0PkZyutHJ7cfLLeWTU
qPXY3K5cMVZXwGM0AHwTCEH6QoHX4Ap5OMbY6/J/uiFbbxVIDMoOJyh3USFNwAII6hGfu8scoQ5q
078v7o90eHx6vzvZSdgfcPw0YQ1g8cNUPI7VRgfJZhh5JXS1l2h0dR4w3ZO4rh5gH0Dlp9wkWhNN
UENDVeDEqCLw5IfQMSe6T75p9rvCu61f+jrfAlh3yPFve60jF0X9mQCaVFImfEkWbSDTLs6RVghq
UHgIxDP0FOWlwjCcjexvWKorJf3zKgF+aztCybxDb6Kko2uvytbyrGSbA73n2U9RY9FK6BjnWN9j
xJFDQ8jRVKju9TcLE22A1XwE7Jju/ibTMGK1N2MERJ4dqOtzwYvb4tKa770ObB4Z1ZmpsB2iwfbA
oTcIJsao1mrwE7GPEAyYYBHMkD9h8KbwVAaN/1vCl6tpzZfWsj+0U/xHanAgkEiEzp7p2SN7icUQ
ft58qyi2Xwco12vUqJyMODqoLWFT5VmL/VAlnSEVQZSs0vHgdbwWx1/UfCNcqXFE+blQ3g2aCMQJ
KVR90gxxtMrThV+z/dya1dRKNY/hRc1qlpUuW7pDx2aP5Ax25DnDhl0osI9tGLGk3mHLNrblAfKu
rzycTrl4E/C/RCeI0blHhCAScFuYOgmiIiC1pFzUlzjIUYNU9mhLcGRU71fl9RKW5b3mRTrgp6CT
I0P8oSrNIKnCFYXVjlaR4bI2xf3GvzhMXrDcX4iEDF0+dRB8B6aukonvJTAFOsjaeoZnB3bIcL8q
2wqKdEFL1RwZpH7h351hfZzbO9maFYPBPXrR5YlUtL6JbOfW6vpJ7SIBF9+V3l9I4eCwIgqdMhSk
4aJ4uhZXR76j2VCMjaS9hN/uEFcPU00aAYs1BA76bTfYi2wPNT1d3L/OdrAZ9+l7C+UAjWj0/vG+
1mdV5QxuSNINW2GX081Y24CIsDLaAV+F9laW4lVTt700J+7DBaek+sNCoFXUXqJpMrH+Je1T+9/j
mQjvfauO/9huOY/DVU2weAF7gzRjTtLNj/pOFXCI4tGTNnLGu0QmRVL8OyRdE4vE0+9zHUYTxaHf
0gFAXAsaM4neZgREmYrflqCJTCnzOr/pgeL/c0Wm01TvzTnAIFlaOMUpXdUktLy87lHRti7AOrL2
SBLQBX+dSha0RxJJF7FR2alAUy7JReT6zmdHLsI7Rv8i/+AOSc4GMtrEHnAqzpotnYE6ZQDGjQx+
oAGiX2u5G/AeELIeAkyLd4ef2ekFy2rJCTMHtfNu/9AmUyOUdlt8280uj1fkRyscYFUHfrjCq5wZ
yPAvo6Lno8iQG1anvnF+CN2wPK8IfSf5Fewo+90eGMSUbU7LNsZY3B4L/2+n+HRdwZ1+NBWErj5C
IpTAYzKMKPLu4m7XhYOntjPke1oSwpfZJ6+clNhWMykupuCAOdp0kbUuAEDuzPxs7qnH8/VMdVNR
2j4LoVPPLBQUDbSrIWt8/M5ZHxs9IcJjw4S0+Wd2Z/l2Mu7TuZ2D/PNGSxUTCZFPuERPyP6nv32W
g/ZTT69BgaGnt0Ke0YvgsMMbEYOHFCctq/XPI0BE5mADE79PSoNoMJMgn6JJcpquI7zuAgXfr8QM
OcSIVY7m/gT7YczuBzo8G54H5ZOlZYoSY/dMWKg3oFOIoOZTM3tQNUb+wkwxCHJDrc6T3yYolmN/
b9TvzPOsewCdvzif6ty1D8yJnDqMXFQwPzdBCY/x3/velpWJd7MaqKVlAgs2ts9XVoYqhdCQZi8B
Ym1D92ZAoeSqQBEPwXoyIMxyDYOUpHy74RvUlb5IvCZ4J6RfjB07XrjA4EACOjwd1mdGOpHJv0w7
5S05y80hLJr0HiZ97W8x5zcWGmZbV5wh4lBJ2lfiPptsRoigqsDnq5jOp9QthuYDUpIsjJNwt+86
374aP+fDNt/4EIsKFkp+1poMhvGIQe/FtvWvi5hdySs8WnpfRSABqknufPoDpKD4V8w966qHHWC1
n/xvI1K4W+jXWiaLAYqyshUMv8S98Id6xZfKmu9KLiADorqZ3CYAgX/vvmglFc5/fA4sTbfq0R13
VAbZ6Mr0oM1YgtqhC7U9AQBOXT17fQyuDAQzUjnELnm0S1p+V2dSU0K2ynmq3FdorxQXWil1b6wg
ZNyxiTnPc90LojgvluwxIcORQPaU8eAFMzlUG6HDnsnr+tmU0DTpu8byLRRewcqyQMhBP+8oyN8o
lLVF4NbbfJVycpPyTls6DhUs4y6qTN/eRPErsw4r9ejMxW1ewh6cNzB2uJhkJc65SQTSDPt+F0pg
1gunWHIPj7+adkD8JRgoF4k9NUUOOyXAGTOP9cvDKx/v0TTNVoMBscmaYrFVGh1tubJBHEhpakSr
HDoudD9G1GqvOywnvxpCUV6bljYFsAApdqLxVZSnSHhpcr7BRgCgc1WFRs606bjhw44fIQ6vpvkR
+xVwft6V/4tWutD6vj14K20BhvYXpa5h6hG8c10cEUUMWxvQOEU43QLCz6SoiaG0aopJc3Vx5BTa
SXfDN1zekLC+kLyy/DbfrLBp4viiKwOWqvqwQxfCeSR2errihLsUOYS1PTbsJbz15hmZsq+4Zvhi
bTSmXxyHZRWsS4e4JfUjKeuvIGP+4RpFGq0Hmmai0zVqI9y8CbHMpPvoPazfXWAa4jZnXBk7P0li
O53ZqPeuDru7FYYIbtb5M7apQBcVjKH+C+kMvutXY7R9jGsU4qCCTfgEwSlWSdzpPBBvhGUfjHtH
lB1UAAerncB09PuoRyucXukDXvGVYSoFmhF1XFFANgdOM9TxfbAkL/Ff/NyQcRojzk8t4M9Le75V
lxU6MorbEA9h1Ph0MfE5XdOYKzrkYGyK2gLNFUS+G4GwYnYAg8ESH1yaUFIvP2xRVQJMY0zMwalq
egez6AaMPUDtP3XPfYcsEhrCEkR+X5LLelsWSSaa0CKKUWDnPPzNvJIPjsJKNSKsiA1MlnPHR3YQ
i+3Judf1uV2BDMVvGvqDblE7VBHADRetbW42xWL3DpPPhwC0LCLkfFz+J8pN81UvBl13wIxqh0a1
3fvjrUq25Kmge1xTfNI2h1D3yvvOcDgacR61l+llD8EDn90trzpvqwdCTsjKjtiXtNt9lYp7W1oO
Z5fImnub4Y1kTFu3MYZWLlWPQoF6uTMn1yTfAgewQ3VjsJ2XwbcCTtvUnldR2y7hTvVhzAcSDnBM
6Ru9dGfFtdTrePIv0Od1k8OEFSGb2WBcan4Bwtaumc6EvcDhJPOHWZp9sXdYwmnuHaIihcGIo354
ZtHXsLyB3EZQFgAZb0q6eF/6m8DHe+bbI48eGKwxe3YA/Kt4ssLXxgyuJn6Vi7sDQsXlBoib5mZQ
0cxwY6+ly3s06X6lAALMfBHmgBnGKcvx3GaerTGGGQXQS+EN1Pq4jh8GuoSwP+3LnxFOS6iIfIZq
+qAGsrb24GnrjIEpB+wQZnMGqgweNxWw1sOGJjoeEZunfWH61HfFAG/0vWDD/2Rlfgd5RIC5jItb
NIwxmd6ix3eTRZxYBNo8mjBrIbSxv4CS+ytHEukBTKfP/pAtaRkG32Mb03A6sxaGxgtKs+iF5Xgj
35mJuxqh4QMHK3oHi/50Lq/Dmz8g++UMFonhhvHrc3oPxMud+nYlY7wSKUJg3CeqN3mZTa3p+GbH
ZK/emIUMqEBY1/zUgFq9VXLUWhUe0A0+L528zcobQubg6FjgpWobW5GzmF/mMA2Nq4I/8usK7GE7
ECjDoXnIg6nlQgrlqo6movmTJl2DIJI2cUgeI+/ZBQ8UEQOW7pZAe+nmvWKmWLRvq/P5P+JnGlcs
TMtru3XHCdDTUhYKnF0DzUJ19o2+qx1aD+LsynCdIpSxsrERqGjRJYI7u5oADyy2I+NOQZpTR44h
G7iOrjz1G/9wISOPzPzFQp9DnSWv/E2BiopN7tfaA9bqzU/Svt7Pm6ZBYxMHXJwKug4/jNq3vX2o
/mAvk5mc/HFzrUiN+P31CkDcri70H4GcytEY+22vQ6JJQz8DD4fs5ccYM8xLKc0G7nDQ167c+rDF
ULDrynq9Az3ISvFVPoT5f7ee4u44OcKsw2hcWmp96pbtQB4KU295cLh2MiaGx3W8Nn5PZVhLM3Xg
W3rvbfLe55X3QH3NpGRFjl2eYtu5HRfRsbO4zO9R92vwpcabCBDKVWBqnMggR4Odmfu7sbNmGHxY
YJJOcfxdRQduN4EUFStoDQMfpUzgpOKtJKCtr6h10P4aTUmr6vBEqYPkjRX5i5d13YIe9T/ckDh8
q8cCvEHBJMuKzItwjmnEQ8PG11IQsDzsiQxL8ULXuSasGtz9j3HPRihkiW72gEMGznjQ5HLSqKh4
KmtVx0k0OWUA8m6pDOmghA0sNp2mtJICHVtIf8yosm+KbsrzKLK9tkpt0ohr0qE2C0AkGxebTOFJ
p3rbgmacKNVI1wQyb+r4KH7c7HKbBt55S8qEYSq6OTcQJPi6Sqwr3KI42FYPS30r7rqm+ESX5db/
zJeMaP06rFkT0UbQC5LMPaxEmINx+pUfrM4axm2Os1WM6dpMAuPaKKv2j3HKWkY+RXqBcottSLmp
A3rvr+Lx+mcFpV3scbvXrknlJSrValGiszX0dXAfD+PqAlqYVsPyHRbsiUMTshcXleIXi89487e2
1r1EU3jjvzXOauuUMVgv/bFwuT76in7rwVMSnjNGux52C0FoJBYhsdkF7L000MQQ7Hq+MYYk+pHy
aKApAFxoGofnwvvYZt7NVAKLjRZyEcZShKvhb8EKqM2RYFCSKGDSYBeT++b3csAMQmSkUuH7sICm
XAirPX7cKHFa9ICFAFqg9iZtnNDMaJZ0MVUox8db3AmiEGYbHp1ln9dPV8yQ3v628Qh89bV+gZmF
1+Tp3xiBRWiFMg0pHPrFqDFbHHW81g0by8n2i36bCVS90/oGU94qm3u6XhMPk/7NiYoO1Rq1wmbQ
wGFvEAmCHv8fcg5E81l1+zVIKLoFjEPznB3Li0UzLtszH+gvqbZeHxsLiNKDp7HBPKszEAqONC6d
s87aIMsJubQYkZxXCfPqI+kEcULEqrqmu2ul1dZji3MbH7sF82LjflmijVaVnj4BT+QvcFStiAjt
N2cZU0Kvki4Py/i5+Eneqp8wSmALBvI/m38I2AYbzSAIsokAaxeBEGty2CTDGht+VVYddTtM2Y6b
l5oAYlz1WyeqxOogS5u20gOi+XFbSZltvJJByoCJuMa00TWMh+6xgdsdUlu1jaKT/Cih/X1JHw9x
cJjxJ6waKoiWULL23cCEVHjuyyiq7UaNul9HVnWKKIKsnXe6TbAcWpj+c9hkFvfYHErc9HMbzaLr
65d60bAO5JlRMZSfLl/LTV650uDS6ItZflLTo5iANFkktzvEx0wqTfFm6OigBB6rNgN1/JNjCFx8
p/mO/GV0MrWv1ql1ds7R1Slfm7EN31n4RBzzQ/xu9f5OtnYGUOfhD+6eqn0BYWdEm1buMQNjcfNZ
Qnt37N8SS4hVjaR6LJYr6LvFWMSi/fMkBYpX1uvTHoamh/Qh7GZ1nJd+e7z54+/TNi76er2EE64c
+9BQquIUtMSevIzLCfe0v9wiXINOP70UTohJcku6l7tpk4grqIxACyxYGL/kDlqmVfBTzaQ/0dAi
fzfohW+lX9xnDTtmxJXeTyI+pZWzQhFyq8IgJrAt1hqnXq7s5EfjRa2XprcokDqoHb0y24F0B97v
kiHupXlLcGarCTrhyWP9c1/2rmUgiVRCVq1q+k4fHLDPtxaj2vXgXXmcyUYNR96FItt7v31vV4nA
d/aXO2zca6ic9oTqQxOHBBOM425UtVmjKr9gxb6i97GUFNEE3P6+D0uJ3rf7TbPxN0XxSYOhgTxp
VW/8tqQwM+6/BhposEWMkpmNAIrmWta7LGZ8iwoPBSDjnMnpxA9u67s9kw7QNInPBD3gG0fzJ2H5
T23IFWQSi+o/IzWIebTSKv87cdu5oL3ufgYulFxbPWUWTXGG5QuoheWW3682zWMCY2h1j+qG9btY
ACTLuPYboaH9SZqSSDfDPMBrtQbG0IhPeeR274vWb9MEwX2w5Ol5sOIF6Qawee3xMsA4p1fjccZc
17GbqnSZ5HL/3BbkafICPAerN0tImmsv14n5/jNAcryXjoZFH8wdgU+HMOnYvxhWV9hmRB7rvCeS
5ln+3P8X00+FkN5H7DR5LTeul7EU1P7g62oTaSUKXwOyamDEOoRpTsGVaZl3rpo7dWNr4xPGWNet
dwBIR2tJ8N6I2US/hMYpYBpI9ljvvFl6I3qc/ykWMgA2JPWR8tlWXfTpTiFjYZDlUxfs1PKbVKQ+
JbErZIXAuMKWtW241GFCWJwJjFj6yAvRrVvC/Wg2u7WWbYt5ME+6hEs/rd92jNvdTG2FnTc5V3me
jA6GAS85P9dpdM0UqY+ee2iM7XYdztEAgM71e5qt3mMEdyPKPZD0KjM/t+NGpPF14efWgPx9sUFn
GUIfQ6s6U2rLCvfrn63PfIu40sZvv/GlzQsKl4rMif9I+QmLbqfB3z+2hTp9NdxQZC52PvU4FV4a
+2TD72WFO5rBxkxFfRAinIZOZ+tNfygt9TfYhqVyuqnIHuhLNLonpGQE206she7mBexxtx1iDp0K
wZ7GyJOBQOVsjNyvmonNlcJ5Y2VIesxD/QfseV9/Y6UL/Ed5z4bfUEFkZj/dIo521qfHeoRJQ4dm
vBnaGjaztYYypk0LlYy/nzF04kM2MBVMBbgBI3Ke9RFM8zZf/zS0fVsSnu+Ya9P1qJ26TsbDGKql
2onFkwdH4heiBzvar5dE5WUI8ZPLr04Q2CqsP7u+m/qbAoxj9HrYJbFIQCrhbRyyn+jLnrknD1zG
5ku3Sxwi9zltW9uiWK7aBMMX8MMzRYACoucnQdFE9Wjh472WB8tkTPyKgi4Rw42AxOMqCzB7YHIZ
VB2nimen98CWabXXE+KUQP/Oretg1VZ7mXF0iY4FA96VRNL8b9LdZIP88rhKfCc3KVnQF+395aPG
ID2D5MZtrX/VeMLscBZm/KrBb6THCjxeXPVcpjBv0JNQONrliuH/L6dYvliuxVbUFUYLNSgwHgyo
gaa0D23n/aU5sIgUJQj5NgCpw34UgFlODvBMrW2Z2LTdIx+UJrq8qrDOJTVGW91y2nWhipd6k8bX
ZjLNQBHShZwyk/EBVYu++gViVODn/Z87l8+xPfAvbl0pCwJEIvbC0VQU0piZNTRZOTlpHUWFIooa
jzKIpGNJLTA0D6xnrTyVEq7g05Dfg/FcbEiNR5pVWanzYbuYSbxagdVjogYgPPNVzRrtxcX+bRhy
RLs8qhXJHVRHrUK48TeBGPPxO6MSIwBaCCisgqIMiZT2Z8a+OhCmIoL0IEFvQWHgfk2mm3ej4nS6
+f2Dhz1fbs8v9kcJrbjx8D8e9Y8cXGsCtlPRZKo2OkL86eI8ZjbSt7CZEd3FxlDAsliMKQZ1CZmk
3Bbaz3nPXdiPMlzlycAVZ4mxigAnxTC17NkL2wgT+HMMUHwTDVON8/+IJevaFopk2Q+Mj6+9lWpq
JI1EZIhqBOE34b93sU9UJT1aq2Rfx5ofoFIaEWlLLWVQxsJS7UViK5c6uvvBdnuMbMoeaEfzFeFl
aKMIdxSTog+h84ukh3u4areJsGIJ/g0XBRnldxb81Ix0FzeDz4sKQABVm6An2BC7MK1XArhGBQKN
TlEEsBoN5HfQ2H4klbwiwBSX2xvHws0NFw6nIkFB0UZSb1+OX1x2fuEFITLa73gZiLA3gTcbw3nC
jT5V/cw/L8++6JUjX6LCHgg9F4dMgZGGXdrMnTzOnf9iNnNzvy3h+gneoxxdpaFcaffh7HuL16ZR
KgI75z1fkBLIttYMPcdAyJtg9yfZe6MSa6VaQV9OKwK8HgPV8GHhGr8VJM169PkW5m7wvu0JnTvH
CXAq2aK1XVJdklZlkSQFdzm8GTURbXfgDz1UgYkmfLuhqAdzOByOlajQJyP+Su8+Dj+F0vQjNBz3
vw4TblCprQMnWL2Ui7YYhxRPwyl3kCyYJ23ZENr8wIiDCno0Y4vsBloaVnZQgJ5w8xY+fvW7JfNU
uwWw4l2U5R7sO5Cc07lfu5P53sWLB7w8LHLW7fhOKrIzdqZLv0W/yT9AhoOCr9fJLfl9qIymYFPU
gC4sFh7zsj7I8uVEhfsFtQ/nAkWWV5cAN7ULzD7P6KiDE3Od9bEeGQPYN6KBJT0RiJ1DBRGZEbgC
YJ83gKj2LqCRjwz6cRwr2dY7i3vze0fyYQ5pv1gwI+LCViRT+/dGiptYPhh6SWSqWSWpSxoxtCMQ
DthJTunXOjggFXD1DanaLVgtL9PmBuvjkjhPW7vkvtjDzUIUzPKVpj4XFIlg0kuUZoCJuOGfTI+p
NCnY6deLUoxMPL7WihoeoHuval+u5Z0/n5qMbA+5frx3qPRpQn68uoWuC1e6K+BIO9Ep59FlhtjE
cWwCymX/U/xRRoOb/UPSx/mwRLZSRT5mZbvtRfcTJ/wZbxuFfIJbqRi7hxpFl4gu3xVNLTt+0Fu6
Psr+rXLdL5VRQogOI0aas/acE69CpDZ8DXzCCFsZN5wtNxBgnQKWw7hVdWPlW0vAe/dPe5zRcRPs
rAhEYZ/7p5iswU3ZK6eFWO0U+FDEYRaiNjXin/u67NkkkH364vPpChsgrFqxeqI1gIhUwDgj0ZiV
UDbLOVKnI+rxlFhd+FV2vt23QrZoHuT4znpKDayc40e5MLu6zBUs4FxBWqvuI9UyBFDKAvfu4POR
u9Iv38yVodJzVve1eklr4YFrxHcet3IZ2hr30lxu0oJxh+jX3LjuQoEgR2lMviNDrekWtCwmqwbH
/jiugPbeCDtZFh+/c9liOR2TzCZ4g87EhoG8+E2a5+UaNIn3HYW2fTjIhFi+Xt2pxXcYew1yXIsu
N9FAX4Acq+U6gXKOQPxTzDRD3PkSWrHABIM9c9dXGuo4asII2ZN2zWcabs/W/LV1gPBxJZppPvBE
csKJCdDYsftye7UW6iqSOG97slD1gSKwTN6KJYghMy3Sk53rkj1d9EyeHW3Oc0sNTbjxeyFw9jLT
8RaUdeDfop/RpRfnm7BAF11Yefn9VAgcLBPeJgwP1JGSXx1z5MIcewCApVsCddXL3e53JBIXR0Bg
OCM30RlIoASJh/KHZlWg9XdvUXadXp2YVpalBCMJXzAd6uoH9cJSYIxAz/oiYKo5LPhzBdClVUBd
cS9VYfqYPOwWmG8KnnuzH7WvDjwWBuXt2IQ3vahZWf+ebZIoiF1SwD75osHDpk9XsRtqPOasTOTa
lIcqloAf0MXZS2nPtB/vGCfUKCR7ahqHS/k6smsViHUna/jJFF0PsBahDax/5hwhp0V/LBo6EDrx
+AZA0aEm6lCQgUnYeoJAvc1Z4247PKAQbUVeu4jnjSPgBY10Ns2WZ2a31JBA4VtyrhqMfv/h7JMT
BnJTa17YOmdv6nfvpsXowmMa3+VuNbPPfBOJWTxA5IAFqnJnIerx2Z6taAXPDjyVNeLbnfPu+68y
ayBqF3BGIZXb0OmIW4YngpU8WP9pAdMdj/j3mD7/rgQidm/Elmdr8znNtrAvwL7bvRSkYGu+vjxP
RJI56BD+Gsq93vQ9/zh/NLpQcDKV2kif+gKduFxMjy0MVKn3NzJvZfix6GDXJsTKpxq7+V9RWb/v
twEmBxG7NL07XG5qoIIJ3GGtZZ374ylMbhgOgs9l2PboDvLDI7iiKHvmZHrWWSMU48hUACwvKiHl
+xBPCCH246+jUn7zz7Ztl0dyUqO5hlVep65UxWEQQr3DL/cFN2Ywu/yjXoE09sK2yOul99X5/fnp
T7snRvAFZAwjpsqPDfe3K+8liFrs0/HTyAVCKU0AxEWKAqzmbR0eyNUiBgzVNeMSaHUrQBfhqBUi
F4zQbr2VTwudpzaeOGTpS76MAooxrQzf5CdwtfMH+/IoyQhSofb+A5qNoj6CGVFlsQKVHAjjiejf
G5cUBOqwuU6a9aJo220waUsq4UzUf9FGY/jSU+wAzoACisUxhvqIuDa2lDeNIPjHGOJlJ/+CQIXD
4paOXi62BXtsmbOfUO0Jw+qY3adW87dty2/z81e8b7nOPbh8P3FXdofjeIQSIqkRBHuetQK8CNRA
AzHZTexp9s5du4Zd3VKScRfdJSfHZ4889DZnmWGTWBRkZfYljIsasGsGzmkafmqtA0Yh16ADqipX
dd7tVaCfdDYMYxrVzIc4SqfFjykJ5Cdr1YBmQKNa+/KofBglPQBtvKgyjIYIcW9zKG7GDlycZYSi
Vgrrn7vGS/9iRYB33PQQTkbx5mFZN1KxKAMsmzu67niyA2gTMEhFEVnf6vWeoQLCp7itTpDZ109/
F4dOW417tvOhQDClfyzaUy8DS5KZPOkH8tkVQ7PioRh1Btpzo2wkNp55IG+zHj/7asRuxAJncTEM
EifSs0eCms8WIH4W4urJHw48FNDlqKi1AaHhMbHvLjEgN+0EENYRXViTtxvP/Yp1eFSEQacq5yIq
LuTo3gaOG3/kgLEY+dQXZsUYOgmK/dRXH+0KhGGtgxFbt8tDL6vEnhp6j51EmH2re1Q9U+QZYiTU
Yr0wUNQlkfZZBOWsivToSntrjHKD+dYRfbMGLDrN4VwQiaDvoE21g52/8kU0M8teZzVFVhWKIvhs
zQ2H+49JW3DHKDpV91KyIHi2+SjdkxZgu3A0t3yYwwNW49hEodjbMXvUXfPJ2s4dCYXoLNP3Jx7a
LBd0I45tuETy5EIK394HfLQQlvHBXPwqPn2JlCpLkquhok/+znleCO+SzIoX0dGv43NpQp3YU5GX
0stJax7VxRS1gXWZa1fNl6LsQDRkB0s8Fwgv+uZy5U3qYxwweoSVjSRrmVq33JyowIe74oiN5Pq2
yzQGFROMeLm2/RSQMTiVd9p/sQ22XZenVvYKGxHwWsxcSNrhdvkg9TBIf7M2lqQ3OTz/x9UdtjOm
N+a8eKxAJTENuesz5eRr5TCgqkPAs2tuVaNWCYVb5hPuju7dt5+Mmu1nUXJ/pQH8FpoUmijM1iId
ppeJu7aOvYSB+i/T/5FqYBae2gY+BtQMIVprno1Cm4xJaktG6jmsWxzY/WTOlI+12brXUacvzplB
d7gGfuiWsoFpuBCoUaNCcGPCumytxDkCe35DCIf0fPEpPTpMjkW40vFu8xaGkP1Sy63dan1GTjE9
B60pkEFP3+JD5bdg2X9F52pQYLzhFgv6/xwWksrJZJ0zaLhmQJHbNBIEpFQvq2tirvRaM7Ilwy08
N6NnlY7ez4Zk9piKb2bRWQYTQRvzfPsiildftTEDg2s4UoudmNHkdT2XifU0AWX11TakZAEzS4yu
aMVvlFDZagaIWAS/5afzkSoZvlDCn3vROWwsBVDkMl7rdm31dVecqXhaWoWYKwAFnHrC93Sx7gJF
Za9rT+q0lsSNtDHi10bYldSoUEn9Zar0EFjHriImhA7AhwZCI4OJsL9iMMLEwcOUoS4DPafZLUqo
XJkuKQGfhkUlzUdEpiRgK//6hvEw01VMza4j2sZGTfqbYEPc3Qt+KK2YtfshJXjGA9AlYJTd2yUO
S6a0qLplgSzArjFz2gfxvzl2NZrS9g4bx4rJxcYqI6tjAtSsb/2oVcccl3jJVlIElfxS8ptKpA9N
5v7iUEbPl5wKt2DI7x75sLQiXdcrp0ecDwAVyYqObwCiJpkyKkBTJdZFUVzQDjqYmkMJDGUIDv+M
fR8+m4EOkvM8/WT5KXZAdzOqjfmAPM5qSni+mJtgvjbVk8WTpSoFU0m/WUJpepIR/oIaZ7I23HOk
JdaovI2GEIqo2BK8tVtwYkCrlk2bfN/1O2qiRfIAMAZ2NjKPVTkRZrJocB1Z825oydIgeNILhiv5
2Nxk/UEnnBjBCVYSK3G59YbQHhL3TuFe9iHQu7pHxFWVfQPmPq9Tsm8y+uogc3wsxo2L3+E5+qns
1S6OrMr5soBVDpmk+iNqfp51hKzwXoiXK8KRT/Q9xjvJ2hRU6VwfgGV2MOvMSTgEwuaUFORUks+p
cgjTKgV6Hn2Lhw9eaiPbJIRPVZPvWdF5SVTfL3C1kLqJ7s6xQeOfQEFkIW7meMctvvw6MQyYvCuN
5E3ml404qNif7RSsQ+KNJN3izyIVZ13qvF3tJrUT/PXJ/rEDoCGXlTxz6mqQydxQrqvweI+kgPiZ
YvjnTwe9hB2nX072Esos6pUrrgTlDLX4lVV2gJ//bKm79wXPm8zqvm+G4NIwcrJ6qB3Elu+qf/Vx
i3SxfLxW/dJINbyzGbPkKslMjua/TqM1bBNdoyCLxJyN6wfInujuQaE5xtynqu2DXgmQ7rxP1C7p
MR50bBfSQ5Z35MNgtQbvEYf2KiztrRTUuG174S4TCRY2hEKRXgZavRYT2FaTJJVMujKGC8wrLIQ8
6uQAgLAzR9Vyl/FhEBrjBkzOTpOTflN+pZWFubwshNk5zaNMHdrsgM2fD+xG3fYg/gMuDqegEHuj
LBZxBPchPBcAZBoQtT8K6N9FkQ2sPR99BsxINaQs7yXDx38JvFVjNqD2fgoRujHkD4+7bt5CABK9
iC1nW8PWQ9IHBp4uzLpGMwNtfBG03fn/ZEyx74glzKcP+tROvHbHvp78hr6wjst/G9MQ0DtikgKm
JrcrGDnSBwJqwsAMRrVhl90/vFUx41TzJB2O42fbRqL7nu9+ivpAw6boLXeKW3pbpmMYb8oYlNTz
Dv43TbW/SsCWVehMKH0iB1YnMLXUJWyvStvXCPksXPc5nNmtPhK/icx3IuBturppxcP3tLVfrUUU
HlyFkUHaxB6yAs+iat5giCY70/uadIS1somKb6KfCRkzXebZuj0Zj2GAc3pZywuI4Xu1c3vaK6Tj
8EhLQI01j8hyF1qBlEA5bx+fX1xSmUW/xOpUBE6KmcQM/HqVGq8cy+2e9zrGSsMZK6qGr+ZIEZeK
21LN8YFQWCK+uCvBEzM9gF3shat/B6+f7rWgtFm1mRK8GDMMFa/SttnHsD3hd6RTvOcWGbmGqQG8
sjFtOlVWtmtFbUly/+0rvB9SGE/CBJRDJA7k+zDMaYEVmeAeM6UtPGYT9s8fRZuiJmxZfYFrlqoR
EyKWPSBqQrDm8umZoy4SZZnoAV3o88XGjl6hUDDMUo57zOkW3xC9rSSnST0+su9gkHIsMIUmC7Mx
TNnI6AL4cmxa3jGi30Q59+MuPFMloPOnHn2Zah/F7dM0Bbitc/xa0smCpzaID4Q2DozVbAKx+jny
fBZVnEHCrKMBIqYwrnKVNMPnKz50tMbD848LsJtByLdnGqrakWqOGbDn1KkSBHgoe2v436SFhGOm
E2Y05ZHkl9/N8CRvNioQrXsEOQRiV5xB9n8sK/idTo2c7r/BLr7VDGHrKrn4nLLcqAAuC4kJlRsE
SUAsqAXteyQ+dw0iHEy4rCmyYUXcdNv1V9yw3DlmYWqRtZLLm91EG2yvYhMX0gdJ7pXgJ4/nAyTP
bClkFvKv8Zlmg8Fdaq4jrFbBCVh659afSMdYu5h4hdnMhgyh0IInk5Tz96R91N3JcX1NkrQaMS6n
rIBUVbNujX2AJinWjod6fvQT6yzIIGJH++PL7yUUSn2qcvzjluqVb6HFqQ66YAHvWlEIidjzeLNc
IgT9Rj+gABhewolUFtBMo6ZDtTRHouWHbqnRs3MsewUsEoP08PPIMEf1292ZY2LrrbPT1ECcMy43
mSYAXp0oBMuSuCuu0efGDhB/cY8Gi27o/zUlo0rTknGvBTepi2y5vzG447lKuYb+/wlrl9Bzygtg
p3nT8TPU371sRrPIC/leu1GKFJaMhsMvAlGzu5I7mhHqgezIybK90OYd9DbcWBhWYLa0RLaog3xN
gK0zgXsZf6LAWnLf212MBjVXWkc/rrtQiIojgmeNhbUzqB8eg9tWMpjzV4KpzX/IvUoZPh+UH0bm
zPs8SYaaUZ+X6DEb+tPmvVP6NlYExcA9kj9aiRNrQfDm/f4DnPKUY+/8GLBAilKyg92YNs9cCCY4
QA6oasttuX1YxoijQV61Ce5csSaoBUdeV0MbMYS+lrAduGu7S6tsm9LimKMfsEsu60LJBdmuUaYW
6ojHeycZxrTvQjkihz9tkzveFoILN0XUx7Co3HxgYZ/7SL9uqdcXoTJ0prM2kYLT3Gcf2AqnNmtA
L9m2GWx1GmgXPnBA1GcFjHM+xokWmo8c1liFKkElfesBB/U28i7Dd09QZpHfQK11BtJFdcd/1s3e
cD4B/r+CaM7B+bAeDCWXmvLPCRwRaU6N2XH2aTl7szO2/V0Q2MBEEHgIR6v8wzNIaCIVpy7bpeNx
A1in1HMVioBu3UvlHmhzjxW/rSJK3DuSFZ5SvF9z5J6ZhFsxoNe4V0HySV6T9v3qgb2ZAUpEgXBI
7f+qOsVlLnYgeJPe5fjxjh3R3IOfko1g91vdTY6nAC3zyY5/3Vsgh2N8iQuBUOw2vgRthC5yDvj2
I55yKdLgO2F/kt/9dckwDWP+KffAndQRZTG5TLpdusr/YzyKBy3OvLgJtgecC8Y5fna8W/qbgCtF
GsgVmqh80xcMjjFUV7e796YGKrVLVc0/dXcv25LPKcAQIyZq1bkIK9Ycsmzj3LVQBZVtLhxBqsgq
uFVQiLo2IYB4g9aHNeWfVNIYshQpJnmMfdgSbkjINGMr79hsyZIU+jp5BICnGdbzgQWOuhEbok8W
KFoBlkbv4u3jNeoDwFk/aj1ByGzCZnTGD8++7z0C+pDTI2nTlVNj/q32/lXnWblha1FGifHQYplW
NTTP7iZzng1w60J1eLk+zhWUhbqYZeeX8QEdE9BCr3HU6mq24PrDK11L2HC7BdIIZasdtWcyON+7
TarDia42FJeCliXlnDLRwiNv9xWuxTslP+XMPHIDUY56hfYAtffjNF8vJV3n6zPIwODcWbPdOpbO
GmdRiMynPCpWA+0lpMaPlMqPkS+W2iicmRYc/wvf+123dtM1rUNFJ8xx+o6XUpJXV8GIwwIewmuq
6dIbn1d0ZJDb3shngAFOv6JhENK0l9H4rgef5kG3jJ2QL+HaW3+ZtjnAI84jLvc6ync7SnJsMMqj
S9qhChR4FyZt0shzWEoE1H+aVbThfnsKE5z7AgsgW0w0e2TOzSQ/a0z3VuhXOtJF5B8F7H520eE/
xUeH4/xJBM5h7L0a84j3mkSSIjPFVhjshg73rphs+Tm5YbfN31t34YgaJwu/2xZ6SPKyyBrJD7ab
UxuoIkeAl3Y5wDJIgscUt21IVmG0t5NHP/zIJND4oHxWbWtIJJw5iw3nNyIc/rta8+QpMorSZy2l
Bn5kO3ApIwgDhkuAagdASPMQOy0ZcNDVSP9V/uPRrCFS3ZDxqv51TEi4WsmsF9tlPzNok36hnZZg
mwrSHnTqfjQssCEmDPPfcuUNYYV5dAOC+l05UhFIc3NyfaQgcmIJaieu0efIUA75sjjECnxs347X
uit0Pc+eIpwfKX1cmwwrRmkA5SVxN1qRrndtyEcaF2vXZlcWr3LybJ5zzC02lJqoYPNKWi9+ITb6
T1YMwomkLV+IaT67QWafD1A0rGI9sFOUsFwm6zAZtWAz+m0ert38pgfuTTIsi/OPdZbMMZnfqu2A
DyqfIr0WZzoHtWnP/dQiKgT8+7l7QE2p745jMfsEmx/FfKmYYuroopSlmauzBC2CHULWSro0FBQG
HiViVqkC9YqUIeM81ZSiuoAqzMuxmLrgJ/BYSSy8Pf6rbaXwZ9XPGOjUgxLidNoWmVd9Q9AkmG4L
+E1F0w65NRvZcz+kcBpOdXVljLTjK+qk5O4PhEq80NtP90iU0k4wa1s8qxQMlvSRcHV+NDSlwVYu
IvJNac0Psgfz7DWT3ZNgH0ZShZYqyyY7nm/wAloN36lMaaPtMp1rDfnB71a+kX0pVYBxu1IXLGuZ
KHuQ35Tpz3p3CBuhNIRPysCgcv0AU+uHguSbxKUVoKYJvvV5EJN7c/wRleCW/QkHpY88dbnyWPTN
RRLU2UJNEXyKKeE6clc4d3WTsyLUpatAzld967lhOF+udfhw32dTGSmYqfvTAW1938tmIbBAwbmB
DDGZYdWsxDPvw1tkaheHF6aecOTsBsE5GXD13JI5Rsk0NHKspE5XeDtR+cPL1DzBXAV7rDIt0f9h
jGuVm6o693ariuBSKY9hWVU0YcyKwgeNWj04O0o5m0nzb8tPcyakdT3jCphAlUEcHWeYx6QBB3YP
q6wF7YC36qbM4Uh1MPrmCtk8U6/jlxun+SkvmYx+DWdefdtjyS1PS1HLdgZvINUjeLdphg1PSLYV
DMMBIR3cG/pRj+vGor/Y4/4PEHoWtxrx3orAGOhgeESs4JhycJjI+ViAExlv/1J4GdSbXq5MTnJj
sp4VuSGEtrueTD+2uKdlubYxKk0T3GlfXCxQzMhqcbyVCmrIQHwV+UvsyHQ/9npN+o9HnSK2jXIZ
avYpiWjZlrfSDP+vBY6VUAKAl+eTArHg3i2c3FRZ+u638HWuhz+tYN73yN0ugs5i1ZElORVs2G7J
I/EntLIeyYiIPuZQznkTIYv29k+pohueFNiiHJd1JpKaNG+KYe5srkADkoe3KfegZZ1dhNUqHA0G
99scEXmNvTgmKhaoAwCHHx/luQcsSn3KW7vasKzxgjbYddh2F98coQUFNl/8eoMV4jd3NPd1oMIy
AxTfiYpIf0eDB3BQetNcn6no33L1o9MqAZGo94eua7ShcEqn1ttd/wtplKkPRgoVn4XRbR5wsdxr
6m8FNkgqICFaIzWm8Ybhf7xd66VcjUHMXFK4DZAoq1dp6YLiMGfVndhxpof0V14fJ6KQ0uk15E/7
+gompGJWcIpd6lI9fLLBMJm1bcuB8qyxoi7qDQ6JFtnAJAd8Fa9eJGO8+D1QuPRi6ANQWEIkYQgT
svj8kkdsB/9b2KQZ1s0zy55EF7cnHvtMdO5Iwdzzq8hBwE9cPqM2zy85xOmXUou5FWTsL/5cGELC
LONa6M684UkBk7KECAsUb/xwNjnnfrc7bmARXQyEHGicZed+DlBkaQW8CVJOdU+WWTuUMgj813Sc
rZWJICTRqjFwAovV1aDClZ4SCLDeBQjJHmf5F7KfC8aHY9KpQ6K3/80+U721BiavTC3lpI4f7pck
59/9Vnxb73iKaRAJNhjXNIELOQeX4sl1adZ9A9sGTvyakca99+u/5E4FvTZp/yINs60MgdbOwIzm
EN3il4U9l+SdPEioabGg+vq8VFL1/X9jBjLjnVwqinzsGrNLYQ400FglXV0adh8I+If51hyH1DmW
VdElA1cpqTHIYN0heGyOAx6addEAzw9tW2V6lOR23RPEVSaJ5nQqg5M/QOsBa3VH9r2p1BET0HdM
cFzbNR/9857TcZhRkxjEKeVKUhoZoJzrY8xZrn684CuISwPWoy68r8nHDYPbXRCpag/hOP90IazF
RRin7CbUKI0MTCEF1g9tl4rSBF/mDifSSDIP70dz/Ji8W+RvpoNnciVNrA3ANI0hewkcO7UgEzxy
DlJuK+kU5ar28/kUWbjRkIr0jZ8Hf4+G6nC6tNfEa4rsm8uJ/G5gEhzhxcstEZfDbpggLUQEoskq
LERl7S0VoxCTzL13dKQqgZ+1MFsweWWWIx8hujI8/0HPMUUXQc6hgFQV0iRSOWegDWXG7jA84i20
ogZtgvVoCLpVPJhSbrnJOUxL2YgV0+1bKGNcbEFgeEYhNpG2o61RiP0Qrfi6pkXvkpbfDrcIpR3f
s0rHVRbOdYcGuSBiOgC5x9FGva0dSOuxyBRMbCu4LmMc6mp3ObUuff782dngub6SB4yWxbUe+vnr
TdpvMAv068XUL4asUv3dfZ1i7j6l1LCpdYuHQSb0TH2UBLTNVLMSU8VAOKVV2W9GkArNK09UWRtW
ecCfwxxH/ubH87PbfAKC6lI3pTaV8ifzSgREV3LQWcY9i1xfQS98Mc5Z/Btqg3xzsSnEiwqW+JAZ
sKlt93Vv9l4p/0JZXCHa+JzQUl3Bt8Xz56Fi6sSrE5A0PBBtF+s3vO+ypU/6tT78tv9Jyy1C3Bu4
vg2NIcO3hVxa3BbreyuqqaDSAvEd9fjdTH2D+4IJNcCMPqjpCAgNCJ6EdT/7owAMLaiq2fKVqoQq
gNRJNdyTxvgU+397A/W/I0yg2YcO4hlYizgy2wRmO1TavxJMC1Q+Vr6mZVCd0RbSMqetr8AzCoaR
VrHLS5G5Py5H2JmUPm991ifjwIXKeoC2QxF6MI9GdN2E9vdtMOlkpTZs14xqPDFKKO0eOnCyj8mn
xjDjAdU6dYOk4Zl5RLmNmzxNAL0IShOj1VEmvIZiGibngzQHuvNt6sutMxUuiJnC6kvkIBAdO5G9
apRwZGx5Xi1NgdehfB1mHN3emaHJD2v9AWPa/ATV2uqG+vu0xN16TOrsovLj67E2V9gVoine/ysX
CYOjInCW6uxLNsGH7iMM1j43rmA76lQzv3X4g/y9H+bVLlK/rEPZh14rROpTIejFP9hAuOqlXWAh
BNP0EIdWBTIhC5WZai0ylbAe/b7LABepjIlKzy0KuZKC32bynZXz7VGTOSyQpkZWF0p1nSf5xPtY
jiI/IurSSKPGZi9z0FVH0ODV5Z+2PSdRGIzhyllxDdfo0fLYnn5lGSmclty01ydKeI0GIEZBQYN3
bsRyfP+G0rmOxiPqoPAYHmg8NHNsQoJiB2tqP48hw3ESQG+mqpafd2X+emHgvtlPHEKxJnAQ3Mgs
CchLfr1xQ+r1GB6Bs5SuErgZFy9D7yJtiOa4EEL47fxhIokKe4tsx5Rw817Ox/D/ncX0T2FbV2jR
jbmqY2FsOdaC+sohw0SQuTyi41bOvffApx7R0WnltmNo/EvCIKIDok1QW37oCzDFKbLhsGxzzMWD
xKaV01iJR1FxcjnL4/wrkaC3sSdpW1H9Fv/w+WCSlR+rhtLGwKMmRa3tSmQ3h8k95utCnhaG5Ygd
MzTlgTnzwSzbY2gDMI3SNaZwNwCDoO9KlR86xuEWjZ2YmtMb5RxoD+VNKGxVngApUgsttXc0hz3N
fCBPCjUkN7iyHsBAZYeuwCg39SwgFtBjqx2BYVVgnSjOmsfvZz9fn5cykl47d4vlL9C2khEwA54u
ujoi/fzrjlUG0psIxQuwiVnAXxZzTH1gLbeOgNPmn4hwi6Gzs6p04nPL6Bt6Mx6ueiVjFijIqbnf
5dzrNhi0ip2Wqyq8BENj3cnwPHxlI3j3GUhddBeBBAJrDpzxr2tcjws7OWlcxYNz27895ns9hzyV
1BHhdQs8OSC33UwWcFIskv9i49ZXhR0u/xVSG5CfsdRca4nY4WkuKxC2ntnyDkV4F6i5ppMYs+6J
hawp0cWGErznPKeRvH7eLs4cHdMovcqkLQy2oQW6yM31eGZLAkkpAQdzWzs6EldpFjWS6Olm5RR1
UWYTg8SpgIyNGqhZTYi3u1HP04N1JIIWxRZKg6SS5lARZ1rB2oricC2N3MB5vllDlxqdFXV08U6B
WsPmjvvaHWT/VVSDQVq2rr9kmRsQvvyAUUwmpkSKw9XearWsbjl7kg6pSxARjfbcFyyMCKxpq63C
idthnGHcSnMqRe+Xw94fTsV4k/rsfcT7JD5Y8wPuILQjNC50UukDgS5rToTAnGD62xRfBbXXdKbA
dqQSUXFIA9XOGzmY9REiIigtzrSbXcvBPR8Rprzu/49jgbxx5KS2kNK4plC0nvY5WPMeEp5bQkoA
kU7eP8CgH6utsHxJ0nkjsmZJW899T3YwZfdoj4vV7AzZCVvqdy6yqC5/FNzUUfrNP9KpGGDFB13O
y5vsFP32PLJQuUudwyZNetOR+LTBu8Ick2u6wSVNqobvaWHtG94tY/g/Qm3iSYL1XYcPds3VsBbT
gnLMwRdOTc+6XIoH12UV0qrUmwDrlsjsM0Xxv9PJ3Aw336f4y7x+OU6TJZezhFbNl8f4lf1rGctR
rmRGZxR57jLZ1GTb3iIZeR+/2JECCkIlrFgX7bqX77KRVawK/Ytz3/Dy5xqoggrOxnZdDUqUYAdZ
wmhliBOfCqSSTiPqlh8s/XM9S3Z/4UaDJgYSURISkB2ufjROil3wOfWt6IuxXLWZuE2UgdMs3isb
z+s6VCgXC6C6iXJWLAP5QsP1c8xjH+kxKbT2j3g4MtgoiFou8oOY1XlUjZMUBQUCpXDmfd7PgteR
y14gADxbFY8aHUMk6L50peAKKAsP79Q+Cu7svPdIuMbKh1wfkpbt5yE/5bawLhISYPTU8GDl39yr
swhQpx8Dk+YonPBwjIXhRUWzpJTdg4XwfBTq8IGPmy+S4tBZrVL7/fLfsz5EwrLKiIGeTcp+e5/w
xXRtM0BAEGYjxsKsrBeKBQRIXbTLJ/+NgCshI/5pixrp/no7FeITV9Cjgh8WEP96PXDQ3fTmmQsa
bIEBIQIsdi/5DEfdLOlXb6GEHQxEnah3+1I17DZm31LhNd84hVqrNf1bnHgs9S2aHPMPcoypZlJp
rRdQvYm45uVE+VwOvA7iPrW0GHwSr8qtSV1ceQcmfzD39+5v8aVMvjBQbfSUYRU1YbytqbiPu8Ac
9SpTnfCTow6yPcxwdCU8RS0J9PP7WymVtczogxwLEY+tDW/tD8MF5WmBJ1E7DtWdcQY15Jd96BQi
5mJiu9GlS9CKepKG394wxVc0xD0kZ/IVOpibDDd2d10F+wGhuvoovFzCB/B3K/qPtZM5r0X92r4P
F1R43DcVx4Ur53L13yW80P3OVfSXHfXcZ3vGls1THIbp1FBpQL/gxQSFG4lk5Afe/uUizYiOHW/K
DHLwA114+6XEkbbFGnRMwl+qWZhBC8oCymR522sY9H7QelojRXY5j36ZsjskI+lhv9PudDjH2Dpm
TUy4eQgx8UIj4ziFOnH93iemKM4sT8KOuvBdl17tGKZ65F9J4JE7NBl+nBFvYWut7XnyKeRKNWVT
goCVIUSr+ho0hAfUKb41+48DI3jDaiLVzqLRJd0moeWnjuuzEKH5bp+kFBGKVww+nMNYPHtVw208
Q1P4RhOKGzPWShTI5CU3x9A3AfEVBHcgh6ZFodkBofBdZivx5XDPvpnB6fGUSNC76b1s5MfQr+HD
UbfLYyj/W5VqOlcUXjMjdVoy9l4Vdblkhvd7VvsWw+fmcWTnwLU4C1rUl681LOGUNp3oNW6A93Wl
6WTIZuapPsZJXOLVmBRtOs5mCXaxPZrakM0EEkS7X/pZ5bLcTZ5HAdCnPKeCdMgQ2LYnjUaTsm9g
NlGT/EAwSOJMocrqYOj++Q8dp7MZxj1f2FPToD2+bbipoJSBYQbpHQOu0m9Qv5xZ8haKQ+ZA8ZQy
MOFG2g+mhX8sfJoPBmUcPs8NMkDqijrpBILFWlsg4qbOuqavxCGzIF1hXsjHOGNwUcQOHevliRUH
Ysr7x39ZssqUiyvZ50j2IRQEFn6xtUj58ULeulntlw1MqqNkGuXcePlFI0FYFppdClbUHGqORLVp
w3zBPjC1OwpJkmmkF6f/JMy7yJeOWERXlvmERpBCjAsibCOgTnb9L4q4MTQBrNfDyFb4Hcsg1g5T
OBsRV8SO/batja7LZWjegnKSmZUhX28uehxlwPy5CDS+YyPn8/f31/qOxHm2B2Y2tU0M9PjW4mT8
g6+sl9MntqWh+yD0GxMWEsQvun0AwbN+fMUXQ/q7n79wymEUFrEHzR/BtAGAs/so6C5zZVDlNX1Z
PmhQceLPcoyyhw5yQfmuwrvT9DdQXqF2U/+mFpOwsq7AU5w3ng46YW8sPfM3D/BpXXbpqHivU6Au
frWkh5bnsrT5mXJHCoCaWLdGxFv81MLR+H5EIGbOjFlE5YnBAIW6vPItPR/PeRwMUH9MoUnLAKoN
iGLUoEQAX69U87qDM3L3NaXDiXXyANXxfWejUf2s5MLnxJMn5NHaAiRPQ4wd5fO95UcP+iEjdia2
6dTUV066O7Hf0fPG+w6l5uYuVW/YEvQh+OEirRVlu0q3ztiI42Yxu8fYfd+90mlbjK0LEmgKjfBp
h2zimfmngOjPDTHVZl8pjNFwaxmepXfxLLZ9KtfFlrxtAZD/bNdWgOjnE1QST97ISSte7Z3iaM0n
PLtAPOAiwpmw/8XCFZgn1p2MkIlEF67xA2xD+SBylEnETD0y5WdYIpqDmDR+lzfND/smZwbYrs45
gxKu4pO0oQRMygaIirb5Ae1IE0UwuBT7/myb8sKoQImc0pOVn23uA/iaxA2fqxLhmCglv8MyPvF8
wvE29Qtu8qA7Kv0s3jN1H4vC+//C0vKPpg/OhcqLen9FjkbtOkIz41hPrBmscpfb6bvb71QASDcC
Vq69R7LTmtT1L/1jjsIKBIz6VkoPtnNY3xTNMvD108+0NEIx72MxtFMXZiqy9P5Le3c8x29O+XCK
ooIxOaK0aMN2CfxsBHP8OIB3jExwSYhnrPj7TGzWFL2x9u5c3mqmSHbmzac55FeIpSP7eXR/rTDd
1DIsqsdGv9Ghr5smGTH93AqyEANLw5R1YrFq3Fg8EJX2LGT6FOa13IpX+glfWR9TdgTi79LVBGlF
NBR0EbJVi+KFJ5eefo6En7RwfILHgZu6gYmnyOYjymErO4RFD0jeaY90lPLJc9/tfu21lkxITF8D
eMsi323bLthLG1TTHh5ttLNA1d3yS4IHR1US3jmBGHIOAoRet4vGJTsKDaYf8x4cx79Lf5UFF6Nb
7aYJGe2lLUXmItmRuqKTZGpHdzKC/n1YqSiTuKfAWZhQaZJdIoyU0fj2KJJuLofGVyEDM03y+IIH
XULSpZoad1r0yHiTlRWCIB5pbukparof4BJwKO+hJ7+oUMa1JPCM7Jg9WyCyLfeKhVZosgwM1Gkd
OdesBseVNYtN1otcNii1TnhBhlcBahIgfB+wpQrvmp70KgKG5HYiP2lubw93RKd1tmpAS4uHu8Ww
DDFRtzuauCUjkZ8FrFoQwhqhqQRHGLxLjvpf+KgFyaGlGAKeI1oN0Wd6zM02fUsApyyXbGEBeN27
DPs+vJDtnFU0Pa+EaicJOFi9PUgL4EQkcMkJ/4FtnAXbtjexlJbyxSOJSApEVPlcgu100GhJQrS6
Q3/s/aAFsRbF2qkklhU/OXQdOatwvjW777Jj98BlzVvszW4CLdWn7b8rQGkDN5ONj/qGj/pdeOTm
Upb5xCiLo+tH1tQ4g+NOCSHup6+FYmMHpg7kNBjojerqM4V1rWsSeSrgrP2KEx+JwZslh0QKuVxN
JjyEoRMNjAnPj6W7+O9nk3hfGJZEj2ZJlrjeZT/fhiEBw+bw56xjhufNlfsUayUuWMcJ4aTIiEIx
ZZRdS3xjUwGmKSWBayADF6C2a+VnCGGpQ8a4j5PDguFrMspylOq5dyd7Pv4sBQR2SAb87c2w5GkF
T/bEY5MV6sf0N7cFmDQjEJBa1EpQAbPkv3Q5SBuWIgcPy7UWx8vosoTJZYpeTNeCoyo2BF+x1t2k
lWiOcAIx0gwSioBWgHgFeYi8oAknkMNwMCAqk/mqrk/WGm2XMMeH1Q3LeT3CK8Ow+M2D2R80natE
2WD3tzWt1lYUic3tMuMDPmkNrWmTeRCBHkhnut5vdI7Nu2xcja/J8bVjy5uJGIQvCeYXwEddmX0l
TGcMjZKbUxiEryk1Zf7r7tPc04kdCUQ8U71MFDklxki2Y1gIt0Us/QfniipjFoMqgM0egiLl4pjU
53kAs9y+eovjosePCkLQwpWJqYRgh9z8+sJ69gLuJINJayH+Cc1eopAxGtcoT6IHnol4HP7gLu3f
uiw3aSXvhFMYQ4Em9EdNOpvs6ovyfvSGHu9yYVGCdFA43tZSLCKe2rgktcCdEvYuFrYnsASqaEWq
WXTebYC0AxLiCGn2abnGxyOaKLb+mjG0rqBnPQ5FXntSFAGUl/cnvJ8xbPvW8peVnnk2Y934n5y6
aTwTTMBOh+yCWdApQMCLw01kpEdIi+KJb7LWcvCZ7FayEVTEuLexoVj4B69ATJ83n7IRmubxWK1y
DcRQm5bD8MXRxN/s/OTXGkpyPVPWECEk8qIbZshDy+l/RJlGkI38n7OP+4IaOsLiVanXgDMVaNIi
JaQHl67szbcoPl05CCaXvOM5ds5M3Y4Feetn++egrPlii03JhLhAlZpwU0F8KNaYhSg6NbZMQDVZ
YJtY2OoyzO5yjg1boeeLJngT5BPXdTEZKQ36k+6b3S6yrA/PEZsoEkZPRN2zF9YE5ykwUvco0NCY
WofjqNq5yGTDPPHDrXMGEDijrXZ+7omvQ5rVp4IM6eoRfkMvpO1tC4bV5gYw5VBBE8qMbyTyjusm
/DLnJWJFJh0E2y4uu5rHqpJq3tO4PnIwsDI+0GVm1VkeCqE8mAZvjrtm+hWWb6xH+ZnsYQ0+9l9g
MBqJ5mKZ4y/VZamPANvnC4sjxT1YmxtGnZz/q0IqtuNV/oBAhl9GQ6wRGZof9PVN6p5bUHY8IVtt
Jh74Psvz1bfY6M52ZlL31pKYGztgNFTFmsamPNN3vrAgaBJvowEKq26o7mfOZuFzfnAIMA1LEClR
Pm8SUeEwm43GMM0hEs781bnhsxRySOLmP2gTI83JrHS0LVA6+DJqoGIFyeZdHQ4LwX/+OnB8k4n9
6D5ypmrZjBZw9X4v1tpJSLnrkfky7gfs5JIGBLHJ+NxT47nqarwFTplNnEd4mRwWU6HFbC5ewyMT
bbUwBWNjW8NM6LBjrUXm3QLGd0aGthG+0pFwOEeguvxocwP7VKlr7hTMsB34JF5JpdTAc1mboyXC
vyQesbBACp3fY2yxgajl2am1Mc7a9DGmDY3jxr+LEeWUwi+WmJqvjbfRlo1VPGQmqT9ZzFj4Ad0O
eqL7bCVv/cwSKVxQNgYLPJjcKsr+KWjYDAGxJQbSc689ZOenttRfWnfR6Du98l74RI+FfWs8y45b
RkClNHk+qczi1iwTwVlbN7aj9vXkisYz6d2U8Vmes5dag7jIGu0EsNJvilB30FcxH4nA/r996uEv
lqWKak9/nkwcljTzvTpj1MisYi88PQcqOUlzoaBt5wr1XJB16sLfP+7x/nOtrA3uaGM8I4qC/0a2
ZRdjBJuY/r2iQd92CqUct9Vhq261pLZm1LLe9T9pfPevmDDI2x6JJsNOXEMiG5HK/diipIQFO29o
iQOCeGsCceg2EqDmTdf/6cMu9k6ki13j6jSymlkXop+8UhTPaknI21B6dwE85FTjPZJQ7Lkwspjl
BJvaG2joy46wKWcbQd8VZ3B2KrF4VpTuXw5q+oiR+Vv9xd3ZmfB61pEoTdMQX8amYBYHJpz6Wp3i
WcBI2CAQtMM55x6F8cBRZV9XYGD/rKnvHM4kjeivmR4OreNbbBUr8bvSze3uMq4jnJY3d3yoxT18
m5hD/ePnY1xzCYeYGatYzm8GDrz2LS+crUEFP7J6DQK3eCFK7a4S8uPcxvYGd+wfvG7IhWeKag3Z
CoK86TdUbe/s5K33Fou28ANJ7mzM6tRneB6mBSGVk0vw0m0HUEME9QTVo1HPUeC2E4kJIUyCTAHM
OG31whFSgj8mSizWiklbs+1MpLYzdYbE2ZhIm/qsSxArtGnxWY5kkOSbWrg0WasR0lLSkWOw8kOc
hRc4MYA7GCPP28oCUhMmhGV6F7vWhHJuxYfqilfHucOdqv7dzaWV9kwoGcG5Vl0xND47fnIT06VX
Er33lhk+mdElGunEZkPKpCqU71Srj2TP9G4+w/kp+xwwn2Zoxn49kMl++/5+DH4gUatJvnoqYv6e
lI8nYhr+UwsOqOhebhSPSl3ffyVdqSOCudXDvf5TIojLPh/I5nsHn1TXsc5WCT6CRL2PVAw9yuXs
aHzrcwAjNcSK8pGbA/jbMlmY8nKuieznQiOmdHkMOidIs9uRjgBdK1b3gFXMMh2QX7ZkH6J5RxoW
X+ERMiCbv3KcPNIhn2nuqFKd7OT4Nk8Su85j/k/3Kr3ExjbXw0+19secA1I+lJBQM8sqT7WIYh88
UwU77+FKkAK2Kfb+NfM2jOiY6ti2mw8IbItMA1xq1LT5+ERYlU0JWsyee23AU5x4dcS0bXJYRcOc
dcKZ3Z99PZjBpMHUQhdkTeEUMyVsS+iwMGMXcpQCysZv7fgbpO9ECJze7acQSIm9gUR/nGb1zcQ6
51+HwRzicezFlZFr/CZtX5CY842KmCClDdYkg3M8sVywsAS0obAUydwHEV2Zxflp8YoPLwXyhQWA
/Aqr9iXOd71jd6hbG+gFYpLJVbZ+JfxPHTxgLBPszSYgV0FlpQhjQCh4U8luARIOAfh7PhIvGNVx
wleNrvgKEMaKIfGerW4VeE2BWgIvCZmW/juoH493LJm3nZunq4wy/v+ZidBA7EQiKe/8nLndedKG
kMPemYvJo9Dd9NXmB214Wo+1A68hJZsWRV6uWLkxE27Zh6SOolajyijteYcgzCykaz7Q2kpefR4n
+Yw1PMrdbevwCV3YlU1SPgqqnWK89V1qxDLj9Ov1IzxcNMSPRcVjN40Ua4Asj3qKS+8hSYgKgz7u
ahx7PlOhUpxLlxCbHo27J2MjHOK8p0/n5HJ/E252on0xd8O9wNaCxn1FLqQGgPWKGlvQb0SdzE7g
jydIDstWoe+RSrZpmzH1ce4pq/6lnXPux2FJtn3qNaFlMqJKaShCZNHlfA2vh4q1zZYCVkcFzt1n
maYTjbsO7XTwuFc2GRdcCNReq0Rg+FcBw1cjBDCyyZAW+6szL+Y9gRB64iHIXx6V4gxDK9ME91WB
mT6ZqncTIXZV8hckLLYOMT7XWMJ0vbLlT0bOqQpnLnmO7jHPk017/RcvR/jGfjwcdDRAJDWwjgUC
m8gjeqQVQTg+bgR6Rf+J6tZ4NP2STlEGTIVnQrTUmWMHJeaLfyWHxfZQM1mZF7+X7CBV//xRVSAl
jSToKesrjL4BiQiL44mnXBbz5rV3SVfDDusFHtr2q5QEleWwyW0UDzjOBLZ2Rh8QH82eFCox5PET
JIc029q5ChMKlU73oB4QhaGugGyBd4V87VtyasdrPpWcU/PvJcw4AE00A2bQSs25k3pMGqN4xpof
r1HJApQVxllOFqTXoHeWEUlrH2lEd9Un2wTYeaRRywn30Tn3MtKrVxraIotrl5O84KfAKgocM9jo
7hhgA+bQUJUeF8SG8W80lEq82eJdZE/mC1DP4BdX+Tb+aSo+2iPwnc9Fll7d+xDET/Yo4vRUYzno
tYB1i61e4ijDCSt7afy9wc2MgkhlBTpQurAh4qu+qRMjuV0Nnb519KyVNuDYLALGsbguuUmZeO1X
x7iAU7tQ09DUdl22TF4f2L3Ivs+4OGirFxYDbOMAhJY6qHgD49lloLW+/8D0bTGn6HQKiY/EJpsz
OmaE70rGMNtrrhbSSSy34mB8T412ZMIJuTBDVOq1PpaekGlEH6qIa1BCQbb/KBjANWLvtGz6NPgD
d0CRzzOmlD5SQGX3raRKfc4noaQSNiF3BB9hkhZpBHbUgd6NiHVFD5N5bhtDoO/sKjTOLjhRmSaH
JDUklsM28JCmBnJxIgqO9puhAOPOxwrF9qpOT9Piiyx1bttAqd8+wnRznKZlrifOqQwBGQPiYdhE
Wd+xkicpzcHFEMh9NS/L4pT+IPYp94+nywwgAnq+uZ90IZpEabtc63GMICE6GeZ0vLOnUQD+wVnM
iTCS9R8d3YumJ61V/rLZjyEhQ/CedI9uLO7wdvK6i2v6ndkuUOfpkrG/JkmVKvrepHrrA7peI+F3
Ye1T0RSdPDaGgjgY1No7MGIJBTFeVs2B/1AoyTPUn+LIQAAqOzWsZ3rjbr/wbJSlzQqhFEDoSCy/
NHwUL0+d/3VaeUst9d8qHpJRJ6jExOGIpXL2PBvzLSNDNGY8yqIhXhywhRT0DkCoRxCHBftt6PoD
/XUOnqtntZxJ/bvO4hW9WxMazK53Z9A4Lt/nxdHb9seo7gOK9P/x181nLSsCf3HxGYOu39aq44kb
nELY0rT0OAJqrEdCTbqFyDbG3nFbtFEyGnGljd8ZU25OJztkzXBoI/YUVzYe2SqLrNSgVmn8Z8La
0YXHE8zayE3fZ8qSv1C0toi+JStGWcKlpFntr1AzGhbjorRD5uDedcP0XgVj7QH02hp5sOkKK2EA
xYEcgOi1saFRDZ+68SbuvxJ1olhSrq2mSXHrlsOxFpucyAg53vFZLoFIamMEf/XvN7KREV9VyPl4
NzJFYAG16l0IVbwhD/EMj08NGpqrjJVKdUiKM/9ja6iDML060YOw+497ad1N2zsvy0s5/c5A8dmC
MknmasUG9b1BwMmJhSPNYwbGhkFrbOnq+PA17SuAcdKN7YXtijsyqlnUUUSYApjgPjQMMzNvAdFw
4E03XmGUf7pwdzFaQSFM0ZRmQ1uAlZqJ+8wHOjOfFg38COJyqTOw2f+hbHVDNjafo7ZMljAAJlGH
WiK3wG3SoFEzdWdzrlSTDmpRdY3OWURm21sDoZU3faKDbxRE93KfCr4uY3Yx2bbJ5okWZh5gq1bu
mDRtshrgRN4WOj85imn6rJ8WB0Um+TBHsZY+OkzmyEHCFYcyb5VmsExoUvUYynRvUQzt1DcFdXvA
HGbZxsck1eVcpeL+NIqsiDqCuPiou7D8yvBgVTBhIaWbJQ9voEAEaz6+MwGkvoq0hrZJjvO5icRj
dGYito1f4LUAjEV/GfjaJzbPCKdENyVYY7x4ELo1ZTSxLlceoI87xqVgBcPoBqQ8QBS1SjPDpo/D
W7HIZgdZo2vGU3JpdMnMfjKt3s085Mxk/ot7/Oc2xiSr9fcYPpR3y3vHJ4xl5h5z0/eK2R3IOvOX
LKc5YPUv4G450FpKP8iKrnVnRa17iDVHZdGXS3UtafY5B6p3K/G64iB1chExVc14mPU4W/CpPUnP
5snjjkrdYnwdZ4+9dNRXHV6wPOF0FGj6b20nuAPejumzbIBpBRASzPB+o8Vcnl4uORAYWhjjMZ3V
DhLMlY/1s7wb0b+R8onnNc3OhYZlvU2qCkQwQiv7R18wvMl1XDkY258Bn3f3DJE0aUR/bPRUIKN2
y5jcuPvRKZnuthULm3AW6Shg1EDD7JNgYJcsHPM/DShCEUdhimdLWIzXn27tdCFZou5TkRDnxCyM
FtRbXbVHvsMd2b0y8rUza5OtR/EXSP45Q2dU2k25XLSDXENzmsO5m2sZ+XQhCUimFp3W64i2w2Ke
u9vq0oVFFwqkSoHmM2Pnlf9zHlK5NjKYsU8VacRQaqeD+z3ptSs+6vkyL4befnMw9cA68cQxtlTN
xpai36peU6kGPQS/KAtmPORml0kZ/8V1co/ys1tq34Y07vXPo865zuFfpsyry/Eg4qkud5u+Bh0B
6RmtersHV1gr0A1u4g2YHKOwRZYts2usb6v5Lb2Ed8CwbdjV5CWqD8BMGke4WvHLfdfcWB4yqCt1
dOAKiaF6gL2jHxmhgeieWzyGvvnx7OBNTvyoheMYZp9HQeVknLieIdFvGdJwwQ0VFbKLPByNtcRS
NHq8pIKIFskUN+0pJAWru5nTSqRNMmHelsFDb1Kji2+tvmsxR77+9DOYIgM+jaWkCi+KzI9P2wpa
p+nBi6e/xhgKwyPv4ooRrw1R9fYyqPrgjcfLyvR/TTdLT6E0vTCecgjHfW6lzvJmdLy8R41lcxQw
NCejF2B+1+F6cj2isgN75oIbtSGJ2LPcFcfSH9sOR+A0LSpjIQugi9IpatuUDeEtpGzBwlFwJsmH
eUAfAiioGNuZ/WQSYWG+O2/x7gR8h3dt9H9PrQeh/RDvFfqcaqqrCOVH5XlxCV86K1dP7zX5x+ku
Yv+zz1SIkOAWIrCpCTSwl31nekU4yhrDDKN1iidyTbnB2yPBeAfAwVpFJOYPe4qFmgSFAJoO73uW
Uj/Qfaj+E9XgofTVpPWETwPb//rvR48h6cabn2wiYp0UvwjJJyAnaYyk9Y6WDut/e2ExBXogQbCB
C1Wu7aIRSgqzwsRRhv2TqfRD5XBSyXjachJ9w7VcSI48q+fLiqWgyBtA/i2yWcQyh0a5JDLis0n0
gHzdflaul90oX7NRWAwWgqeV4nGAh3NUIYSt0OsBNHrSqEXn+OYUmyoiPrO1p5+LLd3CQncktjzW
PxPSGJXJN82hb0VOBb2R7tZnxvcYucv99pww0e+yR/Faj9shZB0r/Qn5JwEmDVzCvUuDfi5pqZvs
vMtocfbejLUT8lMpYUF5/vp3zCDABEinh9WCeOhXYvvjjwo3waoYGFUZpyiEjgz19DJtkh4cyMoR
IGrkWiso8InT3/E0q1C6k5w5T4uYzm20hdC0prlxprR1AFF9sdb9/97EEM31VdsNp5XJuJKATU1B
X3ut/7EynrkWNFTk2rRPJLRNNt3Mm12kDKwk0/w1KXNvFH+v0hbtgE5iAcDnN8ssdqipH05U/Yga
Nr05awajMXUCI/VKA5/9Mjr5c036MFx3vz8Lrf5b9pme0MWCqV7pES8JAqTc88yKZjgWI7IqQdn/
IBqDaxYu37pvRRKYQKDO95Dr/0fHdznA1MlP1x6kqaAHSlx4FngAsQVa9ZOE+fbnuRFajFFs5FZb
CY4CnBfEFjS+NNamVyyybKu4gwuYi7NsttvYTyezd7YXjIKfwYskrE3OXcNEXJUCyEV1r4OELel0
gN9Fhymq+8uPSfL+oQa7bDed1O3QCFuCU85vZzlppOzlvFV56WfzlY9boxuPz7qB0H/NjcNBI0Tx
FBaUhA0bJfEVdZpPu4x5KJi8EtvmfiT1q8GHIHwZdq5JvH5jozlPrbs3t3sUN5NRzxgX4RS15gqh
Rj1iKoZPgfbGJZ+Qnm51UjVsaA/XaN3SDf+TrFlpNBVQIXJnuHCEunLgYAdpYMZdNBCk5q14Nuev
AvC24fBWJdfGq8xvlIvsu8opG05OYADUesOGOP5208rNqD19V3pq5OLZYvYEUzg2aW+RQz39ypQX
oUw36ynDsrbR1zGBlxlhcJm5L6DBHqo4PJs8G69WjBOiFo+rvBBVV2gdsa91upF2eNZRjK8cPtwW
0dHSeMiX1qPnq2q1x3ED1BXbWybkIByxsspyYvHV/UwaCz7bCelT58+fDfR5ibGU00ggeC71WjcE
teJebHIZ1YJ3RI3kPLlrwZcsSMkn8LzYmU8THceQUMQWp9zJMAt4n/tN7JSyaEjYHdaELOjell5A
I6TmSlzYa/dm6kgKpw+8vzrA91W9nvM6tiKwn+n9cfwbK1e+aYs17n46KDArzLRRLeHzIMtuHNpf
subfEXvJu9InBekH/HC33GAssaaAgjUl2GEiWcsHp2vo8TDmcpeccIg0sqz6cIaRqrk+yumrwcRL
DmbKkGgUnKGaww/Q941j7fPkN6oqve00qxylt9wODMoEaCu1hNdNChm5AVdhzQq5Dn1KSk4HcveW
KPC+s3AhFaBAHk1eqOV8Q6DDCZxGKLILsKGKIj9untJv7OZ9sJGwetHjjCfmtvOVssQ81DqujY0L
3B7YClJxyomw3f6vlUGzNKZJQ8w+Ro4gynN293KU5UeJeCbp9/MHF35GmQY8YPI81obckxpluBWn
s8JUnLQqYXT/sJMPK+MS/lwnSVi93y6MC7N6VWiAk6dHZKGghesFSxHT1pJq9v+7YPc90RjGKvaN
40G+fnFq2CSb4QLVjFLJnwP/BpEFxBdUO6ucl4ZgNRoeswsb6loQArHN52VO0BnYPqpYdwdfR4el
6zMRCDP1QKrfBz6khQiaTE8vlE7/JxOGu/hFAEXcIwlyr7wC6ZhwL/ojplFulaG8aXIvsRFpWtkD
Z6uorzFU0F3DeFH6UWZZcm00QPjivwC3fyIUarbVY0Z04Pm3MRDHYDHjQEVgxL8QzvzUvND4suVJ
NDKE4RBcxwo9u8VVHkT+zjsEHaYczuaveAbEITI9qEbTS7XcqN5l/qLTVqZUxHYDKHcJz5S4ej5O
88rWxFtwIcoA+SVAWG7DML5bDKlo3FlVDhMmxaBIuP3tOqkKxocpWCA3+T9e2kFuPVHS1Mick+UM
PvkTznmkHzHonND3XHTlL9bPKyY2jMhsi89v74JxTt/RCKfXIua80u6KCVQ2AEgMAXJeAMk7hwGG
eoFgvKyA2k5j14/T6A2PNUL4WMRAHM+DbcOhG06KMMEzk7P18AHPxOZj886Qmd9gZtKvQLwp1NoZ
O+MnSjmUm+tWFydLlEX4nk6Ow0JrbzZcV8sKgM5dZDki9J184/RvAZ2DF7DryO7E7H3ivHJL1BmR
RqAM13pcyMPxwsnF6Cl7/4QaloEu+y/pn+uEc/QCkn5sVG0Svw6a4yDNVfT5PNxX2lW8Ynkm1rjc
kM8kblHx507tqIgQaH02nnWEfR1Fr1sb9m8LkfU9GEf1Lz2xIci1zcH4cXg8aTdCr3vVr9Dkqfv8
IXdQVy1bkW3IFMyXt14qeV3a7UeZon3Cgx/f6khXoMAXxJ233KbFgUQ/cbBe65L8pzySECg26QUF
LzVG2ZztjgkbZxdiO/t+91aGu9a+N++DP7e4ByDESA0DmvbCWjfXZKGGdbb92ZWxcaN1ZP/Xx/Gg
l58j2jkUQX+oBdnyKqQlhdqlcgXYOwRgRvxH1XgI/KVC88sbjEJ4hc90ermORoAIttl2LNvwH3eI
Ac+dK0uclw/dc/C/hybho3mH3OquGHFQTCXXWDTruT6Ys4hmC2N4jW4bi+Ol+RcwHLqSNUdKyGS1
jnCCLaQvUncquiDOE3WwCxMv+0md23vipGizS/LWNWmKU3t9H2H3FsXq3liH1Q5ZcFQMX3P2bjvF
5FWsRdVz6K/utoMNZ69F6PUjVvrMs2vBcJL6L3nt4T0M8hcIrc0NPvpYjbYgvWwxrCQROsEIxGUV
plq2goXk4ZsnFk6n0Xx/o1YcvOpQI4l6QCq75FJptMOoNmpZtfaDTZo/FlNCqLsT1HQbXrBhjKGa
CyMdS8vVvWCGaeOEKMUovLdI4UyoTMJp9XRjnMdMDmaoK89gyb/jO67LZ1S1shIJFMu/4YfdsVL5
VlwHWyTBSClXXGrEZMU/Elh17pRQCNLTyVgZjgJuZw1RYlaqBf0RMSHbiEVtdITJe+mX4O0tCGA/
cM/rsP+smEZYl5gIms1JOXffRsTUEfzDFguQ4tUCUMCZ0YKY+gZhS8/XK5Jpuic7ufyAAJqpkrbi
q4JFrGxf07oQLTlVYvSvzHfvBtbxLbeMG7ed/91gl6iw8RLbggs/XPf3HTW6po6WtUQFl7VCOVef
wohscZLcWKKf5WAqkYt4NbVM/59VNdflv1h03hzgkCSQvjTwpxs7qsRloVub2tGQArZsF6G1Beb3
STyMgzXuuQVa+IyKl+to01VWGeXFuYiukKpxZ9f8qKTaNNusHZUTODdwvsX9gVGzvq/0X/y5Ysla
zO+FOTyUvASs8DLGX/bfW7EiVY188lZyPr0pYJG/Gw+zDuDm6yxm91EuoAu3UExVYDtyIyvv25Av
DQU3a/jsovUjKcyb5Os93x9B/SepU575sTaagF6kV39jtR3GMJHObMG862bnwlCaQ3MqID+bnoej
nglUggOPaRzBcXtN3HN4EugvntwBC/TKHQ1q/iwzj2hUwerPb35pJ/+1AJYHtXjFxs7JoBE8XyFb
K2YOxVFiW7azcGFq2Lfx6FmFT+e/cW3XxywFlpIbYVCN7oHij0cRu/pL1hA7+KmEdaDNuguyC7w7
f9grN9tsxluc4Vci2W3Gf/dsXwuD97dfwOVlROTLaW6igvMliS0cV5797L72rdtsweR/aO4lx9jB
Lt+X+Gr5icQB25GxAWnjiDdKJQR9JWiHHmpmT6rh91s+avHXjpPfym5sgsPPNvSThdx6LFY8NYtn
a3+hA/8ESCI2FscAxN3tf8ZUAXG45MWtboiIPM2I9RcAN5EmxIdO1xE41QHFZzFxs6ShkhyIAset
es8rHVLxWRF3WGsQZTxCBTOPGesNIiYSEg9ZEDM6Zlbe4NcgZ4ODBucIOhtnm3uBfszZ1hpx18jF
C4kvGrpm3KhJjJCmUmq2aRKa3QSfmkt8zhul/hSW25iJ3hoTugbO8UAaG7diiF4JWeGfw7R8Plws
9RB5oLK8GZmrDvKyKSj5R9ieLbcr87dwhk4hGM+//L+JAQXNVd+LnWIplkgsRPo9BCI57qEtyduK
ICT8itFPQWLFeyZ29dIXfdP2jvWUqqi9rAy2jC8XaOoZYfB38i2HPd7quCTa+8QdrX2Nnp1u5Kcz
YJ7GGlexTrKHLOxhrhY+/z7lQQ3u+AB2KhyjezyG7CYk+7MpuJVP6Ci86PKAO5f72E7klC0g8CNX
U0wrMhdKLSKb9SPOOnjcoLNE9FJCt0rTAQXIMyY0waIf+Ro0Sj958e4Sl/O4dKMk8zkf27cj2pCh
92fhKAdpxEoq4ZqCzqyD0OVGUvHCNTetQXuNJ9kkZze7Z9BtomdiLT0o64KFDNxV3LAaadDT8jYi
CTcJDoXDrKHAnd+UB32uej6QTkNKbQxHL2OcXIgqiy0WTSSQaeMr6n9Gr0E/KlH56RK/Gj2zApyG
g9YkGWQZUzRmID453lRNx8WUbVa2uKjk6vnI8EajTpeN9eza9Jtt8wEMOiUR3U4B1+vS4qjhBSwX
5FKfwvSxQnflsRgMskhdkbzl/iIjSZSaFvdG3AH+3eP7NezS3CVX+wl9ctw7+UsO6K4c7AZt3jqp
vYFrkb1qUzyggnHlub/w2DMpt7qdD0Vl9JewCs0yc3RlkpWDVOKD+vqxz+GoMPhpZRBuT6e3fyaW
yRib/G/qd6dotf02D/HYrzI7D0iKixh7xSiC134nAR3uhD5Dm6br3Qa6zPRpPGoyqPKXS9dwOJom
dqZ2e7bhfDRyYvC+s1ej4yV1QekZuNwwfxM9kEnsYMwb0GPfhO8TbJ7b7Le+6l7icLhE64pK9lF6
N9bf5G1byQ2Plu4kd6DOP0nwPILh56hR8gMaH5T+lk43Jaqr1hLs6LX897znv9/+tRLGJflQGxfx
GUPxdX0EsMIVHHL0/N+DDrewZWkrj/W/ywMafzqznAgvcURwJppnXrdHn4t5wgIxu87B0lOix2Oa
gYbnVwI235+8xOKUntrH8GD8tU2e6ehs9NFanaxC4SPwBJZb9i+AqzIQd5aw7ub8y4++qjMj8FCK
lb45SCB9T30cUesY40m5GVHM4Ays95DbvrvZB7guDbHHOATrtfC90W3N03fz9IupGGfqePDlbN59
H5FjohpuqKVSvH7hpkLTe5wlxirxsbCoEDn2s9izVQvpiNudhWHGFtRePIUaAzE2nus+ZM8tNgmO
UQ1Y2id4/15uKnIG0V5CBXkMaGyNMyOCLZmS+TWR1lUIhKs5rw9JaQWcSb4DqdjMQd7lzeEwapy5
lhMZ9NaPw4nOh22zXJI+gi7Td8xxxorSaU7+oTKadnsF9VEQEc6+5IJjx5khmDqk62NxrSssB5XE
SGwYpzvEQ2Qr3YZ4eXIQRdapeuERIGsVXhzZi57SJHp5ql4d1V1onNp7YaXn+bmqgOak6DVOJWpb
kA5hKEPRvCp0ja5XnkN/0oPAG8zqJgfezWyu/0hCV9OW1SwA03cPyw6meuZqI9x/V05Z+TVESdax
KIMw8xJ6esuzb0+MRVzldZQT4oIuB2ZBkbG9t7lSF/7yXgZiJfjpIjVgKVx+9Qzc+FDxzUXl8dcV
GVf73rZAmf3LX8gmCCpnmYICnJgYge22XJN6UNEjsWY6w5x7wQILQQOKG3HpQmkDT+blxeCQd1qs
frWext5XoFCutEqqiQ8qUj+ZlNrJLYELnN6LLfA8f/XY+6csxqai/R8kvlLeXVUFFpRq52f5ypU+
8B87RvOWBXlwFV9D0H8Yg5JtvlD4/cp0PtWxfKWmlA2DqYHBRvbnLAeEpjhxt+T1XIyLzhhLUhXw
z3Cz5kmdGG6xvAtHnPU4iBJNPdOR4um4iny28hlBPk/xrCACHnezqxmq9GuwfAwaaa6XOL03w+GA
eZNVhOb0q7dnUtaRYa4deo0EspL5Yh7HJYiVMu3J4bYu9i0kuo6yyUXR7/zE4C7TeFLY9sV/9G5m
txsf6WXebPmSY3S3uBT9YnfkqeUWFO2pA4TIFWFh0DBQycOcQP3Q8ChnIsmC87QupTQYdDcXx80M
va138tP2Ded5dlfXcAev+DG6ZgpKOBGF8kqivk5/VBgEC7TR00w167ZeygjxoW5KRNsmb6ud+0Jj
qv8aM30QKPyMuEu7dNkHAqjvyvsPxtW5QJuLg0u+GrzctlU/NSZCFDFs+g/i2D9e5yq/ghsVw6MQ
wu6vAiUL3rsXSXn/aNIGa8oRV52SZ1wc09FLCCzTvwzqjs2prYM/2z/ZFtVrMWtVM0nWIs5JJp8C
3Z8DdrTOwVflRXxy6u8fqXda+UY5gbOwVaaReKs/GnvShzAXADSjRPhoVz1KO+beKRV9eIxn6sGu
CBj+oDG/DgxMh/XiOu7gURnqFxbR/PGg7IqV4rep173h1GuKyn9ZHgeg3BHVlGITkmndDvOeWbf7
bZ07Sz9wfb/SlOTBhlk8Ga5dk2G0sv7U4C0sDUwc5eRlKFe+bFvPQW9Jn1VCD2NSilG+44RRA56o
LkbtU1DfsEfQjJK5sfw9+kHLh0flp71IiepAJ/ETzkexHQRXNC5xSgXQo1CTrcJMTu3Rw7aP4mJ7
3dSPqyOyNTkLQUoZ7RM8Ng8yjRptsd7Xu8i6ECOOKQwfZ+vGHei8stspIaediSXKCJsJwpccG+Dv
TUy/wR4ncrGzQlw4J4nVwHpENoumrlC1COdbtqWM4cAdS3fkAWCLbuTC5+MzxjLeWEgzR1aihKOO
14GP6xnd2SnWZR2kBtfBF7g9Hyd2lkMTY6KYFFwjCdfbwQjgEXxX6rNQRtjU50VtRNaK0fyeYpKL
kSZBFhnOBSVRnYgfl5Zn+1OeW0VIYJcWNtprqVMlQOCAhviz9ex4/ysp9jlFj5qWrKkKck8/s5FS
nlIS9fzVGMLQS/puqpVyBgd/FAM8yXbYESFJnJA5vx6WKE13j/Tdc8iP3ouXpzmGaMo0XNMqyEuB
7EGicj4AWGlg1oHioRs3QK17jodQwZIz4mozoeT31KvsqpDeIFI0uMlbcvGHNAHYKvnRMzA///tB
LDdRH/kJGMQn9PM6SCM3gv8kZ+bPlUdlhW3OT6VKshEl/fBzZIAlddrEPTHzun7WpQ0Ev8hLIto5
INSxOmjjmrW1QpLZxnJI4ODTkhP3iFl1GNuZ82eMHc5/xJTRgbJ/wYUU0SZeM496ZDhJg42sum8l
b3LlT0G56Ky8kFqGv61EIpab2NGukWdxZK+Y4N61kbgRrEYG4uCa2wlnnM2BCViLGTp+9j1VGoCn
ETfyCsYWHPfucxjQ7ozEGrDMGpdP56xnCRoj0dDBct2JzJePFe5hK1yBu2xl9g/1sj9mymc1UPkF
51a2/elI5zQWsM+xcCJxzxVnjBtDutYMJ3aAFjElP7rtFpYeOP5XPU/vK6VZBHRrUKCP9mcSBs/t
UsJUiX/QnMbXtTEXCxc4ohKvMr9YZBpJoOqrdKLdBZA6xqFsOL6K3CNoarwYBFophxh3Xfp8w4MX
laQAeZhkR4eNVc5FCISGDBHYkwlsawb41z4acAgBTho1QObe3RRD8HbDVdNgHE1eXDJ7TkLlVH6Y
0q8ZbS8STTWeQ3nqvoNodTNICm5wlgvRKthMPqCgXxDzrgwILlgt7nORFBhxo/IDihoftwCKTCOc
NQnP4/9GczyWMQrtgTKo6g9ScFbfpDIShCqXtu2Zh7h7HU39mrpWRkfz9fHxJZAd9VcVvkMkgBe3
+IibEnR+2R2yTMGY3BxRJw6k5p2bhSyiJ3w/F0Gvhc+lSAVfxoKibH17ipGc+rhrNi1sxqqf0Nnq
IvNcjwCPpMTDB9m+qkHcNFEbbgUtwUKleWc28I82eY36xLHNzbK7/R0eOMDfGmNXc+DaLacZ9IG1
C9RaDiVXK4O/gPZkq/risOdhJjwZlYimxijRRXyOXhh8jLj2F4ONO/WJIIhlxJ+g4gw2uD6usuOS
Eu1PEU7Ll8thMgWIYdHvup8Kc30v7Hq3abBaKUEpN/bDlNupECQp6gtiCKWzM8mm2KyJtATFGdN/
rVdfS5Qwg9YYIH5+G+rniLk/kg+9n2q+4T10xlF/4PywIOWSx3W8UzErtbR88dWgBoYFUANRdPdC
ZqVBlh34RKEDIuW3qqgqEIH7b7ilyNWrdI5KpJU2eiT6YmaWytI7XKCgWyXxhaXk8u0FXtY5FXP/
P3/R6/UEE21iftjX1NCLqKaWDcnX6ehuydNSYzAzQWFd1rJXYNPW0xs7umgKEV9yyf/mhYpEYXTs
VZ015+PVTWCla7LhD+6GLDf2o89DF8HaQOpvuDdbzhV3cKmUcXf0bocd5xWKTW1miUhCUaW9lbZi
7927oHBiU44lWBdS8WlJuGj7JPPEL9DJYBD2ubHtLJK7xC9ay52bzg8nJMSFSgqlvwa6fLnmoFtr
jy4snHJ3NOdMlnRhgNcjfZoUwH8rBJRKOLM40GnaP/WVE+Xd3dmlWd9lTZxmgPyOsSqAk+aKrWKq
0/b3ygU1PHRpyiBiVGeiyBIMpCO4silSX+ILgofcJPTx2Q/WmowAwQz8gtvG0DNU28w9DzDcoR8l
YD1YpU8WpXDopoJxr/U7hD5wcpDMaaYCN+YuGuM1i0ygZ6impjUHmNetoXQfaxh/r6S9F44OOxcy
U9qweLYJ8qvmIHPWOUG7nkEtOXev+rk+I8vPJ9tWj93ZgMwNr3fLH0MQL7eb7tYJhTOHfPliJ500
+yMa/WFYU8UaQgTZ1tEBIV8VmUGFk3qAxa+N8Y1x8VNhnCya7mKcTZP+G1rtjnHVAymregSJ/qrK
BaxNjUUyBUIXfnn/IfpFMye1fnljteTVxgP5DuAHU6xnaWbskja5syEOXuom97skbCfulZcFjXos
OUyJYlslC77FNelSGjKBHFa8pkywYfxJPB7LLLA95AJeu5wDBu1ZhvLxuE8yegByC6SJaMocx7J3
kiNA//fGHcp0KyGfE9IlT0S9xx9n6Ei1fI931A++e7B/YIuzFb08IJ4wH270mDrzdl8qRs3AVtaH
lv0YSKkhA4hsu/H0U5/fZ/3h/Pj1ukJbAYAcTWYTV1kXPUPo/2gkfXWDAcL23AlZylzJpOMDz+4f
7KrFeOXlDlR8VXmhWLi6cSVG6uwEawZKRYbDzs8OkS/8KjMb2DNEl2oShO7edazkuigyLdMJQ0ox
3EjN5f3AEYJRpQh2K5RSGpBx+7tgMOU0yXrD6CDMZEzLNFKlULyTIFbXJfRdFyIR5umQsUTd4RP6
/danDJsidPODHgin07/l45NcenncO8POnHFWp+umab3yuxAq/OvqmiP3WPgvd/pwJ7RWvv34lcoc
H54T1MGHR8Z6DyTckWRaog1GtMUCpiDVjeJOXznt5Bi2W1bY6skP/4gqMu0jG0gFlWIoCbdghwkU
UQAwnKqj7jALynLRLuuU6EKFCg7HzLIwV/k0GwWMq0BWJpuVUhGGwglfHx/PU5F9ouglKMGydDeI
t3ZWdzyq0igur0PP0mUmWv1zmuCrfSS39wkAK/Egf7AEUT3BDlXswOygHv35koXtnVEmd9wVFNDe
0JhZGJ/uHqQ1Q01/bi95R9oR+iWNeraEnPxRE7u/ooEOE6JKtkCkunjtAxV9BKMonnpcGUYqdAfJ
91CRCMDvzBS+hPJs9EzjZ0w2b/xsVvqq565RfDtpFy+zykn9SLDYBK3axEYw8THiRlxW/ogXI9oa
Trsaq/QpGhcZlo8ki9nyvdwdpRJpxqu910DzqMsnhfv7ALhLujR5CDOXgM9nKeAKG2+0oh5ScOXI
J8tcD2jMT5//Mcvr5pjk8weTxTany/14bM8HLYFbUu4oA++FRS3w2Pmpz0g/isAFRlz8w2L44aNV
7hMiassK95xMI7wKN5fldBQX4L4RdhnLm1EvOBHDiAGTPeUR35U18kCXPprgIkpC/kEfwRwnHEqj
KLIjs1v2UzIopFwewIFDP+j2Eaf8PyUYzhV7f1V/Gg+2SxyjI+PjFG7YJa1m34eDRtPqbBL4cHBW
iMXcxWD83FljePdKzOg26cv3yvTnVchrSWI07+iW5xgaEKuvIlYpSUybKPhlmqCaSKQyC4Nc1fRv
epeKIvSdh0+oRUdbUrZlanPPt6hL9C/AAGbFU9Y/SrmzPKa69OOfcheKH9ZBDTUMxl2KvRs7E21e
IO95E0ic/sGAyH1eWDLy8hnYrreBMk/Jgb+kDJ/QH4BGvmRA0yBnZ3irTKlWk0li6ZI9uyXGoKYm
5nqi3fneZGC4Nqp7FXr8shPSbk5K6NvpABr2qGkmVHugtyYKBOotybbmh10ET83P75mhNvDIXYCs
jm/oHmHh0H/mxvbS+TNsXoxWNsuNBcV11SLFweLFAbuGZf52VSlUwAXwPo7DYkS4XIs6WRba7IML
kaEpGpJQNDORAlNUyrIg7WM38yTn9NsdR7gTpQ5khKef4tYzkgeSekxwCv2uVsWtld5DTsc0L+W6
o+UtEucatbGNffpa4y8rSON0/j5h+tBzIxso5KFJUPy+z4HWVCVGNNcPbGfiXmmqccqd6iKRan13
TxkSnx9GEggprLn9AwM1UX6cT/tErCHuMIK/JmHcR75jBSqInCAJrLI5442mRMUdtWwgrichqNv2
pTLgIksO2m6Ua0P+3h9LaeLUzbEWUMG3C952JKZ2HWxaga8tIReIqtH3oPmAox7d8ujzMUWZFyry
0Ywuj+oc2LqqPfdA1QwdzP++/bOj66sAh8ByW6VStL4q8+RtHHEzac2DWqTi7NBswKcNHRg7TImC
n5VsE1LbUOIEkyVzO3Z6FHTAMmUAvCuemtdrrpMKAOGBEtJ21wWs4s4EoOfWET0qvavwi5SlvNJs
QiWoKefaNGRBIh4pChgURqlAaqlbN0jgW+P08QhAnWWrpqC2S18DOQ7K7gTzSRDyjbuRtxX1/dPj
3DBtn/+RMa+Erz/gAvNeoBGAgQfCR26PJ7Ew+9GmwrxVIL/B498yXIW3vhsdmxW9SvgioJGm7sfu
OEzmZ90AtBr90N5LaC5tUK4q5i8isk/AgkIeQrxL5gxOjmtq7k5wVIu8/sB5TRLWOOfkLDQjJNaP
C3D3zj/MWNpFGV9bvkDZdir5YJ/qYH92LTqYGYXO0DvzqERsSDiQlh7upkHGwk2gg66+pyoV/5mp
wGC/htvs4M6EnIL5QtVvQ8nyeqZxLrxAasNAhxULETVOFjD5bl+0iw6YORjVisf/NbtS16ym1t+A
fABc6bXDvKM8DLSoULTsPCdvDuKvPqI4Xmu4y3wx15mx9CwUWSoLLcexC9Jpoi1921tmdFu/NCH3
GEScEKEmXM4y9oIevyLXyyeafHbw52+eOoL38/bbzoBvssmvcvfQZgqGispH60C7mMxr/sY8RWXe
kqQOmkE1BUkJBGHMDHEx1FrY3wL2UZTV0c4ApESmzFBLUP7sVgiI7B67MJHEJdkjZiv3e1Cf+E+t
TvudqJNePxFRQJ4inn96Br9BvE/xwo+083CVSzjzTwfpN0LupyJ+8j67m1SIgy0D7kNYz8dH+ufT
JsklSfXgcdf3PoAIcgy3d5jMjTEpkL14szkQgBOc0yFcI1pdyjCjLglo5apUUUZBzH/fUq9rTxy9
Ab/lA6l/XtoOVSGuNR4pEZEtfiBVgypUXdRhM5KqBHVKdhM/zqMQ1EkTOTJILgm+cmOYyaaEQN4N
vcVsa/HOmn6pvPE1dCH8ADat1SVbQFpp3uRmW72HvsBgo+6et0nuM1RSWPs/M2G5f+1QhyGpM0XM
g7rmapNhPDS1l8vLf6xfPjIh8GM9fFVrL13kOD0FlrxDWE/vxqFTae9b8gwcxGEF0FO0/a15hFSe
pwIZmfY1l0bJ0vpcyXMBFYt7pvknDIEy7NwCbNXisKwtyexYJUJ0O7S7ju/OzME+xfZQxCn+6Ku+
XsY/2bLD4gRVnukjqedv62tJuaYmytr1PM81Uk5NKnJ8RIDFs80my06GEnsCDlMORsM2WxNocnqw
EmWGsYypPgP2KQyCoEx6ylelb/Fvm6LEPvK6CKZczWvmmhdSaapUUrd6X7bo4a+oNGSRWEMzcoo/
2GQd/E+YrHu7CA5X1F0vymudMU26DW176afAEBjwvKoAIZPJ1BdArpuKcIT5BeiVdVdstOIgwzxH
wywOoKyu4K4+ZYYCi8W/RQ37zHj+aQSOFBYRXwfF/AyZ5CsfAOJIUBSwGHMZKh1A2KsLmBYFgSn0
70IBuXhIgfjdp68+pUYzlsA1H5uX6AU2LAJWGSVwf8zh0/PXtCueNBtlBQlgaN3Gn8F4H4tLL2Vy
8qhiNDc9NEoixPW6J0gY8wbF9WXYxwaSvvk/Dh2LlFGrIrYkma+5hiRfI3lRlIHnK2FiODygsvPM
xWGUEnyGXV9fpea1/OzVuJhezaD45CxaLtOEWmCv85zzSrubhjPgs4R1NtWvNdHKNa1ITOgAKzPg
jj5ij/DlqGrlqdg2j5EK8YgysMtkAcJl54ksJM0bMqVTPftW9Gus1rhCz9Yyui8YsUG2kOglOf/W
JQMzwxZAIm1naenKh9ti9bFB1GXSifu6z4Fpl4BAHUDiajcgMs832iDtVqXpMiI4FQQaJ2Z/u8nq
Zw9nBiNXUpt2JR+e24V3njtrvTgRbcR8vDndbPEthvZTaentbY106NWo4rYO/TB1nOz8C6UFpnDu
X6WpgdqmxhiKVRAd086EcB7x5i2830D2PkUMcHUJSF2Uu1bZJiW7kG4VYF+rPfMb5smlXvjbHGpF
5yDtRlFtwvYg+FSJZl1qCgZwlcGMaL2Ost2AXmi4Ntdo95vSpjd205xG9qrL/WkWJXo0nGzZxg6M
c3bg5NbJbBCBzhmnHd9WPJ+3hj4cqk4l7R95I5tg6+f86jEIcXsrm7TucFjn7H7JWMNZqtgSpCjm
8JAz47TdafIcWk91jD+QXrkCXKBv8D3YiP2YsvPH0miHmldGLhbUrMSJu4yYZ1IVHmTCAm+ZA69u
25PF/ZB0rN4CGhfrhPwDHPQSAnqQM9Yqn1ylM4+fZWcUEHKhkDsmDNkpdvvw/0EznhHctuOrBsrH
L95OD2A228xxErmGVRdfyatNCvqRgSSfvba9SAxMgUu9Zoe4vEPAYNq8yAPJbDQaOiXP0UU1TM47
EUUudXU4756BkJeyHsRhhiyaFf7SfIkDduqv2NMYLcVIrYzAYyW4l8DpH86Oi5GKplB9PezjIYpS
r1HNKRzPr+W0qm86VNIfXQ0CPhAlMwW7q3iCxeBmDsZdZ6KIhz+oHttSqRH6JYxuKbTtS71IWsp4
7943XUkXRpo3BRlTgfcbAODXfu/TBM7eiu2Duxb5PLB6pRgIcALCVZjlEDkMrhF5//xURnQlp6G7
/0h4zw+fh0uYIEXNIb8vsoFHFVr0RXqTuyHW51YmFRPoTTK+FnCzWA02/jt6HdF5jLtTbXi9YFXI
j5laTmvEPbvjk18F4NymDoD+BU3ZrL5X4oSvf+4zicBov7w1vSL1Xj2EA3m1GdNW0nBldeSm3a7J
r3d/cM6UX5xZv2GfzEsEzhg2fa+Q7hUZxirBCynFJ0F4PCcY7918tCBVwyqKmsl5xWZr7HHpeaaO
wjS3g8Z6SzCsVh2zZ7t7g5rjnyXvvJZdA4Rb3wvBAJ3xSHuwrPwj2tCrSkhNHjDbleeRwlKvJ0o5
pHVGrM71LH8cnIQlQfiSDGcTstSDg2akve3vqzf7ECN9SEeRnNp/tb6cb3tc+j3oll2JkSBLMDZR
kzCiyOOak9RozVeRfxsuiv/taTUQV2sGcWaAAwIHxOt7yDxxPIe7qX8aYaMX/fQ7+WlNG/rV+pcJ
7zapaW63dr3TxAQ8oJES5dIg/MfPv0IHF5xS4E4SshYJmb4Z3dY0U+3dnI4WFmLWMCJJYVbKDHd2
6Ml8dTD0XAVUEOb3whyIUUmWM1JMNK85Kr0hecJ+PVGeQcwUOjvxPBbyiql05k7U1nPOvnT0Y2Ey
gh8SOSzvOFuifKWAk0uVoxJFhvzNm0Ea/rO5l7USXI7Z9/coJbuQNto9Q1VXLOxkLa5i3narDrwX
u1qFiK8KtTSRQiohZtsCrJsNNiVAIpz0PnpLN3ELGjJVzkBICvc6q5qPwQ1Cki9BUyqLJwpIkTV6
fLadCBCDMGtbulUwk27d+nmFReInL0cYBh6JI3cAPQAOHLegV3MeXKUH87uCxGobssWHt1zt/aDL
yfDO8m/Qhcl++ZDhJGhWWKRHJH/zUxtYY5MI9luTNO2COXxr4FMdNc9j+U+q4/+fS2AHO/EDQsvz
sM5CvR2AI6I5gAwvUuV7n1CwapcFpcp5TziuJpx7pojsmuPM02Rbi7QwHV33I7hDkgxBFizruCLZ
8QY1E1MDH0eqlD3MoGnoWlPAjjlE2dlXvqVsWx6tEe2jOWKHmUiO6uA41R8glpDOVH6Z2FAFxZC+
KrIMoRzzFZX0bj1+uSPsscuQl1pfx2HIWSfy6KqMpr4zo6qH3ncx9okIFzSd0GlJrQUal+g8RvLs
L1KNctdAVXflb6bhPBDSo56Mrx4p6NMVQ1VTeAmY0OQE4oolZ8Y6CG+9kxob3teRPltn/eWvF3ka
GqzVosjacsRLySIQDh/Fir+y6DFQWsGnJ1ev34vsGsIh5eTLVAOQc7QkRseYCTLDjW3D+8eJLMaY
f2ecABDhWcIPX7gdzyKMQDgv6DRqFpeoAxxAaH04p5p3AiOpwfGgfBDRdazvR210X6iOYRZ3wEYP
4UFbnRf43wtZAGg0CnVfLIbnLasRZoU4ctlGEc+twDnwdSpT0nlpro83vZGhDOI2c//NYq1wUYpz
k68ga5zXFAFSpbvSNJyuGQbN8G+Ehdg/RF/1Nl5e6RX97k2gTF/z3ZQPOfUYa/9D+92gZQ5wNu98
3KXHOSHdsi9juAj/lN6+L29ThYiuVjeusuHX6LeWIcBlvpjhz9JvokLRpfL3yCoxpFkIzeVe/KGJ
RkNUSj/YHT6b/8w8u0x2NYZDrTSbRyVI58b/C+tg/xqF+pV682hMFL98D4+g131b8ID/OIgsDHNx
icSfkQh6kZjZiKQpu4leohR4doChYNpt+PjXDt+8Qf47+xI+deq01fcNYRLh2humWs8O4wK9eRCV
QRkxuxslrbsAsGebncCntytT4V752BzkjzmxotTOdyarCxK2NPfFpzI4S0ank16536TO0OSfBjDD
bJgjARKuuegY/TiqwXTCnppNUitvmx4pUIOBwSgC+XZxRk3cFMJkTVTSfFTMPrqWlXmbDuWvN4K/
1rbgdb6oPCF4tdQE+srEb2jXljoHl4IP48f5gidEbRDLDo77OC0PmhSRisC2Y9yn6GmaSVSED0iG
iuqpVP2cU44uwPFvrDBthMc8fWdOyoAXtg7HjmYVdG0+JRGbOc5Hj2Jrf1PYSE3QFUWDPB06Gy1p
TbzvsA2M3Wef5TPTr7bRuUtPwLx+KXZb/MVKj0mz0qzKv7UKlD1sX2lrtCY0cvxwjmLoRWm5L2qS
Tex/ODt+hQXYHxjoe1BkUuoCufVDKcFucSz5WEya2zIqtbFlD8gPguwvyEmk3Q9ECDh65iFFPtgW
LHnS9/i0Bkxi7/JCaCO5bMb/Be8qIhRSKXvOfeZAGrpzmr6QD4w0z+HJXZuU9BRPnqwFdrfDbk7g
O7VUyvNK0A4HitQqmcajGy/++/eZgNtMrtT4YI2eyQc5R+lz4lrVrBqR2ZKuG133DF9qC6OiShSO
QJUCT9v6mo6/ob+C4TtSkPYhQHY4X/6vIH7FAi9fQSR6OJ1tlm9uffvVtv0tTfuppX8YwJA+DkjR
62FeROyAGTXQfQP2PoUGrkeo1bAHlOQlFijRQ7Sxj/Z9CFD5itbJqOKKStun5ir156RjANVWweg0
ml7bQXEDP9t48Fzs/CraXoirnUNysj2NIoKvAGahjdtjQZXCdlTDQfSKhzP5oP5xSow1PAWu0B0u
MkXDzOw+AmjV7Mnqx99V1Xuo0g/LTbbi03uOWpdeA2qERxV8h418nWp+6y2uxYJlg4uE/2RZdK24
x1ohRYK87MMRabzPjEwpBxqNwSzezne6/8b7yUjVCrUE4f4qQq5zHHCsZmySumVPwM9OQKV9TuXn
WsU0tib3i0XJQJB0XoXHOi16hZ4CdFg9CsTv0otJkYmNblKBEJCRi5C0R4l5ZMXBK1ttYcBGHbed
xHPf0lIWAQFTf2gCNIzXgsVOzPOw10cp4fb0iTVWlS5BZXQhUDq8DKSjVf643lxkUQItpFCFtsqg
8CTziLLbznreU7kD9Sb5RjrgypItiVeGXG41Qeo69Yv6/5MqU32SjJM3RrFiGFnqA2L1Q3UfXrkz
bYlMFLGurwzA+POBsD85sLl/T2dDEeJo032ojpGVFOfkrqEtwA9egEItMyNnrTvBlMvXlnR6LlJz
0YESp1iG+1q8tGxc4uItsnNgs8139EYG5qfMzrPzmZgzdT8gFKEkZpextoBwYnwJJJZ0VoCtKAuA
oaUKAD/t6DV9RDjEP6iWmkiTBarp00yh9nOY6JDxEM4yd3xG7MJktGXMefRcRdRnbT+oiDyjHE4o
ppuwXxXHo0rx/f9CzIUbVmzJwA1jpRmBhinRxxUOJcaakjy/AlYKe6YGL8ECqIG4iEOcEuzV/7JM
UjZr6DDT4K2eS75/Wnj14e93EuhL7bcF5GTvC3KRd2FCBVxNHBhY0LfnN3RB/SetRvCocFOY0m2+
17zIsT8QJ1LT89P6Zb9cLl0KZxZQLV7OLfYKoeyMwxyTuvgBauSEdsRAaxucH0EyEyviVN4BkCQq
CNaXk08L/WpksnUrvpZIGQQ4mklEA18G6wz2wDOCstoI/SGyKNn38xC/t5hxd+v2JtNML61BL31h
/ansuaddb3MAzrN37leVZ0zO/uPnYw5oXKrNmYYwKR67SoyORvCegnuUghaJyjleUEzWEFX/gqNz
2bLYOzDIZn+3a8P6zs29TLIIJCppEavpXGJW9P8ZL+tIK3qpTHgMk+J7uiPrqTTQ3f5NsgBJ6P6b
cT6959VwAhtsfyMhTLEJWjXGUlGi+hqtmI2Brap4BO4uwtYX4HgxNzBM4naukFu3z8QI9YdaFP5M
aEiNL2/lPz7+vse/G8RBKrZPQzHE3+3D2AgLKuZ5o2NCV2zaBwu87IkjfkuIiMdDN+nnLTgzVEM8
TWIbVgE65qb/4G7X8MqjO0LqbeIDzpXe6Q00me216wvmhuaylhhJhBv5pnkdjj7sYMEDb3V0iSa0
Ax3rUghG12Yfx2WY01I4A7ea0gZf3El4n2ua9BtHHW7GpjzJCexg9uL1whanWQnGzL5pko0VytMG
mkAZlFmeOx4DhZMGE8QojpXelZ9AIvQ7gjYRgZ6HXyspV/SAtZmEypVyBxBUNHISGl/DwirxslEP
6gXG26fIA7NO4H67rLoJaxPiL54km7/1xCCSBpCeTHvWUwyCJUcIs5/ETPh6TexR1LWg0xt7mwMW
mS1MEr9B39qLXq2diqgZUmB6di0OYQcxty6Y1gtcrRwIaoBrICo0SGYhfhGlOLtycdBzBEeAOAz3
h5WMjkDg4JmG1xw5GIS7z+ANDkYX6F3+ABtX8Wwt31H7gK28hbcIWmPTvr+cI5uw2F9MkOQ4q7RB
bO8U1TIvUt/QcCW0RWZdWRAmVTtWVfiUBgdZxTckFDQjQs5JklCrASnatT8veZKDGzhCSIE7gcty
zcZWgNHwfohxvHVF+MQ1UCtNoGJFcVK8EC8mGVH5AXtTzXEtHjFpVblEs29ItaPCbddNaxUm8X0B
lGPIiCW0uLN6heUls5ClfUGJho4uiRe7NKGFuouecgEeV4iIv95WXbob5/2Q04aJoOo/1001UD7h
lq20irRS+qHtuuRfVq5vVFUYvOrhKHTYx6052JOQPFngXS8WoMRUgzOte34d3lGfhPavergPI1xq
8RGV9+EYtbz1fMGkIGlfAraynO19HnmiSuRz0W14OhYDIpEiAcHxk5KCHLa8cxphmQkd5visWf80
K3OeV584MleGGlegiy0modEEM+dummJhJVSXdg2XaUvJZ+/7d+g0l5wUWmEN94PYvE4PB+cP8MLj
S3RugUjRxEnIDsaH5h8X4eTSd1pWKIohTmvFsJUKtl4R68YfjRg1Qz+jgQEHthh/Bef1PhUWgW3T
Rrbneune6rxA1J0GGMrJdtvliLkx5H0KBu4LhbolCWCX8u/PN/HqjG2oowUqOhE2Fb4EDLDMs3Ea
6Mh28u8tAUF8PEKnny2uNKD45Op+JJybZnE0/M5gAMhybtVK4XynF1galOtk5sQXWyqCzR38XvTy
gJJ1j8ADFRkh63M8JRU6FSo+dxfN4ap1GZOJlOuXCwKvcZxczs5IHXPE5XEoTTPrEOAtD4dKU+dN
uppbbBPeiGsuCFJzytleXA0ZqlqtmlIiKDswGaiYuQTW/n+IV1FK6bVP/L04FON1O+qI3yGKp14Q
nvP7UcOgpg8XbNXVET1LvBUIxtVS7JZJM8sjTaC3zxcUb7zjRPG+sTQkdY9s6Jmv8/ONz+Uqn86i
6N0Ecs+dIHLtF26fL7cAdBUXtDhI/D++uOgMyEiNUctEIeEES+xHB0YK/LPXW1QrqxJKuIlgfl9t
fb1K/tSVDowcMuJz0z5Ie/xCoViFZYkK+vas/8dvh3qoob/pbh4iC1H+AaX0YxrcmJ38PiMVqB7d
m3j8s6F0cWHEsygMLCD0/I6/wf+6u8W+nQrGvHU+89fO9HwcMFG64J3WpBtO6xOwhLmI6gzqI09T
Zj+pGP2WxwSKI/R/qwhpyaPtpc6TRdfGR7szCH5qv+t+lidWJwup+Zbe/mGrDzpd1kc9D/OoSNxE
2nMC7/zwvfUgTZBhakzhB5LRT0zHAkhtcMclsQcBVrF7Ia8WQHkk+tx0nqyCUm6LEaNs5I5i09Bl
u9nTQ2zUursjKwwfbioTTS1rLa4CwiUEDWWfjn4Wx+FD0UGvBNv7kA1AdgeF0xEPW6LjpGmoZyym
4y+eFALyA1F6LFJ1/L4zlckrY/1LJ770ckTUYLeA8kh4hR+UVQ6tFZ7b3PIAO3erXVcP1DXaRI0u
HS2kdSVMtyzHiaDcTXTHJ4gPdjJ786MVeBwoPNamxGzF7Bvvkqh2pR1zc35AveNUoJjsRJ6dTASX
WxwSEds+DA7RPDr098UTHVECY1JWBArqatXlDNqazx2qBD314YRcH7pb0OX2vcnirMno3BKmQ1zo
CF+A0cKQEGjxJt4INuTtNTgdwjTYnIxc0G+gN5vuIYUniOzBcvB1SKl71zn/R32SYOGnQzpubfx+
FYjUhWqKOB7GRx17qUymyrfqYC8T0dkT2Z/dKYyWpmMyRwsxfxA4RhSUC5JJOubxphrCcnHiHuHq
dUCECVAXRfNnSBIdO8c/2vU+/NTx23voESvrMI0U2fyT32S0TYn0ryKn69ClwjUfj1SQtLem4gbA
uD0wD3QDz0JQfy/V4AmdtrODQsnv7d7UPa7UpOFNzjtUxGvkiLM9TOl1OYDjMPsnTIYdCCTw37th
v7lGmVBGprmsXGMNlXdhQmlLsPqPXiDnRUhoa1rFsoiBwt3VWa155FP85PZE8OPOvleGxcscWAc7
iaSU9RmJwEjUzTEI81s+i2FgbEgkeOAPDix0XH5GsJ/mYpYf0nEDX30PHEBIdK0qrOJevR0z0p/U
s+HiX9YiPZeSrC1XY1PAPxa0K0uRPcvwYb7TaT233Yms31y9qeGUS+i3G0XaJ+FAPJjXBD1+bsLl
jKG7CI1UfqiK3KKkhJEyoAZfg95f+5e7sVEJCvSwbxR3BSPiRaCbRqXM05FLT3X6S9L7jZCZXo43
dA0oR5LNfthXScGm3sMKXv2TVHEn0MjoXCPLfvEh4jvTD9t18jG7CfmeudySE/XvV4ZoRMJEOdTh
2GOdCi4naTIm6OjHUWwJ7WPdmL2kP1/6Ar92YTZwUzosSn6Lm6JZC2FgT0Pog2wQWDQXi8c7FOGI
Xyi/kzyQYQQ5ueEhn7bUB+bKT/GqU3DqVvgktF9zewryJah+QcrQsDVr5cKA8m+3oXCk/9SKMf6F
n8QSj/WcfvGjVfyx2Zxk8/kMHBfI/K/cqpV8kl2s77dUE5fi42FugyGj0+CEMk8T6DeKKRJkzkaz
kx8TzREVkx97ftOml94uTIu+cxnFewQhumP7AcLp6Fh9HvbhKHlAr26wdOnEdxCicMOOfvzAghAb
QMUkmVJ67J3LuwRA1eCo6fFosF0SwpbCUmSoF3VhdEmjAiR0eeWS7v3vGmu6HdPc3B6xEbY2NKcH
u+16oSn6HNe1IJBaBM1h/Wkh+AhwBPL21G/MjslKqZLmtvrjqjxy5r7I10GRocr9ODRDV11M5QO/
BfwpqOXtndScM3vm3SmQZEObJ7kMqkynyA8EZYmeayijER7xOzb9elQETtX/xY9MQ3H3mRIF4ZTL
u3NoZRqzIntGRLzy82l6tRB3hi9qJ0B0bjkwwd/hiHPRGjQSgi8yHYlPMUNsjUNIBrPaZhR0UIL/
zStBA2tbr8M0bXvAYtUOiQ19qjP9zMBZ5gRhnUgqkd5XtEp+VvDSa31RPEXE7bc4O7nv5vh3Z/3Y
BkHLksiD64GxJvpJP/xTOoQxQWIkbH3k1LsTq3XvS2yEmiJLzbEm8nTHcCtw0xYR1V43zWHh4cCR
2hvL0bgmhZuREQuQUC2u6rw6GXzWnnC4yb1LWEOqWSPFDgkHV0BcLlkJMKe50uMJvrAFHh7uAHoN
h/u5snbmtrYCehxiCtimC32D8O2lFrTNIxOK37ug1FMx48rWxhCS8adpve8DRJtpwNX07KQmicJP
4nwkwE97IOOKuQu0jSNpMPo+Mtian9/q/fuVPdpZNmAxKveKDA3pdMxEq18fP+3icAFPeK1pVKnW
C8KL5mWFuwYOptU32ZKWnzvdjNF1L2Ut5ISFmBgNSaOALMGTo/Hs4Tt3DX9y7bpnVlDpDxaRHbV7
M3jIdJ/fwTMgml+kwH+3QRRWu/euJ7RbloQFRu9DsClwJg8Bv1KXW9498nsOlGGdvd86p7kg6wqY
ZZTDjY1gXKOSuO1bFKJKx6H9Fx4pf5vQU+HBWBmL3zPiZsxgmcAYshl5c/V78PbUiCuB7ZN9t+0P
d9bT9lpMhRYfwtdQ2D7mggg9pzRt4PF0rudY7RDMQ7huMDuC2SxzuOXQOLoUVMb7ec6MDoqn0yyS
HQat7L02S3FyZ4cyoo4i7Bi0z/+arKus20mtPtVyF660UwxPvm80b8Cg6EIuD0cIqUO8MJMMMHJZ
iXnQvf1uGNP4lsoz2vgeriZChceIf18Ez5mbajUrqq1vNZ049Hyg7igMEeWuTNnziLiumVhkrcek
oC2tV2zeay7iiyIxEhLXWC9AUr8yxVuGNCc7dphSxQE90GMF1HkM54/iNqSniN7AZA+6giwFjicP
r9Z2AVHYLtxVnfDms8504VFMhfkXa8mF16Sm+rYiyA3SMGxwRYuO41aMHDJH4ZQo68n/C+yWdT1S
NNWPorW6V5oLOFVPRZhlvu9HaxZwy4ObW9OWx5kWqxM3qtLRHo670FA4EpDpw3AJhMDwxLBaGlIU
bY3m5oia2j1h96ucYT56h57qaY30Ap+W5mJzdeJyj0ClXWnaQdEWoPi+bkzuvr3mMUpKoBkxTEaA
ZqiClgMvnjWZWTkUY6TfEi0gYhxf1X7Iwwotk/lFW4boB0NX1YGhZ3qyi27CnNGJPPEBjudU/JNu
Hus0JHk/jzv9GmHJf8QwyTWa5wDnPl+/O7hs+xO1igu1IIkLVx3SdOX98boxQMKGh5NEQZEO69+H
a4F/4h+UwEHQMwP8iOKOSl2GOTP8tKL+ZSDDsg+CEB5pQIt7rvgYpfV3O9ExG4Awf1nYwZPD4uFl
wF40KTNwlOFhHn/YLXNxN32xUoG5ecoPQlQ1vzjLRJ4s4FohVXm/Wq+isLxZGNyo02gGPcqSu/ej
Bz/9jF4txS9t4E5JC87W8qtwqOjn+1nXAVD+578ywUQphYu/vZLfE4GlB5sH8HWnivEFG4GhbyPv
0hm/DbiBrYpTmN6UQtmdae3RvgTkUs2xyNRj1z1X3V4XyZGShffh/eE4O3bQBcGAMholcaqtao8w
c9BJtWwpbP2jaaRgQjkisL4J/ANVfAKztiIo/HuLUAVnkHpGRutlizkTnJ/1UTtE3gYe0YzAFGZ8
QusEBxWrueNYtQpCRGgpfFpHtVFD8cDrmWhdggoNm39vUXcwiq00ic7Su/jho9TrGt4AfwnZ/YWQ
YiX5qGferOIxNr18WesgWw2HIqoSGjeJt3NeAljw1a7ih6qZaNnKfIxQjJPLS9rZxvkSd/3o3XCy
nIIaqvuXPR9Lp533bQFrXeEUUunmGm1bI6Th4oWrlD09/z1UpHDUpVATfimiJvgnvXfFX2u1wbTi
ZpMWT7ESsqBhWigOiRyOpTiCal8QJqbmE5pv+UzrSjXhnK3Jz7WIyX6QcuHWXQhfJvKF+yscpfes
5FyEYwI6zzuK9VH+ckFGk71D9xxWjdDYaPx/wcOMDKskR27dIiZTGYItWHGw+P4W5tHqia47IOQ5
GtFkBc5K2CvBS9By8Gh/3VubZkfL7MMzrCz2u/XhWUlysTZb9UL2kE9NKN+PC8NqQz3znb34tC1S
E+RbtkZTONS+844BEgQVuaUHJ+HmLwX7lqHZtVVqNpXMyADPnZk3djVnj+oPn14DFC0MYpcU3XaW
7LwvNaBeoZsXvQXjiOVbkMxOJEuGaJxu9hLJYLEo07ZAAHqO4pHZbZWImZA3ywkGV42Nu5g7eW6c
FA3KtEJNMq63DtEIrxBxA/i+itcny4HE1Rq8YgM2oPtAEY97FtnsdBTJguObctjRwgXHrL5xgS2p
UhYxmv01943musGsi/X9EA8zVKK7joL7pOgUjXVaoi7cq6h08wCAQnD9Wfk+NI7EHj1UdRRq0Ruy
8NyWu2xuKYc+kM5Adzs7xJMhRX53tdFWmA5AsQN572igyF39Ja04uEefk/D0NsRElyv5mIaU9r31
LcIVT1HMQJ4PFCQriAIdI9UVmgX8n2zni+2SAlsnIxaWU7njkPciNHIxJjNzfv76v5JyhWu8iEps
z1P5PF8I9S495T2oSDPpOsGXTVx1rvPhtZk95T9buw7wT9UsZaDuMw9NXufA1OAZslqFJS4Wy7si
Xl+0mG+LL86+0nXNQKi+rhYPUM0NNa2b0jXVHM4EN/L6PLv9SVsDf5g46iruuCW756bKNoppH7/H
qdeZhaLwHGY5JAXfmeOyc0VW8y8Thcgus56ZTgB6CMHppZ+2OCtiFtNGir/kUIEM+M5FHrzY9VNM
JlgMXCGqozp73DLBH59NJcep34nPP7QyPVt5+faD9xRjUkIpSDYOanAw0RablZi45QYCKjntTiUZ
nVpFrqPAJ7du7CiCCTPjwvaAOaL9jtL2vVtnJxPM+S83Amtz8CRUcSjP9koDTfv0d7OD34heGCQG
uEek+H9xYMdqo16aD+w9SbuU9OC1PeaARnflsgSgChIGWmpHxAajmYmySdQt/vo8HHAfdPmKiDI+
+Bml0WIbFtBHM6y3jnrnm6jd2SFg3WTe4r+mZaFC5Myq6cGRzwpqKt/0zzQshGtiS7GOAmZJ3vH4
8nwK6hY1JccUEvbxGV+1ZhUzYTjz+rBGgYpDxtTryJrplbChClpTGb4bqIXc148yhVfZAj9qXojz
k/LTkvZEZtMJBrkGz/M99EEQKJoeXDscagySe74ch6Tl2hb1nhUSKqusaxvB373mmHn+bbChxuzD
LSopdJAWHxsF3jihdIWCi/MiDf25JUGzwPmqhQuMiy3aO71EKwol7lcNeB7TK6zg4YyffkL2sRM+
alSZq5ctuwkIEPgPaOnBmlcdPOHTp3xjTZcrRSAuc0YQo+52fy42vhSEE+xJcFGVG8RxdPdmhThu
YX+2oLwI/PWQDeCDR0scTXUYb1ZW36pmGns/SZuRog7VI9EUMVhMiBzj+T8YVG/fXQlZy46l0gor
0w5zk+puPUjrHvirN4/C4HjEnLPzMt/e4Ep8+24fPn+p0w/Ddi2xIrztRzcOGS9z/v+2fkyF4oL/
GKCdK33HX7UObrjlHMuvFC265lxMyitoBierM/fjH90EcnsbxtnqsAPAZIxHIsuwamucm+lfP1hE
MaQL6+wjJWUsCLfkSC9vo7eWWq9195rzB5VO3x81+csGIyKYjGcZS6APZsugl/lNYyWJ6hmzlJZ1
SteL4VV3+l0v7p0EzN5B0Mn5RkQXxzLkkntSjFqoetlHk0L94fvUATkhS3sI0A0adHu+oXz2DLkX
RXq+X8ZZP3wgpL+VOBcb5jO1HD+I1LvRq8TvvJwFDXRlgaVrNt6fF0nDFESMEdKybrnBeQQ7K6iV
582A4Xn5ai/QU83EvVLNAGgmwb9WAFjvHKJLFeMbww8Ed+ck+f8ZH/B+T+TWAJniDlR4SCCIZ/xh
xNGWccAmh/phoAP3FzaA2B6D//OD2ihg5nf0eNksGnQ9c6dIU9MXeqpRD3m6BbtEH7mpamsbCGbp
Jo7ia9/ZdQY59Ukoc1pPAKEfk0tFDNR2FlL0e4uOIQDC/+4qNXSAu6lfJ3BrctGpgdrC9mzoaWm3
ASyu08RRB4fYT8EI5GelddjUniGXETZm5u2KbAe398EagRU4yH7nLnyRf3GyMqkBbr3vw7QnaOVN
+9XTnbo8EoQxK0G0i9f2/8JKUps3NQx76sOOF36Vb6DpEAWzATiOfRlsfn7dhrmc3abF4wowXQFa
7C0mlPNWSQnF3csAau72tl4eAM9HlxkJ4TXda0vquVjVY7Z7AI1/6lmk7HSQthwtMdu8nfpx9vj8
CoM1FjFbsN2J2uCQkZa/Z3v/XNz53SSxEc1hS/LWcXARdBcO6badaoIwdW205M9IVRzwMvFfBRER
XFEqaQuJqsbOTo7YG9ford152aUxIFnydsQJGPCUs/rtYkySwlgPa4YpmMimudcR9dbrkCilbLHv
0YRnX/8NDfYBa0tVlJLljO2qoXsu2/UrdZZRWjSqOH7o0OoTvjz9SRV9uTpwV4d29AECIIjz8wDV
8rN3Ms+ej4gdI+QUS6UqTeMmW7qwJYJS/oHoC3wMrPGpkxJOdtQvVoSdhdDyFskRYA8VpFfWW+NV
L44h66EZGRcMAd+5b7S5Z2tYZ1zqMB6Hmv6cnu5xRUl64jHYgbrSbEaJPgF5HxrMStIsHJkY4m7l
jWlakDkUJ2NiP0h9KbM3U2JqzmYGrBylEL3WMNFnY1KDTKafqNifwJa5CrFWUBfszARObdkStKR/
gedvhueZVlKtLpgqrI30bnSwCDcwNG2vT0wMmnLOYgga87RqqLGGwFBDoC5GhE6kV7Lz7P63TqnH
nWFKnkelTpWJxinoIt6ocMits5zfGWkpmpZYIsh9luSIXU6Z0DbFM2m6uSDRH6MnBU/Yj21l/5pi
7lX7DoAv7PTpep4FN6BVzWXqtvWQb+rCJH98OS6ZDcvaI/ifvkTFGYD6Piv9dW1wZhmqxNT3KnSc
vfbvEnnR0006uXHNaKsjwskrVtBKgKbZOEj8jKx+qUFet0srVWxPIE6dpx0twe537q7OFOiucuAS
SEycalq9DYWQBICxG8qF+vqfklOjWBvk0SyN118SpbtteGa/NoRzOfm1oo4WVNYJR9eA3jpOy79R
gwvyy39lBwG97K9CcRnsSm2j9HCE/rB4+nsX9BQfx3HE0t6lJ44yy07F/OcXmR6UdigYf8RIpuvd
q79g8Rpkt5N/bvhmyIDNUYP5VjGM0I7hWUSUSce9Bwj+Tjsmd3KfWb2Paw2hK2QZLQvhpRmUjdFk
dt4Ve89JrPaHSRbZw3ZrlhaBmRa0G/wD34qv/jshZGZeqWdjAWfPU5TNtiAFcqeAkPWtuCaxoT7d
hgmhQDtQB1DAF2+U7Hn3gqml/rKOqWPElxe39nn0fiNdPnM3H7qDMT9rKx8zFKBTHvLuM/nF6+xS
+VzPKCZkLTpqARe70/oWPM7Kj9XygiwkJgBuPAmUgspkx+EvCnA4oJp5Ap47uAlIlerp9tp1e108
6eMaESGfRFIpQn4P2o/TNxawOGnyQMy03HwXQG0wvY2InPagN1nqz94ja4WT2OuT2akZ+yvTg56c
iYGGW0Mo/1m00m9Qay3jNtmOTfxplGZF0N76aUBOzj0APXl3GISU1rd63lQjJiZ/wFCiK7UUyxsV
YflMcxyxalfU3iBo3AJUHbsQ1l7fLP788PeiY1HzatrtD8ngt2QtWPIMt8EHZ4/sxbXpknNXx9/6
+zJiZ/HaEV3q5+EvFzILBdgoqg0DS+Jiw3ZZPvLbot+a6pG9NfmiWIc2IXV3SlRhLv5DYAo64BAo
kcrfxhxsFs4K69T6zbg0ugjKVJnxvpvlNHipH5UArRAvE0LE6cPcWB48JLyHR/IuPeFFy21pqvwd
IXRjbHX1wxscbSNo18WpG9BdNJ6Yk0zhrOVx6pxw2gG7+lGUazRCYNpSxg81oQY3MECLAXO7gdI4
nfvy3F7eSyGHyEADtZ1SMK0JBTPtJ/fWag1GEqdT5Wdyk+HtaDk/EplnUMLo0hau7T9H3JoJ6Ugr
UDi62e5z5L022Pa0vu2MFTl1ifYNpr7TAa9eUDDSVK3CZ4vzuN0g36t6jeEtouVM2PWjfzW0NOq/
LPYO0xfmuxrGqtOYUc1fCBYFZC1sFIZTjReJYKRVeGLkG5e/oIsfomd0ZYE9luAh06T7Hxig3euC
PHVCZxnk0/UVKiGI6TburqQZhDsod6YTBSCH6+fLQn8H1p+2fRrbO3i410td4TzyZY5kDOVjGkOz
ZgAi6RR2tLFGAFDe0fCbJ8zrAPgfX3/yky8mMKUIi0zRxIpZgueskh8iqVv4/NaNzm6NedOPMMf9
eD/SPCtpxENSC8SqfUxEsGoEoUR5smYe1IySYPLTDbPwIKINxG5SWYmkL2HZFgvxIBYNY9gKoD5D
YKg+u/C0037r6/ic2mkwRyYjTBzEtpWPF/IZrHK97v6i7qTh1b2rpEe134ri/AAEGWGz2piQttAO
/mfUNxTuDnbnt+MgYSo6BPMhbRlgyHAUWm8i0GUn8Q6sNPd7EJlUEeW5+nt31BYtX5or7zA9x5Ew
D3feinGBmfsOAlptChG/wKSIjiOcqGOXVY9LgPwhZOCCx15s6BoZv78syWRQ0N94+AzJsH3Jh+7l
j6cUXN92mUDBDoLMzH3PkSKb88txo8pP99suGxdjxEO0A0w4CBWcy1IqGAIYE4ZuTvdzxlNV8SmN
FpxdDhQiS7ubYoJfL3Ss+SuiM9CP9mOJhyRCZfNsNuW1aiPis9IBAb19ZlypA1CDHfM14wPGGKKr
cQJofZ+I+0EREZClZpclmXeDgr94vm75hGYIinAFkY3nnPzGgndGxvSjC5wJT4Fr5eluqFye7a9W
2HYR0WF7N8zvsjTcjInPMwNdmn/jf9+cpiulHzLUc5fKr0th1GVTV2OvZCByU0ivNh3FEEfK2Jbn
/qWN1/x0dKQEnecjfABple6VTUEk3hRLUC7oIV3yuqQH1tcRBxOXCdaxqWXzeJvxob7xiCDkUDFS
kO8EamVSn0w8NA+vIzFnqJ+HqVsvDUASXwlsDNjo3Hhzy2j/MXQZj+zYGcRijJhv6jhNtnu9sf2j
uWM8wC1KbMKQn13AC8iJdLjgM60+qYwAFC5TV4Ucn0wXKsDbvQxxaC1Ajb+yNr5NRrcS47S/CYXZ
4I9uLUE4OePpU6DOuOarW5ne1ejsBQ8mI0jnpn1NsUXVeaj6akFkxZCQFXu+gtyde1JDK+xrXqC3
KX9mu5wlC+csLps4nNShuHd0SUiVIl45MCBK1yJZWra37K2VJD2gaLPkSfICnYqn1B0JBngSeiFO
tBk6F8Q+OlHAMq5xBPb9AyPZtsQ/kyTYz3Mw6bkyOt9x/fUjRA3QOuOyzRLjs0iezi/eGv1ifKZT
HLRRGBLmK0uu7mY+ahuIcZxlboI8D5wfitIaJRR+I1bracGphCgIfrY013uj3S1TCkOAtOes+qbX
C0esUQ/Sg1/KhcvGc/X5OTPrXHAUVqGLud5mnxuiDvFhfpdq/uC2dr0aOINiTNuOJJTq+5hfGwPk
KyWt5TOGxyDbQPQOwDvPMRNc22Rrk2WUUfSSp99jPx5W9SC1dypmmDqWjfUsKoyo4AT/JlCZfsoX
3O0gsKVRK2kwb3xXFdVJGRivu8/jNxNH+apVrRQMiwVjHvtKF/Iv5w+vKX+v+JceOoMrtfcuO8tN
CHDuXSWK1JCIf8M1IVK9IAUTEf9oh9PdNWHA4K6ReYMi4fDV8jZoW8oPKEFbA+bY4T/a1v2pT+Bk
FctaA9NPx8vlfRtUl6hEM856H78sfi2xYhABNGp0SGRk0X4PrL4DBRJUelPmGUcU7aygIGSIAaEY
7wC6dKM8LPB8zCECapYCj/C37tWkDeeV6go845WKSR0dIzVphSX+g5PAbo6fMYUOmZDu/hsG4DZF
X/bIU+AmgTKskONk5gh8Dq9aNRSTLyTyj+ZO7r++Ji4rbTZ0P9FR0WfarefFlZOZzozIffLDD8ED
4Rky+ntp49AqF52Kx4joXiXGFnB4a2QiEh1ObTMiIWJJ9+kawx7kggpjithbb9kz7GBlHR17YffC
KuQe4c2W5exlLElqGsXDqsmczZkZMt/m9qB7uMUknwArrH+mRD73zHl8p5wWfO4B3pZ5nxOty/Y0
0PK3TaIXldumMYIpSF7V8knWAcV9IorY16s/EesA55diMwxLcHLJ/8NLISle+FlPslhG+TQfFMPs
GOrJeA3tsfstkB8wl62agfOm/qhbsuL2z1q6/6dAFZRWJOfl0aLCdbK0aprIKotK2O/Z8ZqiQts1
qswQA64c+gKfq3Ee28fWEJC52VEwost/23AiWKHvz36gAflJ0OJyFA/m26/lqkylAAPuaJlOoNvR
RrXhWt2L7rrU+7VAoMPlvcp4oiDskLmf9MaOJuS0WfFSkhVo2GYQhAlOY66K85r7JMGjj/z5cPEA
Gb6bTYpsQFWmuMKKw2PM204bvl8KSzA1Oq3FsOkIg0EeeoLBmIOjf/SmlVi7Sknb1d4TDJiF/DjO
J33TLQnimjsshSm1wJUi6AwjeNufV+OKSrfqPHhksFVtt2cme1kNK6/wjlqmPaZ3WDsubf2je6sO
rYeENlG0m6f5P+rNoxoCbEVMmunt038aEW0ZfkCW+xCH/0PtsMtKHefA2Vky/MpY9AT4Yrvb20uK
BwH7ueAGaJrDy6Zi6ktJufwzqyWTfVaCydKWHRJ3fy3msWim6QLE9rXY8QW8Wh0XINz19m+UgPUj
LDi4kmxypKe7+AXusrwyM30QMczuxWv8vShGwGQFHbOVgni2pexYGEcQIKIxXFjpZ6LPRfxeaq0v
sN92+gqsHJ0a7ylU5XU5Nh0mwcF/GSO/WIYqMamB8qPF8OTNCs6vrcZ2o8imsSXv6mFcHmqcERlv
w8uewQtN3Ng6ktnBnhebHx/q7r3ekxQztob7JaQIuRQGqFnNsQa6MVxqHdJ10ahKdIDtHn6AnDTk
vveHIVtEFGAzQWrWMvRNfsoJe82haSIi7n/6S6asJhm7Ma4fktc7bDS4KzdiHae4+SFzFe8bC6jf
s8mC3wGChL6xlDH5Ze9ndnS7TGZWpH3sVocM3tz076VXSnuLb8eUo93sVR7824J625768Di5K0Ac
C16msNTEHdSi7VitCcCyKM+mexr34e8NT6/gcc0FjRsvxnkpC6EKYe1NCIUtDxatfgzprioCoy1Z
2Z12czbn1h/mVmbSrBv+p7kwArHuNC454WwPZtOVtjCYfJcQMzgJD9FlT8jLZ9recXjXvvwBg7Zy
hcGkTgmk8lCViKF9oyiK39hTy4Eu4mbjBTuiQ/k2a648qB5h5r8Q+8+XkXRe8LO5QEIsHLWHDLkh
msj/0n7VcubGQaUxGBbGBU+yQq4ZfbrFCtEzI0GN696kz8zzsYQiDbBwYt4Hv5as1hS3/VR1SGDZ
b3aFu6Yd1ojAPq/HUjE1trjNb5ruU3ciMstuclUjCvAEPiYeyCF0HmM01js0hJI/zwkuuyjMDmnR
N40zdEOzje9gengnGZzPAwgAWjm9p2gVlTMZpTA/O+N85fUhYOvSOBhnhwiUHuvQ8RP6z1shcI6M
YmBi7jwq0oFwJ02Eicy/gT8/hA/WqQhXBYtlFscaUx51Rx6+rW5dt0SVBtb2K9JkMkJ245l6U6ic
U6UTfrF80iVIhERVuDgfyEJSH723LO0gbz1ZJMm7k6NzXpMBwPOytfNnDQEa3hyiFpDMM65I1Tlo
uouuEb8uOOz4YbwdaE89X7MBNhvGH3k+GQQajsNc7QmuRA863V3sxJTBQxjPaKMxADmSDuc8+Bo4
TT7v2VZaOFDZzCaIzpK9QOFy/m2KGqAt8d4pu1syEjrwHlZMrQZeTobzeHtwKuW7yEezKeXbQBwA
5Bnkm5qHSrj19UcngJ8632KG9slaThXnk9da+JqPaPrP7uGS5W/yVLlQ0F7HjPrDS4lAeeVHN8l7
hIpzNsbm9QWiOVK0nd4GtKyWDpEsnJckPGacPzoGSPnOzsIMxuqK9kaJtuXcgKu+L/jmy8J2BRK/
I1HsWONWGkwwpaxkqVjh2B/e6FJ57Wwr74/Cbk2h47nEYXZrgWSGeugP1Zaf3PqsZrDkzcbP3Bnf
gl0yukeQEsxUifXNt1jK4Ga0/XrITJk2uFyi3l9RhQHOJJIl7pPmlPw6xO90oJTja6VLIs3nKaiV
qN51LvjzGssVXsT3b7v5FdWW0OluHEvgJnwPm8I1cML1rV3VStE8SsvU1jdjNYKNCPemYzxYAu03
jP2W+7NRarxPfX8yXyoxlCadGxMYExynB8iOvK0APlIFBDQ+Kg5q+yAueerHPFK/z8vAmSy5c7ku
WOzG/N5eVf8UTBWvkOi5ca8I1KmF4uDL1TKCXfYYx6ry6fdh0iNkG7tI6SjN4fazjNd1Smh3Iif/
wm+yBsgu00LDRv5RNVk6SwXFRhMFkoNcyzcP6Mx/PPRtjm9NBzatX6zVDBJI5lzzQ/AwKPT+sV/4
rfk1svxIPEup8U5J7CP0+k5Blx/czkC8q6t8DZ5efq9tFJ+mztdXf6K2EzUZ3MBck0auYK3OEyoS
ekEBSQ2rpBQq7cPHewyr+FOBaj/aGyMrC4pMYCjE+X9Z5wCvkxALQTtigw79tdfMp1YazchOQ/kV
cmNnA0F6KywpvjNeYlDR6rprx+SnOYWfjD+/5ahcomkYWheuIVnRFEg8MTHTR4vp94aF7aEQ+4h1
tx6dR9Q9z90JprQM+d0S54CHyLczKgs+6zTXdWmFyjJtm81QYq8i1hB37RwIxZLX/LptwSPbmtL3
aN8RuoQ7ZmGFvYbnhvmRplMhVo67uSQLLRicylEvBkaaoFbSV2IBFrb9kRHI6aw/4qw7TfK4TgzS
sGWspjnzHqO++By2D+VOFTKDOvp1Do0ut7p4pkdsCQmFWy5+qx3Flkr1CyqDw95LDB3BppyJaMCJ
GcsWUo2+nDDj2XQm9BxHwcG+z4qvL0hRQaTxl3wlWAH/gAh4SA+/+dcl5b7JIwLMt0fa96S0JFQa
FBojCPDZaVgs5BdDivRP7XGNSo3mQfcS4tA9929z1Odc0wrGyo6qrV5iMZgAzUHokdeaguDpJMy7
HxH5FhjCYbbJsqBL9o4hl4QojyN43xr5SNX/YD4OyXAlgSkUrP/D+XxBHXrR/WzG/FMY4kkX9A33
RrgVA/qbr9bYn9fUyBe9CkVblrgEFuMPCSluMlgOr4vKVRnmGEZAFUXxjztqwPXPkf1/bjfVabnp
Lx4avnIou+LQ5EPA2B1FoIp+FzgTEtX//mG2RIdXjsvf/Jbq58NEWpDrI/8HGS5fBMpnwNKTo4AG
wJt1uMDPKxUiLEyRV5wZgP7ag1oX3c5IopuL756g/P3RCsdlV21qqZCedQDrEUoEykUJKgEQ2MIA
5WVSgfqZsJD3hg80N+Mx99eUVPTs0vcjvjc/uqah2tDHZRpsbh2YrlMobMd/liGEnMTjipPp34JS
b2usEEMBuw8+sf9sw9y5Nl7jvhOAhAiPyqf7YA+zBNA6Ii+zbaJSlsF2y/B/r3VHcfDIKNhfPBUa
IBxTUbziwAGTOnI6Xe3Flv9eruo5uB76gbY8jkQIo2gYZJbNmZvcsASB+s8RXWp2kGVufgIMcwMr
yE2McaLWuvGt7sLtHk4z1ZYAbIdQeEk03I5XUfxjySNQ+2Lm5cwgRZT7v+tcsHIeH39ZoEXsdN4B
XQ1/b2DkGQypeMSkpZDGjHX4a5E9A7Xcy7eL300xSeREnZzEOzSubHKxN8IOWQHTQu4v7xqGiOsq
KVNvYkWPTGe8BdjJPdIykijhU6i4mcS+WZ9ycB7NYPLBx8oerLcz+P83g19Zw9sfCA7DvkDHLuNE
15jw0d0VAwsudiFZbjFCP8e62cAhQqeYEeroY1GMVaC7kRVe0dXXnbOY1vj9a/k19pbW3ib2apvH
Y2LADWrri5YGk8rSJWZvjRsVwj0Ujiw01BCCWQwiYQNWGD+3CcDok9uZpSJ4OCs95M2qgTSyDVOh
wB6DB4vg4HpRx7oHJi5SL8FNtIRuQC4Md9QPoAPuojFzp4pveHo298bzF4cFHe6jE5fegV3vexji
N4AHdlxsJx8HA+rrPTjW/ParlqpJV7knGmSzNuIQq3EUI5lRLzmBHmQgUFmB19aRaRM+WHPOjFnN
ScOhLUG6LGilVX0n8g4L3F3YEZ/q3RRj2wcocqxyNuBaD8/8U5bbdoNQ0w1rITgVDIXSQl8WyP2r
v35zyA/8VN0qyUHZ8jY+9Q2zGCIaC19ApAblipFjEqfFwGtfCBmW3QoHhJSNcf1ejGCbQ28I0qxg
doLsuWItqAuM0BigHA+6mQ8zt9dpTEsGIVbzgIeYITjVkJ3tW4WhZLcpFhZtSd6JDGS3/Lcd7ocq
tWSEQIpvxxSL+NicwXuoP967cbsTDvIdpM8aGJ4p6DzCn2LhS+zmuFjKwtZCFN640X/DIJS2yRGa
Cq4VyFCHdniraUA7Pqix7WN51rEuTwn2+4hlo+UhYAjqg18fVbAebCCJMAX4Yo1mUD1rWSfXamnP
L8OTENhgS4IzTNWZW/JqHQrjHd0ridUKMnXHP+N+vc6jLqL1ddZ3HH6wcvLqeAflH3QzEc9b9IGO
6BkB2wNZ61WUcC/aaEc/JHiWGZDbJZ003hcXFrdQrj0X91z6+A3eYTQjezwxb4iydGjupAwyMHg2
9YmnyGtTeYrogbiT4d7UKR8Q6O5ai9TUnD1cf4WaxwMZwTyihvvXFt4C6V2AkqxI0041IVvVCkTv
6ye+GSuVxPe27Pp9M2QkKSNZEZ4q5pBvV7ZxrW10w8wxm0bI7xkCNxV/sw3+JOSkDWpuxsgeIeIF
yYoNvcgJUAZa+AdVtjqC2GnPmMVvDCZlyqSygbEyOZkgg14v8rxsoKONUX+U2QUoVaUHkx1PxX8O
Z8whPivGMtuoAxzUvSKKPuXKXPwDb4MvV8t6H4ZPoLfRrKS7iRvsIzrcpXLQSSgBsC5FQ9ecvD64
3zsfsXWRVav6eJJohK1eI3Z/b2pkzQlkigDjFD6TCkeKuJfbyFiWZ4jwBMAAjEcaYAz+Gobtju9m
w3B2S6UX6Q5b7eNgoB3QxiDy2Ib4/XsyBCYK4vHTEBPmEzHYfDLwYzWUh0wszgvtSwti3m0HFxX4
TtIYWE8koCBLZA21eaS9IanGUNa8BMjUvgJ6Hm3+FB8JUbbOrZK+ab9MvGE99Nfr2dVzlKdKQe6m
pAYqsDrdjwwci/adv63enmGQUJkr5KClUfCUw8bqxybisrHZELZErJ9LaPmc9+6/g6sbgokzRq2/
sDCQgtZ+AZH+M3ImZ9xp5f2eD0yGmKG4wHYSfZMkIz0va1TfoFC069f4U9oR0PAticEh3AQQxsOE
jB+VhzirjPbNJ6+0jY6Tzs+4LYdXbM8BB2BGLzCRNnhv6FC+sJnOByK3ItFHgvAPZm4EVCTvkSrC
48lWaUG4Ow1xwmP5qpKbhoHXslp7lfKTgPORqEZP67cKRoQiVytpW1NpVkSc3f2cQOeMF5g2Wir+
roHzYNdzdmRkxErd0FoOCQAPG48sVvEG0Wm7eiVigcXGZld8qk63456kCuSCrYOl/XSdG1PDFGtF
doEEZloM68mSyykefcYTCIKXC/I9tP9B2deVhG7RymcwBCLZlGQyVe39mYWPoik2CyiDOa6vP6lD
lk2Kfc5Lh7sTx0MmSUx0bVSLG1CNg1TihBIjU42lV6yp/m8F3MoINpZMoUqu8cRWweRbMGyug6nu
6ll2gV44WLV67JGWtOMMfWBWPcIW4H//QAXlMrhSDSLsquxNZd3MK49lYRkc9S6txr5YfEgw1tTE
r8yR4luRstozVk1B2PqAmno2u+TtOj86Fnn9I8xR/ouGZ0fQY/hkPPirVOZW0nd5WHV2fSWdWssE
K3jrt2ejzOSPjIU6UrACcC+PkSVfmw1FhE4UujnLCAA2qvBNYx8WoJQsHFP1npOZDICK0xG87chx
2k5Q99lbMCQng+Uorml1g8zb3+JbFjYWX8IiH/vMy+zINK/uLzolyo/tKmGQ6x8dWUWqn2vhUajL
pMA1dibw30oJdgPAPouLq3lfFEcpGfRmkokkIt0/MZ1YyM2PPXxvEn48ebTivEgiQ0mzblod0WBX
8waWR7m7PE6EQAmk4FIQPAJzOam1xjnG6xHLNJ1JKHYM4E+MpctQNaPM1RoaGc8i3+yDcCD3oLXs
KS7mpRJo/oPrcflEPdkmD8BaSqRVPjL9YDtv8wqQXIQqMzNknqiM8TKq8XGdUH/1j+xKBwxSddnx
FedS7agYmBlWqxJ2Q/61qlwQEkj24j9pFQpfwPsrWec6+GtmvwtutokX9ARBS8w0A24z4BA3Yfim
+j/Xh50RpoIM3/zrSSlTOfaykjW5TH1cpEg6kVi9pTUEmMD39zzbCKvWzCN7++k9DiLyr3FsNskm
s22nVzA6m54fGMXOZvmhfn7m2nT0AxkIBqy9PbxEPnKumK6MAzoH2mlOAYKRfi4ak212ZOJ6DLF/
e103b1SI/zcWOnRLDTokXJY8IWf3TYZA3/Nh7tUGHqFktBZRitT/Y61G3O3LNSq68HvMsPyiSH6x
NqVY3WdtSHqAOALipKxzpA8V2Mj7RypvQDa5YtVoDO5B6h+IJnFf6gVDCqNoKFzMrgCxPpmYusnU
6AwuyrEtdEgNwxTD8dFAUPpa7WouuHzOaytaBFLqfui+I6gS7tbVNK7vRpzrW3+FLpJ0uJ5PM8pw
vozQ4yCc3NU1yJg92Dgr8iwLR5Jk1ABUSiiGKXAlD5/F5R11Bgvn3iFsAIhoC1Bu56T1NUmfZruz
OyrkCyRLHi7tQKYEM4EvVrYmUTUWFGzyvym7Wyj1LDIVyAvfeICV5YwTWEPq7WMJSuEiL1Yr+ntZ
9v2XeYm7nWjyEQQwelYKrMwmEfc6x+V/JslF/UdqZBf6df8lgdiPyRiKcAcgUJgfBUWU+vVs6yZS
Ub3uwEitGSu89NxTu3L5BSbbMIXEiBm0f7U5cwDyLZrYTpbyLfdV1f6kIkdwUq8hFR9Mc9hw+/Pq
zLxJrWseMZsT8+ZjKqmnC29KbXtdb6ig8YT6qUedpTJ/ElRsnN8mrXCf2T7V28+j47WDW/29t+dR
/UyaLsGrxQ1V7LAqhWha1bgP1bRb5MQOQh5GlDgibFMBLx0zc900XE14pqvrINbusVuMMRGpLth2
1e5a/5+K7JIzeP6rvmoWyWWl4Cc6WvupK0bhpqE5Z4jb8tLOpuwCtZorbHXIePNn92IhQiYro+MG
8w7bd1ONqB+xI8wPl23dOYSSYfZ8zaH1w+RBKo1jNe3STx1ayahCajKxnW2V57D2XMu423leTKxS
pw81czLQ57RiEt0JjCoG0+O05QFQJokoIuAQOsqDeb02zcjA9KoTKwzHBcso16sZvb5mi59c5tNc
jehf4H+WyBSvoASLFnNtH68TNaZ9bIaFowlExkX69qwp0cKq4VhPFQOFecVGAIIDZ1P2byo17GM9
p0ch0GmmE4d4e9Xjfxz8qshEvj4oyqt6jKMPXHBhLLkO5DgUvtbO5HNu6d+HnJhC14cmQXgp7M2d
Y9i+rg1wSTd1xm1pi0aS0tqaD9vU4O7xhdKK9k7BJ+HuT4bhZqZYzKWrUxZkD3DnES91ulRwo5s0
lNEHFUgTEj/TsmG4Rh8vJFlp0FOOdzX3Nu2dj19+XzwEyVuanaiOlAcrQuMAAHgZPf1R+zxFDf4T
J7M4Or19E07pHQSNLCuoLLx+GXbpjIT0rL7KJ8OrSU5qABbbgqp5tDEHpO5a1rSE6uYxfE7hkXyc
3mRgjZQQrKIbtrsrefLwG9+tVqywwQ4NhA1esBfsXtxqaEenL+AEdSUcStbcB0hR1i8lj7f3uCA1
nCGoxRYdFT3gevFyHd0NN4TaZvRg9l69MKO+sDbEvDVB5jhZtZVDvWbW8kwoGRaI/2VojXw4Vwp4
H6FaCkBslikisY0Zlwpw8Eqb1t7sS0Mv68VC/8lzAQJSrpn1xipVHHnzxhYkCAEpZdGAKKgZQdu/
o1DuFnD8BcsWmR4bpknrpme4XkkL4dndMjx4ltrJs1xLR90zcfYFG1UWQP9wTP0W3ZBMAJsBBg8F
X9zEl9qE0sgRxts3KzQw8BGYroQxFxviReraQDvwzH3sCt7WYg0iWzCkTseWge3nJM4WQDMsVmvw
T3eAJo0EXuYQbWw90Mf8mmXGXkwwiPaGSK8xy2gXxf0XZ/jvguwDU1R4NgbAVzYRggWPtoFW7k6T
9IQb4q2yoMgOQKAkitDzv8/JZfjv9r/dPo6nQ8LCnr/RobuUyy2UKmHoyI3oAUjORVVL6HcBSH41
MgUe38USu7K3Y1IS+Z+9GMWwZ6cfHaAxK1cKYCTcgXGEh4+Luaml0ZUpRZH01HlwURu3DFvERzGb
hK9JKHhPR4Fqp3MvAVRG5732Y+OjOvA9/UIyKRn8afDSC6g5Kqu19sqY3ax7mo9k/zNrHKdPrRhx
cOP8A6tHlFvxN+t5TfAiuvU6iXvE7U8WQ3dY8uDhkcckrttdJxzzyJkYW0H4ef/HeKdmpl6CRz1B
l6JCOyq31tdnUbrScojwYF1wM2txGu/BHbwzTfN2o1N2xqT+c7TdOr3nvQWBK4vuUtchnr6r96vd
/KlXXqdTLoATufigZkJ5iS6mtdD6Sp14ieIoUZTlR+lOTLjg8FN38I5e+6oWHi8Ny3tbGgomdV7Q
ebm3dRlG/Bow/x7KbOzDbFWCJGz79dtkTlbxHPlizfFoBsWMRvhQX1hu1nAQearLxJb7N87USZPv
bx41VBXE/+IQzN3F72P3E+E1cr4n0jGVmr90lUhmEVrX22Q/x8P/aR3oRkfWp9Uvpbh4Q5e6/4Jr
7KaTd4sb9zAJh8SBywiScvReQ5r83odeqvezcID3pk0LHm6vAJZCmW3tcDzZW41iRFnWSrnGIQyQ
tjG0a7r6SBaM52EE2E6i7VHj5E7MRMpu0tJnCkrjnYxx4rQ4ziDiQSPnwE/TVRnq7HrdBsoNk1Mq
n159xlTeJm/arXS0dwsmyinL2gtVdMIv3KEdn2F9zw0f+DrIRY1fsV4M3UN6wLlj8xxeaqi0gAhi
W7+QxTpe29+uioVxNdMPOp3j6khf59yBWJX/pDhq1KaIJjXV4Rricu0xWNSj/Ufjp20Jq8VWTSiN
SpHHW23eoQDjNqlbvGXjviGiWMo3ed3CmFncJ9+bKHsWH0hKVfOSDHrHg7tbf/4cK/GE8Mg1YvcV
ywZZ/SZ7/wNDDZk5W95RqJdFwA1CjRkAEiaJSaZZ4YZS+yRWScvEWbbdJMSwctKK0cpKaNVJiHxS
sLuuTqKPWneXvmlG9Ymn0vySLXzvFIEeEL3Rl30Ew1NdvT63L+xZG/kon35JAzDNSzSLva/YSnvY
70RTD9bmZl96pQ5k0IPZxSjmod9SMFhC9cvbgnXykq64wPHYtxd16CBFhgC4utmGtl9SKgVRvfOc
iZ5qv6VDhVp2GWCa4ERUOA3qRPYcQUJ7NEW1RBjdcwHl5T3RQsFSQnk4GRktNGKrAf6iZJqoyCAw
x/8T1aHoEkWdx/TEW/PfvFLcxFszuY4RCn44e/qEZDUevrgpn4rkSxcVnnAgvHKrt6FB2zK0xzQz
rfbm+n0cbtqvdJ9K+O2piO6HKDWFwrBq7u+FCZlNpgymt/PEbawnk3syvv3xBf89jWoWBdx6sFl3
ke2XbhY3MyvF4p8cC84uj6LIY41S0ECvmVS72Gwi72nmECrYIiKrlajm12atscqMHhbnzgD4tMby
IRH1o45NHINkr43gCsAkCqaXStpCbWMEtRMBAD7aee4NfWq0BiRAXz2idhFwxObKqnR5XFt70vcL
KQgSRYFPvhnk5uJ4Xuwo547FY4eiZjPvtUJX3UwtWDeschHnHkMOy+hYPnvneQu26FtohO9JpmCl
TJfGRid8qTiJ2/+g7IGG3tgoXL2/37Apm9t8ZokVxvIe5fify93AGUAJqh7xW5oC/AbhV5IURVA8
HwEHjZNedlisPqjMAF0sKefM4wFLhq1Cx4P8iuRdL74VO/9b7t/ZrVGdj6L1V6E5dwIOnRh/Pf1q
Yed+iRJY9dK/f5otoXROYcVR2W8FscrwoEH+jbB4PxNIUf+vq4r7Cwf+QsQnlSuz5SNbtz+W3pG9
GbonjaLHju92jusO560GATkALBR8a9cJchzgZpIUGS7TVIRJrIqDzcZxtgLNK7BcZb/QYcEs3krm
w1BSQqI2gNUZhwwoMmiESzFktmcmbgu+6/wAbmS7/NUjhgUfpBoy6Fj4+3HH4DDMHxrtA23IgY69
8I9F9X4+a3ATewNXlRf6hUrJxYTzfpfGK59J4bgtpQAICdMPYSpO1Ad6U46cm6g2yvnfHc8Kjzc6
Ms8yM819zbGjVmP+vOVVNdFXpzocVNnFbNFUIYMtuvj8JB7OIednyQ9riSVsS0BIlUps5rbE73W5
lXd1DSMgiq44DVlYWkDCA9FDeOPCG1wZotAieydQllL/7nA1+tamgH/2SxDm4x20BixGNJAjv+sO
2fMShydgilIzbIQRW5tsg0dqEHR6MGmCxSSKnvrFSPWQIpjFlY7bWN2HlJYFSA928Uv81teJKy4a
PDcELqdPJJnRCRFD8bmqxIYhj4H6YbBBBxsbt9gvwwe9UxQ4l5lGjPMnDxatPX/UW9Oe/YCR4wgp
STyxPqpVDlS5u49mQwVlPwQbsAVodn1BiaqrwB0QJNl6boAav/Ay1DdM7fQo+eMmiy5w+lHukAsA
xV2T37iTt5hB3Q1u63u3oyxL0oBH5b8hfuwai+ftYZ2t8iZVhZFmOni/3yYAoRgyi6kGW5s0fRnY
LfpqFyySwo597nnnCcRsnqKjrFsIQmCJZRa4Peuxzqs/Ri98ueES/xqvEJ4wPKDOzcRZZUcp2aZm
KPiHhD1OkPQh3mCyvMXGAUevW4ca9MRZTio043FvEkRijqRpMTGFyASg3C18tTAagQQzlBBBVjUf
yDAh2YIhJo1vOldvVv0JnjRV2h+XmEOKXd3Kgu10pHgjeiHa5gGtR0UeUohRF4AEx9j4Esty/2Qv
i5QuGssPu2PGQ2J64gpO9vt4OM2xX5peRQVaBNLRo4Rb5WLWfhocGyGvGBlan9T9AtebIQOihwbU
2l59kesMhpUbtd5N7oQlPqFE6pt/qNJtaonen4S75RggNOEJHN56qaLr5C3WayUERMjlOzjU/eF/
c2fvKRCfB5jRkYLl6zGRfHDeOK8glhsZSluiJuS3Sb5d3T+jHMJdfL88Aly/4fdYSvTvN1ZcNIkw
AKCyCpNqVKyzQ2J7ib5KcUwLwd+NAybrD2Qoqgpe3atUYRmVk9aiOljLW9OR60h5Vat4F6FY9eee
jZYLl7GSj8ExGgxDJnwmyJPjJqMpBQXLKVaHSX/Tchnh+0uiJ2TgdOhvh5VbhCDfAEuaTTdaTaHG
v7UX2EH9BIG8tcDcfx0GMfRj5YQR2fmcOoSgAX7JPOYPnlVktfg4n84g+fyt6L1djypUTLscEAfl
ecFovoxRS58x+7BUOTU5cOnSz78a1LgP+4buC5cSrRzd6BnumPSgIF+Jw+kd/hW5bE6YmDwLddpz
qlZ2HD0ReWmQw25L7fAnZ13P/61R6Mdk7rPMUu0G2mZ7BiJcwNwVt5QFHTF5WyWfW4HHSD+ERpr7
jKOEAOtiIT8ebevEf3U1pwU4Gu8jTt5LD28blqrY8FxOVyR7W4vg45daTL+fkuRXNFqyI11Fxoe5
Lwp5Nd9Tklci+CTcVMSPMFN3v4MQLDsIrPB4wHUB82VmiPF9NLtq6vSDu7S3FvtgLUf8auoIQyDN
eNJgATQjAbPtppKhb+m24QNJS08AqFe3yo9OegcoG2izfjZQD0kVWmlVRNTKLeCFZ2+qOf6VMSok
hJyPhThdLzWkQLKcwqxCZyobM/FuuZF9x1XtBu/TjlEtxvbwNG+1zQ4AvaMyhFHxQoH0zv0I8m2J
VaOYVUGsikBXqebem0pI6trdudEdKuZ6TQGLflDB8/eWWhEylS66QOgHX8QZc2pb48whMm+6CMA+
r9TeVEpkRmgfYetSTZ5Y/rfOtCYRh9AFKPaz+lkn0cwev1ojTCV6Y3I0I9MTylKgufrBHeP6qL6n
l9rS5lJtm5cMfoIh3qk/HinH/j100BUW8DkvGj/eAPP/2K+A1Bx0Xi4YVDX6n3+H+2IWkZtoBvqS
vGxgEd1SjB2MKzfT6wkmZE0+Kk5bg07T0w1nzcGG4UntpXR0VQF+jgBQIOZeqUXZc2KN4MTAgo0H
CdVJAEBT1My78nPgu1dPldnP+1t9xjgzHy1jdTmxcgzkV3uys7SmxI82KnzT8C9kEj1ShepfGeme
EUa7rPTcyfnOLd8sjoFh/A5XJl4cwWRX45W6RZLP9Bm6WyHAC18kk5GYp6XP7esAGSzQv8m0z/qT
kaep+JE7ZzHfRBhdck7NusTEmocWZIP8A6GZ3mpHNRU7KDLy3iKEJQNW+QcPX4ozMekRXX+hKCgQ
Vawcd9v77Hflyk+OGPAPe+t6Q0lUuE3+qU6IBZBvXWnjZByA3SldT6dbNd2pnZoJLDLCUCsNC6mx
lC5qJoCiUiGgAIYESJJUhN4AQWn22sieQOkbphhXIrdf87iXON5ADWv2vD4yEbZe1vGEP6dg6n/J
LiOv00uo6VZ4rjmKAJR5xT69RTge93MogfA5O79T3/sGI83ISG7RbEAkPjOOEPEsFEy0RJ0DYMFs
+3Us+L9V+xbjnJfGtMqOz3K1IaJtQ+6xAF8HVCCHmv/FnZQ3gVCNTDzBM9fNP7Ks2qRNyc/z0rBD
O8UbDLe8QOr065lMM0aKUsQEcuzt6zLeVfrVV72FG6Y4a/SRsCLJ7l0NWPkRY6L3osOHNAJNEDrc
OY1qkABNPqRNcfJZAzJ6n73EImw+RYyn/7tlBI52Jl7zMH0SATxuizb7e+TCc3kmbYBErYfTUx+m
X/k3UygoPL7j1qzwNg0mW7lk+y0M6bpIZ7Ex50TUgUWug2yu7SS4Fw0MKaDW0WeVRPftxBA7PRuN
ctx70opg0Qiau9nMg0565VohZafO5Hy9ffaH3dGze5ICV06j5uT+LCodGQPMr9aX5Dd+WP44Pftl
yXICwuOYY0xaJsV/n0V/LzqragLJ3Ejwh6qJTwnCuvHglyqyPYH1ZcX1wMT7FESx8pSeuRTrEWMv
pUi738lyE2ooUlDYGu9bqp4dO8tGBuzr/pOkajfXGgzFA5o9Hod4deQVO3dHG36Vymo7OpPkqlsz
JCVDwvK2Buc84zd5W7YqZWFZz+SBAZrgGfFEIj5qv0u3VIYvtIAoYCzFcm/namKkHyEsYb8fYcFK
ztl0/EDWMTOSg4ElRdGjmQhfnsyBdxZSEght3k6/MbAxobbFSp90BXPDTUe+dRHJZHbB7z1aOA+Q
TY1pHH9S46VkQntumrjZ8w1EM1xgsV2byqwaxGilJYrC8wxwpSadKiRwxjrmvFJwgrwrkYgzXCgB
/F3RDkSvsflN8gv9G75vObyzniwpdjigFdga3ZZ+BGGs5DSJFbmvfzeScz5xt90nM2hz2HlbAOCm
SMiLCpTpnYUNAmhSV5RZuLBAQDHqyy/l5JXPknHVQIYohzyJAQJKu2ErOS5pl+UfSAFYWC9IP3by
9pFNQu3oV9MQF4GDbUEFulbQROWQZr5ghu5M1c9izm/wFqLOicrcx8eVrON3LTkuBQZnqHkP+kcJ
oWaNPGu4OhjNv023nfhulbTb5+C9la1OmDvY/TmQ2ryGWpFTLVNzBI+BJD7jfOzxIIq3dFznR+Fn
8ZUrRUYcFnsZ6Pzn4xOjE5t9DyOK72QVCOyGfskD4X9CQN2JcMUSfuyvEg34vf9swt0VA1ysSTEI
HXs2mGCqH3+Ei1sfDB9PFz9hc/0ff4zqjMVPh6BjqR9FziQUgR74PULZNlxTpTvqwtJsHe8mUenB
AzvVPnZWRu6oHssmv9BJlqMEclpd28mqaHFeb882HaX+wm+xjPbuLZVRq1vHhNsJRCOYHLcOAECx
8ELq0HLeY0tMajKq8Uoz7CndVysIyIepslPTNzgn43hNNA3TM3uTFX/7RGXxmuHLc12qcafisz8c
8oU6cBurCyV7dr1Ku4QLBhNliX5kL8TEZh1DB4UVbKuepALj1jWMandDgEgxFyjEGyOAGYIwjtGm
VBbujI6yoilFDllkUELhPcmVq3jkFWQy7lGulkA5x+VByIth3RkA4t0Ulwuo7ktD3ENAy8mM1r8t
Rap75Qa6OKsR0q5q7HL4NrkwNiC0KGhV5u+dZWwQ89gFk0Kf1UX33Doijx1uqahUpyAm+pv0wX0g
Z7FTUvAdglOCTHdb30+ZSIO8mYGMBc2XJuB9tta5HahASuxmGs/HGphD/2RdN8PtIzswS/ew640i
0EWZ7mgfRii10LuvP63UxGJB2/tEFCcIO8j1HzO/viFSLiABaHKgugNzBEMb4Y7HVawWYVFM2LUO
pzPmL2Z+WLRm5BZGn/ysMR48ch+Mp/Ym/oXTMJgARBVhF0lzaPGhdwMZ46lw+uV/ZvWjzCLC0V1o
GkRcdpWoKZvpUKIClQ3hZ+hyVCaKHYwYzg+zNy4Fxn8RJiYgUYX/iuPIsPz6pqXyJNOS1rdAVNWe
UQUMe25VltAg4v5y5pkBNjbPk4/v0gtRPzFuhuv1/20Lf8fsnbzM43RRa6LLHBeFI+RA7elO29k2
CPDaGjXdqM2+QdOMHpcvqkckTipKllZ4Ptr7P1YA2LGBt/VrESsOqwa28ZBoqOu/WoAUj7Na57TL
wiTI/oD3E0JadnRMbCjJYmKEVLzMl1rqiU4JPsL0jHEVxazeNnLE7gFOLnJsAz3bVeDnGMFBknDQ
eQ6E1gUCmi/iaOSZaIQxeT6V9w8X2Ov5oGbP4qxj1kHIXW+J7plxajLyeZepm1lpFu0obXv7qBvt
3U0DwTfORXc5w7vpKUBnwW25khME0qMYuJsGkmO3ELTPHFPYTFo1E4FGjqpLuSwe+ps5x25yczOC
LkqcGua2yt7sPpd0i7Ho/Aw7MYMUNtpkwr7I1t+XkftiBJq6YwLPUBF7u6/tAKIBFTefyfFxzxwP
dVJPgrBmyiMLxvWn60YCgt3ji3KI75hW7yYRptvzD9jDD+v4tkx2JACNu3WKyMTXbPIHF0VmjMFj
3eKNSKrZhcvnjSWwhOYlIm/B/rSQTY+ug04vKSYbbKKM+Ka8Z7kZeNqv3EJTqNSrY6pV3haHhgD4
otsoSOVvS1eF8CVzZLtVxTCHJy9DWpj6FUMrLSfAFOOe1AmbAbFDar00ZxTCweJvksV2D1k10TZg
LJwr/BsV3JIbssn9FPXEwJ0cD685O8DTCe0De/JjgCWPtL/jRY/6sXyHzpQIy4mdGq9u6N6BJDAx
kaZthIf3lQeHNfDeKpSwy2z+mp+CYUJywxEJ8UpbeLYQsArvyGujUnOiCITLKWsBQAh6KMI+A6BL
KnUCDjpleHywQu3LLua2oUfSx+z/T7bbpAbcIVMO8NYKzJThg8L3dZ+uDZ1J/hEBl2ULz2+nlszP
LSdnyh2JwUaLdQz47TY4arKJPMH32MAhmRbcULn/u4dMr/h+A3frioiExcItVmMTza5V+V2oDHXJ
3VcbZFdyJF/ykUnggmusyeDfTeHohYSpu6PteFOx5LOADngHc5Ki57CL3/8ZPVgYrji5NwaKBDdg
YhTY9sBvDG7IHBtGVU5a2iy+DcDbYICs8wj4A/5WfrrZt48AdPVEzX/Nd29puA6D9jV5M3baR/Ic
ZGOwOPCcSCm2bdVOdHU5oa7PEZC4fD3xxsg9HHt0mbjxkJkMhxHNlB3MqIihY2FLhzq4MpwqSwqx
16Hzhmd3X5LIFW5Rxx9yl+GdWftyKym/l0QCll15dXdaZ+jOMe59+3R2CKfRSswKHbVXAX7mdVn+
CESL9XaVR0Gf2GBWBql6jhzax6jyyUOZKiCcyp4B/MFQR2fH5OejCauFTPCdqjcIVmYC0yvqJT+S
aMKRThihFaH+ncp07kNsGGws0mAecQflL27bycTSXcudq/iPnDalptUYVCYeMKvjyBycrcCcuJ4/
T2SDCvdj4Cq7TDcz0mgTvLShXP5FX+CUlxaMySW0QSk2Urj/vKQpUZaCabj8ByWyDZRGeVRlVxAk
W/TIfOzWsjyoK1nMBjC1yoc/farN/MZVmQdl46ChVeL96a3O1Bod6z0Ofb4rRaJKjhorE6Ov+x1t
XxE2poEixpXg0j0GCxUj+cQeNzjXE/W3mg8S1VC9XVGallxgSTgpwjTVXTbfYXkaXPBZqVx5Nyzl
ANV5ayh/ze+4SZlqZVS4aFcNEIDEbw6k1hI/Xkzp+KrelwbEe0MAPW6O+fEfkNrOUL67YbKLqcHN
1SZzLx22CqRL00Kb0QLXpyS40BEgsrh5cwBlXN5ogz9YpQ8nlq/5zcxaSKGjGfs3B6rWLJ+Z30k1
Fi4x0Bb1phd2q3kqNUTvsVUhEJTfBVX0ZtZNEqrNeP06x5o1Mx/lGWLGbFz3Q5vS91tYt86pn+jv
yckSWtdOkfajYPidd/1zOwuaanV4tv0d8fDHf69+Ev4dUCviXrCE5yHWVoIg6QQhIW9BvSFKljZC
pzvqofJyb9pvQwZiXRlj0n5c9NkMHcewPbgUUeB91YhpXS5gTUdMMQIaJLSHpqPKoiqDPsJ9+WUi
3fwq12kTy2I0o3EqezSQosH7/j8k1+cwnI3s7LlGk6G9DqoiCKMpw1CfDn4nJuLJoVDIQJklaiFA
snFFNq+Z1QWBOKCSG29qYKsgSDXXMlN1YCN8XsJi5j0VlOoEvoSlRiod1iQp2NL4k8f16jO6xkae
J7si+WlPi/BVJB8w9lkfGrNAj1mKbSjjolJEHMbqBsDapwtClbWCG1Yyqo6P3Rjn6NN2BdV/vvzq
hIz1yYDRcqpV6SR6bn8XLMJfR/LmZshl7FwoxB2drpDAb9LWDtLyZppNbSEjmR+jisWiewpDCuT5
UzR3nLvxQHOYYnQY+MzWDA3T/WI8y2wM73u08LB0CRLCq7YjPKg6ay+zPQGNassrgtLApHB32Afl
tmNXyGr1qnolBnIFzXkcDYPFLIco0UGHFfuK+ZwdBL10D1uG0rAJUr9iGluL2tSp4NpzMTsdrCN2
3Yr3kUrRvbw2T7ONomDjag0/jrt91gf4jeKz0qgAAnh88Jrkfp7rOtM8Qjgxe2RYqCgYiqVo/quX
CcwY6f9e0X8QelOjvZWcZfT/F2thzBkaYFwys9X+T+a1hlkGYGoyNl1osoBq2vWpSD42u6eQ6nml
Lp+RnsyNEn91ibMhqyizGlg5U+PLGB8r7ge2Yo3cVhKQna1rF0VQYV+AjkHpb7VwGa/fJcRJ3lrd
bEbPRYwXjGS61PCT/TTXGkQgpS/LEW/1fnG83mffygzS6YeDtqxYqDxaNonPBbx9uy+W8eCxwYNB
fSyISHu69QQwx8rSCalFbfO4omVHYskp6PVOPqn3ACXXCOXkdJYxcKeDr3UcxZ/OCE9fB62zpS06
hOWqI9Gpbsz7LbzMMbNu+fWDxJ3pjy84NYxowefgAkeUQUlvUUXhKSAkj2WKIN7xQ/Dd5zzSfBHj
ywiZ2LMpU6obhnlGDYPdJ9Oq4MFeXTwtvYbRbTfRQ/QXXQOtTvuGtpASr0l2xGkqguWSoAJXGNWW
xPFMuxWrC3XhmW3xPAMGouQEdICeIMvb4kah60i/NBE7U6NHZ+Ar8ORAFCQPiqI19/dVOG3kcp5c
ArXmuCjVZifVIaBRHDKJa/Qn1ZiJqMpqONh/k7V2cThuM8ApKMw7ZGXygzjR0Q5bv9rm85CSyCnX
7Mu0hFTmafRKCNwRnWncLtvvbNVzglhx2coNCGHPp8CYbT4+Q8+6s/Ro0ffCrxn2UHog32JRsPEf
pW/3oSQoGHs3nx8URx25BYbZ4/iz5oPZquU3GXPIxIPQr8N57hAFFsnhIKAgdzu37vJkUsGhwXrF
Ma1RInB8mHxedKHDlLvecv3HBgAGInGc4mHbVRl/aMB7lI1Nt3+SqXX1XiK+rPfRjbPidy2TXguw
0eSNv57RouZ384BxB96v8m4/vD2UxrDUbqVXBCnQRfx2cLyY8R6Agj2GkBWyrFXj7AUHJY9uCshs
r2OZ+GcmCwBPAIxP4Gm+0rwhutL7l0X2viekjpUfPdpSVz8Kzv+p+fPTHEcmOyvleLqJi3ahhUOo
Y0zNi2pdPD8BJU2fq1VbSb6d2nDgOmLSX1qaOIwavItea9Xu08vc4iB0IPLu/jFGLb89oCbP3WeQ
XFFUzYJoHWXxqwJmBpwuz0oD/63ddpJOnQrYH+MkPZGteKIzwz8Q01AkbcjKP0aYDfa9fkwI3iLl
t/BIjptrLQjTMnlBOJnfHcu0SAo9K1KNW1rT0zmGmtvXoWFlM0RYpXUlspPmedbR7Y2ixnXsBxGf
fQcFoour/t1q5jlDZns9Tx1LuZfT98AdAJjMsPWS81WJvchNfT5kUP20J0y+2H4vM0Y9NxQX9LEh
ysR9ZkoH0jC8NLQTB4ZZO08ht17ACPb/GggH5/vynZtag0YFyUtiKmKL/QkGkJN1B+CCwgpaIyEE
Cg5dsHVVRnUZftNqn3+Bq/q7In+035FDD07645FGcmVMbx4J+wm0jcy07HN9g7P6O/hKA/yn6G9D
9xahNanIONJuKrGeb7Qp9bGlOLwifeEChCUh9MxaUg6EZFSapCTUcF5q8Ib5++9OUCFNvEhzZ+VA
DUvvdp2H3HUazAuHlA6sCtZG9A2puwRh5zWQ6PXudlAk60qD1yeCpWdbTbVoFW64QhqmN5mzfkQ1
xbuTPlC/xSjpc7HhrZqer8CXi4emsg+Zmu1KYAy5c02jxCwtt0HJjQrQRwmPbQ5tEK14j+qJUSFD
spoa//NKSuVTWnB1ff4RyAMBgy4/qBMUmaTfihZmMXBHWmZf0xTAZxyR/qsaQnUYrzoQrF0CdeX8
15SxU5ExTTsDfJt3jv0csEQZIdZb5wwyhzLIcNy4PuXnHou+j0yyvhvatGZ2NzzJZ68sKAzwwN2g
jQSgauOxUvm1ICKd4Uyjy6A8dnKyqrsTBipZVac/f8SqRNkuDvll2/QnWgTLGoQ6taqWvU+fy4hg
Hd9AOmcW4ar7tKuBJ23/AOkdeRsQ6RvuFNCKNf6nBT05JLUM4qDbqxs1ZLtUWajLwrrwEprnYHdh
A8+ztzJeN9R8ugjvtVLFz1hSQdogfyCVSReGE7QbhzjDwiyXKpUJZT/kaXm55lWJbkOnwXUOzaSe
Kux/JEOAhcTSyMJf4OwNlApYNRmded7snBrwOx/F9+nWzStClRCqJFa66n/2fk2y78SX1wVTRgGp
Gc7R66ehqdzYlNoe2wrFBNv//J1fCwJuI52b/tXUg2HIbgAd7VzTJUzLEnsj/uiG8OfmXOyLrfM2
oxIxnyheXVP7eOVmoYwsaGVZOQB3K6yHHL2L+9UwfEalhiNod0wH+SrZyYaXKZ7oH/TJ0UGJ1qT0
CIh8wA32E9w1EHnQX8NhkL8yGd2vvCLafGh2oLFkA3X3K6QjMKp3NRQ42PxEo8/gH8KNLOS7xcu7
UwuSxECaFXdhMAPq75ZGYx7tpsn97RaNpLz5GZRS1dCmNmwrB20z9jMOavPj3sO9jmPJlTLGfp3x
lC3RmpZ4NQBRYqSKb37ezR9x9aWZJX3NSIvLn2RzPGpIjtIAq+BVzSqcjEeMlim0Fg/LOjAojH4M
dWIgRGmMApQscTO0F+YbrfVgzZNmkpjCRbyjWPHf7zh06nwa6oG6SnD0xlGk43ww043FsUouAfwy
jeIm+oNiT1Xj7LWbyZHBj3CnmSd6dpiUlrdn/0c663d4AvECIjoinEXpmO/7HKiwz76nRQgoO4Nc
eWgBNqZKGcG2X5qQFKJVXKBD+UVug+/IqKIaUV4Z5vSTYyvuqkkfoJ45PA9ExMG0wQPmiQpTX8KM
Omsmh71ab/+JB2QpkTbIza1uIrrc8AOhQAJOd1UyTgy9f1ebLxXoDu2PF+PCsYCVqWjI8fdtsGoj
wie2JMIwez8KBCNqhnOZOxBeHbLxb5zKr5Ndz8G7TCOfKk6u3MUGhGACI6lUoa9fUpUAZHMWq7eI
H7o+k4Yw07XS73F8lOjo9zMBLqXif1ano35X1v2xNVytFOOKrJRJzpLYcmWfmJT3a1w4O4GAIPW5
ZcWW25RUS4La1uFSF2VmVDNkIsofKviSDOzin15MtFG9EmlH/SZRYS9wtyjXcLQJoZrFL7VFKrf7
8DfjsO7PNG+LCjfnxDzZAUNEp14C8cJJidovbzwDUIPiX+iqEAI4ADLEvfOB/UKyxx3Z7zGFySwF
hzuau81px3tufB4nlrnYqbduuiod5yiciXGn5W0xSAgsmKR6b8W+LVgTXXr2mzUqnzJ3Wap3+tSP
ZEhQ+kFNBj1ZaRkhXas8B4Ri7P09BNxh9v8AabUyDR6GcF8Qhh0EZH6E/mE8AE42gKxwJbrOShyd
joJe16iG3/mQOVBLAz6eeC4VN1rJGsJOQOl+5pUg8spD9f4RIypgXXSruqVVSRAjj2WE7DYzp6s4
RudSqCrbaPhBOhpO8bpCboncSB/iOKzZDEAb8W0lW98779oVDchRSexkc3HdJbme20xPn60CI3mK
G2KU4fug3PO3MoMujr4YWijGehn7bCxsUq8SkybEQIBC7zHMeUQmak+h8EYGZSf+fzP01Kc0Hn+N
62xW1R8G1dSQVU2NYXBJzRkWykrjuZKWa+nlwAbMfAxiGHU95Zy1xDFJjrizymifz7LArEcYq2Bc
M01zJ15XAmHp+S9DQmNS8ybYLOMDz++sFze3Mq9SNw2cid05BAFXRk/p0h2615kNhlgXdJN5Q/tX
6o2LvZgbEvwkxsu8ID8P9+OfSNhEooQenqM51LnnOs8kt2b77noAOkaPE5FOc1G+7ohKmD0+n8AR
2tXMMRixV/08KWdIETAmih2ys5eLv9w5xUAbLP3Db2821W+x9dHrAV/YPfRgFfxD+1lY26rCJvl2
JMCGggSOxxwy6Tg42qB/BG9YVE7PWzgmdOmEmaBVU9sBZYpisWBa724GMmIEom3i7KbzH/mM9s5G
bP4j5QnIgiHV0+ReDxTB1NnEXlOhhenQfo4xL8WXpmYxkMX4Cdkxx/vwL6UI+LPmzCkPj8XBTO2A
aAUh12BGIN79l4fUcngZL5nVVcTsu53FURRD2CZ39Wft+1DgnLMjRd/T+hk/S+e1WV/4pqhMGJd9
W+l7DcfQhJO766BEYxj3lzPTc2gVXINDXUrCPLB2/d/adTykOI9Sc9SuuG2Tcj9CzueAIhfZTfo2
DUbkhUN611hTiuxOUfVRJyr+q7QKeB2wgR0IirHe0hLckABL96Ut4yA2H/jdVmd5AL6G0J/BVNCK
hQWdBgCmHJ/m6WdvAwYLHBkw0wDP/7lsDxhRiiaRWQWcuBaXoja5GuU66OKNC1P5gfd4nTYlxdV6
MvZ2X1jfJXwtco5sRJXrX7bko0PO60Rse1+eToIDrA3HivpFzWJJNx4yDa0MMD4tNMFiGca2vm9b
v6AfOoBKGBsh7gZY+q2nivBapZNCc0RtaW0QPbkUwXJG9UsQmMDrs4nhn87TYpbaRdzDdjTKzoDN
ob6K/kviZ4wPhpif8iwHOdGke1HdnB+W5ezFXUajmeSd1ETrN3YaWlRyh3AeNZLykPO9zuuaSIp2
j4vz1KWndZlsM62LGRIT9F3f8+/qWzSfXZ9zvbzpAl5j22Oc20FkxdcjCyDY70+hBKSuuSaDBlUC
jUj5UXw4A8y5e7kbXBGkWcC5m9n/PwVpNE2SB3iYo/dlSL0Phw2Bh8keQ93C0A4Y8epOlqNWFXmg
y40V0TUln7Yrz1iCedt2UtyDeshHvxcRlTzQ04iu2EsRsD2adJerBWLVFBDQG+SdoPyeAh+1VuiK
RQB9VjQ0nsoRPGWgJbZnnOz1wrhYBLwK23UEij/4+OZB+QrjF7EJxxbCdTidZca3CFWjeb7w1qcj
0Ih94uankmeGTr0WuSezIEsbqpnsBxkje5KbH7NLVGVLGUqDIEU9Li81ZJPL29n/Tt5NT3rrnIy0
J7vvIVRCxBAREbMBk5BvlLeljkKYqOtS0UZTC0E/5kacGZ3od+PBhI+HoQ60dHbIrx5OqV+8Shye
nH4hlkAN3su58yNTSvk3flV2VLl+GBfUlNIh8x2VJMBn1Q/vDzmMhoBq+LxCshgGdU3cksvbu/mS
3V2oYbMevM4fEIVB0f7hpM7NdSsLuJIUYR8fsTuQEnC/8Kx+Ehcrvyh06w743qbNIj49heSUIVUn
poKtRXirFl4mO7tIZeBxmFipFJ4TQVx/qoG+/4rL4KhwL7/bBFHL1sGpIgqgBsdcdXAZRSMj/QOo
eBERTPBC0Gnx9aKBrphe3UiQ6Jk3jG/xRQVFsLlBeAKrgqABEHy+BVnJdS+CZpPW77hGfCIhIk4r
06bBn1s9REP9UMkNOh7jMCmZAZU4aPXjmXlXvrS2Ngh9Ju6xNaPMOZn9miT69GNjJnsg+GX7Evi3
vt1/2JY9v4Cq5KuGQh19enxbwZ/jsq0UFA5XMmTDrLG4GruXm3zjj+skjwehvYcz7XMlv+7FhYBf
uFuylGxTdEGaNTQJOezpcAyWs6EnJ8FyoKDRVECws/c2kJufOiwCb8X/0fiEl04MPnJVl+KUB65D
7RYBdhnnuuraViU14sANkVLr7Oqjrzk99wKZzNu/bgp57yhk+DGs/GOgSlCoyBUFXRpRbM8ODAfo
xXVLFP8639rK3eJWgDvk41trZwXG6XR8T9SNjB6nnAGZuqA0Wsb+iiZlgRj0NLt8PSKeRtkKci4P
S2TgCgYs5tOVjOfJ4VJLpD7YWBjq13BRlrryW9nVrc6C/1TU8SzP7P6BNOa6v/lPT4N7il1XNrff
GleUCIe2L1Nfkqu3QotnSi4fyFpa1QnDTICY7n6bjN+iYsSYH5HF7LzpON9bsshFujTOP3W3t4SK
qxePV8KE/5/vil4iOldUAGnANj9G+uevwSLqsrYE6p34weAyUroSxhaIDv5Vhhg/vBPTJrkG0Kpp
2MQBYhjFXFXDbSB/3XHZYJ5B3OgFKLLDeCccnqlGNBo5bqfAo91rHjs6jc9aT3ihW+5lMrKttrEe
sgwh2raEUhkHwbqHxDylCI6JLmNCqDcIb3nME3oqNU6+dt+xBwe9DcWznjPGVZ0EHSQnwFZswnNW
wq2fIxDIFpm5vfensGFaidRrxK+2RUt8pEjczCaikNJSiYKpLJQSvNQyxBSTVkSoYQ5nWMY13T7M
lJwd4FMupiZjNVU9Uz7RjeXGiRLlKdBH5avRkXv0Nx93jnT/mgmy9RqapMJUI9WKCzZzhhIjoDrf
vdjVRlthK8El5Ntf3Q+6TqF0dnLV3Q0jPw9tPPwjE3UuusAjEt/8CytiMoeD2wlPou8qSQ8R4cTk
8+OmUx/Vzy+5Y9tUvhtAAKUBYZ5AfjVzH3loAckk6nL/bcr56bTYZKAOsno8GpKbiB/CURP0FYuE
nP3sLkHOH1FMgiRRfozdiU9pZpD8nII/pcKXdLUzF5gxk/1jsYncGjCE4oosyjUCLKLHjj214rnZ
Qb8IgO+sKEiNPLxtIyZ4SSeYzTlC36ARnkHFyuz4kARBGC4aOAn9ctax44UzaqOvmR/N00kYTfjC
IPcyx+mE3+2+EYU7Gi+gW2fahk+5xs3bC/XXIv5p4uHkPvC6cjeXSJASIRiXi+LSJ3cQRUMZm7uF
wpNU/mWIAGdbJczCud8me4JgXAKhSwUgs1WLBrxurIZJ8oHhWt6g2hVcT18AQdkj+26p7xmyTOLH
ymbAjurM3wv5ZCIA+Z11jAuxZdXh03s4tSoJVnnODKyY1VpRau93YoXj+fKFdaOjxEI/13sqphIG
1snfYuNEut0197/WUDhGtW5DueAMBA0KoX4f/sJOOTus93sWCZVUhQ0iYS2JXPSM1jMESBe2bmRn
uC3WToLryZwL7P63XGOxyrL75eAhaipqC3JrDBYTMNqGpuPAeCsaBn4S5cE0oI47g5kw3Ob+vIPH
koGjwelBKfG4CXyzQqMKwCv4qi9uZGFBNm47bEjYLZvZ0CDSL86IcvzYH7GFi4AckxWSKZaZxdhD
ZZ3SkATAJmyhQDBlI1A8gDnQVFvmVcDU8XDjgN9cwwFumlvenKm72wWuYPU+X2a2oIngjWBPVdHP
GmOPND7gcL1rA7IG6B+/e0sepZDin1/4lUzLLvp0Whxu2LdAX45s3+eD4A5iKDDXdY7YW3bImwDR
k9tFNU3K+IBAdAfC+vbyi/3LIWarlpX9XGZy6IPrlw2YEuYW2j3Z5O5RzbupULyFRK6ntv8Pluzm
CYLMEGFAG0D5pHDKAUKGdRUYj1u2b17eMLqmf4UBOVwY8HKqn2F7Z8huFAk/NJlYNodxFJhjqG75
UoSFJWL24oG/lZLE6ReIOvZMZDPOe7QOyp/cNeuURVrk/p2yNLLtxEvwoPZuLj8fsRsqEEdvb5cn
MxMIbtYwTeIP32qifJhUrW4AQD5+GP8OC9LSJuUXxuuRpsdwpfLUafweNSIB3Wch5gCaLtU7CxDy
z6/ivdYXKTrfUdBt+JmpraiBsAuyx/FLKFsAYZTWjM06txDj4qrKrowmW7Tsqr07WlXNswX2qCYb
Aa+4GHT2WvqW3d3ImfaDnVGAehWOxPochZpLCy9G+0BWyWQf3CYUcEnfSLeE2HWHnYcsfvDrwclW
KTLb0WmtbOqHvUPPj9/ycAhS0+803EQUL8dOmhKHY3UNHkyguKFA4SEck3KyNz0vNpnPVseCENyl
pXSiR/Q6vANxcL3/W/DweAlX1lTbC+keMUgRFDHFuaECuZpjNCe9S49kBENdY74HVAh3RkMDvwfZ
CktQjBBcuiUk2GiXzq1zx6dRIonsLqv5s4Ag+0BRURbpIrxMGxkEETjxAMz6ZWjX4zw46AfiZtYQ
yAEJwgvdhmsUpqZP07mMs56dVi84pBG4ZB9J4pnvNH9VVyY+7O9yW/r9Oo7NG4k8pdgrowcAu6/r
nVUdHVfSUL0HRSG6GmMWvTaCwgGdTgQY809S5wJem4yjuZGGg+wM1XmJ5HUy69NkMKmd2heyGjjP
wZ2ccEtT2i0eFlqR75ODh//DkVini/XqBtkes0J+BZ02JrM9NtZ2Vlmnc0ershT252pS0ysqR99o
PDLp5/FtEaTfmODKIt0DQtzU9WNEhzwf2v3JUxYUzeW86x0viLXCgCxTvCjJMnHrrkr8h/fdEMWg
Xjlpqp9zCx7dWmSTVYzkpKu4zNP+9puD6z/z8hG3yynglmaqJ9u8vHy0IaR89r/B6v/vSA+kYVoq
vexk5HfRFVNvI/kldYFc3Cl1hMqUwxsWNBthC30jBDxM8pt68GNueiN31ZzcCKr0dAx1fauLiXtY
bH0A92nBnfCMBXkCUcKJvxiyyFDYiExTYSebzuDnLw50k+T7nD9IONJ+V0BSMEF31rPq16Qvb6cg
j4Hgyo/e9Bx0ikAXm+1XvN700wk6RqXMW4izf9jNVn5aOJ1/RORlGVQwnE/tyx3USY/dUvFgNnnu
a/uBTdvuZ47V1XjKbQMbznvZN5BvP2hN5ADNNYnlIAGY+mYcDBaRx/x8vbehjzu2xLSMICcuUknM
3gbcGnmlExpEp6S/BDy/1JmwoQJOUNbr5AZ4rkRf4Jp46jbgy20prMrYdeiH/QP4eVuylpqujTpg
slhKIGj9Xa2yvYG66SRyyu5nDxcs28YjAnqYi68MlGVg9WGw0grjFV761V+T1WKKAVEhQngYK9NS
c8Q0v1zA03Gvbp0UgdjhLKJnCIWnR5e+5is2Q1PpnFjGzo8OMbUttNjqe42rEMDi5tWw1bnB4u9E
KEa9cruVnnfAtpbev0FNPaIaW8MozzzbOBOacQrlSXI7h0A64y2a2ybt04m3NPSLONcjj+gbqLxz
g727jaDQPIxiGmR+W/9F1ypdQ9aEiXlARecQjeTviBMxvw8YFi2CPfqJ9EKhlfAzaSHMdTXJvCCz
ZzKT/Ac54gOV0Vv3T9cJ56PwpzBC9Ld5Thla0xyyQ/B5doMYun5gdoJbAv/NGU2BDudNkneQ07Hu
ZIqu7emUdbsmHLaG/ebpcL8BnoZ5mu2+RWegLh2iAN/ugh9iOBeNpiiYHqg/vzHj0A0jBcH1yqv5
kRu5oDzp9nGoNqjTrwAJkdFKMGl7kaAPs5hmX9j47TrBPtqnH4r5LH6MmbZEpxU0hMIWiAqmB1C6
zxp3q+c4OW0zqz/rGZ1Cgl72GyEE+7O8swTaRXdrl5qMJGu/ywO+7avZLJMPJeRD9AiQII2iV+e3
+I1r2p+AuZoe4qPNvdniHzMvahvXvxPTbDiFRAb9Hrm/ZO4cKZx2viYx2yqTCvhooHnblE9KvUqC
sCNkucl0HZI1+U10bsEyZX2HmTTnJupC51vaK40koXN/63sd7YQc4g8t6U7w23Cmibfi5ASmP6sP
w+Hh4RRJEdTZWTINkN0vW4wrsWbxMqsMaq04jMXAOIkJMovRsdn8OghBFguBKV9px28BIlLOPU+p
+gkQFt9wq4oCqu1pHbxgossYMSQaCu5Q8RX1Y8seZo7QeggsKxlCfkZ5cr7zufwKFTdSEWE2w9XP
Gf+QTiJdX/G8MJrxY2M1Ph7OFQbcRC1LW0Gme0jthqK9rYupNcliZ7R3bgzZLgtQijFPaRrEszum
66/wofEHm0+HU4c9/DkELDTjSJNa8QkrBtIf5sKrgmZTqsm7oWqOLbWNpZIZIxcptvdOUdd5B7Om
pdQbMmamkcNW/Efg8OFjJ07xmyJtAd36YB+EItuaSodgsBDXfXUqET+eexhT3GsGwEiJu8Jx5PC5
RQNZJyk+qNAQwIGXZ9TPbKA1bQ9WpuQyAKagCj4NFp+70AaJFO0XeVchodhxdDwbgUpo7w82BZCF
5h8E9+TxhBNmRXqFzqjAFgr+jJWNP7vv40yNLtCmb8ik13tDi6ciD65MCuaeY/DHPM1n23vXzyqd
04Vdam1Sfru9rzroVGAntxQJ3g6DURl2dhB0BRiUVVFilt3DCpzwH0UCKeiOSQQ8RglxLazyd55P
pKcxMjc0wZ/cycXQv4FTYaYcUkepZ8Md37v/eKb9+He4a1Ghl5j6QEyQLO7icT40Khefzky7qoqh
7Ezo9wzIUq3xomuLfGk4GvbiZEbt6J8ot6jMGuoq+8rVwdQdPLwPcgM2h7ctPl41kls+Md5Zl7fU
tPIGELKvP/DbCkPaPMRvaZysnT6on/XhCnGPX1wiw7ad5sE8C7HSlL3i9o6hR7fZjeM/YDjkJESK
Qm4z/8RuPDpBLrfpVQVCGULNgjOKaI8lREPdbg9s1WLGcKEbawt4f/2IYZ2FC2Y3MjPrjOKEEwjc
J9SQb9l++llzEUVwZACKby54Nv2SrLuqpkynDJIn+c/V3T36GvISfiVOBlt+peP0Dhos+1BPcrjU
QxZeYgR4nXR0Fh4g+M2FzG3N0GG1Ky62ruo0KKCUfUF58zHWlnFt9gakU2PpCWMFcEXxisQE1YUT
tbY3Ubd6p7eP7cPlZg2LB/vDQjQwGEYlfBIVKleLaNa0KUX2gQvWTUbVeMo2ZJwwM4435VeqDSn5
y8M9a9zMB2tEh2K95Jt1zKY+gAy4VgdQjaBVLpWKBtvA5dGZpFNw6PXMYfvjn33Jtk+xSTzVu1Ym
V0NUrFZvzToPcXr95ip/joYlYaBIjLPwRnp4hks47LlS9Ix6hO6kBq7E/eRs4WkBetKSzLY+DNBt
tSOIXbpOmtYntBHft3pHyVoSXiGB0dq9PIJE+JRjStOA/afzKNSYgUHhserOrrr6VTXP104LVp3E
8Eb9DxWYeR1/bN29I5Mldc0ips4hK4aHkNq4HUUS/QHtxN0lV7QGGGSwp3rfx+P3QO07s0r80c2u
5mu5lO/OotkJlCDoBtxCfavLpjH+3KrZeCM/BuAII4EJFwM94KQM/RwUgDYiiUduyQknl1L7GBtc
zpK+FhuWeF2aCvaHbSbqf45m+4/J5/ZaNfIL9M9ZJ7IJsOs3m2dJCDOVtppCbYOa2fKg20nRFcpC
AEcsVRCdvOy95rMeNYeTpmrJU5Y03Gn1s+Hk+lZGpCbtgESCJpGEJekrA+Od1385ZBfqdVWPVrfC
BT+RYbf+lD/NfGrHT23Ik/uTxmMoI2SdgP3im96bdTK7OAg9ZWQxs30ht90qNb0xkJOezY/3fvtJ
TlB6EOxGVkgQ9TXGK/uly58NYnS7Qes1a4ZGXUk+49AuXbrRCIxakx3yMR/EA8oQJJ4lb//U8vXD
P2x26nBxYD25ckHRdT0z10Yt9lS7w1LO6ruJ9DFmhcl7sqkLxM53GWBxTDOp6+hj3Wb/clYjUz+i
83GhIT9Hcr8R8Fv/lPC4rpB79fZ2HR2S7eOWATC+37FF/e2UjXmzxvwm5cJwgLzSSujKaTcIXI/t
c8HvByHHN+jNKE9nKF1UeprqgYobItkXd5D2mdMzBgwcrI5U6Fl5ZOyt/emX1trMS8sHo3qd+nnI
jv5uwH5udo36Nc3RMA1ve2Q+XpOwnUAKzDp5aJv7o5Oju7uzbzeqzw9OZz7GpSMoHNViOwNUh/Gr
XnofEAP4HBjqRrgERrlaaEjvEFeNi9q0PupOOkGyp7bJrsyedaA47Ue03+3V9eAyvllLXyq4QxM8
B63A/pWwEh5cFoIfctzp4pAdggm93lWywhuojyxbb1ur1n8RdQLeNDuPQRazNrsYMJ+QizYFs8E9
tSieHdTfWSyzmYFl3I0ma8MtAwLv6X2+Zg9izRIJXsrfhgHQyY5noK2GVfFlyWc8q9S7kOKKq8rQ
xDFi0ccyjOaQmswKvDpcEi7QPYgslufK3jg3PnA+BS8ypOV3VGEXU7A5keGrCJEtLvIhCO/iGlOj
Xt8kktDYuMctRrHIV4rtDgpL5OLXAVsuZcHC90dirmnFn2PAHGx14lH0C13KbtCv/fQUSU4mlexy
4taW3EKmGeTYGtBp/XVgW9I83uTRzzpAbHw1XOZAOTR3gW/FGpqO/A/l8m2Z5B8/NVkAKkr8nQaG
hnn8K8LmIGihRxoPMHWnnkiz11H/twn6kSLTJfmunxP4FBe4+Dnf4Q923iIllC8gxTUghNay/FqQ
hv4Zmhr2LKGGXrYJv0OvOgEndtRxwYslMzkdIjAqEkn1oARqvE5igWhQEWVYCKIv4ZROcpj1vIxQ
iInuOHwQHHlWRAmFB/136a3roU781y+s2RjvebJpJ0gEk85LDhM00CARIgDhfp5bfD3gzwdQy2Ae
BUKWF74RhXXgXsWzMiMmNYpANcIJRmyW/CsGW/Eo2b73lcA83LeXPTtfNNjGULXRKUJEXIXetYdu
TWZbRfbc3Z65UIkLRc0FzeNBaRlQccp7yMHcoWgvkVwRmEMNl81ZLp1yAMnsk4/22tYheej/hf1Y
KVJh/knJtVw5WFZA97LbdbepdPM7Ob+CkNgqtvGH9t8v/lskjVhhSCukAgXW7XaHdeASt3P99s2K
YT399zNKFZmrxOuWOcuhDiljZVjfgcmiuwOk3HNHDgyOt6Z8J6ZyErPMNhdUZWtWQ8EyZtKk5eYg
UikW4MGnBYW19WrEPEGcuF1x+YWIXgBx+qOPdxyepPh+bXYcWyEzNPHFKIYrykg27H6X/Q1Wsny9
pifDNxFcZkSeOx6BOhhUL+NV6O1wTHi/sbEIwwmXzLZXWeWLewEtMHXuOJMQ3W6wdTnrLEpMcCm1
dyFNkDmHz3xP51XF2E9vC8/AGDHdBmF/VUR8AZlCKOWV3H6HhJShj0etf7ypkzkipJvSyzjSvdy5
n/OfXayH6EYZ1qkyEul/ckx4gVDWycJxKkC0YjEvuHoDBNxUIuoo7k4WgtfOkl80236WDT0tT4Zx
Jf1rS8zUmXSwSTSDSpq52jaMZiWkdPZRe07OWsDOkZTohbSSBMhiP9hCCcgBslzQ/mvViqDVyJ4c
MZzTph6J90VJsT2vRtYP7+moozMyj1jcsd4Roz9f8jrovlsL7FH7Ii4US/Il/8DgOmTMtjMAS8x0
YZdJpVxo8/OWXIU2pNYHbiK7cebDzT9eX7V5hFWByOkGSC3n3Gp5KbE/DJR+dImMhl6PbCJFBnSs
W98J9Ma+jA0LNl7QXDPv8WxZd2RbxLwxAGhaDHJ4Xq8tHfY31irvho5jW8rCFkjN3Yepxped1xMd
15Ct0mAR6iUJm1wCfYLJiIw4Te10Bgm1jCm6gezTo+GF9/5feIY/PCgaRbTWQFuLxU3B0Gdt/tZd
xQmU0nzvBL1qgsxff0uSMnU5n9g4aIw6ykaLw6SMhqJ5yu0AVTYhJ/eCdzQJjLD87Fxv0FJ4TSdz
XW0nIUvqBAzkNe+z2rlTeDFNgCmTdDvsV2BK/SKCQW7M7EGP4xUmO3m6MWWWXLN8iKUZQB/abtqr
lNU2v3gxXizLOs7VDXW5lZilTi5+edJpAqcAaJNkTKQ+sDBc8w+iW3sGc+6DD+X4hHbIqJzLiybg
IfgSEtzPwewyZqrctS9vr66rJrkNRpknwPld5yWtV/CaWqoRN1fVpk+G69xxbfgnZ/nwcIFnvP+L
WrTkgGlmP04JTDaTvqIr7NlyTnu3b3sAh+fnnFRrlM3jcu4SzC8CuriuQVEiOcjeeEs3Y3jGh7t6
rMex47NPgfaORnWXNSlWkdCfQgn2EiduvoQTTEXF3LPPjhqGO40bGNGHoBuWpk1SbjmAvK4C9DM5
tfEHfS7xdqXp8E96tdfgmETFEFI0Jd3w4d6pucE+0pSXiQOhWdNaIYxNZWVR+sPE5wdLzwMpU8GE
TLw0vkjfoQuurGSJYPY0FPaYbnJyh7zI9wrlurIjka0+Fr2dCWvwAaBuaCegNqu/Rd4WVv8qzLdW
EQxO9aYI1rYNIgClfiLqmI0OrOVg4h4OE7kkH00Z7HIGTOp/acnNhR9pKlt4WPiMDVKHaEBq+rHe
rMXaqru9VEqX9hyVuvJZ2jyRcvzmtJwnvC1FKbudohrBPBfzl4QsruVTJjBVqZEJeUkO2COwcWSA
xg/a5cu8KKKKkUxFEvwQvzBfm9JNjotgph4aN8Nl8RR6dlSCYxCZc9Za0ZeofsYDImft8WukuWnc
ClYQKNq+ZzQPqDBy5PnWb/iyQuvyHFHz+od8vT7ZoxA2s5a3WGElSDfT3uc2JL76rBsR6UUehc4c
U3XXrV/cWLJaFVjCsd4r1IljuYueORfw3bThfNnAfmiu3u8yxrLeyjKMEyXi/LQCOzC6ckoPXwd8
gL3BtwL/QP61pLNRSzNi51b85WjQb2qYIJxl9sWZN9urTZ7JC3pDVd7M77jc7C3JKF/N1w6ooi04
VAPGw8/9osVMeCVUK/gBey7YMrWHkYzqiPuXpzd5PvkJhCgQ04Gt6H5XXCQIXUW8IKEP1RnWfhnq
wEJtkOsWY3MzCOnGTyUOf8Ok99mXegDLljgbkuDEL4IuFY7SFcia4hP0OM33WI/TmIUKDmxBWpB9
9V0SX2Kf/FjGZra82jUhoodVGb40o9E4hjH46OS2H/guFG9eHTeX3QJnpDfQAaBvCIQlTMdWNKsk
056/UV0st4VxA0b6IN0XJSYYKUHIaXIbWafURoyRL55MxJSzwsq7tRR1KrMNFXcca/8oKkmUClpy
Ippbk5WuHAjpCdGP4w1h9W3TEmYQ0UGs4/LqYRYs5GX8XL+fO3EItKoBKTc9jKBjzkBf/2oVquB/
G2/yXAZFWluW5g43oZWIRgZETWxu1hPPjtCa83WxzdpaIdDsbfQGSLLVK6nxdmg7FiBJ4lZj1KN9
9QwHenZlEk8W1yK9cN+k5vZMhVIr/JgUnBwBzoG3PrrtgStFYXdFqU2ytkKPL7vR6MY99nEcVPv8
749w58VELitlAMRreYfMnrSTqpw9K2bc5JdrGQqEllf4BIQ+tJUltk47N77yzXUjDh7rntglNagf
KUe0gNusxJRrMRH+6/5EmVUDETd68kaLyr25PkcdNFyinBbkfKKmmC9fw7CyYxJ01sU4ggS0OpOY
phxNmUTRhGie9aCjuxoQzN33iKro+XbATW4jeA8kww0nSzH+1xjMexWtKFr9SHGmrBqYnwzgxIih
n/EvtiLkPvZi9lPK+zmYDFRDObseyt1PG4QZvOaIIkK09+RNi5ZvOwc6lHwJLutF6ag9/o5JXB1X
GOgfM0cxUU6liIb5BTzQPpl0rULif1T98VnC2typqIufoUS44i2TC69uHBG0/mYOUvH0dhrj/+Wq
hTKskNgbNCyCPOyUdkeny6z7FBMQPJWOHslC12SsJaogefww5DSr4V9BX4tPtcuFDB+psYJ0K4sQ
RKeI5prgLZXGzezQwYksSTBCQRwR/sDTnkubwi1A5IPhWPMmSWq5HLcY344bpChmBvGLcBcLGhj9
sbmO0mdznHxEvRAoC84fRg2igMMPCGLS8k21YEUs1n31vhpGK5OVoMV1ZRVeD32igcauSClfQ4iC
XoHKJnIBhqsEvrmWUe71Jt8ysi9zrrsdHTkez8J/iT+r03jU9NOXzi9YWT3RVPFlU7bP1l8KzJ4o
RM3yIqHcT3G0MG2V8OE+PzgLf6nZEZzYGNFZ28QlYevaKJdRsH7+QuIY/KzmdO7BtNLLGwGpHJ2t
Shhj4wXgPX85O29qA9MsWdofcVKXtQgJ6umhmOz3IxQ7jfHEfi3+WMbTesPXRJqOkzfg+fmTdmLv
rJ5rIfJjYHlc858gowigtGELYbc2snQAT+almkwtV2riAka4TCdKE4AGVOol3dw3E/xrDtZl81Ds
Hhg3yt5JU3rSNwoj/lBXeM92N4wtTdykZIAln70yxW5hf7cEtmoYyVo1G983hOhHlLfQqk2hFbuf
PF+vUJiN1ykd3aQFgh5UXxba0nADoHpOpTwys/rykWO989liVaTqnl9wIGfmQson2vk3WcXGoWkn
rW5cdTIWXaMe4xziyf9b9MIKEyeR+v6XI/Lm9Ynxlm62Ju7d00zEkin3W+rydxX3/GOw0iElwSaf
ZH7/G5Lf5SGq6E8wJBu9/CUKtBrbQKNMj7rIX6rfQv3QsLfhtH2wf+F3x6xxcoqqJ8jeDCMxR8dS
4CpeCwsLHezp3MOuEVu8gMoSZ/rfBtM5wtZ/IKL71mgyRMqJq8qxZ8eIUgZGmPF4yD8PwyunBjWl
jMNoP0gKoMQvDINCkkQqJZH1YjwJYvoVmRlLpZFh5DBSGp47/t9WIAj2ppl7XOgPSg3C6Nv22Vix
MaIuMdGEWbTBwR2pGYEc+ZYD6kD+2bdH/FSKvgjVhPFBvGa8efflKNf4+DcYkn2HnI8hdpMUc53x
4+HglzVqisxiDWQ8h1A7HP8ApSYSrXTaMXK3Ws9st/PD1wxXf3wJPQTIIAVq4E2JNeIpTJFjMV7P
D63icaetVjcuaXOW/1xXTZmJPJahAzJWP1S9b1jqw4H4+dsbxz1sEQdpnnf2rPqDyJMBnmSnhgeE
m97xFqKeMpmRBe+oqieXc0aIZmgbCg4GLHewF/RO3KNQkgHDKrIzv2Y7PXQ3Ovs/E11HElU8EJNT
4W7oNKiYSPWj6YfDgvH6FamspT7Usm9X74Ze3o2y/ddohSNkWpujc4XZMmRMfP0PYX1sVADuk2SN
Pwd7o3zXothU3UIOSj6HUuZXt7ADuMPSims4c6vaIuZNBsgJr5nFIUXEWfetgPac5QzTNhbl77Yh
39ytgws5VJ8KyUmIISTbG8wDyx9fGPnzHYzmqYbz3GihqZcvJJXTvSzG/YSTVlCJ9lwEr2q+0F14
tB7kftyHxybdg+k0cGNyOOugvSCUBSj2LVtgQOoUQ6+NXulZLsqyotpmqJomGVomvXpOeoF6PX1I
7ZZHfv4iy4HDvZGQV3yC2Ug6g9m5oWJNqh4Ki/+ZLOpTAR9sUAFNoizVrNz1gVp+HmFdX4XQ6wuS
fAEzf6t5cgLuFexKqaCWjWJazJCmeONdJaI2BWuoNm4z4QNIkOOMIRqAej3QIdXKLvixYaeZmmM1
4MgQGBjmxZkHnebYTNqnjnRisIxgINNU52youXluVGBwkYmne9W5caX77LNCucnCyqhViCc9qLQ0
Ngix64qWlGya5M58cZikTkq0/rt58/5MFFREUuoWcf2HrQJyJHV24+hiobchCUWAJ7veTghI7Kgt
e6dPKp8HC6gK24e6hqgvVhDcVPFskpr56Z0WIdxtG6yZnydjoE8ZRQPS4tv0tfncWo66b9zjFN7G
uq825eLtnSKZKDzmiGKnqQcTMumn2gF/Drmm+7WQcr9QMQb/spRMwfzDFt0wwnxpLmpTT6m+vHgZ
U7MEFWyqTHJ7g+RH8vcQtEfY6x5qAzpX/LdEhkwBq6OyoEOw2yetLgkn+NWJ0PkpqnKcVZelRAJd
bRfg00YzNeQ0ggdUUlrnrFySJsp6IYqsrASRr32JJUpAxproVGx6IGVBcoh3I20kTc6J6Ci3o1JU
aihQgjIDc+MNM/sV92M3oVllfC7DRf0FtMo5e4PC89QXmNGxbdv8tYdxAw+u7KdoLVrcDEsZokZU
E8Lghyg7bH4j6ZqIMLnN9oi9i4xk48eMh2F7YKQURA8ZxnRoEPnlTU7hXfoGSORwEpmdVp+2zFre
AwHDMUm8UqcxU8fKHtrPJ8rwJ1gpSy4Au/JR62Y8mC73OJAh7eVO+uDfo6h8s/U5rCf/NqIWBvx/
QuqctLiS6tOGInBdm4Qmzu5Al3ttHiDYfGXVdoRdwUjnLqyz5ov79GKYTQ1bXNhanuTcqjJo8byi
RKVPpkBtr7r3JCLWmc6Ms7GSqi/TfOpqOujpGfaNLLjZybTuIt/RyWhdfTMCY20OY+DQtpcOfCV8
EXRR6ohANf2Ns//ZnnBL1hrmHbS3aC2xUrZnmEjl8ZmjRwPC6MndzJY+tJbAFiTg36S82YlJ8SFa
66P+q0aokCY90IIROnRmFJq8RvrO1077m3oF5r8SaFCNDcAsh0mzUWSj/qI3ebBkVVjEiWBYsymO
RUXefmzfcdQLhNzIYmInth+TcHEQIFGHm8BQ3ymUuPJ4qQj3Fjlx37mREjhAKpaDKFYtT6WnH4rD
O/G19t5Bd83ocqwq4I/xkGJWyCeHgCO1o3akh3mPc66U52GSqVIh9gkdhtGChX67hR38MVd7+Y01
ed4sevxAyvmYXMIrYze85rX3mWxULkckXhc2N0adOYVtnlgNpVKUYF6Mp5UjeQG121OK0C2CaoqE
UDgBr/LlQMniLsxof70eBDCT6j7lgGqwfjS4XSEX5E8Otl7UoGmrshv2ZYwJS/1VXmWWNx7sbfJs
W29StmsXvhKWcefI8jsOmNACTqJaZ/cO1CtmY4/ZTVPsrkjh25XiabQYbFpchvSu4ErrtrMKbcVA
Cn5x8f+41pT7tx16eBFVYWMgdTdHqfIhANqx05Z8qy+ITKsrqP4ZEcX2E8YwFXeQo1+txF3OsIyn
t/HnVg0A1Pbs74ZVdNvKH4p3N8TWDZ4ydJqR4pzX6GAZOJnfP8rZobU5S4Qywud59RXWHxJzSk9F
ml9YpNTroXBPnBfLozaPZD4aXpG0gt0RqUvZVfbB1MN2Ur9YbG3nqGtB28J0/l3srhNKuKn7bE/k
s8CjQ+lj17cfMnugIY46n5KQPhMpHXh0G6qhrVv3r2MEkwODUBgslRk5//ZYz1Y9tWtS76+g9YJI
zy0q1LLngqKmVxaTVqzohywg57UlKDp93xlKJVVliLy85NQH8aExg2w/stZqP1mxtDCd9VdM/CLH
T1zVUGeKa2pShH4b0xUtJNQlvz9Vj4wtg3DfdEFgiRlD/jvp46tBtbcjqGApQ4R7hMgjWDjVqZ3f
7Uj86K2kVft+ftxMIgB11gIev2lIkDBr//BSZnqv4PJqOe9ZqgZIzJYvZsPQfQ4QeHMm4ydesMD5
rrvZ2zkhqICLZXIO4qY7Saz20DLZKRPaQrHlqdiO1W07muTY/hs+QzzS6WZ2tl2rE5JgzoCdk0Q2
ZGjVZjrpodfkGIhizs4Ei8AHgWkoDsWiRhCUzp7tFZmLapRaNhewVzKEKWZ4UaLxkc8knz/Y+nCN
06wlYAR+voxIIWLS2Y4lZfTRcWdYOZv0O7uNTfTpFJUnlkSjJOcSnUezw0jQovC8UTPRxx/UVURw
ETZIfl8JSGQfa8IY+FlbGvGLRG8Sb/pwaaoUxIVdnOaynKB1N5PXujGyHcKo4GeJ84k76dV14TYA
duotX1j1Cy4i4GXIB9nwVMmYRXGha8yWdexHQQr9nVaj0cTw3uStoDuHHBAjX7PUDXESEsaABHn9
FKsXC4/e+hHvFsyZ8GJo1GpLoI283XFHwULbNzUkWT4S5u/ZigztqF0ZfnzgNot6i1yr5ColsZqG
vc8kUOKH+eRVD39B06GFFpZDzLvw3Ci3XjpDXXBudxEVuEQkLaWNgBfadB2q3/lipc0yBLnUfELr
v4YjDwMQO779TpfcbDO3eMeGgQ0H+T8yVpLc7g6psCAL2zvqsYRxCtZBmWMW5foQ/XohNG57mVkg
p00enoOv77nKnsyMW8F9ZcpnhKo00J7JzGqhiUcn1a44LTFpFmXTUNVsfiTWsRTlEnJD3jZUW6+s
BDKcUbjev6U41uylKoo5NsxFJALOLPLfnCZCxcW7XKuiqYyb79ENxYZ2BgdbbC0sZs3LL18FLDL2
4kwqSu2Ag1XRPMZt3Z9Sk5fPWEwWDq0hUzZkLDlI3+CEIcvjrCEQ1LD5VDrlEorK7g/9F5Q+umnb
pp5ExjVAefurDUMzPoIC6CY9MtnT+glYDiJejmuLLoCUBLkm96Nxrv/5wIIdy6R3O7bHMhjPtTJc
HOfTeGEgyZdA1IKjnRbTL1R9u8KgVh24YupWQcmxiBGKgzbLO9Dq+KwE60gqlTVr/19o2jqM8Cjm
0Y37SjOcd2DEwlNOwBM22WUxskcIL02qykgqzkfMFr2VTbPBg6lPPd7usHIv4S+EZvRW8Qtw3nZT
MuGiV5J5diyVO5kdXHyKkMr/Nc2sb9Gs3LFNZ4r9+MeZD/hhOr/Hu7+WOuCQD9+mK4gYMb2bAtV9
9Qv/bzyje7N2v4jxtWNk/5ntMt5tNWVzFlb8lXXSjOlm45uKk/476OQmAu/77BkegVOk63zOu/W/
6ddbgcjLlvj1wziGv9R/yreQaAro1AKnEfB6bUV85ZdmIVyWgZzvldPEF9pzjqqCfLNT6A/lnx5B
l/jqTmzd+SlEXb2eO3quNV127EDSjuY2T1gmlj4nNMzFP4U9piqyEoOyukNb/amxOgfgUQf6NvFT
Gej+PJb7v4kRUJn82QamiSMVnljXvUF2rEUMYkY7ChCstr9DZG0rtL9nd+3R4VILGSqgvnSF42bn
yAZYk/E48G/k9BMsrVoIdnfGZcxbXMKSc18Z2jYfCv/teuWK6h0MFkLGpmDc/TOKxePXE2BCkozS
n+9JKY5md5eM2NyvUNzgaKdBt53QSoii3VVWLXEUJRejEnnNiuyp17q7aTHC93vF1dZFrOxoGDFj
Ja9fArMXIj7Cu5TUDdC3Qht+MMXC9/66+70dI+OycxrVz7NnVEmV6o5M+B8Br33a88zgPZV9nIli
LxF8j6altd/qWUyKT2S9sYqZwN09s7+jLPxDJExrq1gaXYHjFp+uqMlpvNCeIDdzIrIpLM4A2JLj
eM25iZus6ydHqVebDKr2h5VKXRBAyRa/BMOv8jAL0PYsgG6yoi9FNu5fl39s3FlZP+/427WTeVLf
eOUwWLYyyp0jvrdFDFxMd9q84qchRZx/ONWKTmJmoUGpzmpvZgCHzxRDHa2WExM3ws1Ixk9KKKiK
Rwg5N1btHid5JxH1UjtsMGwRarVU0DF4nQAsS01J58y8UDW65djUv62UEtIttfR6EwjsvZSsVOd7
OMp/45n9NHMLR+hk6kG9gNZZTqYlEYy/WGS/5Tv9R+kNyHkP3zpfxFsGDpOsHAwPoeKLNclyLKFq
0UU9d/p24JZ5ibTN9zyjqCW+i0HYmLSDgUh7dx6Np0QRhhYbkJpO5/pT+VOSDiUjH7L9B//a0lek
d94DiOPB/CgygIl46WY8tNIjET2zMz1KJ+Fe/g3Jp3wg7XpLD/K3gYbermM3Dcw5gVG/oULXeZ2i
i36Ihdn2Mox1YtWr8/3/3HmDw0ado6lBEK+HG2Y0FkPYBEmvu1ZL+VYfCJpm3gq/gvckNCGF88IP
nZheB8Ci/aPeGb7TIKOp3HoEPur20tURDErwMlSJ8a99JYBf8wfTydNqaVAXt03nEDEcm5e2dwnQ
eLA56jFDnMYG3CJhlLCCrHjDLbOQ8KtL9uzrMWSPT85KchVjjzXhtu57gqUdomDC2qQ1i7uPQGuN
ipnaUsjzIpOhbK+CenSQi5kW/kDxDzpqOxkocmVgPRrwx1O90GjDq2VyyssQDXUG5RgPnJ1Un2bS
Mqdhpbk9KciSkhQRAIGB7DVKykb71EgO8igKvUg/sIbQblgC9bf63mDn1AYGdgOP+x9zMFmKIdKS
UiJQiZhIHtzpWegR6M04SYArhCC8IDYOFrc5GvMnobDSeVnSSWoo195PXfkqYquSDJz58zYop4vX
GOxVbzM7kPwlXD6JKwQ9PS+HUT9YW0ADuua/Pgr1JDdRBvweMaKpvJ8mvLUVV4pCk91zAht9FgOw
gHxyR5byfNNELNm+fWrWbt6hUYBP8kVcg+E/xuQBOwK74ZP6RjHmtcZlI2UGJEOex5dsGp2nJWlW
PHBtdC4FIa+M+iTWo6AF56xI9prAyFxJzmPkJnV9KHwfH3ueJAS4eODQGmiLyhVVy3FCbawShNsa
Eba2n8loj5sigprp49uk8v1TYgdOYSZbunUi3TcPdCRs4yW6Xw+4vd79RF4Ivx4su/6XlHjt2/bu
A5CqxvT8T9LgoHLzRVYHQ3pkT8fr7OllSq2ldz5TYoAOvBmgOw5gPUlhiT3/tmXFtTgWswF5akJB
/vEgaiYkw2Y+yHDwcqrG7VFsnTf1OEVtUrjh3GCLCjP8YA5UI7BLYqavM1i6ZVUTVQKbmdZbqtVv
XfnEyRnL190TVVyMlakUvHgFQYatfvQLz9P35ddYaXoMZ1+r1XL8VSaIT7iLcZDROJLqGfXj1gXX
hysN7xXOPXn0lV0BxvqCed6xajjk3t9m0Bvabahv6PZrOoiQmLFj3t/8HlPbOfBCjF2QW3lxPIIN
VuyTXsA3Tp82JuA8Lro1cGryqf5XTnI/WY28kUINdtR4yV5COZOl46R5i4qJ8HK/VtTRWyA4bvgl
nrF74lcYWUMLPgguvmNeMZrvHW1VjmOgD0MA1C5Cig2czahlNyhk9O1yGdQ0f5s7/WVQ5vPGQ8Fg
EuZx0EjfdDxoNYTB+dgWTpKMeGxzCxiecALAHYq0er4rGNavKSWDoA/H05tuPbHgN7P/NzpYsNaf
Blmv8ETBakIlv5uPtAiu+0ExaibwaP93FpANj7ulyRgyxh+xRmylzYprjQEcdpOpXydChuP/R59f
e/aeq3hV3/TuEnB/r6sh+pq3EFj6NLA4nJHS9BGS/sNIO0tg1y5PIUNQ6OCHC1y8HmGDWgt8ntDb
dWwUiF0tI4O/98y+SN8Jn3UjmsofktVNY7qK2J/TDWXzQX1vEs5eMG+QIMXz7Se3c947CBVTkyNK
G4k+OR3FV8loUEQjiGtMN7ByYMMoPNuyxxNhrZOHQ3iL68y15Y4EzM5o0Y0rWbpBa57hvI4eUhhc
SvSH0R/9GHXCIh5kx5Bw2qrMSuPd77WsSgKzzaolFnoRc//S3AdK3+/LmCN9+3ufaa61vebV+Nlg
8zqivQis5jjasWAuV4w/vTjPsBk+ZAiPbwzz1CQnxuixczTSR71RyiYqWy6zWHbdh0VJxbzYP52Q
MFWtaMQdloAtXkop6srPQ/ZX2V6WGWjO3slEJFXOf/QPOnNqlqb7ZZ6L12QZv4MCtzQG/ZtAPkBz
fReSy/NKsbK/7ccfyz+MZYzI7Afl832qzvZ/EIajZSkwr5g908DeVepxw+yxnstR/EvqswtXKg44
w0nZ2zTn1S2iGHxm8g7CJFPMkVXmfGQ3Svdf55gtN329RWiqP40epfrHJL8TNuVyJvwGtQ1GpzWj
CRaNzPJSY8IIte7qEmlOzWVFeJbXtOUf7elXOuQh2G2E9KvjCKQ6H2q0yRy91Bwzfqf4/luVTt1n
F4uSeYGB4Eht/FQIC1f60dlv1WggAMjtItr0SMJpBC8d5Jyri528rgMNy3KJmYeS0OTotkt+5RUk
V2nLR6Y/1ysaOtS6pxm+EcgL3nRDvJ35cNkrjia3L9NYHR9rp/VJEDTtxvpyPYER9iiRRqx5LrEU
xz55XeBuTO4fwVA+x8xIZFVWxm9yhCuLL01gAwSGUR3DlJtdCQi8/GlEF2/z5+gI/T0tjKb4faUe
2K+QuivFRm2Jbn9UITLq0L5xMic15wB/nC5fll0lZDV9p1bub+O3u5KeHTCwWyGxq2lLhZqUZC1o
mmkeLnDGMmrHlyAFHtUpZ4LeBMMsO/InEqtAXbvGgo5f6Ixrx6R3kgO9d6tODMLOOKhU+voyVySa
ok6bScrnLIZ57TFWAqjbyqt8BPWIYsS5JKhu9hEN81mAZgvT0bW5GHi+MQgl6L+p+NcOo4Grr+MA
Jct2apd/VDUh3og5gH7SXHQEbfPpop5Jca7Q7w3CMQvtMsellZhMBMZ5yKKBK5auRz3OkE85SwxB
4v3RyfT5XIRhkvFypTRX/tALTypoP9gQab804rlFRbdggn1ZqmvtGsPJHUxozbHxKB9M+rOVsSEE
w8iOEX/lrHxtWxNZxaQyBKSwFXPecNzP/GcPWd9ooIqDPg9tZbm6iG/HTpkHNjMnxPhd9R9eZVzu
PCD3ZoOCtlVuvFyQMCxpfbxSpC4Q1sNmN1fJZHbet8g/MO5x2vG2PPBrnaJ5jzZihOonkd8DCEeA
W6nHUhGkOuQc4yJ/LGmCDcuJsxZjJbNpw8cBMFpEEZl4a59P5KPCCepHd4eZziCM8s1ICkXKVXfD
jU5mVyfdC8BsPbwN4GIyBEYOJpG6lzxKhjo2MpAvHwCAYBgz1G7dQmyes7bph4qYb9y1sJTyXbrL
SOn5VUzlSjncyUtx4DpseZEewG01jdeJu+lp0hXUQBe5DloDBrQBr6A4vMHGAbGjg2Abq0UFrCSK
XRX7r3YsQRhie+OcbHMIBzsKs5Aj2CE0aqXdl7YYfa2M/E3HvXGklVhSabJWMdevKSqu3ZU9GMwS
YzD9sAPlUGf3Im9hSlIqV1YHKDViZDaqcd6jQdTHrH27gZ3R2GoSLlbOTCEA55+3rw/4Imx/vSNf
mBdYG7gwEXIYgVNKnlUEmzdImkEw0sKTNOGYqtzhwAZuSi3wV2H4AGgSak+k9X1vcnnUPfI81xcI
x/BpkWu5JqVqhTS+bCttVZ7hVLN31yuPDm7MkORqZ+MDuYEmyJKVqdkOu8vKDxzBm4J391CFEOud
RVbQxu/wOvcK2qdHcwWMFOE6idFbIHXT3IPvdAtXPngABTQSx+aNM6GcYqVp2kdw52kugW+DRSMu
qil0X47gxelazS0grqoyw8rw5JTzWuOv3tStKrxMY01QzaUGO0J3G5tpmPCqPjNyRP3fTijuBiIu
awvTS+gzhqt/Wv3Ls2DNOGlE086owVNgsGBwsTtvjyo/gnZCcj+JkpOpmmSyu47TBRowH46++v45
5MZ7oAs4ZBveAETbc6d/XVphSmU+zLa64vMq18IUy5R4YkO8TPnfU45vu6XRVvCK1ECxEwMctN5A
mgLZYOGUePGHNN/8xvnneSb4sZsYxPKeHJfwUzlegtOD/QeIxannUQI/cFKbWlX4XNramAPxHA2M
efToFdiLBKpa1Fs1HXbeQpOk7Z8upXUTaPkpSu+gEgHFzhDxmJkSkcJga/ZSGukQa6bimuZG75Fn
RyKeg9So36vw1hbWulynD6uz3S4Uom/PUGatogAmBI8InTS8sZEGzXtdWpmCH+mZr7dW+eHBSGRc
QS9wzo2oKgPLXni0Wih78mp6wZyqtm+tCU3+LL7v/Qdt3yo9DzRus/hBonnS2+8qq8ULTpvcaBUa
3nvvPDybkltDpEWbbaFKa7tc9LUxoZicFHrk/HIY/TUj6xFs3XIwatzB01vVhk2eVv2zUy/6pZy5
IPGDBRj3WstS5vCfaxpWns3GWph5t+5wCjou67V5q+JotSHs4QHugtr4ULR8Y7mvbHlr2zYW0Jx0
LT7yaupbUCAPr+0Dgqmhbh4vC1vXUcUKqAYyVijegtLKSXrm1G0O8MRqSDZdQOXtO/iTqzuoryHe
je0V2bKnX+bopt0aDCMb9jY6M1OJDmoruoEO90wW+wLyN5XVlRaIpPFGRjZsSmOPu8HNE/LkWAb/
RPwIckuIV/nI6izt/WCQ3APH1wVNVXxy3p6FVfQsbS8tlioTF5GjI8hOYBUl8LhPmf7duH3OumM1
cMWkWvVOqaWOZxa3Yplkv5jwSri3WP9AZRVfI6qs+TosFW7+k/kypPh63FpZCOr6VUNmTnLFie2F
goRfIuQXoNfXxp200s2DmTlVlzBWzdHjNr16ZdCFiGnoK62F0OxkoM3xeu+t6+gGGWFZPM66DASn
CctSpgCZmD0VGHGEQ2EhAEm+b7sYuFAcWWbEz7twlEAJ95YU7+N9/YYKm7ozzFGgsEm5owrJ3w2Q
8FUI2jqlGAsPgvH9CRbcP4D5hKj2oPDt2nZ4V3mwsapptD+Qd6BJnQ/OqJglbopjkfzdJPNwv7K0
IFC7uBanXjfcTa4O/UD9O7pOsl5378MnbhCPgaNoG8oMVmL8/f0RmyK7JDN+miLOawujQKletcKY
eE875NiHc2WmDkR4HRm8aR/S4ErEf/4dEpIOL9/VCMdnBJY46pfNr6qpQKTNPKVA8QM1ZD3YgsNv
8UTO4zbY8KwkCcq1q14+Qyp0J8P6XAyxyBPt2lF7aON11pFthYmwZtbvZ/OODeEmykqrLMfcA6Bu
c1I0ZEQoEyl+q0v+A5wG9LK3heMD4whhkqyPQBCOZDyXpaPszkJDYeTmVGS3xJqWm8BsS4rhSBTm
gDPLE+Z83AK3L6oPZtPs5wDx5hfW8jvnfwAQ9xfuueoCq0mw0rN9vUTH7SYNJsyRRPZOBK6x0my8
Tv3yEAZXj5xlxXiFnYQXGEnzkDNCBmeX+GnPFXKxZrPI8/qAU3P9TBtfIStRIybweCpBHIQWbeCc
9hlmAm2OCK9aHUDw9VcqA22GmoLMrppkaTk1mEEuEU8mh/uR02iRS8Jw3jh3REwIMTacP3K2/BtT
yMrTC67TuYSOhK30/g1f28+B5R5aDx2koUelizfFEveacdmcmJ2onyhUQ/gHBg2nzO8wJ0VjCSH2
nwM+AHLoxQdHUhIkraAdJRETNp4bAAdTwNVXJQ7MtpM5KTkCBRcnBcOYxYOJkS0s6wDyPFXwqDju
6a6Js8DFrnh23didiz0Ca483sjo58bi7QdAisbdvc5CODF0d4rrUMFEHAffD7+yGLB/w/ThgfvGR
wxojCsNVnJ5oPDjFN0L3Gdu+kghNlufQP0XeaLqZbO7yIRc6RGwtRibbdGg6ywVnfHJG1u/SRXIS
98SKHQbsXNV0ABWHaoQW0xEqAw3AJkBMWEN7SHaeFC5hWvUxHK8jErwstO/U/3+CmvzXqcAAKW2M
Pq5fDDkeFmF54Hv4YTPVVcxKhRjZ1iNnyQVrEC6rIYKCnWCX6TCpN+WA6sfGDRgiUJ5jJvNebvFP
ugI77DBqTDGr9Gr5Jrypb/fO+W1spciHuWGnnreHYHzf+HumLIi3JXHNN1gzsQJ7tTjhc5liAyqq
DzBb45VoyCfkQkZ3/aSttOGINKbMd1DDebrdgJbvigVfe55a5clvjuvGLLYUJjFyLGON7p9CwHPF
WeOROt4His3Rx5vNp6y+czS5fCAJt0OGago1x69VUG0GxmSEoFCh+B4g1U92GjndIVOyU77LCLrw
qi2Gj5Cy+NIbLRD4GID48mBjnWc1aYnxL0jOd72Ee46WNQhbU713OQ9l0GRYOmi+kHZsmjtjfT8V
8W/hrsjO0inKGx2t1cTo3OawfCZ/E+51OSq9jnSQ/oQkoh1hF+mauzLjBumROKH0U0XT3Q/iNjtT
tND5kTrOHPs8HhReLcb5Om6F00/2aVPWxlv4GqVLhUhVfEir+Fxox5D6mN8EWw0ptH6FDldTb6S3
Ainxy4Lw6jeK5NCnIz8PfGCKkZf8XWy7zdfo6zgVFsd7kHII0ogSjR43Gbg9KlaaS9ZKyVXa3qEW
ocRANkJg/Yc/iKyMWLe8JDrF+wTkVtfKZqBQsiUMbTFb0S8DEdSG0w1X4RPMZ/hphHitkMaYW8d9
KRIwq0AD8mtNExiphx5c3/2bpdcBxVyrYIA22Rj/DuI6fBQg6Aba9Km9NJgNMi4Aqt1l64PBuMTm
TpR/5eRzgNdz4ntln6TINrSOhKtc8OJMQ+r59tzg4pu2Zm145O8lICFaFSQsLOpmNyof5Q543a9n
SCqnZvdoJtjWraJcW6Pc1XhMk25XfmXw0cVfSkEzCC7Y4cFVkGnLB7/91H7CbbbHrmM7PR4MxIvM
+8HAuND0/m0YW9Czr1jUaW9os7zInSk5uXBhNGF85W1Mn3bOtUhtMnxgzGu0SD+3VMX9lP/znoBf
YvcPTfZX/5+CbiN3ffou6CUFOyKDsIH/hU76rpM8D0CMpuDXGRB5ooHa8NhFCKRBcorR60+zqFj4
fxtbo14f9rVYK2vug2QiEKygPRsq7Ksg7JS8Ka/pmcuox2A6ejG1dzpCWM2WscYWoWVvQES1zsIf
XDH753GXlBhBY2qYD8lmoMbn3k9ZOjeku8321+nlX2y1nrloL46DN0zSnQSV+b0uT4F/G8xS9Hu6
puXkooKKuC/6+9Vnm61LkVDjoLI7QLgtVOefVM+PdQeC298EQw460x58Euz6YNsePckpPnTWqEH4
iCk+5OT25DrepFl/1w4g1Fo5iPgnnhKvb5HFZikopG57jWnIK8W/vaO2rhc0wcNZVpdY+JvPua9m
3bTcpTqhQx3YTqSQl+qHHTV8fLC8VZHfbaju7hCsn0y1BF5pvMjaNdyU1s6k1Vll2nbv3zEX34IT
nnYnTVHjjmfax8GVVJz4v+Uiwv4D22yddBJSQPs4Zyt472g9vUVgp3+IUD5Qxh35xF949SJ3J0J0
xEbrU10MQI5xCegdKbdnTi9ynXAdWfAYaXN7ftanmwb0/Z9TxkfhH2rrSCXrzu04sHabp/1N0GXh
D4S+Y58glvISDaaQ2bYS5R7Dg5Jrbg+cl/KJcs/qFgCl4ouQ16UjKuTMtiMGTfa7AhZchqDoJmnh
NVNPy7gaKzsqDileNO5/AvGmdgEA/VzsPeohUlPTaqJgSMXq1FcotHfgGn51BZMkFTph1ZMTZQWE
acOMyFk9elZLwfXha+08W7Ya6Q0UbF/snlheaydIA4q0jZJzJhFQopRC+j+jZPclt2R/L/bZzKKK
6JtxvoGli8rx6Vj3yZ26E21lyBb5f4SGbjy4VDNxu+VdlXTStaDKFB5a4sySweFbxdEjb5nsS3YP
3nzAi+XuE3S/eUHqEGxWO7RvzsP6d/JIyazz5b1MjgOcWr5jUyWltb1n884DaSZ+o4upCrMBRqQL
qx4WOloaZZHfNjXCr/AO3nf89eLcr4DvWqJdUED7bWlDSu+0m4IPGL9csfeaYbTiuxGVPCa/3Edz
KB4tZn3IHZJPmmHZgPpfgx4lpPAVILXiWIZoBNOshWoTgz914uqS9KrZW5bVRBib34KaZ5VYx6Sb
wXUR6muvvzgzN760PkAXGxRvXP9bFs44TPBikVDs1tD498/ObMWrClo/ndIMjgLhsNxnBEfK1p9M
X96A/e55SoyNcweVbJXlyY5DlHGZLIZBlOUEXl3CqJkBcO2qKu0vIOgk72QBfdSXZnc/9Pw6GoJR
Ed4HAlQCfetYpIwVb3J29ct+ggHFPS9B5j2sRoiT0rnwKNUM9fpeQCsNvChpGJVIDQ8a+KkW21a0
Sq/NxGKYg5q1gF6X27rOsPFXPbzFcdDIsAJf+QSbw9ihcp5Bli0oYS6xj1lMGa0RVcB6/FR02Acd
NMSzEzdVT6KqfCYvLq4Xjh96XClvHzmLTpm+Y7d9kQijGM06pzr1Bb35pmwi3Ge+z0gxMX5JA/5t
EEKnOJ3Bx+6N/IOntB6n8RcvLSkR8ejcT9ddteL+vhMXfAm+SRZOF844W3BgVcaJMefJu9OSJ4wB
rpOlxos6Gs1nOIFgrCJxPLCzUU8HnRJfhqtX/Vua39SBmZgqollc9z7wxPlojpjzo+Xi+neUn8WF
+TOXQzJZZrfvP7DPTS+2MiyboXMf20s2/3xJZLjmbiZ05zjljnu8kABmapNJgeS+pnxNycvXtCi9
WgIaflHZhZZaSg5cS9HaFJl8f7IKXhlt7DiKVCbtw02AfYeZYiMjJLpIv4fK0kLavxmJki3A7jtJ
QcdkPfZdtUdp/CRt2vx7nzTqxJ4NAGfMp0WRFR/RyZqX0PJSjdE+a0Fc+mnAycgURFi1WV+Q+bGr
XGhoRCLGgTBeSPJ/oXSFVB0+hsev3fI5zgbGq9XBVwRmwwlX7bPgH0USMUQmRo2thhKG/vXxrCzr
iksd6ToOgpI7O+lG++xBE1gklA1+MxxDa5HHbfyXaFA8Zhdfk0J4vYjVrfpPIW/VOn7lKxlOZ+9W
d2lUmZVQ1WNmye30T18Jd1bZs/KDBs7R00pF+cBCvc71Ku81G08QErRkzFBoZIdtTCh2MOZ/emuT
MzoYw0bSz8nhQPZd8gjW6Nlkm7wwy6OpTI15A3xy/D7RM0dohNhGOWWgFYK89w1t2EsvXYPmhA83
b2OSp2ffgsJtyPGKWx1ZUkOZMI7QKb9JYy5NzdFRF/gHe3Kcec16mwTvKBIITh03Q/zvlzSbKn02
HkTiV/MN8m6rWxjK1euz1Ee1qZQP8cmfAhIaoxq0NN3EZc9CZjXrFZ3iJ0KqVGHUVd85sTspDqsl
ld16rVd0nKejemFu46PVpUzghh8Zfdz4Ju3UmB1XmuUth4lMazLjBW8yTSdoPdNO5LnHPNFsKWt2
krupT8O0NdlwzPbbBNsOk5Y0FPlNklYUOi15KJWZK+aVftMO+yaazFrewIvmoCYPKCESJ59pYxN9
5xZN+z4ED9GWpXDejKHKhplVnoYYwcwDfTFiHrjq0+4Oux3S3gblbKvooZdXFfrlQ4K5VLU14bm4
b5wHytmpk0d9eRMprLYFrfMgyoeNo8bqB00IEiz9rtqClRqwdme1F6G35EVuafmOZqza1ZqhHSEx
rQw1t9R+g65WVwMNkP4yOBEG01c7iLOPfkWxQRck5PBEL0n+NslKi+zt1GVUp6Kz637pGl3xarVW
snrbYWoJJofMgt2uLNOllvgw+659GR6yDkmz9OkUZSr9erPclhgrFgUVe2phGiYQyvIq0VHTpSWN
SZtJI1Dit1YZq0E8kVBljCUEZOovR4rUJxNu1Y1NcSHoWSMroXIASVlw3PAdY3C87rt3gpPG4ycn
a9QKaRxE22YiFcMMJ+4QO/6Yn5XGpP3FvfeIMo73ugom84oYkRDovUrH3hNnsAXZkQnKZAbB4q97
utcCszR7+ggv2v+JDU6Gr3xa+cFxPb9PUL3LuiJu3Saj1d/966VNIU8TVJeTL7ENItJ225gJ3RNk
x43nKKlg213izh1SV8Iz5FXNKiJC0XPQBcUqdaS02k2juBeMKRGl0+Qid944009VeyJIqukaWKS5
vinW1nJ5WTJFKmDy8HEJq4iMhKAl1X7k+JehYK5tR2adaS2OeeKhnUUCDww+UaW/y5b5owEQ5m8E
/jAHyJE2f7GUkr4DEx2LnFRsB60hAFUVppYC4qJ5FCSCBoM6gUwmOh0EQUunFm5f2j+u02nkB9A0
zu9m2KmO+hrzEmNYpcdXiqcCrPd0QEyM1YZc71221B63PRQlE4IgYofwjmkH9E0QFWZewD5hM+nm
a1oBn78XO99APQ+o7pZAHeDB7HJGdp8Mm/frxvS6JuQvQT1NTwqYWyhvsL+YSo5vZjF661hRGXhQ
dW7MXsJuT2utRF8rKCCO5tDxzzMW8xwrOvvpIuoIvjApsbsUV4ld0eXqLA/9k2Sf4SNUUPJsDbo+
mLyEM/rmUf3LS3AHjXivlhSHnV4pglnKURs/Et0IWwMI0IlEDh216zUBRIONZ50Q6lcHkzMmSA7j
LSN17HXCA2zcdwSKtAyykUeLvciW23H5c7es1D0rFfQ5oXX7ZARzrF9Ompb9XjeYr4XV4Cc67mEm
4Tgc3smCheL8I5wf+gsrzfXZ5NMaUpM7nO2sPRGUhhIJWua1HEr/Szr6rVqJcXwwNVbSm1++tu0J
tI3s3MnlaZYjmJNa1T0xXNO3gX4zvkZVFdmV108ZbKhNOJgCsEyIw+5vRT9NtelZqmqacH7TaIvl
84r26PYNx0v1Si2VtX1ddHqwyvuu142EnT8jO0LDY+2t7DG6av4SIuOW/OVKo+6dlimZcgPyNYuh
D/4Lk8bed2jipnjlTRlwB/O/vF8x7rsr6BSFg6sz4rzArYsb6q8UH5xNYbUdqEBWJCD8zGP7m6M6
/GmKxAMvBEnYK9wpuCqusmMxn1s9URDzpfFuU8V2uTXJ5EVfNAsXUmJgcWkoMufR6HdjOztiGNof
dUU3SrwScOWZEOF2JTLg9zPqTckoklS27GE2YAqS3Y6h2C/x1IZ+wycXCjZwNONThVP7hgijIEG+
BAkGPIJR21zfFarcr4x5FkCjRsuZiOWH5CNFQZ1tNu8EGdtUd6Eeu/QaKYctN0KBdK8WDHNJe5XE
6wN5llH4zlmXPPLTflMz2DIviLKwTHBQgA/YiQYER3anTrv2oamj1mfw2TdCQZOBG2gU9WtoHVaZ
QtUR1ZOrKAAGBURE0Uj5ZAVJpnwh1V5VCmHHksIIDMjIugjlyzcfJh36XO37VIfzeFqdiHW0klFl
kC+Mf6ZY405L8xYGdg+uBp4BI60N+ZQ7wLms9FeF1y5Sc1Pl88RqI1WI8UOv0zAaxX4pGqOAQVwl
iTm7Td+8q5VEqU/x+MpcrIbT4BDwx57U/RCRe1hAdH58pfP59djFgpEp9WqyvVox0XZuij4YpOL9
IgqwdENpQP2Hq+qJQePgnJhIQdGY6PUc3UlhncOLZdIpzhjxFTV674v8xQW+8jcJa+2jec07fHeL
uj0snheQmhK4Jv+Ac9o+fYP1bSPdV1W2zJJFKuTByf4lK+mSx5DOATtjwwbLgWBK67PRnIajCbBM
qo9ab0jpIgv8wkGD9dPJxzi9DLJaxkzl5VBAo07GrFSD5zRtOgzpdeRU7RHoACBKvr0TAKTcKtcU
OvhIuaEM+BO3+rMd91E1pwfpBzaCrAwu1SjIeTaEOq9nJ9A7I/EXeszZ2+4HWn2PWlirGFELrpzu
XN+d8HMmE3Sw/5qPVqZuv9ht2t1CgW5I4kA/1Kw/kjhgC8wkHr3T3RhqRpegYAqEiA/wqJ/DxiXD
royTWSwKnLLODAOSKFskSlmESN6N5Mw1pH/1h1jlYHeB/VjA6EzTCUm7ZTAxqdrwnxZ1GyB++LRO
abSqeOXIQ3X458iz8VohF1ylbqx39omrWtS7rQj2eTEsehMnSRFa50qHWSsM3Dkt2fvhTextZ2m0
RUaJEb99plDF+ZFL1fhPE5673NaDOqrfgBttRz/CceLQuhFgNktrf2qiq/xOXxvb8wHAfHR6xG0a
faAUAydDei8p9U8r6O2df2f+wNv/LhBq4PVZHdbzHf2caXidzkDTu7T22E8zkygqAXgBNmwMmJNx
N7ZDdh9kVnhY16TbGFEWGkbqCMjCYWWMmDm+B7J62+Eiz6Y6F9K2R219T7IWAg2fiUciHSJtk9em
p9e9yOV7pS4u3uLQeE1dFt9Ov4NfbKXNBFfo1hmflSyPT6Pcv49WmPfXD4RriW3GkgfoSbJ8IqtO
FF/HH2aW+W1LQsxSYNARWoWwskRxvXHiR+1GwLBBtZpthW7fTcQSLWZG1zFW1lSuFsKioX45TrVK
3SfCxyn5OQC48sommaqonBzILfNMZHmkc3HAJvNhXmXbgDyzS++nnTmiv2suUHY6oPAanmPKC1ns
0E3An0ajUsPW+/W2FvvMzDTZvdF4E7Z/jP38ETn1ajj1O5XfOiw+IatinjOML5pDs5qJXNqcfwc3
IxsYwv3bK8vihp/wOHYZPh1M8dQT1d9k7FDuOEZnrneY3eqRpr/sc9KvqPwtq6fOtPgovMo5ZI0V
KmmO5HtnorbYkl/3Ucje7x59azvS7pc7sz5JfJTUKf/MvuzAMrCKGFFDgeQWLZzPK/pJqjlYfe8a
6HPZ9eONfKo4fuyRT4IwxaTAiLBPersHcbLrc1QJLOKvKJKl99pYGXCsXup8tj7Y/JjOBk7sFG5V
NorxaaMtzDgIzELQhJwYbIcZbHVRAzgWwhgiJ2mN7fy9Y5ao9gyr0p8aCsfDNanQ/JgZn4j3qhnB
tj5MllSagnBGIEJ6v8B/22p8U6ozOzuqLuXkc+zq16r+KqvmztbcOXaGPkiYkybY3pzIJSuB2Gy7
3V8vAmY4TlUp5v0oZ3peMPN2UnMYpvbcrvyeRDfsFaVozwNQvFO4CoGlmIxvIGDksgRWve/na6HE
m8kh/5Kxr3QroYyEdmK1dqWvbgKAKiTmXbNnzV//C1ed/2a9CMid/e3K9WQ66tiOVGggKgGn+JPH
xfkcE5rLv1e0IrOjCSR3bx8zFKEUBu+fiFrDF/VwtV4Ayeh79tNYGrTkVbmcFz00vwuzf7smoiLi
E1UbqqyEE9B7KqJKqwFZMaypGFDwYB5iV/QEnEmP4Wf6nhcCHwBPAEFMlzuBPviM09zqkJcAdVfN
nHZYe2LnziBXGZJOFKVRhZARWeLhopQ3+iOIDeBoFNK54sotR2lM61Yhyw7jLtyTL9lkNSRp5wKi
I2nFQ1b4mYRBwqoGAVdw88eZZ4uAiJw9i4L/yoIijKpra5UTIzVtSR7QKNu0FJAg6+U/nk1T9FXC
8WeJt3qtxxqn9+pyETn1ftNxago27Wn9kXL76VLqZ+aqf/w/gke0NH1m5CtXuNak6C4OxK1F0qCm
R4wKIMifCvZrpBlyZaddfB5cSlWuEp9RuKJEWukuiDOWYUKz3gTWDALrsT4+zbCQdoKBXCkY2UQF
Pc8ZNoH0/ukZgWDMKAlukh5bF9yqi8m22JlcnwBi6mf5DZzzgDH0Y/KPztDHVBMUFKoQv5e2ImG0
kao6GCPlSgofruzmE72dala6FQzuf5NwusoxDNtDE2xgFsrA4B5E1BcxgOYYr2z+ni7WHx5mjcBw
DPeSGFoc5vID8kAHO5u1u/9gZssMwtWg5dtxpu51PcGF6JBTYGYxfKsszEhDUjuGleVWfHw1hlKb
SGpdwT0hEy1IpnnJPpyygoqHk7nGcy0O5hL8JIJwG0BcN1ghSQZLxF/IdUL20OEDQ5+PPbFg6MYw
ztc0hIZvhApkwFMDY+mvW8RBABAC3dADTAJiZNURcMFCe1fcBsSkhhGFEA0l/7tuT+o/9eoujW/3
BVcFkgO56l1aywdrFymKGZGhAgTOt5d9aKjAEudgKC2ccRotVmijKxbx27X6BUtHLCQcPOAqnqQr
gJRomup8EnUMFE1/kBnaaBGgLfXV1oVu7L40mDe10HhcshX5ck/QJRvzmcyo9e8iTG/2LagSvD3o
7x+gCVbOtrprgaNmjCDSatEOBuZ+luKIIkIUIg2a6gjsa0GSF4ogKisTUrWTwl7MOWXnWRaH87YX
bm/r73IHeGnS9lX8apTebqABhAj+q2tnOfe3x3/nfjSWIGdXen0g/D29ZvvPr7aosYljKXZGI5Yi
zEdVdp2Bqa75qu0mYF1WWn/Jj9E2CTrFmuGtQUw9pWLJxhzAyZbUsKU7CY9e6TssqVR9/RO0c2Dq
gy4s/8jjU85W0P/d6ZwzzU0wTrLUXVPM0oedCyHWNBhJFNao9nWFgZfUbOVw8ElTRnbP89j5tGXy
sYYVFlL6TvJyQhl8DtNcRY2ogyDZ0ttbXj9Q/g80Acq9SkcrrnstGzwTwtcWikmrQr2qIpIvBBT6
EGKIugMBGBe1reFIPzG4KFPHg/1MO6tWlifK8WwRpZoaQNOShdb+TrEUUcJeyHux3Qm1F83BUwTZ
zsVLtA5YQ1GD7F6JvJSut4BUE6ixmmEUMcZKlnlkgXUZVSnMfti4twZyC6BzXcTs4hWcvGrassFM
hPNXvFaKtVfeXiabCujA1AomWczaBrAAI9ytMWJ0KtLZTU4aB2MopEh3UyW0coPDmjpNxC5qZ0/G
X1dT0t3G0YmCzBZQciV0p308wd3IBjwG7TJx3DYIFDMom3hix9KNjnHILZ21SQ1Iki+T6jXyt7Q1
ck6lNy1ftPKu97K4yKYz6nefJLU+wcLjv+BIaOX7cthDgbRkGOoPzsXNAPIqL2GT81MxIyitCilj
2tdDU+24QttE5slc/ZTAKbRUpWLPaygOBlfH5cOAJUAnnAHzgPw+S07bZr8urrlkVV7it71iRrF9
R9QHvM8rXMyXVSbqx1+3ZcXeHhJJ2VeUwxw0IL4JkZs+dP61iSuB+g937R7+9qw9ia+DFpjk4a5+
q3tVaMQ3cqcpmElYxE7KVDKqJy3c6Om6gdz1UzzTarpaP5DdHRiHjDdMX7WZE/vafYOjtbfA5M/+
VPAgaCmCWamNUHZblIRyuHxi+wGtx34if7J5PcHxBM3MsGDI4BimmedKZJyMfY8q6PdHyLYIzs2V
Yuvz0HAlL/lVkRbhtrIflb6+9WHV+/c9hjzyxy9gaGhzPA3d9HNNQUvtE+13JvVup2q+hs8t+ann
PyaxUfv7zmH96p9w0ISnxR4ewtbm0Ij26MMcbUCKKQH/azQNmBwg+Xa9dShFbQTLN2bjdwl4+Con
BtshwapPLANiD5PhYMCYRCChihO9vxw4HqG5Yg4/Od4t9jhJ9NrCxBA+GHfQcCRZvtyvCtaOPX93
aQd0QphsjZUtm0Mlq2wPE2acQuprlxT678vGenkmbDk7zqWXWCscHgCcKReEB1wdi22oHUZ+NVzg
MB7XadP/LvARNTAO4cHy0Q0IJaBd19JbMBmXk7xziMag8u2vsCIyQzbuT/ukZ/qNkak0JfEdH4cI
Stscn/pnEZCMJLDPJEZIW+7YLa63iHQoa08z3XNzLR4P/X+XkYnBUZ11LUJX3g2XpO+EsFRRAF+N
irIiIjSReeAoBdRG2yzSyefNKv/ot1YEP93VoAvKbxcPyrSaN4g4P597pi21bPL8cbl992DVEN2i
/3Oj6iC+neLILiOjkCvk+TI0jRQWJWwe3fWF8cXsiYdW/ce10olxKnErZP86aC90i3RSHVFYi0QA
Q1kwCiwzN/f02b3adAtb9Nu3ULfsqr7eEgXlC9XDOUdLsN5J29lLlHegOBcOqcs6bfAv347mjr1p
tG48dPoTerBA1TZLWvm0mF6LQFs4FMnO42nfad5lIGr2xAdz+4vrRK8E3XEU2rIwXP1LoE1K3TiS
GxAevY2pbC3bYqXC4j1OwHZATs3tqfM5f76ylr6T4vvVqdR5l77sEKQ5DP7J+GKFz2hnSisoteaD
6vin14j1Xqr0/Bq6U060EwN9euseiTm/o+SKrCUIly6Y3OgV34IL/pWhrOSp4XQs6Z1TvSLjLBh3
d99uFTI0tpAfvcV77DOy/e5Yco+8tDq9nF06KuqvS3oQ51awK4hV6By3mGRH9+iydZNe/TNMQGLl
+pOBT2/R9YUHrU2npxjnr4pSkKQonQwl+1Oz0eUhAOIfvg5C41SIyrJbvO/Dum5eMXzPzfWN4MsF
agCR249NriruczTQGaj0Kg2BlcLVmSGRKLt81EaSgDcEGqh4ryGePJkNyVVLuOFjkXqtFGys/vAW
EtTuJ9M5k3juTawzHmTcvdOHHaOwdXhPzABzdXSSQ0blZnnPVLu90yqr3mwrhGXmSnTzq7Nsmg2q
s5AwTe7+wderCd43TVN9BtoVW5JzPreJ+Ql+ZHeXQ8xKXq0RhabMzA5j4qrwU4CKs+/gcVCVG4i+
jc4LtUCaz/s+eEIsuGkiHUGaTiPLFG54wy51u+ljhSjQrL061V3D5fV5toNdMkYB4Jh3l77vEg7d
qtZ4bVXdmWmb/6lOgWSgRJXnz3MCsqB0D5EacqxGyDKtq+pNy+Rh0PsSFqMLS1tXujmS7NGw56B1
tEPehbBOtEANCFyc3esM5wIi6E7/fhw+X7w4jcXryvK3if68gCqlbisFD+6i5P2Gg8zYMZjFZATm
vnI84ZMLeoD1okSGPl8oJgXmAE5DaaaiVmQaaMJQYUj5zuybhptJHN9RmrwzzlroIqU/s6rvljaX
56+2fsEoVhduf76UkNz/7tw8hAcZjDm2A5lANgoRa87d8gXIzc7zZb2vjsfM6chmyVgD75YgoDKr
18d+0I9yU5m/26zT3WfdYVfgMGGH9lPB/pJoCv0nm4jDWfvtihY0+kdvesa9ZPaT+jhV+me2KuQl
XTlhSlsLfwJdHnsk33U4IdwonrMjMntyB694vXFwGLpzE7iCzUUaS9GjbJttg0/Ub+VTSgEzHNf1
pSWoA7mHEBZr3m700/cMVSiNfCcASNqgnopUYg+FJ2nX/y+eHzQ6CRI67EUBOSrAuE5qIYtVWBE9
ke3qCdcY7WJ9bM1fEFd+Gnng4dbpm+KQudOxKh2PHWHHm//grBKmL0EB38XwwudtFiJIhR+Cq6Em
wGZjWBB2dlKAEH8OKiQLMSVS2/5+T3WfOJBtw6VQclzTggq+8ctmpVWjoRVjzKFTZDxo9nEwsbiV
guYgZNs4VR2CcZlCASVl6my/YgXtJdqYQIVaMcDhgTtj4T73dl/ltamgiOqJdRRGJHWQSFEyAa5y
seq8B3W2cBhQv7ZGkBrAhU7sAZ14Haz7R3rz08iy42+o2d795D4drecWFxJv/TtgpGuuEq6DZxrf
MbCq74cPfLOjhKdhV7RXUpV2zT9RS4EF2ByN0Js9UUkHB7AbUlywWWATnVeKt4EP0peGLPjptPFI
zAju5+T+WDRSiTXMT8gSsrJBMz2bfePy3p8gM1jXcmNpRdebN6Q1CSw2RW+1QFVg/IpJoFmpLHXo
H29LHMbTnINzMDQPPvnXJ6EVTHOS795Af2XnoXkrwCcbVAt45XNRS45MIokrnKzc4sxOqofF2eB8
IZugef43oLW0SIrK3Dp1smFCFFsGW4vfBIaun5DSzLwpxcZHY3K9o+n4d4OcpEIRtt+EWduF9FlP
ovBSLrlqmt7mueZH798+I+2mjTnfnLJOq8jNConsmXHm/bLJWraFwrz/2APQchqKsNKGL2AV1fWG
7nR6sTXh3+zPZuFF7TJCYbpumzeCayMLv5HNHTO9yh9xT7BJFXYYMUuht3H6ZbhnkOdK/wsnF2sy
vTdG+F3bIYSklZ1TKPfgJPBfATEumIn024E/u/0Ik03DKb8oENMTD/uRxEskSRT5lIf0iZIzWF+0
RyRktEFQxoOEy6ge7TGJqEwiRKQz2Y+4NA+cTW2x7QTffjppfU/E/jil8A7/WZCS5PZ/g1Rjz/DC
52gMyjOf9j/wRNpSUD3qz4IlxLepWFMo8GCabmKeEEdwfi1HdBoCS7on5S8If5pTGeo718bM8sbJ
yIOWeKnE+rqkac8yhxQbcdsfbMhmdPYTKUg2WoYj9FFtj7PZIwstUO4OL9QY57rCLW3Jo+4KO/yn
X+NSKzaRgdqI0S7RSsjJJVxbeRU1ea9LGRNEEF42QdvuqcSqH5d+lW11ks0jyDEdG0QVgpmrafay
1aPJyyQk24oOH9EWZmmRiKQuSEI+UhkJZRoSbyPxTClJ96q4ZH8YMK+6hMWGvtyJSOlW0q3bm2QE
Yj8Na8U1uvuqIvHtAzKG8yUcEI5NhmkeWKNBdHknpeRtDq6/ACP5Wt/lGbXWTs9wsC/cxlGFeYfJ
ZpJ2rOsRUZPYlSjSjmc9mVz0FZ3ZIEcPgxEi7z9/C1qRAEVBqggNR10hQVHZspZ3opMfULWEWN1j
VzphzIOo5bHep9fugeN0eHi2wneLyFQpq0V0TeHXwsx4Xs7E/znx7PURaJ6cMrgY5pO+YXWu/th/
VX+jQjaLHfoaWdn3oDzHVDRf/uaqrlfV0REPb2+4ucPB2jA6Hx2Etu1VTYDeq+oR68/oI78nG7zf
RWh6/0TdpXBv2CgcQj0gHF/ukHNAwL4Pu3k3r2wenl3EudExqGnltZCEcl7L7tI0R2ezn9g4phcS
HLRoMx6FMepzfrXrm3QfVsXb34wudzGoGAx2XxhA8yQ8ipGt9GeQ/3vs/dONETTP+r50q42sPJch
n0UCkGOqj1IEgUaKxfhRS7zO7/HfJOkctfDJ1Jdyt0ImhhgTTI5Y72y5VY2J3y/1pfUndXBVG3oQ
15XbZVdfO9GZ62/bkDyZqyd08qhlAeJ/ngVVxXPxhCQm/TyVxZ76OBA8z3UiUCVZcR4+JIYU4ypz
HIum9a9o0GjK3VYpnEUfGXbim2h1jKVciI/m4vgzEMeOF7lS4qw9zflRTU+ymnBJDyplUXWvhBs+
tWLruzVvZRh48YTE0kUWuycqEkCjb0jMUYBHM1+x7r9LDGX9KCbrD9bkkP2xX/xDTFHQ/5xlecjH
rmVzk3Srk1/SYlNWQJ/FJ5zMYe76F+JzyaDx14ouqOwVD2fDp4DoYxfTp61C/9R6T3IkF7VjWBA0
PuhgWBJ/o/iEiDWPUekZYePZyNxngXwR/gwvqGDeCJyDw3q9fpx9BuDq9ZYxIR2RpO6gCdoUdV8N
VCHSDmKp5MqagsRHJt/ibwU134pQzSV6JawNp3vzflPBm1+pA52ZuF7FsRD92qzJOZbHdUjixkhB
kDFOgVnJLu/pTePUcCfZ/Lz6xrN1msHkX40CIv0gxQpVhBu6618GBemkEhvgk1Fk1+JGGpIyuVOk
aNwI6dqgXFPTlSGIL8IOvd3SPMn//BaS+D9WjoTyt0oPJbB8GzdS9heYw0aQWauoCYCRUY0HDbHg
6WccBs0Ku8en5WFASQOPtOFbvxkNBQ/VD8lC7+L74l2Eb/qaHU7ciAMzGhPrloPJogE5tLrUXTwa
1Qc/lGPdMCwU/aT+v1vGzF+AU0WM9F4EiMjII1pL4R+5B+lDLW7yWrkuMDTvQtyIAvk+9JHnDdV5
dMzNCBRm5CEOIrMmlYVXindSST0R5B9aDUBJpP+ji+IfsY/2Ul7dqQKMq4rnJ+14XPvS11uvTuWN
CO6HtV/tX+N1vWu+JfUyZoW6FLHqqfnO849G5x/zYU1Q5JaVy2G+HfUgN+gu19p10SN9t/LQfxxi
xn41A/wqfhL3qkyI6CnPB7d7qgpDyF5FtrUqqIrB+u4o990z4PnWVKZJ47KdcQAUNxv4A0dZg2RD
2pvkB3MgHSQesIpVRI+mFcMlJDz4UBMslc0NvNT9JDKGdrp06vs/1TswH9k54XDf+WYu+pTAaWng
NrpOIwo4K8Tz4+MGvdFdRWlAwk9EoADE+PGYjX4Y0HFWcZ7s3U1B2+Pc9lbSx+oClmeBj6h297vM
r1oJKAyi4Uy0he0KL0ujRd+D9nadsHHQf1sYnpvLrjtyNyHtTz02VOpj8rILvmzU9upDD3rq21cT
5z4zrsDCjJjisYD0YYukw0VmZ7yrpVtc8LFmyGCGMk0C7DPSk5KUJH6nPyIWEZnBvpm0MiqE1JZc
xD1arSCk8iObCsciUkh2xMbX0q1O7+5bUYYzjHnDx1ZfKFetQbX4xGwd+6WVKT5rVF/YRcGPNE2Y
Nibw6EfhMIoVJZt//pUCXipafSjbkaoE7uxbTqvKCcNSHXGK+b0VXfP3WaMNG2lvMXPkwH1ElfcC
VzZEyPO8HfOr8MoHYOJsGpaa4wQXfNW0u9hE7RN3pXYgPx0raAFmkVu22BGHU/B0NlTrWikK+aXI
jQVgArQ3wEd9pPd0+BUhwcOR/tOQkMUOfbwDSo7q3HXra3/JFii+vzptkuvrgTkjYiLfp8aMkg4w
bntIexni0DG/BSghfZNM7e/3p2Y4eqNk7BW8wIBOywVlfDTSYe+MJn6UNNGeMWkjFVMTfQYksHJv
MKgzSNviNLK/yN/l67IWSnxC1dtvFnsFz4+LSzHJlhDXfiTdeERrBQgTM5QI3MUlYw9HP38KXqSg
j0fz5yHrZ5ffbGUZmWCa6sHDCnjS3w/B80VdjJvpKfOvkbTfOWO3ahHbHAvHbUVxx2zqlQnq7ZX3
2IcdPr6+N+CeEq4t3CdhF1t7TosKJE+q7ooDc6yY1KQ/7AOIPAQiHC5q9r1O/18RVYTRmzV6eW7q
mwW2I/dJ0qNpcpBEZAZ7usmczNU7KB/cXjgV14SqCbeauWOc7Zm2T3FluVEd570YuGbwJSmE5GLy
139lPnA+XB+IVYH94bfB+4KRuIcrI4a17VVhCC0uDe+TaP5/0DUYl149IEMXZxkaW1TeJYBAGDHH
AyCPbf7EAjDaI//OVAfdBCOPI/q6UwcQ6W73RZsEIYsrKVUsSxtxoDtnEjeciF1YNKiAzP/yMKBs
6bbBpEREQH7Ncp+u5JV1NBLX9F3eL54L817YNQDWemNVJsNbaefodLbWaev13q6NLedcBKwzAWjv
S4+785yAiyhiviLC4frMch9AjO5IdjgvbIs0Wk6N0AWu9PaDiOayrV8iZmnVElzywIHADG0yq4U2
rmEzvnNECjpINzo5WSYjT2xIrb9IaxRBaXE6yw+X7t2vO+h+o+Yvxl1/tc6YUyZ1/Z7VEcXtmIPD
GzrhU3dNKJWR6FrF/r6L0rO1me96MYi5ZQH2o6m9lD2QXmjlv6Ihl2YyQt7F6zIR4oS6Y2iogzug
Vrnuz69KJcqPB+We4I2BmKMMaUAFbwaEDptYH34md9jh7qyrS8x+3LToz5VxTE/qEFazNPNpwtw+
fcDqgDeMVbdjKFoa8lijuww2OtlfflVPIGdbWgTeijsC3sSeuoBf+tFcR1fHhqsNPndHG/9bZHEc
LK4AbRkU9vlZkpS2gdNmZtSV8UBsAJpZxC+V8qWY7Ig165UmhIMtve20WU74awjTWNF1B/pbb2mc
D7qJjm8JquI2CvAR+glUgkQTvO75fwBNpiPYKNbu4YpJTj3X9iD1OS8Ex5D9vlJnZdDndc7QFEP6
NTtOt8T5oGYknq8S1axjDzEylD50qoBIfsvQnPU4eoM2DTZws/m6felMC9oU20Y4JkDlbU9P8sb2
nhDJI8d/PFYgQgmUGpdPDHMWKdyfcj9SamKKfu6lci0aaTelBVTR8vUh8wxobl+oStMedR2r0KXJ
seYQKJjFsUAs2MHXo0GaFtbU0pPDWJPdU9vZ+RoAFicrnrvXqx0HcBjEUFSmQ+Lrx46yXV/vUAu7
q65f+BeAIVHcokuRIy5dR02C27EeUU9gNlkQhHWHafRKsGcpWkgLROMXVHtJYTarA+vAD4TqFWwY
lfpLZ9dkMw1U6KNen/24UZknSaY39elDzUV3BGHmSPv+n9OOUlXyRH85OtipeByx5/6btKr9BFKK
9i9EGRj5u3bS7eLH1B0hCufCHNLk2DvZvfHZyuS4UmBa5e93DfQdfhWgntFBZ14ELIQcZQcxa4/p
8xRI6Ya9f9UVtEaMHPYM9heo6P8jm1ffrIuUuVk7ylUzSXVyA3FIVTqHRGVO5Jh0IhwOgx8PHSzH
I3c77/45+eAELBh7BJ/r9I1Pt627lBsER75/zDTQi51BvpF1ndd2zzImG7SWV539CE3z/xCJFqRn
PMtCOGI/7nqX4CQupaQF0nLTLk/K9lDReOtR2FfqFFt0C0Avhmy2CwQtXjbL5jKonVzPdEX5OVN+
KcIOSgkMwv4WdkChxAgKOn1PvSFSLo11WiP7HEpVO+9ePNp7bpbTqr/tzBEvkYiVHFhZJvH47YcB
x3QSNbMZ4Mp+NXdOeaWptcmV0krVVas3jflyZyzRjfTfA2jW6ZJHa3xowaHX+kEMDoDGG6Gzv7qH
vQqvQwF2cbOojfUdZ0ByMrHDGHdzXbGABaDtm8Gt/YkhcNY3v/oHoyCF2kLcV9f+FPEoSTNV1BpN
voxnmHcfm5TKlxtVRQk556L6m3W0xc9EkM6zLmDnHuZBTfLfvKRZHL7R5af6lIyBydnpY8QjhgSh
QBez7a5W8bPl0mgrtOF6fZXYKOw2NN6+r96wQO2yegDo6+wLl2Otl4KPUDpFJfllfa+Iip//B8a+
CclBdHPQ6xUkqInKkFESdHtQUzU43aKW0c4yn/5NCghcv9BKHvbl+GkTdlELcRu1nsA+ztGjhHQN
LyuKjqi3u0IxGepc8S/FdKH5Sth2TPMP6zn3R442pPxhObWz329spB2qhLDdkzI/cm7U6QYILMOG
aViKXO4mNWv03OSbmzcNlZF1/n1FMBgyDLY8NcSl0KSzz/ugTcWSzIgnBjMqOtYgs16s0vByBIUJ
l+46fWlkwxuQp4h04pO5uMHYXQe1SLYegWuUjCc71RCMoD/P4pDc6HwGJj70BYv6If5m8Bn3raxZ
pbFA3Ulm7Y8m6r+2fpwinyhHawyGU7Xjbori3Ol5EqeBASb2uC/OMHvk10WcFJFYg+t+8g6bO0qA
zFQDlWgt0VjAGHMvotso/ZacwleRtfq8wSsL/FvuVMneOGJvHmVdZu3MFdfTbJIlx2S8Vipwce7b
c0cfs3+pmb4Uo4DycBhcQYOrLu3kPWFBetvTOnifArOnCo/QY7xspe880ukiEteLmGzKm2V1g/Nu
DNVtjbfcUdBzS763GRgBvaJZY6yh1CwQy/3k4Emu/c0mwwGiZceJDXZstwqaYrVVnUUp4ElMwSEk
2Heo3D9X+6nUhbYpPOTJQa5drzX8Aw9xlzzgJcFM8bt0Bwnn94K7C+W0iyEmCUyAFPS7FluJWUbW
9XLy72L/GRvrIrc4Vr4cxA52RjxWyNmws6ni5pTdTZl8mu8vODhbXIdSfbp1bsdMV312BNMSbMtt
GyKkgKcULBjPe8yCW8jEq3+P5Cn7yo3V6beF/6ZtiW33cRF8c+mvBjR6yjs+zaRiPlYrvWZaf/D3
SS7kHP75rWl1QR/cDF81F5nyNqaO5YTktfkgcrS1BuZC8OFp3sHDgdO8Cwp8tPedMZNYR1p3jQSZ
JUJ8g6L6CY4VVtu5RGAkr7joiuXitVl9w1bf9gzAJCJ8vrzGXUbp5ldLOlCcusuwnRqXp0BO1UoB
NmkOtQUzQQKq2k0X45Cf1MieAzABV5oYwC+50t2GEv7MRPHvrPOgbkMP7M9HK9s+ph6U9l7WsTjB
IN+JJisweoYx+X++z/lM64ZucyMBGIXMRaCB6SHsubfQb1KgDdNPCdJULJFV6igh9czzxK2TVDwB
iCgdkLQDfpgq3nEFJK02e91L0ek8U5VQGUQTx9SpYVIu5nJ81TlPYOhiEoBXVfDy/GdVUySR9D0G
i2AzwDlo+GxddNPoyzc2BQXNuqeIxVS3dG5DX5NICnPsxhIlwUDNZJ+shvO6s4gKz1lpPrVjXT5C
KmFBKCM3M6DADN0F9PoRl1Fw5FJ8cyBy4LHI/dvgRzSpWaOaGA30mDnte6hkHdezN5Dun+lUavyV
s7UqQgUCD8m42ojRxAzAdOLmigVixi9+LCwsGseMqE+/vsaYPZSEYYJHLFMrRPcj6Oa9iTF0mIQM
twkunZRhM+XxfGKlbYqRKqt2gtPDRE35izhDVj5dbUaPdoCxKBJ8mpSy+DzyFmwDwqxXLtEGoEpo
IWq8nZ8UBW0rN37WEKI+HNHUpLnwtPnl6yAPF00mLudUJG6n848X11ZTf8GGVnmK4fAJYb/yHkEg
aSUL4D7ejBmvW6GjtXWluF7Sdv+5StkwwdJjX7x0yRkIkvAlu6XekgtcHlMvUMnvBUMoCv2ZAoab
zqNQvWYPbE2ozASfMiW75Cnx5QTkMQsa8zXeAoEVe2BcNH3Zh6wtsWSdgGTOxq38AkUgtZ7KpvZ8
hM4PD6CvESKt0tG6irlGlXsgXHyHxAqo7fde7Jxrk5Z78eVBoFyc4fUeK54NWs0j4ypnL0LGhZzg
anxxFrl52Soy/+hxsOLCN7hqpq7GEF3ibQkxdT3UnvfvOIyPOruYMRJD8L9NXlaaYlWMk/xyfI2R
+uIX1bowq8KbkTzmL66cWa9obT8uB1Od6xCrtPoH9Q57iKlDhMed+EdZYZLPXuxZFy/rLdHo8VgJ
dct68jlEGHCYkOXsHBtYgW0Ra459SkNbUnTJuUTK4d2qu83S70PPvWuGMKoTVlVBnQRordsamULx
4xmf0thCtxZ+hhcCBwsQk3cKWwLUppyRdlPokbo1gBwxXaRWIC3Eo7C7qikNqkR7f0LQkVICOPF7
OcbwZhCePYprxA5jZ7aE/lRhFPeJ+c0iOkdFQe4mCnnqlkQRyyxnqdCIwuCo5B3NVSUchFNSnHFm
ZVKpUXXJPEEseOd4zdrwfmcy1rVTFF7yOwadO4cGiJBtTrb8gdxbEmTRMi6nSrBJfnKA3760OlHf
tsTwrFGc6ixAgoBFABUwi2kfUYcY7tz9yeUUGkLZ7bWuPhI2jC+w3gaflHWZ/mx9QCQNQWoZ8yXQ
RdiGzK8KS/WdL6m4+XjUKUG2m17TiMrgVYEEesqIqzUujL4L5FnFFHXR8IkU0F6rAjatUZocWTxh
qV4mzDw+Cm5ExEXSZZ2CK36oyPAJVC4EdRM3bT4qL1mv0BM8e5N6t55AVPwo47nFsJ7x8ovEJSdT
D3RxzYpFJgVuycA2Nt5lFSj7xLVO1Jb/yu4Wn1JAFw6pH0EZZ/xdvnC2OG8btu5e7/34Qwf47xK1
gxu42Vrs0VvoYdGhOBhbP0N0kTcPn7d64JBT0lxc2DwoDDPUN+XoUYwXQ2FdEySPa6p2s5gc8Yt2
pAsstOhtPlr5cyfQm7zmmPIPP5lPF5fwSda0czjamOMGXQZAXqfTuFiofmwmf8wKnS6E4rA7e4Qx
KAct8qgJCeEcH8Dm0MUhfbgr98+mJNDXnQg9Yg9xILSzLuv4g+htR4Bw7/ooSuOnfx/njKQTQZfG
EW6BJuD11ojvGbq7A2C2og6jTiW2zceigwTi6m2xB7BTo9j6o0WfwoUbLlY6LhmWGqJygGxdDdMT
RW7o4B1hSgVA0Y7ILisGEwZJyszanf4v1hWCG7gLiG7ESoxdEQHAjlBBr7SR3OrUMWsh0F9h61kK
z7thXud28JNo8ElW5gCH1hS3QYriramdSuqmroN1OiRBqxHINCsiZRyvp6Vlb32caQSnRBF41mk2
i2g9aKMozTASra93+yiLZjHY7Tzzr0S3fvIrpC8fPSeNKH2RtnMp/o1XexCFZpWJvV1tNEwcOzib
yeBlMkF44BOqLp+LJy6zivPB2Q6As8s1IBk3b6zplcM1e5Qe3u8xMnOq8MC5/jK835re3lvZkd6i
vt/lpCzzLUKpl+33cFeZA7Hvelf1pSHx7B11RjTmEFV1UWN85Me5Ue4UCRqUSQ2g3AEIuDCojstl
Rdv2C1G9bLOuOkwHs9NhTgP5s5zLyHvqYBwmXsO06px4IHmvpLQLu6HABQvdO6xwLfSS4I542d8Z
ug8CLz/nuqiNr6hRSNMMxM69yqpd+E3mUG6sVkIsI8Bti70p9jrrwZGnxecdNwKjDy+w2AcQDm26
0jplXV4F4fyv5pofNBer68NZkq9ll9vhcRpGgdz1D6TGOMFBlyh/YHq33clPboy17GWYg+6fiHrV
kKzuhWZ99Caiw0jgwZHzD8VQovCmax/6QiOX0sMb6z+cG3mr3PSnlBAjuW0dCDob0i5sdSeqT8WO
Cmro4U1gowpgxho/yagin5haSrI88FHHliZ+X4XCZi/uBtGdw0b4s3vJEzDsofDva50lS0GxJzex
tuREEmmv2XIUpUlfeJtk6nElF6U6CpN8K9h4EEakWMrsv1zXrmT5fRiMCN+Eimzhdokor9c1gN1I
7phIXvOozjFWjEo1DosfPj32SUZMR76M5EhHWwSAp9bXQBvmvyF0AAb3ltNKavoBENRnOjin0H9d
I7L/LCId24Azgu5SIvi0Ab/uPqgpn1xgOFyCFMc/++/qmBG8PxWrQWUGcFLlrvrTtaMWxzcsK29T
HzEYSDptvJST2F0ajgkU5wbmp30eKdx2HzfhSJEp22H/x7rgE9Qs/uTcEDEka9xaL3Dpn2AR5Jr7
JcGoPRcFth9TL5PDu+VHIA1Ug4W3+FlNob2y4/uFniPhiRjYh9CwBe/ReZvQMcN9N+wqoe2jKA00
fpEnfYxuESbxG7CJTLAwf6tsg54OREMuNVHFNP0QXJMWcDQ9HK1HcMHi3We8zNXP9Hz6z0GVT+xE
eHrs1rQDL5dOl0Penek4ntWJ5DAqwD+2YbStnaUv2itqRFmhxCXpOBWlq8NQ5NqcpNa9dNE7112C
3nsd/2E0nkFt/LTRb8M5j+vTqOZbZggi5XVPO+saRjArB5mijCPwN3OU34FlWfekU0XdQrupeMZf
w/8qRFKZIsBJB9ccZ4gT+jREu8nFWDa4fSK6U+QNs6SZQJszqzQiOwb4+Zcx6cuxIsJl43pIttB0
Nuy3rFeOlM+fGLCaRsgqrTwhatiJRQ+6e9Uqn38FAtxk5eNTxTsbuLKDS9DtkPjyAb1Szm1aD/6u
fAlj6JeA1z5Tx0simfLqpFvb8C53ebWp/Kaixi9Se0CtI71t5lWmlRSKyB3xeNcUR/TMwd/1OmyK
AGZpBmgepS2aO24REDU0egXijlfFIkXlht4HRYqFdEqHl4bIVnewWuGbm8h71oPJdwq45EgZweOw
gBazr6DTXVdggeioeGwbz70p5klwCB1zhuixBGKqApORQtfNkIHsO65rBfQ6zWjiaFr/ko6R5b35
j6+C+ab34ZH3fOXLDhUeLhmgrVgBgf1naroJ1E6zQsiNJq+5k2UooB8WMR6ixt4oiUvzYPvJ3W6M
heoKlb3opBqbklv0cilSC4mx4A4O90RrFzNf+b8q0+YlH3ddkxAo/BZ6epesAseHtdjiC1NA2h/S
bF94wTufPR3ZruAodBcggR888NrM5XqQIL9t3BX7MeNUxEPY0TfbsmFVXL82T1zcGsIj6VEJGPwE
sR92THAzv+ktH8h2ueTXylziuj8rYIQlORKLBvjnsSQ+KXIbm7RwteeXPPaoaNZGSJG+C+biDzJl
YPAbdurFqCg0DgTFPXwHDu7fr8qkBOtFo4h4Ta10wsNmmz5Sv1jFcYTYFwaCfzOLNI98rtJlJdiF
Hv6yje2w2nDMCVGgXR640tqfmUzgqKHBAhqBs6z6TT09ds29t4ge33BFmRn3xWTGZsCR3/z7Xffj
JV0sm9+IDXIoZEh+c0wiSjbBVRfb5ojb0M+rMt/sgNYiboNQM6dLoTzddZ9+lsFBgtm/xXjicfjx
jkzljfRoWfoRzGOE3n8FNHoQwXlCuHzfD8GaLWCa78rEBp1SStXyPZth5VtQ2uImPjFbJOOluDGk
Qk1ygLHUn2FRaiJqQo5YvLVRDP3X8mcx0NfEII5/PgpLQWF2IKWwMsOAwyEZhCWIGAMtx9bu9LC/
iDoo3RkcJoJda4s3gvS+xq52nbEs4JN8bXuloZOLOdvrwxjByGizQ9AsnPPrWuKF5m0jfgVAEHTO
e094VAzyr+SFgbS9C0Djrx+km6UcR07/LwfT8428dS8mI4aSUIQKICza2Bvg6uNeTG54bF3OrHof
pIqgT3A7Sa0KibVK8Cn8XLLiUHfzLx/S2CDJJuE8B//ESFyNonplr6ZAbx+sF89UcWh72j5BqOCe
U9LkICiK/gqhJ7vor21ACS5fNtQX2Qf2aZH4FeUbTZiRDspGVq3XmDJHM8JkTO5htOM8Zd+k7gzz
uZJV8HrrvYjSTcwLb+tlpxEQ/XdS14LLYDKh1AOJ1nZtErwHdzB+Xqj9QyMHAo6mIww2lT7wE6xl
Joebf93/xEac0111vVYvLMqO+WCB1Vd2OY3hdsxHuqqlH5FSVduJrWrOZqnN5vAXgIVttQBLWMAC
9+okIZ2JqDOqveh0oKqtiFaqciGTrTq7+IsHg04M2Dtk+XddHEgue/AqtUtEEQfkI9HbwdfEkSEy
+/KQDu/w9YW8VgSfGWyikxPigbgaW6ejkcbZ7y4fX2yRn0QAbZBczAbQuKOK/y3Unx1y+/3zXn/M
63FQYj1XEsrZh40VXaVGu8EnpwGJZ1klPEG9wy824KL0Xse8WpLJYLSrdq4pnHV9iilmGT4/A4hq
fV/ckjbZ1rVr/LfimnseP0FazjGLIoUQQF5JC/tvDOIKt6CIIut9K4eQcRAHbAgYl39h2SL6LhqO
EzvZS5CdrJEQMGgOYhMrEe/qJQVTUG3CwwKfZDaPoN3/03Hl3Oxb+C9jc7ZukycyLcZDVzkA9MUZ
AE5NO3QdfIGLZWDz/Bcc9F4BcWM45Y5OFCKQpnw5oQw+QUkFQYaZ2rKOtZardN/1Fw+AJOJHdsv0
mOMJYYxN6IOOlKSa6hDxwlSlF5miTndqB5xg90v0sNVMAGC3yUvp02L03Zf6SrNPj3OupRK7RZWG
6k9EEs02DrUKY0sO5zc8pyrUI8Al1BG8MCky9Tt4dPri0fDtdM4lE7jjn0vSIHMZCEOmYdltZvyP
SXuXfMsr9zOZ80VI4J2WBHqJdMs8mUseFL0WUM6rwgyv7yftqceJrTm7ogrwvOhkER1/lOFopYZt
4L9UbnYVegogSvuyog4bBnZGU3hDjL6SuRFeDJZsELzjRwzoEANCPn5NhepfaqnM984p3Wuj4s5H
1HrnOtpqDD8PhRYa2RTPj5btpG50zZGR7YvDgWxAMnzGE6hy7XOUYloSjcTOxOTSIpHcorQvgs2w
TmBSiNnVhVbYC4R9/Hciqohm+9yNJvnzxFU2MNI9A+vS0wEhPyFlUQy4rYOjyDj+o1nA/FO16oO8
cZA2BBfbzhQIuyKMEuicT9b708UuQ5KbR9XS61DUlbmmuocZRVMWS3Hv90XhUGt23b+saM5EzW0K
4Gvs+VxAufHghGMu5UpgMzr8cYEPbn3IGNoYRxPay4CPglyc5t7k+GPRTATzTzTCv74HQdHwexjs
Qj8vb5e7EKBs5UswLWJHqo1Vga5bY4yAoECrp4Rvx3/MKlwo6qeCdDZK5nymuTlV1KBbGFYlfjR4
7kfzrkY19lVkpweMMcclbab+SdV8fFdCSwrc95bQZbuI6Pg+/RUWq+kWtufVqh/F2WfU+KxgHk5b
zjee6YGsDGe0ZPrKCL6xZoOLjMnP9jCNIvsU+hM1DIKGk7vGXfXbNyQ5axlqnIL+/5fvcUf/Fi00
uRMbcGyqn2d5CZkQa8WBfJJuurR+BsLjc8pRgjq2L1SjqgagMDGm4tTWpqoHwZPjKF6VQE8+Oem4
Zd3KTLAYxXy2mycZzyJH2vBWWbP6gX05Vc5vGR/OpTV0A8xHmqdIoDQZMTGUTaNtwEFJz6qidxZw
aF4x1hf+GJCsYcvpn1LWy8eORz9t3mdVeihwaIsOIOUJduyt1tTvHQDEc3Ar9xtUT8J/Lp6im1xC
eE14TjJoxSs1olT+AnK0URUdd0OAsGFmxpg9pZ62tGbCZBEhkU8dXAabx7PGGfz/LH2nWrC3xDhU
PJ8n7+zNDKNYzm8K97iERHEO57WpDpi03a+JYs/6KLTGBFQ4d9JlB+fDkiaVu/3rmpWtVNeJ76zW
eVdM9zZvuzTuXs25HXXA/tjLehW8OgELXX7cUXjOPzJLOcOtwtuDqZWzyEyY/Yy6TYEx/0rK7S/1
1ecqYC4EyZdHxcujZNiRwpKwl7+o1/OOW3RlF8GtUXV3rzOM3lDZtrhy+w2XZwnoNo9nUU+w1Wa0
l6cI+xRe97OvTWsxuhPYCoKWdwq1QvzZfo7+Ebb0yv14xi0nmv+lZBRpJr8JWMEEpVf3XTZGgEqc
s8n/lemI7fgJsUPMfrF9OOPAnLHVj5A3YOi8s0Fh6JlORlmFFRcpmiMu283hyJVWriRr9gcJE4zp
dsXDjfGPErlk1nSg3RgolSxiYTd8aGuK7ETjvkLFZC/pZbjsQnZ0++egJKdkxCZImp8iu+HwrtLU
bH02kS5X6Ej/NjOjd2K7hNQ/VFnEdosxu7XlCt8TPwaG0eZZOwxk2JLqzOv3GN8+tujCB4uOa3Bh
BZ6Fh1rbl7q22n8jdeQr++s+TrLK5DlHevbHOpQVdIDukb5h9KXNRiFFUA2kIgg9fqonXM/kKsdd
ETcAEYdor8v9Wo83vqVHeFeIVX5lViFAQbFmocjOEmKcYLxik2paWT6tWJd9FkkWhZPP5wtF+thf
L87ZHq0Ikc9WNWocvRfRALm+6WWAaRrWHZQsWUNAfg7hHTH6/smBhd2F2FAEnKUkXCORpbX0QWyB
9yR93qUO3dDRQ7dA4aHCwoqWzGIfQvLgtW0mvRYhWzYyUeO2fHER8+y0ydhasTYv8bMQCf+3zj5y
8svrbFrHB8h7e3RvttZLCasuBnBUplCS1ABYhMd4GCuq7DNZBLW1jTzmhQjWD4TQNWnMAYz4e3At
0YySwoKgGECfMF0S6/+7E7UtLJE2gO2iFb7GgP0oc+iWo6mOxckwiaL/Bp32RcDB2uoM7qWsnf7u
aQUsnWr6TMMInhxGPyVhFwnAN7fd0MId7SkDn5JM4AyqA+As0ZbnvyvwNpeVLZpXVipHMTioafZD
QeGOWHEzE3VyrKWJ01zWtdZE854NH0uajy+bL9rIuKlWeNwvmYcKi6uIvGkZBpyDSxBx56JMAX4h
RLzUcwSPALmNZwqQvfpR7KlO5ewt9QYAciu3tZHelM/58moKSb37kkYO3sacIosYP2TBOsk+ewEd
yj+/+ikgYLyxMdbPOX27JWr7qRzrc72d7EQmga5x8cQ6REQZGjXkncf2J6Q3zH7A0juuA5iOmhMR
RGW3ipuR9DFqLDJO2rMVsryXE8XECzHxuEdzt8vKfDQfGnvYlB0d8ugZbGKDWyIT+6V5P47hyy/z
U62HWa9v8iwRV6IDP0U/LRU2xXI6qvDxN/tkQ4qVyFDgP06ZslHTUjmtzrKfSfBoMqVJ05LZDe3Y
nXOoREymLIZISUCP2pWSrA2QuyeQaR+6FmDpvdqpjnaMRkpzoNjE63B7u6hi1aj3OTe+0bRuNHiO
rIGCk+g9m6JORuKTHzm1sUbkmPLJp8Ms27m2S0BWbcq0ro61TrA+ky2NgcgsZuuxXTnI9SnNp7oM
YC7RREhd8Pi9S0ZL+k3M0aHIJNio0PJgnxMMoqYaYlHA63DU7lxQ6N9aCx1ejGK9RNa5BXcxVFvH
BSPyHJrPUM/rkz4JAzu18LTYG5CLfW6/Vs9Zl2tZVqKzDwOIGqNCQN5+aO/kgocIun6PmN9N6mfC
SgL00JxFzMiQQ6Kql4QEWTHJXbi04sL3IHb64W/7Mwlg2bVH5GDcqmjyG+JBqo76/LPpiPbPtws0
PGKDnVs/3nxDZNvRdLjwb9ofU4y23XlTpo0sIsvDbnQ2Ex9QPOAHtRY6kli6vnHWO6/PtZvCZHZi
Qa+24ykeoxBju3sGYlMAOjXS9P0+Z4r5BxRsg2tgKsKvgWFEgil0BDO0duLW9cR7HH73Gs+cUC+V
jt7M3ZcTyWSLozniglsWumUjrhcYf9nqhC1Q1N0e6DzqJaDl2kg/oLQKLxPRPadMmqMkx2Zy4hIw
rf/7q6zqtxOnblXgfeFDD+J2Wn1GRWFzT+IgsjLWbYrWWvMZeQXjbiKuLYKRc5ak5V3/uGX0yFdq
4bSi6sZbbJk1gvDsO20QPNilXFVnouZ1aAKqvROv80iietYiWLVFp8iyKLuj4D81eoloWbj05Vwh
UMLH/nyhRdQm9vnIR1kIGQmllt6RCvZ4aRL1ewMBCCgrgBYFpP7CzoTjfOm8cpqiIWj07v8SGrX5
iLr8lbz2/3G0Sce2qfVVDl2f1Q+bh+fQ7FNcZ3VD/yDnO5rBOPkb2O72uG21iZupo3hLnWS2NowS
CkETjmWLYhRsxC0MY3g/0SN5ZUzzkQTMt8zkG8vJ1DILpeYS5zwuALvunTj4SSoMGncFwer/ASEk
0nq5OaisaBm/DN+INEzeqpuvL7u+W/bwg63XYHjleREN4XhsDdukcl4qeEa8FXRIkIxdCpnv052A
x/XfA++uh6uRBxS8AKQdJu65Ftp416gth2RHAFXUEcPLzJwSKzHRYXAkjxxUf/hsCKIMrFMj9WOg
NgxpcXa1e3ct1vqHvXT6al4nR4CHqN3h4cjr1Jqz031Xcp3jYaz/6GhOZhPPBDEhLt2h7gFJFRbU
iZFP6DxaBIHXH51O+p4QsQH/HjJKYql4mW1AP5NlcnvndymVlh47PI9iYIfAcI3s/gaJO9+h5DYN
hMB/nrJGaM/3oJSZZ5AhWvzMH1TFNKJODHJhO6jZb4KLLHPJ1Vrgzzrm2wau7Ca4gQv91q/1qKeD
8xOtEXfdnqq+fkYLLkbRcUO8Qy8gojylbXHX/dHIOTBisFDKiDOPhWWKYQHFpUjPMUhpHm5X3BeN
BSk+2P2YTxShAOibpuc6f4NGEEYhOkjIUHKvbnUrf6YKSXuMMqGyiWqo2RhGkUbYn8yboXeSLz28
oz4FfePn4MICg0Vl4L2W1J1VAasPlSM9EjJ2NJSp2iaYKwp67FkJ9YEIggtmj0hYF9omTl2huyaC
z6ebVyDADyFhvaAhoSXko5UH5Dqo84Rvd5+OvZAVmaLiTd4H5PFhoIPuB+pr2uBuh0lzFx7puHkT
oKPwH7afS9ICihqbvY/LKvA9EPgAoq76igupy4dgmXnmyqznouweCpBLi/WuCNIqG+J0HYaEWbfp
gt1tRbgDR69hQ4kIUyVm+Bt/O0Q7wVWPdpBO5HmT5dr3N+b1ytoPt+aOv8kqxN0xJomxSJLfpchu
MoYnUQgCOuWBm8X7Ggi5ILkT5vXjaaup4EEhfuGJS2h1bv4M5Fs0bbKamddHu0vOYk2jb+qKCOnl
8heoMXJW5nZz0NM2uz/Ulcl3qlkb0lcpRJRHGN1/LX6TL8q2se9Tp9YEqxCevmFLRPile4AcqrDQ
iThgd8Lhcc3BqQ+fAssWzdksWKvANiiJmlpIL/OgAIMiazqbo7viN/F/rC2hNDnJOeKx+F6B4nCH
Loa+1TH5lXpi3Ii39LhY42cI/Gik4d2wM/Vxchd7J8RwWQbi3DAVjHMySLn2WK4jUIBkKXipcVPK
pKCJ3EQ2TI1ZUKWQ53GTlU69fPt5zUpQv+K2NDJVegcsLePsPtFF5ml9uo03M38JSDuh93zDm4D2
bRjmB0kfQ1T36Iyi0g9iTgmFr3UnzEgzrFqAwiW7DT9pvsX98YY9sKamc8Ue/fmXj31NrND5UQpO
U4mzOWrsLaZgNZhG9o/oVHcgC33/7IKGaV3xy3nq7y2cevE0ZDeNovNraMMcnfd4xwYOmvmjwGpr
Wj3kuXDZP7h8OuS7FLpbZK6HLhbNETv74KiAPUQC3Zd6ccPVpg+oxrjadlZ/C9o5n14qv37Ay0oe
jP7leNOEXZf0neBWoOn6Nlmd536i65pZs4/7ORONlU7Yoa5u7rtca6CpUenzPblM7cWaokiafNtC
eAPQQXVh2N9CmK+k652JBsmolJEbSbwqdjCLoa+wHtol0WmeQUMLRwTG0uEAfzFlKCo4/RgOJXP/
GNZwptK7a6lv3PP/ORZlWQ3Ha1CefwTRcUKR1k8j9nUKEKY2+kYRSOup8oMQAZ8asYKn6l/qF4av
RrWtnaPjmOIuwt3nv+7q0zYXp5PjsT7kkkpR7O1rRXUR0d8sywB3qs9zLmRRElqY4MOPAQgoZ0iy
6y+OUHvwzYqIDzYdhy0lKkve8ZOiT74yidcO+yBKjruqmDY/c16zhSI1vJUYd7IYgCdSqufcMN3f
3jzpDjiJELRRm/ivFdaBmg95Z3pXab71f9dx/L8m1RcqLBiOGmQg9BBUAwho6p4dO2pYyiiWrmfM
c87+csroNZyEMjCvh/7eFjW2Eovk/7dvldc+egZ8ihRzos4sD5IRqm5YQkkYhSO0mG4qOpYG7ohD
qempduHpFibjOhRSs1wMKn+r/6JGQJK2aXltefzonWerInLkMcvg2KfUGqZGNxoyTLIi9eLICun5
LDR61gvY091xo+dDtjKyjQf7uyfhiLMu0AER3Ikjc4pi4GgdVwtADM5KR3G6jdh6ksMzO5J4aBH9
HIzM75wELN9JvOBR1Qc6izE/81d8cRLd5MBS5EfeIxP4zK1+N24SzfeNqMxpPuCnP/ez+jH+6GdQ
/8cuhlrIOmXbDA2VGbjjuRduOfBGZGIIiKNwpTAVMnyXliL9vZ8iqJMOwSMAwM/hDkfL5FhqvYFo
xfD/YkYtJQuZvVzv7vWWSRM0rJPstkujoRtyf1MxASoZ/Nphxpps67q9xEfKQD80BL7OPisJAaHf
QbKroYS+oPzQX7ggDlvLPyOH/kJyIz9Bn1VzeG99JCVVCb5sOGcWSavMqv8PWjd9/LYIJmUZ2rJH
8LYfStiCbZ0RMbShw9onSuGxqRqkcZ8gVE66yk8oHsCkCuyb3wiV0G0a1oD3su4jsGlq8U82VzSm
7LdzPOeAXkICTADJjKA+UBiyrG1HTwne8zv36omdxMbnB8GSirAGdqG5HLNA4fUbZSyjjKO1mUmO
MQMdN2klvMdI5n2sSfQ8OimRglVuZYgoC2Gl1sj1nxVMRJbc/AgufEsEcgeazW1YRhitqpbxnyCx
g4ROfnmnYNrJ0TBYxKWS1POQi+qoXR3F3/BwdPvSC2Xa0wfvY5qoMvsFG+0aUJYpt+b2XokOcy8U
FhQAvRj1lF4e0Osg73vQ6aBEGbNTxiYvL6SuGdahrAxEmZjoN7DVwFfxt0XZXSmcMSDmpX07cK68
YC46ZqySpi+W9KUym17qEQ6gauOla86JGxoHtvpd3wlr/bJhsgwXGbhZ2A1NDmVslGiGVOKPXTJg
ckYge3LVbCLFKxWm8mtJRsJFcYUIabkm2KeQhV5gBpPlTm8LN+Usat4LbpQQxs4+0HHBQKbESHny
5vJqOoMC2OiWIxXAbt4qc67BOC5iOF2pzDXZDW7NhBrrhmxsehKh/HKyrILe5jFUgFQ+lOcHo/gG
yn6TLMzKiLLE6FRqrYlHZxytXF9BZPgciCCXPKX+T/Tl1N4Slnqfi21RgRdsO7lHuakHmknmbzAY
TDBPZ0jziKMUXiqbyBNZVhWZqwIMadt3i0XWhWw4EHwLqYslZzPLgG9v4Z/fMxt+N8jMQyuI1hI1
9OE9mjIezPIE0nsulIO8pN8KFhgevhlsmUpzcfG7xj1Hjx+HUjYfn4h2S5RUSwjh94vDSkdXKZHa
OqwaQ2/YtqcLjaoLsAR9SFr8zXOagHEIIYeOqLYxI5k0BrQQtESW44gfhEjdUQ7Qhm2Mfj7bFF4w
O0DGp/2P8/gOuhXMw7lBorGIvqGeb9bo2wbw9bcKQ3j/7HZw7MIlMGCnjDMznAC9zHlMpqU1OzBI
EQt5kRYhYjEiQ2O9T3TjZiep7EBgcJSmon4iDckCqpwe+kgyqFpRk5cB3tWxYYGwCOPbfm4exYgd
sdGCGolc3NlLyCz8wo3XRSNFW/qx38FFOOAZ/cC+/trkdCJmXIADkuYRyhuSNv8ooa4TBpIMw00c
aQUCZ9B49uP3Aw6mi0XfS3aMrmegf7D3VR7cm1YUGuut8uXZyv5vxFGN3RfyMx9+KHAyebZcy7ba
hsjXh7sHAsb4bIm3bF2xelDj6hzdGL50emOJBYZzavjZVQ4C55e7RlbRRyau3qTGoLcZFlrHNta/
nORDLHhWeiPPdnymtvi1XFtqXhvGQhZYnFnpUvIVvhDhxdzx40scDOMH6kwxAZMc1gxgJ9JcBc8R
heKNYlrFaWvZe1TM6RihgQB30UCKxk3XG6RFddGKt57HEmHczNZxAHpWgoIJVnkWxkCN6izpQnLA
kOElqbDWhHounGVbkr3+HND4YTV9ezeqyfdgW8MSJJUKb3g2laqcW1MPS8X7ylw7VrO9lhnu33Iv
KeZTGi7eoEup65NaKHmZ2ZK5WivSzc00HQfav4VYorQVbJC5fCzQCNWckDMpu53hQix2SZlmiuxG
9mxQ+F8/92dqeccbVLvjn3NfimtjQO3aatd4ZRoGzlbCxt8qCQi5TlBDvIc5xbNe4Ov8wEJ63Upm
z7teuHubuLN9RjvcPkJ2XEGcQNWNqo1RNoUqcIEFIQ9Ft8etHTNmodWPqRHiwolstmrhqn10WqFN
ahZsbk3aawEcjMbe7gAiKRWSGpsj5EEoAuUfOp9qDm7neZdUUl2aDU/jUVpd7o+Z518FFWuYxLxc
DUGYWBqcxzt6pMcFAcoIpRiY+HeHoVraLHDOMBv/yW4zP7TBEUOA3YHrVbKfMOAMGW7kFNOsu2/y
Ogho/w6r5r760Ys8FHKZC92wx7sbRNWys0vGjy3x9774jTjMrviMklIbeytCLZqUMC3vc4w1Zh1X
3RoZjQz3xCMg7ZW3ht9zZQ+cQVsC+hdKBf6PH5UUVbHY1AACPZ2Eid1KhwwzJ1iudJhUl8tf+1ic
U3GUMpgPeTGtmj+aDNR9GTo+45h9vpVIOW6+zPOz+ot5B8GAKyjjMeStcf3cAfpqsDSa7EVYUccD
y5Ksapt44D4r/HfpmfBs+YMfKisUpNi0RQTycE7vrWCYLfJKO+M6/gC8FO5DHOn4GROpdeabjfSv
YBGdFM0hooACAqGJVdlEq+u27S8egLvaHSGhsO1z/X57XdIqYSgTFZqpX6btKjjNABiZGJquPDut
IWj7TW623ISeftjSbvoK00NwOI4zTXeqGKjJS9+gZWrtgvvwMAmier6w2Fse0pk5WEQ81TEbp1af
X2guoSMWGD8yWeCsPSdf38XF7ncTr3WKyvvxieH8tH0RteIxiIzI3nubi0Hhc0PkGen1NwpiA50i
VCbARf+NaTdTpB+cYyobUEZ3/vj1TZl1xTa8UsJDNHrMgBU4D/hjR2l2FtBEyUir7JrO+pkrcjUG
Bfx6KKgKtv2v7uvesl27hMjNFLdAnOweXnhHx3keQzVraAt9b7d8mXXj35FVKzvTffjiyu1YDzHu
dr6YtSKPsNrUVAK/OPENRas30z0vYfm8TTFFR3bou/cs3tYCaPc5KkhPScSOASnf1BelRb7UMLgq
qDLEtHVCYNEh4HSfA/YFuOBVsZ0t26xm1pf81KQntL0L4j4ylqjxypZtyV8FwIzmLi/v0Bo/WvLY
QUp1s8hv1eMEedilbkynE8T/8kVDTvLPxzgRd3rU6m9xZQN/VK1fErKtTUCK6yrJvQl9qRVrlumk
ZU1OMWl3NuVq+CIWWv7uc9qbRNhFk0nfi5Lw4p73996jc98zNaNlZTEQj+o/SiAkZgQCT+gpbXqJ
pLg4iQC85f7KGe7eTJNvVH8QcY6Mf8hunZM2UHr2iNMr/bNMhzEc/MclzGizGdYz+jtkT0oH5aO2
2uPgPKyF08h9HoDytg9BppKXJDcuvJLAAZpP7FqFDIL1UST8JdH/L22YHU/gNYen0n2Au8RdI4K/
7a29yb3GL5KYVgtp4cm+HrXS2NwLR4K2cY0er5WWjUdi0UYTeVpxkNYtTb0vqzAccNMJgDSTuktx
L0rOg/2kyhKpGVd4liw/9IjG4EGZ7qkMb6Z1oQItxk1ZPxH0gp+W252RkIBRiZWyt2DZmVIPaR79
fQtjBcl8KqN6M8baFA5WC9QPMcGW+wyV5Zt0Qt0MbkCJT5of8cLdRc3zvtUlcggwvsDGaRRzZhWq
4/aFqHh+1DR6BsVaFYzLn9YSTwXLtXA0yrVDOZKJ0KWM5eK0B2qOzP/RLIiLxC6P+X46BXRml+9+
JH9TDclsrbWJGHc9TEI5FdGK5dMclRaLFoqA825jxv69T7lYLOsUZHmj0I7w6tUgVzSJjdCxdJ8o
ipXQthYZ3EDQ7kGJoU7Ey8BHe+wdpKDgMVbBeS0uKdcGwyxRrcX3yaz7nbnkUon5pe5srRkZOt12
5tzyk6cFGjgeVygOkQ3SMOdA3Q69Jfn31IMdnE5sLWL/3aLirecnGVphb/r0gDPqtv1q5B359Xr2
kmPOFikDQuXRCM4LAmQ1RmmjopcvjYXMfgerQkNIipzfhzfa+vZ44H2uSSOYqXEUcEPEzmTt12qw
0Lz/VCyzWohmNgOQzqCcSF8uiPY9M+5ufcyDjgZwJEOxsxy4ypOQNJlTl1MTi2qYzKVKqwPPOTJi
brvwD+JuUlv5KGP2iW00OIOxxRzTlakoK/XdV+vSDPWsIkE3qRtz9HCnw9CPGRg7iTS8pNQEE+Lo
oyfm5H228MFD9t5tJvNKYrEmlFapMqiMy5qsFlyLg8RprE4hv26P2AxK4qD/LnlHYEU/8WAV2aPn
VBX8qFtjdpuDJ0YEuIMFN50LBVxyrnRg5DZTiIEaQIdnHXM+MTFDs6y4jmxMhNO92DagAsPg8vzi
GvujBWDYCg7C2bawYi1zu2brhihtM1jDJtYa7Ocs7EpRkpR1VYJAZeXW7YlBK+iSpZX8Pi2yk09x
ED7CUBK6Ou8hVBXSS4hdJDctDnkTOj4ZC9fHf55TI6WoxsmZJ1w+1X6nMVYBAO83v+5v2LNzl7f6
i5/mhqv2RbVKA/EEMD7hRFmkNj8XgJYkPDWu2p8oMNZs2OnwTPkqGIrje/TYnvqvKgpfEedh9GVf
EcDHQq8h/ZEMzfoXVdchFiyfiKplefhYfmNM/r5RDsGp2JqvsPILy+3LZ2j03D83fDpOyuwhrUmk
XR+RmKWW5dqpknHeWXjtGIRyFG9Eluvo4WCxxyT98hJfdolzIrnMLpi5tkR3hPXqQzwyCl3zFkEf
ZKNdzcPIliDApiQFUZ+nuNQDby77sXkT9L8oGC14fTIkVMJ94YCtJGdl63rQfR/Kr6gCM+Nvra1d
cvRdWF+uE2t6ghdNiXyKwa5NIr0Imgehp9p6AocA3YFZ2hiMRasnZ6qqQUKMsk8LT1t2P4FxZYmK
IFgiu2YZN4KmkQ8jGJqLj7viIZoBL4uDRMiV21Pn1TUKGh3HDdilEsc3pxZ3Rn+wSFnVCs+oD02/
nw/S8WcM5BctkMWENnYroBULczH7zhGd9morORLlhBft+DULZAHGMiu+uYCkvkvyWjATM25JS7M4
IGpllwY32jYd0F+DDida9k+cd9RfFuG0H73DDBJxX6WFivbzn2kE3G+Ve30Z9583Gcki165BJ5Km
VPi5PvQT3VlK789r6/4DDaWRkmANgaPeGezkc0dKZRlYvW+6lST2Z9WafIPNrpkX900cobhjK7nI
lF1kJjz143SBuflHNbLHl0+3egxX1iI6rwMzNRzkOzQ0GJN1TUzxd74NgJP+SNiP1v4XxOLGSJJM
0lJOyLvc5iJKmnv9i+LfnNFUQQ9NZmy3jb5X2Q53dGOH1Edpmwinf6S5I++nxrr9HwF14obnIANL
66aayauSGVfHKjzn2PyxgAtxh7d9sr+C4XoYxIqZwjUAfHI78Z+D6pDwMLi3rSjhw9OhC/sQK5TS
dBejm+P6A59zpnSeNsTvCk2I2Lpj5XCVxXyFRiTuU0moieWd9310RFp/nzjkJHf0SUslIm6GrM7T
3tKzCFRtZtsBZ2H2UUM1Youi16uMiYyR8k3FYkxbh7Ho7JXHK+PSHdhN8u2PGz2TijOjl89IKemJ
u8nDZ/2pUP1e0DaCozBAjXDkEbc/a6p1Tcy5JSyWHkl94TeweyK52ZMflWviSjgxS8FyraL3Qny8
yLSyeXVJ2NOrdF0AeW7Ppg3Jr3dNiF7m/yueSqA7f2XDsQsnjl4b/dJNJ2HpFoq7cLD7N2g2i6TL
AzedZ1cddHR6lPlE/EhgAN42maz8Gp30pLVG97rad76vEBUDoy6SkK/1EG+c4x3tNV7kHxLGygEp
5STHo0c6qq7XOUeTtbjgNtePl9+s8ehkIyHp6B1iO6noXhj/9a6l2RlqCeGzSLs5zZkZU2nvWCbX
QMyR9IXaKiXQ/X99cDWxmxjGGZ9L/ju8vhvmemhY4nbqtCUebRWciMG2KPmK6zXofdFzoGsAJvmf
iirPkaYUvQGxAvL7iX2HlUhz/cQ0UvMJhgVNDgjGPq3bD0k78XI/0YPb4z6yf1ZXAO8QQqDgVKoP
/hDaWs/l6PElphvcJuyH8Z5/86iQgcJfG3IRDRK8bHyKgLn7Qjro/XVPVLj6dHZFGB69M2qVeOIz
dAPta3GJwf6mpHCKIQfHCKJqLCcfdmOaK2QIpg8bZpbz1cNsI/XtZuOeXJU03jBhbQRFEMl+gmjV
rlfCPv+csPmusj5NPS+thhFLFYELJToA0j/4cjIXpYHZQyjHFtehh0MMz1fywuTT1wHM655xHM2W
IozQIUBi+13yT2+MLYR5MNDvskGI3jNh+XFcDHqESI0XgP6SICqUIoPUPGVjJ40SOwzMrU3XJlNf
saLK/x59o6xxzoCmGHmMEDPdOQ5m4/eUK4x15aeBnT4hvNuE6pmJQ6lzaXmfCZHX3QXxJD9m5X/o
c16rWej+JEoog3PzAoGSbrYlqa7j3IQvG6PKpZZqfy2jQCZu7tB26jCyByWNWKhGuhzMOixfrfUN
GYwdhBTYE77Qgkl5iORtNflD1bca6qskJCs+fkUAgiNWQxutjRpyAYTNNhH7UQqpcfCI8iWqLptd
porHW5HkC1V1M+C3Gc/de1uDnUj8sg9WA0AJnywPgeNFi+oMSysjbLnVn0yXw8k1d4RVwTqHX3RC
ID/A5WFYJqSD+x/PzrY1jyiczOuMu248Uu+YAqI0BDjCTTLmwPjTdNvuNW8MOUJAQdT4HMSYgf5S
DkkqM51JNgZonpwmspjVmZfKViZl30at/FoEdxBll1szLX+5StiWmg0T5KfeDT22ii/E06OhNM/s
asXQr1kmP8okkGwEJ9433IIIxWSFFjAG5Be7sAADZw9Qd7lLnML+JSWgMFhsOzrk0ovT/ROX2pzE
5RO7TWjBH5gMvkpqUIC0IuQdCkn6DKMaMDNm4ya1Wql+RTf/gvV5b1e4f+h0XT4ZE1ySDTZum+nw
UMjBT2qaqviO4W9bJNp6XfqaO9Q6vtvzfnvGnURTAI33VYHwI+KD/dBMKms8sW7M24QoPW6ur9yV
bfQqw/eA/3Yf5hsIm8jA+BcjZ2Ait8SD41G+tkX7wBlHAkQ351wY1ICEWn7m1MHxmuJN+Clrq2Ne
cc+Su4etcZAyn9F7JQzDSm/cJ8nWyN9bP2vTBhxx4wBn45JokCTPuERGpNlTORgpEQISK65/v1+e
6tzpBg5RF08S2vQcFNu/phhfUQBhZhcMzG2SZUW0MGmhpedLpRXZM5Shn5uf0KhMKzrBfhAZcD85
B5tCRFHx9MvpI0UplaauFeToWQTWFKrC+VzsoW26szuZWrY8jek90hinZWTagtGwpSOTeAkMR73f
FkatHT4kDf/Etqtyy+cnDrRKtkPmWP+AO868m5SLS/e+dwvZjDIPJZyzROCROul1J8hH67s/9bk+
5Js22wNeNSxhMaUEQw9fguysPGPd9FNA8cczc3ETk9SU2oj4/YWQYvvURpYbx38nixCHg7MZnBw6
5ZIdNfPU83ELSg8Yk+gL2WjXmkGSB24UAyJ8VtTV+4p8QbUAchN+JpeyTXPlydx0RqXP7WwoFL/d
YZa4aUcSdFPLtyUTjVIJ5icYut+/7TUxYKqEbYDLsnFjgeOfAOhNZlsq8Nu7ZQOpbDBVGL6MkOZk
TcmFl3NVPIdLzx/J+RZ4LmngqtzXlyJWwCK2MEM8OtovqpJty+cXcUTo8CjJ8M+W6nBJPQ4R/PsU
Xwb7K4cqSK12E88qMRgDra64cn0l9uCVuylab+wd3AvdFbyDJeLDR/KTEOv1eUvfbjuHyfgrR8lB
sW1FGsa9qvRj0pjwIt85vvPJGkakjKkdETrkNQR1VLvwo1nzuzmsQqLxMNySPjhpfAH//UyVSs9W
4ToRtgSCecP1kGUMT7vOsC4wa4AL1Yye46yWIf1rN0tQJxm82fUhUPnkCQM3qzrRsP3GGndS9WKL
A0CErsZQCPnM93nddmUZyHnRi1iuxVPCxrAV1zx2nnunJZgBlNPf1W8wyCHoeFaNMIYFOhZfBWUB
jcpjxttjaCUpnFAzZsaVKtnwr4EtA+rcbr6DYcwAv0bD+k0Wa30HsOQLbDMG9BQW3XLFwPl3DDJ8
khdi4dSochT7zUi7HKsfyTN1gSUr36nR2zHRmPIWrVFL8EXlObmymkI5V4OtvfJP2r9iV/yVZ3Wv
AD6ldIUdpAtPf34fR4fgg3UkXTJ/2/FiXLpPePdCkGzz7V+nh0KMSsGHmUZ4exaLoKiPbhpTPkDl
ziFb0K4OUtx5H2qUKMeN97Mg14QFbs9lLGQOFK0rEPPVhhcmit0OiFaqV5FQ1Htmg2OIj/D+hc5T
SBu88yqhKb1coAY28pktVZWl62sEcxVoC7B7zkUSialkC2iSvBGd30TwwasIDYv1s+5o6AK2/NLe
tXxCPYFFL8EXhBrVV8A+QJcxSzYdrH4iC/aKkTtfmXKlcaqPfD6pcu9TMbaJIQ1oSWL4Al6n/2Xd
xDdXvQQfdJoP60PFh2bNNynUmpMMv2ADeBklyrcVJ4h6dmRpoo+OZNDi4MmnSzx9937kvyQl77Gc
jJPFJ6SoaN/+pGV5tQC1Iw+/g9uwactcDST2PafQnOJi2t3tE9sgibrJv39mSa0e4R9ZJxyNpL8Z
ilI0Wk13Ky1jfePyK/hyxZvkOI4HnrQRvHZuX0/xYgBUs1+qyYl1pVuvcg5boz6jdmamQua2cBh1
pAsHbIICMTJcR8BZBsWFod/64p9P0VV6RZ7+ZNy1Bq1XTrn5c3aFydNX+IUcCiTz+Ne3C3TORbnc
PnSdcid68FpYlAphsz1Ugp+n89WtS/FWwo4e1PwroGc9M58dX9KnjyprH3h3mRN1UvdpipMNByae
aHFQe55SS6Pmn0zmxoJf8g2jfcfnGyzCldKgURwmBnhE7ot18qOe6jLP5Bj8N89QR7s/m68HYUKu
ozuJm7wDDSlr1VEODHhl3XPCCVgxuxZyFnR86wfeOr+uKTsLhpNHesCUrCXMK+dpZdsmG6R6o1ZY
oGVQX6If08dYNPuHajQ5PqKbf5x0XlFhlg+GMT550hnNcLD0y8Ru0CaFB7uVk9xD41bXDQPkXB32
LtVJdt91xa73OMOVoGecxdh3C7cKSfC9N/VsHr3SHuhvPkARfegmYqsCXifi6kZAWuBVn6xE6euw
T6bYX3wJIwjCiH6IDE5xKPG9IN5mCQ8YzxwiNFqAezKMHnu9gPe686UHE93Khm2QsJQzGY3oq1mJ
qQ6YUOlqHLgz+Tmn4qLp2hAyU8OCNR54z98W7Ppc0bB1qTA5yTEqJJHgk9jh8J+1o/FScQKfnZ3Z
ZnbdjIAE4SQLLCr2lCJxbF6EywkiWtEOd6YeO4xQa+7chmJiQDvmdt5qdHlymxWPcfwarYxWH3j/
wnPXxvlQr7mIjNIRKTjJ7JfUgnf+YVSRwQGM/LZ+Gcn7h0Pq3i/JNLFs4hC26Mj9Q1+q3pPKc10s
w8Hw6CUT7vbFVzBG2gpn4Ney1RW2/cNP13sr1gITwtlksojRl2BmjZIJrQL5lifQee2C0jZKtD8Z
hn+1mMeG9itEQcgrvgA/ALcVnPceLc1/SljKNUJz0OTIHoGdZ1iWk+c0n5aepIw/UcO8wL2pJtK1
8UL93Vj8BTJZ9BRUi+ZBxKraHhfwmlerN54xp/J4AQQFR08PRLyZ/xOv6l4m7GEuZHRt7f22CGC2
PJYMKB3uH78LiFSLgSaXrCnC2Agjxzx0vuwM8L1lClCLmqbmSnN4vn0EJpH9CdYUwtRcxBIf4+Pl
qRPRBQgxZVqjog4p8eSEr3MPfLMZCwIpJRgSucMTyDFD6vgrUzcU8vvhGI7KzqpwjLPQFqWczmo1
NKdF+TrG6dnWBAMG44BDGDyQDab0jTVOUjx3viIX8JqEFKnTVlofoYqybdQ+0qO1Bj6Flll5WYwq
gwntRwxaPwqkvyBlsON0A5b/VcB8ttg6y3opIFCzUekHK+IeBci6UdO8e5xygIDpjPRNUS2ZBqU3
jUnLdO7QkFJZojNuCswluu5KXo9jPndz1gbG4FmHGm3x8c3M8BcELs5i55lDsVy/D4dUb62cLKL4
u4P/WM9YrHROm9Zq/a1TYq084CTlmWjoz2ageB+J43FaN4LuhLcWnkkIO+eBGi9rklorSzXGKpCJ
se4MdyOfp2BSYHcysufHqaGGVFDKN0Ht2X0VPZB7Mp1/W5S5G/GaMQHpjby4tBU6YKujLsEQNGzz
Lro0MEK8IaM3+PXartxcAhf9lu/eOoL1TBjqoy9r4QDoWuZE04q2V7UYRPL5Rdkz+AxvCGFL/FNo
WT5L3N5X0xND2JxMw3RowX4KzjHrijwDHA2GDFkRxJeLRaVV27pLwnw5uRkgtZmijMfQubvhO0hR
wmpaEcPPyElDHSrwXfFZ1bYG/9HJ+tgILWgbKXRGKRhin+5byPk1aB4hC85lZ7+m+boijNry0tTy
dtvIY5Rltm5T58josTWmXdW90QulvIKznTOaprnaICMrX6wo+i6FK23SKTRsrXLd6XRC/5VDo0oX
Tx7l0Bx/lkUsB9dI/4yKTTUsjCiVp1OmKMVMXpcGt5mjTHrVeQUw1G6swWYK8txHfw43noeH+CTA
8K+SIQ5d91wmaprf1NYe17hw0hPMHEczdFTvxDaClBvSiXqZE2BYo9qvaQyVIyetZooXp8oASMFC
OJ8YhQ7G5aONYVf2ZZOW/1Oz+UuhiXOlgAdNT56Rz9CZ7aNOCqLBGV0d+h4almbpK6nFvKgmuY+h
ssrm/I5ghTSgkq/wKfGa1M1qWvobJ10no8RvJQBvMukpEkbMJXKdH7UT2xabHXr1kwYHVkjDCG2P
1xub3tJFQwpasDSSHfZvWU7Y5i1SexlhqQoTM1jkTkKBxCmM0tYoXiLgpmMa9lD/cG67GstlbKSs
llFwIxGsJatYniUV4yba3vr5goL/lxqp3ZF2fVVJIpstbTJKOq11A4Ka2gnlpZV3u68pD+cQgz3G
jwGY4+tTsActcFePEFvpBcs+j26hFyUplQaEsMjivXdO5+I92KwxBhBozZYYnTauvFn/v7nh0SnQ
Sj65D8nIC+/AA6OwvBRD4j6B732i5hMADFeYv1O/KxB39O2TJaxflNiRNSRHeyOg/d5gUJ6pwLzc
q8KNVS7oWHEhmn0qoiTDqmgrbuppVq9EJaU4a+I9RC8YK+OtdwUdYRY7mSbBToHwjX6OajQL5mi9
y4tvEjAUKyTDpUpPHIMEXqGvdV8ehpVdpp6BHoFJWDggbqUgan+cDEcxYAaw719iReT6Kniem20H
pu5bmdMgpvaAzt6+mxS6yFOLLDUvhi5LgNxnDU7eaQJYw7QBuiowPZmOdypmJRMSVw5mReDRl6qs
1iNh4Qe67XNktVYlXRwHW8GfZxie91WT/yGiCdKzFW8HCFwxVc+KV2Z8oRfQC9suvuk2o4RkoDgz
wQOuQRCk/Dl465Rbfaj3oYtS9GbNSHSf/YdoXKPF3vKJHSwFz4SlYcjb+Fh/6EJUm6TX+4YKLHTT
tnabBobeZKicSxyyuSlfdaLWM8J+kFBOHFl8sbZhsLBsPMM3WxgU+i3N4xqOxAYGWC7aR7UyX4Fm
XUZ6B+cB8o7zUOrUaE/okK/EDwaTN+BttRWzEFQheqjO1m9TXKDAGf4kOZpX7DXrwJnxv5cFMRsx
AMCCs1BbUOOzXBw/1I6Do9Nc73hDLEw9znRQAkpqMdXIwVXxD8vuqRGC8S19bsnWUN1j1lrIlsX3
DtH6zjkJ2LienGUt+QpOxGXzmyaxK7WV+POuu+f6/aPZXRW1OUcpXJnfQjgQRDly4s80JeUAUSqs
pv//sXr16obHfbKk4kRuVJd/me2GRcL7Qvz3ZwBkpCiglhKpaVORWwRvZtZ0liHxzp0Mid/mLz/h
Iei9Q7ZtrHiY3zBZw5Fvp6UWWNdCbWv7FTwsB0NyWRkhYHQHjAi8InSBN59/Ib9EQRGjW9kpJoOE
+/8p0TAFVlEUJuvFgxI9ImjBrNddom6gLPW7vsYKTSpZfsJdW/eVApN0MvqkE6VzcYmMLLchHSHf
Fdkj6Db7KaZyUvSmjbw44ZzlE4HSGwHoCNC8+yKR2WcrssV281sqPl8qXJPmBRCbl8q+sPLwiXGh
BCkF4tNCXWgtucZbTbH96IYdz7mhGr7sdPpSVkPl+OGbdC98gXdZUWOFGBUtb1zxxwf/Dasy4VyI
9qmFKhiuF7ftpVfHsGOPJJ3l9SpdS7L9Llbq52jaOnbjXo9o3qOODlLuzWXjDW3qa7BuhZVqI2aW
3W8GczrRpVzR/lBYlzxrwqFEwz3FlqG+Q9fNlZo3iaFXw1yvMQ2BnL5umKJdaGmAv/6bObzrMJ5R
B4NYCy1ZhNVeqFtZe6r86Rf3RwCptFPnBRkcY0IhhixHyX0p3dlbTjURPp6DupjNCda+BzPf/n46
Gmwel9a8QkwACpqEcKhbpHg6UOJ+TuOqlFpJEgnFkTUgYc/DCMbWcZhUBMPyu/6BzVSEaTnWEgP2
opFwwXgzScPY0GPeP4H/bfTgEYZTVTIEQ855ky4pPfyHFUIFxelJmWVg8EeINZuB5hIxsMiIsHG/
vZQw+qJkU7yYsBxovNZK16m9BrJsXIkTznTFLDm7+auuHuq7T81+fsNtHCGz2finUhZbP7rEQHC8
M0lPfzdpXy9c3RMCLXpgFKAb3kfAzAGdeZUV8yQ9LxzSL+i/ElXQyqYgvaOWQT7RXpotvaq5uwOH
lagPr5mBoOy+ESOzGyBjJGt/d1C6KZuBEHC2uD7xazX+SFb9o+vCd7uyY/IeC/ZqR8RyvadYOMF6
bF21fV6/euzs0NzErrnajwaXri1K+7PgWn2FJHfvLuYVXsiV08atdPF12YB47X65cQhISmhKV0L6
YIzPJsbR3kHxW0fQqQH/wxMuOHO+dYlSWrNsTBAr5QKruGS300DGcDP2Nrdaq60vMf5pBU7mXThI
O5DKRRON3P8t3fEVGCjdM8U4wIjUuwdux9y5uvIbtr5DRX0mCbsO12jooNBk9YaS6ehU4dSVTMDB
vkE45Md4+M5ivHhHxHF/Zmspa9T7Vg+N15e1o9DZgNcbtMNNMqShTzl1qNeffg0dZktVbNp3rTZ3
9qX0GVwgX7CkQD9/xPV9dMad2OOYfLFp4KsJSLteSegY948k5wGucBhmHlPHt8t4EVvE0AszHkaN
ATT15AgkgZzyNbMKMVcGHe048r9R7TXRGCUWWfHqrp20Hhdk4hoKWzI8JDs0BsLE285ISlsSFeeS
ZnpHSCZ7tlnkbAq02WEkL7K3zYhgyKx/eoMGOVkKLuoXASecb+yh892l8Dvs5XY1720K9CjUj7xO
TlCsPGt2o0Wq2ijwJZaj+YD9VtqIIzmFI1GNjt2XnB+i3E6cqFO6+XnC7u6pRGLSeCCJK9L6Cdrq
Dehpmq7S0eJBwxVZBetuCDxov6hzHm6r/+u//MdJH7If4pWFbxnLfILK4AB4xa0sXkAbxuNgafav
38nhHgbrcbm8VvRW7+G9ImtmM02SqXOKjPfWQIx6WQIq32aIvBkmomLBrLrbwnoTgbvizH0r+lJu
CqoxOyoRaYi+a7Wwo1DPYLbuLhgeGT7LMDj8BcTMWs+AsdwU56yhNf0m2pgy2SQt4ERZYi67KWUy
PbR7AOBBafOP13qR1ztk6VDoSsyHKSqGj4slyN8RsjFM+W00P06j60nKaL8HVspFX1z10wblCFA0
+fm97eifTib5ROm5pqKiMEEkEou1ZryUxhDfQJh9sllQPoaNDk/pkGfnSV8NE11qbzNCJwL0feKH
RHIpLpfUDT1/mTyggvwgmMP7VIDuJztKhqWlaUNejNqDFc00/bmbtbe2OIjt9hgzRVvxEc44l45I
DIHSGIl1E5lJYArl2PZlxgpRjs9RysBGAOIAQxwIZezY0l57EgvvtPQLr7315js4QxVOB3KW9Eaz
HkN3CsUM9yJLNO/UnRPJfvQlThom9+j5H2GMZ4L8Ei77hRK16ENrqVu+ma7qO+Tn4dOTt29C3JSt
NcYq40iuZtT4MmtPyNgtzWHaYVMNPiDF82UbPOu+Jhiz8lB2RPn+dcfxkenJABPQM5eiYKYJ29lh
chHwz7Xvq2zN/SYuXwyF4XRwYEfI2S8HfBYYbVl+N935SgeAO5jKPH0F/PzzQUbHI+vSAwTT9jMv
s2ZI2uhZGfW+APjUG87mT82DYdtn5kAIlOGX8o4pb0MHX+rrzYicFNj4Nx8VMXJjldVpG1niZrVJ
QcWeYdggmAp4It8gLYnSlYSa+URfiuJfDhh8D6IOGZ3PDKes/qYbSNaZM6Iy4O5xYHKs5iScy+R6
Go//uiRBvWMQzk2Xn8dSQHsRLPYL2Mf8qAkqt9xZX6WP8ACvCoiS1ToqcCqjyC0RBNdFaBOe1gFM
+hXoAbFowl+JaN6tHaw4Gi2cyDJ4HNd224BYJ00ZGQA0kJdD7Vs001d9CFVGFpBng1DUsNVYB3Dd
HbSetn78AdkmtT96ttrx637sC+HxZA0gu+kKEXDg/qBaRMNjsq3VsxBNZTxzkGM/ffRJi+/ED0+h
j8QBtuKe1oYuHAek997NJnfsk2NOa3I/BZeioATxEmKbFqce8xMWX6MqF+4nYVWqTm1UF5m0/z4o
MoBNHwVVwOSmcw8vV5uazVjO+1mkPledHZd1ff+/i+YmX3Voy7Dy825Ina+zxicDpkSLxYf/Ftn0
G+zv4XkyX7f6rl63L9QUJFCMxflTJWVaYWB82AmhfNvnOgv8BKNR1zOeafH9Iarl2QFWm7zin5Yx
f6IdH2kgaTeOD4tjsUxTkSzNYUnG3S332s/yCSt3bmmrcPOprWcIJKMtdZ69aTli4z6LzdIEVS0Q
Aekp0k7THqgrFShDt9c4s0vkpyAW1ERRd8jx+0l20XzUJnWayUPIhtNwJ/plaNcTHNlKtM/TRprR
7tzcFV4cu/Af60Mo3TDvypQkHTrt/6VEwixvP/llYcxRIUqgn2mxynQQpVnPvOOXq54wg6CDA26y
RxiZitkRFGBfr+xw8UkSm8qUvW/dXMzQMTyN5S8gfpULUnFepcap9IQCf6s/eKz9fF9hDkm6zCeO
QoK7386nSrxFFe3qJqF+5Ou/+u+Ar9yPWITwBrLbSYgUlzZVzLm2exE0/bCpjc0yFyalNtETO+uC
g5Xg9aCGDmQDElqHcezcVWy/LnhNTC7zgdhXIND2ixPqAN/upc64zu0cmAIXucGQ7WJuxqET6K0c
IZNkCw+DaMWnnZuCkF/BBBHzEdgIZR0CYnwsS7Rx/Tnfc/nf2SnFAr4kqVcrPHjhw+fJqkp2eupw
mzSDUq7EmrJfiz55Pw2T8taeVygNGtTKy17tvBjuDuW/tTz77ih5fD6SNrX7ouRI9FDEaGugEItg
aCmP65he+7T+PETG8UNy8lPHYiCk8etDi5fFMbWDtaSMsdrnCYP/8IE1a0ARPAvKesg2SlGpPgSt
Q9n4Ygxz00KWtoasJuC6bN6vtwanrAN3dCLHc82pvZ3ihI64a1FNpY7DugqFZ2fPHO29RXO2kcWo
YHQvI/g90zyaND8fi552oq9e449w0wnBtxl2xxLhaBBGpH6X/GpjxGZa70n79WHjq1UAp9jZBbJw
+hFWvfWYX9QIgEc0mV7hbSNKEGDP4c2Ynap3PBeovu6j1AgEpkhfMuyHtpimLE/BIVh1P/1YQFMJ
2tWM3ekKHrgOIk9gMIPwIQbzLoQ/oe/t5C+BW9g4VOvW2cMw3+aCG4HOrAnMOI0dmbSsC2HnyNY1
uhsDrxfsWI9wHQc8SwkOGmK+UYjt4Lo1Gbu0QDNgmK/rZV4EBBSrP8ykvizLSoc4ed27+kuIs/WT
kLEmI0K1km5yVF9Y8Ut0ueRXcmeyp/6WfT4uIIcMDbBzSHuXTSMUP1UJNodMTNx6pmY5xwFULGvW
ADR12FopROIRF7ascWHdB7Y+/ZBHZZTudCdUAHS1vtLaiG/Rx5aiUF+q2PzT1+4usLPYLRCgbooS
X3ZBn2YjO9hDXH2DIvuqzz6zP1fIA6Q8ApnL60IdsVQyHmhWk8oS7rJ4wnX4Z3VRL+J75m/Yi3pH
G4LaMqY4qwIBM4IHcWBQaP5I1GAMKqSNLjliDdklUrfzo5tW9rmX1xeNp274KDn3eNPu/d7lO1Rw
IBBpokkKUz9hNnq/zXzctG2cKVR2X0AzsckaHZ6O2J0TzS6CpjxLblscqDJo0bcm6ChNWZj8Rpgo
HZ6rme//rWfBskajDasxkjaSpsrZCyPvODvryPQcDI+YsK1dy3DdxcFo3LJO5hZxNnC5fwMfWxh1
2ds9yBXKBLHT/7Hh1xMSAOyufpffZxMEk2J8vNa1qlSH11eIJ7Stmzl9d1kIpugVp/csxmISzTQn
twOgfMne/pfKiN0FzSynXGFhjPc5PAOJjYoQGo0JGc5+NheNRQDYgke25Ki1Vn/fnD3J85ToB7y+
F/OXoOKNrNqMrcwhTRA0qlzACAKcuhNJ2LtE5DU1bVhz1MSpljYVhCqoC1R0dZBgAYAfYvTeIgme
cg9YtxVkfAeAHRclaOyhWyH99gizMHkKm1lHUxzym47PKLF/JVyqMs0kWZEFPgiPikV8wDfv1poz
gk8u4qwK0r0slkOVImEphiogbpxSHwZFkglh/jAUvxrT9uyOd99yPBwtNNYZMMFIzcRPUMjolnGU
Oj0ERqnFpIOYJDMepel+4FzLlwMfnN56tlRpVE53SFwxaWdRE1V9QbyIRRd6XbVHtGbBVXgRYiKK
KHKWDiKis5c7d5MCImTXV0l/z5+ImLJ5+93VF7oPJuyBdq1QopJhMpyGWBCqMSvWOje3UDTmrrW0
80sXLLAwlJgVkP0bQp6OF7AW5VTcmx+/5JPyXPGWQplKQ9/GQCI8OjZXDxVrS46woeR7ujUMt4r3
aQzWZIa1vKMlMq9tqaQhCG2cPVWKcypZpiaZOLCUx83352PWz1rxkO++Ah9O/FwSoDkwdMTW4Zha
cxeQeZHFq/uvzNe0SaKrY36WehpR0pKqUuLbrTB55Y3QI4SYFeF35CIpLMZMJd7pb0bf4QOIiXm1
FHpvdaG3c6WOuN+/NqEDGxo0JgQmzUH4GPIOs9ASfY4y6mIukZ+gt0Zm1+XfVFYNiGtc5p9c/vzp
4IJR202GGqP52/2fcARAA3Qw8SjBciji3CZm6l9UjLMLa9RoBxN4eZtDI7UT0ws91bPx/6HjrLrI
h0COvgYopuzerKeQ5YST+w7skbRPo99ewdSoOZpNLkvUWb3OR93Elsid5UNW5JxSo15qJz1B1n1t
4Abe63+SOC4NdxaTH3kapitnkmeLedL9dfBnSI4UjL8jd4t/z7mFT+8RYL7HeGFUR3muc2RfIrqD
1Gn//VGmKEQtJE9WkTNLqb0VD8Xv6WjkY9s92Omo2kgk0SFvxo7+kS1SmZjGUW0iyhDXCkdnxxxU
Zeo9W5Ais7X10xWxDJGshvo294VJxRReU6qky+s0hJz/JxZQJa5YQ9mTmMSGugZR50jxzNsaDGyO
0bJ9/VGc+8suXVAr5HFsQq8PQcr3I+VMj5lB9oUf7K1/oCvvHy1XryJ0QApKcC1xaaSZPtj4Glbi
W1lS+k6+uAN2Myg/Bxp95v7w2MLyHo0+AF2grOjaGfWjrhvYwAs4m9UuxqJ+dyku0NDmC7nSh04r
8LXuvn0lLRcTorHt6nPZ9GlejkGb0ViwfWnTt1A1pY5eMliyC+apqLIhvuy92hTG5r90Kud0dn2r
Rt2XNzTBfFriw+z40b/OwCIRZGqasQkIT5uepu6mBFbUyKvOl9tK3Uxg0FVtChud8y8TH86o7iEh
6oYV6SDUfiNs/RDd+4PNhXVb9j3+Qorw6IW+vLvNGcMNe9UzYzaRu6Na4JA/JdNIMrfFqpcKBFPJ
8x5KKx0dEKh53HiQ16WPZhHUBSL5u6yv05fjzW/NXMy9/RTq7CypDLlpEhK9vOb5bY0vGak8lM+0
On+sqTGNPNA6StNFqHSZD34Uzi8Lb7eWi/Hxtgz/YmLKjdLA5Ae+0lv37a6xeTxD+JuZYpkZcJpk
4xJunt8j8wTJI1s5ChyzMGfkm+yyxE0xD23w2XqEyMAlirN5Nz7sh3V2QWkmwFqUPZPN1HdnzAOS
37F8NVOynTv2UL0Ci1MGQTGDGjQHmF5mGQ9hXV5yCQhmRmLEsQlXEk1M6yyYGbnQYWsSa3gPHCRa
YE/e9fwuU25A6eiBbEkRGFKwkRp+KsguGMJVEXC5l9c9Ai9Jf6Vn3bUuNPG2JjTIaO65GBH7D9QJ
S2YMBS3PQPYesKYfJ7soBBAzh2NAYhrMGwFr8kbKxk1oSoa2OE5BcNw0A46fgBfESWt6YH983RMk
kCo6oGCHt9tEd/uIYnBnfGA6h4oQYwDG0Ss9RwankU5IRNQNipw/bIt2SUyLxmj+jJDkjsitIvuM
6xBTCHt3hLpuZZqnHqHp88me+SYLd7Iq8pu29Zof8vGGl4tpQxZl28vSWW+gP3/I4sKDCG98enQQ
nhykYE5yJlJNou/WjBXaCPcTRxm4BWCnmuQtmyHEM3jzZPJS3sY3atMowN+KShVJs+xzCpFeo91o
LxhlYJZR6AdxyhbMLZw3ywq3uWab9/9xjAgA1tFWArCZoF2xEzPZ98BN80o8S+8/VEIYaCKhsDOm
qXawjjxdv4LUUeUf9OKSmXpkgVlWaNqjAwwSnAX6XHMvixqFwpnfVYR5q1b0cJ/CN6VpmPe1LJeL
ZlE84tXBeQGPzk1MyU8ImXYrdN3wCGIW2CYRCiqeZM3m8ct3/wfqDwy5V4sZ/2Ub1oNOj0Gn8Ouw
29z7RC7eOFyEU+pWTM5lDHk+R2L/rv/iF0++sdDKuv5033nrwoBYmzNAgQL23XNxP8uKl6Fcz5H3
8preVmTMBKzl5/4VRzeZ3brtCUAUgJItphssqq9zi9jB0Y1g2GE2qpAwrq8xN2T8fE+F8fTGimaP
YOcZGkhInVa5YRzwtWhUD3VaHpG+SEjN4tpLbXv8XsI7LqXXFj2Hq0yGQH2srKshE12C53E5NsHw
Pt/Zj7FZ/dkHuL3RILTtp9uV6hUThkQtstb0Wtw95IDD0qEnWd6bR0sBSWqiObNeJYHweljI29Hp
/la2Aw01Skd87keq/QRigoH+ORjQ7FGHHu8W1V9pNy6gGGxfCeOXs0L9JUtA8orp1Xki2uoruuoc
ekWyPLar4xSeTW65IhFOWIMKFhOdUVWzB0X9xnhvkfa2oTRKhnOY0i8x2gBWq5kB1zp5/n7D9VZ2
dtJiOzDeP++PX5lrDZM5nX7pri8JGwh3dentix5zPrC+vznoOIwk5mFGVb/4WSGjLKNA5y+1L9EE
ld7U3OQapT2wKDx+0oAmFfiVJj25eSHfNkXjVgOoNy/gNly5aVCVWPwuEbqkgQ1Y0iqCwNox/vj4
sm8ibQ9dRMeJ8xwzt9AFEiJr9w6CFD71caNwamzxD32p2YQgMWGlmyOTh+kXLmF+eyHJHUdH/yaE
XfywJPPlz4vhktKmlcIqYOI6XyORwBJxejImwr5Hb1TrKLWmFuoRzETO5WrppKt37HKhs2CfT5zL
j3z84FSs4DA1NXd/ZvLvajSd71oL3Q8cTdQxN7x+CuSGn+Hr60XP08o2xdvTJN8YmITs/Is7XThv
MN7/gJ2T+kXPPI0BQDakqrxjWOrYr3rWcZBFBQKWQx87YEru1OWaa2EondHyl2dahtrAA/Fr/cbE
XVDg39E+0TcSCm1QOpcPKU3xG2gUG+UU1zdPG3DKttMf4l7kayS1rJ+uet3frm9XGJ/xeI0GgGEP
2CYJUNh23xqNjPzzqK4YNs0Qg9iJutTVPhsjZMOtBBtEj15+Dw2Kxzqq80DvySsRWtlARFUWMNJB
EDHnxt6SyXX0n90K7AE2kCPzARTrX+V80xJVV9Cy+R3XpzA9iJqyqHxHhXfvxpVyGRTFd4cH8gVd
jVWkbr15j5gXLp0jB9F+8a+Y0c/V4cvEwaJ/XoQFY1oZ/j3FZ5VByIvy3B9ZrHQKyih73vPsVFZT
YwUAufoTIpWePFJbxSU1GxUsTaeqPwsJ1/IlZvKXym6ewBhREDlT2vhoCxEqZHyhBEq5vqDPN4wA
CpAz0ymntpU84DgpS1V7yQzaOPfcPJw4Y1m3+x5ilc+4rAff8Opdjd69yumvkVNTYmHf5KH7dQF5
8MxL+2ul5kueHZbWWHBBtYtyeixo5liXKyeNJahcjpV8zJmxsGe4CCqmHf/Tp0ORP4pgC5OH0BXP
/81dz3jkgltNABJky1P6Jbcp4MGuS1kopknTEDPEB1xerWqYqqNzpzBCpWaZjrAElqSj2FXl1ZX5
fhA3r0kf/mabgln7jvEvK3FUvP9rYd56ymj1KpCodyRd/FKTzCkB3nEKuAS12l5KrTLZ0uKoedzc
lvh/jJVoNkbR9La/52ws2E1aBPueiFk8nMdJJ67BEtfSTGU9oz0E6pvpuCybAv6SiYvcr6HJK5+4
czrpullKwtt+wiB1FahdWmLTOx0Ayu7AlpDjF3AZ45FDtUvbsjLWPyDKLaePv0miaU2n2jxtq4Sn
K23HMCDikg1Db5zNZhOQ6f4N+9X08XnC1/NbbEy7IG5wnyEe/8Qx/wP0vHLN3fJPWJuW79pJLIi1
otX8rXiTt2ZhIP1jqzxrVOGvkRCp/mA0qPyDvsQpSe1nFZ56DXhWBrXfImECWGi9DTRPnrcizHj5
n2Ws1Ao8eo3Uw2HCzc4f9Y5eIvx1iMzcsxPcyhKLstpUgtZ+PrA13LcA0WBODpybV4X4+5z/q93Z
OpQQ6zkGzwwk1J0XKfQJV7OgUYzBLzhPfrOfDsZdJZXTNmW7DAOwUfxlLJJ3i9VRzoVrF09xWv54
5jFDS/1n9mNhWDVqWKfg4oUg21J87MlqXiTwPt8dMDr2G6uW8JCXnEXsgkmVEFZ8Dw5KNMgrudlC
Hx7PoPqxJpjDcMAuNjVnZAs/08aeQQGH7VtF8ZRpE+HXipH3UvwEHUYInCxJ2xElz/WSVnL2W2cX
RvxjKDiC+WguT4F0hKR3vvou28pe0lvN/onUtC+24goPw/wVYuz9SGsvQCVJrDhJl4n62CwJtNqp
FwA9rPZkfOL0xN7QJN5CsEqeNyQZpKiPg2tIa/zUOJfzHpFmLi7w2dZkX012ePAr48j6Q0k60feF
Hh9samOSeLZAeiIginaKDG8+1vJNRNSU9dYwBagVZa1tUjcl/zp0lpFeYJSS9yTIcyGIlQG9290S
WboFcX7uIP9l18LQHLlQQxHjjhw4sPio4qJp4EBv5Yn8WeJCcgpc+CsXJD21A7lfMcW5LNZamOQ+
lFi7hOut74KeUe9bds9rq49s+xASQWacvmxM4IL+L4N6N9zzY7MQKOgoGK5o93xbtO86eoyyvol2
+8cB6mxgDXpvvtSrOqB7oV4ktRMVwWn9NT6UQGeo34BCUcVYER9LslyQnAZkZFkuomOwjUfQsF0g
LFIPYcO/HmBxxx6DRfqnPvCk1UWyCM+LhG6+pHCEZe6k2EBoN3m3mrPmUEFUvltDeSX7DA6A1ZGi
kGctOj1skN9Zqhe8YsZeA/8ubn5xGQW0FWjSiYiqK+Q3QXb84Hsn5qZQXZcIkZULktfZNwVz128/
ZXNv2t31VYQU59BCLplPYO8bNlut5/DZB5KDJgpaR00uizvBhp3is8dNznwOUxp4yGMQp+QnF5ds
rAOUSvdrGjlCh+LX0KM2vAiECXlLe8RJbrWp8CTZ1iG49v3BWaUznxxuvOnsAFFDe7zQAZk2izmE
vEBtosYpYUATbybUmBGXR86R/zKaxO3HqgIDYDCo3L5psdC4Yz0Sad5mdbfVS99O/bMlR1cChGIo
4J1/iIUMPD08st2TSTPSjfCS2dCduntWVKbhh7t0Ef52uOrRSTo3PdX5g7w3HMReq7wowNhB7aNa
Lli7ym4zuDEampBVxGc66tFl0VlC38ijxMpywYkoZ9CmUp98VIc0PNclgWKHpxeeD4qP2SXssfQu
KYtqzDWdEDyxF83/dP+LRfvMcaOkb0zSrEXpQBXwzMJ+K1d4FOBlagV5i0F7x6XfVZT9a6ivdTmV
SBBhUlu8lbt5sLMyuzcQlo/9v0bB1b3HrkI1G05xlOuTj8tGb80JdjCJBsgvhhcWe1DubehVbCdz
lkH2BkBrjNA4OYzlBwBvJSWlKfqfQqmpbEx1zRMEaSKxfbpnyYLRY9gQ5FgJyFq/xNBFO8V+O7T+
u/N876S2rL0S86QitR8t8L9MWJl9annnVKBY5uCP2G8PCFIz6RKYRGvr/+gOB/x/1PyA1AByrxqv
yN6LkBt8/B4AnuqvnDyoBhh27Fx7BhgBMP0HQTaLs65cOwFXnJieIIltNjw2gkVN06jD5DWeZhLW
mxi3xJ9yFXzSrRIRogeqdxxK5x4x3H5qRy0ZswdRIKFCxXur8G1S2ubRMCifRmZZqBj90N6G05rF
lkcPSECXDMHMByelN1RXUcj6TnlPOu/nqZoMbop983mPspcFUbHnhJ/OCCQC+/2T4YugGrT/4z0H
+8v6M8U1n0AcITGlTe9HuMr0IIwteiMcLyibrszxXTiFye0V0HTX0MekACgCqBN+sIZRFqDw45Jr
D1VPk8PsCcN84/kq7MX6KWbBF92Sv1Nnle17O8s+ZGVfPERPBYrZvNM+0FSg1PWTrBFAkAHzGkZB
H4VpJjpGxUw32niuA1u6ujmHVhs5vAbJGN+lo8mz/jMUgTZY6h3cy45zMOUdtbXQSpqcNNFaztoz
4TfM5HuaPLVphXww95gjXADtrBDBhDuPHVwfyWdrB/eYkef5lJXvOhNeHLUhqI/hfFb9Z0kfe145
FgLLYhCSITjejHMiSOxBjxzQPCEJTL0gomSAgIJSY2Gm8Ih6DKaPUChr2LicK63+gWmNhni4C8Rk
AfompYlaf2214Dqp9ip6o27ZAyaz+1UM4NylyaUbAjdsNoKJtP4WxaGUIHp/M54PpCoLTFoEyFL4
GuPl1Kt30YVMSUKudcxdWlSCxZhoOKY7yjya87XXr+onrt+/xb7v6qk5lVBFItOcd843R5iMDYsy
GytVxLDyITp5ss2Q5pPKV0nEFzEg9J7YUtivU5KWvmGjkzcPHziHCT3ySzv87z1ksaUcmF4+liOP
YQC8lcyz1bm86QoNY913vJhh2kYYSR8qIxMtjtwfBCVMNsZfYdGV2Ep+N2BsHexEVtQ5fbXsVDPb
2lsl5leJQzZX6nEMzvDYF5VGinYNKcK/EJgyv+XNiplnkufDZ/mmA+YiwNf8f4r7AD+MY+sv0kbc
joIkM1Q+I8FYXPXbKUSPfLtPzicwGJ6yVk+LYCBPQG+xyNkxeYgS49DhC2IrQox1MsLEwHMQkV6I
+3L75NwoToajbCA8BBQWNSpuOqRnUHt/NgCjIPyJlDRTIBGBbaulmu4q3qIkrJ+74DgQrUV79oNz
qez5ZR+fcYrPgoSyXz5NKv/EQDEt/+tKa+jVs6gefAKQEDvenreiKgR/KL/KoN4xU2oufqsZvHI+
sgkro/3sn0mpt2EsaR14RUND3gbIy57M6jlfsSo1asPd4x1+v545w9vmd53OuKem2XagF2YRcl+H
013zZSYsQW0E61Rdo6VS57EHAOzw8TGkstizo2UsRpYTOzuur2Ef7f5r+oc6BPm/ExOWBIhtLO+o
w3VP2wN3nV9bd3jxRArSicQLcKNnw4MiXuanOAf/DJu6XV/tluadE80H8GXRQ1yRuWlhLc1C1xew
k7A/v7skaloxQfG62N9p3noPLc3ueXdUAVxGXJEiMlBGHt6/1+KwF1xwSEXMafFDCIPh6uZtImnJ
205BkSgbxWf2xLSZKEJF1wEk7Ovn7W1ns2ISUKVgoowm05BErZtdHaHA93tn4hrGy3iuNhKcZ5jF
ArNNF9tnbQEnQJwYjFPEQ7XLRKzHGJCOxqLF9TNokqRL4m61j2eDUK2kcBroKmcgKhX+SAOXh8tg
nvSru+gxSjfrL9TS2qJdkIRZwT1BOsM7TtLWxQBw8ynsQaAXmtYObBb0+fD+RTPJz9dFwALaIWT1
i5JGnjVOK8f5WchAIDek1ZJ4jokhjAQ0bNbWZPj20K7zmpe+Mos02kmky5SUvh/snT2X/4KXOCcS
VMQnpVz2I7Dk75Xqk0i76iGviRK9Z9jbfOLW+pVHC6H43erd/P4BakmiZQiE4FPEW6p73X81flt/
80550PbaFQlR+D0/kDmxnjKsEDTX2zssWqWr0Jgqjk1d2Pjra00vJG4a6tsWlpWGm3swLpumgsta
WU2fvn5MvLr6ZEeHn9O8MexbuHRt1+KsFrT5ddAOXyFjWzekdcwaE19erIQtvcu0ykakRvF3JzWp
Ous1j45j8uTpu6OxquKWjRdSicp9cKxCpiuz21OgYWKBwpvTYkv3XGGFQ6iS/jVsJgKgquAHFw/1
VRTuk8B9mXOjMvRj8mFxue8UYsfpNxfX7LBsP4zMD2kNVSOERtzijQjOfbwTgNyevBsmvy0BzeWG
q/F9i2EUUD8K0hRI/y0E0p3Ma5/pKshT6WQLXtpBUqHoJs9sZ9g/LIlfeDNQeu+IXqwa6WLEvzmH
V33inzH9fkHQoZ4aKO8ZQA0U6Cvjk1dlj3g4HcyQ9auK7BsD37CDfLf4/S9oV0E9IWZWtjp2r+jd
fnSITwFU7Ej0LHlY/Hf0DWOqdeuuHjh6sVQq3bn5XSbx6AF6Bqx762N5xoYjac8XTAyuRNIa+njx
SuDbpAT74+d61w256fJi7tmHedWosCJdGj5D2dXJXHT/pr+0MnZAUK1SZzJNms7V1M7BDzK4rmxP
hea+Ptr7l20FZf0PLm1zypEhXevKR1cCd9SNvjZh+/9afw5P0n20R6QlC3AVnqp60oY1kYalmo5T
pGkNKW0iVZa/RZ8rlzczaivFv+nCTPBOxE1xcI2TWWHAjCU8mtUX53bUSDNvptml2JxlAQ/5upWE
JNEmyfaWd+fcTLPI8mnhV76ny62i6N4pgpUtNVTAy8YF59QvCyCZqA/qsix1wu6XKVTh5JP89dHg
lOV5VbJFBMZ+4eWgWVitd01wZLvIBy7F1DWnQ0PJ5+o+XnQeyXPiPnng3z1PZyCGsH2eIl+zTNVK
Ng+eSJno0TwI1EwBYWStsp+tGt6GvvLq3HxE1Fg9/8AtOqT0JPfPAcgCgDl4/0pL7kV2uKG5jKZ8
aDVZzNim8A8dkYcKkBvIjxaHDmCZ0l9kiFPeU+GNfVV+bgueRGBNhw2b84A7rjNpNoqJQloJBavx
2dU3sGM5dhg8PCOJ+73udP4zycyTE9WiQCuJWG/jyb74rrwCnIX3D+ns2HeN/GJh76JEBWhjYepH
mTQtULni4LrHy/LJEhl8FQm4X1kcg8IV4hqowEH69s1l6yBZybwb2uVSkunvY8hsdt7WshtW3nAJ
8C8RFMJka0xroxmQu/scjmuvjhWo8ERyQkBc4IcSQnFz7AuXhvuuU3Cp0WPJXAOi4QjWXUNfa8Fd
U6FWfne9Uzn4tg1ejgsEAYkveU9e2iN0dcBi96hU1JolwQOY2DQwqAo90tijkQbg+SPD7822CV6x
VqWa6DifefiVqD5tXsGkZlXNGER461s7yn0qnkd1+Ok9RYDBbJ48konsK3tTbN9zCA9Cb0gv1mEQ
WYkPx0CxrPuA+C2k0L1wVDvyiHLQRjsntrkMqJJVPTUrQFPoxoplgVNd0CmJd5GSlkklpM0kkS/T
E3ZrVCybgsCb9R8MQwXBbS9uDWDnxcSuyH5TC6J18HnkRU2EDG/BxMwJm8G3xL1md2MHL97vBsWV
pAWvV2BfOm7EK7Glf2/mZ7gjGS2VwgX/pCLJ/uWGJ7vepZUU047YqIzDvCd49chQ+wBJW7Q5qzzx
QjfzXS2bNe5TK5JSD18gYhgx2yupGyo0Pc7qjFfkUJczfahx7yboXZeGImxFLjSEQgsyATJRObnO
UAZmHIcSJ8xp2iX/VhaveRn+LHjD6/UZuVyNf1AS9X3BJzeTblTLV2fRpuy9cRkgIuunefhJMJHJ
hROw+b8/4z83dDjYJuyJJ7glCxH3cuQnH3xoiuaKrq0o94BwiDbdyo/zMP2mwcSrzrphaulW4k98
heiTPI2Jgy08f9Ue00NNPClVFnfuG0BvtP0gHcgaziLF3f9hRxz+jewFwToEl46iUqygW/1CgsKn
vecMWvXBWslFv7OAcoFm69vbhNphw0hVglnUp7R3Ar2ka1FbCjxk+f2b4i9Bcuo6ZjQN3C36FB3Q
Np3/0jzu0mUz5vaDNJqPSAQkhYIZbGF/hZhmHy6osK6BnP6ZQKNY6sm7P3kU2jsV25FkN+xvbGoH
AgRoOvB3PiQBnOUda0Gb+0CgOs/fij4MZWTqVMOqLLH2qVpLchB0isCuEvUTuVkRNDOoKZFDfpkS
+ZzHlK8QRPZDBSP4lXGVJcmV5SxQuERAxtfHeAWiq417m0dycXXvFI0HcTVoh4zqdy3rgZP7sYAI
LY7ZLQ0arv9W9mfuZGrkY0qFgAd3wkKGz8BQqIYGLgK0HWPfB8iKJjPW0UKnXvKRu/SINh489PRU
72vjF4t9+U7YR0Vj12Y9IvqLrSQ9DBbVwDG9RNOkFN1zBH36UJdwMe17Uiruj8P9vztzhhQQGy0K
LT/EYEt7FdE43ZSQCREYzm4Jk3n1yXAAh9utSAGKl2f+zmHaNmMEoGUy/BCTJHcJMNNAX2H6Cyzv
ZdjaommM4DFES+M5A6i4Y1DoIxskMuO8KlYVaMqvRoIO9HIx8PWuNr/5AFD8BiOIA18/wJZKps/u
Q4P0NheXBS9UJx/LddeMrAxIYYUNN+CiNQChGIjXlQH6yLsr22LhVIe4YprNKaFLSYI4cjZccPAD
aZ4+TFDdjIxAFxsP9MdJB5CMzkn7oDt8DpRBLXn/UFD5fDm8ZFR+SZQOoSqF2o/WHHfS1yZQYz3G
+ma5WLquOzVUjShiXqjtF+CSw4w9fSUPvA3WDZowBA6bpDiGzedGhnBjOBBICmzp4P2wMAGsISQQ
a5WEqBZNbHPAd+CuzecJEnx0KBJjZTgF0o/wsqfiibOXn0WvLTNVQ3qXGzbNBwY6ZtuJ5AI+0BFx
gcxGciTISZNqisxrdHD20BddiFTXzzna4ni6c4nRtlmSSpia7EBY0PEa3+jlbK2+p6spoZPrhnbU
nMjr8/JQotOXdyN5/wUmItwZhOH6ym4GZ6GaqXEy2stXwwFyKSKmWNO+3aFAK5eE8GTLT4IcdIu7
XKnZXnUGkXnOE++VUgMp4oLA+m1OzUhGsTsz9hzjptWKQbcR14JxGXBoA8EGoIQuPnNdGsM5tEq1
Ljy9M/VIQVwlJZCc7MYsxENiLEHNq1pTWcZfczCTMFyjUKR5pYjmrTtm/qfCQ+XsudLGMAw7WsZw
RH6rpyB76yqVt2DS3/KdDuJBxDKGKIB0uu/AEHKbBdXMlWQL7iU9COWpFD5z2ylbx69CpYJ2IoQ/
trpaALwJZFpZnBSV5OV3Iu4QD8HPIEsLR1NR658IYSoJnB49s+nPPMWlgsUbgZqWro+oPgAMZ8Id
VkD8sHX9SK5o/ZKgDjyJjr5FAlfXRnwxAUBzsOxITfsEqk2TD86GD9Zf4F4Hz39JSqnBLXGmsqWS
THF7oG/1emupsqFbSFzXp/HUJ2ji8kKZM3zhmGKJYa/H2V2MHIDRMjzCAeNd/jBPML26GAA//2ZU
K6/RSPwOQLKo6+uQ0KCYxdOyt/u4WFzk1igUGEDgcoHSfSW2gy5tvVP72kXHi5y84fjortXaE70F
p0bgkqUy+qHj8lmYA23FTiqJ4+9WSSjFznI1yyi/0RzIKB4T6U2rPjrZ19DUAxZkqgK76qy6wnxy
11N6Vje/GjrVwoYD72K1SLczKLWRak7uvXPFl+sLUE3nAOk18Kq7E7fLj6HsdBZHbjT6v2wQodjU
L7OXc1OIFSeSGGhtJck1w82QQz/EHjWuBIV8nK/celtSUX9t6JTHROGDzQfoaT6pETpRMvVbtwKq
p14Qwxwt3TGT8iHTcTGDK8jcy0p0SruAEiKASNKIe/5Nn1T8SO1S6rf2xcz646wXgio1KK+BXn3N
Y5Jnde7uF8euxLaBOMGStr9dscaMst97FzTp5kQu7IKoKhA85y59ACBIxrHYAYyg2+NyuNkQjNn7
IVDSprhWwe5vCmB3EfaN8D/WPhgTQYKvPsDBtMUlr4QsE9OL3qLVB/YUsdMQzfFWk7R8UN7rl16t
6YBUUE6PNVHXN9ub2ciaQO155TvI9jJZsWNNEnxfCKLNAuITdcEziJUWLVlE1mfR03UfJzM6VzaK
4Pc+L4iW+LPG6l6mehjWFiFQOQ1mk/Ei5M0fZBgXzdyEh3F5nTv3Rs7zuS/XjRJUVUzLM8z7FSKy
8lUIKnDk43W19ZH13z4lxxVDxqCZZzdbzfzGzyJbVU3RuYAVlkE5fVz4mAC8qFrpxAn+tFUufsz6
HZ/8GS6cL9VkSwlcVciwZaWSK2gCqzMmk1p2i/1aO8YbRk59iWdIHccSPq5rW5DIgFc77Zql5Lvq
xD4InBOGjpQCTt1YZYebyyjcjygDMeTq2o91oBHSQXCwSOi+akHXzG6RHAVlLtzhZkihPkUik8Pl
e+n0veYljjb1Ukom/nMfJouUOt3dswF/Zlb1sI7QAzFrC1sHQ0iCHkV7JjKPUrQgCV+7rfF7EPtb
Yrv2J0DsjubCx6Apy71s3wjO5RXaboJVBaug1yQvI+WgooVhEnKvt3mmGxk1ilwBNi15q/jyJhgF
tqHTO6bAUUajzTgTFQgHPHcfRYvWgZHZcJ5343AinA93i5vXV4wwKlm4d33lsi5PCJIe/gkQLCU2
hIhg/8f6qmezQDoSXrfarYcJF8MD9KOpjUTwHspoBvWgl8RuMPsCSJQyQs9z6/U5TVzx1Q5/pjpy
qpINndy+iIsUYuv4yRrniugDzqJwXRdsTZnMdeUWcNXFzrcSNkzD4eLbMsk8LjhvE4wF3lTJNMXb
8cBKL4110x/De0WbYWjsj4hxty3rEe9OqnU+Jx+kUWVECrgfyOGMFFMzE7DxuHnN8Mp967232KDB
mmylgSCxPBSH4sthbd5kkQxxz6ykajv4TZeIoJ6Pb69qR3RmhpCiurd3BNJ6GLTCi9zrxm+rDyY6
qPFwvNNrg/VnsQtHeHaHZlpq1prPWfxaSqVFXLuMJZHgqTFvg5VPwgL8k28wlti4lyLj2ursdEyJ
O8tH7pmD9mWOTo2lhYKskHh7LAM6/09vz/gQrNfOpfOJHCcpHoUc3TaYofaWCrawzlyIdJIrjkLl
gp8FwCV3BnySjlCOdBAX+It0LXCVw/Rk1C547oHwDrBCqhKtE18tpMcTB/3nZu/EqoYJRdP6yQDb
4DP/y1THs9eVW3WbISrPn/1twKi2yTHktlMGSaNcPBcFlhe0gUsSqwc26z+5wrlxR/taIRlqYee6
6Srh2M27YxvI8AJUyfXt+VJK9Q8CCKhWF8VUGpScZrzoOBArmKJMp5A377KaUdPTg7S464gkkq+t
WdbtuP5AtICsH/HyJZWgRPYrVc4W2sr8494P2SxlQyAH5gwUPEuOIgpI9wq2opYNcsj2RgitHLHn
HpEGSQzn/yKIW+KJU4VZ+WymbYGF+h8af/f433OdWaAGlxOBHuSAYUOAEqwQmD0LDAHDqS+d593O
PdLEMCwOjh4tkWT2kuNO3AFU3aZa8NJ1nqa8FFFLLWSLKjT4+zjkQ91HIJsRXN9WWjeHj4+OsL8G
vkLP1XWJFUuqc/iJ1LozclrVBlo1BPvs0y8aMGRlkNkD0KRm49w4gSekgc+5RzAhphsXz5LR5nK9
Z0KEXROTsQl7yChdGuK31IREAoVVm7Xd2Abdx93Y00XQIPKbsna3/cai9CTRo0XEP0GEoW8p2SA2
saDbZJG/wzx6Wu51tveazb8dU4jj1bBV1RRzh76UfmgfYuJFj+KmCUxi9SuDmmNOMJljOUfrfx7Q
fUenBWWjv29tWLRd5PIP4W7gEsJV8MDXlPCF8RvIEgkPlUdrHGdsD4IAOuble7/1DN+0UCVUQ0l7
UXrk2MncPv+l6HLN1Lionnbefc7O2FVwrXOXtVZS9hNS9pEiH0U/JOioPj0aCi9bqSu+LPR3SiQf
18mJlAR2qarPvpOGW9B1f+Bn8mJXq7ZKHnFduP1IwP/Zd0OLxQ6c8M8VDk3ZkXEfgj1jDK05ubhl
rN5p5X2czizM2Nzus92x4xoptpZaPvhrmlZKhO1UXNWIHIL02EqswZe/iUg2wZmoZaawn8UUGaBa
EYyPnu/fPAqL9kk8xy9hv3j+niGyH8zp2eAqSrwUjuI1Vcv1t1704NObRHagsrImD9yV2graSDn5
6IG8Dqmv+GVvH+5pS8YXAmqDt8kwOgHK62Lg+f9YQ0tOIVwGnY9g3Ny30ZHQRBG+khqA+yO+1ufq
QSAI4eLo8ohnsvpeFreWkgNU46lgyktKynI56R84MWxqS0LOq9gPrPzcwqebi0EHp87jxXoythG+
JZJBeaYgrJ8NDrnEvAhONc0JOgvx6yVOmg1QVgeqwzJeVeorL/qbpuERtf7TAWm6FT4176vgiBsX
a79ughq41Zo1ALtTtNH40zwrnCBdQwjwA6w/PKouMQ/bpJguiEjesC0W5+kBR8FETxhPIIMtMZMH
0lMWoWbcSWpmZ+BTWICzRKhOo0BB4+C0ZYguMds4W74CTwcEupCdJeI/P+O0mIjwvxOPYGPVANgB
5qNkZp9U9HjWfHA//IIo6Z9uee3aqrcvuaEwTQi0RCt42BaRD5nsB/1kBZCR4eIKLgO4rHzQT/Ka
kGekqT8bYhqhx1tVP8qEjmhIaoydec5jaP+HlqC6Fa/agnJeTjsNo2b8HrRx7c8+9o1zXOPHQRW+
pyowC5+nUE+axzZFFyDFJkiKsyvsk3XysbEoBwNYqxQgNAMM1y+OWO5ypLAMMS/q2tgD0l16F3ti
IpUByj/vTnXj2hLV16bqxtCIqVS3yXL/SJgZXS+IMT3Pirck0EmpHWM13N5A92rANHOEvRxEF3gu
bLFlLQDjXdspnJBGmSr5MoAAOm1Tktv0WOMgMwha13+G7OEUriIn2MnnZp6hPNVrG2fiM2Sxhi12
aKDP28gqejXR2WCn0rSuqvTKLLCvpF/xk2YWER96oIRAs4kt6L5kG7vFubfCirx7mayqjY8nCC+3
z6By2qVIF98ocnB0mGZkpfq2EW1XNVPyU6+bLu098D+Tj65IC+0UMa7GwLyza1oWYsub7YDl+gpE
Kz3x+fejTbImTX7LpOcm6WrqDpCl32zCUWpm4aJxqiKkKSlsqWT1X01agZAy8zfPH4kgRrXe8bTQ
SBtfwPNHsbGs8S84/0COryZ6MVAZbwha0ifw6odi7D3a+Q2iMC7KJ5w59zsw8YTfcxhsr+n2s4Db
aswU17KbjA1evvv8fsDW4BwdcSUVNYd3Oapx48uEsi1ukX9AIq0aNuPmFAh+fI+6+7LlMSLiTSum
He+ez6Z9sE9n+ZqOLk5VItaxX4d5NkMhK7ibdiAE8n1rxdQkvQup4xHtichb0Ss1fl0lDv63sTDs
E8jzY86+XWW0qSCf5iuU31jv5K+EQ5qHS3mimgnwq5AMHCoBH5h1HHZUqsBfG8NFEzVRoVRC/STM
/7tgUAZ0Hrd0ND6mxZaSPeg67RzObscevTh0o8LYxnZuNyVx+jcoMjGOe+x1XfFF7QDqoGII2SjE
jHJvqwLhLWEjUuGTDvAmO7q3tqVU1o7yhVsWKHwhXQVR+rMBecwlJpToEVOVKPhnEP7VJ2HvnmZG
nS9jRVz897ekSaujVf3l3nnb7Y2CRxGnolj6m/jdZQqPPBDEhtYSQ7bmUcVmSa14+XogZZaXnXEl
8zZyuynCIIO9gkWeoTeu/po9W6grgrC/Jr4VEV1dq02lcZ55QZPmDfVpb9/o9kL7JEOM5sT0+m2Y
xBqcUtcJ55v2i0XUgQNuzsBNsWFZrhX3NTmju8xvXurOSwhluFQW4Qs88LajK7x3TwamV3R7BTyE
GDIj1MK2pefIr2yeQn2GYKaA5qzuv+47AmBSEL/tVlWvZM3g7Rd8VYpXz4f14nnx4O/I21gXaW5r
uQAv77ovGaDXHz0Vu7k11g9t2DHFaUao+90lvvc8TBrpDGzCNzFw0RDbrVBCvoSnXklfLBkbWh39
BST9omDy2QRTj79zQMCHwaGZW8O3hzYLiWrDvvxRO94NBIJmJSuOJlBrmiA9oebqaKtsW/xKZwFN
RF4gUILYO0fq/td/yw2Wnrnt3MHdVcTgQKewTcSMFZELo+uy8xLPErIQ1JX3HwRoxjACWAdTtZ6t
6648XeZiOODKsXbA0C8e99aN+zQKhNNxZgZ6ojdQeZhEtiqSp33nGkVtb6Iz/mabijIjTenEPqjW
ovEuvDz21jYm5XOuyxaN4ruaAri9xuzxgdr3DJNH3s6aWhOl3t+/azgz6OpiPeAXwbMVBl6TZy+K
Za6DiJuY8IuP9VUuzB/fm6zVzXl+jZQ8eyOV+NODK0jP0KsXz7kF1injhX2Oq40L79OG8CHYIxGg
mqPdTcDbX96XIxsagW0JNFy9vhgW4lHaCMyfKg4X9Jd0HS1VvCUAqHs342ESoaawIb/3f5OAb5js
3ohtqYxufY+Ml8TChMPyb48qeMRwzJuX9y5xhoyB6ZsbjOzdG4zwxw4wqrYlewPxIthgLz0UJY6J
miv1hq77kteclW7P0sl2qE/TIE/YHSAI7xzU9YSTUm80g3PhC1se0DIKC6nXGIh3zEbsTASaqNU+
7SjOayMY/6qbrZCDvbra1KpGNu70C8Srylt8vXCa+b6LDXy77g0q2Kwpi6XXuF7qWc6f50dCzKfZ
tpSSofBptvixkc52R0T18yqQwo89VeQgG+SfBjDUVSeJFgy5xPnZEaaA5wPjOHRDvpAKTppZgNL0
DJ9yzkDq0SEjRWTTD4rVeMsw9pFmzHluypSxGeANGbomiyk58pKL24PmWXpBXfvj2IdSor73gfsI
WMVygpPN7Zs9eKDGjeW7BmXnbVtrcchysmLjnUEIvXjAsQYcHhQyzu0dNldUXgpviDFDMgDcgDZn
20yMMt76YrgECLV6Fs19nssOqivM78eSyZ3lJcClPHmI2tyYxTJTxgLtbm4R++d427XuoueTHRW1
mj26EeloQCXQBXQbG+G8n2FH9RX2IA8BBOu5Kw41d++xDtSSvtRW6Lg6JWNxgkQzydnDQzz/YKNj
+cyTF9QVg9mGkLrCUhVdUbIN6ud5FYc7AuS6okdEoSmWEdx8QSR17qIp3TRE82gjPda9U6KQ/K/R
JiBnYU81CR7fzY267YtAArwGE11unBZwWc0a17CAk/t6efwEIFIMP6jdYkviTMuM0hZs0qA8Ox0C
zPn9hEwk8+KBN1+ayOy5Vpw5jfwbe6PQDdm6IHeYDNTNMEQeuasWl53/aJ0CzvmV+pucnQtmiCMD
PWKFxmDexNuSiFeGrbbOY42mYLQvmakPCKTOjw2un+liVNO2Z3lhZr+4q2kpvmfQoMb46rNQoBBf
pRYxX704DsDA01w4crb6G+N4sfHcEkWZlLwm4g31BN8M6WyzjTN2KGIkF/wSMDtfpUuQKcOAcR86
03QK1ODSVevfxQ2LX8DXxBBeIxOp/fakRivw4oUgPJD9PImVupTwQxaI7ykr8q8rVNCiE2jP/1/S
xhD3gi8JJy2pWjXWFTbrOiLnT+IzWWSAMg/l4f6C7BAddBO3k9GnXmkS4Rev8WGHLcEPET3aLgKC
nHnD/+0g4TArnb3046USHWr8GJTu2jFY6g/f/oRKMUd1ZHFmFnJri929bzn9QSGoCOtxF7vcQ//7
LWnQ+OMtkMdCYNuUMNTDdDkQbP8uN1LJAjynKbxi1vL5t5NDM41doiAzTdFEzFgKwuvrDJosO7GD
swXL0/oDRKktk64HlW1z02CK2/99Pf5y82igvbW91stCp98ix3PSR/xWuCdA0qIDcnKXUCmZ9Ep/
CFXXJTMm/AxWbhWBsPau7oFgMCLwnbPc395oYoTPpP7l+erYf9AXkqIlPf+Lr3bKhGJNAaPFqbw/
1A2UPXiFa18f20V1KxnuADaBfw9XwfFdRCbuH40qPECdCoVL1C3AvRUgG5vqNg8jEGWy/iAKAPZS
XIxqdPKOv9H4OWhX1FmHqATzTYPysS/Dw4ACICL0tXSKosBljEDBiPVY7es7P8IziotvM8zXL88G
GeKu/Cvd0ZLUkILb7+LDZHWMxkx/Y6H7xvkPdxoNB2B0EKgICfbTXYNJXegY3BlRtxMbYHUDU9v3
LL+FpcfQYWPuMO6k5aGGU4yWSbzpVHCCtLQuQB+AiZDqClU4m4kbdeDg6SJSLW03RrGeenw32T0F
k2Sk1DnnGlfCjJcp34a/FxPodOULzo1UI58PWIokkb6oxjx3g+G5uz+TADGkYu2RO7I1DCYUgfoK
GZkW0SfzEfhV5kVRrBOjaJdSx+7O7rjupnGQLpxr/vvHqcjM2qJnITClpqK1Lp1jr/G3Go4laWd8
FEodUqX7VALo+Ea1panYSPhuG0dxNRZfmIf9rs1ndwsl+huD80xi/2vYZVbJ+2r2eWMZdz37t6rv
eSV0fc4ZRv6ewX/eodxAjxlF9akM8o1dEhvgtppJovxUJymrvRD4JA8W6SbiZPI9hnIGYHnORBmi
83sD+q4nmeJ7PxnQoOTUBGV92/7GRS/8+lTsCgtzjkOPaWTLKfBJlxnMvpQH4xir1Hn1/haBNAYC
MFzOUEHPia5QySqoJegufZVUeDOv7enNGCZhio0pu1hI/Pq1zAblm7YqiEE9/+HnQuktMD2RzSVg
UhqdHMBM9ZbXCO775JCepeyM46tpbew3qwLsB9k/vIu9+4TgayayPWXSdjkNfN8jtjAZFIphmHES
NwW1uyv2/zJQEbu5tLWTPSyecBBB060lHtAubSy9EcIv8oPKxpRtI0xZtX7YCnTt2JzwPgo2PTIL
M5j8z3tYXp0NJAKrbMr9+JsHmRCul7hA+E14ycO2V1r5Jchg0zHJ8banSbZ48rfL6OuQM++kZzvE
1eolYdizffRmRfuI5JlzuD9lAPAhnhZI7SarhnRL+yF7CjpNa7ZQHuDm7z76sPwtioCagiKEr7yS
bSSpAvt97bC5X2p7oACa1PuJIPqe4kvxml6GoYI977TLeeuzLFteiBd6UJtJ0Y4vYgEyz+pnc1K1
BSTJTwV6M2QJaGkxVr0lHli/D7fhXdpBpZb0UDMEVaYucRrHUKJhCdLMoAMZs+duN6WqkgxqIVxg
0dv4ZyxNfvYQJckESwb80EjJns1XXaxZdS+Uz3Yx/tYSONSjqZnivd9fDK3F8IFbVpUm1CL3vJC8
Y/qlck5Mp+R1qN7IdJvTB6MBV/+rts15rc9J+tEQUZ2zRUMqnUXY91C1o0gZaYXcsIbSY+dmD3YE
Z49ckA4zieljUSot5CqjYgVfV1br0bwR5Pm/u6S8HqmSjtOY34cXkuJ23pCFwpalPT00XwPo+eq7
uNh5c2yryhDJtv+jOn9ua+rZPn9zx6WyVYVKnhRfySewnrRW5MgJqCma+0J2k1PR59bYbLMJWZ1b
SzSJq8+W+F+tr/cN/1mn7n6lGaEEG2OEBMcliFf7/GcIfkGlTi/rgtR/b/rOP7A0SKvxC7aGOomx
8VQbMEKXrGRqWplmHHzRkakVcYZPDuiQBQBvKR72gRArC3L+aNxblA3wjzfh1JleXu25wJ2BSzhE
07/UYHZInDosfZUkd315GdOhd7jeLBEF5xOoyjYVwZa1REkbMG6IQ1u6KbubBedCvaBqVlhru195
/RM92sdanLWI3/AYkJRQ4SlB/nYEYb1nxhEztnHcS1/KWi8GNe2dwJFEqq6SUn6DkNzhT9NdcX3X
GuFkEl8cvgYBBIy/UbNVjnB/p99Ob26K39VGlNRSq62gubxdRUmNmtqD8N2AHF8JvC0KCnWuJSqo
EgPG/WVIpNk5JK0I5/pcEBuSZMe12Jnf+KQw9SdCvsneUnZk4bva41o6dSo344q9sjvTnTilahTB
aorPKkiT7Ybi4xeXKZGQg69UpzJYFgSh16db6sh4uPHvmGPGw7oKnqSlx1U6DQVWU3lWABe530XC
hR104Jj0DXWXWBsAUHB/J1GmgfF/TZJwanBH9XY1nXMGTpAM7farOyfsE2cyPcMpj/ldA3hvLwVK
U3XuB9A2mFjYq81eQRQ18BBUvtfu2fulOSwBOASvbUN2UXoPIU8frMLZ5CRb7qJweQi1xscSCx7V
Ww/7vm81Iebkh9daNs96WSfjwgcz5jkME1s1OJ5M7PqPp2ib5j7GFR9zTGcs7VxFC09qj2E8p3u4
FL3LRXwd4LD0I+S5ySZ9sfFVXyHANOXNEgz2MdTW+8vAY0kzXZOQit1NEYcSxfGp+G7j5+bIO81R
70DArQZabtH8yqbNf8C6MuQZfNiWxV4GFH+BoCULIiu6Ygc2D7jW64f2TGhWHU70pG2KIllHUyb2
YaXREvUWpbNt2gpL+moN7ygWK2s3aNttqtCBS7KR9joFD3ziRuuvbum2YRtVYtPzJJlyln2O5pFj
F2YXzwvY3QwccxWwrzUFe1cbqBB+Uj/5B3aQhZ/n8YxyqqXVcePGthbLxDnfPkvOxkFnZTuBzj4r
m0kz5SP0ovfEN5RtGYxwPpJrUhseHPRbpp84lfWrDP/5tsKPJBCzm0v1ww7vlpVZ/r4rxNkbHdU4
HGTEvmXHXe9qPK3zcv49WKCeZqrE37yQE0SP+w9rtgaipNrqe6wKB2aVcQLfksSQwNGu3oKLt3vC
h+kEGkqZHUwkbuEx9wN1U4fHG3BzDKk8r13Il5tLpdf2Odso5O0QQy8ECSdGmJQKGzw+xaFvTeyl
tnMjIVcrn3CQdqfRRAOz9hkVzFpjWS/SQaQR1o+Mwaq5jLDULXGhH+f5O/w/WirTWwmXsVp+j4V2
xi4g0mAEr0B5qmhYPVcze3NoMo/fKHdSX3hvuFIk3OJQKo6sxDznHFxPwlqnhjdmvysVyR0UlO3j
6wtfuF9lnyZTPZzshZnDlkKF6ES1xxLuKJXbV7+jJxTqoS3E92fEg6iW+wLj3DrXsSNFGW2t+nPF
HR1HpuCdLEFze2f322i1oJfSjN81MOHIRLpXb9D7DfaSyTMIW8DboitvBN8saY8JzaMeYTAI3e8u
LoPna8MGD387zy4VVzRK8fdsYwkDJ6hYaubZ+3BKTYHj2ZPTgbOhRftV97jkHGIEvH9WYC83hnW4
MEzsbm8N22EwQbW5UtJaOlxWVDFqkihZxxkK+7PzmzKBudHIBZPLqB44wVNov+dJwWI1MUx+rHmZ
zlFHJgNCTNFKlXWBuvNBFuvH3izqkeby/1v78uU9QYwGikkyxkuvXtCAyKApFUkJOT/J6ZwOluOb
eBfYt2ML6JfQEiCkT1P5wyytEcnyaA5Qlxgw6HC2SOfMZxmcc4kESNtyxtem3qaspWKqHZ1jlz7f
dXlF9lVqpAGey6UfwLrtAj8EMrXe8l8B4rzAjxQZe4DmPL3KvDbYhWa4minP88oEBWg4Bvi3ezlh
HeIc+zR6+E66gNc/2Ox2NQGsWWOjaxTEgZ6PhHGidUg0mjhsUl384+xZTZwHaU9v6AIE7q659xGV
ShI5x/5DsyL9Hn6a7L0R3M0Dc+4lbG5BIgadmPIDoXNaifBwNKnhFlUIn8kd1L2/Q818/ItfliWN
HrK9kj1t6AEDl9qEv2W0Vp/sa5AQZtFO24mTgFIVJK7AJN8cqgpnGHN5/+DlUJxbqd1gC+6g7JPj
w1rpsPDCIVWgcsUMkoBIP61weoYpf0WvZZ7mxDh/pzf+aQmEGp/fspjOD4tBpLBxyntYAEBZSL1Q
dtISQnHDlSmJMXrJANnPqIHHL8cvLOOUrzWaQIhBv5KlOkCu5RJ1DG9NwH+odvKqohlPp4tkK/tw
ymeqNPYsvOXeoYea+LhFZGGNcvwQeCE6PcqhrSLD2lp21tZkUucg6WXh3AjdcxB4rBlv0+Sna8GO
ergbFpSVDGT6A8S8okaOnt9lZ86GwQupufCPY/57itY2KFZe6Avw2aOVDwVcUHo9MTBxatIhoEh6
pie7wZs+zG+G6txJmUtJo/ifJlA9p0sl2PKFF8huVEvKA5QMVJswAMBVKEGudR/cXAD2zN4KyCsq
FVOrJT84f9ZtgYRcL3frFU8oVYr8jFMCG19klwgG3NZdSRrvTlDZGMv63GQAhHlSLRWmQIUd0riS
ND+EP8tUDkz8rY4UcFEl9xlvpoMAeSX71VJdOixokTBlWkcaAQQYS3Vab06DrLz9gG1ZI9FDn4gs
p0mwJqxg4eKVnVYrYLEq+13/0qBHvdN6TSJxrw0MILZTUB2fvDVc2cRCGoiWIAY77qagCr88lN2U
D44qMNm8xPTTyWHrUfrAz5MGjK9MZPvXM1m34Gi6K6VWmZyAsC7uoat/xd6X8J7KzvW6uB3lhSPz
1eScT/gJakmHcrlljwNC1vbU2To2bgOIJ/UXl3xUh4Dyua6lxmWcBASGy9EZg/sK9vX5ggck50Ix
l4dXrTeR/z3yVC+yMEFQoYVEl58Ta0cprv1Or5fNmiI70jdPJIZOcrUMJZ3T9y3RCwHQKx/brUa/
6Snmpyk0ezmVd/ctXO8sRmkhqEvuGnr9HRS3YVtwGACDXUD5GnuuLs+VV3mvCcAvYLyN1Dlon4vr
s8eR3Jj85/cLPX0b2SyopTepa7Wewr86F25MomcA37OMDtimOvyLvwy0kaFDqdb/5N4sID2ewyoq
b4P7R4XkKkHlJVcI/V62nBTwqPVzwKGhRHBYYwwM5hFcD3Cv+W04a1jwkdufzWWKNnLngpvFIqt5
rt7QMdCV5D9VWQ9BvkvxDliBFaIhVQh985No+3tmzyQ2FaJteH3fBJ+wwg6JFyKIhC1IUgImXFhz
3GsoMq7+D7KBJVHTlG91TtbGDpwoi1iMsqUS7Jk48giGkwOZgzyWyCWT7pTLYKcUoMyUIp2Znqpd
IlZsQoYN8kYRJHNUJU3jQaNfu/K33zIQ8clsr/jfSAd3yd1SxJ4wyIeGP4usiBeCBKP3bDfpiTgF
x2a6G/oZfkZXvYCfTx83L9Yd6q//SBkVfDYyM0zg/BJq2Ro5PywOPZ/Zlrv74ipJpyeevlD4tXQi
HnayaPINVKMDIQDMz+1VwMs5K2BUDFf/yDqIFAoz43i0ft/7rmAg4o11aqk8nNKwxvzcVc4TKT/0
Aooc2Wmxs5WO7LwlSfyfMyWfyY8IFVrbtL03HtiU64fd4NfJY3H2Hq+mFhDyhAzclGFnzGWmKISA
8VQDJYxx2s1JaXdlIceIxPG7+z4TK3G80YCN3KkK846Am/Di7F6a+oZuy+BkZ/AUdHK9irAG0zXq
2ofmT7KZqggKEFdOkDsqz31GhkrxiImd7pzGr9uYBXO3XR2iZuY2y4aCzQYPpnSxeKtNISeza1tU
W+881pxoBKl18ZnTMjtFU+KCIShl7PlIrs+VpujApoL0Kn3M42j4sjhKAVJa502Ni8b6kVCh1rwY
rQGPIcG4Bs/rEYBZ498RWR+3uBrTSUHaHZzyZ118uUUWA9N5C5Y3W6O+2Eq6f4eww8wKz0ZOYCt7
4aRtaFlAOYq6sE8BIYej+gCjzlHRH6gSvuJH+0PiQps0zEGPGKmpEFWShWqqwCkEKreqvz3hgq80
+NInlP+CetkdBLd7rKnReFuBY22XqkJdFIQ2nTlzFO7zEzA/NLc1Zi4Dv3yzBwqADogak5yYCWni
qm9CtIpYCoUA1W2y/DZOzoBHOFLl6mKd1vdiTVGZueIVp/xUsqn7+vn129+6pAWn+kxecyiEb1L+
qGae3HQbSsxRL2Bsop8vr5xjJNsYBw8ZD9yOrU5DI5EqxqJrntBy+YvvcBRbkVIh7TJwjSvmWkYr
vV8zGh+n/u7vgE7aHNqeRHCl14OfC774w/Jc+tzb+VkPwy2MlX/jA8Sz8jfV7d05p9RO/Ab4xuf4
pSmNSeWkKN6oONfT3tPIPItAhjtrMsKaoPrOSJCDXiZLzKUVxSH2Z4zAQMaGUEZLIT3vJ/kHb270
p4PLcgvH0jqLZZAgW+voigHkduOv3QMIqzD2ImZWYbsWzLg6bWyIn09m9j/2Sfw77QYPZn9YKMo7
t8NSMuy4XFJdEFh9Qs8x/ZlaYKNzgUj8pVfka8GVktR/SKfBk3ZGmwfqhX9DBCaF+wHbesktzD/B
00HPUQe/IIbCdU1vpYI+MxpFuBDkNghgWmWU6sMZs7KrnE7S4xagwz1lIDKRQlk0gXwsFy5BrhWY
3A53l71Hl0jNx1e5XZo7QnuKrVSOXRPalJJlO9AtpXChpnquHRhCKI/hjyr2W9/loshCq2UkZSo9
9h2SwMWgyhfnux6VOFokehGOqsTX7ughtta6YBu0KRqiy1jx4XZ91hqysaWWRaPne2RIuD9w0SVv
dQ00pe9BSYXuk0X98dd5oujLYldPc3oeAfsMX4vSw/6guoW0veQKOtBDZ4E6u9+Xed83Js0U0wh6
4LcPEL/4kA9sqvu4vnZJCJfFcP1muCU9u/jGxP6VbVw4zhiuKMMG0y18qKPAB9bJ/DzK8wql+Che
syTBrPg6G0K6vX5tP7Nz29pprpovAS07Wnqqpc1lUJu/EKIIiILNJ9JJWxQYkljuKIqtTiJsU2+W
AB9qug/1UkqVSvGvAG0h5G6q2WucN900x8jfA4kFBI+nhOTWm6pAFSGUVoEr7ebD0xWeuv1q9Z74
Thl4cnT9RfWhuUZ8JMVEPHa17dKfLHYMWmJtsvGWYenDOpPDZR7sHhqtlJuEysIeBAJp4Wg2zC0a
5vHb2UT4fko8pEK+R6Vlm0oTpz6prjV+sCKLxhPAal4WgCZ03ZE47TNLMxNEE2ZhNx2ujFH4P77z
fuZNELGK+5/h0bBSAqaTmtTt5Yd54brd0qbK4wkLfnN3s+R7F7mMEbDEKmjkDbA2+x4Mn8ESM2Ne
dmGzdKi4tcmrMo0AmV1b+s8hFwq+Fzw0iSrSSNzZwWIunowoC0QOV8vUARw8bNUJUHs3oiPUmTwk
DNfd+tQI53xfwFESbb+p+xETD7DRCUVqnRVTdZbohlGee9cmfGShOzvE4Hkk/czurClW1p+OFju2
cnu5VArV02yelYvauC5dq33dn0EOeWwlft2zF86qRiKSsLfRetoBWLhx8U0KJojV5hG5tX2I54zK
sX8ivzQHKy/o60xBu3YbrUR24BbwT6YIUxlUglDpZFwYKR+mu7qeRAzCezTuxZw0kghfgEdSqHUL
sQ4z+x88KwOv5V/EbZstgpkq8StEtP/6yiu12lF4c0DLVZsaQ7utC6YXeyS0MMpIJMAfUU9k2Clf
yIaqMgKR8s9ltm72+ic5wOoCHR637HIJeQ7r2TlQVxtatfW0IycEwTCZVe5K0Mu/e6W3NWfxedn4
X+0+G4qRUzLspKEwNKc9zjhtKhpvwxVK8C/vA8oRBkdQTf9DnAkduk7GH2t5NN8Q0yo28tzEkrmu
bYk9Q6MzIB+srOV5JrQU4cZJGsEF3vRQD/wW7cnOJnKVTA7PreCajk628nlYiUcxP+wUAHfKkKkE
UTZR6rS8UZfh2sgjR7Hym+f43hN9Wi9jR4mwLm6ll2fIg623hac6xF9PCsxqa2G0GJGpXGRPed9t
u2g7hoHdZMho1f/1/bog3UO11HF1Wt16cTwuaurvco6rv/rOfRd7YiocKvX8nE+yaY/czM4lT3jb
CL+DDqdTIZDmnMm2xWJYenYjJK1iimLOMdjGFC0fVUaA2n8FIImTQMSaqfNuFoJsDjdo620xuWIK
rpWH8gcTOjnjR/V5/784uMDiHd2gJ3NV4MfWquRL4B/CEjzdWCsZT6tmOUr2XJWLOAIt8vBFGtHN
2x00ysYpGC0/gmA0bkDehmenH+1xxf9ujBNPwKIePG73Os/5IeIvBPy1wFbSFAKJwSvUYK9iL3bj
BFOBsoIz62fowlXyZ9yHl6gkUcTERtiKFSX3IxnlNZBWbigqPv4h1oxl5ZpluHmia5dQhRwOrAXt
d6nTZN849WEh489e1lWxgoBWFMv6XvyAVT5GZ1eQkIeYi9BtnzkazOtbYT+KThGwt7S94hXCGZ+n
9RdfvzOP4W115yIRtrk9BFLYDTWcrtgSkWE7eSeJ7iIsaAXyP0e9FRJQRf5NivUr67qgEdYH2jF7
I2VnWeAldBjXYhJb7Yf28nx0ov7QivY7gQMgyn24q4NH5AktVoJD4Mt0wOrwcAKsGBZ4yBZeGetD
3EexPTv61x9HK25bKorbDIHxfyZ90GElfmtnNoajzDWSlbXlbXiLheW3J7Gscpr5B0ii65NK0+8/
b7uKV8XOEl8Ogk/ff8eUBNTyki9ue/nUZ4DxueAfhxC3eFzD5aHoSaTm7cZ61WXS3iH8uaiaLCUf
AGdYiblz5uxdM4m5pLwu5eQVF0KYufkianOs2fFwc5UP7JPiEK48ub6p56eExGJyYVsyR2HIYOSu
hB9oepSx2jQNongxnpg/xxzmeb13R1UXMm9fhj0UUAgpZ1v0OQIX2OPlQcn5h2MjmhbWomgDeSWc
XmezS14THiY+Tq6TTPvIhTm/ZXuGVUyeMXSm4Iz1BoAjCNetf+vWEz+6H4We9pSK8+i9j6k+Sv81
zbFLdP1jSz5aYoHhuB9ECQs27Fo0zPUirdOOfYY2VxUI2IqLVdTpFx5D/7ZQVJB4o7joDeZ4/5yS
pSBmu/m7W5Wcd5JxA6NSwfOgymZDtwbK83mJZWV2d7WpTZnflg2tI5nGCoSpWJyzKnon/5yk5zmK
HL6fzPjuahU/M+Twqy25Ud4fsS1OBpJw8m68KpeuTkwNu5KBLOsD80O69BHD8ifnzVzxkeKxHC/2
yLAuf65RtO2QrsuNENIxg8UytksKbEwjxJI8ZqJiC+XIfcbaqFATFO9tujgUgUNdemnIJmGAgecT
1jtYb7CNxVhUSob8lcFhabnWKTQXQyIquikyNifyDDPTrTGUucOD0s+jj3e3Z8weQuZNmewxvYDX
KAo7wpvVQkTF69tIsF9byi/HNlDWa0l/LEsLFl5a7YjdkGlS61z1gBxoLny4bBGEGi44dN0/lnJ0
ED22FNfJBylPU0t3wZ9340bNvavpFOmOnryRnz1I3C83hTI4hBbqmv992cHdVxXJ0ZER5RflwY8w
pwh2mlsbLex3GiTIhHe6hGbRvIWVAxuECVMf2mCL7BWBLjP8svYL10pbA1Vobabo2tQ7aGQuv7EA
HfI5r0aCklK0675ldJ9neC2LONQdPcXTApG/FuZhDAFUaiGEzAuO559cGV4B/oLotQH86cnvSyck
oYenw0m9658W+nJRMtWy3aXYE337vOKkbydUYJjIGF8PNrFERGj/8Thdtr+/kM39x9qa9GdfdKzN
cIqmEveF+0e7UxoZtTBXf66QYsaivzCYfNmoKzM4cDD/QGzMocEAaZnBuuJIsJdiyt5gkmZZPihY
I55PNhUUfSA2eH/K7T9LT3r1YTv/cnGJ19/cEsfmFgmkosIbcP35g5B3NURu2MKub9m7F3mLBk8W
yuqZtfkOpiPWreR3IG0pJ1ON2fGRnQJFPYwfLhpkktZMGb+2aXwKbRon74qPmVCisXSxRQQGAtBE
8KbBY8rcm85WX7UvjtAUdqtfHOR3hYSr/xLsFgkpjLcTl2BwdMb9Pu+fnOkZdoj8XMOIIJ2Lr05H
padtJSKjE4R3QyI+PkmfsYdigT8Nt6vM1rsE47eR4bZ1+wsn5dvO26ExejP/OE0FoChCG0xAnu+a
Ru6E6w/vUEDJp5aAVvwAo0E4lX5qWqug2OawicMnneQdQ8SSZMnvkZmQ9mg967WWVLYa6GVPxxqF
fIcBIu+dFltWlb4uAXJR0eGqY2DlvXCINSt411Vz2MTiWjDHw5qCbes/+VHScBbvfAee43JAEnA5
rEBi84GkQ+w56ejV3Wbk4rvm0YgBGUUvgT2bgGHEVomWmzQwyYMYalfG6QUDmls7KUJ+jzWlU78f
WWKlHm+OD84RCqtaHJroVSGnh9UQaC/KW/3epsxuJJupsyGoHgXSGDQB0YoyWGyq3TXSGg6WriEs
rpkRyp0mOMzh/y65Pfz68H2tJTSglrz1nmNi338W8lWNIMYVF6Ox46d9T/pQLgQJqN0X5sk86+Wb
VGKsmCR2DGHwE1McrouvPWaxjaue19mhd4IS4h35ISgpRrfpQ3mAzUMSbacA7dhpuhZo30Q/kyF0
ApGG/86KBLZGbnrhLuuItVKip+BtjuxT0X7KO+wlsdkMcchlkjo90HgG3wF8F9yRsno30M8APIO0
aD3RGWxpBXs42Ps23EVCQOc4A/bzjzKYi0x3zoovwvyxQwIqskFwiw0aq5+05zkHZXEa7yLjp4Zw
EphIzhVLPtHIAv5a9AGa73cVFm6XQxmij9jIagh1W4EFBhkqnscP7T425JE53rlFNfhptJQuvfrC
QEemawHVXYYpMO3pVt/qDza5U8qbepWU9PvYQAhwokylIUPEUccNIAYGs44L+2hz2v+kdS9Lk7+/
MS2EmCQT0f5yPyAehfv2qdSah9UAVssH+JSkpUCg2DyfRL/kVbzuGruhsAakyLPXExPvuwKPxj7l
MdtWgtv7OoZ8fe9b6L/Equgrp8Lv0Y5Nzdpj0UDh/o4iEtGDEPErDaDBqwD6/55m3vFIJ1lss6j+
QZMquwg16jhhE4Dv3gste5CX7W9404jmN9+8L12X5ew/QxB7dqtfIpQJGW5OsrVGgCJ9uwkf37V2
LGHkKPUpu9GQ9BiQDMOA+5+9t9+jQXjT5W6EHjLCEH+wfojg7WgkIRzBSsaNDxlW0RTYelFgl1Kr
0HzzrATxsSdYWvzm15QWBTWM/RH5dbUuNE4GvXUWF3OqIEvKagRCJaPyDe3noSmlt35PMSgDUqUr
kzkUTciCy2J6cPx2WgtdJUfCeBkEYJfKcJdzrn+V3XIJLtINCiilrWcFJK7lWzrAqKXbyz2MXmwq
lZv4cNJ2YWTv/brUnMOCS5KkIdAr39IB5e0A4vtFx3MVhaCKlnuZebdtPfbPGQFKkYnSO2baw/y9
YaDfwBMp4wmWs/8fhxl7geo9gk4PgczOsPg4zx6WL5qgakAADWFLEEze8Q1f1cKzhQ0Zjl/UkOZK
B+0Z39PIzR6J2m3a04cJ/fgtYu26ThXvJIBGPkCXwzF0GzL+UDmQ9txEqGHXtot6CL5LsZcJdJ/W
PVkQ6Yx4tXkWMR9hM1YiriL29bEQTJLv1rbMh8M0WPJnIr0dxaRaoXRRvC4TnnZeKMSXMD0SXjwe
f5xDwIW+j1IhoKXNHp8QSDx8L0whJI4hEXkAA8/+5Rp3AQNAvMqwjj85bXTgOt6ofOHo+tkkd+Sy
c4wiudQPBgpk8JgHw0umZgr9d6I9gc7/DLtMqA2i6VbCVqytvyGyZWmRd+0GOIqH03kvxQcfcpGU
M+OoVNe0WioJkNAWxBwVabRd2gy+t9wV7Ov/aevD6r4AbUJMKopjD7m4P2PEyNtyW9CVecMhcsVe
bYZBKArOvls8JtzKYO1ewVQnEeWMKvvROZc7SxkoUgwtSW7QNbwQgsbG2yjuGZju0p68azPkZq2n
kI5zOBOXdWpOinnIFnGKbAgg8dUDcRftEKawpNGV2kCN9ULF0WmyZByD3wCiB7HZm+Gm9ALXWMmy
tZpb7DDHfzi2mf4LqxOabpJkvqwnuTU8HSm7gbv4I9Ku3VnU3nm5qJn8fem7mHnvFENrAjskquvr
nW4mu797I+pPe4RE5S6PFvH/MwSXKcRCp3hsSvtZvT2GljZrmrvDME8Cdcw89p+K1G7xCe/YKFvs
KOyyAlQgxGMQMtWwxj2J2NQ7aFwqUJUfK4jwSqBGZy4wS/Qf4B8R6iFIZBIWFIA9vXWkpCKYksOc
vjhJabxfJpU1AYeei6YPpF9alR2d26c0wI2QHkT5CKomm901i24Q5j+c0stnoUXpYs/fMiPmkDBc
HXaJG7EOAqsqgUf/3QO1Tk75m8lS/NaxKMPcuIPzDegx7iDznLbEmDnbBTidXcCNuuY7AOBzZnkr
OeOyJaNUgkR8bXY2bb7iGwJdp9wEw9iyw38JDz0xyzwfthChpJfr90y6jxCFs6rsHlIphDvZqeCY
6nneHM7CqSQFWCOlBYkwdVZxacItYx4rQ71GKqtfBfD3YZoTXnx7ceCKhL5w/vLDPwCTuxXIREo2
L11s1EdxD8tJ5Z+cSPaajGcia3apZlwesLBZ2ipRARS23/F3UuQYvnwsIYsZS1eLkiPND6IXtXrJ
8oXbtZ2I+I6zUWVQaMIJ7lQjooKvBsEIzD6PmEZRA9NAkl4ZeOVAOFMX3L+lERpO6saCVFFBADW3
1ERqrOrKWoo9PupL3VX/olHcNxIWwr5AX9xeJyfmI9R1Yy072MGy8YXWW0ub0x15cxSoJQ/pucpW
ukgsKOR4frhpa95oeP1OgaG+df3LlZd7vH/9YlZBjhz3OE48sxI3bPoG/gE/hsJNirIVCy2BjSRm
RB22xc4RfDampyD0JVp96oLfjKXQamryzm8ffWAUFF0HDJagw03kyn0zUYl/1a9Au3EF+0bJtPzL
K6H8kLwLQOsgMRPNlNE8dntq7imkFWOypvnuaKgxjt/+nnOErRgn/gxdPM1wR7PYbU2Eoj+wax1i
jZAM0pkm8zBDwJ4Luo50dlmd3nojnGiXOkT+XFi7HdTVsU5XylPhzIdhyDQLyEw0Lj2Op4pImWeM
MIH7y/QYJv+uoz8mFIJdhP7L+fdsMGZMyJLM56YhM6QuisjMsNjyNGT0UGyrR8yovxLE1mXGNR3/
jbYzpMV2yyqydLodl4Y5QDXpzkmp2juFtoy3z4EqtiNC3pwG9dus0O/dE7Wjy2LRGD6c0xACeYQq
tFTqdEsEjaNAAi0H3Uu5UDtTRzpAxxFW67c/dKi+HzYJL+Ylkgn8Ail/VrCGJV+oGc5NEoj9WEOL
4ckGs4t11atsdxiwOUEYDaOJ66kG//ixf/TaBw8OOk1HoiQHzgyvkJDSKb1UXpjTBPqmGFyX5KlB
xpzcrvYj00QR9GxIQKHSEgJTRNLJ5GSvxU1yXbEjAsrM7EEiEl9Tszr2SPj7RhbWU8FGou1dEhoU
jjH2Dy9HmF/OdG8vpOQiSOxKYGNdx/LzH3tiMkTg9V0wNx7mvcm4ksbQ7U/jb2+2fFLnpPdfwG+o
B4PnNJ2qx3yKhve9DtZo1XnPdaBj8tnchQfJaVTNV1oQjpbOL3JoPG+KZaqFytbgHlC3I+eSS1vq
6lQNmF074eLIwu/+5PgGN8kw70Rcn19JK1r/Za1ahc8fu46QksKnKZEzdORuTOuz99DI5QxfG2RN
U41XBbQSJIX5+PlUXLOofT5Ha+ImiY1/VrerHcn34oV5XNO5S6FwGv1zK5dq/zISsm13dWzvy1es
ZnMP6cGA6oWNRPV51CjaDikZVnaX7lIHgbWo7fvXrFHYZaiFYHORpc9SgqGCOjweZiuWbyzhASxa
s4jquzkOnV12QTUL8iFyAXiSrzKuk2uugnDYiFeDup75O5wBEiMJnZ02G767GccdEa0csZ0vpn3t
/4iUKtfkS24D9Defs4/nAZJPsCSO6ZQdOJ87I6Fbcy77HGxuTZsis5pWLSo3xFmpVzfMjRa9HUBW
LXNzbZN9f/v+8XUY+pKPFMrTs5vrCF691quH/3wiS//Qn5f+7Vl/2Xx1ksv8g7vJ7U7B2OWEy8i7
WYGI5qLPn/SF/5u8OWPEshljoPnvDgHHUFomlS0r+wMMNNsFQLNKAQrcxMAi5mAE0gTS3BZPBYdc
ca/xaFsq0jN0q4INUGzqFiyvrVQgg194lf0JUcaGbLSLSFDcz3Tcqi6cp324iiOIR2+5canuO9ED
/YjVwcdNuW7Rp8gT/WStWvV9AfazZHPn3RpyaER6vQ+91yXDDD1Q7wv+hfNMVEmLmgvnRCL0ddBD
VcHMcN9ZWl1S66sr3U2YuyWpI2r2uYpFyz4/pXrmTOloXZs/WjrjRRgw29D2vhsqxqEc76IEDoVr
1aciSnw7WAJe/rNk6UwFAXvvgzP2BzT/u6Dm+rjCLt0X9a4n/E7Dl6CGW2l1MX9bM+vCEo38ZNBx
yo42HZuyDTBNftkHUEMVp8SApLV1QE8WqgkWftPjkqKrRHHIKB7VXzAG0zRU6WlXrORNgotxECcF
EFuqX6RICqhoYfl0Z0T22FO33GArugcMQSJ/ohb8YBMSS2J84h/FN3JE/WvDslDrl9nboRrGGhUq
UfI0dSQfBBRqMMa2+3t7h0mo4RacARWGQTQmTPpmWBSR0gFnvcElEPTAbHQwN09owUhqpeE1EdEC
RESnbOwip/4LS1uvME43UH8JQFvsYOTHfT3ETuwVTu2qFFc4JOgBbp4JOK/FY93zA4zhjWnzhwUq
m4A2K5bj5AjBzwWz4tBfweUXqEh4UnWJnn87uJV9geUXeDZ6FFQ4f8n/J8uunoiyHRviJsbhIVMs
lsvNYOsMnvYcGJro8078KFVBIdR63QhQ84rZXnl1kaa7JyisstaC7Ny5taemD0aKnrSxA0FYPBQv
n4GKdTEJsHQ4wK5xTfGV8aa0141+Z/wkcXKcaZltvJAdNiypx5a0gYzmNGiG1UrHYPq5AtIxQiSw
B+1IR4Z1BcYnS1ENkpWQ7FP/ZmTHv1NiqogBwLQLqtSYXsluXr0A3dcH9dQObohFHXAquuhZtYTV
92KbF/2eZV2A1pUUJijv/3Btf387cA/NrmBKiXBcvErLw5FVL5e8aS5b0of30IlWJAnFG3mx1TZk
a3q+1Kg78pYeTXoNK2CCaqvJGVIsx9TzazVSZuR1VNEJRUweNJPY1UPfBkFasm0Q77xLA0rN2ICS
XBYIZoqyQ4s8sQr0+2QUBvh/hHtNxm65w9RCJnGH+t/UmDSZvoucuxmCpDEDXsKQzoDDJkr3PktV
8QBmCldyEDqvJXQ0R94foXu21rEuVt7Tf2oaYTjuZZoscixgH3h+duNgQmrIDUS8vpJYoBoGsjSv
Vdf5D6a1EDIWnpI1jaoIz1e3hdhoAUPDUtdkSoXLkPziUiNsZyjONcofCM5V6GqlPF+XbpyNNl64
Spgfrti5n8NrwGpS4yfOvuuVgbK/3ywobgb2DdTHkRc5cf/sO+wYwk4ZlLiT7zmQDKlkots8enil
Yzt9140TbjVdIhyryBHTKbFL8S70cA05UPy3jKhGbdfs7ACZZOAM/gAtCsu/LNhEeOYDkZojf5Gs
1lcvWoZ70Hjk6nxJBbuE6RYpM4jI9qNJawr71dRVWDzaSv8tkdzysu6/4pSfztC0jifp7tSGwg/8
o2gA0emrdBu/sb8ycEUYd9oTHBr8zO91sapmJaJjJL+3z8IRP/Gv8I1moPP/zHGmy/sBsRSYo1LR
PfzH6/Y1ThfFSDIs1k8tNBG0NlRe/P3aqxofj0vCwTLou8ukUGBH3aXV6QNjoGLstRBoVPKLDtc5
tpYeFE7jmP+6snUzcpzmX7DVRkukeaZb7Ph0iAjlgX/2UFx/+WIcBVjV1p/ybP8Ely8WSDDCnMFB
oWtENCeQUGw2SUi6NL8zQVUOV2h0guAD64LGMM5Hm1Jhh5fIGbJycPzQc+8YwvdannUlEEhg53Md
macz3fMwt87/iEE3YfWTonsasUiwvwLED0maJt73B6uyl2VZUZRpJG17lqM70vXLextSl60AZHs8
E4++eggC2jSrdOPvj09TfQpykcKIG7fLLV8wq5ej1bF3rBqxXohLRYXIdXwUFbT72b6e5syZH9Kf
XwYh1lw0/Jl4nBb3G+Y+eUEKR0Zv5be9EkFL+jCbTxiZmZptttdrCBWFkp6XgwAh9RbRXvm9wuoK
usRhsu+4ihPGUvz5E9ttOYt0SDnzTYp9LGL+wD7Ezmmp8MED3rr+v6Uk9GGMQCIJDAfz0ViM7fqH
h0kSfdjQHzpSA/mAYQK2sSMurRUFWT/Ym5PHkQX4fOKSGMXzQLUE3whBYX8g4zfeMlYBNFNUls7N
kfwArGkMwNS149gon1MJx6+TfKgSR/r4pW9OR1QiryemDvKXUVZ3X8wTLx3dAP+SjMOLYgZzJwKX
EaXssFs+Zw3pq9JIGexRvjIp9qNQ66jb49vkIEz4rsfq2rVgEO6+UsZzb2LqeoAhR76M8RZsrzLZ
JG4Po18XnAb3DOA1OkvwzwZO058pmUYwrboZ5WA2Sv2auof6D2RkvGo0oVH6+CTct1upoyjCQNX2
2LSlbAJrRdHrcvIteCzB0DmG9tCI8Vgom7rA6LA9JfCgcXloFP+E97xELNjBUYkHvaOu0dI+S6+9
Bmt202n8Xb6+wzVjiT7iZhYWKR1kTvx/QPH5oMSDQKltB2H53gfPI2xhL07qzIIBwT/gj6Z17B9+
GCKAYffvRDM9eb4wqSAfab8OHYtbp3jMGPGf3NkYhPimamUFh04RKdvrm2z/o8gdVmSz14KwvE+v
YIz8KlSkep8vsQeW8eTo9w7xakZoyue9WUEcbAE5Y9H8zOEQDJkxWW9LxqA9NmUX5Y4m21tEwEYh
HVK6zpidqhk+Vkj4UO7ESrOrVZR0aQMVFNvaUiCjvG83ZdDs2nOzgQTE6dfatJxL6JdOJyB62m0V
/MPbqhVIWf70JNSwTpLFWOOp/a33JCo7MDRdZnHfvBP0E+GXChE7crpS9SGIcTVqUpH8HwOPHH1d
MdKSe9M9Bttz/g51omKvVdYkO+M4b9DRP5xkkCTGeK1PwKHrtiP2wibKKVhj57xfuzdNCnZ0SHXx
PjQJtCwiNUc/6w5MAAgwhEe/5ctHWesmNxKOYEbqSlikbY2UU4ugP7UATJEJxCCSv4SZW5Oy2Whx
cPgKwP91FbBhHxmjgStRLynvRK7Fe98Is2RzDS168sKGkv2MJWq4WFpiWDOMoacqC+kEG3PdkFoA
wpR5GNsNLiC+IrLTj9kf5lEQWgQpQKs2gdnqzh5GEt5ezeCMKWdgmTL+SIbJPL9yCQWQBVEp55qa
tGFFidcwV2RRG3o7U9CxTn9PFSpdSnTifVEbDVJCNodI/j7gEmEiHHQ2Lxk51oFtoXfvMlDS9Fro
dcf6c9sS3SMjpevIfhWW38ipkGEBdt3RFhgPpmonlJ2VnegtmG+M1eVA5adDInWrOcYVrUv4fcOO
2qIKFW6+Ina4KjxN3+v8ozbaOJhKZ5CnAJD614V1DYbFGKONAFU/EltUABRVG8f71czFJCWqAJ57
F3PgZuA26I1ow7il0I422ojNZ/epH1RsGRb5M/4GV1Vgm7ZBBEnIwsZM+rCjXqjhFqd2htjEjMaN
8x9Dzvkh9+F4iVSEIUrBYki4ex5g+G1dSl/O1jKXGCsHAOdK7iRZt5SuX7vwbvCC0WvZe+PafXUP
OMAW7sCJJLnJm6b2HowPMDS/EpNAeHy6c0pv2cw+gmhIwkMhWXEJ7JsesUZrlRsyqyDxzYwdxuP3
lysWJzLXsgqmkKSAbE0KIE+SbUZQVmyGxkSZp9FYSnFCQYNvMnG+rmk+DcDlrpd88vQrtXSbITDp
ODDjSbO/ifqYdmOKRI2aIOvAxFdI6moDDx/1l3wHzMYETCpN0UPbd4W9Av+s9Z3AEKOtHbUw7WMD
KD5Y3aQRHXiyZRB0iBuN5ogmBgl8F+LcDFRpjc7RUdRq1SMv73K27CnPlcI9jCltUfrW8ljxNoxq
HerUy3axJMkHRY8vZlTsYfNJPOpug6aw6T+Cp9wCEEQZeESi37UUfM7dM2/jygcAzm/Q9jJ1H6S2
qq8rRUeVq4+9d2/0af7FJ6Vpmf7C/cqUIIq5udluzQ6qppZdQgHHY2dn6BTrYQGzsSYTvGKehMjD
bSBySG5B5jynpVy7YvsAf2ZI/+ZADp6XsMRoGMHFFho7qpzyQ9yvlmuZ+QDFbXP8aBPOxanUdaiQ
sXA1SeA6HSs+LSp7PNWsCOzSjhwz5hrtg0tVgliJJgiJjxki1TOmiwAke3XIOwCenvhgTfTCCVIY
u2PnPY283Bby7gc2jlFYwHclAoCXc9G7mW72DDmoniMTLpCximGFBmycFHe0BvwZeOfaSkiiujPg
7yItFEmADi/0tMrjnfXRXgUuX5qy4pUqg2ZGaGCnGR9AnZ9qF0mrFqzcoQxW0W/Mqf93Sa7GFvve
l9aWY85mzRaDNdARl+mphcJb2XgACAtZJRRd0exX/xsaGfmuElk10C0JDkGu3uDQbwUQIvbWACkk
buDJbfsz1PEqUGZUg9lG6lHhezWjQxJ3hBkDm4gWf/ttCwX7aQ613RDmwqFvkkBr5JiX9C0tJ9rx
XBYClKOzC2Rk5654+cCtz9ywN7y9+EVhs/NmX79cWuZgbESBT9elEQ7fvxblDT2eulv1OpPyaeT3
iOKhMbzg09fkwJdgEk6Mh04QjyiwHAVmpUFXxqj0ZOw50kzavh0UoKvhbyOHHKaR7W1Zx59hij/M
QSXRDuV6OU0+Xolz2w6uumibyKyEiyJMia8BSwTmenH7rQPpDLh+Oy8xzu1BYwz3SX8DKbVvTT0E
DzC22OnDBOg2e0ryRAYRWIgnBjzin1lOSziHKElDqQ9l6J9MAZAoceHHpbKvbxowgCyKeB/WEUgG
Umr7TzMLhhYKG6RZRXapLSus/fFT3Ewv6ckpdMyBbFEAIBV71Bj+PhjukuEOm9S3sUgCrL5gWlIB
qkVKExswhec5zFcFa3hjyZRDeBtnqj+TYps0Faj7Baq5coyRUzN3nxQeYOhrlENZbgpKjtgqYPnz
8ekxa33yx0Gzgrs/iUZfLizHKNKyCdZ9yw9APK3cElryjYqOxU14rD6Ovv5LgwcU48CAGLHiKvaV
oaksBxCHikvn9ino8v17wTtFifi37rAiotKj7ZQTmn5lCOm3sqJzwSYwWo8V1tuR0YUWz3+efahg
teEv9kna7juoyJ4YPTggMCWDdViPvd2xjWaqG7l5sIWNo6CEviUvBR6g/VffoabqBjAWiEdNUiHa
y1aH76dTo6rOQhrhUsol+lgH2IprBZKL3zd2toUMi1+8+qiTDeY6sZtAkCGJztphwIBnxu+CzPtq
hk1WkVRfFOVgfK+82bxiH/HLVw5mzT9ZFcXjqVZSeYJxEayJaCCYPPiVKjYlzHg551bj+8sWBJV3
VY7MspsP9GlplDP8bT576UWb9wA55qhlSq5xe08c3zyDN/ynijOr2BqIgroSxb3XVke9J6WDXTlA
tnI+IjYXzeazHaruQxKRpN781VN3NzwO57I7BdmYeK12jhXseHr8/guFPimcz7J42/EdyhbT/dyf
UhnToDU/MLqjIbZgiBA7qIEg9Or4ekJfs6lycq58h52VPIRd/iYw65jFYnKanhC8HCK7QdSNy9jh
oLI3xcePJPum+PMUzsBGXT9HD2bQi8YRmSPCq7+o728Wg8BhxIz0oxrporhJLjZLNw/G28qLPlGL
5Ed8Rp6q7j7YUeH9gzbtedl7oFduHQCE8/D5v1Pb4uFO3kRpw+qUKuFh9OEqzSWSjhOmWHW0htYa
1XfyJJse3DAmKfv2bp4BRYuAuqf0UI2PDFIm64GR68Y6c+15+LnwnwOmP939Xn6KzDV20NEYaNv3
25KU4NGKi7zR9AZMBP7GiGm4Sqs8omqjEQhQ01iJvu/xBdFrW1ei8fTC29pLTl1ZprqdW1XXIH5A
hHuIcJYhzq9k5plmbPVy1AhZe6ulOkglSfTIPXmDPiXzwzCgV5SHb67C3NSGFjFahBS58IMydCI8
HaZRnR91e+ZkKExWtm0dGvm0IKUgEH9NuqfWWHZcn5i+7GDY69ABsuDC0H/S9P6fUx/Uqorazv2K
hbS5f9B7rhQi7fKUg2zkBEiAAdTbiNSSFqVBNjY3CvhBzPr1TffOhXIRSj2puOV5ZvnVFZ3i4T/5
eZu55M5N6kulNuOoIdp+56H2ES1QTiR9iPfysuUlFL1AN+Mdy7+M2LGsfT6NJ8zt/nAXZtC96pif
fg79K1ZSIKMFEADiPCnkMW+5tvXZusVrjxz+gJZucFBbouUtLJWsognv0bzVfMly9iWwTP/jX05e
6/Tju0anZVJHeg/ywrz20ouf1K3HXzSl8trYsjlff7nXd5Ejj0Y9gQaCwfFi8JmeJ0r+pN0fBxZ4
Hy4VCX3n0nyhoiV1qTAZ9ss5gIvHon3BYHhg3ijnUmspvVMt4pAz1ZxuavPwHcXIRZB5924fysG5
aryWUq1PXxMSBb0dVVJnL3OKU7m1edpokZIDx0+mqN8OI/Xo70w3XcMPR4FQAnFL0AMxRAHdnNQp
VibENgaTZQJ2ReLiO8gO0f6Wo2ZZC2Bkzi/rbrMilUlVU6y9CSyyiQuXwhS9HeOwoR/3Y8IUyCSg
YK1r15vTkpCgrCV+iVPsMjTCUYL3ASVIuXjPBMfd1bXK5FZ2i6+JIB74yD/wpdW6QwkL4Z2wuiWL
FUQsq/Xu4n1EmHXdx+2u+CmF46CpxTY7NxaY69ACMi/5+JEshZL0VBhgNdkKfNGcJm4JkqDGRfWy
cizH586psfP5f8d8aGEDMBQKf1k7nWjgHuVrnhH36dkjuuLttDKsG6p2bNW6tb/StMw39XZYsc49
apt54D27QBY7AXCedhUI3rjxS+JVUbxNw45PWvwQvEjjhX7KTlBfqjzmOh+Fs1pe4QhyM8yWCVov
ypj3RWMQaRJf8wt32WmQr9hC71ht3hUynaEuVTJveCwBDUX7G7KU2P/Splf6y4iArETqnd16GlHS
eskTL0f+iON8T7wAGnjB+Obpr6JCxPyF58Sje3LyL2DqMcD2KCCYGbg5TPCsM8kyZAVcte4JrQoz
lCmv4lpinE+JPMmgTvnKyeB4vvOSPR0zhCEslNfIaVq0aeCIbdzwFItgfJKqQws1R5ug9OkjHBQq
upuOYClIqZ+pASUT0B46hEz0WUZr48vpnp7152Ee0tFE/GmEo34aentTVsJeYEpf8Ck8/rIDTUwY
kkVJ6tvaWXlRYslwqOao1kbnGEBxmpMxRX2LDzOm/LrwGI3wLwxAE5y0HRP1MNJwEr2gcRlPSWeE
LrTgq9aFDTK3S4m0ORkPG80RP4E/4w66+MYTQ+kUDG5OoRzARbrmgrflG2c0dfcoQHKN2hkz2SKm
VyUqA1ud7xAkZCZ0Vf/ZxABbgvrYtjT5mI0txyNYoDdINMU2fnPR2llulOtRTniNiF44pABVFgza
poNmgDqxrMYzAZHKZHezrcmg6SrOfr682qZqur8gxUdZtqPGiRb8d5G9CE+aG/JEO4xDidTw7JBL
aYJJsX/zBAKbKT8PsTsSR4gVXF1BQd40FXcCjEWXYokBQZgL6rkIV30mSEySha3QtcoaoPBKGUnI
WPDJ86FX/DPKy4JQUscR2RASMtb+QrJIagNQE980efTM4SNonCcIplDq6XGmyqrKtz5X+WopU0Bz
dYVlMAQVXX7Uc8vNrVuYCpopyi1kREeVMfpGc+lt5SYnc+1eyl5JTUHa719HklgUzddXD8N30DzJ
g7BHZd8fNKlvsrnzHMTZjDatuTnc1r/wbdfdvpOUpH6Ajwc5gyytabuNXIPvC8ENHmCTYcmZ+T/n
u4Gkx7cntAOFfB4UsWPnDjqsQxKIJD8a1eQzeVW7qyIrlThYSj84GhkiEUFerlJOwpKx86oXn1ax
FK9ATHoWcPyTLNcJoEj3eAcumXWV891Y3bG3GYwwKbWt3LtXe9vIH3wHxyxz3ecp8/gX0J1w3NQY
Nhdu3bi/pGpppuP32Z73rKDm19m4ZU52f61YpmDYN9JCseQrt/5w/AdoBGw5sa+hiqLucwYy2nO1
hyTSwJlAQ801j8Gc5E0TUZHREHS9zyl1uYdgoN8Mtvk7CzKaDcNs+Iv+5Ev4EaTager7bH0R0Cbq
LeIaA3Ad6gqNsy3KpNIs+NqiFRPXXlwAeERNwHeDZjFUhYKzE3YH1qwffqbc+kyp4i0/6YBs1FdO
6szIAFJTUmy8ZlOe+9vZ5em7eNucRi2WwT37PhHBomAUgmp9gE8kZAaC4muxw/SJY3Gra/wFaAit
e6ORJoG9fHVxEQabHlyK1iwTLkxfAmBqapYRknpy1TyiqHKHjUcxHZ4kaxXcDsvw+X9CXeLkR1zU
VRPyakMv1cK9gHtenlgEnpuJTj5p0gRwqNqirClAiHefWjy8tEqi0BzwYR5kxB4bFuRU50xe4rLp
L6pqSO6goxZrJAR5aXFoZycpruo7s2TjI4WJh8pJhvs/ApQmQj8Ybq6b8cICI6v9hoLy6nghmUob
wiQeuKyf5hh/9oNwsG7ndaM57RzQBGYMpwuntrwHx5Z56vVcsHwVuQmBAhUt22rC0p41RuMpc8KL
ZtgekiXK6BjSQ4Ts823GEh9WvwL62z8a4/1uN/BtQB0EXB+9qTNjh95LsM4jZ0min1tVLcPJPM/I
tlu0Zf9srUiisj9XBzyZ/aAF0x8d9KRTq7CbkTQnUBAr+W2Q/DEu3q0btxroLyGICD7Fj+7Q7Pp7
+x7F06vEyfyVvAzriOWSNOVctKQO7BD+1RdYl992mVyPVJgSlSg+hTtcTTPv+j2O5JoENNjJXq1O
c8a/KiWcgsuiAHZva/iVBRAbMVzOBDw89km1yDaSpLb+ke20xQv01Bd3SClBBeNDsqIumLkD5inV
/VOnCbCSZCT8zvg0aeDFaObnOYEBRtT5WabxDaDvp/AXvY9bnZCibpGBQJ9/V04UfAB6lV6mAUb/
VdsLZHRAS/aE/PnfMRTPKGGTUBefc9TJSESBwiWPUjWXR8wDu45Wx7DRU5PW/2MrFh0Rd5TpNzvP
k/0x13zC+jqGJT5xMzDeRJmH/3es9JO1E5DWGKx5dIN44RzODVbfkqS/oYpduf+0WskCp3jStu5l
EqjDhDJFCF2CHjQZe2W6ti5da6ut7Fp8vYrakgZfMcTMzZdaVhKr09uiHeJB7F/c2mniEhE9lEb9
R5ZpV/n5hzDVnpmAwe4Jsredx92/DVGo5OliFF+qc/Nl5sTFSfTkxfJk5RCkgRe+pmgK1SFySBsI
hPCAvkwUSdy4XHJDoetlCgg+KVhzyedaV+06zv0QA0WVVH1oAhR2NIsLMe1cGai0aDb23CjZWjzH
rVX/zP0LZSUNSXn+/yRMskGFtXVZAIUsI2LRzhTUVm0CRVoWRhgEvPEODT5rNclMujTCRQwzmw/0
dyb8b3g63a94LeC2gMhGlrEeFJkon07r7xGgckyIXT8gNexQDiomcWEaPalcKOxJUOOvt6UGeU4d
zKAh81nkf65tuu0tYMydQ7Ld3B5JOblN1u2YAbylncyEVGU2XSEMDRGQBx7sflSeNH+HiOeledfO
BL5nP2wVJSjlXMUIE5VLyyLJRNttftiwzzira1OmilJUFwUKfKyqT5+fe8Dx2Io7WxhvJ8GEAnyF
ZRsHURD1sAJFCfl3NB5phbu23xkEONsWI8pZSI5nMzpkhgFrG5CYthOqcHPFGWRkm3g/sGlOv37t
uY9ZdubaMZMxerg01BxzDaQpjeiYbJSvK3oWyD/c+ZnLjudiLduB+iecbMhNQn9F6iwQik9baPAa
eKln2A4TVOp2C/RVIWKsauSqsker97Z675thNXIx3849jWA+fvWwb83Sg+5ARCYXaRf3ih5lliov
Cdt/GzvtHlDr4UnEg6xE2cNYFK8TJ6tEgL+1RteddjAGUMhffeO5VBXw+18C+qJMhr4YEIvNlyhq
kPmIgQuwKyBKviGRfhCHDyGemM88gh9yrcQcorjWVnER7/PPowHY44QOk8NzgaGIw+G25rq2QPau
7wnY4dtLBBgagx16Z2Xbu/j6YipsgRCUd8zLfEk9fDXVZsYawCEZSaJQkVCtLNV/JvWXSKY92GD7
G4JpbywUIzMKfxudDsnbdW39vv1GoxbmYn+XtsdQWlB5OaZpFFWBc0eNwK7MQvFIYlENfS0hSWvv
ZtgpVDhRhFNiLYgORGZQOvdy1SCoutv36Esa1f6FvpvPu6Q4x5i5hBnFY7hyeEgTgJQ389s5+pQF
95COWwunYegLqisKMotZ4D8bzWfwfh10rtE8dmshgC52MdYB16K+qYS280tY/gr+1gceHabruszZ
ed3Xxzfw4PhWF1y/rh+o5ywnSPF1kVfQaWE1+QMhwkDmmaEtOZKFoG82NbNmIZ1W8p6pKcC0tpbe
4hW8ysi7UkVJCVb6K96cezT1uIrj8WHrpS5Po20t9nOxWGWvQEeHMslTX62T0p0QHCYRlLHL+/Ec
U4ShBTQJzjCa0pYd4fU8OPxDZvRHD1hwa1Pm4RHLh9MQd8R2dXT8XH/rzZk8lm18jH+9H2CWdghR
fPIg+ELhIdJMf6wdFgliGEaiofZNxZ9rT88OgBNmqprV55KwoEfNfTsWrmiXf1JONMmX+oY4A8HY
y2MGBCpMz7TNHRfH2nWQxw/yCZr4C1USnXcge1SPQcosg1O3r40jiXlCoJBbBGdM2OU2fu8lM3id
BIzKcOygHqvcH0Ez2PdLyXBgUnrTTjy3i4UcFtydVhPXDQOgcJ/P4UQlHUAmxpCttdoS96q4bH8A
VIe07fJ9zyN8KnI/35Pnl3OsdqdpLBBYhV9AK2DhIn8jKvF0SpQDOBOFj7wCYzidhIfPjVwYC/hy
tMXkIslgmzmChF3jdcelTjkHjdoMxQG5FVA1eHVg9d2PzjDr2SSGw4FJ1FUqS3FNGfsT+0mw2C0o
7mETkVC/LkHACxlSMcj7J7V66P2kgn/ACZ/QxEXkuNfrJQUDfXf0Gi/b3Ki3VTV5VF4GbBL24huK
8taNBejDCEyajdKxOQ0mXTE5DADxIH8qF+Zc4ZILGFcgQ2ght6KFRboiRYcbYUP2BqGXZe3QRaJy
Vwkg1pU8F8QbPVzpcA1cWlSV78sMXVpyUvMdHqjDcVfTkyZrb1H5sVJzTHqm9Mxw+zHOkvvsxaDv
4624pMY1Adc2c2F32cJ9deDtfB9HySeVTKhx5k/Hg6+41jHbT+HQqTO1XA3b596UKrobfC4LHZVa
a9W2vrVu/J5gNi+G5LCnHlwsx1Lw4ETJ26pCO11ZQYSgbk3eT5LXBub9yK73URA+ZbPv7plKXkdJ
5bvi90g7B6MgEimCSG2hb+Rs+aFedoQLoWLxV38or7foO6ClwtN4XHZNxpvD2d25OaGW8SYz9aE/
SYhZi+5+94dJRXGOp9T1KkKpA1nK6RLH5VIMUPAfJ9BGjw0fJElZ8UJmg55+jTVBYSCmjifvUafz
cJ9jRV9VtmPpxnH5v7IXZkdwxCYpmWBsJjEJihlRaheHcbNScHWoHniQSWdrmnZg7dO75hKaokyT
oKQJaw/zRdWwcnXe1hAWMzc3wIHdiphOwQ3cu5/d5jYxBuyj1MMFOYo1c29eRhVFXNlfrU00Bq+S
ba7PB10DT9YgF/sFGS7KlCgNKDBWJlXXKmA+S5zF2vKsSknEGH8ZEQfX05i65tEVeeeAcGUiGP5K
76beSLaEGb7yg3DALgU0uVTSw6VTNLPphK7ZiByjt5BdXFgyu/ZEVkEnPm8fmap0QCPAolGNeMKJ
0zAI9h1YnsWqot1+k3slOTThsLlWozxniY3pZmegMpt3bXPhXsdJh8jzFBq5uiuhmD9VeVpCSkds
iNsBBTTmnMX8Z1ioHf73eYII16rpftNnPg4RjrEVNaU2J3HiowHiU+rT33mKFC+4x3Trkp3igvkJ
m9O8f9Y1mPBKjmLMoLYsbNdZnhFbznJGvpeWLZXARTZR49ibRxz8VT5qxgMaHMSvS3e9grnmOWBz
HqC7adVOu4DwJuDEUp2HY2uDpkurT+c+5SW8zRSpyhzbtGo29fBOvd5YA9nINWrpPwPrtdVMU1jm
JMI5p4s2ZuEFB8RKLGTLl0KZJgjOJc5vN3fmKjIk8aqHUDL8Es5CcgI0c72n5cp4RuQVHx8rrvso
Hqn30WOY1jvbrNAQvgeCyEEJ7Su18BPtiSgtuyjw3L9kQYweT/qhEmv/UsHru8obXOG+4qGo5Ra/
o8OF6vqbviqtVsEv4HsCNQJTDGI1xSp6aFYMKIpM4Q/ss5903MMSZqjPfd6BX+5UDDRFjliHB4Mi
vZwgIMkZiV4pHwprQUYX8YQ63rFV4YjC6hvXt0l48KLD//zSEyUHZsQsjiaRZ1ApBBvJ4vUPvnve
IukGOURlGgPbzwWlZAueVN9J35gyL/ML8AFsbM3+U1juN0QBhAqZIWgoIRrpzDyNRIi7aiqmvdpt
4KmldPfouH3HypgqZi3CmM15QXY40HL5HZRXIna8sA0ynGGxOMZZInQZxeEbTaH4UB4YLkFgafPw
mSa4hbRBf4f+o8C0afNLbRbMpwlTf17P3Ju+sPDli1asNz/Z43+SH8/oQEHsdGmrbZ54X7LVmsh0
p7g6SEzhM+jPPPfhuqOgB72spMx06+TNLjFMxL0DTKmBiXXCBn34mlBq35ut2/q94um3et+2dQzN
cJs1qCX2JOIvNQiODvQ3Eed4qSPdNhAZEPATWz6LQF7ItB5e+hd4IBlE3NCFkdtS9PSYqJDwhyE2
eWsf05Y4dCtDxODfsijRp+IU2lBfPKbRgbjM1bvZa48RRm/nDIjKUo7TS5Cs8ni4BZ8WSYaRDBs5
jQc1Dknha0Ho/wXwNjojW2I/PaGbQ5DLoiIIp3QmPOCjKVu4MBrWNVRsBFdDKhFG1purRPNs4N4F
YaDb+Y0LUwCSuQ8u5DwvpRNOUb6cRml70DR05dh93f5HzBHqSyYX4RZ+L/8nMXJyt8PyS9NL0VrG
o9E9zHc38YSbOICNMMnAaMNE4Gz4AMKeHGM0V6uxPw4Hb91RBVtRjSn1MU52w9M34gktiHyh6lTP
uOzpEHAbAFt/utw6vBS4jneOeY+3OoRxPujL4SfAFSba+LcElXIYLshxeNQkRaILzVvdNh43JCGb
27DQdYKo+0muphBDrhE5A3QQLlQjfkVFrob5ENSZQTEKIfuVy1yg3wmBaI68msVsoj8fklMei5SV
EGIBWUWk6K5OB6QRffga/jdqINp9RBeJk6d25yMIv/B+o/rKwMyRQftv7wgCHtr53ZYYLOsFDYrj
jKNnfMMwgu+l5TlvYq/09PRMT8dwTeAa5MHYlMZ8dB2Duf0s3RtWEpRip7Dt5EwkRJyeyJycfDtr
V840wSXQISlXTRJNaQlxE3mjdPzSCkRmmItP7fJ24si1elcQKvXFU1BsVw3jI14mpczA+oNg0FqR
hf3Oq7oNsvGkfNcIvdFyJAvDsUxIWTniB5ESChXn127Vsn3uXkr9Q6SHI08UG/KKnUED5vFIxcEO
tVy8R7xMokcRSaU+ereySVkLeA+X999DKFjoZJRUkEduyi7fsBX67FYbzOa3oS2UBxk2b+QHHEm0
jaWQx2eddkruo29qFtI0f2VftTmnamImEPgBi2o/8ZX/mIVmvcCahrV9Z+JTYVq9hAuVLp3QjTQs
yjGYdnt06IPLU0mWfPWTX9kg1tKsULRUq5hqbh0kLEKq6KKn873fgQ2/AjLTjiTmn1JKsFgTaATF
ZfZ/Ha1QZM+sK8Vk7ZqA7sOyNMLbcgebuU1/Ls48/EaBRpNe8LzgWYYcug40tzA2eFmJdMMBH2/f
KUOCbfUgy+xCmTLp9qE7tnvtad7R3zXCuJ3NcYCL/YY89ZXRJixjOap5L/9jl+K4X8u6PQtr5l45
VI02tPWtd2m8yKn22JmQPoibQOC//AfB14nFxflgyXKE+d61IVRJb7QdHSYYr4X03QEWx+nfmQXJ
Y59aay/qw3gJHUlaVPLH+D+S7TaHMlhfUsQ0nJe0nu16V7cP0Ooz8+VPvjEsU9HnxKMavx9zga/Z
GOwQO+K98I3YukQHGia88Q79mfHU8bCApX+gw0yrhw26pg0/gB4GuHwQqBs1vjHvulpJYG4frhsu
TowISh7nqABgHhlPAl7ifmIQHoj1Vn7Zt8Ft8+Fy9IxU4LIpFFf8C2YEDGyyGBqd2QYPecjU8EKK
eH+B04TYUUGcJBQeHjO4ks5L2rKFS+JtdtYgfL/yuskP2rHCBxLo5BaKTs3jFuYsN8Mt0mVd3OFt
0zX0u0wnROV9Fx0opoP+lBo4R+FFIkh3EWNSW/RBxmDeKYTuC1+5Hzo+be60ki0aJI3cngfaM4yI
Rbe37zWnAp8WRKt/Vq7nfj5aNRl4451EbhGwULx0gtjmXB+lGJv5ICq4YgBR66jK1PsTIlaKN2G6
bZ/plQx0hm1HdLQvSZ5DZQj5CMgsDCP7mXKIU6UTFLmGwzEEoOkKj3omij1fNDpdAjCJuUAhQ8lt
c4fGyIjZruKny4lbEINOPBtZV4u1T0gjR9KsQDrMD2BWwO9g9bEypbmFKk0BOX9MwV+UKCMn65uB
tIkJZo8ENYkXTW9h2D7WNn4k+UMqF8zcseWLHf4xem2RgEIr/l9pMomc8AJK04fupbzTVB3iNshs
EHy4IqlAQtDK1o82oe27oglJtenuS8QBCJx+SGUcSHeCGWKqMyU7ZbWuZ1Z7Z7X9ro06y2kA8sTW
mQ72uTVTp7qjLyWPHjmhHMy7Ym/ZbvR6BIFdMzN2QH5Piq3BPGi2PXppSayoMwX5WKzED+IMhAt1
yJwwbbwIDT1O8NDFjZ08t8qV/8ALdp/v10+tE3wXlPXPtUE2Z4Nh8Z3HqscKdHOVzPAem5L2xpHG
BF/SYMT49JkiHsLMOG97aKmuMVURl8UYkbxN7vKq6/3aWZG1cQJBf0J8+7DlD6kG/1mySqPRsZYx
7SGUTP+D3FzFJFW1iYVWT77yIltlD27AkBqxhgWi1zdEXpGpc8OHkO4onvyLRoYzaCKZ4RWztv3p
2Jkn92itzGQcZsz5WAIAhS1yNaJc0pnQjF3ByY56nWtA8KWPLWrlkSvikJHDaqNlYoWouEBekudz
LUmMhC/zHJTObtxL3z0y/QZYX5ADJtg6AoxWZs43MruKIUfH79eQduHJUm1xzV2AIH8lmsXN48Ze
MCq/q31pdG6VD8W657KiCxBy5y1MLhM5nD5qezkBTM6iSDHPSyJINxqDET5oiBtDQ7bxCNzhl0dH
1X2tGLcCGqL8hHZjNXNWLo+xFL6uNF3JnFjp0XUH4KDkC5hlOz3mWJ0B1mR104wOwL6I0rM+//Bw
E9sZo1E6UnIpgKyCjm5Sr8WrbGFjuVI+3/jdAYkar+X0eLDs3DPc0kBK0h3i+XImMENZW/4ev0hz
NDKc/3dMGGqfEenah48aTLhBJtC9nTgE3J/G7PiIp5rIsD1QSTQyPRqD0Y4GRsDW5TJh1rgrqGDR
weeUhwpl7ncRChCSVZwNC/mUTUb2+yoiNRbK0ihlLdy+/wc/ZvJx5J30nkyCdz45T0Q6YBrpXnOM
wDl0jjR+PKBzPN1noNfcl0Kt/Gm17EOqbL4L2kITayqK+4Cxw2ZRgcwWpo7GMmNPLi4hqxkjd/Mq
4O5ee8D9MPvuXoPfcuepcGekEwsOFRSHzEWXANrAMvTt4lDilYv+UjiAmePp8BvkOIxVzRgcKZqc
gjpdV0PoMUvPxm4aHqs0jgggXvEVdrM5+cf6c5s+WXdm+Xxrlo7SoKAZb01cl9KiFXGQdu64nQ78
Q+IGs3oKv2JIf1ypmMxNXI/yq+6D8EsGtewmRQH8XELByTelIFGrzhHE3HRd5/gS/DS+ReukQlYo
krpkFi72Q7CUS7vPqH/8RuZCQo0JI2NXMt+ELo274Ra2dLMMaGVeHVxUIxarn4a+7pZrAx8qZMuk
DJmKv9B2ATU6v6jDAP6MQWzQIGmRwP+AInNW2fW1fydRxQ3Fx0F0pfciL1DdkFhekaHHHp3m0ESV
8qASNSDzx0DEG0WLhoSoiOn8UaUJbL26g+s2ukU+yxOJ+TFJYvk9L9ALRu+FyW6k8edoujrwxbmD
Z49dngABFMRE7UUD3E7w5d9181j0EEoGC+kt0DP0qd7cd5J2xe3WJ+nqHVqQZRKWc6yR9ATdRIpH
myvA5b+bXcw72qT9K8hmbmA1+FOUajKDr2Pl+jttzfV0ytaQjkN1sw632LxZakl8L73kGpk3154u
olvyA1ImPjM5suJaI6er/fAV1QUgo6LdhPUNkpnJbj+owbrq160g9ZoCS7+wx1ShsNMVfX9ztXJJ
ep7mH3xnXSDnwM8hpiPFaa/f8gBeCxj7EJhxawAdIxChRpT4qBvbChMRJbj9c7zuDB8rX35eLy07
SwqPOX6rh5a6OoS2pg6twxD26xgF+fDFUXQLDwgejonIlExvxbUkPFun6wh67iI6t6tKt/hq3iXc
eZWLMz+B+nzCh9BFcpqG7rw071KthCLZ1+oZaMcTC/9Nw5HQIT9XPYG/0GYU+2R8uxyYqe6Q+6zI
Ev9yp1IfIie6wjHXMzXYcql/jo9Qsvb8sTd77/1110blCC1F/IkS9EIRCj/Ykmn6IMkVjC7o5rz+
z9k47Cw7r7GMSKp0LAOplIpwK8sF+l0mbGQFpQ4Ks3nEGW2Acdad1I0H3bSAT7LWYKGHsNWCyQkF
GPBLGRCbMagUHkG7HKGc2I4StMvyQm1zZzahZgg9klvyE9SGHtQAHZPltfRE+IW48Lnom3uvOPyd
/hwidLVUukO6DIDyTPZ7CCDbdU1pvHnnl7J34lQi26RWKRRIaQftmegd9iCaVQsjp1D37BId6As2
AyCDotgg+DlL6PBUH/S7jmm7ls7SWyv+ERQuEO8uVJ/3FsffhP9FTI/E3Du04z26Y9SOVwhHQ3U6
51WbjjVqa3LGoTJb1aLmAOkltKSaMhLTvgdmim4v9hlhPfZ2qyZqfgce1IACTcgbAdEE5URh01ig
XFCcpK0ZREzYXWnByuAqier7UIsYzJZHgKlLT4Bf8yCyFMODL7zv5doyLgrQHsr73f8vCai+Hync
RebYp953tUTO8Ml6srLzLpWgPvMRGwRISXLBRR0WFuZPRw93HPPw8j8QUmjl4fVJKNFeJbTygDMi
5ZoHvpQfAziV0GnvRH9/OLF+2/f8Yi5wOcT2w4Q03gLTB6Z1plG5uMKNw0wzmRc8FkqNhNlVhXn3
7/+DatbqmGem2Qvp83mkHwHIl6ud+VgFJA3VDsYq9aA9NG1TzGtI19dusZZ94NrVAAByM6kOLoAR
iGbxgwtz6/gcQM0ncClWkfikEcC/hkMy5suvFRDL+SJtdUOQ/KFmvjSuLNC3l14Lzg/TOVK/D6We
5CUFsAr1WZFl/vIUdeyeHTVwTBiO530nxdrbwDtU40SK4VABRyT0a/KedUDSpe0+Of4zmplLDfeX
2ztoA8ozhbvtTI4OSI813m21xZplewnPwxSpqQtBMiBwLvBmp6sHBYJiJ5vMm64wbfW43vSlas/J
61OGsu2EIXGQR9MOjEfeLEnPfQupuc8bD/WgpTNJtPnW4pY1/YPoTmALRlZ853Y95MNvmZ+dIg3J
munMmV51OMkFEZw5IkWW0n85CIP8K99GVsOg9h/4glVM8zOvBGFQucUROCMvUnGs6NJLt2vL6C68
J6ZJLC5JRDXYO0r9a0ETk07YVIhFD35B3jLsBGd0sj58nN42gX6VGH/BdUMGLtMcHAmeullfe1/j
nH01XYkYHufvjq6HT0Xjdp54IQh+AduiuEu8VbFgJsY6GiW0+mZL7zRBE4yCdf+/INDvw7z3A39z
XckvJ6zaz3kYvU0INQr2k0xP7CuSruQI9RCT6QnJX+hzONrMdjH6dMXJK3SmHjM62Yf5DWjjT41T
HDS78JBPQaBiOUThlNnDvU8U0HIBWFXoSu6FKYXA2hJe2LKjBYtCFAoS5B0ZmxtV63N8xcr1qMk6
7PwTVjwPhmTO9I/4MH9Hg3rwBrDgqn4b0JSCKQ6zFuVj3qzz1XgSENPHmqrtP4dXZX6Rexj3AOzx
g4ajFZUn7v+zNw6maX9LX8ow3pYuiEO9mjW6Ft7J9wD/ApZWR/57CL36pOhGeHe6TqCXjNc8M5xm
PhIzqNMnhXdwDhtYZH5BKPRTjpEcGqBQsJ7uxpv2v8v23gn/kFQ0C0S5V9NQZExBZUfpgi+XtLpe
noqqkBa9yDHvfDmfN2EDeI4eUzf8lL64HfEfF/pMTgrY7nY4KsWegFi5x/a8IEN/npAafh+jDIdP
Sh78TXgki1YEUQfOREuK3YLYyYBRWlq/GeOMyJCgj1VvX3u6aycXAICNQrhL3x0DyudMaLLRXQVA
aIevjjFUrMaR0P7WfkWqjcdVOoCIniyS7HnxaWVvlzIsAMRvKzI8qQgrD4Br5wv3KLsOaBtyzkXo
jZS5x4nahJmipy/piS52A7nWcQj+ylS3jNz5sQzKM26pNkoAwnBfuJ07/OwThWsZa1G2TT3O+CM2
qbHnTi52US7gb1GJ6C+GkfWu3B8hVP11DKVd0Q1NYqGGlw391y081v/huCCMvbjqzyExozfRPFpw
GpKAn7BrvkofS/hBpPHXbDuw0xn3jvzFpPOXwfdacTps3drYz+wC6rMJIPxbY7rPv2fkbgIrJWqH
wYXtOdr0CqKLVqRuZI4VbCU5ZSJthnSTJP9EKa8T+1GkB01D1v4UuJau7jQSVeV2mHMAq0aOzBU2
U9COnGVc0p2GwayQFPK36euSr3heWQL9BKyY6IxxI18A+l+SRI/Jkddd6B4OQ6cTP0QNe5vDqq/d
LkGLMhf4BkO74vwBMYDOWYP3UnH/dgQctzpp09WI9Ri/NkDB+jKy0pZB17POwG9KERJolL8y21VF
XB5Ntsj0glbayyikat8tuLzL5dAhQZvKLhSxxnk3x94ocMaBRvSnW+5cu+VMp+GXt5PaL3z8TpgT
uJRffMiwcIZHgBwe9EzECzHeb0k5hJ9bpJNep9nKm6WhknWiYxBB7nmQ9XNhnY7XOcs+H4BxXPNO
K32tE5cFpZXk8ivGpfQtt2Gpow0Xi7Fop4Xapg6FCLNrmrf614nBon+gpkQft14XxVMnUhYpVQtW
AVjUWi00Dj2P5G3JVMniqoU9VbWYW2DoTHeFbRu3YlrSOOz4gGnykoHQ3xXcUjgpWQMVD8LNqzSd
HbB1Yxk/PUuT2tzKy255zLrHYxckarFivF+7pA5cls4NL0x2E2MkiCijQVXPnyVZVROSSFP0vzks
qU1yDvhjms4MP6R0t7D5jtjMVDvJW+EiESoCL1F1DwN4oQ4ejMR7rEuiMekDdmwagj6ITjBsgA4A
6RTAQBf/F1hQuw5rmwQ6tssLJ4iCY4otgJIYlghLspg3UIbkg3MyAgegiZAaitsudtDz93Us1ySc
OriTJDa7ESOGiR9kkGnGwxiRf14fMElrJt0UT+88iSS+hJgyfsmBnsrklZ9NkmEK2HU84H6lCaGi
UJjhap6vvPeatTpU8le2etifD1Tn0H3a+QOi2gxLvJ9ats6M9t/VIjose+1z2V+E0fewLI+txzJI
sBTuen8ZTjmN8ce2V/aZzqE0rbP6sI7lNfoXsbF8EnX5M2f3cdFhz9crcosp1FEw9L0hDH4Q6jyy
ZlnC7JJr/hLAU+QJSAvYeUHf5AqOk1+CWmtuDSspvwzlc4e6c5ZU7ycrHedFykEQf+bxjaKVGnZu
ojKI8XduEfj73T/MZozP1ccTYOnn+VqjH46zQI3hvY/XFLXrlkbljlKCjaTfL+1KCXHDySbVRQ7Z
Gv/4pVs1EixQXPF2Lu6DPOz6+WAodHiEgk9pI57z06dYJnwxWXFLB8rgT+OleNf7fDp4OIgRSLVB
yYH6VC5oEWpvdB9+ij8wMDe8us9ufIl3H9kzDbIhewLsP7GpREDo+Kmd1ujWPGG6TGLT0mlYQUFU
Zbwy/7mQge4tmmNYW2hAlA8fOfa6U6rT2H1Xvv83vEvKLpEtF9Pxoz06okPXpRlVVPXX6//MrLzW
S3KTlI+FCMjUl7rJ28ETqxOBtM856FZq+GAJ+CS1Yl+MZLP3gm5ZgucfoL86/OGq2y/YqeOcRXLI
UxnZ7VLDwUsvo9HXw4PqyuOK2Tm6dQAyFZm1kg6bk1tsNCABskUt74NMUlIpWf4nUGKi8E5tUY1D
6i3VSE8KLPmfH5v1NOlm4Mi6acXA2wCwxL/jSW0Cv4MnyBHoifMl9GP7O7Tj7+whtHvbfG+H/7a+
T1CUzedPlLYY3jJVFSg/avJAvCp+WG/3QAe07jwvGJgSFkCouAXhqM+/14HmBsM/VNa4MOWs2nAD
QpwAJcSDWuP86vfFTxCc/N8W22xTp1b8WEovwbELrOEJg0D4u5gnFxH8Cw7YMHfiqVsB8r7BYLiH
vryfjsEgjlv2j/WXCu15E2edcv2EirY7R3HK7Q4shxWkqe7qz/fNXoBY+p+dH9RhbgClD4lBZNZc
tkyalBi0G9IOtA5z03YPzG3s0KZQgSMHZSA9toGQYBVL+bwAY+B155TbVM7zOXnIcE91k5vi++Au
Ar/FCqEDArDi98i5YhMThNmWB+fchRrtDe17tNBcBTH64qcAs4f8jrreV32MvbUGxtFB3Y51bYuA
qU0H0iURqhnfV2/gbnfZgHSBeEtAihQfSbZWvBaHGkZY7Ai3hSve57JCT75Avlfm7UO9ATIagrhM
w31xrwO+Fg1SqbmirrP5ejNZT4avldyQexDRrXeeNH6lkPpQCmlD+NT9yvJlJaQKEnOTDpgY7EYy
uQeJAOEZtWyPKfFBjHf8zwdcq73nBgPXpav+p1MVOc6tPBFOhKjh0usvYVyo9K+4ZgRLF6OL8KOy
ewWOn8MPyTW+WAb7jtTYehNBkxIw20jJ+iJJL9kMZjsTfPuQ1VTx61tnfw1slTDUnsfCVps/0nO4
Mv5LC8yA03cnlschNiK1MUMYe9F6hFQ8rhru99dGytzpUr2OcnPOXZ461DYRBByR/Vy0Cv19Wx06
F5J0k/HQph+unDP8ObBXzxOLQ4mFZByPg8rqgCXl0XYIj879n9spZG7sHPUdSF6V7FsvuCkcj3mm
BAaYkb4PHEMjo77bjKDZP5h7t2P9WJODNmw4LUgBrTMQg9TnAhSs1HDdgqAe21LVfMVuXWTe0Hhz
spostqvWNpCZUBo4qiA33d5AOi41gKTdGTICw7wA1845W/4CWIxkwGw64tOWgE43Cbe2V4gN9fYo
Cdcq6T2tZcnFp+J2qIPbqC4cqSkNu+EvmjwADkDbZ5dNQv4BufECWbDtHwNecfTmrFaV6smwUPil
1fuf2LZDDc8Xr9o7BTJFG/ZUmGFTgj4wBnWJxlQkVfwq9tHTh4cWHkaFBfDT05nrPQRDu0zcex7t
dvY22ZaQnwSDS8FQlrVq0T3x6Rr4KkxOhHxWspR0SXw5It5gOEQRhmaDjXfesXbtWfBeBbk+kmEb
0w/x6tA3gSe8494j9MfU+DaNEOApWnraFdf0UTMsudVXpelXR4noOovHdZMbX969w3p0//JUcXQq
8jyl7qK62EysmG2LAhxBgBJnWq6l2rXE7/QwOuUNnmJXqIMYHXWPUk6FyUaoRhonvkaET2u7m06B
wKQInYLbDV8uS+kNwEH66v6OePTaUvHIu071cvSLhhZVKeKLOBPUXj6FZaBY8955kC9MCz5CcusL
55dzzBSnxfSHBJXMYWmm1xi0NIVyvT5JZOkhu3VhNmY17fryDLluOgur4SAX6qW6TqP7Lj0LNRj0
OwZmovNd3tyGjbpOqaDezwYbTgXuKrTQzYld5KLV2UtkRwnVOugit+AEiYY3uJqu6Do0TQn2Btm0
Rdya/K7JRSURX3OxUrKrneFM+CctVOXZ/uKFUpxp2iBiKGyzvefi55vzDEiYoDUtncFWN/gI/xvd
nb1AVmt0H7/Fp5p9GtRNnBvA1oC4xdRYgN/Cj2jFYg3QJioPQMp6JtjW1y3wk7mk9BlG6cwp+XP1
jPlQG7SHp2U3jpgi/HfUqe93kblqvOdCxrnYNZ4r6kUgjVw2tBN1No8rPAvvNKU6a/y33qhF1lzc
bU9RHYmpVsMdU6brdNNw1yyb+84foLQ8dboJ+1fFL/XUDxufypQLN1i6FjAIzfX3Yt+vPoRde+2Q
bIfpbkv6ZOHXsE4xtokp1MFgWMj//SCDrAf1hHkgKuIEWIMg+sCy/+mdN1dWFN0Mqt7/INU/JaeO
I/R2cW/8uDMZM9bkJ/zH8+n8RxrHhgnNK+G2FEDcbqoexUFUjtYakOLY9ZLq0Lf2wEwsrWdYNud3
NOnHPmEgbMfYdOs639ntffBYne+j+6Bm9Kk2Ig+NAGuJS+vMpsTCXyX0ViVW06238DR6YMDmjKXG
fyonf+UiJREk8zp/Ns+yIAK8uHFqBLHBYqaVNeq1O3/mhqTTQ+VWsfjuK+E54HUwCRyXfhiO95gB
kTc5CVbYo/1LwKRNCPyvgx9AhhWspxz4hY3uGdajO8QaAnT2GwS6ltN8v1Y48nqgjtB4chwmFUN/
PuBwZPkhebuSmG+Ce54hINEpe+Es+Iqkkayyw+w5A1OTfBKFoHi8iew/wmrUoi0pLhUg1UIRrIt6
z6eqVC1uRr8HGN4jIQWxTu2WxuAhHdsDXWH80NgJgV/wHw8TNdQMI5Y8f0XEeRJtXWjPAA80B2PS
K4ZW6eXrKOE8CbGDQoERTPqHkLpN/QGMKZpifG2VGesQ8xVqc7jM8KiXaN6t1Nbco/fgXfcHObFU
PavUvB5g0h05xJBYYFaYti5jhx7MAbOonv4/3f/MYCmvWVw3ZLNHQicZhKoe/nCF4YVUEZelcAig
PA0s6DTLsdqf9+hjq6IFqaHJtGPtkY8Lr7xXIstGTNLd7e1OXiIm1SXi42f/kdlrX1cSL1GWONu/
c+dclDkUnQfstyNVwj36K+ngT5Vqd5a6E1/wg/LZLO3a+FyGu1qT3nSFPw3lkc7CVcDdG0247naM
EbAUZugLkUP19tXoD6et8SprzhXRiPuz2jc8xXq2Yyg/8Dz4hgjA1aGzAIVV+p9BQBqL/phUFZqz
mysDZdPhV2ghmI0LUJos7S4nSfAC/ItErFz/7FwRXxoXeW6Tw+eVIGUCUNynOiG0xcrikG9J16EL
yxllbg5bXuf9E6djJ4eHbbKFtHLduMTvzukPZ1Crwr/Uq7Db5kRJqPsYpXo8MotAeE59WBMUah2Q
ad7E1YPY7AzwkqNcqexl0X/KdfVGwOz65KZbrxAuIZ0u8oIsTmn0kqHmRk8w2Y5cmHPTtJ0My0RI
pw1gcRl83l0hkpxCMblAATSDSj9g4uqf6l/Yq8deT61DOZi/UU8sb1c3b39FPomMYQJWxVU+ynqB
jAF7fF92HLkX8c67NiqQAuvNUJlkR85ysR/HNBEAYH6cVkDyVWxg3uvVIxWX94d9Ak93t4X7rizF
/mNihIzoFPKh+pecZKllKLOV+NW5ZtG/ewoffbMbaRWztJC6lySMm9m0h73p9WV09f/XC9wLqJCC
99tkmGTZHGjwYlJV3hfdWeVLjY5l1uWvqISsfEL8z0nMh5f/sHPe6aNVV+p+NsiRIqo2u6sAk7W1
9+0Bmfldl6xnZEXIOLI2ZYMghfLT/sTrf4V7mbYrcsudTcjb54tRumnRjdVNbhXS90nsmULYb85C
xH9CZxzSD2p5fYn3z+sN4q2xAP/9c4VBDyuDTdADzRbPwZAOnUhyQFzAsAe/aENZ0WLxH8ozBb6V
LKgnrY7TOcmR42UB/fyYdOqc6fa7U05GTw/kuHsPnIX2paakLuyRJo4OiQbo+eQV0vT7YHavhq9V
YsNt85/HYruTddfTL7KryHqSG1Kxf5FJphG+OxhuTeno+rsggQOpKxn6si28r34MhvIAkhzx7E6L
GCRUiLSdXwkPfd+jWXHLqorcbWklIIziq+OuVKxs2bLpSGRQ03WcWhfibJe5/rBYcxvcK8B6yb/q
mw/mXNom2+KNOTapI3P4CR2Zk8IiACEMfsQFOHZuAbQU1QKYUTFXLtFviCe71hb37lgTZMtFko5s
EoN0cBJ7P5oj4dZxvDhI9LtP6jX7UjdX51Nu87FB83YE2tPwq+IdZYVONmt7VcEQRODoFg0lEoe7
8aC/Hexal5WJt0M3JmZpQm8Ze12byGrX2yz91/Cz93RTvFoT0TM1MYVkjPK3hJnC1pc1SCTLFl+/
Pkz7PYrzO+1lpbf75CQYQsFObHeIIjbSAaHJc4ZowZ4+FAck1O3Nclp+XkhwfKQXCuaH+ez8tk4z
2q2O10WOep2fzyHZG7JwC9apctIYaZBhkVLaL+J6dUoVTUOza1TxBDPPkeiUfyDKeV0dP5fJLKO1
MVfsbbOvvNeXzRERlsiSp1kLlZfoT5oihcZuQncIzNVelKvNgpvUfwzMBeD2sxz9vf9krSNWrfR2
6LLyWqGxvxKzIqQcc2Eop6jzDYUQuoeMEdurjtaGrkZ+mt1sctpLIQo0mRUJPPKQM+QGfTknJL2n
5ogONwqHxuGhDsqaTnS0J3DsiaCaT8+eHKe3fnxDA3pWDGBTbYe00sL+0W/RenGRWw3/l+F7ORa2
M3XnyJy7mY58G0I05OYxspHl7lpUQXRcQxwbEBW591gB1MT1CVky6t1VigwuPUJ9FYaqXxFiYPv1
keAA7pM1oZ4vjJwz7a7MDP6jBVnpQ2KQiOYSG7pble6T4q1cJvyznM3UagS97BZRzJWJQL6LTKet
0QOpFAKh88HEOXje+gHYPZzYQf73/BNugrMN9iGH/TcB4TkBu03aqmpWP7572hpHcMYx9kCICIF2
gBhuxxiLsQgo09DkbZTI23o+HKn5YM3iMSp6gs6d7COdXEDxaayK2D4c/3KtbyEjNQFnZvc3rfAC
LDP9fiw2NbtbeQQwViN+0VZn/Ic0R/LQDKMQyjgcL8K+DrD7Ld0JXVaow35mNEhpXR6V7eScuq1V
7ZTarsur13nYJpM1T0Kn24JyJzZBev/qSnKDXPPKH+u0vxbhYmEC0Oj/nsH2dWeUZjxCATYRNSFm
8FTZ3qVy7Nyw7+I/TUPbB6fW7+25U5XlGQAiu6BV1xKLG82TwS4sO6VLLRARlyc+iiqraI8po2ev
OCUeOE9SEULdN9rV+Zmc6tX6TYtM3zaMJF44UWn55Q98YhR+qoO1Y0i10fwV1waKS5Bwf8WqvuP5
fX2NQDBRNFmFyeS3K0C/btMgl24Pb9GOkYLPfO42/em1OIpPFfbbmLqXib6EEr0++Dt/LTMJCpeX
49YzeG5/4PndRE/iXlQwN7D2/7OB+vmlBfFlUeclV14fjcuRz/jMhuoZGDfITkPbZTnonv3Q6InR
S5m+0ZvlRxFi0obEV12OqZj1z4DOm3QSD88n6zP09M5ZhHL03MzwQMNe50HCHVXyJ+XI4p6AKBnq
El+AOTFVPUKWRdTMeii/zibX6kdIxDD6iu3zCjpf3bQxAD+vMJ3lkX6y1qB0kpoS/jF1gTsgE4PC
yUCQGE8uWX8OWKRE/N9cx0wRr/2emjjwpsKTEW4hEyOiu9BX4El0BS77R5ZtPvwXjwH2oE3hr+OA
FOuZbwQp93G8VyG5YhPpdlrb2v9ZhSiXipDZmYqw6YCuINKiz/nBN6W/H1u4lobJnBGfsceq/X3N
tNd1b7RWmlIhFBuHvows7G9+y4CK/slqedb5O1xVHPEG2CORoHgmjgBs2YI8HXvgevUMM8UsO2Sj
fVS9jtbMmP2ipdgqThIOw8JX7j1Bel4aAnnuxyLkKAKgoR52zy8KhuEo1jCY920nruQr5bXxWx4/
h4p4ladaimXhRpKYgQ0IiluO+Iw4oa+rHg6ytr9KiJcMXcBEflr3lzAE6OJ0hreYq7fdtO/zeyNE
3o0kKaaddj0Ej9MN+tTZC4OnS0l6Zh1ZAh7M6UVlbsqQWAC6QwdmFdU6OWRyyzlC3EFeVaeMBA+p
PyS5yAfB4EnFV84+ImbIcApJP78n76y/j6LMzJOCutT59gtjp9RPVAbQp18iBn4weCTb6jm0O3P8
1aOnDaNdem11OdDk0fHymhWNgEvn/okcJUcexfY57xf1Xvmo3joP7ww4184P2Y9izQ5IlQyo0pYa
UEeM/rKZBcWkw250PrfriSqFUxHCS5wG5NJV4Q4TNoIW5iek/bPFUcG2tIRqWnIGuEBLv7iOEO9k
nEIZq0TIfrmkwpuJke4gEICRtFH8qGxhX63BX1iDmWSusMyEqbguHbzzGWHkTnh42g+4RqHFEHfk
+xt+ajTVyZD+GMIb+NHSIyfEkaFdMETXEfxMpH8hAwwlZ8oxGPJaIC9LEQvv/Q8/WLHnkFCtJHA7
vlvALAkfpsxWkfs9s6LUD46zADUtU8cHOQXNCZNA0JVjILbe8h5fv42qMmDSNE7ywtpLOFrkQCBG
9IzwY9bFgcqWNGWx5/HqZHTyLl4kariBuFJztYcKA1r4CLiEGi/egF3xiJdbC/Q0h3walwfvOLNK
rV1n2jqeZkuxB2uweU8ERr+v5gT3+OaZx4QDn88pHPwiUa5fsHUfLlwtDvfJDTtYiFF2Xp5ntnbF
ggspFrkRObsjAiZ7xhC4c9I9zgEKEHoZpQ9+C0hSZkYbtQvRANegEK4AXUsxvHSp9RE+JdLu047D
GCV5WLP/Mw75uw56Tw3Zpuowk4tUNnKALBLdadR9NhqeQqnA0U3YX4WsZCeRvUJXULpf/tBTp59y
igrfI+cenVAHKw4iZd1fxsErOAKEYlR7j7jrxvOiuFgVZqHFHK1dTzPReeOuNZUYgEEBDHqdjM+z
bKcbct5MB0dURjgT5jdc1hR4+zLszwIA7lvy2lXB+uxRyTrNSjYnIudArBTsaRN+8IMyLEc3l66F
GS6V7x3fUEKLf6jjTVNn2dIk1QiOkUMvzIRijrNsEcWVOLUbo3x9RA0b6TIKbogwculUnfjWaU3z
tg6LOuwZ3n+O5XoUPShowrxOEN9e03CFsE7m31pTDnq41nbS4sc4CyhLZgEYaEZlfRT4AOuHhDPo
NfGK7mzABEdzPT0elHWENbVIPRIQpxs63+No0oW0AEPIPL1g4mualDsblk10ZV9CeBDGp7VICM/I
wnuqmW2wac3P7lfyzcGk0lTdoJfwhGRY0MrlRYY6r9TZEtv468VEVxiGJwfRDseN8CoVaI3OAg7v
qSLdfKj7YtEXOoEiKl6PSVbMpbtf5pXDtu/e8EdkW3VtcRPRxAlb1Qc5zj4U3Ucm02lq4HlMDMwO
x77VBw/hukM6Cv7X+RcYAr4rU1pem1KFDJKxNWDC5kEuOCorIves/Jy92wo6w/L4yNNs/k694x9m
ufBB4yPFaDuKWD0n26WFML6RJxj/cIbD1UoWyIykPiMBRgfkGf/gKHVCj/0ladGmEPYpWImjleW+
+oxj0RBvwFCEMCV4JAH3oEfb958qlqwKohBiaBn38G8905xMEzjXgn8ct2bfRwDQPs5uBQ+kjhyB
K6CEjF2JNCdn3tHnw78I3JvcfxyN0GZxG+2pcXSxVDFBHz/4JvbvNoCh2ZL+9LlW1zfOsWjeoJ37
1DLijBZ73sLyhgEuGXz4tqBx1V3aEeuyVqJsQu56cc708+slhFP7Jg/R9K0BHV8o3cw2p/cz7drI
43ScmUc8Bg1VMIF2j71tPeRILqbMg8FUztIxmHJynZpuTIP5W5sML6lE07EaKvkWEpTIbEbVzFmY
SgMFx5UfQYZ/YDgpOQIGTl5MVd+jiP+N7UqI6N7wTkLUo1s0tYjsbWpLz5JSp7PkpdTtQ+t/YUON
j4j7BaHPF/rFnvAJwhhiju0SszbOJy8nxTlZsWLZk5/YX73DflbAt33mYpSDp4bG7tigB+hHjS+3
sbPzUUeX5hA20Q38Ptut+IWHsK9ulnDh5pmfhEIBCFD/4GFaHnMOE1K4ZxMFKpxWw2GkClETpUeu
caaYEfbK6cnQHDDa+xZxYn4nyPYGRXddptmHu6f8l7/C4owCXor0RLd6ceNh9Cax/Gajny+fCygX
WS0C9W9Fzc1pk5/cTFVJ7y6T5vo5YF+e0En43CRXfmcFDJoe7loue8YimDsJjl8VEsGJQWRYaX9p
vf/PgrJ8qIMhPcotdp4cpPHc4tBiJoEszOcL7+IDC8rSQgZcRzDgadokf3cPkykf7RQfHYwGRW01
TqlC4HgA2B7hLyVLa3Wa+Zi6eaMHi0JHs4Xlwu6k6smx7JRyttwJaGjWsqmMQL4KgU+rinOFs0I7
JPm5TIzUwW4jAXhtRdi5tNFDQrKT3J5UBQcdJI/worlhue5ZkXwwSXhvSMhc4A225a8R5RoXYg+V
rNGN8yxe/y3sfSMzlYeK4hx7F9SUsfu1F4pfr8xab4yx78w8J03kqy3td8E4s+4ysVO0ggmn/AM2
bX5pjNUcKEHfdDZszwtu39Dqa0Tztsn4+uEdb+HQsT15YeWpjf3qVmXfXPiw6PKbLVUgadld5GMM
LL1s5j8iSh5suoaoRPgymKoynHy3lEN67E9Ek70mnDQQp/NFCizAQm54OcsxQs+MzCBrWfhEZdby
CfPxewpWUnybsqJosnfA76BAMMWBk/dS2K00zzo6I3P7whrKPYpdCIKa+C6eFMK6FhNLBk5SgQVF
qC4B9FvabDJnmguTo119qI9+ARk1TchaConBzfYFO7GtxLgibLuSmSeztbbp+Mb6FVu0Jq/jy0GR
gdhYiwAlwzgXEDgd87oMBmol4RqHX+3PXCt7k/lSbaayVaSYzh4Ql1DPvqDCokpiNk8tG7XNw2Zg
lZvFczNKZge/f7pP/R4UWfRaB5dqwwMEMvdFXeYYfMo0FX2JM+vC3hv3xUaQ5TsKt7gbSD1/ALB3
rtTB3I3/5gJ6qjbkcazP4j1wOQTfPRHxp/i428X+JdxHqJ8jycdCHeZM47/O06yQlU2jYhyPuQ+H
hXHjIPOBCRN9uJapmdvMEF6U85TNAd1iVp/8iBoz00CoCj1WcXvIs46VftlNzsrbJeJQNF2wgQfp
0oNbz/A9U8h3DlKltTDvYeSUTPRcGwyVIDy3Wur1NpuRkakdQTfeXdms3DjTRvl7oVaM7sVsfS5u
lt/Zk+Era8Ixb8ZezSy69KzEKOed/+/R0/dmXmcedQwU+5g7lPPJNdOWqloLxQoC7KgeV1yMu6V+
79GU2FwOLK5n6idJZmz1LIfTFQtr0oc7ROQN8FPX8IfIEUvnxLFyYxgxhe8htcsLWQ9aNYiOIR5a
Plw68T4/PpO5QfWHmtVEurkQVP05eRx2BUV0T/487IavoIAw+rtz9Os9hcodNo7YT/fc9scnPX1q
TBNfi2vODAO0eNb3gAqJ8GPGbuwgc3RhTcaCH8djQbx+HlWAaAQazPnu6f4fYl2rsBXY1D/lA3SF
b4/y4TpOjwOPOgdfDLzgWO/Tm8QRNOxDI6LQ2QaYwuIRV7x35hniFta0ChEB/0JYSs/HpEYo2GJX
ix5UhuAuwAcZNUjzf0XRZ5OmwS1ojai9fhYCMHdKbEqhfF/Pb5WWsVAMx66/FpQiQPb92m6rjqlQ
EBXkThvZ4nHI4gFsXvJ2CMJtQ9rCjLERKj6O6sBT/z437OXkslaR4RFDuKbbuVgs/y/ahJkuwlBq
4ATNHAPQLSaEjhYRHGvKhqANtny3V4pzU3U3b8zxyGnfvg29VhfNKDx3PAyLjrdDvrtAjBX4HAkr
w98arDHpZE12Rm2U47ph0oNdEl6zPfyDv8nLt5s22OkjNAcmgM5UaVIS4JqKW+bIxwR9rI2cKqGI
QSFDJCkgbnMOitogbm+N8odrsHNqd05mm7ibJOtFZlQdcK9fVFKfBlsugtPoMCvIfq/9cFCnuFNh
QmAC6lmBlWLXx/NXc01T1UJQfY7S27uHcpfseIDlqkAE45lnmWm0KhZ3C1YvAOiP4dF8xlBoeTwM
7IZiw/ZxkO3j1fPDaL5toeKXShHIRDUuUfiFbmjs+BFXtQ8dPSyaF4jhTva6py+aE/ZKCTlI6bge
2oLBWcQbRb6Nfn1qAf1S0LnVemRi0ZJo9dSUcw1UaC74UdHOIU5i6dG+LPsFNlM5VbC+1IchjL8O
wKPMqSRDwOSex2wIt9bndBZ3drmTcWsAduB9F8R1P4KW/Z7JFs9X+zXbGzEMSpOhf14mB51a+klm
Q7up5mVwDsQgFJd7EjFm0SChgZ7tfxTyAK60WA/xvR9YoTJWI6YmXHwm+yhLhnEY6nXCscsQwpb+
JW0XUo288uJRgzRFlDCMSmlKGS7g0TsIA8tZUqD7ft+PpZX1voI+NHrhmR+ExgiYyuoVQa+VBokh
WvzQ9K6z3jBq5nNBwAAOi4CA6zCmf+P9Eoqj7AGLOMAmG4j08gpvBsMmA/+R8aM0FTdME5Os3twW
JYH1u5eZrKjSYFqZTyo22TYt0G0bm6o2LwENZMA3hBLShEtOmRKppgoVoomOpfsozVx4nCpwtGNE
pj8WB3GPIBF341Fk07OMY8FkLsfemUWt4uMQtvfB4kJJ2I/zcDjuDb/L52jUjK4VQCy0vzWJi5jx
umF6Bu74dhEvgGuNcxFBKcri3Vps5DalORORSEJtCSlXjX4i33ybXcHYtCtJ26aWeIYGyNsKeaPu
vLAWe1zW6n45SqxzO2Q0G4QmKyvaMtDzhNc4OxGf+QDtnVE+cge3slGMmgdL9kBcP0SPPhA3fjXT
w2x6+dep5yvyNCFUqlLFSp0tP9AuNbyZGBq5LlzwrxjVmUACiocDTGueDDmhgv6rG7iWcVIU911m
7VL9Grt4UEPQwwmJniKjrWg5J0nP4q+JTmsuj0BIXLktixcOSDgA6ifbAYf2S5ThX+4OPY2SuEKx
9YleHBeGvCXEXXiWUeC5Pp4lGoUR9DTh+5JXAqPpVS/yIjhCmUqZeImFI8whf6hTnemADzC/eLeC
uEhJre3n/PIhqh4s0KP2WnAzgBd2yjfnNiEqrjumZNA+9Wrd1xeeV9nEY5hYJkzZ0t4qoylWMaAP
jokMVplEUFvStklpWYjyaOcVdmM5tJHzp6FojbJscXrg7bhL0NE10vaTwYtxd+BeBAViri+dLxx2
m1zh2sajHvzvPfxRugL+D0Hf2B+aPxr7JnR+5UNPqYNQbtnrMiidcMzpMUVEK1n33VuqXpyk8IMN
4grL/C5vYDOgoCUiXYdLBpL07RY4WZ5wxIPFunbpWuHFbn2n3DfbG+YEVzNyRoc4FTGn1fgR4nJF
mN0S9j4DQrNhYpJS+JVrQmuw0jjL5rICzKD/MArQYD2C9DMXlsmOLkdxyIARRY3PHHGmNJLnemeF
iOLgqxfq/8xu6+JDRnxuoR0pFwgnvHqAHYsj3EhkaWhjmsrjkAEBXiBdEqyUqiy3YYQr23fPW70y
m9LjSPoi6Vw/1ChPA37tZJgvrCq4lbQoJMsg0vrJXAq8CnbmXHvg773j49IuUKk9qRMJ06kD0ZrD
7ZoHFGo8/yuJT80aHQsDjSFBNHqfavgvwglG+9abzOK7HxUHDa7EAifyaIQr4hJXxsdX3X5LjC3w
v0qhoxntZD4CFD/L1N93obfbaxgkFYCxqQuPafOzPDUfj1o5DtgeAF8fpgb0NX7bnhlcNyBwzYke
20rWi+g5HnTIgEv0thSHkwTez5WkC40vpgM6jo5Z07y4mqC/um1LJPU4lbWk7/u46fzlkaDGESUW
m8jYfN5Du2vWhyLt0/saAwpgme8Uc3QCC0IIzfejVJnLebsrTU17oFWx7/xyDwcsmHjRzTrNwRJD
3lJ0xLXGfu3rT+sIf0pDfvBOkyGzEu5xYMKyyM3CXXBM9oMHoOSmmYaaSFxkXPa3wkwGCnMpsUcP
CMjgvz9yXhzwx+dtHcvQsPIcYVLbUyW/THvx/DAc7b23wbl39Z6rcHsa/0zADQ8RsXbMfTUqSrC/
7KNcJ1FNpSVzpibAbsGFf6i29FVf1KEVkbQy74r2tFAW8yyLFBeEO9+TV4tJfx2d55fC7S4WDZmt
hAVJHLhKkZSX4IXSqeVop0Dej8nLVwvgXDrB1wkrWJyYq3NHwgSJzcW/J0fyirbD9L1mWoJ8qL6F
Z0mUqSLJCzLlkWzUJ6o1IzQH68OSZJNb6CtX8O5PgYYmNPzR6xS7vHHXGbDqBpB5SsPhrVJtEZps
SVTK6QX+QpAK1JCkWyqjEMq4zM3MBak+6tQnBMTXk9lCC0gl9gt71gn1lWPElHr7pEsOX3W2JJYs
Ygkx5tuAVRkIZ/bVzColDYau3nnTUB6dnT3Uq9BXQZcNeOp0YidS46vOzIk+FL/djulth29w2QMu
5bGQQanRB/MAvr1VlBnLhYGPG3owoT+JS+Ch6/tTLqcX3P89ic1Fc65wWZ7GcXOTQFLOwLTDIvPz
rxsPAWp8LitnPBEzmbnB+XSms5Othn2yWovkIBtIIC/Fe9ppU/woQqMqYJx2gn4i5wmdu9aEri4o
942xecdw+K6Cf+JUgm9Tb260IVRyLfBObuzhJ215LIRaRoRv6ceB0jh613xBPZJX9Ie6A7NSG31F
drfb5BuhYTcYW157UAtFonlSvqlvJ38SAmMY64CK+E67x94XTfog0QDkERX//28XY3yZ0ae3ETVm
UJlB6o1qghrI6Vm2rQv+LZf3j958LtR5EBUBkZMoCLDP+/r/x5A/PEeEa0bz+opHUCDmd2n0Qe/r
gFiVrog8bd5je5x7BH7e5tlL53aRfyZuths5V684dAhveoQk21UAklSYxqGAL6NPVQDd/CfZHTuv
MRXa6qD0bfBQwg9JjH9tLAjWu+GVjKMGHq6BLQs6sjHmhgVaVfMAbNt68SBIQpBwQD0v3CW7D1UP
ITdrxpZj4mK9uBURA+omUz0Bo/BjwdCE6CF6NoiHBZAAZoe/67s0f6nQ/RlU+a8D8oFjKmVcfp9k
sJ12a/uGzSIseKggOJz0xhVCF+fnEhD4pa8lHOrNWJ4N0T/7bnwHPwI1tK6tUWoE6ON8kYdeCuae
Wae1gPCARb/s0wOY88YPGVe9dpY3qHUQ29MACIWYrLe9C7AMPoeTOcn01tpJr36ffra/94JBsdPo
ui2y53psmYy0pzOxdKo4XNLwMPZEzRuqQomPfXmFzmQy4hGP6mbWp81wjHt93/a8c21W1nSgHmjE
64LjUS6lrDYAfs2qWhjJyk7UzvbdOdtx61NWi0YsWAEVk98wlGuhowXOKe5VVF1XJGh+aGu9rxSI
u3pe6uLApoXxcEvE6zhTjV7JdsVdewmiI7BTrohyigdJLtFsLExJgjF3HZuqqjsuy+urm0aJOjQT
nJi2jaMz8OK/ugQngprFkj78pM9vKd9W5Er9lflzdkaeOZIvtp9nhc/GA8DN0q1QO+CfcLUNZiPl
2I/Vx0QEZh9sF38wNdYKyH+xjeuqK4NrBtZu87dFYUsqhGrcMuPGqQK+iK/0Y1fnd7yLvyLMi5Ej
ograUsG1fx7SnTtLq1dUakVpQ9o8lwZnDcYSXgNhe11VRlGx5kM1Z8HKKggm8Oi6VgcFyi88LSdq
lgjpYzFM1DbU4zvzjcpu+bH3pE+AvOsCOYx4XsMkW+mRuFlB5vHwrkp/RiGB3A/euyrWqOtMOWVo
aOkXlLgw1QDsVeutdDYUb8ksxiCufBZT1yNBq2UUvG4acVJQdDcwY02ZD04j0qEPs2aHWiSrjibN
eo8dySFpwe/wk2l37nc/r46Xk2W26G09JGrkHDiw/FVNlROoqljGynnfo3fyyIMzXjJ6Efy2EB8/
9e7GEz2FZhkfedL7198gGkcA61dXJy4O87DvdltaV2f98zXl0LsCGrWrwui24Y09gxx5cENf4pIE
mTTx7a0yHdeOVNS17mxFij993rn7r6XCnfygQFvQx7MevB1wOKeedw7IPUWyBoNXdTFxStXcSN1K
WHrAaFtSCDm/eikEHa+GTsO5bklf/cbl5zK3CiOY5pCsiYnqoHok9DBNcNdCD0P75ansNCIN7n3m
L2V7RLUBHi5KVBYSToObKmQH3hXb6iBX58DYeK8NJxw4IVcIkgXimVgjTLDQSae3//ccJufUnn52
Q/1Rw98XsiFBmH/YCrbC/lCUFPl9X5fWlFnYIgjoZCNGwrArq3UT4zfuhQJPAvx1HaQ59m9HUVBg
QqiagYJW3vcCSNlsd9sOXLWS1dAsSfUXo3qHmLcFdEy4Llh0JZqp8NRAglETL+w8gU7QefSKYg/C
MdlE+vAwYYSehdiwZzQjjWsLakanuPCttRsCe/f96/M1evEBq0wgTe0UzrZA8XkLUakyHhHsr9vd
CjgujDcg1TJx7KXhofL/+0PzY14uKGKPtI1pNoyyZUfHsERjWPFpuDyAY+6V2m9XgNulEu/pD7yO
QInrfaSNqJo8dshWEnmRg24yceeEEeoAkh33+kERMgQpU7ptXRNACuKtZJ1C+OdDzk6NQZ/ziwYB
fKglOiKi7ydxBm4AYokUvHPy2HdBlIjt2PB15CuoAx1FKjmPpPlfk8pNxJg20TuiMkjigd/YRQjl
66gPvzRBsi+NLiVdq/zTz6qXUoz2MU6ZlZVjogG/Ol4ReUGiS3pmpQC9nWJaxI9LmuBp/Zyg3kzV
JkFi8BZRTuDVKlL75cc5ANIvO0ob0PXFMS1ebw5KmPZPVG1a1PRubhS2Szt6vLa0PEEb5KT9/bak
BHSBHb5xIX2VxcL1qwdGU38o1I0PAVsIe28o47CF6JwrRCQG7h19L3GRy/LyM4Ole3S+lvOs2WTm
4xUKCUv/NieQxqadP+ZGrM+7xYdNTwJFhCHIGgMA0SYaofoLAJTPxLW5XAiz2g0ZXHJB2339ap18
LoFEzdKAH4rHdrszD6TD91lhxyadM8qn5A4jQCjvLpVPcFm4iatEaMnsT+BZwky9itwd5CpidQoK
PVReYttiyzgoA5THvDN8C+aMOTT+4eYpsMRBM5Mf0BRuuE/56ojOpMNQXf3L8og94+PSSndH6GCu
8zb5eNYiFjq7pZJ1MTO4y4Y3VOMBtjhgOS4g+AHdf7h15hm9xuv28/T96QexPYNTAT70Ua3gFqzr
H738h25ZleVwqBr1Fc2RMZnPk7FveIx0ylJjBSOokouT1ltklckpYAn9ZWAQOPr4wvzEqi3U+F3F
yJKWhXzHWeU+YToQ9jpCrPy1Jm64YlHg3FaeZ95hd7L/4ffjYp/sjpMUoT75kMiFBgbxXOXXr7ek
qSj42W3++95s2GGZqYiJyHzGkhmZMU0UVAeK7AmJBoXZ2aHHwjql5t9Hm2EzRmLymj2JopG1++Mv
atVD5c4O5pT9FQcZ8o5BPtLqVhQp/zf3scODVUO6LLayPZ/bfmkXWr2yb/dFnq9IDEFyHw47VQBP
TBd9AzcOffBam2kZY+RUKfS5m6HLjVpaD02IZI0b70nHztn8zawxbEwG91qOgzsPBRLYwUTJ36nV
oBtz3hTMSgxfmoS9xod6zsI5F80757vYz6IyAB+YuTcSI0RubxaJCVTWujjGmEgAao6fFji0kvTD
fle7JoP/mg7jUdEdd1OaIhLs346hqo4IsJFzUIM1Uq49DzgSW80JcNsMuMtMfeuucy+XKwOIjEfH
dx4N21tyo7i/96Pc3kjE/MDO+8Ej2GlAGFofeWvPuW9C58FwgKpsZVwlB8PrvEZVbvef92z46rEx
Apn5GN/Z8Mz9m9iZZGOP8aECBwKbFX+UbsZgQww1WMiC+yyr0kQrb4wJaaQbAitfpycjn+JbW4Fb
HizI76Xj3IkR+AQbwkKBnPuQSriLdMiLon3Tz/b8rHonyheGx8ObRe4lopMxGzp4rWgGOA0P+UoC
L99icWJQmydoeBfyZRaoRa4yBYmwVtlinQliD3IPHSU/mPOwEhYImpy4lql7GKUdM8QrmIfWtTvH
1axR04kzj8SDwG5Q98ToAYldMmlCEq9+w/j3e0VU1YQJ+t8WKNg5BBr6LeY4K3utn2LlFK/3eFmx
6CmLdll6iW78A+hFPy/vm2Rdt8oUW5yULiv0coqx+HWKPS+xIxUJb09rbOZL6kaYRhG/JR9awuIq
fvbvJQfGCOUBG3Wrx5lWnYbph5n5+vNi9frwDpImT/Of/c+W3yZHz2ZkY4vPVjriDYuOunsfCCRb
u3EJVwLSSBvHv/TVjVvwCfIoJEmLX8lV0fWX6CNeWPmRUmArWBT+VpIfXG+zfCbhQu+6YDFKlgmN
uwtvjVcOOeOGlSCn4fIbXK8nmvNXesyzfZFRCo87eW+5ZLp4U3R3QRNrKGiwYgZ6mk6Gplc7MX7m
dFp2albssU0YyLH40+ns2N3u4m2dpo/OgjCRS4FrAurdfowuddNYDu0eKHaVwH6XwKGtW3+YWVUd
WrlF2rEEfHggmWheQgDSaFX5zPbtT/FX9pummLSVvNf6v17OvxCDMr330WbfGemmxlUoW2lwmpXq
E31xXb28kLKExuVmXzzCNQFRpjlvPszbDpJLlxs6oD2dkVKjgd7Ji5yCzLDGHPF8v7zkdcUg735B
YdL/0Un+bmRSCe2/twpiZtEWxtsdoee3n4+Mjr/dfRpm+9cMCIxnGkqRGFORHtLyK7N4xEtXJX40
6GnBtZqiFzKW6J6taIsGwYAP0dTIAb8cMl9EoqxOW1MsbJdso2pLkahjvhMFo+oVYUs1tQ8Nsdqv
5w4TJEmjkp8y64zvwT9Dh84p3o/bijSKOxNgviOlk3qUEYNs2scVQHO5eLjYQAoUW8wFcDFKB3Gv
DgNRg0CkAlKF9b9Dp+ZyHXSMtmBgNcClfkYOE1qSzWmjVIk2hx0OIR66Cle+1RHcSbT/+/LYxAIl
Z/2SUX/iMXwLVGrJPOwomr6b5wewLIo3WBBOXviWeKYda4ArXUUCuP0DxtzEtaxUA8Yc/Y3Sz1sM
REP7m7Vh/6GGkgKHwhh3/ZjtfTIfRf1AgS/0alyyofsOU1wPVA9oMaIYYt9PuoioG2Ka/xipf/AR
gnf9bI2BCNu9RTgeqTuAisDU+WS6W0bhLOaeWt+eNdNJD2M7D/+dFzUT9yrxsFJnqUIig46LPnOO
3SPSsYkHbt4YgW/Pw0d9i1VKouso8NRng2o/GfmICILIGXbcX6FYS6SAdXT+rmjIBDP3u6y2KnTC
DjGVPHvHObTfOkndZrqvF8/Wfe2wQACvE3Mri3EAwZGKGLRcHFW3jYBLKYm3+TTky1iTx6P4B5gS
FWLKJ/DvUvdeci/TIc+DxxBkLInvVTZXDX866t1tYSO/EGU8v7RpC+5PW2pBlVempbbW4+Tg4xUU
4ih3SfY/FB6Ev/zanT7dT8CJFaJ+Vdy22oOhKtpUVvE0VzAhlEsELYqC/AJFLWxKB3MGmE1Nn+RS
i5TpixEs8QSZVBQ40lMmUx1PrT7R3eEPEbuG20YrlA0QNGhvXhgub2cwcp6eH+wnUIJB1hRvns60
MwwpPNAFfJvh3Zi40KUvFuSpxkV/Y9h8j+MXtXwO5ursFJcYC06rn/PvgAJIyYedvUxkxHLitPQl
ZICA4I/vFgNnc2sdBrqhJA29zFazTXGvykVQ6wm2luoeVYo/Qosdpqiy16fLLOv9ebUlNqLZsGrF
1V20Zqi3LW6bpTMU71nOJZ0yGK42rRB6zItUU5Ig0R6jDW3Yc0GooiPMxmrzK0d6c+9V86QJdxzL
JvzNMiiq5Am58aMIRine4dsJjfCC4DC+REztK0f/wO/aulS3Hj7ys4zB4ljJhgxTZws7ekpA08up
8BVrmI+iIVRbJ+3dfA9ewmq5CGt428g7E6iK+OuNJ2Yu9yoBmnQ0q8wy1tJL8EJ5ulGqrWg7ZKyd
j/VKi7cV9v+NXOadYnVXwNQHgOjd57KHC2zhZhawfUvuQNnUgVTKwrKvIPNhVevrhNCTTvLtG2SK
34xs/qrpzEJny/PTE2Ayh6R+7X2zx8qPO1vlQcWrE9YDzgSAS9BoUDA8D8TyXmICEhzvQsDV2MNa
1FSDshbqfyGQm11VsyrtpTraxlgcCZi5xQxPwy07k0n8YVt6k0Vj8FxEsHlxBzryhcDddujIpup8
ifsG42545ZJgL8Qh7Ul3WY3fN5Ul04nQRW2pv9pg4PN0o+QOvWS+mnVlyu/oP5oBDKcdGSZ6qnDq
yf8vLuivecOVjZx/CUWlQmCqWliXG6CorhGF7P3V1ZwWBX+DxzTjvNZYldPQrh+vzqDnNl3c1qVu
kR2RkKrXpM8Z8fTw08NYfkc1p/Aqkjouo3o5N3JJ5EYclm2VQlzCtoAZcG2yCoxeGNS60cuIwaK9
Ta0EYs5rGA7q3kOS6OfnSRHZZomYuc0Ylw4k+MwPpauHw+j8GAwm5fgXXOULUYbCF6Rq6+V8NPb6
VkRAONWTpQ1rKrx9A5DPhHLnFpbHnG0SN0DUq2NzmbEAc4rGIjTBdq6zSTa/VCecUpcXc6+eUCcC
sds5dxrHaMEPwmXae2GcQlZehuZZewUd9FAnhRLFp0S1r7HY+V0g9OMYxYnM4UP3XnPcjjGPT8AD
0wASH2/fInMgYHmuFPmCkmj7FBWRZi2wYdBCdl12ktCoglSxNsXyNlHBacXhtz82KiU+2NTLVzaI
Shato7tmvjdMDYuyMPYgsryCUJemACjQ+qwjc+lsXReFWrurvQ6Yj//O88Wr3efLg74o7k/a//Nb
QuB6BeCECyLq9tdY/R/ivHQJFcnzFVwvVzreczut2S7vF7eoy1aSg8hxc4Ow/V5EgrnPJ2mYn0Jj
PBfx35hUmq4WDhybSv2ZjbOaNo3UY4RVUbuwwzf57DGD1gzDgvZVqhTb/dx2RRb4J9ucypeemXr4
v/y6e0F+KWob8yNbNYmqmlzE2/WUu++Hb7yf1tYSChk9V1+RxNzIN+rjZlGLj7IjF4ao4xSxaUd1
yuXh9dXWh1bgpxQirM5RGeK5N1rATyIxbEweMUaJCIPYkFwSZyoU6xnqrz2/txcdMPHzKoKVuUZo
nNWS9hp9YGaKIMvx/0MDxrW9e9QeDaf83PtFnsi1a4cnjHWWlWWyLzW+zTk1q8Q6W9oiU/MGt1tO
PA2ZaD/hl4kFy3clT4P+SPOT2NuMy3xsB9ZTDmxRM9E0qfomTKmUXx5mrKGa0EqeHdhSZpx9bRwu
afAVk4KZsJTz43ZAKyUhkBozcS9RskX4WsfxaiggmyygRQnS+7+8VTzhZeid7tbMZXJfCnHK8WC4
OiOo2IYhnBPSZ/+ZGwnNF8zcQOJdHDMo5uUa175csRoeiaG2xMyKC2UCCd4OmRiU3tWfY2MeUwk/
JnNneWCO/pvakXvvJzKIbpo/7V5vgk93QQN/bTc9lW1QyAJZShQ3DNgYRiXPwkOMgGoYMfVl0oCS
vHT9TqHw6al047XxhB1ABoOP4pBLj1HNM7GA5TxWQlVHtgelaMrKtUmLeS0yfE8+8GfjgSpJ4Wtg
ls93gwMINeCGpwuWzHdFndk/vjDeF905pas1SRYjP0ZU7xt4GOmFjN5AxOS0qqADULm4MAboWF28
vZrSBlVbtfDJC7lt0GUctMNFD0UpdCFlMqGbx9WOjquEmBOuCnEN/s4TxnUnp8ovHNReIwY8L0S5
6561mKuPhXKeFpmjaJ2evRk7RW32PXO1Aj6yUN3uO0qc4eMvVLnhDMq/J6PzI63Pcdx9glBw6J13
NSuEfGq4Zk+cuPqPd9igKoxGbmAP9KwSRG9hig7jd9Eu8Z1HwGhZqfCJ7nVtE/25gkTw3Alkqu0f
pMcEnj33vQrUcJPbFeqmyc9iOR2kPVsXbt44HYRT7EaDJCUMrNX+sDp8VqiA4+m0y/0JTG17h6tU
/LvIE2lnF/GUsps1dn3LZD5v4uzQEbzhHus2HeILmaB9R3z1ZisUd6BqH8UnLjnLxbpTkKdrL1qG
VaSLwMZT2JoqG4P9N2/pNZ8giZIToheqTQvTosxYg4uQVzg6k7Lc48i5A4FWb3N1Sek22f2AiXoj
3xPIuycKocltOANOxlK+HcS6EJIy71tP+iaCUx8EklnxFF3zL+CNGj9Tz/abh2oa9RgIkb4wQjie
RGiotNsx19ntO0e46Od67EwpmDy4cspZREepZXD3Fma/55cxReq27PYjNO6wxydvslAaHt6RDflh
YHVFSfEcW4rYKb4kPwPdBMLiztdES63IaO43PRNfhIzoY014UUTJ/pppjdwu58NTu8BHoW//QU3J
/kpI/lOndR0ETjNZAYgR0J/Bb50tvNrPQ3i5vLbsxK1cdPg9bAC5Ws86sask2rVYkxAOoJ47E8MF
KYjW2Fq4NY6nNVQjVtbsKUnBXMVIDtqCZMLitCVd4b6fPrnqxn3KL0nZp7nFxvunO1pk9XS+Hdke
Fhgk8xMTerpFtpLtTMqwB4F0P6ktVoNKhTmiIYizL4s372IWla4ftlYGfUcs9S5jbMhSWYbgmr3F
NwZ4znHuwteyRP4mgNgf+NAvpzaoPF8AJn9/A+AqDp1bYXQovW80zb3P4p19erwzpmhM1f+GyVEy
BScV5/x+O8IieWeMwnX4e9MDnrOz8/stfKpoP+6yqn23yj8XjQyc1mS55hYp2IBQiiVhUAsTjzoR
Y1B0Co4G+Dv2mThSnVGuIiXzkpLRor9EbnTwKCXDw4nw3SPlxi82TM9UrZtZEip/u9hDhIxfLAE1
Y7TgHajx0vqk+Av3/uDrSgWex7NlwR9J8AKbggrPIuQ/lhSpyrzPYRZCCxWpUIRHsjWFF9q13Giz
7akgaSnH5EnTITQFfwMKVu3cwoQYKeIRR+TjNjNNZuTSIjKUPH6zsrYHVKDIoPgxdF92WDvs5GqT
778EWuJmuX54m/YRrt/ttV1cnmBANCwRtcOTftiVhR9Guc91O+PeWXP88DCGhfklNftw+PXHnmzi
JSahSiPCtWXwg27+UWnjGT3tDQ/TBZW+VA0lkWkkZvqi6+qhxABMMgmAYW3ZCwnURBap3DNAVpS6
RodA9UHEaKdsJr0XfB6oMNDkXu31eFVxhet7AM8i5Ue5pyyKQWZ8nK43wdlXMQa8qijs4dpchjSu
juSV6+KFRXuB+svstcoHVV49kG5a0yfOLDqY8kLYGcoOoMuEl4EDwjrRl3DFXTO2Q85V++wjWrZD
Ue4AMPPFfCebHSLQjI3OOIUcMSLgUUnKQHZ2e+8H2me9/k8MbXviUh5RFsQiQqcE9rLFdp3Iu7w7
o1eXo8L6LNMn+5B1Rhizo1sBSDMC9O8LPa3X2UUQd+lf3F6TftZYVZ1GSlBEjY4Gt4ZYO752c0gO
61mPefINDV1kJ8+yExAY/SdwVccJqJyNCFNHlCQcYbP813BT083pzhuYykBcHVbD+eKmoL/ENH5y
W0HG8JIZRXbqZBUi4ukQfAt4BZRMmWCDY7m0BPG6ypt4SO5M6MFLERfKQ4Pqt3YnpH1YwzM9Rqqr
GhotB4Eydkpv9bv2R1wHrQeyuZL5oSyFPrfL3ZCgGgaob3k69lnB1mzAVUeNbc+Mm6L+F1VDRphU
s+hAMjlB8Rv0L1nyiGxuJiJl+M6c9+Wj355SwhfwqoVRSpr4JaJ1rsZVpGNaBsBcdue8/JXN6pLg
UDr1UvI4yGfF27VxVq7Gy+MmMFPyvDAiXQL3j2Hsj5LiErDqzdikYkZYFiX9ZqrJ0C2SnmLNUELz
7a3z+nBAA65S2ikrshLPsk+KA2wxZ1kzomiocQCXbi1NIIvkwrpdvqLLOoTVXZdlrfzCsDrTyhrd
xhTVTQ1uqkYm0vU1/4rnSOMTP/+M3eJ3vEUbVp7l7eDrEgZKC2UM4drRtQVepSA7NqR/133JsQUK
AN7BPtnM9LBA2nQIMTtSlVlYT4LJ7Ke8rzTZahFe2h4+0bgv9wKZ7XJewTJdATBaYkt/NR9SJXNV
Olys7NRirCpy1T6G5mRy+4IeJ4QdTOlkGicRaiS8noYza57g+kf9mJ1RyjaGdN6mWCH6loC3f5vE
2bnk18SBsXYEDcfJDirDbH6DDsrBAQD/38y+aT4r6v8s1u01ZCpudVE9hA6iI8HyhiSJ3nLOvftX
2d7SZgivXbQyERnojkE0Dwye2H0GQAyYSiHkQasYWwvP5E60BuWnaoFZE5BJ5qrO8G1XTgpvS1zG
APG0d0TbBziDHl8sgMTUgF2WbQw33P77xBWHDoLZ/q3rsIxfaMcoqwaspyN+LPx6fiWAgYkDHcyX
tFrASkgeEsK6vhTScAYfwWdv4kBfWrQtL3P3VmFHnqVPVXYspQ8i4W4xjQzbSDJCMJs+3VNSns7h
3N1P2o1oceyw0v+f7hegxrUIN+U9jWG41H9X6AoHrzD1KdCabPBfQ3LyM6E6Mgy2AYmI8WZGZPCk
GWS8kVEDVYOBxKFfsQL3F5skc+q9s4dPcaf7G5up7XKLvNFMwwwyOQTpDPuIYkd7d+e5p52ODOwf
+v9PfUmatYa1rp/OPWsIPWA98MW341e9jq/w8UXsWbZ6JlU4YebvnjikkzJKMbpTUhwHCXjsO6VQ
CFlso03idzPv6+pqGTeyyqhXCMqjEP3AXxEYRO9xKDKZGFiiMrV9qGu74JCgb3trrPyKV/7hF+e4
/n4yOL3+LM4TvPrAnxZgkmz+7Me01RI9ifrZdkBiW0zLAcDg2YXqD0UzkIdpK/AshIBWIbk9PMVd
64C4OgAlsiZqaQsWjIVrKIiPvfcibM05lJ0qK2RXJU/FlIfJlKEH5DpNEcc0MSqRnlTl6YG1q9iN
Qh3YBxzI2/vyRSuSz+BWWJXGn4FwaNjZzdHEF/+iS3LeIV9lR3sfyUYZiP0vJgPS/MiLpap3/9Hz
vGqWuprVuA6UHJ6keQUXNAu6VQWTbSZIBTlaeN6EGbSUv/ayv66CsHJAtYSjC8Q4sp6XswRVbof7
WI1tsmqZr4FOt+OPY/AHVAuvoLrC6C8x+tkHkxhDqRu99OeBZy5d+g09MdpqkVRVD/doXXLqNAiP
t/xI5zCcoawED/74oQaIgTQRqdWyDsszP9IJKsrxELUkNcdkGfxGIPGnQlQ4xNJDhRBqLS/Uac9K
Tu5xDrtywfONSiOz7TRpgfhNHPiBAWtdjNsgIcymJdwgsPIoL4y56ZrCq9LQo/qmaGCgcnDIIFbM
A8dZcrVV0hdH1O4d/bsdGFZzsMehfACss4nkkXZW2itB3aG1D+rxL23iDK0f5/066/gCfVqcO/ym
sSrIon7GlX8jVOrTfFJLKOascSJLfW4y9K/1srCGymhMaHY8cZHyB1PHPEJeDlFU/Oa7mbkWibhX
1ffTQFobKm6Gv/JKXlEc/r+EC72u0VTa30IXaN686MPcTZs/mXdbwn6dgBCDApJoiL7ONWeU/11Y
edeliyOqRNqILqN9TRiJ5QIFX8zx72MMOYpKNnw4tjLnmo2N0nKuoHv/RDQf6BiVIQd8JNOXLNK3
SdkHy3qIZDrNNCPBsm9zIeldcmz18yhR7gEVIHEQ5MN5RuGxuwWYJquCghUvn4N7xjL1WqMlq0w0
z++R4BfkYcpCjUMGbl4Ta8+B+XELFG4NAdx3HofaYLMOCIjEceuwpxXFP+Tiqa87wwWViDgTbJEt
0SLdHuiIqfDKazsvHXMj7OLyUZ2sVUIkx+JKQQW1WLFm8YYUsGAXWQnkGM6vJdZkLncp8RS6gT0X
J/nUfUqS5GFhnf9MLEUIwnfiE0KRXHWBynVoYnHQndE6SLi1g+y7GKK8djtZQTvRfxcA0d2/y7o4
zwQxgbmtgpUNtgVot2fLLXMCWNDEDoeS529dpnTxOLOazVabkskr+iAms9MjTdJ6oeeSQbt+aDGN
RlSy4KXmsgx4pbBEsMw3wBDi8M0/g4XogO6c+dp4CxCvYDgF/5H8OFf0W3BlhM1AEizXk1bP77wI
gxDRReYU7FLxPalLXxI8aGdPkregGRxOhc8jAebnLcjzZvP4oJwaUqpZSoXoAhnjjCb8WbmzEyOD
OzZGVXjirPZXGluhgTa0XmKzDKiF18OyMUWIwdMvAbVQ0kV8/z4NmJMfCMpqjpFLIkSSAzguJG7v
M6Bkr+F6xAWV+Cm3ho0DKUmTFsExU8gbDRSONs563rwpMErQxqUUcsywBH1cdufvFPQEuzMiYJrL
PpSf+ubbSnXhVwDPqYWJv8ke5zl4+fdG3HdlFp2yxRc8MHiWIjjMOftK0HskWWH4L1XgSjCGiFdM
m7ndICAHUmNb7/KbTxsc3ccvouGNkOR5zsAr7PlLFo3Bnd6q4y4xFZOJOrRIyx7G279taKt8Flpm
VwvlFpTGyyv7IOj27sSD2vZqFIF/1mZ0A8/YZfPNAlnyACAwCz7dlBDlMtM00Sh5JaXV3xo333sB
9kEA2ndMyTKAOmsb2GOMXzEic20Anhqp3zWqBjdAINKzp8i7DTXegJrjghWcy4P5qljzygWzNba2
DuHo7YXnMWnXaImqKH4vnJt+pSSAZOSnt7mggRqdic0na4EXHgMk5OkFLURizFfBM4cDdygEfZIA
J93pZm4/1SNNICQ7PsbMnrM7Riu7+l2zT5vhfB6G24sTBUAuZBBkYwc26C1WzC99jDSOuFvLDtuB
cgK7vXCgmm2AyRQXjdf2OekkSHtGelxIK+HJIg39Dsf29fWHJycBtZm0qYd/NxfnmSrZv7JcVfIm
2My87UZO61Sfk/Xs4bf433giKT21WfqA1bzOrEKih4v3WDgweXfWmvQ8EJjMLnBsyNy/9PyvxVyq
dUur8KGovo3qchrjlRwoTZsHlditEx6G0CVtbaSI1HEV6y2gzENmC6MfJVUS3AMJtGfASx4RJEqN
hL+zm6L13wqpnJyFVM+m4nfqEwIbhuSUe8w581PIBKBlqgvcHl0MyOqnoIuAg/KHXzbvTgfHd+Bp
juiM2zpRWcxyIM2Y0PIkSzUBqJs/9Sk1aEswrh2h6W66r59NwbCfo+Y8JHg1eVO2kmLbRqygwyQQ
7Ozs0UZtlWoQVPyqDp6u79C1k1KSI4pBQRC+GQqO2QQnx63rlSr3+YQGMec+73beg9X1nGOdqv1m
qXB1Uv4gWnHVdgXuuhSgy8RCEdLGbxe+9a65TPP69JLUhwPxCHPGrq1JNkMUTChPKXxhdennr2rK
soeDxtnXI833kIQw6S3lufiRyUFJCQzPAntabTRUVh5cLC6yygIxGqpqvXcFC9gS5uB33W2VQAta
BKtDdInKnWXStA1pL5NnAJU17GhjyCUUB56zuO9OqEUsaK1DIWgiXLIqvXrXFXmpj6eRq092o3QA
+CG889qFomjp970drtaR9HF0Zi53n6CT6faQ3z6pnE5jtvJWjtlo3GPe1SVzQeCVu9eqxcrpHh0Q
dlOrve0HaiSoek9T6GZdOCOd3UQrYEXlGVANQAHD15vo/G9pDTYHIdQ7NrILSkmH8a1EVn62bJ4V
DbOfT4S9kko9iJMcNGEXvG3+KgcKNd10iRQMPi4Bt4/P9N9tPVU/jf0hGMWVuKigrqd5h8XlpBI5
s1VxUZiUyLUloiXqrEkiymgAn99TPKxTs/0EalQavj+s12ZwKy8ZnzduA6xan9zRQPNthXdJFWr+
J8lRP2L/Orxdx9XQfvGVQModkg7eBfPipFhkPWe4AraCjtmHCLS1pSNmwp5OYYgp0n7idR4Nu6HC
wnhtn6fXBCW05yCrtW2as9ZsD97u4qK/R7nizpAFoRID+cMWEwxLWCdDyB1HKiV87Yu9frAenAH2
HucKGr2cmLrzXMZl4as0nWO7b+K9LkZ5BC7pf7FRmqAFv5I4TRj6uqEnzHJpavGmfeDXM8ACfjWU
233/eqf6MneTztH9VAzH8J0wvbecss/jW0wDjUYHk1wNsZ4KW1zR48ahAK4EXM4mWBjQ8Bb4axex
VQsDEKMMWBYM/6nj2IXu0s3r/ePh52f9oUd9vWjxGVZoOeRLfY512TcWkpBV0QTTiCsnbtz2Fbbr
of498wroxXW1obhdaZzQpp7MXzS+xUZS5+pPM9Gm14dxtR1ObDhCBzLWLoojxD5jlE0dbep6zxiP
tY1ThEevtOTmfMAGCDrQhAUsKp0I+2NeO0t+iCMhgoVFPTd9CJlxANn7M+r4/WZlnLx88NaGNr9c
MacbiWiWgrQGcm60QcBUP7e1YgzIrrH/LrYIFPfvJLNf9bI/eURmHSGNpo5a5H72wZf29OB2X48g
sERYj31MS680YJZJ3jzkNtJg73/dnvgRdSL5wMNzKwM4e+TVotvIsdV1d6M+9tyymdPtW7Tj5ZXV
ZGjgcNVUVYsHOdMTxXCOWNG1Ie+S87uIhieMULzk5FqDKv9iSNnwi0nx6DqjFH3qKFpOdHdRdp0M
dwAlEJzXoU/2+m+C5p2kLs/5EHkE++B7v9/mYZoPFji4kYgANqhKhjiEZ6yBNAxQNGWUjQ30DRWS
9AbquUf2JtGHeprgMnZD0ToVY8j7utWoEbmFanbxlf2z6i6jlsfG47TIR9YPoeeamj2yYRKE67Q3
cYdmsGQ1AMvFhYYJmuvwyi6qqhpF4rU4MGjpYOy/baEKhV2xVTP6RDaCGUhNigTaFdvLHxKq2xyl
dQrvQr/Y6iU02vziZtYEvqzoDd1o+s2gyhH/0JqpdRk/VpAMqtQ1pzSMIRI3pPxFcyD8enguEqpn
wDA5yHuuAm5OFGAjiycGJQmnp4yVH/lymQSikt6fObCx3gRSE0BFgDrWL07VVhvxWR0mQ8ow4qtk
2Jlg/hQnglZMliH83H9YV6ZrZiUJicMlLH5EpFHWyy+otWUUgnYGoei3LfYbkBKMIa6iW5f/MqNE
7hrWMxqPltztkAXQZZAWfUvGueNB+x2E2IGu2YZnVnYdp2DCdgqDTuKoXL4NOi691oZ6BCsgVMsZ
DapxIywF6gy+afDWqL99oibn60G1lhtd+D9FaUfwIgbya15lFJU/p0AfnK+26dDDnKX+y5pPLl2n
7rloxjvm26FgOhASG8cdEIzeXEQuv4K10sf1PJM2XUHSOvqm3i/wdXxz14QTaohEEDlYktyDlaVo
mux0BNIIVd2mSm/P0F2D2WQwt1n6L+zHCVN9YW/cA8kbh4bgftlUAf5xW0a7qw4cvw8yycgYMRYK
mTDhi0NeeUqdrCqYR/yai2QNGr+Y64vvR9pkfkEERNB+usvmD9QBd39FekiKFG301kZpvVM0d02M
AOPH7mihJfQce3y9/arkmRDWJrqulcsJ6/Si4eiIl9ED3HeGdEj/WyKYEQPfQtufGdZbx0L6laKb
0HuiBmaOUvTG71bUExbJcP3J30hwB5MFXOjobZfcfBznPYdRGY73b3j9uOh1ybu+D9HM/JhrCMPH
YjnWK/OEQUmhovr/ZsKRnr1752njVD99AXfvmcA9YVHz//Lvwn0Ljd/DZYbi3+YGtwHiTKQXV1jv
pgiMQdfpSSLMi9ZzNMbEy+oM7lagT76KsSuFdu08CvPwqm+x6ey06YCx1ETZP9pwflgoFjrCQkvK
VdmXnTjR/UNLplPsxYx6QO3GleZ4+kqqZgn2l6ylbyRqvucCd1L5y/ig+0s/G/7Jcgi4P+6lCcDd
TRSUIcKqP6ERMeNNQRZGmaFIYWMbPWvlJZBhkhf4Bq1MSkcRX5ka5mgjqK3frb3tHniSYlDPtj2H
iLbxo5GJJC0589vsnlvQ+zzQYrRLmRRTtJHRWjbJtwCn5mjrES8Tl2ZighIJjNYdIQ6IfCW/PHWu
70Rl+dVWPreyXMxtgEiV3yn6f8KFv1/0TR/uMFfKRqB9BaZ6kNcoIQNKh2UXn1nD5raxO4vUmBoV
NCmOC4BNrjp8X6YVBzko8tcuRgw7+udKE/0y57vJDzXQ6gd8NEzcPQJufMlcEcq5nvS+nETghYMg
6rQwUDgAHVsSe1aTwCuiySvVb5TGawDOu7ms1AKj8vKhhtDzyLucT2sIsyXM5gKUX81lPKK9xDzs
J3b9VJxzqK8g3N4RwaoXkGgzNeu6WXqSfzYAWJxCYaIAg6BC5fhD8+oZG1azoHAIdTFMRf1c9oBb
G8xuZzNXqhjxxTs7qJUP3HvEt6OJykOyEXY+QytrY2s+B4TvnLo9+zqdX1QE46/NVC2UkkCIaeuM
/2oet/M/SrZhZNVWfp0OZDHYKovMmEz7oBZaTpQulGtLTVpl42lBxcUlm+UrbKX/vu62rXaUiPcJ
APpEStfDx5xVFCLi7PKjidT0ARkyXbS/c1qIUsMx0mDGNuCj8Tne7jM8KSldSlL16/K5UikgABam
3tkDBCdDdrzidNilIl1d2MzXimCAPe/PmYvJWjNI5/4ISzU//orpLbOBjU9gkWz6zHcsm9jJ81QK
9u/WYw+yTTGGaPOFaWa1IlCyBQnsl4HDvkTeyaELDaeaJOiKG+OoKbkZIL+361UtyOzFi9FDbzAs
HfwW43pFYxLFMpT+LkWA/Yn9+r/GKegIZwrNgbNh812ZUScYvYMqwced2eFD+ZvRcfKwTtsoJ/xF
hCF4idFNQCljftNoIxoxCcHwFxNzYIXN4xExDdESxUse6VeU6sGCyrF2wlu4+slXGLvQwciDgvFv
GlGmZO1mvjhyj5I+JfRm7973GDF3TUmMk9lFEtBXr9M5REkyXhp9hYjzy2m8Dym6wZpMvNy4pAk5
cZRxzk2ZO+yrOfnZ4FkDvZNss0oVBX3O2CzELlnN2gFaLU10HJBk3QFHjkczC1N7dEXUXKB0Ov5f
V8ASuXrpAXTbELiKaSWR/EnrOm5shE0hlyJJ0XJuI0GKBlnRCbdvuLHsVH7AHh1Fxc03zULjZUuD
TQe1ikwpn+NcSyIKGCIK5o+pDnTnpTZX8HZm6aDb8ZhpApK3d4CfRJzNjDBRWGhHsb8qy+i+IGIV
sHyb/YEbt9LEfafM8KqHOKBoW5W9kEMj1PitRZ+fBRiK/4jqHIouxY/nshNr8PhrRJmb8B4K99A6
KkYlxRq4VjvuQ0ZTBN0OypHeQJsh1SQBwLehxSoMCAVCpbJe5oQzFxd/8wDyb8ZYn0fL7qmWYzCT
9kwu/2NuFIIfR15axgA2i7OPyOIWqdy3G/KyzBzdpnPrr0IDQMq03sGM/B6NGCLAGNZ9tTswCNq5
1xA5vgTJdflEuqMElVQZuGiIxxiza8kgxiRlrztS6ffhGTrdgmrwpQ+b97Ziq6EGjECRpOQzV//K
SZ27A24FaGOXJBkdKEfhZ+OsXwwY395uB19VxBQVjb2qj+uLdywPjjG3F4rDJ5SXzbfRLhXQLBrb
ZLdXKb7xIBWiWkeeOi+Cx+3wYYK5EKCqAC410YthEE43UULDOyKXG+G10XBLA6dnASUz817e277/
BjsTPwUFTM5xswNJbZv9wkjk2w+hv64z0ICwg/zuHrAeGobFhk3OjkBm655+x2yeV1TG5VNnsJRU
C+3PScOUx/Uqi+L+1Xh2BW0FZjdLHqSNKwJoyhysfESc6A7JQG29WpHx7ttU0LfGepvFH5GePV9k
8okfM9NxVTIoWPWY8tSLDQoU0V82u5Xy2UP78hT/791Pp9h0t0eTICAKTVhhmAb+1cd/7/g8znvp
0QQOpWc9PvoyJbjlPu5vxOaq6h+1JvSH82FRQsXRJZdS5uA252Ib6mbtOHDSa3cV+JQjjF79z7BQ
L3DxtLlroXpTP8Fd/g+WKtb09wjgNCRReCEM7UlcnkKo5mwDF0S6zii7klgMG1JhlfTnFhSHFyAH
T4FvbRDoo1eEgsh3MwolBwYdQ7IEz9KeAdleIrbyF1RGlhGorjU7tv914sp98tqSB0WSL2Elpuht
nHRGciWgSrHpjig7RaCFMCYMvG6A0lETztCs8uq3Y9mmw7fBgjMX9mL5nqq/Yvio25jdtX7c2v/O
rRRFJbl8zunKn0GoEvpPnzMQOBX6E0fpthnh/5/Fz1AMe7uv/lnHeDlHmFiHxrAWmZWWBz9TPGzl
KvXNU9onPdVMD+a1Yf86SCZJwBEDkVAiHoR5AjjXUmdJljJnFwIzqOxGp/OHY+hp2ctjbMezV2rC
GB1s1JWUxc/rDYKFGSrIm3z9ZIShK9hQxUbGStqb2D8GNCJPhhf2yQICE/yyQbuAiigvnNIewvCO
JzYSFTtSm/zmlXQou/JQrGBPfsWWnonqQbySm02AwXfbNGFD+Qeg2URnqaLOa+jgON0rd1kvSqFR
DfHsQhZsRCSRG9I4PLeeRrgxs1v9aYIRgk1pmz92/7ArRLGO3FMWtAD2Xr+z7Bmvw6PIjQsjJSPb
miQCiZMQvbV49ZQ1N7kbUA5bnIS8HyahAFhvPh0dim6MKTUcVtWn8A7eTQ1SQ0KQpfcddXaA5LVx
+GJBMmNH+mN9CvczDBQO5/9Htq+IKZwQkt4fOtdH9M+o7fef+gV8HlLa/uy5COS0RfYwKgfsUUcm
FhzdQg5IXyKBG3+S+d1DeSp6lRXKmlb4eLV4TB3x9xqvcd+X/+f9G3Zo6eneWvX7VufIk6hhg5or
zQCD4KrhvdVQMsHqiOapb8Soh5HFqHNKP1oUmYgrIg1Clhv6msXSEEVKmdDeBBg6VDeiGM7nfhWV
Ry9d7dmYFedSUzak1V8P8UvwlbIDxRBwTA7ieCUs7d/z/+6bB1NInLTrgHnSinsTBvhMPFvt5cKr
pyjXAH7b+Abw41CNC5HE9ZIFcINROmZxr7LWAB1+RNNTHlEgSsPoHv61SIs+/QyCkIq1zo25AC6f
FOcXx62YQUH79t9VAcWvoj/vnKO3To56NIepSzf61/6wp0x8Tt2MD3ti9P2L05+LOnXa3VFDybZe
mgZYUJ2uOBV+Fs03mh9hIKSK6HjBcKBYH2+GkAym2mH/SXA8dRv/IWDKtD6jlC9EAgRFXWO+tOmf
Phb9UhRYLlUVyuc9e/aLNst9YC7Nw3aIykFp+Gx/jQkHMyaGudiHesvXtXHr1SwhcUX6IuKDmGyy
IHNl6tc7kt2V7isIp6A45TAvUAhwS7seoEhOAIb5njdxvD5x0yNd3phlY+W4v071FTok49j9mn4+
ikvzNx4dNHl5sbyFNeV9TRBM8yrqn2TfGo7KlmrBE3hmV6asv44ezJaMp/nrGqZP1uTjkJ7jonns
FJmec40HmwAx4efx545HhQYGiOOgUvbE2+ZvchCwvYCfy60gibBNB8f+vB0OxiR06CuGrBBZ/zAu
wcWpzHccHFGgONFQlP9EUG0j2fTE3OyMThZDYW5/TxhL2+b+xbWXRstxFZsj1kgjPLcYSSMZXWlh
5HOXdzLx/XdCzypuEQoq+Clcr66dVsK46ry0q1XxpgEh289e+K6C2Euhxtef1m76uF4jkxns/R7P
rhlvfxg8aChLlE+D5eILsNo3Q3MynpiMAvsztsoyZGyy9dU7mbizvB+D3xBQuZsZKbe99ds7BRdd
9bwT8yKmUDD/RLrSi99qOGA+wf4w9Fa6R5oDSMRR+QylFP+2wMGFKRpZLseBvOoPw5dqDqF2tP2l
ivhvmJ/9OkCNfwhbyCfF4s0ZxtW0HBdXKjoxf9BmtNKlrQZLlDjc9U0JLz098l3+u8AeptYmOrpp
aoSkSOJGQLPOeuq1lBA9NS3TcdI87cNHNPBBDWBiq67s+pv3aRfFpfIAaFPV0WAq9S34upLgkh9I
6hOYLBxwUUN/T4YB1syvcydLc59mB6hhazgMyb0TBuptMVvi4MTjEEOT44qux6c4gwr+tzPqYkXH
/fGBIWJ08kLticElWAFxLjg0xCLHp6rln23YYeVGEQ7/+GDvJAkdTU+ISV2DFzL5MNZJhvaoej4Z
3B7P/wUQ+8Fpe9AdSnAD3BDwc0LCQGA58Mkm4TVccYWEKm4QcsbMBLfgOwcgCSRuBwD2UXvC2XtU
EqhdYfS3hCElBUML+TDXtciOWr4perVZ/QMf0RP9kqEHspqD2VVh8VdxyCohkjlY2GUwAnsO7LGJ
iI8gxY3AMwqJRfNm5oDuIrlJV0twvD2/oefSaAMZMF0DkAuqbov6uarPzwvR5gJVEHafkCLclbX+
j1guXSXylZyVExzgqIGgqo/B2DWMBOUPkz4VylbJT1/wDVDGxCm0cccxR4X5txFXSyTWR7/FYSLr
qoDhZCWnijNSZcun0nJcUtcVRxYPBNKBqNhZJ80wFpL+cfhD2dJmWor37wZn/422ybzX404Vlvyt
Ik46DCS9ck2pv70AoD7QEIqfE8Cuhhh8ImQ0Lsti9Lp1oHqN8egm2mAnjfYJ7d4Jk9S1Mb5+NHdd
XHHfnJgIBd9JYphwBXQVWRLmDwhwdhcI/+FV9gfVYQd2uy4R5bEBba+8cnwJahZzT1vOzHByXLJZ
u6TokvmRPamlg/xv4rJ2e9HBfrREm3h49WjEPw/SQtdBJqsAU/FkrvH+DGs89VSb1cSuezYXfRMg
gmg0o6tNrUh+JPNkeyHs4KrUWzwB1tWr/gSEAunxiGddh/9DxhJO9i9bsxJ4YRVGzQ/mX+fQS/nz
JJ2LUOQEktlMeioQbG26Xh1n0A2E92XydrRUfGWpltPf+c+4ykhCi8OxKA6xm/Rak6hIiL/IJeQj
1TeMnmmmEjCLumz53iSbEZShw4/CMoWiu28K+TDOv9hlrGjd7eBht92UDEDXOL6dLm4Hpofe6k7b
p1b3R85wyLLLBFbh2TqtS/ifjGuyUf/F7OOrawep+UfUC3IJlqngfoaqhXEMEy4U28j1JmPWmY10
jvI4v2Xac0z4iWKial8JzqagPK1HYJXqi/E3sufIX2+8y+VvBRRaRpgdFHwqNxyr/NzdOQkifCyF
PQAiJkpsuDENReMWcHy2pdt2cXXewZSAhMIFGQ4SLk7gW8f/9aMoWjolKZ5Z9cfgwy8ZItdfXSaX
wnQF122L5Zl7kO9OFAvw2m98DYs3jVj2J1RM2VYqXqzSEUUIflbmueaz/dO2xLIQJSOsTaSHLWL5
1D3Or3DRTY71pzsQY6YXbhO6W5xKI0INHCF3mI1nxVeRiMB4BhtWCt78Gox10hWysvotjMMELlhs
nImpVHgxfbd0wIwSqQKVeBwqr9/QxpN/Ela2k2O72lEdE8wnqQpdR36qrHHFvyBRhGiHR6jRwcnI
1J8qpwx06u33SllVah19Wpjfxwhnq23PkX3SJgOw7F9d93abjkLP1R/REuTPUAmQV9nWmS4h780O
fUSZCj7OHw/GANPHqaOKjMgbRe3LlNjMbMGylj4EYcPfOiwIZv72wT+EXDkER/QeH5/NxNaVWz6L
mXqc262S6ZvX9W+QUh6zNP2cLovET/sZTCDthg5q7/n18HExk/jefEXBt0Ii3wqB/Yn9HetZlulw
iYHOx7nqXtnefd2J/gWCQe5utG5PrmJiNdoxwH0dgAsm0NubHQcSU+o6cRsVNpvYZ6skIUrFKD3R
Qy/bXW4nl6nOvJ37wqo9/xcqyHPzfAm0Q1cz5apTwzjMIli/3ftxE2y8BLmHVhRKQgqJK7qdCTHk
AC+QeeYmBNdQY9SPeLpG8iWlpLHEWPqzCOEYcB3RPkJVZxVUZmm+iFO2amCUwec0XnCS2Cqglvwl
v2Mc5RBN6rWcE2yYP80EK8IDtXbXCS5f0S+EtPpL360xBLh5d6U5NdRhb7jzke8+gMjJvOtzQZQM
eiZ7djPj8ulEY9dxoK7S3+2lXg/XYYNXfW7jrotjihDFUPB1KwXcpnAPELPxJ0OzOpj2xsB6UH44
S2DFZHD3oDMda4jIt2as6JGmBUaYIZu+GmWhY1eHRKpc/c2qyKRvrpEBTo1VMAr9MuFbL0yvifby
cK678dOK5hnGEpV9NpM5FHOommtJYghh9mO0SGGGyA5R1in2+Qon/XsYwkrNImX9cWQUcO3WVF1U
XA940ctXR+Si4eSQZk1iwqypVnxutmyTpsz7TwwERj8cMj6UmLxIHdA+Ui3P0xP5/hOyXIDKPftX
FnuWzOByQEUUBuIiSGM6sM6Qk+ygnqLAvqFPT0BUihD3vP9s8zRJov7jwNh66BNr5p70I85EKDta
ji9mnbj16txH8dT7ZXuUmUWWYRyNpw9g+jq5nc7WBatcPUX0hOy//2OkMv0ffyGlKyyXCpLV25qg
/7lZ7U1Fzf4v0g9dMKuSAbjVOijE/SzCjvxDqIzMdBAIbu0zCZEsb5ir2notk16/S+nvZiBWYVd6
q8t6dpEmscJzRpzjKFjGfMP55+jjO26KdMYxBwzJBqCY8imfR6D76MCWSO4nkK//LVXtOqoFzqIt
HKGd4vX79J7iuOPMS5R8AtAtGlBo6Q8ASvrO8dluFWQKRp/CHcoW4u8YXfz8EYc29lsmgn+jtZFB
/4Q7vA5YDk+8DFFAgyJV+Fgr16YT6c5ex07OuLDVWCfIDaiz8E/frpeBUiwYC+p90vgKUstYPECQ
9v+u0WkNj3z8Xl0tH6Z2wH5LlCSmjdLOdsVKhpGO2QxOkf0y7j7DkRFiu5R2SHGH62xMnZyljRKe
WVqzP7Lv8l1TeH6vaYTGL4L5tihu6Z9LB4QQgyP1jrAgvo15BMNrD+HjQVlDQebGqDqM6n/FrF3b
k5Wwpfz+OxYyLU8Z5sYh2hT+Lv1h36WmjXwNgzNSrEnTHpuTIGwLumMnlXgycKgKZtNjCa0uGfHo
5cWsJWd0cYqRsuG9xCJDad+HRfmspusBaHi/ZcMKOstZSnFsC0186m3kCwrely8+QBMFe9tGVoh/
cCjtltjHmp1K0lNw3rJW70vB4d4ahTh3VkcqzzPzDAIchBR2EZQ5B6sq6EPvFe2ZWfsnLtoE8nDy
LXFk2NF+o2GY06Pvdq2V7B94iVQ4OikRamlp3CI8JRQ6yMIsbsJXpWh7QiSpNNB+KKLHu4io0ZkX
3cinHAOD4Qnr2+HTL3NbpGWFktEYY0uQ87YMudjBS4LdJGfimHnTAYhSbx0WYXrojyISx06bwfDl
JEY7cRv5vRQcTQeDBZ5OxXWyVGjJD0jvqA+AeIQe+QwBXiUYEIYwLgAQfCHNydaBd3mV/4P2q3KX
VK2FKPz73sXpjuWPiQFShV/o2MNBhxJW0WQmMDQ3ZvXqbMRsXO0uCkGyfMhH3qiU6AcGdAdFmo0o
nEzpM7pei5Nwv9ERHVHEnhG4KjN1kGowpXyY3oe9QohvjalHBvQIckovPp60zAyzz+gzAezHn/ex
0bcRwimc81ADrXovXTnt9lDptc7zAn5kZlsdqF0qBv1Bvg2ZuOf5Fs/SYrYC0WuAy6goBBuNVaeu
+bcJebOe/itQ6QBnsf85SzlRxRnNoenMmI/xsa/NFVIZiweLgzkgJ8aEyH4swaCSEISCCMuzc33H
A/91m4+i2ogwG8dexX/aUtCuRYWGiJ/BPtbJdu7DsQY/8oSApWmoxtK7P/qazxXGeKRu2sTbcV8K
FMPZTIMoPPaAoY6mJmayOC+1lGn40l/sWii4TnjqKd9SnxvPz4sw8AwYNL1eP8gXF83Tbf0GxOHQ
OI60FPZU4KBGRLftCPgH5rYoW0sSlp80yfZLaw0WP5c6XSwEtFPEpgYTdkLhX/zPyAR+MPwMmx8X
Ij6fqy38zgHgMy1mF1RFRfEizxhSntO+9Qdzv4HCYZ07kwXwRpQg56bZKO4+7Ma73+hPdMwlm2B8
0CYLnoqLMk2QZ4eLgtvyEblBBuC3E/GRNseWedMI/q63VBozLv87Ngrt96vN6cixhRYngp2gfEC0
e/whsSFqxBWLFVM5s+nBeHDPa3ccjQY4gzvQpuK6UQj76Tty2UzDhbbbw406c7sM865zBtRq67s2
5iIRTBodchfYisgpJNdHnpFSdcOcLGWD/7qbNKDyqTLusD57w0ze011ZHodNYycTfq+er4UtpfPV
6hp1erRiYTw/ifU4z1KKYFrSNOv83XBDt3rLbZrebwZ3Y6OMRNENhCktv8ZyoXVavzI8zIKuTYPq
2hpGdjjKceiiHl6ZLQ+inexhCr/hbOfIJcVHhNxuj0oZOWisjV2vVFqdTYClXLNy/Z5RRPxikC0F
8bxq8Gx6hrwfM/5IPh6SV7nsCIG3jQltrLsvop7DS1/jKxLG5BOXWIM3vIrcE0sAvx56Qmh0Vj8p
ep+3veFdLSCWr8rV4DoRMxQQKuqj7mEjJPu3pDw+NRPtS9Whp6FvUy0Jq/EW6lCfxemrNytJWIJm
7U0S4a0XBs4Od/KSqh5P9dZcODksmhLJFR7WLTK7N00bpQPcNrUJVFse4Mdm8b+90Bx6LQ0t2Q+u
TqCuCYANGytI4YIpQaQXp9kq2LL7kLC0bwl6ZAnIdJpMmxhHpw/duDXofY36nGuO9pRy3r0mKOEj
LHIHqZ3W15gDTwyJxDa3k/D7NvkdQehuP38w6nediBCUHjcwd7ZyGJd6Iel09iMqcQyevHJDYJy8
Q5Q+/A08xh0UAE0dDzBvmJC9zZSpAJ4Xhy92GCbDnR9Nvwkrhgl09ZpfhE4EsZlfmC+x0yhIcMuE
nxslmil2sf6YFLNFOANmOTCTjH35htmS/BmgeE866WN+krXfFU7Rwg5xcOoQeQlu1CYak2UUFmXT
hwRd5QXVbst0eK/pd4J/oYL6tFOznZgIKVvxsprqSqES0zR+ZRnrIAbYJ/+u5ft7FBpkGjSId8aI
aCQSvimv8L4RZT3fz0nLe8WmOEdNNegjtNqNgATWhFysEQ8s0h9T4I0zT4NKJHo6daVCCDDCEnYK
dev0goBFHXF0pjoYfSnXiVyaHhQXVRZfteSMXU6915012mig5Hnc0zQql0x1xvjutBJlRz4It5VY
9D68hruOZwvTwnjROP5ZgGqXRuNQ5bumOwIGNBV/zjuwoZnXVYq9YF3JhRkdUk6t8BTlu7ZEJe0N
CPlNxFcWhorKmITjMrfK1pAFq7IZYgnLYjnW/EX2l5GIGlMwivwMn36ySAWzW2WuErru5laAX1tj
8ntY+PCcznRzbXmutSyk1kcONUG9eeBAgjYiVHWaQKvKTzBFq5AhjEEjehgbFtQJ4AcBvP89uTCx
gEBDrmW7DMoagAfBAt9g8aDPOIT8eTlTEsxcRIy8SzWmVIVwMggtIizaG3Po/NmC2YrE69ul+f4j
qzPwwkFeu3mC7GIecMmioyrxujflw/XYF0g7IPVSWKk1XpR7J60vcaom5wnl3bLuKJD6iFN7pTpW
K36B1P8sEJa4cUcyDJ4YQSAt2rnlAJWJ/7yayy+s8ECptWefRmbUT2L3cKsmXvZpCNYHoQ/LhJJy
uMiX1JcTs5ZRgvVwu8GklMBaWhnUsMnuB5b83Y2bpng9tB/4RrIm9ymAXlVx8AyPead/n28wuxWX
6XvlN9DcOkSCh42XNKQHBUp7cZEK2T1yhnjge7b7eASf0HCrawnUtCzmUr4Sc5x8/mTQeVdlhoVk
klG1BTd4GuKV8T0LyYw/yN4aCAIbY72mS/T5ZiuZkChyTe50sbj3KrClAf9IBpQkRCzBqhpbPYrd
JUJvdtkKYMUCVWYTtuWrSVhSZJXGWFVx7GqSjXNEQie1lD20eJYbIFYRQ9kD8I2E7sKhW8GaclbJ
TKWsi5g/ejL4fwiRxT204+WLpVAJSpenn6sHSrYUj0M3vt0buKjD9lIB1/z1NGZv1bUu6uQNWE9Y
g9IFRhVwL8atz1X0mlCd0V8jZM5Y0Q5lwLzbfmBhC3R3qfeaFa+3AGBNwf7uEVdrwOua6a1kYnod
30BRY/KPvZ0xyQJdlHBRH1dvL590K9QnX8V/5fcx/QcEF3dE4MQYraPQln+STSzEqtx2sp66ZDKA
v9ikioG5ZWcUg2wf9efF2zzPTeyxt5V+Nup0VvllkHF2pudrRtSVArlP433n1FFEDfu3Qr1Rnx8X
FNal1tZqRqaloX+u7oPSKg7I0pQTzXbW1P26XFu2eNtkZitLZnVtffVMaIFvnx0YnKSf4YIDxCFl
4SMIxMktoc9A5dk/AfBVQ5L8K/Frt06zEANeFPGgBlugDj+mUZyO6mhJ3/j7HWcNvCEncQ4OyPKp
jW2afkROMvFnude5q49yi72NVWXJQ4bhXbngvv94fnyeMMqIjMR41KnvqJaW+gz3JInGcryFyDa1
9JeIzokSQw596QaHiEA25qkKgSXQ11X1xL/04dQ8raK5rQ2kQt21ZQGcxTEAOu58/jHMVOvB7STJ
tBlanEThdRKFCdxtFwgJq6kkqwQnl6tR26LkmTYflNlkmljz9e2RrFyVCUkX4oLGosUWUwdG7MJ+
HAEft/k1DAbfo66Z881Y637IloXJWZhgSXf6PUIxGdHT35FzbvKrwOwWeptQbQHDAoO9qQcgJdg1
kg3Tto86SdmKLDnn6Rbxw9I5yNw/KW3nb2dbMPSDT1qURHwdd7Sa/z+xbxvURHLhYMxjTlVeZ2Rg
6PLYs6SQ3+3NTPu065jslNVGQD8C/ZlDLk7D9MelAz7cOz4QE4edXGstSesvpYsUk8kYJHEBHRKz
aiCDZFN5NVqgraa2kSTneH8lTj6nL4RGLsF6mitlBMYByzz3apizK7K1SiJL30KkLMI38w6K0wtu
nnujt9C+9ZgqeeO6aKWAw6UI47BMlcxonoO7KWEGP/jO494SCl7y/Jdy7jwRnpp1kb4G6PTocaNS
JJ/J6NOEOIxHcKvF0UUS5Ui4WKIReLIDYN3iiXIEygpRcfuGwikI5s40BeK2KQJODADn+liwcRtC
Fn16VPCRj+5wT/PG5OJSByDDo2Subgs8OGGEeAXS+sUDiFHQRRSwZN4L0cTBVqZR9ElIUrLGMjrA
xWlaAmdlbCfbOdX96FvVs77VVxqUaYhNs3/a/Oy/uqcMjTx1FE98TN3PdziopXjX587ON12ykO/y
Wqe5HFcfL98HKMsH0owAvupNDbs8GLJbRjSo1B118wDGGOvkKCdQ832/YjWANP/Tir9sAKXFdsAW
CG6sf3j6b7klZp+e285itGnHqzlAF+RjLIb09ClSI3j7RgAnQYxLYwRhTRY8C9FoQfvZc5YCu4Sy
7hoKF79eUOZFOUkObFfWrTD1PUZuvElvi4zBEQplDlUrSHpkxWD74tDeNboTdZ362Lb4QpG7O1v0
g3kHLZ1/YGFCF8J2l6VNsyp9pTdROaJL614e8Zlp5WYkOOgFWNj87gNa2tkeOmNqd+xMl8BZyaIF
AVQsFbw8lZe9+sQIPP13HvUukRkf/hOG/p573A4LHUbfj8bJnynOIaObZ0tMEOHvIfv1/QsZ7A3Y
JBSnUHMGA/F3lQT9uIAs+4iHWbGC0dMpZhVbQpQMAH+l1w0EnvXAIewIhU0FRnkw+atgx41Tg35a
20mzP7KlvsUWfqHppab7ZEJJcRrd35yV12nYK0nJYQ4ptgqivUHg1ZVLhnGQudJMPsUt9hJISR6k
VijBeGBpYQGO4Ka/ctSu9ILMw1WTPNHFEyndqCQ0r0ejRhKxudYFcfa6g2JV1k84XNaWyK0VIkNW
DDqTIir6F3HIpYsTRfDIYs2blCaKiDqGrNSnaEEtLgWvyPsPS50U6WNBQf7MD11795oCreh+qdMc
wHEzDb2b40ozNMz05QoSIb7Sm4ZcswxT+IBp9/1mf/vfYDzLL37A7ZRQ4Q3bYIqQaMk12y3/sBtn
+6OXF/677OnPu8iNUN5uu/RnR+0VOFXEaayBzzOhwygRw0INPh4zbP6Td3YtR6XbzoTEUoQdXFiW
aVnnIKLigVXHr00fwUpIYsqG2FOf1YiMjZGRTMB3ZdVPWSMZclqOoZtJN6C+Ow6+1KUcGdB3LIEB
aTk7aG3Kqu1Sx65sC2XXAcztoQzDVMo1gGcpRMQ2Go3xroOVBBiUDiOT5T9+So2a+00BdmwcZhsn
kVbo6wDzwgUXkosM8hBTEXGo3iKwhISfH7YcNSfabTUPrReESJN+6Ok7/qGhwG/HTZi9S8LNHRPM
64vOxa49isJ9S8AVExMcu1wUhZDjrPQmHlw8yf9eVPab2DJnegzVE8Uynpo6dupmaQN5j4J/6tFW
tu5GrQVpc1YfkCowA7yLmqPXBSm+2LWlZKgopX9lyWY/eXciM2EPlCxyA60SdE5ONopBqVBMwxDo
JuIKdX+zrYHbD0QruOONECm4etgOBIjbDjNSuiRjVGvRJknoQSCd/NtLVhU5c7BszOzrvKnePkUN
h2EhwythJA8x2Mas31Pc7xVa1nhUbFDuIJ8Iib4y98u4iaUk7S7XiQhVcmjjQuuPa6UzfkIAj5HH
pwS53gZjTCJPxCFQ23thZnP++81Gt6kopVccL8TOz3EMc/4mU6MZCVCu8OOnMwXbY/DfEF26oYcl
dX2WPRV2kpsgEZbOq09310nIn6w6wiIKRWnS46tt6IqUDtnrgHv8RMBhfpa0gidoaJucfHUdeerD
iSa6PMAx9z/ZHieNOW9Nft5hbnJ6D+8cgo0OISmbSXRUT7cQi7Lwx536hx2SZOlYcGYTfHYK3qpf
vqcVDlc5Jecf7+RfAUpUTkUzv3G/ndoJz90nTUQGVzlbFH+Vv+BxzWebwH2oiDvawX4iXOdT6/5M
EdOzEHOe5E8JC0zjIu4b3SCHPsbA8seP35qECLD9CnXpzARKfUuv6QredxRbLZoZkEwuKOR9ivoV
WOvVgmAdlHdklip5CtPPIJmKrrtcb8ttndQBR924e5PddKhHXbKDFhYV2P86+T6ggJoyBIrDonoH
qzDxU3TU6TxIvjZSqbTvNL/eJZgD5eaaTM4wkOt8iYhmtwYv9vgzAfLo9BqS5KcrlCxm0DbYaG6c
YSaTvUX+o3Ik9fr0oJzt/sbFBX8fTrjE+WdxtBfdwLjLobq2UnDJ3JV8q2S7Vul/nGwe1NGQb/ED
1+QyImCZwGwq8UVFuIJ+v+n9FoeNiBYEd7xarPhShuUlN+wQbXTePDvgrlNyV9ZOlcfC+5YVv5nN
JPj9/EmYFe1dFfG0435HDFfuq9NeDqoF20PdFETwWPB8V2jsTS6Y9+mP7qjjGonQ4PxZw8/Ah5f5
XDVx6rrXbkz7l/5WMCm6x+/yyC0A72geL/Ob0rjjlBW6YFjdA6/lZOF+GnX64zymRtdHGDRZPtQS
XMyjfiQdjEih3tJSJwPxeUulEqwR1MhNwATXEnP/WU53GwhAohL5Av/N64ghQPPCxTF8MQErHPar
JnNegisAlKP/WOw9QVOR/pAg+W4GThlNYvhqpAh6rDaJmIPYcuPuM3rci/N1sGSkBnxnWKfcHY5A
YaiJ7I2knMKLedMVH65WLzRDQ65cI/3fJfZ8HhtwEQS7OuUQEVIwZfqY7GvZ6u4AdY1O85P2IqWd
ijg1Cmv5G1Vra8vQbyBNrSoj65LeU55pF18VKFS7WGTkRV00tzHAlV8SQzU01Mn+tugVYCyu8cqU
7Mj/RM2PTbLdcxIri8StCfPf9onScLOSxRYzLuSXNA2eoX3B/P3Yx8VhoTxNPY3Vcte/ROdTJ/Ek
eNidUtrfnXX8EBtbMB+ZjQxmEFm7UKbL4eMtJLH9OFBDw973E2Am8lg+ZUDOa3Ft8UR20/kfnKrA
2/jG5igUJT3yOeqsIYJb89Myfy0vHiq1iORuew5V6FbqQ1l0ApjLOenmsoSYcyLyF72Fxb3qN5WA
j2dqmUk18Ris4ZlWhJE5yXtEN/jAYlekdXQes/DFuPb1rcRd/N8aapVaPUqB9CLF6Noz5RbcwYIK
liKDdpwSSUt0zySPopBAWyYKNW+NSOv9TB26YsKOYaj2zkPkuElUG3eBoQLWUTtF3r+T6m/lkKHl
wFGgecMECG3sZOYW6eifNovVb/uxyaRPHishN/zAZOOE6Xerk6B+WcwHXWeCmO0G2+B7vx6nP44a
uVx+sUx5ZpFBzksiK+NYNYMhsPdyqWqESRZ1XOqTu8691jvYQgkc8KbnJKgijXV56DRqXbsfuOas
/OxtK7cPX0b8AOdxcvXLh1Ug9en3UG41OoDsxG5djEBZYEXyZLeUJgplM3NihwHVBYNUI3vQIooR
/hZqLOY/HYmK65uHPxVeeOrisd8SdfCs4fCTKz1dCmz0ETg3KABQgZkUZDi+DFdw+q3lUSwEAxvB
xR2gD9tZclRF/tjEaW9cIJu8FU5KV7URQP6pA19Pr8U/atsZQXSH4ClxadsPT1LF70uXb7Y4SD3E
dzNOGFB2hxoGDWqM+D7okHzO14p/laM3zqbruUkIrJ8oMr+WIZQimSLufp1n+p4ONaeT7nhIYDdp
D94GavktnHYZbdWgDOntSx96oIsMEAFGDi1Pjq0ehSPuSiCe5pld+J0SaQ9vt+JmghKtvsVxIHys
Nk4jMK9L1G3kHVUCao7ISvpAYlJbICsrQf1H4kK1UFLkTpuH78bYQgnb6XABpirtoXL+qmuPOjqj
1eWq4J3zRkOTt9KIRjFy3W/a/zTAYORUtgY9W2cyjbBsj8DDZOvMTtNnJ5F7Yc7ATsOLy6a8jedq
KqWsKrHy+2eGRLC2vOZ+Oov9UXfZJPuw5kFQ2aT+Y8aM1Oewd+1fvY4b8rG5OhQyaG3f0KIr/5tj
XsCw5qfsygaW2aUulx/ex6EZzGXN+o68TAx7xHNBCGZpj//ROFEQJvctEkaORVZb8FxcH0P9gGVM
Szhn62NoPrldD4R50f/KRhhmWH2/0Y1guFUCX2tSb7ROiUjfJBKcnteqX1iHfgkWAwVbSly79i8t
w8do9ytfFrZltqNOWWLyO8BDt3s1zc1HfSeSQ0huaYxycrN2P8oCYY7jxrzrf7hYDqCJUCr41MKE
UMuZUyFz+jTTJS6yuLO4wwdv8zKvYE9lVTZximTPO1S4NB3K16KvhQaX3HdDoOow4/CD2dqN1290
N/ZhoTOzzLKoiYBeBiSDZoePP/73WSrbSjpyL5X5uDo0ZUaI7jVbzKMKMY8IFFwVBCWLzSSS/Mp1
jULgl5z+PoV6IBguk8J7U0lO+rDRgrfJR6wQ2aDImbNWXttb0R4qYZ0P4gzhLyqO1w6Vy284ay09
qs38sZR7t5vsg3TWlHh+GzcO/p5pu+v1ElFJaUTNIAyCpLX2JR4V6bc9a0KgMp119gzhMkEvfjbF
EsNCa9wXyhb8TN3maU9/ThuumsOiWqxOnZYNRMprfy29ytGiLD2ZDsRvJqOgHAv4+D95UstUEV+e
tiJOJ6XcAZnRX7U1OtzbR8rwDS8MjKv6xSJ0ffMP0+EsjeWem4gf7WeNrQA370TcaiAT8kafcTXz
liU4D02tnJIoKguGYVV7JMP+JTyF2v0eJOEgtcjqi9s6k8OodZ4CpHh/U6y3dMsiz9B8lTT7I+Vf
160lHGXBjPBUtyqLqNzLPg4KSIIXHBo/1aPCiMMY5GRoT8cEa4mHohn6Agx9DoowW8keZd093OqR
cbwXW12YI4rfmgFo/ecQ5ixs/vEY44INgvZ42sBHTUaJOrq1pdrKahXIejKnqhc4tGBDogJFKMsp
V1YJhWeom1cKmoiUDhCWpV2bNwNS5Wqy6wP1JXrmxsHFVXyS0ewUIqBmDV49EJWskVgcugyDRX1G
AM3oYfbZ5AHl3ZOxZIG9LouH/YdJy8NjE8DHjaODyZ9M5sT+UcQOsqu4JJ2HDi5gS+cP1GAw7f0Y
DM9gYPFBGMZkGvvmnqrfkWbkg4EhamgcLa+6Fc69jkG+vMBxIBJ1+FXCHnDjstb1qC0uwz9kSw7N
X1DD4RknPW0+z1MMEX29HsYOZObnO12OfuF4Z37tny9VVyfMymGPrXIRj5OuDwULBiKSXmISQ258
S9ZOZCxNtY5shBpGEYDW+qYsJcN7EBztnoUJ/HAjujXPdSfnSsdimqgg3YhO+6EyE0CYe9aioVUf
Et4xmtGFJ1kNYFRr0VWZ+vLplMB8rIb3O5aDlW/K7mIdaVhNm0tW+Llcd6vEQMzlcx/mzecHvi32
QxAu4MLoLB7jSYswqvurNhhcGanS3jJWSr7Ctlscv4E8NN/T/oS3lWqjNRLzDpKVZybGtPCUYfbQ
W7iwR7Aq9OM28z60YodIvuXq8GXxqKzvPBNN6k8WkKD54KUVHQWcQeMfYgwh2nzxJPK2tlHx/Jxl
CMq9VhkPMFlgUpsy1DL7o+UWKTXg9KjkC4qzP/I3iZrOgKgKjwqmd6whNuPc1JTmYmVz1ELcp1aR
HfEZ+PA8M+z1Rv2C8qMKvdeqD/9OHgae1O0CzR/pPwA2bAhhwuHOBQesdynTEimagOUcvYXV0Bq8
B4kH0iVb//Wjc8mR3vNntVKOQPGpcjGorlpk394CTG34xYwrvqmQkXjWdUdjCVn25UyCYn2v79XF
FLDE0Weag4S4DDNRxOX/E6KWD9s7NTiVmhvmxZs1pYAv8i6zX5iqCelb4BE1eHNnsLBf37fpH5iG
UyHEpV9d4sXiAl5iMk5ZQAk4ixQnPe2qUvHyRXmWJlj4cqjQ9z0hsnfL96lF2N6QEXEYAzXbkD2i
ZJ85BgucHRSqfy3AsCvTz9oNEEZJI9PGdrwSyJhEAPL+47HBxypPsXXMxnX169Yl6HbXQWZSR4GT
DZSJksfs1ytoo4AYwzilGKuZEt9cdX5nkJs1/OUn9yUjZWmequeGDmAloow+i8UB8LZnxnXUjAWr
XbPWush4oaKPfDYlZIxvTSY8MVhGAgFVuW6G1zl/kE0P3Gw8Ic633xnOU3lAzEPorWginMCglmPA
kUsN9XKz6JbU4x4WvDcLBrBV6f+w80TZArkS+rXDGNdtvdHzTl1XW8/1Q47+2YoGD8vUQk7jrcYa
7bCdBvpQtlwu+iXoX4/HBaoP89Rifmjp1iSzjoxB4KBJyn3hqfr58/S/jZ4Rs17egbuSQlcofRRp
1lGxW+++GNOdfRJ3qX+hdCWFO+Rw5SdtC47hXf3OeCIc30lrsqBBjQkrLAGxc7OAouSmAsIr5Ths
elLmLrorpWo6ayNvgq/m/5+yAbAOFbJRfsvcgcRb4VSA/p4UOQ1fUgkvC7FtLf/YRXpPfyiWejhI
s2kFHOnuQFazZ8QYkz/FDJi6KQxJb2piHNG2k220WpVhdjIdUm5LHBDleJy3tOji68nTwzUyLARy
rLIbeTsKA4F9//uv5XDxZLePLzZZHbIOHZIeTMS9y4QB3xRR1Kjnvqf5HAcy6AbLp+AEpImIHmR8
GeZ0HKDYa5zPhfiaxLWtPQmHpCVztKAKWev9HUCxAE2XRKAqUR6sOeOjdaG+oy5Wzx5wOC+YCi/u
YrPj8X3zrquCgmYlw2vbiccjRbL9H3jBAULSzzJ+jrnm7eO2G7mnUzqkDjBiknvRZAOBkuQ2A0Yk
9y9BIZbJ7gXeq1rCumKzv/40CtLlQekdUdMZ+hlAu7qG4leQQwBP3phQ2khu/fSQ5534xsoLgiJf
UgQjFAkIgjaZaYOi+URirB+bwuimOaoaZjuA/t1X9Cp8S1W0inHDFWBYuy1sojs+oamOFrlwhJa/
UojTuMGFnRzFsWYvdSWVezyuNsgn6L0sjWQiPYLOECC0MwTRFCvNKYcIs0IoP2me4YHlZp5KvJhX
eaXUjaE9Ypy6cyNjHkPjeW256xEVb59h4xy1FJDUhRklivVLzuPI/YxC63HumFQMz6GJbq8CfNA8
NmhzozCa4kNYJtmsB4iPu5uiu75CvIXNvBhZQORQ2JWSDcd8F3mUIutslpQaTk3yXsm/x+t/a2Aq
UfYTbW7dMEVszSjbVHpFfbGE8jqyeeIiRAPs95HG9EkaUj4lmaVpAwE3/NcrCuOsbhsFMzNPzNB+
tjnE1vYqLh/ztv8TvPo9CNeXWIyZTWQi7sIkgGcob8DH6dCOieJiqY5PhkZ5G0nVBAD1iUXsBfSS
IdBWmVFEFgx2AKP2pzmov0juDYtVJzeydMK/7MSHnJxdNxQ4YUSoIR2RfjoJxdeORIIuLtIzULqz
QrwYpT/YbJpjqYs0pE3FLjjlpznOSfrLoz04GfvHryupm50xRT340bp0onRu3FjH0uoKjgtOUQ6V
RgA7i3PcrGVXC5XYWfgx6Jn2AuJmuHXgT27jiyY/bVSul/imQc7w4e0YuRpPH4mH+foSFTS3P7Qi
2wcL0ybS+ok6zV1W8F9ysRxVwhoGr0Z4OJz5m+AXjdn+VxqQq4sOz4DkubEbk8XemqLtY2kO6zcx
vhJFRKdxR9ZKPHhDsyUzOJOHgVte9G0LL08O4l52d+CNJaLgPPlxd5nB16isOnXvMVQG+nil/Eak
2wuMEBBIrSJHKw1EBLUvb3jG8FQ1h8k6g1e1k+t0kmmlOHV8y6bl94S4hWlags485qS6gePuwzVL
DapmJltvQ+fz2zCB3C80L3oNeQGVue8A3kykAuv+gWEfyvZCBonea9J0Lj9u+ZkWJQRhJNWgb7Fn
dIS4j3sPYy5i6d4AzrCyOktULZypJJBUHCEDdsEPt5Azx8GGaOXl4sqSKH9SD+mjqW+ijVndLAra
ZPa7xHnb9Ln2OwbMsridFEj2XFh0YSSCTm2O3q6JvtKHGLabq907TUcSWny1VxLHBWt3vjfXWwPO
+ga2Uw3TZWbP7J0y0nXjaThvmxjkbDTNnaR8fEZOFAGWRwESHrw3EpxfCnosRbUNipTKptJoHMGc
C2pjv/KZN5q7XqYZk2HA66OuND02jfuzIEwmYPqzQFtGJgjtNqgwal2Nqr1HvnO2WrNInsk+kTLo
BTS6eNcRf5UA0G5Iiope2fSyrNakpTPDcJy/GTqQONhIjXH/3t0gnjhHhAL8oPb4jfmoKKNZ8xdP
9EKJRft1zeLeaggLbCau6kuRO5e6ZbgMfJNI5+7nZHJ4cJqLSyfPQuTrTXwATLrMy/rInV4JBY7Q
HwWg9Ik+0MMSpqNCkRamy3XTTO/6nWjVXv1XfsZh2OIWC0jEI0zHH3nzn1swYT8CE+myde5P/bMK
ZEL/XuTU8kL9VqJjXjvYQ7oX/5XcB92QiSwdekeaPS5QfpEf+fPVlnkLdVQBZVxRUgR8H38KMmRk
lFeGkAjwCj1wo9rncu8Omns+nioWZxCytNETKNd8olhSVTY+X5cBdbUCoEzm89YF2j1kXKwJtSFe
oo3YLS/UHeak5DGWsP0JCiyDbYzIDjFNtrBhlm4CEJe0wvvkjp7o98fLy97gHnqJGCasbDkb5l1D
id+kCtH4aB2D+f6e/coo1ku/aD8T5sWC6SmPY9VgLZHayDFbcv0bnsusBgj56+RLyFaDl1XlxGv0
EsCftVrnINQaK8ZziZK97llHp1aCVk8+pc5WVaclPJLX7cdZSjgRWdtaw1k5KvdGQn1xHiNBWLVq
GqGP8wBYR11XsRNkCKjum6XUdW/M4dvNp//f6oesL8VM+mz1yhUtsVGZlGmPcJfTKEiz+M2MlEnM
qHAuClu2h/Errfa8AoE46Uw71QeqD2PivRNeFXPpultUCIOm5x89danDFGB/8UtuUIU+NbQhouTb
VVvHM6NwDDAwgpSPlwP95ONf+qAMV0+BDCRzCmAPco+JCLOcbWJUFgTG4Zhn+m61aL6LRuMBydxp
rxUqoDJaUa1sKPEviD/oIg7s+rIzRvhfRynh2QGE1oej6iEB8J7GYEN+IztBD3I0mOVHZgdVgmsa
164m2dDdAKOsaGrWgEG3OHqfwlIvmyKEn1UiG8lcjLPgM/nwvjSYzElvfZJkKy9g+VqcnqcJpfZ7
2ZA+p9IFjPN0k6MdYl7jLsF6+9H7fqFy16e1W1HEFtUr5rwpuUkxuL1CBKSGBossAKPPTs5iuMyY
cVev9I+9f9x1b721gdNinZ998g932Q7I6j7AMgA1Qy5Bpcm2KFZQ/tV21Rq9eUVDWAuXh3It/rqx
QcvBySl7ZpYtppMwQil7007cQAqlyf30eE1OSTMvx12ci15cUloOqFPGCOI+5sCZElRPvjX9ZeQl
Flv72nza5BUc2hvC+apr1h6tePNjpyPIdMdnWTzmXFA9rC9GOXzJ/7kBWi5gyH2az0N2TKXI7jDx
qNDLSStjcsd7em3zZLzalXsXEsZhzXxpb/AxDWt8q5hl+qzgMBoIGI5p1rfHFJ3PEoVsd3p8s2Zo
RNP4WC9APus85TWUrhOOCwNoVq9zEfTrOAyOQ+4KKfg7ZTVDwwFHHuMIP9LFISmfvGpmBdTLCA5z
GLJ96EDUfWHtrt6LUEWQedgqxklC/IDVwAMUvZUB1Im2r6ZG190bZOrBVwoJQLVHxxM1RoKU9+Bq
p26wXxQHum/7azQljottS6jKz1ZWo+M+veLOCq0xQHCB+xjBUaDNTOy0CQWolyQr7EeeXdZ640uZ
BMwB2NutP4YBsbGYaith8AmMPDc56AFahAc/H++ewgVvB1/ON1aNY96M/1rTwWyBe75mh/kck6AS
65aoJZ9QKs0g0oMNZU0AZEkgV9ekmh3lRhH82uOa5l6PdwkXhPTgZGhz47XJcpR+G6a/mb7vJM31
QpirNCBXJGip1tONF4WRwdUlh/A7/OMa/n29nn3lj6tdlNk4ZFkwdmzQnT8r93L/jQfRqobNhrTM
mecSCYIyFt/0ebd7m+X7c0ClQx39I6Ob4b4D21rMmK67ZQ9osHHoNG6NGtXv0svmT7PFUR/Fg4C4
In0ytQ7qZ2n9NtmtPjEeRQUkhCZGYmTM72iizBl6px9Q8wN4/aFBUndPPpozJ4wG5/sCnLTjlGvt
PvYlyy1WpYz1Vh7sDIK7e9HISBGF3QUmZ4oienwGmo3JXLROcBK3ktsu3VAL8y5SaeSgePEGgUmn
3FpzKN0pTRSTwx4go5A0n3HrgwYpd57im0ODyUIo/9uTLKYP/A0H5dEakiOCxSrtOaFCXbSStGv0
BCpEOUZUwY8bzdc10BkhqbBE30WZ62WbEOselWp4ZY+10zrt+PuKnNVtQ/0+auDxa/Wv2gKwmGS0
dKPccetpL4ej9uly5oSrKjwI2aH85gcIERRVVWOgTH5IO9nWp378mq2JcJ7FV9ucCINhklp2KkFd
OosxHYRrzNXbfI6qPXBNMUuueP79BYkZwIWmfif++KXdbFyHFMHbtp7KlXdQQqeOI0MSayTPUx0/
eUm06c4SQw9evHunqNUXJ6L+P/RVkiEvTNi0DqE4sJyOvcyhitvNIfn8NwMYKJMGLbSvuK/VR5vw
WREWfHuNeQ1uIV+1bzqZMsublq/CQgFjlx8reidC5X269ZUsfqWLXaBCnNv3ImueJVN7wXhXNc1/
yrzPlBPF2cfgOLcEBZtegERzxHWnkBgty6jCHH7VB5aw4FJYAK6k8d42WntzafaJo/zW6g7QiwcY
ICaWcOom5lLP+EjWXQ4OFTzXt1tVlBGyfXk/gIg2qa8l82RhvYefH/6zMzHnNNiJ6T8mDQbh9kEd
ayCj/ynUrqtsC72SYqkcX0Bb8Ibb5YWtY+I5uUYdhFESlz79gqhcN+iS0tRbV/0mmCoWcgzsVSNm
SYz3vGD1e231m3GyxQAIyIstMyeOb2Gvvp13nVZsd0Ag0tQiwPBEyRMelbOn2Py5Hwynh8WsKgn6
4cIJHiLFEVLIJQNgMwx8zw6/eGshdM81MFZbAL/QaYUJ5v9XJK4iukvbUx+eVGvfYdpUdA2bdXPO
4QsDamZbvwTSU3jqXf3tsm2sTZrtIK3lo/3qApbV+G5q+DtnZysflDVa3d1X44vJU1J35xjO4tmb
ZYjoBrtjyL1xKzW6bgjBe7cHwigMm2If+I9RyrZRzrHUaepBMujAvE+EPOvlKP91F7ZsFvNMluYe
munVcwa+w2QvdIH2vtlQ8RyYUZ3ILXAwd7MlPhdqd2idp4AVPXttTreXtNaWADmUDzWXrK7EhDx3
Pf+bvqKyocQlRm/A66mCt9kG+SMHArjuYT+piXVi0z1joG63UItKgG06T3kOi2OTjsqvWmdn+9yw
/FgF4DUq91qhTiCHAPvWlgCDt79KxrwmlSVLzPuwOIMvripHLSYNcXH1IzwfP0vveWmwiFm7H1+W
a0MYcgnBnXcQlIJzgiMeITxZb8BtYByFiE80FN+U5P5LkZaamUqp5prdgo7a3TIiCAlBZ4gtNJUU
IgmmzhrGzA3sblxeeIXMD1e7db9jv0BbRrItujSYyKy1v0P3jglvss+Wy9uYz3HKslejUY6rHT04
r/5sMv5nml3CnSoGh8IhwCW4udr6LXDPrLM64xiO2vEkm9kQilp5AXBabnq/1gPnLMtRSDp+j+RG
rBrypWzhipwqO13dcuGzd7/7w7CukEPQc04XiaFDDnnJfk7teib95oovjqI9HGv3qES0IL5IOsKr
7zqzNFeFL0ER8rvls6X57qS9W+UnJk/5YweCHMmDQwZZGJ30YpRpf8wVX17K2B3Z29AKt7a2gN+y
4sK+lHbMBAZ7gInLoYlE0R0VGQIr+Q7zO3pumjD1EdM7u7ldTYuvDHpsZXkklmfwuXLv93yy3xNz
ZY9s70HCZz4OyZEBhEwQZaApLSQ2V4Adm3hEdP8F6GA+UlCXITwiS/NOaUwSgAK6x8h6Wgm24s2a
nnisckzDnkeMv3oSMtZQUGlu8QVISMui/lXhLgxM5caQFIaYILwdrgj0ZPHVsvSY7Fkt5OfkvbJ0
WPAdPF6uemvDFQbVUR/Ls95x//ouKaG+47TqfvzOxhLt82T3E7YtCMOO2d06B6kTyIP+uSx9bAjE
daXgV2thY0eWuFwHguzt96boB4xofrenTb3Jaa5kAIKODxFNNGffDoJN0EhShwJqQg6qVvfJxt7E
hCuV9WlX+QQGo4KjTaZUEXBtF/Rvyy4QH5KPCYk3ZX3aZ28HYI9HgVBMJ04yp/kSe2KL5F1jkHXe
GJJrRhE9qU0Ijp55BLwE/fEDj2XlrDNxyJ0nwkF8/SsOPHqVn0QrCNwUqAITbWh9ZcQYXzEb3y0B
cshrWd9ukahVWQwqN+vbHHg9oMZ6rMUMTGiu28as1Nq7YDQPL6vXHHLJDV3adLDSgBwRtSnRrB1+
VN/2ZjfTptq8dpeA6Pe0FQWuytn0FJZkisF0j0qdnaOvHO2t0LXUMod5GMOwkG8PO7OOhCGhp/dY
w4KNeCq0PhPmYE2GZRsPdR4l2Y0C4KDSil0NXskNqH6iUay+mEJIhIfmCKh5su6COvCafq7TNFlk
cZZczeAPRZoVEqwWJ8LAG7QYpVZDOFHuorWE9AAKwmcXQeZXvk5wyK0avMCSiYeI2i3w7COFU595
8G2gf1Yqul0ZfVdth1TFW9bVkKUEs/exFese2VUr/BtCsCw04QmhKJD2IX4TvsvkkBC3oZeaqXCg
/b208cwBgn5KC5IiCo0Bp+eysm8pjn5Qw6/lqMVwyNKDqdCcclDAvUnirfTfefJ2IZn4y7IHnCCX
QktvXs9e6X+Dbs3PH3+1Lztoa4B2zQFj8y6DYNBcWyXRJWE7RlyV/RB/gpXLdT4uCax3CE5EaeVp
di46dlSBqI40t81UYy+guffAZ/5Xcp7zGMA2ocTGbznBSEEe92wd5wS9oBJOTAqwTWCVtYShfjBG
DDpqTK4WORfXBpL9iLlOSCbEXrXDIJlre2/QxKp7kAp3gP3k/GJRAzL6SYyvCET4IEYt/bYMI2jh
7MEE5bhrNGCUBYxtS6y0ouaD7AS6BGvC8lXNFGCmpkNJ1n+59uGrxBeMuLi8JEKcAjfXT4iSQm3H
QvOnksWopOeZIDTbmO/JmI4s3ARYlZzbsvhCVPwDNh795AUhDqC2VWkqfcfx/Fo88ZiYt0rabP8k
C1MVmpcI6gpl83O9BD/BldW9FUjlXMvwCEXOsmbs2BxPwNGXgrsvo4GRKAbMqQFjXH6YrikpFFSr
lH3tFXUWxWtEZUt4BOdzGaLc6N9D9oULjQbrMheUShwqoFHjKWxQIAsXPvTOOUesKkrM9Ol+LK/D
91WLZJRj7BLv2heGu57OLC1PPG39+YJFwZuSMGJKzY/wghRs4O8x0gYWfeon3Z2XXWFv30d8BSy9
yiSsDkdLfvijVBDwjjg0qpyjy1WJA+k8Z51a7KupI8oyimLCVsv6h/yDBkTIHutNRH9SmSbXfvyr
VCzb9PQuzcRf55yuUDMC8aWxx4udr6ZurGS6bbCo+1wSHhcz7sOD70deb1OXqmLfUE4zAoa6K+Pr
n4Sp0h+rMCXlzbK3+wdMn6qeEyDi8viKVk+ekd6S1OROXls4FN2IdK//ZS571V1MU+x6ijWVSZu+
+U62Zo9lutbA9HUrq/rKkFc9S7jwM1qLmuMtjnTapRmBIczo6Nf0J4qrM9PJ776N1iyQQRJ3s7eF
puxNhLf9F3e6kacB8IVOol9wB0Gi3p6EO+VDLgV7Ar3EhWbAqnN7V6i24zqB6plqr6Nn7ZejStuG
oz65X+Nn85N51ktIRBYGFk4qfFkop3MOuFCWKFQ6xqKFe9qXcotnHLJmpbVAPHRE9yfCf+Ryb46p
pNrQhsCrXuKUmcxOw9CL4BqRSy9zGEasdceyl4AefAKjes9KcBKiTim/kznlEsskXyUqREVu9AoH
Ui46b2rn3mnLphucmyyfyb7glsZql+19BV0HlKg6bQFiZrXYWyg/phEqYo9plB//wvgk3lrAdZRv
VJMCU5zGu+MNdmQsqqahcmgkVnYD+3zi5ym+/Yfu/sqb5VIVgWmkGdr/437rZiafprJ76lYMYCa5
rWnkyxKbBx+D3a60hi3T1G5wSsLbxzuRjbQeAqOAbQLHKGXynl6YBImKNNP0InT+ozJPt1Hap5x0
Kk0PQqpSsOiCBDHI59EeXWlVbsYaPbsTwimPQHkhbJgMGLHaqoOdXSrQfNTZ/sPa3dIZOrjKSezo
X6K7edftKnCyNiwcZE/dn8I/tTPEQrbsccqKy4AajtLH/nx6HiL91sBZhFOcEkMK5i1vIMX0znND
KMn1s8vg4lerdaBlsWYcjRsfevB4vBqr6tYS9Ky6W1q5MWh9ZaLe7BWUBP7pr+5Xw8/mGDsBCBBT
WmAJOmKkgOQG/HbK1vts6PrXBOt0kU+NXQpUcnnQJKTLnk6/zVbC6G4UAN/8fZAxbOjypy2s2x5n
Q/VdlbSZoU5Hjc82KBmwXAscMDhsysflwcDKD3ZEquk2hu1j7uDYFhprOt/nssSQg8/9XmDk9E1m
G6mG24WDMq8g8xmj4+FCRrTX3guw1XRnAM4UGeZi6YErrGW925sj7jva8ld5O9CqxavUK9tvwuV6
PtL0C2MJol/FpMeeTFyrB0hNQ0haXFCMKHSIAcKoBK3h0FXFSNxWwTK1/qGyJUSUfVbMTwVWXT3c
/Bfg2rkKI+9kjc/yO4s6FaLmEQ5lBjXIDetSr1nc1OsqDVB9gtyRhvZbdfNb4RDjnmTSsl9d9sjL
aML4V6BKaaYEqvUchpOjgzhMava7bJ+MuI4hbRXSLoTKpIcKCKJg+Bhou769CDUWO6SCycPti3n6
PI3aQ9e9SdLEZU4vJyifdmGbI6bRA9Q5I26kFeOjGSa5txMikTps67Bt1F5CiPGXB7pQH9fHR0+O
h/dkQcOvAd3HMebNMyzZBKTNHhUFv93/JNCzLORWGrtaZ6pM13/3pNPOFsMBtb86DYO+HkiLNd4m
x9Q7ffr/Lq1CAm4ICrdx6N5cPHZ7E+rQJXWW9hWf2/MMB+h8sOdLg8xHh+Xv+iAJ4syAZsASWCnq
bUCeZZBQ+eIgT6zC0IMQTRZKV2WHIxDZGHzG8N4tOb+kHK5B6LHYXSwGLnK5F3Wu5WRQq4y9vwCt
2MqAv+UcR0ZctZYTexFzFh4nyDiySgqMLestkkX/ucYo4LCMD+kv+9jrR9Z3UppabGymbVGuPcjv
DWVDzPhFoZv0yGrenpqmYYcYA6hA2S2cP6C3BjsT2Ne3YOaiGJWCiqfzwT5B0jaVx7RVcN80ntY1
b59fYYD81wTrOFgwLAx/ucnorVuBUSmzONXuA0ZMgIVk+xIj5QiT6Kei/BQyEX9x809lOnq3ran0
/kXTU95RkkFiZaNbtt1VNEawk4s4zQvG7re72X099MySHFBriwtEUz7xMOTBoONLitiaQkSamJGp
+I3CU+oGXDCIh+vWCJ6YzmZudk0kg8C7PXdSpIifNZnTatCPy4rEkfzQCQKUKBk/p+uRRi0Zx3nS
5F4AQeEtD8K6SaGPrx9ARs4L/JRmjCdeRBipdWw1esHvhDD0D/dHI9v1RXbR+nUrwjGbxYqgjQYo
OdjCAQkiGezag7wuetjc3GRk3WEQF9tX0J3NONv3QHEHqFgNo9xG3CPSfs4W/qwm0YnxSTZwXt8A
bHJeBrxzVRBEloGyNG44tGnyHSIvncOfvuKJicZjVdyhTwn5PDwiuV6yyTX56I86kxSOtf5+qkhp
eaE1Ner3Qtj6OcimiMKh83VK/FLNFJHnVn7L73cMo+5MZMi/OGwEf+Qj+KtbsFqr6MvQPK/DCc9Q
N55+Yb2rP3HRVykRgVgHIJrq/a+C3U+ktc73ioNJ9ONAHKPnWDArDdlBV5lwdOnOb4OC4FjG7hJq
Juu4Bqz1Y9res5uMKEYUaYzjjifH0ymCuEFmgnhFJkTCZ8Rwx+UOcHiQ6PQVG8Rswzl97utBmPyu
xrrbkWTg1ybCOLcFv09AkExaq4htuEraXcIxdCKkrD9e4278lNZ5omZEvXBrEbAMYn41YOG0B4YY
DYKvFbMJV6N1cALwxL0vBTZAqI6qGoiZrVhf836lqwJBbUDYyDlcdhHZ37WUhKdxGvuvNm5sXRtV
ERRIY5su6snHQk13B1leVvj2oE/l41cUTxOZlCOlZ8kSQwvMdXQ1NWiUMkSVAy/jRanBSeC+Q8Cu
SjcVzuj0pkvSKxkkxKR6j5lhcpD4Hdf3lBbR7QeNuL0rydiKWK5HaK1Ht4dL1S31YyKB9Sh4EjL6
cCTjxYEY7kKVslovFJIpfN+Bxdn67+jEq9e/GaYgvJMAsXlyeQCvhyjRVbwiDKuitKx5H+2OO2Ac
xZO+cZc9cf+DRNJdiwfjwT1btVWTTn4/cimn42aHbDb7hmgmpo0MbQy6BRUaW9TkblmRKEm2HIbz
dmjvQvzCK8kB0JxteMc2goT9kYshdYGyieWYw6i2QfSfyE5eWxJxIoEGq5ZxJTlWHXfUG9gZC66+
ZHLOFt04HCJSgKb3XNztnStXUuvHK+GLn9lZ+zEZ9zTC0A6bZg9TAItM0S8jNS5+1Th81p/gIF2U
I/zYPcktNMW5mYjApk4XVFy24T31CP1hdVq+IeRhajRaClOtDshiFeDxqqHGWK9d4J92lTht23/N
wyLAl2FtrqhoW9Qze2RK9q0gGlhD6JtrIAw88m1KEZvMcBTufD9rxH8GhFe4Fj6gQ6raIPamavCU
h2FwH6U5vopwqrgyw/w5TWwcegIy8XxoCyhQ2+V8uZrypv0v8sKKD718ntkDaWYGh3auiU83NdRc
YRb3bGwPiGfzWfQ22/ggOMCe0DvlzxIhnwpxWvylbTvZKHGa2TLyIay86umf9AQERXzcfAfKjaWh
4TJadvWG4qht/+9LWO4dHI4hWguRnzQ09qessCW/gZeBtPyE6uuA/q1Wt9IVH8U4kSMJCfsdb3hL
wSJy/HqB6pw8Z+K7pICXr8qlEjnAZubVp0daGBMo7/lJ2efnKJHaqLeN8uzDixKUKGtPGBm0dPjc
RinSpKKTxJAX77U7PQM0w9H+l4pO7pcgmcknOvrrBszUuMqU/YNxcJjUovciuvfxk8oxVUaMbkxM
J7AKMpgfdRr4EnqPf7Pz3MD1oTrfs7pzo77UhbfiqhXNYLXM3ihZdQkTdTus8bSt3sivaoDRgeW5
s8VLZ8uos5SyA/vIcbDVCEJOs6YiAhpKP0CH9Bo113AmQDGw0mnvrG7BB40NwlETOOTCaN90BQKR
hn4/HlKG0S3+/YgP4O5qiX+xAhqEP6/otxGt8QjR7I9v7yqDFRhJsO04ymmKXBa+ijIdeRmsMs2x
phYoFJ62PPB+NDd6aTfhik6inpU92eid2GoSTEzBWLTyx7RKEfqfRW6qxNKERJDoZmF5cKWwY+4W
m4RM5K2d2XDfm23uOthf2ne1plRTM/Uztnsp5Q0NbFy1YysToT1ilcS1ilABUU/YAPoKx80FON0p
ImO/lgW/OIAGeNrIi7DQ5PjMxycUuB8niFqBU/LVAfBZS61yW7Bx7rzI8x+vWQLZt32tvh4nr9EY
8IVA7TnwjIzoZ1o7nlDevZUC6Jn9OiK5sAUey8RDq5Q1TQbYM/IZ2K/q7NBN2G0rRzlHuXOkiR2B
whcAhehX4tTuofuCqHGEkENIFs0Xo0OHeOLCn0L6HR0PxKwVptRxp8W3q/MIBRTnxQntUayjS5FJ
0MeuP5ekVXrQAG1bo3M7dySemAVmvgG9syCTHy4Xdq+HPdM+PncqzuGGVdz2wXeq3w5UqZUAuVzq
ZuSAqiQurQWDH4C97GB9/X3oBDUH0+r/oNzQVJQKNpTwJE5iJe5NamlWx4Lkz0/n0B0UAbn3dBLw
RSLJizIW2qqYYhdJRZpUkiLXFHaDDTlxHIYJqsnb7Njq+4q1z8qvRUb2ieilDOpl+fIsRWfI6c1g
ZKq87Fl5DcmmGvpOAdyHczvEYQv5iFHcAuPKxqK907ezg6rJoYUgt+E5dfpB+Zv6JnSdTrNC1PU/
Ydl+TlRJ0Ip8mzgAbAKztdYwzyXnR+L+ugWyhV2P2s3kXTxqLyF7gNgtE6rRGXeP9UPtI3QmcO4f
AHhjUemy8TqVqJ6PzIt+qXiQD97UZ21f6sfMYtdkr0A31o/KOXNudHVne7uBxZqH81FaRwFQFRNZ
WMaRfXUjuncBc6/OaVrLhHglW4LNng0ujg9KM5eHOH1CiOcBBqZaN2x64ypAcBzW0EuS6tRj1kLn
6KTLNLHVeVwTDqA2sUNRBlYOjSG+jret6nT9TFs5mmM+MTFCRsS7+OwNwEKs/NLWKBw9TP67/juE
l5sHxUb6QYkH1OPaUAq8fLM9hZPzRvnrD29LDO8vnSItDuhAS1wk554iaJzBbapRM8KLBl0UaqRz
LrvQLiMwf28ap9k3JxGMiRhCVwBXA2lY5KKLGt9v2WyomvspPAvqBVH95n8kk07PGPoMJBBIrsAR
8WXQAMCpTBILXXYPjNZuTQpTbq48YHU1+knZlNUEKJ/W7QoTCuuGzqABuKuml/LCqA+5ovSUKuCK
0cXNz5ViI3ZUPd7928jT6s0WsQTrVKQR5Z5Uw5OP8Y9bZuGF2807A5CQzJqMqyfFa95q+B4TGdAI
1ixC3M8CKXUNYUv6/htjFB6jla6B/Dyq5PRyGE/L21SpkQlEPSrx/hNdgWqxcPBmYjF4lB8Y7inJ
3FAbwJuAn3J6k8pIdT8sxv2aRa4V9xLa9wAhWRaIbwTwKbqhjk0OCmNHjVCCA79htB4/rjrF50IM
eA+EePzdRUrdhiRrQirT+JMjCZYxzIqD6jUfjgylvlt435RVUMTP0KPc/D8hmcC9ZcDdZ8I8IP/H
90RBiYTBOubJPvpaoS72nOtO4YSSYpG3W6M/PGLDaJJhqgCoOmZhaq5onRlcCaC5o56FQvDZ8YaR
f7rsrIbvcPUAbDEj/rnpP50TR7eY6Kd5OBoNeTJQD8yfuhUbLvNiv3CqmguQPDxZpoYR3Ks5fRs9
Z7dtBuEHM6ZBYZg8YhftMHuqe2vE4/VEJ1qodmvZApYwZE2/40T++oPTzOsCMuVYXU4elveJuPNO
Btm0BIVlvJLRVW9FB/qwO4TPzN8+tZeqYq72E9d74J86Y31aVOYqMXh+dgM5s+VZ94QYtGH/anjB
ULVsLCw97oxLTw+uI51ZTkG2PoR1NMZ2QDCujuZ2S8colsI1BIVVAeYFOOm1p0lHhZ707hipJq3D
gdc11xyEaOPG3Hz8hUBFJix/Jkw9wbtF4fWdZmFiUsmVhVZR6ZkwrH7KNRxLnIT8TmPSa42BW5My
sBAj2ok5v39hh09Nfx9rtAZmJvKX4O5dgpMfz4vQow6uvEQCcSxSzZDPdpdgkOeNQnO9LLHtNruI
GTRIZ/puZRxhaKtTasG4fvArylI9IckPe+SpFKW0E3ZspQpg3deltdJXGzzQ58jvNDVFWbBnTrAO
rxMPkLtghtA3EwaOfKHVVvC78Hbem9FNxp4Nbs7fiy5i3e1kw++Q5lHY7xru3mvESnTP5nzO2fzk
WCNuYzHrtJaU/41Df8cRBpiY/3WBLYl/S2xrrB6x7/xz+v1hA+A6muBiKhI9K/7y6LMuUDh3n7CP
C8MmxeZb3dB814sz2xo2QmPKrKrlbYC7y7nF4qqoCDWucqDUIYBm43dUzF5iBqBUVarpapdVuj9X
9P2IV+M5Nryg0KBvuFA8HF24grSbsaC7p7XHPC8QOWL2c873LeDRIwFoygdSWtj+JJ482aL46HfJ
RvIHTPNRj/IPwv3n1Iwu3kMhqquYdass/pa+W9jMKOBZOU+a1z+CXft0DtM0+ztWIoITeSdbnajA
bVfn+LckQfrMG0Jqh1Frg1UbplOSKgi63hL8LIBFnisIG6T8CYV1Sw7BHvz3jRAeB7x7T013RZkR
ByXjgyJLWhOcsu4Pu1BcZ05hYVuaD0AReq/g3J4pAKGgtTcHrXNnlOxFpUiO3Ge1CuhIThUPap1H
+cPE/I8xQ+Kzew4kzogaM0uApTCD1KI0c48Axtq4Hrk7M+nx5GEDo6t9lC4dDo1/JT4IFXbxNuSJ
yHhm8qSQlB7e4+CdanaOWDEryAWlauA0yPiv/L9nD5s2d0yMrq1qwph3CsoOIP7GcnyXcGDRuO7B
XN1b5Aq16kjdZikvzhhMLeRUAR6e/Md1d29WQxMnJITm+LTrQLxp3q2A7QneB/qzLFYXNQi7LRCk
lAxKYHWtR9KfGBWFV8aDG6eBdh9XGoAuGt5cJA//ddvfiuYiuxg4ysW510lOIgRXXjlscxc3cPRf
nfA0tCRs6vz1Ikc6BnFO/mjeStwXdKkTuqdkX0vKZrT8lESGDZIBpFOV+YgelYufxF1zplCkdlxa
Zcvg6XFRVjrN+8khAwCu2eAaiGgKMD291sybtsg7ZKYMRIcKjYCfETaS+LVDDsmuDeHVdJvkUn7E
9EjDNHTaC8sqpXiLtBEvuRF60uA48DTCNqZzINzKTwuP0NFAoDhSH33FTcUeSEkkvGSJBP3/D4b+
LuauOSP+yOFw/EO6k+GfBEGK3e4wjUkPlziiOHSsKVc4JwKFdLC2bbVA/hXnht0BoQ2qH84wYOqY
nrOFwscg+VM26IoPEEMgqkI8b55PKGxkzGFfjJ+EwXGapzDOI9JNwlqWaoqFAtXXsYkPmsYRzlV1
Og+5Qxj9g7TV/DcADOc3/pQtrYxGdlzoLZD37QeNEabj/QXVrIT0s0gYpPiDxudzg85AMkCTth03
bhSRpJCKV97OHPX9qziDD18sUlLsO7yNwt7OqLxGoCYMPFs6SvbOZtKV0lzgiMuBZNaSoaq05fbF
vmVjTZ6wLB1vMrhElndEKWGZKQZpZ1aOWJRUfEYbhLZU71/YRkJd9TdSXKYmm4jrrnpKMeRasQ7F
RTAIUoTpanJR1GSrN/b2Utx7CesxwmG2y3pGSwaPGYXDukfXzft/vNHjNMYnfG2I40UgHY1y1Vqg
qlR6TQQUZ4QOiWJIOoWLTcVmXNZEER2S2I0YW71IwtQHJ+xwrTMMQXTtXjBI2VfLJtvmblNQ+KoF
mCyW+BJJiXrb1uRTahoRIyL1xYOdnjESmLXEmY+hXXue3/C8og5EEtHj0zdAIaG37PLesSNT51NH
7Db4/rARZAQOUG6MQdEaMjidg4DCxpjuJ3x1zljSEn8dZtgKUWkXnnoBksxEFyzw8YO/RVs8mg6G
Ii6G4UgG+s6jYd4+cB/IvSiK9FoOiMici4urB3ewSIlsi0JX1c243tVpNXEYC6qgSaBT/kqWvxjA
VgaujHOkI0epRq5q6QzoIlX4Gyd1oITiW7iyKHvCyN8Eye8Xn2jMKnpTO0qGLE5wLPS/lDqUmIkp
IfnQSmGrCQKQvxIoQLD0SN26WJyZ9ZfTQJvuKVdnqgqt+pBiYK/4Mx7ZgIujk9FlVNwLT6LY7Aci
7JelWy3oQ5/8EnDNUZkI5+DaEZMk9dKRbT0A93ZT87yHEtnfv1wHB6OURh0FSygQ1w8uaK0ei28N
V/FdD93X8y4/Ugiku0z+/8ymb9ElxKNDwBG0h2CF1JnrfTSFxrVX3w35DO+EE/bOLimuebkN1Y5Q
TDZdiDIAgjTytNwZ5JBmU/5mKIu/roZ4FY7g/V7wAeKb1WhIso87P5pco4XJmGD0fBoppD+CscqO
Zq87fbOgEppa2GnzjcUpLHFD9wwKa2Hz41P4aG40PzgLyzEKzFn8yqRj9yu4YZOiFhCq+ddX9dRi
E0KFDSaR4+1I3sbFGv4Dh6Qb8oS6yG3vqp5HCGgwwdtmaDcmhu9eiKw6k94fuEco0WFGnmGulBAM
YJ5WmvOSJ/ONjTPPKR7RmuT7ZK/b2tNS9gFaECMvUqvL0jYrwhm4pYBOhS1Bgv3V+UmcBXM3bjlf
kF5WEjBLH5mEnYyh2+Lv10YfKm86+2t+DvwiSusQ23/yJ4sohZcyva+jC7dUGO3BS+ICYgxTs7Fc
tpuRsRIo6sYuUukn4FKa3PqG7bnjjtL0X5vxPt4yhF69f3v8+ZLbVVlqTwCq/CVGXgifVqYtIZtT
eMUQidB1cSxBol9F+dHFOowC351JCKpQypzVSYRRHKVhFs4vbnKprAiLaaD2RTVaXtXKK+OnHc7N
Yb6WZtMGLAw2lN3pH1hlzJL29tfpDIkgCt/afnMppLUxftXTMEL/MTtVdWsQ7GcrVPa7d5E3syGY
+QvKicKduK0CkUEpL4PIRMzMRqoWfaCLqOSYvR1qY183SJXaAc3fR/InjT5QsJVngwkr9jyw5HyI
KZSreNpnPbGPFoJipy8AGgxA62zlaS4+XjVKNjW+IzBArBp7G4iQ8k5aZtqtPYOIBAmW4JNRigC8
Mgm6rtNCgLG5+1hLlOB465AXZXpNFISKuPgix41z9ejFIuA5jShvJzK5KV8kXrqT7IUz+8Vx9en7
7Sr/e6JSGL9cecwyJkcTk2+19xrDdFqL7HrU5+dP6hjqEFqQNeAZ9mWqMazfIS8avRg/dn425eYO
gz9P7uXIpnFynJKd0ll7BPFlxO8E0AVf/78XRmKAMreMq3dBW+UnylqDGbS9YI8qlGsbNyMLEgml
QRAqD2qWfq+s+kVvLjjYDSlwJ/o6mD+RbcbH6NjtlWtgknOfggBC/mnlzUYBK2QxBHpELQn+28sk
gFWUAPl6zf5rb2MGp+Hs1xBt1ABfmUd8y5BAhRZ3YzJ1xtGeY6fXgMnNpz1TeWLExw3NAMRgyp8C
uYG0/squzMTj72RtS7Ks6EO59T2cK5gBPOHekc4Kwjn2vLe1ooACqTqRLdeF/oSy1G709/zhB5Jz
Kk46528gPuZ6QvUeJ3wplZJ6rs2Xt3ZV83HbIf/f6dvaJSlBVVA6SOFiYaZJ7ZV4WahlsXoZDeP9
cVvimwFIRUIDzGirY4Sp22J1KQkE3J10RxNZ2bEqW1RqhYmBpVsw2XlUQPv5Dl+WqiG4qdX9YdgI
vNeh8noN3y9wrx+OLKn4LcUrMdVTTW7TcggdkiBFvF1b3ZqHMrN+tB2y93Ig6SXJeckqE+/KDnnI
aospMiNIm8zhFS4YqkvmcVWns/axanJwLn4cLWhvEwi5GztEcFdnJDzNVizc8SdkPptwXCztraVS
sXjekiBKyyaP5TbmGy3IBTX/L4svWF91dbtO6PKWXlnmeIbdCYzYhkPGWKaGtsNbRaxeQnX0C0/n
tYEkTLzEvkFn2mli0xsZYDmjq/c8oEb5HvJs3l5xQC3QJ7/OASOrH4XVTV69zLRI8B2CI5JqO35N
EEjE1dvIB50pwihof66LPrFWi4WUMvqIRULGNcfQEc8LKQ6/i50KgN0oPZpdwDRsnYxJtq/F1bIF
/UlQBc3KlJO9mTNqhJjAVq7yD/c1rXcfcypib+/P0ObEHsLPmxr5lxGjDScMcz5iGsmogTp4IUUX
zAacpEOfb++yJXNRocZIL6W/SPQgYuFldZPhOC9nSy6E0g3KWI59xhuuyCr1ogJDqO0N7230XeO5
nVnOwy1WgTm+EOroFpDHIF9tm0HOAQ/DFyWEfJgkbZ0bfwaQVe/P4MtGZS5j1Jp2FbiiMDnjsxls
b8fde/0JO9MMx+ceq1aW8cmndLEleel1j1LqvAFt5O0WS6e5maMGqSTucgEAsA0raUBTkZpvyHvf
Oce4Gtw7Xr5Ith7iONV4n/rjsixmH8RYapfPgmdN6lFMq5cOBFWv6UpODp6VQ3KLN3+3UbX4dI4U
n9Gz0QsATtsTnjVOnOKxD4uPmrE3ow/4uk+h5xgC+b+HhSr9fznvLVJjtKXBqdhJC4X/imMgo7UI
f86puE+EABiG/Uzvd8Nj9+J3CWQKNSZHPRYLW7sKq1UUMg2K9Tml0464JLwpPJ0lXVzdHbTXgXVk
JLBjvDL+nTZYlM+3T2djJSGcqq5Vu1TlBtiG0Y8NxFj8NR0qaWo+VoiLSqhNsHMelxmCv82+m7im
/47DqkLWeqJldhTM4haGXjCN5nHf/0wn2xDIw8shw8GwG5dGF2Q9t6jNpgOVdr0MRJthhOoLC5BF
LxDMCDoC5pJvPfm40QrcxnzHJEd867k6eUmJ2+L5bNjeMBobVqluma6wBue1sLOxuq/X6oCYGUW2
BtPwdqHHDDOk7IV45MePnSxkLy3CuPev0bkPZSV/wpHDcoLMTsp5OmSjSfog9VIhf6YLRjnHEfF5
vrsUzMyztn25SiEXnVI5A3bDqoTCAU7eOzlGejTsqdGQ7NOYeVi/O7Hp1VtQLxa+BZJkOZm6gwrd
oiiAyzK0NXMp68vr31BCLwVMlcFgxOS8Evbdfezrq7mdEIk/9BfJpXbQEeD3mjAtM/UbbvEVWkWr
dAbKqcNjVNjo6Cm/0qtqdMflG1Ycx1oW9hHegIEH7nlKq5GtODQwUhXUHDYxWSqF3Vw/LkzJPMOU
kcMgunrugWso7BJbihjHA1jVN1TgOesESbomEEIhD6jCAFfIfReJm73xSHANbYmanYZI6wFJQf5H
/ZHkUM8wKfv5jXiTF/lQAPmN3RLqjuJMrx6qM2avYxwbLVaNp24Yp//+WYydeTYCSDLJhrvrpvmo
+DCnG3ttSD2NHTpsqyGH6yBP5FPKYWMqHZ6oQGMwBbjq3gcV/jbLF5/0UcGxTAhdK8EOI/8Y7FTG
Vzc1sLG92WE2YxalfGMPKA0WVdQkPNfi8zuOel/CuzsSyQnM60U2i6mIHOztymcmHDCgRHKSZE/C
t2gu3vJc24GZvt8iTNL984NtdaA52YgTag6jlkaRo/1F82jxsyyvEkiqrnL8MixX8IilcaHYazlZ
xwYg1YocMADOa4dhVhddw3wZDHBXcMtWmkGql0JT9flDNkRLazWUQEVJ5Xba8Kb0+lGwtONr0+eq
OSZj+CtNmVHG256LizoFap3l++9l42+LUX8tV4pew5sTyXH0wj/179O91Lgv5V6gDDHf6ZUfsVqQ
6koXkUw+zDh61bv93pyH3mYXavf08WKH3k3r+sBZxMSJXTHSYaOXiDKQ20+WNE1+CUwGvB9aEq07
R7i452To/f3H6RKLUKtaFrnDoOXDJTonRyyb6kFL7gTi87lnrNZvwhuNf4g9coDw021FxjgIGVG+
xJnxcOvBSHtyBVAojp/0fcZ1hZPyzu9oTKET9m6UFkPIfCyKS5965eSXCq6gBWBlhizNr08Q3G9y
3T3dhuJZl5BKpI+7CBu/HGcLLF7452taihOcuJxQDGeWusqwu48nBxMH9kl7cx0QISMA1J+mWM9t
t9e5PH0zINrhLH+ygJD0zFvg9Xb9h4feVpBZkXGQXsMQLqiFO64lHSnnMozpaV2FfGjmTSNfiugO
773qUH/JtMRt+6YHhd5Y5hEEe1GL9FrNmDiXcDSqnSlvJTUsI2maNyRXnYYMKycs/wJDXIFXaz3V
MhAPY5xEgXCqhS0hH5AWtp4EXzxWMOPcbrqflPkrYhVZLwDWzsuyn3oEkN+/eDxEgJCLuPXrVrdM
5FRDiVD9VoLouWUzXYLUmhxYCSeAnBMkeIpcAf+q0AmtEIkVizK9dTxNeHjnucQtc5il5VVrryc8
xp/2jKLv5VHRypRDOHZQBBFHX/FgoDpOx+Lfl3GzhNASAMtG0UjFEdboiSpga9eYuXI6gQU+Fje6
EhpAsucusKD0hqXgWwm+6y1oXrOg7nh3wCd4t0Su8paqecr5qMkw76LCVPZvO+o7ikd0gXc8yjug
n6acF0N2/vTsiOBOsmTx9QXbj7wgcUL+rkl1UEt/vy0kwOA/fyV/y2ns9u0DZd9fA6d4yvbOeQEK
4TBAiZNIXMgPASiGhdn08ToQ5hmXyFjv1QZw3h/Qjp2gjzr76LozycH6Q3QudD/RjW5mRbFC9h6b
3Ll+TUmNT3dZO0jV8QC1rlHkfdkBqO/r0nPVi0XZj3AREuSg4ynzJlQrF6WM9jyH9IMD4II/9h33
YXvop+2jH5g6PY/vIF8RkqDnIsyHSMOcJnx5O7kAh2nWHYE6tdpUEAr1rh6b56Tye9zPCPS6KiqE
ePiLYTIQRN5Lz+CwC4dV31yoOzMZQhWz46RKMtxrLoMAQH3+7IJ2IV+g+b21iHO2lawmXezU7dWf
awu1ycaMslgIGhDYLvj4c9czo+75+Rr69XrhCMew5Xe8RacgTjCqhF6masAS+Vt3Voyxw7o7h1Lm
d/Bt94bffWy5jQmT6DzfpowkM1oSju4YoEhReMf9U+g/Lcl7r+/WUJOjSm+lpN/wCgvA2mIJKozH
2rJoisrlstVWs7Y9v+nVwJPd9QFy5ank+dlxw0VDNYQeXrHKbmKhR4Gl9g0FoLiRK9pNtbzC8NZI
+Fxh1eDLOlqEicL+PM6yinoAk/zgqkhlCOs+UpK/Xg8ZWezjCOfo/D6SlFUwQOvhxSWGD+RGtC7T
sSTHXjeNMAd29HNvXWWLRksAhW4evn0v+0y19CN4UtYvponmxqxX3DSA73aJox2YcNdNE7QEdS2F
26H1i1geqPCIwtkDSBTOw0DweOPUZ9o2xSB8D3uIEOFTdk/Nuw7IRvzb6XYE6+zRU1oQEIGVHJA1
KSvBZrhIVPbICD6udTYgGzyeuszwNbDj5HFEvVfKLIZiVg/DexT6MSCXQZYFi/rfNMUvYbEUbKA2
JASKyqLIsnLU9jM+J6PDsgCXAiTJVhQcQdkenFG9vWvDQbU3TxE+B3IhXRExD9Kpq0N9FTJh/zWV
ZpwsUGISaIjnEiaeGAlq7RJYn7WahWtAlXWL1Z3k4LV253f14b08LJrWoVCjrXXSzaLwXx4iLSMa
i2rtH4mXpV0UIuktCb/L/jBMYhHhDMKaBZn61t+LOSAYxxlmw5ZieLQjratPLSrmm1rZ92XzchBR
NcGtu50Ws5EJYEbeYBx8JRAUxzevGWutsIdDxczVYi0P7MNwwlV8djZfv+oJQTFK5rdYANLm9p3U
VDXhhnX8pAm9ASMXJdyEQuWXF2Zb3kEbmZx8DJGzUHWnXyoBHsHD8P9qiTqK0NIQ3y57bcWMwdi1
LXQ3tasa7aIHyLlAoOAaDW9SmVCaxKL8FBDLV/7Pd4ZPyDrGdKMAYk9CyFeawVKAOrPdjORQRddX
n4r4wnJKZOjAekBEZ2fVNievNBTEwIQ4AkGrbtxK3HEyMaPdm5sdx9HBlsrk4oARKeQrL31QaMEk
XNPfz7IYzPiNiIlWlykKnw/uD3wTdp5i5oqdorIqtIeEpzmGZpJKtmvceI/jb9K4ZQ/HoEbtWzz2
x6xnfuddn7YCxD8pGgc9DEFS9nlfC8tDevYGQORatxivUZediODpG+SZ3q/0dE60xpr/k193fYhQ
VsV1DNfzxTYTCe7wQEfJ8DfXPmCCaOzccZ+mf2TUGHxYBelBXqUasqmqn9qAK+goy+Fy4qldLjot
bsONAgwQnb9RA2aNmzOfVVFS24MIzNN0sJeexpvJLenZ4jxo8LD6BYJH1JhQBMyJ8E/FxkH4EsrM
8J8iSnkNpCE9Hh+U5ch824DCwtQPttYgx4Afr5AMAx+GD7e5f30QPfRJT3JDO6WMYkMgd2ke6mHr
m9O5DoUJfl2msajmVGJeWMEW07CZKvVKWGESkYcBSBae/OR+r02qZ1JsdIzJOJY/jdFdGB45BTia
a18RrrYCL8U1+kWAEQAYUYcA3efWvsAZfArIAt6Krt3TcYd+Q0hw0H0m0o2GF851oNhD0d8LUrp9
+fygCNQQmwphh9Rt1C70jU6HjDfWtAVnobwFScxGiMPEyFUmpGCDHIp82GU4EvvuyQ5Gi6634img
13OvmRERCCzfKNe4tInv6bkCDH1vM2aSsBDntDZSkdFuLReAdFv62KW9ikT/uEyT4agn2covQ38M
/u+cFpAV1z63dOp8j6sQXzDYBV0dQ8NNxynsTv7yPcIiogF7rPcb73rNw+9Bgo4hCZypuATRB3zv
ndcCbbimK+wpNgZScux4tNxfGhEAliNlruLhF0jZHOkC/rjXrBN1ItGVKWhvRP+26+15JY+3+jCx
ntFNo+arHoVL79+v5S71TColSSFElW0LG69T5BMUljH49oSxJP52ojOdLIiLkCVQvVCbpbjhWzLI
3ykKsLLLvIiLnW/QeT+443ykMfMeLVCB6EftHdE2SaA7nWGWWYbw1704k6lHuSO1GFSDLNF1g2Jp
oR6bpryHfkUTyVAXUukgmz2aVZ4PDj9eMx/tMYL77uI/WIVgC2VbllEfrRSv68B/dyK38QA2mhDL
ShRwhuDuG879rY7TeKWKtGE4BxHDqPLDViGOWstnAqg1GGTr76H6avcr5gCyQxf9RNeOrHBprE3G
BQXQ06gak/EGvKU57QEIGlLIM16tI7b9m+14wcU2RVMN5v2uyuEVlh3UiRwuBSdeu0p0A2FpBM8f
FPisEshlr6EmHesVUFYQOtsG66De/ZC0kLjU4dKgWfSZY6kzfedXaYk51hetFyg2H3EdThpIGT6x
jy9GZqlRHKEYpAiIqFf3/DBgqIqpR+KM/Q2R9zaORjTS8LQyrL4M4tKDBc1aAXvapD+WweX51fBh
zHpWGzzzO5um4EG2PC6EPPe43+Z8F+xwhLznA6W3rfkReHePGGPEizHoGZx7wND5i2ORsDkKzvt6
6FwV6+V00V461zFpiX7CRJcaqmPfrmSLyQNfKrk1e3Mo/4D6utTManJsIrhqRyyA04Z/rsqtGVQx
HAZ6iuRCZ/39hOoWVSOdggT6t7BZoxUXP/izysxoDiUZYjvWK/TX8NzpMo1YI+zQlV1WRQg3VvJ8
Hy50irOrUNGCGXL5rnKFdI+ZxAznicQRH4F7fqwZp0f+ltxF9+9yDCB6h3DRewL/IPsc/FVClIER
fumxsZtuD4Qe6O0U7bkTjHW7OITCn6PecFM2Zhfn5tLSRr8ax+ZOPjgfH0tE2WYS6NT0csV5SXmk
fXzpm9JYaPkI1/HLRjAh0D/8QGgEr7EozzZHWmoweKMoglKcaqcRyp8l9PGq2lu70fXXJ/XAfcaC
G4JnI4k4iaDltGEICmDIKJI93UmIeTbn7v6LKMJ4dlc9+gbhtn3G8m4kGvJwZ5Ivewk5hm7q2oFG
QWsG7M5eKc0xy+ZhZXIuXOhLWSkcQ/4KuFZkixsvg6J0jZ3hQyFs/u5t9Qt/Zph+PgudTd2mUyJH
H3bPqnLq1NgeSn+G4tYkjNRqYcikTLUIO9iLQZcRaf0JZ6pg9yTJiaNaP87HoEFk6pmXz3x9fl/f
hU3aYHE/B8W8AkbMf7NJbtDbnlqkJafCZcJac8vzoYBW7w8mPr+/LQmatujU/eYG2DpyVhHrl6+e
YuZhqgvub3meJgfyy6HEmdGma70qnJ6MSGz4lilYUiYnkR3MF6jED3FvO2bkqGpHB3cGW3AabSC5
qVRng9bLzedx78nmXQqnW9LUE4+B0u8LS5CWlFQUrf2krX73didaG/3PThFtPsJbWajDpfrLnSn2
tw7PYHgcBfjgSuLKU/3sehCraiRBSahTAhW93C7U43RBytlU8Ygtk9RBQnb9LDXZktkKAnN/B4kp
A/crvDuTKxEIOmxRJBIZmONv8CErDejRRloiIRMwS0o9fojTt7k2gR4/cja2Le7mc078ZYhRzppL
+M2NgF7PQfvfl7spQp9uLXgmD0DvViQWrVDlz8bPFBMV8GT4SCxAjz8feseYaoVdL7VtN7znO2DT
wMUUEdbmFMuycWiaMsfgt15NbrgvbaKk0u3GWUqMAjm2SYuOvxGBTWKk/zsxB6aic0egxRdYQ4Ov
Weu32N0svX86GWbTw3DawkzV5DeJ+RFgtNPavVneEbROBjQFUBu16k1upC0hzuptDLOJ10oNqvpX
If9grALUIJoP6RV97LFYjnRbnmBRm9VgudW/MVNRQa9n7HtQUN/kJOfqUUF7BJUqqpNtbNefq78a
uCgzc/9fEHDzmyiMromK//AfTSMMIjVGsPinkjpKCUektuSssvjR3sGZWnUhVyKNsNqXAy8IAkrk
d+8mJTkGvxAoaZYcy3HPXlZ0sLd8HVA/Q95jhbuQsnrD8epR4NyHn8LSOV/172TCBpP/BqCP7g2E
rMPcB9ka67RDy3A/gTqGhb2gO0mzUjdXgmbHMQ02VzJL4WLFz4vZCyzMOT/SLnFs100Dlpjd3E4b
+KzQRouok7J0EvJCIOU+SbWeT133H8iar6sCKmgDeOL4vVLh3wg+c3SYFckCNtRniOZf3/y3OVhQ
qNsMvJVqZFiEAlq0i8RELXzcL9A5BzSCw2s2MTSQEGCzVlj69zze6PulUI4hmtIpom1p9GQ4lkcv
nxZEEOTBZqbsrOf6sd3XIHJNdjfSnCyvalC8cKwV9+ivx0I34pbzb1dj6HEis/ROth5MOptkDv4n
DBxniJMqs+ANCTewAsERkr+PeaCrF70nOWR9juDBZUzGeE7J2bpvcTFOlrMCkri2zAwBPHOfgxs7
EFs9wjTHSjsBP3BPP5wNhbcVXDA/Tehs9bEJ0vriMXbrIhDROGU3SuGY7dKIQ1Qskwb78r8TOE8X
Yy1sQtx5Wohqfahg3Zbe0das7BtPXSeR5Vwi9od+P6GbiEN5L4KqEKmPFXOMyNnTmgI9IuwxMyuh
hhpEHdfukYf/ov8br7wKA9DW6XwGbj2w/5UtJ8MNWTX3QPPnLuZoQS7gzxmAiFLYdHSJJXWR86T7
wcZvD2HHqnH27sdyuFGZsCDNOxIoMmxOPJ1LwWZT9ymwd1itztb4iQA5d3OQSNyMdkW8okXl4nG7
v4Bx8jlJrDsJ0UNtDPZJpV+XTUzgqGfHQNcxUgJN1TrLRC1eMCFmzqxi/jkKhPVVaYR8cAHc6EkT
Tp/rGoSXLodp+7jYk0Bpo5ZY1ymUApJDH1QPlxH8FqBp365Su67vfTe7KKJm3BzqzDouMUtfzpPj
XVbRPdDlA/7LEmGv3M2l0Mq4MHP+u9ekWZHdUvMx/3x/4nhX+CSEz/5S2SALmDdEhkyxIAB3im0j
uJOcV0q9yXFNSKY2TZxkEQwUpiHx4U0Lmo15mGvRkx8021Hyv65Sjp01Z2eTtFaNQJaNJyfsM3mF
CbL0UhmoYdVcGLV+9cxt3wFMWHeZGAn50ZsHzKFnL1cujN6IZHmpeQQjjoTbhEqbffbbcSL628kj
LBgI+NPKJ9xV95NepN/tnDmyXqXqM9BGoFLmcGOyfmcwZVwERHu+2PKDu6pMc0kyFR88NzrQw+OA
wlWJrXtKBt0qoM5fkNDq5Eivkilc9wuNOdjudxqh6h42LGoKzjfNWrIMwzzW2512HDCOOwDhOtFS
l3/GJj9Q8FMPniLCrwRGmIsQljnf1gUno5He2+xkGdWplN+xlgTZ/g9Xzz+2J4qn/TtetqCCM4KE
s75MXnT+LEsjlWwWm+km9ccFsAW9xaYWbFaEJbWQHTyLUgbCBWF5Bd2cIEzoOyMXiCE13BpW7n1C
CXXQSvhbVmvOBQbZFGO7oUyAl692ShxbU6xDxRWBKmd+hHcbm2cZLK3p9uR+/EnHsumPAo5jZ5ir
g9xS6X15Pw0xad95ZsWdin8nGkN3rVLdaM4zaqLNgyVymCRhEqPpWUtp8tLvS5UDaXBg2n9PSpkO
Z6S9t1SmV9kTqkRdAA6EW7hNLvBKom26hn4UZ72WR6ck2JJRdrPmr5/XTivKZiUXPpQiXPcYRwep
fToimJ0mWBfaAZC4MkqlqncO8ZyP+BQtFg8O7cSy3ss7R+Z9W4pezAmk1/uRUDer1Jam/b8b4z0J
xiHVGJad/VIuKQHWoLcPGHj8mjWySfhU057Gl0PM9V9Mio3TBm4mC+wLtk47R/4rkGyu0xrxOA8l
w/eZWNLwtLjStZCf8ncjztr4yIkZDJ7Q+7V0QNMyYswjSu750RJI+ZJO0l9X2uISWMFW/GksJgeP
m49hptiKjlgdRh2ViM9aVFNuSFjcvIk8jTQsffN/tde75HZ/nZtfTSWYOaXP7D2ivIdj+DKkb/Oh
wspzHZq0w+ktof4hL7qJBzAd1LOSOCe4YfmPX0U8NJzAoDEkcwe7o1bGvN5sEoA8B5MHl3pRekgW
SaQE1k6M2a1doeKY07g0QnAyfDgX92mHnB0N0FynCccol7D9qUTBpKDHtUTYlApNnTGDrNdXvZlt
wFUBjktl+0LNArXpkZG2Wr1bIhZc68ZVZ+83lqm+BpxIaQUU5AWd2YyPQpfy3CuuzNbidBjHd2cV
ZRNNPjc6v49RxKgh/81NAa/pH3Up8cLd//Nrhv3MhHfqO7FOdXA5Mevs1RGTIzYUUX8J9KZ0z+hD
G+MyMJrazxe2dvucc2iba0rW1A8BE+da01wwwdbOpY8KMaBuiGlWYWsXtFqoNwEHPjt7ZvycsxtD
db0gUgEgmMvDbMnw1GBs826q/2I2CCfc4LvLY3OFj45qwZlsx98KszNLHL46Ely3eq2EBhdCoh8b
riGQ4MtKCp4uBlHCaGpAFfywnytzVat/J1B64GuZz3mJV++ltRyxXew1gVjceA9tZlfWxnxpW6eo
wq2K2f23EqxsR2VnWeZRwPdgZHCB3sFZ+4ioZTJ1oVtDto7y/4AUCrWTOr5q3VDXVl7YaFh77AcT
Lk9LJtRLnngvPz5vJ5gck88Q9iMVKVFHLFCTnFXfxOTW+YZR7Gpcz+QlN0oPPUcKcQfN1UVSPcLI
0BOAWYygf7U/VUvJWRXGbzPZ4zuOohb9kMggk88PvgL/OLk+1bvTlbu3RRFm8bSbGSACztEpjQxw
kIIs4QLGCU1kXRCMy+nEbEJeohOTOg6fL8AeX5kMJTCTVPEOQraFMWtENYTn6Q8GgjXOz8wgSlFe
/mLajBcdxkK0RXHyhnXuw9tf2rXYMyBV5rxRBWCLi2KH/kRTzl4jZzt3FRR1aI24dAh9JN9F0QJl
A9RoKq7sUqHA73/lGvffTa8Q77WqIbSpoqMHSOuJ/Nv44UxrcgXXgMwV5P9QcvaS4Qptj6k8oopX
0oOVz5DxvNMHXOgIKwgkkJrMRluCCqkPmzZ8VpbUgWOVaMMHKhpsey23AYM1a6I7JJfmkWfjLJlR
pUac2Y7IqiK3YlErkS6f94+ZLdyraJbgxYEL28AnquUWMTec+SJ3MSGSQxMsNG1fxIBGXuiVrWwN
ho4wYRA7xuAmzIDpeH1nLKW8wDqHt6ZxjqA5Yw+NENW/bFaaaPbOCfG1Z+oZiAWEoKtG19t6/PsU
+ecZgVXBt5Ln5IKR3NkQ+DAGo0bHKMGLIDEZH9sd/vhcVBEVWXsbcQ2nzjpvJ8KphT0yyovOLiz6
/zISRZOKcZBIJcNrKRDj5mtbvxCNUoSvFddymAw05Uqb1z+IOKFW2ePY4vy9sAHcixJsgA0MghHO
zJvvqTcwaGBzlHdHMu+q5L7LwDjCHICIgvtitJEjPaTInGeavo2vt9XwGfQFyhfN+47ggFQinbx6
tx2mu8cY7BSHXiHPq+7duysOTQGpEh/GlxtDLP7Q5kntil88sUikNnYqa0NyS+HN7USAJCbFxsiw
Pr3ybRnCp4v9L1jerS1c5LPJaqRTicGgrRyRb88r74SyGm6xastiXHRYp8Be+TSDjbApJzhDjDbz
8aXaL8/jzHg2E7Rz+CyB5MGxYwYJgohuHK+oXfKB1Zj3RWOebkodeMOKgDA/OohYF4C/UQCCvX+G
GKJ2VHxFIcBq+56muuAXDamuRuQFFnU8EJaNe71coZQz0oHS8qRfIWsUfzLn0YyyZh9hpEj6cQHJ
gS94bCuKSwKHTyGiKIN3M8cs8aZ7QbTJmESpTtjkwRfcXmx2ULQxhWDA9RCYqBLzx6ZPvg4/9n9G
uyuN77E76FGVQQU3I+zRld3J0CgscLccrcjg7OHEFmGC55KFteeY8XVBY5n2eMl2ZTiACBsbFW/o
8oWg4wzCyVrCHyn+Pzt4YFK1gyb8Y9ifOig9Pq6HxeKPQ3lRdAFVjQcxfYGd+mV4bXnCU8IRK+CV
eUl+f33UtEXP9J5Sl/ay+FIxZBxRpFNd74fEseWWCUOPcCyPQDY4oi3GLTomi28Phc5GjG3nzfdU
U3oQdq2PUQeCCg5SGnEfYwf+etRCcpVQ2nHdwXdhVZJiESGS0Bl39tl0X/qcbWGFdtYZl/ILWT9W
UJ9Dmhgok74aQtbJ+o9yr0gsRNrbK72sEE9c4HNLwEzjREcXG5GMQAKzktcbOydMck35PMroPeFm
wS2Z7d3IcXVRc3oZgpckuwgzftZo0UvoV9p2dHYaz5C7qXxwOc+AI2HdSxl5E1pIQxlLOm/bNP5l
Vpo7muv7DBQ1dK2MtqvzhMWU8aqvH7aXvObDert3pqpNeMQzNmxXaMqagjBS0O8xoBwhKPBrS1T0
aT/F1EriLjzAg2m48H94OodZHQ4N6+BvspQsP37Rnlb9sBD7LIedkDJVl8sFKFe73oBpnPvVepXd
XfjCps6cZvDUO8vAX/i+FqDBOBz44SPiAd/7vlL29g7RHQnw6q7bSwZ/ntxvpDSmHw0oUPS/Qrqf
/5GHPv0aQnEuCIilmZGqc2/h0Xvz1gdkJU0aM2AQbb6JDyMjHMmjGNZmI5qNRi3MvKJFxnFlJl6c
eGw5ogUSyERxCOSWd4jVu4ecMTpWggM6dFgSJya8N5tH1zGIeH4g/L2F+ujb10aGYfM+r9WScgRh
il0h8X2A8czzTiMdhAAeK+enw/EJQUkoEDpGnHH5jy/WptG5bqjvDQht0EUgPuaWpDAp7TzX6IGd
O6Z/zwXHhEPsgKszt899T7jJgZZM36FMAXT+0+n77qGCPSDVUaY296aaEzE3Wsgvg5wWdnqtL+7m
u53Als5B+YBrIswAOaHUJd8oAjHOBBqi72j5tiSOStZcFIQHKjqkGKoVnRnDBnDWhmTTvc7zRhqk
9PakYAD7mt1lKl+/Y3rsFHJYmHp6JqB7WmHdfvFX3YhcfyOa3qXksK9pTL6Qmc+HPElPwXedUqND
VFC8dS0RFBhViAg26ai1YQzoKF8Z6mf763vWVQVO13ZE5NOVkaZskHtrG5EXDd75o6jRnTR0ejQ3
dyVy5iZgTI6M4282f7rlnuTjSD00zI5bLa92EhgqviLkg/lCylT9TGcQVbN0hkND00QN0MBj1J9y
k37GqRzb7sgdxCavvphNG/1EbZQjnAVd7sKdlEaqDK4ah/srgPDnsTNU1UQYBNCjFh4RZJ7E24qL
bNOn2xQ/a0k8QlJkaFh9sD5GZQUkVmuedwxml40nPfp+U1mxXB4bDirgtHs44RYBlVVQPK9WCZc/
KM5F7Ys06dIq3nizK25WX04X1c8DQLZUTWe+HRpAfE9d2isxcrsMInlfBVzjx8/MdjOpb/A2i8o8
UALX7lbItbAeQWqDp7c2HxbDG+0xtSO4kmoTftzuLlAzU22YOjBjFK9oB53UEO+yfNSP30mlAepE
ZscnfIh/XNxrpNdOTIoLP/FgG6i/XlUX0Nwn1riVvPgJeLyZBuMZ3gP44cBnvbuxHxMs4GQz7mhb
A8vmaTdzQp8Egqf7JpLrYZRUeiy9P2No5+TSTyVf+wVA0LMD9hXSySCPdjUYWElrVEZrodovEv1Q
XjZuv5l/V6cI0knVF7hJyFqaziJ/8ID21TfOj5mhNouzEx9Ca8BQBID7UN3kJAkbDS4EfKu70Ju4
fyK+Hi3XULr3fVbGkP2YsbmOfebCvFw2j0AcMIMBHkNeEEdFL40sXemZ++fx3H5jRXnnJ0oObTta
HNjUpUNeplIUDgD1PMHQleB5/AjB0ZLAxe01wfSYFRHPZUmDPwIuHe9Z/8pfYHyDnU9grN2V/V5j
lGpHQ6i+n/HsFCKNjf/p0FWLjhMgWcbfusc3pvxcy0aPk15/0ahNeqywFAzb3vridNaBBoAxbK0P
UgwO+OAgoOWz9XlnJ68hjebwEDDO307MVp+TiGmCj4gN/epYyyFU/kIP0x2Ba8tA14Ivd1U6jClA
T49zPefCqSA7j+555jaZLdsHBMceNn3lW3My+vz+kNCergcNe1HRYu+4SPkl2s6BL5/wxWyts04q
rsOV/HeaKi96Af4QFojPD58x2NXWIC1OH5Jzko19NlmzVstqlN1zcPCVemfOYWLCvfFKILfFQHQV
hIQxe39iETsFa7gMAHNQGSGKh3k1g0AoEj+CuA4v634BbBiR284ZEQaZGLrYPlqtgCB3FzAeIOfO
SaMsqabFy3DvggipfO2QvSD8UAr4LcOkV7ychC5j3w6lsSnrrJ5a1RGKYbOxGQFht1Op+4hOILjR
QqKW+nh8uGQo2GgKQSYljDnXhlGqhnxAUOyHZbwyAx81+4P4+EaU0WOqZVV//67QaGNUDEolfaCq
JYGisDcy3dLFDc/jvwX4vLrqYFF4Y9aI4d2QvVl9YVb2zFFv6oZ3YQzlTxgV0HSYKxzmHloa5CwT
s4R4U6GBjjjR6KT7SJO9vvJhGhtszrqwcSA2gHRBBtWMnGv327895htItH2H2z6tz06+cMWyZrWX
6aw7NIwcO+L/Z1PxGXC6+5xgCFNoPcy9lAoOOeRS/e7tpWG0yfXNJo4TZM18wnvOsyytI0gVBx4Y
4XiXHISVeVwYw2BMx8sxW5X4+0/An4RbLYIb6pRmxJfT9WQrYjhfmZpUf1R/UFzpRmJE719M7cgh
hBdg1gZE0hE6CAP9TQnOSyatxY2R8xrNQXCUMOo1gz/gx3ZkLPhVnzEPUorsslwdDo38gT21gxng
AM45zXKkEExQFWY0EnqI2nEkXa+cDBSOKOPUWRcfrBLkww7XyoppjVKIORMb4AuCQ72rUJKqtlJX
PcBVn8iFh+7TeWWl95i6TXDvHnEZPTw+S2f5qcpNMzxP2Lp0Cr1LaazVLolW0IFslecgx/k8M2Rq
5cdiIK9M7mJEaUahpckkm8tm8Fyt4zRMiJKTcfiIP9Yx6CQc0UE88xdqQUTuY1XEcOfrClSMjOkJ
taDccagtNQtXxI96GCi3QDkqsVev8tEjbI/rzQx0doRv2sPcedIp1isUTWb/+13EeoKZRNy1Ekc0
76bOsDUgCavLtQ1JMj6sYX1/se4jgIShww+cooSbEE9m5ze0WR0yPoc0Nl07CzASp56Pwu35FAkd
CwTddgJC0dzd7WYKepWtXFm5YnuCZ4LmoD7poBAYnDK4c2aHaOyslxQ4n40JgQuSOzKy4oFpuV/i
CtSU88g2ccvAZO5+qnnWvs8lWenDLiiBD0ZR3yi6u+FYbHnRWfyPnetooQD3A4026D6Brt9AFSRi
4badcSFzMv/x05OLwG4whMs8jF40xSFU2W01YRU/RSUCnWrKsJD3kGPqm0ldT4ArB0dnN+GMHqHC
023osxCwZJXYwVEDwd/FVBw6TBPXViY8yCxAJD4KuY9wW3HNLvZqNMDp10ntMzyRzuCy6oZZMYNF
00SVE0bT/0D8X0p9V869h4rV/Xuyf5NtFogCSpIsVZl9KIUoy1Kza5FPSenWeyjGnXDzGmJEig+V
QGZNSPOOMCXdaQvH/nQNXmky3ES1pkmZggcIKlorI6IE/OtGkd++O7kjZWQ1eC/H3uv+IwTU+sDa
//7r/to2iFTqIasyt6mAlbvQplnLb9AXgXZuiDd5mfPrPSUOUeIfpLiPTfKbi4lDI/QAdgqRJqej
XMlBOVLIg7CNw+Vn4/5xZt/Uh5mvEGfAj7KPasNLu234PrsAox2JEXBbXigJ+K06WXG16AlYez0f
V5fQulWsdXMVMbc+6bEdvTThQHfaWg1dTJ5TbkDnBPNq6BqVnJhSp4JAcJutFaagNBx+h1y8Wnpp
A4ZgZZXbzUWzadkb2gkAtJced+i7Yhw74I8qQbCHr4wQ8PgrtgcpbAQJxHQ4ckuutaFFBQYu4zvb
lECWHITTTgqmyNrJKi33P3YZr+zka2vp7OJlWnXBCrA20rpSSeWRKcirWzsjsnjNW3/EiRSWe1j2
VieoA7M8gnFzimukZc6pVdA9Jo13sOJ+faYrseFNdIxrKq+6ePTilAE/cm+rSgDP4ilBxltBxx31
GXhKND6YhTnc8hgEhL742yLt9rdDEiENMDj6ExEKgHf9UDRQSiGUHRxVjcjBoowIHH8PE16Z5LCX
oVv1PQjHCDkH1qefylnDT4cPI1UeTVGL0sOM22vUmN8xRxOJpXDK4vWWYpQhwTYrOhzpd8y5Pb7P
omiLl+GDrEXyvwcE6apKvTldyTRMTBryVTAqi7jO3TblQfdPJ7WYSn3a9Dup1FeaDy+6WRcfLJBM
dzFvBh7O9XdX42HAEMpFTqxBKs1hsJlKygLBqNRBD8reXlV7pijtElBBh/13eFPcBD4PatIMVu1u
RB8XFth15N0QPt+wmMSjrNLGUJvcek6Qw/X607wGiTwNQX4GdvzWL8D8sYjvKmb+LWsgvvqcczCw
7s32hZ0H84KooYq9v7wd+3jPMwsUF4Md9u/GUEM26JquCsa+sG9vQ81Ce8JHgnbvaBXzIQkhMw+U
NOGktMq4TdNIxDGpqDXtL+cADtxriyLokvsz6OqT6qBRWJ9NkVT9CQtBsNZhARoq4VUAnZcJWjDz
KTLfjfiFkyB4c8UUmcZgitaQwk1SA+korNUY1P5BlEzfGK3Hm8htdIivaIBFrSkRw4yHDVpxS32E
LukrGGIOLwMFOa9S9KHcOfcsf+dfa+dfKm3dxdyxyGIzvesMtYGNJlH50ocEsPVAcWRCyzGKK8Ob
t8m3FkieplaG3wqu8Z+hA8277hPRdwU7M7EouaJlmbnh5YcQZ7m5xInYeSQxSPmGpRIvlNrrhDGj
FogFUOa6zyqcLFARjhODe9z7Qu4xLKVzZBHTZUvawhuTORNl+tID68f9tHs0Xxtxi54sY3OfN8Zf
/qyjI0l/CcEHFx4/Mw1pjVQD0zgqSb+efwO84lQuq0YkBgBMnj8ROcv/4mi+H0tNZEZ9Hnlcok+1
IySqjY/B1THmODwi8F6oUk8qZ3CF2vllnqqIYHeqXYVAcCordjIYeGbKgd/ymjiNBGRXI7XVvAkU
wa7tcEVSV2FIwgXjFkEzX/vWhBevtL3FH5c1vbqLpTDJ5qG1Zw6lXzBD7Z8ygErtLsxP3DFF0GW4
TBz1sj87jolBLSqnL2PZBOp9GzM/elfUiTQrEuhhHwE8u8jrGibTuiTVCbt6uirNLeJUlYhHC2t4
d2wSPHeOoHJnhzGwNDbkECgF5vOREGvHjRB/1Im3mNrU54yG9SK6HuVnAIJBSsW0EU/QplausWS2
6Gk3Fj5+4Ovnxa/CZVrOdpf95exQaddwmxjZUzBWBjqz50cZkjC8I/VkbY77WTrabPzqlzAUkAYA
kjS8zDaosHafn+q1P1UdCuL8BIWlhD5qQ77FjwvX7AsP/LzcqsdTfoCH/SLMZU57bBAzGUiBR29+
N9VZDu98/MP9MAMMn7YqGTWMcX4l2wFkmZ/8pbRHa2mKwTg7DlNREzs325U2sDPEgYpYiKFbvZ6Z
Ly/0RY61xNWqlBNk3fQt/hO3b5aLJtmHw/5RM+NqMbqJEmnf5pPiMIuOf0JFMZsxju4ScVpvDgpQ
RdUJkVjnp6mmMhRa3y6akDz7KoxQqZN1X1wREgA7yvazNsRxlWKYefqxonnBwYnqulcnvNztQUeY
/DbwEn+eii0O6jr2HqJdHNXRLRf28qE6x6Krz2FIfqrRIkRqtKFLsTzjkgkxv23jwHO+6MXv/QA8
0V0P4DAGNQ8Jz2GP1OBdxgbquU993gw+0FpQIpAufAvdnT9PDFWZQIL5tiAek6J+mlUd+vBfdITA
T4kMGhMAMCdxOob1jvvxfJ6iB90HcyxIGP9CwCrewiHx5j63/PdTE2NO6Z25RUkwanPIOsAD8Ebc
DFXEeJAZdGFyz1iihuE95ecKqS5PkeAA52rWgXPvTzTLzIuqZpPii8deWkLJl+P3Rja7tjCPYa/q
g/yjM4jNkpXLO3BaCCOcAIFRFkRPKWWguZyv0mepOqBfdG/oIykL1CaTjwxCgYK+qqPqW/2ZR7PI
glE0aJ+ZCs9EPfivKO5d87HOypsR02ia51rR48f1h+emuWF8qXQljSz928Yf9L0sFP9atLRwMAgd
PPetzmj3QXbpVImyYdVHiCOxKzt3F3p5ZORCRCVUU6M3KcjnTBryf1Yq7j+QdrbfYxocidk3OkcM
oUsDxom7axbKQ7Zn+LQhY9S+dQUjssa1TySwh1Y76nDThcXGo2G8wOP2K1hNX0PEL+FTvg/+TtUb
MUoyqvFapK4ige7A5qnOjnn2FI05jM8PJwkRCInJjTPlBZ++l9lA1tqoMZNRFu+khMQpgRgXp1JR
8HgaVXidcaNWFi0/prjCDMCY8RPPZWEnUJJrNt9sKgUmZ9pcnvWwc7NriqZZwmNpINIrtLqGJgOl
c006HjYXg6tg1vqm5kzoyW0AOnN7Kr4lZXKmLhXsem6uQf7ZdSqxUNJ36Hzrah4bWHQ/h8/3U0UU
Fm4gKLcuQCZFBsYjTuqZ0B0zVxMbfw4i4e+wK2RFS5thQpkdAkIWZdrDrNaXlE5l5j9VQv4kkSQQ
vA4IhCaRrXyWZ2oGMP+ikX4znqC+sEoygoZaodlcfkFuDKgRJYuavzEReUIr6HChipsYxzaTN391
BNcn50GO7k+ZO1yMgKcKbWo9KnnMHTFj3Yx82/9ehjqJiIIJRl9nwDQATe2CrGeFEtvvTWLaM8NU
GdpPuG4wmmTElAU+XzyDourFz2G620zx5Vp636C6T+KmKxqTjvmDV3msXfS+gPgRQfzd/1wJHd6T
Dv8k6/yklSOjIvIeKmnYzY5ZnqrsarIfHv2kIg9T+LCyH6OtIXHtWOk4mMfWtmxPDbqk6vzO7Lsr
0Fs1aZcPw8aB2EDhc6La7GRFnKQge27Fz9LXqNW+QFe1824tCpCxYcByxuAC83IRCFeuNHKrcyxG
pkc5dIcuCx9YketA2vKxenKjRZFF0qy7easbO9e6T/h/FoEyYz7KCErxJkJs9tZxyf1dwxgGi6JT
Bkj03h4KRsRIy/jzvcVvBtkGRR/UDMGnDUKNlU0OgxErSF+7AZf8G7lniCBYIFifYtTaRql+CHnl
tQKIkYxB9v2kl6sQ1qHcta399ngizfA8qoaVu7qXEk/6xhS8Gp4VtQUbSLx1+hntyaZkTpaoMeO4
3Ap/CIX4/78nQUHPi1VdRimZFb8reM9zF/9O6XIoGtG4D0pz9J2VQ5C0S7nr1EecaCvdrYRTDwNQ
ERchU0gurEr38np9WFTTuZNkwWf0zDL3HRBZ1ZpNM0dPtpd+4bwROwxDT/Rj9Ee8lL/MaMbBTrVv
kp6cx9P3bbOELNnR39EyZzInnlz/aK8Gzx3sgnvwM41oa1KnD4LqfrcLoatrcArzVREuJyuQpREq
bK/036epMsblEUdmIuPZaqQ67QkdLkbITql6rCAWbrNJwkUGAY6QNT/2N8mX7AJaO5vT9K1WQOoH
GNRppIx5mQxX+tqWP7DslDvTzef2VVYOezUdk2g+5lNoV8kUkuA4JuRvSJd0aOgxXO7mfpfMAuzG
95XJGh+RLB6KoroIB2YUegoRzRp6ZcBfW6FGbbpZRU6cI/Hey2tp1Vc5Fge4tZEgFPwg5Xi4yXxL
VPu6T5+wDJEQUTrKhVvIDbcsea++Lld6aQQRfqKPLs3hTqjavp+ftJvkEDA1u9vZXpnNmh7PqNXu
0yCjlq1nKsiQbmJYuDo6kh3b3pIaXyUb9YYQ6DbzqWnYOxVcl4fGUVrWr5FqgRpGecGraT9wkoQm
TR7mW69llG0f4iUT1WnHvlbA1BvtU224RRKLjjeAZd76kwocBBDevxT2WCbXfIyPCgjw0kvIZ9jh
JpNNYdxFYa3/FlFTex3Yvmt+/e+T7E2N5UAsjA1KnSY6V2rRk0GKEkaxMOG385Yjeo25etqRoNEV
gEyE45be9hTkyZ4w/WmMMK6esGmOrtgUiWOAPYHWN9gpMd28Lcd51Psa2yrM38NkpwrYdWyHB1Cs
zF7/uaVbNMz5eadW8bHuLF2RguCoCtqlzMU6oa6jO+79cuMNrN7ue6UEPsPrC8jSzZcia8CiMwW/
2yPUVdAwU1yx6xkSXHQMh7d/5k6/jq9cRmrXakoo9+/W0z5j1L+9dPAbjIWw5u0QacTic0TURPp8
tUZWgsSu4/XXFN5G2MfzZgqlIQLNzAfHAwNTGmcljPYiyK6IyfenDJasTdkIkbGZG1hQSuhzCYs4
Xt/1tt4BWWbS6fLvvtOVjCXk053E/70qlVV9jAY+wXjc0/WH3ZOABAXgsWBwnxKB//5TMEccgphh
x7kvl+LVbGmwVSMtImoYAzi2N42scdZKkSnimgmJooX1f+WGemkQwI4lcKJ07hxJqO2NgHgYqOL1
VbPcvI3W4YQoxOYcmSLhoQcVyWHIklFpgwcHeGZiLcl2zVjvqHYMzSHVUjXzwUqFW2LDjX3crs6b
9xr/LD9RqgKVjMajoOPKgio1RO7kEI17e4FEnNdJKaS6uHPTW5xtzxGqX1BkZqpgCVrtemipw/vz
mHakHaG8xKaCFUxdM4hVDCNwxowMrQHpszLZeOGI5gBqV8rWBBdNS7s95B3copgNNG2ZMqjHwh6B
5k0GJMKIK1DBooYCjm3js+kqwZSTyzbPN1xp5KC1y9HaKmNyO3GETExB6Yv8epmSIjK28uYNEYDg
5xleQ7Ycnoec46yEK+WcAhmtc0B49gdf1RVKzSeMGuRQzpoekp450h8rWl4Nu22dELkaMmwq+ais
ow7N64FHeorUdFSVadEgIAl3gQJ4TM05PdNucgRy0k1G9sY5nLyK4atU7qWWgeZ4A7YDDZnaicKP
11cZj9sJyVuLXkfBIUNneYP0kUV04lB2D4ygxIKEZD2akGeEC2PUBKqVe+OE9WMVr+Xd92A5bAip
AAw/VGmwjVEF3SFd0UHa+DjMUR+HQEbHVm4ZQdyQJZlwP8uUNJL46eqbDQdJwQWkjqbiVOGjBecv
92qS4VirL8u4RBZiDdgzAajcwsOSKXcsqJAAmaVvz+OxFu4ghmK3NJkZ8CD6AARp/sce2Jm9rFNs
1avQd57bKLwFZ/IgwXSW0vBSBBkJWv4FJEDFm88yOGPDduu245Hw28gR8Jb6nxTmj5s9feuVgstW
asN0OBUpVv1EdKjA05rpdWV72Sl5ya9Tbj29OyDgr5xE57xCHe2H0v6S2mtKv7Ax8Gu/aKqj6yei
MC//8cSvvP41v0NcALSYfxwR1BRzczQg9HwQJAP0iuS4Cuqh+kpXjO4jjiMBgQWWend9Zv4Orvyh
yiKzoB8HGHM5OCuB103ISAoA3TmQv8iRzOKoSDAfQYQj5/lHabpnpO1qHqeF2ZQRoHRbX9WQ1Wbv
ELfnEu2b3QO/s2h9htTBEWRqsqGez1Em1gv3WUX3e7lRQpMy6gvIam5eFIgQ6NOZQekOOiwnlTmS
+9h9X4++FX1kHQ51bVWCka37KzNFgPHRXS336fCBAV1o8YSbR6GXYAjUqoYqPwwod8SWor3kczLu
3mtV85UbVG/xq64lKqJGuGNTUMEzTuwXV/Q6ezQXpl3f0cmd52zpUNcYMI3xqbiHysb4yjP7o1By
c/btciSrcrq//bO8QAHfQ630S7SzWTr26ZS+dDqkLX+Kn44DjXmqYRLKWFsvMDlYM7irlW++w+hc
BIj4l22A7V6VTVQrOqQvioyt69rWI6Fh8Ji8xLA3gWNpIl/wNLlLac0lDeivyqkofv3TJ6SuXfU1
Sybo0VXIFd7/zE63CyY50dBOdvNPpUKwljRbuIR/h8Oat8HMOFpqa4SYOZzwC2Yr/YZTw1jAhwtz
cqRxe8a/2D2MAldTY8XDwUMJEDxBHOvdvES5z92lB4PxaYvKzIzq/BSVw3Eb3LHbXukY5IpSqVVw
VTlw8O2SdIr7KOWH74s9Bobz+berKrGwTxWtf3Kl9/1W91Y/6LEahieazk9rEB3gm+XLsv03tsXh
PyP5pt/7F4OUOWa0p6AKfYCfh/x6LtMVtrvRCr+SpNVQM3MHwdc4J/X0hTBj5a39VWKLgwuHwG6B
YzXBOmpzcKSZJY2B2yYJ56uDoWwtKPeh/vSNUndzQ84W7puSQ4TBaDx2AkONdWKRhEJgXw0noBLn
zoS46cx94XPeB8gQEGt3WdVqlqojCOEJw0zJ56RKYBilV6pOvQD/rDwHVSxJXG/V23oRzCcMB2wQ
782o7wNgCY0njnv6P0juvAmsQ5UtwRpmq+mlSDTwq1QJNcuCKLL8OQ7ZNYIR7njKA05wZRFo3Z6H
1dlEh1TEl8krv6qkQysHaNhqWMSCfs9JKcCJXFgSPC5FqlsOgGua9zM2wGIA7Gh7uJ9GRIDGcdTO
jkp7PPx4bzeWVCqqFycPzXK5H6sgruXUblLXKy6lTYvNbyfkOp3Snws69PeJcpVkKzm8tO8sJfUF
6WUPqVvijj16qPFRv02D1uv7Zz3rhcXEshTYrRdZHBYHXZ8z7F2Th6A6uUGFMxmV5o+x1YqeyiQO
/rHy1KtR3rnC5HGDBmN2pNtwo6HSLmovW4Fq1zuNJXT8CxHyVVgaK7ax7ZNSe1Z7ZQYeonyA4AlB
dCfQ6GgCkKdx7tt2SQkL7bY0OxlxATL0WwYpL9TWdzTNEb+m+nARSLoC2R4U6px9CBXW/iQiBnhj
ZK2+zEc1uf81reE1V68VC1rtbfLtZLlK49J9IbHjGkpNp5anwfjFHWm2yB5fK5YUdfgXs21bZbkq
1xwWC7r4NCO7JTenx3vqkx5HQPAu9fcqCDRdvZQLzYwDB181bI/I0d+0+aYn2g3jePMw052yfuIk
e7BUcDfJFNBjjt0UQTVIiFL8g/KQFtr9Kx6rkfsVbzp58rRchz2dt971Fkt+pBuT9MXi3yzYzQO3
cnFLN5wMFEWk8odjyyBtLM4JFKOBR1IRD1t91C2LqEQroesnQ9X7quPmCu+/YprIGPi9ti2LVj3N
mTiJ3JkW311tFSD54xVHkPzWhnCHX6mIP1Ep+7S28Fur1gFTzncI4r/S17tzZjGAsTltgkhsUb8P
drr8PhcNg59wM01JFvsBJkvlkfxBpwnABvxkJzhJwc9wrdv6pSBXguoj2UvxT5KuUukuwGonbepY
EKYhQzOxLQg2JOyxc3bgXOJZJv7w0KHbdGx6rJBg8k340oj25hiskfF6ACFjiDuTmKqLq+pizRkc
VXzVe2TyXPDJ7MXlNvgGSD1vLe3kw1om6TnWLtrXxWrCud+MnXkVoONr7S5ZS87/vgrd32oFkmCg
RLJY83LZURHaKIva6RWRG7jOhfK4hN0x8i6AhnQdLoT6ft3h96p11n3ZEnhZwlHTLFoeWBN+0qdm
yMSIVVWOIiILZI4DNGCwuKoRoVaq5FFWO/PB9mu6Prcxp1D/NGtzeAW1vm1chB3qpRbplvu2jepL
oaZ0GgCp9bRAcIZ8GUymalmv4rF2J+sy8xly46O0qje0kLqoI60L9Ok2SuCheoaqgNQfj9ti6q5t
uhdStoVbUaeVn9BjcVT4pHqR4FRB1Hv+G6x2b6liudz48TgaZJg+6D8V4gUI21/IcqBF3n8OWKKD
ZDtyuVDyJDZU36DyN2nwnRbaP8O3CWNkm5XRuDxftfsbGH3uaLSz8zjpyTnEhwiyHD0ryYEjhQgP
O1Vs4PyQCSTdiKXeAOJXT6MgcplRk7RwgTtb/aMGrtAP9PInmG3mEeADad+nkApRffdvbpDZLXAg
sLtCyfDai7RxPUCI82v3M9Y3VN8nrT4tdO2y7M9FAx1Zd7VFo29dkP9BIWQnTaiStjTOuwGGFCbK
vB27voflDSqtdYUM5teda7/2g0+qokmJI1CRrFNeqcW8SqVfJYnd6tjTFd6hnbsXWH7z+I9xfx0R
zIubCcnyhDEEFPvUZvj7HTjqGdJSqxyodB6fkAuNTWtwIb5u7xcPF4kAMKnMvWZKnCjwsVimIXRy
tKA+h3UlBX8sEltJzvh0pWpukIbtc0A5csEtb4EssGroQnWnA/CYNGZ02FoUoceMI1n0Ya4JV9AZ
SJcnOh9ItBBN5r/9/H7tuLrc7Sa45JS7cUTEwk8P1JzvN364Jiw/rfgIwkG2zBqJPi4Kx5D0tRYa
RsTvqFhT+ZBe2ZtRpclZQIkEqMdD2WA0LWqx1XJ8yb2w01oEKQOUkKKWQ4q316giOyBr2giE20rS
qtbMivMYHD4s+Pqpw7yh2tEITHrmE0ivTaOVj8I8V4gq977ZxsmTYKeh4O06MIYObPUL5oOpjlYL
w41yCDMmBk/1pSA4aj4hFatlM+k6CutU1dxD2ZZ5RMXm7rxniMRoIvyxtX5Pgm4ASUw2XeeYIHCa
EayJtbxLeM9tIToGjARXhqFnAEXJi4W9Qqiuz0Wt/FoL/RMFwGoLdktOOs9kVlwM60/5/i6fNB/3
6cbW6v8DYl2b0LmaptUXqQmjrnAawtYWeZMfvEhY4+91ISyel1I5q6tLAsGF3KmowAF6A8aCrfTN
EhxkKa2xYtXgWK5iSgbSch+6Rj/zcitc3siqXrCY3JIklK0yRphgfBNlKDXkOEydbSQiQQ3fcc3a
MDiic4/Pqn9Q5Orpyo/TvLVyBdcV09jph2A96DPRQtkDJ4+WjmZUW8mwzcOCa5yNvZFmBUPvHWcn
eMCSmWg9zh3tnNqyg9+1EoNsgekuG7qgQIH6buZ+hBpqHAzVGKS5Xi78HbnR5ubFvR3v5DyPA3qY
dl86VaraFFPrGT6uccE2cYgVoS+yZwAfz8d8GcNQYWy4+RaPpt/VwO8EiXhaJG1oBq43kY8K7klf
H3ZZQYLzXrdjuNCJIkyfbJCp6mE/86L8lQzINiIRVRNxqFzOQu6ng/P2nptEcAq4Ty7LmhL5VWpn
O7EhxHJupmvpSZjzQ5brionWkKNqbZGqle3SAUALQTtXf7guulZacvfkdTCbVq7g+Mpt5BPslJaf
Y/aIeTiZdWuSavXQo6u2zWWNnh8vnuXrnsanS+D0CfguYl0lbcFfmUr6QpTISqb8YIloDMEVfZTP
rnC/6/C4KsnlMpBbOBFms+/AcdiNfBk6cm2BrKNkxa/NpIkOj9YeVOjIifVe8X5ShNfb5t4T7DW7
EBdkrz5TumDRrV4HfCO5YEgg2jqftz+7TdcPlhE9+VyZbjDdmNPRBGdEFPVb5825tzvuJzKmteDm
yaQzKME9J/2ZyMRWIaDWQyqGFapyIWl/24Y3LscrwRwEylgyfuvhx1YdwSpldyDq8WRR0laWMpWk
CN0jW+vMYqwp3RI1SyZykF/ENYLCfyyzDlRzC0nsj+Eq25QsbQwy3kkiBtSRlVO9JNsjV+LDd95e
QSTlLvaTSS9Rykhb6ZFO3YO6nA2cI1+8QwziEakfMkF+Rbbs+nTNbKzhgiIyjQ7fan8SIIjG1W1+
YAPwCkpcl733zUonfK2KYi85q7rsl3LH4/rpnK3cL1aH/tES2NGy5eSeTWeEpPjLC2Bhbao8lOz9
8z3Trmvv6fSmIhwU090zvxneiZePjxDuNjqnnKzfHFLN0xyUjxAivk/AoI3sgq6WcM0HBFVt+rbb
Iykngc01wyBH7kKefxJYKTDwfGDwKdDRv+4daY8VpqLRZzMUxUyZ44A/tpbHtLVhSoQlhDvvQyQm
NO3vF5Zxa4LnwQjT6hpxGpTPjr9T57pXugTXA6zZitLaPENR1Djjy4ppG9RC6xRkWLFwQ+INRn6H
ODNxQf6CDsvRCvYgbxQE0vO2/bcdfe0nqkbqKh3WKLVhUMHe41cL1begfQBMG+wi9vOihFKJtZ7D
VVhFGdnyt4Bft1ac+MoBy/roe6CSgExuoXG+vClQwxsuH3e1xaFHN9Z9o3dIB5L0QBngdyuF62mu
B9AuYe8cVo0ig5pR6M8jyvP1nSODOd4MBe+h6f8MwAeWq7xt6IDOXurAODopYcD66NSdJVJldG2t
ZVICKrv67FfLm6IBlxLQ2ykNqyqEophmrT+LbCwQCp2AjJRLQwifmzABXQ4Y90/2sGgScLTCXC7f
2c2hawUzVPe7DEdmxff7JBehu1DWhKpiRBlUbXh/anFeisQrJmqf+01AZEUgDf1Ecnq8ZYJFL6ky
LqlcBRMPlBsQcws4b4bUkXCK+n1AK2vEAQfqRFOkm5qygynZXJRNEbFhcx3THfMx1Cry3UROQ7QD
/s1KnYF5LlgXdcw9jRtdG8FmnPJbj0EcJ6LF+6E/CVdP9xeGrhJnEubydmA6OZPlVqGi+++puh32
3AvZMsWv/cYVcpDcOmI35nP8Qit4qboofmPnWf7NqVITayEsMfm++ZOASioGoSVabpnlT/rtdH4E
NwxZjS+FQcQgXdw9x/GdYv9uqInpK7wB531ys+Qyx14A8i3AMpGYRSMUSl6Bz+egWw51E19L1Ome
XvOh7hGTfna3BZEU6bF9oJGTyhM411tsL5ifFWkrnk+eaeGMRVRT3g41glthmziCrV6i7KoYYU+0
HwdxyL8O8Dp7m4zqpdW7KYx8GIC3Y2Jx//MBVBqz/SY+wNp8NZBBhSRI+NmsBoX4R58DT+Tngoas
1YGU/bt7fnp0TiPfQAZStbYnmylY8S4bfh+kU0G4XBDvqiNOxKundYXaV0LgSgiFcZR7ZHcAi/au
QDjeHWmY2+2WvgW9ezfm3I8WPy+o0TiWdfuIL9jDGZZT1bXKseadPT2tA34cPr/G2AR4TVD7Azdj
yVu8ZkedqPz2Kcgeyp/QSzx8kkbRzDvq9ecbvTA5bh6OM8sHcQ5MAbB4jUTFBjcwKK0/0pwOcQHb
3WHXulQVyQpBf/CJ207g/dN/TGvRHsv6A7+ShJkxbAoQF0eX5TiDKDKkzpFXk5rgxOM/oFUdO2p3
pfM6o33gMQmshq1amw7bS1TWBhB+b9lbWfqlNjZnp47uOrpFJAEZy1m/rCphvskFgyh3rM7xoQUi
Hbmqfmo0PbRJei15Q+r9t0YmKnvvLyhev5w13MoMHD4ICZtiGd+5B+/jNcK0x9q3EVAb76U5RrQf
IdqIJ90mOa6nD35EC+hyf6iViWwXNWDFxeVBOJv6Zht30r5qQc/CEJG5IhkTevlS9xnt8er+Zg+3
kMg1bm3z7r4xcLD23mzoulhHWSbzXNtlfJ9ixQkB0BuxF4ef2i1b0PZ8LNhz4+9Z111/5M2aZzpY
9ei8exgHLl/+uyLbj0eFDN3QqcZuBGQKn6HCmzOVx7G2KMT+4qb2HQUI7K46WrSSAW8yuIc52jyI
VtcXebqeqbKzY/G3TPCxmMs9L8MTOvyKrfLJRRSA4DlKTGr0t3VvrN3VfFaRdO867Yw9b9YdD61y
r+/EKJ893lQIdvYWvToaXlahXQvtwCSd0BxhQL08fxyodXeg4qorXx5O5trh5S4kHqOC07mUJoqO
UZ8iSPAlcwoqbF56H3Xr9rQwWoa+LZIJHqs8tkvWhu4s1CNXFwhDvidDIqr+GmdNw/PSfEi9YX/2
a0VryZ4Jmmms3MsPrzn6oIPcDjZZ69O26H0rgTZudtvaKAIMrDaBMLlE0J8qDGBCOcmPS2ygbZ15
uKTryusV/5uI+S6jngIWw/B5gsMDkvGhlnQhuyoEg1sSP2vhZJHbTbUUKSozVW2X/UgCEc6WlEih
gb9Hr3O/Q8Lc4HlWNvD1mNE5npWpdYtAEOO+K0awzqssk7WW1oTjfrdQcr3hAR/eeokXzOiUY3mL
pPmhFxD829O+QEDr6j8OGNbFETx8AzAucI95KY1IqoIbUrrbGt0ONHxaMR1paGNh9WJiIDnn0YlL
6hz1Xf1wZnkTfb5oMb4pNqeMf22rWPIuZcTU3lIVJfmYaIIF57rcYq5gemC3YukfZzK/c2+WJE3N
wWflCRMnJw9Ofhl/RarsK6ZkDDYywc5KvOOMf07z2TEK7RYyvMVHeVTlWoMmOnv09TCPmd1CRaGL
P/0QLYGf4EKA7NRWZMJpGULnqgNXXw9Q6+O1u6wIKLvF5rzOGwZjuXtZSrMmyPw4tLysq5Lel7PS
cd4t30IvOyX+K5dbWnOLhSvY0GosZdrVTmQtmqzznIfTbqiYiumrv1zj6DK1cL5m0mS0akaf8JAA
bALJkRua39lrDak+MPSfRKMZbObj4bJwznem5VA4j7L9X6udPdHjP0r7KAtkj11kfZ1dDPsB/GBB
ycZzkZgyrc4GryCWSObQMP+aG+rwELEIb0zE/wZAi26YxiPRfwHDOSB6yCIzr7H/IMJdojjsITbO
HB1km4UW2Natt0ao2wJkC09aChe1wT9cjNfDSKDitKkmgyRy/EUgeKdI1M4C/bkyv4L6zZCkJfay
84kViC8VrlvTQdY/ubrHISPSBh7MwIutTnbadtTu09DUxYBXeqWweDfhQMCjTsjPqcIaiGlh9ttA
bUx7rY9GhRfs6le0OZIZwokrvDI+3UNwwumHs2YzApGFqU+eY2pWUPhKO3NfmEeGNyOOHyNjf8B3
saLv7LbTAj3I7sjqe64xYtLtC1ReOQpezjmu9ogmjaV1NQuz11toqnw/BkzGzVCPTcmtypG3+ib6
If3+o+jfyHp+WewsGEjmJRm9UqGxxnIznzBzXtwFg1ZsMYSA431/FzEthjeoFm+Nnaj2AGAL69G+
bhMF5Jyv/J6d48mhLp8VoldYu4lbDYehPES+VFrpAmv68IetXukoQuFiW0UoS0jp5/sDbKYHIHL6
ERpMCnk+9V3DSwgpV70BEjv2WPuRorVPyNurn1loDG+Ujeeo8GJ6ooUMyKKJh1Pr80NshthKvQ0c
n8ZhmJpPxcb4KJD16W7zRx37F5NTLBrW04opeOLQ4PldAvsR+MJzd3FZ9jMmbf0BESyCSSlEM3p0
Ut2lAU+YRvcqvj9xriUPs+eiPz+2AMZ3bnofgEBn97ia5CoAuBs+o2MyA3dLFDDt7kPeBA6YiIlb
BFrFRBM12qBIktGqyAZqWZ29nAgPirsQ9/UwwFFTFVk0xC9r6M4H1l7ZR7JGZ9OVEKXjjRXDIvYc
aInbS6wiLWdgYY5uPD6yGsOInCbir7Q0ON139jT4yA5FdAORTRXdxX7KraqubzPVfGAHMgHrZ5ql
H/C5VDQGVOLZQAq3rKg6zWOpWRi2pm6ClzOjZSujyHKJKH/9fe/MTVb73GkPKAaJ9e9GPUvQ4Zxo
ic+LWBRglX3QwzioDujwbNVHjVCPtDHNiLVWuB+ow6yfn+TT/6c/rue3Y9i08DFsFKd50diAcuTM
4H7vsZscXVPUEvjWsKcLBn9TK8zML15mp2p2Ze76TDEhpIRI78i83hBGip8oxH+Q8SOw0LgBYms3
ibGwjwc4Mbii0fNxjDB2dps6sX9viNlYt+nALWK2zlMtK1ilT7oGWt84UcfprqfdJ5gXcnC9xJGK
4eTYtD/5DroAfogokxLQgveLeHV49dVNIk+w2z9zbS/aLtus3hKt7i5I8CWcltBd8vEjXWi2Zf9s
mt6yeQIWaY8olWrfgjagki1l7LriJGI8m3Cm34rkiw7nE+MVKzr3rxuViNq8pdT8zWhDA0SymgPJ
3qRt3xBH/KdT+Yyf6vu2apnAb4l89VWDUod0NEuhkdoXv/IcMN9Zr6bm//eMQCjKVG/Plf5Zx9yn
KDeyyKFNkSbbuOalm63fg2IrvZ/o1TVDF8TTJvqYrxRPH2HrZPFhhAZHIng9JHO/2pnqg9Km1BNl
+PqU7+s51x+t685K9erw+bUrr2jW4aFB1jxBJ5+/Z3h6om4Q+l3Ldky4kWHu3s41ovqcTGIAxryW
K+FburSCKz8Z+J7GPuYa4nHGHaT+sloP+r37bVbSCPlOYX3R9XBQTGe5A07mnZwnUqmaLT2QgB1n
ibifS4b8cKHkXUdBlHhlnPP218iteos+v1vb6AFvi5cEmM3APl58LkQ4bMbb9axLgzQgE44a1dSb
hHLTEaFWTXHIfwmGYfurL4eNtFn5KaTjub4rdUGTHsTl49NIwPRylD4j1n4l36aHIR4QWAvK5MmT
W+I8m6ouswWloOKQJybCAsLo7bSyECb9aWPsQ5kZh5SMTgKK0nUkYo7UWBv0LfIUN6mUQWPjG7Li
vaMcaR04ZuHTz+U/v49Lwfx8d17ovieF0RQiWOudQIBIiaKGBsAr32x17NUzUWOLYa66BE2guCLN
treb+PgYkdCTQGjFcsoCHjk5kMP78dbtDP7ff+L1ISRmMCEDKdFNy5zlQ6Xsoh+f3SXveUyVh3Zv
xAQyd2LwniRUOwp7BNjAQtTrv86dxIim5p69dFw0zRYpKPYv4tKqFt5l/8bOu/d3jbTBrZBQl284
zOMtSBpaI0QMUWI3AZuZtspYP1rYBFNzNkohpw0WqH/8VVOSzhY8XPqxUXD4YINlDfsc8wIxwVwF
Iwkm1r37DsZ6m7Jwm7qz6orRRb5dgpzMgLHhnm1TjtHq6uZNk1nFZbYadQrNH7Rl0Fb4p4BFhamk
FOz+o2+G0kbmL5LlhMZAGZ7Xkh3XcBfS6Y9UMq00h7C61qpv7gV+jxY/J7BpyXK+six0pM3HXMJv
58fLQT3hbvh+plJxho6dLYvljzM1CObjITs+m19c9/XFgenAC8hr31crVCKBscyhET11tKaQve0S
0S+suYPg0a8eZ18mT9Xf/0Qr63J4yauRM8ApdqnI9MdSUVlGX9NZuCBsuwanZJfoJZrwAf1dggIv
yHFCeV3Gam0z6OeOaUQgOot2t0CSnNHl1RP5WTKjNWACkGb2u8h3RnUqGk0XctKwDwlS2hzFssGU
SD/F4tJls/Lo1iZD3YUq8tYMvs2B8vCmz2KdstIL+uKZmV7naEXwUorjVg8N60orGh1OCit7P44J
HM6gS6Hu1itt3Zwtkyno1dsXCer61Uspmekfy3YIGYfBoEpdO5hmUuQJeSoelBWjBY1KV7fDuHZX
Sm0GMwv8jdvwfrNFJDRTeSQw2NCSim4/ApRQCOfMEfJdpwQ4dWt0ATCfwMRxrJdy0Yx2YWyBENFe
WtNWEN/WIBx2Z0DiD64qG8u70fejUO4GuW5zjcVMVfNk5Dc8VCqK15JCdc0AhayXj+3okDPEkr4L
kLO+m2Ikvj9mXrXg+rllU/L17HBIfXWr3ME/id4up6XyPWtHcQ43by+I0oYr2aJZnBIevZzd4Bwd
Liab2xP3DD4XNh4Md/f3jjq4yKAYsvPVguLK1JlIRc2Cl4OPvJ4CXsrXxdyB4o8GIcBr1j+e/1P7
zStYNHgomjU+p/EziqSiyj/9WGVONYiLPQzDuuQJ1+IkItkkboaiV0BJxU9TRrTIJzPRGBpMS1es
kVlnnR8inrIl/kh2ib/GvaQfdR4n7LwCgN9Jf+FpTXn3Bbn8S+/V/BLpUvwf5UGm9/cy+Ktj71En
HxEfyKRj/L8+IA0hrXPvd9ZTKak/ZrDNR4nMt4ayKNIWEcdkNU1+KMzILcKeCM/AepV4IHJBkwk9
JhPs1fUNkJd/SUHLibSLqDRzwdo/vV5GtOLR+0a6bXRAM0uSHK/65LA4y4FT8t8+AiAKyJJ16AVL
LxQZ66DHv2kH3U6x1BocdoV0RQ7qkt/7K0dPFG0mk3/860tjP7Ms0ungY64peeCOCzfm2Bz4GTB2
9tDP9LlQoACQvyn8tNQdO5NEy18NdWHbhXt2tFjBevw0oHyenVcqXUuCNcHVXsqY+WdeOh/bXiYM
/QZrOXKNPaP7m15+j2KVE9P1Z4tsYaLvdKJr4KPo7jszXv/Bna9SGGk7e2p0DzZIqYwk7+ortMjy
YMC2lJDLsrCq9F2AhztncnYWJGMyNXDB0wm5xXN9lehHmzrf/tq58RRd4yt+Ho0bk5Y9xR2titNB
jBgmUaanb8W8uqBM+WZGV2uXWVzgaL46WJWJLJSF0mLZBSBAR8JbMPpxg2vICfUYRh0QL66EM9ya
MOA3uyNVq0Pxz1q5uI+m1FQe9hHHP0vJVMx15+nW+AfeSKuqEiwFxusnvhxExnM/CF1u0dOHyb8v
qX6PAMW1FwI2ncUc3rFF3EpxzaF/XJSO028WQL0q07Bfkbvvzx2xKyAzCbkRrB8Pn5ZqSEoUqAK3
PdQPJas8wo80bYw9btu4J7LVSpGph1GT4TP7qszGsLcczNIsq5xuXjphnR5x0ZAnMnbK0/yPycAw
9gB4cQpGb7pV35BUtdK5F8HD0RLp5o1ITH7mP/XoZtv6QgKkcsT1PLvrV9e82yVJYqijlSebiWwq
l/8ZxK4rRrtW68pVisnh6rEMuASJQRqi7XfwKEBES0rhQALY0lSV/mXw+DOYO5etFPJNraUlkd0B
DYZRB4aGi4xMyXGH9AyXj4WyHGWNPrSlLG6ct0E/3r6dpBv+lT1oB7oBLQEvVXjzIcNUwdKDCLnz
iGtgpH+5ngor1AHesLdFescN/PpWCgYY8RiPB6PuxozlUx7tS6GcXGaz4aaLK6GSREsQ2gl8lAF9
32JvPK6Qh/BFkGpzkVfm2jNbT7Ib6Whc7SEllpVefuuChF+Mbx5pUbBEXbJBIexsYkFac6gxCg9a
SzaVxw7IK8aR7TMw6NK39vDyK5M0f5IniActwaAFXy8gloywXVmgjPEj/iULcNbEZhEqEc6Dumnu
hUnftxxz2cKegnT+5TAJov1VifsdDOxEqAwYq0/otCL2mQg9WAIBn0o6JUk1YmaXj9zGum9eDuoq
pLH919eV1+csTiKccyBSiq3Eyo+eecLVtK5nT65T4rb8QKpPmvkMyjJllqRy6XyNMi0MZyQqfo9J
mL2/hR0tieNEyC+6pXI5t/3CzrKVJ98IwEYcPr2sGbudlr94tG1bFEjneA6DkfdIqnyW7vuvNheF
0OQ2LgZu9FM9Q9Q0pkN7Ex//Gu5P2hERfCpbDJ6UgOdGNDVnt+5oc/ua5pV0bQJNGEHtqLMZtOs1
JSq7SR9T/EzS7dYsSJpzFe/ix/+1fI8AKboOEEv1Nr/oxyrlVr8sq63Rt9VlCxwUhLrrYQtDv1e/
sVWxROAzOWsQf8MMi1V6uR8cPVJHhAryZ6sxTkG6FPYpdmxvYzQvGd6mx0vZ1pM78xJ6Zwuvebeq
wSOIz/9ZE9dTrGaK/+LE20J48yBFIiqvG3J1Gsc59nekyr0dkrF1qPaybrwJArgB1I3vpyszqCe1
STJS7kI396BpdzA8nEe5pL+m3CUpYzZuE9kOj7is96Z6ArOYrEnGlAOUBb7mMRsN7UpYaw3UXECD
1YSi1+TC5jZeNL+ozHsJXD42YfogZ6XHewcSDnN6CGE1KvfINMUhXZI//4cFIqGat3NzUyNw4lSs
SVoMlpugAbfGVviXPudG7X/jYey+3s5DYKcFsgrK1rYG0ij7BqnczdB48Nv2GjOH8K92GFfV4Mnc
G+zMSEFIvFOkWdB+29yxj81qZYlBed6RTkYmB3FUj54MPi9KHfZrW6qxLjQog/Uw+wz+WnulRB+O
UhSPTiy4Z34DO/HvrO2iKAaMV2X2kOZOztbNEjmMtRLTikKSwQaGi0ujwJtelYbznK0t/ZMe4ia5
RGgR0aaA7jBNdL1rRUa7gGF9sT87OVGeB1om4ahE/KYztPlGr0lL4Cxx2dbAP7ciHvY7+VTSnie8
4R8BWS0RkqsPY5x6irbwQPdDYjVe4OSHAGBl32dv6l+d6p7IdJLYNg1NUsF3YunSeRxTlEQti5S8
CqxADyQgkDgAlxv1YY8gRnvF4Ztu3nxmqo2Wr9S7Jhrw746qttsweQIy3BDJTBigkmD6DfnHTd6v
W7PkUlkuDbMhZZdKWyWLdvZedUApIrARtPpGIxjU1jc4f2Y11MGn+1/1L3Uk7U0iAJoqNrO9Q5Dh
xskIw6HILhpu++sJAxd17B4rXrgHfqdA3UiTbt3ymdQAl0JZWi0sNUXqu3Tkdb8uT3xqvha0AvM/
3m3b5ZmE2lupHdRDmY6aBIlC3YaLRoLVKIre0AKF+AtD0hE/2+bccG3kghfVKpZSs+7xbOCGWYRB
/9rLJqv+VSKoVim6sd3p3WjvYxcU3sw+9OJaXTHK6RY0p986aGqzrvfAabhx84keX8hKYT+kk5AO
kHQeoIXJbrhtVGIOCaI7mqS3M+h5VeKQwn71uku/QchOg3XI37fNU18OziUJqKIyIUD46FlHfUKA
4U0q5HZw07v0IvzkonWN4DYp1CRKi+281z7bGSSRvimKtEpXieO8uWF34UtVzPAx+S/JM/OWU8g0
hY2rBi3m5WTQX0T0jc1zJZuvFk6U7fVcU5aL2T0T8/HszvTXXbDykPghpn5L8o5LlAQ7hWt9ACRI
5xDfVhcdktyoGBRNa0Xd0uaU5H3mjycbSpVTqDf1LqV7Tra9vGCX7Ao5Yk86hffCkQ5DnKF+9XcQ
FuMS11VD3eFfLIIDAkdjZs/8zotq5W1mguzuInDDUD1ImAarNNHmIeRd8vWozYe7jHX7tV9wYYqg
bMrHCdhS6e/mUyxZfPL3TI8R1Z/8h5W6N8kwxtZJlx8cckJARAeKlw8LVnYV4Ajuvo/QBnNPXnif
lqduXtqhqRamYXKU2oi7LjiSxmFBYUlPD3ggieIidDSA6gM+6uMs3GeEs3v9CGabP4gdeRitMA1c
iFsvw0NvSjQ+8lvhm8XlhcjvNf/kXafMSvYaluHrpaGn3tp2spYeVCK28UtNH39hkqsG99KqFpPX
Gh0tme854VdrCIO2NisV3RfERObx+h4nYqM9z0crkWRU3FpM4hejdek9CI8hIuInG4LB16uZHeEi
CCefKbDqHSUd1xGk9o0dwcYuKThd4aqtNdyC0KNuALop2XJc62gDTCjDdDwqhnL+XExUx1i/Hl9n
8n6iSlm5ExWIdSjPTIsRHxz+k9MYh2dc/sJGJewMy4q9SqVZ5qVoEUZgxE6va+j8zglDF/xAoyHN
cf0QX0jQbSmw3xP2nKc3s8gKsEHkZDTy6rL+Onmb21ccfzRv7YNYXQ8VCx17pG9y/AzwVepK06BK
UHEQSq0v3toJdzJ8wjLnxYGGw7WEFaNp4Y9FhhwAJzF0uRqfsPfRLk/hZ3cfBddR3ZWcYqcWaZKl
zWLK1fLJk79yAMJ2KtRCs2ceAANqZE8GMpcHcwamb7hSMGFt5TwK/rE1PBxp00Xrc7AUGhN/Uy5M
kePJdYB877hUh59owi0xainRxEhgD30GqfWITf2b616TuwdiKVGq0QKVjPxDLpo3YQd29N+8VUf+
IrfYFJCGZCy6ty+CJGA366RKbnrLTgXuUKT8uuC9TDDjMKT2iCEgMDppQW6kqvXykVhw4BQw8np2
ZkgPoU/QM0Abwdl6RStXVhY/1Izqpt+tociy+zgercwpr223Ksq+t7Z82ngm9qni0Gim1SDYvx3x
bMgwPY+2JJZu5Jrkwn2kdbVO4XQzG3DRmL9gIsKubF9LTzKjNdtioYo5N/goJ8zTxaSltIsvxvfx
15fjXd1NOkmSi20VsIfK9zq/Bk4ccgjB1vzkUeUXj/mHq2ZZG8tbT1V5bO1icaf04d1cHfTrPLWh
fehCxliEBx55j3PuC6QOfKa3p4mL+RDsYpFNew9CPRfGiaE0C1ocbIufO6H8nCYhHamSENgHPmd/
1KKr2IcnRFjeUSSy2VlskWuyf+MEvQ5mTCwrNhcbnBYdJRfi2TEwwJVFWUWnFyvMpltkJnEQUS+V
LPQQhB9jsQizjSue6ybrenxtBDXzMZnxTHTJ0knRWg2dPXymUvPefo2U7NOE4bUwXe8BUT//wf8+
A086bFRUrE8ANc/Kgl94PicxmIRvHpUusmh4Lebz6Y6EXmIl7ulA5wx5ZdctcxTR5rqng2mzs/l7
pGMaWC5HKp4m44AXh4QRJdNL15ykHM/SExVFiwPv9zvY0uHS/Y7ZaN0Fonc2KkAbMEwyzzRAhqbp
4925qxTtVtqRGtwaAQ/uUPXzVcJuTdZtkyNcDc47NCgY8PDaK739UCqiUiCHF+sTbO00wlVA9DMv
ecV/UUixgJwjatTKB/xMv1mDkIamoUy4mhkOOVbq6zmtB7ZZtktBo/ChcFxC1lMy1f/lc+tIS0AV
JO+W29X6EyAwCEyFVr8JUDSvwXKVyVjpoRIUYtpmGl/86y7MXoRzUaUF/PvpEyRgcprNv+wOeM3N
Feb/UEiOuOI25UwtI5rIYFTOJ6EYHp7YLCizMQhWR6ZWIY/v6qV5bEn0uwKiBRpb+Pk0zUHf/16H
lQ2hX/ZIthsijBqWu0t95MNgl1ETKE+qsRjJxvqRSaFRSS93MKZ+3gScomgsATSDoqiUGgyT6G4l
e8gCCW7JmYrGlqDKLrgq7P0mrlk7QNi5yS9BrwhEo8AB7NG87wQtIezx0aLYgdSjQjksWp8pe7z+
9CeXtdH+JnolXNJZ6XRndbpZaA6dkbRUGS7ThQUr0vniqXvMeN4Chy9UUJcZ+dsXzTL5PRQJ+5kv
LoGHt5QfXLYXTZNO5HBgWP1i5P2uuTa7tzrYMTTidaK4nSZtWv7+fyXS9NqhOWlxBjI0CvxePxR5
XdFGFC2j8YgRYlDLuaJE9OjLulM+atZcHOeiqxxgivWj+ffQ6OLxLjaloCAtlJAnUk30SGMluRdF
XeP9VQiwz0/CTvPTnvmggWBpBSOm28Y6GqjStsHSSTZHo5JQ+AvtqKVzS4BOcl1VkQ2qbelkxk9/
qAuyTRmAmV+zflWzKPc5hQ+d+1fLQ+jmQpMzBtoodogknUuzIr8jRlIz5ciBj+onF7FAZOUObRy9
54/C/Sb0ZSkMYtIdDBUDGXSTPeC60FgxsiJKlQ9dwFjwd8JqvSgYf586ImmSCsgfgtCG/aGzu7mZ
skCc6vHM+L/C39Hoen4b/XXJVDR2VVjz3+r4Ga1mjeRruDauIbkFAFrDGQgmESYwFWaXIU/58cVx
fJvQCFNHs8WMhliHQ+y+Pgstt6hIJ8uWLiwvTNwAOrDeWnjtx4XCabtT6LAT5L7EqZjA4QyDrJ3w
W1Kix/F4WemjIkDzX0099wrrcSbte/iTGXAOBc4ynbLydPdvYwaKWTZPd0QFPpRAeQnZ2WxK1FUK
o8rbv9WVxDDL7ZGuVNCqZmU7Mz/JueVZL1J+EiuYkaPs8z6eBpQweM4ER8Vt8vtrJ/T/EiZPa1/d
M3RFJwgmRwwwoGhebzP+M/JnE1O9x2ssB1pzvBW7w/1FqAWx4ttiCb5itTaJchkFQGD0+deO6QSc
XeWcr9Lbhmwjns0vGkg6qfSg2BCjwDZ8Qzd2Ujd44mhLI3PV7i4SJBs/+gkHi5AEzukMHDqwJj5k
PGJ4BAM1fbpVn3DOp5mH+lf6QWptyKtO//J3qnanxKAJvWVZev9E4U5taqehThSXrahjg1ANEA3r
mVekbbCl+Q04EvrkebJyH72bH7kISRw1fgQ5ryk3gtWneAxaz82cXjFGNMX2tAmvjuVzYF7neEWt
CAx8AaXTycjfZMB4wYkxsuBCUPb8A8XB7F2/7kj6O8U9UjrNGrhOloXC6QixZ/Ec/8ESwaY2XLfM
HknCitqt588Gi6vaQK6P2cOKVWFokCEeOiZ/SYhCvMfJDeKGHPooE9QpojFV7H8plRdRLBn/HJdT
N8Xir2m3/8xr8RzsJZhG70dDoL5P7tx2ATvsvypeoAwlAXGeCjFfE09WQQV+1djSq9EC3lbWVGhS
ehXzMNIJEirZ+BAmnNtiV+G9q+4XeAEQaWNYNoM4Hk+OHGmXlSToGH4x1CXGVHqJ2iWzsL2JTo1A
nILKiL/mRWbIX92ywMtqERKVEj3Hg5/RJ4gIFSYBsMmRSw8xeGPJRRVE0XSqo5Qe59rCDZ49H7X6
k8sFMyjsvyYLqpCBSaAa1fSwRDRgGDinEnnvL7rbmt5IGlIqV77sK5LAfgVtwtJhy30WtL0/nfpG
EPaT0J18jOwaVDhiSBz6j354j17YWYg6M00IbzgZ8J3tfLtHZH/n95GTihTeNkjVkJIg8Brnjgmt
yGdgiyY0C63lUsLJdzwWeauS3jji5I4gGDluOhbDuriHdxAmYZmNoCc8559n5pCxVJTRvuPfKkPy
mvew/LneaL7LuR7eejiAZrEeKk01EjUhmBoQmCS/fvV/NnRj+f2D50nGdv9Qnoh9b50DK6+xr0wm
99LJ0OTknhnIKk4wpAKJk0BRlZlWyift3Jw0Sc3y91JU5T1ej7us2LdRiKRM01iB4gY5hGW6I+cW
n+IIua8QlHaU9xJOaemFVju4CHEJRU7T04p0qHy8WOvwQRkscdBESckhhyuw5Vv2iTg+SN3dyTFA
vorUve1Zv8ViM4P8TfkqtjCsAfDeguQCxayjHMWZubp4J3mcmxA5UCZIOd5spklkHUu7mJAE6ott
oEcB5JkxQsZPIwCT6F5FI4cNRHPrhMGOzUJySpp1l0S6n/+0RsX//4ZZ1+eDmZT/tBme+Yz5yfqG
C4Qg9tH4DnN4gvKspWaYbzfa/uJj6Opo4g6KCE2aq9ha6uorivUl66yj3xbnFlku7WRYzluPXgyg
Quy/hSdFRe61JBn7aSmiroP3ru00KiF71p+SE7HTMdP2D2C2FxNrOxEcLOH17F+rMuTfTJKtgOVK
SaGkGlVoaEiAPNQtxaFKyEKeRC+OsD4Vm+tpvR01Oei7+gJ5//Q8UFnm6DxGb8ScokACSoCHnC8T
Bm0YvzR4wpWLcyrpUGBlScOfgD3GXbLI7i+GGh8D55JhP0lNxXHiChm0XDVxoo33S7CkshjIfnI6
1EyBNEzEQ2IJvS5twy+sFl1Ox4L5NxOMdLX1OtUI9BVwrKrab6F9VZbxdsjHYBqQsnZibyuO468A
slamo8KIuHdy2j5U46ciWtOHmd19p1leh0jULGHWQ1lOUVk+FU/lQHVYRzUQZP6dSNWwQK6Ek8jg
CL8UTxVqTlBZqpd1y55s48wH8OTibfGSPvMxLO86OdJoQrU01j6b68EfT81GKhpM652mvYd+6An6
IVhlp+2f4xL5FKngjur5tX/h34ouXlOQ5RBPB9OBUf4ir6AcBF8oN0wMNQFJeeNkaQOMAC5RfJ14
WgFNXuuNDxkI4c5RTJSLLJqPLasbJaMfub0sfO/tvup8PIs+NGQMAUiuITsAIPTPzylH1RN3oNMU
Uzp6MB760ohibJ9zKaxFkWffoN8PHp41iFFeL7sBAyxa45LqrDJ7JVfbgW8p/NmdDt7oE2fzVCIM
ypMIwuLUlZhXHQC9v9DJb/KQNxsODnjkVy96EKwQto6yDdUkK+63OxlB+CK2ddXZ8LiUValULdTY
FSlDKv+vzXI0SOfZJHRnVWftmDijh2/8GypsYKbQV7mE6kqqjo22RJL1x65eNd0+BQUtcJHGCG0H
Z9UeKwGpfbTnshPzxJ+/rxPJZjhNZyLG68/dsB4ZIfrzriLxULlfmjmOQZZ+0Ri0HAp1pBN1Bdvx
JxIUIv4BtzOauIG6WoZlwbjFj/+OVtXpj1nQlZbgRVa3NDyzC8qmZnajNnMshm2CjWyAbgOyTnaa
UBP9S1i/n3TGZBuz0+Ex3aLfyL9wWcbywPdJYRiLwYpau+xO8cVr67DeC0RucbxQQkOiXCCTjpyZ
A7ZxeWDK313uTV3q6ND9lu/0z8Unqc0SvX03OpTGg9yVvGElyU/NdhpGmVwSfdTrAAqBNHCOyF+R
xAnkIqYmIoZKR5X3fXRNWA9SdftZ0z+qDGDjlb0rrVjTQr8gX/AT5IjmJxtvbAPxaVdPI2Y0nFaG
Fo+ulZVFKsJGYs+01d3Nz8uwzJh2urYYSL7NQo1AO68MGmjqv82QnRVO9jzUdhDjXSzc7jXdt93C
f6ZrC/ux4IwQytHRdMXBKI+ppKGdjeKZlLXMmploHf8ytWUeeGmKNOxyTPcM49STtlRIzD/Z+eff
LctIbrip4/Y5h8YUR3s/D37PVIiWTnkOK7glzrONP+5DrBiMITAQJem0QFW3tVfgbv30/ZleTfKc
47fhPdSSQ9XylPRtFSRLibFG7rfliYhB+LLLQK5sgYlQQfEyDJJi5DovMa/DQSldVI8JI6s0tMAr
yxLNTXgYuPIxit0IYNdllEj4AYZmKarRo7MjBhRTny8aM5YIjJLCV00SMgmqWjaieGupgqKYHiHa
uQoUYuMHp3Sl1d0JoE6OnvMSpIKztt6WBjMkOVJlFHrjhRsINrCuXwXYDogRX9Q1gRUkNps9A3YG
BmmocH+68jv1e+Ji7R5eiaLpxcW2OL0HqAGEQExf6rYNek7ymITQt/nU8DVxHheZV2Bug4Ubbl1v
p2TzltO6CoT7KFXmgh86vhUY2lnXNJ2Jsovz5F11rGVDfG8jtcCl5d8QLb2KaY6NpRrG32pOHkO/
XPeK2KsgrKLFPhID7E4jUr6ZdMn1IGlUYuH0QBv0S5eYYno6PXrOg4eB8hHMzsUAxb4WjSr+wvUp
4g4g8Cyxoek1hIi4J/Bt6ibu7vtmtrBnudcr8+p9JAz1+RIRrse+jiKyqJa2M2IR78iD28/JCTJ1
rUcCX7H0kBGBTJ6N7t44j2ktSKW5+2L2vMrFRIcdD9UTTA/NmWcprWNkGkQXODgwrQoOi4Xhcbdo
neOkuc1wJUlSbXx3acPq1+qnzrMJ2b6c8DlhOVXHP+jb9zb+J49I/gpxAGvSN8dsSqNuLA3vIODU
daMiRsW53oJ1jpLW0jkJrUNrvtMSYMoJRkaGRh80c3Fh2IqSsyJJ/4vw+1m/A8i2y8YlgdgAgzqJ
Vr8TQXoJAJr4bCDdQUvLYUmr9rfh/J46K0uslULG7GJXdUjbzE4aeuEVM+Hzl5U6PniUpbEFmeQs
f1iNIyyJod/W1PSyYYsOfy1CqPcqZcMGYfNugVJyvwaMVM9/Xum0nt6UNU1eCBerdRQAcFydse9I
H+QTgHLLADEcH1z0wT1Aw8k7/mQBZ1suij1dKzgk0uIsjgmfdquBUTMbwIhO5OvZBJNW4Vc6x2Uj
/l7g0dB7x/+Me+8yh8OB+FodKgf56/VggyljXAfFUIsn7zOMXie0TgB7YJvinL3OPXwtvn2OvHu7
pUcE7hKZE9aF/K/TXQ0ww52d+0hG7zI7vF/i9LLHC35zd6zLV8XhgtdczWFToDoG3oYwVlEDLKpa
3TzJLOzA/6r3Gh1s46mxM2nzBrAyDxyAvQ1RsyvI9x4QqjFAh2+lPAggKnYlzBk/EpwcXEwAafg0
97U41d0bgUjdzy9Ftk75I9/39QiXTsz0DLBFeWdza/NW8t+7QKsEt9IiQcWQr0zTm3u9IUqtOj/I
+JCnlcw6Ig9+Ov8/9MibqTqMdFAQZlzox+x8Jh0JwOvVyKzLkzMugYLxQ4Dmma8TMjP+NqG1Btop
gKyL0aWHminZXtSXqYwmJkqrpURAPe3CaJIWjU3otebgbQoQhWRaqkzAHyjkDlNEApociWQbuBxA
hP0kypntku+iTggrhdaJx1Ue92KUgvXPrdXpNFnuWmojWD0inKAzAiOkxPAyhw3T0rD/LFkgA4gs
8sIt20GIDuz2+N0uEBN0JKizzIa5HEdU7wdLznK11w+2it+FqMje1XidsLxFJJT7miCaYpj6ppcK
WkRwQgJbwqLeJi+swpUYD9tObTcAGFGN6Doh3Bi8+oBGwwQ5JzKMIM33lZy8juQQ/gV8kcILHmHM
gj+vxcZwDBEbuKZ3UwrjGaEAIFCRGGENxwvVLoFluWiDoc8MB1Kfjk6LN6I+yK3uGjziNiocJBEy
lMfVMubWAdX1p2kzlgJjcQMhTzaSbsTwnQtBvlFr9AV86wO37aMxrEPwwzS7IKizzJHoQEeWCjSd
nHYkneBYGhY1RpqDdAUieArHrbnaG3muZvqu7+lOwbBU5qhQaJClO7cv8OnovOvXgJGS6mJ0BQQH
xq1mrV3nLaEOOfIkIa+bkyMMKkZKMT5Xl5cKOHCRxLIz1CTesT9rrerl2e8iTObK5qJK7sT9SPh8
xsIoTsg7AboAi8jUZQt+5fwug52D9456qEZ4Ph7aOFvibhN6yZXCYsbbErqXE5Wy4Z3wt6+NTNu6
Eyn0JXMtARPfSQKaQfSMqTWnXoMDnzr4rbiZ/OhVvnn1gH36lS5lOoTecROBS3SCxJ6vsMGe/YHC
9DqrTrHNEuB18YhHM53imP3YJD2M7PI4dGywfpHRuPtJkcramwOstklNdon8pfMy8zNJffPdH+xl
FAO1C7YFY7A5cEDaQCW6zcr2YEgF5L3I8SJNG4RgVFkCUIt+5wPCJFl+8SU4+EX4SzBsdn9noIYX
dzjtk7CXwbej3yAnC8hcbqfk2dewP0/V2aOHGzFIpS4ZFwBybwgZwAcUFyZpG8/crfJtdWbZ1Ec5
JT4mP7ReV04PzqtuW9hWRrMMfqGptBGUGTgOJv437hJxvbIV0EO4/z+myeBGZTZvGt7xa9NmqHIj
SXR9w6fApNwldLagQqW5NVIG+QS8SwS9vqGCp8hP2OJ/SNPWxNfEVDTRwkCnNAJg1Rdgp0hACKur
cYzvROHvZfQhYLTI11hOZ9KiKEcuZJMC2e/Mu3p+yP4xcspFUWONZ929Ay9RMl5gWnbcDMl0Sh3f
5VzftETxAWUd62/qNOKdc0KfMDD5aXp70gE1lgQX/J4em0ATFO/mCIkkRsGTdIc8xAXGHKRddhbK
u3xMA9V7guNAas3ijVPNXAMXJJI0vd8j3AnEVxRY3tWzp69Z17DUvGoEGnLaXZ+FrIhYxw1MDdBd
9oFumTjyXA53yGGjoeD3unQsKKCrGojGcgBhgIyXuvuky/D90ES1rCR5FY+fIfgvuwqZ+gDVGdQH
JM1hFMTd8zlDfJQlAQkvXkW1BaPL329GbYV15H0rHsN2tg3EI0s1J8hJtUBR+rSt2zzjxRffyL2t
jVBSpRb7VG06UWDXYLWV3NvtCID1rfsaamkx70EziRfboeeq1CHNgRt9qRpUqGC4VmpEFi+E6tla
l1J2ThX+kG/4JiwVc3oXZQSG1WsMKcj8UxTV2axOu7xp4kMz0QT5s5z+uKqQP28Pl8Qw+M+X+uDT
VUVXF5yTMw4rwvAJpcTgqICFD5v9EJ2IdvWPvN8MSSfIADSCEMUymMw5fkJPWzEgxHtxervnmTAA
5rPZifruhAxYuRj/Ppx7hd402Z64KHjnT79WffQVD6OTt7Yb7Ach4z71hCCvl+f2JIMpCnTu1N+u
yQR4R3R224xcXymzZi+BvTvkgq3HqpN645AaDvs8nDL5USVEw9FJotb7cQA6MitSRUDD0yn7sCa9
Upynk9BJMWU714tH5yFO80zv1MyGusfwSM3FfwYLFMyloTckzEY0mFINgEwupcyfQgCenYC76fZv
kIxmQ325P7yZg3/cVrNK6Q/yPVkuFqhVSJAB4zDDGRPA9FuDgBQTNjPDNXe0mNFHIMYXfV+yd8vv
PqI6SiW0D1UZ15mKcnvRgS6ZBsV1isoZ7opfJH6XMtnxFq6D/siXkhCQzfJwGDxqQrG6TCqIdwwY
JMyZRnM2iTS7C5EylkOetPVQH+BtMOeI4XxqzRb65lyqarplkNS2N0JxnwvAU6cwYJnKuP1bVQOX
PF68fhwXgTsi0waOH6OXKFzFlF4hQ7F1BrJsGD6uWlh3TbnLyct7EfZuNURQqMbqT/WlJFS5/xV+
zJy/C7o/uDPdrv/sjNFZdPRI1xo+sLHzqME3e+dpr7SviVwoHT/h99tkQ7Zg5ZTHdhe9PJfaRlMd
4m0aLujyVZUMbiPEtOExaeLaBNrQjIX/8AHuSkGuxFIa/JQV5638ca+MNIs2WcA9ztboRtayMt3S
lvzJVKTYgBOuXFyx+lG2AtwaIIQXqam0gNnJDH2sWSTB01pgaELIochjs9jujLaIE1ZSOmK0vrhN
WuzbUnGkR3Otv4OQA/YFGIQZjTcJoopSRbskbK/U+pAAVloVHLMUlZFcx6M8raU/QSX3gb95ZvDB
syNpRrvqK5e3FTwXJA9Yv63joPrmbuCU7LohvbKWDbbXDQYHlCYS2GWR9A+xio+mMum5uaDPoqZx
bRvPo5gw6da2VMIX9bKkgmPOsqtmOoJFFr/o/Q2NIJjR6Beg1m9/NtDaVP6X8wQDq0ZG7WFpAQW/
EROm1KhCe7I8ZUhbHsGxG53i3r8F9hsjM6TKBNeBsgE7GRc0jt4imn0Oh5P2+8qx5MOfaw52zNkG
foQjSd6011CShOivrqiMvZpCQ7+NkBCf33gcdQHqdcjaj2993OsrZd2nfwe8DvsDI9FZb6Cc9rmr
REBvhPNeSVfMDmE1klBjkRe8+Q2aj86kKqsHVtzd3CMCTO2uz5zfNRtJDwyE4OEtMDhwLaP/7GgC
JvmZyJ1IVwaJkMuwtTg96EBFVJlGbtHfQykN0+AH1kmGyuUA0RyEI6t225E5OMXkd9jQJepD7Bu0
3Z6aW9e+W4FbifPjfSnll46bU1macRSFtLGCUpz1fXemRf60DZE85Di04DGXL+RLaKezzDdz9Nor
bhG1IB+hlq8YaSXWhnZ38yXJf04UYfsoQjtNmrRfkNwltTWylctvdHelzoksQYRoTuIQNacsJB7p
x+7bXxSqiPwOVCWpcCrEveSN+8nz0XPWiKA330jv9nFwIGyUAVK2yGGngqCzUlPx0vWX1Y4KbsCk
h1W2w7zAd/cPjA4W0S8lMBoG4LSBjFf2boSpai8lYhjESwGqWv5v+X+x7H96UKRkYOCrY/KEAgId
hxDY2p9vF/AMbPJlJU8Pwoopwq8Fz3Ob052nqmjm5d1R6Yza1ktR5hD5umn3aVOx2IQ/VpMM5mAL
e+OsfGG8M8i4ITeJpZ2gFZPTkwSY3zGKMUN90t/c8JKvGpWmEp/MSaYECciRvda91gzJpTkKcpc+
Ohvbr/KnY76WcJFHQ/2bVktb1rm5LAUD3eb8r1hbKjIACs+ZChAAnYhq633J3zFRmwQXDBzkNw7O
7NbifBDP3kqc4qpcZUi3a0AEdi2Y535vDXbTFe3agOuKB1JgScU9YEilr7MipzBZH8OyECogPG2k
GR8uzgc3R4tSLScpbdw0vSWQv2BCTaMFXBvynQR/B0WXdlX23La1ST5ETxIcDx+nZAohfOkGq1Tb
VmONuHQlFGQsRG9TpmEh/19AK8l8y0IE+/ZfVe5bCVnVntRU8nrvwXJ/xj3Z1K22Sk+w3O6AVpWW
OjQtEv1OpoLHiWBth7AWDB1SVeBcmemJ3Bhb6dE0q/6oaYf8z2SxZZRnsAGjtlqBhASqxN65dSLX
OrFVcfmpizTdXVQkGAu9WREstEGokTyesXgaejjNTqKROyJsI+q/cwCuaje0Ac2JneBzUg2oJIde
wyQ6nixmQuYldKmiNypnMWU1qD+JTVZ4v9VHE5WQPhVFGie/Y+a1bivQFDYtT+OyIe7sxkca/sQB
P9dla4FzscRgWKsED1pduCKAFWqRAk3gtRWrU2NyrBek26PTMNvmUPEM3nqlA2LiiHXrxC5vEVqH
WyNCkQjeWWn7xLHfOsl26r4824+ZcYFG3kOwdLjJ/YWVsgeLMEDTdkXt9EtXa3dTO4NtVfn+jf0d
bJy3JazaYL3geKD3e7YfRkCJugcsYi54I4y4aSfoZ+n0j9SWUGhv/V/nLOi0xcrLaEzCSGs26cPl
DyjHv87FkeDywwQYykGp4ephkzsE9fZzeXsaRJQjL6BhFpTu0IZv9p9cw0YTd6TMkkZ3Av2Da65O
36mEvnMQXW2AXe+q9qiM56sAM/waGFTSET9eklVDuRIou4Zo+JYb4oscZOGLR/b92rKoX6a50Lrp
ghK/pp2FWiDqgFi2V5piDgi8bkSOGO1ZjfugPoQzytnBqv0RHwqDE71AHEJa5anySu9aOaD5k3Le
GigawrE6MAwpN6Gh+eiarqKy1HwQFPMTG/ACdxKPma9m6eOLsooEzMUlasyD1toKLl9/BzSoJ4tz
VcNa6ZxayHm2coQDXNRCgMPPX2acC8Pg+GrmUTLh0rOF8HG8yhOaAlWf7ZS3RvicQIDO4oPd7BQX
WAZcQIcVe/A0e4LWGVPrUTtk1m4+g1wRehU+ygWoL4wfKVyBO7J71uCO35SOfxKee0R2ksVMUTId
m3KsS0+QSP6ZiuAjS7SIGeUFjKMtEBwRiCW2wVG1Hpr1Q/afTVO0jUnsGbZB4mzDXEXR01/7SpRc
e8FRr/y5MLNsvRpbID54fyx0zBQEQksfWq9qXY1dvAQ4U2k1CdjupFqxY81v7R/6GpZKiFmginD5
ii7b/crrIa32Dvxkou95yItSzxcLy88rY0N1ya1ShwKqcHM3m9VlIhMH7WsMSTkuc2Vn2lTMevHc
B9ESYdNf4t5RvT0PsHqcLzP+TiUvz9zKn0Z5mWfnTrcxPOyZNdGf0OOPxPrhx0QHD7QH9lSae3dd
ixhCzexKj3JdpnpiuEEbM2jRqgc8W6U+9FkZGtcTzZDLEISEE8Gt1QjVF/6hLdWBJML2Kr8TqBCV
E9Odf/7+WAbx//HtbVNubwtIjWN7o67gnBWqKdR6ReI3BVoF2yWyNa5lNt7JqqRi+r3gyPf99MWi
QErLAy/0j0YcIufP7GLmF29aElSGTcPgiF1ca5pgI6oAloUB4WRyJyQVpZQX97liKY20k2g2KtvD
vzbKWHwRv+fHfEOKvhZ7pEDp4yQaRNiYurOADWE1G64maO6Vxj0u+jK+M91gl+msveeW3tum6syp
8QrK8A+jqzkZMZV60nZ0/FIa9S8nxILsmscA4TgK2JdL91SrELm2RfctHGYADiM4i21lWrx61mFX
llVPY0asgTivJFCDtmjrBDL1ruK/ZQU8DCiITTMYQ4L3CUcmtXfLES89vuXkyi1u3x4RAXJKwKn2
ICPWaInVeM6CjcEQz7fLCv0wGmld27U777W8jUCvLNYJ8Wy1Nw8C+zEMOL5l0f4p9ileeekunH8M
h2isDCZhjgHzWwRWZToz8dqmPetR3AAJQjKf+X4yyq2BPLXRfQaLmbB1AnOc3Au+5hXwigRlUl7Q
47/XB0X3lFpZsKl2R1PL+RrMKfXbWhQi3UJlC9ozU2Tl55sbpQlNdnHNdA2Tt0ppI+Ec9Xkbgsjw
iramAZJTL4YHErvlQ7ms/zC8VDLQcMOQuPWiOOTl5fpnt9nKqMd9DlbWQ+9wsf29UppKnVjZ/1of
z3BS4GC0xskLPz0LAJovpl2bu04iJqTDiy1Ee4w6bycjFi5nCTo2o2Ai7qaSiqsXVgs/YOQkkMPB
4BEPPnlfs3PLbulCLAuRvOzxHltKWrkK56Wh32UhsveGnwvDdV92bRhp5FMleHC0+UzZx6qtHQRG
aKBcyTxOtNqCI0TiCT/WbdOz/GlXa+hhTcRw+cjaZfbpAkL1iCW+rYEYonWeFDeTo+lEULjFMxhI
XohU9dlVXLWJ+nW9oJ4vtRgBkIELkrmqN9KIf5/t5sOLljg4rLzTCdvjL6BSJHiCf6Z42wgZEsAP
NbYcRlNv4mczKCJSQYqNR6LTIe42JbV3nbzMNp5eRCCGFdSsI3JIO8M2208/fgc5ATPi/XtgEh3t
iWiPC+0SVRNohpGrsn+R0NwFH/p7Vd34ySBTVT+u5vGrOAlGyol6ybD+hz80mtNvcDBO4cHP4pgS
i//83J97NQf3d/Vb0FZodVNly/FZ3xnF0XgEXaxxNniRT+E5p81h70FyBJUYksDwwxWD3Er4gB/P
3USxYB/ekTLjAN6uNFfBSuBwwWaQCfE0MW8sn+WgnGNYNE0/q+PpMGSI/bY2F39qBf3BihYkhmdH
alwKzq8rP4GP32pAqNZevxKUNlfB/jR3OElukJ+TkjXcHSBr/ZL0tZE7npHgqxUrdpA5wluCJMYu
kSIJv4EB0Q88tJbmTj6Hpcy1l2apg84yorh8yX1YaCT1wQct5CRcLY9vJcX3m/fX4qTsi/07cX0E
1W26vF8UIb0Gk6pfns/qLqyXNivNUrBftHbY4xKZ0s2bQjfNJUgvmXSj7faVq3+kBO5o+hBg3PsV
/TFWyxn5jnmDbVkBdEkRbPCkWsou06boqxYRctM25WAUCSweZSGNSLAcQ0LTb0ZXWXUJ9E4418dJ
GzorMyeLre7bW2tQUMeJXDFogG7U3nhoGDEGSt6zSu30stkggjxrFZMnzYLXuXJ7zOXUl+s593jB
4rZWXbNUFalEG8Qa/voijTT9fzpNGdH7FdKK3IOTZDfTVe5QkCYQKJhB3Wd1feo0P8z6EDmwyMMA
6wkIyOvmz37av/TLbIolzARbdbZOdr3eDj8zgo46oXZKM7xvV2f4HmfS+alNDYJZwmN0RkyprCJi
YOSFqBu62kpjYSzh3kseKzxjPJlsttdd2czWvtwpVzZRzIRF1xwanasLMUWgpxg4nofca90YZeZN
IxG5S8b6OAOcO5U5CbHucFgKsZ4Cm2jRpRNs4/h3+x4IY5AIG5/0HGr99AhUnb9+3/pFsFKU82r/
DC5I+Y+PjLOM01Ohl/Zqku430ZL2w5xxuUEFWUazYO9RciUrEiwhYVKscys0HcA1WF88pLzN2zNs
kyx6soW5M+8KiXQ9XHbk8tnGNEbEkoZhGdT7zN3dLCtUhAwmcHxAGPkU2/AiYKqywGBe3YcbRUgN
PYcgLILxXbi0EYe/HisagP4ZwzNeJK9QmomIAsC3S+CYfOerYWt+CHDOJ2buf+pxbht5KfzTrxB3
+0AgW0BjH78oCojPB51NkakSZ29WM1rmqlQfD5Y9s1/y0tE7nFKI54zQje/NZcBu3U32ttCh/VdI
FlTFuqsoTn5qiETQD3mCmW92G2zeC0MlQSLkgcLnFt031rWyYtpX6wp6z//OORHZIHTRtD7JGCdd
8dlpfOB3mgMqn+cf8CNnPE54aUB3CCqBi3wFYxAJvh9fKAnUd6krcSW4JZEEGua6/jCaunDqkxuV
tCa6zeMvrtt0/xuRsY9lpb4eIkS+SnPU4tt4U4KGA9IvUfYYewbw+Mek9+d4jpSSfrXdFCZ++MKo
ry+7wm277lt/WZwmkPCr1bdMAfg5aeLYYBRkOSlHHehbsr2+yUNtSms7zRJMn5Sn0tt4ILlbhpkE
yJ0L+OpKIDxgPFp6lDa9tkKIRTO0Po+PnXWLhXKxo0Sn8i4nYMEJbmPtxw3WlNVh1cOKyqNb4Yyw
lsf4Fc2DAO9TCN0lXsqZta6pCWFrYEfOn6T7/ddGUe8/yET9dXY0RNvGPtbwZixOjM0oIArIFBHJ
ZPid8u+2cGejJspNC0nD5hKiC3CfbRgZHj7862BNFJdd0nwB/1CbwBDNH7g9O45j/CI1GzzUvuYF
3M11rwmkRvVUSAn/d2DEN3qsmTfg8iAzECCfLocoTL9lJMEIJo5XtRKmB5QgrGiH3njFXw5/c4wI
DXMBgwGKNN6kopo6kSsHlRm2SJzIOXlmCygew82qdSAfyQAFC48i0nx8e2IvjNXkAMr4qMta956G
WEh7wfSoDQh0TQK7LTuVH5rRXuX2Mdz/6C8RzBGd/N6nhnEamyFvkbHR4D57rByCe4SAtnr+Tf+x
0uhzhGpZziIumpvpCerQVeU5/pZWUM6StFiJFeJZiayThYd/Wek74w0vwAVAIphoXvtrK//2HQRm
4wjqXSx+ByOP3enm8mEg4CbVEeFqSzF+TUFLPi2D+GMw6vbYDhi7FIlvAltHju9l9Qzz2tS9yTJ8
HVsigkQAggEfl9WQ/FwVuChQ1sABktQLWEdJe+SDB5pGidVC3ALEHUSIB35h9hAsNbRAd7BFupVf
NAppAnLUCXKmPghQpu0b3X6edGoS4niljn8rlqrkqBlKEOhGHqVy+RiqxdsTapATvpf1nQhsWc8g
gNOu6bo+wBqPfSAo0sHWHS/SWqFyNP4oktgLqxTT1vwCWBj9y9Hri48IDOw86so0Nps5GpBQtBuF
8eWiYtj2CaYYmHNUQgpXLGPTdM5hSqqewBWo1h8AcOBy2AR2UM/LlvE8wYnXqumEi/lWnvt9rXEK
rqCEgtTcY29fmYZ5zDin0LA/VO2YiSIIh5ajx5hXD9/zLvYj/9LF53J2SBZ9hzRosvbMps3fYSfE
F63h2IGcBSmNPNkA3VAXnRvqu2DRBcLf+3NsN1XjHML/qMpMIgMTTm74NTm1PFppW+348xM2U5FD
Dvo9omez8yJUVdAi/k946e0BABd1SpdhKraIuF3W/PN1gKKXMyMV/EZej8FCzQ5Pqzwy3J6kRCn8
UE6HOrYJLMbV6aoP+/GEOMUeRsZh3OH4paoJwR4mYMKoiKPqV4H8aZJujoFpIBAgj74pZVpVr2+P
eFcLXVOI6/rcvMOHORaJat/sCDyooGHmKxI10tcEiWjHuuGnkJEry/QsquXHAjxUw1t91jKzR/Xr
kLXyiwatUcdAZ6RzrE12bAZWcPMiDMpiKUGf6pzb5SmpLJh5dIMALX++WT3Z/zzmGWz9yRvWej9b
Cj9SVcM8JWDytAFd29LThmkU6RhZra6yZg5l39vSBk3j9J+ykl/Bq2+WmZWtWb2udN6gffzdW8ie
pUfqpjF6E/rqjAK/r2tBjlpnzyTSDjIfL7iI1EDs/QcQ8Kvb5CnUPTuCcjy8hCVMB++9LgSgnTy4
I0QomeKmQKgz84ADzY6E4hZnDJx9E3P/t7ZocVHzcuLlNZt8z8epGLLuXtD9jX4AzsnkYWSuoQwW
vtK0UBFc8Ek/xkKBBXJTEoTtgP2bdmesRtoV/+Psg8yiuyyRJ2Hs2by1qjWCzVVAKXJVC0jRTiVU
6f2giKb94Gs9G22cV+dEZ+wSTgF3IpEwmWgkXT9dtTwzrcmvSpaG/Fh4Y3GEt5ZdaAxA35F52MeU
yjF/NfgfT0vo8E3XCSi0KYcsAAiOHnLdE7hLfdfOil0VmKCrh4ob0U6xv1yoawRfigeTI0Ksidv5
UNagyX0GRfudobd9yc+DLurkWdbxkYmxCzP+WzZlqE0uU301WRMHFdrc0ZzL7LGaN3sdEwgDZVXf
oBHpp0QBrl4vH0lYcj/UnUB4WA0kzhwJimALKNNl4OJUi5v0+A7KTnZUqUSTZ5YcTynSE/fM9cBq
7XujEJ47l9WZQldpjuKaevX+o4m2ffV9IFZ0lzxDBnquRnvVts6qGo7YxQB/YPl50J9FC0ebq8qf
NbetGU/NaosodvzkkYhPqBui+ztYM3pBupbwrEesUnFa5mG0gunvH0DIz3QoBDAsZGefzrjcoHwf
VueTH0iitQVA0UiMlbzDwf30dXAwusF+zr0Vkgl7Z+K501zOwyn+gzwv5fdyQ4p7/4dcJsHLAcbt
ScRJRk3Ziy8bHkJVaeViiMqDRVfDj9LlN1bGqwGzO3M5633HS3sfP8GCo8+Ljofqf79auFp0Yzxx
+a9AOXBGUtCaW/w0dfpNgLBDgo8DomCiF9SfIOgR+bgxWW+DGP7cK6dAC2LlCMbOHJNXds9fUdnZ
mmXqlvkolzufAoJggvGh3cW06os3jCPOE8lLDiWWDZTq9ONjBpyqDYTgIsCN9kfkOj1SyT6uN/os
eYuOi171Fe3EkoKNH2/wR0P6C0wkidl3m6tpygfKjtXx93jHj/FCjqbAIZz2iqFFDTVKrYMYfd0Q
jieI62SM0Rx0LRglqWYef/QFKdky2/AIP7TDSUz8tQiq8doHn/GBIg/H1yOY137YsLF8VB4g5cAL
VwIvGnl3oTGoL1EZ4cqhQxWPeu4CJ0MSfEKknlG07ZoScnCLKLnpRRrl02aOReHunNaySIUq8tPQ
hvKWa7UlNeN6H/ZGayXEoNu0j95J7SYDLZOhgFstd3PTz+FioifEPJjMEjydi1GjJhndyTIKizyc
te2kv5WR8xnytogvMac9cIbaVPo/E+LSJpKyh6W0C35E2fhx+dUaCPhON2P1KcYobPELRBF1aPsB
yt+KRI3Ypr+Tn4QnP7MJvFhpxLWJzwpumaqs2+i3wVT5XO/Mb5VGd4ehtpB+EPLQ4vXBiC3aWmOi
G4JN4+Ng+1pGl7gv5LILLjTzq68gmHGlCap2+QSgEuZasyATPkcKJ65ac1oApW8BFM/ktHE+gdbR
Nxj9pw/Bbh4tDLsCEpJAlIU1uwg60lBgiDjyhkHldJU4QZNgEh7xk8aH40Ns3+4LODHyDXO9PK//
W5YkHQP40pecV6pKmfRWtJwuRIxSPbKz7C0Zj4gSMmaHSKYeHOtqKTJLQFaYZJ8p74xqYw/O0Q8y
cpHFnVh7um5ziyBsW7gz5dYBiVIcf4K63mb6WdicdEBktJdZFnwMRnxYMRi8JkUCjex+OId6zpH6
dYPcdcwddaO6CVmROll6hGvk2p50Cn2JDXx9vZFSVIgoxsIrZ7AByGS4HhZGKnUVPgs1PxsMqeVB
d5KG6l45sPHRonle5Rd1SBhUxu3d5m/PxyNyuhwgx3Hm8XjXTw6niGCnaJ2JQ2b5rU87JEJI5PML
3rzYk6A4aV0V2nYe2SKM7RLQoeCXJpFqOIHKUMiexQDeQ/LgV9K3WGLPJvJjxKTn8izcSWYJr+zs
n/bzLHENvNWUGz3FIez27kzeNCJ7/Zkrq9+WIyLFkEDHbBUNhWFMRuMCxIrL7KCdGT638PVSw9QC
x2QCobdhzqLCgIkhltfvoptyC4Q+uh6YpF5UgwFdnIBTrPvjdYY2esYNcL/v9vvT92aLTJkjF6wf
ULJeJ1Bj6lpuuI13rTVf6IvDXQ1EOYlStzIjaTvM/gOTRxu6RnKO6Z452REKKMNeVkpxz8wuHvGn
vTKqvcfI4Kl3Gg2YO5mk3jwsguFLksRFq4Jc6glDiCNu+FYFn0mTFnfLjlFeamDf9S3Y4PjDCYBO
6u3OAHGQe4XJh95xMMYcVDXQaXHd6ZBwtiKrZ01sfF6H8vDM94bcW3mH1YvmMDEmgPxAB5nCZtwG
FEnxZoioGOQJl8SaH+HT9f2/XMVXcPw/4q/GAeE5vuntXs+Y4a+dyIi8fVrJ4UF0iA8h40OlhP0R
XWkjmWvqpvAic2okTdp7yK7fdyP+gSAt+7NpR33lFT6WImQeGgQ3gK5UpiSSjj+IHV/1UozO+4V/
DLb9qpNR7hrnBW89u/Cyhimli8aT0SpZd/8YkX1dAv0y1qKfP6onz450p0QEXcTjC2Cv9Bydjhd6
Qw+oX/ppOoBCBathCtFHi0OXvPv3Coi2rPfa32NCltgAOYwSVACkg7FVmluEduhpj86SUwEkhY/I
KjcRZEMnPO/B4MK2WYO5MXxZadFaHjcXgygAItvkwYNtqD5qOew49oosad+aHt9wnhUOuYuuQAts
pr8wP/EwG8pdxS+LEPTeQybOtDF2nzYD1lH8MWsgZTfOIMOgfbfkZ6cmVBcdJtz13eKbTicAGLcd
frLBMa3vXx+SOByIsKaF5EXwPz52JtVO2VekkIAdinFuvdvmHC7Pq39gRevkb7WAQde8aDjRMcv+
y0PC62KU6i1QEIPqRjpe1BIj+ZjEkCNVfX4uWq1mkJgm/ZA8QgYtCPgFyxrbukm/SOhamUc0TmTY
SPN7Oc1AlbYGpSEQlrJ6lh/9fOly70+1fIXbHZgOjV5dj+SKhTg9jphXjZnZa+wafNGE9QzU40yv
R5vRBFZNrfq8U78fHlaSie00ousboce19yeQC+zsF3QqHwmG7e3Br2E60ZR4fZUPFdcVTo9Nxzra
grE31iYAgERyJoViD1LgmaX9JuUkUd7NQFtgdJHrhuCUxxRv07/LMN0bxj64P+G3syFruMG4cmBP
VbLDaVrggZg7lF7ezghOJhU1rUhxaeWeDpezl0JYzg/QZCJcuL32/E9QLNAzkp+qcA0xu4I/PsDI
4HCA38QW+4jMmwODt5kRIw/fNG/vvspWLpsYXdAVJNBsb2QRLyaSRYgtAc9/97SeeuBkT4gHS0pz
gfvSBoBeRHNhn6Tsw5Q+6bJ8zSqXEbm2mxfIdhIRqQ7jkUSQdhqcs1kqlZvRybA5qytZaYU1LuEO
Z9usAHl7bPnIzxHaajOn5wzjm6IRnzaWnxAlVeT0AniQ3FcygaJTHl1ZJOWXo7YtiGl0SAviQs9Y
RwGnQSDPQf+Zyb+XjKd2IO0sckrewlStzdp4LP2lhw8+w98bYqOSw93UGXq580Y+LLH8zL0AVtsx
xDP7ouD8dBGAtJPqqpsdtMdRPqGLPLNV1KYSoktTY5MGoo769DCfcNcAIEKryQbOOKzDxipuLzUV
WJ/AJcM05q4/yFMA+Fcs3q1zww3DhpwucX3E9pMSBVL3xGi3kqFEfh7qECbrYFktjzimebjFgvFs
Ba5ee25nwWSPB8qAtgNZoEidU3ore4BET4KWdbWI4gEeJhuS0R67PtqOi9uflj/Mtwzu9TXWYIuR
1f1nPAkmoi9Tdb9Jheb4GN8YcvbLTY5HqyTBuMkoyeJ8CsS+VZNARYSVsCGzEn0pydcXSN+8//2N
tY7gU/NzG01XH+3AiYIrA4LXmSxEE8mH42dbfHwfm9GTXriT57w5MKzqC0epjWtNlAOrOOvJEctI
fNZM2Ymu0Jx2Ig5l2tREKF53xoHYsmrHK5YcVHEwCzi03S5s9O61/t74Ny0mda/+EL7ZxXHUOKaI
HKD5gADcrJmcoddLmkoPCqbOvF+D34Cwy/QnB4Ln4Z+0NxmnQd0Si1w0xJHmSiHEPW/sIyux4Xpq
EZVksteoQ46+vklGlYFMDv6IoS7LVBqtIr6WPG2HFglHGg31TBwuI6zIvz1rQz65Y5EzyaoXu9AE
81EwZ6Fo58F9VyXeSZTi1YZx6XI1aC+xmjzieJn3I2tDYBV7M20ABe8MzLH3Hpzc+gtLMe6PFu6p
e7aoKisY5KAVB4u4BuNUXtFHGGC2+n2SF9Gofy9EqW8y/w8Lg3eq4NufoHq3VjtH1n0RR43CTBIB
6pIo3YGfmyhZ/STNapzfpIuGnDO6fSn3izlR0ynN2XF61I8wXsn2x+v15ch6d+0UZTZxfQpmXBr9
6KE/xgUUVdNgq45a7pZmOA+3ATCX7Fed72HGLasEezjOMOu27EwX2g3RMgqVQmUhPAhkN87tyg9E
KhYZSaueOqj3E5R85IsYQmpWR9qsPqoD0lL13GQbUv0yOX1/De0kv25vv3Dp1aROjeMfswVlTfvz
0g9zTfWVdW0X17HDuggYlWKenTQaM0PRXWlNZGXYrz0fDFAXuz5W0425UeqsvWPC3Jm77y8K7aEJ
CNACg3S/5xebEU/EAvWazHzbJ24AJAD0YPpS03neT+3keUrjM1RzTJNpsvmcZdZMowosScQ0Y/aB
N+3J7TI5DdrCXz9kWHLCsx2EpEIj/cC4mKtW754gFsap2OyhQKACD2eVRUSG62GnnPK077lndhI9
ofo7ZEAwMnU3aacLoU56QPPpqHFJy/GjGQmCOZzY3+HQZ+GO9YWJzgF1S8hnHXD+0s28NqE65mxh
IIu9EfH5meaXeiUSiyi+EESHqsAs7iVl3Y/vLECLAbJTuC1oI9r56x+oTy5t8EQDqQigHb+wbHR6
+xV0+Ztgs5eWOh3LGaSVzOJo8UxEi7zA1BiUMTe/B6ZQTBae5z2Oi9Lf7mce0xmHwY7mICtrVP/H
jjtjl3NR0mubJVfdaN19raBZmWgtkJaaHY/yMjVqLU5djmf7aGawrkp+wl7wpghCycC7YSkf0ejr
bjQE+mMT3l1SOgbzeNC/tKpXKisOzeVkLWzfzelYq4laNDuiWIkQVj9kmRBVFrPg9Bi+kV0nif+F
TtJdlLecZD1N3SSHZ4m5ICkt1Vux/b2mBSs/NMa137qUSgctOZfFROufimuh8Y8KrsKoDSZJyIoE
PMsGcwyeVZ87aGx4JbElEs9ZNPBTOWUPgExHQ74Dekaj5xZMBTvKGqRsQckNy5IF4VRs+Axi4c/R
P8auqHGKc0+Uysd7akhG/SZG4TpcJUL81LvLC8IJNYHcgqtY/OrCWsG9xie+K7YT9g37PfxOTFCW
heONC8Pbv4As6ZtkjkVPHDVuQfAtVdMWH/0RmnH7Cr9E9bKxGNtlvKQMV2zVOtVRvC0Rf0FHfjon
h4aEaLOSBrZtFZKE0qSpErjqX+NIcRa1XFvjzy78yMKUf6YnbO2bIkLvqfJo1ruK9RKVnUz/3Exj
KQ7935ga5uRCGQzauOCJPxUNwYGag/Ca74pA2Tgd0XH9QFd5AGQ+Yzq9uyNIhEshDRUujRmMamjb
4FnUDR8kX7ckdNOR5gePeEuzbZK1fEPzWL+CetJlctSfmxBQvVLLHLSB+34Mkz45Yuk6Y2bCZZpG
RUzSekK5AUEg2Y92y1qPY02Yeg1OmylD4I7pi3Hb3P0jHZVkjLcOX8FLLOvmAVtTtPrY+pK5sDQK
fnTLdPzD+ycV6mzuYRQN7Xshu/mZNvM5gLWU0UrBl1aedcY+yFPNgoh0GMDf2BRktcL3pmei1L+R
tjG+sG+fj1nKLpZiRJx7ysmIZm0+knZ+NeWdc7aTxtY0kT0iec5Tsiel7f5iFpywK2/c3QqPW8LA
huNh6eBd6e7MPTyEXZpQDGFj77qav+ej8a0mwZynN2gvrSCNKI8kWp5/GWZpVBlEdBBXH8dDpVz5
/C92Z5GbCdJv8bu1ryvEfPFIQQ42YGZu3tk1c6KRBQTxlk6ENZet3HKW9LZ/MejsgZwSI7TqMkOM
ikBuYD3biGofOInQFhCV5i0agc/vI3/Lb6pTyhfof4qFhxuStIMnuZD8Qh2lXAMmbw27vbSxrddv
cjTC6aEdRZkYslGdFJIbYQ04q/JgYm/movqAVLjQz1SmLmajXCJbht4Y8YDfVLIjfOJebWOCt8bk
5DsLg7bkITfCn1XxrwqzmDuO6WqH8wOprEEcPZQcObISLa+NbMDyGyQfrJCIGuwE09RGR+K4Dnxm
dTx9srmhsRC7wIJCbLXS4ktjIVra1xvoDsAvzM06KrpaCLEcdl9PphXxftdoRh32hUWlCf6mZPCB
FoR89btL1DCzaIcQr6iQM2ukagrUPKAaZEEJUUBydrBSWzM7zf8xTZZGhRRzRXpwi1nSC3url/iW
t0Wnxcbs36IMbZkiHeVRt9hbgtdXFKg1yvFs/+1czDj2gV3qjhvL5ak33UXXBQ276fET5h9OyZQT
VCuQvOlnP8PBOIgH42WCm6B0nHECb3qmfjAj1ZzTx3aXrvHFy3X835PeHU7zXZHNshvjOi3d/H9o
84pSBvYovrCiLnpMBhpAXMqQ/+glZq+bjWWhsVf2MCBgQWgXZMqiFYmKMNm+Zkfu/NproTzzWXUB
glnffpFMfeMpkcHTWcAK6hB7jkHxUrOUuDDh7MMqt/ji27Dff13qsF1eYEpduuyAHHEbhGQI6wyu
vcLJn4BJLPOYsKarKBJmWcUNPaJNElr7hXCXOuufpNFaHOHVlI0ePR/qTP2NyZrwiM3bqDCnx0hB
Q8FQcOB06xH4zWH3JF4Nl2zn5zq2hUQdSN0ID4XMxRryLDkuy70X71uZFLKMEtkwMLuH019fIYcQ
D226T2OscUew1xozkmac5uM7+MygyK0Vo1Msz0Bprbd/4HKfAyQ8WY0f9+QuPmwxrhvv5k9FZlgA
UF72JQDimE3dpxWjH4oJ4jPNWHJu49+fjk0Or4JjS5q/SeB30LHhpVjaXd3A0yslshElTPuyXt1T
/bt6Sccfa5CAbUBFdPbaU9z/KON/5oRxl4eYAnQIrtAquk6ydbfsF44nYnRXoDnOu8fZfBKqXGZW
O6w53cTyGuJYoXE93nn+chlxeAIf2tPnG6LcqEm0w9ji/aHFo9s45y7JTcQWRn7utvtbfg9edtyi
Kj14ydUdUtPp8gkUF7Ba9kgUKAdPwnOu40mt4QX7RTS9PCZY8L7N8t0A4by4w1u0XjGRjTcEmfLn
GrJrbN7Wt5TsaLZeti/0HycYOkFF3dI+G/b7/DFsoA3WwaZ8mBKna4bs2uGfi1xzvx4V6qsadP/k
ttyu0PjTui/LzBLkFkDH3389BpvAZZ0yvNOvz/48hOwHbSCxetvLy8rYdwv4+ciG9nC/ckNowG3W
SCGZe3Z7eh4KxBgYGkkpNPmuy/QBocqiQ+z8/Jn7biWFJ8nSzmz5xvY0p74rGDURntkspo7NnbSN
KJ2HknmjbEoPa90gfsj7ULhO2j6XxPRLs7DJoZIx9jHDji9ze4b6FE8Mi3iI52WIjmR0BzxJeieb
igTQFBzjhmk4qMl/otGKOVdPv+q68nGk+FCwD4ZGubf3yeENmn+7bShewD7smYRraQBZLvmhtJLb
FQ1N1qrKn6wjs4+BkxdPsejdhArMRhoH56sfr4IZBaaSRV1O1zhzy0EQhxqVp0Ws5cR1/MzWpb4y
TrrMTAKjVy6/vZd7QNHYKF+V10iguPdrRkz9BVVvzacmEuZYI1PWjdoCz4ULHQ0uvYwIkpLySmbA
+6fpJSaB8CdsW0EGM9yhIQo4nSkafs4q0AXHQnbCl8+u5f458Ecc7ud5BnEGeebr5Fu25J164q21
1GLTwgBb0d9Sc86yzxNXhRPFHmQPwj9kY7EczVo2GyhCFAQVeAjowQX+mhNe3TtcstGNCA6DyqqH
wHE6Hvd0FJV/azo1FE4LGOF3Hy5S2CllpZd0vMKKfF6YhIWcfApLneohNZm0nO6iJpy3yi/7xy6I
TPW/TiheQ1wWxfPK601N/xPfhwVKW50M+aNwKZw9AiQWVAva90S53XfWV7Cq27pIYBQh2Lr+BuVf
D//AWTxC+7IrKtQgqFoT4Pf1+zoxhMjihyc3pA5DYh/JO60p+DOpgU2rpXM1OPJLtBarzMlgcmeE
oEYdoazOJsk2CZwXZ+uCG361N3m3/1gOfeaWCd7W2o79az71gXOsvMtuRlsxwuJ05Gwr3kvwN1H+
xjyyGYsPR0Ik8SbBXWx6ncEJ4QTDL4YSVtTCG1iQ5m1K/fPIA9DvEfVKPyUJTV5MlUJxvHCCL7G4
o61OLRBBg82KNs+VRFxce0Qc5zKGbIyZ67W9LuB7EQEsfdt7e01ZrUVg3jM4dSzooaZmuSQ/kDYE
mTryiZ0if2E1qmraWl2Rw2wU/BPl0zUIz+Ik4aE8UiRZP+BgYQiQzdM2drUdfII4hwOJ6UPT2RJj
U51ucKoe1RUHTA5FUSQiXjCK4LsWld6g1EE/qXCUPyPvYMWuB3tnFhgJT33cAotrf8Trnnm28xNO
gDNcxbRlFmyM/e8Yey+vxess+ZTKAI+7OsC2UYE5JAZFvgdWbaz76V5CDoVmqVS/zbBWoyV9emXu
5dLmDPSyLv09Jxf1kIez9Pcf5h8qX4avHKL6QLL81jI0DF7QFbHpQVAoI4l3A4P1PfWgwR4lKIWc
nE+VngS80I/4Jb7WQTxQo793Dmp97qmM5s+h/DhxpK9DnUQd96n8MH0deHqVDhaSdc+xdA5unh3L
lhbr67Zwa67edzpjMuVk5V0wSkdqprzW4Or4tb4t9Z7Q1SfTQ0DbCQzO68IOhX//KLAobtbSopyc
9EK0aGtwFXQt5eFZOI8yBNLh/+y4VPIrDQyNQRcYSlxBMdnlZyulLak4pIfz34ecmJoSOJGkJryD
V6Buo/pQ5DfgVmbg6r6IEvj0zL7WT2o7WEBueJdBIokETMiuBNEChitWXawP30tTynBXpdXUDU5+
iwmYpZLEqCE4KSLUq2lVDd3hU29EuJQjEa9VmqMh9d/NlI8fZGxQru59V86h+TFCI5tI1oDQKByI
tSUnkA7YTUw/UQWVrHX/ye5RAuC+xEnxHsHLoX2j0thM0u82OIJIkAJyhKeCVLVIQXlVfAiJymQX
Zrd5c0txY4B+ktdBBL+3jm835hTGfoyPlicN+zazhJ2am/l670sArCZ2DW7ktW3rhMIbB0yL8ugF
ZyRo9yiuaio25+mRbj8xa7KDZ6eZuBC+x9PSijIp7035fWgbfL0cIemYljCPLnPvo36nQWFz+pAw
S0AtlyUdy5aMVx1XqaAmB+uV64GKajsg9vqYPm4jo8dQ14qoWxfqEmKwEAH/F/yQ+QBzjxpBE6c9
l1WUayhx4Iai/e3uIjuav5p2CCR7faIJ5FEw5Fmdsd5KwPhQDTCpsXKPuOEKWTsymvfpxxMmFk4h
wnI7WmPkiT+4TYFCzLpghesC3hasYnwtBe+0xPFiR7gv6To5YXhKvcPLjeSWWxLokI4YsPiBPUN7
mw18hY9+LzceO5ffIaH885RAmyKT6roSpmLXg5c/Nzi9t3YU4pc5fnvYDZgGnRQ9b2oH2fPxU5UZ
6M/g+6MOuVY4H72zTt0LqCjM4wfun+RYA0lg1vzoShwNV8ev8YgtsG7F7/yv0ct4NN6mU89yr4HK
S/o+/84CxzpysnhJ0nju5FiF2JMP4t/g2KNm0IgYIFhNgtQXOIP11bBqZmWfyxiEk4itHNyf8PTO
ighPXr5SbKWEFyglD9ZumhLGcCiw3jFgiuaK1aolnCgXClAaJ2qzbikuTpMDhQba683usgbJY8Jc
EHuzqdtHJO1538RqiHFryKuzzbr4anl32CNP3V7f1BFkGlwiPnaGKHDDJ9deFZXIMMncQq41y+ld
3D7mHwJWSX+G2FSVOT4j0uQZ3QM7BwueIrlnZNG7nt1e37f5FOdBmrDcq9ikKxf+xVbiust8ptvA
DFmzeIWHvFfSi53Ei19/D2e3H+mvKtaKvCARNXmBCb7UYHcw4TYxrRut8knQ6WnUeMddL6Za77re
p2JvtSzCFoB6iWL7S/XwFPIfd8S4Rujx4zxBBlGSOKM4DT/2fY4Kunxdxncdhz28jynVZ7VJL+gR
3H3uO4GHT4XEaVOSRIyf776P/49Bu+Pcptlyapbjw1wT2hnmzPEepuES8WPo7FbGD3b8y+thlucO
NIP4OlLUok1vRiphjp7dmnee3N+T4sXJgATMzXGckd0Tg1FFpYTsobzgnka1zMOD21N8M+J+ZdvF
EayppyuN21B3Fp3RrfmdNWNwL4uuqBv3kHJc0YniLeXWbgM0qwhQPACo2qfKxSRnGlWATHKpIc//
TVe8ulnjucqe925K0t5C/DgSZT/yHG8Niym8VPQZGlBxf1+ST/N338uMUHutKNvPZ/REUsM9848+
XGkK6g/AfXh465jPrxv4uoooojUu9y7TxAcK/gPcC+KcYcu11ONcQuN9+8X/+83CQBNqfQFjGNkJ
MqvBrAvq+w+/YCGxUHo/IuChdltfmJGJ5d0VIFGYJ/yRwxJnGtAqHeaqt9KqiB0Vc1h0Q/xAPvUo
DPZABfc7lvmJcSBJLsb/jcoVAdoT9Fvc306btORxDxxg8ma9ne/ge5V1hfAkKzr9fuskLcn4NsxZ
HsIwLuPjcK6xZHVHG9igHwEjJxXw7Q4EtPv0VX66v8eJAw9toANrZCk2Ztm7VGiZX+tnyi7kOEyK
o+UDOuiZCX2COtjz6R2Rj8dBv8HYuDH2GW5anyeY6MNMZMVZaHWZZ882ZcatkQQi7avayDXBPqMc
Oh1WOxKB/iqez0jdAJB9SZKgzAmNovdOfXBOJu5aoD4GH8U46qvDZtpIU473oVVGgBkiUD0vOZPI
KixMLuQUSRzLsGQBYcxyxu7cHl3BW08nfWMcEAOyB7X9xh9k3Y3OliNgCQ2ibA24fljjRGD8SSEP
rnmkPIJYDqPQkew0pqF+1fHiae3ggxtz6byFYBPfp/q3nYKNUprOOOAFpKvy5BmiZ2SiN3SsrM6I
JSgMA3ixe0v2gm0Juj96kTjMjlzuRyn3pJ/hA9MtjWt9rLTsE7XWNauMwknTeOLnYKpZA7FixC+L
oHR6sYvAhEhQCavVOLO7tXkDufjJoP68idIioiHFtjKlxxxuhRL8BGzo43gbtYiVlqL2ZvqsanWf
fF8jm42P6bNh9GpzdTmjrxgrv61foUBOmPyTDeffRqPqQ8GmqMx/9lkrKQz/OTV5CCGE844XROjT
75Ok4ltAVfzac0ce9nv3ygE+m5mskiPvakwhjIWOJdxI9/idY01s8jUnUOJcMxonuTp8ixPJM7zF
840V+NET5mhHIionA91/0/MACSsM6ueej1W0ADLF+uJhdtZyxixFIUz2F3IiCRvkEvwDM8ySqtVc
hmT7kl2icaV45cNT1NcfEuxd83E5YPfxbVHkAMotBEV33xFJkCuyyaw8UdgP/4oQUhGmJx4wwcVN
0+TzdIVDExICf94WcaCuIFfNTLsLLjgtW7vkVnCJIkrvNvMVDZwhPeBxIuudpfudBkOU3rbF9Hge
teXxGN1+HP87NaFk82vS8R2oFSFlE1OxLVa/WH7AeKjUWVAGSJYNQkicUWJjOYmHzir6XZ+9FBcN
l7HZ04serVj9xQ4pSDz9kvKUlrRBTYnyb23Hzmacht5p6LB9jBtVpr/0jg7Yqhe4KRjkZDN9s+DI
G5ur78RC5d2M+ictWcoW2mQFw2kM2fcE7D3RLrGmEDAC+z0pFipv0tynRvO2ddNuDVqscsA9sTTm
c1GWSUpVZRDRNQdtPdhN7j6iQXlUUsuQVQOJVzqiQdqdhE41qGpKPV7ZFqNIjRrwwS0/tAqHdlrx
BEOIbnG3fUuuFwEagC0bJd+OaIAlw+OI5aV0nXZaB+46p9vghhdtklJCEx0z19w9V9O2o9fdD2XC
UgT89KVk9/5fqANx/UdmcjyLofzf7bXCZmJxSFbxRiruPeKXKXfSVWfOON6gmEAaeXDEYsOZGQkl
gyrs9P7pwP8oDh3IQWRpEv6uBix0QLDPh6PwWEr4qrev5sBOFwU8UbO7VZvI0Uyrx3aY/MlV5b1F
JFlnjqkz2ZRi0pjpmw5b9lxhYmc2doFIi1V0kWUtV+pvm7M7xAFmzzF5uDIlNcAXGgRhU9YKwJ9c
YR36o+BQbRcahkUdQdG0kb8Bsvo53ZszP8fwEhYZVma6TDr/PavybSdwzGT6usnn35sJjxN2WCvS
crh5LCjPZMNEOU7ACKN1IrY76zJZtC4lrfN8Lspve3VaUJL6l8SZLjf3eaHz9CBNG1RaBQbD0yM9
rpy5hZwwL3E725kNrzvbb+wurg2QAEdbA0qOjFurJ2vcGpvyomyw7KJpLUJXnzv6XLnb2AXBfwVm
XKnHEDxC1xie1+oV26HEAahKgatbmukxiBMLrvJeqPnsQ4UCwCRmPGds+RWxQLh9Vs4iGyp8xd7s
t0Nm/kMJNdMQkews+HGbcThYamIYqJsexsV7T6EzStvJREepTloTaJ/TXxZd+YZFXYvh+2YC49M4
XB2wsDd8MxloB+Xfj4eXZBGJ675AZjbaPB+ngwkJlvN2aPuza46lNJNTh2w2NchAwAqjUHSqi3+n
i9iNW3AydkW8BxOJLeuStOakSNq9yfoKKYgjN4YbD0kAmQEdDBiAj+bXSZS87teGGN/WUuZdNgQ9
gWE+F5D4YObJw274E8axOcnfWExq21likBQ4wlsVcs26Q+7yPLpXcKdrUAEAkorh59DBHhGaqkUS
hVbU8ppQA0xSZ9Sl+UJB0Y3cIsazEV4O1JsZFtZ4wCdzcxiDbhzitI7B9OffB8EoJn0xqVTL08fz
1cjwVooCx6TeUH9kTZsoJbJAqDsKlfVxy20LlGepe8NGmWAAjB4ZSGOtOgUKZM8w/oNkEIGJ1dYp
Gx4omYwtCSXPs14trQOhdi48eX3NL/wINC6M3jo4PmPfFW81v8RZKdE63bc0g4kMdVniRqESnHOh
hjJQn/Vmf+AqhCKISK/pn+v7zLkfq6hrqQRhy8Ga2V/yZN17uMDc+dVR4PAoZNeOIvORCDUm8CAZ
Uqd8RkA48nFirdOLk+85rgT8mU+IGs2UZ6L7Y9gdo8XNNIC1uReBIH6A02bStOMNUCvN6eLyffmX
VWMZIkTuY94r7Iu1HVijqXqNb5hK/7JOir86i7sRRfZREmVMDcKbh/8bhpJVcJYYKruDR0CP5fzP
190aqqIqNTa5ctZPeIZLxeuNEOFBo9r7o3p9H0sWAJ+LcElB6H2u9SS4hZDBHgOPWPGl7ynsU7t9
/vPPo6CQ5+L41HpXwZ52q4c7KaZzMZtQK7ZL5BOkE5P4Z64oZwYRzcgkLmqXC8Q4NPGz4sbmPqAg
JSlFEy/SqzyN1bxLcVyct5pelzaUHFRpv4rzpG7luBttsMJ7kI733B+PSh0lpT7/O9NwnYR5paSI
I4hIgYBTNd3jm4a816woAnogukbmVoKxxQkI6MYzgxPUqu3McIBMMY2rNW31XJ2FznfVZ9hZ9UNZ
iw4e9MO+ZDQybVQOKVyzor+esvkMIbb9KHvp5A06bojiEWNuGpIID75T4C8cqjKw3bVTJwoTHEYQ
rDRRyHxB1Q2MKsBtFz96/vN6iCSgQqGsulZYglvju/VQ1usdg/JveyndN0M77CrAnCe5Gn0Yahis
2mTkTbOSAR1qGu49jPHJMpcQACzs7PeD5cKznxU4OsSI2MJHkLQ9yAqkYYaNH5/B3Wj9pBf0VIWb
+Y1ZXZ012Epix7jxM0Ro/qd1m+ulwhkXK6IXE4pahTyl3Nbx6kElqCMYuyDDHzwB8ZoovqHHXtYr
6oiFHEvsPtNWZHy9k26nDXnHRfsfr66vbI00fZma9qhivzgaFpoDbZl+jPxmFgHtaCcwHN5o6Had
NlyttHireYGaxrCyX8oSgwtwdyH7Q5zP3ydHNRflWCE+qs+amuYeKRqm3vMHintc+o7+H3/ryeps
y4luJYhtTRPCSeQdBHcCtnsHcTmVh09yjQYWBnpqhGc8Wv0mogqdXX4yA5IUNo6RsOxLeQVhKXKj
sV9e5jwqsTG9uboFwxROMAYv4G4vZnIECsF3ubV0eaiKmIXU6n2lk2t9Gk/YkNsHFXMNGMggDTgT
UjozbebnI86FItW/u3slVGY6nJGLww42iWVreNLJYQmL07tJGzns08Wpc7U+pz4DalGu5UYdh5Qu
wcxkqpvdCcQjBMb74fvZ+EX/N2MdNosmCyLGqcmBd6dltgeZhTV7SeWPbwSOSVIxP01fNr11wqdC
VkNK9YLi5GiSngAAVaOHjfx9zDx4wEy1dztrk2WYb5TxuWc3UM+7WirjSinBZYZHw6PRb1/nn3wz
MOG/1WfMiIvuQdeXvc3Fh/FEK5t8jT5gYX1DwgJtP+0RiwR8DuPHG/O6GI5Jm/Ev1onycef6gnwH
ycYQHa37i1MIx9qVY4g11JFXbjJ6KNd2O2Ak9SF955LmaOuJ0UhATKcMDj8IyXYToBTKgHfnc5vk
YJoeQadBF8aLqyZItPCucOeH8O0/oHZbGktTyGwU6nrTlgKiQSZeED0Q10frHHQaWRVysV6c0c7y
jacP2ITI5SKsen8JjqvbeqRlKaMPs6k9a8TEsLmcLOxQYYtlfQefPznFs7wgXVAzcxjGwOGdW6dq
mXwj4h5OyP8hWVK3qDsJUTo2FoRgdIrTM5fcPRzV5blxfurcZ5jIZ6+++DcxTnvczkpu3zno7fDG
JvLlILkt53WTCbdFZ3604CbwlEEf3F9UAn2brlb/PcvA5MARvVU2PZBl69WC+xtLvwdfR6RuLex4
KkJEO3roJkDssF4otB/yqKuJFoOFcJR96wk9CPiHPHp64Shjedu9lUc75zNZfoR2Z6E7XYHHL60p
Wv3jpFexBD3uZ9YB17Vg84AkmYif70zztS3fyOX87mbixi89tGlnhxgrmUX8c9X7L2yXkH4HWga+
Pr26jqXhrs0Q8gXqi24nOZ6+PT2sCWa9AsrEjeeK1d7Q7eJexzK2pE+k7cwSh3ZMyp/lxRzvnY6v
UBT6BiV1srcWJRYNYtxbwggDkwPwe2zvD1Sh7yp8feiVLTPEFOIFqWf6XfpoVVFGWDDUdMSNY4BV
ZIDyKmccXSz21JSBTyYoRBJOwofZZGAVTm7ZoA/NvWo7AFdZGZLrXiAH+h5PAiS0VOFjmiN5K6Se
ruf28xgK2ye5deL0ABT7EQpUcPMT/vAnnBmu6RdM0YuGrMEzdz7GqWlasIlJTl+dlaQj1/MIIfVo
RbutW88ti4TMD05uJNfddefOx67JjN2Ox1mmx2eCLF24Kwze7rt7D0RbHR1K4J/2k8vyIbruGLZA
aC0lYFyNQ/tcz++jUrvMf81tKhwJcz+OQFX9AhwH0zykapVNqB+XXnB+wa8DgRWUXl7xiUsHQka6
b0T37zNoACxp08/dEJqkqYcYh6uVFY3EHrEXpXa0ZnaFJvdspR7syNvbJKEjPxZagPFtl+jObpdv
KDVhqzC+Tu4RqSnRT2O1b95RCS5HWPcD0UwKquFcaJG8enZ7f0jmp0aiQvFUzomXeVCfXM1ta8Rb
yc1pb7QcxNLGR+wWl3sEIzIbatLtKyuZxkPJaW8ZBW3RahpfzwixnAkzK+eIoReVFiYLme2u2TDu
WEy2ibzfZM/ud/4ExM80BnoNFHVRWmkVyC2jJg0Iib97qcnL06ZWe7/wyIo3KdgvO5ZWK+aQGR34
N5PcsjyS6Y3OOdOKt/dvP2CS3SQFzPoedFK1GcYgh+jCD2YcVaQaWBM5quhoOzyy41lxjY8Jb1sM
zxrEf0HPsBf5ikKn+QluA4FluetAtdN5K+EYfh1pX4xhdp78OA9nuBs7fCxHPjtvWF8p/+50nz/6
fECPdFK7ZmNFEkt/AqzxjfYUQQWNNST/GSQIKe32oDnuqDb0VnLB43yKBbUWsrEVoRixJFyla9Vj
akgtBebqfVBDBR6XqSVCxl/XgOWNpmldnM75y0UBBwXs/NQ21F2D/KB9aEuD9wXRdlDetLM0Ywm5
ehHrsttMJDeteNafG1Fjc1Dw2PNzgNXCVC5OYQqJ5E1XdTSJqsrM6dp2Whu14ky0iU7baO68ixvI
VvE2uOX5Wnlq/sv0QfnAHutAeAEP8CHgSgEAwKa0s0hO5tmRTitFuJOF1PMGAv/wls62ANP84g4g
EzPdDF/xQnTEUWpD1/DrERD+bx8YX55kbB43tZVUhx4Ar9t2xXqr9VVYNT+0jV9z2Z3QMhM7Yfxo
eIWNbiEtkdXQVLUwIiXUOqUspZpbmrU2C6kEOa3A9KBKzEFsUTmqOtkwHT+4cqW57T5nJ0xn9+Hq
n17xHd8f/QdsPpnb6YjR03/MJUVAUdSNBbyBn26n+ladfrbjxfoCzZZgaZzz2sI9epU/oPES/EML
pu5qLeSIAwMcPsIS0Q+8ZPIUFNYzN4gTskBMq2YoQB2/kgw92g/hFaIASUtXD7L6GWhzDM+xHObj
vePLaHfOkfJ8RDI/BEkeg413eU1qD8qY5rPHmSniH7CUYZMu/czY31JuP/br+sv7o/HSNum9ITfB
39OsuM7MQV3B/om4mBu1adKWbqclmaRphnl7I9DvWWSaiePiqLG3loMh/2fWbQOdnj7LutYzFx0f
9PrdTXFh6HuQzBpjOVVH+tjXBI3O4kLWY+6y+n2I8KglorgOGnovYa8yXyMpWPxZsoqIaqSL6U0l
Bjs3DJcGHldmtA4Et8Z8xUQW2F/mtlCYNQLADVBLi/HjDSC2+P2tspQzDGFK29YarbkrhIxC9xRq
ukFoXN1TvX7wh4bMRhUzJNG71dOE7en/pe46HuTanhsH3fiUo68afMYBGLh6HbZjNazWUNIbV6CN
Hs9FKUH8HlYidfjyFPuCSknPQWgMTJCbXsV43Pkt8bWu36BXzomOQH4RFit6rlDj4qEOdiz8v/dZ
ISPCnYf0aKJigHE8b+TFaYWmScD3Wt/jtqshTYp/u0GMiByWfzPFYixv9dD2fH/SR2AfhmvXLCcx
gCf7S1PzkxUOvZHHfLEdY7Nx2fDHj3jaseFMpuZK4Gi+F8uHw1wFqEKnS0lo6NsmWkTnLSdQHKwX
sjNKz278AZZXlPAAxbkh0bpHBShtZ5bxOdcXg1YdESpHuXSNzHRPbn4Dd/qtC2d/BKpm96LXUCky
4cgx2SzfLC/FIXsTYNZblmrU0NMlGm+CYQZlaxYePTil9JIf6Vy4VDTYhXuYj9F62xIWnrnbtwy2
0CQYzG2hwrweNkYe7JSFtIRnX9e0TG3hCHFuPiJAsfXkSyxtCX6WRnh5jxZwa06512y1SiPUwpV5
JbqQKrkZNHo3W5NBqEZa/JgGNjEt1QeMAorZA30PE2ySrffbLvmPDyyfnFLLtA6aMwsmij4V5rXv
3YyGJA6avErDVn0cuSyM5ZhMmtrPCRid1lVyXj9mEo3kjC+6lzCvBexoF7qQse3/vSMUtZTkv38J
lm2Vl+dYMsJ8idmY5mLWFSwWRTwWKCQ7uQ32NaCqVTALiVYgEtCFWlwFzngVUUK0d5ErCiNn9wAV
A1zdFqBBO6Cp1GhIDnXfpfwoo2+Q9+wfUGEFLmCdSdlOVQjniH/3rwyxnbvuHnQfrbpGomhHMRY4
MXN+TmKnnWEVdWh8hvaCI4+9tc+VEASw1e7HSv5RO8WCiaRqYQS5+7PhhSXlTW/ekIzex3ZLnQp5
iM2hB2X5geYzEymE0PgXwt9LS7Aj7KHegpO2QPrzKKOcaPjJ1NNLJPR/x8lSjXP7l8EKR+cWb7Cq
siYD0YFsTx+d0EGM7upsqZKYo89AKKEXtHHxbzEsUCYY8GbzNDh2FLxlPC70WIm28HcW7m83YYeu
hxc4vopqQJ8cX6BnO95gGZNhFxiU3tIqfok+23Pr3xEZDk7ATn17Y3S0rxQXzF2Mw3B8w4TSMRbV
rBE31+eU7k5oArzJzuCgBCm/AwcTibThsCZGgv5ZjwN1ys0Qaf1v93rS0QsB+WQJ1/JOmmhRoOHH
v1g3r0RaVIR2ijj+ZXf37+BxgLsl1LVZRocP7o/W0nQFl6VvInzzxRVbBXjm4xjhQEtYVR837kPl
HfIC7dL9434rmQY+TPoNDvy5TbUK0gU5b/sNUWLQfrMhisbV/3AXQNZ4bh1RGBBPwhENn+pEO3cV
Jc9GxvCQUqtE3b4DAp1hS+5N3dwD1aMvJcjVSVOgem3RQlH53fh0lVwiC2d7l1WXzT747pch9ars
JNjQ4Co9VfAGI+tCQ0OmKnRA3oN49AbQ+ZZ4HSbI6t4x2oO39S2tLKg9y/4P66fRGRRda50pAel5
SiBIcX/aXS0NE7rI2zc7x6/mtGUMc9C7Tq9LD2aKeW49Nar8/M3PGrgneXdOkMffvsDrVxqj/KFp
Hurzjr6vB61usOEh1VY4Otu3+c3MxzbeBrK+1RIw4plIZtgjI9f2tXZ8rECFuppu/3MYxjx+Ipa/
SEYMWfdmtMpJHFYOnMDgZEXWDWpA2nHx4yIwJAYim0otunCrrYChB2TvG6jyaeo19IqOXEj2BgBt
OY0PaexnUvCpKy8Mg9gZy8MrWsGVTGCOrOKixUJxFrbhPrbAgIMjKkZgjWYgLcSZNI5tMxvFA2wm
wllWEn9SNolEO9H6vBI5YAEaNhQP2FIfYoQAuH3uCInxMK/WfPoMfxudFgcdoz8x23+FZBLzjSI9
G60IbFAM6yx8rg2lbXD4bT2VUv9mQ3nUMC5H2d3esGvChF1qKwSi+Nz8DraE0NHn64GsC3Mff1DD
7IubR/Af7ciD8lQd1Xz8cX91MBTEUW4cB9klS9rOo5Mz0IRmW6g8EnzrBDTccBVQ0e87DokvGSmP
irLohAhSnwJIgpDDpYsnH3nZCLTK3Sjwgb3IRZ7xwFmsNb88zwE+GXIa8ukl8nCogSIRt9Z06fG/
GAhSGsmOUZZU8ZITeg3zNfjgGY7QeGkO6HSjyYm2m/bEvqEV0Tswepd0yUVhFlp8eLwYzvumianD
U6srJ5C7kvyFDF87GpBhNs1vMEW/t0QpUFEDlv1f6Q3awMzmi/NooDJTR+1i21mioS53GbMQ6Io4
qKYlFvbWRGkFhS7aZSXf2NAken3WDod1ATGyxaD4FE8CYrh0Uq6rYi4Xh+Sh2ITD5VK8ds2dEWCg
6JbrNpqLuj7N5+uy8rp7OzgPxM2UQrD5Ui9dIgUQlg48w651/y1Bbcq9CTZagLPOusvY+xUxUFYd
e2nj6yiawkf7RfTeufUcFKkEktR77L5C4fI+2HROvXgWsjd6ZetoIZUifCfc2IasNSlfuUL7/x0y
2c9a1KrBqIcjiOTC/nkpg+SE6tRRSY6ESomZh71Ygy1htdqwkCFD2hDY4FEW9B254qea3u+eHjsa
hORx6/k+8pwUady6Jp41nSQ2wedqub++I+kXBQigkkMTGJRVXNp7aCQnyxhGJkn9dz8VVmKq37Q5
Yiv0j2lcY613Kv5w7bhiPaoqpdaZ7SKeSL2vFS5oUpGwNWZ83qTRkFWsqy9gcnlYr3uzzTeZObXc
lFmlHTm/U6UkuIbnGuzEildAGg6ZIraSvlbnihu6tnDXkJz/GF8g/ae/PyYUoVOIebKQnJaLLHxx
E8yrDur+u7CtyN8MK4Y6DrcmsXT1CxZhEDoGUQjzZ6EDYQ7quqM4WCLjtEbtQvxGI0XhT4+7q7lF
I2WgokU98vB7PplMlCj0nb79HUqCKimkBLGvklTqS69Mr1SO+biatt0r7vNmF/jCFWaRf/8ycavi
dyMTUk7t3JscuKikrFkJzpNE8mvUrgVNX4VnBYVuJ5nJRc28suMWSGl7+cGp2B+KZPWeAvHvmGYy
V/qggtiy2Nol5yuE3NHLCuYZCoRbUIQj2QFKo7q3olhP0hHDTjN+8VVFxXKvLUeDXHbXDA1yAOVb
CzXeeIOdfneS2iadaOn07Ewy0/9JtNjiURI8JBNSQ8aoJalzmvIcoCvpruVSfyPBU2p5EfevrvND
LAYRcoh1xyI+2sGlbJvE0CrUwCyjsi5/7qi1CDfvg0Mqvio0Xh8bMEPDKgiumedn64eeWeSo1qap
bTTYjPjpkx4Gbd1yFFDXkiElBVomnZMo1JL0uHko2vyWjJ8dgQ6bDxHUNpAw0ok8S0GhwSnx7UoG
oUOYngTWm35PuDgZfcu7dKsU8Hnz1wuUHhN+o7eZqcrXvDT7WRO+FU6F19sIE12hAjx+MhANzyaD
pYND8BtaDNGYHam1+pJ3hvgm1/uRXl8PKX09Wxh/DsSFcbuQtiANXkOW70LlaR7aNutxBjHQCyiA
GAPSb0dQUe/uXITBkfWYbVKV06s9IU5eihXiyOhJwivbecCj/66iCHHON7S7mdHdzyJYd+EtsLi+
1REzrNIu+rnvuGX6xJ3Wk8lKHmxoIkFWl6IUVEx93OEwWia7nZJMZ92fjHFEjxNC2HZjDX0rL6GH
E+Ra7gZEa4DT9bzDsbj+59vM7urE3B8N3bwQC6WzVq8aqCbwT/J3NPd2VhIMptd7ajfEbpiFIvxP
ycNXbdroZ4ovD4Y0pfl7PkvN7CIKavnXaKwhaVNgqwdSi0sf+iINEZVnhDMS5300BpgNFEJ4i0Q0
RY5ePow/hg894gGzFw1xHcDxsWUrSbBKdT0K8tlSTTZbY4MtDYeMMBie3tHf3UVMiQE8hPTaZVU7
wj9Y2U4QKpF8729QaGdaCDrg/BAiKiOIhBotGXaPFyAvt5G520PU434up27QuR+5K/awm1Eagq4E
KHY93acpcC1suxJSsD+IIB00r15kD8LX1ocAkCVKmhv977GmY+fSVSFyX1d95E12P1JDpmNzCFTA
fv9fFijHs4ovUv2mHZw/zBu14gcWYYDBIjIAiPGiuguo7jnKwSl2ZUVuJYg//6pTAXP5XMPLO27s
YnKF+isNSF/mkzv+OIFzuTQjUz8trf+a1vVQnfnp9FnM8acbwbJz4Bo9Op1FWi3P4TbWx12/G5GC
8WE5MSm9v6500tmp0H0ZurI9df2ZrB1rMqdo4G/63/J/p99eHv8rOD8FZYG5dsSJuAZYAfxlCQqG
CQiQ5uqqVxKytN5PYpE0VQoAHngCGb5CHstTirkvdjUr1R8+Uq+DYwN16sfcM2xReZZleVZzVpF1
9/mLHCr3qmXv77I5RKWcs234kowiRgSC336OtWq0zyRNzY+yKGn8ZdEq6fkPkxwiiSURfQIBMEqH
j9qL0wMeveyutzI4Pqg2bcoB5ZhQ02iNUpYmczrQPY8giE5HFv94B1Uqe9nAiFWRvAjy5pXYJ0lF
VBNUBO6Ql8NGgxMNw9HGffH2X6sKVum0ohpkkPmQGNEseBKSlFmx0m1tgVuCP8K+yzCNENGijlPc
0nPMMX0hzBDPRWmeVlrjIyDWUO5QX48p1mHlSTEucKPLuIU4jIe53nVAlrgPAEn8uq9YV1GFoS61
05IyEgcDXDHVaFFydoTVpxYWAoKxmDtmbJh1bQU8YiNd1Rx3GgI7yAP623eLQ+xaUOJ2xoeardeA
be4N4vUbXWgNq0Q6rkg64RLAU9WInnNFDa/Bvw4SzxsHowvHoRyQVAU3Xf9cBBH6BWwE7JktrLwp
mXHdCapsuRogK+oZ9A8jjygXr7348ryMUd2s0TgeXE9uJf2RKTJNFENF3alfPAbnVfgOXpXfJjYi
E2z6G6WgBxMYocSxPplpTP5JnXSfbP8I6g9+dO0H9I4s/0l/Kd+t1c85sX03i6Ff4MaDG4ihMXf6
7nbuyqULFgWZacajpTBCaPIwCtEF14XHw2HqJYfop0cXJepZEA14VwysACOmPaqRrf1yQif6jqwF
ovrqHgSe8nU40/bJiW+nipDx7ZUcyDpJkpguGpH9n4+OJguTkjPZ0pTWZPZeIonFIBssRnDiVGSw
4LBw7uf0Fp0tkUIf5O/Q9BQGm9xqKc1HFMbAgI2l+LHIG/TtKJdGqxEkyMDM7rLkQOgT2u3ZfjCP
c9ZVLaB818TOVlubhhFyGESWNzH3UTkHQxCjnxp0hYzVzxTVeLGS5gKkkEXB+mq07rVNFviTOzi+
C50LbRuupZPFYo6qWZk+BeSRy87lXnsfqae+VTmewqDemQMjA0WPq7+cM4BSlhGVfy6ZR2CnRxQ9
+5bzzr+cia9ALtpFoFHbydfrGns7Nc/dcsLvtFZbtNS7ZNpxU5PzItUmJRsF7z80YtgGSxUMjGfb
nG1vOt0S+MjdfN9VKrJQCz9qrFmF1FaxT6Oz/NDxwlaqbXYHUm01LgvolNcmOXTwgmZVCiw56WtK
Y6uuwe8UqKt8DRnLoReDOyRHpd5SI+63O2KuK1Z9SWDnOElPq6ZvWX0z19/hvI+y6xZYRvNB/QJl
q2/QFsqMwWxGaxNT0h7YrfOdrKKzO1Qzvfc5fp4sp96rXNwuHDCJN77mLk/bW6qMHAjo/0jzyGKc
fUsE/8JeYKHoR/PYVlgUMAAuQHFEXzZr1BM6qOuGGulgrPKBcE5c3qDrkXFfSyaTLoNEzrVjFR8g
aaodw+fv+5+8wK1amMWWccdj07gj34nl3M9cd3imw48Wh089fFf7VgkgWCihnDtoh8QY4dSBZMaT
N7g1ok7RPkzXjQx9pT+AY5m2SHgTVFArju+o4jemQuvBO2K20Q0DpV55/98GwYlSQtO1S2kLPoID
u6mKRIdpORIn2v5AnOC/jx+YI4yjcIl6jLxGq0C9lHAxktu+h6EJrt7cyOQ2PAEKyABNBMwfk7RR
waT6R2sCCzAN5S8CzMWP6BN/uZBsdUCaxBk+vmQ1JDJZp/fraQjj1d23ZMWBgdHh7q+qhvPOpAg6
5nFWc+GoLZrXOjMRsmDXnIarfHwUJCc/KkLnT63hHs/quydkTmksIOlChsYqf36d8cL6aLAgb1Rp
X9OnNG3+SdlyHrrerzuQ6eijzJ/OMO8k6tzq48yuRPZmJ2D5Z7jzbFB2G6FiO0zKjS/UO8G62WxR
qurmzl1HJub6iDkzlGPmFBkrRNJccMJv+GYp4BUu8xA26/D8MM0FEIyhNbPxbetehYIZNcr3byh2
akkPV0SdhU3kaUOgWuLiaJ429EGUmhqlTHuIsZ0KNA1MG6CYnIMfU47bHDPRcD6V+1KdYthuQbKV
QWDbO3MsDxat/mU/jjH/uGFqKYE+GGfKxT1avnK0Oa07PbbiB89EbnN9/Tu/lTnzXsZv8I+/FugF
eX3/f6eoSQ3Zynxv4bMDvjkZ2n/NGFLQsLlCwO6SmfJs4qVkM8d2T6GBddGbc4+Epht16+Vadfg8
aiieG2RjOG9dmyXaE4sLw2CFw2i03FQD8DmtMRCq0sz5psiRC6osHDNs9Fexi7LxNLkpYssJ6fLr
xaqd4cH+nr4oSHlxtvjdz4ipY09TSVdcAXocur+IxA5UL798FjK9oV8aOf5k2UmbhMdZXGNjk4KI
BAcmlOTIg0MlpuMGQjD+JrVd71XNJSika9KUca8PY6FOu4qOP9MP9igVKjz1oPKX8XUwjOsrU2R0
FblhVOehx6v1ysYzIsJhD0HF44iULEFABlKGLPIz+cZd0c97RkJ8oPhXzRMmximVUcYx50lodMXS
4DcLIVW2yoPe2wO8+7NugjtoMtPR0nf4n7fcn1mBqQ3r907q1xO8+ChDlg7rifRcTmPvNqjl7MZ/
dheNLuxDJpxaJlu+ySeBsXomQxj9UhCKqpqBK2xuS28KN9t/lSNqYyjb4CVFAlkAzEfz6XqweYQj
RPCdxttvWVIjPwOODPeXRBK3QCmukOl80X6H8h8/4PHuZFFrP5S8oTk69f7TNMcoqYtJuEUNN5RD
VcJEJkCnhQ46br6g4qcKaLdfK1+MDJLG9g+W3OuFOjdgUDtqxKo1Sf2Y5q2zIK+0WU8pyKlBD+5X
6G8P5E1KpE93I3ITj7JRnzShZz9YyjS4NI1rpY0mfurHaAX+hZ9pdtcyA47O+1y0TpxV7gO2gnpG
73OubR1lkBUEjFO2HP8dABq2eFkH59kzj6DV0kwQMBaDIvhgPLlPqfT7YbwwHQDxx+UDh0W4LhKe
9DEm2eVRUIDtxSyIXpmLfEV/mtDxSctilfz36Au4SlCBLxVH49BjUpdlSspyYNobhDQss7HpxoAi
ri+Me9XK2qZK4/Krd6UV/7zX1EdbuUH8tCR/lwTwAmMdgmhFrMRtdtstcd/DR0W6mGYF87E/Psw2
ZmOenUvO1TF3p0LunswbHRk1Ml5qUi5i08QDF9G9ncEOQYCtd8xhFa2kC5b2ewYFVwolH+h+y9Jm
jTrTivg0E23ZrXZ8LrdDudJuywjWzXE0J1bUnIU4FdyCITKBgDoA2o3xB577fG5W4Wi8lL7zbrY9
M0BTMd1UbciZUCtMo6u6p5vfluT9e7+kHEhRJpRygyEQ0gmhSW8nwFgLUZnlJyDI9xUemidxUuvv
/8VQ34npId5BI8iUzgnu+Vx0A/wXk9fGJ5MsopEadaQ8JVviwv0wE6jxbk0opsb84GptPhGAQBND
1FUwK3N6K4ZZ7umNs45riP7KOasOO4wWE43MwczQZzEc3Zfp37woJ0nBv/sXJx2r5I0l8AkjHmyJ
l6kdkQzVL0YVZmKTtcjka05054R4h42QnyRv4QGQ++Z+H60+oR1el2i7bYyYREdPkC4w2O0a6Y2l
E2EcFuqc3QBqB6dn986SP59oqEQMfESnCP1daEUvD8g/nZ1WY+/9MWKlBMWPD34/NHDz3hTH8aGD
7T05b2EjTz1DWZt04xHlLYMLMBvDQUXEM8+HhyXjRqkUQPwLQQGYehZi1qW6VUfWn9i3TIroxXof
zL0VUvGiy6C8BiERa86ruH5ifbgRuWO+QLkt9vZcpOv/lYYO9uj6Go49dqTpKMf8oSafSbrco5ez
Axz4e32EAxJKrvlhMrrHh5CVs3GYPpbGXX0gii2/jhmsavmRIvsQYLJpiN+xr3BCxjImNNnfQJ1u
sDG1wxB4vDlzIaPcnFPw2YsSxv2u6Zi2/eAzxqa/cRv35vIF1JFvRxVUvyouFLFBj4A8X4OoFH/x
3gR6KOUr35sVQ0tSoP0jVR/53QxKpPxQZnAfvndoAirQdWjmj6laQUc6E07PC5lWmuKHxUOZ4mC7
MRE5yQnYCz9FNDOTFMal8NHqyZq4oQrsJ/LQd4MQPplpwCmedSDaJVXp4FRE47c1SCqrIWJqbcUL
6sLtzAm4qI3xJxQCTPEVzu0pfpboSovaGjwFNdq+xUBUJqCHvQEXmf04gXz9AW5n/W8ACst4gniR
EvubuNXFpW+uTM5yipoqOkK76ewHcYDznZubJYhYOCUG58F2dL8kJCiyBqEDYahJpEhzf+JXv3SE
2nCIqJIrOYlyTvoksCoEXsCcsOlW57FJLzYtHwqNwfuXJ0XTrp7L+BQZb7Xif7aUGfQ2vMRVRCIs
QzQREu64zteahyzTIGqK4hk+xPkAmpxMg1yhYf/PybNjO1XliEBSzu/c+ZdhGts036WfPglzx1Y3
S21uEGh1CQwb5XbIw+0Zdex2eR6Bc/09tBKWlT0CPj2smBSWn7Ax+cMCz3k/PSr5IJ9Hcmxp1HzW
1HRsX+EtV6f46DwCwLrPZ0BVXzWMHiEksw85IH8gFKf+A1imh8YvCShlhZhcWf+rvE8W2NKN4clJ
eXOP94cNgnyssh1hCo+SlSRYSo7TXQBPXIbJZOaqnFCnKcrsFcqI6r+e/6XMaK4eU2YUW7y7RhON
2DB3nBO7WJBh/EYa0Kdlo6S+bGAMyE4U9Qe1TMfE05RyFTHNpQM8/IBWDZY5bpW/VShiTXTe7czY
tqzKeCqwnGuF9EMIXoFBA7jce8TlmXYw6Z1CjjoIWQg8dL7UwoutFJcibrQ2XeEjft81QAKp5Cf0
TZlFaKcH0BbO+AKenToE8MNaV9gkYUqhYCXPGLyltmdKSpgON5CTXnjK5q89v1v4APNeCicM/Beo
PoN4XIY4UzDQ7JkUzGxF5JdW6jTQOlr2seZVa2mgI8FIWgCoaD6FfbiYe83QXtg4lUwfTUPbtO17
nlX2t4fYKX6MZxP3EXE9dSU7PfrNXFYcBUE0iCUD/Ctii6q3iLf5owLGWbYtSv4EUmqPmtDtGfEN
z9pb3YyMW2IVS0SUfrJEV56qLo77/kYn7Mfl1D799EQp6co8rLCxb56GzTf9bt56R5HJqzx9g2bn
/wWpUIbRw0bseYCZmM/UhDmVjvdDTzDVJmW5llBJjdj2VT8tWEWLsDY+OgfqLP1EKdJ7Z8EJvH6T
oKKXARSPxrwer7h+Prd+idLmvQIIryn8a5yyCJAnEQzTSQTRPBKX3eKpnU4SGg9SBNebeFhu0h8K
6ZMp8dlOPRR5P20gQJV0ozk4g88xSWLk/M0O8A7xrWN73R6wBsXwKdQ8zl4xsdJKrr1UeFL9PRuX
r0zZAuzrikWUEAvyHoLJ/uRitOJT6NPTa2FYUlUIpbETQQPpbA6BQo+h4FCPYnQw2a8DFc5z9PWH
l3QsXkywjOmAOHwfakwEkzhi9hui/Temx9YFyk06ZvcziYPQPbxEQ7WuEjayyKqeCHSayfkrg3nI
aKc0A9TbSa0quqU7H+bIqi7h8OdLYZFTj/nQVM8unjsrbYXJVm6buT4wPzHjLow7ni2zn1/Y3HJw
vYw8f9KCoUNc9k6ufhGRXmtoJDPrjhad7ypTqQ85/haLN0IvrhKWC+RPlYMHOzUXTm6WAahcloC7
4RGiEB0COalr6WOzlgWfh8MXPCAM/Lj3saGHaShiLvqzTotYgW4cabjFDj4HbDLFN9juXw5AYVng
Z3r+ypED6VTr63VqPj+4U8aXTgbhIJxh20Y15+Q7+m6ZSO4NEDofuObMCNqpM1bLusjzXtor2peC
M6JbkMtscJEMvYsJSW4laNvmN7Q727Ekbz0d/A06EnM0WMXPSya+jIkO1GhpGQCoJkBZzn6vtsYx
THiEXZi4PriI/MGSHZdhpgFchsQlFahQ4EcT5voUt5zH3seOc183WjnCIgspDHLN6NDF27xWkWHJ
oZC2WrctedPjnwatNSguRaMQuWLXG8kRpikDoZqA2qY1gfEtwKye6ma40fba6Y42WAwdDYZgshaE
tLgv18aVwphMrTMO+pFiCvtZ4mD109b8EleFbeUKpzA8QOzaWWWKVUESX6nywmKsH8c5A05cK6oy
/NnNj4A0Dxyci/xZln5oXbfLrsv72aov+SJwFiw7mg6zIwucWCfyZuau1caiJaVXBXUqI8SLALRQ
+a6CfNxSuhWyB3Gl989Q3yuiXI0e+AwlfbXYRAYLg6c7lA3byw39D2YZkNoMizJ+MiLSyr+ITud3
k8om0uj9OJRzKzcj44sYmAOBBdj1d/QDDTxyoTt711TnbAetbZ+O+JV49pFtIb8z0sakcbkymdIn
8UHykHUOYfvDC8jLvyR9bDqaY43gRfBHgWHt4wWVTFR+L2C4dCMhlcKjF8em1Csexur54O/NLD4A
UK3EwL62aE7282JPVA7BxxF2k4S18UxXBLiv8MIxHcrwBLhyOzi/lRbeJISj5EtqJqC70euDniip
Sqm7mQjea+45bfwBIM9z7y5lbE0mEDGW/jGKX8PAR0TDnRXysZYSoT3QAsDgKzewtYUTiWCRsjzR
z+E+rxX3gWzIWTRBuQOuCHnULAN+3pJe2dZSbxwEeQp66AW6uRQKQT1IFkpE132I7t0KrVUEbdPb
6O+/X0nXn2MTQAXWkn9tEl8eSqd0EVQoqe0n4aoZbWSMpgWJncMqX9Q5cz1x+N5mrUbykeKgnE69
IMqq1mChG1bist4Vjs5BvEPc6bHMXCnL8i1YVXUj1s2gkaDJeY2rH3RVw8PqHtpQUM7wY5rATMEy
mga9X270wsYXZBK5teOzQiucB1JwAl1rkcxLCaOGyRLdScA6u8flgtCpVdjx4MadGkdmX+i5oGfi
Ypj5HRlq/A9pG5d2YTUO093xqxkczSu2OZzCi9hn3aCVBq4P16brbkbkQo/rMrNzjv8hVWO5tzLE
Rs6tVKS7+zfB4xy+z9Dh1h9EYzJzfTbx01R+ZJNyy/E5iAU/1rnRUN5uYiQtI8wl3dMTjxUznE0F
CwEoBWm7ZfRYtXtYiHrrC7Vrk4++uh9Q5U9ILMASVZGHReh/r98jUUbvlEe2ilrW7B/Nfii4ZJjs
f8Ic1grVOrpuhdsbuxf21g9GF3mnISOu+Jbr9jpRzf0td/LVhmiE9PxqJa9xKNJ2ssA4dVqxNv4G
av2P4aA4d05tbTjMS0yRbxYo1CXxWMPD+/QUnho3LUAitn3DnyJbuZKQbH2mA7IfDS9BYCYLQfeq
TAQwt2pYlNiWUMmAvv6LSI/bJsQ6CjsGdR4CZpzaN6y6p/lOYoXB5Mp4XhLMcpr66jG699zez8Ch
wjXcU5CMAUsFUvBOu6UKBnqVKpxYOYaNV7ZBa0h5MslQTj8SWE6J6gjx3t9hTm1oUKk1kQWzoeAp
C+LMiZAkClzs8VzbFetx/+piQve3mYbFOZQo8Z25Sqesr4vxQ7hIdUwK+YcOAzkfcJAdVKQGb57D
LiqEAcJuDzFZ28SuYEYnaZ1Kxb94IGBCE5XgiIGRNHpJq7Ix3HA6COm+w3osh28jIY7ZpQ/J0EOE
brUbrx4fyIZo8mQnADTrqFlG1fup3aMOjdAylxQd1zeVYN6Rvks8731gwsUl6H/mgwc462QtB4dh
eOaXlMabPXcdFvO3RUYXzYupB5PxBh0xhhiEsd+Ex5RBf/Bfxt2fgjm5JJ2PP9EXpaKPcn6aZ8kI
IWIVy0CkRMuYaAdZvSXf4YmTuCx2b5tD3PP6lQtuKXHLL74VnybNvdpIKweO7yOirwPD7h625X0Q
87E2CyvuQMfxYL2+fwQXsv8bLUSoiCweqAhm58q7Xp/QJThMkmm0gHx8OrFOoTWvplAbkMyAUwZk
p3DVLHCgB8SzI6CEa4wGeeMRwLIgPSdQ2VmMdtHE5oKX1LaZFtsigR+i3Hrqz8GAkLf5hGRgAJuW
QvpQyirs5dmGZ8Vsw4zgK0WDH0wYwJxywchxdbChKHX5AGsAEhYmC939qTaL7jMl4TgYwPwK0sxP
I1eI0PybFRQLg1h8wvP/vGLYLryy5hlwJK9xvQeFnRD0pzQr0i1CqAeH7XhjdfCPqLt6GRZs9a7G
T+NDHJ8eTXJeoNickHBolqxh8ScuyF/5knlIFlOD4zEMnCV8LoLO4TCYIo8zUQ6iv2hF+55ppNmy
gG6vr7/85oI3wFETczuBkF+8Zv/UAeYtImJRQoKf3c4Gltotj0LHWQDdp7vha9g+AIvJsgzrpM2g
/OI/ous3P58s3JCrlgZ0uLd7+8IGHS3puQAENcCajZfatQMucZT1Yl6lyRxcCUABOG4r870APWXj
n8oQgdF2Pb0jc32CcEvrM8/MD8JlgfQsxnGCqaQ4ZYgoteIE+m6zKbymkPrKegXafd6EY93YZ3WY
fLQ4JMHfZVdge2mow5OaGrVQEx9VhWEydFGHLQsrL+1C+Uklj2pFxLb6x04JhF4YojNE4skYsweu
EpoACLchuVhocE3Iak/KCgeFylqSh5dnlfpc48dzeqmc973YxHKpNRY7/AfnuVYfscM+d9iblK66
lvGF3WEOeKZjejIKWFq+lCNSiNKTJuTU3QLZiUfpOU7cgxh7KIMi+cXCs5R881jShjV6uS/umaJE
C7Bd8hrPqnKTo2GB20H8O3AI4reAvE2s1T4hEYPGIrPt0TNcJz1UqYeHGncUFkUyEq09q6KHcTbr
42ytgURTS7pruVkUTo4iOJHBUpQ3MgjEBvklkIbNUpUsIgwuClNsfZIdewR+JKSB2hCpId67P/mj
VcemNBgy/J5BMrBZmNb75Ns2v8+qMJp9zHeDKuB+lpdClOzbLUbLrq/Ek9LGokcTvjrD+2pkNcyi
IwMROaw4cZzpi2vnBdEpkU0/kFaSoHoXVnscnhKWcQpZkFqCzR9D87JT+RoC9BYX0LsEPATgKhQM
P3Vz+IasntfDpW1l0D5SbZ8z8Eg9ZlQhwAxmTTTSx1yPLUEM/LGb0bkbMexN4LiCCNK5B13HBIx+
QFCblTEbkJ+uctnuiG4ZImGavWJbA/1bGAz+6+RojrMUD76ID7VUUa9PFQZAqzXkdrygRnaRAMPY
4Jx1kYpmhMa65LGm6/H0ZILKjhY4MX/5+Gl0ZID5NL36yiT4r+7uXuLqKrNfN/Qscv6bo6kQo2Ih
IbrjI8P9JxKO8GM41kbs5p9FyQEMouEGeMBB+zWVY54Mo+RX540Eusi6Lp5STNAqrKaisoiBMdii
QUNzSlz9qW5+/EZDy817ebmvotgD7VkLdwDTmN3hj/2WlerYhY/JARPMqhRNKRl2UsABwg/cJgda
gB1GgEkdhO+gG87RfjcmeKyoB5MjjF8ZvN9qbXVusOG3rHOr6hPU6Vp1Ak8b7VkffkKLjTzKjmKU
uSDDWHTBEOFI5Hw1/0uOS/O8bq/yXRsrZNWTnWJ0KoE0qYcKSug/J6DvCuoMlYRi7UloChwQVjvK
XBTnuRW15GkL+p+fjcqDU8SGaHDyHT+dvU03oRAENL0Yr/lW3sdPuyaBWu/2VlOexpa93K2sADC4
lKBtRz/VT+npFvvYqomaITpQeKh3KBnqTnuDtq6SevWibzFO+EUUeeG2N26KnN7Q69r7SGc1EC/n
JL78UyhUmVkbnYb3BBtbWWC4DWFNJEtQJwA3Xbh3swfsy9sDWt/K3W2mhRYFmE1738Lnlmi8RrdA
tmmFTdWWwWVi9IijTk1aQWTvhHpIGpy5b2X8FUqIV2MbvuWOuK8Uu500xlKUpgnZUz5DZ2XYAX+p
L3Uw/oGLWw6zolrhLtknpihSnj4LvSLbpErvyjWIZxxyKjREDkLjszqdpYG0FdRTQD2OljdJ7stN
h25k2IkUOqC1E4URLMFt+0MK0AbjcsFV9DFVXSVGwC4wKG48aFj6aft4D0xPlDdmrAJO7/yACHy5
6UyRmdsdWRGhnV3A3i0gqP0gt9Bs3RFuW2kW8Wb9bNuOFoCpCoX8Nzl0VdLUE0w8hcol53iKIiPX
58LLFXNzmWdvx3gfPI0U1KnG2tUeroG9okfdo+VcS+gdqFxG+tPCPAOcM/nytbfMOQ0NmZBYWgJQ
TB+hxMpQTfTEDEpjDkJu2dzSIBEQcerPq39DhJ67xiiaQfkrl03ZZjVtUgPfIdK5VHPa+QadT1cd
DJs20KFJuK8hUNeCZVTH9UB4MjfRiL7zly59HFPr2LqyFP8O4E6CJFBYG1IrV1Q5De5UjpHKHuO9
cDP+t3A9/9mtvUFHk7nkORpCA9JvOpNwlanvXPei4bPEh/+n+5WRmNDOH/PafiFTOp1Tqsq4HxEd
AqeR3YLFiFeH/iaNYSZ3BYTIuNMEZXbD3WzWmbWiQeyqABxZPI1W9z1jg8bHPmfPVArNFD6VgUGk
QkNoLD53sDGtnX4ehyo6vKE6fPXas034HtWX4leSa7uKFFoxZxVrCP6JyMbaohbJHxQQQEVVghPs
QHTJzExBlJ6/t4yfPXKOZov4EwmL5lA431RgOGpUpLGCpKxg7nrtMwS+tufaw414CMs091hJyl5K
dsTYjXJP6I4U9HGhhwDra9gH/kLgaSkXpnHA5lXByPoY4/LV2iDtDGQqZ3kNs04fyAeKo+URmnKp
aTXLXhfX2xpmr/opHWB5LnJpG0N1Xz+XPdHchHoyJ0PKlPJ3soFw0YgFUDdZUhtg1hJh2woV1eM0
vlTph2kMGIZkvtAgHn+84/RcQVudNAeVQbGuHz/ufOktKF1PrfED4jugfTVRgljnCyWM3gXRBRNl
8X8tdwn/2mSFqcEAeOxFWjAOq3Sb3NIggSiKeQhyvuzEChQy7LEhWXR77U5eLgNoNqFzzjc6F4oC
C4zlXvKl41AN1I/zFoF7MEEjwp3GWWe25bzrdBZXv+CSaZ6WtLt5xdURsC2qEn+0trP2GiwQDfGA
8Q8EzuizllYGnmNOtxi1/v1A3DvL+0AlrmbvTIPFThfbDF0miTTsQHbvh3UbZM0D0bzOB2JKjI8S
PB+NQeJ5LvOjlOXchpjemH/y8tJeS7jDkipnVNE6slxbwCd9AT/vbNjNMh9tBwLkb6EXiQcozJCt
lvnsAlpQgj8DcWQpmUywGgBY0rG47PCWQi/m6wzZ+4DiK7+s1TnsShwY69vWvHFnRwEyd+vx4KEg
Tw6Z1bOnfuhCqJtEllynVHqxU3Ar9g6L0hCN9GowmnpYVCbk6JrRyucHdT+QUhpzOMsshsYAO5ms
pgyX5TR/3tVFlAAzNW2jPe0GBpRzUrCzt6ZvIfQtlC8nN4JWhzeMF5VArRyczyMnjPnXhSj6peaT
o+5agrdfVRhOOqas4eaI9i9JSKngXcJuLSVQFu08zsEXvwCng35DuBlP2xoznEc8MHmSgvfZuvyq
5VZYM5tQ1MKx7DiHaPIXwBegcBfJKQeHkKUzwas8sv+Q5D0DFgA4kfFcbNEjirqpOBu94w+4iUKu
TiHPxJulgsSAA8XS1XP6KOroA448V2MNj5q5jz4w0QOK4BR7M3uarTtV34emCIWIXGkzWbRy+aeI
9JjOMwTuE7tMI/8c+VcuccDcwdmf7FpSCQ8/mP9f7thxiGd0z++LqdrFWx+Gr70F6NBnreuSefF+
fsM5JGqGbGCqb7VFDckCt9GCVi47I9+ETePzOoPFzyZVC3v03kNg7ovOIKG2ul0zH24gsyueHD+k
yS+bKPne4V4X7qex1+e/DsNqg0r2D7TTEGtzbRoD5sxNlUd20hHurKWHRod4kt5ZPGDVqxlsEdFV
qJEKbdN/pimf1f+ZZmiDM7N05xGp7Y5P9wICnXHUey6GwmDSlPQGRNVmtHO/ZQ9+Shm6x/7x0cgu
EJCS0YWV7viGnpl8Z8LRqAGh2AfxL1cr5JA2FwkIqRq1IkqeXQ2i/pPHKW1/KJ4hdA42cb+sJoZz
w/kEiHvQl6U09TFe7Pw/YwFU8pKK2dM80PKHfYrwmvZ/2tO+QlRbKhi1afdiEulJFFjZPWDy1Bpk
IJUkDqe7jfikf01GWZcBGqyUnaFdx1/AiF26ZJO2UuOv5yKz+GItEDUVEewJp2a6Ga/cWyRCEqSW
dUCcAweVL30sbayicOIX0bSiJsQO4etde16X3kAlNYsmzCscCiB0zXF0WZCNW7ABkzape+IUk/RB
5RSxoSUeCXaTOG5miVkEjWWHU6XkGtPoVimrKaM9jJEkICICjFfQ9T76IOr0BmT91Xmj7DzaLK9x
bSqkQ65kHly4AB1kA8X+/Ld0WyEzUHFktd+TqAaMlBqdrDkZIAIioE44KR7q801KZLEb4b1ByytA
4pCTX+uz1bsP41ANozkh06Z9ByfOUYC+O3rBI7jQwFZhF8KJSuTidPFNvKmCGEXKESpEvhB5gNC5
ebjO0/3OLXjLn3MzWcX+nvsyJ8/+FYSuwX6GUoYDSCRLJrvnYOK4OtnMEfCUBOfREm0phgq1N1SW
zc+f48fuymv2bg9fBdfTaxIwo4DewPRxwO7h/h324NVU9zq29qfQm/faqChwImXofdoQvj2EG/sf
41HL+xrUkOWsgmQYY4/NEUKBroIkTEPwdyxI4JAzHWNK7xf/oM2wYWq9vgyA4nn2xKBqh1AFCX48
VTEPqUymKfo6tAy2qBM4mJXVbl2AZ2CQLH167N/URDQ8TP01qOQ0wuRKYo6mXPM5GbNzICjoipYB
QiItyi+LNAo5xyHjPypngbITalDAQDvd0LYTLpGGPuiApAjtabsy7lruNdEZwKb/1kOzIgBoMTQ4
v2lw+R1qT2cEh6GdGxDwpo6v6fdrSNy+vav4u3vR5CEsoUdwaZscbaXrBKdgkW77hjCdUXQS9cGs
dAacrJj5ZVfpsq+9j+b+Gdq+DMdU6Q9rQ9gi9hTKobM4m9QjadLeyms6sW/wVUVGXIWnQ0fhYwcG
eBKvyVzmfPLeXbPEjoWR1ghqb+wctiasWKFITE0U6+fKb6D8hN4nXILYEIyQhY/nj1y3+juTAIqG
fPKu8s9xHOTTcbGbRuBtCm1MR/j5f4ivQpXlqqCaRs8VxGvepmBtoNCTjv7hPK6mzyloATt6r0Gi
lWraNqj+gqwATHV3+UX9Tf3OpO3SdPgVT5v630x9/KieUhawqnQIuiB1mVcaESPRzgNpA1/r+OMt
sWqSQ17RtPPaa66VkGGRYId/O8ksDFF9h93Soi+SVKZCoN/qRxbpjnAAbrzMH6GVdWiC4lHTwdXZ
mPrDrHKAeQ6yKm5ukouxbJwKJusa+mBbsOU7m3KCruzql1Ia8Blyn931PGMuekZ4QsYGoaUHSWFG
BQ2w7869vxYp6qRBAZ9EWHpiPanbCacpEYXxgZnZrcIH3wAnioslETV+N3HRWTloUtsp4ZnIxVx2
xgAIaTc7i6VhCi2k89M4+8FbIJI/pin62EUdShNuhVE6bM9pJU0DOU1AsVq1P04SGKzQ6bnilZVm
BU5saJLK7GMgB04cBulmqTQg5b6jEwL3KLDGsuDTa2EdYhnWCfKaXspbDY9PXq6i//X69Pg7Pg4L
YaUuEy1FjPKBzRNacsiIrrAXBwwbUrPwa8izK8od+Heti/xiL2lHfmhld1pww5cZG9/3iMTXDn8Q
NK6avIaeVTeIq2EQ1ixZfoVgf/K7+XB9pNKW1ngp1CHbfwJuS6jIKSCUMDjgLP2DH/djYms/eOaP
z9VUVtVXuE9uV9CaWcGAfGvvZYwVKmS9QGReEMtcFtt19Nv5oUdOCQak/0lwokVl5xoX+F/mZypn
bJcJYGUkmX2Y0aysSZE2rKSu37UEiTvuRQZNMLySZb7nZk+pc9G6ZuMu+/cl2MVSVre6f5ihnpYL
3DNRy65nhVLOqbamu9UdWIiZdnxM3C1lIaWU7jqKoWKxVnCIZC8HVY16Rc/oTb0taZa7EAp8Soqw
966zwB/DJRt93YNoWkhvAJINNvxlCxdlFVogN/hRW/FEF3/rjINcTbUojxydv3KJrj2VoL8DCqZC
HaAFJY5r6aKa7CTSnozZeMkadWDwFi5My08x3QxVuFbyM03fw9m79rAI5yJ8EieZ6+WKk7yVZkUt
jVT6x9/pU+2BB2Wuz2kTpV43GB966tu/53D0G22JmfsfpR3XjfZvYDsyNSe3qTYti4RG4KNdbjzO
8gZf3l54jrY8wVMrhdBKTO7RgvfEnPTbNiSl5C+c0rfmcAk6fhmvYjVqcN5nTTuNwKBTtBp7mDHx
Y7JOux9d2muXd88jvDqq6yRgMXL/majRmaDnsjpSnE7B5/999k/ctT5Ow7RqVhfkGbx6E2Tra+tM
As6S8l/wAji4hq+eXWSgrGtnAOLO3mQfI5wfZTV1XsnqrnPdWrX/O+OILNvbv5y3jNQeRf+L4F2b
4Ub7k7ThbXMqtSHiDiaVZRmaoyAtEhqDd2saDDA9TtD9LHR7ncRzqQFYHRVEGdi1q68HqHOmmDuA
R7dwHtq88ZE6hPFF5E6bB5+El9lyYZw8UOX7KOUWK9iPbrsa49cVwg7fOpijObOTjMFx1qO8aQKt
GKHz/xgmK0h5wouU1mWTyTt11IlEYgfNrd3PcjQdzNcVT8wCFJb2AFu+rP/52YImNN+fm5zVcU0t
C2V4ECkUUIungveoaeNcFcoAHpjMGHKycr5aehcP+vV2AwoOyUkI9Tf5+zyxgy9ONkpEOjBmRbkv
2soSvcxZ/oUmLIA3m6XvPxrXBvvWmytsbnWOVBkpkDFL6OsN/0RvVb222Fa7Kpdenzc3676KntHZ
bzVAasTET27XZm5dSDJGikp8UCJqHuxQOzncfFLZsyHYi2uV2iHP8wOnEfXpBkQXnj7t8wP+1ShB
hVy1orFUfndfQ3Z72/wDaYKZkFHsX5a5Yjw/DkvlnTv+hMkzDjQl7iqdm1XzniQVOF3WivfnQiqF
LuD0P7qwWIyRND5dUwbanQAiVysARuRV7a6f8UgEc9XC3vrOLD+9rrbqEUIf2AGL7aZR+KcJKLRU
4VbFmcszrQyTB8vzfyU8u3ODLPp2NuD0A2Hj1bXnIs+NNcYyt4AW61p1KgaD3IiO4eRkDphyXoKa
nHE392hyJY8Zi8sKIsaPEf3wmq7C5gkXjfjcaFbRJHEGmZdJLbZtDpayQWpXpn5jOBx5F71w/YyK
4NgHT1y4RoDFemJnwO8scJwfi1v+LP1/+sjGJFEzmc3V2xeqrAgTwpRi1yk+nk7OPEJQseppqMLg
dCOFLIaN4T1P3rPZWVjGKK2qJogkQlRHaZRp1QjUI7jc9SJOST8c9vbh5uiGBPTuNzu+foLjtF+s
SneDz4d/ZQo5bQIymSihfUmeCtuP3T0bMFUQXtAqbCD03R3ib4Bjp9hV//HkGvPRVdYBYnCciity
GAFabv8eI/llgQuKGJcntZEEpBa4Fy09ZjvnGP82pUBV+BIvUDIbkfdCDJ4m/d5nX/y/pp8/FBNj
cojbMxpaQN++FjxLnYRrPrtfKnW7Oc1MK2Hk2e1a5+ExiKXtsvonbFGI4WebQe3D0uOym5aqx4je
KRxyR1tRq2zEqfvsFwCXFEuagLCQ5gYZo86NPNiLaLZY+9cyvsQa8V+PZcDp6gDWwrf8kqpvZFit
rxcF9bnyrs71Zcl9TEHVn+rPLO4dE9KXCHTE+lU/T9RAJJG4TwdoaHcL/XsJQyJmVopvJxJdgL2A
0x4Mbhzql1RXHDn8TaVQnYTGv+M7/ppAR2GM9n4b2dHHT1TLjNCM6CjSPmRedmEQ4/0Cf4+BudSA
6Yi5DBaQhaA7S7nQe6i1KxT1HJPPuTbJnaJ4bXVeiKhErh2zATajDiuJMp/8Zeb+XGhhH0e7L8df
/RrYRvawRan+f33hFj67PdgWkD2DzrXQOTlheI3nJ2L3Y7CyWT84eDsXDk9GTfrAPuQa9vdwSNB/
iHNt48EREGG4xVEzaOHDO81aFWg0jD2ODr2nnhZFx0PaCLY4pR0yrRvoqNfSx8ubzldPUjNmKili
v8jW4KCUavcXwp6dobxPNkeixZr5cMGWoDSrGujTJ5hVZfL1rwTP0axZ0uc9a0Ql6Svcveitt5wo
b1xi36nzZkCaIA4Z81XCaT3hIswSIqnoCCf0+fR91ITnNIvDqaNOCkmZ34QjehgKg7jx1ew01XuS
9fGv14oGXyIUbiZYCJKDc+0STbo+K6As1mq03qb9ruZ69ai3OfuTQw2k1WW9b9IwGdqY87nL0XYf
zan9WSpL0VC9BaTAbUT2+LBVV5T/QyKajb6Q90X6mxcO42Z219zqTq5ALY7a9QeO8xCLa2zjIhLw
D9hwTybGSylqwKw7xUGncJuHkHXrGgDDUuHMgnWR8gEDYchVntmhdUL8/fkGxf0XK7xWHSw7r/A5
wgIugyZPr1gpnoEuYSDFxfQM6etR91XrdB+AkPx6iM2EfL5miBGKCpnP4O6zyRqeCnPSqpya/mK2
iRsId7YYjZzFf3Kye2SVMtA8ErZNMlWPjto54N8g2gksaaU5P5e0+bQvBQaJkg9k9djWPQlamdra
x19noRTKwFP+on8ieD4oTGyTrMGoFAiunWKsnMwxVFRHJJgEOxRNLi32K9cck6DU5qNQybLsr+2n
DZo293qml1dgs4Fg7PNZRiCw6U5M2SmPh6h7JPm598lJHHHPp1FtsT+aKMi60urtCZE7bMLuVV8n
V4/uZyw+AUj/C7BzWq9y7Gv3lWLolbb9wAaX6m0e9eCmlib6AlKTpaXAMG3ZZM45In1imlY+jNnD
hpj2QqPzOlqqA3JvTUWkRgcVyYf9iZ+pVH4zO6WDOVMJrOVcOL4R4QpgLbKHOugWhwObUapYq5DK
OxR4TpqqEbaW2vxdJ4+i067CooqOrVdud3qTlHaS7ghpjClOonq1Q/S8eKWLV4mSBzVypN6douPF
K8vebsfrXs7z/ejzAfPWUGL8y9gQ2QC7ype8KI4llTjkzuYlgd2kLC/oskjbvRKgGzN12/snu/R3
XRmRWS+7UI2CrugttQ4aN2rl1t3FRCN80kWU9+/ATLGE6uIpkYAO/jUt6dYECCRSH+WXV78ZiWxI
eK7DfLwdkmcUFIARM3ucnFDPXBbADAI4QytchDlui1PtKa3e4OXEKsKjook6aQ0DTosfxUQ42KEg
spbL2n2EtqcvPwCql98Qbc9rN3r0U9qnQwb6OJ2ZVmUhkKfigJmfqJR8Kt4BHV0xMuzD9cjNo0TU
gT5g8myCBAQezOLrI/Fe6+9cwf67vHDP00JsIQR7dXk6269t0mu3ZXb0xj1uMbU+sLp4ShEozNZ7
9aE8KNzw7es2JcsGbqqzfI9Y6xrJK+5O0mny/9GhG4h9TH8HlEnYHQBxENNBvYF82UJoKd3R/ku8
9lQA2AKu4r77Q/ASgRcs7zh5jXmK7FoEsZpw6Nl1LoCPlk+xbjNKzhKafomFRT8VCF/OUPsDFG35
LfMx3OctN0J+gCu9AIYHxrLfSiyPwbgX/wGc5Jta572KaSqoTSROP1zzIVsLzCQfQIMNFNLmWLWq
KKJNlbHZHjpgfh/VO5vuAccnzJZxyC2KoNCw6q4sDvWtF7yAH+flrFChoDG4fSD0vyLq8DzGeuaR
Xu9ESE/kTiAG4PtFMdCRM8Ahzd7siosf5ZWfXAHvR8eU3qFv75VbmBrTVPcOhknuKHT+ob5uQoCA
TvKU6pHtf/Mv76sFDazgrah0zvRlgZh5WKH+1hvqnySoXLyBTP0eNnzYu322QOalltrqyc/N+L1C
ngdbp9Rqs+b7RqyBAyAicFHfuSQR3wy3gzqc87hDAUN0MZQ8VxfJ8rLM0E/V20n2VSc9hjfjXfkm
ycb3wMbR7bjKyA0BxvHIUh8rL2ndTeCXl2qFVG5MiNZ/Tf7d2TqqwLW1ZwwitSXZPMec/yxaIh6g
MrJVjyhs/eTAVsyjJHx6e0jyHTprA07qeZ+SfXR72Caq3Os1tt7Ryy4X20rv7s1ctxxCwnj1fotr
KMfRruUG3RvfND47Vk5XBOaPVHN76J/zZ2F01eKY5BfqLo0aGo3OFDpsvrNICujpwBKHy5GM/7P8
ZobJIAZeXbHZRP1APmkCTEw3SbdRe7adHvxbaBkDrZLEnHyRunXTVYzB2OfsLqb7mM4qLfxkBdXU
8lzh/WJGUWx/xHwLjSVnhaB2qIZIBEYQAaC4uKupkDHxYvdXmVmLJrw3YXJ2OYGXkyn1xU+YVarj
471ymvIJdkwH3HwNrDbq9BgGn5UfQf28F0Uy3IEpK0VILu+uSNsOT1QUbXFqwTZB8tnaST1x34sQ
Nlnmjq6F1JCk9rhKYmddlGWkJsPWoBb3xJXS8tbRcYN9y6Ay1HnE50bFkspKLFS0iveULuX9idcO
kBWim7E04HohPSqGpIJHn2BaqM4NttmEHtVJqEO6Ze7+UCjFrxJbNynkhfHcSkcxH5Lk55a+axg0
pJUhflHV1NRFgDnnsiiQFSiAcAvYui59K1Amj+M/dETNweGOcRz5OvNQpSxfWibV3gRzwgXTfrbH
EFSfy65N/GV+RTivKaRaD8SvK8HZDWpb6wTCIlBsR6ua+GVTqOR/kEmdcD6A0e3TpEQQSjJW6ksl
of18TjZ0Pfdjf1tnWBce+J/2/mIT6WjJGntAJy40EjA8bR0qvukFd+Q4JFHd24+jMembXgcZ5oH7
dxOplu4NUymujiM+KDz8Tn8TYBZmqFiPKjR+I5zrxogiSNoD+1j0kXNOJoZtXRF8qhPCV7cOC9pK
0fiVpaI9f3uHpFYhXDXkIWcb3UilPmkRi6rFCWtrJOMT7Ox4hDujFAF0eYIxMh6k8WN0FWDIP1OX
ixRC8nLgSEw3FpzaxARq778JmPHEcBaRq4GWpDsDWSexerWtXVoAORBNjmNmQNEPxunmXuugE8WR
COWjYz+gw6S5S7Xb+pI93cHIwV5Cq7Ndph5SkHObrjVV9yUEjP73MCiS9qfCWsjq+m1ZZXPyfoGb
6sYmCGY1e4jimgcfaZXq/TYFD2rEVZt7zg+37ljPT6JxBJBIalmHprBzHi7kbXf4T1RcjgOlwcNL
Begy1J1TR5jW4qsiliXxXnACYB4dpNeStzNhtSMht4g+K84nFf7tATPX6NtWdSI+gQFShHSEtaCv
0i8Xf1NbVa3v14vZsGcI1NA7Vue9PHYHcjUEQ55QBAjaiT2UsSYkgzq5QxLgt4hZlzSRknzPuoTK
uYdjyKaHpvA7EFQcRtgJUgtz4pnZAaDn0xemfEWOrHJ+Yz3IIz9gcmZdgGY74ZFP0LhDWHthfpPW
zbzqQOMuOqWWcFlLdC+5CvRFx6xGKCbRurRiYmCH65QWLLpRxzsGgAyGcVg2v629+Z4mVXsNDsrC
+P4FCt4kdAHbxNJjnbTkSZ6UhGjwNjDb3FADIqgQY8yZq6E2eJfQBrNPxW/y0GEWtaJHlPaGqk0c
F5K0zS7d//PMuABQH/TLYQ1KB8gaGQcZuumz/aGGdwWTaAcgxsE76Wd7A2gT50lFgASqdfy9TpyE
5coKB0g+tU52MjMbnWVttG99pjAdK78rHbmuFdibgSJ1EJJFp3+HI5D70sQJr9E4ljQLtNa1yMbT
rKlweYZR3cbAI/V+doAFD+ZZ+Wta/uzNj6sFePHsRF8WIJN7zijttLREKJ3TN7tMlh6mFLHw5Vpv
Lx7Iw0Q8HGzzxld77CUtU8HH/1Ec6LanCDX6owSH+zxE/eB9GVmnBeWyRp4oCgjcLlNhipozcW5d
PM/r503rEnAxVR00rtBvws8LttlQ4kw2E2J8djavxw4wOL8Z/yzMxirJ29PYfxt8irIWm1nICthf
4FAeKI40yVG5m9Qfxy35vtJVpo/lx+hNWGkNukwddHLfQT36sdQY7JwMtaiOLu3QqlXOq4uDn8JZ
hTtuP2goJZSS1gmDIJBGxkXACl5ovprkeRPbjoFzLeL2DDwgv4akJVChxEZUqBUiRx3/LxtrF43j
Q9yGB+B+LyQ3Xq0VVArGMVcQRxifLuxh+vjflS7V9oNzxFJu7VlhQTfSR8ewKNP8+7c9oWvuxVSQ
Pky0BNdO2wbvAKLEMrr/zK43WmfW6X1MIp+dcgQLwIUBXzrv2sN1WIGQ3dk+dHIqSorwL81JStGa
HOHGWMchiT64hRAcfGaTGMP9nKcvsCQsBN7OjapKJVx183U+SF/Gd9pUmGc+7sUkoI69zBJlBi1F
PkyO8ratlL357r3UHRooczMlwXcOr9neSjAxV2y1q+vpwXxICvTBixsWzK+QjEuUeu5YQexmgKvw
LgVndpnMCHN2xAr/rrzDoQbSPq87x1vldAThgVVFBhgLIvWb/kr4q0yWtwmSQrKixkF/gEv27pf2
1ztA5bY52FoTjm2aAEzO3lXYg2399SKm2/QSFhkEbAJNH48xWjEioSJYfyOIiwI1pVpZ9elrOkSh
fTAHqX7t/ScONZN7gCPr0nivQ2H9lTeEy260FzRxaWZghKPNaiR41IEHhzZaUe+f1Z+NNVE4aDcj
QZn2fFhXtZgVppMt2/M3E7a0YFceS5fCR90L8oCzEuQx6jOWe9Eo01ZAA6/oJhTQOd3HdctqIN2o
nfhIPNhaDwN055WKdqL+8X3Yf2eWxqxANPXngnFq/piRO4zKdcdjr/DtDAJHepoDtt0H4cM+SMIl
3ykBCwUCtjjJ/Dug0ibfu0hSBq53EX8GtpEg6/t+Ct17lKzZxp218RmCBkb/1vuhXfRFzVHyfk4F
hs5Kc9C1FwLuV35szR94n2uRqRZ1A/kP0+qNxl5CL0YPq6krMm6ZtHYBE902O+byKXCS9m4U9VkT
RLBJAkA199BzxF3N/6fvFa2LAE5QfZ27aWw5o/Df28TxQN81oKMryP2lEJsdVgRNYPuDUJJi8Cxh
F7WpmlIyV/5VUQAUw/cJ680uUsYHA7GZVsT3QnRDlz2u0t/5zxe8LFM0P5aAot4PINYZy6AuSMVc
jV0W7+W2b+WNyApJDao1BmfMMGVjQAeTb+JQiGtyQ2yl4xYSBQjSDpTrIuEaS+ZZ1q7eqxutFW3N
uq4tAkfQ1Sg3lqNiRBZPkQ7pRAjtJeVFgjPYburKlHl4Z6uJLswg8ej+ALDg0GLcmR4cy74QmAm2
KSzFYeIUUq4kK+B+6rD8Rw6f799iSrsfJHP/Ysx/gqb0ahTjPR2o2u/mKpe9nJMdKAcDEc/oSMbu
/q8a2j8+Kmd3/yjuYPXKlZPwCv/6Z6/+50I9vQzvMgeVenadZG88uV7CNq6TZZVfrJmTznTX/ESq
E+Tm2b9MDz0Wd+e6gYAS5BF3gOP5YUauzUlLeE9nr1CFJLaTWwBHF+7MWXtwZrQ81XqoUmLDs4Bo
mE4hhe/jCJTPHgCm0cDJ9BaBC6d1iH5Kl92EQKbNEZIKlNBCtjR2yqgFl+PqSE/fCD7LK1qKjL9h
kuDKJK4QGFTkr3vV518thWjnQ1c2if0L5GVFiA4dJuY5D7LeG4vtrQHBZjN3yk/WXy/RlfwxxCHl
pnIPiDHgzwJpJyndfw2G3SIfrZlzGoNTp0wUojMwt28HDhMyRZlBKaZiYN2PrM/RUzohrYFV4FeT
ivzMm7GaS/vXJzMBqHmybhVkwt2AcFxhXXdVYa5ErFeqTF67i4mPFDIb11UF3a5r3zWf224zsq/V
79RAzEPyPXC5og4b5cZoS2rNtKk85J9Uw1A8K03yMaG3ksOf6gHhrWxURa0srYNf5Sbd4s78PtB6
9QbCb8M1V0yEseLzgBrn9gR0Gy7oJbo2LhhbQRG0uMY/Fa75Liii1GNKuRSJELVBvjfv2+7zRgM0
89IQ++SRbbVwx1fooE41YY5ijW6g7Sm1eFSrcR23QcxNKaxWW9PZMSJWyVWsluDQlb/IHKQxgC4N
YmRkqnTUM6zsTa0FQ2t5Gn2kGUBjj2LAQmHyNlg1bupqn/enTU6zNi2gIxwZRr4lL5mGeJtczPPP
H5PGPKWRgF9l92EA9NL74ZRl6tRteECNz7GFDpu5Da+uSY7OwZIKP4kQjzsdqFi8sGWM7BHM9Tp6
+t6AGXNj6Yljdykp6O600+zQWrGIMNK9od6OajJ5BpeISqC6KACAR6DDqsRFsiA6osr/B8Cg3fdD
k3BDw+D6CQxPQvIdYKyShoPMpDPocGL4I90W35NoX5Yemm1HdZld5kPKsBcxGmQPhG9zoTxZ7qp1
lwpL6hMXe3KmDUy8FR3kvw0nxX5WTBAwa3lDuF1nILa48o3Tr/qJd7pL/tU/lgnZ/dv98uZyBkCT
DDqLSZkKpiZQlv59crSiFT9knMh42/cqLL7oJj6VT8JgsQ1m4vCbf37wUcCu2oV4gBLy6uwtwhc0
VTtWOGjpMZ0uTLXyolZRtHIwsK/K3doBiOgofzrnjTYXit7grdXc/4lZJGtUzsB5BmvamQsDy7iw
KR0OX7rdQF8/76i++Zk++CqeaMTyUVpByx18qkyZmU0+7v41InUK2j4/1oWJ1sIjxkn/qXJ+kzgF
jOJdTLtGwcmGgRvojGVBaouPwD1OBxS06aShN0KSdNxPNaifKUOe4oyA5rO+/61ZyyUoBfReaejj
2sYrbAWwTdTS6mg1/l/JAZorve6OQRJitvGMWo+6eE8y8l/OTOVOcD3meTHgqzjoBFKtVc1zAS35
jGoAMruOHUmUSACEYh9L47BBulZlP2KGpPqJDph2XW6RayOclo8v976/9acPVlnzt4g+fC4POIhC
ghVTV7cImHylfjuQduZhY0PjyDdtbjNis3Gbxma0GtidHJGyQ27UlC8ki+D65URqwTnJNC02wJPZ
CiWqhzxJlqCCucS+/jVw7CHZijbAVPEzMo8WEbPxHrBxwlSx37GhlsMZagkeDPrN+aenTN+OdM9O
+U4jLuXHxJowA71UzK5bbu1aFU1INBt46d2fGcDTxxldad7wi3rsO815eMtYke9zFAtqIK1nAHTn
3Bkbi4wRg6jA5jMz3EpU3mtnwgjUuDXNY5Ao6dBrmUpEu4C5Zrtj6l8oTb8W7fwYC8olqoqYK5wL
2wgkpfpiKospF3+G7Wx5Ttw2PKwCfhJyIFfnnBWtmeDa6TXTdENAYVd1/1MHJTTjkBvQ2uuHOGTl
pSfBMxF1w7WkT03kmo+TOOTsHAKgmuAUmv+nrcY0U+OPTU61kOZXFe58zI4ht3bVZNjQdgR0ESbi
k/6tmjbXmsRa1jmAfNZek/pYdHbIgGztGOwxVvmcG6zKqL3wyVk7gCC+BiUUUolOdiEj54+irFu5
cwUOX65bq0eEJDfPauFis+1/e5KM4XDx5lCzO+iSXfiGZbJuhlwxP86GyBE+3uIEfMax570GKFqh
N3LUtYTIi4VUQBtsF+EuFr+XmS8vEoh/FIgdXpbFqbZbc2U30F8KI8a15VHCzOHC1OqMoRWtcdvr
orKixhKmKj+S5je/AEQxGFBdIsXeBgG+C3qxXDwUVOSOdb5Q+Ek0mSVveFEN138aFSqKTLWjqg+T
P4dxOZlvnKRS8mYZ3gfQ9ziF+kYcu/Db23ZkMPHFnEFsHWz6qHeZiujgDXcaHCeInBlwD9ELsu4Y
x5VY5VWw9NDTBD45FeYrXjOxWuSZ4b395uO/+GcJdb6j8GwRrnYuVkfH6A0St/Xl59jpQOjf+7im
7GAqzRVzuZdU//DvrcpuIaoxh1LEXxQ41CSkXV5rEfX2B8++KLKNr/82y6qRHKyOzZ/bIQsqjV3+
FmRFLm40lwlarLVgOY6mVVNYAJeEw88ZMYmIhTeVPSxBe27rnbIFUDfCbWInIOlJZRmTsdHDoiZ+
IQ+Lr0JEK7Dx/mumfSmO+7KSGW6plXnnQNC3k5ys9Xmuwgjp9PyhFZQkjEmW7ZmYI/Bi0De0yXDi
/RgB9eb1qmIHA5EDG21oIrR0arFMNFO4CzhTaYVvXmwBy8jnVSaKGCFbpLFlI9alg1P9z5o+hEFw
KmlZ1ddCl9QLDO9YFz6D3i52H1uFZJt5S+eGGYyD1eF3qsyuQk3UR5XGP7p4ba+pmeDKr3lCthtm
UV+L2ya297svfEuly3IM3HqOu/zyqORL7DPLzZNQE/sfOozfcLwlzASrVmdbACPR7FCJaUocun34
anfL3qdlZK9lrhJyNaQ93HbkkPvdAIrDhwdKqRDmOSizPmqJz+Dl50V/ECOASc8Wtf3KHy3pr6Rx
D5SH8UKu7xQeJipRrw4Q6bJIyq9qXuDhAz4y/imttoe/HBGyzXF3JIP+bW46Xodb1rkSIsT6RfF/
6GVK/bvSGVFQ6Aoroi2EuNiTlZcW7tRhw75wMIrggzkhutn+RzwfD1H8/a6/+nkgy12cry87J2B0
+DyG67fkYnHesuN4PuxTSqOBjCr2DnuTWQHgpp1ElrHGSZUyl8ADy6lkXxmlJU8gUDkPAbyMDWSG
S2ESSY0ov2X6Y97zDbItUY9/gI/HiEaHi5hfZ6LsDZoQn5sjY79g/jbc0i22lUO+vyr5/u5+Da2q
pzOHTVxipJ1lpLJLNEbEnusL8vWMqUTPpqf54mwac413cbE2g/3Ji/svCt7ES3BVmJN030xEiC1m
+FYF2/g3Z6XfZbXSmKHXVon8BRsVl1GAIwuHG0+FYFKQnsbohFifD8NwpFP/JCHa+lZwHnQAyRmy
f3tECvR/RKRitfw/5YJ4di1tY0flx9ntWSYFQ+TYhEO/ZhxudEjwWNXUkktPSS2pChE3XVriA4lV
cLkpoSqxT2SDKVQan+SCVa8UlYJZON+pitggTU137iilZdojNq6KhErL0YdzmYTFPqxp1pzkACi2
/5Jf+IHEXhCUGkf4fF4nAQ24y0BD6cINYpjlSCV043edyDY9mvZ3SZ20rYFqMKQvCtodwr0kmaFX
2N/mD9YPLKASVoYLY8VBN0HzEJkIBPe2VUo8LgwtdhEjhPGWhEMWRXydYGXp3xzBKhT0q6RDuiXX
XTHjScy77Bpyk7FHeE2OdYOsbP0DK/uZ3ZKkm/KzuY/GJSA3aibl4wFr1aJEir4ZDGSDZrn5zfMT
Xb0c6poFGO/qtPviRF1Eqko7H+KPx7LcBuzkeqgGR+H2g9CSc/Rwz7okqDxJeIAKU7X9mFL7DIUC
6PgTO5ORJ5gcxdVlNhbuiMIjl2rYwPR7t3ZxNAlknUdet5hvoLmTnkliYwYHovQptmQq8LMu4ZRS
EUE6oSkcr0+lyok00CK7r38gOOAf1idAWzgyRMrBDvHGdLoYDV/WRrZZZfEjn9Yqm+nPdIa3dVq8
7pVPsutsSeGdMsMnlQPVe4v9BBPnX7mUtywyA2jDfMUmW0sqlH3sp4imCrwc6WRiXXVvvtyyqGIB
aezUImY8DVQeFA0IOWzBZVZJU6KOMZwdOzk/Q3VgEzDsXrhbrqt1ZCeAwe+87zhFKlNpCrWhwfLV
1jBXIe9cIsXEt1ZKRlPQnuOsk7prBHpRtsAqHO0SMFv5KFdb2GtR7dt3gz6gao3XTtcL97tTz8X/
765UCo+aBVypoOhMUa2LcZfvDA9/4bJd9Xh8T/lrdGRuaFXevbPcwBt7gYmOEn1OSY2vqX1Olx3R
08MbLaovL67Ma5Att8XuEPbpPklKbdYWk3NVbMsxzUpx62jCS63I3PgzWa3//Qrb4H6qifeheTmR
SYt1hlhRZG4Ew5DQUS2NQqOmrmq/+VNq/JKJKHm7XzWyQDBLlljTt4ImLzLYmlm6PNE/538xh6MW
RuG5qSxMkoQMI6UivWpOdCrLwtd1J6zbDQI+ivkbha5d04vlSPQqZVLuLpkzDETd+69XKo5UBH7j
5PfK+s9dnX8n827G2y3mU3FLfxG58nxoVEKpysvUv2DMGzNoTQLbEba1nuP5sFWdNWtQ5MOimDII
Kacgmmv8GAmApNq6MTP9d4nxsMxVcGc009xaGrj8108JAAevTWkpfiYtzBt0dW6RPNoYUXHk+GjN
ZSUmFdX5gX3fHoRXAIpMnIdYff23iV9lhM0rLyDYQhWER68K+7AgBIfI5Sgn2rSDt3A9IDlpb0AH
5JY5n6ZxHJasQ4GO9LbtXVl2JG8X3IRI1pjihYzMPG+CZZf/W3CelAsDCPHuPHuA7XT2oOg1rGVS
8H2QihMGP8rIa1Qb8bmtQXtMYrAQPn1W1kd2h7GN4YhE+3n3T9NRyETQELwsm855TARjZcOswVK5
hko9OFqn/3EWkClHKkCsOtxjR4wcoNAFd9zzJg5G0RjUaIMidirTG0mAYIlkfR5E+Xo0XwMG+yye
mGxxwMYNAumgIJJ3ZJb2TRNyb+v40Qk5flyMwoh866wP01VfHaAks9/cOo32Eu5Bnidpc6Y+mvlj
skXURS3Ud/eLiZjIHUnhhOeLNnxuVvprwMpWm1+BDSIJDs82/as4RPg0aqdobB9vIKY0vWTdi5qV
wW7YuywFSQsF+APUEaMdTj980lYrPcW8TmQ6dhj5sm2c5IUThUZaMgyzJfhj4+04OgIiLSYGnvrP
dibQVlpv4NGYUosHGHvdrkraSvGEnSxhy9nMiWPdpfqk3Mz/q4FHZkph1ZDXPzGaPFb3EPf33NDW
aRxNUEt6WEuV0yzXt6opYyxNr5kF3NjwM0hpLdVL5zyEtzQbjYZ9PlzBAPwOsm1bqoapZckkMRiU
Nu0R15Jd3zhJwHjxiUp1c0pp2OTiV475TC2nf4BnAH3P/1rb7kYfM/F2Una9DwaeYZQiwjIg3lm9
A75c36HUBo83/HvkcsZD9X7PjDh74D6AOFcLd9qEUk4neYtV9q+5KDYePiCDyEgAB5UPJAQdVNG2
PPVqKmOzHtPjN8H7iTM79ENtouU+IPijziKlbRdVlAbLLBJNzUQiOjH5hNk34DR2VZialIVNINGY
XvY5ZGHzMqAwwt51w5XxB/Y2bvW0UzPTKIcvb3Lr2uMS66UvdMSYrxmE0oYQXb0Um2tqbmXJf7uI
u6H6Q7vokzakJIqbdAsvXFaAn85DikfAZDgv/7K/M9EhtFBUWQDVllppbbCVCnQ95IfpjpFDIwoq
Bck7PLLUuYhwONIuBUC4xSh09db7Yy7+1fYgyF6VTexUxRUVnDnls54Tx6W/dQqAjUyB5MlNi7RZ
Ifv9je+uRb4qGY5YhU725YemjlMxwTm2m5creXf1L4TKTW19PbHUs0Qy3UlHfbt5r54+rNkBfXyM
7SAseuomM8pWThYspv8R5scaO1C9kP8APfhUDHFRYI80ScTL6sZM0pXjKXJYD3BAab8IZGX92zdt
C8zaJlFX0iEnfIZT6iFleWNkVFFZ5+od2WuT1q0ZKFBXPBdr08NNq+CiCoRGXADyvIYIhbwJ9ceb
A2X+U3d1OE2GavD0fqsQOiCO6z5OEwzrp3cNKgAvnIo7zNPQkEKk/4ASv7fFDObNAfyXpuGeoHk8
smLtuEJe8DIczOj0JDBu6SGnSRoQRpbqoJIG7uJJ4y3ifbE4SEcdlOQpFdVVlJjsOYZPcNRRpcvy
dGLxAnedoW8VYkViX5N5nLJUYbnHFOZxtOkWopHofHJiXM0cvEPkU1iEJb2gOoo2xosBcUtXSZ7g
vEaZBZKTG+090H/nRTQKe29UWqSXQiUW6rryQt5GrXkuHOTqVdqGg7e0CrhMLDUrX2dEoFfnKFJM
tquiDGMv6AAa5Zx1UkscqB4aS2MkYKEvRgd3lZzEQX8SbgOyGo1O4nc8iW4cxjSUyzhbS+eyV7RR
YE95FZRR7xMdk9osGVhrH8+8HtziMFwjazn+g+cFcGy4mOm7uvCKgZSKYgJ7RBlRggFtVh+WZsDx
7xNf7K5yNeUIz6aLlsOJCZhocF0FqwTJRkXXFX3s6Stvl571ZrlDq/hN+kdl/X/iN+boPm0CmREW
87zzL/y6FY61FlDmbEzn2jYswFjaf94LLnwsEdpNGrpahbPPsVMpzOV7w3tcZmyWmq32cG/7ll1/
C7v09DB2w1ES+V9lkrGp4/FFCrZx9eaiipoqJzmIYxlwicoAMUww4i0TFiLGZ31IF1OLNhhGIIYk
0GY9P2ofa/m/TQS1t73vKu5bRajm1eJIFd+D7G2Ybri7xRDZrfgX6bVdCEM9f3SWeQH22yNFR/PF
rK0ZQrwoYr+bS5azGMtStgeFw+orDtS03eHhObYBWz+C7MtAgqVdCa/M23zom90T/XfaE1DnMRT7
o/BSaplR3Wol3mMPwSrhZFRWUQ64NjOR9vUZPRfQzPsSSrjSSzzBGQJbXK0k4NjEUWdKFpYHZFn7
4E0USksjfMc5MODBLk0DREA8JIsR+GPetF4fXf1PgGYNK7xp6QdyTt+xqI0WJ+41GUkF4h5Ws3R4
4R0pUXy1EM//XC3XUWe5hKU679MJ6+icoXNNQC+eNrPMIN/UTIZHymGHdR+3zLwWn3vFf2GEdFYH
MzG5xHG3kTfTDLPPswM+HphVTQUTqNJVCtRneV2cEkU1aKSGWe7M4YSJbIkC8QrwDkq9br10kr2g
7GGvsMjp9x69+olEgpvPYFgxWwPj1OXUpcOG1hZHVfiEpd9iJx/YOC+1Joufmqq/e9fOtclmEqJC
3pmyzBhSP9t9DxH5oX3m6q03wCqWxXr2D0NcMUwYjOEQ84zMOYliZOGs+PkAJwnzwMaxF7xD6Ptt
Ie+Hz+oVzy6zpe/lWQT7XAoedgJqIrN3R1/AzCTgRYHT3Zm2nQ3nGQqnQ34vbgW+LhYZSsbVLiZa
/pJTHghlysscmrkGe60g4jONZxmLpVmHFKA8gWkmTDOTMKVggkurntGOltsJn+SoEb9iUOX6j5t2
pDFcLLcAXXkFt2fkVR2o2hHe7eqpdNVxd8jixyzwK5eYuo7Jxu2vjnN9yonu80HCKU7Mb1vClcqi
9O44P3oAE0y/HSs0rt3hO20R9fXlkUMgaIxEf1NRnEF2mZWToCKDKqKDpe3Jy/7j3vGQr4/WH+RW
7ZECVMHVvz7bx2xH0YvS2YorrtNDmVY9EBginICj5nD6KZ6hrrkBCP0RMuyHqmjyRYSdnj1MUNjP
+vMC65le3izTQihDywjJP5P62RJmSAPaHkUVv6KfbuvXW4M9Gdy6dY3CUsOv+WUkiCVhpTWZvbOG
KM4kY/lKQ3SiItaHM+aLaDgNLHAnAYfKRebZFgXFl/52Ymfar8eEgE1bR/WC1GSE4ORjf5KZ0xF6
ApQpsKrQXl+dlJeW42WT+oU2dcTNl4eHIMWJp+GOE5r+sNXVJTc750z9fStx+ePY3j9YXgCTJAKX
kSb+vzJE2n0jjcy05t4JEjVYi6IY/eM6uuloZoKipmQswbjBZnErwWoLTMiRGH0qGJPqCctNYLBH
XqyPEXdYN58QoqxRVyI3nJOAQYFJ+S0aJy5nlaXkcoWdUJnDTs3oUbTwJN0FniVmguRPqUaYO6vy
xdSk8PFFI1ebPqHcAZkuFUPf+9rzcqOYNnzMLWi47iXhD5qW762hxolqCRD2m5gmEpWkBc/SajGF
8euEuFUesdBs54ih1pO5DQxzvPYy4OLR9+W1EoOZpo6/XgLwLJCkTnHMW0IvvW5mjIZ7rurdT5U5
cXY3a8OVConU9g0uUtLn6Wf+sdPkKfHBtr86unmMlGFs7h5bs7De4/H7dhAQRvi/l8BV+q6/V34+
B6erdvmbV2uvqBN4s6YPmgxG/Ws5KUgcisPNNqogQ4EbScVAHoJGVPMx3iHSXB93ATFA72lwJ5jp
7WnU8D5tzBLcl1PHE1jN+nMUasGb7mO4P/YshbLazbNDBFr0DMdaufPrjq+GiRJRf2Rc4dkVsSdo
uTs3bcyXe+qpbCumGzA9HEBzd0YFscOZozwiFSMXozIm5qOHxe5kncgPPW+PQz8KCtOQ/F2PNIJm
37WXzow56LTHg/VAdqwhLhqV2g+wnDlWsSH4gRPFdUNnObwZj1Zt6mERQ21pkm8CrBc4eBlYni7l
R++SYKNxQwM8qR3FlTUzSWaWVV3b4a+fS9hAox9HQ62tsRa/MM0rGZO76SNA2LPB6IRRaf7yGRJy
R89vUuUCvoCHBmVYYcmwSN4M+0uDPGoRoXJI8+03ckNNOAwJVb/cAqGUdDIeTVBl1zVpYPDYxH9G
8cayXJBgF8KhQ3sSd7g4maO19qGROcQdbCAnhlBQ3Lozdua1jb2oH3Qc2Eyz7F4eRAa9/PsiNt+a
cdl9UBudx5xrbh2Iyp4ZWzcz8/8KQWtW780R0xHIa5G1/nbYEXIOuiSdx3HqoXgzFKcnNdMoO7S2
gRuTAIPS88+fnM6+oSu+WB3sbir4O+/cvjdlOb+JV8RcWMiOuva4A3kcZFBQZxZ/tYI7e6n9KVNp
GcmX5RW9e+0ncr6WTo/T3pvXqDzUgje74XPMv9J5PCM7bjVcl1JeZ8ereRnzNMpL2AUQoR0waz8P
zgwANLrtC76sjbzLtp192DQWq6LzRCBnFlHLSTfuW/DMgT4O2FCjwzpTam4e5AQHC2hD1T2e74bv
vH+q8Y3vzXO8gXKj1EhhuqcEFmCLqY/AW8Fu/820uDuDwS/7VYe3t+14KJnRrpbTbcG7HYBe3odh
V7XpsxSbwDiIzsByR/2eoPugQw8uwySms7QrpIOaHUoULzkJrpgwuQh02wJ0jyaw1r39kfjyPF5+
a4atzaEyElwFPmRyiV81wJEM3nzDCmb8yQKuRH1ZgSnrkVPFR3wp4/+duHJB2lVNlav4OT6owA/Z
ssZp3VTLtQbdJaSSZvmKfsdUHkdxJw5EzQl19UPPUth0/U6KYqdcGorQ63CoxJGQ5AE9dq5WMCHw
Kk8QM9FkHlJDqayrt7Q3YhhkpEMC6mo31kc11NCyrA90h8ZL5IgoWl6ZNUnIAl518NoDJyYmCe/G
inAGNgc4z+eEhfCiE7OCALAR7DiB12KI8HI3457Jirny4A6evY8vqmPY9b9xJ2Kyc6tFKARQHsB2
KBvdEtWrCT/NiSrSiCbA/Cl4QXoyrHKOcQmtoAJka9CHro4pqi3en/BPHcFdOPxB9Nv3xUnswM2b
KvPU+mncgBVoDZNYuoh6w4gXskO5RHbY/3LkMfWVkdVX1/OpaZceR9RSNJfQr9E5pztDvgqIxjEK
YdCJwgy7P+/2ldffMXTbP7ENItbhhKvoJQCOtm/Zo5/IPCXpf5gkQ2bxAMe4qZhxmxmZNuTdvt3R
IcaB6BJqXaGL4TMwuUpRx6doPyKm30yp0yeJZGr1dWtmikwtMzR09F+cYFe9m+JtNn8eQttbeT0y
s1/b70f0xH09DBcmgX5ryZoCZRmXL52Bn3Lsn69vHLVkcWetVNR4TKLt62Q8eMOQl/y/WzOk7JH/
WAKclHxzmSjEWSEZg2/Ax9y3orIb0p5IP5qIy720wm9N49bBoi5kdC0o9kLQAYmWBtJ/CxRwvj7C
8bDn2cZakV3PwhjHnbtvPGCuwn70jXw0LnyXo5Mn6TdG2hS9dCYu7yJr0innccsdRT6AtmEYp1zN
TjwLJ15XgCKC0STO+bDCJUpYte4Wns/AWqaQfpWBd2mg8fjltixpYOSJ+LyhNjnQAorH4/+vwW9H
RKB2VECmT2In6YNU7ssaHzSKVI5a15aonJG7WpjXEqMJJN2qvxwWbe/VnGonbquqkUskYilusgoV
KDDJ4mT4BqybaIZ59jHszh4bWkHwLDBEEgifnScQCItPcCYaJfNMvd8ZJiSaUZsJb/D10sklZd3O
6DriyK2CGG8SCtP9JQcDBbS4P6piuSV6xIZJIEpY/2dNVINI7dY7CuHOjrAVmUXA7Aq8WVwYox3e
FSeNH3VahEglk6MAv/3r+DPkMFX+vsMzDZ9PWgN/8X1xNv0PTbsV/20cjg7KPvBfj1C0qmD/OeVG
CUzO9ayyvtT1hQQLQPtuoPEPQ6G2ix18S5ZqLddtiCmNSPuJGGjNTy25MnGSkb9nBEU16yk26eZU
Bm6LJbdRy4lKad420KUANuTrx49OrxNThGnJ0DAX6f69FLvGirz7NdaV0F1Em11o56H7eTwB2NCe
gzIDevH2Da6KEDdxnrVzsBQKpWRUuZhV2gJEiQDbtAR8EhXEy+x2U3vD3pPHSipOlfPEKpJSowyd
l6K2PbC9Zq6B+V+gkAouvi4NmTZttaShP2yzP0jBJ0mUJeHu0LUZtoeSFDVfsWW8WXVCSvK95nKR
kZZ2CwuoSXiJUgIiR/nRJ9KtYJHZ2dpklzc/IK7rpM5w4H5nsiIBR+isO1S6MOSLZT2Uva3HBqjA
TcNWpBmTHz2wI5lQc4e3dRFPFM7d4os+cmzJvImqOWn2bWujVyeIVnyV1L/gvODoI08d+ASiRZuL
o5lEI/dVGiy2kP55OnsLkXZxFsEW3mEzGrOhxFYgnrXM3FscgFiRiwtMIXQClhP13bVzuFaQR4YQ
hSThZHVksvu0pzXphFQTnUYSffcOD4LzP7cfc/WT5ITRAGehFsQt7DYtXUZBlc3qql8C9FJvzh85
4syu4Fos1ZlywaAk9GpaaW0A6VpFcVwAGQT9Vd0iZVtg6ECLiN+8H4CkjRs8eZQcqJQGsMGQsnVp
ps3DSuMc5zZl+1GqtrjKAiZAgfI8CQ844NpW0KmptfI5JKY7XYwDqW4zHk5Ax+vMxTuGFp6UFZEU
xxIFnul24v4yaUB/lc1vcWX9rxgEx3KLwue78rqJQdNdAXdBPKFfaD9De9Zbw43ZJ+mWWdNn5YDX
loU1KevjYPJOpb6pWY3//vQoidjYBONQDDB9hPHXpJlOPQa+yqR3Rx8j95trjontvwxDmGMyeHdY
hkaybs0stNroGlymsDVDVo6VVRkG8EZv51DONX1qmcfJ7vZ1ucDUZm5IGcq0MOvKAoclywMRs/uh
R1AFPz3QyCBC5oxGh/Sbb3QlYePWdqpZvV1VGwSpuZwdWWPwGejoCDzHlzonrLdhiMAfDgop9nTT
4BPgwTy+e/BuV2UIGrnPld35oY/eCtyTUkGaev+OOVw+TkWrvFisDd09HlO8TGsG63udqk0HdTiG
aRMQtn+Ovo17B+WIWJhXQoHbvi0KlF+BIBtKuafT6jCTxiZHMRmHYsaD7qp/U9nzANhBZDky7fdL
7nTvKWk5eidZwVrnmwPY9A1qfe+gHQGDFHDNrozg9xKSLSreoOzUjSQZfaJhKnB4WAti999XB2PL
c1CWa2N//cy1BCJop+u0frVrNUJyxQ5LPmspryyO68Zu1fqo7TIeVaUSm+DRZG52fv1hS/9TupU3
tpvV+MvbRFRdKBgimLefcDEh/PVMCCgmQnQpSGpjKWLLEAJoFcGxWDBTendqSS55bFo/PMylj4Gd
i/J8FgKn6bWGkz02Lm8R8bpZW7/s7SKL2ce6xZo/aK0OhnA+GL1FlyfZDKeFMv0liqvyK/t5zheS
lOO8NuslIBvA0K8J8N6gyNBXMpHBB25UYBD2zNhjdcPJ6UvhBcFfo0tCbwgT1DqIxNtvtVdqpzx1
5tzXNs/SYfDdYYcynJuvm8g3nbeMRc1EmEOg+24AsZd8broKq8xeaHu+Vd9jd0WV39EEstkFuiSv
fk3Rs4HSkEtTMjucvlFNiSHDWPpHYe/z9q77afVK8znFEm2srU15rDKorhQKz9i/HEHtmKBqituS
NYmc3qDp2NBjzryDUhvzUDVP/wnrAQF4jhd1AoA8TUqp/xr0y6IGC3hpVe06opO7zmDbhB9BGO7Q
KAMvrB12oB1i9eYBytsaJKtpBPYiR44yOKc+Hxbu7Skpk5fpliZqFhoJnnnW2pSSuiCzl7IqNMNu
Aem222VMBtMIbzFgxv3Tq3m22hOTw6TG0a5RJs1VG/sISYy5yiglqKvx+s8+I+rFeRNl+bDPuIaf
x/HiBu+5D8uObfecJRo1lgAnDaX8dTl1e/AAH4xih3nJ1WJplP1ihVqDAafMmpntmVGl2tbZp/eZ
maBEqcxmaGnmr7BeaYtTh3YOjsQQSASSf0L9rRMCLybk0kZDx/ndaBzc/88BjeQfkO89QR26JuQ2
G8eq06pGvG+bwGbSVcatdg62N4UdsYlF+CL9+VLdZWNUxZcL4+iQHJA0fceV49zjQj+o4rTwiPYi
CIFIJ6Xp6vA7L2MfPQHrojZPMg91yFi/e/ucTIgpJlUhTjjkURcNoNyZDM8bOTZ7DccuQO+OkZmq
YA2zTHU8MKYXFsQbMEJAqV6ZNK+yWOShmrC3RskMt7aJR2PPWGFm2bbBkurh2+eH0uydE6eCog0U
Zb/0Y0Wz57svWK37nb63QZ1lJGvcWy/sBBoHweiTVq5MZBy9xcVzfaY7tlWmaRD/8kVbeZEgHEzZ
X/qQ3epBdJ3U1R0f0hJq4Bu9cZUSzkYHoyoV6ZcML83lGHUfrif5y3J2ww1i2lXN6r6x0kVkIAYS
PGoCA2f4BNfvfy6zeN7cJK1CPrTYvlsNWfzcGMizB8ogx3GNokPVc9RrVADsPI/wkjfVcr8Q2Sol
dIdwCIIrZgd8glDt+eNMImENnytQVCHhvMJ8RnIk71so8nJ1962KTV/jK1usL3wQ1cX2kDbZrnPQ
SAsihTziFqV9LwU4XxNzVel6nAcCsBst6xE2kpoUXdW2zMmibq35ZLldPOf5IijvPPHwsDXVMY3c
H2Bhh3a89Q3NrjXpcmx4Q7szQzgtcNPCGRWSM4lLserZoow9IkTMcyAgN8JLg7sD0eWI4RCCASIi
SQHwSe9W4cqwAH3UVdO4ZAvkFA2l/KCKaLYKjCBjYTSxmvi8gv+/xLG4+/TFjYLgWj7XZ1laaBpe
iqgAbUrdoP3S1zmEnmxSxLA9Yg/Y8iKmMm/6u7AJT+c+UZoH6xU4mu+/kMBWJ5FUwkHa+8GGZnSe
XgMoYYvEGKEMUuZOwMigeve+XRSjWEDngM8xvacliLwxdby87kP3/F+ICwd45dfuLWBN7e0Lh99w
RD3l+WkjKvzB498j4VpHC7pcfbHUCzvi1QAkqSJiwe90ORjIPS9nFeI0Qw3O7StR40eeF7OEkYqV
cnjhfMjmlC0XjXu/YXUJ1gzX9uxnnpaUjsDLnm20pOLi8XCeKGV505Lo/Zo4oC+y8HunQ8NtjEME
2VYzh+uD4s2/Uts3fUJeiJ+q59HLmEeQqwZEGG8KmpAQJuNpt4uVEN1xEbeBAYaCfhK2ir5bM2Ah
dg5ok75mwefZ/wpHSW6W8gIEcvTjPII80LqfaQgf5MQlThFguWjeiO6WiI6mCMMbeHPzE/j7kpmy
ZJmvR+gWBgfYWFKU7/lAP8VK8A8RhNikEq9Zxohd9RFtxLUXkVj05d+PZ39vCuRWYvh2bVK17KJb
XoTQfHDswlijWGl5zcgwDWyO33lGaOfm2X8rCM80vDNflDN361hDOLjnI95BKCyp7IFQSvFa6ncU
iVRILgL954JCAgeF0WHEYds3Vs1aUpqup7ocOMYurDxcZ/0cmFK1C/E0g1pUOOw09qRxCS+YrW5I
V3e4REUjKvzojU6jUlWj6KDhaiL9aV9fnv9yo6VWWlod7b72mrAe7eU/erN3vG1BB9eS5VS1JM61
IDlUX1zQkAYWDdo8vYXET9gvpU72lSXgSgUBN5cA22R+zqj6tBxWyTJ/BCqlmKKNb1D1vxlLlClI
tRxjkMeMlrFvk0qlMLakuffr4eybvtzblflJFNtCssBjw77rHnryO3djN4A020WITrj9Bb5CNmZx
FXZ4i9p0ORqn+189BSN/W6IFlg7q0ilgsTdFrRyM3HSBhYtp5y0tvyz+kQ1dxT93Ia21bQg+E1lX
56NqjdlSW1ybD4E6QyPhFWitVJw9vcqZ04RnMkdtqjNSkDkSgyXtVgSDTs8KXTHKCB+M+gaSaW3t
RxHWg0A6ZkbcX8lWoBO2CUrAbj+T6ojl9JAWxNGdpQdb4WBq3c+hsa8Ogd/DPX+Bk+Td6Mj/dXgT
nOm7osAe97eMNb3+NNcyN2OooOwDaBcee4toZJ9n4S+i0oJ9KevyzsmpIv13L+kj4VTt4GIBUrB1
rVvBxcRCmDH1cz77EbutlwcfDGt5SZ7oMLo5dj/C+XpBCPzcSr2xuqTWEIwJ2Wgczw1Kpu55YQ+E
8iNKUlqpM4KziEGWedhJ3Sm3hvhP2/aBZ4rclooMSNna/wnTfC+XVGaADZZtil6grIHN1I0RBQ+O
yCU7c0miigmLGKBQcrkP3shBHRsq52ng4NpCF2K4LvGSJ8yzqYeURYUWxehJhiT5u+Xk37hIeDMH
wazlvvDDSrBUfM5vFoqYMZPV1KirpjNjqPwfyc/xU0MLPKP5/jpoBltBFtB+ZqJH+4YaUWWY2KLs
ApWlrg6J1ku/R+8cT0Qgg8hUSA3qmwgRBKCIxrfvIjza1oe9UCXfBkFwkjXN+j8h744F6/zuf59n
30G23hEYrFIv+2cZzEkCT+JCVXzLJXyz9O4IjiIW7enlu81x7qsXHgJsv+w04yrcHFEosuFs0+6v
KFC4giiE1Ub3l2/LRcJdHYvl6N+MdKoHkmGkC4q7VISE7hACtNUNVI8wz/6satPFuUm/HbtQDx5k
flyDbubSRCnxItuigKmKK2kyrULlV4sL6BcrS05Yuh056ZZPuutgrBwrGdl9WkodjxAST5CLQDv2
4nDSjXeHZvFDbMxmqArNbfXzVimTzxcecMKd+KU8bXjWzT/oRCbOZRVJMeKFewWf8gTSNO8MxR0o
d1+TFP4eryRKxnm3hlJh8m8wmWXypyx1oF/L2mGjf+yj6+4TfZL8kTwCn4mC8scIUDtjSMFTD45Q
PDhJfIy2v5fcFc9h7s14njKoQpsV0940JhCDAi3UvmY6WIqRPhWWztLZ+A5bj0ZXNxqEH9MLHilg
Dp8m7IH0OHGuG4qEAJSq+HI2RfM5uRx07jxb2UukaKBaskLAGlvFcfinrrJ0sjkcmaRG87sYMHL0
jyOESlgrUKEjSywBkNUAWp18l2+wD2l0+TIASD/tNFKe/BUowYGKB/vOVyC5qGiUXj2jqwjUIDQl
RcvNZhBBbijWzmTo150xd9vDH9xtLy3wYSNdHl9fDC3QDA73NzzeQCWjijA0FJ8e+fjsVKlCIR1O
OxI4wlxRcQtuayl7202oW0olwpjpV8frupDuSMSGH7SrvCoHG5wgMgWTwF7lAPf6/exhk/UU8SQU
kH4hHx9GXTlDMhcsscg+yBT+64Xjq2M99jY/uR6Ff3zczhjVzIjf8VuSjyo+Klm5ZNmiA0UmQfgU
LBcRdX7Ii0/djosBimc5vh0o0Wfdu2bJe86Eh9clqwV/IkF5LyM0o2Xz1KgRQBGxfJjXsFWe/dgh
wMZYMDdvRL51TfdA7amyfxD2wHgKb8jKTtNfck5AOwEzO55RwRTuyTQJAbdU5yonJrmFPKJcVPtI
r4DOXUJRIDM6nkCwmFVI9cVSxZH2WAWiVxtFy+lAUMFFTy0bBX/5BsTcmBrZlmJGXB1Mx9PiVePI
JKDsH+dNxo+9ju/VuRUHli7Hik5rPSAKgEUesAXi/Ly+mpUZE6y78rtlxLyTc6e2F50tSf+7s2qM
SaVyBhG7hva/doHUR8Ji8sRv2zmIDZlLSaRm53F92Thj1zL6emYuRPG992o4dM/P1h7aRkOswYne
yrKi2MCohZs0kfPcuqFlyf7imG11vFE29Aionopy0ehutyiIIxMrUT+udi7IT6Uv0rjDpEZ2BpO/
tSdlfoqEAdrNQvq/31AVjkgPrZXl381lFAIa2Y1BXZOSbj47/xL2st/cpDpihmABfygjZ8D27zcf
/3lCVaKWsEKH43WJqn4x0QdkkpsECuxt1Z2QOI/mFkF6p6NTSWcwOLqbVxsSjzlsHf/Vq4xXvLVz
gV2VxRQgqFl+k1+vj8DFIyRWNdjmIOL+dYeLxJhvJoLEPMYYiUMJKyBH+6Y32m/qVqnCrDykWf3u
9X4Bp8Okb1JbTQDBiGiTTF7EKtpYdSPJUpEl4qz40TYM6s0MPsCpBuUdfT8mqyQ3Fh5jaQbUjE8f
BY3QTIlzcDFmFfjkvd1oSrGx8qoVJPmRDD1SmRvGcbCWeXRFF21XHAh/HlghZuoceec2lPeGPTGv
YNAQZ/RkfdMujfHPM5zWfbS7EaxR/DN0cz0fE/CeNnEUfXI0sPZdZQib4IS21MASJ1C+FgA0umrl
tF008D1zIoIubZZKbTVnrciH2KqvqmMzgs+Nl0AHWewrOZVEuCh/SPDOzJMSXvvB9nA6t1ynLgbF
isGMyZzZalJIhQw4BYqnAwxtDPaFYJLFoYWnjz7A2tubu8crT2exaztYc9Xmnuzpaxxsvb1qelc4
O/XQR/WNG58vcSJp4HRQR0O49VliTHiCpJ69WtzmKWarzcNfOwvum5iCROD9r6lgk69+ruIk13q6
ZQ27Lz9DDz0ipZnvK0yCuTUKc2iarSsSBUARSH7ewboch8ScnnCIAzRDvJjKMbOaJ0x5bkBDFxMJ
IxRvEUKAN9EvaFfNhpdYP/MyRCtG8P5mOg5c+ZnU0w3AaoTgjamJdU2gLm7EFoBE/+6jj36+sa9K
8F7rNSGA6PMxUo1OURKxZNUy50/xsBbJ6tDOqA1hC3ELZEUUSJYsAnjjw6DSPCSdhLeSpmsE2N0G
16e5QB3QrujdICS2EKoT/2IsJZ9xjG3Ts1dUF4+9ZGJZlZsEdqLK4M983j4sI77tLPb6tM6KzMXd
5kx0Wuri3mCCkj60e4/AAOkUeEtf2613OXzMZVOgLRBiJ7XejD0Bumjb2Rsl3b8frPNyn5noPwnQ
G/ft17G/sp47KHsMMnrFYIhcnXoIwjnEnyr6K7BwKbDp2yxaa42b+nVsXwvv7hfSLwOH+B62k25c
e5aENSOHQOc4mdD5cwtrS0fbTpafWL6JrdXgWHM7fLY5oVwrBLSrNlkWKLJbQkrYMq0wt0NlgQbq
BFy3xdxyKn3Fh84/nAiEt9Htz1X5PNJYVDqHDJ2L6WAgRHYgOQHfW6RW7hvipQzDuqSipBaH1jQT
JU/SnojWF5hCWytoXJsi9IGM06OuRrO8yUsmqwQZO+IkE1PmL4RgTLIGu+F0gPF/U+C0LI43KstG
6xNYbVIS/cvNqJE01vy3km5vgYIWQNXlgQHrwRGLj0mTYBLBMT+OnigcLh7mmcHhm6pFbij6MP6C
gsGkhysnMHfrin/RZB7zmbWl1XASATRixue2e8oi7mTRjOnpaSrPonHiIsqGKLl5WRgcmabyVcwd
YaubdQ7agNwXa+6pBlBc7sE8TIcEA8KBLdRnApbPXQlBWB7fnWGwk4530oWrtBrrdf1NEq+Q8cTt
rKsHTnfxKvHuwsuGkBgAC5Jc16hX+FHXcLzAVHhTQ+HPtlUJvLXeCyeMHFBuqt4t4HaUwLv0jnMa
73iyCu9i1K6h0TiZeoYuShBYl9qpYz70qxgoKi3Snmkc7Jz7ZskgnggvVu3LrjhSgZE6R1PkxlqQ
MFVKHKOk0smyhuguCapPtidWnZXLb4rHNExpjQXNOvdhBH05xEiO7vFWP9B1WGwam+3U7GU4zTFu
R0KwoN/OYOK8G+2J4EzUnO76wdfsjA/IapaIii2OdWAKPDCXSuM3fkNQ5c5zO2k0O9iWKErQoYxV
up9Jzb+nAGMinHfT3ux/DXaHvi7FZnV7f7gbRKoNzPt6CHXR7yamoOIGT0XlKIjC+xI9p+8+0BQd
hCZ/BDFnqhiPwSxmT7yywMRe1WP5ZfMSpwqxUWksjXGxUZ8f1sGd+ebKqNFXTlfgCbPv2Acvfqxc
WRzx36PgzH/KEoqcxcKWkZ3owBLz8C/kyjsKtiNw8gZKxltGj9wJWcuUX9n9DvwCSnTyGQ99Kh99
6BeV5150Fk380jvKCsumH3NnjlhhipDGX3fDgtK2tUNmuWpYosUyoHv5T+qcrkrc9o8ZyunAMFaW
oqLBEW6HnRvwcAbvG0LsXmZpb3bkzKzHXV/BjDatzz7Zq7EsLLPuvwYPxU5dHGLu17gogBtCGqnk
zxpx5egNbBj+hDwgAeZP4afm29PydQXoU9ak1vZjEHVMAYuc0ckTkjkUT3Fe2ci/WLAV+lKI0jhf
byXeVnwSjTb6qKheDole8BYQ9szi+EWZvDPTy6kYd0QndLPYWXwCQYugKibKD4x1cZxLFbwkhDoz
VQ+/HPVZM7lEFoJXZ+0UQbIppuT6KzkY6tHtVL1bg2SbbCvTp31KKKJb+WN7p/HH5KGsoqgpRlr1
73yT8HzpKkMQbLgnyT/4+SCZYpi8tRydeGC8ycTtjgqBgq2Ra2FDSnlJTgqrHwBxipoLDmGXhfaQ
oxuLLWZyFso2FRzIackD9zUSjaOySFYjaNgvL3/OCR7ka1QdTcHF1nb+G/Zu6r1d32yFS3Hx48ts
CHd7tcwiemhjWAzfRZ9xq/ToFllJRlhqtzkeSOXw90qL+Wk8WV3rmEEeO+dMlZ5ciFNSpYoGyDKA
Gjv7iXe9ztX25nn+H66CEBdGZJ2kUOC6viWHrqsJQhrE6uVtgan1xDuqXBgznPNSn+vBCQZbhwR/
t9iKaxXAWoycZ7RNK5vOLUn09iZy+ORPTwEQHfyesNwp28CG7L2YSTwBtQzQKNT1efa1exLhQwdM
fO0YUztDnQHvoYGjh9fCMTN5MU53K+4AbeNSJ9z7RtQa68C9VJmUa8NC0Z9Imi5br2Ke6Uwgm/DE
4W1IYRTJ3rauI0sHEfv7K1iN2Yt0tgu5fwIc0SMlcznNw1nAsFg5+mC4caOMf8xMbta3MpZ8I+oD
VZDgKKBjDzN8Y31egz4QAYQZ5Fd8gzcbjp1xsCW/8HpCWQPL+Pc2Bc1Q7L3iuH7YvuaK9yaAGqru
Ub3Uo9KnOsVxpjqUvG9K4z02v9PORbHKEnw7fbEuL84OUzD81dzKu8RuHR0rjBgcm6i4I+kKsW2o
ggHn1c6H8itP6s/WG1XRx+rFn/xws4kV4f0Sn5lxiI75e/VLVBllB/hk152cT72jxoWgzSzstJzu
NdI25UpG7eh4Wt8TGF9rGa+MDVz8xk0FBbma5i0JIVQbcXC0vLCdxPPxINrT5gRKBndsFIqFq6sG
ElUJ+jU4+C9EJ3rcqvYrbUML33D5l5NbPEXZjRBwuDqIR2k4DX0g6PPZF6tE1l7IfvyFVQusaBfl
IqBNOzLabTMaMgxK7dbdiDxz5Fb/7yMqgVwOJhAxeDtZ/htDJ8SK6r3n6zByxubAdp3ICgQayK6Q
AoXI/3XYj/B2y0ulO5SzZJVK8ikWw2ZiY0agnCNFr24J0AqQbaXldEPcN1YQoL1hOY/syOZR0wrx
HPhU12oMO6lTG+DmnOoNTuFvAzGpppoOt23/6UmRPkoOqCjpdO7Fj1yPvX1IezPg6vOYIqjDFQav
PgrV5tFzlpvRKxzgI2dWtbVoIUn9XhfodPjljQS7yWwXGmSGVa5/VJkjr4VoJjXQlaByO+5mUAOG
YNm8Q6Q2tu0361ftbbG9Y1r1nOAqNc6SNUwyCI6sapY5IFf3YMH8yqu0bEgbOtFhc2Tql+2bDy2D
WH2jlD3WkhPnuVxzCS0biZfFyWXGUzz0OSpAwUseRnJU2AWfXuMG6vL0Wy9YVrchCBcsVHJroZsr
mqUt834XVWv8XcljHg+UBtN0u2TqeQzTlNEjScLxuhwljiZJICOslYf/qRlKf8wIasa/RP42ZSpn
J4B2LLlpQMyc6ldw0bFjwZoSGTpqYgiQLOkqhzA0y3cih26LhAmJNoRzLmcjbNNewqvycQaueVih
aV9Y4NiFq6HlpfVYhg1Mo3azUhas+cDVBQgR14RcuDl1P2rHoIadGjHo9tGp+eLxAlFjZ+1gxVKE
nnGFjhCCCqMMaEH/ZS28coPHPe5aVRrLY8E1QBUjkTX42eLeFnoLYUmeeSOuRNQ7FrqvwaBHelCM
lWOveafa9mmUogMZDJiZo9u0kQh7UAhZ1jW2i1WKxDIW58ce9wZq61AwGYqz/nhfhqa3B4YW8agt
MvJHqmQ1raL7bjeUhBNgZI5fESpJqPN23Ev68CJDWa6Ky9b5bLHshCaXJzfQNGPO0pwCI4yJckiN
16FPu/VXv3c8PJzkZ+x3OYtQ1owwF7EPYsOEXmCAdDZ3TBa1NaOmq/lJ3R33y/8iRlKhk0ii7oVO
F4Q2cmlF9GKER9S8TlUunnaf2bCIt+AYTbLaDSgSjA2xRpsajJU1oJK2uzKQghZVUeTitSLu/bse
/OZ+MHA/WVAs4esW/eTpIckFYHO7UemAkOmO6uWlwOwXgdp7uR/2u+Y3JtaXCF9pvieJ1zAE/ssa
sYjsHiB2Iq4zXxiEUVD9mhO553GwmvvWYv2Sske1O3pQ191mWQLbWJPR65vO0wwP4N0QwQglkv44
7D001Vy/DEH5hzwntxHehejwPzJA2KxdlSMNPrNfsNyl8rW1eW0PCWKlggf8ZQcYFgXQYB52AJbU
63JZfOW8FvhIJ810kApKKHbs7hETDFN9B70RPc+X5ySN39wigBrzi7NgQIrhWVdGLEMZY2DxmC84
VACJyQ/624g08k1RYj+/w6nOoCNV38fymE2oODzWUdasUA4/SQjX0ddd1sVuOER89Af+41EXJqvm
zDmAeHP2YSY8EzezxOAAmC+qH5iCP2WPEdst5LyLH0HUDO04ZMkm/KJMOjhBJHqMd8rdbxBYzSy7
7Bde8zVnp6e/jrw+BtyjJlx9gQgS7sRqcSWOJBlGQykAz2aYJ4OF2GXzdzOMF5UgIfdS56Xu9HEU
QVoqVB/1nOkTlZPE7BZ/oka2H5ceLwIVujK67thxMtivjszg8H8JVkNzXEw1tKjsgWKlK6e5zW8E
k9Wba3wwiTBGfevRgYOX+16X/RSw9QdS6G6ipvS15ufO7wxF6WKVN6Q3SpUb+0OiOvkgFKOOqeXa
7yr9fL6ZCioNdUcjY/sIR/GQD/U6zeR5O051Cj0JybYZ0en+KCPbFn9inHtVqYjwqhn3Rf0e2uD2
6vq09Rq8GLqXRpfJA4KpMm8xSsofNrDIsJkhUn2+4f6JXnY+8wL6pEog5Z5Cv6tDJZmhYaP/ZjNC
H9KgFMc52FcKbrf9exj/ZtnEKq9+DhEDmqVrTMOeLRLv6AkR0zlKqo63ofVi5HQ7qtcJmzc1YTeg
ZzEEV49bcjxnp4sy9acDa65A6YLoJzAroBinVIfF4gycJgxIP1cy5u/U7UKF5YuLX0aDaF0ZEv2t
Xw5SfMz0OpHdY2fowjRd8Yj3NIDIBqVjDtuiGl6H6meDy5groXPcv9q1dsWqWILXe5092V7/8Y6G
yPP+kGj68aWVN2rOeOlABQSSf/i2xNTv26nBzmF/+SzaL70slFqkmAPNmquLTvgWarZvwOtC3oET
t9fwwpBRL0/NjFgZw5je4OpAmXdrVeoQ3slPMT3OsDjnlPRnbtsngyCKz2EJbMPPnlTfV3IjhVAW
nxLhWEx1rNOed58DvGlABnFHTa/Ph6tJjX1sMpmNvKPkbF4+Aq/YteDvSPi+DgugWrJVrgwIbrlk
hNQgAEw8QbiW2nKVnO2sM1/I6M/QCBPnSi6Iwe2vhpXjBAHkNkZp1lORnOhAxagODywraDYtfqLC
5XbnOTiBgfLnEi4m3qptDploFD93YJxAVmE3bgTFFFoMK5wXS/UFCB3MoCrPGRsoUaiRkLvXPRPZ
CIyTYnGwrDN8DjuXcaMQ+savd+E4W02K2ll35bk9es1ytwpIo3lFMeypYkBVjs2xmUntCokTEHeI
OgKR5KJk1G0WSe8zVQ9eK1NzMkqHqxvLGuHpfuTjx0Ou2u6o7JFIWGNEejpJVC51TvdFzbUWvpzp
GV4mR/fbK+94GmhJepPOYOJ6DFH5KOze7qZWeKubFD4vgM2Ac7MMAUt+ooYofdwml4bwNQjD3goz
hzehwg1q8scXSpiklD+Y9QzTU4fAfM/88IWO/bWG8xQSK21nCogEiSlTOYjmSdFnyPYXGJvfHOqz
wWvq0cmlfsuEipCYIMCd8OngFcVRZOzSVG22h13FOAtsOqTcC64Vneb6cTDMHssWv0kLDjY6g+ko
9f4cW8Ris1KXBQ1FpfjkS7gaXXZtOnNAmAFnaHiCKeUW7ffBYjXWstMrNYFzOBLYGT2YpDmASh/A
k3zWzG8f3fx5soLklkrM6EQ42PWDgnFZ8GBA5ntbEGRPwCcObXYpxa5Mh6G4dexBXYYvwDMx1rXC
ktZzu3Q0n8VaGS4Z0hohDQQAxyYNn52fkrRCLsj1Cx8ojkGzoGL9DUBuuaDppcygu51g3kUbUh/v
+oBeW1WS5TlFEXp0JXVx+M7pvcAJQbvvjUYrvhSYyzBYNrAANgugryPi6kT+MDLJlvKjt/G5N5vA
g5J1oplOC6PlOfySxP14vhojG5O8HHm7NkfraYzVlHlRz3X3gks/2th3xl1ixNVNINaSRghZuwz3
+r+DOp7oBVJ6QaRcUeMrB24qxpc1f/m8EaMGbYGfsCBaZ3VyRd2VrFOYnlF07OmGAYH3Ed/S/qOk
FSpJ46ZMsO83icfoCMo8WcNLI0XuZFjBvWqWssEDxO7TSYbmFHWzqq8SjLJ//AVZ1XlZQapWRCkb
uDwIa6cZHZz2jcQJWp8iyWTGsuW33wh1ZGJBJQhJ9Tnd0fG+cAsIHSvJwZjXPvZLktrki3SLWLqi
9Wip7A9Z1ccN8pGYKMPsa2dXGVqxPM+hJ9ka3TvBz/Q2Wr/USAXe2p6MQx8V75PZsOAq1mCxJtcz
cBnCxsQeu7X3aW7MHQ0pMciJ/H78xRn4GV1Fmqwik/cnQYMOaNMC2AeHK/1vaVxYQd9i+HtogW0Y
NxeMA4S4zGJBatqW87XGsv4AKHiv2MNIj2CDMgCgTaw0o1ojhpVHOx7uvxOirF3LRRfc2ASwn3sZ
WvEZYwTjpQfxyEpy7siFkbX3pKRGW6+bRrbPv89W+IZ7iOKEOhlLCR3z2qM3jI9OxowSOPAdTpof
zGDNlNJH6X2vFrk656899zzvTxpr+PTO47ijD8KnPdYEfUBqz3yZK4THRGRZ/5LuXt2bJd/wC0K0
ePHXoZ1cJnTSSBn6JmYzvXOTNSUD245qdR45TPVkfx5SnOM6iwzUSwErLRlRfIVXGFaaoU33RbDD
SiDS8NP6nkUp5G7nziQ+CecHFj2Jb3DGyxudsvKl9J7M0X2FnpIT4VXgZkOeqrOZT/tM/CRi/egm
HRN90Wm53FruZ4Mj2h3etO9WcBIX2s8YCfaYVGsr30BqwVLkemN2n1yDuDwxi+kZD0Yrhw/UUdmB
h1hAiOpWfyLjQC57omGHsmrgTFl3gsLXq+m7njinYDP+A8UM9O3rUbCpUCmI9J4/0VQ67Xo3wy9X
r0vYaOzoIcMj1pZhEaCvCa3RY7JqYNvUAXHqJPHrLRazKbNlioHphW6w5sR3sj4fW3VFW9HslnTg
0QUoxcTTxqOphNNkgvGFGBDY/SJWd7xu1bvjcsJCg8Q771LjdDLghuaSAETbsuS04C3/c6OXlRIO
nhhvQQAoFevU2ZsmpPHngr7+A9sNwwaoE2cXOl5429WAMG12Ux7VXT23Ac/KlnqrjHZzR5G+N8/Z
q/7ASnMPxmiQ5qUEi2tk17y5KEzcy/w12FBzPXhTLIlTFmGu4Ha0/w2/sx/CvPcuI1iGhm+7Y1Hu
JXE/SSbXmRZaB9EcpZAY2vIFjFTA8hph6FfHoI/l+6Ht4TAL8mMlEBjeqkfj8j/nbM0AZ1BNXNEH
+XdD2M0W/MA3N/cVUab21n7TnOzPmyQV/ezwvzt586UIjbJEIlF5nZ0wcJ3BeCldOuu1gmcbYqyX
oXZBA0k0lt6OwtmIXyAUgHtCtiGknCYl2WsTQEHnRddwGazni3YIe1Awe6BNIRhUAOx76uD2soUh
Ud+aTVqzst2mr9rFt1cq1zTl/wwnMu1B5mW33guyWjt4riSa0rYzMN005LnO63NfU01p7eKHx/1w
hrqhS2p76UArl1EY4Ak0v7Ek59vbziZwkXyg/5iHDHWZC2Q87xVBwtmrB0Q5yl6jNTN5NHk03FT2
5CZz/VMi3dEv4/h+O5vjN0Ys0iVImX4H4wysddrh0j6JSxWh41aTMFg3k970n/SPNazYZwmHPu22
T4uA73EPG8gsSXXk6EOxl/ba0UKi/O63e06sBAVr4HGsEXMPMd0/6OGoQoenSUZENMEzoHQ7O+zj
co/gwVol8QBcchPJ8qZA1PFYzkNaRTaaocCIbCbIBhcNh7sVIZoulXvP+a3tF1kIqXGSoqRROepC
LZ6vaxWGl8FY5An4QPdHGfM1nl9M3Ee8vHeLHzRTnasAGOlOp2Rr1b1Z3SwSenx2wTCL8F8LRiRA
r4dlulx4d8cOrulVpT7aVgfnaI9uqTVuE7gH5ec7zv8pEofUCE9V2tihK6Jeje++7drBRrXTQtxe
9VRP8PR6SUXmnr4c2j6hMSgZPPSa3XpAqoF/lAVditOwoUJ9In6h06hi/wvw7Jb2q1fe7liIDAT6
xy7yN0wI44KDz4zVaTvHb8KAQJZq6n12Bfo4YvbBXcuhcmOgqozubExRrbM4+8xHqHlEQafcLVQ3
Wkmex0T2cxXC0bz9eVU3zzaJdHeutr2pXn9yYM0/GwgjGkvmXKiFmuoZZHBhiPQdzh+kcfT0IjBq
344U5QEHnxfROr5dmONP4Xi64g8C5mLUG7702QSykzul6O38foMCK6H5xmaFhEyI9U/yq9S4P4n6
JievM2fj0lqV39siMW/C82E6EcaK3qH/wQ/RE44IsO2BvzsQoEr3tnqE/RK9KlfCZeFEFBu/suEi
yHKUSfh7kldJoSmLvD+bzLRp9jUCcxMtmnxQP1y8At+Si/6Ote932eOpSxoUxJYa+yIAlGQQnf3z
ILa6BOgDz5DaJg1cNF2Lx6tbazoWW9xnPkXkIoxCBLmsGTK+05ECsLq7zpt0wPMJaf8Q0eIFcqyS
ztY5DbmBGrOnx3Oq8Wc7iPJaiUiTvWTm2zXFESLcpkX6P+MfkLmTmE828fxJ+mYMw9dnOOZkxD++
etfW2G5gjKTiMvlf5hyyTyU0DU1p7kgPKpZTbf4W7CQOnusPCgnQEL+aqAt910M4GCBAH9wmtEks
qlTX4XzeuB9VJKVPfZFd5t71R8O00dOWSZ/uQhqbAHX4/SsmoGJgGu7krtlrBrqaO0/moMsn1Kof
i3azsqt/AMaHROXdoAp03WL7IjtcsKb3MG8rBSl1KcfUtbCBCyMwrNnQASTSvWYE3mLDELDQftxO
PAvCshYVBOUwE+AJfg7YQVsEqj+GYgd0r5uy86RVb5QxYzvPUxWr3nxsRrNDwidp4xGMe8Xc93DN
sk2tTF6thke3//hJDn15OAWwViNcFTcQJ2RjetsIx4MCnt+j7yWRHiTrwsWOVH5pbe/ZLCoMWZn2
NeAxUYHw1S1GSIDiwmH1ZsfrXsy4xxaVyHEBdJWGqrzs6BTZ1g8ftZhpOSjoJgMazYFlrfSRiiEq
eM5wBpFDdDH3g/aAvhbnTNYAG+5IfUrgES29tVgXdL+XWyNTG2OkrhUJHwqXA58ooRbLdWZOIASv
k14+Xql7wDzqOYLf5LvCwsI9l6kwwRRVy6gvfeuvRn7s7vB6mOOJPph8z9nsi8SYtv1BLrRjSmbe
k1xXQVsIhZ9O3GuI3qTRV8GVDpB3KpjpFDzD/Bhv5QnTPXQhdh7Yt1QM59QvIluLLibf7HJwlLIX
0YIx0xn8jpkuzAgxrzdu5KGbqKIe3Ufe7745v7MmOE9iBQ06ALMHdrJXwaJDEn8HYkupVSFgMPlE
5AL0Yzr7HxV6KemIjz445qbnhP/9ON0hhkxzeRadHC84dQtEBN7zMy7z4GTBM+I1xZPVPz2/NFDa
qrvPw/6+CXq0CcNVTNLhCZnAWscThoqUw8T3kl8ahMEFD9Ut5vf7LjyeReOVexsF1HHBzyP3/q+W
6Rajejn+iR2Zdn0vQZL5yFF5bH0AyX3tmqdUiWDkqntiFpXGWocPlYltEoujl2OCEjqZsrhPNSWP
4XObfz4zsmS+LwvQ2FTJTcNOunvPGCo1L+iCpq92DBUkQhSPR68LYsFz+BBY/eYdyizBaaK9bP/+
efrVo2o9xBo+7NVkliDbBlk+d7eORvcl9SuaZyRBdMnheQfLSY9D1zMRqAgZQS9xq8lSXyN1afbV
TgnGFlf1Hsd4Pjn99RO0GuZZC9ShBDXpJZ1KSsoLNf40+hL+G8yhtdFO98B5QlVTJiP7gEC0XEvg
4W+drT82OFncKi06rTLTeVwJfu+TMqUtp7uB14FYktjnSNX2LaGVBu8ftaKUqq0qmHPe5/eYaTET
t/93Ik2Pw/lsCOZs1Y0VKteYmOFkRwXtZjYuTMGLG0JcnMyrJ6FbZEXVolwgKvgGEcegSj4cyw/4
Zcu9VuBu47znNinG8N/F+tvmb0BNlFa65Ebj0n+BCvVX5Bms7dz00D+mJX17gEnuXPOvxorxjfXs
FjK4HSUer2SztTmZWQqVkV64Qo2dEzNBTsQ2uNmtWthda566VT942qy4L57idigUnGWf1ZHkaAsE
Jynxyve0UghjkwPYBTMj90o0jzrRU1cVt/2oJLjMBtcasl8BmojLxycq/LGo2FHATEXP2UpM168y
GIAbzsElFWRfzMPbbcvoth6J2HciwQKy/PdjuBHreYn9mFEecWlkULC8GH6WCrwnu+2b+IfpjMla
Q8W9zrlZRJ8GHHqaJ4shfLrcaittZ7bX1fOyTz+EtLujl76IzBL2to0zHfyztGOz8tfOHU4U4+Nf
LeDKoe7MZ/kRfTgYx9A75FApje0XaP6dL0bylgln83/+g0QLFdx+/BbolNdHdNoO90Ykro0hqKFW
ZRbzmhGK2IhEqsyacs+cjcUpI4D9bOModbIRt8CWMJl+z9AUbgxTvpH3j1bkw0S0o40c9UK5CP+p
1o3Z+NCQm3lNdj+yAzIF1XQ1qpVcQcrFieLsuAm35CaE8qzaYBzm9nX1c5ECEu0JRs01JdbAawgP
6FbkweB2FReFlnUjg9KlmEAEQp+Au44UYqzaku8TlKND0t3CVf+JCSAM6Wp4RRyFdcHUTZlxmm1P
EQfJFuOvBAb7xbLvg7uXTDwUycyhTMG/pgsGgKxz8yvel7FgUqBcmiUeuWOHc9QClxAsw8l1By/L
/3VEG/6rQhccIyZll6RQfA5B/BhGM+AkOjw1yzytyEuz5pHk19NRGdBHfrxbndDHdpS8l//drk0/
t0rla2clRghOsMIkql4UZEKCQNhd/Pt0wFH3q7kEpbWKpjpXqz0YDvz6IWAmckHAG0JSY5Aiyq5w
yBGbImfinXa8TNxlResPctziI20EOvYF8yGMTEioggt6urk0HiSn8RCuA05yGhV/oPWJbfborqeJ
rVW0KnMe4n2P95534zUS2ajIyUPX91EUTjAafLTOVQ+I6wCvI2U+EtJ4bJL1PGDAOY9HT/tTwkKj
qhYBg40hmuXOQVAWEdYIPSMI4WbO3rwbwveW7O+EcPCCAg+bb0gfPUAnFg8tolLYypYDh23hzAFa
3GzquryYOL/8DXggn1VR+JkrryRuBQnNvo0wbGeJp7yCUwjp2Z5xnYTy1p3E6WSll7a1/RQUM/rT
+gMkHPtC3ZpvHiFT8+6885icQLTchNB5GT/5BHWfXXThopKK3fHRhOIGbUOmAl/VlJX6ZjP9npZw
mBozuks14qH1eFQLITokIWXIuzqNsfsqzwyTlwPVzy1MIW0ZuRrLnKc7RygKUdvvGe/AesXROhkh
n1cQt7g1TjMZjO6CCSZV5HP/3NSf3fBaGGSMXL4KlQTVKa802TdbMvcc+SaKbD5Q5gBdP2oe0yrk
FB8ZMhZUo1MnYwFELPaj9GUhv4a0a/wAmfUqvdt6h2vgByWnJ5uwmPm6O4kw70L9RZYoTEjP0VxC
U2AKW8oQYEs/T5F0zGooMGsP5fUZtUD5YNDSMlbQDhDyJx/VGyB0bOvu8a4QzKBIH1VmJuxz86fx
1oGoIDcSqGSLqQBoLgW17rsWtsWfo0vPTvbBP1qH7Rii0Su0qQS0eGU53/xyAh3XpZfIOp87IbCQ
nvMjQzpSX8WL4MI9KcSBXtyqBKQX+pZjmRqUH+1vMHNUkLDr4BLy1SZyzbLxLEqh34SGNrOEtBS3
Igp6hnbsmRGr5rm/Nhsz91flyKCktH1MkysO1yA+vnRuU8if5cRZtNn54E+ZhrYPRiacTbCnF4Yd
5tuO0Rde204ButvESZrIdFSx6DKEg3sVALqXNwFe9k2BxxpQphsehCqE5GaIUfAUECNXk9TFGN/Q
1OuLIS2rZyLKtSRehK+nNALp2MVTd72IKIRqDCe2qNiYX6OZUp9N/G7Qhh0FBNUdFUPitYw1RDep
CIsJTIYVvlZ7XGw4/nz/g4pxxIvTQdfrljFDC6RctX+h7Zdz6CWGPwyAAWbaSjnhroqf9Dw3Eisl
HIczUH325bk5w167ZXGSarUx/aAXcFf3NgyWCo5e6BSbHa4/oZNxM4Wvmkyl3CK5L/o08jDvmiWq
B6sYaMRioFC1LDeGkOrBnSlSyEh14RgsEx3D2sXEg6D4SdlJ+CnokXONnRD0ppYtoDx9BWA+C+Kv
s94fh6qzllHWnVKnHLMIeKCtH+JrgPKTAPEC+Mv7cZkCBqRaWyI69doT0P4nVf5v5zGp6dbtUOAK
/LNqag+qtmzp9myDxL0ahQs+fYpPTsr54keiWrS6n3S39X4rH4eo96p8SgO9kRkS/KIiZFQQKpVF
b/Cu8c1S0FWT8O3Vq6F4cqfPtTtAld6GYVLGHLPjfyLAuJX9rt9QQo3ZvzozN4TrNQb+o5LxbNNp
U3oQFa1TQH5I6F7ctc/ilbk3s4uhbGqOFbC6tjZUzB3jdPBh5H+mR7yuIBU8wa9M7FOO/NuLYCsh
M0mhUVSw+tejYysePX8vk1u7isHfL429cIwiA4nveSgghLFjtGrMU+z2unIEpj1Ihvh8Cr6Sox9v
RLkpeuHW4xLj8QFLln4UOS4ScKRqz8i24Y30mxy0NrMAc4kul9sbnorqKU+MZq+oHppAwIO9WbpH
X/h0o+Wq/94zXvdRJIFWM7/URq6Pri6h3/TBsbGwsubLLP9SEVz6SHhPXVaot7/blCpOLDfqM0Ey
p+buisZYb6QxJUFuAvI4XgUmLUl5Ijs987YscHLotasLE9IDjnlinEI97ROwOv01VCMYefuXSkmB
Up4cF3Vze4/ZTlFBwog8QjraAPWTCn64kdm11w68D8e4IY46BLI8bz96STEZDMg/6Ngf6muwIrT7
tyJKn/ybuhwt07zM6TZM0NZ7mtTiYP24a3dgaD+JjbJFuvFFqN7WL76Vvayainc2IIMzsmZGmxvW
CJccqbEG8sWUopyrYCJVrj45f2OS+BCmQbAXPYjC+YFwDG3SQ9fRElQp9riie+lI0CreSbEZ2Stu
fYQ7plSX3lm8P9FL/gpSFisnnqDKB3TjFrccujDOHcgw58PJ6AXUf+ZrnpgfNHveeaKeacmLxB/8
DRurDeQYv7KAJUJtrVB3OTf/di7O0LWPnwD/TW56BagHUi1EEUQLpOZAzg4zFozrsLEfyT13Gudt
RrOGxdJ2bFif5HeyyN7MC59Gnl/8Hzi46ARFM6S+jhnueyCBjZjm02+upYCCSNrWlyj7wmYwQIRK
LLtC+HSbJbOpxqJd8ezA0Q/C1JBW5466+J1WDe3MeGbNZMAkWKD4uwi40r4vSkfPN2MnciOg9ArE
D1c8kQRg0kzJQrkmbrw92cTbQ0WkV3peo2f11zu8cbukiCmARDwSH5U6atGH8pQWD5jlUrnU5Jne
Q8hJpim+x5aZlf/gO0Wnnnzgg2TGIAKRpnyp7uJizIfzerdl8dLjTOji07cZknwHbU1KlZMuHgHi
VSFHZlWL9g45eWo00hQd2+g5sdWmt1C4B30p2T54kAkWKv25Byvdr1lMlBJ9dBUvN5OPRFC+wYCD
1diCD3hqMMLpb9gb3DXBBcTikolWnwJPt6qm8Od2reIRDpgZFJVoo92PLc8CsiBU/5VQ7jinVmS7
ggnL/AabTTnHUzmmkUOIMY5EmUjDrxU7Q50O0d2rStbeMSZmiOOQF+HMvSd3/Bb37LMKuk8w0Xat
AlTaEy3Sj0zaGEw5rTr4Gg/CWVIRO99HH+28HGiPMfae2/TMsQxaweQIhTfi3+DdWTHmybV072V5
RTFhisOedYUkbSUyVaz+4BIVZ1bHe+WSGo8s5Pso4KfSmUvCpLtOcVKiq41/+c/ZXUYD/8449/qw
sgjV1ncLXgnnyLDpc/GEykBbCpfKXZlSTGqx9Y0Wme0/mXg9nZOIcbcrSEt5bgnB5cytdhTbF/Fd
0PZH3dLYjxcJEOMVoWjbQZ5DdDIBlOWZ/PmE95AjEpfm6J6Yq57PdI0T8lf2AjStk3EOe4quAYtX
SeaI5AAf1QdR4Vnt6Ny3mzwVhvg7Nrb0nEtxhOFerIXQ/ZJy1mMxncDmgsYKhE4R2D/+MpSwEhyE
fjntsfE8hA0LnTplm/UG13zd4XpRAQkS4JoH054xYM14q6Y9XmBsWKm+AduQCg65Y26nqTARcxbA
5c1c3FlJRdulwcV98fJgz4MhkHMynyxmKbzuTrFt7FwuExgHf5yQIOYGmrXrO2QJbfTAwRX6DuY/
C0kmNDzX9/ARSUDmuLs0D+wCtOSBnAqwpRZhTJ9T4mgjjXXgRztytWDB/35IQ0ZUo29TZaNwGcNT
Qz33xpwaWI1JmhJmoIFCO4Nn+EwtP6UqgzHhdPYaDOPrlw5EcIKlzHE//LpbS5z77H6m0wOjiOgT
GyWIDkPzOfLOneNhHBNBmxCDjEtrDeFMMdEQeRVefTNLmZ2OhFtI/gvry0zQbw5tv4OYSKNMAGSF
kLfsZCRKCrM382eB2vPDPFt4iT1P2g2NmNO0dSB5wW4PU8Tucn5hymK0HsovDoyOdF1rOACho7XE
4yV/vdHtv6FD9CbzI53vAYOca+kmOdUCwj1YFJa1kjoOuorMGi2QkAkh0t3B94dRqK0LsoOCm4mv
m+zUBK4jY0W6lPovrLC3LoKv39k3wGpsr6tunId9vUUtkq9vzKH65ELrJDxRD134lRzEx77q0Dqz
QPvPopAsbyiDcmQHRsUqto+B6SwT9eMQNxI8p8tS1OUPrbD2bmi/3T6JaroP9bB9hTyjSfN7ck81
Ka7nsDxReWtHzosVoydLJ54iNVdLR4Lree8TlgIIMSz8/aYm7QLJgXznBItdDbGOqRJXsAu9kPBe
BK/gmspYo5W5/Awr9Mr++f97piGaG4Q5i43Ap+wZAVfNa0TlUOMqHHwz8IA4GjLHz/ev0unZuRyb
qJxwaXj/AeGnAZplGgzlrmrtAGQe6SlzxJjBkjrXt1lvVC9BnW5p/7GGUtdM263X1WteV9QbLPxp
zHueL59GdJlc3E9OTOl9fmvGfnRzq0u9yT8x0wTLwhi3vRbvBujIm26uknCy17Rt+0AP/pqYFRJW
xZlFlUI+AuPIc4mJv1nQo3cdrw7yuvYVtXrGhoUVGOgbaoL5SQrlJhL0EV9WIpEABLmj77W8/JRx
4SekE3xpTDMZPtO1Jvd8MC2URGBfMQFkWTZEZk4D6mWNRktpiM/B+1YPYBuw8oVPKG1q6J13+K6K
eFW1FyQ5AxOHEpJ3yoDkcSB1hu1d0KXLG/sKcKZ1LaG6OmzOnWGY1EKZtxk9ofBcAH+H30+dWmDs
X83JgRdQK/R/XuJp9LPbPIteUZ22xlDKAJmAZO6eBVKV1YGZf4stqGbnrh8qdaYZ+mzG/M2iHB4p
J6Kdv3kowq/BwHBCl5XXPz5XS6ffJVEe2AdICR3kPECIfXFRirckFSj8P/QiJClOrGYrVS9BSTbH
N4QZgYHWYNMvgyn71s6HSnSPblXTqSapycN6S4ePaKWCiPyPAiOIXZx+oYvMZ3/R7Guk1SSfA/v+
14H0b3quHWTw+I1aon4SR/P3bC/+yGG/Qgmrhl+qPoPyRHC+j8TEWB8CC5b2qJh4gMVaxzpbDPRi
ILKLhf9xFPUgHSCVc+dWR0wtP97HfAAFqSqZTaWgxDauYVAAxiPw4xLGlbg7venukWkudXBqxOax
hJAHb1+WQXeIIS8GmqAfVEZop+mF1aK8kAMUrm4ZqS/4a9XItsm9eSCD0X/57zLSLw18P1yf7ZxF
wgHgyRSdf0id32OcPu6N8ziUJQnt18jYCJbN39CT44Mjo+cCVrJq/zm+8+5Uq1vI9OH7MrqlxwJW
cgrvWiYyAiJLsib5EV1mxUtPH3LbvxoY+tXpYjDblwKlRsi3FBoJ1nqs3gZAJjmNFZIlSBmvgTYN
yIJDhpXMKVNlyBS3xkM4Tufsi1qbrotR4YMofMZpZeJA7JWHx+5wVMMBePlyl9oezgrb2fVPxqRZ
prBeqA6X4FjHMxmXaxof+ZY+2ctQhbygac7eAZ2RJaP4vWXXr3koh7xZZigEfAGcclhwfGC6gZ5j
gntMhol9RawkpX58k3jS7kkUI0OipT4VLpbcNpgBtMSr6r8Ri2DNTK87O4hIMVOsN9lGTDgCoOw4
/Jtd/M1Y2/ZfmZ6pPjav++mpPD/cAXnycn4CbhAiitHRtARxeFftIWiHdukZbH15MDzAgf7uTSy3
iRUpELPkufrPqslVNSE4djBAp8qU355LY+WGSXLtbl+6RuO4IN9WTOQvzq68EqyhVjE11NLmJRzF
9Py1UeV4n++vbcuEMk2QLUXX/YGh5ca20fE3IZeB8hA3gI1/VJjG+COHjDjoJwpeqhy/UvOvrq1u
8wsPkfuZJM6MzAqTuC8eVmLmg07sLxJ2RisjFgp0jKZBZ4G+f4JXnkjX5BRSG40RReC6DB5fPNMT
9g0S4Xp77slH/bGWHdxMezKYPa64FVXgJry0s26yDyBL8bmnwTKBEqY9A9V0PW4MeDYED2XVuaPl
ZNnE1kOWcoNTIaiUbr7eJsZd25RRKLhD4F/fv4YhS+ynnJ/xCzY/6JdEw+WNV8MvLqQmw3Fbn9lM
63RVy7O1uDcipO10hrH57qgrL4Uij6HryqEZLbuWLDGL7EWOkxTdGIcgS0wtJUOxrHTjjN4NhkMg
Em52+hAVMowBqf13SiE8ckx1OdpPyh6iksSTDfUBwFegQUmDOboYteoeJ7HSj5jQ2edWwTY7tQYT
jGq68r6Q2djrhaPEy0hB+50yBLeMpZyVXQXbmFE61H5E2nqQT6eaV5qaw6VstoWeDrCvSZaVMiAR
1o0WhzPyxJBMJdU/3UbN+f0wh4D52i5ZofkhVsZKcSOGn2hQaDt3Qus7SfVjFIlgRmtj9HEVW4I1
QRV4+lcvG+x3KTBYrNdRRFCJd+WKI0gtkeN9uH1lZwPKqJZUF80rxMwf0wHLFIqJWRU+J+7FF6Nb
RRfG07RBSmNTalDrHN5mBfPMwFnB02JFtt1prgnoTp21/ajnMVEW9m9pspWsCH2GxI7NEVXUcgGE
OUwyv7D4dpoECMG2IsvF8whv5vaT/We6x+7rGSmoSqzb5BypzChb3Sg4NtO5fN6URAQDWJeJSdUO
7ClqH6X0s17rxtSSW4NXtFq2+Ce7MK0hSdYZJHfsegoXyxqtkL39IUBRiTw/FDGt8TxFBl7REGxj
i6Bg8oKslkf/4AEJZeOLYEENaHOdwaun7VgcBe6ZAPl6ZAoOPzYADRHa9xGZ/nhqBBLQAqRD+mip
Ab1K2PEViFEErorYPw5aD6rDnHIz+FFTywBHBAnNI0GGsWndtlxCqyFzf+8+wzOj8llRqQ2WCvRe
5WZ5AlJiJzXv3xmzaYxwjGKILR2woY30lYTUoJac4bQNadMaRq90w40hE5jTvWcdgbj2tGwpUaj3
skIGmJzmMOmZTBkaxM70CSLAYpp87ImHX7pn3yHGpBOdWD0RS6Ds2QV/70Pim7RAY8tnoDkI0VXg
T17b0ZmPxrf6bc6KNIco6s26hpt7wjx7X2Pl8DcOCJm0srmd6Eyp/Xv11FKknRmAim8RPA4+3tmY
feNJAr1TRcGan65fnftemY+cDSS5dAdMQz8XLHq+tB5NuKxrpawGj4Pg7WGYXdgDml0u3w5ZgnHg
Z0WtCUVOnUBdV3SrWAFKrVmVcvWtVIQzdNrJNrBBCsJd/cBHEdaYmMyr1NYhCKKAg7+8XxdZ2+XB
4RXJePevn4/HVMfCpEMQAp+5KmkBSfdTED68Clz3JYMzJHql4rmeXbS3Uv1jUT14IjiM6x86069b
Z1VSX60Jn2yM5PWZiXHyaKEojZgJ7DvpDTyadHAxIdhF1D0EIMNuQW7xPUSl+ttkoTf2DLKVxRJz
GnZXjHHzGrMiA94nFsw4Mo8InDPLiKkqlP1nGw+dyx/bRNLJgyyaMIYfhk+OGLZdv6HgpQ06MCPX
+VET4feeg0MVpo3AE6tKYHvgavu7aafhPINCFg0eERx22ewkMn7hxm4w+H77MofA9qh8sacDfSY9
0efZuHR5IYzt4HJcVts34CTDZtjHVeX0rg1HNSCLhtIC9fsw2LxFky/3XuVcDvcmlqp6ejUEfZpd
37EC2Fa/FohBVwDypPqyQnMxIWGG89JBpx2CKI+1uG6H1fyPOAvPjfRQsspCT6yqNDniMraPvm1i
KWl040MSWMHxvUuIGNGftnlrI4jOWhYSbTRMLSOCKvpRhlaUKd0aG9joGAhOsVbbHPxl2MvnF5RX
yUv4gYDcKi6muCXmwXOcb54m268Es2D8obqiZwUM8Ka7ngFeXxPzLL2eoAWOOGhs/oW7gkVJ5baf
FhlBavMSHuMAoJ0fjO961n6z2PK8eUbagwNYA9OGqw47Iy5e6cogw2jVhSgfUvFWWA4YdZa6U8X9
BX9RXgpmgJoxKH/yjwssfO3qbWfQT8rmrVXOKzMrghRNkp+1drIBrrPUZr4jXOdYUaDtKZT3Agys
yDCWyIntMn2q5zge1blZG4dyia/1N91L0D8frLNvIerpqFMAxDwiJLU3VVagZn3LMutV6x8yldaf
btCfGjSRAMY3C6mr7GEq77Z9bb4XLTuQmxrGAzn8elK0InOFMI8if1LBqy8wah0HVVNUFa4Kk0Cn
pnEdsjZtbGUF5p0MOhXMwWNIf8ze6W5CABOYiKB+5TyMWPFiwM18nxnMe+Nl0LvR4Uv79RXdmral
gtoxIyX+4NYm16YcaJ5gnXe3hS/smstikrIU8XkMskJdm701CY3C15eg7FIhuKA9dfMtDms/OlN6
9ICz1gJyVfu0NA9r0dL0LKR4sUHYGEdYb+06oDZw2B0bJb22DsSLMvlxKmaHsqH3B2XWiZ5iLeau
ji+wgp0nwPt3vcXYAUV00y4oiWWlT3R2Xk8pbaDGYSLJCGqePgy6CCY0YwTtQnNwX30UTiq3bY5C
3ExoZQA5QgPHyYRyB5vsV2mjbPUheHUqqNUhiVutzZvpmUMY8XMSt7S3Zc7vK2qLWJfXrnPTBbFh
K/uQGMCpBUWxoR6yliB04PWKJzuA95q+Q5yb3QR0HIc/fM3TZa/ymlKGR86vn9Kllq2+E7TxJAo1
bI/mYsSwaLtMzD0Gwmpb0irOvhIbYea7voti13c8jm2muXyLUTMxNtfDswC2Ive6oI2LKN6Sog6b
zNp6SMZOpVdJ35H8KCHbN9WGLI9s4rTevZgNd1BBTVlXDJMtY7i+3MRBFmiOB9Ytj8duoCAtfNmT
iS5TIR16NRCFgT99bc61IpDyCtpU0K6ZDh2Tn8EwIEczuCzXBHnae99QtdsSfg3yn0eEnbaxepJp
zRQIKRv1GEHYi+AWq1hN1zg/7YUVubz9FTWgA+wa21yGXKUIf48GTI7JT30fuHfDQOlOBxmo3PP3
y9BxnJp2TRFZj0UsveMePY9A40VR7L6QJ9BofqMT/UnpfvLgity2FTngbUGsmxqAkIDXNoi3Dfrn
XQDquJa3103btyAzT4sg03gkbjNHXTxdeq78gRb+dMtyUzqrvV3XdHyKdtC7eG6IhKsvw5U5EV56
aMw6ticAONwALt5fzbXeXEhwT276QN/yowxTDK8jDU1vIcfQEdQ+QoGdSIuWeZN3/uiJJ5p1N95T
d7U4O+gpxF8sKVMBNOVb2wkuGna36l76dq8VKyOuJFBDLmqH8Zy0QNgS6tWvux0AfRWRYBbof8nY
/ZY60BG1K0UrvSChOEHMHXYMMuHlnYzgvkMP/HmHlw5EzydF6SNAEK+ZZfW/0uUiqeQxn2386jCx
2ryp4kxzP4bboyZLHDHpnNyZPb7seCGNLYNT10ncaCgPuwQxbmLhvD1Ee/t42MQognwYVaBX8mZv
twZZjc4ndVkYn1Ooof23b4N1fwu1nkWkJXoL1narn1w78HrH2pRUAacI5stsyResMfxsUqw3AxeE
mccoyKOVSkPeEp/caNLZShVYkXA1EBlxCOA4CKqaeA2BEI7fi69HU+kI5qGnG5wlKXcHbfZ5Nivc
/rygzjR+4+jIv9T5DNpfq3IE2GeNGN1Fv6iG2Lz5fRjxIaYvJ1ja2HKyPn7Ui4IrfLtyAQHRzoDT
ZORUkIFP++/iG9Ct07qt2QIR4fBO4k5VtByY2ehFb3NmPymoyxCYRr6Ifo4WhTQbvbXPBl9THt6u
1HLZ5GuRLEKfJayWfBYYCiXtxl7Gkrfnibi0GWJhEh9DY6ZuIwMRqwAJbULeIDPa8b2HAVTPi3ws
5tcMQSZGvFRor+xhU5uNUGA/nkqACTtfS+p1NoyEZw3m1ZbHDLMS5NaUymT96CaZOXDFZK4spSw/
YtkzWIbqRtODtdjWLQnAgQhOJZROZWR10aFwSCJ/1qPWpaCVoknJ3wNH0ZFQxsLg/kysu0WNJva1
tXl15WROYurVUk122z/RkCZQaYxufgJyfH5Ok3RMzt98/4tGaUytu3CT4OIyQFyQ5AYZXyp+NM0C
oIla4GGUTrMx9JtO1hu099bwuX5uHlqHmwaZtLQzkBfSfGQE+GvJ4b7aPZ4PczGsXI/MhmiQgXQg
HNDWSsPgkIbtXejydWjbwYOgIWejXMsEOAKJJfY/fyDfgsD2YLODwEktmTO7x2WxYbpDzhF+J0lf
bpOZIs8GeVOO/ExecvWprhnBLyXmng+yycyGrkwR8nZAJEKbF4sgOfAGOmdQEwVCtT7Y5N/DOAP2
uGD6R0r8Y6pmGz6B/Y9CuxIU7cBA4TX+z61vBjJ2K+nA5nwXIyOUhlHroQCcINGNIXtBjdB2G3IV
brs63fW5w4eY0EML/nqqWZvylYSDqa2tIwEhxYBhAnGKGFwVS4fgGVE+w36wl4SsjE9XTd+Cnrq8
hHJO0ZVYLm83KR1rOse3hbG7cBz+ROnKsVh751zstuHxN/9/hTYtt/6uG+dNZUW5VrJ9OG1mnNPh
LN57G6vA7yBfhQnRUH9rwKqmRTakATmYzrCW1TOynGfjWhkjo9suCDQEc4M4GmQMs++aet74as0M
KRJTCvKFrd9d1KliTTbboOKErhiuyl8TyE/tzGLqgQHrIUT35cmBcUJbEM3yMIVBpxR+MnRkKhiv
kjmEEED2MPLiL8z0UpTQfJ5ArxyjGM0tppqu+3FMsakxsJhW8EziG5WH5E+x6jN1diLwbkESHylX
v09TlOQN0genR0w+vu9IWQO6IekZ8fRJZIn8NjC9ZIYOe17TtiFeNb5WRdQ7EpYj8V8aiiy6r67G
zQir+C4NVRrvXXgCWpuLYraddzZr4E5S4WsCrr9AEge3dGvSvvVXu6VZuCc/3en96JKhUXLmxvA9
+GyHjpqADPwdK6e7xol3zEvnusgS6O7V+eLSHQCZj5xs9ElEG36TOijGQkUR2ham+1Cgzu3eG/Mk
REXDvMvSKSxh9C1x1/1b0gE/wS7a69NmnvqmYkElw+H3GRCu7E3br5Ssx94XPPuCH+MYxlpRdTZl
MVcibMng+XxegFgQE7zbnba+6OOwqq3ZAFyMRJuuU5l/32wr+qj780U8ittIi8nyp064UcFdxkEF
ZWQg7ZdQJaRmmUO1VFyoUkzvj3h6KRw083zC4cVL1e+MZVPzH8JuXQbjP7UEgOSyjN7Y15bepKzF
Nb+RmnKKUUMPBcB8pr9FFDb8NTI34FPffwniYBvYO3RrvpVXSTcf5QZazM4lvk0LIk3+yTRgkHFp
dk9GeXx/vJ1O6+AmWaaD0p6C3ofmN5amzpyEmHm32ZKc4C2D4mEquIej+o5hACmCLtW2y5vbePKP
8QqmZh6D4CoZsGyoOsDYNfHvT0oA0wGEkZcEVVfAzLemm0IWB4xL7L2bGJoLXYYdI2Wnps1cofsV
VH18Y45AbvsoDjtASkZL0AxxQKz1/QL0Sr05zq0ybBNraFVfL0MDKbbMV7D/mnL5Wx4xnITM4fGc
20UQlHYGS4m4Y9SNxi10B6TizfLCZKQ863WQg9NvK0l/3/igVJ8/BiQo/FQ8s9/P0YKMUthyOpzm
aJemMN1Gti/x9k88GIemImxR0G+teAAXj5PnhyttE7I0P4M8gTRAEnCSE771LUXhOgWx77XU2UVW
BIox3epcEZFlSmVqtspx/klTVXu6TtWhmO3C6FQ/79idgcSyjUECVX8E5L+JVuBnfssnkGm9X5qz
Mjo5x8pf8lcTvb6qQHCpr2siicC+NCU58uxKv6Khn5YUxxuAgOYDu+TxS4Ylnbvsb5TMIXU8iE5K
P8C2fZtx25cQ+K+vsXR5tvKNliNv/H+RyJSLOnA1wUozk1AgApLTtJ6tMsbdEPpziEoJq3aEStDF
/I9B9kU3mZllddhM5P6yXjYDBbviAvU5G9mP4uBCPzTah1eWvUdRFavtkrC3HYrLdfrv+UxsdFoX
ubHcsWoBUa0nq4crNh/gDhzpBxCnAxUOOPvzte19jUxyOFaua1DLVnW7pKfH0zmwvpJlAjRnlcs6
Wyeo0ns8DvmucHr8DCxvt0cKeaO1Y7LaeVZV4PR5yA/ZWFHXQzKs2JsftBuaBVg2S9hp7Xj0z6ae
mA8hn6Inq9NzZVHyVTbUuW2f/hxTjh8HknuQkkdg2TIyTqRtLfbpnpzEzTcqOG8TgM6JserU81FS
3S4ahzg3KbGwBlZAQZHiVtSFSbEUPobdkXq1TV8Q79mOlpCbqJCJhrqzU1KOb6AAys3ydKtuVSzo
+g5EQDFXtUbhyE65dfQ4gARBTkaxE3PvUitEgW70N18P9VSBS2a3qENpsaPpyWHx59JcY2rvKwNM
pwMonZPvlO3Eau9nVBT60ck40YoQVZlvhwr/U4lOiJ2tGrTNm5+ctH1doTRwKY1pT6LgYeRGkDG2
HN4uaEsXkgGIXE/en25YcY00kpj9bAZdEe7u7iJJyKY0lAtgJVkq7PiL90QjtrtPlSZo6bbl1sZ2
sPbmKJO+cELi06QiLnhX5jxbsVpR36jX04iLELms5F3Map0gNZvinFbFpeXqaqb/eVh5hsvPKVFH
TUsHkI+f369910ujZ5zaKlWJpJfHz3YHfrMyFo+Lb5Q22BT9yRSEyz32L4C42mdIbIRZWyXj6jDO
irwAfuPq2LhkC9O3e/+HRR74l1JbZ5Ya1iKnmK2zyuuNODs3O0IdxP++LDM1WZ8JdD48vw24eUbL
vnKvYxptyRST/o1v/mo8CIVt9G1YGWzN8FiwSo+NwbQhYU9HtTf2tldOMXFgid+OARp3nDftxde5
W9pI4PvVIzXWBc2Pd39pY2c7idkfnL8jEtYXFOg5i9Ru84aSCvYuQwr0ptDNWr69SoARb8stxQ6f
r26JXRB31aHS1ukxMqS5iqCuWKp+zy1HxV6nbQSGoq7cKklPrXbwGJ9kvLrsmf4kLH4xbbKTxyBG
v2OFo72O+IRPTQHFJ+mrpmpv7q/qz/lHQaXa4H99wciT9jkN0Mzy6ww9JZK750MxfUDkYMKw8rFZ
Be+hqa/PoDMkwHXgeBTPxv/VinBor2J/pwByDI/yB22ODiG7/e/6y6pjZKnGzh4rzi5BtU9RPSkq
nOh9NEO48W/oiWVFf/72of22mb4lA680HwFwOROPCuCTX++1gngYntKzSXKvKluxKvfWFyGSg+yc
dJWSMRIdFQiVrYnccU4ds9zSPuw3lik1nOD1miS+f8H/GCrbb0G268ij7hgorPzw0OLxhbmO4s3Q
j95n4DKE7MMfrvujqSwiD5VYTd5eatMbyUh1kn6Rqp+OPInrm9dzz9xXs8tAWrrrV0l3xq6scqRw
dzf/oph2c/l6lpeUHKawppbV7OUPXjW4X4hQ07aByj5w3zMk2zhfCWWKEFLtgPZ5qLB6CYVEqw8G
QMq8H+c/t5bEmYjSAJf3vDi7z5DnXbeiyj128VAt2RUsBRUz/5mFiLUvVeijVxtR1CIdbB3dEn6B
Bja9Do3GfcpcBinWBqc2G+lrXrCj8OSsX4PGK95Zi2vEk4AX22KZc8JZHcf9KwuZfnD9sOPPrOFc
CpyAY7ARBiXfemMV/TZU/IhhJaDMBH4RHDnX8CKE+aNc9gL7IF8+3sN9CSaNkMTUKwv/m4kBqOLI
UMdKursOncjm5Fodjbd1T13TVGkScSrjHNl2Mrnwhv8J5C8MBWFFcsaqy2tEBHIDuM6N9qLfR81F
Mr/iq3uXS/dufYaN2f6K75AKYrwRAo/tfQSq4zpU6owu2v68ORhMKpvE6zaHfmf1RPAX06XZbvrE
cRap4ccMRsAkBovs3UdmtHfqeZoe6TF9/agqUyiPFsfpQwMluZiVMMocbajcrOawP/0VMr5I8Hop
dhSYFnHBp2iTMo39VZaIn5rgZLmV/qB8AbdIqga+kBTUHZ84aqeC/5ML7gPT5+i/0KiHw8EoMu2g
sZ03M6DZKsHuJAl4g3964ic1bWbEMh6HVZrQ23ZmGQnYlqIqLLpJ1sV64og8pujWEavPqFvGjyl3
8k3Cv0FaW/Zp10ZfQfGhJTc+7vfFb3zOA0y9UYRk5UHHOxzq3mh5Fv8cO5rko0Azgflt1oSF+VHF
P/HG3aXdEHUjh9HngAHCb1e3S2a/tEL4bsHSj+XVzOUVCGXq9Afhowjnoem63KoJEmWtASrsEMys
d42DlcyQP1ELknQN3GkI/SmzqUH3rALV8qMizUY8yVlCmdHzNKaB9ScAfm1x46RT8Jhx02xT5JPw
Qu3PIJJUn6niBYlI2QFTDehqwZt5GNnVAb5wQBNyTAwDIoFl9ienvZucVmpuvjIv/lEf3TUy/3BD
DaxEFk2+rj2Di3pfHXzEqWQEpj+qan3qiylDG1Q8Pa8DlFvk5ynK2X5RkTPPGrx8uuHo07oErK8U
miCcK8FjXbcxgRUjm+0nFyGROoKmAg3sIp6AjPcyfOXhPLdpa+vIANw0V3WOoM24YyOW20xr9KOe
4desLvsbOkeaPdRz2CfxlPgD/PGyfvy44my9trm0x7djtnVxPIPquJVb6qhQzwPpBPXvpHnw7EHH
tuEElzoHUrFscZJasZ+nTmfOtdbaw/dkoEiU+shTwRjy8dPKW9d5ysI846XqeJQeiuXUapNucrEo
WzuOJ7+H9kxSWZg12S2MvLaTM4yvOtMoOd3Dr4JNkdormU5tBAiHLxnstnDfQ4jkAnBbcH7Gkiqi
wlAfbTV0bEEiW5LUXy2zAqkePvextA/UXVeBG9nBcRyhFq62KFSqG2dCrVG4Dj6dH0YKSCmz3hb8
DOCxObLxDX8R9EYQvPGqpEK8F/1tX2WEwb8gHtjJMVDtVZdBDFlLCgakjt34TanR/MHNJy5yN1tj
ZsdqY6ssNyTjobJu+VI2LG1IJRrRJ0H71Nv2Ob+82zxHU5NguxplUYmRIklpY4XI7q58aqlMc13a
ZiJ8NcOmxZQ1E9b+0fMDtQh7Cv/Ljjt9rB4BrY57AapzvV9nUnGjB7je+r3doDBxeaf1draGYOSM
jgkmqueLczmekui/EqZcsTeh+gMsPrxG4aBUqG6cy2hTAlancBxP+R4r6jX5p1ZQzwpRZhhCszv5
FB8BF13PztFq1jWnwehi8Rbpfa8R+8ENbmeFqa0WB7kz+TXvEanNdbZ6GlOGIxy5NTiPrQgbGSk5
FxesoHUnPEJpG3J8nhM0nrVmKsWs5uB200tvIhjNlUCaTzSKIdXzDFhhtpMd4r0P2d8cUQx10iy4
ec0nbT7MP5GK0FAt3QRP8gC+o2b//qTVLpm1fhmxKZIAMppVylzNho7egW/Rwk/w+CzQ/N877mJS
o1fTPaXM5KOORgPWl0UInsLNniOjPjjkKNeVrt1e6ziiuYRZ0qrFoRaCASAtsJYJTqVCGLWSN6cA
nmUe58hPpGzIdrfKjeOcQLQCGdph1UEar3WXCQrLXzuSCaMuu5G0IZHI9WcNbe7A1oIlieScUD+z
k3qw+2+6lgJ6RQBXNjCvkZT9vuZY1dDzam/vvnw4a3Dcwx/DZ6ILDe1bsSElDWOXOCWLH3UqNZhe
JWaPKzgd6/FPTvevMlS6tFG/UbeqvRGNgoVgkd/oq+RKUo8pdJikpfXEc2SSbN2yHAAOkkclYFpI
TXtrZBWyolN4c6M78hnkZZjxnAHb2x7Hwan7TkAFqt3uHVim/yZDTqyqnWJ+9i4Y+EqMg94rvmkE
5RJM5CQ53Wo049n5zxpU8XFX44iDxxl1/WTiq7tPsLJxtWE89/5tDBx+hwwQDF8BknvpLA1yVRre
UzMhsd+v69Bj4qTr21QS1Ae6HXHijMsDqvTHYJeWKpTTz5d/sc1i+1irQOF+fYpf4vvwudnNURXA
pwbHzsianQqlQbZuwvWvr7lES9JzmWjaJC5K4eu+5SJ9rGY99Dd9QvTPXdqrCqeRrrH8PG2aT95f
CgjUZa1Mb4pZUTQSSp2VQj4VTqFFLHdWo09joy77Gb7028jbwyT3BQmgARAZ2OW7ZjlvDEMXE4RV
oMHhZaITaA55MSfPQ1y/mpA1CdjhifuiggvNPOovbixdz/M8D2bJWwN7FSIsOovkfyZz67gAXVAX
Qz028s6h82fdfZYntDzc8aBl4CH4CGUR+OwMLVYEay54BpOGhy/GX+Tzpn3xeB4Op7KA2GaVYs5u
mNNYBkji0zLuKgASBhVfiOIBpLZTr/hjoWUFxpjd3OP5r9H9Q1ztkDpp+UP1s/5zakYSfaw2G8kz
xSZSlTZWSJeAQGc9tzfasCmhDdReLxSvp740RN1j572p5yLvTW2PBmktHbCrimu4JOp98iqO0c1z
MaWsDgsnfsoChW/qsF+G/JT4qDehCiDCAxm0NaDjXpzJsQ2UouyaD1QO+ShBKhS7Rxa7HHxr7FpK
/wjQVqBaljveVTqF5XKM3adreaxYam8h2/AMTVDMVc1h95WOoHeu79V5WzghVci5iI/3shuVa+rV
Ol+MYm35QV/9AI9Jr3e5yrNJs7O4T7ylMdTumrAo6XQVrsklFZPEcxUQ/yzLh/wkJpbKIZJq17NQ
vZPFxWdUc3EbMrbc2ohDle2s5SpBBcQ2vz69Fu2nMILBsv6uMpHVM03elhcb7PHPxzm+3GVRT/lA
EgcxJXjV0f+tLW9TbWnZyKBxxqg/H5qcM+zQBFhdZxdUilew0L89XN5WpP/T0KKXJEsLPFb6/vka
LHmnThtsNPM62bQcHSvnCxcQOc6fpjWYSpaoX62o8s55G1OvMw1biSUyVOQ9EU9yCXWUcdF2Q4Mn
lUOwC3t0ME54FgHs1YFgqb85vO6X9bhL7t+TLfev6eJF9jhoFndQW3QO1wDm0RaU5hlHCgEgwMpC
5TeAR/xQ5m/820WlZCpIe/4u7bx4Fculwk/fIVDmliWhxiampFuokyK+ash76ldBswtS2W0Z68XS
pamLYZdQlB/XmFg5qig1dl8mnxC9lgek2juoGGaOIKuLGZ080LsZHau0UYRwTHJLQzULf7comXQq
96Rgxb3rgBtRm4/zjsEahJboywQtKg+NX1B1DmFkQwf8g1Pm08F43vceonu8xgXDtWPWoG5M1rTd
a4+VGLQS8OI/AozbLhH6Z8C+UQEynGAdDNYadNet4XJTiq/fH4xmMRbv+wuJB4jNCkXKHvrbHIuG
Aey22H45fJFz4lLtMv+s4928uH0fFYt3WnOa3BQmmAxhSCJix7ITD+YdBvVuvFAxAByMcAHO7L3M
vyvtOEcOXnYLG7+cMduMpkFCetxaevbf4TteIG+FxUUFOnwHor4ojKRRI4iTcdJOAMcTOMyZZku6
PP2QxKOMW1879YJ2Sqj4oU5pKrdLMLmxtwPEkUsQI7FqJAivWTRm9E4q4QsZ1T30OHhcl6sqUXZA
aOpEC71gsgH36KGM+b/oASGj85psM5CzHvfa92BqF9YHPhK0qohUSvcakWrYhIramx1DZLb9eE2W
ZDO46sY8yEncU83Z2/A8rQEwQTawUIiAIjyAa2dFxj0FQaWhdENlwcAOtaQZuM9UbV97asXyxTum
rwQGoEHTeWX3PJrYXLzlRYzcbRhNW/QqcRRAL4jrjbCRjyhTAncNpTo/nNeIB+/0vpoqBX9k2Ws0
6buYkrUBh+WQTwgF5IhrnBsSLtrCSg9k7x5o+R4Ot/A+8+Gg93JPCyP52ikUzwVAIq9QSpzdF4jL
B6EVIrH5vxFwGI7keIkqNsicD6jC05i7gU2Ls8svBNKTNLtd2ggST9d4BsK4KQdzGD8JUIYO5+i5
GUi0+NG4XUOS3alBDbrwt61KQQo52PJcOZIZFRpuFqFWXsllDgIUIhInlPwEvctBFJ045sg06JTm
u8dnF4OwPsA1kejFkI/Qg03F529hcwF79VBHmzVpAeD+pLCiHkzr4mBmx38qIksUN2B8ulC7oNKv
hzZi+NLJIT/BE7egjpgK4fB4sFpNyWnL5g/+1t+3/jYE7ZMXrDjoRhIDM6B9zPCzWwIyDX31IUSr
rS436GRX0Xdb9+nQxd8YfV8SlMvEpm+ihknU31RjbPJQuoCu7ufOkrIhnsadYfWzRvi+9ryWdH+/
9uFLx8nJBKmnRyM046UA94pu4n4f43H0vHCg+pJ0GupGmCU/WriR5qIgEYr/T0M/FIgeTMndEfN+
hUEHkTJUTJwDVtp7LCAtETAxMkpixnCtSqGNu0UJ/MEuJ0R2lTUuQCZcmBVrR2deYnyeDrvAhx9w
blwSLLONDo+GPyOfKa/0KoolEuDSemHcqylk3Y/cHely8lx/jAz/XeHBJNfYUqLd1xIA+nTuB6Nd
Hb3wfo7PZ+T7yGCVkiUgKRWx+Qcl3XCPZrCsf6c6rN4/pXq+YGwAQ5s0O0KUV2RvbeMxKxI7MHXg
2JuiRGzibCqPAXvTTHUNP5FSGqB16aBrP3MNtW+4Q4696MflVe9bBY+kRB3a+CKQo8AbLLg2kIaQ
bBlKYmU4iPB9Y+wmRUTkj4aRbY14HWFzSGWZo+gIlCsTLkyjT4gpcUGPiit8mJj1NkTUfBs7fDR+
wiYGia7Ue0CHBqllyu1uwh57KW8cnCDLmH1yEsyfEhIxjFf7oaVgPe9gD7QEBWG+UwKgaeC4D49+
nXD5eltMLnLoPz5iKd32oJV+HFQ6yE1CnAaY/hKzcPn18WScQFp3hrXmgk9W+SVP1M75rE20F8Bu
QTk2Vb+1Svfzbj7TFcTPl0VfM/OsUKlR5GJhCi/OlCctEKxyYLsU9JSDQ20rb4xBP9738Jw5ue+7
vqpKIFT24nb+kxgYLF8wuQ/vv0KBBxqWDtr88REPwjcSPar5C95jf/P611Zifr6wVgtmoefndZC3
RFNgwThmpUEjIpt+sQNXB9oxYtRAXzj+jkXaGcEzRMbpkfFa7bZH9/MUJSpijaDj3AMdxWCzjHU0
APBha4r3j65HX8BeaBtIVY1ASGw1TWPkTZdj99tY+lXujuN3p4c6+1uBm2X24D+GbB05unaX54zG
t3qois1QflBQP9CkqLJU01VS1BK/dOUwpe5BbRg3vDt7Uba2nAqrgqqKWNd42E75OUGCDYtbR8OM
f+q5hpwn3sjsCzJu+yB77KduFPqUBzEaI5FIoOrzYw4uHpGobZVtAzz+iRQZVtv3C2zxvpdMa+p/
4RJADmEGeAf3QPWVf1XuirqUARIfagLXKnVoJ5ib9oEuiLu4DJ7EeLhmvZ4dEDz+soSspksU45dd
JDgopLsYHptLW+ElGq+Z1RVtEwqlr1HqPtIQ1W9GdHdUSJSFsHvQ7gh1r3i86oXNJPFUvUqjUv/x
RqJug3eKJG++y8Ua2Yb9LeSVnMQionDKWwUENbAC/QcXN11pu6lQLq0vVPpjaGlZF2pQjC0GFBxQ
7KIP2Ha09mwyBvT1SSiWDXd8hgAXvuBNtVqLzX4d59EvKPUw4ybmUjOlCznz4lCcbq3OTpFgtPZk
LyuBeREoLmxKLe+TvM7z0D0aI+uYBJ1Gbk1s6WbKuaIpIE19cdGECH7EDiFb11Qej8jE7sJOVnqa
iwPOQoz2ylLrXsNUmHq1IAZ+FSOYHizQQs/Yjckl7yy8NP9rd14LiTaRHxtHKPHiCVGYM8zEXbC/
+yo9eEhNCYRv6HbLJbVJjVPDils/wT09ZoTwISBLSyTUIhjdJc6PZJWOcHZT4yHdM+T9K2st2x9Z
iZ4ZBHmTFnMgvt9y1mkk14F3w5NsvA8OGCuJmgQAJTzWN06PZJ5wPTqE+23BeC4T3pgriRl6tqLp
fzVTTJGdq9kMKE4fzLf3DCX8P+hHqaw43pKtLKRW1Q1FINpZXqVPLBt6CADKhzgfNj62FN7B96Ag
eBxX5DygMN9D1JayQXks7uqG/IzjthWHMyZnl022XOhC0sTzxHGFOwd1BucqznZ2A/aJcTZsVXUl
XBY1TidKCp/uZweXNjyzbnE+1bxBl7o6uesFHLwdeZAqsjL2IKwGZW0cOepKUvkS7Eq4tbqEFDTE
gvLWcF5u3lRYuvi8o9/9dQ/1aMnMuXeK1p+atau76WnHf0l/66PnwXulaxjo8dC7zHAF7fjF6Meg
UYTQNgT/aW0rKBB9KNMFSh3R5AZsWdKGT4txUaiy1s3dwVpHLUsJY4B9CeRVzP5znA3NGALnhgNn
6Qt358dtlrKMz6UIgeat5AYdVLi64jNIUA7ROApWe+ByqW2MgnwlbK42cnARMEuIffrmq/zNXNa7
/Q4zByF+xoXKH+89Udth6oXLAsGAh9KkmUTOzUJ8yaxcgNn97wieFXfh8lv00QU/J4z2tUcvtMoS
z62s5YpKxngGII7LTKJFhLiyuYYM0z8iazBxm/+GpYgmgKgh+nBEBqr3wAwXxwuGAG7uRN4GAnw+
lyevaOQHS/WJESA8lvGNxNwJnV4+6oV6tCO0hWXqbCXD1h9SMDIDVYmmDMIaYG4EnN6cWdftg22P
WeRO5ZeKpPSz+xOTZsXV9bNP1RzDs+0fPg48g3uzMpgAeKMHPJBhL250bcSEOH2gW0p3LrtLQzD3
bcx+wb/QgH0tKVrY/1rErw2oTrj31mRXpt8IiKRxQ5akyEk/Ntl9kDPkv7Xb0Ax+sou0sXhVHGGh
hfAkftmD9gO1ujdgPdLYx1Lg6pGyLP4E0PXVlUg2XAiToyMrQcIAI1n4QXUuCkgef1KB1yAz0Md0
ggKPMWrshhNkq3NhubCsVaDwy7aDhNdyfbHBOKiK+Zzm77WmuHgopElmoRLnH6eaWAiWmZfIQqYv
3uBqDJd6gaOHEl8K10DUI0rnHdieTuWoT2MhuqhY6zyYbga/7auVQ4vmru0R+j9V4Wlfxgf/YG7V
urmj2qH28+xLxXMuNYLNM3oYM2UUmamMHN4xdrzm+4dWvOBHEWY3XFAExidCTAzwaUmkkfHTOlEL
ZVe/DwAEbIDsSyxkQrFGW9GNcLkqtoocQQdBI3Y6zdltzXWFPcKDvrXIEWcIW3y8INvEm2XxGvxJ
Kf3A8FnXVIgZQz8ywG+vMm6vvU4L8I2hUYf9UflfHRLiZT27breQExEvv3ukKymkfzH5khvlLVih
/urU5kgxFxhhvI+4bh3+lyln7oy2bwZWxmTZqAVrarHEu5BK/VNEXKAP5v+43bEEQna8XiMfyr4y
3X2KZlBeMWEoBr3kumRyGANuvUjXl55tl2bvPYIB0e5NoflvbX4y5AoHzQuiE34mEEUJpalD7zMV
jArWeshq9nz+0XUBJR1HUxb2+ZOTiNXG50no9VK22kYyZVdFHAasz5WJgC90ZhOX62Pm6IeaSQ7A
UsR+oBkMLhWTvROJpKFgxNhSWXtOas0H6tYrU5UPbpuQ6HCtWQ+5bBkzAgj6nSH4VQTQwVktKdOK
VoswCE9OLhMnwens0/8s4qWMR2OQEhmUnDlvHzt8UnqANCVq43Eo07dwb4sovGkO4wTwuvqfbIPs
ms3WeaxJAMqi5ZDdNBbV//ag5YMwUGmkkqdAvuLNTZ95PqSAh2sJdn+STP5eJ4aWIMFZhXS3hj43
gV7Sgi78DBJTFXLuuSqNSG/O+I33EFrep49eqayzOu7HSIS+PvhjX0YUCPJGF4sc+2OTWGMoOQAR
XHIjJtn28KCkfcAL+qXbz1kedbOOLKBKYkdTAPfsmASBAPCYJdFBXxsVg9b7RJ24e4JQ0qjodciD
c8v4JedaPJ/42vMNU+3I2ntmIb9VKqZXiAfJpGmMb2y+rStJfGXJW8H1bMkdwLazr2EgAcOVUll7
l0J2491ZiJZpPApn62KUHf9TiqqL4hm0ioLaG20hBgtW952ZKFbRDb0eQnO+SrGzQ51O2zyzfoks
tNhXLyqXKUrXVANkchEyzQUqY0G4sledfUljiMf4Zuw8U9RdDBPyoWBhcX/wy49UQIz0yUyPDEq2
28RplOS8tpUxKLoYmIi3E1lIkWEpU61P6g6zxAAhVWpaXd6zFKjYrz4g8tqWq2I6Ol/0MuzxeOtA
XcJ3XiX32rsTBdOZpkhbkZcptLdgKl9RXO4faZb8ZeqwRsd7HGCSXvxT7fDXvFjIjO8V+nFAPwMp
ieHa2Ua0qEiUoybBxForIwZvT1WysyKba24tlzEc/Rrb0ECxD99AoGCIRcvyG++ckte6f0rq8Bil
B8DZB4FIzcc1YQV7ztu1fa92on9vAQd8EFd+E+mU5a0KXq0LnP5R0TzLy9y6DyfIiMoiP8gCEN81
+rezRs6mEeuNq08EmtDyUniV4XlG/xemQETxa5MouZNojjYo3JFOI2z1ZaFOpETG4gz2SP8IZSlX
/HeYUAc9FcoYmtiTt8tLzOEAIOcUllscakLYePS1RC7w5BSilBqegOW4vWIcqSjzd+dPYREsQi4J
wsaSVr0G0xHv/iwF5FaEIZT7/ladzChT6Ge1d4OIjmd6lFzTIBEjSlhe/Fv1QlSxucREOmDROXRL
OxbnX2OmWa/MiML2EVqKasc28E914S1Ty7iVGDcQNZn/4rChjc9MOSP1C176Onh2MRfc+C850ccJ
2LT/qQpwAfFnrszJAOlYWjA7AOUQroH+Uo7ta4t99Pdef46smtLO3UsrCjA3Ke1hKEVQlNbwUW99
eP4Pxbg8/v++IGgwCGiRaYudC8XAlRl8RDiIqPh+i+iDR3Bvs86AwvfU3WHoFVaQ0E52N0KBe4RS
dd1N68kG8FtzrTnsEch2vnpBSOyeUyFFPCKkePWLxr2xTwdetWDxWRlbU5GsaWIml0Ty/kVwQG4T
2mVbwenvcgLasSV/mN6nphu+HT2SefHgNIodACWdsrcbStg2MOmwtGjh8lBV37s0H/H5bwSQ1xOO
8h2EmC7W0IqqKygS1wr6U1fxP7Al9Y+3XZpaTIljjQDpke337Zsfyp7Zey3e+xF93e5739Z1FlCE
zF7wTR9uFneppnNXOdGR7iCci7dVg1dLKU7z2eG53xA3iahvb4+1lk/HrUkK7LEI94hljTDVtshY
dRjNT/roemp/E8qjvpkk3adgSMXaj4h28w1fjI+bpW9GTJOYTi6U/oZLCG9p6oJ+pJQzz4EkUb87
jRmdxCYdMkYyXsqmgH3KJJ/7Z00IErluger7Ji9crktLf5csGzrWVjrGxyvYoFPHR9/OmtEz0o5Z
s6bfpYSFldjLeSNHx9VSskqCylfkEQZn/W/rAxX0Gq9l8WFzULrN2yZ38sUw1/mwNGg+av7LOzly
yJmipFNZDF0nfc892Bn6pjtJvz941LW7bCI5gXxOBW3b7wNzyWkOhecFsl7wP2eMYIbvhzo67nGr
ahsDxG9o0RAVBLW3BFrCyQNrIUd8fBSyuz76ogvQ5oICmR+hBDX4OzdgPvIvoBPonugYEB4QJBoC
ONKDUutmGvNiP2aGmVNU11ynGU7TG7A9G4+aI4YkjFhKcQnbZ0SSeUJIyT0CAP0gyC/G36Dv7wvI
CCPZpR8nyo2ChtoyGJsFAwmei3KFkiBlBi1nOzfe+VVDgrynWCQ88Diy5GMcaYBkFy2CiKwIjyNt
Dilz+uZxTlfYl7GShv+d9Mu7LH1bVgKszZD0m02p4m7Eqg/uSp8xFQ/0sJMxOJrv41wRU2OUkq7K
JCYplsUaNCZgdSiLPK7hXzld17PqhP11Qy2Cye/+i4WVH/XQ2Q9VbklhGttPulf+vlAclStLg1ek
w0ubf5Dj72B8ykT4TkPgw0p7x6flly1+q8KgPUIPpodqpRkc+zeZjSHrxQkjd9/dAaQo0s0KaOdb
US5xVQfLuT3kZsrBfSj7w4S3zrwalTectCknWDaMTEdIBP5oOl96a0h6lgKUcK30nIhFSqFaAl+v
rBPKvM/Kko2sF+NygiLCxQuxX8bVrBNXVyWEche43IT+AJXK/tUgXwwwI7nbzBB9iKAokCvupsxY
5OZAufCE/zi/ZalhwKN7Xi+op8cVMXNl5LmvIabbMIPOZRqpdQoSQvyLMUk0XZqNFeMJ7FCvbA4W
OeJZdoTg086BwL71XJj8j0qRzS1PhEJhuJ8s9FLxkUll1OeuBy6YTLbqRBa3aqM6ZHhr8ZIeE46N
X6FOpn6dIuCoE6x6qRhAPtewCkj1JhFIiejj0n7RSwOsK5RkhvbLM9oNHE3J3gEx404hq1s67BTE
XtJC6QYcnop2PP+VMINJa21tVVChDm4J+njmaEAmtuq9Mf6XfKDg8Z6MhOhf7BtvIKOvJi0+eRaj
JkhcKPSE9eZjBTxPE6vcFtkSzgKEteVlHgqf+jH8AiMD0jHysnNPQ7k97AiVd8VxTkXz0oymofbm
b8fody9qquj2o/c+NEwBckyv+Ul4u7Vgn5WaPvXRtiKlZi/nFn6Ihl4kn3CX8XPTZi/aG1vAL9Wm
l3opJ0DCoGZk4UFY9ot6Giq9xb68Ajo+5Ipf1SgYIMRG/aG5v29bj9DTnfjeewv5l0/KPKVm1oPL
9YtT9vFwHh/wUaMbMynkgWOmOu5MlUjhRPT5TLM7V7g51PuwXSZL+cwLSNPH2mw8nuJV1pB5o1W7
dcVAUvTU2S2C9/SDo8XAqErx8uoD9qVEKy/C2y8lPDhDIfWw13DpKGdOb/vIFL0ePByVq+RBDnts
MoA93OLiFrvXGKf00oKZm1mj0ieMiMtsQs9ITSmGzhvfRFKjnjAXqBR4en7eayRMwbsmFzMEIMkS
ef0+BiQ1rsRuPqHt2LVpAfHPV1VwIg5sFvjWcIAf8tA6hPcdX4+92RgEtbgMMWW6jaK13yRFpn9K
+M8XbkBjN/GWrB9MNwYQ/zp5nBmV/ZZCWNQHla0Rgx/alIqbZiLTDyQKViS8qdF52t+8wioZXQMd
gdiGB77J74Kue3wQSocu3izYVZcXlkyl0SM0c+9zQYik+vzQg48TNx2sV/k+NRV/dXvmyHR9Wkxs
H/xmdluksEbTDDLwXP7qgdV6qNCMXZ1np9tpULqvGlNaD9Gk/mej2G6oZTdNj9B6VHMWY6DRArRT
d7NS4SvYbG1SGOQ0evzR2FTdMZz69qShrQHeqXqfQX1kN+WuIz4b3PqmkfI3z3UGpzgSvQUlhgQ6
r/0OknVnkcX0qbFm8RVua/Nct8blKvHDMP6sfYuWBNu9MLAPk0lBXon3PFZnjrVyc37n7pS5OIui
0pZmgTI5Rm/PzYCC+kAr+rScjy/T9HrKt7en9bZPuoQxhLp/G9SLupNJqt5OKYqsTJJSYe3qc8Ag
luDW/C5f5N3BkEttSWjpb3Fnplp58JINNusxNKaXSSwrRA0esd6WxxAdY6xMEQ3IkOSu5UTiltW/
2TmTR0+lJI36s5VgaFnnxfryQGPvx5UKlOYfnC54G0AsvRrsokhVIEvNjd1oXVpK93MnzfvIxYtd
XIS5Z+U/DUBUBX7O6AdLENYJM9jyCmN8qQl0fW5zWPfymG3GV+sR73YY98DuCPC7OjW6W3luNgRG
eqrjGFbRtsRrueoHIc6NvxLGpT/nC1s1Pc2JawwRiGrzIvnvgG5yTM/5Z7N19Oj2qNH9xu8zTQe7
EvHxptMa434gHSzTEykvySL7FqdzPjbeklSVPgTGcdh3UFSgCDpts/VnO2/4cxzXB8O4lK4POLmi
oSiakrXCGq/YEaaP4g5FZifbSrHeS4aHtn1Dz1qmNfdVy+xVx6VYOHXQ5i7xREQlZOD/UbelvPTv
31kYxihn/0w6/nkOlAKCjw1VOxKKFs2YoebH5IZ21REkAtmo+WMZHcKj4coSYWAuk4TXRd81/agl
sGMdSbwoo+0+IbzjT90bJ2b7r+MP7vMTLRNEY+9H8GX2BxtEGNrLvWTwlKZHopAyKy4sHm26Pfkx
G/EeHDyaB+oA7UwP/wh7HLfvqI5HVQMNyIApiyUGs1Llt3iSyymigQ7l/EjXud/t/4OVp30Yy+vX
r4Imke7CoUhoM0M83RSYOWJuq8l5f/LZA+B+NzQFK347Tt+79ka8Kw7tNWsUu+1WhX5ZNpyVQzTO
A8dTGEsmJ5t3Iwf4Mke7EYQuJnl7h1UrRV3gksK3BQmxpmYwnivxzAnlMkxfZPmoOUe0WBopctvn
fJmZdnJIs9sXSOV1IAviotocF0inOx0eX2tNt3uXia3x7Uw/Tujnf8epcGBvqGs08/8u4kX1USpx
giqaLc4nDvKG9ZPhL1xG3+ZgEYxd6Eriw3RqVFK9KRiCOOIfZInFZj24MYwjviva9jvWRaDf37g+
CUkbIYLRNEpff6OYNLVXkmSWnlqSBHHtzErDPLNB4YhdU68nGqqoaiW1uV4GWdF+feurkRhVQBNr
MAN+XlLLp7FXBgl/AW7krx0EdHeqgGscOSjhN5ffXSJa4yQRjfqnjEMgovWgp4YMj8qDjT42zVk/
xYOVcVsX08PegObMrjbV5Auw5tGdn/qNyOGRHbwgUOswol25bSx7OwPkZFon/DJMrypp+/AtOuhV
SGegG1Jqmhgc2p9TbDDYgGSzY3cs7jcgDxDI6V+b4fKl4jmu8heqbOoh/MYB7olzTihOwxTQxXm5
ocm/32nddHjEMsuPKzM+MM7PbctgT310bfKUrACRpxjl6BeqIbxYaalaxtiVcAyyJGI7LP7LMX20
8C+1ScymOqlpTX89TW/eNS1TzM/HLIZhGBBF1YhZowZ/yMmYiX5XyXz6krsVfNcBCs5+1S6h6wAq
Bn2vKs5+xxP3WJxZYf8F8G1Y900gjexJQYGR1SktA/nzkz7xhGWA5bOTj2CLUEKA7N/StmTfwT5r
FZEyLUcoDcXcPJv2AVqJ6BGAk2NCj7KjJgUlscnC4ntJgJs3cVhrVjnDqLMhrT3StOBOOo0v/PIY
Pmd14Wr5PwHW+0bQw/G9qvVMtoOL3PbSJIH0hyBUcLIFdWJd/4RPRtVtBUj58/5NOySEIo23A/16
RUa0xBJqdq+nG9ugci2FH1FolBO2GEZ3cvfpPd+9zvIB3cThNYEY9UumPDDF2UobDlyggriu2KI2
+96kWvokG9th8e3HZeCkcDOeSILWSXciMHtoSN98MsJ9U2X9GGTQvq+LAJe4/97N7xBcyvH7DZ9u
FW8AH12YTxRvb222yGsnQnP+pwFOgBMu5AEROwkx3EBWHZbWMBS3M91rcb8STp0tplW5Fa2y2wIB
YPQUVmZnjaoaRtxZlKDAWhE+vpDDG/L/gjMQN7obHqn1nMqcbhYaVorCrIyIoJ53X0BCA2uQAHHP
c3P44NV0hEDWIRcNx3RUcwxZ7Y1duQLJLxGy81P+VJO0rADgi7k4W8DyiCpZMs678uMFO2QSj07D
GU4A/uvLzVXbcJeiwTH0F3XkdBzZcpcOOrUtVpjgPogCS9Csi00Bw96mOGkKIujbe0prRliI7rKh
UxALyw1VmCKdErCyyUhHvmmiwCPAq2mkklBo+i4i5kUYKOf/ofW+JlmmGu64u+9Q7MJIL2kOwEXr
91g6GreIFcKL/LXq4ftrjZKDpkmCe/uQPWGcx3fREgw0Bhff4b7Gs8jqVnUccP1LUxir9g3jT9NT
0msQFHsqxUbDC6HWHwyMlDj64nNdZeieJzEwlcCk8g6t55vtbzMqF3Rn3dx8DpIW2vqg0cikdrEX
0V7R1FW6/vgwiL0FWQx01EPMaMDRxQH6smx2lTpt1ALgWtNJlC42vK3efahvL20wwiqQiIRpLl1h
aisap8EjSAaQ0SkvwMDmSxT9Ef+O5npIvQGdQACkcso4A4iSigwzGtmQwPPve/tPRIasqLAausD+
+8jCGVgi0LMPaqYfzvVLHN/nKWKYWTvayzLj5oha+2FIO2MygtODHTk7Qsth34wb0fn6BRMYsTGt
4PCJPJv3tUNxIxw0Peh5FzaeezuWaT2Ws20s7aPVU8BHB2tVrqjIW0EGBO/9QOdPOweAVkOek0vc
PRBC9vbczo6x+tqQPmvzKRIknHNkHBDAsPRl3LGviXsmD+E0SK5bv4uISFODGDnDF6XqWZalwLZz
WuBhT+GiDWXDgVUGYvexD3uJfvOdTJ62Q1qG6X+KxLxu2jFF/wGXMZTPckzFlD8qykJAvhCArgOk
rACX5q9bxeZhN7SbG8Ddm8gPbF8PxcHb+7jp73qjXw4PenRKNxJtEADpwGJ1jafxuPIOARPrRHlC
5xblVcOiHaZC0wQi2o06eFvR0SuNlKGVg614WGMSyQDQgC/fTOoUljO8eNmdfws7O0rAmD09ZKsI
KmgBwr9ZFDIPASXXKSYnUHoLV1L4LnUgXRjHVJlAfyYNVILjYViHJvwQcdG+5rAgP4NJ5wJZDMbU
0i0lwehE5bNmCBLDbh+kV7YXEcqNHxdaT/4Zjc7nupDXze46r1fepIoddyUOp/P+prpH3ICyeYy6
vS+Sx3/RObGIU/1NQA51CybSEwBbOy00kPZMskM/cIW+qFRGaV8/3HnUT4ZSu6rMf/kkfp0Hbibs
0dDeDsn9nvSGLs80xOSl92tdaB9E++6Mnoqj/1IlRSFjvd6VayJkK1MctXEwmE/DJV+vHHpWY1T1
ixXPFQ6urA2y2FVoY0nGEBUB+rTM/Ub/hp3ihkaaXJmWRrgIfnxhnFmhVPzn59sIQ5rkeoqUGymq
uyRi7gta1lawHuF1T2wB3tdKkKv0YjGV6o6lMEOYKYO+QIqi/U72EXFFzLjl0uB/z3uFaRPjFJY/
3p83nbo0ICC+1zOflI7aYU2QNyseFsXGWNiPb26VZHuoFZcKnDC6oJu2RD6WHgujXnYMzDjp0DUL
SG4HaCTbamFfSbdSIukNvsNm2dKKwSRlDZVE3/WdpN7+1fWK2F8AkF3X7JGMmHoQGrWd7+n0mweP
muP1jHyJgVGnfjkwquYT3LjnluGwAfnnGPXjgntQ3dW8xPgdVk5fksPArzj1Do6C+zq/FV+NCzy2
q5HRqS2vya9/9vptqpa9/73s1ONv67WhgIctUouVzji+COKI3Td9Pb3K0NWrms52DdNvk8u61DWS
Owe889qUZgKauTyoSZZUBqwQ8q3iwIT7ZtkQfMHsHFFq3e7xzIS+hEXziRFiX56yA5uEntzWHemM
u9lr1vMhFSJRZDhTUifza5lX9gWrnv5LVHeY2NTGJgi0EvaHt8RvIgXSZ2mWFcjuWoMFRiysMggG
0etitJHeMcT751kQ3ePm0KmIvGGMIyOYkuQ3mR1pO6gaRszvAsClNzO1l7nb4ajQWXQO+0AWNoyT
CtMdshjyxcprLiqe2OAn1HB+93pe5nnWvk99fytcSvqpZIkLjml8L3Td7+fAQBGlonE0N2TB6cLF
4nAFiGE6bRuOmW0zN49M66evPEbgyAR+gjj7Af0SohuuapkqrKtTYNKyn7fj0VEDeCTAZ514BFR8
btETaTADaF55SFdEc/oqDxke+mCkKtdjHwQeT4qN2NOM8D0FGBxZSRHH6HPJg8UGaqoVcITrTb/+
HoZEScddkjVubhs0h8CYLXRlsj0NS3uj0xcRcKzBOv+rMmpOqWhPHaV8B8+/v7yubV0yO9hzH+sr
5k3ZrREYANftOf8EJJbjhQqWSa4YghkQPiIOi+jZk6ujvrEkMUkRUj/Fxj8xam4FcsXhKgeQvRu8
cxMfCnCpgid9s6dsIOiAotBgqzOMaVtGPM/lMVoFtL3PTspp2q1skjsXEshrmtBTZfSpIWqHxFS8
bhl7wO503GbqpxTVr10Qn+MZcXv46aY/O+I+8Bp1RgvBYirqE/hQ1a9tqKxuUlngkvr19pE7rfUE
F171LCQnrdb+4TOFVT9/LZuNgzSAZ6N11a6kDoZctun7I+t4NI71ko7jv5/qcdKwahkuD7yan+oO
53GHHI/aXw5D+hiVM4uBKrlNgaS/ky0QelOqsD4SZuxKMH7ISC9dP72VTccVNzgGW+VWHDFX38fb
6tgvFSl9+N6VPPgwrS5M0wLBj6E/DKmb3teovyqe811vaPZc3hz9Llh0keAPLA06DBY51mglVZJe
QiudANgTQo734N1kHyf3ADl+PXoBDKOm2IruHR1x2IU2rrHwhC4mX+5fX3jgJV/KtjEwYu4K3Kal
hrXrRm9vseLby1IR6EV8qI7W2Av+yNiH18ZXVU2bFN8B2PFDRDS+zyyPVfPkcVZiPYljBPvYQFYe
b2UpF9eiqL+UG7uSd3yGTSViAJOusvscTYEt0gJmO1iLvRL8Laxf1CkpfTnoG4zRquO/AIQbuWFu
4TnNTluzTNFGUYwXW56nkHAamN2qUapwrfVxVh95vDjwFrn41HCYMDAyFkISXQSr78G/6O65LVCK
6YelWklQycV3bfgLNPoJA6RtdsravIg9ipkKImfBgjx6AFdPNhNUdq+JWvzCKYXUCApYkMIXgcWm
CBpcVvpU4lRZslDCFMW2/c4S7KchXMdkx4hk8VcyvP8Q2FSV0n+99hzEKtkTiyNF1blU0aCRmndm
mEYBJYoRmtTSeA7R9DA/0Ybfv86InrF2nN5CNMYsObh1FW68AYixxsR2DTRGSgYnzeMqhq7daFAv
0oYGDT5bCvnfgVmsoGCV+fCBb9VbI/z1If4naz8BTjmq2gFlOtqpc9RpBtemwOwx5yxPhSseVGHb
S+G40hgikzyjFI8oVDkG53LkfBhzyCYm7Xmo4vpd1JwGgfzNQWg7T3gVjT5Ohih1UtncrNiiquK6
qi3vzT/bNrVRITl895GxLV09qTvCRFc8YqagTeT1EGQ5cTGIi2SA3F6OClsl3U+yWMs2UJkxJhAf
/ojIB7KfGT/sc75UwUAijgLt1E3ti8EkE9OwA6J44aUBUCuhcJmWdvyLAzbvOQaMFrJv0JNerkt8
iOos52MW0aJDaUiKt7MP8pjSylpOI3xURfSMjImXjR8mTesFpLIMs1XxayMFPJNpcQIvROFmNaVN
CTyV6bTZCvQsuLmIEO48rLlLvnLlfPK81bW8saCpH+7PKlmdoQy0G3LfQwf1m6tKOm47SQ+0KAKX
NKhZ1rumCNYxgF9aI6Y2cvUG9wJMx47zwcyv9Veahu8FfI1vjsSgEwkm80mJaJSE5Msz41H72Dgd
CreWzIy8a6fSOyYY+fB/pViE3ijiBdj6nLt5DYvy/tK23XaqXgihRBMCRCq0+81JCdN6DvV8+uHa
FUZgthA6ttlZQuEpSGkBEcY+kBcvvFjH3yhfuomQVc4DVwO9x2gorheGlsizAiTlm3huJzryv3YE
jvHwnjT/060yPjja8eLmOt82TuanBfUD+K3kTSXxW0Zm68MC6cziZXVGpsf2JrTyqNYxQVteVeJW
NpXc7Ca9nbIs2VyTriZOTJHoVGAqwaXJnMwnfgglsy0u77bcn6FQRGHh/+DFJ8ttmNz9WhEqGuvQ
X1FexC5//Mb9n/cSB8h/CcksjTH4vpuGN5aPOCxJOlTidZr4jL1oXif9uY3TLuyKRcdvGvjzhbZN
gEjSmRBYheeri4I0/k98AGe1haIAvmvnCElwpRqlPzM9CNdyEl9u4fPY6GsX824Di5UDPCXocUF1
6qpHpOUMSx6/WqJfGiAGj/SUFCjO2W02Qk0iy7fg0My5JlMkKNcWdfDvKpTIQ0+IycDql11g6lSK
gHLnNQo0QbKLuDX+nqQu+YSr7glgbVK9hgT5SNUymWiKkh0j8LnaDP6jhm3EILA8slqFwb3Lakn8
AhZfEtftxfBD/PKhmgeVfWtXBJjcak+DtvgOZRKXD2AhYxrBAdn51dqv2qduUtpprRNqcqo+dzsJ
qhY3SLzrwJn7x7h6qT0gESRdU+egKqDTq+F5MnsO5Rbvcn5I/9W9FPl55rvKOWw3SDuFqfrnYJRH
b5zonHmt3a2OwnMIb+GDsgSm6h9fLHtc7h7OfL+gXEQi0gk2KFMM+uOXZnPy5I+nCjYru0Vzr5qD
8t21KdphNKsakgnn7CaCG9+G0J7kU2XDV7FRZe00qf1yh3qBa9wMT6NL4PTZxLH+zGpwXJrOAd2g
frWA6YwPBrAPVQLtnRR4cCaekjJ4M9OGxR+nKM2FMTLzwUEyxkjKWQKvpotN6aDqBGqiwOU4PYOA
urayEU7AZvE9LCP4hesUSuAeIDe6wsdSoSLTamw4HdXuGVSBnwsVrP8PKtiWS+8TeTEET/fGSxaN
i5WNlzF9l5OvPlCa9wf4YRHDRuEnbdJPGn8jKRGNQe7GtjkZnCuOhRx7L22Pv16JhPsd2oD7SzfT
1+eB1BKr4E0fEdSsWUzXoLjW/zAwjnyzLJ3aQ2PS0UFtWKKrxibErF5pwlEGMXnJQaOgltyLI2WF
qRU3Ha+7QxHeNQG3fkZT8tp38G28AAex5amq/vtCDymN7EYWRSzHRdqMEWk/momrz12TlW5uF1qy
tcS7X0IHQ1J8QYbhQcNvN9taj+B7rw/SqusOgXii5Nb20jTeLyZZLQAcvGoJHozTwOlwW6BASs8I
RxEStihGfdxG/B9fVdedk5divejyJpHb04Wdm6ImwvflHr9tvoXhBa9qQfJqg9D4W58tVnqzu21t
ugyqtZ92hoYKq0hKdpB6fEnM+UgoJdleV5azYmz/2tRCNHLuFIlhtbJn+PjYMFDr5PNAX8aLHaBB
QHr88cxwtbHSjAOHspbHQsroXR4Nm+fuG91rFKkv5voac96AbCymY5MYtDzCuoNDxqT3J1BKqQLy
P0ZSIfE31nS+qoIGFNNhuqVIe1Z5JWPMctL9wRytdWcz44R0yCY4LuDavu/lyOL9XlODWa9d9yVu
uWgxpQ5oT+J2LmNNnChH7aSuH7JdFCgPofohLMovaqAURxSgScTaePI8yk5+k/ltUEPyaQrfDlHY
J/Q33htmoA2CVEEukzo5tGM68RqUQcvwgc8ZAfamExroXYlpBpI5IxWYoazS5M0MTNdLQXukSToI
gChChtAHjtbd9QQcJTbav1JOc/fshynKKx6wWsuRhGl8RjO8UqTTZJ7qQTLPakoTjRyJUKBjxbas
veIYJM+kO2HMGJOnmbO7HH8avT2FQTEgpWXUK3ZKGE+Hve+7uPsMigNetxvmOJo53A1erPnYDcCv
PM7Pjkpbr1+/GiSTqppC6E7WqsNdHOy8hvyxSE035myV5Pgc1Ivr3/riwwHTOkLrBA2ENPQPSqkP
mtzE+AKj3+UgB4XjqATmBEkq3z87F1TzltRE1ER+ZO5bXgnLMn2JeliULtQ5PyGFj5xzGdsNBIhS
6XXHd51dcUV0rOuOLosOylO9YIHegqU4hces3cVW8lxL/94EnaBw8wnMykWr9whB22jLiJPwIezn
nibEhMEjYVdEhel9Zuw+VUZMNLPimrfC2o+WUI6cSnotiyMbflgQ1IZV3kq1cn6mITS8JIAdZWSi
yN0fvDgZsBIt0QBlWusE0v5F33QpRGu8xJZYfQaCD2ESsrHua965O8hycL0wd1GQHCW/wEjVk5RV
T7+h2BkYHI97UI9qfSMF8IhXyPcAIB9Rud1noeySGhcerJ/P2DH7lRbtCS7ZAeDa7FLoBN1taFGm
FgNNmihS1irPpP1dlgS8/ddXtW3bDVUtwWO6yMQfi6ET+RwjSr7KRCDOD2GbshLdM8RcCQ0iNb9D
3HuAHObG3Gr7aWVkJmts/i+XgHBgzqIW5vz4zYrm1iOVV9CKt0HP5sez5IERUf9B4mMG5qMULN25
ledPBJupt2+cAKGOwjZpszQhHbMZBmq0FaOKCJr0/sAcx2pQJppmfrmMlpGtINLzReddycN0hdju
D532ijXrASHPDlRRetswZuz5aBdVvPrmDBT1i0y2zBTlQN/QXIOa8mpKrszYyxbRNHOwBZGIHHFX
C3BxEzMDgYX54UzPY+MP9yuIlvzbt7ZwkZIZ3QV5nbQaYhMAz4wMKnvsaTorI4fFGAFdaThObHru
Hn/sZn8JO7qrhBef9BjGkwmNkwfwOQcUiShofrFRlIImO4VG1sBU0nHLDTG4ghHbpruz3i/OK6/0
UrNUySzUCYoFRg0HMEeEs/xS2uDaAT7jG7uBqqcMl/3I3PPv22H50EexWgMXy4cSR0tPq20WqJv9
aZlZNxi/fVJQZI8RMaQneN1Cm5MKxiRF64Cd4B3n4OFkXdkFMxnYI3oI+BCL10pwlMnfqoDWBVN2
+HbyVeVcR2HYkrzfLcMstre/wNQ5U4pNXAVaFl3uHPO7U5DA6VAizaal3hEcoAzFsLPCUh4XSAkd
eOg2tj8GbAJnVyV8jjh3wIIfG4yGyYh2PE1DBiflD9PHGFrMi0+GPr22m3oUoEYRK2fZUzHEOSCz
vaGn6mC6Aohk1vzrH2xrhAYhT7yxIzgvYR2jOaP3LMug3oKClsseEEbY6ECYA7s5QJnyJmIMPj6u
xVm95kPnCqZt9qMpuCiUwfbgHRTUk0BhpPC7WG+pOqFpWYERVncpDrnQPjPy7y+k74lxViFaRfzl
xm55FIQGEW+aWi0q6FOEMOB7GmcRzWIFBZABryXDJfNX6Ba7bVZkEin5V7sgzsZROf3RP9b+rX5H
C13T8HFKNFd+ni33LQmWggMY4D56fY3/Zn/y50UtuyimugykhzBpoTjI/wwc3e9/6aSY5Yfu/tLe
xevWF4N8Vt0edcc/nTpGLmIQCHM2PF4YIrmJ0qiO8McOlTjgXrrVpnSULlzjygMsci0mGjMkaVmK
OzJyMKauhlQQm6wOJpJyklV2S2NQUiuzIGeg7vFuNYZibmLRwpMJzittvHq96gQaroKm//Pn5k3h
kfNZtM6InUbMCLAULwlbnJAloTYxY45Q1V0Evs8sx/Nzbe82MnDPdQBli+WuQ05Vcb1cH5psMWQg
Ovi8QZqF8QvWjTZGwBfFHkLsCkUDShHfdROlBuqUUAnge3gITN2VTJ6ktk5eX8+aCVo/BI+vqTeN
bnZ53rEdtssQapbF0JXn/tNviFw9TJfIOMQpWmODdQ1Om/YZk6rb+j3AY99n6YJM+76UhfxvkGsV
52jjHqxBxN7kFmf5TqnykVbHz49KL5avc/n44rNFd0BrDWj8Ny42ixrOi6wuUa3ZnB5/OUSXPWCF
JS20yFNDJTHheRJK5a56ntJEsnWun2NyDZnAarpEP+5p1oOB/vlxh0L3XxwUFEqafNHPFZoOUhXu
dVPlxeB5PSinArpLNfdV8IAelvI45EDrrl1J+5NEIcqbcdSuXfKnmWQtWHfOdq779uI2ebhBV5RL
8DAuO5/tkB9SDgYq1Z/h7vEZhqee7yYyKXq1+QAyaGerLrdb7XG6iqbmAG4Toez5lLAPOF3uownA
yikQTVSYH/d/pkOJajjZnRcX0b5YTNnVjSFZ/og+bviEmXE1xcj8SkP1/b8QAj2q6arzxbddu9Dt
vPlCIycWiZs9cksAPjcKlOoPqI1cCBB7fgOSM5tw6xlFUKJq+eSNwfuVElB8FY/XJSJVBpfDIfc0
C4wA/XqFMzQE9SBFQDmMszEpXoUZof5ltG+FtVJ29n2/T+12n5iQSikyKdK60VYCK0oA5V6ICzxi
JT1Wza/tgSt122VcTIe2VAla9iRjPxptTSoW+ClqAzAB8W98b5zPFC6p5u+jkBQpAhsDOq6GO3Vr
4rcZXWY5xN3+5mwQAFESwWHliLK+vvFRjCVSZzvUuW3IIXF/QYEcotA+cmLUrPozDfn8wTBkxC/a
4NuOuOTkxkVpn9YXSSRSHLyZGk/x9mAM6/qQAKgJ97Vc0B1bX7YAJexJuo6N7PqvMeNSfYQxZx0S
8zUyLOqlDkAG4TWnh7nnw3qDgfSv9zTuWIp5Cn198CiEift9+ciMLdhdA+a2dSUFwegY+r7qSrLC
pvNL2pLZjyvZQgu1/LOMmCNEDHZTFbFGKrd6GKwR+5pTPzQV//jhHLjVSTFYokVWJkkjXycIB2Q1
v9YP5dNdG5m2GO7yFneuc83rRnNUFVj1OWNEBa3XJZjF0v+KUK1jRiBQJKJRrxMWdO4oRyae4dOy
YpEshqMbdbeOA8vyos6vCrfOWGrMHbA/gPvFariTbnieApTZAcxh2ctfjw8P0WKWUynuRYm6WqTY
jgv0ELAa5cJHPZnjdShnLsyEUNxM/tY3ZqhBFX5rYXJTA8b6MnVtR8DulNhCO+UsIGo/yHR2nI7P
Qw6minuT9jfgUVC9uP36sQtyzcszWr4lwki1CdmcefAYYMODcAnW155rbbV3MieewlpVjgx5joKj
zJVCNQ56/92x2ofNNy6GMex5uKVaqR07IIk/Wh1YWPwtyf+jF7tqDtGbXGEUpDRLB+EuoU8xYFre
86B28J+GrX2fOD88bSVSgz52KDJss+BFApXmIVuhvfa82b2lqiWUGsJJb2fy1EFW/zvxgRCp1O65
+BBIqg9SadBV1kqTUHRTjCZCzo/N9Dg1/fbTG1hJz3sjdrXPWF3BZ8rDCH7Mb4prgYXdAldIiJac
mLr9I8EOVM+qpf2KkcYc1v8FbQTWUKV4oJTKGlycnIaU/E+OEhIYfQ5IsXCcHtpkpmOoFaUxqDRQ
uB1Op+aTh4O4HJil5eTGZD8y8oWpUlqSd98AZZCrw/apcHFRkNxNBoHfHpGhzPuBRzmr3wxoUR/0
ecXrV4VQGGoBbrta7V7keXc60Y3LVzn/vJK9aWt2MdKyW47ILzKPV0byPjNVWerrh/73ZBzDutZX
cMfykjrl6gUeU141NyAp2rGqJh13x1szD/S6iBJAcfyNM5l32O+TomN2aMgofAEWEPCOzOrJdMrh
dB9OjZvVa0RX5phPS/RyENki6YRKdo10Gx+p6G1Y3bFGkpoD8GUdhy6aYqX9SLxh3EYAiKATG37y
PBqnaV6lA0xSol38XJzzXus9QIZkOpjjx2v+mVHrfm6/nTw3hRxTCngA/CA2SxOQkeXT91J9GMSS
o/HnxN52Fj56YlkS9URheCzYjhTInI5Ix2ua8pbxU6XthpUFIU99TT2dsxbzhAlYE1t3oPSYQxOt
IPQ6kBSooMIUtoyHGUgz9As67HQuORUvxAPKB5IbZcb7w8ooyaxCX+V7fFqBx0c5RI7Mks62iMRF
oIvSncOlFl7soZNDSDDuzdWgBosFgii6Io1LpV8H77DXUZiI2uXzf39FlZeL5DykmF6ZCPZOF2d5
2ilixeS6YtrdL+M6YjdmdjCWIcNa/7WhVwvHfuIC4uwDlEGvNF0r/+yBinBobMqU9MalX8R1V4ib
Ob62yQspOEKSIY05bMuJZnVEdJxZsWIOmbO2Zj/4x8BuhEK6HFIivUXqXEKEV623EXx2WaK7oM87
F25QhTlbLscaxplszS1HUflYoBBoG4VdH6tOwN62hC5HW15oh+7Qf8HRaNN36ay+b/Rr7W1QvsvS
FHX/zB3EQoYzImiOFtpPXA0TY/NLdkScqCFxXDeUny383gc7jh92PTBbh/ALBNVgdfDxBjBOa5JK
wIWdKxJyBOJHt36CAFK+4jH48uPZAfDo9o/wawgYug++zClK+2gsp+N9OS999e7fLdWKwSmYEsYy
46ol7ot8x3GzEMEBhswlGzT5DinUy9csaMpLtGj7Jwk9P5VMAW5fcaYEdlZf+PRInTlE8hlvuPIT
nycJb6L6uVQ6tF2S6Yx6F43OcJ/xgXfUDVbGRx9FzSwjCYl6IfiwclKaeQBJHirp0JlGTJDVB4hw
y+GCMsmljxp4IJ1Y6MDEG3gih6CI13NjQ/8oBUHQYZg0xYqvGtsZ2ShxmVRIhtkvry/Jwp9+4OkQ
5E+bA/8gRcstloF/gSUEFQojs/bvrcgQyW4KOw6ZnlOs8XW2EZ/9FgKzdLxXj71xRXjwQGVPbbxG
LlcOdEnooIsbbubKYfyVRGE8ZCVnPPtiJ/utk1xivYIK4gI9GQSrciZ9WzHHzvj8Mi3KOpAzmv51
z8uVQ8Vk+0sZjqtTF+jMw397QopiJ0LJINxexbh9W3NsnZVIWQnTalemUWF4W2RnKLehHKpK7B7Q
BlxXI1SgyaHPHCQ+NVuOLF/+mNnjaSJcqxT9mEUqCOWUvlaLmwH/+tFK2B7b4AYxkl9CpcTfEK0K
lMWYYdp/Z0atCDaDBZtwVgz+KUk+JtToY29tdAaOjns3F+EbDzFRdENjBXngf67CPKuLRLJ1t1Yb
xrwe7hlrAgO3jjIZqTiTwbRFo2DhStbmt2XfPK9/uVa4wFA6lfLY+WP9ZFuCNZUsnzlwlMMCY87S
duBIs5gDHZ389LHr0zuu/oeMml1kK3nbkX+C5vLh/0XOFyQhphYqjjggFjYO0pXNB/kD26J2YUiM
9Hq3hbeR4IijJe/7WJFGhq5nIplanEzfETBob06Zztmc6+4uQenqBvEim7UZ9Ds2SdBdGMQlR3MZ
aG2BY7Fbq2eUJR+YaiZ2F/tGHWPNlvjmGsML8RPWXs4S2XsbkHWtugH56iJSULbQWPv+koVxFB0T
nVMkXEFuXyNcgKKtEuEAwtHg+mZRnWoQUXv6Y74OwZGxvx0HPOiaQPaE37udge5h6P0o/6hne3i7
ZQuw0BQfmQLVNCrMcK+jlGEgnpmN7svsKOGOUQ3LAI28uXPrD8RlzjOelzSJ6M/HvnbahPp3QjN0
Y1r8VL6C91+Yl8keb7McGnXjv3+dtcvxG1wM1pFYD52kuVsdMW3GP0Sf3tr58OgfcR1w0Yq1Cbyx
NBk09dDwCZgNZfaHoulJohB231zjwkPmfktrdz08Z5yotrDytjUOGX6MDDA809NhBJipYQG8eWPA
Wu1JvKRjdON8skKfZAsTPI/7Z6Xv/7QdA2+u4gSUPzhX73kWrb+jRDwT5xzNO9BHj4CbbIRQSu86
3nZiEKsgxSYjbvp1/xUjcYlz9pxptXRvUF73yMa1OzIBlBK8hlEsETm8LeiVE4pv2lntcKQ5T4d7
D4SkHlqp1sFC3J2B+NHqNX8Jj507MvxAci8GGbxAgn9s5N1C4G7kQqJtuK6mVpzSVZetLC6WRb9r
EvkW8DnMZIZr4/VB0Mwaqf91QRhaP/MSTn43iuOdaZkapF7lnFMOTaK6KlnToB43FLRnJHSIGgY/
mQKglzJgLPHQq8VugeGuDAvEME8El316TETJ6aXRYktm7cyYRpZ+BWXiWXC+NsI2G3RgaNN1Vgpx
T4JrzF09+dgEmUCmxkX/HHViQUmTk3P7NmM16NsMECMbEBd/WpvX6HoUvqT43HDar11yLdmpscQz
JhKIekDuQQaSOrSpJgJUBXNAYTLpYbvfAgTTdyA1VR9vbpFCjUbx1hLx1CsgQlO3XEJPuz84XCEw
wRlAesmc9Xi/gktcO3vAv8NNHPHL7Nl/nd1G09a4w+s5WbUpdqeY4duUDDeTQpeaQy+PV6fB2KO8
mkURcEACh4b70l/G6+a9cZrmRi/DyTfgdEHPkZNqZ6ib2W9QvZtHKT/QIue+nY2nzOLDpA+5lA1j
mZABrJmd6yEdYWV+E3S6XIbeJfvk2jxXeDuVF7qVSKzXv4nyCQTXqGVMRtlOFp5hyHi1+l6myii5
nFZOJwADTGwyuQikQKC9XeQmwLnAYj2qcMOVC5m2fdEcbNGMkJgTvQMk/vEa6n+QC3pYvroIkbcr
DXIjcF9+UxrbCHKoBJjtuJ9njHzVjtSmbetjjt2Q2zJOKhqOAJ/8exUZHNWo2uXj+Rfk5ZqXiA17
tc9A+1dQb8XDlCOrm4dUQBnQc0Er9Ij7/4IzkjV4wTyIotjgeuRqekq7XEAKFOSwHeQCafOcX8AT
mFXZZwrpZ5hlw5QwF1wC/z8N4plwuaGrWdjn2AhFxoUn+J2rFm9TDODqbhw/yzvo+N8/Qspp1WcF
9zEecONaeqbyUhIX0bGlsfMPSMDIsEPepxUB5BurkRFNwx+w8nttecfLSMP/O/1mAVG/S/PVVjj7
H0vKpujIMJ3hvcdbCKOWDfcba95u1qCGDuNuB/OkVjDmSb/zyGXIiXlHKA38myvZ7MGvOpzcRzpr
oIVRl+3PAUMN3tDtRq4Kfp4GmFnMNXCUxCRo93kE8SJwr3fI7byyLz31NCPUggkzI7saPhNGLgOf
avzCKh7U1XIDR96I0YdP8ZIdlXWYZrj/pvoaLUohPlpdGXjw3/QOhFL7+wwNxGGSME40CxmLOalr
rPrykpjP+qPzoWw1TfuNH8U/GI7S+9fZkebS396HAbrRsxJSud+KWasnQyXWJyqb4AiueaLTBgBN
dyAEt6w85McQ1vhpCqH/aS+T8+y68BaAqD4jowp0EDy6ePljGZQw96vwnkr0Dxkb/inl98t3UNWl
WsFpwca3MYZoOaCtNeHFmuWipCjqahmWiQ2lZOB6GnavkViBvfft8ydJnmIXPTILYYmrkxF+W7Z8
LQlwIy5aBQr08cs4lDr53324pPtN9ErTkxj0kCfcMOI/U7vYpOCZTUZq2NouhwekfeZWoXa+72Lx
YT778J+obxvnUryKXrCG9mWGJVJ9X7Hr5TUKfcUqRENIeg1m9PeBjacShm2EV792M7IF4k/sQoAB
kE1oSmQCTYhqb4QP4hXmVStGMoabhPt3A+QiiS3b7mgQdZ0VeuSJl/1mZBc4rbT6gpb0pZC05OTY
Ilk8Bjl0LyGcQNOnH+ze1j3sUtbMHiIwhXG9etxXosj7dY7js8nR8L2sIrOKeCmYKPZ4IsJMN30y
pXytftMug4IqM/76BG384XfZxxsebhn4FiVtBlG756Zx/FOz28CxuYgRVfkHRaHcSgrHifFKAJIr
HuTXG0Dq4K1eyVEqSn52axJn7bP5xPjEgshXIBOa2aLE/cGxfeDNc1dU1H0bXphERqT+o3IqoUdB
Xck9LVjkE3i3m1wohdH/iemTRsYl0L5bGzNGGuWL72SOOZs+TjKieMtktV6BTD90uJKyozVVTlqE
cm7y3fxrpJm93f1oo3NF1EuEsA5ZEWAmW3FqDG22w5Ke8cGg2EmiICUgmcsz0QUnMNAI3nN9DuQ6
KgDjx0UIjsV/r+oVYeKEjm8UAyRQ/FOokGsEB1FGGMWbyroXwBGwl317DqlvxsTs3K8tVtA1u/Nu
5m2gVlYSABtaSFwmHmmcFSOcDryQpOO3YF9uWMzD0zoK/pcfI5QXj3co6yXrAc9NhpAV8dcGkGr3
QHIwo/5VlDzwKKwBq/FCQFkcVOCOajU5Kg8Q+tqrh/1W6tONSSTQvZxyMubJXe2FPhoBRW/B1RJR
O75iRIr8DwY7rXUhaYxwMHW3knCNAzm0VkaQmc7btsitdk1UARrIZ56lkQSE+M1AzN6MyVpoR1/0
tiSe+mnJt/U+8DIcHHiEcM8mUvXGenRe/tHHvUANJguGnH9xU04A2ZE/niwY3mTuakWGKc9v2KXb
xGRibc0ZRoch7E1R+jbnp08LEGtrXNVl+qtWM7GFP7U3UrHmOolbc2HhWJZRFO6HmO4qDdny3H92
xOpPOhUMn6Eh81lRckKYFOP3awwagEbNi25o92jCXUWPSEg9gn77jYakARp/yO8GFxBcEgsINEyV
OwsZEK8RaPndKxhoAoqUyu4OmMp1aNXmkxSekUIYzeOAs+/DuU1+QQ9TR/HelZq+FrB4tZ4fjU//
enFhfncaquteYN88vWAIvOgbCIwlBd7RlWQCw2/FBwNEyQ9kbDHH/+rCcyhLPvXo5QPkuxUvQuQT
WeA2Rvh7XoaprnZ81kXcMnpzZH67VKA1Z3hJecCxQXLnp4YaheLnbRHMEhIcsxuE2qyQC+ljARIt
HrvIFquYBXoBOWtK8xnblTi2oJkqQDFfXkWSslfLwMEi4cUduUgkjosRhFWjLTTIXt3+bYnCq+Da
DI2a9VlRTvz40JGuJ3TbMizfY/+mDVAKN4Hos/o/mouuSamZAVB9qOc8iU7RqSs1yw/bTToEs6/3
y3LPvaXkrcP/9iLkh6p7HhhPNlnszSUk3+LkMQ2EgDnjVVxzba/y4zs1k4TGhxwr00Mq8DdUvhW/
8pbWFwV81zXeK46WoLEnOYnJFCPr5lv++q9dOD+aDaVw+ZqJTpQxB/IK3B6Cz0oj42ClsuanKJz+
zgmvX1DihtFIswerFDN7KRT0DqOLKugJ7OhymZLt1asJFPK1GcbxC0kNfd0r8h+R32bykwq5jffK
nZ/K1Ud608bOkQZLPxe8GST1/Asdd4nKrnWVOy9hmGAevV2dU2SjdH+7hn1ZMOxhjKUy1IuuQ4J7
Mhc/suJ9dXVU/UIf+aJGwb4jge6Q967i3/eok+MNUdylx39W4kuqxvQVo3KXQhJ7ZgfRkIQGr5mG
hLNMZY51WhZ8lRXZ8EB/qhGh2gYF7SAR9ghIwy6vuZKpx1fG8cKVMBzIbF2dpWp9cYOyNiEvwif2
dwRb+WvBzEUZD+jGvYyF+eABk4dOxt6ZwnSWda4CFxRVqvddSM8InT329Vt0rQH4jFT5kMmCOVKS
Ieak0yLPcaCxjTzjzizWCj85ZuiQ6gzrB43D+LhUPgeMtkaPaRtRr/y72EiOex9MhLADdkPZF99j
mBLCpzIoWcZ5+bLtd7KGz4jraRTk0FlyzCVDLIqJIegNhiBN8SA8uh+Kcy1WsgipfICQf0du6578
WKHtgzHdZ+onIFRqCTnCRSiHaCJfco0ETLJNQ+h0SzsasRhYfnh8YPJCAwyBkrZXWA01nLAY/3JO
0tN1epDY60YUh3GpGPAJDzEf3nWhNC8x/M42p3cuH/6ve+B1YdwErzKpgD9g0KmgI3u7qQgUgmww
3ohVOy6vA2+t2vokwXzsaLgqV+//bl4NgvU+Ecdf8iRe7BtSdTiU0KHPkvxq/zVdLKI7Tl1+KKKQ
fuMcEgIrjm4MdPIrgag/3dk8Swffh74ngXQtB+nDtGIYbu0TkDFJSx5siGkagGR1lmwp65vvqhlA
AcLjRn/SnSkhq7s4qVOZKAAYmmOmVhCW2AeZSeE6Qdzvx1deMcp7ci2uu+2soa/79/TbDAwxE/Ju
UvzgnOMP6srMiaGYk0gOMiiGDkpO2U7/Cg/5qx7uU5Oi6mEUXuV7o4ETkrlcKlxmcgsT2nGdkznS
fbmPpsJSTEqeS1Rt7v/Co0j2Ny73M6hOyWED+KRTLUolueMUdwyFwZDu/ANowsmjEjVjuhWLP/f/
XzRCbWt2iJ9L0efEn+m9xvcARTLstTLZ1qmPsaG2GDvDgp0DHIY84+eLTpmLxn/yI7wuafa3SHzm
evFbgHHKXyxWckHpJLtvvA5qQIYNH7hOsO/R19NFUGtgSvPuolyJ1DC0aMrXNrNAdMKtR7LF0Ofu
mkyqAIVh+lMMdY9LETklhzsa20ypjtwBHDQMY90iH74S2v2U2GVGVHXbiVGhXbCAAQ7weZH0M5as
jiYsc1y7eZtMgHTbtxwtyRijs87oV8Xjw//9BSP9XeB6LOCJLn3vOme7tmBNHrm+wxIG9OHoVJqq
HZOFEzGyGqrN3OJv/xpwBR8RVPhXCqOi36qqPdc+RGjXI1fzNwtnYbpQSFlhsVcISPFMIZzm36LQ
2BrggGV8hilSmg6SF+PTur0se88TKU26l8G+OJRMjzMbsYYZEnhtpkZM+Hq/sIdEw8+sFZzGZH3+
YXNNLH3lUG4bAua8fUloGTwb7ryAQu+ckoqM/fYaZYfj7ApY4tcYk9UW7HAmwopC8ZDWJmimGfBS
DwBnec0iSZCocnTlJC5q4l/ReEhK0yZxYPaWOegXapji1ESbV94CRSC3fkbAeZ973A0pu0UOAJFK
6IL6lDIKHOfLavZ2MOu/tl3Alh2T0UWPvtA2mTbMA8InaXFYlkgbo5XFK7Wb+6GSnLRXYsBK4rW5
KhYd8SHxfqKc6HNnWihdYHmkvHixBOEBowCnyDbUPiLWNnD4lbhUVXsTkz6emDPyhdzZUQXZqe/E
B6WP7t5qpxfAmerTQ/jrHaZXdCaTHFOyMmypEYFWIWZBjVD93O2rDEqbl54AM6lZV/hklXpBi474
UgKohQlHUkfhKLefupq/sUe4RRYJ8vn3DKz1pZV0z7Ubv0HJPN6GAcUAQJOjjHYxvm4BRRJ8vWMD
csiAmI0NXiPXRbo0ej+iGwW/UNdxNR+pFVBjUc9uhfV0mYW0SWffRWjRPOmvP+ktrCtvKWw39GCc
U+1QcKffwhtcOni+hk/KntBJWlG1zAKjrDVyro/2WrVn5l/kIMp/PoPGp63ifkRJ2p7ldwVDakOJ
dhRBmXTR+rY7vx/12pT+ZUGGa6ElqS+AzZM67u2+jV1OnyX8DXY7L80Hc+DTT5LG8Pwfz9bEjAjv
xc3LC8oZS361jhWS2cpD3Lnt7KtCSkMLliIDncOMy2syP02u5lGFZLreodBoB1XU7qWdzdvwrd37
e/CqcvcuESqnJHErYdIMElGMW+8hDjxd6cxgdPBIUa6N3Xq/Z92MGFonaJuLr7X4B6IlFIxcfXV8
o0f3VZmL7T/mQEpLd2ZMbfJld4mOvZJAHY7+GBglOGjGkanBRI4xJ/OU2MOwkfqZbGPs8qqJC+7z
ufmtNxyowx3/GJZCeW7YgweDnuAnN0yt8v7rrfBulQZlHbyKMJC9p+pIBhmvyHbC4eRDDREom59U
fwngCXxR/rst6lqLHQwZ7wVaHvj3sF8DpXoXzqJJWnRRZc/yVHXBj9qLcjkTeD1kD5o2OX1Hr8bo
jRHucGobp34GJa+595okK/eIdq/8m46eQXQZxi2s3Xz9hyRuM3T3mtRPfrRr9O+9t5PbvUaPvkyU
BJBnDGTyzNh0ZeFj9LsAmXFQzQe8XPiM7jaXhEsIEeJSO09x5gj0yoIbnm7H16KacGb3atVWRDjg
TK+w2Jt3gMCerASqHNh4ffhd8lKD3OR0Gmqs46CQ04SmwYniECfryL/+XgU6r/sXkBYM/T8iOUze
midrfW3aBrgeGq08ZkFF671KJoGQvY9026YU8xzAP1212zDGDuY1riy1KosxuYGFx9bbAWx6pqHo
XhWoKbf1JkNuIIdPN+kUlFdD1cWgRxy8E8RdB2hgWwHpf1++zSdss7iim39GerUYZVx00v8N5Amm
8xwr7hf7YwcpvL5+7K+CGsKpRo4fL1m/tM1eQy6peA/FWGVdMMYO2NP+RfTmOteKYIGx4NyYK0YH
gR7hiz/ZJkfQKMrlM2x+4TJNgFcSMEvZcfSJi7hC/lbkSu1wYLRtzaAnzPdge2t++mqkHKMQjtXH
1BMNhG3/ByHMRvhG3RNQZMje0teMXcadbjqYycAkUEi+wfe8EHrEpMGg41/DVMSdDdEbH3BaPOHm
Ob2TqQDWzFuKZkslGUD4nWY7KGq5lw5uOmWxQzIArBcXznvZw/tQ899v2v0mNGGVKGGe6azs8FE2
antCtod2P+1uvdkFNR2uT/332DwWPyyI8s+gpPb+G3PxgaSC9MtaVK94v1xsT632q4D7J5sEkaN9
44dgWypCRlSAvqhCBbqbN10iRLhFGmCExUffZ94mgTFPgJYI1dvy1sB6zwl7BEGafupCYhfZnKcG
XC0kY17SSC9a4R41pGBANws3t8KKTFeK9U+Mrr26Smb8857fwbXz9RxYbREL1nB7WMEljmy/Sd0q
nTK/U8u3FNhjmHA9mSXKWW/Vl22/CZpI17EyznXLu0jCQ+mkL7iNtW7rGxzQqF9zTp9+lbygL6QF
9hDeJ2AuKbo0+E2KizijtF7U+QhpachKqkKE4/JMUhy74c8kO7GiVTEGqZSDrSO8dBGSoXGcD2qN
fJJC8n1cLNhCIryWrAY4p6meNBFhpuezWGje6cd61H6ZpxHjMBNEasM2PLMCObtiNo5fbhCLnhA6
gRP3I8SO7rlncdQwOc+vXxE9rflQ9Xd61IQeKGiyxIL92gfLeka29Xtt8ap7syoMJCZKYhXq63Qz
DUrybJCjczxWJCYgfaWTUW2RAXTRuaS6yU6PoPZHxa2qhIyoyQyt1gkyRwns2JwnjbfIsLFwpMZJ
1Wz3vhjlZlCQQmlfxhtquyo4WB5ck5ikrbglMELPB2C9t4HoYjNVuih4mujhvw8zNVdWH8Mm+MAi
oFHh32PeToXi9IRrzF2fuYY/RUy9yGVYzSwwKA3r4vrqIRPC+WeDpdOftiER3m/jiXQEkLI3u45s
pP4IFnrFrDg+aRHDtO00s9Ins7DwKkF+cuPvv56Pi8nAoMwoeoQ5s3Hd9o/YTl/JOOMK5wQ+5ck1
eu5xIT5CHAOX+S933yR4BmL1HTQSn9OkG5m8gp+l74jH+Uf3IjAU6RKU/i/y/86UurMWViTmWdCy
gTuhLUbFbidi0IXeniMe+YYKnRZi/Td2d5cfKaI0llllaROpXZamAfYUXFWgQ84giTLHfyyz8yvk
9MUFa1WAtI7tFy/JdQKZSpTa9+gfDykzfiLY/TMC7VVbvx0PmCuE0Hdkx8T742daC3B/EUBAz4av
Qt0nxIhD2XrYFfT9Z0vSLAptSRPtTKcMU2e08/ExD/R5F1tb2P3e0l4tFGSk+Dd2nsONG8lFTNHT
VF0+kaj5/K1S5F3wXs/rN4hVKbmYiA8udbRS2rXP5B0BQVKW2kMek3yTLLIyEyTFxKj57KDy+q7W
pl7PLt7RW4b7qNQKku14HAINlktKB9jDGMzTKg4TXGT0SsNIed6541x7SVvn4DVgRaqBIZu7BwrS
xeg4C/6BEtY3RHdbMXjNL/LoKb+xzxkoZMqjPTOrwsNA8clsRSDRv3SwfUq8JOASt9/G6vDoIW76
kEVriPnmaYWR8KbohrDv+f2qjxdkr71zSBO6FHnvACDe4dnWoGaSpYhh537UbtTx4+mMgr+DjK1/
SJ66KbSIRPRiAplLjSmoHo4guvXB46ziILUo9iQSy9s95llDOKTLwITvN4aZZGTUcOIDdWRybOFt
sIHQBCUYwPtIkKQGl9gjKiXQZk+DGJg8jp0OSJllKIUxa6nBc6wBIB9+jXlqDZBY7+/QmaBGOHIh
msCrvM3AC6H/sqPiiNNN4q1iMsc5sIZjPfylioCCQ6FTNOEuuJ6Ni7ahv36bV7+nNLWmS3vq3CVd
TOORhoVA3zS0X4APUMO/pCr3+MXfJSBEacnGEtncZnQZ0n43Tqcn5cEaIZMjCWe8MF1c8KeGzCyF
axv/KVj1KKimLjm0xvvf7uj+HTNrtC4a6uxeM0kOkBe/fyonjqMyWTzD32XXVpAlU1SOsexf7lro
ZU0/BGU8igpkUcom5q5+bdNbGZaYsGIaZBFnxS3zQeDE96LuzOVa1M6NE4bSbdRAaKNNstG+uJ87
1LoqKe4D2SjrYO8euOl81f6t++WEO+oDnHkLLvoXrGH0iJvHuVviuCKhL3L5IB4A8d3+vUucRr+7
HZZJLUBqUqITcpQ+iPqCmTncNYprggG6alCMUT76KM4UEggjBWh9ItUBHo0oU3I/gmRuZ9IH8/If
VLzK/0HSbM1h1t6MKxtnxAz1K9Uzsq17mkjN+bSqvP1bmvgtqfViyRnf6xBNqkNw5wIngJ0O7lSd
VtZizN6R5D3dgCZ4ttIVDuDBy6nl6j9mz8iyjjPJqWxMh7Ztl0XzmtRVXgTGRvWDQ7tD4gThx1Ts
o57HWULDwUJF6vvZ9fKGzYBTsZc9WgV3PxozI/O3gu49CKF0hUUiRLqSOThJhxyXBBpyt3GF5PSK
1beE4b2WaydfmWMPoKueKcoAi8D1eSHyTp3UQS9bOIi/huIome4CwgAdvElY7wMcLXs6vQY2yeR6
ug+YhZMC5IUvx+8eQb7m+yGdCyGpdxniAxfISYLIq221gOmUnol4n9FTUK1x6XToN4SDTWlmPVaP
HgXVKAdMF8Jq0zuWmSC4tjGtquNLYzeIc0e+FUZbruYjGgTaxkkAXnkdiEMb7xBHqLzY9Gbk1AIS
V8++baVIUs0s6QSZpRNO/X5QdLW1Tf9vGwc33ZYL3bz4Pir6wCJdFww+ySG5xBJ86mbVJZERqL+p
c3E3XkmBwFgViDy3h+vRAeAdzaGyBHkF39JUpv5dDxpPSR+ixCIy3uY1w/124zLl5nLksLAWcVPR
/kLI0JSa1pGKVKIju0ao8BXz6pmlMbno2kPFqqtlPG+Gnni9bFhGCrcDxO4+Pg2TIxtEZKF4MRAN
6KSuJqV6OExkph+p7XVFxPeW6y+u3XNfybtQ7lVNzRfxPMkx9zy9JgjGR00TaveyyUQY1MHF8BUy
548BhKxoSkTDh+zEsLTHm+yUXuuv3A8GUXAa2/J1mrH4MNtQypMwZlUCdh/Txz1df0+Iq5QRoAo0
IQte+KP7+YPDGZfpbaH/AoXOEYtbqTrlioV3tm1tlyotQS3CBwGF6AN4K3NL/WBtmO466uakZs17
3PHTB2yBzAweltys7z0LS8MPRt7cF/1UsI9q7acVVXavwxDJzvu9KDq0ntDGjg2AoJstPUu1msds
IwxEbyQkWXjdh1JiJlxMRrpKHi4950nNdfZCeaLwiYCwsBHQ+hmdcXCtxDw4Z03n0RIVF+rceX7Y
JaLy2fFCr0p/b2Y1OfM7GeRmt89XbDKr5WIhMzjYZwnLvpeTAcSaORvsAZC9amq24zy3FqBqJ3Ij
xkCxIsiCxX/sIXCPQvNGRp+pLAloC/z31de6Q6VOwKSFUl3WViFbeLIjpTm7jGHNi+272RVOyEgv
NPmVbuvcITY561qu0IOj4CZGii2sqkcMSd8BsVHsQbLSneO5UgR+Ka9EkHLoG3Ek47hKRcy1soaB
9q+N12rDEvHAjg0gNXdPamQ1QW4/Hz3L4BEdeBdb0DoAJ8yYLH8pp+tZ8xurqr8MqDEIPZ0F4gnZ
0UHeTy1e91XFdhrWqyaZJDOlquTzQGFfXzZwoHd7SXGPU3/dgKztq0M1YLhFk1u0uoWk2E0mP1F+
8rUgqRFMGWdkGbiaH1tayj6ROxGl547mMD/XQkctgYoSUSplx08qvxshZSdcjB5GrLRIid+YpEb+
fW6rt2CxL1nfpjvmCXytWPYJQ3yAir8NlhrGyqmBcSp4iFbf1/2ccdgyHUwCKckhFqVGH9REMzos
oPbkNk82N0uxu2CuQdXu+BOrT0hE9YQNAI9n6Y4h1w55TqOfZ/3kAlglGvtLzQ6WgL86sWTkDEuc
nOu3jtxiJ1z5JxVItscgM+94Qb0Fcfba0VnFy6pNGeRF9gDSAWiLQKQ/gXlZOq0wTtQp5z+kyXNW
TfYV8md7GWxn1pTjX3KZauI60xZyFG5ulwzo6g25PdO3PaXSF0F4LtKvAj0t5w+mGTWW1U1iCOga
cSWQHHsGcsgw7a6DyEfOG1vrf3RcKy5KOEs0oMaCi+GVECq9VeHXzUznaHYh5zwE4Wa81+JbfYgc
IeWA5ZBKzhXPmH2djVTiMvBOKiwC+3VP9dGin4b86EtTDvJW/N5I4m7KVnj+66Z6WV7cSIiKbLSv
y7PrwJveeHj3yofmgSVOjNzeeKlo6md8VFR/5fxTK1L2o6+/L1GmdIUucFnb+SLx+Y8o44yADkB3
Ec9WQgdWusAFl8wwr6Uu+iuZLnmSWhoOqUrwCwSm7sICOKNblblcI3sJbNNDzEG7hEoXZhag5C4v
t6kLPz6HpmK8sXjHik1NSqBsqJ7gRRmB7euLbLMuhR9cpzfjMBeMY0+7JyXw8S8sZsVDqG6+fdnO
T2VyrBe1iDk0pUMb3iUDjBWUxTyVLpE3eIGTvGRzwIuypeQw+d3BQXJOC66vIGO22fdV8VVm73qZ
kZGftHL1lUmvXDl0m1AWGicsO8qatay4+FQWVpfuo2IMo0WGSMVYHHJjtTqY1VL40/eTfEGyKOlv
pHaYXc1+A3K/koXOyF6AokYsNYCCO2SWiS9RrMDYLSOXDaTtD+tms+LDBCP3NPt0XwvDpa3eAs8G
is51KWyOxHuj36q2Lam+UA5Gd+07JtQkrTqiGI1NBaUk5e+cZm+kF3RoCCYJVb8LyYWHjaZIvXEV
miQxbFKt7wLSwP/bK9iKC+KtBL5wdYErWpRyGr8ES53/w4aXZSuGfSUb0A+KS4aTv3/l5iRNx6lO
rZeWwlYVXIapxR+ce/jf82qOGgkdH5UTxpT0Y/p1RtRy8TrCiY6apauNICrvcdLCRS/fBk1hzF3F
Aj6Hbo8ja/rgbApmOPyu6EoVaPGCIEjwbs6l7dZLlHq8bbOXC7pPcKKroCiUCcXT52OYmXNHnQFT
7JGokHZymsDHxQ08s9uJaSslsfVuvqwSJPz6JsZH7byx+NzGF8S6pKgZlEs7U8a7Zh91RVZwuDds
dL6D57lGh2PqIIBbVILTDleuTPiiC63TZe0EWXFzU4fX0TD9wlOW5FCG7XIxjwRBpO53b01ZcPA0
g2s55eBJDQ/LkToAPV4VwsKL61LoqTsdKeQJpv8Naq2MypET8LfTadPpXu6zrpeTjXd6IvY8CPUK
G5poqNMku5qcutnZJ96Gi6AKdinb6uljbU4bBmZOzlQAC9jVmD2YLOOgZebJ15uXUX8dtKIUc/Cs
GDkz+uhUdlkHDCd5bGmHAg1fnmBfXt2gknjzjyH41JHUeHwdeUQhhN4zg9yD3NfBpkatNoVA40lK
2o3OxHeyftzUsctqL9omVzev7++N1yuAvlFJ5LdpQgYM1rFb+jbMUvMOF55h40yxu9MeObP+OczJ
3ss337pi86FRZoSQr3Iz9ZyzDbrjJwVSqrQlNjIsbUioiCHr10zmv7ZsbqKq7TvxGbGLv7VVXvMf
zEqlY47W/LRMJgneyNt9ZSL5/YqYaqVsyjXVjAjlesuQtS54uqslX/F3/F9igS06bxwqPnqIdDkm
hikkJ4sKG/B0EBaQXEdCw3q85utwOs/afG/dPCzkqIa+n40o6RoUaBMgcFkwn9NkNait1/u4nNt9
M1ySulJSiP6tFqenIlCJvWqFDFDQGG0tc1NoQfgSTYZirSsjeyzTb4XAJ9r/h1EF1LccccloNPeK
3I1nbYNyfTjf5wELokEwYi6O8htKnFSszkGznsTvsKNnIWpn4S1HCgBCK/9U91BUyHSPVOHGx+K0
TA10IATrUMqJ4Uw5U7O4L3zGCxpRzfzKwvuc6DpqaItbkg+TvOy5WBzFicBqjyIArcaZTGtgPWpS
K1Lhtv5+QMRgRS56H5dcOdERqeD2zFjnyX2ppZAT3hMLT8GBEoYXZ8VXXm/TQEEQEoGyWx63JGTD
Se2ijOtYSOrDKVDoDLosI/Jxb7l5p0Zks/qXO0sqAmzH6tK4Eo/vElYOC97daT1hDZGBbW7Q9hFj
7p6TtLU4wEGQ64FPbdGvewSlFsEr9jFdVJEHB/LQ/ubv2yub7JyBFjRmo0SsbVx4g1MjBIcEiom2
BfIwdp8eWpZVN6kEts+06dz2mv02/QDUQa/DpDrvqdYQKXka1Zj+5J+rNVTJxrTVASMv4bzlr5vj
OLv6uP/xRizQP1iesiyzxGV7wy2xo2hFmZcwL7lGmNIDE0dG+24AiwDkwDTnGyO33pkRRCNj8RfE
awHK0xdnZWICNq+hTQC5S3PdQ7xRCU9tFOAKxfF1NrdxtpwHl4IX7kbALMR/s5nKLw6Z1zp+3uMS
9r4jwU+k4sJT/yIKinI075pOdMD+U9X4u48I370AKP/XCkxRkCRtPbwkEck8/u8WnYOhR79ZukQx
RrQhre7zZC+mzjIjibnsrGL/Ru/CAuPSSatWn2yWeSj6MD1RF3rfEAsyermp13x2oOGcLJeKIG7e
vkRu0JkRRsdxikUpk8Mstux4fhdtTYYt6G7CeFhVyFgYm8fOBgnIDn81s9JmDxfd1EPgnv/YjL5+
fRJZ9e+yjhKQsZR1SgX+R84GKYrYSPJn5q1vdp0R8sluWjsPjXnizZJK4ZZMmdDRZux15fhwqyej
b5uP056YKwDj//JQMDDSNJ+msGJwriAAeuS0pFHda4a56AnYFgzr0ubwmuA6I1YdJOkxjUd6DKi4
gLO7/yYc0KfsCSC8J6mi6vxcDt9PBYIE4JjKhWB00SpTCknFmOhhHGRDcTWBiDGz8eANL4lP98zt
1AEiastGWoyxJNWfv3sWlwUaiFzBSeMRaQ6xdoRzYYNCcXKsLObiHBezLw5AUx6f+13hkyrOGbKz
Bal9UNvtVMN9jRzvKPw+ITZ8rvmMEyLIzn4hBDR4JWDmmYnwKuaseYQlDK+iujYbt/65afwm0N/H
y7Mm8kb15aB+jsKPEFrPmFx4kR7zC+yqs0hZ4/znHGGtOEIZivYmxYRhQHJ3Kl9/PfiBEraGCiRP
1uWOV61S62XQfrEuU3tBtss6LjlStGgGO1nGEyg9iBjkIsA7Iix2UM1Vn5KK4SMs18cuU9NsLrqz
3tgcedgDczi9tyN4gg8+Enw+G2QNpBOtqYnZn49GjD1caJPqlmrVLJNWyWWauYOvmg8eS8o8FtPS
kQggZyzJgXmt/S6rsR0M4AkxlKx4SlIKDCDry6MCi4V3SsZPUZzJcpag7YKuz50q48+D0hWTgwIO
MQ/8nsNJBN4KVtw8t1ZY5O9Fp41TOeBl+kxvdP2BUbf+CdB8xrfAfuEkXT7POU34HLNxC6ZtV2m2
q9PNQHNIUJTncsrgd1ScQmTtgBmHnYkclaY8BIrupQ/J6lDgVXBpxk4R2ziHmIDouuN8T50z63E6
1TC17RqqzNPfDfv84T6qPrSumaLX6KdDtEzCbnDJQ0l6fAV2Nn5y0FzJdjfuXomr5pSPCLNdSOGP
MtLMwFh0qUAgRjO2/p0zoQ6VJp5WbkL0sWwU8pryvok8NBWjqHrNAeA0oyZ3hBFPvI59YkpqA0ny
B9aJQ/GLjLZ+gHs1n3GWQhg66bjdquW6swYy2ivLjbGFe60zJVvH0FMF8ih58ZOAsfjjRl5djlKj
90lB6pQ4bTDRoGGIz26iSUCKO2zFmWHGVPNGduQ3oqI0QoAxtIjjq8Kya5Rra5CH8InucTG47KPz
Fbr7KZ0Es3zAlLFyH1pJVPSVBWcImr88v0ZJPGOmpe2Kviq13Ep1lj/3ezeOqwRyn+88RWALMtxq
/06oSC7T4C+NrwlMBAOCC/H5MjOQ5Dk9v8ngQLv+S+XYu5zlNyEVc05KjYwyDNIWlrfzsFcsdrsB
GM/S7oL+x4hHsQd6ZLMJBntvbzK9n/tcTyeISUMxAZKGUxafKp1Ev6tQLY7TX3DoLypMu0aoNZ1a
VNfyUo2ziABFShJsCBc2IAEpXqXj3CLtTEkiajchmlnPRavI9H3G6eSdSnFox5aEDzuOeoQR9m59
HQzgiFYBPgXQ2oz/UJsZkdXHKeDGs/KZHW5Ev53I9s4C/A0t8HSUFXmbH7T0yjz3QUPyAK8vXWFp
+1Lv4wg4CQOtTJAxKmsN7h+8YEelAsiMGmWsVF0/AMAwMicxiF+JabbbZIprA3b6kRG0fDD0S/Bb
ej/639nMnpc+b/0+OOWEBWzHxY/Chi3KN7VuNDl0VJY2Ni8hl1g6j9C+YS01SvjBDfVKCV9AJEJZ
ZguaAzQCDae90D8nRV6+sojv3E8teoRBfhFfkP5mowBs0e+F/1yCGVBh/+rtFBEDrkE6rX2Tqt1M
8u2OppYpbijQEkAsqqNafXJrcNnUT9WwcEOZp/ZjY5I85hsEJSXwEvdg0CB66rP9Kz4JrJw7J9yE
cuIILzZik5Cwa1tYaJ/PZFDDTJukMqN6sq4ktipRYXWVzpceADiODnqkEm4POLEBYAo7//GBVIit
acWHrv49uJFeQng4mYjw06ERXF118CIRZyQyDpLO+ALmjPkm2XY0Ho6j4S6t87lKBA2okH99M1t6
SPyuxLpjVaX/RIC4cPhL9C/ywvwupm/q+1xT21CKuswujTXVEYDL1R6hfb0ZLqAuzG54LlNVimGH
1KXp2pOEVpkpeHMCjL7k+2J38wZqSckeHVV834JjGQpye95NPzCFUgeCaTu6O+10ZqYhw8RleapU
Jj9RbWq/SgCEH+rZYFvuZCcjospk9/P0bqnssxVY6n/gkqPRn2ow+q/M355dfqeZgSuE70KQ/MmD
m8qzOOV9Tb5FJ9yqks2adEh100GhxAJc/IV8j5rXIjq8lcwmzpWuHSCZuUG22UToUrGewcio3epe
32PS/TkP0qfDyrnzLIbs23PTTmfJzXD92RMN17JQqUaueu5x/0Yr+Mnl6Mc8TYibPIrIM8M8Omnt
z8q8ZhDxdqxrZfqSiCE55XRmdqmYsj0NP9z2TNb0IdZ441iUi65MOFLcxGXBXmONVnwTaACn/DEj
Rfq+dFIGn4nhIgXwUqBK7StamdgH+j25yraLvxGjvdc6xmsxFTYYSftDHM7OT74KmLIwpBdHKaaX
IjGEzrxSNnLTbSmgtCuNETDHxhbrh56qKwsaHQFFxxMsZIJaHywUU7/4ohG4EEdyBtKxOaTQnH32
EB4wmCKYASv3KQ7rVl7yx8Wrh7yrjsx4YOKZOrqgFiCssZSDVXe4NGyNgQSoNAmXDlbkNfGHZRCR
kGeYOlI2OycuIHrZAuzqda9dmbRadh8Ujm9hkpBJLqzwgxaQNoqIRXgYHqHsl4kEcmiMJ55opKJG
/tUpN8RZOKx7hvC8cnKlSr5ZzxfomU2fmLRaCG7HewME9E2hHH+NvjtF+xutRtfOY4cEwcvqqZXF
KoC09dgETXElFOyMJnzWDYj5pFMMBKPO5FQuV3SbiVtL+prpS3Ah9m5U+/ORt8VEiR9xdEQdbhQk
jdPJwbc1buX+8kcqimC3xNBXCeVM90TH46JyEgysfnXbMTMyJ2a7DeP1fhaGWRJbal7zjcrnMAN6
xm5VpPbiPe72u269flgBSVPRAPmtNcB2tzbFUM6Sb5ME+FZPKMqg2WFXhdsp26cxRsPB7AqAAOq5
jFn5/H2JFc3hL7X+ZhQeK0/c9UgZ4L57BmyvmbxVHEHr+mAN32sEf1T91HZScrjqhO4a9qFNXzws
egJRmBUTCmotoOFWXI34FWK6ZIEK4NRlZitOWWnZKH+xyExfr0bjDR0xsmAzmEfKpqz+rZKWzeYn
D+6piMEMXrROEbvYGmBRxSXKYwGZZ3XpmYiVyBH4hud2xNZTx+Ao4iSh9lxPcaF/HZB63n7La9Hk
kY9ZzqHRv3IovSC2zdBeFrFFKkhMVt1Mg9d3nQvnlrMTM27lJpyLU5vU7FME9Jl3GUj54uZU70hO
+OA58eH+8eIUovTjNsRsypEYH8SfyR+wun5sVIngWr7PxCd+NfQ6HOIdRabS3ZmegUZxQBAuVGyk
LND2WlkD6Qo9gXZPmRGcMvprYkm6xXHwnrX1xCmTu7oLurgUIu4zE4uNbXg5WVNU88cUElUWJLmt
+tYMrD8zndzCk/n8wBB4rqvYfX2mKYyN7rq6WMPLGJcjgkLRrurmHf96Ig/DSGg5XwIWBrNoAL9n
wtrks/3ray6++DFI48xB9vOG55Dzo2LZOGuigUYN9SVj9CGwVjZDxAnjDI9hGdX8NyP8i8ak/nM4
E5A8DM3PXDVpE9M90BdkG1bidqWZ21m4KNR16ApoCMLdlBR1YvPGyzMtqGtvjtNkYKCXtbdTI9uM
+SDlY9eEuO8WHMjGrMm54GmtbhsVjYvZS01cZJlXSjTEBqqihXAxttNavQe51HVj0jvxfMZFPUqx
jY09af7xhvQwFCLPxil/QCfUL6ZYZpk8XzNXdMAI3HTM3xmYZ+8INq1HjKe+rwPJvHaWbQeOd5//
vAi2pIfKDxWr0ztcOMJAxkIHKU7xENP4HvsB+utdjxIgBJmuS8Ooy00BxWdIvB1N0OcV18MqCA0h
R6EYfZMHQ+4q9zktPXwi9asyG8ALvs7HRLSkRz6bQ8Ml2+8a8jwkaY9qaxZ8y2EeuFtxjkxAEt1o
niyU+9VZ8oHFboFrhjUkK0xDLBglAaOcwoH1HowUlmQeKtU4qXcTGXb7/dL9Un+EreDtbsXStDR7
/L7Iydg1OimAg0bPdRcUHs5kgQpD490sy6Wjs91KFaiAc+LW/WWAZ9kVs0Y96qmHhNuxEWKlKhHQ
2oZVqihUf43KG5KhJyw3vejbPTmd9awpx8fBkpAalot+DFFF98Nr/V5f1W8pxjj6GdkoP37dvba8
QyGT5Ciie/IzwLXpUCSLcadeSOqYXKdGeqEq3QSadOinJ1bPVlnXdKgTVII7yY5MbBUXQfCrbYfQ
rvRPRBxLQ+hkIRIvkam6OgzhO6hrLx2mGW6MZiqbq4n65CMFo644bpDZ179vpHO0ydlzthmA6DXF
5Glz8mE4hSIA0lzO+eDqd6FAkvcCi5I8eKEtTb3YD6XV98kxTqX+gnbnio4Fsh1m3pi2K9heyc+Q
alCIFm2scBOZZBlgdPTNP6q8RKQeEPCNhPyk+0fzKCUaz9dN7jDDWrzS4XUdeXP/SXSbhbaKE7/y
pTjVXvZ9X5fbt30gykbTP6D6vntw+C6JbpFQ38ggPvQx1cNd1NKDbC0q9A92zkk0i54E4gB/T5ZO
IaPICOyf09kfwkq9DW0CZttjJ7l4rrT0Yk4NgnosXrU6as3AIvkYXGcSN6ecGX/llh5HC6gP6oEW
ysqqrkF1uu70ku5DLp4RrUZQjuF6GCDPpvYP8MmekSF6Az2kelyZJSHVgYQzf23ahkeo8WsVebKr
cGfoKalAbFRtzVjPRSus8cNvqZBIXH28DMkmiuBAKxy1FtsUaLA3ei/aG1qMobPv3Wqq3rFa+toG
uSoTclYq9JMyeAq4qU2vGpxx/q2RLbWbcEGkGXzyi/EEt8rkSTU9Lb3wzzAZnTfBCp+15bKGxhFC
J3mnUbHaTdVP3NsFQIOUDEjYGB+0foSODCa/7RyttKpWw4tEjiwnEaO7ZggN9tBJk8+ZUXsLM9Ga
+PfoaoDjQZY/s+ISNn1ozrTHrnuZwiQCx+gEZ66zN5zNycuDWwMheSVpuylCBXTjf5xlbHKAbcBw
CPbblths3cLeiVyFhXCnBmCQgpqXSqNmyiCHWuFTN/hLyaQ6LTWnL0p7RRrYJJNywc4KFymbT5b4
jQ3ffrX9tkRDXgIm284qfb4LvTG5CyO2LAsXZ4h9ps3NyKQDXTS0SDrJzjQk5osVk5ttRwE0+/Xx
zG+71kNlfv7dsXTuBfIMolhjbjT6vy1RoQysEp+0Zdx8U52mVFXPrSintyUS9ShEUPEaAp8fxoxR
qnDxt4Qk+uPehsZStTlgGZJFc+1h4qTmtNyk2ctzBYTVFaUnQfb1RmHPwpq5C4ldQuZflLxapPEO
p3XkN1oTkylXm7uZo0OiBaJst4hU/aoIHdLdQlFa3Wmsr42UNaoEuHzfio2fHE277vSuQ4DY/Idu
B0dZA2AtRI2lMeRRu58yctZqDUL2walE3j2lM/ysuhAyKbCNPn1VTp1erbaGDpzMyAeKAjxhW5vY
4OL70Zr6EiLFdE2RrDiSE1DJeeIJbmUsWpj6wtpg+XU401JeRZ1ENfz3WTERyVIx8ccVSangJDwJ
XbOsZw6SjDNBGsHvMdwqzIENQG7t9yOXXnlIZVNzBX/qh7/wcozTUqRxNz8IW7SShr1UIm56eXax
KuFp2AuPBmINxESBSYZxwCkfZTdxQGuEx6ITcgrRohJ/IGCSv8S/Kphp2Xu5ae6DGNJ4aDJl8lRc
8+Jjyg8pTXpRyIziZS2hyDsn6Yrl7T0d4yoBHeNfxW6As4pHNS4h/RLDC076Zn3aB/nvxdbzRWKe
KHkPz5XOsRS88ZZISMfr2zV4UzaHO0HCW72/OCh/ZeHyYuxPBlanr2wEBl9B6+lseKq9VD6nmKxM
zZDA3EEI7BHO2WL2WnLKeO9Tg4i7qoe/AaDrecbImQzZ/ckuF+llumA2rZDFGFYtPr/6U2XmzTCM
uT92KCYVLmBuN8EJL78GTspzoWMDE4A5SYiqtx/dDgGfi+o36RamUv7WRvXHbLfWrlnSy8RI0uyB
WX7oQpXgbreF6WFhOihHHHbX7LKKrwRkCdRdltFZlkaFhsi+GwfPkVgEDD4Af2pS5i5d7Q//vt7T
EnqZ/7hGZZjiKbda6ATjHnMPLObgUBp+TmeIFuu9injGGM/8hU3CztHBaDs2OmA3FIMr2q/rfYbg
HIk2xKlyE6WID4jRpqBuD5QVwMRw6kq2PX0tBcANiaVUC0dAtHcmbHOiSQOOdi7zseyL2kPu1Uwc
XBeHSS5Rfc0EYlRGxFyxz/GK3aALSzjK56pBL2H5abIl+WbHgJF6ONaUhskpJQ6iQgRL/a22minj
23jBN4ObIuBf36oOnpCuHCsuxhjlxW3BJeGnX89/R2/AEgt5k9RLbSbAXXySt/UXTU8jJSCQNBoQ
oxfdjpiHz8rZ7p9KObVsVDN0vjF6Lf53BX6grMuqV/UGXn6vz+J/Cx1MyiyfrqMKyJfcCpD4x7e3
wabhXwSJGGrSfr3pbU7RXPqY9hUzsjTQbeyh81TDoJdjfiPqCr30VChys6YtKmlLsjnMCGETceuh
zx+a+mVAVwRaRoNb0M7WbsY2ruHzzrPP2mALhD8P3kXvuVbXg5DVXO2ePFa5TyM8A2rpB55H87TV
VaQsrLj2e6afbwYysh13P6SbuX4P/3Rcz3zFHrhn+LWM6ngG/aEk4oN0tFBlOD23JlY8SkDdzdEI
14orEWcuvfteZ+zvIR05FD+Hx8GORM88ox/J+vrTTCcdYip1U+kWl9gfA2JV5VzJhbLpmN0Wp92R
pN8zTSe67AuRLfFy81XqHhBMQXuoU/ulnm7b/wskFrIrUYeFn+GhgZ2x5Eglwg3DuIJp4RPjXaLK
v4IEeEcYFf1hpHnpW7H435URlWwNpweqHyh7IHXo9dhPx/NMflsAOdq4aEPbvFbdm1DQAzasAGX3
P6tNwVh63zefe90yFQKB2cLLiAMgO8Tpfv+lx4UbmBOJXPYCVifH+4yH797jgyKiPCfhRzr1jFtC
VTwo+/Cej+XMtWlpq63pIF3ozJMwwHuX3qTq6tpnwGM/fDT3oUun1izOLtn4l0WA3qdEkWHk0+ym
lO/AJxz9HnsgGlGiBnItazFbEXcfyECNgscd3Nv/Ls3HBw07AASucQS5xG8KrJ7DD+eHs4VvZW2X
PqittAvDumCMbIPmO+GOXjtyVgsejhtklGxvOG9Ou06VkLOSSWwV4WMcXryWp3roelrrFzNK827y
z8un3CYEUE4ysZSoZoCTyWhDT3aKHpYWIRbbAupiFviH23k8eMtLMjgQnC+JtxH4wR1bJUDGsRON
8z1TRv4Cdka35nbFjNjtPaCihM6n0VGBjz2waLBpo7qz+qmCDqt8RzJJlewrf5ZJm9TA/5M2npOQ
b40uDnoLeMsRlIz0qC+3tjoBEve2EEEQv3p89buzM8xdea4Xvl7S3FiIfUynuhRPrkXcPllexZhe
BDTTc/ned1hpLJWvBJoWljyLEqvYOjmdepx327KFGSGYd+/10W15aVMdV5YnPfzgSbIIpGxsWvy3
bXq0Pk2IlSbRyBObxf4QPL7HvaubPzHr62gIHNH0RjlpbMGHF1289EGh0ug4ENyu7r3Mg+WN7chi
0U1PJN0toa/V+guVp8Cq1X6mT4njdzdMNSW52P/LDS7vsZoKYoal2XwLBHt2nCObC9eEG76BthNP
8Ageb5lqt16HlaOTlGGC/MAAnrt6Odcr6CIg5HBP2Xy9omaEJu1l6Q1tJRniiAWjx3N55+i71NMX
Fw1mkFCbzzR2g+wO4KEIAF5lNqIjKSVvxN6omSv1bvBPiWGdA0ajCqxcjYcLChIFr8Ikl40NS7Sd
nCe6tMbPc6tZF9wqemU0eQgtlhWj/FGpCC0rMTVS2F64KKwipW3RYeZfmRhGlTnoG3U8L7lwa3d8
0rIwNyafCkV4YoCfU48i8lx5GjD6HzBbOt/v2f57HMcJsfDMox8csJ3qyIhQDu6180s/K40wp9q9
w6GLhPshSMT14i3n2zHM+eUdxphKmsuac7bhqVbuPrw5SRYUo23Dv8QifJXMiaMBnsHDGDznsIoG
2m5RN2Srs7TEckA0SxFDbg7ZnA/2oeKRmcnfM/BAz+y6+Hutuu+VXFh9qqQTLhQAvTa1vEtqZaL/
tImOtNuP8LDMASMeSNzg/uO0vclsN3Ej7x+7JpXGTWP/NhRYMFk6E0frP7TZtX93rGQmaANHgd4T
4o88uWEMlsD2sNOSpH4zXsVhjuSyXT+oqjD68nIqWUF/kecrEsix7WW2r9Zcn2k98Sh9X3vxqkMV
gYIGHr3vLculBvYCRMdB7/kjVCvsSadgDeWAyQfJ5g+IZNCaJW9zH6+EpylpE2vZsJNKsbXEid2w
z7Eu/Qr8bv2UmM4wbZUFbmf4Yr/gaU5n2Zh50+kwpHx0a1rrplIfwBDVhbmFywnbAWG0yCAEIkoJ
gJgWkpd2/yp3gjqaqjlo1DPwghVsclOpsgsqciCRVoUcNKu/D/PvPlNLE2ZMSv4T8BajP45xZudD
oA246jxlnIxlZ7mrvx6vyoln++q/LWyhPGWb3hTnyTmVreEuNh/qzbURUA62TS0tTac11umaP10p
qy7FJCS2aKph8+kf7ARu7FYfCWsvDo2HZHEdJ/FNdit/trn4TFmZQoh5M71aWP4b8OieGGbZOl4Q
lxV1VPWt9hZhtI/GXDYyw5BFBq+XkXDL80jKqiMgZ9dCMwBP9WDQENnS064BCQPnQPba1YMw5yCC
pRW9fwYA2bZjWLXEo/XjzYvJbostj+3/m0YMb/UGZa042tsvC57Hs9WfbmUm4rf1njg2GXeY4KOU
St8yWNQMwtwKqcnYlCMlIhwQmKMk/dsFU6RJfvB3+Gj+5TtM/zaIyQJcfvc7K+KsRJ9wVgupGWIw
0lQYIGm1YH5oj754HsDdgP/ogEAlk/PW4mKTKwhCUkgJW+Ut934afiHFsYO9rDVQ6WceU1rzDDlo
uNvydkmN+6H6NGfIeHf03NA/ILxHDTmATZDv0z3JlwqnsFzb6mLbOnUoWXp0FaJvpXEGJxYfp8pV
HLs+Vd5ylRxRVwAK+nXlZtjzmoc50x3B/zv/jeHtE8HY5ah/4eB53GsZ69BPlBKQ58g2ia2aqVLJ
Bn0UC71du0mgy1kTEfL4i5WzxUyFE7l2hAJymoZCaLzjsqhjoKbzUGbuvH/z6dSXX6+svaK1b7wI
RpxuR557B2TM6yqSrO1o5y5REVVCS5wlUu5QPMBKWCI9Q2QabuSu+7A3Xd73ZTpYmbMVxyXYnCJr
fYggxRXdBHz+8A2+oB12OyTBIhidM5m6qkCHuiSGkx7wDHkoW8zzxIFWsVTH89DWVkPR33n4/rQb
0aeibCD76s9vLWEGdcX3lThd0/bDE0NIv48jEHMvMUJPtb6rj0tCfMl+xgBFyFWVO1fI6S0vStXm
fFGkdrxt4XXcD//VihGJJjeMd8eB+9gLEJrQPdMQFrOMoulMv7Wgwvfk6MMH8FspbGZhaBBa1tCF
gDZRb8MpP8bQhO/G02dv6OaUIG5Tk0nJLeBeTQ17m5uXaSJRnRJzWQQXQkUW6omHyX8hIsw793LQ
YJXCv+v66vS3n0QlonnIPSzUHLw91sAWKjQzQzLIzZdoRm6MbPq37w+FbYuGK1HL40t5aKJ3EmHI
7QyOm2BMQVXFhVByQ1cqqECNEDul+Q7/FyyctJTgvd8jJulg7z04N0xrlTOBoEqw4e0cyEWzhIdE
DVWYLaWbe+fwy3R0QAuvv55y1T7RQgxefNaolGI5/NV8DmJMOPFyfgtAN2hJkvUrcxa5eT1vYydr
8cUgo0bhvcugzKxvWlJW0AzZqkUrRGGgLatDykZVbFNzaCxPNGskRsDamqJRZITNjAE9C4dZyBa4
XiaRGtrNdkKnOBBoTUqYqvqSI8/2Sg33jmhRNnNQ2g8Zr2CgosmqDOsIljFXL04NWvYWyzVVXE/x
xCzVq6ci8qJ2XLgWdFYqJRWBku73Jz603kIX+BcNIpXgTl88fD+Sqtq3lhKMV2ZHlU2bXkmMyTT3
XUOuVSiptT0arQmHx9yp36IVd+xfJi8TvAgkAyFRqbaAtUOm0Txa651V6aAIjs+Rw20FJ2cNcnYw
KBOtSjz+jwTCykaJAex2BWH4L1/gmj0kDJHs9ijA0ThJyRq9lP2zcqqhS5ub+ZJUaWdNxUXuhb6s
9Gx0EQ7AVy8Aqks+nePvECjv7ipZazdZyMT1U0fngiDkHLRSfPzOA1U+F5z56WkNBC46LXe6ZTe+
6EM/FvtDqtETwxnc/bzNyHQR6CVFvE0j+8c2ovfJewan31vL0Y4nbSTsP/4a8jvbYDv39np/A3HP
MRX8BFaMeMZ25wnRnqB0Tf3xALprDNYkPmJpXU/og/dhd06yGgotJaSwCFuE80OSphedoprwBygY
sljOwb7dQryA0eNU6BxfrEWXDwCe+wZ/Y8vb+8wmDM9D/ky/lCdf9MouCZEgr1iO+vqKYFavlVj5
6PQHkEkQKUO1sUinriaxu91a5P/dMzUYvHzYmQABu/h53I3XwUPSj6o3bGC/iPCkR1/wCAidih41
VnYQ/wSCK2bdZgCa0o1TmU8ok8PNCiLylCSXXtlohhK1UT14EkqCJgcIo+OdOuvO598AWn2t70mu
he/blKtsZ8CGYOUHVE626JaMRgS/jn6f+Fyke/jyRTb4Jd7HGGRZxQVEDo7YlwIGHQQCbCsxNt+2
hDmC5XFjdHWI34SMJPhz/jPhXZfZDI5cSinXIMS3P8MgYyHhgjybZ5Q9Oh//x1yFAv9F6TyZqwVf
B0OhtUMPHIm18StHy/fchCEepjZawM3rYaiAQO2xVVIx3eurjhG+1QkUr38CiizDoeDgGydWiCJh
dLuF6RF3EvfZNPqSYXrOZbSUrkmEQiLMw6vrDJLFRNuNSqhv+bNbIdR9cozJFQhegiAo9B+patue
qqxaaBNH5PrYx79O6FIbdwFcb+5xZyYTI5uHvTTA5xu6z3KFivJ84FfReyeSHmZq0EDgNV/Nqvvw
txdGrCc88j+RaISFDH91WMD5BGI2axT3+0Od0ALqTnjVAFzf06IOrU0BuR2688LlF0XU08pd883T
QNhPrIdYaxqfVcdHpmZF5zY+A3/o9BvBgxp+vBHBgv+qodrsOlMX9CbX+ARib7O0XHLGGu6zZqOO
kLb2FgHp2QnwxMJkxAIuCqBE/p8QNjAUvAHEq0R/aaVL0J2Kyp3kt2Wt5eeQjARBmxOBKvu78H/n
DCGM4j6DJfbT0iVWuCladxudbH/ibHoUli+MEcC5mGEiS/5PaNePtsoZ+Z78Bmju3LKIEAcXKq/P
MVq8hqJDnvC5B50e3bMdCm9gd3ZllMvJeU+7MB7kHuJ0Iv72vlxG5tUZxL0K601UZIF9d/posu/O
7u9SeE/op5w8PeC+SD625u21xZoD12Tv0O3SJTbBA8MxkpnxLx8zvUaReUeEuXcNO+hwv1WYg5IQ
xy3sU9yyZcearycHSHBm5ZhSlRAsPXSIqSgsz4CihNowtlX3wLtx8Yt/rCNO195PnN05mDQU6OkH
S6F3xbU5hofb9gUnNSR3iUf9nqAFnmFFK7zH2WvJL4N3Ntzk6ilfZGISkGT96YWpHLd9d0hXlA9H
ZbVG2PS3ESie2Lmb0iSrWAc5nmtc/QeI37/dk8o65yDhgTG/JQb6lKYi7QOSZ6KIJ4tHLty82Far
B9KFBy5+eicG3/Gb9eSSSUXmLiUqbOcTd2U9F4E9Fvb3fhs+9U7XBXFQUC8019KKdSA1IomOIw9D
wgWhXj/0W+BlYE+lHQsL9ZTcGPeAOWoqBEngPn9Nw8upyF8fRl9LgEwlLgE4qAqKV7lYJxEwXT9S
2OED6l8KlOTPWESY8tK2OoUoOld9gZVb9yTkoAhYfu/vC929j9G16XC5cuseavShNVxhCplK6THR
ZEnAPDO3m3cx+H7q0QEHidbO5XKj9UGJ/GOb1j7W37uTmxe2dDYykE2eIDJ7V/v0fc8FG35pi6L3
et3RYVNTJiUQpD/1+2FcW4E0T38pNKKQoUqeNyFgFokT8cLpXoIfoBuWdp/l+jBXKpoHCwXWITnQ
7FUQFXwXbXvaRBWm2597GndniO3OvLlsEjRk4Lhxqd8i//5TrKDMOY1L7ZLBNJAW2pp79KQQiZxN
1l0FQ3F6tC45yzVZ2HwnHLt+1V3tBfs4rfq6X5XnCCQ3OQwddS9eFMd73X41D5P1J3cNki0A4f7j
rmtRevcfwb/arVLgheYWIBHsaxdtLJJFJ33Fojcs23JTNBx4OYnwzxTUOKUGP38kLx/v+Gjh6JTb
qdkFUhJZ50XmNwRwxuZ5RKJMAlKLT65+uYLXIO0TcobZDruJF+NzS8A71XFSrC2KLW9P5e48J+N5
YjiS3Cimb/kQx8Juw0qg8G5+RDxca9bFOk8XVrccDzy0aVn72PaGLshz3xJJyMEYIBA35GQ3o6Uw
+D2mtnw5xq1ZQnbMmo5t751IGZIW3ZOesGurFdNQQaM89Bxlcd7RcDNeM35MFy90y1M4GxVdRHbf
qryqX1MaYG5i5FsJQO2ziohbM3O+Z9VpK4RhE2GMNjRbhIjcl5ZruUcDpml7V3Y4xbCv32msk1HG
TtoAGR+GkS807zoYFXKc7dJwUQ7jupArFR56DBc5R75dZgWnMe+grQ0GaD7SoSALQIigTHkvOgWK
8VK2xrIsMUocuYPz+Uz3nKwNloEsztKADNX6UP9XNAh+KabGF+7+mI1ZeDa6Oj9DQsr/96PWvv6D
IxClBo5+2s4yEHZF6hKKIT+NLOCWTh0ZCilKLWcYwh6vBq8I5y7RCyjkf3nFSGE37Jabf90acbNg
CmPgZeGLKWWdoWoQAvsZ92mtAUB1nZcUo7c191jLUbSiiBh38KkaH2YZiwLapSTOaTkPZL0arfmf
e9whzpUTXZ8hvnb411iic3apJnM8EIy1OncL5CL35Nv+lqh2pEE91Qw8dDnkS9d3RxEjc1IOlxVN
2wExEgMOMgSc6sNVkyw4vP9Td/8p6SpQuvnct7dW0lopTZ4smVFsYiBjvNMZs+v8vNthNRwgliXJ
xdbVk/JWKSnzAFdKmWvmo+6SXO7GHxlRUaV/Pmi9uZfyPv8lwqqMRwLrm9lXbh2ifLcX0C8IVHG5
j8HbGJVBh+ZEmQ0kf3FYdCdw8oDHBFT1YQ2RHWnrfoJijTV4CGdOtQZo9YpDZ50q2I2aW/kjRDdw
JdAC45PeWS3+NLbTWtoNV6AX/oQy887fgL4QSnSS1oYo8L4jxrEb+fq98d4JuOQUEEIKcJUGxSSF
IOMRDPAY3anbAyXmVORW5jxx6UY548EXQDnk0vs0jBpeRUFjg2+6x05tq/EICG1Ord9eCZ+Pw7S6
nJVI/RA66zz+QyznS8/o8U9ediu9iNuXfYYCByHfxh2+A0kZrfqVNmtJl8+2NAFBjA6bg2+lbHN3
FDOFqM4VOAJ455lj6HT+h6W8/FkSsBQVM41GjrBBRhaSsPUrCcZHBUW9FPrR4HoHCcFDfMylsvHj
piRKj4wGWTLSvxvDuXuf6SOIPc27k7m9tsn1ZZhkfNfCi0PwdDDMYM9Tuyn5y97Lca/vpxBY9pB3
Ga8H7a76qsFpNHHqVShP01eX1Yw7m1UbNMtUePirpOWSlzGwELW3wWgOXvw2iS8LTL+fE4GoEOQF
D4eSGVu1Q6oKr8Nk0MJw6qPzo+euUaYBRzEF6MsQDwN12DK556HWZrklCdaUePMm6M0Rf8JeJSxL
UeeMzqqQ5cUecv0fUxxZZTUyBMuUoJ9lzB+WWRHPgGoTznX+zTG+bnB5rc/psd/KjcXfiyj33u4O
duYWE2EJ/XDeSwj6gKWbGlk2zK5lEdfnDopGrkZAB2BDFwahHT3GM00YSWoetbOcysyNrsojSiRo
oVc4RROzWTgMIZke/fOJE8RGT8jIzIelkp9SE9igfKGXUlSslBrZJIDtChQphXnlWSYFIv1DspP4
h3iz3NHEyOx4YuZrZL2NIeK26v4qBJOvmaly5KTnqRr1J0z1gwc3QMPleIZx+BMQH1+piLvqHhkZ
xI9MKKRkovseREWhpOXcGEcSAPhWtXKtAgL8dQxLoG+wppZeTSWNqiaKe/L1tNJEdUl8ho1pDT1u
HYvbQ0OPK7e9aA17UQINdbooNvXdV+HSgi0M+S1hx7TEP9YRSaOJ0GUon0HqNzLJ6AA1tmtz4c7X
UKX+zbkisvQfLdZyLRONYV63G8v0iNVUcmHdmNO09tCcms7DyS4P82ePLBJ94pCo4zvaXJdnuket
beraFQBzah/iEkSdkg5yupEKR00baBu+v8wh4Pi+NMUaqiTqgmb8tVPLpm6VuCOlnN/rQV3w+HVq
2ntF9JwRoReqRAgBBtUCw3nF0/BQ0yhEyEr9Lq54rg/+PopAQvlzp8QHBEPPZI/EcIuwy2RJpu5s
12JhOlMFAUHzAR4EC9ANahnwBSTLxYX/mAn4diKQOUdQ97L+PNnM03D/qdiNh6NK6njExB/j1gVv
/9vHF02z+LA3WvHUC2kw0is6AzOBESKdccdhZ5B36vMqLKeyhMYztB1HzmAQQWgMW9Ud43dUAgfd
0UlpeuCRYu79NxiKdGwxS+JT2XH0fk/JcqT5pFDoaPpjyXm8aZVtmjA6/6TLYWzavPRKHURIHsq1
nkI6s0N6xad3CZ0suz8f/ZBELERIsrYgbEkJUnqueIpc9a5DMpws7PR1LL555FmE3ScWXmhHV9TT
OC/TqJDtpYEDDbi0yqtlXtEq0nQ+elrEl9sfMO+K1TZMFsfo1fgygs9/WNDPbfTG9p/U08MXRPbc
bcjO697idm/d+gdZGPc+omSfIaoNGfMVOG9Kjsa+BE0nqXvsFWWYFeKNdpPUHLoMoL5zUspQ0dck
lc1f4TCTaTSGnf66FmP0Kx2Diu44cDLYIw2FT4wjIzAOEaG5rpP18qU9O+HTX6lvJo+MFb941Vgg
3hu6ukIGigBBSxVZuLlNHKVhcBf0F/Es9sFdY22UCaLbyYT7pz5bp0upnPYVEK7qbXviHtm0UHlX
/zn7bvY+sua0UtB7IFcTJgY568Jj2uT+oGPn2kMnMXQDDRd3ecT07FMhXaaTj9OKtcrI9axE7ZeP
UY5ximJq3bIvRim4k2bFNEBOE6KX771uo3z0I5mhd8da65L3g8JkCeQiAZv9lzSnf00b950Fm0cn
EAH1XQlJwh57mIZfpREIMFbbJnk0C/CWAcaDsrQRRBRBg1BgKjfJV6ILbeuJMG7vq2DCQa/mmrij
Q7oLFiT22WxdLpj0CJ71A4Ap5WEWOwQKG71A+GFoRAidj9YkapvzEZRxy5LYY8/8KVnDiMSTMgoI
ogSVgYbnjvpdQ0aKjWTklu0clb5jXgRtUtNoAGKA7ybUAW+o44IX9tKgPE1qEsejsKhByitL69yj
2uhuaG9QRNd2AVAG/xXVFXH2OqSWvVKHdTlaXx+WK+Wbhbi9TbASXR+YFs6Kv7rIXt6GvLimKClG
yJpNfhyEjM4jzeKQ8xeuwhId88fosr4dVDxbHvHF/ue38nJctByYQylPDXGYbCM7Hm9MEDNQO530
5ZPdISTf4t8AEq9GAYuqEOgX+2tc31wolXRI7RdL6rMFWHXJ8gEhAtYqPS8ZIlsqnTWAhzT67NdB
r7UJgCZ04mOOdJ+BM+2FOeEoZ91oKI9/o3c5m7yklpkGnJ3rO1pvqeR4tML218x1J33KLwgYM96w
sqVNVADUJx0zh50N+VS7zoUYSDs8dDyqsuZ5NTkqN+nREM/xz5ZW/CU5g6F1uEg27XjnXTOO7xc8
k7x7qZK5Liq9CG1Ot+dTd4q9O3yHN39Jltq527z3Mel2zKGThuqwaDUwp0YBqnhTPjXktMg3nBB2
GhjDywi8uVnW3Ya5jUdFpIomGM5jrv8tEgUSfAFmnjDdTJh8NYbh8jQVMcJxULd9mFKQ3Z7gtoKk
/QxVzlj1PiXGi+vbWsg4Ylp94+NwGA1ukYD9FysPl2PU9Zce31mkKdoLo/8SrBAwVis6RTJPNdhj
lrn3ubNZOn25w0SaepcSu/NUOehst8Wd1rHU9NdkQ/mmhQMrSJdGV594KDnkbhPNRKVhomClaGZR
ymJSrBCGyTz4KGZmNHvhDICoPEVFsE5WncWDLVEVPqVGhFnZ1VhFx508uO7j/mu5OmtCvAX4vQUF
su8+J78zDYoL+ZbLPuGyLqI40g1l7kRP4Lyzzguy4CYKb47gXE99613oxAYi1HDwGpNS8xvu1RpM
4DcACMC3cWM5CKoZdGy8QeztkS9mg63ZzcBg2w2f5bU4CdGIX3EQe4aRlfHPwkz2IFy0HH59B/r5
hzksPXjOvvkKK69W9c39Xwlqd8FE4FwmBvTI2R7xBZEzOm0zO276TUkztNCSWFcMATpXRCyMdxC3
COtgtYYOVlgzlzG0B1FVSwlrFzNSlata0LqAz/m44TCQ7WNtsAuiPGCszNwM9oDAqy9QihueZhdG
pwVxMT+KjcD79qrl02ZHj1OWhKcmKE9j5cIwA1kw9IJ7j8dKnUzAqj2PtBlCCTRpCK4gnHfjpVbF
zHj2bV9Nv4nmhs124g7hx6h7Ac9VahiEXNieh3oV2+7rtWWG0nl6wfPSxzWNgq5GKIgR8mxodfWb
s+93qPi6JhbFWwUgPvsCMRAiZQhDhFNMJuo//3nRctD6bLb/czLVH+wnyV1BcjUrlg8XYQdO6Ny1
B9GZ8qBws/6Iwzia+EVWv6ht4nHP99qAsMOvfevx3dt+CFlG+09arpYjuxrPmvk8cPZQDsa3cWPu
eSDj57Dz/YTMhsCPARBCdwXl5sF1+YFPIKb3sdmI8EER3gtOr3JzDp4+ITATSg4Jo4xvU2+vKdlD
qbgviuB/AuVoU3rJ2gfWjGi6aaMyXgur6gx0GrmTWncutZA9kzTKXwgbBB2klgNp4wcWUTSlXd+z
Mu06eLAoQ4aXHAfDpWcfEwNdNrktV9chtFZXgrKNecWImcOPf8ObMvXtbnia7trD4cPpSS37W0vI
GPEc3P1l/HjW5WAlbWIcfexVMPxeo5YRTmBxYhXHsm5pzydgCY76vdaGKivOGomdBl1CKhTV2c1M
A5fFieKK0WLk5JP+Tzx94yEFKawDdOksx9Jzi9a9UzIa8kePutj9IFiuuxhyYVBdtQE25WxB3pcO
6VlG2qK+KjRy+ND+OKrmKLIzhiqCofMaLrK3JwMeVLtNlPFO+PAv1RQmGsrtHdQBFZR1JZUmzm/i
lCxMWxA5vrZUXGjfxBjPGRRdagMCgGNZe8OeqlQ1Iyy740flx8VAS+QVE5erJ3l4QminSEFG8ydI
FsqVdqB6MKFVh/nbHsgC4pvj5gf3bcSFMOLl/tNf8sU7GZ0Dob6Gnoge8rln+5on/NE2YbSqYYnz
Tf40QwzYDs4EU1zevova1IbBLUbVUC3zTld3LpMdxhq/tCisShxziHIv7N/RDF+lLtbIMc7STg4r
m6jZGxvsyQ9WyyGhcoAPD9QumkQzabRwwmC23Q+qFJZ9BhcPuZfzTJznEscEXFnv2qPhcsVsJT9/
yfkVsAwY3kyOK7F5b5NXF5+Yd0YhAbkCS6VVbeLpUfG15dhI7o2t162OQ1TycqogbG1BITx1v6ZR
JF1T8PxlXsDQH+GThDYUWW8pIJ1Y6+YzQHiNMnvBH+JSW2mBezEBcp83gFHdnxkBJFVTbzgZ1sGZ
v/rcJOKNQSore3tyXhtzFwSEZoOFghI/BW7zY3j2eSbaQl2DZPaZXWH1uLx2kHiIFfQ80DewSIqH
5znYsubjD1fTeA7wvPy/zKxqhyvZh/LI4CJ0hA0zNHazre+CKDfxGeFPgdA1xgG5iUzByxetRXl8
/FSUIBEc8q7Dp7YVZj33SSCUnG3dY1tWWrrsol97NY2FBgxHLx0V6H+bAEPwTpcoavD+lsaKIDSQ
U+cT+9+tDwCTl/1IGiVihhazbIoodmTDDPPhMXK7czndyfOc9Bm8QtX/v9Cn4YEcPwNX4pWjwhlR
TThMrLpNk7o80VJa4/s8wjJlVUr7JwYT7W5O4OcyQYCPa7aT8T0TL4YZVxaySe66jzy8uXlvOTIC
Mh8yUkqD/z7LthJ28Zez84EcW4jeKWZWghFKuM54AAbWT1o0ApfQigZnoUszHhXVkZGW8+3lO47h
1qJDwjl9Xiq46OdP5+23IqLPJjeYaeXG/AaDcJSMBXtooFy0kz5q25grb8QFdX4SRNT9Gs3YsFuV
xZUS5CnvymrcvX1jiGZKWGOO5xHVTwXS6FYq0NXrPW0lmO2626E1aDxqTpxkEeaPuQEeF8ElGFQK
IKHg/QRC3lJT/SIUVyeD5rn+/4U6PUB4eraKUomeAGm88a1qugx0+c0s894GY2zDGVPXfJqOo2LM
58/8xhHbHKSoTIXBNh3tP83+a7xq6HXcs67jPOaRe+gE1y9ya1log38/Kl0ppt9BUDH/5/Bwtvn1
8HHkPW4p3eXGqeHQAABkB4dIZQJ9yjUCFJWj8rrB5ATXXIQvaTJJ7qYZPGo+Plpj4hxFMp8xpS1D
w7506Ey363XI4N4+LWpDSM1IqaCP/zRUu5H/3OOFNXdTtiV6poucW0S74oyoRA2xsjSpx8Wv1j4x
zKInu+iuAJMH8N0Ea7bA1MUAExe7u5dloqbfmjKxdu2AHVgWPdiOPU3ARJ95FLQq3yOXWXHQ9Qqo
tW0ORevTHhGlyl6kmHNkQeQNlOVo+27nitPFctBeF/nsZxO0k+qT2WbU5mTh315dBjXAkwKkGGav
kpCgw94lop51jJ+ZiMHZXVP7opXTJaHCaswbXkG/l7UqUBkR1VxZNhYKxmet2Z5mnGDg5CEvXPla
+R4FyKSFkg+xLE6/KQzUBoYpOmmdQm72Ls6J06eCUAqGsydBnnLBMUsYJyw3daudu50eKPqk6BDe
eAxZpl1icAkmzT5w9YNe56XkUHk9bN3Lm9Z5uOr2vViqXp33A6YX9IeXCs9cwV4ZHGIUoKTO087f
UcQ7jCMp2trYmFqiFaVbG7POXhg398rbWRlj3dBVZ98IGTFHxiKjiUObh3KIscNvBBUZTvu4MWr7
iQyp4hI8X6n5bVdIsUG89DVbaXreOtZeU66Ilr/F7aLN1/KwVl70V+zciZDUl4kOLmAia1VXKHCz
Bg182KlU/BBap2J1HdGV0TiVPom0r74RgvRV/nXo1A8jWc5Bz963xJ6S6ErxR5Bcp9zjdzj/A075
6Ik3bI3Hpbi9s2XoIxrVI2ojj9LM/AGbwocFhE3lE2PxnDPWVuOZqxLNs7GdBmbgJYHNv7UcE7iS
DuML3o+8N6X4KvKLXNXSYrGUuwww1foAxrXXpv+grpLzz5WSxOBoc1OIl/oInbxtBGRo3MPsPY9I
orpFlisjSvmMzX6CpuFgmajHYNsXIYdfNbR8ckEHXG9QFmSMUZ6aJguqO1GsRtMDJXcCWqN1+dSR
RDyWB6HbG+kc1rmtE2oHCn02dEVtdpuVKSkwu0o/bhS6TQ8URfrVq4T+FF9hBZ1FPjZWUG0CTtVU
6Uh823npZCCEUA3Pns4cSrfYb/ecwZGJYxiqf3FJ08nKN7qiBY7s+eHJGL4WUHTu+EwLPtJiKjDQ
uYj3RABNVJe5osXrDL4qg/iZEMcI/KcvVoEueK2b70/x1v0CalWwocn1jPvrpw3h8kMHXu14qDU0
x+aW3h7wCFOjuyBFsTMRPSeD0Dmzn9AiHqFn/yrMZvXmUNLRUYTjYuPIQDdcXzyihsKHukhGYXeV
NILRBWtfIZFYfj1HvTFS6c2Eti8O6W6e8VJ50pENsAZXZy13NQS9El/O2Z3yvqpNX9zOVW2cYZ+k
B5AGBFI41lyXGttERhB/QfhD9Fa0bjcxnQZ1GSClAs26Vs5t9jG9ROKx+8KzTREBT8k+5T2XVORl
KRfuqgqUED3NFYRu1L08kEbGudv892GG3zlp4AhL7ih2piWrdIiUKg3u33Vguoq/FnjfmF0GOqTw
MpjdZUSLOBvK6gGgwkxFg9giyI5/j1uJALzsqxUNY3jClBzLJ0lWXmXW6mydxhNS1WA3fLtjXexP
9uNvXQZd7mQAfUdi2XdQZemQNprIeOV/3ZJLmLhCKAQPqWUwb8t6O4ywBSuhqlTNZsfecQPzDZ8J
QQFeujUQgdBn8ilYdIoqcF1tNNrm+Fs9x5/WUrll+6TSmlXEtjs95AsV+uSM4bjeuAgDoZv16x/a
S9N4KplMXjBUdstowGbP1yZ+xCa2BIWvQ+lGToS+0Db6DlUvWSIyjWVuBy5/+Z4GrBtvqgetrWBp
pf+5amCxJ26Zrwzgo6sBN4ydtJwyy5Z2DqkrpD634GBfZTt0+WiwDypX/r1DEwFfqISZuqctDjKQ
8ME/y+w5QYTb2u0UzQaX5Ga8F16nyscUplmnjwWdVt+ku481SZwCd54nhRxQvNYCHNC+3LpxP3x+
qdnudiksb4E3NdkF6pkHV2N4gSCeQ3QcXyMNuXtrpeYN2sRLVAFxKurEqk0ybDlgoNO2rQFf2Ikn
+W31n36zXhDiTRLkjJiRRX3xxHzOq/cpFIfgRWjOoArHLxwUHibpv7lrBsC0HuvRSY0m0VthtbpB
4LOX6bXDOZMH0JINOdSN8cLCJFFpHhUPTKrsjatWm1StpLlL3HexYYzyz1zdtSA6sVfny6yoIdvw
1mmVZDzIEA6zs6SyF3xYbkT+bz9zeonNASzne91iCRCgsCzWo2kFhmu6UmPJTISnTot5G8yYWk8q
PMPfqrB5hFvxOwI7PEvO1ll/iOOAwQbX6SaE+17gWGnq+xZM5O+GChhz8JxWZ83z6SkEWWwXfTMM
adxDTK9h221nXA1wKuw+vq+kKuO7plzAclaroyVa1iWyZ2EXBFfLEzz9+R34NgkKSoVJC3KrntNy
LIJ6r5M047SR9Su/SDW2SaEaKmMl4aP9fr3KVCqMHjEisgSiQ3H3jiMBcdJ/E3qPZFMMgpmHqO4M
m/6kvduI/7vkeTlq5cFlVcivCOW8+IYR1nTAVyxunpHXzj4uBxvFmDBWw6fCQFqyHTb8Xad7Xokw
/hRrICw79MwfcIhIj2J5fzagmaqX23XNKov8fJapQk5/itqV4LIQ874qtrgZK+in86oywInZiJ5h
xx5usyHIAbr3Rl6t5IXYm/EXH84GzPUEFNHagx1ndMPSZdamEe+7LHRh085oW/BnwQjKFBPt4fu9
oUVpAJTO+muRRH9TeZ8EM8eT+Ey7/fSfk7KO7+WmHlfbzLIOgyluFqC63Ogj1WCTXb9BeyypQVda
U+50mdUJdgNrZ3BpGFt5olxkYAKn4Wc5kydFJcaxaUkJPcttPtiVGB59khVO2zpf0DEgzuWgLZB/
NWOlcHASdrIUQWrz15yxOb4CvJruvykk58P0WD7RsVsEes3++YbAvr8Nx/5j58g0Wn36vfuco3iW
mgxalK1VKTOxWKGc8adNeq4x8430DQVfkourT5dyCv7NcP5JaPAbNagGNefMxX6XuVxbFfzOgnKd
XUm9ij68iu9oBL2mb9xBpMTf1XwsC0Tt8PHpxejXZ58LPXfMUr8uMdbqhl3quEPAR5nWubzsgcQ4
BKWZpqfhq5ZQ1jDKQbDKwtY7yIic0XnMUTKSh4OuuAzkDwly19rCJAhexFerulHra//dhxhU1wSO
O6LJore9saSjMOHhE/2rZ7aaGctDb+0IzC6pE0/Vj3Gow0pzrjbZvHVcVdrhsUu3tAyQYqRB1aJd
QzvsAs7L+OExHNL6DQ7wbBcp22eLcAT6uCvSJHF7LTGyI9EZiyf0YTfjy1jL/dmG5QyH05FnEDcP
m8EKt+TvHQ4qhR0P9AqABofD9DE+vFFH/LblT5x0de780KUe5ywAhI0vZ5rVEUf24fhEkzSbcAqT
lE9qOoSIoWn9DSubRbdk3tpUvXW9oT3tQBCzjhBnvCwmwTX+v/H3ymULsnwEbCVABmJxFsKlRhoP
eSB/8CieIaq+oQSDbaTfaeF2/S38fuW9admngZFPXUAiufJJtfJoWBevrq6Wh+XgC0dZJRGa8tyL
PQdjKy/jF5gV58waKdsqWA5RuDmj4FIHcMKeVjnKei6uxIOGrXS5Aj6pYzQkMdcOImXLEfT4Sk2x
CRJwtwRiWH/+RTcRqQEHDX+gb0suAMEFw/iFRhP9+08AyXvY9dhFrQXlDQvdPE2NcoqcQae/KeBD
SMWHYiPFsCfPjP+hfeyYQYe6VWtNIe2pPKIYwByXfVUHxK2gTdeim0c/6ILXEz8cN5jtv/1mmOK5
qJ7JY2057NPhrBhgVnNRtPK7QzcITMMmkPTz7Frrc3fhfpAXR8tJyqqmq1pLm640LKCSLGRPw+Wp
S3mz9Wv25eE5cXFYjlyfnm1ZhkIUI7XO3Es9PD5D6DWEFnwYpNnRwKQNJTIVOttWHFdugLJm6HlR
6BVmS3yJn54vYl6zZy56aEOVzUT176a+1WNCLlqjMYUmgJII83wcS0vtJj/yJZTdHxxCBZqosOY4
cqbjp0y2zdg53j72cIgzcVtxa4yHpQT02EX+iV/TgADuNRQBGoNsJGJNpR4x364YPm/XFjFK3OP2
02bTTqkd/yWEK8ZjpjoQiCiPWS/rmUF0pj1RhdMwNOUgrmbc5hMOCZhq9dPBl4/vSZSW8s8znBw8
/9vO3wCIvHKJuuORvAQ4lz0yNsDdm17C5CIquuW0CWN0RwNm8QxPUMbBiJGxGfyOFJQpItNPn7B8
VXSBhrPTFja2ss2F1u3tki5JRrqZfUIb7qX9+fAcTaFKUXaotemBr7iddaykV6DrZieM9XohQd7r
+o/lAGdT2C/BNoTUdJMYVmddNlmQSN67DFv3cZJe7XVIW43EY2DZzD9sWd2nETotQOi4f6d1nwaK
w2L9hidU+8RasU70TKdz1UXlugYq1EC6Z3MlkNKfjQDT2mS6+v5exm+UZTEUIm573dWevHo205X9
364aOQGV7iy4MTqD6/6ytby6KjUikAwp/MQQy8JIoHtRoGvsLcV1WcL5dCvXZFmygus7rJR9+BSA
23xKBzGkX/3boqE3YToM72Dy7bf5M4x7RU7CVBck7ZvqRuALLMXKUQwSXbwKNKC++Riw2ExemfJV
bEfKSAo/vdHU8jqjuCydhA4OEL+NJhr95Q9B9NBogda+oOv7RFLWzKPIBmCm+NxxoRHxBlA9ICQz
ebOVxc8bSPeoWhGdOODFRF1TpIBICqpZ28aai4EOakI9zk6gkhiU98ZvR0c7Rawo+MS9mSM4zNy5
hHtVN1WrQPyg3znlr7zUXoltRnbB4lAv0yoKGIiGuecgeKlex5/jYpeLrNVdFcUyRzIgK2YKRU0a
ERqR1HagR2bB5Pk8S5ZlA9jAmjOmEsUGqFiIZgXOjcspMPMzEyuInOMvc8CWXeujLbdt0RCKTX+U
9h33WUbb1avfy/ZjEWjBcQP3A9fw/L94MdDZAKacbMorw9dfhIdj2JdA1CGAOB8YHRvE9Xk4Wtd1
55icxrW0B+YC/TQaR7zlrKtwziR2F1Ah3n9ndtuTFpwZi6u/XEFFnbzfip/2n4LjrJbSafMRMsg7
VKx+8pyKkfUhYI8YMgAoBGmHvxKc0+9l66JIMe92F//Gdfl2N5gbNCSxuEiAub8MgN0pLOVnLytx
jxlaJFcbFQ3nMT4vdVhjYI2p3NKlPIJimw7ksvFs0t9JAAUQUOLn8nZ+qQbk3wNQeCDQZPEjNTXC
dBBfM3MqHzspjthWbzWzmq2rxRUaosyONFxXtM/jMThRRMkyXYg2gvb4G/mwMgllNHUnfOCsFSEZ
zPSbtcsjatkXV1m3oODmLtZVERIzxebnNhxnhKbsD74H+elwoV3Gs6PjrQLMTaQ5R7FFIMhECNNN
bDRYd5fMORB60AvmYxJxU0fIcqTZtYoojTBsU0wTL5VgmV5Z2M1krfwPAukI9NQ0hBpi4TYOHcRu
16c6sGoj2N9SU3h3bsOFZ6nuC9GnbzVgZeVccgsJSxY1bCnIBrZJg0j5xC7a8Z/nFw38fPkBPs6X
cRhZm9gEwL85EPgEG8VKpxRu1ZlAQr8MT8cW8sew2amzLaGpznpyPKvRqHPdKHKadZtZ1FROigXM
sycuEam3daEAueUreQbXCGU3QHu+YBpKpMu+Dg5ewNUi05nyemGsnT6ZYw5aDnnMzKzygAaT/Z2z
ikr9xU5lu+KmV15rJ/BoFX0lNwej0dln/s/Nofp+D42fMwMQP1CaIZqIgI/aSglhFvKAceuS/moq
Ji/+lexmnddcpHgCUKTenrQwsqPDTkruGNsQlP7dZ57dckBa7AuNI1W8aSWyhn7/w0ZyjfOBO75N
wmoPMV0MRU2RcCT1R+DmyRyG8M2gsvRudrsMoJ8u79tMvgSA6MQzXmUAUxe+h4FcZiyVo962Oxov
rN/tpOPEJmwOA8Cd4gZFw08x9DZWmpbzjrxFM7qp5C5SloxPfvxQIOhtjpmnOb0/EhV9XxkNH2Cc
Hcuwa+Lmipxq9O4k+DJBGg0wECBlTUCH56f+9dLKDmzA8kfl4utcMCcFv+VHNAeED+L31dH3rrU8
CZh7UrpAJr7vEhFmR+kdAg1Dyj4Mfv6qEEwqTUTvmd3ktNhspQUb21IQhh9pDVtcjcJc92TeMKrb
1YsBTJXhPvKS7cnCj3vKTBzEE9GLUcqugE78h8hGzgNuWloo9tVgkR3g8BmOsV0NIrm9uz4wmCDD
LColWfNfz3wqRVsTUkSc3abeA3OoqidKOypT45wBiyAamNJRVocbBypM/xk78QPP5rW1kffjm+Cd
JOLFhibVE+zaPaJj3x2vTKzbp35xTBUuGKkkpk2g/GBo1eWQPHLCFYAsxUYZc0MCrw8Px9UBX7j7
wg2URkRAfbjigOz8ceFM4zqCrVtxW9LBNa7GA4+UuhpvBTgRXMXk4zf4i6gt9APkpuL7Va3DlDtE
HDxMn1nM22sJ+WBwG3VZ9BKJimdpw8MmrX7KqBH7Mu4OcdLWCbaLyOT4s2dUY5XtMtJSgkMFiLLl
walgj/btLSDV0AGdQjNcNXLcUfnXW7Bts6GrUFfNgfD/WZI/mq/+R+dt2SiwSFfushvVOLQx8EeJ
05G2+EpSirogTQZfFwApOT2iHqHyjM83jj+GN1p2f5zqIzlA9MW6OlibgE0evKW3U9b3jnyeNrzJ
JuAzS/r3VohjgkSMF46ylWYgUP15fkLa9/8qps9P5TTGhIMyhqRS7/E4C6f6DnMLe/X0Uw9c/i6X
2ugo9j6qWEXVBrJxn07SWy5n11AIGCOlyNHhgZa7Q7mDoIbVvx/IZZ4mGaZW+h29Mry7HPW7wOmr
ojS2/9shvJZPjQgH5+j+I/zg2k8QHsn7jcTk095VS9Rc9vHf3JQjlnmC2phZrOw2mPnmj2Vc3Z0E
w6q5A+nmkWAjKZJKdJbtvrJxWbdKEQlDqeFDyzsLxzJGhKq96S9WygqlPi2B9UhJSb8X9cUvFYP4
YeUNxXW5RNc8iC2VSebGGZOF/0CvXIlmHi9MS8vusAndD+fNS4ZaodfVuZlqHTlusy9FwMXfBftQ
I9VLqtMVLSlyxxhrRGOirw3ry+jSydcmYeAHB3bjR8+gO5NyLT79SP5pdat20za2qZyPuEOkOyDN
zU7V1VGChBmL3CTt6qmIQXdcEQiv2w6HeLoNbUJPHZAWIBltOqpjkOXUzM5EYAxOc2ikz7wr7bjS
4W8TVti1MqsNs0+qQuPsSBuDf1tr9tD3Tu5d1vzH1wm7FqVAQ3k2r5PiPUOxQZ6iSNkkUyaOBjhh
yxWCwoj01o6nGMs/ZQ4u8PGOpANH6Fr/mHoa1vozW3xuVHvnakU+3HggIJI7q/xTlKIZTG+L7UME
LH3IvrKPpmrek1RerCuPL8SW3TeJGYOQM9aF7iYBDRrOy5vyqYclQE5VH1edU0LgL8BpT9lRTEX6
Lnw5hhq6WLTO0nWjDJl5kzT5eK0rlTGUnEhT/IF0sBWTiYqGcVKvsqlpLj8VP2UgTGWhDRXQU2r9
LxU+ZlvE7PMvBfLmUhb9mRvh4a1EfdQ6TTpP/WoJpbpv4Lp1v33EbWCMkxhH0c1ypBJqq4I4vKYO
Z76CoMfO4xJxK4HXcelJve64VIj5x/ikBtqMKvWI9tilNrl/DAdoG6DvIqnoukTtt5mqqmy3T27S
fMpLyZsm0gbzFioM/VywLLwS00KQaDIGWx2QYz6pR33cyc65OFcfXZ8iTYqR3/YPtzx6RI/l2xgY
3zOTJzPuwiglNbcrwWD3z9uYzQ8OioShI+53lPTbWqlaNhNNXhjC7+cHmgxPhM6uWwRiy4AcNzMg
e1uqdhLyUSsgeJ/C/GNY0g827fC2ZSz+B5O6mtl0yCfEujoTybXEUt5pBHsRq1eW9M44lqyjETRk
cx619D151P1oyuELUSqzY+o+1yrXOKYGVOOyJFLkhhp6Rv5Gf5ana6GDfKKIw16zBGyv/CvC5TVH
VeWk9vJhDYhI6l8ebC2dtMpu1lA89dTyzguOuubJl4+etMgqFngSvsK8HAh2H2DSFaumDwKbhorh
oj7pCRuZzqiqDBWRypCZKNEouua5j5xKAdYRM/bxx9AIYFvnflSxohJwj0fpgU5bdCVY+3WT8tYj
QduJWwfA9zRBq0Wpk96idNTKG8MKv7lqCS3TGKgeY25Ie2gjrkZlleFxNw7kEq7htitLTJm2Dakm
4mUoNyny2ZJ/7Qwjli7AiUOM+WwMw/klZNoZeEYGIR2wIvIZFfd/1rArTI/4lmA07FhlYrwOuY5T
XZyyKRf9ly1BUEdU2rFbaWgILraQwE8CzvolCgdI5A6TPAwsFj21NB/6NeGW0E9NfliVd40LgzVU
Ae7uMVlDEJotC/H4n+67BmRundNUcWUEFFBt0BO/rBYZmsyc01dcvj9UeQBx/zoK2vJLoOSuixqa
cIa+o3sQ/xuxnRzcZIfF8AVWVY+heS1k4WDpiyDP+Kgb46xEb6x2Xwol+T3sX9kRthtrrQ2Bixvq
K5zW/mxf3m7s1rF/DWUNJt3/55Wa+hBWNvERT27Die1nHuE2FBTKkTmg+NT7t6LJGYANOacS4DgN
xLxmk8RQarPPapHRSTFF9c0aOMa/9rNZLrxYhjqyhBh2Fqiqg8cjS1TgfMOCA/TWBCt8R1qrfLqr
y/KzAH4tH4d0U4Fa6IZOsc0A/ngPtoeyokOMFTbSV6Ha7bom5ai3BN40dkeW6/t4jyq79/kvc6Oz
ocs55FFx1AxsgTcfAmTvjRBhinLrSBHRWsevmtd84saIM/XEYjH1Jkz7+O4t2aUp+UDjtFjVl9G8
x3xadCPywHlQWnOdbiN+DJRh+MZfcsd02X8eb0ci+Tih/AaA9fDBH0Oa4nlxeC8RIqhQZ5MOkoZZ
KNnMYa481koWGAM+f6l636FExy6mhGRx3+mjRcuH87m6GU0hVCU62QQgaTDVUJK4wF2GGwXnjApU
+Bp+2JHHA2FycZShRlUu488JxTs6h5MRJNL6LlZYQwiLLbmet3eNt8WTukwbYgIZL91MSrjwR98H
CthKrWBrbJdtvcziPzH2tOxiHTH1R62xiRqlAotGe6L/pkeqmN+pdGCNO2UYECQZedArjIypp8Rz
918tThPG5vBPtm0mDhI4MCzSTMxr8UgT9XUA0MNC0NYW/sNHHC1bciHnPJWAbIS2WXW8PRnoodeE
1m7uzB9388nVaoZT47HdgpS/rFvDpTEAsCzk/iyBaS8Iah4ninwjFKdk6Z/qWmE12glKjP3T3l17
f0drErJRik+jwmY1YP5rLWqjRA7FvGFVtCF9GmpmjUWzVaJg4rgZ/s4y/EQzFQ4Xfi7Kb60/X9xU
M9KM5yc2fzSoAgUCd6B0vAz3VIoUzvElKoJYWCONbXf6zsYRfcZbRvuw/Cx6BT7BfkBgGMEOfB8q
wq188r68mPILRmYHRewHnCLgsozQ87VA5NDZEgMASNvNBrQ8ou4vG7QPBoUDyy8TLH2aikstY0YC
tjc2lxAKGR7Sr6yYM1Uk8ZE+E+PRJ62vCuvKqLuQhtHo3sFvLZknjDtg893qiusnYKp4K4iv6uTP
/gI7Hf0gGNRK1Xz2ZQQRtx0nsSc3ANMvMEYUwKOLAQK+jVT4NS5QPGa/PoVPL4ceCG9bwpWyabGd
wHODb5GfO8boLCEg9JOQTVkhmHpRR50ZLFVZqWbRDP9SphwTrG4LAW0CaJSn59hQNKGvdDX6qVYH
9zTWCFv3ks/lZHpskuaBm+YQPa58aBV++YRuZjuVAWFBnk30sTHmEFOTLi1LIUvQY/a1glTKh1Qt
NTJNLmy6F3YEvr9ictECOplsEWQscjOrLmkuxln/6ztkPu3N1Yar7m3S0J6K36yqou1O9l6yFHTr
Z3/T+5O3u6OVQIvkWp/k3nUpUSJif3sU6uT85+/lE6WLHdOx1lq4HE9Q4Pj3F4gI8o0AKB6YKW4S
UgUTgjVZfLNRplhrJaAxC6ADqe2YnwX7NafwEITQp1C8X+bKMgiSq1qwseXzizQX+P4TrVTtfQCv
Zc3wYPlYL+jyaEeTbTNwWtJoWql3ovrsnzser15Nr8r05y9YIkfaYjKJW6KIpMy4xxG7XvL60+JD
vA7kkXrPH9qhLKKmtX+AF3Tj6EjasQZdc4qgsVYVO55FSJQhV9+IINswhhjpvXnOaniCVTp+/1Wf
+R43t+zfAnDvzygHqi79xmp5DrpEq98iIU0lw7Z/emFB/XfybImXHC+gWgEmoXhl3HJE4Py1BwHP
BYul3gfVXhGxAvfnbIefB4M6T/0IrSzGr8Cedwrw8KnXGtjfaLFjSIKlDyGavc9Qh9t+hMmSI8KX
RUHbQTBO1NXN8U7Vvjtn7F+HxUvjyOy64ahWIVnn8Fr5Op6Xn5W+uuh6WyZTrovAjUuNiaqXDxAT
aXbI72gudrAVkXUSN+5I71rlSbunW73+vP1T4vwsOFSBXOQlOF+k6+nK8YT9+JbCYu3EhscaNPSv
nD1IbgC2UjWedRUpsuOHrliXSbOGwOw0M3RPNB/W1x6hZs+xUprgrSG0Nh2rHttV6Ey1oTsw5WCO
mzDQ4we2gkSXE55VDGK6crNAsCqBWBiP+ZKFZGYl76NdkUubEZ0V57sq85QPbdNrqeqFw1PlFGeo
RNa8Z5wKCK2EjYcKwXKj6PxA5Xj0O6MrW+Q5zIpuCIKCq7cpmzVi/SijKBvr9ZbqrvnKeblwMDl7
QspFyWGoINrtk95G+ui8U9yEivA9TvaD8RG8O5Ig9lfsELLwYdBDM8WjFF4HgdRxpA5hqZczOFZC
y0XeI5f855m+2WyEGkvj8QCL6XtVJ01HfYxhfktai4YR8szNf7avQjjWJhURwdd3AHuHkh8mPLIJ
8Wk4lOmkpE96GpUGPQolQyqUaHEI/kY+m8vQ/MT23Agjl02XWb2oP1hfXCyM2k7SkAeh/XQ3IRp6
0CY0wT3quqZUAi0kA9GZzO4HPa1MK7nofpKJW5sQ5cImvgcISPDIppJCLNBUYdfHm6+4QrPJdNzp
juCqbKra6vDakwUoNj53BHFieJubm7ERXa/q/mYEZdctO/6mqz1JgsMw4NxSB/jrXV5jhipXozMu
qXaNw9eg8eToV6AGXkockb8djw+6BGJeT1YieNONalccC5a2V5AdCOUTOOY1D31Ek0EHBdwjqHRp
i7gvu4JDHgkrNJpuHcj9y/0XxR5zQRS6qtelZjbB9+rNKiLq3Cj7mQfB86x032XGKnJCLQKW7KBH
D7hIKnZyy+f5Zj2qi86t4dNMyf3AEf24ZwDEg218Pgwg4MqPKhVLhrJLnzuONjn+mx/VqL4ZVhbK
+fBcU3tO0UIWoVU6ZsZtnoAE8qAoGUfdtGNEUTfpSF51D3wbZys8KeCMtmUyzZtHo/7V5Ucq26/L
e03NefbTr3Y+1Sj7DE+hCK8t0JDX6C7UHjPaATD9tYx1MhSwi7///O969MZAL+YVYK5G/tSKRSVx
lO1jbgsiraAN9sAmtO/xfPRSZL+0QANIEuDpMlefwwXNcm7VTEbUNHEVfJTPj6nvEhJC7lSP9wwU
uCrJ6uSTikgjEY1hTAuIkMxm0dwRf3GEcOZHtxfaBwpnN/OiorkOQ5osJOFcLNUnEN89MQOY7E8G
5pGP6jJKAhYvzKOHsaIk0T92USHFODal7/GQi/C+QqMpUT3kL6d9qqd9M9ysSesBlglN95ifukjW
zZHR/pGBw08wuYnROfrY53X2B5+irqB5LPhmFgWDfhvJcF31VoJRTcUPzTKQ9lje9/NKuiDD8jn8
bgif9d8OsFkgLFkO7Qmxqd5oaCJil2gRU9xCp1F+jUCfVJ3RCh5iaWexOzdmlPHE6UqDUjWwv35W
k8YVxgwhyGxJ49l+W3tZ8+04fLv2UwT68eDLHEyteRqq2JOhmsG25Bxgri41ib+g5el6E8yel6yh
Ltk6mEGmrdUubxCTVTMrz+j7W2msMzc7GfVGpW72Ihza8fBSeNEA3fJcq9xxoocXMdLzlhvidZLE
pfLRQ83tNRBMudtoGG0R2adXd0vcL9RvD4Pt7FfGLFddwZByTOkXeqDZLN/GIMVF/mjj1pgGHRE3
tZDI1Q2kRZwLL6OVpDa8zMJfx/leBuzXwgJ7PKCRf6moNxopR0qUre2C6Q/AdtpKF/DNCOIKK8Z+
qwzBojy954nnfddJjEV4Ovy3CILFeweDwvK073aa0GxeyU7hGz6OrFDKgor4u6xAzuWXBd/Nm6ZI
Jjyd4iR7dCTv4v/qpTa7GonPXuYclwJjnioQ2hz80AUO3Yb6FYYoHfIPtUbXAaiB+Nyv+TqEKQjZ
UodAaiuKnlFqqUiTyog6mzkuGrQrV4Fpl/ugKfmguiP4AUGPaxhhZDnSdTl56AUo2jA7vj/D7g05
bYck2aAzw9mgP4MiETMBD35VloudgCx/nn71ReSJWedaRmH4vB1wW8zwiUZtwnDkdZgpRE372yVf
SNt+OSJc/BWDN+YE2lG6yuPycbwJqI+PEbjK/BFcORR1MZQemzMqfPq5uGBbiLrZTfOpI4COF4fq
ClIYYWazQfnT08HK0t67xbtQDwaiCR9xdYO/m5B7dcOukPJLljTD8VC6JepxF9s/gQhsWlBG+tbc
6KUz2LZdSLnvGpTlkGir4c9M86zmvqZ55lpsjUI1HGkc4+y5364y2E1mKFJihn5EbGUetP9TIXwk
ZvxJOcfkfgFKwt66oe//m++uAMhUC9IKXiCcP76CrqSLhyV/SNKKyCxrTuvQkiAMZx+XrJO26Fd7
dynOj3jhdGvuEvFxnJCZG480meDxFQR5zV/SInWalXAt9k8ATubPT6LMITgaQQdU1+Apd8aTXp8U
VQZ+3lWTtMKg7l09BT7yxDSFLTmAnUoaU9iWLhZU8AvuRGFq89TXB3MEUXwFvruEgnFzHqCVYYS4
Ny5a69FBK13rYZN78qfKGSTj00aXJTG16Ot91o9L2FEd/uWaomilE3q+5gdQawMGhZAAE+mfumAF
DGPBPMIw16PdwD/ZWgWIF6Vwp68O/f79+L+kzn/4RIjIMXSsvkUR1eSiLefghmSHKYhtfYFDQSiY
EUN5teeVswUhuoikwgUPsIyrn9AOTIVHRl3ySk+LXtVhTOTq06SXlWPhmR5XfJmQ41yce66xlABz
wWyPiQ1CPIp1uXgnOENzqIpZXgNK67cEuhxvjcktzTmPQFm0doxJMIVprRUEmCBlS4HKefXGhMf+
cfabjE1GaIF0nGaugHsC0dPJ76NVrPyW2MRMlujBW37PWcXm+eSrd+BtdsbafZSpjFxi2Mxvpaya
RP7I1tenIHTTRBQSaiRHKhj9asmbQFq2F6EHoydrkvEDF1lTohc+ihosBqG6UC9SEAvPpgLivBDR
Vgd+HExOByjGQaKDTosLsBfcHfYG/TaTF2PjqmS7nbQDVnlo5/xqBKxchd2C0r+GSGA8TMDYaqpa
yrS37wFbAyW/CpRhiEKa9ckCAohBIHROUq9NqCTNoQ/KH0Sod9IbPshZxFN/oUs3og1FZIQXEh/Y
VF7NVT4IMzgisMIQnewD67eOYSShGNWxwLPwqBYFY57ESXb4vXaWcsYBI1hVlUpYL/PQVm4v8dyx
eO5siVdfEzYcQxDktybUHesz8lW4sUqcelDWO7Im2W9+QUb1BBrSznZVTZ5XrCnEAhKTG2OZ3CxO
X2+qJnTgITrAbRvxNoykuaXRwR8j441lHSoQA7ShLBWoVI09BJYcT14ErM6d9VkZWzwcP3gq0nhY
xPqh9Vh3/807VWMmHRLwsNfx3HT+7Mwg1IkKwXsYZjXgeGG82/aKI6oMb08SNlE45I9/8Im6/I0u
Xlpz58E4T8Mi5KMoxAfzWl4+X2rCWaAHpXGNllOETQImipspTMTP/OsytmM9lKLwyLyy9p5HHppU
70cNAcF4YUU/xzDx7KOEMhRCsVrwlAB/mNk+s9HA5UVGSc/+bH3AY672dDVCU8tYKpRoE7wVC29R
hfroxuSyBpzMDvzlWmhWRtbhhgWs21QtaCcAgf/XKr3Ft5RXG8olG+tgxPQsqrYbn+vuaTMKm1w/
zB8h1JZSrj3Yw/Gf1WHeTvG1emyWSX/mONEJIDcV8gH/GGDbUDLaty4oOp0kWaej74WeSXMwkRak
/nxQ9WW+BgW+r7r9LLL+tqh3gVDQfaKauYtIJ93cE8RC8RxN05Tnkop81CScAR52SdF7g+1+z6gx
AB8t3U9QqN9Ad3B2h8mmL9v4fQWt+wLQPgRe0ZXbeP8qDaAp53Mas1ory3obNf9XRM/9+jUi896y
vGyMNxSnOM0wSkrlRcwLZwz1r8miATU7D/JLE64MCRmNZubTzDFdNi5v6ToTkRpRff4HC/HzteHd
krmdivbLLFfQyxqzaFcQjdVwCA5cdBtbV8uOHZ4ny8Z59m7fsxJ3ppLMwZ4Dy3cEBuSxvCQQVryH
to7C4YUFVdxcZPBpbM+nlHqgZF+LD4aXuAqY/d45bPZvZm9bLcQLekzrpHzEnHn658K4/5bs+PCb
DCFkGSG2wj010iWiWEjWRhPk3PN7hqQsg9baAQiDWF24O3lOa4I6ymu3tuioWCDAohlBoWn6/PR1
dalPJRMfGmvnBQ6sY4+YR+8U4IPKm/S22BFir58pYb9n2LuJ5Frc3Lw1M7WnQcVfsVkOSlOQiPbA
M4y4+sPjnBnYMLV0Dwr5o6qsypHpL6OVqGlyjQGKvwv280n6v1EuUbFbJHaZCbILMmYd4F6NlYMo
b+J+JB5xXPETOYaqI57jB4FOTm1DolIIKJwVi85nahLukejNtuTh4MT6InAtNmUjxnJdCgf8VPQd
munlSB4+R1lDCiy0zY88Gbk3R/P2OeIyych50RsBmkwGf01ZQvrk44kCmhj5kpOlgKTE75lkqXf9
9SAqD7c4OsMXD4kFjSTtesFNVkH2FN0LMA411c1hw9FhEh8jA4fStasIKfxiJEOAmWV8/aOK4qlx
5y+dXDKE28oXXgmpcYNpoDIVpbABH1eQllXVmkHHehplPLx78FquS8yMsNnqyyanfAaAGCszb+aI
zvCYxSPKIrtWnFV5K9kVvPGIo8u4J0m1OwHySLJFnLyJOWvb+jw/UtrgvnPECwMCLiDrJtEfACsW
HYFWRJONV6m0t7QCYax0pWtaRpa8DGGJEkmJWVpXs2Y2LYgQ5Xdrf81uKK3ZLU5zSNvGEzBhjZYm
0Ge2klyMzHwFQ3gmdybz6zfacYrHJbdepP38I7qihI8di2s+nA3hJkguxWDQGNG1hlKuqgYG/Ko7
2RReRZsbB/MmvAsrjKLqvajBnmV8vkXa5pJKohflC1rXRQtD+++tKGK8Gn5+yGPbCk3nkoqCZr5y
iUWNuQgvIaSkb+Pj/whPcBqSCfNHJTS66hXqNAxgUh0gJdh4RogfheM98II8i68Sn7yXvaIPJ28v
hcsfD8cofUdBB8jQYr+1c1UOV2JJJLS2B5UmFhLTyeMYKbiXRafdLoPCKl3LIGrx+132GiXGAR6o
Xji7/uDihPp/6EM0DnOY/AQINwrxPEKmUIpsLRhcXCqRUOs0W5i624VDzkt7kPJpNNBOWSXpvv/N
MLsiL/X8cZvRWhLrm6mB3WcMIopcPalt8+fHqdLPZb+ZRi5Pa9UxgOmtV+Ks5pWMVOEvKO9LEe6/
2DoY9JBwIzCJEaEXe3GndKPCFIfPEa54DxJLkGsKbzXBmunSTQlMvyGzH9Fj9iDbO5lO0eYzBe0v
fjkT3kGqzNo+G5ISup+CB16synrs39vgvvhelAhM3ifbKJRwff3M2i3BpfGpaPyuAYt5H0+X0xDH
C4IBBhka+wqubdGcXhLSNmwUlRawCIx61VviN1tgVnW5p1L8EhesyO+JazbKv/fMjE+eWVkY+4AN
u1OMUL8RZBid0ryGK/5osjeasU2osZQpvkoi52L960vD/T5A8wolUIUOYP2H7tUVYcO2oQXsjU8Q
w6gNmn6Q7fW6wbdihF4dSMs2jcGZM4uQTESoujUX6mhgf2upThuimIjO27iPkQVMhMtI1emIQ76X
fKCiHEtGLAxiv3kIiS1yi2RR+RUfsVq7bU6myYM9SISb7Z9rgXgekobuCREt3qld8nmMJrdVYfSr
qBk/bBWvu7htKLWmrnDmBiQbHg3efYNWIDzNU4Wf0Lk89Po+Wv+SySDFb2g1S16A7aLHD+a6xAUq
b2Vcip0J5dsl3MnLT8ow+IBXTshIbnJ7l+7C2ytGo6SpG4h0mg4eNe62DiPBGvHnIucSW/Ae0sST
v/htHLs1PtP0Ly39uej2zFiuneE7ULc6B/9VKw4O1pjtPhLWSl1uxaVHGKMzCN33P4NPUcqVgBTA
bENRC7EkLsJoFSrw1oGfSuha2zQWuyukK7pQx1z/3FATwT5n8dfI2OKmL8/RQkWg5rpfDAuaa/r/
u6RjbpV5nz5bGgL2zqObO/6ePM/365s5oT6POGY05JZapU76oi2/4cVOHTob7kQOqZpQ7RHXu40N
QjVFtqXqB6fjbNjBx2r4mI5ZnkrnChLo0Vb7A2S/978w6LaRr8sFrhnd1goEwAPllrSyX1mfLr9k
OS+DjcvhR7LcyMCrgXswMwE6W8Z2csQzAj3CHioRMC3oJz6roxoqs5ABdngBWXu6Zm7mlBKu9Pmn
8FogtN+xU6u/YZmGLHZShPu++mV0om9/N5/qDqc1eZDhZnzzLV6ipaawq1LtkYLkukxFsmkJsJ/J
/XdCZQHkNEc821tQQBAylfhjg79PckDBSYIdMw+sfyI0KJtkEmZwTRXQlLJnD176BM9PS0VwWWgw
A7SKlwiEJzqNb60a15jZKN1ikOjrvJ75CHuUUIajlzovsz2exl0PFQAKbAu+hNSw/XkAulPRE83d
ZAZWg9z4J8UKEKj2T3xXBioake38b1JQH9KZb6ul/XfjlXhhAYvYDUYxL1GaRZ/mb43ZznXb2uBJ
UNc+PTS7HQcKlPGnFmi3fpBMFh/nSjIp2ukUPQxU5e+b3Mop7CRdWQFSaN6zrFTGPvx8LHU55yDD
TGzjjF/vYF/nCVaJCx560Gu0sBoaj4WSxd86mcx5lOYx7owbeI0XRpiBBkU6Wwg+/+IGj3ryd7DE
rPEixIaOVW0uBXW8I7FlMob7en7XIxthVIqIexhNrFMWskzXCdusQcO74bJWFbAC2L8WKGaMJcuJ
HChghz1dRQw3jXbOhlx1sp84/j/SN47sKADfPqI0pETwsWHcrYh0l1B+aisvvu+xFmejn5A8Cn0T
2qX1SyGvwdKUf5kKQRZapq1b1Taj53KWRyAZCaShh5wKh3lJXzVM0CFJtzjhnotutNILFbgFf4Hn
iFp8+XiNY1oakdjCFxhi/fxWDtkk/q9QyrW2McpeKO7v89FH8bERnQqx1mcTkVhWuPOet+t4yb1z
uwmEzvFedU0iZwcaBARO36CakTyId1u42W58IEgG01ZmSEiFUzXJpCORfoPZk2RbFFdQA5RpYM28
sm/11dYq5qS1MGVa0jOx/moBU1bt+3afCXaGgB+NneKEd0jYAEvxJxmRHNPz4hn1AecpFeoT2WDL
BG7GjANyviHZCEcBpCInhuxm+SwuqCgPW29UJTQnbVghilARP49PvjFJkPB/+GbM7RR+Yj543yYi
U882UQnHgm6+uMKotQ51NmhbtgtDvG5BnsuYN/JBWMu+5DhCS2oyoyEW8RR7YIm6YTpnnAbDMEk2
cd7B2GEPozlKu44WbJL7ado/7RL0H+zX26hYUw4sPmf5N303oKMQ7etztcOw2Cs57LzMU2e9ncuT
ZBbMTGJwZDuF2vK9OfAWgELf+ECqJem88U/aL94QBvqdhPJXRLNFcicsWxqi0dIeoCau+lcdo70l
CzlVOLBV/FKQfyVq8XiaovB7hGe9MmGXea4ZDkPv0jB5uWojKk8eCW8jwoBYPy3N6H9v/4RaGRdS
qTmuGhUkwIVON9KwIWVGMIGOIyP+PFNJ5gtgnFxGB7ylmmAqKK0xcKm+KBT8NrARDXJRN8OjxyAj
h2qqWPbAfYmHDfsQuB1R2isvXc8TuyMU42FgCSm99e0x1a4admf8j4ezSqbLJ2QNogocqOqoFoor
ghvieGfzT29kq26amkN0XsxrhseWbrUXgj5YjQFr1JD+GScUJl44jd4m0i5sUDeKlxkUqI46uJRn
1lt9iveLhRN6+u7wmU1Ti1GHtytXh4xfIfNRYDoZ5L68mOJ2o2AGBizJk3HT29n0AITUBKFnrKRQ
dyIi4IgvDckRAFznf8McI+IHCU3iXzWB2zSd58g8c8o84XCrMke0SmdFaxQ6COuxnekaP8aiGqtx
kayOqCuMzL9AzMxxm7kNZ5xq30P4/UkLiz4hPXtFItszK4E430Ga27ToES41cMTIrSvhRE4gAYBN
c4J+2oICOZPlAycWusvLmfNFFNIx39WStLjW4emU6HTANSDyVQpM1K7uWVqqwNivMOkzcqfFEhgQ
TMKLbDdX9tUc4xb1BwvNrL/U/ViVKFpAHgQ7LX8PO8UBula0RyiU2vsP4HXyUIz7FzK0nY2ky7eU
vYH+71BJzgzZb2Y9wtngWvYQuHVihTeSvosDu10Nsh0DOe7GmkM/Lj7/E4a8k5GfSC333WwMZ4fl
OxhSZYMDtJsK48LYY8ZcyTFRoQu7oYF4CpQbO2neHFI9bR/ljNZ17aJi/hZ2qgMMORaavz8fOyCK
bL5nQTfnN/00d2zo16E2as+cYnn0cEZrDlxeHBfjyX6IMUAeRIcJOUo8oZ8UPXIktuDXfi2lDyXH
KscF0VZOBnOnNeSvoQbrrgwKCA6+1n+Ujl04HHh9Xmx9ShYeegfejXZDKyiiDAdUXYEoT1GnZukZ
ClOCnDuzFk2eYWsy9z4OjcX4zgGEyADyatmP3ThV+9lLGW3h0v6vzheXtgr78H9G6hbOm3RQQ/SQ
yRuI/DMY10qr4aHAtupUboAMJLG7nanrN7TEmtSIrSrOVw+g9ZCgridB9a/dXC8HQfMvmaAVztM9
s9rIrZD0l9zchz5HB3Wr9SF8PqNsQeZBoNoFizY1tO7XwR6UGbzafc5tQok+Vl0mOXDxyFG720/u
zodS6nhOqLjbhoTDikMsSclx1XNlMwGE5Dc0nuy5+UurbJ9Sotc8T7HsuO7Ld3YCeiFZSSmagj6n
9a15lA7wYnjkFa4vD4xlti6h4k5W5PmDwOGtvt/W6q8JYcFH18+7Dowa6tHmMyTWWtktRi0fk+lf
ToXQiKChF5sm3cnDs6/IOEvy5PxsUlY0M7fPeTqYY7x6j1r59vWTbR88bpv1mThUqRL2+rS9JFG4
DMG2jTAvmrqizH45M0Ry+5gnjKKH0WF9xocUylc5Ky6/3ta8IwSc9Zx61q/sr9t9xbQwV0Q+Py/g
M+ySvBcU2EaIX3HwKZcJ4EcDvYusiP3PtPdsEwkjPyExEXl6qCQh7mqMYZd/VuxKK4jaIHZL7sa0
/yOZJfvv2n2F2EfEYi156Cw0C7DyM58zFZ4YWi1/hPFAO4V471kjdlUG4ojh8WT+0X4dp+6n+qCd
HWCD78a6v/BPFj+U9A0LFA9zao2Rk5m5dSB/gdwxgRX/b9Tn2OLt+OkaPs+pbJ66FG9Ov6DrQjL4
VyoEhF5yM530t/cxLhV3NMBTVd1SV288CsHQEe5TD/HRiDRbhxauHJi5Llab+6no8EuiSbk/rrOE
piv/2QigiLa9LoAVp2wpEeuiebFfAiE7losv5oUDaRT8c7BL8haBOyHlRDqvpvoDijpdjLPrZ6aI
tOiI/Xk/n7LhXHrSbvnEIrQyB5E3H0b27PsBvx0ZxmqtdA6Re7pwBqLCkJ2ln6E9ww0hvSkzZQxs
HJU3flBAkvIZMwc8pjD3BrARmO+4MQNGwaZcEew9b8YtECUXJ0hjIX9V2Rw0D6a+xTddKqxa3r8H
HBQe3CaaXnjE0n2pjgWzBkWPFSfAo5R11r/Xi3yBgGtUM72zc4clcfZ4e5XfQtUyqjW6GDtppcKP
PV/ND+1bk8C8GWkizD31VkpCw17/GYGHMDUx0mOl8s/OW3voNRPPiCVZ3XI76X7ps2xYbFUGxBSV
NY54D6XVPxq/RND2xvy+CyQrWIFbK8EcQvTGw0f5k3zDYxcamEZzDToRnTvOa0+pImMmaZGO/zZV
G94NXpLEuZnOqtkaaAy1aFXt/wd7RiPIXhiGaGNyp0I7hPfN+cxcBxbMR/3vEnzm4eJqYi2TtEBb
H7kQYTWPvhVoMKa7BKP6TGRvP6E5iYUMJsiyVGBB7tbThQ3ViBePpk+eL+CwbAxVCyQY3RDvy+M/
HK69bKcl8AfajIbuJl2Nwye6ZUcc4Gls6/56E0SWAWByL+7uqKJkH8f8Q/+5oGc0pTW7oTtqG4Be
dyQVPjw9E4JdagCNRdVWp8DkhvU6HPzMQeR2xaaBgv4qPg7HjVbclSuWIC3tsh0rpYPTU46IRflU
fim8CNyTxaaWL7P0BVv1N2uAPoBYYdoZbcOQ6DTY+EjXZbBpDW6gwrGisnF2jn+Qk2S5GlQyRUWW
bm3NJP9DJ+ripPg0HwO9dJHKYmvbOn/0jjpLpiBmpY+s2c1qxly107PUI6ikf/W5wiw72vpFzvjZ
JrrRiXk33FZ8/M3vKubx+gTLKKZScPQaIOG+ZbnQW+ZWjSejLanO1jl7+uYFbRpSOoPGp02qp0N2
SM1XCtwbqIlILadB+kPboJwoRyGEJFk6ylI5e6B3AIMMtnc+m3FqfdaI6uxoOVVQlRyJbtTveK13
byfwE0MWmwSyjxR1kMSiiR/tjsiRt7Y94AtRKyvVVM6T9pWG4iV2urNaBHoSllxOgKyu+vJShV9R
L+Ls59XPXn2kp0VG987xS8t3T1rFfq3qknldKmpBcTM4gy81Aehmd2a5YhRzv/D6Ej/Gm808y0vj
EfKAH5Bi/jjAAYlO6uY70Zyk+CWHr+XBPuAMySi833sz9Dd5XIza/p4oS3adCgCrbj1qVHaCxP+2
VaTvowk3JGIA5ghtTcZ3TzpnCfwihgjDDGmCYoed/OvD/0ris9ONK5PBD7UOvBTMXJNXZv+FhPRx
ccxP4BN8eMJ3d9jFkMSTZvQoEWSf3rqCz4v1E/ohjldld6sjbJ4HGw0xu2KrHlU8mf67oqnzfRsH
qYUl7lUOE4SP6EWmzVV3qeXtVjyL5o31axLu8rKIuks9NxwUBsy066h/rGDOJ7Yn7mZ5iLp8v5NQ
XWQDuXh1aBOH2D6X/7tvTbcteb6XH38gWjeiFBG8Fh629rOjPT/IM3ZepnU6YxMaXB7lCDktub+P
wL8oXFyZi8rFugYaB9JyFklx9DPV33Xm536BK3EibYHE1drLWEV/DfeYterXicAKrrwtJZ8hWFU6
TZZxv6DVZ4CW2kBqEhT0OO5oiEz4vF1xxhYYttBkEskY1NFDX6i3d7UoOh5MBBNug5adp1YLkYrc
fpTGuliz9o4AvgCcePqf4OdGvdJR41cZsKAxK9ytqaXi87uvuskE+eHJvg9AT+SDy/HDPjn2mgZi
ZtreDfiK6oYSPfuOY/wMFcWrnyAoo5B8GEsd91lA/sEd+b1Q1tXxgM+1Ler3WBWLzyO1XvYRueLI
wfyv3vSaSDc5C+Ufhx96SkI7lRo8BzxvMEk8jg18Q8Edc/3cnB9Pm2W5TwgNlj6OmWoaPaj/mn5u
DFHwC6DtUHiQgH6tUqBFswEQsoetYsWE1JPKa7H3nAgZ4xG0Ldm4CP86ESZxGm4WoYq5ZW/psk4p
y1hZHCz/1XWtcMXt4RmBGU18pljJbzkKSQ0Fv+qs9t6ozgekG1bpIduBU1r55d5jXr+cju++oC55
VfLsGsWMjWBhaZOLo7LlZ7h7VqY0SD26/yzq6n47ZnjntmiVgSb3gZFHT3ziF0t8Cu9nGLLGRz6E
lMKUcCJVVOFBAeAaHgatIx0e7pNbpbhHRyUwSiWWLfDa8kPL+/xjAFfCFIQXenpInhdf27MsJ/c4
jdexXEW7ROrrRI8Ly8d0e+GQjgjCpLtKo+4hr5yNPNGiTx1ggrpRidUjdkvPm5PyfIcY7rXRFz9U
DqR/gdpr7WQVaSU7zT9A2L1kFFXS44uM9HDLjbiUCVPWYqFBVwOYdT0wRJVgEQjYD0W7/ZVDCEG+
lPRvD4Pk/0sSwLATW/9x8YWCeuNS0+3s5iMPPGdyuoaSsjRQCUL+GTFkCwJ0PlHZBLfw5G32Arnn
dTZy6rkMaVoTCOncFrJ/XwX1qhhLQ3caseSEaYNLrDaSLRusOvKcKZ3sZFoqhZNwkI/IawE1FaLq
jXCXrEyrmHh3lnL7j6Rl3ZFtM2/sZMbkKHElD+AR7HXDikvRJIvaN6VmlrY6OgEIyAKfAsZNzW1X
837sMuireQjrLaRqEWZ3+/Aq2jP0oxyBJUBk/c4kJFp/TVBhY8mbs0zUQdFzlWHUDafZWl1kBNWv
Za1KK3Xc0XQOlc54MdPwnev5laNFZB7UchkfbDwHverywGir1E9bcc+zB8azzIOVouO/gunnEHcS
zZcvhPe7l21YuBkLbLVua9L9mtz22rtz5VdOIsOElaurVn2Vig7Y5NaViAcGR2HZXVqBR+2uO0dw
ossuUCjKEl3hZ6LM8WuJnXPzVmPjaXrrhS+7EYt8Frx3jxedmDTx6/XXUaC8FYSR37z9G228HJcS
Mf2o6I3CnCl//CcAJ96b+cH+bOxnBTzyHe95CEl8pc3zw9aTQJc+blabS6HcauHguX7utUYtV6cd
SgMgPT3kzcvcIrzgNtaIKImVa3R4pU+Mtf5PN3B4uhloCLWyYlFrG323cJFJpHj25bMcuvbob2q0
q+RidNNmj1JCCfPBF0Ml2Jj6CctK30t61UxIVKWMZAIcAOpY7epHdyzsqnUwaxfB3VQ3K4uulZHV
HcgFzKJmI30HTHBGJmByTBuO6rQBw0utsY+pEgWcvZWmbKD/gHY84S0J6XmTAg90NGmIZV5RzMf9
1snsiwNigjhMIypjoaS4RbNF5soBkcjOxT9YlauRt0V3IjNl84rKNqTXTI+BwGioty+lu9rPJ6gT
eHSAxeLqkZ1hsqLXFOkn+eUdEKt9Jkhv/5vXRP99l+eZTrPFSSUZfMmxP9MQGCcFETAGDZ7agNmM
XaGTDiQtBa/44nn0EfGXmZSTPojhTTHtzDBvWF9kyms4PRUMJdzHs7VUoZ0qXodbMDcMUHN1FLLD
MLTY+zT/LQc9EneI7ll32W66X/hu1AyKFREJn0stJoKo07BMnsz2sZ3+waoVSe59N/Xx0mgwX3q1
5KFvZQOjDQLEZaxtP0O1C28Qz11AIyp1Y4Uhmo0+jRwoUygXMJrM9BkKS3ASus6daA6m+UG5XlZG
m3UOYtil6vL5uvdHgJFGf0cJeOzxHPZL2WlIdG0oIVp4QDNYgR1TKBTCzU0PaVayai/n9kHvR+HD
VTGNVc72UkhvJcJmU9vJH8/E9DR8Wjroi/j1h11QcUAkO9U8ucSo1CPjpcc4RjQNkT08gOApSgux
uARVLVxsZD54woAJd634IrRXgS/4sGJ4LHCxTB9w/3BGOiG5jvg5q8uNmyb6MdYondQPizjH9tSc
kxDkb94Y+WOFEJFNQzP7ArYmomeNHHCvkcgUcvqhFOHHGF0YieQ1ymkJ986q5t5DIM2DgY7LEFAv
y+t/7nwsRvJzKB+sG28zXlFU/D8hRsG/4AIHgnrpmZPmdhIdzFbidZWMx+mqUnSkLDXSrKA+20qD
Fggt+VCmZrb3xP5cJpEVRXWWg1oHU+WVAd2wxBTp7Epk3aejm0OvUSUktIDHUk2If2l8Kt/6M0Vf
KPF8RIjyeUkZ6Awk1KHrySufh/ZPtMzcY7xaEb4zI1XtVxDG05ZaparyxG/4PWXwh/g4YZXs+VRX
7Or9fhly+N9AImSe70qb2L6A8+tsKDfZGedHYDOx+Pg4b7YbBhJZRZhTmo6v4PeZebOi6gjNB6w5
yWNNb8NjAVydWu/EKnagHBJ1arevicD4YGMNOhinr5I79VBLN2eR0jSOL32BWkAgRQY1VnI7av5+
F1FJJ3scfof+b8ft8YruYzA5BlJ/YGLyw1o5pXvyp/wjDNavEEQHJzZ65FJBeyD0T2kRS1NIuLs4
aY6jh/N+UNzuqUowI6nAGIpNslvx28LvlyMTU3A0Q0K3wvlO5rck6gFRRzDDd214oJqiOhuo0GyD
pbxRYWlu4BEZkxOMFKshNLQVO5UkotDcD8w7GU7ATHNEe2k5zCovTvKUPz0HrbCLzCgz7DOn/XL1
TLTMIBwihgKwZY4xP3qipzMMdVP0KOuaaKnQxUuCiYWecaioRmHWn1WNGzkiqfa1Ayp777SjIgKG
IEZeIHkTpFuFYcjR1I+8YaZXHO4QQ43mk3eDyig1xYpu7t6xEMigNlo3drlMUFjXIhHGwVy6H5+D
HP9qdxrS7QhE6tkB4Fxn6UTlmqSp5HUUr2oFdEktPXyxIZSHQJ1neQALkjan4++/rdgUl2cCGPtd
LIYt8KpMOKTp+7n4QOpahkZLtYzAqLp55JOT05KdxHkg8uTZcZ/fQ3Qlo3zx+297B0T6hZKOVYAr
oDDupRthAB4PxqLQP+6whc+6YcEw01oOPz+IzvKusPZfeKqDVgxVchw7Fcf/7WSVHGoXdninqbsB
aRXooxpeUYMR/hGKei4lWk1BN6S5fjA8/ps7BpIou1hRIym6Efrf9G+bMjw67ik+o7RB3K6hybDv
Yb0chmNfj+jvVXo+5qijFMQ6odrtuLlXnxX4kigyr7HYf96sIO+XsZIb1sZGYIBu3jKBefRdBCqX
C135Rleqx/4ZCdzifh9A7kR49nlKUrWkPccAKfFn2px0Ce22HG+Nl96DbqpVjyWci4+B/4sJ1qj9
iPzFMR2EDuEb0iIlYKkM6ztXxpJpSxmchuwNopQWSTLLvjr+CH91J77FyVcTqHtPiJrnZL8te78p
aK9tpJHpRQBsGb4U22NjWsqWrsxESpIKb0pVLg48w9qtm4RxcRw4BeblceEwr9K1RhnZlvPT1N34
rRftJZvA/5YdMTVHa3bztktTACFVYoq//lCgSogehdLUQlThtFo9iT5rSImCnCpJ87UhN8rpvk5A
s1cWAgBM+w0Bsq1xEqfAI+LvdclrMa+aBmuCOSzn/2OrxBq4SnvZM+bRMakdVGmNQxKweiX6AHQo
DKTNKCJloEC4uZJ+WLdUET8AAZ3Ju4B8Juz+oXQTVhrzHgqQPa/W2NUadwikeA2yMXakR6CBJNMH
9lBzcBBN4M+LfTcUYdvPxHmPyeHI4k7N1KWGxw2LjHLwXoiQXseH+TpTisl/sjrXcadSyavVoiz8
LKwuxoUiAPvma9k1mCLE1dSP6UjEXFdakK15qcBbqlF8P3EbPrN8NrG2/FBEJM9QbMce/PQ6+ANV
O703hn3ej5RKYsBkSR/3s+nj4QIul3mpWn6coBOQmv+nvxA+FgaQhIhPF9VI6N9W8J2RB5qQ4fU0
rm1bW0qHsBw3uUXabZ65Z4fQBaNzr8wmViG0lToCEHqFdA1elQHpCvBswZfNDUHZ5v3tqvmTl8O+
hkStctTaU4jMLQ7BDhVZ7hkC5TqwNlwHzk5EgHLbCDJu+UE5Z2Nq78Rq9lno9ZO7Zce6IH3MTuw4
eFq7evlOylHhRlFeABrr4v3q8MjMHASczZo5mVuzNu+UpnJn0nyQFRJJH7VgK/gRPwO3J5fMotYp
4SZ+XBFrLcGTPe9fBoQp9MmBzAnCIRlfSlxjaxSluhH2VlM8gLNA01FQLNR0C/DJH77qwN7ciRDr
3a80zWWmfpT/Z/YlfniwkQJLMzMEn1Ygqnz9crKCITLWRbKjOBmkBKtSY+oBFbemsn1MgWqXODMw
5/nrd7y19/MkVDhlzcpYVwYt1r9TIAgJ9N8OsX53r8SzzbZ+zYljgvfYBM9HRXqKlsVVFTENvwGH
i5J+8wkfzTvAIsTpZ1KsSshLLWGquX64g38vtS40BLI3LcXI5lLKsghBaphrbxQrQWWJyvLPshYl
xkM2wSbCHOaASpP5SojY0DFFRN7yG3SZPa6mj2OlPC93nnZ1/xE40l/ezZx1F1AaK8NOSBe0Wkh9
1z6My5Fj5k+NDF7QbbbecliixYShDJ25Zqy4DlN4QDNxtJGekadaUIipsiv3gseakTvOzcD1qTlU
HDg393StSQOq8RSF3liApmW6EfnF+3VJu3uZTuEM6epWr68A7ePzu7ja4iQgSx/vzQdSZENlYxJY
pGFTp9eMHvJ2tegdP0Tvwm1kfbHbhDvlo1LnRDqAeqqEpaiHuzJnXgmFNwQ5Twgl739tBSO2wUXB
pwvVUqd1o2uja1G5aR8K08W1IwGEsYjpvvuplssfJ1Q+wjudLyQ6iOCEMCgmNrxRPbAfSBqaOrxU
jFBim4SHVZ3DKwvWXnDQJP6qGRJjffH5466Wa03I5D3THR7iaaTEG+K42Z9nNPVEEI+e7LSG1Do4
RPijbE6aAWZbffZUHXRGG1fquphOejnlRU7pYBVvKilhatQVb/rNcut/G2KeFCkV39ktfLYu6j19
JC0NqKzVLIPHhi1nQpxPegTeSpUXRHniquyKwqNaaAEOvWapLtEcwJ0RgKEDxkQXSCFez8CxgH2Q
limDc/vR7dCQDCgxfliiHVJHGpImWVnJmAg8cUVylK4NirMxokXj1Y+X+Twr7lP3uCWvl/y/T/RY
XZ2orLIQ57HYXGdB5512BZgOabmHtM6KHuZKxsq9higdDB5TzTHEy0vhlr5JrC6wXcMT0JtaMzEi
U5uzetUIv6Lp263qiUwyt3xbHOWpsGIwiyPzYMdFzHd6AU9A+ut3jfYCJBGx0B04Bfin8+KH2J6X
7zj0y5LMOtxlXcB/XIYH/sd55R7j8U8asDMdhG7q0WZX/Jnmz96HlP8jX2Cb+39YssijXqo1vXIR
ySpV12dwFrWIyTOll6GLgmzf73KohYdeo31QXZ+RJPVvwli//yAPD5wrX8JWwu5X3tVH38HwCq9m
asX7X3WVnqImdwMCWDtluSREY4nzpKS07tLA2OQeUwJqIIbpCtZhoWhfyo/3iS/k7z9mGZDaEqtY
OikPC8obJV+dS9t3uR1x0w4zkYw2NJsfBcv3bIAGZIyXq+4xyskMpHbGU06fb1Fi9h2SWZ4yroJz
aXQL95uaiKUeYXgkDwVhdnnH4EH7WAcbdcJRxZZT7f4TISF+sbEiaEy5k2CUi3Oj44uFB/oCR53v
IQASYLA3Cc3IwxHl2zUUhNJtOABca46qFys4kh7y1PVsqDBd4doYfeq19g3HsDkq7eVhvzrXB5om
wa1DZ73PqnNvf1D2uBxNq4vNu1Bb1JgPh2yrVwlsbrV8gBzszS1iHLg7otCThAn2xtwn/SeQzSbs
EEJS5i4Ua9BDIxywSND2iRo+IDMTBWIrAbNgSvQZBq/wINFOD7c/ffPd6sefQPYLYgW7XpxN+lfC
iX6zKRatDua56eQ2uMAgeJb52wGTh2/W+3JobOLxRY8P95u0K1IH53vAlqOikpJIT8TyE+9y/Pw7
8YO/TPPQJViciAtvW40L3VU0Xx65ePWbSmVThv8/FnlydC9AEl0Q4vy6nH0CGXJ9OOE3v3t+qcoP
+RuP43FnPLcdmN77Pl9HXm1Sr3Z6ocLle7KR/gnqZVEp/pe3payGQLtrI5mQQF+VOBoavYpXp0yC
UzuYsum4/Ozwf0Si/ZhRDDLbfy0CPioNUcDC8jYVkvcCb6mpagthL4QEkJw8fEAB2Ob+0T0uJoor
gZBpP3Orcr/B1RNA9/9F/XsUAtqw9ymAb/1A7C2sb0H0gvpAaandqKF/B5s6/CEk2dTV82yzBA5N
BXJDDWDqzgtfUnrH+UWX9jAPaaQosWfFEQg6bfapVJQd5x7i+FAafDxuGMzCrmc/UXvXyA/L617b
kwA5A1T1l4lzmIE5uwmOVNs0qZ0QH7DEienqbwJOMrJt2nK7I8rqaJzv1GB5sjSNRjMunJ8z7YG4
i7xyFzGPU6OT2fVseMLUuWow99+yT+zJbdS08MwZUt5SHFAbjxaeDLEyMa3lRBfjO3Z24KLiNo3l
l8xW4x6X33bHe/Xn+s/W2XvVjTI4t3Bf8bdlaLxl5Slud6xWpsLZpbrjSOM7ESbHyA293qt9/H1X
B1YNp16np7qYODlGm4AVN1s+0Ukpu9fB9rEsE/PHeBN4XXKnHE8DPIVkH4UYjXmROknwZTIXlK2M
UP3aOXYwbsNTQzyffv9C5zuOTp7qMN5/W9f9Z9UGwH43yiGyblLiNrOnc9l/GuguTsklzfMYNJSu
gn4hi0fzbve8nRUfy251VUVGwbzaOZuCvOTKLoaePyKTiGcsh9qOPm4XokJrnd/IDGy4NjIBDegD
lPtLHVQhUILeoYla8mkLJ7tYVES7o4ejSDAx2yd8IJef5MgY2urA95VKIBXg3OmWG9aCMJHc/Ia+
tqlUNtc7/Io4lOvWgtvPYtZOd6A2WI5xPMI6YIU+m5SbKBOMi6hxA1FKJNFSOLRjs2wYAp2UPPkM
TuDB3DM9GxdptraaAVLLb/c/QYh+d5PK9O2+o4lVT6Mx8SKoTl9TpC3iSN3SbghW2NQEO3DSL9EM
qlvq1d4LKivVygLGCkcqIwqqUAXTAbyKK5KvkL4AB9cIHUZd7GHEvDmRt32bgFUOMttTs1DaWjv8
aW6QGRxABIa464oqZOFkS7tzHkG38BJMmb6xXe/kzDfCeI3SeZ/rXVRzikxask8axlFaXZ2xW3kz
mOVmJS9mi3ChEOTOX3KEqWDfA9XbfFzRDVr8EcY9Ob3Ou1y6wUvn4HUjHWz5qKYwnqp4AypN5BAJ
qHHsRVgPR5PsEnwxWJTfR7oYh/j8WwT0NQoxnOKOBMNV1yHPE15UX0PW5ia+EO1q8sd/Jkid2aTb
dKPIRT8OONu+Nki/uaxRw/wNCXv353k+adzL5/zudDrRr/sbJxAOAovy2dI5wGKfBiousKpYj8Rf
1ROO5sIgOsu1AdOY/uID5mVsIi3K2KQf5ADxUS6GIWsc9+nonOs5PCjNoR446rcYGU/eQBEzWo0/
PXSXJrl2409zQRWYd9ueyfngpT+78XPzwT9ualNxUoV0bshWIWOKEF+3wmLkU5FvhbKWS3+vrWuw
72hrBt5mV4FiqO+o04T+S1FiFhUgPahrnp4EFabnfdrApCJqMSdkTqD4m1BhxOzccVpu4OvMcu1R
Tr37p/iRReivmF2muzLKZpTUFSIBcRZLy2jNTNVoSTgDo4a6P/vSGN//iPqi9u567ZLU0JhTwEwt
S31AHADph4Rpwe+1rqNtKhd4KigqAs+2s0hY/AdJg/I92ADHOjX5qhtV+tC5Vo6kotY2V3/6IF/B
JPLLshf+QiK7sIE4graXcfbu3WfP0ii8+th7Ael4zMrbsWy8zl7LYS4BqVtZTtFJdwaiCOCXdj/K
tn4EZS2A/CVuSiE3wJBImS3zkfHBMx6L6Tmk5+bhw7ogqFMmNJai75mh5Bv2u3Iq2tWgrv54R6Ur
kX9Lte+NTRhmiY5Fh5FqGrxklDcQn5RkiL9ua2d5s2oTRE+IE9SXuKWsxplb7GE76G8HGZ8jr8cs
p/OJWrHScq4aob7z8f3yWN0FtDUC3ppAckyVQc/7iZ5fYindn9NLxN775RkXW/ohELZnkKDnDKUf
Sk+rsSKyo5VlHAfcC0zLrSvQi4KP9yHbMCB7X6acWeV8ERnDbt5PzbtR6Y5RlS4dMzhZNTcDcL/k
/ayawPKBaBnZMzL9HoaXf7ZJFfEW/Ewn8G659mQtIeqLENHLsy4/xiTfBMUR3F0DUGlJv9W0dlSt
80yuqr4frVA9pK9IJBfjpaEUyQcpNdW7fl63j7a2TToYWKQYGoOrD3A5uBgcXIvcf9dU9wBaSVsn
Dpn7q5REWokycDTclf4vkpcFc3E1NdYjn/FdCVKwp2IV1hrBdR3umVLe4Pn7+OW7spP94wkyv8Il
Nsa4RU0U0bdXMRaG0M7wYDNTQCjpacNni6uXH6+8scwHpWjwmU7bFSdoHxaMj7XaoTsrAlvAiBbC
LqQ4JRZZXxF7qD6djUA2n4lYpGNLKgFOmk+yx9OgEbHwld/afzUdT6BScPPzzAHyf08crMnENtQS
uhuwHQ2EE9DyJMffz9xiZ3mza+TNxA3YjSTPoqUq4d0V6jfUmM5faAT5d1mbIaNaLtikdm5HzBJx
NGpBzzWuOJlD9425xgrSqbrWrjph03582H6xRJXjd9xcB6Fl+ola7KYcSvMlN8bjmgPRXkYAKH5X
y/doI19H42ptE5g+3TdaISj/DdVzqVzKr1LVg2A9OYj2TKdSQKNF7iQpwokoCtCAhglCMU7cIrUp
xhkrKW6+JkZo6gcwQzQmpKREEFF18pBGUWcvxGOBWv7ZWfahRZ6d0TSccomZDXewXHMM+A2Ps97U
nKiXcYcPxL3E1cExSY4/0SUUYDXhiduodc943LjhzeSQZAemQ8MToF1dttAWUAtszxQW9bLLVVzK
7LrZkCBS+Kg4OfzUiPMrGfEHeyEieE1+UzopMC+YsoIUp22jmGRn9NWUbfUKOCqQqZIYRIyderH5
oSo+ZVac7hGzcUyA6136FjcLrBa2fQDQQJVL6k9hQQeJH7HZYqTFXIK6iG13/wclODUXnID6lXi/
rApTJj1NZuRQwWNBKfA6u0a8Ea5CKYdi0hY79c7CwWRnmipluvzlu4xcMWL3oU2g6I1G4Njcgg/2
M5VQyIE6I/D029PiUgILCk72wYOSkHeVmn8IcX4f43enekZyK0+gqpjIxvirQYm+DpeSWwqmbNpx
iLleGJMf5aIxz4H8Hn7nYu6qzeGea1l0pKJdLRXdoQZqAH4EJgqpoxpcvws/tBdandPWW2z9t2U3
JoW0nyJhfnQ7ZW3HVC9+CR4+aVOxH4Plzt8ftHzs9yh7yaNXhr2Lu95684lvANG5AdEx6/1Z/rf+
C9HsFYHAnVb4nVC99YN4PFQrVg39OkOzb5itQm6Mn+jWSYZD5O6aak+EUVdBW3zB4jXFosgs8Prp
odUrBWVH6sc7S4C4U5ikKoVNkF67we1aVtG6Gugy/Xypmw7CZdTTsl1xaAuT4bNcwFSazSfPNyxk
Kwiu/NVBGnwAqMnxoDqMyzUTSjKt/EXYj5U14hKBYMQUeWE9YoU9OIaeIvI6WwQv2OA47zrURPMw
20NNP0DUxi4u+Wewqq6N9PZ/kyex/BQTPW7XmQAtJFcWvvR77VlOpntmI/YNBCn6opSVfZ2bjek0
a2/RYI0yBKdj/0EGLY0K0Zi3KnQyWuu6iPI6pNqX/+LrwMuQt9xqYV6uZxMH85a0GPbGC8NWFJI7
NuuAYiAwLTkneUaw3svfun4PNzQMJF5avyB7DqRuHsE/AhaqxZQD3SLGtWf/Qez9ETUJplhBP/3z
XrywEUR/aPBsj0Kc39QnMsVR5XE2FAysN9dViWq4vliM3TIXKIO8g5ePofgjM+++UdeIHdkJMf3Q
RRNaNh/AVuOK8j9fQY7hKPphuZUI2PFZxjHHpH8SSR/CvMHztHkE9J/9RdzHQATh7EWvmIVGGX6H
+R8Uo0udguQwh39dJ1uG+Q+NembRFzoMc4mIBp5APz7Xp3/G5IAZo2I6s6ak5jjdex/LTNLO2kXO
K0xmVTi8HpHaoiJmN/WyVTsImUpWXfXNfvWozgML4nWG0tkjfCDUSLtgO0wLV1T5xKGjkTABVp1R
6X2D2rn/Nvc9BDbJyNfiixeuii4wpZGQ67Ae5+bMrJATeYHwmYjqyCx0sAHFbPJX60KrPPxBdbxb
nb7dd4W5R8px8VCaLpq9AvfRwgOvXpBYHp/Li9fd5ppAzGEHIgxW9HgbSA5MZ+o7TOV5ckLLljJT
RXJYsxzuO2oPXPg7n60hf8amUQIcdczyPyQuI2CF69Rnt2CuQyWdD5vOxQmzlVzkTD9ugCdHixye
LKi6whiK9E1AyqaWnYmChJZJ2iDCE+RRos2ZyNDwNX2vhIipUsj8bTAPlsikcMmI1kuhh3/hktv9
pwR3G9jCiDRIWqpjmmNUglpsUdH86z/KGT/naVcIzA2Nu1qQaG23ND41aW/Mp9ufdc84s6bZ3tTy
1R8jAs5JWMCkWY7FvoEylcLBv9gy8Y8TXq7d3d+PuwLaItPmyLQ8yvPy+gkvRbVo4uNoQ+VrJYEX
u9DsdBqNSNS+P808SRnLWL19YWhCqfVvsAal7CIVZylXYSB5wBeiVYfbjVp+ybr+0SEGd/DjSqZY
qIr4Lq478cM3SowynoZHYifVIdnNzRHkvVWU3m35nrq1kxq7jyqRjSbizr5o1z+5jjEPPATwLbrE
/9vq870tb8hcAZ9jAnaPVagIW6uYNM9oe8Sy5XQh7/V2jxLDu3K9sy51E2NbCR9RLgqG9qNIlEuX
pBCAFcKAgWoamLc342bbbP0+gP8mZYtQYZtw7Wf3dbSiw4vE0LXH3mFr9LeVzQ0+WEbuneAf1EfR
zEDSLCO6GiiVWR6a4wqA1u+pnZRx2Hbrc9MF5IEKpqxLw06KpWfgaY9WuNiY7aYMaAVkGUjDFtR4
tcxwyB9eWWGCq1reWdkeOX1vIVuFlz8Rrgjjt45HkVM8GkPnt9NxFx3XOF5JbCB97cOKY4zwFVTz
RFQ2FXCnU4YU/m4yiSuooogyuhnSNEKMr80J6zeGpwKhZXCJm2Xf6OazOrph+QKYXdYL+JJIhM0B
4NCwPrA/0jKfim2QufLX5/n30zQsHlowGNc7tYskoOppjaIYXhwRG7zjEek+hUGN4qxX8J42+gDf
RgWz6zRBoIbzEPAwcULNY4IipEg6q8JJRms7CCT9u1RUOqZVCfAo5PJGJwgy/dW3vBdC62oFXLRH
Jl/TIcygyAiI/6+9KI83mgwm8unPWTDXSkknmGVii77hlr8rZKeQMjPsFmdzhxf8FJfcYN9RC5rM
WyEts2IQzI+TwY2tv4mxo2m2ducbAdoMpFchhxc6PCuYYZiIvfdm3SvA2Fk6UAsoU+BrPjD9Abnk
ilk8gFDaJhwJEUlAL2aeLjpXXDKgRABr7wOOtujwyh5CVjTsllgL/3HZdid+bf2EmUcbL6/Pqv0/
IZZllMPcI8pBun/HIHz0JkiCTNhqrUKaTI3IKWfc7UqbygqWVEUOPA3StHk27gX2VFPWz1MOE/gN
v14u8HHg+jf6CpFwWPyq6c0qIgr0zt1aYwbqQwyqkUbiQTjgQ0dXvJAoPBp6dJvCi6lDN1x1+ro8
iOIzCpy8sds1iQb19hEwx11UQnu2rc4tUMZvp7HAZtcCABNMJ7N+44iQbvB+Y5XD6nEAhK6RWEuL
5mO1+c0A4skpqpp5gaQtuAvB/hNd1/1QEHxbboV5jDUP8imYVeEeGSLFPhFGC4ag9keiXqOhNJgH
j/jqtg0jHx7rTcTuP/2FXebXgKHxjsN5aTf/+e4yNeGNt2j4gbBvtOKubow4x7AlFNYiBS/bDf27
du3PDPW9Qhz/X7yzR7IudlGrea+ZgW5GF8h4Gcygpjw3vsFrN9ATxdEFQzoqt2FJS9/2VpKmc77A
nz1NkNfPMIiuUqXM0EL+dNnKW2LxUgfuAT/MyDqEqoPqGZ630+IaSSih94+KKVKQQ2WBNq1RKCmy
tLfyWQYGA365QEpKeZTCvczOYeBB/RA76tE4CgK8B0E6gXsE4uysf9/Zb8J8WcwrpgE+MuV1+TIk
fB1C6jqPYAiSItZFhPSK9P+OYdOth8ImjW63Jp+OHHkDUXiEfjEGzWr0vWEujafDy/JoXFTku4Ty
BXrbOG9ADVaiNT+eWzNiPJyT/3fNqHQfk8d3W4P6nVcylsnLa4K/GAWmgz/IN89NBxx5z0ejqrFS
df2levDTqTDAGQiYCbRs5ZcwO9RycA7Q6LqF7USPyaDzpu87Wz5QJhU6UKSiAoCrUFk4ZopjLeeP
38QQD41UmMxqqEVgbKtzQ/2uwhOUaQ2UMfYPscRAmZVK1eE7BZEge/1XY6LmmjAL6gRziIJBBh7c
0RfKyy2zcvxZjZffsFUPprpyhjx7KZgw1MO6qJ2vcqvjlM8TPuWwozCO2jRtNCPxU+kFI+KJsnsh
8lx1gTlrFJmeUHW7XNo7cXYBRlDrIJc0xhW4mUGuswa75KqykqGI8y81jjcBe+BibrGtCr8jIleC
saql+sFPzaaRp6D9QeUdnOAIbsUiKxVg3uOkxJ9Jl2yBVeDKEmyt4WdH/Vhzln5d7kYDZQNE0RAy
owCGHDVuH72oYnBFbifzCA8bMFSezDEi3LxFCNgM1W90KDY9O1kVLV/cLRlxXAKSYo/OscXeiHwN
X8izCfVPxriQno5KBVzdtdKaytjVsx2sI0IwkZSgDsfSNjG3ULZL1vndLdTKOUW625fp8zbT+qB+
kZs2sxVm0S4rByol+lnHYM5iRoAWtaOeHwixnea836YGQfy8dA2Wqdcv/lqE/Uhn6FHssmXsC27v
AgVqRXQVni35ureDZ/9Vje20Ug22HMZN2hupidg4IbTj7c4TGOi3BDIPm7CM8dIFMMwo9Jxuo//c
27dW4hAJ4UXN+idC3KKFafn5HdUXyc6+EfEOSNeHyLt2grBuL1hSlnpsHb/3ZyhwnrcXp42g3U6V
1qpgsRGAJ9q6g5Hg/WRWJs2JQkcYhqG57jAIIVn/TMmThWa0a30X1sKpWl+eee/T6x8rGWbXsgnk
w5OzmYOmPmBaa1kGYLBZs9Z+gQS6CRWg/z8FrdPr5hA4r5Zxef25RN6pZaRNowRhIsvqmoOJvsW0
NFK5LmYQRx3Ltjt1pOqtCBfsp+mfvt9sz/JclzFBI6ZilVGIfg/3Pnmf6pcLhHjLFMBHDdmnd5Ww
lo/Gl7tVqWaWpqur3XhpqSEu1jTsoMc6eDBBKYn+7ZBTSNEqYv5bvYE7aPzBLY40H8tlKByzmEIl
So2v4Am+96VXuENJXbuGMaLe/tso/x2iymv7jXAuVNY+zsfq6apMqKQIQNhv/yJH8uHjqAonyvuB
ehC32WoT0DQT2ggvkkQY2hNoZY7SwIWwuNHDtCrxk/0holf1h7PIffcqTtSvry9sFNbCtw7crtzZ
2YwlTX5HLKjUIXM8ogMd4A4RRsqLs2M7Hw9dMau1SkgGC9WbL+W4QyFpAlQ/SIxubMdVY8BAqY2C
LZn+fDqYplYSVX6dv8ne9Xc6lMDVZJpn8nq9rAblRAHemser/K3phQWOwBYrmjR9L/DZ1BAQ6SAG
hSuB08u4b+2/9PXYe0Ct3uM6Lq9O9n28DjAycc8HyxfjRyj0M2XmvXVPE+kiwVlIUtTiTnk2uXr9
ViBWPKNiZIQAV1lehwKzZ8iggL1oJS2jPg665yFBh9DIfjNgh8wJpuQj6VKHVomU736WXSgL8VnS
ps0cu4InvWxAujvsR+Cp76Ui+TRnlPM+15DnTF1f/aX+TtEwwwlOlGR5qwkCKDp+a+ua0ZyZwb+q
9DTPlCKEIwgVH2cV6ZwGMAu6JjqfqXo88Ld1HpRn28/Nnvt5cFNtlAYrR57VOduAywkv5VMKwVdp
eSmVeWf8o3hEBGBM+n1kQk7gxUfQMpRDfFrO/4WObyc2X1Csfx0iaSLw3piuQ0AucZdoOue1QeWF
hUxxN2Qny7YmXrugs3uV4GQnjBEDZPVrW5Vv6EJwQavi2rTLja3ZUFppSt0iqlfiMWs9E9ZgRrK7
zKqoz0kvYeBTYNDZo2YjPHD+vLHCdVw89q5JLrfjMMKiayy6n/pUr5bb/VCSgE4myDob1vfSkvBI
QbVCxuqUKQvBGkfBfqck6JVMTqMVRKomB1Xgrk7VTRMuIDRkyWETLEmUATo04UMMIkl+kcsSSdFJ
GNbJm8LUIpP0nQJsXL/Ac6PCXDFcTsGFQKGLt87whjonVWglxlwrACEfArsXXw7uyFn8H+FpOPsd
arbgrMMcq1br/nF0Ilkni+YLxopIC1y7YyUsr6wUY6i4cdVE2yXyCcDe41Nj7AH2jK4iN1S1AMm8
Gz6WdufplDksJVMKkbYvpqnCApaE49gWpq9ECnbxaQHQ+tOFmWUa8DC1RpgF3PlEGxADcrxhLyiz
vWIvSpRW2bAVU2U+dk17JKwY3PBDr7+7m7IkPrxW8QV9r1lTUQ0gHecTLXYJWGAJj4b5tQYPIJUm
R9CDikdF0ZHUDUpHNP82awt3XKdBtUwstGK0VxmwxdPacNpZzyCpNYOy6dVl7FLC0xQLp4y7aEW0
dioslaystqhOhPWGPsqTTkGlsrAcUjTiL4f3A7Bt5onH0Bf/MpuAtORRkNG/R8pzu/kFnNARjibs
ovbxF2rSicIroB+KNFu/mIjZh52OYDYWcPJVBjq6lYGJhsifIoU0rpTI+OZmJPCP/uqrjDkeRl4/
V/6nGavLNdZyGBVGM5ZrAFNjwJLiQnZNBv7JKkEV6sbJPcrmaXdwTBuMeDbrM0Qdd/L9fVKm79jZ
ELNorBGAvcPI+0P3Jzlwi2yjoUp+yv9SHIkOSknZLwCcm65KAiqGC9J4ZE1TblLP+/LGKgFe7H6B
1OVSmWKSmIlcqwRjNgCWEkuS3JozhjmkB5JWX8jxF/bK9EV+ornQQCDxWbOTxrubHgFg9gtLicu/
Fct5pt+HEwGdKOT2nDPwXFjMl5Rp1HeYhOumRMAR9xfU7qqs5ruqm3/rVx5bevMvWDWoPeQqXMFB
wYB/5hXHV0EIgnVdEwRceG0pCYFQNZuCEVwYDzOKlLkIudy7lyJNOcE2mq3hC0ZSQsizlZxJEGN+
/ar/gspuJdvs2xjkOwMGAbeZ3VFe0ewU2PlkscIeRTdrBZWKMNEeQ8WiHnmJGFBcRIbHHjinzZjz
WvvmAu9x37pcQ/PzwG0yQP8oNHUW1TRQMAFV55jdXI6wAV21RBd4n4PNp5LUdyHJllzd/7m7YYwo
t3d/l4VgtBkSzaxd732bnlB99v4OhImkHCqtQaEb5WDxMKV+gizy96J7xvB8nWjWip5zXau12NGA
AC8/XNu7RGkMSoQzUhiPe4+Txibax2Fhj7c03WlvzcI31Qcg+slq1qzAsS7+Ss2kLNZL7X+hlbCt
WPpxlEODOrL0ENBLtO0DI+vPq7OFTHdrnkWnGsc6PXDmz5KBYYdG1BVAFK9ERH9mU6QNWrJC4JD+
+u3Xpj9WmjRqKYD4B17Q9PASQ4bUsVYjAr8SL9l8mbWsqiikgZZjGfSzPkfBNKtFnn2TZx2WdJoz
ckjIbV25JgyCBIIFBuqPPSkrFf3rU9lRIgtKOt1qnQTKwn01Qnjh/hg3AxiA0Yo8fx3XAAfOZXiz
cA1BgSvBb1woVWp1xGykcYxWV/jTZKah7p4lf8ShjtFtbKF6X71f/TrsqliCICAWmGZ7xN4mqonf
tWJNo0Rghiz1zesw9wqEeHGyADPjuaecB0H5TiAbTfyNwygMPmnx+ht0uDOM4h2WJGMPvNZWdRw4
gQvdbA4nGTNvk38Tm4QA2wDsRn8BTTKNseMeKWhUn9aApUfvzsXg7j91WajxMBEHQ4HwD9RPhsGl
PAYnts+1N0XBPAct9uiAHDpnITvKf/2IbrxlpXZij3amroNrLPKSqIcSqdzXmEa9dLkWuaVig+Gz
wSt9A3BXQUF7YfUFbmY73b404/0ezeP4hpGSZ7eYO1AZRW251sojMchRre45DAe7rMI8vlNU+oQX
MlO/ezWb951Ukn5BLrynceJbTUOoi5VWJmzsyGA+7vIOZ44UUsv/OrrP75dAYqZmUpCVHM8J/2nh
yTJTZ8SJ7bH/iCkfhmjzJn9brMU9OnQBNTOj3CZ0eTbeSlf46veh6Me25qJj6HxW1tdDAS+QXEI3
nLf3qXPp6N0Zr+DT7k/kiSq0pk9FdjrNWJRuHdOxwtB5Zk7WtUXAzjSTyNNuLQHXAbY/m6zD0YTM
KdyV/aK9QY9RH4SuUKyNb9IIEm76hOTUrtJPHA2WA8LuJnYM2b71C5b0DSZIAn9oGki+QbXexrw5
bRhsUm/sxovQFuIuV7J8eYdMduAqkanlJX1BDU+CXQCvGHavWmiwTHlO+1sEv0fULcoeXvBuAo6P
FJgo/myC0dWFV/X+JQVxFNHziW2Uuny/Et3JbYObVl893em0vcg0+joLt/hvsxGtkxROOdfF8uFq
1kd/evN1ze5fXjaD5+5DrgbEn89C3j8A0+AGqYuZJJb7/wjlg9yGFVAj0rsqcAuEkRoaq5SEWzqm
6haQSFmpc6JMh/Yafeg6AnV4EmxNR/L+5Oaz5/KtLO2MJdTjgdYj4GjEwgX4oXWvqNJMypgii8Gt
yPLaq7HimkqNyF58spTMoNA1sTk3ZxjKtnIJW/yQF8M5sP0oe9GCpUm32anZ8x7KLy8BMgOYLMSt
zoGSai/En4NJzsfhzIUIaf0P3ehkMuXbPY5reuJfgrO6qk1rJgeEL5vgk3kthhbCLZr8K7vkdKtX
n7CTBmlI1yM2HRAxazQ2TFtiZXF2PSTwEEfL5KH6jvPjvxJfyPJKmoLMhsI9yNDhbGf6V9lHSOHe
IyE9Ick257SrJzXo1FrBTZ4L3Nzntw0U2gLMcIDvM3XWem2qwwXdQpep3fbWoDvb3flC5TAyFApF
sLBYGXZobc+NX02dhykRpIIPGpbTd9HT65tn6UHhnH/ZHYKl8UwHz5urwn1tXju4XNizJWKiG+lQ
sh9Z3vPC7MUFDWo4KfwZfV81HBlp1Z9isXwcXpwZNhzgfbkxisLyEgLEs7xncbGuamhqXC06Oeim
1FSq8dts66cIAaix3xYz4EIcZqA5nL2cMxeSvh9JxiuudYQha6dUX+8SI08fPmQE4ViGnxs15HeX
kI0S7V0ETuY/IdmLPk9N7OCwwok2mav7tIEuvCB+iDAsFNQDPdJ3FBKZS/SfiGgK3JGkar/TjyTZ
d92hhFeJ+/nUtcHsG9lH9TBGAF4vR+tVhhtkJtnDYxfBj8YkbFOPckIstTOOpdiS6Jg6V196gw9J
NXqFu0j03VC5n+ry3Jga76LYRdxYQAGQniVwbPl8paKzTks5Cru8rF0S9l1nUJ7miHMiiutwMA0B
ROyiGZNj3pmnfxwTvWtMaJzTIE7udeMR5wSUHrau0vZe1JNZBC4eZCUmuF9OiPiLmX6aFIdIi71J
JiFAbSnJa2yzeS0wVQagqMjtEqBChRd8UoUv+u8f7vgJaHnJSDoSqR8TwVCCMChqTG8x9uDfduDt
nh7aCEgbFfDck2waisuQHeOR48R8Y9M0MwrOGal58cIcRSDZf9G/7+cYU8I58Ru94IYa/tl1tm5s
jhSzMYTaFL89pRtJwiZxTQ+e2xjEgbkbkkU23i1ePuHUjhzHO9Pv6aQ/A4/An7hQ+Qw9wrWOj3v/
n7IiIr3i17XX75V1ONCNr26MU4DnqeEE0/E6tHd13crv1VIH63cSvO40R0i/FHZyHRgSq4WRR8j/
x1AtvF0Vcf7KbYbXzCjW1/8z1cICW8K9ucfLPTfrAD57hKmazIxv7rtzCLQPZq0SxDOaPIdWkM60
M8DBerm1e1swHcYK62fbDKpOJA6BDkd9DlgbamxQtyARuNthofJlrO4HMSmpsxTeaa5Ln3uOcy4K
JDSxJ7bhWlkdSXerkwETMjBMglmwq3pjvtzKB3thpa6I26OiQJWhQqvQ5kordrNba+x21Q8FD+8K
q6KjLFlKO40k4MkcJZ395FH9VJ3y5uoxwJfgymajKS2F1DACLiJDJjmPMSzbPR0hiRaWj8xUzBmY
u2KmlGvyz71x7VQQ2g5pbcGLOwlMkpy2juuYlEue9cYH0VcBO9b76sOpRM/6tz5DtLnaasmvOsiF
zJV/Yitj/5DywbLcLXHHBms3JZ/k7dJOPZZ4qxv5M7CPPaxqnpNoXBcg6GD44eQDvVXi7NoEfJRC
rfVPhFV064RT8AY8eXP4B4fQNJTFhO4cu/cN7lp6SuuhwDrUjfdSvPKBK0URUw+2KVISM71t26/B
w1Bdlql/0X34yiRJ3+Q6kkOEyc1GHFwc4sajeo54wzUa5tzppvawzxUtA7imiv6fle5gzPvpSfNJ
rvwxHHMEj0IRtEJVXUicIXJSd/sgDQlW7TSdOJTJ9nVYpUDIoWoc9PBTVVzPsHnN4s1/QvBkF92u
F+JxKIWxhlYOyNeAgOyVxe6B4KwmCqtahCnCziiqaxlhmWaNoU6I6IuJ1fMf6ozf6TEtF+iSbHVb
zvGpUUkY/Mmtl4lvd0BVaCC3d36sxoEJfMEpFPV5EIT2BqzB7pxPse+adsWgYEfQXH7KP2MHKNzr
PrixqMHY7d2TumAVnFgbyJM7mS+i6/RaFMrW+u6UGLYyBA4cglMahUIrCd7FmPOisndtnaglTUbk
1D5bU0oe3s0cZ6dzEDpLAX1q8Z/g8sFpjyNgn+vewCSvsU/IpJgbh8LmRBDWf+uUM+7f+gCrhe0I
bCG6rpc8DtNDI/DO7ydDQGFIIHF8LL7AsyMdu8bymV+J3RFdOFOTN8qbf7g24YDk3HZat/dxaxWN
5HvJnkV+cLhJKe+dOYbXWWT/6ktX3ZWNzcar/5KswFIIuqPoBp4CnHTHOnjw8My9lRHLPqZMBNH5
L72l76UAhKcFCiPdekxH08d4SjXwpeC2NcPnRCukusrH3bTqlktmqMDXFxmfkwDNqLpV8kh/zkAy
dL0FMz6b20HhJFEStiKXeZDrDSXfhi1WPiw+QqPqeRUUcHR1iCCkzbGUQq9GoHtUKvR6ALIVA246
YH5Gxs2kW7RGNKDj+6hiOamzMCSs/m4xfbQTsW9vqW5VappcCbEiR6rWc2cGRBh14WLju0uMaRdE
xgdIxhRNBLf+4kYpfN/F4Z0lIJKJu12He00r37jNFAHnJCBTXfhihpMZx51kCpZep6ywfJd47cNT
UvGh5VHKFIS3dRvd7YNVrBCG8AloqxWmtywOrhDD/6sx+pJ1LHOMvDzuEFQiVERhAVUS1b7w62bY
CcA9KmmdJuE0bpmLelrrg+bHxoBQYtkCG0GgGhhZGmsBryPAjleMdSpi4Htm+LJRc5X9ndzqmuUX
KKdhpCzgL2mrxUBUbNKeH6QYlxV7EAUZqm15EewvgpEa9whMjkSaMEZkRZSTx5L1h0+Ks/HGQdon
rN6Bx/XJ0ef85eO9kLPjbUgzRI8Wnt7V8fjf84M7qigJg/8OPA/ccCwNNSwA/QJ79e0fUrtov4U/
q9CtqyiJ7Y1muw9CDwPEKPm/olneLWNnBQJjy0RZHeeAxVntEtnSlhTeoz74z5WU04hvdeF6BovE
cVw9dOWO/G+deqceyCXE0WQBtGBZZRKZD39LinWd3EYLzoRfE+iR1ZUr8U+o0yi8fbucLq7/CWr2
p+lCSkdTjo/9MyWWfUqiUI4Dd3yG5s6uKnismlt8+rD9T14jQb6l5yyHtbRDMq//lQWGRbH4ZiMA
UMjHg5b49JxxDDmCW5oDsAk5H3m3ufhMNzpCcmZuJv8ib6zfTWgloJjdoFfvI8xvbVHUcoU/eLRm
3AWkbqBqGZZ1ZgFGLv0L5CK9oRAYBSxg/X5/4d6D9HZ3wgf40VhtSOePkS3vrxzZtMBv2mp7h9cU
Zq4u0bvBIswp6xfcB+L7wrgD5M/iWl5zhGU0/6fdMkUp1WdRhr1BEOt8E4JuBtT42QCcADPKWUuJ
GoyejfEeNpSPKO/jKVlowHbQiNpMPMxfaMRJ44g19pDG7xJGyA8rj4xbnIEW9dWQ+LnSNFNWHZN1
wlDejymead0fLq+cWpYzD4esHgVhukob54bP3W0tyQywetizgwqldT+KzTMW8nc28eCpxmlReWP8
Gc+prdUxt3ccP8w0ENjQeEA7mSDCEdaXe8o5FyIewo2BEJev5e9ePD5zCfxbjVC+BKCLYJdSmSOU
AtN2wq0mudGqFXW088usXbxcUDF4Hk9MO7wTy140dcuETCj5fjuQSMBElEWRk7PSanI3RYm9qYnL
kc4/BbuMApfA7XPfesYjlv7lJTHLqpXvuyRegb2QbqEfG7/9XDYUzdVHtEAuwUpoHVYS2OGbJlBd
t5qJvKCdpyZBhmg4knQnpD9Rg80spg6E4F/Wcs2yF/sY2ReMIIn53f89ydp69G5xg0fkbSXqKWY/
Rz0BBwUm/qRA+cTlgrurXRx3iHlA5Ct+9Sj0I/REDtXI7oyfrBM2PbmYhHiGHw1+4GLymuAa2UAy
UCQCP/bsa3dMbR5yuhU+mZ3qchrQ5Iizx0rLHcY07qio0caZoF9IAVSLJ6FEgUHgOsqBwANLa0AL
XElg8IgCyiOEaMpVrG2x8FATYwmdccU4ESOneQj2Q7JRGrKmyBesxUVV7E7W/eYm4EJfGmj3rMgm
BS4+43b6xV73cOZGaJeRJuZaOEauW+iCeddD2+SdkoK+q7NvFwDdiPCZD9H95KAhiFoNErJ7U5hQ
0zdHMmt/0HLDmCtvz1xcLOW8NtGHrD7evMcVmRnQmc628ejq6d0tGd2gGQCqpnAoZs2gGoLT4E11
seUT5Xy6e0LxuPRuz6jcTnqCH3/twnT57iZrrRJr3N1iQZIBy7oLMr7N8hVNwpnCQZ5/sQmU/yEx
WM9ukeKEIeaymrOUhj166f0Olt2x+8D2Ha9czNZ5hWciLcyPsdfRxeKJsbKEuQ15qaG6zwtDeROr
ZjC+Fi9FUwAvhaTh4hg+gx0wpuMlx5DAFCR0LUYJRb/c+hNFfwLaDA9z1AlhL0NJ+Iqm+IxGtlsG
ICT8T3sX7c4Wr4Zw1JW8FibK7/c0QUFKiKWzwLRHT7I9DTl0du2TVfUS2tNi1ugrbKtSt9UpXctq
z4oN3XIUpVd+PBumX2wMN5OsuBHMPp3V50VSeIDjL4Je/CR/tgRpVoUNkZZZJ5Kps++GBQRCMHh+
NRHnPJLS5HsT1Qqg8+b+H8xu4UztzoUq497GEiC6r6P1ThWYief955riKsbkMYOOtnp2nKYXS1nQ
9EEsd2ALUQ6Dunu1s7bzSt41fw+OaZtrUaAr6q7P513u5RAFmaVmCo0+Rzefw2zITV1KhFuqS+Y4
gkw1I5B/gVL6QfQHzpaiiJKzIbxsBvQcpqjaNtDvdGVMgLBhXowXWXrUmJXZpa0w7k00DWppy2iG
V3cjFQ6NFp8JQgPnP3I5rI/tZqxBu9KKVJA+q/a0PJEDV3rpTZUoTnFI5Q3JAYujHI76aEzPvB+J
uI2+JLwsbxWFT/VXuTr8JBdQQR6Pm6mBTVvh1T1IYjzsHcqqYSIKLDVbKe1PwhIJ5L7wM91Q+WAX
4Y/d+HNdzQWD4Ofb7hhWB/uCbddd7SaDK6GBKuHqd9Cd8at+4aUWk+W9JCcTtVkH0hGk5J6yUl8v
0knELF8pSjdJmXtyruHV08YGAZ6o3M1pfZSOLuOCrJC7d1O4E0L2nVCsNG4e2pGt8LdHbTDM4Kqs
rlPBvKGfq/br6erdZTTfX0xqLkBMe4gf0xML2x4DMmPCoHhQCh949FpBUyUX7gkOscsx9FVnMWpt
7il+nv/MR6/v7N7dZlUtLZ/lKTMk+sDMK/uZDpOqcs9kk1KLVLSixgWadYSEIYSx76vD0zfWbV8s
BjeZvDToK2SoOAjUK8zNnfNxEU2mutzZiAW+5+mF639iouQpudxAOq0VrM6XDqjXGgBQUEOjKSaP
EuqrKJRg1hTiAa6cTj3deifNDv9xFyWZMRS+UMYyWlR273ztOIim9bnEDufho1+Jcxfe6vr1UX07
YpR8e9ffMD+1/8x/Op/6eJoPdzGTJ6KcBrHt6RBMWTajk2C2XKjL8dZ+/T0GLDQiziKTW9QAjjkv
9nDrxW25+Ar5z1ubsOKNQ9HXjHKuRdTUE6/waT5lRQrWUbSZA5f9YJ0/4YIedfsH8x4iqeD65yFl
e+jsgqRPTVQyTTUYZ8UzLJ8JkckOsKp227ML8Zst047A6FtxUJA4DhY4Ekhb+62mY60oZuORHpxi
L/+bnw7PnWbTP4/NpsvCQuYdIBa8Drb5z20W+39z2n/m+FfGwGr8/TKDByTzYG+YCivyc9Qkk4AF
uCsxIYyg6Z5bBKppJWJ4rXeYlhHbmikgrSWwK6cXuolCiZf5Yk+ICAKmm8RHdIOWqxjXotT/Eedx
C+xC5CUjDjcHaMaacT6Op+dKqmLqE8OdcqoXAMYBolMwQbYvDE/1pd6M2vJDhSm082lslejUFpyd
1M/CtCQToYa83hsIqlLw21VfWiLkieWZHbAakw8l8qfye6paIOtEBnhPVUuhYpHEWyOcSflmJppc
LtgL0ZvYYvQ2GuJ+6rMP6fMJJ6yADN0R8lBrNEZQ6VGHOYLaybdZk00XGBWg+v+3D4Rcds4ID55Q
ZuNZEHvBsiJfLCSVJG7j75gJbeWd+IPymXSrjC90zgIQsbya3ahbEunac8c6qLzduxY69fyfTTFa
CIRAmmAeIffAoDMS8DZKC48RDXxmpT1EwAyngRTTm6YEf1zxumtDV+ld9G6oUL1p/QSjjldsaHgv
XwtTYB88Fh42ltTcAf3APZT7rQzqMd0W0KmeXQG3tAFvCVWaT9jGuSD3bZ7TFNL6n71xJRHOxTQa
R/2YQm7RQootdpWLKODBdJ7Y9vHCAiwMyLihn0/QuSwAr7FI8izfc9uFXl4XI4nz+TfIbOB2oxQN
fxZXIkmD+oAtyyNVBkegVDxkD0pDGclrS1xxjmEsEwHK72fzQ4LfcYgxjHADqmmPlDh/+URER4NV
khGZTZVGzf2XlI3P2eF3X0++ad69FHUrTWUrgELtW7Eu4CBUEu47tVYVGFSwpN60g/JxSu4h3GNT
CfSWQ3jRcjoynDrgPwyIJq9IaKjhlg9nwwV/UENc1cXs/xSElzBTmd3XzWg2mfI+k9t5gIjqnVLd
27RrrF9xmr5zyaWFaO2U9FN1BHXysYIL3lm7IIYSAp2ObYe1c5TPe+hT1jUK6nGZigOkhfETNDgT
0SDCSo3NbIxNpDzYMxnjYymAMpsfW0X4IBFO96ZbuO2TNwe20x1vuEsfBSVizlk6L7vQ686GEUXB
BOuZganjg+ytimikcvGOdLsswSca2CTqsEEEmTigeIRgvnzCFxm1QCZZEi6zXAEg7KSpr6FRitNm
YioK8O4otSREPJQK/cnKLn3opAIQ7oUdDbbauZNEfCFJLZND7YYGcSiT4PwNgDnInTZaCRXm6D37
QlN9XIW5+/QimdYEr1k84vDT+GkaV6u60us/Cg+Q4CTnvTIjjfD3pBDpynx8/lClvFmhKdnLZ1Uc
uB+ZcYoHhcut1i0/IXH0py1bU+b4t75Bk/WzpAVyKZlEklpugwl+JyKzI7Gc6vgX9DoPCgA/LRRu
zEygYn+OiVU8ksdnI7AQG933mjQMRzUFp86W6imLBwBfdNo+YjxihvkTJjXOTZAMSaqUEELI9tuy
GnmkeQPtMvd91puc1Jdy61jX28gKziSWB+6dtaDUDtWYv/XrQQUzFhHxr61B7ccerqsIkzjTyIv8
QSrg0CwJK5BvOK2vfMCuzK5HEay3mCvjz3hj9zH2I9AaEBmZha5cEBgeb34KVm+zLyrhhW3YybeG
jICPr58GQdy5+aRx0HX/gq2bjdpMJDsQZOzG+yW/0IMZvejt2FRwpF95DYpWPp2NabFckKjV3b4r
uKQ/0H4/Zrxeu3WwjEf5AbPi7T5ezI7VoludzoqgarEJpdqHRKnIevJAc+s9NijQhZmHs1crZuOo
QmuHj4SI5NZk0WJNG+c0fGr0tOCfrWkIsnGUMJ0kNt0V5Q3mBFebt4vsWC8zGcAtgrO+1aZmWtjs
3m+EZU2oXDhQQ4ot8wUyTPAADxX9dIUl05TMM7POAeVUv3Z0ICNOgN9/+ZPuiLV4/s7bRcAsL9y3
q1HaY6z1abXuisDj1RQ1XXNuzFsoEK2OqB9ovVl1QT5Y8ahu+ymIkMLOeSrZqgHnwc9QZODSAkFL
ZMR7Sgg0272C3Bs0b68VscKofo3ictF8V1ODSilmN/WuGpr4a8r7A0xdxasNxhmE21cWeI6HufMs
RgbcG2mRtB8nYxOD7BYoDrPwQ/djgQI/jwTu/gxRGxUV1aHoU7He3ocVgrcRGS0rX0HYPeUvjif1
qhwYfzLqSuDByVIfxLzGE7cPo9XzNOEPzjVJFttahwC9jcf5D5Ccdcylaxhc69gQgIwPQ6DeIWwF
wrnt/axaTlnofy1UnYYqFUsrBu1BYVbAfGpkZGAE/Q+e63fpeAoHdU8eyc0CCplLgv3sK0ysiGHD
8bRZ7OJubrpeYJZ0Xb33xNrXAkOgvIQdYZYCbBhaBQrSZHV3Yu+/42gjr3hrwfRAyAhnHlSJV1fd
rZlVbbmZuhbtK1zthVqQ80767yE5OGsxYGMMhmGcFZ+yk5wR0YZu7jy0iSqupCeoNq8PLtMZppmS
0q0+XQa0wByT1MwqFJHQQe/Ii64sF+IRY773UE0NunEqWzgXM5T9YUQe16PdmvcU2/jYujI6OZC+
nxBKE0GQL5tXxbiVvH+PsZHUb8GqS3uqknDQcyt9JuGq81pPae7QZyuHJbHNr4ntj22nwBFWEu9r
xYkVHSbuZbsQNNZzsBm+oeGIcYU5gThVVYXAQdEs2Ma2wTerThhmTt0yh2t6SE+d/Egdeg1rB8XB
cd6n1uB8Q5OtZMZc/VbcatmJ6ySRq5CGOLwVy5WxavXNBObtmzZCSuD1lZMs2CWQWKn6K6eGpSG6
ZZjj0qzn+uF43BNfFHLIlZpe68r6ZFEkGgCQIQyf3Eb6PClnMH3gwKD/I+R4NeS/ZrQzvf7ImBkp
hcpmMcZwfIq26sCke9K+O3KNg9BmdRGj0orCKHOxxTBI5VKXissrlU+2Jle0Tn209sKThLu55dD7
aunt5SryYCKQ2OiozEi9dl5mWVUIVGpgS3CDWw9RhNwwwfBzHvTbw0AhcTJTsTXjQYNxtLsQsEiF
gWIrYZ01K3paxhAiS1FoHQgGcz2CIGhveq9Ba8dlkBiJ1EkG6APZC2WmH/BH54rPHhp45iBgDJ0E
jRWR/xXgMGdfETSxKQwKvF3X3WGV2MEa5yvOy03dbcKlItlS+0pxOBbQmKUPcG1sEm42/r8aWw8r
oV6ziWxzpc7HQKid/OqncfnOP8Pxk5GPE5fEwP1LykSLcfXFxMgvp+NleH5wJDfcvo9TEFssVtkX
bc1RTyYKy/lgUTdkYOINsUKH1tTxAiMMTRdksvMLcMcfhx6/vw/uWolvIIjofQqu05gqhobymw1e
y3aDpdaZQ/XKjhDdFaDaPBFcc/lHIhRoOk9KJ+kn6wrbeQMpZ7+bwGHBPkaYHfwcGCHFL7NENx+b
Jf8rrnTyjTShMLXeAVWzi381FuOOnxDFDnY5C+H8mVa7MPtKHG5PW6ltjZUgSjiNOx0OAeArcsne
ZG7zPbJjRjSBoLKeHCdKNNKDARHjb54Cu/MuSPWhJ3f/qEeup4O6heijZp13RuluAbT3qWmBlhzU
4Pv3ODEwUu9OPWmnDlM1ydVTO9dm3FX9X1MAzEuQ92WCoQVOz1NNTQ5grO3+KDZaomQxgJ10SxUv
6B5x5OISOJJ3t/Ir6sThkT5qo/AyCeSvdzp6qvx/MME8eJwcQ5DhC9JZN2/kskhaS10MNytwsLtr
KcWpBf8iDh+wPb21Jfn5CftMe4mD0yb381rv6UZcsCNJz6YqPZCeKg7LQCMysuKq3X58oXOuo5ow
kO90trLoa0/d4EuCC43EOH2yPNVdoXh1C+Q1vROapMOJzweey8vWRJ+dfP7ozTmQ8yI8xk/BC8Wt
FQ+uHJDupd2u9C5aSWZ7Y1VtRXnxNm9WA1mwQ10Qe8f2EmgUNLeSCoLLEECxFHQCK9omCk79Jktn
pduCiVujRCZoAHzyuB2uPocFK6xtUJz42lFIaAQ0u98S//M9pu1/gD+zCmFVhx/g5oGvle5ytLuS
q8cg9cecdDPfKGq5mPt4+7Uh9BzhgSwInpikUhq7+41bxQxMJYPEMiCJaJcG8cbIm3OGNXEy4svr
ubblolnSo7ieRZTiGJ9n6nKRxYheok214sBcNZU0bkpnizNoJ3Y/9dHvDMqk/jPWZE4HwKx6Wa4/
/DZeSUQsU8Qw3vULbrB5NQZoiUmIoNumam0MjkszR052IoKrNC795aObnotHWuXhJZG/PQV6N0hl
wJrKlo7uG410V5WdVQM0+Tp918i2Vxi3lg3NpjLYpTEn9lfFlYppD6dge/RZudIa1MW93hV0uFFU
WzxE0rLCHhtdQTmjsyt5RUuYT4jWWnSKEJRVdHk3kXcQFw8zsFN4uNkqQrRlSbAl96g8w7awfIuF
AqRL8h6T3X2L3+/WuMYqcfw+WsAO7y2EaKGTgsRyqFwYx0TTDKkLCuCDMoRv8EiNE6DB74ulwsVM
azbW8U0nDksPsd3ZQ1ImUmtYbkSAkudBe2zYeex4rZ3kNazZCcp6JP56VJy74JYzNqF+gez2U722
MArR7+wIVOf680rzUrJe3KK6qGjR+G66bRTYbrUiD0kOCCqAjmEuoMJnIcDfkVefdqGPxresPU88
7uZTPSUIGqlQmsPG9EX+D54fvphhiTADgD4PbZ5f0ntpQd6eZs+rQotX8kf4FW0BLyRRmE3AqX1x
0c6yoD/wCPIAVlnDvMk2l6RFRxR6zxenDY0iwZ2G78rOB4Y9HhRvZoB2Zn+hBv+JWI34/wZ1blKN
sRJNmS9E0GFIoRDz9RN5CTprRHbt137eVrx4oIZy+E3adgfOGrqshT4uhT5kW/zXcbZ81mewU9o3
JJJHnQJzdd1ldZYUyYKWx+o71MSFmdxIdhYhHPTj3uYhmOlLFbcW4vwo299lU2UhVE6HwbB6MsqS
+vI6jJBoAsII/jfiG6VI8tWk9k8rAmkmEWM6a1WwGi2xIICnq08DF3wMFnQykKRFIt03Z79BUblu
4rDZlqVKCQExx5xx2bL68AW8iZNVTTvkVNYbqkc0ZuVl6oX15vKZ5pfq4mjgHlZ49QyUEeNGJQ52
xjHE0NY04K9n9xFWo2FtFflByxhXgQ5sc6UsPD8yL9d9tOGCfp+++3j8r2BnIHoecD1Zs88iC2pY
XdRakeqkwLe9IlYHiIGMgFv32lHnHiOXo78/M2fA8WJ/rua5valB2jYjsONN2CHjS5BjLabzvCCq
e+U7SNYKOBxlt/l4qDb+GBCsGobMtkX0Z6+n3zyQuSxToIz4nuPuyhF/j5hInqD2Mxzih5+EV017
u0D2qBzYXANjCnpNM77weDvXB2rXoPv2GRFJr9/x+vdI5GXhqu7CM/EhVLmJ/On+mQ8Ofa11fokS
p2Hx04iMJlMquscSSxo83Rq+EbdygKKHbO8ovwR0OXsEAXjg1NOKXAYkgmF6KO6Yh/jnKlxcUht1
OElLyE06RCSLhCAE2uKFFcLIquVcCgJb7U7E4uN9WIto1X+4yi2jy1RUAwnmdllG0Ru7j6GwvZkX
/5OnLP7990vmRgZuahY/KfgthpYQuwQt9WTrjn3rw+h/QL6zpxr6KaewPAOzCADpliqlir1ed5wx
8YBvIsCSTJDb3sgeYplZl+Skg+6CnPOqy1FpEdDQY30wg9fExB8vKQZyhFcBJpQi6Uo6VSmjLMfF
R2I1+JvUQhWGHIxUjfA5XhSLkM93hwzM9S8S5Gt0oZamPGvLJJNepJS/1Woq+ZbvacKA0/tEN1GY
P4cEQOOwbrPhDFqqpQ/hCJemyYW/32C/0dT4FEYT9+0rVBaYPoMW6l7FFzeEp4B/FSykJpaPgaUs
sFtwIoYvOkWQFNgssZT0h1JX2iMjK0x034tLMzTtvAzD7bsoKWHg7WxXhFipNvo1CDxr0kYy3tkf
TRYWhccSJKygEm+ZgAt6Pw2xx1AGI3W0zy1beyxjJjOJNaMw10OC4ZNxzJgFGQ8Jx9g8/fA5S0ov
+SoVpHCky19lKj2VZK7bO8B/zcuSFbFjH9wQJzDvoGC8qBFkdXwLw6mViAtdRWRAAPNa5jWelgms
giAaiM4GN9GlTcKPoxQF/FuBJQTc5nROYwFII+Ma6I+9xhNS0GZoWBwz1VAkAvZr2wYzAtArTdtK
0B3dRO0gfhohDdDf3YRP26LbS16s4UPI3CPKB7Nw/srSXJRkBZkUfcYCiQbMJN0Jr8H1b7+nX/y+
hRbpInDfNKq4PMwI+AmalPIFdKSsPaMxFMKbNtyxxmc6i89OKXdOxL7010vb7BeviINKQdHMYXkj
2V5HksZj3DUGyjXDOpWP2UeOFgv/aps4ZSGLGLMWovH2OMe/mH7nk0yRv1Cb6cUndIZ+hT6bzxI8
mKQwFdLFoK+aD29CMCbqB84FC11ax5bkvjqHLYVxM1CCkiQ5FAaKnFVrgcIQRF96285PWmpe+6rz
xFJSSoAyHoZjozFPmo2DNGERYW7BAn1SjOXBDH4YJ4vtsbTrmeUOwHXt5RztrIMdQ5i2YMsMiIJ7
z2kAXk5ncqSoU67eizHsJMbJbgQobhHbDFqkKqDuFO1GHtNLOkQvfkLkK7QI7HJSxXrhqiHZjprw
RuyrebgjGahljKBsqziozma46BA22HZ72oyP2dzJzn4puxSLzqMrpbUsI1IWX9/oL6dsDwvChRC6
cvtPbsLIE9iY+RolDf4NDM3caqsLIpnAa7XHzNpyo4CZHU2ednERB47zj/qt4mbGAl3n9SiFeR7l
JD02hnuthRdtL4WZ2Sa+HH2fLeHjHuVLf4gc42Lb6nHV6qpiHVkQ/dpThucXcgviZItI6WCX1Uw5
5b6wC+DRhXen/Rrad2BlgnbAQ8J2Xbkx+iEQyJhb/vVe2nqroXpackRdK7nKY8qzAoM/iLzTZJ3F
YygsOaveZ3w4QKbMZ5O8iIqj1UHRqu5yQzELFAXY1OejQaoRZXXb1OPjZ+ygq6PwpHXKh1FWYZx9
hYcbshHjvVLGzNJZXCll4B1kPhFjnfRa+RR8KubnYFUrz1jvN5CTZ+LDWZZAgd5q8qC4jZu+Aq9j
6/0/lhGtAkSUKNPmXYIe7KKt9ly+kPDEThQVPOjq/tQGOk7vVlZ3+NclCs2HwI0olyKHW/r5sEwg
urf1CftLlGnsocFY7cleH0WxYi64O2tdKQirwuRgPpQBYY/fUT9/bfBwjqZ+rG+I0rlQBjHwdyPX
MOyzNEmVw1BtyQRtFMhtIa0+UY1uo9Yqast6GxN78I/GSxym9vpCeOs+IeZYb512RViT+Oe3KfHv
UCIpII6gFbASkyhcnBX0svNIEnUTChT6JDHJXLJwD23GtY4wqS409EQuS+ZlX4P3IJxyV+XUcO4M
UVsnezQrc79WJ1kZyluxZZlnw/QDhGhH1AVQ5afmTsgJEYg0biroA9bAp85ekPff2EpKdOWExOjo
p3zcVwruvtL41NeBqZJiDD1s8y/nBTdCVRk8c03dL0HtbrsFjMLJX4Y04EJN2JzVK01w9J0WAPpt
1RkaVgXIq6hegt0PJf4TTLy0r77UgiCi+1veFDgW3hzSc/FW87BUVzLillwG4moaWZx1Y6BYUJBQ
NYX6TIgCITkIqQ1VmsayBtwNpA7NM6b1Qb1qhNaHx+Nz2AWixYgJIxc2hz2qrTjC5wRrYL5xaAIl
Cz27pL0U40D6GvGZ0WdujcLSVAj9rYrGKrGdZi92zLpHbThXj91guB0YLc2eXqbtAifoPlXZNCU1
PyJ5QMhVzIB7faXqpLHHiheZ3Zoq4M4fbp85KElgwXgHEY8VKZe2vMg4XQv9rKHzKb/eh7n4IklW
Ri6uRGKShX6/zwYHdOZAJ1qqkfoGP2caX2qxa8K4CJHpbivTlwtdFC8CKT3MAUv8mvs5NQfI5kP0
et0y9ylb308FVMdG/3BC2l2qy6ylLhMiSJmnx6OC3thZG4/Jyt4JQ69W+PxCDhb60ZTBUQYNuowH
OxTAIMb4Qg8THsHSZa4uIEqRJd1KmRR/xF38iMoa/CihuzYIWNOJaxHOKBvBy1douY5lXQbaIEqK
QNwoiki7ZzOhPUe6ky33gxH3s6NZeQlk8vtrc5mRpph2bbkfLcXiGEfIKyPvRlxOxQDXDb+ZM2yU
MxA+OTKon55XLXS9lIjp6pSZ1jD7+OTY2dRaNA327xJj3YW+WV1pEaE0Gfmdhea7D19brgmbJogj
uCDhZGR0iW/V4CSchtwrjYDdUkKJfnZFzgIjg3WnikBCakDFCdTKoyETsB5U9bMTvF90kYg6saIU
yFImNgRYs//V3fKpCrBsk3oKf1NEkq/spC/lldfebke9AFdJBIS6Qb/KIQRbeLAcinBIpMn8rAtv
JD8DZkHD6KewoEC6dREcQsiNKd7G1JYX6LL5JoO/6ipU185B/SNuDsJ+DMlvRe4lTH+O85iPXQpb
vbgXo1BJD1jrcr/U5YDvzA8hEiW4yNZIo4TecQagL2T/gwlhuuJN4S8PSACzoW1J3wrJNmAfjCXj
2LVfxqpL3bKEt17j8LMtGIxm4GTNHArWnrdAZ1r8mnyD5k2IIODzo8GWzUpkT82DbSYKqqwNH467
z1kVpmnSREPOoPyYK/0kfqCwIHRF/5F6P6+HZ/7Bwyf7buZnEVRToVJr1wPiLENs1O+J2RekZfES
H09oAwH0NODnHS9w53aqOuxUr7USADPw3vFxDUzqOOc0K8YHrMnOwvuogMlTcO/CMv6sPSrJzeXX
ibg5z6YeF2ur/57nQauC8nhhzREx3Sw2XKYzY8EG/7ZEoVVvU4KP2RNhQaDfcCGbvrMIHM2PPIKn
qzdHsnCVmJiT18mZAeCqxZdUXG/hVYVzlSLuS1qa9Ylx7mc8Q7jy7huawGp0BqS60yt58hpS7QgW
cpJ79mZA3KpYR7vRuKKEo0xwV2E4od7U5m0wTQvO/XA4mj4VNK0aLWhMeqfg+gpr3Xd/qr47l5uN
huIUsNjfgsmZ5tMHe8o4RyHYdOEvMrkfa3DBzXHre+oqDhOfCHhN1+JH57K/XlbcB/vYyElmdzuf
1jPkNRsNSuGJQRFfNIiK2Oz49hoFLUVEpCdGPP5NpRhqWVO7+iUR9fbLhMEBiwQu2AR0M4WxcryB
rTLrLbPs6nyF/kWmk5pHlb3+tTLwhXuDxuAtw6o7yeRo+j2K+1mXebhvH/EAZQFa/0Uc9MIUm9vN
ct5ysSO3MctgqUFCkFAjTqtzQUkI/Kz16fcvmWH2x4wOL7VUOtsgqA58MiXe993pDc2ZAdd0v1qT
zyARQ5vg6YS71RYLZe9H2VxHuBfakW/nHZgZubIsspP9bckNaK/TZEfl25wHSyO3dP+fZQVODW1w
poYB0GXbjN2wIOxi6pXYldIYKLLYH7uPSnCDjplHlBnemDq+meTI2xY2rmyUu4u/J3nD3LBtzSgf
u7L4fDzOEgwPL9AvtjtgHnmSIX7y2zAxh8Duc1aBK4d7xuX5T/Ns3oUEVmjJ0li68xwoArCTNNiZ
JcBIvLMkwNiFY4cGsbGRBPJPp/vU5VzZBdLbfq+LoFsKFXkg/27vJjyXiWFD3YiCYFq9g1UMALTH
/B4pNHH+2MTZArHhz71aiJsGdf8Apg7SVoQNYOpj3VYOqwInTuJDiNAT/7h5OvNlKnN0mPF7UCNJ
fj2LPB3Nls7oTGiEkZPKyi9OcNXA4HPH4Ea0UuLlo6NX3kljnQiLihFzux79fkCXT5LS6K3ycu83
MLOVwGm8Uka4CIbz+x6K8eP2aPm3RkIWTLMomoneKcESPT62Oi1ZIoYuaK6GmHDiVQCoeGCZMS+Q
CrmgMKVc+OZ4pJq56QblMt5i8C5LeC+hzS863pw5PiemRNXH3Edo0wMtFmPh1vekNVm/1+8K3dbQ
BO9ZZjpilftweHxqaivVV106x0cZ1zURxASxuOTpjGh7fbkOA6IMHsijuWals41bFgwNrx6ctO3N
rDSl/L/uU/sWoO16RP4eDknkGE5xEX1Tj8N2XSrXlcDdID9VFmj2twlntUifKYOYbnzoxAs0zNHd
zn3WmDzKp59jT1/hZOOk3EfC3M+7CwGlLtUehFBMgfS4yvE3DK7JSooOIBwAUUKf9jJLck9ipo/w
xEW90GhCwndsgnCEZp8QDgeAbUTYWb48XIRoyaFqIdJMwKi6zCfDmk5hP61Dd17eAlELgRrbEHWc
6dlrGzzkHmtAi9mjqAP3c4u4nnNJgldP5D1tUBONLMVwwCg5jZ6JBijPgkyq/R+S+kRzQAVhT0fK
BzOFs29FzccFINUT6yJPVkJvw+1qFrXk8ncxHbmkWbYXhJCezAEsPJCTbry8tQzmC3UyTYO7OAFW
7Y3aTdUa3QcZBE9GVtjybVY9lOouoxr7LLfWUdMwhWc2uT7wpKfc64hfKPzHMrhraWGwOH4ZzMO+
NnHKypDkKlSJmlnk5Faf5mkh9RmnHbP3dsOYUN6D39gTvip0pjmLbLGO21Du0f+yJh/+hAq+Lua7
vdZspCAUI6fi56+lWSGC/tpqfXee+MFk8F566IKXOS9sBplLV7U8AGquvI9Yi34Z89J7ZvnAfnlr
4cCmiCS+lNKcrIUAIFZdPFk00cic98gYstLoVew3tDjAWkY2wQmYFfkynjZP4Gq3z6n+pXoT+iLI
8pAL6ptnLoHNxVEVf+dF5QMkvk6+nLwMP7+SUAqT8XuG7YOzvHuwnxodb4fDIrSoZcN6JFoYeCo1
dYQ6bMkRRtOngSa009UTVt8FO35SMpyy2ebT3oUSfUEMr+T5TEt1q8GpcbqfetLJnN7sU5kOZwV7
gAMV9d0yDOqAuRbOLpivers3se4eK+crXFptVCP0v/xovdNA5vDPSYQ2yTa+dC6xgtfOmxCu8LJ1
oCA70fc/o8vk3CzIEm7cI1xUPHLZdVNbyj3jhNUx7OEZ++hTc/p2Z+DehGzi5HmwrOCgbEMQ+06X
b5Qr/O4jtIjlpuxl7wGhq6cO1nT77T6TwKKl9t3fDykN1zyVFQy1PvJYGK0GimqfFGbsz0eBeJAI
sx+6KIRziE/eG+/IwtH7CZGK9iUBNZbdbe/fwJte9fJnRQ+cRs9EypFGn/dQVifrC+O1UEkeKOPh
9QkrMhOtnK6w86xfa+I7RNVd82jBQrgNiGJeMGqDaM9W17rYs2ZTQbV5DdDAGooanXNdvSo2g3Bg
taYBknnllns6lxc3P/B9Gza+k+Xzre2VYY9VluQKLxDThCAbRrO/dSQBlc9QWjVSeAb4azBRynXd
FR0DV5kuaM5FODigfxO8GZgqM7WscuEn4D4NIXflNfT7ia28YlN2px1sgnO45z4G8kmAWSApH/tt
7Li+HJ9UYz1CaMnJB7+LfsmNt3MoICerA86uzePtPHffN3R7JBw07+2Yqen2ZE6T0ClJMe83gUzp
eH+Czf3RAiJRORT3sasRk728hT0LuBqiF0DQTVpokXZorTvnKoQJTDKiCYQoq+xfKHNxZTQLyyro
H3N8EZ38k9wetYhiwvUpNfe5XJVWisXX5fFePuZg+j5muCsu7Bjk+lFevyr2vTnx6ZAkWpEEIWaK
O/a41nyZY16MI6oadld5nUpjQBAqLouAGt9wZfOLaRm+GIRSQPmbo5yx9VxcknyT5pO6l+FfIKHj
voBcPMb/GcLMeSu6oegHMRe7nnoEVTlJGkm/qyPzdqqH8Boq959C7q7moSYFhEA9/E0PF5k3Kaw3
iaddDEThIAV55xo4klQYROpKWtqo0WJcfvAVinsa0k0N5AnXTycRxw2XcyUGVgTEkAuAUHgYAW2A
w+Dkube9FcuPsesN1FcDpq/nx1cuWI67LUYyw5wp16xkD25GGwTYw2K5pZmxBrlRMtjqzB5XaXXz
slrVQZIi8G5F/pG99DPtrZQpyTdKhdm0yLLDLyAPeqWpwixVHJxPi0d7OMVl90VnqFHnNwdruU8m
Kekv3Z289DM2w3XP9geepi1BnvIQBfhM2Qyc+gRGl7bfUfgJi3EXvlaKjdcjCMh98ma67FS+inn2
PwRSizrOD2wJoZQMUJIXXkVDfd/pYV8uQNlskgRRuvCUOzToQGiUdxhwAXln4FKRfBysCRVjSP+Y
xWy/NP86kvTGmbAGPzIvx0oyDV47p4A+juoLeOVOcyyA1Y2u5jFro+72mAK4Yi701vSQrORGwyoO
pv9EW3Tg62wIfZV6XSwKB6ArqnyqGl51Vp6VBm6IimYMISLFIQbpThtrdmUDTWtQQ9m46iPN1y5g
LTwgY/IpgD8NIYlPm0aH5+rooWjLM6+Af92vIhsbRtJwTMUPQGvhKRxFpHrok1fB2isBfaItFNnP
U9PFizBx7EiZQgV0CDbjDMnliaDE/td3GNKsQRLJ9dG7x9DGoJaOmiYgMcjberwL3aE8GxBTMOMl
StsP6EdJYm6hV8P+tZG5g6E87Xn2GrmpbwpvmHh86/k95jZWxyCJsxfPLqUOU4mfbaNj7FWYTzuk
AR0H+KJinq/G8RJjpYYBNo3u2W5Xo+y0tSerx3kcCo55i3bWF3HFx4DU6wAs3a+tdwMBp51Pf/SR
wezRySOmDT+x7yS88r5wwKye8frOUowhofhue9dOTJGZwiiiOG+L+HjzPxKzNviS+nWpyLRBEBpo
MwH2pT0beDYzqZ5GWNIR8+S5ExmRCsTEj/bTq8UJYYesIK7wWS8O1NPWgauNXv/HpqKIrJD5GnQl
lUGHWz4bQXXgUoZBOsPAFgmKGWZyx8EvkMEp/OjXAEzKuuSMfQF4srpN75BZoKJ6ot8G9HK7lc5f
7Ds26g8giS9fAHe2fpkIjp/Cwsd3O2nR5iskGfr/DFxZK3T+2MsQEPbVhypMRaTo2JzkPyRrAK92
/lqbj/M1MMTi+g9zGMW6chxV7qjKy/N5rBJCR3Ahr6GLU7km83f0f6RoP6gsoF2klhMlG5f1EJX5
0PjcmDiYujQ6ZFUfufyOViiATBfdYuunO7lrX5nitTmA7HjOyoVvAbiPFjE/8ilqEaOELWtnA2Jj
+4a0zaT5AqsbvMkDKsD9ePvUUfyrNJ3ShDKIqODIfbmgcqZw5jRrHjKwQ3CxO65xrR1jZGow+mh9
L22BCfq/vvZi06SgsAwe3fDILPU8F+SpwgkV9snCHY955zn51V0lN3nI8mtGo3n2G7yHur7rYtWk
bnVeprd8EJqG7zFSt88PDg66btPlMvXxG8E5/l9L/wAl7b7PVzjBjhkB70e1Bg9vTVcsrmSSJtYy
dG/NI+eF78dI99hjbabaGDswdbOeVZLbZ/2samaJJPRfHTbG6YyJadhIxt+bHZs+Z7rNPAij3kkt
BC/YUM8HhaAJnVCHOGJgtLetd0Ka2FmAcTdc7k4RU4EpwxleWHi1KtnHOVN01g1xkJPYOIqJws36
xODeu36u3UEOAn+QqjsnoWFiPlfvpUUA+2ey9hpXrKfzuYvd/qPc0cbSYFS1cXbVNm0m1CuNbfMg
dE/KtdL9qsve71UukM0Ki7ZDSFyIVvodtGGD9ZgOzFVoyuCTkSGnVGAbXvdcORURJ66xXZGfrerq
wbXW04jTYHBdhIQQwjJwRbh38gXb/43gdVfxvKqrnp6vgZTXfGHiypxco0ZkV5MYJxle/TlH5ZWK
RYGX0UqxChsseq2tRMPnjfsbNJPbfDRA4AW3EiN6BtXGzdVEHYniwgU6WJtZovZhYWdl9rZQM+EB
bzdavCZ7739gwarW4ue8CQaGCidON5grCyUY+g+vdALwLUjUMW42VI2XUi+QWd6AQJqqWZQMRDep
SM0svQfV+52ZzeO6XFUlHxhcbnZE2TBiP2jzrzrKlWltOJXLMoxg070b/ZcRcZNtEydQKN8LEwXi
z+HFLHWGBp535622KOdTkytIMPrm7urKOxfuGnze5zxA+Gfv533HG5GwUeRfFILUTP1OUK/Eeg1H
P7P55UklXp3XghXQo2EqJEA7G+qaavsKea9BgfF8ZbJXwBTUqgXspZTGeWwxxFFMdNt81hrH78vi
QpdnZ7nz93wh3uo/lUElIdIewMUUoMDPugXcv+uM7PxRzthyS+2ApTE/aD7cskqHMwKwWntLYyxa
db6pGfO43dCQrpQVs688qvmTbXs5bfeG5xRaQiEkTbsdaPiZ0Q6hSmGj9VJh49HzcplvaXhY62cc
Dv/X5NxCx54IfphNI6lPk8tANm+YqfcY+2+r2L5pkmrZBNQfobDwLOE+K79N9fvvWPV9KVs4FPH5
A4NmaBQb9smkUiuTxA84RjNGAxqrcxYpdjR5cvw9hBasK1Tdn29SoAtiCXL044Ux7nZVTbiL5zCy
NR95fBqNLvPh+fEWmdiyxt/7S4VWOTJHRZEgcE6RufRCK3ePgw70acnzafcIwH0WqsU8VZrwzr5Q
17urR/YDBe+o2XdA1KifuL2XZSZjHeR/OqzvTyX3SjAU9DRPMy3BuYn/zP8+bORGb9EbMVUkgDZ5
Eclt8hNWSjlU7J5oJFo8STcnqc0vATr9yQ7akBEcjbEoFr3ghOu8zWSiB6gr//SWNHT0H9bTp1O4
ZZZxPX8vJaOUGqg/W/Kn3KDx7KA6jnKGcKx6tdryIvnC8nNgS/NDwasW2PFYYm1I9grmDXJbD59i
mv49f56NbVvycLZtyWJKSWJTC0CULAdZXxEaGhMG+WYfyOewAzBZKMuTmPzyLECgiPuDGj3B+qnB
Oggaax33fb9UbjSYqKSQ/B7cqKOiGwa9fQ5VqmBWN7oo/38DGFJNR9gjF5TuY4j+UIBk2lWCTeu6
XfuWyU+SBUrxNkH9ukAn+jvadgLwXnTu8mEeForIxwpVkQW7g9YmISKY8JyEwG6k0/9+WIY9Gx/j
eOTU2reIWuaXOMkrM40b7MAKZLb8Oi32auNz3bQxR/RGRsxOpjtqZy/HY6lCQ+8HzBNHP8mndunp
Ee5ghinL+/3y2X2cYws2LuU0RH6+nbeMfV+maXDFl7L/cJAxL7NsVr9IdpU11DxkH5SuS1kUpBYL
deuUO8Y6sVBu4F5CdeR/4h1PR4BIQJV/+z6+/wwX3eQxqfKOzTwEj+bp8zlcXCOgBECLIig5Z4aZ
6yIO5vuaWDxgwsmll8g9dPuXcR695CQ4nE5A3/tz9BtU+b5eN1mgYwCe0fA5K7BjIH4VJ/PqlMhl
6E1aSyAs22O2My82ifQSp++kj/+PpZIg6MMtwcVVNGRZ49pIK4xWMJ09NSE95Mdumm/X4LK64/lO
J+ap7gbuQCgh5sAzmlNzSNLHqna+0H+cXBclkyJ1GNL4YIjMSyHNIPBF4yP+ehlX/pgQJuBRSSwe
oWuAat/bpb2TVr9lSKUM22d+mkPOFMQltyO12whPPjsjp9fHsM025JaWnF8e23SvqBF8Lxo5i9rL
fKNCcsvng2cqOWEhcfeboHyrqH0GvakqXze1+E0rwRyXI6n3B7Bp0SNdW1VkDfp63s4MgXZlRZfA
qziHJ2vFVb7JOasx3jfheTrFYS/1UTgJw7aw4BFnCg7zoUQJbpwTk2Tnm8WfmKz30EA4KBzxTKPh
HtyLlPpAkD9o69FLaBY98KK0Ar0uTIIw8N9fs04vHaNFlu5AUp5iBGg9vAlRynFCLM2pnQ4ipEGr
N9jh5oZy+xmyvAT8/tU0WNm7dA5GE0+432Ff0cWgBmDSQxTUUr4HJDO0SufW3ownYEpb8MAAPiES
hfUPgzNFbOizcz9fecQUPCKWbMt76x8ht2VsmYR8nWQvBwQiwUWtIXa8+GuzxBwXGPJ2Rkae9ocf
x8af4MQMXe3Nwdj9zc/f0kG7DQ9f9yQznai2r0tADiOA+1fRxRHLzWegZMt3zz6BH5heksIZ1n1p
jTEnxavOkta0EZEiD+RbpPLATh0SrDaQH9a+8XhdcF9ZfvEGG17M5o0XGg9yWqBvpISFiq1J2TnV
SdhVkN/YLueleoecWXSjFwfFm2Q4/6B/oTB3UxlJcLGxgXwKT3bmMF0hi/rwoe2SHm2BnRjc5V8A
eoQZDcSjLkc2t9rBat4S4C1byYEUVBuuGSQSdt4T75arj/faxeOeGMoD0aqClzKai4ICGABHVkDZ
t3bouCQlj+p0s3aueKvUhMKX0IcAuQzgNDRW91I7mMwi3R3I/b29A06kWqlX3aSMnRlfxCoz3HN1
Km+s7kAF7EAuKP99ofYT7ip8KrzyUDWhkqcwg1Ky6Gq9jPW/9t1pFLlKMpMJMYyVQp2nIxOftiaA
vjEMf/9HqSkyUm2LDuqW1fxo314tCsPqD4k0LXcey/d5dm3LoSVgNU24UabMAPLfSu+3fGKZLFht
2C1lODFwzzUrg4wptg1S8djUbOFR/KN6B/qd2HASfGFkjE96x8WUtbDxnMxZQUkfEK1OPF1t5BQL
1SuuDyA2+Ojvbjp8pK+DCZd8Y5S1T2Ode/y7OklDbTgVkI4jU6QMU1iemnCWzvFC34GK5GDifW3R
Ev/7XTg/LCgSQvWzZyJWSs7FJatCqYkEnBvaGIf/18Dj7IjBCv12DzfUtXE1cJfnKqIZ1DB3kDBI
TI3+cM7SN2rxI6igoo/qB4jHDG0Nyvoc/ylE8ICFFT6CunjclUb6HbWmdqdpkvoFsJMowBIBAiFm
0G2CQ9FvQAErv42H5D5WdbhnSnUx7QJBeHoINN1CRE6yBmRrRQ9TfA62T7waXkUvhCY5OqsbnBsi
gnbH0Vh1fPuxhXGfbRFJxaXnIkPIWRL5TC5DI60vBvhswuJ3xokMX7EttHn2jEFAN1ijRSwOI+ra
GU5fd89s7SmhlnygeBGkVyxnqqmr2Mf2TMkK71g8/HyP0zJ57jCDXqJ8JAuUDILDN6mWNIRLglfI
pCN/CfymAlS9OTqBs6zlQ+sRPX7jF8j0Ox0fYhicimG+jS7Nl613EqzBWZu/1tZlzZUK7MKxYyfx
OjZwuNY44dkGTWPXICQZ7SrbjeiAg3nun+A25AQtdgvMFDJzZM5kAA2Lgn1epXvD6iIYMr2Hc1Sa
jQgHNRSwm5ngYpJu105EJJo4NFbIZ0VePpR/6rm8epQcHSa2kak9UfIaEoBAvJvdTaO/8uJwBEyZ
oKWVcJZmGHR51bCtGLsUD32Gj0PCq3R+uq3mEoQZkWFaX196qClCDbztS2QbtBG+26a9xECfSIEl
jvqiHgxDNUf2YDq3MlQKDl1ZIAnRwY9E10JSbzGDsWNGi9/LLugQRwXVpArd6VeYgKOnL6glMtS8
4bkyzveagPLJ+V6RWXPSLO1N6rQAl4nA8beAOkEy3CrtzEWo+Sp9vLOggbxTazKi/gGzAMO5+y7C
1Wb/cEs5AnNLy9cWlYQWdRxNEhMkZeTkKk0l//0A/KSwmzDv7XHPoGPk/hVe8ydg8jt4lSrn10CL
5dJfjf73h8hVcMyCuaBL/LKlAZ/hX0YgnsNa8jLKjgnJxBt6kNFej5zIYekbjbzu/EGsUgbYUnr1
iFwwWXlNFh6KXJ7n2a6G3xXme83ps39+aYZIU/fHBTLtBS9N1vufnav5kBOw+W8I/T1TQO+GMKi1
MiP68xgYXz1Nj2e0CWlUckoHXXPJYyIDZfpZalriqZZ17ccY8CrLOHcLZaR543SNvNXB8jgyqpsg
CFGuBaBCLbA4+e5qsMYMUO7nPpILgAHMyXDvT3vE1jMEcKPTFTYiE4gKg9RQ+8r+I+9umO/nEC+R
PhwcPuR9/yUESlPR4f9ekV0Vtkt1tqddO225oo1TVPufd35wAwfenDt7dug5LbX+Ch+2lVA7u5rN
C2LVRLyXZAE82aPUKVB+Ufhv/xJveXC0DVlTR30clt1IRr1mF5EGv54w6l2cUuXjVm5WW6rnXr3D
62En9eStDfMN10bfGa8djtZptAta/jya6fn55HY0sDlbQtFH6n3TSu4et4iphIvHLoo2P6NohegG
Hul19DdA/Ij+PzwKcOOkGTKndgbOfWtX4DHHhZc0Mtlo0OzeWQDHSzIsjcy9JvpYTVFiulrA7afJ
C3gkhehyG7xvmUb4VRRLZqaKT69qqisKxphrJrRsJkiXbrhnqrgP3gibaXF5Iec6TBUJyFm71m72
kBZY6UHMI9JtLrvGtoMceimA/AiGIe59BfvmaHgG4k31bgiecZnGTmfvhLQN32WvC8w54FRf3Zoz
vqh+iR01P5TLtuJ+MwCMKHPHqIEkQd1sGEWPi133Ee3olhHfWkNKI2wW5QBP7TITT1MiKPryQvlj
l6jk9zYgdS/eTVzCv9lQTXV5++ntVW3ph6+jcjl6iD4mKDA6k3ptj3jVT7qXuO8UZk8hplNb7QU9
UXKgICef/bvHUDfWh2OS6uprtRc45M2JYzBRwV2x+/Oqj0DN4FY/FY4r4tXKAbGQGkCr1cM59H9h
EbZAubZr76CPq6dzLQZFLYE7iGlnA4ABZcVggKQ5Ck7YHJgO4fgCkiu1cHl/QXj0SL/2SKwDtA2r
tdm0NjDO498/8Q74hYMJfXYZRvnLgAJMtibWmLy8t6EafTDjx2ajAjWQ1biAFXOERPRZPP3AUIfD
EhvosRxWS5Sfm6ymazF7oncvTarrqQO7Iak7izqw/yGYM5iDkk1ynQXc8lf7SLzZV8/pEGfk8Rxi
LqFs2e+nav9WG5MGFcIursNEjVMEXtFBzh2eKnbV33GuSQ7HPGWOtD9lVhcwQw8txacMaHLFclfF
i1z5YyQje7yvJ3x1uVYh9Eolv9blnQ9Zsx/mI4qaMgz5+lA2IAmlxoVigxpjQ/XzjHQfq5Tu3MpT
bUjngyl5BtKUlwZy20AtJn9tDS/xlBowHNUCUYh7Ab7TDWjdxO8sYVyGCnROjI1t9QlPDf9FmaOG
0+dCTrTY95J2qvYqplXx1KKNBR78ROf+OcTcpiz1b/Fp9mZhLqZq/sYfB3QyK60c4ltRllr9gEQm
jVUF9b87G/4l1IJV90SGfQlj0kT9Mm53dHffKirVSoKucLjmxxbZj4D4YRCzMzjLxhdio3Zewjfn
un9n4gFniNiKU61CHyqqTacdwQrlHarAwLXcYxcaHDMYo+jr+bsMgeIQlwtfqUEuOhGWQNWuIDao
9jlDl0vg3y4fzchpos2cClE6bGXGE/FaEvesBjy/Z3Hp10kt44ZhBCwViflzCz/iOHuiJf4mMWOZ
XEjSVL6yhin8diqRQqMZ/xtDWU9aWZN/zwxJvqjMqJcdrjrJEvl+5XBg6b0OQeJ4LDoZbIAaJQqf
2zRc0yilcpoi65uZP1K/XHWvxOTAEVsQ1GOkunzoQgilBCOZjVbqQwAPPiASO3ZPT40WWo/jpAw+
dxiXqv3BoJdgZ9hk7FmUuQr5nNVabzBLrEznca5r745ffWB+JtVthZ44U8kgkof9wrsvriR+FwMy
kGSRA1Kmb2p0OUJZeYntHONf2PKui5fOaMGmE3m3+7tBxItSlVZtUx6qwMFzQIg9lUOGOCCZHcaE
LTq7CMjl4ETxZfN4rWq2ErALpEiSgdslQuJJLevNkxpd8iKpzTaTBMbLxmQiraJYV30m8H9uCrvq
+Quw3FJprfLzG0GoqIWNpGZE6hErirpdzg//mwwcBHnMNJp1lRTsoyjaqHnMD+L3vkpqMGE6AJeI
VuWceRlIvdnu52R/uN1YkLpbI2XZbqP21hEHaed8k/WhIact3a6O0KaX3wF8rvy6m/i8oyClk7sU
3BjIFwgrCGsurJnbko9NorCFZGF7bMc4bH75/O95IvDcMURF5a1XnRGtt5xbAyBlWt10vRi0HxIG
wYktcR+XoewWGUx1GiOyyAWAyEOvDDE37et38dt0fOLKCYCzmdUUfvHyE88bSfajgQH2L4BAYfgy
aKE3zGmbQivzFNStMa4Cu6uxiPqrOQYg+kIBVFcyUKiD8wErV1HgSbhxOXv4HYwjEllRTmzizN0O
9D50uBaOnm0deX1p3OfDyyUXLtG4+W1Bj7tTv0FMUpOpGyUYahhvXWQhOBivC0M1EdIRDZWZvwh1
h5qSHE1g3fJK6vhISUEBxV+Xlu+NrZlNfoAOk9DwloJRj1IwPXtsMLq0sakVuMLGBmLCm6FSkNHX
QkHbJTovDbKyKlUoS7hp/oBnonUQQ3LIWK7Di3CgAqnp5zqnNXf/M+8UuIRnWea13mhhzYBQkYnx
PI0/CQJgCKnfoNk5BILHWzzPKqbkBBuz1JyzposMEeUVxVwPuwWKC6B4Y/pk6+M1BmUM9YY0T7I/
9fysog8PTkhuf388+2L+xntvWrGvYWM7xdeXBDf7BXX9iOGq8cmSFkEIjB/2/wj2iI65m0FPvNcZ
jDw95w1H/k281Unl1aupiS36EQkxLbYKtTehTJDHyvJZy/p31ZyClGDUsVroVf5L2LBHkuucjGUt
lbych7cfOfpPsDfjf+3EQ5tnhWlpCjnFiRSLruXCdlRdB8F9LnJ2b/cKplBXJvC10cHF3c32hMQS
kVGN0QS99VgDAgrfrf1Ni4YXPlSvDGnDRYWtqd3NHgSUoyhKxA0LA6jbyVAEHcz6qmiBdNjkLaV5
FjewtgMKVrvdhipUyGXaCgEeTtfVBuACeUTdeqAoLJqZVmraKrWvYpr/fGJk3qKsLLpGVUI7H5UD
UKEzEJNYUro1kiniwH9MDRekqPw8aX8/vjmj4ufvTNXTrmQHm2be1bEHyH1XpInZEDkjjt9VhNgi
O47p9l4xutXRLFtq3YKKfQqsqf0tfk8j9/77kZPiZpSCeMmEZrqpUiZFSdibI8uCfhY90d32MnXl
nCO1kwVrTfZz33gTxeLhIgAnHwkwrAEtur7dIBojowcB8H160tIt9SxOG89K/AygL9+ui9SaEdOo
WcL9WdYEtbiMdxRVrg/JQr+epYWZ2/d1DRi3U3Of8S+fFhImNJ3uQCcZUOQIpTYl40MhHdtq2OTw
PAEu99W2XGZrdMJx+DBBV/WHwaZmucj3IY1FusB3/j7sA6EifQtJFFHDCPEhCJYnPDIQK++V+Ntk
Mex5lTsrpdYbqA0QG7oJEep1kmMMCbD1RiwdNaWHnFBCFwxgMFXSHCzuuBMSJ843Dbzm5U6boG4N
1/Vzyc5kp8jAT+aTTk4+oi2cUnwpszlsMnVzM385XxrLlgjMSwMe/mBe19ir6/109n+zB17fj5RG
livJL7CQ4wAPBSxYwCkSAALyqiA/a4SP4EkHe7x4Pc/49Cm1XNwhwBMux8u9zQ/VKQjoQnOXWjM5
tFmb1tXEO0u1BakETBeb6G+i+xcJVnpkufUyN/epN/sSCAzKBtDbj2CtiQ39X9VtHcC7lyb8PLUp
rLfJ1yKaoic7lEUU0Msb2oDrFbGaJjwxw7Z57g/qA5T73YpqeXK8eTCAnfmECEQGhUmA+b0gozjx
0blOSPavMmt70coyG6IXO+eleVl7T4fRUScfTJp1G/b/S1WVF5n7sdoJZy2JQvvm74xKoFKSKzrf
dtXuCF6fSIOPOCsQ+MZJylU6epxCUi9Y1HhhJzIRoYPqTMnTc5OOkKJpu51NOZSn16RzjD0dtKAO
elJSRJ6tCGpwrRD9r4YaPTMIbYf0ZaBe/skg9SUJ2E8up58m4Cob8TbvnM0jWcUAS+2LM1HL/FRC
tnd7Mx4xZ/7oVgE6xSjaXLvB/DVtTszdKoIPemoHZI7f/lP38C8iMDrDqnMZA6MAJRpGifkvjsHi
HJq5tQPagwQUiIP2wZ3mRonjkTUFnX/NE4DSnzrw7++X1Ki2eLwPRQ661/TcI4UUyYcTuO8r+IMl
22vmb8N7y8adpH/gAPzjKyGWvcFJXjF21DOy5Qjy5WpTYeq6X1qSNANpJHALwbA0aiF6/NalLht8
BIr9wjnXvvqoeiMJhcNGlLBsvbu+dLi6I1ZU526PsR4CGqQIXzJnRbB0rVnHQAxa3sa1ejW+KtCN
RCKGRlQqGSYfIbSlVh/KDLG0ulWjvSmUvxJr3t/QOxEC2rAlZ7xAnEjfieD5Lx2+0CYSVx3wgYT6
gu/Y43JikKTyBSQa/titj40jrH3U+6QImAVVHImlUlqVgMnfsolmnVMq2iYbCG/oGlB9N3A7bUFe
rUNgVQRKYvkIdv6Kaj6eVSerZyiCOup0ncAQfseJCca27uI0tQp/65XN0Ot8g4jpkC70+NzBPukj
abVavgEIFIU2gkLDuRz/FsYVzFKszZ/Hg5GFvbXfrROx7JkSsVlw6v7ioSeIbtGvXYbxDRfYY2tM
o8kxV3zpa5NiC3qMYds0iVZvpVm7i+zlbh+EimyNQl5tcQRpF33qS7Sy2wLKDYY0JenuYiXQle4v
6nFs68k1r1H+3SArVkh7QjIeO7NYk5EBnRJJ979SQU5wKIIWj6ZEI8GNlMbh9XTLIH9oE+rsaoRk
izJtyl7c8S/7p7A6WjEkkeC1qH1L4wY9dp8M+qAeyyAcobQfdcl0ormWwOu0MdTvUvQUd9Udm5mk
tJ43tlW7Ha0TbNIemIixS4ClE1elCPZMjOMKKMamZWl3g6EfW/JNxJp9snR9VDmdHhapVf6bBadm
DFEDD+HbyXUo3CsRRsjhPIF5W0R7844vuSGYe/qrB7fi8ZDL0IASrS/193tRnAw2vHNKDae1YGfr
LlcnZxOFaGwJoOUgmrYRW8Lu2GoX6VQst5DkBG/DFN+tm9Rc4syF7kHy4PT7XMDj2vPVnqhQR1la
Ypv8YnefJhdtXRhO7BWGMEFp1TzobMcf3Lo+I7p5P0BVGR0uWxOyDkwSk8sCK1q6OR5CSnG4soOf
BWikP+cykGE/A8WGV1t50C2FMhKQUZ+TKv6AN+7uS7we8SRKdzr/dGDlsfFTYB0fmxL0SdMP8AAC
j0SI9ZYSkWdwtFIbfo/Hq9AWcQTK+P+Tm+8SukgAoLm0jg2gJPiN9xyrYN8qTYtgqSwd9T/e290t
4rZgR4AalaeNUBqAYprm031fadE1LGS+NoGm7dO5LHccjIXkhuOOmw05lP5q2zZNCHHE/p7vyzYv
ZqJ7DfL9ziqf9W5nQavym/c/w+K7KsjWDbdzO4AAuh+FOuaSrW4mOoUwYhzeUGpRPaqYZ/OMH2a4
ZbIYtR/cI2lqoieWS4pdP2GY/KtmbU5SNQDjD2dzCd4OAWOg/HadUWbKBP2Ed5L3nyC0Ia4jOsLZ
OvQSUlDWtv9Z9yTTtm9W7RnZTVOrk30kCYdXbBjl0DYIPBsGiAT4/lpRbj6tSgoS86gQwnDCLEVw
sk4NeW9HcQ+MElvFXfMychRyvihkUFBIPGJDSQn04oDQznqflWbLzlPn4kcmPgZzqjjRsksLN7gD
scZd/gGDRGPy9FuxbkXq8s6+/DrNOWP1kz6g2bpHRInIohdzo7kL9CxM8PvVhI+CHQ695HdA6sai
uhWWdC6JTuLwo+M+67kojauLTAWWG2Boy5tCQmoU3n9qUjlvb0/EhqLhzSPKUy+fmw6T9u35r+j4
gb3k32OJAgHkSEmFXNxsC6Eh+QKRwrNbwEN047VeKQjvJ00vb1H3F2maVXNOewxjMScCuq7y33aJ
uEGdLdQAINgrecTcez3kFv6xq58CV2gZsyQxbs8/hrxZl25ppfVos20nv87KTuw3yHcfjGHYMEmA
oMiyAkuKAWHE5EUh1GIVdxT9mPVL1zKmizNrxo7Osrwm0V2yHuubwxgmYfrpHzOxlbr4bCTye9ma
2TMZs1/I16J8ZcV4cUvDSQOTvILZBuDm2mk2a4QUnSC2b9keCZ9E4r5flgiHp5Mzw9ruu3vY3u2d
0IfYwbcEZnoK4666RapQ33Y4y1JlK7geLovY2T8HZoXSCsm9vkxraMzprIegO8uT4I4cUmqN50/f
cgrHCi6j1t7dPNJQClN1nRMsSqtfxQ/ADAKRl9sInPZyFbXWl7nrl39akrSMBV1kHbL38m/AVAL7
VCXooLUZO7d9GiVGTw+eK8VtWVD6WRD7/DDvOTELSUoyj1kcJO94c0vaMtf9lFgWv7CV/qcJW/pj
SDyBl248aRg7um+9QmP6jPR67SQZwn2afLUQb2c13PgvpHRsblT7y+nWOWZLVc9Eh5LlCmiDYDG2
Y6aiwiRHkxUsrsAPQdwgKBMCqUhmyLNds85rRVOql9TT6R9msnfiS1dIIi8pgH0mfksro0rFruWN
LYXsSoJoTdLATaFgsGc+F4jXKXGbm9Fwi9lX7JdFTzHmPnYfkTVbmQjXVMrLEvKGPfV3vR4Y2tB0
eWmgyBe9T7Iw8uNQuQIUQW+6Djt5F90I5HL9V/szh07XQjWx8Emdm87AVPNZMXSekQjXkjTtPCnt
FENe9ePtUWJdPs4/OfluklxLKvDFk060xqDlM9spq2Qrvv6WjgLdSMLBuf36i0gaovyt0h4m+8JV
Fx7eDCVO/F+2TQpI3Vb5GhrxyoZ2GkgxF9dDnlJNpM24NxMgU7lwj6MoavOmTHOrDQ0lD3wlLAdA
6Mxy+bJ2pgLyZA2fVIZzVit4H+qKQomK7VvxYew5+DTzWpHkT0skteSICtuLeRYPC4C6nMsuC1Mb
hY8sNrfsPAnS6g6RcyBFFJwW+ahcOh8Ynbd1wAFdw5IbkeuHvS2Hw8o7RI3Gq2qBv4kMHvHz2zdo
gMW+xaJBerhFDp/2HpyWwVtFUP/mWwhbHjKitIPg/NrwmmJMQq5nsgAQ8MW0YwBUA0izTYp/25eq
t67Iv72pmPnSPGXgIipzMuoBGJ6dIdiSGYnO/8p2+ftWNawrvyfuXmyRdb8ygNtgnFeyKfGiXJNS
71Hu778+KpaAJHzoFdLtp3HJ2i2ARavdsIeiPwsHSNxBr4XdzrtzM8vSrVEt7+pxwCqO3Y+ZM7Ht
5lpjqvrzHgpW3PrGQW+vx8wdwH+Jc9H+6lFeuYtfQXNMHQUz/WMhacfHHI5ZLUdp7R+VaojSBDNv
KoFo/tZb48WBo/WcnpcMK5fjGpeGwGts9wRXZZNBqoP3EaJpmR6BJ7UHH4VdMBC2rp/pslJH0h6k
yRw92bq5C+n01fb7nU0255mbF8UlEIqnlzj+01CRDUMEXeZMwCsfXnL6rhqwtZi/sS808eYC/5SH
wimQOEh42+Mcao2yFbXSpA03JGfwVdCL55Is7+Bks2rQRcyWa64je/yP/Z/MA8vPJKgrGFIZbN8Q
y+RvHWNstbMa5M0ZTDsSLBE1EY/BfUrrgi/VxeoXdcHbNOvIAYS+f7zw2ZxYz50rB7YUMbaNVCeT
YdJWMrnPFe1wVbagHJPeD6OwzaC5CBG6I6R7BSB5k204L0HJCFShhxxxR4Gpcr5FmeUOFyrCmou5
yZbt9H3lyKiihg24mDI9yEpwi0VAia2N2GXlXSVD0vAzrBtZooBLPOqZykzT0jj5uixvMLkPg1WJ
kgOZ1NeGZvmKDRKAJagWhKvUpieRS50PXSlHv08ZjUqD1LBmAvXXZL8Bg33ezDtaNrBt8Fdrhod3
r9yw4QL22PXTjQSpA/DjjX5Plj9KYO48WX89KdEy2Mg6O+fN/AEr6n3/2/nuzT4AKxeJ4to6TG+t
jvTwOMMEi00qJsbIHXZIUWa0KAz9/B8qNFoFY9SlcggaYVsTKeogWT53d74ebxE7GU3IBbM02RVG
ey3rVe0ZBFdLCk5hBxuSY/zEbqMEv8ToXSmdRIOoNlwyd3HiuSARCaV+/p/ljBqOMSYQ3W2Hcm4c
G0grp45zbZujmza4XyligB9EHQYi2re3MpX69wqjAscC1bsKaUwDSPsso4/UOexiNaol1emoqdRr
QuCHnnuVUeB2qWvbku2BKxBqB66W/iIIIL8JjW+yTT2iebfoz7IxSYNcgtrubJFGA6eyeMw4Kc05
+WuZ3XKG7OeXUgIUL5zuLMK1bDMxeCKDmRXfI+Jx7nNxr0w5cRbmVv71ng3FdJwWpM1eZwAihsrv
Rph/Tu++PBvgS3RaF/JJOoqZ78nhmLybGQkkR9TeRv/3/LgMcr3Xoin22836u8Po5ZAVbYYvco01
xaHIj9aYMpg6cRnXMpGoo1GzyE+82rC40ThFjy5/c52HutUQnSQPvJomr9Zf6tVwpql/uxw4p8z1
Oo2Fc9HRW3dDQYpS3bRJs2kJftnsEfacX5GPiUpxvUYBx+n4wpApFLoKW/tQbhBLEevUE+lqgwkj
NgBFuwIxGXFKodSJdD6pFwU3F5udz/Rh0wws0l+CLrKJWd7vTboEI0VG46iv7aMk5biZG3Frc6Uq
5DH7w/D84ap8K6rs/UF9d9Wy+U85dyq6+iczMmhx1zdg2TkBb9twH/t/vRaeyikI949vPMVWTgbk
wC7jQmSgyppz5jqLp5+lRPMWO3fAiHfOm5yD80pMaut/kxMQ+Ad/9zCsP+5HiJcUnPdstxYK3mSS
8CyEYcLtm/cwATWuaT5Jd3QHZb5mA6wb2+l7PSvETNyV4OlFvPP/tffpS/2dZJdBiQssfv3hKEmD
ae/ZiNaiwh9Da5mjwUiqLnKyMPzDx3b4zD1mURw6CcHl/Q4hm4xnt1qEXpzrN1dHgQuCxveXm7NZ
6OWrqanjH3dAXHztww989fakAIoqfShBs/Yus/5NhIRlRGNSNN0k6k2KBtKyC+aYcDEs/wUsOuUf
EOWFvA2X0d8Xw1AtmFQLICp+rOm6AwiOVEv81umC+oJpWhFbhSoLqFogUzGTFEMKnsHe1bIgofzd
O7DLCW62A+90AsW7mOW49iWov93vvjB9myIuzi0O31fyI5mPs/56uOR8Rdl2H1QzLPoQDrNiccvs
8WQe7HtCr7lxyZxgdzUi25wVy9c0W6HnHHd92GS/PrtWUPEBGH1Zyt+2UWArlPm9hCI2lDP061oV
wFfK3Rblz6+nKbbFFdYnir8oZg5HWPSSpWA6Ub9MVRM4MGrf27aAiXk6MhiCyFJr+TOzuIlIe/WE
97XYA0KlVVeP5iiqdjtFH0jHMn4Ogx4EeGIA5+Alhl2ZtTBGl6ihJX2f7qTq3Rg/DSyU50NO4LJ4
FUUCxUAZ/ZZMW9lJP9t3YqPunRQkBme5l04X06IUPeQX5DfPCTMpsMHTE+MjQiP8REFhdc8Ahvta
ciNgIHFLMawCrQFrjChZ6aYbT3JNy1LE+mvpitmNMp6lxlIZSB7pkWjXfzgMj82kyQG348wVbeto
5HNDYoXua2CwvyuGRn+f4p+X4nUBaFLVgXqr8x78zyP6kVpnSsd7Uy3W3bIMcDvfxsGZTHh9BQhx
Qg1pXGNuKQ/lhHGExNZbMbX8Je1HrtXxDBl46nrsWdRH7/4pUsDf8qkIbgBbXMHwjdRnrvJAp+QL
TkdyEo5T1qilsZHSwPi6guq7WUZsumfcy7YAStFItyCJJRxttq+QhBofHwZjsEUdPnQJKVlfShP8
FfPICJ1sdfklxmX/wf5TuBZGor1IGigM1+nZrxWypNrLsKtwEobrwcgW78rIRCnF0qk3znSfBdW4
RKcmTJXDkMK1ZzACA5pkwzq8//nYkwssSxivVX7rvxer2NrMQl9Xml7lhQ8rO6l49lSj5CGvJeE7
G0xrPm7ihdmv+Q0p9gGtJ/vENTNNYlunoGdbQLpFPDCnP/EmphyjR0lSn9o6Bvwyxa2BKFuv3aDp
DG48r4vWwo38aLAWhLqGdSIm6ksHX8z5rWPLvapnCiyvtr5hhK6F2HraHDaGIwfXfzyJUMtJ7p81
a3n4zUh+EOa7HD7a/6jlVuAFoJdWX7xqk/9xseblRFex1Gq+zEiAfANFesCILb4OEUTLgNQ8lF8K
ydPmNo3WZR+a5Kzb1g3LtBuy37dtHF6t/88Tz5ocyuJZE0e9OJFTGukYm1tbY4i3iDR2Zvx4ZaiX
rH/avLUbUX+hDu+4AUioAMtHyqtN7GlxOSHX7Mepl3JJolGvmj2yCqHVCbBAFanV1mJAKOVjAK4l
k1moMyNDKCVPjJPHZouzrgcSvZm+kg4QM7HxbPwxpTDFRjU6clfe65QeDSwMXmK9G1dO68INC+kf
e43RAdNGUq9DNpC9xihglmFjq6fTOLmdaOf0FVrS6YeroQPs4jlmQpcrKdF8RUAJ5TZNH4K5FFGp
wEtEbWI4cd/J55pgRt91Pw5F134DDTgAE9v1eYkojADEYKBelIoqF5s+Jyr9gnNd0nUS8U7LHyjD
lYR2WMXuoepMpsoNaAT4z/HjOpSNd2t+raE18/rmw3XAlZ0bDDFs/CTg8zZeuGq6Dm7G7PBktMe1
u4TocIdwdxRu58jHy2Gyt4sj1Hf9gbqPshPryV3/VA+FPqxykzpJ9zXKAgNFW0wTeVCxsjkkyplS
2bfyrRjDAYDTGO/riu7iq4UYbAhGzHEGWqVjgsdfVrpfvJwsl4Ov/hrh5b1GQHq59csd6nTju5yN
rN17M9L+2cOpuZUCrnqrTGf8k6gbmpAkT0K8U5uHojyTZe3pcVb/HciqNh1xHxyNP5h2Vh72zrIV
lLCA3hlZ5m4Bq3a15VvLYi/SVFPFTbLn5iLmNyVRS5NKMKh5sOKNqWVCTdHlkzYJiSocry6Tvpmk
66LZIj03VPYGXUiHlz6E8yUs3TtMlrsUfoxTQb8MCOEPUu4xgvOhx/5qO/tGXrh0WIsX8BivWi4u
I/vBB7I4168yqj6TNbTd83QSrG2hC3p7t45IeMD+nnn8l2hLE8Q438HVWQMw1x+TXQoJnMvxDKkV
J2az5o7+sK00pfk0Vid6ylx9rqR6+6MqwAUvy62R5KitiYL6g32ZysjANCrJhkpuoFZdnofX+Vnp
t6TG5veNuS6BgwNQoTrJG+HMKC+QCtEuvPcmZ4JCBkBX/cFqZ8GG+j/EOJjoiYuYMih8W/Ihj/o4
gyI9G3dB8eYP0dFteqAGN/ot+FDzGgXUmU4+MpDBghR6WQkxbGX72s/cAAalwVfdCwS5RenFz86B
jDD7gZLTIVXfdmTA/9v9k5AdOWCGLMVhUDBfwOraR7ZSCB5TDvLCX68W+/7ZUS6sI9uUsoI+XUeB
Hi9nRfE3N964Z00mRx6gII0YUbPINS0dZpU6BP9sXsg69iuOHfURLVPtgR6YxaIie8oEhrfw+BbH
ywbWqfdH8EyM40/zuzabuThUHf0PQ/s06ZbtG61htqC3r6MgTTSKYXgSS4xs2fZqVGnXJQTtiySS
Km6huOIjGFuNdpdn+49gSL3ir+M/ZW5lUOkwnnQIph2/R2Dw52uQ0dwpc5p/VXchvcCyXT48v3pk
XKPO4GU0E/O3IoQK8PgD4PMoICMcdbhpmsZchtYa55raPSvJ+hKPjHXltd3+0CRaiygY9/xbgTPW
kBANy1eW+M/2kRfAmS1NLXXDBrw0VWS6xV3dTJDdS2CLW2HWjJjcwGo09KuP8uisVpvBdGw+Mt23
Wf+fz7lmdrCgWm1xG0GoiOsotdq0+X8gyf0q5ij+MjsJq8h4SO1fRGiuRoTFYWnrXyvAUApgWyr0
zB3DGwdqHuorhzKf4lmNGFw2tLVo7lCZYr7WpwOqQGLhodTPZ1dt0y25DlbsNN8djjlqjgTUfgEN
tuBL0IHd07ZDZG8aQwxET6cK96hE65LP5tCuvoOCAtNxHXatJD46t+QpPSxqliQZLoX7yfmc9fwV
kkvWO+g1i9N5ZwzYvy9ZxoJJXKTL5SrDWyc+9IRbh8Cm5p+tzu6d83z6gUcTXTixks7EIzv6Uh+o
3X8yCKVXdgFWRM/XQ8nuD5ZYBifjOly5ROEVFA3AjdndDXZqbfBReKfQgitb6GEUE8Vvq/ptLmcv
vdFpGV2AQTF/FguYXTTgr4svsDaQoTbdFKESuTCo+lRD4AT6Qr1Ga76uE3Td8+YtziAsLdL24sxT
K1DXJgawt9NAiqRWsnW4EcqNk3//W3Q7Fbxk2QvAcmQF6l8YOIalxExXF3esjVT3Ng4hSmU3U8pS
4qy7lNgy3+BWfRLwj7eqVMAeTPazHAwmeiKdTHmlOAORyXkPu6vGI5U+8Cd9SVnewxUWXxOJ+/9b
cbjrqs5cux2AOrZVZ5bICegNPMTSwAmWNDDfTkz0Qzi/0PEfDwiIHYXilSko6K5C4+b7d0x1HVf2
XhoruKaxPxTWvuyg39cK35RPEeMtezjxYOhE3wHs/19qAogF4ZLSxth/fyxlRd/B4CcIqWEw1oTq
5yZpOh02miMiHQ2zSN8TW/SjVKaF1l/5Eg6zrsg+B8eMqHMLofERsge7o0kPIP9PjbOTXp5FbL3H
JAIlCYsTWwokfbGux90PtoEXdjqY1/0J5HTfHyzQylCuCPFXxpYqmS8kUG0Vjq+wD5LEMm4Kt2Z+
nM+Qfd1lMIJ+GQ5ReEGGRaI5fd2dlJEuGPLIxMOcunQl95QU9DIMukWKS0+AvV0efCAo8SfmiFDC
d0duQtTc6MBtS8CC7FH1WqAvag+dF1RxbzESGgDXZ0G/+6EZyMhadyqYFePQoa1Nvi6Ja8upVG41
LORKSFtkzwhhpEdV/MlAIzlyXvijoEhHwNI/1nhomOsbiS63fZBIGXFsM3Ns/rh8m0q0Yn6ip1fa
9UvP+0pEzbyf65fZVe9Mh/s1YoFd1W1vsVYxVnf5kEpbU1P2iV23oYGjXVGnz8ajIRqU1pdrsLfP
/gIvQYwLaRiqsFXeT60EtO0jDONN9bqBG22264LozSVt/nMKxJN15yBioI25nfq+omj0WBLwAcaz
ygAXnrtHQ0jElA7HxyS7tfeNTBkum9VkCggFcyQuqTr2USG1ry9eYQhkQNvXrnj4PEvJnAJShie3
qKgvoCIcRJuaYI5MogM6JkWpt0mSgHp7ubQehikRMCkeOGDiGiZ5nv4Yj51JyDcWomCox220Z1oW
RNEiW3+Jw3CVpXTEGrWwJeDyKzhXBTauzbmsxPfW9A3K0r7JjTLOT3W8C9IwN8QC4zAzHyjQJ7DN
iLj3A1CKFBQTgsbf0U8J+Yk/jrdycp+J/wErUlCGuFTnM/MZ+j48lE6psiAFLN2IzmQjny/m/mff
TDbhMM3grPjHQEmFFlPt3DjskUCPBMkxNgk8RGMAyb/LvRElOtjbp5YKXMm+/Cz27O+6BaXiWMIO
1W/5BXoV5lJJjJNOdiUM3mftXnMT3UyXDOAPjl/jzdkzLJIbKZcEAu+bVBVmucvji4jnEeKyPfSq
/naW7CUzZqEYBhJZ33hXLAL99a4CDpEiSsnz7a4QmPWs1ahb2FZKHpkGw0IB2bIkqSj0SOVWa2ZV
vSqdjUte8Lwg+mY2VtEyico6PwCRfgnKWBHcOWtuXShk8w1MZLwLSh+x/859IorQiHyO33Z2jOU9
5NK0p/iDtT4MZ7yt1icbGNR3G+v4RHWrJYlwJQqoc4Prcn6hvAYLa/M/lVVPi3X9xJOocYDg6F3K
nnmuHZDdRfxfwXvsqW4OGmiQhp2YdbMH049eFgwjhUzute6oRr9NIWl5O1WFf7qk2iwIppLaPGiA
8h6v5hlwYwLs09BGaYxtjbmSOUCPVHMn2DlmKn/r1mXe7W1p+7FmJdpjCNwjE0Y7a/oegUgXEIcB
qxGaLsz8CK77GmWomIX8NOy+XA2K3BoxaE/ZtRD4fxTBvRM0DsALV8K+AWvhfW4odJFWMteGSP3V
kRNy5vkly+NI8Vs/wrEkhlGb4AfTi0w0kgaVaN+Gb0DPpJh574ihjnmTRoy9kn7MSfgK9sAJhKR+
dVVvppVOnQLFtu7T2cMUipD3rR86RAr5raKNfca1gtdm4IpMpGzRbyBvtDBkRckGhY4KhH1xjE4T
nbaTlIh8PWf+o99YCnYH+tt5edyRx3whAMHLoC2icUmJouJ9NMKCZnOR8P6Y2JHLrMF1zzdvNMVi
GPbut35IxdFglzufiWWS4csGp9U1ArOX7r1D+RCXG9gmKZORwWl/jkaEZkXw0/IU0wwu5vpq6Y/6
C9IsiuJEpUa41pll9DMZy9Ce4/zxPDdbKntGzX2//aPQRgCfWS7CF5wyZ69QG5PrGrWjTaNbiMAK
8BZXBhT6CFck2K2t3teM5T9syHQCwK9mDAVoj9QNVUQ3RV0Yfdr4VKndiijb9Cwf9zmY02363XlC
1UWMORbqwX7dtmbnllHYzrAoMe1C3Tlb7G6CsY5S6WUx+7cqUJIlh+OHEhvlwlFe030j+7Fdqznn
ZxvSGaNCvT0I0ehC2GdcuMFgdAYwPhO2k8JFn6jt6djiOv4rI0TkirUE2Cp5wwloHBKOlzanMqfJ
JxpYIvtfDgpuuHhvWR9A+a8wlyLv791Q2VyX83rFeqHThfFljziV0iQOp5R6dRxpH6Oe1KYbrzfW
Ga/h0cwbyXwF5KVcRkivhCltoVgRuUdKteKKiQdEALdaYssuKDrFqP/O4m9MdWJCsCezPYKYnS+J
DK6NvlBFT4aEmWY0V0L2G1/tPvOToPjMoS6JM3eo+YP2CG5h9yrPETBWkAlPT5+K4tk7418oBUqh
l0+VVqfXF9mglBmv7C+0p2rAdfol8uVYENOGQqpeeVDHMORSu39964thC+8HG0Q/pX71THd9+Czv
WynkReHXySmyo7+NLlUSNmAl9uQt3qmV23NhRoQ9nzUOW3Bjd9l7ztNN1wK7WgW7Leklmccdbw6C
FMxHtoB8MrdN+gGl0BaA6/Hr3A/elnQdFJ0F+P9N1LeSUr/Rr0v14FA5ueCK/lZVhpLv3wUXElGT
vfkLoOTfGy7TDtk2VLTlhe1JFki6GGCRD/aHWwkDug5ZTYqZpE5UfOWdnAuB0C8Yqhuc9idquuAu
8HhToJAx19xwJCPndIYtJos7MJNKvJS6ryxg15aGQwsJvCr2wQh3p5Q5v8FZiPWTYvEKOu+29ofD
tF+KhXDBhilAu3zrmN7HV0512O+QELi+JLD3N9azWTlkA3HVQechbmv/Jv2/tKyqHfOOqcYlqESl
NAy06lfcnk6z04OCjMDz+rDMF3aFjb4w0MzZe5rZayetfkGW7EUUPHcC5p+/0ZPcRuBPpmoqOFag
r3rsODzmxjBoFBAFNgH06kMndvkH7xN6l7PixWVkdBMjKhVxSR41DgmNXIxZnGVb7R1EkS3cvA5l
OTCH+L0SXzkPqKH7k3XslfkD3SOyfldKVCKW1CHgsu+9jVYf+aITRY4l0AFLIa5hAYf1OKPd5YgD
DvaVtU3vum2Swtk+qys2Dwl2Fd/pHLNQgeZK5+62SQPiiFCEY2jCeVU0RnG991IVcSfGrGbqBgcb
oCy4U0WwpbehyVCJNF103W8VNcnfsR16ChYkVFUpsAs7tIhLa32AsoH8dSckU3r3noqWYBQBd2rL
16ycU57bJ/PYh04a5tKr/8J9yrMk37ybM767KCDUKVMbvKmPwvQ4XdjUR3QAoc9grsk7nCEG6OA7
vtuxRQuhwN/ynY5gPxRpufWiLA/X6TQ/xqy/4eHxTsd+oHNAngWQIq3sf9FiWGyzR986aO3RHNO0
6H4XIiKeEPCp/SR+DfJk5r/DeniULpgXb7bEVTor1/h4VBis31gehfjRszt3gK+sCuwUwvicHEcl
flSX/4iXCiJKne2zPxQO5NQ48g5rSF9gfToAtU5vQnW9ygGFrGwAVzjSSFyjm2birDKyEljUUBWG
KW3jCgSiFGPF+Ia8pyVYLXtkpImb7lScMddeee6V2Uiu48i4Bzyr42wRo+5cesdidyfArIP/ebfB
etwphzpicZm5vB7cfzFnSPcnZzGoxRu3YCbC9pdXYERsMGT4Nk/xt++8GH4is4UNlY1YxJH6VoHv
J/Yfj0sYj0935iv44HQsjlpioh7Bhehm2eM9zLS7H2dfHSZOFkNHAZHhvJ+6jd9lMotOnyiCft92
5fwL4USRudNimwZ4J9jp3o+0GLWM6DS8vAzccHdvrUulYH35foXvfzj8+EPd4ao57e/i6PFWIrPL
tZU6KfQhtUVlvCQ/F6XuaviQy37YwJuGPOromMH0B5ryTwy/BpJtsWWmoGeylJjGljd2clzZQTWx
VPCo2bWwDs33XOhT1xzg/XuCogIpBSZmpqr2SK94w54+4N5MlOh6McC69RNpqSNSJTo+JGFIWVok
oheBVe0Mvrk6TQcph9I6uVXzinDcGu2GIVAoIAGk4tYA4veRTvWBBaSS/et59PZENJYhXLsQdUUl
Yr1Dhdu6bPFgbOWfS6VwpbzsUGyG9zf9NlPDi7ZKQrthgcY5xNHi9RpBvnQtLWfQjV1J+BnohNa4
QJXxK6b53fu47a68i8GzDNRK1fdmIuC2iRZDCAwwJOthdC5qHfFhiL5KHsrLzgDL5KlYBvz7WyUM
0sTaQNBPHXUzeh/ouSfEdquBYjm9q44ohrlQx/7TnBQvjgvEH10Lt8hVDxWPfc5ilzuq9jAv/xQM
7oETYfM1jfGEL59LfgY5mvf8l/GAGtVbIoGKOhpw1nX3Yhsr42AeVk2+aPzYlOLsfIrNMuydAlGY
SOFahXHsihuKc943r1NZutJPHjkWhKDfQV5K5vsUleIMMAEhSWfg2Ri3vc/tJSI/qFotow5oKokQ
R6l56zDyEkNlkkZLuYP14KK8Li8LBgMcoB3TckqaoGJVz7QJFf0Fsm39gYJ3w7L8fF1MA3bMAKSi
GVqXYISLvMyV3ZwZ6Dp/ZTxJxk1ckJoe/pI/hLfHb7gJh0/9SzRDtHxHsJwPGhTXFAnTPVQduDqA
Eom3xGmv+5ailK22clj1rJNFLrb/5hT1EleBIDW+59hVxEJfuHUinZMKyMsTME9IwjEIxclRrhcX
diYdMvUUrrCGGZ2e7eJwFz7vgeX2N1jRlyh3Ye94K+GhxzDhOEfj4dvXKuZ52zn0LmjwtK24kT9f
W2WSvCANpUv5QlM2scvA6KYNQHpWpF1ej80RFwOGrnlGow8izuiwanXkUfdB1wQl2ZCE1KfwdiCQ
snlPiGAgvEkF7P8avOK2trCisXD/AqymgrRaqvNr9oYdWIGxw54vG4dsOqwzjsb4eeyQZwjmfXQW
IpjKLPNRZhxG3i9gGFIJolM71kUFTdK4gtZxANelx1VNUWXXHHxMWsOv9k3RWss4rzac7ow9Xuzb
RDID7oXR7HYF5qHUk+3qMG5ITkmRGzwkEgJ92MuJ1V8DJfCwgvlZENZv/aAQasbPT4mdNhcB7ZvS
Nojm0lIwEUJTlZ8aEvZx58dEXlBq58X/u27zIvTid/nf/hnt8yrvpe9wZHIGQQBgnHiUAuxsDVMU
IS9rC0oFWgmXopIe1ZmN1kvF//b2fdmahbE7j/FG8DIncnX1iXXV/mappMWDl4RHcQOS5Us3hxrB
Rkra4qyHeCgdNFoAVsYNt7p9K4FeZ9O98ii5Wk3K+E9yqquWANAVT7f85Uqv7wcYLKMCiA2TuN73
QcONAUdd9gQjG47XYMVwef4jf4K0wyTi0Kbcg6/iQksiRc5+qSjvpWbmb78/Z+R57tT72xVLbvKi
2IQvJwE0J0uacoQFL+HfJYqG4rjdEtfLxTqYV5LeelNOX4yoRG7rmn3iY2K7XM7WBeaC95TSpfYx
k3x5fZw2oaQ72ROUUP0SRpq/0Ulwnbs/hmRy4jjwhuhak1tLlDuTOv6HtCZdvMizXr6A3hvWR2Zc
kTGt5j2T/p1QrSHkANi1RkdyNJ0MRoCR/uvF4bkZW/V3b8L1HXuO6Yy0qNZZ2b5PBNaC1My1SSgt
e4vTk/F19A3qHeEhm6w//H5mMrcrBBuLsepRmQjgJnAMrgjaexr2S1NHxd+/b1AUPJx0lbVVs6qx
G0d2wuOrEW2J+fyiGl4sRdFCZBaOpDXa5QAYsmFwptLcO2QpkouhjjqFrZs96MHWkj3kebOtjKS0
rFoC3ocvilrktRsm/fIQOMohDSbXDjSadsk6GAuh1oJYlonWEqtbPSBqB8xP1zy9KxYObrGKBk0m
8tTOwtiKt1OsSkFnz9X6HbAIkg+gUFe+gJkT7aNe6iFO8gh9sZigvY7EYC5iwvWQV69Gnu2vmNON
8fS/Crs9Jcawp9LdpW1srcUS6NqA4Oe9eSGdfGXChiauAZnxOoy1Sy5cjy61x+EUpklQoFLI409e
K3k6olx3eTFE9zEFp9I3AX4tAdKTmpCW5e504AV6rAsZ3aj1m+LxqpD22kAhpdOQjwXaMvdUmHkk
q+doP/SbG/b1d1kB3YdLxm/2qjbLRQSznmrsT+dHNzPYnQUClZqUETXYpfpZxnzYzet6gAgk7GOS
xmsXWtuEmAFsEqflXi+KFP3eHsuNwKPqeh5zq42NPm28ndbb/F6FPCzu1ah5DE3UYvfgyxTNGXCl
KHvvO4PwiuWtaDEC1PS30O+42lR+59ozk+1G0d5/qUQqvCz7fi2Xfvx4i24O+B0OHij/lL2VG7s6
XPbJyAZg70cDopf4i1uYs3d4K9IXm2P+uPKbbscMyulOjsSFc3vSeF7jddTLdcYMWFGJ5+a8BcP7
7Qbt+6ARWB4WLnNEvflUSd2EMz040rHzIlB6AhFQs+3xWojV7VF8KW4ORmL5QkbOQIX99p3+I3di
ATo3E5WJP5z+O2tkeJtwIVXPifVhdbkuvatci3RYiKhwgOD1MKw6dKk8qyY9UhR6Np+GMtkkcFTU
aNFBya/vampKk/Z/P5/4qZ+21x9Z5mgnNDHCcWRA8vH0GfakfsIpsxgHB/nbBWisJ5/qqEnJdjlY
7EQ7ef9zt/sHSwmrL5HMIgkS27t94SMPx8US4P/uyFmzpAxFe6gLN2BWkUAecJA7tk5Sb0gYBhrO
gs9vgevt3LgXEUvGEjw+Xzv4Q+hh863eb5rNptaNs+O24HBs5zqZG55GyeSrZAGUHjiATLlPsrjC
RJDQS/j5PJ8YGEr6qGFQKsE+60xnlHgJ3MPNHAoeUPmUSzs5yHSxeZZunikLOPaOipgC932re9vG
pWTTWYMZcyluntGfEsbG34nwHqfzP/oXDllntT8ukv5QdrUbqkdj/mZg3az4FjhEv52DkKRfoZjj
Qj9buHwptrnWFFDenutUpIv3SB9TDhCm8n3/3TBn7REQpbj9SOkKcVCF+zZlKbRNhZslHPGOYXpx
x1Juhvff6twmV4ZjMts0hNkP7x1BydFX6XQ6ZsNqjQ9Ew43apR1xjibM9qH9/Ckc+MJZ9s+bfGyi
bt6bRTxCe2wtOsa8F7ePC7uqjsaBsu45B8vWqrV8HUy9h7XWCzbawbU6FEiBBhlrhKSXqUGIZQOb
oidIMXFY76tUOgYzmcOXy/Aqlv3h7GE0voPgLSlPXAUVwdvCdF8ygKvt85jFoeX3J6olbn2Z4mz8
/MtF4ajgJTAxdTMrtCH1pacRktHaYH/yEM1jq+HMgD9wU/Ytn/1FIM90YxKTHp9mB6qBTLfmI8cs
Lewmvx1Awqc87eSlK32qprngTKenHPvmiJ5HalM2Dcf9yVB8IUQ5uhaG/iZyAR0Nhy5NX3W69EGa
RdQZZ8+S0674i5w43HKDiIX2LnWp8qx1/tInzIzj5Gryx7fOjRBo7kKcDYzSAwSleTUe5wRwKm9B
UzmMlSXCeg3+i+EhM4aV4IDSCFdSyrP/Mj06WgBC58htfwry6EvR7VR5HcLj8ePZODRtfQTWz+cg
oj9SEXhAK4fOFmg8Vhvb7907wJj+Fnsf4ZJv+muruMX8dm9QiAGbRkTkcCB2HuJgXKtY6gV1BOF7
fw7won4x35hK/8FJMn4srdRk2bsb+5sFKPf15XPP0k7MYBFpqgjtrcnR/uyGVbrN2AJQWBuBdIfw
0LylEPUAAIMNtCzmcFpWK7PdzPxDPl5xW+bneSodr4vrl27P3RHdo68lWXzG3k39oXEXkZT+iT4E
ZB5nvJYLUyhBmldCwKUzeF5IkziC1Zi6FzMT+55W4Ix871GtdAQpxDGewjhQyVDVm7Ctdj7MkzsA
F4izhjJWztyYLTwitCQqjErz7pL0zJ0MUs5yJOfWre7TBvM27rFYBfZcS9Rx9/JKp1MB9PlDOSiS
DbQ9FCFGtKHS6U6n30FlxCl4BrE63TUQUqdKC5JPMVkB7VqmEHS78EMfVUudCL+i9VtXEI3owU7n
Q0Eb8S4nklJqqwoJ+t378Km4IQsmEtv8Q7oN7Y8np2T9fcHb5Nse0oXgv1A3l2WnroxdfPIgkhQk
2TggcyAGicMuMU02XjA6IUR4XmHbUZvhmkoHxIv9QZakFPWzsyID/+ysknXw9AzhFM8jcoU4euu2
/DY5RXmnDhe8WvOr1XDPxYTFGpNg3TlpL6bkYTMWnRtuetofYHdunI7m0Kanc1+Op5rIIxsPMEh4
glFItUqgaHODRKml+N0NSIAu+VlnGksBDH/N9GM3a1KNXaHRfjzop7SxzuwXZ1Rj/57GOaKbCe/p
+JGCjtT7yFoD6bRLQ6g2vQBT5YuO1xt2v/mWuerqt+9vmAl6ocZYr5dWiMNVW8bkVb5Q0GK1x5Uq
42L2q7DPPQXWIrjH8svXZP96zHYle/1Yx14dohavlLlR2pOt1gWVTjKtpwrx9e1j9mGPlVGTZCvn
8vk+tFjDVUmBxk21+qbHxPeRIZIHRo3y1xnKq42fuNrVbSxfODpvgaDOWeGOeQJRFODxzFY6INkj
x5n6i8w7NnE1AZreU2KxsSLu8SvNIjLvdDzn0G8yAp3J8v3M9JdwYwuefB0hgw8cwL4Jsz81rhmY
/8CqPnYj8x6Ab23/Opo4icBmkdm+/9anph9vhbh1g2djjJCX/aZwUJrrI45/bZT7Vp5v3zHHUxGX
BIh2r1Nt12NmEMYfMTT11/sIQ8ObkU/zagayVjHrgSIk/brwc/sk1SPk4tSx+ZYX6o6VId/3STrr
kQlxz8A39TSI0AD2slBu+L5iafofvzaXUCwkbr0Og0js8dQ6U1xFVJ4bpneVZ/P8RP4u3uIzJ7IQ
b9mHNkalaxdasz9GKDK58f7fuYY5ERpKJb4c+tK1yAxTCK2aYOBslPq66xrblv8w17XqlSmiVP+r
A85PHBp9ECyNp9n1O3rl/i4h6VwdRS5oKwT5urgckO+nxhdI38UNOcYS2l/toMHyoVSPH7SFCpop
A89xOnePIELXf+dP4kcY4WFsy6B7TRmK5ACJUBBa/R2q+LnIuRzuS66Gg1UotpNPzQ8v99IFQAQn
fPbwjvqd3HuBcj9Th+jTiFKJeV4ce7iqTvSYLmwUdliZXotJTNFsD1BTuy3cvOCCd6IkjiMUHObe
CeKmnjm6U1HJDm1pZG4LdxCv0EB0yeGqfGmZfzcP28pwm88uGMozdEB/VXeSAdlZ3rqSsCQ9rgmq
2OeR/XldJ/dQxgKx/ML2v8ZbIsvh2Tu14ZU7j9561XgLThVbvhBjpGsp7zcIg/WYMhnaQw5xev9n
PiR/MPfuWax87Y8tNsvElDHnUHtbvBSbkFQiRbUyP+88dfwW50gpaq4tamnp6ffakD+Z3Tn1gnb9
7qPTNZ4vBQDVjC6FNRnb6qHL64JVPxbifan+KjVwoRXkN/eZe3MElbBD3tePI32KJ1+M1T8D/yk4
f+exJsUTGa/xTQJNjtmJ5KrMpVpgw78ahKzvvICmgiN3X0bH2JeG6lBiPntqQMnkNedbZWgwl9+n
lQqajmlxVgASr9xS8rJnquhbVaTgjMREkgt82yW4xtHRq8d+U39J4P5SD1utlstk2KWQS13Q9gbH
G183Ok+GYc1WgHSgbBkgDGx2dJ39qKrPjvKd1j8tJb2OC+p5d6WsnwUOnqv1NW4RVv8EFeYWDgQi
m+M10Ms+zN86fdLgYFBEG1KDIs5JZ0kThyGj7KjKwnPeCVhfulEX7fLWV8DX5X/VV492tzdrO2lw
U2jCaktx53WVfu5Af82unl3PwBFY2mvPbheSqywqG7bXdpNFvetj9MplBlSnTT2CJZea2zJOKu6z
49GdpMg+J9ViVr5GCztxlYVmWvZiX8gUN2D7m6+BTFBO4ApmClQ/uaPSiEoYtaaniJvBIP+tEW8I
D/iCuQwkvO0vJdI4uZFStZiUVorH3khF5OvMibfexGGLf9iZFRRcfl4SMfZPp8qY3ccNAqcjxUZ8
MBfuYOWuazrN6KaMUygaUGBCHIvw37M6Sf2wV9GLQrQgArj6iqEFD2ffuG1nrwzihfOeiEiYaDgd
JorzkxAYEY2w969imV31sk28DTXM2s/qqUXzV+FVFYzieoLKrNRuDFKX46EwYZuoF4A6pwolgDip
vXvKUcubExdtNqiB+LACyIaAlmXdU3JK2grD1O0eQOLEJXOHAtQUgjvkoHOxlfIH5vBKE1aeAZxM
esC9s4XM/A8NrBkW8ajnCtpWvzhUQ9wUPsHBULhLKSqdEanfyqOYneh2adwDUwDiNYeBtOCpJJpE
O1moNb6XBtfUyGfssptjfH4fSD2ZcnJ06B3IW2noJOVEdcloJ/BFIVbC/F4S9vdEBGd8pbP6dnth
7MXXBFTL988KBJWTpaPkKgc66SvXic71phsP3oVKWBLq7cyyLCBb3PNj/K/HKJrFywhc9mAyVUOc
mDYvZgf3y7V0agfR1A32/5Lz7CAR2n/OEcrBEUS9+TrUglgexyX4b3PQe/ZBq5zyPXtyI9lAP6RZ
xRksqEg1vnPY8ujV2iYSn4+v7yW/XiD/tfGFcf9N2V36IIMxOQUXmNbo7xZwSydXHpPMWv9Y+mMB
SeF4HKW4VU47nyqwD2baYfGYS3Ub4ZBGlp6TTDvNiZBCOHS39C5Hq54H2cAgs4Bx28FU1ErXLBl+
FZPzenO6Cs3m/4UxDht9YOfZsywV21SCNPL+Vpt/05zi3YHiHv1lHhKDXWuaPYFhDkIajIjAcFDa
p1RA4xLn/cIykqhug9yoqbJFp9+RynsKMzUICd7VGL/b+psUpjfKCrV3SCnBPBsX+TnVNC0TdZPc
y+G9SsLMfK58/s3PDtk+wShBZMurCXKLMpoQGZpRvqsMKKb4EwERgytRicS1ozCPjym5zNa8FSzI
Smq3u0UOz41V31pZHt9rpvjPkqqI7S0N5erczsxt46yYPfe3lFzZRI7TFVuR8zmFBAP7puW6OvWf
nZt/VWIXiD7Cwt95WSDLzfXT2A39ptxN7G4oEGey6tXVZ5nuBr9sTQgA6WsmEXDf0GJmhaOBeuIq
dNE03nCvlywelv4yJu4HHdSiQ4Mr1djfuZbfjcu6jyMBBg/Te0Ru8hHnUl/pHfmd+TCS58WkFhgO
Q/QtawTwMZznKzAMXI2wiJxduNJKXFvHBTgWNGZZUCvBYXZtFm1kuPEvzmCWcdE36KOdzqwJogPP
ynioyh8FI+C9K7Mwv7/lY49rx+T/bDemqngSqaFDJxoVmrgSc5cYEYuRVq4dsbBbzXr/LTgxg3iy
enE5Qh4Ldo23jBeOEh4oHQEhk8hHVO6+0mgMStsd1xwJw84NiInMQBFibHBWsDkNgU0ntZ40s1Ck
0MSjGj6Tiu805inlTrml82eK/1vMZ3h6qugAsPNZYnQdL0UfVYx85j0vb2kLZYUBzzDuz7S2wApZ
LCjnWXD0ppa8qNdfBLn6OEiZxxNKPlvehuL8jpkcoiNHJonaSFUdRwoCu8mXhl04tSBNjOkBx5pg
71ktOJ+SgqEDFgujmC2/NvIQcy9P6vpiMobu4sOgGDeaJPa4ymUo0Ww9UHyoXEKiERTf1yXzbeGG
CMCah5pYvzj1TH1BQr7Zvt6VJXvu08HXZrfdIFI4CY4DGkzA6ULxXVA4PL4i8NVHA1RDKvbtcZAm
mp5RveVxojP7dU7CF8QCCCPamKIroT2BkAdwqNO8dAHo/qaIzanN1L7/qKvbPjoalH+94KgOojAA
KMjT+2H3tqYUw9lZ35/d99zlJO1pURx5OBkWTSjGf+Cm6FCnOBG9+TovXqBz1Oe8p2aipJLe542b
nJI0FRhDzZK67Bg7uWiVCP+/xETHWHZ5oih6VkgXEo4N/puEqQ0m5si8vAAKNUcvlFeiNbbrW9bb
4soSEbWX7DuAjd5ju/5Bs/ACy2jZfSqLYahZl2iGtFBVkO7SIxT5Bglsj0Zu7XC6k9BPiz2HF5p1
Spx1AB3+b2rYJH/GQLEEe/O/TMGq06P9Xe2VnE/veCyTvLjpGodmx5ZLLxMRwmWCR0TeT/CdPPe1
9Qu+hH/SMuMSz7Qlri3I7wQYtgthGLQ2IsgSKnF3zApn/9cKLPRaD0wpuKgkLZ2ejNSHCloTMb9M
1UDu3oyt9uL6z3/JGVYuSYf+Le9hVO79oR1ICxaEq0GJYbw+TzC1IfdzUrck6fZzXFKw3FPnPseo
Eh8sfLfoKhNd7qWaOwx/cRAwOxYFiBRiDhMmyZSNItmTU9nceFq4o0qTD7kRgDhxniqrfFOO0+rg
EA99Kev6D9y0gLPPYyquU4vuFoUhGzuE4c3m9vcCSll2Ydak4uYmcff2X+CxT3hMIwNJ0qirD8bs
VfW7BH+zbasdvkrTDjthySqm4ZggOuRxxfGZExv2zJPCPecODGqUmkFOENHHD9uAKQsDJJ+m/K6u
SB8lWWabhgM06nse4i3RlHmpUs9vWJl9F+pDSscIMLJYh3jIjRf/blzmzmTz7GhW2leFHrycIoWV
eujBC+ofxdOAK6yxAgzGS6zJmPWY+8YpNAOL9/PLuTXlZT+nVVo23DPkEB0Vs4ed1NCv6NzlQEPS
7x4IToUAowVjQ5luOZzSnWeNKzJdZBo0YSe4vjZ1McY0lGLDQnlQgPq20nNSGSfkxw/0AXPjllU5
R++VL+8496E0vUzCC3tzZXFFmsteOSNPX2gKsrGA93sOWgOERYwYsMDnPf+oWmRl+VAMDJqz7Na6
JPYQdJ5v9URdtCfMqNLMUs5T7hQC3gfAGFqhPboNPZMkBG8yHyfkLpLVmPSX5M8vNTVTFV9y6KS1
F3YiABCBopLgagjkPXHJRimyyfx1EV7UdfyTJUbiGVYENLUmzmY6K00RYrYMGt+fSIh4LVY+fgt4
3WpUKxVbK88DkuHRiASFogbyKD69GRCXKv20Au/2FUjVQCFtJwRqkMJ02gyJ6YlHkFdYdaPBpE+A
XBblaF745sIAsJ/v44mkYc2ertSyc7KaDumS7GDgWoC4Dr3oXAWoEXZ777OwAyj4SOFRSWOPTwTB
PEfDjmt76y5yKNTOZ0n2uLJUuy4dUBpxTq2aMxAJ8PBjmD2OumweD+LdySWCXidm4Ppiz+7lX9sf
uZoCCB7SnSZWQHGOO3W05OqQBXx7aB44X0YEUIiVLqUP3TYAizkbE7TXh8oeCLjDySp8knBu2lnT
wXUe06DjbBaQhQy8rsm6eAdKj4tGPKXMe6BHpp3XZ3aFTK+Zg+fLCblIAY95bdl1tQek1cZTQ4hm
PPhtlferd0QRDmjNNu4Tuo1CrDex2RFykGDIR3kOzL4I6Cig1MhBn/VUoSBL8Q5gL4grwRaD7CkP
fzjsO3Il5TitbSS12NGz967YOMtA+ruZvo5FuYZ1LOdsCSOnRXFUFDrwC7IoU5A4STyo5KXfheVg
xvHSw8J/KNHM/jay29q4fDv3HHuSS/0InO6+Fz7cpb9MEADH+V1kabribPCdN0qlbGcWcHfJZt92
Lz1FELYMhtctKnvNRqfyp3B1KHc9oSygmXKMEehDCftAvIfbKGa+xqV1xtsPnrso/I2w3PxQhv14
bZaG62e+S4RuSD/uAbfPvq3HLzs94Dr7SCC70Y3Q40x8IKpzNmIVta1ZuW+gttIaSC68sr0JVcp2
9yX94dr9xB5Z2FmlRv67y9vPVDOJ72CfC5j4vR6BSFgUPjuw6mzqiF9lcDY7x33+MztcDDExFo0M
bTCupFyuuE4EvDoQmWiE+KRjptVa1TaL14+0SykHrYULWdJ6F8RUUsrjcZLcH5iFrMQBo92/PNhK
bZ0H/+AslsorptFeeb8y5WOsS9h3nxHyNdRuq8OdlssuG5cbOp7vWy9LdghyuDHMAOERYv7NXdW5
pyMsePAuKgmnt4Wsx2iIrlk5eQiKguoKhKDMP+kwbGg72AluXnEsQK3wzlDUny+LN08f1O5BP1I7
bqI8YPQLXm1M6qpBa3gKd5/jtWpKt4rcTE41bK+5NI9YEayX16yi3W8SJqYBHbtvSne1VMLYfNud
ZgCpcO94AnXbvN/YbCjhq0qjdx1yJoHtT2JRjI8EYLhSc3tvGQl7aeLlkGOwnGcRkBzco2UeXpaB
TbSSAyTx18kHzKvNZ3EcvnUtQHyhsEtg3EA2NctMfY+qLtr/SUTv00umVhT6YSRTUkRCdVcxSH68
pCTX77HzfY6KouceiIo6K5nmz9c2WBiBZzNkT++kFkH14iS4YtimuY7e2YSMaA/yG/GMgpQJ6wRy
MSb97UHRKLPmyOLFC5OTfk4wuE/Ls/6VnPTjFg8pDS897/3PZyzYvjFmGsQMCx0JFTtXqi8AmfhL
cgWp8K86xNctrU9/QeRe94zGRVH0vjAT3PEqYlJ8A32xfHqq7r0gmLqPScfku3U/QfJfuJaTIlip
CfuHQazv6eNO17A3ZdFYR7G4zNANDzKfeStEN6i1J5WYomykGZPOEPgPEsvex+6AoIdOyWYnnZpg
W3mZd1SkCeV9+soz4jue9gjXXPiESZcsj0N+g/4xC5idFSrrQh7vkmjddK5Kn9ZqAV0E2I6cjoD8
EDuDoEn96UOjy7+z4SMDTSlXbeOpNQVn5lo2R0Qj6SVnH2KX/PfyYreN1I2d8obAEvv+RnOCU9Cv
hijQXslEV1seSaJfHxun/TSe4iZwQSHsPLy5yXtMQ7V90pO/9zgLeh/pB3Ch63Syc9aGCR8AKa6G
xiOkdSR8plbvjn8TFGNnMbphibKnIEwbatrrIcYtKoWAyW80mGTLSYEh8jggjpec4qapQOiSGUAP
dEUdJHtKz+3Q7QXIKJgjuSuRhxVZxeClP/YU6t6uE2TeyqlHIsmyCXkEQW9VW/kiDSGwPQusuIxs
PkUJeHEw/17ECa0j6j32Kg3ZOFdgoAdIurpX4ZQLlJRKAw6bsr1RrYSzAcsAILck/9GFolGhQER6
eJAyWZgQ+BEKJIbqcbS93Pu7aElqBUvm2U+gw19O+M0BmKVY2nGLfOJcE0B6BeSepGZvAky21KRI
/6qxq+Nav9ugs+hwQJ915YY0FjX+vw3hBZzClQeb78Ayc7HsfMoxbvCqqRPJ/nyfdmMFEVWbJbMR
a2Yqw4qtqa4DkhMsOioMreLr1BBrYbfNDr9s6Qd+6xG1yjhHgiVsT3qeK20Lv+dRdSvBWqTTwHk0
WZ19n1zxSQXSslB0dbHB539UIV/t9NwaIyAGTXuZ7ncJKVG90ow7ucoWpDBxacnXmuIlfYaQwhTj
kyHz9zbAlAEbS0J6slu8B5xhblpN7Id6pt122w1nNV/zApelHsjEZcqZkac486u/l9lt9KvcqqVG
OZ1Yd1OQZaOXWk2H5I/g/pRTYcZSWgQLTGNhQUhgbsZdB12ZT0n3eQU47JTOTpenvJc4B6bufkTf
O/kpxESm1zXUIBCFnr91pp3l+6gASE3iVdyC9l6EfoERGAlTrgzMc5qGLyFeIoYBY97GGLsvdfOi
dMQiWcHKwhw5EmihYb9GEdU2PJlGJTbdBQVepvSx/m3yfWtONkG/enV3jCWg/XkAMI1gTr6LmX/3
fMhmP7x3TOk3v9evnPUx+gMVFcz4pFiqhVI44khJbYTXmekvDgpEH3p1CiDLF/DVuW10cRWVsurd
UYHfKoV0Qsq9GuSzxU1uD62poSFB2XgZAhVTG3S05vVUEH5UtzbNWAbxxtBQ29m0LWJwKbhSFMtG
Y3XPyrwH0foOtvYROdXDN5IICn1gr8WQlUdv9czj00UekeYktzDLqKYljo5224fyArr3M5iRG1g6
/XL3p0bRn80+0Er7VkvQhYvgBPOvCR58U0oREA1E87iQMaEG/7tiiZGV3wAqrzKw/a57UJ910LiA
budsz7RNmrzOzNygNDwvCF9evGC4/tzfgQLX/Z/CNfavJ9t39n7GnsNK+QYWXyTfYxkeTKKIlDUh
/0VhhbZn8lDpPhPqL3eHwPSa8SDLVlFFD3BPUPqH+5gzxUeHI0Zbl2iwwxPJ4tdJpT/wmE8TDc03
xPxZyGew9TK776o7Z2WXur0/Jua3nk8EpoGnouwTaW3Z+r31PUmx9IpcSM2ZWXfpCN0Kl3/O5zr5
dumWbkIhKmtskdV42uREy1uSBb2z7FsGcF96WRkadM2CzlwohTejWvoMeptoxV18++PBjAtiIJ5l
5YdQ6lMsqB89mMuGaOeivqTI7yt1rJcT0k19aIUGoQ4CfGyA1hD/oAR7UQqhau+1VKkHvt8jw62E
UhrnTLNYT/x5DvRM/MQGklIKL8Nwip+a5icVwXANoZLF+hRrjZnT5exfJJzyo7IoD6GQdqo6ZPDb
lTXYICrEaGVehMUsE6U40V5zHMApKbKT4XA+EDeX4YXQi0PXUwLVZLYHTc2Nd43Si/jZTmYez4M8
CJduJmqCD0s/SzoHt192Fv+Q3baseqE/omuUsgCTwbvcxJhsOQCASuKdBV1Nys9a9of6x9K2zTBI
8h50WfKn0tHRMK9PRqGCJPNpDXSRsccWrvjEKZMp0fzbwRDMA07I3JlvqjAeM2IWHPx7HdUsOO4g
c7vh7uvEy78ykjFnG/wX72q95XQDMSGYO1sAUJEC8i9d/8z/uGU0yeAnfSw4wK88BXT5nELTm1pw
VrAdM9BqkOL9gnpgtB0T38/koFKq3v6l/wvagnRsQHZnj0COAGXJ7tRAqsdC6ze/B5WrePbdodtS
zVQYiuxEXcRWEn+yAUQukSfjLJiOWj3XQ5KcbOlEXMnjwPgOTxHSaEn7tpUjK1TdIl+jBT8iEZoH
FZDgX8w2PgYgep1ijV0WgbOTxszrjgBMM9n/ObB4wLm/ttW+2CxqGQ4StIqOtARIY4bK46BS3KEb
0kPSNngYBtW0OhnZfeHGRF9es2g/AqZ2LIOiwjCJ3xhdrSURiawTRwcn7615hKmSOPXMlyFydrQi
BbvQ1508n0uF6H12jxhg7buIdnQYEHKW64M3plotPg9MNY7mQXKL9bRuMV3PrCYy7YC/tEYzG7Se
edzz8+C5psMvJOv1ZrubShV/PFECD6fmUfzvHmm+kXerYYHGJZhQ7aMhkxBQskuT92AR4gIMojP0
m6L3fQlB47plH6iI5unTj+Ae9A9PgqsHi0d66fdmUK9yXFG1wbKXg8I9v+U7esZDCHokejdHhO3R
ErAO3nHHdgeBan0WdWNH74rdncqfoYIsNkSXuyiyz6cNWLmDAFKAtp1DvOxDmIR6UC4aUl0SD19G
x7tbWyqhZEPS/K57wZJnGBxCc6n0EgKD68tOf9fY2GBB+UOB9h4KNfiOaTvhaeHsXq6Msr5LgXCz
uAi8yhNep3bBa5IceIJi5gZoc4kXMFOyyB5svZK11qVC/fZcg5Jhtx9eBuTW4oWlo4fYETOAN3RZ
ve6G7AVJ69XgvnTs5XYK9C0nnr7yYYUG1DEnwUI41PEw8Wh5bJutO8UfsNyBjn9fKRVXEloYkWAS
FR9zT/EpW3xEkOXUbqbB7cG2vT+9cAGex7i4UJat9S19lNWkSdsJQXojd+1oWYzhKv3wH5vbuvZU
4AnJT4Ki349QvuIvFkKi+elkC5AZClQ+E3ZUyxmJwo6Mz8PVXcpuy5VQVZt6dWHQKTf2W3u6qtuu
s9GlDIdPzPNB4dD6BNY4j1EJomGWdZcI++kYAqX9SM/aGSMM3ZlFwQH2GnpemdgHdrT2tlCPWMC4
YEvQC7EIEkRXcZeiKQaTyMTLOb17WD+PkiMO3llYgtB8bdE1PCvDjEDlsWWu94vpz7qZeume1AzI
+cdGjXWBQfPZpA9gFQDiNkm5rOx8NyyjDelAzzN3TFPk5lrAz6PwyCKl/dyVpDK0AIosqIM3/qTY
tDETq35YR5QqtaX2t52NBWHgKaz5b4lKyDewmXldtLy2YR9Uvxhjsm0Hxq3JRhvMcFq3QQsrL8sN
Hn6GW3s3lGcN4wqazfQ94vIUTuCSCg9P0Deaejgn6m71ASMF3WqUfpEy9atkPlNNtusNLTxOagei
ETHEzzwp3DBFdFVMjqDLRX6siTWgT+0UvJPHyWI1Oc8oe51xQ/+YDbzMASx443iBFqqXLr0rtNmY
Cq3kl8dksyooCr3hdFVP9nnOe5yM/sYugRrKMF1wDVk4hWJeNpxwFLX9isX3CW6YSwZ0ihbmTWtB
NuUwhRgf8J7IfMQ391ULsQLR2wnv0tN7E9UHGRP5YhsSkQQJtjsn9ZEVq9hBbIGPR0tOPZdVtGqY
MCNacXbO6D+TNZF9RBjZE4Sg4IYBlS5ZcqzXXkHa2NNjWmRyTfKgQeyJopHukCKjQn50cTFx3HzV
Fm+REWPCcuIcjAmrkDrGpeG6yLdClp2gT2QwlLan8d8bPM1lNz5gIYdPrAoZLwFLaoF8HCZVccry
jolraZq4HTYZoIKKK+abn3TajVNPv17ZjsMRGx4zJFnevwtJRYUesZ0D1Uu3p2QxYpvhX/m/6kTz
fg4PmZMwrIEsQznFLj3NJViNk/0PBk+OcwTHvdv6REpE4mrdpA4VXjpnHCkvVipgg433Ql/d54f8
yGf4ynllWnAPPvJtLoD0UDnJRCndHueiTmkfHlMltsf4fMgZAMy+jSYRA3yMr4RgFY5jFrFLOwqu
rkG3bf1QsFaQ5C/oM2yJbR+ey/C8IsxPcyxqLjlg6MDRgwglvQnsKSjBw3g8wCuKVWhpAfW5My4E
UJooc+Xo9/6/GhCxdKwzA6KH0iqAJleQ2mBWW4N2Uxmgi+7CAg2vFWSwl2iAZ7xkqUXjCjA1zPCJ
rQvjsLpvE36ibU/+l+sX8GpnG4oUa1PrvbIjMYc1weqWD5YMYXw5m4+0nEnZNb1t66RcZE+zSsec
ImvwpiK/0eZ5ksm5fHcx0Vu21BKTVAa6R3MUJtSFexoyBPtl/oLuRpGDVBSFp3DcWhqdTzO9e/y+
7OKOl6HGTShgx0nhX0hCWhBfFb0zepXhKcsg4ZFWnhfiUO1CdQvE3M5ClDisst2gbMZz9elVAoNH
FaVLy6Q4mtwUUKdP6XqUwh/e1RjfJ8DIggsKbaZRLiuThh/PJE0bKaw+f0ItwSswO64XcD+pu8yL
SNPDvOsVripkBefJnhFkWQBtcd5OHrQjKN8X+L7pnIoLDtZMa2jM+MMYuKGwcFpQKapoykI8agC1
usePJGrrfte30wJ5R7Z/JObxGoaelSfcCn0A25tgASTGIJXlyfq7LPFeYsf2b6QnD8Ija+BKedrG
mGHc147SagbWDJ1UXlgI1gEpQQmxt37WDB/i3Em0pGvRICfN/gJGo+cHOfbGaM6GhEqvvtLyMeSy
nAodokgvBw6RD/7AucVjps+nqw5rKQjUUVcjE0DnAGh2o4HdTjvyR6uR+EPxqImEpouROrMYw1Mq
fhZiM32scNkhovVRZYC8HvtYYMC/BQd60SciWh7KDKuCGUNnkz+QltI5a73T07iQgPMuZ3TCb4sw
d2AplwTl8JS88VvT+l+K85cVhbdCwznlaYU7nCT6+N26ngMe7K3obexlK6lxl6m1qZzRnHsBjWOH
O8k0cAAEbFTTOX3gRH65yKcRDsJose2RpXPfdHiU3OhZRLleIrMQsqrnRQPZEZc60FCPGaq0/QSn
Et7HGl+YSDXNRIcUzn8hLlq8VN3LM1uz+s2szkwD3/4oNyT56+i1RiQLHJ5Q00YCBLJcZC5uaNAP
C/5JpZ9KP3NZBLP38ye+Cp/hGRgjPWzQfsKc2rybs6yUH/uJlFTuHu5SJKFKX28ByxIifEYkBgVp
wUogDBduJocDI/Rs+/fE3LA5O8sTlCQKBKuSb9gAP8lEva0c0z0Ak8edDPc6YGrWCBme5NO9ydkk
4x1Z/IT4KlfFQocpwyIcNQ7eemzbtH5niSARP1Wpy4pgNrY2dA3jjpceKTMG1UJiTn3BwUEx0wp4
dZiTF4N4b0ZeDK5vHw2u4bDU8haNLex8nhkPWrhFveo6B8BmdQreiuYmn5bRvnHWlZB/1OFMMtYf
+w2U6oPCu+OWOkEfsAEaOtmZB6sH4De3xxT5cojjDTxg8SNQCfeUm1bXOpntgWONBSE2nS4eFS7n
8U+g2mSIx+3u9fJ9M1vjvCHYe5gIWdiE3okghx4OO9H8KJyJwC93VpMM9nV5Kz6GssTsYelHD19Q
r0ArnQvcztOAXFwOw/MEssoD38hpEPoq6dQhMz6KCc+3b6ZoiOrnQFGACHSi7tFvvIECfo2qqTCZ
ppDOdkTZc82lep4tQuL1XdFV0OPh4uVTb8qD/jT+GwwhFk5E4VdJyfezOGCDxy4WmnvAgUCIRNkV
FOxvcnc2MviUwpYp+nayX7O/34k/2J/d5j46XC/56TAXglRa4D4bh57/yAwQmvrATcXEaYptGp2S
aYer13FCASvXeA0VNQffVCOCvwwNKRd0UFbNb3eqidS3IWB6M0tl63ilB9n64ZaG+nYeE5FrP50G
BDvWRqv+nUtA3KYrl8r30adt+VEtQo+G84o9uJirAjrQKTOmbyqHZANIf3a7gfuZ6Rq8KgxCPnUO
BuvwrSaRgVgqyTJJe7CjKV9FH8s82zFlVuWRnxpWZcqZBH8z/ZgG02ZtkEAjuGH+BKI5bnd0SIMA
KSoIQhIastK1G7wEYeY+LUdhjinP51QAMNCDej/zW7dtm6kBglIeOlGN+5QCfHjOvkoDQ3iKSHkd
9g41SzkrGKpNQfv4cl+CGkRqSO9vgIFEEtoSPjWH+B0sOD5GiBmomFPLeGjl8nfBRYxH+iagjxtL
hx+xaenTovzVJOuXg8xiLpxS72oDFBgXUycSfYDTImy98tqpNskZwXJ++813O5WpmVJasVgVceM3
ZbyqAV+pBzqN1BlM/Umedj4+hI+woGt5Y36RAnxg943rcnAe8JfdEn+dd2J23HtynhkJd9iCNNX/
OitfDPLEVRIhaRd1l6KoycbWEjGBu9tYpf5iUzVkVDrL90kLSDGouDE3zhxwA1op1bKS6QTFJJ6S
KB0rr1aZlZU9Rbs6lkT2hkyvFn0RQV/XA38jzPW8B5l1ya+D9qDU71D/rcmZ+Io0Fgwzs1JJmvYv
oRzYrSTWD6ptS6MZLWqVq9C5lEOF8P1jsxUXkddQ9uAvh4ymJkD05eje23RFo8K8bRsj/D8HljAR
/1xI+VHdLh2VGxfDe49VRAZjn6QVl4U3bf20ZR9Jb7yoXyW85Gu+RtNsQupRVutBAI322E2tThS7
8yUxRMBCd0I+mdz7/Q8P5FC/mZtROSp9bpLqvHoRpzlKCaQAiTP/ieSy8u5o/q7JF8xgZYvrOY2V
SHzF6dx8+tpwkjaVqiqwdITgZfO7K0fotIouM0Tu1feHy1EcuBUF5Z8pFv+EMK+O8QDMcTuhUVS4
wJHFLT+tY8FzoUXj4dryHV2mV9YCmhlSbsSMSfXNqEw24O7OM6oJk22O9koBeMy/ry59GNgyMYCQ
16nHUxFosCbzzUP9Ifz0jywM1jaM3zYK/mFqqE/qvqzwnRn1ZcavpFofNzPfItJvah1pNBLdWHRp
oq9mq8j/zArayjTBIJAjjnLFSF+puOBGsobd0ezlJl1iqgyzzo2GFgghpjIzn8rF0uWLIjZwmFuC
qrcKgj/V4I9aotDEmGm9nsEMJcnvTbip+rOUPrVhkSl1CWc0MNaSiF3S7O6WsAZCg0ItFWyXj36L
All+JapEsyzZc9Govxq37z+/800QZUJEL4Qh/MQk+x5aLL0DwGh1jd9b9TqiZn/2bIVEQEOToS0V
gYMisMFUF+ZLmoxmJip7+OHx4CnuYlRlz18nUtWBxg+t8uyhivmr0vpjfemybW/vIWL0Ns6YtCYQ
s0ftgLBevukQ02+ABlTRpLhEKzuM4ZK/t0lsIpv2UTSSSWO+5xDxQtapg8PYJf+tVokiTfNZfB1C
xEFDQq1YGys9vCoFS1NoPdXBMuzI07cOKBQeG90/alqePQGocmHTYhk7nW7aIKvfaD7HVxVCCanZ
SnV8L1cMk/q/4jrXA7iPzQqVwYpaSnZF+j9o5G+y4nQwiMEJIxmItopyK869sODEdqwBkNPZZ4Rp
LcJwz7SDuwAuY0YY0M4ueSYQaCTwldlWz773XgfCOd/11swFhXdtdg2hWLDv9uDCz/UF3/6JC1at
IEpKYNVahB9j/xwEmCcoUupH8Ff1k7PC5vVVJLSsB6l9Hl0YKiT8iTCSVY+7AvuKWm8fU8ecf7Sb
BI6j6EEKvtQwfIuiY7S7cQ20N6KHGdKQ1Xss6r3KbJWWijQO2EJjON+L7eXL8bo9af84Z1Re04G6
8RPsx+Plx2lcFYqliNIMSX14yX8OUvXv68x/ZSqpAmNdOxL1Lqqm/0BMslSbZ8L+cx16EL7H0Udv
DUQRJSK3mEOm9q/TPsIMhT4gRhAuVIqpKQqOxidOdg7Bce/XvWhb1mEmrjFlLAzHalO9XMwS25zv
qLIZjqrpalNBTuSoEPe9fH67dbsA1y5HbQpyCymK1aU4yjm7pUv2jIhuRUC1KxSU+7cf9k33mNXt
OqzvkLa58h+TEBTwq4I5QqCUVg/+TgzixEX8lqWyCcHnWVREmP50GuwFcaEw0HkCW48QdZwtE84W
6Z+ph7VkhBiNuCkqO9a1XGCqe7mQte5rCbiTjPXxFAckz4WjM2ZxOw2U3EwJ1w6oQDme9Dawbr4n
7WwdN+ruQdIH0HENBcTYULCqANB0r5JUddQIMIYdBk2lOdJfwe+DbsL7o8yu5olIFcm5whti933I
++/SmIJAlCIUL2oijjjHI0sgggGn5qbl10HS4Z9JrUhhXQ5iAlHJ0MzwwuUzwJ65Wi060lU48Tdg
/jGP2IX+2tjzuvdUoK4JOSc4v2SCbpVRvZgEvYjNsVkWZFBUlnAF/rkKjcrlLLH7bzjNRal/vYgy
1T9D4q1CZUPaZFlKsJryD1JrYWPl/1YTer2V3nao6rKkelFO1l4VryNa/lBUGFp8KyFK5k6WuyxE
Debfdi3plxwI567gaSfmSyguBWSpdHQBI3ZmHJ1VYCBWgdfn+8Y78SEZmvT9eV7/9e0EM/5pjHbx
dtyteN5Pqqq5EuwlluwRCUADV0llvaDyXH5KOVE7cSEr++UuEvi1Q8TJw7s/9tcrpJTtXy9uL1eC
csQWvM4hBrSnBbPIPketx3WPdRICHJKBngOIVhk4thDMObbqAfAxeLzCXDirlQRgQmPtNB+wYAvI
H4izEw1L+LAqOK37e/Sr8IHYEUB4DvMHgog9UEJhJBfKzKlquOTHFXKZ9Ii4e2IrNLFcgr9uptz0
tHAx7KxFQlk3QsStagJjKc7Wm+KJo3cU4R/sVDVr1Y+gmiWTs7jcBQed8j2dT2aLC13crtdEbR/7
SgkoQlNSQnHCOefrsABRp6uVxaGZ+97hFGyLMU9WA20HGCUujn1L3MP1yvQVI8nG22KAm4fockrs
aD2Zc+AP2eOVVcK2a1A/hdY6hVbX2RxXoJ+5uzo2238TB4ctugf9kW3GD7IUbxQ3Cd7CHFaJ5fbs
jdckLv7SWVxmWcYN7YpKFTsg3mM6FV2o93urFP2OVpyfBWZX5C/aiVBC7ZofdWduo/fv++6Ob9A1
XNJ/xaUnzX/APEckOGlAV/fgBbRgUwS7TOGkKaww+NLj7zuctHDs6Tb9bvqhumhzSftTNvKUFB5R
VJDwG7afW6aYrHsxrsmfGSvdyZ40yyakwEvjDAH6Kkmkbv0WYk3jWZDJaz9AepamvzapneMa70hr
qe2DOwD8KTRoyayuktBPcYN/NWqf+9LNiX/wbEMPPDGamLJpI5Fpjw6SXI6v6t9n5cTeXPvMyput
b4gm+L+fOhzPXRNwbe/MGeMOlKuPhlIXPh3kC4cozITEs/WCRM+ciHuu+1vtMI0DDoOafzJKx+Ob
nOwbTBw8Q7diSgYuStP9BtSridKVlEOzGE+/7x7eX0GKX3w+Fy/bwcawBMo450ky+u/m3aJLpyhj
mnax/PgeflhSdghj9lohp8znoFG/rn5FYNiZsl862JRcDqwEXdygxhQJncP7/HZPAoADzQEPznb/
DGx23vO7sjmDWvnYtpEWVcQds2zxf6cvDRwRyZ90fnPgOK7PtVqsm2bMmdGqoTk2eW2/370/IWza
36aMa0Hh+wBqgEatt+aBBc1v0O1YVRvBDDXUdIvmgV4iOCjk5So2rgl0vRKC2bjCJe45hoDZCsJ1
w0QreDoc6bYB4w6iY7YfldiJHVpRVt0L0fJ6JHQJBsz8WMup3+I3ujgMRgqQvY4NWOTygmDaf+kz
Ryfk6QOlH3WzrvXCDy8BQDxaut91jI9lwhWiTlQbhddwcM3Zvx7xzZq++MJK+oY0yqt/MeUxbYVG
pfs4cSSycf2CGg11Gb2FEq21IqSmhEoBBN7ywO2NnmuHZcDp3SzBE+A2cxLQIfRlwuihLVBxh6PY
rixWd65yrlZe2wlCbUOSf+Zz3WMsa4660WJrzO7uqrhVtHG44Nnkvd14fxAQ3xNbDuzNOZs9uOOe
J3PAaMJw8dtV+30IqIHEPUP8+4a0xRr4ozVOrGW0icM+l52C3scKCMhtU67eE0V0gSCQWbDtv3Dx
cBYgQmF6O+pKq64fsNlAyu0I55kWw0yhsKe1m0c623W4W9KQ+WWAQcLvas587FGYGVsW/itf6Xgc
9dFx19mBcppjVSvgvDP1n4vGBh1wYBTo8xjmTvl40Wylo6pcGiI6YYgC+ADbhqJom91+BKl94+t5
+5AA3pt9OP7Z6pJ0/oDRCd33/ZJOQxxZtCV0Zl+yI7CcDvV11/lt4Rbt1zsMW4kkvS3RFYc3FYrF
yy0x7ewbVCNtmMFA5Zh4ulO602i21ntyzcfQ/aelmNc2F7Lfi9imDnxWiM/i18Un9yMUfC3L44eZ
DhuUzGYO9RFhUUH0SaK9OREFQsVlt8wfEep+B8Fzvci9UfOyriRQm7ZtigZ06AYnSf6ldW3wH+lI
Q3Z+ryPaldCbnfyeIX46UtriiPlGDwijsVv5mqsqA1MCuaq84xMHsCI5c/XW/TJa2XxPh9OO3/DY
0nurPycqrRAOMubFBsJ3N+7OOMbfXWDEq40zr5hRZuBxPi6R6/mU5kihdcsUJF+zmqZFsM6vnJPp
HgX6zDm8vWOxJ6G1qvPMNcpR/tJkmla/brEmMBA5390/wbpABFF3B4Cw6zGi4SLEczngwPSoQlB2
nve4Eux91XTJVJAWgp4sMOWAiUMwc7KsOu1dc6Ik9tm4NMfwEjO72klfmn4QtC9sQHMb9v012Mui
fIeK2gfBG+WnZ2FLtKvKArRTHksOy3iLGKoQ38FdFuRx63u+i63YjIzQDYvYIs+H68exX2LZxGZJ
jg/E4uSzXQr6NFpLIVmGlnsG6vtSA7lTHz17t5QqEI7aGUhLKsSzadhtrF1LNF4vQ795zCNfn/4U
3GSlo9gvCaOFhuTHh0AZM+i5tDalcYG9ZbC7N4slkY1U/CWnav6wJ4sHDctHS36vZEbEzbULlzJd
HJ4GU7yltRhHpXswBDARFVIQQ76j080iZ3iTnKZ+2YcFqswmPajbj0SYWrrvkgL3bclRPkS/ao6D
UuwIZ1y4RbnzHqhVVEskbe+8hCYgY2ERPniIcuXF17+nT1rNMJ6lB/ybznGIAUVQciAu/PU3RTfN
pI7X51i5OZlgrQsFWTcIh4lFqDpPmN0ezzmTJtTPAG9W2NPYuyjZDFxXigNYzzXFBlU+CBReZYqz
TsdT595vTjmKja/qN83IAzbhj1XQerK9ZYlPSWWjKpO7XRl/DkdpkjYB0mVNYsqONsHEJr3pqVOu
5R2dkYhxBx6L6RXr31caJJN0yHlPCL9Y0ryYV/mY8IF7m7vt5Izrqq24cYxzmNrDYwVPNpH7dXqf
j6fC3qsLr+HqZBwQygir7W5vxCoptCoGfQf9iIu2HnDyUbNj3kSD/YInN6lSiIJl+VZWQzJ9wBWD
BT+gPaDtRDdEsYsl6buG6/doSO+XdS0OJyEjvrxoh3dNA1swj8piK5A2Fg9kaQuPpgyD2UGW6Vk9
J262lV/CqDY6DbuM0e/qqBEINRSWAj8e6XmbUPYOhwaL/zN54iMX+3hX3mPRuPu9yUrzriTKSWkT
0Ixzqgs3kZeiLsNFf2KgO1PYYDKViFk5AQX/UOpWoABwcaUu9iK89MD7QDaX7JA3ehCjR7A4IM60
XA/o5+W8xt+NXMTeqmG+Vkla/E/M26qESJ0Adm0bLiBmKMNmOcad5LwAriYMJfBtIPSyQEeWrLwr
HzvYo8k0W1SM+0NLV1t9KmUOpezqBuOVVceiv9tzZpK1Ifh6VRv1ETKGYr2/5L5WbY/EUlgzrjyw
bBCmRfPhacTKKp/mH7mWxX6X1j0C0GPuj78GtTItOpo67Z0f+blnFv/CrxwCboUQPGHUA07dkqtB
3ToJW8AWpgIw7Bg4J83aiL5GB1PNjYBlInEp+VOoH4syAiRHTGhzR1YGStxSk2RFZbwtasccPbY6
C71B5h9DPW2msdXU1U1IBvJXS98iAzkDwlsrWCglAGv+9imU6hy5l7CENhB6yiE2+fIS4XQYK4KT
7SfHWdDiU8zafj5y66+GxJR53eZtjM9GJ9zeo1tbrGZfnlW0Ji/HgIK1M223B6uMNRVneBI7TLf6
zKnPxp/hmtrfvhOo8Hgc+MwZ6j0EdTCwbdZK8VvCKABlU8ghTEu0xmC1zZNOFWfmzWX2pUFDJ7gT
PWkd/h3ndrk8Qnf9p2hc8Hk6Yj4UFyzNIUB7ePQeCacJolZXxBIyG4f51nclJkXNXw+tvATINBFB
a+wDNOHwWSOikPK23mb195VyyMeByC0cjyg+huiDZK03RgVR/L6oVseybq+boHOz0ie6hn4sr/AK
2AoM1jQ1hY1BFqeXEU1fITJk+fAudugl9qVrFiVGZ/CYDkZcqb99nE8ZcM98dMoz7TQ63K1jfR48
opMdNrLaioFa9Gq+OQVqjFs50bxtNb6tszUwMKMT09M1wrRNe/6KucnqA9t7HLusqGwtpaFuF49q
Gi80Wtaz1afHCMSVYbSWTwfGnDjMju6pEUepiHDGA79QROjd5Ps5q+EmiA5a/YI9k4b+A8fVT0si
dcP1e5OIEQQXcYxYujvz2enYKhMf0NEuAziXwg7amtYkJL+XrFZMsh7Bxq7d/hkn8LSrYQNYUZnW
VEH478ob7zyssbV+Cxl1tAUyMJFFk0wWo911zu1yeTvp/fBxE7nmzIH5BLtqZA2k12ClJ6HmgPcs
nFzkoy3Cy3GotnQpBE45OASK8XcYtrU6V/TpSAHF2EIPEhzGUlN+RFk3KkNC1FldCGF/OSqJhDPP
Q7O/yyVoiKW04vu8m0izjM8XOrDtakE/3yOhe9UEBh0ow4CwoIBjoWchC8hOKVzUL5jiM0nTYfmP
CTylhdOvIAO4yEtZ1yymemR7320+v3E+0ZfhkxRtvexK0O9kBsD0E0Xlz7S0TkA8S33rq9G4dVpC
hqCaf5qV2BYpODrng4R+NC9YX+J6rm/STKQRj1PXwXKQdmUKnNn4OSCwgqgVGu1gVBWbKKbP29fU
KJbBy001s9Uj2PC/2x1yLa1Uod/piDFYjT3fI5IoLF/UDGSBKiGgy5Q0B+L1l0RhHJXjeF7VVYhs
MG1Y4OWkD2Oxt58SAY3G0JIX5pfh02oyLzYB7d1v6a/tMQJvCqMGbEecKZbEhVWimfv3zm+y7rPw
EQCZMCb1LvzXcmJr0AFjo8tCSFG9Pcepj7052qk6yO3UpmW8ERBomElAvHtQahzMgTmBD+pjL5qD
7Ahxn0lbwyaHxjpb4WpQK+mo1LMnp+S4yjFZohW/Fiv3MYMSXvTiAdQNrcsKADEhEfKXRSk0RTSY
QrofzjfDPb6JpDX/X0hkwGvvyHnXB8C5FdbF3sw4PghY1MLyBQnlSJzftyi8ZuY/GgSAidLcY/Ql
mmRPOi9Hc6eIXt6sUs+l8oQvf+r1LVCPyw5o/yfX0PSTCrdWfAVY2ZhKbMoUeFwJKd2KxAjpUlDy
a3AjIhDY1oR6otYcXAbYzeZJ3+x3UQNqAUmpueUm41F3xgWYsTkRPmHMiiXHAoQuSYWwNFzOEod5
GdwMEGNs5jjiISL/DtUo1ilyq/kAQJqvAmuERb8mUqhU9L6fY2CaZprFmlnEnSTHowO7qpNBWRHT
gyV6hopY5EQPrRR5OZ4+1BOgSlJf+9SSfbxwm8LiLMA6IjXb+6J2QeJFmU/61eHu7alWIoGNjer3
Le4DtrK42eQwUgXMVFvNhmZhZqDTCKblw6pWTjX/NR1ezt+p5N/yyogbFyfnSk0M28OmXsfBabPN
Kco+61Z949z/VIgmbDAuw3dzBKhaT0Dj5ZMZ2aDAHFLPDOHmKJScLxaucjJo/E/kV/2+gWrq5vxT
1glSffvTxkrmyfFhv3p7y8jKa6bFoTZPVT5MGowDio/kF04joOdoPSgvZ841ick58uQ50Spaq0LB
27RRmAjnPwgJoZDGm+vmbiXAA068w4Mc+WnFXrYIi1QEW+wiLBLxtBdlEnugKZofFOyoIUaCVkGM
RN0dn+ZXxg/fiV8oLkNVmF2QTZJewZpoD+cep0Thxw4g+f8vI7HDv4a5JQJHinQ/FkxM7zON5V71
uWRX8sw8lpEGULH0j+EiIyvTLZ9V2yfMKydolixLQu0kbaPB+3z/khexf0ZVt7MXK70jz1VXrPtu
+BJink9dSjQr53OwYjslNvCANsNoWflXK0ej+i1IVeXA3MmgEEgzt67OWkZxPQM1kdZyHRmVakVl
z+WeflLIOZ//WYn446USZx9scg0KUcYy8aHFPh9Ih39hH5iYVgAJgjkBmgAaO+7nUMIrCSQimzkm
rNe4t+pj8ENB5y/FtfITwEUVjd4GKHPt0hAykIxFxoPIywcMC1UsztuRH3mxEW2MYAMHOvbC6bXS
oO32SuR3uAFuP21KF0vcJKXm9xioDs8a1C5V29DV9qlNmBC87GjUewj9YO357huXZ4VRfE8CMH/r
q3PuJfEjeb1f9YG4f8CYkX02ti0dY34OP0h2UklihONJB9bsD8Azo4YA/pBkRzBqT+C4QPlgGW+o
XsUEp4nknp8Tg5X3c0FyncGaPaoq3WXMy5M7z70IECTJKKnMx3EnFJTLXRh4rCmXlI+QCZ+PfSR/
iXwijQwg5q263RwVpbaQc64TZnquQn4C814P5K1JcfWNRxLDRBnahYaKef2YeteBpDgbc0d7tXLX
O3lRLtdo+DkQ7912wpzowjNqbzB8vWEnZ/HiWpTxZHBy5q1qUjv9L/nw9Wilo8WUX2XBJ7BDO1J9
rCzME+8bg1LFwFyWSH/AullkHxtA9HSVI42Fe3m/KM5pnMN5dfL75YATcon4U1KvgOQAroc6PZRm
U+Ozz/oQ5qu9ZTqzL6ei+KghCQohk+WVoh6xR9zWlrZzfGnxLrKFdx0kF9M/7ZKLNLUDoSMCDcRX
q/O3kXwHWIlgAheI/em1rFHtcB0Gt2uhehkf3moAiVcUztUnbbtCPgMlTPUdnvIDCb4ErtcuKm0Y
pQc8BoehQreC5Go0qGni01KJYf9fbDZU8sYQomWeSR0NYnjfOYrZ26kEMIwxgWrNU1jCy2CUz+bi
mUing7tbRXD8LzXou9pyuW7QzPY/qPN0OxmPlYDb33IoHWjOYSnlRRb/Mj+RwXa5gcw6VLo0cHCx
WhXT03mIKAqDUezgPTw6eMW+V9k+lKCKNyaER4t0/JvCyXqKL0C0zRmzJiJOrA/m0D9pS4c66SNi
dxJdrQKctrSH1I1C2crOyiEjXgoYN+11S34WUp0REgXRuJFYcTCk+QgydynYEY8JqpymDjLTLa4D
3fSLJcMSFQlS6XuCUWpACMbjahOXqIFOXCowyOcEpdftZ/T020UXcJGdbKZ87IZw6DlzZYhd4WLE
DVPzRrD7jaFsIH3fpA8TWMj9EQzsqhRTgX8Ts0mfmn23VUcvqaVsPZwjUTmHRUGJMindKQ44HUrv
ypkuW8d8XkhRkrU96CEkueuK0g7dWqaQ/dr5IL3xfZ2wVXNTTvzVPXclg6lGu7ra4XM0j9PuXELq
UIPr71M3v7ew6mUlmDZnRu5XSg6qOtuhX3zv1yHnSfNs3Nf09r1LGkcyrVWIEAcazV82ByESx+D9
Fwgyvl0sdHUwLmIhKvQ2HSwGNcTudBtzHfp6iW/8kC4O5lNa7+VvrYfssBx59YT8eo0Pg2FfrW6E
AyJs7ajj+JqYYV1sWtgPcsUhMHGU0nYbQ6izm2/3pmvuKNHzbWkoknrjdHRm+oYSksMngXiALuRw
wX9MXZcoxx7PuAErbYCj6hVYH2aJRaWfdG8WX10We1jhFV8snMTFWU7XQoX6kqcfAOVzeR2D17pE
bMpXwlpDD/EBQ9/nwSGbQF0NeMiG5SEiBtXk5WuO+ZdMd/f4qf1A8hNVv8VmJDfoPsjxA/mhBjrF
mHiZeaN+0DHq0s+7inCv2qe8VRxNr5uUVZxcx+cNfzDWzlHjIAQnEEJX4FxPDUfeRH59ASS4WfM2
BcSfxG5Ol7zg9lfww+1F9CJP8PUB7Fx+AKmNocmk48HBh/kFrHvv85Bj4V6SeYK5phFMfF9k6QDT
sX5rmNEj2s3jzHg+yKWhPIKbRiXIDiK1TZBQDdL4yGuXNCytXmMrF3588sgOv4RpZYqUr8etLDdS
TGnwJDYz282Qoeqr5QhiBZOIm3WkAHUydGtNlyF6AALdpfLn5id/wJNLPCfGrSd7gu2/nODYlraQ
jdMynA2SvU8VuwjdRioiwMuVS/KkoIVvezQH+lTxk3lTWyTGqxQwsLUFjSZOde+v+ASX4hXfmiry
zlCONaNvWJhdUwUh3/Qz4Cd2H49bbRUelhZmzSHHUg4WR+ULRfu1dpZrqV9VGV66oRgFAdey9BVI
rj7gtpJ4ypWR8bfCQ69gpPakxtRUxkwntu1czNr9jcYH5OIpo9E30TPCyXVrpS1CyminUj+rk7tN
wyv3Qt0ClH4CIe5j9gh7kPYkTGtdaxT5z49CpsFMFo9q16egqmjT3LnopikQBnWEcRwNfQbz2BpT
U8ExpWUpz+jlZ8YABrTEGDQzYv/Yb4UMBTu+5DAQfTbd/dWP4m2/RZ3a6KSQsm6DaCRY0PZSIq7U
cjxONqeIaH+OqgOPvarnBFFJ3R8iGVT69HfvgHvlDaZKn6UN0WSOkxPx3tVppueshzqVoaAsUrEl
9GtytjAK3By30XQm5as5LCqi0LH4LZYnQP1gQ6sEijYSepeEjlP+SyeZIbSihbG5YiW18HlOdtM2
aCYGE7khXCsmf4/9leRIaQDayD0PwkMfW2pb1YnuNaTRKCic04t+9OPmflTAOi9IcqGP6LAkct9I
0gt94C4LCJ3KSgnAY6BfxbPyA6c8VoXo6EKolU7p67vquJlZUHcNqmo1/MsxR2MV1ZMsg9fzKLJS
dhcGVyYMzGs3NwLoEZnKuR7KB8iE9bXVCTIHsd2K//U1OU33OHKzaA1jEq4p/acpNZKLKHZ5OHXS
FkOTISvoo+QG35MnmtYJWbPDGS0IK8TnU92YxznsvmzyjD+0wSwdUlc9ir7UJwGCp4bFk1AbvpfF
rCALsM6vfWTqOFJFJL7MgFtupaQzIyfZzjJuCs/LSuiC/04MeBlvtuhgmFtqCGfG6WyB28fe+HI3
uWRDT7kdPYqhVFuO3YX71l6C0yP0Lm8wvpoXAT9Az5TygrEYk1BY1NbfX9t4v92j3DkrOdNzDx/L
rcIn7jw/4lsRWLXMEzoqlfj8wff7XGlfk3QFjh7t4ouO5X9IuoDH6XDa85zOb/phdYu8FEQnYUb5
bFgsx4YUnPlKOt/jNuYe9BJ30RwWfUDJVgZ24LY0br0i024cxNt6WV3zNyheCQdSOKExGbfNjiWx
cg/1ha3XkXvWxh4EmpEtVaLhWquv78wAm6b4eHPO8MCuBgv7THUlTGftZkLtyvTkIjOHg4aIfzQj
jljgWPiY1THCqeH7exHBAg36nYvq7BAGpuC+N7bwdZZ0JM6e3UHsgcF4FPIqkRQslLFJqFl7CPbo
yQxtNOq3S6VLT6SF2JJR5+jelMMw5d+P0G1VP9LOrDZ3ERhLuTNIW+/iCcxgjHAGlIx9CTLp/Hlz
c1v3wmRIc3xfGMzbk/ARBKwlBNmH65j8wSVvEpIuq1mASpdDxXaWkoCCBtyWIajK6U/3IlhBF4Q3
rvTpOoKIplc7rLJ237xuYqVXi7L2OgsBNDjficD+CA6lA85u5KBPdV0sKHX+Rca9CT3VWdqHaQ+t
Mhn2HEJtv6aVg9w+Bx3kpRwcs7V+1GoZw5HVDgmuBmwfaJqP5xtXtOsAvlq/AFh9/KZ2uVhHWyjG
+jxewEQoz4IGeKWsC2isalYy3dG/FP09+1jYXhUOERu/iI4xLi0IhGLN188F6JrmYyH/dmUZnYVd
VJMp0FfzCHETZqrRUp+ZXKrhjb9cQeTnZ82za+GfQqfnfBbbtWpUHimEGx7aW/ytPEuVeSA6WPyM
xW4A6WIaieDJFtkwvSmkjhfiHZjGiqwFPIQ/8wHpUBiWlC2o7a5m/Xy0lUbmLoZVkGjT2sbnJ7fF
nwv/i1T+jTQYo9Ge1ZENS6/4JlonpbsYMREXPbOdBkSoMmMGPq1LyU89Q0MqEhz4Y63NAUX20+zZ
Gncz8KCMTzKSEOTZounn/LestBGhm7EiD47dbALKfjaGwh3kRoSg0T2zwBNepC9OLR4psg0LQ7BX
oFmgf9xNRVyzvqLd3QZbHjEb4DLQGDYbXioLzpPJ9fbuX6rp63YREZfcWPqk1DxMbDdBfb9C68iK
anJOLHQreW64azcdsERIvWFdllboAfJCb0MV5s2gIkA9i3VsLZHlv8/Fo/gaQv+SRGvp/nAnuouo
1ui66bB2zhSB4hLYVb8vE62ccRX/612UHgYj61hBQg7rJq7eFaCiMJrayaIE7rxpECx2j1MKMgjT
08y5+pkfYDoV37Muhdr+1bfQjuRCxhpclocOdQULDiKy8duhokRuY6NGCJzLGrcD4bRsllcO7jdv
ie1U7hLoq5EzEqBzbmun1h2m3pL4e3iD9SDg1zzHrmsF04T10ffe1F6TVehwebMBnriVgMWYGMMW
WVpILIPVdJr4t+Dvezsew3jG3fhak/4xnnUfXVaYrXezm1xzOdygUSVsmUtnoPp2q1fWh+74VMST
JIzi7WqJ0jmY6gzivDVvKHIfKuOCWkuJTTb7s3zmbcEOjuSyMpb68ra72i9iBdposwsLo4t8l0fY
5f4SIjzUDluTHYxbGruOxCo9yFjRLEmuhggC1YN43xS5q2u/T79k+NYw093r/cZtpTl8JiBW6AZW
y8R2bcOz/qNjVKm/y8Xdvtt/0aJBCNJuslrNybK/fAepzjyNbMGWoRJNb45mkO+ZhlrJaS/h1VII
JNgOKcRPH7tP+4g3p0nbnjlCk4aSnGuHUvy/KRq0AjTTJvlj/X6+N9iT3q74n9kBwX/Lzt7evner
pXqG1tUBnHGKQxQhI2bQx+jAdyT6H1hFaCwhgn0zSSHgTJr9/nTN+wduqP7/x4iNUCtt5EM1szUo
ML+xtGhQSX06Yt+TYkuTGRKo52LSi2EgR7IJ4SyeJCYc7fC8h6jgFck66KS7cTCsyueXHy+rv4ry
HGPGFXgXA94WRhGgx3zj9mbI6YY2rIoQF03Kj/dmXsi+w7OxSvWbhS0JCi5gUB5sXc7GtE0FAQpD
EPD5GdD3LWUZ4+D8+Qx/KBTUBv/O6wy9nRrXY6jyQ6dMmLNpaEZmrYU2AE1rvwBXmzJjpKjrr3Ys
Eiahy8M/gFPm/b9NA0TEw8hyHNMVNwYbG8q06Vum4pcXWcMlEDQ5rbil3q3hgnuIhARsX8f2wWGH
6F8EkMZJYYucybbvOEfoCKb0dwmRM2fpP7SVQOtSY7AatmlqkTSYCKT+MGHoHkVkG2nlsqKiBGIu
6eeAfavfdt6GmI1YuRrcL43qDvb3XRaD2wfSTewNKm8IdSCdfGuwQIWtUPoCV06XULwD1pj7e7f+
eB8n1nVIoaWK6TCcBa72H3Pz+gbL0BKl7FiMUJLx/fFZf7ihTeHPLOlt0FCFsXbpD3NtRfXk+R1v
u3/1eJN7BWkxLFkZQw8F2l4ZloWyDHWmudx0slorpuqRUew05AmDKY3xTfwy3Bxb3G49B4RhIbfe
M+ukO3vF8+uLC73yIQhm2KowLwNp8p091Ag9UCQkWkEh+Tx63+JvCSVFo+Xyw7vqG+vlhcMmhx75
CncdJC6I6172R0OMmxrqpN3ohH+jRaYs/asdEYSUipLloQxyuxXITebasF1r69YmisAjtT9uU2my
ficEz/afuBJTU6uB3H+uyzrmyRFeyPvsLxJVjx4R6T0IJBqivFJS0Y8bGybRIpGdUqoTlJitn/PG
niWoxg1uJT+E1FrVe9S5eysac7442sqxi8LW2r9vBmeQ1JlcxsXao6ERqsI1i734eQLOjkMCQNmP
XTHZbnOUnDZDx9gQuEeyJ6ljUMCPubMDgRYKNy7PZ+DLh+l/hndWr+BT5qRoJKZOGyDjqXujQfUk
s6c54fPsD+5/IDKtL9aGhecZT5PIYwBDJc3nkguRNVyx1KkXohB4P6idqCVvsn7uOMl9ysYF2mZ7
GwYbvBZumlCebS6nJAb5Q8dXr5JHDtGVuZfzTSFL7SROz+HqZ7TrbHWHsAIkrijWAwvwrbRUJgJJ
RqfArU7gdEQw7rDpswddefx/e/4oNJ+OK4k/ymFJxKylPd3z1BvqiNOAYXSratKxi/+wQanuqpD2
WEbsZn8cqBHz30T5cgJuKI+zKKaUxpfOf7fkv4rAOZmqac5AD5LpMDsLxnwFdVnO+OXdPD6uHI+2
h68sj4GCMSvyzw4GTFku6KdjxaerJs+xnDSKJkUAju/6c6/W5GC+/9SogsP0+BSkV5FC/nCR4FSE
tACzgi7hdf+9GelY1NLxQmXzec/txeDgADilnqA4rB64qCsPyTtQvqNhQluXZH5lh/rpqUM9wDNR
GoJU8OMud497NV4hQ5hHhyn5n1JcDtxDsPULHpMV3wh9iwiR7knkJoQEa9QWMONovFoPwnCLHbPO
nIISL0pwYgT5VW1+bP1MMByZelTjMwWN5wP4mCgDNGYQkjdWWW9PyeVh8Ep1aHzAVDvn1wFJobH2
SvmV2MHVPQE6UOP7EDPnL+1fV5GpeyEWfddh85AlxfJkriYhEA5mRMjkpuiQOZIe2hqEjlVj4Vor
uRI00Lt0q2pHGErhefvz6VwSDSpUcawIl9dD1U510Nj6V2w9amoT6vWPLgy9cuntgDJt15T93kmO
zfZJIFsE0h87wDiO/0aZ5GvVIPU9Qdwc6VO8DxkoTdQiALH/gInPyaQqiVSPP2FPfaHf9n1AzXVK
/OXdsjrRcFe3OYw54a+CwuSWfsawSxcTLJVfYORkDOVABazRydiv65T3si1D+f1hxewOTbE/vMZi
QjTxA/sog9TZ25am17tw2nfwCPHG3rDzSpySL+zr/dleOG0o7f5t+EGDwXye5leJaKG8qPua3Jp0
lhyy3oauI6r3rtq2bwQjrBamNTnqdjpqpLQTCdh5xWVIgD+gsmnH30mZNeaIleSKtvBpIt/ml/32
JsYfI6BtNLWv/7x/YKmV4uf64jiXA/01KzrKsLoHmmplqzY3LJADePs9VmiBwFMFtQCTIwRwKDwq
+znIyjK5Mv57kcQuL5DZd2/EVcjPWVJU4Sq2hD//Ap5xmvREK93KwreWNV4ePiIBHnqkDbO37B9N
hfYhJoLwvH5IKg0B2Xj4JBfxbOtFIb2GZNOYoJwTU3WTWe+W3lG6mHaTZAfGSES+IMnzyfuYheK4
knjQD6mJKuda462wInwOeviwLu2CYKxasx/nKvzLyLM4wBDkFo31ECHM7ULlH+EEnnPvyDT3u56j
/sgSLEz2e00ktLUJ+T3njm2o53osgaAqAp/DwWGQZXrgkgcFJ1b6nydp6FLC2BbTBi4Ohmvr5SLr
HNi8CB3AyIryClY4vh0M2uSgsnXuTAW90zNx9u656hrZ3XGa49UBstIcOLia1rq0nqjvNWUt0YfI
YCrfrWc5VNSkXW8rBI3S2dTpbok79QxFMiV2Bn6lnWDruYaewdf7sJRvtgCJG5yAIn0zoXjPcfB+
0r87gzpcLeTt6l8a8eQ33HixgGD9Yw9t8WxfNbljyOwTGK0NXzAmDsoVy6yCMBH2536FR42XWvLq
1qoyyuWZ7ByGpYL/r6/FyeQ+1B2j3qTGB+I3ZZoNruorQi7ih4cDz5z8cdZ40JM3NAcfc31wXuqV
0UrF8XBlvui7zXWxhlvqsvCFrYIiBqW+ZRQU6KFStGsa2QyYNeHy0QjJ5HXte1MmpLUr+f+UUlQu
gdLYCCwEU4RcAmxAk1Vr06NcZyb8ibR6QNyF4yOVUiKduc76tNRUQpSYsw0VzYL7+sMUE/fN4sm+
rkGI4DqDnzYn8NdYB/G5HZDHKcIXqjmYgdcIr9nbvh13YltFl3UY0V+B3rPAeFzQd1iuKO0pp2/e
e61Uk/PC3TcsY1iq8xoGDAaH8QqaBuclkqQO5Ybadewy6l+Z1oTjSw0iqmGCWwb8VwQvvcwmbWgF
MpSU6i2Ty/eqZ5V7vgjY0IqI4pMaVb1un2VFPNxxuyhs1oZJfM+cP8J44hsbaqZhtItRKEpDu0ZV
+aBjVimyt9vNeBpOI+DhswJJVejMhkvicY4bp4pnUWiZ6Uusi/CMTb7tNdLe7RsGpxZkg8bCTLFw
6Nc1STz4vjIbEci874OON8MckRD9IKeVd12JL7sb4/CqI39PeHZLUy4+97VHtC930N14x5aYDu2/
ANRFyEDRFHcqa70UKQ1QgMLF2Fj+NxyxFhHHnhgogX27kyiHatSMPiiLRZNygTu1UjZMiRIAU/T0
lhsXzAIIrHqlImOIuyIArUMePCQnW/uZ5108qDWvaksbcE3TQrdx2Fvve6Eg4b8SIKV2TO4tDFSI
kqPR16VDFfVlBm6DXu6Tr3zu9GNvDWAGyI1z9niJBqwnvJPIzHQFWswfXFbNHDFcsaqqNnphcZOw
v7Ae7ltUXpTmHSe4o+g+iXFpnoGIPqAZoUO2Q+zaWswU26QZbZzqzcrJ6KOMqQoDnmxXfL7AwkzN
STjgmFvCPj3lIB+91qlaWC7qwBe4No2mHDPGPnLm3gqsSn5s/QWx7xdW/BGYIRtcLXvsnxhjg3vc
QTr/Xx3AHXWhT+EP5JFIDzGCzvExMfiAE2vSNkmh3zI7y73fR6LYh4y3LfbHGjELS00mrSjVlN1o
ft76Jo/5d2LS/fi9mvAMznmTDd2JkfPRZhS/YgigW5INFpjFKWmTBYNXaqm6Y2fRwWMSPESJ7AUH
tEZNDaRL6C2MycSKodo63GvrdoEK2D1c7SVodrAE/rrnjY9CwhiPTiA33Ylj2mPjq22UppFwssQi
T2Eu3923CMUfPxbw9sd4BthAYO0DeYTFL9dntJEbnbsrBLz+zDkYFsaAzsVJKc0kMLRCwTKiIySh
Tc+XVmvIohlXV/S53QXaS1abWFwB7ReCoPSgfDJjDUtY5P7p72WH32KYGQ7OVFJ3HD8zqsiLrlq1
bCEG2G9TUx/XnrHogbqaGmAsMfBPtQbNRa2dOaS3069i4MmZAYUzt/CdDTNJNqVXKTXzYhheXhsc
aNR8G3eDy3MN9Yrw+nHZfNJTgVWTdyGvdOFp+3oWW1O8mGUN1Jh+2nQ8lCJrxyYPIcHlBB2YioyP
xQfBljuKt7nT4mUc8MHBDXlJZmvP3qFyFMNyYi/aTHePFZ61uUxejh9Kn2/Zo29SsFlZCZt1RZHL
pDvMQ6beyDq+Al85aSnYp00Dza65mNtH+XgdqfG5/Wu0hYiwwNluXpLqyWOQtzBDRelL1NqeRP+H
VCJIEDNjx86zN2O4HYNo6BnSpmHWM4ppFoiSYzvjEhQK1KUihnGsPTybMOXGzfsOsD97UUyWC7YG
VLcgnepUt/dRhEe16kXwGocAIoMdfoVBSdTG2BhqwxSIKw2+xRreVcd1YrWaX71FwvkwREgKbAj1
XI00fxwWf7cIMs0tWWxDeLdtC7bxESDfBhK7SYo4mKxzOmN9ksO2Psi7cnqQ4E/Dd+CK84Mw36lC
i6V+CwkXHn2+OmWgp4Lhu+faNHiLTH2QFMtRtFpYpl3pl3NJpE1gOvqhiUFEw4N5cuzyGjsGA8bh
comu3t1q2uwRKoZVARz9Zx+fsQIz+NhgTGQlG2jIbKlQIoVqf4HbJ/zgi9bBNH4jieMHhDScENeH
+WtcWeb8hjZefCEw7OpNMHITMea3XWfiJcHFmJOJQ2sdyqZjfuaVzafIkTYILppy9cpdzACqtzCL
CDwhf/Jx7OeQfg1991g90gosZM9pize8VI+a8BQxJxrcMI9Suna7wx7UGbYVMoMa0OW3sTiBCccc
ccIyHO+eCNE2ug2ClkgIUlTb25sW+sombapALDv+BSuyCpecACDB5KGyDV+ZklS17GOiApWa1a+T
OW448kP3dadF+RtTimO+Ye8UVQKQcYbojWFglOoyEeDkvJbhA3TMqZpCv8gx1Z+g1i9a2JtfjvS7
sHjd+4ooKTe/8VgG5xAFhP634tCgwc2uJT/GyPM0f5u3fKf4Ur99DX8ZyBMlrMo1lPmjqjoEcln5
L8FwYLDmoq97V73eH2jF/+wJMsGE/WhQAz0hen2GS07NzDzBi302ebErLgccJcyeHK/ivZ12Ugcd
THdAyZBElA0eFKzhhGi1FFE/AwrHdZAlWXao2zKl42usccb+O/JdGrv2AUORn006vcvnkdpj57IT
VpdYwU4KYcif3dveFbi9+0OTnXYTY+Wa04JwGS6BOnpT1s541HrhFehC43rjznUblkR3PufNu+Wg
LDXHsX5dP/xOoHK9N7snMjjQ5PsybAHH51UHmwxRRx+PhzzkZ5Ps12zyorFBTxg7v2tLAy/u97eD
lKDiZXxiDffmJqrV2uUh4gR52BInxMsj6O+xO4Qs5nWSzN6hlqn0rYFM/QarAkYC4EDED2xoxbbT
v9gfdGybi2KHE97Bfx8fnuOH7I2IgYVTHoBAUWuPGGGnbmrp6nUQCUyn7Egt1ITUxNMALsWW4Gsj
hp7aXmUpN2g5pOslU0l1nbYbZXSPSffBxK5ZcwbA8CE5cJM2TJI1ZjrbTOn3wMYhjxKXzmldiiir
TQJavgTNP+YYPTk6EqaRPQ3AytPPSAfx4k2Ra7ZRp/pQrrPny6tZhpkaXD6iNE+aY1zYo+Abccqv
tUL2TcTFL8hlJUQUSG3PvZ15EQX4Czhr/r0rcGewW+GYAWvH38G1lkZsaFJEOgZ+NjkPhw15qBcx
rfm/GCaIHbDYhS9/MY11TVqoSrF9puaChIEmHhERX33WAjHg81fHk1cS4d7QXozl/VTjhAM+8r1Q
3u8eJoDvRe7c4jHPyS/xf1I5s6osZgzTJd8wCCpzegjBNB/RcWlwzmWn6CvsXMqNK+uU0fqSUacB
AcVympNU3h2Ur8Fwwtl+PVbFENy0nHk4NJjZxmsAzMW5lfPVBux5kjQRRQ5PorXrO0hgV3AMtBsT
OP2KDUspY52Jl97IQ5yUhvvuH52Bl3WsGPrsNHZDfYrM+/Md4CeM84CVT9m/zXe3dTqyF30tWx0v
B62FfdRCK4nhqu9a+fx+1rJIxqZrrWc1Qjj9944EqgHfxyFW6fwMihmTC+8W+tSRFnJM41DohAwO
GoaScztOekV1i2O3tGgXhqq623JvURj3chy4HTq3D4IOmxDFeLiO5QZlNtscf9ZheRzzjk5FJbH0
+UrWUbgcHjcM/p3gY5OOK9C0qSeC9YgXYUjR04ZXpfIE8aydxOWroUJXMEUXA1NqHqP0Y009QJdg
2NRQWiuhhp+uPnfuqdob3GTCDQ67J5hBTirdNOyqYmovqOO49fSUbOJ18UGM0R6ZCFb1i41Ik8tz
Ss3BKhKuNt+CX+/EcWWqFORx6uCQC0RL4tIFhGHdVfls4srYMt3lBhutgNYZFNCFa4VaWuUaBlke
8kkk/q1uW5UMKdquHr0l8YT/l1S5xhz+zhT71mzQ+GDSXA8oaBJnOWumQ/NDzfYAiI7/BlpV5Vsl
JE+BxE4ek33L4eUKOSl0g/HaR4hc+UvDSeMVFL9RL0Oy9zFAlgzjQmfv1twFD39h9Mfz0FQhct8Y
GSxB6LrdcUSjnT1Fo0wFxgQU0X+PYTpuRE+XqMVT19bZtGBM6rcTMpIbHW26nhOHFXOp7W/GUoPO
ZVgRMa32p+WHY8yZMnj3ee1Y1Tbrlsgm05dgh1vzbxyIxRDkGS65OP0J/PkUnCbIaedHX9CW9lN1
CsOu8S44Uuct/7MJBmqK4GKU3SdYg0NEj4ejd/4JOzslfIPqgqRZOWk0HD6PjKqsKPhqWsRmJfUO
9B7vDYlEzcUAduvJEOEgYA5+BLby8cgXRn/nqXiRwIIT+mValDH2BlteVrM4nhzziaF4anu7Neg4
v5c4QykC2QWp+qVe10H9/rhn3P3v32A/OXFRGkZ5oHZXrvWnFZEBHIBo9kMDobeKqtDiJAtYAKkH
nReBzOLO6q68SVAgruQPvZGeQwDdW95CFGKhA9uofJoYoniv26t0/MsgWuvqO/6LkgGlnfp4XDIw
t2TDRTW8Q+oT2IQdjpVlctiH44usPIE5tGljSzgbcu8qADC5j0PKxW7sdHf5ftx3moqR36qXnl5O
IOH/x8Ua6ixkfy6PcZWCeRyYqrtNrJUmi34msxVy+FGx7DADorLVqApx1Lgspq9Krq3Smn1VX0Fo
KZ0ROlbTH2b4MP0mO4HhXdyN3oNCP45+61Pg4LBKkcAGj0vz6pG3sKyW0akG0kaA93woJ+6wNMsm
Z2+RZa8FTg6FXDH3kmd16MN7AFlK5Wvnwy5ltSrhDDlyNWT7H8NDxc8oN2i7IsDLlJ5XgOxHCBx0
aEZPmPkn5PXCe8lAlztO/sNdQQs7lejEEY1iuIynPXtvu8hfR8e4JURJmnlfwcTMhGSjBrX/TUQt
B9/9VPPklu9V4XOEcsqEv7uuDCiXpXQK1jNEBKKsvarLLj6d5X7bC3Ie2targBp+eS7rqNV8RATE
PWk4W/ksijHNRT8kb46cw9dDtiKbj3/4IvlHiJB228/eh8bLXHLA5aczGEMAE96BfaNhZ77UYUkc
8ZGZckWNR1vf/vu1f1TJ+D6BamWI8xnL+NvmEMgPWK2wysp1fpbzdlc3ahSlp4om4o7Sbcw58VVZ
XvV7UWM24XM6MDWQ1r/a99Rmyfxq1a3y9XnbogceaAT5Elu52GRnAIYVU1Mls9pCu9pxVg4oFLAD
RwAgdkc18AtGa3yOhe/Hs2MbuVKe0Y6Mc9YcjQt77hhJLQhY1Oxv2XVx7Lpha9+i1DbG0unUWWqk
wYUSLMECFAVXYn+hnLAGfqUp41gOChFkgWXDMDiGwNZTfzZmAfAYkCy/aYZesCM7HTZLD+3XZYP5
1ozDeBRcExmbs26iNNjFCZsMHWiq323v9PchNvYxDLelAniFO8XPw6MbDC+KJ305jHBZeLow7k62
q097LLPKwIx0XT4FupHXXJ6mihcjyM2RFP33v9Q6ofclurcmmaQDIyRyIGhNjVsuKYP6Y2mCwpCd
PBB1ykY4nfeuGzX8RxS1uaoZCSTDYs6ndJcw4UOmoFiCTK9SJSSShTyiCeLxnTA2osT/nz80xdyN
XWmnDIpxvoylDTHbSFXSnqECdfnj5jQL5F1nX9lG7C+MKCLcPhqEnsSzMVb7j2ph12IDOMOfCoSb
RWTFaDTalgCgS1PYmwwaojaC6CjWj+Mm8Jy/v1sVwmeajdpvkDqwbwkAKn9qn/LCzKdooQZY4P2W
4R1Qvz52AAWdB5vR5vDFOQXLMzJqK4ImWBPpHbBrHd8qDjJ3YO7VG2y4B+X1jrPOzlXH1YUOk0Kr
holhAQ40nn9kJqVbA9KSJLH1X93YTmPc2WhNoYYqzFHcQyNOj+i/I4jD856F5feYGF2pAuAJMzE/
HFKzuYVP27VQs50UMDtiooRUNtfNS6uZwnKqTs1vou+ldpEPgE9jAzZ3wnnDyUOpWAXjHGA+Kw1G
b/EhjZ0sz1ShqhQLTrUjzLxMWg2DYHiXWL40A+KDWAbYJsyFMrHZCz+3wazvO+qvSZTkUqNPoNTp
cTWKWlEyzui41eXEKAKqKYQJ4JM06GLxLnwDMAnUOD7506qRKDIRkGSisPKuG1+nhrU9R4BbyCTE
59HIPbI6Xt0sVBVmZ+U/U8Q5DVh28D+s+qknVPVx3307gcnvHJ5ltcSn2bXQzBlH9Ccfwv3hrvR4
0ukbpYx5dfz/DqVymDLx2CszcZ8SbXN2V8lQqkBrnsVlyFfV/JCmvI8vUrhE5RjUVfRZN1aTeUnh
xqC0ikwaPB9+2XFL5YeOIgnvZFcQZMHGWiH9Z11PYCyVkXZt2EaP/oS5UbKdJ06oYdTsFCRwSA9P
6+2BkotfR91YM4vcXYqIFx3kFHOL5tzbLb6pxr4+HLiEZ30v67mBiZdQ5wgEsR6fuUDvHyPqEtQX
U2YasQXueSBgymI+zJnZBPNmaB3Ym13ESKwzRwjtRiz2apaOgZ/4hVzgdTeS+3LiAFXeElmY3AoT
LYj8xV+hDQ0L/At6pSavGeKJI9nxwPWTI5nPQgdBrxXTTtFDT4Ejtf7bWo9TGBCao8/ZiCPsl/0s
V52Kr/kidqKjEaKItyLlbJ9+rX4dNyaBCLIpcf8fEsobRsa14VoDrVCuhPve4C4tBfZRU2tvoMAm
ydzMS/fD0CZqPRSed06BHewct2nOt64rIOQY4yowM7CGUG1k2VXy5jFMuSDsmoRFJuqO7rYxh89N
xgETO6DvFvJO1ZWfSVLqmsFXvjTPEnoAvmnCIcwe7zPacN0kpYDtfp/wedAFCvKiraJujymeC2sX
O47cEA3VhvRWv2fWciS3ZDXLB6zzD3WSVR5jJht1882esHHFL06sQaEdeJWNYt2bfe635usVPW+8
NFy5Y+lN1tjKbodEmquS/ieX2TOp5yhhe70eVR7DcN2ziiQrl/ek3SbeRM8UruQcsAJPDtdGL57s
RsqxXsgEEO3Wu4/L0HAJywni6Fht0GJ5dWQmOu1CQ+fooVv7OT3yxjIafg3Qogde7m8HHBd5zgbP
L17jqlMzsBT+DlqnfKl/pmIgekfYErnRtvynngQtVyJjEl2h9oOiiaqAOrF7UU7EKj7ZA3LNPaTQ
ZsY75JQJ9HYyk3XCGrjzrem9KpT66nA/fEVSoT40qjUaCs/48S90BnySMsCXIvinIQ7XrODjsdVE
Rt40wIkkNnoWPqeKYwyt1lPvt/puXY3F3ETYjfBdjYME9Ot5ox2iL6CN/k3iXJUGC+QJ9+Es7DIy
IwyGc4URzNP8eysh4lbtnCmHFpctZJI8EAh/eQkqpETvVOUiYXqFja03Spv6TigFoDcaTkujFYjO
9gQv2sda3o7FB5GVQ+HN3AlT7DL8UScHMFhHKUuY7Wj/oyUvt1DE1SQ6WmsSh+RVvrFRQObMig/G
RD6OF+GEoTq84gugFkygvnDSJLO6pqeHl9hDFQq8c6lpce3O9QBTR9+xTSjYOfBW6xyHzNmBehb5
YrvZFKMiJVZJQXt8iKYKC4WwIZtrKFI5jhgq5CMdTBettADc3yOmvT5uetrkEsk3qOSMB/pPmuug
m3AYn4MYDJefD68135gyKcjgLH8eur23ZgT8WGWIJIduipc+XpuDoBi288ukeLlyI79qZBYt37zF
34+QtISkyqcO2v2XMTuf7m4cfRJWVxQD+k7tR/FFLPkr2mk23QlJP/81CPRByboBMszPdO4bHCrT
W9V2boxYWXOYcKSS5vBIAaJuXC2lvDHcb51xMHYI2XQVulZir/xulk4qmFdHW72d/KWKjJWv1ubN
FTO6sRl2POqy7fb53d+q6OSl61zq0Yl8iXD0Xbt1gV4ZHry89ofAW7EUrO1RO7LVa36aFcaUo7BH
814sfiVHoyj4TXcsZtsueeHOqJayuNke+MerZ4fCaM+rLQYN+f7Oi+APJFvpYd8D5Z8JJZ6yF4o7
5b/8qbj/PhVHjO8d5q/lb4tAArRVR8D/iAurVLrc5ugtnnS1vmdNRO5amaC9sroDQUJF2o4SsamW
pYy7MQQQKvI4vjYYShxykjPOE653zy0ny9qCrEsQS8KtC4RiKck5d7+E2W+b4btjr5FWrRTbOKE3
ORiscfI53G6YFbuAFND4fIPS8WwZOkwYQE6w0XROgI1m74xZeYau1e12Ac180L7huOZvpYidbSVt
rI88u+L9y9S+BBkt4rgFhI6i6Ne8UrCCXWltPV0nuS4hoArSv349q9VR+Hu2TganfdiylOQ3hBsX
7mLsKKi/q/xkV+O/8hXAAe7Pj6GFynsQv2vwRDQAoOYMdd7qy4YXUm3sRoILL0sEB0E5NBpt8PI2
OnlTxvKUoC6LmoJk2fvhWXN3RmiO0SRncBKI+cASAt5ck8sxkoCK9/bD+uIik1De5/2Jh25UxW2g
YX458TOFTuWVDtg6JV0qJ/3fvvSbFKrHd14vj2Z2zG3cSNTM9nS9LY0SjtV0R4F4wiExAXH3fdNK
QcUpPL0dQyiFk/kpJTU+PkQrl6nB4p9KJ13SybwPIt9wL/JMMFbrs7sgH6us8iPV3s+FIdLRM28s
jYdG+ES5ymLATRutRYrQOsrX2Xi4Z/fHxrKkAvgFlxEnXI6h741MSxwcBgGU6s9niDzbO3hchHMt
Gh+0Q9QjtBtHfjEhPhFA1zlugkjK7/qtkozr/Ie3K7k0u+y02b+KtZY4Zzd9STtg+csLmwIOdgn/
0/9e+hjchOjAmRXtHEiP3kSmk0lQ/U9BoplyXKGIyc3LFVZIL867J3GBoU1+2Q+6U89CfEPNTaws
HuILhiw1blIW9i3ySeqO09C3COuiGIkTXrHCNbIrVaMiOPekA2iaoMoBiW2OI5STrUesTBIY5nUr
JZoK2wBjidzhFJCZ6l22d3V97y3c18+uiqAwSXw4MX6F+L0QJ+I6GqrXcbsZ7GGQlCe4wzc/WAd7
UuzUH9ud8TtMub5vHSxdKvdXarmYuDy28Ki9qvGKS9xlFVRqThajjUTE9N6V/7/tH6HQlqlo0ROf
tKbOtLmc/QfRCmFEMglScI0JGf8rAatlaCI+m4Aqbd3T/zWwaoQ50bTgeRVIiJtfF4c0r/2j+y/Q
X1aKOEqBtK1kG287Fzsi8odo2a9lCbwxp2vtjMzaKGvi0bfcfowXtyphd3K9VX/hGf4uK2L0ctQp
nutRXRxqjPbTzwjRIdvj9cMX57tUqR1inN+kN32nr/nwddNX9yvNQCVPWiS+7TZVBpsDL7EkXoNU
DG5jwbj3rOXQPeWfaORYru8lY1bflI6iahlRLO0Urc53TZooPGvOEotWC0+F5XN+Ft4s5xRsCxee
fNk5jAkKgM3RnsdE8V2uLx7mMZuMHapZZL4mZnLonqAUOgG7Q6KJYW5KswbzmRPjhKGfMX8i/HSC
Q8BTYX3NxINOzOe8tB787LW4PMPLeh/qvkjcDJF3nynn7Pv7sJuW7q/ep3Z9R+KATPdA/gVUf0EQ
7xVilQVruhHJgUwhx2ufV1h3dtUIo0gZyyEBfXiCzKyUfYLw+qGlmNVtMdTaPUFofS7pCn6OQHNM
zEbtrbmK0noHWE6UqZm3lncwiuBOvZDa3DzU70kx3WIphLdXNLBzUoJxd/2ZZ1V5PdiKddwVBcTQ
5yWg4V0T4CXghQCOQTraSChrls+RcKkczKWHFhG4LRDFhcI7stBml2H0RP1h8jZReHu50H+E3fFr
QWEkPXg+ngENh1X+EJbXKlBNIJa/J7HcCIe56L8Z6IOFK2a07A/Va7Ev45GgPSpDADqbggMZFPU8
lWz5DdecvkfEkZnMRc3OMmpmHCbOOvKwptKMVY7zOQOCC5uxZbXFg0sbXPaTXLcyTmmAbkc8kOHD
tz4rsdDuQNzFNh6Pi6aGegIdpXUL+bYnk9PBAn3nKML7g1ZFsFzGj4+hMHHonfsbGXPZ3T+tTeBT
riN6N+ymasBD3l3MW5NH2s/x/CyFqXZMr2JUs4UjvYr4CTkMJpjFaJa7YX9UWwtgh14/t5PbWa59
l76fDAi4rVRnCSAvxkFYMGg1EC4rfVXbPKOq/4nckYV+YoGcXiPxhHPOcawm2jA1WcQ8lDWVmBvp
X9n7qeuYETIObw4FqfgoYXyu22iKz4JVclLy/3LMg23DojgJS3F4h2IkBTRKqrHToy/e0P14/ySf
aErA8HdShvzdWKxup1nzs0sp6vFBWoT0GDSvtAs96YMR/ePgabNMGt97fwwP3vDdhY4tCTbcDE8L
IyazEXikd01vAYeZXYI8Bqg+o1or19HfwAcXazsLhYlmxPuZh0g7NBff1zCzhjMiRHJaFzR71zQM
lhIDkwLON/RCSmF2WoL4HwAIRAFZJAWWNhktcBxzKtEf0RK3JmpUrpI/We7fR+lpsyzGUb7W7wOc
sVeB/L6f6EpPCBM/og6FBP3Arkwxu6hc+PdBcwXfA0Of+cLq2cYG+JL2nPw5lPR13m+HijIpwttv
EVsrltlnXNnpeOqc3l8dVk2C4oj7TSrDxTq3u9v/KrOlRNx+Urq0Nx+KFuuQccJGYcIlnjS1TPg0
LePtVr999g03zF4DpW1eZVkv/IQzQ//vSsJbOzR0jg2yCKMexlpt8LQgdc3q3A5luVEsr/3GKn8d
z1ND0CuRTXtmkNWb23KH2CWkmI8D1reH1W25VHXZ08qSji2qgrzbw22rnjZ4wbH7KMKoMKa2UKdK
Oz9afT5upcbmUI1adzfTcYKjbXGXSWkOGa6Dc3DhL9roqjfTPsgjA0qN2T066ugg0xY1OUvXzTz5
aLiOgfrz3kwDqoqGsFzrEVRv6DNOZeMsy2DdNaCxfMjaFCtdgNwHDdyDMj1e7xmVEqYQMO8oRBfC
ep7qHmFRpoXk2MMDQRXk3nWtxbYPYVuD1RhYK7UE0RPF6U3xVR5IrgHLWbqhYKnmKPnRtWhRBqGa
SRb6jC+qR7Q0Gv555n5dIa9OALAcalqHSh+AIUDR2nXTIOEwMtTx71AhMVj2pwD0zegnH8iXl3a8
twBfeaVovwdaPr9E8j06IdsPeaoBRfmteuX0l5UOIidgqG5QMvWCe5Ykmv+IIeRRB+A5Tnae//rs
u500/REW8u6ewEfi31g8z0ZAfvFdvLRFZWVD+ueA+cVfcVJ93MDQdXrYUO/nAd5k9eNI3Tt6kOFP
/6moG1s3RWFXXxQdP2EIHlEp3NwPsRwpcGUghWzhp93geWDPOrHWN+pe1Vba2Au3558UW1EGY/uG
0VMFwgBZ9RRqV+P6XOl7TYm2+28ty/cynaNvVoEl4bp8NcomT7TNqPQj/iKzxeOERc8P2EvkqY6v
3RFo2PTMBqfGu8B45ucajt3RJhXY+JCT1hdqvVDyY6Rw7k2Plneu8BadJX0FUbmo+aRHx9ZRCK/D
k7JDQzQwFs1XXvta2CVOYKN7tEOeK7okrw8brY9j2Y2rfOnWmhgr6XN3lfRN9xyEZBZjZuKRS8pL
dtojQSPOW+I70Vh2+zMxCdaZunGgT7yiaYulacy88dGUO6xmO50js20a2LqgLDdhzVompG8DQmN+
eEUz9CEgC2lRxUklMWy+4JpgBrVpt0ld2fAz20lARlpJ8wl//Wl2cKo/KNPURpSAvWjTs64/fnci
Uz55Vd7Tc2ra161NTs+wGxEKw+5AprWnHUV2iclqMSWr17sWRkgNqFlhAR4daeb4RcPevPAgz4L1
YcNhlRv6xx+KWbD3us8AAnnQSsFzITjwYfgRfJWOBwmxSyJoFLYoRVXdXpSBcqi7am+hsTPN0Fdp
3I0ziGiy8w2+dWHXYapNN3jBWQiGk2HhfpQWMvoI1jxvW+jm2QmzHMw46rLTmhvDQLuyHw/1nGia
rpuAAuAnMrzOR0dsmtNPcB1mELGVCPYZ/ESWcy09gls9UmAP/XI0FlMw6dMYNfn+V29y2pqYEuZm
qR5V9cx7Il8WGx4jyEMmBNdasBQ5seoGgRz5SsHx09v7+gpeMable9OncRCEZptZ4xtVay/dC7wn
g356bQ6BKsd/yX9l1BJ/8972Ku+6tD3c9QNg4hJgGCzkUuVfnOKz0yCG16O/Q+qiUg7gjaQoAYxu
3dC1Lk/8TegE4Zxzs/ntEJWPvy4A6/gytiCiOjixE0OGUPXY68TpAzCdO03AOwbVgiTRKw96hCRU
zxS/vxhlvbX9/PMH0Q/1/ePsC3a/AHENqZuBfJpjNeoFUboEkOed22Q/LH/02q/TyyZaV+taCdPc
g7/7TpTOf70cLJmolR7qnu6s9DpTIq/hb232JaaKllWU+VHbHtC66NvHHkkEi/Tu/vG3MQOkeWaG
CVR1KDaGNNm0cU+u1NXMd5aZkMtdQfvWky1fSh6FuQMwdFS1bsOY4ehvRoplO8LqLV+zjtcaxh0b
Jwm4R6wVwHxI3o4+EXp6r4C2kcgS5Fom+cKwZV3wGYZg7hAxg/+XiGSrN2l3Inzhr2NKJAhHNpmd
othWTg9Zu2W89k+1fRMjVQsWFOvnX6RAYfRNrSvcFQIsIEwnBu0R83/KHHNC+Z2Phz+VIi9L6Za0
8hBNDo7WVgnmloe6HnbmMpT/abZ7sIhb+bZj9RiqTVdV05wHIvamE40dyVmes8PivJbVcAlNNef1
HeqMCRcan2n+fQQZn29s6IQlBZOs3viqMmq2nmcLwfD9VcBBDGCCWZHEUy5rYB2uLe4sM1CuEwJ4
9xyA7bMhA01lA4fSabqY7M0bnjOwDG1H1t7UBoB6JctLPMR6BGn9BsHAI57pylqBgfylZTIeGCWI
HWYJvR6fcBnZlreJ9sc0eseUjeGia+vsznPgCkDAcz651lZE8jgFdSeI6JznkaxdjtPiZmEM7OUE
I2lYvAdfRZ93q4JPcP2oYx/hnxusAX7xIOLF9im440K0QKhEUKrryvBI8Yig5/gVOlWovInx8H5A
b93NuUnf8uBsD6Ej8g1oG5PwGudo1WRQPdKOcmNDv3gd+zf+ViiJfv5+pkmpzpnAgf4E2Sc5fu9x
pfDvtS99n2Q/mQTKFMYMihkT8wIqZ600eSC9atEgKO1m1BmwgQeZlYvhdf65r6vVgMqOLo2Rhezb
+xqQWbvoSSk6AxxDlHZzho88fYwYaV8hTNdgrmHazDQSZWdhPE0yNaPflPFux9fxtnn/HFkoy/Rf
dYZrzxJTjGXAwKipL7D+FmkU2zth0XvLRH4IVwFGsoVfYVSRmuMsIhf1ggbnS8mLi3NQ4moJQgEI
PC99VlBsVxGYiKIMu0TNL+D9KFRbMiv7C1gqVgwZHwmq8tgNlPNP6bgedmhDXGo3cpksV7WzkMQw
rQH90E8SNZwD8EdEhFXsNQMhuduAklH2/QneXdPgsSGkhP3iNCIlHtH4fvDHjonz9icsJN7+Va9d
zf8l7oJsI8KSxBNr28xqAJ/OE9Z26ilc27FWamleSVuV+/cSechEz7fyfxVlNN5pPKJTol8mxlgU
5YbHU6aIaudOcOAAc6DO34T5HoFdc6dmZxgjheYCKkX5VxX4cLcbvFPp9tudzmcQ/i0YVkMWZ7Z/
ZeErWHC9Z84zapSjHzRy/JYN9xBV/hXIo7ijtmysIR3xNDjJjdOrm+qrQtL5it2cQLA3zGNfDjA1
gYwOnjEec40kNjlo7w1FldGHT/cHY7DxK6OIAml3er9UObSvEttXBMsbF7TXLiheo8Z/LZCkMyAo
hSCcqMcZ+LNGu8xGBgHDayUmITKmjulyWKgoOYJjgPXvHKKxC8DMgwTELIap934j2EerCcc6Ko7L
QNPm2gq1swGYKGomfq8doznvxVSXbc9zx6tL2uUe03oDu+mPDK9rMsJbwZwZu8LKgz/vCS5w2dqd
PM/g7iWvbahBhmNkgONHJ5D91JrhOdecZGjCujI//66wVnT5f2RPS7VTs9lGwFB1zD22XpxGNqB2
O0vYpJQ1uWTDZJleWVt51j2eKA5lox+AKlk5jJouIE4/dy2+8CMzttDAJP9WzLVitOvRTtbOMDzC
j+5MIAC5PVtWvS/6IEHB7TUzvFL92RM79OBSGkOVM2sATXMSImmUYgN++0TdDv/NJC6Yr7mgtg5w
n4ouap4rEAZvdxV4MW2jnr+nn0cc8niVzvkIQ5kkG/h0jHM4MAlfd5QLe4BaSLChe2gcJvsBCv7M
vGBh1KFJdFCL2MYibRqJi8q44vXPZKJKuE3cXHtkSBebaPJqyA+u07HOfCcQh9wGFeN11eaj25Ry
lhbALZwfnISPoOSjPHMzIvV1JWIdVV62bsuiw6QDMwx1TgOZladYwGR84mmYYLQDjPpj8BYPhkkj
3XIYJ1q0F5gLGPoC1N+a3zLmWC41nK8jFX8D39CwhWhDfVkD9ZPGb2yEF0xdI87X/8G5m73Vrnfn
V5QvJ4wEIdkCYLAx6WWXY4ds4tkur8C2qabkSqzbdLiT7aenLC5FOQdNAsd2mZaoh8EMFr4FMR6k
9Gm2fjGoOJ0SA088wyXlXpA3Lb8kwh2fASOmksNuMaFt/lIaSrZrJ3mBAe02Kf87akF7RUhXM/rb
lji/BwFcg1gJ2DI4bGrSNh3qL1utD/sJUnWR+u4ab3HfHLzIV7v0dF3A9VLWzzNnYblPzBFi/6Mz
n4mAfFlVUvZF9nGWnT52O4veGkF28t06IVJQLwM/KN+vXqfi1ZdEk3lUkhVpfADzbmWJeu2YgRQx
gex9XOwyTv5qLP59D2REu1aS0bedgAn3yO58fpOgjUJTD+cUZYlBjUGgk1Uk/ITnzGD0pYyTq8Pd
XASucX2NjRRsYH86m9vf6WL7jVGmnR2NGTG99M9F94Ef5jlwerM9Jx8hUH7fm6cL9/1U5RziB0n2
8/D0BEnLlGDyukIYFARmagCBB1LbPfCYLfrywvML7b64Frq0+91ABWVj/jEkAee/KITDUOiFAy17
1U93/COIAXzo2FxRtPkqrUNsHxkiXKsT8pHe/jDPn4x14El9g2cG7amkdVSTahLXBM7RBgwmZlos
XbYLcTnXA4HK38EQSkBwknAoQGyFcz0qAmwZwYtvwLjDbVwlbKPMJH/1e9aLXFGbqk7xl1MZn1iU
WM2YgscYh2hXioJY/4WxDuz85DvZeIJKg0oenA8ZSlZK1cN+/OMG4zrDAsDvqXj8rEKm5PlG95xC
454ZqGMqgGPEvvAA1BwZH6VSCKS6r7llnhfSVOkMdsIjTgaBQsKjeWBVLOnxJz3HqJvXm9TO9HfX
MaX63JvV8mLsaWrjl9wDVTjemvbQ4inn2HcOgjFqx+KMPr+SuLgpMK2knjHdjGmN3o/B3hBfzr8v
sHHBXZnFhK0cW+z2HL9xwlXtVL/rYzXJ8EWwxb7r7V4TfldHriZK+UmHewH8R/cANunpSCkWt9q6
ldjsh8ssONHJwAyCYbT+ONsJ87mEdCxZkEw33faz01vCESP1MZuVlIpWB7DY0bBEphnyiUOQWWnS
bGc0BRlBBZ45CUJa7dzTW7DmU3WbTJwJq1Qxti6+YRrKerUAa5lePCXTPkm/3MworFIh/nPOWWWV
RMR7hngN28URMwEBchELbvkTdVPzSHQ4K1XsG6SNAqDozbvm4f1oR6h0nzq7CSxhIEpMnYol5zF0
UOqNuhZH99+CGKmsPwkQbUdNVnfHjN6v2bdw5jzdKnlAVCGE9qYkmwEzH6tEkHAJdVfsxYFs9J/z
qwyhpLVi3aovN0HJAcCeZxB1/4bPWQREMFo3F80HW2+FH6Hp+vJlOLkd9zlCAle9cT/U08InF2XL
/sA2j+6AF5mRt0RRFQFhd765f7adQBgTZTfZo0NZHR2SJlKY4j6KtU4hEaHYa6G48RPNR3gM95fi
pwCYdtCkQ9nvIzvgfaHlU0vGaQHoUZQvHUEqBDB8MoicErnuetSlfgzlznjcShkv3X2TiAnXTsXl
bRxCP/IQ00gkVsdDhsA0D7BoypfaO1KpxO7s0TkOVImEWSyOSxCZ7QRO5DtuUcRE4rZOKlyATtGB
5AUnoU4iq8UZD6LOwFxwk0WbuaUhkJNf50RWNd5nlGpzExJ1tbW5unPU3aBnrBna4kQL6pbE9CRm
y35o/muq/Z5ve5aPzNE95n50XVhmKpoGq4goOdRpwRSyyAY8JoGpt2MpIkzUxXK4XqdHlATxANvK
rSKP+2l9UcICnHfFDVR1DXNYzAXehW0+IlSGVXaScqC2n4AtyaP2mU3nsl+81LyciGltM1AJ8KfN
LhEHe81ErJrLEy7iTtsY2IsphC+Sql1q2if1If37FoZQGf8NOadzfE46UAXIxhd0yTnzpL/IM7DM
vPQK0s48++dSS5/EmT6FBEIK4ag+QaJuDS9e39Kn66dGHCHxhmSj4XE3j5FyE9u3bCzahZVWArbh
orfReQGp5bUNIREnZ/DVeWfyBFetTXHpZFWkgIZ5NX3wcZvwFFEpoB62SQJTlGtmWL9dgFFp+Mfn
J8bpGNI12ery1+W0B4TVB/Dn+hXQLHWibA5dh+kbroEDOZczmRNINqy7+b4CGkhIYMeK2z5+Ht42
Q2Ls1YqrF277uVLfIbMkzeGoo/DT6jUZabKA+WXjf2hXDGwBjXlMPQCk/v+uy4X0Oa31hLJjSrbm
QaYt1vFEX2cKP8tINK8eIoUAL1c8IGK7dd6iL2GUi8K/eGue3GipOCkB7TJU4g564IUl263zt/24
60ax47fwdCOD0UyZ7I56DH6XGd9UT/dmJCfALRFKXxCwTChKki6uTp4uvZpo1d42kr4zC5AJBr9R
7g48uApLhdXPBl6zm6+KcgFleJRiVYSp9czMadyLeXS0Nq2KYCbRS1a18JnsmWeteSi6VmtWnXUb
yAFPHyydJD4qOJpf6/Q3qAprd6M+OXkp7QHmIPxXQ9k8mkjcf0IJWB0G3hvXdnAN3bBD3oFqKJtn
8w+XKVN0MFNKpG8dO/3RbDAJSJoiiJI7sxGO+Rnl47LKXrGRwgWihrO9ZLDxuaklsBcikNklzb4x
Y9WWHqkpeO9jQBSW1jQW8lCFQicpouaHW+rHgs7179EBLKFL8MvPcxq97IFsmjO3Rw1z1fBpcGep
Ny3AeGQtNlXpYyB4TPJxkrSSs42fOqlYf1CnkWVnzbxglBFQCQNBVZAtaK3w9Iy0caUFit5cDohB
wDL0JKQWNgw9M/UOpskWhvpmhbysSC60b5DbZWCJ5wpEUIZbuQULcddOhXQU2NK8k3niIB4zNULG
95QOKztYARwRe/8zLJYFng/7noRAFTw1lRUWduJAlogCjp3tVHx2zL2eVXTQuetbi8nFKzt6XoXu
QZP0LTRfmFw7A138Lv48GAABvTuw0/OX2EJdFcx+NApFKKL+LNxpkp30i3wD4nvyYK+umq6FRv1S
ht/NjEABRQGuIHFCJCwb/jsQgnIQDtQ//HjQU1MV4u2WdkYO+Obb32OnxNvmwVSGF9FYV+4yysnO
bPkm4E4XRuThz5fD5Ezia8ueHdjhgGKwf3L6TiWd9/azIJ5e9IwgrD6LQ9t3MxLD3r75hCzgXrs4
ouAGHlVrIfl3dfnP7MKDJPWSxuqnibVF5lrhQsCLuxPwIxlHhSkllng7euaQFRXotlsWHnAnOR2o
1SCe9TaXjvosUGUukfuRXyWQoWAATPbDIZT0cFUFewAIrep7ls+Iyqb2Q8HmxwabB4v3/xrl2qHi
pN4NZ/Pwz6aWBfDm/d0AN3+DpBB32yW4EhFkuIg/+Y8I7Sgfvq1YIC74JDMtEUHGfTHnJAz2DZ2K
eYadmEEbT6EEyHq6HlW9DPTCAcLSvH4d9BQ06RuejbzOtwHaF3wxcztmogvwWK9WvqeSdvGvkFGI
jzQkiBBMHAYsVNbOcu1FA7uEMM8x+I7V8Wogq4bUVtCwIqYZ/MxxVAKs2b2mPtr7F2SnzRc5viWy
vHuFMLXyFl/QCPsJUIKUH+xdNejMkRopTwibodLzaxer4sFr3eywnNl2zxghkyIigVp2eXclamUE
SQtSZIqSAUO2AoN5rA1hq/xbPWjcqNKqHDLSofDTKLSa/e9dKkHjleLBXujsc7tuHwbNptP+AOh8
BrQ8Y2H5BN34qvSueTPfjxXAUysY7VOswUY4Xe83fHXfubchPiYzFtosK7l9ICQfmAzb9jT+SpDR
F+L8HgLlZNQMxsndTuE4DUDiRb60jyyqE+93wpg2fc9TlTl/ey14Ylk5l02qkSwoiYAzGALXMJwh
5YSB2NekEYW/Wjebd1RO6uIrAhsCUTR7lR9UMCUbMboVksa7EAxYMfBIXdSyUnaU063DJPN8/Dv8
I5Jm2SVLMackrgCtj6875neuwTbW1E+kY4Ha6jt+Y2ALxQ+OrhOPQNMOsJe9HyAmzhS9/qb0SL43
G6xj0ljYNMMMS1WdRnK9+EUrfC1wQ3kIjxM8rpTGdTjHFlyJ5iCISNwcFzT5AZIO8Zy50Px3V0eR
mOtE98o2CK7TV0Pkkx9b6mxJ5tuXhDbxW+8+SQ8cIxO9E0vLa/e15PM1Fh5z+6gMZFwERu9lXhT2
LHg9QV37ZUIux9JdQ9zVmq+QqMVmMh3iVytTD51zTKv5U+EUwreSA2+DvK/BW51pZfQERlgq81ZK
veEHSBS/53A4jI6BBnWqmESNJ9CEKWnoEPBxR+Umorlo9t0QSdXun0X5wch4cbheu5sK744aEAy4
pbyq8nrfNbD3LWGZ1oOAFPpDyO4oFZc9Xq8ohuy6pSCWwqUGnAyyE9GXuAYB+KrDl2wPKIdttpM/
FmhrQrWR9YL689KS0zT5N1MDhmt+IqTYvInXswhHMJksAxiuLcjs8mgA7uWTWx4bXWFl0lg9meWy
kG1jffDRNLNVWmoE/S3IMqstECeskHRoPhyByaxki/FspRtykkcnvFlHxfoaxP15J4qNajDPaXwq
5Z8vwHsvX8YLzhK0B3cRc+7mG7fH23aZt58rz/F+lHbduTODv5uiunVf3YSVklzTFAUfCU/W/UTI
DjsuAYA3q81InOK11qONlxpCtt6L/H6p1JSZxfdzYKyp0BSS6YQAQiTmnE4cp25IxrkqAW6OuFOo
KiHQQ0Mk+n39HwwnJwiBjzIojXpGGRvUI7ca6ps1qFZQQ4imKfH8QhUCPQ2xCivGbN/XQySyO77p
aLANYQKeXQHVpJBJT8JISC1M8MCG3K8fo1VptZAk9lTn3yn2Wc1Oj8Bt9u9/E3aKY4dYnhLRrB9o
Ux+D0woMXocvZmuonUCrVZBJEdUcc9GZuvt7CDTwOswWwChhhi/7dZ/Y8dS6IsL6d4Iod5nhGK80
SU0OsyxdE4lB7aol+eMuORZXyUVNjdXUfLO/xV3Ql03dUv+9YZ7m0njEqhRMi23o4mmwwQIIhhLE
/GhvX4ORRYpl4dIN6UacGg2C5WGph+LlU0zZr+hn/LtkEP1EmS8+h08lCYQXGrIFUHVn0hZSVW35
O5i/2QuuKC1nUf55nxxb6LDgephGGUKHCyT2AK+cwKztdKD1tP3ZgnWUd/w5jdU+0St/d4H8w9nP
U3basbdkSn9/n/5xHfKBMzvDdRw3TUoE4Do/hrqEOj/8UZzfQ3eyqQSGttkEvZsLZbA1MAupcAqL
kkEXroBSvIaB6GK8mrPjVl9jQqCwAmbjWXuYQugiu1IbJjp+akdYDl6YiUUiJYICfkQja1WmCBgK
/UpgHphKMC+v7DGGpTUZkpHBAAp9JoLoQnNRA7syJfoF89p5z4psBpA49ReUYaMChpAJP4cpVefq
8MboOaIrZmzVakuFaNdjppuSHFHCVNjzzmXypaLLQF6DsUK0sNSfVQg9TJQiR+BeEHFZeI+YDLKm
q4fEGeSiWU6PE5h9y0qKkuNCBs1R649WjHeV4UpYLhqxRbVKYxG2E6xSB08tc4S23wipl2xk06TF
B1ZCAJnCml3naNJwq01TZLluVrk6l1EzZZms4M661g51/Rgi14SwCQJ43Mt6xhotI/zfhsD31rhB
v5y4waCqDBEwph4+JHrvU4pOH0xXeoN7Wag+mjHLVhtVj0beQUok6cGIyzQSxfcH74fMCbfWO/Md
c+WYqBCKlJE9ZIdE05Un13zkOhQZNfmXqOGNeSjAwFn+lYpTCwV3rKRYtj3sF01TAnl+cPQaSPyV
Pbu6YcUiLF936e9nkzjLiJhRHoi692LsYjb+XQ7Zzo1GTOoUp0lhdqcyaqacaKjr7iDwk5NRWJVc
igRi6UQT7h/oUQi2upZULXrUDEOq6WqfC3mugI7Y6oJsvbwpTrmkum2djKPOL4e3pn1G+jARyKyq
+xJg9WR4lcnKyBvEJTTo1UaLxhOPySwguxuf86au0mjOziRQHbGfD6IoqbHAKCz7vFG5CAR3Rybd
XmgXwR33Ch9Nfk5grwsTGzY/Hz3xzGoMqiJPTliRlu7U+qCiByOd8NzXq0swiakfVtHwvrLYusFX
IAohD35I2AzK0obFT+b5j03ib1RyNAuFQyA5IP+luU0bIsdJLTi9EZyadNiBx3nU1N9dDPE1ZIYM
UYyoH3Ekg8yBd+6AQO23YnjtRBfp7ZiJBzgj3dmIevtrdtOJxw819X+XdmxRp35VzsuPHYymwsY6
+nRTC+ols47IenQMHSLjjUSd3gddpm/zvQKUk+743bc+5Y9813o3+kCXv6NdHlPuQT7RZ11/yoZp
nmPLjZ4lD0U1e38RUy3gFKDR7BsFKDNgaGmusQyJrVygNWPsuVeJRdsCGQy4fFegb1CoSsvUyYoW
Ve5tQa68ZNiNBzpnsMQfpJoZpImo0CkM6qYeYIzL6K4C8NDDkIp23kDpKGOc3yTXB1f9clH78jKB
9wSUC9pRTXyS8OE0s6bgAxhos1gKloKjv8zXMIYLCVKr5IT2itR6j1HHJ4tFJ7UB77DCr69+d/Dc
Ahd326URzUJdR4bQw7Vb86A5ECIj4L5QTcazmBNwPYA4eHAFAN35GSD6nHDKL6fQUQE9iY468qkw
s12bLBUZvbuS/BS3xALuh8PaY5qQ6RElwwg0Eacd8dxYUFU2PpX5FXkyE+EPfxJnJTzg3XoW9Q5z
rmBdRNOlIMadIJx9nPQWRpd7AjASCCEWujzu4ayaoMtTJUolH2NfZh8MhFq8OAAJCdr82FlDrcMV
qfjFWr5fPcLZRT/l7sEZymOfQmPSFyP4k+3Sp8xYmBfkLwqGiOzT4kAWh7hyy5vPkfmTa5cBg+MV
rxBZkf5yLPDmh83aW8L0tqPF5pwgYfBtpHlgC9P4fXvHCKQVuJAIfBhQFe5O0IIS20h2gT1NwBZ5
zV4t0hsfVwSAfr6N6j5fZwjwCR+wzBNQ8B4AM2Yw6pv86j0lLTIRQi0KkP0tumVmp+7zYmeIZMp1
BQFFehMf59rtGn+YJFt08zHGyNyj95JudhQfBwVx8/BdBjNqr4Kd1XhVMrGEpH/moYJ/YMxRyyyR
PT+5/lJ+sN3Bmb/jue8eL15eTV98f4xexmvkvX8nEYM4Bz/sNcxAdVfHHWdzE5vYnjO8XFTd7usa
dSGqE69zqNM/SHn5R9EIGAyd0vfwSwMZIe9zBk73qmlVZRQ8PAKm6MK0wfqcWSa4qt/kRETAJG96
JGv0BIOExiLaAx1VykM+kdcvAE92e89m7lXU77JFYqf3Cc3rN3Yb+Aw11RM7QyO0p5poqMt+sO71
m9MMHYE3CJ5yvEKIPUnScfwDNT7W/hAdgegE6NUnD3YAxEtUvKqo1vQ/WthdCn+jlqLOYiLZXdRV
A3ycspC0d/CFrs/FQRN2y+7TFeeaNyHf0LOwuSwOCCXdKPycnif/uSL4XRSwBbz81s/mQBs2w7ZU
YXVesCA3I1cqheF00QzCAt8XrDgsOXyW/qzlNHRuhWv3c+mGNFO1sgq0XcctBFWxktob8mT6XR9n
x4C1GbxK2GGUjFcc3U92bSF/gpgNAWE9oNJtZFmiKjpFk0BTSn5FEUaB00zBOO3buVo8l1WvgEz5
san7mdT2pQ9mX8owcYIGBhlYW3RQvmqovqsGehTl090OK6phG8EWIAcEl9JZBOW5UIWEygFV+nSI
LvJ1dYN0qj7IQB6hXEIhFppzcT2YFgHHZi2nFoUfNFZOEw+MK3QgQdJOUL915tYVb9AOwsWsRKIm
ZpuTjJfhGHA/C44r0X2Pb4Dy6+0pSsAjFzmeOM5eu2iPnEU7+x+jrL5N2mcbgt1Hu4Y/sm/FOivL
RAeluHiMJgl1VKSv3OoumKZbW5H+B2+pZazULMGZ3muz3Sq0JGo6dMtDCMw+aJq10zuiEcO6zQCJ
AOyrI/lPaK8SuBplAOpK3D8lmVk0fJmlo0x99fcMu0pQ8tEqSNatylgU0WYinebT+AZVsnnqpEyF
imf/ZpBHVsGRRXJXTSkWbrgnHv9WIby3/5ebEn4H/a85yr73c/AmOTZrAYtuNwUYr0C6aaMwKceY
XS4Sd3q0G7ymxEpmue3/ivh+RaeVDV2AhLA5WQD29M2YOupLH3CB429rPp0cJrYIIrqLoMksQkz1
aIRFdG1mJJkaXc7V9S7m1Z1ubXx0gt0GdEGdXZ3YiC0hpWDgH5bmhqtA/++76qHyzBVq2R6jGRvx
fBsYNPzdIccYqLKRvacsemH3pYpfOndgrofMMdtGSgPXowPSHUnBR3/Qxq6rME415sBy7vnYEFpw
HaRCDvAnQdv8lqsK9e66T7ZuXDTt3UHbMPoHQAYP0er05iK0xbk/66d1H5BeGQH5xUv0CAtNRzEJ
Av9hsI3Nj4GSZKRiLWuf2XwUAual5KuIgJpzec9CVCygSRZbRjp5XzZSj2ztwq4FE12rk2NcELxO
08CzMeFUYM2Qe6m6Oyx1Zshn1JMxvCNmEyJe1syoZBCsg+iMFGLl1lgWCJ6/o19TldO8x7iLSft9
IJAOPMYXxJwYyaDuBXHvXo/URCo16FOuHs6wuPvl8mwXKzqfPScXarNgmU6ZKjyfoZxpwgXrxWv/
ZJtN2r+lcGrSH4Dj1ZvU2P4ICjkBQuY+0ePjT4G/FgD5xuEIlzX443Lb0lydsGIJ/Raco9wAQVWC
joV31ferFzIOlk6TT4okB6zxFvDQ3SYPN2Q7qDdrl8zBUX+SS4I+HBr8jPYy7mUBojXzxpw4vGeS
ZX4qyV6tvZHSWuOJtr+7GXAg1k6piq7zac1w58CCRIu7rst9Jo4Ra+pUOml48ht+BZKryy4ZmDT4
ezp2FbP1vZq47Qhp9ULw676X03iLIOCNRzoPPz1lmRBWCmLzUk49Dhnwl4DFXxIzAXB/egA5XTTH
gIDql9UtIK9gYV0soSYM9W14e+l23pscpv9YJiO3osAs/Lp6Kz8+vDGby26+a3Ij8dKPvlMgmq5O
PJwiCdDm9LeVSL9JIGeS1tgnjfCVx81Q6NTGGU1NMsA5tJelNHD8CpYkGpPQeWnM7TSq8/jp4pKh
4QqTP4J2D1T10lWtVA9fWBtUtYMyl9QeIaoDFfXycj38Kw2pc/yxFLPAjyZHWXeO3KJqtF3YYbz4
MNgchgPXeCWukks5Tsp3l8K2U52/PztKI25Q5qozeqnvHpDiRbXiUe8J8Fo6RrFpVrT9B3TO95cy
kjKEwx1oIzZusFWL2EGkR7G7rgxYqEtjGww7f6Pxj3Ap1xlnauO/pyKOzCnDhIkL9Gtk+nh1vNVw
Gb3VFllGCxMj3yn/BZIrUZ1EUepgRsI0qZGJsipDIThtSZh9FZcPMzaC3Edz2Mm8skSOkSkqn465
KP0Ug7EHrYBcD7QR7quGTpCryxkWVzPJk/v4qKwPIsAhRfkhxxeoG/b4fH+oViCZyRQ3FV6oXDqy
LMzWRt+1JK658EEE2NaMYbY5q3m0Uq3wyFk+l3Z9YHu6Thfz8PFRd1tHaC23EmJaAeVaumamywLC
czYdjWrDGOebMhqHgYTT22q685BjIZxEkOvqXtzjKyd7hqlTluLQeRHetV1F0VMbSoIbPbB14JQn
db0cR7iUu04qkX6RC97a5HOi5QzXmz4MAAr5T/RolFI9bg08URXBHzXYCwI8pIAzhvj6w0kgYoei
hpBjnw4QUl6H2DvcpryyHeQy6lzDWn9+cAU6RtWZNCmKI1g7VyKIadO7P+SfwPyMRkcpYp2+lbfV
3GkHMoevAve3vhZL1Ch+vkxMLLtv9Yk7vS0oHYVkDrh6zBnwArpP20L/EyQ5wvY2sZEBW1XatJXW
zbS4J8YdVcoTUcSGmX9flw5qXqr9YUw9Opw67egJZLe/o51Un73jVnHGCR0tz248PDTSCwZlu4JM
RJr/VlMuvRky+xErre1nsWAV+3M6m38qvD24MdBAFKR4w2i4sUdv1Tfwymm4ExmU9BUErooqS+0n
jyiCZ+Vq2rEf68nXHw/MOcaKt9nWIH4hfr8HS3/XJUH2awEbmjc+Zy5j5AJWp4tM3cO3LWVK8cwW
GNDLnh8zrV34OUMkT/xgOP3UzgKWkafEQu/iOukKzVCs19WvF0/vGq27vDmlZSOzYjSn8tZUjJmN
QpLWY1S8YIXZGiknWs4g2Rh5bECJs1NYVgnv06x8LkhRSEz7CRK9mzxyOJ9rLb5D/WUp6Qh3QI8o
kHtAm1vfcqvVJjwJOlafLIzvPAnGMrkpn08lB+RlJuOWypZYz6AzTcVyD3F1tjciW3iufL2/tzMy
LG4SJUTLZeCUckEKvB29uwKkYgl7PWAqb7a2xa7Fes74Tbj/2ZGJJtbwNb2vvjDj/Pr1GnXYS19t
UTWAv8hPx81hWUVU+DrRpscD1bUWEToGHXNOH4Peqz7BmTaialB8KK7U3JufWCopCxKaaRV+JA+I
pO2jBntKSQ8BZQMSWRj28mpmRYyN+53KOZq2mXLNlijsXQuGBCDioGhA7Ny4Epv2lVrTPmSJUKhp
y2yIQxvwHvxV3VH40BbNHm6aj3HNB0GcB2HijPvBecP03urOzHz1B27W3/DIg4NhA/QGIvg80h1O
iy5mVZG9Vj6zVlmZvb4cJvxEkMOFFWmpJqZVa9uSffVyl7XylJxVkvhsAkE0oFBlBpTWP33cv9XW
AFTxFJ03Trwis/Xz3uLoWPprp+GqB/wGkC6zfoF43VgjswxklOf/2ExWBXZ2+XCGR4ujqkYaNTZF
GsmKT9L0oEMkGCqxlo9STLJGIxHIx5tkF3VYWHkqNFtgnmlXiGrw9TF9t/tI54mk04Gzp0yCXRe1
CX4GE7G5T1srW0i4l+wqwXO9E/NOxp9382imL8vQrqFqjB9v14OidvEBUMKpUCXUlNWfPrhLJP1+
RO36JTtqwGmGPCobk2eKi7U2xfxA8VOFN/ckhqT6vsTvpIaWFyoZvgJBvjj9iLi2RuP33R/CIE3g
jKJqgVkF0vFTL+R+0RcE/GsN8MUifZQcMTd5/g0D1qARtGfgycVg+0xmrVTimS3ADAARRoKUiJUT
TivET0i9wGILZfsxMocrjAWORAjGTkXU2ETx8t9J6F6pR3q8fpru8BFaIwH0hnQFTMnORhiEaS5V
Okh21XqLiSi58CIQbzbrrW1cm/zWn9JdK7Tv1loQsgquqy7TvGLklwdpRf8bjpIRLTwIyNg9Uuj9
4y0AiLY/ZPxaNNr1rptfqLnz6/FnfLpG3dcKpfceZQlQ/Yon1cZ/6LE3bL5nDfi65wNrFl3RZGUI
9cRpku47ikxplB3ffjC47zud38QNDL6z/7VdTphWk4dDxuGG4mZXnfzRDyRV9uozXUGE5XTlTiSN
MWZxOGZnSntnxz1jvS7p+EBksQ58EGLe3P5WhSdN3IAdgSpFQJeWmVZOCO4cT9MXo24v8cOV7IlM
PB00qSFvJFsY8ncYOO3KomcVjN17C7LPe9yN2Sk9iyi0Px0Q4Tlacd6qj300t3zDULgxyoPTceqr
IRNWA0Jn7mjINQ3H8yGgR19GO3mYFG5X4qh+o6d0ATT2V8we1X5QoAf9iHfUHbZH2ch2hMDMBUnI
Pyv5G4SLbbOd5MBeXUvW3wGWJT+5YdojsXmv7hxJomSvgQ5u49zSj7ckIPcoZoiFy2EsSwRqu3DH
aCYubFynX2aQSHgGGqLoYgsw4Fhm2rIL2bhfmsTowYAanhgm4pn4lYPUU54GpxTgqKv1obkRNx7J
7CO9wJdfk5UfGUZoUK5j3Oiy8O0XXPiyxbwpOlLBwQ+2rtoxLEhIY9btvoa2xwcLrIHQuI896HEu
w3383o4DJfjPc8IreALQ4lexywdhmRG2ISV4EWityGEkjMxUyjc9822LsA0hCQfn2MudD+O1YFIT
0ajsR0tFlM4AFzp20Fxe/wu4m43HaxDJo1r+bJOD5frMX1MvCm63Mqd40cbWL88j06R9jiEX0BDN
xo9oGX7DlaGyTTs/WXTScJ9rROYn4szSKRHv/SuRoWpgOrKVySGs0dTSA6KPYpCEm3H97kWBK/Gy
tbPzhnq2SHC8R6GO5Hq6qlDfbgVTK7zym2Qtl/WYaRiBv6TY7XbIyKty5ughf1ky8iSmez+wMpVL
jUeieSsBZB3U4itJkztntuAm1A8BCTL7C3WegO9g3A5cPV2I51wFsLHgkJ+eUcztfV5TLJDM38Cj
U6+NEGJ3Ff70IpOT1fvENx/eDHf1ciAK2W+B8OqsA6CXWPR8CXm8Iptd4NeEdOKfwgCF/lBB4qJ2
PSU7LyxUXkSydIm7oBtkiQ3O8u4xhMCH+x6eQRlBWiHXt9vK+XR3ion3vMwXcffGX90B+w+TC4h5
Q7HudWdk+HeqvCefgrkDNwFxYxgYi2t5M6u2ZSPQpUDm3teoodS5M3K+FAaNn6lGmXUmC2p/Dz7l
zfXJrEuxu+JnzWBk36R8ceWxCGCclfVCUJrL73kLN+fkPJwAZoxONN6+0ZPWQoMszeaA7Aq7HSHJ
wzynegt7L4J84Q/sr3w3yfq48+R1ptvZLdWpsWpD1gEg1WqmP8MiaWbSlvEPHGiMkI9haFsplnw4
p+Pl7QSbCksfEq8pgwc+HXsg5POYuuc1V314p5Ga1V8vfVLbpsBjXeQy3cpm3lsOaVifLK93TSUf
JE7i2/74Bf0Akefoa02i29BFTP8C0Dhah/xkP8nsHpAf3UBnFd1/zG1dNWEn/+sGJgEXU0itLFxW
xM1Yc9FU0kgUexK9gdcXZvOnxoYB6dTX69ulTSEJtxInr69W0kbhZae9IcdlVQV5t06WAPAlgrw6
AifByEIKwk3x+EJZnf/sTnO0fI36JUjI+XP/VCab0HaWlG2bD40m1pAdVbe2ZBV7heko6KUtxTAJ
AvJa7oJSa1zml5YYCOmKflYmAZn8p2166KU26l03GQoTeg7lkzzdq+I7MQv3Yq676pQKI/ak7Gf7
ZOzZvP3QemSTqkcqtLwWf5hOTq5lxjd+ixDkmsCmwuo3gG0gXcuMvzra1ECOf7HSS2WhO1BYeAEs
1vHliVdVmxUn7BlARE8wlHhXE3TIB+gwKyfdNKbnjGP7bh9CKlWr+PGZBl2y0pRr/lKRhVtPPvC7
DlMZNglP72D1xyoCHBLAu2XUC42Vr+fwuMVarSW432tLrSZwQtPQ6a7Z+kMaAVbB6exsJ8AkWZMs
m5k9cP07bPKG+ZvxwTlzOWce6xTIpo2KecReDQpapUGH0TN1N0QBLDRN4YAPTVMbIaCqueRbuKsa
Y0duoM4U2yhIdEsX32uSpuuDIKt4/UwjYyX3T5S7ZKMAvFZPwGZ9HB5mOeBCUOu+zMBw3IdiaR3r
uWf2GW6OzcxMu9cp05DqDMpPCW7h82xR4Jvx462ollex8uAf3PGHUu/auWWzSQsRFIb9KJYPfVRY
cN8Hs2vEJy7VX0xKRs/dm6ipl91+bjFcBzPAOGUUbjEq60Y2SmUeIRAnCN/Gr6SHUkriNJIKhj69
q7aJF0NfJF+xxOrSa3FjdkHKReoYQm/squW28xC0ZHY87xQ/4/A2xp2xZKr8ixDfmZePBmtQh6GG
Dd96JvfEnrqF9WxaFXtItn3lPyAZin2pzp3oqB3FXc0+02tUlSodAzAHKHROE6DntHwAUIBwVb2v
UkME6adBWdZURaY0DQMSUx7a5HyaGHge2sstyjWQUEK0+DQ3DutnbT9A9WM0S8b0OsO8P5H29lel
8LSDSrHoKjbID67191Ss2QT37+i3tMU2VPcn8c3f1LPzDkntu/+KDLE/O5L7qzsEq+q3NEGnwhYy
2bPk91chtV/RWEPm7cbDfgQWNsoNwFkz+0Bj3VV5UjnuMyXyeBrayrTEwbQCp+PbWsswdsQAVkxE
uSjvMFi5nwv3JfEfHEdm/gmHydJSUlDnBfqp5IQS8jHBBL1dpO5vUuIbItS4wj0g06nCNobcfIZL
T6EE/GofrLXls/UWaoLoMdOwHTposMJVIo0YXZVeX26pKLE6scgR0F3Wt7PqexQ3ZHl0t7tzMLYL
l99/uQCjnYYNCyU4pUj9e96td2ORpfgfQukxw312net5PI7I6p0RtJBNHMmOcxzhmzfZ00q46rVV
APEguW3O3QlWD2DqzRC8BHqLu11EFhu3YZORaDjomzT5ts8ZSONiSaQyuWa3MtjRYULFhT3rbcnN
Ion77XtOHdhLckR8wavYoPCQ5BbQGNVIoc3zh06nXos001F6oPmA12zkOYivsSIL8K2DR2dtRSf1
wlJhNi7V9+OhFIfeYmxeQnbYFwFjm+AtedCSmeXUQcPQQkg1hzYzYM2WZNqS930kueOFw8WeBg+v
PKpd6PQ9S0GCGG3reY+gqQAacegNKhHidEhoUl1IxdOck1KDVhn+FXqFZCuLfc8RtcyafuB8JFQX
wOeucj/qiJZ4iqaYsgLqmP14GoZT8XBm1A+aF365PRj+f0y5H0mbhU+RqFGLp+cEdEq+pbzxlwK7
TAWf7n/mZRUzcoFQ72snDXz+Wy41lEkR91a4kl6v74AIH3oyFN1IFfKqlueFztEaPhcaNjh5ebXo
2OxhJ+AsSgt7evRd2ytthdeZyGJmOBVN8cgkl0ikayCUMdWLKq96RXSLhSbEzk9B6kGSW03P4HVo
W3DB5eQ3DXRXYx+i+deXYWciBHxu4WhWf1DKYQMbwXfXXs+KDIJMXdPEwSTKafTJPp+h6HR0qzWA
hRd/CKiG//YH1Hx+A+g7P9gAWJkz/2SVMsSmzLFWv0bibfaw0zpyTdaVBJ+b7wqRf/b/8FFgYidE
rlHuBTvKQfWbtnRVdej1S4EtHTHfMDTEqNgwtS3tev+I74sfsyBcwSdlXncaGB2GRpfkM24QrPze
Ns3tM101z3I5ph+IS6hhHd5DGh1wgjQ6Bqq2ewab83mvSwd1JNd0VNEul4q1MTtDXU9dOIu/yjml
Q65F4EAcM6iTrONqppL6lWBcH4SJlKjwkQogojK1LhCUknp/zyP26Km/6F5j7s0K7NRUQ5PmsMNR
Ua+3OUgRHfhqp3HIUomKnTI7GXB4/0yL538gTNGwqW/EBr/w+FqTAoEjcOVV0vtwskHrKTiqLMmZ
Zj3zLzVLNmGjQwdoUcbv6WNJ9PCComWwjQppaO2sHAOmY1z7rwiY7o5I2631924RsE8UGWSEPodV
zlhspdL9zsT08U9lnqVjboKZHe5u3bm6M5do+VO00f/ykxhPskqb/mToz0NLzg9DIKf9ncrlM3se
j9nTHflimVpRJe4FOxyG4g8d+LGyjsoChfq27UuE1jOt4AWxm7zNZWdhYq845teo3pNuqbaibbES
vFIg1GIOiHwcPvFV0w87+avdDDooBp8LVMKRw/fo1O+qYLfkUSc9VYfBEL/w2HloJIYSIP/tOgTX
PDtv93p+CIkCu6DHVH6Yv3gGGPFZtRfRhXMaGT3h0XTcVlvx/OfRu2aaO9eB85y7Nd6IV6NPxH4d
iOAIreuPkZjeiZFyqlJOG4i3IVxEPMOzugUyqTf3H7HQlD+JCs1GhNld1LcHI2wPGPoMVgcKb+Fe
V42RE8zxz0zqeXo/ytH2MeNStegt3LaVuhLB4jpLjexC8ZR76YVocUTOO1CdEK154Zg+RtFZPyO6
oQWJXNJKzAfFd1Op6j+0mny/CjvdLC+UdkJRb8dvt4IUMRMZ0hTrhT8gscvUuhbsA2ou5UmJujf9
v+yQt51nrCxCFFHDlpEuyHeuC4VA0WbuZQHTxoFRfOJ87v9wrmwKhBhSIhYTCg7IwTcVV8Ym5rzg
sluCvPhihpnP4oWaAQLzXfp+YEht+m8nXdUfORBf19FdTqurPdHUx2mzQFr2gQANwk2GWhW0RK3M
FEIvHWFHLrbmBubBtvy2PaqjzTuAAxInr8KgreCrfFvJvrHyasAxZayelht2dJwSrdesOSyhLEUh
frhCdok9y9wVGxbdCMuoioF8FxTanA+nlFHGgrYFuhDwb5a6W1jLO/t7TLzeg6JnWZQGKo/FTKo0
MhqJDKd+WXZ/zhQNMHz/OIPZwQyvEs/DsxOdabeuD5PE5iE55Sbr2GTLGh/YYrMVFjsYfjeiqfIZ
5yMfln/xmCytVt6To5lnfCW0oaBpFTQlIHbx6WTLhTA1+Fwlz3uynP0BJLNrEbJiLll+HUlJclti
n976aURoRM5LZVtBvydqKZgNqj9wNVd2kzyLXZ2V0PV+Qe1vHuVa4Cw/8kwlMAMkZWnn//rrHmD+
+kd0qD7U+WwG6HtS+TsFq6AXjl+zuujTlcnufnltqtRWxHaMzMUzGEXaLdYqmrZmae7kN6fiPiq3
2rwK24iq/aqZp8bBVWgfJI87vjFmqJeRhowuKi2XQCQCGBHMIaStKYja4ZhYZ3AxCrCNDL33XoLm
vckx+a+DveA2iosThXPFpBDGnnfkeMuwauZ1PEk2octSzPaDh03z7kuw1DzkKueqHOFGPdApDjyH
bmyq8QOTbCORW+eZz04FFcavh+jcKolQGfJDkSNJYkFFB5vSkyGTa98t3e3FKYQvCAgV3V6oWI1P
16qlkU6dVNM3/c6C5MB5zj83Q6J+20AJDkcW5bJbV6R0jfQG+AZDkS3uOwQmqvdrKUxX1ZDRIp7+
IepQ+fmlMwD+kgl+pre/WeCQih9JBp8K04uGEjBKkeOWj179q4GWQYG3pnJOaqqfVkjl/vU4KhOM
/T+KXZlI+My3xlxwJaQSsAhCpEwRPqukG6uLmy2lqBuNt8S8YPC/UNvYNNibo1b1iMNX6nZKN/zd
kLU71aNgADMTi0Qnf53GVuLhaYQs1uu5L2bOEJkTnhH0I1HLii91bTTICLd9va61/C9vB3Gw2fLz
nPjrQnsU237/9nvfqZRxTNhDEtDjZbYBmIz2vGwTJ6uEjs+i4MLzJfzUgzsb5CeBXdUrSvU8woZQ
WLoi8gVy5tGTwEIT/rT/d9Ja9C53o5KtpqPAUBOsF9c25dHj5QcPvRdbJ+PIsYmZEmXwlSMhvRv7
wmrJFgQvBLS7by12e3u7gPRuYTwYIU/P7M2WNRIQ5IIqokRAw4EF0/MYz8a6+egxaJURZFajMjYR
/fyCEfLHNDqmdh9T30oHe8TLu9vnR9kjWEEVPvCBMH6hucAqUJuKtHxeV1sOGJrD0i5pF8e62wKm
laTgetLFL+yDOUBKhP1Bauy9tZ0bk7adM7yyYE1iDWfnXbVC3PbDeFwA4/wjUMQRTGyrRLY/AAM7
NfPAnpFo1Ng8ejWojPjKO3vLID5TNj2st+dKGVvw5rTn+oqkpLkhA3/JzlQZLyJFnKCg1ha9KEkX
ZNm0SOIlLUjJhcZ4PeeqyP89czwvbLTpVUZKSspgogpQ3Vml6GqbieWbkjKJ/B1Xw6KvRditfuLJ
LQVZjIzvYiFt5lgLpc35hyA9ETDO+C+ecUBUtktWDv30B5LFW2RRZmLT8gHE4F4ABQ2qOFlwREaK
dH6UweUiaFds4EL4pBU5WPLPBcEeK3KVvqhT081s9LQ5i9AXEt/vKUkThszpmsgOc1elEitI5LpE
KRb2l9RT8wSxzXc37bW5lPgcG3JbI0GemHGygSG4AjK5RilsI9+YLy27JbE1GIXfBENkLSl6x0uW
9tPiU+R5pT5gdlc6N644NUJsPzruxaMQSFHPe2HliRmnYNFexAStOzgDIJ4IOXmndJBISV9v988R
JRCDT/ngAwS72Ras5A7XNgDASaybAfruSyYwnnc1h1EgiSkJ2d9XGpjZribAUdAmiSOcg2rc5CvC
+AdOyHKxT5xEgTEAhFmwxWJ7M899SDf9BN3pbK+0LOsb+B6XbLD8gBmmIx80ol9ZkmdRQbPdLLtu
fkhj8b+VrkYyLk/hFSg2A4djGB4K5biRgmZcG4HIDIzJNNwhgpJoQbamKxJx3bNU4X/x1qaVAe5o
e9nc/v6zXLuDYIEik6sl4szjsP3U2uJn7y36C8qauzUzTVSagI1Rz34MJPFykOobRAHPYXN8Dn/a
gUHzPFzMsINvWxPsvsekt2hVJGjWi5wDGjlXQXFgIUwFcFQFaICBmTjtA055HJQ9BlWiymcMx+Wf
hbnEbTvaoOOIZ/dz95shopc9h9qLzKXS21MxNWVj11G+FoCeI1zFbHlrGxufy2bFxs1YXyTGGo5P
IpRxS9nYhTnHNmjzrP3MqXXDHz0SLTFdLncQP98GgbeqsFhR64X43laUjruxuu64AiVrvh2gqD/7
zoEk3cedc3eJob8jotCVH+Wh9wULzdx8Lc78aSouJ7VcZ+LdHSplKfR+Y8hgOhRBj7eqY4RgGufC
4MlWWLozOP5V4rVNuDqkWKiNgyEOFQEt1xolTI9ZJs9rpQVc8u2XyL0+IJKwFMCCNKrd7JhKZOFk
478GbGUnglclYCBKoNjUKDK1BRSvLh6jsLLU/cnNaiWLuCaylGl3Yd86x/LFDEi8iY8sgX7QlG6Q
LoiQQAYKPumjbN+Yj6f+qz68fORryCyPS23rFjnfP4dmCdncR5p1BWaPOhapb5T0ypLfViURcmb1
l3XalcLCjBTIxrY8Upj2RRLg9IPfPUto23rBiHp9ZyEIoFVXxxS4vnjCnZDbVTtaLA3h+oE0P+dc
BsDeG5iLawnSapnXsHDJvwC52MEzA/TRxJeN8zLZa466UWjpIBavL0nh8GQwXrIoUAe3Zs4eJTfX
qwD3gq9imh5AM626Z7bZ7PXTY1WlEJoESNvE00o/u62HWdjwYWmyxX7drC9oJHzOwmLvucfv+5t8
GLA/4W0b51Q5Ow9mM1HJA9aojBa8Qy26US//rbS2qfKwEPH2jV1dAtOZttpVdus8Vs4vzSNW0fcn
B8/o/n6Ptb9v8dWM5ZVK65iBz/6Io6FAphUxdv3eYaYfvw/ItUHpUp6ANBinO+hhRXzJ3QZr3+Ol
kLPAdqxCwzoXamonypsoI3BWXTX9saRvCcNtmElDnYSH8jzkM65e/AeFnwfnZzCuVt55sRhQ6Anp
K0ewMdB0me6j8J6N7FkPNsU+aPFkDiY/uf88tg6iaQOYnQYk6y0qDA9I0pg9PFi4rudTEx3i03wi
0/FPjoByVglCgI6tPWu7MgKxZodQT1WMspuVsI8TowuTBwPtBOwwJCEJaGWLE2Lao2XQ48r/mcvl
e+Mqq+Q7zwN5dE3ZtTxvNjnja6GlyjHv7F/gR2lQy8ep4gdsKu8mP2skuoLG1X6Vr57q7Mftp17W
OSVnle2u0yvY2XQDOv1klscJTqYbfyPnSa4ad06ysKDc1r/MFzlH2/VatrS42WwvzHwR5q8r34ek
CDfwgAiGLehCUhipH0RTbwyx7/KqfwNCtVZIOGeseJEmeP+3gQFOyjNiccBcKEGCDLcYoI9GeN5b
d6TKARqNCE4MVgeWysSR3HPTnxbdm8sCUwljeiAl4ZGpdaf6NuD35iEd3HPEatbZMNz4JYNdcKWc
whT2/YZ8pxmttIJ6ILAfGYalvesb62WDyD6tq6a9sK/6YquGywGdqcE7sNFPZ3PgwSKWaKJ7oMq0
i8hF62nl8vbo79NYq3dVaGCXV5lJCETdOUbQImBGtbOz41OXL+sT2/tg4fxa55s22CV+HHL+PhKp
1mssrdvvQ6u5zuOwFFRPWY5l8VDpRlTjvErnKlNlYN+sCuwKddCCAJjh5Z3PwlZpF4fEYi1APNuP
5rZWJFu/BqlYT/yVXcliNqBeBGse/TZYCEDFOhIaqrvtFKIzOxvSRYPoCCJ87j1rjJYWlPapWPtP
nUVN1KwbuJOux3oR1jTfejSRMRD7Detc0o8UCfWsDoZuLQeGSr9upibyyB6wTAZTjiJIzTHHodHf
S1fu0uwCmVTsl+KqYb/0cD3qqCewNR8/OnNUM+9AQX67rupSKqXXdBhTBFBz1ytxPMJLRWeryQJn
kC9lbpdNQ3o/MEBnNvzovbRStNpvxyaJWXdKQ2g6qQWCimx96EknYRGttGmMce2H2SW+pyOo3v8n
PZDaMPE7edfzd1BTK3UstF7kHb2rJOZrJc1SJ2j8+XdFGSfXavEE7mSJaeUYOmiBkFUe/e0KAWr5
AKtYvXgm6Vv3SzcHjPeuUP2m92A1gUTB8bt59t9yzoraY02JcnIuq/szRAmVD3mQcQgGAVU+v5wL
auxc61jIiSWL9pD8DB/ULcfSe3A3M7MVmOEvqEyRH7ydKHN5UYFCks0Wkh9eFclZqYXp0Yt7RyXD
4QvTMd1tjur3nKEOGyeW7Sm3URC3raYRwF9DUCOO4Yp3J4KeMBn/RFvo3GSmodThTPJT3r+pn2Ba
fhyf7qyK9ITZB7D6dz3ZZf/52+bMqapSOHdIiCQWVjv1Tl4/6O4CE0yk7a0nC+1r6D3kqlWfut8T
GpTFIAl+fR/YTKzb2QDSqYT4eoXIdSYpvIA0X/br60S0KZGmFGqnSnk9hgGBk2aOEkSOJu6gxvmG
ND3lBVXhzb6uJyGGiBHZdYIOc5+QSMjgWryaRGYZL5EYr2ZxbzLzDWa1S3Ebve58Vxdp29Zue+Nr
9nqxkJSQHUOnJWwJzBrFUUemK7O2juTU/qlPDTQZT1aWAXTQgiH4q11F24J4IVjkt8sWbgV7S0Ku
MrP9iPu81SrRubGoqc601JwXT8ba+srn7RSTh7K5zT0FRdlN0WaxLYWmhvMn1DXyTWAYRK5tkHCD
MLdl7sUwPjbluqOAMUVjJKTjKp8ey4wTihVyyjR0WtwTYIODj4lHJSOmd6zXQapTDJQFG2JdYGjo
0w7g4wtsY/+e4bGKPnRucFXb/kqYP9BvF9KTd4W5qkOgFH6sQDIvL3lCcRVWjent19VstGD9mQWL
X2TcU6JHN+rskDmachsW7IBjuxgkVVjMsgboUynQaVBiGuNAayAb1UrX8p5J/qhrsNB9uZwnqS9R
Lhn50jr59ShOpou1x9QzUiUGiuGuQSzAZpuOsca7q5ziTw2+ZpZQRMZjylHR5W4Xwv9gl+/IFxhT
1Y4FKpRZTErtApVzeNu5u9MF5KSeyKJ4EvVC8CiGROn/1BzYRtcoOI0gQMvFK3s9naBOYtSP//8n
KOlrYosaywmPinwdlrdl8qlXpacEKAVpWyjqWfkTMIbhd3+sE3mOm2nVYLO8U/cdebbBZ9d1MVJ0
d7WQeP3ONqwAfiUKjRKctQyYf63UaczGloiTkLi2xs3kbH2Hu4HusxiTb1AdRjJvFSKbuzoCFEZH
ZJHM9UqlL1YmAbGry4gdZ948sH0Hcy8kSEQI0uvdvHbSBgwR7Jf6MSRQDO8W96+nvyDBuPZnL8F4
11lwWkhlBCRpmO+BxsLLNkJ6HfxrGXZBxFLA0XBJfXXl9+4UhCHFPLJHqz5Pd2sL2dRVNTNy+h+6
+1VGu9m8UMwb4FDKaSOc54YXZe51MQpqCY4u6K4dARxdqH2OylRvKeMwlrRXA9sK/dilnqjQgiL9
RhN4whBkPn7988+EQL8oYB4cTai49gEV4R0aRRQuy311utTnVK41V8wrIC8MgrI1EOQVM7IT7oI7
Gwt4zaGFCgvbZHaf5axMXBFgbPEhRCkuV0Np7u5Bw0xQKTeggDyvTLtZ/65/LV/8/hpqbBzI4b4t
mDdnzjSXs1ARXge3QQmM/SiznI54M3N0J1ef94h2UycInTCk3h5tii9oP+LplILcORashYQ5o1ps
piwf5LKx9/x8YeBvWXIH3qBlCicboNv/ATZXcQ46pzhEgYjt6HSxgckeP4HleQTU0SZpUps9s1n2
qcLrkXFUm2Ln74zubr7368bNhd4RuLQiCC+Uz6fK85nscaEtl6F7IAYnA6F2j1olxhKfKaKzP3II
lEtO7FdlDoyJT+7bkf0fSd6ZVWsf2rJlMXdoSeym8S0GzcyW084H+f/McfUy5LYfxA7COhTw0wI3
u4xyXkXmf7RKhJO6dCpl986fuNJQBJR7EdNIrdFYTV2yCs2fu4DnuJhu9k0rAuzCJffFJ2K6nCXx
74UPixZYWPJdG+rcIM2YbrYo1XNPLArp/j6wVtphDwuZwgfzSNzMUO+nGvRU7EcAJqufE8ocF9bd
kusTGdU1Ixxyibz9M/fovZ8iahC7VnAxYgxG4jw3SOwTPfLe6v5JM4BYEXKcTPxKMcn5BSPn9L1a
+HpP8vIv0vrwPcbfize/LIr7RQ35Hr+h6jMSTx4qR4VrcbIl9FiZ59S6qFpIOVtaS6qRWuf5pdqS
Ug/ZkU5/wpMAfbqbW5Utdf2X0iJYKfbMZC0HZ3kl7Q//Z2a9872Im5rq3ts2En0LsN1UuaPb2Fam
YGGrIvATdQ4wVyM2j9kQwDDaB9ncn6Su6Idd8tGusnZLb2T/5Jx5ukT8D7rBy5STa2M2Ie3HTdy/
CcN8XZq2Us6+81cbYQ48SF8RHLBVMDfd3894jMuCf6lI+aj2+slrIC670fdLAUDzVRFVynr0iJGU
RudxMLh90HswOqaWz6G63SJ9AozsAKOCBH5VlKR8yyOie6fAdaiYaCrzECNZNakdqpwtGNnhMtH2
LQCEUdaw7ziwQ6jF/kcK3bi2tQjGNGg6J5fdj42chRqh3KLIQbo6PE1KOIqKX/FC8ew7Oobz1HjZ
oajbdM+A8Pk6ymOjuU7VCqKAwpQIOEz9vAlB9Vzivi1e0rgx5T0/W5Tk5MDhWm4Xs587bLqbVI3p
ydsFA2UP2loaQmgNkzxJzMayUeBDYKFBzjOD4M/tCbHpDTukv+tuI9gBVFWsHUdO/38eVbpuEQZL
NuZhNplZwH+hfFecxZZDnTtSxY6H8ggki6u8N845SCBiOerJcUmtbVhuDZHmw9b2sneK8uVXYeE5
qIefJ2I3qeZU1daAqEaG+jIzYpvw5SjcWS/FdKEI/yjXU7HmvnuJoKUDIl2STwnVo5iw6M3liBxi
jigVZAoQLo5TjalcuoMa//JqpyglmgY4KE2OBNBldLjlp5DcC1BMUf3bm8Lnt6Xzxx7Z5m2sy60t
63/5erfDEJYAIkcFGdrFozh8UNRMEerE/gpAKuR2KM/heE/WJ8U7M5vToiqYg1bHPQFAXrIBDjr5
D7dHm4MYhawEIL0m0RadcgavXIDDaBxCyS/xVDRC9XVvHgmrIJeNWMRJCWHijzVW1oLGecr78gNo
v/4j05SUQhumYOGp9oIGblYh3r41Ky1iqDdPCEfD8ZaOFE+YG7eGEDIFIMWBMH1NvGQSC74jWlM6
w2t6fw5kucr6B1kfEHqQB+BVEHm9rm8ce8B95O85XS92d8SSY9G/QSy/y0RmoYkNJOXxhZKLslRE
iGtTFUlY0uoRON1TtVASNqzmfB3oMIvrwMl4K1rrEMgj5Wmi+nBQveYpiLwbduK4hqI8zwsW7Jeh
o3zpwBeryVThPqgE0aV4WiWmryS+aZRGi/RtrV2oEBy3FO4hQXI/3MGKg04otHUPfjVDwUfVFdJp
8jmg5X34Hwjovf5W5Eba2bLv5q6+1Fjh6Diq1dyLiwmYYXfhu+HMNnZ9nOhKi4YbayF5/1uynwA/
2d0fBQV7+05uhlk3OTvtu8siXp7e1/dLUmbJy5LZkmVaTGgokn5ZxHNSY9El0MjFrhqMgAZImgZd
xPvaMVwpvUCmTIKrSSx/QiJ689/VkqrE0HalpogZglSaRRcrzFGlTNEmx44IUzAp5v2qyrLygb8v
lPNv4Xe14p74CcipjJy5rd+Qd2CYvM1W94qwDu44Zc04D5tRuxTsHNQ7OYjFyqMnAoxUSA2gzUZj
0jbyudRsca3jJz9M3F8r4YxEHwiAWEBYsXKy15DtJ41HdPjRzAdP5mjC+1HcJp0Hl3d6ADL1tjGx
nRGrVhFweUCUnj+PNg/VRWXineOEq/z/c3EWKwHtXiyw2CodLIg16on4UEy3F9UDggOqi8FdU3O7
DYiSh+alfXg3as9Sk30PJWZJr4ntDK9EDeZuABdWKtOF+YmuR3wcSZF+y0ixmZE02WAZG9s+zNEV
AL/FuZ+0mIWqsgw91x1gjj0I0xNHZoan9vMnHhQzBRfvlPusZWzp+I0xggVdYsPgKww7UUt93u8b
UKePBXEovHc6XaP/5VjmAy2wTM+shI0SXD/uxl/xk07XEYevNN3UdhYZrlIb3T+0LIq25Gef89oD
pOCq+XN+PhIQ51qxA1pYKi4uRroSUaEPSwDABUnstPPtJPiRiCwKx6ZOczAqwx02eob8ZHd3NThT
mXjM/m3HAGoESF4ZbOl/1fkyXqgcE6lFzsQrA/a3yTRQ17iSUVdCyPahsKFpWwThOn2xxBXEdBvS
g2t4XIKN6q0b0EqAEtSrJGLzUieP6zrv5Mm+oJvjJ5pE0MSUr8fa0rqxPv+UQ31l7TD/xNHd0Dm7
Iln3tt5qzX3G+L4USd3FurSqzRh+t7JAahLAsm95BFGgfi3+e7G5yU6hLHA0+teHoLrF28k2ULK8
3lI+zHWHC4OdcKEur5NcS12NhlGiLMemTYcwlm7GGeXTtPO4aDB4XEGyyG479FvtqD+riM4/omvP
ZxzDTLIWZoKWOqi3ryLfQtT5qJ9LVl9dVbIB/ZmjpviB+NkbmkO+BRx4snne9TCObWiYaP0RGepC
UjeaCa3K7SZgygQIKTHP0JS8GD6gP8c8XJqZBSjmP+u2lnYQ7b2OgpVzJ/2H45BnxQZJM6M7s77N
c4BtzJypCd1708VoZ3++zAFbWq37Oy6z0PnwZYWpmRK0wSK0yC+CsALoVDA0qzGKAupOrWYaUTWS
38QTPM9pHevBEKRv/4sXc11qrtANGPXw9eH6Yb+Pe4cfokzGxRfwuWkxH1xTtOFt2wQGcFCO8E8B
GiFwBMfv641Hw6UmhUawEOH1mpEgygcKk2bzzWrhiWUOPxikIWl2qofnr44PljFzofgZ4cDxYuzV
1SZ/Y98RiVKNph8Kk3vRnWOuKAdhsLHSMnyeUseVUunqaYuZhM94AmhI/JHSM7r9UNjIBmq6tsBv
ZXaYkpCNZIw0e0gglyTOy2PecRFqVXYf1CL5MIenb6EOTQaUTfyXxmzhLwNhNwP4meyYVClKg0b9
rpg21fd4MIMNhNeG6m05xva8t+wbZdL+GdiRC+T3mhIarX6dg8ZJ2U3Nt08pd5hAeNSLQxbHrVOz
5uiFsawJNCYjkIOY8pssQ7XVoWbfLZsWQplaUCaGC5zqWOshcfB8R3JUN7SU0GJFDPDLVYY9py8F
ChbFnxKEJ+6J5HpI9awbR+R80bSZqbmcwWoCbxPFAeiQYjdwhc1p7b1hKPvDxfjZQwmepd4PWS/r
OvOfW72PoBtXqc9ZC/3mDK4EGW7LK2E7wua65F6HL2W9Oc858IiztJipt1sTfHL2cp1bzj1RktJp
7Ru0keiUNU2lbEKDz9ZWJ7x/rEXELjHrMleteu3X6kNX1sL2by3Irb8JgJ4q/6jIwiilQzheLPbe
tyEOi556ZAF8iNDq0DEwM/uvlCcu6rs3isEwzlkViLY69Y4e0L3/awTpHiKuUOl65VBN/WumGKsP
aJ2s4oYM7eXsDcpn2lCyYqeVJEIi4wdlhCTxiHfL5CgWYvlbmhc4LQlRVBRCxZ9QzrhGzP0wI0f9
mPZElfAIh9jw00uik1Ocs5BCLY50OBsy2jak4gHHHROX0X/3C648Atf29BU6QUCsuA0e5m366z1Q
36OSDgcjVwWuKLDsPmesHRqy7lY4eQqtcY8T9U79feKEVji6IlelhPo2qnKqQPqqSsTPxXUnI1Xm
kSN3J/vjfw0a0f5xO21zxjd3Flev50R9Cjkt1H84Wp14zdUKO3IetZ4JAeNNQfBXXVxEKOk+ouH+
8kmip1Hwea5wh4DwUX0c4S5TO5O3f4fsocxRZgQcSLWezIbJYb7meHavhlFL1iSt+jklQDF0vI6N
xa7/QuUTm1FFQVJ1AfARVrNZXzUvHDIdeN+ZHfMkkZfxWMfKgsFMjdgTPgCfFPis6LWP1XBmW9uu
hWWtc8sTqe5UfHjTsBI9ahQwyeoyl15JvRzcq2iU7d5NPyrAMyNqjfokwc3m1ICTGM9cf81khfFb
xIyu1ckWAoZyOunN/PJU/2wkoFeLdRC5jyySRErw8zv8MCAbNnLApN1478xhNueW3uN6AxXjNYv5
zFpQzxnoagCtiW02VF/P/HhYlsvbhNtFKwNlToz2xUWj2XIy4RsKCbZHskBrprIteWF8jufHTHcc
pOpLAXfK33Ujtllxx6eABaFP75hlwZEzkZZTSXiISmNh6JsgZanm6Tgbhp+q11o1vKGe0oUuSvnF
13L8QSxFHfYAyh3doVdpE9SouSwhoS/n0nG5aB3BHMjiH9hiw4P8cctQjJJPYj1olcDjasTnpS6I
hs3JS0SUhU1WkuHudiEhJXtM/yh+JzXJLSLIR49phLOLco6SiPxiNq0tWalz9imoQWKAoNkoDymD
OXrwlKqL48MuZxiAyC0tCMQNnSpte9aV+4W6041cavG49zCxagEVl47p9VUaD5iphG1rtUtD4cxw
29mFUxrSvggn5Qtnky4KLtUeR5GcjyG4KnNgTRA2vEcLONK8ztGOshx1pnkC+CetaYaTZfm7uAUF
AbtilzfleXihLWkZDUNclo6e165w3tC9VIw5qcg4h/beZI67xXZtZ6u6UR43pGIPLZk6Epcw+nBD
7DK8jDIBvYnJPGmpvoECCHU9M+S3C0xEH6Sxhl/Rlz7xVr+k6nBXdiZcH+vzu32NB36IPOC1GEdk
ARwxo8HYpVkonaoK21QIEh+gmXuUZKXY4o+2vApJmQ5kAlGIR+HvJZ8qAB5rwaAuunxAedj2xr4c
zdAQQfV3a461AOP4nW36NBGyueoh7ylE5p2WiuUcrIXJRuiDlDJy5lb2MlDWR0MhAxwhXKts58yy
ZLsyMPjSTDBAPpV6IrZmbQS9DDAKgph8Vz4iu96r8/HvqOqmTsJCn1hWOQ4Ql9oR0mI4F+FfDKdx
BTnE7/0ReI7TxJGpLtOBkiW6Q8Z53lSQT2SMBb2kiO4Z/ZN3967QYeaR2B1N3DUf6GDsA9yZMohN
pY8EIUvRty/OV8hmVG3+8k8nifVAzs5IZJM7YCLs/l5+Z22t392ltVjL1Os4wU9+O+3qwKCnvreR
BE9qB49iou2rtaKgBAPPAD7KQ5mqrZz1dSsp7taxlm147LuTBr5P1AR4FGFEA3Du2fFS8ALKQysH
OyTi17aDOkxKaG9iXp4HxL4XpEL0kR7rVL3VD0svVgt16RfzU00Xbw7soazaDVsOEc4d90bjTbac
k98p40682qio64HP2/hIf6W0yuWxjR+Awotf+xrKXdjUcGg5CE6eI2vJzrE9UT+GrhPHJyvv5JZo
pKJ4QIei34Y/9+UtmikzyDY++u5tXGxpQkO2sw8eZKr20aFncOG9Yi1oVf19ZytjPgfUoC0KlGse
k/m17u7tHzOrxZ66aocAX2oh/fwB4i+FQlIdIxndwjFTies39b3b3F2iEHsXt+i/StwGNj0rujSK
zEC2ZMXIU8WNshAKC2FGKdx4heytNtNUOlR11hF4A8CoH5nyaDs+bQeLhnlOnmV8Q8bLrslaCsL0
f579aGDlE0slDuXrq3jsBzwhpuY7gmYEll9S5tII6QDWvguiXEV93+yJzxgFB1xkbNDzECvDbz0u
LAt0v1yPTeU6G8LkFT6Y4pyafcK8Zu76vuxDmH0iOPfkHXa334QfqQXWhn6FsW99bNze42Qp9SDv
I57XYd6SGa3e/9Qnn7JYN5SbZXHJ7qDO2wNmmuHjxPACrUBeEBzEFZl7c5mQ3aAwn80tX0kUL/xX
rQXbY9byLzQxns/Qozo14b7KHfF/DW5rHBMT7gjdm99IFapTIBgN/IdieCy0PdtLpKDP4a73pTXA
cTS8v63eYYVI8D2Z0B6aBdf2ne2TQHK2kgpwl2QN93SWivtxwaRLVDNHXMY/3TkIVdN1Io1tq52H
1QMy63C73aBZRkHD19PAXz9CUYXQQH+PDPmJ7PBXFLzA2fLFnSJeCok44N9VZJiW1HHwn4qQ6mAV
4dh3ETqcH8HLScjzYPHR/kp5XbLZQqFHa6sb+RABL90rwzyE2GFR8rdMNXFi8HGflG7LcoLX/ged
gyUHrD/WCJ/FGJVdLA88ggixFtvKekTAlQEAwr80dR2Cs2yOF+M8B62duzTz43j1L2MeHbpavvx1
kEZ8bAgXYzDhlbje4E+jBNj8xs0ETLo3R1ypBxoYiLL70/4ljBGjPcJCbkqY4TFx19UAN3BmDGFG
oBciTSQwe9g0zBld4WAlSpA1koxAhNpSSBhkKYmNbi2jdPhAGTsdp04HDlsaAPvA1ibZlSw4JInP
1HGAlJxkaQcHukT2IOgZWCphUq/kyIRdh3llkOuYq9aKxPY82W/hXg3Q4JRdfaSRW1B9OqFp2Uag
ALP9c9CPUtALXrMHEBH9CTDEQh7RywDFZ34KLCamuEUE0PuXb5eaKm7OnVz81hqbNJ2dxEIePnhr
SS2Wdi4y4dxFxfXiupre4GtmaCJx29fZzyoQwnPAZgpyBIytwuVOMn5peDf1t+HkoGIUL9EmqMmo
YVo5cHtknAE8NiyggX15Y0WYbRcKDjT1fxB4ut7oeIsGPYsahb2TlqQolnHt1BGnhrNGN9l4ydPY
SWQLfKKM/v6KC4svHXGXINXKUfe87X04/WClYi/AEs1uLtCBMe+5reN2RZBrq67gZcTfksK7OdAE
ux26R8gfEG2NK8MCmXr/wscaGSuqkvXzf7scnFmu207vcNuDOA41KpBHtaNh3Zljz7OlRY4Q//g4
FtoXG/n0Qrs0nCud9N75nAEstjbXhNKjlJxAVobKJeRRIqaJOoN82NhGzpiOf0Ajz2D1pe8LYf9p
uVezCJmlSsR/JJEoo7rilvxHLxIQQhWW98s+jmTX7PtZZMS/pNCZe7wIeTBsCIRx3RUnDNSULvqL
X8dUBKWbVUzyDLk0LXMqgkEnX/cajl3FN7Rps3X1cLDUXLl+pKhedQPz476RFPBmahu2Dy3Ztftq
PY0G4zdAx89FTpwIYPYGh9g6o9Qdn+3n4XcyARmgGjXHgHwpmwnyXh/LPzGFArHQ/OdHUY6kt31m
cYuqS41flgAC2pBXtzxm9zFQmGRyRaHqdoTw3HC/0CfdHaWGSzJPsi2q0Sfm9HztAfTA4rjIh7Y/
lcSzMsFIa95MG2378GAfG+pv2iSm1gFM3JPWb4BPFD/JkXkggmR15sNM0TqFcRuqTTr6krxWVZ5W
C5pTub5Jfi9p6mGB3YtRonnFXyge7ycyt5lxB0/A/zWZSJwtRhaGkwhwq/LV/80JplyqXjVAep7+
ukloJb2z6iAAmQWnn12VJlvF0x86BtlyusPSqHZAJxQqpl7iBawjK4RNqYh77rzqFmxZGsfueIhv
eU3IFLA/ZNmjxkBOu4QxQKiu/F5TNdpRau2656y3wIXW+WdTqFkn/ZeOBmtdWkl55+vFkLeMbAkr
avO4Asxmtkie9XaZSFGeqBYT8+Z0J2NcbyDvSAqR4bpNJBg/PYtEaWyJxEZt0EY3v8IuS0zBUfiw
9LN+H6UN+I7wTxj6lkd1Z/b49zR5f8Lg/bsTN36K+Su23bPg8Ab6UGXjosw/O6JOf0k4XttqbRnV
D32x8+0oqBbp2dOpeIoEev+lyBjv5yj3L/LMNhOkbm9ZU8prar2wrSPp+2GBbTI4n2F/uTopLY7C
u95HJhMVKmTPP0Jno90Y4DbT1WvCHsBTxVHxqF0ma0xvASNs0R2Ek8kg5U1Nia3E8sKaw3ZXrfRo
VNe5TbS94Q6zEgxmA3pGe6LyQKAnqaniBROEgHcJglw5gL5kRtrWnVg/GqjxzYyhy4pUNeiounyk
k8kQgXi/ZvJXuHm9p6G8ptPkYb7Yt9gP6hL2AW34CMjpe4xNJdbJC4cIZfD3BkczlVRfpIRDnaIi
LFXgty9s9HoZBrhrxvZtigvebar0b95snx6+/HF2nGCdYdoWDNfnJ5Bjkja6SgavpfGdYr/u0S2j
zdBP6z85S0m2XlVmz2ksS0zQ3xaNDu2v8slMYV1yDXlsPscXG6GXZjV93f2e2Cg+WlJEqJ6iq5mZ
V8PQ80VAewQPHGyLtgWUrq+J4wEbF1yoI5KZNzSOwdJlm7kNZB7nLfqQYvq5vhujiqjHA6ZJ+WIN
kzqaKGOiL5E9q4iK/DGIAL9S1S8CfIC0iZXBNGJowTCcgflOINwEWoVACb/JVl9Hhcrr7GqDBKOu
Ye6nHCvQvCd0VtVzNbDlovvXdW3hqMLMUKWh2TQjdHDQjk+TymbyUo3MpsxY1qIsNIFj+Fg8zE+H
W+MsNJTv2mEmIEObXdYCvMg3D0BN5Wpw+XpGaD+CnCygWIgy79evSr3pF58e9fr9pcKrkeY9aJh0
qradGjrj1Xk+jMqsIPw5xGrd153MCtYF9BOVU0ENrz6WNSRh1yHaiCqFbhWy0aSng0Swpa3wmtv2
we8ZWTObBOe8dqC+SokraaquYV0MCkkVXJQ8DzW3mUB0rMWIdghe1LWh7lq5j0oVFrFT8p29KkTs
RaR5W1cKvFui1lZ6zm7k0kb7CYy4MKvc5aS06izDz10Hx/zhcaS6u7cFDLZMawVuxOKJnG0DTvNn
Bk180H1CHCuht8sp+DxWBV5x0aXG79dajlHA4J44HvqVVIZcL6idXmhlV4XeOqn4FqhxcQeB7gWr
1I16lWwknwUBN1D3R8aZG8StYdVXxfXLO7F0Fczyk+fBQcFBwT8KxJYZH4iv8MGZaeQK1QNMpOPD
EMmrXg0i3Ir0INc2EYVLsQcptmvbFbbQidAd1YimTWucQLDvPLJkLkWnf1LTOAPz7910fhVhwC4O
fu9jq/0Wzh5jXIR0/I7JpQQVt4kc963lf1dIZU23bk8sxI+uNSxCL+ZEJ5bEmdIOrHGq1TpF2j50
cxSppFR1xcXUuQOhzfZG6QvmZ2fK47r2C50Q7iBP3a7cAyMOuLcK2Ofz+6T21jN0Ul1olisZW3IQ
N8cOOeIqI/Vq7Rar/i5Y6LEfBWd3/0p7jD+sTJ6yv9U0Q9pZAEAvKSvtVZzeJ+njDOtxXd+KwCIr
nuo6F89dtFhBii7quGqyfMsAcf8oEkxZq9FrbQTVvyJKkFxxopXQPVszcHjoZQAHLHJxnpowp+Nx
PN1xD+yUBvdwoYnKBembUQEAEhMtxr1bPXiST7fuUMWUJbqtR1u0SYnnb3WivNIYxPo3CmmxOCH/
SvoyVHUmbO/5KBWrb+eLlRCAXvAGQWyNKiwPQHBkYywWrBxvPC9BgxSJtq/i1BklCAEEl6fF2XTi
moQHSEaEZ8Svh7h8MCYIxjQNrRd70B5gqw0jrgSRavDJFeo2alq7Y4bEJsVI6Q6NUP4HZYNdxtVO
8bwH7eCsQjxS9nZWvhxTIjEck0t6mizfs55KWXpsZJe0Al6egvlUPVrI5GjOD4+59/ymFoWMOTSC
6WigxfeFXDUoidyOhqk8k8xdYzdOnW9NLGvcHoOoLsLvrNb2v6X4ERPDdH6sCvhA+8RAwQK2pXDk
auxO+Fh/WkJBIatFUJ+mCzGUwsCYVrvN+aFQwCNqKM++YpB6DfCeffnWPh0oU+Tsg3WB9WHn+rNl
aG7onG+htC199Q8e/SL27/MeKEQBHx/nxs9/0c1LVLdbQx2M6fkfN0peTnuvVywji/dY+YtVIjh5
iDYoDAkHcONBv3V94vfI8szjNnsnQiin+UPwGDFLuRsZrKxIUSEwA4tYDhhlwrVvcKANSvA5fFjt
FsrO66SH6xQf9K521oNBOlBAGVUDz0uZJQ/RH0k/vrPRZwLvQS1X7G5Pnz80jkgQ+JajY4Mf4Qsx
SMsAXmhsgsVxycd7FNKNvHJAS8xSpzKEAZPJONbGyA+21xElPbWoQ9trkaKd2vK2MKafUFw8FCeS
vi9FYiLbxYu+4Y8Diwc5g81LhiylTaV87tphoZj5iqf1KeP7dgMpGSOFP7LhczNNuIDgZYgNPqbV
cBjXcfjq+F6JsiWAH9wXliHqoXt/xki1X6rFLh23v8AE5Tv860nxHRWdGQ2WHR8MIQAiYlVPnF8G
K85IAqX7MaQSBHDgcKy9U/yM6MC7vEr7rGHtm1Om3uP3NO747V1KNxJSLIf9jiGCV5FNkG9vzuCa
brAVP8IG6xU09azbGqLseAijpp3UtdnBp5GtXyb2AY5dEa/lq8+/UB7ZExdxPv9V7D1K1mDEumOt
qqmhI6jxHFbQlHi9zkFOdYGS5W83NyWlcZEeMX08od+n4j1A3wqmjXMRBbzekcxf+8IhMKKpX3Oq
pqlzDPGCsNWzufkW5OuvGVJDmCGj4PyDq5zEeIq/rJvPGb3eOlviO55smKYxTpcKOpUA8mohY2vw
v2DVYqAf9415aSGwEm9qlescyo38REpvS8RBpW7VRVQkkKs1I22reXs5ux3B1kTuYXdMaPphWyee
SzM85Mgir00PkgD1nEueFT8P20fATZ6bG/RIzFps5nhFdgaG80yNgT5Cuz0hcN11E9qLdkf6m9rm
jQCsc6hHTZZe1oBmpXgTtdGe6Bd+8S/zOxu5FWcdCww+ck+cpy2iEQLTyhB39jBOiyhYPE3a2mJN
QQ3E9xgYc1RHS+dglJhNAxCDfvd7dG75UekK/orHaayKXu5eK+WlaJnYzZySKFfvmDCr0pKgkPG7
9Dkhcc2C//y+dnGfv++Hct+QV2bErZdvRfaZ6SBLruRrF9aWXqm/5jShzNi5UQAF6h/VZAyzZ9SK
Xqe6NlpGO4NKWZnfrm55LXEQDk4EH+vuKKxzPTa4G56/M2FZ+ayHooBW5zCty5VvJC9qENB5iBOv
kaOtq7YnZ9WQqUmEsb5pRsPtBerYDzhi/R1qGOsvMNSn+z+DbJdL6hgxId6i4Q8T55xyfbfADBGm
W7BsxtHWWCVGAGNm/D7aSVkdBu3tpgsGByjLXRteLBfxCjMFrAzDGAahXfUqixY2o0MUK4uuMfF7
haJbyZ/BElyTpBotSe3CF6/dvqbMaheOUavQZraut+mKKg3nyxxq1GvXChN0cvAFqt8HymHx40cn
B0cEi4JEa0w+sHqYI2mhqL2OMDMEjK0U5IcoVpHvqOQ3Lu2W00NFedKVt7DDwtQl8y7J5HqAQZCs
zDQU0Pn5lrGHJvjk4D9FC4ngw6GqcZOHG1gdyhxZN2CrN0n3GsU+6H/G3M+SOcPHUQyQdVqVAPDa
7YckrAiQAVkNI1ygdwItivWHRl0mbnqnkw3kitdHIVRjyROoImxqC5UTOj9BlhXsA2CYJSTBneQb
835bYm+Q6GIxfd6POJI6y7HBlulEqNl9BGIDoKj+KFpzuvNaZ3ep+RSjNiG6Pngewy/0APkSYhkd
HYgmyxq/vbV7lgd9u3XYt6Ks302pbnvk3tuwrziF5kiB5WXu/nd8hxtn1iLBMlOK3ONjTm2GFd6U
7SxKfVehPnuMlAJW1urxInAynm5Y0WYu3FzwwWhE2XJvyUWyuAhPDg/ycaxoiPanL+vmgYg9U0Dg
vH4XJTaX44GrBxOlzTkwLxQyMGwgBkEoVrtmYD0qVkUeJoq3APtCEWCc99fkH+5+SALzM+pmxZXl
oeEQQz1Rt1M+THkISLRk0MMmhEYDn+I2b6e5GpI3rVBBfWqcXoiIWKXCi69MHGhijyUHDvXf52tN
ouO9p5CESRkF9205I3XGU7fny2S43tN2WETMwF5QxPOKjsVj2p3rXEW9wqnnoiLePvQfDmbiUfRW
xziQXYtj5GEBGdmTvaKvPxq+M5sFP3vSdp4wcF5DCgnxyctThWMBVtRHX/Gg4AEAtoQgXDViaCoK
Ht0Jbsi8awuH1pyBpAyBTfTO2C69VUT1lxodRmn/f80In7CMy30swjU00xyBnbpJnhLnyhrRTQnD
Q6kkjty1jDx3ja4qGQrELZP9yRXLKBD7l7QBg5Jwl+fbLjB6LQB4QH18Jxdukehl737pf+RloJ2c
4mFcewNgFTiRmEKiW6KGxzk/ZfdbEHpUCtDokMziE1eJZWlyFSN5tAUmv//dGYWiaKg8g8PFF2St
RCoL+89p1QxkcllrTqBza4CjBxJdKfuihbUFLpB9SjpzHnKwmEwzgPnegZHvaQ4bXN26CqhrOysw
ZqH8tlfSTg5TvfNCKsedtB8hTN5Z5SChNFWZEcxX4zSVW3fw5CH81bgKCSePiyN98zbZj+E9fW8A
APortILRrsZ1zlLfmsAgYy87Gij7J9xgc8tioF3AfHmVwvG7Y1R8EwUHYjv9AMAm84QPKmsnMp9O
ygncF5fW+sPdKLlamW6PZGrGEmgK1Ex5NsHgQ/cn1tBbwz6fMxbzu8WaRuFrx9bmAvt+rCfTGfoS
GmGJ4wlatAaAGuudi+HSdd0UC+lpMENklPX21qdTz1yT90a7M83kwLg+mpk6e11pOoxtPfvA8+AY
TOFcXwEsrNRN2cxQ7MIzwPY8aw+63ZQ9cFkqWZJwZWDzZsTlNMU9GuIE2D2NMRxUOQvGtGpBAv6Y
T+fEC5Bqt8hHnNVpnQKSL1rPkE+/f9vqNrdl88jigqYqSzllP0dAf5E0DZux2IuEAseYI/dBYppQ
jwnbIhzeDCSYzXgGvG/ZmSkbM6C62vAL4K6tXGq/b81p1rlhQmRPbVlL8UDkiLihfdOkfiLsuxHw
kXZiL8komwkPoh/ahRVmb86S1C8jp9aBUxrwKYqhKe3/G+dtuV/zBHuhcpsgQPAhWIx4QoHpPx9I
SVf5tbnvmt5K+K0wUiI+5I3TzS/uk6grY1z5/U1kjLVkfJLt+jjGDYjWmTva+FhmOxoIkmy3h0ps
Z1YYKuF9L6uhJFK8slaZJPOi12Mf+3jzVkTAqCUxOWgZEMr784TYgEIVJ79IdeP7PUMI5lYi8QfO
QPRmi9MdgR+6Y05stuDcvUV9qymys7ceI1FHPeaCWQNbxw4/SscGwGWcBv5rCv0PPe3wIpipj9GA
5t1KAiR4aBjPxyk7pMb/f7bRZqaW2ORTGYjOVInbHPue36jvJSlKqwNJkshXpziP20jKAH+HTgZk
9KCoy3OGUGqpL7K2R38UTNYwslhzlBJ3bn/BMa/7+9b2dnxMzb1feP4ZFlrMAF/1AWrDKUKPg4Al
fPSvmmi5rL6S/puaOoFlQGSfS2PAeTq6DPhu1JHSPrAABNAmIyRLsvLdsqIAcn2xIQtecfgZsx2r
sYDpL+Xvl/7paNy07qbVkYjrRMLyt0zwZvPliNnUFSvI+pl84szu9ZILMWR9OFKyQYtK/wCn9RXg
B1Tu0mYSeVMo2igtVEoQxVj6tNzKX9XZNxzZkxnBtXJZoxe5Sa+Aw0Ybzfq3iwajNWyDI7l3ZZs2
MA1vOUb2AEjoIIW3DRvO2PCUE2hSgn8RzvJKKmercVsGKKU4ruMmddpWsQL0txA88Fiy5p9M1cny
xq28W/UKlHC87BEfQETVwIBk1/pucRxqRn9glxlgX23G5H8jNmEzc3xp9JJURu08TScXcTGp773l
WaJrAZFnnC1GLrmsGP1srsMgCvyydxXK29dIHFTZg84pE8M9sJX0gwefw4wheDs7sCY1P9mT6vtw
pKcFMrePK5t6VCSsw+krERCTXePnzBZD2bP8Z1sU10jf4RXDWrZcuAVxaywaVXtt6T//HSakjt27
Oa3q/RZwaQyBT/cDxhtPjrt6HGjvs5oyRpXOyxodIWnqzHHETO0MUKG9AqbIG2SPjSN8Apws7Bjg
r1E/+1DPTIIEci6RN0qWOg/z+e6ewr2IATMbTnq8S96PYqsWQ9VIttlkukHpyJyTpx7F3Nf/wBxG
X8etV5Iv8vbYXkOZrGioR7L2pUt6MNX94S5fJqyY31iRCjl1r5leE46W0/E/UddSJ6NWbza5xC//
lr/xrky39NJ4PMTUeL2/tuKjfCZ39q76p/aIhHXHYn31dVlhGt0JggKK7XtzIe3VNBd1rmzs0Ngh
15H6z/K36PZi13oZPm5bznONThpOz4EEAU8jKNtmshVN4x74DgX53Y6t2BS8oEVYSzUay9YqLny3
jJqNzXD8P+euqQLj3LLvYiT/pyfhUWdevWLcCJVB5YfQ/dYeIIGAERsBlAiwvvKm+Z0O5tSUHr+q
0vFPUYep+Zuk0ijb4+oU4P9NweLYdn7yMOqYTKTtELv44+EruakWyhvsWiXvOpxRvnqqzJkLTHvT
OI2/iIljtUw27Xxl/u21QrJNkV3xzVKk8GDuw0PAvAMruGipPpsDfR+nWII4EAOunPZAJnyy8MyS
G5AlgAAsorxm/yPwz5ExsCqUBgVRIu4jKDYLpr9IRa8HYG0elzQIaTiBCavxLo2VMbKOkFmc1vSe
WaXLmT2Rhb3MsOKnuPSuhXPLDAouz6lkFhnLWu9swKXtqFCfj4Ou6OZMlAc7SPdPPd5os/+ezlH+
PW5Ar8dxANo6M+4N4S7afFJJvzGn4k+H/YpZP70jB9D9EVv3GKscfXxbLLFsu0vKbo2ATml9wh7X
vcA5I9DKhr2ft6dymHhkDsL8IWriFffGRp+yHBFXbByLV9tpVytqblIKHb886TMFkpgke/6h93HH
Jh7dwfEubXnzVC4T+RwggJy/KwFdtrB3iQh6cJMjY3ZlsumDXIfx/GEge/iA6fTKCO5BVFtpn+4v
PEZSCp5Q753yHdEkTdFeqt+hYGEsoHBCe+aBPn0TJ6G0Wjf3/mkH3YNrSglczaA1xHpqif+t/3lw
N+p9hUtqfyOwCTLZfw3E+dHg2sRt+W9xL1010yWptvCrER87qbpv8pIKi+aGsMGbvQHQr4hJBRTm
UqTzqo4AcniaJFHQaynFpP/kMW6sWGPLKXXO/8Ink1eF48zPTceG/Qm2EaOqZuki2AGJYxJqMGgS
Sk4Gq2frra4Ly2pNIpuRyqbs1Mt8x7jxgz/BnD21O3vr6DS5nZ3XAXv2Mr6UaMH1zYlcmIIPEi88
0rUUmcK8r2Oi+w0StxcfAYFoIM70wWB1ljuJZq6eXMPCFBtrdodzdVVcG0ZwEUKm6By4lePz9PgB
fGdXbpvg+reqZ82JRlzkXqvsF/JW5WE0gEvVEGLqF9kdFVgzU5dgxGL+Fs1cX9yyTzcTzvXgR+kV
A5cOhvRQmnCnas54tp36GIp4rbtZTXQ/P+AqVnEMjzrCsasCGg/0vZLz5VwwQJRQpH1eUjBba7wX
Qj6EppItk7MTseb+0j7zUGkEjpgD8+iMOa7igFzphLcMKu9CceJ17pqlPQa8m8o4jjJ4dzGQ1tO4
smCutWcEFE8RbVRZQHPlV4VXG1FgddRSkq2AVqAnZd/OptXWP7awRmewiL8B8YIY72RfO1s6d+Du
7L8Fg5lix+QoE10dVjc5dqI25ZUoc1sgqnNuxEFx53ylD9phGah7ie0DLnM6QJ62G3Le01U+VrOQ
MVyE9xG/Ui18UtQaLa+QWP4FZc1UNR8w4Tx95ueYAMbaJCRanbDS4FKoCsOGy5qr0Wj5n6E3kgy2
4gOHVARB7Xg4EGl+UKwVc/eixKnf3Hmgu+IsZZ9TTTyWHO1CHUlpf6aG/Go4q3QDzaDtoLxyNUih
gIlQrxr9e5aQB/zgIUgvLK+Nss6Pu7jUjWqAq5sWtud+98iMiqFNKuRvkKIof+QqeH3IR1BKzhna
HK829TEUwHnr96kZQRuSQLp5nnV6sYc/e7vnFGp769twSz91W0Vbesi5MkdeQnPiBG1PMuT2N8Vv
mwpj3NgtM87RLZdWjADwMUYgnts/4YElnm9YjJ26ayLXpatSSerxzROwcS/OXL66HllU4NXsmSba
4uLGdY/gHRAhJqXO5uvxpFBFXOZpApyx2CjIvpd6Y74WdhZIxI5jeHwmcbnM1v4b+5ov5CnPnFnY
JADD3duvIxaVih5LkKXTVp5H/feQ5SBgail3W508UT2qrKFJr3xp2N5x9XoRoGvUYFEU7nflIkxI
YbO8MRe43zJ43rI4l6T0TadN3R6+6O6jzMKGcFOqdVnTiVvPt6ZHn3SaM/QjH5vK75mgHcwY2+qE
tolT0TRTq23MD22ScRIsaDIsOQPDIzt8+NHDCD4L2LbsSHk8DoXVXWxjcEx+q3tCthDzD++ZwhT3
vmJcx0UXLsYb70KYRSY3d/R5w+Zdy4AHEVlXZN7FGQkhPyAyPV0eIcQyOjZhRAKVEsuhpinTh70N
tcD6E9C5QWnJJ3a7HdY5WQ4VY5VZXROf4C8V6HmO2/YQV/8lDx9AZeO7nrF/zNtq7Vm2Kw+B6NKF
xCLUpp2zvy4XYUUFahfOU2MBKTu5coAc8obxN2DAQttzGD1RCeH5GlguyTx1+u+/wuEYnmV2N6JC
FR5VncJYc3TUpxhf7Pd3XslLTrpjYrMsEdHezkdFaR40pnd018w/VjR/ksh76T31EQQZ4DB3rqFx
NIPGwFshS4cNH3fmUIt0ZS2aYXwmVrIDMUPze1EkeskOOhq0AzbD3tj78b9n5BbbRnnCTFghMX6G
gOIgMIuVKxX+DggERhsGG3Y0IO5hbwzGqU9wd5y75lBSbiyp4bxKg1HuHx/08UcXdPRiTL3xw1ms
3IzeDVXLFcuiIUgVHkpQJxw4ZCeH+Pk/IdG3AQEDmvByf3Wk0uIXQQDEUMM6BAJuydmjygosWI8a
Pt2kw3JyISrCCU5oA9pgXKn5OFxSSl34dY/7LTwiwY3TPRH69oj4PPXRqrDTLFxpCNuAOrlw5CR/
xDzKW1eFEUzvJP3xXAt50VfV/iytY42XERgBZQbe8+0BsGcK3y6CfRMCmHhvRNo5HFDmCIl5/7Ae
cTaLwFzWf351uWLYM2kTTKcru8HGVn1rqiIALlU+JGyoh+W/VR4yXDn2uvh3LIXhQrNNXQwyKXRR
/K1jNWa9xlmrYga31oChgy7SunArvqUENNN9WqsQS3c315B6ovgM8al1/VQrz77v31zyxpXStRgU
vmDpVpUeBAu/6tldwSvHAlkfn/bncnJLXRYbGP8hQACyB4fY4wwnfFKPbkU9CAZCHAtZ27kcHch9
hY7+4xIOLZa+IpajuZ54XjBZ9zi2YYs+Bz65UwNMnyk9YQtjVfMrFfmw5cHGz5tKb0wpAvd06Yk4
iU/6Fad+nWYYFceXXZKMxmwfrtEYDwqtcNEBmVsD5LJHQx9/Cs1MPg0NU82/+NK+BC6UNCkmTHWA
kZM9RM6a0uk78qlwnj909M6DUwMFjKo9AOUu/piWYy78PH+OBEi3klnDxI3l6+3SVHa37+AaHrU1
VNs9nW7p8doLO8TftMmDyEpFylQRLYQeFQIHaaJMC2J35hq3H75aKkk8MUyiIjnO9PNZaOY/3Agb
6fMqeHRHQamCJUGgh8LXAEV8oBLxsbeYPPZ2up75RWheoTAEUoQ+CxFjRNw4OY46au+AgIbug+VL
b7UhX6ojoRNmGxVllFW2+HUJY40cUNey5MPNQIhT/QbfLPkwQJfgJqe0kmHKhIURLDnmeGykysPE
7ch+rrRe5z8ocIUyeEeEcTf7XM6wCxHXb32kwseHnkrOgR8gwMMlVpxQ3kyuUqOsmTFpN5Tu1ENl
V3VBY+NWslRxknpA4TnfDGwNQBExQMSb3OKPNh/Utg/mKL9he9SEwKbfFYD04UuIdZUTx9tMn5Mf
TTFQX0luKb4r+7bTPVYKYpwQOzKgSMSG9fiTHAh35X3iDaQDZdwJkfPpcpR/Mx6ugV4SfTgD+49J
orvEW5299oGJF/UMEA1k8CrB0jWtQlekXCaaACi1S7HxBfJs9ED8ljD9oyGZ8xtFlQdtQXSbVBXG
54cURcrKL0IMr0VacPl9sLRCcrzWVXPYZYc2uUBdwwVetTHUVZZLtMFVb4U5wbGufMSWNEU8fubX
fW9ZV1HRyM7aiMKoXYCa+bijlLhhKg0Xnl4jE05CWRgZcq26v1JsFG/yqrFWDbBZs2r97WBGBUfs
XjnSKxqFNhEfjhQRMLr2Q0VHtYX/Bl3d/b5ulIcY8tarOQbDTALAefDyXPwmJg2rX3UxfXkXFzXN
jnSv8X5SsD8Mr9RfUYiPdV66Juqcj90f6QBubA9Il50n6m+iHkTz9l4rNes1GQ/2NtTGXoMvcwR0
QZ4FARW3HF9PepxwlSvbUHUe4tkPERPimXMnjy1UMOI82o2a4dnzxJN2dmdxw8ehCQjBZwszq9XF
upblDQNFiH2rLKZic61OckElAdFSA9+UfMw5++ac9qX5KePE7Ow8gl8va+4WMwS+YhhFHXql1BoE
24BMJday3NtLRwC3f72mVty64y8bEp4pEYtHWzKcPVsY+7pwhL9SRiwmesToTtky8WrWBpOtkxjZ
wCHYCFcwRWnN4M4/qw/RnqixUL2nZJs0cu+nYMpboUQbr1W5MYumKnzIQjfSFstxTsgWUw2XgOXE
IXPVJk7MJMi7NV/Nd7sftnHJtBNYiqQl6WbNPR+ociXi93PNv2oPRgiNQ1TsI5xuuvTca3U2g1tC
rHNWkXIMtHuv9Y//txN92pks0wmfckiMK7GNy319sEAGfbcGrzkTGCHbE7Bu3Epfwg+K00exKQ5R
AtgkToNPPOIoaJay606lkjmJyvTYeppH9+mVpyDjMpSCRYJKyt9YfP+kgobBKRUzFV12YcTHw29b
7h0em3NbjAh6DVR9n1VY29oTj0g0k5XzA/ziGf7HM+uGoDX99oGg04543+ACuP0jo6JHA8IMslKV
9kPk/1/3mIzQx2k0nHc+NgIi4Oj5nNz2P+jfJw8Gen7a7yr+OWvEai+Yy/0L0t+wCU+xM+GcSGgP
rMC2GhJl9eKEwiYOZG2HPYv1ZiFJAiPriELKR5AJ2HFObGYR0B0WtsuDPCpxQaYaCcyAiiDR7sc2
UR6US1vd+hQ0J0joVCGwBlSMdGpjJLtj8Gte/sah1G6/r/FezPPFyHtxQUNasHnGBsuOydNZbQ6r
KT1XidsCn/JE11FK4cIUNu8B+qzVYyfo/y0UgwJRRvdT0SiXEbKsky+0INgKrVJjv3PFuAabadn5
L4KDBHBO6pYpT8cMZV+txrMLgidkNvki8S80kasERPqQa8VmSe3GnHG8Lg88qIGXY5Ctt/BDYxDa
J+0TC6+/t96szDtUnHSp7vDIYz4o6FKF2bP759zuyuBqt+NMxfXAqYZBb2SBheeSk14IT8Q5Sfga
sBtaZxIYF6MDUrxa6NXFnMb6CYa0+glmhTIvlAsumPkhxOTdkCJ6pLFNHKE93OZQlnIJl3M7TBtm
+3pFSJaSGDU5+P3nu5c0edETJNbgLwGXaPa41vfwTolxEf7KNFhBvdwQxSfVCq2HFLGh+oKZepT8
fC8iM0tCG/937b8AR5NUlVFtI3uaHIIA8B7S36+MNABduTSmJKWua/5tq36+NZt03iBLxyp/zaB+
/M3lUmhI53VFdJHFgZ+VFRGWxuDjOkew/1jijddp3KYRKa2UKLqfMwlLqfGAVHbSNLVkEQwuv4sl
nLo9TxPp9ybG8Mu6EnfPYsCK/vLrrKoi7EOAfd9+H5m0h4WmGTMXiOcTDyPm28OLNcE15uDVVS+q
7TL9NvVB7KTaoYKRiZVcULGWrRheNqgQAQRCDLCRq+maB6JTkNnR3ioUZGDCKiKLCbyCuqZ6Yj7E
4bHtHWoOY4cVda7n1PFgRnTuHHR1KMSlMFUxPuc1wOpP/7Apr/7yTulbUQo5B+XZhIyuwINlMIMV
rNgdSMfl0YTlTN/LysVUtscIuPpJfCcIvNpFmCJAH9ruhUd9FT7aoFQOwDJw8ulGUhtjZUs9zdTu
iZxUWfPK9ikb/laxohnlc9xOY5Jc2sEgWTunD8kLqBO0KFS9bZK9GaWbtgzBEhAHS6tWXVDvzdOO
uYg7Jsz8JCNlQ3+WlVjJKZw2E5u1/zDjiAkjHgArxVj2abJ/uNXlu6Ied/ks6ogM+cmXnxHZDAbO
5JxUIloleLwmr9bnMG08jSsQ/5YaEClwgvylZ0ayRc2eytBifz8yqFnMcvJanrCX0XKpZHNIhEbP
HAdkP/X+ZUkfNDy2/S1/DvHRsEQcZV+jddmjXzO4Y6Y80hXHdqNsSQ5edrgeqDO+lzdyh4qlQW7k
5scX5V+Bg+LLEARHcOwMGdEhbqUH+FgXBCoS9tk/oqETBDV3JF/eujI4CeSzGQOiiYRrAWDlftJr
RZ9/1cZrAZ8jwrBmeFohi6QaJk0KijTWCn9qovxczp7ipV7i1CKB523hr7SvyEiGhLU9LcUK9+uQ
ESFVU6SaSYdJyOmceWfMbTh8t/4PKohbADab+VE1NCbrKADmT2KSp6VTBbnA/ZdPOZ7F2aPQFlrU
nNiK7YqfBc0UNhUxqtYDfeET+G2xFaKLaradjquRFxWQ0WACLqSkl/oFmWrQn/0UfqnleQccVqx0
YkW4dC95P33Z9rfCoQyDuqcAgcWjpsrvr8Bt/Om9YvYUZgVw0caJd21f6kAEJIICjbZepcSeCzFN
9zk9NpkVrOvGg4iozjgnBZEgCtKYLQa6H4IyFhnAerqAnViiA1wdH6rnmZsTgoe2I0nlTX1MD/aR
e+uNy52WGVHPKmA9KyQRDsLNVjMpxxicTYQ3j7PevdRX/YjhkFh3DuZNeFYX5W3WmYRS1uasAmJN
ZF3yXoLrytNwa2+IhR95sbYeUicmYgaHp9R8s1fENX86DhNRc/OeBstkJ9egfdBv3SHa0pNlXFUZ
2eBuGyaGwwddh3AOacdABH0FQEdijl4kp2IsX9+DJYEJnqAaeRaUHMfROz9LpGeJoyTPKtZUQi2r
5x3UOLDivUzsLLSyNxh8XONMcdv1cxT37GoxwdBMlFg6b5yEu4gssTLR1gAZ0ijJLtsp8ZoYKXJB
3Esm9bpRmw+Uf7/+4IIWijlfyorO/d8/+1BOGALDUhWC3IdOcYtMIqWzybxkbjpRVZkgFgfHi74D
I+JH1n+Vm4Gw9xxCp/s+i35pwATItC+kLdAgY6fuhSkJxgk9rb1ZPv9qAgC5jVmYn2Ms9jwETwP5
Hvvipfr/Nalpl6xOj1ur7+/h/jJczpW4AE7tejdYzCP2BeBD+Or11I9zwM9t7l7xdkldkLLIBt8s
Qtx2D1CKr5nSBxH6P/O5TlEf4mdf4LCn0553oPAFVdfXEp+E9lTHDi+GnclN0ySWQS6Qy4+XsaJl
QcP57h1ukUzIEex7PoeAdzmhMyqTHLRa11KPiN9Azw4k6r0q6xV3lU2CdXBauv8MF83SIMCCMULP
f/DqXG4YP0hYY4ku9RmTCyZk167kQeg25UPdlH3r709i5pIrw79HtHU2xlwUoZg2PT23Y4uPg8Z4
BWwgLwTeBMQJFh0Tn1YNweH1c/G5c4NbhoNhCZGru2MIugrtASbNuIJkIEkR4n8bbLvAIvv4QI2g
e/In/PRtiszzvtxSFhamDULnTGT0xQsgIjNNC+CF3cAsBpqAJN6Lw1UPaEwA1bU3jJxff35ClIXg
+t7mhcX1qpVakmSAeeWe+kyzt4YBMfdQP/vPHYWl1mh1AmV+H9Iasu6ymDfdPAzpFIkoL7AuWr/S
uRPVatj+2HmWJhNw7Kb3K8EUV5uF+i5esC71h99Fea22zs8yptM0qHUcZ6Iw2P+z7na5fVyG8lbk
sJDTaccYgnlA+5uShr7TOJ6xDFLFeMJy9MWrp8coeeQKNdcxjb04FyybM4kJ2gwHyUrggY9rffx6
1F1nKnb0RaPu761MOCVsH+8H41wj2PKQEtgWXIHmBFXYBAl2z1RRwWpSAdiDZB15+fPXPvXPUplD
XRMQYLocdS04PZPcCxJlFh8EUeVpU6kj3ueTFcWZ+Kdi+I1hsKILiqS7jIOrVM4zJCN0B44Vpajq
/Dq2LpAtcBQcIM+HFd4C4VoNSmAJrP04m6BYPjp1hMmONnbKs8oDvjvGFvRPPp23NI+5L0QUCXOQ
oOM9/l4J5kJd4dPSRH5guCwQxtWxiLukNHw3m5xsmC3Qmg3Ribc8XYGkX2qcS5UuxxEVRD15B0U2
muNuDFkMimIYAUAt1WFK50HjiWoPlEAjmoZSdM7YpdWYKJ9MgfQkMQXzJ93J6Jh7w5aNwslFVWgF
kqlNFTO13BLF3RD2DHuD0lyUSvQrhdsMnVsZWhy7CJ/TMlJb6T3UpD9FtcNL/WR7KzZV91eUagLr
B2s3hjY+lN9DApOW28Vo6vmxs0Xm3m6x6pRioz1QPRe/WoxF5bljUaoxJ3VNjkScQdBMfsLunuNx
WmswxK2B95u4hRTIvDDN+a8J4mxkO0/IkXv5oIxsAEjYsNfLYQd+OWovjxO9zMeVGbBHHg7IckBy
zKF97RUCYau5ieZqEEYR7HGDK+2HD0tCpq4N6r4Zd+tSUUVj2ut2+DoWy+uB+m9ofC2+9YE/7Kpo
IeHg5nHdDmE92Uh/ah/FM62rxwjAlRKsMTYiVBnyAWxvT500vNERtmrbV+2rf+U+HS/054vcCilj
1lYmHaZKzYXHklieSm/85dhOHAGJvgY1XG3P27a9b8sN80XKXYRToqcHetrnd3Yz6DoeuqZfgj1Y
V01nGctBWXYf/oo/yyIAxlbITYwDO49EZhg78/87nEH2wJB0pVpcZr8CC5j7bHbgpo+sb1O0Yhs2
HVd3jgGj7YPvqpxaDDh2zxDvYb95BZhqEw0grWYQHPUDH6K0lLs9f3/PSE8rg4u71Djl171Wm0J1
qJLtcustc2kgR3iZFJm4pcqya7djosxiMcTqvzoYRCV1cEocqjzt6Js0u1RItC9JcMy2onbLRyHi
R0G14a3JKzcSRo5T0NI/jMQ+eZ+z0O2ZuC+sk4rjSArRdsSPXZ44x+eSRjBmG+UHIoRk6bE0MYcA
H5251B+V2NvRhrr7wmBeGCPCoO5KpnwTM30/X1LP7ZDk6/7Ds057YqPoMYXxMsqr1x0PaJ67VPeP
ie3aBzleGmYGIXdqRZdExqmmElgjV5DtqfMxJDq/D+sVlFwp5wN2QMS1QuHspMbnwfaRNCt3i9O0
VeMMskvnECNaIZYEJH0PgVeS4JPrb44EmvaSyrLw+7XsNjottKk15qTDN0Q1L9n/xMH4/a9G5pgP
m9tX2ZjW57AR8je7GRAo9PzAOwXNOhPTIiBY6s7Ao6W9r0NfYSulXN5cCcTEWJfkpT9MuISY5erJ
o3hCewjZJ4Tqt1iG2DmKCibpC4jix0rzbKAgwSX9sQopG2yyD0w3JfbLiQdbF2qE8Ic354BG3HvE
OTkDvnd4z3LBnaNAQ0ZO7NsUnSIv7EelvYmFDb/XwQ2HSl8nQAvnbVBJ6Bc8EkhPeFc9cLvE11eW
su4Q49Qsa/k6grzR1/usH68hVFy8spYrks/NH76k48UzZTPt1VICmeUdFHU2dGxstOcZES4B8SGE
JSC35a+O+dWbIyzBZivKP6XVQ0A0RSwhufDENhlOhoamhhUiULg1E118G8VzmHm3/fTByWmuVPv0
jwkSjDtcB+1hNsDqrxAKr3AelPCNrPcmC0SkEWeFRhIMW0QtRCaRsV5tFRLgG4n6yBA2xCjbd8gL
CzDNfoHF97VEsJgjcB8pKNNGlq/AVv4nmptMFiik5Ee3L6V9Jb3gbyhDAU23E1B0UV3BLOtK85Za
YhZDQ70+QX+fN0exnS/9AKNF4mzMi6bYT5yhyUvJDMyEp7OfKbaTSa0LA1UI6FdES39+8TPVkkxZ
4ARpe3sSnHmLilF+TBFrvbkQx4pDdSgG5wB4yaNLC8eM0IzSNjNV8nOYNhIsNXBZh1VBB5wtGu5r
ulR6WmGeJdb9UsBrUN3vps8CWKgiMSIdw/YgCOyfFyHiXw1+Dcb4YM9IJaTEzEaoudHiIpVmneBI
9oVznkzLUICGCNHzpJl6/g9OwXaYNX8+e2DWMBCynZGhA4IIuV9YHXcXaBDJacgP9hKIdmdUc2r2
j8ChMjRtj0sVfmNKKzW8c31jN9U7ACM7bJO63cWTECorbMp4f0sfDNMehsd4gXZnYJfnjS6ZbA48
OPUQTJcjLwW3mbZd4l/Fyohs/TX0lGobdlAUSGtZajvvpkJVLFnmOXylFBUwIFdtPzCBKIoRYM2h
Qt3vSdAcHFiLjcDNElfMBN7iwY8BX19Qgqi4ZnXI4zU2EqufL1CItNnb5Bf4lr7ZYUHyrvFKzqSC
mmuRMglPvupHvrFqgu+hsR50qE2yWY6iE9BDMcdn6dJKEiHkNglKnafUvBV18yqymYkC7Dw5Kb5/
mbNMq7DEtWf0Ltjx1uKzW1g4cL1K8wwhUGjMg7iLgaNNG7ZbNyuQ4q1aR6PsJzoq2FWHyN1pkClp
5Jk0QxoCI3pdc5F4h4jX55kUXeW2i0icQPIDrd/x2UtppDOw7kvPByxxUDRjZ0HzD7i0zfN+HUV0
bogAaTpXhxCSQLbM/u45Ssxe9KaezOKh317tikfIDPYapad09FTcHDv+fSalQTEN/y/LpuOAh5iD
vKHhurgIKDg3/D4iKu4lFOomzMRjNhzitItHvshzw0pMTOU9uMltWkxYqGDit25yZwjY7DK5I7bM
bsAFg03J8pbtlD/ZDhjeTcr1+IDcoZ3hEqI81ddZRpv4+rwzMcCTeseIFJo71ellbSBZqaJAGv/6
+WV1Pc/PWFONzoX6w+doQbIYH3fmhVHKIyu8p6MYqwIQN+dZ2XQigWc83tLoDnJSpMesS2ilSR3Q
2rsS1nIc0WamJ0XurAWfCvhXoom3/Boh2cPgCWrEUUr+qXw8k0vjKqvao+PJnofbtNYW15cQFKM4
z7pfEmRRui9JuIn1yRk1u/ITyMYxUTzt5SdrkgXyX99hA1l+LYniCCt1VZ0LLwEhhUS9+96wJU0l
IAw1k6JAXvBMD0IuBgfduEvKvv2YWnvOwew9ChmOMwLAUN3HB6DhwyWP3/OLi/LJVadyi0X6e5uM
B5FbbfNZpmVpFngO2xrNdqT3fORFLi6ji+2eWi1+gEqdLGO4GwJkTzy20dGdJ6QslS5FpejqFbTd
+TBeepct797svKdDQKklYEiQjOlqreyIUWzQ8BQbQalHHhfM34NF04hU7L54uc7ybCtmY5RerNNt
hgSIthlAhut19eIxbdqempMXXjk2LLlPIwE29aymYdJ7v9/KEIUFue8z+MfF5VacV/6VZ3Lna/jV
ykZQ4uUmVw4S32upSYoJ/SFg3LQn+rzNfD0FMbQ3LtHXzgFS3SHdGPGi+1R2VT0rth+yjyXVcfSg
GnqN0+KsiX8jdUdZmmDQ/bP9o8FLcH1nPC6cwxmxmGGIIDIQA+iKcb3UcvNvOC6rundcglUB3wVw
N5Lv04dRotSC4bK7+0Fw7k+H5tKV06H9EaACqRsZ1wxlA3iDcm5AmikuOfN0Xvq7C9y7aoMjTSUm
dw+NS+gswa67RbSbZgrXBKYcHpDt19C33kR0epFd2kLfw45LV3hW8fV1zJea1LnbFJTI4Q7JFQps
4O5nxvPCI6pqXNxPnYUd/Gq1c2s41QhS0xXsA30V6N0jh7Wh9ssuRlYU8pA5juZI9n73MpHBBgGp
AXv0SCt9BymhtQIltzlNpABvpL0ZHh4gWIIk4Ee8C+J2Myw1q+OYO/Z9IJvVGdSa84UXCfgLmgW+
YTSKxUjYIQWgtEiAZ1OK0S5TGjkiUXCvonDXBTjiL5oSMXxu0zTGyzKfUdQipijjOadIWzWB6tLq
TvBtHI2C8doCOL7Ler7ODGn7qqssJJcXX1ya/D+OBLodzmgBXFLmcVOKLS1KGANMutgf638rm+9E
rbSfirUIAd3Ues2Dm33pYESGFPEc8KCUe02WxDCTaPryG3PSLULnjX33mWQ3JbAZnjD+DmIHWbry
TZEF2QzVoZGRjoU5h9WLRSSr41DMz92G5gMyFLLNKMoLqQgexEOxasEcazWH5hc+LxiJnlxW8Vqc
lz96Fc44ZUM6e46jdxFABc/vB5gSQlv8W/cSU4edLWPFbqipTGtTCqsHl6UceBG9N7NeJVJuvEkb
BBY2QA7rV7mQfgNEWl/wce4S/utvZi2qJRDBbgNTcF16d3rvUT7JLIxwkm3EL9UXAuWdsDbxR/mX
1Nh30U+Bhrwnh4BFR6P+/l+kUkC0gxfOyb/V40ewN741v4lj0TmUVdXLL9ptvjP7D/LnHyH8K5v4
xg5ugMcXWHPZ2YNzlfN0r+ssYiokZMrOqeuBDwyowCKYemv5t0Gn1ze7zR9koNbLi27zU+g2Pk5G
MgGE3X1bVG47mUuOU7BpnPE2tGNQO/e5Ug6hBi6GDq5GWR9bwVV4klw3pvFE/yYFoMusY2JP+wvx
pBb+0//5VSrEb3bFrlS6YS2A0ZMq/fqxwpWqCFdNt1YKH+yVLOnElycy+uNySDKvDUo3PriFXy7U
RKydne8U7i2C7tq28Ac/cNZ1s9IV93IHwqL7HMxKd57ifNZ8550fo8CCyvt6tYVLiD6OCilCavv8
Qg+JkLTbW3ocpiy63rlzyOCVW791yI1Vgr2Km/dybVlGM6/sPnTXjyqk0in6tSkGW1VSweTRdaNK
tlEKCzqtV0FvaDv7FimXfW1EGpWwTohn9+Td/YFhxLpLlk8pr9ma7Si7fNpHJsulk9uWBPBHI2mQ
VxGwXLTZro+aSxJqHqCDDbXA/jkToD8yDtoXRylwhWN6EF2X9mEpRSF/nivkaQrYi2462Bk2d1/U
ARZ6Ok4wCD1uhtiGzeEP+gsxF5yeCqiIm+ueDS9RATYx9iTzYF5kQRly0JoDXQCMGGkCDoQ8/Zzl
b0esSrJ1fL2hAevNj64wibgM44b+jbBljiwCagDzltMXSeeqKQFpOaBQVtv9iGrAhLCKELI8g8oM
zmxaXGQR+PfrXt+HXjV16PvkSKGKbgEwdlNv3YVjerI35Wy20d04qmSkGYCLmDXRmJ1PXIIK0dF+
NcUf0w9dYW18VOLzXemvcnnY6mEQgRUs7ejRqhBvlsTYulPMwwS8mHXAhScHQlAgjYjb6p20ckSx
yl6C1W2xslaxs8JAkWa8Flhva96B5cRcqeiXVm6cNRNqFSLUxGJsug9U8pZSu2rbaYInQ19bIc+4
sZKAaYWYZ3Rx9ZD8zrrVEDTjwsA/nm9y4PdaIV2U4o0d2aZB3rcrvOUHTbaAmFPPvwx6A2C7hfxO
GKPPGUIEYWC5gkweICuIi/ergyFHLhKXm6jmAY84cuVdgbgoEeQGdum6q6ZT6CKpAq0LIy0SQAkp
Jvjzrfe7204sSZO/wCUy54Cmfn2ioVJCEvSOvz1eY+yFhwdqHJ9D9kFlff7r1S6To6L42BAW9kPM
du+Q/nhXnsfdVAKKfYAQZ/wqoNlNUDS50N4cHlsfEZIorpjmuxw5M1vQiHnym/UEpXAKZR8/4L+o
oI0pVRAYgcXGJudHqS0eK6ZRe4XHAiknX/On+1mJrR0pTMN92BIdf2xfNxAPsBqPUHySaKikh3bQ
aRr4cKwPqiBA+E1wvQ8UOtRiVMll9oDClujRTpTT2sPiQ7zkkYO4Hpc5KkXUvBgvL6xd8hNPn05k
pUbRZrNNJ2wVLK+0BTEQV0PWYJWaS68+5B6jcKLpgRk8ejorxWdmRShFBUOpXTcpCTy+qvoG8ixL
xL5X3+Z+KCv3a2woFRAs1pBUsMhd9rSeClD0aFkdwh5fBCOy+037fatArBENh6rIXXv3bwxlw3LF
nH0HRYjxjpo0/GV7daHMx7bsp8WTD3D3E8fGEEhV+NOZv1r2jKEH5iPXKCbKQBzPToqe9C/L0ubC
pQGbC0s/kym/ZG+/SO8u0GDLDHMR3RBTqsAgw6eBSeXsgBM3uPF27m/GNxq7nCg3X8DmW5jEH3sP
vGIusWFPzoCx8C+ikEug+61d6cbFWp8OjfAIDOGMBInoQRztB7KjFVjYGXG2dbw0SBaDhkvL0raU
aujGQHqwR8AFNkLSirGOLKIxDsygQFJmiYv+fm826MsHz3XvyyRPj4+OVPErM+kghSS9pTo/srQO
d2jXdViPOhAwctxJ3TzgwniOSB+gQkd89Dqb88hSOckMOs9ucr0nqJW7JLpwUDZhC+nvrqAMIeI0
hGp5NimBjkAIZt3BWlwDDKdhlQHFTMqAGd0+uGlYmskgzw922ayOmMVj/xM9tqf9OWqDvZSOzg8D
en4LWXPynTzx8NnUeAddbp8xwslDi3PjjdlIQ7nKMvR8MsW4SxQNaL0J5S/5gIWE6Ovhf+m18/S1
+5CmpW4WZhqecDeoTnNpwvF/+vOzeNMpv0Rad6o8eVWJrnBlAxyBItWmhA9pAUbws7SmHG609XXx
GKCgtgn4oezGY9TBCfaD/oK2N/k7toBAaI2i9QRWQL4gFBDF+qoM7WAz4vwpQyFNKdNRG2etDIiG
m1vDmVpFjiFI0SPHsmaUOsBujplIdoTA8I4wmTxP75twUQ2RDLyp2/Ra2/QtW0zBvFDD0jU18g+f
XDrPrDsYLMu5nPcMJk0GbZCAN5ByBwOV31/F8BlricG5Hp2eIuLjqEQoiRBp4I+LwILQLvgIKT6V
D5ambDIssWRsNla0wHpfeM6X2K+PBSeTMlpG5SKlUWLOEpXcTMdgsD3v0Yq+ndSq3wCWygShU12p
gie1BBt9x9Aqrr6Y/+F0sumFXCeBUAeRmNC2JhSxQ19NENSiTzFbzsvX00dArXcqdL5kKSLmzom8
IYcgJP7qiV8rrpqTuv2jF9HNW5extNufMsrj0YoqnDeSQqYTa5lOV2qkqSosILKHpj2+3Xs/a5p0
rYZ0Gjq5ZOCQy4Hg1pSDGIHNpeSgCLyGxSjhn33Vbfw+eH60+yM1I6DnaOypU/HkX4aDf/6gJu6E
D65pf6Q1EzMhML3ti5EEejU9bHiEiDG5W8wRFxkKRdPQ2pNTbaGn9W+cGr5US2YKyHF2M9KZ27SO
lHgpdH8OoYPKpzrnu5MiqBCiCW86b+uuM8NWcr2zbqhfMW9l0wrp4/gUL2AqBC6B1wfXcblkIyB4
qR0lbKagIZ0XedqsY0OVsM924qIIx+kf9wi6vjoKWcFMHKnDNUKXgW5oJedOWW8YOPRdqkUjpWE5
Y6iSTzcqF8ix9w+4n51LJ0D5oNAoIqpepoEDOtDQD8ftYgXcml8lrLZ63pFFqm8wRH5KsFyYG9Ba
ZoxJ22HhBbeXHYClfahbwYNhT5bAVo3L/eyPQgsJEqgIwkOsSUQX3ZhtCZj7Fb8bOmTbGsGeGnYI
jhGuGmrkz+WTyg/O6v4UTd4AZ7x+86Z+GzBkeID89rbkkSfFB+gG5Cv0IghSCJZ0VXN5RyeZgs5T
oSL1GSEL3ScQyg1EXFBfZsJRi6YZjxeXVIiA4iYL9dL6NPe3ifjmXMx9zDKHYDU6du2X3z448sDL
14/vri3lHwiseA3Hy8oQeTimazxA6WwOcVK40QpCE8pLGEPzWcnq9BZutySIBLjMQ2aXwsMmxFXn
p7/oh198HOehCwODbSMHKVwXY5uGsOAZZHe4I3PzUOmkXwtIt+AB5XmzFFgmW4yDfPmNr016GiwT
UQMbCusON3eH+ZYLx6qOVzcYg5rFXv+aoLkbVcxtQWhzX5tmrLexQPutanMKuz/fBsBLs5pQbOki
C6Pu+5ce4DnRu4Z0g4ktNfg0D9qofU6WK5fWALIhrp49xjGOhaU9g/FKBTo16uPSA+lhxL4lKSfs
CTgCRUhyxh9kVmGnJ0b53fHnb2fv1yKj9gf4KK0rTLycZN5GOENrqOSsNKDLDIJA21vfXT0FZ6Ln
TZgKzPspTNNSL7ojCnSJqJwY27XkaRwCDlOzZF0eDQcmQi5ZueDkhVZHO2Xvaxt/YVf5lyI3GcJM
5oH7DTr6ZE1rgpBkNYZXLlADdWf9Nkbq3cMAzrw7/p0fqIuYbVNDTQRn/519wLkd0cRxe346rPep
B50rGAw74gknKLJUxXe0UnXhkZhFb6oaTnZM031zz40rhNlsLTV//zUznx6X9Jm71YqyeNyiA16O
wXt7r6ODMqcsRB6iWj4UfX+5mBismzWcxZd9BXziKevZMYyBdomKg/Yf5UCH3dEQU3WrfzBMAwNN
6FvnnVsdrJPNCbzVav1B0p7fZU81SesJDzfk27BDsWR2Jqz6bHMdOPXi5eeUA9xWxw2MfdiVeL4B
cSh35eiyJQJzsCPKMYgseBiW34adh1DCm+Voiw3Qp5i4bOZ1KC/X0ryIAjpMHVOa9ZE/5szsf6J4
i1X7ixARmgAkARguPbwg9YYca9xt2/ca35g5e+npeiY2AgsA876lkjOWa+WgNdqpg/+8kv+u/5XL
kIQFTGgoIyFoevWoTZ1y4H5LWwLOWyizBYkvkhk2V/nrBxj5hgN1NYFtk7Fv4/4MpUKcrohPL09q
vCLuQ92Drh/Q6rLBhUi4tcTs6/Io2Wl1gJ8HVBBiCXpMjDVPbDyviF4BKSjbKpAWqJKBaFZUzmhK
fPZEXdqu+dEBXa25NyxklkJLuvwxtZummeIuAl9aMJ55nUgrTKwHdZ1h7qVUQq4WxMj+RQMUs6TG
qNZm0bWL05UnPI0YNsci1KaQMGxtybz8zZ9fzTH7miI6K3kP0FFH89fxXrU6RcLrlOnQcwH1v79b
ff9dvpOCvVXDClF94CaeWyrzMnx6inhDrDpdPF8NEGpx7mtT/FjKOEUGCkZfR2MGwuUk4DFPM7vz
zuh9kK+9UxhvoCsinaqqNIvlth8xk9ihWn88K1Qajl05FEXLxK1hgAM1+y02Oa4KPRdTq5pPls6G
ZMGYjv5619fE7xo2B0uSeUsGKeZo70kCGqw5V5FqJMrH30LNw0jgRwE18J5sTybyAmQ3dyeYyly6
4hg2DSmjWoW8OQSKbnbaT48Lz9vQ70EFMtRN4NNj+J77ID0+ngiUW0dbHmheHylyDk4Rn7PfsXr2
uJyjPreXtage2Lxv0ZU5umswojQSRW3mBhW0Ce9QzfXNdNdtAYSOBs+H1LJVSQMaS6NQw3oNFXSH
tZmYQFIS61bwJd5NWUS5qCW3OCS+P6WjIAlvr5lPy7Osb78523a/ASMPJPi/HyAe0fYUoIXBD/V8
YbrVQnQnmtfrybLygHrCDH48EC+DebYtbs/XRkqrxCod3Qb+wUfRNCUzV1nkj2c7UB5awtKvm+I3
Y7SxO5SafOalVR0SZ7LEWxyaki9+ZTx3yyPKsqrWV4H27Kjm3f42SRvi4bYvkjMsE+4Bm9cb0q76
qqGI1U74pWxzdIk6er74v9CeD/3+iCSp/EdoyWt2RdPjwSyqStteeGCVwZWvwEnZ61nVqF8RytQr
POAWbAHROrdkjtck1sVY9H8v5sDEFlUT0v6CM9RSBswP4NuxZfR4+eToueS03UFs3/ftf01khtrz
O80mMj3ok/qx6wGB8TC5a1i2PJI6noe3nzQCA/WmAiezUAsvMavg4G9FAt4qtD28dY+omutciwNA
tM7nuld8u4a4vMVT4FO0GqLQyHPALrxLpa1O450rtw3F5BvakjgReiH6G5FAo5EHQ1GKjaaitD47
hysQU47b3Ndb+kg285/4VFTLQHgXcLY/CYQRLrPUJ8d26lM49nq9BkHTpHek/QXhNO0KkmHwmhLc
C5gi1pIvX9HB1MfTcsRkz4rVKxOIMfd00rHg6kEJ2UqoQ4C3OssaYd2DW/njH8K3YpfNmrN+boNd
v1Trm6AhE2aNqkdeRDtEWWAJrayhwoDI/yrSj4OYC0VZLB/4WW5Tow/35iwYE+TNwd/tyN/Xh3iI
HWnpA8eSaYaBPg910zU1z4aM2UneBOdlBwBiT9s9d1P2Y3xcTvWU9pSnFlCrKOHR9XxXZMiqEXR3
1Xs+5UNKFzvrzX2Y2al2vpFvkRErLxShwIX5+xOQWw4+6Beduz2uJLyDA3ersv3XYfSdQafSJH5y
V7dFQxVJ1MtkYDMBM5xbxpqzcCEAYVJcMuZPK7Pi8FAV9Y5PaGVzmi7r6ccibCggbMhPW0x/4kK3
u4QSMIk/fIrQQb8aQVJDQ8LJVPDlIpbnv8nP5m8dz8bfIY5xhV6FNZikeOCnaXjUqZHmR/RDyLcS
QP5+i5+lDSLwQy/SaH4sHLGR5qQnXPpW5+czygyoyCJIqxAK8R6jX+I3P4fka+NdnqBadwzgkoeL
yrpA8eM7Ro5ATwJOgwwNf2LgYudZn+NcUcSl12OfKSWVPNnSJoETLUzH4PDliCi2GQ61yUbLWS4D
alYfnw9FyV5k2pIYXc0Myz7i8mDaW1gbIxhPl1bf0UKKIBylwHjS1A8q2NSXjGF4LamEIyrtCKZe
VXsJOfr4lQHsksYjkmkJZxaKoVq1sJqTVMfBUOlq2ta3nLU6mH5clvvwlO/YFc49KactiHrBTDQj
z6E9lgkBwWzt35UNESW2tjQIcZ5I57ceZh9k1ZmClYLt/C/JaRFT1r6a2ZfUFLiREbTbC0mcwWqZ
Ud+uTcYLnPIxyrm6FSJ+phgGzdTpJKjyyg6k203IGqSxzvVrgmYNXHN9jO/Du75M4rGhfOTqyL3c
wcOj4hjBjlFj8El/SkoV+EkuGx/o6NPTF90Nraq4LYoa+dH+FWTW9NsvK19YFYFD/zBIvU15VjS9
iWUQEcJnFjbdRnrTasCvvQsBBZY0YDsSzSvAMRXnGh86CScPepo8ebe1CHIx/MOBHZbTF/umBdH7
E/LPnv5pIzwjIVZdQ0qHzjCzHW4MOggVCXnPldh3FDz0Q6kARobvS4PBG6lzf/vvG5vvUCYC7+dr
V6/sdmpqvtafSrMW6ERrLp4ivDBfvaPDC375NZU5K1AbE391jcjZPe0MGlPTBngsw7t3V62VKCBk
jPmzLiqpJCeSTIY/z8BXhuRlaYettX7voStf1xslrteRCyHyRXJ0e5+0uHXDegO80CZZbSht8O40
KbeJ5Om4O0p5JX33JNFzNWAtsKyULgBlASVxQPj9RZFqb0HVFSEEb537+yE9i895tzBGt8uXysuG
zetsmf2VJIjJlVd6xaqjmnxoMlvmOsy/raDVvV8C8lTvSh5YbOi3brouNaP+wVN1h+pRRkgQMDb9
Eye5gzZh/BhOugr6prcUYSQLjCZb6XtmoJ87O4po7sdd7CStrD54jguJY2JmMg0k37EsUUBEXI3G
nBBT6U69lqQZyX6JS5GWiwJdUh2byGMXjtcRo5becHvVepq9GFuIaQi21MnD22JnVylz+hJXIB7G
5dXBqepH/dN5HLUbEbCvGDj+k1HWrmMgWA+tlumaz9P5RWt9rhmRAhYG3ATW/V0PVYEOHpitb9N7
QK39nFMCWt83TR4OkNBihi6gTlBXhP7Ibe6NffZyeTh4/s4mV+vVtdKfXDyOth8KAjiCzxWyaj7d
m0fL/7MRob1qo8yM7EedytC2oW5kAKAgO30syr9v7MFSLGzPaV1v0SMQmCCx65FcRUJz9xPsOc+p
hq8oX+GG8SEMZJz4GBCMnSSMCW7kJmBWjakQKF5OF/YZ5J7sqZtGQEUQd1HvYoWYQ3bwhOn7I2Tr
+PDh+wra2HFCb5XhRiFuB10Z8iZyd7x296IX0k2ygOKucqbt9gl4VgPdngxGgF9SD0DDodQHh6si
fF+sRZ6FDi+XavuPwem3oZozhx2DSaizX1we5HnPiqLMIw1Kc9auh5vWk6NwV/chXU3/fJCthmCT
NMRKNqtl4On7BesZwFMoGAQKX8MPI3hVTQQwpwpX0bu0JsL5/fIjcJpOVNP4P64TXsDAbbQ4qok2
NcxwBV3S6SWv+nK7Dyxs08BEees6P5VHt7ETKicUUKgIGhUGJ+xIX/FMsQTfiWUTlK6Sdre0sI85
u+B1Bdqk6a7tJjVHXk9EA1Zxwh1ckVQ7Vl8NCRYaoUL1NbaNmbnl3QbA96QSQh/lySzfwcvjMifF
NyBk7sWitqNDQ7allj4osFB1uiUw7PcE3ok6AbQJvAYDKwBCT3Q4dorE9lby16BDuIXzaHjqiOVf
qfc+zKG7yU+E1j3jiuwMjbKJewnkMxDM5CdRBu6xmrpCQSXeLlo8dxMHf52kvInvN8BmuPV892rP
50+A+7aSYt1H5Nue/UWuDmK24P5gVcZj5xJv9BOiwmMZX9ssSazkU9XcQHI5+ZZ75+OUdDbGe3Be
ieaVYyKX7VjKQuAV5Gn5O7D6gg1BqZdKDmBv1H11TL7kfqpS2Tz+3DG8U+WkIQ0lzav+i+kVIVFA
6zWIUQezFb0DwhPS4MJgp4As4guoi62Q+wZ9iuCd3yye/LzYaDDnIw0ddbz+Ok6GU7pk1hLm6PyR
PPWe/9ctdSAeKITRHu3CB9dl+nR/d34GBg7tmXrvtCLOgZjGHjyU9EXtdSHs1dxrAOuIpFXBBaFH
ODxTjwNLTNGZAsVyjNPcXq3w6UP279KGHXAyM5Q/Xtnor9BW/L9Yebfl4CXOHwo0HJWuRZWc3f0q
8ZiDSFO1+VsfhPc7lZ+8/dkLuHZOpuir4KHUHTwl4IpMvtoogLtizwRU9zXJlYPFmNJOGuCaOWeI
a/icZicnLx5RHPDMxu11d//HCeoXZdVpOLI/uSgqYNHrnjfXK6FlPtEMtJK2o+bjt659EnaF1w/W
xioUapoFvsUk7J2gO1EYh+A49+rm0ghQEiE5gHPq+mo/KC2KcvcbMpxnf7CbDYnbwqo4jMHKkrhL
BNnz548NYxmXHD6M8ygoPKFhBNe/JsI1XRwnLqD7Czy9a0WG4cO8Sma6qo5zdm34A5LL6FJ4IjTN
Z9GyxvbJiiKWoB9G7F9UQ4c2eDKiPxkqQcg8+sL/JuoqZID5p2zkl0HtF9W7dSKq7yBNJOxCHV/C
s0qc1TvV+lTQMn22ALX1XFTMCMy6x/+U1VjtNnZtVV7y6zjtQZeNQqqNKVGqVXdpW41cEVmkRHJ3
qdekH8I89vc5PcSvE3UY0uQzP7kQu7uaraDgJjLhlvO+8ecH8PSs0QvI9B93PfzMID+frOi7T584
08QaGEVxsUiN6xnvg1a7gvJke1Y912eJ8uQmSKAGvlG4ABUfbKsZDbvnG2vEtFcnywCG3EHCpPo3
7pXmD6gJ1Lu8QiEnyF96QKV0HjEFk59+WFqSab/cuo+++1ws9eFv8kvABsbxjc/lFUYDp//YqGcj
OUs7EYG2QxxBqnF/9kLuOlUSKazCe+fpoJrrYjUJTeQ7FcAZhy9rYpHRCBZdsfCDydpYJjvKs8fX
iSZWKVWSmEBC3YyxtcI6Q3MLIJHH/pEfqk7FhIzhMhR8657zBgpedr4NurKjRxFIuNP4DFs4Jtxb
EAl+MGemPD2O8D5qkTiqOAlNpjWgNkNEuIxvVP9BrrbXf6MN0KIBYzdd3NZ9BCjuGO7RScdTlsVg
gYDiwSMgHCF25uVhYJr8trXFrS3Dx8abREWq9Fys5E69Ri2JmjM86nULKCjZMZ++b8vLWxxo3eja
W2I94ztm26gy9Nl7ecLlLqMYOqopz+QMisUdx1hCSelkEICzyD6GEWb76LYCh3IKUmnEk+rUJciP
5I+sZ2SyTRJnINPcI/EQ+qnGnOwLOybSMhnCWvJW/kmZ2rKUUPj03TIGQyQVr5MJhj+6mCGUIExQ
Jb+/vZScYgPUbBPChFRNPIfcAcx0x/kslr+7FSNLSKWJ/RvBs/kDUXptxX7QLfsvYGxYKnjYTmzN
h+CETFCaFIom5o004PDMj/usqVrhXhq5l0d10Tqv20ksGxyo0PGyabTLLnmEn+J6+j/5MtWaPnrd
tcl/G8nz93RvL0WgWcVxzguHMckxJO0rNNjaBdvvDscNBoOdNvCvVvrNqAFDmmRnbkxTJBjg0Y+z
i15chlwQ941eP3ed0OgoiAaTSw1xOcdU7lNlbju3uaZkUKRwVGxP5boeSnV/asBzpB/IepItm2hf
oyZVYNR7TQEmJJdNU+S2bd6W5PklkW4sIXf2M87rq2LtgmD+xo9GdgUO0CtPc7lRwS0rhCHDgLNW
lFjxkg2D6Pxmbf0KJmlmndhWSNn8hsfcluKjrE2e7keKmTEUhvAAzWSz2ivAAnQMD863a9PPojEL
4Mjzqob4MWfWXXc0L6wOLx6oAfz1yfVep3iWH0knc4/LMMOBc0aKYeVkOCvxOIfYruPUVm/9KUHH
fl3k/37b6yaKmuqdktA7SQjPJg2l74GRKaJlJVdU4+FfD3ik1gL4N+klim3tTYiUIumpCHzc2STn
g9OX3QI3UmN3/twS1JXK4hFCR/7AAWVvZm5RRMuNjSSc8UAQ25x0PgGLH20BJhmLAAG4se1h4To7
4qmZB6SSCXgHWwg4bLIngrlQSjEpp05CeHYNNRN2jFXrUdIV6RwaPVKhohdaF24bVz9hink8gmVF
ZSQbR/q1l2ZG+aTD52ACr/pHdyxY9XKSA3+sJOlgyBdTIo0P6y1xe+qfRTbMg/Lpk2VirR4Af8g3
3Pn1CJ6/Pa9CEmwwMMBs6tuU813yFId2ekrI+G2BQ3YdXeeZQGRNRsZqBLvzXp364xIiELpKwgfL
h9oPAR9FeOCgSNY2GxqQV1p39xdeWjtAyLrPSXW+yyFw89csr4+K9gL7a7+E1lP3DvPjoxlpssQc
CMkRk+L8HjxldpGV/dRKJlsJtMRQyXnEpcKPoFx4NhwoyHZUzJo9+2H6q5dJMirOBMbKlot+8KJ9
NA1RDMm2XBcFD3RDuhJP135Xzlxqtlf1Y4k162eCXNrIo4mkBQuzYgNfYR0wJIl/i8cGzx794AFh
75eg3do4L4HyNs/TrK4xosK0suceUTQPumWCij09CeObCWqXmKKNDqHcz66g0YCmABmFzYMiGGr5
dyfACulHoTwALQOqL9oL5ROsWfJjxCiDJRVE9gU5wv0kOyMsPbBvX5cX/KkH1IIUPe4uPDlE0XBs
PLrpuY+LBTMFNeFosgOZn1foooVQgNk1M+jTkwDwoNy7UoIOSsBHBYKuzs5Bh4CwZPq3moEaj3Rp
vllfK46ALpuEh7dKAtScSuC3yPKRxfyGvP2wxeLphulfDX726o6pmCyG0HSaCyses0TDeRj450RZ
+uz16hNWB8qTQj24SacWWt1+Ecb9tFalmr9sZYpexspKUupXghJW4HZMWkBxbxT/nlI2iwZ+SQ64
JAcXrzO5YKEVJNbvZM5/ePAfBUc9/CXZfB1FOBtai+b+YHXv62U7ECFqPQXZ6bmlfptsLAA503bz
DAZGA5ldd8VDtLQ5OyQFDgtK989geW7bmf/He9nVV/i0382mjMSBuM0MbJFxQxQa9qYx+Qke91fM
ex+0fR0g/5rwPoN9awwCvFM74TZJfdmqX2vGYtE8BrrWGs6mpg2BfMhIg/FjivfqySPTtkmlBpRO
O1Ipt6c4cY70Ljexfe+tusg9/r2+T1Rx6nnnHiN4hl1bSniA/Pq/ETK7sGKwKaTmZlNYCcAFiE60
U8GrxgSYOi0vFsNHm7kL0dTQkG5rwIY3v7d7dE6lewjPLhUIvme6feP5W3tPQxpfgsWmVZEDxUuq
1q4DMySlK/Ggq7fN15KZd3Q52mRNxm55hJsWlOTq3tQfvOIoyTbFJAhhDSR4Q7Cns/daW9bzDRs0
RybwNnORkZZLgzG68ajTl7/AFng0zVbtwh8+SfocSG9Gg/r6dSRB1ivfRHSxMk+ThO+gUPJvl9W2
2TDztxdqP9EGE6gyFw0uDP/8Juqi6GbdeKzQGU7xtzSBHIMuQu6qsbFAWMzmaaWyigxErfUhBPuX
+1DgQPxblI3p/fD6QQOmg/YR9e1IjJcwggPoqy2azIUmNBMDUy/6iLXWi+HxwSWVBsZd1jaLoAE5
Nqnql980AUO2EFxAle68cwa27gyvOW6k1QuSFt0PFJDHVjuvHPThDeYCks4RxoRGYvzVcWIzATgU
0YGW0g28Y88UmUrqnLrofhpEcQqpkDgfIH5CWPfOPJy69sjDcgC936mZorDPY7Dv2fGdKMH25nFD
yLAHR0rRie1hALNyKOxKvvbfIbQXI2rMw/QmsWHnrK/QOTV4SIhPN5sY5xQYNJ1VVyCUI2xTkJ4c
hRpKI28WlPjTBHEdxMI4qupc3BJruRpBm0yk+u6RU3yeJAa0d2HFaq4oAaXq2F6wp0JFpuwqhgai
MwhDDPhWiPhYpL/9rhgouqP/srJ+rB0jfzPFKN5byAlkQ8bbj82AsoQjiPKw3rqVOwi1acf3M8//
jUITrN4ltj5U+MVb6D7CY6UfLlehl0PIiuX5vHXgIJtnOquHIBBuXApz6afVLt3stWoAW7p/1Zmk
fs+TDoeB+PivP2HOc+aN7aTDroByNFSnZD8SM1o/pmdYnB/8kpj8MCsftPEw5f0AAwaXxUB1dP38
Z18B/+OWzpuh9QT7JCtsaiSREe2yUyPfUzWTov2QP6FEJ8tmGV+KzQldMCiiVFEtaS0z70cyAcXG
2Y48dcrZWV1kVP/lPu8+qdRbXj+QIKL89JDMK6Q6EBCikgNgTPLkWHsOKHBF3rG61weOHRcoq+at
8Lsd5p67Jmj4t7qHfEPE4Dz7rKHEaTrOPLTcQCX0z/cfO0W8q+XylMl+TlT/ao8f2PILMIJRwtM/
1tpQpMD9GEw92IYw4mKcZxC0s4BSN66BhKLNqHU+CLLIvZJNyAjJfMlWXUVOoEoM7u6YMSnlmjK0
DIAQjg5NFzyyFTM9YwpHo854/gmhB3Z1lq7Xch6isIvBi5n13QRT6Pr9dK8hMirArXMt4X+RDom/
aZJiwYBf8IE0KA/iKNt1PJGTZ2yvZ03I/PiVgI9vUf4aoeHgEzWsBEoNQWjKao0s2FA2aUq+8BxE
mtnGVhrShLtXbeMEXywi0IA1m2pNk7BppgNFr1bdIPFsM5wE+MeftnhH3jZGfjGkalj2sp7n09Pv
oRAoK+4e22pBnlBXzafovUkt2XCfhmyqRUzjhopu4vCus2vPi0OYd1hw3ifuXBKd7TOx4QlcBo5T
ujfRFxSAWX58F+CrNQ/xD1FQj0xD/JFHYsfumyCfyeQwmikbWIBoLeghZQfuGbDcoEev3+cKwCIV
1LeU7jzuko5IHNr+tPoCuPHrTHO3roJu7xCbRELbPdHinajNG/557M6EHcQMe+u+ZjCi/Wnzv0gv
VQzvuW7JR7IJ5VHlkKXEnEMA7CavcvtXLZDtclLCWGtp8pBA6uGZ3oBr1gab/woyAfusifzl6aeB
OiwhQdZEToNdmkodC8B1Mf7fXZz1QHTqAKG8wpj+6R1hUEhgDCX88qHhCQeAWhNMHnEC6rm8ij76
qkQusnUy9RDNE2um+4eFa7f8viHPU/0h/CAqVA/SkJi5cI3lP3ZXs4gleKjGbEzA0NGNeaUtIeTO
qypIpEj5gU+jZbK9FFgKXgv3vnFPoXACudAOHobE1YdpwXvn+rs8OUli6SEh7GAr4pbX04qhsClM
BWl4/ZEnucc+ilgzjxF25ieQ5x8zI6Spy25hcqWtCGHHGlekidLIt7A739rM9Jx6qvRED27Brbrf
uGRWlC5zMPSNHkeySO8i+Vt1tGLKnpSSlHqY1wJ21612YfLL9XSo/wlJnpM6vun6AU/BEqhPuB+r
4joDCd5E3or/05oT5JkoCXg2PRpaVBSL28v0GdeA6ky6tRkw83cnIi0WQ65lCge5anaTKMIYjgNs
ZFU8f2wgiDjql/tuuBSXrpKYMWyPAOIRVgbrMQU+VstxkjX9vYBx952594RS0Vh/nY2GGdYKD4cC
/SVAQdDQ2bKEWK3QeNDP/WoB7KGD4NdWqG4c8EPynrt1YTQtQNqn0aD6EBzvMkANvZ5562rgxLN9
6v3turECjFdjgcgx06UJtxVsn4Z9uazMOst2eDVWvkv888RnzZfTwtUWSezdkhFupqXeYahni/9R
FjKgpicMa1DAyOUjqXsG2G9fgwIc370T5zea1513J8HkUN1dyAGInKJzX6SuWafOMZehH9yAOuT6
sli6bja2yjK3IjmfE7BfdGGJLvQfAibkKFVIVmuOL6h9asso5DF/i8GSmeYwbRTkLVdQZ0S569OZ
QIs/X0RX9XO6mrQj0vxEZABWB2+A1sb74MSoqXYj3vEIRQaic3rGoZ7t8ffTWCRgck+X4Z9gl5XJ
GYoWIaHCjm4LHRCtaDTVIDZKP+unGsX2S1zHPN4R67+WvRL5PiRQsUUo2ZA7k1N9UiR+mMemqcp8
BOjOoGyxjDEA5//UG9PpZwEc5Iw26xnGOhxIEPnQGSGz3quXHYJ9H9k9i24PCof+awVSzBb8P6zr
vWZoZi8jiizfvwuze5fyklAopIhZbUlJgFk8kPf/QLXlmdV2y+AbbGG9DD3mUfGTygklnkgurSbb
TJ5KBs8r1mLm/B4/dx2FXU26GzVtYumMB4P4U0zQtFDjDYQGMGnpTJJQazZLXl0vxVGV9g9mQdPF
E5NyhTOybQNpf6wnWnFit/S8Rra3tTfj/xR0/5hgojiXP9TmLpAurOgOwwvoK0FPp7jsreNA+YWt
AOZcKQPxsQUTwcLRK4aYyBWX3s91N4antBN8N2QPy8h+vdntTSclTZU42HY6S41l0/QhgpLraJyc
eb2bSZA9lnbZBXY6G1PnBvmDJzYj7ZrI6OPyLFPF5BHpmkRFNgxxvmN+oui4GsBU1Y2xooCYtR3P
MrryJXHn4C2F0kJXQDkEK+L96CJwc3hlVirHlB5qBi29LppCzEjJOymbwhkY0/W4qPmaL8sqbOPB
OVXzI3Z3ae8pq9f0Aql771hPq84Z3+E7tXkqlvVpGJKEhkEl4SW9TinO1Jb+EaqiqFgGoEeE9xkQ
UbdMg/nKKQPJHGrEB4QJZC0t4wM27mYAu1dqK9aGWPFS+Irfg966qP1R4qwZZj9jvradtYgRYUD2
NMxcc48lkvbGYATRNawNrOFWK5EvttvdBsaHyiO5TbJAMLmbwf0pB6kn3a8mrHJ26TuW6jD+6arr
eI831f/N1j3VRTYWwpP+BPy5moKWPDOLciqe7TWTNVt7SxQnQ6T3JI3lahk4gezDRhzdH58+Spvx
yIoc2S5iv7TuNVJ3KPvCSeWckYfrTUdhTG686gVsusjXHR8B/Dsxm4TMImU53+7gOfFhWHIt3Wu7
z9+/eNwFGNbbJbScR3dtneS20gn/hVT6VZlf7WShxy5Z6ewfj9NQQqJZiWnUbgMPxmtx5mRWQO5z
yP94EfKqbj3eH8HeYjsiftipnaV74oYPatc+gWUJhp+QKBWRtgwgpw5xmg4RhT96kDHKfPpTWMhp
MGtlQYc/2ZNggqr9DCnf4tlPuD8PvGPVBIwjBK5Y3dKSoaHT4P1K51hPjjub8N/P9gQ9VvU3dARJ
otcKFSChzYaLGVc1ugc6hpBC5JSU1itREKKTZG7WlB5YOmXPBkkOg05I8gypsCRTA3rto0GT+bb4
9ChVUnWSOVwomJDaZVNeL04dUMSezQ1kU6Eusp3BoX8y3+fAKGmO/0I5mZh+Nw4XUzcz335nx4Bv
ky1TDILp7sAnYvyMFEl39I6SBQAyL/1m4j737GFoOMPvG5BcUhoznV5VbYPMM/B5yGj94oMJyhu/
T5858RzZjXrAKzkTSP5tCucL5DQ7BgictM6OsgyqpZGnj/HZexOFqk9tlysw9TnMyKLC+KVvgiMf
rNyKKAs4V4JrHCceBLCjcB3H8Hypvo6hk6gIW6yTkPf6AgygHbct5BvoQgxliJprHVImLnR9Ha1B
a49HuGOqUyf18hmxjd4ZdghU2P1NZ4vKEIpDCD0gtfedeykS1nIxkVFKN1fPiaRw+kQ2oDMEQzon
R/pRHe2Vnts8a18O14Q99ukiH1xmNokbtj+99P4lAW76YaqyshnSfyXb/uZDQAM9mt2wfclW5shp
04GdnOEfPIlYIElOTwPppusWrFqvVb7GEmJfaZsx5GFzLbqqIaQ1r90Mdqq279YN/4T/kdri31k8
Swd/tV7GPhlkeR47WGFLLXFspbuDUz7Hsv/iR2abijO4BgtiNKxngjS1kSJEJ71qCxhXlZ5VT8q6
4I0YWw38Py9bS7gDNn0hCfOvtH8v+w02kxeJeyasv/ZThk6rjNBRPGR490GnyznIHFHDedHW5Hm/
sVORk1kyfushrOwXwHsAWfDfnXi592c2OHFIzz6EKJvJQnpexzojlAb6H3tbgNXPFsJe2O1sFF8T
O5FT41MFiKdCptfKn62s9In06n98tQ4EsEOapl5HB0lTYVh7b/jwSNZzkQ8X158xbApM0PI4UAF9
yw137iaIHYJR435ZHDchuzalcjSSmbMVjO1Tt5Kdq72mIXk8OmrOGQv/NCX1F3Fyxy7Vbfv1/1+H
7CRugYff0GOy1w+oPyT2Xbnt0i5qvLylSYIj2TyJjT6Jlz3CgktFuCxBGjNxQ9QYZQyvW8k9uwfR
c9kiEDNPMxojC8/nVNbsCmk8y6d14bn7wu8DgW3pjuw+hk15UhpbAMlf95O96QGeqDDNcNC1SBDP
R++wYTQejsj5njcG2eu2K5m2rRMHz7dvFIgAQMPdQ6vzN1FxgrmxlQOsiSvbRXeaO/RuT/EgUTuD
tSU8CUHOam33AjktZerwR/XhEUDV6/mzEiaYiu8jwMG7tpsFDm7YcfMM4bhFaG9tfYAtK6Y/2Dx2
Aq/E4tDhdCc8bw2PvtFHI9We0BzYGahmalRrqkW0W4AMBrcB/0Je6ljCqGKsAglEIVb8Xw+7tCz6
Gg7ULN00Pui7kDHmvUhVY/3I/jC+zBaT2iG2Ya8jcFm9mJgAP5QEnCcWcVQq+uCKdcFCcijIP2qJ
Csvu3xel/+hX/tBUXkRI00YWSyaCimbCfZH/mbTBcTvyyOHlbduZKDV+8IioGxcwCCxeK6idEC4Y
ytl8Lp7STQYc00ciqqzhFzHvmB0DZdifasbCMaQGe1MQODer5lN0GnhSGNowg+KTQ55rUL73NtiX
dAlGedGrHffgOy8chpOFRyP1arZ4cH3OFfgxYHt2Cx2et/Q8QDlft0gy4ZnwB99P/u68/bo8gsYh
kHEb1cACWmHW1rdpErqsWnAsP0Ad0hpfpUdPKpcs0c9QYRDWLwFxzUZwfrjCMzCjZsfmKwoB3zKr
Yq1QMQ15b5MLCaf6J/+p6izJxiy2o8IpP91vWjy/TX8w7Qlds2Ln9hh62uLGtX8jWqtbS93BrT27
wwKAX2zrL1ZO6pFuzARt9up+SbLYuC0RO/EpTvyKIvmAeexgxQtgsfA8CVzch7hK+RiVrBW0UR7V
H8JuBgSLdfGwvFXTxFkniY6wFla7ASDQOQovzqNaXZgqWIg4XeckbaAjX0B6g1Daifc101BNk09p
TeHA/YbUOenuZ6yjpCxolDmeChu5HO55xIHpqBz60VfPpqMBjw3LCSQJv/hzDQcmdNOHZgBKsC7n
R1BbsXIJlP3Tnj6rCgtvFRpqAqRVcNqZUY33UbT5Ssn5aXTDUmEECPIdc3P4w+bTWEwPMrhlPN2m
LPaFHRJo7Ad3sO0MDHDWTl8kYEhDwAemAVjBWn88MClTn5fgz2PAy1ZbRyBkgBepBn8VqXmr3n/e
NLYkr/HNjmu6rJ9Ow/Pw5cl+FETRgHpmvTX9vEJy647dUgC9DpuGi3VvLTC4/tCT0yXx4gkmhWoF
45cA4ZcRh1fxcwm3+RmOQ1sc/HRoAUK/jd6IwMTYyxGXktJ8GQNaGNSqW8s1Ek2FxsxsJojXx7J3
VCiw6qukF7A0rLo25HVrOgKd8e2+gw40/YQEgNaIAHdmFRrdRkpbYdr/Srz/vi80fAWFoQaMY5N1
HEjbY81LohHpjACa56PPI/E9SwrZSC67FnvJMPt5DTgOgwDMF55bVIRq0lgthVfA1nPV0amRxP+w
WGwiZcX/aRXcI9v88nWkdv41nbpN4cT+CmpekBKkmnyjkEu7w3aozL0baDT3Yrki1x6IO5+DFz01
MTO7WeT6njRBtKcYfQ0L9UUBQd4UHajELZWeT4u6WZlQitPfn7Yi8cV3thIwZifwRu2GOJaPpj43
C6lmT/eV0/4cqUvSWPqsepgwL48lDLgasDzDInI560fJxx7IMYoy5UH0MhJYRWA885nlkoOOEToM
DsbxzY5p4r40htiS4qqwgiplvU0NRb8WISa9UB76BhCCGS6ZdLNLnWm3UqUsXi14hr6J60ScELgf
WOSL+5+2UBYuo0xqUEbH0XqoKH+wiG2cBBFOSEjwgVQ+VRKeI5IldwKK/PST+TECqEYGPWGocsQ9
Fmz/PG2W8tneY6w2etpCNEsj458GPZZDEUOd9Is8QekejSfVlG+H5zptql73dNU+xs81hjHtWc+k
CAQbHSgsGKm59sPxMm/8huNHaEnbGZvspHj9sJirfDu8cNl3ODfVOhvJ0WOcoQS2ICXhAyNwzCw1
1cA09QoerEKea422LgKwAnUWfIAPnFNwfLn2LFKsHboClj+RWuFn2q2dIl5ZknSMTXSCYrl38L/F
MVqX3fb6fACN2Ep0+lp91DlME59zGkavfBAZntqIVq5ickMPo9KevsncCvRrjB0qESxHMk+Zs+D/
vDb76tDvH7KVEJvzrhTwlzxNPsBChm3Bck+TLXUwz2T9mfUI3w6nnUI3eQsn8u+nFDoe6y/4NqOn
c7+OtE5AzvZ0OmH9Hh/TEV1lY+L3NRo5qR0jaMvUqLWRPHW/VMHr1idivEDIbajR4ZUcYb90kCZr
5vpUEuWwBf1BmmIKEDF7arm0knQJ0adJHL76D6l51C2QH16hQ7aOuXjN5AnMnsRTW8C+h5A+kAtq
psRM5ppi3b7KNXDjpwM3LAAkDENjLVnS8xDWWAZywEEIWJtJ0/V9lwe+gQG0xBAS10eQzT4KLoSW
3ioQcTy5/4+NCLm8biUB16G+b55Ta3+m+nGK3JkkUtl8FeRWusY2dq76r/fwKDuHYfbTmmwn6O/l
h9tuYMi3Xejbjqn3bQW8vIAWTAPfZgRSMJFKZHstiK34R/S4TkGCB4KgiloNvxP4RSrV6tL7M3qN
QoLqHY+izg+7s/BGzmHujU9Zod8LgVVqQ51U2Z6AXKM+J0EO34RyHQjWdjapJCg9AUF9ER82Ufum
9Kg7lvi1BrfL1Go2SgEyKVwh7aQcQKKlaVP/AE94DYmHtl7ldeGpqlU9vBVDVBbSMz2yDYTqzaYL
Ohw/VctC5WDG2WLHuOFdyXsqkKZiMOX+ulGzBz586a5nk8+tLOYyAhdkNtGz5OtoURw3WIETjAYF
wxYY/rXwayXTmE8dsBK6UNdq2D2JDUw5xswMLFA/AOekUCiyXMIJmI/GLsNdejwYLaotBhOWV+Ne
91QhkxCbLbQCIVETSCIkeobVB+rT0LiS/IBwHQMYoOXVFHVCIHB3ckHo08uHCDMmZ039jglmsqM5
q81wA6Kpnyn1Eyt3rvyM6ZD8PCGn/ihechK5Kn89x4RD5Ay+iRFid5uVshP3e1IP+iPujRw3Hp2I
tHbmpUwY4lq9wsIkgRJliwZmELm04wFa1shZqlpNNkN09xkQlEa/apxLJ4bt3BjudsJ/dHB49U9/
8tQE+Jr0dPHvv6H1lUL1wpBkOM6G3DPgRK2Mo9Xk9JR2vpEUraT6VxwvO8sFnWYu5JrkH+VwyXBQ
FMupTW/4iop/05ohJ6eBWMZAlRKNrDfacIhScJ+gEdp6d5Cw6BABrEzOgp+MhJEdIUUF/+e40KK3
rg+ztze0UlQZOOrMvgYZjg2erNT8TnYRRqttLDx90E8qBK/nepgTmiu8xVPIc/INW069jCJGie3f
Awv1F+b1kUpFBQqPBUy70TcN00OHWFEMUNelTqDOqVgjkrFdll31wDr5HEoLZMuB5OW42uau5EZW
x+QHKtGMD9csxjMGCDHIKdqF8rGFng8fFRR6c7hdrMe8J6QFppM8Sd+fh/gUJk7z0tG5Uu8msM7h
9ZY1KXv73xC/HxugoUmT45oACi9RmS8mcoVckMSmw/4mZmaWeYcXbHlONXvyKMqvcA2GrMOKN9BQ
q7SgxoZQ8AUjXXHaArwsc5ibmx3RhGEyOBtecqksr16yancHlVwftVySXawdwhP+4QY8pOdODp3K
U/AxnWiI4QG4LkTm9ciWUGDCCuxh1/CQAlC35RZBzmh6j2GmjGgC2nLy20MqnrFvCFRwAeEbgr2A
EPPAon0wumr3S8IvBSxvtHDJSdDro+3F80hiA8tOtYYHWpejCAFUKgEZw0fimFv7aoCGb4OfuLGZ
cAz1nbHU3NLM4upOBXmpuknuYGRE7uDzKP3W3VYSsGnyDov1FasUdcbBvZHj58I5G+obqz/MLLyq
iAT1TYEy40cBcFr5scAB/1Vir0G6WR7VJJwEIYo0/g9gZcW36UDUlLlmNWFt4z8eSkkqL9Hb7ODQ
3V4MV6paHOFKCskKsY1yG4HVc/tGhIgcZyia2OI8y9N3lxBPO7IGxq6VAtZDLbybO4+YZt1xC5dW
8DDyF+wUCvL0ejEkRtHEFZJjz/AooX8/Lu1JPqBr2gOH0t7E6TkPabwhpIBgdQKJAOiEmn8cX4PR
DukEvLXUfHHK6MAREHPnarsAXsptio/xqOc5IiU6sb5R4tllGgg9gxvRidbX/aWwNygHRtt81nHO
JpeT8WuYWFDz8DrQL5+4wKZYcpw9ec8Dfzw2jQEvBJGiJ/8wItD0vVnITqcCsmVlPYwGTTvooqaJ
IuIC/pV01zgnsY7oLmoQtynMP9FvECuG3RvhTo6HEI815Ls0NMXFS4mFh2nhmsyE84Dw7ab8Ohfl
miYBUB2HxyIw/Opup4afaKH1Kz7n51mx1ThDO9y93isQfFXxyeULfiMG2GmP+2auBvgOH8F3SCyN
+9HVPZmFey0vrMoN+DqRNnLFv/PbUCiT92rSwS0mHNqk/7chTJv1KTfUV0kfY7p015HPNZi0lAq2
cimVfW3ABmPJwXDVJWLsc5S8kj2xP5jKWfZpMiUMvVl/HNr6QfDnl6l8Q9uZJg0bsTJ6IbQjD/PI
xwfYeJuYbuhSJlu5bG40NyhlujT2jkNuYxMbnkkTDRideT+T3e7tCtS/MJBrOrSPww4FvOF+bdTY
ROE18gXyBziNYGH7Gv4+nWoU4ipbf+PVqvxaN718nCrBa/5XhGDW/Ox8Y3F1S0JAcJB0LRozJrAo
h9g3ABtvNm5Wbom7T6q8uY6X0jWtDjF6SQKsCIB75lUBHykMQzPKI1zGn7gkSbNetSiY+2Khz3HX
3ZSpstGuSs1oMmKfjNdBk8t69FHuhE7a8fCuJ+IECjRLWl4ODTFGLyuCK43oT3X8yFGp5FaL6K+Z
5LdN6Mbyl76XwoyODxttxdrN0qAip9rBkKKymbu8HbRSoSGqmllyFxrTQDpKo4/6Jqb2BQZzjlDG
z69NnPQtkGiY3BoSNsuKgk6ypvSVAlgq0GMEpj+qbKeWSNgUeddcOQugj4jxk5Ju05o2C7wdOMoX
hH45+2i4wG6Dn2Mlj7SA2gW0lQyeFJ/dAuxbalb0hQ4wZsxmfYUVML7uaZEx/etSXOIPhQF4uX3s
d3sOLIYaiiVC4wWgu6OqOtvnVGBedpLqwqxsnLx0IMqf37wgl2fs2ihY58hfFS0shduoh45D0DMX
fOkeU7CbybkhPhAyZzKZPvza8M0W9w9ofevKF8NlStdy0MdJS1f69ZbYPI88uMEtsZ+pt2QbtRhp
bGbr2srTxaeP/VXTBbIvnRwp6sipjKqQ+5gJeSlOkaZH1sBj5Jkc+7ICftRfj6lw+olhM1Qd9vC9
YSp8lCLCFlm11LMjzYNO05SYpnvkZPAVPWPiwP1zDX1o17IUJDKZbdVEZvWXes+tvLfqFVWGYFa0
0beq6aoLB/Wg9Jd5JMvFHKH/IjkhkIC4Xk4ZL0wZcuNe0VHz08VFHNa9sF9gq55srcH0r/FZu9Y3
yVNMssN2RX3NwA1vooQTEuTuFw8vCa0eNSiJYC39E5tgBgZHeyXzZX9UI0eXqv2nFnRxhKKiYI9q
DEVPtie4xi8v2kipwL3q6IVXYJaACmM1qkGsXoqu6Wblu2WqlY5HnbZyyLBQsEY7x8teSrVHP0Mx
vXL3x3AHMxo2Wj2rQL2wK/IlMVG8w4Y50F1pWvbsLvzJVHyX969TJI0T+xMLMxp9H1HgIuDcSBsy
cRSRfku5N6wUibdKfPtJWUc4rIu+uNeB6j9pvEAoVb//XBaI7JTojSkeLL7BZ3ZE9zS1O6pMPrK6
MI3AnJJ8gA9UxCVB7kWsD6uPUn6WsZnEqH8Qy+XFilxLoVu9TmV3u7vYXZQuAHmvPH+0muLrKYqV
6ODv2YB/wEZcpCZsI1mWPkv9Mv4lOMtNdUk+dnEijkt8y5zVdhEM2Sz0KQ0ffKOimKc35G7A8WqI
9EDuFBB0GINpO5DWX6jC8AjaMqzL+3WLxML/AEFqCGhdkrfFkRpXvWM28am6c/fQ62vlJWSs5Egw
2yYpU0i+EmkWuy6BNPHvE2MzgLH4dxNbNjZO2g+G409W28ia5qqrnd9VZVcTpZpBT0/YLE+POf9F
zgN+F3yH2RlrvWvQwB9sUSEeot7Tqwo0RhURI38euyr5Z7n0xQ6g7v2YjkORF1CnIneXz23t2RH5
EeHW9HWYOVbqm5I2HP0xTG2iB0RFOf5UX+FpfxRXdox2P8iRoABaF88NBDNG1RuyQ0ah1GibH24F
s4YdWycXlbDzRIrHONOAGO5krZSca6zZAbydiL1Np2McHki55ceK124Ggab+DBLaUyuLWFeBg308
9tzmUX1HAaskelmqzcxtjMlhs9chdOlh1wPxWeTl4kS64kn0Qv0BGmFpYnsqEZe4LocVuPKgNkKO
u3bP91Z9bBV6uWp3udpX1w4ZQUAZ9e3vQHIWaxsOo4n70PN2MULH19BtLsrVWdxgdK5R1zV95U7q
37cP/NjtoYrrM87VR4gfYAC08Xrc7lRDTbM4sDFumtWfi8b5TabTy3C1Z5WTUXU2q9lawf0eeOJt
Dj9lZrCOOD4rlnu7Ps48nL6Ex6ownbKhqFizN2WHpHTAdb7zqamgSaIwnU7uzgcFlqtsFr9a7unR
vqq64N4AWxX30/r7erg/SrH7sKd66VGLgbu2bkuCxb2CS+3hoU7L6hhxf/2TNgaqxU8j9Z3HJtmX
myZcppXkshpyltAXebxY7zmrA03TNlQ2gBAgzydMPp9lYkN5FC8EcAhqogK7gV+xw16kCM/PY9eN
a3l3Ua3aHBhSqG5zPfWNtKybdjnclR5IA44jqLeh5ImZchTunMcSxXhdQYBm60dYEszgEOa99jTw
uP4puLyOXkh1781pWksC26OSN6tk1nkAlceJaADHT5FaOYfSL0Fyt0F1swk0+QlugMGdKE4lEzuN
tGHvyVX/2PQP7o30pqFRRgH/uN/KWX0TSUP2aJ6oHQlXnZe05oHlJ/ukozwCEAdLhSxSK9MwYAX0
aQv95s7AJzHOAbgqOhb6SVKhINkL54zI6s/lqY5faKigdomzq4VfFV1Jjxe0V0LY+E70TOCbgeXG
Y3/QYLxn20tO5bHzwQeGTA1jrTDwFOdGZMf5IzBfB8UQRhiNCHsI4Kp+9QNeA5mnmfREZYJCqSM2
sH25PURo95todvluc7qmlFLPrBM+/aUIS0raBdmmO1GPhTyMmefWXqTLPi1r7/4eFVetbxjwXQJn
UDc32DaaiYO4Y+PxTPb2nqxH45Fjjhl2oiylJ1y5Y1IkOxE5ur4sDVvI8CQHjbzl8KFuR9/z9Rvf
n7Y0x0PvCj4BiKFYidwqTfjdMtr9Ue3elABHm+ED9FYahi+h8qbzXJm2XvWlvCrIUzKh4TPn2kPp
drQ9YPxMC3BAK4h5OTsyOD0LkrU6gfw50EH67RQyS8cLRZkHph8hRBENuGCe6oLcv8YXYrMHgriv
tFU1cElKPQ1t5FLy2f30yqra+Z6dyWumnXo+6ituh9NPM5NzOAKbXRVAElwrSa43GUs1QCj5+0D2
yazcK3JbSTDXsCplP/25iYgBFd4xwl5k3sRUcEnMAAXWSvBTm3/Sc8jEB6OR9YhvJneJXWUdv+Xj
w0mprXw++BqM0M1dmzNFhSZA/EOGbTyyn2KQLhoqH0iPKA5keDx8xvOukiUPQyRn1D/iHbqEqqmD
NEkc2eciVp8yBY68UWsxlU8/WXWbIuIDpzFLHT7+358ksezu7SEhHPrpP1OLN3Q/ulgeRwEhGpN7
zjvXAwQ3wjymrX0nNDAPsiCH0hAeECINxnO8s/VcKROUoWqAUgW/R5RyqFAhT7zWwIojCA1iswQI
uwKedbA7OSTSqLRAw2kBvMXj+7oabSNN9SadssoEK24gim5QEHMB91DyAmLFjwkU4xmYEm8teif0
AM6CGkv+BDbUgRC01Q0UfB3ogt5gU01bjDPmJdSNyKKQORrASm+xvlBDPPSx/QxDSGUJu9k3Rw21
7U5bi1wsoI0AItasgQPMxnVN0tx9RhVw53ngYe1VoTm2k0HNaICNbwKuD2+aqMnhXc9r73H6oaYa
UO/qViNN5DabpaRaB41lYirkmgkmmc/Vzels7kCtAxj+evAFIi3aw8BehVL4rSulOFjJipa2941s
YUYdXvvpSdBqsVmV95fGDhLLPPVkAcCg5IXx6nopELodh6IwAzqhGfRE1XAMg9v94WTZxNuJcVXN
f6+XVlRdNWtrzI82tIFPbErLc61R9lsGshAAEOD+7xnLJq3ffPYF/gYfSPKyCcmL4YVfCuvxiBC0
fbCyoN3Rp9u4W5VccT2UqmhWQMcqAkOUAMFJsR00y2ITG8p7H7IGEBs3XIf7bRmxt5jvPehjRDD+
aIzrap/p+jEZ1M9AAYKsXKFQ8fgJXAZf3AuIZpIs16JJnbXglVEH35L3GV3EOqUXDj/3I+l+L8R0
6lZv4beWlpTreIjYllfHi3koWX8j0nHQ46fGfTya8cl+Cs9rwbh+ilAtJo8c3XnMzAvopU9PVYn3
58MG3wCdsz/Q5R8Yye03jWh2fD5BJI3Y8jxeSQto0jMK0E7keoMcAHG903rSaeTJ+QArr75SGCpP
zDJm6+nzho59AaYB59f4YHOfFifQAbsfFl7V57swq9mE3uJmgEreY87Ba1jWyl6tjHszC+cLVrA6
p5Ct+lCnOKIMbDTKl4adXGsBFNCp3ZHhVmDkfJdH4yG8Q0h9j4FPOc5xqkamRz0f0Uavsr77e3jW
dErg+frrMhLQlkj9Hl4p5lL6xLsfihJdTC/2Io+dmP5vlDW3PkKsWFcB3T2JvyjOi0utyOv5asKo
SIVcJ9HcCxNBmJS/YlSJjchthglstGhdeYSLTe+MRyeiU6RjGk5w9KeC95mDAwzyO7LVxmYRvoe/
ckNPXetunrSa+aNuAveu40OLuT85y83tnFAdLedU/KhrPPmF03toXISJdzkush7kBZoYUIQYl4TS
lMwpvlxCIlf/0uQRfbrtzq7HHvWxT2jjIvMcnechjSni7RYRlKcVR1KOICTJq/YSPsme2o34U28m
ACsrCygvKNBWf8/UMkkkBYfF8T1ZT1i/Qf05/GyEOVIxvKLCGtdKcX2g2ocwzOSR9FuKe28zNnT8
tbvPXjYinM8iL0vL/WgCoPT8N9fBSgwnnDscrZrzkXfWpIUFd6HjpMzL0FD2A3cscn8LjWJ12Kez
lMRNSkRoWNm+30JGSo3qa66z+QZUX8U+2wlCgdEwhWYWw1cV5oPu9wutVVvw1TU+4bUOZJsab/uU
NZPOCJcUmm1XfsqV/dsVcDDQZ2JPSdhcEwhEb6lJWDEkev3KPf/OIAEAhLtLDBywU5ktc8/koFg1
JtfmEV7w4A3qXKhNWOBBfMXJrevxMOXaMPbSikTA756ID/RF79uK6wUzjD6aA5RrwMgdy6c9N2/2
jRrZAMwcAEScgcb0KNaBXjSwPfv2DMDm8h1vzFuBzcsA7J7tPWWz9I9sR4b52CvOA2mMiDATTR33
eBEFomKaC4+LB0R6o2oeO6zImwndBMCBiy7j/IzXM4PCy3NVmh3reN30BNcvMSEtuoy5QFer5WCU
tGAcPWbL7IqBEzneYbtjigTsYO6rgGUINUGQfDolSz0JW/IRKOicekdJ5d6rYK6av/7XWO/wu39W
JjDi1bbkzzViHu2iGBM64Cis7QlACmXj0G80ZugGnbQtY2Ikj6JghTloquRynT0DGjaAziDt0Vcn
DAtKewZ2o31vcNTedbTy+MQ7NRTtgV3n6b5rrSIDa0g6+YRxatzreGRIPRxbfzz3M6MMl5rUd/o8
Ts7aHQoYnFHg4say0BzFLXLnau508xHN8U4cSlo2HbDej1cDxjCc3064KnMsN7xKxn7Ka5eviru8
XBVrvuodcKHSKzAAuhNid0mIVnI94D2pHnotkN0Tv1J8DqLbvoDU2zWSjoJxoRvwxu/W13+NW+in
B8z2+FiKQmW0dQA9EFon03pVwN/JuVsKr7xpevVgnOIfbP2FjZ2s1fmvRDNCqFi0ux5msTksepak
YXxfD6QP7LoFSVPnQmZoNCrR5QvRRE5SO08FFan53rjz8Qu9J3XoAHY4oks9zuBaYoYLakJuR9bc
LbEXj2HFsUCMYcefYWYtp9dSumLLILzqw34HekYCoCFPGJwgiUEh85Gpn9h/Xgg67SXTDvDNooeF
o6MWW2KjdLWqfq2Y16TYDx5kxr9ylD+1bvAh4GMZt0KywXNVmyBRWZCSd69kIlVzLO71h7l0kqcT
oPVy7dd4SJWpeaDa5KdMeZzhX8aabZWE4kIL8v4bpOzsuE0skCKDri4Cae+YY3TaJKIEME6y+bei
yTLY7ASOuvukfgAhPCsjcOMmdYmu+brw58/i/HU2VXwglvrZitvPmt6+I2uB7fxkypMcuwRzYKsH
fEpYNGbUBMpa7+WMjLyHGpJl/K/yv9e6/tp5ocLjzTGpzD86gyAu/ovZechjZhESpEuH7yyjtDmH
ox0ZlULvUMjJRc3JwWNx5Xp//hkA79GlNCBjQRzOFv6KnRGas4bu+F8nHDwThXJ3sCt4VZeh9SKq
4zOxnJDjRPkCRNQQUbGmBWy4A9H5XnNV/57CDhoehBl5Mn+vqGimXdS3n9bx1uQufubhBBXuxFfa
ZLBbATVh/S0t2MiEu3ncImbzYLhf8BMkbzaSGBJvVYk1UdxotH7ZAYfxT1kl2qM1FNSzXQ5ZQTrI
AEhDq87MPc04vN77XQ4Le08pnqePUO3ddDowoVMofJpe7YEmDjW1JPN/Vv0FwWS9rqp/KCKGrlne
zWWkTujtcrdSAEft8OkvoY/0t1iWxtFSoVRfnNzv1Ho9+eQrOEdEQHPG16WAOMPvngXbAFS4dpk1
oFlUpdoqI59+pyuXUjeGQd4K3JetUGXNOzHLBg4FQUMXKoRefA8txiFbZ7hj/Ng614fEeDobPdR6
55vmOuDeld/EgsHe9wJ73ntiDrMgodPKKoFgoJ74u6OaWypFjCGt2RmyYLzQAXCoTiJC98hlElPV
o548aMTOQbqYsVdq460KrW3MNg7Yek9qEV6gASpx4CJx4iZZMzxxX4AGS/5t1vsnN6gzuwkzeez1
Yj4Emp27KCrnPCnuT2EY9zxM05bqk+d58V16I42kZG+n6+aOAMxxlzi5txsjByw5CPgUuV52+L0x
ktzj75vpPwCIFTleKouGIgJjhuGmplDoSJfTzBgrhXiq6HMszrYJFhs48gtk7MoXy+1E2WtXyTpH
gN/A+PEcuQKXmVrVw/IlT/JFPpEounpON0l1BreIjEIXc5Z8JGisVfcVjDcVBtpFmXLemjX2txix
i4rhUvi+wvHLDmQ05X6qo1Iy/b5ReoCPTXF2PZvRzU98frXXRfatBc9iTUqM75YYHqqU0WLoyTbQ
17IElOFIVy4snbxPM9u7PExtXPtD3+O/Kz53cSx3ID+Rz4qDSoqqmTON6fzJFSb98XKpPlC+0KZ6
ORLBiYt3XcSEltC3wPBKC1Towxz7PDE6+TU2sU58XSi+/w+g5BN5mzjokf1BUE13QC8z5aTYth/T
G6ur+c3YEo0oKuHdUHbkJdlNCIv8mklkrdgtVIR6w03wx7upjf7vQ2JMV3/gh2iWoy2usRqi4oTj
3SulohU7DTQkMTdM6wCU8cS2bQNUabdszp2jtrkqDfNMPsdoKYd+eaDYu1l1DdpeaMP6ULFTzf/l
gnBJeDWD9b6VPSylujfOX1/pNdaJildaJpDGFNGLU1/32meQvot1H4p8BqveBOcVQ4ta3Y49w7Le
klUJaae4vH2OmFvkltEpFwZ2hONcKjLlNcmY0eyUZV8pvkBvCDbvNlnGd5xECoXTajRslfosIabT
oOxOoK1M820ENIb3GJRnxZXfFfthrx2Vf10CKZALfURuqkv+gHu2xyfY9aevmmtVfIbHsuX0n5BS
DcniNph/gVbHP4M67OtuhoBn2WvA9pLrmBcDLOTSzUcZSViqIVi8FE+zvcjZsqlERK7WtywBpN5b
sAn+ojuQi9uFou2QCGRDco5RA+JIT1sNlLkDNyppTGMUF0uAQIbyteWVd19UWSlnwhbiEURLjFEC
xf8bahMms6m/JE5evBYfCqT7CNv2U9APpiJnH/gQ3WNIjRlat1tjXYGhcjmEVX8mcoCbJV1GTe7R
1r9yzWcsASnh83vdGKjSuIJYioaahbvtkj3d7DSeCU1dfe7iGRRCQvjLnFbeKfjsEBfZ135sdRi2
aSmkAz3wbc5dvsBAVzbH81T5ZxH42nEPwkLw0L0dn9eXFQl/dKi3P+VmJN/AjOJhZNlrQzVdvquq
pXxpecIkRMaC11HjJ2qeWc4SwviSetG7fj7dUci8nR8h9iAa9vqxyGsBcHNvbsB4tJpRD/libtKi
l9aKALVIo8bVhs4EC39Kv4ceN9KPRutT4gfGzsopm0GXLdR5WBr8reOvZBF1pk170NL7L2NMRKiR
2pzFNbchStG1vQFDYJBPRuQjZitnszk8oBsAvUJwaunt7SO6l9nSW96BTnt7nnyw21p9PPXzSa5w
/aemVIJCCi4VrbnEErfyMnCiQBw3p6V/tFOXoMyJt1yjzKT1/NLh4PEeKmCtsjgZBh4XTcqwSenO
nfUVyRViALhN3PSLqP7giZQfMBg0By90lnYizfbfLMNVyUFQwXdMXL+e6SCfe5kwqdIr0w3CFXLb
VUdvWZya6W8AhOFYDB2QkEKmGIxWpi5SCE4zeywD0amcXzgUmgX6u2AHy3MnmwKaQYta/aIp2r48
N06ZK3O3ANpJrx4eHY5ro9hUXP3XOUFwAYI1SUCEaMxPFbNLFpAhwqTr1mqUvx7xBuQRct/BSD4J
uZmo57z4BOgKV8gLYyg4AHqqERGqr3vEhHc/UyDd0NgovBLv5F5+KUa5a0KWPWcDdxwWt8tcYr1t
2+tUrO1GiBOpjWIBaSnoaYvx05ExBFtp5NGpFduSF9HCd6GNl0DTE4xfIjhMc7dDptCsZFfZjbQb
FS7WZix4WKBn41CpWL/bg1bPigyalxY2739kouBH8/7eAmffb5hPY78UBKHROX5jUL8v0sO2fXL/
47tdBkMaLjvWPQryURrBg9l7dI9ORVn/JO8tgm1q6VWlwIZMB42MoTyRycArOpZbO//t83MCf7Ul
S3a/QHQG/o4/6sONYX0bc10ZbMzQWpR4rsm3H/qloQRaKofxMokMSE/boRxhOwJcjkfuasKTuzUv
gellivDiSp0tkZGeNfBQGMV7SrZolVM8bwIzt1gjzjf4+v6tj9d07hVBiSG0xhLQ6UWof1p06y8c
ZCfVQQaBPzVv0UxKylDii3SvD4TUdY7CLt2aq1jyMQ132cIEYy8jO7icSbKLv8IesCPh0wPdY7s5
UfWc7/rs7E5KUgLcFQ8XCKn+Bw9aI+lUVB1Xm4e7SBUsOstmsaA1LqpSJ1BQh06Mv7+9Orhi3jN+
rbjR5Z6I1CHDt0rCsA608SRR1ZAf4aRoQB932CiluM8rET4+LVZuQf33RMbuyrC13Vlxfli0qzFG
bPP2LlKBYQ/ssYdXiOldttKgd2Lif7pdvv0KT3g8JkaGZhQs8+NSIT4zPgpi2einJCgJ2M/cDbUT
Mjf6Ly5vwdgdvlavbMa5Feqvq/J1cxzxmrg7yD3OthaWoVD1LzewnRz9z/Wp+/3vyNM0uHnLICcI
QzTYThC55KxpicaJZsoxeTBFL+eS97pintLIQQL6n7GyvSXHHNUKQCvGZsPeoIGpcaFzQf65nzWt
cW84uTiHDpPsDBReBwxrWyqNf8pxbopVDFcAPDOvRv5gD49LQ+mfPsA3q+HfMllOgA8gugGygvMr
eVqpgEYBkGfuTAMXyVH1i0mVGEID61ltikpWb3zNBqUsVXdW6JNJlApo8riB+NDrm2wk0pGnFBad
BYF+Ds9Da9Pcle4YeiLUYDePl6xR2In9pM+6Vcr3OwtshaMWmwxUHcapqjGSJ52amI1RNJ8H+dej
aAzBS74/yv5A5SJBMNMR/FMbuqJKpbKZj/Q1LmE0qIMVkX7pINFuJgm4XP51SFgDFkztTiKgSRj8
nCCacqdDCLEiVYFWoGrAUHj33XwjccuIOLO5vbQRgvyYn9ksv8l5wm4wcMAwJYHisWGFyiFMDR5K
80s8fkeZzBjOPQBlEGYcXujC2Xh3rIIbQBE1OLGU/I0YdlTobk3gTiji//mB5pmicRBXReYgcT44
/cGbUwAz99vcJ9UhX8camUqky6b+gbzAlloUSLatHpLumxaXk/f3iZ+mulYd0o/zXRtIQ5o8xPCM
lWLt95vpWidJWKNotVf9fOhNhJLi5jp0P8sEtVog8cSk4L+hriIDY0dfZyRU+nA9iDOzAXh7je8b
BHOsqhcfBb8jJFaltrNxDwrHhBIir/QCQsYdB4mPho+7PTTHQey5xezttdQ3/dThW2excdcPbFXw
6wi9rUiBH9t/lzQOMaUMyMcL+C5XXeD+R8+jMZVMkZEXQZZSdgz+68FUmUCal3uiWKdbnq8LLVDM
C2jk5bDcTtpuDrDyazuvhLd1nEtJGJTIOGevE1uf5k54qldneYvM9L5Cppgb4hO5MksM/7ORzbPR
OLd/2EPMm2CPdf/G99ZmGojcvKwiimCNefHLdbRGi/3ytmzLx0juIe0jXLDctCj+M5arGuVZJSWP
f5+X0tql2aEROTK9r6Rd6fuXiXPeeHjDwFAuXICIK03k7DIVfZpx+A3P2XmiMDZu2lHaxbUgErj9
6yKM/ap+KHKjzcnugbo+4H39qqYYBOyI3hnfVZ0QwmaH+b42BthNG0iHHrPDy45d2hs191E9hTg0
pVCh2SAD/VXpj7EIa/uAS6yUl/TIJpkKJGiPFYPp+NZdz+oiR4Q2QSuidsyrb4fdcR9ui047ZfWi
xkBPcqPWU9lKylHKKholDgjLzdeBBBmFnN5RuWul97GK//k+PBX+HdPO6kkWzF8hIlLzrd9UmDAg
BE7XjBBdIIhU5u8ntd5d4D0N5LxqqWjgIBrhhZlIfEPP1OhOWa9GMbC3hU0Khy1Tuc0wshYCDflx
8tQbwQoWfX1po5x2uqgdAUIP5L3QeF1IW595FDbHaj18hVxOPLb85Y7jkcf6hoKicGx4CCtfOC4D
xXouJlmdUc1qzWkCmTW7n65TgjInZfCRxIhbPsFgewNecFPtX4Vq1eD8Pv33klNjI3jcKav0fNbv
MUcbOkr6elediqM9TdFnVGatygr3VxAU9tWlWE/ITe+cO4AKLHYEEo2nzlx1r6jX63P7wIOKbPaH
6RRNzrKWsh2eiIsWHbq6Rp4AhjYouZOv7I6Lxhd4zgYOEaj/2+qQx7OPtdousS7GRFXrNKHbZ0hm
0LPh+ou8rv0li2VdOaMewunGt2+bJzxQOnzyDAh6ftT83oEl6T1SrRz//JCeLGL4j/ZNkXO6FPcO
1wW2u6xtTuXe+8LkdO2FW659snziJd/EsBkYVWsEFbs8XM8QBQzNlKA+CMck0fZ5ZOJh+eRNkNn2
cbhWQk9CzYfdgrfEm/POV64IFEigMtVuL9cl6V+0E1BJ22JAr26ThnPVVA3n6W2u7rW6OsEEjWG+
rmxC7yuRehavnI9ZyWBn9UwT629ys3cIhb2eB6e6AIeORaJSNdZY/5SwXz7Azq07E7wB3zr6G9nh
IuxMQX0Gbs9oMlWUGB22sXg92iNxBPAgx2Jf3kisbruEjKi0k5M0AL4k0Cer9OcktcJ6vBfSjPhP
xvl7um9EAZ+GgpY484PfbYQVN/o1YRMEz1IQtJQxTBkkMQ35PEt/6ZsEtdNh+mYeN8Yy4uvm/d04
e/qC6x6R8sV5/EsNJfK/iNjprPjJbRh3D+EXja1SyDD/5gquVumw96mSoXkqzJmrEazpzgEO4O3i
xJpbGKa5cTWbN1npET4p0sYt2SAqi7sS8MdRKaoOqEDxloq4ohDkOmnzgB+PDJ0EAFq+JHxpkH7p
dUiy1eWS08SXuubnqSx5lrXPxtswIVF7a21y+ODNIhUsUkKf+Dk3EU6b/M/oVNmNa4BpECiOeMI1
b507mUmma7BW+TZgiGmrtVXRgIxKq4VR9b/8z5sfMKMNcs/zXN+YpanYEDfxTN/HNrftzDNDOXKV
kbUsEgz3synX8fvec9ILhPYlsnuz2ScTcC5EMwcCDz5EdJN5KKIfa/gTPCoXx4aMMn3Mcn/qtDlC
V/9445S7g+eNqbZZymydXd4f2S3vn/i0lOruYg/ViRafpQQDPO+An75NDa2Kq1lAwofLjqXiKaDo
VNFV72AOUuG+E1bsTtyN+zAcs/p9QLJG/9JdiGocBqLVaaFSPCZ7DUkebYfVuVPNFw6T4lFbbdgL
xDK/eqC/+ujSugPwoe3KCd+T0XQGB70z69jP2qrstXBwexMxTJBg2MablOQxivBxwOGmeowWDwFs
snXx+96Q+633TJuutmobg32bEpUbUrsO3H80KL/yrOWV0R+x1GNAEg4ayM71Cfee7CMBSqqtMrOH
c13a7FbQUewSFC03CximjwuidzcSdNdhLucO4ZjjFQ3bDkikw2BgyOKdlHp9JebtDdxOpxVaU1rm
w5eaP4LLB/H2sw0UyY+Goa/pz6JmF9D8bWtrP9V/abqkUA/1UOZ3fCb+i7VhUoiv85j8EugqBBno
ZemFHxlNH+igFisU0BVsrem1TiiKrrBCS1HpK3Kq7Q0MD+S+zh6GBLczyCspVHi0aUzNJEzmnUFv
NhR+AqWG9T87uFyYAdjYVl0jd+Pr9DJi0sgtckbyoQfy3Q+PeEcHZdRl0+Qf5NrX2wPeBRRHFmbo
fTOEG8XF3L1TOXqsKAx92QoNFgPG0TTyMAL/qKTibJAtpNdmnwE7KYjPWNSMyICfVnSDpv9aoBtt
HL7YNhvlTt7y0lgHflSlmRKCsz+t/j/Yszkk33xI2Fbzeczj8vUMeigpPFVeJ4SNQ/feMq2ycpsK
Dsp5NtCkaUDDT6Mqrj2ekK1YaL7F86Z7YiqEBVrjxN7LuMi1o2ViNHaJWxU73tOP2aajjQP0cP6X
oulfYA/XZ4g6pb15v81OYJkDqjd1rlNM1WJQ50YZBLlnGxdFqbpuwnT+oxg5osu7j5hEgyy+L/Wf
NtubACxWKazljlVEQvOa8YPG+uQT3uAa4MxmwQzmV7nH71HJEyIHUGGf2omBlxyhOcVyEez9WUMu
laZ26PvNJs1ljH+MNxpW+VpQqZ0jPb3zzaz8mzmt8l35Cm3tL04jsqpOVDaMwOAafoakLfLFq3mV
l9KqvFQUF1SVB2nTzFXcuABqrqa6am9P3JDPVOKOJbgZ90HQ6AF0pcpRs7cxsjjFKzMvsmhrNne7
eWUKjbMWqgV1YZCEY0pmt40fvbaJQ0Upv2+b3EkIVeioE94f8e9e7tBKYKP7DFmTiOJ83gZD9Z3U
GixqO9am9SBwctK6bzXOLPjSDCBi2CnC7QP4m6FHTO3xFDuXb7a/Kw0J9zUd2frfcWEW9/xRA/Fn
4Cma0G9x7IMHPb7gZQP/vBROS0YgrU6p8Zm2dIAPJMKWIl5tEZ7CMUgx07hHgpStjjGV2JC5+Kyu
oJBgfulq9EwFu6iMsdRhRd4raPFHK2fWocsG/DayLxdN9DogCwOwttWNDuZcJqCOxQWICxWnLdoA
siu3XVmJsZW3FfNHyPCsQIilVi/M16MdXwIirCtu+OyLL0j3UQbXyOetcr9K6cYHTUggyzb+of4N
4FzC7hbNDrjhqMzg6lk33P2mUuRVUgjdLsaZXxr3QMUiEje6fsq2LkioDbzvh4eatBbUOnCtNYoD
Y26zBmIhfRNtMlFB0Mp0Ve2OQL1tt2Q/Q81F/jl6gQxXKWIfXwZB19uUPEV8t2xwsqepY34fGuak
n8RLyoJAI+sL4N6Psx/HZLK7fDwr4PVAx8aG36mggeeWKJ5HxqZitWObWklNNr3YLFL23HEi/wQ8
sDwCJaQk25gdMYf9vBgEGYnz9zqDJ9uuT87Jq5xQgAXpUOf7l4PhR+sW5n0FJd9lkXvHjo9aBNtX
PDazjcf0VQoOZiFrdcFBzgwrQF0sp0X2fO1ghltcQQhrXUS6LKwvBFaUsHZcz+vo/+26su9rMIPi
Jj10MLyIiLGV5TCqkC+BuS0MMkz7jSP6UMLSkwmi56/sUul6Sg16tBsgtNBviYXwgD3cUF7hOQdn
vmwcWd8YDBmXpL47Qy41ho4kY2K+7BG3om0O3mzvcl2mLPWvbyNVgUR5qq4HbHcqHDEu6rghntTF
ZSZHLVaCHzpayR6cwkVCaIXeztNmLf6v56hHJOMOLefENucjdJV/P7fXSkBnVR9JIQUSF4BV+JfX
z41+OLGihDeTL1f6XoJZh4fvs6zPrnqtZnkVwablz4QDtJnZDldU22IFVgID8EzuKoLjmynWjyho
3QNh3uapm2X39H0qjR5BjIdycCiyAll8C7sgFmOosuG3+msNpJkz7DdpodfLISxy2KUiBBGv3/Eu
01ThiaBHZ/TMBWarLoz+BRJ2Dn3jzDCh+GszyX73vLTAofUtJpL6pkqUSBhvlItosY9/W83WOu+C
oe03FOonTCkk2GXwr4lvizENi7LxuUU4PrbSPR/M5E6fMq68N9a3nOnEJz/0Z5Fny1h4xL7mK0eX
NA+xnm+QhMVJ/43CY/wbbhL2ragGJP3vz1Z4FAw+q4ic4LYowW1b2xhdGTrP7wp7PBFvGZHkFDQw
1NuiSdpUav6e2g2Oylh4uonr2y28k45Gf3QkJ1prH4CMNMiv3T7ExKf14NqSISMoiBJKjVa70H9+
kh8Ldrp+PPTK6ssgJL97CTD2l6gDswK5z6HHtnSzmV/AirS7Oz3zCrf1htT3YofOx5CJtxgFghS+
iWypttD5sbG/JjhcOtz31NUWTi2RR18pAzeimls0vIk7TAhJT8woy4mE4GXb3f/1KbZ1f+nyEBDT
kB/BxFE4i5VYEzvM23aslZW+QjFom7eDyMn78SL8FgClzNlqQ8yVcsAoMAmnoBU3oxHtKNob/8pE
ixr00nugYMGPIl7OEs/zAHVoTronmCmc+8yEDjoUosqZ7nqBqliI8WG/e1z/9iYNmv5kenRSQsrb
bVRM3IsGHh3gYzSgIwu72qIiCyTHv2lPLDOieDcjGBI8OWc/FthwNXitDa37npUFS4pDur8bhawj
v7fSI8X0WmAKMWVyxdvvFkzmKk/qFJiTVKJVVNTAboD+ABfarfnxLTgSwEmi0bglhV8SvLQ9hxb2
QtyRUNDJwz6ltuCJBjac2Aj492ST/AU9gu0OF2mpwR75tIhymVuRtVdbW1JYXGsHGXV7XqrtPc3d
5rcQAfI7FZneuZyLprwVVDlTBOXS6zuSoRhdfC2oCizu0UXmkgREbJG6mcLiMIn7+apIN+ASWjMD
recgeyZ8abKCoPtYkV0mfk5tZoOu+kjl4iMD4U53pWftIk7wUusfJXlbtllDolZO9RlZibpCFfNG
eb8cyBHPTuYItTbr32uCUate5ADOeqvbpx577G8RbEMgXyZggokfVCqbXJRzzTvoB8tnweK561y0
W9jWi9O6EloXUJIzwCzlLjJXhW21OJOdSpp6Hk6A6rhis3y1nHrXwDV9XfZNdsOKUo7d1LXjXPX+
rlcsvHZF/lA/CxE+Y/UN1gqnU6aFQt5BtJo2Afmi10qs3uhzWulusfLDnvb1gmOzMo/sFOwkK+zh
K4tFfX+GE6SxiluFyZwfw0YQCgbuq2Q4F+5zpIv7hBmTruoiCo7WyC/AL2gCOBdTn4+Whg9FrZlC
0PNz3ApazcamojsR6OwxZpW7cDTMCMFkiHM2Rbyl1c8qQl3SlTx5YDsKtdeF5a/WcoB5nWhUrWHs
Ejz9IxbBhMhDHUp0JFKd0Hh9iBHWlyctV19kikw2XR0Pnz4YHNEYWYNnWdKOI7avFbWBWumi4z/A
wmm7JXQ3otOW8PEeBA3tos48aeSsLqPYAhCU8WLjYPsGUL/0VZt25kfYwvoJMmRiQoKWOH8zJ8qz
hatiXRbN7ZIlrr6vK5zkdLyroAYnrJSp8xrZtQnMSDGJnJS2T5OkeNfkFQsAxqakV6i+Cz0twnVL
8jSi2hWds41B9V1+q6iFnjBKpNMSTCfgwIxeeIs2b5rXjRqSZN0oBLFZDwJOSMIqsY+zAGwfRhvb
9SF8m8rfKqp7AwViufnNOLOe2RJpONKl6tqgl/nR2mg8kPAWnstVNuSmfXKz0sJYRiIAOilO+00A
uvitE/NmmfYEREt5A3hMH7BYW4xTEDJN6o2xRQxPoeQLuuRCRVxvKWqrj+t7B9Y8Hn2XPIsdcKFn
xpLFKFK9jTbby1LkihlnWYdDCyBytoYLqtz4EGm7eG3fWcupU+f5LPtb/xiPyPa9/NiE4Q4FcE2k
cDjoTL3VRdlLLHGC0FZ+iEiSQQ0D3ljPxoru11B6rJ8AiiatGWv1ALQQ3SnqGEmc3Ad+PIBy+pd1
SydRDAW0BmdPH2s6zhHV670kD+FDbxeiHo089L79Kma3hZrzUeaVYsrJFtiZ70TjA3zmLkazRQYj
t5HBqPYIkHXhXkjMjKmvfbhmKG5gNN43MgM8OwB9nBykzXnUCteKJ2zZH9H8mwo7JUYcY2pH1L1h
6ddYtPoeFYqfdT93pKjivPoJgCsq3dbzKKQ7prtK6GxKff1VkDh1/C/YEM42fmmJRJxwKKVGpOmu
atYgLRdxl4FIgEzHMIiS4u/9ORr57zEaqwZvZO+T9A6lukatQ6TPeNVPYINO0o3kD7J7ZhO9S9ga
pigtwxDXdW6NUmKt4uuXPp7QGlzRwK8fj+ivDYFSxfJ4pLXVPG/2g2DEipG00jReilgQ6JdGV8ff
W6wu/1BhKc+4G3DtNGDk7TmrpCywfM/ninleesLMiXmgxn+mufZjJetHrvFca8n5Ipe/thqkOrCe
/TsnnCNsBv1mEyOxuhDSUIYVjvnic768in+uBDgoZO9DndU5wyULhSbNQBu7YSt6+s2ojf6LSJxz
GzG9XlPV6VDK5yCzEEulbbTdoa/l9cpO1oQtGzFTNcXiPtYM3cx+Hpn2MQMOMK3HXYDT5pDMumdl
kKQFtIpY1L9NNJ5Y0NYkm0ga1Gr0C4ck8+KyUxENgMZ68iJYSwWpDprJwBR94H8Wn24MMJq6aHaH
QlZBcIqz4rkou6nMEFkUBIMLbOmQZKChr8UtcAqOu2X6mpqLrKqtxQmnUUZK5GSZmsxbqREaTQAJ
73VtRvfkKIaFj7NLQCvczyFmkO2KsOd72DEB11BwQmQMUTBxxrab5ZahKZ6XYW6iJgdo53gsnubD
bfQOIHtFtmj2IO0Xp0l9cYQuRwxEfY4VTgGfUPDmotAKqlGBWXuP9vwW46Z5JzXWBafLV4DPS2Gc
35SYnaM4gvP7K8RtM7tiMqo0+GzHYS5DKc5X1IeiCW1AKaDxnpjO44Oc4BaSUpFsulHABbavdLc1
Aw9GlfOwe7/910EEdLXtOuQhfRzChxv4ujD+lGKhc5A8ebb9Ni0WsjbmudaMljZ3MlmnfAgkyYqc
gfSAEwBe84fFj7w6gv41cRzVDvOfPyPladfsz+uOGyniizzXhr1yH6uOnUJ13IVzp0OQn6yakRNK
PnXNoeUf9QbGAQEthFD/1fg7uqr3WscQyqEvgOcF3OWrogxc1KWa0Fz6X0vIpaJmHjqKQwR3cJ7W
5duI4KahYnF6QYX11wwRGFTXHrUERU2sM3rjid73OY+oQ+kzG+kjdD6JSPmkk5izeZqjLsI+1vg/
9XKNqb/tUAVVroO9GfOIY/TTdYs9z3hEdGB/gMkfwZh2H9LoI/hjGBiQxicUk9cDq7WQ0QVujcO/
XiZlBGFndJClc/trIfzPCHe3o+x+YGeEjuafKyyFcbvO/YfFFxPyFzS5bt8N+IViZXSdWrnuRLDv
+SKgfjwwTlno9NErjXz63OXvRv4TN/Vh5jFTPQmE1Xa6ZsB1fw1vIBHrWoSKgUe8LApQvx2ECjjl
X24KaDy+NHPeF9TlGIBBrSIqSURkCTF3Oxm7ghInn0vu7CMHe5mqMHkltGrV9HhDrZpIiPb6sMqV
ybR8jnl+EKtTohJpJiK4X4YABZr6fLpumvXsUnSHj0nb5QTo/rmvrj73eMFbZLaSyAxPpZviiQUF
gFiUIOjitTpPuNfSNlULWnmhdn/we9Lu2Ri8m0yOI3Nr+E5Le0GyTZZdx+PpdQb6+xRz9Gv7B8+E
dtf8sXJtDxWMMCy76XqjZvJGbGFU8+yJlHEXwTIhHG7Slf2WATFIvzBYs6zC7ZYfwoXmfHMlffw+
w9ju2aPr0W2T73QZdSVtT25fawG1uGsYf75DnNJf+GCNTlPzgtcxnk0d0Hps4WytLhszICqV4zpe
AufbYFc/p2xqGSS873u2/5yy44hkvYBG0S3cjIdYDIFZuS2EA2bc5ErrmJ0sV89jttIUWrOdaMih
FaWgOu2UnBZnG8y2D3dpG2RciqtRHeCID0ZioA9eUM32lBLwhCYZfmboUQjmVwAP3JYru3xZmFwR
4KKSd5Tad5oTLkMPOjNc6uHYLNXrjq3gMQp+v0xyR7+H4ws0RBXfMLj6kXxGM88HdmCS9SxuhCGg
sXtiZF8t+GVLTwwV4eit62faL4V+UISKak37/3QF85tH4YQF7KeXGkyJl3iy/ygRlEK5mIAA9E3g
e8dpp/6fwc+RRPDdSJpN8myOyvvNyn9zZz4DMXYfnV2qAhiZta3FfnX12vIgYKmkjRtP89NWvsFi
rDcSLXYayPBRjqGsU51PnGS41CjHsXlWmwEnc1/mLybFlJL1NKvl6jyI/mtwvBqgIYH6nN2xXN31
eerrkIoXFhmgTswdUKKsZOcpztMLzBumGT2WhH/ZMH7DC/eW3xTGlrvz0h2iM8Ru60K/4dd7o7Bm
iNx7y/zft04gYwYG4XHj60njXk//KiwFMY4iOgAZPHeEeOV2gqZiVdicRBbmsJ0Mx7ckTTIT/4zt
LphQyPRKh30qrXoBTjWnLeyoPrMvThw3HJJ1LJpDv6FXCfWNioO6weWQddNIqs5VFx6e9l7LgLzZ
kgmf5GKPuveDDTxWBY9AYte6f+dLIJKw3PHzna0OqqTQHoJydd3jfO9jVTQYqq8By8g4vdeUFVH5
Qz9xAbojI7IcracJafsxRFIbQwoxTwMGTPU+3l6X5JM2TDT7dO8CsGw/Ohmjnu9tBjiyXKo+e02b
HNBKYU+TtMfX7rgTnENC3fiMWmFHqaK4xG+d28RWa6HaEa3kzqrWIh69bV8YXIFFeV641mgDqbQ0
axPUNM9q1M87KCizs3JxbMZZq1lAI1l2ZC/jFgoxqEnnggtcYfWkdk4kbGUT4uW/X78jfTCs0tQM
5VBF5TAGb9uXloeJ4frSxegmblm6IlCX3GK90xkwUCYAKx/N15dICJJlwY98BkV0RPwUSZ1V+s9a
K1mN9b5inbLhSPhQA7e0h7CvgLWYQMgpOV5JJD0tePYuOM9NGZu+ije3k/BoAW1Md0d27VhBViuJ
VViXmFRkZgJsbv3W99ivb/OAgjnCh8Wq7Yjf4KMp92UlH5WkindGM9KM62a3gss0vi/mOMiN0ErI
yEy3JimBbjEii/bE+zD92nApaBiZkVAMZdOGr3hMwon9IoxLpR8NWUu3O5NJKq/DB2ebz5jgqP3d
pD/O7F3ycYNTf1twyrdc3+1RPgOaPHO5Yzf3MoF0Lu2r1IRleonIV0QfTPyf46W+jURD8ovZOdvi
22j0tF1kTTD3g+NOjkEFKW78oNwAZYIDk++/Tj98WStPrDiR+fhYpw0VKIWbtF3d5N5FYPg/O4Zl
M427ip/rX83lgbOEUnbtgUX0Ac/Rn+yF8msVeQiITlNesIQXfwgUhB4HRZd+af33zCiuu6QXiF0y
yxCKK3zjs2Vognz6HW1s7HacvpWpxVzcN8TEIk74eoq1YN7eQFWUlgLEfKswvj0O9b9quEcaYySa
fzklUzdWXeiDC3prQ+1E0opFNDzENBlJU8ZmZ2H9GpR16bqYNHSWlQ/Dxec6sMj5QvYMj+X1SoNy
+OPnMJkRU+hg7s1a557Z0vkQuOLEcIidQpvFTUDeW76dgjv11FTEvOO5bCFXA5JECxK54YAqSjCn
Qycmm5CPXDMGJ4HqDznye382A1Ij+mKOAlUf3GW3xSe3ERKYDhgaPXzfhmwwbWY4Xi6NxV1vVSxE
APrzMGa50jz1aZIBdEmk61KudWNK4aBW0DQLrIfMamMQir4TZV7njLJIcbdB+oPH/YAjT2aCBCbG
rBMwY6C/lYgntAeI9uJ4apUp88vX/arVMYyhby7FInGRGHBiPFMffjyo2qgvGblCTv0BS/15Wf30
N2WDrbqoLC5mCyvhK8p8/Fh9B/m0EDlG7fl+v3GbCGnyRJuZUBn20J8SlxTLtQs2Mp76DzwcCvjj
VrObDR+/3X/1pUHKig/lTXDPtzi8nwMlrEQfgxc873dngKbzYKfaSNqLJego94SQ4a6IhxurcRoZ
HxlvGbWbr8GNQP483p9DOgSZcAKmYPaZupFp0oeU6TJNeeiLqf2ZcstYjj8NqlnLZZP23CI4e3my
CIIrUllUUFU/A1yumgiGj7dkk6Tpj20h8VtGrocW/No2XBvmpjqUpdMF1Tpym0V2PkM+odqOFxeO
hMGKLqd52TPwwaRw/d4AbX+tceeKFTHVSdT6aKxVV9ISkAD/v3wr/3pufYQUJj1mfXIFdpdabgjE
E37y6PW3P5TeBZaI3sWdydDTUElpXcFJ9Pl8248Vuc7NIB6eYcPNkluVXJIqDdS3KW6Ud8w/8jXs
Siytw+QDrodWwXj/799qOr5MNv0FTegM5cLYNvTY/B5d4UNsmDeav1EAsvAUVHZSK5aV8Bi8UllJ
b1CP+UaB7H7WLd/slVCqeJmlhWveKWFp/1pikb7jjr0YqgaBTf5KRYUFYi5ONjtRl1vxvdUZLP30
5T7jlWF6CSnYU8uOJkafjhTtNTFSzJZJ+dHQ066VL4VT7fSJcN2VqnvEK/SVhU09utlLB5pMz44O
bddxIIwoEUo7bVFS2EKg9a067hGpNpOBH9uHuabKuQVXFZPJTNZH7ItxcluxGcdmR9hUgjEh6o45
b9fW4mkyp/nflNJnwgufFsdlHwe6IiEawwsaxyrmGDSUfFxtvGPcF1YQQHl+dlH3i+5O1w87BF89
Ex9JZ3TLG5FrcATrUXvkcj1lf0Qmy831QZGhlCoqM0tjTKI3iOnGXxbPrOoKIMSwU+rgmrYN+YH7
V2U9wjYGoOlRCZ1hcGi3C6fPZ6tey+kbduksRQR/6qL+3kSsuceuSRsM5U8GqgZZPRxrkJ4nqGyt
udd+Uaqq1szuIhwhejv+VxIery2p1BtxRDkxMbFv6VbajJM0k4xMnG8dZ8O8abo6ephRtVo67OnP
T5YfzTTL1GLr//loZW4KD08Zr2AMzR386NcpdrxrhSzdtye0i343JkanA8QWVP/AMUkccoEpNJiD
BQ5tNfBhjQFRG/AibKrv5i6T95xsCdKFu5M8jjHz6FuJQESdF1kCV3iYaV5fLTiOKa/xutNAWqaQ
nQcgmvbjQUi5G7GlLmSCn5RdXA/7N3BvVr8/58L0kqsR/vyLuIfWqBi9dzvSjyFS7vj7QD+1dP9B
jCH9ksdcgvR88QvL/eMYAMuzyV7ZI5/2UskuNbfOva0CjguKPPWD+/uV0tgCoHQl3q6Z8HA+r8jy
Y2UexPn+9c/D0eU2t3j7SZfqoB01PHMDEsptL1mh30ED7wMXKi6wBdooBlAbhWSTmI/d5uangRuM
V2aYMc9glsm0N9N2N22OhKAjj9Yx3vzyB8hTNWLNsSI9H+gcJ+9qNf0qM5/1er8ftPXN7nZyFMbi
fVAuTs7zvfSxss/IxbmMlS7U1hC7G5LZfhhu95lyMRJWe5IgyyRcqR0sHDjHFP0JGv/2pCe5HjWh
BCWgldBREbnI6p9hAluIqOBdf/qaK5sC8GBprVi20bB8kSG1OzJUNVtb85zSPlX8+IhZV94/HXiE
lFOYtny6UVL+qJ985eioQlE1+dc/eKSbAlq/pPYnNsYkPyV1bxy8pcdi8+2BgBdWrL8z9T4SS+Jl
z6V9WqLuDYByYjrmhZHKzh34YDlBBrLcdXgvCZRKlBimTngK9eJfpA2QSPg+b5xTYz6FCDypoiie
vvJBJAcXzIvVoYVrA3KMcxm7YVnaeC8BeuveSQUafP6UouGOyyr3umpwt6FpDp2Ds6rjxfIjJsvE
LVVKdxiwJu2K/A6/LBFG4ATGM/PtkxM0JRdEWUm9MJPsdYad2kIg5hm26E5GFJQ4TU2Ij5CllQBT
ZIh7U4ldsDGt8qxCx3odH66TBnylTIPdvsc5wwEOVpHN0MTZ/hb8PtLyL3keBsZMsYOpNIaqJxT6
EVnpvpi2oLQegiNFle/9tQiOOJX14WDxxYfsvt08e45lLyDhrMFUaxfcSKpHqahXljIEW9HQqAtG
yMmt+cAdigIOWP6V0RF5En0yj8dyUNIC/dUjnToXEce2/dWKImzCoOOgiKJUtQ0Rq/s5xOATED2Z
6zbwWHaKVrQ5foUNBVW/jeG1CvLBX9HaU0gkpC8jFU6fYIeztuV6H1hLRDfphiwZqYmcEVRyPr3E
TtNBvxJ1/vS0fwmkRJ1aTPb8y6JGCTJAtjrXAZwb4VBTt9Ye3vMJbBKy1Tt3CWgXcDkN6XujlcVM
HMl5L/wb8umkZSuZPaY36WzNdYhWRJ+Fywmn/dBYNvVJHoqQN0V9nO88SiNar8BY7W9RCqcMFHTi
ujrUN3mx0rv3h00BBjg89x+ni2F54fZdndZM+XCG7ovVn59BQZEEA0uGQHFBbACYLIrDoYdLGt35
4EPm/K0ZbybA8MgZMKXyY9kZ6QJ5x8/L3HaI7Y7fVvpl7wjGw4SZc727xBlgB4yDBHZrxMErGsCw
zC3uRE7xIvS+65HwrYJRNZFCGAfhsRcYomCLUSmjTFjtp2ftM5c0+B9CXlnlWoWfseg8YJrn2czc
zBx3hkp7V2BL5U1DF+yfc7Lnsj0R9pnEyynCOq45rUMhdD0fwbk+LkW3PO3TCQ4mju+IVH9Zo5/o
ifmEdGGbUVR0PTSybqCitjr/zYibc1wnQzLoig+QvV5/TGRkRZMa7cR+ObBHjrMeAukvyfXt/Ab2
RkZV4tCOVhI3p2bJrvf8EQt3BmxcmQHh1BXR0JYKyKwEC0OKIXjwSxjXzn5GOFnXVKwp6mzsZtGF
voDxoGgS8TP1zfclDK9ZGcxVKQXv89c7SgJ33pSHWK5OQVfBwlsoJ1y3ApKd3mpMcOjPGqFfcUTp
4EQYxPoby3AgW2jhQaZSYggfxaktAAkS5vL9MGbpglj/Dld+8JUhYJducxmCkA7CpxV14rxCgTf2
LM+e+a5HsTui0rJOX3sp4Ceka1GLi5g5ZQ6QQmlIIZhJ7td3YM1+olUr6jZZsAGPl0H9PGviZ5IA
njv+7SJaf4xb2UddzfbQ+00axzbfjFKfArjKE0gf3pyPmoZhLG1siDLn/r81I6qoTXlb06QbVF2L
CnWraZD/2mXAPTvVJyYHJBwidCRfRFWx31A76nkEH+uKoQwChEtkhF0khj6j3HT+X7vdbmBPJtat
pgYTuqz2y/V4enyOnNsXC96ST5YqYY0IHgxxvQifSHQOYtLy3+LBT+FsHI2I4xPLq7tEVWhWqSpl
vP/+MCn0oXJHk8XNvKXkeyAV933p0jS+QdS5rSOZKL+Jo8CsnkJqIpPydsWCGOqVpGWaL1wp9mBL
4WWl2sypjFgEwK/Ncuq06ynY0poItoPINS4k+5aZZvKBen+1jk6i9Cserp/3mn1mwZPH8o54mSuF
rpZ3W1kBYiPdC/hTLWU5Wo849xxbQnUyhFQnxcJryJ7jx1/YCagd+pwRJ8IvepJcs69Kl3AOljri
c2jTOUeYA6jDzrDjFja1Nr2zfz2HhE39dvPUARxEhUdkTWigOlKx2mGhwiRbwGpQ6HjfszwBQ5X9
m52LFp8bWXMzcbrO4p3WO1SNDGMokFKz0y2ta/odT62BMkZEaING1v1DnkqhDYlkd0dP4FpR+Clx
od6t7maZQp54I0adEaTUH6prsughTpXxA+GU7G8Fusry7Wes7zw4z/BfJfk/6wY5ChJ+Wu4AjSC8
k12fwbkyMa0zEwtqiZfi8QRyi/0ezuY/JIjoy87ns12ZtfV3Hax7XMBHfwh7s7rRIavMZM9gIU+g
lNTW1UAY9R4ztrOR5krtRxO+AGYnYYLs3UjCgla2xXnxgMVdwfP5KtZkrJ2ggRGeUoZev8/WyXRY
5fCAPb4ijaHwItgAjCOWAxp/nrXtVbAHS/R0hwfiNtsduo1uF+kAqtMkJ9/xQJCHG0DKOc895YU7
2V5AbhwkZDH3nCFhZlck3Ml06mAp6RBViLjrJkWqvRok+kI93BKMLac2Bw1Ou4EYCeCnI+elhcQQ
1VwKMiiSiXgt9Ep+pda3eJXsAoTPxclaAE/3x8doO4FP498dZrt3nZLnJsdTWdOc399Ip5pTAF8W
yjbKBk7OzSVz4uUWPSwGnsBRuyRYF3J7ZZO98MBDEG96ndG3wZVt+TQLcgg9dQJxdWLg7OYFDTzg
jf0ogknC4lXsy3FbL4u8BSFYIx9CmAi1I1P4z5ttPbI45cqdKPHP6QUntuXILeuQk8Bu0B33Vr8V
sA/aqwvT/a6sui0eETySGx1kmYpHQs4sbMUQuGeZv9nv1xipQ5dXb2FDjquN+hE0A8w0cuig2AcL
qZQq+eeW9X1TZOgkUI3PncF0p/dWKTV4C3OTaZc2XTPDhnLMYyTnrkLKBcbAvt5al7oLZlHxtzjJ
mSJSPLKY0xNju1AxHo3z1gkkYk+9Je+cqkpgV42mb+BqIJgD1bIcfU7vuQa/aWHCdyBr7F7kwWEa
glMnEFGa7qdvBsNLHohJeG0TNaJjZdE6v82rfEhlLqdD8wHJT0dU6kuz+gH59R0C/ctYZXpRF2VM
rfCsZ8NreB7x8UUPYQxL7YpZgd0Mko3rCiFy1GN7PFwguQnd0KJ8bdIEBCrCyrf1AnJaY2415Ym1
8f+nTPYC6b6xBRq+uoLlCoLx4vn21LDaZPG8BbeEdxj19/4Fke2wbQPEL2LkxgHobCm+ORmju9NU
yiyCYoB91BHL4BYxFbPKdPLTDGpnXKvCpuDq/M0034TbbpHmBS9jk33ech4G32uOaHlN9AmIAUsa
bauTBdQkgTB80pPG4Y5R5DFgvjmgxYq7z49tSpZRLyqkaNS/f8Bolg/sJDrYPaT9LD22HqzdG82E
Bmg2I7zu6PQ7ipHtPw20ZFaGYR2khVmNbGajEkW6RCth2pRh0P4T+GJ9LwHEiOlpgu3YebMmwTp1
+gCaht0uyY2+HlrPaQvhNhtWqVhXXH78GE+t0Y6MFTIc0yG/r/emWcSBYm8OGyWV6naYUu2sxW6s
jNsTfGOUBWNmj63gfXdlBJRXQLFjFx0auErgNnPpea/nOWsSFR2/Thh47PRajV4nsaY9aVYLeXtT
XVZPgUTO/Wvon6ogGFbFnkfETBrMXkTgyEteGO6SklMXYPIONI8Rr/Yzjt3MadcIDyQghGtOWYyc
UD65ENzVjAuoTzxeSMlBddbWPYHhfU5Lccxdzz/xUfFomG24z0ZL7XGulzkAKdZkbQb0smTARx3e
yEeTUZmZWgSnsbTDQpNmQemKbfgdBp/BWABVCX65wzh13CUt63JYL2d5i+ZH9ZXcms1wm3UxdybL
dTNkxwxSAXUDZbwemMGuyKP31l9tmUpiQrb2L52YNOSaA/W/Y2TJQZhUEQ0bAXzw0SyxhCfkGTAo
qYI3zJjPCr8Bsgq1P4vGMi55Dzm7/FXIQIc87/CB2xOSgz4FIh6UIPB1oPW8OaL7WAdPxpOEGXac
TESn5USZI7NIbu2BPwkdp1BNCcA0r0hLBHChvq3bsrAnf81RIm7+NTbbl/TEYSv9+Hu1bPnG6ZpE
QnI4UizRa2Nyc5NAcMgVBi22+JB8wURtOUJbSVY9Z3fl8sckmQ7AjZT1efte88JeXdesXOD660oC
mBJhZaxCtxuoN9NsUEkmXR/PLGo8KSWBTBp/zYX9H0jGNnrsgdkJRwSFwntd1ayLLMqPOExwGKBT
WzcIxbEcmk8c6sIIAjD+YtZxtdGD2tuERm1Z3tZcFu0RmSrPXTW/M4ex7hMkVHD56OGz9P2Fhwso
dXaQMsKo6q8WIrOzwjSCPYgHawJ6UMxK4AmoLSC3X3XOWa6l2ycRKewbxGIP/FaGbK7Yw0EV/32R
I7NdyBgvDGvC3lsDCEHgVz3SG3A3zZ0wxrK3dzLWLGYhiv08ftrGh1yj97N4ZU+wjgFA8trRX+np
eQ/RYh9Zvmho6VjO4sSFRQNJmr+a6jDQE9YnahGno8MM+/F8z/lIZPTyM2qvESTo3Wn5Tpk9XDDj
JwJcvpauqXm1dmikHK2KSB58+Q6yNhgfjq8qsm/R3Z8RcuFK1xw/EMnTHwF7ocFOWDvuCOZoix0t
T1CcVvWEQebLN/Ka51zJ6tDpRMODHPlXd2gZVsk6zgmB7fdmAMVbSrRVbW7H5/U4S9qIFyfyCOTx
zUVIobjE7Bhk1LOW8L1CJlB2ePsz35B04fpdvpdyyIicFeTfPvz/7tzUTJIMiqGl63HYRq28V8DR
hX+reTzl59nm14Y7HdQ1FIvH6LQiUU/1X/rId080n+c2B+ch8o9r9/8xTcgG76gYYi77eotst9Or
m1SLBpPes6KrYObcH20MPLOdcAMk6DlJD4R2bmX9qLL9D5HWZZgkZYa5207LTJbdGdzK9obDwNOY
gRCd5PsGvilj3CXYmBWBB+xbv6j1d9RHXLvi9qHEMAk/j93eteGZv5t8Y3TgyJzyEroutaVXsu+y
YdBifncXgw4m94rkN6lq2+XMBi5Ebphmot7wAOxndUb+1HtXIq31vtM/zMWNwKhIOIk/wdFQeq0o
HczSG0iW2ngSFbB+sbzNMbU8V1Is2d/s/wGjt8Q7nm6wtHmD1RRDySgt+dg8bTmSs8hv6rdmaA3R
2qgtWBzjnRtB5sd0a7fIXpsIe6qmXSgMCpMG7r+dI7+FvEq/5yNui6/s27cY9cJqfgYwSOniCaQf
Jz6Vx2PXAE9HhWllqbS7lE+9eAvXng2XFPXYd2ZjEJe6O97DIs2aVBjkAvwqnLXhSYPREL12Y3SB
Wfu9HvMIhlI0DImoxpPRkZVZTnoeJ1rNOIIvyYzCywgOCimZy5aq76SZpuTKYPjfLzKqQs3T9IHR
UecAb0JLpXy/8IcP32U3CddJOmE4aO0GBx3Y/qM/Rif73xcAS5/E7a8V3lWFvj7/dGQ9diOVellb
9HP6M2Z9cZJZsS6DForLjFgNDImI9RCYTfqC+dqxRiqotRJGTDsfdG/wlGgxPqES0sHFKjGh3ShQ
x4SRyDHnjektYJkWFgJ/FYUTxkanykU46O8n3O5K6aAssxLjRKlTL8VTTXyk3Nl3XKvG1102ADn4
lC28Um78J6U5HMkwOTCbxa9G2YYGAvCZnl9WmA1veqZ6fq8MMru2HqA4iwcjxkekR7O6UVdVO55i
mVqmXUPkfh3Uexw+BDyu2KeHy900L2d9ZwuxWtDhT9hBytdXplvWXXbeYnK4fj1Si77A4mVWzTQm
e8lvXtaQkZBccO+mnNI0zhUxLg9DrJe9eSIPL0i/8UPaC8qhAOwMDivbKMQE+uVy+bkUI6ErfQOv
fXEpM9Y5BbsYuJCzaYtSy8wmchzCvKKM2K8ZZhC0W4dTSf/+DQs0DgYO4BnJpRYK1thbSP7r4i/e
uWVNSpXnz9BF7mhVJEZgReW6M10yO+BmXH2rXqtnA5PQ2Sg4vSJWrpGdMxvemMxrZvi8bkCmBuzj
du6jz8skbiyhzOQvTIZmBpz4+TFp1+wgyyrwZQZ+TWsKo4ksrguMpo9en2djGuf1Ma2DcAtL6l/G
d7WxfTFigBQBWPi9ldPgb8yuF6HFtJh6iLdW5JcPVz+5aNBV3G2+fKlqtmoTneiGadoYHkseQ3XS
5ZRRLTvHoFeKfbSFFziPwzLuv04vOGhbnvTFVPP1UkDT5O7d4GAH4apumGepcBVb4z2Olo4QnBVb
BYlEHrR0+XenJV/GA5CtswEyS3StN+8MbujHyxb4EXDD/x4ALGBuPSASUELUmHvr4SZrMLHiAXmP
ICn4HcTfSxPoP+Iv1S04k14mZr6d676bfaErLUWKFXQ5jM61OgkAeXCV0Ovt0O/C0ggJhGfZWGL/
cQhqxd1SKpqKlONhcq/oNsbC4YDcBc6WzdD9+1IWDGAzYenCpPQTOzb2S3ZEy8ZMVoELofh1m/hm
WoX185WuNc90qlTgT7XvpaUCRD7+Zlwvebd73TvYYbDo0yl/uUkKg67cbWdkstLWiVGeQ7Gz2aBv
SdIG/0J7IA2XgqePpAetrxKD0O/74tRkwi8IyClIvH/Ogx+RKvPql9Sk6fvHMqCWw4qo/vnLgNqf
isrYS4ckSZNlr8Im4nV2DcO4fMTV9RW28XoOPw1AdzvNYIjDh5rnYX+n71gdZlqTBTXpQ0YeMOhV
ybgn2N6PJ78kCo8svdZPMFmH61KgZ45o+HGq9ycesh7TJDYkJR2ilheoFNEuSZcPQc48i9mnrK9V
kE6JbnO0a2jcDF5PZKDIujauZ+1WHPtFBBoniD1bHrDNN2Ft9ewqPITIy6hWWmZfYC77aGLT5toh
1b/JdNJ5Qr8YXqADiVGctPAjrFGDp+7VfZdcM6tvLCrwHK9HIMdEkhEkQZN8CiPvmG39P7lxZWMl
ktvRXFNS9eUyljK13vjOJTUpuk2BXvkK/Dplq/41Fqm29J4tTj3rwE3YjD1Rc6/05Yu7o6Wxn8D1
18//ZaAc1ApX1UtnG/zFCO/7iqM4rpGSZio2OGIS630kKR7uiVYkJdBRv2+k7GqV3knEvVDbbnMV
WC7S1yKqsG7sTII4vYk12ZVix+mXo0xFGZXGv3gkiwCf2V/Ysxq+qzXMo/2HzTENxZnnfp6dHJTz
Zpdc/6JJeWC3ugQ+H63Jy9tq30xgrz7tObVVEx06Xc34SPz51bqmo+7hXbGcLChWqrH+bV1ZMSMg
TLbxVRa6hKS3g154iKfpqsCRWm/1gfUJCTN42f09J4lqdDDRhQDMtOkomUfvYwFIa1Nt4oMqvjKg
lD/dQRVCkrRrSsdndIaOo9L0H3sVVCBwKBsNAuJlXsRJ7LJPrKgkgzDahnncva6KX5713OmANOqT
sbg4wovfwVTyPd7SrzxfjIXuqgodz4oyRSTdSHDe3Fy7VBD9fyDBbiFrk1TNsJwl/cMmNCVJHPG4
zpZYKMsnoLjPdU3Fk/5kdE/ZoGh1KTz4DX2YbCS4/TGhp91MsfcTLbzOlkweMcRDJF9BRDa3L/B0
6tvM9CMBW/7fX0V947u+1D239OYTX9FLTv5HHzBQQKG1N1qhAKGG3TVxoY3SmKxVjOy0JcV44bzD
Zuivv2LRYI6PTSsWfQBSMwf8dw6+xwSAJvJsH2uSiOU6/9vnn/b5Ct7HhXuSXJkpcYt7auiWgKWN
gsiZ7eWc3h5dInPIIqOpp4tuWgH5B4+xPnOcnRhiBALwPVPoj2vxbGUx53uhFsvtfsHawXtX7Pu4
pV5O6FnptPAAkt14e3WyyzsTZvHb0Fi2hZahRdvGQgIxfk8HgDuSzYtVah4sVuvmNnNSj0PQHIVX
CqBIhTRvjw8XUolK9M3objqWLW8oo0Ji2zptN31qtqh5eov5XdRBXQudmhYByIUSsRW5awnVqKEa
FkSWO/mhmtEC73QI4Ixdopb90llu4GtULwaISdq4DMI3pSVKALnSYu/9QYh+gguYdlk6pcARV268
VAOFG8X7pyCrd9b52psEkO06OOQfjkTfFpQ9zxRyCa+AHxLD5XhzVT6h4jn28vuF+HVTncALpBEJ
eXdGVm+0sx+EOuFivtgYqz5Xp44p7vA+jxxa7PD3LqcuGIB6T/JWH6nANtzhqLR+ezXws5Ilcn7H
eIfLVgrz2/UIc/iV7ldPcZFnIBPys8KojrKZaPCOK+cESELq7NPeKv/y/TZ5y8oeX9Tbxw05syt7
2tPfAXiPV0MxLowx2Ea100Ak3eD+LSvEisbjez1EkWw1wFMabCAGaTOPQeZO+MP/KKG8TPxhaRRi
P3eomjTdEmmdRrtPzpIAduNj9ZFKUyfpqre5NQqcrAz6k4XKV7qNAoaiuPGg2pIPG6SnaJ5X/qv/
p0k8gTyAFYjwOQI1/O5IJfAxCY8z3FR9LPUFjo654LV5R/5w2rCOC/BQWhQGdeNYnD91m1IGTRPh
VFSsRTOCfag+4rOzmudmUJ0fFJqPylx8AUHbtX5J3Yljjl2JsM2zjweyOSTInmlo3WJrn2cyntx0
sf5W1rGvFapDXZ3YjRmEXPB4rMAybPztdqou1H9CXPZo7xA00RbUuhYIQ5V96MHoQE36KLXz+4iX
1N3NKzAAkZtlG4m2iQyhHIDeZoeLevQdZJJcrEHDbrb7dYDRcgFDoiUfqOGFux7uHCtZtk9UxSr0
NfAdszspOLzQgeJaZ3E0Tq3Z2tBjPJP26bfwnOy9WLCCfdcMl6BHt2S/LBsZoODEMr7gshxqmIAw
76VvbD4HDTCeBXm5jMOlh+i6Gk128hG3deArlOWzLraIY3BHPd4AGvQF1rp8wUYUBmrgP0PDtBfm
nk0tSvkgMWE2uH6GZUZ9mxi1Uj3X/iLbbGQfw16aTlRcGwlBtB0tDFZN4dN3IJgPprfB6lu05uAl
nQJne+ykud9d3TviFM732I164x2wzlgJMgYNdnTOgF8YQrXvpYnq+OLyaGXeg4i6bQ1cU+xc6Rcx
Kn8dliXCqZ3PzzXohVAtXlewFbgW4gQLylCuUSRdddLyiibn7eQ0xnyjTaAGuxQBroU7I8OriyDc
aWRnu0rLLtMpVRqhfMHz7r6jvA170Q0ljoDw0b6IzyfUQsTOEyQHNnUJz9Q+oFvJZT50tLtbMscC
xLpjNimmwZ7X4X/pizoA+TWt+iDe65kUNqlSZyK07d0nd4d0KRMtcvhzTXRf0C55HxDnz0ZrNdGM
qQpbcuc579YZ0JrX91uT95avzB5251uTMY0lQR2TANCuXyE07IoRvmCJ/JUBS2xnc8uJ+FdfPNiw
M4SHyeTr6oxWD6/HVK25doM9KA6xVzinWWu0+IB3cDtdjqQjmhyA5dsyBFQe3s3Ahovlyg0u04E7
vpc6WSnSJG+A0ziKV5kaqXEtJoKCADbvZ9hNfw+qA4GeHj6SXM+APtSoINPAbU+bxaBJyknJKv7x
493rXu9PNh6xUOCU/Q10RxokXgA5XSU3V22wQimc6dge2dDpnNHTQvUaao0QX3lEfWRLJ/Kt3zwn
qMYSGfomaP4lPJlGLlOPBAO6p6AtI3wMQre+3+9qAToYiNag/ys7c5dIV0n38lzZ2SjRWKMz45/b
9CJ5Q2ij7bFM1MeIbrxK0fMxCV6phSCT3hj4Yd6KU2F1WMnjAfxeMpWZpUP6Uz7U01jY2OBtb4iM
u+C5dB1fJ64scpk/qcoFVN2QrmeTKJjqdwEfXtqlNkHo9sKMpE4NS4CtRK4fJah73/SB3bTX8nOd
AgLfyuW1bpyezOuj7BbZbEbT/4/8ZLtCc1ws9f/9QNKogMu6JvyEXQep9v/XDfZgopI3YXFikBvt
NxLgNo3scr5/0as5kK3f4y+9EEyXOkIvydCtXWoW1vgf+1VIIcXaV4xZwt43VV9BengdQP/soCcb
vrSICydwMAYGjxlTiNeM0REhnCbkCc0rA8ZBVArKxVfbyN1DTA9bOdbB4sGDj7rDzzz7fikPscJE
PIuItXPc8RNtjVMMg7a+6QmLDc9UfrwFsDHvgt+LXBX+brQMCIsnd2XG0YOHdQccBQzUNbtF7Dfv
Ja7miH+0qi0iIbrXJQ8pw4Plqc4qY+/SCVu7je+5vogTTBHPd45TAf6rXB9rolbEOarMkj+ja/1q
a8nF0/q4Dh8dEBGPZNy3tCuqu1neX9gCSfAIa5K9U1aX5sFt1lc7YmQ5MZeHvVn2KK1ABYm7EhGq
K+io+zVtH52bQhiQL2sbwkq5TRWtx+fvJ6H5BKMXCymDtVk0kyxhwuycSfrQcofoBZpwUXZiDBy2
071OS2wH3HktRYsjBnFzCzWLNmsY9Cr1m7aUsKONO28PPOL996f3gTFHIujfsLaaVO8nthXRmhHK
xKUUasRttkXM6oumwdiAE6xEUsY+i2W1rr/UuXRGOTBsd+V8Jn8P1M0XLlDKriFqhn5593NqMNbc
2jqeWrJnAhAMzNOAC8CMd/gaMNjWpmpxp1MFHEKdNM/+EZ3tcGP932U1MVD2ktaAE2ZX2LJKrakb
M+s1JQIv5zSkTApcSkY40/gy2eUMrHZ1MyWw50UIQ4XXrCh1BApC+Nozd2Ytc+Wso+ohv7v3qypU
uGA76fBIzcuqXHBVTQgsFYSUfKe1t0F166bnQEwYbIJNb2vMLckMqX+YUeBwpwRMQsR+tqUVh0q8
3FxwIAg5CdqsyPfVbrsE8ld1uP8Sb8KbyKLQ3BKQmBNllxPNxHlHhD8kyAAtFN583CWj6xKdkMh9
P9lXB+2pkbCj8hPKqdBSffXgbxSqVCmRhRWTTObyY4vlWo+rjUmmQqsoUIjcFtvpfipg3YQHe8pE
ZadUk9dT3WXlGWIImcAhFY5Gqh9VSAXM5unWXmFeGJnRv+VmhUtBpwTAOZSObxs/llWwnlnb0WKs
tHrvOQOZekSzAueeupClKrBXObzBdl/tFXshJilV7UKcKJe13YG4myHrMHdqTNwMWzmwkcg2JlLJ
RyrfscPbczW+1abdgY43tHTBDIA3xPBIhLsBhhm29/wisG4AdBobMVgbCdpXh7HtyLIGIsQJrgyb
rEx5JZYr/bfSMCQPsorq4Tg2ZB1YqVT2zxIltbRzaqGc/YjtN3ZET4uPWRobsDz59WgA9SR9PN97
HD5qAmuZ0XZxKawW0T9T/Em0GlV9U87v1O8mKb7CDJBNsdEoVEl0Cb/KTMrKyh2vCTQbZ0gomgaf
GTCvd2JwozR0pLI8z5Te8dxFvplwxj5plWTHAlRjXq3sXH80cg/1B+wMu6Mxh3wb30Rk8YPYy7YM
gzVk1OCYH0hE09RFY7Zgnzj/rFNTkn/bRb0ludiN3eCDhxvTNwdRjQa10DmEGxYrwhSkB4K3ff83
SZUQpEbLb3KQnHem+r1pmWsIAxtD3ScNfl1qNIqLOeFfGynVo1kjNsN7+n7tNp3D6pAeomVSrbTw
ZLVZw85FJkL/olYfGYZBmwMQu6ZJIo4v4fvfTkc3KUdFjPmCFtpj6H2XV9cS74fuDfdcWizEllYU
U64PzOIT6AyxVNiltYnz9+k0uiFPPo6kEJCiaCVeYejrhmNhVfq3QSbHS4VVqJh49KyqdKAWX6Km
b8SSfRV3IT3Zj7pN81Agf4jNI2ib1/ZAHi73fHFQ7WiwTF7cAWNninyYlQgO6K+OUIWqgQsQxDor
9Zm0o7EPP1o1sw9kE5mHvUqXqp5ocILnQuW9qhwDcjLdfutNKF6s2iWggGy8VWAZK64XVK3F85K9
7HAc4mys8Lkdzy+HZVbDLx3UPIQ2PalcabZmeQSkU0FucgHXYufqluko5pbvJusmYgMTVmZ5PJVC
yfuh6CLhqFlHCJ6ldQrRvZ26QikTevocwOqiMq+erAVSyhtYXW/7WHVlu0GioiEGQflJLM+ILTRb
eT1bFex8hjxH2OJqYaqtCn1X/jW0nfl0upCuROj9w2CRpQ9EljXyW7BjpZsMwpvy9EPT0TVdwDmx
YhOmGKRk7rBqdK3P5Fa2dW8JFKdPnMovECGfxLkOxetf3Doejk1mzOR8HP3XItU8pOfMiLBpX+M8
R5WGQc+a+paukNJVHdNFmt/PZxslxxk208gifmUowzn9sqTA++ONsb6nXGEM8nPCjEUMmF2hil3x
Q6mdWKZJbI1FTHi54gVWIlKXlf3lXtq7vZd/XRKWXrym7tGMgC2twtWrtom+hqsGOGF+dPzfw8TP
yArtgOKzyouGKhhjBMvherWBIkS3siO+WSz8T663bBaBFd9s+zmoxsA+JrHY2IRY8Qer2PJoSgBa
N+/CDutnFFLyjvF1JHFsMbRgpRsLEfjOx8IxkdaqPaEatZVk08Vie/+hh8QFuqnGLSymW9toyp9R
G4F7wfEuMOdugNsNH9h4+iyWP3ovczG8bryufoDNWZ9X9FPixSUjC1TnkDznpRdZBQbq9qTOGcUV
RBwLFQbthl1HDXeuADQzFZWc5ZmsmiClyFdNThAvFG5dK4MCfSO7Znd/gzrrFpYDLL1n8t4Hjuz2
hFgrTltNmO5LPSLZ4nWtX751tHxOgvj/f6XPOf8hgKotF5fkCfxcu/AqGFUcWPm9AYpQclaxUhix
xQuKaBfFiPoyu2CY/U7OI+9cy2svJNqvNu8RjIYk+VTZLuqZJemC9NXTjAl87nzFz9OyUzdcJNy8
fNL1HVVgY3k0YgU0+tI04XtwgJ/8Ez3Lo0sbwsIolitx9fRuHdnowFeZI5En/p5yZtgV8z2FXPE0
3g6oyRAgNAslPOeU1yD4d1pKkcXYoKpbiZDDqH8gWfct4vvI2rxHE3fDkPbGaJNqjYgLOrxzIqzP
CXfwC8Crb/m37PBvXX9FhvkpJ8PxZaVgGuCyw6B6R7JksAWnE47z4FNtrn9iWMh8PN2j9tXvCqvT
BuWJzuyJuIJVgH+gMXwZ/VGRAbJLY1M9HVeOoS6r0R7kkAAP2aXMEbBEFglQrofa8EoLvVBgiKtu
KfZzRGOYY1C8urp1HgssCLsom9HRsZj8NZ8ri6BCmvz8HiunuJOocAu/0u11jIn7hSxwu8vPRc0r
5tEX+MBbgDhouVrYQFWzGt0hxapdTWAptSMILGYTgJ0AhuqBZxS868oejr1L9Oxdm7jOCKnKpHI3
ke+3aMa3cQ7P3IssxqIDsvriHm6747pOGcy+qSWDofo/9iBMpj/WH0Rf8/I9s3ov0tbzE0ZL8zH1
/FKsm3eOb2XyQea47nu59Ujh8i2Yllmm/5XT/1TCmmU6vJ9iRPhsktP2ZJJI3pHS/hIXYwkMvkeG
I21y7NWCB5rIKnz+Sy+0SKoR/RFtPnHdzR2V78DjMwNzp/oOXbXM9cWMeDDs/eog56VqFrdTAMFD
EY15dr/Ltweo0mPqQ6x7HOOvdAzLNYRzeSQ4mN0xJvAXdVjKTVEMCyWmwPo6cqYgm8GUOsRa9pDD
Eo9Dfk3wmP6u3xf8/4r8SlY6EXE+sGtBMqvOvpdgddPZ+Cp8hdV0PmZ80C7RR6AdCOAghmVKIv6S
YdoAs0MHGhoTX/BvOBu1BxBdwrSK057epS/Kh0+q67Xgkbhf8EL4rtzKAv2QoVhTI+g2lpz+f0SF
PN8KW+X1LcoxuNGgDEk/NYuYhRIjh+ZrO2T7XJNXC5Szb60Z0YVciQ6tf5YCux+XpM34sP6tg9RQ
DAhnWCgVE/O0bEwGHK0Hm98pF6x57a0rn3lRXp0jGm6E15BOzOo4afozxBe+HG5unhYntyJvXBR6
21KP12FgTNNCwvYVJxyuSs1bFB/qwD8jXFdppwrEQdn7qFFwj62ygckBr3iL/ae7hDrouW5aggEv
Wvf0STTj+A3C7HATHjT0y1suebNAoq35ash+5qsl4mb2189JpUsISovK70369QMCMq+wt4MVl5yD
tyu7GeMK/TqDjQMe3oYzz2rAsrmaQZ0CkrVZheNaRMWl+0tzAmGS4bqVJx3XCPsTp0sA4tKI2VfL
w7sYcbRrzzPM/4ok9Qb0EyZfn3Jr6UWBuy2wgv7XNictqEYXDfQSvm6k+Ls7ioawnmpFQ3M6NC02
878368LYYadNIC9YwmsclypSrq2dkBhkaNIdJwf29NgFtuyhErc6o1rK4ISNlzQ2htBkimdlIEl+
PtlVRWgczSMZrurTGsLfHmixFIaHanGb7cUJ7DcuK6ELK4UUtfr8ndhU8ADtm8euy78haSa8Wa04
qbdtiwFAryBvoeLM/FSlDPP0HMzSdo+pRYf0qLvvALED0IVdP2l42ZYtyHNzk+JMs8y/Kd+r+q1t
6Mbr1RVEI8A4TNkgI+hcBDt73t3wxh94yaZqxzcTl9f+MFTIHD+H+YH3Q+XwAyGhzFaXIMJHMNRD
iGJw0HYCaqxaA4RoVkCKWS0o+BvaJ0vk42aO0LwjQq6MDPR/iGkHFWC82GEIM5fFKCCteZm8L2hT
6Y/9OUzUf6GPsTOk9tgPy38fx/LvByuuGQ8FReyVXlI/Js+KBY7fupsSbqGnoDPjr+V356o1xHRr
Ui92HzI4gdR4JnHWsZGzsVLwPAZdbksvq0/R4txMS+i6G1REcw0W/CUaCSZuue6acuQ/te9hwcLF
g6NxOxhE9sQNB+uQHuafBu+OcIoUG8rfQJdDnYKB+xgUoJM2N0Dw865TykOZv9fxyevH/fgdIWUh
hl5uUDNiSmfB8GbcgWxTSQlJSXZ4rea8mV0clZ2tL2/jbYyiQrdpImuMyzAc0Oz5Wb4ZyhRgrqoz
l6BFrhqTJNX9MmWVdmvmzkFezT4ImDVoU3U9CTLwnB/jMOqL69rkAuyQDQMm689FI85BNn6BFzb/
lPV0x3nQcDKOKV6a/5XT71tSD9ejiGZIfEikKb4aGTIArjhoSZXrwWAm8sBzxcPhtNUNafjci9ig
P5mtRVLPG9jipuO65Ng7N2DZzmJwE/VM3dD/xZexgZUmY+k57LSycKsir0RQNofeTHgnBmuFoJO2
y3x0OAhxAUdJ/Yk/0SPa9riceUWYkes/OEW4zCz1D3WtCS3ILQfv0RAQnzuE4qHTzHZjyj1PFdpn
9Vs1o/ogwlrC+UONFU6zu3kwxUI8uRcMpQXNsvI4oOpun6bT2DQd3R9aAhmYqUYqAR7ZDVeM9Jne
gT5Hwzh8V2y0PzuX2BlJ/HeF2feuPCUcPXqKtO+BHZ8uW7+ZpSGfgOdZ+zBuSUOru7JT/mCW07J7
DAphPf4UkrDFIv/dIwyxY2DjjO8Et/uUdv1i5rtR+Lor2siXWo9R5Lj7+YmxCbqtCN0RHaaSS4NH
Ifd5e/7peVYPRpk8kWY8BSBSDXd//ya3IrWUj81dpAfh8DOWkMymWdJf+ePOh3jFB15cjsFGeyIz
AZ6XflFMs9Lg6qfF+hPbv6ha0CXQMHXqVLZntr9g2+eUVYbXZvA8eWODbH5MvCiZpltacdBgy01I
lSIN6GgZzjmFlciFlZLmQ07HkypG3s7dZk34wMfGiuZKxL6cJl3ugjloqiEO9jaiHyBZc1LBTuJv
Loeb1i5SBnkK9Iphj/ZyCvuaAGk8UkTlSkyPSZHPD0wkTNv6njldXHAVbURdbpo35Hs0A29KnlTo
g29ATWD14rGUo6yJHj5kI0Vx3vFbFNWtzJGFWpJxVYSm9OynSnfoFv/2REg+lH0FD0M6qvAWHRgk
7blnd7UX6AcZ1b6m0q1B5l6rL2icdEXWjjSpU6vxnHLM/nWC8pdTDmobZB5C6axzNBSgEqAnVlyb
wVfrynOWS4oERUvS1mVVf1XTTFDA0NpB2UrvVigFsT6w0LWb/kd5QKS84yucANI8rUNLEEroBYMD
OiW3U8rvG+rwIP1bEh1R4lw1YFEdfzi4mqtE1t62iR5bDkAh9IGx1428yvkEEIV1TQZqxuCJAHEp
uvNGkNhK0B+wPwNiQqEOpEX2Vpko8xdq93DGFsvpxbkYfNyZre0VoZAuR+qbuyz2Jo+bDsYfJoor
1K+8HXR72E8hWLc6j0YqBUp7i4IMVpD1LaqErtm8KYasYDo4bv1CikWgNGLwEsFnIMKYPM+74xNy
LwInTe02joAlnbqfuwG62ghZ0bWFuY1rCtcOMNFvNFxPnt7pZIzc6PeruLDNmEcwm10OGm1IAAIM
3mwrNEcWrn6hdpN9BalUWO7TjW24RLrmjIodvyMfz8a5owWCH0eQTCTyDLB7mnp2t5Gqeayc9gaA
N+9i6cfNBwJd/BUuh3wTvFN6wVdT5K1/IY27T5qKJjmm+8MCz+nYXudVF8RK8mrwivLPAVQz51j4
HKgwUU2IlbhPpVUF2ZcIhYlHt/+6usva92NXax0oRnt2OHwjhU/AJQEy5cAZ3LrjeUmnGtJTraaE
MPmWZzaWp5XZ5sRChvuChD2vtIbSKfwzCCqDd9GiYb8KlNPjLSI3JenIp54KVJDq+Zhuvk4E8Tr7
snpY3yIu/ELgXLgtcVgyBs/uRdP7hhK5NlQA58ddB36ELf3huXlJ/M5SO6os8EJpnTrfwymzg1k7
eZjTPUjBPcYaanmxtAQETb4V8EFej8wBf9+Vg/OgQKo3IriBC1EVnL4J0WYoYiqwF8DfRPIm43J8
91jWITUvuU8rzR2v2CDqSnCPd9VHb1RG4rrhgttAGioJJnAGnpjAJ60HWlUUku9ajtdPm5A0eDDT
ie74Wrj2HRbCnD2tnwU3sCmYYVHQz8r3qRKwegFwxB/d4/tAKgupna74lO5fDz1wRRLf1GgvxLkR
65+mx3umNxmomooByXUM1UgVFTFQS42a4A5TW0c6tAddt2xW3jQ3VqeXcI0d4Yfgh2x5yR1yUCAd
0PF2gxMdNptvmmj+vGCaxzDx1IO/8dpxOZXi91B70gfXixuvLReMFKTSG1xvvE5J9ZWm5B4EbX6H
jM5kv5pRLr76rSHXpvxqgO1ojWL0RP8jKqpnuFEujeDHqjfQosYppyMLYo0l82vH/TfnPCO2OFbI
03ywnt5Z4eFJdOGPiMKiC9M6JKkqBidEen6kS9uJ2y7gY85UyE+LzkVYGgw+I1I8XQXGhNuNWn3k
JzvVW7O0W1BDIVOgjuhi7GHYhZgshXotmLov9p+7o7WwfC/EdAUQPsS3+nBuP7W+j9QgkxU8DGT/
XcthLJl2//4tQTl6oIw778tlLmRpmEX6TiFCa806gW9YG3S+inUNVFDDKugU9thmLMFPsO4HFlGx
eDLe8Gyfc+IVSSWh8HFvkaJBJsQeHX8FFezFbF8vL8gc8ShnC3+1hi1Mfg0nn2aS/0pIFGrkXHyB
344VcYExyfO/PtFlUvIPet/48Cx+GD1AwSan9DxghRgIVexPTIaqUthqsebzQ5Rz1Bzt88xjN2Iv
JuTS5oRfojrX7zQtD2saIPSi14Af8apJwZg7fh8L9VifHDFH/BF3QHSf889Caho9sOZrReGN2t5p
dRaQbUf+WSOR8miivl9fn4QfH4NMgWUKoVG7yoZPDpAdQ8Nez9PA0sfFuJrRhvtclWV8/QV4PPd0
LJem3gttykjISpbUwqc1/nVDcNfxhaxSdTEjetTLZD7j+x7FBDVKri37T55NMMDKy1RED5BA9eEP
5CehATV0oys89BLyLEzY445qOBGfa7zdrQg3ukmqI1AYj/ZdRcHzsF0aRD720HczFbLENp8u9Mw+
Dgalhu1/AjtOFSk+sYAPaidj7E8sC5cRzqe1wtgVGg342yo22SDj89BKrsO+Z8aTUfgSIqnquan3
O3r88L3tWIt5iVmVSokAa1qPHrr7wVXL0qOBDuKT9JV36utnBUDusOhgYz4xFRpyOrnbEFOoFBrp
BG5vBR6Uvb0A0UddIA90jVeIUNNcpruguTmX7XiKfNQHMAabCg8ghRmbwATNACBNg+VmYPUVXprm
+80PM21tVdpFVigrRrApgnbaQVexEtyPPHnUzB3GVVL/uhX+UhfoIuYkVhf2js/Gq0noLSbd4UIo
4HFjc5QdDWREU7ag+KblPhni8tlhksmDwc7n7vyiOVvubswLXohGJ4CgfShIl+SOFrKQiA7iD/Hd
JXFPb//XW/eN4pQD1dl4YnF7PwCCfibuc5ecqYB4TPF9ur7h8kqlX7EtYE1V+tU9geJdcBUkrTfg
3MMaO5ib+kKGqAZT8UXT1rGi4ZpqkmQGgjLSVSlDQn8lgd30vEf27CESF1EHj5G/CBPfXJhTHa4a
Vcba2i4R5CAf0m5F3/h+h6Zcrqwba1ZVhHhIOKO4Z9vHONJ31JkPHXVHkRrOA4k+SHDMNms6sgOo
SpQ4eIfHOOH3+95juey3TGJHpTruVtorR42fk+90DqA/Ph+mCguElwdMJ6g2Vfw3AYaSQGXNcq45
i0zlSKviOaXRJwnE9txB227rBdlBwroOjewlvOCLp0uaJR/tXxsgZKF2DJCvUvmMatrfw9wQetWN
RnF4MrSE5ifdqUlGiIfofE22OZ0vRKYmEfpmMAzRNkklncYWGlksipEuACiS4Nn+ct3+91pqmscO
hQCGs96qxDZTm3qEVykf5qw58zCf98phg4LwBBh6+4HS5yYhktV731CICV7C5XDrckfMuGbk9GZa
lh1szwr7dim9yqWf/uVq3V8hxIDWMf1GLzxijc3kE0dGiq3yoQsPQ6CRHmhW/xRAloI+djKOmPeA
weQdCfWSc5RNM+uPJu3hv3ubummfDdXmvQZH4r7YIvIWxQ1mWv0H/C7SOeHqtGLJ6GWBkD/BPZag
qy2tHVYEztURk3+H12WLI3VpaaqNddJbTr6TGioTJPbIFeHRU1dGx6eAcJ3T7vIyGkUMIgc5CdCT
b798ZJLKd91eKwVyn7gb3gFzQbByC7C6XAbXxUWSTve9mvmW1ymMBfe8fxKmZ2jsfvQXIMiUQ7NP
VcvsLlHKXJqNCopUtQR1Fu6MkS/rKsSZczpUEA0Gb456XHbbshNWyHTcedsBuAUz4UShf5JfVCgu
kV/4qDVeoXhPoP/rtm9UjwU3h3FZpQmTEja992YMUhnSEE/hDLvJcrlaLNKTzThI2cuwqLe/OzY7
3JJ3fLZ5VxlVFoT3EVuhy2J/nxst/JL5vOZLEKrjVs9hjto+nngAna9SUzWbxD/pmAccZa0b5scD
9W9dxzhxe55cYXQZt9Or+anIKmS00eCJU5dzVUz9Y6KAOlvz1u/2eaUcipXeOuvLWz2BZ43D5t6k
qbzynJyRrebfN88b+ucdTi9RHlbTs5LMPw+vRSOZ5EVWF92X+Y389a83laLaL5nCJuf2gNOJs0M+
uA1HhuCMNQD1AJ13agWjMRYIZlii9kgQM3tvRvS/EWXMrdGBzRtSDfx9PVOht/cvWT3Aup6Q6qER
2XWTUfHe4CZ1IOmhqzEKlhM9QYDgNDRCyS8A3Qm2gprh38F+syK0uQ/ERB/zrI90XKUoqPW0/qe9
9Wv5J7kw5NaH75x1+DxeEP1fQeS9/OrZp8cBNGl4swavsPXhD5bH5IcQ0F3h2SXlxDKmCXY2sEBU
oGWtThymgBR4U0e6PH2piYULdWmvJ00UIHHauN9HENfez++xZIBea8Md8/WJid2OaynJifrLS3cW
WNGobZfCmcBCOremHZwcAmJh2LVSdbxDGnebOHqGQyxRrC32fFwciVV6cw450soenurt2vKdMdXr
Hnidq+6vKRvf16X2yms+rS1UORZxCGQxrOCQ9/z/KsGJa2i0pxL4/pyrOOw5UyB3te9LubN2Uug2
RaFcWJWH+eU2qIo8ZwkdP1vyXjQiX9z9/Zzg802KT6jTK/OBxUnwGOKPWWNcWAHxQaGIwqV9RS0z
fQRNNVH/kgGnowubBI2gF4oWpQcbl+9X6NPtV/0Tp2ebwHL+dVnxbdEhFcHLERgyzsSj9wfEy3RZ
E6NWm/gSSRJ8B6WUxBHSAADjsP8P7nj/MgXahS3cC5RSQTUE7bHzJt+WgVr/VlbyMlf0mK1Ky0nU
grajjB5vELKvz8OJUcRZvtDEJHKSq6cqbmMBjDjciEmzO49fJFVLxlpTDqKTVsGJcOtTYf/idTWk
tPDP30YEBYdi8r7bpb4Di2j0x18eAIEgrLWNNTJAXII03w0KRhFpqCqq3v2Mpe3y48uV5tBJvCQk
QDX4KEBTEDvQSLKMF49nG5WljUH6NJ0RubL9DRBDJTH5yUkt4nZnrtWceM74plEoeHWQHRzJ7BPn
aPRDL+dMg72TmnzbVb1mEfR1hZPKXK9QKMO9ByoEm7xBTOfHwt7N6V092g9ys2ZUJEERRff+AubL
KnJO3McKJw6jFYUG0m2sCbOsnKh9lWJsVXoAy4B127/p4LIlwSLJaz3TT4wy72m7l9imcAEQZr2Z
YxyLVuFTTiE3dEFTDOX5cM689b7IpnzGOICFFplpn98C1GuOHgV8VCjw+RwJOkbrChUF95rq9tsr
ffPyBwzbgGXu8N7CiuxRMFOIZmGeRoZOTJO0NM+Bj5ANutnJRFXWGjbJy0gw80rezv9WgnbYIAB5
y1eCrtn7su7/p+RkwQtaUJ+4QklhxaDD7EzNUIatmFJeTktIx72kDVEwY82ryZqmC7cdU4eLP5R/
szJ5gmXkvx1myu5AnRq5bEnFqGsYfQ5InK8TkXpJh0liNRY9AEh2wzQ8UbYK8T1/w83pWxgcZD8l
byZBsNcr4oam+Gt5k819WNUPSHvP3ltTD+CGD1AeUxeDvDlnj8T94pxJRDvwILTC4jVTLyDz+/AT
Cd4WB679vhLDlUNR8++P5RA5Xle7j8PLXcjG6/r9f8fn0Asuu4X0PQwJF7qGouwwO57yGqfDMciX
gGEBBLr4iqqXJnz9DdjxI7NmxhfyVAD9gaO0J5n9blF6lqWoX+waepUVDbaoI8u1uwLIBkCnYyLl
gVFVxa1kbTDxKZ8JcZTdbe4qG5q44RiLBl51CLt31kFtoIPoC6fqeysk1peWrlK2J6vmdzdMVOhF
fGGX2U8ADAAhZHjA5AnkP5aDl+wfeWkHfQMvhuXhFT94JIDlxPM3FSQNU/xWjB84G6u6yb9KKPqE
kmZBKZifriiyh4hVqFuTL5ww7KgsJVQ58DjpAQJ88H7jwZyVDyOueGzv5+mb+EHN6QXVcZoVH6/m
P6Gv0kHrjqm+XFP6+5xDEq7TleGXe7qO/1KNYAeDVO80iGnejgh2f2+87Bqs3w75+zQ4eta7sxLO
OLKGFnHGTlSxleIP0snj9NEamBy1g8iWnW+SZQI+gOqPilPWNzA8q7TYy8gvZiOqUQOfN1Lnzu+Q
O7Buejdb6q3BJbK9zZISZ3G9xgpmSWIOxdOwCf1j8+cllDg69stIWLRfa8o9k2XzrBjYEDN8hh3i
FSloraUV33kRTIl3+5xBaIkOy6Og9YjSByTxCEDT+USr9RwviIBq8Ml1Xgs0ORreEAuhilHoqjNP
pxyIuw6+TP4/kiifV9oCZoFWnjwL0D5OvFG7enBJ8RSD4aPiwkMzrbeEi7sdVlIW0fJUctQLMBUx
uvnh07cU3i/4MekpmL+rf+muGDb24B3VQB9pRByqDqv+rCl6zZ1XOxRo701FQoEjIrt3B5PJvh/F
oRyYoAW3psgZ3Yzw5QL+1C+AtrRPhNgCPcGhDR6aL8cXsF5oCp9+Z+HOnAkb1e1FkRiB3Xsgjpln
3UTpEAVMiqeeHc0HHPpzec0vHIBdmnZiYIT5UzR3H/Hw8NqedqJx2sxhqyvMU2hx+ag1uR1wdijO
aBN5p/iXlj//gWhmAP+1eqXKz4yXnbwHONlYwbp3ZjObbAi8yiEquecS1QwdqOTEVoFMVSxoJ70k
9zhZaHV38pBqctlbC09kiXHjcLrZB3VzCUCMQbXUArInCWvCxQLNE6MV2RSs6F1mBmyGgoxdthEO
Hn+riC+AqLpD3VDo6WKceubWFoRSEMnOpPSZq3u1B/nBDQUrVEyiqWK0SbLPxrQt7FIycmDzyNX/
lPNeUgWf5o9qAAGD4lPXsfYHknvc7f4hdvUYABXoRASA1piczHZWI3MBTFzCE5eCwTuZ9odRYm9p
jurH18IrL65RFVMQHBHrh2wNUwFs01kl8BAb304j78D1H898PWngK0JCcEtFEklnLhKLaHov0LEq
C14gomaEzzVDV1ENjjgJsZoGdCA5lhege8lo1qeBKFClh76B0iuOJAXIrsLTWlD1W5V4KagZeEpx
RUwz+n3vsVe/u1t5ejDb+vxF2kqXO+1Oy6Kg/AGSw+eTvtaEIJ4yGHgyQ4X90sjOqQ2VdhiEVyu1
AC7RTlywEsIBIMv3WR4CD3ndvgITgYdKb8HILlCqsmNwSBpFVEwRji/4zPjZwX74jpVoLTMXRz3F
06QEgCBBIu0Wtb0LFu8hyWmFTeb1vpHFdX5cL6rlaljmX+vnROJP9y3/wzPVr6xu3jJWb5qPcQOV
GPoWJ3cvXOJVjo5jyWnT1kFPLLM2bnAhHb2hokoRu95A8Qlz/2fZUfhmmptOvbdW9a7b9F8YZN/0
1nnc0qKgZuwxa3szwgznHTR/4yP0cZS6jTjdyNG2nFxFjF3p4qGPkuR844ST/S4DJO56DH8AF5Kj
f1sYwmxHC00vpoLdklWnUbsr0c4uDCUFfb7itOuouxB/NwQ1O7Hrr+4QYJNEZNPPHocjIKbSOouT
wgX6QHqSao41BnZ0WbM47fKwVG3kEJGZPaAfqO0JuuSvvpicvwhR0hY24tkdfmaooI8k4ifFZVr2
AJSGxgXDclaFvsSxXGV0LwA0nlNAmFSmECxidEG+A8W/Z9zDlXamVWJDnw9zkQUPA5VIaC7m5zVh
bMEeCrLjFGJ4Yjckkuvg37hiqohAYB+bddaaa9kvI+0htag7f36Sbg3mgZmDBHUCzK29fACMglWh
SQ45HQ8UkDaja/zAoloEgy5A/xP+auFrNeRP8L0rirn3li2VfTezgKPDTzo6jAEOz3WXn410O7Wp
eVNt5n+hfknBxgPDWxXB2EkmnnPWCuVGlcQ9wIxqAekBcKjt6kjYkOfGPDwspAbY3cTWfW6TCb2d
bzcijjBJhfur0hR7JMMPVoJ91fQpDmdqGPie/zlJcFBxCXs/IoIMi+66BVOvjEJ4KpWWkCDOWTX/
IPYlJEDDZ+8LZoBNGC/W5I+MtPYwsmXz7+nYhynfJ9vf2JJ7F/x2sgUCKlfFcAnkiC8Hs2ay4QCH
xlpqei2LtVDyUcPvyRr3+mO1LR95nY1Jt0XM2ZmgZUCcFLrfgvpvOCjTTmMtyE0091LOdWc5/9RN
wOPRvsM3CJTvJ/qST+LD6YMDq47OWuuedAqEP1OQ/+EBYCm3J32rgWcv0DayI6jWP7S1uhWfOgUZ
zIHsrER0YIAuA7KmluE3RCjOXOesIHc/NAwj9esnSMC617AeoMGvQLmFPZeD0bZz751O2hhrovFX
XgaX6CpduQzxjk1E8nvWYO47FPum6JS2jun0HZczbq59yYPXNjXnNixr9Q1aRF517LRwUiJ9f/D9
213jXylK3FCCeixesZi+pzf3nHmn6svswUplBs1H94I8GWEPebJ+wbn8reMQt4fAG7rbKQIg19Mk
Q4Uj+rL9ru+edxhVCGDaQHtuvD9PbZuWGHbqGX2c334dcR5a1ACz/3MNnNZoCbPihRE5Xg/4e2bp
wTHBhjMEHGQJQDA8A061dM7pXjl+W74hQ7XRGXiom/ShoVlErYWhDMZ3hpLkqwlKtxjfECk1JZVt
TTX7Fxg8ZdGi9xY0AzJe4pJupn3W7iyKFxsC+qsuJ0iUfIjFUKCn0BxjkRLqrc7mQBpudUZJjTaP
khnJjFoUqOrtamwjGtcR6U65nqEor2LnX3lTnc1w5B8wv7NGG0ptn0nY8B/UlORK4A+byt4+2DtY
LmSIeA8Tun59/Ya6QHTHAMtwaKYpZikti1R9XJLmz003Ta+UIsUEJBb+FiJoudUfoDKPxtnAfAmF
ZPknapNdt0KNq9k78l/ZYCgjGzycokt/qqp8C9IzuPg/NokXRD7R6uVTMvdqPHmQ4YW+pZRtjDH4
CEpgO9p7JhB6Vz19QU/EEvQk3ECRb4jpKpjdFJ9Jw8LeQdAdVmGWw+Uz1bcyK0Z2gfy8dC3iP38e
ERFcYjkYsMcal3sxqUgrllti+jEfH4DxLw82SXYrahH6wY3oWkGtFTPDdKf2zwi4nMjdjWj29uo2
L5MrMgkfHrxxsFom1jb82QXpgO7Iajel6d+OJUT6ikt9Ywp96F2oVvgPcCCPm+zRpeqdCpcksEO5
Qcqmoy6+Jmf8lDZ68imh4iNKhJKKDk7lzd3NKhxLRblzJPCJAZe611sK4mPt3/9966UjDyK3l5k8
uXGVGT42aKaTGTxmiZThKXDuQ5dpIbthwTBpphDTq9bGxowy/pAodqSsBTZzP9tdk2DDEEUhXAK0
fPVG1EVQJsQkFz8t7MjExr+5SdZwS6c+VCbkeJyob7OSghrQFhFbD3fcI8eTYifQBLVhGjndNqqr
jzUG0r8vSVe3sLLt0BSukK9tI6l4rf/yHkCoXsPE4IG1d7sHmmTFHbBPEgPFZlC+LdIKFHIzBlLf
iPFcwwClCBKQcGBE6kZGbPusLfgqMwQvJt7num51sGyD/QS/7SLaKf9q7p4d4HA5fCIjcMfv2pY1
6zlXRKDUX3Q+kh8kaezf+CypvDIGC4gj0wgz91hIaUJOp5d9j7ePLFJbvY/E2RcLT/87RmAyOoNE
IOUmQELv4/w+If4Xy7179fo1Jg3Ia6Kg7avO9E9e8Gu/W44PJMeiyIzzdtg+0S1wIrceCCRWREaB
2qhDnrzPjtuakqMemIZ+f4tjSus5lRGn5K7q2adtTESMhuG0g/jvmEABUUhXbFs4rk5Q1/SterYH
sMAU2gFNzK3KaBlnndDhJ2nS6+kORuGmyjLvYqpW6AmrhSRd0B5IUvReEUQQg6Vy6aJbwEwr7oem
kjr6LVQ9XfHc5QmioRkEPe+ArC0ySsrczcEgtVUW2O8lUcLaZ17V2QvCFyTYfBJDst5K1Aj+5+1B
0sHzECJ+P+S+GSTu5SyZ8jQ/67iqHpi/fHT73sobmQ7q15f2k/OGMP+08qgt/oiedv+YXkStnMkn
Z1SD4wgMSKn8JefIMCA1AIjeIVKByYwkfPC2ct0hvQj2HoaOFuuBMPt6il7Vytjzlb9Uorw0sWVx
F3MS3YXWIXle2fGgoxrMfUhTYBjr8j1Wj98I4OWr+sr7iOTu2ibDOfHO2kTbUmKEd5ci+PW/e/XE
3XjzrJXhmVAvq9JXTqnCEUT5gJTOfs1rkFoRPzv5jPBVge/r1AmhfwQqGb7Txgn5qaY98BSkG8HV
3lQeCrTnKX5Yfzf1xy56o43AFAiR47TiwOF5Vn6giFPdvBTByIHrMobacMIya36/yHZSxFN8zavw
FbXEdtEN3cbX+yxNCbEylYqjRbkiawueUO5QGmYDnmhLoN1lp9Z3CqoBmzASUG90jJo1RWJ9qiz3
4njTb0s9ZCRQTcKK9sAa39guZ+1UqiO8841SKlahaK4Wjznl51oDJugvSEnvJPPUhQX8iD35DiNv
boj4UJGJQS/U0ueg3UbU4Sz9EEhO1GMCII2LIH73+dwDmNoKybyEBl0j8Qe++pk7EM7ofsNk4Ynt
lIEJIsYUMBtw9X0BjXckmFaMc8FimZsuo6Vi6mulfaL6eu0Ilxgq/taCRfxeFt5+gR+VVlWbBOPG
Fa1gLrcFn9wuWnY3qP3hoSHmwCTU17xplvcqvbEoxVuVx3NIold0scjBXkWuo6EXQqpZH8fbAZ+M
y4iypAdrNKMfU48skJLaM6CJWBzHzpQHsTzH2/MkBE6yxtM4UL8vHXgeaRiR0g18k9mJKp4kjzm0
aMbUd+8WTlqFW6zDhAPS/cV6BwgBMLebpQPx3hyZXGyz5Owrad1IWpz7Pcrqvbq3xDvw0b8J4vt0
V0z6KgdWAYnAZgdhq+84+IuqLq7DvD2x9wrw39z4cyveMqe/5P5HLSD9i89CRCWIpCjQKSY0T+ce
15Pagg5G6XKUBhgF2SSXpFU9nJeFZQqXpgnowrFpf04ImXsH/weO79bQyQk5ABmdQFu37SeA+4vg
hnfqtLai42zLJZ9brmSUQ5uwVYuEogTFRw9JhN0tCLip6dBChi0DzOfLw6DYlbRfag7y3VFBVFU9
oHBgnc6Gh2Zi/+8RLj2Zc6HvtpIVDtXIT5qkmdjIF4+XEEGuKw+WAIKQbPhDcn4NRGSawErSLZJd
JBx2T4JxsXUnFtBVwEJHkyckckcAFb98mhIDtCMBEH98J7PijGWqJG98aVD8NpyG9x2hmp+VvLvQ
twYx/dF12Z3HpzDyow48nKqJohIiYs0iwh98dbXbBqKaDsElYaaLfv8Zg62vgzMb1jPod2UWG9da
Vx0G8XQeLSUZq3KogdZoPqn9yFaDPotGobGA74cI+1ifnq+UJUc2YknEkoIO4fqApo0d1r1ii5hH
2BfDZPBFw9ulVN/3jfHCPxp35LO0xLnnqqInkSXgQ0ymb2sN9ETgygU8JH2u64b/31bF/DF60PCL
Nt9cWtFPjEzRflTECdfSuScoOsBjPpmpaWXpWkjSkucbZ46rYnsJaAmCZd3vc+OcMXiMrv5XgEad
X72n1wPlaPqz+9EtmGje+MirxF1VPnlg/FICHkf15kHs3wQvNmDGyY/d9hoKMs6ilpPJmgSd650k
xw4ik3cv0oVWHCWGj0zhl44jbTblpl3ZEZBlvkP3OoU3Yrw7INDS4PMoyrhQnnNUd7/LaR1BmVwv
B6XFRXurlEWi9p9oMGlOiKpKyLrrLMJysy7rL5ouoiZZe0HYDudwsPQwZ6L5zhTrmbtkatZ+LNnd
s4wOLulu3VPc/zBE6sLDpTXEIbSNfYQOYEY94Rm9BMKr/BlIxGniPgfXGsWtSbpO7fkJy/30CXrL
mWq6CqyhJrb3ZBs19srma5pVmzFf2KZq70+4rarssvbv+htyG+oy76nNSegNpw3YGgWk8Od98qwX
gOSe8ZOz8MgBqpgetcT6HLKgR7wXP/1NTQjQ7BIJjN8lspboWMNDZC5MbwbomQCL5zU+of0aOhse
QclOuhqc08Y4S9EyUy/thx7g+gQnes2h5iA8p42Oww3rIJM7NZtmxWWc8JwcHmAIOVqerOZi9Pl7
ZtZu4TeGNtNAnvRUfHQ0rUalbfuE25Q7vCMH5DGklhPNfmDkHg5PgJrFjijcZStrpe9zntEYjSk2
8HeLG1nvyeTrevmou1yYNqE64l2OFragSlWDgkmDEvTJTkn0fJRxorL1EtFgezH7+h4iQc5R7yAV
oDza/kYmEwGJkADl4bjb/5S7LBMCDnnwwr5wcQ8scRyueZw+Oulnp6OWkZjOAFqKkDPYuosaBbi9
L6mMx+Sj9rUT+gHIoA4NcJMtX5eJ40gqWTAE6U+dQ5AGKKVjIFBv8zR288W5Rpslafx7fodAIlAn
dRGkZs/BpmSOu1KFDRF9yKmUQYFCxXWR+fJb978oLgltLAYUZL1S17JBqqctLvX3RvOV0zmcgApx
uqlRdSuyRtD62JLhO+cdsbOR78tct60gljF4GuM5TgJcNEwQLtHIraNjD/evzhyGbZD3FakQFeii
XBPZAByYWq+nR7Hf7msVDUHQKXcA2T5MB1uCibmPIyK+sK4AFbR3dqSkqc3Ox6Qpiz4ODbA0/TkH
M2UVowI+WL0lTg3RaeXqJ06OwreIHIjWU1A0t+sdR7Tj5a9XJZT1MWhAJP0bSKLjXiLjI5Lo2wen
uoJ30Hi/sNo/bMs7DgHNH4Ej1DaXvyrvQ1u18PSzfDdKbdYIO8TzEFAEWaIn9qu/30V8N3FewwJv
8M9oJHx75lljxyI6gZjPy5OhMLw1wefLM3icPkJSvR5nQr9wbzif0AWs3bcbtdz2E5GILWpZoTOj
th8oXTiUPaTjCrjBGw9wRlM8cTG5b4A5DLfWn8K1siaMzApKJDR2896WsIJDnPY3zF+tbKsmeMPa
F5xbQSwpxfYWLyWQaD5jVfNqsAh0uhhslrWu3xt9uqoV8Jng6BaPgeEPdMZJczBLtdfdA+9KJ9BO
K//795EgpQAMAvTqXtctIljIxniJFdRvydLzKaJYPNDYHpNSMmUCIhbY5CWFdlevkt0wgb0Bwv0y
UJrI13xvdxaeb2HCnozZGcyjBe45j6xn1Yz9fB4WX3f71Vy0GcjUxWxg1DusFNy9E7nKYy3KZ0Vo
ycHUIBoTdA2nbIldaGaL9M88mYtFmZHL/H3Q1ieLLR8etNskV8/D0f/szh+bNCylLJ0QHzQ9vE59
CstiOdsNCHcSsTNrOAKqOMtmhRC0elJuZ6KaJ+7+YUAMcLWGauBSRHpbRSpXv4HJ8V4KDQQGpjjl
9RKkktwCYJjKZ4wevA5scFs4NZhPvV2r6tRISIz7y9ZbKsGS0vguV1e+hVFtdBsIPphOdbhzDuZX
TX5PBSdO9t6kbcL4+WCtW8m+Z0Vh9fgKBwycAQr6OeG9uGZofmXJwnWoDFQc3JP1sgtYsr9DaL7a
NJe9tWCXhLJ5Qx60KVtOn4FYpYPvGgU5vUcnzitCWRXXtwNdu4c9krUN4dp+YNe2Vsm1VLVLMB+x
gKVceaIbvcQ638FiVVQw9OjfjYTWLE2zBoETqhfM4VTM/AHgEwPyMyfFuCImK19ojZ+rXrzmaoHh
uZXCPVonCVfYvsbj+Gk9zf4TcAPfjL9sQ98dLRpXkglP/lPn6U+nR4xy7TSr19ei4qv+5Nps53uW
Sj6HKo67mkX2hrD0bQp7Cc/wBDm+4LLMDSq3CagqrInplPwuwM6XpNTd7IqqwaewCGdL2MMe78gn
jNpp96MEG8zNS+aVL6cutmBV2RQPY2S4kopewSsrH6rezWkaHnFzY2BD9QUa5MY8hPcGFTjsEOc/
+CcZHJGyBeVM1F0tH2lDtwk+c8/OgPJOzO9ZW50LWqBQTw4oamqXCZBWW/oIGRibTx/K1Y3hIjC/
ld76By8pyNUtbveIHC5k2jzIsQZ2MdBcuN7ZhlnnUB6DgInfFRQLzlrwHQlRsCUNBx7dBqI/xpOw
m6D697zeooVtIn79Q2rTcCrOlFWSXb44+I8D+JQrkTKGBIdSJWgSOCXaTfK4k1aI/a7fByOR8smC
vq6o5MVv8SdwKxrkDg48Y2agURSj7+zwKgarvF5pyRSkDOiIRY3s8Ya9dujBt4quCKwYBMZE91eq
+PLa0JLom3YBZzc0VFj1zYso+pPEb1qWV2dZLtnVTPKu9vtJoLJpSDF/SsnNXPm1i84j/3ts54ct
VE1mbBuIUi6E2VcKREW6HqHN7CMVtq40qHluv1g0hfsq4HOjtUZRDG02PmiwJH+gJ2ej8XnNeqVu
xvdOncx4bWSJmzLO7p7Xi2VrqFYh3D05T4LHsgNr2H4vEYc/rqPNUVq7yf+xFFzW/4p+4yM8u8GG
CBEqbDoGtq5LIrvr/z2QEGx/bD8JilmXnaD8bFVtr4XVIOURmrtpJp5YDCzFozyaZNgNze0qe5aS
VJwNjg/zqm70flYrmTaDZ2XftkVd86oJ+xRFHqLJWbc95Vk1WoTq39wefZ6Fjg1vPOVO/gCflPSj
2tfl1VCQ1gScrXINpqu3+aGW1/TK8roj4gzQJm7fMWACRU2Ga4k/b1U5xEuzJBr+oHQ0QC+Fjgeh
7HwD1TwqAuQ50fPrZ1Uzd+ZTBUehuF/NO5SUTnngkJz5GndKcj5nXKUzHX6CuHa1vpnrKF48Y/zw
Igp8Fns3rrw3JSCiB2QdNTg7dzfGGerQgEVKWZIi3Nu4Cp8dyYvyDDJ3yd/dJh0bc2OolsPvKstm
1bqKeUdA3ZSV/KxJahO6QCyU3PAOxZ+otRyi0cxt+MJLvRUHnWFaSrcfAOUV9DGhRJJ07/pIbNTl
KF7nXlXMzAYJrM1MkVUxC8n2Q3CS3pATmgsy6Ay+Wj0P0cVIQZAoXE1ggwRr7YAUAVagCuYXivqf
PjdTMSGSn9dkOIAnA9Pt9DrKtO6f6tIFvMY32AMH012Y4BUeGe4ubWqPsEAALexRFji4Dj8mIn19
g6OTWBC3NXo7g9Hjmpyad+4H9KsZlGriRkPduds0k19BL8QKFAGBROShFM4C/oy2TG56Zfyx4J4B
sAuVUFAImGP1tWUBucm+BbFO5Mv0V0f1lUsrAmVa+0fHZMDv/MeqXFzfwzQ2UISkMUTrnFc5MIVS
acpKZdD0ABqCSwuIxa0CSMTxIDDEcsvDuPfT3FUdrubb5fbVnqr46BmSbCi99v8bGQxuc5m9ZdIv
hoSswGuuPbzoxS2YHYOP6u7DDAm80uPm/MdI5sQoYwubod+TBjLpjekXfwIMd9mhPdgVDkJvxaHH
zfZuF8IvUwysmnJgl9KShzqEY2ERBwMJnnBCbpDOGCCJWbQgSGflBjiqjHk7aQfFOEKsPdp/d0Up
8GkIeCBSMHaqsneHhbjg7J757vI/G6s1+/XcSvjqZuhtJwRa/6Hiekvna7O9u2h7jbEliMI6l6ih
3uuiUaTjb6S9xZD63ZWn0XGe/9WgGTDaiv3Riky46q0BcoXuF+riq++wcpiHLYHC+Zr1m9ifYXki
oTLXFOdIkgHNB/1q9TUtb6R7f9UZgqq4dR1eEb354jcL+1v/94tC3cAwwh9KP6O7UhHORJiGda3I
XuEW7DiC6CuyfmvO+Bcf1wylVibPIZOkiOZMP18E4rW1Pz/fF+tVLZVqpkNireJkeIH7G+DnwGkE
Vgk3+Pj26ZygqjCgEoc6TIn4Xfwy1fJNkJKrYKCS2zvOc4QzJDtGRSRQgDrSkJf4+Yu3/s6A9yaW
ewD8tkWmNIMUoG+FZdLttmqP5/YM701p6Aa9RwloOZt9z08Mv020PczcX8CKdMO+eUe1H5czb0o4
GWs2DNT/ggUoyzhcysnJ0f1lV3qL3rVcJ9zVh49aVXJM576H/DHAvd3zSLfamAUqMl2LEE5KSzhE
LKkFStCr01uz2O69BCUV/xyTLScIbde/rOP1FePmIvo1znhGRXdoc7otVOg5DUXT2RyNNx3iDkyA
ptH3+Yl7co6BhRijTaHXYFlLzstd8hkOvmV66DnE3kK3Gt+OS0XwUpI8lHJnuVIoZBx7NIqq1WUf
OWwNuQYzexWDls8kja/YZu0F/7KAFUj0FxIOvQVPFFrtt7G2tBFTLICRjr89gw+Xq2o+xklbxgWr
Ek8pU3YYcFW/c01TH/Y+I/+auUrxZNTroe8/9HvoW8Sb8QeFtgJ/BQ0/gITC6xQqPunhAPjYVyDm
mkKnw0erVbfMT/HZCxxou2qfxXExTH2jjtrl6Oq1tO8Riv/8ojdG/x3oYqOQIOnL0VCTqBMEUFcp
9atcAKM44JqTPJgwFzlGizMXBO/4q2igUHgyeZmuJj+s8Uju6TwCf/sXJqiSpmlkKZ7CsVlK6Wzh
JFsrZisNdIxyCT5vu7f7MR1+cY4qdrmzuuV5l8hB7N34JeBufwtVEYG0IRNAQf7aoU0sVqz7/T4p
N32XIiq2oEr3Dxr6c+VcZCMr4zrIM3KLVlOoxir9k2Chs6lWMMYeYLcH9B86jqHaV7nYyrCf5cm0
eWAcnSvPnvxjUrImlxcNpBriO/mWuSy56CIG1pAoSGMjPCAEVfXlHjYFIvE2LwRvo4DNZz2hNPxa
R0nL+HCTY5j2cVXr+EYTkeEUV/DxaEcYhfm5qknVUdS4/bfagml9vGhBhzsuP+eXOd1TeWax2Doo
87/fJjqXvOiNR0KJ6WI+hXSk4rNj7WRO05dGkli+KhMwEbILOO0sak6JPly2ssdzKyZcCZll3bGp
pb3RtFyaUrOginHiTBiKKtb5vWiHTuHUWsHKM27G4qmOqTD/SPqyPogNKPV9i9aq9CAq+ZXk/D0O
CXp24ngNvyDkmgICB0KzqDYCysfkyLZahroNXzFwlgc3ux2U0bKjoyobVz+OCjo/OHkq876XUKt4
bnvZGfMbBljR0OlVU22aG1x+rM9S8Wtfsncd/V2dG+ystJwgPtLsN9pwRXPHT+iyV85Gaya37liW
/VDOX7Gk7DgwC+mB/DZSSE+PZTASvwyESIk/3u3xPPvMw4fREethKeCqEFAdpL/iMXpbkLShko6g
KT5rdFpiZuVAeittcA7/90l3oLAPaxtaXRVtmcCQHBnz21sZayjn6NFDPvPExZSn/Q5Mzq/7x74n
8uaWvCYUx6IjdlQ1mq0yKgfh1Ji8XYsgaPhMJckHP2xYovkhKyJxv8ANKoKjTcY/NKrOapqboEij
Mw9GIyJj+JDnAQxZUeabe8fhzMPJXSmWGhJoYzZUvbx/j0RX6Ko0SekBN0ZWnu6eb9Thz+9pL0fG
Z9C4mIXH8wEmdth1fOUBVZDoZyeaw5kxa/VMvVlMRNsy0YbLZ6hm3dO8E+185I7pAvUIAmx6TQMM
h3fNzCSEn5iM7PVb8NglQT/scquaDDz/+cW186OUqlk0MlzAUfQSONIW5DMupN4C4g1iBO2SzEML
WSRNPvYKxM/sculqn+XThHMtR0rdVAXJNNwjgQIj6dCEPd4aSXlBPvnQOWXTXyMp6Rr3RPbQn+M4
f7WSVVRCO8YGeqcLBekq1G49hIwp1t7jekCNhqOPOqrcTMHw/WyUgJJxjF+KioOIcqy/HlJ82/HK
m1/mpyhVg0FhA1hWcIAzgJfQk7LpVwknLLNbvPBDYvuqWRH94ruI7I+XdZWT2lKF91MlBZ5tRxxb
OPp8pPm2rpOYqQcNBLho/lBpVUjFeZDdcwnNZZt3Q+4F0WZE+lE6vi9RQoNfAGQZ2fzTKlLytHKF
f9BVDKSj9MM7cbO4+xMLQ6qVlJjejczXHgZxKo6m8w9KV5CWpVgSytnqxVuHHUu8UXDuFC2EmlP1
bU1eE2AlNWnm9NhI5zXILjkz9MGOTLJvCEVHG+agtfLDEyv0nGyCFSUGuhNJZbf8+W/II8i2pD5z
NrrYdEYjaNJ55OoDhp3Jk93Kl4dju7KrJtbviZ7F6m+GnmgOSlAlWRHPeaCzwVVaXBsoNPf1KRYQ
9zD7/QYk7HVyYMTgX/zs85Dj54s89nyf0UyttIW5geHNPegixS33ViZPavk5oE2hvniOLS5JCmrI
4AltwkRPze5LZTjyk2JAfAbjCTM5qvbQ6Fh+upmu1XFcE/Pjs8ReCzWRl9IQEbzuyk5V2PoAaCeu
HHCQiMrBbwnQVvXvy68jFvcpb98SDk4udSgD0HKg9kKureSomnbwdjca9tGi4+6qNSDQZOHrqjoc
QU2140hAsAiMSH0VICseamjLmTPSNaTKWKimt3UVruOeQCtlAUD2/lcYsMGlvDBtWVfd1DwguapO
svE3RBX0czyCKRqxuxlpHmcfx3Qrjy+YBrtFIJPNtqIDHVwOxJpkojScYtXScuRSjLwgQ2pru9g9
IRg3PAsJgu9j8K49kT0N8z3Nzp8WLULUPyN/7AvHXAHERaJTZHsF2LCv8qK1584/MM5lKCUhImQb
C8U8HsmgEmJMutBMRMin2VWT2T1xDFx6CzkDtQTudCzC9c2UlP5XYF1kDSCj2HWOzuOj5xzUyETn
W+Zy76iSweKfrwVTkqJEGPEwJO/R3ukpbO1t6kx/Ues7f5MYbfZgUjgd5WlHN6d9D43zjp+ZXPbI
gmx1GbOrwTSjo4RbshPsNAEwe+EtfXHa9fKmfZ2SRCq8XEEjtx/r4YuH83Ls/8osZGU46OS9iKVZ
yU3ezD5d1XdI/ErQp2hPrBUXMcOKCsQUrR4p1mIQL+AVbxAEwkAZvi0/597N+hDme8BChmc5RM+B
jzmoLbeJAPLvVCuVc+BvdMWPB/M966EQzOnhqEGaJLjkdBkNGlA/GPLFV3Ex+W2IPFwJJX4DsA07
CMG8jgy75kF8wsbagsHxTux+5bfwE6kxBUN9DpHtMZVSyqSlOyqUEuHUav09CNFDlAXHOGekg5Ut
kTCnuIGJtLb6DWrc5iPPM2GlvaDYdUG2GQAlCmjG62/MP2PCPwX+R6oTzUED8oV27R5LKC7HHga9
iBYgeep5ytujBbvm2PqvvDByn626yPRUd7k+fVt7sIF3m2JeKltRrkp4/EjtyQAp26mYdpnqsIr8
EHMGc6lUyaR2kj8HUR6txJ0+kFgDgkc1ouZeBQpKkfN7aLevbECZ/xhLcvXU/76E4K8+f9NYv3Zy
ezn5DNbSq7GX07sq2ikukzadKogzFdJs/ogQPBLeH/h/y3UWTfxKloq+pn415U4DcCZ/exoqakur
7Vo78iOJJSQpwWf+zlfpwOsT9Z1SlAJaONS2Dx8jIPqDAaoS2B3a9TUbyz4n5gXtYuv1Egqn0Klc
SuaX1yQoqmQ7WifTM5V5+wuwClRaRQN43wChRCvibD9rfJm09B1cvO0+CF3J6tyCE4DhW304VXGN
Vg+Z7ixndquMBIcXjA2zblXV8cPI0AF94UtLfHXCXB89HLWp9QW4LztbNMDD/p7r70tZvzRIsUd3
toJeR2Efj28ogi73IcxUCnm/YTbNYltkCY6CYj+YKTAfCWPTLC5FqMkIVZEiBgbgRBa31E9RNIN7
sct4OXJWkMODyprQ1+ofPUJdWKT8e0FJxgFmlb6E27PP8hC7gTteNRqKvCCCTCnt9JOjff7Z6CTZ
iIuleLsMbgqpYI439T7jh2Halp2aL7Cep0lMtjywilPxaoN+xj88HVgQyjZxfkdtX7y6Vl77kXJp
4NwXqZBjLuJNPx1RIhN9eJ+CYxhaJ3nRw4Cxv2kDATqR+YmkcTe8++7mQUSsDtq5o56HrqibXZd1
Z7FmQQ4QnfBva17rK+on/NoqRcXeBUsybanjM2nTlpaL/eQmOROiO8fNhUjAvx6WIDzbBluy+rJL
fC/UuwrFCM8gjQ1+P+SyDXWNwzO4eHYzbebEvvgDYSw0FM4DhRAHs2Gn24JDmQF5f0qKM/shgUgq
9S15dLVHYDCiYQPU5qvB58rFhz5ihavadlUp3GL0VhHCVopqM+PSrqVvj4XPgDZ8Z3QW2KxRVOPT
mveUJ6QGoLqahcsIegSFWBAORXGfrC6Z9cj0i0Lia900UgQ8BV27Uf6pml+PybOe5oU3GUW+H1qi
qkyfN2SdyJ0wz3gnxu/BYD101BZQRN2QGV4oP4+cHDccSO4TWmZ6WWNuI5wHuKEncsz7jU2LpCCy
AuSfrc+fvhX+Zv6aNseeq/bLSg5Qssma5PY+AKAlupccJOH6FS38NIIu6BBZ2dxEVFOfr59K3Nm0
gtA3biAs8EDFXKrg29kKKk1FclKEee9u/CdaKrmBnXKlXLoeoAoNZq2AWZh82Bt55BTVHtVZ8Y0S
ZQpVpXAzw+x37SwLSOa5NfVY2RrodZumZUApW9qRRO5jsqNfabHEIxJYNS+2PVY2LfokwWztWuaH
kDFSPn+lg0glSml4f4hXw4BrOQoZdTz/6c0kwqBjEg53dyJGyVoM513oaEpLuvQm5oX3Je9WhxBa
UO8KQDsV7mm90e0apEjY34AHXmMnEIuJrql8E3px2bZ5n2AqLyk4fREa8qtGRI8xKrqWeARs/l8Z
HuypDiu4fFAyZmQNalCZSb2Nf2ngUNS57gTATqAZjq4gFOJ8yVyVxU3Yee/rT2+i/v2j0U8uPzrs
TARYwV1EB+bSIanKirqkrh5RfGSi4/8TV6B/5SkXOrWr+TA1Ipt3zSnp0czMKGQpoMzghK1g2eLa
6iNvRQq88TQOj5ik0rs79qS7eSBCebpnzIbFls3iZauKk6Ytx5LjFZyb3rJIgB4W6d4EgPjh/PKr
Wecs5ZTNiQt1SF0Qg+UDJVMyJhovSFOvhWo/KDVorJzeT+QHea6IJTMNGuI62DgcwAzRinxBe0G3
QJ4yJzAozr9l5eiv7CdVuKRr1jczURd8p0KQ1mKe2Tz80RXWZ/kfKpy48yehuswP4udmAoT1zV9R
isocxDBbDqpoXQN1cV83CB5AuSs2LzDERcEASKeMaoVkXNKQ2a22w/UvOQdr2OFlpD4BG0ZGKQDe
aiKS3wsCaJMEeQsqNkmBoroJscDc89aWoF1eoXu8wROozXC5jsUvKnrOduztQgtFB2IJMtSy2D+4
hSG695L3eqLDP4WYYontK9uBDjC/0M1suTy8Wj2o4c8bSddM6Bk5ZWcm64c/de6JFy7iUqAlRLEN
qb0QssF4oN/Mw9pfQTR8hibmjusxzDIxGACxFTJtLXtPG4ltzsiaopPgciMpnyd9RMZM0/rXFNyW
U8Oe+YcMMmM5kfVF6orx1t32twN14JgmzVj0O1PDu63jTtAuCX1kVxJllIefnTng6XYg+/yE3pfE
s1lgSPTVUpyk6PYBJwXyQgyRpMhldZl+lwhRrmDFBp/ic9ZH7S3wpygppi78ndqnJAsEAg2NzfWI
l2S6qgFkrcBfxYr6EJYniXlalh+VBC4qm/HFp1TR67w/OzFVYtYphTHMOzDLJnO/rCfBSKkr662j
+OEL3U5Q853wMclIdGY2tvTAX+uP+rhnjhEU3WQ4j5zWtr04IXch9UFP5g7goSiuHF349t0WFEwY
zk2AUpX9gFbmp5NXPnwaBIqwyHG+BOq5w3d1X45B45GkL4wDIaqc0BkEJWaQS1z3T3ByYpauxUov
v1CARqYv8gYxmo3bM20a/MKVR+enJUrJw+R9NVmIWqLp+NLKWALGajjPuEq+uDz/LmgVr5391Jf2
axsmI95mXgrAdVSAmYqWEkTqxWdnQVIvEtZCMEvq4OSvCBJgxlfI3a/aAIHA5AYRo1YQE5XbAq0D
Xef/OhWl1J26mG/yKicznJJfQK97fMSrsGyMhcA4qiJ5/v5NW6LLLz/KIE2uC0uLPWAWk0nXME0X
ezku/hFldwzHcelhQoFLUMWHcZCrS4AilQLdlbtgg0KlbW9BLvteAItqvThtWkfa4QgMi8gwNy83
cKkIGCQpNyHDk9eaiA0Cwp7tF8WuGqcT9PLdHlmH6QVtsRz7WOFL2HIFm43oJypQN0lJw1saZb5t
C1W3o5wocqsfL1G7LcBCEM1ABwZzFN7uOSyiWOM4w2LT4r5JKw3x2fYoseXopQYQ38XrE1vn1JrC
W+xNPt03y0qKc6WrJWQ92E9h7Xgxk7noz7SQnvo4nHDvs2KOm1xen7sDw4BOtN6ONeQiVxQ9tLnC
AbbRniRRmyu3+5ICWy7UKDkqt2w3fGLHYadzmnmP2y6nExWSIz+SqhtbzgecJpPIK57/U4hss4zd
aa4HLub572mEz6w5NXmqFoklGyTts9kmMP1T+QIM8oX5CaTnwpS4R/+MkI59uBRkx3eGDBhB+3+Z
9tMS37VYoXsLhpLscyuwFQa0fBB0acn/cbvd9PQQGVzEq/PLRYyZY5eCzPV0s9jAlmpAQBl4rpls
9lPm2pThBF2/zzcnn+CP66te0YaFzJ6ipm8c83D0ORDnfpPMrEdkm1M8Qo+kLv89SmMdnmRepjQP
1gKX6YtgIRmWK2RAtzMeU+qvjzuQDeVP4o3nQaSKOcrFgknV32IYHl+2AfYqxzKd/xCna6tX5h7I
fvLeju0dB2d0k+izw8ATSAgCI+YeAVmS3okCezX/diWOZWCBHfP86rrRuUyhwrtxfvgsA/Hq2/d5
alBehybfkiFTPPaLSUj2z4HD9Hnr1Volq6Sbt9h6IoNUn4LjG79D56CyFBOs7o1MDr6S9JN7rktN
rmX/nazZ3+ymRkK95ruCR6Ln/3If/rfKM+0adg9Q5xqPoS+CaImV/Vbdlx68iJpZl2YZzDeJKqDA
xiVdD/lJYbC8/sw7YKKiBfW0URKAj45fl/QrpFReBw3gi2gH9c+cYYvUEE4iu+w5H8hyD8C019di
59zXZd4rG3vB8wliUQDUF5Lv+v2/nxYtavFZQzdxWLUr1wzBCRCBhrME8iRZa+NcwZVLbpAMTHGM
PQwMF0yV7UpfUEI7mYHKG7Uzx5TtAnSVfiWcqvaooSYH7ECejoRA2jRkHRDpmYepb63izvKS+M0/
E2O1SkaoWxEN+z8HymTgF5gFQFGErQRVLJ6ZfT1Ns5QDwIlDnaOfx2ah95pLqQyAyVzLczTrxFLi
baZ3Aau8bjil+21hwTq14G0XQg0fYPbMO2o4Ofvi5iBvawDG9DrdVXirgALdziht4uk7GZD2MWCb
ViiAKlKjnFNH+FqLtJS0QazqINsKFzSRV8vADB5Met7En+uiz7wQklehIVHc47/IXmwthznY31oV
kmRsVmne1N4cVpvbyjZYvZrrLiRq5dJrpQFJNwNZWU0/ZMHpZ71jxUJryJT9wTnxZOTHrx82JFS6
YsEzRZZK6/UMaxaOdttIqyQFQUW1hOxrsrr9eUpEhMk9vUo4ABN6/pD0+FoeuY4b+cq8pjAN7bq6
a6ZgDa2tnqP+uLbESd2yaqB7qz+pxHJRgZGYf0tsvsmonkZvLCYvYq41yH4gaRZ9B4K640CmpPRe
UAUOL4gKzTUuhqGtmXOlsuK600kDnE7a8a6GZVxj/Y0C5MjYUEmxieN1DG9IFNUHgDjAlTLNoa/4
vUIsurYksEmZqIKvkY8oeaoqVy71U3BxM3KgFtPZ6du7KQLBB/lAUKV90C5FqAKnLmEXTbSf179q
7iltu4AiHMKK8S6GT8hKikXAYh9qu1mZgMcjMPzV3Y56NVq1XbgdgLztRyP1vpQjM27LE36JvNt+
eUUbUtkoeyIvmeV+2uYZc1ZB68y4B6nnEDuWlqhw9QU3PpdPQZ0ucEQA155vRbUXQ0/BHvJeVmJc
+mlQ0W6BMPr5oJAnEXwyPj4/aVjns2V2mZhxDI73QlnyyXFny2ZV2lr+BLVh1egTTfeMUtsMm1KR
e3ccaNdtds/1iUhVX0eEoQ3ynenQ24ZvAFkOi1fHhA+feNOxe2lGhke1pkP46T5XlARDBQ2SYOdu
j+5ENyjxuaMb6hpC7WyMMm9L4MvaOItQ37H+R77GXVhFv85iTXx+hZzzMnxKCDKeX1c5K0HyJh+R
DJkUhurluhPTGI7gc9/CIJVikCo8ZeSDQqyydAhhjplCjZKlhjn7Seq7/kDVm1c8OFwvBtG+SvMj
hBJdFTOyrF8q5PjmKFtixMLrwqWwYdjL1WXjV2lp/UYWdUjqChrje55JE8lBZbGiqIEtl+NvueIr
6RaPchm+oXtfdV0W+embv/9OjP8LaAp4A8IF1BjCru7PHEf4XPvW04H9FaoKs6sb6lljbBB5H8Ie
1GJNe5jJ46L2XMxWDsa+ctU4DEDf5py+s42IbOpfokx8u+i20SL5NlmBz8M2ig6XOl0gC2Wzu6Qp
muZ/SkrWeggjIp/FTT+eL3zQqRfpuWXSGfVUKMB6rNk7FSLR5pomSXgnVe8wy2b5M6gVUPPrVv+r
EyczRq3DCULF337X2zkEaTJ/ZKodp6MpFzMcrVY/RwVAH/UO4G6NeLliIltOE/DtWuMcm7d8c2iL
UFWO9ypWFIqkvcnGQLiLNEe+sgm2UPGlrT0juNYDZLLbvdWerObL5yjWcOTZi9n2JFqeQP/keDEG
DkGrjR0squM2L18gGhNIk6qrStxdV+pRVveQ3S9eUYcjHQkaRAyTWlSriLC8XjoPW/sxGxeCRPf2
ncCx9wpux83x4zrXxGlMY2k6aCiN73puKNSOFY/aXwKGVd4NAkyGox64pSmc2pevcNM6hwr6HpJi
TeD2efnogCISOXdT7Gr1Ako+DZDk+dJhUKZ5Fa2XXYXD8vAEX8UmdRBa2bmgxbko60FeDOZg+k1g
g8hpxG9/4pHED/8ELVqXT2hJRWXDXSF2/Kq/sJ+l0AMQJAJV6rJi91+BZLUAEe1LmqR5gLu0JIw9
FBO0FSzn0IEOzGar6aPEfb2CPW4RL2fOg/qHy9c8f8tstxLmXtmmQ2DqHzYu4uyirECVRyHlqqJt
wMuOAL2lwO388KHBxWoIy1TwCp/21qKP9cWTXP/y7EI8vMTvJMZD2sifjV//85EOucqGYwvL5c49
hRoTIA5Ee8+6yw+TiCckGLZNWbodCJSx84E+3hsUSv7fPcafn/a2z1FfTt2FBTvl01xvTp+NYw4M
/Lvq2Vds/Hlt59knFon0E9pNQqtHL1cmG4lQPr2ECqXNB5LqSnNBhhWQvOSViR/54mOdCG0yoeK3
gk9OVDwzCsBfkkpybjtmapKN4IwGJ55qqyO/fjwV+R71/RtSFV9/x7WFA5m8wQb+ypq7RFjGI6UW
r+iDwd1dOdBl6+Pxc2DBihAB+lA600WjlN3LZebYPeOzOakuDo1twSr4yHSOtaZ7f1Gkt3D+zi6f
tyaoetY/b34ZgXXrQSVaeLtD1ZToowXptPYSKiALMFII0MiE3C31C/hmHat72cybqXxdl9U59Jut
D9Os8UFx57jVzXJzY/84zsH1Da1y6CV9m2dZFGE5+dpEGunx1WBetHl1jQgfWfTij+3cvb6r1xim
WQALwx1C/304NLcvPx4ZGHnTL5ofUF9Dj3yDcP5mtJnKG8VKGK73UbMSScP07HNEP5X91T9iCck1
rpjdNzx4IuJ+w9lYbs20ZAXswHPCWr7cO/Fi8Phg4D2aA7Bir9OU9hi2PLFJcadIpMC8Bk7vPPUm
ZwnOoe7B7B3Qb7JMFPfPHcjkwPaNhOGwzPgJ3jqULZ0Wc1cCi7MDQJfyMsjDTVl21SMn0HlLPqB+
ODO5RZiWyA5MH8qO3eZ7RT3094uSHSc+1qaSxQ9ZcuKYcZ/gjhHPlxMIC8f3sdOJAk4c6zZjvY7V
cIGUZBb9AgqPzZ5JVy7lSrU0Y2sjTNJG4DfJn+uIpw8ZnA4UN9h0h5T0As9c2ZZAtGBZTwvkBuQE
/1bWWQCDEFkXipzjzoIu92imccM3sXto2mzt7LRg3X5zgj8kpchG0J7uqSbVcxfI4wXvkxXld//M
gv/0Mh4Zzm2Js9xQyQb7ZfRWC2LBWiqcy3o9cCx7z/JLAnZJ72G9HDTZqBXmL8dvQKf74S4IVMWe
/2N656WP1fl7WieY2i/3vRyCZIk5IM/TE0CNiZACaf/8cDRHJDnXnOj9qifTkXBOsijOB3uu8NyB
A5v1Ky1eSlJEgiG7xBVYkP44Cei1QIoINZCsFD+jERqEfcqvCDT5VkdGnp7v8eVqkXhtk20W3Xe6
NtfuwuMNKDVCYt1OlBy/jN2D0UlXMw56zTZnK9fqlF6ORklPBaRdq6wwd1Il0P4mMaJMIcvo3wCR
LFHUnVHRsJuqBDR0k1XZh5PN9bXA2b+M0EJL903MwzKlJ5mFRY7X83vczS1Bmrv6lm1T5YAt3VmO
D+E241UVUTphJlQhX0Jq8+Dlf0YNJV3ZaC/6V2ptCczPsVY53qCNsUCzYR8UoCUh0eFdCh4FQ+p4
dVhZhydywF7hJN0KYVfIT7LfYCVH7wtSQ+xXKoGvDakQURYitwjCAKPANkrDDMO2B+m/Mkd3iv3S
6Hs2zwLvrBwGgF7+rXZhz5+zuBFztwzotlDolybXH6dJHWNZLGq8SVGSXoG4x6xIRFjhbLc9E+Xy
ejDfkLEssvE+++uxMM2cnJddc0Bc9mtpSgEBukYtZSAHDX+g0rhpE42VmGl8gxHJVu46PbIeBR9n
U7YkcryLVKo6nWSGiTRaaKV8lRFswbjSke1/tVPoMLezjCTD3FlTfVIS2RB/VGZLxuJX9YIGp5OC
I6tOhzugsh5j2Qt12d/UV6a/gjPtOvJUqwr+71oo/i/T9SgjM1UF7yM3eCl82s/aZYd7AkFq/DAE
VV+Ihs9eyCaTqxxWxDC1nUQ015/4eyUswgIDfrh2gEYw1Hls70M7CzFN4jKtklaAowGDwlCZfbwG
Jf20I0NvBf4z/N5iC7606lRD5vm3tOLy+F7ZAYJIjkHnHHNvtgczX2G7ltI+C2EfB+jjBqUJvvMS
Zo4VYzRUps4aAqIYYUvHZVq1L2Ot04bwtK+GJ0qfJG9ASc1K+nKszxfdd41Mt2qhb1LgZqf/NTZz
opI09SISJ6XgZ+WY8Yd4q/NarmYba0y5A106RUazSZ/SnZiBI+2A32iONV6gy+WX99ku+4ZKI4mQ
F5W3L2D3iO6GhRGrbugHkylmCGJrIFzWXWU20E4aATj0FVnYzrGXdu4pyEsYIBb1fqXcYTr3sTCb
SaG3pbB4UXM+ANCAQroBeVF+ctTSGak7ubGJkFc/jb+vOWz5CM80TZTvxlLy6WX3YjGJhQ3cWX+K
CxvVdcJ5uHZj+FDZyJtYXDWu3jc4lTv5amSZtjoOJVjMQUsdp2ooOF0jhnhlLWhXKHOCLW6wy4NW
i8AVSl7YO2HWkEm26MFc64E8S6eIp6GUyCDnt8jQCnXEeS10GWU+mqqn1qPGnrJsZbnwvyhSXTRE
2VQKff8VHkXoYo0YtpTiLjlxzKQGCRHws71+zMtwwrzYdwyKkzQ29V02Lbal6T5L+tEIIZdGrTnD
BfPORd6qRGYKa8PEA+RU5QcNHSQRIMgkbubx43IoB/G487eBF3gVf0HYDWOsPnEdX+KF3aqirnl/
gck3wpKvs94Owskacy4/XDiOgE82sj5D2HIgzE7jG4QDNw7hsRm7WqFmeSMQ7C72tmFN0GZ+ycmt
f+Luf9zKu+2kNv/3KnFuKuiPku+D0QNDpDH0llwwOT8dvwjnoFUHZYixcyz0D/YMzDyn3+D8EE5m
xxk0+7EVx/4PCDOLDcn0XU126ueScklr3gU/q+zNOUYib52SsfAjwCAzNhlmeiUU/I7SsNz4SiNi
tRjQYmJeEN088ZhAfaGqWYxOowP74Ujd0rTFoRcJwkRo+y9+Rody25+Gx0K047FMhwRnWNsh1NqU
CAXqnoVvqfZGrn1k3kW89Lmr8Jw4ysGx1+mjBysZ+jzhBoUSHffM49vZuOFA+X18XxfpxqRQCvXT
98q4rw0fRAsaa+SApFE8ElcPc1HskmmKPoBM/4FbMn0MSIlQ/9ipdz8K84wZp/8dFLj5NhGPFXph
Tpv5ubLZyZ3TZVLpwctX9pF6hPiH7fWIvHbG/C6XHflyudWjIMeWsg0gdxohYR7r5jBiZ6oqWOlO
8Rms+FOoMHIclB7TSBBQd2wDnGXq9F0VMcO2X7Gk9Tb4XbUM38K/QuaF6/R81N+1aDlN8dDbmqgU
LY9ko8Bo7IGP7/Rj915BsjaQvQm2lbDE2c96mAEZv2a5F61OTwZXwzvT40dToVUZzWYSDYw4tPJw
6G65UQVOoPQVIcipPAfSRtzKurRV/0Bk87gUDgxzlwy9wxTSGMwGOR9KRexSacfqNtdRN+8aIX3z
+5fSTHtmUXm0dd8YKUhTxOTtzpP+YSo6uhkajnjSwmNJAy9rm8F7nSYVKwEsndOU7NUDhFNwg3X+
vfTRsphT0A8oVDD3OJrtxEL3o+uKiJ0jJIPQk/winiN/indSwnqeawnsdc/v02dwwKH+Mjbf6/L2
ZDprUqynUiDcncYVjqKXmRaxtHtneQUz+AY95Xr8uaVQsPEMuMKWt5jgdMXSG3mhtPMnpL5el2HC
eJJ48MO5/kEILRniD4yVLDdnbyquul0eMReowVgNspYqbAJMOkNBvS2BRBZHBcRqSLxdo07JorVH
03IU4PIvPuU1QW9ttSNB64ww4BVvpCEMsaYQS04uZM+abwEBYtid/tDAEEEHDR9oTgV/pAwAV3qb
tA4CUtE3+UXoOCeUWFpead8NQ77DK16fT64rJiUe0gwahWo+nyFDIKxXuUbxQOI60U8BcVVIGQC3
s/X1KgUoRQlnQAXip/MJCgSjkvLHOvF6cEquTSlhII4m2JTTdrixVdQQoMo0hc+T7OKMEsrG1wK2
VsKjDy8vOeixjLqLynjKkgNrTzSdqs81P+RmPplebQBAmX3by90XhcKUTH6nvMlsuTxoMMwvUFSP
IMnPJV5aK8mssEoEly80Fa0rMtMbXNAVGvrfvl16OwAS5J5jT+skU678wXVr7XfLSXSO5e5H3mPb
CoCQL99862AycZOu5HluusFH3wu3n5iHstkwbF4+0s+19BPTnsod7JlPCtuPxtEnrFs4p2Qg/WgX
QSttPkztnPrDwV10MwwoPA993QuUPzjenvTtYdbfTB8CCd+mIikh/UtBP2bHAU3NqtYZojGzSuBA
GmIYUkH7RcfbTQBI2S17I1j7D7ifEjJYBWD/vN9d6N2o/spmvj20h+2+v7mQX2+4VXBXGiUMkHqX
lEBDboskn8WjCBShnHz8EAA5MCnRYamqRuHLh9k0q4cpcEWGcS4MSsSekkc2jm3DZ/Y/42MAjPXz
QllB2rmNKkScxs308bjzg0Vn6bqX0fqKZ7E2s9FFf1fo+2dIrpp/MofZpseZIVRFBLyxhri+YJAN
A+Dg1ELljmyEEiZO9di/IDyHSCag3+G95DNdWJCaVECTJ3zS2k6+JKmUDfSHNH6TE/Tp+Nud2Dt5
RyGlk9KHW1BjpfMmbH7ODM8MvPTmkifGoRqQS0WtezVF6Ag001+QlTD8R5XQJT/+YHYpPFBPXIps
nwXsgL9k05PRCTJKuhrY74DV/k3K/48uGZLVxGqtRwX5auH0kFtYfp40Y9Irb/F67UoAsYmKGDLn
i9P4huaHgbCq2WoS4JXQa7sfAWmryRfudJuuLFg9a/in5Nh0sdw18ehzN+3ny2Ukk1dHbqlAVvYL
xGp8NxnNZhlNH2oCkmpigSeFZgsjmFBZJQa4HQCQbNM7AP9Hj1PAM7MOkOiLfVoAMQxKPSX+WPIX
J4jJ1E79AKWNm84QHlu9Egn/jKZwYT8LbeFuhXtpEMF/gpZGXIWdvxyIFnlqDVMHWvYmFh40x7o7
GE/E4Mm7tvwc84jyOIqLcCmGLTSHwz5X0slGHYhjGupjjDE2aVRaHUeKQMdikGd1ZRnjl86KTiIE
CxPV/IJ5MT5SgQcMOsYMQ5f/I0O3qEjFjHgx+oGRQ+e9s90RBNbix8P3zY7gGeCdEfNfHOg5L4fT
A27vMKJs573uqnIGw1MaSULejvnj4PTRi6JGbQ46RSWl0w5xoOgCEa6hdu11B0GdpkDtA+yqVINX
noSFmzKE3uD/TRhz0rOrOXyYbvCLI/TS1LAYa7Fcymt+e3r6OsQImNvAQamYqc9JPgv1xnaWEWPp
8emac7toou+j+0FZc9yZpVWSUpDm9rDkAzYB9rE6LzIlz7XveV1gQGH+0D9JUM9d9sadjl3t7gGM
kAQsV3gB2llliIx0PIrgVK0gfkSJL5gbOM+5eUUeQwNOkia0N5jf2etXpnml1ihAbHul4rJgfO/H
laM1P6QHo5jr0CPCF1VFKycl8DlXsHt4R8BmoRVx7oLs4pMukQEGWyVafcHwxnprpWfVRH7Y7Iw+
M8yoyIyKkhlLFh76O0WhOf7lvBck6N4hbP01bYHCOBkRx41t3gTjjuKjyAGNZek5r3ILjKg1sczL
j3iCRoiWS9JuRGLyaUr27C5Y8tC51Q/jDdQ+XTiAOCGA/tFxO1bMU7mxlI2aBqDS6iAeUzoCHyXC
nn8BeOByK3cI3b1XfKDREPwvI6+SMSfrvHEZJ2AkmgzQ6wveDmX4JfultEFa1eM88fB4EaJs5A25
jCeQaCuv1huJ5PbrzmaX7T9TJMdEWTLOGqreeH3N3FIyPaNOyFdsIRMI18tDOCN/Uc/AIKWsunWC
PU8DTTvOQ3nuYZuNygfcitlwNmaISNXcMwred2r8U+5r+NyNlwgCuryOIiTrn4/q0H3DX4cUGJLL
0+C3Ovx8k58N+LaDo9pIxaBDrHkQ7Q2RKtGPsczxvNoRv3I0LJgKWPCGPRFVV/pz2KthI1YXkp5R
EQv7v9nvfTYe00vxsLQGrW/PrJePd7JCavPUoqOrasQ2LePmnB6hMiNiHYC2QUMZVwEW/EomlkYk
+Jj66LP1UmGpbYSc4L+ar5b9NVu+VPf8xDtdq6OTbZbz8mxVcxElyghAi/rbRzXvep7k7rnPpWpg
0hYIHDNWIUWVIhuedBnc9iYcVKVWkZdaOIe3U80etA4v8DnsVSflrQvfNnGKM5H9UW5VIVCgZyGx
lSRpJKB4pR+fQgChhoVtTLZwnJuVRTB5v8TDW+brYRAbFdfFKzTCBMSxty60Z6h9EoH2XaK9Ieq6
GnlgiWqVaBq0KBg0BzuUdUxy1qBgEadNDXfyIl6GdU57OwhcsAEgtEqMEldSRGmRapYNX7fwcazi
DvUUszA22tGxM0/BKD/iJDLg4EibIsRBX7G1/fYN9Ox98fpE/Dsg3AbHZyWJ1YSMDwscFVL2kCfq
9yh8A4OR0DNcczyMGVvJetgEJMSQAYnN2gmxckr2xneOUMuB/Qr1/yjocGiRoFdLR/qZWOsNVCOF
teKbsLOegnYPoKlCqlOYZvE5lTV+ZpemRyJPRiXF487HD9IWEaauPIcbteVSeoLgBIPKir3iPbau
NQxXNYAW4Dx6g9h164Vni1SwNWkoo9kj5CUxq8OZTIcms68wnYTMSJkjBjgKSgCVP7e5eeZlo+dW
BqFHbdl0yti1/fT5po/fCUQqShWOcVZYFcPi1iq4ghc7NNw7Ofxub0P+tIxG3i9OVnH311OuQ8kp
E0PZB3Fi/W1QydUeR17+33CiyhrI7cbr50oJDpRgz+T5WHPk+rPs7YuCaTdfPbprsyRlpoXcikSO
4BObsuMqa1aW5D9BfA0H95WuTy8rY8ytudCdNjuur+fhwYj7vqx1Z/fU8g7n5N/IuKQxbkbKXPVF
icVgGeirqYhubIDav70GxXvBswFAJDg+uvdK4KMzo274gcaymqovuSE1mTRRz4CSuPq1YqrAAQgE
51JHiY0dsLkHZK8ViDFDBiqtOQyUo0xXFSM/SQ820/iSyKEt3clUrz6ILilJlazjPIX82QqjuTdJ
ChL1Z5CsiMd02ixcJ3tTlVGVUhO8+JkSti07Y+gNPc2naCei8+2rJVv/MFcJAGAhG/At5c3jHdGe
jv1yd3qa5vU42eBNmMuyBVFSiqzFfpX3hQ1jHDUrx5IrFJq53MrPUYzW3d45KYly8OtZdxB9UqXH
aNF0+fYqW4Cs3WVCNFYG2siAjR5TMo+74gyU8kG3kBQ3Qq0nLsyOVvr3JmELqr1YhTDV3RKbu2K/
GuBOknBdtn8QBMNXbMwpEbwac6Y1DwrLxzzIcqBDI4Z07+G3sL3aiysZPURYqYNdaEMr1A+JDEuz
BV96i2VK7N3CSNUHWe+dcuNxNykUoLNA0v/9vxbyqnGZF5B5fY3HqWIneIdY8VAYOurdAs0Lf9DE
HJDiJwAnZjC42+aSH53kocE9LE3soTk3/eoggJ/ZckD35pQPQT1STMuTvYAEkc7cHOZgoSvi8HY6
lS67paD7uJWPqlVjnrxi+6IFpAIDGWMmySggKwQMwXHCIoccthvkxIcrVKZ8dyR2nyGLu5RKRW31
ggfHnKDkFIqqExP7JC0UnQOMILYHssRfhYoyryKEvRVKpq9lDj33rYB2h56fxVNk4hw6gB9sBkDf
YiP8gvy5h46LENsCz/SanfRszRRjTKyAX5DfW+cnJW/ii0hBJf0VSCf8r9U5PZ5z6ScZrcdAUoPt
Wn0vhogF495ub4GM8g3W7K0MXcitNtBcvlWWLqIvG++s5sNdu6UQzaUqhkMp7AqDR2UTidosaEPp
kC5t3vlRjSttcr2AUjzm32HoK0BBsg7Hv6jBx4X7+hmOTsEnr9Ii3csW9wkWgq3aoN5NZyr/U+8l
geL5ZArHJ2ZE1vnenam6GfaW7W1YicRfPwwL1YMBsFNcm3MGEYe5EKqybvzI8MJwSux1vS1h5E0z
Q2z2MTGuKbCiSDL48C312Rx/gSiJ9Yo5qSA0mXzWiRYVEAbUoFUqxqqHJp2vAk+kMiW19sHpg+JB
MbI+DFFWKywk7Atqt8XhRkxt9z0YgJ4awisEYvEO+81WXkLmikj+Rm8L38WxE4B4wEvSNMPaMeLU
PnZQh89VDhdtuA0Bj2WtMZ/LBnYuKBrKk2t0zZkj12l6ssF3/Wun0tREsZ3V7QjgsOjfYKRRnLIE
Rys7oZiLLN1hfqvpBzKVM/8rQpGbI3DphkXqQK4nx8410Dvb2ZiVCkyIxhdJPs44/h1qqzciGONm
yKt8Or8/EpJQbeldYTZOzJoG0ASseBzJXqaKHtVQYXa4Ga3gtkKcy+uUlEMOcK7qIIzmTy1l4Rel
5KPbLDs91fzHzENHK6vSj59zfSJdc8+h7Cm1W9zuGgS2bbtI6tvuhmX6Spc6SXDAIQgZILsk4DmV
HiVw855iig6cNi1IZoopWPTMmqfzhnGrrv+1snwK+6o9/iLVUSLukoZP6uLceHjQSDt0KxGR2KhD
NzQEx9hib/34eb3CZkH8GTGj4ItEbqfwMYfJPWuIG7bc4WmqIWsYmREJ3f3k4Fz/z2wAlrqTLmMg
XV9GWjbqDQKgQ42bdQrFx1Q6a7kEcFMzAPHya02NfFXU0xdi8uhjtDuUBqmKoePKFQhuciPPMYPZ
3RNcB/ez6i1F39P4psmFXur8By3zQCy8kBIT5b2Pphv65yXmEPYdpVTnv+TzrMWPieMZ6LH5sxOU
gTUpgsokPnLhxaVqKENpmnri8/eANrNAD774I5vzRR79yn7PbmgN3+zJEom2T+rpkr5dZFeu5TdA
3z/CiEMxp1hjq/FytJ8W4RYn87QzpeWuRlKuIh1NYff79Okt4NZ1yUyqqHmECMwOs+9Xsd485M5k
rgIgfQTiHXsF83ng2ObpMZcY47iujx1Q7wKLscdniSgbsVjHY75E8vXp8NeqtyInUiQZjySpUHpn
r7xxcwIbvYwjeCyHcv+ZqvWbH8JTP//dWwasMKADJ+okgCyfYM5iKRcasx+zpeQgjxqDABTQMCuD
Vb9KvsBRl1rI1JaEpcKaybaCWwQHxWCAJbOyT2pDPlBZfik2bBbpNQdigEdzGEuKYsPLHc+OXKY0
sQyTS6b2txS4ozxuZXXxJ2AaJRKOS/SG2Gvnu28GlWlnIV/EwDT76Mo5oMayXlma36XvcGiddAWZ
wh6r8Tbxu0mSAnKs3/qXG99Pa+2O0yzq4w6p3Yu4eWfxhlXfJfDshQ12hekts1epq4ifpuI7LkPD
zH4eMfC710nNarfP6hpvA8CpRZMuKzqS2tSMuxhVzNqL9of0zGST3JFc+4q3gR10sPbGy4t8s/hr
NeDx3/kMVwxSvLxhnUxDzwgAnvbNZxQPOwedI1JSwQ0SQrpLqM8A9WVf14yPcwYMuwaqohV4a/cu
cLbk2WuWyXySn6+p+FW7wPJTEJaXd39or6mD9t8C4tBBRgPkJop3l2n74H8VI+4DM2yTSX90wnhP
8NV/cp4bE2aaFABr+LYTDAlaTnFwyUq3G3jfEHtVmIqmCiRRArvrdb0tG2ejItIzZdTgRX3cwEuw
1hOgftL84Us1Q9qyQ5I75yvMKFRWrWsVIibHjES3sd13RkapxBf0Jh1R+QCG61XoglUs5VMS+7ay
c+0DT+cJmT/oJkQ84PK/QMlzEjhAnjFeAmL13RX59t49CMwiIvFdPw6YqL1KKehRPypMwdJmexYz
sDfVvBsocdjnV/U9xyujv1bp0PCSZcg725/lDnCmDed621taOpk2p7NRojIueWDE2G3gUqyv4lEM
u6m7ziFBl11CI/EXZfmcVegt7Z4as54/IiA2lorLLmacHwaGdi3yzzWevN1idswoiBQGKYRwH1cL
frIJuQiECZ8Chx7UykJpE9IBP1knWJQVZlMW8m4y878WcJO4OxbanTXv4FAxxOVPK0jPhzducEcB
RhN7u8k2JXSKGTi7Tp/aXObxoZjBXJO+bGrExBRaN4e0DrJ9bpNrn+YypkIXezLttpTGuCMM+eA9
qv8EONXADNqu/RIGgpn/xbpaU3Uwy5/J9RaTmfsMkiTAxmWhv8z+m5X+4CH0OyuQp4QJ72GDnMfA
p8hZQlIJr3QKUp+8nqQ3ZhPm5oXsUnx9MNEuu5TAg54+flrP615msTJ8YSHyKmni/aPzgC3mm9Bw
khug+etd0HJYKKtx/to6zPvQUsrmI8+SOS3uS6NFIipHx9+mxxGXr8UcubqvuxlSoEXCBtxgTFtg
1PctfSQzbOmA+4WSBBRqDdiEKneEIi3oE0ZLN+OtZK+RC3RTKFuBzm253xNRrIJ/NwY0abGtYN6J
UDsdHRIQknr+3rWo2hW23/XeS9fyrehg5g8xQOOL724AFG70Cx3qULaI4iKbp2gAUeWd9ctLnt8I
3nIEV7ratx3wNwcVdzfxVyk0BkCKjcSRTkl/cG8Djmi6codABWBlvE+lAdV0m98DGDDwSKkG3u8P
kDhvA7yGrWCOcemcxOIfxlGDBb32MNSmVyBavIdmO7Ptpp8/Wv2jLR5dLxoDzjF2RxjE0Sxnkr8R
X500O45L8/l4B6ccUhbwartnWyQD86PQ5Xs5mwV6pQ2ShIKFuMlG/9hPsnK/jxxPyqRERvoLl1sA
03WlGLG465YqNzMDzecdq+rZBYZ+KGNvhOga1LJj1kzNIUOmItPhfSjusTNwERO/VXY6iQ32csVv
kIKaxvn2dZS3r0f5JqeNk2XW6QS/q1dl/NTbt30kDeXwV9MyfAI9/Vokick904sLmxawy6qV0bxJ
mJYj7L6hFZ79yvL/JRt4bYpBLtHXZxCst4CKw18kgz4c4Q8RrPVvBh8QuLOlGElW/IbwZkZgV2H+
o84y3ygiAqVf64Af3HGMVaAfylKBl/UkTs7gSGJgO8mJXgQOzYFCM5ufw5ML5HJqqSa7ra1gZvUS
N40laKL2o+SQXNQfQKHyufs6clbPN5L+FOUHuh6zpTWODjOLYSJiaMhAFC50Ey6IhgrFBcAJnsEN
YccO8Zc+NfG1y9DFBxN5SJ2wtLQitQ7Y36+uZ5vHI7xmqFNtAsqNXmg4+t+DTJ4Dw+H4CKXYxogB
18yBNv0DIIhejTOsZ5v3UkiTHKxK7HtZ7kd4DSUMHyyWYE80Owd0g+TwCdH4BWxdFr1K+Uh86MWt
H/opawOFA1Gj+1OtqVJF1jDliwWXz3gSA23c4jUaOFIpsJ+QgXp3Ca29MPR8SSJzwLJZV/JoMbTf
1ok2sO1rkizquRMn1D03h719icd1VVusNJagLAtXcrVA+mKekcbfenTtSUQfRFPJ1esvjccsbq0C
e9vArv/fBH70TJ2oDi9VnvCyQ05imdckBXlRmtJ8qPqj8Wf7rI+E9P1nNiX8fV8dUN+ueJzQ8J3M
Hl7LSFG2alWHN3ksBemyDpVphlDjCKIEnKEn+G2CgO9HKm6FugSMOz3EhW5lOlQx7A45VZwNUB96
t7a/qk1H5KAUbfu3VUSO4zWvU+j39sT4beLc6ddf/63uQZK4dUaJsZA0SSfcnMCc9az29UsrtaWO
W19c+ilvlre+wThcGlLUaHXI3mA2QEUragAhQhpBcVz3ediSsTxjFapGdA5Bxy+zg1hPGXbfmCro
ZYRVLiZOlGdLBttmPKgdWat2uVnZ7GJhUId2qIydr5Pqk3zUXT/F09C0cmKRWMDShtGP+y29iU/z
jWGiCBiDiNQPhu7cJ/bxgcZtlHgMOAi8otm2BqG32XwuD1Ysu6poWek2yb7zIssCcPtw52iRJ1iy
1teyIXOwKPhpy2Sj6hOJNCL2yyT5/iRo9COub6xJQHvTt/C0nWIQuMAZU6SKCrlk5/vUlXI1qXs9
72iGE0Repj8ASNCGj98W8VXtA142ZDZpOgPbZDVtUrIOtbNY4hqzTojGVS2TYKhBPhNfUCyDdApq
q1IYmMoiX2jiWvGBBLE5sqdRLGK4Jj1QiZZpwF0igvuTSknZhrDZC56Foafwbsg/GjjBs6020wl1
VycNpAgtD7FXM9jASaV1GRyyYMG6Y5+DgoARvx8Jxgl+EmLFzSgXeFmyk0mnbBDY6Tr9x2zJAF51
yukvRFnTdddEfO7Rh66QF+3q1MrUaK6uinwg40N1R7xal/FerFFWwlVALjT5bhx4XyoSoz+mzBoX
2ixCrEjDisU1jpabq4sODASQv0JLM8ZekrWDZkgIKZHd3AeVzkw0FfDzMrWoubPs7rlgJuC2Tkl/
LJ51BajfGhJErd63hqNqI824m2MBOyckYl+MMzRU9oaRavPtmBnkabB2jOxw/e1qVCispZRvupi6
mAtnb3Sv/reR+y2wAEQzJJesn8n9uIb0SgC1UR70s/HZrEd7ByqFTpt7//bd6C5hxlhSeP4UpxyA
tKWl3sK0eqOeUSQgJNvlOX6hEuDPpkxTWbe2mMYtNHrq32D3c2oc7myPi5SzS3MxkogXku51fRgQ
LCXJTZGkvwxyhpbN9Y86BkqsK97hNQT6iFkS87/gnaaTgtNKpdr3wi8g/5ml6I/54jpNbUbgvQJV
/BnUSrY2ezM4Nk7IKXnqsjh6VaDly64nRy8cz7Kl+RYhbwHSInNlbbYxnTwg4JRmdSlX7OHmw3xc
r7AC12g0a7FoGzIkrskM9zEWgmCuDqp+/l7pp1XM680Ymg2Yrm0F10Hy5pqTCpmlaE0IjoRe773x
X91Jcfa8Qdy2C7by83dwufrCzQfLqkXa4QVmi/ZOo/DX6wYj5qdUBIvs59J7kS/vVtXGmabz36uJ
e581hiWRLx/Hy9Cesgbw1RqeAr5HyS3B8gBVtUZbKO0Cu7SaHeiltPk3E8IC6ad8SgxtJNRzwwjB
FtssyA0s2UJfBKqf8wiQFLlhAMCcH3HMpXIskqVOKW2JTzlpjgJOIbedYlVlYDw3ytjthtJlZ00p
QkXhxpbQbZcQf7j9AzGgkaVBK5+ZEX/A4i0SXI4ilwSGHlzYKYj0IDtjSlE819hG+qCS4JB1O7pX
PmL/7c+YG00k4k3QEhD4OFa9XOOYknvvnBGChOmclYk7ok2IebcEH2I4o/JLwhsldfKI4lnFi6eK
CU7PZESuyjur3WbEF29mXQukhwLb6ka7xIH66F2S4bNDOC9+U86IwTbwJnWma3Xwm1UUs01tYPyN
5LFZyCSWViM/QZdxOTs2JpVjfgHSgl6RBo7FkLW+lE8VBAv2Hi9RC1ROrGcDP/TmrKQ7RLVnOMh+
0LNST2SYkN73cyA7E/xRbCrFgLXeDa1nSaE/2W58XNOJHGq0kyWNMSMRgOt8yeQTK1twWfBWUbAi
+UEqcNpOSTAvEMndjQqBLgRgdI2zqJe1Q+FcCtpk3QWvQczpvEM26dl0ELns53c0Q7lupOyBW7UC
koy6gh0IbEiMKYqociitC+AcZBbVbt7DaKZcsOTMZ3I0GnupZ7tVytMGBahM9p8yfPRdq7hKAuU+
SGUe89ZasglQ+6jR2O+RuiqXj59ayPzwUmy+YpDiZY8wI1zkdu17kSSlMHTFZfdvfUvCINcYoeli
1pvzeNSeio8a7giD9VFvAY+ajO9Hwykg8wZ0Rk0DxqaRZVoWNfkrSatz4wlrxc+dIPYqBsLHRUcW
I7GuNnGj5fPuC2PBty3OLGSQeFShmnwptk9yehipH6TZgNeDIbIK1A9hRAC9RdPHWUCFdAJg4BEJ
vx2LuxvIIiEeUVYOST1t3nAh48Rh9i5C5HSyFq6/UjHlH8JKEXI3ACJuyaith0uAzUVdmDMrhpwK
xAdAz7suWJzZeIWU44lO57HNF3UN9sCREmf2kltU0xzcyGAUFhG+WX1LNPOMntGfR+6vv5f0cnbv
LBYvpg64dNEFsTCG+Za1JTNfmHtNiLCY6YZyOs3Ig8aRb6kHyKmNsmdZ6a0kHx2nks7Nitr9PRD7
6MChWu0nGJMQo6UJjflofJKN5ptAkmAjuz2jpDqvhvPmXE6OXmGDecZQA41HzAsSz8aAHQNbsxyM
qyzDV/8x33lqiLDBxkG6g5ZwiV2frKD50AmMa3NyCBtzolbc1VP1NLdj5c781PNXn7VUlnJ7zTeK
RVHTeNen32xikf+QZPZm8rmVKmZSvUeZ4Vc+DUwVIi83biyNFgWlJ3+GY40LFqvB6/eqXpwJrd6p
Asz2llf5N8DotEZHdTPPd+mOOYeiRsErXlC4VE3JcOKtqaM7r3b7rJgFURemI9Arl3+rGYmFGuKq
jOsBGQFZhpnmyob/T3E0KqCiGJuTec4oUbm2R48Zi6dx7yiNS/qoDoT3AL6zRQ+FLOQ2lXp2z6Hn
sNn61nkgKDtFmpp3bsGWtysyrzFX3i04FifnFE0mnjZXhjk2mOsbo2fDZoF9xU1nCTbi/D/GQgKn
Fbp4jg9X2xG4EPUzMz43ahWxYxqh0w+s9QnNiWn3XRBlRyOl6YB5bzGXwhuE1k3VW7vpo3G0wfA7
jZ9+u84M5Ei89ztAls2BzAWxlO6IfyL5VD00g06vSltKEou3B0D+UXgig6g1OSshhW/pO+KvpJ+4
/MDIqZCSaX9oFdSTkrOtBPLhj7caWxB0weueIz1GUG4U3JVsfa8y3yTDZ3vrh6rZCfH8qCycl35y
w5B+1686CiUZmOhOuZ2R4TBNoHQrKIB7m0ZotjqLFai/1dcxoSA9+gPruUbJbfFf0vL+2dYeD+nz
/ZAPp/f9OTbSOkka9iC3UDev7drIUDD8A6VQ21uZXrJiIMT39i82LZ2QV28rfnRQ7F7LRNA5KcJT
iQAGKSqkuD19WubTrJqAfjXLjugpaXDeX6ppQjYqBO02P5E3ovlDhMjJr8TWK007/rgZdEZo57g1
PTSqPOQ+NprS+o9yKBbE8YTgtaBDkBcc8DUNkSm9F+zxMiwVAo0JQu65QCEErqq2FOvx158JShpu
vvcpQLxLej8V1niR7hH6nXF/6fl1rb6BIdNZFD9WTuIhQIYyyGQflwEVXgT4KE7rd3UGYGWiTtvj
GDkZUaP/OmNxWopBM1dW3yulVETb79RN7jzJDNmgFQJJRLwiHnjRZ125bRjVHnrgwNW3VPFaZJYs
f77sbgev0oIfkQ5299Y9D2165Jxz/8yd06s3DfuX/XbdTWUItEkn21MG+QYNULhF6LNo9QBjxGCb
Fr2268BDnzDUIsKmED0P/e8iwIBVkdXhrTqiH7w20VIMXv6Nproq0kO/rJosT7L6+eiUVTkEUfwu
ulcAM/259SDcTgGVlyp7OdmCgsK6qM2+HYa5ku8YaZ2sIo7qgL1o8VOuwm13ev5wDkkfy7VSw1EQ
nCddoEVlqB17lYWdANi6GduQcmJciPCdHpqXYTKMIPG5YGBlQxBa7zhxlqbi07M9rn+we54n7mCW
tdld1CB0RPs4dM8c6q7aUZArVySUhPBJcqi0zvtkP8vMy9c6b0+a2gvGlc0QftoUEvgzoO3qgKUE
EVMSb/nUxWIL8owe4yRe3AcqUaaiSbuYKSKxQc0tGYaqAneX3Xk2bpDBAjOuXSroCfAjmjv35N8/
3b93vUnR1XWUapkRQ0W61cRrXPTu6sXuyaHilfjuk82a4ZlMO5IVxEzqim8ovxicf9y//gPVOUoD
V6ubGuWELlrrSKsAZKNMZvW2kQX3gu1iOBmGqmPjEM657W/9NnaCyhPv5ud7OvKRmwIUHhkjIaJV
+8N0oNq5zps4DXxYY+CvegzgC14SYJ4564ag3ohH0Av+sWc/+G3ocHYpW2P8z3Z9DC+WqzGiSZyS
bOOMuVQPyRXWX+T2BZPaE+IPL//eQ/oGpG8VryOlVA1rKHJSd51vtOscT/txVyaMcm27tnXC+gu5
5Lug0Jb+0x9v6mmM4wzm8QPdtBAKkbG/48s/j5awr+wYy+4wxmbPcot+pCQVGTBqbyOBTPDoGkxp
jXyo1Yo31U9lHCEfihVfKtvLQXLUMfbpGP5gj/82rACVIJoNphLdqh8r/z/GmHFQBUiQDY1ckfKv
DdbEmOzlQSt8y/xEweSZSIX+Q35l1pk+ODL7J9QYyQ6Ybk4f8s5to57XmliI+ZP0JJx0cAxMs1/R
4yMN+fwKC63/kAyZzLgxC9vugSYQhnuYjbnfKIvQY/FL1buxgTrJojjBwbMB0fn7YPHC2ggOTtue
+iYlWOnClUm66KgFECBc0sRM3faKmf4qs8BpPVwiyGRFKtw2+zIqwNZc4eskueQhMhi/MO80jdlt
T4B6SCfkLEPSKOn0GPlRf0Sha6o9QVW2prAd5t83WyvP8+XTnq5mfviDUq2mGSqPuLAKfZV1g33B
sDAFG1+DueCFRbLHi/Jmnv+jjlrpi9fRQdfhDwfHeSpY51+9WHx2aelOlZvJV38ydEZmKOZOIema
LVGFtOqQ4VbEYHlyoUR9KQyfJRYWH8gkr5p6Wa++1dbtbkb566OPyeY2o6kxzsLzfYH00pBHIVqW
ArQxA2pYAcf1XnFtyN/+MriD9k+89DgQZMP0SEi4k/j6vUDEcAW/jNeRPy9yTEt7lKdXZ+I2EqHu
CdmKwQ6q64GDocNdght25dV+wcr66Vhtvnxo04YUQ8bSjc55THwuwDHcUQkUCcO2rqoGAlwSAUr+
B0PRubYuE0Eu+8enYIHMoAkJr9aowtiQZh1OwPFKlbyiPJPDpDHYysaX+9dtRbjslnXmZk+pdweZ
dozyjT+V7xV+TgKBWkQcec8YA6N8j+u+vlI3Co26mrwo6UQZ7IxiJ4kcYenFTJy4XplITaZLzR5K
EZz9fphWN63kXNLztKXRrzSodxYOoZ2oDJkPX/TtiZMqghbiSLfKi7WVsB+kQg583Hdt6Z+v5M2r
QxwwKGyxxT7EoCjevwbN46f9JkQ03vphG2/xIKBJrR3jF84Z1ruLDVMy73dsJZaXAu0vnaV5lg0F
XGlB8F1Sy+Ux4nW52UHuy/JCuxBhuRe1aJglj6VddNPw+zeHKVtoJ0mJRnkrAxyRc4zUr02oy7F1
I6MDtX5iSYMTCz4gGExDey+SZSzdFRqlYi/N/B5JX3AeNTHmWWIeE4LWmHK0jeAoGJUY4JMrv/0o
JRPbgk3nQ09bkCRrAzJmbo45Pty8lVullBXGkIgjk1CACoWJYWVMHai42NsH2T93hYct4fePgdeC
Yg98KmSK6+WrBf6nnuPFZEp8drAMf/D6G5yDmibxU6LEdKBl9b3F8G5WeorpkcuJlDcyewZBqiAe
7w/lLpyKcTfP71n4/RnAXfhxgaiwXM8DoE7POX3RwJbN4jIgHOB1pnOFWV/n7BIG+56Y0R7Ys0OW
3DVfd8Pz79xtDvnt1WAOQRW8y+LJx8DbkLbXZTICcbl5BPD9JhxSPPk4zcMJ+M85cOwBjnKkoXS4
+RtqcUjWE31+RJSQVaNc5sCyf/+GJTvpV59iKvFWCp7hJ+jAFrrCDia5tzJrkNNWeQ658BMFH184
ZZ+wEIcOJzILi9VjxehoarWdPkXa1qnM8gCVUm13CldXd3weERwYuUMTgCKlcbqje5ydchExxVNp
fapyL/NbmZ/helrC6gxOv/oIt2Qp+MP63E8dpRO75d+OMC4xIKfd+l4WtODwOsqH8rYYEXGhcyej
C3dbL3pYL6I9rriiOhpMqMAI90xYDEqROR780TTmCIh56ws54jIZOxC3x1BzTLLfK3cL9nzCHMHi
6Vg96xEBcVA0CPM4CJCwxv6jgk4/wN2n39b3J77bWTfGqaY+u561XS/01fbq7s6o3jP3o3nCMOtI
EOt1AFstcLDD0Y2TVx3F0oVUJencryFDH5Vorui6om0/wmDwfGDgRSlgqjAroPPFdl5XTAznX2h9
SH+tUdq+9Z9pzYa9rmfn1VMk9UPz/9+ER0UPG7fOPNyV6r7Ik5rx/PhcoHKYmECPb03aXekRrHlx
3btLBodEuUwZVtGM1eYbuvgf4ajAvHvWj9vMKgWy1tfDMvOW3b6facH2ZenCNd+rrWGYEK+/uVSN
7CvZ7hsr2ag/TujcV9QXU1kMTKCQVpfOHf9Io9BBoetF7vga3ZRmO595J1uUO+0LZpftOqy9aE9K
UwF4Lu91ISJenRRHOvkv7JE19gEnBd4CiOCyR8EAQRFSvSBU0xl5U2GrCiCNDoHJUD859SAZ90QG
XVWZFLmb4OAUWcUwjfxzKo6U0mGhxc7oaKdWJRmqV2F5s1LVsTJKsT8Dewao8s1uc97gdB5HNIeA
0iP+b0YRzrm3tH+c/pZ1hsygW9xRWgxCxE2KWiSSOQaErEYvJGPBOwnE+EWJQVM7l0vZsKPOo3EP
pXQE7YgKomTcO9bZRidctTMZyZotqm5uzcvadmaK5E/RHKvq9Gf1j5iXgc572EKeSOVTojj2tand
1ksjQsM+3HlY2lP05rzhCICJ0IRb7F16ZcPecPhpR2Sr3i/rcTQN6jP6Sd3HBHb41pISxoJuFbXS
aBN5znni+TdCCcxY4EC8CLbYN02uPPVLQyt8Uw7sSU9LEWoVX1fLFkiFhncRQkKXlW2z3HMS7bSN
6IPaTurvHUzkPuIKXc2ylSrjkJoHIZWMey0U5qQW6hg41BpyZVdxDIQOUqUmtditOtxp8ek/YUoz
sb4uTYr1cfZCBfSk5gMiDCAhvAsETiS87Pu2GCwZLWBxFeVcYDKfx1ZBwOgIUT83PEyISZjntM36
OG8wotQDnKhtGpJsLy8vaXVurxkmZpqMnLDX/lPvDxePSXQdPN2rzBmfWQwsRPIyTH/xi4Mn0Sfl
fytefLQXlJIBhfCa9Uib+I+755gcgLoE2NVJjRsVTvKLw11dYGmFfQSQ8ZM6U3hPYLPKsAPX+FTy
izXtJYLneFNI/C36grhewdB1b2AEws0lQreHz0EQLx+ugpBv7Xvu4s/ZwRPD/3EryNEvwpjyWi8v
meexU7ImdqJ4drtOp463579wT+nbbCymF2Gcw0t/4TcIdE3clZRmks1DxeIR6Vz2Gna4oUH8msnD
DNuhl1gbKUsEX87IfWACWgaFJ2TCYx1eMNAg4iwJwljopZNG7DPlTELvv23FWwkEJpXhpeJlNcFM
NHSPDv8KSjF3tyqCDA9gFMQz1gYHySIVkoW3ZdpXHK9vqUIRqWTxXFaV2HC+Gsa/49eFKR2CoPOW
AQ6wTH9wlY3e/tmQFgW4m/jrvE+0S2vQIgezmLYn6gdMsViYKM431W3FRoyi3rSiG9OBrWcEmB3y
sOROwCkBrJd4n736Bf8v5lI3KSZOMR3bmBFf2iFHW10StyBG0rkh+a55SRvUeMMbmV87hSGzQwv3
7BqGpWTilgZ2i0LR3iNSnk3uU/qTN+Went3IFJ8Nz+/ishffCmPzmafziyJbNFA+bCZKiV4yWm4f
siyVMSfvKEWXQ4E4YmINP35D7ZyoECRjOqTOXVM82E2Wmrqzd3gi1A4yyUTMvUYcqOgOnki6gc0c
Q6bfNZgiOYF7jc8CWrr3ys3CHlml9lcgqzfJGpvTZLSf4/FnsGh2F5aIcvgATr2x6rZ17IYbbW+h
wqlAtbPuyc9/I18b/QRtpJLuUXwNYxrDPuY95CHlrvxK4wm9n4JgMujTJ5Iv64XWVuXHWFqpv+pL
GyY6C0Qd9PwAt2Nu0UlTJOUqyV6IHGn2DtvGK5/TIhPPZXYAjJRLe+vgJzagA1p5jHfBktkFAuiP
FgKJ0FDzSYSe9EsM3kojaWYEJdMTE5zLbkyv6oUUwg/D7zUFUwc8vW2Cvs6fDD4RTgj5awbHdzNZ
070L6WabdcnSZ2X6ZCn860xdmuv7XBA4LFvP2450HNmXrVimZcuq3RKtPC3szheYDlEJ1IwM5e/T
ujfWvloFVJwAOR1E+/WG+ZUl1vZZ05M/993aXNZ9Z7QKTD8Ylg1EXNVLUNqdENV9buxMVKgvkqjM
Fup5/JAoBv5ln9t8V1G2BmzYXZdfC8xuHwCtWnx//PzyZvAwEsMdrA2r8lNr02RPRzFHX6tZgeHI
ipoZ/hdIlCKtlHBnbF4MWh+AdmVd3+ZNx1G8wWfzCkhrVblqZjRvuENsQMXXZab/OqcASzfckg81
NPlmcZuVD5gb2rGWc7mxgo8BINKYKdkCYcR9yuCRTDcc7hwwZSrk8v3iy9yEIzCpTOhWMvS2lOLw
N111fPd40nl6LwIo4vl4XLMJn3wZO2pM571t5ceYlRga3o9R+Gd76S1icF5lNAZOp7TaiFtjZmsc
t4RD+bTuGXm9EeIRSk71zBWu9WgfTNs3qWmP72kOorO6uCOEefV8fJIamk1MC0H6Os/xKbnnihag
QIR4/3flfEjtrCFgcXRdKu9VGeiA3+th2bf1poGpGRlSWpndzr4+KtMmnn7Cxwm48I01qrriu+XM
DAxNjBQpdt3ZTMq6qA9suGsT6s9705S6V0p+JGvdGvR8tkpIw4k56rogRVpZz6uLYrNkr+TquDnQ
Wx/Qv8tclNTW2J8Grl4enk2dd+lPe4BQYgAkWmVI3HxAi22RyawO8hjqpJ7tV3mN84lesPG6tWxH
zMYN1Pp+nK53NzwMfWlU3iHbM5PK+ElHU8eSTtJjFBzz83PAAU3ajQMOpGcEjpB8rSw7nUMKK4jT
UvklMa09SZipJ7881Tb6o+2xn4Fwm8GZpoBltC2ZM4cbdEsi+y3VT0EU/jevZrAwtKJKTLzPDNXo
oHFCiriOyjegXNJvRZzhfZpJHQxOyFRqdi+bx9mdwjOLLIKHZ2nj0a3zREFWtdP3JvQgTtA01R7z
UOfe1WDsMfg9E4wGJUytyGifQSHQIWJgJ202nwVyv7BwO0+9ErtuAuhG/6xs3dYTxBqQnbh+587/
Zvi4qePfBaBVKvD2jKHauQelHenbiZHYKI2Gdv13UUJFtLuoksGM5CXK28CaMRdotLqJAnCXBVzT
vxZ/uqfATLZwY0mjScT0YcWEIgKZVf9eLEqxZ4WHQizaFj3zAm4eBsFiHBDRWJWr+HlQOC0sHnPw
CqTeW7Lv/PoPjjZ2HeybzKwDgqVmH8ydMLbbLPtRl9nEgnnR+iFO0YLZUytTtDY+sBBYswNMrtl+
LFiywrCZ+Pa3a5oX2AHZOdkLQgtml5gn2WXAe3E5mtDHVu/RXAinNlJ1Ofumc4ljCkeXfJsQLdS4
oTYDTpknrCjEqXCN4BUntgE7xUegPxdzGa7CmOIGB3bmU2Y5vu25bGN8VY5Ds1pkNFlOhZjjnj4Y
DhD6rBrOmPK/walvsb1L54AlJ5dingRcp1xnLdXAyvWNZ2Ao0UgTW0b63Jpm3BexKbj/+/gJi5l6
skxb4YQBaICOSjcOHx7qDC5fDnIoDJCZYW0KuOOfKBbOhqfC6O8HQ9KAm1XgHHsh/rudwbP7dtKA
O/5PXHJ3oCC2yLMJFz4qSCkpCy2nbL24PMcx3FzpzmIxRbxfQjvHHb4zfE8z4bL9bzhYbLx/jcbM
YFiLQw1EnU8HVF1Wv561dwhypFLrbb7E5c/hWnhyJN0XBpFjxuIcnnGCkiWPclQs7sBPE4P99fi1
b35pKfDFfK08+g+30QrGA+71fCx9jrCqFeYIw/w6PK+KXrlOdyU/8G0xta0nQTa4fnv23L/7cHL6
mP5HbBbeIH0cbJEhs7HSaO/IZCDlHEcF7cyLjp8MBBOPSPB2qsGayPGXqqe+lMjxyALyCHQY8kr9
MEdUKixVr+yR2KaSi5ull3fPd64AsEpf4qtfkU9bhiGRbxPM3ELdFjGlKFMwjZxA7hXhI/3RTJ0x
3uW4z0nVJ0GZDs9WAmlwscfzMytKO4TErb8fu99wiVoH168/TRLdtax2wn7F1Y9eN0vi8zLvsOLr
7m553WpyQXIxKtgLczFz+/kaeKLG8E8DUYHZJFIH0XgHHMy75xra11i2Fu0KlgchqAwhZIdi3+kz
sg8HRuAy3YUEzdI00FsS5ivMcV+gaX0BMyUREqbQcdzOLl0bJfXroRGaA/6JFDlaT9yrsbvxCdOd
IS3zziq+G/hMPUBsA8y0QxO99bt/+gpoS99CiV6LpvaIyng/ysZC027gb6XiHp85d7XZtVyuaP0e
t7Q92N+ynlGQFcphkBQ5PFqjnEzwPNpsBVuEvTP5o+90BxyXfJNdJMUWdiA0vdGkChaHz4mB7h+D
sAtO8qXqpi4wGpD1WQYmpNiU3v2GY1keI+JXh79Hwat2ISVqIzZ0I/2diWCjlOwkSpajtmsVgtTO
0dyvFEvL0xm+r5jC1iGQdPC8foGycwZpEcWyESZIJCNnjebf3bxVpe3OzyNgLSSMrsxbRfSPCy0j
TPkeaAOKQzhqzKY/8nUzso+OTMyZBdZGjgip83xOksrf3OanWUppbIX711dBMMzwaZxxNmwH1RIA
bWsKT4NCHgLNCau5dO4CmFi7hKrru2rvZfTqy5IWAVCYPX1pcSf3M7KgxMgCrjnhNlUE1bH/uUaO
qu6u9FFuJ2Qb8Z3rjYVT88+KPzb1rBm1alWlSRTPWWCkbRplMENhxG7BS+JIKbgZcI7a9iKyMvT1
JrL67Fankxv3AJhO9mFAkNHyVFQB+K5yQgLe7UUN/HcR1TU79fa9YwS5acR0l5ieONVHDyYL4MPJ
CRO2Bbz+dSoHRISxdyCe8BNq9I/XvyH4jyAiQDfjTzE1e063JEbljF4r2SigFb8WyLKZsx2ir63B
xAG5OP2kKNVkmTvMHPoKeWbYfEN2BXHT1XE8JuorUFFlmn7ULTXD/7u0HPk6J9cd7ZgMJcw40NsL
kbvlItw64Hf/m6u5MiIow3JwM4MFMvWxvHQ/ocHfYbRN2KHw/lY5PPf2E1YljxD07ehByJiCL+LL
oD+UsQIRy2oEbMD9m1tLkOeSrR6iqypUQ6x59zEp0gr1uPWO66SDVuCMnH8CCKC2NQRmvGqKgQKT
lZeKwCnnS8tqwxigIzQRbb1bOr3aS08jz0paytf/Hm2PjVGLJlEcAkYGIsIPqd/Xmv0vPjmeMBR4
fVOnRiwMkn22uo0V3lAuEetYFGVDQg/5G+zreH6z1b0/YE2bnbFqfWwiOm158EfLydM5AN3qDFkT
gWiQmvJNx9HmcuQxp0dAgEB52UzM8sVo30wiwjkaHz4gko6wbJu8z2R2hp4fN+VRNC5978ueOz78
ICcZ15DduRMpo1pnMyosak+L606dB+yfVvg11Ax8krj1l4vx2XKptuMyOyNHNpgEUEKHF1m+Oh2j
rFmdC7aqMQ3RCpPxCMy4KOtJkSHocDNcjHoKo+CNnUkLOCtmAOvoyELLR4W/MiJfasED1nf0i9li
g84o5cLmuSkldhhNq+d707RFNagBExrRcbPvs0oJyNCiChnpiC2r9wgRTjYNEBTXGIXItGOjhzTS
EoONC4ZBUt1m5tHfCExpq/kdyxl3n12ewXj5JjAiwKSL+0hX/kMAINPChrZ1p2C4GNuccRRRPXaS
VpySL8yMZEFiUTwqig1QTYIMNKoHa+mETSkewzDi96H843tEL5GGhgzIokyzVR8NKXlHxDWKx3qx
pQG5RAkfDDBEtJZdMfO1fYYvNsMPrGuckVdNkbtLwpzxEtc9diq6Gj9atP9KNwv6v4ZhwxG5aQpx
AcbSXjl5Frvoq9mjhyG1LJTYNa1vuz6ZkuUEJsSCJ5EqtZCa9iYKkrwbmuiR5ZCWnTBNn3xyjiY0
/Vg98ujA9NnFasQ3W8E+aEA6ak7WPjS0DuLWH7K9R4aetMBYw3yTxaDJ5eueWp6ewVLmO/zSiFj9
rtbusYJCjgPfJN9vLbWPlF9bvQ9vTIW2k3YY33fmioEvaI0AMw3XXqMNIDKY58/9K1+1su24ViOV
Wzs3e2jm0gLcyOcmdwNYieZg0QSs/oQ31hyeD4PveO2hMR8EE0fNCUMAVmBqOhWHPiaql/PzjxtM
j1hI7xVLB+OGMD5RGUDLvrhwpFF9v+VlbFsXQD0SjY6pDeHEmK4zlwlGAL9mGPUR/ENjIsI8S41z
zXEzSvFVgO5KAiuSoWmxFnA7yXW5gvoxa7eFEnHm7vNO4c32TSF3MPb1s6bWc2XsU8sLn03uiNgI
JfDthSO5bFrlEOTLMN40Kls3SlN5v0j1x6aKNC4havauQhlWeM6Et0/9VMmPCvtUw9eaLNvOq7ry
1fWyQEq8e4Qp9hhAFd7NfQ4Jhh2+AWgWe99aOtSWWmeCNQ2MBhZtY5gMdPoKCeUNRe2KEy25MbK3
2qvt2Fxf1ohIBPALaeUH7mZG41nMUcU3S1Rq9N940jCDD5aTa5Brn2eeFQE3mgX6I0GNOesGuzQV
zNj/Naz7WUu5puTIR94VrywBWtpd3DRuRtMesV8xXRWhL8s0YyuunnByzbuI46sriGiTJKGyV4WK
sfrEUrkatAPrB9A+wG9R66PMwiXA1V9KcBkidtyNRJ+J3NE3Sx4Fi3KoWWQm35e/b2QUcYmDhYSK
fxzkHte+2K7CmS9h/Q6cf/Xur8YViVmK5ZQL8s0xfEFUHsz2j1Z0rLFl2SPD/mRvVf1HRGG16StJ
I1hDuCEpDAmEnIc1iGq42CquD40Oo4WgiZT5OfGpSCJFbkBrJVfr6jah3OKvcK1iHvPNIfPVky47
c0YV1GKUqiXst+eBgXFZ+sKeGaH5rIgYawrNO03P1KrhH96h0epzI04pK77pW5SBavOQchrAlkws
uuYAHc9C75b8a8CpSiyy/61f8zVFaZmFJlX3DxjoP/dIZxIHons9nzyg5Y4B3kOMZVaynSoVczIZ
Es0iCKgyLXkB4NOw6BDhj1bwFSGAUU6S///ilJa27OofdxBn6s+rpOpae6I+klbyHw4Ih5ZMr0pT
hp8WgjkiZElwaHd527TXrRY8ekoHCClu3nRCIkqBpUbpec5MtIi0EbckpuNf7eeb+S22lt1dVRV4
Qec5k1+HpMd71XnbHUf/C8yReMesw8Snk9fov31NXoVvo2Z4ndWKBpCIL5ja+FySbNBYxx7pAlM1
Mf2aT0cO3yZP2P2P7+khd3ts9PcJLOCzEhPBGtjrsNTKFs+wVr+kEVhUPgjZyUJKA/1tb9rpoY6j
WAlZ1qJ8XPqWuWgoDzJzMnPut7lzYteeRslctlKqkC5A7vIWv9YFlrq5k+f7VHMDr6z65bLWVB1r
wCnT3Hx7nHZAB3A4b5MQHOZIFV4wj8BFFt5eI/vEGepIZ/TVzUA+ys8ntF3j3MOsBtA5v9fLfRE2
8JWy/ojwIg8/LQjOKtwb7GpSUuTKShQ//zDUbdrY/1mGQyZF4mez6nM+DSDZQKV/UGZbjHZYJTe2
0ekrbEMqSlq/WYPHdqrh7XC6BH7pClUKtGbHAbFRgwlT3Bio7C2MPQaKSoU2wfgOPgF5YLcC8Mte
GRqaEvWM5BkWSfbRHQpEVVqsWjMUPB+C+tdyZ/5VizZC7f0aAy572l9LAfJgzkrkeqWQjzKjKud9
ueKu2o1BwfN9EmuRDdoX6F2FcS76HGUbMybI4egAHOu5T616WzS/LrIygpstQ86VP0CMxufTZfR2
1v7IWos46P1V2gY5GdhU/7sPOkLvB5MhJNDsMJQodiJBXgWgbNmGuPu4H0KXJwpj6iMUkrW+vKZz
iet/CqXDR+4tVE3XOI33gdgXCDbCmzF9Uy9JydHXO2HiU4muUund6xXkxbYC5VgP+0aypaOsU79X
x7eWThOEEA/9xIjlRsRN8iZwRSEbSU5meC1JsCWkleC+JJxY2hQWU1VvjAoj4m3qJy6+Z2HgEXT4
Y2JKR5x81VRysb2p1yZC8qNcNuyzanO5yO2OY0EZaXWcqxbjMJjtUVmVwuTLrqLJJEO27KvkN2Fg
1ovYuf2FgTp51IR/W2bEuyuL24GBPAq3MBxqrYy+WWFdZUbD1omXSFlhxZvT/7hU0mkFczJ/bMQ4
+dPOQY7Zbax/fCEjj0lq5C1eLgvbU6WmSRQECdxzeatALLeFCbitdEyrrLSM4qSy4Tpu8+Yb3du1
KxSm8MyaGMcKwADQMYkSisqT2g0nIyz4HJPEZRLuDlf6Xkj6uYv0ALRw1r29thXTf8jv9r+stmUa
88ioM86DvpnHuwwdMBErc2poTWSe6sapmXpUMukdw4smcO7/kuug66dq9usW4C8zgWpxfIqAgPI6
c14pDoxRH69lKo5uY5N+OTfFPnYUgHbNfccNMFIovhQKvG1VCk/PbNiOWJ6tbmS6MLf74r+mI9Dv
VN9WKHtSem7m6PYNuAAOD9/iXk82DcQEysaCnfOoeG2oZC5P6NzkGtTb4mVmXk/FdywAyy/ZgtdP
u2li09atlJihZKO83BNsy0DiuOuz303UN8gZrIRxHfUCwxLr9adDPhZ5CQG9jO7sXcSArU25Ba9V
hgA3QwyLzwjsUjgMbgXwLD80AR/ML2jNrdY3VsuZFQJxA6kh4GN/IpYKICT8rdSdI74C00aOL2aK
2AFEWmHf462y0UkS0y3PYZjQ9GpXaikXqvDjOUTfQ5rjV73DXw42++yTk0+DD4qUBS55aEDdE1oh
9AwS8qhnj1xkxouGcWAv5PwjqP9e1V1ksh3AA+yySJrZXntV0XkeN+Wdgy13HiI3ItaynQ7j5PsA
hB0YeYolqKhhA5TW3q1HZiaQ7RCwIEoRRrCy148mLvtViJgOrIR/XgHKRirtYNI1ok0izb9pUP2U
UeVxrqZSp7Ott0nInuz/2Jmg61YbK8SeCy3MLVxWVxU0t3gFOOIx3mGziaKHwyAFV247OVuWIAKm
wr/gjn8mTssuPvX2uPPZfGailv8Jbjq/3DaUYGyg3bduFCq3jRYc6ni3O+U+DvF8ooHqET0NBYum
yuLDPGB4EaYQdPCtZf3TfKTihFgeyU3EK6XVa6e5tPj9DRd7bGSnuc0nrAsOJcvRAgpLIoDLppcp
glsCnfRZr3KzBxUZ/RvpmvFlnWOBqaGMExKLNSJ6loHu6ZL+aygi8+U9bj//gnGVZU0mnxEEFcRR
b0NDWLX7/eBLOo/J11Uw72ZryxHd+5B1kV7pHBUkbFs/T3vB+IIT8xkYLwPBbXe8uMv+UveAd3lw
FAaOyi4uLZXDvgerKyF8Np9CpYORzD9wGA87flA1H5rFKb0W4Q/Pnw90FapAYI7G8/i3b0KzjHlT
UY7dPFmV3n+MdLUbyPDo0Mt0TMv38Z9DpIBfEUz3zNt0BBIaxkHQzEihni9EK+8eTICluy85QISE
TIQkJ4IjRmpXC2z3Sxjni4PnIkcC5By8N3jqGu+T+yLfp2eS5hFOrZt11BQGkqFBkrMbSz9hYJnO
7QbLUji3QO7R1ERVp71mp0Elr2deTg03+s+JbjIRgT9TSS9cgvn993j0hS4Xi+FopMyiIWg4e4dJ
5dqglOhvt7iaSOuWmY2crYLxPTz7M+0Engvw28iRCbi1a2NOd6DCEGP/C3Lp+klLqxD4utuwFiOB
ZE3XaAG0Y7y1MtuvGclWUIUhTN6hX+Lc85uq+aZrj03S4I624SxMuMHDGbgT1S50npJcEpN9eI4s
KHIOYHXTx2mP5YznR2TmOxeDdVc8Csv4C3+FPHfi13yqtOdU/h6TtzJf+GEgQ6JEOvHhDtdNg0JY
ojLDBbcwR45uWUIc2CRULFjvx/jGksjqGbSgC7+fzPLQLC+TgnUuOUgoqgz9W1hHUfOIUQLMMHEj
xB/Pxkodnyuu8tDSHchW4bJY1lJCUp0COSZWJFOUIGPabcnDoy9beO4DsEhlKN2CWw2+bTv1MzNN
4hPmoQlI7hjuGWdzD7f261rxqKitmMe63LFanC4CJJ+mgTvWCEDj0ibZdZuNgwq4SWX0aiTnDsyp
JGpzZfR8jtvoddgOD9PRKFDWllQOIuPTVsdOLefWQpGCn6lK0XFB+MidiLrDiEyTn2XVS+mT8AtS
ZeJsTN3B6mo7OdSPdasA9oPzt/1cfmneCQe0+mphvYTK6y7VvtUI7FaSK2cdir76zFWEH6NYfnqu
mKnUuGvvQ2IAe1GE6UoBciNXYo4RiCwWjOVwDRiTXlAO6IDUFOA8x3sLY24O0mGdtnxruS12QDue
qW9U87b3uWhEBhU+2NK9sRIrhgJzgspcpaNbqpOzk85uCN1L60Gy4+OxpiKU5Co7FbU1UuXsjeo8
p0Eq/zvhrQPA79iBLCxCYFiZkZJHqM1sJBi0sWEX7iC1Q+48t3DN61W4RewdtlnKvZY9q4u7pM1q
z3PxmiQBz5nwtzYkNMyd4/edpXfH73DAzb1xl7CjwKzC94oszrcW6Llmr9tOBVFe7SMyw79GGBxb
0zkaPrtry0mANwWUuJQxn4isbJN9SRJTvMyZnWAn03H6E6BOQWh4h4AuZ5ZkCJSrw9EFnP+VY6is
THjjR7hUOTKvJs6UuC+3yxiqbkS1NYQ+/pH34Ys28QUK9nWh78BFYwVQBzRlpYNOlqhNqSUZGN9/
4armR6RVP+KLefGAE3Le6pdytJwNmkIXMvEh3Lp9cxKMFchravhv1Fuy1NOd+1glFXUQjyOXlCKo
0tqQZH1Z8tDXm684lPOhmYZAVRG0MXyz+Gx0JBlXa9qhvm4De0zEYn77ArkyXFyjZhrsoYfh/iGk
B9R1TL+/waWJH5VmmG3DecxoWuYsl2YJ1bDJ2HJuZuSz5VUqVWXegnmeXoQkgBb8nKIiJ0qAvIzQ
yDhSI4Xkdi9EvOrweg6Jq9bUiy2Da/D1KEWjbF1zBx0sNhWrxbgASqDiWP3dAw+jqGzZBbsjhSV7
EHAAq5jZ1JqZYC0e1n7ZxRc+nWvmP1G/YqCGh3Q7NrUZcDSCYDS2031BwfQSYUWw534Sfe597k7n
3zPOOA3ayPOXsdmgDMQPwtYjE4rqqmdzKEF0cHOKWhXfuC5It8GKz2a6+MNk3wAhpGJdpw+tm5HM
hgs+8UrXKT7YU+J027Vtu38UudFaHDjtugdM8oath031tfutjMzlHU3dXwVKIUMuRmneuH7QEPjy
0nzpsWvdGNOVNaH0suZle9W1Qr7ew12WuLLRxfWt5p1z+CwS9iLxNhUfmH2oCJmhHGojNHkZmY83
IC8RKKvSNDUffuLbO8bZicxKzF9uBVpk3u28k63RSKAYffKbhZJzQHyTy3m7O8TXsFut/0ZkinfN
1NV+otcO48hIk1X/rK/UHbTJGmkuWALKQtKdHxHM/o5JS3vqu6gmONd1d/ZFzStGZ0/V+eczZYTN
f/J5YqmSissP4xPxgYTcHZIx7kFh/pmXKoY4URDwKNod/UGOcTcvgVN6zr3olL2vdDFKyzZEjyIt
MVX3/+UnmUsCwvFAwmbXqXqxgdrNpicVl38F8AnYpbQDmfVEBMAbaoUbR3Z0HUoekWh+3H1e9k85
yg6ppKVxxQN5nvs/UC0te5NbRKzsAAWiy/R5e/j/F9X6tII5xBHByE7NdzRvIJrIrAC+7KKZKbQb
3yDK8p0D/+W7ASa5oKHCGBv7lreU4xtc467gD7pst+oG5SET/TO0U/SdMukauVuF/8OklMBYEy/J
ByfMUWmVJj594a5QgNg+p1cgYJVukYEPVdSoZyROOH7csrUMUQ72f1YdR6ETbjNqpfuvdnCsrb/8
OhciDgzfxnVTadwPVKMlxexMspxQege2k+/6vfcHI6Eme+J1n1DkeAmYRgdDRGDGHy1nqe1XOH2D
631ZzJ4yvRQIKKhc7RzWnTBs/fiPO5J+jHI2l1HMWgiD6Rrj2HIXIRL+LiwnFPG1GiFmbZP6sSzg
VAhh/I3hEvbQkpnMFZIpf3q73dvP1YVgPyt9Rafzp1OnsGoppJre35Hvh/Yxsc59oRrNlQalc1NA
pQJQ46xEo7SIJgVByZgZdeje8a+I+U03xq7Z1TN/aVwFlzKDmdDU0GD6Re4YE+zerr417WKVOzXV
DI5kDIJC4/lrTBb5a3wePNSkubzEipMFHZO88FJgCttL8QmJxgYyOjmogtbGKavUReTwjwMFd4Hu
dr/qdoNwc72qKSguvyOJLt6dI4LIsTpFNmP/ljLG3gMfK6o4aA8xW2ikBOCVg4WpBtONl7D4x3PW
bWwU36tIP9jqV/kf+HCbzX/mPyXsb7lRFzM8fk4tkk0sXskJQHVj57mfL6cI23TkxUSDlZqVGRuM
zXj92fv5NfN4+QG16hv+pkmhVdhhbt3A3tvRVuIObs9on2M8++v0sS67IYoMwMF/Scqef3z6/njS
8R/1C+z16BavQSA7IWaqWyiyp+djjK5M4UCfVHvUpIXVa79ve0fpdHbCHb/uz82TBpl6Mtta9v9P
T4eb6y7o6yZouHt48Mp6I2T7uM9Blvb/KdUtJv6mLgH4laGdXy9CANfvMq+XGYY2qA6xLqjpl8YC
gGoLUtUFG9d3vO33fUrSA8oim9FV54AfoU0oHghV+Zm8Vue1cqKDyB00CBBcV8yzNJmcDOFuKosY
Gvei1M1QuVtPhWAIkw5XTQYUgzcZysa3XuZ4g3SbqhG3WctK6TUWEwgnHgIiWyOLj7W4DfWbLzJz
UNkPRf8z0l7+/gLIs0SzJLUP6Z+8DQem7zKBVoA6jfkJYwzHQnLicKfu89k/bsBpiRsPApSLHsFy
QnYevaC3sEBfr2S99qmD0d9i+/iVOax7NNwpC33agOgM994wYJimCeE2+iOeTDNhBthFzyngoeJT
edvgNxzfVwGff4AS77rrHmYKNh9LDCh+Ex5Go7qr0E7XYHuueK544et+ZH1j+w09yowOs/W4aOvX
u+6PSNuDtPJtqNTUWN132jIT1+nFVTKl9ci+YWzUatHrIULeczYfAW0HIkX7//nu5HMNL9TMaQBH
frFMoxUYFv0wUKPw4XXDXLQLnUrqr3WIiKZyFXxRH/Fv9ql5w61/VSzd98ACKs3Y7cIoZtAvMOtP
Na374BND6GPhx/CzRSE2D6EHPXs7nba4K380Q1nLPR6b/EABv2UQ9tEyxEo9nu85p9To8hWjlgDt
qvJqxko9tKI3Zghk1h7TpJmLwiX7YWsaMMbCyQS1SOCBPbk3iiuD1AvgHAK5oXP7iBTWPpNPWkBz
m1p5xN/hVow/OTLl88aKupwvHlyMnsWqv50YmHoGDPkdCwIsTI12OULRgeIOw2iumMVJgfkc2H3s
HnbBumWmoXprXBDP4ZF7tLlkuk3U9PWicsy5KfLOiXiPoL9n7kz5R8wvkw6Dr+jDirf1SC7+iVgG
fhStyJD/xnff0I/OHpT5Af1mhoC6QMARjsmuYdBhpKWqi3pvQBzeQBlOhZhcFpKgz2AEjd+KOgVM
tnHG7xx4lEbkUzkDXKIniV0wF09MC8ZtYiKX6PNWS/jqBRM16ami/PbEV+lEg0oLe9cEs8y/T7Ny
yVCY4XbJSkdNjnB8+yET/5IIPDMvJrhn/S6FI2pvQsf5isOyRxUCV/a2OzQKKm71NYWRozVJZ/0b
FauR9GaG/HaLzx0PCTv7iTLho2E4QuhmvcSA/QRQc5byEiNj/lnZKWYN40hfHBf8BABpPNIZbNRo
yCy4sTcFcDsNUid7Hzro87XkGXsiU59HjtvchewZNRI8UBVDFRO2JUE/YkLniOQ8xPGF/zUACrhr
8rkEGqkHaYKCcHAvjLjwBNlZm6bOpExqJYuAZnK4vsyEG8gZDAi9x5/CqiRVL5oF/MlkiHdUkwG7
ANgy357ts2+6QCjZztV/tvteO2H5zCbaceWWFlI5jxQULp6S+xRmMTz9DT26Skhc1O6RpcDE0LvC
4rUZ6EWnDD2xwmOrQ+WUGiMvBtdItuAB8IM9XYlJlIbk+Bb7xLFpHo8eFElkaXktf+3bycoZCc2Z
83YAuEFowpRMQY9lBu+v65/KGa0GewoEBxu+aZA5nSIqeXz1/7YFNBqm9LPmRTsBf2kGLvA00SZ1
XoT2IQsO4dqEaDQX9aKuvbKq48xKyIDq13ODPXmpYMYZ/N73BhHYUFiaVlRjIV1uDYysNOulM7Im
WRZMy9PmcaX+M00/Ox3QaRRoAeevrS9RqGMaR6iosIu/AeffQgTPxxdiyUsOK8tEjktc8PDWFIKu
DZ4DPteEYENlmTbpH0r+O9J/hC3MHpVcAavHt3+l7Uksmyl9hCPVqcDsWDt3gL6nP2dgykzphShy
cwiB8YMM1I7a5Lb24/lT+/EBYT44y/H9p7gt2lkXvCfX0vix+v/e3D9hIxD3yTZSPkcd28w0IG5C
yNAUcWecX6q7y+imfo85+TEyB/gllduxKxRkyYQQSd2hjVXluTUEJ+Vw+yYMdvVLL7+VmCg19OC6
tPSSJzfdwyfhwKucfEnBksd71Q78KKveDZwO1Q/fABOqm6i0Rs+dVHQXXdSYKvEFHB/IT9fTQSEI
zmtzqBe8urJK/WN9uajTS71znqO1Bv8zg5yjtUz0/OiECNbh6HGBnBITQ1zM08fhSeME6JKdPWsc
GTJB7GbEkkYCN6u7acG7KYmnKxq6BWA+PsY2h1VUL8w7syNfW9afs2I57RpKjuUWkNel3Vxq2yVQ
rnU4l6FXOiuHXXSC+fO23fZMaIcvDmoK7g/S3TLaLRyfYISJQJEluSwqewLkiFaPcWhDivcCMFl+
vyvZFu6+9mQ1Yu405Om29sR8w7uG8Zvel0oXewpjX8rdvaOxBsnvESjN05zXJTyAWRl9NwSB2yNJ
Sw5ioCeXBaik3J9LD8HPcTz5a9KuXrG9p8gT/25yW0BWPePF1nYdaHnkZ/GcVYsUBd88/0Gf6tXC
ii+UpE9VciKdPnXeGSLH+RkNAZYYOllOpFc0wBtO60UruDK7Lz6QhswpEd1MWS++MpLTX5NnPCIT
GRGnL0ZOnY7U68ey8ZsCdCn59A/4G2jydsyQL00FOo5y6yzZgGE4olcYQENHqJsyCbUCZmFONVca
wmQjH2RMf5cBeOiwNUBL1WajFLlx0QkaXjDI/j6mKVNSuQ3xgT08v65cWsis5tWFXGlAWScHYeLj
XaKV4LulyhYjjSVQi6uLv1AY2WdhmrXf7yc/qVqbaMcmw0u6RNnYt370au9P2YPF0dw6Xbqqxn3V
IkrlcqX2ZX0DuQ+Z2wmmMZFrre/lcDlf+IsFAUCCN0raUBK8uU24yPpoepSZB6K0WkHFPKyh7upX
QQWCqJIvWhWVZxq9H5nqWbY4dBEE4eNtro7Cwflr00QR1fmDb10rC0g06jFxzKbCD/Pz7ed94dnM
vyjkwbQzUSNKl/lt5QdjswIS09JIfApW1J7exDFoHgqBzis/xrnfCpx9Nnp7UsoNHOPQ/bb2I7o5
gq4TBSAmW4/FuAQo1lCqkMvF05Pyd8LsW7kxYFVdnncWQ1ZpWg7Lfb5hqpVCREqmaXhXdjDhRBUH
esTu5PAHNq22DCgfYLiQWwEbEM/TV7PnQFgCM9vSbgNYXvH/bPKkmN/KaXSpn0BuposNPRNJWoCj
33pDhFCLOtGLsGSuJAhSJJDcczliY/Iv4Z2adBKkfMojebgktqQYMRD0geHoa1yCNAek1mB9tho5
K7MgdlUxYlQRAUUTAGyDFjmysz/BQwfdoKsKC9htcMGq+FguUUgGYMKHj+j6eQVrV3mZ9m0uC/Ex
+AXbXxFzNdnLVRWzlpLKbAAnuJ9HM96kFi9f6kkPkN6gLWlnZUCpr2xYnXa798PuaY/Y0CXumRpa
ceDAV21+ziWRUsuqplWM8E38cbCEcAKlSn+RUeUi3Ck9Xu/7yU2QFIcIiMDhyJnrzBNgryhKH1RE
d0qWo76ZyN1XH+kgTFQj6dfKOEr+TlWy1lMAJVvDL8EXeFJ5Bk+lEP/yUl2YopF+2XtWKTRvLo3Z
mldg67jNzz4VTpIZhVBiLUigT9InB75H6X9UowNR5XytoJzrgMhQWMgtBy2SU5EPjSjLJcbGjEiY
UU/VdzemvRstsHnYLC5qTnstmyUeHWpw9VGYDD7jPXjv+uf+aPSET537l0a9MHUyS98X2cMHWt1Y
bx+c4I48EWqsxNbzB1ttRsFfQyn/zVzaJwORKTcz+o0xlydcwCwUpLP2TvzL90k30STwk6QrtBi8
TFL3tB4N7rYaZBjz4YQvG2HkCju6xfqHPtYSfd3sfopbMGFddgmEzEVD6sKgyNwGdZdTnUngJOHY
cCOPU/UxsHKHzXKfKBIHQGdiE1P++BuNQn/A5yJYjsX1N5lU2W6E+ZCgim0Esd4q45SP2l6OyR1b
UgmzhgL2hM1nm/geUPdJ6c34raah33urkkRWpZixROLk6HEmGOhbCBsxv5+ctU9e063c2NiEmuDZ
B+AlrXOycW141hKtr1uk4Ow9rsdqpyc8qXXRrljCuvhjn59DNEj/mrG/fRw2rFTotzKszB9OS+EC
HzZz59rK36dwbRfgGzkVMDcTe3IfapVroueygCxNy19gMfkB19rwBVXWo6vcIgKqu1QafsKkXvtt
TV3eAOnk9yWw8uiILfh6G3SdS9PAZ84ni6IRDDH5INU2XVKCQw/w9ktCeCMucRpqko4xJpoeW3Nw
zaxfjn35eUzjqt8ZlMRi5OwZtthr0tBD1LidFNcHCGsX9fdwr8L0+pkEpNmFyPO6iNhrSXMIqv6b
XPwbnfWrII+Q/dHvy81rVkSvfvNVuuymJUTqGn/Pnk4KEicqGAqZ1S4GRRt8F60o58dOwD2pYOmT
G46Mpy06odJH6TkKmfhICzo/0Yjb7bqwmviMlwcX8Ce3h0B5/qD0vYSVRLdp9LPzYOAml4+IaiKh
9N182BgMJqm6RJMtpMu/X/i0R5L42WWAdmLL9vrHadT2myWfQGEHwhM+MXy+uuWkBS49DgTXOmvS
AaaZXHDEilRONZrqMREy1Nms7SAJcfgOaJBQ9m5B665oTik0t4bB4B5vSKs47KsEP0sZUCT5KH4n
7lSnQzkY1J1jLXucKbkSfDni3OQ+1PtIY/EP03Hdwv6nx8ioYqmsgSPI3jvhgyZnomTKJIK7CaXL
Ot8sXjPo91IK7+f/kPy0C0bv/1DCxKM+JtHIiX5/FZjd6Rau4mp1h/34YnIpxOmAmcVxssrGygRO
eCY285ZwxQWXGCZinoqOh5UWwlpqYmtujjqXBY8D87Krtp0XB86uclxJR16EBMprAQxzvoJccryU
r19OMeelcx4l+X8kGB7SA76pbV9ub2GbaGFWE04jCnuNymw0lLEdIbVHSyddi73Q+dP9/Tox7ytg
CBeIanMgHAXJzL/aoCOSnXyznlELiH7ai2oS8oe03pcUXxFZ2dnZ2FkT2ERYbov8X/Gg/d8A2mD3
0TjdpmWkrCQKgHeOoy2dltAx4vEVGHMjshTQEPvGKIY6rQMnzJ4Rbztwb8zwYyI2VX9tSnu1RPM1
UID210HvMNFMgDmVOPpwPzfLK4GoGtosWL8xladKr0FVsSP36tQI7COaHaX+/OjTIt+BDvF45Xtq
M3IbSpzKJbfICSqMDT+YAoJQPPtKsEM7TBOlC8SBAfkkA6Og0SAd+/0duI/lJey8k2IqyHrpdIcv
vNc21uNdtPcATj/ytO2yAsXpA9rmlVE437Vps8oxj00b+EzzGmEH6ZuRac/qbZwAYdq/WXq/T9Ra
fS+c1e8RlIbh7WG/RyOJAXZ4FSg09bLH5hgRiM7Ks1uO9UE+9C/57t279q+TcEPSnp3lgpZ30tAG
XyC2zuFLj4ZS/vlNFqo7fztcIxwxVOPAyrUcxlxAZeg8uaSxYv6zuEMzrC4d9Bxpg11chmfcopXy
ZUtt8KrTdmUGbhPeJMWjAJsEWkuYQRBVqDOl2hAJWEkZh4nF0hf9Zh2GstKIw2MFcKnzEJTreFel
n9RF7p3+hFmAakK3FKiBh8UlbI0vzj6AQ5Js0PHLyReJduPgQCnFZZQ17ySU9gqNQpCyTThrpeMW
KSYCXXUgBCVeOUzCiolMXigWya/B8Rf2+atgijHH9xiCGrH6G/00zNnAxOIRh2XcduguW9RlO6BZ
YjN1TRU4iW4zJa5JQ8Pp/sEICkiuOw9WgeMgotm7T7yglLvQxg9wr7f4fPi9Iy3GmNJHEKITNwY+
0dFSK0H98JsgjVgKjxv1x3xeJSvBLgC4pJG1B084rzjgsN4JuBZdZ9+RnTlE4HnDUyCJloaL6d2X
ztDphc7OrzvwZeZDxMb4BRzywEGoIANW9/7Mc75lkdx+JXipoFZjf0XllbXVgq3+6cYlatscnfEz
TwhT7kz+1EGyOn0LIG4wEScAXbeTNu/8ELxLNRG+OEcZqs6G8qvcRD8/++GBLAq6lZzDyCxOiW51
DcPJS1DfSiFZ33xBIIhmtqK7yyy1HiYQM7Qy2XngLX7F/LxCd1ovCAAmhQ58rZ8F6JSQ4RuZNBa+
dzLPBu2L+3Abfwqvzlpo3oyCC8CmffMRh4BRv182+yVnIZaEzwiRe5sDKhRzXCVha7SgnNjIJTQA
2i67scGbgxlSkx+wlyHO6OlbU/eGTftg0C4Ed0MdRy7DZy5i4VXTtzysoXgu9t2tm1Ek5Xq1Fcl5
irgWx4SUG5vcimHAqLLPshVXPArEw0FaXpnwxtL1cnbAQciTcK6cUfb+FE5AQs3UpaIVUEslM9jt
NUPxoxOmsQxccMKF4eD+Up0BJE5GCO7zjHcfGIF8LkmwxE1LGp7mgpr0zdIhl3UY7jHwsfbf0MVs
KM6udfCtqfRdTU+48Itf4uKg/lN+PJXYF/OYXbC+W2YuFLaViQfB482UHEV4DF/tJVhHM//R/CEl
g9rGFNe91PXrDaU=
`pragma protect end_protected

// 
