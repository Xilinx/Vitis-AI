`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4368)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0ksq0VlzKtEIMmoGf771SdHoUCBE8KkGLwvgxXVkX07yFQXPGu+l+Uug
M+f7q2dV6Fo4wPbBb5yMhFMFS9PgOQoOxo8KZcKrZyuebpGtNvUiHhcAPr3sVqXSOObG03U+O6Lf
5Upx5QLDgfCZA16h4Z/ZfFo2XXqJU071d3CZympJ7j5+tBuBpu4/Lg298bOuXt4mik++aZrIZzyQ
EFPpjenIn4ihleSVuNFbOj3IPHl53ZE3AoGFVvkg+XnpUPoK6gVWUMQFdsoXIn0Ai3DbeSzGxJN/
aRlQEGoo7DyeSE1WcY/3uYy7r5fr/r9+lXthjGqnJLCVOkAHWJ/3xVCK9JVCUOfHGvxIcM/etU7b
IAHSaJHt+Dc3GjGcAMNJ4NNQw1upVHYq+7YybLsPRhJJEx7vuJqThHVSbF8MPl6iK5CMICODjQX1
EZ+lfE+7GIgK5UujKK9iHt0PxRPevhxPco9Rrvrse7p/kNsC8WYX8SiTjlOYBhT3tnjmWwLpjyfR
Wg/jNKuATXZJp8G2+wjEW5XT+u3UgztDzbuVzKeXZ+B/EYLMsO/Rh9otYHZnsWxvt0jF5WjxKVfL
ccxWk5mHesns0fPg1IxVweVG4LPN4ZpjOFx5qIlo2v5sgmt7WlJ06DrI+2VFAAQsWPeIaATtDxuD
SiSAkCw8pbNZNFa/3thFhfDlTRC1BO+yJAAJGspKKSGhSlF2qOaNAHgiqyB0em29Gg2N+Nxyqkos
Tz1bLAk0gJ23kNgYkUhKNM5RnWMry+4nD/Vqh8V/Tt/T0xjggw+dg1YR9o+1WWMgImJ55VFUwDEA
5JesHKh37W9+1bZzWx7xNJmLk/FQVJdY1WrOwfaopRIEa3Okw3OUGqbqQATIdyCOeTbNbKVYuEXQ
R31My1L+q9WBOgK4FXn7VZxPnRy0YEsGARxdoKSpfr5riL33NOgqWfiuqMt8UG9XO2Ubimxv/vQD
1NwPuRzCN60pOmmQaveJLyP6S8mLx7E/hB4X1SuO4ugxYQSiT+VjTMbzLkD0qfQn4fdTRK17STPj
Rpy5Z8+BZUhnN4biASe3a4qqcf81gwmqDRxNx4XYdOfX6dd3qqIcjtdJIdrhkGMoDwFS/IfNidXw
ApTT0/gtd9XfKoVH8VfWhIAjhWBH3kzbaMAi2nV4s1SITGKdBYcL72lmBZ4r6gCAqJhhhMUaWnns
B/srQD1YCBieZu2isUFwj9JLsOYSB/kjWtX97yRksm4FLq+MyAF0gABlG2Sy1R+kCC9AJRWiuE9b
klPEB2wTaNteeMRSV4JuRIpb6cfubJXydQB2ZHyFaeHfO+FDSpSZztms1AQZ4Xk9p4a7CVs22b+d
S92+MDMq0wWebPjaPai4fRAKH5K4TsMARY5A1brP7c+rFsh0bW+RFxEZwVRLTuVbxvsNaxynLPyG
DaGsFzPywUTaogFdpG5m1+B/8bnGyNFCWDxccj8DibTtEGUTudqFVVGxE4qE9YXZNL5XyzNoI/Dw
gfbljUy4hk0n0CzKYkqyIyAWlMXGMiNwY4IoO1WoEqFcThu/khcUoSFr56mIYfypdg+nwDQsb10f
CTitXqAQGV4KvwUBYyW4O6rrgC/bHO4nv3fK0DWZ2d4pLSoFmGNL8qY3rpdAJ51TwDbMtFB8G3if
JDBizmnsUrTOMVllYn2xtYkUFa0kOFUgvT1nLPAERWA43RSn+JNDBBvFbvmA/vtUTNU2gTviTDBQ
lrxF6DOWeZZilA4KsuD2OCXFfJmYEW3Tm5mYuPVpkOvQd+XJ+VdySKYxaFzHwLTn3Sr5U6zwCsZ5
CCyp8RDYTpcUaJGgm0I3rJjbQUqjgouHJh5HAX8CyWnCx6uBA7tKxFhwIQH1rzAWm8mHNFRNGKLN
3odkqnnl4IRLdfU+amHvqlTO67j8+9yO4xOAuQ+7GXi7R6mfwyFvlZJ/9wLIEyuPEVnPEYDsCXML
qXRkmHZQqVeKjR9FiuLfNZFDNhTrSIU+fP9vVTBPezLr1Rab2uNSDKhn44Mb3HYHOqIfn9n0hNLj
cokHSdztDNQK9wvm1Jil23huQWb3i9rLAUROE/Jn//BIQsiFbfcCdZIWLNkMYD8tamnIvE8WLGGs
5GHwoMY6YXVPk7QssbergzcMko+AJQ3MyFuS8MZP92X7Udp7MDGprL4aNhKGQRv6UXZalD/s0Kwl
Tu17+7PcIS5aYcITu5oroLtJBvUTllQK84G2HxSR0q9zbKP5OxUJsSnZ7osOOxIBuRY62Cw/PwGd
azdoA7qPx8xxa/5c2rr5fcLb4RpHT8aSkYoCS2oyCO8qSKeVN+pUMXrlp8TWTg7UezGUMJeT7daz
LPgSs6WpSagYv9MGTu+9P0iXH9BZ8ty12E5a2Jm1aFYLHPxi5VAw2G3PMR/DRICgE0ovx5lUSupZ
5r7dIUiiVPUrxLhaFuM8IhHh4AKHCa5TLN1khKBPIMOdhYI4MCWCkrlp97F2Xd+RSOXRWH8Rey2n
HNyZBx/5D/2zwwY5vStGEUAe1U2bnx1H+toP7yX0UYXAgN/Xx38ERaxDVkvLCkMOZziPwt/dFL0d
02KJ0SQRoF8sXE2zRP3T+l+KAuncRbPe4vlEP5YBrg3MadtvwlHyFPa+bB03euBmb/fveHKhtGef
Emr0v1ckJLXELS+Iyt9H+DUHgxIqXA5vhnk7L+a0Cx3OyEbjQ5ytYpXiTgGXLqlobsi/p79fnpv5
AVIM05klsE8Wzuk9ZAHFdn2wnmJz9SMRalbTbHxUodEYUmy3KSV5YBJzBpY1wCn5DwQ4tH3UGu2m
z+57MeSogkyJpfQy37HTWqbFcbhEneED7AnTfIK5lZU3aZfQPWtjmKUdwja3oDII3FnM7D2P0wQC
Wz+mIf9eeZmjOJL/42K0+gyyoLCNFfVo5VcBt+ze63EnX1oPMnszQ1YMqa+EwOO+I2lY/zM7j8BV
A5FZ2dxeqjwfqqUZytwGlL8sluIs0RVkVhzFskKLwR1yPBSmRra9ewCSeVZD1141d5y2UoEdB55/
fiK3CGch9Oswzly6THYaSRm3+ihZueG62Yf+SBuO60JzM198Mmjwin20EOcFFk7aPHuGiHJkSxJM
mQMr13uthvzmWUX4H9GZqybd5so7gHduBvZoOX9KfJPaz8SpEavXdm/9FfQRKontrmw3f5TWoLHS
4EcGBRHJfu/i0Ij9r6gBb/nW1y8x/ugEN/BIlHc9ZGyEcwoDx1YkacKyz5thxGvjsW3Frg1v1tPv
Guyyn+fw0ix5MDcMcH9iaT8FF8tShdRAWpMbJcwiDLIlVfQ9lTtE/WZjFBrZmctAKJbvWPBn2Typ
uLbkLBnt6N3PqkrQIerGysLnz6qynsjNysfDDy+CC3EDGx1WYpai0YI4epDZGKe05pOrcwd9//+C
IghEnzEJYCziZlr88MiPXhfqZ4YKM2RQl0aKFkdU0nEG/CsBAysMIQ4lRt/gbuRvE4kcdDnRqWYu
IanRaRkX8g+OnfKArrWvvQClswt9lWw1UopScDEqzhdlHM3WZJCu14OoJ9tCzVLwxbHQyOUHoj+1
SxfTESkqRlJanfUBrBgXoktUbnFhnqXAl0o8bBAl1m2YxHzuMjzl9Q1FyRUmQZ3PH2RtRkF+kFbf
VwaKeK9yFtfni66bH8n70S2243IuAxO31sSQngd/4oPuo/ZKe2/oVfpdZ51UfdT6lNs9rfpqqQjs
0pWGEEcOOPI+FSolN6rHgGQsPD8z2W3IONfscFVKQaf+wsmxItUR0wsKkK407HdK4EzosXJMO1vx
OMLk1ZapDeWiGf8qs8c7/GXCIzSxf/xE7IHIWqafcX1mqxErX8JjJuMPsWVjzT74Bu+ca9BJefey
Ckme6PDryVnsjyCKzFbRRaOvRk5v2S+RCXs+qfgWQuoiidCmi863Z6tMVVj5Zh/OSBGxfKOGjwgx
dkf4Hj7azhYvqlUZelz13yB/mAXzsTNdEbZxPaFaGahxOXm20Dw7UxDiVSa/nWta8MmxJ2vRlAAt
QYPAGVU0rYMfO52OwaqScJOhahv3Rf7L6K+Q6jItdFO1feyL59DWITnkdGlxaECUjQv360pu9KAw
K2dIfBJQ3o4C7aN5wFJqqmDlNoi5f6NghI3QREMwazyss2L9P5D/VhpJumAjMvTQOjXTbxaA0MJb
jIFjC/ggkCOQ1gc497z3yHPTGmt2yJP2WZaJugQcXQi37HLsoBL01eLRzLUI/q8W1dWrHBKS8Cgj
3IVqDa8Le6YEseVa9tnIAJMGNWm2Pq6HhGOltnwMvqWOAfCllqOofpVHMs2ueXe0YaBZE7Jua3GK
KaOdKrR47iJ/nZOFLro9H3dz/lQYv8N32mn36mlPuUqcoZWqwOsSLIvAVd862D55mKn6Qz6RYSWU
sIetV2iQV9fhKrWsKxHWxgRqMP+U3wuPdnhXX7XPZWIZBkYTytyrBpFy5kT+5H6Tof4YRumBdjY9
M10eHRj6WCb0xtheJJSPesS2MkHkZfm1S7seaFU5s67x65My95qjmqMPyHUmO3iqZ7deEx//0VDe
jDZjsk7Pm3wOxYT5gzeBMesZ6e75RyQZTS1lukf25ShkCn+ZCuKTq520p6ejylyWLA0+FH1UmPyD
gf6cC8nWvf8O2ExEE1yQwPq4ErXDIyD3SZwkkK21CHLDhTZzI6FG+lIfTL7cPPUYld64mB6Y5CjF
iTh9yZf9IvsiBCx81aFo+6JGZvYZlaj9h1AdYc1O1RPHYBnjzl+NGUdKFOY1hlwoBwnVwG1jztqC
6CVBhubonqWVVJP5v5ldX53SXdpQ9D+La+cYzr/VojPhMS6LYEbe+IAZya21QPKuxYT1AOFLZ6yu
uAK6B+on1uxiEbE4YTR7Wc1vyMFRVzhHKVMNIrEx4iN2honqdHBpM6Fv/g+AGFKjhc4e5liujCb3
UWtmjFU5K2uT4j5Vbn07yiirkbqyZqQwm9wI/5hJivbfF76DZCfmKaCaRwLvhTC3ivz9vVz2R5ww
6lHOJ08f3xujWmvXuw+sIuiLej/NxWOsmcJxxzR8PbdTAdL0Y2mTp5KgPaiClhW4DDmVIG0hJOWw
zpnRk6EQ/McarpqGn6TmLD22c3RkTC+EtPhZ4hBWF+AM3H6f9bZxfpC4ettfTXO7mnGKyu/jhoys
68pnU367MbqkSgpVMsyxleyRxLIQN5OEX3pq/jvHvi0U60P/qp/8+waneBbUmiun/lPu2MiiYbOb
fdJwl9nM7sbrFNqjjWIzlFpRiIe0lHi3XtmZ9zUKjM3WO9Dmiij83tf/aueI+XnJsaJiTjkRvJnl
M6HLcVRteDMEM6JD4Mw5EJV5ad5RyhOC4EkmnXY5+ag4Gv6eDayXWQnf1M5syMi+rsBG+fUjCo6U
wLtwT30ueo+z01TTXACqX2Iag5gW+RHQa/e50GFor33AB9oWXX8yrrIBKiW+dEaki6ZJ0IfPDt+G
PRueqSIwU3ZMMqKJZUXPdKhUOhRIuZ3QXkgMJhPERCtI0ypiiU7b6kdDwWesbSO/0/UFtNLHWHme
1NJP6A7k+wnRH3xtgdijP6VqKiTzZ9FR/J2HbO+1yvqAqMKo9AA33ERnVUYxg/c8WZaik9rZtc8S
93jrpUjpM9K4knFndK/pAHY6Flq3FwNwaB8T+z+3F5TvIIfCXg3Jpat6T1XpycBVcAzLxQ1NNr97
5dFZrW2LsjmMvLmJF7FP8oQJV7lij6mnXik2MobeabeQp9BraM1G4JyTDDNZZns5Ch//fyV22+yH
ihWyeIhP2Anu7M26tEIeseZ/kT76m+oZd9UnagSTouQpMVRk
`pragma protect end_protected
