`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40064)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPamfPOr+rPAO7s8fOE7DMw165NnF4LypmOhpB1U+tn6mBrzC649bsMh9+pSlmtwcve+o+qYc
4nmjBm7sZhu41KI+g1iFFgcqsfbWK6dK4Z501tYVfDuygWlHujHKEdgbhvA27tEXcA/UdTh34fc+
TD4Qdv9SPKn4fcnE97yWBCjTKp+9l1i0BGJ5bAkAhEJ9gBTnqA6cWREbgXLD7zC7L0L3QYDnINcH
Bh7Le3/TBrZNHLPF3jqOo5YYONAHbu1EnWJlQu4HY+VClONBrQWekV3joY9m7Lafrb45Ea8ART+G
R8vddqRE/1qaqFiPwaeu8D9j1TR6vYoHtnu9E88OwZjqRwq0Xh2PJ2sHcxmO8isB7wO2pfDdqiWZ
nk/uO9+8B109s4QDXyOTh09T8WMf1NDKQjX3LfTyyG6lAiotxWBA10YPtLU4qfc92k9B18ySD7Z0
xzoKsEcMQdlnxL4hOKCtAsEqP9nlz80XtuHxo74ovd7XYGrRAz2aehy00WZsWwyyI7QhhaLm/Ctk
qB/jwdDcvoOcNzoQOoBFgYelI7GlTHTQpnuhjCEcsCyg6GKV1rkjghLnQx8UvYChJdlY4Wa72hQT
CeHLAW6BlbMy3fqpVK8HdnplfARAx6O11UDj96kqjPLT23S/OeHO48UXD7wNKsevRXrALwCkkXRb
hjeE9YoLjFJmF41yyK2H94LiWf4+vv4vvMf8NSOGBF5ZxeCgFil2/VLH3LU4GmdOVIBFxYxyIh9H
ZUGa1Q8jGeoGDvxEhNHf+VZh6wQsUjv+hu2IwM48YQyufxHCTOXNX1PJVFSQQ/7+2pkpifU/n/wN
Xe2j/Xy0vpPtllhdSaHPI+iZvmqu/W5DHY42ooEnJjwm8UycoGKYxJ+knKtQF3UbpQ3m0ZGgwTXN
WI2UG8c09PQZaKVFzsY3cGSi+TUmJQNJGi2vvbJjJtt4su8CD8XSXWtbrzGxwm1Oy5+bXb03vlk/
oYB4WFdcEA3WIj4ffQvb5TkqURrgPHxkirPGFbKYWQkD0TMZnXT7vtqvEz+XxNSJJGB6q6um1w4L
idnvNgP/S8ucohhwDj/9Iwbk4CJ5Ck+TB83GU0Tic1bMdOnQwP2TiSniLEeW5baAZIuhi3z+sDlP
HF3FS4wBR+jsxD5KBSNP2tNDAz4paoDEwFsWuu97S6RDiZUSjc93IoqKzZfPFVGXC0sSXj+zlJS2
nsiq2hdIvT/oYTRn/Htg0Ju7vTQpsET9bubxkDYdri3mT5G7Ft7zOmCaaOHeC8e4Yqoaha1NNegi
qMjYHlxAD3otUtM5oJpatVMZCDwjbskG+iUb3n5aABTjc081HdAEqRDmx0FRavdicwGGF3V2mrdL
lxUd6JZySdZbKPVZE08XFwglgR0qUXBGbbG+XaQFCro0qf8N5NlC/MXedjvjCCNcfIdrTLkgVATa
LaVmgRTIwgI90nuf+j8ti1ufAwxaU/KlOk0bb7dorYos3emlXN3+YeZDgHSdvFRGStrK5btfLvf8
nOOnSNq8PbJnZjmzLKd9Oiyw0gwmszk8Sr6PHJoHu4Ja59xbS8YZ98SGGS41Ehmt+h4RBHsSyq8m
HEwVOnRulc6D5vCUtdSmcRHowQjv0nTbjiH4uwvWa0RwgSKa7+hdMs0ypcS+LWgitHwrqbBxLfuR
SGMY7svDy/Z7G0oeWDZou9AstPbZcWFvvHzOZCTRPcN+xrSO6wUroKxZBFocbx+Qwy9NH1s1GQG7
nsS8lX9oOuB7ksIlF5lc0HPrONh2+Z5O1qeor+wztCGz6InsW6DZMiU7PO8PMCGVyPhmMROtEl6h
vgeZi4n7BIfGNXNJ2MSFhW4mrnbjZBUM9N2V+q2isoqaZ7mc2lYMbFvWa64hqBh0nO+lEP+5mkcW
e4Oe6Jewd36dMOWOKB6s/PZA7ACd17qtB5N4WBCpn71oEMkPB70HGIk9Wl6Sumd8ouqhHN6gYe/B
B/F4za8fk0lpKDZnJEvrFs89sR5Z7GQDlGQufrgTRBrTWhX3TUTVQSp6e8MhhRD1z69VgWtp6RQB
qpsl9aPnxz8jQ1/CRrUbtMBIKZcCIvH9kJ/Pggabdr/X2kPMI/EdKNA2xRrbQLVqTdgNIGjz4p1z
m7Uq+N9hzwW0R4k8Wjxm4b/CVNnlj37xUyJaeTQvGuXG8WitivyZDVtIw84egWSI+64IC1JjOnUn
Ur9fT5QoNRvBqdExxUeWG2hRkZExGiZ9u/f86IrjM6blact4a+bCH0nxLPWh1ac+tRWfDkKE/1dr
6u6Qmw31P/uc0N3ZZSA0IgohjItdZ0b4FlUQ3s1ZTVgdxadVCVBmyxYPKGqdjAAHGvr2dO/M2Ylw
DTIgBi99qdnKDJWKOHV275016hzZb2Xq90tZn8un+zu8B+E7+8JgiYJAqExzR2+/wZlT5rGzrCix
Ec6ZNP7DG/voqjEomL44APwI1Vst3p7kxdi64LN6boyVElKnT143EV3zKes9P3k5Q8Sms9N446/h
SupDRZvv3IDqM76OR8TT697JAfd8Er+OFkxInUA1BE4jVEozS/RUmohOeLK6vI9aJ3vc3iMxZV3k
0b6/60siWwDyZXFw4UuFJk8xE8VWyAUVoLoxkHBovo/wvW+j94E9mnML62Robnm04igxCftHn1Hi
w7qnsTuO6PtU+by6sOIGrGqaMUfM+aJqKnk7VmhIGb/rosLEjbnzKgMhF0XwEh9dP27C/OlOsixN
0qtrtuH3wxr0sFZPtyudGMApPlRUVJgBMf/YGeXuz+xV1R7TmbeWL2dsKlisdbK5zrwot+kAJVVY
T2CK01jOsaJxC4Qj546lJlN+9oqN5Qc5Ura9oLqev78snP/L4SEJ8fqKhCK+tfmWEr3bn6Kx7/C1
zTWqIM8nxPBenXIeAO9ucn+tJYEWVtsyXRbMOnGC6LWzCU8Tc+PiZuXipzH7Wa3W30bz2MG6ljul
t2npTbNrLPwxprHCUd7rGi62IMIPPgfVTPIo3si7TRDaGynaTjyvLl8Abx0zbmiZfWfM7mfTOmym
KuCrOu9SZ3SP24o4gxFLUws4me7jiSK8oSmkz/TT2pimCLySyXtKzf8qJ1kYU//YzmjQ+x2GQEZT
+LXEj3EL/mOFhXna2tFloblmHE+ZA0am8SlcDCFYNe8Rb+DqiV0ISctvtxNgthYQorvsMgL1JNXs
cVl0OkVXmXkKv4lC/d36q+Bv7dnU7Gq31nsR1sYIFAyb3ShYmUWsPUmMTt2d6CSB/SGKGheN33VV
UYKpqmbz2DhjGWHW3DJxcfQQ65JoX6RyCwK2mgMk2x9AqSTb++kOfEFF2hS5hg///xMIwN2CQoSh
oChSgEmX4DWJ9lwUJXsPdPQbPlPTpjyuJhGgmarZJvmLhNk5D6XzYTr47vz2S43Nn135KYQL1tpn
HmBg/TjXVuBdLHu+v9MKaegKkiic0vqStp6f77W9zhhNDu7dFx3oFkFTPolEPmijNb5EZjsSRYAp
HB2WrrIbrruwwMlCeT932t7Yc45XfJkN/dFX+aWWgq1YctTVsto8MWl1FaA2jXsK+QUvNy/4kRo+
jOyLt4D+iaDE3RKj4gSLuf8RTVkQtdD+0ZjnpFqVsqtAPeSdsyDTke8ZgyWkPhZ+7GBO+7hNIx8f
MsELh4XJqPmar3+sl/Xj+TJ2bbIjviRNKeOx4N14bWQsvLbc9BIl0vc9A/fhW5S8pMnXVzzt9FRN
Y7KTbw68FrC9rSl0qE52gskHL4kuXYeayLltPUv4tB5DRovTvGmK0qglfOs4uiixncmwXoWUPCdb
7Dz98iHmfaUlGjNQ4ATqXLbgC2JBKx7CdkRuvSw4U0yR5irboDPTlF+qmLTxRJiy+ndFKNTb/UfR
pvyohSOee6TURBA/8wWjQZILpV1TmCRlTXt4Al4sfxn16L2ZYjHVk6I7bUOFRSBwS+Sc2PyyUhp1
TkbIrjigszJVn7hT6du9sVBL1YeCuZN62eeg2wrLW71Fetbse6UHxI0EzPcojvMKAYENKdIcf+uE
78hGrKpEQYu4S7LiV4aCUywE4+OIWwMmPchQhteliJuG+zNybmFXiQxOFJxoIS4J/vMW88VGfMdr
2d3iSOMKJBuyjRBd65YcZuNpglpp5DjkWyJYUhm+O3RsesMijRBzF9fyOOf9bM1CoOCaQHwHmdMM
fb+kT1ayev2GPoYB0oEZf0Ic+XFaFdhhehYMqSpAW0cosBDuRPyabWsyfnbRZ49eFWk80QNhvcBT
q+RglHCLfSOMy9L+Hb3mL4X6OyM38Pr+s+/zemfSAsiI0zAYiZC4ve6KGKF8QaO9klHXsarUvlBM
b1KzQm8Y1WQMUAO21WdL6NjQ4uUINEWCfLqT4DOj+IKuSQT8JS+acVd2RJz0EnXxc9W0Xhn+FgbL
eSznbEiWxtVN7+4357NdFN0vIcPZqF5I458J3k5LNXz0LfMwb240m52+WTZYmQDaVqt6palxSxLX
7qu5W39ywx2OP85rPJM+lq/JpU82p7AP9AtE6IS8heyPFrjTJK5xB3hU2lv3naXjlrvYgg4gsBCN
b0LajpWtg1hWsjOx9OCv25CnUnpKvKRws/g+lGtTaweulg7ZxJiHoGfumejnAh+VhmA6OVVPYIdL
qjxgj0VFm41CKok05E3xp++FwBpsZXHf1y5tSYfgzINQWFVk56H5dQhXFj46TCCo8b1XMGKu2lLZ
hDY3fJxxp63k1Ywrx9LZCZ1MFpdOU9SadO2aH9vlVWleVn13yw0KRSPB1t1QnPAXUSz4jnZXD3c5
xPtPlJe0y7+Uons5pVl78lRn9Ms8QK1vtdcHBrPSwqIPCigLLb+slE+9VIvwKtemvLRKKFOv3752
HwTTD0E3rH1A7w0mg7pyYqAV+gajKYnB5hLRYEDZz5qr5QP6F0m0VmilLp3VWWJxRZPB8VYB0S1v
p66KgXQSSv7b+rDQi3o34BKdVOhJOtajgJJH8EeL99KmvEcNH6GnMRHazr+0b6VS+6uzqHokNGAA
VpZFfpQuR9E+jUt4fzbKNNlbSdK7sn1EnKjMxZcG962ciYJ2nvuPSE6DtcaAwK2TZrIB78Ris3FF
75wfynRsA6f4hpyElNty2im8VZZbHHPtJMZPXwQXvxq+8mJEsK1XKgd6Eeym6yp4297FGVH6TL4u
TSLZcXk3XTdSnqOoGblYgRdWpKKXYumVNPTnKCRnPAobEqoTC8QlP9VXpijdAmTa082nS9SRvxtO
T1keulJVaXqZZbNXin9BpucdsaVxACbbLyHnlCTDCenzmTEXtlErSHgn63L8DPD8Ygjkuvn2AV3H
L0J9wTawzPK36Efp09pcG2i7ZaBfcWiXaSHbbUwreJ2S21YSOxoBBea8Q2zJS0IjrGRpwx/oe39N
pnOzGPuvLt1XcuruiSVWfaGi8wPVraOSoAra0tW1gTKn9PL0PKLTU1AzXZYfpRR40kOPpS7K2YCl
+/4jP+2FIqpHkzF1BmZkKSXK/kiswc0B0smwq2bUXgg1mPRRpzpBKFJrqCUpQnR4THxjMUkfJi5E
+pxSXo82ElJBkk3x9TqIsNO4n98ZDnJrJinq5lqxcBJyi8qEWvlq4vmwVO7IOCN5yPYcnLBenfkS
98mrKhy6BDZDH+X5w5INbKeqAhCqkwZVcPJOEnwI27XPGui5qxZfW12nEsMBQjxPxFWWS94D87zG
nD1h9MVNjALX4uYHK1LCGNxhZOPtJwADtyfKizFJIIs6kY/8YG9KuKT8KPP1lfj8j94eHpmk1KTP
pcNXBODAt1lDW9UTdIMhIh0i5UH9ij+P8SbviheMW6Z+h16oGJrDuVmMt3ZVuo6H1PfLrlJYnVyE
BjtBPZSJKBzijVVh9xPjPMFVykkJJu+EoHA+uoTzZkQJ/2INbMeL1yt/Ljwcq9DrUu85GkyjCEHo
JOOwNwRUgJog9XWzg5YUbcVZ5Ovi5sDqCh2HLoEO9fQQtAwpx/OFzOubj3YvOeKQ0bhQS7VRwiPa
PdOdrf4/gINmagI0kWc9cfglLa5uX2G6CALYQrW4jz+UCa2XsvZ4XxIFOOKDs2vqx7gu1/rkOTDh
FhC6PtxYRzkRzx3jOUB0LgDmWXjT6DYwfs5rXW9c4PZRDfF/7UdzY9nRNFCM5/PbKo2tFuBlobh+
z2WX3G/stRxVfd0E0wC9+DOe4IdekXp1SS+u388KXB4h2tQ+YC1VRYaPYE1JQiuyXOiRe+h2H0c5
55MNYKAiekcUS632rVoxL5RxflEV9LChttjFYR3wtkLq+DcnpUOJ9ioAfUNM1zSpJEgrVS932Szk
XPkO63ZStutR6JDj/Gl2GNJU3kuKcZjL9RBOc4mBF/6631m5s7X42X9f3t/PPoNl884tR3M/UiWs
uBPuZsNgelkijd2G+0kvn2hnXTvN5GPfLtcJO77KuLldgGRN4fMset32I9aSR5x2wuaZSxDg7KYr
PLd7Azp8UpT+mXvg3/L8pD8Um2sSAhUZa8fvu22NEGGj1aW6HKH9iuYkkfdu8R6NEo9yUEpqc0nn
P7qArXX/btBX9zrXMGmjotipMjw3nqf8POxcoZtXcRkE3uTZSDJzC4FS/N69SRAu9QFt1hIG5vmR
6CxgoEeR07wEk7/uvGoEEVXYEy8VqqjIBNrXmkoAbw9JwE/C74U3w+qn3rP/uxVFqhknh5zYIXCz
hKKgSp0MTIAakvmNaQB3HKgjRp03c6U0X7Lzja4cEDqL0y0o6CNCjppN77zwHsn9omfYHRMsWlvD
ahF8KLamL5C0+Wx04Rf1kOFs0oV0NGbu8ybfG1xdaLOXkdM/DDIEgRo2ohzjjE3a7hdcm1C7oMfH
WNObkQXQUEHDAPMkdYq5n3um3e87e6FsaKdvAjMIecoSMQYwcbvDc62CS2VzvOuq9sKiz6vJNT8J
0ppMLdzfofKYutJxLD7vxz3wMUrh0+c9O5o2sKTRqF13ylzi7kxTGKf50fNRfUGbU4npvghB6JHQ
4KIL2Nv6XV/RQFEDMfNvP2OPyx5qDppY7gXj+AP1OZTMcA42Dvya/so2icIsGhg+IO9KBtxPEIwt
PS93PnC4sG68lKFQCzJxKkl6WhDVoN94FyQ4rjwdwFYovobV/iDXF9a1I2rJ2NdUO8pHuv4afCWh
dDytDcS4prEUYMJeyATIET+VPFtyMc6uk6uE1Ww0mjt+VMYbeXv+wahwZF6ZHO4qdzXQ3makH+JO
R6zOTRevadHPt7x7BZFrNQpfNWf+IX5dNrJavBwdBNKCRF55yXU7CMoyWzIgWlK9pyYNcLJwRjPa
k8eMEjtVxYEkZMc7C+6GYSAlx3nJJCxL72YKW1kNVKhON3C/ICrpVWS2uU6QUecoaki7d2rwB4t0
3V0Ia9PVh4wjepbLkVdWZKRpxY9KPmmZgnu9vTq9efb7COVNnEIZBgDyAg4Q481Cv0j/hnvcORNg
bytn+ELh0jF44h4ifG/IZY6tTUNBdPJai9NJwYMUIG5WwpkQ300v+izbnYxUM4+HnfU1866pIgR8
6meSay50e54mkk280otzg4VfCqfMo6CVcOW7yR6agvHqvymeFMnVQbjbDiGHDKJzFlq625zAmQJI
j2/xSOo+Z2DTRpMjZzxtAKxxJ1py1spetbX8jof+perH+dfilvAPf7OA+nj2WVjh65hatMe08crG
JYcOVDVateTKX37qXqQ+Z4ZpnJ582YTKD82dPabdMp+g5TAjN8oU5cNLvEFf/IeRulVSjO++v5u7
42pRvHQPuOkTok4lu7KY7X3DRuWF19yvyt/3fbA1FTC4tHQMTrSdfROKBojOL48JqPXMq7wkpLY7
ewu+1RabtF/CYP5pIEU21lyu8inG+lJcNYKVmsV49/ej5YZ8qeML5T5tjbqy3+RvpMcVjYd95yTx
CD/yzjZtvV3poZnvYon08PKZpSlSg56zrQo9NiWS+w+zcXdCLELxkB1+HCvt0ujvIY6m8BdcpJTP
tkwFyaOnKHV8nR77D6hRWtU0QHw3GvSZv6bD5HqldAJCr77S1wff7bI2HkY7CmjaGwYknEajb6h5
sivHSWbbr29Uurutlyd1nt6FpdXeThVVHZ+865USjdkb733FU2xEUwjzMzpNmI6pVjBXW+AdSvcc
U+9u4+eh0kNRz7kOi+IN4t5wQQWeZuXJI+jMKxS013s7koe4ON32bU+ElhZOg6/VYkz73eLBE2PV
oWi7pHPky/79mMxE6zHWxw0oLbDB8fVVanfpvk+Rh/jYGAouKgGvHqZA87fUiykamW6w+JRJjozZ
AAwwYNX/AqTPi5VndbZS5RJ5/a2TrUdyK75eWCqqjM6acYcWlcwG/fYcVoZWYzvQQ8woLUYKWhxl
muBpc2ZSxnmceUe2KTslEMHMTEajf0jBIVs1iiNQFdLHAtSDEzcHALszeflPYzm9NYprfkuBpcZ+
M6ktXtolZS0vsAEyFTQWut8Fb4I4LCe6qImzIuV45jVjNq3VyTRIYHJTp3UVD0bR5QZ50CKg9bwF
1kLm08C9ncXPuW1d06l8R1h6ah5L7UHLTsvXzEvyOh9Q3e7+dOSFDDNts1lUInrWT5Wb+QMGfL2Q
YaEKhvRguKIP0JnKO+P25aA9CLBGn0nklA/3xr90MXefAEutTnh9EJ2bCdUYjcd1AD7kukiqrLSA
V116AqA/RlMhmIW6TB5oa3zoTsvyMqXxc93o65bkW8ADGj6zjsS+itEVbTBi/6FxQ5YM7CZXlV/h
xauaargEPlXl44Kntiuz5BqU47WOmCpNMrHh622RH6Gv0JP/rZL4LtiyNHJLNBdqLJwl5Fhn8z/Z
GQITPaqePM2FpX3/U4Ypggb9OCrkXvNJ/b+6PaRqdBDEKZUFv3Va17U1oPoOqr4gPvtvNJ/aRhIK
mkj/mk+mvQ+UUUKUs8iXOCcTahqSROps9D85zWC/Hyh4zIMqfHIFNSVPJpBEZZBRcZVT2LgauEWh
hJN3k8P0yOBCPOX8hjN9t9k7Vdh2KXF36APL4b4dhVEsPVn3P+XXr2Hrf3PA8p710IlR1bRUL6ws
qhGJniI3J4N07Suk2LN9N0NDisyvU1kqerGPBmxzE624jARYVTCAtWR/e4G8ooGaVkmuH1pNn1Na
FXCQK9HfpYTyuWg7+t2A2+hnz5E0/B6aWMkwBCpcLipZVodbjO07l1ZU5ggIMXqpcCbiJs+2gJMW
lS8QDJhCrFozPbb84r0Ve6Cx47obG1F4yUINlulKNal5pxrB1ER8j2DVUvEdnPxEKEISJTVjBNW+
eyCOfewgyEygNEp20LwlR38aRhZbh8IQWJCq3TP2M3OisiJ+0kxUkFB+s5A/XJ9XgJeA1kxgost1
rnGg8zYb+dTM+Vzm/Arbnb6TYE6dlv7Q8CA05PXDCSoYElDnUbuh22ctYkugBoNWM4QxoUUnQ8wN
QLlUgS240LwZzMplDhAiST/oLBgtRyvCHmjXwmJA+fFs57bpr6KI/vi7ABEH2/3ZYYDYU6F9K1Bu
WqCWnpBKPxCSqt5bXB8j+h4ZIIn3mMEPXCWTbGCrR1YVzFOwJRxemlpsSKrOb7H95JI3GRVdFVC9
+pjJsX60Q/3mV/sMfGqsFbUgMbBxSoOXsOIPZM0YZz/mMnJkvgPsCKPp3Ab7cEJIb3IoX3HXW/Jk
cVx8TGpLwUjvMhHNmYVVGecsjFu6dDwh1NxFnRs7ujgf7H95mnYNLkBVBb8YDFG4VWoVKo2AQyqZ
OYN5ZDODhSAigfrETHqGwWXowzMEUgLJQ9UCP0Tr0+sqF6ydouf14WBJuTOqBu9I3XPrnHcqegqG
LzdNqnoKxLWQk9u67dvx2HiG6LCxbxzykYX1Cs4u/RUJlj/evNeT2WG4StkLS/Ycg2NfGj72w2pF
b8/Rwfmg3MmCVFaULydD2HXQV181LbEKzIgFNmm9uaSll7uO2nSOSFl/mEayvBFNi6NyOeb3Bsjh
63UHnptzMAmAJ9VgiJK/ZjYTLVOa6KcTpgBdeBuOiamrf44IaVomMck/3GUpqhmxQfYAZj5/Ofxd
5ciO1Zrs1qO9lMbbTw8RWnORXd+olpd2N2vVpdfdah/P5rlAlFPMM7QPVADdQ+F89Lbb8eJNnhuv
NoNRvK4j9TeHnG91FOe0zUIl8faU8Xki6ae3XxMWB0BJWqiWoFEuEa+ccmhRD7qqBuOVWGwvzhs9
Q0RDbuxhBp4OxDrvsJtN7tD2xBndVlDF4eFSOdIXtPch1L9vqpcZzkE2DyKubK/7DBExQMSob9DO
OAxcLzBx+NQTSjZnC+SeDtoxATYoowg5A2qDGRI0MDDMh8iV5ViwhbVDRIOHpN0IPrbbRXTAN1YN
zYq+CuoCWL/U8P0323+d7bt3YFsht037UFMmhk5UaMGiFrJBNwTszESXvmpp5HpxyJnD+l+DtsgZ
79YhEFJClHvK0ocBtDHFqBeFdL+ibXqT6Ebvu1We1baZabydNnUVx4hHLce+xjwkpos4AHT1Pm8S
YldlLl4LHQgzBbWwrFOZX2I4DaTb83dOyyH+L47bV++BgnG6JliLiafFUMYV6mROVi/wFlcI/nuD
SCgePVs1u9dTtNUF/L3d9AcIpfPMyBb/tfbec5uNwzKtRAe/YqowNBmhCjk6j4ZUmC7E0rfr9vzT
zjjd1+hOfNqNkp85ASL4xZPbOQ1iKBlUZVDZTSLMwnPZY9bmbBY/IST2rKWKBKf2ISSfDzozREP7
WweEKXiX9BGpEAuVloBK5pKfFPNo520xxl1vNSLLgIvp4I3X1AQYNVYbs04zC6ms2HRlbT8Vf21a
fwiJsnr62cs+doOe9fmNBL5EW+tkmC28dA9CQMjR4SMOuWd10htKIJONw6nw3dxZO6ASQ+7TcTuZ
jWEyo8tkc2ibqFJA49CaeZiUUKuvifxHeo3cOd5dT2P3Iklo6RWiCfq9X0DKSQCW5axC07noFj1y
XVUrqCsNJayy6gaCZYArCMYnmkCJg7DbPSVdhTwN19kkDNWJL/zEJQDiH11UO+n7ChNMT3akfmNE
8JLhxeBmVFff87JmdDJaz6ATkd76pCCYgxglpTboJkDEuuB7ejR1frPMbfhwFMCyjnImoDftjx80
rfLu3Y6mEHC72X7EEMN1fBH/nJARy2SpOcZukCRVENG6hGuJHtEzPjL/sx2g6T1m/CAEzRnyOxKk
lJCWZ4f2bwGtbD6pWFavwbjdHJ64v/Lxwxe4bmL6LnVAfAD2eRZwIO7L2+20yqPLRaNO2GSFKdAr
QeEq8VrAqjVSRrIRYWCUZtEblJPOfX9bQvlJj4LCRRpj1RtR/kCIarTrFn7uett3GxIyRMrljsLg
NEE57mYNoB4WaC6exMnLWuxnmMLF4hUHClBbf7WjSGyW21Z5arKtRpA1jufSVIxBlYTx2bp7A7R8
Z5+MD0BDsJWDrHRulW23EdGuPSD8Jivg95lLrxKdFwZdQ/vOHc7pDCQhHZ9a/Qmoe/6iqtVBGY5c
6Rz5iK56vHZTgrRi00v4cHQ7t8WPYqN3n7LY55xIjjWbuxY2JEDei1cRqypWwaeMpXycWFuEVIsj
tlaAaOy1Do42z0xJZmYTYnAgjNsuwfjN1w4JfZs7G2XlzIO00RczGVyBqDjhax69DsMsRbcs9dRh
WPcF8DZt99le5Tk/n2ePPlF+ZERqmgrCfww0ZNr61GeHedy9Z86Athq0600SM4bQvfPDo/MnCTyz
wHlrhFRNzFkQG5avo80/MgDK4IZkYR6pqLNRnKvID1SmBSdrxpV3DR8J7aIJgTisF187gEhBJqF5
4YmF/krIQe/mfOijVWTJ0tFN1Qqrz7BFgzEIuTcYaN/mdkFKDS+TRPBcDeFDlgUTH4uE1HQLu/Ii
7ktphF8wxPjsEEHBnoxnDtZNiMjc8HUxi9wYpIQV4ju5sv38jszRiYandwCoizVXcYjkkl6FH/nh
cSh3hpAHk5lL77of2vsOBzrF6+h/CJ3M2W3VuU1q+nJjEA4Hv9aKIW/06z49oSNuQa1uVseTd4/p
YUXikB2tYTM9P3L2BlFV3hdC6UuTw7RxD8cOc8zJsrpxAmmvRanPDsyvQfra6DcVigsAUSnm/s6j
6RTo/YBKDZEVC9w7WiEGYt03+YCXkyzxtyH3xN83FMxmzSmxhmLsB3qS/kfY85mfXj/83B8UtYj3
reDTddY1u5H81AqGWFDtE2sKssdF6UKoTgA1z9N4XoCvithvvKkrkILTOoJp/fvHmeiXh9BjfrUl
uS4CtsG5XHNhcUg3Lu7qohPaDtZkBfIwdw1slWvUxZH0HU+T2jXS3chcXr3GtgRI5iRkFLiiBTxW
oOEZz758iMEmskAegLsQasM3k9fTZMfRdNIUtEfFBsm5oprJBOa3yXqmY/EPyl7Rzy5USH5lSL1Q
Z3WQI6DOGDgkP7qzR0bskdJZ+6KjhqjKeEEW//kUe4E4NlCgJjo/UbogU66xG2kCkaOyD+luYWFE
Vt1YPbnG4zNb3K0WaVwXKhkNq76J9NS/tXm1QepNkMpnsY3QxpUcdmIE8QRq6+mXNhmr3XEefbV5
tfXbi71p47lxUNYPVu25/aMZZj9EM0w/i4trTZC7Qv6KtP5Ep7aVPAhQJRQb13q19C0vsGfQw6t2
qpRDpfz6ylcjtFIdm2qpVI1+wgHlb/v+i0SJPFCqAF6pymZrsFfVdlCmvEqIH/zZMp2yqdgNp+N1
StYfFft3dpZ+eBNAeJqelJtwhfTQscXsOYOjPJ6XH8jAKZhv2h126P2jBMAFj73DFan/npxdwa6c
Hxxqjwl7p9HyXTU2yBxgy+uzJ6nvBE1iaZw5DDqeFlhC5U3WT02fnACV1cXlZK5V8AYV8eiaTbto
YgMI7E693OhvG3Papb7ehP7E+fzeocGkZ7MC64tpfCZ8pN7r/E2/Y9YLZsqp+QZaEaGpTNIUD5ow
ZiWGNkm4J8UWHbIWHFi72QEHp9KkuuwAY+xzm/zzzrd2RjOl3mBtFtGbIx0qwHjHEp4QQYrvO6m1
2RJhSzzOdOwf78znQmbh9/FdXC/NVGcvL26kY3RbGMtQUy6ogkd8/BCR6KjGxPqiU2rxIdanWtjo
vcV/784lV2ZMPiANw1gTgPaKZ2WuS2LetxOnRdmaOhgxJuMzUt5jCs9KhgRr3rbp91udC8fkZfYT
GyaCJMx5HQz9pPHTgyJDAPpY/26AMSPIXgwRpzukbG2u/O1EaeVD0fHvRQ1jF8VXB9aaOODzymBS
Xs+pIjdZWSpuZ1mkOVeMFGM+OSje2K/sFS9gTrGfgcjvSgpCW/fWXKEXK18aBqjWhMJJwP+fs0EV
XA1r3wYabl4ZFpZWOWaFWieC9hEYK6RtKLoNXLXQPd8bJ1XT6LSOlXZV2Wy8LOdDVoYairTVABWf
EYMwhO+PEGG65E9PSjzGoyS6nFCd6MxyDKlVBnnZuBWzyTldaG/PzLFcdEpjn3o4f+VG1Vq5oFpg
mMDh/1AU0dEOnpwrubFcrlb5nzKG+/MgGdBebZ7tUEIuMIakqPe8/gQLg5UviZs8U7XcTTo6uQpu
OgekWhWEEEuKcAy8Z7RJT/eepeRKzZsBSRqzxMEqaf1Md+fZb/1ENzSn3OPh31pa8Ero3CSsh9TT
Qn3VzM+hzxaPP1wbw0C0dGUN8U0ijI0LGQ4WdEXies3wD7KkKFtfx4rIt9ES3+5rzSzVmoVbzFar
h8Z21xb1/krIZto0qufiBvTEnP/POF2PqEM5BUFuy0n7FNWdQtoRW/V02v4y2bCxlkEZEbJV2MeT
m/9Mz5KTrPFNIThcnB2kA9Q3t2z6qjRp10x3vIBGPLTM1sGBmq5jJigBl6C7Hvu9DIv6da+iCOU1
PTJnLRVbG+WWIIfJrWeR8FVbmWWCjMAzGXSXvr1OnQ7XNc1ObNKjOQIL1DGbbU1Alj+h9laCGHSe
R8GPia70qUq5QCpkdyiXf2TF1zCG/aXg+yuzrJooEPS3XzgfD/3ECLdoLIvrvYPVvDbcdI58ioZo
S3nh6EuhgGtxXV0BGWC5h4htzIAJA7RJSqacLtIxS6aObnlTNG79qP3PlK916hOmn9DQWxC/NWy0
W+9qMRK0MyX3l9W2iKh/BNGv0WvHy4vlNa9tHAqyz33Yrx/rHN+qN7Kw3Ks6CEQsW5D8Gr93NZuQ
1MNLbbxdCfs1EJJWvIkS8XdP40LudIYNYLQR3RDKEvOzxf6PMD2Z+aNQLXUf3Uyd5dELLYJb7Cy3
UEqzl2KgqDA1IKDDepxVyn+saWXr5oU8I4G8Yg1Ms/F86cIm8qNHVoDmBVQYnq1IzcYf88fuTprL
aUDN4DwZoUP6lzLYPdAq2yVycOEIw2uEjJSNy1G7VOgpgyvHVLFvkeMvp03PhVFmYT832ozoJOv2
IQYkSh5Qu3Zir8+B1nvQIxEqraDM/63IgtxIFjRgbRQqh8JI5mI7W9X74vgXlhoaL1PFJOL3Suup
O0HEAfLns7Ki1J2y6EKECZVkzzpcMHuTrMmrAdBQk1L8g4clIDgT7yybf2sWoJ5hJ31Aoofw5SPD
ogm3U3BMzZ1IPdGaQL99Mf/hbJJYBRJSERIEAXPWGK1EVZzzGgURKOObdDRBKyLygHmZhaUtCbG9
d6/UK9LWObpe/s8BnnUrXhApvkb79/1go8fxO9/RE0PTnv3coTuNgf3QklGsEzcXr74TzBNEuNra
L94+NLrPaOFr7vl+zLCXHEj8NKxb4UZJY4A0LjEnqESpajM66puL17QspWeVgfUifRMWmf2NKL7k
52IMLjrSyXeoZ9HR/aKTinVQIs0fjZOwb1KN3fDZY21ixbI8tdGUluf39fycnAq/YawyR4J7nTt/
UHQyAa9SmhWK9q+Z6YJLfBSpRsXIexaIqFZoW7Qs6ZNIKva3oVExWBay8k3QrwANsXCRaG9g+VZe
tSbJ+ndbUpMISqn2aI+h25xsAzlD8J/3M6h4Xpbf6UUxk00IRqkkSEk0gSNDIJr+72RR8kWaTED8
1cWlJ1H/ov9CTfZK1D15x+dkFwUBHvaZIfUSBJsHm6TDFlFSCuY8yoRIS4bgmxJ+a1uvydnK2reJ
5XdWkPLgzcoRKIZZRhVDi3c5kxNykjm8mF8fiBkoyX2Lnm1hChpMlWbuBdgAGZ9efqMKaTXOM7FY
XFr1OV9VEWVEqtoqfZudz2XVptPREmA9Uo4qf22U36kfKbwOhduJ7v2ophda2q6yVwAwUQhVLLK8
k0i2vE1/lAZei1HS9z9UMmQRH5aiPVttzXFDqI+Sl8lNRBvi5yzemz5cQew9YcGRMun7avvnCo7/
jnbzgyLOvmOkFgI3Dq1XRFiS1SjWq54M+9xasOKcm8u80VHHsdRqQD2mOUUGNKDNwo/NgHJaETS/
v+fr5ZqaCCXs1Neyq8k/hs7j6yhgIOA4KIA1BoPaEqyWhqLmD3vxl+uhDtz/UH8V0IZ+mrtCf5Fq
ojd3X9LngU8unOwIsvvLy9LVe5YyP7bX7yChF07emh2YgFfesM1K0IiYjeaqQoIjvdV7ZI6pgG5c
bczCsEkDcn/n/c0O47QUGyRAwJFoa/so9/kDDurqEZVn93zqzP77qKyE6lUQTkLgTLQO2BUDE6wu
6oALCvbykTaqO0ZMYdjgYnqWCXITYf/h9PDqNkx3Bt+HfX9FokJaYCuBPR0EPvr0j4Dkw23+9s0f
SUIlEhJx2lUy+Pv1oKKf9lp+W5wHBiZMj6/D1bup2PZ6qQD/iVssaDNPo48QguiZ/nxMONOoHhkN
mCs95q/xvd+djSzhkUl+k/9Q1jX6riPJWvX/gieZjJ8K4JB83EdpctXXiLcfJdQ1wQJZirTKN08v
lccDRKnqvyci+gJFcGiazbYqU4OW20OrzywCx5wb73hD5dENtpfZcbBJQi+3nj0JyW54fR8YO7qI
fSJwJ5TD6nGEfD3xF2MTPyctck4kR0sO1LCpcW7BfvXOxS/HRDVkXtn4Thu9STtFDY0M9oPK/m6j
2hbGZ2zUsHVwc6oHXvy9/RceAexZPcKVMgvvS8cF5DxdC684m9EMGuBWXkGbS6IHN0ttNSTbIit7
MmeWgXNJkOwqGBL+OY1vyoaJSdBwcTyYIGadrFxc/zmUwXEV4A0f10jtPS9VTpvK1eaUk2wBI4bq
WYaHAF/K9010VSzHMdJ/ZOSfEYWQRDxnLt0RLB2xGoKDzhT9HQj+fzhsN5O4GRTq/6CwfjyAVW2G
1Qb7BMhltlHLeNMogFlpGUgiJO+sUXo81itRR4RZHHax7b5w+dS15KpjowAXbMeac6PDjbEET5rg
WShiF2/KalfrFF0/EycLRumU3Mx43c9o+TLo4X+08kXhAG9xxlbufnwiIiv6CSw6PHpaEsU0IXZW
0tps15Hk3Di+MuZN0KqoY/ncjtcMfDTrTAlr5BP/tJeFsjRJSx57650/2miAWLp2oV31FiXhi/wW
k8qIK0PuPXSQ94VC4suN2/OHnxxASmk34lslybE9fBlf+Nzzrn2zEzkga9+NzrTpvnhVSIydJWDC
Hkqj/i6trVHr8uyHktTHWT/MYPms1arHYsvrycclf46VyssLDppwVirY0eB3k2y5JD/MrqIHhOmu
tsoXNbkwVbt51eQU4PS1Yo419GBjjWaiYD6/3Nqv2x8TfqvbN2FuSsUkKWaRck2oFMkJGMyvyGoE
Vo6gE7WwrtQcdQKuDRqoImZBnY0vkf2+lRUUp+VAVnwRgrirBQJnFZGe+hLgNR1NkNzIkADb7yOl
OTH5DXyLVKvK4WjgsmcEMrGdSroZ1DzRLb9RVMcIXqEtiudlKzxl9xGAyZfag5bj3555qhqXy0G3
UfHo3SCRU+GGBLfzh4DPsLzZPzzElmEJhTEY7pmIpbOgXe5JRoroTjOrJqc6YzQdmo4+iT32Sb40
BTrJTMKcvuxnDws25rl/zCI92LAG1vBXAvdegdhmFk65HoJTUD0WO0FoMlHiGyKFNHCX+qF4IPBE
IhWeNs2gUhww5vgVJNOh9gely8fHBkoN9WyvYl/fG5PgDN2rsJ2u8zDOWuRtOTR04We6HCDWfcz3
SWxxQ8nuWa3i74IlEkL2Gq7B+sOrAhruRi4n219cPosM3xJHG+2LWu54kHLtp31MagQGDUU36blC
0n++9m23su++vqEZmcGNUV557InHQAhmo/T7mRvAjzhI+eiHtdRQMoInIsOjFKtz3kfnmYMdkFka
WKi3y4TTVeks+vwEW+jGhf/vgJZernND0/tqmSdKZANB5BwIzkfKo2fZVswlUuoR3S4ytDdvaHni
EfeYsMXhLKcaxev0CwWrzItLcMmUlIO9IxxYRorWvmO1ctQFSIyW9rIwF6AzdEij0friMxfjmbPH
ybNide7bAKcqMGGMfpeEHIBhnm1QnKPKAR9h2QOmgqSZ54TPx2ceLJ5GljOQPBF6dJnX+RadQGpM
DYKSwgrwg0REgffBILHPkxxXr9T2hue0ObFtHSpAUvLX6htkGfWEoNFiFs97jxxpkrv5uJlF0hZD
4GHF7zO+JiqROx2110y2MotFG8vBp9lswm152hieUq/rrrHrCdneuwQrMDDIovJkbrenkV/NKdMI
ge82zCeywctlohqR1+V005j8ubsprJsRinWGrZvcWkJ43tKtfOjgTyvsw9qeLafZTtZcu5ZpCqCV
WEvnXOOCAt+CNdJ0W4kG5NL7wuRc2t8s+ZKTIdZKaUQEz/MVlRmgYRJuYLbtJmhN82NJo0px1+NQ
2gOD4l/ULMxhwqTOFvbq4HIuKJsvKM5B+T970GRG/SxMr9VUZORvxhw7TGFtNWGk2GuMqTixZozh
tGkvxZUVZN3a9RHDVdZ678z3JUsPvrNbkbvDzRVIlHKVi/+8ZP1c7eLyP/W9CQ5W9BS00PO5QFwD
wMiEl/Mpdy8xu8bvx/51rsHQfXgIRy//Xee85ymF6IFO6DYp2PR6ny48vA/Ei8h0I6IfZS3hqY2y
Lbfh94WMCzbwgbDCxHyILstzHKDer8g55UVE1GUCJneGlIsKhBqeRM7aTz9KBOMLq82Ki2l6UTfD
O50L+FCsRuW5yKSgGtlY/eUTtDxzKD/x3D1/A6Ch3BCme3Ci/Nzphe/trGILojWOQ+6w7AOpAxvB
mS7FfPgxj9skPkHcauP8evDhId4DeeFRkkLuFAMezZ9TQDbxIMoEpYBZPVJkjhdhrcYBr/wl/CsP
JWegaqrvy/DuYhyk50ks5l+VRTUUfjVfieoII5IrmYVdibZlHyt2Jmas5EixJ8rx2hrN1XjovKoR
0M7tUyXrWrkyxt5Lc5D7ESPda3LSsjtQA5k6StDD0uyT3G2UPT+MjjOMDCkZ8NNUdyMjuWbykFlz
oY29VsFXNJIhxMJXNwPVhCklJaSX0wDqVisMF66olDHbigzSC7tGZKV5DHoWeu/JIsEBfolouiCf
4oTdfoX1oyspMS8nuRe2ABs8otUD8mV/d3EdPSg9VPSOZ9KsT/xMOEgb67RlSdl/QMVvvensfB5Q
6haevxyyUDgNVR8WdFLlALbCvoLidIOVTI+rmqUXeYhfoIOaoe5sGMVyBeN6bhzw9PBoWiqGAjII
UMnXeT4TKdVBRoR2j2jRBjdfq8bLvhYN5Al44lM8FK8XcTcCOf/oMdW6+G8HoKbHl8LobwDTXMWZ
++XrRL3TkHRQWPcIKo1wsIyjbOG2d8T/QV0VIY74T5qfIufIEyn1gtjoLHfpU5o2dg7nnxDjaVD8
v3M6xyyK93BF9e4h6xrQTgysgSu6LKM/wq4MRH/SVO7Jhg0uiqDrWXxMV1QEOkrBjese6Ot8Vi7U
oCz8klsDKnhYLnDaFhIwsp/APRxs8xqyGt2bd5E1bwhJ1W0hu481K88edXsOk7QHh4E4nY8GAsR2
6KFhmKSgpsqLRIyRYiZtQOoRPomcIRm1gKRwl7FZ/ZY3mWr/M60ZRtbSHsmBdq5l9gBRVL9TvWsT
5XJgpKhk8ojBcDlKIG7iZ9SxPAlLAWiZmgCB5DTXutC/eaebXlpwhnIzupJIsIhYq35HJefneAg9
uO6pcUvTsgpa5D81QA5sXR+ydAPKknV+kxgfhSYHcU/c1jjqW3FnjC4ZhgSuIgI4JnAX5oN6KY3J
PwvWghlWu5lUQcaDVu9oy31krfta+naf8syQzU0kkKRBh3FysbzCcyIGluzDuni8tbNVQNH+YK7D
ISdfrtgpCts7RhpX1UhjwSmVr3zAHULMMCRy42cQRZxBnIh5pbMsxv3u58LCXQh3Me55xLgVtdZB
s8E+yj2aPLQq3eMWHl55xesEf8FJd63LWJeBkXxnwLVxleTprz21sYrRiiZx6LLJQcNnKNmdgj1w
CE95tWSJmsa03TESYrGDZDH2voM+UbcIqxDd/4PalIQInWSa8PPmpQ3hV37euZ3aolAI7ysM76RA
N6OtldTefI4QUtr5xP4NX9wYMVYcp2AEKVSbYVDAdQ4U26kF2ueDKS8TlPZovKnp0//YBb6938V7
OdO+g4uUVwbKqGl679BsGl54IEEpKx6PCIQrH2sWyCG23XCSf+Bbnxp7+CmsL+0dKT4DZ0mv/nql
0Tqax2Jt4rF+fzwwoTd3V4PgUh5EDwoMK4/74Fh+hWcKHODt/TjXjBY5fxnhrhxmxMm0LkCX/F6O
yHv4qoMCasCG8COPRCzGHnb/fnxZpVzdVnzoY32FVUUDGMAl5+tlMg7JQF5jz1WmRtyBfZLA5Naa
B0woC2gzipkvN9GVH1IWNheI99cyl1QK2Rf83TJXFHtaFARLIwPSJnWKmRTVhBfw6E4xKH45LJ4U
6d+bLysPH+h98835QRhUAqZqhM6fnRB7LFaqOQE6lqyenOShX4lYsj0+0ByCFNyt/ynROkbEvdKy
Zg1GMOzmr4VeIGhkBiC/e4XvIfNrEvNCeGjQzerFlLxN4YA/Cz//+1GdO+iYS4jhYY6M/aGWpH1A
B/Txn34mk6fsm8gXX4WBt+xoOmWgZSLgK6pdw7lMqN5w934nYJyEM4hV44yU+QR10KGEnktVp5Ua
8v4VPSVXXPtKvt+jOWx08sRgJga7U9YxFwkyXT6gB8vbxXczmDZWZ4iKJZYtuPdiWTnDrkDfU85T
b3wEI8pGKyC5xVkYxEnYbjHCTPN7QDTfXy4uQkIHpCF6CpIg3nA5WRQXfpJkz+yWiVpIwFS2Ia1C
j1k4cvTuINqRy93CHM8+ZAnvk3TC8oIZXZuYQxjhrz6KcufVRfxr6xl7FYzKpZ1CIwYo0bWJi+qt
uMHluqP3uhGrYEWy2+Wta2SXW4YKfXddsvLAnSFzJtwuCYgUzmhUXlNmQA/Hw/2cI0IoG6sFLAL3
guGCIVx6ZJKLHMtvdDs3x6X6gQUXIXmRhJDoK5Sj/l19kUeEDTN2MATc3cGJlDOW6fmiooZezBqa
y0fRiMGr3VrHD+wOrTC8TkFwGE2+PFflh7y3Q1hE0g4EoGVd/7N9h2XfYgz5VA0RSd8XZo5XOM6Q
JTtHsL6XRo5k+5Dv28q70TZRTfg7g6tB6yPCJ4TtmZl30DjyDjKjwjYrah+X0iVBvBsvM3Z1eh0R
PgvVWXrSQ8A7hlLxwBfTWwuiNZ4tBSmS/cwOqNw28V9h7uTSQO6EtCkN+IIngNrX1m40/AqKx12n
kwjRW8UqmTW/GTaGAvs+Uj8MAMeWdJIckD/R/IFfkcDlsvxh5asUL/FpddQfUE0YYhRxkOHBYlog
rOmw7nJnd6V+GbCKx51au5oWDXLVNo2i6PiySteRyGqZADFn1mp/2NukFMfCzMhBmV4TvL3gjhXv
b/uql0RV1X7gHPn+OBOvVu7P5LpRn1kNnzwXsNuH90uqfg+0rkM726+9sP0Q6wlbXsjk/1f0f/mH
OK5DPSU/T58nsuU/XKiSROohxdFA5/Od5pgvAAZ3XNw6DacehbamSO+qljaYoAXIPeuOVrG7l1QT
Di1+aeCHVRP48q/7gha+5Pcy7aVBMHuZS1miSIwMf5mxT0prhB6zcR+qw0OHlZIeCNXTidLtncdw
74YkG5fKng1Lkp8Yj3zS2zcwMWdN7Mo3ic4GxfCLQqOncph3vw5PSDTA1WTTl6lXnWp6Nc5tpcuH
Ws9LZlJ+eIdhJ89tlyEgyVvO82nyqtsBRmfoM/CCaX4yLKWjpG8iXdiJh0o4HoS9MFaEVdToPtbf
8lmsDaMnizBt9PriDi4rbD3XR8qhowhYzOiSvcmR3hwEciZbuJ3GFtz+pJsHz/Vjs13ausyYTPCc
DNB3J+eOL4CZQcIwfo39R5uyI3vMBi47f5W3zhVGWwChqmWCo0dn/oSAmYF4JvLgO8sLijkfN1YV
w35+UbRj+UR+O0K7+vvVb9NmEIcUe3Of3i9RQcm0oOehh0+KwpZhy6JYJC9obZBZjQbyDGA7M6pk
RgJFjP/2/AYpN3rHcPZTpebvddQkWKOD+6Ssj6DhjgeA3s59AAGojWhZE2ObPo0Id+zrXGGryUSx
X4hSkJhmQz1RN13BqXSxxGxzcKihFOJFNmSLrfsj4shXKyusdZfe7I8wviJuEPmGHvlNYf0Aa+zh
mAxigL9gSqbCm5NAHbpbotbW5ngnV9uzBB5R/jyrKguOs9b8AzN3cn7qDJVmPV7TW4lhse1F+dHz
McGod6H6xQaojpDM6Kb7wwZgTIfrlTa2T0ZaurD6kXzU4oazjQV3lMlGaCTAvzia3WLQ3jdF4d4W
aPzSJfN40wY54G/FhZaEzumv50KW9bTsHGADdCvzJkkUnVug6ooCE2tGE3wmg+QFsrEu9Pehjrpm
HWCGVuOWTEhTlTG5OGe9+3TOTNFyDwKiR09MReRD8ehXbhPd/K/20NFksTIPwBw1Sa/BmCdxj0vd
GMHSg2cCFNZfy+C0qLCRqvWCrNZNqDHLL5Xed5WyyAJYpWfqH5izzrCfVM2WYpi/o6Asijo7dxdv
0nWSg3HYKjT3DYWK5ugIib20B2Ji3EU8OnjFKGuWP+YRuJBG/8/rtasE16SoSwPJTffex+CcBD+v
1WK/UTnucHgzkq/4nwJzJuP3YAp1jpT8eT0wa9HL9slVFAXwF2VxfsYQ2rUGMXoDWAibcAuDVAMi
2coSBlR3dFA+aw0pW5XnYc0BFwx/yCz5GDXLpY33kkQgYrLIhVGN0m5QsrIDYn9+YGRZ7XtOVYZt
priRjk2AVOf9ti6/D6H83JWn96gOTWYhWEpimHVErUX0+9uUonV4EiLAsWrP1ivOK2qUDegAf2LU
n6hRxXAsmDqrE2NgEYdUL7Q2I0eZ1YZhFfq7/mMXdhPtVffyHmg8Tn4Dd2PGJDg1oUCsZ5sSprdB
GwSpinfny/dV+m1sbVkxdtLXOSp/f7xlqx9WRiJ4yGXwGonTytf7y4lL4pRPk+GvP2s6ttmtrEer
F+8kLexM6Ib/3MR1a2o4rnjD6YVwAJ8RgEBTI1CF4UTmzTB3bKdhhCiwRQltc9lz3DD3MYK3hv4O
leshAfd4ZWlOH6zsQ0YqPp5MA4xvC8bLZR/na8r0NYEyyJG6odYAOa+3j8ZC50WZh4cuUbYdqqzy
PF+ppzyFSfrMnawL8ZS+3IEZb56ylrIRCbO+Rc8BjKpBi9dBGHPd94xGym1wpmI/Dr6gm3fbAQ6o
VwnjNVU+piktF6iqfK2DkABxzbAs4OJodPZs4xWDmeWJRKzOt8g1EdZAdL1Vin/Cbw58lsdKQoLV
VEOI9cnwYR9ec3ExxBqlDBqWEFuwF5b1HowXBoBZkrIAaedpnChCae3+ib4ETzTJQ1LrY1S3SeyX
ZY70Yq+tZMMRoF3Lh1kAVwBA3CJFCSpxGAyg/GgT3WJnPd2g+KqA36+Zrk60GckJfoavo+0EqWk9
lepyF/jn+b/q3HeXx43P6yFOQOOqUxhtkUutdEX6ISN4iGqm1O6JyiEdAkiVG2i8XUUSexJY7Q/l
EKMF+zGdYFeIOsEC/mSfufdcUDuVhAXBehsNStu3749QWkVXzxvdvQ0tQnfj+n+DO1KmKaXMBSUa
Buu7c6ctAj0GjyWn4N9bFgZAaqfzqKG5onuTIaCVbkGrqNgA7rSW00RNotsFDKl2nOBcbg5yJYma
YX2H3Tnt6Xc99oHEgjrxGbKUBl3iq3SWoX0HrqhwyUCC6OXp2ts4anu8JbAMIVJ9kvP0uiZAS38I
IA4osQpNJKjH+Bfd/NXP+0OaSKNRIlFaIeWvngPaUQR5DDHK409SAcfbWxeb0DzNJPsC/9hhJm/j
KwuS8VqxU0bc/xZvaVOcXT1XnnkTGpsnV80CKbzKblt4x5kHFm2FdhmFVLhbtjFvi0pLDKkcsRxY
a0CGcXTgOkXW+5bn2YG5MWe4nw98bSfo4EXfnoMOYDdafimnQ74lW74B6EvH/gphDeJBLvkkgZjr
Ah0aHsYBll842dYsx7ombIjSA6nbns55hitOAYRMeuAjHJRJ9pOKhRaoo11R7eE9q9OKYWLTeHPb
2JfXhO2RHfhtwHyeCIUYt2WFJyeQwab6HaO84CutSwu3+UfZWq6qSf+v7P7IRHoyminvTYcCKVMv
VjAQcnismoY4x1cCvQ1JWdsehdLAgKYJrAumB1QFbSNrk7CZXCEr/+5DYIRGWDt3lUVpmAZj+pTG
+j8XhV8Ab7awhZNgqovvvFW35FX+G55mvGsu2ZdMf/ZnFr24VDQn1WDVPgMglwlgF5wSJniLbmuE
zySK7i10YNUBO0kmNzMCkT+vn8mfKWR4NI+ONLqJyuhtNbVVy5McpBhOP7ekbDTmEDZleNfr3Jae
nPYIZnxV0q+y5UTk+bTbOxf9Z0TglTYspWitibKkjqcMwaOWUNejWyW+NylIQzD/kRsxqbJuBIiu
eab75rA5HjlWMVwOoTZMcRCkpDWwlz5PJ1dre8vASP5aS8jRFdjiLFj3JIeQVYccpzO0/rgIPsas
7B0mRrUKCk+fZ65U2GTvqjROqIwl27LwMlrmDHYiMOi+SfNGVU48b65LEIrRh/+dnJvXLgse4zy9
M/921Xw1sZgV5qJ43q93wqXSefSxnhjOxPiAIhiwrRp7yNJjHHNhN73J1jQCoOWPkFiN5C9G6W1w
S4FPl8F7oIir+I+koV4qAVrBKdcw6Tj2zwZTrzskOJog9Sw/EcHYRLFAFHT1PllYfj/XMxfIsZAP
YEEEgvyGk7Y3DgTmbjg2JCASb/OLSRpLTNoy8Eysg5oOSzS9U10cMptNw1TSfSsCqODNLkz8//Ro
l32rV0dRpE4ksyuWWuoWazlC8QFtH3lWUZTnNnNBG+eYT1zICZ3NfJu0Xd+kEulGhOSwEtzRhM6S
DTAn2/hGbvRIUKeJjNKntwWmWiDWNC2zrjkimf00DD6OpNh1mTxhY4Hp4KZd40eYwLikzTIbyiOT
GL1pkO+LXZSxjYzEMCnZABZzuUWFM6BeR0IYAkFbwPr6QfUzw6YNp/4Nyw5v50b6Ptd+PPkaPc9V
C0cnZ4mLMb87oCtzH+wjnbZaPJf/wY8zpDmfQeONso6C8KwfD6ZkM9fH1ZesCn5VvGrKdSso+ubp
sPNR/pzxO5JBz+OmCGBPynTautS91KG4FTySLA+KZNBfvcGbI7KUevyECtLHlW33k0bEGSZZ6dud
se9cUzdgNcRSoGNmr55/mxAV9hHq27O86M2dst40MLpMr7OlFLugf2+rEYbBJPsiH7DwjxVa0rje
hTYlvbdT2Qgz5bQD10JCW/WoS6vNVA8RNu0EPStljDU4aSzdAEZJE+yZZuPD+WWdpr/MzoDGymH/
9pfyHPapH5loV92jYLBAQpnRpRujWyyB/ULs3+qT/NuVtOJeT5kkNnKm5W/AnDQvabU4R8PSD4Pw
ZqVz/5nAEivC2KoT0QaVNK3+lMTPNiU468cJrb0jwcgNppPmc83a1axGKN/lLtihaxHcuOl+Py8h
TIcvDZ+RGsd67rQeI/0CrqneHcW3azD7hB2JpIXiQCO+p1eahdkTBTCar1ikxgbkuRQJNNR2qf86
4RKKXdqaFEfqw7o/U0qDCj7aFbLmxWEXlh2Ywqcr/SF671rPyf3le6Hfmz/0uboNCwQ0B9zxn98D
0eSVR6MjZ/ynoJ6t4LujeI7SdioGy28Dcwr2aZtaT2/BQSDkDW6eXbL6zHIHYk7o9CFx5rI8mclU
DZG4Md5+SGGIN3EY7xIU6ShmlwIVf2oVrTYWDbRS9Pc0tIQLoqGhNNeh5fa78ZNT6TnyePbQYZ2i
u7nq7aX0PA1HOp5wqr0ikmmfAkev4H5mhJgIJu+9V/zDOc/p/Ry4YBaOG4BLEu3mOH0GAZrBx38l
4DzW2crSyMXLWhR8ocpkFnhJBft4rty0I/IPGokaS9aHUmk8Ks4RikVbXVnLLrs/pzbWwSuflC9I
0WeQdzdiZRrQJ+Y56gQVqQ0psZnfLSxsYjqgCZWVKOhMmtIQL9UMjmCFbBp7pnimwfTHOBkINp0n
M5DOmZ3bTd34K5gXVBzYlZqz77wzpH3tM55pLEWmowW2NVz1Sqg0TNOpE46lJxIlSRVLaPHWs9Ki
GNbGG7FtWi9D/m3rcTovGhGZM6pBkVwPli1szoC55ZTSKMIgo0S2p7UN536Eunrg7kL9y+Ox7mVV
LNjtVkSTYLN8fVL5eCvtpAtMsdkv7F652jgeYIRjRDbbV0Nbm6UJwGTfAa1hJKjFR0K+jiHy3VAw
P5um8UTm4kHBAhNhpZkSr610Gk7rMxZj+jcXVdnSugCo56MfmwSk2/jhuz653VPtyiXJosc1ltBn
HuCdJaj2Mwc22QWqJPYLLNRnimsmv5BESmsZW/tVLGdmnT+C/fSujXOIvh/fapwUzWCXhaOmE1Vx
C1p+u0E2eH3Q6X1N0a8TDfjyzun7McWDukcGzZOu4FB16Ca+2dZZ0gt8VxYFw0cj/sysrkh4a7di
VcOIShBq0nNvYaVzlputSoCisaGno8WhKqJ8Xa2kWGSt8pX1HGfCLAluPO2iHDD+0RFdKXhne9Rm
hpo48ouGHykV1g2MjeWd1JtyeENg415aDt5jjTMXwxNCAFbLp9iwgvVDKehJHNeWV6C0W431OxoP
bYBinbzRj6KZnA8AGSgb5omYlD7e3t5jhTVIgVUdNVtWWvUCL5FR/VIbCGH5Uir/9uZcvegXlV+y
BPcZ8XzNXHa0mGgBDXkNorY8VEzj6XVPt8sdJ4YmfsObnKbMYJycXICqjzcYS2g14puzuoMTXZg+
wsI9unQGUNZSysyU2+GuG/UHVdgJ79zBlG0s9KAGGUa9EUxDIBSnUGFA0OCFPeY1Hig67GhKzSNV
fJyVDgA4S6vzOZu/GJSPkAa9JvaJswaStBAQDNWyWDYb5iprMA0CFirRq6YghQYbylbrvp3LKnXZ
Vh2jNYxklPrOKHMvNx7M7Ydv7lvMce75dY8tlw7RbybjEQEI0IsNB0RwsbQ1s8L7oJT1eTP0DkAz
MDwaPP+DGJzQurwWgcKf7/3wrEoRn1TW8g+tJJv9fqjI3cRFGPUicT04fgg4ax/gwnlv9fCnsHL5
cgBu/3lMU5Kvtwe9l2LQRDQW1mqbDF2KFQbuZ4PHLQZZ8AlyeiV1PDqQqcE16j02esyNrhsLw+lH
0cJUXX3+2X9WAjfNkJ/nzTar5VpZo8QZ+/DL45MH8ZuI8B+5F5rI1t+T/M9QBFfjgDCdvJaW71Qb
7N1MVofij2vd2NQjU2YT8EIVtW92Prv6f57zjEcDrpsBP+/t2WMViQunEafhbjIHHcA3wLn1z74O
8FPoPztDgcjpMSANyogz1BMAPCSbSXzAM+1gvCLzxlOV49AImMy+DadhjP5s5hNUyfmZvRC0WMGq
KmM540M2THP1oWqvwLR+EYVDphXO29zzt62U0ujzudo00tY1T+fGvovbRPagD4EGL3weA1Vc1TUg
/dWagYOiD7aFd0DbnV13VQZOUXCHO4ZrmRozmsN6eO3veHit566sJQs26VpBZTGxHiLFCVl14TW/
B9WeD5u5XTFTQ7U2bFlb69I+79GfZJbSkiJG/5tzJbUhdfaMVrUZiRqEIlgQl+gpjOWDGVREVRb1
YDhiQXqaGRMS3ti7jPT3F7WpgMdvo/UUF3gB4Yprx1p0sKsOugCWAthl5m6HZ2EOm35rZnoOT+95
+18tYIdxC2FK5Twdf4o2jN9j5fynXVOMXuPAfilDX42Pmkag44Wtlht4w+9kwnRGIDfEQhkxrLrb
XCaG3Vn4HHWv5OgLxPS6z7dv3jSn6KbCSqWfuaqdHaxmW0GBo+noMbNwhNg0DTppTgO6cMuB1Unf
1X3Tr/F7eal8e5nXp1FMZAyGutDwrhg6iU4no4RWXy2aGtjif8KwOH3Ls9OVNm6hsX9tV+arM8MK
yf723nkDWimn5QiXfjZWs90o+Cn0PzB4TxT5sFhQS/+SYe9sieMR6AJBopTDw0On1fBQqdFmuMTQ
syj6rPGJp8HLD+L+Qn3by1tlq+WATwtmzHVvJDbGn+oCrsR3DYAPJ6dYUx9epAl/eERPilXize7V
saAAj6CjpleZ3n2OUDcvGUFuy5MNxdK5VJTCEL1C1eyRU/xRsQtV2o1ZVLyxFeVQKZevwhBmTfkc
GEwOZFAZzHs2SN/38E2Pvmkpljh54Lj5M472W1BGf4UUzGDZIBo7vkfSJs+oPp6Kb4P0Zoo9PAhr
ICmzUUtTBVlRM/MI4mCnj2DpsJn9xX0UR8rTAalOy2qkxHUw4pvCZ5pJqu2KBYnX+J98rxKxCzEx
AIYmYadAvsI76FtWk4zb4rGs3ULQUCOTf8UKDrFH5vI01gb8eK8v0vOUQNOTn40PnkFLcbCscxyg
RjjRBEPu20Rr2f30N1lKbuU+M8z4SyMgJCb5s3K2us8Ep8jveFYMWPPOaUZCaL+CWIF/X/vz5ROb
n1/l48723KAH4GLVsMs2BD5zeDZlhfNiyJb3JrBUjLjPoNdXYKLjfIM1yjfbmwZsUNi4VANeG4NE
tqDTt0PRlHcItcrD59wMA6OgzmWn8pa4kck/1bZMIWInkx8ZP2fdhy0C6DZLbCZRoBCttOYRL+bi
cbSyBmW8XU6EKnJKULcIoxUnaNiyAKqXym74wOvYp2h8Heaatp7qqYkb8bf9gOTbrDE43H/kUisX
QpA7VhyeqYh5zcdm8byQN7Tf+tQxEEwijTus3NZ8l5IuqtnRWsfMFBEVp8mpx3WG+Z++0gJHB3HH
qIsbkecLmnNW/hcvHKTZ3EkmhL/tqNyHau/lmlfI7GAU/RdVKKNRIR0ion/stXCosNPUc5LoFlBE
mI8APDzFl6KMqUOjAFpndb8qCOlyhVjfLJuIRPrgcG+uPtRPAWv3mBLYt0oBiJYqNnBP7SBiXj+A
Qr4+B6oIvElnQxzJRgZ4LPqW9uc6Z0VVVt+gy39at11+zW2LYESK2CfeBYlID3VyJynYBgoneawL
ACCMHdivJzTtLtS87Z+2SA/30xiw2tbVa7/L+8rRjD1uF0tkk6qlHUMBg9dyA3nG1ZFSk9eQUlm+
i+YT8yY0QUndWv6VRv26Ir+5O9yV9HhMudi+eC1EynBRh0TY88ZIY2KHj8o372CxBUyjs42y0rme
T+lVHyGvrE9oXk6ELvRCY4OZL3QA5z7bnAqUrwlqAFczhAhjik1V7AcqQRolLxZ/4XA/ULRtaL88
9XiyjoBReB1+of1uFB+u+J+bj8mF+Z3w2o/WSXmV4aamq+F4DDX+RGHGLLsqk7eo2beoOtxiJ0Ja
GhwZlf7dnGp8+N6v0JGkOpWY16alIqLIoDJXT0rpaz/53mue9tofzBS7ruOBXvZUgNMpjZOCExVY
EfUl0zkqIxHRczTSduHyAO8qGxDJJE0yQpWQbKzHM5LqX+MEWhVARplSQJZxdgYbbpvqDH0FWU2q
O604nigmlH13EUr1Kc49sZaFqpl/wIdquxTwojVOPdM+Z/t0g1VInR85e3u63hVEdoW9BA/JQZfT
nuoCanBXzisCQ2wqFBjRCzMkLzzCHRSUrB1+wc5PN68Cv72suoTnZA+aP5ZU3pqZtN94K9JoLa0G
Zn46XSeIPI5V9pGDoyMR093gtkbHW0CokbcehnCeFWgGG9sAoh+xAfsd+gOFNqkHIaqyfLh6DYpi
bFowlvUDCGIMwVi7oPHSHJqSoqkOFR9g+XvB9mOnGjXmrOA0QD4mLwCIGpSpbvdZZmTz70g6SZ2q
J9QMRoTKXsNv0+jkSArEZaDiIidEaz0RD46OWdtNHs/0u8KIHOoAJVGikFHKV+sXsSYfPSs0uFE8
6/XtHGp8dJJOlsqZhceXeJSuLFK8quq5eoKjoaeLFzwMbXHXq+4iVVU4VxV+LoKzyPitQN5TtoRo
ARV7P+mPMw41GfPyEXCRGfWc+SPKCtBMpCu9wRf8R5Mu5JayCS8VkAIPv2xSe1+WDVmS5n2v0TyK
lGDJaXEQ+nggHnXRP8XUwArSLCbjGGdy7dca5DleCbZH1i9Esnxi/0eysUzO8WES/CsA6nDQm69x
acv/cr1UBLMbawtLVqhtTv17EkNybl6dI9SzY8MdanCOuVdPtpK7yCozR8lRbNlVPrOjie6qzBMT
DAe/b8SxB1s2vZpGMS6FZ0jQfdLBtGKjQVXuq8JIoyNsrLBo5GdKd5+2daQjRvh9xGE5h2cgAaR/
oJH/dc6TG/1rNET2rhRMCE9CYAtM/tjO5NMgjwZNAItmnW26ooA3Ye37xWC+6NjRWB8rjLVxa3kj
67u27vpSy4473LL5cw6ZnLYPQaV4KfgmOp9b9K/g/RzXyJPWvZEEwvoQBiuYOhw7MGzBlzRQhNui
N4OtY65LpOTxRkkS/Iw2RhfvVxM2+yKKF7k7wGOlbfiCbn682Tr9VxpJIPEd8XgpjhJ3PdJfI1EG
z8kMDN8y8lnLaxfa9rpWlos6N2Q6yAVrsLMTZ/MJX5nZQ2cXOvkjeLPziaXTPEP172VSTIinFjaA
fGGzXOvTr69zXeplHr5YMeh0PX5BtXzUZ3UMzUIZRKactmM8EEjMfgNxnZo/WPrpWwlu56JkLhQc
tcIC5qELltDMJ2XqHAsMdeba7Of7w2mylwUXAcM0L0i2mlnlPoIupRstnLpklGIPhdv1YuDQCEb1
NK4w6IvWelZ1A9ifzRx8yBGN4o0OnMX2ky9yWPhKfRZVC4MPqhBZff0ntOhSmm53pPVIW5S3wqHE
YZ2XwrA3dGQgylDrvZepQO+kvEwU78/Fvx9lBrDmam1S5qfQcDBl/9ME7v/YXuhl2H2d/KEtJZU/
N2xUjZGl9L1WElB3u2reTDdo0EPh2nVff+TBRNLCFkK27Jp3a83A43ttTDl1IruL/SAxo6arNEZ9
Yx+ba4E4xod8CLMT+MsAYYuDy4Q4gSQDkKlU5E3JBomhj9zzvsIPUuIc4gQcanOKrhGEJZ7TVkIM
t0PKdlRdGzWBzRto0PGSBDMrRTU7g3gAsreX/EfdL4WG8pGgL4GNPJJnYkm/gmY6C5or91BzQ2vc
3XOkxW6NgkTxuLtl3Gc2kev7+QZINAsosxdrqZhuxL/iN7BmfNhSChsyavC0VbzmIqyf1nCEUixE
p0faWuP2emFYrdxkd+gK3dE+/cHBLvobZ4tCWEruZ+odCkv/0QCfihdbLL7k94bVj+r23CeDgS0+
OtdpPPdJw0gnkYDm1cDzFzWsYHITgceeklzcYrHq7d1qXumibN6S4CYbKl9s+Kj8TJZgKVab9npK
650QoutaQkFHIPz2jeJQVdlg9+66khAFggy/BZPtfiU4bqCUjpqgYiI6mi4FiD10Ig6mgqqP5tyG
gkuyWBEiE4LJpdQiQZAaduhjfUNdV20M4VVAk70oBCIs8fVNj5d05WuS9u7SHH7gdQBy2Wh21/RB
bu3YsXstmHc/vap8asE/ak/u21XPFUQrkfO2CLtr1BFJAg2O9Ddi2Gqi5yetCr9B3yJHo+oHKErb
2ttW1wPPcn71uBpgZAyOixDlK7bvOz4jpzdhOus4VvhkWsIOTfr6aLs6fUPZISJgA6uHcv2u93pw
C9bbrNdP9NmfUtmHvxeXNh9mV0Jn7cE4CqHMO9tKsOCsdiQHJuOha/8k3YqDDi5CubN2QacAJ+fZ
+StKh8n09leFAuUVMBSnDGvtkJxKeA700tN6HCpnhtolGC7w01/OVew8TZmdRbJIhzcvJnRgdMzw
EJXuZ7NgMesyKfYrsBPVAZtFhEuf66gPbu5Ffzc4bpjUJVOCDlGgJ66RlJsZhp/GKCxuEFLOxsYy
y5bAUcxPoMN9dj4L6i2pv7z48FPVTEju+jh6tu6/c7/co1gr50cRu2MUnmx9lTnrTrIfibeYdTfp
5Hq1rH4gw7z88T53poiKwYa4idbqfhpAktmixVpgLWOh0KDiDZ7J6SBKfs74n73EJzDMwx3Fnvlm
WTz5KidBU0N6j3jnmeKt1LXxKqWhB03c6rM9LoRU3l2zCxklW6ZnGViDHjuyqF+uf4E1fToY/0W8
sWxiB5/fgBF7nSAG1q6zhJGHaLkWedv12dmRP39RqufqvYeWPzzqQv2l9q8L8r06YSzjku68TqSb
+4cSQg5ytxtTEABjdAltEBQwup47ObMP9UxCiq/gQqCkaOSKTs2FNGkHxE/3TrinFN9v1KlbrxlN
Fw/6YM0RNGhTvNewtgX8iQuOw4iw67T/SNEVhQMuS0wT388svlETgfqf3MDffIr4hMYFVE7XquG0
9dHcRChG7ly8O0k5YIDXZKGHeuqrmt3L7K4aUfs/FKzEUt3gXX/IuHDLVjI8fB4svbxt7ldb1Zvr
VKZq1bYDUcaXNKDfm0pnfzy1EijEtSV4j4gvd2ghsaaZtQh2kFt+srfJxdoPSOw/pz+ydP8VoY/H
a+QDw6tfNK09nlftbAhTg2wDZ3/m9qVAWjeDnnNgAVi+U1MpHMqSBPpz0/nf35a4KaSLj5bjzJz7
CkWGOk/VOSn0VqllcdYdw+mCjX81pJh5Lj7VMMC/XWipGUDws+qpvbOQypZ5rgKFWyXp97GaUUhJ
iB08+7rI00HxS5vKQFcdduqGTnZAOgPsewTWXjIGJGSROy8JORmtUolD2vWSVkle0xqu3i1Dw05H
BUb4m6Ll0qaa1Q97spIhu8LHUO8vy8ctU/wY3CjajJwDIyaE1NsM37WlHsx4FDkiUf9FUO2wWuSy
Fs0ZSFagvDxPr0K+iyRbqasRLWwwnBMzCmZ1WgJ8cnx316Pq/y00EPDJF7fmXLU5jzso3KRujnS4
KHl4s2zMLwujsnPBdiAAe2Lt9hCJiNmy5UJqI7vt6kRz3TmbqneZ0h/4KAj6VXDzuebcmQVk9fBv
Cyw+DVnqWXqYxNjxLVJfxJhfxg8b1PymJN3KqmN/AVj1KAB0ZUomocSZjdXiKZkYfknKU5hAyYOx
66D+Mw5rPrk6S7NufYUAKnHg782evrc21QOVpblE8c2WwndxA4nXAi1FdzY1IDxbgqLVamd/IjAN
o9lom7n1Uo3nMcaoCsVwMTIvyFnVJfjKzS6Ah2uAR7gKvd5atg0wNosmOmK21RaSX8alYQ96NbIv
zd0nFBJ1+tSc0CjVUzH71c3NmJ7LgkW89HGPGcVp88RNFS/6gA9Po6bdCzqo56r7cjl1j4GVb1IP
mHdqVm8lTOkMbCDmWw17sHJkwNngLT+NVndadhJCOn2VNmaoTfGrf+RhtbxQqE+okgjIxa1Ygu9e
b0gd0XLr+w8Q6jEEmDAgiTMITGjEsRwCV+xwt7lGksoWggquIMdxvjL7y64rjsbtoydRkpdw1Txb
dA7OSL/0AVv59UmDgwyeLhtyblqBeu5PN6RysVEqGFF/WNwB0z0klUl4yNwI1kIGp5G5VJM5zMr7
+SlMrcdktbCssOHeumCdcsMomeI6o2uzZUk0nFpvNecTIS5cH1touc6R8+nXEizFXjy+a8FccaDo
NvYRQm+EslWplVsuTPsSi6wRcVAZDT/Q04gec3DU48De14TZrUk90zo6HDCVdzR0kNm5JFjeincQ
SBJQBywr0Ugd/NDO7ZUpZDc5eYy3TAJ4CJqLI6I5WkL+Hyf85hYoLtQXqOOulI/E8ZK95J3rJ0bD
vjRFaiS2yePCi/U8O5AOIXmIdodxkg9KlTiUEAHO/wYqK1+twAK8rLyTRIfhuQeZlyZrjS1mqVUj
tAkGt6GLqaan1RXRnUkLuc8oo5hE/j8Hfvq+RQXRbTJrcC9Z4Ycr3L4Dp6/3lxPOO4NdoBWh3Rn9
LDPWGiEaeuwGV0J3Ifyunfj09MvGf1/NVw7pdHwtuFr5zFKy5cL35No6bhjRDG/HThwaWANpXxCS
9yC5j0L4rUcoUEVgOMncF+DCl88ZRAUpdgpPdjtuVUEA2tpv7mVxL+bnfP0gwddwrZeehOOVyPlH
EwHez2AMgkog5KGnrr34X3Nuk303VGmlDELQLDzEU0QzBihljFwsmOhqqG+F8z9M3Yfmnpurcw3H
RcrUlliznZ5fsXqF2d79shTllE6Xbtd7Tu9/XJfukuDKLBU0LlqPRgUatxkJT6FZqTrKJ1YdmOvr
UfUAblpx+8IsO5eCeqTKKKNuGQEFMucH1OEtqxf8FiNvBeN1IbbbfrP1byVMCOSh6Xs2lBuR8wVR
ZHaHCOBPZ741hQ3rJa8MrGKqn6X2Dz8TqMjWZZD+a+a0/naMFrQX+P16xNu0XnRGx1zlVwpn1eEa
pZQ49pcuM6uhQhCue/jNi0xOuX6Ok2+pWoP9Y+jierf7GzOTeNUf7rw/IPp0Fjo/vRPL443GzMxv
Vi82s0E5IIBxIn5r31t9n5r02Jz9G2R/R8LYrmK3tpgxJQIaUp2jaTntsB7yHatS25Hykb2S31LI
edPzxm1NdxWF2N/G+t3WoyXReesuJ/IxOZc9bFR6/QKX9dsOucFF7hHuRqzAzlONq3xd0wWhn7bg
Sx/hjlBKoPW6Sid8Jf6eLbmHdEr8/ykbdVPvPrJ9Ewp54JpzBFATpsl6w0WUPF5+F+1f5/qeWCVj
arY9LrEwJXBnVHFWau1F6pilSyP0fYmFbzOWT1EB9rvvVaQkFGbjHreE2HV5434D7/6PGIjtQJxI
aLGItPkHQ1uxJUEeq2b033RjuSE/3j7Ewv9FQSCANT4M4apCvaDl2xzIzPcbuuSMfzvggzLTM0v/
O0rYkjqCm8Qhfg+Hrh2pA3X80id6TuiXkFsQdSiN7Rf1qsjhXXC+wbUBgCyX/Bb3NXvPjbJbf6fI
maTdyt3UxITUMiLqukD1gFoxpYaJOjHFsJS3eyG/4x4tiLu526bltcY3X2EEZS3+WOw1gO2LOx69
O4d4YkvIgNDq9T2RVym+eCHXFgd5/kN/TRcymK/omjv/UsIB4AqHZvqim56yR+aKTCTTmhfmwkNE
hGnj498/adTpsvORRphICFUXEUTO8lQiRubGkmH+LzBqycTj/hnX84wdcekNa5hXI3TA0htsCBIj
zJOsHgCl73pa/hbrpmSU1lpyClzP3vrDgjbJA+UL8SnESPZP++BgUmdon+/6a/F4HUi2/o8nIUX6
sxzgxNkr4h27Gxj8DjMlK+CrxWSz4zoxn0RcJ7MJrits33O9KcL36v7eTtSVcZvDpsAOEvVR0I/g
Ks8HKAnPT0jSLZFEaA6gTz6dNZVCdS4FRLmxIorTytXR09Lj1LFfzdOnENnD/uxYvFZNZJu/0YUQ
8tmKmWkQzNCt2K6GVE3qe8hGrxtlBgXWbSneC5x7/ib8NYZmHQrZKLm5X0k66eBAYbN/yadOhdvE
zUxIjiNk5A5CZ5MxQx6nczKMnmqAaN+5V/We7BvPVHuVyquyK8DncFdE+PzvwNSX+ctExaocwvwn
YFtGmKYm36Vkieghh6m0R5tb5llntyfNfQzFpMqY41536Y3A0xL+L4/DPmujCGFKpgh3XS+I/pUH
gNRLwOjSpgrz7WESx06maxOqF0JIycS0XakqtPVKO5fXKkXDfAT99jiG1hX1+aep5GdfE2FDynmv
dY9/h31bzGjDheSvr6SAga1mDdlrXqiMkmEMUErB1I3RjmwZFMDj1gEyr2dmUBv/nNziK4kMOxzC
5l4a1HSUtMGH63Omd851dcr2PN6DagcEZX1Vxj4T1rlNT077dgSwglsGyiWegXYBxSs14tNPsLsT
1bb8R4w2eXf0QI1xYmKQpdgq8WJADU1MTQbusYnPfrfxJKExixO5oVpTnVLge7Kh0HFr57IvxYTh
m+cvv3gaANMHY/LvHriR708UrWw03rRbvFloMBfR3Qivq70nJv9p/9lG1V7eJUJq5kdREWXVgLye
aF0IwrxtqMlU10TnjTJXp8KBYLCwNSzqeD4x6+Zhrq09KHIGgcvWxOE8cH3ZviTFVBGu21TjQweY
oSUpdruFuJxSKYTVOupxRuDnz/4nNtvfSOcsiYZwuom9nLqQjuldx9TMzp5c1WQZWbDhbPYTaMwQ
rvYTMVMsqCxFHZNATtKgmXQvcBXznmQAnA9sXfl5aPPneauVOuVAMi5rDofwmzyLIu+N95Zf5hn2
ZXx/MhKBGzcjkANTtw8nBm8s+IyhlhBgj4n0ZkeaRoTmIoB3Bx6LECRuETFIiRJMBjl9T4k5fB6q
zJPmG5odCAbZANf1h/szdAc+anBjRhHwSACzAPbL32F5TX73638CwR+95/5jTpkaO7FDpev1xu6E
fpFO1oGBst/82RR6n1KZcS3ZsE6Oy2QE/wJYrSjREo3YoPXHdwcN/TwtMw2TSiFqwmH+VpzuqHQB
16/VT8bgGsJBBJnmzMu5Esq3qBPXobvYOjq05x/qIjyi/JfpsTteqDD7f5W+Vsxm4jlYW/UwxiLm
JIng60jOelMgZTmvEfdJtYOQH5ESsGB8UKloxqHGT2wtVdzKsbn+h3TwTlN/KfRgdL64L5ESRXOJ
xqf9DnDgLY15e6w90r7lAcDPwX02jPNODxh0BOtC7E7Dyr98pPuZWUZoIxAZ9S9OzaDFINM/CRuU
9YmCTn0J3EELmrzmQalS2kEdqyFjOUjndlNpJCkAAt/aZ2Ea4RWCll1Fx3IObQ7ALV/HdDY+BMdQ
R8a+MTedtBlmJO67pka9cnWWVmvYO/Ts/Qeno2mzEiXjhymmNo3iBdZbPoyulDE0oPTuEGOXED/y
HPzgBHJdQrGuld7zokaWJ9mdVMYVdvZnQ6o3BiUO8Gg8BtaZ1gRg1kuNtPlrzU4ah3Nu0g+3+DB9
2v1EEgFKBrLYDexKR0VyDFijnti9RxJHr1rUF+YPvY8dqfv0/0OY1e2c+LUiUgRP4trw1Pb4+u5+
1mC3wkigQ1yjY38jvYHsxEUuHcA/3S1wNkpsy3Kml9HxDigrOKlZi04lPsqGTpF10D+kk0uI1WQ1
h79mM1watQDqTBxI13K2u73GlQqNGJa33AkatB9i7H5ZJXbFlEmQh9xmZuFT08N32aJQDqzKKyUG
RCzXOCx4hChN5uzrYT2WRpSzRA/pj7kEDiVXWTJWaxZ7CeBEZ0IOy3P1cSlAxA5cw+w1oNiiSedo
LsCZgciH/4H1Zd5GM5lZ7ftC6BRgDLgZN3mW13SRQH5rufc0D3h85ySr7/joSvrNRlqeEygMfmG5
NBVh+xDC5rtIBMoam+K2WChTP84SeUueCEoC1wTaiMUjQKDzFJedWAIS1o/jC1MgqOhT+DCoKKYs
ngUC5m99cGlqrStaqNWTllq0lTBEWxPlcc183xSbR4Wd1mhdAdn/ZxXI178ICoqR9IPvteVTg/B7
xHgwh52D+vEnmdkp/79h5IA2lRlqoj28PCGt5YiAhvnC4BYWEkOejvpco0gvfUJKI3PSf5or5DYT
mYYWeTDYDPOcE83yb/GtgVztgoAiw97NfEEkHEomrY1lmc9QhkSyxWbERlb6Y6BhLt8h1gaDj3HK
m1yGlLMC+KIXqv51m+fRZ4/DupberfniWoq4lyPYzG27zAprbfrjuooJJ/InFLq1LCoW3R2U+iz0
veYTJsOTsc/DMtCtoPgjrKzI7wBdAEXjfRIgyK/u9uRMOLus5w2ChGjHSstLUWkOlKtlp5Gp+e3K
C1xRVS9nTRY8TYKgxahnxTzDmnOuVmCLwELFXJjEb4fvDuByD0GuVCpjGIeCEJhaibSjEylxWeHC
14lEuvAo2obUU2oCU9hbz2JsHfetuH/ZPKiVE1v8iEU+QcdkEbyzfPaeHdqcsdXAHhqd0D6TD8Q3
jxoUy9ZHJBjrCXGuleHdkeJqh+dq2AXalWn5aqW903RD1GKplwc4AIrKnghcc0z/p1I/+FrreoG4
oEr2WLRlBfgUW0M/QMIczKPMtPJ7oMVJoWJfBz1vhK3oEI7TNXz5ALBQwqsYI98xbZYJ5EzAnjom
ojJXwJrDyqW5zBv6GN8zXnIugwe710JJRlJFyUpJLs3rI3OgEhXE/dv3vGhnILBOLSqKTo5w30ah
mE6fjqZRyshYbT2Jhf6XZ6Dc/tiGZhJT2Ra9H2fDBo+iKywqModaa3bSl0yOflVdgc9gm9e7qsY7
Lk1+kh5gOalX/85kh6RkMQJJbAaMM8BcgLUDtu5cgqRZ/UMHfJLXf8CexoYbJPD9fflVA7xFdyEl
phwANSc9uaLNJO8dX3dpXTW70ALh+n7C4/SB5nkiu7+K7NWuaRYVYsIuCDRw1LMj1H3/zEZFTjsy
fg040mxDl+S3h6AQrJEGr9AkANZStfpe6g+OyGSJCzrbyuLbn9rlKQQ0V2N1j9gRjcqlL9vUXUCE
9dhXM2GevuLC0l4jrfL6ZlgZrR+qtsExLy4c9xd/JS4G0inmSmslrPf04aidxmaltP7RIkDt/EZM
33r1REUI7/nY2SXCDDSdd4xDptEi6I5OObO9YxuSA1w+IF/EJHsumPHwtCVA/Wsf+EHSsqG4oQnj
92mWlbbryWkmDjyR4L5gxdYcEufbcAIwL/i8nFXh4TZISXkFWXvcC6yfpKjvnA9E++daa331l9nH
eT0qSll0IFrtwcKttSqXZncEjqLvbLdxejY1rA5wsudNWPpFvHKKiHQkF2iMtXHA8VESTauDj1Ne
6rgMVfg/Bai2U6sDvSDwUWw/Oq1lmMS2E4Cwaog70ldWz3KCwN5eVMPyWtBUy7ihjSa8m/13T6LU
/gBidmvnvddeoniNdwVB5JglFWabeIkLbabHVREym2VbEglREKsGluKZSuC08oO1Cu2YLLdLXcNE
IE2xbJTINnqcFIWeWxfvjr7QrTe5ZiYbGxp5dGK4+ujxZ9W8OPKn/q9hSgdKivdx0CRbaIDA3zeM
P+TGZvLzTnYohYkc1ww4zXag7obyTJJJ8kXf96PlIR6f+aX2JdeydRA3Utd7X6n5uABYpYkW9S6O
Z4wEsfVigBcL3+F3lBJSgWVjK6kQ3ze+3VmtoXB3+spAW8vPmuoqT89vciVVm48iyBpmoSaovzDY
jpkSD4ehBr56fFhOhpAS9XuosDJ5QNLsYTVU55kGGv9Gtxy1Yzgd1mzGiJZQvh9g5qk4sB0D34Sy
VyToem6RoEXohux0bIaxK01Bbv+X0TfGzWGvLtThxEZ43Kuhf9Z0VA3OsTPtH4r7z3Aryj0WcGPW
IE2z92Ae9i3sBhahtgX/y22J+cq8z+jzwNFZsTT1RpkSKzA/VkGT/XLzPxpEq/HS9Qxpo9wDVuXn
hscBCDXc+YLpz1GEXvMcEofr4mqmoBMobwf/suR+qFigxLEEdBYATeZ58jhF21hyI60OS0lbRrZG
Mr7bB5dTprPB2pBT2c86MYPCTva/N5k5gz24jT98Snt/kyrKMLs+Ls/OUQYJy5O/Ue6zuqb9zZ51
s7Q3+ZS43IRaKe+9lsPvs8aDRAUQtGRls8rtQDMrDC9ticaKTyqK1cOmzjSFyddFQOdBAncg2nkE
n74CB/pKF8PZ7mtTPrC359Rc/pr4AOx82nK6L/HPt511JXYIiJ3oxWnlExIwg8pBcd6lhxk8z/gs
H48Dgl4Ih+ie6a2tMiFehfU0MsGxq0wP2s7Otl1Kr53bfQOpl6o9LXBPPC4FEgcfTGL8ofpoPgFx
5c+/uyk3OhaZK3z8MJ09HExGz6zuFvi7GufJNqrA6OEpY6+p5l1W724yGkBefAYsmYxAeoZpEJpf
v8/itolKiykU9ghoxuc28iQPmauf+C4ZV2FFzkbcKRAtxPgOsG1L+RvNHX2JvWJMa4zwZ75v+V1I
/8cWn957yxKepSkurNnsxRR4i2dTtW7AhI5imle60zCXwMiYczcsS5xtYMui+BQveJIArGySKN2J
ZCVzn5aKUIL/cO0tUuhTIKqbsJx1ZQNVxbeBEPbg83r89gFi4735WN5j08mEuJdLN0oHcy8gnlgZ
rPLXZsUTi4zEx+biH0dtV1GRXVwJWc9B2E7SRPT687nrTUTw9fp5ZvvXDlTtIxX7GmJdyVHg+soB
swVVSjuQHSZYvIEF5q/G5+1LNbGaQmh+H/Z/a31A131G1IzQt/z8ZSr3sAF/FrB2FCWe4XqXTNnM
cckOQ6+D2EkhZ6kxESUM5ea2jPbhVmUgZnLF7NDTLNBKHpNrs51edvfZGMkqC+hRCrU+06iTe3T2
D0PQT8O9jA4YwARPplAUiw6yebFODk/n9x2YVIvP+jw73+4qn3faT/JJ7Lk6NKFybtaRo7LjniDV
Jc+ZIgsiqYI06XbHHfO+XPMjY2GAP6iNNLbUU+9O8s4M9MspSScIkrncsL+NoKy41Yn8BXxtd/Th
nGrvAB7S7suFCJc+nTL+pjFND9Pw93CnbVZyixhYGR4rnEOSlFtnKdLVfmXLzJSAF0uBKDmjIBUf
1uAmsB14E1/gW+rQdglaB+4u3kjsOahFOjLQpRCu2fMe2sSJ9PnA5tdwdvKKDRa3UgCTc7eh4K/d
AkM1px1c+kmcBWVGAz4cxj7NyUS+ASPXupbSoo5vhmnPjn9bJS4zSqxrbJbQB+3wuEJw7gaKl1zO
nDu4TG2rmxfNBlLbsqo1k50sE4XegGpoYMSosX5tKOOGLn8GYCowhiYtOr1uBqdDa5ZSlzdulDS7
dMpamHdkv1wlgaAkPudZ23cpYr1163K0tZZIpLx0hMt3dAOxQNvb9XHD5hMHT8jQBN3Hs++9wHfu
TXO1z455aMmX64RbO/9VxuHc3ZwbuBc9Gn+11r7jGLaSGEmUKTg+uNy2etsV2bbTFyC0oV/Rm5vA
w7aVXJ7+mGwacUPcTC/YYLwRgeukNoGhuKbnvZtOgVILlF6D2GlcaQcPcaFfv1POZWm+4sTz+0aG
AEUPb738uxSFqeZF/QSeoWpg+xw6Yw+21Fks5NAavTLz6srbKLZps8dfdkZ3uSTDNsTWwWYzzq4r
sycAAWfjK3zd2vPPGa9ExkJxgcQg4Kyq57h/fRZQS/2fBLMqPXh7nt3HcrtHgryzSsOIaJIDQVNJ
m1TjHYv036r5RqAzBAJKIvzeDturR544gbkGhMo0LLe3QpCkz5cL1//zn36GV8rXGQsAkfS7SStZ
HV/J34z/n26h9773xY/QVFnVh59ko5GOqzI+690qnumSXGt63VWrcMY61EWcPGqWbxGaPkV2MgU0
ZvohvTP5rw/ZA8nwiCDfaiDJN54jnkvTqyqYdiG1KZa7Mem8TYsqiiucsYFj1zcBUFNuwky7/Bsm
GpgiYG3EyEC7KruBhTHNsGK4efXSQ1A4v1We13Qd7jZnmtQMeXCboVAAg88+S9ftcQ14iX7rDJy3
9TnnAnjm0Ht13ZBRAQLHaSwZ7LRbrx31WPvu8oVbQ6dX+douC7q3fgvlQ+/OHQrLnHiuDinxLo1v
8VdatN9r82jKkmtCBCR73NTby4a5TBuFPOTYbdl5+L2ABZg/RG59FOyMDD1XIdfsYexTFWkHQDPS
8v5VjTCPa6KKfFVqOliQqIZePHbsjiRG2namQu7+dE221IB+VMwbi+2Yg6WBuSmpy6xyUh8YQhfN
sx2B0MjRQ18ul8zDVVPNcV/PR5vj8p2iLfGy4O/FMLl4MVRDiibYVfUUW5S8SVKt+pPBE/iyz9lh
N8CaAK3gz+pbTRVj3HGz3UOXhu4WZ8ya/Sn5fZ84S+DKJ0vfy88534CwuOImEgWUX/v0ZyXoCI9i
x74k6lWUK9s5Ot3oN9QapSefKsmSOEBBH9vC6v1H9LYBYPDTB5PRmcXjNNfIthrU98qgBEgmTGRi
u8jfgDPWqBK6OHBPBxUZu1qCG+Ofdq+hVgEC6Q1SPY9ywvHKxhQnRWoFKX/5z88oTPSYXe3VjFSx
wKPuvq8nBUSpgqzvdbQ9pRy5UaUp1aluouvTC4t6/S3lUc/BGN4UXBxD/sLvFgRAPVQhW0X//EvK
txZEO5LOCh1rJC0tlzz8DXFzT0QPKbZY9VGk3YU3ModBD5uFnuJiyF0gNNPqSuh1RPMej3adSvVf
RfrSO6SUoaDBH4c+ZTjJL6ZktRBevJ6jDLsnlgFbkKXTbchRalwccJrSq0EryVOmzfycPrL4Sbki
qYdFFu8wiJ9dosxOuJgIb2Tu5ZrD7sPsTxGHJFADQlrwGHNuvQzld/yr7hDs0pcbqnnH7aPCP0um
/x9iUOwD4xVD+PDDLwvfbMHaK23ZDqt8F+1VHJ4k+60YqTE+0UK9QAVWAmsryknDhjKybE1hUnBy
gIVqHsDqZzaSTU4Y3VWaGBs9Vg/+hzUyf/8h57MbQrsom0uKF7DbRr3k+PQDatiNEXF2Wsl9isIX
7ye24djWUFhqittjJk3JZ61S/tY3VqPV7gKs0ZrnTTnB5jEJhUcjt7B4bRzIcUNsyqXOLVbOtwoY
sDlHjjyHh2zD9oJk3DUP31hspS+11dZ4XrxJMyEz4NQ6V4IQ0Srjd1lvB/qjHT5qwxLdVCCQQOhn
ejMPYwzJPxY2BQ04tRyLSFPCKQZiK36UgWGx7zjWeZws+MEBs/heZebhooTcR0tXYwLQZh37OckU
84/ATJfCrVJV7ip2lKTlIzV0amQRIxB3TeaROTXfFUshMi7VTnLyxxRwcAsPFh+ir1ZZaC6ZajyZ
nVrEKWQRg3vSRpwTom8d4JRUIY7eC1XlBmsP13x0pvQwq0AaFSL0+8U35yRiBe7BXU9DkIbtp0u6
RuhVVMAGG4YrYZmb2bBiUmSVO5kvDUbYI50W3UV3waZU+v0Bz2RO8OHsEiv+PhcRHfZb3rRQnmqG
WDLAXWjLrzGtJ1nojkrhF6sNGQZPBelgU6yvNhwt1J+Y6C0llKztFPNVk+yx4EdH0RWcmWurpgAt
VbMNtvjhcgFd2pCBzXhK8d7L2PsaEaqM4qZOWSI2qTl3WlUuIdEbvd5Z3zK/Vr5sfrtZJlH5eyxd
aCvrfuk81Gx1MlKLBYQdQHTRpsO4nAUfSzdMBJAUJGCcqyNj9vEAMwWMsqK67gdCUaNQrQSQbK5V
OqlTWRcISB2h7EYibw2o0fZUWxt6oT2SaVRm3pC1rZHj39ORkoENUh80bQlRwI1Fz4X8Hdoxzh0t
vhgTWGpYEhjmdNwB/jjHXLi8kliwF3L/uyTcFGGbBm3UKt9uT4iV1DU8gsxmgYQSZfOIoN9PWG8/
r1SsrNTLSJiH3L/hXhYyxx7KkhOcc4vw4/YmIlfp+otQ+kgr64SDGZzd/098kgqaFllryaGcb/GO
mlafLmkjWdoesLXmwXB4mhkUgJvf7VZ+DJpnq2iGm4eRFi7QdmPzTTaUK3nViCiRBR8UbQFu4JVx
gGyq5TBk25Ag+O5O1tBiEGKdYnycV1AyFATL9h3fk8HLR73cMgNqQDSIP9rLXGj4jzRRv514ePAS
k93uO6Qjcq8KJREb3D0mP+B+qgQULFitYx8D5ZxqVH+lf227h4xhHMZWNsR7zy9ZlIx3HRVMwgpX
1ct8KUID8WDIbTVbfBE5xIUDYPv0rElDMQHYB3ZeY+0n5Esk+DXwZGafKc1U5KnQyctQxvJPUu3f
7HFJQ7OMAvgeRswIwaFm+55gZe9QMmUJ33RfRtOtcC1YOJUQga7LO6IK1rqQn57/lklp2FIAnFPB
Lwi0vKRsRhRewT/CAOtvb5hED6aFsv71R5tpdJMslsQ2S40tVi9+11q+/jnO0uAYWCPL3bz9y1mG
JgkUP8V2ewm+nr3c/I51i4dvP5cd33I7TliCMzDPZnCSOoVFE9dlHb2SFsFG0qOKSW6tbmYop52n
wKzW2TmSdo+A8JOJTiFLPQd9U40Z9DcoOGqx5EbthCoTCKMdhIZx/8+FFZS5CeE2vB7r7vVwD4An
QC95LYjLD5TcACPMzm076sjGapBaRnYcHAR0cInXtywoa3xRheEdKMuwDIulgPU2jQMtNHj1aajn
OVsplxW43NA7k3TwpmeeL05PErh2fot2xKc1XPVnMzYNLIp4tO+ISqcM4A+3gnPJy5oaJsl0clEp
3y7zpaMS3wdkPZY+/Z7mySxDttdtdd5Q+chFAYgBAkG94BG50vKvhbQj1Zq4ZWlTURD59p9xcbpB
DfGGwCj/vPXMp37t3vhs3xov+E3SQE8FwqgvyVuKMpexmg5Q3UQ61KgonaToqTvpRvMibjXi4lsh
pfJlbZ0kOFPYFxBCrdWj5ERuz1Bd+qiOw3w5VGQrgT/0BvTOo7mx9W+tCXxE45ivjNK/MZygGiUx
EJnGwwx3L4ttVcY+M3LWuYxmEz0vBjrLkskuMmm59XXuPt4LlbW0jNilgbAtJHtZZ/ThA8DPOnHn
CbT7BGuQRyBS6TMivM6XifJULvD6V0RjxjCh4K5YF7whWWOqVfCl+Kqa24SU5WwA98vcQCo95YMG
g9k4YfIRC9owsfEHhMcZAMsJO/YUq/5Hi7WfVeyfSMh4YtigtK41gp8AAkGWQsqPiLEp0Huv4MJA
oB0MfAEcIa9sYM1f/7Vp2KfwTFCktHtVXAuAssb21HELz7+tV/+AW4iAfIdUSeIphOT/tWO7j3f4
J16mCron73hPACzPo+Th4QjsWOBYDoacEIn9OB+hnnSaLqeSq4NzQp9aoLpl+KQWX3CgEQYIqUrV
AYyDSHbTumOV6otarzhCBjPPUzCJqaAWKC2Xk1EYT5yxGDUqzcTaWjEYq+J8JLn+f4wgshtSKCLC
BFG1l91c5RKgltgBAFdHRgS9Ph+6Q61ERxRdSVTL7dmfJ5wQzfImFcHsUDuxfZcRmfvJ0tKHEQHE
KMhD+KaVnzI850eUWicsPw1NugoX8cqAdSOub0bLiqfMSCFcS27bwlY2ysdCG4XPrr6cnNX35kyx
NzGVGWwhGKnp5dRcj+LxZw+qN2gtCHmYbPZtzdMxckeAH97eXnTyasIGYemNNOIyE1SYBsECgzGo
ZzrInojK3shdrLVdkhiwi7iNxQqZRfLzDzg3fMNauwZS90g5wUW+z6F5P6vtjjkHHjOi34LlhViq
5qlt8mjtr18bxE+dyKtA83T8jI0nhAenGrbl59djsu0yw4p9/A9GRpVhAFoUENYZgfmfN38bWQ4F
MdB69Peso7EI29icsPq79rJvylbJ0lsln7UeseB0Ktvy4Z9zdTDeZ/Cta3c2IgFP/7g19zHMLV7Z
e7K6mJdVdg417lEh6c5FKBRN9wDrCe0CQxH1PQZiKjLR/vg0Ke8F+MY2qPOg6yXCS6wtB6o5Zd11
Y+KHybdC2Tsj6P3kVE8U1nfe00VOE9SIchOrvmGu/UUzyXXyB+QLbHUrtLXrAcGqSZzQPESNPC0l
+JbPEorTzZ1na18dOVvojZEksPiV/0YYSZJs7jqsprl8GtEC3zkOYQankg8whg2OKWrhuVNY7gYO
sVVU+EpNf6diZV3nc4dXoMGvpk2ewg3/DNX5WrBVeSANSvB0v27SuIZdTy0vC0fB9LNgh9UBXu8U
1oMOsalSQEzniOKPdSwcXIAmLxjdbsNvegeGpqy7oXkhSvGfbLGnTY8rsc/3BdpgLeubx8syJtDy
r2a5CzYqhZwyzrrP6p8DgCK2eu/E1b1qIaQLbd8jdBojQRadkfO0EmvAUFQHa3q+wfM+KPnzR80M
I52rWbbQy95HSxuEiyaPcUnSWERWEMlUBVdNzg/h1EfX1raYBi97EpE+lIH8F1r7rMwRYghM3qRl
NFPw5Oqd0+ogEBebMPKYG5G5E8u9sw7lxUTw41/ieaO49k1B14Rp69nGpKUg/cEpBxfJKHrlPs6C
BPpJ6vTQRqY5PwmJS8zP6sCjzVLz4KgOX+7XfRtYNn9PAlnccoB8MhYq9HnK8b8Nz8cpMZS8fhKT
9OzE6BapStVxlnHxsMIO81Mf93ZE0K+eL0xFEJTfm/qBzgNOHD3n4Wnj9sW3/qqB8ygh2MVHNxQ/
VqXeO7BRg9oRlUXiACb2ls/zbM315byP8oUbZPt6ExVg0i75MprPz80K6NjEMT9VFW3f8GCBiFHZ
9uo6ebCMftXqExJY79zCs97IFEAAyh2bafC7F1h5Be9yB5AX860xyzX2/OATuJGXTEToC6dui4p3
idqG3TZZXAAIxW110CEvdeLEsqUNZxNiTvKppszoRkjeIqMmENC1kueXpO4tJdSLoeG1lMX5h3wd
kme7o/lefNvkwFFpKY2dH8NzereuFTHl6C01jbM8zjfiJVdQ7dbeKmIWOt8s0UUeZq8YgaEs2x+4
zvSois+C71QBmAfqcKDhPxW5ueak11dx2cUbe4855AgyeMlOfmvb0EQ6wvslBQvQ5CLG3DptzVZ1
8lbNOCHPG7VXltv1eC1NQP/9NT5bl6zKY5/2Uz4j438G1LYgtn1sV2Z/PjI9U9MSmkCDhGFBEwxL
Vd91ZaNf7A18KFa/A3mkiGVHKounQJyaV6tz7EG8mXB5tlhuLbZMr+yGAl/9uSuunwNs1aAY5pjT
OJlnSs5egeo8MVrB6q4L/vcIq/KEHJAVbg5xmVgm2vk/gIgQ1a6KxWUoay5Qw1LPnZiBORABQmOG
hIdOglGkdjAX1alujhb0mvepoRNdxXHEtObqHMyOz0HcCy1BIBTSdlFLtF5/l/7H70V9ax6gN2Pr
Mxr7ww0nTuDXu+Ud1SDcGXwIzPIUdYYnrs2jc0knwjdTx+dKO4AyzsBMHO0b9IKs5VMK9f3XNZQC
ZtQJDV5VNIi44MAaBTCF5J4bkAzVRhmuxoYwd4HsEwGyt/pKHmYhwzcTDcs0d3jpfSrP1aXkliL4
imKQjfoZs4jQVe9onYCVatGGOQuRNevC4whwbSQSAa+fYrKOB82tMrqbUdKHZYXpGLJmN96C8Acj
Pr+j5WICSkxtOa0JsM1Rp7xUGmo1ugHYF6sLHH2kd7yibqbntOXePBQDXNO4wbShEDZmyehLZ4Ru
PaEyVRo4VDxiolYabWqr/J6Z+QPn0+Zl4rkU+Am4tgZWUkyskRGKNcm7x2nqjqoscY0QL1xDv1Fe
aAgUbgpvCG19Lffvfd0WJRyoyXpaKoDy6ngH7IXBIEuUvgt535mSU2aBVGDFB1HGTeJ/y4gaytGq
WWGzrKZZCNu7KYn5/yEeQrsCc4wY1sSa0rPreGQ3Dd3pARD7yI5NxnZR/6x2OQV7tyjSjp1hdebH
lVomQeNjMIFtJKjEmJOqgmJtWQksBGBbomGxFxpCIydyQsWbmZTxVB8M1WF+f2Ka1qbw/itzKlNj
IIP4TvmsYKMTLaOg03NZF+pk7cCBpTCaXuGenqIoJPlg5x87mR2lLTyPJUrucoP1uStIwTpZ15Y6
3oJvg76YDbjQdCEdtr50MEJyzSFSS/uw00/Uftvk0Dy5FzxNdiLZ8Gh2N8DewmjbGjLmTlsr5Nev
mT6sTYHovGZevc6bJ2y54+HMvUthnb6ys19UnMyWUc6Y4fDdgVgeNQurWkNBwkuGKgkIpW64hYvK
gLn+IUFlt94JJ7DWvhCPZrCyHyaGxqfVnLpVgtOJmwJMmCeb8JSwhudC8h5FZCqAkrHruIWw5GGz
NvyllgH+LkWOjF4AzQ0KnOnOKllfEGJpXBgZB+aYXLzup05OQpsubEKIk+8fRfc/iVxtKAke9DhC
IFoaltQ9UQVYYqEgIdPcjt96Oa3UoHdCCp4b6PO1AfVEkpcDloan80xgHzRTuCS7GAENGDJFJ7ms
UGvoAv3qrllg0Vm5Ttcg4rDqTY9toj/lDSUKqg+tERbaeAtmjKp+CE/tlEldJyVVmobog9F7OvB1
uUUo6rP+a6Q/yIltjC8f5u12dMmtBJRkaXIGS/VDErZlcV5mS5jQ8qzgFc2TidRnjD8TOuEBxHDY
L/mxIbH06QMvIjhWkD26BC7ceUkg5WUe3UWF+INBjI9+5L6/82TzebA8mmbd2YFuaFddBsG3t48Y
NY3rjeZRt56JJmmoNftveGwUqn40iJuVwQE0+XPA3NpPvSKUTebv9q01eAesd/OH9bPDzCEOkBIX
yogrO3smIiXUX3B/WM7g8y+Kh7MhYZMhx57LnDLXpc5Km6LFWiunxjpwbO1CT1uOqE9l6MP4CSUe
8dI6PzFISnxStH/Tyyo7x1T3F+6E4C+D7Datu7nCwDtlIwDtwjbBzbgBQqNg2mlPwqBVn6ZWeK18
r/dlZ1q/x1mjadpb99w4azsy4YJXhg46liG1HCvc3wmI9Z5FX8rJcjZEWn7mwofabbDa1Bf3c54M
dx0LTN7PCOSutHsvvRT0CIgAlw2Awx9V2F08OdEsM3hBYHnQk6l2urDGG0jUrKqIQILRA/okmGi4
HgeMTPqBjqDWvcRT7S2zlse59eGsK3MUFCVh4CPOyxUR0iCWUveEZaDxdBYn9wre5GRLD1YLttL0
B9F7mTIiAmyL4FI0jwrDc+fuWc4PwyTYR1GuJ13CxwBmvKquVnrSwgcj0JCUnZyf3XdJ30i86BnK
+LMbtUj2h705yNju3cACxS/bKai5fE3u7ar1K7h3C0h7/I3CTatxY/a8oJxYBbGRoQubKB4tpkc4
IVSz6Q34ArVGtbYV6DYVgX7mInQvQc/E2FgllSWFv5NNBFTfUPBFfqiYBRZVSSy978TZj8IlBlWn
xbaw2GJBO7uSn7CvP+rINBfANXg64Pztt5C4bdLe8xpLq6aRIS71jp9WlvGIx2DkbW48PSedpbkn
AGRG2eLXAxluc4xaJZcaVl0D0sxQ+UcyvUO7f8KHrit6LNW2rbAsSwow01nJhKZb/0GymJesUs3r
2ZGhK//hO+6YGwN2dPj6+kRZI5HZZ18ftXfEcGvFU2oMOiBkv2LFPhuf1I79CinRtfBmuUda9tjt
GBNUCD8xe2ab3S72K9EO0M+FRu09LkWmPWzap2lZggsAt4ZHOve3nomrK+amSfLOCw9LgQeHy/F9
KpIWPF7LZsVCLc91F0Z+o8RMsySDnUeu23RJMJ6/b4a8KPFP+5INaN7B2MBMHwNFbIQxqbwRItlV
tnE0b/QEoBEAwXgs2GwjHAV+NKC6wiQjCOXHIRJ3XvM1kpko5qZfCCm2aLHlI4NKoSrE/mJgPc8V
UQTPvfh/CN8BNNUOJ+sWca1unTnTHOlQ5TGqYvRWa2u5tBKJX+pFw6vgz1fs3pW9HY9M6+cUmxzZ
5k8OsJiKIrbpxL0UWJVWu0YHZC95Ij2V4nDb2XWDsnZaa/LdoL5VW3y6q7SOoidyw7CPhDBBlRBs
FXcXdYLu6cRZE8gqKUnj/CQDYf1dikZFCPkguxpMZc5ZYRktuAm7xelIQm4u9SZ9rmMTQkyKVjQP
Z/IlK1hNgPYJZZbBpp+jWSRxsMLZ9bSj7thxIk2A0Ck6ljKYMPy3UX8GOSH1aITZdRpxFh/9YHY4
XkZLNTssHdGo2GpPDdHad6ZNuSSI+8RD04JZhW+SZ2LliHx/LGYYsmz/LohmNfELU1SkwPmZwion
HX8tdIj60m4tkrAcXBEhWUYZ/jMkmfp9fnGkt8XlHnTlGgQvReWq8X3nTBH9IKF0uAywdqaECfJv
tD0C98FjunrqITZ3CuaiE5CL9W9WcYnQXWTAy6pU9bd4ju2aB8tIVPf+X6n9tY/EQSgqFDA20nd8
mHjHlr+R3TYgtDH8nF4ezT2LOsjgXTWM5PNpW1tAFkVusk8nLOx1NWbkEFgJaUy5V40J2mFFdyBF
MPDh7+JuERhXC6wQ8ejKZ9ECZOlepsm1/9PAtp1SbUISEKltH9r2t21GxinPx5YFIcxyo1mfG8v+
HSa5oSDS+WKWHAD/pdMBQqEPyZOQ0N/5qPI5BO63caj/4iMBN60Y87Ok89J3NQrcqGNL6LBnjmBU
1sDTjmcdf73LCd6FYXDQFRqUaTXUdE9uEl1HdvjbvTHkOWoSyW0ot7kxuv+oUelnshf6vIS2JFS0
+P6mlxoStK4/Cz6/1L6DvXGKodTEAecbu0nmsVVviiLnRD6Kn5YV/QMI03DoFuERlyDGnMOfsqeo
JcVJ/61YT94oFH/dPVM+A1QOt/sni80MEirIkvRD6Nk7Cq3ksriGAcwUs/iBptCDjonQZeVodlzk
mGmNzlYp5KuOW8Lr4JOTTmGeaTFVo85r8QnTr/SZTFW+2iUDzKFVV6Oe+Sks3oedsNlc79yZ4I6O
g3VySuPwx4nB/hg9loxceQai9A7mka7axZSvqd+8zRR7tYd6rhuf3F1GMQk1blMm/tbdXDCipd5a
KnAYYUCc9Iu5GFD4WXiAQ8mNOL4c0bPHeL9PF5eKtas7HwUvg63g1pDEUoWvOzuwRHenNFPAmnzF
QhHf3gvE5XPOU97pwi45b/iJBId2U8OWp903a6K4yhS8A1BF5A7pu4ZlM5dIhG9IpMk66YG95H/u
xvIMc2O43NUyDODOOdqjBQapDgb7r1zZfr2wthZVrtoG5ZDb8soribRuH/REwoihhaqqhlo/o6DI
33ZAD1k4H2xngjtS3qvL1KVCsZQzKwNiV5sKOyLsEOXG6Oqxdg0n1pLV538hv/cE8WBa1Lwgx5MP
Y1sFN5QnvT9JhVsl58eMsk3CMoK/2s2bsVKRn1HbCI0RJzncBk+rtFyf2JHioddMO4KtaeKVxU/p
sUXMl5q/ZyDoA/9VkSSPD05LnsjMi/8i12cVvAO6vFGUlllJ34gowwEKq+kP/OLWwF6Kf+cFRP/w
yXFsjFz0mvcqQ2cwj6d8UNJ2zgS7rlSZzG1m8YVHfpcIqVShVBff5HzaZrExjp1cE30JjQA/uqlK
BRhODzNVLy0Q/rSg454tGNm4ek+kFcfjgwQuig5PgR5lD//o2hERWSM6W+HFV+sNS3/XBivILFbE
qxgxbniQM0XQH4dctqt89yTsifmLW4N1sYLQYQmi2PTJK7GMo+zFYyJHPW5r3SC9MyHrmSDGaOfd
5GzPKAfkoVeMm1AFDu3ge2bO3ISuWQe92VKmZCu9NOLESHXITO45tMjUBoWDxYJqS9MOsCMkIbuS
vUVignAo+wLC6hqHBy7WtRv05aj1uBMVKExKo36AosF073Z+EaWpcX87Zq5tVa/2b667OYODjFhu
tyrH27aBjmj0pX1ERNz2tP/z4lX6dvH1QmhcGcMsGwr8n14DE0Ogh6+JyOeN4JJf6HMoUmVh3ORy
SJR0NrqBW9jenTeYBozi84srBf9HpZHb/cQVXaxj/Gcoztl1E3CuMLbi5uAGCQy52gGsPBKyKUt/
fU2YLpbP/OtQ5vPdIHYU9fR1NiIiH7wGq/L/J+2Uwknm8uvTstPU/ICJZJQ5HUkqtIKqSDVo6w3P
g2TFZF4zgij7SMnlKol/R7Clsz8YAz11FZWTchbhT7PVBOYBUDH41Q1MI3wEQu73pcTPrIwtqdlJ
546SsRBTvNX2GT6OesGmkTVTb7OaqR7oB894g/KJ7aa7QB3+b/9UFg5HV7+BgQWuylQe/dUevfhD
VEs9OTL+ahSlhbcILZyqrAF9kfjQd6aH4b4BWYEGoMG5MGnwrvNo/PA9niiAaSKXXAaxlsn5tH1G
mmrN2SU/crSZTIXeSh05c/VP0Rbh0Ggf7kuz2i10vvRLvVTOiJDTI1MJ89kO9c6gMUXdIr64BjZ5
ABT3p2XoZ+rgjI40o6JxoGRfxHnSpCmL5TRt9zEypvdV0icOxoqd91AlxB82TZdnfJg8a2ovpCbb
QBVyH8dgt63LcM6M8vX+n9xIqDhqW2jZ9sp0ZKOL4pDWLJXWOCmI6XZSqpu8hh2EswDpNX+fkMwG
cKxH4biadXeWSNABYY4Wv0o4jyfNfg6cw3A1uo9vJUxSdzEHJlIx2TgaXSpIk8lKfxBfyTUeGaCC
idHufrMLbIvX00uPHXWlflvA8gUkq5ZqjAdPB7qCj40lOqAZqH9oPT8rw/ftDuXi9wagZkB4917r
nMNbsjQp7/4RHC0VpK8I3lEg51OatDnjtuE+lxXGycYDOzgludLTJGqOoueups/3H0IFq+tb0iuJ
Uu6BGfAYwf+cUJlejpBYrSWqN7M4E7uG5e018XDtnlbVcr9fi99lHMPler/v3Vpkz08SAH3jebIO
yV85SyCeKpMc/e0a/UiniRwzRztHybgdwJxtRxFGVJZrx0NLMezuXfIxA9yLRZLjvyTUJU9z3ucN
9QYQmSqtfy2TK6BtOxDq/GXKCUcJEfJcNcw5+NDvUmi5P8HZPTfCr7bECXtj9bjs+spV0SAOGjVL
5764t7FQih+CrBem2M4ZKvnBT6Dn4MLuQ287ZvpTdyMTt3nF7Eq8iA2OTn6rNjmehGWfVO3zbbwP
ovmytn9VbfbMxP/7q7GLrWxkBwgt0dPgj2e+80SsFRwDfwX3rZtmeU25YCN3nJOEKSMHOxSthvWD
mGEhcBC1E+eMCtCVViTXhqpBl34zp3+30bKCADTKqRmXrNbfcPwr7uvpuCTnP67b0GYVtcH25U1/
jF108THyMYIOwzuEgUqTwRjP5DH12JzZlLcBtUKEADpJPa8f83ESrFn2+7F5FRxSWHtmXkr17PnJ
1nZv91FOWZQxmltnSt+n9+JpxNlbnhh4aK7CL4JeQLONi79SBqN3KqqlzyM9RbNugLzmG0N2CA0V
26ZfnhNyvFQAH9w623pDg/QQVYDjykH3HoiAXVqmducSzRNeHmcJNqObiTu93PUfTI3en+95bR0z
NIgx1JZ+MBIFbtf5yVtoTaPr980GnzcOIFJJ9KOKvTqqy5dWkPi0+HcloG5vLMHL2FsanMNCmvqc
imy324g5ffxIICfarX/Glyb+Z+MLS4cwQhPs8hH9OK6vuAr0pj/IGjSZ+iZ9wbsRJYddj67B+E2x
H6LZamT1D0AAIuBdGl/vaiRux3PxhdncGaMvQkaArLpq67+Gcs8WjHQ2HE+alWFC5jo4SDMLIB5p
puW9w0J4B+HKmDo8w/fZw2q36S4BtCtsQG/yH5KGrgA6OrXGybsRNr2yuJzJHlBY1EbzHJle3EPC
k2c3wqS5/9NgOcvIBjqUw7ICpO+dnJsLmSVZXmjG8rAxGENNZAXWUDQJl3nxTgtrodhPEX4R0VHz
8KWEjbgNeGPE2v0Ieo0U3VuIKIyrL7BCzC5IDSkjvO/lQz0xJV/1F688dMY+PgFwaZRs0PPBJ2tI
XvbtL8bDa3bBHfO9OuTSx1HM75BchzPEKqxrDgk5Ah7Af3kN8FtIykKq1sTNinEC3rhenOiSknDw
s73M5UBrUpsCIhiT4IVF42ePGZ8w+ydYUUwWo8alcwLAxlAeGZltuYUBrZYKn4kuM1oExBo4YquZ
LbOu6d9Xz9agATLsIJDpXr7ir8/jjc0E0ZN4i3Mi9bwJiaRqmb7E5DmhUI22f8MOnpO83j7a/Jgb
pDqQL6Lq4+Gm/Uk/3QdxWZxa9Mn/WLqPrehJYoiWWA9+KH36TK++1ztayirlZUFX215UBT9ouAa0
DZZ6B+CwBt8Vx/oyxR2gjw8DsUNMfSSgxMqiZj2StTGi8iCLgZvstZ2tuvOEhDqabgThqqNquhIp
JANxpu9QYKgYah2+S4ItIT1psLTSvzw4KtjvCNFgO1OhaFYfCjBMJIJ/7PS+uIIbONi2a/5y7dj5
yq40koo5vcQbK8rw61JCcc672oHla9mPn0t3FUD0FdWehRn/lsfDnTVak3D4y0h78Ji/GfxRyd23
SSbpj16X1OjLCVL/hYfwK2KLLGh/LbAAQkMqqNT/AvVU1IrXxCpr383fM9sW7sDJzgY5mcQHycBz
Y7V6A0jrIeSwbwLTlPielKc76FM+RrUEJDDI5VNC0FX0QvuloP7CPM0r7iPl2V9jZesRAnjW3+P3
Me9/wqEgDbiQXcbUisguS2wvAWtriPVk+d69dFLTZHfPe8losbehKxbHWo2o09VTYnHhdcMbX3HR
aD3uks2s6bJjMo7qh6TLQLJyYpzoqCGwmDqV8dbJINl3558ioHeDRKcrLbinF5j3m3uiWJuzpZt+
WsMGh+sy+ttwAM/2A5bXDSuPfcOTQ3ZeK/qkOsuVT9UE1w+EVnBenPThGWYWpFQ/c1Y=
`pragma protect end_protected
