`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQGDi5+1T0zt/Jw20/MosUf/BG/H
bU1FHIdsAm6uft+7I5naFNkYDFv6fsxdnfu/MX95XWwn1vRNirzvgSpKb5hcd4QOYknPGL4xojGp
sZ/5G0qZehfOcSBTUwqBYwtM4gmLkZgrLiUWeW/+FNXWDn0NY2ltMbohM50vnoaoynLxGMkjWGST
+ShwzZPpZgxAGOV07TAjXi7/AwOrnFMZ42eElNF/pf2qrjpzbro7vBI92w+dAWBMzWukXzhEmwut
jw13UrJgojX2sEuxFo5hdMbs4WPWuAazJVuoV+WCj7gHiwxyydAMBSX5dIq3Jej9VgA3S+zzpnc5
d+wPMOmwtdFIiLZcNPyTNAMx6qjH2J0/WThErpMXHrGLqBxo1qT8jy7EnyeGHoNcNojZfgGTcfNw
mmuipBcHNXyuxW22cvMwwsVLaOMgHUQaFmqQ9MwN9veMI9y8cKHur9qnQ+PMeuGpBMkzHr2UXcv5
6z6wt1uey1jGm7dDLdCGsoKPtuIOq3ZvzaF+DRlzykJcUcLeiaoxXqWMCPx42Q+i/zQt7dOYV0Tc
n/P3fKJtCG97rYi10xedhHMH4zamBw3b6go91m/j/DG0GEQN0tCtsRB1o3QFnyIOspkMz22oJZjQ
dbOyVQUY4fBH2Cl+10DLWmJana0mSoyjp5RsnYCCL7WEFjEEXCWSrwJTEKWPLwwT/bepLcS7tJne
yEctdDCNPNJYZeprdHWBRqgmx5N2GcKyR4EmH6J6mPunGae7jsUJARSd4EbV+ZCAVWwXl9LH+VgA
j3MOyrPDfXAJDdMWRj1xfojSIHQ6jhoEDiEZVYclSMgnmdo1Ztghz7MOrajXCDRds/2C6sGHFogy
i5FZd8tMcL0ffsTEWMmpTMFWsq8TL+4wUhL/U0gL+7yHswOQsf3/Nh2bDQunER3F/E7PkeEXM4Mu
DqOqz3CrHXfbtY7fy/yd7HsMbpb2pYQ28zqbx181zuYkibc+pl92wYSxjKTLao72Mm7yDqi0LRWY
PjtdZjHT4U95tZ+BXU/WII7/XOL/a52oFqrQuCkrPluN+EDpOi6aXDsohS8f+y7eWE5m4BP+8b1Z
vURXZrQVKrCY2JW9WST607NqBRAf9tRJaP6mGLkV23MAHt4bR99iLJkeRAPh/u284XOd3sFLBQGe
6QAYw05AE1ndFHQYoqWAjFPgRsMWIEScZIDhuLd3pRzHHwMqx0iawUeP+lO9R6Hhk7hMUyZtxsIb
cbbdyWZf8FR1kJrwwrox3LpJFIRB5n1zslCu0gZkJSPcKFgoKJwWwiH8J4OmdhctwVs1xJVN6uQG
U6MSHir47PBaygU4GDM2gUyrzKGuG2VgmNm3VSq7iiOasTDe0erkMipleVsJy5B9waRced/GVdTF
6bfWvRbJwwOvWbV8WI9LeD99MG9188XFQzLnKI0SdA5BPYlG0nq2hCwZ38kV1e7AmCXGS82TSDOH
t7DnVgF4N7MpUcBDkkywcWDV7qqHA1GI12xY7TgXiM61q/bWbpcLSmAUiD7ci8Ij3gT8ZQPUu+1u
+I0r3SCOtlWsVA8jtgAGWxY65mzxwXY0xvQF0ZBGlrBxJ2Anw9zoTES1yLNsDuwSh92YLpPX+lCY
52E11xcNxTVQVqyoKqGqzh/txbvXfhn0oJHtuzqChpAENDtt4HJe7u85mFSbptN5L3OfCJwkgYfE
dL3CISmu5PZV/LZ53tugf2Tmi69QPjyQagxjgXHo56tOqQjdWYYZNyFn4N1YMJRaNWeHfzk91Zip
qKglZ10hfhfsB/c/IUoTI3xICFjUXOU+lIGZdjgkxLRaDpW0z3+KGQ9JtQRhD6kI2M8xxBqbDRtM
aBB4uZ37BY36vwpKI8uugtUUyyFl1+XXrKwA5DhxskbZvKAVkBO4iv67Vcy9lX5OdMYPcwZ4wPow
iUbt7/9jz+LPo10aWf+67wV1QcuXtJSsM7LBYxObW4xLbv95zXDXyErPQJuuwDtC4CKerde+Dapq
aCiIXI7o2MAnbNSzX73WEiyhcKwEoeHUXkLp25DZl4DgF7vuVNULntUNf0uF/ybtzybCBDENS08x
D+g3T235m9USdOo77/sRF/Yzf92xK2XqSROP18iABqci9yO3V2vQsp1ES7/D6BwXJ9SdVQzQfuaP
8b1NP1ABQbN1G8djjBx421ZwD7bzOYl8YBTJHzQ8nKL3ubLzY+PCdDDhUOjb7qTc7YM+34Cr8JEC
S6l3ca1YaCOH0hiQO0shnVCgCt8QMj5BJL3H9I+bruI6yYtHKb97qb3b5OitEiOdWbY/7aTHEN8c
FaC+y0K0IKgQrgoAmVJnZ74RAAwIFK/fj+D+mcUOywZo/k5ZKZkDtIBSM0YJ9OrYN5ULJ1rhGPxW
8d7liloKP1WCMcoR+0jimt24EB6TJZ4J1fwJkYHNSagRKiawCk7XWKtj66M9GdgOv7EAOBThJkMu
KRO5NbzHtv5nXy4mKj97dAekYMjFbocVYKsvMYlEq3+c00pFUeQzHrDUIPbjuuJkFlHNHRPWL5Gx
qAfRJjs0AJVAy7qJfgQav52GbR71mlyimXBb7kvWxqsTOK7VsBoKZB1afteNV21z6hUuLoTD7kYI
20CMNzD7i/yxT13zY3eHrdiYGdQ7M690OJntfhc+UtEBM1TZoTgNk30W6sU6zg63rMBkgZsHDhiy
qAx7I8S0/qDHiwpWUQ9COu59bAyCVyrfNt+cMxQUs/dofXU+v250sXc39tZlkDyTJdlGpnvw+u56
Pd1BuzfVO+VCuXa/ztoTbFfv89YGhmAjsYofocN+HjwU4bU4Xx8J1PuKbmi2ijQSK4Yj1ljF+B9s
vTEZ6WDPCX7lTgZFb0svCQzIjj+x52wfpc1bB6y3r5ucv707ScuK+grjGcFeALyesvCM7k1avhfN
kYGcVRFIJ30jr+ncoVTp+UueMRxJva9mmJ4Dx8Etxw2EFohpDlgMuT4rSbINTq2yxi+I63ZZV29T
vx86v2bgKCt0SDTKxNB1AbeoBTDRRSHsdBn8Y81/D/YTUkz2/xs5uDXTw+z3nqCTvfstU0Sbo3Fq
lzcirWj5uEi+8jcAlJu06gzyvVm7i/rb/IemydRPikFXYxdULwa0okh3r0Q0l0ryoWyrEWHEqAiT
b98xZzPAqnZshzuquITOJagZdMi35ULZbymu8bUfSbQ3bEEC1IX10CY1B+sdJJRA64/vQTP2xLeU
EO2zHD//rkzhE7BRxuABmcuskg96nf3WcBSM7D61Ma3xg96KSVJcR/g9Js74U75uS43KoK3VSTg8
/thPwPrwjzdv6celYvB1bwdqUmiDXn7/CF7l5SwhoClvesUKxp57dtni2JNFBVAi5zB1GY2rsUgv
oEwcU57PMVHGDG1x+xFBtdCVSbqvd95mUCv2+hq4cLRqRO1mq+kPZPZC2fDtcqU/EGieNM/EyG4v
BGzTJim9z2YJ34LSEg8VkHCFYfiy/hxjXFfbmGYjS1wp8osmMq8hd1axkNm0zo0qiBBO+H9K2YHP
V39kY8oQ7p+XQ4kRkOqgX0ShYKOvUXZRE/np9g5rYEZlWf+f6uhSdA6WNBh5Q7kSfCAyPL+0OYdC
3kNbgQtnC11cTSmcJNgs38ae005MCKBSsfGnA3e4kxY2j3q0kjMadzBGWM5fb1rJ3hEivBbDfa8t
sjjnauIY74ljEFrSOEkdiI3rfC1KyRQoFpInQQj2s+cdVJ2cNACorg3jAdd71h8HeX5Lix+M2KyT
FtuwoPrO77rqOta0f+Jy0vAvgu4iPfUqrlOwljtbRc6Nsx60kheJwOkzhBYcoKjOCP188Mkz7zqU
UqMhNw9ZTy606TT/NppVJoWuuzDB6F4p9bzmvE0HDpaFwElchZnkGsqxie35yS6UorJ+UBtR74lF
YjpVBpEt/KqQBg5v4O+Hsz/aCk8hw+t41vMRefce77YupZGC8DuAGmeG8JMEcQZ0WKr6lheKNd6X
zQw8rhy2NVv5OVXg7uPj9hC40BTS/ntmNkiAaxhjg1ajzzHLpHm5aMpwl/Oa+k60dpBp5b4O2dnY
wSru1oecczvez68F3VTbdeM8gSMLmUUxBfrCj5wBHI557yxZEF1NH3HENllUXh3zOuAWJaUioTrF
K+Tvzvo2VrM7USE3B+7qPar///ApaDcrmoi+TYdgBRqZYxdCx0Ln2CZy6Fbq7lykj6iXnxwJO+9U
lQfhjcWl3fFBM9e7pcgy9AJDLXnjUlddY+D4Lxuh1RbrKMVFaoTY4xsffo5iZVOMIEtZawuZT5R5
rgJsw4T7lejeFulP3AcrE3/9pq5ZZ7cAqMm889PrtQBK5pxoeQTvBeRk9NM3RvwuSA5EG1FuCW8F
QWji1SQEJOnNPvmQZ0D+ber+kHIc/sf9oxlqkpJIfE0CSbxPj0KV72u+5kww+ExqCs7vDralsTTr
xbRArTibMwilSVLjHarNaEFtS47FGWTIa+om/RzvHI0gabLCPwM/MlU1X42P+zbVEAT/mfDorvdq
CT3wICL7h0C/e46g6T4Sq2P5y0NGeRS0ONQlHUjcFMQ5tYlZO252tLmtIKqjO8BlfUxLW+QgVbtC
Vm0ncrTD7TqNLS7y3odCotcCj7EjDz7h9KFD/yYyPNOAUtnN0gae5InbrnG/5bc4GnWocAQsGPWk
K0PD8ozxaZykK8vqEGj3uHiRwx+gWmPOlkXFNvhWEW2K98i/mUNEFETJ1ghz/Km6ovrjr7sCsFJL
2UkUr1exH+tnjg28iNNfnE/DZKgT0KGWFpGovaKpkgmBV9/9J/mhJsjurHeIhPU4pymJyFEz2WRP
RjhMAM8vFA9k7wFiCQ4GjkpoufcUXqdQzLZrNM6tek6/tTrHViyJq+CGUl5ETOlYvGrXds+UuV99
t94+X6T8QpUbqnE1ZTB6k1OsS/8As070cXtr3VQt+yVdKrj3/jhBSg57Y2210afieIEFI1AJHvQm
vGSLvqqd1UwwWg2PwagsNkt4n/66Fts1WXJpzxmq15zyvQ5lFkdbTTRBxSvOb/q7jV4DAWi0nIio
eG66K+S3rcOznl9ZhnJP8rCTZjWh/sZISHkRdU4oJoDND0Wy7XHazAZbYSnn6Iw/V2FSVHJXsxX6
Y4MLaSnbUSvri/zABZ79ctRC+M/M0N+sgZhw88wv/JSjK1tr+jHpQ3R2itaxhzoNiTbp5S/mw2PM
aL0pWB/MpAAUHL3cnj7Ts1N+5tSDZGI2llTsz1lcLXWZMaGvtXC/wLr+QDpp/BuBLi18Sxlsu92B
z4BGATV5PyOkGwGQyZu8VgkLuzb8b39IjbCfxfKVIzZegFMTfkUpnG28zYEIi5v53G1O3EKFzdIr
ALMVHHGNZuKLqr/LIiYEzoNtXW4AUs9PbAXGamHdjfGMXA0kGfPXuiTypDdEN5otR7D/3nqRSBnA
CiUeAoeoOMoIoZ/oZIK2Nz8hnbM6EyNfdvt4m+2vm5fbV7Yr6JF3gQ94tabP4atwJUQyCSFoXS78
6KbUxQw7lhIHfos3q6j4ZCcSi1eGW0mzs4gRuO0QAqml86a3Cl6LKg6BUB0cTCkykMI4HRvJJGRC
lPVfQJtaKG1YKJgIM9R/qvyLnVEvVixgpVUHiKsTBDiGnfHv5shT+Tb2XXtJA95ASEmdYxVw6ycT
6rFJKaVzCxzgwt2DbbDS7ypsc3DDXF9cjeSsrl9SEfWJRegS+CSnsdRuwZCFncH48PVzB3lFz7jy
gdcY8ySI4B0J2gHY9QTk1UkgK9+zobjc7f0NdV/9nP4ICUdiOmyCnfEJfLEZFFq/yKgOtHeJiLF3
WejOtcFyq6i2mlfH9Utuzpu+PVUmIJxX2AwokN4QK2Fdebzqjc9ODbHlAf87+AcxG1rHJQEoJlvP
K0hw5XPlIcpd3TSR4BrPeESemcXfQSLwa7ngAQ/RjlzTmRcMEGxFdyELsJBUopVmXQd20SJNvKQF
qZ03WeK85PLA+lRDB1NoA1/AgMGK4M5uvTy9t7T1bX/g2x5/S1lwVugrkMXWdOKAbJCCJ9Qf93Tp
Vj9PCt69cO88B3em44z9Ts8Rr9clm7CSnZTUxuw7tPha0f3EU0WIiNBlUijrRYLlckcXDvMWkPUT
nxRr1ECAaErDXf/txBXgjpqePOFKw6ZSUfmN0pw6ICI1QKNo3GKo+sU2oamgrmUdgo01u2DAQSOS
hWxM514/XoQIY+5+IzWyIJHTVEAMJKHIQbnILpG3EcSqdJaFqpa/3Qa7MBYBJIvHQnonIUa9uURV
M5btviiTcoFmcCWeKBIXBidMwvKiOCP+mjyX1otHRwTZEBXQSXgVCLFd5qevdwgrxSovZubBgBEu
iljyy68aTWHabhmteyJpiU/vyGnnwORI91BrLuu3hg6ENA39A8afAMX260JbAX02om9L9Ij+04gB
TahDcnwSP3MbwwyDfjmmdp86bGA57i0qDEE1TtKGm1RQ23SxokZ6rabMDjXURf5KEzMRKV0NdjUD
2sE5MkWu2Dm/HC9fledKBJV5n2/6ZpcxQGXZcvD53gA8Uoj7prm+irb3XfU6vYUbsXR+nW0pXxLv
Vq/OURWKsVHL8Qqwyk9bKRlTEs4HoAJVxGuHc6YnF0LpK+oINDylw8P/pjrMpdUM/otnf7DAVwY9
G2vF44QWLbR8tcaOQJODxkbFJlbW5yDk0TM9YI5v0zyM9MjXuPWwvDIETIIzWQNaZ9BjGHwkCHb/
vQ7+J626JPmiK60Hg9jvXuLWu26pVdf749PxzPPfmznmrEbpDR33eo4LmMRWxU24Ngf8PhkvBWKI
GJm6H0s7Xdtds6AA88peIOP32Kg264CDzMuitG/aNuARnqc03lN6IirGbJtTBFeta0buCs0O835J
SDRqXtSl2WGaDfA5iwy7Fm+VabeKgZEQmz0N4K6YbBaY3sr+fXeq27VY0Ot+PYI2hJbIHITzPMxr
txI0EPez8xFRSfjdMJY/1EqMV85qKItYTdZZPED6ZhhDBit2pa0uOgw/oQ2NvLLMpMVhehUDp1Y7
e5+NFQlrWvEyQsx+4DYQol1ra7K7TBVf1kAoeqMAElFBpeDdz2y05bZm0pwzTWOIsymRywg+t5SG
B4Up7veZgIUu9nKowx8icclKI1JorJUKczQ8oZFLMzDj6vPPUotEpUcesgAkTZ9Mh+GqNs+UMA0G
1Tvc75YBTdSL6uzUbdQtnNHbQ5ABubZxwRtyLeOoQRsIUmUsV55eyul+oIHs6W5d846r7iqOZ1YZ
JXKrs9XRsnGaUO/D4S4ZNNcZf5Eq1cppzvCLHNZRiKNidZTL1IM9WfaAOku6iS/f1JjMPXHgAhbc
mDvX+AVlILyfLumr9uc7TB/T7sCVvBT89eLmzUPcVpknyjV9jVAVx9gxdg9HuHKC2fuG6i/4utG3
NTLauEQeG6koeJD8OntJOnnvZ0gkYABs6/vcYtNAdsTj9wDD2CYR6o1eozGqTH+A9cyGaVpNdChN
AcGS0VZwT8/7L2X8eAXeqkz4Bs/RKQN8ga9NzykaakQAwA4F+ym2DmZxuuRo7FcfC55RSWNGasl5
F0VdBZlyrvAREITE2YhaLQIESWi5vpt9bHcOAdM+ZFK8NcY4/7ioDBkVYc1BD+8PgYV2kWDckfR8
InYxH7sMIR/tCGu7NtVoAhOgKY1XppOE3P7ZO7Cjty7V3J8hy/YqXHAmA6qPE49SfXBJnPa3FQ7E
Z1EidZTScn9lUrPsl04k0ElrQhVMN/d4CNACfPmWyfzMzQNV1KtixvVivQYDkRUJIGsbZUxRevAU
qPQ1d7VXd7w9ZCUpAUgD1LkR13wu7Gkfi11/yK3eXGKID/CVZhj9GhTirzD6zqitoCcXAdOXbVyw
vVLhlQ9+UPw4vz27aCS6btUdvPOcx9fSquH6mTmnvjac65KJYQXHnwaZEYeumAuMlPtyJPJjviBU
M5/3f4Y2/CIkm5JXSHb2JYvuuCChNI9r3lRS5PFRkSdt5ltkaaMLrBTOpTyjWng+8hWbpA4aGdq3
8rwOtBBBN6EJSHr6lmt+eIxVepbwZmnfYQxv6c3xlnqrrZKm6GWFzMhqlQDxD962trKkknFdyTYb
Of8Wa0qOcKRJj70WHd6XLBJXjr/TCquyAReWt3w5d48NnuSejKk9QD+rAzsixiK+hwzmTp/0kWY3
HD4o8PhM3DMMc+n0uqImFRczm7D9GnBI+d9vQE5ZjLOFkGJ6Tb2BciG6vsrE58ppsMfI3FKzbHr2
tAVo1ImISnfsU+vrVJjsDpwqzDv1U8e171zV95S6/t1RcGQ1AvXpaK00gVWETNTRFHNVk346MKZV
fzJRd81ognoMq7SaEWnoWa6stsfMnSj87l8xmYpJzlccohUtD/CotW+kuvrbQAW1BhcxTHC/CGlC
gLupfqk+GNQX0RvdRaxShXWDiEXp0SJ2HVzU6AZrQ6XrNu6fEkPQuMuHh+sFEwubbdvnNmlZytat
wxRzlKMTQ7wATiS+Usqas8f4197iFilpJ/mIh6eTd94aQ94z7t4g19Yed2skyFxWxBWE0iFSw1De
HOtud/uxOYkZYhWVQTlCd/SQBMF+Zl7d/yG2tZiqw8HA36qgJnR/65zWDoxIancQezXbYEewD+jQ
HjsubVOCTZtYaBWWGPj/Ip5alTdOu0Z6NmgqxnUr1+kood3iyDI18tnzXAgdyB50nKFJYHtd2ehn
FcA2uTp73P5B8XqeeU98bLEuRqFizVCmcYaVGPr3yYZvnYcyb1MpukBhotWjolMwUIvZGJcAo1kf
oNRREVJb79NW5ZI1fJUIsqJiWZ1nYpk3xis0WxNIfIt1PNbqSCLHIzKbccChFKsbTyjR2l9l8KBg
1MDT6ZEoyTPSXeLL3w3mT5d0fvDBKfJVojA/4xXHHlUivDR/A9XRpo9QcJfv/aOyWr09Y/YTPFv8
QXVhaMyD8DGBgtbZsWMZ6kUzV/R6cz7SVrpQzb9tgNrqzo6dGcrgpj0Vg3ppLJOppVjlnOK9icEd
Yq2PjDqDF7EUQtwQv3C/Oi4VBJwR8Ez9ZSLlIlFFccbI0TTCSG+blsl8JeHbcDXNCdgfGi9AtLaJ
Aq3ETCRvoNCK6IzuklfrlXvcP/K48gGJ6m2UFW/v71bXd8RobJy0w2Z0rCRH0sMYzgg3/AhTheGb
VMhMaEk31j4ANNcbfYkv6YNACj6MICTZXJcon8Pdm0QkdvDmbC5HEQdfz4Aq590yqf0nC9w7rLr0
MBG4lHPB/pZlYibEyWgkTIWJ12mjK7cXKDZAAPGbDTS9peYclr0Hw+vSrlnhNDcwBHqnMFkr60M6
USvpuMLpk2VvQleIOFh3TEUI1qu/SRx1oW9A3MwFbNotheUZwefHrdWoEO3KivVVSjf/sIZrhlF1
cuSgjSV+LNimLwGjhGrwiPbMBkOOONuG1d+Cwc8xdsutzwL7W1nq1NmGYGWCZhcgXEEMhqI7eqiq
MCAwezh/kAPD80aZYXUTWGDudQrCCmIVcDXAg9NhSpDeMZsrOLDiZB8LtASKCPYGp4HotINhw8xr
7YvA3oeF8ZJSeoBnV7OGiS8M7+0IPcnVW3qmqqfUFkg7ZcYCkXbSf6lOJubdTlB030ronaoF3Wol
uqIHLbX1d7IRuHfyRxRbebOixk1427C3L1eETom5i7qqMjJfGauvyUqNhsMgxVVoYG6HORkUT83u
yiFaEycqyIBpf+2qdopwVFYIj3QyvUE/u8shAOvuYAQLblOvmsp2xzKHLYVPqTdqhvrD5wrbq9Zd
EVk0aPzgQiWEYNOkhldTlMknTbO6dLLE4no+Kg+Dc/8itPPg5CG/DVj2O/s0uQ0X6RTb0SPJBSpo
LPA09tGwc3Hq7mSKklhsm8xDaMfEFW9KIg0M59NpCbDwv7rjizC6sdmp7qrNhNHvcVcFIGzcbTI1
2uKemKvqQbyR7bK4XxyRaBldwpShd20FmPlSQS4JmXOxEAnL5fPioiuF5oopP+pxZJo1w9cJVA2p
RZ2vhpkXP01Jlubw1NXwdimZfjMU5HNY3CeTAVAByDtPjYoQQDNum6XKFWG6GHi4X92xS2yZP08u
W8N+SwuEAn7dg1R+7dsdlDD3KlNt83Qh7sOCBfAcgFSEJKISx4mUW/DrDqiKQBNJrkn5/GID/Q79
3Xc03FZaN/ViuLaoTp/jmqFqpBa58vmPMKhdxKrcDropBSK5NsABg/OqCX6nUwCbAPevTtbdiCma
bUHW6ns/A/B/4S7MZoz2r11J1pqpnbALVAT4aRIdsZQZwuckGrQmrxwUEvjNJKHtxhZLc/PBGuag
tM+aHWxGQ5vTk0UhAanKEOzyAaqHoXHvpIArhGuMHyHQu1u+eA0j0FBk/zShSe1jw773COAGYsvt
xwnLybhAdqBuSJ0spYAGE3KUqmMESIeV4TWphI7MS3E8WwEo3dDdiac+a3U4J1Pyi7ecxFUcXPzE
HFhoS0x6Ub4y2Kcw6hegC5R1fJHIw6M5ufDEgBJRVROUOcLtU/lTAvU8CeBYo9UWgWEfUkSUUV4j
kmc57Nzo5CXjmiyHhqxH6dTplE6a5xxBqM7ZD9HBWRDwYxkBepym26S3ac4F+wkBulYSehww3DSO
zGYW/HbLopPQv2USYY59iEkwery6iMJ6vuhpvyqBFjQy8ACHnSy9HC+S+WbzZJMA9q+O8m7iy6ci
4VgG8ES7i5krvs90KSUCHPVSXSWHjPzKTVpNsiIQehsGMHtdD7TvF4miLdIvc4wP2l5AlLFrDioO
VfhDzFadN5Syt82csfoBtvpKShJMPKcD6zqRISJ6Svg77vvLUzJGWRuYdZRmFIumdZ5koAgBOjcP
++J3XyNM2sb6j+Ah4tG6xGGOIbdlAZLW8pRkEcbU35AohiIxUF6U7ehHxmFSxFBVuwos/4+PIwUS
Eo3EdCcsFvWggaFXOpsw0Hz5Hkd9lXdvyQXr4ebMmxcpz0TH77J9UXA0QgDVJyZzqrdji4sRuQI3
BSjmSD/tFgo72gPjYjo9LeeApv3R24laPGSnfVh14SepOc7TH4+XRKv+RlTmoZ0ta+zrXBCHmyc1
IzKZ2SID7sR+Duijv7rBqwjQzkUIFh4JDoWmqc2xmbgbfwMp7sBxnSebbx9Op9Z2gql1hv1+tqTv
TQAfV2clmkxcjzyelpf7NEZtfKPLotv+gd6/mRDwrT5+yqlKxbGECEZbRcALGyX5VFTYuipDROdx
8TgaOKq+HYx/oS1Dp+XRfze7vyrZmVln4xDSphJP1juQakfBBsINl9i6i2xVI6uROFYPZtyj+QHX
lmTXTa1f/V9bG3biMrPTTQfyGNXBDiSQU5IQl1pyKL0r7zlnj2N2JRzMOz1HMlVDphd3NEsFw0tU
FE7pLYMlBJ4AqKTz2UgbhVlAVG9giWsCAlhVK48+YOCnbhQUIPYJ05qMNGkkpSFfzzrXgr2j9JYX
H6Wa2EbjfBfPdhEuaFfHb+LaW71Lyl0/b8D8Fu/IhdEazPeAfjn3WEwZMQP11uT2QLLWWiqDBp/X
CPYh62vAQO6xaSHoadZmA4ou7x5R/B/2lJ+AtBf7ZrafQWQl2nWOBsOqiuBPYxiVZEQYLNE4q+c/
je5a2OHBVpxrvOUCpcg8LeE/C7CiearodsVwKadDwLj2gTU3liHmV3YBbSlV042wwLa598LC12yE
lVQRDNbmCaEkLWiykMPz6lXcYdhKm67bAGf2YNAHd+7NxDxB7yv+fgmvUAzQQWBVKqrwdgWRCoRF
I9x0Kwsp7F4zeDkLDM1N5dxSQGu4C8JklqsrDbeaOq44ND2rjfMrOFaI+dfkWZ2UkoEz6K9g3hx/
6irZhgd9XhYdWfq4YvFvQWiUxNhqVTi+H9b5ygzAd6dQfgokIPYOVHnPxh+SevnZrp1oqOUMOiuv
vcByLgRf09OdFqTktHPLKEgRismN4ej1JMLB6x3oSswPGy3UsnZBkYbi7F+yoof/EcOEz/kL4AU6
97XFZr05NhhSP3g9C6ezoaTojY5HCXXQEvFxbhJsM4cs/znb63xtp53+2/eH9VPnDwRzVy8J272R
e/rrtGluZ8VaEU8FWn9GnNK91dptTKlxlh8X+Gf2oZul+2fpT3cd7GjYZ2N6ciB0wox+8cZaQHFb
hfTny/gcbgUN4esAAonhzoDcMTLIHfzaL170w0yilxSTKGNoBnO1qH80RRqC6b7mzzaQBuwgthWK
Q+Lri1G7kPYlb5zZ8T3GX1Nc4HwNOnPpiGkIhQ62WiUyumS8TfMZM2cKyOI2onyjndcPD03wL/d8
H9kYFF5FrjsPp+25I2iYE0GRJVjFGO/9sJLxi6Cn4xvp3bzB3HI87ohsNxhLD+/VUNBIGBlFn51j
KoEGekGGHBisXOqoqUUBz81OdRbpTfQoXhQveuZ9FlNtNlCGVkzT/oQGa7GXuhLTYs5EOVeZ2hab
9fgpmGUMeYwsrGUwqBtnJNVSiG+I1oqsLW6os+Eqsyg0U0mINRcYC6ruI/5Pswi8igMkCrzdOm+f
m48Efct/YINTLbSLw64Ug3IY2ReBdfEa4gGA27zpvbTs9i0KNddCY19+0a4lDfFGlqXDr8F9uZ8Q
vGtDUsvEOGA3qXRixtfHeAMBjQmObKNQywrjncuQtsVKJC5osy/qWJTapETDnJY9fs4wBFwIAY++
8Cq7u3NJBpbejfRzI/kafB80z9EKOPM8E4r8+ywE7PIOt+fv0L+7Jf2kTz7P8Ja8oMLgtAf9aNw3
AFObvcMFV3spmvSFkQy7h1B7oMK3kEdCi6JQEM/El/qZdb5ANnr4sMMZEPtqAiAF5YoucGFeCAW3
bSohjE8/6vx1ZQp0/+6CHIlQ8Dh0z+OgPv9QzCNn+DSdAtJFKsS5K71ks0rxUwlxEyQi7D22YLwn
DyAC4gS8en9FP7bA4yYH13xQ51QGZhnITeo3ToWOw+WYdziJY2C+0O98r3X8s1/qahTksBw9HvA8
8aUnqJ3rRy9cU5c2XaIwjQmHF6g2dbh0kStxp6ozYhtOJYpfyi1bgBhzo7LhAAsj+Wtz0jP+Fy6x
WeBMMRlaVwKSU4Q0TaVPNeSkiaPkPkzOJPH2VmcVaoQgANxrDlSlBY6xTf/IP7WyjiDpQbN8V1Ew
HszRfDKR6k1Li/H34/2LGKxYOKJ0ROxBte2WWGAxFvNCbLCjrV2G/VCAliAv0OaTtSXpl/7W6RMZ
ShLvSAAS8QXJfRMRgDp4RJraDKK7oGm0phQQryc7p6Y6IgALLYPe45hmRGGLr/7OInPPAwUkRbvg
nXoK+J8H59/sIjXEq4SOus4jsTn7BDpiFPqPIASYFslwZpRgGhqzetT4de6Uveth1wB43ThRPSIX
+te4cBN/bKyJlyGHQXNbBVJGXn5jpEg7wPk2+01gXn7PMvwRorvHy9gOFK4kK0mx2r+ZIb5s0qZd
d/VlHpX9UftXdmttFZhIXsVI5TipnjC1vH3ziYR5M2OT0kX3eJp/LG66tFUlEusX5lO2rIC91Ukb
L6K8AUjVwvEV8huAGf6ze2aiT+oi7L1ih8Xi0hXgITHHkP5H4XsCTOHS6vKmu07aZpSjGQ8OBMos
Vo4y/J+W0y/eII6MBRTDgCDWFNscYDnvEHXuX5UaRyt9jrylff8aeki0CGJ7nLpaUw0Y52/MfXhw
zKeijeIbsi6mhjg/tIc1MwwRrAv6t3/lS5o8bc3yqiVbet1RivAqN0nx+ZCVMpr8HbkSOuK2LQvF
Nu9XTxAnUfXXKOi3n3JgYWYpbR+BMaJ5IRfaCr2Uh/2OBWgMS6uLfGSQmnKiJWMLRJnUgW8fLq1X
9C4hR5Dxxnj4ucpAG61ex/SE2WQQ+8AM1XIAKTlTFu0RLkagHl0NMSsj101JOblKWJC9zUlC8ya+
LzDbSnWz1lx00hjja0TPsOXUXnAU+FfeZMoxLl67i0wg2IVZ49JMvYw+s6yeTE743Y/WrE/P+zPE
IQ/oV6UCAEy1jt7H2ArBkruFoavsogVp+Kcmlel2AlKT58CZcn1uaFddewQne3/QsVzHiIJbSWUq
ZnWf+raDpvhcuwI4PBmczm0QGNlzoa3DxdEof9mAnGB9DwOSjxZ9ygn8x0ACrhkRWwKYGT4DfFHm
IdepHnJxREkQf1aRWW+0vDFHV7XN0j07mA9VVKGrAwmQyQFkDTo5W6NA/7/sL6w7iVgCOxX99wv4
XrM/nVaEN0KHMrRu3AFYWqrbHBNOqKOuY5WV8tWsSBCt2XxNjwzpdX/7PcXjR/TAbMTRdeu5Iay7
Aa/tvVgmDytVxPjEUEWK+mX8tf3eSFS2GIWpvLmzXmrdSxUeuviHk1sV/KCDT1/pbjtcCnJT6oDQ
LnwYfIV3+W/lb62KgGnsQ1f9pYnIIWna9RKpUCohFPVKaLAF8v3fM2yIng4nYFmeP6mNP+NQR3Hx
qFgQA2ZoD+lEufI07dZVcO8G3g8MeI3hPOY+/vHoKJwZjUb8AUFoRf19cjoTkL9+QJgvqt7dAWT7
Xi+covsvIiHZPfypb/op2Nk8G5g+BvPKzpf2OZ69q5m8N/ATtOll1aGrFXhl+PjYi3BzrGiEr9PB
+D6SEg6m1xepuBOUVawFMEQdOaKNMTj5Hc6c/Cd73B8QtXC6R1btSspJUBEY8aK137IZJl2/kjqg
fj3cucVf3D+1f4G6OB4zRjAcy3MAC923w1cugDuS3o0P9TPVpDSm21Po+jAo6HCsgkrwPC0b37BS
lst/3vjhzaop2dTBc/BGQnklDRe318A3kQGuSlFd6fk+BtEOULEwZ2IFDD/f/ajxqB1N6qIIUFMD
mKQsiBTvMrUYQRAITa8S1NGc8HAjG+3h0dzp9otJhAFlfcfXBXK8d7ELpw3urvIrA2A3TfdqJGnx
q1GZbsHICHAVpFIIcsxk/6s9Kh7AE3lzO58h/g37u7rEUo8WYmGedt3LOUxlSPG3wYvOKmi+4+BK
dWnt7jxqWz7UkLH0saaumPQrnJ058quM06hI1TYTIqZVgPHY0zxBqmuwF6qWJwyL6qgE9Q/KmAKk
qA+KqSCoMigGJt8YCbIZep0HLLy27wEL9PL5Ev9ppLVEvmYuR6nnv27IT4gg0Nf+npxLyTzR/0Rd
8/J5tVNyGe4sVX9tVKXebgI+44cvVT6hqCbKFDJF6SjEBb2mjEp+6NZlhdsaeOyp4qVVHBI/M0lR
EjxRevVPZ8rg6FhaatqiypHKLc5uLaJ3+Zi4Fwje7lK64eyKjpjYwwNygC9iOZESlSMCUZhX3vKq
0Wh4o0WbeOAAKa6KgOL8rHxn9U8x+DxeXlF69YMjnpfonfBGHUu64BLzHiTOR8qNws8JpIsigSH5
qPS87lLpz6UxjnA4Mr4NCgkQO18edyxOY+ezmgRfq0eu7U3tTgIwlGET3ap0kDjWIqiwawlFawMm
Vw6xO5FDdCLSxRhS16f0FAejTeHFHmUv0DuMzTAqrLsyTY+p7qVxq5YAIZnDO46rV9Z5voyvzudj
27uwTtQpQyq9Umbrl2U8p5UEE5AXve2CIobl9PA6lbAyy2VDPD7M1ymXx3gz7Pr1OMwgEsDgcYP1
bucL+DtgGcM4DK4v6fqWjwkVFxj5vr9UNZkQWWMbPWuuwh1d7YR9Pd9lYNJqxmRJUD90u8FPgbDJ
fH7VbFDtHZ8x+/P1/5iJBoe2u0u1lVXLkUXnicxUYLNBRCZ+VnXc5ZDOdmnwMClm6HA5ZzdV+6ZF
4KiZRcSVMP6htRpqcwfEVKZilzHZ/204nHOO9ZFgD5Ez2swBMozctUQ+TVi2bv2BwlaiZDv1RoM7
aqVTeYMFruVpFkO5A/TKbAPtmlugezXkF2JeSfcgE3iJr4keGNGqrNuooh7CEcAtv2dBZ9Ox2l0I
TGQczZFYZf60fMuAGfEgStoFnDWF3R37JhxqS5870FL87Z9MDs9KnEDYdDNFwNCg9CoyMFfqGAkI
XMhk8cKx1IBclPQiMWQHOeyf1mJhjWwS+FA0IhUnCjJB1ru8h4XuM2rVeEV15Cy7u2uNgywKTU6I
Acp584X+NxmlK0Hnb/L5n8v1OiVVq6V46xS3uljPkoSxR+rUCRpVnjVnEYBbtqnx4hn3FWza72lO
Km3/a/KFP/Wj7dZkWWskEJiHmEm4aTebwb74yZlVwoSspnKreWiiJ4AMhzN6C9xLtkxebZ0mz/au
TpMRgcopAbi2ZJWeFbfz9xncRTfzha8uHTnCeUw14m5ga6n3Ln6eE36dEXEsXVladGasyApHaxYF
mFIvZxmNO3GbwbWvDPBYZREz1KmitGsgq3POAP6nb0Os1B16OzvPcUY5a4E1KEI/tluIdKPxH0FS
U6mmqPq2V5jpWxZDZrhbJyiPOI09Khi7JrwCeUA7nRH9Q7qpa1d5/ROPEaANYhhs4/Du2nPpGw8H
UXugMlxaTg5kE8xLuQlc83rWIrBLIUy2OQcuBJGl6dgvSum7iwgFNLQat21GYl5S/NR+v7Sr/LBK
LDqnbGOVP629OQ6aGUQkNjbS+oXEP8vs8i2DFh0ZrT6cNrHZwzJJmvkXTsCe/qZxWQUTRO5Kcy5O
FTezGvMUzehreYwp3iu1K/JEflPgMTcli1XxPdxKbQdBuZtxSiZe0IAaikSu2YnVeq3Lx/6cJEI4
A2EcrFwjS7Ds68j8cWafDVuv26MDHi0LSSChC5gDCyKqZFqXivIG0nsRwjqe2nwGog8IRmRUMXXR
gkP6RfRTahkhb0vkDgrPtHZMG/5B6TlLgECfqSA2H87XcBTXrqI5kixXK6L1xRNGkmDV9HqRKDks
zKVWqoCXgnUSwdMY1pGiTxUBZM3EiDM30iLDCEWVJjjVYdgR3N3F0yZWWfbXHR+GIdsRnEbXh/us
Ps1BiNt7eOeXH/AndYWDe4yP4lmgQ+krMIbcmv0VWa26lmZ2tfMCLGkydtsHUWvZbyi/e+0xeT1K
HE4KCBGyyZUUT8udyhXAbQjap0OhU+v9qZY3UoqOP0BoTN/eq1cwA1eqr70vIWBPKFWpWKtlGpsy
fGKRUT/2iO2xcwhK5zM4VQ2tuTqDirf7wkU7RkDAP3akML0wlGQlTY1VKqhidP3O9xI5YMrHrxNO
A/UGa+8c7B9qP8n4phWkYoR+mQUj7SX3xKbOxQ0725UrgfsOcBVLg9Xaxr7HGgygDrznSZJ79m00
F+5IqdZR0mQkU0PBVw58P7zqIFcPYlUxyK3oqCTMLdrBgh6ZzrW49Vna3c08hw9axGbnXP9zO7oq
LWBpzASEMkD2z8lZRXzt0BzVMnQOp0z+ACjGi7w348UvAgYrs6IJ1AAp20X0KM0NeY9kVWgRU61q
zeYrNonmH1yKOYEltcjNFY/edLDhK1UONmQcNNZCYIahTAwjiewovqWnhnYMvjaEFHG8qkhegAd3
5t9RxVv0nyVF8mKPOuZi+LLLaQgtYEtWCDAN0sY2/5o5lwmqA6KG5PXP/dnk5En3eCDggB5RACX8
NaSHlwNFW+0KPpQ5w7aeSOd8qu1yYovGWGkCiBnVtTaYSMmk1rwzlFFFG/5welSROILm1auKXw/C
z5EppSCUDPprzLRoTouJ4KSxFLhGknqbvL2CqYRlo3tei1JHUIYciJ6p2FPpmqlLICW7D5eJFg/B
WvUTLbaEkn26v+livqsH5SWS1Tq75BTeFUnzLXAJ0BQC954BFXwzuSbWWU2AMhVwRQ4YI+RzDD6r
T7ydRt0dLjXr+IHpLmLBOQhrtk0H1ex8AtmfVm6dqUPArE7R+YyBfXQLOh7+SUl33SzpdYgFkd2K
dYroGZtjr5unBNhfoPlH9EjNZ2eV9j9JlGuE0UVYKp6zxjQGrnqjrXxhozI/YU6G5ZaRdeb6wvga
EbAF/s8bpUh4CYEGpTRGloVUdFOCK2O6/hcOgrfEdPeURV1yF9GUayc5eHIzOwtpYrCeVdV4DgRs
GVGvNNb0bZaqqV3qNP2hm7At32vRzoqGSMlYdZpFRAF4vy+hCeKPfqRQoJ5h+n31uVlpHkBwFmQg
80Ww7ECXyOHBwMs/VNglYP0eUiBZjH92N2x1ZFECyDozqzOjrlUMlypkyX1wC2Xq6dVhitZ8f3fP
i9sBjsVk1esWz9+aN/eb4VlRLE37yfLkN1QQA0hs2d/mBFchikiVPgklcSjqMHg017mG8uEHUOTV
a0qd8kDG3vag6AC3ZAXeEO7SNEFs51qoHaGmj+YoYKz6z6g1HMTNyLn4oZLQ6kXb7uEy93kXdk8i
98pn6TnHdw2bxpyQG8cV6pEVCeShySi0dnZv8PGtCY+e1kY+wfzh7A4EjxNW04mYWYEPc/JYe353
nz9y5EeBCaCC/vJ3zcYj68lNZmqIEYtMrpNWNV9Y6kfMozbZjQldq9SoXT2zmwTOFKRS0Z2dJXVV
VwiKW+pfI3hcVY6TMNoca9E8eKpZ/PlPTxs3VZLqalU34PUAqH3mRVqyBbx+i+Hujs8Rg7z7DXJ+
jZ2kV49V49VuUVOQtUCqNxvKXTlcWlxem+U4UhF0ydav/ZldIHAEotLdYxrS+tj8g5ft+pW1A+LB
IVCxH5JYSUfE9i9+/Jo+n5t3TAnDqnuJ8SystIOjdY51WmsRbO75om1S8bhyO4A3R167PXdfS2PV
Fx2bNDjlLX6oxDfEXzVg25QJgojlJt5+MoTaBnmYHyv0yYyf0tvSJkj3EEe027Os7RaVCs8mnkdn
HVE28qx/0O5LvhwuK2mb+5Bp6AhpaljGCEFXo5cO4JgXnL6iP63PQ/dKj35D1zgLBGz3CyHBOXWS
S5Mt2Ca6iQe6wZHCoqZI4BbJgi/m6G0HtYvydcE6BVGbxiBG4ZaYoY5F3E9+ZEZZdIpwNUOCfPKp
XLJvE0AjrowdQvadxDk57jxxVDBlS0wfbCH2zE1838CGAERhSAfXaYBMcsUig8FvvQ5/GkR2iEjw
Z1WNkhVP6ZHa/ReXU/JCh9TOsT924kKg2J6eIhl4J4sL5aL2XjEDAtCVLPvGn1dkFdbHVqdsjr8D
vHRRWvKqCtigj/5b5UTVOO77FVfClcB8Y5L0VNkgSwIr/hG6RJ9otDaiQnUTaKbdaBwM+NZFOXnA
AEFJiYVF8kLIRVDlI9tXD6ow+WrQkE1f0AW5xZUL4UDK9agGc575chjmN0t8opxjbaHqKoXkFZYI
47aGvKT0UElSZP/g3IXYr2NB7VqG0n7mHG1RadB3eAOvPN3LceUwat4HD6oKcXFknuIKEdlXSqKo
xEFD3AJ3sSTfE552zDS+7jjQMyLHsgXf5sqdoyDLmZWiUiVOjfjgm5i9J5p8f0oQcCYWtimVnDb/
xAZccg+MKW8tCwZy1oBcbCJEaXjvh6+2rsC4+SQLOTvuOvZIyV9TS1x4DJtSc0Ec8SglVTXutBZX
HX4hE2BFgpkgIAZvIWWFzKB/Tg98Tl8BvmXJLtfDVvrpzUnlLUABL1J6x2RTlp9p2FrPnj+pntt9
KH8jUHbJKn6fhwWAo2zwxytH+LYkyzyRv3gY0A4rlc1go46DLZLrJ4GuqnECGunANO0ygYhmyAYD
UbGAaJB8II8UBg5cj209rof+bxA5B+72xjYJm8HjU00Rc9/k25IJJvbiAOxGLM5UoLdA6r+y8ljV
L4oNSlbUs/5v/eVbo5Hl04zgfM5lXuvGV7vfeHxqb0S3i1tGDEtwKncuZzusGTKfpodtCM6r4jTq
xZHeQFtg9vOB3zps7u5mcv7A3RrMxqDdG5vgqCEioNW/EH/BkcKliJVKP9oJHSQBNlWRHzLpe2o1
E9L4GKUaw+H1mrTdhdjNgrBsIipcV3HphUTpwroI8dupsb1CTV7NheGYmzlSav9dGLVLcqwZ/rtN
x1vrajFP3fiSxLD5QrGx7EfMugthVqo9Mh4pMZumTqGCPmmhd7XpkVXhdCgI8Vvr5B0jNtXI2HID
ZwQvNDjsbp72mLaM503ebM0SpyF5nk/sNlS/GgoXoMokhf+7kEPsfTQnTY1PDQLdiPndmPGUYdg/
x9TF7r4QNwcHQxQtRfry2WZHafrBs48m7xcPD90FLvPRhOASrhVwFJZCEB4bWHdo0PuGgM8uj4L9
MH706vDRuq7Jqmkl0SX9Dy7k4VaOBge9KpfsBAlA3qmc9auUI0J+1/x1PbIkH7YcjrVf2sRubBVG
bG8adiVbERJAc0dzFM+PQ+Gij6IbuywOB6gobfXYIsVz+oVSq7N1OILQGbk4XMnDtidxW3oKjbyd
Hmt/KLJt9E3HuLkc8ko9dgG9Meh0wAmHTlwwwk37sMgH7E/sfWPlzVYTn/Io38HKLC0Xh+XPy4Fz
hdA5ctn7ipsYM/2osbieGDeUmDtTh8soc0XlttBLYAKp+obaIKaH9TKrdIjRch4Ly4gVYakM2MZk
XHF+pTEWNToHjRjBfxs1G34mCXN/Z2eryswPPBaeU0O6RGzzMcBEBM2dcZKamxIkm7jnxVO7LOdt
lPluzSpZ6uJ07Jk6oSx4oXMAAo5kaatbZqkzJIYCkTAq9C5PjTAMn4mHmBEp0L9CdHJKDCTABCfU
n9sUsJIZJTaf/MRXSMJoT0YFPTT8I7SPUZ0x4mzhZCAqLWoO/jBsP2qjSDMVvVZPe7ZDGjphryTu
XWSm+DYxPxnn6bF05kp2jvmJ1tCNpXF5Lw6SXvcsqm1CeA/5+0ibOn6M60k9DGuLJdj7QMUvtVms
yAqe+046c1OPWuocC/4hoGPbyurtcFlqW8gU4SK5DKR3VAaRj4bT/iVs8fhoOcPyahgGXLUXYIsL
RPWQ+/Sw31EhrJeHOAAWKsQU+qdHQq/xWROs+o1hEMGfSInRZSfDsu8yeCN7oOfeSUJFZlY+6khi
wymznawwsJeWgl56JmeHJFzKgLrAlDBP+tTqmKDI6EicDACrh+QVFHlugfhp+W6R0GMAHJQPvgTQ
/dOxb/1AMdyugc3W9wiBJ/7FoTx9xZGb59ikZfqji/Oc3IlPGTrds+ogcSmI9bwnQDf+kvY4ORTF
N1b4zBN7ALFukafX/FoDp60Zs8VW6+IyK/qvonrrGaY2bzATBCNz8RaPjw8xId2vlUwqWR9vqwpF
zSaWnadnSKpY6rwyLPFdDYnPFoiQPUoWTdIhR5hVQEZsseJE1u7sz4n3EkRcLAmD1YotfAHDDGt6
4O80yj4urlbTIHsOiTwr56EiNToFNbvzvbqoIHoRbDlKkfzTVrB+ogSD/t9byDxEWFrc4Kqrhxt3
rG9dGaRr0pAIlwmb1wJyVwZUkwVkhihmsGo/pnYuI0NsQ/g9DWOdf8P4yQf8/n1JZKzZyvt6Mcwa
X6cWtmKrgx/uAauv2mdri9Iv1/7WNHah5UEZcwu2D/vlO/rtITc8g91e6/4PxmlPi/65HDe/oW45
inQbx3i/o1YUQoKakVC2AZYIWpETbnjsEvk2y4aUcF7RHs8CXsLY64LBI3UcdJiZxc7EInJV5m5d
d/OY3jwEXiujkJWkanpZjl5uyZiSdoF0g/u4lvvMCupc3Sx74vc5b1lVMRPM1JppRxTLQxDz327s
jPw7SAgLXc40LSc9uqGPg8wcQX7VMb8aqL1uJLjFHp7EkNEdznaV9ldIA+xkfsdq7VennEg7YUsy
vvqbU6cbEcC6PVtJIshQFrRgbRmvQ7wqWv0ws83E9QMaCYZFTlyG5LsUePDmmKq9Nwo1FvMPtaxi
5SWmxfU5vrZv6h3tsp7KGHCpNFHX5ji9ShGa+TpkxPo/S8dLc747EHpKgDma60ea20DHvNhCKdLV
xv8KGvw1Lj7S50ulrWBjHZhy5jtdV47zmFw3+KA0/ih3K9MoZOIF2+WiGYHH1biyz1+QA3JeMaW1
UbqOUad/JSC987dmlBP4h/qPSYNT8OneotTujguJOhUO3gnvNg04JAAgbxwcdBV/3S0YunBcRFVj
LvLA03oRNx6xGUUqq4Stg25lH371emHumXQn/n59GUS0F2Ji+D+m1OfRrxw9Z1I3Pf0+vFlLP9By
RHljKk3Q2h8qutzqUlfySrf8f0+ZKqVWc/hKAbBk+XcpZ2DAUrNylQYZx41Jx8CLcdEhvew3jNKP
SdFQn0WPh8cau6pm8TJxYuqy/JBH2McQ4yoRXfJdVXd8jPGwgETr2tOivecidYKdrxq+llWeZitC
3PavnUsPL8+IqykuaeZwcVfzLOYszmVUAt8RDbwut7E/h72WelABEDeTIkP18FwqiacjA+gx1Udi
6gRXCFV+RAXN3MTeLNpep873ozUtNW6Nyq9B6BHVZOYFAmb1+/UIj1otSDR/x0rymQXd/CN4EI+8
nMKgQp0nI/66v8A9u0nyj7wi3LQPj+Irw6hKSypzgFo9ZUjJsIH3RS968RW4c308ytyrSdnQdvUJ
dsWjHkemCjzNTuuwBPmisVbTJBO6OiK3H6l8PqI1aRv2G53hTreIAXxxscQDiQJmqLQNwM/KY9bb
sW6k2kkLqgynZsVGoJiUkuS/kkZwBUFYzwWyEVFucAT563OBL6vcAlbftaGm9OK4AAH3SIzhY+8o
4DZSI+GZdHKURfNfvZXJ60QtTVsy6GyV16WJLkf8jFGPwgvDjwJb1KcLawXgYf2xU/nONe7XTP0C
P0VoHML7IEmZkNOcaQCQ/cp2F/NvlC2VfzASI7JCGonJ7ogr96IoBGLiDIL1FbfPe2wCWDQtdnqg
jP/Fd8FqbUf8mrZbeyqrNj4GYAMUAYBCoeU2VV9hXlC/IQ5vq4X47ftVZ72dl+8TBZrW4quIhOsy
noxi/1jEB+IwNgxCVke9U+JyyTpJMzYdelEXjwR1/t6S8G7u/Jvme2Eg3C+qvuc0a/frgypHXwFW
mmfGfEP203tuE1iEDAXCXrecTD0+owk1PsNjokv0wkpwYp87AdPMhBnrcnBP86B6PC5oWF8T9ycz
ucT3KLVNQjEh69iHPwHBPWzwb9Ggk1qGDccfF98JZxZsUoxEr/S4osWtsR9BTrUOeSRUQNLOwDam
MYDGokTf46S6cAF+AsauSnnKkWO4iVg3SBcrfQ1gBgwjrFyvGKHpZlvFU/n3Rt0VUcqavBQIP8pN
mhtZLlwHQ5YQ2qkAQ4Y4QEjGT8lZXe9Quw9J4uT3QQgElq/faLe2/i6T8BPy/nPJMC8Ghw7NSjlP
WOLZzEqoroDvTcRsVsIakBm0e+aFXtzWobEPQ/p5QoXAS7bkH+6SvP1QE+gPxTqzZTe3VgXugEJC
t7YBpsp6MNuxFM4dTcPTC8pa4/RS0fxj/0Q5irbqx7c9RqDpxBSaAE0x3RwTyZLqUW0BfJmsgKhH
QE8awdiwv0O0FALC6u8S5gjbjACWRE1MKrJ9crC0qvkreweCWGW64dyJjet8wO7uzaZd8XQBZxJy
IJIkyXhfN8kYq/6Z+sI1KsAT6Y0yAEYW+ndxEwWHtTRtQXh06cLh3kXJm0U2jkeGfVkAimQGUG1Q
H0wri+Gwr6XZ3k001IJbDXiYkbdzNqgH0q+kpGJO5JOjL8cCCj+HdErIhVbynZg56aiwssCfXJKy
gvvb0Cf0FjN8BYDOd+z5Z8rJoFlZn6X68vCsQlVteEVpfYpuw8Hht9QX2kbc0sy+i9uzh6iAdTsP
MlcK3Bzg6EPKRmtL84d35BprXrvTUXTVODO7yu6CoaqjDeb3qC7D4C08bZfM1IDQFPd7d2w4Nnkb
UpoWEHABJBUFntfjIY7IluH5lajf9X8oFD0k2qNoWKYVhQyK7vLTagT6IRi3dx2KpPz1QWRkzjiI
ZjpPKMI4LdCz3l/MZ8vkwo6zxHJc7BgJcEhmiPD1LndM3PBdkWRWhGQCDeViMsZHUxCQmmi38zCD
twQ5Bdp1YlNB3ntg/SxWkbo2iL26iOcZsFD1iG6WLa+hxHl7pC9+CpO8LdcZMSfGlxLUWej53C3N
N2jAouDSdItp3v8RPh2bvgrF7sDZjlFej8DhppMHj6Q6K/J4qkb3Sff0UKUB45tLwVQFPh8J/Rq/
R3U0z49Ee+yhkxXF0u+BIVYPeYGOVXtlZ8mWKg5A2/MU8MavcgZJXKXgPOHQ132fKtXKWHE8BHQP
OyewEFAO62YKsF50hy0pZngVTtz0Mix72QO0yu0KeW/l8jXOLUTCVBVk4db4LAvGQ7pbbDIUKsLT
K83qPhgXB1nkbMde4so4bjqii18DZs2ARhNPi2DYFKLYlvNNrzFzgwH6fivHvs+Ss20PoRtM+vzQ
EyTsqdcofrvFt+dajtJss0pVV5lcbaozD98KVNuiTYeypLZ5CvVpctSWdJxY2lZ+3Avdmw+x63Ll
KCIvb3bqxWVpigDN9ajR4hMbC3LIaYOiSnBMSdkqxXu7FpHb2q+QcqBob5KqHvZaDbaDfjkXYG+y
OnsvBSxhK96IAakAEGQtDp69hcyM0G31qOi0VepTOG7Dl4kQvDhoBRKaH/J6vozj23fIFtJPFWdy
5C5Nfayne0ArPwektusv/9b84acnxI2jFk/s87nzhdkmRmqCIGy2PkHUczog1fEgMB2YIkz6JG1I
0WLXwNGOTKEP1N6hdlA9DjdAJ7zw1mQDEO80AmlVMRJP/WliiSP6WayA3gmo/Y6LrlM3jlVuE+jR
bBX2lWMBWYnVCLBvMNdCjDKWN7xPrlH12HD6GJtzLtMZXr3z7r+LU9lJQAQIosMQovU/gsdRfHA6
SUSvLBNSBYvvPQRe65H6zH8enqqGaztWTCVLIgIWg3D0ehy5rItE5qeC+y5rObvKp10qr60EWQwO
OQr/7tBTHQdt0gSDaz20mEDBuAntJYpDMmCX2BAz6oq3rSVis473uMUN2qIMNzIyLC7zgdEqrFBg
b4f6qna8ZWiZtTvyKJ7qRUpSifi0KitXGGSCOkR7f+6qMca+TTKK9/+bYTCl/k5nEb2hl5pqf3j/
FpTv+mLluWWevSAc13bZ80nRaNFDCz7amZJ09qXP0iR2w/AAsFBwncPOYfmE06UAxcPZe4pbI7TO
HV9ONopAP3tztsbxaR/tEtniRz1O69MGAZcVPZRCEyvs0eU5H1/VYU+DZdI5mBlbGZz7Z1/dbfBB
QtHYRwCSIOZr9CySvM1Pp1uZplM0i9Q0OYkGBi2jB2ST0Sfgq56Crq4QI2OIkDGnJXjUH1msCLDV
aVN5g3L2f0l1lvwvPGR5jSXLOmYPck+KR9kKhdv/nSTUl4jXt9A+GQg2EeZUWRJjtlGSuQFFUR/b
/ouPIDdyf66P//HcoT5YoTeD2YThYfL1DPtF7VKwM23gSK0jZ2X53STrBXI7fXaskbCmv90fQTfO
SSqTRI0wSXJBvJUU9sopMuXFJa2aE/hjqdazZcRlAaznPKa+vBU2iTNxiH3mKMQ304PH0k1x3YVF
wi5UOIJqUvwCWqNA2w9ibjymIM3ZtAEVozRQxI9R86R2gZhpb7Z3uGDYxrp/9/n+8Y/GdaIWnPsE
xnlIl9u2ZHlKkeERdKmt22G4X+RwFTwOA1mC4B6PH741gGxu8v3j5w00oHeZqj3pbznQqBLqEmi+
a3kXuwIfKoLk5+NDtBQ5W0GXQwZ1TAW55BmBdkqsKKOS8STCf+/4aoOF1FRYiOGV7E0anxgGS/3/
gB+76NTFlAZGCm9bhgwLDFGz1QPXcLlG4wy9DUwFMU4FEw1fHvw4hJO53J189jyp8pelvT9K5cPc
Gx/rUOeuFrOSGYo2ofwL3H75SLd+gYSuTpiPkES3eqeNv0yGgDk75sPNmhaKf/+k/sb72uEhirSb
1wsz4sEWG8+fSPUDOQB6HnIwBpFw1tjcRbvTjng8D9yRFi1mWcxCql6r26ipr3b983djOG0jgQHY
zO2BmoZhSDQghpKICKsqK3gWugJynLhM5TnIUgGSFOAU9Q4fZ3A804ruJmBFhT4DfGvg2WU8Drix
pU9A0xKG/tCnJDJr8kQBUfqfKmnhwY/rygq+FAKME7bYMqHihenzZ+4NkwMcgJiCl5TPbQBrnDXo
BTa1r1Yh5y+PLTiOMR3xTDYDPHzC4X4O3D/q5vZr9L63EAqHAn3RRUP8Lj6Tm4KZKWmrplDcItK9
pn61JQnV+7pM216oiZTnsva2fLY0Zr8zT7cpUx2QKdgT7x+3zXYz0mMlaf7KDFCJvKmmdkWkYc+z
L/iHw9D4TWPH4c7pXpHI5w2qNaJ8vD4+tVYqKC/M2J6OaHIcZY1U+m4RFdEt3HDyaRdgATdEUrra
p5HqOhe3rxzG2id+BFDkKtCOU4E7c0URc0Xnvwmf6ZB+gfDHYG/j3VDygDf75aNTqpx0UsvXYzQ4
ZnYvMyFlkTQEArA53vGJG8VCwXZQVQ+ofXVAPuGeEGlYEmArKYZlnUDkIDQtswxHOohwYyw2h+j2
zt8M1BcZzcOBVVvTNmO26jf5DPNH7VG2YQ8ti2/gSMVgC/KUsCQ71/5cJ4YC1yZXTGJuxXxD/bzS
34ud9Cy3D04VlzucWjM6qELMEaMZwMbeM8aAN7DRKF3uPTzkHHroKNg43P2UneOzYiDVjpVPRSvw
VqVxbMcB/AcLU5jIUKzn7j8lwrwgsIY/WTSZ72w1YOzI2iB1p6TDQLLF+0Rrnu8McgHUmhyA0HK4
F9dkeKo/bmGMFDNcQr6XOrGNZHhJFHPKMYujnoKotX+D5eWWsvzSzAtAaZk+UrFaUH/sZ4q3wE0a
XtQjp2JqW70JhQgeyd8jpfLIw4Aaa2lVPfbrvxqDAri8icpiLBTzP6lo+pvfiqUD0Rk5SaNvAiIu
+sS+X69eqDNto5Xmv4tl3twqSXxe56Jd4RiJwrnCrqeLsaCAgiWEJSilP6G9HEXQcyzHuTVaJMr8
uBHeEQXJXJyDqoCKH3wIL7pkA7FO/FqEq9dcxWd/xAv+YbR9TqjPbqsMTkBoCi5QxIywUyokm++k
5T5dM6CQ+yYMrD5CffCXiMqY6rycG/u/o+fbOXy+mom3mQk9tWh5saxCrT4MfKP0FZyLlsq4TRwE
QoCiFErsx7j5PDB3/rqC2oUElO6w/Mg9cZC41LGVGin9HcAamJDUPgEuxixK0VQ5GfW7ESYn1DlG
koO3MQmSVWD5GMJW7nQbTlhjsBSVt/4cyFqxG+Gbjnxg5xwqqknWP9cmJFzqvQSvnAUYNZ1cgJiw
2rNr2C6UFPO38Iw9evS5GwuItkMCeceq9b2LN40JLI4AszAkLb1Vez6fjJbZpGPuFlNU2GwfLdjn
4Zib+7rTpiDGcuphi79fVWv2Y6l4xQR3G0wBwQe7Sgl6XVq6bMVomJXaFXtYQJKmzNPAmHFAwmW2
JIqtvd6kfy27Fw7i5cs00QyeOE1xI8VEw84pYFGr5rvdVYSQOXnelWoS5uOT0zvmdGCDDDOENK4d
wpo7JASg0YYJybYq6yIR0esmJxNEVPeenyVEZZmotaZl63o3H8PvdzHDofVzC1Be+K3k2Z9iN8Sa
KMAHwnFtX4k14Uj8lydfVx/mNt97ECrKGxDPlDvIYAoS8ZRfRHZTRFxVen35S1ph7LB7eW6ByjJg
pq4H7jAKG8J09lG5kTEyyBSiPRsTZAsE+XaCrub/pPwRmhv4V9SlnFXtBbpO9xGZnSIaGHGMYwZy
4QRdWAjbpmFl46BZa24TY80xN/vwQ9tUrdrrYwG+G8ZGV01M5goF7PYJ/T1rW/NdIcf44gQ58BwV
BbTj0h8w3Cwq+AU5K85QLTGiOWcc7l2J6cNyN1ELzRbixuVLjBhvndYaWMm2GpJmZiufaDVU/EXu
xIG1z9kMeMNt98HJ7kZfp9nndXDtnct3IJvX8jHri3qdXfddceqyjrObmh1fpG/bzfVHZ2ncQRWo
KbwceFzLzmQHE//J8VwDmr++vaURcdyF+JalopypmJP/m/yxYeXV5Ne7KX2vARLI/IXjcZX0Xg3h
+UpRXh31Ke38Ik9UYer1a7HN/ozcBpqKygk+qOLEnbmxfzruapI4zabJUVR9vG1t8U++YEt1wj1y
O9uF0P87rZSFCQHP1Zf96dgJksq9F1+sVtheee1y8DL1oEpQpNQ+M/z6RkX0D2eEaAMyE9PONZ/A
wFUVl7m6kd8B3e/GaZIy2rh6RGxTYEOk7wnf/VxbMncThmzFtkd0+SDk/5CAu2jd8LfUXY6Pkgve
W1pfbgPNsvQdG9p8/c/4IwGRXJxM/Tq3B7YiVx8qHuyMEqMKOqsZmsCZPnjYBAtrCJuWrA39qleP
uMcuwQN5tPVp2qJu1R53dJ/3aNSSzIXr2tk0RKojjZ/qBcaZqG/drMxuvl90r5c2TYh7S76E/D3M
rfMNo6B6MAgy7bVj1epWBhLQdQC6PUeTnFjzDgakh/yx4sris6zFP3KT35FquFaTYAWqTY8PFLOd
6sXSVFL4AZzATdrnMj4RQlMWWAYo4ijhGlhA96SkUR2HOgUk8Yc6QNihlf9npWspcODygAy5sbFc
qgkCro3dCfcu010epK2vCze73q+KZT38SffRS0quFmAGnHK7tOFB5/gsG7BoVW1cg9n1VJJw3/K+
/PBJfeN/Iz9ToUITKyoABfzOuyH6ZR3WAsp7UQk6o69kEBIZ+QZvQdLrCazbg55DU+TKNTrF1hUm
fA6/ZNOJtjHz9+ne6DJ4piWiqspq+hCuY9S8ytV77NKtMUf9RpjRPbw2VRWxUfJBCyM+FBSatQSH
qESjPGOFz45PuXDHDFP7bCGoqGA060iZFZleIZMZ8KWeJc8/GEJcdDYZ2M3Vqy4EWimUIDKOtk+w
OukllONzXY2TqYmWgnxDZouLyteGy+qnKgwFj5dvbuNZuQLvR26qjmvDfiNdIjnQdnQZF9BjGeFP
p8vKv+KghaigiPYmjQITgA6HCgCgdtGvStAmYoNlLfgjXacGTkd076Nk9Yp8cfWIr/4DdV77fNM/
9QedDEmxuJF036W0h5yZSJPcksd+bTkRLsdQ3g2FwioGm8klDlBdpso7LYjDlKBfdljkn8ihu5kg
MksCtpkA48ERpbXFCoFJNDltkk0BaH7S+YfzKAA7ZiCdwV/i/namx7u48Is4Q2U21qT4NTan0OWo
CA1KiHP8BE7rl41olshRG9iMO9x9s4uoVUtt1vE3/2IyP2cKFd/4cHo4XPXqNSkb9/E3z9CcNtnL
cGMmQ94d1lNoyZfMlCB4AkhOhj90sMGSTTAJjaFvlSszbX2qAOV+UzkCVKYWH7MDhDN5qDVy+Bk5
Zz68Ph7LdRgJtnKS6N6ER3xbv+Yz3z2iuGdRKDEIw84lLjeZ7TDMNMzPrZtzosN+3vp3ZhHhmK6z
C24mKx9HmopcWubIF5rqv1sv6dVVih3oes+8K6dSHO6f+E6Nv/Z9Tb+pblpvopY4nywAyKWntGWB
GReXH2UWmoenOcsbJJG7u555O/m8hjcaXyeMeLCA5lUyhSKTJ7fOfNb+KYxiH2gb3nzS9Vs7s4x+
JrLY2A5lcjHBBXRIxcjBwSpfH6BIOLS2vUzYNcoKio+hKwIm8dntbsH+SzD4DQiQS08GlLNj6aNV
+WwVosSeY5pfQG0aKVLV9rFGnUCoLkrWguCBogZrxHQ0H4Xr1+O7qM5yXXr2tTQ5lU00tFehhpu+
JJZRTZWPfbS0WM+qoJhay4nX8Ov43Fc8T+TKCveUexBu7ltxwt3/pkWTLdnwDivBN1EkMMONBU/X
P6YWwAgsM/sC/m7O4didqYV+DwoDddn3WT6WR3viBIeE8Gn8rNskYXc0fMzfWHpLCbV1wQo4NvIm
PNWVnf5xSvNkGhPNTNRRcsXWLFU/nEXv6jQNT8nAX+5fjQ/ILtP7WGwQuer4vc5rVWkSxO+g+Aua
/1Q4Fwcx2jNaS6cIZcbLefgODnrWsOZTjCx/tY2pPWwHHNlTAb3FgVJ3mtQ9pYRLI7eos/WLwysF
RDCaaaT7amikJAslBkH1D8UDLC3CQvzohWa8ZM67ATW1y0jvXg3n9r6ZMv1v54vdfeqeISilISzt
ccKZS+MdNpFwU7/d0Zgbh/Jm+mSiq4vMauHJP+SsVbrwBqYiJt5z+ifL7sMW1J4dMF8xakw=
`pragma protect end_protected
