/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvl8/pe97suua66uGxJvKMsBk8px5Ly1PbBsW3TM5Ur+5Sh8zC8FxmIrz8
bpM/AxDLfUaVHrSOu0lYVglVr5wAaxSw19nQvMomszw+fORV92hKGRaH3h1W0VKPMk0cqu+5TIoX
InJ6rA7Z7Dw5OtCWcGGFCfBAhlsTue2wp7b8xPZecgVsYG2fZ+lWcHoCdLL6SnzmghyL2m0c+O7A
t6DyUup/UtPebZoDMEAERECNtHdNAWo5WRCKuSrhbBBZikMiibnq0rYqC9Zd6cVtt75s9ZZT4mD3
BvOzRtAQ3nkH/u3ZXqmKC4KfRwPdLrpY4Aq1biaICTfhiEnqb+9b9RR4+IM1bS3hUqT5NZBXCcDw
kcZOky6V2LHyJkdlupWMcUyZHpjLEUF1RTRJ/VAhC3TSdq/FvA2o77/1UyXm+fyxbRAf/n7Pgf6Q
s4cxRrRCriUKQ/AegrFp9cw8k+fpIxO0cP/a/Nzk8wys18mvUIi6EUIB3Il/za3cbZYZKvfBVi4h
IH8ujr/Q8tCWsu/+7ldmdp92fIEiFBRV8Z+7EgqvCldMuLxqPP/7QY+MGQBjLOUf/qA1YE4dMdj/
dYAvEuJo81F9LcIC/YitBjeyA6Pd1cn2QkolFwrJGPioBBLUpPGYs9pGSxoIRDXVZMbXZ1m1pNER
PaCARlvuKAploFA7lZpvVGEeeLCEOHqyOAh6XThZkGKQIEaq3ul4dL4INcAvTtJM48/uPl0P3qoi
nqxADNSIfJwNvZ/4sPoVmofWUhXVIELSCyl3JjNPF5Q1Q9isTAXKU4LO57qjPwYt8HjW77bnLFwt
JElOtogEvXsY2dh7PlqF/wjSpWawO7y2UcLQeK6eYGVQq+CVh/KmfR1gqsDdkIlP7LT7gMCPiRUp
+b2baRjOSL+sVtJKycrqnWUEcJ50TNsaIcl6vp27O5egqn1cvHQuuMupmW/QY9Kn46hec6c+Gkyt
em8vo5CCMz31dXTJOHCIHNwUwwULDouF2qhGgGp/OMlehjiWckrTSLDUGakP3xPg9OzPk537iDnF
ndkviiKRloP87ysQ48fkHALm6YD+ATi+T7lXHNgLWAg+kRLkcupkGOjNfpNpy11dZoi1eLDSMKfB
DTwbuqm9fRS9eE3OvQpqjPgY+ztdQAZ4T37IY/x+t9veoVXHB8bB8QFB+/fRt+zxxSP65kCnfn6t
nfG5io3Bhg18pH4+1c7kr/AlN6cKMJ5HbSnMvKMpPuK0Ne6aL4CfIp9a5sp0r72Ehw2Q3xzZrFvp
xO6v2JEV1nb/RDYPnrj2PtyrRZ286mGSKnOCehj0kV0w3ctlfAZCucROpLl/m7LoL1n34gZa7g5V
I3Tt7AgMUSn/2NBqFNrJmnzswyQjzUjZ4Y8y06R1D7uCqt9Cp0MNgClDZMVMtiES7Nh3848seN9E
sPYD+LEVcolJnlH6cSebeyBs0Je7HIQkZRZGryxHiSefBEctzGrrpVOyfo8lewJeOWhWoIWT4C2U
CzgAVaiU+AyaXbUAMat0hMaSiLDWA0rBVpBmGr8vHgD1c0eAr60HhVWBrTTHrKA0Mq/4rv+syBcR
YTWYiUFfqcwz/3eoFL47Wukb9TdgQ4tg4e7jOCRXH7AeP+C+1RSnVhmomlzQKPDq/fHatgw956M0
JZwF+3AFaCN4nsOzasU78idj3bO3VlqvNDxSZGTe0gXru7dKb/oQhsKIk6MuS0Wm5XZJ/yQICTtq
TzR5KlzFj6vZjFH+jy9Ijr/8wgoMafcUKK33iNw4WjTTligiv1Nytd+PKICn0VvC/twY8a16dxFQ
D+ZChZaI7drWl3uaZViB4cBuLYn26Ul3nWH9oAXlQVeWn3u0nU6j7q+AWP17Ed5yuDG48SGVHIdN
uuq9GLgb1S7uVTCtE9vf9nNnS64VGux4hsBgrsDuqAKBso7UAj04n5UFr69D8mbrTN3p/idcdb7d
rlJ6Och7XMbmynrLYMuc4ay0j+Otps1MHMt+wKVmTI6eWEwpEczG6AGl3+4A76PtzcKqikYB2gjj
++uB+0YqHUFd5Bmnbgq6Q2NWC8E0h1JqV5tykfKAEcf3ceOrumyntPbP6m7YC7068JzUEp7dCb9k
H+emMR9us/QsuXyI51pgaQGRz64F5kLA9iciwuXZ8InnecfVuj1v+ZJXyiCEI4noZECKYoPAx0BE
jFO6kn+i+ESypFet2RDzmEVeb0if+cG3T0RanXRO0VTDr1TfR+jlWo94yWETX/CXlpCNgD7gPp8z
EdVXefH2mdOsY6WeLuCMAzv92Z2um+LmiVnp/7VO7ml+QQuWjY23pUCOoAEJpGE5Wc2Ksmmczuij
y6UuIwbMliG/iTyRhkORtalqC6ririw/B0ebm33UR17lz2VjzfY4RWPMeKxsDnxbcwVEh9y14Jh5
NIOMgnharxpE+INxANmaXbDzbN/Uk4NayOhX8ILqQrx6ukDjj6pcD3jiugpz7XYGiu4QB7PW1Dcc
r47LQXqXuHjA+8ykDMOUpNr9K8SeFNs7UWH0/faRsm1BuNCDVRMorVRekENINQDDVxvcR7qJXkt8
ghXkOveBY7Q9czWBqHaHS2/gjg8WzeuKKCcaTxg928OUlAXYHIxYBNT7xYsSfie7s/E+LY+SZFcj
1I3EwC74t5nyFfIasusD6uN826tSFrWPpkQm+IaaI496EI+0fMEerOQ9+pTmYrf/lGQfEVKGmwln
GNXtOo2+Dk33uKVFpi5N7UH94msIYfj4Fcatgy0IEre9NuodN/fJUSc8sRV8zVVPTDI51Liys+4R
kDFHjZEL08fqaXFQ4Mwa51anKi5WhKgWhskCjcfMVvqlCFadgSGYOXS7uRUEYgqTmF4i7yYPUjrN
w9wUTOjqn6Omn5dQyID9tnM2lTZV+wpghHI9hx/aMxuYJinZ7mu2iwZ2TBa1+pwUBb2n58Wf5EkH
Cg7cNpnY971WSwZ5vnzUtECiEz79tX2dnTUOEqw0DFc8X3D+51aqCOAonKMJ66ajl0Q+ARupBXIX
w5FNTQgyinLrPho2Fg/cfIoV3LoM/vpmeEnhdvl2iIJYIhf3Ag0Fcd8c9NZtG3KZQaDw88gloRaP
SlYg3Vx3aMQNwJWRaelg
`pragma protect end_protected

// 
