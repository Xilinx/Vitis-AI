`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdFxRDy7LOPb/1kGDW055V2dEBLGWTRbWOSlQlxcbvKoKNuZod0Wn8fYEh
JjdRGlUxdBz6/b5rYk8PB43c9CEK1l4Oo8PD5+FOAB/QPLkxyHsIpCaF+Q5t1FCKkYbu4uFOve2o
XFFgvkIxFlciphLEk7Tq5p5gcJJtkSfaJJAjw5g37btSYXvcNqe+8oMsHGiTEbVNVVjA3Dj28Igh
wpwAjtulCd5mAHHE0pOHoGYpOSsJ8IRgc1OzpeoXnWfVCbK7TqussdLoCgQKp49OS2v+wQDu7G+K
w3DP1FdnsLqMpEeFcT8qrYn/qgNrawBkMzq+mRyjsg21THR49ACCCjZTgaztjQSu1+dZxmipMyJA
i/xWjdxaQdobOwx600v+/G14gKsrxHtxiLUqestRpAHddfbDW5S3MikcorQhxmMbbi4M3Lqnp9m6
fziiwi7kRUftl8lWueq6aG599JrEX51aRpyhMAvYifZ3kHwECvql/TVry1XcXpSjakdUb1zUKszZ
MRDwUQAIk1DBrYdbH5iaV9r9c9g01X0tKPieLeinxWN9b5C3AsebDtRaiOokThqTKg/m41J8V0oP
lyVONjFdiRTkBdvb4r+/I/ar8s7wV5mCnmTCnHIwMBJaJzwSDbVyZLYJz5WbGQNDgsMp5gguB9xb
Y8ENu+nCvLF8TjLA/zZsqpSZ2ctHzBDxuIyl63ecoGC61U+Q7yqw9fXFwwf6gSXzuLxHUG2rFmiu
eHChliR/PPymJmAnKbXylUiyT6D6REWxg5tFTBH158MD5mO7GXDW6D/UNLdLy9aelzQyoB63U5Me
S9y+n/ny26NjdpG+K3lyQQzShc/+/OJCLQmw32s45M/nl7m/5EI7CnYxfqK16Yw6xzp4O+wVlVan
5aD7aXv7Pct94vRHHQvD7g1QzMTXbd3tXHDuZB79wEDQMUaJ8Rvkuhpcy4IDQx87pGrP9n5vj9Ql
q2lGlE91mvyaqzdG1HC97AHc6UZg+hdNZZyNKIZhy4VP6PgsYrGbH+cIJJMC3z8l58T7EFgUm6ZW
fjZpqRcDl+18nPXrnEH06p/gW09BKGilIWlBMI9AlVxBD3HChulWvULBKr7yPJeI0h1N/ePrm2b1
4j23pmNffhAL3HM5R3HOlwsY/sONbw7j03Xeust7qEAd5mQqFQuPteIB+2UT4HGa9hem3hNikdEA
tAOqRDa6NZ8tlaBnom/Qb7FG3kE66WBar7BaiEwGaIaKo0n7Tmvpd8dWGjewqdq/R2cLDSlQLxm8
quaEAPfnwGG3iMJ4xIlpLiz9LvuOz51dcmEyw321Nq5elqrtwUF4a1aCCctg3B2SV5tsvTwP/6do
voDtIkz61m1YUK5yNuM5L8+ptBd5Q/Od5tQkUjkSGmywjnWkP2v5RjSx1kvv6TOK4YOJpqWxaY0/
FIr4SBfGrs5ueBUH4y3NElqDgkkFriQAzqd4+69ARWkoepaJGGZza1O06ErJWQwcS8sSauaA1KTV
5EijAX3vC5YlTDTT3nggze31ozNp0APk4glNTeW5dS3ATJx5fXG5VWKyJGNDTjrhGW63cst7FZFn
cL15sBwqujHxEWAipkYROddZGAqL72rZxV2ILHhxmSe+ydi5zyTbcGKyxhbQrc9HOmVlxuaxKxil
WLGAbyK4Xjimgy3JGTt3YonSsyDY/OAIMd7Cml9T3dK66ClbzDUtcjaQ/9YUnVw9/A7gb4cnA3hL
pch1S1t+YZzTxd/nk6PGQCuORdcc3aeaozMkkjBLsS5d+kFZeAJJ+oVSj50xy2t7WIXXFtlzP/2g
J4HH+NVT1dqvuwWtDUv3lfQkqDGEvZKbPq/YOrOHfXSwGq2lBAckQjW5qOarWgu+Ad7iKxzVTn+p
ITJDaBDe0kyMXv4o31DZb8TYQuUMcEeBMxT9TPaxjL8aUJMM0yS0WMKb4hDNyWNDFeL9GvWc10Ss
xcoTkZrH7VUq6tWlobdwWIuIITEuDtJ6ONTTJS0Qfg99YgwkAb5al/J8Sp+kjhcP2oOr9uJQDa3G
Oa/2r71ZpcTV3QQOImTOPF96uznhwyC2HAk8qxox2S1sdhq0xyqxVcr9KjAUFjZTIgTPRAmPnkqx
+EBmtTswG/EJXJGtnxYgTHQ4+GqmGKBOyV9WAGe7bJJSJkOzhbiejmoneFqOQIH900mN+TKjd3pF
763WXxrtMeQCaoPHQ4FKa5YSmUjUkA1d9L5YxPTjia3X2Oxt75r96Y+gf93Pbt66fHieD2Pu7bi/
EPaxMkGMhj3+d3IRk2nT5//jATgYV3vEchbX8rdTNqnbdhXG87pNrUvawlT2YCzvOuSu7wMwJMVz
3D55A8Q+k1V/re9Ejl65OWUgnzTPludq4Gmeei6k7V6jLaDjlqaJ1rSsOvt3f1oKDWg+kvNkyIcV
lsFW/nMrOIbVAo3pMoGjFRWRvOqh11SsPJO10bBM1ryEq2vDHUUHtc5cXM7q2AzAp+aK2o/Ie1s4
mgJJym2a8n6vPmb6Kn2m7e/hybqXyhTQHnmH/JjRZO/lViVa9vXTd46VecVaSf7twpHkms48/RQ4
n2bY/p5W6soRMcfBfBc0tmFcj/kBKENpjYbDN+jL+DqvucjFUIa90jaauUVjyFnzl4FW5aWt/l4z
d6wBy5Gjf2pVHgszGPQPAgZ+CV71HOu98GBHEv7CSp48RXFlpsbfwS2uwL/Aye8p9PrVnht5e0a5
UyyY+2njZ1X4kPP2k9Mk9nzY9VnglXhN8vZ12vpRJAR43aqq59MHsvDjZWA8rlawsW2xSFYeWmfT
Pk0WJpxhkDN3qR3Wv0Fjz6E7zcC33+OLKe5UctCZOGIHRIwqNuwGUvp9gMiUuRT8m8Z8XwTBBof1
VjwVTE2iG3jwaFXFO6scPPCxU3MEHk5gA4h7wbC0n3ZstVtStKo4jTbdMa1FMixkV8gbgVzsCQtx
/bnaaFmkPKdXIi8i1vYmhV/tStBs3kEQ+wwSrns/fPc/LAufN3wb9dOq+1+60qMDDLdWnnze0/Wq
9ELwF+9J809ked+p8N5HYjGnqM18NLXUjfwwC4pqA6yluFE9mn4ZwlpboAZj2eB3GonP+FgAu1rC
f7d8EAOjJwM4Gs05mzv5dy9GRf5lClSpyyGJuaZD4mvnMSylxIMZH1JPd04ceO5nqKiXPwbO6XhS
2R9usHRr6w6FBs69CtVMDtdWxgs42dcMKPQjJK2PwpFduGdZU5/2cggqEpAlkEUKBZwKkXxOJuLu
8FYvXF7bmyMjZMQ1NBD3OHV0SnqvSlnO45ydVNKmlfrvcMvd51fsdYDZTlw6OBrQA2Ns0G8Adm9l
8lsie33M3YN6JaW/K637ovSnG8biMRSdjjcog93IpqoRRycr+w50/LHXOEfb4XbUl5jUGEOHrYmM
vrsO1F/EHpohMqvm8KOpdkykLG+b4JCydX5B6hmhbroS8ccSEE6fp/0aGXJEr07Pt19UxhwjKyD0
PH7pe8D0x5GppyOsC+R8NGTgBYEeAot+L3PfKZuQ1ospAbS0viUDtGaia7e39QKUPYIVGm31FXUr
Jq0l7bLTRShtueZXL2SZQAIa0SkFKlct1H0T8DDavzIY34jmrKra6br1IDrtgup/VtKwXYnp57gZ
8LC6u1TSfWMH7qo1gmQFD7vt5l4/+54/4Xe3E47XfebuUdS+OsRlid5Z3hRMNlBbNFwr2hyYW1qx
kkYl/vaDhv2RixEXC7Gacq9C6bdS9SxACoLNzCg92ObC1JRd56Fcwhj9SbRilLNsDbatQLh6ILis
aWxDZY8YvREXCwsHjl5vhkD+BVQ6MF2egfPdSDKfWAo0MYgaXYCqRafCkduvuUR0xqnq63KdttvC
ulvvl4Zk4B7Xz298tEZY5EmqIf4VJRr39vqTkbA23MUF3yehkKmpeIF070/5uOHqqNbBxSPD8Yb9
hTj6tTGsGVmYnB1RXHXRFdxfOw86NUMiNZZhwXTeDriOFLSIBOpVsJAFQ8dx3RY8K0NOVvsDQYhA
qZ7/1bQBxmIwmRV6E4To+PKYR/B03bePE5BU1E2grRhWKwiz+nuGu99mP2DRrcK17qo+V9ZC538s
v+mvQVa1x7bqQz0/jdYr7VuvVgYNPNdR69OgeCZAe1k1jsYnuexjVMkJ//U2DUSlE6Zk+YoAvM1E
C+LfV0V0Ut3krneWMPNHQSBMgEbqGghXHkj2E433S0EZqlwEiQEB9j9oQKQeLXpzGapxM+pE8Oo2
XcgjAvgKvjxHOYDILzUs3JDRCoSvLiHIzCGsod9uJplLvI/koqnWVqcUBSSEU428SQxHK61Xo0nr
UOSW5u1gLV4shR9VhDRn5QvEQlPKHUYxXpBpl0mLPhELC9vsJ9WsKp5D7nyHqKTPs5qaf2nOjFKS
OE0gsUKx6uJ3YeeQOSGUlivmOUttbKX06iGxAbL/olFHqe1/kST6r3gyiiF4YLk8jN/cA2q+7MDk
hPKbgtsZq/oPVIGIrSVd5mOHYmlh4OptWAmO0KvObExan+uqXu4EmascwnCSbhn4xRaPRD95zXFW
sOKo3NIfs2/iCVrE3wCe+EHQONneJWGjvLjZnUrtvbrrZLupbbSGrzNLEVxSoDKdmnic0x6Rr5TM
5ewQ09/8VL+xeKP3sJstGFf7tRFzQO0GPSMVQNWbeprr6S1Ylo3wfXII+jjVFZt6Kx7/iH/DPS7H
W7rC7StHdhsrZ6nM2uJcSZC+WQZnJX+L6iBKPvFp2ZWJ78nYyysx8TpYmdow0Fq4clMC/kWjL4bQ
t3UslrdAP6oUrCKd3QfB7Ouvz27jsZEdWNszvqdn21+uOJVOiexuCfbSG96dR9HESM7ukFFH5N6D
NfzujuCvOK9PFsd7wWBMKFHJZZg9LQGo8b4RNmCr9htTpH6JLS+EW5Hgv8GYAlexMzSl6k9hGV+c
s8YOtX60aFlVnrdSABviDB6i+OnFs4GQGMKjjK6K3i3tjSjAZ9U9yM+kBVz7JVZfxwjEGHWsxxO7
NwVL11W8dJXbORh6kxS8lTRX4C4wEN1TWf0j5ixEDrahEIDxf9o9hLskb1J9/hJ9nNy6f/tkrRIM
/DYLpjLG6hyaM+DZtz5W/GFjCP3CmXGkogwc3yMlmD9Wk+yvFpyRr8YN/68zvhdoVPsMYyPk7Zku
AF6FrQt3/u3Y4mj3PtXmczECoiuhmJ5mWz/+Msybm3zRiDKcZz8bPfIuhtsqcj/M2x+u7zmV5fbc
f8+QDPB/7GfneVaHhXrUvgJPGZexjwAvZwKVClIrIYHKFTob/qOVZtdJsxcBr0MU2eaus7AlLycY
JrSLOOg0CA3PUhzqAsDnnj6hTTkEOs7s74rASA0//xcaHky3eMWCLeI7MzHoCbUDroP5bx7x2RyB
f5GdxV75HPKdqp4VaIefUwz5Yb3whAo38YnmtgjBnQ0zIrNKWIKNgNGW+kbicX1XjJfs8DpzbwH6
KpStKRGGbDKDmmziMYTfwb0ZZFBJlR3Bg27VYuOkk91/gfay7He6i2t5ZsFHbVwXMjwdesH4o2ll
tc4W3RrT0PSlwjn2qHsjt5hEgAFzRnJl83IxZuSx9NYI/waUx4H9LOaV+QKBqzQwamAtk5zpQEWP
AbmAqxK/WkK8ep0atZ26D24pZ4jMYADlbvcEh66eTHO9dngQvoNJ+Ntyw7vKBfEZZxjLjMTz+Hr0
VGAcX5fBIVCB/Cdhg7x/2axAUflXoVvxuDXV607NMGOAs2bUoHnFWbS6leNJsF0y8/o96EMk+5Cs
vsI21KG2bK5EOMqBcVmEpANvPGxeeaO/YAsqZc9rwDrmv+YjjNuPY0QqtpEWZbtZEY0cannvDXhk
HDBsIAlfNoIYv4IT6brgVxQAJ2vc77EBzesEyaZEQnRgRKZpe8DjPNwStEsjNCAweAC+jwnld/sT
fwkgx9RlXSKmWELxjP7Otyoo+2f3zpf9fRTi8Cyh1kbQX0wOMfjVBVLO97g89ri6i/uj3rMnBDLY
GFY6f3HMulRtIdQCPxKewj43HRqu7sy8JnkH+FTBq/64qWSGLTQ3lRlC3r0Q2DhPVa09ZjfFuLjz
31s8gMGBHp5O92GJvjZxDkinjcHuavjdX9evZr14yQHAiH3rfRenrsHHBYwUxEO3JuyNxvVCJSDN
LoOHgkc4sLTX2yqoN+Ovna6x3dW8up9gU0ytlgJLCafYDvVBj4RUEXU+Y/s6PnUsOIyUSGGJoQdd
Qj1k+beEYjpm+9ZcDwReaXhWIgmE1fuHW7k5Y6LMv8lpSH5FIwf4shU6rlaY+e/Tg0Vi0Lgw2qIB
77OYrLNxuESDBUkizkWLz381nTw2Uh8968WLVTKtv7taFRqRjzGoo6Hjxgvnn83fiNQukCKD6beW
UnowX1vgFIN75bkCtOxzxG8Slw2MQgl+0xkhMC0lTidU6p88+MR1RM3+TJQmSbRyN1ycx4AV5ukR
B1S9xRRJmzPxRKdh1Thmc+NZw+jU8ZVdh6x6vm0I+r215jCfwUxHao6wha9aeHj1NE/HBnZYpDIH
ieAJmjPgHmg3Fpblb6BXgsExAHHqE1zhT5yyfarWA+BvV/uMBIX0MbAAdXw8vmXrHUFqOPOneWdo
3CPC47VtqCcjYG97vMpPzvGfnNoqqYEqJ94Gst36vfg9gQpE68y4eTN8fnvHCTmH/w0HHdjflnXI
ftUXOPS2lwNKk9J41KHHiAPlPlRvx04KF9vP6ckyEO998rKnymaXhPl0tYKtbkPVGBpN9WjB5mT5
TrDdCMy9wtMk6gDUGJ5JpaWp8vkKWZFZSi83NY1vuwju3qW8pMXZOEtsJ4JVYSsKCl60JQntkRAh
AAkw8fjjs8MzBBPTLjBUMhwKYpkmRC5K5XC56MGob7vFsCdTVJVmOJv5cIw3dMm8nrZQHvcUeNlX
RdfimQ4ysmQ/8o5qvSXJDL3KMKzFIrSQjqSsHfIPnL1DUp79aETuvSfdFzemniWpZrIxUSuAXoDz
/Cz5UsiU9YyMSA7seRwyShoQWXRnJKqIOnu2POCrGUcBhPcLmP9pQjVPU5eYlY5FHSBi6pL1oWQL
CHCIOLbKJjgNaQXP0F8+rlKU/vjHw0tk7pyZJJ2W0+akIMbV28BxANObZ5c7DS82G7pvspXhl8Jn
f6l274YoKs3jFTSCU6L9UzdtSrw5Wcgxu6XzAYDElAT6t1EvHrGNpVbUvIZp0BjYEL2j3+0LHi5Z
3Q4klO8bG9RbjLCa3AKROITBwO66ZDoogj4q3ynVsPX9hKXN7jKtgZ9ev7vk+ErtD4ADwrQL0whG
nMcyU0ch6Hh3Rqh60LF5COU06JoOLQBzxO4eL7tCa4tR8gd+0OFzflj9kSRf3oTW4rU2wB4VYekl
CCxvFUTM68Xova2kSOOh7QyTrZGdMoE/7KcUtyok3wuD29pAYyFPWnznNyLFfpqKWKeUn8P9FqkE
kggv0dpA9XaJHpOC8T08VEmVsHYIBbVwnjSzLYTmoFmt8O4rfWmMDA4MI5z4VDbCcfrn3ITzbZg/
YtTgEjM=
`pragma protect end_protected
