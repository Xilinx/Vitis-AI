/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 301456)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/3+b4xjRU+4LM6X6vvP8fEfvTOErl1eC91ncjy3tYz19IsnjuJRHGV2N
zP5z2l+PBknnkJhKjLi9ZY2hUvMYcrAW7vitUHU8LsfqNIrdwIn39QYxtQjNs+em+6WgtrbTON2n
Qebm5Xh26xIkZ+okReyKefgxhp8t5DFDXpkpAbfW7GgJ24mHc9rwPCcsitlWRKt9qiE0uC2DLGdc
SUPozQPVkcU0RoDQJE/vwrKhc0XoW2ZBPpigcMsNX6MLNac2tadZ5XqF2QUGS/i8zYaXQMuSv4dF
7tqbFjX6jVAvWqMR5RekHyGt9QpzbxwaDOHsCvBGdVGS2QWh2793B+P/FLt6ckxQCytIJxHc53Uy
2S+Hc8yI/0Nqt4/nIpAlmWeba2rYLfyshn2mdIRDjp3ct2Xn3O9YbDaOU26sEclxs9wrL3r13erG
hOtn22FkGsGWR6OQRDivqFELuPGunVpo3NQxhk4N5hxxRBVeZLAVdMO42QDCUUVOpeNt8SnNC6xW
FIRxB8K6rLY5L8MhmmFw9sr6Js9P6VIrpvSRtY/NySA7TbKwk9lsOhfgKORnwRKFq3IC73RIlcsJ
A+NeaXZWHlW6lSWIjLXld9L+rDXFC3iSyvVrznQV9Mp5AoohA/IqzPnQVPYdJALciFq3jodC7NWl
g2hcivHnXVNhWpXWBZRyI5YHc3JGyhOlaNAvzmH8VGsXMCkudg0302QAjzYdMScKRPRSB5ZksLvQ
wFynFdSKtx51068wKbGUpEa9QeV7/c7gUpCqL+cyywDwHYuT4jjrio5priR8U6hXr3h8trOU1NYz
hZfsFyRT+0E/oW00bEaPyOtr9Tsu2KA43h+r0RBpAk94X1TGDKNOp7J7kZtPJAt7OD4W2NjbY1PE
Dd6BSO94w7VNClHLdRKXoB2OZjC9RW8MWb2jqcwf5C7LAZW8XZ6tpDKdQu2MdMEbbe0yY74BMLva
epXyBwO3gJtJpSgMS0iQM6bUgxdWMsGrVRyWWbL5kEskGMHQ0Nyf6njrfEy5bcYl13/10oofzscO
m9R+zffxZIhgO2AiVcxDbyIINobDoOO1IYT12EcbSwIxUX+4xW8Zaz83o704WXJ/3zjlK7Y9Abwa
JcNv4YUycgE+a4LpH02wJ4cAQ1kecIH9vvC2tA3OPI9i9UXb1n09o37M1nlcc2zYUL9963KE5hL9
4Nc7op9GpbapHRIQPglxLTFpUuAvjVjqKAosY6YaQx9raWzz4QAw4vpciQzE61J9D77NqXeKRBzt
yAkYICSCOnB6aUQIuoVxoyKTZEKomf6tZM15hZjGeLuKciwhlx48LoF5tO4+3UReAyFK062/jrAT
aeITxo3eizgr78Po+HMHFQipIhITT03cL01UvsdIyHgtxODcbZ1zKviJsW+rEfJYTpWrZgO/R24n
K5O1rfxWbxMI6uKdaxoqz2aEu7UO1QQPbiFwqUmgNBWjEo+50g0ZSVOgorGzUYJMHH8O1zKHr0sa
PHTCJvqMWDzlmZdbh6XeIKhO3oBz7JS8+nU25UdJ9QwR3kS60cHnGC9L0GOzrPMmhMCc8Selndx+
h4+Fbvj2R8y/sT0pPaOy0nVuTR9/u+cZT5pvcdaE7asHmPGrLQ7mkDdlk3Ku3vojB67N5UDYfEa0
Pwa9a05z6e94hQCIowIYedSclyNzcKlgnx3lZqkiynJX52mAVIztnpURra+tU5iJeMffS+Ua3Wns
Fk0m4zZTfXcq8wm0oQJ3besRwUBP4UzaZRpWThbF54FuebfRqEpEYjs+Q1Cxw3yFcyKacd95YZIG
MxpM9ZbKYQSIcURLElHvkKrJ/VNLvuQEiqBaGHdfJXx3qm3HG8diqcIAi1QQWQvV2OzdDcWzWqxK
B9qOSrNJqHihUbvunzBYAU6a4Hy/qnhwN9AKBions6xfMTWdEfDmsMGERzMOs84SXEPX3wYCly5T
bTJa+EBXwJAn3AuHIGId7xuKuAjmXg5GvmnUUfFfqjmHNZjvmgfHEzZzGN7g6/6YU+v3Dp+rN6TQ
n2VEAmr5qO6GIBLOZcBP140QI6zsGp4KiHIFITGYC2LH/XEdjqj5b71LT1Ig2BQwk7LRnJbNTKiC
0RTeO6/Q53gHnLbzBHKrKjGpaHE3zBm3jY2YtggNTslnicBxSTmCLL1nUXqXv0si1J8PeLNFgfUn
aaZZy0pBs5M5u21jEws42tcGX+ESlS8mCtOyKI6aToo2fqQeKVlt908O5KQUsfui8hUQEBLeanBN
Q9zBLdgrJRWlaTl0viGpNAER3BJTOEIBInzeiwpWKxFdPZM42x5a1/REqTo5RBPqmfzbcOeW5tIY
ix0mOA523lA43PlSCcDlaVAxLeGeGLFaa5iD4KEJzHYlSgADXTL8158cmoY3hMiwco4C1vSP6RtC
6Nfj8P3zG0Ul8O10WzOShAJ+8fHPs8Z6fcRYeKUFPAQ1nsr6QVNxk4gpGPfv6K9TzrK8cL4SU0t0
OG2ebHzw76CFpkl6qUlJznvdlhNsHvNW+Idx2TK7hyYI2Ti18euO8Gs/Dtaz1ApXFzgIv0Ko8ZSQ
BoOza9/9wp2SPccX1d51/0gCSqj00IeK6KO17QYseqD9Qsq8yGCZL1CrkrE9bjPLVlJW+Ztuc526
LWTFuiMK9MrIorn+JKEwGNgt+3a2ohhJJzmsFCpCAy6qNF6CBjmC8OY+WAeiXhr8IUSnYb6FSMEx
5NAoabl4D+DsvVOGEhPIcEvR1EPaz3a7MMjJvTUXC2kJf4tGmaTKPgwF0MeiayMMtzKJQWaGWPpT
TiSc/T7E2aJTcWYT6w7SfAuJQ8f8CEHXFUDRgX3biJ9nY5hYclG9xZJIUbWJrVf8amzWVWeCSerX
1aWaGSKJPp9yGB4DKpyGJoNMLsKk/UI+lk0KalihfmD4XF3LodeJxUbWZn+YL5tMR1HEJBxjcDbi
T9rXt7w94bKcMZkXhi7NUEw+z3Hg9ImtbLoj/x8qjYO3PUi65DROYMJxSnL8/xU9WNpNjdW0io0w
7uA78JFWpHLHkCUtYe+40uoai8xRZewuJN9GPtPBRqg6xMHxLygmkiYMhDY2HlGV7XvjZGZT9V58
4wYcW7EyvtgjlVSiwf3B2MZmI6xju16fe4hxN5Ej3c3wiYaOl7I1YsNK/D5VmLoBJ/LD39O4CoZ5
03UhNlGfCilQDaSuSz9xLDQkuS5IoIq2mjNrv2hp0oiH8uLsA2achcKau/l+6BAwE9cFHNwOS8Ik
H1OyfVd1bR8D/CSeEgDCYLPiJ2b/XEG8XdtIg7iQKOEo1vwCveW0ajO8z3mjQdz7ZgpN2Vldfkfz
zG7w0xHw74mx5wzA9DCWqtumpFXf3/BiH1dKx0KTB0hwxU8q/TRojmcz7kr2Pueb9HgzSPAY4rwz
+6kk7f28uadlihLkcxw04qbGyalwrisk6T8IQdURdjbgVEO5DdSyODPGFhxH49pvlC6baDqjKZxY
IcdAKpOWbW0+ym5jTtaftSrxr31/jm1Hll4PPb2maOdzCy+dBGjoNpd6Q5XP+WK/G1HydiWy3B0U
Ddna8nBkCkZJPnmoc7Xts1gapx1Mj3qRFLGqmAStu9+dXZWT+04y9ar8WbJvOZTtllWaN6i5HyMY
9fEfZfWjMQXNzPqT9XvWK9yxQ37CHsw0/PiGS6OHqOVTHRS83apC6GUDASeTg2hAKP9NGE2vLKDP
5IWK2ye3evfs0H9qZpPLStskfsVjuenMAc/alQNdlOQDaW11uJq5uoB6oexpkXyy4XLGP411wNa+
ETOUnyXOQOPYOMpVJhQ8QDnlv4NrARfYF3LckPOo0AwwWEFGHSxFDGmJJ0JtQK6OBm6tgfRBnC4k
/FcAE+c3nR7jOpDmFUkiU31c6LUKfOpl2JlFcaAnFiJvkMDqBPHmrwOYmeWe+zzdqTY+qGIDWChW
hjuxv93JpbiSDaLZdvBjs8hjMGbeOEoBN1mLruIVRYWVB25rrRR5B+2Fjtbxc2e2aS4KBpWNY28n
QZ797VJeIJiHOJ3hd78Kd1vTIQq1YzPDcMfpZlhsH7Ws4Go268UOCMmy/z4d9rx6mPPTBSxlyNoV
6D7O/R04cj6TbZaHFmegqFExVhR48q2apcDKdUzX6TsPWEd/A/wu8rYCTrLpVXdhgfF3dRhfkXMn
vaW8Qbiyttvv1+5ZgyHKrjHuyFH4MkFSkivehlrkYE/NvV8cc3YvjvE7pHbmblBlq8rUdWByFNec
m8/Icc+glUwUmohPsm6vyvAUo4GqriE4vMb5UtQn6NhnAYhroBw2HhvYNf/tdspxm+usF5cr+nev
+1siueEYnQNvYw/c5a0EVqjCX6O6539Awumb00Y+U3pwzJem40mKdfPziNgzIH/Ki0ejZrmjAWgq
D83a4Cw9raxkthL2DLodEvihDSsN+yoRO7LUd5w77o1PDh4WY7NSuLdvDLftIhj8Cgv/hxnPdL85
1DRsqXMRrtZlA8P8IxJELCP3sdcaRfxNE0sXkvyWNMSXfjVMbsV5+xm0JQP0+71ZsbL/NF2iw0O8
Ogm/f9MSf/x85+DGXjaGoioxTQ9xO3QIRFWOyhFIZRiqagmB7URZlL417C/+27qLg+YXIUHakg23
lLWTGSv5JatQicFDejzS2hqxswMCk70pg2VIHllIUyDJg5ZybbFvHTRQheERK17iA8Cyo460vQMQ
9zdCgrCVrqkq3DD7Jbf+X+Wr7jRSYe2DqIQgUD/GDutB6qaMqtTKTG/Hq/ljboDEMshyrzf7K1m4
80qGiYpJSCptVRzVmESMQJdSzAgv5SEg7Dvv2PgHnBmFfCope13Tl9qBg9vL+S4y50irkY+p0hr7
vq4UYaUE/2gh6S57V68ngq92JaIWI8J93Vgo5ZYx9QgBzhCN6p3THkJgEpb4dSHwI6AbEv49YWcA
UNq+zZRqV6A3/v3OBVoBmgCy7D9CMsIkY7GDkcIjbQlalTtretjuwirt6SteXl+ILiNpweQCp+ba
uKo7DywHq0IPYS6nS4Kzyfu4+WlZGCAH8+5ysGQgxPd0zXAmrEa0/KEbvB+Mkt0NpLBko/uoncAc
pI2wLb3d2v0b/F/6QlMKGULbR5h8rGwB8tFYl9H+irFn/nMhJYMO70HIVXOJFJPi/m7ce7CLrih5
yrHzb+ygDkPvlUJcRak8GiEciMC+EKjtqOqmc7fcgUcW60zpo2lznwyeaUPejxGfasz3mnx1jWzD
IyRqPV9SD1OQRR/of9v/Ljvq+7yDL905yQM33BkDe5JqPugQkLNaT7fUEfrxKqdTP5b4PgrCd8IT
z5rI21TAmq5jZKpfCmzghq9WoYUghhj1aHxVTBCFLallz6kT7Wrusye1VUAuowrXFCYdgFB+tjmK
dn8E4zzyXpO/tLGSHu47R36TOd6Mk4iBzPhSo2xSMwyvox3EdsrG5KwLTyRQSBU3iBfDS+lvOCA8
TzpF+7PjPGOMq3bi4JTptL+6xZxXtp/mi7qWz2Th5BN8lsUXn9KCCiX9upk47BrrCj5WkyQqVNYK
BzVgxTwd4WnKu5Ha9+Vu+aiVlEtgS2QNVv9zBd5JgRSpFT4+YCelh4lQz5jMluFRjMNIrnVe4gZM
aGSpCo2co/KEkYPdsye+zJdPCTCtFFAObMNT6gTbOASm0/BEDMnunPwxXOdyQ4owzc+QTCs6E8fE
uD+oeavE+OZFhy3dRg3lB7E3Fbvz5ULjVygHtXFmmyRMy+ndnmkHuL3JQh9NJwrB8zOp0FohhWiZ
g1P4brliOlJxj00kob4WdbK21Gxc8O/VTaxVI+yNcz+8zFQGgvawfTPdZekXp976oFSe1Rxjp1Xj
GECi2ZL2RkAe2oshzNfE2X5tr0P39fcdfDJMMQDMurKSiNEfh6V7BHxba78axT/uLR5/UZanCIdH
dNB3eDhdaIuRKR3Ruk+0vPvOQTySSg2AzFXE07v1KczVIlprvEfA4WoTzlQqzM4h6w89PnLBpr/M
oAzeCtNyRQxHnErCcZsj6chzkT8rIDYjIAca3xKEnHB07EeSQ45MC4ns10++0+VLd+FJC5rd9FIv
94o45GQPTzAUBQdnmXc6N/FfSkdK9GqvzccHjo2vPTDm8qKmW82JBNODh/kPdbQ64HC5CNCULCKQ
aez+0lT+dgg9OCzYWxbpW5Sl+6A/h0wLESEgvoEnAI83gJ5OhOA4Soqltbm8Xrx3UHUVuhkalqkf
ZLgFR2/IcPmlUysQ09rToFblPiuBbMxF+mGmiRGFQ/JK88WPZkiFZFAr/Q6aaS+buMm/GkVDiomJ
LDN0n+pjYLwBu8cU5/CdZEOmoRZhUBk1aloXGUVWesOB+PHkqrCGq2Rmih/OQ3E/UEsCvGEvot2d
ujXyLtx0t+BE5dGRuELSdYyMpJHVd8/aJ8UiOrgUGJO4BMDNMW7d+9DmhY7DflKCTApemZbPkoh7
Qyt6Y05cIG+0u4YoSzqfeUq+ccxEDqWnb2RX+RX3VyyaKKajZEfI3TXdREvdqttEEqMk1tOOgOq+
t6gCIiJSCCQuZuk0ht4bgaIqJfToVgG6fsrwka6ZbKY2h3Ymah6joJPH93cCjscAWyy1bb0SKOny
AAZ+PxMubBV+1oN8ZB5kEgjJTENcsOBiaOCLOb1lOUVmi3LtXuQqG+ymevJhVTTPyVrWog9VSTzz
scIoVK2nld7BD8yT0esyx6l/UpPltolPyV74li998VuAqGY7mGL3ANu5GjtaafVb2Cb+IxJIGLRP
LIhml+ZQEJLk3SXLSA5i6JKAljyA1p/MhkCgkzSSVCopTSS+g8um9s0ES7WBLs68iYoHGE7ZXWpq
pd9Yru6hTQ98sP2obc9YUi7i6wurBg6GmOVHWrD+/rqJY3FzNg16/jq6sk+HZL4TdY7KDfLFAtID
hnIWUng/USwx/EHfotseklZeyWh/cN2nsHWo5P4VX66pV4b82jhWPkNvSKLnNkwrY/9weGi0J+Oy
P/6sjsPYn0/eJ3DGusNs8s+7y3Musxq/fbatU23QODEm1fwcthckz8QtKBVL2/xjlTNQBO1U2jtx
v/WuoJ8If8DsxZA9z1di3CRZJfJTg5PXNWiVKFf2jYw2/3BcVsBaNi2XhGqMtv748Pd0z7DodFTj
718FQ2sjWbCNg2oN9Jez1K1ChEsib8WqkzSVS6opHEf5H4qUeXLUbHh4t3S9mqCHoGI2nocQKhwH
E3x+FqtOMllFXrUWLf1m5CntY2l1KZu8J1sCJWCYX383NVhaUwX9gbFZZ32De2cR8MheUsxSNSNd
sP4zspgNV3G65MuEkClHKWILyb8HYQiBFPe+uV9LK25o/7r9KjG9GBw0Aa/7owPXC4kFxB1B5A94
cb3XjfwJ7kaTnuIDEIDrq30JdW/UgG6IdCVBdF+efs10B25VFezOd0Q6/Lfi9VkoWVR49rSW9hYX
ot2fwEmPCZyeqABFyZLfo+wYHJ6RiLMCvG9n2xT5kSYisDXENN0B9Dv9A/9a7i3UayBwwfNeZq0B
OiyajX23CGiAAzx2oK5oBIPJA0HE4k/mjbrhGKoH53sSvUH58vVE6fEmWthiTR1JR6q/iNm660eV
PhCWjBrtzFwZ9qEdHkM+Zs7v/tkIv+P+MvS6Ca/cucBMhkvYvXKFdXJj8Lpn8X/qW07poWK0g7gW
dOgJGc10JmwFpJLtDZuYUIX2zYoxKHqnemkD0LnqHvr4H19ZupyujmInh0W4dnkYIWjwdBX53Cs4
tmAQV/US4VKNITANwsy+mBEwwUD/mNnlAZxehPG401uAKUKHKp1OANA04AST3oaPZgm9JuHSIDbR
B72ZM9ulI7K6Cpc21Ch+qp7bkDTnE9RFc0sCpm65cp7d4Jp7ltW1DQWU3Ow99UqwxAIBn428IqmO
o0EGJSQ5B/AT1FMg2aAAEkjJLbldwda9OnTCutzjKjAwNPnx4fbFubNxvcoUQ9dW8p1pWT/qycMn
fnT8v57rbdqfwkjV6rbX/AmMeCoX0Tn2ufCHTpVr30u2rCixl+poTOMkUamNY/Y0k1lExtvSM0DQ
td7HIuxL3VESKubx0gv4wLCHRF7STH//r345/G9md1d0Ttgpw+pd8Vq7M1b1rgcMl82beq5jdnWQ
PQNzBfSavU2wiQceOEOBp531u4oqYHY+luHmDgTGBVl7BXX/r8Jrdfa9vPNtGMR+9vm06p3HDHmQ
ner3J8mZ+aREqmrofx+KqAfTaHzxWDLwBlj6tove01OWYPlaeC/doUovy1G/qiou9/DZqCrsC3LX
5VhJjTSIucfImXWOFCxXmYgdkFm4r5k12jjfA3IWx5XNFRfLBVRPu/Npq4YGuVNKnyaqHOZ700kr
lA1hhDuNBqokHGZCa0m/5NKXxiksy53Oc4bvg9tib2ru0t3RJpM8EhKnVehG15U6sgLxum9R4qbr
ajd8TvWV/jC5vaYNW2YnoZVdOFOyowMSGM+VuEeAXewNr4dyjpJX5jTkyxLdEZBLJaVXzw42PHxF
G1bcdTPikbE5jyn8HOVDl72sVr4hpT/fO3PDoZfV0UKS9O9SO0PbGG+bRaXQoJ6vQ6yHOWROiIb7
A9vU9MK8zQrC8wGeuUpBQzzK4S7EZY3+0Ruu/RF1twcJLkaTSDOH5rT85ocd8QVT9lY+rJF6I/98
ecnf/ncDDsO6gNCcVWLoXT8N1GgIO6Vv0xCQROaWlRLVrJqZitj07GlJ+9qEBn1huSjwMYQ0HnQG
p1GZQ/uozLqL8YaiKmg5s/tpK2ACyEzRH5h0Z+elXqK87jD/bADtpklQuwbGORyewvt8FICuDMQq
/Wri+1NOHPCB/72TnFWnrBKBd5ZxzIrO4FVjWeOvSoIAtf8IqvO7E+K1li8vJh2NmeimRHFi81Y2
pJxJOTeiwUrhLRoSGcqEBTPNQGpOAQIxsd+VrS0/OEZ5SeiwdJCKuTqAcZH3/NzYbpXjWJvhcibn
gX5+5F6puHkiJr8/L0SNt9lTXkk6J8EcaNU2l9SRC4xVlA3OxUsLIfKLatO/tkt+yJBTRMKhNNHL
UYorVdOs+GV2vw406g8nYCg1oX5/U7992rRuwHM/BXo8GyGU2dCNwYGJOZCeR1n/LNsDJE7JC5o7
liySHB2IfH+Nv5kyaYB7xdD8LpKA/lIGwH+zlTGQKyo5Fuy3/QrVb0e3+9RWQHG+guS6w91Am3xu
Ht8TbLI/9WOZ25IgScxrAJLxnTvnKlWk3scCO1pP7Jb7OqfstDw5NIh1ZH0Fc8ZczyeU1MWUbDIL
JGLyduv300NWre4e3bhGIMroF4aMGlo2oSXp1tG3cAy3KXknr3kHoel76ryPXjjEwUukhwNa1S7n
brsS2BDi8Cja1M/aZdPWPOwnu5+C8YTsCSkkG0mXYvsS+CGi8rsFVmXUvZcmUKmbH+JOuDdfwxLF
MBuxl4Ce8Sc7gY37XnvxyHseMBiopPCI6sUzFeKx7doEV1F5IE+pxnb657GKbClMP+yNFlTOaWK1
XhF20DCIAQc/Y/Q84pdaAuk3pFLIrChF7RsyWIUhUDRa/9C3TRJ5SVrEjf20mo0S32/OGS5n7cWN
J180gVTIoE7PVbFuUSR25n61NGskhLj0xU7tDlqDziUAcWUx6k+48gqzEeypoRemCy/gyzGB/AnM
JQPTOJ5gX4otzQhtWeQjL+HC1vvAhcJgGcZ0kEuykehMJuv0A0A46b12USoXr/ln28c4T+qX6tHt
lAgH+3FQMHc68vDrOQNcVCmyMOUx2rzCMrAMdiBC7Qt27rTGq72qd1qctYVs+FIuFJ6nFFQYCqC7
uErXhEWv2mLdsPbIhfzLrCV3Yj9Dng3DUUCHQSkVbED2jlFyxou9cSdOdiud9zMb/630FaEOgc1h
Nj5+qWzGluOw+PfkdYBs9mYeVfTHiqZ9vo92gtm7/qasEuVC59z09y0CkYjHdC5HudILd4Giv574
/CQUhIkiuwF3UB+EGv/ZR5LkrVw6C0wFTPf1Ub8Ih5KDWFNuRBA+Z12+ZNRnorU2nMCYGJFdye7M
J8XWGCd0cVYWWlenaSu9nXUPQ4kC6XMyml7Aco8vEz/HweWNLuOcBFS1qwrmXtfS6GLYC4AhRZLY
FExpJwT4WFjpvz7VKTjU2DInje2ve4QhO70kh3ojmIpqLSZP15xQy7K1RLXCDO30qNjQ27UkUUVC
X0tciMpWJpVa1lnQVuDyxVI8DQz58CiJnM5oArXq4NoXLpv4reFJsseVzut0iOS18Rf47SiCfvFY
+o1sQbxBss3Zex8oftt8QMAvbeCucxnlQwjoSw/CBfelEEqccMYKllmXwYT3Wxu9Le+pHR+8Qp8v
/uWjDfbqT6OwQZMoNee5UjBv3iUzqydK2o0dTqw3h+OZQQ/1+GLNr1/Q2OTkhEDwbJFUPC7hQF1G
hu2zQts8tbebGpVoAwGddnM2/PSNc2Q25IxioDK9S4aJBf+mIY6VnCYOHcCNwxqUdwOj46Hp7g0w
zBHu3YRJ/LjJHeLXtl5n1kZg6KoN6Wcm3Plw5vf2FRMZyZpopYOZBd4ggLryigS2qWTZF+o7IPA2
lTGxK7DcDg5VQf/FPYQa3rdQww91ekScatr+B1MNnTo9tr3X+2x+uHvW29n3mvz2Ahkul5P/hWQP
12Bh495PHIQ2nac0gr7s+pZAQ7G2H2a5VhQcqwQrNCBFKJE/zZ/Q0U1Hn3WxtlCpu04mTNjv/Jtl
Vew3Hi3mAMP34u5ZE/o8mE/ZfnkikKIMoy0TzQaFsIKPrSEmI0Uowg+7P8jjPD+zDAI2f3cRcnIo
3q0HFIKs+5QjDzK66txa49UPQAguVsC3+lFGqyEeTnT4qnCsA2Bc+CH5qx72sJdde8dsA1Ge/fGF
0YN5AXyU/IX/4VQyDEkdBOeM9Vjardn+nI9kNFQgZR+wlmJfkmA9nG18yn8vF6D6BH8drVLPeQ8j
rTUi7AfmvXnvdMayH496vrgEhdRtcdsFgSORg5dQhIdFgCnUWcIBgoqKRFu5N2R8tpYGm+Yjz1YR
Z9BOmHQnYibvWfygiCzh85AxWkO+nmu7yErNBoTZKgeh6Kr9QonJh9/HpSd3o1LB1qLn7WTgCIIh
57CUem/60viAgxXPGuwjBUOP4LYmUVJ999RnaC0A+JVCalXiiCeweR/rAkFI+ADa5GI5I97f13/O
bEjwFxUBzDqmTJzwg7Adm3xNq5EvjcjNHoR1Ymi/yuotF5y8YLr68TA3fFZhSfAllPxhP7ubQ70l
YLIUNEaf+nVtS7AHnSsiGiDOsVw3Hh2objrranmYSbbC2wM6lGFNp54WV2zGZqaOAnHetf5qtlWE
Yc3lnD1O1OvP26r45dPxB+7TsZP9LORnWAYZVDV84DM1psjbQ6REiVl9bGee4A/VBhzAWFP0dnCd
+OthLvnuBmkfIiSLPvezC+q5wxb7rLJnuVyrfCcIV2qF52l8C2bcQ4l9MMbemc3BpI5ayaLQCjY1
vOlNE+Mmg71Wp4bzKRVmwqVyNjUw1VqjGFpfOEvfqq2vePa4aNmD4whkRt2B8z1/1zgNOc8bRCyQ
J1bnyJE4KH/lEBiVBvjoFaMol5JDMZy6bk1q9QtMfUsc8W1BXUKlcXZhjYaos0xEvJueNyUItDRT
cIe1myfcAnXmYUIwzDp1nwKkiqPehK7oEdxgArCiP2SF1O/8qgmZEqtTl57Az52bo9Us0VviRzCm
cPs3/MspdEvQNmHdEuLQ6ZPHBvQSkbI3zyswpjYbCwWi4ffIklmu0leVelHISaN3OSXke0mWBZ/I
coXZu8cok7vebwd2AUv2Dr/8w95xWOB2tKgbQqmy+5dcSJQmHtuPvUy94qxU3pUQ1SHwPvy8qTHP
gByuaZ/GgA8ZLhH8cX+USSs49qwuIF+EnLFnrSNVho+mKFI5fhC3ZJgBbJh7R5MvIh6ZyAxzzPaR
ol2gIXZvsVXDeRMcDNLHMKqjqkSaNcHeaqCKdIF1+WGhR3zFkh/r2yJHSE9i0W7SC+hKSCGcExAR
124IHfXsesv1MlWAJyejAjWPG/qDBf4jjRRl2n7uD+j3fZqlBOeJhWF8YUabgt92tkVgVrSEfMPT
5Jr3fCR8vGUcSV3qfpkHEBLVROMfr5JvCFup64E03/6w9JIw1AbEQZ3daRPQQlZIfQ5dA5nFYXkp
XowrRLM0V8Q8zfokTsnt019BVKMp3I+3a+2qyoZ71xV/zQfBxvU+N6sXNyzAvrIuCgidC/BFCpaf
2gWoCE6WhO67qaIzz7Kyi0o+Nz/TVbuccRAQVTVf5BY9H3TZPJ7vQ5fBKHj3n12TXM4M4Qym3QF0
7olptD/IszCBKY1Vefk3Byxc+B7SNchnAoMzGff1LQVAUrJjwY8axlSGEJ8pQTrw5FqhqGrkXTUD
mhv0/jDOozuBmzXCBXh1js0Q6UBYJdKOigwle/+V8hOchmmBilwiarei9QWZDskZx86DBss8INng
BQK72ppYfIPySvHpe+o+7wNFRz7YIi/yeDt5SpG2c3TEyatXMYC5sXnvPRlHDUuyZy3NEYDoD28e
H9SWvhdL+2+83P2jHw0z1CF2hZK+avSVzm4m39sLukNVuboQYh1yynh75KOh460bqqWim2tJRpPE
l6M/1fvN7AYHLmx5X75q/fVqM8doGpSf7BygC/ixe3FI3emdpZ1x4gRBcSe4dWnhflucSkv+ikPd
Jh2ULEIIUidUl83a4/2h6xJnEQsXeCNdH4ojnQUHVmD+E6f1iTXhZX6l4i0VYR1KQUWjwbTNyv0P
LGbKQGSNZqiHMrcS4+8WsC2ocBDifqOWVI60tqLOkSgs/a7J7vwm/q3pexiV2eM3a9+5BG+bTSKS
Mn/CbEVgAwgV/iz/0U0UWL9SsARycLb02saj4nOC7y3531EHbBrWqTAe50IyCXmzpZBUaqR8Qeqg
hwGBv253p0GIBn9R6FHm+h+CFGUDLNZxbiUplKg+Xvhj+WBQOzPO+dMLBCF4fpGEssM41gSg1FmO
GsR7zjBroNldYJ6iey+Y0i/7Xy1zQyZbOFVa9oLqcvmkg9UXuI4KTLBbxwJA1FVB66HTABRcfCsI
NkD+L36iVxjFKm4mpOvECJ1dv5yEQU/jxox3gaBt6oaKaBRj29tZ1o/3/DfnJVXQqBudX8josBTJ
pzCdjZi8rAersVQz6fMajstb17xQ2Gs8MQ7k2J/RvhFsn64yUkBesNPytWCVbgGgZZQx566sXAQP
7ge10zU79HzJJ8BGkTWzFW0P4PwfwfKcus0jmIpPWnhDFIVp8yZmYqwbdXQDHiAsn+G6YCilUYTD
RQ8v+T9ntynbx8I9PdGmGMjmFqxn5nX3rPIxqidmMjN3D1tefBkrUmRvRudSG5+n+GF0zEq5jJeu
BSH0W1O1ztQcWQsdWABpqUiZCq+5WieH6FsQplDV2d1qk4HVrHcH/3S2r/FiARdrrguF7xfXf079
eDu4pTXEYlRYdjkyCf407b3zWJtnb8pUo8AgnvEUe5aVXqgiYW3Ule/459bZp0ubqaPl6AaQS7oh
TxydNHk+cKgZaxrR9vN0jQwq/1j38J3EuZxO9rgvy9S/jQadruizggkQKq5xxB2H6p8tI181s77o
2lB+DhXPfVz7x8QaTqNYLM3wyhkwEvEOw5OCjov2aFwydRbdu3x1kGXw/dLzr6xw9ILKAmfWIgOZ
UpYB2THa/mT6BqZCg4IeEoKEMqQ9a+8ATDs1nK2V4TO8OuhMVxk1X/cA1bz6wLMRwGUtuxJ6LFy3
88ZNT4NcHIKTCYAyThVYRu8aC189XCFc781KGSMuPbem1U2YepoGWiyWARXimWpH4dgoo4v/iONu
LuYF/7rxTg1Oz0qaI9CbIigzt3hulg5hpcX50cHwT1787KkKH70Yv/qWWVLixJbzMAWvhEtxsJNl
mXFn+tA1CZg/r2g2ElY3CZKBKVvf7mvZwLUEgrpGv4FP9SdYcgfQ1/bGkfEWLwe18unsAbLBf1Dz
FJvRybrqTjqvFZRLnyCIPtRVOUcm8eiFtD6cGnhb+1WxZdncyDepxHy9xXWwZFOC5Qtq2R8nNauR
y/sXJHeHuc3eSMOXZxMtp3tUUsLY6ahzFG1l4Z7IEdSUYfamM+Vs9WR1CzDj5CQ9+jp1YnK5jTfO
NbFtsivJOV4XA6RZ//WqtdQQVIK5SwqknsT/X7/es2b2Mwh4Um6vGWHHVM7FOmVvy3ZNq44gwC5p
yxT/KHr4MfMlMxMSRN+NfSx5/NgCLtX1+yLyZhbTXHdtpugPMsmyOXAh2TqsI1lxaCrHYIXvUEQ0
MsHkdgtt99l6Rsjl/ZCiPZVPlpFsEyUGr7TH5y6vT/AAvcm5/kkK2wJUV8CBdAjwu6LU6RaoAI82
pKGVPURU0XnnufuOTqhcYxVXBcmuZNxtT3xSgerPp4e3n9HzTofrKrNQ5yZs7Q06D+0jHspJosg2
Wud9wRgxrbqYi017XGoO5VnkU63eP5sEBpC6vkr+4nPUgXqCgn86qdfv+zH3u6GLxDfcWbLcB+G2
GRvTmv4+0xLks5ttOIKPPRPEvMh8cAQTveKujBmwWvbFOdfQLyXfJLJZRqqGAZ9ubjvgknoc40Si
tmVrOE/a9wCrZFqkLOeq04v2UkgFq2HRq36pfV7xWq1u6Y/AJf5DACJqCp5RR9vIgTQbvECLZiPX
8XFdxnnWT+VDtevTgSMt+6yF8icP+JQEM0oEiSAfKInX7ue1Qby9DEjgl4tMARa1MvGF4dxRcLD4
qMH0ydmoIIqMdxZxBCVuY3zj0Inb7e3AcX2LrtX7ER+MFgjrk7sDO+v7Ldh6mjK5+ElUQ398rsbZ
pI4ckdYHGk/UGnBDUTFCk9TEjadP22hBeMQ+z9UNS8nidXDvy415AdyWQa+7GE9L034oCBH2l9IA
nEcbPZ3zxjtTwdY5rRR1HBUeqB24pUAaAnyGOFmxtenkMv4iWieKvviwHt2V3A05JdzMNEm2n3Sb
dl374EfrEXg7xTpg++2IFHSfBBz7LdEJsiBnpiD2GsntuPFnWCWKFQWeYfTlfTwQyCJsfkJFOxIg
PbCROo4AN7FnmbEM8R4okVL0h/zL3YhNA3DhAzDPg3+MV/ZP5/sPTcyGvhAzYENHty84VuAkR46N
X1Bi6ItI7nnsJous98X1vyyx2wwF6G1aoxT2nohKPggoI6Tsg+8oTAy8oRU+pei9+ddh9/iZMyqz
SFX/zaXEJMeYZq3AwE1UzClWp/z5R9juordlGmwZhiSiAgQl2eRjW6yGYKIQcS9SbZ4Ih2oiXVym
t9rAsNeeNzZ/oW72SqwDcIKWfBloXeDI5MrGon9o8RgXzb6amGFHwT6SmTlTtLxsIiQiO7ZbaivP
+h7xZ3FNyZ3bFGR7P1IIxo83aNjGpoDSE1SoI4JQKRQ4D3AMloFOmAcyYMhpVqLFZEdBYgVHDXe2
viLL5CwtLMQi7FZxFdQ27x3eCxeVLjOyXIEgakjvQaOfDWa0lijGoYLIct2On3aEsNys3huUc/1c
ZAuGYVfgAx4FGS3Zoq2kfsVcOxeH7mN2XmypW/YCDg+wrQ7zAPhtRKnaOJB1R+znOVfabwJhVSov
vHxpL7FKpqPj+Asn/0PZ1WJ/9P0zE/5na+w0nOoDyr0YQ+XHD8p3nOFC7vqkaTRP/seKRiLWlTIC
SaooTZtbdEkiHX66caUPcnQlpdN12RKs/X/bDsBS4MzNN9Nr7qcfGsAoeHNwDSHuVqNDVZTX7vCV
HzxVVk/VVlBDckPVZgW3GCpabcZtcbbtncvOgSTRzGnMDHY/8OblPDWCv2k3DzEVv8u0QOqGbjsP
tXeylDVmyb5XY4NEP+tovgycWqGnDVUkHP3w41fZjr3Bq8+CEKNeOgqgtawLmgSglA2Wv1WoSiGw
mjwPRW3bCacas0/1LiupE3jfGC/E8+Eqc2TlDKC6ur2DxT2EpraoW6/rpGhWBPjHnu3GSSKUgnYf
UepzLz/0VkZSx447KPDduh2KFMRyIpvnJrwYKl0oO3LjjXAmoiu8oWWRwXJSwZhJ0fx+fujAy6hm
mucvKrFtvRQ+RE9mxF/h8HQ100m6Qt0rfoQ1ES2ky9gf8O3lvTzlmLtcIOuwACP1CQi66a5yw8Uk
CUiz1LP2KdM6h01bGTGk91EVTGArHcHxmy43WQv5XDSwpzPqq91GJbJF3+/c7H5K7E5mHpJ0KMGc
Ja9W6XdJ7VYKEBeJ4xn5b8yqQhiBBpzsC2Zf+oDUQ9qXwUItfLjPyZGTLQ+SbPoL4BzITz7P1fWq
bcU4Vj1yQPDlyjYvTMtBTRPMm/UbIrb0gLgxLA2FgJdsB0xT0a3EkasPg2s/CXtWg8FKUqY1VHfr
p5c45PZjua9nukcGvI2budULxzltoRPdzoaUOi+bCwgHFzw7tspQCHLeutzPoUlaLBX8L+Zb6r6s
6HemKBHjkcXqQrZZBFTA05Rz1YlLj50umD0tBMU1FEz8SertQpNSmnUh65EEtAFTkp97cW+mSqJG
0Ne5h+BRskRaH1MJrNCrwNkoTnuMngKV8760knEE4CryIwyHt2V7Uw/h898ppgauO5Dpn+mgA0To
1w0LjjhHR/cQ4Lg+m8tAXDsbUAHRcWRe6fNOdV/hKukMoSCMphwoEgzfPljDj5jA3nXHzqj1iHf8
7Jvcsl41U2mRFU8PMxSF+qydBsxRJnne7aPOowVK1LV8RGxSF7WMRPBPVj/ArLfwHVm+6ZwdqJuz
+UU8QhWKrU1aEP3HX9yEBVb70UgoPcsy9Xe7P/37Er2G4wSXxYNsyQaakG4uwcljU5b3EaO1LfjI
0cMzRRQRU1tvYw6bGmQJA+CUmxnhomm6xSLHEdV6gN/SsmXyhvcPbWZq3a0TRtzOhC82STyKhaf6
V/hyOrt+6mDxbwzRJnSYE2+aemzx3MS1r/a0seF5Gjo0uqWBh/xP68d3vWBw6KFF1GeySb7CGK0F
A1fitD6gKvOQLWWLlU7gCdyKQtQF49o74C4enndr4mhVy1q3xVtom5PzghTMQCeuwqPp7226MWRn
nIpwKwPWm80eH3YZl1wvWJTEO++8tK2nSpyQcRf73d/lSdXVzMySif9Gm/gfbZ76V/DE0xGCQpN3
s9cuhizvd+xmW9wmllLy1MMlhdM7fNoqhDvBDGAQyASWH2OaCJlX1K1Pm+MVLPo/uyRfJrtOYgnF
uV2/kPEWf4vV9tUABNxW1M+MOkikeuDvuj4HX1zDIr7dTG6KgH4csA3V68SzUwr3Fhqq03tET/Py
fexBM0Gw+JDJRDZ+1x6xjUN+pjPWJc3LRU5QujJ2zswkaDehedeCm2skw3cKkJ70IaYKiy5a6Dq3
mBSOeZGTm3EgsbhVX8REzhvyQYllCuS9Wg3hjbZM/+HCrS+w0gdo0AA0YUqlEqHm/1ebFVJ19EMP
fnRI9HSNF+wkFbxkhbnBSu1WLyua1WykvZgo6RCB8LRUpBiH/DZ+FHKRm/HnTHLCYGWBkYeoLx9L
YDxT/sh+rASjWI1iBTp3nzYVsTOxVsvbu+ZY0K07jTSUcnnvtg56Fv9INFFeT6TDndvomo128H00
kwtnnX+5gAMx7wsEmeomctRjGpFO7mn/NuemLBe3aTwKfDD2uTy06nUvj5+OCacybcMz43gBB+HK
1urS5eDDd5mHMmv0pPioUj/cDwboYb/HtO0LJ1SUR7DTnvM22SbVTW1nY/R439/6sSW6I9AzLSgr
hFz9YWEguR3Pn/rR/uHw1TaArAT5dlm7vKrcu4sO0k7a/TlzQQPWmfceUj/phn7vNY/fQXFC4b6O
eLhFpMUb/QtbqntDU+ZWnAngzRKAM7cBS285V5Fz5cop46LRtXcUjstK8+aeH0oprWSbTnNAjOXD
c/wjyrC6bxAEK2NXBuPuVfzUSYH3kp9lVivPvcB1s+nWy/Rp0VgWvRu8CfLSYC4Mp/q1vOmCFcR5
N29WBCER/DpYKzELqDCIuvTYTD1+OigszZCSwpbIQ8B5GOlAUB0GC2ZtrVMhDAjZTnuMp4cHEr22
/iJkZLh7OI/iM/J0Ey1mNJ/1wqx+7on1HDnK6EUOm1sc1e+x4x1bohf6i1iuGWDpP6itEwFz0O0r
Cc+nDbcWT3Ft519XxlFDFHFVgr4Rgn6gOZHNuSk9dXCokeuH2KDen6EVH8eCnEztybOuqu1xsg3r
3w4uwUpotS7As3v3dWcVlXgFGK0tAEDz4sKSG7e5oj82ob2KXSH2Ax8fzBNOz9ok6O33bwCyLde3
7hWymOCHoXmO++MuW/qEkhHX1hupiWND77duP9rwMmp1aV9uuJ2xa86suGHJCILEC0INVt3PZ7t9
PjYgPgcu2vjXQTTYvloj6tOyixAzbKz6Nefbtelw9CH5egiOMzk+Sdky6pycwk50IvBSq4tIqgJH
+ib6d1OQsGuEwecizRPOE+fzvYrtMS0bamSOa7d2HigcilTF3cb6qboEtZLXqhFyCDRHhkTJ/PJr
WeVruPqFePsOOYX1l8WHrLVw6FeaN4aHFUpviRMIJx4y4U9JjNX4FeDtrtpT0H7BdQE/MJ5MqBMl
Rpzw7leFkKmTb8F1sUYYTKRXSSL0CG8OY0AZATnFXBh9WynWqQokQ7hdsempLaZqCE8jIFJEsyO7
pPM/AjX/kKuZ0GS6B7+uqh9zll4sur+Yh1kdy7g3Cq49760ksJxynHXhsabdkr+atO5botzVTJ1E
Ih9WLWQ//y+zghZzkuwM9k1YMqjR9bOEcsiCYpJKdfekKwmESvU2tf27Fk6Hm2/6NgGXFrtLxp8p
BKXnoo7u/KeLDiHoLCFob/5FXFgR5TMHDKT8NHPI+4rIypluOrmnJsMvhQw3/4XHxShXsKSrpyyE
ndCUENN+371spneOMNMLu/jUm/BoQLhb6vaVEkEEpycsZyz6FuQ08KBYXNWkT45A3Ob7NgsQ3oih
HWpyjFTMCNv9zymAnKFjiBIcevFTD/aOFP3y6CgECd6kxOQctXNJVHOLmG6kgK6ISz+3AE12JNDR
1UlQAPeftQ7zz0e7Y1w3lUldo21D/7EBOXunOL5nlzg+F3jny+YDnB12h64jz8YlFp6eF8pN71eK
JbjoREAm6Ydyzigk4dBjvOCfppYPKAoWQuMr3Hr08T0PenkmoKmMb6LIgAS5Se/IOw8ZzwUUCpgg
MDpZHBSXjYmDtxLJS5B2+EuhSSOdHQdalQx1D2BCpA/gGMj4MblrOEgw2LUmD2MbSwohzjRPXjGR
Ft+BsUBtM7o5TYRhrTrjc5mYNKPu0sBb3moViuG6pR3jxovWouz53PYk3+PET/W20CBbgmZRVr2M
m5jZDkOILBKH33DwloVb1UldgjeExjkyB6m2Hg/vuAnGNXGHsV6duNe+LgS1TM1w8xl0tFddcnkp
aRSjOTDbqDiov5CVQ+BxJP3L2MCJf+Yb7JDIOXuRy1rRbgtEbm91ypoK2d6Sm8Q4RP/eT+8V8PQR
MsUcSBzJccdibHR1VJa4lDAMdSt5CEjraD+0jal9Gx1aXaF6nikmuSaL2aZNizVTkWj9KWltXGlL
fZw5QH3qcgUHxEI2XHlKIMfy48UJNw9pOqq/yykLchteryex4DJXaahymLoyXS1bX0vAN86ddy5L
NecFh9nfQCHT9FCRm2YsF0llY5BJXlLuO9ieR3eIhX3WAQmuUgtdgABzsU0aHdR2aoBvrgccXCbt
O5Tpilwh5pCBrLRoAOwau4yCya/Jwe+JHIgV0IGbPO8UNEUe6Cb3T8yRRIL8nos7D4PtJqwif5o8
FKCH/Cu7aPuwKF4kGYMcFptxNh2Na0qbdtzBMl7sr5pbyMV0vScCqzxKdGMwqWLId2np6+PYA685
kwOFbsoPXynIB9sBzeAcpWQs+DhFY2nj2jteHgae24rkFUmIjhf7/y6huwFBia0xD6OATASKIHba
PHw3jWMcAKd4aT9vJwuExw2I48o+2+a/gX1OdB7NDEt6yzF/NpETEcXZhm7GWbuhjIAQBiSNUA7m
35KDXvyBZ5mcKCCkTwpxVPeFOo3U8zKw5Tlt8/T4dF9CibQpRlPwG+xTZKfY+MWXCY+RgnEv/uzH
ruG2svA48mDnmobfuK1OIKxdE8w7igMiZBQ8uxbJve9JJ2EFTDAXkrAHvb3/qmHptKw8zDUXwu0K
yuvTqnIGdWNDwpYsJHteTB/Gd3o0jiEaxY/yCGyY+9GbOvpHYZ3MurkSF5cKF6myo4FltD9aejXI
wUGwnher4Ay7akpHPoIxCbJ7QHbfCcLsJK8kITfMove4YhpWU9pjElP1Wq+zTWZQibgyupPGxAYF
Br3NvR0V+MKZMvBLtQrIGj3NM1YTFik40ye48ywt1qQa1oMF5fZTQPty5W5kNgLB+SptDzZhJWve
v2loelfgC6J7oBz4xNB40Lsq3OMCXDrjUmIqEc8g6y7Le03K2uDHBSDhrL88M7/45iJWgTRGHN+3
l+znS+iowL6K2J+y+A8xprk1pfUNSycguwYdDUqe6rPL9Jy2UHEaX7HORVpjDnqWx60eoKZRmKWl
g+mLoeZbGD1U1AUAQ67mLKp+ejWdECoh5jyqUjbilHV+Oiv4egq2Hmd5VAn5qQoOHXxGcyfUWMc7
n8n5maIFDqOaOABRqz6VDufRvOXV/KeUSvgdJ9uhPgqP9wrMC765Zv61fV0DU4nCCRNc1k62vOhD
uFiK5AF3WdxEN12thYaJfGuXEzALHovO6oeNjM/0AmxZvGN9OTaRpnKVwA/iuBKYYP4kRrqrOL0W
ua9ibpEmO/rpRDqw8LOyY3PMuRKQayFFu/AOP0yITXtnU/AgAdCU3pV0RBxWg8N/M3wr7OZbHA6U
aq58sF7LoVF9CCTPxl6MTkBCuDWhbjj8GKzsylbiD/vyZxF0vmb7iMDE/qwYzcPz194+cRJA7Kzs
tdsfVJbA9nQSz2KFAk4ZmpqHErc4fgS5t8Vn85su0m+N3W76PKtuPvDsZottCNn9lzNzpAgcKC+E
3Frd0DjlvyhjpjHBDG2/ap7Ya6VSlfauUzFjQfYKPPIOWXkiPxgLZALI/ExQa8TIpsKhdUW5KyWX
toJTdA6JtLaTUwwiJLC4UlgN3f9C0PGfWQjni12AD+CggegygFE2weRor393l25ZagDBQ3mTGFyQ
sc1dSXE8g8L83vHvbr5oBLG42OQ2BjXJxElvUlZQOVrUqFP+DN+IMIgnNvV7s5n1X67shdunpmra
rswMnrj78Lg4kGoiumhX9MW23bKCXnwHymyIvNgo/8S17lQdXK+euCvq/zzMUZ0WZig2Wo920UH9
2kRcZBTtsmY807hyuPIjNfSHaBvXOkNp1gqCm3E1EJRhN3MvIs3BJrBdzUaPB8OMnnNZedtLdVma
cp3ycePLIGjYt8I5YarAJuIhweda1jYxv1fUemkrqYieH1rK+9A6q2cbVtHHgInym5cx2bw655BF
Kulc2azIKJKTYXlZujeiGK17kzSjhyp3yBkL9aTVQ1hKCeA34XS3USchs9qVx8FKil6AhVPbNO6D
XWuKIO/BmkiI6WM5OxWYO8fB8w2TYPIPc/4Coo9VdNQRh9OkcXlgFED6dqm2axmKW/kht1sSBlFO
pMdsQ5QcE1FPJMF8iZsj4Ty8Cig0lsREDib1oCud7fyLAxfaO/ovznHqwogQQ6s8YLWE6fUfsCze
rqm2G3YHri8Tb4AlePNRpI11sEPF7kLEmVOQcQ4G4KiNi2rjmXTK+981ZrgCx8hXR3+r12ExYGoS
BExUXOb3bAeynpTNTYxwW2Rj9bLMGnIM5yhrOaBZVeZdZsg5UlGjcXWmjWn6Xm9f/ud+Nn0lIPW+
4915MDSW0dsjfEEClBy4wELs5TuCrUu3/ZqF7n/I/9vjjUFZKk+uKxh+VkELeT7bOdcgMFLNvxIE
cMeWrjFYEbF99xKStBWRlFY6veD/1jYZlk5eiJQ3EQcXHKeQ3NiBLXRjzpMGZ6VCUSykJC5+vYyV
EN21Jg4MGKQ5fX2i+VZLZsxrptREc8/rmPgsIsK3syl/cuOc7FUCuNFad6l6HkJWChtcHzwUj2yW
TCMtQtDOxWI9kpEt/TMl8yzoZbYnha7zW9KSyvvaC8suxdnuu53aNagwGfxGVElhXjqT7uTbaFgo
yOb3OQbKwg4h9pHKIGluiEbdUx4XbvdFbX/Wn8XvbUAIpRi+EUYw/T0tyw2wmEp9n7BgHp16Pubb
7ukf0be4is1sGvX50cg5Ic4mHRKqyrrNIMwy5hu3PHV9NMZYwb5fdORczF+uuX1eegpoE6W7tmwH
ehWuS6dLp2RXyPTEQnAQM0l0RmOatL93K72nPiC/O4ew9BgTdlxyt9PPuniEKMZNJCq5gV2hETHX
BN6haBsCh5spxIEbMJrqjHevxJU6PCzgKao4QySHAqYq4NnenpQ3S2LO6yJh/PZGlpa532G38Ted
lRSkzP1PZ7fDsOM5wL6e20DmzUDlWopkg78NZqBa9ZiVrRWGEAgFbIfV4V2RYFS4FqVTt48H9l4Y
w13ykLW19U7kWvQ7N2FADWSVWJMdCeLfnF99HH5Hiz+F7ZXw9StK3xG9GuEghyMxWTX0wzpdL9J8
zlBb75rcomQQv8JLyAArgnwV+omW1zUUlQEkF5nO5G/TE2wiZR31CB8Qjr0pd/L4p+rh2KNsaKgS
LFeGJyT6aVbOkGmLp1YnXvOO/9oWEbDhvCBZ+PgaImLCujiPBcBCrpkGAaVJ2jzCzJ8fHVoBbMHI
p5IRjbi+E6TDrI0NXRwrUOXTzTAw5rF7pTnFJzJPQoxaNcZYPeYKfcQY+XDvIgpO2Y+5x5MNU3tE
C4cN6QmyuI1HUPN+TxyYO7WvvzcSjCGy6BQw9fO/LIcQVwzZDtbeH9+kwo0dQMkt+IlF7GviSS+l
pTrBdBkfAYzKIkUepEN+rPb1N0NJeMeKgmWOjuulB03wMFT3LXD4ZsYUqZTrD6KWo7VmnhqLMkE/
tSxxUWHbeYsiTCoGI8woLL6TYdveG5N/trJO4ChqqdlO8X4AcQqRxKhzoWuZxxyk6+rAsaZjj813
Lv2HnUlL8UZnNWiOA4qQylDM2bFFpHpdwOE1uXpMeX1DtYmAZQ6q1K8mNAUKLBftf8gWdcVQBm7t
8c7TEaBknbt9dO16pOT797INAzhYV7MCDNPEGYJScCd0bdG3BwZDVXprAe6eT/kwU2MTCGbzxuLC
3iUenuXv3UkmOJkkrUsEjt1xYJW1RLRyxEjhL85bycJCwfPSZLU4QtsTYrwNEUuymTPq+VYrGeG9
hbZs+NlovBBBzHqm79Coozns/Zr36PStkZXvDncw4aH8HNFhPDK2na6I+ee2RLRkAYfmAltd5VxZ
8JzKRRR8qShg7xnwSIIkUkLLPnrqqL7P1hsS48InvxUr7+w6ITUFjBNg4RviZcyop/XhiEC6z3Rr
czgbKr9X6X0k5Ibm5FzeqCIydvReCe76ImQ72SgUdVCSzcTfDQvVMewt8tckBj0dZCmdsycM+P/P
tq1AgUSx7Gv6hdIEyhlaIt8sMwzdaWG1O2pg74nd/qqKBRLBY8PAalCWaTL76zd74FRZOy+UloET
93nv0jKueguB70Vyk7j3JKXOCStuLKKeKPxtZmp9KREaxXA08PIxSQgD8iJ7pSaHoAZMQmBNpJTX
6T6MKvPgMKBbXWzafP/7aK2Q3HItxkMD1l1ANppsHvP7Vblt3K8vNaoK/8iZvSwr5JLzxO82byMI
hRbzCR9F+a56MiG5AbChI1eFT1i8S8Ziq4+YHjVa2HAHI2SLGwUdRelt1+ijDmKoySO/QwjbEoAC
Vffmw4KsQVCpy6Mg/vqEHjY/jHO1AESW0O49UC+ThF2Is04zMhUFlUjA4B6pxwp4oqbHGQFWY2Ff
/Nkx5K+ZNqmCVSRffoQNP+SdIZrCnt+mUDg9hdR70Ga6hRXhqw7XLvxMZw1ht5U4akxaKIEAUqDx
GSv8qWEwjxVP7hbGlxP81pRXPn85C2xzwyh19WdWRTfB+20EkX+nbRfmorb+Y+0lwJYKcWa8/erp
BEkvAobvydrEAsDtWR04HY+BALkGbEk3HfPYWMwZmAABGe45AVEpUXac8g1Xip7o06CNZcAk7eWz
0jsytPIzl/V8GOrqKXoBVNWitmq8ivnEfOnGslStoNEN++16iE1RTEcS3vbw/EfPAj2nzUX0/gXF
VYNDInydOjKnJXTFJSCnyzJLgNGRz2u4z1nYvax/4H71wRcoO/Drv35a2bzZ8ve9uvJ+kkaDFidj
kl+A5W8ZgzOdnxBeGchWbs0vhfZ2AxDA/HLceT3I3wYc6W+hGkTUaPiMxTOuWJDy0XdBXrFc2Pxk
KpXpmPqYdaEJPp6bUzXWXSD2MUn6gn17bxZS0XUY4nGSgfNW5Abc/Z40xBSK6nXqcnasUHhu2RH1
XgrndcCHO/ZgBu4ANyowd8i9sss2Bqz3Llh9ZvaB6MlMXopZvsgZHuK82HzSBxTUbpYu2om7LdXi
TRDT1u4oQNhAMNatLNJSWTkVOx18HU+hKhC6nZoNaM6M1GjLaw+5YmWuot2mRjSBT1Icl7gYBPz1
NkJyPDtjtypFISmGhyu8obWcXTsbDM1JDxD3KrffiY1K6rCeOoBct8mog9T+fOZIJnv8aCXSH6Gt
sxfO3mnRwn0gfTeP8r+HPIBfMIXUkFIDrDJxx/WbIlF8LKVJG8/T5iDkFKIvTbBkp33H4kbf4dHc
sX8uWPGfxpd8MU8q+cyVprGxBO1aepZw7NNYNzsmQ0hWA5Et6Lw1KAsiEyBJHWpT1P1ng4hxqoZv
0dU2nVBJRWJ+26cyTIjJULUhkVGFm6+qrtMH8Z06MuyxWX8Vmu0aPlaMwPRafo6kKFUQ3GDDkG6f
ue44o13NtWdWSIDeW2tVifXw1K8takOViiW4TCpDMxfBdI8Uk+PSGz6askUyYPzaoEUK+xp/i/G9
juEamgJXBDY1tIx7T4FgduLWrmXsxzsz9auRJgDQfYmnfADMy6WDs9/5VFlHHYTFCQ0VIToNmt1/
eebKU0YRhYFxv9oKDES3zJzxoE9xL93bLok9zWRXRlEupZ6ndLvAVhkSOwbyLV0Q0NfWP4MgNKY5
+nVV6efZDicmQ961spjn/Q6z8wj3His5dwzruL/c8PI1hLh0r8MC0nd/rA8nC+qIOqJOkvizaqKi
vkWzs54FW1dI1kXTPJgA76pxI5mPFqw3FsmKvRc6tdXIYZKLwIQQAVvc7YmQAQlTdm8YYD+s2wzD
ZQLS1UOUHYZj0r/eTIInfmD0gg43+k8mJ7nVaoQsyg1WfTgKWuMMorgknZbrvVzCoeOHwpCrqocg
NuWhKKJ8nPvEtJrsZEMi9x4RJ/G/aTkTn4sffxhZbC0bRjKCbOlqufhBw/KXf7/fi4usR8jnwRyH
QRu8EwEp7F8U4FI2SNXBwqdoQgOolnnflYgaBZ8Av6hQEObmdOuU6zQfr7RX+lL2tnbStHeRPQd+
wBS2okooois/qNSh4YGM/w+KDiZGMl/IG4UHz/vILHXI3SJI6JG+i7BD5oetys2VHCKCvHcsQ/cH
ZVANcJxhxX26FK9YW+kLOREY/185OE17gLguyV105pd7wJBUzbA9kPDkLcHgXCJSQaBzJcBTHjQf
5XHZRv2y59JH35noW9KGskLjI+qjHiptOYk4zOq54L4soI+dFV4m21GYNxVbD/SKhpJzA2sYVfKU
zgCGNHBWOOaWX4aDpULQI0i/OoI/ZtHo/VOJaCHddjTFIzDoeyFkFdNsed2jYjULyyntOImb6m+Y
3PsxPtEU3RSg++uxjN81YCe24cBitGxJXFsYjuIQIgTFQaIC1urmM+9EuHdyNNQ9UsJ7W+gpA0ee
aJoQ3jOzhxVr5ZudP8XxvskkRjcCk9HpCg9ca+aqnqZTXxwdXZbt3rR04TgS8ryQNe5W8Y3Rli03
+OknJdteKdiI4BYVf+Q1cJ2fOpC0gzQ47zaPcckK5xCspdNjJNyK2Bdcv39mOLk522K6ELQfDUza
W9NRiJHFgmUJV3F8UK2YhIhJrUdjHowxhVY+6Ty/4xT74HdLHhl40K2gOrUHgKJcGt4zBSAQhtMV
GxrOmtAaLqZsUQ8d3EPupvk07k0//9ju+BfjomNIbNS1iDbybm/xbWESFkDqrJw4AXR8Lb3+GIDk
s0x82f361193iMXm5DDcv1iSn8CvzUQV4Eb74Ja9Y5sQQIXGJuXIL+O3bAZhZnjD95uJldaWiT44
2gatbwVewTUoIWjtdhQGHm0aQrKVdE+04Wt/h5EA0T0oZKTNC1jNLW9cqab/rCHbpe/4SI1mBUG/
n2cx1bcA0h1m/zEu3sX6x87pXbY0SQMlje9VK61fkak1bhCb8QiWY7dPYNESffRAQrZ0bqDDjZdA
hDuzYxye9bZUsCKpbz/7NN50LCG0KdG5+QdxJ6ftTx0o/HfxQmObwUhTa7x8KUYKSSiI9+u9ZS08
D1cClnBN8lVW3mL8jP5xzUHK/dWLwsVZZr/SCnZ4T/dGTZJjvjGjb6913NSEXh9R5wVECwftZ454
AGlwSQfyfm9aNaFznPyUMsZWn01eZ+QF4XoP4KdCP7oMOv9OyN05/mqTKN3m9BBiy5Y58soMOHCl
T9Am9Ev433ArT4qYYl8ivsHDD+n2F1J5XUxQoz/EVCCdSXKf5/9aBBrmSfBs4uRSJ/GwXXviDTEt
c3toAclPnlo7XYmgPaOhZoPupqzyYJEzyIfpDxWQNfsl8b/A5QzNyxcBPPZKgHn56U183JvMvI5z
GoGSFGvN1tqo65jouwkHXgWSn5h4HRizVGej9irQCUyu8BrJwBSv506lrs7mNzoYnrNDK/7LvPlU
KZn2GimD2bkMa3WbsopJjdAtEOd5m8xhxum62EQni8WPkM1I1Lf9okRPmqasUJL7JQXBHWFJlpFz
UacQM5LVEdUIvO4RMCtY03Q1wSthBGxKNC2+FUcufp6r0WCmQBw0TqxCl4Oil5+7y+AFP8qzBJ0R
Ob8nndBNmx1C2dLCbVJiWpgnMMTiEfUxS1qkbrbLTIg/zGv6xBR2DmxDk3KJztYOIZPheQVwZrBB
crqoZnQVtF1T09+XPvrIjmjZlGqBd3lFKVjChTcgDftZg5bJxvwjwT1lv1MTypQp/PoxyKYr+pIc
bvVg2HMv9fSu9SI9nFSkbLBpMkGI3MvYwFHR8O44bxBrXAbl2xlkf7d/Q4SuIJxaCmw6QbemvXcr
ae1Zb5ulYx+fFBS6RpEhnjxwodl+BaQJvKsVnjqi70bkqT7l/mE/n2v0EYflOJMnFkxHQ5VOYV6O
pmWqXKz+KJtba//y4QXQzKUA6pkxP1KyzZI16OxSUxe0ZBZl6bf2luSz1Qddnen29K72ONVodg0/
ENGaZsQHBK9ozJ1rBoVS/z2KW49SBUQ3uarznOC1EfGsbw1SLK+4bTTA2v8REQ7yw4naLMc0ScFK
9uiRbyB2j2xQ6qpO7dEDVO17gqMQ9m0NHyOAGDlVa5UnQTXqpUeUJh+d13iLBILN+jlQBKF8GRk9
U2qwML0ZIsw/f3vZ3vyFQlh01qqMdK9pgFh2jj2DXIpif5NHdtX/5Ri/rVO8zmHZWTJPvZavudYz
8q2/5SiOQUpU+lQjZE0gWN23wwVXBELIS0bT2njQ/cbHELBWxmgThX/nlJ3+6Y1Ssf6HN7Sadsuw
yhtuJtWg0yVLqq4IUf8LcOaCiUmLOjjS9FEAxzsVg102HtpjpfA3Xa0bTP0/9DN9WJgDIEhmC5lF
rtAq+nvvqLo1yHg9NwC0nemvPd/eHhsn195zKQ/WsP8H5x4xijm+usJ1Wv/UnlVAsHEj5fPTneq3
nqznaz759y8kY3a2vpd7xpYJ3uVksdPeLjWYogo9v8iH8YfcoBduu7Yh8tRnN/UXMISPJYy3QicF
GSTGmmnIRmawpWtwkgSqlYB+BP7r7u59UC1iEq35R/SaV2GGJHdBsPpcZTJMEDtdthmqGW/hsvCi
pUDMFOMBmF5CGVEKQ9mJrtv8WLkGChNNY9Rfqau4rmTQFrWlhX2wcjLq+WBz5MA5O5vGA5RD222U
/fEyXrR7T9W4TzPoW0lLPSsdQHtybFwUrQuu0eXyOgy67YOtWacq3+E+7q5t3RjZUR3SQmI3C1TX
6eRVHdaZF69xJMap+CnUlkSd4eTPBY6tEP6F9tONhTqNtuFJxx6FRWklf31cGUCeM9l0vABwTno6
yjCVZ7v9+mPe/R5DRdluq9EhN6Eg+77TLezsIEGKlEjZnCEW1r1M9g0NY2nQOE2hwLEnb7Pfuxqo
5iOEWc0jHUpyJC5Hjl1weTcMZ8NFw2WPF6VCr0sWkbO8/6ooy2Ji3suaGD/mAt8eMS8vK1x17Si+
8Af1TbNtDoUkqvBjXbiBR+nWa0OIBKrLKAgg9Afir08F+052Yovt6OIzC/wDRqN++JTRGxyyKHFg
fsFkghSRazJU1EnLtaluYVhzEfmEEtXhVbrAPkCsQLDyi9WKkoFUBXGLH5RIUsvu3dA9mVanZkJS
oVYQ9/a+StkC/ONAW4I4PYDo4ExHBG8FrnHKqhX+Go6yDf2s8H3lJUhtmvevQrTqvfpkOCWpO/Ka
iWCJMTnTpqcbBq3xiJa3oeTiJ/fuMGPKTwg2MIOTj/eDRmcwTlBqNQQJdf1wkpxKFCpJjNGBWZN0
+J+qzuVuwqNaaGEgDHlgGegxyOTQXB6J/0sXBy8v8ZI5px39KSWDgWm6Od6jz+EsQVeqc4nWV4qV
pHGRvPEHNOZnjm2gYepL1kW0u4vuDf77bPIa5aG5BpQGvbtS++RJ0xOrrus3PQjh6X3myBdZOFb1
sCRW4U/y71H1z3fUuAjQme3jPOIg+tmi5/5U2TgHIEBBBRAYuRp+GKgFZUkGrnbVtP7udGt+piNa
3g46jbuTE1DFHvWjJiG+vYWjMgdoWvgLqNGDMC8PTfNcLB1gFBLX81gtdANahW/QM3hcecoEJTHA
uCiG3YSqxi9+q/GyRmGHbNkCUN83XxiGZMhh91LfjjwP3YtL6rFK425vZNJp5SRZiKkp1C/xzsGN
4gpGnttStzjVgTSqJFpBEw75AQ7uQT9uIxzLB726zIUEoXMqdwgw+qIEsdYiozsLvjx4vbJRiR0x
Imuc/njWo7TTHw+WyRFWQQzjjXcW3GjJlLhMpkbCvR46BTIcPRJI920r3oBLRVnma8ghxlaXA813
PSTl1zI/V++QiyWHFF9wjQCraytWHEAmEGT5EUyBvlOP9L5PPGStiSTMmzSpk+DxQXOK7Wq33jg/
0opSNBSh94FMOTpdw3MGHYlBu+ns+wcdM+QoKAhXq+ILL0YKW+26qOjJj5FLSz8h41uj82eflMGy
8U5qv1Pz6pLy4b6Pwegke6Pp5wyWzA5ji+cvY/HQPNN/ezjZ4K+xs6Chc2BeJIQn++mIg3ihGoQz
bNnfqsJNO5w9EXkFHzDlJY9UeEIO1nPIPvJGNR5O9lIj5Vc/PdGd0A7N1V+A7//UUzmoI6Ou8ESq
nwETtWiwwtesohIjQEbDxmPgBgtvWIbR29AcJNe8cfddvoLuwyqXOyrnMOGgLNXCvAOKFcnR2lyO
u0VHzNVJu1uF4O0bzveaoMqf+T+EQVmZK1lpc40HVrrv82KngVnxcz6d8XrynMlBfqZ2lhgRdsEt
F09bBwa1qOcVpMRuPehmJ1+u0/yzH5BnIBGI5oNL7iBGtMd7IYvmBAzEl2J9QKWaHtWVSIk0RTiU
Gn+F9D/I27Uo585dN3p6mxmhOOquUadLJAERJZ6kBQwZbbLKWZXbRV1dPzatyScMwCEGoRKnLKBv
hcyMzWLm6bQPXZlGA4GsIdhGZVIol65DwlY4Zyb/KtrNxni+Ab1B1C+Y+IiWbp29EhngpXK5i2M7
FMZmvKSv66x/eZv7xui0pxWu6O5k1c5ipqvneG7WDKokrWvb/sGGLQCm8BvK4E/5CYmND/lRqhvX
NzGiXG4p4QWa4ZPvel3CAF+0cNol7ez8ABENllNozEZNU0P/3w+Si7bxuFayVM1cPd0O0en6LY6i
Tgqa8T2Tmm1u0saae+AwWD3jKyN5+Pt3sH/9QaANXwLHLtM2zeXUfHuneCoc1p0LUlq0kD+6JRBa
PXvM1FuDJb9A4RWYQIg+ld2ebCvStZe6SWMgFSi8k/pGNXIyGkyiYRmz0NTARf9Kuv7R++ClC2o9
gH1XDSFna09UU9LVjbg/+y3eCdvGt8W9+SHtLPPXtGdThdydLBQGQ/vEDkD/C3Spm5GXLuTtJSe/
zJz3pMRnMpksP67ulCMXsun/5tj5BH8UfqEVBz1GAPu7+VysAU6Uu/wZ8l/9bdWWktq+5IYroIYo
QD96rrdS/H3Ga2eZHQcxkLzLNeMaRQSu59WzI5f7Mdc1Bvi1/48wu8jBTX0xa6QCT4hVwGJbMyjn
qVVoaYtLcbVsNPbQsh0MRmo8fmkMTjyoS4swIgXTjBxRDT83sR+6Nl3Ef8POFtBkFEDsxeT9/Xjq
oELOh8pBR0f/nY15A0GvarCdfn7dFyFYad07A6psgwLvNgFGBCqBVmaVVPBMlMatyooiLOtjIcHu
ZdO1KuYIkd0vEFyzMb7eWHZMyTbJD5lGQi1npty9eZtg0Y+RqxZxr5+Ae7A6UJt7cxKDQstiflai
VgaOPAnUJsCcvH1ZY/4zNlyL9oNue9AjlLWZM27YNeQVgQMNX5I8ymGUNSUrK8UyaPpZ5rg51cBI
SGFPUcqhGu8ghwqRqd3o9WB+IlMh43uqsKlKbc9XRfH7KM2eZD5VvDn5hyr4nVhd9czoGOvgD0N4
LIGC8aVdhHusredtpZOk00kzrcTB2s2/RZQ8YB6tIKNLAUii6be4oQobQ3ljkG1dc7as1F+BtToD
75iTBHtNsAlqdNndpostiAJbG40QEo1d6ssx+Gr5e6N1kxWLnFiwTjJzlSfYSYwlK8IaxABKScTb
z3XML+1JerYSxAgHEzSYeZhSAo8v8pVvLOQXDSX4oQgG97Ax5y6SiFTirxvLSWK/bIhNUomUYiMu
L2IPK6ur4/khOCM9tpn/tvra9nTygHJAaFdqmFJgf+n5E0KN7lJcNjX3C/3EuvELFbV75l+YoEDP
7VFA1NHU4ox+miLNcnz165Mk4VBt+QeOOI5NXqV3jkTqAao97oZvmUGqiCWep4H1yveLrryKHS8E
ACkMrBsE7pmKNUwzv6fH445OUGw1Hv+vkmchSCy8LlIU5rmOa2yvS/2Rvjkqjrzf4JkD+2ukRSSU
T72kk8RqMsAYt02q24XRg1Ka0zapcyLaF2kWkzl6YZKC/croyU1iGUh70lqmV5wcm+04jgK+/z6i
Zho2+agFO7KB85jldx4KhbWRaFWgZfri+TZWfp0hlulyiBjLBdd432MJ7OYnlSYTgMxz7nvzLlAy
Wd3h8c9c8AdXaOaau6lF6sdvqdvZKLaV3x/JmbpZsd3SQMoszMkujNuSDbX8PV7rj1EFblHY4vDu
CM8rl83+I/VzblhE+TMDQumuKcYYf+1ItIC5RgYMQB/95x5Zhl0zC4DA0UqPGZFNp8ufKZCdYpvV
gsEBLhO3hhzNTbJB/4YEaIb0DW4SuOvxaYkatM3fmDb2uw3ur73oJd/WkE29TLnFKbjna1KRvvgt
4ElEFnVC5px4u57ppVIy3LQ3iAhPi5vJs+Fc3p7B/CGrp3eTcjZmecqIcBs+HZZT2MS522OynUr2
3k8yyitiDdxImAAAJpvQ84oAY9SyKB19WUltx05nfBCSfJAvtgebcbKjQ+++fEGLn9vw4bpoAX9N
l8T8GiS5Vf2CrvvUAgrvqD8PGrdmVYFk/26iHo+fq98fTL5c+gS+pscA1sTOnMYAKUXyknHfjeGu
dd9POn/5LsLGuGGAYb5Y7TRQ63Cjfr8dvN7KnC+J8+ZRTitb/u67zZMGchQ3D7Fz+Ya0sLScjaDR
LGvFV/lz96QwrTQhGNC2/09NXLIHou/2Fa/bpmkvfzoMfyE+y3a4c0axKI1VaYi+2bNhz3vpaSsL
+s2w3JoNbYqEaWEuONMhtcuWp8DaqO49TscPoHEGPkLzAu6Gh0cQwzHLyYwCMcaak1nXfBvBxmmQ
R8cBYOIK4ck+Ya1S0VNPsmt8S/Q57gXF/sTUCTGZuz0oQ2lWsjKgdlcdAOljZFek0uLYRiWAK+YW
OnMlX4GJh3VRIbnOJ3WIh6kshSeaVs50bl4AM4mlPmCRDpXtqb9geOA+8dJKd4ov/Ykd1GTU+ZpP
nutYP9PJYvJc1maLMM0f0u3HiGL8z0a2APmBXl1JCGVeyzyttdCon2Os4ywjtC0hrA3r8i6uqMMQ
87EYScH6a0wxhyX46SF8OsSzvR3tSBFzfa7aShwn8pcRKJ+ARhcQUOncA++aQ3NJn0JD5yWmdb/4
8wTZJPWlLknFjCBK7VY0RZurFZgSN3Oamct7IS1zTROM3+ygiRo+LEGjG7klARvG7z50JjylQnoR
/LWuRI0z7p4LX9UicLdNe4gUreVvm/6yHxb2o/Vxnl7dW8bCcF9WvIJSsknbAgqs0cVz8Q+gMyhc
sF5tLUfoLbBHaCw+t3IAu5J0c8f0qvadnpjdl7zZD/UyWfhJUsN+KOwvy7JqqZVVET/MvW1pf6Yq
cRW8ymhywKEUyka+8db5RckMDhVhw+jSL5aVm6M0UX1DSQsCor3yR1EEplETEblUvKtj2IasCye2
/kOzLCe5J7Fvv4oOiEYtNR3zGQnrg2n+ZGyDoLgCcy9HyVykLHI+riPGdlUwjliYrw1Q9bF4WwBK
9yBqJBEyDaETcW7Stmy41KCWdS1CvfWrmWhgC1oNnVhSYsy2TW7lfstwskHNaXY7a89QutfKp1VX
HnwChM0IeXzSNT4iG2BIfuqeqoaifY5h+V+kd9EgKxr0HOLawJOZgqy7F8XizW4nlwNaepqcNBhr
wPnenB1mlA4BXS9PK5Xmz3fjiS61zDvNCCm6n8fXf69pN8MtmZxoG2dkOHx2tuFAO0G0blLOHWT4
1mMvfc2L/qvchRj7N6ENVZeO316jCZuqK1L0uq2yVUGbDvFAgupm4HWzlQCx6wTgTiIsK/6HlhFl
j/kmWsL7heQOm9mp0601ylIPQVt5Iy29AMoK1n+IGMbzfY9BPshNl9WGQW59Q4kY2/H+683gJU8B
NFhgjU9vvk4hSYGKd5PQZDMGH6RzIF0sfgU3EIRCF9Il5WpTf/G6XjFrJCme4JfaFRItTrGBTsiq
IFqJA0AeuZnhPPMz4vCb5RFGo9vewslWzogwkhrNrtdEuDf1IFmVUyc04/8LgaR0JqW0FLidtbOv
UbxCMFvcjTpO7viE/wvjIFVdX+k7X4ObJ5zxgiLT1CZJoU63meRTJ+YbXtHs1UOS2gl+xmLpqqex
oolSaEgXLZqSkfh97miOZZ6/10RNeE5C+S1Qjg4v7OYlyD0zd4weXedj9rH6wlEv+r4kh7x+X6Eb
e/j8o/X6WsD1Q9fXnn/CyIdNo9fMXtj1BEH4PTFU0yQYadDNzRIqHQzdYEytmZj7kJNrURkB7QUc
sq/W+GTnUzkwrefpFZDXHa9hFkTNo3Wzbv8/eLjNgJjH5tKaDTyBvkFNhdRgGeCBmw9L7nE8poLy
//wZaYpD0UxyvnQp5R2HAZJ6Sz+jIRKtfgyM9WS29BCRClCuJp7aPZb7iInyt+mOULBWZxzFcdiU
ZyvaPsVe9nbvjdgt43IX1q6OIEEDRIcCbKXFaji0N9xyQxMJHTQR/5k/uOvD141MENtgzB+/QvQv
uOKKphcjLOrtnTrUz9Y++/egpSQzJc1utm49tLwYVP2/wkMD8e8S/QHjviLJ1yptuiwwwu3PbE6L
5TxcAwOyhjTb5Djqral/GTwJEbf8UdOOVQpv1GNY6Jc8qxyfao8BpDULA6cOTF3c6exQ/Itbwj6+
xDQWQ4VxEwq65eWfD344nx2zduQZbmBRqT1ohhjnDnA+cx9rnFKstukgujj5feV03H9t8UqNAHYo
q2w9kAH7ydoBtCTYCXlMqqzJB2hcc9g4LCpfoCvMjdFGP6K78zHQZl+QQ6H6u48H9/mLz4/q+5VB
QKHa/uQLziYDHgaM2mc1izMC+/jGKQkf8nwyREyjY9m/HVSJniAs6TN5cOZQ5/mp/XlafoccQbFa
9i8v0Vf5w9wWvZ0NZsuD2bhWFHhvh2TIO1aG/1y40J4KbGVWCvth+y+lD4VEfbY3DUgsGkzS36Ek
mvhPAw7mVQEdqA9RtENJ7cls16FRq73iGEwpXvoagXw/ae7KRuUuArKpexMtc14Biaq9qhC+qfUM
iFdGP5IJ3SWYbCY2QGwWhOnNs8DXI4IBlznS5h1loEBy0oNxrZ1jKDnUKsaDD5udMnZpEVb/+EMJ
jArNGCICt1WMwdOubeurC31mO0ZIc0yu5cUf+2scrJH36gYQBRutT0fPGSI52VGxXOVn5Ij7Ua2T
1+Ta5PApT1vXwGTEJH/FSnj9JHhwghK+odD+7sCKKVqCqEHuZWAqmdjGPrbI2Kh+UHGsu4ItUSj/
FG/lYIV9b5SzOO+e3ivRS6UtlW3V9g8mbOGInOcgPelGu5CXU1elUMK7tswvn5mauFXfMn2KhjyR
ZM05g5ra4zKRg2RU9Xrc8t8fLgtQWUrXXdFou9mQFLq8aIDNxQr7gUbOFB+K4ZNHapd8MJMRd6+s
+60YSAk04GLyFrxOyYhNg3FWGA+zHTON1PKoEx/vG56xibAdXrVK2D5e5wbDUrl83kCbSS2KyFIx
66khT1G3y9vx2dKBuljr+73jc9iteZeLPY9cAxLjZ+2AqDc7RjEVKUttRSPajyEln7igHdT0efEV
KugN5jEqiraZi1wQoMUtSmU0O7USsO/8lEuOp2SsoicWwtpTKdSryobE5RZOl/ILSC/1EPqS04OJ
62mm/4IalyehiI+HJQ5b0BH5dMB/PLXnCkvxNdAFmZZ/7jhIN9oUBFKyiQr8BR4qZ59xxp3qHwla
UQYJTTszjKM1IW5DXfgFBlpfGXpTKqW1SuI0XurlSHhIUEu6n8+8sjGxnDZ618Oej2QLk+mcVv0M
QJN9QGho/SsgXiK7Z/roXBMm+eTf44DJFVekdmRJJAZ5BPrd+uW6KneKLE1Ki1LN2xFnYhMuYKro
OqpGn/3KcEsu/yMggYhGWhMKximPuNPdS5+Ii3lZ1OOFNHOe/i522ewiB7z2O9g9YD/PNHtDw2A+
78Z+1s27wb+5mhRSKfM5d8Oq/bATKMEjWegmDgLbnZMEB+C8JZVRhe58QXW9qq+tnb2NFLUZkki0
kNNf1AZNLNa7cTXAt2XbxCpBylOgCS9Q/lHg/uRdfRvZupHUqKar+gIoLaw+wup+0t77j0DeyJrw
47dlZcQUBQS95rtgKXA7PPd7ml2Kz/E1Rd8ds1nH4WAV+1/kEIFwYd5yEqV4XpYSSWuZG0RR6Xsy
wkz6ZHQQRJBQ3X292KHJfBkO95KMR33KpB9MaorDo4Z7k5Ca11Eo6CNqXqAlbmp9tZUygCRk3Bi0
iariJ1tp3CZOwBJOGkRME5+2iu81uLLMQqpPDx/WUdr8ITgB1j5xQPcHKx0iKPWMt3KvgMMTktMT
dICTYh/bAGVXJhVeZwrY1EXDkLtJlI4BlORC2tvBXpPIJq0xZfmE6x27XEhlzRExdkW91Aqcd6Em
v7YrAFWJOqovAhYoV2cGTf0zPPDvfS1UqN32R49fx51EOZLT0hW+ktQvnZ5ICuJDQ3u5YqvGZRY3
24qzSJTmVMNCrof0xPVDlZZK69u3rU/q6Iq8OpUsoU+fmLH7SO+ctsAURXHXEqocEbPhndr0RM21
PqcJ0MzCvORYfnk46quwV3aBdRO+UsqyA/DZBN4IOmMElQIzL7vwVbqr2bhhjNH9LWKgUZDzmAmg
m5oFBxXkW2pf2DY1g5PfHafPZyafPZZjzUSSqSNpfkDoeZSgyBbw++YP8Bv+TYV4qxfGt0pzKZz1
vhZWqUInBHjAMc/qJzMcNHixgRpgIsimQRwCwuONYHYjRSNpzeVHKiENtwuEd2S/5VL1BylHqj7H
pzjIIsR90MeYM2cu2DguRjStJihIycvn0zFzcV1NfZTKEI1mkQL6vFLszEp207IUW9VGNgbeR1LX
EcT5NtFfNc7wVccf/E3JbiqNJJNMGvwnxxZzWCdCCsBrYwhbLeKn+xNCoezbDYJ8m6yvqfBILNDs
Nss77+HwCzrbR2i14WjBwY33H3+ByqdL6PBHcW/KdHoIB6rzIKhD0p1GzkdhVemvdmvjksSkoNYx
ExIB+o0pkHVAy/bGwag7rt/aZAtiW5ALqtHR0Om54CTqZ6jv7taZix+8WTuoiPoxfeu8wJvDyAvK
sy6tQ2NsPc6yPK4XtBpx2mMs1+5tkdfdjrpP/762K7uz/Ex6HAFCtKZ7FYpZNuniHxnqVec+bDui
o3x17JvmVpazA8P/fuTu929GWAdiOUjPa0Porbp3dudM2fkGR92c3bpstWzRfUqvuHrbdegB6fVM
fwoVW58sZfYAwgEWVJZU7H1X4www14EUN2PVkVON88AKZ29yhyK81MYnDk5t0YU3rSnJ9DI3h++E
WbSls41/DAqPtrEcmMiOBKfWbZEILJWZuN7+vJpIlqESbJldQdLtva+ywKcjunGjDNZGJSCd1LiI
DalXZg1UoiPIiLImhVapO150EhQfCtvO8a1FJiRMuzAkS7cTq/e3CIa8XkI7RJxeTGVexT1JxyC4
BSuwSLGNk6y2XuLGa5H62rmbQNFZZCsp/duC3YwaUkndd+YW+HkadAW1e9uhZwU05YsakmxWIkPD
gHWRi1K8+A3Zhe0bEX5MZZLfPw9iq/9lvxyZqORNpSE5EwcFd+a2zxVE80kPZzi7nxZvugDZFvhn
H3TJ5fbp7FKNAsUs68ZEASaPwtLVzQfI8j5COzE2YTiKgmoPjqLhpsDdAbEwWoFZ+9hF5QqGf5Ll
QFn6yafuRb9aJou3YPWMo0hQS0p4Gtj28dQEKFZZOFqp/Vgi5k6o2izc09ITV7gws/xdEI696Kk4
dr4qX7r03C0H3yAnPxUqGxXLgk5zTFygkKl4b2jhIdT/taJC9TzfdqO9mz6LT9uJIshv1LfsJKDq
9uZlZBsAx8XW1N3PHnI5FGnmUIkqpLidMxmA9EXpwcWmEWa07wuOgNDiR3KtJ3Hcb3nkgtO41z59
elKhslrlMVLU6oaGi5d1POOJmgws5g3BN9MD1uesMwOPBePxOwNtDp9JJDbDokwAy10GBbZxArZ/
fnp5vrgv2xLNHa+bxfJOtgJr/h0PG4Wnz74q5z+663JN8PEHPVcCIoPMpRh1wlJSsA9Ofl8HC34W
LnZpGvQ1i2tPWoTy1l1gwU+K8QRRuEYU9CRGCFs43anjMOzFhZTmhBVn/IPVeRJcwjbLC4DUsOiP
X8Di/MOED/2ecasuARnsw8n1TPnt1GpisNcw/bnMsnBIT95irX+eYVnY8I7vl4RjFHrWMC4xfaWw
bwgeREwoCc4D+70GnJYv8CSgs0mOJ+bgGzrfu+kkzRmNBsiwKhtC+lymp7+BctaLjCVThI7sGaHF
+AkQhsSdOrh+dq/IqtnSaIpYk9Innp2eJCtNMWp7Ur0ZxjSH5rpzQBni+UM/afPR48KBoyqHcHST
+fRDaqZydZs80id38gTPobGfPW2hSoG/Qu93xqWx88qO0M9dCehUkoEhjZZv+TfBOWuIjUYTtV6/
ihU+vB15zkWlZ0FyMocXoSQuRmJBCq+VFwpBK+e7vHc8bYnyZfsiIS/0R8CHBSltcD35Grr3nKEs
czK3aeddg6jxquhUfo39v8S0wuRWklWCfhvoeVjeizhKhDc7XTRgcljzt/hAnVtcbP09akmemjzj
btAvKpogr6SE4syEJfwOuHFLU0KUSD8IbwLCOsgeIy5h2sqEeUCQVFinamZspjcBEeD+u7GTCiYJ
so+9fnYQO4vXkaMKskocp9wUIlqAYwwTnbgiO29rkYjNY4161F/7rtjNtWd+wzk+qECqDJDudyks
0P9aZJjvfF/pD8HUIXINgA6j3RKGa7UvQNcM2LOR9jVYEy9/WuWsT/JHNSHZDXCkzzvsreooeTsY
bAB7h8zWm93PNF1kmPjQ3FSDUpjU24hr2JxnBfQcl73/A1ilBOtRa8D/dtZFih6SNoReCgWQjlJQ
eP4MuYeyZzJAOk5WyjOKESFkzF0GstSeDYARzQNmnqDtKdUPr0l4N2zeQgxuFjEVqZFSb85+I3+4
6KPWjX+vXy/HQSSFdlZq0WCIy9jGM4avxQbT2rdE191Zs3csYaSIvmuZhGjOhC+6N55Tu7mItkGG
9oXAcupPn1M3wx4Rf4XbG5iAXzY9Wyan3lWI8rOGBuM0F6vFoC0oj3tPi34ExwHVgl1LGUc6BWOe
lmZwYImFCurvUeR4r8Wf8scrWBeGncqxy0wUnV7ZY6Ji+EH84gpEKmBuUrqrsttPWZXOnZzw5RPA
cuZQMDKPcX/VAYESNzxgqwoScwHGIn8DnLiDTxGEhIc/xFQPZTSzPDoyqodFfZI8vInuIDn6HA/q
rQ89ep98Mrt88CZEWrTyGVCpbXzQgfH+0xScNlOjTeRKJW8YIXhj8V42AtU0tJE4U9uw7xanKO7y
IEJq80HKCAmxe+Jd7pC0BTaFkwia630r77wP0H4RCFWF+1f7pGkXgCaQt7CMKKqPXvHR5mKbzHHX
YOQ9xMBnjuOXNDRR0M+KQeRuRtdOK6vxMBtb4Oc2p+VoB4CKsvVlHf/twm3D+wkcN6Hyg77L1Wni
C7cw3UKLQgXcevql4Q6qfengxN+Ydgy0gctrBdtJ/XWYyUBaTvzgVxNjGBO/xyffoU2nir1T4vu7
smMwFqdRSNj0+31Bdipa3xO4YkuxdpEPeDr3K0YfcE3VTK90dHcCSeWHW8Q4JP5Dvqp2k3z4lsx/
YoHp77hVPTNUECCTuRT3fWeMBtlhX6SjEBTarfB338zoOYUbffasK1RIk8ZSH752VSJHPdwJ4lDD
+H8yWKeYjONniQ0nM07IjtB2LmOzhJOrBjlrvVQi11K55D/6G6KQJivLpKSYgktrhhhY8P2yyIxK
XodVH6ioZhKxXX+GeCy65rlqpdheSZLm4MLgsJ8fKwRYOE/2LmKOYXFnhVOkKcMfr93c2oHl5ZAr
hzpAE47Q4BvR7jLkeMKfxajR9CKe3uUTCagMe/AjqJr58XhgFcdR0yR1+hOpClzB/MJ4Tz9nBQhi
avAHRosrxfb36JppjW3snEYPP1wrxh4CDbq8jK3erqUkP+YObjuTmbfhVZd3ntlGxvibtFWb/5Vz
Zwl4oqHwqlkV3kAMkPh5j1K1R6EcreEvGivMjKNIRQUUxdXIzQQhmjzie03xEX2nRdYX8HnP5X0i
gDrsSz3k356FKpKmpEKXck1EH6TKnAesNsXE8gzslRx2z+Oh2aeno7pGysm1YWWqsUqCb7fpkFC8
eIBeZT6rZOyalCLR6KTcUxRxlVTKFjxGhZJ9VWoZKwQnVf0sbJFw3N7USpRNqgwYC9yHwQAlL+LC
RIVZjcwz+5Mimbj/IvzbPdwh5gL6sNoeQXLDCmH10XHG+f8Vnww//Maj0hRXNkFJWu4WZuNlQsAw
Hg69LZx1gHpdsQX9y2vdqNuiQ/8c1YhQ/Nbju9mlYc1y/R3FbZzA2oNyDtM1mAvh5cLA7UvSK0CV
tz1ZKBH1DJ2lYAYrGApEWuUBmNtumIrFzovr3BNK2VjNKGxEqKimjGT21saA2gk3xYq5CgGyvCx/
gzbWq2tX0DdwQi5FPuRPZmin9sSjzoJ6xO42YxRdiiu3pb5mCrQgm8wEPdWf+NBhvwj2u2uC9PeI
orgBQyHd7RWNV34izNcMG97UoT2PVmu1aexU14V/n7l6tx6PMK3LJNObOinyvA+GSG9fCscB6Txa
FSNIi5ya3BjE9b+czvsuwXjsLU3B36ITF8tsdCBavQbEOXiiBtVrc+AsjzgnPUIFj410kqVzRQuW
sHfk8xkGY66a/CuyE4qQE5HNJWJKET4rpNC225//LcRWEum2djfoz/hDaCT/rhGu+72QHZW64B29
DVwcLM7tg5Hxr5ACcPlSiqQ+OWcY1+zNS4GdHObHcbLIU/RFZl3xPmTPl/Ka0fUDOH2o+yd3QT0u
tvdGC67Nheq6wMB995U62wPF/hpXbYW8ToCYML3BepCcpohOD/WMi4B0p5BOp9zruJjBLeLW6tEz
EzIQMmfjIKRXyv8tR5D0HnFgVay2qZoIISirJVqilnvVsO51Rj8O6GDQBioBNDsgikY6JMQamcaT
SMD/lawQnZv9W6o/H605WUBlS4QIz7fMweoyx4kFkXR8pgN105pxY8qI0bRkoXiGRTW+Zqd3HgXn
bpgDMLBh6UblMiMXfiHMxd+NYlWUwmiyyBNogt5XA42RQfJQ4pwxvsBPrBPTzGpPyJNNEZdVzuBr
1jIu8euHLx7gP0JimXSDCCIKkhYlPCtBN+HnKnWrMJWqxb8xPnrD54ircGPsyLgwaZBoOi5PYA25
oX4PGu+mmsaCz6NJAQqoQTJQQNWXu9+ZAlLWJ5+0vE+8ye8ICH8krupQdY3t2bU+khY3totIiYrb
LXGbkKqF9+o0W9EED7u9DG1RlevfLVRjWH7oZev+1EpbcaXu4XZahIoOFFCPI0UIyK9q0JrSQEZE
HTuavECxEn4ci2jSaLabHY6bDQXVOrmPvqGosHCuT5MKulpCBStFWs2/7PBdB2Dn6HC1AyiLDnNe
qSvQ5BLm8sekC/oudNymNtLXiZxVJbjiXXUaqCm5sE0a0mJ0pGUlwfn9JoexTfYT9tfJqhUy3R7H
8Io/Epw24AjWg9MaA1p4tHcuiveC5LlnM3rz82l24tYy9Eu89AVleV2kGeroxmqGdOJ38NQ4MTdR
ryh9jzg/MBXM8bY1eba3mz0pGM5nobm9J4Y962iVQCmzVK3IHhR6fwvdrOBSOg2+7Gt7tPp0BUQD
a6Q8hRcvAl5sV05pPPx6NqXrz7yD2+TJZF6xjtvVh5lsL2q7zFIAjL5nYWjY2LzV4sfkFVQ0eIiY
JhwkXmRkvWZyG9DZ2ZGHxNefV/wromivSX1ksOOYtivZDr7VYnCMzkoNU/BlOovp6fXN43aAqITa
IMYxH1f7F1jbTKkYs28AUsxehSz6tMVvhFIuLQaKQRnVZysT+tiBM7ru8NldGW/20dprZG/fBFXt
Tt64NveTLJ6wO8061qy6/VYvDOt1+fhcaDAv3UElme49Ap9rt9oUcXIirZzrjpFI5EmfHefkKwgp
5SD4h4DqfbjI6VogSKmwCGwv0XFzqBHeN4zdanmg4AnZu8Dxc+xDkFY/ZtnfvsoXRz4W+W5/+7V2
DtBVKBu3kDa3Ai7VdjMgcMElt8HUpsGts2wH7iALbZDA9KDlmAq9lIcfUW7OU7RmEsm7QCUwdcFG
vkbf3G3U6QNUXedmZsB+dzbXkc+qBXhRQwMySskX+ttk3lDA7O5k7UtV18E5tIgR6DsppWeTBCCE
P4gzlq5ehqrpVtT4RYJWievVpa+SU/kMiHQU1uyiHs5L9J+z1/TdyLw01U5laVnvM/7fsCs8RMJD
+5FuSs4pHtqbeJTxIRqyRR/aHspv8QgTQSCvc0A8+SKzc/Zdxb0gJSd8prD1XRMCYPK+ma4xctZb
B0HLZoQtxRpB8+7cNbwYBLL+XfybcvThfdJo8n7fQMMukbTVias1hHgGHxFqyS//hKja+iv2YcnQ
vR0OK9poVSaV1s2YL81sEANjPAL4GUegCgAk03e4TP69fMN8B5WTHGncRCqbCpdVGsSOJOVigutz
eeig3pCdiaCnnx4JXj7NKyxVkDxRsXbe3OKgAnY/7EPbQrB1h9xWMAMZHs5V/wYfjeqCSkU3lJ1d
xjRQryUQrdwi4Z9+cimjIrrLPprsqrFXtK4nxpBizU5npaMUR8LEaHHQCpnJcdvjbZ+6y7QthV9V
pUnWxRMhJwcE2dCWaord5p4F/jW38cL6rGnKpYmENr/WTfZXD8JzttJLRB+e/IPRsPc5tssDVAJH
QsHsdeKtKwOykpS2fuVmbiKBbXMxQfDPfFto+hXvcm2U+u9PXcCFCmnNVvFb2UJRIj3FEBhHfcp7
BZ2ETrY8m1go96LVh9fFsLVaBguPVsLofhWaJvkYO98Wn+DxOhyBjrNKDPjTTbgSRcrQnUtPJt2y
L3p5S2mY5NQNwzPTcl2qSwJY6o5zh1tiKZX9Sx7zE+fVNNQecCJ/eoGeUDYaMcsVssgkg4Twk4NY
LbdTNFz1U849VrY1ZJvdjVeDRA2cnFhJMTnsa3nMwLEdiWxIcQU9UwtYRxbnpqFaDHfBv/UMVG9D
aa8USRcLchsti8egWKp6lHjYs+/la69edWSTvON8iFXc5UFFG74sHKL2Aj6Q3Lmfjp9u6tQY6Jr0
Sg3rETZ7wyQfY6E449+fD067hCSV8ECyJY8tkqbslYjvBVMaBNo3fN9VEr2tr3K7sSUAQ4XLC+N5
7ZCuEn1Y4G1CRWM81Y+dB83lAsxUXNqFliNiB3FUbITAJUiFvmUE3P8I5PKANMbme7B7hD0+U44w
SJBuaSzwC/YcxN/XNyU1DqajdOh5/GSU1Nfdj4OPJ8AXudV2HNRpsYBHrdJVNSArRy0JtAcf7FYK
ofJWL6p5kGGDKsq+HEbAG0mbk9ZIHNw1Jczt86sWUKtoXfXHsMhI2y2Fm9pFUscwBsdrA+9tBgZB
gazvrzfVCi4DUTFTr8J0fLivqFHnX7f/tBtDICrQerzjW8c0TnaIXHGcNha5J4N2tT0SVQIjYyNZ
kAyWs2nLW4zh19rBCc6c7of7T5rirpNqrvyrWrWBSV/EVZxpJhh6RquRtYm/kO1ILGh0+4x9wuuh
VnDgCDUhgYa/ANI7w98jyeTNHOe23IUAD0opMfSrlfirY6slUqWBpt5a52QQsXTJTJB14XQxNaEz
2AEotpWV4Oo43UkaAKPz1RRGQhtJwxQ/5AwK/WFiDKdouLVN/QDq6KL+NMIXMJkGgA4cU8Rghwm4
V//QbP87zY0CYGQaIQyETCXZnV/ykqqqmuP8B8FTUokgvnXWWEW2i6p/JUKOVZqYqTZwj2MVUWr3
cae5TcxoTmraLlC8wWp67Bx+E/AMWRgVwGipdOTnv8o6UX40JKre58ZD8oXSlEcR+021901dsICQ
4W1s+fSnNMA7iKjy6o2xpOPhzEj1s4FURx0NIbJGOpDhKAMGFXxTHkwaXye+VZq2ZK2odI54Bxc/
2Q5GFfvS2Z61f77VkzbTjIlH2e6QHRFpJocmJNZ86POfIjQ38d5yhCqwR4q6rgiod2U+bbSZCyKr
fjqCibOlQm1Y0AbgKI3hEWMdas8v3izGGQqEqEA+urw4YlDhuXlMzxa9Sw0qP+KGRh6am5tc7hTR
+Cd64yVc8duhEmv6WmgPDh9k2JgSEBokmBdWArhGx/f4FR+2YdR8WJXEEshph7ePW/uBXytsrKMM
zFz07Gwmnv3hny2v7xvqq4ZYZIFgDehATJE4N6bmo7Xy8j57V4dXG1HtC8SQcD6JwJHAxXTN8Pwz
CngqgnSmsxPkczqEqYGhvt7RutZ4myFBRAR8HNmrjjHirm4rpi3MPa1zaA9h80+uJiRhnHgmIUi9
PJgtB1pH/tV5QS/MVVvDYckgdDkqNdJTU3dKql5PwqaVRq6LnfAlnjyPfWZvx4xko9DZ+DagjfL9
CsoRbBjMdNOHbHxZ1+rT8B8fP5OC9gjP9k0X35WUd7iviV9AELYZ2/eE1ibNyuhIvCthsnUmjOgj
weeXTluosiidPI8w4ASMpTgoMLcRliRSBmgK1s6wOD09Fj1sMWksrvGtLjQiUxMZuLJrH63a5xMt
ODHYiXbad0D2t/gUGQklpvw8J3KBl/Bv1B7I37gLRk+kzMq3J/w0+eukxK3xbMQsttDG42jolWwc
/LL4Qw14pdbpVKrKTmrSnrIZ94Vx28mx8nK43t1PM9weqtDYNzZrpJh9PPE6l5s+77zaIL1rzRHU
GugfFt2fVAO/4DfyI6sMCX7xQX782yqUvAhXwN2O4L0+m9f4eAJ3Yti1T2l1+EGEdx1dWDQIDVIL
pdiuUUYwF9yHK9ucVhYkmf/rrMY05KBvPS+C1z89vMHzPTokvFPZET6ONxiDx+ihdNatl/ZXj72l
BjOFvQo04vm+pke5nqm0mN7qU2DzHEa/jFUkmTfHqScIHUjTn0/9pEWOzQHvReHfvYSm1iBnYLdY
4iwwOvxztk42NbIgEw0htb3zIOo9YyJTtYtqGfGrluTpYvjncA5BzzoGs4Sei+vVNwdLvZ6TJ+as
l3H9TaO085iDy+atjnrg95Y3pQWQaETsccnrbpUKBYZD43q5RQtEbzGSzn0iprXJvilyjVaSMigS
LQvOGBdflukuQ4lW5A+wPcfxKAlCBsGFI4ILVcdNlRl8yWF8xHKlNXrBPZUNZLqIdxhrQPkvZmD+
TdSX+ImZPc0ZKCwbvHC585jxl7P0rGcGYkoYUPaM38jZSDRgHIIfzFoCflVti4imNMsKMwzY1wXD
raBLqYeBI8JiSkUhD49Zj101BNEYS4vlSdZUY0aLBii7Dc3UWOcQAF2FIvjzUXF8N3vKk3Kc/b5J
oLK1UyAQqPhT2jgnf0LWHRNb1Sg+8hWAYTgewuy6YOGjwS7PtkyUGhxL6CskcaZIYC3RNp1fZuA8
0DY+HsN2GTHNaDldIb/0jov0X0j10u9qXf+dETNngzHPwuwthB/fS7ktYtk4hFigb3uKa2ttwS2/
sBjr5aFvXLTLmJS1Pc73ZdnDxOtM1WxmaUIy4FRJCXoCAru2j+8XSMT2KLoW0s+O8qNf0qYYn7Sq
LCdNBFWCSqrmex0DA4iAB420Qkq1lQXnyYeYly9lKIFbAghwIP1sZZcB+cLfn0ybHlfo9b6138bi
0QQYMwEDfiuaTUlmzuAE7lCHgiQhV+CrC3ZEbfQVhOFWy+OSXuGjyhs7eQsPK25ZHAgLC4Vl2Rrn
krBy/Mgl3JQRm89X9KU39q8V1A9F8DMrouFZKjYs9d2bqmwwupwXI0jY52HPXidbinYV72seBW+s
VQ8DqfXrRDOy+3eVwt5gU0UbmDZLTEFayAAw66x+8ENtnz/WDx2iG7Ew/kXRIA8R2XiR44Hcsd23
KTxrboMxRMfznRsfBYpvMMqP0Y2BR3fqMNgNwKE4U+IJ5XSIe5zngRiZkxrDngoPwWDsGy9wBtZ9
6r03Pc9m1naWjSWr2Bv83lOghW+NZHwh/CZWG0NMFUyemA+P38p8pohuh3id9yaCI8X19eYPIn3U
vew2DrtvzQ++cSa8v0b84dpzYipa0Sh84aDp0qJLAWPC+5lpw2NdwR1OCVviYyTzFiBVHh2JFoBl
hQ9T7COLOVAO0E4cliSXwR/eW4RfMmLXuUiqY1gSGyM6qvuVOb0pKHEQRLL9gbpgivVHuk8N9CMR
sWkeGIVrpCv7W+fWguugnTABquGTlAT5NcOcT5ShxD3tGu7YFNkIc+RxU8RuJLj+I5Z6kMjxdacE
SHN4t8HqzvahiTe5Yv8grWJ+PhKBHARG9j5pGVqLL4DJXX6b3k96NDxlNQ/vfmCU9XtLw3hwR0an
+0K9Rg6kvSy9O5EpwipSsj2jGG77sI7QxLg1hl+1LNFz/DDqCOjsvVbdXZWZEpFB9UFibS2qwhjK
xv89232yrVK1HpTwJXWcs7pNsRHMHJl7gOA7zI2LTcwvf5YG1UUaMc+4a6j4xMaOZgXevxaThcxO
face0rxjRBdvVswYYz6DJs4YRyB/tewDAgZ+nf3731EnX+K+3Cet8hYvQrefWQO7UOWtxnTvw9iy
M9HpzpvXqgYHck1bcyjBlaQo/YBjeu20olWqavDUk7rL5Nj1F/6scvOpi+J45zm1/oLa0A0JuaFL
55bHZsV5qk9MWk5Ja/WJqMR9qo/E/Z1mu56RFDWqUy2pzcxlVhgGk9aCuuQDv/Tm3fqd3dvVe+KM
JGbROxOyewp32MudfCb3gdbW63eHBxpWdNyq0N9MDkOCyopsssaLkojmf3kYiWOhB1FTBJNJAMcH
v5gIcLpINK/Fs+ZzGPO0Dh9qNCC1bda0K+4qKD5245ll2xxirmf81Au2+uzrr47TtE0rxl/a+WJ7
r1Y/azxLkrXQMenLYSYK7tUEX3Ywi9KfEmlRaQTW491GVKa7IfSaWbO/6b4TavbDwnGi40HatYri
KBC+TAXjFT4e7eJymzeyLCrJKi2QrywAAGbByGF8PXMIJo6QhzIbXXYozy1JTQatJp7DtApANHPB
7Xa2TJyBkwUTiGXnZ6s79FknJXKp7oAgicXx5M5KyH6PFJ3KX+I7DXLcKjxuQGvCVxUoMd+BUwSi
QAUW3rns0nmfsSmBmdUhmXwSqJOT+7PDODkXmnM0RgjRnuVXBrGbUkWqofvPSHm6ZYKj4BhP2EHB
UktspTljFyqXB1jQl3QTQh5ApYpppfFp5SjqE5oIDlsIuUxpApHJInWZa13HLvIigQ1H/Ia98lU/
B0UuzVNJkp/5QS2ilII9aauT49NQH9QJCvDJHz0Zag+0sf1z6evo37H+0FV3XWMIzr6RDg5gG8rl
1alYoUmt5WcRcq2GrXcPgcniGCXn4zkr4G3/NLe7vOP5m+QGe9QWiPyGBz6HINEsjJ9OEZg0R3nu
yNVV3H6TH888d1d+36U6XJw9az4UzSXFPf+qWkOY9endhHSJNJiQA/GE+N51RzR4c+TkJGVjFnuT
vidTh5akNFGzja319fLO/UsEgpuK42lqTmrafBv6Lawo+t/org2oF4Y6JUar5B856/XkkF2AfN6t
Pn+e5lultufg7FmWT69QZl1k7YbASleUaq60SvknLUaoo2qzL1KKxsFrxi8PR7yFm6o/ml4uFuQs
S2nfCjOpHAZLugyCxuomLpbiVYpCS+wG3mf/NJfjRQpvZP+Ap8Uw4EvdVC4Gyd8P80AxVR4mF254
iaV8PJLbUZn4amj5Gxk+yOr24bcmDHPanepWySeZrtYKXgR09mw1MdyA785jiww2VDVwBa3G4nCh
aY9Y9sMRCWveJo5853/gZI70vkm+VMj1k9M36J1RAHC4tvdhcbBcaCrMWaPM6tRBb0TTW7ONvRuT
aPO+tq6DOVSh+T5dLs0Xx8gl9+KDOOdcPtJmWa3SAz7SlBoi4Sr2JD1dNJd41rdxqD8VP5RYRvhZ
7TjysVxVghPceQywp+8NqAKIqqWHkycI62gHxqzix4o+h68L6sHFdQbAZk6XNS3BXHr1KXSLJTXL
5UcdDkjWLilp8GKWTe7+2fEQw7x/aE5fpaJLBcAJY8C2Zpq9MkXrU4u0+Hbh/KFyKUCcyEa5IOtK
WPhTgJxfRWwcHPKWoFMiD75vXbq2lsAQpy/UafOEm9w+Fj//JxXmtFr2n6Tl8TJu0ZIoDfrEAh1h
zhhHR/lAf7+lBK98rJark0p/zm3AgJ5aiJzWmKVRGWNrdAvUMr1PfW0wLJBR1v8iQ9I7KoGeFmzG
1V0zhILVkbHV2SEGq7Y2/PnGPWeZoSXiWk6QGHuDr56/fkTr1vDWQVFukcQR7lzGSPH35C7e2DV+
UY85+3irX+umM/PwLgMEY3JPbv7LWSH6hVGCyx7oKHLcX47mSIGuzTv08Xil7lotL1apT6mnqtYV
oQoJt+wFLrBnS44TiGPqrMGzpk9kOKuTq3J6PRJH1e24IecItxEWnEeA4v/eYPtRWCaN5KXoWin7
fvwZ2FkIWlszpmIiiJI4LW4uZ+YlTUzLcVCJDKHtSmIR9UZzG2n2ZiCFeRpnAga+xKU2+akw5nkA
qGo2yvritB9oNlS1ZnnKrOVEz8kkj9WrQk52NEMyNDhYxJhVLZw7IsR1b2tt+u5ztSLbSYm5LHny
WNKbxkFuXltwfNdgkZf+ehd0xYWOTLtIF4txwSujsnvjrd43o/SEmdscUDGikcYRDrgbHSictF5P
eVcjr35GrebQt/lV1Gai9pd718hjVaSpsnJ+XsgJSXMvnf859j4Yb7KgmBEQFJ0G+RT6pBF4qEem
udsus01PBeZ4cJfLeTuni1HW8NxazQB0j4Fh5PlEtxmGTiGADAiNiEr85t1dnQcOWl7JRfUDHMlg
q7a1E5kJgNVEwaUEPUCjmlVXCa+95cZaJIm63li6NFO7WHqwAAhdwZYlvLWCD3QIBqXOGh+ZPbFP
GcOM/bkTYztiHon8EhW+qZN9yfWb63c6L40giGX1PRViPU4itb+REzWE94EDXqGpct2PVf0Igv1d
i6uP6zuhIrWU8brCVvJDSFeCtjGY2LdHrygjvomxTwdQma/yTOP+yvxThp16EfZDN6eT4ld+eP++
WBfHfycKoiVBr4Pfpzi8qxmVedPrxlC/KEisyQdug0g9lP2H7oCZtoPGjnsddHYQF3jP6heNfHb8
vXmwaGy7MK85B8aJxaXKuT9/d+b1HfmhmCfoBiNSp6tMZwZrUE72wvX6GZS9hJKm5kY2ueucfiDm
D+N5x4a2jcdgM+5yY6aXWqOjlqCrFc2B2J9w7s8DUgmHexOMjwDVuGuwwNmwirZqHQMYGT3zv/+M
1uEYUWZtvUcnemJ+MT9BqZHaUStFluMjEJD0uuxWijZzwmVw2uFUjtYVZ0zft1w1Uvs+qM9l8Bbp
bu3Na5MIugj3MR3+2TAbqChj2avL1cKA9tql2dF7xknNfQjdMcOYVTVSu0ID6ODo8maHy3KhJ8wL
lrXpgZuHRgttyaZHGOwzGXZmnO5ER9Jp/ELFxfh07kYp9J6cRrbXV86JeTsAsGhADLc8m1/N52U7
YvgGHDBa8JiYn2SaK3t8J2fhBLnRLurDD2rsVTFOcGcx7Rcz1HQlLmL4GejyQrTulw85uzzGEbeF
m+6CE6rcbjrtuKVYRSpTA6LlnNbQtQ+0dUoAzGzdilMV1skc6B3LxgROvCSXLqje8snyRZFDvtcW
6TcvVylDHXl+urFDF+blb0mnW2coywVQVoa4yv85rmxPZT96Q7EpKGySKj0V1rUAhLwKgkHGzkPI
o4EMq7vdyusMdL2rHb7M/abZgo9ypKAUrsHHcODEivIBWFvhGGTkva/MlxMlzu/+lfocWLc7Izr9
f8IstoONrMy9De3kmbU5luDSPFghOL0G2EpKDhI3qQjwm8FpJDYlvdnMquovJFLllg5i7fET5424
qN56bnDGeV3svPCsqZz8F21Rm9Pg2ExEYw/B++5uO+ZhHZgoIQvbBFYF3sbwsVDDePqyzoTqMY9X
WNfCq6kufDf1OMWC5BJO8wCD0Cj1Zo543CIttQ0E8SqSKk/Kqw8iw7Z8ECodOD/zeRXSJ64mfE9S
QUS1kT/SVTe1PR3UuySkc1amTEAQKJjrnQ6UMLkjwEyqUx/i523e7ZuA+T6yo1ZxDjtcwN9UN7ph
BQpASgytLLeUmPcD+cUdniyrJRb6tYwK4vi62a25gYROhULqvnNJPXN2C9p8tv5NpDN610IeaHgD
ZXFgcaYPEbND0XAWXRg3Eap2LYYVqHEafd3mwxdCtzqAjerPKHNN9A6i7u3YdxUCsFmhJqcdGPrk
tFePpypDqJ+npWix/NmUdDB4qTUQ/ozVY5Q7H5rTc6ZXXvzQevU/SKb2EkYJj1cpcFFT1gAurSiV
S2sPCKL118GmP219sF+uuZnI3QmCBVEj0Bcqm57wBa0/KH07U+f69NLbVzB/ilkhwg0YugCZI26r
frDZO6ylj8Q6ErFZhV2yzH4CC0+r1Ib5019BN86Xo9Ud7mCbw91minLfCsUdGbyofx0Un2coiy/8
hjpY2QYNGLZLPGyEPBtisr8ku5p6jBuubxEDEtm62Wkgbp2vIw41Z8HeBo4sCjUQNDYXtaFxMdSO
POm5nn7lXROm82jPdvg9p/bDVL7WptmWCi3x7Tn21mCaFl+f4soOYMYOFHcN3XCZGCysSwPT3B0c
27CvCQ2cRqgehfjhIbaSEA+EJWcamp/AXMCU1/ksZyT9w1+zetXsbS+3qqpl2WVBDbqgQI5YAeG0
ugx01nEfUVZ6WccQJJGsxXbrWR4UqyXjuFkDOeqZYTPYKrbTb8Nnw2Gx9leMnWJn6HDgcUi2Tgue
OBoMlJ7L5hj2S52od4WmPF3Ps5gq+0AtEcBxC6T/l5o8hGHseD7ajKd9+t/IUI0RbOs9zm9ONaNx
TIh03ObI0rsdaGDY5UN757LRGM2DyPfyFbep2kxg4Bn584PfxylUaQ7QS94X5kbbL/cgU9kpPNo/
od/u+UfERI9CamD+kZ1HiNDwLJ8X9pXIjX9nin5Lrv6lCMebOyo7ZEATMYi3cWYVbN25HxfC1mL7
cki02IYT+ztGLwkqbmfv+x3/TY/aBApmdNAX74OFvrRyU3GpWComB9SYHDis5bwDJ27Xpa7/AUX+
+MUeGC5ijtUE8sAuMMLua216lwvWAtJy5wXzE+3ndx9x2MSHj6dJmpYPgwyCuyZ50IzwunDG59TX
LZwgon2fNFfuHL14/9/6JRThJh03b7ZklZJK7fUP2ALtN0Tk0FBRuIf6owotIZ7Wv3dqjZZCw1fw
usa5QrqMSNwTld22v54uQ5Dpm4SiQePn6KnUtRX1iW78ym28HMBZM+Gpk3QCbbZa7UWC1n/c83mb
vvuzxHPz96+i7DdkQBB+ZTGw0fToaw8V9U8KW/FUSLsEs+nwBWPyMvrAwiOH4izRX3xW469mFx9n
CZsgkb+RGoPl/+Hv7kxqqlWYIZDc82V0uHVqzlUJ/Pu2hAbwIOSK1P1BuK68ic0FSNJLQRnsLSKq
O2iYxRWZXnjJoRGHYMZDnJnw4/5ucOft6SYG2rdd3bYwxDifdNXhiBNdP2x4Yv+roIgI3YyvBsFn
gCFyS3WooJzrXfK/B1Dv60F373Sf97pKdvBlsURYfC5gaJWxI1mZJnmIIHeIdYXgRPtdgUuZSrbt
hGUmul8tvdF2pM0O13Z2hm8zmwKPypm/skWW6mxhQpuWJ2q7BsY9elwRHOgKOhNK+7r5z4jra6hF
ekNDMtoQe37zMd+khAHY99PL/QJdnsHZ+U9UJf+ZIGM6q2L5VkIi3J0VRe+9TQHnVrGWI9tyPd6M
Qk+AWu2tP5VUOUPud3jrqFBSsthx/1npi6YjBnMt5Tjwp5CZReFsHqgc8MMYiQGOe7ZMPmuABuH0
82O+zMARj2AzXPq1k0PAg9TKVq9P/1S32NjwUNVJmY5EzgnmWHwFa7OXVqseTS2MO79EyHizWDN2
S88Ff5+lHOk/mSJTsFPIIRhaTvuM5/C1aiyqeNxMDMGo9rs/I+1CFNGRCjQyE9dGRkXD6Khrx/NC
cqtFLsMY5WtcCfmwnJCRpz4NGbmzN8C8KLQ+Stln/ikmEg6mu4dfCvl+230pW0urpc+dN7hG6zdm
WGLyGSFNUtZ1fu6sx8URf7TG7m6n6nc5/hoaFtmW0zbQOUnxJAuehw2s35YiknHGvPuQRkzhIKcB
hjBNTTra4p/XrjgutAOM0/2OBlgCJXCdM/r/mG0WxrJX23rOwJlmRrb20V4kqwAeHkGEfl56fFJ/
xkiFhygu8EdTuGN3D4cJAEPQwlzyHzxteFVViu8iIzdi4R6gUxi6kMYyTZ1gygft8zcqbdncfQJv
QI0zziJHWzHVitMIVE7tPQtAgvGLcKSAP0lL7VDTueMh/qPaRlYIDqUmSjln7f1vbW3NDdQFi7tp
mIOXtZ56YrFayFsj59wGqpbnum+aDD9iiZgFB3Iz6eTnOn6nqdoN38jUg/wCctULkV0110OqyOfX
yrvsUhOezXfMywEPSgMMYFWFsvUX2p5GzZIHuB4BfutljSBExPGsl1CRqIgd/r5VS2ZCyxY9wwpp
cbZDFt7iQOIIBRzWaRO8qCg40JaYcKmc3W8N9YVvltuhGqC0mnNNgzgISM9Ml6ij+Jz/l2yTQ7O2
LrIxMSYrOxNkIUO1/7z+aXYzc0d0RK3EnWbsU2F6clL0VWITp7GoJqmxy6KmC+4Ss5QLOdOAOBXD
8x7MoUfma9NO4bj+soNYmvhWQushfyvUIqUFx9KvtfvTyRsasL+cgCGfgelXDL+lJOpa8LKSUisN
X+Ml4tN2kh8gZPQIrmjbMmYMF2Xcp5pGIvebnGgBnYFT6IH1brNDAvt/WvqUmrhp9Avw3Ip9HvQF
dvUB8i4RTvBlGh8mG5gyVfjCNEDmBwJ5G/X/tjigZCL2xb4TJ5f9xJp8Pwgo8RzlHMdxaCxm4hkF
1vvQ/4XnG+QkFjzpNcWzLD08GCVvV85DVGryTs69oNP/4Wk2zCvZAf+dpdxp0tT//bM/5ATxUzuh
IBDZtkXUZHB3wpjy/cC22xoP6jTtyv5ealD2vFcp+YuMNPzVHqQu7LAio9ZO7t+5eefHuIy5YEcc
mbC9NStFxJx/DIQeRrBxU/Qza4KTsqjHsEiZ3o+se2aCp20h+3puf6kGhABkF4/UG32cxcF2GOpa
HZhiRWr4+VAeg8xYx8ZOkLoAfwqYB1LvZ2vMJkdZnRgjG/ubWAFZbkKBwqGjo/p6Y4RF0Kxq+iYj
vbNqUJVRt2h2jfLGlalRQfeZh4qampxCxrxuMnb/RQG7PMGbcdSdSv/bfK+ZtkitxTEgkmPTU1L+
rhIYwYiwxA7J51TKN2oJRqFCT7TDKNVKsevntZ+oVkyKIR1+d4ZabilE4d41Zdjztb4A8ZNxzvVh
yUetRUTewwidwUyOhPs2NXBqJXJyF9Pl5fQCtrxbJlR+a/Nn3UeYfiE+kRnHdKmEJtHSQXq3Zh2M
oP+bFKGC/6STdsYirqwNMHBpfu/kLKu/NWLDAWM3ejdG5ZixkvIJEOlcml7y7FF2p4F63DqCNT9x
+5ySmSrHebC/BtwX6ljWNdpc/OR+SSx2ZletWL+qB2rxpowOtHrMjyJStLarl2k/pINh2kBpgv6t
nl1tGj+G7+ws7K+s+atS12ERpIsjmEFV0n7NFBivr8tInOpg1wlyI5mr3eobodJHtgRX6sIpibCw
2DoRtd94IQRVQrc6+19JzppfNNn9YqZEP92mDMh9fDfEPt2I0M+q95ERo24LEe2r6yqIFZWi2pKF
1qQiNd946f0cvJXQnqZTKaJeWnLFDUlMGqH88OxZuDdpMLd7UiewjLUepyedUr17pjXK5Pl9vUc1
+0Y2usfLm38yNGEiWo07cA0xHIulGTjWpS6gszPF6wfaVJyBvSO+WBIiktcQ1QxOhSbjpO7jK/B5
1s0F0P7qtWv9PV9/BhdQTl714GIclRaz3KfPJ7ioYXXVaqthqnu92nkTyQiVDjeKMVBbo3jlJiQM
f+4SrrRTl9Lzgze0VhIfY1HwfatUXnL6z5Z4cHHwWU1GQmN6Wo/MNB3+4KWIOLtiAoOYNsgoR+YC
/rKbiMG2LRN9fMdtu6Wk5e/o2jWbs/9zkTdY4y1pIoWJB1/d0zyhubgXVfoUUGLWhCX3yXj6fvN4
8wELNJdaPlQHCnKsIyi5M9AC81tLZZvkbDue0jXhX9AG63d/ZVkA+8mY3D0r46Gw6jAWJ5PvuTXE
9gmovvLppoTC+d04VdX13tQB/OvfJSIjK/URz9gKpWnsZtC/77rIc5ZTrpFjobppAKM6F98dFGZl
lVU4wIiQ5pLqysbMhBvU10FG5/8RlOOoWKAsHSpYZ3vWeYlDCHF8cYGGntlrISx3NKSsnL9fdDhu
r+xgJ7e3CjuB11y4YLPOP2dkNNhU4pji2pYeWwDjsqu/X5fKIztgQGT5dmyo668K28TDUHJ8sYai
wzCoZeIXOg3wX8hHAwN7B29XRtEWigm5AZDunI/Fe4TRmzBeoJ7oGo/1twPsnfuCjut+wA8r7rFM
sY/RBbTrvrO9Tp3mJ+Y2TitAJli3v4auxJN6I+D2TJdTz++rt9k68XlU5mLF7Yl8r9d98wV3u9ic
5g6Shftl91EoUpKXMlNsJmi1U7Um/zLdihLJHJwg4o9f0lBl8bXT09TA+1Q0PAXjKepOWaXe+zWp
3M8AgQCaxvdy7r1+YLXkiXDFXlhLXKhYWFeeLOIXSz6WrBiWZVm+/bvq//r8zxvwLBio1xsiPL7k
O4T6zw9ezG8i9Nbj6GflYNb4y3XO56g7JsPDdAkZi2EjDSJaELBV+nte8V8QBbVPl9folUy8f+qx
7xAC9sm3W6MKBokdipGv8sLB8PIfgNcE1mCfQnnNOujcRaPMGBj+ZQmRQf7RIxF2xQHcXly7ytqb
Blxbno0waGVIoVHWmIHigCkLIUJAw41smTG3VKYMDoKWZdcWwll1axUqiYRboZsigHgHuiCws0O3
Bw16gFI3bDN2AfJzzhkWK50edI7m1aorEjLk080kZ4UVWbpujL4A6TCFSyGJycRIoVY4C7wL3TQZ
zrjR21vhdz+oZeJUxT9rUS9l9web7Sd4ci4mTFYGeDDsa0EwZyQgkTJqlj5x6LACwfLZYk/CDztZ
kH7x8fmMe3fVyeRWL1APeozaFoSs3ipmSbi+MTJzy9w2JaZwa9sZy5ECkatkoCmZDgzeYR0SQ7mV
V5w/GBAunKOnTKtPMdXB8rdHj8BTcYypHABOWixpO257QiYjqZybAZvPVGM5ALSXnP79jx3SrMtw
adEn5JScrFiQLN7wcyuj66k0VoM7T1GfOoiGFj74MLDba8TyH9RC67gMUcoN0GiDmvRqpqe751S9
AeVJ7SXdROPy0ce8Cjmd8zlJjvljuWKvxIqbJ4bT1pyCrXkL4mjfRaRpfeYJrlEeIosb3f9UQwHs
XfFRM6JC2cO962lO0RRM+4cfuwY/UD4hbNSXyI22dhEqIg/Qml/BSz0Ai2yxgB2qFOASEPUidng0
aE1uxOVkaUtbS02zknk3otWQqT1LwR69L8PZxF161AhdKXykk94E64ZDBE3O+tnQwmphEclBkJx0
fuCQWlidaqhp5lLguGnFb2mV2I8qcvtv+HBgY6arza3OZdElS3FSQvJuKaXleozh7qVNlTTTEU54
PAngZi1tNgSjllrXO/ip3PhJ2ecabsthnZlPQvzNIC/IWP/kpi+IeD3y35Todz4xaFY6ufp60Vp6
G2jv95lCQdfZOh0kiuVh0642EvHjvVCcpzlJuPYs8W+5F+GUn375Lki3W8ZCo6ph6uqhRxxECQnC
Be3FHg6ufMSHCO6q9Wt27tg9UXqv5L4ooMQQveIBxMpjTH/zVL0NZH7c91LwtjAvKLifsZ8z3ikS
onCumM67NrcHMqs1/nGmKaMmukCm8ywbT8eFPg73JUnC14cK38/IbDvlJKshX5gnAHrXd1KBvTpH
LjDsJke3NH2qqQBHImCLlCjQ0cdRD29012dmv1VZtDHllW9Velvx04rMNcmSFyxyK56X6hVfM3b5
mm3DuzONyqYpfMQWW2Jtufq2Z1BLYm6SLBlPX7R8/fPg0PJH9Hg5ufnGNipDm42XILEe/8PAeLxD
Z/F/TvgZFdaKuYWhbOowp1OLKgRDpsiEnolCelWr5hELjNKgTDzN0tWy580/JnLQkPZ5LheITGQU
NWQRVJfkTFPXoo+J5GZXii/MqUNMmW+q1atzZmG0MLub1nHqtLqY6I5XhpuRcD+yc6V28JUuRAzB
QU6tZnc5cgl38hE0UFhi7sYqs1f38T53HaKuz3E30welt42PStkvCa7yJHr9vCVGO3gzuac1Q3c0
EL/oXAIdC1zrfYqsXGHzuKkAfmNUXQOkGLZ4RkB2SqrjRUF+SXiSMvjK8p2akE6akDmXdeHmW6rG
BvP+xu9XsdU9D48wBsuvYUyXRnFpi1EhIF1MzBOymW/gvgTLaJ7eKJwCIUXC9324R5hM9kfavSGr
82Y1eWNBUQ359KTQNcroEW4RKmqxi8DgGvY6ZX2vfBMPkpLisNLlDJ2ZcaxJ6ZG9GlSxiWp1r7/0
dC+FrRO+dQvu0goPnh9H6ZCMqnWsI8X1LIIr0b4RfZF9XS/XXihADSQ5sMA+HDavmlbCYV8NxYQA
tXW5um5oA4GFxySYC/N8UiL/cOlwCM3EapnpJ7U4IVBnrgs2pUIrLuOPXfv34hzUxCziVYNxVr7B
lhDjlI02Ax+qA73LCXN78CRr+DNsvSoSyvNNN//01TO1vcXHLar0dsmQbPXp8y4KAphiWnzEsJDo
Ee6o9Pijj5jePxE6WngRbVno9zu1ff8EIp2yj9VAe9M06xdgRGxzNJVf+PCJ1qYWewgX2Zfq2gsB
Xcp8OpDvLEES4WDLeAvtoApql6MTSTIOFJJpgDMONYNZSloXnSrA05a/z+olmxYD63yyQobWX3ct
OMmA9RnzoduDsDr49zUG/O+c+AuL/rbfUdp5nehKM/pLPmJAPcjfqpI7MY5dWHlZU/55/vRm1FdB
5yPD5rDFisZ1axz5IlZPg3HH0T3+8l067C5BBQ/JIPfa6wBVTTou5gCV8K32/J8iVxFia9T+oiu4
Zbx+EdUlZs917yLl3hovlyFFTc4Dz7r0wyV+riB9efK5zAwziQQfRLF7fFzEFIcGPd2EoA7Cse+X
mxOE7aUeVpYuVtw6HAJ0m1CWhD/evd+FQIRwReE6GwGs8NdAvZuUADXDvcVfyo8VmaeEh/q5/Iq8
yDY5DcLleHMV4sUpWnXuFVdqrbShVQD1wQV8jElCzFAkNGJlX8nkw24iWa+Fv7VMddH4JJcgzLtu
PBl2hQNdGQLeoIBhF/ePPh4DWZ+ui+/5Zki08RRKX5AEyEwfG4PeQx066ZEKB9/DsHPdAFnudQBu
34iCZN8ilsLdhPYUdpqzJKP9LmVZdOxSIQ5BUzkXm2n1Q6O885UruN1ZiIRhbyzxKvvr90EM+129
UxevI07ttnokdPOXEvw6ZGDouM1rjtjd5nQbMJLmzKqZm5x2miTSg/BhpSEyPV8V8C0rQbY4TS5G
oOixIeIvoleVdW1xq6bnmGWGL6cBGAyWad/XEKi/+hmG03+Lw11GxUQIhyf+ToBkkgXbxMNovYrP
JCna8ebQ6CKGI66khkmHEzPO4O/22GVWTFS+T1jzamvPFdpudpNoR9SwB0VUWXMNZxFJt0es1T+b
YazFOdIsW3NlgyY+jhUgmesh049mlJKu6ojsfHufQbBD9YpAW4SBuvOdyCu8b/rAwZ/kXN8//1Fo
1RqZUbi6W1XaUhoSFrXD4D5IgldA7KGK3OKK2aMfLTNhdV/vbBIkPf9SRfnxWHn6YGqkmP5jRORS
j1RYJvnWFrCrc+OB6BSO9U9x69jNkEMDPFjuqqYYlo4nRwRPaym4w2qRyXDvdHFZD83+LMVQOPIW
32Xi23emvvv8aC59eAgGnZ/bIz5EsCo+UdER5H1wzFisHmUk6mmGoqAgWd5fl2pEytvqCW+OwDaX
k9g2K1MtVJ963ZKHR+t8eRmVwlFlyckknwzPzxJMVV11qjjC2Wm96xW+98TAlVQrE76D6TrXlfYq
TL+ZzOjWqQxj9g/1yFNWrIkMMHnWb5REx8Gqzk66F7x+WpBnB5ho8nMfEStJT7izjBx6M1UKfOyl
ssd0obAk3DJ0rZcov4e5ApPbB5+vfmSCKIInaq3qq+ntS5wCkmNhI/GYm6jotorZqexGaVbBOQvH
4e2R0/5e5MQrcG5pAsxaRLBv7p9etil8wblN5zTjnUs+4PpZoQHjDaL9u/iR047xH8AVCTSnl7SU
RVFXKfj+N+VEFNAfRzu4go7WTIX1qZztnLWpqzAS/CZ5jAiaEOBPWku1DuNiTEGQDejRiI2uGY2k
fUVm9FsSOD/agDVrnTXllFFyYkTypeOiFsqmrIMeU3olZds01fY+EN95DBAFNZS3DLgJHcUFqcy6
87QIsjSlAGxWrtprjgi7FBQARRXyfXPnHDRKvGLPzLPyrAUDx0am7YR8tjaznMPN3Zazuayon1qD
NhXrjWMZ6gg9Kw+AhNV4yB0dVDbB1/qLpQ5wPl5FWDybTXwTn0l52E0Ger1ArWL3PXaaHJ7aNLuo
Feg2B6Bj2kQCi1ZED1o1fVeNxqt64p2s+BCsgxfLcxnzM6AIVOvYJviK2u9sBSuXWQzq5SejqhOF
c7JE06riIu3IOcyKp4SgQbewuKsMk3PRyvvF6DDC4W5JCNfue97SES2/gA3hXZXd7e+L6tntAlAe
uku6ELlHdK96AxILciMh4Hz87MYm+wd7gTh8bjNDxHmt/BM4pgxdimIVJn4i2PVurTg/XB2P+3YN
6/5NQmD527zuVD5g9K0rgDrpKwHimD4LBN4uMRfZpszoePuQ3JEW8KTdZzOUNrjyiS+2Cw7uR7dX
pAbF3yApOYprhh++GmFxr8ox1zObmxVMfIvQ0/S75teKDkiMsCbXsqMdzY88d05cDGIOX/JoDRnc
RcXleu5E28TsOxn4OknrXgebZcc0ia4E993bGQ6vWmFn2VdPYi8rteWHxy3Y/R4HpCGdFEI8TNHk
oi1Ez7AmsPYHD8s2KtZq+rkFbKt/SsKj63bMtGSV+X1r3oEYUMnPB8CbD4Luqc67paJbS9MkCPu7
A1wg86VUUZaDm6kUyWby0aYuYo34aoenVPlMA6WBbhJt5oPzVLHGNr5nQneyWHwM4k7txZHBhtW2
ih7niOJsF1JP1rnP74MwwiQ9wOGXK1NGeg60oSIrflJutlfp65R4P0WMuUu/eK7p3GEDMQoCl8qC
KYWgv4DSwNJWsV16eVX/qsPLAYzyutKBieDv2s/Trr64j56Vazj7fE9y6Mo99/xTBE+QeG4RyaKa
kAPmFFkuELtNFmh/6vhRSFibrNzp0Bqey5PCgp3eLSnujWM7GWZLOrpXJejEdrGR0nmJPQlqJICn
71wrp8k0+dtiRlDQ3eD6XzyEOEaqG5MQBWBfVWCfZFg3wuTJzcgTXR9Xq18L3M88OgVp+Ip7+v5F
JaGvALR9DTxu5PCwYTbGQDhLTGhlgnO4Aukn669/O+ZKjHqWPcexXYgVB2HEVZvfiPKnJtHgFbCp
huyK+n9IX+T0gGuxmuaHt8GW4C/sDeoyTL3sMShj4GkPQHdor2j5KjovBYWCwZcCjln5mVNJHnxT
6XvPvXNI2pCWpNn/pB6w7oekuMqKKKTZInRhpiAaI1bgykAU4ktlkd69pntBQM87OiYC055J8LXP
qYSnWITyTfwQPB0VpgmOvQqjNE+Ifwa0pqBg3K8uiQBeytIz/goxt5Nrj5KMMxCZxmJ3aKKKVNNu
o/5go1s9Aw20hNILVgppa4bse8dvSAxu3Ey037oh+bNVcHnCWagfPnBVcDiM/0TlY20NVZ2pwCf+
RmnfF6kVLUJI+9iFgD3LCRJSF9wzGdooEA6MC8WSypXfruiSeoJ1w5GcJiNrqQu1mLFZ7k9a2VE+
vwyJ8UzZHvw4N95JeCWX73RX4G5moLMyrKHLF1VilDNXwTi8y6MHIxeDUp2NfC7SU6uxCK2d4R7O
saYPmR2HQJqifbSlksbHWol39FlOz0DLc/7OHRvnn1pEgQ53NAJnGnDgC0djsFu5SaSFBuacQgn0
V7co/GbiQZ5g1/TrdzysiGKZwWJ+mYDzUMO+fotSC7dkvX7iU6O55nbuj8RnxSYzWWRfMzelb2XJ
UCMAbwutf7GgxeupHmZwD5bVS7d45Fu8GEZIB793Ly47RRruiRieUjd5w51FHvtitXfG5vrPpKlB
/gA0li1cTFDmfakVrlLx0/1K4+ZuMGa5pZ/RCBzlh1v8YGIzbq3jMlro/dC5/GOS0pj+KtdBesgX
lnHuksjP6GbCM4AkK+mxsjJAa/e0Wyh/L5/VDYEUfrnTD2wvknaj3fM1PqMrc3GidUVU33rgyQdX
jJQc0rU+raS87trR23sSnJGYBN8bXahWSeWmm4VICZSnLzOFuZSojEVe71Z9vNe36K92tSC/29tb
pPL+h1JM350Rglt5DmcluCymNM2fcJseMXMsCcx9bEy2Qd3ZU/HVVPNNMvl3PXrVqrf3rNjvySEX
fPKOGQ/ytNRw816CSqRzs6I0My4YNhCPhxBtEQdyAos+Ht+lLsIMS5nsKGCQpxpSDMpA1hbWng7V
+22CB+rhHhpagA+7qW19cWL0N8zLv9h9svxGWAYU6BLLLt/GljvNaYPmte6d023qFT1viImkArzq
SEAH6njgD0U8y3Wj0+T1ezmpt8T4b5GAXeue03Hc4AfP7NnIFo/VDxLhVErLPYD1DT4TLvszpm9Q
+TY1i6+wgJIa4Jy7OUPXUBeMB8BDqCQmYg7QIQj6WaYjqGU1RTx+QLtkaVzCMVgEIMnu72wL88DA
CPwU/l/cg379hZwT9R6l0Myd1ShNgCN0zbjLAjgC5OVbz3F5st79HmDzp2nxg2lLHixZvEUERyY0
0djSoRIQhcJMXCEZLZhStoKNxUSEXCsmG3ZJ4rJdgqCARCmwMLNmxZGXlWPQrOob9VJ1Wy9SDJI2
ZE2e9hdNSvhfFjvUv1s73hcbpeJdEgR+PpQg/KwUugSJDwoAdHizbHaySgm0ctiQMp0ugCkFFX11
BeO/d4H/1YU9+dLHRWxQ7kc4+oaW66gyoIAd6P8t3CwXfHqDrZzOGDVRkBeSCod36Ktmd/H65DfU
INNbxrQXWfSNHyzFuqgsvxlwjdcaqwsR16ywdEnjmgv+gM5/QkhTiSb7qjDAOXVXtGB0eh4FINlo
enF7aQkYDb63B0j6bCvJb42VRbUTa5UOIpMD3Q/67gO7ZsTq7lNUxGiV8DoIGs5fxIrtGBKgxPDZ
CKSrw3dk0GaP7XrDZ8juFdtJYi95xJGzOVtMDTbAV+cJ0RtTG4sCHpbw/wYTtZr69kNV23ftC5al
JRTzjZe07HvDTVvqVsfww4ByzS9CklsZHppmrh+6wDn9kGhQ0a7sMVWOZkvP5b5xb52rqcXO4Twe
p2hmZDsH/gL1Jcq6SbybTKgdxNUJZ/BKF1rjex6PGN/SauXjXhSe504GXyXNi0ECZa27N0uddGEt
n3I0nB+TFkC9D3ON6kWzeQ2Nw/6sbnnO3HrMzT72kbzN46dM1kJ9yqnCrDWPi+5aLn3CvaTKhxuO
E23G/gkSxC374XKVj1Q0vU2c/9PJ1OnDg2c6lWZKOCOIyTmPYVVFUmq4LY4ENNy/1SHctdiHF6yt
Da7OM4ug0tE07/AxJRndr2VYW0CDpP1gh5+LgBJXB3xTE/kj27xC8t302dXzulMilKL5DsecYly5
c4I5pbbAUiwMua2QVVK2LIIJoOT0mh6DKpT9ifM4bEVB+rOl1mhExCNxUM/W91L7OWB0xidcWlFd
tU+Jv6Bu0iiFL9tqVAOUVwQpfWOEExcJ3tvcZcEh1lprt4PTw1Yij1uQ0LFMCmSLnv9fnoYrVPH3
jlxH4Ja/pTzSRkx486xDAY+5PqVQsGPe4JFzJAO//ho7k9PlpyQsoIsCreyYHeOjW57JVwii0hRo
0mzC23Q64s3HR0SnymtL8CKVV003Wan447H50wZ9Q/63O7ozHUMVhDpBAHzjLeeoAFTEgxalCZsc
PojTyRGhhySnl5ZUKNQkNaDLih2Ttbiq3vFJ78ZWS8oLDhLZSVBK23yImMkMXWt7jhhe3OMn3P+Q
5p4RKuCiZp2KJSORmMQbX63mDDbGAwmDDlVxHE2P20yI8Xc2f/aYGl+AClWPzd2Dszb7YNjSsT3N
TMCo5gZ3wMjuecrNL4Z3tdb1uTlzyGp+yDIzKwlMtyAFG+04P9C9SvUf/xATROKgZbz/wJUEE2d6
Sy+3MKTQF+RqAlUE4E2LAdzjTtuFgOGB5e+9Nd5gSFJxTJ2GwubZtxRKYYUJDI3ED3eN0ZrobVBr
6sKaV0TOZCfH3OUkEZmMdXqxbIGXnunCAuBqLKk/UY1Zx4DOoUBXeUHzUFX52zfzzGwUnCD/zmHw
i/XPEbMQiDhB/qJdn04HutcJu0LW12bfeZVTKhSWpBab3SNVDXxYHJ9sBuCzC1SMG9AfPmly6lpL
MzdJrfbS2KB+ikX81yNqLj1wykqqSc6m4SsGY64dXO/Ik0xrHf7DaajNvozzP33ivUJSm5iCMp9f
AaiR+MRMN7//QhxvQbANLs8PYuIXvIVQ3L/YCQU0aOx0xDidthakD3WcHnYwJvSanKENhb9/J2wN
89GybCSkppa5sDoAc0uJfuZdZLIFkU8UWOsevWF7vhsWl1CTv4Gcin7wjqDcZ+CJJMCnlg5D04Ng
iNjPhNLZ93dTZSyHTp8qo0T4O/rb2lmIwhVVzx/+nNe+BO0bW4A/bvtHQ/vX3zMwGUvSF79oVlY/
IIXjybCiBRwRlqWbn5XJi0IgBf47rhcfWRpSfxTbsU+8PSmkB7d47DEH5NR8n5qJko5EO/wkDHtb
qMdTVqz9P8p1lVLKE6cRJmKuaKNm2ZR3A/If9WPZakNTd9KYqJKEsaValqGFZUC4H9kZ0HXSWajm
khRoWed2hjrUzqWzfhMb3yBN3d7xLo4JfvCGhCFlbxG3Z0pRu0xtbr9+pb721BJGeJ7xPPdq+N4A
lEVA1oyjfEzEXjj6juZKSLfvaWb9OzOPw/txcHttW1KRxm231cudbr38uWxHfyaHaQtlKNuDGac9
w7Vc6w3ZR6peN5KWLZGia2TKEeSJqcdBHrn7PQy77rMz91AVazwg53gMDmPyi+tVJtmQl7f3hDgx
x1XXvlkhbtCfCJeVuP3VfMhmnh+evofDXWEJtI8wvtng8ctCa5DbhbpBB3cT0QoOg9ZniKe6g+8m
q5u6IMTferbQUIe+NYHhXZBbqoInJA0NxrsWV0uTOl0yvBAHL3yA2GC7Q7lom2EGS0vIY2uDB0LJ
nyeF8s5dA8Ggs4/JY5r5CDNzFt0zLk/CufxtjLWugDYqhB8wK+/L2lpL9VCukOnHxHDJsvpqpJfT
JvhkmyOl8JyYNcQZpPCopAHZMmlKs3J9iMls3AqFjD0Zv6JkWkrGadWbIrxhKfMF78xBywwrW10A
lz5SNoZijoVQXKWbMoqTjHowyxYE36z934VPP2hlKTvty45dK1rU4koBDeQlNmdF1exKaP1+nHuj
FYp18QE4jf/N4gxlz++cCIaMKOEu6VLY4jKTJoSwdHXF4yIm5nunS9KejyrGqshdZkrbhhO2JD3z
pKkx/NkEZbiOoue+Mtg+ICCTgEKLepc5ZwII1DiaaRVPtJzmR0p7XuYtcSl6yz1z5h4lS13ibWCB
sZoO0/9NnpflfUvvz0fgEkJgTSX5fAlnrd8Y2yp2Hvrx71TXs+f+lhYVGxmnntMR52mxeRDcf7Yt
iniNd/b+iZkzTNdcWhRsyU/y378obqfEe3qyTAhjgG31ECXEhvOGeWlT2uNRefYqGCCtdQh5vPX5
DO2bkO19+vXybRlzCTLY+VxEqSj4QUsEp9MBmSo6v4OV6FD0+gZZbxjBp1cu+82ZqnmK1smPk6eC
OEQMnwhN9FnYqGBwLE0Pp70q6R+vhwKzEOG21+RL9sdLxL5HYeiCQn5LLc9f6OT22MeAgUNlMv+g
cfuao1t+2PtA8mDX+hpfPx6AQEUPbyJOAfaBUNrA3mbzCpgtywtlas73cFGW1LIOzeGaW5QwZ2v2
nPL0R783tprePh8fcx1fcJMlNADcOtBNVT+hTWjpm+XtIyQLnfZyc0QVUsIiVoe/bQ7PLJ9tZKzK
eewfyTuOEu7OwIAgquUPLJQwSfiK/PWxXjyK0gAVAB2P38VBPUMFEPIJmhilNKpcU+W6rVZS38dA
xvy7I/ScIyeN36P9hSp7Ulf7EuRuhR3rNe+SLgXxf/Wwb9Y4aZIP19Fv7UAb8RlS9TYINGsIlMLL
CtU6dWJjqnhs6kdRXO1X8Pd8/YG3UVkUeaOs3Fc1KV8woDaXs45CTvfODKerEjBd4fxJ1T8AkvsU
KUPfKlAel7pbk+JjvZ060YjrfYGIAmYO9jK2UQOrpxhBLUve5522zKQd5NpFRSvXFqtakZfv8r4R
c+WqoG5Fgx6h/gCgqCSUVlW6a0ie/XGc/gM2WQFG2c2quxIm86PZS7ad3Og5DQJ+0SSQTaAtUMw6
DeYX/K9xsCqiQGmVSibpVRbhU5Fk3RZEYusrfyCZs0NwwquBdCh8AOEbk+/5jk3paMwzh2ZiiLLU
UhLn47PCBOMLQWMpvxBL78uc3rEaDXp7l9sJqt4diwIF4BgDkgXibn+fDJkMTP6jO20D8B7UiMP3
YtabfOgktXUb5kyUXSP6oiqK0IDZPdU3IhU+Kp01yyb9uUOTxCXj5G9O2g6x/jszzGbXe+61fHqe
AfkvV0Y1cBNRNZ+QNytVtzBw5l5+OGPy13dPe0hEfR5BDzbTLtS6BfjUFwvMime/IGn0KU/TxOqx
eSdYMNtJqr8W5JY+xMZ55T2Xnl86BnepSGXD3/IRbh6jmZWQWJ8oOW/DmvX+Vr/ZQU6bR8/L6bZB
HEUN0/fS3MqaWf+UBFDDV4v/+DCpgjYbukKj4UYPvDHwCp6MY8buNE9+fV6PLKmiFhuUJt4nfC7n
BGrTvb57a5czorLHeUsRfybZit1S1wb6kdTZxaBJ8kSqQjoA/Qb7orzbH83K0OqR8aIe5M9crbos
gfV8lqJh8imDjuU7Nk78bnfHfgXe1teK8jzItSMgxXzCgE7dl7kP1XNJaugGRfU1pclPq3LudHQH
ABSlWBQ0j7SqNxeWIY2LPKUNhGzaoINAVAEffbUWKM4dp9bE26Y1BAQ8i3XPWFP5PCKGgbHzUFd2
374rBxTz6xA3mRxWNWcvWD56lDYo7NG4ojzuLjV+Q7ABWWaNN0X7CnAxkt8OmhsDmm4cGzw4l7IL
i57vZRjw1hvtSMcibyIFJYdMBbBZFKtUTiLhFudChaTIhOl2HlAxv3pRIcKeJ64tNb48XaAJTSVL
GQTjT8Z9vm5jlAubclVf/ZEVW7FFa2iGKo42lA5zGcaCy6SJ8b/LfcmOOvQTJQRJ1ap8tXqnT5rn
0yNWk02oNXag+J83TPKIrdmHKGkCUyRtRk5lqq0lTGhNmx+LYHChoi8d4pvoIEn+ylXHfesVezyv
S2mBiWtn8/wvw3f68opC4IWWh+tsQKPDFlaz1bbq97ZmnVwLPWaOpYunwPmV4TEMtCd+HAiAer4o
GwT70ioyMk3l3SDFuqeeSL2D/5ySp2bE1Kse+iQl/D75YoVHhMqeOdxLz4NmvbChChz83jtdWp/r
ug+r0YwgniUn9/HvkDcu6njRpLTeTXfWXfUaVM1olr7i9NZctNFY2B5MB6SXg4RKi5IxgzEiiZJE
ROqr5In8aeTL6Ni2Ux3XO8v/Q2V1bkbni/1tiu1jutXe7AFnRYoY3HLC+VKP4cqAsSZgOH9BQqwK
zKWWdXTgj2dXPKeHe1Ghxju64B0hDWTmF6Wld/GqUAB+WFolaKIMCAn+eGzbGHNZGdioiHgxXYq8
0+fI54sLTuzxSyoO5E/yx3fxU0wlYY202Nxtus1yz0nYAF8yWmyMiJ65GfwadzA60jI+cHjNbfJS
Tdslf70g3XeWKwjsyDRDnDxkUDJpVePcAbMM+WiEvfeoNbrjRuEHl3maI8HcAXBCL4Ym55VWXVwZ
5moLmoBsmmB49dZlm9jwP0HEVv2HbdpcnLIZNfEjeatEjsxQ3gBPSZ5VUdb5Dr69jHpY0fWY9rI8
ROQKCL2PiSEyMYVm0dw1zZZCGFoNpcqGNgGNpHG7xjeZNgfM2D0vEs/ucbq2z60ZtCBw1YQObxpU
qJU0WN5L08SzTznIyroTjK49bLobhLmUP7EkQu7Otj8sF82HZxg1/nlaHDw8t1z4A+GCPyRjYGhr
vWDMpvedFdZ2vfDym5qjuWttAshF/Jztu/Gpy3Y8ueaR0VfjUkZNUxItKrpm5c5Mr5PmGS4phCs9
SFbGzz7s/ukb7Lk9FhwKdfjnWtbymB40xJFlsgt8vCz0rtUWNKYzfFp+vHnBD391fr9bqluAhpev
DZeEgHADSsTKOn7dDHFtpZOI6FoiIJGyzkkoRHdw+7OoTm8S+y4Jcr/dX79GAPWP7fpRyngXyNj8
VMr+WQ5dSonT+0BQXXt1ViqqtXJi1QapJ0xblYIGG1vmSldC8a3XBH3nFLuCuqhE35MPbeqPc9qE
C/mL9HpLQehBJdQ4s3l8EIFLzqhTULr01T9JkdtWpcVLzsuLtHE84gEEmKEInylec6GvxOfG28pl
J0SB5TV70yiT19jp6RuvgstPt1E0qbeGyVNCsf8dlEwBtNkYB24ceqGVuwo03g0zoM+gh2AzIdax
OLmNmu8Y62uOyWzFFcBJ8iKRpE/UUF0vXFpQfk72JL/KCTSLBxlGR3itXrzhg01zTvAs5b5LpIj4
yEALlVEIsBtVmX3KsRpo8MLG2MYd1mhQrgqb54zMmTJ11rIchAOcrFNXcqTmCcqb+4YpAjpEcFRO
epC1X2inVfBH6b6yHjxpwrV1LAWYB+cUHxJJ/2zdzr/tS1JI/xv+rwyana4Zyt203UP+rRLliA8B
vvy/gc6ilsn5clyH+2mDQvSSaSER4VdnWUZ2Vdeu41U98XM14wDlHE3+5QkW8wM8jsi6Qxj9psql
0kmJ/DlureBCqJmB0tP2W3B3yudBlvwrQGHNrH6Y8YJ9mpJQ/Qqrl9Is3FnoF5Of3vLX/QDaPkTt
PL20DQkMXu3ZWMuBlOxUozebP4x2EEpyRdlpNxwudjeGCOgP+LvVNRwf969GQQQE5G860daljNKj
PTupYeavb6egtCoRCplzyio+L3okjIJ5+cwlwDefeqGd+9DHcGlOF11dQ6+QmyVyKXhEPotyYAys
y/nuCEDshGxca4aWhPj1hDKNDHQCZu6IsVt2B8m80tl9Vo02PwFnHOlmvlWeebp4GtD+w5IWmmMB
qCaLRpdfQv6zVL0t/iUwMymUGF91+rDugsvQlMV/NO7SEY+PuMIIFt3NcXPp00tzN89h/3mwkMSd
nCqdRp0q7TR4Wy+Ean7+HKH/0KDIg5P3CFLEZkAPvTlktO+6lhkiS8W47KxBxqU+yUtPNDEi2C/A
MImTYfGAXIBJuz0dzmfdFAjFlFk5tMA+dv868TZ/kXmyVAe/iY8WBEthyoU/yJrkmR3tcClSZ6rg
yzwphbHAwAYMr/LramJZX0JvDfMvxaAGIhRiXXDb6y90qEFsiRHuTSoV/JJkXM4GH9E6nKmPPXjq
5ov1KPyKrd/HbLpI1s3CltLhmSttQENErveSP3scmn+J+njMV0i8tsbrYdN3+rQDlwlK8DbfHJSi
nFBafG18P2KI0CVqtfn2aS5VMqPT6j0NaOXuSrvHdpfppcDS/uT1Oj2ENzbhbp2a6+HvlchMpmC2
51x8WcxqHBf82d5UnMtSVhOGS2cuqCvXnfeRqp7/WtM9s/bA/uXqDdqvBshzBjMDeba3U7A/+65B
OaDLTBmQMp0Bdp4LrB/htxFzbjduTI40LCPiG3tNak5bkxB8/KndOAJ+7YiTeTr+4E7SdmyF7EeT
OzWQny6D2Q6+yG+0azfl4rt3OCrxCuwhN6gR48dCHNYJT8b7DawACmsWHVY84POjq95jaDj54iyj
ImKNe4uTS+njerdrEDLIs6IQI+8Lct/29Oq1SAzcmeNBbJi0DCXnv9w4UdrE1/otGDCm9/Cahbe/
fw+Qpz7tsue04f1DZfziR4vSUuDra4Hz5cxrNVZpz0FucwffFuqCufKE5JkSFiprvdvXe/uqfmcA
H6XpIaAdBD/s7is8Aj0eoMEsB/0iQtLq2LXXlY4P99uzA8bwMF3Pv+/5GbkqUKvdUQLykkk65wa2
AuFs7njNNDK0L1LcN8xNKZ03klZXO11ws+zJe/rV42kxf9uTOqgOa3Es6AMb4iBuQ6lMO5hP2O1X
XTFLcU52ilTkTLVILtRkkp3NFr5F1JrulTXC0ojFMR4zr/YX+3cwLf8+QIKHeDCbEeXk5Q4nnGrv
CEV/26k6tAu54WoAo2OFYBS2tdhtBoFWerAs8YC1xehaq4c4xLSh1dQ9AMO1zD8FGilL6/MvqPHP
/3Wu+Wtsapp7csyJpegpkKbdEl3eIEHSabzzj63emKs8jDH8s+KKfGCs6t1UdM6wE6daYalQPwAB
N9swmNhCw6tqL0jiuurUzQFMD/o3ht5FquPAOLTVWCCxk1Yl9JcC9shFf4hGEHnixL4MOqM8QL/M
uUi6jZ95TymJWnRaKhUkwTTaeCtg0EWeGq/8ZAwGEuSB4qPTZM1I6FOjL/U4ZBrCj4AsVP2iqT3R
msBUltcEOZ5VUFCrAiobKGXIt3sVBN6H7tJAMheL1RK4EPwB2avLQWHOOFekZskYF5ci8jbhJ5gT
bM31sXd2TTNTz9QJHFyKVxTi9KK220WbPRDLEY+CXHjQbVphGIJqTZefQbFVzeGHzC76gifpAh0G
Sh38hUqFCl2nDxOTSktZ2jpnA4wApmKv7Vv8FV6iK88atGI1hYZKDIZ7jUIIVdxD9spjlw080KZ8
zLs/5yvog0o4LElN3leDMFp/SjYPspBX9dB9rB173Wy377uZcVnp50YVlmLbhf8cmlIf6KOJsrKM
apz+1FWtAP/r37H8ma4NOh8/VJNHKQEgTOwR6pPLGIujREEGuDuisi4xxeY4UsAKfzVVfHIOpm1F
fotOKFW/rYg0Ifh8uPVg4GcmBpXQuslLs7+fkzJpF6FXZNu49fEqLp0TarYk0RQYJ7KhvWulAAXf
GDByWlqTEByhRPQ2c/L5XLLBVasf33oyDrKEmzs/74pCigB9D3XwoE1FBmrWzEhL82q9YmZGDD3o
MP3n9MWjPACrCXs54azHGyoi+G92UzLdybPkPtTwxF1acnFn1jF1C8AacWTpkeKbIEZ0XAEStAeG
PstxNh79C+Y5DzFvd/j1J7FtYg9GZxA91NUiTWjEEZqr3KTycJG0LZPQKGgWSCJ8b2FZzD3YGRTw
QYzzr9MljcpwRNgU84XvojJYkLdnW3Kvol0qb1C4NINYbR8HQYHvUl8ZLHmyMBIDjwHv8KyIy388
uAwGUEnTlYdNhW50h8H2yxB89OmY9NhE2FUZCmpbZEi/MHyh1sWD7Eoi/vD5IvWCMU/v6PywqJkX
5Uxbr+C6UDEr/5PnqeRfCPvLk0Z+v2jyFgblKnP383u9f/UP06DsX9ACGI6rRG1sfEDPcSP4HES3
JPocmcGCS9r8JzIs3aglGfpqg1uOVqYqpVY+nnEcEQSsgsVi46SscrL60KwpvxKmN9GW3ymIMOo7
R1RJlQs6SsPnMWpm5AOXuaQUXG4eGGdhd8n9HjR9CbscQ5IFMVIkXMIP9q0u6V9JiwwPWFuEMdzA
ipLDOqtAsVgkFJYFBTyJ9dyafnaem+IM4ZryRGPMVgeCpyw0qVYwigZIurk1dsdPhaPuhrnVzKU/
i5NfDZLdApmM3DjLJv1K1TSvsLp1u1p8dl2/iphxXCsisMNc0c1e5MSuo21FJOFTJ0M7UE4+nm1z
i2JzCTkWrxlL3/OarHwPIbsBR6McK2k5Df24b8URsFjI2ZgAnyz40ZnCrm/zqp4CvgYTZN+WBw0O
pgjaiiMpai3e73zhHbBGtmgtAeU5OI6R6TNyH39hDr2ANV54ESBWFrZGu5CU4CSA0rF51pl5xm4f
Vh2vQUheBX5osTFOrrm1viq/iw5ySzj1NGJzvT+BWXwfpa9Tps2XzrVciO1ImxTBiZXA4KLjlva7
439BSm7Slrvka2ufcmDNAPXNDmwoZOChMpNkCiF+RAOH+li2pxl2H8br/rqR3z0lwSZZtXeAGlg6
/Suo9b+i+nUp+dw2csqPTjGR9cv4XplutznrCUfTs9b1wo89AiOcDGRzgjqcrn+G7qV8+3MunM1j
2iThLYzcHxGP6OheiGbbV6AwZt3V7D4mADWvPRx6cCIe4MRp9HuwJ7G0obFXuotyNVkYiP70JMPV
k3kpKY9RaKUrIKVXozzKthUeYAA82ellvYDsLhUidtoJtOOC+o1Mzr9ptlUZL+dFWa+MVaCGZzdK
LcuZ/wlJpPAFBCCzl3F0xIhmG/TPThdpmh+Psf2FC23R2rQvN6TzB0wnkqPCS1AtRKDU74Q3/0BU
uTWG3t5Dq+WsdEr6EpxXI2XsDSaRIoBu7VN5XVR+MTve7Ag4U1YHh7BThsLTaYA38KUF9V0mcp1Z
kYsLtX4hiX602QUoOkqLb9fp7obr8WnG34YDCPotWvc2gyXUvGYyqQTcCUb3zVHXjFsZHSu8Kf4g
pJbUHWvNAAc/6/3rAgu7iDsJ439JpyURSeGPJNiLIk54Yql4QgdJzrGXB3mP0XFSk7FzJri4/9bf
Ohb/nuPt2b5+ciAVhAgSB/x3dfSYYPOcKbJdkEjdUWF+K3wAV4KOEF3ZlfXPymUT+8gGEXFwpe3K
nD1r22JmMGnqHH1zZ3nWei3XRB/uONZyMkVK6B/syQuiNed/W9vsJBtYqsdJRdQ51OfubkaC+w3+
D1ZQ5t4Wq78i0cgBleOSr1dbm1aVOG9AoZbb7BLCL1XF6s76rzROGhq/KMZHW1kBJL+GOKdLMaii
vEmCSpl19ZZtxzJ9CDyz449sPw/8dBT7SJbn5zKcZ5ynqGSGZOeBxRSy+EKYQ3xD5qJldU9n7+u5
9B1Zg960PeejLlgJh63mLajYKf+OHgx3GDLUbjI4KUhcdrYRC3BrxrggOORCV/11TiwzaUkBWJXN
eiQ3ynjCLAIYEyfot6A72xDXaeWLT+sOmaMy0VNiD1Xsx4/MTP/Gthtm5oInFActpQkuN+JnMhnT
4pIEMpLCpBj67XMvHpQZXovOp7NPyg0ZgSMX5EilA4EAD6M3TpeTflMovVBbhGa+AC/VE3PkuRmu
qncINtYv2OhvHoDNhIXjRHN870ckUVWaxjmLQC9jMnR3NtFvJ1JWjfG+TOYpXDTjHf7UKhe/L36i
TVv/EEz8N81zCAhgShecBX0OdaEM1hckB4pabs73TlYizXxRCsTNu2Wjmvp5OStTO5XKY9XxYvze
RrzjAYyeFIr8phnOY4axkg1ASRqn+kQd1v71OYCrf5sjqBgnC4/8BizDJsCnKMMaCgaJ/kbw+oLZ
xCphpE0jTKJQ0D1wFqPkVJ7NV6BZNgyKy4you1MI+ZG1ZjhHJ35eXoTRv7plfVSWrzhTb67vNuG/
PAX4xg4V2bTEFY8g70DxLKHRHnCv0E9BKNtKQ3+FzzrL7G1gVtEF6tt95GuhOm2imZP2z6/BjUNq
vJr5lPGi/ag3FC+W2/OtWIv2sdjmTrtPHOuS0g/o9xl64eZw1NHXc2UteZUxn7hoHXjjlLCizNk3
SEoTLl4tDcnRzXJ9tUDcb8ay3ACgEr6/9lJ99zPeZYtgBia1lpBg3P3tEpFDjrNowlpaJlGnC84J
31M0rk/GbedGVk3UEW8/RLa9bpw8gDZVN+yF6peL9V0PNIcRnsA96z08XrztOLzSSj6cYJ3oX+5E
VAenLocV0orh0dTqmwFfe2IACHZNJIMFC6f/Jtf03UqqwJv7nVIKwDTjilG4YhRtNgjZeafkzjjy
0jpu+4TEhd5n6AIw5IThfv2haBaOl4lmEGgDflD6C+WHVQya9HFUeYYPsTVFYsFqOMWhWIHgoqCy
3MOZdQfsFQy1OswpWCAYH5OMzenJsapwxQB3NCbnigs0KgraRstEZuUrgl9557o51y8w1PDD5WWB
MV/5sURv1fc/xKurJe4EokKk9mgHxh4BFcBhXTrTLzJDL3XQVQnLXkd1kg0z3CNQNkHelwlwu9qh
nhksFi6Jixxg2r4XEphKowuCYqz4TgZ+yLh4I/HrjcswCqBebgzeaxQAA+Ba4K4ZmdxyjZ0OuhJD
yUktvhQOVkAA3ZzGvjMb83bpL2DCekHMSiRVrEk1z+/D4APgzY4A8oaSXzsH7BzMQwwA84Ks23Zf
kkdIV2S6x7Kd8UfXXTGUrYN+b6jraHcfXZ2lNP/OHsf2Udfq7YrETSTVqcAtk+AwF7n0SctN7dAq
s+jUoqKD57usfAUUD2g4KYM6LNTmJhloILwVHDVPZEa/QfHFWI6lFGosVJP1kOt/9qzZlGaddm9K
cFHtOJN1UrOoII1kNMyRdEhWf/j7paAgElloOoKu+cwSQUrcFz16msRtRwfLk6moiLNo/qpGXkoG
uhov8ruNJ6jKGyfVJnDfhlkqiQ/C8xM03IxMtKGftfcv5bwMKWMK5RalyNMNkBagqCMFGRqGo9Za
LaUiPnIyf5vnGV5vGOmqQSEEnwMTQm6q8sYGsYS03XIAHclM3HJj72r59NinV9tB6IUxa43EECxL
TV5I+ycwozz+CAYUzcMwiofoAtYMZ/oEM47x5TRxYfZa+TavHrTrvYqtKdruxhlvmjtrtGNr17fY
NHV11J+svxAWcEs3oQn0jloTzESA1xZ0n4jkRo+XD7FhRiuRfYxSFhxKWfYzOaYh8F1WZqQTU7sc
vsLIsX/pjBZFGtmY1y6LWdVFnlmHjNqjd//wdUbU262/aXEHEw0Da4gBW71zvhOlX/84GKxPghP1
iW36w57pFARUY/ag49GPqE9dfdRuU6Uxm/KFtJtI8Vj33PW7g9vx1yUHOdjwZGnuiOjAnGfbpM+e
D4So0Sf2tJmaskNN3Hg7trrak/pzLgRHALat0JsVe9hoZXftTLrYVWtEeqAJXMjM8BND1Xu0jzKz
TUL2+7KiMlgeItdzOrPbPle4N0LPlTTXaLirVDIIJ1VH06t8lu+LGCLjFVCdgBAY/+PsGawTgGRU
0zy9yNu2t1LfQ0tkyOyb4/qWn40rT5k0MlJun1ULMFAKAsSO+WLZEnmjXiPFHWgDTje3rlywQnGK
hR7H5Z+k6AuxztlJWdc1PKdaAKWBgfZh+0ItcDuSLr8A8sWN4NoCusGjOEXstfZvtO8vZoyjFaMx
WaUTUi6Rt+7Lj6CGgfQdcdSrPfo3HAeHafT8sXK0oBoOqzCag8Tcy3P0+dA2HAUvYeHPzKxTkgEa
KZCqjveJqCxlwg6P/CxgzdKXYss6ZRoUCtmdQYJIed3bgm1zujfcMGsCy/OQ4sO+oQWgFKjGZ0Xi
b2xB+fTLvipGwqbPM/4QqQJFUBE2FExvjUbjJdF/kjD7FDoyCsf/rSMOK/GUHckyJIQefXdF/MWT
D/o02Qz10F4bjXMQwl0337VZwC0Pu8eA+5IFyqednL3okvfEJB+IBNHTTg7el7jelAwCMfTgdG8n
AbZeKtuU900tvwfTwED4VXKZpr/Ka8wf6xVCvxXdKbj+oenkmwd7gNeFdRtRW/51Sq7ZBw6HT4vJ
VQuHgAg0Ip30ZY0qSO4/exYUnP1kOzsQKdIUX3Me8NkvJuAzxkOrJDWo0rja9nqDK3u35NpNAwHn
UHiQwP6rbbqiC1a9BMNHilNgWRRs/5GZQOQRX+e1d8/d5H+++NCbqKBz/F99hapMDWTgt685POt/
xcZQAXs+mI5B1kqILnTysCvsK1SH//RbI8MffFdBQNS/f/KHA4VymLFW/OkbS3Cq7OQNosXhALQV
WannN96Fw2yF3UPT4TfF2YVFiSRt49GE25TjRDuc+LS1yru37TEs+nA8+OORBsf3Q7ZsnvwsVc1p
uopY19dL+jp4GmhsbbNZ6muxPr434wNKhbKVYuuA3ZcaYkCfamYikGhRupC1eD2ud8Ua6s466CEx
tN+EF6pMXRV0qttAaYVaVdRxJiFAcUZYUvQiIQwYilDw3cqicF7KYD8DbaDhZW8VTKGI5b/H1lMU
ASI8T9YTIIJcNUOI74LOT1cQCqjfQQ0awFIQnUVukgQ4BVRj+2e3TmFGdz/mj8Vy4RjY+biw63Tz
Jjz4h8YgmpC+dRvh3nUo3EcA7J6JjGQkwux6Jb+b172sEuWOJxHCBqmEXrrcn+9htALBUBgGuN2c
qFBz9ZOTrOI0/gHVSRT9ORRJS0NbNSeDh/dwpC7slUdmCHkBRZo5/Nyb/gnJJDvYk305WGoctuoC
/scYjTHix7whIQl5whZ8JsCq7WuRVZ9CRKBxniq9JYuX8789fb8FoiprFQuFLcTKy+knGvKeYb3D
75VZHkKlLik7DQV8XGXQGa63BYvIZNSDLpPaaYOJAIoVUUfSQFq7ACHqHdo+SCUPIcFlAOuyJFPe
CAP/XYxRPcWc3fDfOklh1k94O0zAlaPyo+ozSjMp5FAuQXn90pzp0P/HDJL0BmFur2A7X2HOi3Dy
TyAtryP/59teNICE8zGmU+urVBYIjQx7A2IdsbrdLi2bZLAGl8Lfve/t1Azwig7TRcSqsBersifx
3gDO1+t6JJGMAYmcvoFb9hgamMjjTkNIWmuyBJ8m7WOa3Ox9iT5PVGk1RPmxOnVI6jMdPVL5d7U7
NlkY1naiCGUXND+nt9WpbOlaWNSS2TI6+MJKw8XBncFPLwyr+lXbn2w32nAcsrwx+UdCtMfC7GLs
z7cawM/YxcokR0cUm5IvS583zUzaRdgv6DwToSyHY6xLuFnib+ZXMR52HwIEq2O4dEP4Ylmn+XHs
ezJiG+k2wtRdeOVGPwBrACeP5SXs3qM+HMp+IUSHUTkWE49av84VB4FHRvD4XQ58FMi5xdEW9LqT
kVbHaehXsgLpMynxrD2Fv4MaeLoDC6TXdiQGcv0EymEaVHC1TXiTZXeW013WXNIbNsr3BHV3P7wQ
KiZ1zUxcAbVQQscjf5qbr4YUfmc8yx2qJJjxzYUOcC5/G6GM6bqK1LXmA+RfJ1mP9lIarDMdicHD
Y730P4Xc3xVM9btcfHJkGr/H/lxFOuTSM6tyiYGNJnYzMCG6Zpbmbtf8qyz8oDKLsiq2Vy+yDHJz
DRg/sSe6IY9s9AGQTWdH2ezlSJCtaxh9Hf7sstkfe6d0Mqp9LEj2yo/ElFVmH1+B54tGgwqupyYk
8sXzLWNL3TXOTYM7Y5Vh7MKexQO/9SewDDdLg8r9XvXBVJOvaCP+lxzBW8s9o4+FnHPD76X0iV2B
+W/Tsye9psw51Lw48Bs0/hiH9O28dbD0bGe8apOjkaUC5laC7YSYOin7Eui/dxLDZYmOBf92lB53
q04K8iyiaA2GMOdGCv51zigBarSp7Nft6j3jghbLrhfKxnKGwrmsYxfbvc2+9AeBOjXlyC7Fj21K
3BDQZs0KZ6URxr1B9cDePKcBNb2JNuha1+jrhBvhj29DVWYhRCmJgB3WDnYOJ7YQ12xuobx4Xxd6
vjovPZcmb8UomMaEzALNz168Zb7QBVMdaolK8SKZon81rI7iHErahTv39XQ/5DBDXI9m2c5xuz4a
oqa/ACOmSxxwRMIRzqWgHOFB+Pwyz3vQum+7nPWzjW2/+2eM3BSYPwnL1C96WKRvxvWjstqNRRW5
s4r/GppnAPPV/Uq+IabnjeMD9cbW8XqOnefK1/hYeL9zHL8WuBSBQj+ZwfttrcID20Uf8O1LhZGp
xlXGIXmzklcHOkqi41dIeq3m98xBhn2QJgrGnwsM89tUivheTinlp5ZejtXt6bSsnRareCdPuKcM
2oAK2yPJHsurcQZO59LsIII8QWkmxrwnilNt4xpbTWcB647jgzlQXJkW1+xgTytuS1/J+qfxZNeI
j74MZtJwfIphIM7Izjzw0XKRn6yi3W5f6nLvocPAxQDLmYjA9wpp1XdOLcmGnw3eWRUtgHibAFNF
euLBe6HYPkQ3Xbd2p/PKarfFyI6ehNB5lYl+Zk9cfBETB9bMVKNrXIXNY74y2KR4QiQf8lQqSkdT
3xpsfWeBDhwYsVnbnBji8l94FAUPRz0Pd8vGDAUFflpmL+75Na8pNqYOyvqT/jTVU2WLAAU8kfHU
q8+HZ7HUQ/HHNq0gX+dAqYxiC9wV/YySHScMHeyZaNkwO8kY7NZJ31Zxr6lzsLwJZPLBP3W8+GQ/
JV6MNRaPHUqxYYQDde9L8VP4U+F7JjCL0SQTsEOXyTg9Hw9rbRiRjeWwsh5aSVJcE4GPI2pVwBHB
hQ3LuZnWpCOle6NXRZYyLreclTuc7QOILN/cRQQrsIzWQf6gqI8P/DUAjU2dxVBA4WzATwPYo63d
Jq01ZinsNkuiSkcSnxTgr4D+4ZVTsTFkBJ9InCd6ieZU28NoJ8pxmJpNlJtJ9Ujm8cLc69GotexI
NFDlTUHiJ8brlD1so195i4s00tck4/1ms7MUVb5A5NDVmxlqneEKh194zQwD/6YAWbACAc0YQNHK
4jCk36m5c/VDDKAuAGS9oA4ftsTwm1x4O1Acyeb9mZUJHweyv2Kb/tjjI844nRZea4fiRXkYq/hc
K33lG8zQquY6C3iN1UatBMWBMRyhx2YW29MtdfI1xDNJ7gDLdN8CwtyLP60CxRgl0naO1MevefMU
o7O2Zks40WTnOcJaNPQL+iUtHNakiQLH1sbtNK+KNnckpryXHeOPBkDFFzc9daUYlI0qKd6jawo0
21/+JsdwbPuxiz7mXzwzvg4BynINctYN/uN7MXtg2Ge4HmUGhYS3UF5Z5ChUB19d7S/d5VjpFasf
W5WYlmojTyHa1JUpNltg4a3kASR0bGJSmAEX5Fdgl1tgxbbKhTs/HY+dakrBJgZ7ChlVH1YSn78i
lF89GHKqzKyHPCuh/Af4p02ijNbJX/tdAuQzXJ0GzfEt3bscMFN6mVYSbanx8PtwIRV2V7YbgdQa
ikIVTM/Lj/Hmqd/xQDVGAZNGLPMpZyrersQB3pCjYuh57MnU+T3kOt6/ej+ANC+9xIW4iCyWSYPl
rEMh72UvpLJ2E4iWpFH2dT09LWlOcmHqxBVjtH5gWggUepUjot3ieI82mThJnnx5RScdccZkLq5I
dXbpJTjD701k22/544rSSGMJKOjRUfVVmVoRMaUQxteqFYWPx8f5ILfOWkce7J3rX2LaS+nVPxnq
r2JIFaj/SGLEs5dtkKdvZtUGe7VJGVC+DwSiPZEgJ+fmR/HkuQhNgZ6Sd3SbNIf5dTnkXAiCjXg3
WbEjE+O6FV6qE87ZmSYd2wudQKHfNsRSKDme9OH+N6Xb5JrVswJCblexX33MlRcAj2hpy3bomtHM
iYzlh92enwNh+h/S1+L7tGDkshq4EnpmyZfbbtBwnmf2Wg+EEpWW9+8WWAzXX96rSbQbUvYBLmIY
bGrXnhPB4m0AFq4MCwNzxSX4xa7n/sNGtk1S/44c4xi1kXm0Jz5ckoslkSQdF+7QnSjlP/Efwgjk
l7arRRnXDCr65wZEpJkOOHciLEO4DB9ziUfcwEXQRZ5adt+H1s+r9D5ovtAx5RlZc8pDpf6uiKft
DrFGQ3YFKXEUiBc639YdPme3dDpi2uYzVA4SShZWKPJ0zZrcgN9nsoc6NjiYmycCV6Met1JJ8LMY
itBNfoeLe3nPQjYi1cO2C1gyMkLvDMcJkv6Mv5qXbkYZrWAbsZntabkXQDMHUC7g6AePdkjoTwsd
Tvt11QhOGGLWzFkkM9oF3pWD6awPCIhDltgZqMnAcrYz72UUzPk64YmBViufSNhwk3CSxmrtqYdk
djnGMhM/WF6uxAWxDMqEnpI0c62YnoQD9PeRCxD0NkofLNWJxGLj5S4/ItMXf7yNhqxlsO9ZIIui
q8IWkxekfbQ+tAFi3UMyxJG31fdbJSh8BchrLUStsPtDNe4zY6vxxpQC5YoZ9CL53cS7rvCot8f6
Jd9mW06sVZfplh5U4sFMVqJf4uYmjDZ6UhUgBS9FiVeHR5y++A41REvSY6LTCJXOX8nYhoMslDeZ
XZbqjLmHHolLWWd71vSW6ojPvmvpWv0OXPvXv0u+ucosnxeBxVx5SZU63UdsY7bNOq0ku29YyWHR
mGcoMfE7caVX7aGZ+u78s9gc64WQapecy0d4+JdjRZNX8KaXUYxqrmqRH2aiQUmUXHmOzGmYwYkh
VZdJ0UyC0IvmXg5XlOJzQfNg5Ah/VderkwzMgUxjDSmQ/vL1Q23JcdG8F+8b/ts0ObnxLp6x5RwC
1UlX4ofNmoYEyPOtOotkzA32jl96/0o+VBpmgXw3ST4uN3mI1bBqE7PNowgrzwnruavoLYpnPM5k
9Mb293c++BSUFvH9xh6rU79KTuPDTLJ7wxMNWHjls1MeyfEHpGIQ5DM1zINIac8Nd8D57DWgwgTZ
Jl5O27bTAZPuE0Oqm9h64MRKG4qKuV+dsEbcDhllG7tHjXR2sa9UbYwH2rvDBtrgZjdjx0JbceYG
M1ocNW0ZDjnY4GbmEKayzuxb4G9TCEpEmGAMPUbykM1t/831FFjT+rWWltxO0bm+An46eo7ZPaX4
ij6oBhsRtm9SiLniB+tw6WAntcJ35fzxTRwpnt02WiBmR3jxZO4a81GNJW9jZ/bzkEhvXI5G5pVV
rDghW2AHa1MxnvMSTvc2Sh9M39UTbYQNr52P2PGwuTv71jh8b67OKnbAomfr2IcqCpDqNWVcBoa1
28NV6WubRccLQ1soho/uIdMHQ66ke895vNji+mSrQxvyQmWiwQ8OQIuqD1zCve8z4WpepxusyRGP
ow+qSswrT/Ia9k97Zwc4tMZznrXkcSoLF+oiSmYeE34qxAZAUCRaf2BI+QXlMM7V1wJP2RobeIEf
cWrYtPu9P3CG4X/L2GMQoJLApDWXtATGV+cUEuaxnNpIvQaLjD3LingBJs5rXajR6/VLlC1/jDgk
8EMiEGY5fwh9L3Q0RbXUJyiOOXTYE9tXB2RPz2lux0JRGfAVebUwc6nA6qRaBMFCTXZgoskSFMQw
zP7BLf1YRZUNFJCMdkZ3shKhfEnc8ZWkMUOT1WxSKhxLlQkmHlKw6s21920kqaX0Izbg/QiONHgD
HwJqB93Qrz3lDRFUguVi8SZ15d95+etsee/BzHXxvycMBMkNine8Ra4YBW5X1JG1/bCjJPBn8BsT
25umt/FGsLD0Ag3YPVVTHKkjrWaTgN9NjOrtPLzIMkLSELcp5mP/hhIjiAJrSf+Bd6zOu37yzgl7
4fHwFMBVsqy6U5uEfhQmkHQkxxBbee6WBnNK+KWCxwmN7FPqSULelk44/54nEgEhz9h3hWxMROas
RcBTyoddFlTAgrAcmNBOu0S1y7iWAwlTddc/YQEPhADvn4EO4q1iYaVKn8XutiIzizzfWz9Nsyxx
81f2D01lDbMOUVaKIA4DlIiBt1L1uY1SnZ1pdKc5cCVKcZBLdGcAWAeI7dUUbPXuRPNUsVksog4y
jtCOMzTl6mgwJM3q8Kt+OyeKs1Pog9YEhYgxgFDpp8a4oQueZlgJj20T4nmU+jr+muacJys7yqqO
EPTRAFo4Zf06wK9Yaljwf6/X4BKxrfhHZhEKayCz3yB/3TBssfWnnF8BfNdULML0/UDv0jT9ZL8z
Gj9yf/+fR73HHPMPQ6B+95hoiBR4qkV8QojghhSdvg2/yN6jj9H7Hk0XPmM47mNhsXeR0+42ztw9
d9DrqYUYJAOGjZQP0NqH1Y5d2AbHmgVEgUbhDfdKvvBxiWISfCiXOtQi2mmit7wyDjWD8oiC1Isc
GW5eVYEgZ8W1CaAQB+ALgJdTleCucp9uvL1Nca6xS1nsJ5KKu+3MJf46q/mBoVLUsWaH0y1WLFGl
UyCI1ZIYJalOj4KcFNCfv6zc9bgXuHxZ7R1uTjnOoK5q+XdtW1ghUGKjnPdz5V7QCzkRXNgepAou
dX42l21axtV4W+s/gi9YC+qY43FIusN6TmOBYsigBPyBMd31iK35OIY20krgjP6RqvU1Ci6Zp/Ml
pgEJfV6643W9mivVUiXF+OO5W0GEwB+t357BAj+qq8bqMOEgBvFsU9CWXyXSVVziM4UqQO6Gcd29
j8Tvid1gGcRCSvYimcXh30AusHRCj64Ard45B7xtkiE3CWjQHVX5t161IG7O4Qrzb3L29fCSKxze
9t9PDr4nK2lLrTS8zZOI1fQfLaNi3gXBCkIrwLjNDg8Y3EPqoX32tSdrMeYItHfOWeyldvwvS7ze
nD6MVWpvmwUGu0076+/Jb93bwbLKrFTDbw4gxz9FnxQkXLIhJ+TYbaaZQQbRq1e5BBCELqN5Fz94
ETKbuJ1YmvLw5Wbmz5CRBVZnRS5laOOCj0mdC3HexF2SSpBuxkeF/EDGUwaNTzquc7aSkyjQV21u
2mO+pQ7ZGnUFmzUaAsBfc85jaeFxA0g9yuQMJ/CX3+YAWOmxYdptxshL/XK3Yg4JmKnD69ZTQCgE
dLToJJ3exnzshQlkeIClPnMloE59PX4YskCGoWSbIgtdVC+lSw6RS+RJyVq0r4D3mSUiUzUrnAtJ
bkADL3zQ6OkqfHl6pJ2OV/f2zkDovSfiUsDL4kCDp/J2ny5fK98rltueirbrC9O5SM0Rjc/12wdQ
hhpgnGi56a3AW+8iP2cjRQItTYaL7EQWh3VqvaObSvo3LBJsxIUgObk2p/YJ3GAAqzuye2GjR4yw
n2xj/2cit6K2X/ay/+8wz0hQqQxmky2jZab/2Ye3yzDhDdXYo4ZOFRMZiga4lYn6ewaA/16VgVkb
QlFdj8R5wvWnPwzG09GqKrKwjLBKNBlBUdwuQKztb4joElYc6KheADN3AB6VGO+M2Ls64/A7B7HT
ev5LTHHTkPmtLa1p0+5kT9ubY5JuZTDimeKD6XhEnotmhmplvKfSXeEcUzv31d7IXBuOewsX0CeA
CC5/x7wWGjyxWV6NA86DrMptoDrZlWogzEdN/W1Jm235XYj1IrLkRlPf5IF6xY+Q6uOXWIY2oMmk
6xqYJhN4lXIWPyzbUFkDKWjZ82MVnZH8QRbFg0wjyI0846iDvRihJFQeK5rhLx2O7sY+8OUyxmgd
TWPSkwnczkodw+oV0yT3h+Rz9i+VXwRh804sUMuk4rZ3/0P98tjx4G+S0SaU713QKPuyffDYUjFk
kwUQYEDN1hml+1Us9IolRM5ejx4FR9hzu0KGif2Gl7VUdMZdHE+15CJ4INH8Gd/EhUcAFymDJmNz
C1Pm6zk8NALDLW+1gmdefvPmO+7muBzcurnuXI+fswwXGL6wG5iE6c4tKZzFf/9J7Qm4D0WDKWbh
rbs5ddpznkYAJyYpP0LNwPjK+1wOvT1ojbQS4+mVWptQQlpO02fzBoINgtBxE4T6L7eOoeDckRBH
j/pu/U7CcaHQPasM7nQQrAJlX7okJbYS8xiYkDI+Bj9wOHRWF4+ZgDscySg/6ExHQomjSKITuxv5
3zM35yO2+mryXSvUYqXw/qKV6I2h80pVsbOhkHTp40yfx0V5GBsnZxfnqIH1spYwkti7b8RN8tfi
xnZhqTgIi92aUnhKIiAkWWtflNV2BwAhtKj7fDO7UJ6uwJHBCeUHL8xgLu8w9S5vArcJ7m7pnrOJ
8zXe6PCq2MtgWjyeNCZ//a89jj2Qwbt8wNcdbMLJAf0M87m44KQ6GnTJZmzVaiaPaBUnsC6Ob3UH
npsOvATj/9JNWtE4HdYted5lUg+e8/aqcASvlVaGPMQb28dKctbmDYDbsrRzugygoMaNUd4NGGTz
ChrVAYYJaSYdSAIxMkeTorYlD1fb/WhuLJfFUxflqLjOf2KI0P8db4ynoSq8+zCwerQTSPIWTDQK
ay4mOr656rrZiJu+3jcjA6XUvtPlKdw0k70ChdNN5V1nc4cUW2IeeLTawXjoePJXT8kzRCv43xSX
7nB3glaDgSaoxYmnQSnu8p2/IISxZqn8d1vKuIijhwh9aQafsOh29UNHhT0lpJKcLMiBnHKq0eOd
K7CSgE90PglnkSm/UIGZWApb7hmABnGuenwNx7/RsqeY+ggXmYfdPaDuWxvjzcKZl/HmTF4GgsMS
i8ZAWNaJPFxDh2b5mXoZkk8AOVD5em8FchdlVn13rScI1+ahNXXncH9aA2iin2NOxzw8y6ouIDad
i95rtajex3HaCLIn5h9eiuy9ywGXUA76w3akQM7FXhAP3TYvT04ZTJc6Yp1qwUt4Q5QOJrzvXB8b
lUk1Vpwk6+tN94LvgGUv1Y5IX0gGNBm0XwEMuehdK0S18Q+rH+L3qX+PASBjmOWooCqsNLeqbzbG
bxQzAAnP1Y9t+thXx5EIbZHKb5HKxDwpEwOY/4bxChxVQf664i2Q4weR5EifG7OKJslpGuILlzqQ
I/7bgzjpuOMsa+JPTW2qCGf4orYI1bTh/Taag4g7RpOyw7M8/VlT3EEiLX5CQqIFGX+QrrwKFglp
UXkAPdmxXOu7TC2v5Q6Obh7AePTebkFlEMpOJuO58mluZg01vkL81/1EI7W3rbNbcRzbOGU/7/S+
YyO2jnA+PR3J3nCrQSQy5FZp4YXF2WZ+KQueQSzKl2t9KRJV+GVw5ZDCy8BoMKDtLekT4Ku11gkq
BYs/D50bHqBhifON5YDW/Iq0oCxHIIL7ZquBNyDKPxBSlVBdYjE0qQMbnKL6WEkK+vLdDsxdNETt
nkAvg+RhCU1fLmMPvFf5a39/8wjzdbGkY014T+zO7lqTcUV+RVBByOItpFUMEqZz6pTqdixN2SvP
do7gyjXROGjID5Wj22WDXkWUD1KMK8JG1u2Hulj73Y4egQYS6GYs8pVNryhp+iNQiVv9srus10JA
nWyfCjjfd7hgz2/TydzttdVRBHzHki6I3UPtx5M/5vfRqe4N6GFlUfohwHsfSvn4zCHQztxpwDQd
0cYc75ewN9O6Gw/gxaPetFPVfazyBc627iR/cYqqJE1Yy6iUc2PMxVXalHrPjp31wXmFFxlXYDju
Q73zTqHSsUxHqIqW/76fJMfM63uTLX59Q1A1Iip9CbuCy6HYIbesXpO11qcXIa99pX9aMeiLLETG
TYCvA2+S/1xUKKv9sBQ7Cxx2QOmJT4hYVjBzBn7BS2Pn1Ywh4acbjD2F/0lwzUbwEKlDrf9OmrRw
pvz/bP73NwMLi2xPojD9Oz7MqS40vQ2uopw77l5gK63PkRTx/+TN5hHWArSCBZxLVWQHIofQHrcr
pEwXFJHjfwvXupVVk57XTGk7Gv9q5mkDcGlDTLTWhWmPLCnQEotd/O4OiE8lEv2eK5pm+VUSornh
8jnpd60emjapJi9+1DrxH+KKn3O6qOv+5avCFCDCREo7ah6C7ZyDh6yFQ7PkKr/lH7VfUArPqjUh
uV9Vl4H+CJhKLwdg/bgTRNLsIy5MCf8ewFHkm0mE+GX3HRXHaiLzfMxtKUJw7WECOfuEBqqkSQeA
I0Yd8yrdLGAQGx2DDNpB+cMMd5xvtnD0CpxEFSgglSzeyaatXyVqt4J613kL7RT5cKpo7695Ayn/
cPliR9NZ+sLhumwaCV2R+vjlUODGbUrARPUuTCD54ZjgJUoXWlMlSo6znnuQMWambAMRqch8wnDP
ZYdGrA6c5zF78LXrNVub3NXbg5NMe0iYNXb8YUeif638ZHPCmu6LwM62DLUzLuE69Eqx4rtxwe9Q
2uPzoBKLNpmHab6wJ1kL9WQgCK3GYl8MBJ3CctogTDkYpCFCHHn/4uMIrQdwR/YjfmmYagNqOzL3
Emdhx57sjhmw6aO/5jkoPaxEYPaqZvt0d3Ikic8siUrKnKweuOXSqAmHu3nJaX5vyNLcPBe8Uf/S
MKoRWg+7cUJNOMgR7wMrcuby6569RrUgaPltTgbHU/c4ev3XSlGhJAkEp07PdfBk0z2vytL42bhl
UieG1V07ShYpdKtJS4si1pshJif6MR/ijpmtdamKgyJtjPIbU8agESTflzZ6UM2hC1q55kNn9nuG
g4mulL8u9MpNdKUZpUrzAfyvEQ9+NP8lBdQKAcyBJhQd0ehnLybWtOlhalFgw4DEnoPuERMewm3v
3/VJGM2kcT7SahdFmFmGpQ9ZZsjyLgTlKDx3/8IzEX08FBKde8eAMZ7fjSgc4aT8hI2IgXPBSccE
sDJFlVaLhHTO5dmdyEpkcGJqPonEQuu96lIqFTP3R0/8hQx7M8BEt3mxf/knjiRnpmiEvfYnI6rS
RnTgLJeLMMf1c7JsiEo3wvKW37SBwR7hVtIOtlI2w9xj58HZHa2nRh0gAEDMUa8gnxomLtA8LbM2
fXDhLz5s3NgQCr5a7iJMx4MrXoiFeNhvb+tlyfXxrG5u4K//+I5ErYsW21B3C0NLI/tXyAPeQuxB
BCJiQP9Qa+xyvC9HlVifKKgLW63CLA4bG4NPvEyXJ1A4PuuePvA2NyQO/fPGkAybDHqxOkrq9oT1
md9BtzHi05XPystaDpnmLOU2WnBYpEwmtyJ1B79LzrD9EbHmR3Y0P/ICPKgnETKGufVi/iB4zWPJ
iNsfGkIE9HlXqtDp/HNE8Ny96rJkYhJinJO1HxABMXirfvnJsV4eDAtIsAY/tQg91HNquakLA7Ym
p6hv6Tb5TLk3jAoXrKUvl1AdPv3VlLWZxwFcYmeYVf1amF0ZjJ27f/niWAXVcUi24/Yjd5IfOgIO
LOwhISFyYKdH4kr5G78amgD5ORNgordxO+klcb0aX7KDGuRG2GLSVZakEuOrluNkdVDzkxmipaDU
2sZ4OKCzmlG3cJghsHbtnOR395PORz28DU25lDhfCCN0zBahOHljOpEcGwXZMFWUQIga8Bw4+SjS
3MLUrHhj7b5QYUxU9ET+a+6z7iS9o6+bYj8ymzGvGpf6SU9/dvwXgKLxE/1MpTNQJRNUnW/yKl8Z
FRP2n9kClwzs9JAmzbr/Nl3tV3xJT6bIT0iRA3QNGrHSFJKbiZkFIlmzGYaIaNb0mMptOnEQ3lXb
PepFASF3BuFSZ6YURo2PJ4ILbTlFI/g0mX5uzV2gwFZojBw/XTvxmJgCUBpg1dh7q9/ICTcpldg8
QNFpPWojmAp7U/1Y/40XM/B1HU/Z+LropPW6edn8G4oJbbRqwvYezFAPlF+Ssrvokl/Ha6kUriUV
1SziaG4V/cVtRr4BtSWCFlk1svZxxDhM57VrAHvDlMPRFxyS+lMhrBdSv1ADM5pDWT9l6Ejx5oNQ
jRf66Nj/p81BrNN3kerdBAGS8EjP+kw6YGp3UKd+8qVf3jqSVbOJpyuZiYavYdEfb6RAxw2nfPwp
JY87vhYKUTPc966AxeIsq6HQEEl27f4XXMf3tyIfY+hd3Owu6l8RplMLGVavFUt4lE2Bv8aWClKq
RXkYy/FrdenJuEVBxDMcUxq0iVRqj5j/PuvjYdDiM0Uhn2epee3YmDsgFrfy99us+d+7YLBb4fwH
Q8dUzynBP77QbJ8IX3XrggsV8T/voHLH1qvNYbSxyb402TKNTodZEdlUympY8/wLqHTHBpVisybs
RGc/HwSQOhhbBXBh8Fa96f5f6wqLPifX2SE1QYiPeoGVlzm19jvI51KaH2IA80n5I3OzsopfbyvA
qQlujYCj/RuiQiSD+igBPLTElf3YRo8va3fss+BSGB7iMDuUM2Uli5k9kgs0LG15WHc5DMn/wYDE
uwcUBEoC/2L4mw7gUog0e3YaSh7OJKus5uuZqZu//5Sa0OvIAwzRJH7tuDnRg/CjzOQiEhzYnd5t
spo6T/dm4LY9VQXqT0M+jWW33PmccHYqyuBMIrj+p4np5TJGQNYZvzHlwknQNrEGC14WInfl2s9j
BLNX7jubQJ5RkU8WMiEJdxXGo3OKvgEnjoo8lz8S+bg7HiOhYnyTP+I6e2VUENJ0qD1dre1ZgT6H
CDWD9jfFDRdQbt9GMHXYY384qIyHpnC5QRf0ndXrX31saImC9HdAO3OSNkKZGxm7noMxGZ5R6Gpy
QeBAJtbskbe72mixkZFQMHFDY7Ri0CED9l8I09t63YVbM8PZ6isr0tGgn6DDkqfLmyzaj8hTr9Do
Ind5MGc4ppNHUXHc+7YKmUzjWImTfRCuOV/3bF9RCQGykEj5fONbi17jZr94d4OKWr5pTIiPBmLY
yyWy/HXdL2EWqSBkcI1JL6jOZRaHIGrHdz0tnt4H8ZV8Cwzs/yBz/Vs6eAbHT8TJARw+zhKw415d
JS42nvHOWmxBDD+DrNf4eB0I6xO0N1BXn4+C04h+6lrJYiC9pjHgrkymgaxYTGTuveefL/vLCSWo
w/34Rs049ZI5gZgwvPeyBmfYlFMXMgXqnp+jM02o0EX8YBMhO6trfav34tZO3C7MhLCyITkv1PJf
X9qrTrVmHpb1+wZNkoatRcpZ4CCc3Tdd/rFcvQpBg6nNRVmYmVTZlaPFiQpx1qJyBatOYxAixC60
L+KTqKAgYen9W08G20qwovX31fKeiZk4ejdeDRkSfFTR/j3tYeKaoNz1b7gDQhxnHQy9YDzRyEH+
SdrYyLPH9w/j/rZC2lFlY3takCk/Sc92Kg9DZG/3BZ8FNo3AsLmaEXdiPPwEdohg6kSLluroa+uT
deJ+rfZVL75ATK+IrZXf0Pek/ay2Ydg52eX2jMhq+e907yHnSrxLvDgKNVtFQtQe455BhIf0aclD
u74F5WN2+NUodMog3FqLQCAW3WVH3m7+P4pDcMbObZo3h4FFC6XaChL4neLEMlcwU7x2AVMsk4qi
xVVc0s0ylqW4o6jW8lAU9vKM9Mqv50vGjRxLnEKK0xatSeiMATfzJiOxLuLpQDzIrMQrvbC71lpL
HTTutt17Vxd00fZHM1XUGk5g7zfKFld4QAB9EpByAyEwsopi1onH3vwj7a2nlbj5XkT8zUltyI6j
l9Cy6NvgOEbs98+wTbwzNh7zZV01+ww0MbHSc8c4H4YkUWvtfy/ZiDGmILa0Xs1FG0Ly/Mt74tVo
+XjJoU2aN68MJNSHzhokqmG03LjT1rmxhhPCxVTa3U75/Ysxn53Xr96FCslEzQX8G+U0YBnbe2dj
uynZfpf9xGPI1Op0zhvHCb5ln8lLw8aIxZzO/DiMi89/Ah7j1YN2X5BBwUDwhZUjBm37hJ/K1r1O
3g+WmTGwKTQddUN2CtWnDblJdDim0Qluu4quP5h8ZKeLveHpdoiL9cxCi118Ztjzj3LQrsAL8CMx
ox08mK7ABX4Q6Flwe21qDH74tojVGeE4AtN+/L3DsIiTd+m2Ge18gYgRA4ukbWxAK/mfCAnDQxB8
Ej6jrW3HG2VwVhfRW9CJy3GAVzwdbxY8tLwGvQSamAScpkM0uYcNWnfP91twxzeMKRjzJgwzZgVl
kXFlClEHT1MTmK2n8kNZqwx5S8fdq8jmx1j+Lbf++hnhIsW1Pe4GdZGhQBWuRrBJYdwL0ivCCWR8
tRkXLrLvb2GjEcqBFgwIngF3/NfXMhWMobu2T9INmOoxqJgFg3uEaAyiA7mOelhZj53Du5zoTQPA
RXE21sYK7hefHeECv9lCdJyl9BnLeBLQKg/rX0vs4eNERChNFdNW0fHnxaRe1Qohj72Slu93HH+g
GVdw0gw8c9WzzwQHaL+88C74HQk9csDrogMg+yexuKUUGv5L9n42dd2QF70jvqaEcnJEDVW9il3V
xrqCL3YlZx2yTB6/X729vuWjgS/KQGF+KfRwygS28FeAbwl9YVSxVQqmWhLZz6FRhP/cGj7bIaA8
ttcO4cEqnr7wciYK4X+e1hia2rDwLBKJD6rAJ6TWQfoJ/55jvXo7kb07XbWQe/y9ft8g/OAJ59pA
Laht9SBVJEZmGawC7uBUz3HlDgq7xZtVD5krzml7vi3FwVmdGPlpRIN5TDEmrKrtp7wXnFmb6lyZ
iqjT6YhwkaFPLr5pIEB56P2bVAN/1xIQCQwOlr0WeHwx56AFnuepQMq5h7gNPX/vbHYt7TsK/16m
Eo0oAP73WFSvNfm/YjD+K7jYLKZcPCD/0XX6/0pUC9f3NVoqUK3RTIm0VwPGlRK6X5p3lw4jmrL4
oy3l0hKrgUQxfvCYgoGZzXK3WE9i7Iy/hVd8HCuhhoAhkTD15OLN7ii3MFVojwqiHmj+tdfRSkEw
Uc3Gr66SZt/pDRHZ/axGv2Y54Z6Nhf5relihon+vgF/Xg3sHAo0lFm2hZxW7gJtOUQGA8qUaxlKh
nyrlDuUBDv7wqoWpNE/0Lwef+WHQhvRuu+b+jBFTLsvE399sG6m01jrL4VdfGjiQRFosZGr26LpG
wPMW3TLUwPRbjeIHV4WuJAvcJqXwVCkGY51t716UqFkRJIyO3BT419Mm+fOBxcL3DBPkSdeLV6pT
za2+am54qrO+STMhrG9kjC0c60CKqjidUVyK85mPGWGTKxqo+GjhtupB19fHf83okAMoV2/pLWuy
oImDP4lmYRni6SNykQddtETUY1U7ntZJtCMXXWH6WxEP5PoKkkct6d3Z7yfyZOPKgidDD7HSg/sf
CsS/p/hs8+AiBTGpC1EFjN4Hv+xtDMcmZ9l+PQukERrAzuAH4TYObYW2L16cG3QubWBihyj7WUj6
/+Etom5xAY8l5DFNxiT652ykpTJ2GVwvan/Bus4bEV/lNkuuT+bOMtB65g+LUTB/mF7cj1uvgeWY
NTg5qWt2qfHoOco58Tn88wmG4JHtSVdi8OuG1LSMCvp81SCER+gHQaogDYgSnbCzGvmpZqmH8YVa
PSO0Dh1G6BAVfj/PvuS1r9O2y+gZqZkmR0k3uptox3gOXEjoSLwJJsMWY5/FsgBAgi7Q+cnqX4n9
2c6GohEXEl+ZehrifnSa2/HDJ4T0SVoqOJM/6lkgZPffF0lChDpJvmMfUFABhosP4+pwxT+YUWa2
sgy/8Hw3VW1SQWWhZ/Vo48lvCEamW+BsByRQotgngMzWMmNIOiGYtWAxnJTjHqdDF4SlOkBAwoPY
zFGe+0EpSjA1FpgubW59sgiQkGDcTcM1jLqUMyu+Q/uH3aKk1G18FsCvUYsGCtSoeCYInrHH27in
SYDQHNqCjGoe9ZlWwnSSm57mk4xZ+BWSwbtwXWiln3dkYXx0th/SnvnkNmT3b84ZL4FfrEVJLifh
uE9oSWxs7GVxJWh0uHTyhlDQQJ6lT3tPV6vIhzcDuCr/ufMh7GF8v/Gsq1M1Zp+iQeltn5ClAln7
BU3AXjkeZ2fJH3sFTFM7ME0r+owtSWk31Ur6zBozv/QC4Twcxdgird5l0yLilvUklX8DQrPm7JRN
LUUlEQ/UzavR9nO64QJAfI96dgKxr59+Qg2EWaXziGPF0ZuGimm/fFZqqpB/w+lpMD2UCJd+nSMK
w/2rzLPc+hnealvXIZLLypeH+Zg8N2VSprd74Pwo2dOs2cWfiP2uP3O35qFs4aWFLBka3NGMwT3u
+2XHLOMjcAqNBgLVeuhmhVlWX6W9p2AgR8tNExx/AFUW6iiTsTQuYknKH7tFUnaPWwKSMkz51V2H
DGtfhOg+zUn+yc+zpf5OwpsMnw8GuL4AMJLGZyrDdBWXMOyCuc4stlGrTVHA94fFxoz9xYqEbac4
wG+qcdTdKi8Mu+Kisce0KCsuOlyf8x74C3D5YU5caSf0cwVrB9Hvj4jZUMEQdhPecrsRP/VxCZom
ms+e2PBeuX350qG6P+6RWJ2eNLrIG7hzAMzHM4vnTDtJqY5mHBGeU7ux2K1e7Jyp3nGcbo6iSnIx
N7PIEA7VPK1fXdtffYMcUhUALz+PDDfYLdiJcNohAqc7DRj0ODp+lG1yuGhSWwx/jfIbvzBUoNWL
bkEbVoG+pXBsdXYVNVRsDn5jcLYmMzazER6Ohg/ZChaTAgM4KxUQS/tMiD47PIkdR9rDhDGWyeLT
LYvWCRJFrR3gHJG0QaSIm7Bz86wEd1w1QQB4YjQu4ncDXmOyJa0n8Pj+TE16D+LWhLFPuENOfeJ5
RZFl0gwMH5qbxAXj15E32TxECCrKSd6iOu4xeevmSEZKVDzq1kKE4EXYUaCsHRUcNm+beuchjdya
UiHdQhkWN1vMk1ntOjm0UUTypbJ7TnzHk/GPjC8n6tGrnx9mZVx+QakvrcmC2HFiR09nGDVANIBx
s0hOi1cESIDjEXAAcQinDEH89wV3CIVeGohI214MiUsh2PQzIdFmCPpBTX68qo+rx1fNH/CWoszv
LNYxJzOYC6kfGv+ro4aC465fGBbd/4IzFWpKMbSTh+9RAeCXGL7vb0mGomDaGD535p8blPJSHu/B
3E4PA9ztbHOChbQ/r+1LcjQU7omyTMGP85Q0jlwiuEvAPMLpEFBOhPUIPCnQKamVA0gJg2tpuSRo
/YTZ0F0ZxY7zWwsHPbD9hB/Em7Z2WLAxWOERoP1j26XCa2jiwrsVYquGryAW0Z1tOs+ftaT2E8g5
hkbwL6D8MMMFv8khnEeMuxBdBlxf8M76ui0jbJ52HWHC+BZ0Czd3naAbSzjRGLSogI/6MRV8TUZs
7+3WvGomoy2GBW/i1dV5u5/twZNl3/Tfru3WckDV5nPKvvEmJQC2WWBszGD8W7bf6PurkMF4qsCX
+pNdA9O4exOlGUdoDmvRHP6q+OsfxfKjo27ZmhrVQ+B9QhZroB6oT1dYd7RvIcsRovkR2lFYYJNK
he35cXnBClCYA3ajDryalkBvq+Eu4tIAkS0811lJIMX1/7oRnk6ygWKIt8u2LoSR2cShgoMJjNg0
j4DGV2Y36ofvZnwLg5PR7wA8sOQh/ce+q4/CsPgoXx+Pl8iApsig6boErse+QvsnR/04+mI4Dgpo
c5xuNrufnxn3sBZ8QVVNMOSNcgUcPO5DufBHsATjGWZ/Rq2pYqOPfiqeHDlzyxBEkOnQ62o9W21S
gamtHWvcqrGc3lwVw4VB81Rqkx79UosAJRGp3tngQi8/fPH5N06JWO7cb8pEhFElC2YAv3O1GmSi
U/VRNZAXLZAmjrZmOd7Kgj//Banyd3vCNshU2X6aLKzepi14QtiiSMwkVUWJR8eUZ5WT774eHI6o
phoA7pGx8sB6h+sreQGyM3+jxGUQGTG/mQFT4GcG9CQKqmg8vKPERUXWYSQX+f5AeDN/tj4AojqR
1MMYSEcLGPwEtKvcc0krAPiWxw9n0rtVcj3W76gyi43BF793P4Xxl4Kn7OpYE/HMgyfpYAIIpPD9
WwBIH5jSwzodWvlJVaT5O/1mRnOpyINidB4QJeO+D0dcm7I0P8FdoxQxUYNPHRfxLWK4PDf6iH+a
NmY+hRqtel51CKhn8qaN0QnjYrnb8dWTD/H2JFMeBComNDWT2TEe2O0G/jFnr3NqvaGQOUCHbDcw
2Sg0ybtAf8EoNMj4oF/KK/YAEnMvR24JPchvtflhp7BZ2JxM92V24Z4v12R2UpAilvtZH+72Zuau
LOuhTkNFNcbfjuycTFds4WitagR+spsSoljloD2fpjaBk8MfZewUgfxAEscDniLbv8MoJ3hc4j3i
AlBy5OwGepRaw06UkXo242kWaZqZHKBMnA2rCdz7TDT1CLxjGLJglXdC1r7XeI35HJrPa/ei4MLh
d9MS+gs4iIzQtWx8Vq4D/qaWZSWlqBI4KG2Yo6p39rSBkuAFexwJ9EqdQisVy07xHAE6fOXr8fSa
vYpmtXaFM0ms5zmY/vSuGVUtsqJEePL4s9P8s1QKH0GygSgCAbjWx9lNb7X04q2P0n3TYIhVaA9t
XDmKv8pFu6ObwmrZIO4w4h8P5UhAe1QKysfboLvoVzo2CMyUQW78PYViEZTRPoVgQpCbGOc+ZAwz
awySVdQQT9EOQOgmgECaIAcigFcHx56hk4w0qFL9pZQVNAgDnmWGoaSMJ4ZacX+ZQc64UmcLZLCD
L08IF7hA5B9TJmIujhdSsYWj4WvkLDkNGVtc/dpb3AoOQ79zf15PJydXzjvX37dP7kEemSNSROuQ
fEY64jOXwtMJMtQBNagIOexm3iT7kgWwQSSfAufafqUD4DuJZW9n1IfROQ+6PJLgBi1MM1Er+P6G
i/Wr7wl9w13Vi6JcGhlVn5trWrE2rv57QTl3HnMeQwCgDDzDiZaj9GVv7cajy1zg4MciGhIECAAj
gXSwAYWHNAE13OJgcU8YFt4NaYWJhiGaVCTSaVdCjW2c1Bqfq8mMQ69eEsUEyM/8b3S1P9JbTdNo
9Ro9XaHJL7sazlWziN0ahmHYWA8a4ADcsgWkDFp/oYeiWma6dq0LMt1JUY37J7y1L16nvcvM9UJx
VsDU/OnBJQn5RYohAEZLIUNRT14Ay4NRvYsyXl6maoSl0c8l3Ch2Dn08D3Zq/3/ydruuXlnmqPws
Zk2W7o99VIRAoVEqbKA1rYrxsz+yy0Qo9PakuIK56EFoN9G9cBjJzp3tnN5d2CEVIiut3ScwhLBF
9vaWwjh75PtnjnP4rASLhXAOb9VPRMBFBcDIHOxM5JUlJoeMfp2eax/Kj8eWY9HvJuHKH3YfsiVT
pZ3E9NHpDO1BujblaiZ0utLdf8XJe5JO5QDu5tvMoXIup2m7vycUd9sZMhJbWhslGcufuwTxsYvv
aKoRBgh1+C9qfgRcLwy+tkAdC2ENAd+n3U/EIzXOiu1oi+ARzWx3e1cxqrsuJVngFWvmHE/PMBml
qiaj22JqaAVceGxffkBNCedHynoxuxbLHvcdBDhGFSBnk7c3lKk0ZoYi86/o/HIVH9cJOTUDQWtW
mkPCD6sn+flMLMSZgzyKN5pavwJPnAkPnZjCKmNn0LsFYvfnudPqAojG73LUxy8pEvQ0Zd6BHSmc
sqhCNH4kJD7pAZUCCfpits4bRIA7YijTp3Jc6MuJauT0I6tFwylUvObTeCrVi/Iup4rLSpNFMVg1
nDF3q2IahZZKNGeTVSvDAQEgZ7uZAXCf1NGTCZEiOv5EfnZBpwdOYls29gAPGxhF/lEnLcVXH9uh
BOgHEE63iSfmDv9JmsWs+4Npdd02hzs8GWorm0OOQFxjNClSZ1biva+spxxflZI75m73vDpeBcJ3
6f5PLqo+2s+633PokGPxxAKUYrGR6coknt+4BxmvlIrD79CLqi56IkERxHE6yWsefJMLgZEAYtnN
9l2+PUQoJZRaa/ml4zlaK6k5wbixjQzVmdaRj/myuHNhnIkUZJXXfoNE6/xN225B8lGOe+7+sNrr
HxAETaQRIc+6gPdE70hgV14GHg7D76Sgghw2heNYiPiRzgg9XRo21WGVLiu53M60Y35nwLMDVB6p
VdgzOnlPKXydDG1hC5uPTzi+hTEI1EMsaAp8mPfqS7O8ajOP3L7RnPeQh+MTA30VegdNKOMMbf38
H/C4wrLsOFe7dSVQnsVkflY5lVL8DRVcZp5AsedBuenhtSW9vk6RpN4AW/XaBbXWNMqRqoPXgxGE
VbyMQaOoL6sHd5WGZDdGcdD7YqR73+23aWuOKrr6WJCHu3obHppz21hO4KGPS5kKTHNbf0VjF29J
X8WlZGKjz0liN+iA2C7UHRuvlYDIFNYdV6fp6/2GIlW1Dv/B2s1IT+RVXxGvJgbgNBIiCcFzJocl
3uMKDn4MUYnaZQaaNl/DZgxEgyYdOjkepzTRMlps2fm2kOdEvoVPgwTtX5BJPkn25v4yTCHJDnhD
MT3RGL3w3UwMneSLKoTvcwuyeZxtfE6UiULacTzboTQYYqAV1u7BPpL4mZati2EJOtWu7W1U5weq
2G37cTbmY1HYXmBDmD83iuujLOmV28CjoOdKMpxNAwFfXrObAiZNiaJ4UcwYXovRz9rBzawBGDWn
aA4gMKKcoWpnkQWhx3lI7YUAz20IzAWQ2H+nDit/qw7xriuY09sSlFDsj1KKvQcxvM4xOpxwg83b
VVWboCVog0kopMFfVyb9+c5brGiu96PkA5p8Yqnh2YQA3lyMvN+SFAvbZk9NgaI9d8Vsbaiwyxmc
i/rP5kUhyLMO/svgprK2jeyV15opJU+HGciMhryts/PO+DmkvdTdI0rHZgVe3zr4w3Fgsz2H7OcX
1/7msRcvruwOin4s2ACMXhokwcv3YZGj/fRSkxZdQEYOU4QWYXXuEqT/oYFoI+TUXEmfQM4m4D8H
TiVXkHY6LDVbJf1t+PoB+LhxENezqdzoLct1Q7GRPLU6IQ8aB94na6R+yQZPifyPc30D+ntXOfjX
6Y5hEPx05AUcUrjJ4nnmtPI0qZx5JbehZCXG/vGTPyl9V5AdQACgMYBiyZ5Nt+LcEBJOqbqPPl6X
OK7ZSeCi4XaJ1HfBMN9RSUpRbj+BQw2kzHAwSuf4trNQ6HbsjRotVHR2gCXmcMew9GIyjALAPtzF
XDkPDAqD7jjXP9ZN6tk+w6xXREa48uIgNzvIMzHJQF748dF2mRfWKpKgEdgnVupHrMT3HHxSZzdn
S60rnlAM+Yf345EgFXAk107o4OQGxcRQaTfFGK1QXed5JxZVwR1KloStBRoIx8dY2nEFfZIcrqNs
pBoB1uDJG6fMBi3+EgpBSXLSQRR2gZQpZPfB70ZPqa3CdxtP2XOOLtRbfMJ79C9kKjlrpAm9ijk4
LHo/Th9sm1JIWMjuu7oJo2rVLNKkdMZzR3JuoogCQbXnu3l1ObT+wVr+TLFQlQPTYMXLZgRMvApo
vrt1gI2+f3qvOqSLZrRAUZqkqF9qBwgcnlXvyeijtJ9vjnt5YeR1VYFkRyQOffBIelRcY0qFWgjq
BQWFEpY9e+60stFNNFbx83sGACeHtJsjtVE9KRVebJ+mM5564v0XyNU5BqwF0Rg5GjL3wdoMMk2F
grFZHBA3+5puKd2ZcIJxBpqLmfjZ1Q0zVHgr9TJRNc1BP/pqTlMJtNXGb9G5vXNhmXJYpFPkEDgY
n8cQCb2qV9HRdyfIpfOka8ca7Qj2LTyw7SiSiHWsR2Oew/vTU5nd4tnGa2KnsEZMG2tbgvyDzWvj
uOOE5E9N0oeIAfjy/Mck4wlk/Km3MIiOSOdbJhwAnDQMs8YhU7ORC+9zFCW9AU0Ra0TF5yvFO0Q4
60iCfOn1P4AZj3gf3Im2ViqEwvdXQMNUuT8OIUS8rOjJBrUIkJj0K0O71RMQWjAehCGl77v1u1Am
tZV3lcuRwhKa+eCFwIz/ZsFa19agjvX5g4VrCsrY3O42Ld2c9SnqhqKgQ4uKMRplTDID007yoTC2
G3gUF+h4JbRvfGLIBXxGCIKQb/JoovdaRojsjSc+MzFyub5+NJydn6V8DTykjgsyF9RHq4/kbOHl
Nv/Gyfe+CelSZu0Mb6k9UtbPY7LxAVR4ZVaLhzG9SgmekqsReO6nNjf4+l98xYbhOCiIdD73IMLS
VoF8rmTdlWS6TEAVL5I04VMEImCnVeQaFmNVDu6xJ2GNV/JwvKy8D+Q4B+j8hzuL9nuQjs8/Y8kl
raghYVWFa2V3UF2m7pVIjQX+mF3ZvGhIE6dml2O8WuBdawD2wseiLVPqAMK4pUTwkNGEHSUoMwGb
2fX7jNP66a3kQiXNxLwouFRPpi0Vo9L/Av7ua8PUGuCIsYEHD1ebTCat+zMkFakRRJi0JAF+CZy3
oNwiq8nWxdhdGVT0cjNTKdmDBd7D2LaCl3yKpAvvsFuhuF6qASSz81Lwob73jrOryJfPCfdFtxSI
aor+Tpaica9MN7Z/tmvKjnQs9qhthCEoLcSIaXnEvHndFDBYwYwHtxV2QOPTWUO1sDqxuxW79HO+
eSxVaspeVJJAe7AF7BHy3BWeh1TsTqNMs0U1/E2PmQgMOk/GK1mtgLymJknwtKAq4Oy87HDtAzjw
8HRuSFH1PIUm6gx5K7J53kQRH7JUN6k3k1vZOJK+qoiAP7GKWCP05Ns5THb/oxHG2bFpselkpvTU
L8FtHeXJ1wLon+HdPFpATZY0mhuFWlAmyiBy9WOJ0BhuX8n8fo8EkGuZn2dF5EbXjzv/oPB3XBW+
n9HmuUSyNISJFe5eDUCnYQW88+N58d3LvwRT4SX+4QjUgavupLMpiVTHQP7A5we7XShziXm03Owl
9Pz1WnJ0ZdagsJ1Lq+tX0aaMrYce4xYMw/9kHk7HXorHMcDgKz6e8oidfo9wUFsfKs8mHPFVIT/1
w4WndivRx8vdfL9taOKn764/X/jxwzVKDBPeTuuj8Y/fNGA12HlnBgrTTRNDWDYaHbkDsh9OotdS
12aMGpX+/KJ2IZ5Bhw17g8809RugCXA5+7PIxydr2yxRABvfeIw8LA/c081Ia9kvCEtOYnamEKQu
CGvptbehQ/cTKVjnohLvWpgxCoJhXENoJQ9W8cvN6189H0RnX2uflSV66Im77npx0FTCW6dac0ok
fG8suz+5okLkOQ7eZlHLr/RJJwOgmVlo1o+780sW1HrZhk0K8UGm1pkut1cqnwpHR2uV9D7hSZib
n1OUiLWoG47u5Qw6rDtTN50WgZ0l0g/sodLVbqUXSdzjDjJSyjo2J/PXtQG0lHyplEW+WDTn3qfp
/edKf+VQr6PylZFkhCpBuYQE5hM/+Lrwnw7ln0LAkaUrgWlofOhCd0gdESGd9mMpK5LU4OocaTOW
uV6yq6g7idksTzb9jIe4v5B1JNw1GBQSkAaywjzkR9/MmYKsFEf6pbmIBiSWNNWrxdaSRBjIwJBQ
jVIsSm2yNowXh4aXMOLXGzHLyzSUocK8r1ren9E1BRQkXlzJKDoHFueuN5F+BxttlTiA3JzLVmwW
YzhOs2Tajvt59+YyI8itREIGzyP64r5cce4Tm/rlTBpyAppRuTtMPN3mzLEyShbynkmjBAYdBzoc
tXg3lQ/B4RnL3WY8uLo7f91bEBCk4vFcXfJn5a0HB2vGRseUt/yVjctWc7jLeAkQTsZoXq8AjgEy
QIYRn1ILPNp2LELVyxxJPK4y2bBJLH53Vq6ryLmhJIidP9/dmk8csYsvNcCtdaEcjA0H72G0cUH1
/pl0sv+WqelgADK1kSbV8lhrt4PeOBA8/XjQPp3VBKec3op8Upv9GIDDXaZmwzsJQXoZpst+ff6d
Lm2nq9KZpprW0J+7LlG8rH4ozwZqK0ZnJRxuOKqPCHARAKkSkqAnoTSxg6jJLMDrTWI9Kq4fsU5T
HBuOOEdCdJFDyS3ONNAbANZKP6/9cP3GU3YeNtNnmoiM06jjFlZyjWp9D3NlzQxiuiMhQJ9OfEb8
jUdptPsXWg1l6V1hryJ3Vw501VIj60LQ869gLUYCzzgQoa6I5/jaaRGRNEEboYp0rvSQ+X4ltHSB
cFZXYTOzbb2CadEUOiAzXyidvRDyhUshAsUPt//ih/gauJNQEdUq7OQu3Ec6epKq0Hlwx4/VfACd
8O+Oxqgbnm6qr5WfkLHwCbV6HJJDRWcHQZLQUWaBX779J/1uZ/q1iyXUgoFc0e3HHc+BcBD7kv5Q
MMb+h/tZBaPiorObjBFxXq72d5LHzdUx6HO1UtNz6wdbYzLd5EaO8wLHwyaJbAP31BO9DTVXTahw
zbDX8UGycO23MzLO4vlaKIbzNxynuNAvJbvr8DZA2s3lCFSnevjROKSRItkiRrgj7D96c5/+2Li1
xPwkVvTDKDNAHC+2LbYW11Rwk1T9sZnUuJT9eLK+pCdOZ9xVhH4PY7ZA/mDk7yI5tpNVbGtUjgzt
d/1Ibtxjnrz3BASllWSwzFfycZi+Ix7oqsP0HJ+eqbsRauxrehbmXTqkWqO5ZsqQHYPUhfHGVY4v
0+wzNwp98FAvTDvz3Jb7MZwwy5+bHsa1aLLISftsEzEThwR7+et8pQDLhcKjFReiKumDFPJkoixz
APifhvu/uWR73G1zSIYsaq8lcMhBjDrAKKwltWnDwcgLG2ak4kG21RlQVF4Ed+CYHaHt0JcUG5M/
ZYT3DKzrLRcemNQv98orIg0QUpapFZat30IswnPw5J2mt3MayTJxp+i3X0q8AL+T8JkIfmwcsB6a
0lm85C9etDtWw8MyYKRE+ysYjyW5LhNM2UmVNF/YgHhi83QzJtQOe/va/OtzuMcB8bLcly72GFBp
Mmr8OGSVZ7xmQWdhGAFQVL2UbHuiMl7glOxMEweh0nTVl7kMZ6THcAl4dH2V8BGnB6vVRS1X6duG
FX1XbWm9sJ0tkXnt+/2aaFn4l5V7DxvH0Y2R/LBxjHi00EJNTwjwfKKtqVj11oqMajiL7PKnIQQW
ftfZMMedWsea8ItxaqrKRBLZfpLaSUmKbDJV5j2/VoOCglUOwLRoaqvtnhqcVwPULOfYfgSW6bZV
PJzwiIpCYa/tnydMx+mxeNqGbc9gdcSpHHu6cGQcXOJ89+uLh4rbg2clmwVaibttziKRosT46ypR
FMXhYmWt8EJ/XxHGgaBwtpOU/A4aiMLjog8Lla59/lauH6B0FrZqPM+BcZ4fNdoSFwOVYhgZLxzp
l1eyZszqM73vxmC1AGbBlWDIi++tD6/ijlwiSfA/2J8gBoMFFnLswrGyFK/M5zXoctZFDMBqLeff
Kguv2oqiDGPH8Vuuw/85jF6mwJ8hx7d0J/jr059jwdl4o+WnB3ukfzOHA6bXhzWsDhT+Pah7hVam
HT1UEAH2R8onoKcSY/HsDxHEiR1KRpkVzEFKRNuKBMLPAqC2G6J9VYVj4xdrB3gccKo9CqECs3Cl
4lVNSEV3prO9Dr5vnih51QlGKxoTP35GuRSCSG0dmE+dhKmABP1/WDk7ylIDyLoR8fcQsF0fD6Vc
ZtkpoMjvG7efZ4A6EQpCI1oUZDLhHjDqWGe5UfpzUT54IacCnjr945y5a6Azk7A2rh2dqRNu1T9D
cuL2t1ga7cV22TunCWvvI8JR8lM7RX5G1/qhG2DNC1HCgLEOhxpDdg74+MOHtQDNx6CPoySjP+pn
JHwgLuq1U2ADtlfsjRuNuBIb/EN36YH+ogA3xN0hRJE9jopCKg1SvqgzAsAoKUWI1vm7wGIJscTp
EdLrOKi5ieQ3FxePdAmGlH2H43jahXas0Do9taKBL4yDPsKjP8fM4V5o6BLdScxtFRma38lFgTPh
GMUsxed1lg+eayRWF6+EO0BZWzozfGY6PSIkA7dGGzLqO/9BIZk16RsRizWoHO+cQD4565m4mlbb
SCPbVcUMGblIgqiN2rjva5TE9sGYVVwwkknsjo8WHd1khwpRiIHqPBIdWJrRoEmGFSStOaPC6/DX
KK2PqKGy1saZv91ska9h8fpVa+UfzZttURJLwB+B/oMajKB3EoekEWsDkMkzbfsEISUyshgIIFOp
C4oSGsfGOCMhotnS7adOoLMAvmZyVQ4lRqM5tX7AROo18y+KVGJR0eoE+aw82YehLCs4urzjcAYM
vPq7kNbwmYu9XPEgBZkFL8PdhUJV8B+vxTVpeR7pm3BSVBS2AFwFHBLOcmBF0GoN7N8Ub+bkD/Jg
CRViVzQFr5craGnscUMbuVV/MeVCmQsS/02D7dkKu8IkXRDSK6r6h1thDvg8ePgfzUwCKUF2nYpH
3a7uJNEeMbDFwBZwOf1Z9MyS1n7TvIBy0QoSpPrdqwimxYI7kffDXJgtTHmdX+eYP7JrJ4PG37ao
0VT6hgabVzpwPZxy5lYEWixv6f0WM5gWsEvgYzRhZ1goutquzmempL6DmoZpPZYIhmOGEc6d24te
oBwdiklr+anwwjA4AbB/JRTb+N2ZT+GW4MIv2KFn0O10twFsmFrJclkfwrNuZWgZkR8U16zOoxDz
Y+Ff4wcerZfmUr7bEQw9Kn+lSS+C5CbsgVuq+7mkuL5IirqYhCEvzB2/pv/UvvfwB1Own/QyLbag
tYYVMzlEazgnZV1QlEvFJtVoTSW2+dVwWzAJfwrPKAq63YL4dQ0Hrqx2z9LtDUuk+rkomnPPvcU1
6JRJNE12bctSFSru800ic0YKTm4Bb4oZxnoc6/FIgSX4uF+pQ/vBr9aZRX3s3QYIdxDo6NNZz9bI
RCCBI7JVRwcA+XDEy1pZNenJtE5IiBBIBvLQamiLWLp+4Kt7SokKRdCYL0hIwZo6Xs9h80+J/LWS
ymnp1yC+mODuh2g1q2TFtkEctv/LDJdXWrPhKWAZzUcdcQlr8WMXHfR3kgckuK7g0qCu8uoHn5B/
GryE/LORB4GpJDQhiEpABHZLH804X4+/c6cmIBRlnPg9h7sKOEh2O/B38UdWHVSwzWtx/YL5ySFC
kmK5hFJ8/DGhbb4QAo16R8xJw82BeUvzIK/VyNAzbdU/ZjZqFM2ceoyP0H/ZzQ1lsY7PpALGRZWC
ir6DLihQCg8UrGfjT7wKfeErVRbhB+Mbw/3Ngi6C1/uXpf82wk1QqfeMQ61cRTvkFe6+7NLXC9M1
pEhhFwXj8PJYGYgRu1Mt80uFiAkl3T4eGIZFRoQ4hRhXGnssZlPH8NAH42rhlQt0TGWl73ndzMlr
VRPQf5LtA3Bpy3EekN4xJf9TwoJ/+qapUcd0cUy0qtyufLn4XCXx/esLtr0/cLwvwKIsyJZDMQF+
rFHTeJABIs1iie8qFVR104tRvyDYWqi8szVnbl171Q977sbEPh6Sz2PTYu4ioGLegiMz0XsKZbg9
hHknLhs+k7aZa1NGObX3aZhHfYBoWx9z1T9eAaRp5oDDSrNzZ77IswZMmg1uC/+Q9+cG7QSRYvGK
GuIFLlWpwdSzBNkQVW95hOMYzKULj7olLJbaABHmkykXt9/BqhRnScM9pK6BCHO6+KlQT64h8IJf
UXOseiUJlxgk8MhRJfdCqV6uGrWS6JuELEakGBPKDsYbzBO/IX3adAa6veW16gKVaGKXo/Ya6Il6
VbR9d7rySH3mQwC2h40NUE3cqPFsFT2lR7+sXXzKo35Eu27wUUKR+QMJKxO27hzPErFSy06vl3tk
kuIPsPfYFlbEuhIGVwftnILL5rb7cDAXIUlnXBhO4oe703yb/jVlI5fOdYRCN1PWup85Jtj5BPsD
75dGXzNNlnDGuHEzir9VRXWacrB2avy8kNgyxeNbSqlqLws2D3/QeF1MqFOpLLsS+lyiZOiDg1yF
/uO5qRww8ezykilym1wcd//8DhHWquAx1wMOrUiVgS+XBbXDwbiugyDPhsGuV19sBeFOk2wRH+RW
/yPVwLzfxj3ufo+yDhd+XIY5i8Q5ue6rlBRz6bzPQg4zhFTzDC23+JiYODViyuHEgBg3P2fORSPf
7JcDmoSBBLEcpxoVsjKiBcOZgCappdL67b1e7EmzTVe5fic1maQCE2NWaDiW0CLjCCkcXwCTTIVm
DdGIxe2rSqzp7m/SFmqNAQ492+mRx95cGtRRyvPW73VWsPVYHQa2PG9zc5u8hm9Pqx4gGHT397pl
Cf0z3dPVfZ7FxevMxfyY6bqDScdOXKW1hkOAim/Z3DakVfsUj/p5nM9EbYm9anWWgZQ6lw25rNXg
u6HPi+8Zipi/TzS3bcC/ukXZrY/kySr8UXz1lnfKPtN1SFy+/LvwMqBFgWbC+ShVPBWEUZH2UIYz
fgPNN1PWd9AYudErYKQ2pfOKeAR1a67s5PLH+TAouk2BCw2H5Khg7MUjMbvzFmibVzYTbjIEF9bJ
SPr3g/TVTtOGslrp0gGR7NEdV61gJ3aA5pNUa/Xqg13PRGiNM7v5StM+HQchj5hdxXIqUL46sIt1
mT/GEahIhD5jNDVXlx1ZbOQy+R/N7MQWZc5iLgjlfkMC+JpotI5THGaRVtJLQ6r4vnjyurMSu/YK
4p7wjMkK1R85nJ6mFz6gQpjM243vRWfZHAqUfuj+Ps/hPMVsW8IbCm5QYAfo7Eits0A+/ISYW6iz
L0qn+SOVmT+h2/mUD1Txsfbxs9KOWpL4PG7I8JyhUVSYbzeCTWMTtkylArlOlCtpRo9xWtjMKGA+
xuzjVaBu67i759l2AX2VV5Gwe2B70ZmH16P/K54wP3KgLNfXrUQY5YAhN4tvJtZUTiCuMmoNECDe
ml2Aj0KUawz1Mm3IuPp5zgg0DN2h1JOXhLVFZDJyHwwc12mJHR43Au1hwYgj0I82RqqQoMmF153h
dCCCW530nlWaJv4JJB42B+JgCygjkoWdBdd2fZucSA9CtYe/hxPJfxrrH273xmVniP31TBs1G2Ta
Vie+Io4tDwuc3k9Jq3eOEErZ/i8HuNjzXHcg83FM3EWE0S6oIgunP0mFE0vYgxCxVepCheezA7eh
Y5Kg+gp6O62Zb1KDi4ViDrU1YGo/4g+J3YoWxp0x0LlDANPtjv6i3ROlxaj3z3/VYcKHt5auF5wM
yFskBoafVTjtCoDHgE5XpAZKfuJfcxVgo06UQHykIqp3WoJ4LSohOyurIbvNA2Fji3a1E2I47WMa
NQ80rkE9JZ8skQmqrEqcvIdfGba0tcQ49nsulhBmiflXyAvKm4z2eW7Y/Qa3+oPq+6w1RTrHiO3A
2VYyQtxnU9uGeDfAV7o/R7Vg05xREMr8dX1WHxSk5j8dDzbb3QCvr0ifVs8cvjF70mRxJQNAa4eX
XzHhLARLquuC/5Ew5AYdPkk8Yz3r4wvkAGZLya4/Tw+wAf2bPfExJEwKguWzMTWO0QC6LhIvjkN0
yQtYojmXlRb6ayY69mcXhSnQOCtFB2uiQm/rAtOC8x+WJeUVCbnNqFwDEmBbNXWiygW8jljFBNku
9OXY7U8n24japrYS7c49Vw12CKg8bYXLDYrqkRAK/p7yZhigpnXkIgynNtyi6ACaQ/9ELi5bnF2e
XtQPPlxskTGZK5zcOSo/kYMmWif+9udpqkp04jW3BiP6bTUe0/phz4sDS2VhNjnSBhy1Fyvpeaai
gXtggp5ZlmFJ80pQx/1HQWSBrYPE4dMM5CGF9pIIPBpnHXZ46qF+VsnHUOaaFcPkhzpbioiDiXF+
5+MRTPAubfZyH1gwuyDswsW+Ha6eyQY++7srwamCEcIMyoIC32rNSh2Z2fNRak7lMXBH0kD6lcNc
Jhapl9k2k9aQo4T1Rt9O8ncI6xb2ixiyVtgTF9ek0MklxbRXz+SndAeMuV9HPim3A9jYHlg5SxVw
rqi+MFdRYuabRg5ozX+GzOcuwRgKPsOOlyC2l1j06dfEzHfqlpejgiY8JssKuY+MtVFvD6V8Waeu
t2zW1z/fFQ+LY7KeSvrgMON51t04G2hpjFD/RNvYZUfw3SU6ZEmqmLx5SrRSL0PjdEPA94PfYHup
v1B+k0B+DA2H/Z4EL//anYGzEsGTjaeXqRaUTTB3UiTXS9yLDo16YVcRYIxXhf+Fi3gtdXAfR5vA
JFbHJ8mVF+n6qPA0lEJS7KXubb3J00Rf27b1ys5EUO8eA+59aP5BeYCCCspz0Wrsn4FIIwLIaz7O
WYgDJyCIhCMjQZOFmUkBSEonF8EU0bVUu6GnvC7EpkDmjn3R8+bK5B1lAgr5pZWXddY/kwwky7sG
cuGmP5g1HDvaYnbRyUWRodUJPoWEoVGVBz6lHtRpNdKRMRgdKS80xoJ8+xPNTFaFRvWXZEHisN8/
GIAgvmAwBUA3dYAUiUPFQhYDbQibySju0b9oFp71uctV5uYsb8eMa/VROHLc+87YtDHnsJSAe5KP
MSX9d6vQGoJSW5ljBNZMhw704xLYA7/BDd9xW21QY0RM3Bt5qWtX3ts/5GotTuDryrI9rUynwOX9
mI6y7JpMc+NYtXuF+oG5NU6obJlnQeBuKWinNrxgRxDeZyDUQCptZkmM2KJhgD4LL4A0sAE5pnSw
xlq4MCstVgkUB4n0/me7LXQuXys5+di8GrqriBwiulluGpl84qz+yG5pDkRUH0D/6mOPzC4DY7Ju
44C+OlA+LXBImQvfPy2L4ZSmuu3uyqHV57EyOWf611tw12HOlxqTF0mRlTPReymwAb5xIRZRNDXU
DTYR74/qTOjK1gqq7tfLbVxncHxJY4z273pkVAwK4Vu/poJ4DSG5hcnWIPqSK3KSCbow+70DinBn
4d+XIwFfoeqLQPOBH+wj37AG9SGlXX5V5xFVnDkV15a5g7UqrGV4jxoBtkfBZsDXAYC5vInoDZek
dh4P4/izVAoYD3tn1v/dC826YPS+r/Ox54wLq5Xsruc7xXo3uCzCE3J/tjHbohRYor/olTBhZbBz
dj1IoYFLpXkImE6XmkOJlYB0K64ystkDcszM3qSbLAH9vTu/FwFVmM6Zaq+aPJ+5tS+phLh9Spx6
m9Sqb0LB8SExKF2czMHFyHXxPRukVjKrxvn/7E95J9i8kgeCBR6DKJBckHqruQyh2LTImwfJ4pbM
cesPscsVl7+KWEhwkZk2PgPGcXW/s7ZS7Wsg3dBoKV5cnHF63oMPZ7yhBZAOCLAJnXTp1xhtgz2P
dGadokaGUNlgr0s16KcOIwlfHw/VMsVBYvbs74i5AByYdgml+UtTR4Izy3KfyEf9iVgEXMMNrdL8
Ndd7R8hFr0DzFHOuIL2h5/KDyqtZThHB2nYGkqCYs2AVq2Fw8U6OTudkKMwFirozZCY55uce+4O3
oOReHm5KnOFOH3Y5Zexl/HA/c2wk2bvx30yPlCwh1O3kK5/DUyln/rrMD095+XZ34630VLR15VWI
7c5bVlJrMuSVDuRc/vAL0yN7eJPjXLHlSwGlITKm5iDOBUfUjfDshGWZJLPkywW253GZKhsp3EL9
FDsv7NEsIDrBQjPgIQSCbkJOLGmmodzrB5/DW+ASIU8xGgdzYXeAciq4iipRT2PakVoVFruPP2gE
Sf6z4pWKAB3ukd/PTFSGWCN5HdOlOlwKs9T/uLmssY5E0Tu3Z/3OgMysqaO61OSgK3FUxkbSUTsB
k6YVXB3MUGbvFtZ5eX6Ssqi3IXRxyxWIIDYQgQMCa15kob2cG5Nb6vg2ryeJwOtAa4mcQ9r7QKX8
Qg5/eO9K93YRAlHgEIuPOguFx8vGcVU0gPUUHQnGMus6t/i9Mipb8eNJkB3AkD53aKw/iL5b3E4g
ul/eRtm3OK2aqBZ8XTJ/6sOXS/pwAV9G9ZoJx2FeLg9SiaE4HSQnBgNkt53jGF3AMlah4Vo5v4rA
OBtc0XFIsQe2aaiysyZsY/DG7DHy+govQCtdJK8S1uCyKxIuLVxQepc7653ULqfU/DG6M/EssIMj
h0zUU6bOZe+BJkL1K64ewq79O0u6u85Ra3k8PkCMlDF7NXWYAgPCo02WlpiyAjiAoIXLlXEUvA3n
cPRFEvh88jBD5v2YgkAc0SYvQpZN+3Hm3B/UP16pymgFpHRoVA1RGxM1SsTZpDXEr6EWNEN3JIp3
3RV2WEzpWrS2GVuXea+RhVkdCpgvYpjcjW5pJDAxi8Wi1WnukxMngIxFl/wD2GsPbQ3C3i7Z/8ue
Dg3TNAFNVo82xJnTtkrJLIMzsO9bo+cfSK0yBl7cnnwMlIEKuVjiV12n6r0cFB3aADVbv9z4H8dH
XpB5cJ07y5+NCQsB6xCAcQEe8a0fwU2W05q1ybrVPKW0Lol9ViDPJGzRcHN105d9dGp4xxLW5Ei+
aEMyNrtwAF/Ka1XfL/GzEHSZRL39CcOmJxdrfagECP3YqmMUDxdoIkF1gdcFz89EJb+vqSSViLI6
xez5IHHToVpOPmW8NsxGOXejW450UZeL1s3YdS7Qors8v5jDV+MsyTCkJUZEgwD0uCnJxSFq2cHt
9fcGJKgdWyJUATkWzGydIET4ZCUTcf9Qpc1d+qreEuokl4U3vXjAXBdgtik5oJmlEauZqbhOBeRe
tsqRPGTkRXjMH1CImE7VoPolElnVO21HzgOiKwoOlhvsyL5RxahGOu/SbSUHbncMUn9d/4PTs9lA
rN0MxKWX9V1GKzdZ1N9hhmqfUgr12ykFf4UbLbI99sP4E7C87Q4qsdkQ+HFASAjRPTuULhMlNP7U
GA4viJXr/fEX787wdUrNCHg9QFtIRmYAfkcOAt6o+NWi0qbSRf0W/w1mMEvw5lMNrIWnqLIAeSAc
K4RQfugE9Bz5cB36OGEGFiJm8ud7aYocLWBhFrJpubsIE1Z7YK3Smu23wNeKnVNzKFOOhFvpSb3f
ItjvLkWderMQt7RJ5sPZEFLq/t86kwCGlOlTE7hmYDSUdoRpHszjYf2lTc2MpsSKq+TzVCMr08eQ
ZS3hv7rFms2wpvY32QUDcvqpgtAh7Y5hcKHTlSOKDRSkJkhChWLcyDwpKKgDa+jNIaX1tLhz9Q4A
UO/IibTSDfA2jGCb/Ot7Lqlehsajst+6+cjvKrqjGVx5Pwmt0L+MybRWpl0o9Tvfk79PKS0hSspO
mOlj2Mrnd9HYImAwa7EOfvWOYr1McYT8cENiQ3fE3MAqDb0PEfeR7PPxAqB/ADfqrF4HLV972txV
nsN5+DbWu8y7bBkRSs6yCOzlcgcla7QNI0B/if15KaM63ogbBuGqU+yllb/ssL/aTJfmAakLpUEi
91ZfgOEYU8Rl0gGYK9mIxRc2Ha77D5nda8ucn9YIVj38BDFQAYB4r2D7FI80qN9EhP2U0W1IJHme
vLWve31r9JtMMhjBuXESQwvnpYpttvEEyMgrmaBgkVjyuhkqkHfcdGNRNDtFF1ARsPGKZYcxLv5O
nLPg6r8wOdf2xolrVVyBi/k/b81UBd477Sh5oxOKU/YG6ViHNuRtTSPKqAmvESLPrp/Gzt06AUpZ
1GiVI95Djw7tLa3mCaBALpfU5c1JqCZ//BERbluIrzcA58WwqTrX1b6vTujFQ9vYa+dtkUcl18OX
4y0AZKjgRWdjkFAEDqfADyNwnfH1XCT0hMoyVUaTo6/DU4KKNhWWJBvHOH5pVUXhRtOnn+lAquyr
X2wOKw4wxfUQ44/vlJPpTbgdNADqNwmBhlfjvMQztzuXHIjz6SOGCblxz8ANnRHpIIcJWpgxuFrO
cHWPql6IrZ31q0fv2tOwL3oICn4KFOvPy6MYPqH/O1BRf7XmxAj7bSuJeLo80/zMMPqTqBX96D6K
/Osm2v19JOi1oX1+9pNPHrUL8ckUFaBHyz8+b0eIbk4hyDNo48WCNDfi4hCCa4la391lLLv2njaj
PqdjfyMq6C8jr6gzYtCdAcOx/0H8z1pQM3w8NhziB+JFXYGDzbz+B9BVtcId2HmaycoTl3AL+bbB
B2GCotGWaGbq/m+DPUspD7p/EE76yoMuWr8OaRYJM50IToQ3A5ESawnYKWF7+F3AC4ouH8saDHEA
hqL4YkdMpL6koaRCyZPMK88IuD+cYD1r0dM272813lqf1TESSEasoL3fzp35NCX9B3QFXKGniAcF
3EcsR+rIRpu04avtwyzusUmwyMzPGyMJxn5U85ElbIIMReDPmBbR+7sW/qcJVSye/GH9S56PeldP
bYBXDahoJ0aKZKRsT2fOt2DPl98clGRnnUZONqZwCvETWpVSY5gFItVLXF8er7T1Qx5bYvO6jads
YXGL1OBa4WRlYdfJs0GkqqhdqvcbSBPnoKyu5/NVOjg4IKrKo6VFf83il55NABKWYHqdtYhQDd7n
hZsigdhuxyPN/a+zyNjg1Hocl86qMuL+iCAjFCv9zLxjTOA/ecrPoBGw+t+SFPceOyQxSIsLq0uq
7kc5L+EZbiWbwDChQsqZGoBRxjhavGqcTBsbpjO0HjN4CBO4/FYk6//brrypHlZbrkSC0wIMRYhz
GEyJ1+xOnWsp+ful9ju6G+ltFy38Zz52rPeVby998l2dKnfzUZtB0UjqR0O9+xH4m2Rh5P38i0FZ
ji/V+30NAIbjgSfvIDCGSc1B1XWlfHQwRQn9DvrZT0AGBdK19U2+YFaf5USBHt8Zn4rchUHeD9vr
XMvksAJ06OeuPVDQtbBQKuh/WNntj5JHGpzdYAsEh/OmqX25XEh20fYEWFcdMAvVdJXffruLkUwa
WHsFJpt2vF6Lwkr7M37mA/r6pu0IVfH56grCJsEblu4HVkNIxFYK2RUtUEZRJiNfJyROeY9GA80H
u0ZspAlhFECzIzIQjrK9O14m0HVzlFHt+opMRST4XBh/TadKR9M5xz3+7c08QJP7hG2csrkSnayI
S3nuZ1S7dK+cD3rX9//0TSHgbUfw/0/AmON/9E5+YGIcpkrnQ6zkiXm768qf7XWW0F4e0R6rAtcD
mXCZ4aSx7i+JoIIw4DuMZN4vPnmUXK9UQifmta73ScKGVymu59JlLNOsVBHQlPQPxUR6C4oyewel
GdH9vhzU74NLLIYex1L9DfTBEji7oflfO+dp9galIfArzdn9KyAjNOMWEoO42YprH6KuU37cjF6U
dJQCFf4kBdbWtt81E2sK4Lrdp8aJWNutaxTduFmf7+zjbsNqmt0XWMB7GkyoI3pgab/K8YyS+vNt
FYC/L448AyQ/cBrnINfgBxYkZDdcoAecDMbW5z24OCNRtjYdcyPnX5pZLDiBA47E11Apda5w2EEb
Owf27OeNV4ciWAHMX7QaoyQRn6KhWwB+yZxZ43hQboOmwMVL6nHAFooW1o8RjUUr4c0szHCFIdtj
Ned29JyC3EPAJBZKB16tThjVM/vVHArpVHnuJp00RcveZ64FT20nnYxqnQyi9uuSP6bAMXpMwchC
iWYJlOCLenJab8lcXtBJeSkcsGaH0fZ2tXG+ImuuAzeXwMwqOqf8LERc+FkWqM4fGRhKOyuhvZSi
ZUedrg3860tQE6lLXxLGUc2xGV5Kf9tjNXt0xZTpXemjfo/BhkC/y3eXNB3DMbKspf4/tmS60aua
9kP3Hn2V+OiMqaEVTyg0zp8db3yhxQMgk4Bw87xbmkPIccqdNMsNerh9FBzjzBEbu1EjIx/qw/eZ
643F9yCN+xF8ck0KkdFeZW2R3+Ng2YDCXFEeCxSiC9zd1TD92LY+DijmSC50AN6lGRrj5C6M+ek5
Zr4QQyh2r7INy0tJ6zhC5nCv4xiwMlEgARnbKs63x+3SE48UTdfjxcVaS+OBUjIfN6UfD2xbIGoK
r8kdMgywHVeCIZBZJ6mZrt1ZpT5dpOGe0KS+NiLLoqiUuyITf5/9wcyRMyCeip5NXnADma4R4c7E
QUxr+pnBTHtb+agAR638I2kOhjAyp7/6PuFhcd+QPQkbaCb19Em4Ipl8YkaGPoqexKLuM9yFSaie
Zj69bN3Mb1rW+3wGpXuqe1xPMbeyINVpk2BtAeLr6IvV8cBHyLZUbVLVMg671SoScn34PWkSMT5E
bnfsnj4SBAEWsQW/m2dLaxFMK3qpZwAn1FsdSMqFp5jqCz7vAKMQXAvRXNv+9m9xVLsMrUQdxOiB
9hVJxr5XWNPH7Ey/5CBfLBrZPi40NHS5ZOlupZTyxULH+i+Dr/d9z3PThdNth8s8A8Hpj8ApgR5V
1MEYa0O511/V5DqGmQ53bstrtT5Tcbpe7NtdDmd33HjBd5yNe87CmBj26BI/4RMUzl3p8j02Gf1w
dFZYePqxg0o8804Enixio+eap/1HzjbDenEwxprnDR3dDYeOJKJ9vaYy1bIro0jTrQUxuUbQ95/e
YRDNYnL+vzzlnXcWkL4lyGM4W6WH8pBdYFXrXCEirPfsxUgpx0JjDphC5PbqvLpJW+DNR6nzgI61
DV/XFG7YrqjPjyFyeTAciwWLPM9XumaSoKy4sv2/+Qj0pJYmSXtRhymiqnWVPGqu/1urTjhPig+G
MRH9ZJEc2GG+gwXYVz8hDg2dTMfJtU/NOlGw17FyTJeegePnPJVz1KnL2fImP4hlfMv5GPR5q9gX
elaKz4DKW2J72j4KZWkd2spDy9nZjrI29YxMPYBMajQ1sHooNcsnbQHn5QAiKhK77JLuK23oZlLl
wmMmMqrYcq3UjDZkniZ5XDMKcRo+4D76qoacd6bcm6q7Ev63mvccsboT7Yr3dgdTwcMluoa1ZSwA
HHoSIfELEyg1Q59txMCpQcH0jYkYniXkoMkwddMYX9D2DjNPrsS6vv/XKFDpOVqp1SERVDq6F9X/
voGDRzin+ONpaD6izTHXZabaGZHIjMK5O5P8afpUUWF/MJbmAwxIRibXk3ytprZXI+cZ4ngoYnT5
FrHeiXeuSGI8xy2CMwWYxuBqfac8MW7FdDOhFw9PrgHCgZqfbjzgiQfjCsn4GUVgFCvcoC5PPVUM
MlO/aOcGVvFvks8mXWAd+gvtst4cRsFhf2lOY2f4Q7gNMe0kADRSYZbLoMeXzfIzK2l81HFcf/0l
UHihagRJSairdgZKNoRoNIVUIcvEYB4fjIBp9iAYpSKPm1W7kFkpAFjj77jt16jz+70uP+lyDXB5
WLaaJQiD5xia6aPEGNUSjg3f9R4OYoCQozwDZtylqFFVabZOCV4cWEzzYcn7c+cZmJULwqmboxob
ylRAE8TqmqPdlHegW7EOtO0HHGIsEikgj/Ea4woEzxtffhL4OWC2cAkyZJQA3LbfFpP14ucqw05+
Y9A+9A0pqy4SGfAkX1AEk1nNSpWLvZUYylFJv0RpFZ9ZawL2U1XIyJP/gCJIm5fSImc7hFsDqxGM
3m54PHA9RqhPEM5DiQpXi5rZoeQEvJLsiZzSG4Ugrru4GfbxtvN+CEW4WcjulBa0OUaYb6UQgQPf
ge6B8EQuNEEF02O5sZCgteUfkEi1P5rIzV3Rk68VtyDRj2bvqA28C2fXJdvLuXSfANJwPwOuZ/Lu
g8eXf4AnXZycI6Yd/78JLq/CoQ/NFEqHF2GqsKjoQNB35dVtRKsMmDTEbd7wHZ3vVWnfe0ml6nLr
dwv08UEAnw3ydXUy1i0cY/FtoKkiIOxl+uc+eeRFu/rC4cbj0YEQP3q1LR8AL4uwV8ygXXVeku1q
k6Yq9Atb1ZaTvkTEtsq3lO/aK9CuYSu7NclaBfC27l1z+rGJCv6CqsC+hoosTp0uR+6dnpE1bhjo
GwUTUq3qaqO/hMLU2xcfzL2sn2jD1Cp5McRG7haytZUwQXsWQoeJ/1LgpYFsvk8i5INMtKCIsE1N
5Jtp7fHRs0s7AbuWHKtcY8jF7yTZs08Chs/Z1EeaUo7keqTOHJEFPEb/4c3qR377UMEBhOC9T/LU
4Y2CTA+99xlrhZ77Z4uGTjbt9nxdb9dG3elATra0QKGE5FeXhooA+lFTUY9Ct7Z2nczFf7IpiU8W
VVFYa/3Rtn9Gm1aQZzJJgap/F3Kck95IR/oWYkixprbcIg6IxIGESWNIDVRLSWVAM1LDTPZx/kCX
yLsoIRoEkqyAAKgdAtfRte0US2A38orDy5vgBSAoMgBzU6aX3nDfB9B8VWDVZH91XleTeZBpIzGy
fljz8L54TxlplHtNAxF6T3rFO5II3pzu4G0HDd/hS7usvULgkDkD8/hw3Qfg/yJss5bXSjHTD8+4
JiPX8B7+7F+ugchLdMYAqzaM//hBcd3HkymhbFPiXEsbuWLW2R53Mlh+tVwh0zMRGalNsoWNSdnl
y8D7ujzFfZynKgQqTIIL7xy5OIPuhV0S0oy+gSbgpQIDlInw6bEEKS4mjOJlYgPWKBfEyDgOBmtb
lYZ+Xx5FkdFcgjHdfeYP0NmHh4gIcr+FDxkBz8CfbKze2bKTXMsiYMnq9wkHooZZvwvMNnt6cPcP
VR5WI5VedaA2INmUQ2HJDUoASwsGF5OHPQ03Mr0Rw3puDUIy+flbJzH0AohN1h7Z4uBhOHNsxQMU
sN7zFl2ug75ltYllaIUoMcmwb4YnqQ9tApA3JK3TYG2OVTk4z/Xd/LS39B3/OI0rNz44TMI01m8R
JiLTmhLN9wofI0bhttupbBJCiR9Cf8kciuiJwI9uBLC/lUP483GM38dlBzi5P7TJDQ9DrU0SmDvd
CwblZEa8xn75nw/j+amQxZolDh4hCF49kD0mFX+Nz/3f9gccwd4b5YhEB1NylKw1wjH5y4CVN0uV
8mXwM8kCF01fpogRZkKv9+ClJl4RSXUIC7Xo8wNrjfjcitC8flnBEQURcbJJqATUoWmptJ3Z8p7t
9fOIIFvWX1vK/MLC7yteDkrPLtskfRiX1vEfmRwdsUp55mjj646guGr7SNIcTfUwl9UZYZ75ENTh
SUuB5F7KpBnqvN8CPU+abr5Vbuzlrz5DBUEEcfmoG3BypyziWMOOBoWLpXxGh82DUkW33dJVtb91
mpD6A4tVB9T3Jsd8412PNnjMQNepGbfsag1s0lwdTl8oU1PavUiejId5RZI9kUOgysvIoYsQ4WMw
IDGmORZA1MLsfTvKpWcnKiAjaQ41yPzFn0TWNQm/Mola1e69NIG7QnzAFkdmFKaGcGuReJcz85kj
phNFM3GP56XRrxpNu+9EktnSrndGVLXUUwPq9/2e2QZZv1ZOt1XvlKN528gY/Itz+q0C7K1qWHSy
KCFpF8ci8FFUGz439uNVbnqWPrtymy39xYry5+zhTn8lMC3/m1IpTb7dlna1BK7j4t/jo7yIjUxh
mexyBfdS87dAFeWZr/3+0+FmHMfMBpAqgHsNkqLkzB7NfqMes37x7p/yTS8J5i+MvIqe4NmQqjsU
MVx89eOk0rKHMNy0J0CtbrL/r/w/Q7Xq691+uz6EiO7HusA0oG7FzV8CZyQnD85x4M9kTpOgMNwr
qhUyXdx5QvZMQABJxBgBCgGoU6sCA8lAd2I4wsXyVKKg3ddrpj1kDl2zwyKfCzt7jow+k3+TNG9z
VWRxu7VU3BuUxfw1myQdkb4La5O8irWTUDTidvVR+QzqjeZUEwzKNcFlnoSMdpicGWFfCorL1HlL
Gl6NG3apWgf34LFnChUy/nJhh+fJmV0f8I7X5nXcJ4SKst+/OvtxWq9cEFP41JBtltK3UIexhjbE
sE9jNbjNiNz1jyvTf6nhJSGtDbrnq4ljG4r0YiCX3VPv3MJQIUx5SqdtpGLvzFZTxLNAWuoMf1Bg
Hv8+TDoEI7WHOQawsLgo7DqJYLtl2BKJoRWJZwnOTst0WTTIL5TLIB1EguDs7zwt9CIL6nh3sj/Y
KrTTrw0XJ6lthXTg/qA0VxJcUffjo6WIK+dt9Z5DXJmWxrDSNyjp/PU/yJSSoiwmzJ/hsKeO4GtY
p2GbGf/E73+fmLPhqciyLq1JApuKJ858f/HwVQ6Xhndy7cBa86PEJctmuT9QaDt/u/Nr6ovdW3pz
MtGa80sldLUNYkRnB1kNMk4rFuFI79BIEKVLOYcpP3e0vDFbB74tOhmZxivsESCGt5APDcqE+9su
e1vRPP2Af1eESEvEXugsAei1ZUMx1Ifq5zp2ADXML0AAnQsezzOJ1TJuNWCChf0eva5M+4hxaBVe
KvvEgbgeXWa+Acz+cBcw5Ic+qAL6hWfAZgr+QLlPNcaHdtfAT8IpJTHoHKU8dkyvJIEG6RFw8wCX
JAX6hNGw5OW2adcWQ9/zMdDe08znjoXG6HfzJPLUFxHbazT81ubB1VVf+wdbtOKL5s5Ragi5ej4Q
x6M19tcagbebbK0pcSICGx4PnCmZBuWtoMeCQVIZ8ZCljMws4f9c0yEfGD7RK3o1QUtfnW8330AD
aRMAUPdhyTzf+FCcW3BrE3g5uIHL1gpYzScNGehhUgRO36HVZUuc3iErRbrQXd0KNQ5FjVGtxJC0
yeOjNhvISjp0yXEryorx4dGQE3+sOHoEiZ5zIcO0O+1PRdWxE/QM8vovfbC7fDvPbFCkfO95jJPy
CzYf/6fSfTO9avxTraPE1+esxsMXVNeNK2hJ0qqrOxp2sw+ixsLKfYmaZDxa2b0XvEBE3azP2hWW
VdgARd7MEUurHdTD9+sTEzpq9iNbbrNNNCGe1HcAjTk6ifybLV5B/ZiEF3miHjdzA4H0QgeVPh1M
jWWWdq6niKm8axzk2EzKAu+GlVV76DaHaJJc58zvM1yHAzPq0i5k7vHWKdPFxKUg56ROJOTssgke
qugPXvu+mVb/5cm9ax5YJ7bwVNXq2bKvnagsSGLUqcF0KWDdIaMxaFIpHlUNeARJXTPztELUJWuV
UphwIEE6k83jOhBd4G0zCgWLyrCAa4tDV6JxWG8ozHy3AfqbIiauXqYy2mMUBUzN6kr6f5Yr3S/p
yeI4Q2SNmAQxb0f2HJKl8wQ1MY15fesIsVzalgINLQ9r3JcbhtjFSUf6gSCBkVyszFsqNZSxzjmT
PBuPFGulo4jJNIxquoh2SdcKZdyla0PoOIf2IVPetZCDROaoG/BCkFlbYYQtaT0OBog2xkLh/tZn
qmjywATvLL9zEfDkPw/fzEpmwHxE9otucM0O1BcQRN/T32XGD0h+Cp2T9sMsDSY4S3QCFEqM3TnV
yUH8M5sNmJs39+SEQgFTRcTV9fk9LusACHRDvXLYHLuivcf4AeQ/JE4LPRUJPkctLSdKZuSLkFVm
vBqItC5z29eqph0pIaJOLxz0C3Tc/MeVZxx3B0WNJuPnKl0WGrX3pc+AQcpm+Gd3Ehu6JDZxKTpo
bb0rYGG+MG4/0VQIpAtHUf5KBQ/SaZFtxK/cJeBDdTKnLoT+ea0DFlZ22p5NOzTcDHA0loD1y/pL
YvxkiW3lcAObCQ55IbXWWULAnYT+YTcucc/afg3Mki3x1QTQ4nUaH/GWVZSvpP8h10zRJdK+jwUX
MW73oQknl+CXF5Id3GZk75isPcsrDBTiGdTp42zKEYzx+LrTp8ifXs+YelNZNclVZsh6+lnqZLQi
lqpRcz01YCHrDE7za6gxFSAeFikjY+vbLt8i8WZ0BFSJRXGoPeb4pFLKxBtQ+v8R2cay8szmnA1l
g7bJow8csByYl6QGBHVOPu4PXLGEB9IQwQYlbuf+RSc3BEtwRCdFiaVbJpR36oK2DO+V/hSHvESU
zgPDZ6iNhWGdq4BsOB7jeZsWgZM4CqUF/jUSJanxhMl7HJ9HwvcDzkTyL+BjcFpGHoA3PsDs44sB
+wn8449BojsNLwUyt+Kj6vbszDoZJtYJaMuTeOvP+0cIdgF+/l/F+sxHHgt/GO2E3n4Fcj0vsx+W
YWMI6vHfep/WtY6PTJC+Nxm59ADdMlctoOLosyZlBOlBHZxHj2zLirJ4m0TZWaUkbzkvXLn9yilP
AJngmWdqTTg/lHLm1w5b64nFVHYqSSGAF4lldrzzqs/cdMmAfw28udJpfuDw84rGjUqlqy+TiNA1
mbHAT1IYIUhzba3F+F5NJmosYmxgEmPBptGRFujzza/HW8bbGbOjkya2MBLPW0VyEXGKuGfiXOpI
/p7r5rnYD2IoASlCvcOD7PWtMc07hBlsHhEJX5d81nGIaDaas/lvMybs0LeIzonNmb7xvc1pf6qa
L9PyknRAe/eUcsaysXeCV7+xuALntMamgHPRAKqfzKkMTrTLPgdc9S/ui8h/Hx3f45U64DGJtNrO
lv4Ex0OhjFRJNKjPM7L9mxYcnXOziQOIoaCcGK22Q1WbJ5gZmv5gio2XpJFiNNHyaXYDlM/i7GgP
4WnqUWa5IzHICa1x1jzxZgGcdjPbElsi7BS+H9fuSg6PzFTtghEltRI9BuNUYUywtWEdzIH4Sy/x
82FeVUZCl93OLgXxiRaKyFr5rWtnKuVYiAUJCe603Ra1k6fYnYJDtt8z7OsIYXy318CBuus8dxgY
oOnRasTvPwoK7hkROm62SLLhJjDG1HK+RHYQHrVpgQRioezQXQYP+ocIwKuR8RT9pO20G4hWeOCK
08jpygnQ64uqO2S/YMX6MgUvkNg/a+0+laDXwun37Hm9E1TUy5TS1hLhjalifEssMObhRZ79Tr7V
Cs9fAPHicuce89sGZrOQCAH/PLAo7dyXimbj6WmHSiQr/n/oDPNmz1REzlOO5oEOxcQcpH3/Qi7G
/bj36/YVtgg1ugJTBcWwA1v/UUThKselQt+x1PorG8HZytQOGsVVJ2V6UXB/u0nV0r2qDJIFEcg6
g/oXqYwIPrKegwVVZpKOhbpXjA4sncpi0EA4qeRMYDuCJsddOPeCCAxkL39tLtEHS/fmjriRNUCt
avivCZG7/fhZmspSHG3fL9cP7lyQ7xh8NI8sZOYQjxDVUPpwKg/zBXVRpk3tsGmHkVust0Z23nMI
/3XiPo14XiUNWdWl/vSeLZaCrUtTNLn/Gse0GwAgxLvMqsrWOJaQU/EJnNL36RE96/KddmCvbyV2
tVcxVfawPqappdkUXqnbW/0E0P/Nrmd/PEHZ6yna6JqlyZbfeuhfXyDvzDBwSHzrcgYWjiZmVYo9
Raqu1wPcS8QwrQsurLDR/oogqYTQXpxBonU22MilxoAVNdQUd3zV+4jZmJLPE68ndTD+xJzgOY4e
HECaEWAYSGSIcVQ3CXiC9pUWtDSfMv5uwy8rBTlhpkQG0SvP8UQ8V6IKf0j2D0wRnqnfUsuK5540
3oIpVQrWEDg4Rx4lnFnIbZjjfgxinAasjRU0zBl0fNy6kW0Csp4g91GtZBeeqG8uJ/+9T+DDIRoZ
7YqsIQErJ7yg+Cm8F7A96QOounROJAL6e7oSOr2rR7xQ71UKhJyJhxCqWI7f84Aa8uih2FGKLSrC
fgCJB0oCvNE6Ptu+Emftw/NlkCg/Nn5VbjQkabm0qJseo3IT5cZddyvfnmcma4/EuBf0m3pLrnlz
Z0KjZ5G3EQ5AaWlyorsbTK5egyoiiufwJyn/3w2qKVb0ZoRFy1n2Og1Mz7IFIcPLbY8zn7QcwLzP
+yz0H5qJZB2Z7eVzoZbh0Cub3HySRczEXueZEqYDNL+g8yA3UYyxuOqAdiJ6NQCm7kPaJNBUWAgA
gQaXs9OohjNkTORlevDmXgz0iFtU/W/78G82rN9F31iTTRIUgDkXfug4CNCTBxlUcH/cm3dIGwi7
Fg/Son7BEX+DQPzBmuedECjXvkLiiMHmjo+6vKV9ZoezEQ3xm0BAR8SVci76cjBn5CATYN0NFu4v
WWh11ctc10UDam9XnmHGpFTOaFC/k2AHTMtv6yFv7+hbFUwXr+hqKlyU/iZcdlJZeSGY4AZKpo9r
QubrZz1kunskwhjZb0uXY2bz13mCzld/YE2GRdYjgW7rAogsJOkA2tvWec5nMpaQSUnD1PzTCa68
1em8ZFgOqW68ROyMjkHl+XlAWySmfl5WbWZ7GX1s/cJbYkcaB4JzjQjbvKzREENuDcPbrWYs32Cx
dq9tV8gdLDsZ6g904zKRi93d66D6Qd7uL7ucPPEfXLxzNregIu/SXSABVGyt5YN/7lhmxCHCDHJ3
LLlKKfUwQjx1GUbzFcxe2POka0dYqrLsB1pP6NLK+4cLzEVkDnPs8qZ4AURt1QsWFoSOEce6xOet
QkiSU49kexT/2OYNTW1xH/IE9aKySLdD4mV9lKfwgYZi0HwwZnkSxjgk7hDKLSzr0KQ0dm26/ItV
bBcTmi1aKqoGxGRC37Qy68GfKSL82BTDEGO4NQ0yOTi6GqcpRrHGiyQWHakloD/poG39H5JBj35r
pNTerQ5na9yPJQxMQZSxvem/1xXX7iLJ0csqZKfSi16LQyMFadIF+WxY+oLI1Wqr+8bbVUWL8vHg
WFlEnZ8BruVLOMc/Pji9otZIi+i4iI+462M6L0VR71maDyscL0Zt1VPZm1Cpn8sspvM+X4yw6FxY
lPmsKGJgyXpeimSqeFrDIwBFlGa6/WCzCFJp5apIXHy03p5wHzA669jV98rSsUf6hLfSs1uRCmuI
F/AdDFih67n7P/D5Vnlk8dFYQ2OfAx8cFoUjymlQAKc19L3kLaRXJXc2LBQYZe3rwWM1DSiKaWtp
hJR8SnM8em7hhOI4MMn+8X9sukmFOgqQJPEpxisW0aNNmfTLEf5IucS7rZ1CF9ftZlicki3fnFGK
dTDzOLBD9fmGW54OtVCvsFVTZIf8aSw+++29yNsO4VnEM23PfNRex7d9J82hvfLS6T8rkzDkAdk+
11yqq2JcA4yFbnwndnXJDynkQYcXH0cHUNHyml1NyxUMIIH730qbbaOwOshHP0Id/uniULgaWykP
96QxQjnbvRR+p8p1MrPrWhz0yvcgikFCVR5c8IXKgrNw/81xstFKEjWblv366/pDdObOcxFil6AP
U8gOFQBAM8m7OxKYW7JR1f+ipy9Juo2EanCHr0JAHkVrzyybOQlZem7syj6cD8S4Ysf/OSYbhXCc
ICD7JOiom3Yo09nVHUF0BCm7UV4WyRJaGHbnLX0kliZWPHh2rOa/vvAIew8hfRugFGcANMoUrS07
Y1ZVJZ3AGuq0Hys+sggFiexs9huuLV0qXsW0szG1R1YEIdFK6yl/f+xs+QtwFZtIeScvQL8QrH0q
x7dSBljjq3SjZXKFzSwZGwBKW1LcpRren92AdNj/XaCb94Z/2jDyjTsgUFkPE1WytbmYBAOgMZQ/
AZ/nFcMO1seiodOqrU6Pfe15BEyd074MJDDJssGeLsvvISUSzAI76obRAWbD0fWeaN+XbWwIFoRD
QFK7/awZzU/cXD7/vgClNzDaHs9Dthtc0i6edK/wa0yBY7W9sKb4WeNj52Od+WrRMUhTbn84vyyH
LVcMoPWxIy7pIRf/lhvgy9IyZZdzxGpssv1uCjg1giHdaGWkc9Fxe5XluERzhXf/AnGE52w2EaXm
PHIU4CHf7fCd+MyclWbpxIafC7uo2evMqWZBdK30hIe3p8YKSxEcJ5T9fTkqy7pmF4PIB9dciIMK
XzzcN1+gRbgHkB/rlCx2uwS1eCdlLbn9XrriSylRxkAfwwQ5kddpNEk5FQuSK3lDIbOpfde65ahE
6mOHrPLf16p9mRt0TI+JjLcWbohgyiYfr5+Xg1SYrzccWprh6dM1DeBGcKebnc57Nj93uhGQc10h
SjLnPujXQmQu6+9MT5XaN/+ydlKKnZblI5y3hET3MHePWioEVOO3RHwBWaVcO0cxwG6zfJBA48nu
10Nj1mxvw1dyjQxWYdXJG1kUJDQ+xi+wPrxQFOypN0bT+R4CBGrTfzVGujdvyWw+3GU0PXYIoGsi
RF1NO/kFwqdGMuETk8qRSfeYUPmNbz4chDGb+hu9O90WgBDUvscsWAHrwrECzbNQQ6bHmrjQMo9w
peY+eX4o/K5bVSshhY0jyLvADRdMMy18+KHPVGaF7Gu2HE26n+c+UAfstvYcU6KDCklCFqQJnW3+
CmxJN/Pu2G/0Or3Uxi8NUVvR4fdN8ks883aymuFJRlrjbQXNx9OpICRKlC1qQu46a1lC/kIANLTU
IhAK9ungWVdo6pq+cKFY5nqGYoBFV638FOIOUfDFaDSfBK5D5pwILDLWt98Pea4nlaD8k8ZxnTmL
YkA36NCCf1XG0QGbomRcNgH+/BWxU21PO25eGddv/9TvDBUAQjqvhc+gSNZHawxw4sg100CAzNPq
iUQwhHIwks+wmVHbZdDcVNWY+mPXUPxVH+dIYkl1Khg6+P1qYgxRPvD+BFRRAKR+FpLe9GluRAd3
pNcctq65NjyQqqL61u1DVaBfd58HnK23H9oZ8sQJwR6lzuXVkM+QN77hwNZsKfF5IJiJne+eigE5
NptQ66mngaxbkq7VkF1A3PuzCZQSjy1a6vfXnzzPncnAIXKkQtur9M8TQ7fdOrL5Ro9yCPk0ZSM5
U9fmGZ/OaYPwO775lFSl0YznJn/QB2i8mC6p3j5x22bP8DA1b8UmWKZQdzno2Z9vLpdsjDZzWVuI
bcaKZyTUf6Z4wI3cbjuuXf93lIz9nMWY5ONU7QLUzdls1WxJmTc8Y6LCdYB2QBZ/t6YeKERgdaIx
Zaa2osnlqiL05M94DgT7trfAiYiVeBvv0nruqHE3LwDpyAR/bw8WtTklHBceHlgTwKUjXt4Y8eV6
kwflZmuU2JdRtuD6TAfjf9WDUpn4hQna0kYcQm9XiuQq2bipXuy/7x+O/JwMWzgFNUVfS15js8Ja
A4cRNb7QXTfN8YV6NkoEfLTerNZj0vN/BmQW5o0SZYs9ULcy+G5E5J9Zv/2POqOAbagws3r5tKjq
+Ci1TZ/1jktGsdiubvycmDKbaic2YWoIdycq6+l3WY+AjB0Fd03+6XPEvcv0X+AN1RaMnXoyoNQH
1dOaWRFDo0iESUpropVx/6lQHhiFvu6DT50G2RFmLMXsizMt2ySCaTUY/rYlWM2KtVsOfx2Lt2bt
RoGcoiFKOPsqS5PvCiCg+EZWEz9zaVnQCjKO7KreQ8RfEM0EwGlcZcQx5j0vWB2srmY94miolp9S
OWumdH5w8GEleO4SaqwOgWnlY7bOT4kbOg9D3xp/Rxt7RedEru2QjO/81qKOqnW7RdArwseCmE8b
SQ+w2gKLDhllnYVZamcadL45QoSMCbEzGZUmHbK6U7WLBCB1rP64HClEbp/7xgHYNoycq7N0v5n0
FnLQqaGK39+6ACR8mjkzev4mEaI+/mCXg8PQglX6mqpK4ba1g3LUJKUqm1mqFO5gOz7I5tu++Y0h
gFtLnJrJs26za8gz28k7aLywUru5K7z+TqD5gKDMO5JQQMtg19hRvIY/gMrNrtp9KDjkvVPhJYWv
6R3eLzxzFL6c8Zgb5oYxN9zuMXIZcTS4NF7vWnboTpSsyaG4cdgpwqptRewYUF3/o0cRalQc4q29
6cUm+poonzN9wwaZYR7WA+OPXA4YztYYl0SkwzZnBGP/f6/7sWZ+81gAOQh2+r/xEpfLLThfFXE3
jYL3YSFqPDhJX9ckmCWr8IylpANqRDqznrsKvVaeH2tAoeETjBkA+rN5X/nksoVadRzVxidOJinx
xrHMB8B4FH7sss9rzHs2eKKdQWFO0flZyQuVYcYq4btjYYckIWMjcV/2QQvaHq3zt+PMeYRD0Y51
qRr6kwWRwV0cP8c4ks+kADOB/Ez+ckp/wKfwdmXt+DY4751fJWDeTYnT8BiZ6dy9wdAIwu1YSZa7
3OAnYVrR+8/KyDCF6XMW3nW2/b5g4wEGzpHG0lg1Q8vuBNp/xx6OBF50xPBMR373BjN+bCCIrwEe
3tmLeXLRaamO5QZJMw1sUe8AeQHSV0mMFq0szTpR4WjtNnCjkrK/YAcBbhGAZ0KEfnJ1qQ1UiNAt
LW/wCKeZP+2iGDlEgA9MfSaAaPchQrvRRFDlchkm7vhJT6oUi5Jyvgq61t4A8aIQ4jzIse78nUe+
efisxXfy79BMAn9bA1rh4N/v8QwaVD1ODALQlBke0xMZetOFYJ07jO2CewNUEHwW/pzj7H92sgxJ
jGLMBjsmK2AsoqPcVimxKUI+nZxM60UO22qVFnUj4aSRGnvMUtGWaOuCAq7IOGF250kjvs1hZGdW
NB+LcdxWhTwDzVNqfR9zrEChs4+og5F2LM/JNuunS/ILQwdFA4f8be5SM08CnIeTwHIWfC9O7v4G
lNpuivpXcchn7GkKEpjlwAuEjiIlhaxYPE7Y4vxIpc1uFqW0eL7ZP9IKRm3hPv7mPirgTKLRj1yw
8/rdOcRIONcmwwFNHz+J+tqC3EoW4znCwbNPAycVv8aewBICQP59gmTiWHXLQTR4xMYCr+B6d71E
m2lseT4YBn9DUviemWlxcx1z7pJQiWr99eMbFnYc0LeSfm/M2aPeJ/ojL3ziBrT97sgrxdJbvwzp
O08asndXdoCVDxyJtGjvT719yebxq4cgZt71f+rB4M7jN5AzGEYhqcIyhnlye9cVpD3sgnYCf7Vw
LQW99LQqBIBrbeYS1WX/ATdzq7jlvssPemJoO4ggj+IatyIHbcqgrxXIcHKWCo1wekpvcYJv0oXT
wJtQrkiZl99TOq+28XvEW16TuumU8SATEIVZ7D3Q72H785YtOctVzxcQc5bs+0oaxIKFoe22PqUf
34x+ru0JqPTwGbnwOVzkMce0+92CCHcsZ0x9GA/p5pTq84pEs/jGoXRL6Pl6wXhW1sSoWS1v/NXU
bmXf0n0qBR+ScfKnc62xIOG2O3I7CViqUhaRHqntsxK3d7p65NCU95U1M9u+ctrC/NrtGi7JAeHz
cs+hpqL62i2o7GE/d2I3oX5VR56pluYqfbRXW/1WoO0fM8y0ALrh+Zo2l2g3vTiJaZ36CqxDS4+2
U7mdDjcZc0hSM5xBUKHuqb/w2OT8A+PyA8LGigZSQ5vctWSsx2wa6VvLW4GteWNpN+14iRZWLVlh
i/B6aCttzIzDAJGqkT7SMmOPd854G+3Aj0v6M9wmEjPOSo/+Br4AMWkWQljYYfd82x5FKZ3Kaw4g
Oi8hK03DZZyGIQqtSLP/rMr8iS4LlzxUC3lrKTUnihrc6vQCPpErBRqMdX6yeZrH+4hTA6D5vvEH
YEOhCcNuNDrIlvCQLQPnSuw/hiasxXwIasHiIRGwA6rYLm9+usaXEl7ciwSrINtrKOzDvNFZZU19
xUG3QKKi8Dej0HOpxtZiTO1ee7BYRnTQHm1x0Q+VKCo6U+9A6nDKDSC6jAFVtEP8mhJVhIfVCcSD
XZESvzh8BOuSqv9ty3Poux2ChLRVC9yaQKSmNEPkhsRKrXpOY1kYj7puTd2EDw0gJZF3/WBY3vA4
707nU1NL2m6wK5pjSvrmf+OfTSIrSE20rVdEU8ImNACbtRyNH+xlNgPNBUenbWGDKrvu0ZUy6PZI
qKNFnsX6KinMxkXzr6F0L4m7jXI/UIhs7didrto0Bt7tAt63F/MVtcKVqx6NokcGTc9pyPlOdLSv
QNDbvOuhy/7jAMFCJ7684Xi6ifI2dSr3kXDV0ujOdqbODxobonXLxrmVmtGJczOJKp+aIqTqm5In
OJ2pND0pnx9kY6/MZIDcPvSwI+OXCYu+e9OoCny9NUVRev93+BgrDjTE0GK5xaaKiFnkd+e/VvMS
h3nWkcXtwSARVW9oj22VZPpc0m7FXtvM7UfaV5LX1hty9zf6fZlJxzWZD+PJbcO0Kut+PgIjnq9+
zBsBfAJvEQ4Kc8mYh1qXp+n592D51kRiC9p6ynXJg+Tabb9PVaAS6FGFQlqg2QqxSFSQhcTD3yDC
Osk/1kUZAeWei/RaBrrCxuMBEv8PP0OgUKv+mgAbe73qVEMrQj1klNUqUpafDXXYdrwt/ndcD6RG
Mdrb3Ycggk+lCqRsm/1y7/AnH65TA45fetkeqxtKfp0RbsdHThsxESzjrvAfYQ24mxdo09ThL6DM
31VwybIR/hu83YrEon2tkvR00K+Ws5C0h20eYNQK7jG6NrGgsQYH0g6wbhxehdw1OybH+R44JR3B
0tZa28u8ftp4V8DATsWCcstEobc9eDr5E8zDU1mNhGWjduwjTus0lh+jo9QxjEeDUfmZV64xCKpa
NZEjpEeYPU72bmHJT8Wi16p3QXFSS5KesfKbQIq7FBP2RmG/1ojINJN3+wfGXA0Xzp/zXg4EOBot
VSmoFIB3i0BwF1Hc9QpUPD3Vk2Zmyw6hnKhbwD+5ngoxz8tMJX95f5gBEg9FtiL2FWyTFJufJ+Jl
/ygxlVvb/denwT90AdLn/q7JTd1boCgovBUu7/ZIepFKwa/FhtA9sIX51obF3xamF9v/s1Y35zUn
gxAsh/QzdKQiPdQLaZ5ydrRuhWvf0rD0tOLG6AZ9fE2UDi3ulvE6ZXOS7O6OGNb+Cp1PurFKKxcD
Nwpm3ae8MFXuheZfB/zrCF7ZbYkp9ZaFtHN6u0WSe3SC+SQ7T0aBG2/W8hsLe4wCYcaNdJKpf9Uq
5W325psR7rBS53uy7ofeUfU1jKLhFK0uTdGGJ89qvJch2W1c8gRdS/pTK8vIsnvvPpJ1LU3sybSF
1QpMHh9HkfloP5mTdNgMLS/ZnC3gkvZMwiIYZsG+AKVDyeFw9V1p8VBNo4v4fLt4sZ/Op2KFZE+x
U//muHO3GodYzIiaKsPiI0qXWK7c42pJmnrNuhkBQFzenlYHjps6kpK7hESLtaqfBSoIlze1aXXJ
oLHbJsaPJ6mdUSVEMbvprfE2b4MdJHUYIIQqXU6/l4IucyBf9S1JKJfHcVGlaW8Any2ZwvoH6mg6
SDlMFtk4p8i3aMkbSAlSHkLkUNWwccufi0Tf7SFWrbP+BnNyPa/ZtQuRaAy+/kSuUiSqev4lkhZS
uXLgA/3MJeeyFZI4E3XFo0c1h0D96okNORdb7c/n0mrnMsAbVbHEIBzhC2DAyWnXCiA54u/iluRx
Yj/vWm7dnz21ZzhjBSJ24eT0G40SduY31Y6j0EQ975ij6Bn8ZECNI10NsW+I9hzq2GNgvI2auAkZ
BvD2gMxRDfESp+30BhTg1If+5lCfXrECqufP1UkCxRWt058Xo1iQPFspcy9TR9I4gtx1JWEwhV8e
gwdLprdGMMafAzi1QzcarJu7fciZmrdRMGKf1NeFptLyPNo6pjHLPLnWKRL7MEzn9qY2swrmVGdh
u2kBFsgjuZ+seRu93ZHwWTeqrtiqglvW4Zj+qZeqK9wn3cFPL7riJMd0tXupCBPqgivb8wX3NdT/
QmMmaZ57sXtZSY42tWPM++6fWuLFYzzXa4HZ66QBqJ+GfPjZL0W2NDRWuSjvDaUDYjOyzeN5iNvt
j80+r66TL3VIDyYUwbShEt1nFQLQcM74vL8w3fUfAdhSEIUmNUc+Q9bskzPQG4yQj90CTuu8z2/B
iUieQVkZCPX4qVlS2NhBWbdiSH30XynYD0SuRCQW0l4MiZv43eCJ3/ltYeSfD8+F0LDVNUTMJ8az
7JsnwKvsdx9tDIUb+APu1VjrYkwNBT+/n7hiFT7/7ZM0fylhJ/hkMqbmHlzC+yrQhL85NDCzOAF+
ZNPOwyMpD7M9ju99YNmCEC4txOFZU7yJlQeAYkDkBMeor7u+lIJIjZHwdAAt/fjVaK7iIJSNmBC7
aMH7bPBlvVLIYaaOWnD50e3XDAsfxvRQ9V2wea4/+YJ+S4QYQzLp0OaBfsAZLs1SAf5CPpz6sjcM
1NxLUuNb4n0ppRsztgTLaVU+TXzEA6T6Uv63qu5PKBrVgpwb8IftplVkLviAxM7yaSsxO3lqExDk
1DBIY9aLnx/5CSGn/z6iRfgW96hS/KySy0q1qO98HOhPaRVDjNtNvhp39wBHwT2ru+bGTD6fxrC4
+nPNfCmGH4ibULZZ6yli/PdxLNw+46B3zHZHa4zgNmHS7KXFi5ykZEFY/+sKon7J4xpdeR9VXA1o
PSaXs3DsXfCqOxGpWsuKy19VDpvrMs52FTGZ4sKxbx8g83BhoU3K3TB6bNXWOsfUveU0Cyv2vtiX
EMHRqR2BAzCOmDqDEyF+e7NWs9Ofofhscmvwg+LND9m3NwZVUjJQM3+gcisisLn9bm64Uk+JXHSt
24XU+8h+PMu1xxCzKwWb+7p8VI8Ct7CvULgcQQJhg0v9mVwk3q7DDu4MeNDgS8xBOEspwOh+d7f4
Gfebm3PlOHAVwr3MuKKSWkRemhgVko8xVPZsM0FC63N4ve8umb3SZVdwUyAHlLu12/zLQVUm11z1
xf9ZNSDfV6H8jGmQVGu5GD9bY5TS5UFm0DrKWD+FFljBK8Ru4P0R6fxG5R7HUFd8ScVQFabORQJH
dMWg/H3h/8eLZnN3hdVgJbh6OKZaQJNZQih35CkIxCz97fCtad+eEm8IpDTFzfLaMoo1kbc0DaN7
aMZKqzFgXUtmEpmp1DOq0+QLsXV1Tzt/v8A78k6eNxJ/BVqujvRMkm4ilRGvqvzHOOae8rz7GFnj
65HCw7Y1jKVOHjocmZfopRajcFSrmjhK7dr2XrXEim7/gL7XYepMUzamJ0AZhaad0OEH52isWxpL
9gRoyU67AkHYzaA8SoAhpPs++aJdojJD49jq5MsyJDuhCe5QvRpnpCvROtnoBaN16YIzzZlDcmD6
Hiz9rMOmnO2e8npHvB3RJIr9oKKDAmpba2Iqv0DILV9d7t9/ROhFPWGD6vRyaQwhNVLDwjl3WVCF
wfADkykFQmx/Klavu9RH0ZS6E512KalXxGTS7CqwyJksLb6J/vJwfSLQmzJNMwSrrqW0r9LFh0Fh
rzO47AWLbS5Zz5A/WZWwD17PA6d2MIkUNwwtx0vGCv7FalFQExQtC9TtKonoATeh7aiw6EsKx1Zh
Wcajnq0Tl/cAyugW5Bt2uEXI4stVe0+tj64yBadgmXj6ponQbkI0k1lDLU+pYPWVjDl0kFY2J/dH
BLXcjmkQnZ9Ue9J0QiJHaz8D3yhhtibf7Oq2q6rOGqgqmGT7ILAS3Nd9XeD6HxadNdDPybeQeKVY
6fPBdxxr9E2CwZA6h3Ilgx2KJ64pA43F8JIV6xGyI+D+l0NNUKpFn/m07B1aFSNbmKad5aQghAi0
y+ASJ8wV3uEugjPqE0D5yfgfwSxbCAuPp/GbjnP2PfiaCAMH/iU8I+/HeY+jTAHm1fWTb68vhZHZ
TpEiQDTflwVIzXu1MRa1/590GrFhtqVdys5bjez/IRmXX/oEL9P+rPy4Pr84nWDlfMtgHrqBMPiS
0yblEj2X2jaLyQ1jol9jin72RycYB00Sm8N2CDsgd83FGpR7uSo6HCFF0rZc62VqXjp/DQY6trdB
a5OBHUvirtZ7MDEzRnhajZHramR/DoyZHeR4J6rbN9/5gJrqHttXQMpvZOjJswAzKr9y+aUm+LFA
crAolp12qNCz2z3fiIjdgal6HIMbSK7XpyBGGIUdByLodPdrRjwLCXMTZaFj0ZQe4WTvF6pmH3hK
DVgAXub2pSrdm6al0RP98Rpt8UW/i3/hF0JTUntHcOM6EG3ocr2XuZO0OsYKlOrYJVvARRzqSOGN
MIMJzHEzdxZszT4vHRQkB99b7vJSLpgR/OcVpm9axvG9I9L/QjluK6Ym2Qd59nPIInHFMy+SHMaV
yFlxhQMXz7FB+okzVRDTmTGOtyueWu7lOPxQx4YfDIrMmeSgZfKIP3wRv9SndcONFcvGUGnV8BOt
+C+LZT/j5YzZLVgeMnNx3EwW+/liYuVJbMXDI17WDtP6+CoB9JRryInhR2v3Bz0CjgqZlygaK7uI
b8nubI/AWIzt1ifg+gwMZvs+13qI5uyBEAgDSZ4Lo6YrFGSj99H5DiO/BDk0ZAQe+Rjj+YyZIn3l
QI5YvkkiRgOShVuvZ3mFso4NPP9F5nooI/yWY1aHmVYJyrNYXO9K7N+xzixIRGARUw0nxMGtc72A
IN5yAssWlg6FGnoe1W6dCffuiSoS1QC4CsH6z8WaCoauovK5XcIVYBK2V/8E7Nt0+vKa9pHalFWO
GsBCNssEsA0IqnPaXfoc/sGVL5M/46Y+yKxm9pUaJ3AyZQ4NDSMYJoNz7uxkWazB7ocbIIWsUmAQ
/PHtMrVBtsmoPI0S4ZgOnd2MGN/ROIrHrLvipp4gE0EaTyJ5mXawDiuhzT8xJgGSsh76y1wWlgaR
Hv+3cf7lOfVnOd24Z8tKpS4zwrbaryF8SQ+Hf/mbiUmGpMXGq2Mj3eOljcm+0OzMzE6ViSDeguSj
wPVP1LmOfbRWCaY+AXrgi017uKRxuaCWg9Js9HiL2bsTVL1UfAI7e6Ms879ogV2EQfIK2koGVzRg
skjr7fYxiy5Wiw9AgIaEiFXi6prQfEc5okNSK2Ogsxztz9hLFfUodFsmlsMT3nvrWM9Bml7a1mzF
FDXc5QhlKuq9fu8ZViMq/CEvsalCPkHyPQVnGlzYYRl1jASJc+heE526bvYn9CbCBV+ajaANex3I
sUQeEF//aNyAVKb7qsTksNeqz8U5gh5rXeGgBgHQHetdfvS43fWALCfvdbMX7f5Jcw0ECuln8MEm
zXGgEy3W3fL8jAvutLayYp09iwlo/Fg0nsyKvW/GZiWFG+EFAlwsBlXSXJnkA86efOuTEH2ZiEEs
hvSnPnTwRzzE7SMY6acSZOub7dB4F586FUiwgfrDZVVSOjAOBZz3fnKs5ppjcbuk7GQJ/tUkgvhb
w2iY0my8Iwp/VOTHuJce/84ylVgw+99qybG/PZXodtz3QeuJzUV3d/Pvjn+hysHVqwjw2K9hkpOQ
ZTsIBJMHXPLWfFbEcz9LFHd6If0tEkrhpSzqNTHzLPyJbS3AQUkL/5Fn1m20jOoB1CBn5c1MaDZ0
NNnVR+owm6lON2hqMFF0tJMkyiubIS8vaZvPxmkhW0B2510ewCYo/tAsXJDUCKe+oscLAKDV8ymF
twjOgSBFyOUhHh4abr7ILkyx9gSoxn6DzPcf3+Z09wFl+oXJKHAW0tqqOdOPJgp+XmS09talKWGk
DLTpnfGcS+a8JkLhXwhG5Ynz9CCWfTmMLKwiYwiCSV9ztBCkiSXCtOdGm9qV7e/CClBSLJ/D9sPQ
9DwuoodhsVd+H+shJ1WyNJYvgM0736oPz7G5IJKxyyNVDaVJIiuPJ9Wjo6dh2SfXUeBovtuNLQm4
N0KVc2G/f9TLGRY6GYRp1klpfsFEZYBIMPfpfd7OGPs9+t61Ty+9BLaNRdxUmlpEjFY/9nbEJ2/L
pilgu/ZdRjgTA+9yLPzhQmI9l4Pk6t8fiyI2c7aHzlvMy6s6G59jvA6zeXqV5zuoR8au5BQzV4pS
XckiwkArhuwzClCYOuzKm3hNRyWqCzCaPwwJl2qORzrb78EvGLf3glaVcffG84gXvgW3PuZRKLz/
cwgDTz6+6fpjK7ahNdBL/Tv61zp1Tvc3ME2Md6pcDL7+GHlUEjy9e3UaEpSH2+d1E7ai7COP2iY5
ea9RTIKFd82B6epPlF8kTS8sC4xc9tX8nNhIMVA5wZh983DRTt2xK7VuuBjCmodvTM9+f08IV8q2
XniKf4JzIZU2IWqowbdKpnDwKzu3ScQmXWLbt+5Ak8CCoTdi8NjxKaLdddn5YAhDxSgOXyXLaUUG
4BSjWSL5ujBr4d6a2qHg+x11X22k8zbTNGbWkEErPKQnLo7y/d8ICmT7GJ26OwmDRdvZj9lKPYuO
YwcSUl9fs86HCOPbS3gltlYDt/1qs/xEMtPMKOE6anyZYjyBOhYMNnT1njB6dwUcvOBxZr78k2qf
HU0T9XQhxJBdzHy2IFYOj8l0rYfSTpJtIu9kwtXP9Ue9KGn7UICE36dIwg9Ka9s95+m6tvs3mmNv
pSYvEL14m1iIahGXzYgEqbQrwdAGY9kT30UxuaV91lSo4b90fRtOXW6UpV/qrKHauM//ZHh41S+b
Tz3DPIsj+w9VnVMy33Ll2I3TvaebIgW0qQjuNoSvFS7SuFVSSplXj69M+hDttgMHpLNIUIJlYrn/
Q91cBYHf5JVWq2rnxig8UZ0KMFvQFKCabOYb7TD1XzfEryIZ8FwBOrmaNzOHtHjsga4k+jqBGi/L
F6DTFCI13LgAsxuc0wgB0m836Z0IX+9YVy4ZJspesHtU1n1AeMp/GuokdMb/sRwlVJ2jH9WxCbaT
/Ou9cgiUhesoSkGzSsPMdorgLyUOoKSgjLY5UwC6e7+Spjp7b7D4HwYNkd9lJ87xoZdbGqwNekik
N8QVXju4IbGhJWuEGpyzTUs7vopqqZuDiSag8UoBd0iyxGDqLTKpU2iXIqOfK1ZKLq64fDeCcQUA
3760sCgOynSIVqp/HtXy1hNHXoVkBBqOLzScYaQTJABnhJxvrLxLs1/eunlqC5AYQ+T0aBcTKBYi
R0O+6y+/pW0h4CVhW/GxQsitkbBXnfE0M/9G4uYBnxcKxv0WgPNdWZhmxNShqJRhYpOH61YBgTeS
6Yz5x3Dte9tX7H9kXyweSIW6pooADf5aBQgD686o7nvEjsh0PC1dbOK3EzhztIA9LsL1AiEHmEDQ
ETRAavn561fbhp3ypLToItCgfv47/78FEJT9xwbSt3IOBIDRW5LHK/r2h1GpaW3+kKUThxD28Nmc
qgVj8JvUM+PUM42czaHNf8DQSoC3ZVPuUqh57saBs2e/XMOo5rhvMs+zTGssL9qwPl4caSZPcW3j
BwdDobalLit1WvE8+tHj+h20S3LALi8nOZMJFLZAEC648Ds6mtf5CyOzczc69ZWlajdVvJyTFSju
QKF+6bI6uUxHsO3+Z//4g3w+OODze/sM2Jkq5ZdPN459YCfsdeK9qXb284fmy6K07Iolq99B8EVn
nR/y91AeYRTNbVEpbNXPlns2D+6ZRmuz6Wgzqf0OZ0GwD3JFAIG+DLAENDJgzzotGcYgx47GJTJw
kH9Eq2/wARjkC7Krcz4ad/QHDAxRbtCpdTN7E8B+NBkjpCgnBWcYxIjgXYeL2ZASFlcjLOntSakQ
DEhIF01fyD9A56br3XkgpNDdMHKqlwA3GJZrcMklKtEViTvO8xJowgsfLHhKJEh5YxpZvckBhfZ3
gfrrb76NpJKClpzPphxDYrSuXumgo/oeF9jC4HMLXHtneMTtYBGwzYm6tysb7qC8oQYiInaDmtjg
tkDSpdraBdvTXO0CsNGgO7l6l7r3A87tsIxinrCz0PAbJPQG1HCNJ8xpe7E8Cav5TOEXWsmPWKwj
HDZMeSyYgGEtW2lRlMF36lmlvPnodBJ/nKqCPsK+MYrwTnsw5wxgZrBDGObvYxTks41ShoUdSE/5
7rkgHanBfwortuez9ExFln5X8edIVQGeMFzvsU09OfaC0zXjLOSTvQSwDI4BJW0L1BH7UXPvoxB6
GUcu91UuGdkm2lNKhOwqps9WIj5ZbMYSMyXupntqF7BdoXsSzvOw9qpTDE6yfg8Rw8dpronG4+ph
XprHS/623w67YKNCNsvxuAyxCdEzr8YyQ3gnPMU9iYFdZyab+rKThudD+e7AGvng/KG/XW6Bnxek
lGdoj8hM+L+gxrOLy914yM8/SLpq2fKrKuelA0SPH5RvyMTiVr/HcPXIq+EANnGYOYIuP6fLY2+1
JVNy71MDBFpDztcjT4tpvk2TtkWFBA4f7QOUgnRFSZv9ybYvaWgYRn1S209OEYx6RB7mRrNS5k9W
yDuo5+IYI2nAjrcGjyx4x91pv51f/Q7H284Qfr//QVloPWx2WItA9d6lDXQ+79p+wz9iUdQHSXk0
vrIWPqvL6dwHTInD6X3tnJI5DtWfwDDiVV5Q06n3/pFLmNg6W2HpRv6gSNsv3Alr8836wX5xtZpj
V8O035iodwNWmvR4851aM1T6rTiS0Vr0wSddvDheel+8yCeNnT2EmQpGVSIZ4rMHw1tlrygxh6eH
15igNPgWaXfsoHc9j7EAJFHabY82j5A2UZ0wqeyeDhacYMz7CgYy9jw6sFH7NhkWpWUklcPnhw5k
SUnXVO4yRn7FvOAQ7JIPWVdyahr4GQsZVBtPex39XKW7rGo8YotvPFaxiUi0LlMfDryw1tbOVmMu
8UomPTd4UYfjLQEQ2qZE8OCGWDwJ7dt1JLD5DIouplgtjWGmKTD91wp7lRR8R1t1T3vrvri7lxsJ
GIDjP+iW1nBkFO6DClnHGC7WEnZqZMAWzM07/wt5O7572kCDci7EHIUVXeN+sAZNmusrJz7mEqxM
9vuFOqrIfVN9IB/Awi6LCtX0dgqE2Gn7WB0u5xGrUWHPgwSBqfQGboMAdTsFCEzn9MwXnD/equxV
P7axdMtoi6hpqga5aToXx10egDm6EzMeoFa3hakrFu7nvAiQ/dvlZQqo0Tu7+O8sRqnClOReIafR
S+zXnsFAAybwvwcW/DafjYtAllxTPo+PBERmT4uL0ntSlCGgYXNXFiuJgWL+AqdaJth501NfkjRe
USOSn6gaOxRcAotczeyIwkMcg850O2MEpJSm+StUoRaVNsOmj6jOAxiEex55Ig+Au4euU9kxEJg8
9EFsNzLu7eabN10tkjN+iw9UQPihwSOerEzB0eEmK2yJiTA77D1bKbIt8Bb8xNznXkdCTuaoynCO
Tl7IS0tfxLySQlIuit4ASV+BZxyMa60VTScW6rKlB335jr95hqbBZC4P5KS6LCy4Tp6+i40BZfHI
V+bMrJUTsTKF8yuiDINbHy0jaRve/Sb8J9WrivX2yQI7IjNtzJj9klMqJ0jBdHMYIN34Fc634Rp3
ap/YRd4aUCegAz72pMZl4gylBvwp+kBBNbUyKdvR88NSvgeFwZH6gyAJN6D2wUVUoaNbNrRLzsQW
pLSUCfnt+V2IQLyQpck1Shpdy1z92jrddHuafIq2Ix8+1xuWJyhQt1TxBAHU8mxnJZZpGk6Eq1TW
t+yntfmqamkGN9JW1JjJJBmBfFCT0vAnTeTsLiErMsQs6b2WVumJXU9VKeOhmcgDV50PcHCJH348
TgtSSnDNGGvjKhFxKeVjxUKjjH2wMSU0TYjgqnOL3V26Od5s7DgPRQknvi6tj2xMt4+n7uKnnKqR
8+kehDgawctXWZ6z5OX/GF8+YiIGzpzvWZFEFqdpymcsjqCoPhx6Fgw+4UJVT0p92BzKnUPZi3YN
ggQVhnfqRpOmPp+EzXew4qOixkuYLXdz67X/A/LdeRcghNxvdw2ykj1OCjObzXBAKlRQ3cDJmRIn
kyEsR3igA4fLCp8vyA6ovkh8UDysDIXXTAmv14V/mwxdeL/VHDtHJgJFS7bOlHGRaX82c+3twt2p
2CUZfYAn1uQ38xglrCH6owkpGEz146vwfFyWnRMaOZ6Ub2i5LAoJlgXqywmk1O6JaRsRaqj84gLG
ILR4m3MU7a2qMzbHWKUiVYKFu9GFL9laasbxSY9rGBiG0fFObJhV6iac+Iy3qu4+IcmUqVdMSbxl
s/dv7nZNOSmFJUYvce3PRC17w5GMbsmg4yJofWY2LXYXM23Ac1IpOFEsqU3xXzZVeX/t7NFr5jQI
quIY33mgQOpGORCpYHGaIoVHVsAbrQomJZ4cK20Jpmxnu0tkHalLljNTxTczzB8x5vOXU/VruJjD
aCH6wz9u3ZP+QKoCwc4KyqgMXg96QAoNSvIFP0GMXroqNq/A8ehj0xltp7emxzKNON8SMIUYfayl
xIDa+uX2P1l3KQ0L2tf5RKRKBL5H2NOMGKrmlXLuKLZMUyXtzyh9IcbW8Ws6iCoNd+vdHSYnYm8q
FH/tYadf9IhIW0stZj5xGOHTICdLclhC7AqDdGEsLJo2hAX8ev2jMqVYG5APKK0SD4qtFLD+PQ+B
KyQLy+MAXUiBm3R8oVBTMzotMUgs6DnymyVF4xdfZsMB8P5HbBZkCDDhjFXR72nD++I0LqmcXOdJ
TVo1FHJhTOlkrspQ5A2FXXinzWnuhN2XvtQk8lqN1jOyN+wVbO1V1q3g5wvRcKIIlfv+LgB2CemE
7g7QKc8vYLLRnFGsCktGlEEB7NMwzSjWOL5MbumQXieILkoGc6bwtQt+qL3o6GjcyFFChnNLiF97
0elk+DmummdmOKhS4q1nBdKo7ZEesOUF9tHDJCyH5fzjbD5U4LX1WQ5Iby/EJqbyPdy0Mm9WVb8G
br6Ov+XdjOTI+RaWMVoJc12vwqwEmNTDbSHR5pBLtrOKG7Sx+xRCu54AeKmm1TAOo5uON6nBCc0V
Du3axzavLokWnGEcAgIKHD3MDzqbqvM7ObT61uUk2iJGtizVnp2jPUsht2nSNw2hrdsIykUI5Qtu
v0LlkUtn33upFw2kIFcFlti1NkJ73XjZaFoha0UadIBdj20FWKcU9MlMarIuAPhaNh2Sef7/omTa
NjD5TgqZrS4cS5yQ4VW3DBuzTplS1xoqaOJ+CuCFws5oMIfOyePdsaTSafgcJgDncyYrYy96B843
qzCKF4jO+nHfCOHaHFrXO11CnYZTNQgSOxeHpHwpvdy90pzTE0kn+kwu+bvG2o32wbor4FighjvF
YHiOUe3ByPSa60HGUgBJRoUKlGJ+QLvEwJ6hnWcIhxr7HMqTAn2dsXWhdDSfBhGvW/f3hCo9qRlO
qwI8mByVJtjbgydRYZ8Y5qZhf1fA0jvCFhZHUSVijlNVH+G8ti8L+LfS8BwYWTFIGiUeNrmmg+uE
h4eTNMBj0wbxrACBcBo0GcYnjxXVTsxvtCW3W76c0adgvfM008ZOLIYOFg4u0AvDy31VBYnsfu1m
BD64xRWUu+CV7RLemekjqLVAyAO7Z/8iWrpUQd4wNMAvPw1uagEGoWVCGpHYqKHpkL4/+sv0DSjv
dPCvWx2iJSu2sU7OZp3jRc6V2vaqAdbdcN+M6iip8Rd3SuIIz1HqCeK1iOhrvWxHRSegMYMH4nL3
ok9i4syNnlZH8LbT7i6CvLW+/NDlCzpcBe8pXzt9i9lvqgzfQ8dgitoR+sFmczjBXCS4Dg7EJL8R
o0z1g6ZdhpILyWvUMiZs5GYpAISC8LSqiG8lU8k5onO3Q0g6AVfJMuTvHbaD11mPSe6pM6mPNC2D
Xg8YsAAzhNs+fEDhwvf/jxHE9zQvHVPVliUpZ7uDwtP/NKpxEd4mHdCSI8gi1w7xoJXHV004kh3e
DE+9YHTszBJILb1OB/z5ZweHhjjjGQwH19Jdz/2IIt71j3yCx7Nxf3Tz7IITyGnP8CZF+kora0G7
nZWfGva64hG8r6jGJE2Glkee3MQO0AvoQlDRpa0nypWe3X+cRW3jmVC+m7cKRPXb+YeCmLitYnhJ
x0AkHhVOpW3d2egmt0MJ1Cj7Pjb85obNl94C3SDW+pegTW2ee4RkthZ3M87FKXFiEaPfX5qRxs8x
plAcACSWFa0kZKAxVZwl2JqIfCI04hzNzF6y8KU0CKnfc4diFGiF+sx8E/QRes3/Q39uZ62bGGIX
+nOhZzqUJ96Jzz0fTyUfVccwKApR/5S2s9v42CxRveeQNy/7kJ1BDcUcerPIyyZ8qYJU3U23vA4x
O6dlm96CDWH88SqgMQq+g09AKEVfWQj5+wfCu4LtdZQS6wJDxi5yik7QLBfJuWk6tWtpgFvYEKHT
0ylbp1xUyl3+n/bSFgyzlxWKUV/g37arwaVo3GmnhLuj66dE2CCthnzMWZcf4Rbe3AX4U93o1VPV
Asmg1540ocBqYzP5JvP5UY5XbwLIHWGleTv4eYqz8w6zR+biX07p9IDHgkcq9g8SUXnJWVgVVMh8
XbxUZ0wnfprj4Co2sapsAAlk+sUJFfNVP766LuTyZru3RGKfDZ6O573g6PJ+3BTNzGKhh7tIoGYr
MSkRValhGeK1DChh4jPEe7JKZUj+RUtUZzGkLQRbiBGInXpBdF9oDm2gaosb/0MEA/GsKVeSo75v
7l3LZtUYxAV6cz2/YFeaU8WtvR/M8Xf3kUe0BdAx6ZbZh3L3XzJ6FpxQKemiJiO81VL8DuYvbth8
Pz1W6jg+HX24iVMme8omIaQmB84oYDcUNoRjYtkS01GjbyI//7OytjNWGp3GVx7HtQ/60Qk8z3bj
uHkLenHoEKEd9+HbvhNtYjKjQtIygE93dyKZi5sGhnCJ45MIaxzroTxlfMpNuSksAibIeye0gyP1
CMqNrZijqFmQ8nr2QOB68vcTKMjmnBHzuHeq/9Bz3I0/qHA7DlSdNyOLJkNIfJxZ7/hXIiDhANhv
Ex5otUVtd0DXVQeqTjb1S1mn4QUkJHV85gimTv8yk7M9HyPbpJqnkI7IAOBa/qkS6Loieq5woxJJ
O8y6sRAt10NIOitej02saWmaajvwfGeFrD9Ws0G7tfdBWzgNTS2RU0PhRIANfGKyiEYjMwUSTLZN
4omXFGJRzYdyTS24C2SLLowmjreUqjS+0JTR+Aq/XqTGG7yiuW/XmeUgikhcVMp0OjkWKylngATx
5hWlMuCR5XDRmzWa6c9bYOeyttBOqUaa4cndP9Z1sfku6gxyNOFv8aXNfnaYCuO95PqXs7+5lAMY
1OuPvpXFxmqIGSxVIeBn+yOaP3VY7Ipcz2nGnObuBad7JDph3mdhkuU/7lD865L8zfXNZg4M9zZ0
tEaPm6CtoA1wE36i+1s/3ryDcmkKeV74QHSKgp9vzEPorJIJ0WYabS+TtEd05VS6bh6GlaZaPmFi
aweaVTAcD+2z6P0+mwtYZ2XzaXHy3mwC+B5CbwnXeVzQEi7OoMSGFKDWhVFtrwthJsTLbvj+i6Xy
tVzeUwjr77kj3UdADGzWB7qgkSC4QSdlZQhkELWrCOJZ4y8AEKE3+GgZUZMer/eL+daoGp9ne9Hv
BAJBgg1wKjnCnFyPB5SNigNkGLlMhisXKAJ0EdoStGBHIszC0Kvm8vfquntw2kkRTmVNlrjUmdrM
kPsZFlN391g5dVl+x27L5KFXqEqznl+N7L6GdVlPuQenpjqUL5NkDNIDzoPNsizg4Cr1hrhDsbhq
Oqvir3qrmCjanthZB/6twpKKwhjMb7R5eh7tHVFfoH0JMA70Pd9UVIrUtDDps3qEyp8M27DcrI7u
lSR6kYwITVE+NI2UNNerVEsp0mQxXpKUA+ZUVvk7CGGaKrQcNODbWCbkt+yBRoYk7dpqOVVHPJ+i
LEUuo8wT4nt8TRxOYT+61FPgG0js1bYLjCEyQGqpX4+zHittHYY3gzXhMlwwkCMUA7odOMfzP1PG
PuvO1VpKu7dTj97PTx+rbtOcL0TE8tYty5K2NwleLI9Sp6NNRtrsdYjE9fgT5pwU9uqiFVkWTlwc
aj0AF7IcngbEKiXV5cQwrOwSycpNoiItb99ytyzgWd4FLtINNKwPS3ELc0fXgLqCAlCYB1D24xyV
vZKx8mQwHEz7DkNZZhlJSZ2BOJQRQx7V5hfyGNpg0Plrw0Hc0vfNMrUD8DdPso3CY+6tEtINIjSb
oIEXjPTvdkM3gRAa5O38tapZpiurZBwh32U7o3n6OibyjKTyPXUxBL/9rQreKzt33q9/BxCRp+4a
T2Z/Wl21Q8x0y7rgpT3id+DCNZRozMcsaR/LnwJlbvyhFGOqT8ZNOfA6UrqQXlkBRk67soqY9st8
/irwyOFm5x9XxIvZVJongK4tK2Fv4s7OwmbyAZtGl2imeLO+/C8HRpZAsGU/FIu47kg2Sttzj0vz
c0ohODGWb6qYYvgIlEP3TpfJQtis4C6udm5dlIGyF9EmnLd0nWsJ1PKB+/XYoWUbC4eswmrUrGOb
awkXSXFo+uvkgItMHWI14WsgZinKamIcA4+r9CzmAZrR7CRmG7kGSnGfxeZr4Ly6ztuNGZWxZpQ7
cKr/Me/EeSvK5eEJWi1t27as9AMro9RxkIYpuqPTLNwyicBDX/nvPT5T5PIcxHhWvM0sEof9zm4l
yFjqZbBFwZSj46xfJGlFBzr4TVjvP9TTPBc4YIHIbLEzLHXG9ZOjXhBbm2p/Da3YDTAseThnvYql
Aba5nO3nFdBX7svycmT9lRILMaqv/PJqNsE/QgmlS6un7BtV/PLdSuhqrCTIH/aIBUVhTsWFds5c
/qn2n9FnX81GLS8AM4KxFE52wStyqnTsptxW4UXRlF+Bdt3LUZ7uEXthTiGQegGfWJgc79AFc5QL
n7CMDj/zguzo/umAPAWZI90CTn1fumeAOdMXPo6hLlMD0GeA2HQ5SIC8b3L4o4lGBhiZUWWQr8gr
cycc1ClVqtiSjsZ/vI70C40aIcVEBEw//hrikzCYSAcnd9+n7ErvQXM8OJTuNR80gbRjhE/ywoU2
p0OgWMdeyx+HQ/aFyPdxPe2P4xWG/T68ZiioFOPrqjnj9bZEOXGKCiky/YGGNn4nb1Tnm4w8kOEK
dhjEuxxnKYsttH7iFlBOGfRavu8AA7d1/mD87zPXT6FUkvqLvv+UU5lbw5yagVIKFEqg2GbIzOyW
qM39Mkpgw8T57BGhZv+D4YFpzi1GEpqA9ZBbiViFSZeunJJZYz4T2AJDnFljxY6FKfhqG0JMR3zS
9JP4kZduq99LY0lvONizBgmgMParfEm6PXd6TpJM3fDPmT+4xbYAw68TzADjxqbpHJvYjqkznK5r
1rvZ1LQc4m/bTCLcdQFOl9umGVDMqHWpZ8ppDwos3ZWQS4JHGMzBX0s0CwyY8PreoMTKWMdpR92C
KlSenMnqNpdcNTGfMVLHMzxvYjRYRSrM1gHYOd8WaDCZIjy5OTLvKSazX10+7WPdPi244tRwdDiI
9MDzfUjXd5zRQqZ2vheQ8611kboCbEpZMcDDPl8ukLvVR0wxD/qsvuWN5tvZtWeoCIn8EzeOsLmo
+mGmWFVu68vflSY8IY9Avox0qg825wFaCKq3VRLddDcYKc3hgf0F3vowZA4T8amYuMn432aDlQGl
bZrq280aJMZ2RWlMnqSc7jT3XOk6b0TifbR+yYJdgsijcC9ScuasYx9fN1sGBnE/x+edaR6/wYnE
XkkpDywJO8cIITI7M32/5mmYndq9bJ/33wlS/2R5ZPaNdIc+Xk0Tl7QUBw6DU18Yre43T6huQ6U2
WtrZSxHKUxtby7yY+k1FHFTr79bV6hn5aCfRQaIun8yDpDya9NE0bvXbgM45Qfk8y70pWYgkRIRj
kfLLPzKRj/Pm0M5RR8lexbehO+O5yvoSYfnLvW4lzn4KUZITOCqLUpXo+CpRtRkauKgzMY/Tvfsi
nfPplSNQ17dgHkaGiWedxZtet+PyKIFDgumPPbgxkBfWZDYPmCylsMcyvLBiUOug3KbVKWspaC7u
7uwNo+JU2HUjK03SObNMWBiRowCjTcikSC7JKEXDRz6lg4OzEM1OkfqvY0nqxKmTsC9dHO8SWyqg
0sBGUmuNjQXKMYlVcsWkPS31tijwKHGgozQnAg3vu2akNgM4CSOemc44m8oYElNB6uJh2oZ2EEBQ
B4wejPa+7jHFZ655bXFmP3RYqxUo1QvbpaMZDp/zMI6uYa8UxIvBHJ7Z20ZHVh0tpEPidueaQg5V
CNfGL6WDnIfHdnpWw5gDHPCn4MvzIaxGmzrez5SyKUBtyMKuo59US4MKeLS3Dc3quz6FSgADlcuw
2l/IQt9TUh2imyQWkZ11xzlzgLcTSpBtAuaritauJDA6NVZ5nxQ8Z/eUrhXWk0bUadVgVS+RZF7d
nIxWHcxe0pQv3zPz14x3anOrBk64OwLiwCNtgZx5DH2HTaO5rqGi/OAL2axvPUvUdOhk4Dg+zNJg
J8Tm3QaKth5jrZqnCShwEsgRR2FX+FMqk83i82pjQDnd6c1oDy4dh2CN8HpEtSnF8cZaGknXcCDD
baCTYjubaf4OYMqPv5BjPbWSr8RFWiG+ltgZHNWr8R9PMePde9ty5idKwq3+oYOB2KRmwlCX8EgN
R19upGxu74lho36z+L8kd70DnWcNjvi563OL+R1jA4TGHG0XscU99k4AEHwcsxaL8JroIB8VRVPA
LHPxerMGntd+o5Mc4hwq62gdbEivaAipzPC103L0QTMSoaLmJPFz1QGp2eyg+WV3P93V6wSENhgu
/rbCuLVFw98sMYKh1a2+5p19PfDTzXbZ1/1g4FeVCf7Y6uxwiEYjMdYZUx/yKQMeQMvN2C34EUmR
+LJBV1+dYd3CjnPXDwDtTDqYaV8u1NG90JKtn+9kTOtyfgqL/efGLjPxbll2PhdDfuBNXxlUIdrC
tHZq+rwa6IjYx5AfhYy692YJ7XlxzAC5kfVrwrSu8Sn/2K9uAuUgkTQK8Y6w9iJtLfRcXLtPEpTl
8xkzjdvAAoj0K+ZyO9SqUDNHgCloI+KpAwwP9OYj4V+N465nmrcJy8lrq0Ay8dnxpcKRL6sujE9e
wf93LlnBm8sWEOgnXtJqwc1jQ2qqp//4AxZxJFCiiAEQQyKUKst7UnaEfKZsh6BKdc30bMGYkOId
v07ucowhFFnz+lg3ePyae3P8UDwh6MTnCj3tZ8biz0zZmdq8g/oITDp3u0Y2YbEGc+9We0QUMwbr
mXXFKvnfMVOzTSfI3V+3aVBeRWSWySa4LSav++BZryra9My86WOoJRgIfqoKK8WX4NpnQGARhbyG
8/ysHr0CqEOh6bQexRJH0CuazqYr2ZRm42fTkd0W1WkOfjOWJHvTj8O8a04JI4/zCTz20iF/am0e
0QkPzMYSDDtoNkC/n/zim5/g/6WKtEPodRAReEA0uVzlqWnNJYL5Q2JykCU1uo8rrbImxB310MTG
vq0rTbmMQ0+lCyuQI6S3KJYF5Oe8sBNG7UQ5KsjrP9KEW+jWks2LuImPwZ+rtHUO+NRxX9TfVF1A
bE7CNKDXZLbevrVCzEZCQZByfV4UxsrnLMqSK/UvIiXNBbNhaoHnAYEpUaeImx9Yqvtn+uFTHWNy
IZmYUtF3JNchZT9q/XKkpAsWkK9HZDrMXW//svPlBXAaLqYrCn9VJ0noBVQ+VAZtCvMm1v39X/D4
1+TKtSwMzsw5pWojRlUS3oD/CCXRrq1cdByVyUaeiGqFyJYRGqFRnDsefiMEmtDHliA2Juux7car
So0l3OZW8KJDyvU57f8y2Ed1hPs1VojyYeF/ABxSAUlCQQ6fti7jV1ACfksM4TcDLZc/HxNnK0wy
geR0zCB2YmhfnpGNX/2RCZfvDgwxoK7QCtFm1fZFZWPLCoR1vvPKMPlumGJGgz8NRG4P9IvZslGG
3ouPcyel0XWUCMEcvgt//15pr5vnkHp6SNxekoMxn0qISY0/DU6emINW//66JkOX673ufJI2qgbe
CmrDCqDR3yuVdKirHM4QvFmSBVhG6XzpjZMQaGAUcDhASOtbjDDuMcmCqg0Mq3pUNhBji3RrL7tw
yhhtdUPTH21Cgy12E8HVxvciN6PjvF9XTVMxFFIAtoXLOzZeQJrZ9u876mTqTNvT/HT4DzpXYjiS
NiTZfJ1l8cRIRASt2ujM+2fRtEtHjBshFkyzF1KtPqowk7tA6E016aOi4MLl9hu63+M0dOoUUskA
UsMBEM4m+zUrTT24UMQZ9u46V+yTXcdp1MsV7hlmA7vIurHpbxV4g/H3UbzzVKwgsV45bZa6SYwi
Jn9crzPfgDZoyf1NDn7jAuk2TNvoom8MurQQ8X41tk9QglS5+lVy6R2wpwd8ifsJAZO4qUFxyVIK
UeSRjWR8VxdbRuQnAtn7OpCG1Vd6KJZJsNCvqpr/hzvQXhqSL8Mh0Y+0wR836vFw7qk13NXzz5Tv
oJIyVey2v6a9EpTj0VvRZomDsFH9v8ncFvvyVq7VtbHjYK5DyQ9vcdqcntvIwfjUa2FCAHK+2wPx
Lnolj6GNll/DkC/S+4pEML3p8eL60AfnaIqTPAka91VA0+WmQuhZBul3jGBpvZAS5zA712w4ApgQ
vIwrNB2l48kJgyM79/u/uywIXl7aqU3hA3n8KfBCZLM6g9Fdysf1vmM1FBV2vFyDbdfMyrLH7vCL
iscaMH6H8nBvqaUQzCnlcosUZAJ3QTDN1OTE9HIZbj6D5mSyHpH1/K85yIInT9MjVMyK8mBtYGk7
LYLTIdiy7RwtRbuBBNuxE71sD+jmpod8b1vmFMLXeixKm4BcNJY1zNbGmYxt2zo24SEQheFACppV
CzVz5YTUqyMQ2Tc+V6KB/DlVyBrlo/mzI4/FnBpi8OiBJv3DfYf4TEDJS5xn0M/swQWXWAPfkS3c
yQCI7jyMoQ680cY6nySka3tj5ZdS664LSgE9RePz5Sh3fNYzlkN95nC5gnW4HGXA7wpBwg/S9s4n
zRji/fhcV8ZOVgVAtCzxQN/Beack4ZWvYf/4s3ONcO2qqoaedo8I+BVFxtxK/aNDFUk6vHpjL4yP
TS/7xPhlMn4FUBdJyXxAEiKAzbPjVMV6WiPIuwO1mGgs8jcfVaWI9uDdd5sUJUmJUTJj6gs4rMpn
FIoeDUvNFlgSLFg5QBSsBdKS29rDlVIYrqFZEcXsO6Lc90r8Gy4n8sp79NhCEHlbcGZlG1VTxrbE
5p4TWT9h/Ul0ont049G5xJnfYspSbI/eEIWXb19CNXqahJm8ZmUXOs2f+i36g+Rh6IpO65+kgjh8
uBg/C1khAIYyLVug3tgnHy3w/vgqePSusoM0zUSRhn5ddntD3wMfcwyFhzFZJGNpoIsSWK0oEVOd
RVT/Md88d1Nh0vlCigSPZN0EZsmQpQ6szIVsrHqYla8Z3JVwpIYwgogU2WUrvy7yZ09RcYG/WBL5
OqNXkBUB5Ip4+PUpBvwD6nSt1rwUnVBwvf6jvMLuvarpL1mVDOO6npwncxJmPaccJLDUGqGV2OSg
Jfxo/sfgo+hIoVgKRA8ENHi4aE5BPqjjlF8n6n02L6JPXzMnIaqrhzH0J55sbCBYllA+U4NcmbhD
Au7Ehsk66mm3YXiod+WQRNW2ceO2t+a1ZIM7KIwWgA8b757rgttTbtoVIFVpzloHMhHpfXT61nLw
MbwJhoe3fDsiQSGBo4kvysyhUVhURpfRiORISHAEua0NRf+ZqojZKAtQ1fFr98AJZaDdkQWQfUlw
3lnwWdgivK0b/B9cd1jMIwNW7Xe0hwTEcupy0tSs7SHJNgMvFqLKSZduoAyfeGD9CfE2g79GKMJN
uMk+OwORxNYtj56GdLJQa5Fn3y5dR76ae5OSi1soT439H4qGRnkRLwhw+/EP+ixErAMLJrZOaBLv
896iHDIv1p02QBuTO4dklO13yoURSZlM8aX7at8Ft6mAMeDAYgY4MRBae2oYxOCQ5x4zksqAWHEN
Xtp7acDzfh4P1cG9m8kO6ZPRphDCBWgiO4pSRr5fYU/VIRozcb08/SxaY9Be0rhW4hEgbDHrlc46
5TFNyDu8BqRU7nBuspAW4TU1f33HsDqzYzKCHtZDcxSOqm1SxnbGbnQ3mMxI4IiCOmp/Xvm6K3u/
+i1/XeEeySKefpHGlFYlXoVe+bZvFsT8w4cVo8XSp1LOXbOd3N+8jNtQC97f1ccmBogDkVSruriO
S1L4yhV6eQUxY+BbkjD9RLnYRPDORSnRDvrFBsOhhuddMxUGozZ0uGJKM8lnSf81OZjKKfGyYgwC
A8EOK0sCEBryymVQlkUT6fxZSoYk1UvY52M5bJAxu5uhgt+RJRaCG1OE7e20wmcY7MAI+y2R1aDG
9NZXN04CzB7qlx1Mfo6ifBhIkKyzoG2XMYL79TqXwXaqjqJrgd5bE1rqcabfl8Pdr2Cv1BIFN8Sf
WhWAfU8Shs0SpXmoaiKhzg0TasZRe3MoTaB9Ml3rBPApRjWINAiFUrJf/bLzemYA5eKkVa+W39Q0
RRS6StsN1l43dMjwQGSejlpvTrgcWKJyCFouUAkrMChg0ST+jLQzkD+BbbZvxxy4kSZbtSRnLwGy
GO2+j/D+HXVeIxcAXbddt8mC2vmPj7Tf3VPcoxekAaQcORULiyiBIE3vmNIouCFFSJarRDusiIQ/
l+IimUO5xNw5wliyx6XEGUJskCmYsxCO67bDg+sWbSexQNeaBJ2Bo4y+ybkNrbOLiuw5JwCGZoy6
4SQX45daxSfNQGQ759VbP2gDNvHa3Ghid8WIFmYi4+7py5ZR9ppWU75ofzjwF3Ysew23IGtl3TXN
jxjZ+9g0h29K2mARosGp5lpYJlw9cEaSxZtSN5ri/akScmrPdx2X5T4CAT7yFdwsRt6Dmt7KiTWn
m9PjEo8G/pltwJNBF2frMrUzRLykF39EIEnMs9EMi/pcpmeZG3CJYv4fLq3VOQpUYdeaqYLN+OCr
gK22SdI/4k3yOt4UON9VhoTdNXYz0I+uOBotcJ9oFrtu0Tm7yts/i5mm1MS+kUz0GNM/dfr0QHGU
SPSggNKRO8OwUQpGE3+42fjPCWV/HkOXDPboxDlfm9c8Rv/xO4OYkLG7M7MzT/ehGYq5YiMKD+vS
HqpGXgexw5W8O5kmJNPreWC+dLbT1GnLJyAiHCcNgEVIBeDJ7VqNTnUGxI9r+SU4vbbdxyeWqMM3
E+Iu7FkkdGRd2oKJIeWf3qENxeumlMiKdfaS/K6a4tUxDI/XjweTMg7bjtZ08lnqz1DCD6a7AyUk
s/Ywv15EqqB2uCY6KvoHBIdkFbqnx0ZJ9qG6YQnf62dLNg5R+kAH1oVcnc9NynH/zKFqeyLDOvTY
VwAohNdY6tFJIWeW/dePkNWTAqP+LYDrXCmrM8CojHjjFy+pERab9DXE61HYb1NKyUbPmsIrBP8P
HjtTXFs3j5J7GD9HxK33OMnIm8EffsOFS23DrmQvQApfjfL+0vwZ1Udm6L9bwXuGLhayvMbFdKzV
JKpDHN6oYJg8PEXcQkgmhxmQjIAcwXX+6JCjPbb823YfynBXAyMgqP/E2W0rRNJHGJ7T6MhY2OT8
1ESLpIrsfWSpxYEEEPfCLQ7nNG1G17DucTTiUuyYs+FslydpEOOvh2+swIMaCJY14iroBo8ThicI
S9hCk42DKDlX+92ydP4FkmEGCVMyQfVInadBRTJ7Uc5mfghMplWL6fSd32WmUC+dm2lUNSQVg8Ed
KNDVMwzIGDoyyslyCpwyOo6OH30jdYw4hyln+Wb4iBKdPUaQHjX3mO4Wrwd5iR0zESKmfHh3CD8x
LT9x8NhF18CsyTokp/1H2nP8ARZpU2GJMEFJtl1qUtEv1f9Rjhu4c032dBmXAqff+fIS8YPjgls9
kppXr/tjFtQ3ZPuygr1AxPKI/PIHeqP+Yojly/EY+xr/6nIBlSNnLpdbOtPFOn0CRunIQwwK6Z1q
KAa6MfLQTJ8QwUSBfLKmDo7fhTE5iY18PqM0A5llay73bs+0AQzlsDmMZ8atnQID2yNB9N0ohrXW
5slEd3KbVakzHpgDnMSj3dYF9y+JwCk6qxtlUPR7AtOSYjXkgiGuTMsDYJvant45FrvlOYjixNHo
C4u798XXZIWmE6idCVUEsqrDcdCa4/VP6eMsnSfXQ34amEX5wf/rtW10vL2igiITeDAMzirY/92G
Un6jN55gq0jCddB6TFE+LnfLSdiQW0teBys/8Sp+4Mmf7eMlBNJq4DhVJuBInmflmhw/2Rc3Dq/v
vAFpQYOcA9wSuXUXL9UA9wN6d5oHHmvYST2/YI4xr8pPXQ7+ycV6olhag4hEhaJcEEu0F1ZmGE0O
9J3ANlUKkkJkkjObOho7d8pYIbHg8UtC2JdZGDdEhTlN6WRWGyANfqSAa50oUPCw6z7T4I9Uwm74
Xyt8yXkA2pFiXxVptuuIEtuUTJW9lWk22T9UC6dGyXWQNi2pM+4Up/WjmNI+5IijschKO/uxTClE
BFxQon0I4GohBJKQ5nZiZuzaX55NOFTOKSVqtiG4TV6PA0NMSwwa57b6xhrcV/Zc7YD1fDnTWsy1
V7JqpKBVdGllqFn7TwHBAmF+57qls5Lpzb3Yx3N2T5iefv3Cwq/LdwbRNU8ZN/IC+qB0gg7n7p1n
sx2y1XQR4ipJEwyuyRjAV55oRvvYtfaIQdEzCmMvTTx8xyuawdSQqo5WWefByVZMwNeLZReNixOh
p5iUk56v7pi3COYUzMJ8j7mmgXbYHvok9iERwsx6nz+akq4G13csi+DHIK9oPMSc9KnK5yz7LKii
A/GmG3lGphmhCLDZuH9vblwYmRbFNU+9/Fg/y+gAgEdGRpJNil2AqLiPlPd7s4RFgNk8WZBzaNzi
A3QLShTfkzQ5+M+ub+dTU5pdIkLNPKfuIgenfF2nyjPGj2yPJKmxZXX1OBwrMXMwkT9T53sgDylV
bwRT8GaUQn7g1jfmnLUl5LOxiWPJF1gKga4efBUyhho3yfK9jD7UgxebZu2QoUzNzHLTVqWVFluR
UZCB+5HVdj6F3ZpvPdruw6xJ4gPtW8OLkKLcUHjLHwBChTwA6oq+NlcHFhai7waPh7L5DW/qUGK4
f9SeZHukCY5GxX0SZIxYBEnUEz8JkYPKexhW9kBUJVjl6yjFcqmpYuvB9rmFK4KVjFFl15HYfrVj
y/rV+q2QWHClRGOGreTSJeoyWpOfQ6L5nyeSSGM7uXdneQ5tXZKANwyicGDI5P8wADV8mcMnzFqN
nymhIvA1qIyTbPzWCijJJwuYewqfd8ch1VyYQF4rucSl4uGP+i5kBvUjv0FpaW+bUedgK+ZXJlXh
M/b3MIZ+ckxniBf8SQYx9OmKvAxupAc58Kz7X4dFbRG7KJbZwnJbktqoiiPMFSsUUSTvrBLUqDLM
hlbqxsmtu6Ifdvj6CwtC5nWHD3iNwb3CxaX90fGPsRuL1ZQ1QQhYLcewq+6KHAHAXtEMh89cfxXr
Rg/dNhWefSnPw0ov1zGpSBBwFby5ohMiKbhVPvPyjDONMWn86gNuxCa8rfVG4R55gmiXQV6yWxOF
0wQe08PrYzh5xVo7MV+YynEJaurgfJkpfHd2Ml9a7zvCGhhmHOHSAjL3mHjqqXBqMkX6EJRchnRt
inSWdfJNIagL78xgAerYsIfxYNGPHz3WLMthuWOUMZLuSZzZlb1GTiec5Dem+GvLw6R+6DKGnP+c
czjyfr8m8L/3HVPd79TDN15B80GhWW7SbQu8vsHUU6LUnkDUHto1cetc0yll4gmhXIwxzWM819pX
H3xIxI2Xqt4yrYZn/CkEo02AHqc1HUquTbvDLR+QRrT2wBn4n5AKDCq4Cydi9UgoGhU/1wsCxZ43
ZQcp2m7lCQmZ6jZICv0LXEFoMXc8MeT42+b124SFhBEgk1LHY+9UCkva6K65dRzX1oD9ME16GuFo
S69YrV74rSTuwYtIZNdnaPvqUIM6gXMCORsSp0FIA15BqLeL2quMP3RndqXjg+nfKIR9+O8QMMHq
2nC+RJNUaFhRylCaHq6ihnacoVBLmBcwzCGN8RyzcGfqrG6BrBJ9M1lCtD7c4LKQEZnutc7cn70P
X0NuE1pMdhCQpuWStGVIFuiabTyKqiiYw60N5T1v20EdkNeJPZmISzqx6zddEeeOWnKuofx2kVKx
VZh7Yoefaq3RNWPV0GnHpg3gNkRbDfkGz8TbROfYBgbf+cfcXvJ1BEr17aEQXHiHW0cgmLi2dMTp
xfuZx4/4FaXKgHuRN6fBewopg0SoPUKd59WOu1gjdQc9CmH0Z6+fnq42BmDy9zMAtRa+8zGk8IX5
XTvB5gvt/ajCXn07DOoxXkTFdDPAo/EjjKY8mY3cSEyuyqKgIO461CCdoQ1foFVW72hlFWEan17F
QMTl51LZCn3XsVxq2P69qyfiTY6kpC7gPjmmmCri9CQJvdPi7xkA9UKHlGpxUr1bhDHAyRRI8dqZ
bk74YELTS80ffSr9yCkV3uc3YaKyxXNJajqaj9BXiiPNjSj+CC73zz+qzqQ06YOCdvjp/VyW3Jbl
0XxHq9Lq9S8eBA/mexZWPswIbIxGuSlNaKavk/dOmW8gpkz/x6y81Y+ztw4R47TeDR9kiynkxhvQ
z1L5x9yQCxXOKl04R/9HHf6yd4pP6vHsntuvYMSUQSQmsMIDGKmuecXdN1NDvJ8fD9S1gscQbxHC
OrASQdqRDM/2aYuiCVxwzzlZvRiXV+YuZ+gOVwGtOoCmEmZlW7cOsPcoTygAXNfPAWkfdkO1So9L
xJMOQ0pBd5LMK9QwIIee7rFoKxBYW0ucbMVsJC+XtNBCwCdhuO+dqiS75lBDbHsVRmKEdBiwdRjl
d0mGHKEACOJqufNF6P3uvYEwm2Ek/N01BvYhF/ZXBMFfx59yxWkNEJJPJcOvQKGaozLzx5+qNatA
Tybrx3GVfy3ys9UGTPviEodPP3DcIgTL76Os/axXXWxvKntcOVBAr7whhsxkMLrT/4coiUW16SKc
zgi3WXvJChPPqhXBF19Kxlc3jdda6gnU8dcyS//56juCgWcEGz1imO0HQRvK8son0DsOMzvCa/7G
fhjO3iesmXPm9BiesVl92YumsxekdUQhlQnvaWqYOAiamN9Av+MIp+KPYt4HvF5X4eY5xbM35cEt
V0jL/pRIj9iHUKBpyuCtxOIU2aGB3EaBLhaKifchRI9CUs4K/fmNG9TtBv3qeMT+AIYE0aACXebI
EbI8P4ZyAvWve/WP6G7bIW+NbvZ6RoTouim2c90CsGHY1l6mUiHhvtgL7YYZmOhgEOHsQAvgVRmG
vryArqYuv9NYR4KH11pUePtWlN81fPERk9iQiZN5qr0PvwOirngjjUyBEbHyv3GXdoCm+0BTDlNE
XC2pGMOl9T9fee7lachfGjK4uXkTXR15mVg2zS95jrGXG5iXLLF3APSnzC884feBN+vbN5HQnvB3
O7Hpvf7SK02Yptb4lpTL+LYK8umqg/Yh6/BIb6jvAiFRFycpNY5Id+hRriFA79dbtvntRDKMIUd2
LpoTm+KUV8bC+xYx+3E+wbB2i0UbVs0qU700yFMwoXgCdeVjgGrMBoIxmzSdJCWJQuneLjtD4MBU
XsXlDCRgeyAutuIMZMvIAfpOweGFvpNoQdtFZGczOS/yonWzYo7jUASH7yrTX7cGofFDX7QVPKbx
kVBaAlA6CzbfWLVOJeJOX5Zdr7KrDNq9zFsWOeClGo/L39WKuRC+znSXcthLM24t4zftZeF2WaiJ
J6lFbUadl3w++sOKvFF6lQVSNfVoo3ogkLBuDrGDeopln2LhIm+cJFgYHf8A2njNdnUuspthG+qD
rVM2yKW9jJJvrQTX1L2L8dLnFiKKMvwJlvc8bxwB2/xv9whXyF6OJv3v5KU4xSw0Uea2/52M/8l/
OVfslJ4SMe7hhyxlu78rpEG5PX+7QzWTvJnvIxPL3kXc/mH8fWlIwFJW6+teMXyM+tF00mwOLGtg
PLyGICN2FSyA9jLNwk5QhuX0xv0fenkKdHA7lvpG4UkmgK4Y3zg8pzHyQ2TFPjDyiNICg2rSUKJ8
7x9FVyS+nDz/M9FZd4R7yod1jR2U+4W3+JugKn9OtHqF3JiSYrBG8k7nkiLGdL7ra9tUgGBQjWMC
MB+6R/2ULsTtQr1W/XVME7+beMsiGFDy3i/wB3DX9qNygSj/tLo63C5L8AnHK1n6B3QnAxufJLJs
+J7Bm9/cfjcqXdvrwxrJapBmBXmheLIv+O5cai5tc6zROGabzylf8jvoQJKj8KjOIJPliSeXWRhp
HyWXV4J/ap1dSWcHAIAOlFr8laQOcoGTqtWtKA5yPR3uqQR2nGJw3DTAmijk+UsNPWwghsW3zuk3
ZerM36+IINGLuuWbJYGyIMUJx+YvuigYSLV+mB7TSvdKL/8zA+n0miLonDaXLfx0WYkpWbgJ2hGg
bPZubKNvpl5hKUBwKHq5X2FrNymr485ry2NkDb2Q2PFkI3ZiDOOXCiA038XgDo8VWijdWL9geDz9
fSGeAc/k2wiF4UO6LfWwHUhrnF4wmCM5uWgUnudD/0laiCN2/SXvI7nZXzsL6+a6Hd+dvSlJ2uve
Pg6H0EstDTfA7vbyGiIVoU4jsuoYu0FBeF67BBblhAKgw6q0GPCw0Z3+x+lpxaVg1Md0+Ct5LbTc
gwCDs5OZWPuOGr14/LB195LjHwN1TJNaHk/ia1E0ucO/5mC2d8+wyp8l3xnZQXWGc1+hGFJjhNxo
8T2L0u5CqA5rQb1atOgA9JwxPHl/aahWc2Cp8IAEJ1m4zD57PejpKS1aLB3r+Q//WO02hpkplgKi
fKIPOYZQTL4H78UMYNQwZdNcIpWDqDGMyi3j9JNFWMNuyyXW8VXl9jaGU33pDdxAOyr3+st8G+2y
7gwbJTkiiE2wG8NHmdHpzf3ua1FDdbG9n1+JZRCqHlrX7joO0RwRmU2/6y1FWbJqhZpPWSplaBOS
HLI1Hupuo39cnn/C9AmeS0hikqBtbGbrIZWJPjBLtyPNT/skygQSCCmmxIC8SMNrI70BqeKY1WCe
3wbZoJW83ECdJyof19G57qDrflVRQNaz/3zrhAXVXIQMhjGNhIyoEFXBuV6NESznBUNsvkUIKb8d
AxCwf6Y0RcddfUEjIXXlr6YBPQPRyVUQDUrgdDGUyor2RaEoA4n7I96h8di3RglaEh5+x1TkVM1i
z2Ka3op6opyzLGs28z4v5I1dxmzEqhGS4M7OmkTasdo9uRnCoI5KCmgtaBN3etpgOS9jwTz0WgVR
gjWn0ZJyaOrEhhW/GKaq5bK54ciOMNW0gLqwn3pEMo/xQ9i1NCwcFuG6pbYPRvrC0cma571VOb3i
MwzZnawDAW2Vpcwp5n2P28gHJNsYAbkmvXvRTbIud65ssa5NTECz22/KkWMiskA1ITAaq4KP7N4D
TWcdfElGGdzJb+DZYUAEYMuCxz6hPXXgkWlsMrry/BJnzRBI/SwaZQHnBBEcJN1LcUCQLIH7rIxk
rrjnx6hKoM/E1StDlv4fdr2mpC2HGC7kBi4nyO3PJcREab0qafHeNw0V+AEUEIq66bNG0CLwDE/j
rLOtQpPwDzQOhpNwMk5ICKdcuqjzevqhoUy1kl6/Wh6CxezPDZnpV4U5yWbNvalbyz+Pm33d4y/3
jCD/reDTvCjmYpZrInh3/C71cE7SCToX/4XaqHJU3hveH8w85psWQ1wK4hzvzpDjLfFDgS+wsdiS
DtdnjwMUot4kBhXUh49NxzexDClsV6bnBnauUdkYxb6uIdM7JMT5qjtzvUQ+Y4QxLJ1ccjOI2Kpz
KNcMlplxUzLwSLRU6pYyVpPEW1rgQwz6pC96ST/D1+GMNAfQybOcJIDbyhKGPx7BF81OgRw2FSy8
ualN7z5XbRDkTm32fNqoW0jom8eA1JLe9Kno1qY4mAl/1hB4bwZLZGAuZpP4vf2valpc1qv6AQiv
Yl2Ir5qeo0fu3a6MMS06zFRygsemwMHr/CIKlkpmsdOvKNEZq05scUL092jU9dvhw8VkaQFbQk79
G+gvmLQY5TV/i5QUnSkilKPHloUImfzuuxGSu0A/qZbyWchtu1VaEAntrxydbWv+C7DoHXuRTdqP
wiXCrE7EDmJf4YfX2rW5rTZROXTDuwXVvTBQQnC+ODnrRg4ga1gSGft45kEF/6h8SKkCETYaSAyA
RP1D+UIHtZQuswmPZ+wRSpC8MNsubkesCNS4O0e3gG8JKVp1wr/+/ljeagUUBZLnOmyAn6V+khhJ
T+wJAIPCi02D0nUwqnRt5/7c/fphPAViYhYmbhZamNc/NJ8HJMW3iS/YAyWoAsq1HI+KL6C4GAy4
rx2f8H/ZrTCzwFHiCmSft6UP5oplcgkmtXuyxG0DmcS7WSFDjmtUEGYQPkOgL1kSXJb8UY33eppH
xNZzM4rl4qKxTeG/fv8SsZuLx+XF0OwS+MtXqZTT/rA8kcNzmT5/umkxl3hc9C3ZuLuHd+Y05U29
4gedcwgGUXJPzJtgQow9e6sVRQOOhjZvFhNgv4POPb+up64+kaBXKk7Yv+Uzisv6L2s2YTiQW0v3
GuTuZF0pV6LnCKVdnmUrFmD+Yb57MmUmON9dvq82ToTzWE4A+evaE0IrArGZntnZSCwwOp5f2or7
MEmG89Oj6uELC9iyxYXSShyiLOrgm9gwl8PYq35BYIq+qIEaC/xIxgUXbHhK8A1u5lBm5urpVDJ3
srrRbsThSAIrmacZHfWdVFgRL+IqWv9RiHgV1vefQZccFBO+245ehz88UROpUCLdTpWOCfquQnG3
Ef30YC3zQUw08IYu4PZwcWUiGmaL6NFPL4m1jVVrHp9gowfovdib7VP7vLAHV6kSvSqffCu0Q4I0
Srtp43HPZMINzN2yfj5kOJ47OJ4RcAnSeSO041Dopnx1PmHW3Jgc/4ekqrEx7jDkEfvkRBd5MIuh
bFVmQJ5cVMu0eZbcdp5QkUrS7JhVArB0GMvPnbS4OnA2CL8enlKJAcOjhEr0qZyV4I4wo4C8bUMa
8LRwhez3gdiXONRRMYasDzrZt7VEoUUK5BMFM0bpS6okruoBf03LDIHT22In8/IHR9dIB3ccdey8
T2yN5RUn+s2jvrcsXVU0egopFEs7E5UdRE8RtH+hDlAxa2s2tmqFdZKvwjwQDsDhQIlvHn+Z+JlH
CSJJ+uCnoGduMD4FH3O5HiI0mVGo8TAkPEN5NAIMk7gHR3QtsTMgUXdZSSf9Fy7s9OA/69G6x4bq
BB1ohniWsPUwozIC4LqU8ZTCHW6esOiohEYqx0TFyLgjq5YZVFod3fTh0yuSloyFY4iF7MeXHR2i
EbpZ/tRIRm/+HDtVrK6bY2DrYzHwBIOO73BUCs9B0jHoNIgfETGxR6BJCiL48HHbDGfoaWjCW2mY
pSDXYmEqdaLSmwMwTDAI/kS5drV8FYsuBSjcP+CU6U4EoRBMhpFp+1YN3YjT5b38iakV1gn7JTAW
ZKpDXNFA6ALuhdw73Hf7o8SRn1rGrca1EJS+dgF1yGCs4j7uuKz/7xzRJgMkRcKEREjaA3fhhA+B
UQxKscxeKO91oVkPqIIJNY9cAybPiBD7YTiBLZL6fvd8iHQrxESKvsRTMHp2HHKWc8YyQktMsjmE
5FUKX1Od14hVvVZn1wF/LMkkk+tApWPj72h4BKQ19F8EQKrhl4acp5IhiAnWCjFDB1ADgcRRGPf9
v2jg3UZcjE30tYYmd6F3wR50+oBwQ9q0KvqvJUjub4Cg0fzbjhixwfB0rTy62hXhA4xyqltneD4F
MJXaR/9JPQDnTolpacNeeLFxu/y56SmI68bHAVNVW8dsg7LhLul5SsMGsFYHBKpUdZ5YdW5pfCaY
0Ky2Dudq1PIuf0+9f6FTDWj0ZDmmsCecVD4Tyq3ePi7YOl0Pr907XSVCCLZcbJs8ZfMRYoC+DoiY
ZvHuOp6E0dA0O4PWNJ/gtjVzPE5Y03VkKifOMciTlniD6R2J3e6DdJgTbl/v/nf8VkUktJbObZqg
vh/rpNM5eqeGsz+gFdlPBARWq1u6ZgSl9lCQfjbouJo9Q0XNyNdTCRQJypC1qRhsw7x0R3WI3X6x
PpURVWcTApNFHwuSkn9AhYpMhZ/VlDF/2Omp17KFm7YGLbESI6clJK9Rps02t5+Z0hNUEWX2Cwp7
hi306jz7qf30ubb3RqotJw5N4yvozA6/g+IgCEyUNlxwnAwSIVolFgdyGI/pHbDnfGtpj7qSodj+
3StiAwe4RgNoU+XjSexpEwR9Cte4ismZsiREyq5Kb6l4s2peKy9ARrf7oXZa5/ybYMrCeCSOJXiH
n1rCJq5VgW6gsBSb1WSOZtmRMTo2kguCj3KYCXDZBAIu8RdN5QtvPCz/r0Pbeh9NvGg6owtHRhle
lCbGYCvCzoGi8AsWs8Cc9zEP59V+WCXlKFyvWKt3tC6x8hT1nmY35farJHOOAkEUMhRZNFuqhL2Z
aVGDKVlPjFvbFXtWID5tMWS8DbkXx7WEo42M2/PrN3AnGBEeOCW3GHvljXA4tRlxmXm6F2WjklcS
uDSTc3W0PdX++xHT8/dueGqzX+Mvy+L3N6UQ4irIh0IeJvML11EwLR8pUB3tDTZevTKoXJwWECgY
RHBjhE5ByeCiwSFgmB3f2E9nPgZP9qg2MIoVlpIkEg/kwvdLUjk23ZiWGzKhL2szsRkIF7x60zhN
T9eb/5cTbg7V8dQod73r37rXzQ11Dv+nCfHeOL8/1yIAhPAe77V/UpuQ8D3AmWeSjsTvsShox+PZ
5iyhP7GUNTvbH6nfWcaiGWa3EpDbk63C2PG6ffxcWs6KDRk/GdkMl3iv0WAP4IMc/aDDCOdvE3eb
Sli8UcOfw9PpO5PeTayrC2NRLe8Pt8WiNOeGZJQ6EacrJDUc16gFiiv3DftyYVKBJzQAmUNcZ9o9
XpU531ewvJSLqX3Il5dbeKe9QNojfB7tWJ2qjM3YBEkL1+W3gMWfb/R7tsw4r+C1+gOUbYPeDF6O
cIbs0pbIEJ+WnvIhmKdWwDn9EjhOoJxNRJbkcM40e50DTrJn+pPbvJhBiE5UyL6w+lN9y1KL02dT
7gj3P1PWnL9b6YfNX16QXeVO3FB6rIL9Fi7w3v1C+XNskZH3r6tyQJmYwrGnlgOFzyj88mzi7d5b
SK7VqMC+Owlh4YFztNwL/xh21y0xp0R8UcmcZlGBPEpH1YrtYGib1tuKwrLWaYaL5zo8K6Xo4r2K
nniGxAjmUZnRRiypMCKcF8Qln/5/zUobKngrMv9i2gVboKJ+r37HM5Idn9pWYgB0UZjVTEGwI6hb
bOumKIaWzKFWSmMl51nsmyQ81I7LvJbEmNw6qcSiRGhJHq10MABqrSckGiqxJjFDkLQS4OjfFrUk
NOVSiuuNaLeBjmAUstbq3/wd4kc7okQGkvs5V4l+HbOtsLmkzvXHINaGlt7c0wUqKCBDdggH/Yil
0QrNJVY+/b0hUTT8rs0IDd1bM0G4V3K4vNFfEk7Yr2J7m3e+TM1xwbvqLwoK9hl9G70BFC+w+2/g
K/u1VNhDZ80gelwi92RnFkOabJrrv74BJfkaEGYfqU/lUMKp6qguDypW+2Nwvr4xjQugTB/epGn9
51C1gMefhombxjhxkkISoDZz0b3FDI5XiEsYbKw+elbpnRNC7KylPXl19FAE+PftmSNE/kTwJ9mv
lgj4nd8yr2Ll2jaoajuLOehlwuRETUH3aKinugNLkZo/vA7IcWmM0MX3xIykXIpLVY2BlHjpiUv9
zdWR0vBZmF/hjad+dz87hfQJ60lKFqWbypoNCgF0nRIjKPqyMdjK92DsDo+ETXWsbT4HiL5dHc5O
JmAbSDOMBkHoECnGN/A3t+HQ7+jOQuYBcuXyQWrFevHOuixcziZgDRftJpHJ+S/9CrmZJDyksliG
6DqhIKVwn5kOIngC6XszzzE31a6noX3CMKGZMi13C2HvQczPlOeL2H5JrzNrqgHb/EPz3TPMV+LH
n0w24e8SQSkJzG6cDKWdSo+pC7KjG9eBON9N/VSZ4ASjoRa/1xwOnHC4A6+ZKj/oK2vBqpyLcGJX
9YGVaoNukBpm/Zym8kWyQirGacRBeDZbVjDowQQYAdbclPhFrURV0BjcwoPTm/Jiwt3tQlzV3Ahc
iw+h3s9GQXa4BM11WZ/5dwV93cDZHu89J3ZVbFTWD6UlR2bMH+1m7tFA+H5iLyq6IJE/gHefXkzU
v9ibq1BVVg/fiPgtCEJ+frpghenzNICoWH18Ucte/KsjbI26hhq270iyWmM5p7j6zmS++sx43FEv
+cL+8+TccL2+TMKqXORwNBLUBDYTgn7ThLLd8wJlPqF1c0ivMB1KyAnGLt0D6JxyavsZuxEBBwTl
w3oK0qBeKasw391+TRf8Foq8FZbyUv4mm/qfuFmuLKPtYpqG3Nez8osab84IOlA7UTdkn6slwuT+
YJwrgjyE7jQ6DsdYqT69RgAWp8wndyojedtYNwvejymTN6Nw4tDQXmCxVNrRsFvyfNcwP8WizWqQ
hvlt5AVYL2yczBSAYk+riT6vSHrxMGy+TwADFiDFR2GvY4h00NOpSLtOqe8qChOLoR2M7KBRz7UE
ZLbZWeB8OeHNC3LpZRNsdqXXrO3SrD2LqKukEsq7J3tM1gRWd1yL5ejlXfKASsLp/e0tTIBrhCLj
sMMmVWdQxXg2YuBD7YaTQHb+Gvb8ckVcYkz0+yKU6nEW5q99OgCOl6GEo2sukEipsqWXT80ZX9Ay
38Kh760Oyrs1OruT/TcbRsvJCzyd0DwYVuWawY8UnuQ2dub6AYK2B8opUnzsged2Ns148nV+TPCd
FLiuTm71zWlJzmm3mLgtQh8I4N6y2A579UC/uLqEPSMrY0QGF4++pS2ytQJis4ITvg5n5rZUHQWT
48chvJ/1WW6psZJiBpwGmO7FoRVuKR15WQb2Gy8yJEYVEB1YVICTn+BYno/prRK/rMwZ3ZK0TJea
hScVvFZjgCv4abeRv1Qa+Uy4RXomxRj9FHpql0JjIHXgnsbW6oX39G7mRzpDSRe6vR1g29WPeARa
jE/LIT6wVu1JGJWnMiMbqRMXwqonv2i85MlyL3ickwRK+mSVcSGrMnr+NoupidfInB/8CQ9IGLIj
Tv0nqfEMLjYA3rxKK8j2pOuZM0diHcDKQNWJORNv8OsJxBQuDtH3KIBcY8hppjTLEMX6WEXfgaWr
yioCm1wU/s1zNEaNLZ8eSWZK1E72atOuMkpXN5msIKVE7IWUxxML0fB02JcT01HqOAp58+NNbfOG
wOM26Dnteko4QxDDvB0bAP70DGidWX/0AAyVUZczoNcG6hwCQLvOR3hZNQMUgVCEmIE722yRudqj
A18CMsiq4r73A9qgp/OZOLe9x8QxyMGKf9f9fDGVjGhVzBnvhdoaNktA6D8XRHd9FZEqUwYfXwLj
vuBhTPdYpwm+nBK72cARwkk/zya5aIBCv7UEqOiJRwOz5PdBkXe4RVMG2eLmArINXSGcxpdsLMm2
kj7XOBoZ/Vv/t/wVm3H/AjgpVfIr9lj1V7JRx6VeRNzjB2OFqcRzvI6ECQ2/NYCedocyS55L08CS
i3g+fKSGNZf1EmeXh7wqjpHnBGE9kh0zDUOGuKXpkssXkbA3SsHy1krsrxsV1RotLFAx4iANlcCq
tIy9PTkRvMjs+VLE/M1l7sXoryDex+28C2jiPmKB+b3IDgi9yR8yvYLuwxKPRaNk3LjNMJcgo+Il
9r/BOZFdmZncRoYyG6FfCpMBIUemM6UdZLx/T4h76GoocGT20mDexAE1zHdl8zXQEtoYVin6hgx5
mIFZtZe60j+jRRb3JM1MGEnSW57WLikZTkyfcPCsoSggFM80fzs9qShCg3WasD7MSTBRfUef77oX
IrkgrkzksTbdKcXwbPyEmCD8qQgpVgGXzufZORaPUy71chD/aagAVW2yPP/j/tAiGGcj00/hMeNP
Uyz0icWNAfUrQ+sk+O5nZnXQdz5TxC3Bspk0VEMvyHWLbFB058qqc4I9D/SoPx/FIF5UpBjbKrYD
ZriGOOU2FGygy37TkKLjpLu98Zv+GXEsM4ZxgZ033Y24fgui1Zdn4/LuZEKh8DvFoDr2fEEioYXc
TvL642TDFOJMC5+f55SDD8K4pRUY9qgdrJDrdPRbVrj3uoQ+GAGQFYcVa7MDjQnwGJt2GJPUm7f3
c22+VA+zIXeFcF7gUDDuh7FIXeVeYPrGA2XCVWKx8j3GVPuskkivAbvqaGFfkjkE90tpqBTSieZI
YN0j/nEA4c2yfAtzK+/l655uKHiE92a1E2k5zRF9Z3AZuGuOKA56PcDrzmPNjjBsg3kxJon8hLfU
qdG4cSsvEHZbm56gakg8in8nslVsXbm2DO8q73HuUTk7BVJ2totjzcYuKbB5nQmBWZWOPqDu+goN
wEVhuWP325l+7Fq1H8bco4AwZ0FeNDfQhKQOijX6u+zTey23e1SmFaWDUNYneLFsMZwrFILCP7OY
Ud434sCDnw4VL8VW2r+GTfHVQLm4f6K0TYPh//t0yGnblWnL0YtDeDv3l5OMx3LCn4gfOeECZUfW
sJjBzp/3uw7fDjtvwyxZqOfd3eBKpY5keKOg760q2/Sr/xA/FrJQTOFLM0kaWh2Ctaz9Qolve7nx
Kd6vfGJ3W68v4qugTWYxMMGkjqDYdqI1miQ+ekETEkcL4CGZbo5Zzo4xUNfRK7tekp5TeidOJ3e9
ctHUs1yzTpSBxZE3Z7nW+HejKmR/C/08nzlc6n3NhWpPT6cEvFwvdhjbEy5AHA4JVBKAtruU9HsK
PRjPXAgjZT7D15GCLlr/iKNLo1XstSI1sNWPCOweUa0fE+eC1qg1ANuM9exdpr6FPzbfmGJEs+va
YNzQALffMle9UnRG5frpxCR6xpKj72AaA1l3XbDTSPbS6XTEZgyrLW/TKv7gUMYunCekCY5aoPud
Q83kDgKLKfzYtuqpjT3PhkCoQFOCRCeIKNsbh426WMC2YUqYMCCnVxu05r6p4Xz0LG7YSOhCoqPm
6t3OCdlcLHTfjwfh+memKTTjaCcuBtzwAhvARROpwoVRs7Pn3NrIQyBaba0hQmChabjsw0Igs6PG
iZ6A8XECxhPKk16kBP8SX6wMZ9lmuO2Z4ukuMYd26a7RN5bkai1YtNGjvQJXOf2PEJbVCnh1aeUr
kSykWLSh+wV31Zb+l1zRi10YEHRfdJCW2PM3ZkERM2IXwBiTTRAuONJh2dgy6rO03CVcr+Skeqcx
ctAjer6ioVHBMVJFjIXq379zirMMo1YWHrA+CKb82MawjAbyR5zsJUA7u2n6A4nzTBHcnHHOBpRr
6Qs4VQ1WwbU/2KcS0HQOX+J6mH9FLPd3jOzvLIMcOH6FVIsuZFWRRbBqeYfOx/9xaUnUaDyffJg7
y1V0V1URa49LO+IFgbL7BhRv/Wp4A4cU+BCmOhJ7/ii7CFGMfbZGBSeWWuWdMJI0WAuG64mSCaOA
RpzGSoFeNHjYO/s/+iYzJBfyMQ9O0QA7SccW4e2KjGVuLb9WMR38HYMvhyWmHzK2wA0heQP5e6s/
VRn5qi6GXTfPxQaJfagScmZFMdg8rsZegeyRWBILCEyk5CnBOG/JjLgOqkRymBKDpwhq5CzKeQlD
S8DkqjorASDFmnbBI7EqrACMraeNmv2A6klHTVuSOi7IcPJ+yGHaY0okJk1pzk4lh0zBZU/oDhPG
T7z2OSlyusCNq3i3vfaPnPBUlSDJibPRbVNuDUEucZnzpikFFJMj1bBOZXFlb1EpheARaRS2xZRf
3dDFclY9fzYYZ/RlqlNTaKOckUh2XwoQeyC+yGU1urSUVNnof94tn1LsWQNJgoNVbHVxDHFZ93Aw
/qnalmNAmdRB5wAkpG3tDndSmPAzM/Wd3AB8ixwvJIzbFHnCCvDVMjamzf6yolYfeufnTy2fuNdP
OwHN6WDli11G5ft7Bo21IT2tRJslsAnNHec4mnOPl/7e2DyYPl/9gcynVQkP1gP90opxyCoKUZct
Q3gM33o4q9U29Pps8/ezgzA01oawiaT3F67z4aNVLwyvbQR9eZ3ZI50qpBiMycu6MCtk1XrTAY3y
Dsl11Jsa48siax2n6n6804N/rNkVNM5flOilBtcZd7WL+p/yh7cSXSzNypGqvclj/hacMpEzsTCt
lcJK5P+LYo7OKwaXti7bHV1EB040s6Y2RXNEu5DyvjmGUj8H3ucgYwkjiyaNYBnn+kpUshmEUTjl
Ec5pOPx7AAtp2gfSNu/Cs384+FmhBegBV7SIYXZf1zS7kejZUNr7arkFZ7XwvNhMJnwPfLXjNXkr
ZbujgNWK13l6t5rzFdvwcjScK3O70mGoiK766QSRqCCM/ca6buKmTIKnL9QCKj+oNxF7dJyV0MxJ
AL6xeAN5Qm2gVNCs4gcsbcwdDlAYrq6iWoNAiESrn68COfOgAmZpRJ5wi4mj5HILOxKBs4j0QOay
9RAvpcJvEBOwIh9WcDHwJebHwsA+k778kKd0v11F316v2/arqK2CltJHH3gQEMdrytzSBhqR2xw+
5dQgR08LG+hoiz3D1jE+DYQq4e7Yw5PR6m01InEYamuCCPIOOy4xU6DWynZk7bcjcXF8ZWt181UP
plQcHr8CVxaqIQPXL3eMS//tMyiJI/q9OLhIcJ8qfPbqg2ikghc6lcgZm2E7zy8VbM4OJlNN5dop
q9fJnnoa8SWOQ0GQp6hTj35scu8P62wdjaJ2f62hJz5aSSuvsiw1rR9RFhQPDTPvgwRDpXsY+Kfb
E7vsr0ynqCyeSNuc1bd2Dq9bfNXC022HXhBClVuvn5bl8/w0JTMxdxab9AQuWvqBmGlFzzykfYjM
3oTfEZKYECMxS7wKi+S3fkuR1vg70qa8MJaggCNZ/Nlkth5aKz8wvscqzuk+nTSa1plWfoQBb6QS
3rKB4jKIBIdz4WPHRce6M6da8R4ec5j+heux0yEJ+A+l0Htsrch/cE5aua4qT1TnQFkJp3RAFbMb
YahhgpUkNwMzsw/MQKImV7bRvHIwctVFabXd1dtkwlja6+/WIZovdCm+fRn+XS3qpcs74omc+Hda
MWeceM7PP7m6RBFwJ0uTO3Clc741WA+etdfNyKl2PQp+AlopW43Ru8E0xCIz+fj+1yON68cOHfpB
Mj+b0zxwDEaakJvvI0PWEya7BCzOY0989zBOeyDsOX4fCIPpr7oE04VgSk6dAc55LfSpubeiRVUW
bZj2bGOydpBuBztK3ea27hjIAqUSW4tGUKdOp48TE2jqyTKgCPjpUbt8mB+A67zNi0Bjo8Teu+1S
19K1PShd4TWGu2tFyrLQUxNZavVYLe65UoaZjLj+yze1GhxEUhlCBId+MMlRhK+q1LahGlSH5PCg
yjUoV/c13CDOS7ph+5rbeMfYPkq9t656dYGZ7bAD01hMy7hq9BeBhtOcSUm6u8TwMFst3U6hwQgB
MC6+MfKDSR+qdp9YmWJtqXzEBtHiCPSFWuF/sWu6sx2YDVdEQFri2Nh9epYBb/sRQVCNgATGkICi
JY4rLO4ot6gDcLQFAicsr3PIh3bpn+spcq0YfzH4WukY7rJn5sUpkNgxzQhD6X0WAhZK7C8MqZrU
ugdPXzm/GxbvJyFfLemJjLXmMcKh3XlJ1ZVegU08DS5teK36Cg7xHFuboZW2ASYrEx+o/7ugQxif
4vdQ7fyM1MVvZI0L7NxLB6/vYJpkjUx6Z7uxiEtdUnwXjlo6OPUYDoT1bwsGzF7sv7h1YBaojPeZ
5YuFDyQOoJ1CmpbpXagtJRGaMYkug2NG4ex0xeEQKFae/sIojMSYV1E3ZstmQW3x8br65dDncP65
dkti1TCopxvo0TRL2ltAxk4YAdNGj1i4qPthM9JHQHHQWsLhWG//Z5w/bRhdzmEQ1A7RbdfbHVb5
4wo9Mb/HddWNHirLTAo3DHQkGss2qs2QMKzGcodb1wB2eqS296MbUps5ByH+kwIj2kYlUq9FtJ7a
HQFEiECuz8h3d1hx430BEmdR/SnECABCj6wodFnr4GC6HMd9oqzksRSAO6YHSLgISwIP29+zRvWe
DfxvnItSedid4qmOuRISjC6VhnfyyvRm5fjBdqzoMf0vkSDc1pTQgI7kjZnxQB6JHuq1anzk/aBs
z994BMuTf1Qkbomr8jWJC/OVqHXxsEryMUpy6iVdRX8VO5WSWrY61EhEz3Gozc1pFpgaMv1bzBE4
UHbRYecBY36LQ7Zxfyb0r+d5+N/B/q70Vi3jNAMq+b/8HTTsoIk8hrpS7+arO6PzZ+LoU/9RU027
+xWb5w4RpevgEJtDLuMHmcebPMDNtDJ2zCkm9Pq1skj45klSuAqvKVbDcPAUxT/sxAYrU+XSsIcW
OWjPCS63f/H9tm2DiPWCsu2ssW+/tjkDdN2QBMoBaW13y1I2IK2FDriduj6+Rp+qU6H8Rar5iNJp
hY9FomlD6aKiOMNEWbmKzrD/Eod5bF+tYUv1be9Cfco2B0CqeWWcCjqrO86D0l4IOC4RRkegu/I5
7DceUxfaEp5a3WTXU9w/tUjdRGDKMuibprIuqAa9XiHNfTw5gFrBEHhTdRuAN2V3zrUS/gALrhyC
NgjkoBb7fGbO0Pd/LAOy1oA+CQ5wibSh4m5FwifJ2lDLLhdeh6xK7Ki8mwsJon0ld0lN864oFJoJ
csoLmBMlbhaRmx+o9lQTWpFQwqpf9UGQdwhpcFfMy5gyQd/YF6jIWUZ+US0EpTanaGyJ3u029KOt
hExp158LLwTl8zaQ+twT61Y0/R7tscY3ltS9UkqTr6LlXAC63KaEzka4h4nZYL8GTNL03o2AuDGK
fS2l+In6vhFjQZ30jA9Rk6ZEkRUieJ3z9Tr6mk6O19KqKtfEIJD8lUR4tNWGX/PZrChIhfwn/51l
TmAZwWx+nI/6xBqIvMDvIj5aoIUEpi+9y0fja3iHEJJKX9/DWIU6W1UcQPODZCEQKS05ZWSVx/Tj
5W065X2Eq5D08cdzk+KMNTh6gt7miUG6SQuspwdq6SQTCLdnVdD7IPQRpfwjPxnKkhYRy1uxnWDz
+IKFfKAoaEE7/g4FqrNWsgXpRtokDavcNfgEBi2UlSTB8QivnKjNFDahRoxlL9M5wgkhUekDfSAY
x5vvLtBhta0ezACL7lN+VJI6xv78cnswqTh1NZXBof/Q9hEmPHX6h3/gohhxLGxTEQcI6hPE/hfc
2VmDZmeX1KAUjFztLXkb0R4xZv0flU1zHGZyQ7oRcgTlpzAXgHxvpSFaJVJIcFOQzgbiKMsEN9bq
8ZHaItZKiTrK310vsXW43YXUXXKk4qGk+SxwnaAS8COqNr5jnL+LR2QUvVw5YTTgSHLjYaLSMQ4c
lQduJXPVutTIKixXWi57fUC/f2byxEx0w7hKboND70bgPPLoL7t2CSmhvN8QPA/XOrYq2ZFDiMtr
LQtN5KQjwgErjcbfrkY3OnrDONWdI31WCBT7+VTcgM+iI5wzPmD+IjrvsFAlQlry2wRNg7NSdqlU
4I75l0OoLWowu8Az7PO+XkTkRU7Wj36PYLXho911QTbxOtYNFLoLXu31nrHmFWCqN2jP2dTkN9Sm
O3oVzlTaMcWW5g2tALPhKuyKLvSfrFdvxhaNTQP4SLJrwottkvuTyC1ywgJfFPHIcWGjNemC9FY2
kOz+EcrtQl9tEH+BOb1eYQNXb+ElpIaHdLBtXDDmq7plalZJ0BfRg7LEBi5K7IMQJbsK30zLeoQe
W6Om3xXmQkeMNzvaCTimKIVYjB9NDX9Pc20PvWJWLd/KYKGFCftwtVWAXqTuEAGWurXC284ljz3B
7+dFzNneUXdA/aihzW4wHq5Q0VJP11r1HONbvLZ6CWTeNZufjdW32k587Sx7BRJcZf3k4WlDnmgf
d5G2rc9cAmqmjE0AZZpSqrAaBjyOYjcwmkrmTFR6cKyw9GhWHunkZA0X7xHXsdWEXTzzdsiTk4y0
tW72+pC4Ccg7FwFIXWQKDs+nghj2KXtABXQpvNjAEIT/mvBvRRH5EV81pMoK6vhKjqZtHcAFCWN4
6aFt0tjTMJot/hOueppoj6O3ST8a151YujK7RuGM5ZNp9THBIMANfd8KbPbDTAD4wYefPzcvuDSP
RnBgiYwa0ZqxDthnJqdYGjs0HcZkRkb12OuwuARIK2BDsBfAdm0Q5MWUEhQMbRs430bZuUfIXDxa
myfLEJYKKyszmMD8kW7u56d5XfGhsZfRwpGa9h24WrQj481Sjt49OJEaLqA9iJCZ1SC3FtxTmpOS
JXypdD/Oz5bbvbPw6z9nij6A/r/xEER6us2Yep41ABWHEJ4O6Pb35JnraiBYj35iLVFW9SU1TYJY
r2V9HySchhvcseHiW8bFwU0MKPslnEYE6KjKGuN2ZMHzZd29VjnNP80zMSbq+xPSEyKz6i0246dx
+A/jp+Rpm/+deu9qCJQa1j4Zumqw/j3BspduSWQXk+LsJZEcnr/WxBz/yBSbZsiDAaKXFr1vmgcV
EWHH9nZOdJWpQ8n82h3RzkeFbQFr7+rliHV4ikqXQ63J2xaECDhSz9SEgOuA9S/KwdqRg3EBMs/X
dIScgXtitr4NGEOPHjvsPRA08eNwtiv75pPLowk745UOBliU3VBbI/5blNIAvlKauLV3xESBUCR6
Gs1Yq2V4W0yxilPGHIeSzvCgNB6MfCZo/k4YN/VJUX3TSqu5eWFVhVkoTcZkZ5UNmyTMbTPWCc/A
+tEsiH+YAILxDyP8RPFfgbMe1NdEBrhmTDE2IlVEA5MJvRN7Cdv3kGjs+SQwZAzW9MV7UcxStYhk
IoA436uqZHZZZg8OUwgSc05X/b/KC3lqj1221rF7+aWRlAl3QH+sT+9M1L4/rwjHgvJ/BgTZuD5t
d08z9OkZ1LESbFmWbI/texhtilAf8vCTljl/zXaKBcthHphka8IGvFrmbw1GFoNA8/PBCUmGfk6m
5Jh6tfTG58mmnLFm3gYPuN5MfjfTTXS74K4BmKlQBH0LGNtYscs1BhC9c+hT5wPfbTBGdDA/7g50
4AMkjEipEuSbC9FD0/a7zi+4hOSjPz0/AElfuV69amoqoJRCG8NGfHBnT2uIfTNiDO0XM1aTFEF2
AcPuRb0OR5LcOHEzZipxiVI2BtX3mmAMu9uUqUyB+qHaxfFULWT900rrWJ0F4l3wZ1XqDtamfSBj
aFu5pRmdLPMZW4j51jExN6J5sAzz70QA3oyon2AcXxJrf6WGrpshO5SQ5FHMscHwBWorsFMB7vYQ
Xi2CdZu2bORixaIcxcXt5KYzVpBexCMNuy8DPxOqmGUzjNI4u0tofsCBJqRCxlNbaE0DPYaz/GGs
J8eOrE61M4juYeQk25Bch7DeuU+yMiFtLtwZAIprFAjA4D7pzmveu5kTHd+xw35o+3nmPNqYtovR
xGtI4gxmcrnxm+tRVInq8ojZ/QCE9tstTtIsdcjWTLNw6Rdkr4l3+ClCzBgaYzsY0iZrI9UGRmfD
dxODx1j5t64TIhC77InOvQ9aCZoJAIuKveke3rg7xZCshEY+Wqphq4/epfHOHD9q1L2o7LeojK6n
JHorBKmx1yziVSGhsmvFNMoFZ600WCCyOBh6Z3uFwEPn5AmWTb69HAoNXT4cZjbrio94lnI8HW2S
u5LOcPbfTWVMUS7ahw1wm/2i8mMFaQwVUTkVxfFNDfo466g0A5wV96p0d+bAmb4OGNPuYhigQO5a
4FglMvLTDxy7Lj7yXhsD/wC9dg3rusrb0jtZ7PP3YNhAijFXB41bAJD6sKZKYwCCNSKJ69Ci1BTJ
kyjnxJgaLl9kTYp5ZiuA89Oc6gObvTpgJbUf6Nj+2CMBCE+IIFQkmPOFTSEMDqoWnMWZvXIl+xrx
IOR8AIfbhqqrgG/7UxFOZcK7H/VwrYfsGFoP45N8YTTelFKj+b6vc/ScmWXPb5jc8blq7S8770Yy
LC7dFrQsyX9Do5AZ6+m6o9q1UrIaZuyxO9EJzCmU2ppD3PPbwxEdwWour4BVmWJrqxYiVG+zdoFh
XXXg6FKH/RubzdR8DoJls7AEJ3fipkfXEbXfkhXxOpICE4Z5P3fiDqET3zCKX09piGeiiEWgGYhz
4+lyK+iH8Rc8uT3lzdxZNkC1p1aUWqoRpJLyT9MJQLSBacrM1xQk66QZyb/YMFmOuhR7nisbBOIZ
J4LhKCcJSEGXwPolv1dGp2exCHJnfFDSjNWMlnrO5xdcp9lGiiIQWJ9EqPHkeAFedg0zlf9Tl1t6
hbaX8xD1XVeAZxqTDmuNG55m6ZLbgQdCoERmw7JsUMdJog05Oc/DPEstP+ff1iyifHgJwI6XkkvX
twS6g7lUMDLTRRc+cbnoW4KQfVc24c+230vkS1XMgyAfYnPUG4rZXObvwiVsrW4EQl7cYcKnzhoT
h8ytFrQoTFOoNjj8Uyv9hOdo4EHkW/+1uVvALAAV/uOVemj53tSNxlWs46EK9khMbgodj2jV1LBZ
gss1wzjk4W/OGXu8SZqzMkh9HmLXtHgweKCLW37WIzh/LCx80qkMnskuCjEC+4ot37kgif/JHsGw
kW+h/zfPgKtQVKvcQCRoBY8hN/pCCnJ0TFUbq6fsxJrsugpQwnf4aYCZ84iyMcf5fFCmpempY0E7
DVQYKGQ0xELX+S16JBa8czc7kSqaq2qngx6VNReks3nemrNdFjEQWHEjruAlaMZzbFf2oBdRIk2j
IF9nB+k0P4Og5bpElTL/x3RstMRD2rJzLC16CAUIq7kUrhpVJRLDZDpPJoMgw16wlXeweOo7HLPK
hDXf5btrfu62/d9YyQVSZqjB1Xfqyz5BxVsYXogJexCvLHMd253qWtW7+cr0eCqAojV3JCSOl0cu
6iQQDhaQA+4oV0/fGYpAJTjg0RMaCYDTsf3qPGav9d+L3LOXLuOXEQMkW7T/JeypZbccuDnms8qZ
QrwH51ZvkeaRMFzEWMAB/dDBfZX/es49mg4xD/zVei2QifjNWB1zmhHMnXwqCkg5CdcjWdWKSF3b
zbeXOsHaQxi29CtQziLKog5hyyct8y64WwOM9KW/Tb4h4VKgFlN5n3KDed78kCX+ypYwV17OLqrt
NLVTHENVv0zHssqOBt80YbMgPNtXjgEGhEbWSj2yyEa8I7TecnZpiNcBgz51RBDNhlCnqS23KUiC
XmYaeBZE06H8T2WSvWyzTZD/WbwJOiEPXbQGMJcmpeJ8PXHwappLBOm7+NwxmS9ObQPvSg+c5X4V
l+4oMKauBoOikbuoj27dbqEqUclFzeZF774v/2PEw0f4mm9qNAfPEp9Kj/cVAm2r43kefgDAPaCS
DIrw75rFnTqvC8ENClYyww5Pk6jHlXiCCQzvUaVK660AOUX86f4S4MV53aQzUZIAAGR93r3d0aVU
kj1kNcJ7Vywxg6JL8nSBme+gqZrU7ddVXns3VimXHDnzSM582LXYJw2mZGpBYkfsX4AQ9QVPo1ZJ
Wp6YHUVrwF4hHKp374k3VPrtO4kVFONhFRMMLrUyJJFI8wBk5v74fswwhZ+HI7CpGR8jLJeeDcX7
AcrgI/VjcnWEokPi1j6QnKOoE0LuaMYNUH4JW7LENF1E8GEQv3Vu4pyxuh96uTBXTN7dL3pBbIjX
atxyrTw+O4r6+wevzb6qDCDabuKy5UxQkAlObg94geZhuuPNUECHj2KkOUWg5FW+HWtZPoX6Rs7o
ouKNcYv94y1lcgAzoE9me6LNZ04q1U5gtZY4RzawNET7aV2GK26hJHzmtTKUZg/2s3pOu4AkquVz
5qCc+vRnJrcnnyvyjj78jhNnd5jE8jpbOEzvQofBhgrrX8aU2rJye8j7t7xfS93pCU52AnbzrHiJ
H7rkp9yYmWqAdAm3n9oBte0VNNyAqn/Mi0q7XfV0foPPhcdCWReE2a3pPAqrZ0OdxrSMT2hJnSkT
ZyDIPyj5Zjd/2OI86rc5MT8hCEjAnkif0e0E+4xDOGlaPH0HBhKi4CsR0jpstiSHQP5nspaniqmY
l3lWZaaNUbqZ7+Zc6xNmTcSxrbh0CCDlMDaTIA3MGG4ppYsRbjxSUFMPvs6dhwIKyEWYFrg9jDXG
xp51XuWWWHF76Jyyf015B7BMppWyOoQMocQJz5hbwqf8G7YM6FZHmmwmJgsL683v0elPzQy1zCqD
5hUDmnMO/a+XXOXfqrABTXmuJKTdlqKjAdpouIQdLwPqBMSOccOCEwsxTk+zsneEENx471qc1Mgl
w6GcJaiTpcQltCUAAS2cf/5tfmnDQuEZhQC9RVLql8NpMY4eTv72TcXghVgW/vnhaxaI9vT874Pv
/k2Y8UaKJ2ojfSbuFpl9xWLypqPwDFKNnD/BlK9Hdo417mO/XArCrz9Ei6eRDo4It188thvxik0E
iMC+UOnA2U22a2yezyLF9lWLSBW8WkLeSyADDCXYLfZVgUugJYB3yKCR84hnXhw5ckl8HXg4Ak0I
t397RFicpskmI2rGLjZD9JYZkqwhNIL22ymkIplCbFedY+zKKd007qIwzKI9D13WMUpSPen5et7G
Kt7oAaoBs2KGPdZpEF4umwMiehun039fuMadoiM8fCQYwXX8C9WWYWycIM6kfphzvfnDid4/EXXJ
wgNW4Rp4bAYp7SvBt6fNlkQnlZMLtZ8q04yXt3BLp42AM9zrdwDUKS+Uzb7IpMmK2qr3yO45hFHa
3u1z8yxmmHhUJKZ8ODhS4mrBCSvejI8+juVAiKdSbjnuTokZr1YjKz0hD3pRbJGyKaK3eVkvuhrA
5QkiRBqBZ8VFRskrA/U472RWDKhvYgCmcCpaUlPGAtLgiQlFKqTW7LI94QpiG64AmdRvygwJ3CFJ
tStNhy5j1BYNe8ic7QXzoGqI2bs1mGYt98op0y5/zdse0Zy41hFP5nbApSBvFxI+FD03gvI3eGWr
yr+Inc/zNDuTJwy0LbEfqOxwWnOI0uhK1iwHwia68azVdLqYt0BBiFz8Bh7d6LWYhWwoobmZjLka
qRIfjhSzaf/rfqgtu4+vpppnSo02Vl1rQYASUC+WL/sn6aApGNDUpeonAs2JOl+5mRGvFVCrhOe+
4glsFzLfrBpfhi3F71Un/gE07EEGR8XWRt1WuwlitfGA/XR8fJTzlp8Eq3GcP7Z93zr4qFltg1ho
9dOkAeU52oNBtXei3gmHoS75Nls9U2xCu1Yxp6+9OrP7DrOnKFMHB2jDB9J+XElr9NipMXjxYbQN
+UUoEDRzD5tW1A6aHRMFmjTzZiINRxYfSLBoewI9YsQ4Isi/gMKywhRtOIcVZXWYxhRiAp0Vgomt
x4TqYciAnVY4vfasyTjyZoGBySbcLL9/dlBvBJw5CbgbjQtC78oQ37DskYFy8MwXiBp2mkNAvXuG
15pfSuPas/ADCnCewLdYpIP6nN3oxOgsH7suLc6yoJW8QWP3kpQ8YdFbAeOz7sDbtNwHx7B5reu7
z/Y2/tH6qIN9/PMeA4Le1FGwSC/FfFKziGTOfUutNbzlkeHNnjZlZM+rPDlU68TTLI1+lJrG/rOo
22SoTFhQM9m9hzc+5a86uSBO7Zup2doxqbBPL7Wg1dV+L3gSsIigCQ+MQL1TgHfONfUIl5eVQvyD
m7OHRamqEfKG5KqeFIvxnLXsq0Ucc+KUZCpQU4ZuX/JUYU9bMLzJFmghvUxOGjTZwiPNJN/CMx6S
Ebh0FfbU3CI/azk+E4g1t1ALKpoWUgNmwNfb6F9W8K/JnPnlqwyRQ2/4jZt+1VEJEvXJ6YZ6vkGZ
SUlXSyOFxxMyl+pwZDKWF/ge+X7ZYiWlgEsMqrYHy8F0IQSL93JpP2PWjgNxwBY8Bf+CP/4RyUbG
OrfvmSwFBPdoC+TM0UHmop/tV0N4T9SOEa/PKBvC4XLqDlwuDwtQh30cxomJAhQr8L4MhE72UkQT
QmuyxyuUEgoTn2zBtETftaNhiCM8UvszK8jHkGwHnxeOuWgLVpTCcNka8p1/zabavwlgLs9ueBRw
1RF24Lq7VBD7Yk4lRk/sYcTsiUeYltT0M5HEfB18abLJVUd1uzGmVf35QsSIh6pdGHmygaa13BHL
i6KnZq+kyu/VyrV3rCVvG3bcBgwt2D8RnIJSEw+eDAMlzIeLiQ4nvZQqHVi/ubJa+MYGJr7xVJGG
t1s4/NjIJtXVKCI7noSTH9x+CBLaYWPduNWwSGG++8dcWbyWOpmtyxRPEcONLU1kCHDnqhs7dPmp
EsvEAhXo8OZJdZ5Cij/cWxSIepYFuFSzKfqyQeLD71P5ziSkf7aJAh+xkMYKnB/wMKgxYmIk6A9R
hLZr0R9mhelAdp56C0XvQNTPRrSdvh4A0IEv+TnH9R3wnGCipVVZEYVXzRM+2IwQ2nlpzSkgAwiA
43oI7qdk7slB7W4ZaY7NOoZPrspO23MPgcnSnfc8LQeL1kud4MdaSIDOuo8Nx7sNvZbWuFpahyyY
Z9tYrsTX0tSiHAqgZ8syY1ya/pAgH6FMwiudq9PVyCFv29/hTWz/QENzqqNiVx/y3PgBp1Led1Ih
trZkhkPu5Bml5mG2xwPsS3v6mwjfNHRGrNSRsok27if1QQeO+632uRnc2Ic62OL3Y85dHE6XZyh6
wHUIMxDVOkg1BbGoeVZjexK1oGcPFDNwNdqNQozg3qDG+uOZhJ/lfIodqroqTL2ZekTK0xLfbe32
dSt2a+Olk3iDndpkvQvdqi+rhOv0CaQWuxGvomfYdtKY2g7siwtNORa3HK/yvTJv7gFIojPHhFsv
oR5LJJQa6uy3tt6am5BlcEO5eDYeIs+LuFBxEYJxAPCy5gOzbOPrbnPuUL+upS65VvVUtnFvfto2
ELYl20z0YN60/ML2MEoqF8g3bhLpDBXlB2sbH7eHtuRHiPsDxiwNQcflSXb1xnPF9EyRgjQl5ft0
iJxIR3rDZS751okAIftdRsubF0VbcZ1PJLHP4wqbQ7Xk3DQ3BpELv6Mx3ac87Qj3zQh1mJNcpIU8
NVhgTcYrVAagKjbcySVoyWatGCyEa/YiQVo/kQtwT8Jde4M4KRgqxFePCLKDrSj/c+UlFQUhqs0D
i0GV64F6O2C1iUC7ee8mhp/2672zbqAsPKU/v9FVe+KPPxAKUKzqs/cEM9sQ4HF5wTiYU8ir6Ti+
jeYgF7+5tu8fnn/fXFXeKwRIeYITC1Khf3BEA3nvW6Jzs1+PqSJgNQbYjt7JoSbpE/jieRKdSZKq
jroNhxNOp6A1BykuLiC2a8MAONd8pN25pmopNo6BwELf/wREckFtZudFlbbmL7amTI9nDN7rr+O+
yqHfeqPCBZzKPWWFr6bvZqDEPFnLG1ghkibVSlzQnWUIufLOYYMmH2TOEqww+m/qo9Cj1lIFU7F9
CkdhEZT8C+WrvGoLSRR+YBdXrPVQxi2E0t+pDAfGKt/Y9BRXwZC9zVzZ/R4qNG71mFjb2Or5uaon
OW62YMEaVgkh4ZDC31iRXm8O6xsOqwc6QbF04qsYT52ORZtdHCT9JlASIL3lNUqs2ZMexYmTfFXF
3qTCYCTlM6W7f/8vEURYf2QvL8/A7nwLf/NLaNl8YcbE/QyklE/TTMxuMR3lpPsOvVdKMdboqeU3
KgUB0PwtrHlSzVL8tql/MMWsCMAO5p/gLqfH3OtP3RjasdeNA2SGOQ7gLhwmgoygD8kDwCkpSMl3
Zth2hkytJDkPWrzwQ8K4DTlVqC4IivEL4ziKrXVb6wY7sfZcwxUYHUKbpo9OtMi/Jp1I47/clvAE
5mNYXw3HkZ7qGgu6El0zwKzaqrsjeNjwLBSW+YnQJCEFVUswzjiQ7h3EpZdcgDQ04UZskbmCSTEz
MmpP8KZoOc6c+4LLxozPA4i1UsCJ83xosDHZG2tFM494l8A1FX2ang0uuAnm/8/4ZkxMBpUXEbYK
eSILL+d95IxIuq90ocoqoKMdQhKfg4KfMsB1mCGX5PCaKuqG8x4LU7ek+O45YIkQfIr08efhfyC2
ccDvK5NYLjKywL3zhZ7UzjW9hu5SqwDPE+Kn7FNxzYtb7s2WwDnVDK9GHPxd1WC7l91ppsYVvSAD
hVeB63BfWSbOUe7JzzzRlNwHGZVuIIIDEYzjOLJ0ZLb6P3WQAGo3OtxRl0luGopOyYqY21t9bJm8
PDrY138aI0fsjpxpxcJ8jb10dEe51lRqSdTw1cRpGCl0TVpWL0wJL1Rsxw8iwwahHbnGrKk3mtFL
3ExFPLP5MdUiQVvt4hjoqsvJuO+hqW0BO4YlzzfYxevvd5aqLe6cRlhA7mOZfkvaOR4dac8/VhQF
re2EtvQH/bWWj2q2rTLJ4ym/tK92pasr269ogwQ4Ieq9plh0wUvXl5XIU5TAfmPcN33jIlg0+khs
k787ZVW1SlIvnZfTQGIQ/Pv2oqLzZyVGGVrJtEubOJB1c+egT5ve5ZS7pSHIVParhFEkv7m1irlx
Q8hHfq3yIkFUauIFd2Iigovw4Ucyr4reVpdAcp3vlzM6kv+lmbZDHt+0PqkO6pVc4/eU5T6935PF
4PiVwVkD9PeWHP82wNOPWlsF6lL0QrorH6ta8xLout2gA491GhD8H7OebHYN2cQ2fRGWfVW07fkK
2JiGZl47lItvHKqlyqQQHiMpJtmE2o99JceIiJdAxgAxxuNCl0uA5SNGoAIZYMSb9szdS5t7wwXw
Osw3sOYDY/c/oULwOdHTssmanDKWMrp0CAbCzCIop7v7UJWD43EDThrpNtGg4LQGcV9oajyG6cmq
QFvnosk+hY59VOLPjpisEs+fa72coUhRmGcwudZFrr57AtUIOEaMF9fnNmkRVdOHH1ujH3H00TGo
sEczzE4ytMXmpKGfdXPIO9wV6yOD32SOiIUMl4o6AuxVPHxTd9jQKiR3xRrHP4HbYJWE9+IkJ2Sl
KJFFHiPhXlRb4WZYoRBHZ8XpMpimfF3KXTrZMdIvt53EIg32sfDbd0hrOHpPMq3JwcvO8Tg8GOVS
lXEieWJKHgOO4h4rd03rMOdP2AKF3EzI1J0ijL6Z54Yy8+ukAngq6bQcjIjjMqSVFHz+7QITUJr7
5F9tKlkO9UIjEU7lg8sOifss0yvAi6fOQlBQqHJItLHmAV/zea1NqznBhsCUXXl+pKQdBD6NvXH9
eEPfC/pUkxXOBKQYRe+yKAZSSzSE7A6i/4RPptIUYEDczUXYCZw2VlTK022+P9Os1xA+KWLRcWUD
Mfw8vpWqELLQ2tcNidX97ZN7Sbeqv8QRGUn4u16pi4SZjZ/fibwAoAcA6yA5HYJkuYgzq6dU40RR
rAX2OV5a+dj1HCxoOHlMnhrgWmXbnk9JQTAAFzZc9t6Ek+VsMXN//T7zjcHiOWT0efuID9lDwzkm
vA3s3KRHUTn77hXIpf9zquoASCi+VMj5gnsHcvoiSBZbYOtmcVjvVPrjfb3mdNDJ/HGmh6RLu/G7
FrWwa19a3kQ8jED3rxbVxJVm/Beb/STpxsFU9xiYHs9Z5altVw0PokDd3ZYr7SXN5BZNu/ke4N+Y
nlEE5DiIO4DjsWczkuCR8rJWjpqR60en7UbgiI2MfqOq/j4B8bT9twU6Rf9o1/LG9nPmnUJbtxiz
V4DwBghNptcKrYiPkTvC1kpQ+CNw1tCY+X+ISuumScwnvJ60Oe76QHzOX6zsbeIuyIN7Hf39NJ/3
8+dlYkgZ3MnHqbO95bXCBsKr5UeLmik+MzrR2acssJJCLVGudGb4qdcwbv+9OHIoQaxP+RuBtHjK
xQcCbn02yruChv3x/+fuKi7LvOiJ+OOpRwgyInxP5MbnW9tpuybh3ftFewNeIoWxEYGqlOwVgv/H
Fq9ZkPnpU7wiKUxUy7wSgjtawK8c1hWpfJlrS4ZFg0RHkRL/pV8TeRB9eZJxluYYITGTw5ZS7S65
4re6EyWa26Ts4+CWS07TAbWbG/kbxTsBgfE7pEfrBS9Z5khOGgi3iwZ2dNLxOr43YNqolnFmtnSp
9uaagu1ttz6Ow32yIIvTzU1MV/9bgnwTEmgC9/wAqRiGyQ+UyIrNxtLolXFeIxzBPtZ89b1vtV2y
taVbJ6ZGRQvsVSPvr2PGL2VmaRssBt2eEfEhpBJRJbraXEAyWX0TYnnQjzr/uuxk2hMpOO78LoFb
bhaP84zGGa1WvPF4n8sFisB+lDC8CXdwnh6Bd3w6X+aU69TkGItdHaqc2MQ5sSCY0ebfnghggjBt
VzSh0N8WJfwBezObrJrjH4K7DBvaJoorEtSwytSo5ttdOzhKIfoZ5caMoNS06494siFo/KW3yOzK
juAwNzSpQfaVdCMYV9RSREdVJsQkuWqnzIuX3q0IEiJmio6wzn3JgEGVQ7TIeSqbolbyegEEQcUW
3ENahZfHNyMVlPb1dn+T4nVSAaB6ryPEOp0Q/MOonW9gqVwQcC2KaY5UxlWseOWOvHHSuB31iM3y
CoSJXRZEQXx5USqvh45ktvOAMMyqD/92VxJWxMTTpVYSgVkiOO24y1vpl7MOQB518Cf4mpvsLso8
rhJvVbmE1CqgGVN7GKN79vo1uhroWnSl5tuCSDjLwiqJ3KGaARbKFxZbhZf8/atRDaZaG2S9eSwY
o3ECRiQqjOzR6DYGMq2onThp2JFrt+uQnedHxiK3IwVMXNWmqrE5k1Yzo7Enr8fkYogOHlC50Qea
/JHcJnZhs+6JeFUIDDfpqqlKbKJ+hPeL5AeJHVUaaT97qwbDS8Uufc+VSyVJDpNk0ceZRJ+xOMwR
V70K1UHTmUDt6uX3UZK6DlxlUmkGZJ/R9Sn8z4BaJT1zl/v3EDaJELjx2iHUON5CJabpr7X+SCZe
wjV7lufhRURnvhLPm3Oa2i4cC99nBpIP53VcTG+w0iI61ihSDItWpE3/+iSsIKrGa8Z+Ta+1Y3kT
xliIDnktygmEzks+ouSwxQ5VVZZkYtA+iFF4bG+Z+OJ+6CJjyrICFYCgMtMio9F5My32RrMkmpip
yk/6qgKQUcHAgEHifBqwkF9l6TAAiKh57gkWeF/0ZtHj/clhRJrGXX6gIgq9pCAE+qog6jLOqdNs
15J48IKka5ACykRKmqC7r7zMEOCF+ReMOfWi5dgyDuGW1hFH/Gbje1ahScraPn2Yja6u+0yBnx9S
IhlCuYlcHUhMMHoejQ1jKp7WnBnxd6mvE5l46XGE2ZQswoAhWK0jSPK90A+GaaOiN59X0yLParJ1
A60voZIsH7NKygSISZ84P5u/LML28fEcwTwsMEUn9solo7ta1bYZy900LKLwmZLbdechrq5jF+aI
/cY7WVm7UE8CMuxIH/DFIWYydx4ZXut1FPaU206fnll0WP45MI8DDG75AxQFkUnIIYI4JsnZfb6r
+nUJhI1QzcqxCY7Y97VGfLsEdxSv/tEBMZsg3b/kE6Kz7QLN4sVFxwiXQac9/CJ4jdxSdUAWo3zA
/ACML+ZZXDyt9VCJCVzVqcvCXr05waxYXL6scFkPY8zHO3Hc5IpHjP665+oUDoiqKNNz83JHl6BN
3qdOYefv3xFE6I4SGn2siS0Ci5pwRJ82TDpUzUrg4iB/QuwMQ+usKnvguOXFN8CTT3QgZRinNKkF
BroYhMQpZrNL+v5TxC1yBCuHYKONH3tipwWh1s90hlAh/aeQpCAFplS40q4DbQu87YSVq9mT2r9Q
JLYZovtJ/K1hDNdQlZdNqM8BOxWgiKHgVPEI4JJoYNcmQnHVdHNp8x4HK8u/+TvZ1f5UyOni8J2p
CxSOmQg9GS+9gcykryhqNhl26iYCuL7PZDpVBfvIPUDX+Z4d/Bu7lbe5EAirpSCv69/1FYsot9UM
LB81+Gjp4/j1YAglBt+M4cF3hZkTUp5gWPzsNrpVBZ/hXR7Qy/z1vaCB9f/vSwyU6tXItc5oARw1
srR8VpJkjMkcV9bbfPMAbS1R1HTv71oBsFvgGPqeepvSeXW4lI255dR/kxmWRb7Vbotj783LDx4S
0lT2BL2im/LX/2B+lQUw9RXLHvWVYRbrj5Hpj+TUjw5szllNjXnZCcWEANVUMvd0m/OQU1ITe+vS
BaZpN51oss8D8G/rkCeP1/BCUtJeE9V2dAhKTV+mrgohDb/p+MhP+2Ks5wHpTY/AmNirREe9XpWH
dKoiBOdmRJ3brtihK1Dr7yNYtIrKllOsci3lOBW+EikkzIMtZtAJzGirgVVF/SqZTDUrjubnzrLB
TMIYG6cwo1SEEYF5b2Z5ICP/PAjicbYb0ZWqhc1Cu8VQRL3yankEwGp73wQiIwxHkh3SrP7yR6Bo
uH8Hdhw2A7e8qJA0xVkBm2T+ltDd1Kyiqt1gKrrZ+R9QJAE2EjAg4W/YnLaEMvixcQTl9TuLjRvp
6ZOAYqewkhp5xL4Zq3QchQM3/KzqZrqlAoeUrMhf5JB5YH2372SdFYR5XozQbLCS/WqkGTSPPHDg
Urdfln0bhJ4Bh/4qmpz6Me3oeI6Y1vYzjAvDXEUFQ3k3tRBPbnxIrhLQleu2g14qK4ZBIZgJnqMl
FnFffMdfHRxdcR79kGzoU8snhttVam4b4QraH6qSzSxzsq+Lvwbmh6f3M1dpmqc0Ei75dIgy0FAz
we3jU20AP26f3Pz/ZpeI3R3NLn0NqEDlLtlsWdOM5BmciBzs0Cy7kWt2p3enPjhWeOOXJZmCrlVw
zeF3l/F0y0wuSF1XtMRmVTJCUUbLq5L++m4/MtcmTZ/aHlbTRzQGcar/uewRSK6bxrZhcB5zFDR1
pGog1q/nxmGorC4BHH84kwoyPjSfMScqrMsIL6kTiqHNbw+GZPSOimQ1Lg3VVmNaHzaMU/6ZZm0+
56Mw4nGKmNB4VuAIiqrS4dH/0ft3oS8LwIXO9pEquNgM4RxEuGrSChx2hC+Y+RtbDJ/Z2VWbFfBi
CaIpcF8OX4E1UR2tDx/osTKsPi8bGXsCbtTeGMno+cYQzPPXtRkm2Va3DsCuS48SBGe9MSLB9zzN
zSuaqJtuXQPmQC7m80c2dUwVnYKoJ6TXW3O5mI7sKO3NusiIcouJ5o5ncwG5UzfhLyZ8iYQThPBh
7Is+lLamZjWys+g4m68csi8UNQBhHdq+2Pggq3i/ZQek/SudKT4KoqAt3LQslLqU/8huOPVceEiZ
L0sfLgnKdLslRRaQAFs7Dwkox81eYBcFEE7G2IykPEj/ruo5JRrtC9CJ1gWc6bnfHmfG4aux1W+x
BmuAsjS3lA2YIgW6XBEyTKjavraCYziyVS2F6bw8xhX/QgkoVJhUc1IS+E9PGZQAhh1ehBSLCSb6
xxM/t9OzjH1eC+2oU4WU8J1uechIfMq7XVpQO1tqqeV/gPhFCJNQnyiWx1K5YzChu7oRhLMhfJbo
VemcME+r70dm0XqqPjew88t3ZMGQCXr6AS+W9GgTER3Su8FdYoK0SrOlmzkrKhwZ9MYX8c6xo5Gp
jMHz8on1kjKu2IHE1FhcanaeIfGDb1tq0dAcFvbT3bopr+X3jc5H6xRsy6CZjIWfLQv91DNHZDvM
qN5YkyfNzhmhhUHblf7y2THyR2UKEbdtIu5GfW5MIPD4kHnqfzLI0McyJrdFZuBVI9u+KuidGBAd
3gGSKU1+vdm9ooxeJxIrErRDo6rqea5RrlklQVkXGl3sGD3auwPYf8gpsMjrWmcje3j0C1ReH1xt
CFySnDkEzAl+iRV2BFi9D9NCo3x9g1loTNfT2DYzRpytPa9dKyMqCGDE6TiOhYCWB7dDsH4jQgxX
kHpBJSUnUABEuJWExn99XzHHjmH13Ms5/IHjVgOLF6M/ld8Nr/4We9TdSbUpUhbUud/3MOvrxrTT
l4xeOdzmFt8YlMBNoq0wPAWu5P8KHoydskk6FhN+44ixKrR9kISd1Y+XpIT6B9iNyQpU0YOKkaN1
fch8JzlIyi+ksvfjQjd0gscc1G5T34lZvT6sVfICaJkTsMhq6TJF64ll5mnwhvWKIehze+D6wPEE
uBjpmfzxwZQ8cGmdKBxtcXmypHnCue0Tt0Km8NlLy452U1UZ3FB2cXE7TRHp16Sdgu7iuB/oiIkm
g4fkUFdcBE2G8Por706TnlF3baB5pfELvnORPhRXrXQrFMT9qwQhSLgx9svSEan5afvq0HkIIedJ
gOHN9xOU5KMvmTcZ+YgwYF9HWJlwVSvspFRG144ONEPLUMBzQX2LMcwzn/kO0YT6TTBLsg6jIZF6
Xi/xTvsJ54tqvJXoBm72MVmXueK7tpKaVGYIxRwbR6K6m16cLh7JGj4wAIM9d2ykjHih8DCAEMbY
EC1p1N2ooyn+LURrJJxWJ9VW06689k0ljcezrBEt64TkRR8k1MsfcETBsBXOK6A36+GME/ID97KB
cc3iQx3jWr/NAkx7mmA59gEqlHd6r8mWmrzVJzcK6q3RAz39w5tZbQcU+MtUr1O86xpLW1459yvY
Zpro9nJ9t0LSiqeuO8xnWQzi26wn6ZUfgNltq/29MvMRAE6Du3NcHl4lMegdWtmSsG6So3KArq86
JWodhJoQ8LCBD1w5q97z6lFrxh9dHsh9/yKz7jZ3OeDolYAgQ024It2r/xIqZx4QRJgHrnsnjF90
NIVzeMyHejWKFWdz+tooer7pT6C0yEe/v/JiQrvvu3Fal+hhABlSMQIw9i024j7AyI4ksMZxp2T/
ZwEX/1yFUFvfM8gbqIblH1LXV8yJZFn5StHOmEA4Kr9E2bXGLxTuKCiapo0muyX2pCXOX0XX7jgJ
RVhTFqBjfWOR4qcK+ANpNYCIlUt/Kngkzq+/TmdjdDtP9/3hW6CR1EpQi1A2l/7Yp1wKT8v2BbIK
Q7BIlvNGpUfa95cxZwY9UrhdyHB1Cg6Bi3C7B8XEnn+nb2ihPbI+1epsHjOLpAYBOW7T/IBHAjFR
4HzcJ/pwnCvMs3xOefyWet4ab3dq+27VNtyqr8SVliWGoCFOQTpsK17K8WgTq2UhFg5mrvy6uoho
I1iRwiqeOThhX4opTzc07ToAzf6Gsc14f/Er0hdE43NGiJ/yzD+GN1mPf/qHjxwFk9OFDh6MFTxv
75SdEo0tl4GqEZKVK1FoZGXpCpGEw2439nzYnNhjVOR5RVCYEbgOGl7+EJ9F35rHGG9EuByafzSH
W6yXIVCXETV+HCtIYX8XldBwHkCggg/oWZ1/wM7TxvGJO4PdriTrhNmdrprPDKBh+BXJsQR1SH/m
tEJ4jIa3JfHkzl4FHvPNjQKENkHYMQWujkDYLj1pS7ctuW+yHTSxVq51sID6sckGyJyyy3ud8S+3
UIboKdb0Ex1LJsuy1Mv78CawMTdMiO7qtccsJKpQTehjttIeAknZMjtXUXREVAuhvivMwwkfTh3E
DYNpQ5gU8zeRBfiA2cD6UwDY042sO6vpFO3q16PSd7wIlh4E+0k/31ydGk4/do6L5sYdheHoVAYD
04FUC81LQHGKJZK1MK4DpP1sWski70ScVQSXX0fSpcKZDWsXExDjdIRw8Ol5oepe7G2Pdr+rv7F+
Ad2n//007CEbV4t4TwCeB0iQSDk+oIkYDSo8jvtUEvLPQFCMKnCo3j4aKAKTCx6d9ARDa5i2L/g9
JSZggD9FdYZm1htALYgd14AwMBoy089S9mpYvJwluo0iZXycSR45TXDNxDCcaCmU1g+mb/AfRX+l
5aWpy/gKMN0VnzDfSmorLnpEAQWG57nO5+fsVVThEMWVNbMagYsLO2n/qh2rTMpJ7kmzmeqWTq2L
uFtBsqCYqBB3OEy87TgC1rctJ6Cby0sfmVg1QIxkgc+XHcfCLCOcp1BOsABIFiz/M5ID8DUyaW16
m2Xa0xniBfOMEG/keUDloDPENeOMXnzTgfb0iPI7Y35DNc2tAub6X4zzoYSndkB3iICK6V6lL9LK
pNH0uX6XxQbzdMQVBPpDT65yFkV8tB0/9dHtRPWh7wk7dKjV4We/ghXm2boKzLQmyos6PE+HzyJS
PFpZh0yAOSagabGycs+gG4/VTcIVFN0dk9OHIz52ozrbxdTvPnzxDoPbH45gRnN34MO4VvXPqlse
Sk34mLgH4KXoiHB44DUhC9iNUXWgzdX1TGX33LaqGn5vnN+87Yv6XffMu0io1WaT2iNuu3Smmwr0
KelRc5CSesDI5zhwTnbYIaRMHn98OVTJuryt/Hg5vZolmiVF1JYEFb4mj+hrGzUDZGDGn7PFUUNE
DeX26dSF3iZFDrjSCU56pT1HkxKPy4ZW0Z8TU3cK2FWhoN313gZzePGRo489rPUls4Mk8hX2A60f
j0hfCMy06Vx3nmgc4bJUkpAuu4ylHXFUG+Bzu/atMTH6ZN7jv9ll1XVh/KP3P/1juFR+zQI4GKjl
smgqciP52Rwdr2bp9+dTyvqNh7yqjcoMdz1uvyjvQ9Rpl5GKHBV79nUL5WAVuet5AiE3grgKCwDa
NnjShu+26aX3GhfxG1TVtEq30AQODZhLXstvTyOsXR170QxfTYeiowJNcbxaxxnPRXW4PI5M1Avx
eeXKmN0FoWdr/50b6zjtkmigeN9ezbNGD1+JFJk1LM0V8mNG0C4XSpmwqG63fERXX+hYXgx7+5WM
I1/mQ88nuGf6lks1ZCn2B8/jIyLsz5X12vNj6b9mvuKtZLKJilwM63ajSXMEYt9TWovoPeNWqdzW
Y6yodFsFqoOvOO6gzIOGTMVHL98AQQZ5lJfaYzzMjtWnfREDdIFruQQA4LUBDyOtJwLgyJAbW/td
sfk9h0PjF1kYQGSLt8/V4E8ghzVRai0ftWRUNc3oz7+X/+0qtAOk6+ysu4NKj/FtUthm1FEf407I
V3SiF0ZAaZSFEYXUt8/oECKmZma2iGWfcxPTScYjeN+MR5Arayvcogb8QlqCYXiHpAhfGzyQxirI
NLdpZVe6R+PMFoDm9XrYJ9NqcMImfzbqX69GLKvq1X1/FbYa6ke7y2L1X4MXPpgbMp17jIIjz8fd
O8B7FR1mDb4WaXV3fkZM1nTrcxwRtySybEFVH9TNYYONHaIRM/0uVKd3KSKzRDlkEgZFFoFR3csD
1z3xdpjKDQxettaEj1tXnSLKBA7R3fTm8zSnZ1Nf+se56H9iGNLP6O+iZofKjP6P0eDHtRj/ZQF/
egdv55KcVj2J2QVo3xb35qMtl9L1XZPSYoRVCsxs2bRTBInqcNrRSQhEpRzlT0pV8h7sieiHa9Tb
ysFfa9p9KjdY46dYg2Jcwt2vTYOHDvCxOio8eUmIYXaHTtBCLh3ahBA7zxInal25OVUk4spcGstT
c67/sTrNiSwx01K+iyGWA9Mz60nxRkvMN/w5+44C3+uGoWXfRK6sV57O1LNevokAJ3ldOQm82Vbx
U3dC/C3FF02I9xWE4vOvZyCgmtN24v3L2uPtdtuXtzGSEuH6tOo1c33J4AxnYKV7mdbyB1PqnAgy
3UBe+vwXeYcsnCIjb5kuwGtvx7aBkk5oTxYo715DZ2ToRRXjRM+aEL/fRkkejlCpyhBt1ka9SKYf
Vk3AUEOQjCCkDWGHRoD6bEVRO3M9erMSvR5V7dz3mKnZWe1pHe5uw31X8NZ+0xV57xMeWstNtojZ
i7WRwnAmNbLeJEsfz5y4A94AsLv8S5lMbCMEbcwtka6VcpLuttBhD3FCd8T+R57Kvgp6KEDCSff7
051EdkSISnSeW6RDsmYAWhqMmqgb6BxFvslsQSyUe1jR7YJHJxqfQa2dH8XK4phNYZf6vO1fVkDx
kKfdqTxE6T8Jl0BB0124XY3+0GDba+ZOGwZvBNXW6FgjbovPTF5Wp1kCbggHplK8NDF2tYRIvQLl
Zq7pcSIKYj3Uhj/SsUNDYh+gNswopEVbq0H4OfvK7N7WI9hY80dswbLKxHfPHHwkuyN3jK/1CcsP
a8+efVjIilTYf8FWE1o1Cy1+kx4TBbUsOSWOB/InlJKlxVMTc7iH0qjxRsTV2Qz+OeTUaR8NTSW4
coW4Q3khjskSyQaMJjdCSUeCDiGPImww4LloepilaumtPKxlFLkGqLqkxyAc3RXcT2/+UxnrsBER
4c/4ayG6O9wJlB0n04lCD/svgAe2IWnQUICAKmwXUdNsIUpi2f3e0Yr0agN1fB0AAPWHYrEA2lVM
jzHzVwDnQirblD3RcYVum5UIzH8kQ1q5N3+LjrNfj5XjMWiEG6gP07rJAz4PnCGI3rY9YTi+qHfY
gp13hQL+fbffnjDMfOE/tjzfhnnh33rzqn8wR+yOKJXyR+MO3yyN05Nyd99ZVv/889kmsWptorQ2
9h8UbKGnahyfiMh//KOCItBA8axNdUXtWS3/kx2560hnwoD+1wRr1fUamYFuZSpOublPHklqp/Ca
LA61jfnM2PigTSR86nzv0Qsqt7u4FExemra6CNp6JAKujJDZe+PWbf5z7QNhxZO1jvNXavZnJO8+
fHCsPjZlYUNvoA+ZlnRHnAVnyJAAyVLa2oOajV3kvU8U5GGnoX0PBQznpwfjIx0TZ4GWZr5OGqw0
rJnq9/gj+un7L99RpNRY4N0glZ+oxrLDsQEKn50nIVQeGVHemCeyng3dsVhmFVyI4LG/zTzg+AXe
oDqmJjNknpiXG0thJI3UlZ/o21WLLXuW/dugLXD7QF6zfZXOTogn21ZkWcH76T5yaxRQXS5PYhpN
9fvSU/uKRBVcg1CUV9JgFZ4nnTI6fjbzBhMiMnn5bE0JbmqX1H3X9dQUJY0kp9gDAxCBs8dCv3/3
R+3xwZT3r3sWq/Gne7blJ/jSIv/erhsgI9WbM6/4k2Nd680kTFNRevLVBQvsPLaoXMVGGeJYOWPq
1EhXYnOvs9iqp+cVWsfN/xo1b8bvR/5LDrp7MJwhnGOCV8/h1VQlBuadf9QPR0mXNQezZ4grYWwF
u4whzfT9Ux0J6emSGvD9naPhwb0LVvQKmfKJiaU7GgC0gCQsDXDUa3liJK78lxChNZUyO5/PKtk+
Qmgdu6v+XXCLcxE5P6eC4PclkAa5ndyGHoMZ0j8YqUzoZGwOE3HyB9+/sccpKK+bRlX2OY2gSPik
Eouqio05mkuJ2Eaj6pGDPDzdNe6FNoK2KohBxiZQ+VUSKZbEgdM5XjAWDv7Iej53pjgGk7InlShG
MwPE8UZYz+Wjc36ozeh43C3xp1jQdSESLmlREPwQicaR8a2VU84xvPI64tEtA8jGwY77/BGrEFhX
llbF2JvcSjCKfpuoNdTCPxKBA6Cq5s2IWByHXvjUgPRwPbGhWLv0OozACjy8IFsfM3XTRPaZYQKU
25vCVt1ZM03Hmzwfr686yT8saE40G9IqHZWaJivF96+DUvicdpqRlh8XCQlVTD2DyTxwRj73QsBn
gKp3BzcZex2J02JCw0q0OY5EvJLIfXiHmixy5tej4Rj4IR3+OLLYU/oAO2+elM9YIIewbjr1gnyj
8RFOH5xMaHI9SqYCFRkppWFBIrh0pie3r2R9YltH1iv7iaDXaDLk9yRIdub4apReJkTS8lb1pXdJ
UDAyfSdn6H+fQMwxeitRBMsYV8OfDH7f8jbUmHZ544zMH82d+iS+d8ICeeIde29KJjGneW8vUs1a
bz3lJ/OA1k9VkDsYB0kAbTiavaVrwpgqGwbrNBvwb3W+HNpJHdC36ocDiyNKMMXg0esqiUuUSMbf
gjgvJGNU/ESm1Zled2uG8s/R61FqGH9BGj1B8pl9BdN0nLeMA9mFgGfjorBtt6Hu3G/O/wJFCRJG
UlnNRT3H5/zOdymIujrvQrsbzXYt/lU+I1OV4mjUsNtOFrw3nWUJ+08KRCRdhiBya7seKaXVN1cc
Afg0qIsowV0Lh+wv+LMOd095DBFR8oIYR8P3Kw0wU5rdFyV3QfYNB+uSNgv3aPiiSnuyR2ybfOKj
tNVDsXQCt7xDeg9mJyhaTN8vxC2munjl8sV/xeyO9YPeakRO1HDPm+Yk4bZ64doZVDtKaAtmDtSN
J4He24AcbRR39o2y9Uvt0rWXqiGX7I9ibn4ArQvGW9Qjeygfaz1gnn+DFMcLrU5kf7PM0bRiRYs3
B8QSr67LZixwcRCqziS5/GcZEHJpxoyKt63RluoSrrw4H2jBpwVgRkcU2uq5ZdD7ijatsEcOVw4o
wMSqoaXQbTvgR/oHok0cJTRFDbXkYcd0QJan9kyVh+7sqUDmeAb1L+Ge6JUaLw3l6y6rF32AyVVq
k1rJTK15jmxg854HXqO95TjtAOvqG4ic3/34BLSuIMmuKuwp0Hh8DQcjgkSslK52tCHxoM6Snjx8
LyccwMNENH1fuD8R4coV3Pv5yJkJzlvJQfQB0q3TPPqmkEY9Cq8/mef21/bwHVt7QtnQsxM6iXJw
uDbPaiJg3MFjTTCBwYP/6MWkTdZAKamNMkyS91GOsId80JpGY8hJ4brr+TJVHSvRSQQm9C9THXec
jUL9ZCwx9aa5VwPzZ8G7qrWJMQrReJnR6OOGEsWTp7MCTIDJusCgWX6jqO6LXflt9BPsTrvqQ12y
cnxary6Wjjd85P3MSH0aM/Kezzu9jacbsI49fkU5DSRT7S9jDqBrJOFrdqR7O6dVIajG4Q1tlweP
oK+P4Gnt9ciA39VzFy54wvI8VeqlmCCX+CfMwr7xOJF0moRwmwB4yxSQB8Yt7MVrLSUGqQQL+sTa
ZpAAAmm0+JJ8A+qernKlIDWL6HTcU+SrY+9grVabs5SUkJgTwIqcbGXgWpETtK7xkPnGSFN49F/j
1iWtHC9X154UZeAf9tnBk8xKeR25cdkYcfA1oLFtH1F/VvgxRv3Dq53k2qRTA1JwWh+uBomdXs+h
aN5IbhlRYLFRGu2jcHNgZ3vX0sH1TtTFyMYj/Gb1nPH9ik1E9xH23Loo9akNycKOwwHZGu8BaQoF
XBAPLw7TIrtJt6+Tz9TW5oYoVPjpfzkhAmUERLpU6Fq2XtkhTx1nQVgd7YtFqlDxD764+smO0L2g
F6dJr5sGt/CgvgVI9h0boI6CgqW+j7qpgY2wJqb9SmNyAQ3K0xeVIFM5ZysHOZS9ovAPLtqTTI53
E4OtvidHQpF1tKJYzqJBEMoaN3dEqfSPKrVFegO60D8iVhfH51biW3SbwuyEwDrSY7R9XNvwsnAh
WcNCE7OS0cE//35E2Vvup6bbgp3k/ml2yqdbA5RpxPU8BE6TVmFu0qKw8pPnZyqY7fW6t39DspLP
cWosQ6C9KMowac9nFPblPFE02KZ1IFav739lBGdUvPM2sKOeXiB5nL8p/AzmwLH4L6ywx0Bjmlk+
JF2Lcbb1FY7co0mEfopq2J30vwTmYhC3LG5wcfyTCHgil2gVHTSbbyIvtocQiXVYW+hLQxve+uok
Eb4QDQ4ODzT2T4oT25SAcbmudQQQ9aWd7wlOOpejklIvum40w4kfEeL07BWWEHHW4KZs7+e43qcs
El/jguEO8wjc/DV2LpLvrw/HLQUP6mLS7kM4kXsG9JzcEQZdVjpCydtzx2LN0LCH9ljNrQ+pa3FH
vAe4ntJxjyuQe7+92Qnv3zg9zORCrBQmxU2sRTLiWeE4LO/PB0ATPHdcJYnW3+8SFULHO+TUOHGW
R+T/XbQk0mlsfGldx9zZfDdxSpXxPewAHVhyMROizXgUn0+QOjRngYZRqcBYXLWPC/7Z0B+UoCw1
5JY9HpF1pFDFCn8lapTkwJph9ZZmZMQkWnLlvTKY5ScOHQgZaGoM9eW4RglWhrd3tWF/lYgD0gOe
+OWTQPUzJTakXuga5pTLQrF2K8F1Nh9ojjwueQp0bBqfdXgcSp9ZvmwxyIsE2eVBQenndsURR8gv
jeBKu9pW5VYBiQ+b2zD9/xah6hJcqGtdgIlNa2uD/yAtZk1eVuLyx9K437VDloSSytVd3TXveMd8
X5Q5t9RKsziR8GE/s0Gd8nz8nkUJqMC1K/JohLOGRDyF3ThS+LathUSgbs4AoihIygNLIljJ6elp
VJLjMeaOgjkg4bdcFrZgabBp5A4nvHLAV4B/dBylS1QvitkrlBQkpOWVEr4LFWGj91zNOTR7MZFv
unEdPW0IuyB6ckqn7yxRSRQo0qr75HhJdjod66DS3xw5Qcn+RrtEIUMEnEJz803g1YH28CgdQrq/
ocA1l5ycBZE0nn9JTexQ6Ecf10kOK4/gOWUd+ac3MyxQz4cdunI4n80jqILxJcsNaOLVNzOW4tLX
eFKuy9izGUA+1BxmtFW4Bwunmb89pELQ6xc78DbY6Ouih1lrEnApu4ahM7BU+cXHGZB9ucPJYntI
gK+6ZIsvn/QMnGvTTdsDDDSPtr8G5eBfCCx9JdfZvHr8+ms0f+LyRv+IDqw56r6TTTwyMnreJWJk
vOQc8bsaTk1lvX20UDSpI3tRdXSspUU1vegnSVUdwd6mxpqeMyXFHvispkHYyBEB/NAFa+icigN8
1X5z6IskoMHr59+41e0JOB7B4bIfz1yoj5/W5FR0gScJaXrhgcpkraokf4tS0E4kZUoCLai2s//2
xkyXjmCg8erS1jX76qfdFwHmtTwwOzxXzHz8/Y03o/2xvM3ClfCrKks9Hro/E7Lj6v6sho/29il8
h971vyDdlTzgKOv0y4sYmFI1Q82PvZDWMQdjAjZyJQa6wYzdmm6mtpV3tVdJulXlI+dDfI/i64Qt
SxQkTk1xaFbmBu78dVdhuX/HJfkt1zzebWn/BCaVoB7XQITsbqMqLv7Rv9ZTOSekjs5dVh6Ldor/
tKri3+7TcaBmwyQMNiaK7qaQP3515rblWKG/SFEqkSPQ4TwXbodLwc4VK/qFJiICLvJCXFE7657O
5VR1oXmYUWsHDMOY8c6blDX1sF1y6rOY8dlitxRIHxYHrgwUZKA4N3A2g2wfFdTIbkUeAn82qpcb
TQ/PU+IerwBoue2g3vlTn0hK5lRamln7uYqnWJqixpBNWy/Yq2Yw37QZwJyuqN2V8Sx8lZ25cD0p
mxo291GLrWyFjuqd6J8HqdoQ6pp9oqNb/3Kp5mb4b1JzhT7zCktM7ksZr1ysqKWeQvXawIBydiqO
ivIETNE7szVQqmNIWYthdMlkKf+aKFx7555bBgn6VYpAB2Dhgioky5RbvRFiIWh33zYQtUQfAYei
sYpPKeZbqUUqFe3slhGlOlfWPkrjmqY8GqJPommoxxvc6Xsa1mLQDkgV5mcsjD6rO10uwjstlFPa
yEErax5UFeeDZ2ETV9QnNRE7/duEAXNEdbc6q0Pqo8esaXfrG+tlnq9GF3qtGnyTyyPOtHXf7vtd
LmaOzYsQ19o5cGL/rjKJ+vY86zHDJR7B52Cpty/c1tjXCeEL3rfE57H30+N+NQnU3mXY8Y4LLMpU
bMO0jvPsZn123CajS40RRhXjX4UnWmpypX6qAIjOTE0wLHlYV+X9qfJM3+oCUXuYcXoiD1kk5xfH
amL55AZDcVsC2TBzjcUKAm99wXgq+Rxa/T2w3QMZRE3VtNQPQgANuXLXJ38DaQ1VZG7vYBGbeoGW
JgV6/6QPu8v5fk61Ru0WsbZ/5SD0TopfPw55ngsbZ+eHdifWb5AhG662Y0reIsQV/w8sXTf4N/KC
/TNIopusucMq7xrFIZHBXRf/2JbsBVyQWHP6aZEvBWnEbwi4cYKFe4acmr2kRynL/IdYo8yfkj68
9ioX79OQtHXf07iZIl4ywQqpFO5MRSLwR9Le5ZSHw9/IkssaOYEASQvfgJD2NYvC8phN/GwULbK6
VpYeEYL2SjXB+ZytYsD+y7JDBbWtbUEQclnZph4AuNJvBbjkq5ZmQx7A++0adr73niP1QI5kpnfj
Tqq7sdsolUq5jSvrGMotoDfRcJ9TcbyPbHJ2RoVEIm8doU4oiawBXhnoW4tkoYOA950yL8Bqcbs2
p8Mytqgo4GLuqrKN+EF2Cl9PX7bq6SxTpFKYvV0sRTZGLOu+R9PHmJ2nh/V/UrH2BXKnR5LTLT6P
sKsJ07j5HiRkzd334QqgFojcixMd/RxdPWpL4i/xkY0OFIzUt9HsK8ydku20UeRgQJJE81CXpZJr
MXTb8Ukgq2W7wEqrPvtCIDeGnNeqtw8Gpg0prRwU/E+N/FZmnGYprxscNr8Nm+xOL+4qekSNMMSw
QALfHYrZipDdHKI6Sd1tOmCc0a9BZG/m/N/oBWEYJK9MaadNJhkGLEg76g/CynJhr9Fb7AZgmdOD
Tii0MePqgNiK2di3s1Z2JXYZqXjvFEUF3UHE/TVzKA5Zzfz/pEBiARvG457yow0u2/rEm0xdEDwW
xXdvNVlI8mxMgFE+sykjXPdunmyQVOQKUnlo3/8F+hqfvjKGRFShdJ+usenjVchNs20nLMixtSCo
zcla4Q+70X1N7kGoPTBI+DjZeqWEpjXtMM5jP6aAA9sNoP30Gu7AsDrMQDJCjyTQNLRxsCRxRhd0
pJPnE/MzfTN1qkx04aPHAxKieQh2lF+ZjcZnqb9svFC4Pri9mcypl661J5Rom6CD/SGkmhdXoggi
vJVN2SM7tnjo2soUrBiBhN1QukZ2z26cKARV/9m0eDPw+Vevcr+LHkVB6Yr919miPrFnOZqPPNAQ
KVMq3ouuyTQMm/OmUEn1BsQcLfG8+EbJ29LlrcBmTgBcX1cESIj785ZSCdiRrTQWyUsxscp/JD2U
T5tWlPFggRHVctgu0+U6xDqJlNpay6x212vjMK0I1jB1jjGS7nCGvU3TLLCGqqLBZBplnxPgXpZ6
kyv7CCTWj3ntzSnS2jhV/udyYAb+cXHs84ROHC/tPDW4R7pjvTTfblWTQ072wc7p9606iU7+DKEx
W2CL+96VPBUG1It1U1RZgSbdeUboM57IVTlv9Cl45oQ2RlRP5bxzeY9M5JUBvww+5cNpuMiP7GUS
ExG0cSHkQo9vjU0kkqO5Km+tGIt7hSjYHCs3caJDf+cpRBvA9evBzPA4kf/3F1Px4jWiVsZg9ZPY
qSo5caEaFIrUIK1cP4RVbVQzK+KPfkdioBaAFLz7LX/jAMFLk8Oc+qozcxaZ+iC1yTrBj3D6DZyp
vPVulYbnW8yopATpmg8ChpMPlZ1r6LhxwBp5pr/ZYZ8IgOf7tZjWApGWt+td6QyIfFNJP9bACW3C
shmu5ygJKil8ZaznXTZXnDk1tBW3hZ4FjbnhmJQud8ddkH+WC2kVogZdbbx9Ru9M6ugB1YGIUJfA
UEkLE2NmTJ2UHT9m6VFBjUucxOtft3Tb+1AqipOziWpOdxci6tcvAguMrjxf2ziH/hf9CWuFd+e5
zcUCYVJO406CeqW+S1yzR0ItHxun1V+S7hCfyr2x8UGjhEJdbQTsj7edTA/Mq7vonV8E/BCOUtGc
kp5L2MuEZNruxmC66aYqmufAdUvexC018JSCFEHEtZeUXb2VmHPsfoKO8ah7APzOfgk2HvFbfesj
3cpDlut8l5pV5oi2gITZsPkQ+we8TYDfw9bXq7b2TDjGZOt6OfOet/Pok5vE/7xyeOaVD487qHnF
awvITjt5KciZmLBo4HnksODnu8tJfCienBEEmxyeYISgT1c/h5Cxn67Le9oo5bKA9xVL+e9GWHY8
1j0bHxV3HZRZDYqy+8+Lxbuxhhd0QxfzTGGEbT3FyjDE/GoevEH6P2Z+ieM57LHY12ByDCSaRAPx
Gm7/fSJtmrTC8LPe6hNE9D4qPCB9/dLZb+TbsEiE4l+i+/YLZv0KbCBAFuicDDfhKBH36cLL+6zs
wEQMqSwAH6KC7lVbB29GaKox/L6jR3r0y3Fw2RPkerRptQUT7Xc1/fcn/EqruGw5NvGhLkPK/xXY
wQTnqu/7d4hEkq+ukxdxIOgPFbcguM8MJBu3tQQStVc/gVjF/Bga/9lMpodWyfNCHNZ46XErJX5m
cRcW3tUtZukYFkdhDga7ohZZW23Y+W9rmp8oiMWQqecgFhhym2dGA1ZsO/xoroB7bi5PqC0gCS/f
Oeo+zxAhTPzhFSs1DAeJpIjGqr2bvg5UR2vNdI9RT53koyMaoyZh992qVLZRf30F1eBCuexaa003
IvJeXKf5z4AWfxjBbttsa0Y2YrcB3FtY2JmNHT3OOOpvgGTjcZrZRVg55NcwezLV+pbTDjO+6G6/
jbSYc/IdMVndIRhwJOb0vE4qdesy1xY2MB+VnztPVkTKnKIgfbJjO2AXyWQhfIKsfwUjiwKPW3HG
W2x5+FnsjKHEVoq1PU9ve1/is0XowGngo/EqtnZAm7GxQlZdXI5Vg38qgKcWUzFn1CtTbLV+UtGE
9szjGPPzUWH0Bi0bZWadJyNL48SIcuX2SWpA+x6S6/wmcWW1aCynjTTni7gNP+cHmSlDqOIpjBrg
16uPvpDXVZd6wKGOku5X4qaL3K9entxCpim2uOmsONBrgqaV4WCVuaPxStx364ZpLzcQh6fUR9X7
REY4OaoiUZ3kPjf8QHUr4aBcnOdnmmn9cUSphCkI6KyIGrgeLwrdbNT+rhgKldwWYwEBr3hxZDON
I6DdzkI9Y5vFar0JC3gPjuFFPMwZPJnKiquRnIUg1J0bBeeho4UXQVtoYNPR+tLUIuoZQKDDNwOB
qjhe4NrBMU/fsGt44zAyOYbz6f4I4mgwrPE+tO5Y8+jAsgHnenSHqmv0VS5WiT0wKU0uh5TcOy9c
HaqE5HBP80DkSovwdj8L3y6nfg69jg/n5IQ3tjDfOXbOh97hvy6DPAvbDh2NHiGr0mQnNl7WPv1D
z0K90Wxu0xzzPMJnPRF/D9OIWlmlBX8mvd2qROw5UkDXHV7/DLDaG+XQsIY7S2K31ioY3UM9xcw4
y++c2s2g3bDMH1eUSnuduFrJ8yLGU3+jaMvMVOYaV7U4Wed1qJaRGShsU/+Bs0dMoL5ue/cJbX40
iqObAV1Ziw76+2OhyQ6sgGe3ss0KWHRYA01C5TYuNi25fwc/LQDUTAyNdohVGAal2qWDxS++nq+K
Zsqp9sKzOJHcOUhwhABlg1vRu0qQfLVXlub5WC3YBpYEEx91CogmPNPxMbYn+/nO7XMQUntDX/vj
OUuJOYvnk/T63xpaXKjgLyalFzWrmcMmSnXpHhlC5WBVug9uPI21WodzXLjifmOnSH0xo5czGxRc
PVmCq4mINnYYKtVh2EfRW2KxkO4cgqhfOSGKJr2ZM031qfbrmNlow+nMwtEzP75RvsB1fqltG/Ae
dlANcRLYq3NAC0CeNdTRWNaoKD368BDXz8jAnBlKx/ZGnii+d3HTCKAUGKg3MTquU1GPGvbPgufk
P+mfdnosWI2pPQCkDih4VxM8DMsRP3aEX4EtQcCkyNnra37pHTRgY1nmMjmLVeXuITivB+C05NcO
fRp6q8mzwSTuaO5bt/BFyfu+VIAoNJ2Yhc7fi/VyDkZnCh7uDVwbYUWitBNi6MeAMCfLgvpZXWC0
0Nn2DiqJl1Cwl9NJ/8cnJN4Wudykfqsz7nueodIb0nncvyriYPcTj4sGhjhImg6xR1qLF7dZ4fYF
wXUVuUXlrlU1UrNegdCuvA4MmnkFqgh0CIssxPdoY9mG5wCpzeO5RCiE4kD3Dxe7bByY1j1OLlqZ
4aNHWwmfgsXBVG56THJkcvNohMp9zPVHcscOXSuT0PrRa2PDeNFf2Up1/NWvSUoBnn25Hda8umiL
/XBgHbbHwpesnZhoHvIgAulQXXHS8px2gzUF8bsC1Pnycdxm3SAEQTBSP/pPl3PCygHgwX0hPZ1k
wZhNMj2gcZ1I1ufRvVIwhp8CjxIZiE9036AMvf8WDDCwJsS9749FgoH/JitjnG4BQgxcag4gwh9Z
vyf677Mf4NTnbVNTYYznPIwAKGwy8M4LB58LH9IksHmn1Xg42MAs5wm+h0Ee/JmR6mrOIlAaQa50
5B+yzl7RHh8LUcUt7xSiigkto6EHiyF7bhIdBXGXvikj36ZNVnhQPxgswXbPsHskZPkcc7N9swdr
uch5rQMhbvAz5vAq30RozVsNCK8LfN5kHvAOHxHEDD96/fSRZ0Ooj0q7r2s9Ky8w+X/2udXybZCR
AyxwqEvgtB0fw+ciOE41Z/LvU2sJHlrCDoq/UqCfV1IkAr1AGXKYwk+FsDCKclCP+vb9j1a02k50
JkD55yiKJfcUBqSggKsz2fnMErditLQJdw5ABo1JufSLtszTaBbjEWe77woEOi1ubGX3I9f9pEdq
bu0/P89oXiC14bjmo92AGsgqLDZvyS2bgghnjmdA8RYQDhf10wrtWNw8HXCALadc38Epjf33UOjk
KQMu3gC7P6wQFBU6iwo6pc18q5dAOsAPI6/jgjtNdsubGnByZYxxxeKHoWU0paVtM2ybLMU6WPNt
GFHN9SRJrq6V++ckmIwREy8OGIPMbUQBQMpoF7I2t/f9GljwhABKti+RuwdePc0gogtGZlCTVvei
JmNCXf85h6ZWCSmO13ADvucVNV7RXa6TPJDoMvodOLzi432ZC3jMJOV5APGRmnalt+TPoWnXDDP0
vCk4WC1ZcjSLsjkZ5zT19e+b95l1ygXLPbKgGAar5dE8fLW7wwLw5SWhwLwq7DN0gtjS/oncXHDt
RI1DrUcBh6BbX5bvrHTiCe3i58PK42BVrqhdYl5l+PTdcL4mzklxwG+gl823YID306o3tZppdrdx
H0c3BLqUl55HaM44FHI4VgdWkFXuupxTRK2UxGwtjJY5GN4mJS19k8xLksKuuQOY7djc1JboqgZa
CS1fY5HgSK5Oryq+8D/yb61rrX2eXQU+EZ6AbiBMsSBPj5M1hS6n49R5uLrH47wvrk76QdRY4fiE
PsKRzh7Lvd3I105AI8TEU3VIm1HbBS8QbdAryYw8907DxJDppG0mCv2wb91wP5gt/FWkqBHcYmfm
nR69tVfubAQpgeV0H3VBfWajIOvfYExaACUbJq7QCojIIvMxzzJe4RDYw80rzkDVYnZ02oPtsRYs
S7ftn3UTOXj+gnYwsGp6ebj2SkWOCKflllG5a/7z2USwrFx4poxX4Ox/8Xsge62/2IOGHX1UaZyR
2kMOgAuxAGQfBcqZbSYWlvA6gw/oXk3YLT2Vrd3/MbFRldVyX1GfceMStzLZBn/m0vUhl6Knh3f4
4JeYcQNCjw4SMLBV+b6XO2F9nzv0aVuwRBd4RiwApDBsjU17zajoK4Owa8EyTrPj38elfjDbBfdJ
6aH1aDh1+awLYrGrtMXrQ6QhQfwY5HRJl8fxjIWjYqhG8an++h0eUw2a5lpYmiqlnOBaRQHNir05
re35/JyvOBLmn8qybZaRMJw4MsL5i/m8yfeDA5XT/8VE8RCtdb5yxebxlV/xBHqnF03PvJJ9RAWP
xYZ8HOgFk1iblW6oIg7acbxbPPyOeD1HnBKl3bdTJoHQuMQKjGrahzpjWrmC/lX3SI1F4tKZPxg4
aSeARzvCViM4kQnfBEwaEzXQkJNna/j8KBx9G3kjRS4CF+EasEFufqkcTaD/YOYDJe4KGnpDV4Rz
LhkDgC8EupdLGWI9SQcEyzv5kI+mN/QEBhyT2Lb5rIxQl3hjE8NbYWquVsDobCsv97Bd/jqpaFDd
kNb2NV5syRhIkv6W9dnx1z46UpMIHBCns3d/sBzcNUTm2/vMdZSiDPjRTTRjnkqJ4J2M3qtbYl2P
DNtl6yWGl6+QISvjbhtu2fdGK+mFqBryhOM9UhZ5py1vBEEsGZn7OOelaSKGtt3qF9lxj7g5ffoh
eIegyCtjEYc7Wm+7FrhYip0/1W44YTct5L0MmPA6jKPwYZ8Ism7VMnlK/AbXYg7YdJ55S418WZi6
3ZPB6zvG7suEl/+71V4Abvsx0i7KpdXnt8P8ADv55JcugjXdwxpPciK7gqnNJDKDBvXD8N54t8Ia
+SZnTfabP5gfPcpau6RFBykJLJBuOjDW4A2cMsKqZKbbGh4tpoFwrgroaU4bhvtZfqGjPMui0Eeg
5L7ChYJfPzVAVBGhBxuaz5luDtZwm8qqIh6kxyL+en6c/Tyg/hbleKURl+yY/gAV0ZfDfnzg5eu6
lTgLw8hTmqZuOnuN4lfUU9SM+cVg3Bo7DVXA5fpzlAuZELBS82XmKtD8o20txCYGMrQpUtBpAMPF
Bmk6iyTrpIagy0XCa5hCTVyaQJHdQ/3dKKhED+ACbFudZXc4HNl+CH1pC344a/tBqkw+QikoP6LW
DM4Fzg9q9Dunfewi1F/vVMLWWCDRRtVVZLlmUdKK6s5Nu1RxKyhm0v0oT2yLqHk7ZCPkGyn5QH2V
6QvpBl4OmohkO4BU6j22oX/UhJtvmHfhdKUdeP80WeYbNXJAPaMXQ/gvphVfBQxPi0gGlbcvsuNd
/QgIVx6IcXTl/CTDxVH4AJLMZT+dtgrO2goEpsy3w8i35zrIF1ctTYWoEGy7kGC44qZ5lFw8UOHL
8FipCSHWko8b5SPtmPSySok20V5Z4SDx1BJyOx92nIAisE0E+Fd38AR4mZOL9trf6YBEyOHvTHdC
I2p1kCi01iWVsoFGvzKYLih3AwuvHZ4PdiMwqdVedZJ0L7IuQiEaJrl8s7qUVziWXeu97/c6TnOh
JwiTA4nhskAU98K0TxHO1EvLkLgIsEq64YZPhZsh7BOyVI3GTUj4E3qZiBAoyMfnRzRvNZ3/HvQQ
fFYv6i8QEIdjvvY3aw7c7ufmE4FlEv6/gCQFUEyqlHPeJzPM00HvzlEXKFwZhpQes3hEFCwS9fy3
gxbjEyxgYIbKEBu7SahrJYor4BR5O7Hhoq2OGuvJY6ADD2Jck6n56F1gIUvGk6VYvBfsZ6NnoE/a
JM/1h3mOuT2/UfjChZK1VCdwA51ISw7dT0ZIOkMAAIMbIG1/S8uPttz1+5ViAcZrU1BYG0S+gQNa
XvxHJEM/k5kONduYUQxpLVt8A1N4rzroXo0/jzYdSYB+bf5gCx8eM63aX8XxO90j/vm+lszdCKsq
sH3ue6Rz/8k5IEha3jLdPtFEv8G+lGHijneEKH9g3Op8n4ChWwWzKU4aKBzBRqmCjm7NRiEjeqW1
NSUFPU2yQ0Hx1ZKUCT6eB9ippsba4eWxmRmu76OGjIyeyFDHNvmvKdwJyKDLyC1Q4LbvBUxqCWU5
J3m7jgDHdPLUwpoi2OINBZYdxQBeBTtN9QAd4+k3wTXMBmPncJ42C4Atl6HHhcSmSlFLE0dZrFa7
2EwIw3t+L6mkPkSsco5RYtox10daaPiPZw8MMnLCHVHCBHGl2lAKUUTU729kJlyN2AH481bf25Gy
wSEq3YwqOfOrVIfzSxtsFQXKiElkhxtb2uQQcNg+67FscHGqeHN4C21ORTZJ0R5ZyiV/B+k1Dw5t
kbYd3nesr7xJQfie0I7+53L4Rs9lHLULdF1y9LKTq262ayCjXRwRse9PfYFRv9fCtKDlBWBJX07b
52gN41CoTvdivJJN1pGBFHY9Fzbu1gt7gYetawUTI3zO72czmcZ5/x34yrAUpLvf1EyhTGeRgvBL
zKq0F/azWvgKGTAJRp1wCQSWj6iq9QBYaz3rJBlXsR2VzRsmfF6GdQ8dxf+Bqyvv/h/SFS3Kv6e5
w4K8PAU7ixEn5vUX94+rf246fWyb20bRfNhpdk+JuMFB4AAzNCfU3WGYvQwj0499inlHB/bsO0GU
eENj3eNemTPxlDDxo6ny5g7sYoxxVq67J72cI89ZVULaXhVt/0RjL/f9etxHnsfNMdfe2Ap9vBam
Fa8dFLHBnnMLWNc4a54TYAyE3UdpF7L7ZMx46h/ebtbuFP8Lb/wCEVQPs3pnlYMcVqV2D23ePR97
TttVV8+aLd1yLlec+47ymJXdJQaVXGCr50EHgw4iG0odEGIBd0ChLyWoDUcOMGfjRQrlMbzUtBB3
XLOnGJuz0yoN8+adKMW2k11rJGBdfVEB+fefTsDlNY4s4QQZBrmyWM0Gv2IRw0MNgTpCPwvO3uLb
kWAn9M1RDvYZnI6xbAwpUsKXxrCsAlU28VvuKgb3+nz8eiqotriA6BvWN8HVn+LAergw1U61bXJm
V+q3wvG6EGtBTmL/MfIJ32lMzHnrRUJp70+q1Li5fDr1FnAMD3fcila9vYTHdZ3N2u/4tPGyydTp
qdVf9JQsrGf7exTEStv3M7XPQch30qtKGuFCNymWBNwOZUfgU+o4/y+o/Qq9tnoBa5p1XfRUfBmA
BOIvJH+xHGOmKpsA8DyBYZZhvdeaDOcVwI9qvfQEBe9AF1vzk+QCKGWAlJsfkonGIFgpXK5Wb+Ft
kREQczstIshRfpXJQ9yf7VLTUU9056uSiXIgeGzPdfUIjF1+eXl2PwcyC3C/Ep6cPoE2JXuWTpM3
KhTe+6sQHmdGxR7sMvSH8CiYx1jIHEYirT5KUpBOlq06gxxIBTKDlfWBig+eNJm0TCtCNAwkCvwt
tgst5szK3UecUgvBqQfz4UHncDoyoIG5Zz0SXsAXAIwCAAwDBZEhFwZcFnqc9cWeyf4gw0HAZvs5
hCvSgnh8TcfATmES9WN279CfrndJwY15AGJW0w5sreTmCif3KhpOO/I5PWWg4qYidHB6OQtoL1qm
/AHtFQ9FzGUQacetTlEz5pqNvI6w6Iu2DAu46hMPUlTVS00QzfNN/Cgj1TUcedi7R+Bnaycg/GAB
f8lVSYOwXlJWwI5YQyusmfa2fRstyrRPHoR0fcBXbOuszb9WP8cqIq6CQau9ltAEoHMa1U2QMAs2
sgsL33RgY04jduKlLtFn7dYraUh4WAOOmVrzVWBgbqviZ95XAzF5CJPiGEstOgaPT8d26BUkkbPL
kY7TX3cR1lPsnq7oRQd148f5pYag9Mv5vSKFud6b3l67sEmadRSIoHFNyzGdPxtf/M50CkPV6LQz
PVMCvxvxEc4t+7ClVL0jco7EQFjwAYf+Ei1stgD1W0jO9q/e6lNDt4gUHnASd2UW8ubBVBMSv1uk
3fBt80GzkhzoWv5Rqi9sdpjK1yzolju1YP7tSC0ximLRC9Pva90j8i57iR0TRaZvzC8spz/sDWpj
fNRdbMujWGdIdweBhJ9uRt2FSSqfCa2YIsV2xhNmP0OpPOu1EEYHfGiI/FM+CdBYRZoDPIBSC7g7
gsSW6N2OzIgxBSWouqaOEOa1OfM0/FIN5WZYupKPHmaIdyBNxJ5Euc4948VDZjnDn72UgUIoLBXP
3TUgxEJGyrEJE4t2PcOl0eQsZUD0MuYf9RLRvioW8G8T+vii80DPim5rLe7auEwTfMwGbg+g+TfY
9ykhgm2z0dnTcRRbswtqz1REHQELNhYdOyPUnbptOP2i092lERikIS1DGrCVH1KEGxBjCUTdyJk9
74p/iPWzj92p2Iv3cEUuGRIt47ZHeDb9Y6yCRX2dtsTJbO9KWeopwOfAd8o0a31T5rBSepMeMoQ+
ZaFMsFJQ5p4buVdHdzi9ia4GTbWAc0NyWWTj0hBiVzEya/Z3y+uFOFmtjijlj14MksyC7/RJwj/9
EDEEzJtPwl2835j4XhLjWdzW/+FccGuJ91cvwVDlNDgl3if5cTEQpx1wCd+s9i+CARqxuuL92oFG
CXSmB+Aq5fp3XKJ8jl/iAuP3KMrQ/opdG261GsWkMsdjKmYLidzb8wupV+mDeAUTq/n9JORQr4aD
95udjH4gRNaraPzwzG44ZJsfgsobyzFjivzDouF5NhJ7i5r2F2SrMuwkO1fhb/QFlD1S5/FIIOfw
4DNZbR7F8+0TWVXL4JJ2/RKFHfbzfaK68o5rEhyhl7qLOvlSi4HZTV/nIKx3AkkTryVIHH/al0Iz
a4GJjrf5IzuMC4ne/X77DOZOfmGtyvnaWylAs/FYolGkJKpceFYsshNx52BHygl4cDJRKImFJgJp
lloxUhcunX6rQOisM3fTYh4cVdVlXzm2QNlhivgxMXDIGvEdnQjx2foZbP9NoU5e7shcm3DlOJvz
ISK/UlTTOjyTIt1CWGp4BfItTU6zmwYpsCyPz2S17qYqK5Mc3sIOz9ygKpxc8zNTnK9y+jc4lL1A
onmW7T+tdfwgmrBX2PYvbtDNZ2u9UJFqUvQVoEbtU7qyCtcHTlbd4q+C+aHLDVKDGOG7PTWARf69
64xBSV7c9Jbfl7Q4VsE9bt/IsW9bBMCnNTWtDVmp7VYSq2HetC1XvfNlaie1WIgn8aqz8T6+1vSu
nE+klfWREM8PDT6XbfKe4MW2sxwCB43xX20dQvdgVSgr7gikZgyz/3IbFPGw0m0uHVidYN3ZvRcg
Mf/gwc80iCqsPi6E+F8s64taI1d681ZPht6QZ7a5z5HrlJAFTk710EisXCyFYjbr8sGGbXE4atyP
NOXIYuST/nwXwfFOagx65ts/h696N/tMH6TdCNCf43w8jZRaeB0XVAFQ/SR8NPp5d6DUafT7AuUf
nZob174lq885IqoYXNGJy/SA48EO77iW4+KSasDN3DsnuuA8+2TSkloGBfb6+zEaBMjFdHveh8em
eGgjQ17vY28J6zlFSszUVICHTWKVBkUgWJ0hElQ5TXGajjVHreV//KDyyvsgxWHXmUddiYcnpAI+
BYfxfcyxPR5gClot+NANpw4EiL0ju7psl7z2wzM9twxuRQjvaKp+7t6wCrsvd8JjTNakTvev1HdE
1E/9fzjOF1tKwzu1kNvIAhuOFCkX3HtalnrmGsj8lionUSavNYRtY7IrMTUp7L/L/1k8bG8N5Y51
11+WbI4sfiCcUvRrb5cExcV5slmAc5iXYzU6nJsy5ularq6b3mNSINMXFNa4qSnBmRwiHcB2Oq0h
Lt9HPrdFpAJFbISvp4U8A873oe8DkxYORP4oF3qcBI6FTc/gnkiKefyqjcUv4/Rp0ij8H5wYz6fk
BE80BCHBE0zCjwpA+NJxNMaqPUpHbnDPWtsUrST2ouR8oFRApp2HgrIK7NFlwtGyeJro92f/YdxH
1lL1ec97o1n4+dQaXpsNNFwmtWtPlgifPZP6rQmfuND8Dz4LUBtwlliv3Vw4VGTiP3hKhEzH0HNQ
In3LC3JlXdjgpxJ0nIA4uhIClUtjK7EIUKyojp3i+Tf/PEo9xq12ztoE3QEBa4jxmc8kDBYhSQmw
0WbZUwV89FHb2TVquX/tH3AF3WB/w02vyFsOvyZ9HKLnWwuWAZ9lwf66nAK4VlA/D0dEyuAhxiVM
BUerbItjIJVah1ntW1ZA/ETMEeJDvvDt29msstqDfmPPwkPJeBP5B6UdpcZdg0IrQzl4Ef5iNcgX
I+m3sK0+uM157GmTlD01twtdmzNlhUq6LNhwk3R+mJMJvOnxF7wJkKK8RcJEtTRfzfe8s/iIpEUA
e81kUsGHkUV+h6lc7RB0nj9/BOdcrs3TDFglFSlRJ2Ec1/IMyj+8uzNiSxu5iHx9YQyB7CKMd/jT
qAxAmxATGyVOT04BNVO5ibltI+DgaFV0aEyZ2y8lb1CV0sQmfiq48hxsSnpLFG3O6rSmFVW6WhK/
6mFMUimJpUSYz/Ik6tpFxIPvxZnqWMoF9JrSMQtVoUFiNsP+KA1PfoqkWKN6EY7+Lco/NNeVQIft
s9qp4zipPq2e87lI/nODfik8/au7QrVjX/NiolfjhojEsJA96t3ZJu9ZO/+xwLEYj7Ib3nv+hNJV
FhiWsK9JE4z4meq1n2iGBYhGC+GWMKyXeMUXMdZXJ1IsGitJ4FHBzFRvVHAFnSTI2ARHRyxGBC+i
X9YSxYKbMPymbpegJDCPdQiuzFeochsbU0u4EheDFp/Grga4iME4YRvhCNYFgOINpC/iP5F6moq7
/qh1ztEXrpm36AgnK2frymFgf4JIB2QlR/FHvV3sg2sIXs7+S8NrnwbZMbabNZ88dpUI3tolVfrc
iXXeq4Zoc6RFJ7V89Q22Ht+Y+yAKoT+Ls4dOUdQBltpAz9A6FGAXtABqSLBj+P2ff3YqLU7Huak8
dGlMGbV2Jw5ao4vWkDJUQ/GGomNRx+CqMlQzfHxt1qh+A8rDqbMty7VNevcFU6IOJWvsywEd9MVn
u7C19wepVYaCBNOst1zZj/QTfv7tfI4Q8yrY4JEX2FOPt/Wh3JkQJAbugxelPoc6csuTUlRIN4kK
LNEr8fHfFwMngJ4SRepU7nLqulhJSiOrhqJrSAZW+tkBgGHYeXo06jFn5C/NRwhntT8sxWJByMus
rutetrcWXDySfFSqh3K7uIU3anp+d3qSXHrkFWshe9LZqXmwGjGS4hdJb3O/H/MuZg9mQRE8Dx1R
PRbsKvSlOYpAbNr3JzRlQ3KGYsuMabVcl6xQWEDqEs3TkDbkUe5vOk1U91qSMod71eBQekXBinZe
0Ael+Fy3NwTDa2AwaukrxHl5xUSF3G09gkOrp7KHPOhHU0y/X4HLXhTsh20Imdcr2/r+eVxRGXft
vmprbY465Gs3BpJHRQ5KcyB+kSSTed4jIBjxM7ka4ROX4NvJgVD4N07qlVeX1Dlal6Mlt0iEWFrv
rRwOEU+/wuer1xw0VVSBsSnnmHpcBCfuEPYEmh8dCLiQ+lBoQRMSIih6BmHCwy6tEWWjwFYlxYgL
RmuiaayPiJ+e1iH1mIYzSZqFBYPDBHs3ZxT4WpWiQdPs5FGVFnovHwWvmRI5Ds9ha9DDvbK0jm3w
cpCF0zhPOxg/wfQ67KRZdqgt3my60wRPOAjAHE6J4zU1bKrs1CW/yfKB+M5IbMySfF02FzgG+P8B
AVjO7yZPPYtI3t4pgsJAy/QMEUuMMlRTJxQvDuHjYKMKYmpADaQhu2EU5UQXylDjFb27FHB8nSYh
UL5qCcin9TrwX2w4BN63Kc9thr8V4bAiEHnByY9PgEUNufZ5bQWrXS0x1wHIivEsQsWlrRlS/S9q
SHoClwnUGvUZ9xihl1ZxlOw1yIXWphJ2jeA/g12iv29LVUn0u2dB7PA4NT/169DNvW+GUgCh6ZlZ
0Bb2FuW6RDLkvJzXy5w7jBy3cx3D/1LXyX7aIyskHAULzHZ6U7Q9t5WusBsqPZe3iAVTEnKkyWcT
PjtpM2ISxM5K47GBs0hdgD4pgBsZw0sEYWFNOyG5SSWpmgysRcmJU1ChT7PvZFIg9eC/qt7T6P8e
qok3rj4ol0F5lVuaweyHQiE5/b4ExMxgP8+G9ggrnmNjFGznRs56BTIwl763DQ/tXWDjdvFVlSgN
2TkfdroEPNWRkn3gWHZKDghuR2t7wJK+FJxzMouEzsfYZmDhKHcNFNM8qMoxvLD/lY0rtUEDi98v
eTFmO/3j29vGyRbvpWWremEcgZDahTRVLbOCwXMtna6qdMBLB0ivs6T30tg+elyH4i+/k1uWBGU2
PtAa0nBgTjHdZAX+oVkrZiSiAeDigoalbl+oOT44QKztT8dBuB3OrEp8xkZ6nCyJY0s+3rlnxHAw
FLlVR5HG1NEEtfVMK68QS484C+5g/znssSarGni4vBVYfOVDj92yMclhJpAjvnD54V2oyiu6HaXB
KtybbkIloxInF3BZl5am/ScBkY3sT3XXrgj5E2sfE2+fkxcTTIzD46ZndYEKlpo/94muDJCoW66X
ttU/yEthr3plYIxEUJ75kLLnNtS4WnY5pBgdodAsFmMgTXuqC5xKU1PWd6Rc+f6MpcYa5xNi759c
erpzgKvUtTZvqJWxcDp0GpGB/DXnsJY4mMleZym4X5F5ira5TDf4LuN1YmryLPC9YMoi/IlgNVQy
NtAOyWHYbhaaLsB3rD8HkVyIf28nCmU6PjN0T3Ckgt0RdFyRmeV/MbfXj6VygXHlXvgvqfsHdAIT
GcZtzXEt63nwDcQ6foxfE7dA5A2v0IOshdPvZimg3ZHae/AZgwt59GHZdAIoRahvqMkxiUFDRD1L
HrJFiy7dp4pxwLOYSk6quZC9+qIp3WvsN2ZLBFRkrpPzKHH2U83Z3/aAQYYLsEabBkWDfCKvTR0L
5EcOuneJwWnOZduVqCODDNKRdx6SOOuFRELVNfM6BKs3OQQZPCx5J7LQJOqPzXjPA/hQcuwupkLZ
7a+gYpTyKiXZjdnvh2hAEKVOHuMsdJuly8UBtNNpshiDPC+lrdYN+sI4qjecP4tXUclvyzsySCvu
RTynokPlQXZmjNEpOtbcesOdQ8K1fxG/7WTSbYMofVVp8Vr3+AkUYchEssORRInQ8ZzkPGlh8uBI
O6k/8kXDStXXfjIvdIQgHCFrNTtmDY45D46YfPerSPfpB3ySaY/FF2qybmUbJgF3Sj+Ra2EBHzbk
xuSg+qMcTmJ2S/5FIXRJkR7fj/y6zFjAVHgFpswy9F57xig6uXgx7Lq3TsObp8R5bFwbozt22y+v
tL0PT+vfn5RRVyGNvPltKyjdLZjOOvBZlLKLVK4hI0OeYWj75ho67V9gHtKDdFCQZ1nmOTHfO9JS
LpkFM9Sr6BNmI5hmMwdzHCnsIpFQo4qmE0NPkDcYa8JMAa6EdSyhFvKKob25oCm+nKKf6UpfOqkT
yUPApV6C7g03CYbwG2YOC+kvG7Bwq+vvuyK7nQc6ii5dCHQJyC6hNFVkrD8mnP8FmkC/z64X9aoQ
Yx58VvKaNNjU3+oKj3HL+GXXc/hsFi2+5RsdD1CcVN9q/F3ebxHUfoTULFTQAM+C+HERMtND/vLO
Kyt13cbYh/YU0jzrs5pG3M+Ht7yX7Vr+CHPXqlxo2ivDvH/FqZS8/qSr90HCFmre1prgf+ilckFa
kuZ6+/LOLzIeGaZKHRZvzHOBx8MNAgoSkz/PVFcPTr4rUKPzHiGvh0gAIh/aJG0sU2d/8cOgV96w
6A5d5PP3/barNmRfEXbC25FPspTmdvKsBRstDv7ahk2uHbWzKwab0lQNufpQS9QSilBquPVu3e4t
lcbMIlTUfSyeEaBi6CkBlVQ1xupBLSYvuXuwKvVDEi7Mnh6VaAWc75/1r2v4Ch8L8cxeHBdeUzPj
5hhpoAmc0dIYDcvImw9BVL4h0KSeEi13AgKbLC0jTs7RMUAUjGZHzmxhWB4jaOt+l3G4IpCvd6S+
LNpAlwhlfMmAVsOx5bQvyG2c05YGrAapzbYSegiNjwZSURfj9VDtAD4IPRfX0iSc2CGjDX1L9sni
g6EuFRME51PjfRhL6b9tuawmj8xpNh4U0258Ux3PKCYXAwre0GKDt9hbogG4ll7/Jq+jMtZhmC+f
urAkxnK9UFVjOVbgV87GCbDhjSwAlCh2uDZ0G8Fuk41ngSmIF2SrEpqrRIVufYC78dth7Ve+6PTb
x26vLJQ/uFFjKizYU6MJzP1JCKnw5t41DMMWS3/XjcFuBhaSGwn3tiKkTS9nLme3eBGA+HH9E/iR
ZWP1LKMQ8r/V+W12jxtTVWUE8S0aJ0pio8SMHjHqL3+HpbeO6OOCLl8sCEl5m3fz6MBL+ZU/vqGm
FxZPfyXYebg5ksMA601GMJz9CiOEfzcJw9W3prgruaCvh89vfg520tpuJMI7oaReEdzNstrGwXsK
L6jf3H2A0vkGNFFDdT7nQkmkD6jGwLg5fudSFuQpQrwxgBSLngXGQw9orQqaY4ITakJL6A1cEYbA
PcwMhZUz9tNJrOtCqYekqsYpI4OY/WDEJDsQFZbunLL08CKt+DwaYBmcOb8WfxuFrQRftFzS/5si
heWN/NRfu/7/WXe9cB9u2sC3ynSvuKPdu/bN15rLki3KAHmywOgi9CquwYh+fdi3z/a3T1mo9jiz
Nuweqhg8ZeHfQ+AmY9Xqi5zscENmjGyxK2el2nHGjGVxhR0ct45y/xOUz/yUHaLPu+3n3G5vGFPn
+Id3FA0Sf/oUGcWeO6JJozMHEGsgliR5LuxPAaTSwKYJOeEYMHBLUqorZoUfKukU2qFne2RSxXJb
4bf+Vas/a9+ISqP/fzrLBkZkSXtCIojruik73/wNSRg0RWFK08BRYOe0O3Lb9nxZKY/B4eHfGDCv
1ER0Xihz3S7gV2LeetTlLRCcI5rrDRFW3yyAfBY3cTdIyxl6rqSM/cfoGZ8ZiNmBllh5Mt/xk71B
/W8mOzb7AcobigLNudC/RocKIPvrQ2hkvQ288Vak50esjkqX7YxUIHl5sjXV/+imxWXTy4A+hV1r
E29njejOmrC7BlEjMM9mRfOebNXKZZHIf9QKNPYT4wZplijHQP1/4+fBHh02gec3vbHImk+zCD9A
ZMD5qdbEGKlzu/Wf5eEzUN9T+VMlSn9sB658GGmqvYkMtJfA57yU83qJA/PFw9tRoRyiXf8BXPhB
Auh5/NidkKJl3j+U9MD5hADkEz2xJd0Z75Qm4L4s8LYT5fkY++akwrKkF9Y0kCI7DUdwD2AEv53s
ENwpeiy7kwJ9TzlLJQivWA25ijZfOap/vbcSCQlzQZBRoFzDX8ObDEveOEng6lze7Hxb1JSf4R1k
olcxojSlq8kP4kitlIxNB5zusfSJg3Z341TMavbpY+aeNnfHrnHm/LfLHOBbwNt9LS24bmmj5lGh
NO5+UkxPmc2BlaQEXZaXjFR/P9ypHBQ5+ktNYtBhd2CVqNnIF2fIRxkYpXEPmZtTIaQuahlnS9Kb
qF//Ev/nw0YWDX77812vs/NAB7jWdnNo9aU+8pJITUGFyXMW4zws22P91mEQnPqfdd89Vb8n9q2H
ffzeS/SMZ27nCTUfBaZt21TEqjqO875XTl3MTv4FHg1qMOmLALtHHO8jswq8mdOtGvEU1GiS2g8J
eKdDGhqko5ZOq8f58q0omMZwSRsioTBRFxXAbJtx9QC16Ka3cgEwawe3ymp/qOhdTl/hgm9WfIFi
N0bUklOCX9ATMyJJ0xB6xCgoPuoCupxfVdE8ZvTsef8UEGIG1TLww9PfNLUSgMUL9vm9YndIe70x
zY/z5dOpxeft5uFQ7AAnbSGHPC6IcfoB3JGe8m58bRWfQ/YR5MmdIe9LVqs3MAJ/rC4Sl3njKGJz
mrkt3NZObC0eZKzTk5rDhPaRgWlB/oZIQzrLKq7vwZHmMLsgzauZjMkYqs22olSQ+Ense1SJRHXo
jp1di7Iz1usX2AIy6x99wyHEVDjoZOJkNO1wiFpDYno/eTBd4kYADRv82JKk8n0DkIlFFWGPEQoR
mqqFmvA8JLFMG3PWx1Y4NIsRPjXPCLGFchTsIjGH1DEvj5J4w8anJ1qQj7rd6/2DKxNav3PtFw56
c8bhLnoAzMgu4z7f2bXKrmut+Czvti0915uFyAVY+xYwYmq50t3XJXHUfvhstdzXKK4ieywoFZw0
tIWNaJTsjVjBHgdBTvmFSI/cnSNZoxo89VQrZpB8ENSVJiVlFOCLSWS9mpgJaNHj06XuSaJ/N+aE
ACTtO031I3286o5eGf7oNYECJwdDD3Q2bCwpUYZ4hvo4kgq4P8ZldO9eS57UvPp+WhyBBt40pwBQ
EV4otyb0hzQv/CR+EeziPsN4eJaffQl545IRGubfAR4awpVamIgA/Wv9XmeTNTBQLzM/8dJ2DHp+
dtFFZoaFIl/LLvrnSgY+kA61/+qgaqiUd8Rvp9s4gKb7XNuNI01xKQOUvlkNljSWLCxwYpMV3DZ1
bJnMKwbvi7V9Y0hKfv11c7wnZ1qrsQLYQ9ofGYI+MQCZVf5315xW93j6OGDoDGLViilNG/tfq/js
IpnO2/TMdVMqPeZ5fgpuv5Qg+yNaJNrRnWgPNzuAJaUNZriA9WGzVhlWgeksSobM/h3LV+dA8mt1
yqfdxXwimMITZ0qipPoWDO63jU/Qb5j7tA29zAsB52FoAxeC/dsDxB1bTd7VnjNXAZpguRkpjLCR
5heXbBGbAtwt8KsbQ6otwJFss0wqjNiH9MXuSWXF4LmTkTNuOs0sUX7culUKi6gtRBquzwn6yvUg
Zu/5KejZbVvJEUZoxCUXiyFiCBjsfDWz5XNtqisjIUwpb1X+oKtzqUi13yT4UOBRyf0y2Qy8pr/I
qzSZOnPmA1Hy0WCjUeEdvv0NuZiEdXDI3crSeWDfFW/7efHqeb2BspcXpUH5FMMvW3bGAJgZ/a20
MYuEnOpsUxUJgZx3hVQpYx55JLIJvpSz7XFy3/ADjpeET0vFl4oGtQs4rP13PsD+j5TVm/hiNgwb
oqIW57cR3tr5DzB/H0JX5KuN8BQTqQrgUWDl2bj8kHHf4HOReQn1FQmhEwanHyGY0RWWeFIGi7h2
Qua2jfNz7IelkQzNdVxdTMkoNOCZqKPzz+ISGFxV2Fw56JhjICna7tSP2MdV6xEZ958OvEOVgLLN
LsVEG4rjp3ki1nMCRuM65JfcCP4XcN2y5HzEom1Qkf2b5hnH5/DKdune1PjwfFL1KMPbUYKGdFN8
20Opw/9B+XSHijAztZkaGZDN5vBCESXcC707QOTryGsBsttRgFn8Uh3KQ7YJzBRNvBxPHCtj56Iz
wtUOJkgCHg1JvCNznLA02rObg1fvqm+t4H9jNtfpWvB732jT4+X2vV5bDSQFjcPhhutQieHCgPAh
3o8+CKCjmZqtKwNsDQaMOihd24VEdgg3Kp53BoKdImMJZDnXmp+aoN5tEHXCT+u8Z7vOi4kMk/op
nvlwpasDVE12+BVkmNcwJMkjPV8jksu9O1jQxmHoGo8Ym32MK2egUgqWgqxZMpqpFTjHK30WOuSB
3siXhjy3mMO/ulMe2EutF3f7MaMFZ9XkSQ6WTMxKmiv3W5H+jfj4l/BeUmfowrV1arOLrRTGoLc6
o3CsolHMlSmseK8oAm0G8Qd5mOE2dQba1jMPNcQ1ePIHnXVa5B8w5Vwufpp2Vw2EWIzeglaabFyD
VDipNhoqp1P+1/841sFMARPaeZAUdGuY+sZA+6WIglcOc4OWR8vazXnLEm9wgd4hPyu+EJyzKfTs
/GOibAUawEFmugDYW3k8imtbo2OLs/Z0GDlQNDzFTaCvhaTI5TTMhGlnNj9DnLUquFzDagdaGblN
iwrYwnopqidZTIFBu5el01wXk+pg6pH4+0KUtiYTEattM+C43aIXJZs8KvLLb6nYg0c2vMDs8mJu
oLP38VCqShkHGB4xcIAjhMpLGG29b4VjpbXAb8B0YXNZyjHiTcy1kvk7GRrC8AZwl/TjqHiLnW2n
Fy4yR2gs/gOBM4fv5tKXxN66biqZ/jh0dRdmULzjk7bcg2D0dXf9tZW7E4AMNTQWy4TMpgVhZqk+
R44O0gtSTnhdM4psa2knig6T3gwSMCbFiTo7rsSTzQUa8ttlOnpfl+wRI7zgQWadtEfDZ/goF5mw
jDZ+dBXZcTEFphefsOAWIBan3KylvvE+2VS4/xv8No3VpVSY3nVHCR37PguGYTAgxhrb8+dTaaUG
yOzobbwNWvPD4BeXHokXAR+GyW8agiNiJ1fEVQKWPDqQcANXwurZ1qPou7eA4aHf+jZeWaeOhYj0
ySfgDHuid3KKTvymsOARX33WvxcFkTShAje7aRlWOUQCFq/zKc65e/itO+BwrptiM8UNKOc/8d4r
ql1xpxXppJU7SFLqXm/nVcJ3uQ7tFCBXdpT3is6vwiBAsceI5fqKoaosGMQe7Gt8Mc5cIaB/J9nP
ILjGbvKPyEvOkQKraU21c6aJDKGLNG6Zte6XStmPhv5IsBsxTrOO9VTrYrWxDSaK0PJPQpQp+FL5
ijwNVx59XFsll/t8sW6ACVg24Yl4lkHi5f3TDXS1DL09dsbdJuJ4mjEEBGtRiI8Ym0dDanO/l5QU
bIWt0TIHTUrDBX7xibiOFGh+B/T6PoSLvmDllDudCVbfoPaRgIum6T1e9/3TkkBcC0fnGyJGsCt6
+RG9KPC6WydIFvMVvAs8sw+SenPF6qxqoJzeuAueQoKOQW7yz5bPsCzJnJTsBf7tQ1hf/hHpCd0G
+0EAOp+tBVuXWp0c9deKm8Jx+VbhRXH/ZwiGWieA8OKpCFai1g+TW+ZT1BMPw9AOIdRz0ArC9RVP
SyMqZ3dZbcE54Hizpxdbd3OnWlPZZwol71VF+h5lvsGxcOiB43ZUB/r4kdPv7efVMDoe2HTX7DjR
o5ZXllnaatBweljTXMceC3tHg7g+2Ct2wclprC3l6VcDUq3TdJBT/LPsaKyGpSm9IZEhwRWq1GAm
qiS0BxO0nL1qYn7UEbk85z6qfag1E9tI6JxoRkaeoLVToqVLlXxGhJeQYCJ+T3JHAelO7P/zXNMJ
33zFsKIAt7CVJAAqIH2/v54VbuKpSSyZHbm61/cuKdUz20rPTbXmWR6nPTSn8qEFajTy3uZeFQqU
ZA5B5sW+PSgFe+sbfrjrfpHx/7yMHX/iKXagvoydc3x/ejkkoK3ux+hC5hWYLwl/ogKy+d+jx2NV
1odiqzrIbJDWtroOCYEbf6KKtAOyXXhc68fDVtaYCcRkaBQSLw/FJH/71zEqrww0qqUmhdBlBdZw
vj2AwWyZf0jK4ZJSWv9y61gGr0Qb+yMnglRcpNNW5tnDOoUBPlGLjxtxuJNQADYNXEqvxmXquwI0
zbtxym0ouJcWlDXeAAYAebE2M7fYJXX8ghUtWJB5O9efFFJ/0GtAXvYhfM9XQMtA9s6OZuaWBOby
SnpuHZFvwin+GA9xja+M9z5FIbSbIt6+w7k4VUz08NZtDphyUr/iI3NGBj6gup6jWQd8kNuotVRy
2hTpxFJW2BH3ijRZbZpLsGZ0fBwApN7FJDBVzvnbNvHvSgzffu2tIV6H/KbvDBFzfatcw+B+Ef+Q
HLJBYafTYQFICZB2+ebgf9pfW2z9MhkLbmj7f0Gu73exlcDS2LkB5FHXSJ5V8Glwt/T3fuYICeAn
QakWCkhglMqzpIKPavpYICYOoJg3StzZJuNjTpwXxPUjdYFOzmUAmLTKoYZ343P/Fis6a/RI+gnA
VDC9EoTsiBHL99u07drF3a1BHu+xQkDZVj/LtUA4WyQUFSkmLsdhuwkfTRj10+l6zJ8fwvToxE/k
+BmLcm5OB61WTpdO6MLrirCHDy6QqlWJjhuw6P1UXvxLmJzLIY1bvoyV6IgCxgMWr7/q+znUSPQm
F67O6auVuaBYzVMadFyzAQtyWooQbZZaDGzLh5syYMXWP8OWa6ZIiUCHaDhnXnrVdhlBF+D+FVtt
Ss6L8XFOjYAJMqTIss+n9qT8oUeOaXSrBudqxKajbuoLWTQWlxVuACdCh3uF69X0yPYTZfGcKqh3
NbI6nDzp1T2u1CPNxnoHlhkzmvU0nfGU6mTnBzuKfYMrZfrzKx9y3dAHre3mFAS3nIzS/+5gHZvq
tg86mkLjzyLMlGLt9rb6FYfFFZ6H0gARGTAAoFH2PsQL37+3q3QqSkPUuoEwZidSlpd3pv6KdHx4
fG1YCdRtiLmG6XoOEqio+fO4k99eqvfs9BX+zWBCPLBYIDvNLZtLlilINybGgv4zNJqkDHaVMgAW
+3QGhnQ/CU630HuNJIgM94r+LfZ60yFSmk1YiU9dQ+Eor+bZ/vTSw+y6aTgU3oxt1C5FH8cIvJx9
HuAMerOZsG/0rPaX85rdmSJl/AIwdjMG/ae86245APJ/L03vYLINsQwgsKNrs+wvpttfLT9/ofO7
UJGeEujyV3/btRoWiqXmR/yYxQ/g0Ru7r/KcDUQBW1Oe08t//xe7iVJHpA5M8+wDWMrVFFpR4QuV
VaMQzFZhtwlPIa5sEebXsCmxw1bQ1+3KPQYC8Y8H3rK5T7xZjsGeah/ZUFv0zp2t0/6f8BnjHTGn
x4rUkiTy+x1qjGyEf8jl/TU7e5Pf6t0UAlhuj6rIS7qs8NrrfHGP9cNIt6keJ+2JMSLaPenAA/xt
73R5IKOBH0mGEv5ankGzfV+0eBtlySlcBD8Be2uJORcr59lN7vzBhNwWcwLQhN8539cV6wWRJkVm
N2roYloG3YHomq+rX+0c5IyQLVmAn81/nVgNi4m9diRi4AeA6be1lRuDmf5h7DHIJEla2QzmGj14
sDP5l3LYhztwdfe/cvvQw6eol9CdyA9Xwjj6QFF/2+rxZm9nk1nSOG+QFwym4tI8OpPm478vxflb
yg5u+bKHCehj1XnNrCN0AK7Okfs6MiCC7lyd9vRBVV6pzg+F8ODDvVOlaWCudtQ2YdswOVX9+9z5
dzoKRf2Eljh71+XkdTYH0t9sf1NlNM5pld6gcb97kGCtGCoxsiaw9xALvsI7NuCiCDdyYv2n9Cf0
NGIVknd8OI8hVO4JgS4jCatV2XKP895ThZDBYft10ZTYYxrfav8uislfihogjyCSEQhxeSIYZlsK
tzqsXo0FgY79ZYGKi23V7zDprwQ3do1V7kZ+yshxZsNLh8WotoE1oJKoSVHqHyfklQBI0vLjiHkz
r2H3gU2SxqfV/rO1Y9fkYs+a59tVqs3gBbprkO6SToisi8Y6X8wLzZpmukRa7dMEPAGXNVldfRj9
T9QJBkSHSBfAS/JdeaLl0DzcisSeSaNVrp4Qeo33ZrJ9ViDSSafHDhJPNhjZ9pFMDo2Vkg/YQMEX
uQThactPmgGb3mSn+8GekYBJIpIjcx+ZBjf6PmSlSrSjEjgdToxdhoJOl070LEcCAjgy7av056eG
6dBTRz++FxaHavDnmZauRJAjnY1x0bRPax6Qj1hEuEq2lYo5AwenbM7b1rdarxuHilggLWoZM6+I
q07J0go/QIHBdCbhLF6vk/HT1NSphPunaksNzSecSNIYClpWK8NOvB+cJXW1OR3ZWDQxcM9HzN/M
xus45jQTEEqWFxjeafRF3QkkfzYH6JvUKnK9jZ6ZFVcF5N19+kL8A72vtVgVrQNNq5s/O2o//2lO
fkAT4JPIjkk5sbN60n6awBntoq5/YLRB0MeQwZv2GB9DHJH/vEWF6M13jCn1k2zDwCnU3xz1tgiZ
mqHsvvtWZhDCRI3phTksMD8r2ly+O0Pq43d+4K5aWtOPMqHWggdQ+1PfsTl04DoXrAkvTe7b2moO
KXRzXrAiF/kbBHguD3eo2DQG4ISX2/HdiIeg3IMVdck9myq53+5eWP6SJr39gMT2oj9Zwu07IUOZ
c+ZfQmCkXLqDZxEhXD4hCMtdVrMBxpYdM2BHsPCiApiuMxWMVdb2Eg1qcQpvoKvyD6qoHNx+hTXS
3ZjCmkeTtFEIKBvy79T91dsgbGV0Zw2Uy5i2Tlh9YAKuYwnuTuDQKDohsR9EhezC0OZhJ75xeyKq
El/6fH1C1AbKd+/+WF983TJRFZoMzV+F13hnHSQ+W28NfRXosexeVE0ZVx8PT/H4LVw5KbpjhSxk
V5Wii+m9zWunqjDmXs/7v7PJDLr/CRSKocDi5VztqlvSwILUeMFabRhV8qrVllug54xAnJk7A3Ph
Qruqqte4S/tpZrresh7UfoIT0BGy6mnctD67OXtmHvueMIgqzYOePUE02KD+CDgA6BDL2LyOrX6N
O2ak3BHrr3SB3cHd6vOKGV7S6E2r4zbvh4xCudX9WVAA5IS11fSCa7z2HruRxS0nsEuRjCv+G2yf
8RZ9WPaOms7IkCn/bgsambP1gYNhkCW7QkEBJbBBNhfZr/aUQQnTWhuDMxcP8zu8L/v1nclmV78y
g5obEKracPGt22ynQNxVnYiFLU2/9Pjt+z8tnLzD/ZAkmTEicxrfb1mOj1o6QmkXUtR99lqEvGNk
52A+NTXft3NM9bIX0OnF+OKSR/hoAomXmx409jGwAOqDZlXRLjwM2IDhvv7cokQ8rctA+4oimHjs
Q19KNlr6gQ1W/RZScqIgAqGMQVuUG7Mkf4tsOuFVka3g6u0K0l1mKQ8R59+wfRwkf5VD73KLQC8C
ii2PLogDQIprNiS3DLI5CIiZRYtbyPSFQqDqMvNp8ceocrXpZ/+mcI5LrmxPNBKGn+gHt2U9QQwA
DSEJ9wAvRS77XY6MOlFaOqC0b2K3gBrZetbP/uybQ8jFf72O9hkoHods4itjbWo+aCJC6vDkVIjk
UcAQZwfpqR4oty5buDCne6n3sIK+NFHM4qzkyr0DkLNV2aFA5+8EH1z92Itqz8LrSrU5qmN4Gy3T
LMPKeEin4TpM2WfALGW3cep16A1UW3nv1Wn5eAM2zZVKjFeb0jDOek0RMWGXm1ISmt/ifVsBWk2N
TIBVvFONguanqlL89fdfX1565kj13rbmByz9spTvdDfyZWaRLnm0jhxmgzRY8ff8DsFEsnkNlAid
56VzgV6qHXSbXL1+Qx6TDt3lahytJVoKFGx8C33jisYTdFbNy0+8yS1XVdpyUzv1PFQcY7Q/712x
hhIy7CbvoSUFRJmCA3IJs/YEXkU1DToTfVnAGaZ4F+QJiFCAe1XbccGHtUF6k9PUkzymM+tFNeRZ
VT/hF6cjL4IVTuX2B3h9iPDySd+FkMDtR4Qiz3/Obd/qrrohFvUooZ1Ucy4a4pL/i9Fv5Mg9Zmkd
Xdy2Z4kYW5MeQyaRG1ARL9AEDhwNQ95BRVC0+LMDB3u9ZiY15/EjL5hm/BnJKcWPZKFaa/TvPFBg
JhUw3qTIEEcnVPPdhi6Y80HCx+SarwiLMFp2qPLA8Bqasfnzu95KotXCvMx5Rc6Nz6MKkqRdpeMe
DMAQm/QYjE1dX5wZHafYRj1JPC6qAys4iBzk04a4aIeDDmdlD/fAVZOm/wjDUN/t2a5vuQQVNl/v
DWj5vUKJk/c3Fa/AFx54x+DRxV6CyVdE6a4KERo2zdp0q0NIGcPeX4OYlXARlP4hAC36lRDd063Q
gNjzUXbd7Q0c8as43F5a0R6KNxc1NGnHh0zigG0uxwmheIv2oiNNMrKb800foKbHEuxt5BZEKJAY
Cx8xiqQGKqv5m9zfwJ/O62uV67WyKm/Bche7oY4o6N5jdVcFEUgQkoXeqsf5bft+QxzGxhZ9rqE6
BxsNVB8ud/QT3JIwbHVDGjto2clucy5IVf9BLMF0NridVbAg0AsUEzCMboHgHVACoK7Ne+fsvmcz
l33DCqM+fQTxRPSSIXQQrG1EtxCviBQn6WsVXELrvgMFKlckhzgxtlN3ZWj8DgWpEf2zVBqD17zE
LHxrY5XFPuGPXb2s2S9X3RApoy5UGQkVd45fr9i481K7ydb1u2kw1mjNZ33ZEAXr2ElexgYCQrFf
6Hys2WPhdjlwXJ7gPZYFLk3KuoFqbZ1LrfoFwY1fkDqAc/2pVmrP71itpK3L1dkugSmK9htUy8+h
I3kKC3Sy9hHiMCC2KEjSn5ypi+yKW9DuDuEB0LxHGTWsSoObS60fmznfZacTbM0eTEEYR1VMVAhg
X3d6wR91Vv+OeB61HkRq2Qoq3zx6RL4WDsurxbbDiKZBTveksX1hf5klPcxHW2ptQQ0JwQpYo/Zd
eEIYuYaSX2quRwgqNd1S9nSHoEIu23Xi3tr7tVHjkJDKmabH30QEgQPdpHlWcuSwHmDYxbSP/bAv
DaxV1ZOUKDYn32Ps9Zg9zfPF+1cO46QB9nO3i0MrzTWsen3MNwIL2Jg0TZcLeL0QKBMqRv5NVV70
fJ6H3jut1CXqZUTCI+r/kXwt+a1hzvGgVTX7duzareeH/hJI4JFCreBLri6BMJ/cR7f8PaQyc+6u
vjfPMBZSvXY4hF1dxR0B7irRoa0p6eWKdW60JqYidqfJhZ8cYB0Au5uY6BcUOBWS81ZJe2l5J83Z
YVJmzGbaXgP9oVfSFoq5R648Fl9diIglmydwQ/4PgCJ4cugqvdgh54rt0jNaZPJIu3Xb86y2BXgc
3Bx21SSNoCNslo5btYXeldV40mWEMYZWXDDmp/5SJ8FriHzmUllbaaUDbZPSDhQTCfBDB5UFLCeX
FGvlS/XMXwO8eLG58C0JJrXT8RW+Kv2xeZTg5aW8dLrl1CfP0Giin+dNVbN4hxKroltrxrUtc69G
U3RYandrYQ/NmAlopCsczua8Twg4oPxhvJYl1vhCP+QOuMOaj8Ma3HETWr57iEIvFpWCAJAeX584
9JEu+phoj5/y3Jj3S0ntOsBJJWuUqp7yFvvjxcA3Bv9bvIy94wew6TUz8zi/oAHJDfLzTYS3rwpv
N7fo+NXnjdvSqyxeCPIMSpXsYwc3iY1C/Qhpit7zG2JiYeJPY9+vG7d4STLUwnxf50+rrcXXubux
rlajZKIDyh+sMLB/pGIJbf0wi3j+mQ3uzjU955M/FyRoxDLcFEGeAug21AthS9WgMcKFaqWCq4xT
2pZNzMNLpC1GNomfh955KyV2ALF5+Xq6uG6t6hj8iePPc8GFTgbSUqq2sK7Bt/ZJLNOltx5XEvL5
4uHdouHCdcRdo3n26OgkFq2r48eoowR/5D43FxiNmmBRPtyf93PKIS3iJoi1IjcIc1jYUsLHbvSL
wW/qju/Utq189g06mt7n7Sswzjdqa4c9LK5dRYCknreD/PH3tBgQ9x6LnvkpWvMEJNU5jbMeb29/
BCFTD033Lj6naATe5XMJ0pm2ufY9gFkgf8MHtZIKoL/fNscvuaS+7Y0IjyVsk0U4xDfpypTC0v+I
hMCegJ6Y05PMGnerjf9s7uSabRiYEtKagWx8c02blN3TIJAlcRrW14Qhg9b6rPqlOf8OeatB0ge5
7Lg8Ad8eTnuguhdLFF06xLgrNY08vcsPF6hDkSkwDwEX3M1mVZdTf1+/Lbg6fyGsZtkjvS8xqngx
izuIonuNHF3+Rnlnb6p9/xeihO+q3G0L9A94/g6R07lDdXCA5l/ZlrmTR1uI5iUAuqDR3V941aJs
8gXOCZGGy92iokUNZ0M3BmjU4u7boEBEaNWu26NKVS3jrNUqm3RKgnT/eNkCvyJx8XApsw6GHKfk
l20VbuiGayfNJRBcg9NuLtgRv2IBzG9U4yIhjrMVluAdNfHfh+yKJw59A5SFCWUP/eit0s/F1nYI
XoMw9p1VhunCEOq1I/ZdKXyYVRlxd/8t+cKo+LdWbBTI/3bjfIJxjLcI6EHYvve6NQKSpZUIbeQA
nXTX5QZoJnp2z9uuVGJOjIjux4MaYqMIxVNYl0f/Z37m/jhH8+81sDY+uejQFYizoDRbCyegZ7H/
zfC2jaju1u4CZ9QmZBoQlkYf98rSf8Zbfjhmxn0ne6GCZ8XELnce/XtRm+y9gChOsRz9p1E6DgnV
rZUu54Clt7HbkMmuoAvpWwnIujC9hmAgMpRqT74uBHR2MeGKiyUyNWopHWx7ejXkJmKyjjJ7pqwP
iamENHVfOBK4Q80kztsSUOaimGocNHFkVUQBMXvSGfW0cfpWa/9/OqZsRN5TcH2p/ec6YTfOROnJ
rRozwrZ4f/Y9HHPs5cZy6OMFsq1Tryy0DXblrysEXk+y+4TZ8YWkvLnIcx1BGrilA/pMUOLP+N5l
bhFL67nGYZoFQdbxNQa0PK4A5ouzuZZZOPxQrC9pMW+0uiXfQN9A3/klM4rP7+PXHM5o1k6nrEiC
Gyt2K/+wP4VqBy+g77ta8UxUPS76l9xR+xugtCca4PQKNknSXfXd0yHTyOc+Xw6gI8dEByj33VzZ
JdBY3bzxdDQnPhOHGiF+me9MMMtJstBgLjSgk5j8N1N265isRBQiCrgMFSCLmihEVAYGncUgiKGD
NvWMLq+KoGi9IkdYrC4YPQ6xOtLAZDJzSJTSyWg9ZBOpwEaZI1tZeQEJZ862vVVFM7sS0HDm/Ft0
oq1Z+YKI/PL9RH3acanGEplIQnQLvUCFnqhLv4bBo/xOoD8FKp4eEV76b41a5tAa87wQ61znGcdk
JwTGgn4KnGiG/04r4BugBs6fnblO1v2gy5OmABrBhM1SWjX8oVunJ0IG9+l9vU3n/UzldCDU0MrV
qvUpCbGK26PsmUyW8rQf6ueRIi/X1ogsD7p1RYPi8V/U29S++Tl6F2dGGBQ4dRy4+uCtlS5fylWa
gpIeyVQ0R8+buNOrHbCXtqeKiB1R1I7cEgipn2dIjZxtG2xtmAk3+RcAnpB9DSyjnRJxJ59tEIYy
/RGw/Rwaev5BRjrQfAeV0qVHZTPxrtbAcB67XH7OCbhXjaQZU5jtJFEhdp98Qn4mXv3N+8+BmfEA
He8L416qQO8rXybHvHs3TOQzcMoPb8r2qXfwx+VO7iUFjdnH6793W4B1sH0hYbqXJTxAg+jJsoM4
St/wp+4fshGsYzqLWcv0VZBerHclFhFahlbSVg47PPTfCy94313XBpLOqi43anuDbUjUGBefmGtq
Vd8caZEl1+ETHe3f4t3NFiRn9/Ta7Hy+bavvdQJxVa23rj4sDHd9zZjKVxAXqU59CBkc59eMtMX+
2Rcvx1YqYhkyAwPmQ3nZ+CpOJl6qECT8kcJJR2z+sk0kIJl7lm/0sfyPtsFJxVLuLHHf4H2KTmC8
+FdHobwdZKbxaeavLb+kmt75RjvUpp9fB8EvXl2JJ0g8U7IVkftnlkHTBKIRFJoWUrTNCDdpaEXs
tPrWO22rcpr7ONs9aw74CMjUdJ2gW8bZW6JQKbtLAtpUfYmOFyEXVjcBCzHS+VxuV3oZDsFpcTJn
Cy8iu1BPEc4hKoac6NZRsLi/ZjcMAQCakEc82C8cQR4kDfZPlHRjrI0X9UITq1+aqhM1MFjGRFSb
qnpC0PjQWW34bJtZ8EyNA6q873I6/PrkAPYGerJgtJiNSOjWMmM8f2zc+goBSNy5GaBQb/B766zj
/97pjwZYQ4IkjaG9FLoIl9ujfzDzQLE07GiCeQI/qPMHKNcVW4tXm70KIL60pCSAbZBIhtGiRJf+
y9jfUeNxRYBYs5oK0aP7TKXPyAURvQhAuK9miuczvQxosPE2WAXVNr85wklDIzRTxL/8gCIsuI8j
SaWEsMDKIg/ZL/1QJDxYFvH7mZP7+mFA5Yxa4Emj2lNnsldf/jDWTES9IRh6h5e08pexEoVHZygc
ZJJp/ApDPA/RF8Hvztjs9jxLsyIksZyvH00Np51wAZabzAP09UEJHZhlSXQ5ybeNmk8FibFWIuQF
N0xY5e0mjWJ7U0YhoY4QmfQKcQwivOUETZzR79FejPHhGcOocA9YoOfSqfrnYPLLhKiAiYtydYko
ODxdwg7zNfeY6iurwvS9lsDOSEzbzfkmdNiXs38vbo8fXNlsEzkBFvE6fsuQYRcrImW85KBfaVEG
igVGl11S9N3jp67lBEEjVsD26Y5K3fcWgHaHJ5+OQDRQspw5lTMj0vAXlYljUD7E5AWMu7cngF8N
L+bjVenphJR6z4PI20biC9Cdlm5dQVaMPjyj6FywnnlAhXhl9SJw32fqxmtCMRwkhW+vXRQ8XaPT
5SlssqMdRYnpVQEaEqHzHo3ggS5oX7kQ2gt6M4G1MNohwJVqCd+V5zUI8XiYKTHL+Q6iPNo8mX+v
mo0EcMnsggHXR+OAHkpEiDyi3rTIVBiEazQU10fWnFzWjOfURBKhu+ELim1W2bNIrdBKF7pP/PDv
FhJrbDv1dY2a5xt2XRMBIRBFRHbi/T7z/VGvOHLzVx/yrJxxrzU8OpI6mR8EvLhXokX/QmxV8SZ8
BK5Zf+tNGd+ajzBrh/m12PYaEcN2ekwgM7/dVFzYVqOddNNtrkqo4vgnf0uSfCCnOvlhosjP/pTH
2E5lnBSVvU/rZl2e0tmpSv9osCuEurFnOhS8vqpPGpdMwN9wBPquaMvQFyyTb1dbLRXRypsPg2Cb
J4L7dpkf2FAPn2OBCKNnKSECAurRIczVireVUvLA1PuQAAyPD9wyT3b5ImBVE3rpW8l14WX2fJIk
Idkw19ZttZZE0ecWHzU7ZXqtWmaN/9RHR4uPHKbZRj2JgY8j+GnKKyBH3JQ6CePN4snsr2EO00oZ
eFU8JoQnTPxaUxOk/R/8YGQcF6ZnFHyixuFQYeYMYSZVMJ7+SjoZI/qVMrj+Em3WdRryX03qW5of
E9yBUOp6MFGQYJ/IRPi7zRncbs2jB7o38JmUQUGJFuGWTn8KyCFdJcLmW7k7OjCPyBGFT3Fc+P7a
+OzYXrZ1IW/hqAH5bXPKXfcR7yEZHj2t6naFKyY2RaSQk7Kg99LfDEo9d9HoyuI9UC4hmqdRQNtQ
HT2sM7dvxqffVL90lxMJyuI/PrJQMg8kxG/hqtEpJUhr1S0awJw2PtDYn4NuQfVhTOrJrfW4fzpa
XCKQnbrDWOxFRfh3BtfKRcvlDhtamh2YpaVYb8NxWe4A9ydObMZ72Q2CYqHesiNOh9kippVeumCB
tdv0nsny2nZznrnuMH1vnCw4olgGtQ7wzMPre2ETvdxkRT/jb/PAWrldXcvXD1QLLlMW4+2UgeG4
x6GuQw//SejBE1okmjzCrhrbKWdlpbyi/Aboay0Y1N9kHFYTNggQ8NiJvA3QkSdoGVuFeJhhfgg9
zMC20M6ERvDBAlNKFlo7LkewsosbY4MNlaK0EWLDgjDl0o2d3NNlVJgkiB6QyNDlcTtpaeLHUr+U
z04DpNP6imFfcMIr39h4z0mEcCijzaWiql/n6TAKkQYgK0ozUKL9ktEFuWlLwXu7FiFoVVY0gCij
93UQubVH7q9qBHdjNU9oCtnVYBpeQflWP/EqL8aYF3kTroEqEMMSF02wGDHmC8E9LZ6PxNJpScpm
CPRKTx8sv6FGstsFC7q3mwnhUcQu8FoUL1lg1UL0+6hlweY9bLxlNP5js73VG7LZmgj05BnLRJbZ
FxOiLC2TFCbQaSpk9XiS44RrWsolZqKWThvCI05/BuDYot3lHEtbKF1M6SMDrjk5rkLfuSvyLj8x
Y2urN7Dt5yu7gBSDwOi4zadk62lab7YWPoQF59oWNszP9s7mhpnCcMfG0UJpuyBbRtaASOMcTjqD
2KEpQVVUv4TP94/Bu8IcXefC7PUH1LsJ+fvESKhtyFmIK4UH3z3V+Yq+UMqSLh1gryi4mpJPeyOZ
D/B/l4bceka7TxGpOsxuajgRd9XHO9S8Oxx/VlvnhAXOPlNAxCpcQjFTbZJT2dhNzmMiBzNi+7mt
uxFURi8MqJedmhtSwXbR8iwb1F8gR2l8ZOdjjsDIIPleLpsEpHd/Bv6Mhphcu9zHXIw3XAvLLpr8
ya4+6tKt3OyXpfQ8zySuJ5etvPVjdyp3c+//wcYojLKb44DuNUmnP9j6y7G8vOlQxcQf/r774vzp
F5BvBMERPEUioemgz2eXcuUQ1jWHw0Vly1l8/spvaCzU++H3umAoRgybDBmFOP8FlsAIFnBUjTdA
AOnkOynj/ZOnvPZdDECbCfPQW7MUmOD9GlYD4xVzoWo/DrC9bwr188ilhpajfvYqFuFt38c/6UAq
cuOfXci6fxlaU/eUJdoo2Nka4IfmW30DrrAuPy/KHTADN7XZNeBFxVo8M6/vf7eGYG7NpIul5iFg
+Wx71mm61lO9AQKOW67jOi2AVKtQxk+SEkPmolZ+dgYKiwzfZHQz797NYoSrHmU+F4N3z5bNpIcY
hvvCeQWd34rROveYsBkeBlqi4we2e1Rbj43lVKUhiGNbRa0ioEUlj2DYW08qm5l74HVwEQICFFtS
SSf4KonAb+N/EWVutdFZfB60kcXcqiW8vXtcE0utj69nimcwNYmBwoJ8eGDfF0HDA2soPmkHcGRu
muSJXsVLZN2g5OMHVNGo7B3Xyd8N2ZCi/fB1PstXyxmdbNUVRv3QqFYMfiequ22q6eDSUwoDCgG9
OFaCh4Uy0ojYld9ZJ4itTxRZgl9Y1SFJFHaqSoHzVFOWTT0j1TlQBcbMrNd8y0kL9rd0yJKOnBNm
t1BPEWrUGyVh1g7Fk/ChOYMJdY3tssLDrAn3eigfaqhlFNdGXxexH9Yu7FSWabGWaPnYidAKKuVM
5UaLfU0TIis7OaX/o40sz/6gmd4CXWZ5GjC9qEnB4iejbcfRhH4NiUHCHg8AAlUFefMsQ4/Zqp81
YluA3g8tkaeVtWGUVBvw1Wfg031AAK/rZriPJdYBtncOnxaQQpXzUIY4ACbxOYv1iY67CqO76/3J
yLfNb1743trBy5fqoT1g8X8tATo8K4/PMUewOD8A3Pb6QJnAGvabhyPZgtR0SDh+P5UmCjRxjUDv
a56FhOFEEGXadliJFIzvGs0EoQEr9i3zjT9WGLuMKTZq9paLWKcCFoAewK+D9rIXUBToS59k1jhL
rq1iC7eJNIird9YYGCpd9Vu2ccCqiINa+guagmmytqa/cLR+pk55FsglVRLXHtPgQKU/yY/mcZbL
LIjoYG9s/9bhhh4JSCnsZLShtPNhE/hazzabTlpe7uvehqZUkZ8ips+9rOpyRQ0UpE2zFEwImEex
2OWRDqMchCIm44dEsyXvWheNfVlrEI9RtGvu3Umlic/f1j/KCBlQn0Os2lAlu5aaVVUvj3+mYCNq
Fzg3BlKGidAhO6E6HY+Y1ONA3vyoyWpg4zUOWAT6wskQAfNJ780H/8ONBYRJLZ5exogAyO4XM8+W
7+vbTojDErFWYI2YkzbNi36WMafJqdnk1i66aPgDwp7XzH74ah6X9ODrlMYmIbVHzWec7S1uTl2M
4WcwREDb4NjJdn1S1+6rUlbYAt+IDWmgAsXwSL8LFuWeCoNPbWFOy5OGn5g+Q4bSVtKl8xLM3kdG
BdZzH9jRnP+Hu0DNT8F3wIAftJlJ7sPbDGq7846QI739OpTfgAX00PX+zPMbcNW061oXIpWx9ZDf
1HkglEmN8U+ZnGnDjELZfXqDGKfURhREABnwBk4jfqlc5fKuL+TciFs5OVomtIM6EFLp53avWz3H
oPwS/VefuscAWunMcoTKXpngVn/tYiQtbCqEuvYQhF5f+7vdqV9oKVNKT9/l+58S3LuZ9giBTdDa
gcEPHCxxvrW+NslmKKmOK9XhLKHKy09hU9xRchfil0ut6Xo0QnMuCym4+JxluK+VlODd6umtpeX3
v1IN3ieVVmO1Yq3Xxo04HBI/dQ10RkINHMZrMlUzGpys//7HV20MMcxqH3GEiVOyR3eXJuccJ7Gn
6ye70KK9Vk1pZCHlI9/rxIJrHT5x24HsIZQ0axPcQXkY8QqoTxwrGnBAuSmv4shVowJgJeYBOgfD
W9YuzPeueV5h+d1tP1sloN+klXhOyIDYnUlOmCzzLUzOgBla99T1gLohhg8Ry3tXkIZh8ubhlmuz
9Hy6thW/Rmt0X2DAJEtwLBHqUKcCNj34B+JHmYKLisz/rc+13viLO/ZddjpgNfBOV63/d17+Oyzt
PrnU1reb0z5D/GXPzpeXd9JUWhmKj+UBqBsJI7aaIYjT49tEJ6UB7X6hCR01rimC+x0p4Ltlj2l4
Hkck2LE+U7Hno2W+4zwP7NSKTjxLMXG06WGF94a+Q/h1HWy8Ui8OeT0ye0CjxrxxNrhNfs12+vqh
N3mro/K1k72vdJ2enLOA1CFhy1cSsRH+8f6v+bNj5zrq3ij4q0anhIgWIXXiAF0Dcgi92L/m7dUX
y1l6uK9i1Vut/TB4L1LkxRWiDSI8alVjrc2jXGNy6sIrirpM8dzW3ny9nCkirJ2Tds6BdaNxNHYu
QCPnnA7rn5kHuW8Cj3d9rX7PlI7CIDWYGXYvU8QyNCVrjbqYhkhG6IWVhZllk7n/fiXTgRvUhIbK
m4EEu6nPARztXtIdudaRry1BETkEeRAzh2/uEprfNoZNZMsKkShptBMLZe9SNs++BeN0CCAs26bj
8GxVWDEvWGti5caiulXcq0lQ9Tjq/orvAye9ahLNef73X6cDv26NAj3uU3fnoiD0RfwvWVB/+j8Z
kWCjck3BvZjBT+js0iAPTUnLFp9VHKNwGzaLphX+vFCidXFoJI/GL5myfdASvqU9x6CchDVCS350
vLnNT1Srr1nGEw2jrlxHxRPwa2q8XxnG6xwuf3p8n/x0LOm5m0f5Ioe+qujYjbm89sgZAdQoe3WR
2mKW/TWmFXCIDSZv9x9NFyAoR7Jxi/f46JvoSPuzEbsgaSiYX8+JcxuVZUMzxXAjbFcdMeunl0F3
Eq/wjt2CkjkngZLel8EZRmLnGyZ/m9mCgFgnofcxGkXz3R3PVX5zVtzXHhXRB9fnqFs1nzgMDRlx
v6blW0uR2J65A2GBXwesntWKm/yIiI99bo9oknp4CUWKQI6P+kXrhWd53TfB53kF/kcCyLV2328b
89rIRrwtgpHsIXxQKXKxjwJB636A2BPvUMhGcOt/NMMCR7F/iQIzTzc4DT9hlryHDQaQA8//nwU+
EhcJwxJckHzDACI3U9ZvNpZCa5LVWmM6CjIbeKkpbJzsnzNMLMPtJGUN7zmFdOHUqjCZAxRHqpxj
2Mx105VmiwJzG1DM7NycDONAuaRFqMtTVykGFpVkZC1SNX8k6vWnxbo0mqW9ZxUAmJ4A/QQti0H0
BCpuuIIZAbcYFbAKz7S4iteA+ZhfcuIUCPIIabQjnxNVErklCig0BD4fl0sfPsUUzdhlPNgkXon3
jl2ZfMsboKnoVIVhRgVOTmPUiLr8QELKgiaXatoW3vGPO7aZts01UIeDUYRofEUpJTWVzcXS2TVA
0q755FmdYD+I/J+Caiz0hnHB53RgvbKaUVJbC5AB4gL4iFB7FMYgvoEGpNIaEm6UYFwQ4+2+Wn8e
atlAqSJ6mgBHHKGXfSFJ1c0wyhPuJOIIHY57HtQgHQY4kwQN2BTW6ZS0E3WS/rIxlj0c0fv8LdRZ
9LREPPkmp9wdUDRVyBhzuhgL/J4GYvl2piSHgACGZbyKAOLltPCL6fTHI6YYFUqq+ZHLjTKqJLyt
WVVwnNBXIJbpFAvHP1ydGvCFbaDj9xztKXDXtakI/sWjLR2W3MbzyxwG9qSBW2WSu9N76UiL0Fza
kX/16Y+yVcAV38f3gPdCieF/F43+/9X8XYUNkf7Uq5NjfBui4Jz0bVUX+NYZxazt+OP4adZXy+IR
sxIPkGILlfGETurAJuWGjbcaLRZY8IH11+Eoq6oUfUmzihSbabHMyYCkb2Gs+Aj3VOij0Fyh/xa5
RUCJswDeJB3prn5bSurY3lQi5JNFqv2lbprYcjyTrUrzdyg3T3rQa/N6IQXX3s7+yqSkZ8U/C7lG
uzQViCuOyjpTyencI9ISOXBUip61b+tbmE2gyI7LAJHuVNNGJnOr1KCbsiB9tJGN+v0R8cTBUTuu
9l7vb0drx6Mhfycg1U6xSHLQrBnyBRde6vkhbZ1muMSK/hfumnu4EFW+IJYoAWKbqyWXfXrlbDMP
WauwkMECl9E41yhT8fmn5A1dqF7DOftFWalFz9ozPMXCSLdOzvS0XEi0dOzrKB8CuP7W2p8rQanh
AErr+Yx0vmVo6krlWDbcv372643MLZLoJ7jjn0Ahz/C1LiDmcJsvmZQTMKTAAmNCdgjB7IAXjUmd
1wjRt0BtMQ2ptNh58Ny9z0ucMv0rgDEyctgDMFUepECpxOYVPa9+t5dkOEhJPBUb9yJJuAzmPPvq
zSqYFiz/N3o73wUytiOgYWIFszJpdO6nvzqPJr3DPUvFMuuVVCAFRJHgtyqn24PfBj80/vRzAot3
+mz81rNFwEq7fRZx+4brQUOymXTSMAuoiZAvPKfzho259sBnsOsBUUu0mfVuJWAgg9uz/laG5Vmj
KYFWQY9eT9FNmb18iJyKP2lWS6KFp/80FrwI07RV2EcvpkkvrmdaUx+9waYKTqc7CbKjRSJ7htgh
6tVIpp8nklW2RorGd/1ij1vJpg20xVmm72CaAp7qo5DC4OBxUX9iI/QCYNBNvG44xO5Y7Wk0uk90
I0YPswP8b7Ga2F3gSWE+koLQjud61Ugp6fQZqRUMFkNM+XoxM/hABksi1AfNNkaxXqecDOLkAdCT
nli1VieXmLgSw5zgo3Ef9/Fa8V1GBoo75uEurSHjO3zVwlY4cMv0wYRudxOjlIYGE+g/L6jHlSWX
VIuGvZ7bhltDh7nf37TK2ZMFJLWkdPKil2krmIonWrO1TXgTtCYcNELOEXXFGdRc69HlIlnvuKUb
V+uUiNSjD0sDuwv7hHTmCTwy/jT4rIF3Ccc4aEjvDIyWt1iqCSFpt+5IXcH6brvQIbqTPL58VJOz
UHw3Tqj2pexKJHDXncnpXQmGz8Zi6PPaajQr77oEr95Vd8+RMH159oa6OFWEkwYYse2MldMg3laR
hWVQQbcYQ0WmOMNCjk/LCS8JzOXqjAFmnEodWi+Ziud0RI2E9Ul06T/uAC1PkUwVJscQlFL7ajYu
G06Kgzgti6/RUZ84it/qL9ymO9uCwV4E84T1br3nfYxlF0xWy0Mp8ABFox6UQrNcvsP1/hUiwsEH
zYr/plbIp69vWUZZgjvUH0YICuy8C8mxm2l/UxyqFFsbwgh1KWQxqWBub1FCTwHXBjRY6IK8Otdy
JgmmGNKehr6KVNcBOPLcNDBGUjzh+Xk6UrgPQH4E+ZlIw6GToHiXV1R/NmZehw8RYIBGgFQsoDpD
WmDL+97tZ8V1A/5Jwccnbf+V3ORFueW/xv4BLujijrFQfv9q5SHSBKGafgUli823Hw1bYWHWomaL
dvkeh9Vs7pYnWQ6K+FPxXDLOi5ETk6oxEH606iE8p3onkNvevI7QUpjxpLlXhdmuCAPaeqLmnKFc
0rHHv1jM+cLANyMGZ0d97aBeMzUAE373n9GxiPadnVI8WiV1WJuC21EzjvJmOzCYeWzgrIYEzuwR
AQxteE+VmDPVkWli9CpYatMWbD+nMg+u1R48FLZofGnaHRcKjV4POjXSRiAk8OQVk5Kp2TCT/cVn
Isa3DNEgBSrjgU4z+4SfAAR8/A5jmE8/kfDvMBBQjsjdN+x0/Qk/Aianp7UmAJHxMFDKu4PLoUkr
f0Z0sBuHzw9E1GSLsXUyC0+mW8NpNOL1HBAuD8b0k00rKlXvNiZBIncLM17TnFtfjNJ8Lo7eYD23
3mo1FSb2ncvpx7dDNomAYubovBw7FR62UNL721o+O2ngAPPZkHxSopEyoKQv1pi/V6iSiu2rx4zh
U5mtc7xhIC9bW69Rkdl8HSgqIE5AgcZJAzWnL8KBdeh5WOhtjmdsZuiIS8VtOgoR886SYhO4sQOf
JFprypIgX/JsgumgvrlnfALDh5EsKOOU2pXdIbJvrlw6zdE3YEvyh231A5+ucCZ8kBW96KPln5sq
ASkt6SfjDy3s2NJnFAOZSCZEisgYSfZrlIeNLNfwlfmD2EilrJAQRr85W+0INlm2hAW+yh8TW3MG
LZkaddBxsk3OzKGyaWPjIegi52a1Ktz0YlEdCoZahBD9FYzOyew5/2I9CxpDtRJ+VjGEB2mHli1d
2dZPN649WMvun0XWKMmqdnaw+egNRYatiFEQmVgxGZe1D1WeZGMVsZ7YRm3Akb5OAQCQDhWzyclZ
WfKJu5NYkSrdmClQMhB3/v+32gCY2FS2wluj6vS0vZKOGmQsOkiEgCHVWAojDva3bl+NktccT/z9
di97PxC3sWAjzpNcUR1ARsdkDRBmKThrNrZ37DIsvvLziE8nOfoD/WaUdO6/3sRhAHo152Za6KpW
sA3XBacDAnaPjWhT7UcYRGePCRddk3Jnr8gOMWUYtmPEl6GQWmJSQL9nex6rD+M5yz6NxfZubaXg
vzDWbEHjDTgIN9Q1/Pz+BXET4pE3td/vyYF7ulwODVEPPqoeIC2Uh1W8K2Ht3kG9c48/FdLRrTCu
HN4oduWBpHgujF2S0EyT7jWuk+jy9rQXOQLBy1MgmRgiwPcGKtjlo2KOAQgbrIhsw014KHpuG9Ap
VwcFLxrcoe6aIr0uAQ2CnJNEuxjWAf3xVLsfOjAXZ2DUftNmTr2Um0wGYKiYLmyLGoUcAhnrAUSS
2mp+ZZhMorvkroi16CLj4CchKt+7tExUYoB6HPPLgU8fBRrTFW4RFB72WkZkNPa4jhfaWEec8mut
S+afQnuhyiCE6Xy1L1pwBEYUapUY+LYD2fo0NSNKXolyIS++7SUPcFuwdfNp2wsOtDt/hAn+appG
51KZtcFtNTqSYjGS161Pbqs+ocyY7z5NniD7spJXeuVIkKU5qbXrozVCH4RhVeQqBsnEmo7JOfNv
hElUjk/kgqASU4jsaNdHAzXOeWpnXEqcVeBbs2zCLWAyNdyW99RlUA1zP0VS40GX4vXXX/yM5I4t
Y5GPREALtZPft9xrgZUiYjaXVkzrHvtj/esWqbSOqi2y640mv1ZYWmbnvIWl/yuyjeG6MhpdKhp7
dohh7wkVzUTw71cIPHnnCaXcXL/v8Tve9YAPsMw/MiYIOQTihYEATL00xBbB2+0kfd+rViig1CDn
u4Zrip9y7g9TnvAktVkK+O91KS0fJ1jeS8wfpsniwxeSCrA4K+BKyILnvFWw4FPVrgUM+Q6Q9k8l
CvbwbZs8HGzd5jeXhuViVAztkAUBGK2DZ8QF+bwnzDkcxxFjJa6RyKZNIBs0mkwZG78jLdX9yT2z
asScR4a9tb5VICuDbBDP0lT3L/sMjq2Z/LDcny1Hy87ZV0VPg2Nx3YBI9RZP+Hm9HlxsdBn7OFt4
B4SyhPiikxje0L7/8NAr+m0hAW1J3Dow1Buk/rAW/fTQWFhKDIBlPvT84IFg0cLZ4X2Hu9EC1d/r
TK1RB4ffXQy5ZfV1Qo7bKye85jDnPvJEUKCTgC9iNTum5NUQFvB3uS1FhmGmfSrVXxMCyC+3U+MV
rs9SHDuNYQwPc9nPjaVdBoL7QzP8NKe069gw5yDOEkCKQqekmJEIIgcrBl0NTyfsIl2o7v7fxTE1
qxUg+mkg0H9rUL0aJ/QlINQGNS4HdfsSZqJZ32amvnQAqcrxXdzpG+iK9N2r3JRgvRI+KWhCGzzr
oyA7cN3xrFuK+rQK69SFBVaosFGyfpfevxaHE2D9upcrrL791s38Mj49RGzLkt4HdIeab2OfiirY
+Zqf3/BneiLruUvyyD+neoSPm2OYwQV9HbAFYkRJxutgDwIkjRUrSVj2diKUB8x88ic4RRXLGHU7
T73M17m0brA+6LgAZzXkUJYg+w3SMUyc+iOEenBxrkzQ1kvxK7z009D9G0u06A4rXFkc8dmEGeKU
oRhv+lAYO2a9CTGXHPlQEcup21AHa/RBTkANMWlkBBvhRdYjTAyd/G8WcnTt81NNRqWyjs6SEwtn
jW0zYbye/HMZqSAdzu/RwA5pINgFIvqaxc4cs1TLXUYuHuENUTCBowqc4d+007uJu1d30jGTzw2P
873C0LgvOEmES8YizK4V8IEKiK1N0ZCqRYVakGxNtcHHhc+IuqF61hZc16GTud8fqb6lObJ/M0mi
K2SzlOxH/mfJ229IvfBM3BKa1zIS6A7d2PZgxGw81lNhWQWc7XSY+lwr19xF4Cw15ZSIYrGK/sNJ
opEiTZraEir3+Jck/FD3xRmcrD0eitaiMYqqINhVcqTmvq4plmtCvtXmN5U0Ll8p3shOS0RCYV49
zL3YGycIlhZks7G0KishOZLhDcg0uU1ruEwdJ+zIOuxQrq4k5EZwvzvFqEDULu7OAck0DxrZLTRu
e88uMZlMJ7tWVkW8zJISNbA/orveC6AQ7jug8Ic2/zSAI9FdyYtiLPB2JAnbqO3PMMnF3FRCfB6Z
u3xWUD9qoKc6vJ57/coJYKI51MJBML+TkxBH5UL38rhyYRS/32Q+TY03ZY+wLxhdknZtxcmsU8kk
YToXLT/2uP2tgtikWtxkEQZPHL4sTv2CKmRrRc6B+N3H3P6vjIzfGNPs5AQ/Hlq11bXhk4q8YOd7
ijVbqy0K7wSL3jACs4E49BAjFgsOWY893zbanj14lncMohh+PPneaLrUNUDr0SCaoW2OBWJlB5eS
HTrm9BX/zrBOOauwoe5coJvyMYIH16quGT8ypj+njzQ3vOmD5ZCJHx5UhfYtf7tzX5mzfhgJ0/BL
VHY8z946t5DBxJKUIe0MsbPy2syhXxDNGYv6K1VwaikMsesQa85TBPGXkRsQWMAZ+sUHAyQHb2yW
xKljZCdVsQ8kHb+9S6G/npZ3zfa9hQGRvN7yDCk/CqjSnzadIXFD3FYD+iNqWv/bWjNYnnB9DBt7
/suKyydXWtuSTO0Tgl0eao9ncitLZPFmRR7u8HmoM9G91HGnmtHKMd4aEMDguczAmhf3/tx0hbH7
WzMHJfe03mwXRzjXasSA7F86dGyBmFmZlfhLyx5CrM/CfamnDzVDvPjcO4UByIf6ApnExlXjmg2/
/OL+MIXhYk/IUUN2QTHnGUHinZYZrydA4qmc5PqzlwTnm2ag71x6iBQO0zvN0nXzVujDAdKeQZaD
u3XqTSw/lnNl1RGCvL1sXlPQxIrcN0ktwC7wSOSHy0JTnG6uHO8tD/lp1DGzYQMfOOOsIsjIvPDC
8YNIh7APpSrdVvhwvO6/E6BABHW6/qrQwMHewN3B0GATn0jASNSpJ4V5zoUuvt449pHAI62pKSfv
kwHN0oWlxcDvEI0p/hVjDans39eBfzwv6WoU2OJAMEtlCRGr4i+PRG+t9wLZs/8X1bEVmGrNg32Z
jciyJwLk/PIwrxO3RJyUDbSVwsYfKPnzzGowS0IeahXcSdZpvC+XJmpO1xvwLhDJWrZNDgHLXORt
n+TDOBP+HPHKSgjy209/8p3JVyhCd/oRBcdmdEIsvAXI+ikuzmGBasYG7CpSa3GWcpKblfOvyNLY
dVeUp0TLew6ucbXvIiVDGN+e8CPyIcZ33w1gcJHvw8hPv7EsACONXJ9T/acZBC7GaO99H2lFko6X
jcfMZLBlyon1x+MvH7slN9N/Vs5niMRMj2Rf2OVwyCv2GGrPWiifuFpDJUa2FS3eZEAPQefizL1j
gLB4MkSQ5cX/aSWoR6mZUbuLWcJYudQBwXms+IEfEh6qMRlrPlZZGk0fzG5e5mUnINg/3guwPvu2
IdksvsCdW7jd89KwIkfFX96E6dk6Z3JgDegDVIud30v3w1OiDE+HXhLIm6R0v8MLQ/eySuHpOLBX
FKcVfqQZCDA8mbmlgVb/Rs+oTaQUbU/VIoLOiyzH2w7aGIFK3Odf49wphuffN770b+Vjw417QDgr
tjWhuMEEidjTK41Rgu1hr4bkkLiO9aSC0YJ44bGRNOKilKDDWacj9OC4ZzfzeFTqXBKGs3zYCBCA
LL3GsRaOzTSYg36Q7p4DgKW4wbDJtPq6dohXH5Uso3GppRvg/CSq2d11+B10oMppg5mRhNHMNxUn
aU4w+ht2SkVMt1yRBl2ZMjNgTXh3GfK+O+rmZI4rSYclAYLaiFkmCAwtc8fm1rfj1k8JOje2P5zO
H0jS2zHV7xyYohBzNW6/S98kwwYglB7/A/9mYtp+Z4jYR26okTCRiS8n80rnKv8t++oWFRXfTV4f
2m/1So++9TgwmuzhACMVcMPjk4BdyhqgfyJ5Bc44XufKKEdt+bjyAWb/b6flLHoCDcyW9Ywjk8yT
W86S1t/3YBE/x3B8Jmu9yynZiIxAbq776wtajoAXaPO+4lKlTUlaHr30ej1ltfz6+8p1H4We/6oC
OXaWtOsr+HyHJF3rYkbuabhvMp9isMt3uufZn5Pbx8sFm2giDDucLr5SdRLJy+avRKbNs/SGRYpw
G4SKV74Dk0W7/tKAd8GhLxWaFe0Xt61bx0MelWtKFJ7ILBrPeJd9S6y2MdZfkLdWphjPVcTxyeLE
j5d8pPlkLVOSgdmRQCvp8yJstfhtjxinWpbJbZRJXJWppfqlcBZUY7F1mxC8OXbui0gicdbXMxJw
ve69SpQFBRpzpzW67SJAjWSCYhdzP8NyaahZvdsrQ3/1PHJSjvsmiJlhs0Nsv3ab+xWtk4gtjhag
T66XC9W9Dt7zPygIwSbcYGiEZGallDswjXMpvx4UIrzVbAZbbK374/t29W6cgsTPxcjK5AWEmJFN
MT36o8b+M8y3f6CQrKm85felhcOEceAVus6uN+pRaSbqbMUfyCVk2VGcSUYZc+n3hn3EDhHjbsn2
JUiyH8TXKLUMZlxpkJI82+lgH6Y46tbumQfp6rxBP4synjLqxnmPEXVC/0yT7Fa8DlNIOAH2zaDq
booJcSS3H+kei2SkKU7wu87viEJVWlkmED27TSfHCHA3f4ODylBpDHIX4R15dGFSnC2ywgQy14Uw
RyROQcrHRmMPx4zs3j066WnTOYQpSp1DpYK4yyAhpcEbbh3W64Ke/3HmCB7rB5FOBTIdElUJCjG6
DONjyxM6GXjksgkx+jBIbuwm5V3StS4+rNHDf7se7jLgxAJDDf3Nc5yfSVQnpLI1aDCVR0zcS+an
wq6tIXKPgnJguIxDchiM9jEe77jf2Gr3u8QgysCuDEpjRcH5Egf3BXPR74NBRJbopwNVB6MuXjor
bY67C6IpaKDmqvHRPYfUW3cfYdsZnHP/HqxIl58QZNtmgihsyD1MEKWIrDsZlTRpvLEHCiXkKoxE
RaZE7zY8gxISlPOAh6MyqXgcftZNVKUKoV7x4PIWBKViJX2p4NTWr1JEWgIwOstZQIZyWas2IcNU
BINI/TnaFss2X+ddbBFB78BKqTQAXL+pE6VtViFzQnuCN9Sk6JjjAuE2222xMW1k8HnTx2LeHYeW
oKx/Povk5d6spB3NJMcYef0yrc3zp5PGwb9vfJ72a4r02AT5Tw2c3GivA90us0o3CB0Iq+8cJzIl
0CpZkeA31pyso8kpYL1L1lTuiKHAh8UNp9dr4EjtJtuTGFA6Mzk88IVZNnkVcVWCVQKNyG/sekf/
EVN9ssJlqIl80F4kKkS5gOrickNLIOhXTeQaxgNrPmwIVjOLUpHhEX08RANoLf0wNJM/aPoy9KAK
ZPyY1H88YYlwc/FFkCWAMeVQAM/oRoVggdLGY90W+JvRJ8SQqkg48o4diUrwK7Bd1/va5ENQ0X21
9ir8BbCOe14pqLgNKtMqLSP42OZrNgOWDMTIG+lhKB7UZdWXszi5FTK9lntTLX76rDQXX5J/+Bnr
k1AMr3wpHEvc+PMK32AWgg3GBBvTOxdS8JUMzilxYowyOUQfr75C9q8QXd6gyCPDtZNkXYPZw/pT
T4UZEDC7HKE6o84O78PZSpGeChlDv9H+8VcfxZ8SSuqEG7+Q7pGQH7J1wO2XTTqOJqc2Y7rWURG+
74eRWwhJk4QjPF6CDqaB77VYh9UlsjrFLwAAcCmTQkKeOJ88Zj9cgJoRL/6WFsTT1DGYmjK7ZHle
R04oNhBKUVPBaz3KRZgrXNdfi1losGJjqZNQOg+FO/kKxWpaNy+llEPyOW5OYOshE8tIGf+/Gkek
fxZd5sd5XF30Be5VnKm8/RNXNDHDvV0+vllJE+Gx+i1GH2rVKPzFY4+4OF9d7/6cJaFc3CZJaz7L
/D6+5Y/G72PIwE0Cj6Qf/FTToad7R/yEXGpyqthgaej2XzIlW7bVb4hSX6Hn7CM96DGBDFVl1wh1
z0fae7ywqDEiAxpCBdXXtHvAdoinack7+Y2oGCkQqlx59wdIQGPyqk1cx26XZmu43iwsqPY9/lc9
kcHrM9jmgmy31NyYiux1xld19w52w9/06R1H7jBquWhdqK3FdpCdVFmduy0WPaN6LqoiVhB9oZkf
QSrx5nBgHrUSBl7BsR8JUuqoJygeT3RcPf3gP2MbF1zVzrTA7xcRs+mzvmqi2WcuPQuM3s02KOQN
F2JrLoOgjP/nWtsv6rFvHVpJHELQyPY75PwCb/hz4gaq6YaUS58xfaC3MZJe5MHeVf6ld1qJHciM
PuTEbB0z2pznmBTiwE/XV86j5hD2XzkQbGMkxQLsyijZN8cCQ/o7oYUVPQFvgkweep1yrN0iaxTQ
8lT3iOwrp4M5ZDvMBEdmVKeWyT+irDe5s0thWvBSR2bki42Z+aYIE5snQ3ZDFSeM6Lu9TVs0VWk/
RuY7yBLQs+0/6SRT+OPse6jGKL9sX9HhhruZnVUitH+s12lv1tslBAJxv77C7GEaeBFGC871mm3M
Q7syHjUyoN9dhkYzY6/xh/Sw47CQJDwm8cBpBGpvLRW6bfg8/yjKDqlGzk2pLlyoy37W96h2CLxy
nEYyJPzDDXHDjicITe6geDLDxQomBHwEU3EeGRRk8IEeyi6JuOStT+wsAGXqozyefmVWo1qJW1uf
SnMV/jojbcsOXXF/Jpl8HNwM6oQ5jgxuv/oIolM3lvaDZir6w/ndFafBGoKe9D3W/UJmG+nO8Piy
ekiLq0h/v+H9zio7VRdBtVTRPMsUtcwoPBL/Z1N1DQtsh/1c8xS3PX4VMrwHFjC66xQMFNUbzwR1
Et9Qng9w/zYghEkzxKAfS4gxJhBJ4f77Z7maruWWEZ7bPHPPZK5tpjB29tLsSG8IlMteEIC2WM2O
mWb5NL2QVRcddg3xKpQrwFQCZEIeAwbyoWnOCID9n81aWJ1GQKvpdmaoRf7LUjm8VxJagxyNEI2p
WmeE71JddpS8O5jFux9+xADuIyGtJloDAhahmL2/R6t5RSwH+XeaXOT9a5UJhlbQ/JGH9+Tgtt5P
D0JRQfvZMODa53v6X++QZBpWmhpuuLC6kcNXnyPm3d7F6g+Z4rhI/dJePcyXB/lxBjlIOiBZQTVN
b/pDiVG1sO0v6C5Flef04IbE9BN3GMjQbtn5bvredF/3vLrY8/U6MH3VXcZoWZxAav8+6zGqyClk
QkHb271aCepG6E4LmvTl3AJcg3tQoChDFPogbB0V5CTUj6dvEdEExovSsdbDlgyBu2wLduJTe9Xp
JHlQI0UdFYPsq2HxDMSu5Q7QQk3piOreuP4eLM2BU1BRdHsEa+3i/sAwFl52UHq3B1ThK7Pjkhxt
sIyseWxsgmas9V3nx4/4Zfq2JausQyPgOsm3Uytf6pBs9Ej+IcpnX6vrsf5GslwON/nUz6rBdDsb
gJzOZsACiCfZIOVukpw8pt4pITZNgmc/X5k2ciOyr6PqDGB0RnO8RdcShCmogu4RlqrtfYxinGeZ
mUqp5d7ZOkClKKQ0d6lUV9IKF+KCzVExDVtBqUP4AWoSKVN4BqmW3bvvPhF/NMn7HWR7r6tFQIKZ
uUa7/UmitdkdSK8Q9gA2Ww6r/yIGIsj/1MKu0OiVTiAuhAwx7VcNttvrE4xOVR13DQt7HtcC8unw
nG9ExC8bNopexLX5oQU3Y8wlVx6MFo+opJV6FqBBx7VEH844L+cmfU74bumvceA7oiubEYw/+Cf0
T0T8sYSOttXMLoU7qgGpqHBvAJ3/Xlc+5A81J8BKhfhIKRarCVJCpT4w3HyP1LDueGhuAj7ZVk7W
WeGex1Nr2vEKvh9kFl/kmW7HYKuQBOkhZAqp+ER+QTegeGKbmr+n+AAFpVy0dWcxjcxu9SeQlXdN
8ud9mIrF5exJWyEnbVIIO7x3IXAfVopkbTQC9VIKCJdWAsGoXGK1XSdb4BraREyirhsAP28uoAFB
1hixcRgKs2lSJtpjCWICtsUOxfRBEKMNR59S1dimmvqNb0aZABBDWBNWWrmxbJa2268Lv9WGhL6J
OBrcV8GVypifUZAVV1xlQOVggt93l42HMW2XMleVttDJwWXBJfhO7ch3TbCk8wCF/6KzuHtWMIk6
dE7znFkw5SCvZSkBAKgDWG1f6Wer9cqZUC3J9+oXTpC8jSr1je0QrHdw/wCTp/60fnpQn16to0N/
bCuJvP5ZzayZPPS+GDzs9j7iJmkQoJhPhSK/rtyDLka+HfaKPnMtB+0h4XL+1EMqpW53aauEF5Qc
DV02xF06g1kyv5jYH/NlvmhPibv5PVdmKnAz9PHTqeyW+LgE7qlzxkcBk2FLKWqMSnDiepG7rX93
SzDU3sRuwnBTa864DcRwIwW04KKPXxEmoTg1IU4Q8SumTImtcm1Mph+NOM1RY2u73Pb0d34xXpg8
GvtNMxiraKOHfAh9mAh4hvGvW16Brt6Lzml7393u3slF6U6tPq+Ae8AbTpUDOzj50lu4PtDmCMK6
P2AMAhgVPdi7lYO/dapGSWnw3LC6mVLXBqY5dlKYjYQBIozu9SBXHQwHekQUYsI1GP6Xb/xpBgu2
8p0VS2H68z4xL4adqgYdWdLgtoow3qm2H9ViqLXRpdqaU6wq6xd4F4bgoJgsNqxqjz5Vi1nBsJuV
4eoWRpZkLx7RS1zqZ4LeN1wUP0d1ynNdXpwtg2soiGIEr4d/Wmoe6cjLcHizdPOPDbC+rK7By4/M
aC9PE3KDlDNVGaVFhcNOtpUBo5eC2gB3deBpkFxcOBh9rnbSg4vgSj+5KnNpBqiwUgMUr2hxXXOa
kRBRQ2zBUnrfoAZFuar6SlWlsBK+Ksorv2OBTlWfd+j17fk7WaWEXwBVSa/I5LeFNapjV8ccRMwH
Uv/aKP70sLMUi2U1tc9a+FVkaotnYQ3EphkQqjKpeDnQWM56qMRugQRhgOai4mrcyxxtU64wZzSx
wrPH9jMUntoI0O37fLJCl+6SHpEyGHeIj42docTGsaPbaJHhOb0ByThFGq5hJHClqdAixNZNAdzA
Utq9MBX41faM8JHzvDWG0v0othCSHh+jYillFhPn9Cq2tvw7wHJCp5DRDxzCQAuFStynJIs3C6W3
v9aOQySnIMRjsBHveX+cRG/2X/jl+aPvUDMm0LPTlelfuqb6CmACtOx3XVd2HwPLHNUBursnbAbp
piR1T+XpmcqRXD4UjT1K2qPuLPu0CuaZA2glM/Of/lecbSIUTaUhMZmSdxENDrfxeBzuVWJae3lV
FzP/8gSof80M2lF0iKML8d3Fkiqsd9Z2+REID70bVc0n04Lj4EHSl8wPBA+ycMt6UJah9JxHnZNn
K3MqNXm9lkCoFf/bO8UiYx0qi7/RIVNJLJJe7e1d12w79GGxmZqReMq4Ty1rDXarQ21uWyL1o/bt
ZPK5Hk4JrjkBmfqly9lEMzJGwMlGrv9NJ9CAf+26+t7c9kQRX0kltqTarHxg7+Gb7ImNi5ALqFDo
SdVQmF/r4xHaC7V9lo8sy94w1Hhvbt5lk+E20dvenuzdv39E57BG9Us7RCF1wq6BCOW66ngTXmlY
vAVjH2NZbNemcbOYOergB9PDxL+XFXWLRSdMDFvtR76qFBLk5FxUo6KFq4qIl0oRRZcwso4jhpz4
4fEGHOKYO4p3YNdps2/0mDo2k/6FzJbEhImI3/g/rpKTxFGHtgPi3FZfm58Y4ay9x+J/qrnuFpgP
lR59jSEscaogGiZvnEfEuNRP4+bulDqHTCI5+IgPi8yJAdsTNM7VDKnMoSkF5UFsZzyFunp8pCgD
TsoEAJn2BSPbHbisl0be+44qXqoAoZwtAtuIrCRtTAzWmTIB+dDAQc37LAKAsxYL1xgFbhl+3MnS
sQDbEW4r6vORdVQEcNdcJvnMkY2hx4TUA6X/6EOIVu5gsN6LkxQE01MQBKH5IRfDkaqoyKFlhc6t
2B6ugQM0ykPRRPVabtL9JKG5MJCwRWPthbqUmUY1fpK6oYfXbxDmT/d3T+5yMHrqYYLXzX10xvaE
c28wDmcntjCYDTArsRpFyct7XdbSrjCmsCwoavd+iS/m1WYe6sfZ1i89YVFhNUJg/lWajig0SCWO
Nf/Cn9MIy8wF8fCaywcRKC0MhMLCjkk91ykBW0iGgMh8ejI34oN74wQWYe08GRQFGtWXI3caWaF7
sSyES2LP0h04IroZZStBEtjNzkq1v5MGmj1h2Qp/ou7yOYYbxXuQYhPXqAnwgPqaJP3r/zyMrLob
lo+Eq1mTZ9thRpOaSof+mEHJN41VPa8QuQgBXPpxSGNMJRmcRSS8MRkRI2DtOe89Lg2+oMop+itH
fs8wowIXqMo41kNUFcCG8M1xVfk2e0ixIT2C26lAxT/VeL/DhLnAEzUn+YBuxMhyok3y0zrHL4+q
uHmBundNApehDF9xS59tMK8HQIywYXFAyRcZPCHa7UMonbbqUVdxCzSt47FkVtaOOJEUMBSZC3JD
oHbeeX92/dUnh4ktGFIU2Yn3hdJrZBKwcYBVHGekumRU/ToCk9YlFxJDAvkkE+GJ6LDas33ZgalM
a4MoRAq2Tlgs4yFT5DprzNWPsDxEs2MAIRTDvQFP+10n8IPE/TkCT5SMchOSA5VlLIQDnELy0DXq
HL6hmRxl24DnkzOoY/ylYOPUmAE5FdMg4pdaIpcrokS+66r2S68mB8e5JUuN1xf9B8azMMyYVW4w
1YzRxOk7LG0BSLjZk0+LwPdJAF0GDBO/dpOKlUx+y9OFGL1zBaHdRCGlblOmSkQugVSHHWrjuGyI
3hHIhyzAnt1EqFhyISNtaUqUw+iNia9K3IgQkMDUDDxlEazcp7PdpIWsQ6ue+/lOk7g4v5J9TGpe
eRz/ne41jr0dcKq5iG2Y+lUScXsJ+OZQNannlDbESEpOpf1QX/57jAnP/42XNcTBoyPItXe+yJS+
GAOiPM8bIelb/+yDULCXmpn6JQXspz8eC+iYNYFaw3sE2qQl2C0C/odynRGnb0wmeu2IHKD+uk8H
aIccc5GCQPp1Jv6Y3IAEKQZDcbRGgTedKr/O18uGfm74yC97OUWQ3GmYBWIGJn6DtK8KPahtqBxf
4mVxoeKbDTxw1rj1bXk5rQNtbQA+kBJ8yofMhTTAadWwh8Hi6KbCugPHORBJ1KsiGvNcHhZOEjot
opcFWVp7qd9ENQeLQHxzxnGgX55RiIKwKBqnWaaO/VVPRDODXdSB7FDNiYsCHDPmsdzgt6W0mhB2
4NJ4vMuckG0+z5Adh255y/9zIBoaMgoIT0VAzv9OSJYFM0ri0K5lBQXnXhgSSVq+6+XavmZrWUVv
kp9hhstSS+nmIX+LMt/sbRoeH7FDAFg8Peog6sraJzewxxjuwP4WLbUm52LfUhTwKvbMW1lQPcfa
jREyJfQG666rI5rpViv3tDQVs/gZPczcjWiXsVCyKVLS0LKHD7hWWXmE5mWqNluVf5SDjnHQ3Peh
aLc/xd3lmXfgb1uLwTaSK99wW/QeQSs+BLYamm5oogGlpfBYbBXhkdUw0J2FAo0xdhAU/fRoddk/
COlYFPjL1I1QR7oFPViATmVMmt0N68EkquzaOzb1F8T1k3wD+pFYOJOUgS41pX9BJLCmCqnLpU1W
67NAOoWd8BmC0W4K7a+TwGDhjVC68jrESFm6b6CHe2hH4xJtc3x415o2rKDTs45VMXfjoUfbj4Jz
8uuY5XiFu+1pxqzmKo6XLs7SnMkUI+NJmbUJpiXQnJlRJFWtQrYfXbb7cPheYjLc4KI0yXBmWPMy
TsgHWJbNuSDa/qu0JQjJyQh+/6dCH4EJlphPGlqlaJAiMmAkMqUeSOGrSgyb1LcYb+yF/0RXOnXz
gxeoGR4sP2V9vdJDRNMBj6ROf8SIeoJbW4F/Fj0y6SIftpvQfrETv9ixJ4b+OZtbXtvsx5PsBlaB
nIQaYMQTNLDFvR8bq/SmFZWKGFCfYGY531TX2E8YGphtHDmNQ0rklLRim8UoaFhPrRqr3ZvThgq1
UDDPD2Hf/4wfx4cv7QYMI1V8df3MPztA7+opk7uOqqvSGf6gO7T7wQuACzbjtTsfqebgrEDjHgFD
ZbJRiiJAc+VmmLVslqqZLMxRg3wj8LOaKRq8Tz2Z2t4U9ziKbuLaAxz1LwVAcvKgNTlBT4rVYyrn
BYgD4CRqJJyWpueXb1sUJLNKZ3ar87YWle3SCpH8swPBbYhI86YQ364Fg3g3Pz1ZpIaiwO7qN9Tk
rUQPGPlNLyILldg0yd83dYiOzY7OBcT2voTY9FZqCih+qydkzso3fQ2OxmckVUXaNvU0nX7dojlP
UqzK4qvtt8lksccFg7pcsSDFyiyOtql7DsFdc+cqJ3goR2pOQ4KwRqXk653piRxMp++IwZbboi3Z
ffu+S8JZifSPPwdqZmuDo0sdQVCnAeoYobR9ybTEACq3Rz8UGMjMiQ8i5OyscdL7b0XHtLMLxf8Q
OKuXVzvDBZ6yqU22g4C0mvZVseKTRyhRC31mM7jnknEOFtH6gV6//bVcr14OvOzdDnht4l6MQKXe
/RaY28nAZi8pWEfVBgxIou0FSFV3FjsPInxGvJpgDOibkewLGuR+qdpzEleH9hnKOacIcgAy2n5T
aCcRNlQRGCfU7hQqPoRAGXT4aC2IcEzKM6lyZcMBJgQNrDjU8o6/SIcxds6qqZHNbZ6Ffwk4q8kI
ZJPUk4AQhXHnVfw+0H4P95yRdP9GKH1SKsw8vGxa9KfWWlQtHQ9soFnhFXTkNm5SfRW9tfAJ+DUt
daYGcIjSS8I0SalFRnJxgZAsPNHXxSuvGSTrFUwybe2SyT4TyInH6s5AzbSk3odAZ7GfAm5dEtgQ
MsMHojSdmeWaOEDug2lIyvsPChY8V23DXrbil9s7Zme+GcOYnYWaToAVF8kTRDuq8lqXvA/GBkOR
UHaDgVZOEYcR1accUBK8psgYxPW6y8mWBu8tuqieS2QqH88r81CWgwk0648ek1xbqu04arI5rGBX
iYRFkCgMPjIeN6sYS7zrqQPqgL6vj3UAH6/rb98Nn2CLdNEkW4TPH3+PDHQE3Fb6ItqhfEWOsjGI
70VdLrCYcnlMGnDbK7ENx3dTbjjlghmMhlmocj5U6drZwZgJpmIVOHcHu1EcJD8Rf5JbJBYxw6YW
89kevEb+NiVt3u7p9gSTMXnxg/0+a6LrVUJOoT6wMqi+IlNkO6fdPS91pfgIiZpKSjjLy49A3J/m
9IuY5GCp7JvGfyaO8AgX30yxGFln5lKDdX264lTg3b1OHeyxQ/f3OqYH7+F4GO5YscHLh7vMKaX+
BnFVE+6qDSSW6sZ34Czoxk/0gKgxXIAH/NEyuve1tK92YqjR65f4u0UJKkmGlSerGtipS/l0GKq1
XVSw+Z0nw/V5N6TvWXMzTVLftc1ssn4KIWyG/IflPe6dX3goDDM5lQZp8zTt20dXbDh3/XcJ0BAJ
YzfNv8HwtUdVHgYzPb5XNLS0iEL2pJS9i6aKZoknW8am2VBGzZANOfexMmSR/IMAiczlgOHRB8QZ
tj1jYymC4v2d/+tqcOa3xUTNtCFFVlbQlyyT0cuMvbjnFA426v3szazCZyH7q4lOc/JnLSS12oee
6k9b4DTFH6RuRhulj+4wqOFfm85MlFyXjQwaXhf/V3lfUJu+iPNYea8oMX/uRP59ZxFO096peU7W
qRZ5vswobcyLwAv9WT5bHUEE0k9TM9Z11+DdhmCwy1ZGodQ5RSUAb9+sJs2vKm4bxpHSPn1k72v4
JtXIN24Z1fFKYJnuVf4yp1VerDH78/YKfwyolwzhkHFfuTL569uXQG+XDZrpKNZFjQMPHIg8sUEk
Y3DA8wHt/dWKHXwHBquCtrK+/vStPwn+yU4dU3hUFc4WCQ6uEtTRlMpl++N+NeL2GW9eJx0Osc/1
al7Ue1r5Vc9C26EXpuVRtZDo4pajwsNwNNKG9p/0Iq5J30x2BKbrimYs9rmsRx/LJSCcMQNp2pQG
7zRMpwULRB7e89aeV8evUSonswc9K06AaUI1dkFDx1V06gxbJ7IFpnabU2xaZjWdfTh3ndPMbQx/
UImc2QpLG5tdqv1I900OugcXMW+Lg/SWecwTphPbGV/Y2ecP0ycIZcavM4EGakMaDUApyNELtHM6
fB+oqIz0YP1OqdVE6uNyxPDjDZaGwG/YLSpA/Z+tU45atAhpXfkPNg88pTl9pv0H7iORJmqR3b4U
TtS2rNYHHDR+sQAfojighXm/qi1g7gfCz5FJbV0WoxEMtPZpzreiw0ToouLVKiMC3ch6xeNs064K
VGT6rul4f0KxCD1vxtGu2XjU3M43aKoE4XSs7aMvyvDDOMkACD8kW2AHsEzNa77LaKpuoTjZ+qvq
o0ulLemv2AROQFGGR6JgYggm17Mj6y3CHYmrJNCVu+uCb9HLwFgrTlqHd1aeHW0hlRHfW/EksZCG
Aux3rvfPRdiMbSzNtEh+8qzvbaySshvOWds2eS41t6EpCw3sITahWv83PpziKimGpClkkGd1+AvS
yfVFWxYHW2fStoxlNX6xJ8olUegxfLu9PEvlk6viDGVWenlRSb9UiPTh6gpH986AkmONDz/KGYRX
ByuR6pNh+Kop+0LMfu2PdnQj0UVwJvErjVfGMcVZMZUf0T2sKQXRG3vZ3Y8US9eAawD/PlJv+aKb
+o8D4ezwAT/gsS0HPX7STt85+ZoLzdxR4kKl+VA7GiFIrnuq/LZeTi3Xx+Tziw/T88NaCrVXyaDf
DyymCrn/Dj48uURJzGIHKMzxYuTTFH8sX5p6FHvzm1aEOkSPmpRtTH2rpgeCMg9fIP72hADzMOG7
3xKk+XToTIxcVZhRawFaPBBPwgEkZEdRUv055XoYMSBzQO4FVyXoUwt/ZHkxmNP59NXB8QzFeev+
/oaZaDtfcBh6SfiNYSq/gAspJ0NWnXhxOWDvOGEY2qp7JBbcFsok2zZr0H2zcpm50TUGUnWOVbQa
Xv0rPjo5yjCuPvBW/PaNjjKQZDdKh7lEdy0TxDS1033QG0o+2ct+K/+MiPZMT8PuZ4XtBI99VKI5
Wxv91TLRlSeP2QvFofbcZn4l1uZpFRqzCKibCppBmXZBadB0AbwmH6clKkq0XAr4q9eg1/ZnoMWw
QNR77uaPP/s0FusacmZDdPeJSAACk+M+yTo4FjZLtUlEZDfgy89Fz6JFgEg6Y2Z20Vu01pKL9rhk
8dYDWEwMYdOBn+jVrKnLfu5Muy7zq9rdXkf7ix1mD3VZo23v1ZvA/L0C0JUgnGeSJQh/1DFOhJzJ
AWUpwDHVeMRL6MnnMNMb0AY//8IIrgZ0PYpBLhGSHnSXgbrnKmxUK8s9uPawTlOdj7ClQ6jT2tpr
AKSbVYfkrsxaOBzR2z76R+XBUSx27Hzk57f0HUMuA59RRUN1ICw7vsKzo9FFR8AxTqxHiWVOuzJL
yiYJgoVXup5VHle+SdRDDGIQ91N7Nu/MbIlu3PI+1rQuVkYgqaC1cPcguhFDa/sfvG4BnSqznODk
3fSqo3yNkDc3gDqvpoKfwFcPk4XS+7Z7fJNq4rUWCMpQh1N3vQM65Hc3Ex7bAONXuNrSV5zWDpJM
3TEEwloWg7EaXHMKrFHpIC8RAEjo6v+H+GNXSAHQCOl+GQwPMdKY08on7SQ0RCMY7vAKb3VftWva
JBLtQpA1qCUN8Zo00FNuHrP30QNQB7SISWx9CO0Ov9MzkV4EeEU9xOPGrrgR2GZ23xeif4GRu4Ci
ZyRS1dF92DCrP91Yrg3cEPrhejNoOvCfzLAi9Fyhl6j3vEHBuFhukgW/YcTsS9NQvNhldvd/yt7H
zb45jOVex+sRYN81qZolZOKiR42gdKhC61GIERLiX1bte1noENMSb/SBaN8VwSnXfsH/xqfQCDR/
N4JIZ4JS+YUrCBaC6vCYxWDiXahmnwYBcGS9PGBUXcA7zkiy7AptEIhRT5EdU82GvpY/ltpBwEVm
PLawO+zojOYmU2VpeGq6wVLJug8MJA219J072vStErxfXXbv/CxYOWDLXkhDDVeoaq7h/BSFmOrX
z9x9eGtgRQCfznYgjoSJECooy6I/HAxee1f6cngitmDe6H9m7fskZex4X5Bw7Ks4cbbfasYPP+nF
/xWFec8fc+2z3koh+iieHYmQzKy4TgXPG2QTmh5zqIfbVNqmXnoaiaxoKxzWz6Ms9SSjhzwDmXih
etcdNN6BK45TY5SGJWngsSEaWx93H8jiqlUgbQdd27ziuoZLn0OKjQSmmEos0D3w5c3E08Fl75Vc
9fFrj8TempdEqbO+q+urEkapYHPZ9Yy3SLHUhgHyBOjZYiTTMBCovHyBQPv6jxODbJhxCxSaAGEJ
H4I1sE3AT84jwhq5xrWJnltyLDKKRHNxLXKumw8lppHYK312zn+HiQdDLtbEFA2e5PUc01KRR424
DMFeUYdHaD6VdgDrDqFCjFQB06AKrTT+Iylayg4Kp1qXyGvYEwwcTrqYgIzai2dx6sUkaRSBDBmm
pTZb3kreKvrqjj0hWRB0c+vdibJsxztypkcHKFz4IproTRZkAsVYUUB6TSL4/FsiZHYZib7hQGte
nayziXqtlexJPv6xLHjnPcgZPdr6Vmx3t90LRD/pO6gFomvr2PrcFxTHd+Fdm7Wr6vdft7BOepog
07bARW3FPFBWSLGGw2GccJy73TwjSc4lrIhCxliUL0dGmq0SziucbCSgsBF9wvR7DMmCkcn9AdiF
E9cxDWyXEmJDJu/Wu1tFFq3S/ue/7Ih3WvFBxmkCa5SiDvOQJgCXJ0rK+ZsUb+5ebL+cz91Ecj5I
Swlqjb8sCAMljGWS1ORo2Bhj/Rozu4TlZJ9Y89FDNmRsXOfiV89W/UcaEme4bOx4iDvtU0eUvjsz
K10YgRWkmnkw4Ynk3c7Tb0viIuoqB/aUZfXAQSim1yNYrsrYwOFFZfLYSZ4irRh2be11OyMqLqIY
FCzQqyQQPEiLUD3CVK1Wz7e4Yz1QmBqt/FeRuUVvdJzFU/Ea2KMkFMrhKRnz1bXxTEUqGpQKOW4e
j+F0cxixT2qR8VDfhU0hzDyNG6EYwI2ZpSzdR4APLDbJfhGtDC23bl/uP1UWaBEbY8zbM0FWTMYR
XbT65IT/MmYAbo2FgF6pETZ3coeVcpj8tIFMTiaeupAkWeEB4PwKXW9QTwBiccK0hZJD4HXI+O+d
MAhvadvJU0VsuCZNlpQqyNOJ/RmtwMN4DpZ97thEdllJTloNPHSWKwBOLWmRPINRw3ZmW4HLuwjx
u4yeO1ahwoz8zbwms0G7HcYUN/D0mhJ1kDm8keSfGoSO9Dqv73nWn5FMXVFZWMa2MUfGCYrmwm/K
d/4s6ivtlvX8yWI+/GDuw/xwWi5aqBWCB1EYIwum7socfjfc0FkL9J2gKGi9rmrTYb9imFpBeZPI
WX+jG3wU35I53nMyPOEHE1kH9OGrSHd/vhf1Od4A82gd/b8isTLcCuUriTJyVbeCuUxOE9j7dmOw
XD+lJ7VJQLm86MMKXvn03fJJnPQ771bvUuKKafs4+DfRgwdZHi0N/2s4yEWUgBaviVrFJDJ50f/b
RFTsawR5V1I94xLJPlDGJbIEiFdgX2g23OAIzDbv8WnBBHk+bTXyQHI7kcx6JAuFng/0cqP11kyF
CCpnsclBp96EjhgXfktWgEYfP3zru48HTECK0ZYyJKq7SG6oXefzS6zoFsQxRoxrmr/yLmWC59kR
D+xagNBB922H69K6zEWeGFqxAalm2p+LZLvhUmPHnI3bkNktsocjIisWUDkIoZrpq1g3R8uYcdl+
j7pqDseygvTrBkWA0JDaqH7iJau10mFPGil5bKG1iGJmv0MZse60oYIlvJFR4e9il7wl5wGBWnNQ
zcR4mSZMEYE5ZHbB1FzK+3rawXFSgCjmQVKyqkGdxy1m/VQWmwRB3fP7bjft+MIXh2OxlUnnubV4
Zd5v/mzLNUBlTJvw4abMjOPsUjhwvIS6o9LUGTG62J9xep9L7eZFBhulLVLrUQzFGVatJwUcO7iz
qoPv++DYcOw2Fi2fREEiS2BgJxs5XIteonxOkAU134rCouiT114lkD4cKY5rBMzbkjqA2vWW+nCO
StQu/KnPbKSCVGIO5purVeZvPuHv6NOqMWm4TkPL1qQNo21o3v/qXdu/QMFQp6zksGL0bztc2RiE
CVFLBnKHzVhcDAHzHCO/xyauOIwOahnaOJJcHpxamusxJy6+ANuRvZIXybumwuQJVdiKUy8btNfs
Bx8ajKvlZjkMmQQtxH8TetNsQYyxuCpCx0q83414PqmWPrciDT1g2WVm7nTm4iHdmxQ/KIGupY5u
5GdpatTe1sF/qAkqnT10B5H2r95fZI7rDcMVstSDdyiGA5RfuvrlnNdMBl8b/Z5IDzQfO9mLDDJj
H6aEwjTP4W9JVjm1H0hTe0J1n+/QOnTwXw7eLKhSzXxdPLlAN069vUyrlK9RV5NBKOPV+SX40xGL
rZ5zcsEqH0fqk+8zDrSgeRQlRM+ZjdfJU+xKGfSfNL86eJADCTq5L2TwA7Uf/7+QcBzoxSf11rc/
qECLyC6x9u5Zzu84xXlC1ISUytBMin3gm47MHoFdfTYWAjZbzlEFGzvgrundHtK/dNKSjiMIS/9A
kHCIArtmwznG3Q6BzlLGbUP1HpnCRGcWgiTZd7RvaRURtUNQA9hGvkyL2d4w3Fp6oo94mLZLEbet
s0tCL93qGlr6YervoNezsT/Iy/v6fY0x1HnOFFKgTgUarRi6kysoen3/KoDYM7vAFfaOm4lrIC4v
2CjiGE5RAg3idCSv2WWJmi40rHxjrgOa+4L8EOnaYYMwoLgp+gosw63WN+/Emf6EbeM4sseF0yze
q3qkG0fBjp67KnYLfqXZQV8HEEhYDJeMCtbZtTfX0ziSNdXAlfd/70HTSwsllUUkae5yfNhue18j
KOSyKDNeApuqyGNCbGKyx42ERCzMNI/jIFz1gwzpojZ4TZPMu/pHtLk79gJ1rF/dgl6ieOriZOgY
0p3ShGqNnSCfPNwzgj8RmFLXANGatEZZM8LS2KpJL+zbrnmGVHXnB8B8vDzWSFJ7VogsjeqMNior
mHFOpCDuOhN9xe5gUuKqn2JGxDm9G/EiQWHQHUeGEC2GLUTeWaw/PtAsN5k5cmyQTGJfFcszXDaR
eLGqge+kcO4lYGu5BqxbFX0h7WGd2VNtHsURNrZjXAvCsUJY+QTdROQfwp4RcQ9bhTNvJ2qY6MLj
3bpFZ6hIy4r91U2kS+MiVW70q9wwlroCBLOVcIXGfCuxQsaXA9EaMEfq0zncS+Vn43qxa+OTl2tT
lCi0C4wdedkUz5RoKxOXddlmNbHL5L/EiFiYIz86mZpbnMwnH3df4pvGx0eQ6CUz4zt9A1zOVRW+
BVgJlKOAHC6/CeN7aolxJ04Y4yPQ9SxaHRBuT1xsFBCrSFjxq+eFf9Zm7RUwSHU8mIIqa+E9rHeJ
o5ma/9AKN/aFikqnh4WWDpd+dPTKW1WDTqJo+yPtjLtxJfOHRdmQZ/yM+3FUIp5gTUA10U2IFeH9
piIdr0JsdC60SK3KVA8ToE+7EqVvrRZ/3fe1S7GmMUnFfBKcOZS28a+V0DAeQofAF82hXqftnpBU
/IXGkupu6QVAG8MBGHx9G/+zSGuypPFpEUdO65DfTI0yrt4gp8WxYiYy7rXp8x6OOxUHW7NeMasj
MaswTJuzihwN96LBmhLaYJ+0TouIHeWzDPPTvdOT5gwHz8VzJu20U9FQmfwaWblMPWKeEejXObZk
8qr3FcRLq9QaVUgQCHfnn4BAAMZghO/zGAklSnSreeB68/GOZ6i2WXmvUFaIuENLHn1RSfGqH2z+
n06mwpjc+v8k0IwaZbyOj0rpXrg7qjzKUjedegVe/3v8/8mxFNqm25VGOOZXFC8bg5o4pmxDkHaU
H8CnRiAhxa9dZ19awM91+QXkTL2FtYmplo0J4MsD451mj72vX2N2RUALWBxeJ1bUm4wYcTVWzX5Z
ldiK8mgftERi4DocYvBEf/X0D3/k/7pdDESpyvZg2xoTs6UmokLkCRzb1IOA6EZ81r1OT5IuZ70L
iwdW/S1x+WNekoh5nKEzqEVITmtbFFoeMYyGQMqyCtrNnYeWaPf1XaHXm7Z5xYiIlIqF4ZQBWn1I
hYHDKuIGanuD/TuVDQWqOEwdmy/N9q0LftvQq42esq9vT1hl4RIGFkAUDZUUfFlV3cp78eFGHFcS
hl/QCenj+KH0X6F577PrxJ90x+hThdbjYRNpMgvmGfwFaiyFOcXUfwgn4L5afsjIVbpIu3fkDS/l
xukbdZqdUFx3vgfm2rrBCv6ey3Prvpvp626t3BedUjX3B9G0ULZNbE5w5MevX2K5MMJK049J0lBG
J6fF0H100QlCuJ+JEbepKuMlbBWSQUsqHyUoZcsv9wKCEi8A4x0P0nHQ4TngtTYcyWbIUoHPBM8l
35WJlo5PrrOG7W/xJKZ7VlVRtsju31lU2CplqZU5tvfHQ7hCc6SoeJyW2PVL8UTdUek+SHd9KWhH
z0vAlWkXbfqGmtupa6HWtMPxPGG/Ncqc/JStQiZxJ2m5BGAyzTMQGe3JwCLAog1y11tlMKYL2Y81
nt8RJvp3YQ2mYfMs5vxGayzBx8poR4JRl3Do62tagxSDqQEHlpcvs9sONuyQ7lVJPH5Lwi/Utfnb
VgcyMcz+I0ByFb57xJVrpAnA6O2WMgruYXioZSvZNUNjFiCFt30xtGDnIqb6JpwL1YohuPXejLui
wGV/94ysAtY2yI8gvljy1RcryqbhS6Ni93HITnvHK06bSpdJri4V2YPRDvgtUzKrTUYmg4kE3TNz
4Ja0l36wfe7ohUbwVVq6OJm32KHrtVci44dlH14UZodskumVHAtd8Dv7gGE5s9kMfa2Sh+XaXZjM
3k20ZCw6B8CclOOm+QwRfu1ynsEI6gyA6lvYmDu/kbdkY2iQ1vDsn+TUr9rI6xc9ZRsswWbAx26G
oVkqdLDg7kDjIWbXKQ7C/2/8pw3cnUjKLOJ6bqrIk86n1hXLHtN1csxvlfzNG0Q8KBYArFkALIpK
DvezaV3DOj8CTfWPE7FVZHuhMOwFRsB58aSkK5FcikrM1Up3bvKqxuI5FQCnlDpzqiYysgy6Jzam
jr0IITvqLU7nAv9QFkZw+Kw/hmck1P8WXvBCqtaGtRV29Wf0MRin4Mwz5fa+W262zsAGpJf5twRq
PRQwyStcF6/vCeQHT85hBIamee3ExcvDpZeTkx1T0s7+VwRAkmoqi97XAqjEvN3mEc20IjH8NFWw
wHOsNadnOAlmaMzhfRZgtqe+Pl3tZ3aO++KYjm7E1EJbKIXE2UJ+uuvIxHwlHnURlQluUEt+JzGA
IWCP3ahL/eJcuY+0GGX3+IMqueS75CZgyl3i8WZw8nZ3tn33EF4qPaOqQ7+zDGdv5OtXGweZhoAk
jM9LheB6ZgfISTnIXnAOoGAUjmgMwWhhpFnriWIAt515lH31/6VuFg22fE72Kghp6/q9qWv2rfHR
WSmwqJMxNaqjYE/A1cpIROfxmfHW6o1edfo0iMmlPBgJoQpJh4R6dMB+12NKNGtiJbBAuamOoC1z
usoA07bvSzfMJVOnljK3m07OHqOm+TnGn9+9IxBD9YXATyV3xsHgqToGZFgtXCGHW9W3zWfn4n1c
na3ZgFPFAM75uOLpsZFJtm7LLvBzVofiq55KlxdKVF8mH34b6TPkYVtq9vzSH8wkTRT9O/HKNVt9
neKlc9JNEvkfisW7NXxeOJ2h7wo7f33bU7liJn3JDa5W8JUtA2n4mDru0ifzdFlxUwrteBmAQgWw
5AiNFMWCVtTMOfxZ8io1zEnLkzFJJahRnIrQhxA5wgT+u6vC2fevqTkU9xzUTaLzHrD29ipYBeLr
4VXLBcbtKaZcERt2vias2A/n6dvgVsZNLAW95wcZRNhWej4T3tzg/wtqyP70T140Q/KdzRadOdJW
ju+OCOuufb2z8LnbGlLRsdM0PBzjTencSaMWCcijPTiCdQpAPXO0yVUU5ZZhhnSkL59DMwNInZ/i
7FqAireGQ8HBUod/Y+GzbzTRSSYh68uja+SZUTfFx9KMZhkUh2OWo/Qu0Gry8jyPqfSbFCcX8Gho
GvvqllA6xfIUU1ruTYI0p6fV8b1hxIbDU/ePcTKBWhZ96eqqSTREOVBh7kccZakiUKkSBHz+4cD7
PNdCcCIbY1VGdXSY5VFfY+dPaXq+QqD2f2QthxTYjJRyUreBDhsG1dvIRGBb8h3RKb6GEz3eCZ7v
Bdnf4etPVBezELNaccg75jGCuZcsQy0rXF/JWzHmy6cm+ub0Iv6jWVTlhFWQM6oKLf/Uc83+a74l
s1tYeou+yYwdcgmCuQD9LgYxtOV6X3hrKPTA0D3Efc0F1iy/IuOSaCprMvRZ9I8R8202mlaKzdom
TwfAsDAQ01XjJJEP/WMKAXTotV7JpkQMbzhLvdvpO2Nh086CpS9ZqyR2knfuT4C2/DAhh9k3JfxE
NShj4KSAzqAqk/cQgiIYPjmYzGj57wrgsN2MQdLc8RyymNOCakOzsZmtt6iPdzTfC44M0iTFzHCf
BHdNGlvjQQq8HPQpzUxBjhG2iNFAPSwxjWDz6xkw1gcbi1ClBGOg6yy1N2mTg3aj7mWwA/+rcB2O
94iFZmwUG/O2Sn7N+iZpVtTgcXKWAzECbCixVPQH3XcxQTV0YS+8+S93B6V/Qbk8VlopGxl+uIIB
Cm0BMPjpQdc1ujwte0QGnZ6fcYmkp9DQoQv5wccbuQTWwHlMesWz7DXsRVWmaMRKs0neHajIyWqJ
Lq0XDtEdq9bztEEGcVv3Hop+ZFpwFhVikmOoB1uACrSQFa0lmI1Aal5X/khBP4+7pN4PIO2Mfxs5
9qycELIeafZFeB1eea4FsTN7a0tm2BCTnpy2405ItkYTpDFy2//mBf53ED22Hw5UCOkX0tAE1lFi
8Mj3BpZbQZv427e0sWboQN3TwTdQsqQYXcfU1bZhffkm3ZUm/0eFQGxKgrfB7Wh24RhEEJXh531I
OJuWh7HWzBdQK14EaobKmIybFV7sSrWyPK6snuAGTcozBRrAmlJbgTRL5AZds4xLhuCLmCr6NtC5
5WvUH5fmhowWDpxxZDhiMXwRFMmgO1AnY9JsrG0SoWAmiDrzhaQtpmmbBcn+lJ/xbrUXnwfwiU9m
dz3QlvYyRHEzWkXyjx5efC78LstJ6fob5EAs+GfXJspD5uaiDHuzGsZJ0PruYd6+sSz1Msxtq/ba
EXVF/4VAjB8QEC71XL2xOnrN6smgh+goMItrhKh0SU0nmkctAmvc7DXGgmHVWv/iPS7io/OqW7sF
YFaqhR7b9k3OgQDJHKKDJDNu2Eeu6Xxa19ZG+EBkzfHPThG0u1Lq2HOR2BkDuE0UDwdIRHcX3mIn
amo+23ArsMjbqbrr+667WOlF4pO0I0/26KaLx6UDq42WqN8tylHm2KW1Q3jpzbJEVVYsY6MO0nxl
S6EHvai8CFZ6S/dL7t/4lMUmJLv5PepUxDlJw1cFvF6zlHZCNtdleBOImxTU5jSK+Vz+oQZS8QcZ
DNBwZarzh6qh+JKA4jia+w6UOjvVrl1ZdCBdrj9hU+wKnszCCuiG03bbjv9Rh5X60CLLvd9v0/8B
QNenBXmCuspnprsAmZOic+JxKsO9io2OSycsdrtHRutjTxG4qeqrZeQyjfwytIV0EUvjHWuMp6wh
wzwgn0xhWjnuE5IY6ktlkBahv2jH86EsoqCQUJqf5Rq62/rqUjVOV1iI2dyJhX7Yrv7oz00cHc5I
oKvWpzycQkOi+sIH4WH701hK8VsjiDBwh2AdmMFPQpI9nsMbjYZAKvx7XAY/4wYxk76h1ja3G0u8
j8knj6X03lRrkN1cE2CcHp4Kmm/tyrtJ/wDt8DvMHKeK7MStHZzP4FlDu5pa9kVzOnXU/knBHySC
4Xz7prA/4JwBVT339kfCTDyd0w/IMTb7rMFjI9RVvGyW+/9wvrKV+fmgLhpJxGNmh1ta+LTcIjnh
I2L5RkbzKpzuFUn6qPHS7sQe0DcX2UZFQDou/LaMo2UnjRDfK5JxJv9WgyQYXyNRmOEmhiNyMzss
modfDLL1Sbm0lVD7aaOpXySi0Qgf+uCgWAaSHRHMCcATQu+6InDJCNFc0N4TG9RVrXyJeDYStOde
uSfWPyC/5WuWHGUKTIHM7XfBNfyIvFGz6qCJiNoW8KXkmCTih1jL4AkfD8CykOfFfeCxBUafgICs
Ed+DHXTfmHcJ42C6hOkrr+xSP3aAkjXm1O2mm5q6rotnRRJ2GxUha596FIMJ1H7RgfTCUEykPSMM
ZDQRctbNHrZXJDzBlApt53zJPBAqP4EXk7d7yS8dMOsiMmvnK4TjlP3+Ygy61iyOQ0vnM23lVj2O
nxmBFBRIqBj/C/mm1T26gYGdwr/WTDMDV7SuZ+g9Dx6etN8NKIJ2Vjap3oSB9hqQdgXw+rhYygWY
rhpKYT9WqJHBn/rPLUyQz+ZdKNOkVd4G01vnglFbnr7JIViAsadgQH2iVNc6FzvYxltq6CfHxNMN
wHhRnQJO+ocZFuSoEFu+bBcxr57hOb1PjfAcU5fQod4faaEW1QWcLDChHnvVkrMoEm3/Fc4Zt6pR
MLCG9FI87yjNm4hx1iZsBwocy9MeVG7Iq8TiVDhWi0Z45NOWRCZW3/nkKVwWE7+vRCBgHWyQ4jvC
uv0/EmmD8zTTgOpWz+7rGJxk3uF96GOEx02KduHYScQlOPZlka7aiFPr3MperjjwVLJYSCATi5lv
DIDGM+HccKSiNwnJJgARKzstR6381Dq+MIyatdEGxGrKa/+OrfrK4wr1sKiHfFTw7XTubriali4F
Jexv03u0Y35m7NbzGYbiBsxdb+l7VhxXW3EZOcTSGrnUW/2jvZcRVdJdCZE8Y9iaoSmkYt/5IJ2a
I7+/qXPb8o3PvgshO7eiQL1opkQOLUMynj+qq6OCPJoS2pqN6o43Hb53378qhXmyJbgk73ZbamRd
sfhtsgld3Kk9aw3QjcWbVrRQsaMzQxKmdjuLKEVgx0w5jFJO/hmkYTJ33WgkRw03gGLt+GxmYtwL
JZCBLQ9OvdwzRvBeuT2u+X3IbS9wTMNnx8AO3KFFp6obr5VptdgKTi6dzmdcdOjKliPrDO7yuAl6
sJen44QyA7OQgd1U3YqFdbguYe46ienYDt1KljY0bBjeIthPwveOZMvjsvOMUaHIXdgySH+KOFYb
ybmVChdwCZbbukbSEIHWHzU2l0djIPOwHWG0qbdYz4VCPN3xBj/9WjeJw+jHlo4p7vDxIApv2tMt
BTJqvD9iv27mfmI4HfU0AtnigOFYNW7XA6bF3YIx+Qo1KEX8W/SleQGos+YQw4wXnmIPVoTzY2jw
b9mX/l6m6FEWtxISfmdWE2i2eGAWn3t8bcjF6EEmsxMao3A3qptzu+815OB5SzIgg7Ga6gz+FWaa
e8LAVxC7MvmRC0Bi/mNxSc2zwohO97xLPbmLMiWePNwkC8fAsQs2Jq5MWEQFj37P+lzB71+GBxgP
UXeYIh5fCUkTGURc3pZzEifZs6f3ExbvRFfNtvtgw8S/UuEDGyqZzk6KvvqU1tckd7nHeMgXmfBH
a8xGxiT+EhXsSgTK3x1xVIwdAbBAPeH1hm82r7FhRd9A8JWkPwFimHR56WJpGSuNLrPJFVrkfV1k
y32gNxHmoU+Sbvz2voMRdNRYtWdGjFaO74blAhbf0F0cTEQBVRuJxrJ610dHTgK8bluaqkQkYIYX
2abgB09IHqTam6VryKwqXcycE+OyBm2LiNXe3NiyWkw7yMghfzNB0WOcjJbfBgFIownxl+0kyhmB
9Fe++1Yhnh6w1jAn6FrrhuyfcRXk4ARv1EC340fYRrKfr2YBdpkPXZY0lBXqPx2ZgNZOvT4z5rUP
+hFNlu5WOv6HfQbVDXbBkeYZa7BJb9OhfDQmWpaZAJtCQSe2cK9PI4PqXE11mMw293VqxdIqU0u3
ZLQVR1KhZTyJPNTdK6fgMoIdLxoqHoSw9Te1aGgcr9lK7fOJy/L25a9xdaxc50JIYFI1mMHKTd1Y
QT/wPThQznZysVQ0eMHs3fqQkyYXKAMWsjKPV3r9ioAqVAiYSBX8LIgRZIqNv+WmzjJGm8RA6dcn
/K9ORUgHjTEJikAL6+AKKU/C/uW+54PQIFVqJFj7JrndMttk2hnGMWVYTagyGFsqguk22Dj4nMrP
5veO5rdb3C2+66DtJliQ2gOjl/pWevVL6tPtBlEbNe0Je2EbQnrk+B4bBZ3Crg2jVC77XdW9zBtG
InsyfiCAPPZGr1mJJ9FOiJH5Q0tYw9sknuEK7ExABamvQbPX4M8MrIrtzjK8lm6eNjHMOdj/gOJC
etfuZY61Fugx9jyTq7wlvYibMFxzpTHhnsQFhTnYMZRU77AFwRibD/3o+N5hInkNOmQN8MOIXTIp
0u1AT8+f6I4E/sotjLzBgoJOOnClEn3ma4PrsjusbpBM1WmFxpJmkACNhj4obkp4KCw/qFa3swF5
8tNmjColwpsMhNWvDQpsLQuI8f3q0YApUPBgvI+dB1GJ4eMQLJPDUglZpYl4o6CgliMCNHlswfsr
bqV+qxq9splCZrLoXFHEL7yROQi5AFBwa906qL+2JuC1r9cpdV017SxJuzadye6SarpnkPFsWSVY
zQvNmoPa0RKgnhEJbfonCifmBq7M5b/6XlSNKtmeeQqgIYIXNHEiURXrhxX54Alqdy2lA7Ss5ME/
eHx6bfIRu6NL3UaZj7NxblwFWSQoTwRyuiiRRcgmx2kDRm72wDqA7kXjU9Qq0Oumh3iz6kpwzKYo
ha1JtfIwl4oJTCon+O0D6rM84uhh03x21UNObzywllWfL0rBj3h3ZY7Bqpbiw9g2xzv4OLI9AIU/
AWksVPqTaruPYL19xKaq36FpnA1xqNGKC58aHJ0NjjgMzvOXToOeVt1FJkP/wsjjl15zFyn7sC3Q
hLEjbBvoYxvsmCt2fqGvM/jogpVHMXaic8zLpg0Y403Fm5B9d2apAvGHFL/KC/Bo08uMTgBh6ZP9
ea05oHzbKKT5eSvF5fFZHEj/e5GDERpjhsWU5SxfSfwXzF4t6fQlzJHtpYnGj6+Ky/z8DDB0Ukou
wuvVhxZTyLEd+6unEo118gdi6afH2R3n3Dn8vCXGoTdndnXOinnJFLz52BmMqUzorp7vnv+LkEYn
NmxbdaEvQQODPPvsdtGkIbelV8dykDt89SeUZY0UO5ml1OGsOAzJpVSfjUCRWrx9KGn5lwSlCxiy
TvcMiIeHZ+tiDC0OgL2VdsxmeK5rBI7TN+c6isngPdhIe1RWEr7f5BikSqEu7+IxVWdS8CxEpa4V
zwD+QQShyKpCCwp/j36KaVsuCr8dUEYLOtYWd/+URnKqgbelrXHrOXq74Z7JYHo0XqTrkKj6zVvX
DnKeYRDqCkG5x4BlqAvX/EZ47gMUBg7GbtmzL8VW2yF6/fe0KrQnBeEVk3SiO99peyTELnkv/B+3
cZPsXcj3XoAFVghK2Kk+aHnE0crcKucGmBnSARuh8xP/MOWA0Q9SBKUBVW456jBfErzXcmSiQI9R
Ymfnvjils/S3JT3fi9Zk4Evi7gHzw7G03lc6Z0JfByG5jl2slf8JZ19HYRLsNLIl/jm6q8UrTIqO
YvslAw3QNWYZeuUFRMF9ZHEgazGw5Rkmkp16aJejC52ykFvkJOk0ooxYG66KNTQD+u0KJ4Oy3/r1
14wPW/G0kjR68T0t3plpjZNIGy32uWGvIgMqeUxnnqQXCJRnXPqusmpQy3/YNhKYghBw8nH5dD9n
YVqKC989Ls8MXPTEyg4kLcUX8P4gLRdSHnS8nIXzmmPYOMpwdlVQtkzdDseiPBD3HDgkF5impK4z
HYDoB9BcnbPMCJ/Js0qHeSYo+2NecaRYhLvo+UyJfa13+0tWIukI35vsoimKDkFLhRMPKN9FkIit
aR1TpJ+9pHy2VRWbK3YK0iA8o+FiMVLxxJR1WASWp+G9e+xakCXsw9tH33tCOwdtbt/t6kyJrHME
Rfb5H8xRiZGlrkCCo4bdeflXYwwH2808pi33ZvZlxAzWrS3MDvbAxfVocWknLxrO1RdHd3EQQGIh
cyamlURyq7gNOrvAAgYWG0jCpwVHm8knfUc5E82eYzycuEJwsYVQljJ+mdypDqUHtUDTfFaIuqMV
OCclBKujWAtmeDeE/dYho44q8+kzmzUpEzJWRc9O/roBJWXPUcpHYXUz3K8VSz4ZYoitUbEN1iI1
osT5OTNOAsqEvPxJw+uwtLNWUmp6msdwlgPlL57V9sP5DW94gILn9d6fgQz2uHjqYaMFrT2CGKs2
qgZCcQmiMuvOLC8/k0jBFXZ5HS4HazXtFe0sERUsKOjE4w07R42fNcsteNmAwLhXYc+o6U/fMG9G
dmFL0X11s5NwwcKFhIUKm9Tz6SuNRhacbEJGSlgJUfEbRBJsre/Apjca9G2LoekSpMAydCao3QwM
grTVWUBHD+cWV6XHA8+HJYuXROD0KEzS7CA1fgKQbz7ltCKNsmrdl417biqnsgma6Xvock3Tw32m
Njv1fx8NykJMs4CfXAQdG0B/WwW7WGAEkOfY+X8ib8KDBtiOyWI9PjZZyF2KNNaXmn6pB5OdYf/Y
Oua2XIsnBzHBW500cqf9WOnSy3PBZrR1kTsvwxcRB25sUYgjXFRJoHJBNB17TNFBuHEy0jGCP1T1
u5dVEUFbSDPx4FGa6esG97O4Qpadu0YmZL8Rsbo5HQemZl2aeS103V336cj+XRMC/tbzYTiREj2/
2lQEdEM7tAxqCVTrvbQKeWZSSSykquCNq4tR62l+xBxN3DYrn6iNmdRaJgg0NAR1Vt51RiUZr7lH
fGL65f11ZW/8G0LwmolbjtwvdJbWKB84vQtzFs/wrmqas5RNAVpk3PVoOkDeNywpwOyWH7GsqU0J
s2p+CFbQ9F+fdTJRePKv3q68RYp0/GvWOWhJVlTuJHCHcM7Mi9qZDOADE7k7wxDDvJ9VP+wBLvEu
SHHiZmqMaCl/0C4fVTcbxx1DniRJxFmkgvBmprW/veXsYeo8tekAK/n8OwnVPu14ix9eOXJ+7E0V
fPMIjJARR9T76nNIaBjLwVnHdwT2Je257ng2EcDr6mfvmsg/svVPkNB/ko+NPB5wbuc546j69YKx
+gZakjwPqyjYDFnGA1XrvNgpEMT+7fO1vh+ln0bd2A8Sror1N0bdqHRzBGXwbhA3ELS5qNqq0U8N
bAa2Eb108ZHI3Lws2lQLiPmyjhUl66PxWlnGqSjinFQBw7DYc58SJLvU+M4EMeu7lUJRKCDUDmh4
gMfG6RHyLrSJvAm5AH0TMCrjjdjpJC3/dEFo0SiAYpxRZRJ38t04MElYp4eaDu1T5SpdJEmekA/r
gTtOBbIS6qPloshyniCbHXtH/6CsGejHbdRywAhIn222XEnNDRlfwXTiv09A9bClTRRDrkfdtZlp
hoj2JQpDNdgvxlCuOzOVm2KgXFDh7fpLrXSXVPez8z5KWqf6F4yrpIzsGkhlpRaiMa3tYN7ScatW
Huu407EQuX45z2QhPsJBWnkafCm9+eemAgPwSsTfOjPwGNhVvibDm/okZoOyIHs0iMKzeROg3Zco
YxZuv2fCYrgN+/eDzG5p7cgVnfKItcr66Ly7/KaLI/oq+5TkIoQw6jXOL3c8Kmrqcu6SjwSOKSdf
IxyvMVuqNUU41y27NmLSzRATr3jmCicsVaavysY6iEJnViUTFeNOpehkr1qCFoqTC/rE+gYkPDHG
aXVpGeQOgmi19BK/N0VE0Y3Vx4B5TeepZ61l4PTG6XuDsJZF+X9e0zZVw0xxJeX8AnAGHkFD95gE
vFdAg0eK8DuPlAXsjNZdkSYQh+PQBaYANmgxF5AxDTI8SkhuSqJBxYNpbRo5Dkm+OnRhcL67EjdO
9Fr617rfxDHY/JqfQ2LeD4HgdDDskXtDjHU2i+iZYicmALCl4wZVfE3l4cZpRhssNuJVYhIzp5Sn
19VaM08vU4wvNB6P9AO2CBHStBH4H3e0eAMOvVuEBNmqnMPe5fziE2UFGDyWK++5CHikEBXcDYBl
uh/6elDtIAdE+5TFOKpdIG8BTKvnH6n4lfLbkGnSM6G1zqap7NXXsXcLzTq3Q+KgT7ptOwq1hH/4
rqF2qT7hOxF3MKxyJAQdTjXeoUc9UgG66VPLRCFBv5qvowF7H/uhEOH68p1tWxDZAeYBmeDxpic0
aOe661cP/XzAxjoXc/lVNGjsshLj+e1WYvicNNV//TuiXDPzyn60YvJyKncyJ7z5w/XK0knocqYI
ptsjihQdOJB1K67d0aXL4TAWZPAAqqSVdw+5g8uQhlzcE0u1Lg5KbULHlaOgnJnxwDshOIyI6Niw
jGd9wSVFK+0VyCXyrd/sZcYLaGTgNrB+3wioQtx4aKkvihL5Z2MR6GqazSlzrlPdZDuYT7ZpYekz
gI1BbtHSbEj+mHQ/KWM89Z0OGPNVUoHNnfXyZw7CrYiMB1tpIXI+Y5Qdm4sqyOdbsRmcKgENixTF
4DOAdsXMzeyZ6Lsra566tKy83FL5xZ9+SPld797mGMnRKSMm8X/WmuOSqAikkhkStAWCN1fe2HSO
nsj5guIoZPIT9McahEbYEP4DKsDYBCKnvqgGxGioZrefR1BgwqmrcEr60VNA5P1dnGTkg1jmWebs
W+vAAwg95/nCQGfT30qy7Gs5i4VfepxtZzzEbmkR/x21FjsPd3yDiqlYwHBYaciBsJcKbn7EO8c1
fQrATU8s201k+kFPgh/QbShxq15MRNZJ+kZQl9bANmB5+cItdpz149zgSBd/t/Y1AdEQO4XFYcWa
AMixy56PBB6ztur4r/Om0lLktCXpQbEhRnOaOIccuDNzeTeGLRGcnSmcR7Jh+BCs91cYV5d1XdxM
H7BsOMSkA2zG1fnhpkpr189gTt+oE3QK5h3IEZT5O++yYzX0oejE2rWns8NjWgyjanUktSb5couk
INRTucTBjN1R3YiiJH/Nm9eAI0kBSktkrXIe5xXmAsqR6PW2aanuYflip9ftqao8V1ucv8QV01Qr
lIzHTpsxvNR2qEjYGxPQnePfNR+OOfi6U02CJDxTBMAsTSb16DWITTmZhlkLtm1hmS1VL8OtWX8y
iDCY8HiQcSD/e6o+otuqPdo/eskvYOkYVGhR0HvGR4wdULutRHHJ4Ekru2dZEndEF8rmhro8M1in
j5bb3gIiwp7qK78ldzDzS1YIT/jCUlkC/iyPXovYAas2HRdc6Hn5Uw+yKDixpinfBe1ApgIZHDqq
muM3R7vVK6CxGac3kAORptio7LqmfASiK241AQuZ/SHjg9FqiyBQhM3/EIurbhjybLXmfQWZTMPh
dLm15ajRholtMmn6ToiS3GIvAjlewHvWKlDJKK/D18P46xwPm5ewyAl0NbT8kjR7M5zbo9ADarIU
n6j92b5PNRrnstYg5rJ8qIxwSKB7cST9HUJ7Ki+81Mw1f9knfJs6p1Lf9JaRv5MaE+y4XDlFbljW
QSL1IF52zT8nZSxeJcgfoa6gFn0F3kBEkUmt3NrUFR6xbZIMjwhKEmFtHZ2Ss7tXjbphEjBXPppT
3z/aevqKAQfonNLP6j6fW+IMkStGuwmningAJm1sGtOh1GNYwi0++BdMjj0XTuJpqxgOyzQ7ixTw
XmyJkM0UNSQ19bh7VB+FxNRWFkdmf2YddQVsi/Cjzfk5ZlBwIy7FDCdxUGjJxpFKqls7Xw/niIBA
OBGqKFntUW+5ozFqsrpzVXePmP8NH9TcP2D+q5t2acEIJbaorN9IiFxU/buYPi5vnKLG4hDiXIQ0
HQlU+Y8jyMVZlga5R0L0Zj4Q82vqfvkG/N6yF782NfnBaG8a0Zb/qE0J310nZRCUTouOH3Eeo1NE
9ewS26EOkNg6dCKnhkLf43QQ7uswf6mUqItAYTcGwPPSJWv3asmWKZU5a/AOecuJKuoEqFhZgDpy
fNrDIsKhJgNPmEILzBnSm7//Njaug7QZsc7ixINHf7H1hW+Ms9iEyXenssIEA35fvfmgGgMj709F
BKSJ4SEnttiR4KpeX5lZIcY1WhvSAgq4eerbn30frSyfq2nTcr/Nx2MUY2/P0iM/nIg2V8alYAlV
f91lLwFcS74/fxs2XGy5C/bWUUXW+/gHuSixBBuUyzBPXGEAOz6mtPrEDzae3tJUadLHpbIGPi4C
vezWltNmHMTUeB1ucyefH5pWn+mBQnLJ1sPbkWxtYI4hUCgCBAEVzxHSdHGIQLRqru7Xc0+AkHTl
//4LDi4EAV7rSRyzuTY8Xrqhw9b+VwwHFE4TtSmKymT5O77R9aLV94ljTBnoVX93sfFhkVVHZG7k
l/PPXh+/JYnUEUMl53hKMtvDaywiIQ6NP9pIo/syw4IyQhvyF0xpaWbIrKm+7SDflbJ5oWdj/ZeZ
X6YuibEnO+9ZZf6wxi9EypcOeaH0f12xAeDv495NWv0C2GSVxeEb/epC8FeU7DqAqC/3g2NeZ80k
JCVJlfnMU+Fm5XICSz9rnLPM7Mr1f0HXTQSeYBffBztUz5D8EhY8y7xpcm+SSdOcQRUBhfETXAuu
mlZJfeVMTPII/AwbwrtuyLNp8sl4E2Om7WiRS4WYPYXFWikm70cioNe64JSnix1H9SPoFU3xrIb5
VdbAMIQvpZVIV7Bg+xivW/wFfv713JCqcQfCbdRZkUI3pK9LMejcp5KpVxWSG8/kxXgXZFwDygTL
kv2iocSSEckKc0bSWb+B9D6+rchL7ahzZ4sPDslVsHllYe4eZquKFN/Edf0M4NcVvqN5JuQuuiSh
BlVOkW5cHvEB6OYrWQlp6zZ/irOiZnzkI0oJaLFXMFP+Iloz3gQbMoeTs99WAkw/kd2+1i61B0O5
saDb51b8mKX+J9tdFvsfJ8vVOAbUwQE5g/uywzSsQ4/oPRCSoUiYLNP4a26hI7kQ+pbwfSa0+XCI
KfhR5C8o34F5vTBrttwbu/PbkrOaGWofQE0WNVB1eLNgsIKVzVEhfuXMo9DrQ6QMZC7lJi5FnVa7
b6HMiNxfROMfoF0i9iQEpqx+b2UzAd7fR/OiiEjH78cg43erlZ522p/vM61//S/eAUKIEZ/dGmVe
NxsbgsGBTBUpkWUUrlJa3W/lM7eK3dbR0PTSmLnQmj/vhOK9RUQdd3fdrqqkjTS+wY0AhRIUWxCB
mRnGzieUBHJQeeJ1EHUiL6rZB63t4NseXiFdToZMwruotJXvzBPP+7+tyxyUGRNTfW6dC+38K2le
X3bho9SmICViso8qanhsz2BnE6WfO7O6oxZ9Jpvuh+wTdzYnYWG/UUWWbulEE0WKVt+VICfFDMI8
e67+UAV9r8ZLyyG/Ibs1vGB/NiOAhL/swXZig511M77oGAOVNwLzwP6mUx4HsIm/ug66rLqQukWe
8zUBS9u6BgZHcOKvTQ3BBYYjQ/MKf4es1jhqtbf48+D2SbLPMQyRs7H5PT7+4gPqTOx64mEMIwUE
YrVwxr3AOg8jhU8ZAwrgpArxLu5+OrBiqjPcMRdGvbImsPKFYfXoFZ6uKczVQrD3nkFCO7TlKynn
8mT+zjCrYMcI+qRV2SOzjxGGr/7OmyL37zsacPl6h5OrNaHlgBYRhpNnU1ls7nCUYt4Lj74OV3WB
r6wcOXQG0qjiuA5epLdUcy/DtbNRnvJjAqU8ZkNi67MQV++4G8nLzSK/l2Zm7Izeq9JbDEiqvff9
Ehjio+zvPs8FThMBOTxiL6D3d/0NGUCrHkzYISeB9wD/SKXfEDhVHp04l3Pg+gF7L6FUItNH5Jj9
yKVwP2PTfK7tDLXrz/EsoPeex+4Ledx0gCCtFbe3zkIeRpLBaUDs7KHbrhqXdKXjXBgMlP75+biO
nJ2kKIXgUXgyXZaCEOpXMGOHt5v3TubeJwhRB9BoF21iz4PuQ7OCd2gYlaZwkYc8o8dD9f+OJ6xo
Ubx3Yryr639/x5GqJFZCFOJ8LWxGWrVkGxuVAI2Dv6AFFMzZaL3l9b9rS+mBe6gxk7nqb4zbIoHs
S4HlxffW8o2Ces1reWLhc8OX+Y4MhQpGuDqvHjmDdiGUuNTAjrUn2gYXTFB28sP7ANpJTLcuhmU0
mphXfBDpRa3L5q1RboYJCq1/dq+K+cbsko/8xfv6c473c2kSmi+NVAnxJ+YLSDpaCRfAPK9q/0qG
leW8iwPIInq+iTUCrKPY+Uru9uh9RRWxeJVydxzxW/ufI+u3fDxNiK81/xLP8/x17dzTnTy9btlB
aWx8PuAKxQHGDgIeXcdU2oDZfipcz4jQRWPhQ6fGWE/ATrw+g0y/+T3caj2EV215EDkKbhYrmn9L
ViR1pj7PADIGYtOYbT0A8pV11ss6Pw8q6OTLoBZo2jsWF9N2V8uZRCoyApwuh+bBTIdOmV/WrRht
7FCo0VI8n8a1zNIxz2+wr5gbY9jZlOtn7W6izYqYQ5+hbXohmJPWFaAuDFVbWkkhDOZm+FxgpX2Z
7t9TdvCx8ss6Ua+mcCMP9WXg04/UcsppJRSFtsJup7dQeEP47G65SOecx7cmMTQBOThsOwrj0lZB
3JYo4WP8y+8XNLdDNPxleIQyN+jO8BjskDKLmH2CjFPZ0BPDHlCM4tyW5P1I2NGsKvB7EvsDK+Rh
+QiZFLjIFf5cvzi4aqXN41xdHrqmRf6TpXvVA4Adkc8BgDJ/OACnz9fQPbSO9uGebnjK3D2i5gWO
MlnABc8XNjof9nbLhM98LYVdJviEzT7djhm8fAPgqG7EjB3SvaYEPBevFrm9MZKLfRoTWcq7EPOT
wYLEuagJHaEyWjV+OxxUyzdpol039V6aYmg0V0qnBovLg3pINQA/DGVqDFeW7dGkPuUzmOgm3BNN
/I/wYAsEITh8OBGPRJ8cRKFaKTV+5SY1+UGNzCgtGryQWiKxa2TiTTbcmSwjk30bkeh2jNCv+mjj
d77dJj2AgEh6MYuddbZ6VkVY4DwOinSM/1oYD5KR5PVAGW5cy3LYym3vkAGmLZmi3iXTmV1mHxJp
7PaIWbJnR5jnQSV7Z3FtBRXB0V7rDhdKRvqd+YS70tBIK1ZyP8IT843G9SsXkxO52YPtTyWAKei5
RHGwuL8quR/ud28foBSyQCmuNyH+xyWY/ka7WT5FCLQdQmSOm9/GMiTN0jZBIT98QR9tp9UAZeDo
H1elOEU6o9tIb3wLlHQyrMR3uWx+oEL0RsSw81p5ctChltf3nFAF594h2rdZ/G15ratHc/z6KLXK
GAXNSkYDe4t0c2H3cLbS8S/IovkGQptZWBlggLg4mNrU0DcceB8hOoU0NxN7LeH9EKdOvHoM6cZd
/hYx6k+b+ivNNzXrnvNYnYz3POfu6+XDh7fKeugGo1EzFlbE/PGy5OShNhSg6fagLlvnoUOIPkj9
RCqUq67EaYSDWPopJb9NDAsUBinU6fZfg+v7eIAhT7VHi7JED+eYD1APshFS/ub1We5ZjxRfRG48
giFqpULWCHMmfL8r0nThG70hUNmpIQUhx6AEvAXKpr7JcTJ/m4XoeNi92Pf/ziFKa/aIR/NA6sfn
HCezX+69c5PLJ4dXUeyp8hwK0Vj0mwtU/Af1HfgNbwtYhhwhdoCPqvBrrtkgXICBVUoCGFiFTLPj
RY1L3gK/fkHcaXFaptUvIu1lG83UUgSLupeqxnxABtJlQIegZhKFg/hO65LCVHnV78b+XCTVIlcX
xGjpuG+MhBKPSzweQeEDbHdoeXp2Mv8zdsYmQq9KgGw/3JS1Dl8zIXwF9XWy9U1p8cbF6cbXsAz7
VBxtrq8KEi5KrjMr7LIYNYTaZEjua8GMNMG2gLYyOPQODyV3LIyWrHw+DnaIbWnap6Odh9ZE6wMR
wZwphvw0XaMUL7CksnFnvHlf5630Tk+I+y1biuy7wTMV+NryAJewqfZ8eAwFdNvVRIYpap3NfkuN
wiRwZtXFEJkXiJy+RsSWlXItFp8NYGSCQVzOAI6r/ftFT4mHsqJchovZHFKs3135gTF+u/RYiv4F
1oEhD1G/AYIUExdOMrdzxRfDDqrltMQh7voc8q1c2fRMzHNOFnz83tftYmJUHAvwkzKRcHLJC31i
WRjDFWFO3CjuwapUX0zJ40/cdZ+GDd7CEYIqXiq6SBTKO8kwNz8zFwgoV9VgTJaRaQp6N80Dqiug
DD22Cen/GFw7DSCKOPbrJSDPCWB4Tmdj2Qy+MzYVQxbpXfZAWUEcNcJPQUIuBKDDmjepZe9PVN3B
6GMYPDDbBRHAJxuD12PSDvs1qz5cZcHjMk0TyHlocSeGjAHEQ8qinYFdtQIfKk2yWLipJIWq2dRI
ceJOk9sCw6IGq9GhHb/h5bQZCufMAl5CT7QMyUY5Q85ZZbQPX0NDWsbz/Jo1NFy8aMmIFNWMKArB
5kKhJccoCkJBQXkygRXrtJeU320lfOfVpO3hV6nF8PBV3Y6sicDxitl5NeCvwDc1sjnskdbry7yI
E5nlK+eNkCvDPmL1lQSzQS11NQ5XZtKSIdw5UIHD6q/pGADSit50SuSHXTCwv6j/APfVAajNOi1C
eJwKfXdWTuuiuJNTYPqXGu7p0uHg47Ylv1L/sUv3hNtstb0WRfU7ySGGPzw4l4JP792UZ8dqgKAT
oLeEQAGaL/lK1LBwiooZ3+BpQqV50aiTtnhOLJUsb/74fkuIIIdsFpqcut5FiNdbLcUsu3cl0kZF
2UGw05s/m2lj9rMujm3csMQ1g/b3JADKPhbH49Na1PqRgM+jCxysZyJv8rJGuJECOClwTG+ZHLtk
raiDWz98BRF5B5srYhYQxSq/DChq4xQCO8oRyHdkmaQ87k+Ax/4CSmOM30FKb5A/nPCZ/yc2Epp/
a9LkJe+HHM0ngGLw/1hWD7zrsiG90gTmI+TXXIUG4d9z5w1KVYapdcaxGgzQLnDOsLheJORX1+bm
3UL/tJZv3FLKadz8ZEZi6svCUDuGeL200vEWZ2ffytK+ascKFeEFfTtMVq0laZgChpSjYDTRgkq4
YWMoy872SN3Xs1zuF2rZPMIhsnnrF+QdnTDtfiEVFqd/P98MyoIGE/q0GMal3sNCiJsTL6aswPh8
YIt32Vi+9fKQtx2nefs9qRkA20iBKPo8eJei2OcJ2ELWwe7LNe2n9VW68uPjMcDOyjCRW5Vxl0nZ
YH8glQAtni2N984ZVjieBDhT2tQbKag6UkyFzHSDTzJBN0e05gnGxcbc/Sp64oZKXTZJMpqtblIl
5jje26en3CWdKDvK7ZG6wiroXL6OegdZtAHaxmVJIwA6AS58M8DuOAjCKwmdpusTYMkS/Jjra38U
aVysZERFYjOh2vcM2nzoWQcrQ5/tEZ/bQEKFndoKWXca6v0fY/F2dTDCIFCv18E+quulOEcpPreU
pvA3nm57F2M54qDHbWyFZc2kfMJUiT0l1ua5gId0cg+nXTxiZNY1KA3DzXpX2L8FXSJgHWZKTtB7
g/xdwJWLDhy6wFOG82oGlU/9gYhUalygyq4jF32kAadV3B1LLRJD2V7PlVhR9i5vWqZ+2Xw/mH99
Ax+iLBCc/t3vUvRkGusFu/7zEC37LvE+zhCtjjfVl+0e995Do51RdvKwRGZvVD2hOIbbcIPSEaKH
RFSxw00gyDPSQu3uVad6pRgsapcDYLKCBtQqRZ9nZ7dd35izr69PDXkIuqTpBG+5msOwJmDAzn4m
iYrjhaOcicgLSKv5oMkYMh/tc0+MtKYzRQQgWzsaOlksSdsRX1XRWgCbwqPuwtR9QGZrhXpBD6d7
hdKL8QCZHrPf1kNP0ZhBtdSEcaj/2/6mlm1JEWoe7HvTv2MW2irAbn0FFsqJUzEPXcwK9XM6QyJL
h8lLRxE3kc8zf5PdM9B7Zc2s5jP0s2tUCuCN/64sWW90A2rrWuoArfKN6K4Tp8Wkvc3ijhQLoeNk
Via+eQ8MRO8ZXAQNia03Hq8QhDrrQ08NiWIyWW7ui/ItFSHp6jm5nccDRGIq8Gqs1U9nCkQO7x1a
T3qI5J3XcAj9sniH4VyBkYWq6sFNThLBSDPxnz9wLAqE/8L2kX7wzMk02t1IkGKzbawqO04OwCw5
86TraDQAR0+j/irCA9tIrLXl0MlpkdgxBNncCWyXWgGPmi9AtT9Oo6e94NBjhHpcOfZnVSCiiSUZ
2WsszgSP/k7bQZWu3CBxlR5jzIa7EI6VbcS4ULIape0ohmWHbjeKTdw6OH3p43Z/TToyOeKr+2re
0DU+jMFhROaV00Et32HIsQ+Myta6JQXBRT+f0htRSPsWHE+FZ+r+5OBgL9Kgl0DEcpcieZxmZOFF
ALKwyhIsZZhcjbGQZpDsai9SQnIE5VUHVidnQKnuXDusuWSNPoed5wSBAPGX2zwmwXG7xA7NeUEx
YNuE9mvlXGG1n2zcttsqSP+4QMwkzR6QyCp0V6UIKgXzY4KddUkTzQeOImGsYDbuUhisn7iyZvpD
Znb1u0neTQB1K0sFbRfeNqLsqEvNVP49CmhFLCOss8LHgCO+/hzHSzPQvDXeJfuIJaVLy8R3ebkS
LX4c3dpjrdhxRWZtJrBqFXU4BdSYvs/vmJwbBpCMOVWHIHe6FW/fGyqshJ/6cBwMLR5+w6lIhTsD
xFfzTIfLSHcD71QUGhQJ3xLUkpdvyWNwEEoYdCPKvZwIPTesc8sVZs3p/ACOwUhJ+VOlvu7+69Ns
zWho4liwNGhVuPPABjdS9Tz3j+Y85udlEtTh/Y8i41fAT2CQsHX11GYH6SHoJ8b8WivOJgRisEdN
hfZ5WnJKP9YwvTBgdo4xke6Wn9zQ7aqQ2J8XkkChwGN3xo8ld+lHTbxXzoWse2oPzdLPxv9P3LYg
tWP24x5e+0HPGSWqqta98pGIShtMlidhHohtfudndeSK7qUBYXc3RCo/F7ojjSWGrrYU9X/x1uuv
H6cl+kESTWG8lnnb/iSbcuzfGO7Tj2PtyJ47oxKoIXeeFFRBZoVqYIsRwaGtsEaa8X7TfaZgftQu
/3PlHf4160anksNkHkhDLs5xZINtxIJPSZgs1wshUhzVwEQMLqFNS7djiHEjVu4F3/K0bmHd7Yas
xu3G/VDoijaX9vjpm4ga0IsfmoMdtf8d3oTzHuOUohuFSSm1llVD9chRegR6JvwVzENqdsZ7Ys+3
JtHzNDmn2hpPKrr++XerZu7kRn/zwQSBohm19DychF84tqPwhUFv+Pk39sCpRbpC0J+nqKMatZI0
lUKocrLrszOpa/c+mEa+but1wnEOBh5AipzcDETSF2kD5/nAvzzmNxnyZOPcFT+tiIdgSqV3YSRd
zoPKHku6oQg2SI8CsmxvPWwGGLOBVrqbMZmDk3AYm1DPxtQGlCVYfQeLsVWauEv+MyJLyyKmSrUz
LmM/5n1AcjOf9AYTunTN/q6oOPIudVrAvQcFcJwXFKGayhndiBzzRmwq3FK956+rNf+OYUWYS674
twyI1xzWAwnpNC52X95wZcvpuevopFywdWmR3tTE5+BRH6cjMYde1ANA0WLh6+tEgraqEEqEmY0V
3bDhpkCytQ5HnLl0JON7vskOCaHXS4esmwjvVs5Ka57phvE/HblHyGUMnCzeX2eRaQGe5yYXOaPv
29iqNtFSK0G20rRbnyu6Q+0xJkWMLbJ35BNJI4u5TMfHJUNRsn0UGTHeZsUVozcntch8Giwsdp5p
YxRxDjm6ccLJ4HcUQZvA2D/hgB2U2bQ3FSsyhZOoKmGtJZZgx9EgjnyYA2ElSBpXi5iIVou4jidb
jfA5T66VTsVko35M2INwYu6+A4jOckL4AOt0VuYXx+cithsPr60gyBB2Sj3EyIHaE4m26LkL/KxB
wtfnqO7aq+0ZxmWUyR1wf3vWnZVZEz/S/fKmJwr3qTwKM4eDsp2FYW0/R0GLGCg+vGxkgK4fduh8
RHbzq42FJuUZLZMSbfw8gyF2c2M4gIvGZU/3J7FvlsZYU9gU83cgbhPvnf7WaLIrJ2wXp9+pNPyX
WdKN0okmlx3g7utCSiexqhHSDEsCkUZ9MXK83cJulGdfhptUB18BfCEf8DkWW6Y2rrkc4dmLAFzh
QTVYf3Qk/Sse8Vk9b248M0uc4cpZsU85fN9TJvvy5Bjswf9Egc8Bahq2nFUCF45WesuMqjeDDHrH
oXKyJIvOB3fD/XXz/kYy3wPIpEWKKFD8mcGH43aGetBlePIuOa89tAh2IDeQrg+J3zfq/c5xXRLX
hK5P6PVWYn+naioWR6yXsQ8uarK65FhIGPmpe/SI0Z2PARpnUg2WC4Y4gHHbRkREK47f1u4RQG7i
M7KTgEZah4O0js7NYX/NpdnThIAWo4mSl9ftmQt5vm3OO90DT6rV7zRccDi0Y5k5nJPHyP/TF0Qm
7rxEdsd6xtnlWrbEt9nkYGyaCQtBDPBKaxefun9Tt1CNh9IY+gklDh2yLahBlYY8XX0jMkrRWyJM
gHZpBxfqVZ2ak9snsUGzdL8Xm/hY1V89REilPDvzKGAY6oX8s7XD4i3MULMx4ezkeDCsxkrvcCDK
Y4UiFNhoVrVC7lxzL5H3stf3s0JbMFkz+j3/eEvkOM4TfuKZdpBm99oKxIvaXofoibE21BY8u5ek
Vvc/Td8R7xe/r6EWp5fyub7rHylvB2jRX2Nho+GnhHtWVNNspSTRDR2EmgVkKmbnOpThqVsfFS9j
d4pyiJceStY9BNmqE9IUHeRWI/s98JYL7FzerGLu3owNv3P48+pNO9+/3r8SoQuCIuCYGp4i4Iap
mK+fTt73MkQbmqk2J6ef1n0kwXYhe+rbAnGNSIXAcx5r6iaF3EDAIlYzrbMxsB2MwUQPhCdPVCi0
Dcsh5UhrlL0rHOYemjRrxsq0dgRJvuvQkX8BZZr7CLuw1ccrLo1kaC7aQhYkwWrN37uFocUEKkiZ
aLES0wpuqXaBC9zvQaU8y42APFbnRkPswyf7hXe1WtFE4sQhWKzwLCdAmYdcczBT6zR+Al3VkSQh
/DyIB2HiOER5pIsmbayA8INLZEeWqs+XZfGmyViu64nefYPAojfQDh+3OnoK+bdGCHsoPjjyGEB2
UIevAV+9Anxkcm4GR+D3COpUOZVvkOZNNJB10PmGuk1/ggxappzDJ1g1YJrTwN4KdEgnVtBBXVR9
t5+6j5WMUx6laJZegXhO8B/+TDI9iiQO7XDyZvRT29h1kgkINl7qm2FQYSJ7oy5zlP0cXIzJLhfo
emQh6Jb9vamZ7OWSz/USuncUfkKwarurAnD8dOaLl1n21vfL/eSXys3QUs73KLdbfrr7Bkm5SMyW
R2oWBDGQ+n/ecfUsDHCskXF+nhW4X6j4GP85D81qgh9FRmYPmtM2L7zgC7ZLmQZahzw31f80LFnh
gEz0BS2NlVuyquca4SlgXzq6bGe299e/6FpPFlRmmfPYa0aKdd4XIjUT8u7/HC7hhwhn2MUBaM63
dfLINMCLG8nO/QT0havRE5kJldPl6HeQMZky/MuBbMtr8EsGcShAmgzbUeI/KKZ+e4OQwuVZtEu6
aKp/1yGbp9xHuBGYF81pket6YbUY+VpIXc9Ai3COzuNDrN4Cw6nGieRKg3L4x2XvnbFhQcdAm62c
xm9P3Bk0z4KwB+PR7mwKynl0D89LahfaEMCQ9ea60l9p9HsDz9DOEBFEhRHfoO0TbJEffNN9rBs7
wX5vMtYJGVh04lmEzMwYhqa/9haxvpiNA9FGuXX3DrTP6FwWvQykfs9WVzdffhF9kO41lNNH7lfV
8JT/nn4gnh6nLgC0Nab3Lgx2YPvaGfBX8+F3+hDj9DIEiiRh7k4lWXOo3XbeYBT5V2IwYf/Q9l56
uPRF/NDVNTCs0LsYJ0SjQ+pBkQ4r8FeLQg9kjgje2wJ3FnY3a/ByKa1yysgKj/2Rz8kMOqNyt2V8
GqooZ/1Uk6J4EEGS/j+Sc+cpVoK5QNMRSY03YkEkH5m0v+G8pSFzF1fOZYguFuqG30w2yu1rtk5A
risKcwaP6dBzu1fUWI9/harZKxvSjgxnmhQhKjowuh6Im/3fXglTCF6NWiHfgtDvnTxid82+OulF
ivByysepfAaz+VFEolJr6vH9i+j8Yyvipjx630HF4CiA10ZlSDrkM3T53YNkV5yvLXEXtUKumbIZ
RMDgwnHmleAdHOI8ObOguF57+qQuoT6SE0+BKoCDIzRfeTfJC8vASdG6JGIGXmund+GtkScj0lTZ
NkD2IcgvXM3nAhx/vxcedZfGJAU4rIf0jfO9/eKhaxin0YlnId8XAZzGnpyhwVNUZ3QEbz48U24j
sQIFzbhOMdMf4O8SiT5o8o1jEYH6Zs9uqxEDOx84nj5HyqBIH6/73uYIcRCzGpeB1+50ea0kgrAL
gl2q7kBq05cjUVS/6EV68XWtn89LuIzTwgDFzHCKfj2iL2TPUczHEvsEw1O2Qt+Wx0l6PBaec9fK
Ur6zwPt9jxTTqmonYjUk/if0vXcRUEUBvvpi7H4t8gNsgwK5T6JLm8FW+iKRHabo/UxgclxldPYn
F7um+9gxecMoXTcreaZRmfPsUXN86Ro4GRowR8Ra3zPE3vIY5XS+1wzcxuc4y3meQ7KGLsCUt8oV
L+TAGe8RF3NyqMwPipRSlHB+5otA7MBNzLJ/JLMeO3rbS/HUXgUk3+JbYBB7Yx7IguYFlkCHfjE5
4qsw0ePD5MzfDkjHvGe5Dxt/Bq2TTxa+/72BmSokyLu1gu+JLcPML/q/vTcvUmIKO0OXP3xMfxns
80lYJogu0Org3e6ugUtZaskj+CBulOQ5GK9255NzMz0tTyT3iHT6V4JbZE1OfIp8ghzcvzDCTbWI
0hQi2yVGpj0HIESUmImcqBlAYpnvI4xplkBkbrfKy/Sy/MlNZVt+YM3l9MinNJE860t/9psfvwz5
zWev6jVoOv1lt6HJeIEjZbj6nNVRmHiHuy+XivOXO+7EyYuvI9PUfk3Bs58T6jrhaREkuwSr2HeK
ISCTj+Bh+XvO5rb7qmOW1/PzXGtPMvL37d9t5O01nMog66ffAOB1jzZvh794tFUA/weB+DdmOvvw
jCSkzMnEEV7MbzPX4jKvyLPKIQj1ILUenl6GXfyqmQ/P7G8wElngI0+NI2GWtW0ETpvFN1uZwvu2
WAFzAOK9Si+2GthAaJs2E89BKhkt87W/Cjxzee+7Uqx2k1poLdguspisQJUen0H+52J6q7EAehVY
EO9VeIfuncKRh5tiFK1qwRYC80e5gBC5QLbebp0b+2gXgrhiHVPpJzlUU8d3KKO1VrFDVEQAByHk
14PQr0Ttr5bNFfd+XdVYf+lcLHiCOWuQQU1ND6M83l5xiwzWiStujuf7698KdMbh+QYoVfupdPUE
atF5eGn4DEdy9KRlbbCRFzAfaUwLm2iK9bti60jxYt7Oemi+dcz41iPOdHX7KtMnkWWguLmOXuba
282pe6xpMYRyqlTrt34P7zrpluHPak4xU1c9T0U70ciIA3zpFWcIBDtQ47zlZemT65cU8P6z0VKT
nLaJ3SnnLACOlAAXMahPcEn75EILlgC2x8As/QVyGkqZ61XAvzLZMd0qKBILx4A5tFGB9KCPuYv+
eVEn9NAn2phVa5yylwXXTMyWM8y7FTp7twAQQEC9j8CND+/3rm76gciYPnDdbAucYWAe9lzyyrZO
EDp7izkFI6vHgeceFU0y+uICViu5Zw+HSdFipgYi2z2UE7JPsmPnyTAAd1yw6bilJVy9DhQ5Yinf
VPpye94VF8Wl+a4A7cyKbXxMP+2rgrQHZJDtfG8k7xP5uYT5G/auJvjP1aLAtWYC85rAz7Oc9Jz8
IDf/EkzLDZL2fj0ENmGYOtb76NbIGuDsm2Qi9taOVHaDiFkbyc1AHh8i0cuf2KrBOkwQUo8ayBA8
mDWMx8AjRtE9jm0kTHLmgVIje16gP5t3t3TDR4DllxCJaN2nq9l2Kc22f68jn8DlP8oLYrOWuvMo
SkYKj5tJlpmrQCknco1e5iW4/yUZ69zJhtxhO/iDW7pcimQ88RxnQJXUdbV+vXzjyx2Qcuu5k62N
TW9zAASnopbMWpkOC0eBRLIJ1xX9Sq1pHdp3wUoEmIS41I5uJdZhDMsW9nevIWatwTL5RFOkYqRC
UGW0LLENkjA1Hm2pCm2akojH4caOO5Vu+ysYmIG/KtI2JytD/eCOdxCCDcO9awfK8QGRZMwNSNnj
I9SQY6IYNe1YsETsCPeLjZO0cEAAOxT60xSVVXS0K6ErDt9m6WbUyWEdCtExmu+Mo2jvAZZn7MVa
tUTbjNwsrMnsVEcYcAusih1xlQZjWPNf2D3yT0IpYdYpJUPuToQxss1i/TEc2fou5iKxAxWXyZWv
y3kBt8aHXHV0PZBpgUwufJc2qdWYg6SrULjYh4eIcteIm5VCwKgwp1AkVnooMRr2gjkojAlcVrjs
HmQGzYOWZP4f8e0MA13hDk03bezL0gm9jYspwVPyLiPhD3v1Wmw9KWuGfjvha29pgT8Z86KOe1J8
bYVQAfTxuccPAS5SpQwBZ4n0jDSl+J4JLww+x3NmRNm8odnwV0IHxOwSykmf4vnWy3iHoWGIjoS8
VfUAjPzaH29sG4z92xBUJYIUlvECetFh2danOuERAqAKK8ICDXiosGdwIAdjTGqp3+h8oOeWhoDC
d5VnlfhAG+MJ0VslzFuwa+sdAwjSjvs5n8WWpoqlll4kWatVl7w6ajEVmIabuW0GefjTfDW+uIYl
ZoR0n8TpasRo+G24PVZEnvWtWkQMGRCZaYqRyNaBRM1DjaLWHme0NJeVoK/syb7DAFd7YBIW8yDm
Unpl0oClxJyaMkmRuotge/0DdFjw5B2WeePdEZcIMBlF34lzvYr1cY/iNoB6P00pI/KGbi+65zwU
RtWk/Ad/qOKWaU5xXSFme3Vt59PUpCU5hh0db7IC0VLxvlxMizCaTAz4jC6M85tm1sgkj1RR7HoW
nCOnjEb3Bre93F4Tcl2Euy7fqKejX1Yxs+5v6qXUDS+1OZw3xW78l1H7CIr9K02HZ9JvN1++FM7o
y8+DTKVSTBpCh+/pDY8vvt4yuOMzO1gWZ+CJ2SSloI4UGBWK1NJ4N0M23N7UczYePOpjXT5nBu7f
2zpgQDE1VmRmS+svTvP5PlCccE5EMl1Wt1ES7DC+6VBEATP0TzMBMo7MxgcyI6NRFGYb4pxvh45x
svmbrfb5vcMWlRhZiAUCyAFjwxlOMnfZwXr+x+xuX/ahRP3I8xByTgd3TiIrITiYRuTAQ1De19au
3Jmg3Ggs5w3IVW01WXcr7P7pJvPDW/J5mE5jVEkRv6+XHVcxwyxtBMSIUVNbZSNBMl+LpLYl6q0y
cEvzNl4gqAKorf+nfZCZKHIIch7zm1JdgT5Vuzj79h1/fR/D2YLpLz3JOIfj09v5k0g23cY5CdnE
5T0JpQ0E8+LdhJMCuG9i95i9XFpIxK9CMrDaYknF5rjKNMD44xGnVtFGhqRvCsZEP84O19q55Iqn
uGvlPvXWmbY8hglTyOPaBUoZZGtn0pW09hQ6tL/ebPzi5oa9Ln+0wYU8Rik5gLj4ttONi5lVODM0
1+9tUPs2r87uQoJrRSzK4LWMISia7uht/yqxvhrWIk8NIjGv/1Q3c6reY43cKQwjFl2fd2ILhJL4
f6Hn2LgTJB29oSR5lQMLiBDDOcmTTQusRTrXhg8QKGfKFoPCiWR19kZz9H9YlQzJhNgJ/3Ap9QRF
4gF5+FHAFw8UPunn5BOgdJV4kTJxF8uyCAGQaH8LeGa9dHmwBLR5lFxC9Ez2M2BRc/fm+8rOEUjQ
o/TLyJs09KVGTOrQAb9hC82qwUQT5e5a9oK9n8AHV9SRu5knAJ6SEgDmZUKHpdUjlPeH/73IVmad
Xty8mqyDPSw2GPQKUBdGOSYhMwOnlmdigCFLEhJm/jQfuln/4t5vRhZDTQA3EnARgg5Zsz04H8LZ
2j3mb5D5hfQpNZmN3UKS1YGWaXtef6oO8jcF6aWw7Z1TFlbimN0MzxKMMJo/93r1/JJet2QQTaca
a+35sF9lOLvcnE6RCF5uzXDgr6xrWF4JU+XMc+RWWzhd86fjK6BG+K3QwdcEs4jJwBx+22aPNmPm
0rQzMBruThBgKwdG/9L4VlMIGeVpCb4tN3/XCjs8781B3gHgDlcy1B7E9GCS+Z06GVfMbnd2Z55T
fTXrAKKzzXpIFK55Dfn+Rgsy1DogoEYq4sosEFDilrUc5bbptTFFC6U+AmwgiJwpvFdZbmSgEgy0
Lgf+ATsy+w2yxGUnOTurV304yPbU/KGMWyor2JkAmvg7kXvE/nrtBzZe7L35VGQ5754EJoi+jqUN
oXaTxVDM8dr3XcwEdYDkl6IxD0vqdudGP8KdRZCdHfovaKpDq2jX4M0sdwGCRM0VIGT5gZfo4wCQ
Rhed18P2G6nyZRdN/LNXvz+wloUTg2mCmHUu8soMaRMs6JYwJ7af8wCYG8Vm0JtibNls4pS9JYS7
6qVHqKEu5w408rw47H9hXo5NucoMUXdDNoscC6BSgIRk1op/fQXHufn1KPJeeoPiyDMN7Wh6Engr
NB2N9aBuiunDpJb4TSvdOZtwVgvqFnMCopPjcdXxDRSWc7NBaYM5hHAzzQn1JYKQencAUHggMY2V
P5d5hnm+p4kwvKNUgIUgQzsQE4g8I5DaSgv7BeKhsdN0SuY2/oNIdHQPA76oCajsJfs0Jco0dq9q
jeg15HnvcLJwTpHJxEOMbZw33oS2tPOQhUtaQGw91oITTpOKS/Tb8aOwm5Fiogq5qB0cHszig7Ui
FGGLBn4snKMmPqeMrmpsKbusAHEYFWA3pYelGeMLO0XO+7o2gQcFhb9LqpVVtY6T2s/XKhz+6FvK
qAlu+b7EgJ7Ty1HefjwqsXf5DY1XGXg9UxgW/JCE9/BZlIQTYqYDTAlaXwE4YXcdPyp1zh6kXl+L
zDV6x3quaY+czzzIKOMte/OBzQIcgGW6nGwTa5RrlYTTT/4e4NXZtoYFDkjcdbXer+Zj6cb2/Ig4
JTZohPCh/0w+74B2w3QC0TeTcaw9+iNoHYJU+mYfTTudS0uBRdTi00Lt5RLSFVtyff1eqc8yTF5i
SxsqfidyUFX+mrLCQ26ooeb4zdR5cTgL6kWZqLTLjKCG/uLWmRPBmnDw3BZGdK1Xh5p0NRT0tkOY
0jHl9ukdZzgo+MMPMEAfxoRZ5RISLQZxRM+/f4OYqGHpapDcHALteyxu70GHq0QnRit7mCFp7FRq
RmdOZeiAMFENSgtVQSmidLOuK07o6QO9suaQaaMsRa7OaOIq6DdA8+qOdAoV8ay3pS/0B4mNXef5
phnWI38luXrfrS3gfh+/L4FwHv7B4OqM8pvIR8cN5R5/tkQ9l2bdTVS/RLxfVaBfolsjRvN18CZm
YHsr2gAhdAIM7T9BjpBpZE5JfHHMYyeX9S5LuH96kKriG1+c/YFAFeKcxgHI+ofsBaMCxW/eEM/Y
lz7xvDzZ44arq0Vky8z+S18GBmsX/bNo6cTImD5XtbMMZAT/20acxQlw/GZ63jRjUhg05gIE+UMv
0NWhFhj5ZWfz4+vh+FivbNlOSENK6mP7+dDHaqT9t2ODU4ur84Kh9r98a/ilroROZMQO9Zk8P8tQ
vWc8CttsgSUN1OivpjSymsUWLg/A+n6utzGwcPO/K/guCmOpnk6u0dszCP0IexYVO1nCqyX8Fc7q
V/nhAhzX3EwBZoRq2eaepGGEnfzP5HxrRSXMGLWNVvfmdPHH/kFhFo/lBjkQeZyVAdX8wfuzrEwa
XrFcChWH8yMZxf5M4ECQ3k3GVkV+47mLdVSku1qXK0rySiNHnbiwAKA4McEiwXjmXAiAZgl/6fWG
jZ0a0k7NDF/M8QA0eWJMNOizbmwoqrFghdTkWF2cfgZPw6FOPUKF8LSiVeNy1AJ2JGqqT08Z68qE
5IFBN/tZ7Rj9/fpGwyv1M9H9PBTobbVZXexZCKSCTkGImdGIPTjRKWWqgvOT9Y70hbrSYexsJV1K
93xogGfUJgjSEd5opwyLNd/UxrpEKLYLJnKmINrfg5ROAXpticFLe5gBjVR7u2o84qkCb/FFoC36
8wLDLcWt4Ov8WrquY2hk24I5P0giWGs+86C8opUxYM1uAWvFqctJnY5KoVQSNfcP2jLrz7N54sm9
rOXOZZQ0NX7OzS95wXJcGav9Ir3clHF4A3DIOZHPQsFLKTZ3iEmdklIB4aR0AdKxirxZGH2JgXo1
lzhyMoAkPj1Z0AhK/ULKz/ELo7NNe/hWFMZgrbjq7vMSHWMjHqR5haofsnPYwhzBv2gr81IZVIaQ
lZyewntf2nH2l0etw+Awf0Fm/L0ZgyZAwXydLjhyvLqrcPITDDMnc8jwbkQQwTZKtsZDDWK37Akp
MwM6doztFS3VEsGZQgX3wI17CSKmHmPwHzrOCJFiYFKsPiQUnWclIfwCjEb8otSGN1NJ0UNnwenr
yT9DpMf3nl5G1t2GP7Zkpg0TE0irBWl0bmCnaKu+jOH67VMKOsn+C4NaZo82tNqyjOg+myrUY+pI
hBqOQ6f8h0ld2vUzIBMmfQDzlrCwHRdr96N+7CTkkN6fAAsYIOTpUKTErm1Y1+qF8MZn2JsWbWg3
En//Y6vYnw8vchB7N1vve2cKIaSCKmWTTm92jiPq9N90bFBc8S3v1rUz5c2urRq1ItJqBtE59zN0
iP7n8szHYgG0Bkre8lFVXwj/+5tbYm1+AAjRs0LvyPP4g9I3dPApjS3L5cCwBpZy3zpCDrLIWaVo
8VRPW8G1oWkPZVm8jEmtBoVRnG+2SrOA7sleKmOJ/f9O/xq/kyVN52yNZVBg0YZ8AH63lykgvg3i
KJxhNvvkFHyR/E5ZG0O0mQ4WhS4W5lInpiltwUMyyPsvooFeJBYK8ncweuDYnBmb61kN7hDEgFIB
2d6o1JIAkj4e2hVWzcEErb7B6ejwVrv2ONP39+l71j4sI1d+WnYDwzStrqe4N/aITK3W0gOWojeP
yTEA4CwywnTPBZzeSOLGE75yl3Tw3rxSZvi8SCpIkLfDRufvqdCy1JHpvvy1DBW72G3HNnCibTIs
L8vjKr8ZZFyvMX+11gFm/+Y1tU/Dhp5G6cLl36JVkjnljsiZPVz0xHZtIJSNGpzbn7mEQYZJx1+/
3bkt2/t4hMgIiUgdnFzal1PfKa1WTchAYghOdvSowmMDs0/7xGtSsYoHuEdKb8BJsM6hsrnC8eCQ
FWsuFcimbjCG4EdopYXwiObXc7K430ZSut2YdmTQeweiJob4EstqigZTqU91Vu8hxRRGhJiTQOIy
Ec/EOKoIAM2uba7rrAr0maAvUFARF06E6bmLGMTg9FeAZ+qDUgwzHBD7fzA3yW0wVP+HTVwy7ftF
pyPAWJEtHwaK1uN1qC9gQ3YvDWbd46IZ8DSx56QUyHRO5xxKfc9lFuOyN2dEMxUvKdAmIVcqzSjE
QfGJgPbBLy57JBOAQnppz4ID//A1X4B9f2W0Vej/koIn0HLH6T+LnUcUm2DLVUQQYyYuCqKfn285
+Y4lXEIOoUb8lTFMzsnd/59TSpoqTgPMIPyi+IXnJRdKDLROhrN/LPmdajMNhnnja193cxPphfuh
WIe9xagx3cpYXr1TZhml0KxhSKWvYnh9E732YnS6xLlv6H5Le2xVKPsSTHvR9L3bPYzZAWqTmrJQ
lHrOCHyX992pEWEO1xMFeswtNi42w0UeDz6+9gPtbSMXQwuEkBhxKnDUZC91ohUpufxU+I8Huu8/
RVJQwaHmNKMyt0lVyJtkQqIX+HJSKk0w1W1Xc6Z5rJHjZPrVLVZyulompFw2+3ecsuRRv32yiaBJ
ySCmS/+xsZ7P+yJvhSM65/nw2bQv63JZr0eFumjQnN3MbrOVTz2rDwEGHjckt52BplS9zVsCxnyv
GnU1bzjH0SWF0nHoKvIOUayi6E1OgP1FKGm5//7iqqxjI4Jrx4WZIl65FXnWwNu5y8/2LQErAd2Z
Z+SG0iwwYcAU3ExSBggZ71amt1LhFNUJA2x+rrTswpL0Fa948ptAX8LvoOcq21WYvk9wyU/AwnDd
qDvQ8iJHL+elG5Y0juTxjwMWUbO8TH1Pox/CHP8yhF5LRDb+ESYWTckphBbTwRXiKSzrMz9Lzttg
Z81azFawUaxZgVZ2To7gP1TewBJGhbTx1wNg5sN4vxqdSo7Rheq35AdOGEzAENz3Dg2Yb6HnA+rv
RC5kFkyWfPM+jxn17oFNusaUldyqDNWhS6xuobxoaQO+w1XA+fOcdiYNANopdYzhaQUcd+ynEqhV
Ao0oqJRbzmew48DEORKvP0mxNIECy4jTHaKsvzI9J09w6uGo0YdTOyuEMSaQS2tkfsRrhcfIjaYZ
n0wTmNzGIvBedc8jqHHHX/SHbiYo4zaFwmZVRQaE1wP+NoMluKuE404aMC9ZiSSNE4jdgwk0gi8q
vAmZmupE+EWdicssR87lL7devNj8a3jZ0+WF65reXUo/SKO+uzKrAWNM9iEGua6n16xH/PPLBl/V
fuC1c81u3ovo2BPB2+Pnq9QyZQnjArW6cQI/j6eyZJ/qrVevfbiIevt7hEfnHUBcZGslKY+uQ44z
yDgpkH2W0D6FWo7SjvoEWUE4KfPhgL46palEKyCIMkE3QBP+5KKuTQrq+sV9Sad10Q5y8gBSoM08
nZxOPh51Nd8fSWFflklWFFORyM6onckGj6j16eq/QhGaUKG98TQzkC9Adtxz2SqcmbXt9ixeGkP1
30qh5bajHlUEOPnJX0TXKULmGxZ8q29bOmtlaDAKtjn/W/jlVko385Yp77STdQSMiADlP4i72nGA
kje/3f4VzDENfnBJX2w20ID6dqdpUnsnEoHRkEN9F86R1QNzrPAMpeSMedLCUDsuNroXkh9jR71O
+yboD4xhK9Vn0AGdtB/0/8I5qsEHKozmMBp9w/LywAf4tCo3nqv26F8SWYHmCatSrjnqZELiAnev
cPTN20r8g5++cpIsoXGu6FzKMi4l7+X1RUpHEyiAHYaLZpnSyyuIBPKSaKBc78zxesUmjbqQYq00
UgDYip1QJ8DQlL6LisrwRjn4ECxAKnKueH9dNoU3F7INha4bdj5mq0lLseNmvYeZOt9NLryRwecT
PhVkwKjbPmDYnxgJBXneKu+t5TSk/S2zx7f8MRzevHsuv5fDCzBXfAMjzovX2+KGYOHyFqFTHGtl
UdNzzgYf8w50VYHNik9l2XOjf36y+rlDnh35zKjSPjudWwYzD7lHTOMYS3N9YeNqFO16bWeRtqOC
+uIn87ogFrQYETmkd5rgoMuO9OgF6fzgQZNkC1lZ1NtaW1KNraz0Rv2BCVQESB/qHow3ARqwSnS5
7NdFZW4Nhq0yZTNOzxNSnD41IYhatlWBOXU5712BHHAZftEy7qKfCOZL/unprttXoZsWbydjGG/j
BbdvzMaE2GyBulRjfSdDeM4tOk15cwYz71TEvV4j6JBLoul47CUlh4j7qBe9aY8FIRz/9wrfePDl
CHUXYHlvlrKa0E3DrFWKGByMEWQvlPM9/5z/fcLyV4Tj3kdVuFUdB7yh09ioM/5zVznWdzurd8Sp
HqkfViSxertO/r80QKWJeab57Sfb9x4kIMixdmsmoarvy9QScQRymwwYSqfSV/+JU93LRPN8vS6a
p17s0etGm/Dcw+vhWTCV61EMvWDGXr88zPakUW7+uF3AFf9cu8Hp6QzVMrC+2bDbPAZPWNdmx9Pa
r5cWlTV0/HPu+47xPBn3fVNPJ0ZspSW6UC8HWj/4Xd1hocrprJiXBftb3r28G9K9E0desYH2yDNB
EnTBD6ycIXa29iKUQIc6BdA7su7FSbgCSLUTRAAXZC1l5mx9JIPD4kdyWMI3GpbyyXLhhJd1QZwU
yRpubUA6VXDCnnSie/vu7/uZFGUkhyh0YQnDHhYLESIsBzKk9v98yPjNNRwsK06rhC2aaO455vyp
WMtMDvg1Ytr26awEhVp2XvalhB/xfO9TqG4VSFmJq4mHvPSLKjo9messuHl7ddu5eDZTCGqBUs4s
zQVt0Ayb5hdVN24XZV4ubojdqKbcOzQW+XeNNKPFE5qEOqXNSwB9qdDYRv2QmjUFpsM42vNTVxzd
4QyA84SA4ht2zQVfClWr/UoPBTN6ENGIs7RivRyt166pqBujlkKq57QpAS/t+LaJS5IrQg6IZBzf
KW5mE8HqI4l7tfhYHOe0GBMgfY0pb+ODV1SXb8lNCyuDbME+nvHnh97STEUBHXW1zh3qJ0SmzYox
D1a3fuCPB9dGNDa88CFqX6z74qaPgRIo3i9SKAqq6sGzJ4NmIzcqbF8jpgrez40BM9Q1zM+OnPFb
tE6QtD7yjr2hVu+w6pmRFSX7AScztuqGGaXC2w03sBRBecBzSM8vQkTf2/wR/cJlk+TtGtjz2Tto
bFFMjOcLBgiuw8vtl7S6kqQqDqTyBc+vK6Jg394AVlkFH8rd0CPHL6Fjt//4n46w5xwxntKV/ePw
//UMVkxxIXkGedV6eY9wJpaEGC4t6mUGU8ecMZ+GeLwTKSObJmfoyjiTTHJkR6Iw61qFh5Hd0H4p
CRgzDpdcgrmlI9S5TH5Gy7HRMXzD3uHpOnoFN2hBuPEHlTh7YuRBRWYIRBx4AY/D5+I3mOGxjStY
4IWDZSaGrezk1pgSZ5gWsd0pKfCerAL34DmRmDONiMV/jjhjSIhRGCijKeUmfhNjmhsjoB4sswZN
NiXWD/wOqqoLFW2ZyV4DMelXPvuLdoYBrxzLwEYw6tP+22hCQ4BwNlpM0a+KBoQ+VJLgjmReVV/3
qjGWwPoIKbmlviU69YwTgLZjLrKqAsYsFAp0GNyIFBTPlM/EuNnBWjzDPgH4DNik+DwIEpUqGYJG
Bn9CSu45W7lOmUW7YSIqZK5I0Gy/J2NnS5VxonztFDQxG0HiRt2DyDPAlh2TSR945bwIQN5jzGYd
3GJRzypisVY7Apcnwoj/f9u/lvBzcHKlES7/zIiL3DsViGiG67LaNFp7H4hTXs5dNon/r0vmTouR
Ke9YxbetGGGyjQ8D1+GQGYjEBKjB6QsDIxYEmafROJHRy5aBM0tzk2T51IQtXJBbwdNZA1mKbpGE
I75cr/sVaDxjc/M/decCZLGQ3RWFVswRv4kM7rFrH7icn20z0tS6L+ABuemFGy0/9ZLRncBnU+c4
3IOLj0d1hnHcBMpRH2M2EU+FNmLtLUfZ4ErPqNrCEcgiVm1fnbkYsthOYmDnJXHeGuqENePgCY87
2v8q7x8uRJv8risC1jg82KoAFCy1Gjn+M71khxpvmfurLrMgJdOstjNsLP3VfmpyPMRdiF+wjlla
nslnNgMXok11sb50WzXRADbiOzQiXlIXzHuUzoFxtTm8Hb2u2swknaLbocnSbLPcCqH+2JVqBD5J
mbT0z/APotat+a4F6uV1/EPHs9bUhR0BHvxDvG2nWFRIwNZqEOoBnTnIyHH/uCMoIPH131nUoz1a
VRTz9YFvapfwuRj/iacqdbLgSnD9c7A6E+HgZ27aoUPWaDCznwV6ft7SRIDSgIjQ7uCbusUs4LQp
rE6kYuN3czj7aokMsGt24qKsG119baQyJGvH4jx4l9yH8K+SSvlcrlNaaT+PmLZni5uG5E8tH2Gq
MD50gKYTyBgRxNMatRmwtUVpUruKEHnlC14wykzwd7E2oouVgeBz1y1NHwaLDXEisNY+oY7AWD48
ovgALdrJuc0/1V3y6ayOn6+Vpo47TYiOgxKYvLIugFZvGxE3A/ENcYm8rt5h8O107/pnKpIKpVsa
+NMD5FsvP205SXoHlyXy1b6ahRWCCuHThXgqVm7nEY6ZMSZHfKqGmvZ1+sORlsjscztJ21QuNRcC
SDnqXL8adFBWl6nbrLOynPQJv/gfC5IpyAPkEbS88OudFE1YXmU8UQzZsSHlFFOsFTMWUSOLR35M
sdVH4ws0iSZOuwFp1iXlC1EqMhwns4xt4312aNMg4SXAgMSRWjriBvYYQlvL/IAKj6vcyoV47YfQ
ry56V/NcqN/+7yaU7f/35frDCXtGrEolLZLx7PspI1z2RuZ+On15L8s68MVEDT65kpURvTWxuWQN
er4eqVIpmpIRYSdtvarlK41eZ9v5d1V4adRVa7arP+ENhAULM5xkKLGSXRbAYSYRJaGsEv/QIO5n
fJUfanCtN7mgFn2DipqFshpUP9SQCvagm+q9eXngXDvTQIZKvLi3e1GKGymEwMRkmjOOQf36Wrmv
Zs8tlqmvALVdW1OjIWHBUt5ipVInUg81j4ASx/c1vokkENZv5sJf+mO6aITwwPc3UDYT4TBOUtkl
ubUjl4hfMFZFPzXzbzAEY6YuIW1V48NVDJakPYo3WasRhsGl4TINaPLpDEwaTiYX1PjKP+Qbz3tF
abtUYK6+8LLZL8NoNDK5oasQzANrAmh4MBncctX90W0qO13jvNsjMSBlkbyHInvt7Z8NIEtZwFhh
oKYculLkUv7yDMxLyK09gOVEMJ7jpp6dtOxB3ayUS8WhL38RWAC6rH9YPq8p0803DMiogqRc7MM5
v7Z2mduF8eCYz9gaVHhXbCs3XuRPj4vrnJWTkes6yDPBfCfYsnpB1ceZxif5ZcgycA1Tvynw5l6/
HXCuY7mZoXGniKFL0FRxmHNQhc1QNmiAlVyGn3402XLG5+oubKU+D26i2mbGN3V+/XBAgEVirlsP
QAcKGJfwR2NWhfSPhBqXfApPOIOYWo9ucgWpCGS0rZ9Nik5cW4TWC3hJMZskf7j8gOHw5SXcf4eX
59YhioSOHY6jEhhPLCkmDCwBoymnnKVO9Z84BP4gd9ElXiY8PjNXA+IbLmnsAf0ptaPpQq9WbkgQ
RWhhpnibY8e6ZgrCW9iTtOKzXVKyBCF+QwZotsDcE8yWMtfu6z9g/Yrm/9o0y5QWd8KSzCvhGu7S
FMdRyas8dKRY30S4rIIeT4kSqf2BNarT20wBzQPSJDJVLE9bSu7VSXTBijN06ZUXgy5BElNBXojq
4NppKSEaeEp0Zum2YFtB2xEaIyfnDXcaDGnfvRabURr2GC9BF+OqFmbeTtLqx5lcE9KQbDmkqB6N
n2339vZnI2M4rcy5ORVBzrIxfHdepH7v/Kf49EoCUA59rYa1gnNpcV0tDivqrJ90FAFFifrFGOJ9
UPV6cdhAx9QB1GvrYNCjXr9H1Nh5ebYkFRBNrP52vsrLhiXB2ULC3TccO8RMauZk4824cCOJQDiM
ssPhKnXqI/iz/C8fur6F+3XQ93Z7Urleuu0KQ6j70zOC29toChHpGVwBqK1amTKIrR83TsBn9LUJ
t9Pv7LAIervb2DZPkKW1hnofor3IY7swmrYEniIF+bv9+qeiuVIBMy5QDmaL3s/CcO7DhbjlKun+
KJ4uoEZPDxIc+VlLds3b584rYa3ZgtkNwO9P53HjE4uMDg7mKfbwb0mk++BtCQG+68Q5/rCBv7Xg
yLioJ5e1gCRIy49X+oRQPDOoHB0nasserxmjHa/9R3k5BSFY3JZIpG4s8jOrlc9HPFxcwDX6wxPZ
dgxhnpZ0810IaJzTfNEJvrCrFKatIgmCFGuTIxvlgzj6FkdqkQwcdfF6rckAUEWuhVT0Ee5yRm1T
jyM5tdzPq4YJuwipengRNaGAM1qBmOZikuBwSdF9n6osmYtocCrXO2W2m82vbyAH8Hzh0MrNFP5l
OI7rtvc0KbjVPrBmS/Wv02OqcH/7pqzR2x4zF2dcRcHQja0/Y5p+aJns0KR/Dq7ldP+LfN7ttRTI
7n/8uWILT108F72UWce4U4aRLan+XGTqFS/nkYODm+CRqjrkTVWC0CJqlXqPNdjMlWwVgL7WpeVl
XdpaXu0Tzt/8vaO+UPIKUGMQQbqBm9qJpKdWuUtEY5E/fYK3SsgwvzO+KB1vM6dPO8Qg4hXpcocN
V1egp9PpJUPb2keeP0tKwvTagM7dx79h7Bpn5WERJmnwQ0+MrXwgI0An7OpiBcDcL/kP3Qqor7Yq
rMVZhF7N7pXMA30SfEVCTnJaXOVeFdU5Z+3vJvqUeM9RjPVzpamx7jUo7bWRakBfT1jqXVPAnYUL
YjQ1yFKWWl2ZWuxiltmkas/Z8pis4qDzHIAY6Iidmw6Utqvz4VHK9/eODPV4/rgHKclHj88DHwWY
LtZGQ6n4E/RFT1YhIQH3cy++BmC+ekp+pQuoDtsT21Z5ynu6kPxZZHqrq+CoxwVN7030e6hi140D
2oiwqDL7MwEsv2syuglGZ+q+SmXBYBK9OHXV14Wcdwct5l/aZcW47lt9Bk4+ZAw34eb0T2LcVqal
9zgIzxX1/F40gtsfb2cb0vcWbuS9nQvnvH8dJiHTY8UgHaKP3QSnctFsQGLIiU6XWSYS469qYz8M
FASG4B5a/xvyWZvaI5xxXs3h7vkcjJaJtZoSOK/5BxSHzDWyQoHUipAyotgIv9/wLfbs0cru+y5u
Fxr1CaQKdvjWmjCsLht4y1i9C9YE35PskrnpBEUmGWXoLx7wYzVyN/cVuenl2s9ArR/r9cF8FGgi
gfk0oIJBQEyM9SpRRbq9nFT9eCdMHduvDYou895hwmOgaGGMxEp9qeViNTRaBy50dLvImmAnMZzf
dGmSL3BhPR3sseyuLdeOvyRaEdyBfwJiq28MIaAbjRhum+oJe1J6rCeExML+CANQqAiEZUIinpEE
8ywUPTWQImOKOnRtceaqKFHCJD/zals95//Z9v6r19thvnjt5bFFqbvsIxhVfmyL6x1q7ajHAEMz
kX4GnMICnF8uizz9dhfJUK6tQ3+fZnd60fSDkm4reGpDOXeeeG0LrXHoOCqW7UwyFZn/lirRww6N
ntM9ox9+jF9dZp5qi/QB7RETy9mb7lObeiMTmMsWRPoBqsGODCNMY/8XUa1jazQ55KeRDE/gTE1C
l9dInsniN+cEYLjgQw8A0gnUEZjyGgs8ISMG+sFPt7MNghi5I2K8Ekpfga1P9eXQikE+T4UfX+Qa
vahQq5xN75rdzsmlQMkh9QSTXjYJHroZVZ7Tk2ZZH/fZKP4j0qBLX3QCZ/T6oIm8xpFhSgn3qHi0
KOH8lpZC08P8AI9K0kOYi6rrgubkbogSoYt+Zv+CPq4dbR71EKT6sqvRwyxJ5OTNb2Cx2cY92cI4
Dt6jWwBqDR01OKiEa34HaojR8VVHEqFrT9CJw9gdDq/a/XgYV/C4yn7cESug4zjLBiTh8y0PfoCD
s3VXwauGIPvlhvZvNsFzZmwG3ShGxSrS5Fanc1gXMuSUYiNwuTkiH9X2v14nZ/P0rdGEsIsn4pMd
CDu1LoOOXS3gm9QexwDX4ZU9y7l37XD+NF8oxXogkd1aTQtKr+vwtHPJhHuHPBUjADxJW0F5Jgii
99WC62z956ITuuReVvOvIForwAPu2AdsRDqaJbDXFhrJOwgoh1PaGQsLo9KiJCSSYkF5SF7XspsA
Pe6Af6AMybVGCavpB5ZHCa/n1izHU+6wSg7DnESom+a3vTR+auhAwSG6coHzR+xEyATf72ZIOuOG
8JgUeRrU6OvcO/lveeC/iaqTOZgsl/oG7GvYhOS1CYMnc6eJj3o8HpuBv5k5P/cdciWRojCXPMbo
RFugFWBOkA53oYkvvxwxhanjE5Vl+96+R8oduEy9ik0y3mcO12PUMA1IDcG5DelxoauEKPEdb8YW
CNAoQmnhMw6c+gfvYKmFlU//2AWi/fHQSszxcPncESjOvp8EIu/7ni9moK6+mvoA0iBF65srGlT5
WF/idgG11UnypHFHBvo774NNp/mTIfSooannMM/UPWZH8NCqC1FuUOYjRlWzw9Eo9FL0/I0wUGZb
A2R/1JLikgOgoH8qzjoiFTrx6uqM5Sv6lbTXdJfIRCiSzXrz8ySRD4ELMuUm8MZNIr5mC45lRWxh
Cw17ABywxQApdih5eRPIYu5BIcr++wW4gRD4rKgbjH8LfK3PfKKVK8wxqXqRJ1XMGGyXju5TaEbU
mYl7JsPd05Tnl4nygCiCg3joeXM+25EkNHU7KU2HDCLx7pPk84BdIa/MB1vSd8LbkG8o/BLMzbPG
rrGOGbi5w3m+W8U1SzF85qzhRUwHFtzDZOhnif1Fzk4JEJMoC3utTwwkKg2vYRFJ1tHGgCZwNDke
jxmx1G7Nf/dPocoeSk3QKiBH0hdysi6czORT4vKGivwX8Dh7sDIpfsAm70QT1bnlk3ARSQuqUuD8
Tl4XVWugiOHPHd7DdEt85oC3VEr9O/lEDWI7flTf8tLLvIOWlpl685ka7O/ryuWpoPKNPT3bgYhv
+V75KiT5rEbEiGhfzrWcy7dRH6iZb+uMiOR+4nEe/9VRRgycBDjFmFwCmowjwhJP+xsWdDa5MJWy
VmGKdy+uaGLUI2WQIGBObxa4c1vadRmtKLXQuPJolQqyZsrpC3Jryel4PLNUHEojKGGN/lJQx3vL
ozV1nMpwYOwHTzOcK8AlAOiq4KGCHqrzCZE1A33xVKOOW9Z/qFHGymvKAhxfFRKwSwYz2RXqAqMK
BmVS0oI561kyokgsS9d/opuzgFjt+SqqgdphHVbpIl2+mXSG97QxPHBpH+Ot9QRr71Hvg1MwIx+s
4hddGV/V+wE6r7jE+naEtoNBRtvlADALKtXSjJdIgkmTT89B/LlCpyHbFcm1/b5bnf3QnpwDG2tw
h+AKkzsl5rtI8fXs7W3qiaVRmSPU9rScH5TQYGp1+NBVWkfK1W9kzVChF0/orsSk5DLf9k2eR1hR
+iC2cZYbraGmRFoq+d/BRRy3tEfVtAyWWUjhvgqhaRzPbV4PP65I7L0NIpsd7phaUW2Cp1jsFjOs
6pTjTZFFNUE5bSJVuww0Dyxo5CeHAyMVZGP4azBxtYHUHfUVtJmYIGjle5uxSeXxt+INVyAzEdj6
LYoaMSPcNmhGokIWwZLBr3sVGABfn7osmC0cuSSXw+7kz96Km/9jiPg0C/ZxQDhnnGh4+MnIEzl5
HeCiNha1Pp9uuOeMkpYPhBcoKshCXGe2+mM9s1HCaje7W+0FYLH+TEl5Kk4wCcW/Z02LSDRc7EKa
UvfU5kVCy/nDEC9Gc6lcXpM8A+IHCRlMHd2P9T5F2c1Wl3/8M+tOxSyVnic0+IA2o0XwG1/ogvjP
OHoSpKa15JFw3WqI+ZHt2Kks5HjQN727yytolEaI6DYvkBZH5zV5cRMnVf6B9iQhW0158Q+4vyaH
tYBRLUEGtgUdky18sVwz2+0Zs25o6U6JHHDY5XEjOStikmXSJxfFcU7YgqT+3i937vOuOXyYJjSl
RtbFynyPn61K3VKxVjm8dEnW5oZjnIULc5AodJg6rv/Qgw8NcvamKb0QQlex61YPfbKskNHmYzqz
KFkm729jHwX5jCCwy4t6femigFCBu+b/Kr3rD9gN1pV4Ai/lSS5Z/8/3TsfcWdH1Edi1JlRwn+MZ
YlSogTTQIkr87Fz5bYOLSg4KWulEFZCp4XYk7eHI3hEWz+s6E3Mh1FniSfV8QLiBCjCzvI4z4Psg
nypN9k/eTbdNQB40CIhpY0SM3CCodjgRKPnNyu0feuTqetl6BMrNTb2mKbigDK5JVp9iGid9kc5Y
yjM/9yWQYLaI/urrPpMsQd5vnwZE5qBOQqr2GJg3qW7MpDU8EwGu6Wm07i3sK/3LbSDV/w3FqF83
DbwmWkPMsG39KvUEq1vw8q9x3/jQwn+8PPb9ZvrMhgkXx+MZKJ24aJm3TAR8MDBhLu8+K2MtUwmA
8H7f574l5O02Ky3oHrwwhVAK2b0sNJE5wMzMCbllvIzCJ+frWM05/cI8Uf0N7Q6KWcRP3Zc6VnkM
f32jiIYlhQv638+1Ehgof/7+2TQG5j1u20lcKgYYU575yGBh67bY7Fda5dN9W2s1CR1xk0E7gfuK
BPia8kr7+UEVcKE+IX+A/GMW8kd+MCbP39FjEEBrffQ2hgYCgGv+AZWYSSJxP1S+gPpsfwY4fxG5
7j/JTskKJkOYRiZQdl6Lwh1oCEHW9hgL5/F6coKum/d2L/9BqbWZVoka4tvRmqYEkt9yLl2UEwHQ
rERr8tymTXE0uZhKXhPoja+z6L5X88pNJhHWClOCRWfZnLwWxB8NZITMIAYgk9onJdruVFssNNKm
k+AJNXhOJokPsqqsYpE8bEBvLRwQa4Y4GF62aTwYtd45eRHJn8+kwuomAhBjnKrnFd9fjsfhJb5a
QLfiyV9Vuyb6YDMeavK+PdYKCNm8zgAz973+oFV8nsTCS/imSEgO/XrERW1yxNMOooZAgl0RJr5W
lFDwfFE4/GfXW7dhBfIqE1XWMCH5NMEbMFW6j8yAc4veVxFwnRfXl9gGDTDJdMyX1uKESZX8zSZN
nhzrB/ukf0ZGZdoQLnV62rtmvKGjKQjyPm/mBbXDCSZ3OYinsOrK9AbG79vXxrCotc2i/npvN78S
zpxplEne7zAjqIdQ8zs3cKCP7O1x+rusiw4Un/ijmuh/+K68hBaxc6Qc2VOjeSjOWOwLeHJPmUui
ij3+97VnN8RaKV8Q/y5kcL97p9RZsmXTKdN8677Ms0sEIzuKH1MvXfYmVCZ6bNHBZRhC+UY8CXLS
MVPvIQb9QJslWcS1KLRKOXXO7EcehU1YrPxWSEv45nFBaaKZMGUMSwvqtn6aTylSO/IAp3Kp0/lB
u8a1eNszxPsNJbn4H80wfdT8e/AlDKOe2NeLMExX1ceOyy3XRVc6HLLrMPqyezDOO8meLk5Qpt+I
DQgGIiQORDf0yPshl6IIFoyZEAJvWMATTghxtgR0SRophid4zWJky6Y+2vKlVU3+e3JUNDHLBboU
/aghCSdvGa3Cmf2HPqPTfXfvJ3sE+FnmFWSl33LbYSD9UyMPWhLtbYo+fHUT1td8havmKm6vLk9T
nDsIbeKv+yuWNOQJKpR+1jvQl/2GuGDbJXWjlaH/W/1I5I5cnNfmz9osnctAyjty31ui3wrzDPTu
xPO+MyM8MNFKLv9Jzz2E1pr6CAUXDTCeM2RAfHARnV1iqLGVdgrjxPQjzacxXIrQzCVS0dpNPvIQ
YUaTU1iqF1XmVqWNJL1kXNsm+cEMYMX7MHfEcWWFo4nTfGZ9DRqciglqVv96Q3oJe7orQ75Sfjgp
K2O9eOgN4BdSQPb6eLConrAlRsiodPWEK1Br8WcJF38Rc5C4hN8ztoWaHM2hQ+XQ2rxEuB2zGImu
FP1MNJHTQ22tdLStuIgEX0nx0GvelhXtmmFnzd7fVe5l7EIa6g6eFL4fCB2np6BO8EYQsqcojHsK
knmuQA1P6jHWOxRQ9xcNVzySO8nVe1yzBSE9BeHOLKx9XN55Sjf/A3wzHc7nRSPSYqC2bGwfqpOO
5XU4zRTJ/x/VIVhc0W0KmWkjZT4GD+9V3gk84NKUE34DIAXCu7CtzHG/Weza4AudmMt1PB/RrV62
6ZZDAfktkNsfoGWaWiF32T5l9ZcZp2ytn6DCOXp6uRAaAbYUzX98LWtyueBvFdPEikSq67Y3LLyp
8X5GFSVdPpyZ9jv8BZIbiwqsIGKEfFue44PM2aQR7bn+Q6iHwIkFwFK1x80VafYUJyldYDn0uHlS
TETRxxOjUV5mCA4PIYr/SxyrCkZrtO1dITKX6gJUrZM5WDGGBlq4K9sjt3ta1CRl6nmZkB3Xf1To
ePELG83cEiU4LjXSFIpotvs3K201JzYX+dMQLjrskV4mHW4vMyEEYbhzWB7P6ASFYh18NPltJXmP
x729XSSbtmE+HXa1dgugiIAQ50cyvZ/6cAOp9PnwPk4cJ8stGNrJNX/jMWYirkktCeLEI9ay/gz1
NTEzM3hP9JKih/to5475SPzHSyEz41C7SQEB3nhvsDzVeB7N63kvD9QVMWhWcrNphNZFuMKmzNhI
pziTtc2AZq57MWeQLJY5UcAyeO4rm8npFh/yxoAwzPwhy6YGGAKopE+bk6e3sLeyAIhUgAIjdHyf
o1t1j56awwnjC3p0DOlTv9GdvfVZitQziOh6Om6Vg9DPWOZ3uN01OUF/wzfs2IwGko5AonolMJ9e
24BmsNUg72HMA2ISDqTetOKwCBLeo4dCzAQO2eKO4irLdC1GhOeY5rKnfdxccCO69X3HkMAEIGUL
3VsE0uu4cxlFbtMJE+2ptWZ9Mqp//Y2JGQGWJuKhwQ+qMIZg9gRpsNZ7fAMZzPFSoFe+3/oLLRGJ
hiNuwNodPc+Z8l3UW8O95ll/NDi6kk1Oq3b4/vemKiTJoKUehIMIhx1AeQEbUMMDf03TPm9KWzMf
XzplEyFihhd3v467Zl5wdKIeh3SRFQ0oPvbuwBsMpLtZCpPyehVnv+9QhHyTMlWwl5FQ1jEmVRpm
dTmn2h8XxhT5PR5MG7x4/HewyHmW89o2jn0nRdkaw9rXsSi2nUsGnsw0cjLy/gtTm5YtG1Pmsv/k
c263bO9kFySH7wE4g8b3uABgdrgKM288xeBX57Qil92UHb7HfYQroaMRPVxs5mXHl5Al7m2eyMgi
0ZJKJ5AQ92DTe3XD5jkt92DkbefBWSE6tVbmEmSPNJklO3ajnyvN+6uPC9WLJwISeV7xKYnidU1x
hUXT7hXEB4aOGEBdGbExP3UchQoxCjzTZgBI/YhG6UEhZsPuND9e3jEl47Xnpz5aJwlQPjkyR+3g
fPnkJlU3vpM7hoTFbHsF2jWg1pMjF2ud8qVf8KDabopsNSLNskWYk9+PG5Zz4MAotiLW3rhYXqb6
0Th96pDYHZ6M4BrMNbP+vwtMRQ/H7flYtx7lC5bv51ZUyY/rZXhuah92oYquZmE32/Q64Af4nStC
Rv6eBG+PUShE7stgDZJh9CXoZbVzcnGaMF8ofOKyG+XsQkXiOVMGn/jWGcRJgFfeQVpqS9VnsbjL
ecnRn447wbL0EAzhYNyxufMqUv+1jAxN7qriKX/NUeRJ2/IIrmQavKczMPJUz2HCS0lNf33CeV3V
f6NcTXcanii5J46SavNSUB61mQ4m9Jwlf2K4W5RFNCfJy5l0v0ejXD+nBHPYGU9CPILS1R95iV1a
RIFvH+fj8/zXWQS97V0KTEgg73bJbMyoXVj/iTXZwhVXE5e9R3i+unicnOhNlVHpEYct5EEFLkqZ
w7hXPJFzDpfpsiGQryiOwXBkaTmUC5JOc2vBtzWO4ODeaGlFV8U5ZHBIAc/qnymTy5in76qteBP6
+aC/w0jVNRX95qC+Ffzrykm8VRaFhsxuaYlGk6rvwWX6uPx9YjQNCp7A6LAcZqHitv2Ipaf5I9Og
HkvjMl6BMBI1ERD2DZvq9Daj7PJ9g7j2+lnpLZ+u0BgCQX1IkuNqm+7XCbsD0+Dt9fH57z0XDmaT
kirnvHXnZYraUF2EBkm9vQMRrpRezNZcNOjMulyD17p68ww9Gs/beXIlASi0BsHpxJs32Ywx20WU
jWJyb9MblzH7pTysaDUFH6J7OyYl21Sg97XYUhZnIIOQLN3ZGQEgSvLEDKJaj/LFK/c/zhH3PSy4
NmiCu4U0yrVu0gEDmyPRoJiIBRM2sJiMk/iA47iE38NjEzHNt9NV4BbSwyBDtnBKuss3hM3Xdonj
iyC+7GMIvK2O6C5r9qnXrT85njgi71Q7KJAc7rBLyfOztnila7ZABHC6bLvBb3lOLkoeHWbTdKC4
Bhapzi1QxNZY9Y4I9JHvs6i/xTMDpF3tYyWCv95NyWMkBuXlHicorwAlr59nYOLDXLmEOds/W9SK
+tY1bkkQbQw6G0GSt+YhOZygBfV34Ba26Omv+hRBxRp1FPB0IBlJPKq4z8EV7/wd7qCEhTSWArSj
xQpNHPanEpzaocp7IScUPIgqzYrDwdB2CkKe+x85oYLFogjtLDIMJExmwuOS+NokGKMbMKdYJrZ8
8H6tFuOPEiwubqVBJA2EUEW7Bugu4I8+I9o3A2zWUb8cRAEngFi1Jw9D84vbOh+ZbbbAk2wYAHmD
L66ONNsqiD3TarC8zPT19qUN4HdgjZfyFEa+JuoGWRktRoowzDXOiR8WgGhAm0TMiBsTMVlieaUD
wQW9gB8qbD9cy11gXZWOXC93LDtrRllBF3fYNoRGOJI02kM6nL478SWpIPR/PV9bWLo0E72jB0SG
u3K7KyO+kbMJaeKaBmZIA7u57BApWYCMo//fDvYuF3Ghqhor2jMogSYYUAETkRhrbeE9EUt4uE09
JGG6/0gk7c1GFw5q4dFIQqnNVEuDJyKBtIgIqC6gs/ecVzBLXD9BL/hk3ZJsxPdD4Laiy6XmUUiW
QiJtGRa+SJE6KgkChGfKaDcVc3ckJBtkXkZveT3IqQu5stixF6VDDulG3DYI/WFV4+jBVzEcGUDI
rMWUeoFpVS5QeDSLhadpfPO4PyLhU4o+hH/kqEBG7EAnCVYYgxUQbDQtLNMIJACu5fjSkt7/yYUz
I81WRNM7vJT5KipFrGdQ2CWg2xPEg1mzAOnxrcr0UVlJg4k3rXd7d5a9tZE+11+Jr8Ffh4Aba6vS
5UaruyccEDirphD+yc+SIzLgaHeSVuYqmgFT1jOSTA8dpJ4rRpO+5dRxqOD3my6+Q2dVSWqiMPnr
dX6taOgiz8JCGD0/vHA59yawJw7yuiCC+U+KljSXfktRvYfssOqy/1djVpABoN0bAtFgDPC0F9+m
wxyCkw3qOvwLCA0jiEjHKDgTniSjkaCMyJmsKQC6+Xu5nzK3ItYH4pqCHHzz4zWH46/u+YDgUcc2
pku2dj+0nY/CG+Im5aZlGWhMA385WpR5zAZaqOs7YgeVS5ULKPC0xIakI+m0bSyiNnyzhXGXAugs
NaPY2ZtLGtMo6gRSNaZDaXY33WNA/kbe3hE8DgzYvLZ4knV6PlsfB9KSI9xLfNzdqK+Imk1hQtcD
lRj5MU7BEclURgX0NpBLqkNTPbRjGJ0qu6dKpfwJK8VqhsQpp5oMPiuBhJOV1N7c5ANf/U9kcXkF
29MjjctwBRWQIE7ExDe1hFbHF+IzOmALk6jpqz5HhBNXwkBDtBfutF3uCO47chKMUixbuGct1C+t
mKEHqK4ZJXM+apvCaCtEHGh0g6J16ptUn+YErsw65DnooyjqOtn2ebZoLQ8NBoSvyy6PUzdyK42o
KjME4T/dM0zA+pg0MBBeVCIdpGrtzNc/JGy0wfSB9vIVoApWgekoZdZZdSa3JyLEUk4vxbFDEqRo
xLX8nUZn+C5h5xvbagiKm+C2+F5S9KZOsRbRnVgVn6J3mtzLFCHEKZH6ixV+7NYJxZQfN0VUACvC
f2NoKjEwq8VCozHlBF6hfUqAyR8QCud2KyXdjLYWL2dFWURVrHeJLJJA3QXkhmCGfEgm7piCRDmZ
fv+VnGbu7OZfh9IIalj5fTAIJ2ePcsaK8+lBQG2iFRV0FtEsTzj5H/ka1WaXO1uBP2s8oTj8ASJ1
xZ+baYuLPySJprzoBuR37ClRp1wahIDwgzKa9Be2EhtBGp/cxd6esK4CYBXXj2GmUMBoEF5dN2gT
a3mminUpug7pCfhIu9sHkpVcHzctdn9gxdXSiAplxgPAcYMKDfZ8aC+3xrveD2bsDh+B/BYCtvsP
Aszryiae+7Yug/ve/rKj5786s8pgi5wtuenKJ1SiIDpajwlyuFQQhBw7a6RE4qC8cMt7PQtrmvvX
7B0aReBGKqXIwnwPHGvMujJKZEd2iaYnDxZy3lP6Jytc2UZwwjAAqNCg2vxHrWmQzVqnY7Km/JDO
ESWyCgpdJfJz2R33wK2NWs3R4/4AqXlt7BuKFSUz9S+ZUUBH9NSV4Gj0niJI2aZGmpa4NKYIt7sj
JpfBA3eaMTWj4M2Fs90T286IKxMb1EwGPitQUxen1blGX7F2Ux7ncAYezmKvtMKGOlm9HUImZSm2
MoIFDR8XdjnKC0aTfVG8m0U/Qw2URt0bjpIGr2KQGbd2UnI32lTtIZx7YHLiv8y9T5TS/UsF7t/z
MHoI2hgffLFpNP5dOPSpcUOoUF0K4sRjzF8S0kUhcTvHq+av3bGyQp5164HtQs2G0cYXa27mNVVP
NcIC/6luolqWrL3Pgo35phEZ1UL3ptJHZaHjYHDW+Rg6z3DgnmMlQn+qAN71B/3C7VPZdRiyfj3e
7QzsrVAiEuYYH2SuiCdLdrHret8Z12qhTAC1Eg8+PgBJ8HZwWiE6rCc2koJYwsx8xi1tnzN1ZOqQ
BIznrAgSh9lMzb3zM1QcOnWdUK6FD3Rp2138uSkXhjesLh2ZVbOT/yFP9GR1TX0POgk0o7E9r+u9
GARFdAvj4hVHqii17AkggZgabQ3T6Q8YYGL4TBg0R+e0JrHfYSTc1Hm5gLCYAnebuVCGItDibIG2
BDA8rAKNk2PqF2hk1Ek36ZBm5X5UsdR7D3it20ja2iJU9jyXZn7oP9a+tryPnWjt+wFMIloTUlnq
Lvzm2aKNvsXDCm+1OTXPvDgYP5+nuaZBThDyIq7QB7Ez8egRoHgdiG3xnf/NQCgDWAHTEvkciiRF
10kAosr9c6ed7dEHEF45R1hj1Cmk0RdLgVRnf7sMT9T79OAYZJ4LBYQCnydT2IWFyhK+S0h8sIbZ
ZzPUc47F2s9g5WSJlyqZK+RBGb/VLtijt2o0+UCuLqjleV2bepQSb7ZbADT1iqh/5MRebRQ4pHPu
rdq9bgrllFzvCvPlxZJ744L90S2ujlEpIVz4tIj7G1n2mJxOFHYdze2RLAxBT/yM835jPrvAYKHV
NGY4ojdfsZ16NHdBTCUWnr+BxsYpKn+MkU5QpILYVGug8F8cuD8uKa2KuNi5HdVhnTLVLkaA8PRv
4a9Vxw5fU81RwXqCanW8HXcyT0xHdtXsC7VALOYXz3yBy1aOqVvRpElxM/krI3fc+PaoAnBx0WrA
MLV9wsqQ6wtGGG6Yh8bG99ez/aqcPH671JEfHHrCc93P3oK8KXAN+/hHHrEj9mF8NGeGMmCK2jB9
gaF+Sq/Vlq8SujvGLONqgU42Xp6Cbgvdv/6s0mJ7b+psTND7rLy5O8yvVtBlv+b3Y2voxgOvvhuj
T2uzMnkBo9soI7tMNslR/ER25BnyIhWD4UXhhW/Lo8vgpP2uttUIdI0JaAa0UitXzyhUv++1Qu0w
Ed/6uMRFk/7ZLsdjFG6bo2B9vjTKQv59V4u/2RJsDewJvkimSWwsENJ7BA+IxiHOM9hYnVAv9+KU
WhCUBgmvOQnhWtFa4L2GBj8Ujzf0GGfm1pN7Odx4dDsJheQDsSASqxvWcWe3k6TYfmEnjVHP8p8p
BDENhyj+IoWti0UdiqK25mXKHX2q8SKSnwgSHQ8MKdy+9YZ5SPROpZ38lGy9yRsiW/u6cKKUXsHI
BGF7JUCzBueqisPgIlsaF5zY2zHWP4ghVBWKG2q88ovb1WHegZvpO2hbsWqUmwsWsNkIebgqpyEP
Y7eus6qbOunre+KGq78TQnU3RgwVT5HW8mkdTbvDM+JqquKMmnCrdV0sN4xDXS5oF/Xi8zV4UUP6
HkV7Llhhkkss8DLh+/BbsGZNxs2FjqqIRzdsSMbof/0Wb9oZpvoMi1vKmYX1SbfaAzBbCoZESmvO
dauuDEgOOftrDJk49YUqtR9SFuFu8vsSIoj3JaQUuZFMa9xKtv3Tcvo3a1fubMRCWWbBYN7AAgj9
KDpZEoYWw5Q3+iZYCGpc+CdFGpqc2gWJeFzjvIqCxMGH1aIBARPnXZcZFxHWWpfMibrmfZvELsT8
ACWbP8H7ViQybZnAejpRWAaIxMmk7TZEEQB9K/MLVEfZfrsOF7bRFqpYNuhJLFrtLv1BUAjM61Yx
MQPE2ZBmax1MD6/yvGExI9qm4bl691W6jvVj70aUnd5emwXmx/lqgl/FVXL8zAiQiaH5VQYHqxqf
1k5drSG7wKvoi1tNHgWGCx3EdN7792pPebhqIT9yjxsGnVydrAa6Dn9AVg+sfKcPLnd4eSZd58S6
RpHwqdV3CMs0O2z9xr7sKkFJ3CU96WaYUooa3XbBMK0KZj7PYkltkNinKjuMvdH85uBT877SrFzs
B7elQfKdTJIvoDWSnqyHC9zTfwo+gGdRj4jRQU2qNal2VTrma36yp+zitLTZ21YMbY8KNWOowET0
Nvb04sdSaFsAVEzucvyNyFRs5ObKLL8HP5zBd/BjJtzAmo1BqlbQaDklZFk7vMZDTmNmcgpN6ORa
LyrOOwtSmzfOSqbUgLAKXsj7ebfk3UP5u4yhTazgPgw6euuloczELLiD25Emg3fqwYRvtKvnp9Hc
yF/85ZNjZJKG0XEh/oAnN4Hz9FEoPlMoag/FmqeqRGcIJNv0CeoEglTgZ7mLTqrrivZErB1qw6va
rvL+V75RIIC6UPjxQ4+mrJGlZzMudtqB6Ip8WANyrD8+ZrYmSgudGjqjCh+tN/tMMvXAM1UXtpNB
YSzj+W36Y/kDiNvaYPdBvNzV4kXRG9nV1fbFbtzcrYH1l9YtGoj2N9gHNTrjZIe/sSqSsKFYKWgO
XxfNgqP8KrrVOGs28btjSpvR5iK4pMKf6INpMsmez//qyYKPURks3AjsWFOM6aSn21EEXYtAMebx
DHdY4DT/EMk5vOg2akVBJUJhFfQ9KW8bqsbapodj83SbgfTZLD3SQuMpqUBYisZIYhznPIVYGmFs
ZKF+0oC7gVEm0yEEe9xlihVWOxmB3RdK9g8RASBVYotktWbjpFFFWIDtenEfFJPwSBDGQM+mtHUg
uMuQhwHTLtQEviv/Rqx2MzP2xpwBp6vIw7B66pc1utMxKXxi1R0K79OQwExr5wv5AwhSXyCgOLfu
S4KcHnI7dbiLeuA4YDlXe2dctdCwmVlIVheL366WIsnua9Ihbx0v4/+6o506/96oZKVSrlfQwmdh
f+tB3caDkUUrzxR+ZYNknKCfLykj/k8l6gawySohQCwjJwmfBvXSlNpsSaxNKiFzUT3AYnWcjN4K
dY9740n7WSv5TD9+UZu7NygC4yDN2020CpteZ6TUnAEZQuT88ANiE9NLa2sYDGP7omyyxhCrl/tO
3PMaln0zmSJFBfeKH5m03X5qrjZsJPWfpL4mLleQ1O3klDkr9BVKnZBWQQQC5EwfTRbc8p66OyVR
f/yc4hfKlq7GP5Pl6qSvf628tckYCetQPyR6omyxfaA+/QYk4PXPSTAFroLOwpvaJM5jlddjByIu
cW+49OnHynUL115VpOuMDQme/DfYGbqbVK2LjJBosCFrhiA8xEqD1Lbjt2VqoAbSvp5SvJm31IrD
7nkPEvq7xhm3PmGTknvgpZ/YIzjwxMN2SLGLyHrB2fc6HqvI7EXUfxgE+9Y2KI/rMMWix4hYxuWK
Uh7/IFOSVs0JnkRKB8T7hPVX3zuXAXcdM6PVX4DCw460GAdbCjbsiwLct7TphC+RhIBQSGmOrttQ
wIBqI4SW5e7zYJ6catMA/syhq69J/fsg6vrnQ2egMJRpIfH8X/yjvttpm6vnprkPXWlFpH0rl0uC
Cu0p14T26T+H+bYOf/STkBuBiqj4qDCNv5fFZCLa/HaJ7wkD/JfqFGExY7Sc579kZFjoXD8k5rwL
JjXtuTHfOUNPx4TO5EQCpKD8k937ZW/WvwcC5y+h7SdchLDADlXiTSU4OfXs3vatDOkQUC+LCLxg
lGBZsl3F67727sLXe+MQkrZHynuZld4aJP7XW6L85TfzlJ0uM4QC5e1YtZx+tOFGH3sFsuT6cCBY
Ldt0Y9zraLf17o3dXrG4wWYgm/hmk95ND6YNWc+WVT0aS77DALOA5PdvXi74AOV91cPGMBV33iu2
UKMbLs9E7n2I24CQtaV5LPjtJcmSL1gpp3BSdVEV3KpVd8q29Rtjx8mDhz6mRtOOyFPYIMbytwfg
KKPP+bTPRtzaEqqZJtSr4z/YF3IOVVVbR69HMFp1hmT3Aq24oiasBHlbgcYEFi++ImQjQZEGH4VU
jz2hI7+1L5KaMnTolpgA8LBEnfA70siWnTJajVohuo++Hv0KUeCiRmeLybm8Xge4v+TfkBvtQgXL
4BoCUWlaqFKcvUXeHMS4TWWBcyaGpsgnMJGSKm3p89112YQR/tXoo8cWUaOj87NwdCMkNR0+ly5P
xzWPudofHp2C/uCAWx+uuyzeB1FP9/Ir+juoxZiXg/7eyE7JjiCKeh8fGluquVKV8QeCqN4QXwjO
E/VMd/wqNAQBnPR1riTixjmjiCvA3tVLrIzw98VHQOICovNoIYkl9YrehhbJgGbIvgbiBYJsj/DR
WwIAmNLt20I3MnZ6zfSzIAWKX48tqAaDcWv21CBm23mA0upWEfWrZcZAczLfrV23TD8cC7CzUI3Y
54zQOwKl+Ynm+x+sAbcemNRfY6o/ZHLz3OHfp3DGpiNuS6k9XBnqFVseU0Y7KS9TEY89WI9398jT
HnQPdFcpm0YshJSFbz+iB7TSUUdv6Mw9bwMdAXTS570oEaC+NtJmVU6EpbhkYZiACvOwJ6vcwWYY
LgkdMqszOlbZAfRDtey9vI71VbSTpS/I1B3gC+ct6FD6NbVKV28SaTu2GmKOgbzvLqcJOVzxLtn2
9xTc5ZPji5RL9ZkSdnxdthpbyNd362qZrzTR3mkndM5JR7Q5Fb6exGSgb/dIln5d2ADoTn+kzRwF
NrlNq6c6saM9Yz1H9Yjeefw3heVJu8Bsdiz6ialTT1RicvbcXphhpO0UEYWzIxHYHDprCwbMmXIV
kqx+YXI3PtzwJB74kKFNeFDOx0TxatmexVObU/unGBnaEsp8vrMEvyi9E1UUH68vDcJGOmpkt5i0
dhRO/sBkq7o4Vp7wzzIGFNVjqfPUogKFyEvYiuHItRxnzQJhE5JGGy+NDR2/Ensb8JnvU+aAFm2B
pHI77sj6XeaEPBvsOmsm3nwGd7ZGa00P9JvN+jgk6FVGM9r2zvzHw4kmSE3kR2gF3I+98ePnJWXj
l+2KaEh/KfI7c0yUqcU7DiyXfjs5T0vsJawXScB7vyHtXwmZEWJAwYT5pXR7fKa/fRFkbhWf0+gF
DyGEZKWPFXEwVA5HZDotIbKJ05rldqYAQ4y11lg5Zpqn34EAdV1VkHLruFKifngTIZz3RVT8X6EY
6H6HMkEdwq3isY+KUNqaBv48DF1BW1R7ImQt9fQAPyMeJBysFfAtpPeYCJUaSHBoHWl4w/ZWx69c
IXbWmVrXVJlHMt5Gy3npafE8I+RR5xNUrBHFWGgr7Ju0U55s+Zo9mjGdUfNIViJgYAh/D6N7RW9Z
1HZR1GX20VKnIWbuPs9zhYbHA/OkjgzBN0JynWcJz6x5kcKP1RnnBJZ4X6h8RNwdo8EI9UzeA4kS
JbPYbIFD8UAd6OhaV4os1s36LPbF7YDLx7y68fZ06aoRCu6wBEttULZCVec5iLF6ZNFgOw/GLV3m
uiIDkVuygoKtFnHG9ObAIGIvf5xnUlgxef25ohpBbS4OukfCbdf0A1/Nykpw1CtYHHE6IQGcTf41
3OnpYbGVy+njTThoSEcWAwS/TTHv4HaGisduYwWE+cWGKSXk00rWdo3T5zXuV8t0BYslO/mFBjuT
VVUe8uSruvcy9EihySZOS2ybi1LirPgrVHawmyit5aLEynuHDqJVZUGbVF3pWdbpqRzTgDNNQw+G
LZDHFxHhSa6v9A4sStPWoAkQja1QKm8P1/WWr5YRrZLsaYAHUrPVsUcKH743wCqN6eqpexlTOhVk
49+yeaLCrMNJcbaV4EQz5WGhHWyNdv/RizIAMV1J/zfDAyjdNoK0IuOdjzK/tjMKJVJic2DrOxm7
uczM78UQetmVv2iVgZKuxoc4XVY1ieWu7X14wD3UuY8OMi8lcdDxbjgG2af+Hiu5jsRujTnFjyZg
5ecBpqmOJVK28dhUk42xMpz/STkfTUoaBxN4qyqnVdjGdY8dAouCVO6AYfr2N0kRSnxAFsoQRoI2
Gu+dXot15cgt+QEwYG6gQYnTJzRpfzPptu8Ac4gjgPN2dqr052LfLgjzpdk+9KXiHMpnrLskeMw5
oMSTTrA6zuggTeEf+0xzqEtjmXz4XtBO4v3VGDeHDsbes/lNx58w5tzABF704LjTy5cbqKZBAwhK
CGbGSnHXCudk2AGdYM3yNgKM5pz8YUX7JxbHGuDBmfuAqzkkXArWA1TuR2ZTQXr7+sJ9Qy9ZeFFg
BQ3oCr2a+V2WWkx76dPDe5RgHUm+Ez2/I/szPMe6uCqUT8XzyMfxz51NuG/g0OVwqCRfBuip4eAD
nSr4lU3AEPVRJY/awPNiBIi+Ldr+qhg37Q+JxubrTrH68oSlGpvqEMrqurLfB2ImyYxC/TxgVcMu
t11tv20ArIih4yC7n+ZY14C6LAsSw2QiKqSjUxONzL5Py6Df/vPsymftjB2bsHLeRXUI3Ocy0X/d
e0gh4ZIxPB5ikOWqZ8ncKHhjEzZ9sRPSFxB31fJ7WVJlbxqvndUb3RU8tHPOO5qxGGWqHDnSBOan
IG3/8MrJdIF623E7v7Q049sJvNhmeGCRVp5Xd1lvMoKdk1I5R/lgxVPz3LBiDCHFxcWYnZQuCxIY
4mpPfooTOG7K6jP19fK/pRZ8EqXny2rgHZTP/LJ4vHiTS1fMvEJZH6qaj4+uvfnKIlHEg8OSpO23
DPcgre9eT+DvGniwohG6Gld06vHcH9ByqzxRVa3DAi7lKYLMH/44hWI8cd0HmAP2soNw1wVWqYGw
wumG0g5cwl9J0qlpDlVONVG3IECvcLtxAkFL35uwjfa7X5Ga0Tgx5S8q6Aw879Fu0AhIWfKmDuB5
FgzBlwOUp9lzppLEC9DpQcYS6gS7sTbZ1i3ARAq+xpaQ2LXSS053bvW9dHuHe02w21EhFK9DRysy
yamuGoJtnKF8CNxtuCtybCbHQ6xrCWAh57A863oKWTaRLPU0U1TaVDfAcw1l5cZ0PaRFcbNz2ojH
T+F/wR0On+kx/LSqBhcbfji6a01dxc8V2CJlHN8Va0b7XRZEjtrerqQP8T71zXaP6W3Plod6X/Kk
5v2MZNNZAyhYXUtLMV0PpOrPgGvR+tBAd5RgkdtoI4f4o9nqp8+ypWJLUxBkRz1MY1/wkhzX+8y2
7BI/DlVdkLq4Po7SFz54RECxDm5NwMT2SakfDEGcp+Qhplxkb2Ky/CeYIsWP5bZsgqtEXlwooxtM
5qN+8wbA6HERn0FDfg8BTlVA9+fx5dRL1JspR5uaF1eHQrdHohBWYpsOLPvUKPOn/OdWeHA/JMza
/SdczvzkYFKBbb/ayS558PtyFF4b6Lyp6fg2mVqCixYspO/lXGvyupiGcY2qL6MidBTh6o5kdBLC
ynB07+PIZquxnDIvlQk2wK6YR/GBl383mEQNHB+CC5ttLzZwbUe8XLGyu9oM6sp1GsWv7rV0MwpM
yqjg0IEpuoCBWKlomMkFExGQwCbAU3rsJFvcabzltCF4o7Bl5YR6Wm3zjq5dssP4pQ5zXhgRhR0S
1BNrE09LUvfZxwtK5Px2OjuKzb9ol9j3n7hKOzSy1I1KLvHXhED8tZPkm6sv9PnUQBhbq9pWgeX9
w1JTLGPPFv4KMx7q3HXjQW9Ws0BHFAj/DjqI2mGh7eOImcvAiOZlQo7HOF4odnEFdN3AbYYYxh6m
ZCrDkhQyq3bX+CvzLUsStMfT+7JNaRlxc1f99GPc8NFHJrzKJ4W01Za4Mclf8jj+GysNYFodcqJA
TyNJB/Z1YW6x3Ym0TAP61KMr6TD4dHNO/ONYeuO7PTvRfrlZ6d/9t13f23SwYJa1jOgGV29ZjwI5
AutrHGDhw0NClWqXw3MsXlFK6MXOmTjUQlUH3wDLGWteITFpEwjWM4knp1ZuN1CKJGwJv0ufx2LB
+P0w4CDZiZuSCuHfPkmU6/Z3pBr4YEmqWhgAFzt30fmuR5tPSwBS2ZYwff7xCZBKQ/i804Iz+Lr4
WMx9m/rqW8JJuc3NHFvE7BT5+wSf97tQqGGHe6N56/ZgTAyJlMf3FZ7/s5csPUy0g/O2MJYlR2B+
PsfxzsmL3WaW2KWg6xhbTJABMkZwrSEWPku1fApIP9bYwIKWebvgs49VQhRmKHsAYqF19LsbpPyu
tzzhs2DiHcQ2GI9/nznkzWftxTb42wjorUlyQyRHzxHPw79ybAfmAMBKaaJt2mrwy5EhDNUqvo4g
JLzx15Qi+g31hPDzck3keAwmGDJEzpUAyUNbgcKf1TWcQj320viM4grQ52L06T9Rx2+WLogxEm4D
Pn77EOU3DRZP3Ejc1lQfpakTp31MZj18Sfb7i4l39NUoKIlLBj/6W6jzkmNMaircCMWtHlTNQ6ub
Ridtyz5lEyTFkPUpWEWqG/YK7p7Y8KCgFo6drvgKOBJP42y92/DiutE+JWTQmcC3EEjj5WgNeTMy
IVgiFe9tnbNCE5ENy6lu1xxtYbisYbjYo2b4R6I5Nbo90zD5UmDQMak3eWSxdpJxDEAz+YNiA9py
eLM2aJ13KR1ZPCwxd8iaU0HFO1O07I1fTDWQ/rfHkjxw9hnk4irEalzutBjScaMGiDyMOllP4Avk
gT6Z2A1K/0sDv8IisLwvSSqJHug65Zb7g39w/sd6D8WuG6FgDQzayJf1f+lG2NlGGLbLKC9hL9TY
d1S+mBjnK2Ou2kPY/I/FeLueY6+QMhpQkxfwTul4+CEtIxl62vHajadVgTV0LimU2R77OLqyC/co
gcO+MMe5DCnV/M3ukIUHRmWWrTtccYewQ8aN0rNH8qDphhOIwS5cT8D+79ZAhh/VRuPs7bTOOMkh
UzHFj2b0CC2QTZIMRftXSYn3Pbej1PavYPcXGNV3j/eatoOnALkiVXv3gXDKDmCVEvScRXL5R+zj
dvnTwpn6KZWsrxgOV9QDU2w7kLOHMHZgBomgQ1bSk2jhPG8T3EbWZzIsLEJvitiOJnptTNXjE7IW
005Go6n4LUKYEz2Vr8acJopuXxWEYSBTZ7LddwD2fQSiCzQhpV0UdkH7v/rVGbcoTN7MrAL/SbA6
iZuDD1uh7cWHry5B9jUVeHgExzH1nG8ssHur1vdeK21n7k61+ZcdM/c6bkYMmfmm7a2v61Rwid+j
dtp93/GlDN1XxAbg93+MMS7/GOxPaeFoeF8kntoF+pEDqCS938Hx4epGxoP2WlRyvz/DaujhkiUz
qmH4+nh8NQMnp40PIUhz8Tr7F7EZnz8EXg+XMUqBMtm/42O1EfNCyffWb/qgeKUScaLCx3j3lIXv
SYnqRm/cn5mdmG8ap1ZOAVCeSwcoWpzvPzLh1EMnc9pBbLUXr1+Zm/69nmMXbZ1FOuAR5pg1XUyT
byxYOVdVneVQ7hNethgI/2xRb07Zgty8HtkrnwLNkJsIMRR/2/q17T2ju2LJBBa2l91zx1Hvq5R9
BzdpbkHqUjgDxKYcZQ3qiPoccQVL1W/xGBBRheAKfGEzE5D7Un+jDjf1ASa397r9bundbC3EY8q2
MVhO1/PaqjZdRyHbyaySWhfU4tT1iBwuFaEC8cJtoqENxP81pc7RitMXnDmcqt4A1dVA3UzUv/63
9f2yk6zCEm4c3bT/QFzcb3WtDwzg1aCQN/ujpMrTNWRlFdKh+hon3zn2q75/+BhzOx81bcEMHQor
9vtL6ZX1fk1XkcSzdFAvl42T7/ZRJV/er+p6yWyVqbcja1Hw6V+MToQ42d9/PKsM5RQkGPi2XQVA
skcyWA2hPjT9mdo+qRarRUNa45YyOr6YyBRvuxSohThp1Zk5W/HG1eii9cj1gwNQ8NdZ0rkaMGuO
cBPaXr0J8GLPcjei95ovJV/vudPNxYRtSmaHm+RrkcJT+hm1Vxg/YwXjNcrTx+iqQP9z1iwVaHNh
tjlG88WvnrdpkZSnyPZGNRSLblP5nIN2HmTUoXrKbvrnpEs3Pq0jcyfwVsbU4iDSfW5OWoT6ODQJ
oIwBau5EoyZIf3dsDUC7xt/MV77CMTyVWus4vpB6AKHqiWD+jCSlvD2x5GzrhZBvzRoit+o8xFDf
N6z1nXoOW0BlOBDkM3If5ABZVb8k4eba+7cb8KSyi32HVjRj3HDLiRDRwPN7VP0vHgWOhCJSiUA+
QkVDlgMe5rPgfOPvgMHO13bX59J4eh9xICikhC0fRHFtrHeDrvwiZ0MhGjkQcksfM0GNjbt4+pIU
lKQDO5lHtT8DCNdCvOwLNKonQpGy8zX4VYXPCtZJ2EMXCYJQ56fj8W5vKmWVwYdqHDgDeLdQf5Jj
z8p3CYbyr58IzHMa4Ivm3lb0mc4WkIr6ECLglOkfYpF2jucwi2woc51KuTpvT9vi42X5j9NUn2sA
4SkP+CSwMIeZN/wb1hBa7/zeV/HIgyCWNueWiGRSYBW9XjA9+MMtt87ulGA7okp/DJGIX4sG9ncK
Q4w2n1XtayqSy8RvahmV4sppwFSzLGaMamAGvtgHBHwDn9z3oBTGH7eIU3tYsdeUADuauJ+y0x12
+hy66A1WAvu7RREGg2V/chW67WxWYha3kgDB1OKkTLc74rnFDjLbsV0HqkSNE/feTdOenzkaRlcr
f17v882Tp+m6Wr/GBH6xrw5pU+li7A11NbBJy94BjeFPdRxkrlRuweNHZCNyk187qXPaXNA2WNlO
dZAV38ELWZ/zGIE2ggBGEFa0dnxN2ryG+hFmhoDunOPOkiyV/AmBCcHj478E+mLV7PzR97HjdbBD
Yy7wA15faqYDJ/TUuXZUfz2+htNFVvSe4pp/N/i8cmbKmO6cicE5U+LHpT7qGRB0xoYApkNu5EXB
aikHV1R8FJU59jfBF27f1xLrI0q5rQqPOdzUVI+/ejjlsPQLljvClAO7hI3sr6HyVIoDaKJdjdjX
MZvk7X6W6OQhUvClHBGmu0b5gxRP+9VQqHdVRc5NeVyrX1Vulbt8BL1KlMxALv8jiUWkORy5kQWm
2hcseb31DIHntM+OkoUnqm62Nkq5Hir5T9kfaTrwW4xB16e148Z/5UyZLZ7HMVXwe+WEdEu4oNM+
5JmDJXIIt0wlavXsDR5l6o+WkGuFJtgSuJ89UIdWFiq4sSrKDkizL5Ql71O5XbI/YITcZjxMMMN1
ktZs5XFzMmk0VyhvDspxyjwOQ5K3WKS0wtgodeVqVcboLDWnIhG5E2RJFvST6arYkes+3rPDSFk9
y5wkMaaNPGOD6bvuWuC5XpKuAT8BeyQDU1S2ij0x0O2pV4vEzJY+bcr9EDuqEvJd260oXItpm3HV
096+hr7YHUuStjyDG5PcAcNYR9cklcunz91SWatWw3RAmQwfM8fAxpVy3EugSeo3hYsQ2TdnRQZk
qS0YBbK5WAMS6VvkdZgmGLrIjjHYZAqGTYLeCc0PJ42hb4NvE/PJEqI//trnj2sBAb4BVjxIXN2V
zuOKyg3RzY0AkaRwDZFDxgq2CqyTmoK8PQY94uhB9iKYJWHz/UZWAtqI0OM0bnGOQO3nclGRDsSq
OUnbsedD7uGl8g7t6VFa1fcZbGyWS17a3o3KOnhbz70qAlZJs36iH8wFUoPNPy2ILvLsgCfGCqxS
ObR46pFqYYkWx852jd1n4svNLEw+IqczFR/wN/UVLR6WOnHQcZd6qORst8k5qeCx0gt0qTGOBO+6
d1fnG3l1z5hCq51+FvDdQZShsnFhe0KrMydM9E/avZ97Lceuf3E9G/3Ppl9IEy5edlEixaoIcVsh
41e3cdH8hMvxYzmvRVnyQ4lN8xM3Y1VlPcFFQ4jzFigfa09LizkYlXpEfnHAjzpUB0FYuTqFo9XQ
ZQrclU7XoT+wmjucgcFfXQeoPY5P8J5USL1/QG4Y7M/NlxrVAcXyCEPydqNRhh/YTZhlFWtmm7O+
/fcxOhcccOBnBOlNBkKWyj38OChY5JOe6Xw89uklSnyxeyUmiMJXeMuO+RDarsCFtnT6fSJqMR9c
I3gFjEXotSki+W4VWHtyyT6QVkeeVAe6dMKcnD0SRTLqCnqW+INxoqUMEov+0i8+6p2pUScDjWYx
k1cVtfYhLjBttf/gOSVcPx6sf00SKAx9/r2MnPDDemAzSPAqXWJx/6foQpa7LfBjfiNz7upKJaXT
nyyHKIavJ7jYbNW8D4ajOLBHi2Wb/dSTSyTFPfob1FTKIOxmSI1WHGWF2ugu7T/YXYw1lzdMxW8b
DYcpj9vQp+kpFyLEkRKEUtdx7W3S8mWLK9Z/jfN1C7OgyhXGIyG7kzSyawADekJ5kJMZ8nsNrqEW
30PeUZ7ehmsQSO28Htv7yfypme5IbnzSfpMV4CVV+MWXSOOm5kvEbUp5ejMreZkbcRzlMPGXpBGB
2+bUPWeY2OSmBz/PDxMwAOmAqi45udRpJMqel7fSw/U5Gr8ULyPdQfDU3F6BRVVYWZnlejTMF2dv
mrFg/ScgqoznTyOw6QIHxqdmWpCNmhM6nnH1TjyJmPZR/W00B0brFT9RH/7eF3k4ylBXjHh5LsTE
+RUDTeKvzk31wUIPsf5A7a/mw4Zs1QVPM/evotudLvI6cnrBcGigmscFE2zzMsuzPPtvM6LLpVSY
QIEyl4mys0nyEwt29x4S6yt4SQINsCn20thBZZ8qKn5Lwe0nEh7sjWsib1nunxy74REQZONPXvL4
rrBsO3RLwmr7HqsT0MhiOv3X1WHYOGcC9zrSld6K8jiaQIM3y2Nh/yhjGaOc2XyzCh+b7wFLNmYL
7Iy+9Uodpr1CDGxLQjttMug48BifT7s/ioSD3r9TOEG0ROkXkHN8A1fkdCznfVuFq4DkdfamJpF0
y9iilXer8FS7FQMBCmv0FaPJB4vZXTALX+K6Ns4gLGflaID48LyP0s+dH7dh1mTs0UIcmkGDvfVB
GZqxBL/ejcWxdgwTHuGTGy6ldHbCwmIxuCFnakBgIJJ9h+cplaSmA7J6tUXowFvhJWTjapihke4G
2bBI+jloQPFm9W/A7o/8d5Cx75+zAJYBtaNocPBIejyofDdyNF94qId8yakCf7TS/qqU6iT9F3HG
PLh4DKyQUCHljBZXAstYfYJyBgSQw2HWLrPoJAbUZ6V0TqDIvwFE+X4MEJPgy45ApQscQSD0RNdn
ezzTZj3MCHLeXiK8fCjzSTKoo4Vi8015w+4aHBFbevlbq4b+tBcbsNThQJC7izLTMD+DS7a+vl+/
57vpvmVXaYjjy0vELeHfEN7lJGJnBvCbBPkuiZEc4TE50iasq148Ad1YbGoT8+eWNdItxoV1RQUM
yFfnQqPsxijHJLwsuyCtwq0sgcfhjXtD9/r1ZOrJN4MpDAPh/IlYZr9xede3jjAjTG4TxPXmV0QO
Jg8tLr/y55PzfCgZNUrvd0ujVROggtzizR5JbhtYmVMp/vrUJWKEBRJCAb2gwwDrO460boFPwEZw
yQNoEuR3QnD8Z5hQTkbCwinRrKYMpYTjKQ81R01T0cm1pLvFsyusOdZmDxglz32sXPYtnkm7V6Ho
HtbQJxsKo9oV68TJJaj1dZs+ZVGfDozoqKLNwBbqYRfy68W4gxiACXB0M4vdaa1BEGBf9GSXFOm4
cwgjhE9B0+AuiYj3BNmt7HR8p5BNBQD0Op75hNRN+qxGYIcnbkS6/beChahT+lo/W+ZdxuMrmwgn
/oJfFLbJMHRpi6UacXXgOWaH/fJvFswzWBExwwihZBnn9DClqKrmWdFbvYxNEpNrIdRmShOeRQqK
Ha0EZXvqFtDVmQFH/9fUqY3TE1Rpz65RTsLNef9zbB5OOoDJQS66TEd9J8Kelq7GvIoJxjtF2GSx
vyQvfSrb6Nf5zk7G9RWWy5StZrc4G+HdEGaKY83b/eR8gELElfjFvm4t2WxXDuL0LQm5mBDBftlJ
dPN7QtOtGs/q/CMjV7BjMCDudLkmNmWhxrQziUc+F9VjVQfa2Di7pwzzlX0YpPFRbI6fIuJ6ljXn
evTLjsHqK/vARbLkIBYsDzv/XPuquJT46o/2XyhFc5/wAtg//9uLDqTydR6uBq4ev9wNYkpjClgQ
C+dxsND3cR3Ym3fL/4oz7b46eQDNjIPOJwgjmJMkMTs8BhWMm+aqM1KVNM/nUHpsAC/SCR9ZQVvs
HRQQbFsbOKBuHfdZoGpeiAuiWJTmUs7J1NEuYsIsO3rPXmPlgSSnh4YVtDJi2My1+Whb8cCEmQ+E
cQxweVutW/BEBdx6XGbEQRCKOrRjjV5qBBL+sCjpT+JtMgMpaEToAIymvDjwoC2+ZXHtj+w5MCJn
dW/7J2+8+M+S+WL7DZzC1gk0UTmA3+7shSTBzPOngkYoBtMpvFyBHU6X05eyvbUipBje/6NuWQoH
D9igAgUntIhGAI3S9UskSG+AS8omodhtl3KAXJS5EcFxvbQY0oA5U/J4Q85Q2YGKocJ2Qz4EvQmW
qsdRzMZHZaoP7O2rk6Eu9wmGU4WCAItF8pO3DGhDahulNxAB5nYbEyPeaYTezQ7GPHLQqaQAZ6eG
0Tkb8z72qngpZEWembwa+t+nIMoGX88ypPG2ZSmZQ1CvcIzno4WMh+9V+spgx4ANIAxdGRTu4TKx
V9IpbR/ApxABCJwhgHMeOxpgHX5EoDhf2WT4k352BPOJ7bneH+AIUAS1At9i6ws91VPwVndMG8Pr
hPHL+gZVmdqFuwmnaV18oYpw0U7RQVuBnMYbkHTnQvDeTizE19pLt19UC/8Ze2gF35UBYVlfWUt2
xVore+/rHrVKmZMF9BoXwy+NpeQGXxyeSME419TEmD8+l3t97ntHvzMZNtjOWGWzZiR0XjMEx88R
U3T6Ft1yn1Xz22wnMLTizaEUDf2lnc62pQ/DUbx7NhJa21QOSTLF9XbPOVwWv7208rFXWLdU2kXs
PD3r5FEg5DCz+G4W94GoiT1eISWNyaMC6QZqpq7ThvNHsg/lIMylgcXyHkVgL1ZM48IjX+KcuVS3
PtjlvrYHIDSFgNry+ALgaJstjPgL9VX+zV6S6W4AOd52JS/k0CcI8ndahmAeOJHxAg0tmteD3wwK
I7mhFBwP/xu76ausP5qY+KKpGY8zq7VEuisyf9QQweBtRm/y/IZ+Cn8H9ObSO0upmwh792uN650F
LqLeqAfTjk8hnYuKinzpVemohqdKl+sjL7lAcbj0Rt+TN4aMs0DXNWG0LWGj7FRRPv8QR/vYWTf0
9zIwAK3RD2WAqSqa2j5A6D4kNj3wUJWHcr6Q3VyPZCQNX5LXmx1Md1F3BF4TQaRm7cl5Ue68205c
nd78PKPAvuv17IEYs06O/3UuyalWSMZBx4Kfqk6W0lsT8t607+YvS5qiGWX2oDzt0visEQ8EaDeU
93yl8gYjiwrRvbSSPJoDYDdVDGXxyMpdk85FaqPhNUNqIgFKr5juIrsttZaxBbhinzrF1jCJVBqU
Z9/O0TlqL3Ikj3DwMhvn45n+kUZgycG8exCDHCpyTEU+j9BtQ+JamxUdtgJ5I+epgXxASN2QQXwl
/94GAbtEYIvpj+yAm4t5yYMi/8ZdAcQDnoPgApVYIT2m3ScFLeNeddg+xCiZLVYLsByPKClUhm3J
Jp+sXhxWbp6b6daGRp9/uO8pibZNXm7QQJpm60SKoUPlZBRqRMcjXDYzidD8d2Mh3Uuc1KkULkqP
1ySNAXsTJfVWz5jCmaH3hW1JC+N0eGRVNg6CX4yyPI4LYd2Wunmqw9aUwYZl/BxhcV+mPould0s2
kO0fuyAGpT0cDAqofGaI5Rh7E6H8lsz9yhTjEduz/8XXrORC+5Sukd4OF32MrukdQD4HWzs2r7KE
Fi0/lceAdUGSnoTOxvmH5vu2yFkBiDaELadc/at9jaJiySsvs2IPIvLnXuBOhx9OajwwfQX/t6OA
Daafhdk+cmyDm4CveqNIVJD/e+XoBO82AVXsrsIztGUoHgtLQ8h2gO9uuD0y3KidA8DLTPQmGKc2
eY+iL3vaE6yzZGDJpztHpiiCdgOSIL/C3mv/7TangBJx+LfjQsb+VeeDIlESKebnK7ArCfJRpKe9
LEngau6Fwz5Lxb/+DPOYHT+TUz9JtbrUcneNEqQN1ijPxwBw1ySU0iYJd2y0p2TvxpC/k+ZGjMLP
qnAiLpweHop1BN6mxWatBxxWwAB20A3XjDUlXZ+0Ae4Wfs39A8fIzystSkWw8uInVg/J9aH4scoy
5NkTq4lSFRNbPvDtE8yJKii3iPTnAvuZBKXRoRdtPCdPrWm9/cGE9Rlz1+k2uqr6feihp12kURMQ
w2CbmMmBRxND8VqrZXZE92qfAFc1TGpOdUGiv54oC1QBX9QUpaFpcsAPrh8MN9RxRTPHuFonlM5o
3y/INwZNCSkR5S6t73y6Dx/SbSLHpoo1Xl6lm1Gn4trL/ph8UOIvSR/LOSMFIeW371j0qJaQD3um
FSsxzxBEJ/L9OUO5ZrAkWkKQnnkzkDuxx/HESoiYIaB/9Ll528wxRhLHloTyNIQF+9szPpxujtl6
LfTDgcp7kGqBROAVE2yIqso04xwTf32rxAZVUQwqt5WR0fvrwOCfjDELFWzLrNVsOw6vfWZujbLB
mvKT+VBn3a9L5rXCod59LJY+glIjptS1T2GZ5WOQN22Xb0en3hZRePAueq9fWJTKRgyxxUZjgvDa
+p0t4dbzxsNX/AMY+fOP5vPqTHfDOROPlgAbNDTqsYE/4Rimj6m4K+rZZVXboWCJWVjyoA2eFP1+
nGd6LsW2U4axkF4boylfelEF4dIn51iEa8pZpDMqRf6GCNcb4424TmT41lcsQ5cVPWV03S5NAnng
bW74ZORtzHp3avBwm6glr/gvfh/zBboLc8QBpeLoltQ7pCGOrtw+n7PlcsVSRi6TEICo//P0bS53
hQGE6VTydczc3qbCQVCid0BeWNKCHv99Jcueg1lrVVaq+Amu/JHrVMu4DtLQ6eGSO7LrF6x+AFrV
AiY/p2sjlpediTpVQeZanlQKIIzCroINfsSwzoR/TpSms8fMkYD1sQakd/pQTSZFMr3F6AWAIao8
LsHSGsmJkK/AxkiLNSsIxwisHPp7tXkj5FtkxRaySyiIcBTJtndl09aiWRgXzp2y5O28pUiBJyk/
mOfAhQgllPwTp1e6mN/kYsxHNT0PlawS7iTpb8OdSlFpI5c3QNJN+nbZUKGrVjhWEQlaJjNWUdKr
oagzwSDoAhwjjfOs8ovs6SPw6rnKCmrU4psy9q6m0EdYlpkNMNMxPUzSMeKa4bjVirPfUaW1QkaF
kOasdXuGSWR/O5TPgqchHiNh2VcUm1knhpltskyKxTaVRoZwkatfZvc2ag62zsqibLXH7IdGdkWW
bu+zBBMYeIl6CThx6PbbUoZWiOIfQJk3YiVAmUmW9fxDbgE2KwpSeY1bg4heNRU4oodrgt4xMllD
pECCa3hAmtcNq5FZAT/R7p6HbtQIF8HR2Cf8BOO5tUoevBfrRuX/lyAK0ydTDXln2tX3q1yX+RUV
vC3YcnFKQQWBfP2hgWIS5HJt2EvEdTjE7jbM4VfsskkjrsxcCqfQVpBfsP5Lnu8bMmSjITo3m4nM
Ju0I1jAywb5meem+1rx6nGC1h/KbgN6BQ+T8C6NE17yTm7XQI/P6LJtHE1VYwfhVHHvKHta2KQWn
nF+RIVJSV6amJLbsyZNT+mDI+wwRuSDjt6Y3O2G3DG6+L6URRv8TN7rHog6rHhw27lf2fOGkE/SC
Sl76/NTIAzvVTpO27tWxzcl3Dn6UshnYGJnDXki3ksV92zpwYOQKTHd+oVoQW5bVP+rCm1CodG2q
gkEZOIQb+HaXxgOFWX+WvYL8VI1hK7qp3u1SF7FaI/sysNEIQ4jMUPV7KhFVkNz3toXpZ09YRh1g
mHSDDFmMZvNHJCcLzUrVYwXCxMwJF7EvCW+854+lHl7sGQ077RWaFmcufPSEeu6Y1bPbfvHJLHRh
RnHaaYFdajyPIJ68LguDu3+MSSASpvkwh8QHw4/KnA1NLMpYAorDtoA7eHcLr91jZxfgOjxY1HFp
0qVBI6sWfWfdsxith+e1SDpHoG5JvwZhvnxSKM25rMNqZOceTQZQiDxVh8mU8JZZi8IW8vc703u/
6ygrg0iCUjDyDdBTP6i4l8UKDSiaV1TPZO4V0QLYlL56gfa2Tpa4DRL80Cy459f7VYZ4DTdLl2GP
fEd0o2gvKNaAmShCmr+ohF1DWrSvVvIUJGzIpI0omVz4k4R3PutqwaTT5rKkf63WOu8gLsti8Vfw
NERwtMMqolR6u+WKkHGHcquBtj2tlJxZKB4VxleGeSeb3M9Uj43qLbXDpJfUR4R9tNXXQ3rwofvf
rQHzGo5TR0dLvQynp55v4cLD1wddtKtrk1ZbtQJel9vbdp5roKzXDnwyKgdjE2bLaShKkCh3+wgh
cLdlAQoqkBB3SiP84ThCyQlYYrhIz/bWeCyMfMZVPpyvbr4Zd5tfSDeJyxWYIUgKZj9mxo6U5xCh
RogSWc44z454M87TZ3PjgywJaZ3WQXV8PSjMo+inrm2MOBNxKN83LtcRlvFzR28N6aY3GUV/SW6M
81u9ZrX2Za+TDchmoWc20UKOfaaSYcN2Koqu2i9+WMfduF0VjKUm08j33Sq7S1chUHEaisLwEU/t
FXf5yO4XfxNRtRH+DBCmINImRyP/awTJDFC9MV/vtCcQD1D9twMjI1Lefn/WRQjsc5PC/jQBIcFJ
uzPzgSQDyiCJ7oJbjnkVMIlPMeecKv+v6LEM5gm/iVrqs/dSB2UFlCL8EP5M9UT8GLYO+8NcLHZz
YWWoH+G5zRW9QRToASPXdzlcTStLLT93F2jLsJ8BA6syLaoAiY3C/FD/6E8uBo/pMf35lGyXf5at
IY3rHUnp0CuIKhc98nm0B/TBeRleKG90warkhYYe3SULzuAq5FvKTczDn/u2VdosD6qlpWXVtg77
/8ikgOR8jtxSaMZnkikx0CLV2IBlG7vpJ9cxZ6Gx7JFeZ+rm1k9+tMRZ/BIXMsPyb0Cp8z/bZ+Dv
56a6h97MriFsgzlj9r6SY2ORbQ5oWgmESM1O8M6msp0vr2VJ8ZEEFaXRinL/q4ODmeiJRQsSLvR9
AxMA7NJrJbi4Aq3m/8oeGS7C+2hyG+QCcdgn70vgLHSGezfoa/3kh/hxh5wnpRsKNqMSJw1s+8OP
z65pFFOe4Ls7PYb0T9aKKtvLds9eJf5OaxTY403fRt66Kpah6biqbeilwCn8h9AKq0//X2NybBaG
RXDpnDZgQIldqNvJm2lnwM4xN+hzQXwGdXUWJsaCoWZsyzypTSQTrFiomx1HC2DUMOXG3AC2FxAl
VobXzpw/rgZtsjI6O0k6g+vpPUxZk/I+gXhzE/zadpQl59kwtGrOxjZn3XugbHxcnMtviVj75CYO
+4Hxb1/Zr+5tU/BiqBFyMckD5nmfJB/Rx+aWiQN0Vb6M11imdYmuRp+HpU7a4fT9TqIZe2t2lhdt
LTwUo+jWRPVS3GpvFP5aU3P4bATwJwDH9UOk8cWFNLwNza3SHgsci5Lc64bdae3EIrTPes3HOYww
qOcW/o8jDRMH6DToy5IuKSeka0lSzp3v7yfj4lZHjuBQNzx9H3v/UgJFJiBgWC2fV2meyL8I7p9v
Wn7ajQZ10GdWG/JclBd7pc/yija88159Hg+UxmC9PbqU2wF78uOA3Xs8xdnX9Q6JEwTnhxTwayzR
zhN7aItZDX3FPbBQ+Zdej+OplGVpZ9IGebklWHoSCTVa2t+R6C30BwgyM3t4CVYeZEsdL1Fs/irV
UCDvcT/xMETRIeHmwQ7pFL6/XV10eH2EQ0MNMu9jPoMCHjlxJWFvydD1gNoqSl1ahuxX5R8mZ1YT
0CBcvaV3NQCkrp+bkNeJ4aHn/y5Q//5ZXXEmOL4RGWCZ6a+5k1bdo/AV2MFeoAZxAHGU7PmEojOH
vlaKtZm0wsLMy9ouVzWAFRorOn6AlSdMOrV1IwDnDurQd0gihla+32kboCGBgaDgsFvxli8r5DDf
1npwhUvEnb4k65+NsOx6xcscglt4q0PRs6SOmZ8y2ultkWViNu4VT0Mfiq9E4hZhvvfbb0N23zzL
tsqi/E1C9nvA4Osp9CcBOE9r9CyetcicmKBXxP5CQ+krn3AKZvCKf3JyFwfvG5cQuQFjL53uk/E8
FxhYBOqrOyNFRLYpmLyXgXNpBfbpmkmbpV8EDFsemmhBjV1HJxR/BiUKpFgJLCpC4Ys9kefnY3+z
/Q7EJwSm4RSmGGlXRTX+B+aNSVVYqOq2kIbWzyWhBNyPHUIJHT7qkInKYlfC0cR7dp4NxA60R6Q4
3h4V42D0rI8V2JzfWfupji1Oo4R4f7mAglPWHJtdXHVb4tsje7cj6c4V7+7XEnj4eZdDNConTQJH
u5rP1negcRTSFCFSPM0Vs5iaaBbVJ1O83AUf3iBf3yNOiTojWfySvPp9nogZmok+lNJrQnPghctw
hjLgLZENycA8b1Cx1kv7EkGsXJJM68mJZUi/8p73ivOVdtIq7J6gX8ODePea4tQLOAU44yOCgviq
lNCW2HIjh2yTK+306H7/iXVWBTfaJia9m7q4E49LPhR2h5e0CVC6K38lHNVW1rnqlaJsQakZPuTg
pe5FVviufu5Az9HsHHm5Sd5Yhv0Yad+cx7kff1q/SexB+agacGIM417bobyARrKHi+wc7SWL7LF5
RxLyCmratpn84e/xoFmw3NQsz8y4+p3CB+ke8g8IUGDH08qPRPcfk0zq8FEK6KQLk6UgFKxUYYyG
WxPX1lriv1kyHwkGAwjn0FVn6hqfe+uGNNAAbGDylkuAqbT+tZ94NV16DREU5aGz/OSYBO8gxhES
xDH6Tlz94L8zLcvhpvffnSndW8ZsfDrMNH+eE7ZB6CUZPLUFTWHUmwqUT/LusWFc2Tmme/pyfGQi
tKIQvWz/v4LBCj36Oo4/DSAaSvG6CifjQYiBTMNF9d1XVsvAgxTzZlw6eFvHGCKRPdZIZFk6J+rd
3PoVUvn5Ebifry6zHSyCR7D4ctvjIAbbY3bLYVze4K3vox6uEo33U6RjkjxBMuPKi9OZ5DC5LEu8
qVUBxINqrRupRfjGkHZYmhPCZzoZpXC1Y4yjbUjaOii056LyYq+2uubZC01mH43L8b+1GWMA4Brb
2ULlfbSLVHWN38obvyl0+t8v3dOymQNpCTaYCoIhrJJ5idC3n6DliTa/sm2gfV3w6X3oB6PyLIQR
jh202D38JfvTQml/4gCASCXrKh0/9YqplnzU0V1KR5TFwB6JR4xNfBAyaKaGz2EASaRCUa7FaHEy
+oqxnQUBus4S6oLeTtXU+1F5jFi9DdjMw78I8ZM5NabK+Vpe4VPkX1EsoP9pCex3+cdkySlu+oe3
fZWx3k0S2IW9TOS9Ia1wB1WzsVrh+LKU0z3VWYyexekikAa9KHzUTYQNITmk6BjR05hyBllm4Efd
spvJL5McyRNHWoLMP2be7IZykeVnplkuycJAASwo5vHuFzzUEefszS8OPYsnnQPz94FYOZOBL0PO
O9ZfvdSpmXNCSrTK5gn5c8jEeCP4EIkcw7Aux7OPJkFjD0416KgQbJdaclpoLFCapE0lY4imaCCa
Wzn0fDvGlgBNOxvHLbUTqJ4J9Vusp/myxJOM6r8DQvBJ06QKSWZtWv8iO+31h0NSSQm7JcQYmpx8
8D1ZboLDzuM5cg7RJXTWHYYSjqJXnt0Gw468FyGErtZzGFAuenzcM0IcZo6hQLSsGYUyOeTCutSQ
HQroYZx6roFKWlOyi+h7pPhquGx5cEvFDCZJ3pCAMU2Q+fJwzjxq3aDiRexbikD44Kc/4f0jk58g
LZf3O57kQFcxi3hoia5Bvkd/Vplxp6hNkXC2Fe6ql0YLucOJvpblh1eQnb1lS5ws4H8rQxnVBQUE
Qc9Fm9aHDQXimmlPF2wsGu7oaLCWlIZFfB/tfdP+Heis0TrdRNZiYCvfbmIXzKeZQAhKDATJi8ib
tNPxU5nRm9rEZR30XfRaoDF75zq4qSJbWMdcpb+7fCEdZHBhCNTN6hTH+CcqIO8XxHpkIe0rxKMO
mBRpuOzdwxc9Q0r//qWXpfvpyHOWKYEQJ2qOJq95O8NjmsQeiqOLeD37GtxJSDOD5Y1pt1z3PZ8C
HvXL7AGuZRQ78vB0gpH3uxWV6zr8BmCYNxle29iMkYKk7/nMMTSCoy9GHPCdkfNMFtJC3FLYYwuo
PTNcjl4IN48KmTOLBNWZtzKsIJh8t3QXN1LVsqhpM4Gr4WwJqiLWH+GjHT0d6paMFYVM3in0bERX
EdHZsM6bfNg3kmrYCM/olXn3Jn76kL6WsVdQAy2cDR/VjTTzInrKh0fg+RpeemK8hzqzG099C4pw
Z/GHksvLShTeNddVvztYQJlD2qNSQsq/FL2JlTJBTZ90OOCS+qMWBH75ut2cotWajT6Vs59Fwv3c
SvIKFhcxPdVlfxRcY1f+vWPaYGMt9vpu6eWWHRJsC8WxAHvhUn+iTGKrc76PzC7mo+w3Iyu4zDTH
RUciGewkbzuqzxTl8tzo5nPYwpM5QRwtRts5DyV8Zr+6K49pkWt1aC1LjYpDj//lT86dV2Qr/U6Z
Q4IDxuWJS1MTXWvXvWih4ajrXCIR47t3VkBy6PDDkLKJp3YCxM3sgpREmpsS1zYbS4ur2CR4apfr
3iQndU6QJsMDrf9atSoRgHfuRffriptr35bZaxI/UAuggpM2wkzjSf3+2WOUzdBlMrfkFeVEZjvI
egl8Y1oaSy7IvsLui/B6zagdIft4sxN3XAa3H9qQEFURLNjO5uJd8KGHci1iOtHGoKypzuOqJM+z
l6cQxjracZVjjFGvOFYgJ43FWJ7y2NjglqxJbTJJ9NEKefRlAnOzzWHjJZ+uN2KQ3xE37lgEO23T
SMXAAF5cc8CNpkrDv3aeI+/u28CiPOjetP1cc/plH8amJidSt2EFgruhpCmPyUk1d8M31q8IuxQv
sN/qCWlGTTbJEcDzkTafYP3weRAkN3kcjue5HL6IaOE9tomdIUL3NKDiwE/UqLO/cKeD6+dgnV+X
ORxxTQaKo1juTCH/11rEZw6nnTo/w97t9+/GMswAfsZkR+rjF+iamXu4SSllB6cyt118mhgbeL3c
C78D2kg4XzeGR2CWQoS5d4fkEHHwgJemm1jUKai2/b8ca0PdOsv+h6neKw8hfQmBOll01RtPUxmt
dhLF5INoyYOe+A1Nt/b2CyvcJtdyGHXSVx1IFx/zTpxBV6BcvBFFGCJF63dAEh6RNEv5e/5kOaAw
sdN9M+BkhUbfr8h5eW8VxZ879Ov/lYWkFnzuwf5JmmQI/ZP5hLhsZkB/TSTXoIlPoisBKrR2Az0a
NdBBwlO1dzRc5qOwriQ6sHRjshl0XISFfR3DWif35byiRmj6JUBiihAfbXk0e5VHxi1pRGS8psOT
7fmbo6eGrzgL1eybhMcI17UXPIezU/la1Vi8ZU+XPhBGyo1URvCXZfASpna5ucwj8nVibd4Di5mw
37biLFzrdaap50bm9FiynvRblVL9ujKqCc1NYNqP+aVt/H+/rBMfJhrW/MnlpCpEG+4tCqfkfg3g
r8Z1PmfD05TzVc/+lExuRUFKWxkHMEJ1MNLzpc0NFglofL1Z9MBQDIho07ow0Fs88msTQy8hq73Z
sJk9/c8ENgOrmJikSluB3/78jnL95b+EKBaSzBqizbG1tEdkrlbWXH5hKVPhoHao1Sgu9k+/Mpas
n38TvH9XSnn6Yywpbw9N/quoNWk/8Vr1bunhvD/kiJKhVfKgZUH9rB9XqSy/ZmqPnIOCQ1itspIl
xp5UOZMyXYH++VietLq01G+RabsbjMkVz5cwAMVt+Uv9FiTxxwoifONLUIqf7ZIvVCvvsldlWS3h
e0inh+5v4goypOr/0PhVgPwiGoWX2SVw4q/lX2y6M2wrFIBGomQmnyWg9nUpY3NtisTeVwFmazVU
jIZD2UNyQ0N7Bej6GkxhgFtPStbTzocLuKVHlpRTIgzQXXrD32Zhhdi5Li+7a/3IV7os7jyiw/hB
LpT8oZ748tIuzvSHhUcR7+LsXHjiznd1Rq76zKVZvFlQILBRNMoG+nYMNglI/6gAU3GYHgUKa79T
Wbzw9OBMpi7l5nI/HsoOactnSst1IorjIjKr49iqov6frGtJHPcpvFGhHMYSuUHkZCqFlIj0Q4zB
iHu+xJNP5aHmNUWd7Ze7T2TkE+e3Us0rtCnGAdqa0OKw7wdYDepTB2J5nTQbKUQ6x/YKqJk6C3N8
JwhxLtcA6miB2+y6o2rxMsf3jMrys9ZWD1/FjsZ4G56/vfyzDiUEdst38UMsnhpkqZ/3tIiUUJ9s
bZNUSnBv02sU2A4NbS2t99VbHYyg8z5ax7py43EjU65oAfm3fg6Uzi6Xt5K3gMizGjQ/IhbP5ZA6
lbjj7MWfz0PxNN28Sdr8y56YlFoK8oxGmpH+Z92rKIQ8v9Heb+zACQZHCgqqv+yfJ2Dq/rm1t3Nd
EodHJuhfZuNjYcF8KbIH5OIH8SroPgiaZYOedkVuLpJpFPV7aUVyb44J4PhYln2yevevkawkegVV
jblVwJuf7Zswp10V9d/YdrsbtQFoJ7kWnc8Dl7tZUK3SzFpoe5//8Qu5YUfg6IaOnap488QCdNqE
dE2XvoddcZoblNDS9QM2FCty2wsZj0UL0dncZ2tmzIosaK7QXQo+EhNf76J6YVvQ48dA3bdLKMNa
v8AZA1mTwhoNpaolwNUz99x/PHkPUcwMxHTIiSgeghSrQYaYk4/R41pAjKhYs5glqQrYpumFUPjL
LyIEXaOPZc77lK5Y9z8mBmLJQ0vULsoM76r6L8qeiFISzalsf0eXvJEEHCJkJ2ggStpmXd8lUdWN
YiCmaI8DkEL74qgx7TiKFHYnVnYd+CmJp9T40BW8dxKVu09b8Guy/vVW7iicYZ8MyUTQCFE8Jiwc
GOhBcq0wSKgrasF3WJnhLZSLBq9FVhTtKZ3r8jvuZZ8/NkNH3rwM4GUAex12na6BTOnGgT/EF49Y
IYOZhBE3QddFzGnauahwadKn7KrrxAtOs34QQ9CtmTnFrUK1IfhQSJJnaAb+Szia+uWvPvfcDtf/
78EJTlbAaIV1Uw63TfJG9xB5vC+Zb3nvy35i2rSWidIxWaZGnuh5LQe4/HukFCpxA8SHzwSd3MUG
EmA54bKXQRTVreZkCy/I6E5xKaxLrbqfDEC3GdjKWD8k5LHeww71e39j8uyba/fkj5po4mAzS6p/
H5B4JYe2OL0HUBIJ7gDKmQ6lmpJ8SOd++DxYl6kqxg9XQjJJ68tQwAQPRNg81zzn3eg4DZGEJIjG
fIXc/QRrH+DD310fepkGEGHLiBOX3egBO1asJquvI+2sfnmhOs7iaGAAdeRrSARPhmafHse6OoMl
7kPfqQKVEqnOqzAFlz8Iu8qEoIiHkNDN1oYZkizHwODRH8xFOUKmK73ekmwFnL/JmkeOMPXXVcLE
PBxGrSs6ZDwGRgDxXQ5UYEH6ZbwP7VyHK/IeupbtvcG/ugS/tnlykwKv3iMM6cztu6H/MW3mP/T4
OgH3h3OLbSJgXNuKdTn3z3YN5kRiLaN7SNMtDy68oak1+7+1A6PMrM9otgFkPudnqnKJaU6maEO6
FpZxxBDBwxXCaqQUP+H4jfuyYEz87oExkcfXYJ1TJKiFJN2rzZFBfg1EDO5oF0yF4sTRJhl6Ivlv
s+YEx33YUypyYQX49JPKq0U8UglVd4Gla3QoQLagB3zOdJ+sNE27Ywz5T1o8Bt/2j2nY1LW3LWn8
mf1axohJNdt/JhBqC6e7U5XhZBjCy7JFoaW1QhgRno1mrUWufqNlPi2p06wAZkdB0Uu8ElPeAcDr
CE4jsBAHV0c72jB9cow+fXYzPEOY1YxCTvMxR3nd1/43x+CcBPHSLP9KFc2S7s/ZkgAITF0YccF+
/D3ChkPPmkskCgFQqUM0rGhmYnXH3ekj3pl+XkTMu+AKKzs6P8cZz+sxOkZB7W601q9/q0SE+mT+
SE9Yg91vjz4iHXWUMn3rFxhRHItfFHzjO+ZzBEC6iKEkG6YKdVCSEGP2uGQAoGLytWCbWbOL5yG6
uz7SbT0s+hDLVg/r0RQbATeVUoxY3V8hlDcDaSMP6oZu0iwsfk6Rumk3GWD7IBdCJYR7G3YhvmOP
msfy0IH5bk/U6fxAu/e8qF+qzIUy8b1eWyY2Ce93lzhc5A+VyGGM/GraOB1zjk/lzxhyiAR3UbN7
WCQ90GUk76LFihR77v0csT87C5+Mf0tMwGMo3NKLQfyis3RG7ZfFIf8c+QsRWMuucdaWLRPMrRgk
d5jvn4qIuz2vLfem5e7NC3jJv8PKireks4ojLR98SubAUw9c2m8RtFPTJ52EPPwJxuK1x7t51YWJ
PNpmfqRKET1GjKYH5f/i3HYbu0a+Ukr+aVIvgUTFVbkpS7yEtv8Tv+LEGKWKhE4jRPP6zBwXxIt4
eCd5BQGvmUWFjq+zW603ryJ+l2gzeo9ypzaCwmo6I8duzJXZuYbf/+AwTZWFIoWr7cjas8E+0OAw
7Ol+5TgQAQBoX6cz5Vsl+GdUwo7gU6OqSP8aj6+zGRRkyTFg9G7cjujSQbfpGBOT6i5fsFS9ewah
TD00uJ//VW9o8N1eB75D+4KGV77daRmyXpGZIIZS/ETfNbZcarrz02lJP/P3m+0lmjoQsZNgcrp6
qWx23vc5T8H+eNgdLXyHqCyUoP6ppVHKC/X3cxj9+nMH6Y0pjBMZ1SpgyfZLUX44jgyIVNLv8CTy
Nrg3Q2K4t12f3uhJLy+V42bjsBxiVzuCoMPfMz0cbZuDbHfND5tuUJDf+DJtDeWJ7Fw5dHOga4ls
5iYmWbugzzDvvcz36Wv7FPsGq0tkOyMNpb9RX9VBvYu6vsvxWqqEncLPyWtVDQ37erI7tQLIVf4C
AEe154TLFXIuSgQO/uPLpzm8uNmNDCqrq6mACD7+o2Vd9DWx3F1cQ0vfIN6AepSmZjWLbFw6/BlC
adDpTD9dwQh2xm+2bojxMQ9Wq7udNezbJ3R9SPGoH7Icbf8q9LpWZ1G24kvso/ZdWFPQUvC8J5Uz
1km9czfZkgBh4ySEkxlJK0mW82TT7EKOqQsJ4AP/iTMoqHvvr2/PFWKUgDki0sj/E6jeuSJTNrDo
8Ob6N4e21ykdi2TEDgOg5nnvC6MeNXlfYWLD2qgDxDq6uiKq7fMRQ90aG/iHFS+PpKsXAiLugAtP
E9SOx+Lnbac5Diwp1H1UPG+FIY5J6TZmjnE4+z07GJviq7zfsgiMq3Fd2eDO1QO3HJG3DWizlegY
vpQ4P/wfpEh2FkfKFLRidlL9tdrHJg8pcp5a9m/r8FNN0Dn1PyYf3/GRBwVlNxOV/EowmDa8Yd1Y
UqKEItr0Vk4th5gCkC6bVPm8WaADVOsFc8hrwMEFAxParkbZoIADDJ3adO2DiJFhJm2INhu2gqzJ
PfeiHGS6rkZ1O14R6Kr7z/OhpZP2fYGqG5ZZlzSECBqxzR5Tirj9aXX24v1jOMRc/zaJhgDoCAX/
lFdZYL3c6WNpcQ0gF3PcPaM7V/A6nSix4HsR/Mqb9+xqgyH+MrMvw07/z8bDWoWMf72fMraymh6J
RCT1ycvGxstmnwJjk4yfisRd0jtmpGPa8hLYiuCS+QdSWm3R659wYC39Z9o+cEc6zYI0k9L4z8FM
biFKTmecid1sBkJPBD/o9Je0TNsgCBSSP30eiKbxrCwrg+fHXA/GTq1AQv6LBflhTsrj+EWn2tJL
PV7jCPRzZ2RzhZ56202KD+uD5WjGc0rBPj1ISNWhOScxEenH4389Wkz7+rFd5OzCZM5k8BG21Y/T
1r4J5MPfQCloaRY2i+P3h1uoECMPreUdHd+wGcidn4WzDUcfipwyaNvVGFPKEknlwG41sCebwHBO
SEURC9BvdoiyAjWsYF8+FMp2bam1+CoOdcrOj+UiFy7SzoBo6BNcD8ygnbOO18ooXkRF0WRNdW1O
5BDQ1rUXeBUuDjU3cxI4oDd51iFYPxUiYCL3cL/tI1UYWo7K/cUiG8UwslB+D1X6wx6MCSXioZwD
6nLsVdlHZE13qlztXnkhb3TjMGjRkeux/YvJaqEYXanTLxxssNgEjFQ0eyq6sdX6fHUNoMq7koem
X94s8s5RtZ+anc8OxKD+kItBDFthLA5kFCWemzErD1nFEtYhk5mgtw/ai2j8NIyPYa7CgjGX0Yze
POZt9k8YZe9QeJ0o0pP5kpkA+Rvy6psiuL/QWZ1fKdXdtDRFB2irmADJ9GRHsvdJbyW2OHbDP071
iO7kjuwic3JCmYGTHl7kxMaC2Ds0U/N4GmQIXIw1qFpZ2f7M6BARyZb1wuAViLTY+qIy34njvxr6
oZh6DcSnv515PbuskmIV9/R0vuDeh/yIFV6BuYRLoJawHFbL1qWUZZ6Vkf9Nr8e+72UgdX19X45t
05voa6biNfXboKJ2DMYBfsq0t8TOBMzF6WGcUBEXMpNtR8avVdN4xDCZpWsvy8i8tDdWhleUr92R
yZxPShpWr54liFD5DxvOYb1i7TGlSvcF/NpqmR0k/qT7r69BKou+dh75LdaokZzoVGZpmxR7QxK+
DUoCUB1lltwAKrRgzI0QPwCldi+ZTo52ZRny237ay5OW8OZfC8+0h1TijXgOSEz4BPzg7ggCZyAv
0UTKOjnF6QBBFIJGm3AVwfeYp+SdyfRYxIlNzZGYBmnjAstitcJXCFMrGc6e4msBbRgrhnUPCXq3
Ril1ZwXitd04qpX5XBDGoMLfZ7pI4waPlz9C+glbFryOGuZnp/hPbwgMtKdKJFGk7Ebd7Evi5Q6R
XDT8AJ/eW6hCPINFfqaRYw2z7ilPy/BrQnTyhBPj4AEujuJk+M8Xdd0jfykigVoVWEv6kTWCsI6j
SldRJMaHj8ps/TyumDk1/SyEYoBBPyb9fxyqngX1DMTiclECxnl2boKWmOQzFvyhc5mfmMFHxR81
KzxlRmMfka7ERZZwfU+Wr5Osc02iZaF2uCWSjhBEszSxe0rJBR0uN+EzaLL+zo1FShoIMvXM9Jbq
evwt3V+leNz99qmIsUI9dJY2JJWC8JWWqtza2xfbkc5x6qn+PVVzK5Jtzz8H5M7NYKWByOcX1igi
BAVpzlGjlG7aosInKvrvM0CD4edV44jCViZxJOewE4/Chbf+ouPl0olcoihMmk/OGi14/XwfsJLo
Xv84ekqcr7W99DJl5jZJlqTFbiPzRJBVQsCamsl82ttZpjKC49vaHsLr9kS5bDbBFW0qAMDiAicH
lwHqvc9wJiRPrsJjVp+Ai9KXPX36Vzii0CiyL8mUNXsCYraXxEzPdT1pQBYISFHdrNuxb800Hzj0
9I6jRcKSL3x19286iwsMRfGS79Atg9xEFv4CcG9rVZHtq2aE+AUXMCrldC+8DePl6LdTrjK8eV+3
cvjOLrkbaRhGfX9lJ0Jkd2lDy5/CzQ+QNAEokD2u3vPNwZGA/fcMA2NgDXsrakznLYk+y6kg6uL+
rxCmzZtwO/9PPFZJ6jKDztuYswmmAY/ZS5BXPRpQGjsmSUcSxEpbV+LFKaN6Mm1Oglwv5MdP/rwD
1ChU0bieue1v7qGRGqE5VzIpRiES4cx+YsBbVsUQodT9UhWL3NegJ9izA/tmSpIXem4+NsDX6biW
5ND7a6ZtT/lV+z8BhlVsfQDtq2Tfkrh1oF9ZJx+pavSfa6sXrdhrtS4xYXLzfnnDG3R0/H2TyzpG
1hWwTcHftMrp9gi2s4cTxaBu0dR64ncCWzBs+QN0LCxdETJ0oYcTTK5v+cG9m7vhYpU9wiOdSTmm
Kh7KYZvXWEtgQEOAAUu+HpDlthXZJhBoqjeky1lmMWbHpHRiMrEgCSeIfAzgXrmDgZomT9xXJm/X
lnpfBYbNq7o9RuBuVfh/lGaCQYiqJN1i4U4W7oxwYgEVH6pFXADAi8CwzG20FinX9yFTpPoG0RfI
dlgZi8whZkcsVPJ7aGTuJSuiopIkflu4N+7kRuRZFx0Q+2Uu6oanIfvbAJ4dMXHW0YCbRCR396rz
LXxfgV/wKAH81NT5WXc7QB2vygnPBybeh2uETlOhTEm1qAPG8VtNM4TiJW9yZ3EiItXfNLfudPL9
gVtyr3RAueR9c8xOUxK6rPkz1xtdCC7uhSPtRo1GhP+PGzBy/cvcIDhXFs02XbWjhsXgdPlfmrsi
QeEZqT1gRshJmvpSYPpUioC+JeMEwHwBjpuCTY/UP+hU3Q9ZP5ZuxdNuLz3w1f1+J+gGZ0ZRQ2Mw
L99UmFcEWbXz/RMMWJ8/DGyXZwESE9K9WkerO6dRO3qUfuCY/YhYSmjWbMg6ri49wl+P5CP0OnSu
K9TApmUl4/DN3RjNJqYSPT4ghL6viOTzLJbHu1r2zbNOa8ZdQuvP99sUcMkICOfLAWswEw5y8zGi
12ue+yHVpl56hxsr7wX5nufQcBQZ2XRGgN5CPDcMD5JpaULLkTa9LMcPwH442TB8SxzJacN2Qs99
BTzqV1bc4NhrYe2TgJasMPFNnksx23oQa7v4H31Orq1iCu46Zlz1YmVPzs8qhkwTAy5LRFLN/gYt
8Bf6a/ArsU4FGhvufkUq8pUFBHa4icA6YsGUpkhQCGa6sbIehu/3y5QOabd9sz/ahTqLzk1I0itn
LK2nH9j/W+eKoBDQ8Rdmva7pJjIPeJLNkSl69sQoa2C593wthaJybV181VUBYzpoXZB6ELBQJv95
Do2jG4G0nAASlBMqQTnoxGNQ144zydJBCyGUYVol3cU5ZFo/a88tYXv/DgFlVyReyfjcL3KBzEhL
DMPptKwGPlFkuMDepz8veU3yGiPKnM/bVsLFfZmAu4Im5ADEKCZO2fKkcGfikQt8EwKYk2kZtkeG
bAA2uyPejfbQ9WOua6IDsc5VI/z5l0Cyscn5qmnAHexDOnKURgVO1w80IY8PhZHAX84MZBxoIAei
t/uBguj8UUedoOOVkIkQloozlUwGdWTsEP5PlS7EZMDMEZAZS8ElkyuScKyUdxZp6Y5pb0fmZ2Pk
6bdWgq2SnaXcZLuasqE5M/r8DoyKTIttY2k1n0T2u0AGYlmnM3V4vCu4kkXdS2h/PaI4GXwOY84B
eMeOOW307azsiq0TdUl3opW9uvZgMSsYRPYsAuwctHLI1mC7OkiP8eAZUa8F7B4VNQI8kiyc6TT9
iKDWX/JUnTfhixhXPsR3iXXV9XbPnTtUWK918criTSn7A2GFnYdp7OsgQDdJZUTmmdw9gKTYkUft
geZYJ4zEcPAH4If8abWPcYmuOTV90qXq0o5NuasSuuNsMOHKF6mqeo1ifDC8oNZ6xtZ+VEG7EZuG
DN0ZIswoGo7YNpX/bO0sdrWVSsForatWq3Yu/qzFDkvnFSbxRgj3XeFMQeSxiF/8wsmO3gw2RPil
TBAEhklQtGT7BYhVd4iXEdXR9FJ3nhGcUg0NbfZvqUswGzuFeKx27YOSbJh7HAi/vO1P4L2GjGLw
kvAwJoURPIz3AxMQgOayV2MwjlWnU0fWMQEHtzoe5UZjhRytBwoP0oneXYpsYsMdU2UmZeIEouK3
T2cxfo7FaO2oSu6IhZoXgRdbmgrs/byC2Nw9KseviNTUOuAAcXtpj5bc7H3auqZcGKRj9EPpvsFg
KacItjEuStIRLebHnd+JSI2X9+dibCtIcvjpf9yeXKY2VqvG5BvkobG+VTfQx7UsUT2d7oWr6RHr
VHxdTqd06TBYa6c0iy59M89rF+WHBvvjCoqiRbp9baIzn8SBI6rmVO11z4r5rRgsN7z4je4zuUBK
DkGf5VFRTUYzU+ZsKyjlbIrNAAUQDf7cl3HrExJKOpsTL8oAIM+1qH4iGWlb5zX9sZrrowF/NOhE
kidohd++RX81Z+U8+9+t3pxO4kXSX80FZ6KDs1HBapT98yujWns04bdBHPO6h7mRY8YTT/bO+dtN
bBytJCSs9JSFABXSElvJQgOZQbCYLqfaprFmGJFbAbTvgfvvaK1eQE33kml9C7jyDiUsfjvhoOsa
bb8PUC0XDD4fjsCNuS+9H2hC6JN8wR2kGkodWilS/LxW+C1g+FL3Q1fX+D2X0nk4ERPIHiGGPZ09
/cNvUPTfUOKPSt4jdIROq3gRg/FFN7CIWBuVGqgmm7Akg712GUisgEOmusk+iJsO11Dn1Gw+7RNi
txB121chv2e9cCJvZz+avsisZOAM+R/8/EPIGIbOhIIlrpClZVRFnbUExW2rT/Gt+A/WrzXI36Dm
x+aCPD4g+FE3apZDs4AYltVZB9knj6/9DGducH+YiF+qAOg4Uh4DYrbCsC0WC1JHU+ftkKRs+XjR
KGGMeZX8sl0UNFkMJ4Zm7hfwr9gculBFHvSl66gOM6vfhTWq2T4ZoQq1ddZDXzO0FIEMUqoRnh3g
+HsD03cB91yQ+h/Y4Tfl1yFd8pN8n8pYlPs6OMLQ7/jRcSs8N4JYD3Kv+0Q6Xo5xvcP+6e6HG9W3
m+oXVQ1oYYfShIAspe6trOPA7voafUvaLoUsSYZoBKAYeQrkYIkw5x8JxM/nW74GvLELEa49h/qC
j+V6Iw3WeQFV3AQ/ui2zsQX9G0cccwAnHDJjxq8+0KLcrnLZowY1NhGSA7Fc12jIT/nD7BDX75Vo
MWoC6Q/Mcojjz1ADgDG1VOlBxHIr2AZ+LIUJIxPHdHE0T19n4Iou1nmNt5HGQ8Ui9LLbjbUwTx/s
PyH2/0D3tPrclCUCx/1mixm/nd32PaqfyYi+VmluJvv6bOQC36yjVh+S3CXPjZHZY6ckQCCNjsxq
W4sL02PBC5IOoXIcai7fHtjfAvbZgsET2cq63lDHKY4ZPNRFD7hgkz4oSj+Yx+VqFw9kzTSdmpSp
9OP+VC7hgvnbEIUuZ5cQnU6LZ+8rxkX4E1KC69TAitUH16sWwki/RfyP9kBYj4RkTjeygQD23QVO
SnkCBF3o35rhD0Ixqk2jFgmRo/e2T1WRB4bb5tSoJxE18foYQ6vMBSnGf036bYAs/MjEhOaahXSb
o/s83z5nKyN02OKTf/8Vm16gcWQy5BPjgPaysytnUEEILvusUQK+5xTpb54g1ecl/PMxSrX69Svu
OMH6le7x2JkcDB0TN0UhUY+aC/Y8UNjX/6/6UKQIVgsWdtSdeu4yEeTlNAmnOg8GYWfrvTxoIHaG
tiDt9Rt8uz1un3uPmOei9bl+GryzBnXdX4sbO3J3lRoWstIBCtVzG1/S6qeqb+86bFaCINgHPmyE
cI2L2fO7DK3qnivxPb+VQcEZbMedkdSqQ+jOQs6fn6vWR0R8yMGx10jF/26CbtTPWUb3ChYDasP6
KQg71J0m+BV0g9qUgQ+35JY2MwYNOJPDFmPXF+mzUXytIl+srOhvVS9nelpoC85vWQS0IhsPpoCV
wtO38x2IY2/kBib5nx9U/tBsXL9Ri8WpRafOzYexC/P3Ma935ZXLsNADh9UaxcGj+w4bpBBPHAps
tpDnPen7IaMoIjvhLDVWvLJn4dQj2YAkXz4n/13JvYH6xnkKBNzu6Xw8PLprqWyXwU2gozoQfHfj
jfKP+Fufi02YitRYlUIwB8WeJIxS0vZSljxa/vVBwde1DdwLuJOeKJqJGo49cAsVSRQ9u/DN7H8f
JEr5+7MYPnqyEoGmYGeYgOzedisFW3+Qks1o5UL/TZuw6ZvfN2Noe8sk5AtieVmTnGA0eZYleajU
+YrcDJqDReZSwqEPhlBJFSYYJRoF3YcHxTBYqDrApiW4+LVBejjEEz+8NToSglUvsZZnZPk9woYX
lHz3GtmZC9RF7pijLwZYgu/RIsufcK0GRfsp4ndvMMTvkRpVfegksLjt/LS1HceXyASUAdPHHHEL
F14SecU67tvJmihzON4AtKlQN+gbqo8iOyoiR6Gzf3/ki+rLRaIoLiemqCSaP/G0o7qOJqXpF6GG
W9+rPY7jZObCdE9R7AoaZB42a9Jj13m8A9tcYJ/uuretUYaBPfLtIxly3E9elqk0UsA9h5k+MtLD
LX9wUumwwF2kq/Vn0yxgwcAGHSH+J2cZBanBCYLeb5HjeHSpx2XyFz74leC5XP8Z02lWRATWaU7a
j6CcefHDrwR7bR0wXZmhYmIT4mEe1H7Cr3GQ120lfdfW3brDPeVIJmKC+RZLyoh24FWY1/+GMoAM
aRMoX1ELp5MwbGoLqERhjCcFLKAlq9ErWA3j5x5QtfV0SaQD08qy+J5YtcSMGa2Cz73fQc+gCVwR
h9B1fbNOJS4+l2/6ZgDKg3BwD1h188fQO3E7tWU/9PzkHEaNU64fbv1hTiqeUx5ckx+1Iw1dCA9p
NTeSiBMdsbcMupzqyc/Vob8ilRORxc4YnSwJctLKD++Eb3Vh6CZt6FrAyHa0P4JIrQ50LynkLO4+
B7y+fuGLJ1xCq0lEUOabmVCnzmbPNv0UdCRY2B2nJODGGK/xETB0d/gnElAIzdHSbnRwAwQAPkBZ
6k+rk4qOyOnKBanZ2bDZc1T98/r5+m2KhrtUdl2ZV5KXvot/n1JD6NnO54mwnUKZ64210bP5ZPse
Il7R4i2XqHBGmFu/3wC9gSYTeJE3uou+sr94iueQ+XP3Ba9A0EHKYEx5CcLnnINtRniq/FGuoxW8
aTZOiRzUTmSq7GqubZax2EFL0t72lgQqEdvlPSDkXvFOU+NLM1wBUKtihJTMczP6p1t2A5/rXf+k
w2fjqrK+F9/YLMThyHvuffSNu9lFO1Htr14h8lIEN/n8eKc5D5Tm2x1Ju7bdbFmARXMgxGXW6SzX
9Iyx2DXjdw7YigJR+JTY74BFkt1dzir48JswXEjLrI82LcIRNtL5d127/aW+sRMt+YRnp8n7glnA
gk4HgkIG69v++IY9WojtRHKRdGQgBV9rHyM69/BIlMR8wQh9QU9Xb3AXXEf5K3hCP2Z5fbCxxb4w
b6xlxaeM53s4IZZwM+YkH6sjujARJrQGCd/XC5qxyid0S84uD3Iq+THr5VN8EMDd89ShkjUKL5tW
M07RBv/iY8mIRNvHWev8pqYJodlJVpuHSKnGfLePccj0AKohbqNfbguAEZK0067/ly9Vi0goxCLF
MYDE2Kl8rjSYqsbwXGiiDFY7T4ZEfsJiSrWbtoEQREjxZPoTJaG2Ml4zUj0YYT+wAul2h679t+fX
AsPcVFfYY8vv3bFGHxoNp4xO363VZ/yduzCQvpt2PN3BsVewyIHiy3h3+qScslTCUpCQLZMkdfw8
V1aWT1OhuXTqCWJqOa4CL+QP6wjFgouRT8km7hCA0ESjWfxJTv1NQSnDoTmmdDKqYZOSGDiaYWtX
7wHtl5E87hzQKk4stRkm9AmBEFI8kgN8NiMRwGOvMUcEsHLkW8plX2aYgrBTreNrz6Slq48bMtDe
ub+EnnZIPntILHufT2625FCzSxr02T8JgIfZ4aSaR++p2qVyFpom6gk9UUxXJbv5hVsY63iGzX94
zPE0cMiD+zzkubxuFQjU+STXm6SwIC5+4qXB/O5s3WEC8zLiUqbTK+AdI+83WQB0/2YizX3rGLmY
Xodsno5x/d+wuxNNey2lAj4l3Ti/du2hGKVP5GsblaaS/k7t9dxEyA3m7RA69HH+bYCZECVSbEpX
paMD2z1jT3/Ja49baOQ35eB9lNrDd9i6CirypX3WbsPBO91cOV9xxttOUQTEFMt0vslDODrrgO/i
rvegPUcN7GtZaGBhlN0h9QM2QugwK+x5EXyVMKq6rvCdw1TtvsUW8+p5D2y5r23jIg5txyBmtOEh
cW2/tIss4d4NQ/4hYvxjLh9r7KGfQML/DpEcY6VgHOuo5szGxqYM9G9jax/VrsANbaGo+014VFeF
lvGaGaliPK1fxaC9/FTB1ECiUyUFu/tybQtFag1NjNe1MqPguNDxpLQlSls6w2qCBDJAAwgwlnA5
8iSY3RIk1vS+B5X2Sp4g2r65fe1utqVePGfutX8tCHOekXf40nqwOX9cqrW/00tdwZTqosKnsOxq
QS4+XqagScwNUgiXYXZ9+Rmk67laHe3TumZL8z+4CB2d7XW1xL2OQY54v79vSY62YgaqQ5n1AO0Z
NXoDdRrf0W1hObp5zBYXXP4QbGTBebaFgDyn+EbDGZLNgC9xWXJ/dTrYncDmfhOjRb+EeftmP1oJ
9GivYmK4+0O3bbvE8SZYnx8HAFqovT6/J7NdkGwnxa7CeZGErnD3dHTcT3VsPyCn+HlWvTFYx5wF
ugpWsxC4O++rW7qtMey8XrfUA5wjR16SZOQiMscDaI0bfxI6terJr52w8um3mXDFSW0JJ9KJ198A
1fHd7emKh4sxXq14eosVFMg1f30zSqffIFunYvmQle1fWt2wcVBt8xQAPCxP19lMIEjf3Jh/MFpN
P6bq4z02cW1ikagP5cfrHjlwMq1oXpH2vlG7Yp+T9eqdH08cAb8/t5QxvjjswQId1o0nrB8Xb0ID
xP5NATNI/GNzjwpaEQSz9zrn9Q1w0NrcwzU7Udc61b4CQx4UyxWY40R6aAXvod/vnjPWFUr6ZIhL
qTSbxMqw5kA3Au8iy+zC+J2wE6D7fwNQLhiVYJ0wg6tprR8ue8VYy2GVTYf66n/DocYq289ccpTP
dwogtIRLWr44fRn0UeG/eFVJC7kA1of3hfFmcP59bpD5d/0RJOwHJjwW/w8UvHM3LhnZeZCvw2qw
I1gc0KILXkQrjmXkzhyuPXScxNT2Y1je/LH6q2pOsOLGkpgJf3+AageKHMbb4eeJtTmjol1FEL5X
4Sjo48rFhdHEcxCSDIsW+tKleRzKFTHZW6+Q/VBWkzRgtXTnt0Q+0lrJpEF5L37KRqSiFDResPLb
KwxKbsTe5tYVTXV/EM4Tj9BIx7PgXmzNnXQq+cvCNqdlGnS9LupW4rW4A9vIYUebNx4mBNxxDRBM
W7PkKk548s8yvRvLX5vSb5GwGGBj58qMUBtCC+BxpH6FChwP7ZZJmumNH7mBWELTIfy3Z8OMJ25A
s9tl/Gvj6fBjrFU23ZGkgq2RJFVQGR2ZNZn7jfNO8awVPd2SB44iAUxLVQIDBZFlLzufFdMu5xzX
PwP3ADVWJcpbEGejQ9EZjpZAa7IflbCXg72QD1Xut1hB/8K8/LScBmXexVIzje1uKBZ3Xi52Y1pe
IHqGTN5pYh9NWJLVABhKH1TDIhy5lNaEjg8ubxkKnqdWmb1APObXIuL0ZQdY8cTfoBXaszh9nCVs
TKT20YfQgI9WJ8RLbqtsJFQrNsNwkKyO93qpYevizei4K9auwx9rzjTVmLTzm4pF4iZ0lk92aSfy
6I+yiYoKhk/ZykhstiAb8gfZI5Shw8cRja+uh7V7jgmIZGNAPoZM2htyDmGgUkOrj9SL0/UitnSk
9XpQPJzdyU1cjhi7LV9BkUJsS7zqFK0ZFH1DtI33GnvOIFPKrWO27lmuOWKZxdmpzzVPMLC+MyUo
Q1kerTINNNDI6y2CbvlwyTuyLPjdkhp0Jbak9eqdjcrM4V5iRf0gybh7MzUGTgQm7ChORRKAr+CQ
AIWjNLz4anj7s4zWjfaFrIVVe6+LRF8CArPutShESbhC++sf8Ksi8+G6/8ECWadakEXwCVulKhSm
G1leOKdAmL3VLaUJH3FwuDVf7CBxN5tSXQaDviF/cDkaQo0LGenjutz6Ij5Ibz84wi42pDtfPnHG
kkmQPzT2moe1YYpcE1QsVQU8WR2xf9z3bhbSQCxp+yq9B82ZNPAcP6901WRvXuagz6hkHh3lFy9P
h2477d+lFnJcBL85DqJ6chQaiEpBrjY5Cs1NdaLAUgQ+bhmsuKXfnXAm3ikBeya9HPq8rwJ1Bsyy
NNKMYK1OVqe3iGTV64h553blDtk5o0tTeFlDHgVR3kdEKlAGK7li0ewXaFve+nZBNXuufDlS8d1O
58qnSsPf8RA8ocgPW4M+1jaDZbrO3zCfEcIOTKyMIBuqTYxs47GOfc8qVdtszfIuQVo44YeX3KaG
5kFLOybbkQ4DqOzOgFicNUQLX9GmhoZMv+PTyfFpDD+So+9faxdFDx25t2nyngxKLYP6mbggyW4k
Wl8xh4n4c16Mv733HvEoqpgu+iGqEbe32IbFUy3jtjKIHjElQMA5ufZ0ScdXGh9n50Sy/lldp8qp
sATXDYplRlchjALin19l8bny4VSK0hbuea6wz8v258FCpnc/UmG6CSlR0DKebzIDn864gXrZvJlm
Yi1oj5ooi7YHmAWMYcuZrsLZi3m7jZYASM+3nUJjOcjS0wt+NDCw8Hu8OjP/en7h82tShTSlpUe9
R1M5kEE4eruv8N2rxOuaLr235J4BvWgezUFpxvujIiacHqfyQJjN2cN4x1sl5nFnM1FokF6ICc5k
r/18qbFofB8qSVTDlHqJ4Fe9fd8Zc/DRb9NHy1CiAehzscZUmYLmbUMgvjkj5G/XoW6jdsp601G8
icUQhY/1BE6wTxfAN/gyXnb6ZSky/PL+HdkZmLOiZCzPubr2S+zLPAuGsT+Am/srU0vI6ShHCe7I
PoH8z6a9xPHeZhRSOv/pHJR2l8U1cW04zKU441/ljtzRjdUIeuEQYY+fQGOJUHswcPX+1vX9e85y
hLo4/PNDvxYvp80LiDr/7Z9u1OrimKLesp2I5sU7tLDCDK9IojuOZTG8hO7Xq1yc3LzIrywMWuT2
0XR1tQ/ymIGeyyEzFCIU8JU+QVotmRq69UiTCzFl0s/W8V+/nn8h3WpRKjqbmSbm6qz75FsD+IME
vmdgmJK56zlv0wwKna36WemzziHBTFkm2g61OaV6wqjilavvL2eyWC/ilGgIxfhlsRN86Kel1sUc
OSKEdVss5yNhWatcsIY9Ve4eAyyooJ41xXAFrL/mHlPfF6k1pbY+QnHUwUa+Fy3BLmMj0UvZdZNJ
7rcBwJ6p5qB5/88UrM//0uZr7pJ7q0Sbc/hqh/RUIMaxwldRxt5cIItL2EE9rQbQruxlQBEtpDbx
AvYZeiq/+Wx3C/rVdJ4sY04vAU0C79MUnlbi95AUaswkadEqlHr7TbVkz0YstEKiRZ13Fy5uI7DD
/VvpPWQ/V6hF91Xx9Ehacz1FqVMfOW/f72nmLZqDX5yV8k31rFjVrbUA/2XulZSUhsR+9KGXE5c6
pIOEvdPnPhNoFDxhdxt5qajGELeAysYANQ3SCYKe61kJFsYDOiPIa2Q8BWeOFLXDSbHa8JS/DENV
lPufqZxFKdHQC6TmdbnQL6gjxiMvaliT6hFdkMv3vbOKYhEVGhCC3ngatjGfqoa/BGpCg5Uu+mAC
j18ibp+qgiBkRANAV0m2rtp/Xy/xLYDeELSdyNXfMN06MggT6JWMxWIarJDuNypgwTKaafaEFHVF
bABqs8eq0ok8CWVk1GvUoa7N3vsF8UNlY6dlDNPmVuktAGDuh4qZlYWz3k48tRo5jRPVZOCstrVj
7ncdb2l3i5Yhr3JuNs2t3qnn3aFWwcju0DfCsfkisHob2vtTGMXgGQgYZ8uWffq6Y/w5q7qIeJyh
RAnDAG6wfp8HzshkjKeHqjKQVggz5GYxUmF7owVTBCwOdNQcPDAL5GIbOIQlbCVBQrEOwL1ubJpX
rHKXgX+32N/w0gKdzbdbaF86cr4WCBLovYsowEKNkd+OVkPIuR0kU/pBvWumbXelBv4AlrQKmS6S
JQLCnEAZD5qTfdNrzwJejVTy+q9xSPUWG28lFooupySIgIw5DyhmcUCte2wyWrMtNP2n7we9T4NU
wBVj9D+0pqwtc44uMexrRiJi9mSi8bDVxKx45lLPDdBT0T++jntwShUH9TKKzr5WFKCIG4NjbIvM
YD3c1AYNJEiu+KzTuLExbiCtcQYwGmkO/UTRtf90T5ndbCg+EPr8xp9eemi2sGqAzH01PW/c/oaC
lX+FKNmfyiJeCUyxkxp2cJii3mqjXN6qOBCxAfOk1JEPqSYJ5dODTBh9Pzrp8YR589YTdHd1MGQJ
N+d8tdMJREBuQr1PaPQbMNzezvx0Oy3KnXEAl1gt3sDpd7LLoS5clm1iEfW+G+a6Wy8SUOmK4rbY
RBPNhwJF+x520QsFyySUD9VbdrCeiIDreaf4nhM+/6JZeNkuzEveZ8RrM84mRYkd2ij05hLqDDE2
OCeuATDf9bAGEzmoKQQyOj+rHjlpYzSBo6gnMzRUNMl92J4XbhI9CSNOUGc03ZdGTEx4j7VyrTKd
IR8t+WuLt22vhXW3eZbsHEFdufkyrlGmI2+eFhvAX+dpTqpVzW1Nbfqq0+cgsD3Ik06wPnPmz8L1
N1CS+bdAjHTumYAtv/2rioBcUvRiDRsbNd31UzpYqHqEXgIH4tzlsGxEWFzk6yFPKtPKUllDOKew
e7DjVxTrJ6ygqw5DblVQV3TYk1rwwQQuCtuxNF2fTht20nsDtxXwfSyr+gHfFqjIF1IME/DW3+UB
+Jg8UUrwlb5ErJJM10SsfXCidwMuh0WZEStIAzFsHZibIxepJmKcyOnPjVkUGRGqYBwZngnZxoOz
PisdYuQw0iQyYtupbwF3G2vIhLMz80ts2j+jjAjtw494w9RhhE83+K+W0HcaN0qYgB8QhE3z+blo
aPvAxcmQVCuakGrGZ7BnL00+n7T57fyJBtb2YOtC4KEEw6LqcRQLI98glzNdmp3ekgcRVr030cxW
1LBlPBAeutcIidcaeJYi2V93cdeHjRuxNeCOdqoZf0dvYuZJtXTixvEOfO3+0jZOO9lpV0bWV1VL
c/bNwU8vn4GAzI+nJh1bGkm3yARvSJBDNCF81VdjNsMAdPvBW8dEyyNeeOVdb4hBdT0/bznyV5uX
eyrAVwZVoE7JR4N2m/5zQmFk9j2kZlB5ySlzkbncx+p47sXKDkEy/WUlD4W6k3C11u/h/ynI+g5X
nonVNd76BSkPckEULDLgSt4nf7MCeDjkFVZ7GZx5Y0QkFKlzSRYYpkcK4XQhf4B2jBuCvwamIb6k
At6fELaWxTGn/cckJTQSWRV5AtLwmc4zhDaB0x53O42SGlIzkad3FCVtpuwji70g+anR1i4I1TVD
fe0l1Yz1VEleYER1qPXX3w9D5j8WxHlOYIXAV37uYN1KvWWWpHvQcYs1YhiCxi0nqHqr/btgBjNG
mtDD4wJQNla1Fy9WiYe6g9B5YUjSsem1gY/rNHO717jXEEFFJPNdgQImELuAeIcvs7/n05PPBWxz
Luq+NTRcDGbI7P/URz+Iwqc59KUgUS0yfrVmh0/VrPzVDkJhBd3eX40SVugT2Ob3fX5aZIN3X8dx
8jKTey3olLFkISHyn6gm/IV/pDNK0H9E2qb8Q+c+VoxSvhHk+KctK+NOUJfO2X5D+w17wdMMNLzs
uCqeDsqpLLQcSVQ//5LVEdf+RXHEh23tvDwdPAXoJUcE7oTGf/esIhA7YWa330ee0wL8u/rvSavl
NLrLXTBIn0uPDlsrl/GRuPngyNWvw3HKsCSE7rWj0r2Rd6qOrFFmRFjrsUVliz8Pb7BedEYLqD5o
OI79sKKRy/ViqKCzqnEY2V/dEN9CpnZeGTxGaBoyBjkfk2I0H4f1H8nSO2grMD73GWHu9ceRJ0OJ
otK362S4/A1izYRx2RsGvHusKUMIle7RL0Xmzaw0erh72cEqgqgpcomgXCbltxHKaUjfrpwXniPf
t3t0CTPf/d2O2XCmnD8SstHTxSd3moCGsdE3TtSolExVIA+DswDvVhKLGzPLczQJow+KSD6t/6MK
6VybBylOqOedl5oVHBTgdBTP/NU6lgR6Yi9+Hg19pdFQGbkU+En2NH5T8SsUKr6MAQ5r+mSqWIXi
gSEpLT0GDPsXAWPOSqwkEQIZA0byDr+sMkzO4JlWDY310NpjpfJbT0pm1VI36Z4HXMOOhmSaWrSd
kz3HIAKuVidUcDK9f7Ri0eV0AuiipY9vTFPjIMOdHie98/rhZnmjj6Gq5VSGmil+wkRxvF145MSk
4BDE6fww7ZE+Lgzy1aRhNQxlXmBBFIABlpUa0kGRiIrF8oi8YDETEv//jrXbsp8SF5hIGxo7rXS+
7+sVRrWTx8Duf0pqGtbGMD+qPCZdoG7y3ypwv7zwZrkZah/XOBK9sHk8bfrQ+G/7w1rBkbWZRAmn
y4oncz6RJKFEtIys/UYyuFDOdTxHXIIM1wGERgKg8ytOfD1gLa9B51MYPCbpoXSN5QUjbTvR0p2b
WQtaKLadvqpzf7g3c09cxFKbrG/aqFp5zucdUvSKU1wQta30ywrAty+OEcZgXH726Ab1NQPkDMkR
q9Joq9/dqwcVRB03Jk1N1Y7Px+OTXLNsQx/iXG/b0mCF8RgjVd4deXrFBL1Bn3PnDBS0mJKQyxye
wwh2s4Fie/O0eO7nB61URs+gAVv7SOyJD3PZY2uZb9c6XH+ZJA7sPTWwh7eNP6CJI+nWbnyV1MEE
TjRDZpi/h8KxGwQ4EKo55V3H3sMi3jpXS+YUZqBiSIUl/5Blp6nSOMgXKyDvxjhLZnfWmg7mkIXb
hOYTnF3d2+5kn4+UsT2mkbK58HoCJellwuxYoeFLyZeji9uT5TPAUV2n4nzjZqFTmgH/7ysftzjV
O9aEc5Jto4yCvrxScWT+Zytzb8rLXFn/rS0I/YCYWL+PM3S+W1EXpieCNKcrSiOIlWk+aARRIsST
UqNSESQ2mvT2fAzj3B3timqZjagr0R6zvvXnx9j6Y6BuutUBcP24xKQM0g+9N1peIEJz8mQup6dh
0piJb2tjOAejZp/BhHznMNYhhGDOJRrjH60MJ3dih7NeKr6r2ziy3MLau+ABkIqbZnyoWsI4iMCP
nCR6QHIFTYlRAkoUv5wIURPc4Zqo0WoOf4YtJnmlJdnJCNJ3aKXGVpFVwiPBJsxogXVJfMrGVJPZ
ahuqzjjZjNRQe7zflICh9OKJO7TkKn4dhKhYmU55QTKJ94/BSYlSUiIV8FhUXGUcMaKDmnrEL+pA
cWw8LTQANM0f4fXIhjtU/T7bJToX8rCp7E42vaxavPnItYpiTanzL30nC7VTXF0By4TOcibW43rp
aH8inFk6yzXFBxgEfwwld87mhi/hPj3mtQmO7iEMWgNP2PdQpRXZYZer4N6xMnaXDXitchYLbaeR
MOzziXmi4DiEbQbzd6EMvrw8ruEi8agiWoE3UkOjxn4dsWQLUP5tiI3LX10ipJQ9OU8tE9nt5Jby
ZcmNsTFeVRK4QxeP/FPpc1pQLe1PoY1nAPHuYQsYRmxO2dtW2KIz+hzzemsFsa4OP/4IxJIZa0RR
xkOwM6yRCAjoa9yhlGdMnfue+FQP0qcQyg47MCTSq1ilodaNmYuaTaqQqLS3NofA9DJ5JRbEEhgS
ihQ/SuwDPyf6E7QZbPdT/eRKXiRLRVXEnE6UnUI1QEY7dWvi2rXKZyWWwW45fJsi6+QNWUycw3tW
7ew5Bq/b7dlPjR9GsStxJIdvoMjnOErQ/IJqfcvmmTsIHgX+NfWh+T5Bb9H2J9IRkSkqoc2LeD/4
4TO28gfLVh9jCYTE8R7jSVPocSXPZNugM5wClSzxGFZ1Lj+pl/p5Epmo7c5TXl6wB7T+bhtti2pm
c8zONsTt51mZKJcxm0/mCfjvjmvQhgQNnSw4m4F+BdgSqvx9LNhReYenx+BEtcyZEPhiLo6wSVEZ
C/SCj8tUpsFsMlFPmBbludqqf+qJMLOcewDg1Mv2Sg722O3JCgt3gR8nOjj7zEO/pk+BNl1172pr
B/gn0/wCph0+2kmTwQx9myiVOkc2T9Ahd80sNIM8DZ+gxewpQvph2wWxxmzhk0OWgte9b5MSaCuX
ZbUvWQhT2Xl06w5eFQza+XMPjZ38WXJd3B/rtYq8Gp2ggW6g7g+/xkskiBQp4IYM51OEMxhn0IUK
MJEUwTBcd6GEkKQXwKyIAv2+StnAnshjiRGpFTa/x9koVJKAx1kIWYWmL2fQ7DppWALDJiyiZ2vl
yppkVby5Wve8MTR0uJ0uzSpcF1KH5JKTqP1vQvlbV/PrZ2l3q1tENOUYH3/gYLpaMesb2TJybAL/
KbHJLNe79dJi0IfYwHWJGxOYPXdz8Q9XuiMBDAZe2lwt4HJB0aK+/MCGJ5fLyzlfhR1lfBuRQXcr
hf7OjHUUyiL/TBFnCXPPAkAcGhuIhqcthseT68tcK+Q6JQilDOE9NRUQ1buVPjn/kB29Y7NEI9h4
aoZ3s+3NdwSsh/CT5c9moO14ICnTHCxsSjCHe4OYucN69bgZNxKN2MHaP3suiOekhGOeBVVb5ob5
V+pP5kzNI5KXwMYP+Dh1szGRkRXC8ti+x+LOKqiDCW6+VJHTB7ntIqwuOYV3v9Tf/AkGrzOXalNl
y+yIa2J6dRdufHLzFjNJdF03tWMCbmbDeMsvZ2L2LRoPiPjFFpdOeujIOUeSLGyn2NjSz3U9zA4f
4B019fsfM1ON6pMODh5z204w20N3O/W2oUuRIM72dq+3WmSyWjAUt8Ip6LmFD9X1bIpj2u6fUrzQ
XqGdgNKRgvi65pBn4v4UwHC3qkEDwdOM6cifupajbhBZpfSqgnjDb+nBG7xiZ7wNw17alHxrxzGW
dN1Xdlf0hWudj38jcDE55d5uw60hWGWSWLGjdxkG5qZJG6LRKMMJAaVeJDE34wS1GVjA2CIy1jo9
Ue7ixgzJpEPdU5yKgrNA3mM8Do9U6RYmy9y0CkgZnKXyrOBkv0mX3tFtzOAdkQCIE8wCqc4/dLrH
CuTGEkCG8h6hlrxHTWWukQjLS8VNCoTEOgDtoqUHqmp6yf1RMwrKxFwWCLoqHLpYhD7KzAIqWuvE
qdpMUx3Kc+pqsPGvZ9cOMZQn/txTwSEecDNixY6o2vyGrb26xM97yVIaq7lCuvic/K5Daia7qc9e
3dae5rTTNXUmx/ajrD4z2eU97g3+00AQYO3OTwcb1FCOfywqL0V2c1X9CPR9I/fzlATjdgZntdRJ
GSyGVf1XG/dDVD7U488Gg7xUCj0YIWPO+eETIoZMmA8OotJUz643ajQm2CukrY8LNjTYW/9Uqs1c
6yf3FBJ6T7ZYzKm4qmaVghe2IbNSqw5TcM95IaeRAE5jiu8060P3ncMtGg6f0IJHYa5x8m3EXMiB
aFnR/asKU7h5sUvIQveN14WOO57rSuY5RCztvwmymFd1J0PGagdfcLjfO30dvAW5jz6cxk0rLiJU
sHk6CO5TwgnMOcIoX1AYlwTJ1A1CBWmCdN0xEy8akuz94Mo5DuEUxPHu0MVih+sarRnXt8vYmtqu
fFrQrkT79UOb55bvpI2qLwwOq5EI5MfrdFkxp/Q8XAbUdabllX0fEFNrH5lmygbD3hkSx9xJAr9r
RDDh2uuJQbGRyt9AvSKkzGc05Y1r4mtCbsrclUx0nt3DajdHJAwnR0eGbXNPwLCf94hRG/2claC0
tOLBemyx8bx3l/foK8oWR20LE+MxIJ3aU6SLjy3T7vdpT9V+ZlKV5cJ5OZX0Ra7Y2mBayuQ1HjUO
YoYq/6YpGpeuY2IKOPgb18wvOmhJcc4VZztcRFW6x3U1ynx1JEveUn8ui3bwQk8JosELW+k6I/kg
e1aZwE/GmvPGn8r53B2iil/MXHn1kmNsta4w/L+aTZYhlC4/8syD+rOLjQM+dNTyslZKCnftckSw
KAtH6UBvIU1UiTXRxBoGd7ezW9idBLuCIA2jFe2inn7tT4udyCXaNCiktptZzwLNsOXIWtz8Ufyz
Jr8UzvAOOJnhu7kuFF5CqMqsbzKXj2RehP8TjMpLFJTS2bbn0MYtea9Ib4XG1U+ETuTB0Gr1GByJ
qPLv7Yzrbh7ymPZ4O1NNnNrIbnVb7Zap4WgFVrZ+TfLJGMXkBFVKlLulW7JDe3OCrKA9I7IUA7Ln
UHIRlUbQtoUaLxufh+ZJaG93M1fC70qip7YCmlgEICOX32UjdB0AVTY/pu9BbLRE86aE7kdOfXZt
WeqwUkybVEHLxLynpih7WOwZjJeuHnFNXI+Ltbo3LIwquAhcBNMJ8FfjtP/LWGHTaJsGFXx1N3uE
XjPOeq1kxUFXjTtjj2w2eqal35xU1ps33nJLqjq12aBkzWuBYy7XCLEB87/8SFwmRdjgK/YocCD6
qoHad/brEhfH5DYk3NazryzWaSag1+ua+VcIaWnJL6TFW7zGVLi6heeluVn4gxnTIpGsw2grhhM+
KuX40ve2L85nrkvd74bFRTJ9Mkq3CU6MKUGNEnF0BTv/LvztKSaLJ/C0kkD5FPyLC+Fkk+ca3ZpE
B4cTOns0HuYs3RZFVQIQeIL1EULQ2irnQEA+R9UGWGJLqADpTdtOfF22EnuKRUZu0yWx3/3Vuo8v
CUgNTKQRGFmTOH4SO777DDniOBbnynoUzHtJO3LX17NPS/SIXWkWJ7frQ4E+dYnXqHCN29Ly7jVk
wVJ3qXuVhMp7CstxTK5dYVe7MmsegkNga6Sq7U/y00kBmdiSh6RfKcy69wlLCaxTJT8nXzLTNcJp
0q/pGwlfYVC2hGxFuhIU72PLvsW9s/g6IXuIofa2dad5cgrVmm6Tl7jLKKn6aXwPLztOt2BUpL1s
+fPaHWp4Ng+7yZI95vnmtPXgtIljQO5uSInThHUE5nWzGGRhfF6c9MCuooKWnUMclzUdly6JfnGQ
9Lenctr+ALgrHhOag8c0wOm+gNzEKiq9doG6g0of/JAvoguHQ0r0oWCnlG4Diizrr1nKPvDpzjK8
/MeAnBzmSx0kN8x10vBZ5q33JqYtRyngZ9cUyzZfBZWSN7B7MT59KFyUiIafZtu4pz4hvqefeQvM
nMt4DRrt32TY2zAZfRS1ibRz/fRXuxiE92cHZg7oxpvdwYxPfRqDdRdGX97vUGp1MCbpqknbesko
lkQ+BgdSt9DNhW0i2gFaorINDRrBzxyjEAKz+9HKK/SSPLGb44iajfjBPfDWHhPz0WbK0mkRpEjI
+ESek+n7REbc+7DUCqS6NLRcuWIIyraU0y1jANNZdJ0okJ1IGuHN0nm6yhGvICR1s/HenCxSI1c4
y605g7AVIV6s4UyiVFa16kI5qGnSO5QPw2iUDrWuuNmZcIlJxluFb8539SuHG3WWfKIZ8446Gq9E
jXwEKUkNdfLDw/+DcsTi3s3afnZfHzn/JXr5ij47YJMh/PDSo96KZGbQitC+HmeVpxuA7/6P+vOG
OSQ7Tcf94PDC2y0F+5VeLT8iV22eTJSZqxc3XBRdjPJVOrXxlrzFcHwn7b3QpBXdmFvlR1cK7wpq
aM0N2vBe3AcTUC9/ZeO8VKwhPQ7TEElxT8OlwEr9bXrU4nV5oYj2zJ6Ff1PwX8Hu33xIdG9fSJZI
hYP0PZhSTb3TV6i/8Zx9Jej3RxR2A9S04e/TVhWSR+cU+y1Msj1ap1cyrxt9s8BHuxu78AbLwXcJ
cIb9/KcqF93wexgq4xzOFQXh/1wtL2V2U1q0X6JEqLXk0wzkCmVUeKp9r/+InpQcYa/DdoFGEPlI
O8+/m6B5Mf3RB6fUzMwBWpNQUHuam4dVbaLQZ/g4nCxWMuez/NRDEPkhWfZpGDlcZJ+qg9Zura3d
MxIEvG3pGPL2br2fd8Qo+svv5UXkjPXSS7ofkV+9Se7pkVb5auSXabVTyxZMixWPgMf3+HWTt5pV
mG5xvWouvfGO2afa38JFWH35q3J31S5ceQvre3zTb9CW2zGaa18WBiT6Q1q70UHz0AXtr+Yl5+1k
c8ziFR+ikNjHNlgg8zShkfMV8rsf6Ny6XGSoLSzrcJYW3RQRuxJU4c7R7l4/muiYLfIK0rMCejHT
XcoAQSSK9BNCy3fORBeqYZuRy+NHaaz3mifHKLCjYXVb0EMFx6kfBPl82afU8z+/IBb3l+N8U0wl
328npkXGjMzW/ZX5zwannmUREz+cFVOQLhQ6h1uQt/+5xdxj8JeUaKDS7AkRTZ4W4+DJUjLSBK0J
GPRHTBaTXVVlx3U708Oq+8u7ude3fPoSnv5Xr77jwr/r4FHAZ+1xjPywqZXrmIZeb+76am5dY1zR
jUSUzv1kBWWRuMtZ7keEvMfdxKHGSBgf0W3ijpA8Kw0jUh+ibw6XCLnud6iqGpwL0mCF4VJkeLA9
iwQCZnLV23TC/xkaSalfYaGu+zG0ynjefl3AhnJroBm/NNQgTOJfWZReGq3UloTK/HEd9Elvp8nu
dY7ZPLt4NgYyIDpkA1/2owa6olwvF85r8b4zf7ZBf8fzmfIZiTjhZKwoQSgmx17lvgP76cTfC5JY
OkiAoBEGu093suoYNYFpPOyuxQyCLJnRd7QD1hVdv6gXJLElsvU8Jy8Yb+uKER31+gMNDJKNwbNo
IAmqgt7LkMmK4T7t9DAsAiQecUHQG97ZQXW5UVKX4yHErlPPk/wGPbDvD+/E1RM//uBbCZhif1Vg
i8ueGxJN3O6/wR1g6o3/ncPqqIDeeobudFoHfU3KYbjkgP9dVP/dR1dzhiVl80/CpQ0+Y3pQbV/e
mCMJULVkw3/ovu7wzRq1AhCRUhT3dvH/U1mJ4sab1DjYqZ6DvAPMfJwYtutTqESADhNCrbLfinzy
xDk22kqZL/5m9iBfA/Sz8PdxXkDeh1SYxf0yllyU1aTRPLOmXh1tFA8BoArwSDhwWo4fAHdbxlCc
unMY6tnmp8X/GKWquhX2v5lOSRkLDn2t8qamhe/hhrqzkJ785WdprF3RgeWvlV2ezKo2ry9X8SbH
n7W1j6Tl2BvPmC+3j4gNlCiqY8cgSCKcr+6efwW6cxoRWJBF0iqM3Bv1elgzPLTm+syQXiNkUz1F
9Th57BVdg7pSYhqpbViH2dMF/3PCrbUjarsZ2Vi5a7Z7bvJ/j+/t9EpvyeAAynn8TYuCtq9pCRjO
r22acREUyZJwBdHi5bYULJUW3Nwux7DLgUt6E2pAtYm3CLYdBKBtWdcLZddx5demJy46RLPN5t5i
hMnVPOTs2i2q/FN1riPD5f5b90Gu0JrRFW8THLFHT3X6o17ZhSDEOJ8KoxUyTcSkvRpFKTO5DH/d
97eGH/0sQdpRb4vI/XSfoFLTF68eicD6MQxtM5/qb928X/hV+peJUWD9AgQ4RXRVLs5ktYzMNLAQ
H0Zt2MAj2M99XYZCUmPRnwI+xrXPz2xMdKrKArhxncfvIoyyh9RS2rVyeV3YcTBVKokuivO6ktzL
vanSfYLTW6xi/bZtWpHkP1F0XJPJzTwrDuoQabkxTsoq1LIGqqnO3E9A4lwbwFgSEEx9IbiGmmsm
VTHTFsXOwGxVHbLH08bSo4nXJrEuwwNsMRrHwecKbhHpO/Zq53YHzRdU0O4e1PN+6EDoozK+N9YM
R7iGn2T/QXpS1Mc60zrtIS3NgilXE6BYdpHE+v82m+Ne55vVlAk43FmYAb+VLr2Tmlwmd9/u9WBg
UPdlsVnTZ5u1la5FjtQAHzuxp3byD10YZq5qLYU85CdFCva9zROVu2vE5gDLtSyNVWQFXFUw337l
p/FMQoE+1SZ/2fihvYb/AwDRYZLywsKKt3P5sd0nDNaXkPumgq2VaecbfgLZttSyqUOLTaDdtSg0
5EDf9opdCeQa+V0iC33MAX9lsBhvN5RxsSpy7uH9pVnxR3z65EpaZgqT0CM8ja3VJHx/oApObdFX
GRuEd6goSRkTzqGa2swvcRON31/TgIMcsZb0cghwD8QR//Z7aDNW0WwNwMTjOWwSIxzUFzk/hf3Q
IZEh92vHYGgfZ2xgY05mMqO7O1xTjj1t/OhPv+1Kg4pSV8PRPDrQBM/Y7hQAEv/r+PCX9IMJFFBx
Focl7wecPNIwT4bBq0bHrzHikSP1oSdUermff+JoVG+sef5dXVYgcSdyE5LmRqV93TlMB9qwZ7wz
ykCR0Q3M+1StNhohIjxoP6JVpPD7xdSwNWAtaeULujPs2e5QOdtWLgOMC3Nz04Ib0vIQkMjy7CrJ
anj1DmHc2/GaV+5L4PT5lXV7LOMUM6eoDOq55hGUTaXtE8q3TGepgZh9y1GHBkzLEtXAqa87MNv2
D36J0+/wSebolAXS1KWxy7cBhWaUgoKb5JdFdftCQMeSLudv7reMMZegMbH8xAPAgFK/kSoQoUZN
CoelC9gL+c1SMDKbeJKXRA8VTvbNepbzibRgMmP8BxvSA3mog5zAZfKCdH9tKgIcVHQe8MvnTE++
JsGVVkT7cnXpf7y9zGhdazfGLeLcq33lawkrshchnniLTkIsO79WAY+2radRyOqX3PIBTeZ159CJ
G0UnXukBSlnyxE1f0UbqWTZZCEcsPR4CM8t1L95TXNUKWUVtgpGJmGHx3MUQXKUjs4zv8TmhxaGI
7lqcHcvESvHCHJB0JQanuQG3fn8XE1rS8MBoxz9bkLV54z2oV5VkUCY/9I9kc13rvQRtHQaYpLP2
ZjMTqn2v/pB3O8LlatIA2gN7K6uH0Fzk8TcY6egywk5k9FWopn+Pr7Aovo8Rh+Dh1PO7Jdupc7a0
r7xAtEzNACTmgEPpuzn8z/KgnLO2Ztjz59qvNRVqrvhlyBOe0n/doFCnPcpO/jCX2m4+6eymopDC
1UVKiF4Zm7j6dQCfQuiVJJdzCz1+oWe+Q62WZZsRku0Ynmamk/ZAXG9c7VFv9NQdO7NvqM5kLo4F
/3nMXSsCcgKADQUM9j7dqyrI37FyqC53ttRXJy6xC9LK+IHu89gkPnNCtQ6TfA2g1Wo9xqxPq5zw
M3017/ivCnzvQnXPCHDpEWGf5SU0+T5AD5NoqHOW4wpY0U/EmpRQ+qreEKUzy1QfNo96KlmlfU/y
wyCAutv5vEJLqPPjh8Y31nR4WqoH5I9X4ePRqOnLNb7A05eA7LTta5vbwQkD9gWPAQP6eoWOMn48
GsChF2A+zpXJJAIrum+oFp+DUJ7SwYCtXsnqklnzhHcKRie/lU6AsCLpHgDwsSKotYwSSuNU45zN
g4pb4RsK3fqNcl4+5npQb4qZosNSf4vCohD1N96wUV14YnO9MfavGamDVovOtzwEuR5TpJXROc5s
NMf+aToaQ3q85FTh63dYFMRKh4HOh2+rV/G8bSjg2uTPtKaNs5AMU9kS8X7/4WerrKyYIW6VB8YV
0Se+qQBngv/yXH+sK00xgWjXMsAT+56kLjmCF129fxuT0rf2+ld5tA01IoFLIq+zEUqqrrKN/UXk
qw/immrHQvOQcP/gABd/n2h/6Q7hOdtwh7GEwUpHeNbiBA4aZ+Hch9T1NMozql0MZWWHFC9f4Vbk
/8awJ+W4PkrrFVwwhKeJBaZ86ybl6+/HIBVfSFUPMEoU2vSP4WaIUnnOTDThxJCwwpsJBu5SDBGH
gJ6krfPPZGX9o2Z2yD0lC8YlaRBtC9DLgF6EVq3PIIBTisI2ysQ2wlBjlmk/ZyMqVe+DO/KI1Has
hjKXEZqtGEtzH4aYQzyRFimSm6EnFdAyM0/3XbVMHqkpnFissIWdfdCwC1ZziGy0jlyR33eatn2y
RpJPW3KwmB9nbaVYDn5didxoeBxW2YA+Q+bfcRTwY5unHu5NVWxsDHcxN0RCNjL3dcB/YM9hmAbI
VBEN8Tt3SmY7N1hDkqkRJlV4qoCV7Rar8vrXxm/pv3n+gW8V4dkW+co6jyKEdOB2keTpHHDMGJXL
xdpiWwZTDpokZ4TuVzSSArfMk2Q4ggXGnPCM0BEojO9VruzGOmy9Jtl+VunVqn2Xx6sdpQQB32uH
XBUlSQbOsO5ZXa1DPtrpMFUZm3TzoJqwJf0Y0KR8ShXUY8VtEQfPjILllEq5GB5uKUOZDvuM9WYC
NQZ5mit7AOEEBLxFAtb/bwBrtozmsCzElIQtt/xx2sT5IiKwQyPp1q5uR8WTqeRjarXBJ2C23XXo
ObzzeJbkgkXHDncAV92luX+Uxr8f3Unu/O+z8vhv944i4r3AjQww/1P68icCa5BJaksky+qAmkpe
xEugIMN4udPHb2M2Zq9HsseHsP9whwtPPHeHfphXafGxBzzkrbcmi/VXSPzWw8Hst+3U43zuEoC1
gRmZMd9ofUh57f+apqxC8KzlOTsxKUyauDfkQr9pMEutyiBgyunn+ZIlqHK9dzn/kiqnphMgGU38
KGIDH77sk1TwdmFEDdLWIOYTeh30Q6SFvosqsN2XfFKZtzviJojuorI64xpVAPfC4cSwBEGDQmXn
vegTCG1zLnw/tM8Xjfq70sKFW6ZpN7K0+kzwBktRKVcAfYcxda6JH+0Q/Tz42FQlLVoEzxHrm1wp
TaF7ZbWU9bX16KrWAFqkIqVy8PJn1/AKCO5FsTp2LyuKNMRoGwrj7mjYi1bXg3QJuit4L1NK2vSM
jkkKeE5vIyp1bfVM4jZBXTJzWCZv25e4rHO+LB9vSwauSscUa0UHxAKCGr/JLfplhSenNaQiR1xo
IGNMcFWj8IEXPAxYLeDE2F+mCeK25OrMrE5prvmExu/HAHzC2eHDImogC0elIu2ILiM5GEZX9yt4
O6kiYnVzWpwT/10GCMWyldPrcrnQB/bVqV+5ijgqnDYGwCRwaRArcYW6mRrWHOhTzYNONNVLa3a+
cxh8UlapS6UQZ0BR0EsOJXncBuOl9kDNOT4On1pst7mzkQEMq0kzWWldPSlm0x9OlF9L9wB5St68
BskqcXXRvZ2Tf9QmZs5RlCCOCj8Zstrh006asYLGQPlZibVV4Rn1YWaihcnoVtgflyQXE+nXlz+y
vG9LeNAvbVRShQr5Rrvn+P91aEYndjSWclh8KVxRGsFd3YxBsOWitzNzA0+cQcAA3dglFHYWDohV
dZztfmTv3rgiyTBURCxSnt0MtBUaLzKAT8c4MVbyOpxFjFbboN1FE9EbUeYVyKwhKpfysfmgeiaH
HJ8tdUn4BwG7bVnxUxEiSqsp/NAqxMZwPUd6N3uFtUrQOXzuLe2aJ2+vYr5lJXgPtHkiz6rXUutp
AdQWNgicwE51kgBJBkbqpPo4i1+wpckfmVro0Odm6+AhLD4lWojDrMoCd/BvrlPyY+q/iTdrslM0
my0vGcLG31Vn9br3pB+g5gTK0tSKRgz9ofNgqHSezN5CW6h9VyveiZYStQ5pxmsUSkGxrBQQkM/7
1V6pqMm5aUH896Bzh0lNwW17pD8cXJLN4qmb2wM3V4YRWY+e/VEUKQXioZeuzemc0YVwE8oquwd3
JyRYcRnRs/1ydI1VR8h8DwfdT1381zsRCixRfaNIw32ag8mgCyA8M50EgNBSlZpHFfWaaKHLCIyk
dt+tfkly62VevjbKHtMGGXRZxq1UCnNgE2lEJxMAHavaaMqRoijk315m7X13J4Bul11wKUngbDgS
aYWEpba6WeU+UJeKq0TdghGcvhfHhYwQlLXDTnM9I7Rb0MDrvMjK+1bBNSsyo2P9fp0FZ/4hjAwt
o2Um+cNa4vuLdnSV205Adn994FmJBzARAPSXuPrPXHWBD8rXB968KKTV86L1fT8K2ojT6cSIn3NN
3wvGJjZVLfJVoUkWKOVZcUpryi/3G5x/7+Iyx9QswTxG3YocSMH3BTXiOGyT2Ux/INcBDkEzL6Uz
+FK8HMFgo2fYQGDmbosUA4YorFOjCjs0RLIfQMyGxpY4+P7y+NTxInKtuRH6CFmTyPrgRzwR8emC
thMZBWbDv9nNtsPxFo1gNV67H2AWM+EBrCdf2ARL45Kd3REBV2/flNUvstM81tVKz/USoP28/g+N
1VimNEj3o2WAbNbioBwuYso2nEIbNIqygup5tj5sPpcom/3k3pjniG7q9hFunwINokWRPMLl2p4z
d9fdXVZbRk8VzztxM5qs6ARDxZZrtjqU5OsGsaGH8qdyENW5xVH+7/eYhesUOV5GxNG41xtoFxOl
Gl/s3jnECgHaM2iuuysOtkoKFG93rFSkjMzi9Qh2qd6XDvg+f+VIqjaS0L+lswsB66Up4eekgryO
THKhC9N+hzj+apGfGiaVW055cZ4N2N4+3nWSo9zlJv4zM5+DVxp7QK5Khq0vfRbAduf22Od9o7Z+
u2h5rDlNNwMm2+MsgEcXFAJVlwUwfOXMvAqBASm6dmBVDBezcfZUhIxn7KZkmswexz/HBr4BL8Q/
drSfe414bpUNVJJGxb6wNPMEGvkM27AK+9qUcxYJUOr+Q7+iX6FA7id7K3gteA60X7UVF7nzyA1l
iJsI+sBPWbkrXYa4BPG4P6XCeKjnRKcRpRyZhkCH6Ko5+pfgtlugf2KT9eLjhtfwlEGFuLFuHTxe
BKIVpxwkuKoBO7XspCXb4cO5Iz2R6Zu2oS3ahnilB5meqvjsmTy6idqcTwJn5dL4q0BlX6ZcJPv6
ro5kw8TPvQDEPKR9Ns4g2c5wXKv40ufpxT7Yb8L8KqRq+5rvFF3m1zudYUppBocJ0l7CpKKfP7Kq
xi1tjOOU0M1c87cetlssgnP+PZYHjn4PUvo4wGHEQanTp0u2N5fwAFDhiDZMbQkXijlOCopNKb7D
qjp9xVrwvYmVwbm31U6oVSEa2wfr6EUkBNXikOr5Ijyedy/4plnoDYox1RfACL6tIK2//LeOSoWB
qtPxmjLixjAoEd5CzWwh36xJcXh5xyG67ew5B18lEkCjgMMQpM5LmXBH44aLIndSVBGaVsUg0uGa
h1KJjoRY7OSHr0iNwEpIt/a4nBbI9cMhLtqjqlAN2kpu7fT5cEMGfoMA0MmH/M0dA/kJUGPaRJPA
oXCkIbZp4DmLw+AMWeYYzL2aXfPEpTdpaO02awhNOFUbbEDdu+XtyO38ihBx8xIeS8zyZUoPe1m/
g82lolzNyYBm7cvLxtaTTiIXwv4DSkf+WO/GOFDd63oJO8R61NZ1WYtEFaL8cHPm6rYTtIEJwlh1
87xIWUCBcFyO/JnznyLGvGuUoho0yoHkMMbrJSKxZWAlVeSRW6FvLk35LMVmYBN7hbl4RsThH9gZ
0rH6yzeXHNyC2IJuNndx3bOPyg4c1sHgafB7/qlS1Tau541UoWNkWFTqci6eHKTr82m9+a+SBXYe
CdtWMpTw085VM6xGmJaq7cPt2EZL0aUdlTrMFPKF6l6iiUlzg7irQ2qU+YbXvbEwYBKlWd/OGcvz
VJmm7GDhtancT1CJZ1mqXitT3MGskyzh1V1uwJn8/slASHRUUC0YtdbpZ8BC97vVPnd1ug2tRZjf
5VaP35NtD0RC4seXiPE+MVRh0YfZDKC9eJq7xxxgDLUBWlClx8leBuHWwdnSLOdA8Enx7clA2kw5
xgqRzonMy+Tyhk9wi9ra73pokg6n8fqJuSqxcs9ESHgo9wmzKZinZaSMb8deonJqNLj1pPGPLy2T
F58C4iduivsJWYLgVJ0Xwk4NFXtBKoy8FV7SGIGu3BRlDfHjiCqcP26YR2w6F7FuGxRQ1nOloBe8
8E9d64hWOQ9Y/KrZhCJvXsZwhjx/d8GKW62OsjJJMYqackQM9ThM7mxL+0iYMig9wcGRm9GuUSD5
pQ5kITcU2rSp+yC9Xst/cWlKhdycbiVbP/wZ8x+K32V3adjhayvX06Xa0ouPDhul5fHO7IrJP0/N
bvnjxJN1X0Y3Pq532gMDDYvz4EfhYLC6LHSKTEtVhYdRAUmzF9K3h3sbaiu8gL3Up2SPTm6swRvW
m2YHDJrrOiHhyCRLLugAiVJIQCpIS2TApnypmxrobTPHL92G2/+9bxAHcaGSECmyfmt3I1fpJjiM
eCuMiNDPzAwkBpjm8LCv7cOV3+LqZjjb01ATRkC4rVJgnTq0Qpf7StYtxQSQ0IdSp9wOcBUmRe/Q
WtI8r8PWHTqbShIeUAoGKvG3gMUUmbWtbJcSGryTgPGh/EvfciBfFIovNHyxsGmuUFiAARKQN0yh
ZJSr+qifs2+A6SMxEO/bcpuSV4eBpJ8N4uq8AEecJT/lDPsbchkON+TiVNtlhZ4qh4ec2iKUeiG1
Lzwc+af3u8KHPSkaa/L0qV14as99BEzcNB3TZaJRn/XKUObaTcGiY/9lBXq4gXt83CkYVonhLF8T
1nAmRuH0qvku9boKhjdDue+PKFD+RGqM5tJFDDqIIK4DsPfQBmbbWTIptxVl1WuO2RKRnzgGUsri
a5xpT8vAefhEOsiH60253Ar5Kagr48MDW5WKRnOkE67JZGNoe6Kn88XR6Dpip7bM8dypSDQjNKro
8tymWkUxC13ZC/uXSicOjnvzP9qSVtCchlhVoTixSr+znk7Qgc20X9Qy8Dd6dPSGFYYVbrmK2drt
dd64QvVimjBlwdJV8pwDNnEkhb41jmf3wIywEgRnI6J9zLU0bpDFuATRe0XyQvgea028qrOEDuhp
s5Pb6sIQasiVfCQ7z5varIdkx02Q7GImAII20yp0qbg8fVXcxNUeEwoGtluP3qqBgMADqnHKepjd
vSK9pD9WSf8aYnP4W3SGDyiXRJoEvmHF0YAvrJy/uk0/PozpH8+ST37FbK6dJ9KXD9vYPwH8NqmR
QINwzZdMCQwVM3VzTtXtTG1J3WjFm7NDAuL+TwT0Gfu+8effzRCp997vhpZHGm0pLjeKIzD8ZOdL
tPRKhBcte9iSMo/EG2kvTjNeBsHzdlqHsNqdy3ZazPxWZOnAUOR5bcRTD6enZ9J2yhXy3SkjVqFP
ccE3DA2wkFxUAB63APOnsBzeteII2o6G7nyFyQb7BMp0M78Swjud70SOykcXAMO5+Gp6xRaZ8vIL
z4jPn9r2e8+CRP5W9V1cyRqOE1y1gdKBuejShL3dW3KxdeBtsvHuHp41NN0nXmbawt7e3xlGKfPj
VtotphsgM+iRKlxlqMZHnsB6uIot9IVBPPPHi5jg7YhD6Hd5sPFGms7/EBwXgujOWqz0On5dI8aK
4i2Hjqcxv77nhnvPsLscgN3jPyw6hR6vKqsA91gxXb+KAYaOMA4sEaB/O4YgSFbC71j/Rpo6fHjm
x2Mk74c+k96oUFVVU8dxDyCIoXxodP4AI3u2pKpQDpUqFP4zfr3UHyNKJipiAPZHBl7HhaJnd23V
I1P9ZyWpgvNoFMfda/zWMWIoo04n2MTrpxTk40PezcjmYyfobFBqcFIJzFLvDfmYCLBSDD8+wUDe
oHjPWITfT+IhYRpxX6716akPKpXsFHQdN7LGJeXoAUgULg5c7go60FJSF+wNNpJ/BQ+DGnynALrm
AAS8c1SCJXLAvqNMjda3BEGG34Udp/PlhSTFkZiOsE1IqweG+yl8vzAVRIXqxL6wvWmWxfJj8gla
2f43r6ALi/DaXGULJlC76KZS2EMmS18/MiOdfcXbWGIII0mJzCm1N+x4CCGtRtdSkRjfsAbLATMp
Ux27IskFXRh80SRq6MUvmpVvjmZ/b7YyvjHOlFT/iborUP65VvAFhhccW04CT4NH7SVJCDs9PhL1
d03xBZAEJvE60rCZWMj764p939N5LMo60FUFiDNOvQa/jlxtctyAT6K6EAoPnza6cKaJl1/9y8zg
uIXlSN/XwjXCB/l2eEc8S0nemABBhWgtfibshN6udgHedCH8sOUzTgMMFyxQORqJduWL87g6ybZ5
3Fu/Gp08UWw7NZhd2LvP0n/ZHxoeSm+mVCS4xd4UDIeUHUvwNC6jmwbkCj2rBKGXOzom5Qu8GBb9
zKMGTPKePXGRdn/RCEIWp2hcV9eb/cxD5Kmjv7z0xKKfKntzaw6MoE84g/UP6fp7lk+aQn1YGs8X
BoiWJgPke7l7VbvPd1un66GElIQocKEsCFAfsyGQxp7HzD8gCGst2Uqcf8za+WZk9tsFzRHvy/pT
NjIXXYc2BvjLurb3zLb+c7Wv4wccpzFswb57bH/GP8K+d913unIuddriUlLjJX60vKjelCy+jIFw
WBGfyYiYu8Oezo55be+V1aFq8E0SMp02hVetItTTVj8nNmPPG5gRFFWZ3oMzNpCGXzvMi5EOYzZy
6egVSS0OOjQpckh3YYay5qIdHy9dy/F8ojrxB4DJUuK5JR0akFrNXes+Hj4L7Z/htN1aztzKRiDy
z4qu8fRhH3gQBsH9Z+2qNae5R39Utq4pXTZ/XG2W0ltInO6YxIlCCO5wiTzG/1mykN3W8cyS9Wz6
6ObdKxInRQewEFBxk6YZim13boFoKw5BgFFOwgXGXNz3xB3Fk43D3scqpn2Nz0Ndp86OGbcgR/4Q
1I1EuBO4eulUocp8gZmMgFTBNjLQV8CTFQZ8kD6C6oez2+uKCok9aa9n1J4JOKZvgXPMRYLkznw3
apCt0/oOlAGyAu1QtbM0aVwX+v3avBiR5KC0im2iJdXc5uStvL+euUg+2x28/Rw6fTa0wOXHJQy0
eNz/FflQXcVevdZyOSygC5euchNL97Pe2pmEaKHR6QkZXUkr7Wdv5lXfbfbAL8MihvHWlcbirMtu
dw0/zRXyO58OcsJTX/zziBVi4KMsZlnoLUTxj0D2wT3KaNzfGNlDDPegEMbhvkkL/7WQvSO7V5h2
4cFBaPHYxH2jr8sAe/9ZJyoo+PpbShZBV/IsmMBwasfMuBwcKaelYdLPAUwM6Ma/b3c6DEE+MK0d
JhDmquBelWKlA6Vv4Jo7wyL6OD+QLRed1wybiXLMO23YZuai4Fb4wK2uo2CVnohFQIx2hLxz8o6F
aBlpkJtzT/JWs80iH8G3bLJVad0E6vqXKri7vRE2lQAQO26cnqQP6pu7/JCCsZABtexfB7D/O0DL
T2xReSO1uBSXqxsR9y6RenIl5PaxXTZTq+NmRXtH5GR7AVH9oaQh8Jhgt2hd/EjwkBBWxWmjVoQP
82zN/2OHpsq7O9gFL5oOtlFeOnWoi5lDhiOdpqHMeKHXD4r9GWX+AILlZc95Nq3HULH7JeW3Dxg1
jySC6rxQNNyHfcPpQCiYlqX/qmHIQji2LDP3o2WY+ZGPG44prJf797MpxzEgo6/mixMY8nGdeTsh
CltvxxJLIfO+yl5/muKWFGcBQDLIcLnRSIkPqP6trRo9QiOtUeGHiLDsseCnmiT4AMhHSNB6Tvb3
SJ4bG7GJUUH85U7dqwZ/340sQyj0Qo94Xm5yoAgAUZJ8MobPeB4UlW0YHejMXDabZOvRwnzR0Ckw
fZWwXTerbIE77EZp0hs3F7gi77j/uftYd/zXjrY5hDRenSVMsLfjMnHTd84m1NGOuQ7h3KOp/jyG
zWVg7Lh0KqIq/IiGxRw4b5E565wt7a/LD2jIgZo48uGekk0XrpQlgZtX+QWTZtxwz98qkJyzq1zl
mw1DPmzPoCtjf6GwKKxO3StmNW61W1+amRmvHpb1TZawbKrvVZD+wrG4cL5Goj/F+ETWdhQSQbVX
H8eOx4Aab/I91Qk9qsVI9amHHkCaaPg57gMrGXWy0f238Kv7wMMOt+UejhW3MS2dhQwo1GPoXbf+
nDN9Cscrn4vgG6Z6+bEwx4ZxmkIeXz3nHO+15ja4O4M67MlW2dFuh3Cg+XiKHDVGfM+cXaFgfLmD
f45/0YRTbMznQw28tzT87+oSTOPKrV6GMj6niRLXO8FKcLngvArdHw5CmYVEfL7xP0tY/oReFEbd
F+qGID3unq8pSp8mqBikb+yoV4NB3GGaKjmZs0z+pT07zWy+WoHD0d5Zl8qL2p4ikdzaXHRwSMdg
kBcBx60E6Lt1eGG5QFKcTnMoSJGswLfxXOFNUAHo4kfkxczLzhPSnp1DnfXcRCL5zwOmJQ01D9FM
8bwh6WL1yZwmSug07OU39fCr3ftArUrlEwxOOiu1UIstszyhLBo2hEdbs38QskCno+VXP11p4vwW
Vp5g/aRIpjr18Q+Fq7A1O/ypt7br2dyRkciG45J0MpnxITqpUEMPKgy6TmVwleGIVWXAWggNoRTb
V+6YioYbtPDxL1KYId+ppVmwv3NrmWES3fh1xb7oBLDS1IgYHynWmOJLFS5EEgyE0WtOzVgfGYAe
v9IUpCHpHk7gZPG65+kc6ay6lAs18rpdJ1eclmafvzWZf49A+v+PDWeeuK3/yfmiZpw1EC5D+Hsv
/MPoHuQr0MmIrOyvscqZR76l9Rf8tspg7C2AoKpojMKtFpe0BqMjbnEZRzE0EfVZZFh2tPY/k5bB
hpXiSKUq4ONBDEa9SXqwyfHVT7AMr/JBOvi12wyTxXpgzs2DhUzytT3sHVLelc2OhykgAAv460fN
OnuBUG4CmhZmVnjxyWNZmuOayB9CIuONM81XFFuCx6a4lJq7KQWAxvzWOEYLYttcqjeCncDUgAKh
HjAPomlFP+dsKdJSY8qjPEnGDGiZldjmhW3F61RJF2/npXHA6k9bZJ8O0JD0UggcWd4qw4REDivJ
i57oG9zz54OuYn/aCBE+ijClNEbdYoqGJtgdWq0iW7AUbDAipOP+EtxVLg2nND0GIYmwOlPrY3ju
wXzmvpKvj9zll3VEjFK0RNVpYEyFV3oclHNwxVTk6xV91AGbv2kj0yXn1u6OGjofH5oaVZ/w5PMA
YmWTKtt1lLFA+J9D5ICjNM4cXTYOn5cEGdpifdHGtC5PuX7l8/aypcj6tQ5igjgxBzLJBH76Co11
JEApnzEKiJXm7WCiwOOC2cPjRX+EwARqhX8DpLhpfg6hdEA9ytD3/TxPeWqaU8ID+ygVeaol/AB0
Pdv5WliVQORn0YzvOM9I+jZKpp8lReRaUZJ8zj6x39aAQKAIrx3rKHFJkb8yV9EhMKw5ropLyEfc
XIRYmzjRI/cWzvkWXuS+b9NLXKkVoJwG4LPvJO51nvPKYh10OgKn5IjP9XmIpSCII3Q/PK2ZYaCR
OrO3sN6TI7rVtctikz72Kwiaty3X9IiZ0FFLx3W6uagnUVT4WiSvSXFVg86CqboZK08EDVwLel6H
wVo0nNt/KyLjjOqhrZ7lZX5lLSVdeXntpuLEY30SuhDGuZ36V+lWwahHuj7g/WNjv5s3Z1rkoM8i
pa8Ei0v31v6ovKagTN3Zt9y/gwVOqCyiLuqjiPMUwS3u2/Bm4mWVdBDOlYpiIW4LvgwrWAgIqR8s
MagbT0nHetpcAdY/+xppOZHeGRySR0O8hfV1WvaT7eP0s5I9AP++OcxD/tPJS6gCpRjrvaZp/g83
piYA20Bd59nbKGQOK1rW7hxaNrL9IgpEpeakatYvyD4zbf8MsXK/ao80pvB+6Z0yHnx6Ic8XCm3y
jYzf+WZoVkMAPPhZmETmaeziqLyClNK5VjAQSA0o/oIQZ0QCfIQOL0jGzjOUJ6UBOLX4Emi9Ls8K
Ddee2bnmxZtFNuSlVHl19gujxW2bTpF+82eOzuvG1mExJf+XsSLICGK4AVYL8xvzeZLCSfz7Uj/O
eQBcmsS3OsUBu/gZCFwIQNlkUTV8QqUTV4kkpYEijoKZxm+hRfZpTboyzVn6YZ3z52SRys5xxXt6
F8DuXDPRR9eRq35n4VJBCnDs37SLAbaLRfSWueWjSLnFCW7loA/lva5ptLl9Q/yh7wPE06LqxYOC
BzXBaGJQSykPzqMWQdGzt7SYX6lj6pcBl92iwzfiJhPENXN7wV9ZAa9QkIv5/uw8pbxZSpg4TBMn
Xf8iOemlJgnyO0qQVphkg2+OT9ABRjxpsuDsxErmnq52t45XYeuFkcdaXEe4a0cE0DVlLjq5zOq3
nug6MKDVkdRlBbHU6dU4vIo2mnEm16NVJpn+QRUCN5qVgc2y0XLtu4eW3R1ksvOvOdSzvfJFzr3j
MvvalahfFQPyO43EzWXDNKfVi7h6Cq3ibuji810zmzvRc9Ct8w3Yg2WdJy6FABWMI+k9tsuUEYbR
5dn5GXSWvOAtzNdDyxXB0VBCgk6hIHTL+l8foYKofWENfB1Oj4CWKOZT3GN5+nkRBTfkD2dV8Jd9
ejCYBPo6wv9+RCN+amph5i+qrCfXPY498P7iRTtE8SC9dS+0Utr8w57aacmqt5gWQUSCVNHVDndO
3WYmSevDyRuMHFH1ctJqbbJ1Mwffw9fUoTKK5va4iZgWqHtErK5jlytrg3JtRb/3ccmO+F+aBSay
IUzhla+WGDXN/DjpImIQW1Poq3grHXB/odGDTdI1Ftzid5Nk7SbyfWBClD6sA4EEDpX2N4VrdX6r
fGztiMsGbLr90GW5KvRiktNQf6jmwlVq7mik98IphbWLq1HoaWFkGq3EJtpy8vPvx9e3ZLqivLyv
E1nUoMPHXN7JkovMuIF6Q5ipEy+wmtg5Qr9rfZAiGEkNUKskVaoY2e7UIeoPyF1yKl9Ln40rDko+
JIwLAYe/PIvCf+h87Ab8sc8miSmqHIzKq87reuT/VyK3G0QpkfY7THLq4RqtUB0JVg7cH6hVReen
PW461QSpOLvAivyfCAaMIpvs7vswa1sBje+AkE02q0WaaJ+B5sNW+OQw4deDpv4AGgSvSmyGNtP2
zghzWvoblgqb4XRfOpOGbQY/FaONNkdXebMalV27yNbBaUd/cNnS5yQkUuid6P/2NksJHV1IKpmi
INWY5ID0BjNQzwhONp0sHlmtVh5VPmn2w/o5eUbinQZZHILw1ceHBbyrSAmUi+/Zoacz45kW55hT
YgsQlgT2RTnPiIEFYQ1I4iZsdhJsRiX9F/ShZ7yb3PSFXBZQEsrc9Y08N4KiDoRuB113K+CdJRTL
ddOs5j72orSR7bY5ldqFLfKdMbe0rizTikesJ5GpomCYrkbn4n6gCT0SzANfKcG/q6grjv9H8D9p
ujNpf68Zahlce9JetBlWwfmGSz82gUc+kzWluRcIpaGClVCEmouATAk6yQmbAZToGRnNexAS0+f/
4RYJi3RunAaDRS6u9nHMtYCWNsSwpjqCylzjLD93F3RiOqFJ9d5oZnhLW1jSLlRBnnCKpytt3OHU
7o6FMTeCxQN5s8sRaEGv0fnYqhcpasUEGupFXYVMd5b5+l5r50OvENCMf0DncOpWsbb6X5CwLfjW
V9T5dkoA86cJ+3GwyVckNbglleqQZ4FomQULGnpgja/umIsDccOKNRh3EropCcitVu82JDPhd/UL
VKCrCzBVbE3dF9rlRuh2Y/5PIxOfIltMmvpxv0+2FAv2Ebey1nuNyVrKXuFqTYKfxxxqzHE0fVuk
jsvOrZwrCke1N0O9/IPq+dLZRplar2p1I/iypwcdzKuq8/Ljhde+a9WA6FtL/Ye1CRX9sKoIlkDA
Jk0x4MSmdBIIcVIz/lOEUwfsHFE1Ep1Yofs9RKhZP5cK/FVifDTTG5wijsNETlVty3wfVS+P6O2v
g50azGDBoNHuM+fUqM2TKn2hJf1XSlznt89MOSuoyHEtKWJhJtQcHpQ+7eT+ovFUgk9ik1nMvUBh
prYVDJXflxcxEgRFV4ZXJiBaO91wPXAx1h+TiF33/U0HOmhP6x1UbCd1ZFXRD0DxiY44sLkUh7sq
z+jzrqX5Ezt4ep5fP+mBnnKdAbE8l5ktPVXjUIZStL7yQ03oQWmHLlPCxqMq4Ljtac/O8U/Owpro
Rijf0dXLEqFvxvsKkL3MqPQ4hujVd0RX9ukEBsFAPKUz51zxn163Gn/7/1+F1yshEu1WbTa6ZUn8
XrdyWx+7nI9l2wq15K1BcsHm+NOPObTrtV+iIxo7GkCoFhcGThC38k2EIgoMy4E/uskv/aO2kp9p
bCETgjm/gptvZ+NuKfZfIUw+zP5MjZ1ZyvNmWDWp9pUPue3kwABOZgFu7xj5htHiZWYVKiQMRJR0
9nzKsLmlLp2Rt7OMIQ7xjnKRWvLpySJXbTtNEkiLgAwlkyN01o4xnwvNtKm+zNM+oj9qWJoT7Bgb
o3iFMMlvkmvwFud0/PBOk936IYVi0na0yPPY0f5ZkwTjvOyY8QccISpaARwxlTmiL/B8CRoZz9mH
zDmrTIwvHCMegQWyJS/2kcCzQYz/YhxT1ymNUD9li5HzckTgkSPskNDtsq1hn+bjM+VBd7S6D3fK
H5kPr0GXwdf1UiqZ/F4jHW1rh7CuX/fAtxLbseoUA28TrEMbq1qGXXfVG9L+wn/3jtYzlLq1hgac
JmO64mzEfnnyPh2cYW0n9yMxEc0FcO54awwacwi14R1+1iv4CJAfiwfaLrCYafTxjWVleE3rkPqF
pr7i1qAskG21WbtjHhqG96/qc0pMxHDj2UAnZ2BcWsF56hwKqWwOmwjuTdrR8trxhrbhcVpLPYIk
cCZJ7aCvjVvnnB9PBUUXti+U34hZQdUTjQiVtfu1+DAu6kmsLY4d7w+0UcuLal6ol9BiutxGVCVx
YkCp0GRFoq/e2RbY9bb3W5gUOmcdLSlU4b0ahNaPZnYwAafNqalrKpSe18Qw/laFdFpFbuxG/yIG
5Cx7Tf//t40V4SjTfeVcJqIKP0knUt0W7HqgVG1sVLxJPqzdtVE/z3xK8/4nZQ/xo2Nvntd1MhbV
B0qKgtMvga3SFczcogxfoLwpNj0+/4Yc97hwJ5nFm3mtd3R7nfjJb4kpCrgTNT8qt39Ocuw+E/6u
y2ghqQEjym6G34aNPpm8dJz7/Gs7ygO5S92LbgcoBpL9EiMTqCk/s6j8rtu1RrRiMI7CR/ejlExg
f+j5Hs2Ej43YQ/KD6h7XqsQJeCXHIuUCjnXHlbtmktY8xUfSOMxSn8hPW57OhgOVl7ZxPj1saifo
X6ddBjgnqwmnP1979c/3Ik92v2iguFOEnG3CFsglnQbXH4ADOnBZf5E7CIkEzc8FZByObkfyqgNE
wLF0/IETXAlhYnN9F+SiEK293Ziew2wgA6Kg5mn/XG7RnoR95mgOTmel+tCo16gyHxQpK3sqUejl
kMlAyGolIAb7FCQD6QjO8J9EFYQvP7urATCo4YUPwXIWuOQDxK2Xs4DR2yTVrWlYrWBiPzB5DTLb
FYneT1CsuurDmScX35LQIU24+/gjY51qKJtwNJAiQXFAwHE6WUVowDtI9QhMnZQnp1YjJPW4zQWM
FHX4rHWjh2UDRavEBl9G1as3dz5auL/HMxt0YDYcxifmFAeTFIMl36ehZj9tDXwEukktTRh5RXBg
yZXcpRMipY+xXHR7jZ1UZddSxrWpv6ViIXHHVgGF7OIYHWyuRHg7SYBsDgo438VsCLdOBYHpXehg
OLUmQmOLmTVeAAUig3Vij9CL8/M8UnjRmFVDDwIXhPD9wdYzFlrOR5Mo3U9eN4pTIFeMMgPlmFQ3
ndxYnlq6tI0PZdXtKKjP4YgiFrFjO+wYuhXHXgQ2tHIMMPGrY+4Z9VPmrv7WNE7xApDPeE1mYFf9
Sy1Dy2PP2WXdeJu9ee8vjld31MnvbJU426rBMbbd0StEJxh3HU0pRGG2oCe/rMNZhMCBkZda/ML4
bd6F0ulBO28pk9UtLKgCAK+lwNDeihxyZnIxJsMB+O5U7KO9lxc4I/H+TxBi/SmUEG5GwDmXSHIT
th6/BbDwW2OPy439ZosGVIxo20vL7BcnmzCuI5pGYYAqvWFJdaJhZAOwklSCewGyLhvFRW+se1r1
a2S7tGa/LqyVVS4fNvZnSWwRZz1bxx/9zI8L32d1WGTnzzWVtbus+pcLhhJ80jks5GxvEV6w/AtT
uVlQmwl0NgXs5C4K6refe0LDyaimBQifHgObW3rwQfQSjNjbG8I1R0hwNfDVPOzzXYWyzLz11swx
fCSTOiSPDh/lk7v4xIBEsvO+XJVe+jQKxMW9jcApNUf1DRvX+KOC6V6HTtBhPkMnmefXho0HPD5m
gvTyWrx9/EgnmP9EYHpub+QxsknB0eiuqCx7XLcG8WIJ63PfHi3jBs13ejfvlOnv0NJSNqjoG4ga
qSzmmWdU9Y+b9yLoCEx52hK5ka9Qzix0lNj3fwmJXHMc3tz9fD3+Q8H4ThRhDn8IoYThkEOtt5qJ
lpd3So5+YEi5EvnppV/cIq0cEVnwAH/JG2XL6xD0U9StTnI2cElLWkm8qOkAThvmlSO7rK717YO7
dTsladEsZvWsrj1Dz2QuC2j1FAp+TN0GQTsSpDXM0Ba8650BIjoDKhFOt7j6YKs3FRlwDJ8GDawO
tHDmhfi0HmaptuqiK7I7CLCbd+LsgO2rWfmJ1Mpbatt81X3nogKHpPhKOwHXvNSY4wPALaUpKw29
9VHZoai+UfYexNgZl47WdsLM3TrIwyLtsCgZhdunmJZF2wbFPCtlNCC8EAOTH2huSqIaoRUMNu/F
QQIl0hRPoJ5Q/cvBGLsop2vFstfluCuCybcjdYFXk5KobN2CvdjezHggWinBvMcULdEcxNcCg/3A
u/F07s1GAHVJLSNsA/S6bfH2XQRwT1z7LmWXiu5m70hR+URlQFknRzd8Uhi1Wg/1CBaasYGP3vCJ
S1WdPeKI5G4rEb8y4uE8fB8eOZpKugbiOcbWuPRxOLTCQajzVxN3vSAvQCmJAzh/3HKwTg9pFc/1
DvBoB0TnjxBUVNmjrEjwH0eAVNedxqKxlsbbgFQ2kbMZuUZlD+172Sho5/pSPZLl6EC3w13XiwJX
0MztnEa7pbgVKMAPtMnCfigjlNn2QXOx/Bc6jRMN3ixPYHBhbQSl6IZDUvPHS+y/DequnXU354md
miEHpBcKgaKe00QH2ZrKMJnuPN/3ZLT4oMuzSSnxj0LpGBWCRIXwz3AN1nsSp4+V58MfDqmsdG0I
7ujVvhIocxxuThWUVaAPx4Ok0q8afNr19ut/46nl5C/i3l7ElcBAzahoyfFBIbqukyvj2cvUrZ55
vjwNkBKX3ME91oNJaQMWWHswxV+fHGMv/nOGX+IyAwHakHmcIsVLR8tRurWoyeRd/OB+z2gR2r+0
i/kqhFShI6iT6JegOYD8IQkJ04v1xs49NmOqOj/qXifXVRnLIss137YdLuQYOOVq5KPBQxqlIAIt
kKGAYmXjYubnoyiCJgGtqiXi9zH1/vkWPyVGU8mbCm45TCwNLxGgfdQ4m+dP0fnYwRH+kg1oNGqQ
YgeQaZ/Xei+LMT99TqkYknRq/LmtBYi0ldUxn0YL7xdi7htEZsSDi1l3t6ihANaN2qiCjDMGL5+/
6H1+pbJ7vIun9g657kfpGY7DAH9SSkMyTo93Xjjy6crV6koqJs8OyXqA3MXEFK4K6NQtI1ztueoC
icZUj7QaE4Nk4aRrue8uJCvJAWg41fbAwrrxH4hETGMxRrneLPqHEM7e2XodGGy/h2t4ZcdwvPdK
0hMV5XUbi6ghnXCEdgP/5XaF9pMZkTFRQelSXyCN8TG3dsxI2dlJY9R+C/ZmLM2xluoPAMwAfYhI
y0efZl/QtD+OK9ADJPHDk8B0SR4RlsB14LC2pEteD9wD8VL+QLBaoaJJqYZ0xSMB/I7ab6kbJrj9
ISocCbHSUMOJsUtIRHj4sOuylSBT4AZh499sxLo8o0+8c+5sx3xaIaF9u+89Gjpsm+DJCIehl9eh
p5fVvI7uJHpr88caDjD3tY7uRxHQzKsnp1FF3fH+nGoTA37X8Gjeicsnktrl4SU/djq2+juzix7t
/C5uw9VoDKm7/v3tYMX4mzf04gPFSwY9UhxxpUaRjtu4eLXmlyzPMjuM34MtL0cHGwvlEI8GqFEH
x5Qo0ttMQNXv/BvxObO/HD3HnwEZSMc174IFau0tABG8XBwbhqO2vUg9aWoAbQ8V+KoqOIDLNAjQ
v+WuE/mClFR7SSZY5lQG91c0nsXOcWFurKzb8rmlLS0HWMA9YpwGEiz3OU4hEd/ERLFiecEAny6C
zbD3Ri9uQfJs61xAY/CXTRCneyaSBVSb9JAd/PxUBivtBqIksYcEeQqri4P86PBVBSr/phzbciWD
UFmeLcYug2K158wmQLNZiaZHZo+SCB/u71TV1Ql43dUNRSSKV/4qxzoVqIsN4CAYpl8gEORaKvwY
6tFxJ051g/GWBYZVjwB6kyM8ZShtfxZlERrZgj3s2hnVw9BnXnJCPUvzzaDd5Bi5nvwuMk2Z1NgP
sT2i8XkOhtBJp+c65a6xuAwLIcwKmlb0ASgv8GXjGupZeU83JvPGgtLvr0Qy9/2ME5qvImsFHMjU
s2E1dGo58EncQ7YFsHycj6MwESD4nbMRxuU80XBmGWW9AZ1YTB2aBUe/7KggR2BGxC74aIM4/1LD
ancFyTLUBRygFHKrEj6EI2j+vqBnHkpS/mjB8gbZxANELop//2b/LUprhlQOO5ILQISoHq0J953t
ZWEbK5tVzYTFh/uZfw60xuCJIwcg2BVAs+RLo5eGWsVVNMqToSLHpnsZGHsy4IO6rJlSB1N13UFy
SCjYA1HiJODTeu8gm4sU0Xq98UpuhCSvDpw2BLzhvTl1wk1uTbRP8GEp1r3DxuVNALHlGzbWHUbf
b18bEokEL9pFPPsswVo2lr3RXte/CdQbrlvEAp9tnEHiQIUdUA6KCSOV9OuqTvo0foB/BZPXlf+0
KLHmTgX8eJCDD+/z/ZM0cf36Qg0pHmCsT3N9dXB8QG1OG/v3hOSyEEUanqkJ5QNdxMDXjSnXwjl3
+Ymc/UcUPH143vAGtrj/E4DPImGN27S+spiKBeCsq1T0MbgzT6JMBmKVZLB1b1waDi/TW2CJpXuX
v2TwPXZDHtESYTeMpuu1tIfF1QPuVZS5DY9C8uaZxk6xNSCfN2w40kJNHsVlPyKHEKlHSkfug5CZ
sdTx5JpG9bL0fyW0dVWMqd9Vg61avu6pZPrWsMu+soI1Q+GiADgJ45igzFDRXCMrAaMN6JNjwJwT
6utqn5vMtor3/egDKLFjbAQacKq7kZ4FhRGewxf6Gw7+wMrk8X2uF9759els+EcL0S3ee4azv1xq
h1VO/lwZeZTz680c4aBjwZBn3MJiWtutYD6eFZhh4mjzuNdvd2j382CSs05QhZStQdl1x2DZpvcM
bvrPnRDVI0wlBYsdzYn8HccljDzdiOfvgRPCJXiFcRrLXv8w0zKQP0id3G+5EVDodh43L0OfbKgr
vGYtiU9lYA54m8ZQdqozSaN3l1eSLmuMxdYFGKEmRhfoyByzc1rPIxZ0Pa9/H7eZjhJmylQEYv2F
i7Rk43zfuZvXJN0aNIIvrOB8E+c5VcF4lzgkBSMXH526B556HIv/rfsSJasjH6rDL8ejA+Q4mEi+
EcAtET85lJgCpvn5anSvGNPDNq9pMjo/TK1jHeUw/tUsDbCquOiVE4vwSfwVhVi7bAkYf6Y/QYm2
EUEHzmELLWXJGgPOtkuQ50yf/pxoZ19TP75tqBGcVBwSbsH5jeUmR70sIkVZGezFOskUoAMd4iLU
o63zforTYxmFQy3uOmZANwVedFB7mq1e/zO/g9dHlMBKAWk4OS7wzdR58D+mnLddzV2iB2htnSXZ
pVHFMG+iRV8KPppm3i1SZZDa7ivDev1wp4Obbz9kTAvwlfiIh1m05jNLcz0k7CktLaaJIrOg80rW
Cj8dHOCoo/i5YBTU8UyShbwhlwqnIoM7dd7JIbpzNHEMIgO/xVIYi6MkTfLnqXopR9h3zLaFh4Kq
TjuY6QzEv8AQfW6c62RilstI/2dTRfBgjx3nxgZKLBZwrfDRM/fw5NZTe201wkt2GjKNC5SVZeIa
rqZs7qrWyYCxEwNS27uG2VP4W/8HhZKe8M/KfxNAZaeHnegrc/eOu8zWMx9Af4piM/+LmF3zrIGa
MsgJuMbGgjb+TpD8WefojgQkiG0pYiXxs0GDcRfHyBRsbCk7ST7DLZQ7WhK7CXmfVQVBPmBjrPNE
ebCtoHFrTiLjsO8aUpu2Wfn3BCxJuDDHVHKnVZa2GtCqBNzA2ORzmcVr+PCkt8evxUf99Yb+MOES
3QconhmQipjqsgnp7B7j9hLgwttzgJY0c9chW7jZOeAa8cewj4mFGZcf6yDAage64KA7+lz2deMF
EJxzYfeWoVHENxekPee/sb1YmYpiBDw10xeuOFCZcMXOqtGIPHlcXGm9yOCgNkgWQQFwjb5te6sg
wknYP6g8FVMGrfS4xcwFa8UCx0qhM/SPOyaxpA6gcIRLs+1gZv4jjLTWdauBFfc05DTkOSNUK/5U
vEHhP3ZmV7e42GKx637PyrIWedJLNlBZdYTLsCV/iM/yoL+b4LJwd0vRHJyz7Sh2Q3r2kVxGZjqx
WerDyUmJqWdi6PShlSWCGxt6IlXki4k7b9OF9ZR93xV6ewAdthjJqVb2t8KgIPVHxal38KAKjb7S
yDvQQzFu4tDOegS8zmMIvk3HIlOqRTRpM+2ZjHygJP7xIpGbM+mm/LOCiS4XYyuON3cpIOfecjW7
rPCLJhQdER0sdwwcu0Kx8v9TFA+umUIaANfYJJabVFSLGDtvlzFAlHlFqtEln2Sd49Np3ToxYD/B
zaJCVrtoKIRxnBypTovYYxl3IwVXM0uJSf2OhECqJvrtzmIx7FcNmnTPa3FaHbOV3BTkcaEiSVvb
kmT4qMyjXyhVvrNkoZcFl1UHgraN4bsOnI16UyxrqEb7l//YsCMs8Jaj38M8cseOVwSlvuJoHzrK
dE1T6b8c9AIAFkGD5Ja6ZoCLuV4/IJvtbMRBypHLXVuuQfJXNqdrRLMbw7NndL4hrtAP8VtZAWrQ
dRd97nkuzeMIMEQ93T7Zy+chtVzJeJqyhMQTfAXkkfX5Wu00ActaO+qXz770K4zx+Tam9dCcLr9t
N1t+FH19FWSH2JCzDbxPafuT0fSaBOFY6F//J2Cd8Kqy4+hMp9SkjRbrFmP9Gh3swtRon32MTaz1
VUYCa31M2LK5nFY6pY2iu8itxE+Bzx1pYzbGgCQrswQuqCrxb50GJ9tL2GOL+UIkykODZ3abEbyN
TlOZ6ozvSBGxp85btNk2MbQyl7pR/VMiKqWSX5r6t2HJHDaELDPPugnu62U8Xd1EyUlvrUoihWOa
xZijaaHOBcd/BdsXshWEZ1mceAlUZ16lK0p0UOukdltWWozuYUwL29nEAGm9Sk+BpprsTj66ct8l
haP4A9JZ2XUSIquPURtvZcqH5p8ot730BXPsC+XkTk8w0AP5XyWB5h0YWo4s9LgkYOvMe8vM3pea
V9eKTJJRCTsPuDJF0XgyB3P+f+H2WEQApqgKoNMh/XtMbzlW5s5WRY6TbNg6ZQImEG/eFSxYQrPi
MZCYN8K4/zDpbQBv06PGjm+PV+sONpqrGKVQzsOJ7Qa5lubGnyPEcwzya5uV6Mf/TOGE1qZzGN/Y
zCF/QdeD5CTq4HvszlzQVxNZ9XU1DZlB111XVjqD2aofkdUloiQYt5tBgWiSkFxoWOk0vI74R8WX
WHtj4C/s6HsTfnn/UbEu9dptRNf1qTpltHak8/imdx+109fkJH4vncu4RYc4cbDFxArUljffhTlm
j4959wjuyJUaacJq/1D+Tl5K95kPCKJpl8EPcDiqcEtU/C0NzZWpLaWJFZHZYXdopKVxsfEh2xLu
h9Ea9lLl8ibPPAfRLeqfq1Qvkv6EL+xLeD2jtoq38V0lkfEpttsO/Uk25mhXHCWHr1OVmze7Mxec
Vffu8rYjD0y/WriQw2cRooZOo+5twSGuVNnlK4LhUaq8m5DajSd67o/FyqvmFr51GgGNUhTmaRep
1/SnxHMX22IQdvJv+XhG69JGt4aFATQpARpCA2ig7uWgs+eiwU73lbNrf9Kp1dtlyuoO1dayp6Z1
dS+JV6+K6OvhNstqlmrU2PC+4XNuqdgeYYHw98h/kFvxZHAsNzuUgvXnX68Tcu5E23CcVRodJc3f
rmB03sxedFHVUVxnTf6T94MqFgEZGFvsod294y4hCHVT/++HLP4mqgpRuzgaJ6XNIJcziU3EGhu1
9uqaMT0F3rAKbjicR0UJdzgJ3pds7Bw1W+kLPsf1QtUODCKp7CvZDpSY1vlDRUxxOGA/4S6hXKhF
cP9K3RJO9TIikDyNrV8u36D5Vxoh3apirc5o++DRr88fKc+oml/wvNjGO1Hj/IZz6G/04YcM1RPj
vV6z0+PARdQLhq9I8IMTuhiWRHLgbO9DouF7EkatAc49QDDEAGVXJaQ6D7DOzaoKlcnDYTIyod1u
pR+kEP7o0+GvyF9Zt3wRScAlrFAz+ynQ4nKUrPs23Rcrhu5zTm7qezPDXYaAmbj1bv+B52q74HnS
7pUSVbY7nZ89EafmfSeeClDROEYwErgbOGSrWjxZtMXhiuXdcthj1uDhM2sxzMs88PR1P156x6y6
5diOp5IVfufLZOzBTGVWl6mLA3t/NHQyRs1ddTFfoyVEteX+ZlFnmy558iZhFgsB28hsiwo8ce+C
sPRGyyP753Aq8jM0/9peOCdVnwNZ8OMW8URZ3aVJ3W7Df3IqYG2IAu5hqdvWEPoiFLeBYYfwk64S
gB/D8N6dAXPvtsasSGyGUU2WHecpC0UQykdUk3rZ8+cTC9H4G6hM6LiPrvw1L2m58jUwke0ILhGB
nIXqJRmWxaPYVDhAq32jvJ99QVNVCKljx+JTHUTLviTa/KuNFXUzpRlwvT1AKQ8+/kU1Cu2M2bz5
QJHgR5X1pCmYWUm5fnhQQNP6toc/pDDmHUTWsnHZ2IRql5ZGOLlS/XAnoXe5CY1WG069scKUWwbg
sk23Anf/HtRFiwsbsAYTgXQHrrzKbCtdamMenP4AUci23caLHhvPZE/qx7bq2V2LQBpHw60RJptS
vn6tULE2y/qF4F7YrGGDV8aV9V4tEQGwpJjgXyTxdtal+ASqw2gH2ZAZesuNeHWkbIyAibnt36nr
FUN8J29ZUzqL32la+jzLNnHzyhg1xM/qyuGSDvK24Py95bpYTA93GfMZfMWHneusSdBVcWnt4qtW
q3o6bfVTMt0LrtQz2DIIUqwdjff75O79GAa+3JTkWouQofVR4OwtzwM8zj9WdDRecedgHkt6dANF
49keWLoDy0TvhXdAjR8mhZF7d4farnO5bhy23+lvKTGh1rT9Srcb4DXDGuBvW78kIvWutggOVKOw
YNuXPT7snx4Tas/+eQlgKZsuSIzFVVUHocUpzRS5q3N3wrNeIk9W7OBqLXdachf9ufAqroN5pCCZ
85lBp/h6fHem0h7JlZFS7Wno3MZ5bh7JbKiETI/K1m8LB7DWIi7o+eZseP/YYyhNqIKv8QRFJzBc
maLiciv1HJZORM8ZU6mhfXP54Cpcd/trb+M7P49YBcHYvinFXjsIdrkOFrGtZSoVAHVFXiliymHE
lAco1vE+BHWWGlDte3TITsN/cF/mTwOe6ytJQl7RTxnNYRptTH4LuzhIVEMdham1FC32d2wwxFYP
KOiSlOLES96Y88olgKtbnf6lQ/o+YsXLN+4kfGbTWdHFUPOlfuIuWCiRSCLA0bj8wDWJlb+WJ/WN
7OEDQIqAyF0VmDReJZBlr5+uZsjMsGqB3zHQAeqPnGtNkrYDO96noUhAHaifbzLrrcUALNLtMAiI
wj/2k4wQAr5vvKD3ezgTMETu38Rg6/LjG0yHwWfGYuFzCAQLivomd33yiNMsHwPMi/2n24yJvifH
XwMvc9YAODo6v8Rz6VMOTEnBw8hl3snm2/hzhuJIKXe51l/If3xPX3KAo61PayczE/KJop6uo6Yp
VcntW64S7yiaUhGGyDkk0kWJoox6S+89MRajUjP9EKG7DLmI+kAjGd2y+/+rg5Up2gFlejDUafcD
fFZV3xN5U8X+cf23tZnoaFe9yCw3BqK+aCO7ZIhnqiVO5MkMmnpY/ldTpTgC6qXyHnPqGePuNyoh
7/x03hFtdVQ0x57crarY+KQuPutpQHeIT/zk3bbp0NtRYaZSrBFQkBNHsvJL2sJwvpFNfKgjWb9k
0N2QyclqpBe3qV7LdYVAUtyVEiKUZkhq9DQV+D/dfJoa2UaYo752eFS2GyDXvF5jRu7LWCmzNe55
fkoJ+KuUOW6Rmpe+p0rQeI0VTX6b9wZHC5GllnQTn0cDJbfWALtLy0Fz8Z+lAaeKdvyAEBsF94OS
wEMsg+yjRuMoMi+/swAVaYzmUHCz8WiF2naWYUDXUUNWXoqt4U5lfhsu3Q+d+DGWdTsZ2pNi7x36
NrFM+5hnbzkdabePd0KerJvdbVtG7kditdd1NkbQRVz/ApOEJFv3NEHlKFw41qr3ODtHLNIlpXWn
8ZsN7D/KiLmqjshBnwCQBktHYpo2H55cHOPQ3cBW4BEqMPPSQxjzpBvLAvNIMttdJ93pBBY+iBx9
HbDmWuYJUBBRW7XMj5ooquVVbM1rQLgwLpabvSGIddQoiSjerm1pBA2f99CDB05OZq/Z+JMQVPkR
uqV2T0ygC9xoGuRYlTnX6Q0VZU1AHuv6B+/msIFHZUpAIWQzdW3f8oGr3Lb6sDDHfv7cHR+zfgEx
sj+NxJg6//uZYLY2tI/1OgT6nk2D0eJ3QwA9cklGHS965k6zI/ToUrY7ycTa7EynXeJe2h+Fg3Ax
vUS3BTLu1jGhzdC9ygLOFyC1CJ9+WrJXSbrV93IOW2KnTuOCLn+bsX2avu18BxS2twVEeaqn0w/P
8zvW4XlPJbT/aZNznyZb0Oi+Br5Oznfo3lMlierFUFYPzzhPtfKKykRvnB2el0MX/lMlVwOPr/O+
Jh4ykREQih0NP6AVM5CEq/T/RED0bORd1mp+u2Opo9qhARLK36Q53jFWlVQCoSQ2il32zN+IL7CL
Bi+3JxLaJlaSgXf+vMNBQIbBZEelEMkHyuziERyPetd1sQFSYZr6BPYYL4T5Z3mjWKbTW7I7TpX9
0wV1hWDuuSkNsC+rdgWdZ/PYKsJbe2B5+Ar8fqBCh48n6MAyDDV4t7RJmQeJrTRj9Vr19LSvGYgz
pJnqcPO+J7+u87pyMoa8MofuhlZsw3gge5j1y+hvvrj1/kvDSVWa4K+LpgODaRjR5YpM8FkpW+nr
jyfT0J4a9i/YFYkHZykzzew9fq0a4FcFpBD1vdo3MY9N8PE2CIn7VWKmeKd3iqSEVhzYKBMWcw0l
mYnRKNghUWRq46BL8879e7QWq6UOe8UanjOlzKOTTwlIPWg5znWj2a1U7DstDMcWpQXZjJbtnaT+
WaAeSdg7XxweEN+eQy8Vm2+UpfQyFbvDJImVMrlzqpTBG4rvOMbefqm4d7ORItXaHczpxgKdx/i5
G/PGLQn0vF5awnpvzwkNjJqmZYu045lX/oKMQONDvzZ0hEUhpPNSHdzO0ouqo8J5Ym1825W/f3y0
6GjVrZyXaKHGAme4n2UgC3BsuZa+LFHdVdSfxp6Tc3gWsgmlueOx8AQM4YJbfOXfmt2HwY8ZFnGt
GMgcCWufKUY5wkO5rEjlCzAFtC1liOccHfup+wVWkTss/Uoo4GIl3XYTy0DXysSRlLPoTPll6Exd
dI61Bv+nMEFWvgYarrTvkvkHN1NfPNapjcP3q6v0wWrWjV+G5wJUj2eFSNQCSeYHJeje4lEf0wM6
myXC5Ee+je3qkHoCEq3Ej65biyjrLhvH6u6OkDhKlzidLJX9spCaYUe4aQNQ50Rms+RGTlEPfOpy
UU+cu+BNlEeDyTeN1gPRYZxan7VORjpbcWCDQe5R/XeBB8GayT0nQ57z5T8bu1Ox3e1cyMM30dGm
WpvWeghqs0FwiEdTltIAe8CirOLjoKFSrrJllZ2mng1tNuI9eb5oq1otApw27CpM03akJSZDSf4r
Zt240CRtSIVc3ygD0FWOw4QhVTIS2+3xZgQD3ISGuM+MTTSE7DzBu7LMdeyP3abQ1r9kSz0y3O1v
VQHXkyzBWDXIvaUQB1T5KHENLqZJYPuoRBLjMK5CgqlfoUlXbM+OzHYqn3myJR48NzEV5Y+92vmh
ZeR0GKybgUsQ9tNiir/5S64GRUUTazA37Spb85Su07xtdej+rQb9eLkyWrpPimCrrHevZ+LK9UCE
g7ikvUDq93aNXUOujvL84GLwuGbN2wBqQ7mu4aT0XJHPFLdiunA0pDTqYutOMK2MFlnqM2e0Spkw
jH1vbOoD2QNGQIoSq+k8GSo0bnIH2wd3sw3U0O80OMRPnc2TZWWyOpV4nc73ieaa3mn8jdAio7f4
NBnMDjoDyNfZ5htmTXOZHBFfb7yt6X0bjEQQf47UCdwICmJ6DRvkW5bVReKRAhW15geet+gwnBmt
XAjQtOY2EpbE1OZ+oSFOLzYLlsE5E0trMGb9J/6Qki2kongaaiE0KFxNpVbchcDIDhvmNEHlzo/C
Iink08ldtl/EAHOisVVAjXV74+jsqt0r4e7fnprfvaBNIuqgEtmMJsdjUqnSMfaGjeAp/Uk8BIfF
L3wh1sBct2+s5ZZKCT5K1ItTovkuFYdV2cx1UX3gbxIgzl6E/89wU8AiK0xYxHGY5TZSGDcQiLhI
ORZ4Sxrds3pzzse8nz7CZ+vNxSmmnE4DFqPkxmTLEA6UQ2yxyb4RVlAuthullMQ7fBRvJTfhMnDu
PHhJNDGPC/CB8X+SVx32HqSTWykievMEHyYdKNEJ8eWk/IP9oP+uIF6/S02e3R/PMrYxcMCZY0cP
lxu3mZ8MKhqG5qQovEpFtUZnuBappKGHgAcqlDNZrMjF40ne0/q01padORvOqJmGAaEWDmFSor2F
RZONlLj5Ma0qFJk1oT5eLJK0b8NW0gyaQu1G8QpENzNWI4FlfpMYkV6wR7Urv4orMQUDVDdx+VKc
YS/BcExU+nJCpXEP8DsxUQdOipYtS3Rp3FCjYwwkryYbtaj92nd7btHJYjRG7zlgcW5QvYQ/HH3k
RGjTjAQ6UqP2cy1W4QcxQPd9vaFwrPxWw8rHTdLZH7MG6Zc3MoNzFdPEvY1kikA6PGjXquiiTvOW
8Iwbyti5B91PY6b9ezQiO07oc/h1nhAlqwwPosmZ58LNG0P18lH/M0rhLYvcu52cWWa659MRIHW4
LajuVNyNklxRiMvxXcIeMusH+gjXk6WL/s0LxH7VwYfXJ4CGOoO5FzYNfGWwdSufG+xNAtREgQ+i
Wn+ABE4YQgB8t3PLeXUptAP3CWnnhptikjp8JMfHkrgJjqXb9vBH+xzqdlWpKHFDArCKSzDCTeJg
bYkp5CyQYZT4PpmOpmdhKEM/LD5zPMeE4Xib+fWw6I2IYP4DZQcCWHsmrs+LMnnfb8R1xygjOzyY
av1YYorh/GK/hBw3vHwM3f1HUI5VqUwoemVxJ/Dne95oTMJJsfXtB0phhghYfr427k/dqe5s5dYu
DK4crd6Yf8Wkd6Epz+VCLTbCT41hZ0CFOBwv5yDMlj3CzOTKQbV8NghONkkStzAb6EmqHqxlHMf4
Trd9dLfpxAPEdZwUgLlgeLzP1XOq4aRoWm9i3z0KxGQdNK/eCmF8U5YtCGDJXhb4EDEKR6JNkM2P
9PIBaLz6w6gqpi6P5bkOs80dr0pUWshMsz/0eErHsYejmy6Kzx51WGfr9FW7+AmekWi1hOzW8MTp
cIzsTx7sNa3wmkLqOsL+nqnSaIZP/eTnD+pp3VKZcfxfhmT0L1nOhtWSSY4MoBFSRv7oapzTQy1B
yqDHy1HZNx8tk52pJegm9uEq/p3floA4KNYYAyFRqEiaHxEdekQn9UMmLBcf4dDUvwzfLRZROz2h
VtzWbzu11Kv9fGfSsnglpmBbba+o2TB87IdUEuSOFPKHhb7sGtz0/Kv0rwCA+1JcV/XGU8bLioik
MlEEOcpjS7p0r+pY+o0YNhdiX6l2N3kcKQn3AcBCT67BmQ84v0TXPlc2RdrhHAcEtTe2Z1QP2Olu
njZ8cKgVZJO21R5mJoA+8dI0H+1H16fBdjLXADBgAUxPWB4AK7OTWVHi6E+xXiAd0lBb49u+delB
1Rnrz9ThWPwC9AIZYvdpMuKzHbKuWEy/Kkhd4jSC1Q+fNqpFju8NzFKRkJF9r5CdZp0LM5LJq+BU
d86o9VzzlByBoL2Bjlo9qHmE/HZKpNAmFg6I/cJjIOjEzgrn0qWO6YgCLJePSr/Op7Xoevbv+xKX
DHyHrAscTbiaeUbhS83WyVYZqUC4vkPxmNs+v692gzx/+jc3HSoYLwIkkKvY07JK5crmoU80Pc7e
6YAibC8awU91dpD5HQ4Fvj30Q5Gjt8rPxO9F+twc0eUyKEIKoB58ydfvtB5UKh9vJpKAxgRkC19l
Gqtdf759sC0W7Bu43iZxFcF4ss08nh1cewUjqsbim4QWDXLFpy3qbJFEdIA6si6F/VXIhJi4G3At
rh4uR5VbjG3ncI+Yan5tK7Ob9dGbnEUsSS4gc6t3rhk/0yZfLhJBu7WGgTscnlVg3BdP9OFHNFO0
rVq0tn/jGax4sveQZbGKpX8VRqaCW56YxOB/dH9+eW3DZYwf6Ki2uez5nesap5+ls6QzmeL6/APU
5+qYdBDwIK0wS0Mode5IPX1ZW6O0DKc5FvIKLureB2yYA1LK40J4bYgAEhgxJbIV7/VPieKNSnXf
kOgFoif3DOvPDURG4OIZ7QRkoNWQfBmkFrYBhBWpT8+s9+W/7gkqLZvCJw9QUngX3T0BgmhAxBsP
n1xDHvbPwP75vDf2PrLUPZVyemb932lAawsANCyYNa07doE2Ey6RgprH0SWfcdTj7fnk/5Dhokbc
JNXl31aMdFKkOYdhvKCjp29mMp8G3jyVgzgFUE597tGwFSq5GNrxfrqNCCSHPAZGs2cTA3HwuxU4
4FxINQRQXgBGTKsURdMGX7Nug9YdSbYJ6hAp+7Uki7Qjw5OXnqvpghf3Zjl39UAxpOVhvc4JSrmD
WXY0UlXJ3c17dwG3mQhkU5bIn29OlomPioppLlooA78Bs2FmTHUA0+phVgf6mFbgFM23UUc/xBln
WPUX4skyVEItXIv2s6yRCDlNy3tEDlquHGZTto+2fCp0KvxmfbIqdCL2w1J6/sHNAwcWuPjGQm+/
r8TIkbAG6ZY4GeMpfQNA90hr3ytImaQO09eNYJzx4sK8po5sRuqToekoH0Sq+FUAa/JH4+MoiqwO
AIP34pJX5rqGFSM/0SEfDGNpuLd66FjDUHp7MtXRf2MoFRMccpYUduc40JsLZCJzigH1YcWNAxLP
+6qQLp5XpuvzhHQK7rAvFcYJGMDvZYnfFMwU/JWJuppjxk0hdcZauelIs1tFAkuiHsPyjMmcP65n
2bfNet7q8Y8bZJaKiAO8LKfauwkyir35J1MO7ruKMWutrNykZvw2bJivpklAsc0/2RxDYficnksp
rBr3QS7opGsO6LKmOvr6LXbuNUhHrupqGePiMw+TAfuuxsp3arOq+fS7y/zqwHwnhxAOpv4AfDTR
Kk752bVDl6Dv7ckFn1AAVxfjCLgANaJ7OztRLJHpfGDgg5p54AY/CHRCa6hNQo9k/ak/hJqK8NkH
PAzr4x81y5bNNaMrrp0xHc4xn7jvR4EeS/+h5ioDDyNX18DDQnuOsiW3KLkhotlyQI9BoqnGD448
NLJ9GipzWlb3eTquwXxTZPa8KvGSCDIeshok0+p7t/N+Ra9q5KFivKx5v+00QDuWV1sQp5R86WrP
DBsLk4WZkLmpmdI5mo65YGtJHyCrHx3lk4MG80qrGa+OD2IR5RpHDCwm+VWWBPuE05DYpmrv3zC+
9iv9uA/Qlzoads+v5UB6kGJVLQkgpgh+NTaIr3ez7rLEet5wYqUWPr7YdZBX8fqiStQba9DosKju
/ZfxUpXBBN1aV6W6ABDYSbho3QYGYlejLX2QUhPhjqbC62vTY/V2bYd1K1OVEMYs/RAnFl5AGq5i
L+oa6nFyH1Sn4aHAtIF9Em5AVljvXJmXcXNKZRlhfj8f5KTpnVr0q5wZTcHoObRDVbuiP7nEpOZP
hFA8xldKO5vq2AMlxVKlZk2qDC7v3KjbJtmTN+90mgEybkQIfehFPXKDEZZFYpcYoxvavnYpVboA
vnP6U1li05VgI+CxNTgo9iJD6ycusiaumlHtvKVG1EbKDdykA2Ra0xNPlM4i3x2IlUQ+OFBjI6i/
1dAYuwxeJAUXOA09ykycjGK7LqX2WKD3MKqe2F1DpVzZbiCbZXGG8/C7uGWb5K8ddDAxrE3PkZGw
dtt8Adsn3SCNgkZfgz6R5pk1gSIgf/xHt69yXqp47TH2k3BTtiISIjMTVvgn/SoxiIs1FIyJO2mt
QtZwJPSLZjA1CrIxR6Q3wXa5ictUZ/fdkS62Sl5aeoR0Erg/8b1XGCkuh9CvGwLtzPKo+3hfGDtP
8mzE58/tEbn0Prx8ouwokKp23EpsLGpWV2Axbj0kKBpbwCz6o87h+Gmi4ZXqw7J9WxwU7X8Ii1Rw
L7rJK989lrMCD+p7piAqLdmChRkBrNyYBh1zFWX/6wxTCQlF087y0TNp/goeV1EOFJf9ct58Ssf2
mjnJAt32NW/1+VRuCvbomcrlM8lpyyTsvTAfytaGpIqJlD+H8XE3C2zQSV54jvboOXzXCMbQmMWn
R0Ett1AHHbjvIPKMkAKTBYBZMQqwPBtGBafT16ma7QyvWdHyqLkoMCD0AOSn+4NtWo+RylqrzXMs
wy+jzi89kAGgL6gHSmUh3kRrMI/r9PyxH0yRUzCOXq/OniS7oUpkncpX/RwXh3rurI+aUd6pfEaW
fhVnMqhMvsIuphW6iKiEnki71VuQOboz/iipRz+4J1afrlLdS1YkLSA9e3x2RX7YbDHkwBv5UqkN
PRI42awORm7U9buLFuH+D/ZrrnKa+AlTHKI/mYvdXeMa68l6DKfipQZO78fOcCaFFfZwssGfoxgW
5p1/a0gzf3EtSjSsg27tgqHkR8In5xe45S3Op68Nwwkyiup4QTzvMfJlX85hMuY5p1kRmHw8T5KR
dtR5iBgVqjTL51Az8f3eYv+Ycr+6NlCubEUh05HAA2s8R/qK6dbY63Ied+xYPrvWdRev0l15z6Hz
uIQi+QoCS6XbJ+6u3I4a0ZgRM2vrHzD8EwV0nua1Qc5uRnYWTlg0Fs7MbdekOQgA6yNoRx/k4Pzz
0qemX7MDaOC0SvQOrNnLFIcQ34XQlSKoTcwmkBSgdokBvh74u4xcvwIBPiz9SCAFQneuUWj1ZNpW
vk7urTQ+4EwGgmySKWzpr+SpUFgVe/bfjlJ5tG0EjAz04IdTmkv71VTf7N56KFFdD2s2w3pHFNLq
pRL3UKtwO62EX9LYoZjVWrbGKzNGsP57Oj13R8FSkXl+Dy+GDe+/cO6dnSXz9zdin+WzH3+Vw4t3
mBWxqX9+beGREm4jZPKdTm8R1DVT9wnarpC9pFsCTL/9RRkduODGB22m+cGn+oOVAAI8EbqL0pR6
qAD+Ua4GSX/QWrzBR8m+OuqUItaWWqbKzlI3uACI0q6zC7C7OpZwrGDNiXEpapC9kxP2vuoYxpQK
UB44qD/Mtmp4/eFMfDb8pcOrs+6MQg1zn8wFebHAuJXmG5PStYHOF5c54kVVIzcC/xel2qF4Sjrc
8QQd3KKffW0IcPTFH6riT+aHgkqWxxnjoWw8b6elPAJHm2RqdHbinUS+hwKG3CbtbwEPoT1scTyV
PPSvscMBaX0KfMOSM73vo16G6qpkSN8t+Eua5kAW00F5rG8L+PhHf634vM9ttxtGiwaQDN2SRWXq
irhHMipGYeBjUnrEHDVAy24xMzId+/r+8YS9Vq3j/Sp0RpSC3dkMCjSpX7uepDRmQTiCGqgstAgY
eifvQfbIEpItWR6ZvbxiKKrfK0u0uzMphAGrgZ1BtX9nXVb9wlC/57kqlsV/mnREaZ3lZ4kuDqaJ
zESIDd7XGt26/2rUlWjfve462UaEEbV8BOyoRGaLVSfobB1bUxP5177gfcL9hFP/0/sexNlFFYTf
Mw8AkB7/Cc/yzN23zy5a3XTPrSv1Ic0GEi0ov9pbUnU1rWfAKXwKOmsyWychzGj8AfCBb3AhkZFU
njQFFV+gmPJWbMFbnxjQgg7K2TdVIhkpyXRaqi9tZTS72l1vWCAT8wc/dTqK2EO2MczaMzC9P+gp
aAbKkdD2Tt82GsL1oruUX8S4oB8qb5+59hywlY0SfY4IMNCcwr0doHJTT96EW2OEP975bMe2tAWe
HsWpEYASBs7qNK9oiJfklPsDJwYrE5nJuKvhof+6nFg+pBngLQMRCaMyA3f3N7dod/tukEsmT6Z0
L0ovRhDZVkY+nfNCr8Rs+QeYXsfRm9iOrLXp1elG38EbOaJQvxAV393KekQ4gY7Vv5Zx6GErxhmh
OvSxnXU2o8iStjiJUXsCfUdzTBjonut1olMI9WkFy774b1etB0/7dP9+6hl6RWsYoM7L08ApaORr
LYXwKrvSz8acb3EtxHowjOYBPjGqw+FilJX0RDK4pJcDxe3GLitTokyUudALSq73QC3Ei4YQBuGW
R95dR+UJi2Im+FsifExn5bILgXDepm8Qqh2oYG21dQPQNwdQPpfBcLuy1mOsru4D8pOR3MCUi3le
BtzxwmpMCZv1n4q6thvZuBEEXMtxUuXvZE1zTWxmV2iH1hak+3d21igStqIKh2PXmAd5txKyk0HN
yWv3O5kK2gpMx0DmH5NraBPcynzu7Q/RXS7xt5SFpePXhEf7XYGngCGieSKfqtbgVY11QFiegjK0
sPmbgkbXxAnQ2/QDcUO6mPWTMxzxeuhC6+A7U6guh2JUfdj4SvZlk147HjGRHGy63bNC59eq7vKX
FGQx0ThZmIVYsUF5oY1nwWWIRBFGZ3lM/d8FOtyo2ZdREk3KsnVsV1ijVZFYnF9E8FYL5w3cxyvT
N+j1NHu0G/tRKEZdkD08jBYfARkQgn5yukDxNSPCOzDovFqwEDpywjcvfoxC6O4b5AhTCEDbH85b
shNqkyl9xfIbeyfRHV/6daZ3mSVMBXCXmPryhorgsVvljSFpmXy7xM+8l7O2f2V76jIQUVe/r8VM
a/4QChBtTjB0zZyN21K8iNNXBgEDVWCaSw6S0gHqhUUEWSf4gcYBXX85SIqEAmbAtdC4h42/q8LH
/guZ9RYyc3NuG5+znq3F/HtDMpTfK1oFxCd3g5BWw7a7oWZEJa7EC5OdntU1ULKFHXe4NFz3ETBO
OdctP1yjGzefYdEYmT2FpvV1Z0DnqXIABuUgcZm01G94hNVSbacR+/McUOwgMwnTFFVCzCNoAOwp
6frVlDBIfvqwhxtzFmM0/GgkOygTfqzyqDsaFsCtG0X6NPYS2DJqPnLZyWMG5wz/nwgAhKne0WXr
X2UizW8rstKhdmoM3zCYJNL0ZNar5OCr7WF/OTY56e38MjVycolSvxjNYT5OX+IXxw2T7aQB5EUy
arWbbsUYS914AQCZbfzGzHjXPmiQCfW30QuNDsO2RZW7Ve3NTkEcI3JOGz7TCeM3P6qHcyncinxJ
ThcJdIFHTxbM932sGGhHj9CmiK5UiAoJYJz3GIddz+fDJbbQsVF0eEI+G+oHMzdA30yHj3nGL7sQ
UDXFPDTMjEIFvGfB5tkCA0fWI/v7urPXE0JRQLlPKWYRwDbozv5pLomoaoj4pAQ9KFh+Rcfrr731
umozQItCvrIgflJFS4ujQAzYncmHI0G96Atrup0AMWzL1WpZ9oQ7gPuvIUV7RCvziA887fYAYrOU
fNyBJ8uDMvVcsRRSSdE0xqEoS9Q/SKC7fnC3uMoo6+Waje0E+F7/R40ab28B9ffKgKuaNRHXOJ+b
+xVnpG94j/0igjcZhgxksvoaF81VyD0mnXHH0y+yenVqHYLTjUDSy5QQKo9v0C70sfznPnKtU8WE
sihqmxMjsEPeAY94DSn0tlA6sNiNY/jWdOtmW9bdkN3KDRDNoENFIUboTwgsfZ6B3+zLR+iPVbOk
LtM/qCfNd6iYB/ACFbiq8IPHzNpB38G84GvEVBEi+OVRlXgTJu3mLYqd/9L1/xYMe/PIpYocEZ0D
M0xI/5azG9Ix+xbAfg+yA0mcEvb8t+LujgpGAciOk4YLNOB3m9C2OIp9x71IBOlvl1M00YPaMlWZ
ragDSTalQJ+B23If48d+94BA3oj80y7Pncc8RMEJMgU/19//FH2dpXD4QnDpOQ8WcHxGkp6PtGSt
BmBTyfz4IMWwnB77ROx/8+bfms1XPeVjacVQuZhWb1RpyvWProvcuHTo3iDWy3ntoTDxe8lo+geV
I+lPDXsCsAou329PHB1NeAjLMyLH68i5U25vlH1f3lo8xLFwgPmlX5sQDM0r+ety3s9kom56Bga4
SGiglSeNGFjpeQMghxZYlmfkShpsS6hI33ONJyGGKJ7NDd+aWshKOzN+yIjvmRvZ49AiclkjrJNV
Zoq6XTpvwYjbhUfsBImqk+I68SB0sHg9FndFdYgic+oapE8PSd570BcXNAhDQapB0wBm59F5nGte
jpbYo5bqS7QlVndCmne3zIrvhvQEWPXyiMDPm3ExW+KR3VvRlV136D7Z/2n6uUD6cWsDVeD8CChU
NTBuckWKtMcHL136o4EQLT3EhtCGnnHu+1eeUbqI+e5QlpWbfla405ao8igGb5ikom+q4+Km0Yp6
WF34uU74eMgiYWKbabSSdF6pCwS/544XHPUcrROKQq7olhNg8ygQn//qvc6+crp6Bk7gpO1rPaoV
GUYwIZdAid+vpCdDDjDPgA3NwuOzs6mPBdd7uM9z5Akpf/tLHB0losueJzA3OapsgwTeEScEYvwi
tRSifcw1vXAQJ7+6FKJCVVmPHDKPQ9t+pp17jQ5jRNgVi8upE/eYK4xT+nSVoFJDPZqMJ+eCTAkC
ma5C3yoc54wjEUXtuBGgKl271ocOPgJ4xo7AotDAf1ZpoqbTjBo8LMUQEIMK6JppucGDEs3sAaKu
c7nLJBmm9kM86VDlglVzVuOqFGTsuzuMdCa/b+w81gAqpNCDXGG7Psn+aNZMwLMUldDGKIKP+Rdd
XKOROwlV12mrjdKNChdlHtWZeCnwfKBfmIvrEvEqlvfKig4ET+d3kIZGgkTASmjPJPcRakb2x8QC
sqfmI5cabzIqdGfpdfPKeDLAWo+/UsICYWs3esGu8N//g+ndkxGYw4hBmdt7q8Fv44jI7XHtJYwM
x6FYS2u09nGQtlsj/doD6XWbvD0XaIAWfBn+IUlPA5moNqgvq+mdNtPQOuSSp4WoWfvjKputle4S
Uvy72A4i9NebbyioRjtEBooYDWQkHEupgfXvFCoIiN7KlLdPNMxMKSAAnT5f6rR2SdYjg8KeLktI
Ep32Cmqm5yKYagBlGEBSKXRkUNW2qfqP/4wi9lsJov+pp9cK/OHs2hiOoNaI1xN7v6RlzAs5/MGL
QQ628Elj157gYCv2hFwLMMhsMEd6o7KLAIjK5HV9ITqWxh9fddoz92HK/A0Y0HpFHeWJsKQjukoi
NN+R19zpcpCSsEYI6DvrDdkdbNE3/zEFc0SLYs/M4Ua0eFbG0CeoergEa1ePtdzw+lzMVpgUncAG
dLiSvnAitdEu+cOJ/pu0yMbkAqCz7zIPdZmDfSRArmixCNwJ7MoikTvvPXjv8UYgXQEXlYfpMZXA
2kiccN1z+YfpsqrtIFN9qU3YrWll2JvTzJc86NfypbncRaTeO8xvJ46eUhwu4wdpPOzSzewvQnVr
x2WEHO0jD9UZ4UPHRIKseL7EH2zW3r52hiRMSLJUT9pwVKNounwsUzuxRRMMZ4LoZ9krPFlviou3
U1u7y3zp4RBVJg1CedThuWaFRvXnkgTpUl/HoMArQbPhqOU1Wkp+Yldm+5aT2DhB1QfxEoc+y9aE
1M55elrGABkAz5qQhnxv3GvNmK48CEJd2k3XEo4u3oYnysMMjcVnOh9IVc0fBSKD0dxNQnJGfNHa
STxzOhxOz4VN3rx7ZEHVMPNcEVjD7akqQrKEZ3rs9vQoTif6aCsI2eZ42HqbNzFaEKqrHru759OJ
5VWndvSBni2bMj6oYD8LEjlz3wIclj/k2L0R00R+y61Xhpv+hIez16RcJio3eELWu2Z/BbMAZ/8C
gbB71l8Jczmrv7sNUmBzbTFAf0AJIfZCU+FN+dYf/3jXDfr0VYlBMe8gq9OgV13hyr453KrmA6Oc
y03eRm6ANzwsZzJxLgelVpH8YMrnhm+/O5DxEj0qssMJ53hvL44JugfzgBO7JfDnirEBz/2hDoq2
llR4b4f7u390nq6XZ7QRC2asgITYSqSNd6XZzo06zjU7Op+AMG/XGDOzYMc4j1utoX8tJmKkDtfy
tVtfvSjNeCOgls/Q+NmSnCJFlYOh2mnwmXueBl2+TdUwKQsUbE5SfpjuVZkJb1mBCaZa+qzglUnk
jZq9KPhn2bvgS51c8SZ69Qh6JWhdmCea12gDBeNQrlCCFa6OsXA0dPbBDxfQuVkdgc4ic9lrzLyR
IygmP2BpApLl0Ydzmagnxph9c2G1xvmytlUAPlUa06LBUOV9vfqCdG84RltAcWvWJUFy4G2r1i4c
dxLtWgMyOahcC7yotrsNkB7rkXB/EjoWwU2zGjIWSUMUgcAtwLQI1RAXq4ckI2Ag3Z+ahqzMDjJu
9KX0grYURUaoJ0tfjFPKVfqcAaeTxjtNtDwKKLm48MxjVF64ES9ls3ZPy1nDtUfW45HVnoxB4jPQ
0OcKasnxMZ32pC/M9dinV23Iib6hCneIYhz7Swhy0Q/7MCXc5CzAn5W/JFyGFDLOagmAuEVpYjWh
R4GT4/qFgTK19MK2piXJ9e+g5azpu1jREbfAVWGbLSY9HMVLNGADXjZrrOB87H8vcnFChlBd8jgY
6HyaWNKYDgA5Wl93nEQuqfZ7aWQ7h5bDuWUeyXzVvK2A/nw1H1909FrTA7RLza2LMO1mvUcUMosj
Gh2mD3jezNSdeOdIfVHefiJYz/Xsmf5KJgxO0+yxR8HLt1IFpwXsZsuPHG9rcjC86M4ZHfO+QqD2
THB2jUYmQJPy5Zs1ZmW63YWtGISK2aaqjyranOc1XzAEfyTwZDTmqtjIxoRgeoXlKVY5QkAaPXgo
42zv/dypngUDC2Gp5EHhaYG4QwyFt8Uxpw5JiSU5H80FLoRHkoJbzUMSq3mRzN5kfnI5BYyaJ75J
W4DO/IBK7xiEhxRNnqR4pGO6Tpjl5IWqqMKja+pfe3xF4ADe0htwrzxsd8GB6uuSk+J7s3aK7weg
w/yJQhHKJq3zuBms6/SrJt9Ysu7kpVED6UAaUoPf81Wp8MijQWo/34+IIbtzMGNC3uxiwBDzMu0c
F32602vEXT44fklaES989ZnOOCoW20w00jV4vyy/fwxi4v7SfTjdvPqloCQyfkmA16piSCnGCzN0
1RUm7aDZueiGsWy5XmJuB3TYAKLHMrBiXQfZ/CH578tGyh8ysM+WCydzNY5En9N+103axsTfp7UX
/pACIGjdawGQGSPhNDXEOf5K5TSIOMgcKRJNXi38zd063oxSwP5oz+kARLaGIAxSJB1/mGQI6oYE
DV50xJgB/TsAj3i0c/AtEazb6JKMS0fXpnzzTVNC6Bz40s5BeP1QtVuN0tUCUkH4wCEsyOhxm31c
VB0aI1qhCq3BtqxBM/r/cZxLUwJZCWmQv7X3pHNdwdSCvuaiR9CHJ0ux0ZHC/8WJdE0AIDLFftM4
fugyRfGTF44NkObwCUFQhgCFPqs+dVjaPTMLj/LuNc9MSD/S+Edci1aWuY9dBhq2Shy2TGM2X8r1
F1r6ndF42zN5GQhg6egmGVeNjF4H1Le6DYgo/yxHqF7cUzuj370F/9FeUmoWFeSByAKdL7IEDXjj
TbI6wJGXVjBA6Lx1oKA5WNUsVXtZd2ECRr2NhjOceeZW7g7KPs62pJF9zNShaxEkBLcQYrPFLiWX
pRBOOuMbHlYzC6os2eaGM0JQVKoJTiHGQkvmo/9ZNAXyWPHwCQQ5kQKgypCK+/5cNfKvuEygGnhf
oDg95repb3yal4/dtg0T7zH4skwWjamytEqGysYXPrCCKX6ZtQzo2gf6bzA3500ukCr1Zi84wTYu
cf0PlPn79cpPUvnibX+8i3QBO+B/DZrPK115MoQX6+s4lNGCk4OJ7iqNdglXEgHxOk2mrhnc5RQZ
Kw3eWOAJWHkWEnJuxfR8wxC4xAHeqDCGcWkXyoxv+BIUltiHDwN0E1x2auw+CaiFbUt8kXpMoE8e
SwgwvIxjVxTLOj6DcfTYasK4jgn1f+X6/bLfWYdovirHFBrzNadOCO1oW0PJU/uptiUpi9HT0V/9
x/WrjxrGPbf9bCZa9xhHZgRu16DGmgiO6wmmaQPSlVp/o9hI8WmoNFSErlqNow3+CG8Ggd6oWPmz
H5PA2bZhtrNfF1Tit78cuSQ3gFAdmT33I7xycZryf444rC7Wa4PtAPRF7dPJfqfJb/8YQNNMtHLn
ziXOMEI4BSPpb23NndAtJi6lNS5Er9sgv7qBxu+qkw5dpwJdxBQX8Kf5pAazmks+xE8aFBzI3hWS
2cjS9zY3kykIUyXEjbAX3eT6DzT0iRat5qtpT5lnF9LYCsdYfZpFp0qzguiYkrvXisiJezJfcWoe
i0Nf2/acuEY2O6kg2SSwOZtJYt9HOsUvs7iNHMYqYQkKQV+Ad3qqWcLxaZDHSkXAvwnlYia8wiyW
8qOAJ7ApXv2FWXvEf4aU/vHKGrjQvpjp2f080crFoTF/OSPgSnlR9huZoaqqGffV/gIuslhhNDUJ
zfTrKTkZVcMmaY5VgRt0q8P1Z9zcJwWbaGHGCGFxTIMt+Yt+bbl4dxqz/T17dzKlDnWV5avCJLy5
ZR8fNVuCfqU1yWpa/P6aEvxKQnSx2XaD/xWcq1r/clASSDUvcCUcuqYtamOgVRWBtZASXRIEpqNO
/tHzgnc1GIXwQ4X//bRWjfJ3PgM72AKPppBICzcOMLGuWbeIfs16v/wUN/VA37Z8NTmfmjkfDFdD
8YGLKK/LOaPDfQX3KeVfZY803ps8MYXKzsx1s3v+ZEyOpb5MA3502w9xajGWMxqVW+nirLDGa6wq
kDq1aNrCzNXDRqDhxEYwQYGIenaMCCJ3OCAhwxrX16E3IqJohekv0TpIeM1vWsoQ1jEwgk/ui54h
Nw4ZBq/ayMzt5d52/Knbbn1iWgDtKE0rbA0iGg+ooJ/Ou8ZpQt3wWld+tyzZDITov6zBmhLrmM+4
WRnvhet/4hrS8z6Xf1rTnBa5B2O6iVIYZ1NuhCz/EPDK/hHPjAvuy5e0Z1uMk3ADr1V3YZaWaGsP
Y0NEIJWojS4ed2BGZWHzJB8wcVlzEeyMyEsajJZ/9eIm7Fs74ge1pWpoVleKtc6720bVWld8gBxL
EkKjLxuhWTcqUX2VdFrB0ONHeJnYJneSoS8QlE/0+tgx0P4QXuXHsPWJzuKwE5kwbwH0p0Mv74Y8
/yNHLSYuxb0IPlUmKdeV8r2vzi1uhRYGOq1qPHhEbxaTatdLrxNtzeJ3nx7gkO5k/IlYpBw+XPlP
k3TaWA5N2bCirQ3RgOHkeiYI/eOZFdDkXuIpMrQqRzPtU0uf8FjUhv60xfk6XePF1QFkGEMUEUqH
GcECI4HH5/jOlBwqPWV2bwyVOEMG5swdUblFG+wNSubxoLEdsG86s2BhxemZs7kXa4CD0y/ErVB6
L3OUXGtBtJiVDKMcIp2HInKgTLO2ylIO5XiR4tUxh3QP2cy3/0tJN4Oz/TXXYy5RDLDyDKmYIOLh
fuCqlhJcC0so3QYooXAx8efp/Dizp3HIVCrlLFUQiw/Kie6tCj5kqhqmTxtnp/AZm5+GmiaCYKnl
L+Zk+mUGZjwgEJaw1oIHA7nib6vu3feSw8o42BSatqt/PguM0g4TkM7DlIbd3n/Fw1f2sObSpuBe
61ivWAy8aonsiWUgy1k4AumWjENT+QVM+neUNnBdfF5JxLVbs2LfnhcBOYiY1Dm4TxYF8EgxhpVQ
pLVY/eJt8ezrb7VgniGNNrHLOXhgSQ0gM/R76VLSDYMkI/xaOzQnhKjoJfC+N5e4zs/vXXo/yrEn
4KmPqvW4MfYrRLPTjCUVsejgtOtR4WaeNR7eAdwJNQVOvVQmSVOjB9+qtbTRNLyJ8WGvE21Yzxhf
ASDxxlT9mmOamkTkOEDkUY9bHS9gBi9KucPxHhVwjzFNgYzCwLxwZ2Abjn92FGob/XXq1lvMPXLX
rWU36e9iZ6f1tPBWpq5u9zXFpE/K3kkUp0/AhNbu10o3w8flzh7DxrYfjXgKAn8ymTDrYClHVi9g
kmbFKmKlN/RE2zXDs/M/hCf5i77VCpwMjnl5bgV8DHT50eZo67Sdg8mGTHAcjKUZ7MahurSbZBYX
0YjCsmwTnmQSG1z29Yl9V9h0zYJEYH3ZSCV/oFz4iqZ7ISWwWrbtA5EHe3ESkJik/IHz8yifrbbN
isr3xFTzdxbdXtkXyyfa+kVOQRcj0W3L7SQQ0Pmzrg6lz9AbYvgG7UMWKwhJgfZ8itW0rEPGl5xg
/EnTk9yUfuWoiANIZl+DFqxSgXjIPum4G8e4RgcUdFJbtRQaaJ7XQzQ7gH0UcvxObH5TxJs4b05S
rB3eSF5XpQhaZpitPO3yS2unyyvY+i24MfNT4sdXmYUnjYIKQs4hgxOCc1pQWDPrrar2NVjyny5Q
5qyeLamSjQOr5yImbPk9oEkDZ9ZsnnQAItojEO/Q2D0KnXckI9y/xGZAaE9cvk3Ri+ifRvdx02U0
sjANyXi7XCvAVHtVYyR+V51EONIYTr3bBvGDZSoXzSm9iSBEmPxVtcgQ1pzwFFCbCyYb7ZPvys+s
TvN9X9jmkDtlqCMDyeyAAKFF0Er5pHg8RRYK+oTDAKaCqewZjmTb9Dj0LeNI7q81ExstaK2vDthM
dfT/q3SX3wDBlU0MCqK+qQZpg3bnonB2fWGWoEVJtDoWKKM7bGYvMMxSd3isnKG9Q+L+A5OGG9Kn
2s9gs9t1MvlcZvCUsIKigFDOSgecLhNxJe5Bqf6sSemP9cHAqiV7KelUQzbuchHlcwdd43tPSVE6
wal5k82rZBD4bDVFKK9VAP0gaH3DQuLbOMa34Ilw/5tXKHq8k1VWbxqL+ODqo7slolkp3q825lxG
NwYCIlECx6brxzfsryB17img8jrT3/H4326A5dVFsDNH/18D2OeXWbhHAidBoHT0gsu4b4NljG16
7dRisdVos+xmVSqTpcLoxAI0eeg8r6EUVW4xbCkGFYirOmnLlYkbf4JHlm3mUi0Y0/VtftJ4U9W/
Q9BVrov2a6oy/XZObhEFp0gwmgQvI/rmcIfPC1KPUmwFjrbtt6fJel3E2mLBLWxWm+RGQQC8Rl+D
YMlceTKZ1WiiNFSQxQCnxIvo/pn88/XOmJb0Ck+BHTMIyJmHSwWCRVGvCVrCdaSsZwerZCWzmNnw
IF10G5436n6xTJIoFUtnV0XmEPybgOdhIJIGS1iOGx3d41GFwDhn7N1S+9BfYAwOMWc2VlhbYW4G
MH7DicJiBHXi0RdO3Py15h2inFwjR1vq8diD4Hi26XIuFMmjwPDZw+VWGM1B0sB9zJ9haD0wNSXO
8AD5cYEWYiH7SeQdBnSLQGkeQ8YZU/db0OPBwOFU7KObhUkUOaJluNPVng8/+4W+qzAbiZQ9rWU8
TXaC1sO4k9Z+svA2Ztzdz7dQpvm+MOLez5xvKZWBXfWK8KYZdVC4t6q/JBWnCarC0b7zER3p4r6I
gBzFBQyODBCpxtipCvUD+YDImxp93oQ01hJGEmcoikgvOUMMXQ2YMhH6zmXYb9csel5fOkl3L5xd
bfX8x69uykkBRm6zxzPPCsewqGM2yn2pvlwwGCNIuZVMsvzldNnhmOdyYSZpDn5rfTTQWjq4VLXB
u7U7IQqcJatlId59k3raK6Kgvuu/3pEzwEa0TjkQiItZm2j+hWbTSyK06EKbJdlnFuijaaJHPYMH
KmcX5vO7u40QzYfhZJkkQgpMTXKOaDZJPnPgEvbpQEVLNnr9hnYN3/TIhM9LR5/FtMHcVehPctiz
dshLwqxQO6/cXBDDkHcmGjQTBU9yBda73HqMYcWMoVvZvPzl+FPfePNDrAtD/HEDYy+payDHhkOR
pj8B9w3l8TyvTLM/MHf4IiGX/p6J5WLGQ/KzH31WFAPPVyVcmPWH34odEUY0CqKCSuIaB99Gyuw1
nAPmnHsIum/MYGLXw/1N7rWgF45FSHFfpMGoLGyWVLyCDWsVObyANoWpK8UvBwafk/a45nYRtB+T
+WdTWQPAfcfVNz00lzXbmNEv7r7UO4EhHfqysVFgnawbB42BAmFpoWHRwL0/+NBMYZWdlcvlQw7N
k7LECVtBJcc60evEmyBOt9fCPHqNOQz50QIknxI28H7Dvkqf0Fl3Iy3OlpPOYRAunX1TgQTES54f
h0HIjO1760o/fu2SU/KFQ+XgspannTualccVhw6YKURGKTYzQFPxLWnlJt1/WQiB7O8LEwLBoyxw
yFbz2DtdrYj5SKwR1twx9sU65kj0JzDJIyY1CcNwYTmXMBHmKkP+AwGaBL7EyVgQg0OyYULSaq+m
cIAZ22Wlx+lrmMmBVStt4b9zmaR1Uo4Hdj0m6gEQJFJL444rkxB42mjbQzzZd25QxGEeCIOoPR4T
oAh4f19IE1CKNCYEIbww59ScJ9Zp7PI/NXzMSn5yyysy5FWMjMj4AcKFzzF1U4njacfX4CSr54KL
SubujuGooFMMVnVnTS46KbOF+sIw6jmXcD84WDEZPkvLtQi246yKx+3cK5ct3NscaK1JhQBxP+Ft
qC87Urnyaajy9AEMbdIdgONSlQy1iDOyHJkxuEbRM3ww7wc5PnF4Y/0IcoHV4gwclDwT8Wp3LY9r
ixKKK2/jUXQvkFfDLIUqdh3MrgPZyxzVNAa5Rx0L+EiKub1BFtN9vRRhAmUuvkunIQNNVLvWj0Ji
zt6IbYy5RRZbYTzfQLU4J0A4Dt0S79I7zfSqh77WI1crMcISeB5aC2CJGHGl8L3lLMb0heY1nA6/
h8ghoExCzHH6TnJ3qKGcBT9uNf8Alh8sUyzrQy/KYsdGGd9X12/NnEAtlAAsrSQS3yXy6yN5hXLU
7AbdksZmpsUYdoiewfiB3cNMVsS17nU4Jqqt9X1u8tqqeZzBPvoFcirtSgEVhXB4+wZpFTe7oH7x
W/7TXNKCpZhbnuS2BCyKZ8VYy15aom26I6q0jorb6RAAML40rqiLqSipcq2PP94S06jqXvrZT23U
051gGeiXpokcopZYMKisKjU+dYAafn8HI30UzbeTa9HP11zi0rDTC9EUrXT08Azdq1nmG8snPjhC
M1/s2Sf4J7uDEIvJGsQHi/0pZi0S/paKfXHq6LygLm3/nkAP6NcWZt8n9FS12Ea6maaQNxX+PyZm
FfJAEbYUYfkYsI5fcvxuIL1UYoHVXO0T7YJqcp+ix2Jg1cH+fOat1CefGTv8l5QAtNV2dqq/eBJt
FFVFwLPXoKTI8INfNJW7e6H7XoFbhPYHMvRqy40COd1oEMLNW6WGsf6LTmjbFM4Gw4KKUAmem+Qg
vlw1/9a35b0oTvaQY4LnIIBkkJ8g+eCXY7MLWIPkI9j7xvxpjZe8uVg7gim6gc/u/ZKG1IzhIkIA
BglHqQI4KxN0HC55pxZl2qrw4PtyTmoGZeZhpv3wP5DcBac3tI0heRl8HV/Q2eFNxjhdEmj1pKgi
4zCLuRVdBDUE7SsFG4+B11sbQm8kRoPtdvbgqMaadXUKb1Kigt2xjfeHUMMQ71DBDzrVI4HBmdj+
VEbHDMF/ENfNvBAoH4V1+URYiV1izXT0jLSpYsaHLxNVJWC3LvfJhnuzrvORFk2+6viaMavMS/NJ
pddAgt49O4tMDXjtqQdj/uPBtIFlcr6bPHQeFjijiKM48xfXVUMunQGg171oi8aShrTzkfIBHjF/
zFa9Q8fmtlyNPcAOVwTskum3wHwuaC7lYIjNWHNbwpMP5mR8wUzJMpxMq6J+CMmCS3zi9gonedGR
Xl37YFK+/62IOW/IRxX6udRVxIGlU1w/ehTDE9pDj13vQtxsUt3mL0eBlmIz7/oCacqn4jyQSj2Y
EVoz+7MTtJYR6lW6DES8uKkRlRyf9wZ/5Ob5MjFC4AU1XGZd5TpKJdoXoUYlZv39M7uGNZbaCNYM
ALPB35wkPYFkZmLCswP5+iDABttEnE81+mYsY5YMkMUYdJxpsVdmx2o6kkgL7dny6UtnW0ALPE0v
5WVgPJwSG+A0K+Z9/eNVEV9dc8EyUjL8Ivg3c/27Z2fRfa/q0lRFr78dzUMWot3nmDtYlc3Dpzdd
kmRJQyjH2QNC3jRnmul0stqjSIk6g/i6sIV4AepveKGRws0gHBwiRw9IdldKcKC+C9yKt41xfrge
i1+2XZNPfnUeeMt+7rIb9M7imYB09fG7p0jEWkmm0gmkuhL7ejsyAXJOvuEEHNrLgOajXjysOMHQ
0GDHE4qSJRj0ktByev08oHVtLkAojpgASvPR+T7oX1qQ0JnC6u1N6Yi16nDvBJp/SndU2AAkpj+i
c9f+gRhqRILvb4/Qbr7id17wsydMFrjugFrLg7i/giemQgVFn6PiGfEJHfbiRiXo33sSbxLIJb6L
06m9ZmQIQY1xoqsjJ3YHkzu7bRSLxXvDZVQ5Q27+K0Xjw0jjYi7mn5rk8is90ytEQLvW8fFLfSN3
FKbzCWOgWvl344aE8lcOEVKGsfMGhTZ+x0MQ/0qpSa08tzoCfIw1rnENSAJCAkGuFaZ7cW/rc4Ft
moQsV3nhoEFjUvYa+Iz1zWUCGUhq+VlZLsWFGosEo3XqvXCxBPwXt5POns7fe/Ld5JvfLixw6yua
3XvEuIGB3ss2pGbooAMCMM79gVPwlHfUykw5Qm5dxh8VNuGyDbTsDqRgIKoD73iObqcykol3UKik
0/av0EuL2B52FR1zJHIW7aUapBFaVYzIcmvdvN788/d7+fhs6H6DwPjC/Foaikoo79zGfcEIHfsr
ReGIygEG1bUddsD5sUW3/LwEWZ3XzEnoevo+3oPFfL6qwPkZk9mQ3xATF3NbTxHvopHkxpfOoDJK
HyPYAnjbJDkbI2K0GavbIxfKmLtdbWXlvz3B1JlfKsgXkVG6xUwJMhpHphxtcL1eIWkgRtMt7q+i
gs5+OPjAgI20PFXR17/bLUhDnqtOHDRZR5PEZyYT8XBIqWPzrypYQnqTP24HH99thzCZHilVKF4+
ktvepmDeHWh1tIv9dsx+dp3lbjQmRdtd8xhJT4qG6OB/BU4y7QD61kT5nMwUC/gu20sxk3OhR6CR
2QBDIKyamv17VDRR6pkRhQx0E21kvyqmom7mvhRJKHlLXtjf1cZs8aT9MgP3l4AoNzf4EFmvS+52
kiN/93NZPzw7CZ7kK66VTyz0zTDsEijD5qNAiEVGncmmJHvfvxzJh7O7o7UgVrq/LlssYV+yM9aH
QMnBX45Yg1sz+A9io01QKE7zR4GSFAtasEZInN5+UssoegPmUd3Cm9OPbNH9ts68QZeN0AF8Rcr3
Y+fjugLeTb0BvITlT5jgMR/j1DGTZmSYhzqmTN1xZyJzOv0lokIcNQKAS3eYYHJv2LZ+D34cpgqz
egIVF+DBdP0TY1sJIG5sEm8+plJ8Jd+KLNndL0xEKalNaW8vcXA213gDrJphbtp0WU61eOKO6+ox
v7E4o4rXMQ/77I3nPSr+1IJZkTpzaC3f63jzzLOYjFL63HLGKxMlY48gOmFAAriGaQ/fGO2mkdb7
hKn+ZotwWBzMXe0fcM+J16omqZkaeSdkaiwz41+5hhYa1VINoGF0+la2nT+w7d6wS2ZCYH2LJToO
mutmOJZrZjvHqKuD5a2wO4wL7GZNs1hnQoHTknpDfu3IHyDW8ILAgyVNL3eJdtyQUmYdqKKLEPF6
8d3sjy00w3rHO34viUqqlkWmU7PQREF/dsSC4dISl2hwQlTnXM702MoXLQyjmblfO784gHYzQXV+
v9oYlzn+eWey3VlgvYIUe+Ph4df3DRDJTASb60elWx4VJybHlE3JLwnw/Zbsh3r65SeSGyd2kR7D
mCi2fhWYF47MsNOvScIcgrRBZGwVZv8HN2Lmolt24E0VtF+FLQ/noxV3RIAE/42HkxfkFvd2qI42
Ee8+5mNorH2L5lNVp3U4vEl+zfRuwjs7MrP4jfjp4M1ZKhIaaVfjnANUM4RMCp8mDVh1KSYmiEoT
wW9y3LcjN71R+U8w/4LMUkv93OniJ02Qm820Lkm3ojA48bui7TFY4UId7uhKln9NQLlwOXhymMg5
QjWwbUjl78pU/s8xQFA5MJT2l2sEYQZw7baSsprn/GPTt+grcmAAcd3vfqHkpa6Qq64VDtbJPYFO
WKdsmRtuj0dmGa+4AaF4EsIVmVF4UQcyEtTA27LRnGPAa84wKByEXVsWhwhtAx5LYFuvMX3iFJJI
4P5Zd3vNJXjTanJEqRQdRWAzKVc9/gm7V4EDuwS8CayUncYPMiW32PbsOGQluKtePF2ico1oK7dR
4eixmeZfQK5D1X9XZkAEJ4/9Td/9Kqsam64xe/+KeVwSfp4JqgmSGTaKkpvqYyVBtOD0X5WEolek
dz6VtlF1SwCJqWVhCJvRHTmF13WFlzDMa1SIzW24RBbOPu1JnzVaNGapdLmDudGkMvs0VsbQRn4J
CR78qrCdxWWPHpMHIdYsQZVz23aJ666zI9UFY2nvKatB1J2vC3P8Gv1gRDlA2h6C5ZMPbJNFVGTy
9ZqXf4IAKNVSmX954Z7jQv7i9ARZY5e69JOEqh3XEHZznBbale+UmvAUcUux7hXptyd4Tf3T9LY0
ol/qZ4ImdvZ/LGKmvoghL4dClo0b5atFrReMyfy9FIij39WG+cA6fzO/F2FtyQeqx25o77MC5/tS
jFLgsZKLSZIYi4nfbhcfXHMpxeM+yH+Fqlb79y7tWOPi9UHz2QjRYAl6N4CUGH9/NcuqyufdXBAv
1Mj7XzN8Di2xg/FGgWcmmnWSwbpUXanwvI+v84GkvBe3DDF4qWboOS/xGpC+9xoOQ08eAjK1iDy8
OGTM8K55rcT+QRJtbvjmsYy2E37H+9B6C2RQ2V9FPlkf9gPUZ/jLMrSgNAzDchgpi1GVD2zawI59
mBHvqNtYtGkIsLVD+t3SHTrtFOH6U5kGPmSoB5EWNOa0Fpv60C6IUpuTbM7gRl7cqKkA4fxbtcD0
uF1rHG3mRk95fZ/35lamIVDFKTvTjcHeqUjlXkDH/k48lMA5cBarLA/FVxqSx4BeadyUACVpP67V
GE2uvrHQ7zMFnAr3sZMo7HBKuE+Pj2Fh1cQGwNQrFHBBYQs6FpYFQ26SADWj/+vICx6ezIuf73MX
rtHwQLaNSK3L7r4fmGNhgfRH9DrJxTjqrcg9pVIkWGh0xiPbLlj4cyqjGxewcIWClr19UpeRZMaS
N+gNkwY8kN9iXV+Vf9CSyR+VbZ3TBwX7dOHHktWIhbDbDQ9Wvpdl1QbKLK8nEgBxDtS4TIWlw/B7
WEh8uXeCCLgVCGC7lXhSW3w1HnMUsSPPb/mF9RquXYgT0jkJbEoGCXs2NAfExzq7VNKoMAFqIuBD
t5fImkxwpFb6gwcOW8Rfdnzh8QzBG6dQoM6gLi+OKz4HifdkweMvKhVG32i2EOTRQ4oWVbdVXq9K
IoPwSqvU/Ypftt+R2LDFtwsaDFXVHjlPvjGaP0LSlWjB4wLHEScMf3ESpN2vsfWiD+PdOOgJEtbj
tComLzCtIT/lPSUw9Ydw+C707nwYS9YkTo6bGQkwwJx7mWPTep0IXEyQ/eTOGz91oHJgbfvOMv6K
S9UWJlKWDMUEj7G3gVThRAzAgy4C50cBT8J0b4PeMImXAqBqPjmP7mJVYuiUKM8zDkUuq2NJpIYq
0WEbiPJV1+EmlYM3ICTfjkRwcCGnAUXu5pkJB+cOybKSvMVNVaii69QOMYhGdUjZOJK+DMFwXRrS
4fyusqrBGwfwGUrcq3aTXcnjwWCNv2/mDbm4ylTH/mowQ6OADAlnMVlDC5krI5pUM/qqp3nZAycc
7XLyInMdusKDr9iMAuVFW78oA4UmGUk3zFF0l5TZFgXr774TaSxrgtJyIicpckQt+nsTsXiFnhIO
QMbLI0zSlIUNfpwTbYL61eSVn/6jMP2yXNtGnMy8TAPNZ5AK7FnY6I81JjK9BFL6Z2bCjLZMEM1c
sIyFmpdh512/DJMYGvXlrZoOHP4khi3W+tcOjB1q4yc7vEdaAlU+g+rVrM4hfNfF4CFFH18XPjqh
Ig1JqJg/4pHsCrCHv1jB0bYX218EdPFU/CVuV+V9Zz91EtIbokG0612kJZUmynOOycnY6QQW1qNq
opAJm7sVXhy6sjS1SZ0fAe1k4k8FqAL+mt56yK8wrIPvd04w7j9Sukl8qEeHyINKmAb485w1yAa4
faf6WcnnqVIgUubGsdj9Y1ZO4Kg28/pqHqRaeGWDnpA4FHn377p8R4BALFiibY8hCLzMPkrUonlv
BTLIRH6Fi1j3XTxzMVgINn/LADb8DaOdS/JplgVTqCch25z8HhOc3aetDqMmibHHFeNvKLoEGy17
40VgGZYY/PqosPYiKFDhgxqO1SaopsMIz3LV05IfxnvaMJVfX79cD4G+baMebuAS/5QS4XbzuNFF
QC9Lc4GPkF8qU8MiqGZ1fO+9xV91mVJEwsJIURPhki/UIBCy/0YqcNtMqraA1H07i/Ooh4vMoEfk
vwoCCFFNXZTN+xI9j75jM8x9ZVuW0lszAjDZvlLp+YA6TLgPBoavH3T6J9F6ukL2gadwpcw3qD4X
whZicKPmS4YM/Wueh1zcfJSGzvfRN2zFRS9K/HRxZMqdI8eTSszz77v49DF3RKKUFR7PYtehtUni
R+LKAgdzXmwXOapEqNjp5IXa1h3N3mRfrfrE0APedurOcLhIVp1BQpOyvOWk4uxKRSzxnwzVI/pW
8iMeNQlZMWvwN7DwG4F/5LYbwPQR2JS3gu/Dm5zQ+wS7Og0qM7eaiIi52HzZncQ9PGiLdR0MKuWy
CSmKg64mJSbUmdD/PBxNBkuwNGMwjs2brr3N2KJYfEg9TPiyVdNjnb05s9LKC3gSfPOAb0nWV7z+
tR3+EiCtZyPdwA6EVp4yyTCCpVgaQ+ZsvSgd/jpIjkLd+nT0pWm/y6mlBOKtQq8hIK+vwoH8gVJG
HHIGo0E4AeL5G8ZqJJzzkw1Lpo3313AkMg8TJRKq/vsS2FmZ3Xgmu/Mtaku8nPlBcDjUe4CNvt5T
LDN6s6FEJFqEsXE9UEiA6ZxYSXhWTGk5JSQeHVpzcghvkjjvksrxb1aj0alil+/hdouwMOBGGheP
XCIFDDFGjSVws8P/fEhywdZelS0pl5JtIWeHU/36pxLBJxYcp5m274YJaJRYQytkYBQPCw66u1wC
0Nbmi634lwKUJ2ZIxFIqreCydmtBy2C85fORo8rdODYg155PQmWVU7pOMD9kOTh5y1FnyT4HmHx7
d26syE4CpCAC/EsjvqwtwzI4piCE77KSf+HFPRFtHfK6Sj9Ozu6GpXgm4UxexI5HOj3+UJPQnW6G
7qodrxzzTAOslfExGqBUBWB364HPpWXm7a45/GJMg1QqDj0fPtdiQ+dZU7l+yc9DiZv+3fQewe0+
V7Zb4xbg15AOzp0gyyJ4TRsTb8p/AB22A5z4OEo+BgoaMk4wMSIQ57HbZsE+acZvrtTAB/TsZdyd
LwI8bWKgIP5NVX2fFDx2Wxbsi5vi8Xpgkms9FuZxSABXQeqUkHrCvWF6hEnwyEWl0rxwZp3cr09Y
FAE6XYywn+/DgID73VwpgTQkAUKQTKwBymcpUlp/xL4abaf0Say0gUo7kfWNT2t6/w7aRLNSZsPR
Or6hkmubNr8MUfAJKFzjVht+tCmPZN5kJM4DIyd1XcaVyYboM6uk9I4VvNxKVghbGiwjiPv7mC+g
i0m0i/l+92VPRHEJEv1oqdSSpqOnhyrPRQNswwGFrQoE5B0KfDP+cPV1eMNNG2hW7/kBvY4dXJdE
FZEhQo4QAcNqYA1S3PTouQ8HUG4SwlPG2sWS8q0g6qZRj6IItobjFWQfVa1429NSLtcwnM3DfUfm
RcP+j7vnfrGSDMfVRHScXM1TmEbDI7prgJEpR1N4UbDBlgmz70cma9TYl4PQmJpXI5sWFsFdr0NY
Wuy6GAQGsl5BaKz2+fAPxo4qFRc3ZciTQfqgookrljnoO4XiEY+a8OPNPscxxXkBGvIeAkY4DzLC
nwreRDAIdGC1X2USCddEvfEyLkGHnS1blWGOe9Spu0Dn5izeCm0vdEFHQgaLAGQ8IdHESMlePWHU
IpWIUtsVDhINujE7YVgR1xxHrbR4BScqQKdRzRCgFKsM8xltbKmt2aVo4Oxfr37kpbxc0ir1JfB3
XB70Vw3PrZN0PoymsDtYdmgVtNaZW8lP7ft3LLTsAGJLyDBYP7GPFN2gEorN6KE4yLfalZFPJuwV
IR2SIweLafyWHr3zV/GSQjk95t/ZapqDl3w79aVOQZeD+kmZcUMZAN+WfgOqdiSnddswrYDIwzmW
340UT6iyoiyrzUL/UYfOb9qgUNn4zH8izAGV1Eicjo/Sel9ZoNoNrEtA+jcWCQLsJSpq2MXhdw+U
rmfQ0xRjVKERlWv9ABNnmb//CosFEPYcXIB8fFyeUd2S4eEHgyLU0fCZWmAGW/9ICqSRtbqYUXcX
ycYzO1Me6YOGOlsLxag5QkoNq69iMwwOeKMuXX6n7k7WrEp80q0d3cvEijd+I5IWb35LVpL6ABqB
ZiJwyiQGJaf2T29H9RkdolBuQ9PK+CgeyWYbZz7BsQyff0iIbkJHEH9t6gCeBb6HU0xJ68oay99H
IlAN9zujpPJG4DtzVmJ4bKlyke2c2hc2E+vXujsk3UlPRiQldv5L9xM/OoQxoL4e6Rjne5HKyG9x
DD/rGsLFVCHw2q2luv1h79Be76ZfLNzPbJG1AbNDMcsDlTkQpFzp1G2Gythcoxf8+qcrzqRXG+8m
NTC5lkPbi+wispSAwuusxUM3cMeMeWKQUPNfPCyR9SxpsYHSlRTK272J2IThGwFifqMUSZB3Xnmu
T6BmdohFudJ5/zt4c5sf5whjjVWQsVveMwi8lE6V5Qs1NDLhpZu7/0G8yuR6EojQB36ESGTwYnou
Fwg6KhQhAEYAGhGsVLW0Iz0O6z+h6RFum8M6t8sdIdoLjuZjDLI/chGD6Mb9+ADHP2cL173moeNh
ZkiLIpMCoasLAr7SrE8mGF2Y6DpKm66esUoj2IabZuv5CD+7AY9+Zhd+8UzemUNaJt/r2v4Ow5to
ObzHGhjq8Qa87Q1E+vfq6VAjlwdwWgT8j/uLKP009GyTnP6Lv+ISBO2cmsaDhMyZsEUAUkP1JwUG
OoBpIwrXKEFGq0D8thFUSwWfKwNLXclmNdl+Co4qCcdBRd3USfDVBqeU4AK0fAoisTpgTHAXS58a
DxBM18bYxJQ+VjwKEHbJZuwmwwBIguFaDoXz+oH63Owhc8WFGT1VvVKBiPzI6Hyu8APaFOE2Nd99
8tI5ac3FfeKC8K2mCqw93Lab3ETx5yVE5nnVLWmifgAkeERnFXFkDh1Dde3a1u4IlhAA4/48Dcwv
bNxN4hFOLd2MOQIM0UZav7Yv4znVXDMGj0zxuu0XuU8T0FbL/keL5mO7jgvOqo7ySIk2WSLG3On0
rMo1RfLnQW00cqI1JVgkgIQWt55Q48QExpSYhYYrNtpv4KKfe0AR3YqPFMfokOpFT/zAr4kC7AvI
5h9WIb/ipTXWiipvjuR48CHXmh+DrxpAZwuYz+M+GBFbyp44NyKCBxENgqb+PwNJrTJAulIQwkiX
SX3rDE6a/mjTTVQOca6ENoRWjq4AAP7xfiHUvO8l1yZCv8wBqAWHOv+rrm2oJVbAQ4Rx5bcOJK79
Vgy6vHiQ/uM7x1a/Q3fPTYSzUZSPV7A83M/hLTYPosptNARj+bOt6JfbeRP8+ki3prD+fI6QUwx5
Sd0hYBW6g7n7paB6PC8Ah9B6y31gMoHeLkwgU7qthXdgiVwJ83/QDHshT4Q5dHu5+MpxQ+Uq58Qu
PJBAHKckzT06ExSwmBpt9PRXb8QXZQ9RswY1dtugmKjgRrmWWI013WzW0okk+JNUg0Q/jdgYWWyo
2ej25Y7bfwj0lYTMtjixeD/gXtqMNrs+ksZqXk+6Ig1p0Q6c3mBN36M0QpsI0q8vOVhQcwFxbt2I
7Zia44MY/+OuUjJQm+wMt1XUwI4o35SBEXvLBuYNNLU0yOqoeuj4ZqIu3NWqTxfgRKhJ8/a33ULf
XHIdGOhf3XvczS7yhnwlBLhT0Fu7WSEaO+rx+ujBz/2n1LzxiT86ChKejW2yRlGyFHHHutERDJGl
DYDxmcDMQRW3nDkmT0ZVM9rwnzJS2k/CACqFGNo3U4Iruir+daj2K5/XE7Ddx7Rzk/qN5sa/8fnw
gVbokHq52rZqmXMpeP7uMzu6sgKSaEOof3FPikHRKUH/Q8RhLeB4daRd1zpbdAbyDQCNRF+VMlG3
wZixt3x3dWqEnNDAwXeEd7zLI++PehRkgyDlp6QVKkz5qx5D8ZVqbskboGU6fD94fI+x3NA+pxH+
mgPLOfb5x3g1co5U0FUJXy2FcHafB/MP3dgYcomDGoTf1FpJVn42TMVDfdl/dAFFF/RfafZpsZ9N
YtdXLcYXrNLT9GVaQNEaCsfu+w4+c2H9OhBtOd5OwX7ywh4dodBdbiG4sfDSD6Qk7vBy6XrruR59
4APqQ93MJU7FgGwqf9w3OvH1K1Iyb9fvEKI9Vl+Uo4x8u45LgLvEGJy7m3DGlN2mmt2bwhXnirNY
+voarAFcWnArITmUox3ph5KiuxYYCI/Eq/GnJz9buveuz7qyfqwRlC8PK4NkgFWl268iQuDayeMK
HfdRhmFrJ0PXGf6bLBth3lXHdm0ou2/65jOxy+4Be/UBEXz9sxaZ+wkkO0ypJP2HL9jifuIS270M
Uy8zYV6+bA7jEuePF4fie1JmODs+1aJa0YU5wsAuJYWMyLP4z4lL+GjzFPY6x+TlP8Fxz/YuEdic
22qU+NifCqukivdzxgysLZL+WPcri7KZNvW/ybiA6kyNuvSI8yayOhC/FcTJ6I0MkThHy/o5tcEU
648oFsrA6NJd2pediOawxpAkHbM8sCV7C8BLYcdaSTmv4dhimpoyqk7JWf4f3LFZUbw1Ob+djd7h
g8J8VM2+vYuxoIK/RjNuIrTG/V1OtW/VSZdgAa1joP00J2r79PZH1dLZADqSNpP5cjXXRSDArLLo
Wg7u2Omb8ajTnNcjQfmTO2AFBwLXv8JVJiHihCk+CaQCVHR5LvE+CogGYV7gRpvR8sE5MfhnpfNq
oaPgcO9FbKR+a89+Os4JeBD1CyKeR/JSDS0xK+IjAqLPoxyHOIvvaPPrSn0Sq10CuGjTX2Z+m+HS
egBKHqeMggl975yVIJuipC2VwHrrbVoMcXFc/aC7BkM5v29uJPc6mE0qBdZwjVzvXsX6qFo3MWJB
g5vzPl9v7R3QdIXoew7PAjdza/jGOWRVytOKpg6GOi8c7KuiwyC1ZxAZmG0Ett7A5MDXykeNkWNt
6RFeXnLXOT6hGwpC7O/J1lHMKLx+Q5wExK2RGv8dWtJB6uziX1l4jT46653YLhzQtqOpX/m4Ouo9
KIj5xZeyz/4cokYRMarSOkYmXLTgtqJ+b46FhIuSJfj/v0F4qbxs2gsdbiJNoJacGa4yEMKpO3FB
QA8Z5yHEUUQjSsOTexQnIiRWbRZON1PMokG4prFQ4kyF30aTQfdhJgl4D//jnmM8OFrNn7zTiJx6
W8UiZqCQZxI2pAqLH23vFNuVCY7HzuHDoO8g1qthiKY9uDTF3IZaMmK1gfBunpI0nSefKmG7/GRf
xnM5vnc5xuy1MhymqD/5lnE4JmmC7vZNzAb8cE+hTA+ENCELZ6FRrcxkk7c1kvXsQwWI94IygBBq
rj/xbSCfzMhFJYSVjVkfSt2tGgsa92yyZwkhwPbYZO9noytNvIbA6eXsjcwq5VGDXjLABvUACEpc
Svz2AdF6NExr1xWSnOVWmL2QD+QXwJ+vCsVaa8gkzZLc253szixpl5d8x7HIyq7V3HTtfnLHbj7c
7EnzpsndWYzEprGMUevAlJCT9BwXhbGOsirjkpVyBQq6zmoLo+k9dPtk47m0byAmvET/8MaCGjF5
sk2+TDDcrrxDgkP+qzkpH2mDDc0L/G/5bnyQ4NMsRkrN3q1Aydt8tDNLHQdt9diR8uA2A/ZvuEnZ
FiJVR0s78WohqJFQnLM6YZOIY5EvyoHURtbho420H5ioRmr4/2EDadKjr2q6KZvmiPOH46trobO6
G0/a3aaccodl7RWpQ3s0HqS/CJACKs/diU+NOw08f8vVTFOhOBtbe/JEd6BugnCJrLuJFeikatF/
3yTPUwMWmL4UtO/F8SnQdLzqGjCzy1JV7GGMcAx+LLy81XWMU/7fYtapS4buWa1F51uOTGxht5Rj
1extBrCzB7q+kYagS4b/Jwqrm6znUKmgHNv9AIPVssLZbt7qvQMiFRg8zHX7MYHEDmt2luDuZuH5
61+7NPPCTg8Jy45bz3AXlBX4juFFK6PP9MSZ/iC9CSh+fm0noWeB7VMWFwhyHaVNwJs2JdVnTgwh
KcGk1ugxzI/+gzurDyr3RocRCcL9o214mSe3PYbWGZlwWp26/+IwBl3MePDydIamIn25Kn86Knh4
aeq6YvVgG48f/ZwEx3cMLi3W189k6JKErBVm/g11XHXcHrkcn9XfVAvlQ90nxMtDXfGLTfZEkXSi
1udWb+roDykMNLJ/hGju/AuRWu5gYmWnbLLWeVtHJEli/w0OCaS5mxX+L8E5noGuFneslUfRRLyj
7Gs4CU4ovfxm3BOHW/8Wex2qD05g8gFYD+tIcBG4xGPvTOADWcthMSJJQzfnl0mCzhoaxdfJbY8c
taZDYLtoo/DUrhihjid5PQEUWjH8KkI2c6H93fwu8RaBuvuyvPCHftrh8rTCdAfd7ORhlcT3nPiL
yizM04XNmPN4lmfP45livTXpMlHAd6GTp11reg0O3KGNuzHYCfxUiOuwLTqceuYvN+yFAP2qej89
BeqMG6Dd98kIVYHA334yG+UkreUIikWSnMbnQxG9FRafBX7BETjVrR40MO+VqYEXpwfv/E3uIcMI
dEd3fVnkRcliJdN82JpBvncS/OMwhClH3dA51lnRc9Bi/MjQfGUfE8pOjT0VxJTpB4Eq87UzZZox
/tMP+AC1uJYV5dxLNA5q23pPryqQWUEbPwPk2vrCR2Er+vqpn0SnoNTQSt6XBonv76GlKtiJgTM1
81pZDeeKv7IVEhSU4t5VyF1TEoSQ59Zm2tMPKJ0IC9fSK4/PzZRSW6QN6ndMq4F8uxmEFxlq+ARl
bYpBq5FEl+WES6b2GROgLkPy1uEgddZV8rsCnabjy43UhLYDOxeTnGeNbHDzje38xnM97JWSbMGD
2/SbQHmflYgfQzjQ8YaO7VOOdCFeO4PWwvp5j+mGpkikmjK214qppBdMIX+S11ZfeSNN5xTwV4NC
owv7X3pq5lceEytLnPHItldbMamJlmBYjWG0kHGcPpT8DPM9dk3+hoHDdYWHxvMIsjjrJLJmZLo/
dGiF8s3qzUuKsVovseksNEJmABIaon+gmTXiyFSwHnGF+A4dJuEzsVXYndQGfCoCnH6mgQBy6m/S
ZxO5+OF0ItBv8la1uld6ENFjXVFhj24kt81LmDJe463X4E9fBztVoeA//VExnqP7LCt7wO7YXRmf
DYlHJx/ERAHNBWovcC1X6l9f+SpnQsC2DII2baOTKMqOINtb5Co3JsgqjEkCUIyB9LGl8WzJan30
N8Zg3rdWn957XZ45w44boLLUjmSn7kRI4IqiVphk0u4TnDCc7YOI/3UBk5NFntBHvF+3ibcRBbdM
cXo0gdg4pp05/FQ0FaZ2dgc9meEOoFkk9DrMUsV7yQVPgCpP3ty6JP/7STCNt0uNIigXugBPsW0T
1f6pHNQCRtX0xb3OtUz46nAk1oK2rRXh7jXmqy4ltv6jYilpB9jOngZ7i96mZb3bwlAH/WJR6o8v
zoo41FAem1OKs0e1lBic7YmheH5ghqmJD5N/fl8krMaqx462ncnOuq9ft/9gCYstR4xNcOUbSBrH
twehmQwkw1kArMbhcYVgcPWlZ33w7BlBOf81Zr+g6Kcrr+k7cqNVgLAsw6cFngY76Z+xP6w+etKz
4ZfgT5oSPscz+wvzREaTceE5ta5ZQyEGB86t+KvfL8beEpf+0apkLkbRC0C+EakM8o9JF0M43E+D
oXS1/0ju8mx0IKaLw/oxAFTy37hl1isIHpTl5MfuZtIJt4KUNCKzx7oRPW2cdgnROefLotb/Cqse
va3BlxT1zHfTx7jiMZc9AbjcHI6DZCcgZyWU6Dsto0m7b28mYm45hGKidQEa/k1Usu7Xmgf2NS64
q2CMTLm2Hq3oFB6jwQrW8OllO/kGesu0jpMk4h8cg9zvRzQfHlIUSMs8ok3R9liHkEBNMcvxA2VB
YBYBgUw28Tbg7CVvnGKmH99Oz6Ag8pfAVfh4EHyMcRDn+uj1LBYKT+NP/RGEIVQj5+jDiIzkPK1h
gO2cs4xKvbHUedifwxbJ/D4o/fBrGGcq+SPZjmNa5G+p8gQmFdVnm7y3p/zzsBu0xsq9p80YkmAv
gX12gs9iUI8sLKQmNppQsMsr7j3F6DZXfZJcQN5++fJf5lfvVYCJj1Q6VGRjTRYc7dTP04IsAIX4
KpymlC9Msgd3lUaX1CTlyBYOF5zkhNJddohINRyiu8ViMrAioKzE7Cy5+zCPwuHYrMv4SVqoTz9n
oLVc25BTGXkJJn2p27kLZ1txzGzj8YhYp7TaUkZLM7ujZlZWujbIdOgl3HKaFolgddAKprjO4eOk
Emygo+T6W5NprEBVDMFGHw6rCZS6vCheo7li4vVe1Rul/36m8v7Rbu2ip7c0V3FPn+VzYg8PLeN7
nDu3wi5APUe9eHOs5/oHaZGAhiU0GLFFEGYa17jO/YVinEbuk6BI+5yjKD6rX1DAv6jpHW3r8/Fj
3Mb495Ebh3FaM7Wokt6mR0trS/tx4pWWI4YtmeV2XlvEznu8+yszCFyl3/jfSjMjK06/rJ8cpccJ
1W2vG2ONBG8/S60aDDTjCyZA2n7pY07x4obdG/CpYoia/jJcFIqKNF34rItCjxWn9hZAp8ZzpaCG
HfMhnNbjz+YNLhC0G2HqAV8ktz2hCZdjZ1JOn5jaKeRU2/nEesN+GfyGU/gqYcYS6yEMkbIrNHrQ
0te+OsKLoUZW6wZA7DYhvX2y7VeyQaXRsp1IsIjF3wQ03eDZlw2vXNGn7GocwbjHopJi1gSYiHXK
Zh9m8PnmKSkvx5Frv3cClo3Y21NQEy2vNaUZoA6tBjTc6cQU+OIyZkuA1P6AdBzy71xzcFfeYw7k
i5RZgFyRUkhY6YImlXJgdXZrg3EMvJTs1GHTPOfybeJGU65UXj7qy0uj2aR6TARpzht7Zde73LFt
uzv4JXssDwgo3yyxTLZ0J7iwETodQM4drE0uArYklljc0dzR8rRIJfuLRfKdL0/4aD4i2bdGhtNV
N7RsxDOSew0tyDwuezmYP3WMtMvjcGS0WscdRjHtjEUHQyAW3bc00RIhdpdr6LVtFlo1OZ1okKaz
Y7t1pVlGBwrxj2FdQxC24bVr11MkV6qtC9cSFMSf2YKwISIEGEMgui+UH8P94j2BzsTZGcNwJUw8
UKx1RJ9F/kap6XwgcwXVkQabVblg2nLaOIQNNgEr1YqRvuphmgsfQbId1bOD2KSCHehpDvrv+bcz
DW7obrs/j2ULJU/ubzPjdoYXWhY/IfQYP/dbgbBR1mCB2G09ysPqLgJs2ExEGDMB3NN9UM43Xd7Z
Jw1HL1bdyifav73itQ/1kuDexvVLEW+L4m04hHC7Y6Gh395bDOrSIiwZB+k9eSkcKsZeszDwSW1p
mAKZgPYdQs9BppF2kVDofFLIOvfCZ/mKAubkBrQQzu3Pkc7LDDqXqK4EuHgTiOEffN/kMG3QKOIP
bXtdZL/PDrbDeCYGizWnqYhxMlUCN5kn9y/bvZ0V4lEdwNcW1hgJwG9h6QvzYbNbv6Li61IOc4cv
cWmovCXAdblHRmVlD0xTRhEMBFEsFM/DTjBPFKN0JhpSLRhvAPo6vauOeU4XpSTbN/8NJAEdFXMO
JyY4WzTlNfkg3AFyzDud3f3F2957A/FkgXIWXZ/O8odcsJNXvwyp4ZbQvzxutxRPWGDy/xeNpAPs
kRKvUtiHjF1b344hy7qeLEcfJW53Loq9meIyxv1MuF9AWpGhCSrCNPnkHrT3OOiZGzDOHJ5epxD3
v3oJv26bIv+0PA5umhJpyJGhY72Rks+GAh+tfHf86sDVfBmYm5D4ejFqR6xkxLdwORPV+4poNPNa
eRFs1kx3va4hu5NrkhSy5VUYL8cnuTURVfI2irLrKfoPlPGM45YTf6p0j3XHI13QwINZixUcjtl9
/a/M/y9EczlXUWokXIahf+CMA5ETHqiYHGXmf1JMiCUcZECd0oIOpk+QRTCCvX3AaM5WNIX1LPt9
DauiRlCmi0TGYweK0aFj5Ozdrw+0kmf7y4eNdi6Dwu9okTPxnB21thrhKqdKoSExoHsOuBc/Wtr6
TAmegaG30uB4gfZm2RCPbOj3bJotHSfGTV19eo6LNQ1+4sP4m40fMSH0jxztGUCw+PCqSvdnAndL
XOZ/isc9eLn9gXXs6Luh7IFE8oNhC21o5AUw7kc7Mh7vfe46z/qwpL6MQu+DDrba11Dqjupszqmf
sMDCue1nyaebFd23j/QrVmJU+aiEya4YTYnsgD0vw6QGXX7Gf9p+dzKqEk4im/H7B+ZZUUdiZqgn
CrxOaIowyNcw7c/VjJ+hpGumjSh3bgkYIRDZ2Xyo0QLmNUcrNhba8GB/yAiyjCXrVhePqwza7yWU
4eSFN+7DzQn6kgCHnx7fXKuREm8J8O9hLM/+BbUr8QsLiwm7OgtANAlt+kBPDAP0NMy2Q8spVZQ/
Z0NMacpNHwpenRcuXxv1QHrX6CED1HHL+/Z+Xl9t5q4HXHVek1IC+gDOT+M4jYgapUGvsmb/BZVv
oZk1kgadUXvjtunCXQJ0BEVZdq1mwkt5dciEUHl8ZcBdfRpwqGenUWBJEDab34FAPh7gXV/oXh/Q
NAzBTZ6xat08qoiN8nUQyM7Kj9kyxzyiS1JlgLuGeIgmmsnwKWq3LUd8WTo7EaiwC2UaD9iSe9qX
T4/HKJPYzoGED0rWR4LzQ67xekzzx76Ggh5aBJnVeYIQ/HV2KPm/4pWGwkSc6fCzGOLyvfdajEtm
LYFx3IJnSYjTtrg38Tf/0IlwGdqqKqjCdAq5XjltN+Gfq9Uq2ldV9CZ46r4rmSzuut8GJsV7Oq3M
dWwOKEOqPBqxf7pH6ZX7CiYJpdddVzGn7hqz+g3AZKUirylyTqh1DGtSgzy/v/naYXqvnpyMFNqn
eJvK24NoDtU9xzR4wcZqFfVHFtm/vM8XBSKhJ6Qh1vsD639/zW15rwUxPYG4MonL1qq2quv8sAle
ZhJO7L8UZT00g/dyZ5ED6pGo78E5LWfigN+MnxCjLUku60CazINU3T3V6fqct50UTI39SDQXHo66
b+Nz9VaqMYrJbvRdzEtO7abKnEiIWaDsZoeyqTdiVVFvSDplnWTRZGe0Yo/rL6s7rcsQGJH4Tu1h
q82PhBL5te276/J9xKkXGHPq3y7SWS2J5fZw55bBkU+9yx/2YaPbJ8FXLuraKNmRTBjycPUo3adT
7mjnfAoOthI74TgZImuVHwxTmpwgNdiYB2Wqq7x2N+CiWaNvQLc6o3HpyW3p5+O9dVfMqYcl1O5r
JaJmfSjNGq8PNHIJONUWcITMDbIn1etAM2M9K/+GWvl5RB/bJgEVXeQJ1Mp6YX5bM5zzNUugfmGa
giLHEXKWJ/CFhr4sh1wmyQQCLevZ5LqftnUtnfndwmbMFsUoF3AM7jHJD2RBRNdePhamm7rOb6Dr
5kIB1oU5uwZ/yWU2SFMp9Z/Slndu221cRrociLhH9v5Bq/NsubPE/sobtSbq02FAUiH5Xw3kxvJv
GKDBLXZwsS5WW4fPzzjh+tVlp04EJSssPqpzzFtk1fYXCLZ8Psj4DBICrFWhHShnhqr89Y+4lpqJ
HXRMMo4CTgtTBgj1WwAWaHpMWRpWd3UbXYLgY/kQ9hgeOrTu7hKF5TQtJFXcrR5xlt7aCrrZFNys
/xfGvp8vUNGwyJmCVHn7o3InFMNJXL6vCHsDQRvS/HfpsTdKZXdA1vsOEyC9okrrdxRHearnQvYC
x/aUtPhpCog7bDG9ppd2cVboByXqBKUZBZwJqp6Iivu9ymTRq84eHYAqBQpGufA7en+iWP7TjQC7
bCMyPZ6Nu7yylqX854E87cl1zXuOSn3ZemTrK7RjmnVCevAYNVU0DAJA8Yw+CmscMcliVEpDSaRQ
DxUVlstfilpEpGBN9M1DNR3+uBEUpCH2snk36zpdA3D9EarfX/db0h13wcBG/ULXoBE64kjOLsnT
vztA3hNfgAja3gAJ10GWucWHi3c1NO6qCKNjr9V8CVP9myDjJdBykghz9hp82PNbUrEbmJH/QOUV
68dUGO8bDn5ULQK4eVISv36tMjLBJDzlAiZizLymhWGb96ziQJocw6PRM1dNqujOvj5mV5bVoHvC
FHhvk0CuGg6ll/5mhZxt7VbTAzuc7WTkwzF/UA2jJJdBxSmxfl3NrQAY8Kkx/oAOgyA5Q6mwAmwT
D+Na0zpEAPzG/A1hptWhOtSGpokSrsFojtEjhgSI23HyfWuDMLZvKjhRWCwg1OJUwKoVk4O35UWb
TWB6pPOmd5+owEhAZpl/qa5dlB3mT9Mex9XI5zTe/2AHOLEKFmuYjiJnOSEb64/srZ9gpfCvercU
4vYwZ+7c75BQhuLz/mVCRRyb/LM7nIYKFN8Xdu/w47us4QzfXoK1m7FJiAOu0UlQeDiKS+z3YfgF
LrpStp6ru1Zxhw4x2gXqJ7VURuTKK/wv+ORU0VVPL4ujA76Zjm/cKXimHJhP+vtuBAliwduoNri+
GA7MTheqAYq779Fgkml8fCFzRjrfn2t50TsUBbDEiRWR6IsV5pof2dJ4wvawpA4jSRatEpyxxYPU
JidcwvdztPtA3F8wt8zkLdnWNaGYTEjRlGjklQoPbfJovBWMd4CWqQ6B/U9jFenC8kUlqpxV4wzB
LbkOZ1lbiI+h3glcIDMzjWBXdlbh09kbIPQ2fkp8MOh5xTZ4sZWJd+bOeM0u6WEH8izwzrDF9gVK
LY0bn4jhThxGr1mb4r/5OSPNFFfbjRfawOFj/F86ERFtbTDhuFErKWnH+LT1O0cKy5toB0eu5ccl
EscUF8dhs1hwaGjGftV3WCEG8Uchd3chY+QvKl33AhriB652TNAAnTToMkDkychYY2Mb6Kr1OI8r
fyxSCBJQcDaqFGQt1WYVJZ1vharQeQedTEicKYK5zrbYQDmgAfSozYOv+1ZdcPD4gV3Qh5kyGKyQ
yzHR0AiOHnPTa1vw9aGLnkMnk4jgRKIN6f2Zf5baCcNTkRau2dybqiFKlg4azyqVuJYZjdW4R1z1
dBcRcnW6uz1KMiEIRXTLkDxP1Kle9sC5HbELIUV72AA4byMaRruu+WWivNqGoAKSRbokPZuhKDCP
JGINxuyUbfFFI3BjfdRwM0RlopMmgoE5aMB+W31tf9e1guFzwGAmis9REVo/Ygb62Jy0cPdCRh1Q
AcgyzKh1aSKyaMXIDD0SQ/QNyJ9VsfaY3Y5yKspwYfSUS9acgSZyOm9x0ilxi2IVm89A96+VNa3j
1j8HCDB4ZGw5A+2r+9rMUQKZuoo8TWy4mJldHnw9Py8vKHqaxSunNOM545f5b/VZSVmzsenq2JZr
GaSw9c58hCDtfMM79qZiFS+C0y//PIr5xQR+1ii2QGz2C/BSuPD5iQKdXXRQS7Z43m5THjSR9QkJ
0oV+Vz5Zsm0VFs8lmYRpvT/rWly1XUSjclbTK5XkCFAWttCjxpPhmVBON/25cL2Vs4RcL4uFgly5
s+obTyjHdhVX8n/2kyq9kyISZLbXyx+M4Spwe+lecQx8xNnSi9+Qf8i1VIcc5uZOkqhr4twvEkyd
ioiKyxOJLebzvUad8zmRHBwMY8WsGnGu7/qflGLORoh42FIIp0Q4ec6y5UFxoqbidbWY/4ugZdR8
zzm33HE6kPzzx7xBdUBMiuslzg/Fl2bwreuP6ONN7gSWuIipCVNb5u6Iq2UAmUX3xYxPz2L4ITc1
BEcQwfZhpkP17VUW2/XHEHyH1jJsJn6vC5tYi5xs/c99AL6HxxuF8EhETSjE5LWfsKHLDjvmpa5G
ZWtsTJZXGgJj04MiRhyhwQTPnQGcPZSqnwFKXGd1mHcA6hZGGp77s0JLRs8OjX/9mhNfSTBTRj90
ZivwTsogofP1EsFIV5t4BqenRmsGpZN26JMHs+Adcla686R3rAUCIlgfkmS/M/rUQxF6rMGazr04
5ddK4c5tSYYUvhfazJYU0zQd2iz9O3SLQyOp6LHGf2rpCnSr1mf7VXfqLftrlyuF2/AaSTjPkRhc
w1pQCOTUtz83tGhNVPBkr60zbC+4YlPVH8DTl9N/LhzWteoEk24vmO9Ri3RptfV4GI/f/u48cqmn
9cu4iL12NhcN3deZplAR7ndvT7zZWN630NjTacbXnkZs071vz/SEUB1fV8rxYhSvgeFrmcFnZfbl
FAjWOtaH1tjxGdhb1FpPiQNS6Nut2IQOzoakKBJRSjNmloLLF0OoleEK65M4m8c29uoRVx35oBrT
FVJLG+4muJnW+CJzcBhavG2lveOrtgOY8pQ+A7n4YZNC54+KoxUU26aNH2ivmkpMf+6It4TyXyql
XfkDxqTZ5pE8O4k4rBUoo8DksHyXsyqLfzUnfg5ypFtr08yKB+pukwfzfZlgQvWcYi2kpBAu7mgZ
HhnJ6QQ4tjtPqc+IDApvc5lVe28nmllE6cHDQT97leNoPTNHcaMAluHX7a8Nf+SMwDvO7oQYwUFk
ffbNam5USlIZnXZs6hmXs7xyqO9Sa3pwHIbhqeB9yzidrgOpbnMDJutAz9d5uTkbHjWSe+qhfL2h
fBFgAcHSi1mqgCqbvcgyh1Den0U+lUfALpUpMNUGRlkn5zn7au7GW+beOUlKzNkTNGO2IZeXkIbZ
D4kzqaKLKA0j9brRjsnJK7WBNrs7iOYuxJyu1MUXLGPXXq+WGbODFKysfOhc3I7Cri1uBf1tSSHY
yofGqy2Mj6DSEab2+Y97pur5zIs+tqqwKBXxB7Vhh/oQm6br7c3SuMTo8OcE/eTOYJvc+nXPYaxH
Ujhky1sDjxiJXK3WxuyXOtiRE1bb/VN3m/ZENs+j3IuESEL81q/qOTqFudgRKbVkGmjCYDW/+YRw
L6yw/lFLAtQmPB/apjNLyeZFrStDjebFtq0D7FFEj9sH2kHLLedWaZ/YakHkjQwsDv6NVD6S3OwW
RzZ9hPaxR0PQJ7pj+bjTF1NjPWJI6Mea6T2ekt3Ygx1QSO8VknnLv8wouoxCggzauyzOndx2GJPh
n2OVW91/aoUtAWi291JvWHXLpx3W5OZbsJhtTdQC9TuWrxXJYL+9YvG8iHC4PGxBQJm/GILi2gB0
8eaMjywH4V8/5u0q+wjun1LoSbI4pDSuIlD6nSCaJoizN+53t3XHVDajWUSOLHmwilY0tgdBFnmf
vrU7LVFXOxF9KD2D88Pl/X2hPolz4Mw2Qu9hTwI3gGZlmjMOfFAcGlo7AmaOuTqI8YeCf8xTxVJ4
NGjEqYmvJwKInMRDLQSovOs/Gq/DWq5Ag41/gpsnVTzoqwqMSrlgbHpz+vnMKOYPlgR3MqbPqQ3K
oYaQXQvS7nhtg69RmGprQXwLhmu4la9BWXnOj19RiLVjroeyFZ5kNkixLAxTdzqlImrzopWAJmav
ONbVli2An8z/dAyKT2yR+mfvv43m8mEO+Ike4PmXyLMS7gCYWmYhwgZrigeMRctqj9gljHN1hDQq
bgunWvGsX8HXqax8eIeR48Mlcp6HGK7TsWEfWyY5d+9OaJ9FP6VemLX7WgoUmD6ej11tXWK5D/sD
5OMM+4jD/mZcgu4nrPJv96E/Y1DHEl8Gdqoew5SmiLtIpXjzUuYrMAcm9GArC6K2tOx7FYoonPRA
UDAOJswiGCr4ZAVA0zcn+wrWEJa5XBEyoO7qnLTdSNqPDLWE2W/M0FS1nh44XX6LCUXwxSmcJ2fG
v0RuTPs+BdzfoaVe6dk5BmVjf9yoHM+2dmprYy289NpQQuRjrJd3tn05HOWWD2og9U2GvjTE0yrT
fgiUtTq9yAu30zHonGcJ0Mfm33CeCnqkGP92rMhoVBrj65YMrhk79ypYUzThOLaCWD8AXamsf0op
RV8njB2gG6QmLZWXUuqTwrE9cOKXsK3bRjxGhrqEDaU0l8wcWbcMsUdAMxWf9enMrmvjAipRMCb5
VHadb6MQw9/groqqrJDSxDx3pl4J6o983t5K7XN02O5EtXTyniRsgecIdnvdqHz9RTvtZKT4XaA5
ZRprcpGb5Onfnq9BCMiJIQ3JMWP3yFIyrQ+2dwwqpLrVEXR5QPawB/nxZmr5wpNjyN92tSAM5Pif
gVsbQ/sg4l6/VzcUFtQzzSyhQjfrUnuo6DrUUPS0I8CKX7+VdeyVn5mdJ7wh34XOJ6XnjbMapiUM
4t/sKfhZhAhW96hmVYUfup65MIlwdamqCd70wKwq2vNGFlzikGP69Xr2rdMTL/IzASFtwYhKODh4
b7hdm1iK+SfqrMwesQmgfAyfLLeXK4luClzCl2zbPcc5CLL+rBf+x+d+aLNYRcIg9cX+aR7MnEEp
F2Ei+gMplUke0VpI1GuFO+zpXHDkIZKKHgg65zwX0fxhoJAfpnt/fI3neejbeVOFODiUG58Lgh6z
RRexRTms4XLj9jTYenNJWKowA5wE9LskZe6kUR1mN0keLHdVGzcW6A==
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
