/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 303744)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvl0D/RJBgnBBfFHJkTUlMQQqwBE4i56aP78bgrlGzyskUNWBOunC9pjig
Vg71OsH6KbgFah3qmk9fxLeUxC5lWFu3PbhTdTAOsgYfEM61LM8Y3t9l+yYKBHcJ558G3oyhu9bx
IajXyo6o5nLG2fYedjjtyGxTLvnP+P6SuveToUTnlfpEmhXYySo0MSSYJfww/v3A+gDkLJh92HW0
/pSaB1Rdj+T5oZ12Z6zVIRq8dR/qcF6pReAbLdR9S8qbWH2eCeKk2mnYX8dIPspgRiy+YCPsD7sg
g5xZWuNuF/cXdNM3GPsNi9RHPqQwiOQgTJII/3Ru9LFpB6A3eXhmtXwNlBr1RrNncF6GvUqvfxiM
G/3CnFrbK2xpXSUuo9k78Y+RBkdrHqYnw7+VTBM7/WXIwpAD51S83hnW039aqeZFE3UxVjlwivD5
ckZ3MvS0aA0GpwTW+9U9UFyWNOq5VopLPbCvg2ZgTuBoKbp/xC/r20tW9zmtqDCbr54SvQBm4RwZ
FrBQgaPo1kS03rbYZq1OLnrMTnad1S/75QHAMJsZ8BP/xASB5wlj0xxZwARXMxC/M2fLIsEKEk+T
OMLPq8AVRHhucuCcXI+Em6L88kjTYkJYxtX45Y5SOSBTdeYUp9jDBogEYcgumRvXrdvJeTxz8ajy
2HaVGw7Oia+qdwajDxAtNzpFMW0wFTgpqznSY+WZ98zOBIKEj/kQqJjyBr6+mxqqjASPo8u/TQf8
rirnfKzPdu9bFS2qPE5Bjg9ZacgjD7a2SZBwSgeE1ahbWyYlzHfw0xvoGM79kyqiznNY9/7F0Trd
kIShv2GvHfmCQB5zboxcJIz6idoWS1dv0yC7ZO+e+LIIqvzmmC+THLbVsFUMo/8p0rS5BCguysop
p8rBjAnz3kAxzfPwHxUT0lWfColS1GV6/v0pMzFENd4i6jF0BwSR6Mfw56Yzcv2dLB5oucgm2UOz
n5ApNBvhxyP9SFyUC4DISPLa1twFGz6pwK0g+cQFTyDc6L7AlFEHfCeh/dpN5cvxxahzcvGxqBl2
zzHe9rONh7OqNMnEthFT2Qvynk9SjSrhZ0Cc8LGnUl+ZpX5Ih7OwhVHHVPNMEiXhasyI2D4q+uqg
RQNMI3jpfHDecVqHE8vJ85IwBroRXI0MBgWmFMVjSRDXGhgKMIZw3/lt0OSVqFIySP4lflKZt2y0
pDK/3HkIcJa6Es4MDM+UXCNn3AhrhXsDFqMYoj7RQvbpbzEaL5jczmCPpoCaALaJ610+YZAde7k3
YasxfxbIio7oLwzAESVKmw52soA43CI3ZSBxP7QaPmPhUKKXmv6p6eCovBvgsC/MRIljDYDPz8Q2
2iQ2OqjREPpIa2hvigm35poRQFD+udgkWKTuhof0k1le7lD16MfD1TW5W5VhbbbXu/cTjc6AGpdv
384diDNlvxSn7JNKf71PY2UcptW87L+kZboMjBzwYERoW5sPQ+YeoQoQtFSEBWSpy6zeSP8rrjN8
C0D33pjzdXyloQNpd2+Lqipl8gTE6FVf9X+18/+88YsfFTFq7JLIL0jY6pupgBnQIYOzmCZPCNm7
4POchJkFB7GYMizmPA+gsLY4Kr5JoSb+d70w8I/niWuHvjyfv9Xuc1hNmWLDNkmZYxpi5KohGWYG
8L+eqe99Bw637i0v386HbKsPoUndcPaKjtdeSyCBoFqIzuCpVR9xr8uwFkmxoZpppafj3KN7U0Kv
xvdbdsW1BFi7g1Rc+MrEuwq7xqfc1mTNJMmFnEXvp9BNEFCwAq+qapJYlS/8FXHbMlq5+CUcY9A7
Nri4BrPPasOoqBH3/VsoW1ruSSfk06nXaJv1qyFfoLZihM6lYFCiqkxsweKJpknOqsowA5SkqvbX
d/j65JC+PHdlFrUat51cCx0WwegRvAIdSffDXMvyxJd/2yBQZtdeBUKdrRZmqm4AaOl9f3Y9JzOQ
E6+Op2YAI6O6eIIuUxJLYn0A4PmfRdWXH+huZD6AErlOmo/Tpjg8nZzPtPedoCaxiCgneutUxKe8
c7K9DGmnl5E3i51eTolqOXRAYZt/KWmyBa/dA6jm6ufiX9yUTR43GfC6fvWCqKgYhn+6CnAQmCfF
NBJF3TTkekBESZRdOUfKiHQ9mEdQH0WidcRKPG4oXjIlsdlafP71F/q1v0ILi9sDYZrTacDKUFu1
Ip+hV4ualROiwndGtX4tI9CdMEzZ4H14fNPWrpPewJPJlQdTsgS+vW5686TP6MI8TT4qUDh3WhA5
oL7u15rKSEXSzkkzPXOTzoM6ETV/mJ6vSkhd1BIOtUW4LYQ1vgassL9Q0Xz/HKuksaW+ZBFAf7j9
n2NMf9LIFS2qTs9G8zqd1OHjqWwfQTLXQ5Ku9FV6d7Xvu+XkI2c1lbgvx4c03StXKRLLcm6XtsKj
8skTjVjJppAVKx9d3W37CbTV8bEPyefQxafpfxC74dGszwLOMObzXgSFnLLuwFmLfVunI/rlr2tE
nVdeLfzv0oLahXZrtBCtEq4BfgOghZtga6e0iPkh/KtlOwojZGRSYOikpYp3Dzaq5M/5fJ4rEyD+
7e5qxA3XxOrhhOjJyfv4miI56gBRbT0ZxzYZXtMjkKm5vAcXBPfefj0kdXfhasAXW1riH5wCc/LQ
/5Bf8Ul2B6b5+WUk2jB2zoatcwy4T3nLWEsM4b5MTFhsQP06h0dc++8w+zxVp7Ig9M9n1G0+0NVh
MGjiQTaRh9uxgxwhbGDRF3RA9Mwq+wkD4Hi9bpUYPnT8WFw/GY/3GUYFQJxgB1k3fcv/8V9dgOTu
koevsksp4uI3FNaDqNbjqSvz/RJLUI3kRhvPolnrr8vOrNJIOOtZMb1DiggS3r0+aBswnLzmbYsK
9w0G+51KWF/KJThhwctMj88Sc/lwgjM8PqQktGnGCbcmObj0FM87KXAtR99WKLwFzDo7GW3XxMRY
Xs5mCYJPu2Ox04IhdiRjoIbPwK4yrFlXOP+6NniscwkIZcdSz83jmvC4t9w3jh34CMSaQk4feYq9
e+8vw/sY9Cp5ad49Zel+wdQ4B5s6shwmK2ZkV0kxUaemWCd6aY0yi1nohe7cwGHTSady4y96KpxX
UjvN8vjlJNTVRFuCL6Yi1irHOUK2BZJcNcam4OK0PCdustozcj9i7o3jUCnkA3KESGUYZ3x3Q9wA
RIBMm6ZA9gakrcWJvntQJcwUm3swVyuuazfE4Rv5B6o1kjwgheBmj/gbrTUjTBFVfLWJUMEk5ufE
8+QhwK1jNxZlm8NTKnpI8rZ6vrUNAhBFaRLGf+3WpZiuPRimrxDeLm/0XVrfs8Qf4J6LvdRfN1Ev
akVAop/gDsCFdYqRkd2/PG44r29USgZd38hvHk1SN7i28/NaDturdSD2uRIALa6VN/DkAAYOlYK2
amJ1YZUQuuphOSW/BL3bBX0BXaHzQBd/I1A7F6bvWguV8IXUb0R4WfkK9Y0XE0CFthIK1SiY79NP
Jk3eIfwbijBiYmKXj1xJcvMxygDf2FcCf07QR0UErG7Nz+shOYGrLhzsYxDGam0lLucn63cFshPL
yTP59Ocn23kwzdKDNdV8DKhD/oL+dTvWg1Gv7DZAP+H4fiT+i8W5GEyoiEvUNoWpz/xCQRFFZrag
L8asFy0bwBXkpTCLZnhq/80TXdbA+QZEFWlc7XSjC74dD49uwiADijV+MOFE0n4yDjLjiMFdGR5d
uOsCzB7kmPtaJXbRh72WkdEOBbymdvJh5ELhIsefM2kP9ZjqEaAXsHT0pweO7KsqFCDyLhd6kFtA
OU5TYVCk2aqU1OB0r8NUm3rEkF/B5QxqX9pSn5KY/CDnypN+eh3nB/rYD10kXVWc9xrde+Zq755o
kHpQeGN81mRw8qKO6rr3sFngbLMzUTvSH38LjAcMmCXQvR7wJiY0Hlpen8TuRTqe/2gYDE/3yLYH
dF1k+AgVitD0+WIoxUmM3S4m7QAvCWlVe55zvFDLYMqqgX5fzfdB16hMaWUfqxfnseLkd1H4L5PM
Km7BAZ7jkJfBX9TVvmuMYCed6Oi9GIvtOBqamw21v+CDPJkIQrzmWTOr7nIJnCBUu6JV7UyVlCwR
prtVi5sbZ14NGw2AIguq5eKlPuPPlD7yOGeS7LvfYJrDNwlomK7ViAhLY6rnGpHqzRxZoJDGvwIo
4zEguQ+P2jVAjTkAnBrnZ5IooGmKXMfvy9ay5G5RxmOMA2vcnPSk6cwNSIewD5vKsEaJTH2DokUY
llzDlPARVihkbLQLysjeAerjmTHFKdilZxkltRkIPpaC/q6a1SbkuwzTXsYkmnwdqpIcLsrEvqW5
hary0es/q+XbRbjDOWB/ESQEI8CjGiXY6791O1hW0YJK82sq24Rb69egdzUQUw0SPYAr5TLyxzW8
Ov+AOgIC9Rg0Rm98BOLzMbBZv0tbOMV3Nl65HM3zmLZokY+pCqkKLeZPJIvbTOhTnhhzkFw4Yz3J
4eoEtXI9IEGpVPhac4EgB5/QlDW+CVkXFKPhxbIuMYDUpedC0poVshvsBrxvQdYaWGoDMDN+JYGy
NOq5fLg/qQ6I2LycuG2tXDWg+jM+83Dz3Unl13xkoPOFsYCHAZEA7sdxq/zk/ihuhIJiIdfTSEOH
AN6yIs5qRxfSJVRL6MaWwuPA42UelAPSo1//EmV3y1EbBHz3BIkmoDrjmXxjPCFEatUw5eC2EwUH
/b5Khr+nfIrXy9qihGGMMzyTyAVnRdm0TBtekb38kW77jdfo7+OE3GXF505jGIHbE6ZV8vq/EJZS
rysfhNVqx8zZPrTBoMvSTgqpFAa8bpgxNnCrXKrwAsjzpBQHKtKaAsCR+Dk47DuZFJTkMlyvYHxl
X3xmJziJi7Tc2WWj68XLbeKWqlNT1HupbRc821DPdfuEwX2kwhanHwCyoRQwsZ5Cf9ns63ee1eJE
BU/cg5tR4/f1m0vLgj7i+yGHcs0XOIAZRfeit1IUckOuKoa06eP8W1PmuqWeg/lr0QrzDyPtyolP
PhqVnHA75zc+MSjma6aOpqADWR8UWsQX3e+SKJPbyJu8v2PzwxeoMArSAsEBi3TTlwRF9o8AGIOn
G3TcHmNY8bJdFsvSJVfX/3MRaMZDvPtzh30uasOoE8egqOinix1K99ZPnUifafCt9FfGr4ayhuJN
k8VQUSBcQm1MuGXSp8ueWkqDOuwItef/qBewe3j/7Wo4cT5fIWQT/UlV5iCJxsI8rXF4Bauih0ww
tmkmW1zrF4iGepaSuSSG8wiou9+OKwpZLSc4MJxD1iP55FqeHXl8tbdiZ5KocsqIt8suakzuq4fJ
gAFalTxS7SJhFn3xAgv66gx77IjpqlsFlhFA2RP0y0ybIve59E0J86csdoySh+7OaZFTp2Fm+3pm
2hnptuVJDyC6XCzZufidvMq09KRL6iYgReBMx5eEb1DH73IKMcVP+tdJEHk6zl9Byz3h50Rp2TDZ
LrCK2VS9B19Y6+3FUP0JcBi09lvAkZ2pQ03LpbD+m51ohFPom2e8iamEI/u2lVRHko/To8erAfW4
fTwNNP/zZFbR++cd2pk66HXoD8s/w8ySCRnXym0h93/sVI3seBPMLFUcZSVUIPC53kMvRRejWd78
LISBNtDXXAWeDfDfiNsf9qw6bMJUFQK9qtRYNAngNBtkxA6TIkfLfJhZGMSZEbOA3DeIc2bOZgKI
+IZTQ+7SHfHcH/H9FUF9toV7r/pof+4otTb2EfDPW7JLbFkTxoGHJNWFSckyKIS/rUJrYdKs3ZCV
+syTxg7bbN/86QImytQh+G1bxSeB8ilp4F+4b9BQQU2Pbpkq7IUG4WmXY3RIg/jZfBArJXb2/nh8
jw/TqH/okpg9OVTuJ+amUXDp7KgoyP1Gu+GeVUi/CO0PY1reiHPeg5H8431CYXeIvE1Yrug07rFE
rRn9j5DdHQoTAyiKqDNsvGU3C7SjdBTw8BOQNJ9co3liaBoC3rVnMxeSQE/dIqAc/wQUq1RnWVqM
noWAeKdrvOsu2mfV6Z7P9SuDMVh/t6v+eKZ4+afbvhd7+DiG+7akmrcfMZlQTNDYoPgWYYXhY0NN
bDNmovIOIX5EqwULUzp/lhgsmo3FyUy4bnksJHIbRVhQ10dlN4iN5LgK0hYh0LRrmbxby57/WEv2
lvYm11+ds2t5VV9yuyLOc8q9FWIFahqIv5YACofK3UYdFKqiBg8xDGi+M8w/2pKl83rwX0SdZlsU
+VeExTdxHw7vUDIY+8ZeOouEFWYia1TN4idGgv2qn45AAGuSAdQaSeetHWOHsynRYWogQ5lXNNbQ
N/ip9ohzwu5YzMXrwbxjJG7/nBuFo6l+qD/fa7R8gcVcFgpfddSDl5NA6FKujt18KuSIYX5aJ7PY
gkdwO9uhiedU8SEm45+gB3IwhYO/uR+ocA8fU5Sxh5kZMkXzg8WpSrplSGjtzX4AUIHUZl42ZFOH
ERS/E0eDT9qwIJV5Q6GgMmeQU/CzC/qd5QtvJXI50OrYPq4KhoynPnNGNd62ygYALbyPe2zSxG2Z
T30gYj0XKGIV+igUMschX0ZAPulMMx5UbWS1FPGfPbvsOuJ7HAxBfvcxNLYPrHuZuRJ7ZEauXYD9
EjSX1WiHlcecUHsEGM7el7TLJD5cv7mlxP1fdaExz+gBPwSuDpgocYG7xrsXIn/lAEkPc7i8mC0c
Cy8utyenhJT3ula+T8PL0c0FhD/DU2yYMLtuOw4egN4s5jjQgpEVph4CanFEyxC+AwpmSvUI+F2o
YcE315pylneTgqFjlR+itp8KFCCgYYnHKyUrB1Tz/PRnO2FHJV5Ll/jEaZj4nBjrx8M96Y9FKVNB
3kveN8fOmk4iYNCTl2FDCDQcMmr9Mnv8INWcCg1DlIOWMOfYWRnuLznsU/rEVYoKug9ou7177RhL
BdKMtEtS/wHrUT6bfbuPyBPl7b98FpS52c7RmvVhfDzNhikvWGm6ZFxYrHT0mWs6Wv81jUxQW3ah
UNk0CoCB0izjkbRD33QnA3pAjNhA9bGNmHUAJvCYWFOI4RWi5BLks1/hRl2GuxNn5v+1a7r7L/ED
4KnZn7s8IWFb5bds3dFrVuVG2yFo6ZyLezdnAxeDJmyNeFETJZSrD0pGYixWstKneA2LJIokUqb9
SBH83rdmeREb38HA8z9yiRHUHbFPVFXLqA3HPnmfgN5EJdfdlG6ERe31UzD/UOhuuM6CKqqC6paU
magFXNERK70xTqBAptrOg8Nn9YbMrun8KOd1rJPn+PO/4Ltqeid4wGUytqe9VzKZVU1o3R+ROTI6
FmEvItUud+wRlNJgbOEDrmSUauDuTINGmreLGmCV9sSZTbVTpFeDa9L22/BvmE3M8/lPOr8XEFiK
sbyfA8/+9GWyc3mz7QoFuSUuJv31iwMPEFdV6bSMOq18YH/k0f/3xF+e9bCiO0nk7IJiPJ89lzKH
uYLGmU8LykYD2Mow+yjOsxupcb43cNHNnwgRLKnpl9J0h/7/FpKPXdQ6Il1nswpctFGwx2qr5RIc
MtO67XvOfuNh2XPwf7kYhvLLmdJANB9Ix8u8QZ0ux6QL99iljRjlvu16HTt4A51RCJfpczOFIq+7
75f7hCCwE0qZvPiAF7k2amLJqPZL3If6ullQbAuPqpTYW9zf892B8mucwaT7WPikDVBy/A4fW2+P
oR4r80h67rJT/zwQNdh7lniJG68uhnaYXsoUSOczVQ5f1o6kThOvPP2nyXGgfOUhGCfGm1CuNTb9
8q9cMPCUr2YiCk/HfFK5LiCddQeXE6fPieqv21SpZA47wVsWBADLrFMFH2pL2gK/hA1D+OWhTyh4
Zv3a2zPO3NH8ZA8Di0VNZC6iWDifYkjqKhJEmbhthc9QFv9g5YGiQUtyQlyCEAa7CeRR4x3fFMVs
MjcstucgyutFtKclMdiUGOjyAVsfulNZlAlW+P2F9zLfXiIsRqh7xu8DMq+fQop9a6vxoCnDxxwc
IfQw3KD2wIGT/s3hTFRf/3PAekduzrphYYsx/ttlyCZpSYJ8/PdH2b1eNhNKgWtdjBiuGZcF7vbm
eh4Dfe89RiaOdtdrxe1gRZ6z/dzJPzsDAmKlOSD4x7anIVR3Qbhf+qjd8ycmpcUSctyvxO8YcbQS
AosrmXAME4CHwsizNUnP4Rh+9cD7ej57cK7RD7IrvLLY8BhjvdWT6sqCP/wXRwyJL6E2YdNCTidP
MaDdU8wwxwc7YEJwFcDE/qQLQqCjPk/1UqFk268WJw1TTbDb8Y4xGoQidbRuSk98eURS7WqGDY+P
IBYdP2lsJU9GkU0K28kOVWBuBLawiagO4nU/+m6kLAWMn7O/PX7H65ePKrmIUmk27i6VTR3uoP68
/TiKvI+ltnh3oOBKZdPXEGcp06GNSuq7j+9L+9Bwir1PUcFVxg5JIO++6NOdG1w6jSUDGGwZnd9G
oZxSiYhndzI+pUNZVkyc1NIyxe+uNDe7hMsBb6JkOZUzMZai+S70tjlLt13gUrYqu3n7W1Y8pBLs
Ubv/MgUR41mS9q1ECruXzgnQZ9njL2Ht0pU5ur/8WZ+SXoWXbID0FJMmFcDOJOVkuBVJ9WfoYU9O
ObEbNBFHOo5VsGexxxpI51KxHHp+A8RG50L52w1IIaBxpb1D3PKNvad0ip4bjKhk+UUM5l4uGcoa
9l2tY7cxERxCT6BsijpB+VlqSVF7v1K0HnCFH1eQTGqcKo9RvgmKIAWOKuhYjnGsFXKV3Fq5cumF
cqrhW4tLGG7kyfzyeJ+xZHrANWxeiFdwPhoCReXMYq/7HsqoTQFpiiwEAYjnljYSDnbKlWiYzFpL
HLWD+HXI3aU7DCrOn1m2Sfxo91cEycXc+IjYHJsZPzPkXB6A1jcssSgq9iEgvwxUOIzdjAoPtjlb
fvPbtjpZUL1A5IQ57djgxxFtS0lR31Dz4sc8Rd3vnjTeWqfOAz7Vtwz+3KyX2C82dLT1Oy0dQrNF
eii5dU++TXDppurgklVXf7nfGyl+bN+UjiJ700ETU/N/BTduLYqrl6tpJXYnYyUR0gLqD7/mOJLU
qS06J3qCa/rZdBPdfmiOGMa0pj/Dsm9r2hkEbb0tnyfOK7gAcC/lm//gNceujac2BcITOV3NmOkd
4Z50NFKPy5BKl/gSGGJamWopRR9yGTvdCyGS/cZyDMycfoeBBAhavLOHB4L434468cweLbBKui37
ll888o3PsAcPAc0ifZR5GIWPhNni122WfIP85m051giLy0CbSQUj8zzEOwRgvEGNBudrnLDKUrGZ
yix6yZZDavd1j+igH4HHMWKPiRpj/Jp2CAfBw3pNu+vbypdL6y8tI9d5dvtHCPZSjlwPGth+cW0Z
u2NVK9KG/qOVJckZnZCo2ljEb7fqIVV/FJDNg7bhR8vnA3yHtrJW1XZ6XhXcGT1rNU0rMolHS4A4
tMs+ObzWbdxpK66k6cXxhloLJpNiVgf7418ZFm441mnW6uGYO4h9346z6PGCOEl5kKQFpXnnDkHu
ffxtykJAmgiEpzExMEUhTxYaO64G2AfhQJcpVNocfGDeTBnjHVlX4iDvM3iCaM47lxbpbhoVBOdq
8MG/Wrgrd+Z9jG/iubr+InvhXtqgD3rJwyHwtL6fHAsMwjBo5LIxZxMJH6tVpUqzqQbEUnex2oaU
MsfH2Yfh8Fw7OUFS4Rqgj9cP69OeAbx27DY5tGGn9XfmTfE2Y3TMXGAp4cjPbRU1tyFMx207GpAE
xGTiOO/KTO5Hnl4yIZm9XV0X+gR7NVOb9/CL6Hk2wwpd3KOKM2jRPqjJ7cU7ggpUMpu/0OByStGI
MXov8dJ3EDyHuSZs9gUcMczYvF0WUN2CT0935bf1O5VjCeQuwizTLeIeLncbb31j0XUJupIQmK9c
HWGxbAD18tNqEvXmyEuHsJ/YO4cPr+LQynQ/31tG52mgxXoMLYPfCaA5JiMoQ3GXtWnCy7Kc0lD1
uSvhui2o2tnnOdJR/GikWPs2SimgfzUmMZxK58u24x8L6UFycw/uZfkV8MIqej73hFq9lrwPXcD7
WwCn/J8SrvJkIFQb+PaLW2sahi63+KW28tHEnSc8Xtt1awV1gzFX/AGCFJsh9Y7OzzSeUpBlxHy0
0ujif6MDkBB3obA7xbxwoIVMov/Xki6dm7JSPjhT9Rw+j6EiTtg0ZtzOd6dLmLK9GVCJAZri1kGe
GWg5veO5x45UUIjkg9gdtSKbiwOPlStsJYAZOXWhcMmE7nupC24SYqqwPT72r52muDD1X5rqCHlz
rM2u3yfIbxwu/GoTSwHzpHrWkoBv6AO4rVWDBtfDqB+BJEqk6T4y6NFhOry4KG9ekHTc+pIY4Guz
t9VK5dgasI/CBCBxHxq69YZS1biVIDQPbpQtEIkk7J4cFfVqQXv6x8ltHP8IfRJWRmg7vIocVtch
0mKi6stzXi2e07vC1V2L0Zt3g0ESIzGPsfeMnYM08nw4qcLW7ZYRyaj+uKFboKhnmWF1/A9sW1qk
5WLjm/ZuONNAaO5WipCoHEwhWpsJNmSZ/lMu+NoFXoKs8jLi/0XDnRgb7N0QHMGyqpgxQUQJV857
vPFMSSZPPiF6/IyvpT25Vopnhu96vRXcbeLJwkBjOAx6x7Vvf6slnxWLJOOsn36v5rwsoOM8iIT+
JRypEQl3NelGr7z6NObJVbWuBm7rLYt8WaZmSqrd+DcZYlRh5xHfSVUG43XNYFXpKv6IGv2xYqdV
sesR4RHPbED5SKr5g9F74lZyA5iIurn5qAxJWB9Lf+fzz6XJp+ZSbWTuXgC3O5wpRMa0peVcc8d+
bkfGiMMB28PYOWDFhSVAbE4Bt8gg8UOWM11siA/GI149iq8nt7GJPgwREzVnIQ49/LHGTAMWgrXo
iojUa0lcGiju3PEmtmP/NDE69Hbr0ihadSkbfxCy65r+igse5vX10U+N1G6GqoQeIgG3+DR/If8m
SMc8DpRIgANhcOMCDsMgxSBOfFem4Qfy+niM47jrmslXa+k2mFC1YaxTX2NEY2oInQALvHRnbChs
F6UwUh+nrg0x9eAHXIRadhUchixwfAx8y2uPMU58EksrnoJvA+1pTBj2kPIC133HEgk0dDme7ZL2
ENNU3n/hI3G+Dabzjx81pZs70hDTGpdCcA67qwJ8K+z4mOb3YnrTaQAwsHZoOSdtIWBt7JdqKPIh
4F4+hUpqzl3l493XmIAZhNRYOXNvjNNWC2PXI3s3AdPjrmV91FfXmHHxm3LG/RF7U7VXhe41CB8e
qgNRo7yPtCIYuOrZI0oF0678LN9yxKc/GEhRlQD/OyfmKov2jY1cooZz3JySutx9ZnvrUbzTYSnQ
ZPRDdQ47Xep+TU9Mp+L3zHNM4CH/RlGG9MqdK/ayraR1TEuBewQAYGohu49hk5+EorEEx+B2HRbc
Ik9Uho96qAJoS1/tPSGOCOw8kTz0gzcCPbJCtr6DFNG6ZpF/vtL3XV6nrxHBixBMGw3YrmytQeVW
Qw4HWvjrbkMmbOLsXNjCsgDaPzg7NzVJ3kIv9mfAqUbgZvZVkt/4uNiRkuxgQeCam6ggFz5DTxJQ
EeHa4YXQf/M1JHNBMp8sG4dZSC/1ESyAcB+4IgZPwMwAtLYv/ETRTScGXMF9mfUs0Ku9BYpqR1OE
yvRXWThzffGb+kALKxrctgIVriCJgCdd9GSamMtuiVqe6oRxisJCK09sqf4w3Bl5z27reMjmgs8U
rdyi8q2IDGSgE9OTYzM40iwaG6BzRkhUjGoVWyne92nlD9sVc03DxcdsoGGilxhhhEC0JM7NfgTZ
b3PkbauRbnlzzz/aEq17eM8Wd1e8m2OTw2VjFjKDYQnczcj8Z4+PHIQB8+gSSQFivgG9JOFcmlkx
EF19ZJ9W9p5K/EsgMllGryGNO/AxkGoDuXcw0eNtyujU0q5IprkG7ugInzMOWL08f7LStOGMc9gO
XkurJ2U0cKjmX5llFXHOuA9i6HN/vPArTUed50nGSEnOfZpMer8/xkgfgv0Ne+vsRublAo+FO8Zh
dkFNSfsaon4ePZz656ecVXKIlj0qLwXHSzl3AHy4jQ//dghuK4sSm7TQydIwtRERDuC2mFTgXSDj
RD1ZqX/ydWE2HjLEeTGLMH2XJzem9E/XeTrPKUXzYkvbl95NDOvHgEJfC9/v5d96F4aqqMqOiJgz
jU57L48oY16LWMYUSN4uWjkG5AVzDMB2sIK3/FMxoYSU/mqsBsd5/Roi+/vDF7MYpUsBNJ1iScRg
evY9KRPAyWW1Ua3FDowaEBECA2jZ33x/h4Orz1gc+uGlMTfe2wz7jbktX80zPWOfz4qZfNjpSIuX
lCtVQs9mvDGZBF/I3b8xHSCM8oKqZuQukwRa5DVO9IiKvsUrlUL27eV4I6MGuQrsZQZqzApjyPIl
4bEcB8GSS2+p5CiApKF0xWcvpaN9EKQVUD8IvKFEgZlvkYWg7XYRGanJ75MgdMFwU+uOAfcuDJIZ
pbmjG33vKEHsf2bVzjM6tA0fmjpByUh3lfbUbbVhuG+X50l54AT6p6Dj+RVb96BXqxoy3Cefcq6Y
9HgLNAPaovgNiXCKNDFeLeQU0w19MVIfFqio9kZdVvGNQ566h98n7hEJjI785Uhs5bIxAWfxCI2Z
1POOUUYJCqzQSXfw3BcSSrZaM3+ielx8VjOVmaCb+hVTG8GlA+7UACSQJ8W7Ag9i7m84abYdRFTq
c0bDdhQfBKxcTKN8+FXYPFErx4AGFGrmVSm0HvimbXfpv4DAJKIKheHQFw4h1fzfaDXBRDjYZEI3
a0tx/HP1S5rZyR5ghWJSBy0mI1RUQuVw6+cpIr1OPz/Xh4b1x9yNlqfqJx32XR6ze749H7hm2HpU
wAow3HGsVUkhZ/8La2ohbqzFKm/m8uSLBK7EvlSFkNOUg9mARCH5Q2Kr3EwRUoBgXTWYphKEDDTV
5pmAWrhQqkSJws+ca/SPHDAxWLhA+EFmi/ndL1OA7HrJHv7cev8/CPi1uN+u+nUMKxovTKPyXoqC
/ue99iy6JW+EPc3WhZ77sqF3MV8HOjkJ+tDzQsPWIJPD2ENoAEFkEBGEjPHogoXBSeRXAboDTLZX
0ZV/M/pVFn/1a0vKlbP+1swZCewViWkkm+izZA2jIF5bhUX9vv8VGXofQWM+r6H7iqPCaBPkPxS/
fY/lV2q3YGZZIyo/w9yr+7URIMOhoLspipoIun00FtdURo7wZ9upwxJvelGe5KjSCZ2LDPVwLLLj
G9OnJIuss0LLIY08/1ONyUegFcgTenTuDInmEG4bCf6a7yNkZvy/tvJXMCAo3h80rDkpDxK44/Eq
gQhixMqQ/VRl13Su7vKD4Vuotj7kZyRihgvsTM+JwTlD72PM7Iu3E6kYS+I0V3V8nH6/w0/4hkPP
NFKIOgByRW8TLhHIt4mdQJNcVse2DqhZQEEzN3mVeRYYWxHMZ/n2VgTiU9UpROj5MLhGhyY0wV8y
KODD7DToXf7JziLbQlBcHqPZ2agXUJ9Z46gfUyTV7n01NOKehdvcJEzj7EhoEWTVZ00qdpntClix
Yx4X1l0fJ9kNrSmpKFI1z8cMxAT37AmlQf4NIfmiAKF7r4iCpgTKCvU4Ygcp0NMvm7n3e56mp8oi
1mkqmyj+JVs0Rc9A3QMiBKjEoasNzpNC9KcCktmWuWYp0fvXz9gKfafdIaZrzUcnC2VUkkMZqxMe
V89ctzaiAKXVPWEMYle72oNCxnFk+hW94qlpdzyrhsPi4VznkW016/Qw2hk/ULR6x3eyTRzu8i0K
gNs371K6a05clEQq8QnsvKqB59SscsBhbvUO+0/foTYpVEsxr7sofYCR5NIAIgViWWZb64LyQcE0
TfHJIOWg/FaIn/I+XG6C/bdqvGfnwEUy6+cAmURU9vlI2aoqlvhuw97rlrejSrOzGH6iOrGGD0C8
b14T37UpQOWfVRf40WPPzvoXUlzPbPERQU9ddqnwLgI/IxhqeEKUUMeJjqRg0wsbHYMal3Mc1UqQ
bahnheJRa6TDk1UcdSukFwKrV119Ovc8WPE6qUcWubkv+jjQPVgflne23UhlaYEiEG16bL0K5vHK
WvEwSuEFCStaI5vm3LqR9bfWIT7W1aT6/R9KutYfWsTWl/tqt5p4Gj6QNCpXthJbw3Iq2nAPJB9N
eb4GeW7bxwBht0jvWmXdSH01HP9SHQEMWqFcsT/nHw57TYKvHFLT01R5Yoh458987I71ujKgKb/q
n/lmlYAAIqQA/x2fNE+paKyyLGKX/B4NFBIrrgfduWdnXIgdL8HIFIivDCKoNPT8mtBkcrU+HaeO
jvztRz60D49mYWwmSVfNdz8dNLGef4xbNsP7OJcJCQm3gxlN3lA8xOw1hvqIENvLNcS32w/frYgN
0OTb411U/zGmVe1XhoKerrRLPNNl0u7aO/VeQWOcO7vvNcDjvPmxiiOMpgBzuOHvp54oBjjIkDP0
x5Jq6QNeE53kRoeOT5Z0jXy+hQlF+Fa9eHT1eGG0yEnghV+w2FkDFpEQE7W4jV2ya7vtyTFLtxz7
YwzJbuczW14x4LyFNYFsqlmcTj5mqIICHupSdXDh30+1r9kdbqh7jKVy4T1xwSN0tYZmFg6VgrOK
rue1Q1oprv3BvW3kX3OkRXW3uMzH+VMfsB8lwmJCvXdkigFljj3qeij/v+pH2dlSWbA5f48L8GuQ
uqPuxKjzDPY8TEVsRn/RnyCZz/tOt4Eb15OqYb/GIv7tkpJ/ROVa1d5Mk609GFn85CE1qtcsY0gd
2lOkpIDmZmbzclnoY9v+1XomUOVjx3IcfVjM8yVpSZCAWWOBAKvaCOHJLKKa1WUrdgcSWHO4LYh5
0pC7QvpBsQ6ZX2fa3G15FkNTZ/aAYNqfqW6myPEmja1aci6U0Bxu6Rx9+2e9I/xJI7QQqJyQKiZi
LffGm5tZyCYWQKqwfdIDC/twZ25Ph2Qav8JTsBkvyLdSPt8MpckPDanx+YXwHbezzXPBNDlAlAq6
FE3GGXAD8frtCgEgS6hDuV+BxcBnifWy9bwZTaZ2/mjmutT3BKjPyAaS4G4D65xV/27fV/flCQRA
gfqS1rCLM2oEqHwyYDvQg6HaBuPn0AsdbPoYRK+o9Hs7pJbs1gy3QCvtOKqt+qTunPQR2bzOb2aI
i0HW03W7EimOKOkKFq6d16VXRGaZKf7oixlbCoYXSsBRn8+PULAevlvXKfzzJfD0gMRossEhiqgc
4SI9lYgwBL+mfH5wZMHzZnzz7zNsTOtFt6p2fHBCxc2dQJfDKcUHQPJ6C7u7xgCNTV786Bs7Yb4O
8s+MPhc7nKAZfMWS9dL7klgullk7kKmhIGD52xGEJPQdOL9CBJEYb6ClXO33cQP+d/CF6EN9yMTF
b/JXNfj8fdtMbKCc+S+y1uON/ekGcqdDAsfAa+E04aMRAKWyHbLWuSZeCEuSvro7wbEw1Z+Iyeh6
5y/GTipmQgdQUNzr4MvJx/wDLOXGFGINr8Y8sQU76xR3wnHnbQLCutSGdw7gZUNNpoKVaty5lou9
K6NqPCSZlHUW5FW5E3AqPf01XbuHI74jsWUpVPVH8ZQ+JWEs1uEIRvqBeD8U9RVYceNYy66CAM03
WxHh3vWD4QX7WpVwpL0E/PemdHK/arz2btCl6I0np1769tyaLNjVykPf8e62/J6/gdPH64S6rbKh
mPo/TvqYle/O6eV5nhZwqWVuRARBf3TjR4rAsKXzP787andw1jIkwVVl+UVaOoqY0c/2Vp9+PMWy
REikUw1yNDgSfO5RM6U/YE/gD3yJfC6+2o66FWzjtzIDkBEfHlgoyPMzI51uaORTEBajc3NhChQ0
qMC6sk8H9Nha42vu1epoh8JqCMi0jPA7gjeoCH8NQUTSq0EXj4iM1hVBK6NDuIVIpcW+CsASO8DN
XQWWig2u7mNHRTm0jab4SFo1fxfgP2WtG+NE7UwjWENnCwRNpk9Ag8VdnvCaOkLtDkCt3BgYmXQw
xC1c02gWburUqDGy2xmy0po1l05iwpAjiv3B5VhQhUcXFvdFIGdVxBxukcejs7H1apMcM9VPX7yA
2iMZqgSAINe3oTBx73X4mg6wiMb5AvuJahxzLoQ+97SHfpt3fDOcm7/73KSgS0vcrrQyY3XKsndV
+JDvb6ZVi3QOcRpP6Guv5IQ3p+thVeplxkZD1KAy0DAC+2ZJX5xPSyI0/yAU/CCtsNbEypV8muQV
6xmGy/n3G3EGngWtWKfp9jAjSgVerNTTwB/B7JS2AYPoAgUsIoE9/uO1MUMJ5MRk6ZoEdFpdcWB/
MWQ0I3uh0+9lSyTCFt/LoLszylPPfoWepSlmQrkCjIUAvcVVN2ccjkjq0/fZ5vJLEM/yhACi4VjW
QIHLuXNiLOA8walfIkfLV85ejEhm9qMDoQz8sV1edqIm25IAofhekkmvO9OasVP/r0QjreXyKrCl
byvzg+kVzngqbiJcf7GN+F+fp1dAatAA+enP097yzDOWT+IUMS+UEoL20+fFOBl6JPv3ZFT+yu8s
Iwkbv/1i6xoO0mbuZVLifqSrvVuuBnY2HkijIf4/AGnwApqlWlsRrzvfl0HWTy68EMGovf4FKJBK
ms8ibchKWWfzK+SrLm6+m61jofU5/Fi1tfabWOP0ucd0lORb8im+ZT2+kRYDm0B9n7pqQep6+EYC
KJnQ54/jcxwstV96Tm4LPcvD2jSSV2xaM3D5VQu1TLUgi9nishcwjwy2I1nkaxP7Q+0x/5X2PyM8
FAb8yS0mXC2h28YcOuPDd+Li/igsFTo1nx4n927aTL6w6R50JG9TsRQvxFmd8tw5zR5/e9ftWbCV
bqm+kVwrN+Sg1oTu6/I+9Pcz1DRLRpn14UAaHSZG/tIaR86G3Y4pzMrdOcGUAynN8mDNes+6KjcZ
x4sQskWlEJdoSgaFLWuTgMcpVYTcin4enpYRGEEHCJrCQmkcK+AZQH4oMohcW4j+1rQ6K9FbcMqR
ny6vQy7fQ9ivyfLPXotikb/Vo2JRsoNmmRI0eskoJn5x8hpLBQ75vIjPNVBdXSyKEBIoI8+iaAif
W8Nt7hqW1REqTjzGq8AHMTgNV+bIutl2oHrRQoI9VjxQYpBtSByfewcIcrjYqFKmaYXS7WSDOjpO
bvinfjkJM/Dl2sRiSGeZf2A5xpdZbJ3BVbEKvbJN345TYL259mgAga3pecpYMchYzxPkZQ3n5oKk
LDjwLduMapFlGTJAmWPS7EKkN4TviqRfYatALNj9opHkhx6EDtCSs6L0WgC7DWPQHsf1nuWA48hm
eCgDM8e+8T4aIu7NT0bhakv1V/p0pkUSazTsO0qkbZkLXronP7A+Xyq1y0x4fTOJcblY1LK1uKw5
jbV99RoBzK/m3jPPPbfdxJeqN9DOTbKHGeCDOEKBzsyzZPygwXFm14lc+BU5lI4G8SZZsTw9NKVE
rSUba12tK25x8xuZWJbXqDbT1kCbxVvvF2ww178nSjoi8Qxd8Brs68yLQztGCdLIYAUsPGRQC7x2
8koaq3d3nnWD+KMetvgrVjKT/BwtnPutJg0BcVMghe6Oz/EVe0Gpy7X2Ga6T2tdV1WmLprTaMnv8
icKoGMCzkOUZZDxo+5VPdhKAIsiJvvmE/GnBlOVIlWfomizkxpql8J8qLa32Pflx4jWCGP+nG+pR
a5M4cRNf+ha90jEBJjH2ZFjDwTNEfbk5RLdmbZxUYexLYdwCWUu312F0pDa2J52VxlO8aEp4I+dN
FEuxfyxanXMRbMwk4YgeyjHKlBrs/VcK6rObb0eIh3PpA4RKmysqFfqV/wPCSHspA5TMlNYIuDmp
q+q4J6PXYPZBBNxGMNQxthctLzrLk72M2iJZavqPr3LvfI1XOUfZpZuxRRnfFrnPZfDDPAy64NZe
rKevZPc4SbjwEMFq2i8oIpzcBXs6aKnBqELYws0VS5JA5TlBla312/jNlg+vxlfuolq0lQG7FRkX
1VkE7iyAarmKEjZvb1abP+knpWG/exD6taIPrshOB5rHeP/Vc+3WvcBSfx9qAm3fjTNcZIqR9gLZ
xR/Pacs1PuJGFqgfwR0v+1y6HnB3GLRr5y5q2AK4IIC4WZmqUsBK5hId18Vf94HImGofEj/ruiJm
3+1oYjwSzzqPFe86kl03xwhoIk1jtaszuFJCuMnMjJYLZ0QCPnfyh1U4NAw8MsRklloIgKJTZGqf
qr9Ny2+OThJqgY3vqgTs+XehQBKNictaImR3h3ZKS2ihrSGeEUrdwWC3m3yloGsKSzb313sZj2KR
Uq7YgVyoNW2iNOKwWcmun5RtIgfWx0LsCtCljER6Fa+mTl11CsipbyMBQFWnpgc4rPJwTQHP8ohc
qLH+BC7uy4VDQztYwUy+Df27y0wAQwLk87606/t1sa6Uv/DM+LRzSYoy9zhScfUlbIisMXY1cxNo
1iPXCEr+gyFJoBlkJSpdhZcoZC1JLe19x/vBkhts5d+R54S0SFZ4WFgv9WAxtj0eeXsN60G5GI3g
ry00a2Ha/kYc4IPs0vGMPKMnzdbbLeWdCqCwOwfy8DQMIIX9uOC5QhGnRI61kxX1e6AttuMveqYG
1PJjMl+f9pIFTXBFkixCbpufJuLCVgCJ4n+l6TJW0tH7MG725hZqW6T19KcVu04AHAdZHFzr/vgI
DYycSBHJOXHM5lU1l0jaXBYD69qZH5hbjjkzf191N7uifuDzgtfN7aGB4CmmGnz9OPzmtLQBZdEG
4VtubXmNJHKWFJ0hnjVVBnEpUIMVnKeK0jelXLjsfNlQRdVmOh/rmicxaSjCmsONfzdRNZcaeCXl
fmCWMzLdeR84SxSIkqMMDvR4brfWoDB6qucwXksnfHoqpvV7R7aHvax15ascsgLgffzBPN+b14ad
HzG9rm6XSkRFF5d3BmZojCQ1o55BpmrVpbOZ4mG+ZZh4MONGGVrYQ92pHUyStfxQynh+PYD+j3U8
fAs09szoHRT3odU5kQaj1BYFHd8Nc+3tUwsCqsuX+jjHc/04r/Db4ZYkHJNs/wqWWshPzXmAQTKT
cEcK3l9Qh5gOtOz3p3HqOwiCk+/TLMUrJDtP2fE+gWOw7NXNP9W7pRMiGmecBl/i9+eEygfv/dsA
yakUohAxMxLTkykPKuGZTaB9LcvpNAergL4qzqmzX70WXFU6N1ww9tKWa0/YUPZWnw2MnU4qWBPq
OuUNmzsYasjEIymHBxbZoJ/woTo4f/qsslcXDfU+2YJM8l9BdpOQNIrCRtFcj0b4XQOBRhMBpXLJ
jDMoWm1nZLONB0BFl/6QmN34ozZ8boE/KVXoOhjfddH6yn1XMlNl78VDlAaV7ag8HNeWn+bdKtPq
lv1wtnHiAg0BY+/LT2cfoHlTCGiXtLVfYQ63prWOXR2ZC3iRRqDtJqPg8Ee8bS5gpdOY0NcEDY9b
Zz2NpEuS5G2gl4eB5WJV57rB+FqV2xxEe8gAnxcRfOSwFPk1wLs6sGUU62vlG4e/yTYxFFY7TwTj
8yOTNW87/wEhaaFfA8JQ1LerzfhHHL0tZOf/wKVGqwIeK03GGtwqP7oRBsgJoNM+zLYbggLtlsA2
nfH23JuXc6Ii3XAkJfsf+GNLaklzPgmIvYg1dUJ1RFgXVtKXg5k7E3B18Di5xqQtw9M8UESHEfun
IH0gENG3phNCxqhPJg/gEGBSbVmDcqgqM0hb4fHbQbe+kNIh1j486Md5Hu7Ptj7y4RydnIhfo5Vh
tFak8b94erCD4V7L/w/Yju9sfm16222qD7TFFf8pvgdWT9hr/g23D0hwXSRc7i2sBWmez3eKUk9H
R2ysUNfT45ofR6Y8XRKTGRu86Gs6lL59VRxxuyezPraM9IxT6ySAzkzxL0+HuOzHve9jcHFhy4aZ
1XkSr+9az+QRRA8U9Aq7VqXkKzMJDpLDdeRSvS2mGinz9C617NTBivG29oMYbM5uapno1FbpJs99
PtF+gPYIPJ4UKrwuf9fiRz4bnUlVAl+D4hMDkU5DaCek+wRE2Ox4O+0C4R9eTxW8mxfKiglCs9/f
JEktqt0gu9FWvcPKITB8Q5G1BAASyv+kQ9L1FKpEtpv1G0/xdPafG+dgrufzrBEEAOptSfFfjx2Y
dKOehlHji+PHvOOHLhqHiip7vcS/yqrap6Tl08XYi6zBXY889J9QTmeg93hldFonv42chzs1okkb
GZyDj3W+eWTiqE0KmPDa4HpAtI2/2BXEOSXEyV2ScRqrZp7S9ZRDGhpl7wiBfcJsEX35p35PdA+r
Fai4TH+qegMcixRKeMPOHSmHLFIHhHLraFN4uvbVvpxS/7L6FbHrC3xTcO7tM0jRzsHCzsNTjEUA
ukvJwC0AJ33hA2acW5cIPU2pxQSVjEP2kmVUUbB7TD1P0EtMPvbqHhJ32jxViwhV75Mxlpi2y3X+
hfHLdgAp2ZH7UhrNjZUA/O2ZTaPCrBhzo/N9ueI5Glwo3ieEQPul2r2lkB8MVasNozLAEYGjnc89
tKsfL5itzZux8XZozRMnBso5V0N2RT8mL1NhyNILGohNZkkYEJ5DMCA3JE2gQDy7QnhS03HmPrrh
tBC7qmQgnIrIIisrb9xGqmyecj7CECuCJrXJjblV5jZoKb9U5oRWjNV7HrrYSxHJpxpcGaW3hx1X
52Ce1//L2vapAUbeViYN8fZib+fbIgOzHcuD6PrKzU3JE4ZtwMAKPtRbEPthNEiT9jXLtjNotg48
0i/oRLV+1GBGb+uwMnUQ3Sxpn2KhddajtxZPGDxHJu4LcyUo3bgWGLVuuIiEqKx+ZjHwL+FhyRV7
z6Ioxef6UpVurqeb0/Arq8+iI10WJic1b1p/LEbkuC+ZJe0EjtsoWufLWo0fn5B+YEv9mD6IlqYE
y0D6MbWJirBorlSQFlw22YCKysSy5aUmXMaxqb21ELHCMk9nalXxFTiB03sCrMwUIe4BEVpB34sX
yC8bpz9Y0aTT6KOvIpsQPCW2buZ1k/IYpEL6fLuCEQwXFBqYKos4Lly9w0y+e88EIE3DYyya35Si
aOH76M6E+o67pAMVGJso8oziIc4yvsQOqVvbyoOpM7CYzDTQpf5Cr/eYsUXlWTLJNyK71SOba79F
GohWhDxa3GFNiGZwSxpWOuwd5pztSeKHb241VgYYpjci7rSG0Pif/PuNs+Nkxtb4SlGy8TWw1tAa
Q6L032B4h5nBCVUW3Icy+VpJUifmuiQoGppH1IpIl5/44G7msUMQ9dduE3scPwYINXsLz/OY1ABk
0amd+p1aVoYaLAAQ67HemnyIhlxWYdeEbpqKU2NX2JYevoiFrCH5rSQC/Vu//k68w9mE5IKBmDdV
Zo2WyMFH5lkowYX2KgtAn165RFcNolAnxsp0zi0TmMvcFo722/xCffhDX1MwevLV1YUJQaBnIY85
C4j+soTBB317J06cIoWgfz50MoYtWwKeLZXcVmXnMqKd1KqMIXer++zUcydDhB6NQjeXdXWL7tRQ
0Wqr4yhFGgZ+jxF3crP70aIm0JWGGkvO6ONwdUAh21C97b3FWO6sQXgDu+cYH8BkV+jPbwk2W1Jp
u7mr3PzXUofKX6zhviAf81QIxrPnm3mbVuIHJNt5bsA/2VZ1g0ElUAXDT096dngXgr36Ze8PR3VO
s4fhBj6Z6STmr+fNwZ6ql9RnF1q47GJjOyibUMqaCemjDrkLHGVzsrFjJooE5mwcIq1dOuicNMeb
CxtMNDW8WlmuRuBbjHYzCDj0+mjhp0Ap3LDPRL1qNHtUPTwwYzjkCSd3hqaCmjSFlWvx3MSCD7jn
Bza5HEC6UI6E7TCP5drtj8uxU5LQh1DP6i42OMA12LmhReEK/K8LFM1nX9MFVIu758GwgdVPVLEC
YlBC+TDfPPtReb2hYBGMQBcNPGRQUupgaM3GPugjKPoEgzyZbB0uNY/OcrXe6NiNXY9YGnUYu2lW
djj5wl+Nd6fggbkk76Pb3AszbuwKEtWh3dhAvLhm16GGsIkWvwsFBxljIxkDx/KMkq+IXTLlPdzU
ahs4C9tNs6/B5LTrf5acRhXXb6dtTxVRVSUDzaUbbl9c6sUUSgTOsPz+3u37MkdcybnOZvNtfp4S
f1wxPh9ki3UCoCkthEHsU5lGkNK/htZlRwphO4HKqFTNhrvaHIIgJ/oVdYOAWY1JLcIoWWn54DKJ
AIBd4u79lNqabOnkqU0A2BzEFgPbAzX7N7qR8kmPudokkQOS/PkFvdg/zMA7dqfROq2PSJ3/4fnG
9TceyyawbWspQvpcsQEXdFhSSO6ZaKeu1QWKaaxEjcQvPhAZxNLE7Wu2opyNDap6fR8lnOEEKVg+
Om4Q8lazc/Tz3i6tfnf/AHszXl+KV2/lQs9fLdD7T/cI9AhkOyEMhF75AX9ok95YjhAXifNdGbyE
wwLJnuia/N7JwaNynDu7lxriLN9hi/I1uLeKef1ezHJuL5i1rjW2m3+YzrO6i3gR0let1IJ9m9FD
mf+HukDMC6OK+utbhHezYW2nOXC3fqtUUUzsqkUg9cfv3W6ZgptWvIue9/P1jQ5VYmPmLHki76qM
rBBzDQnX3sIHYdsQKkXmJMh/YZzco2dFGbB2ia9ZAwEiW40m+znevHnetVs9gLFk5Xo7YZdrI9th
fDJCi+nwsgUy7ELQG63kiE0D7D1ecCBuJPWtA8G/EbY2Cpj9GiqEx5UNxvQN25HtlAH2y7iz4yNl
jtlFfFYwqxnXq9p+1J9JZ7xB/unXsVTBKWks7H+N6ECjnx61Qz9plyChr+QrV4fYli2fOMQTkWEj
Ulr3+hD/4DiPzTjWgY76vyYUf8fGB+7znLLnDKcx+00mIMKEH+3M5UTGSsRfyQBlBEpsqX7xvxmS
aZ20v/3O17DdKbBLlkiSbOsT1hAvKaSD+NlKgjGE/bX2Q+4g6sRJa+pG9y1rjgNBqU/g3eZbusXk
MrKqT1hJGnRGlSPBvAxxI5H854kAq6ybpV05QuHUeK2kMCztDjXOd8CEa22puzMJWlTlbcIJW9Tr
LLXOe8nLJHOX6y+m3vh3X1QwgPTlTk8rZIuCEpvfd37RDjKhufSzZ3V9qKug6E8L9LDRLX3qNI34
yv3kNZZqVuK1cY9d3bPXdI8y/mlgTuVjA1y+fC72BJKn14Z0NOk9qWOZmpxKQX0QJSgg4/NcbsIJ
gRqdhkOCszju5rNsUTjOLZ0eWNW1Metjwf4HvS2AWqkfixH+n/q7ajMsdAuxfCqrxqQ8yRroY0u5
OzaybMiECu6Vjm2C/dmUAbL4BLyJUjA9kwRLLVMpQQGLk4Eu1C8U4SDOw+UEhZcb8lv/+/XesFDB
bNmsSLvUDQFkoSVu16W+ZAtL49ehjhALDA3Wbl0FhORdqXUzFD1novqE0EW9QgNt7+Kb5AM1tnKn
NspqVymI9Cq9zc1jjqZn20Lxnx0zEKWA2rcYBAvmSHFFz4J89x5Uph8bSHu2YKMyzoKfSY8nEJ5J
Eo+Nepipay2A6FQ1qDWZGjyBSZZV4yFncR4JKf+5IbmXJZvYmBRg0yrbSy821kOc3BQ62ILMhEyr
B5FrPuL6ZUNM7b1YfVookJFRmL/c59Pu6N1r1BsnjPG5HARdEHkfInXwvGSNsFQmc1PgLCSLaEOJ
aGrOoJgpqVIkdsp+Q3YUATPvA3cs88TcpwUUcXdFX/HEzzKevekyTfFtRBleAVhuL8D7X+341SFT
WkhZKhLJHIShKYUA3tbhYPOxNn2KhYQEnOF3g0hyO71oROOHDvlcnV7Kx6ziVI3lMLa+gt7TxKjC
csXiqXffL/7UCkrRr8GIc3FclneWH6mnObFCke03mmS5W2fVG5y8OqUmDjrNyjraGYIZi+wqyDQP
kg7XoMZZBw6WmCm1w2Ry+eUURKx3WOk3A5OM3IozXGFvx8PWiU7y8gTzYHY9xDL3uSennfcJT6P6
CpFg402MkwEOLspoJcKdZiTbF9hPetLuJWnd/KnPBtQD5uGlXrC+CS+aNbT3Z/hnbVDEWAA23TNL
65Zzyaqvril5IBBghmA8eF16wGiyTubqEU6o9FIwHhW18ECXmXNlHXaqji9Xnpeq4+kR6zFlee6h
1xYQLzFmeRkla3LSQoGSXmnyOCxaEd5+53yVcD/JqJn3LZm0k+E32jDfqrvidxqjro79mhydgfqX
y/eWdAIJe4k0vE+X5fjjmmVSjJkNwwvx13MzF6+5a8fO1CFkDmWliikDwyKgnDhd0UuGWPTWPEyC
/khozKx+A30yqvN4iZ29juOW0y6qylxNewt5qIBqLfhbIzWG4EW2SoucY1ZL1jBPro26d9gK4Ezn
azGdady9zv4UIWZiTZYXA5KvQ3nJav+tEH2P2t/e3BxPQgMqVCjg4YVy83Y9hKr7gYeYYQIj1dT+
hiwrJgPTTEtjsEPE/oNfSktpehdpZwUECPF2EGjqshYiUE0tbxTvUXoCPD7lQJSrIHJDPZNR+2eg
luAfqcZztGu9Y00jMDq2IECG6Rk8o/VgWK3Bxt3Mcl/P5Bym1WMcvTZA35ks79VDXrLF7V0WAndD
iJwXkTn80Hx5dTT2+2TQ6svlnO/Wd3RKFCTb26KlrNxNiMYGyJ7B6BGw9mVcxcVcNhhvdULW8Zp1
tLgbC4rFCXx1JUFHjU3hKicV4nzVZCmDl9q8LiwpaEarRwRbioAhzJa5AZkSdEcBJqKS8xypX/py
E3p+vFsmoAB9fGL3XAVl5PdDjcV8Xrl7YBTeOq8AxwKjB086lZcXO4vfx4SMohM4c9PkCWFHgiAu
QbtIw8oBB/hrOMigivACDut0IKgk1e3o35llZ+Z1PSiq5fu1dqbvoGfwk76B0Kc661zfL2t0+ix0
ovjC5c8CwuUrs2ojSpVB/4+6xSGNbyISrkYLyU+85qHChyHd6uIOXGawymDiLSG5pQfZ+dXMcpER
5Rs6v2Amv+idQm+B0UQwKwxnQV+0Dogq81i7npghpY7z+l4I9Hgjan/ykV4sIPmPl+48kJ2ZTdOX
4WrKyZzQ9wm/L8qjkxY9mGHuXRbbVdgGLkPSWFGMApFgA9kmaop8yeugHqzN0we6u/JYdUuoGXvu
3bLQ11WuZEubdelJBEP/fo7Y2PHEqCFQTx2VI2fosdJWEs5S/VjYGobDS73bdkQZb/metfNthPWV
eI53/7IYvue87gU0pWzU2HmGlVcIZ28lQVMFB50QV4xZkLaFiy9IPzs5k9E44HaB4w07Wa4qcNkn
TC96Jtkoz70bMR3CGTGtS67aPLgud/E/vRW/Ttq7DO+ObeXROCOok8DP8rFgBftykPAULy/W0XHh
XIGvh4iajMthJXm8ZFdr1Ramo3mqH6gEvBLIDqfmnhKxT6ZWlGhM5IJR6qyrsE06FZ8++Gh6fnl4
bMM+aPr3B3/8+0vWLmc7Gf3kfKQqLsNLZSWY67t4OoeOHiXmhuhuNwngqcI4r3fpeZbfRl4JoD8j
8CPJOj1REfYZL/diSxGJQ81UxNedYjZSR7B6Vx8YtdNkU2Vq5v4YWDGO37w9IBhkMKZ59vMlZ17+
4HCSR71CpKXCp4YcwAy/v5JoaxikfkM+9I5b8Tp2RoB9wWbQ9V+7SSNtzB1Yuss8C93oXNLoudIs
nWxme39t6yMN1X6JrQ1Vhqa9ALxXZvKhIeHfhnS1xlCKKRHXB2p8csfe88Zz23peK7nuIgH18cJ7
BoCm5KUBspjLb09sI9HbiDE5UlSD9ewROIn5aCeOQJSTyY9AaSan6CXyI/zkRVVBuZb6lIwiiTDq
gwP/lxJA6eFmHGleZr+57dkNO7AFHpF5gqFS3JI5qMc5czOfV2lQy+T0V/VGUPxWinlL47YLhk4Z
fMSEffmHHTneAMcyjXIVSr3moac+rGZAxD12dAJH6Itei+MXzChjVDgN42LCyNjBcucgeNGhA67c
Xstg0lNCfpjbYnNRAEN+rZp2rDDr9v0KH8G3PLQpwbnt3yfVMK+uPP2+f3uL6VsIM/z8Nl0kaOhe
tyPMtGQIDy+kvrPfkIDnWAhS2uVKjWHzIZdv0baCjMpzhvTeZn543rJDm1A/wAP5gld+z851yjZf
S56eexUXG95VFomhi3Hr3xL6angje4kMCntmU7+gqr1A7cs8G3rnKZHJOIS/LD/bR5uS85rffJw0
CCmZmEPjwF1IbgkVOOJPCOAsTKsIWSPB1xlkTqTVNxBj6PLhIt89/eEfcjZcjsalm3sFnjUmT/em
VoYvmKZWgh5dpXrMuBif5PimdB7xjZrca3l9BkUGVErEpQCBO52pV2QOkvGIIifu3AMg1IDURfHX
+okA93yPPMHYcoJ0/ZjpdhjzFALTpoL8IEmI2QykVjl7CMdZFtAZ54QZHAz4DUXRfEzqiZZhPcjX
2XvYOY9SQ1/Qwl+7JbEdb7KL+JKF4ClCELEhzPJIhWpUA+k0hMejQqdRxqqrZkyc9QLQPZVKaVC3
iSGlYgdcNb8sXKFvLnqZLRTrMAUHa5eaoDb25NLLEfXq5kOMAnAOfWSdqO7lvdql0QNiIl8WVyUw
fRxfbhxuYveQc4C644J1ECIR/VW4juTlB61JfS/VaVVfFiARfS37dVJB6Lem7Iis0fS5YqlwJlHW
+uZZwqgX423d663cDFnS7ptg7yqLfivT3CQeBM3bBjxWtsOUA0NuZEmlJ8CTghkZCucFF2oCFXt1
OV5thRDpMmDqdU/pCsApdZ361lswRLdHx/PbMmzxtCd3gjZzZ5JwydurxrILnciFYWlMWUWDryJ/
5BHSl3XcQKksyr0dDQeCi+aICTA0Ee7d9LRyZuy57AYRbMF2oFOQNskvaSm/hdvifIN0jRt0bmpQ
gWOuv7s2C94aZDRtIWv6M2QsGFLDVUl6yH9/DDIBLZf4Gtf2BfItAPrUwb0lWxHc5VpdMuhtuuqj
QskQsADo42ESftiFca54dqJnte9LfS0y9CzethfDO46ztig6prEbyylfuELvA7uM5g9DyODyGGMj
IzCmrrICYrNxXwHzmu/8huFZq3La3ELL3AB9Pil6zrSuCOrn7GAqpmgonDs7NVQczbqxyX1dwzOo
liQMjQPdmk8+tqzJsiRaUtFwbHjSZhmf2ahx+8eSEhJdVMY0EmMmU9OBKLeOhLobmH3F6ThrCTEI
gvH15CAr0NQgLMobWJfpJ2Ynw3Cg/5mDqcXd+zhRsEUlmtJr2KXkxlce8oXocZhgdt4MPiJr5py0
7hez1uuefElki4A4zZ084JQXJbilUV2zmWDd0/RuzLhw7zZHO1llKQFj+om7sCg78zut5dsinUt3
YobnhQpRr93o8kcBHSxuq6GDO6VJQRS34sdvAXtTI1YUc9BEBO5VtpYG0QhXvxQ1Mue9RYGLj2nb
LojdfTBAO7kuc7FuRxuOICfhZyWDjMVL4NrTSPERwMZADcJWXqGkmpOfth5bewYWQ8vOa6FktvUL
uyKojxvkLjoWpZ9FliSuP5ujqUjQHDfZK1ZwsqMyJLn91WqAWI6kf8bM6YA3L38OoaLpA0zJ+XOX
RVL3+H87ocQJSrQpvs9coJ5p8i3bqQNjWeLjcOUEX7zXujmjwrOD0G7YW0G8kazVJK73LvrNXwhI
T9JQKJVq4n/9RTX48HXQYTIkVXsjB3k7V/xl4MCp/VhmRHNGguTpP+q3B58/iLlr29wa2MnoAxIq
DxW9lDnr459hb455vuOI5i31g89Bm3BtYQFvmBqL+NimcT+Jlb4EqdAKl5ir3+ZOJHk9s6R82O+M
6FrufMDwUIP2xzUGWu0el7US/4qb0RmK8pSyVARPrjasvtwFwcgUg9cLVOsz6v1+RGX9/tqNCYyj
cJjkyaG+INmF/MvkfnfMTzqXYTsvC6tiHLxR6aCaN08i4Z6rd51Z9Vs/BtscSlYg0hB1j2MV2MVZ
vQoDjsBtY0ZWv17ywAZokL6DRmcMl78DFWIUlHYTs8No6URwm8t1nVbRzHLiuAVU4/QdSU8iJ4kY
Br7sMZ+iZXweNNQ15RHG2/NmLDqYKnFZT0e03y4Y2/WvIi2ZcCQ2hCmH3LRUkpEh5hC75Pm0Hnfz
fXt6490nNIXic3LK/w7KMreKT5eXa+m73xUIo+Tpsxpklhq0zqzAbS3ynvhoQdpw4QY7s28Q9Imf
2jsDsYQu07ggJ6pE7naOSGqDVxYu4sey63NuYSp1AXSAejmU4vYeaD2wjQtRmz/3CW9UG867vAa0
1oxZ19Qsj8xTLUVVACbtHGJRnQg0em7nds5FWZ9pcoo1w8F7Emselqmc7E8k1gZ4iPGNlD+KadBv
SAPhdeoVmYoemzKKYIn9MGh78YhbHQCOogvvIBHphCkvL8QKu7dGttX2s/VM64i+lvFUnOvDNIdU
t0yKcn9FfIPUjdCn/Iq5/kFHHY5VFjUgwL6Ei4NV1oF4AnH9ViaxL6uAmC9qEsELql8vjk4njOco
Ci6uGglgxfQCs/i8QCFOY3bUGo9/SaDqrekZE7GIEIfjuAGqbERbq/m3VLykmux4gQp8y1gfOCLK
rTKHN24jfB3w3eDpcXp37FVfwGAODghaLOzBrtMnmAVLluFt8EYW6HGwXbFU2AF2dRfoJqCeIOrU
7W73YdkOh8y5B4OQ/vxja7MrfWe6Hl2LEW/ox0Pl/FNMeH5eUARE3X2y7HIcBtTJjoBCtqORnpVM
vxYWjvJm247sDpVoJjIT3s4ylAno3sBPUSxPoLPzilhGu9hOPVXByJtDRAlyfntiXxX/7lUjHTyL
p5udObI4tiJ5xQCNH7LFzNPc/OqtmadASRINNx5eHtOFWmx7/kj55pOO4XUUjr1fUgAziuwua0pY
GmvGyI+SZvGj07Q+3VWDtv+T/CHnJar2eqNfrGFjPJLRrHiTyjz78xNzP5sJuKX2ZWdgUGq5h4Tz
h9YswUhS8I2RL11glZsFStDGb6xC6G1macU/HFw/jO40LVP1UhxVAi0FdlAplw0sVG1V3GKsUI2H
sgOIfVG30asyGtW3iR07RV2PuxDjXo2K6M06D6SNG1iUKe6x6Cgv0nE6lXIZJfSY9eqY0J8LCtlw
RbOfJJuICkseLc+l64wx9IXWxsUSK34CCk7+q1CkqHytmfhzqvl0kTek/ZPFwnkPa1HGr3HS2Vsd
fLR1PcfmLxZojd5E8W91SJ88/XGmufhhZOaKAXT6f4PzY7uruyJ8BOMb7VlPEiwj9+3vCbKZ2tPq
tRSBYSdYihVWhfWc2wouk3YHfOX058Ifl+OnWKAo3IEiT/8hAvCHcgDR/elNo0GyRCap+ZwsP8/6
Kh/kP2XhtUpefTLHZYZtwCZTtJO9JdsZEd+z5d0N4CIT1pVD1VeHxQrrFexg/YpG5eEYFlPJkFQ6
8/dOyQtqD3AzLAcL0TRJWdoRvpjjVdAHYCp930L7TouVOoP3D1sHYdOpTAUbDeqDJZjL+znPMmR8
cktApfaAXOhsjo0LVXZuDIyZEXITBVynnybXmGZBo2mQA2N/3MrFj7J5s0LiR96JM6GX1YqI5oQg
W8eOTGq7oZ28e4tIZ/e3ehLAQbOJX/UdPwjpdZAH+v3uQudL5TaJm8UPXAEPcVoEgHwpPmROj18h
O1PXgA713ijg8Vgsx9SEqf5q1wLjxEYx+8HozIDAWouGF4OegAGess0fUUB4P5+7WMgUy8esoKQb
ev0rHLdJMX3+wihzoJpfVaOZ7VU8F6to+YFhI/HGwbsaKTs7oQiZvWtdomqaoJixbjdiwRO964rD
jEs9b/Lq7/7hpcudfjC5T5d7ZDB7Akc4NLR9VRlTntFFnRJa7+xlf3rwZ261mRPeAZx+Yzku4FK6
D/j2hgbeuXiY45cRkiYzi4bjHTlrlameM2q1OWiEGGs/rsmHGfxzfybnymrLwpbPKg5yz79o8kp8
t+MCW6u50CUUmIE/J0OkUS/8Z05Z1wTnRoQGX8t/oz80nEecDllX0oj6T5t8KvQNG45RMdgLR+Ed
IQnfObTJ3pkgdeLeDDjSWpZyLhlIB/cQVySg+pM7FG1GVEtvuagST9ANPrs4U/mhUQ+/PmMSRYY4
dA8A/SqIEtB484HCXWtbBB3ofJgG6KY6HXIOs716yawycKg1Qgb3QifWBETonuQnAnRLQ9HQK9/J
lDTXtuw9GBqHSn/Q0IGZilCPidPPrsqXr3vFU37cdtB7mDKYXFhZUoI2nLGh4b1KKx+moLRpWewq
EGfXO0J9WOrZtaRUXYrS3pruhwjxWgki6VFbYiBZBfyxM7oTiywPhR6FwAcySSuVG/1u4bE1FpAb
vA+XYYx7vQiM/ecD4NIreXUtKYn+QHpTD9Irns4RxYBEdAML0NYQB/2wGxai6eXCamRlfeZVnW8/
1iOG4ZlzcI/nXVGNfcBJTYJkNf1JG3S9izzZ390fvKy9oQuxaV+9LQ6M+FyOevyVtE1muGypnRev
39JZLi+fbUT1MH9eEfWESmfF7ZSpWGiRJiNtG6sZrFraDG3MrAbBG0+wXDhrCyvykBvzDSQv3Ib9
IPHB3Hoa0D/eTQOo2U8Po+Ff6Sb6Zgkpt+bAw08XQXhmDOKyTYQ3KHtKRPdNcI8Strke05FY18Q6
UDVp/Z0KpVlei8GiZlYtKVrZ4wpnIGDZNPbxm84W+trDhS87U50kgo+yHkUMzx3WzSpgyTs0mh8Z
bypu36fh9slVTv9ePQ3CnkGeDPFSJZr7Q8Ky+zYebWikpst0OhB9AKOOt+6nRuBdmCPtu3YYz7TY
9SDFuIFpYXn6BDVruWqKCGj7oHWuPOcVjsURacUAJZ03iT9eKrQSoMw3WM83pdbloGQJeglQ/HCg
ZDa0GTM5Bv4ScaiMjq5/3hTWWYMbYYz9Wu9FMvy1wmpje/zpZDBso91owJ0bZ8NJ7cXq0AxLmfUE
0zGYRJ4UP747ohs/rnTq9oS+1ZKH7JILxaE8fM6YJmoF6ZgMEkwJgaPRovc5yOzDTKJimkOCHb2J
O7BzJfDzvG/uwEbpqtHqu6NN0McL13hx8qLTmNqobrDgQDFK61CgN11aRACL+1mxwa7IKJ8U1vma
TN23ZKotbgt4F2ics4V4vdjTMEGDiBFrnZw8DEph4dsddwfzyTQbllDikunfAYtA3mzoBui7K3m7
k9u2tWUD0XA3UQA4oHtIuRRbUFF2dJgfSVS2+RieooczanHAvna2fTnlaxyh5TD1nnzrmo8hXhOx
/5hhz2RT6CO5rEJkK2T6yf9Mk0bupVEVZyXCVCE0M503jgcAmjtJY7YwQyCjW/sCuRRWXoD/9y8c
7CYF2JI/nN6KN7K+xuL85L6No+O/Ex7M88jqORoCa/SdvZydIZPhkW+IwiRZwExRw7/SKbUMPXQc
F1QRsigyiv29NcuOhnqa2mdH01q7spdvVd9LNtnMUeRxHhD9zFYFNRW6LJQ14JZOM8FaW+rS+1zA
EqU7ZqUsHtdrJwMS92IJLOayV0/7dqkA/HMdYEGHeLjYZtZV79EJVdzmc+jWQXCSPLiY6MNTFie8
4WKGXmQtK43nDIi78QiLyVMblXR3bILsTUSq5Eae/zXVeVaNG76K/HPvoUEe5tFP9E0mUL2UE5Mq
+K8oF3sbVlPEP2rC8TOJdStfyfLR+QkoC3VeAB+hxkKIyCKhxXLiFKf07sVJMav7kpoC9x7DpXyV
yBFaORcqh4Ep74RP0ZSNtKRpmhBHx2K3T2T4V3gFMvrHzPnbAEoIJh0SK3vV5G7xyt8fG8/iKmPK
PJnNCaIJleMf+t2kr0EV8KtvflNwS532OB9eHTfOoqCohoeMlKRm8WpZ65D+1VpMCgYxlogNLzCr
QoEalH2Fv5TOiZk3c9b01z5n0CQROsAo4+OfKRB1uPf8htCVAr/vmpVdkvoQENT2Xx4AGqnwXxHd
txHBJAvdxto+fUb13rZgH15xzLP0VvWGO9S0Gs7p7Qmog9ePetA/XdJ/vgczEITWHOGeSKL7OenU
J+lFQzMYxveLNdfqcIiS6GAN7JgThQZterXnznAs0S/i4PbVUfMUZqYJSv0NhDCGp4AjjXCwzXm0
Cg17HJLZamebh2zMMX0yPzI30FkonBLfGikFN5rskY4SQsd31t0vnglJwjoUFJMYHRsTPHziiyza
hZKzhhakL7yav3o7V26j3bzyWNNaAINI83CjKxZvkFawNiJ63ynD8i4B2GzJTeAtmiFmP5M+ry7o
6EzggUsNNQTuRO364R5lWbUR058/aV+cVDLAXKNXsvBj71nbgDI/Taij/Kx9SQtGmq2OMfvNmbtr
kbUu8pvSxxt+EhdxnbAQFzB+KOitn5a2iFbQVmS1gl8PMEPyOnj4lkidswGujpW6DPnuoYhc1WWe
opIFNClGOehwKlgqQSHSuP/11ImGAjsikqu1q3wgRmlQPjTiIEPbUoR2/OeRRzDwkiod8vahKleB
3E1YuXvU2RGW5ZVXyRvMAQdCY2DWf32N9yZWrhmArnWs/fftj1IKsfF1fBqDdmkhU9sNjfHuNhYB
uqty3IVUARymqjqe5fWH9j+upHP8DLLr71gkh65P4g/ZDSJ8rWkeClDV1/HqEo20CwO2U18iOACd
5f1uv3/RBy6CocRGH2c93xxfDVT7VK/67QKaujE1BDvsLswuTnxjK24P9pWpcUChjgGjah5ZfHqz
mJY3ZER/hcgGCijiL+tw9jdRm6VwT+VXw1g19RBDl6VUEsSaW5TeMeiQjcKYm3ze4ZEJBWr2upz1
e6u8Vxj/h1WS7yT4Xz3i7UtpCL0wcK6rFBFNtCxfX0MLVH0BGd9zs1teypW0gBPkVF6HBkcF9p5L
o6LXNic0dgzalS2lGS4FeoTn10E3Qxd4eKUXLTiD9mGkc0y0QGCnfbjy4o8AY5BtG7I1tfh2H9Pq
ZV9J6GwC1fZP44OH5ATi/HM8WweHTvFZGYkEm38xlW7+d1A4tTDeBnHtsDN29lH/qViywDnAxogk
wOpKWdwBN12m6i++Ub1Cz0I+amKmjjQ5ZSp0/8z5hMKEJ8r5R5ABYGRqtLyVgJT6he3jO8mBgwYv
M/91GJt7h2Yv97nlOxu7XqhFpLuLP3ZFEi9GwXfa6wdUrFo9JPG4tev3kX21n/LFQOVefngvYVkM
2i4pi10nPoR2kIOVMVuz1QdgBmxNlMYtti3rxHmFBpIEY3ChnGg9HUKuHj/f/YvIYph/OwjISEyt
rzY6P/iKiXcIkylN10dDEX6/u0VYzHu9p40EPbK6+C1Pbo5ZTv5Vp/tbDrMedY9kiuxOafJzaDR2
3qVXTsGuyO8OuOTut2JhVK/evZApZ5/GHwyV2GaBzgvdxIXkDtk9M6TVh0Ug5+/CzI3bJGoPwVwa
IIZXkamVO+DNBMNmgjqJFNBqAEviqFhR8htkQG8e3uFfLPIzgSpdg7J7T/9wERa9i4v93Hha+wI8
s2h2MjzhK3Vorh/+gpDHeRDz/EnkVN46KXoiutQCJg0r+rag9MbqoHTgn4mdoMe+PNTI4xtV1spA
8ABZtndBUOuYfYpju2nOaMwkQDm0+rbcs7llIBirGc/pgqBZvC0ho4OQBTeX4p4FZcfbfFuY4jC2
H9NZ0OX0WW4WX1V6sIQM7tu7r1fuaZnCKRcp0jd32/2ce88uBmNwjBcYWOwmdvvDyCqioWJpSKJQ
a0Kx40zQWMT/23H9Rf0CZoPOkZ/FUlChnCBS8+8KcQlY0F6lzYKJMs/ACGx28cIqS2CcSiKpHD55
afY72dhcnI7Lxyef3+segB8B/kz3E9XJ1cZOegcZXfbbIlXArd15Zz0og8T0T8hW9UBEFKPHaeoW
4PlO+WJOv1v2V6mQGu9cIJaRSN28drVX27jOBNHEygxMAt0/mCQCx5q1STuPIdgZfMtDNYt/b68r
0M5SStpeiOy5UMlt5RRP16ig0dsNjB6k40jJLFhvBwgNeRlmv0OhiqdKcAE90Ft7RYB5dihM1RK9
JWFoO+DKC2rvuyxp6yuGjDyF4Ki8QCwDNvws3f2yvXubk1UiHOFjRQzKOoWRFKq5zIUZBinigueE
4A+//VgN97RAssJk2jECP7g3Mislvmz4Hl1r2SJBp21FS8a5DVTGp+DNy+S3JT5agCyXqnGrZQP4
W2aDUgwLlGXStZrU2y7WYmrrztFT8qzHT5SXmJ/FBugl12GJaPUaBLyVFd//1QvDcWOREbeWE8vB
sFh8zfGR5AWxcWUSXtPZk3YiZplad/2aHyFEbW0voRbKkSwZkJ43B7crC78GtLrude7OEL6HoLrq
8bt83cXsT/20/J4BYnfZRVv6WO6MDLn9flwRrmMQPUH+jwI/46XfVbqXmLQFjT5sFzMfL7m40Bd9
AMqkmAH+fN/Cab+wzjtMkXHdz/ayxcWpQkycB+l1Uta5nGwwgN6xU+mZvbU8BAkRwsbLeyeu9LZx
qocnijzAS52OSCk34t2ylBcP7r8g7bCYGd63a15YDm4PjGHXpc897Bnz9yq4xlxG1QJMkcIIP3+S
o9FYqI4Mic0j9VMnZ+a4+CtA7rwQZZLoZFfHiVC2Ph9qq4W88p/zN4grBenDuu6dxl7MX6V9tRst
2al/cJmCUpP957XXTYlJyK5MMb/yMOXA3sax3iwEIntt6wU7MpNS5YX2zORVG/BzhdjSpyMlhhSG
IJxTfzL4FKO6mYtVma+Me6x9OMbk6bdP98mz1pntzMtt8oI564P9YyEtlIta9U3Bm+S3OuWzXkVe
3L6hsg1eG7KKud692/xDbXr/uP8UvTRxPe8cjpdXbs/jZxP9xazPZszSHHXYy0Ih0oGuNEeRmEhv
4aofLJDS6qU2d73lom9ENjzWlEnuEIqOIxc6G3GdlOY5V3qcdhXWV93ewPXGNDcQX/i+jO51M0lE
B38su0UbCpCUh4ff9qqaADxm6s3+7EOtBIic0KGW3SePF/I3LJJnTyB2tJFc1eglTztOdbDba9OH
sj1glQXzB1DUMObhvLVqvwsuZckNvN7aKOgBShqB1wqvD2xnqJufRerKAgMAhawgEKOCqvvVFId/
6EddBGX9UCm4XkD+SGOiGrS7Gg6ah6LN51b9n/FJOBeVvXPb8kGIbhD2gctN2FFunjyfeQOuKNmh
+gagUBxksLewZgYjfuSZk3IY9VnQkb7O+36oQJ+5vcBI8/Z0i7hNvhSDZAjnwdr+KMpyV6Ayy47Z
8A3lBNKmdRe2dooHRiuecVraKXp32apclfHW1V8WTKJOauUf5ER5v/shDtSuNzDF+NPo8m81E7Zs
yUUG9RbD7Q7yiAT0j2vLvfMXEHhyhlIQtM9IePpDDmiMS63eZwNU828+ssr1wgQcUvaWLE/al9/4
is/+lRO24ttPgzF3XszpqBenOcU0eqmz4bDfPCuyASe/ilEb0OqcOO6iL5WabqC5HoZ70IreqxIR
rzyvNPw0T1HhZsEH5INJXzCmfz//EX3Gy7x/vEH1dWpYmdlEcQZWxq53vGIrELlLAvcBfvq2ZG6L
c6D8Hv3QnfbAAWPWh48c3hiRmWiAbFL8LPr2TEoGu4vpdxFNVsrPEeX+zMewmKkibEi/hyq5Jmqg
tLjavb0tlhPA6s6Nr+LKYl80TkQU6URtwOh6OTNA/MYZUIwUYnDpZi+EM2g3YUwoWG2kw8IV1HGV
4AtY331rxfqeCLTMCPvjuii6OcDzgbKf9SRFZ881xGpbTHrqS3PUK07bwQXnE07P1niP9EXONo2k
mnw3ty620OrtV8DXskOb8eXStAOWvJBfqu9N4veAutGKgRkrOLwISoqWuJcYv5/B99j7t9wSUMek
ecxbl+6Lr/V3OShyPAZ18VXgkWndi9XuiyyEqq06k8G0DxyEr7u4lqLfYF43Z8uai+xOWNhsOxwh
LE5/fq4Bw4xPeekku+Nb1Q00SK4ES4lAq5RZBmtD++cXg2GYM75F9B/KkKkJXK8q7cHyrcbT7dyD
Zj1oKuFTS1sa9sBApFntKwMCJLIIDrnOLr2E3DCle2VsigA5W4H0IbK8QTePHmqcNGrTKwiKQIST
POtC3B30ITbmzqNVljBqasdgEdqhlZEsnx5DAym5UxjR/gLbe5rQ27XcjakQGEszdpGxN8DZz/jP
QeoSb2qMuz0rpUTsXzQLEiXXeIbPUkZs1B1W4+e53/9EY4ML4GVp95KGOkgrtKW1yJwxbdP53HXs
os0Cu4wThyvIMfqm7LOvjeGUwDHEWKGR2bB2Ig1mUNPtS27u+ZkfQk7DGZV8KaOLQ2vYJn5vf2vw
U01J7liC67zQJMb56Dqvv8xTNqQTzTNhZzHZ/9Jwe4e3gNEHvDxkvbykBOz9MavsMD02xcPFbFXn
R6FMRVkbscCtW6eBf+rzcpz6OewQSoU4NgqIZ+26exiKMuU6jv4AUvsbCXp63u0O/1KkV/DcIBBl
6XRb0mz0EUk1wz86sl8LZh8QW2OHc0qPza8ds5lJ4hXfA+VulrN/05IyGfXaJgNM+9ZCXRKxym6L
khLVZmfmr6yzxgV7nNmOwZq8wqpeCiNSsbHgQOsxVbBsLaggo6Cvg1nIxKT3piRhawU8yFGtsDK/
bq6pyqVPwcJ5TbeulkXur8hM+9M6IscDofALXJ06fjrSnqjLZX3XpXl4nnHF9hbI5rTRX4C1WhU4
wSZh6b8EPwalm3fY5LrtmEgLq1I8hqs6bFokiHVyU+HOTDuWHkzkhV1HsAMiLMfk5tx8HrX3osjQ
NY57RDTrmPRixU+zONVWdia0HyRyEYMs9ty3l2rndX5fTQ+QC1sSwi99sPo7P3Xuf+j8b+690rTu
vD9rm3vbujOvQLimoGib2b+PBXsWBZO2cRf3Ay52u3Wv5/LRZ39wmQUds/79uyzFp38iiQi0gAO4
nOBwxbZSfnSDWlhj7YLMbGBXLhPjzdE+R4q0QomQGnUE8+jjBEp4pyCoqDzzudjJAaLYohqU1kwe
5DVg9gcZdaKBYuFc3JRsItJ0f/OVx2nj6YnzHYHH1SwuTFvMmmbsf5OIDDo3Zx37MHDhzw3Wpo6/
mql+G61LA5P55E3tEnq2uDoSgQ8Jopej+Yr5FqpOzRO4as4FAxq5h8JZJQB2g+3RlwdGmzefCjlM
mXN79BsW0lfTi2SvWadseBNOCjrOClon0HlawYitL+lSkI/3ZdKPaJX9c2g4khsIwiLERrW0sDEH
AE1ydNipZD2yJXCBk2tdu7nrlI4hezZZOYwUWE4tHeWcVJFV/hwU2cTchPdhiMkgwZ4R4TYBQDyp
Rn5uYcGKxvV68BIb6wgbFBpFDbrfw1Dynvjx8aroWGktbFq2gas05w6joBpR4cSLlFRy57eSKPl4
Gyi9+jY6DnjCWCNlsBO3YCn+glemUCq5j3JT/Sp3gRiBhJdrupR4dns5REYPhcW17E1xgTiiIwrI
mijVv5SXGuW6ahS+TA/y39IZ6vLbvV9b2/HhosBY+Pl3GrU0aKt+fR+bG0YOs0ScCZIaGjM1ViRF
22MHlUuE/YU5SFRF2QFC/hm0XAar6+8aOkw9uCQESs/mD7v5rH2QhtSqEpP9F1g2MkamZwEQqYrN
DyD/EK1K0sSWLvkV/xeyOUJcb7Ky8gJra53bpIIO5tHHQTz4K0N3WG9b+zWT0kN1PpEXMD0ByrPH
mdLVsVkyy5vfIQhIoDwySyIYTC93HpZ/S8FMJnTGcPvUEIWjCGhz/v2W/XQhGhEZQN3OrNVhR8Vv
HeThZxfact44fs/qJoAKoX4Zi2n/51tV/FfL7YykBMCtxF7xhSMQEewV7ZJy/qQtuDB7XMwAen4q
InpFMKHHiugovfxPMndzr2SYP+wTjnhaBo5NHUBbbp5e0ShCKiDm4iL6I0FNv6wi3snUpLymlODT
5C3V17BSMoQtu+yhnTVL8084SQHoZLO2JBgCyRTsSvMFvizpV+7uf9kdogOtVRi4KFKtELHfsR1V
HCd+DEHpTRdbvysdBSckZWlvdE96UuQpZwt93lRzrxQSiJbenhemfvX6w/traA9hiB+muUJ5oGva
HjLK+pPu5/Vq4gG068Cwp8rEeek6WrvedZIxYXkScEySkBwYLnB7rEcCxFbzfe35fPm7RLPuzA2R
2omluQbZnuWRuGWG3DcoQXgfRo8LjiE80s+gM9nu6ljD4Jn+dHZ85VJTOz2YNW4GpILr3N96WoB0
nBoHvesolHwS6TKC1K2I65ofOxuZXanILrQirqf5TdAtZzz9+BCycVkGYmZ2JgxT7AtZw1c4x0GK
WkCTMwOi130JRw0N1GnadM5m/UdhXidJTjVJt6j+hik/dwdyP/lolOTo33VvohLiLcmtSenD1648
yv9rn6EjbcdesK/vgn1K7I1I2S6pVK4y7cs8mBrwma1odV7/Y77aXLlBGB8H9ONoSlWdECswaaGf
EB1FoTdyKfLuxILGtsQRFzyy7VVOxpkJ4F17rUtIeVeKEH3XyLhPQt2+LaiQuDwo3nqRFgy19/85
ngceL69fa/gPmFRL480Xzs5yEqMxiUIrn/F1TQ0fCE/I8+atDY65++lCFpoyuIDZMCfgkUV+adff
jGr9WmFSscfTXus8/ZO4joqnxvCJBuW65Uw3m6JhRewJAVsr35ccblhzrB8mH8f6f7yfAZKLumXf
nR8o0ElqQmIeZjQY4KbUb/vptVz/rcvtalxNocxoHqfXicv7PZ1uMx5Z/0J004pqJOVqVWdX+TxG
D+QDv25y5gxnjSy+6kJftCV1ifZdr4oA6oRlv69Se/bX5D0O0qzl7r6qh9eIlM8SZVoOkkXncq0W
BY5+w0HCoxgnvwBV3UvwhQtvggEfiYGyRCM3PY4GIItmevg4FWGRZf2VAk3mP+WbuLFbGapAlW9c
wpGRN5rUHDMelX+Bi9irik37PSpTnTh1skem/hG6CA0MGEdQgPdJsxm7LQVldWrF9rwpUu5rYmei
rCdeuQ1/untE8Inn2yMtLmrI/s9mY69ZUNs6uVMCeNDiOclfaStWaBibMrSxzOjTKrgsKJkOnPxB
dsAXb2MrdiKcgEiVgjhBM4W2y3ggbrHyaHGJeSQfdmvCErZvrtJqiZkT4Ys6CF6tfD9CDWD4RV1v
B0JrAnOCfj646ybQbrVBMVBsYtZ8EX0hylyFm9owGk/KrZW0G4nfilw1WoB8Ka+mnQX6mQ/VMKBI
Zur+MzoUiV/vxf9vzfiDzfq9jH4Qusl4euZsfgSURCGn00r4pLS0rOyU/JfrRnRAdJMnuE4IR4FC
SJ5EIGDzjn8gICe3C0RN9PrGru7gdgdGZ8Q0iaHLU7Ft0Wh/eQ96/fj+qOTxZT+Th2u8dxCovDmP
7Lsu+h5j3bqnWD6ZodOOvcc2qZ9EUXFfKAYsXA6hm66mXtT7iKUCDxjJkYNHbNFq9Ykia8FkIVMA
PgB2mZFnfAd/zOOjjP6B2mATVZkLbR+2PkfoundrkSH6WqOhQ/9Enovhh6TTvbK2/jwk2UReIK6a
KNJIe4URC8dczDBBRkMcCn8hceDDEz87bhs89dF3mzpRX3Q8DJsWt8T+kk8HNDrsWNmnLtm3eMRW
qoV+M6WSO//sFH5LynwMr9AYJrWuB2afBudnaNF6vSwj4ctVDDw7jnIWnF87J8rf0fsCSGiihiMs
AMPx5LcXfLOWe2z0/tB11gmFoub4i14btKYgL4B1KHs1GkaHX4LvRpHtKrZQ8xUyVEEjL+RXOtJM
RqnBggc4E0rnvmObdHg/l/QHR/Ihvso39nwVOHA1paNd8sSKo4uG440vSYDM74ugrthFRR30G2V4
zRq/7gWa5SkPzJEfwhXeDjBjsHBWkxmhNsJNeYTKPTN7jvf7v8yK1kswAcd4XwQDqvIKwCVtQge0
ujfMlAr5yPqM5xq9+O8Xwwfr8tpBNIXTwbBfRZ2QM5xfWvkeLn5ZTPvR4AzZtXADcwq9wtumNtMt
DuaYRJ+A2fwHbgf7UElNBvcLwroKiZzPL7v3/GxuAZ3seh6W34OSXUedM1fcL4T0pZeAQf6Bc50y
2gXG7dQJFrCPtlpsRdO4leSNiOLFqeRMe5lWBIbwAtVd1WZdEaMhD7PxCd9H66O7vn9dznP3zAYM
XM6sIq9lmg2k4e7vUplcsK349zPtpNqQD2vr1gI/pCxQJ8F2UQ/kZlzAyLeCd6hlKmOhS88AgVwu
5I/ze9cMtCqX4DLORQtZL0e06WJBUrG/U6NABIZ/q8DMz5eIO5lOE9AdruYldCGT9MjSLl2beXgz
SiLw6b+p7joa9rmHGAw3fPiMHtP1GvitXfkRpdxr7sMAFPH+2xFBp1iYzS0reKaVGQroS7cExlOc
xCJuoS5WKvgHAhdY0rBzQ1XjKC3gwBCt/RVLSsU8oPXyYl5FbDF4xWn01M4b+vUJS857XohZ9/3A
aqoqWnqJd52hR9HhJbVIJmG1htDjz/N++4x615TZl5dfsUabC4Cx54SB495Awv3uJlZ2y6YqU7ie
NbVboy/sEiuoUr8q4mz7WY24kGvRma/x5ar3FUMWnHerAaROKRKHKgwzJ8gQoxHcbY3KXtyLjVTP
+SgNyarsH8R3in8/2EZE6ymKCYjt83ypKV8G2H29R6/mTE6B+025O39HI5rdr/tSBcQauTVQXh2b
0HppbGnqhMz4BFU3Rd1O3M1/CiUeYAi6oodVwsIu64RDmF8lVHY0h3xjsoHDhtnKNAswt/p79Etw
XVbWrvmQ4dfBNhnjsREjt3vZtj9WCJsbKmPVAtqfJ8fXHLyAKdZwlVC2oKpBiR4kKma0qvxnUQH1
d6AgCAuVp4lbqyhHrfcMsBegL0ODhvZg7ISZXCr85Ifwrz5LiX41UGQosKF9kZ0+NvySHmy0u3hY
0pe9D5tRFl+bEGSuiImTswMc2/PEU/WkDhOLxGM1bFXC5l7kpE5iSyaemN2E5eSdk8EeUzOw9f2e
TpcZy4PXOE63hiJIiw8meMAat/jR7l4L2YSDi+TFyiV9YQsqvYplRHigpntn1Kc81gXCZqyzUDCG
fK1sgArUlxWbKK5Cy6jvMKgsPfPxhuAhT0NawxXjn7iifq/DapvXgjYzGYclnjEuAP4gmE2pu6C7
1+jSh8g3pHt1M64+tfA0vJSlxuUhCRAPZOLvDhHribwlHYnZ0jWzdiD6kTDMaTMBLrxOIgtoRLso
1DHrajUWXK+4I+oLurrdz0q52Glnuh6lETACgZ0paNcBa2/Oo8hgOfbxXyHgMSWehTWglgnUwTl1
POR8axPHv/82puqjlthKhG+YwWP3VBH+D6Pk2Bf0E/dFB2l3KpNyn2idX6L1qQrF6+SkGZOdILoO
/BPPpROt+6mFfTsy6X4mIMEaVTPkiqqObumLXm9zaRqTAPjdiSif9lx9NYf6GijcSM3UQ2X/OCPd
EtRddMGdQILbTOJzkvZQtMT4ynNklIBRxxDplY1mdb8SDuJz1tg0s8uZVlv+5JEa+WiA79PJS1f5
RTK349OIlvUf6SBNR4EXq/XbwaChccYutIF+zhz6ssNx/egjbg7vrvm89Cke/vv7Myz48Yz/Nl1M
U3msFkB89ZWlePo6g8XV0zLyXF0+RyPUni/G3JheWU8G1wmiGXxfacJF0b0NdKf39gnqs7eqeTau
taVzKvFDww8nSufc/UiliUH9R5X+PEOJRs2efwasr9Czu0qnClEwAvMI7IHb69Q9fCCAjANOGg+e
s8vQ+MoQE3GLeUi1VYZ1GwECHQyJP31Wt/XJdo+ajQVGoOg5c6VEZpZrRWP/pTooPVbWrbbXQXai
4YmPGmImRMPdGfMktCWZBLnP+nwzsrt1dTERC93Rges67ammM3Io5bdojw9lykThmL7kf1dYwt6N
C7e8/hbjNZzBAFZ5SY6vWTC+mD8OrkdmHZvkO1cNmMG8kk4s3yaZ1dDh0fXeflLc4iUu90pcl7/H
+nCcgmAV45gJ5hijMSbiFpVHMNpksIN03knLzhuZQvlKhyttwmLvyVxtjOhWGcNUFt+w66lD8zxZ
Z8CNZrf/ToOIJahanlvg6izu+TxSEKYL2eLTQi5hrgKjF/Sy3rGrw3KDctm5H7fV7uEYJYK11ejw
dngByMXGTvhv8wkxdlR9A/I5cKke/4PY3P6LW8pBr8cvLixA9/ZU1QCV3SZ2JmrCy2eVRLRLEHlZ
HqHsEoWeUFZRdcrZAqF2I4AOiEGlHgtBbR6bWdQYTmVGGRtBKRpTP9qbuMdIt6gqaqyOrRCh0P0k
bY7JSxCyO1BLSCLXZakcrgm0wW3xzQbelxRSuwcUKj6Hj1CS7semUcCX2a4yFMvQOo810qLqtaAy
oxIesezH0tAA0/bRJ0yzEfW4sakRW8ev9nz0TJxeTTm3lcefCaw3AEBYuDYelw9yBEdl2/6D1FeX
326egGPfRCmr4lPid7jHsS87ocaD+UziCuKEehmvjxkiF4YKuqcKACeae+bdoPdIEitzxvydmqgl
gXPZcbTgJT/QbkkAO5FJ6TE+uoduBKsv5SsZGOce58pTFHXsuasCnMHoaISyN8dYJEkAjQX5jXgp
KjSanjA3HRShOVMvGqw4LA3gBjk2DzdwZZ4gJAoI837+wlgA0RShUu065HwU/URnkQTzsKtXMIAC
KmeISR0hdXfEr2O+YpX0RAVLmcXzl8augIWHNmYqFTOgogT3RsKU+z643/9siejsyosZud4nb24U
uBU0ZqslCUpw9EnRHFu8H6epMe/yvpkZqmdsclilRDHzNxoyeE1zPVZuAiN5o4BXynwXSACnvbyX
Y/xA1EYGJKufr6kf+gt0JQ5g8BLfSAtDb3nEkRklv7Xjd57s+wPZoScnPQbsagtLHZuaA5jGl98V
6icDEmx7p0hG7NizzEptfJLARr36j5JgoYoSXgoqQrXPvXDc29oKk6hZbWPC3Wr5sj+KfhYaUk+/
dZChqFAT4S1J4WgusJ/99m3Lu7a7hpptRcRwiFVuYjkdGnMAQqvOMznlUMcth5GC91ylBBbhXUSm
uxjMXayZsTS68vDoaQ+TJGcG4GxezkcLn50bEflbn3CEqDy3qDRw32Yctc9wyEwAnyQ3pR3CRtKd
iU0U7qecm1Y5cx8iacyUtmzARU1kcR8Cu1F2ZTb8jRinv5fjCGiCFdDqAkAa5SpR8JjUkDmvxK0y
RSqTxUA9p8U8vGvY26tnL7Cr8dwjXA0pSWsktpVJtW8MkrXdowNbcbjMhBQ5i4nFwiecg+il1hOu
vNB2otni8BRU6RrGvyFSraepI+8llDaZwem4FVWM3MI/6yLIePTstEIWbVExUfKtzVPBE2BdT+Fi
xSuzWNSHnmceD+nbBfBO3ufNO/sqBQCfX6/qyw2Ug/xnt3LioKmiqDsPmIYWRivdU9MpAWPRmeFo
C0eMhp6QF/a+nBzjKo8sese/5pXrn+WsldegDkitBHMJIbqyKE6UTHuwfzN3jC8Hvy+QgVnnofYt
wUxs6JkayIiWSxt8LVhbi4HwtTflIaBQGC7IWP5C7sqebbMRl5MANArH4rH8+Y7CCNUoUhpARbhx
9P71HKBWS+4fxsnZAOWy5YceD5uRjV+cBLcpbPxJSnoPRv+F78aOM+IuCYBkel8+KK5eMs4gvzR+
p/Nadq6lAokFWIvPnspXBCuebd0Sg7zfCY37F6R/398tsZJB7vgmiaX6wYScot3PfD0xRYFPirqt
ksx+Gc8olXSscDy9yy3W3a5/+dhKxSrQaVP5ewOLP40i5jeD9CHlt3WLNXOabY0CvQ2h2Uz36Ozf
TBGZj+5lFTVaunEuYqJ8QZXKbqW4SKaHY+JWSgUeTWTlssogjvbyu9szMcEFhwhgLPQev4Fa20Aj
DT61VBI9ZcbUh547MfuU9HoM9xMqPiPsPBawn/5fMoECFG1H3vMdO9+/SgpH5vbrypJZW1w7E/r0
mJ21pYm/0UP+8DG/b72UH5MixTuwpeeEViZT1hiW2o+NhTe1kHzYRmjm/oV6qq1wE70lLR14Ovrl
0SNtyaFLet8/VgTsUTycBq6u+D/lJiVr+u/dxFT4+/bJ0n6HzhqaxcqoGTnMqlQytCM82TM5KVAt
eJkt0IjCCwQsVNeBMUhWCbhuyg3Q42PeJyuWMT2XjGOMLRkPM30QwNb9CAQdpWbmxtWBPmpFoRNo
M8Nmuq/M5w5vAJb3gXIuLC9Bu5FgpGRgvGgX91//e/Fg99b5BhLUrKoq7SV4+NgxyRCzSzbUw1cy
HvdZzsNKqew5+cYay4tRXUYPz8baEliwWakcnUhNiEszGD6fRvOQKtcbhmdTO9JDIydvFYF4dVM5
EvO0LrM6/Ah1/XrSEtb3Dy3VHBpOwQtQZ6kUcZ7q8NGHTwVWI/TJhAtufMrPEbIdEbOQMenXHhCW
SWLElRNvFE9aGptGa9tdgBv22PN3RtqmLhxafO8URMClshXoFF84OfhadNneK5p3Y9XK6HpUaG9H
MtnojplwTXJrvyHPTdcRTOYFj8COol+zz2Cn5Xv/A8QjiIcl1WD1me8BDaOg5oWQ1a6akj0aBhD8
yrc5U35OBg8umyl2xBPdbxiQK0lEdfOajXUPg0gUQF8ON82g05wdbGdKcloKhhlaVNNCYl/OTGY+
whCsCV3bJxqKzCVQLbzvpr/dcIGwU+yHL5h0JZn11f4DC6Ng4IM0ZIZQsqKxrfC3xKMP2i5a7iwb
LtZ8MPCqklonA3FidrZh0IpOOl9xeGRySZ8HoqsqcJowuwbhWaElBaap2D50b35ikKZNOURMtFJf
9VEkxG1Pke9HELgAGw+QIAYwODPvP0+5kItIK7wn+P9pnEe8oyVs14ZG144TuTAxcTWfz/Ostn9W
LKauNZ+QTrM7lwb19lotdPA4dhQL5Ik0OCXm3e9yXqeLD1cS6LX63DcBo5m+byiNGUH11HR/cmSq
QOEjVdrKYucJdkUftp+CcqCGAZqYV8nyH++70HQ193P/rO7c/PpAMVuQTyaD2QmbrYYG4ZkUrJCY
H3EXeDI8aLv9bT66eDRGeKpQe3eLkVfDovRF3OW1K9NJy8JIwexCytzUgnVXGgF9CiQUkGn+U3f/
PSKIwSGGEWMD8xv80ftV6nfMCIBApXxiRkMBqpXkInT2kW8KA+/bl3GxW9d3I0XJjvIFB1jt8R8y
OjW4GBimduAaD+c95IQhf8wRDeiCuth3JhmKQ3D7uPQd9v+pAVccczYbybv81edA+OKN4dMhGC6Z
83tHvUCfqKiyzi5hWirCWuBqAkz3UnLW/QHepX5wcsaVQPmh9miLhrPdGdpt+w0EFxhV1cL+crR0
RvIh0MvyLhV4VVEIqOaAfwdQHiMJNpIjo4UD+r15Bqo4fO7rQpClVQnRcf7hO5eGPKy3QHut9iPz
j1MBfrer0/RTwelAo8+BYT0Ta9Ar6Scs+FaJSSmaPlQBGefs18O/zbf9RapRNhTkxZiJuSCSoJi8
XtZcO1cEribkYZjnqWJDp12pXw171PLWnr6kKNqFDznSL4GBLLigsJOJ2WpjVFQ1Q4AdkqDfSJe9
Z75ombq3VaEGdHRujRkbIpQ6sclaoki6+bdbCNKC28YQEQVcSoxqkJ+6ziZp5h94/IIg5HCiKqXP
ty4FVNLysC3gYUVkMyXZfWX9dyW2K4hKcba8g+23QiVLPcBEdWFRx2ReRjINRaAzvcoc7azzC3cB
EZEszQMAdqxmGMVYe7O2iDP4yDWjacPDSWdWGYiXVhtIthpQR2e6aIyNN7fvfW6F9yq7oCIsxCvy
XR6+w6bPOHAxHPcltvRhs2cuFxK/Ohsy1T4FxhsnVIr/stVq1siD4BQP42lL9oFDvnb4PAnHhESX
huhpj2+tfmtoIrDQGtdiNV7xYd9Wb5+03Su9iJr3xx6h2170h/SJQg1wbX1lxLS+lqW0uHU1d//t
a9sl05KdSPDhf4rjbag2Hquifu0A3UqpNBjkKFQQxDoVjOmRHRGn19qX0PpSkI0jFqqVPYLRg3vY
gGSx9hT+uAaVfquXIy3gfUdTvAM/Hc1uU3Xru/pC1cfWGIrJO14aFIFuWsVfV5zyuJywLSvngyBz
5sYo+D1N1X25dxQqYzVSva3Xcysd8mGxOZwDsq4861iHfch3n467mB0/HNui8kcW3EhKDuxUX5vj
fj0dPB+igXTlJJbhV8Xjuq+ccLrG0hwp9DMIALgwQ3Fm10Tp2ZINl907J4DsiKG6nhLZJdbhhASj
iBYJdbuoWt2BBhYjiKjvopoYmJAbekM61KrZ18BL6VM5d/7A3ZDQ1Jznw12B8MfJbq3uHgqtLY3F
AV99NYT5hqbUoAtm5I/0D+eO1UnM04nXDEsd6xT1LS83NDfhPwxgyiHUxEtPflYNQVOUD22X6AxU
x43llSEV6e+NXw1CecH1gc9Dy2mBH70qX5jjKj8p4LLbwr8Lfu5uPYn+0gHtDyGw2e9njNKJ/7tj
RaEN05HweahHTa8uYCMIuifxggelh4b7QqG4Qms4crs4eFiKo4yZX+dJmaKcz0/TlNPYCFvU9X1U
mGdge1RCgajr9rSXwUN/U5pC3ACUeJHK+Zg1JC+vss44O23YEfFP4JiD81LVwSq3HW53XRdqBZS7
zwqKy+C+qQUgCSc80pJ7fDmk9PvTaH75qr/HM/tVoKX+ikPajbrOQJvGEhK8WVb0mUwD+tWKlZsg
IQLVSYcHa6uIcInBoMrKA5OcsGIN/ymcfhisFwKa3e2A3WJtg0z9FK3oqtLscvuiKCd1/Bgz5jGt
njQY0D5jFNBttiFYyZpTWmKvheFI62KI8J6icv269CBCnD7Rp8iXzRt6uqHIKf/tEtxGCrPkbSc/
xFzSPY8I3IuzkwPZJF0cHFoYOh4mlSFPMoq3x6xE1pkrFXrD+MJLh6VAQSVj/mx8ZKrIX5niR4P+
MO0c/S5jBF0rZ+0Dvwzf2R+fMEZnZoTBtlXecQ6fwAgEq3CR7/5yyiaC0pAdrf65yVFX+a9/0cFB
7O19+vrPqYAMTosXmJa6NNLdY1hu2Kt7p7Vn8dfbPBFeZ6MX3dQLacXeG10/517eVRNNvGctfcqi
FXerr1VkZ9Yp76bdH/M8CvSys6Y6I+RZxhFiBrJw68/QNKuWDSn21W09FRh/LF55tOzS36RKS5dw
VT9982cbP+fIUEDLmRoRtX4Tb3ZhNTCkZ155ksgV9lU1TjEhLrJFCFY9gm8cGf2gO9f2c5VGz9gE
LaEQO7kCe6kkQMjdSbitSW0zJ+pXf/dAkhg5MxHrO5mVu4vGTLSVgNduuegYCoIsozephILXAMdM
cNSaz06kBgU9aokRwJBbsyecUcajym6FATzLNL1mqWgFA2AWW2W1VErmn7N0LGFfc3Q7QcDfCPXz
amgmDcX+VZrA/pNpsLoIGf2j0qR5lndfXQHXqUIJFofDOWB7RFMmbTu7wGQe7oDqRb2jLGfGehtR
8lnWgZrjpYds6hS1VYeZ34ZsbWNmHYa98Ge+f0N/zzAOOig5KbO+X4Pcd4h3sD1gF5keeStc6ksQ
3Fc4zuUqKWXoBOOTQ/cAWqrODocK8AIKldfdmZ/miZiPU7vqfLu8hL3sPHHzQ4O8gvcqL9OOovVw
AEYMa/IPhLZ0Ef1T6joKxtEQCVGbxns9kS9lWBFbsQcMnhRIyBUbKFP55nM+jG2uNsBnxFJlWnKM
RtvUMVeGkTKg4LrIHq+yo7QhTED9E/0Jlv8vK0KB0wQIUj7v12ZvvDN0IVy9mrrxq6P2xhygGH86
DsSx1tjOys668lAZnh5Hq69WBq1EvF6GQdbcIx+aUg3938SRHjcEH11xaD2yFZZsWFMnltYGYl7p
T/Toyx493Go3+wkYf9bscEJ3FHiAqjmHZh8JX3S9BGwS8OKgKfKt22ReAO30156jdgYv2oQQ46b2
XiKPWd91+ExRYQNgJUr+Cc8Cj6t0C3drST/Xw++yDDtICdKISgYtVScabaB8tKhaOQlfrfd4f41v
s2vxNmFoO3GBseZnVrcKet/5EWTQjck6AKN/JMe5iK41lro0oNfyAmIJiuPiEPFPbIoBzZ7gcR8H
sH1u+3T1EnT20n1FuamjcX6wH7T5nt+Ne+tV5EhKZapFpSqFwicOX/vmmeq0irHyAf4h0eewCQ+q
lKbDrr0aFVWl6YzkgeEN5Bu5IyPv2mR9eSFmPpuMKCWKNznx/BKtP17ha04gzqQrHbSb6SJqKfMp
j6/u34BLj64t6vTMULDtigCbOCHOcYjkBzm+8Lf1Hg2bwSU4VzZEKUUKSfsPOo2eQ0nwMf7bDT9c
49cZbuFLYAMlva81ai/5bAfS1EsdqjQO9rVlKYjV9ELDFxm1DvtaSWudSIuK8ApkatSDHQ9bC9qJ
5FCrxJgzez919CF1Jv6+PL3uOTYN64wXrtSyj+rFcNj91Bkkb1ATcEsttIzIkYn3IgOx+/CS//g0
782k9Ou5R57pzB6+111hN5R7+wZphiE4fwnu5FiFcoSsyt3b0nHed9E3l30FcxVJQgjVvUL/CUb2
uLMyZuENzDqhhtXPbC+KoeOeXTicdlb4TR3+f12+BOl2/yEPN3iI117uzllAdVTaDx931ueQTqY4
qr2MdBSzSJZiMU0m7uquUB58rAb6YrKZRDs6/DETEIAU5bZ015tLsqpMzdmoiTyLxoIbWs9TBE2i
kX1tbcty34ux3JGW//YlG7ilj2ouZHctCe4UNKyqWc+n3Y8S3cd4hISnneH3IZz81U0Zm3acYqCN
5w2ASIWur8rd4xjW2Z8orntrxNXH7NQNyAxIH8sDj5G+7l4IMS1KkFy6ASkxh/gLQFjDMrDbG0eB
nuQt3lxUIvKBi/CdLDCHP8XSqm8N2L/GrQo6cWyAIuHhiaP0ChkiLYPEFYRQVwnQkKkWJFS8Prxb
TPi4aWJc4OwIFEiKDm5g1F+HE5tL71Wu0ej0zedAcQnYS12VGgWCcVoFqtsg43cLsBTI33WqX0kc
YaPzBeM57XHAnp00HmWlJQ0GiBUnVIzli5tuDJtzasmrvOBBuI4YeegCtankRP7HdhWrQlEUg4Cm
E0mS6xdGKHdVy0HNZ4qCk7PtI5T0/o9bzdQRsrjBL8ubh/PgY/gIxGjXzLoMSmlS+RRE8iHO0Dif
BApfsGdvWTKBvITMY1VdkJtnYTxK9WQ4nJfOZ7DWyiDxWYTdKFT6qku1tviyvBfm+E9lbjxcBWDr
ThVxlWpjCNyyaqQegVUr1wJYdWM50ZB2AKdhYLP9s1+ZwGD0I1L7BOwqwIAdSChPop+4i2B3A/EF
2OWuXkq/tz4Be9ddIhOzuM+vdvxghpjnIqBEYL+X8K3Th2YxXwv0avj6VuAT6W56QWtiaKEIFFjN
lD4of361tEh6MDhZpztU90ZyRbDly2mT5bk1B5/i8i2oiC0oXykf/PswPVW2otzPCA91Iz3ODays
Mbn39EvTwEhaCtRqtdYa1Gg+4PkB4UmFRgbCX+Assedyy9G291FJr8ZDPMA5E8N/XZCES20eHSsS
yeyLao21ahjItF3AZ+xh3fsIChrKUK8X3CUl98Qq/rZ+hIBRKGSTRvikfCJygLnwheWS0bEYA1FD
RU01bV3c5/pDdkncf1drwnSMoQlDQ2VcgN8CldjH/oWPpRfJdCpqyaKujLpKgj+elm8u67n6SuGI
Wm7HayNMsUUIG0gS4sZ8ADFSwAq+rIjEa8KMcT1Plhjl5+kWsQV08aPcJGYQ3qdmUJc7GhZ/YAIO
BbjsqqerfqBTdwbV8kVhf9rUvDG01JWvRcwtYk7Ky6WvCGKI5ub66N8C6iL1xdUaoM6jpeVtnAMf
WnTVUqgXTH0IXKcNc+SrxB9VQz4xkMqrluESTbB08N8xwouygKpA+3rX7xDw3U+ysRUr+SseGFcI
YQ+59sGU1hGyhBW/O9PQ8w/WrWyw/lvcobIcR/KpW0lqf8sPBod2Y+yO82NOT7jZShtmobvX2sFW
8gaOodn3sHmOJykOzQsRtBO7O9c60KYfqqH8GFSHT8BKMXH75CHMsz7OXsYHnKGu7mpd7PMH3GgC
fo4MWE5ysRTQGVmmenaP/X4HfWF/J7NFbBCt+qKDfbrBOkpafQhc//F/+O/49m2Rz4bS6nkKcwkj
Xh5ZgP5s9Y2rpWlm+Mter1Nh1xqVcp5B2ACdJuPHBYiV10ep27MdV/z64S8YHITSaO+h/wbEAojP
75RukGS+LUxf3LjicKm9TkzQnOS+Eie0FbV2pJpASPW+Wrsa3LkndXVuoTYaWmq2WEF2WrHeJ5mz
UK0UKPXnPzOobXSSoQqbRKTezc0CF4xc8J6LbNQHdiqccrurXdiuIlVZywmZ3jct7vj3JZN9Scqr
6KOjtc5+nNsUFTwuleZGnxdHi7Mq2sPjGMhgaawgUwvx222psSz/uu/cay81cYfhG3jfXtHtpB7V
UJTj+KzqOn6WqCKzCB2Yqy73RUXu+qg6Xo3az1Sp+61T+3s6q+QGwio3wfrADGypaw6lr+1ZvVBD
2EYAR1L6AIdIIZ2Bmto+2WDYnZkTJae5flZvZq5/vlTrEVJaWqUWde8EFeuoSkAnaCiZqpxPQ62t
IApnsR0VSPfKgjdlJIYz3oERkRVezlkm41QA+0K1aM6+l1rGwWZ0qNItgww+g6zVQ3qWVJMciCVt
KGnUoV/wlOBjkwEu/mtzyz4xd4vpD0yGcXA6CgJ0hMssa/m1nvNYRoKi9+qZhkoQSQ4yZhGk7s1e
DWzfF3fn1/XywUtSugXctc0rszWiBPyT1NxBCMmv8jtMOpbBelEo3pnEYcDJ1ZqxT6kGWS+nwEgo
/J5MG01iIONwZU5X3q7D1ZvEWzowdBKdDXs4o2ySp+7UYUfUhqANCOiMDAI1KaPvcTHkSOHtcv3m
M4mN5kWl7HyvXHwx0FMZvOdph7AY7IfE3AboYm4c44+e05C/NBBLrzRqRZNOawWy8I3CRSuOjSkg
/JkIuPEv4WXwtUTkDjwWm6UUXAOH7uOudn0mksz7TiYTUPls/1NlP93jhHpQaH+SHQCZEFuCXEbl
+WyuVXT2an9AqgP73rLvbZ2NURYWDs0U3Ng2mIrALF6IH/iI6chRcOyfYsuLRlPKBqhkDF7AaxXd
5iwDvdVs1agC+yxefQfDRbPEdwyLtiwy4HRyt1YO8tEiHJTW5F/+SYI3if0M25nJ5yJVsloeFG8y
T6hkKun3JaNvFWT2NeZKEUYt1FgKJluy516HUhnY1csF+oNThPGKjI+teVfgSU5vAHLSYAwdtWsl
a7SEdVIbkZYWd0rmwTdWsOE3sZjGAUc65KzLyFPx4bPTENGX5kHPbPK/KZq2qSOh4+V+lyQe9S5k
M2gk03ULN098/SfHu8tAUz2Ae4tAnV8GFUujJvdNhhWI4URRvuQVnQQIasuKX6w1ux9RoLcquafW
YPdUvef/mUWRQKjMVdQpCgQdP/b54fs8Si3PDTN8VTbBXFXlZ5rWvAH1tnrKB11nQoHskuo5M9xK
UdwXF+sqwp8uAX+u3CYd5KZtdW3oggFsGr0MlJ1C7jJmK/l7bMkvQA33FkRLxAThhg+q8zGGZwTY
sHpPJQ9lJf1o/70cGoByBMR9CEo4iYgyeTnwmmXzfKyO2uRI4JmEaDnsGVuJs9Ggi7pcohibAJDT
IsI7ak4seVIxl4lKTkNQmZN/Q5VpJcGM/njE9jsQ9EPhte9aZIjdzWgiXwm587lxT7QN8VXWw5JM
GIVuMfHxhuia/zhdjxPQdcWitprJ1ruPf27p/wHDxVLUgS2zlQFRu9Z6JbkoVzC6zFBrSVFVNQgk
0/MDDnLnF3EvluNNV28T3SABa/ui4fNKbpoI5B8BICrfGtv4UOL4/zBvSb6Ua25O+ji2/aeVRp8O
LImsSKzMjJCbsN53Xk123FO9nvPrwbS/EFkG29EJKr7JB+zJdtNnawXpd4WIJWKAacOuGHz+pg7V
ewLfEMW11qTr1I0ZUxh5qvBfsFBPNi2SjHdSFk/mavrYQQzREadPzLp7O4XDk8gSwCzzF6XWgT/u
eZSQ4iddQRY8N/mEGa5RHYgrNs1agfDvS9EHKnA7bXrwUc0Xoz0fZr6qWzFYUoUumR6KQFqkEjeX
dI+/lSlZRI7GtY0BKbe4eE6WM4SH9iat9EUL4QvFCdLK5mPXaFOphOrz80tdiGX1k6UXdS4uVpUZ
pd4mfLGDmI0C1F7pztpd6o4MoD83tl4iiPBALeqGkODEw6mrnGDzYoSQFAYI476/uyJ8acK9FrBV
WbrpS+/NQitaQlRwxbGICzX9hWk6xzCZ2g2RYfdlXxuaaX52sZiz33y6At+l6qGWsYpJ7cI8SQ28
YrC+Wfe/iuv6AwF7LNHyXqaxL6MIiF9Uwfwuqn0/CVLbBl8oZSmQJdsMQEhR6XeCU8VZfYDLKHLH
tpyybYMPYruyg+l1xj1pws7xC9mo/oEWnLhXHUJB+8KFpWnLxHNIr27dtdcxacTnbF7tXEWJ8ZLk
eqArHfDpTzBQ6i8zm5BqF0LiG9aTvnoAqajG5lfRAaX///9/7drhiJ6wJMyPUxYZGBVftz4w1Zoa
zTHdO6GlcQjonSm2SanU16N4/DtmBfOChISnuLwWUYcNjBPPaR0JtCCGHBDF7cm2lhY3L8AZOT/T
TLZ22CVk+U0/JSjOQopgPzJYOxIDVqXQ4rRJcy8x0UeKlyroszoXu0B89FJ8R1ui1AlrdY74QqUg
6N7RqiMXbS2jY9yC1q0ub99M1KRL+v3d1uTfU/WuT9X3DY/IjCwwyi0poTMzn+ZhS0VJICOKbMSa
R+g+zo138IptpBwL79xt7xdrEk0tge54FgzWFjxNhu7lhZFgPbd4OJ3TtwBPqOYvnE9Zhz9uiJhf
HIc/DFsocg4fo8ihYM6YI4/JZrA431KvoW3YLHdYTP3E/37k6H9oZsnHE8s+0VMWBwtbdLjMYMJ9
6zP0flUza8q/zJVNMNcmv+9qhchPT3E2a3gwHw5g+F8wODaZm8Q+Ff3V6wflzVpYvZPspoVuH7+u
iHQpU04XWrAvEIeVoP0lWy6Q2Gkd0xJYxZT9jRjA4Ra2Ar9q3lTi0XuqWLd0MHaYLjeMplDuJdOr
trZUS4e/y1CJoeoJRqnb0HzaiPIxqrBoM03Zl3w4xk3CTCs14plqDQSkHr+PtM3EhVVkXYkJgFw/
4JwuirhDZn0vB0j4s0lnU3ufMHdX+QmKCP5zTotzkHXFunsQ9+raqMR0M/gW46BU/D8HfotRQNi6
fh3VgJdQp4J3rxyiCYrVC5czpluJdMCPoYVexNuBGWr775/qI80FGqrUcF5f8cROJI6DweXpNka2
ezqH5ImVCt3VnwEYEYJ6Tqhx16Sd/+THlFlSxRS1qWTVKTJduyTVSwH8dUkMhvp0nqSkITd4A+wa
9XKL73zW14njbaCy3Kk15HHJ1Mpp76TL5hS2BFNnoEmqZVb+MEc7FpBYjbTehFjkxfIRsexTMOwT
S+zNySx4wH+hma9jaBcWnydbvCvzUDmK7DFX4M1JAYaPqGN+wTpFiyBynqRP+4tG9yW+jRhWeBGX
rlqCdVY63MDoa0Kqb6HFUiZuEP73c/+hCYDxh7RxbrXGqoPrXB92qDIc0fIJBYOdtXMhl+CbSZWr
m1CntpYvcycEPB0kPcxGhSnNZy8/wdJ/P633P6CM93PO/D9hhdvrPY9ebrcKBV4N/Lce+Mui9OAa
C8jA4O5n5LQy6SN7tcxtXDGDwIdOiWDb39yXco0ttSW3ssI4nFP7K6Qdbnf7ERAy5YuKA2Mlhz2r
/KM1PKwhdkQJDm0Pjg5kWuqpKSCGgqvwRiSpQLrF//5YVcYnQWM763MiCTzcPHbkGnkOoZIPKbZP
ZlVRcFRvy9Ta6N6o9y+MihBV2tf/ANQ/F8JNOJ30WsULwuExblwsglTNmW0KQuOiLwdJiIY0uj6+
ZLbSD88NSslJhz0lXCiaJdQXDDEOg/7qsmJW4FwnCQ2VMo2r+rFBHrT+KocuJR6S/RtvfC6V5oBY
uaeMTjXqnTfGny5njboWEXfJvsEjgAE+j3A//77NxVW3heDdYX9UySD9T2//uogPOrnkpud/hfqJ
73lijSQok0iM3VyQ+gUQYpEGEExruk9pcuaZZXt2iGXMBR8fo8r8w/NWCQFnzrqxcphAZ9Xg6C8S
wrBKv+iLUmOCWxD/GEknVFakiCFPfKGzU93sfNR/aU9hESCI51w1YFwGUcH/2FBxdkuRWZ0DUgc9
pGyBRIzKKn4DTWIxMgTtod0e4rW4t0Tq2Z9MKdQxYy1zBoIXDiN1VEgxF7cErc2QBcGPrZV2qRYm
8b15nlYEVfjIFJ8lvmdwbRvr/Hu5l8i1lrNf1L3p0byeT1to52CBxhTLIYmrUgKWqBHHnrfsEzIw
EVdeZDUFoQ2W8cZj9we6vB7fGCK3I9c5nYd4fLI8oxtDdrBTdb1V/rjLqNfsjhdltEB2Y/v87Hab
stK68jKg3TB27uiOKzWQcuOe7ur0061IDIsc1RTZVXwt8xWw6UvggTmdshmQpVxJULZosI6nvWXo
Vf1Hdpz+ZuSgkYWdqooxNxbMCUaRj4MwFrOsb20l50bTChFQPEXQqBELFs+7fWVQAigKx1uw3xC2
Mdu9aLu5pmeJL03WZfE23fWebJbHWN41msor6bgqrwBDirFI0gbtjsXxW/Bs3rEWT4UdOeh8c97K
eH1IRPKl9I8aBsDOGFg4yvufp3Kig90L16xVsOtA+0KY3l1/1/PuMK6qcuP/WLUcL5+ps85Zs1FI
MZZbMVSM3wlsd2knL8bZjsXUbGrVFkUpk5Rv2j0yNIrHroLNz88wksiDRtUkqoVf3QcTTFNQd8i9
x0D0zzQbvuFAkhNqkpfUAvJ99MBTc6c1/10KB6B0wJJI+qyMh98Z2wDi/rQX78rSWFG0xh+c4nST
eW9PdiiwvOkOTA0awHMHlSOQj+FAXdzwaI8BVNHCm8pguvCsGBMjY8bRQYIezePUgT/UsEhDRSnm
isXXb2ouJdn7KWWyNjXLn5hefoEe17v9dmBX93Cgi+iBKxnxVY577TA+duCgBiC1CoQ+f+NTpONF
ieHqFZUUaHFYjdvztFMVH0mp0RtZOqfvx9DPFBSHPFu/UDB7NSF3ZzOnfUgftD/EP4uAuSvHbZfp
UXMejMiOTI9OPwGXW53yiOYhlAUmlhB0aGAy4kH175jaxGEW6MHKUYUUo3gOHmtUexwX4Lv2eQQ8
JPUEPUeAka933K0dl+oSpv3uTWlcGHxaeDMcSk9cWbrJle3+G3cw6QbEUyMoGfY+THwi5+O6/Opz
X0BvbJGGqvRRh5j02rcSnkXMb8288m0GD1GZmP2y4Mx0yuenYTOse3SskoiETPoVXeqytCcmVtCK
lH71SfVcM1tq9Ah2EPnfo8oMnMYbs4/8/tCKPFEdBgtB0A2hOfogYpuOJ4oo4A9uzLrQfdju1nET
MFjsnvq/i3r8UE6fxcOMjQ0rlXyung5C2jOet9aupDLOb2JFOm4qw8C0vLUIuA6IfTdJzGsA5acv
xmuU6HQImbO7sTJOwT8/XErQnMIzV2BOWJo+/GTAa9/aFJsAgCRHc/la1xfh1ry0z0Hfv77MpRgL
CaNZi+BpfDqCyB6XogZKwkiFmHIHlvrwhJd8Q66n4Ox7+aqcxTNMV3EKRjzVPWVDOWm+dVy7hYwV
qNApXtaZ5Ipv6LssNHb4G24c/WDzws3Z2h8CQWsS4M6hgUNO/NghuiqUslfFzqphjHSWRG2TYiOk
PIbsbYcZqcvLysQBXNTz0ntEN2ybNpPyf6M86N5/m6VxxknaTFVTvD1SewjS7Ma7t2s270X6Ouli
/Ca1ciVssgKHvbTzExI5ywzsmsTFkzFoxrABgeJ22LPJgqfLrl7gac8lX32A6GcCNADK+fn5AyK+
OSR9jAv4untm9vZoUoPKwzARt7syFcIfCwuTz3xwV55i/W65H72bZKcnxUDPKpeNa2jtXZKbOnJT
jUmVTJ9hoDwhnbeONOerHVhY2e+pAeGhW69aWCAOnauMaZW7wD7gxjwE/QhCX0+l2M+0vJ5LdDG6
wiKciMm3+WdKFnr680XY7Jc1dltib3RTOsDgdsmcy83zVWcUphUF4t9d5cfH0F2p6Kz3JxMpfZK3
bz/HOMUrlYWLIGk9uR5lbDaYii2skBCZOlxId45qP2U3BDgx1X8XjopGfhwizhmIFGsAGOSqZm4S
5oBgDKxFH3Ddc7cK6CJZ9+yYuD0eeNRC/Ngc6tdznpJdOqmBnoVoJH5uJtfO5S2ctAElBvaSr9vW
T/pqxCEmbeF2r1uYblwRtzJ4Xzx9dAgbCHdREsjQ/7m4djrCQ/m+7JNhbWqsius0Isj6BgAPOfF2
hip/DolF/wJCOEUUqRjoo8e2ZJ566rVFCqw4wTYm6B6juqHLq1YBfoayoXGdH6xCK5PSAqnLvf3a
VmshO2EOoC8xdtjMb57TvOYpSe/y65EmsqeFz0f+Oalo7/3b5YUrqXeFIAnPcHCbZ5QUp4EVy2RK
yhHlGFPENt2IJLWdS350mecDyQBWvf5EEbio7+zQBAxPs1kks0AzKZVoDgqKJl6ewx748xbB0fbj
qqlrSPqvuAUfssy/Xg5MrFJggCjv8HhlwU1cBQr3/iJNtVuKH3p1tkuEsoo690nVZVlndqmVcNHC
VlRwGEV5zA3ZYtOThvAwgDnOGJAIZutXNYPovTZct8z0jxqb0fu+O/tw1zxKgggmONSKD+VFPAZg
ImqB+Nn+XcyTW0LvN0BFVwA1MBUfHIJ/IgPh8F9RMjV62an1dO43dhLdZ4UfF1PCHyIiyEsdtv/r
EdCsSo+rZKgjE8+/rDd7WBgn7W1zmA+z0CM/TbUqarj/OBrAc9eU8uSqhjLFm3c9WxO1rK9AePgd
cMz9a24Ca1OCwearGfQ8CvjCyzuR3pY+Ih9c0tD3S2udKLBCREbBdJ0NlaTEeeOdWdKBtfYT7G81
QsTPfKR6GHysHMcQbhE5FireDNT7x54vPoGUXqsARwhB4hbNs1+CPxeRFiL2GZY1234qPH6bPFiS
I4NCmnZFoF9KQ58erCijtZ9QXgunNncqo/UcgtHop5LtyES5Qfbwl/aNvz88QnxgDxPzXHx16tet
r/dYWC5jlWbD43TzE3zic47xwYpCk3t+JT+fKXMcIQXk28YvKESLf1IwU7mH5xtSlYaRXmSujYMU
FIsjudhK6z1WohaY8M3e1R+gEtxOUWIjYuVkTSuek/75blqOLs0cW+EcYMQBwx0lfGGOV3llBoLX
6fUNVuDUVe8Fc3VOgJTifYN3rXcvTPyqYAbjEwsukquNzN3MeHlqJQvLuLpV53ZtRDNT/ABWsSz3
kPQMO/gW5qLTMIejAjvdToM1D3xGEPqs+hoiLfH/JehL7xOYkzkHx+BphvS4UqeTFb2N3fi5huSU
SNR7fvlsfc4UaEDGdbe6sOhLdlJG7A8TOjNLPCzewNY4c5VhiUIHhMW+49S/wxJt2YqAKI5UgzU4
jmVv+OiltGpXSAkzRSIshmZEOMLHNq4W8Ju1+5ulZaiM95iyrjNC9J8KgQDBX5AQDDz7MZbEpAoW
Ypz/pI/QZkLB4f0l+2+BdPasbS81QH4VBegj1eC0/+QyxDoaT34+4gAibBc5lFSVKC+EGXhdIvy4
4HeDxrBV93T20p5eI6S9+9JZcYCR+vnFs06IRRx3Ya1LIB8KBLBAm5AHAeo67Fu+tZdBBWpeVMNG
a3y56dwc/GoEdSwRMA9QlyYENPtgdejNEzicVzSGYjedxKiZ72LhfAV0yOmjrX5CpBiTuqyd55Vt
JWrUgAzUbbKoGwpVxUpX/8gK1WFUKm24CX06V52smRAl9WoRACmMJGwdVsCoBaGevAaTrJoiorkv
ZcItIZbK4KtBJSlw4PqUMICuQUCIMNwAZzs8ML0vsDMS/FnjHraOl7VRIC6CInZwnSIKKvgDvPXc
KtjQurautwwg199tTujW+goOkqJUOpJYYM8iEu1VeyqqIXns9AF8PH+vivb5qmleizR9p2BkYnk6
ag0I28kzUbDXGZIRqLYBYYsFmQOpDr9SLI8CooKzZwf3lHCGn5twT+J2pL9GSsstTkb0bacp7DH1
7ojCdsUd45w3krJbPDIkZ/pUHst8eeqW5e7aROm9Jn7c+5PHpFCu8zMtroVSGXzyUQar7GttpJIR
fN5y0pet6Pv4gYJB2iPUZaCoDpkPW2D00mbrnp6ZpwUIwypFyjWv2TQ2ghVrCnEkWmwBA0aIthxw
JhlMFXv+sGU9ySyT2brY4lkO1CiM9ishlw2cCmMgv0rMMrpMaWxTdawgDwPTpJLj/OxcIpQZMwHv
kstIaF+IGfP6sQpHgSvvFQyHhNP8X/cYzUzj7FDepm9TZn0MtLIzeJCU5qzMFuXckWfl9MBTf6eR
1oEBR+R5GM7krBN0yPsmoluOJRWry+lwQCtGd6qt16UNRvYheSwDmzCaO3TPFBtlwTqRXiI2aYJb
SYyD7uJwPFSRRuAmyjT7nasw/EuKq3K3j3SCY4r4bGmsUBrTG+64dUGZy+BoCGJRoSsjmG72Blny
UbTFTcQVqatchahRIBs3Lmw0n0T2SWPE0ZgsIqOpVhYG4Qz5hodYLgy0GHUXHfPBp8sO0WpdOPVk
sJXzQw17v+V13/Rt+qEDRmJnMUeAQQ4ARxUZofq83z0LkX5uOiGoHQDM+CU2HmWiTY5lPvZA8Hgu
qFlwVrOj476fqhe01kXIA4H2NoAs4RFMZzOXnPyr6AV9ixqPjdPRe+dtPoUdTPmRtPdjzmc26Yp8
vtTjMYZEuIEha/ulYoilUFiJRMezcZP3rguLAs9i7K6us9NOVbDwsCPAEZknuH3ZS5d2590BZTbh
nY9n7OKnvFgutIKq33UNMzPhLVSqyYzGwq2fVBg4GMbrAF0NFjrJvB9zLB40uM1k12AEyIgctRz8
4TzWp8bgbT4FS21uT209ouC/8zIV+ApMzCmwML3ALOcn8+ahE7n2kw83oNEYXY0RXdRS+PqJLZlq
xXNfVpcRsWYSN+6saIGQUos1wq2pvF3XPPwqL18T/r1PiLcYMcvUlyryy50Dfote4w/XMbCikM42
Y9NvfidjHFcAjj7BKWiu160Gu2RKYx7SVbKJGhLJ4fbzii+b/urAwhU70cK0AxMahBmUUmq5Ux7y
HXozYk/kkxlc5PW8DszdiLTlPdpUDw3P6b6qNxw2TPStdcbO8d2+nXGKHPwVyexvEEl3MpV0csnc
tRVbMQ3bZp55S0/nhFUuHtE1dWH2HitJ2dV6EBt+UnNK22ULI8Q6OqeM3+qL6PZNY6eRJ1oZ2NCH
uXHP6/szRG7NQ7ADuFWriDfvCFAhZ5toZRCLLjmXgZcSR5t9tyb4/3muvaQ2vNSIDJ2C1PxYW3Xy
UbmkaWEpVAl5aqOEyLRI970NlXBZGFQ0m0/1+29+E3l2j/z4f9QfHqkO+wpBrCK2XiYFQslLtA3v
tH9voRB+iRvbzsj12adA7X9v8/9ZytTCFw0ha+IUi4kAqI1eSMoJ9w8OjY5AsUxOCiRxN40SBi6J
/605lRJXwYKaihwiepFdz7f5IJcpkBOQP+NbsEOalp8IlQo99sHUBEnLJiaxI6pLhEzc7W4WliPB
IOzCPjUVEvvDetg6ZxvNhMrHCAIVVNO4P4PGWytmxLNoMxvJ1IBA2nLFP8ituSXsvVp0fbN6o7F/
cVlsR/dzdJUwtjtj3wk7Xd1JyBQyjJPrJUx8RpAiGruRYBuG+a8HXiRV0bahnRDwhIKuxb07BxPQ
K0dV7tvnUC989LIafnnaIDof4hGl6rtFE1vdBmsYTWEiTxZcH2pfIiSmgWyFPNBczXisZaPaa9GF
1BjYyWOZbnQA7yX8eKg92W7zmVMFJgs5+IE0y/p5siHWeJv5qZC8v0qoLH4viGnezRzSp7vz47Ip
gElMRcL3v29sAZ4nLCH+poh74YlXl5bkGEbbaVaeFxwB6Czskp3brFg5Eoivnp/fVrvLskW/6Tn6
LGy/TkydFo51Nbo5RU9CjwVVUMnCA3nuDqGvyGoGrQeCWag9FymLku4fnkTURRffjeervpwmJtpw
aH0HnbQpyTglOOJKBY1ZEoM5ikS0jbW5xuc+nPsd9W9N5PHAL7jcsZkR5/RJ11YlnGzUuOzNpyA2
CcTxaPb37MnVh9ydqzMV6cOxj3Lgt3AhndzmSX/rxG9SY2YI5GNbaJdqFFF9kIWpe1nS5yYw2Bmj
St945bDoidTrKbtpkCZij+RxbWDygEZkHyGQ+RufTOmquayOlhsiEuSeg8mrpgbwHUjTTPGrKwUj
Q31tRYQQVM75+ap/cI7s1yYkNzPwjzVRL96Wb+pf/Oo6nw3ksLPHx5enEEzPFCGHSxY1slyVsBaR
UiJjPUtcHOJIITJTkB6JO8k0jX77q0HFHdloTqIPGzkYwuEG0IekM1oAgUMv35QdoGsKgfJmQjUw
RlkuMZMKePwBR5DCjQRl8tgVFLb6c2ZX3+TmCAhu6AF8BWC5Us6EqTaKv/YGGPozF7HVwhnkMHHN
cJPX0vPUsvz/O3JyFJ4ddjSaCwfxbK5dgC88xTX0+w/OCYh6eCmWZQRHxuFzXMnpVioYzaBemeDy
Yv2AgLWVyLYVkuIfq7TmiveqgOLJv8VCTLG105LUJltv2wvVx1nVuEHZFn4fvP/jSxP37BLDlE7y
iVuIU3NA4CluZU1lSIqe8jQbNEHLolub1uQzdzltEgM579QodA9JkAONSTg7T4sWfXo1Sq3Th5WU
zAgSxm7ohhcJtWKvyEs8nlRCKU8N7zp820U6g1RICzd1QFmi7N/C+eEcd/HBO48nuo+93D77ypiM
R6CxxVB6oE/NjEHf6do7s8YIV2HZIEsB+JDZYTBokqY1eoqphbiG4RYfy+G2AsRaByHij9REANuv
x63ZMvSmBmyyBElyoaAFf0zapvCQivKUhi9bjmkTa8xgsIyZeMz0xE+5g1Sx/Yq7rqf0zX2KS6Yk
TNVJXfyUpjaxpZYCqpLKLIbNgNQzmO0QN5MwKfJRWZVh1Ua9ptL+wRZWyXJd+F83lv7PGgJd8haI
kAkAcTUZopxtiS/+h3s4no/imfzlt76DXFyeNPJgX9S2A4Q3zn2+eCATr4izJ0/ta1Yiq3BSl+zi
tpYwUpT3BzQ9nklxHhB02LVH/QLXXwTIYGRFnFB6Jiryw6Ax+gBg8n0nr8hUVr+2wS4qJNlhIBGN
LmWPeb4NT/aJ8smd0Uru9xf3VOw3VrZS9rLW2x8vMzQ/aBsmsxVqsab+Xww+4t+U9diccm6hAcyD
2qeNBtcTyZLIfR12B5+evqtJ15Pxw92OB6IdZarQLx38ip7Yfp/py5hD4M5nMYEjjG7Us8AlpbkK
ovxLQRD6m0bzXqrs85rj4K3GTzQDDeHOZkKshUofqu1l+ALAKhI4n/zuI/R8HLlZ9GTLPPC0vYeK
0rBl0mJ2ZSz5cgYvMIvAz2q9zvNlGl6QwCsK8Dxlt0otPkDbNwM5kWnWXqqn41jWvepaMp1a0OQZ
RjtDcoz3+OAQ9hG2NWl+9G0SaVBipY6hAGAh5xRGffW0VthBM6VSkzsq5BzpaDrcH4lElTqKZ5rS
ygZNDbXiLPM67XyO8www4md5Ct+xBPrz8VJl4U87c9AOc3jCTREHyFiBwwH28lzu1SvnYcAi62Mo
0m+EBGhazHgSnZ5wl7u6AJD4UqP3kAHbRfmGHEAQK12TEwhK6No6cWcLcyv8WuN4Qs27hgzqiYat
IaDUGPlWRuufL8wxeQvuWhLOhuQZaVQaJkK8vXY2J2VdA41W9vEFLlQqZqT8k8AKpBzvBcqU8ySO
8yFqOeBCtevtHSwTRuvmhhJirWEDoQIwuwZxG60WHkSarhEtEAg1GfbcAxZkDGR8tlgeh8YL+APH
p0H4CWtsaAsUlAz8QJe0zXfQoyp6YNjTICO/JVabGrbfLxxykBhgnYQris2sz510Y1qgCohL+JQ3
gsS7d5MboWBw7Q42LHrdtA6E5mBg3siAJ7SMc37jHkSnGanL8/KNu38gczfQ7V09bc1LWRRH9FrP
b6cqmhHOcxnH2U5tN5NjjHEnxtw5jw9zbQMfUONZ4EPE+fGA30+yd0pcyTmE4BZhBLwLr6fLGO46
akRUKgSEhDE9f5KNWkSmcHoK4URdUA+EVx3F8KEDq5z2q5wW5HGfjhKnyTuxdld0YYf3izSz5/GI
mJxPEZomA/pwvTxFMGNdq1uvRPrUOsUN9r31z1pwxkLwkM7xrzO8Aa1Llt1JRoNnX8OyR6mmeiHl
RaGs5xEO/B3WoPnxOBN/LAu+isXlFOnqOChkloQcm+mgeAAEm3/v7zxIs5eb9v5WNmmGS8yN1Heu
3F4g8c/qSrGkmp1z7WijUhgySXCyZWfOHq+urozhW0uYqEWyjNI7VThS+p+SJiJwALmXlPZ0gbnI
kJPrKLQnqG1MsJ9hwHM5jheYM4wa3QDmdjb7m4SjvvJIMOXf7UpB+SPjHHWAjBwyvZgGSxA7sRJ2
ouBNmTiaYsbecW68LqN5ZXD9aY5hqcdbGKANUs4djlVo6cD7jri9g8a/of8LaoaGd/8dd7U7GjBT
VugSv5a6d2YaTv3K0CE7AsYiSaIB6nGHu7u30Cyx6FL35jzDr4x5P/M3/IYW1yWSZ4LejPAS5jnX
tvDf0oqHpdZDSkIky8AQJqb6mwkGSo2S2XqueRSWLaMP6orrgDDQkT+W6/Tq3sW/q+gZlQuuctoP
91yeCN3GTRFrskvPaFv526m7S+k98dql7zHXAvVAO6eIdgYVTafeHLPOyqJ2DokqSbMGqo5jB6mf
vA8mxFz70YhkE+1/y/8oTEFTpsdG0G5v3qIlx2gXn6RzpSRyNOmbVSYCAteGqXXIX2jQArLTUPkP
uaK9BUbklDrCNswLD2Mr0c5zieTZBs9EOQshahART9dP5GjkpujwATvT59xBqhmJJK6CXLQE78Gz
KcU0WfrWet0wSJGE1m+JOG+fq2O5721U6O6VgXT/6oQeisA3tvwZFMfmy+eUSUuSLop29LqwUCe+
chysWU+KuLBwTutEx2uL/kuTxjcI2qymSWuyMQfcwETHiv4H/XDNTMIgoGX74x/nbHk8aKbtqQQc
PP60Cf7cAuS4fD1c2Bp6Y7IfhcPW4x74DdgXdC+Booydtk+5Z7oPsUGtHh44dm2P7mSh4KwESfT+
AirDaojEDXHdCiv3hv9ZwrOM146bmY3T7H5LLsGOAgvUzkdhlzhXMA6q+iqQ60ZRaLwYK3ycN3Pi
crnzd3yqGATVfOog3Uv6l9BzEBFTwhZOeUxyQwiWOOEXqYpe/X4xthVvNANYI+UjzZdIsOb1FQmV
W1jlUXG6mmg5AeVzRBMU0nxkcKFe/KHqCUicLEW7bWHzc4asHe9eryiKy91bTk5x55m2aXk9MrU8
OztD8vbvEStf/6YTSA+oxmy+2T1DvAwufaOzLMnm+f0nXepX3q26Ecal374c8umyu9WTcde+10Is
HFUzMWVlDE0wdiqkbv3+OA+KMvJCRMlrHHns7Ka5TYlDvjs/9zawCssbSfJq/zgHNYGP6r9vGbxD
iV+oWOX2O1/T39brk5FGxzyrczKxC3+zXA8OSzPIk5y7BZk0R/N/a4M2uaM2p6CpGepVsushN8lM
9ZG4dmZ4nZymhTDITR+cMHUnubCneVxFxNIwjoWksfQnYBdqlHBNOqYkt883IKrdQI9Ww7/5LICH
uGmH4xgT4MJJfxK73GBy31ptty8V6YKQ7MypqdC2PsZttHN6PySF2URsM8h/6658A1j0SLOGbU71
xu9m5Ep3dENCtKMbRZr+M6oNzPIT6oT3slQPH9hikzpPl2P0dJPIWQ0kTTAI3DJRihWd4d9uwFZJ
U6RK5aqUfJxkFbI+ZSb1f7wI9mYT2Ah1PWHruvNz7oOTZfMpcnijl8S+R7Luh7ZyF+lvBhYzcAJt
hJnYLBEZPKzWzbX8/stUCPb9rnBzSshf6ByXb8HoymHJgEZOSnqAzguNhpWFqk5x1Hse3z7d4oj5
9mL5XWQ7QjnGpKZjQ+aMU4GosCwmV648btS5AXM9N92qvml7b4QiziGDN4CyyBUV/B2uQi2G6q8m
oKcmhFNvGvYqkjRIFsVjGluq3P2pLDoJQfgilVMHPlExOL+2xisbsVnyzJ3aYvwW0f+At7lO5IEX
dQQcCqTnKp9HFhrTl0QpG9qTl5pCk66+QkBpqVUKwPnDGD/jJ0sc+q/sam74hOjQP0Xjt0IjzqGN
p4wakUYZg3PjghOZTo6HyLdQUtx+ylUAHNYSA3qEgDa9eBQj0qPkNNiaO/4RUVcZItQRv4SWVVDJ
37AIMTMH1lacx4k9FZsgTBSEehUnvhzYwaqN1fX8iGkOXdVnT1NzR5bquLUGmME454APNZNMtwGn
a1WkiAhl44mGV8lAFPxQ5l/YGZQUXTcRS4TwzOAcD3PxCEshhUq+HkG3Lw8aFCm4KA7AlBrirO4D
PJsAZYdQuFp4QREuPKxm1tqatlta/91WEwmYjE7Wm369FzbSx4cXpAZRe1niKXnpEfU20j6BDXrW
Pg1TKWCV2Zzao61sJIqYZZVOQ5IXjKg08kDImZ2LjH9rs9mk+wCQ+nE+WRRxXCevlb4eVLs2m3LL
B6UALGXPWF3VdQHKqV+Fw5Qw5G1io7X7Mt3IafHsUW/KjFJoWVP0YTSIoFv0v0MZF12EViJv3fqP
XNHyzMPYD0ZomTajevgnm807S3qMJoy3XIvfqC5e2c1J45Z6uP4wZSvUtbDyaECxERw0RRMR/uE8
eYIda/3gLLeAxIxLLLVNmWgcCU6DFl+GNIHqSf5ezODhNQIsbscMyBRHRU+6ro8aEz+8CFfuSnM1
nyDboKL5zDkfxC5cPbiFLpLm3LGpPlVgLTGc26QKoMvqAVe4/8/pH/aDrgn9IELDpMg6VMt4bEqG
2y94ad/MFEKuYGncIit5FJl+3qzzXw5W9n8505Mr6m16xXp9JFuy86RC9eLau9MLzU2DcId5mwpW
5ZoYL+7TLM61s9WLrS0NuQ83qe3posIaU8Rrm2jeeoYxvV0DD5EAAOMzsTwAh4VHgaUFItLzlAqT
M4vNLDKH9Be+x6qMhuuPemqGyQX1FsrafqUlYSsg5Qrqimr4tMyA0uQUslO/Mdy/MW2JeVV79/5/
qVY8LpSOVutUb/0ZDqYdW9AJybQ0nb2IcOMLNMcEWPc0bybBa3ktqRwba9xu1kWwruscP4jUY1KJ
htJyiggSJflxEDJO+FJtxAYrIm9t7aDLVXrko6mzl2S+u0vCgzaE1ZD5cycJKATC9csdhc3dekBE
tSfGUR9CR1nBBNl/iyXswJFb68vPywbH+oa+B/y7fV4X86ktAXDTATS2aFucb56btrRLVeEKIE4N
zfD4PihKW+nzBAWO5e56oUhes6Bb0aTFMwFPq+l1cJwj567TfhwJ9Kii4l0O4eO2LpSlRivd2NPl
NhOvkzeDHKADnrAx5NPiHiYHmu9ObTeZvd+MW/8GnvuglBV+yPyZ9fl1+d6doJxb0LMbTHhwOLP6
fefk1z1NZJssJrgl2ahc6YPMPjbEXLDCbwU/6EzUZcsygxaHQ1zX4l3BSawq7jcVpCjd8w2jwuMa
xnl1aqBo8o6QqmL5rrKN4mGpdxsyx0fUXHExxfcaknh4hVNdk9WkVxCUKOJCto0nora04uj02QNz
SpAQnd3Sd/GHRl1D+BYJrR7niGozyLswq5EoZYHFMgHQOGHur9kzHcMKG96ixB6nhs/KvQky1+PX
DsD0dh+ay4ZzCtZwSftgSurQgeoXZFmHGgckJbdXgHZMRF3/LhTjquqokx9pwimcb5lj29RtRBst
O+Nu+k9QCg76kavEovCtJYUg/PNa5WYuwtBrPyIQVZPOPT02EzGClRfXoFpD0EWPzZuYJaJokq2u
CLp2Nns9XuBQPfZM4hrr8u6LrCSgIo8oX7q3cqbJxjOXgtoZYs4MrPuNtBMYdApt7GmfmCex/0Bq
QwleRzotLwOATrIEBx8WkcM6FLf+RYKPGR1O1+YxHLoSgaq6hxXOSghufNqbvybblI6ZTb0KDvhf
K/vMirqZ4zxzWULmK/wBhcZ4oqehp2XDjJvA3PZy0L3EnixHl+m8uPkFYAAsHUTxUUuja5SCBAcl
+HoB/0YZkck7+dVe4md1yljgO/Q+8wjV6AZDBkwl849TKPFSR0AG5+DndkOhZI/EB5AiNAY6THhX
z7slMc96iGnU9yyfglpsG0zItM7YE0FeaW3/6IgPlW46GiKM7lRzGeSR814QaAYMLaODojyDIJGQ
W/SrmddoUlxCj0C4BISkL798AODrJIU/0e6p2O86xP5Jaex82dTe1OA2Gjp/W+XazyeSSntOB3YO
dAG6xjMAVKLkVfgKmfExsJKbgS2RalQXJMKGJd2sVQBGWczyNpzLCeOwtxTkHscCurMd6gsxbuqz
3/5OYmW51wLUN4qPGVj7NJzr0D2uUp79yVe+LByIehveBk35n40WbikgesT2hprSJ55UhLCkfVLD
PJ3RPij4ZBALTV33xdb29Wa5zz5InFainkc/izUjEG4ktMgO0dYSS3wkJNuogby9TJTIhGPVN3qH
IjyUG69iOTR/BdUSGzyMcNdm7cx6p1S7tNAtWngCTo94nKMAOxxXqdRj8RlHtCcdhmv3CvGHndg0
7VD2CClA89ClTZpN76RSwzrGTYY9STC9kOIC6k5SnYhbSLrOf6N7aYDmFUYD8+7UdiC28LONkZQ3
dUtqGq/09rg4JIbXuS64EfyUp2wSVoaXAsP1QKyox3BBV9aCMxWl6TKFx66BHwiYD0bkVh+OTWYb
5VyNgtm8tr9H41cev2tudNoFIaZEOf119DFDtk7LDlvbi2eW4uhdag6FPWQoo+levry53v2SxFqH
ZlMS51dUcb6ToWxQ5T8ealgWutYhxuwvK9Ye9QEoGMKKLNRnVNNBxUAmvHtfeWk02qOokhNvBQpQ
AP1tpDCzZML9H6OU/MCQyjt9WgKj/OWw0XCi3DHvyeZnuUhEHfAzBFRy9EF8+RgmX6AHiyleQNEj
/XjxEAHNtCFiIWrJRTTIcw8yiXQB3Bq2vFf75rAqMq9n2Hs8nl+yDd/9W8oXpYNxSGaVNKYTpIbr
GFZKV2XpuN19tlrLUzsKEud6LZO2kua+sGBOpJhib4ykDq8fSY+n9uT+hh6AEzGrgV8YpeLQu3gi
HDe+VPqCU3uDfZbR/nhJnpv03aHg1aTUIJ/uDjUYZCVelgwU4UX4NruR7J4oD2LSWaS7yleMR5eO
YzdlFBbdL547JKNq98ozz9sNdMd7bqgVZo0l/uVmUbckxbo89OIVQJbQDPA4ACILcsaiHaXdpYOI
dA4IccboUeqhxjnkp1B0azUwAvI1UPa1C4ef1DeL5fAZACK/wQ2v+ot0A75Rr3IWwFffcjpyp/jJ
wjXSFtIHJ2OK0lnblcY0hFRjvCe/srBZWdMCw2nw3+6F0plZd2yPxDzpLBlCu2CrxzdVZU7hKpib
0oucxOTtgPGRIHeJpPc0kksHS6CCVkjV1zlrU5HcvdPYt6t08RLimqR9/vMI8eV3oPBoW9HsWn2o
9/EpIt9unXwH3jXhGF/pzPv8ko4+ubOtmNzntXbqP05EFeWWEAT+1Tr5i5p9nGlv6T11Zxcmry/d
CPO0VRdGA9xBDF3DSKoWa3qNu44c18jO3OETBugvaVA0mHECSLoaoLLTzBh/BEjvO9Y0IQIThpzi
LOI4aPpzJrDoxp8xlSOrIPWRPPf7cxdUFdfgeB+5tHlPw0N0rWbyrwQHM0WNxJRiX88hr8SNPDtw
B7JiQTT6gb0FCxBZG4VNy2p7y1CpPEBCHQmkG0m8Ncgjta9ULMrQT+z7+B2xNtJTxoLtfEiJ0afP
2Wiw0/vlEY4TKTzvjRONZeXU1EetFrnQvMLXjfbCvor+l9lyLXbpVxZPPIVKmSlGXCPAH02yF9m/
rVmkRpB+h9giU0xLVH4JZMTWNJvyJmmBX/nvQkc+pxT5PS1wq23er6NnRv5Njvgj06vn4hvnls/M
ZitILJHfv+pcID2pNN0Z7swZEr6LoY7qKnl9sglqKmtX83loe5r6wEeTp5v8DNIUWq5ZvV02wRNU
vsaFr/kjSoGKg31z+l0OQ8lADwP8VvoxkfzmxL2tJ/fMIP2GlkWThFzEyQXvjLe/cWhNxWIzoziB
/+v/xRMfk4KUltVDerNpwnrHMPabQsQoUSDiWkKoYt0t5Hprc5rx+TMhMr+wa/Am5wan1iahU4FI
mBPB0Xxohm7LNL72ybBW/MWAWuUcdsQYVVCTi6Y8z3tWbqHeVeyG/k5QrmawwqaQPvAs2Ic1+MkL
WXHtvXPJrpxIDSdMBKbgL9W1nuTR7VzYRgTG+uLZu/0nze9eSs2saO8Y9kzefaX4wcxjupd+KVqC
FK1ZoAcQyNBRUYgeaInRq65YbFvrSNSaSbIQhcGhJuN2SBTOSxLdUMbeTRgLFCyVMYOjkcnAnvog
HCz6IPYnPN6IU18hykR7l/qfMCfzPjCbvXHEKltUvmystEihmZ9bKqqUegLoC6a1KypHcqrDTfRR
rxnSVsAPuvV/Fo292dcMmRCg28KPXHeHynhOBucWLjqlxslankpM9/i0H5+qROLD4r1A9bM96mGI
Y/P6fNOdUulg/YhYnZcuxGIF3UOtIBoigAAJBwNWvbQ1Byq/4ZsqM99KzgRs4TfH+gLKgBbieWUI
48XZVnjGOj0nd0a+aUmMD3ia6Oh7DGfN4ctrwaNspGzaJCNyJ2+T5GHhqIh+y01vlmw4Z5OxVMdA
jhUaqP8MhkV9ynr6Br04H5Y/DDxuGCOIShczMp/HlRL54UQuPzKkiX0c3Z3J4ED/9O404UXPiQsR
zX2l3MFKBYTJzDajGsUKjrglqCcVSG1sBDdZAAlEUmobRYoz07nuk+wp1aPhWwO1ylu9umHwKyOi
g9VO5wHfyYMdo1RzacBVzj+hYFe0lavu/pnbEyYjUcpO5AXa+/IacCHJ9TLOYrDVxPLt6mOUPwAY
JlgF6S2mOVW03HAi764yTM3Pvuu8XaO/JBflOHQSNJUFhRmjfLXh7JuFRcQ4ydaCW7No8/5ZlO8w
6/Nm3G7RsSJClGR6YYACnkPN1VY/mr+V7Saz8g+EQPdC2YHPr5/PeuwrbEztf5JkV6kv1iK+fG50
dzTpQ6YN9S5vmezgO3iIL2/iLEJTxsIURjjbUT3hKeQjCJ24CqKL9PzJKY004zAOBTWtWoPDGC/4
xiSY+ObZmxT2CiCrAW+1VtDm9QcR/78sOAvCthsC2C0Yl60HhUKU/ZRIbiB3abJb2BP/u/HX0oUI
0ri5a6CMVkf40wxQ5RzaANvypan5peQ2Qjax3Lq1pyJNhezaSJbk5biAREnAT6idfH6xgak9rLIb
qk68EdsSrGUBNdio5880U+lKw1wp1xOYLIJUUVwq6a54j3bNz8Fj5fHA42Y3NGS2XPxPtyYTH696
/dTnm0m5UHYW96oyb4wygOflSACHzsXjtfisijaNk5cg/VpW94RZuT240hNB7dG81Bzax4W9pO7P
UOELOD72olNkWQMahiHaea4hP/kj12hKJ1e3v1dlQ911/yKwDqSo8DgxaWG2X0+ad3T4WMJGLQ/u
yKAxfi7ZT+kIVC6hW83fFlBKL/731Pz6RIgeq3i4osyVDR9Wp0Wjs9fIq/EuxxppCimx4Yy71mMT
u81JSeOpUOfvUB5DB9AmTpBcAhEl8VYaezaiHwVjC9cjlc/RLD1l+L3Dpqu1/BThN4yMCoMv7YcM
pIL6HjtdyxHcwF6VgQyEaJLXNm/VhTV5JSpzlPC2f15CWHJqclEfO1I129GTH73AcZQPD4nls+/t
qQ1/1+9TMaPM0gAJ8ozmhqOWmHyxwTlg3Gdfk1Fv5KeVDIl7voFxmq9RCKuCVWt2KfE+Y9WtKdnn
bEhzkGRCH7yVWF2A/KTopXL0s56rYHgnS+xKlqvxIiyAKfaBedWG3XaEErzU0yyHtr3D5pZHfjqL
YMiZ2zUMzZHgpB7rWuksojboiMwLs3mtKpEBeF7h7BbMnXdC2/5GxNk+vxFtKa1KV4BUeKhDC6lT
ynkg774OWrvh59/9aC8eG8HsqvG5X6UyNn8r5GyNUG7ii+uSbRUA2zDXdjQ/oxh7fVfoz0DT5LFx
mKg068nV4uzqiZZWn9XCn8f5hOvt4sJ211/RFJR/nN2B0brjxt4bhKyJysdRVQAU5tDw3MfVniLk
RUBl6MNFirEH1L+AAkGEhEJxpyk64K4LGTEguW5UmG1o7WOhYwAzGhWIne6yjLsv534z6DlqFPW/
E0z4rwxFKqXFWl3rF9x1gd0tEBVoi9DX/y/vyoSiJ1tfjwdUdaRQX0qsBLGObl6TjGkKuQ7PAtqW
FduFFuE53ePSkmPW44HT3eRCdY0GDcoS/MsClToKrqNIW2UGEKJwflgA/SwnrdlqJMFAH09OrgxQ
m0QaUpVx784EO7NwjtaVHuZUNhE3GYxOQzG4yu9kyVKfMIJqsAelpHgchNMdbnSF9oCc2Qm08kvE
ueLcAXgFaDU7yCMygXGkg9YJSoZJYZxV0lbbxtFhgcLXMdfaZRn64ShxWfXdCYaYGJhQwYeD+opl
Tw/ANckK+f5KZh7hZXQmh5MHcbwQFQW1W/uLI42xRJzcLwHj7zpvAQO9NU8iLDpC+vsfIM0xKVj+
boXHeWICZzz/163z8UmU2zoRK+tpevnKgT0fs2ukqXT5dkdUe8WDQWKX1/9yymaY4rIzguFLQiLb
xp2/7RLRNJU11Ueu+MOPLcGRciurpimxwf6e4sNgN6JLrsoFKSMaOg8HIZel2w2bKCYz7KPc4BtC
RvNUPjcH51+ls7k9OmIPzjY+NQIO15W3Ifplo2K0y5ERMa6IkmPGNOnxwCbIZWr4AyslZ0euqOnV
t8/ReeVkuWjDqexZQms4v+PqO20x+MaA3heoOqSijn+LJqE8cEnuOyFsSYpZg4/u25BTfWIYkCyf
U2PDDiRC1XYfuQtXqOxwFRar8OiZibgNsOLUbjZpxsVdaTx7A5FauDafB2cVG+fpBFOprMl9B3XV
O7Y84hjA/DpWqkf3wyxwGCLqjX5yP/BCrmF237CqU+QHVLCfVYfERinfLNJTEgJQq0mDEN/W6jJP
y9RG2c9QiTfYvc5mDHlfdqAuhFAczvOFMk2qLaF0EfTKwHMRuG+mKy3wh/f3j4YhkSqgpQGIppav
nr1DAfu0yDqAEI2I+JWlAW3f/Xo53F+Nkv7elqFbc2dM9vly8YNQBRE0ljbLkmeI3LVbHzF4p968
+b9tepam4c3JBZRJzqFnZiL8l6j+iPocCaZSp6jgBUQY8Mm5ulmVS7d/DI5Tf/xsncFEZZid0i7u
lrc4xTGbn+vUsLsP9xKhe4enyNGUGtTmoSeYaJRKwwgzOPPCgQTDVYiIm/TDIhtOVwuIS6PeXRe7
hBCx2qm7W60g3W7X6oQXNxiGQ393K3VfQ9E7opqI7Zp9/xAk7iD3sHhF1CD9TPvyJ+BjLRc/15Op
//Jn9QG23WTaY/FqbPDdYbF709jaBp/lVm2PmvxTEOPLnDvSkC0G5qJiiUCpgFBJH52Xs8i+UiYj
+vKERmnO8lNHUZYaUYx9Jt37lw5zJKJg4dsDQ3qtzwWnPdh1S18DXUcsBGWg3SF0CXEnu6PSiKyx
bVpvVc3yXhyXLyhTlvsz4TcnztIfG3o3qQzyrBo3rySjqTx6ArfpTiZUimH6u6k5wLvAiIfOngom
UhIPy4SZdXplxy++qgao8Ezmd2i01ZAPRdTNHMaKTT4HDcCR0uNiJscTUC4emGMmp4pxsZ4jLv2v
q6/hzjBJ7hJy3njxzTuTNPu72nLeNiG3Ex8kX/Z4s+HtsfPFUbRlPiEEJhvlZz58py2o9bUquFmO
8KACdfk1BGWMlptgg9TNG56fAJ1K8FkwSrM2fFMm2Pq+SHfkf0G+jZi0hI515ZBEDR71BvhFZrmz
CG/hDHMNuIfUBDBecSkzq/LaxYq2KzEK/eStIKVIiXLZZW7lG2Y96YhZPTlbuO91srJ8RQrGcz/h
Trw2+VhPh5naoeruGi6NzMtv/2fYYeTyN1fFNxSgFXv43LOETEP3wpuUUkmcWMlzrtUm7wO10ZmG
OnEIWNxj2ovQ+grTYcSSQ52lUioRpOEB0FYwZ5C9euDku48BZgTshL42R5+v0YzkK7ghu0yH5CRv
x/j1u4rKdXPSUR0AwVjw/qKN0ONOM41oRUFb0L33ez0AL9EF9Ir2VeMpJDfe5zno67uldAs/SvSp
qaF2EF85q/+Yp0ZYpGFQkPnkS9yIdw5bBNT10uOFai9AJQiq0mEcVnOR3lLH/OCpxiIRSjsyG7aC
VvX6WPeIeKgm26MDQiADZShx8fMW8W+TmrUYMRKmvyRlAsCGgD2ffR2aVeqn8TwK5MVk6C86ztvq
/i61eg30X9w3nFZADLpUNxSr9VlYHPTUOcXo/D+q772rvsLIPW8O+XwohBXhwMnoxqeMbnKrYMw1
gXVpY09Zc227dmYG2sbju2MwbYjl5aN/tyFiSMIP80U8tdqKP/mdgDJEfLPcXTn9WB/20zK/716K
gxRiazaE07CMCIT69bC2gCQ9f4ljOU6TZAZ25yj5iztPc6tgpirDsMgoYcGlZO7IkSZNe4RT/kra
qLdbx+EPxAsBszGFwdjIT7yoUC7zmmEu6aDNMm+T28Ixo+hybdnG/kxRTWbbny0MIeG1rS8S4Zi/
VkaNt6OZHwm69/hzIHQqU+n0WPEC97Ljbk8wtwKk8riSvCalnwbVfmnX8Zqz5cYRrdNcfgkHBHUH
ryn2pd3slTXMtFvdPbm8+/lrRcVJUpB767ugj6zMDERqWIVc33opoNyVILbsMUimho8i6fLKjEQp
RvBIuYnIdDtA2ULRsAblM/1SK8f96RaECgZZojSEd60ASsZpD5/BexK8ZniIjCIOUDs/feJs/kzR
VI7V4MV7CsjwifWOE3iQXEPQ/8+rqX8RHWUNbxkbUmzaNhi9yo3gH99+OvqJYGIfFAJ8daGHWUJg
1khQEPZXrdCcGjz148nGsG3AN1PiW6tJ9ZcoVZQ+KkbEO3j0JsK8eW3pCSSjMDGm00FN3Nz7jkK+
fL27q6to96CYdAPM7Wno6VwhZxPJzS59OzwQe658BJM1nc5rf8DDJt8MET4oDcwY4r1Yr1qMU0HO
yztwuDhpZovjQAGG9YMaYpJgI8RKY4NwrpzGr1OGkZYC1pcD4YLss+rA3KqyNwBkakd4t/HDyb0M
/VPOgTIvQ8Wtr1+3XVCa9MD0uNGiQK5cFnlSpYIV6C0qGoiBLYZzb/3RjDDbjvu19WnuHPqw5dHJ
Pt02h75jy7valU5nTEAllfbJs96jsFzrQKl+rmSoacfuPatJkhNP+YU0zVArFog/ZRmEY/UHClxo
TKylKyiD6KattF3FTureK/2N3vWORHBmYS354YOTtQ981ftwM8P5Kd9MGi+I1rQbWklvCJGs4mSt
/+Wy5brLbnOq2OHjM1obUajvS6Hgmd2qd7RjMTilF6vU7IBfV7v1QbsDYvWDLuHKt5St2QwzRupo
d2KYsN/ZF+hXcpgVBO6Yr+7ikR17RNqs+Mp3RvK9GTMiNRhMk6fX2cuq79qgKjADNeke1Cgblpv/
KDc9CaBxUHU+pBuo3AktteXpbsiHuMTbCMCsBBOSbU0TSnTpigj6zP1toD/TLs7F92SMXUBSKdA8
83yb4W6JwHa2KO0V2fnWHlNLHzBCi+e3aCHimIU8v0fotBgCdo8KYIweAzY5FLRERsdwA57SnNDS
KZgk6VhUssSLuOixNcEx2LHeWZiPHNegBhRsPaiom0nMEofq5HaswKJmb0KdPQGmqFBQRpsPw3W0
eI/LUiE7uMp+gfFq78ZLhRA2njATuc/37Nl7GNIiEgHPYy/647nFOMFvU+sv2Z1MB1yXtnk431A3
UfRN+nl9IGCsZLn84tgu1e2YYRanbCDGSmohL0CqeGqm1Xcd2A6fhtxPP/xuLCIeZdVZwJFBWAVf
L2jJtDXQpgS3BqGHYqxLBeGeaMpPyLx33rgpLhjkvjZXuW7SDqtD/6v8TrjhK/a2x7Y1spxhEEjr
cD8rYDBOlcctlSt9O20mHFFfXhEWxgMNhFlgoftKocOuycccgIkUzvBGdrvjCgciaD1wqytFe1p4
vIYd/HY3Uv1zrGLl8v/XvUb+DwWrWxuvM87b7b6ejcS8uAzAEkP1VquBuekXgIz6HmbDcx5cBkUH
hzahBEe3xbW75Gf/cQTsrsIS32E44p2DD8Zt69aLzIWAkO583NuCq3GUhJkCdTSOIVhHJyeCs60s
E7+9+PPmC15rfDaE4cIJ3CHw+XN9Vz1o4KeoEYgk5enHn+uSpVgGyE9OOeRDIFtgyWRoRdkD/l0t
LumOD9zH/5hBcI/hr80aTyujU00+2CrW3zp4M8NioTxi+yL5IiGg1xX8ndcwKjyVtF+ZIgf77v3b
9e2SVwXVRk+uHKOxNaTKWFOPMSYm4uu8e3zDFWzyan/B01/toO3OanjIpjvZ0LYiLvnrJa+699H6
M6M5OLRuBFceRNDIVbfLEIXq1RqX6l3lqpuMV9WnhElSleGnhsDVOHZSRU1AsarH9zi/NEVtympQ
v8rEDW3wDwsZK1yLffdS0t3FyCNF3pozNRCSM5KsWUlsUnDZ2npzqMShm+j6KEWXhZ8+uvbAbp9f
riGgT/fyN7I4Tr/uvXQr5qF4Q/4kEmeO9PBkHL4ldN9tv2CKBNWcD4DizgB2gsYAza34WkIO5S8e
tI1w29TCRkLrRq3KKcHJXmS8o22G+JkAxORmUUMYWHOdqf2/F7iJugv8RYIpN6/AYK7bv2/1s57g
sp/tXMxQkVAeb57OKcry3ok7TR/57Wu1K5vmAK3WPmDq+hwceUdIJ062jdYCn0knCkkT9svzagDG
bzoGzqg8Q/d3l1p1sMnc5VV2Ra6Ouwirg2ZrC6BD/3hLxyLWJHYoiiHYRr3PSQV4MMmTUVx39SYf
BbV1PUpTXZ8MnGFeGURMoqNkFmPZBe5rt18WS6d7YdAxgxtL4dfayjUmLxgQB8LUGLCateKoeW7o
fTrajNG0O7zCb5LCOXKzEZaclZH4txz17NodQ5QFz1WKR3yqCR7+nTF7ekKh/tfDnFxM/F9x/zbA
0q1z7ejoCnXXHA9IQRi3Io6X8lAk0aeLJMlVlORIc1w5XWKlRg1hab+QrKF7SyGoKc9CtCEChCnF
e1JTfCqYtbYAQj2fsJRJsL7jXhltbsxd+YDXFmmllMPJwsUIYHu7u9L5Kogf5p057s9ZaK/EBch5
LO0QbV7MKb8zvWMMy3ITAjzozcJyL9doLXLm//6o2tYQC47XLThna09QjS02/TWbQw7pga/ND0SU
g9+1E/IRXEwa4ZH/AF454nriiGr0s7SLKo2Qj5cn55dzyIj1pDYl/WLG7j9w54NZW36W7ys0T0y1
Q0laokQflwfPiCP6IQJSwd5nl7RV4atp0wFa+ky/92woBImQQAv4rGggIQ/mecnMXXPJqpy8kbDY
GwY9/nSllvTJLaf9RS90wrlyW+urvJ2agmczLENsLqN5Xn7kj+8ZF1S4GOHulA6ErJ8jJLV5J1Fu
AtkPWt9BffgnVSyVmtbLaKkK/nnCt+V8ZThbqD5QFykSqHLk/TyoctZDNjhXUmewofj+WihgqZxl
tUZuCgrOb+z+zgTAcC8MtKyqIc3mOh0aScBgXxHxmysATMWBuKEJ/T8OHue6Uoe1yfNEa2GwkWEW
9b7moFrHI1XOJ8uu5V3RFwzAsCK+w/sexI5HK0Qn9mkOly7u6ebawQr1byW9J60/Fyb7k3CDmvgz
XiZoOl3lrs2VXINNdThIpHKEeLYQkOxzACA4IknytJFxSMXpYaT1t8tUlEm0E1K2xLTMvAfzhYs8
jhj8D6HfxW+WUUqN4TPiH37xe00fvSUCBeSLxibBV98cbBQBkSgXFkAB+x5K3gzjTQg8fD8OFTnv
dhmcJepWY82RxaxjnT74L4DotJDsM/ad8npCLeg1hVH0KhIARk5w8GWgjdX6Ds5yVofi1BiBBbTl
PW0CvLYKm2NNU5o2B9p/65Skpv7KFnMwT9SpB7y7mbT1YzEyU31Y5pM9uc9O/+QTBsKQ4N7t+8Ft
94ENuvfLXiRbcIecGcfSuo12me5uUhW2Ry+0jpOAMOFySTrziELAJYA30hZTotwSdD7QQAGAb6xf
SSuTvVM+uyGZvY31uQrq+RFUPAfOF0ClUtbVGxrB1RCsiqoRbDTB8MODT3vApCx5Bs+RQnPvA33h
4AV1hnvvBL/1Jk5wAyrhTC08qkuyTivVIbh6Gyf+zyJ5qOgCrX9jeB1bUwsiESiCbsejxvwd/sfb
wW7CGIuPozNlhrSmHWbMaqx2vRfO7S1goiagJ25nDHjY539iT/pN550g0W4oL5PxcoJ0H5u8KO8r
7shK1B3ISGOAdFWG5OOUrpY+WY50afrLL/SKH3FLO8wTBJnh81Xw8GKsVZdULUT227mfzZSMiidd
t6fgmPxFHnFDSCOXER5XinZ5GBjC1u/sE7txc+38sb+Ps/ImMFS/FLPA5My7E/cLISRps7NZa9Kc
ziqywHQj9Pd79yH4I1Kpn4Qg78axBgtak1ZBsqf8XjqDrDan7U9nNuVjWEo3PunMyNa28jM/RGwA
jqXpCLJkw+1lvJPjzzAwr8qj2if92oYCAIRRQDXAciW+2JCeHAxlgi7tPG6jna/9RE+9AwnBy/vT
9SXPXPNcSAjX9d7nFsgqEr6/L1o2I5lR9KGS3lkBAR/25Z7M/MOib523LPSWaPc1B4O0ydzegXoG
2//VstoBvA10eAjH74FKX2Qbo+oYTU7dUOK37QI68jUvjyetdJZLx3tGb5GEePGdIZeBU7uILHiW
WljMZMlhxQSZqy95r1HrFInPGiZX5vrXzekqaVBA6o9PnEVD/L+VKiX4NskiUkJibc+p6P5C0dQF
Eqe+c66YacYuZZMHVoDeLE6z9dUSzdltt/3UOK+xYNa6xptWsicDIXgB7LU08ps/FRNYYd/ZwaQ+
baUatPYBQKtx2sXIYK++krWg9LaGaoIej9JsV8ayOfdPivahPbp0mvwzGJeZl1DENDf16ockYPdE
/MXG+Sz6JQxPdlOVUfuCzRhXqLjr908Q05QOv09AsRYRDYzDMrpaLKiHC4lgRsPVzdn3KYMqEVAt
/I7oEVMoOC39pFSxRzA3jwjmbAyLPC9Jl7wrLnarNTvLx4k0cxB94M9MJuUUTZUzGYr3QVzXIyr5
PBuytuE8Dyl3p1jnk4fpUaVZuYMwUMI7ITP+53Yu1jZAj3EoOZ+gH1skvgqaXkZSC9HKZ3UI4cnS
Iwc1lzlkPP75xcGAeHdAGyhUPqbisUNq6i5BlXTvM3nRFyTGmkQDL185u53gh00XO+Auk2Scu1BJ
Nfo0NopQ3DovpDVAKIN+AX0wi38KQy3h8fncznJ3+J3sG7rJkVyZinQwyGMEkBF9/Oay4YZ2CROD
z3RM+MZOfbJrNHmQaGEDOcMfxZqpSbMBEOWrDSSP/mKYJnBzT4NbL0S+m7femD7ocgfWsq/+sciz
/geY0EiMkJ4C/svXlRefo5VfUg8wrZBt/unvUqzk1hGZoNFtFnXoe/LnCGqHGR9uj4cC278jW61c
Cj9CVuUus7b5O8zyrfLlCgFw+fyqiH/JmG86qBJU6s35Kou460Fd155lmePuOsmPy4Mi44g3XXr2
IaUGjsHbBI+sYACJcFXPcAkasPXwjhAZFGzDSn4r/tNh78PFMNEyrP0cy+77tTA+CAvyU3eMhok8
GLJJgEbWF7ky9k0CoSuRPE4IrYUmY3De2lbOPbC8w1/fNOR29aJMDZVxR7RUjlh+hDjk00T7RLyf
uKxP60kya/EGNJ9QN61THl8GDNHMAc70xGd+Cz0RUCfWboZ7wBztZ8q/Nu3j4nja7o7KRVPft7CS
yrnFirgUTaTvoHNERu5BuS6CVK6kWAcDZ7+7GuWiDpb6i6v40jesDKb6jXxjLCKPFE4KLoeGloMA
TpxJZayzh1T6DBsSArICJXQBC3zHU0EycEPovkI95BeRFYP7rOJu8HGq70ms4Ej+gGg+cGbV10/b
1a7MbuDSjad94j3tSmLKfvi9c7p0tc+xD+y35YrMkFptVPgaqsaFWXZ/y7G53EmOGv9NjBFGTha1
z20ARHRe4goCHhs+EdfSKLRkZT/CELaehP4k5GiAq3NzbC73AXV+fDzu6cAmgd50aC5s5OvaOknH
KYT4Ybmlz2VidOZidzsy3vD1X5OIObm8rGMdS21Q4/cVJ7Tmra0QEPkdo/X+UXuhYzZ5WsBnTEHb
blxzaE/R+c28XrjNB/OlQ9Tv/19WvHldGa7pS9UV5CJPlo1TWs0y/WRSu6qV5fvd+NyvUoDz3oJN
YphgnqnvswlCNXZzvhSvDYUhYj6SQnoX/Ri60Y+qkiuvQOmHPN1odAM1JrKCMgWmo5uZ8VR5+Nb6
lpbqkZXIngWAjScsr6Ehws5oAfFUBrCAKbqGhWL8Ok6+xTOi7AqOHplWS5I/nRQHTnGtKqv9Iwys
k4schanm+3boFzllbvQgx5cd8bGgjTW6ygrBZaU90EcVyUt+l8DUMwrtZJ9fXcZT9b2JEDFvAaVE
TqK413d2iCPl0fPwWjZpBWSeDXfymgr2xfY6jPdVz2aWhSF7Knr5+b4+BzZUSoeI73Jx3NXK3yHF
OXGNTvspNBOr3A+elB7wrntF2milOXlN7L+U1D7q607FwXIUsXDVOM3T9SRfo1ZpG28Xk2qwodOC
T6Xr/NCb2zxh7mM751eUTEuiUpnGbl/2hjESLTS91fprz6YoIEZt0MtSx4PS4yBxapHUpITXum+6
h2zVuBXFA/IPF0zBeVi0/McOsaUslAaa8+aWGT9wUP+gk53fn1ENmXxtRTkFZQHnRIRdbsPpBonT
oqiNeuo2s2QsxRuCuiOMKbKr1n8bOoL9cL1jDhMUb+6245A5egsC8mOc7OORQRFijy1k0IltQCnd
kjXjwq0UMOB2JRauojyF5FyBzxmSx5/NHIveAxIKzJJQM5/VWoOREA+wfi9x/rQAM0c1PvxR1laj
lVeNEIt518DTVcQN4b0Xo8XJOTyY8Th5XgBSIE0zqEmdvapMEr9+hIPACmGv5FUiJ2WNEo9YiO1N
VKU4XO8t1XX4a1hITbqZnpZ1fzfHrIn6by2ss5nrAhelUsRHanFm0PC0LZ5QEp5CBYa52Vq5y0qr
lVxpet5NjsxHhHE3yigeTu4kTs5XTvF8GjqQSDJI6Dt0hinTl08CP1wiR+ODFkxyIwIyEPrjLy2D
UpoCCLhlaPPKpbP73BJwcZ3EwEERyTf5J373b/slcUiPbFAMi4Lq1vX760fcewV8OYnJ7Pt8pFnG
7hTxp6oNb932pLorWs+OlTjhwdmVWnNjXlSuU/zbDrxkVpuV1Rqi6W0lXqSNBieVGs/jzit+vnle
HmvayUHGKoRJ1pDzYolg5d32ZWFlztvEeQn/Kf7eyjYPxr1QGVb96YxBVey81ADTQeOveX+gXaOf
wOrZAESXZ2j6DgaQ9RbWisSSdyumAVKFrLApzFQfZC+QPhFRr5+Lsq3Cxd0oplxYpSG/wN36AheW
9BMQEaqA4whN+UrnAnAFfxUoUk5nT3nmvW+6vjoGTXcYjWmJnj1Pd98/RTP/EltlPj5bcsZYIpaf
w9FqycAxc2NM30B9A9qcayRW5q9037iMsJMlEfT2wnXDX+lzK746e8yq4epkNa3SQN6tryiwGBVw
iSgcAfNrdRek/pu6WKdA86ivU5hYk4yWmgPknLcEPtnEC+UeHgVdJjshsNLOdeYFqj0D7aRAIHru
7kvqnIYchsxInUy4ubq9aMrKFc4Tx66/YndLngb+oVrKUYUVXBJHDlg5Bql32ff0NQEcYte5OsWF
h+eWqrgQbGNNxdstagaC4k/sYoVraG2hgtRa8QFFN4eLAIYU7VTV5yu3L6gT+ixf8z1k0WuxOsor
bWt0fzDlmaNU3Th7J6FEqNwR+m4PSTHOBPlIrZNkrkDQmSVvKD84KXHtVew3jSrrqMSMytBjrTGV
9skOX9teFzEY+HlhjpLMpXcfAKGZ2YIeKEM+2wZGM7n4U/txBTbeCqiEq153SGKknNl4YS+zOJ0e
EE9Bg95YodlSojkzJtclIJAqsuXGR0cn4lfWZfmHopESmoM1I07P8BFitmncvQxBy3VQHJmwVwr0
RXnlER852MVk9A9lfDJyeFKCu8nbpORZhD+sPy5inftb5UP0uBSTtKsWuwKxEpYJEiy0t/SRQkSP
B4vVAEnt8Gg7GAuPcqcp+W06kyq9RfCc7jEeNEkABbIr4SMwTlK61oNj/ZD0tex3YLOS6ykCr5ni
Xq9HlPo8H7oOACornUujBIqcGBNz2biyiB3DaTC70wNsnCFZ1ek1o0nhZNFMjCEUpnJe7gTkQtUP
lu08sX8aU0/xStiDYE4DseFdcxF+YgAOzq9Wt6JZSLW4YXIQWCo12lFTQ/7ntXe24xPFhiosNqen
sG5IKvz+WoUD/AQkUSvI57iP0xga35865ZuSSEDKruAYY5t2uoJJdUrbjfU6VXzL6a66eKnwGclO
z7cVshvy8RxIKke/2YC5wJ/YVdE3vrpRZWZcHNQPxstlaUYW/3mt4UxklPP0bBMrKuPOy74wj4hT
doGGukv+LX3stZI+G951QGaZWRtt93uwbpWKEN5twn4oA6R3bR1j6pvWnWTC7ag+4gsGV+4YKQnX
m8kExW8eW/TqZHDiTR4rW0xCsrP6w8tx6xpVRbd+LNUGLzGl7uuIBWF4rMFhJl7FA74gRTmw1XSm
yJj1AjdWvS1WC6K6w2Nj3+avoEfAtv+Uc9urscGjbiAnoav00Rf2m2QppqCqBy8ylfh756yaJ71J
+jzSpqmInpz1e0qZlffS3aGddHurMklfAfckxk8b6x3VNonueX5lM5hVKcnzqUhkehk4elDKAgpj
GekUtEuwxFPAwTkr8JD2ovLbLy1ArzaPo2px3/DggTn4RtVmcWsVU7WgDHAr1zGPOkGlAHyipMSc
F52d5YD7vVvuKs46vzd+4YBWPDxHQRAWkXqhzyi9CHUaeu8v/fuho2o/JEl0s7xgf2hH/nFP37Jj
VpAx3s+cOZbCxZiUHmapJziDfx7dAO6dpv79uXlQEQF7XuvaqImEWMaBbZUBTQ6NxzlToG66BPwq
d5gObmDU/brtGVAye8Y3FHjJpBB2iOrbE/kQtrp5wcMG1KLun4XaGHkq6x8A2SDkrWSk4+Q4whMC
jzyG+vItTlMD+GIqlP9eZWGC8gqJxUbgNo5QbwIDNRDtbTOII+eCQ4bjUR7CyRdg3HPIxsj1nvdw
8n22iAp9dh+ZVQ+3oXFNCKogqjnd3+K0N2tPPFTTReZDpdMSh2JUZRLvxJlpxVUx3tQx0AwGsd+O
KFH64ZcF8CCWG6yUHljWJnnOFqhPuBLytiUa3maS01/OSKWl5C9mdDfFoovxfgKEm/6TwHW8tuw+
cNrTm0T0eeVW94Mcbcple5a1b8Gn35Yk9xD3vXcGBkXCcSMKNL/mBWSYFWP89OhRvTrwr7lBPLnr
UrCddKkbqFwQFg42Cnx+1HIZBsQsR+v4amTw9O+JD8yCNsDxoEIzA79cGaNvHq4sql/lSyBiVA0S
uhvhVM0llD7aBR4PDHuwhV7KJK8GwHIANM8MMlNOjd9Jn8KrWZn9LKXec5lVcXuIewTJk1wiE693
l4FTHGGce4Z8vBbsLN9aV1VQdLM9kn54txld6+8NZodX7ji2TGGceaKXLKw3g3jcUx4m865OPbzX
iNP3wiZndfey6Y5HFRuVR19PZrhHOyA4XDXrXKGi8AtgKmJK0FkW9EwoO5Dy9rNS/WgKYlRGXIOU
tFourZRqt2Ccp9K+at6AOCZlvqw3xk7hrmeinlfs5hBtNz6jQSFHZfYWCDxMswRINCfdkIMVMnXB
/9aAPYDVqYUUf3nriyCR9Tpp6qnBY23ExWfZJ+7kBliArVWzJUhNbtjwfsYGHsjCJOOGvDsBhE3v
vEXLCNTTmBL2qtXSFjaIYuc6JvP1i3x4JVyxKrcEg1HOuhzvY9IiMreYY6yoj4zm7KzejNDq+4cJ
wxfUzwSdqVA7dBHO/GP8MJ3u/uZf23WCVbTsVGsAO+MJUfLKhn0+IQGpdBxEWKV+8bjPMMDo4qqd
HQKBl8i6truiS/BIip5zHexCR59Km/dPtyrAkMBMh2Vcix87d7ppcj89W/CQc1Wf5ClJrtPft/9o
v0Ipjl755QmQFh43Fs2MnjZi1pzsY1WdhrppMZt4CrEwMYR+xuyucg2tdxxPpuCQqXpzsn65RQVG
rkKpj6JrV1XKDAS2+TVd/HBZCS0I03aHtkQ0oLHiPNohVpEGVL4/+fXpXuLHNgA9cjzgK0Yh4raY
8AMeFvcuM1MAebcDA9DpNh9I7kqPGS6w7mQR8bxDUCgsXPSpfL54l6hWmwr8M00yqcIqF5w6Sd39
bSgXYmb5PnIQPL6FXfJbaO+we/lyXLiOKRDlkGSECA7QMdiueqGFwsX7nGy+dwOQQxs2Fz2gFULu
2uM59oonh4Zr9KEp1OIYihCzCM70uSRUvBNZJqIvgy4UtMk7VZvRp3v+0hF2x+m6jOXYSQ6UsxkY
GEQgfetzegpmO0OaF5NNwlQxbZSZkgUzB3M49mL3dlKdRqY/4K27LLQOMwgaWNGzjGBb2aD4gTDL
OURXOEC8ZJjdM7PSd2nBbFcYNAvQlGs0brJCh28d3TMK1OFUvv5ypT14LkeVT5GiW4E94+GBUKf0
smbrUl2idDSPVAMM/giuhlYn/4J4NgoA6enStSgxHIzhJimBV+ogj+mbowEDOepR9iejrAru4khL
SUZ/MpaRYsjZCuFmEmCG9Ibk+QXsDCes1cBWO0c8Q2LjAgZRt/EMNq7Ds6mULNvBV99BN/s2g4fd
m7kmR2C4i63WhcABA04JqO1E3vEUn01dcfTKTk7z2hfjlwVFKRozzzsG4JEj1KQKUnHbadcIBvsY
FVIjjb9xNMwGa1FS7vDBj0w+iKkJNBvslDRNCuk9s0Tf0D1lLNjadDxEh4QcuYCpTRhFpdEegTfB
BQEP8yGsNQzDSss2yVrqgn/NWs2ykRj9BDwkXXpKmuyIz3MrlMxH8FdpS0o/lMa/ORL9UrIquyQ+
DjiSe8AcTUag1NFNYc0S5a9TWpgtryxVr+0AIuUCpz3uxqjgsBIGn7vGs0tZntaIbZxVt+SKTnJ+
vr/iiAipj70KF4goeaXd0PNSXZ1q6bCkFPPEsHBOP1OrM3KJQITSZ3a1oZ7SI1stuMN+XE3S8d03
02m3O4vulov86xc6CtBSyGBAHZztOzwPos47lCPd+/DUf9b815yjeALN1jnaOyOwEOIL0qM0BEb7
53Ud87KlbiIdTfvw0LXJzX0c5X63/67mPChBj0AR2WQzM3uSuIrPSkYEdEn2v5Jn+IoKl+c0QRIn
jG+Fk3cbo8c71PLeaLJ+n2/9030atcghDyqZNwIOnX45DmhKVZcpqJtSdUU3+oBrzULIqoJleyEY
DE6S7EAYfUpt4H0WySwN969ptzhl45dPTm6zHWfpcWlVO5rKgiWr6xaPJ496YQdzozWOd/gafZVy
Jmz01CTkELNaokYTLDNmJfQXgzK/06amMKpkHoIT5ywJ1THLb6N57ZiG+5wbBLyw8kBVx2i3PEvR
Rcd5kJtwF46pDgK5wECXoNVQpcT1bbqxOnqKt1wcigCGwyD3eaTvvzzq6X2RUDV5GMtEa5z5jACn
kpId2OETxxLXOWVwvfcdEkqJypE2k/rsDeJwEmm2sPKCCJsLEvcQqmx9nyn7c1TRPb4uPVrN6iJL
yztr+W/s+LfKh5ckyWFJdUdAgo6gTI9fS4N5k8kIWFtWKpynBIZ6BnI6gilU1JsrdfT9q80nLT9D
KnPi2kdtT8PZ5Brwna9TKIgmhdXUt1dHRrMnSaJGPwvx7J8i8aOZusaYtsAvwG7Uhi8QLpaWHm8M
+BtU2NOfzanfmK1zZqchYGq5cL+uq3DPi85nH56FDC+uwdF3b9JRcxwAmLMjDK68XYMYYx2/wtWR
dLBNwtkl4MzGTqCxY83ZaftPc6LUQt+2qdehWquMFLkBG2hd5fh8/AYCiHFxfpMKbFqg2nfGeAe3
5DzwUhKEAUyxJyLhnt2urmzYDMGcsNvkeTtgqyyyJalKuexi01DvlUvVcxNECF2Z5J84dJKyYeoh
Dwaz32GYTNVlRrzw6rMQ/L4qbit3Lvl1zWQwJ5Xb5TQCYXBv23pcWqlBvefIVRb+AVbllFROq+Oa
VlEHDZdzzRlScQ7DCF8Q1nRpRhgRJkzBIdtX4t7vpcobQ3P+nXDwDCf0qKKhi8iE0/zeG25peb4l
4tUoqVeZrEqNBOFk4vUFaaNC/QfdKZJ0AmTZFLsP3ShG4ITq3oLx5la47EWf93G6ThqVskQ2CLVi
EAbwOrZj/1ccRjrNI9DKgds44mRia0PwdYlSMyKZfs5c81tUmGdsUfsKHUFnHeHfoxD6TNh/B3Ys
UZvSBaIdADDNG6O6Ms/JoaS6tIJ08X1HXpTAse2Wf97P0bVi+oYdSxMGPflQfsE3IuVy7Ut6FFv3
Gwq+j+VE9q2ptkQvqqeXwGLOAkYuxzI6b15fBhgqotZ3Q3vw6nD6BgDULS71wtQyR8mTjzz8UAal
c8O5iyTd0i2mjC3Jr95wLeQJBBUv8OyaVIdUjbCpo9zVT0ApdDT0RlCR3kVe1z9Q/h5Ji/5nnjLk
B9ae0N6v/n/tYiTdvWTw25MAiBNREWcd1QbdtTbHU7JiL8+evIiRRfHSEf5nR4+F5hbgaQRfCcDx
9Ym8F5BGV8w5G1+9JuPY+UsvLnLJHXOQg5iqNsqL9a+1fs6gmBxJ/QtI4SRnkqnjMTzst3ExJi8u
A9eFAekXo3K8ZiEbcni/ZwzrFU4PPZipHzEI4mtnmTiyTtE1nZCoQyQI3M+w+SUnd5/goZ46zs46
4xZU6twHSxPICfN5TpuhDQbnWGgaFN61kg3jmn3eLp9FoyUrrxTb3nttPfUvffhqsT9Sn6LsGUvB
KSBEHcYvA42ghgRfneMsrogPEJP6X8PvTmdxhod0y3jgUsBWWetFxaAQLeYkNyy1C+7mTeulveQf
n76AmKMbMKJYsikNDoSE1p1Dshk5hf/Fy0YQbYhM0Z0faGJ48EqcJHQ584nChKR8rr27P9fGewsv
yCsC41PxIVxz+kEmPO4mbfnYh3MPf7pecAs1tH7PtH87aPitOLP1urHQhEDED832Gn7AGUs46gNC
6i6IzMxHwuJxCfsTNBhy/+gOQjnqYq9yGvm+t2WffjpYEMcOi2sS8cZWoGvpYX/ydETm+6KmKWDU
YjIghyFjvALZPr2vXeEYKuZK/lNj0nTjk1OLyeM1n3mO6ktd+E3mM7xpBwL0xLGtzL6bI9asFc+F
cc7s6CiC8ErklHhwErogQ492qKSmmIPtFfMc6nPBoIple0cC7oOemdtZ5CkY472mk8BfEUj4HyNU
G/3ChDs/yEhq92uyeqGU7OI7llXFQ5DIzZDT6Iq9yOPN9AJHPsp6yFA5w8Vl9qKwHF2NZeRGKQCh
k32Yh5GctKG+zRV0FCbaCL6dIxv2pT8tpYNnaOrj2Ct2aeCFyY5OTGJjnVy3NbhVb6VKGL4ykIsN
1UZ1k0yOez1tE5fs0NqWnpnTOpnSWhYPeXyWi9tUXQqMhFC4Dird6g50SzdJSZfAaKwHGZ2i2ysG
NV+2e1j0aV3tSco6l/u/Pm3rNVu8u45VUMVkP/nExjWI+ffhL6qS1ulFeWAozPF7yxNVHpQ5ZHJ4
Y6yOWFsMAFnSJ6w5B3K6C4x7QrFlEZmZXoYSaanEhyYM0a7KfpIzMuPs1Vtl8oPh12Tte0uR/5Tn
ZVMuDiHhSH8gxZqvBB0Rt6ASJfSxglFkYtMtp/d69ckTfatyNbFaSW0r83zWunPKGDptjVI2cmZq
f8iv8p0r2P1vQrWkfs2ZsP3BBoxnMTnaZux0EQNbIG8snbz37ZILw4UCjYVAGgxZRW9agQ0dsko6
qwHDjLnBLOT/QpkpKlz3h/nA+In95i2gg42wa2UZ3ZZ8+IQtHy5/7FWmrC69IPvHzgvjD2Lc45Ih
Wq0xutpdVJ8bGigGG/KB6bxzRtri5tH8un9dL2Rp3EQQGdYFEt1aiWrdG5SGt/JXk7OyWJ2GhrAg
l71OFANRMFd8UtUNX8FfESXSOGR8DJPQx/bZ9jWxQBw9gN02dbdWjx965UQUPDFlJiCZ9LHLPQEj
bZiJam7Xgs+SvZpd/q6mnEsjtwFMBgreLYL31PO12IBcUR4tV9wB7DlKv/uY05gJkzmgYA0gUBmz
nVjofcEgLG0eizx8/nQy4zguh+BTnxBvoVEYbt8WNBiG91vTdgefzRC7qb3tpUHXFf1mzmXmCpjv
4V8QDCZMkPRDqHO5XVcPTnCltpQVWZJFi59Fk/586ZacRtoa0Q4hX1S9iJGwLNQVLx2aIrFQkIbv
yIpm5JDel77xOl2/t/AFjYxafhMzFUJLCe6GhAJt6pn4WagCH23XV7VCjMnnyxTGmm+Ak/WuyT4M
TEp2lsWqckIKot8kZ0HIPRNZPZsHnpScWpwXArxf53POoUAK0s8sazS0YchTMr0FbLOfs75jZgNZ
i2hZndHXTiJDHrOvilqyP8TGwwlehqI8sgb8xDZJr5Oy8+8vsrFtlbkboSbpfDZOtq9Qc0OupEQp
yBvApHLgkwEmYaMStl+TCmfjxCsq40RFO/ZhdSa8QhKGUkeVBDIs09ovGtFraMcUJY+seTxl1nU+
hwMoX7bpzeqHLpjPjCLNd0gGQPjbrOrTsPa5wb1hyojOVtbbJMs1dpXFrO3hrmG1RVMANGTJabKx
lP8Uxiy7lRedNKyptDLSWHVx1epLrLhDIF7J65fh1H4daP8AjYMBi5JlZO0CC1Z40u0nD6t9lGjd
g9FNwO7XrofVn2EmUtjklveMspANnzGkXLl3Yg5inCAOmwmePJswB/8X7AD6I8zWj209GD1P2kEK
TqUmqs4WCdPlcRKb716R8sbtelM6znZNqb+Vo0DmMrLl55JI+0fTVO/XPIohWpgB4YhoLyoL6+4r
XO5cTzxSQpChXOIRrAFnnGW5dnRc6y23Xq0bxGfhuEQoxZqSj23awqnsBusboXvY0o/KZERAzx4C
FR9Vqt+wnVvKS3WsgEjYOl1T/7Df+r40asT+yjqM/7F806nmIf8CJJ/Bq+oN7EiUE5TwMmRe0NAn
2rBdDHkWH3HpBCCyLkdO7oKzogBvtV89ulILn0UwJTrmMW8SCRA3OZyqbtST1QmACh443PKxw2A1
bBdLijpEkFqKoXV7kxDP1tW8jpsjNi9FpVG5KVSce6OX6Zk1NrkMFw/IWsjV8My3OxFqX6xMFovF
2Sls+ZQCy1j1yBGU5ro6x+uodJrAotpIkM556TcLKWT+7TXgyUqSeZK6mVmBokft5aXzilN9JAbO
RIE0TJ2BHMU54An69NzRBL97ZBk2yG8Zo+bQ13yo/uoSjKpBJThUs6e6PzovGrs18DW8pVTjIMyW
y1yxz+zZfNOhu2dcst0NQw7mQJUzpfn6AtR63YtQnJbBbOMPjwOaFWWxclri4YgG6tm52Hp1Ygjh
tw+S5DKKx82K9/1NScSjJOIkm4MURpPh8s5Oo3/w/aA0Y6pQPbwyypTJL4+yGYHDrBTjZfARdsii
uvRWf3zeh0VeurYjGvnXpmaIfN1SIRvq/gaQUkGUkND3LazLKeSnnsdZ1v2uu87Jkua7M1wIMcfw
nuy5jrD9rh0ZldS7X0OP2hlqDN5UIP8GXHDABc8SxCZkYh2a2Pf5Mvo2AfyJvMLmBY6B0c/9CQMY
DieW5VO1kAElQ5+pBEW6wO9ylG6rvXKReQxSSZO7Cc18G05jVZQLiE7LzP8dIzyBT9vndobLgtFL
PSSAv3+ebXMhHp9/u+3LFaWZwEncuf6XzgyOb6P7p3h75TlCEjiqLoUZiuZ6oTGYfI1hO0Y0aQVr
EXE9l/Xlo2fuLKx73xmjg0YmaXYkzMEGOvEmqDSqdi+tbFyGVoiuc4phEj9q0iR/ck7VUrxHiqy1
l2N1FyUkouZ2dQF4Qw3qCOZylq7RgcLhuXWHdKdQo7lWwxulUVQe5NtzJdCRR+hUISsvwv0nX0bM
B3ESFszW6azSuEKsRu1LTtiCdH5FsQiOxmmVkekQGBo5zdksCQ9IYRh3ZkbfqqZVMhuG++qfx95q
2D1Yd6qqdC4nhDh/+tlSdr29Q8dGXJwP/a1Izf5HkA8hJjlkD/X15Vcr0VW3X740oCy51bV/WIfn
ndiyzc7x5KegIT4LrVvYMsZA36SqjG8aIRFM7IE3EP38EPjlzPsm33xpQJOtUrN1PQmypN0UGSxC
fuLcVk5+/YOsEbDC327kcvXdsdPI4sJy24JWYTSqnn13g87AQWrD5cgFvD1YDsX/TZzzdTdqiXKJ
+A1++zMU41QcwAjPCO+CkrW99KsnFuxKM8NWL93D0NooMupBaYbOM5Qe+SBCyAoKwxYAYP5odrEB
T3KW+RcToeymc0plt+iDi9ystaBqZ9rchYNIz502RQ3oQyPxGcv1BgPbHhrenObrI0qHCMpWIof9
QkKqHSQxG1x4fKqdX3q+bGSVJQt50FvTKRkxlemfxmvo+Af9hOuxZvCeDCOx9FNA2o0avIk6SuXd
/faldc3dG9z76gJqIeeiUQ7Q+F0iq5DkidJmre6TY4mw8sCWF4jLOhwLnUfBWWgD8YHXvP1iYvYg
2pKttcO38w2/m87DBNwm8ETR/xaxDkT8O6o+eGbCcxjFZO3pkTbYJzWauT4ywzBMwvKKfGKECrEs
E1bUVbIZjKejaHhn/F7z9brpAwLlNWdt2peMNc6QXSc9uUaHp1umbws8+PvisMowTEgtm876JV0q
OcEBJf4koK79rkaAMUZyd/llIS9rdEoOBBRQhCe+7X+8jaAWfl67KCEAsJSrUDj0HAof2v9TW/S9
Pw3SgD6VHcninOWp5D3DnRWFPYWubHn+0+J52Oxo1nvoyBaHptfhnUaiY/AlglsYb5lFnyqLt+id
tpfYw3BUN4a8F34HiytuJAUbLSVdYQSEDnTXoKbnNHxytHA/aVyKJ4EbctcCki/tSa50psFR3WW2
YMsudbd94zuiFPnEMJb3hHOA9A3vUlfmbvN7jV7mr0dbutCcUFl77pqbMb4cJ/koCGC1cdobAW/Z
C0p7ngXY3NcnLxDXx9ZWaBwfIWIuFDUcRGsoRZZouQua/c86k8QCTre5sMDugVkDn70KMrDu295/
O/f0OCkyL9RUD2jh3Sl8O+SmgF2yItZ9Fkg0RG2Y29w0CjcGaocSwRHfO1c5PkqK+LwijgymgDVy
XZiDhIcLHVMC5ZvR6supbSMUZd4coCF/VgPMtXjzdlG6d5VYsQZaf6nZDJI1uclsPp7+si9tbJFM
U/dIneUGeb+ckfOcpKgynE3SlDi4B4mXACtU4j34yf3zgPMJ1kt2TKgFHDy2Tk0fBM/FCaMqhY7K
X3Ic+gpB+21+q5bPEcE6Y9kvV3vUya9oHASHnsdb8K+IDZ2r/5VHFSOVVsAKbun+0vhQphsRXB/e
4XbXU3QI1dxpf5QrZDbGEqQ742UOwlS541yFx20mX2tyS9hPi0qiffAAPJsBYVBsCfnQfC7slbQc
OrPqT75HlOB+O+q6wiDuRQX61aekuzDYNEcpMwytbWWo3L6vaHN8nZt4TFfvYJ7BvrR5TPsqLkSX
RwJSwP0PnTm9kxZuonil3CyLJdS1RQPONHj0On+xCDFEd/6LwTPbOTeS2j9WYe4jqq9h59xsdWvf
2HK3wztcEgCu55QGpSdUa3DIfKO/t7Fi7pP9sTvp2JUziNJSJtq/M5L3pCkVbqPF96LDyk7ceVAh
K+iDJYTA870DrdKEY0jEcJswcFFwaT+oxtMdPkHywXSDOMkByzdPsmHb+azN8hujmA0Vosh/cDuV
fLWvXdZxsnNvkAP/nw6UOOq1bQj82DA5LPFz/+pr4EFxL4SbolzT5yOJCSvl9IwugazQpsk94FvT
w84hoS7GMYMjE/CzRsnCER+oVjAaau/TGca5sKXv7nH+XJx+Jr5FI4SHk3T7aJJ/OUVX8VBhDqho
5hvnFUrjePERjruGi01OdZbTtony3qhbmihlPjXrx2FAMp5YsoF2w+DlRvG7uXRWmF6LZ2Ke5Nl3
hOOHnXyn0cKAENnOXWFh8ivW0YxidJ5RvO3NSLMQndJx6njwRqj+IaHD1l3Qya8u3zNIWi45vdQH
MHMaHnjnCyMr1ZiSLIlEb9lJ5J/7ECSukQRux/FKCWit39qPxeXkT0k7YJlahBbN1KWP0JzRaQhl
s9LFQSVN5OKnEqcHQOgv6LfGRaOdJ6UU0G1B6Kl265F/pSD+mjRK6Lbwgzgy8DfheQOExjS3uO/D
xoeesMX8JssQcfnriBYhsgUuGo0eRWuhmAhhJPaiP3snbbKb2dcWHr5HJ8fbDg9EwDYyzqlFCxUw
kRa+wosymdLwKGq06mMzN6cNOFZPRtsKsssSFXFVLUKOkbuKPB9DPkOgMxUJPWhF/rZsYRQ8Yc1a
j3WqiTs5F71yKff1i2y79keUeUnZ7YnS6OWbURfq05TP++bH+RDhFoldlRXxa5oYIj3YOJ7rZDOj
czH3RaT2OWnd256LKVwidi3KikmrwxrJXygImjvFV5fmoXLPD9RDC/Kk2bjiLbBsMAeES/5NJ08+
YCR1KKcXDIoBK9eMq1Evr7quOD5VH9pYRMbZVWDOzi1Gq+GJWnSwpVxU4F6C/UmhSLGX2l1jMZQ1
t/EQkgUWQBnaGVhti6tjls4x9o/YEdvS/fdKVwW8Cf0/Frq64IOch7cB4ewHgpYB82NF4K/yG0aR
ZIoI4juq9PEdXzycVZdhCAndSwuV5qiy4NsZGwi5KtiEkTloJYjCqGF2mNWHxhA17g+XH8QEpyrE
x1NNcupnp03MFFZ+15JjTZlrVw/CXOWNOThw+T70FDXxTABCJpufa6UD7qaNFvk158sRzyy0Q5kn
3rZaXu62qdHbwlGclnnIPpG2xGVkn9s/6MTWMT/m1u3XPTx1JWlaoC1XlF8Cdaq0mPKg6+10pr4D
2W+B8dDFTH9gbnD+sfbpIxQBWdChEJjJEq+rtelfhfcPoZIivlJZtPUxJQ0UeV2jZLg9MD2FPWgD
wXLwQQpgwfrExQ6ZTHHg87d6K72bV6anVqz5WDLr182tdCBaPa1UnEV+vPOHyPvlCEqUWPuIuWXm
odXRM1Q+XIAR3LQB42CMj7ITlEujSihNs+EChEIqtcUh/aRL3NqvwHOMHF9+oPEa7+UcwPEBtB4Q
9/lzQz3Xeg6LIZHojWYP1q4D1BbPJPA3syYiNNWdpeGdMbooO/QAOhHkgewdJzIXqefjYrxim45M
IQUrpDSADiLVAicmU6or7YNI0MV97rNqDewAJht/LOLEghmRQoR4lAlvgzkA7GKLEDwti2KHh/SV
WgIYftl0n8K+iiZIpK58TjSETAxCQCs9BPDfYRyw8RbKmkm0OPPWnJfLgIHRmePI+Ixzjw8LfF4v
VuRRK8T+RFmvhAUOccFFfTzKv6BwMRq4g9tADELxJoLOEpJJEjVTyIl9accxx6zLurC8eazsM8r4
gO08T0pijQ+cEwm5r+psHSHjKgrIyn7qlUjiB9nGnke4k/Y17NWxLFLiqXH+29/fMjyEsdE0pl2L
rEqdcAo9zyFP7FrLDsXZh+RL/Nauq+XWflkYhoKfdW2UvxjPiv3HlkIFYzbNJHZzN4+9RzmDqy7H
lemLNT0dkH+L5hsO0DhRaC1X3sT+uCXzwChfKd18aZf8peg8R3qnSHgJ5aTrPxnHe9s3/+iRlj+3
SkEjJU/FXXdfi3VxUrEkOg+Eqa0CaNbdV9qJCAJWp6HoUGNZV+BYoDa2HoUmwdE0t7J8eJZAjAgZ
BHJCi/l+pPiZL6gZ1iaUcEraf2JYOFGbDyHXCJ2PZgr6IkgXbEjgaOxPDkYFq9iVPImL79JTggek
ddG1Vc77sXH0uHz8z152nZukTi/CQQJC/3wWJJ9CGYFOHV4K0WmlhpmuPiU/KZBV0e4l1ZXaKX4O
uZh5QWgbiiCI/GkFu+koSbcgNj2yy2V2SmrsBTHV+e0bLOgo3rPwqYal5fT34PoVJ7m/7/kqDQTP
/AeukYGKsKXVpQ0WevyJqKZyJHjzcR/5IPzI4xnlfAAwjKruThONGyhmR8eBy41ug6YIBkPCqTn6
b6CjpP+FSV2BB1Set8bd/jWjKgQoUigO3NpuQFkkWFULVEbQVrxGI7Uf7NTIPLiaD/t9bF6ucA/2
EcoSG4AA//V6RnFzPO4Wr2LZu6QOEkYw35cwrIj83qOSOWNP8yXf/rBjwcQINo3J+3OXcmQN76C1
sLlXvF4hltdxKlnuAE9hU8hKrBe9kCWMzLhOjSIloFL8HfO0S6q243ZsQ1Erngl7T5mY1mlxXeNJ
BQEvVWFwKLpUO5USZ2ss0pw9HL8wJweKRpVv3/f+Qr4wlAGahpnJcQK89pm3HNO+udO6f1ArMBE7
DcrGaru2Nsf8/E3nUo27NHquf48k5jcoxUJtC88u3uBvH7K5itNz62fE4PrbsNgQAKc5Nyrkhkmz
vvKZ6DV3uG09l9VDo5jrO6CSuwAHgRIOpKBM66gyBnJyZE2+/vRu8mPqq6XtmCAwEQL3gm/Yy0nS
FIPNvVfXpCIKJkB0+m9N1w5EYeGySXpc+2zUEz7EMSAQlRApE5W1bFKccYf1PffXmoPHiTW2a2Ig
L7G0HQ78s37dQPwGQ78BWwpPAOo+CZ2njKJPu71mF0UhHU49AWAUzmqn5kLx+VJeJt5rtuEakMsh
nvzaLsgCOtZ6JW5QfLl4uwTQK99RgUKrgOWukZ2lqwpqAYpgRsPQKMzqKRKoP6Y0RJC7K9Sig5CQ
Rq+tXrDcDWFxOQy4Ty22AjQOkcBdZ3kCd6wa2hKD8mXNhs9XMz2sKFINGUyuXQbYPrZxbXOiMIx5
wfdEgFFIZrFHc1pD8RsnbLfdxEHF1z89YnEjCO67exAOYd5qsrH0gpK2gCLd1F/WvsVtkWnhVBdb
XrhHuRuAoCB88ftWO5XEf4ZTrUtMmpf+muApeieG2iQhZLmCWb+WwoA4Tjw5ZS3XVmbiidqsEnJX
1bcGMpT3zeemfle3lCfAAs0ZUuGAViPzkH0aPXKH/jkxFTY2xbU2S/81onFL2p3tizhXvy7GGnTY
7vN/2mTTTJdARA9ayNG417nyhUFsqB+hEPZncnl689Qmo9I9hvtFENvFdfOBlmB0tln/0lazmv9j
A5sdKAFv5zud88DQ+t8ggMMyIb6zHa4yNXTtREB4LvmrX3I8bqgiO7QxngyogQ9VS8upZyftQ1fv
wYjk38Xp+n7tZ1vG5WCKHHnswTB70aT6h1JQcyQV0bjm8x5rlphweDEoRnbSXVWouD8DoA3d3sxq
p02HwFmtCvPEmvcvJ7Y7oZZ9IfT8nfO251d0lkwRELxto9h9RRSOOq+sQvSNhF6aViqHs2FNzmyj
qcTr6IqJC0eCInFYOFdrGwOzWDnhkFXRwkQF2ODF8lDe4YqJ/GcXzoPGfiI+4Dqe3u98V4uH2Fqu
QY6QB07Kw/DR+sdFbWcES96RwzxZxLkYQpQ7xldxiUyeDPQTyOXEKGtAHL1TwbmOXNaZrhRXaxeK
whX70oBTkWI7rlCrlNyx/kDkQP5dfu/a5jqL5sWoh62WtVGwUp3nsy+y+f/I+iyBQUu3YWYaaotA
CF6DDi+Ls/Crn6GFZR3q6qhdzLmgbr8+VnzLGIIQSzCdkFbL/FUzH0QWLTZ5e+I4Vr0L/3ViJ25k
BYk8Ucpd1nxulP4+ZwaRt6MQywBdhSVyOoIUfbMzntNivHM18QQswnN0KKl451qCFe/9qfrt0z9N
pZwWoJfIz8IZ/E/PLYuAIPKpe7qRX6XZEXQW2T6fDLZ0CqffsTgPOK1R6wHSZImH/H4pjPHmW7Qr
9EjXD4WVuVpsfNoTllMolnSdnAaQShdjRfGq0st/U9KB3vcsu/lfh4gV4wYZiXD52fiMBncY3yGi
31BGVQ938nNmLTFmqRHYcSb50giEYlgIK7P99H/z7JUgY7zyEyx/gXVOEwqoSVJCLITkvYE9beVN
MuD08UQHhaSWT4LmLqudUICIejFCIR4/j7VrhEcFEaN8oIbrdfGKJBv3AOQdgFEUN6aQmkobuLZV
OO5/X8BVl0WL1QyIJsPZijNG/db9BC34WlDMB6wX1SJlksqoEUrRnpJp2g4J+ZbeU24K5bLXXKGt
+qcMFbxK0Gw6I8gvfN0DIn5+DFbVQNMkoe+fjfIxB9bb4XBkgKZ4dYtaVrc1gNk5f0/Fhz7kfRsc
XzG5G/BKKMkbaAO4pzdZk4N6NcNQPnEaVjEl0roVKSs9bv+IGkJCFqoHKDkCWc45MTY5LesWWJ/o
TMcyvXomqY9c2Cy0I/3t28sEm4aBz4MAqc82GxQE/A7NPxRklodNvLvFCR6iYK8Y+dCl9/z7NUd8
s8mw3IV7GTLfE4JraO8E2Zd3PYerlXWBgIoezuKGZeuk8m0me6+lDR7pR3qc8FO5CzxGa7omlgUF
5StARhQNsAIm4crbR+eVWipHFvfA32w9FvvCjCzODIU5gBptcJVMsMbLuKs/EoZiH2GtZds5qRYi
jR3gGz9NJV0TJ0LhRR6fhO9o7045I3bZ0wALxh+/YcEG1ukNfUzf3oBCL1ckkf8ljLst8sPSWSQi
irfUT0mBa2d313MkGm5lGdQOX3RGtWRPcruaM/2XBYKE0ZUn9ep4wctZ+yK+OuodNMZsSAyaiURn
DLHAqvRydHDbInmrN4tMatxHZv6KIMjZJI61z4WTEhVosh+GmdijJU5qROs0oMue/IkoM+X1GNf8
kLsHRUGLQXYqZTMseVNO6vB/3pECrJoIufPUGaFlXfec4t1+3PAxa6JkqYSFCto1oA5tkMI/5cmu
9FT4MKaM3EyzzyApI7mPR+FEZtjE4+6QTULyUVuInk8X931yBf8VZwpmrxqYPbj0Z8igtD4SDvVs
OYMKiSsTr7n8dN621Y/mNREk5JDFr0SI71IMATO4J4C3UCQt7OYE/23YBfU0jNT0qw2VknljfqJK
IAPrXA9BT41dP2m3gUPDxIL4ajeVgDb+R4K/BV6e22g91BLLJBxCxuxVUvxgOVCKTrHpuFlu0ksE
RbGHzzVSFHwWwQ0md8ZMSxqw/uPExPWyuAswSV4drgU5BbgdnpViQspv+5d1IrHhZjAl4ZYDn/pY
Htm4HwLlEUI6DaCuwj2J0TjJmwjIP5+BwpRUfKGIH2i5YAe82AaocJfPzUI0jzj3yyzTRwH285wY
EfuvbJWG9FxfR6lZH/HoArmWMEmMbbBHKPzu2nOWoi9VaItqqd35th1SDJop7ylM19x8jjdPpNNF
lJwP6ojsdyeZlWk9MP/4x6xf/gn87j8xztMfn9g7SmOudWC9IOGkUbfYNC32MBKSMBMmVP8FNXCY
bNDgmKx32i/wbWF9HN2XANkCVa4f0PsUiWQ97hx66sIc1LVNjffV6TxFD5wkfRMe4pqZYdmd5nUK
4aoD+IPXZGZEe/HENUlivywlNmEOaC9Zy4RoEkx0z0GGrGoFq56uoEAvsdTaD4XzyiY7s1c1o7xe
GNXwJQp9uGURfryt5BGgIHEPjoA3LcfuPqZuZahehSa6I7aznAOudcsZuToE6cahZjTGaOJT00mT
i4mUon+M51F3vaV8GHtSHdFayH/nAHGJsvam9Qy4HOASQL45WCEoVHgzkubdAtKj5MkNyqnhDWFM
oHScvUyaCkfqn0HPkMDzRMWld/r6GyjlUdIRIMefBD/b9KBmb5nir5k0plHVhhMvTHhQ0uZjuHJx
N6SbBLyg4IANencjZg2bpCzKnrY83lukhZpaci16wxPeHtyQ+7B2MMJZk15DEA3hfm5FQ1ZPFgtw
949qg2IM5odDWCKwq2xbfusN5cW7lch/lFgui56Gcz9piiqXJnEgdEmBzQXw5DOH2xQWl2OWaTMD
mFdb41trZe2Zqt3DG/sYkgd/AnqzEhyprluLpk0Opv1G+wKtG7iHyW6wplZBN8qX0YA+L2ji4y26
qKWKuG1C4svj69BEh+3wNAaW3s3cByNrA9ISpfJH2iPBsLyCY3JuJls5vD0B1ws8ojpmxyG0zgLQ
/bOPYtUkmlNMUNcfHRJH5ACk+owv44ryQ6HKEY8nMJoB/fZn26vCzJc8en6xeBI1OnYT5qzvzr4n
5yZfrnHBvgoYVbCDpiTBJFFr13sIAeMMHo8T4o8n3/RT+Gs0Y+CQBGyssTwWYa17gFdt1Kr1RJ+n
puEHdwazFhFuyyDZ9RdSz7uGPu++VPEziCyPuh8iG3zWAqoTjL3VflJ655muxB17B1vsIT/BicQN
+y0Kju92gBkYClaPQcvXKt1HxeLxJUvFszgWtCu5GVyKMR+RVRap2yVTExwcqGe8pejfQnviTxc6
6U4cTjN6nvzLfCLFuzKzWil2WVCfYKlYHohUyqUcjFbZiwr8OaeyM9wy3fRF449Qp9nPFn5G7ylz
dOn5ftATm7Tkc73znx5SyoeSc/MsWHtCrie3xwq0jWCdrhB4kiYvr65c3mhK1e608yPaqj/rXKzY
yiEbnSTyCUy/Xczb0ATsi8KU/AvucqmkfJ5r1gFjaECbw75qXkIukE/mUY5kKDeQdVpC99ZDoxhA
475yi4IlfrXSgaGalSnp1dT8Af+eeOo0MKAxFMUo5juhC4fkaEi/rVTCxcK8d4wQ0gO7LAZIWF+g
2nn1QodnFmxmZfTD1kT77Syvv7t6nnb38a55yuVz2WGhq6zssg9cBW/hdI2eVRlF0O/BTRJ2TvFG
79ijff/exCpkVUCV9kEcXItbguxsOilYRi73fHW4h366QQOj1FrzHAt5j2UZUFgAzrwBSobncrTm
7pkmJFW7PkyOrs85XM3TnS7CYQhMmHcC4NJfp2sA7A88A92Rq7MBgJdLjd/QeEJiYOeH9S976ceH
h3/biCDJeprw0YgzX8E/2q/gfm2czP5bA0lFB1obBi1/YAlqc2C1nxqi7qT5ZoBLqHzM7iRhTyiS
6tuxygL0BUJCkQHUtEqIGsUYkqnjvpcHQrGUgYqbCc3o2cWO8FCdsRvHeSHk9htWoY+5/X3RGJdJ
2yaJ9xAWA/8u9lit3c914UdDQNK+Tq4q2rvSutwswapAZBEspigPoST6ANIdt6GPXOciW8pC/bbq
dvKkbA7k+m3j9V045uxRzkbve4xh0D2gXRlU6rH2JJXuDbpRp4YxO7tpU5ag0V1d1tlLhUafhzaI
/4MtJQ2fWtPyxUZqxCdi7+boxSXKEIxmEBiRE6wKo0SjDGn4yQsDut3MdrYpIH8PV5vF5iAcxrHF
Te0SebQqZIno9qZD6aexGI3mOc/LcuVmfuAb+9SXIOdoymMaogEJJ57AiGpnmabZzBKZEWx6BFWB
StHXxpqHJbt/x5M9sO0yQ84ARjNMjFdMpOxm/5KLDFN8un9J/xdRPcgb22YnyxFRx/CkiU7A5Zed
1SIcumuvRPR5Ij2MqETMiAl/Je7FhZfvEmW96Ve7g01XEyErn9dyv1heUHLrlVWfOfOJLSrNerp2
/feHl8dEpbUBISK4mYhONcNbCZFhHsmnXCQse7Ypsw/O8TtFHyO2Fa0X30G+OLyVFG6Dav0EpoG1
ST6mAlOGTk7pmS3QGzaAgeQ/HWlowiSsDDDuVVSYq9A1gOsUF9kGZeefEuUoBuM6nCF3PlYQflwS
9jCXqc8gKPwG7hHpsposo53Y76xCGO2ozuzMbFlBFtyDJdrAJFUFx929IoSDeEw0g+vDKg/qlieV
6lAdzJlF4kgtKc4UEp095oEWgktKjhQWcAmT9d4iqrtpdMsA5M+lmMuCcuSltk+bTXHOdmaT5L2q
5UeTmKtUZncETvbH1dHFqoU3XQfLZxHj2a31ldXJe10rrETlVu605fV09Sr3H9jpy6j5+MTlc/V9
Ri70BMjtkYuAavj7xQKQBi/+u6fHA/dy5tLDPvRkwm6UewQN6gmDKktrzUaUjIMZ8S6vGNsDL8qy
OZjGSnQ/fqJqiW5wIbGD+Tvj6+iDSGonXLw/3z0HjjZOKLzizUx0TJqyK9lawi2UveVoy8ujqb4i
xMD8WEQqthiWZRU6QH6CCbRtq/sie9TwjvvPw1obbJBEHFIePqhbruWm9y8MyLcJE7iwmP1kWe81
ertck9nlsO1y3e8DAZHqyfuT/7JNITVWbOGnpkThdw6O5FNtthJrNFn5TkjZDl1KOEEcRTyNu21t
6a8co6p/9EKFU4t0kGFAaIO5M8S7fMADqBpJ6qUMDS6t1zsQAKN+m1sBs3HtOEIw++g/xDwI/vAq
CM0YhQeb75bCC4KzSXJmi/J8SqzWo1DmvK01BwyhHfiiSNuWKr1zJ2YVoktmjWeSIz+JLR/jEf23
pYs2f8rYIBE4v+GoFiJFvi+K7J61SFFw4li2dhiPxrHxMG/Qf5ZqKcBwL1wMjqozfignXNi5OoGm
9CRqtXwe6d8EiYmEv+s0ZoiqeTatHK8+viG4DopwgMjaDuxAbgemEJ8OFXC6XXa7/3l9gC1OeYzd
8XMf6V6J9VOr0KAtMgoeh944l6x0Xd3VBugTNxP8ghEaEiH6ZwSWJ74os2uD/c6r+EKExMhYd3NP
4V/HRka0ZdhOaLPGMduXfRqWKgK0GxU79ipHoUio0JpRcTJLd/xiexk55oJX53rFFKJV7HwLVl1G
cJ0r7zPcNa/Xm/SA5HQPqysC1eEn7RX8CjqaxnyLjyb121rc8zhNPZ7tSqigm3PARnpfe/kN9Zcy
5yR2a6m+iswN2dmyHbFkQqB1x7/sRrPBq6rjlY6cYkGj9Buma514T+mDZo5o6w91GsnZ4u3IiHmL
/jcKRpWXal5rYhco2Hy2HZfmto7HZj3cE09pxrKfZjCwyUhRXrFEnse4pe/0jXMP7e5PW7Gw/K31
d5PzCnblgzvqYkoaZAcxVB8vjLz97SqhmIvsZgk/yShrc+DBpXo0uJLk+0I5JjnP4VcsFkUPjZI/
HCjLutDAVsSDXG2Nm1+RepTzMvgo/2y8Mwgd4jhzN8R4q3yaBEVhw34pQ8YxyvQTlz9aKvy6YOqc
xxEAmOdOLdHZvcR7w4zdvFy9Wr9DsiDXEC2S6TsnHJHV2jBFNtRpw8NpD4X3h1qtxvLX4bawc7i1
qRZnd+sMWyAn8ceZskd+R72YIHvrS/xCqjLthMzpQA3qnltUimft2bORAUnOvtj4BKwuHes6VoGN
luMawUY18M6+XfvV5eo3ptnmbe2t24GIQSnZHBwQRS+JfSj/iQlXl6CaO35J40VQlg3qTvVgBfdK
Q8Bc8QMZKVbS5ynejTmQuTGnROr50pRHigaFevkhdkAHfleFL+4H+GxfoXWfIhLhn5/0exusLPXB
ytoIJWBCs61lUED6VYWztyoSv2t/yKRMS+nKw6meSFZBr4CkztJIMBNirRHoBIxnb+pGN7lQsvVC
hJ6/NRYov4P9ilsxJnn0Clldotai5hdDhQr+DeOQ00xMo4Mk6eDFqBPa9zJdu/oAbQq9ZjsACEkh
d/E2n6hc/ISzZZjfaEXsgvuzbgFQ3cndkkwk9gO/RSS5MiQ0gB7bqs9hDnJSI5fu6l/1sg+RNvuA
KWhQE47wSmgCroZG8FkVW1HxpXoG2yVu3KLeaC95gz+XQJrG+yFwUlQpHbJOwYubrpw/YHbMwby+
8Owpcr6cByqnUmoLxqRnztmXGTwqi7qz1ssXR1pS/VcBCxieykurK++qZLY8nYX3aHp+cLje+2wb
DPlv6i5LTXUHSDJQFQ1NNap1zqjI9UGXLWyNWOIACCrSGFQcaQSerd+ON2pTe3GCyfGsUzKhMo5q
jbLMmmp7LLoRs8G40G7rvp35mRfWSYABEd/z1BhNTTsfzev2Mgw+xE3hkOtCf291bolv4ccA1XUR
7+2sGK8zNVBR8Dq3RY84UeA4RHqXqtEaTSbzyts1uWCwCsXW77rlmGlxb6wDV/v88A9nJyDNx9sz
bMNZeOuw6VkAG/gCXhvtf0/AZSxtQ7z9wvLO9aOEIqjXglq6pCHFAmBXiQrPsrIjOofozBRobb/8
6v/YOlniR7h5ZVKo0/LRXglE1zpKnJdP7pRAUIgJmnjSkFwJRc3Xzpq+tfM0578my5106Wdph4ji
VInARgIGdHznQ/oCxRSvZSp8y268bXJ+kHEhBenfidIPPPqhATtiXf06lWILNHibwMuRmg7U+hsA
oBpSs0qKVW9C0jUVIlXcpL8wLs6O6sOIRYAJvFvdu7VFyXzoFjdWwjfPx6YhapiQ/3frWDes2oKF
GRHLAEXpq4V91Oo3OnCDNRPb+hJTGjI4kl3SfFxIBOKo8DCC+VpFUHnFbDZ/aeTzOyZn6GxNfBdU
j2Y29lPqTd3L+TcXzL3U3omfkzmx16n/yAfBMAK5WcXkZzLa6A4tFYg0Pcl4db/IJ+SyxjinJnMS
4PlWq/06daHYK+WMv9ngsGwfMiGRIzeI9FMGrnPZRf/yl55G7ucJIGdvuh8kICwVMEHZJlf473dc
vkbmGRcaGwQ2PXEDZuMBKekjmgxOxeEsbFqM4ZF65oMx8QlAxXuySrIYO44FEtk2SGqsfB+rOTT5
vpbRk3Qh+4w65Gwv3kPZzNbt63rS2qo8POGs2ETUEzqxPRuw3thRzT0QeuUPKuGzsisiRFZ6LwVW
IOGIpr9nJrdaTpEboe8c5K3fWZaiDndNJsNnH81bhQWgBCMVJ2ekQvpZckZTBBwM3WIrqlU1MbEQ
v75TDdvah/aEqR9/97Y+cG99QT4j8L2Nx0ARmPl2ndIsBN+IUBwNEbrG9Tkb6NjVU0xbqGNng/oA
4CdaCRL3FnqDvWEuCfs72mY5MVDPv2TQnyQegFvp+9kB75TB4jxs2HuZcF2UyPMM2nU08E0My3mq
w2AO431ACTf8xqEQ7AZYH47oltgdVq2QsImHkEGaYu1vm6qWxeO2NeqR7eLVWFPxNAHKd+i/63R0
RJa4Bsuqk6JQ9dNxro920/BX0bdHqGcOFg8N54faug/WPukUIHo+KtQ936HK41ilIrjbcqNHnC5z
Ed77Yy/KI+B9useX3FkzZLxja8IwevqxC/qgzCTWgQ6IiJdKxBS4s7UwCC3S83tY5XWl0L6mUwkc
GgqW2YgvUMV8iQqfFuJ4kS4qKyT5wOVlK5culzGhzAKH5daG4mosAsDu5tV8QlV+NjT7oZK7yuQo
wNxKncXWUKzRiObOgFc1vv6Qy0Cmoj+mqXING3mWxm/E8MYCf1mEaj3T32IMt65akvNKRZAjW9Nx
i9VCt0Isx8bRGbOxdbkBo/uVu4czs5lrM/CIGEfqchejxRij4igtLctw1YLMgtjtkFQesKbzYCS+
6FNNZVrj4Dz/IOYp/M3bYPvvp2aLSV6dRmjv6H4vaULINOcGRGu0rddeGrYfNejqDT/wsa5uF1B0
bzakuTZSZ1pgKp57q/2JLaQXXCgzheD9idHShUOz/OeTL0IzWoWUzYtWlzjJFFd/OrSWzXFghZLr
IJ2pVAzIqUmo7y9x3f2Nya+JFd6hWCtMMvoIv6+gk34g0hwK0N+2sKssWB1Ny0fev1uSvU1xIGtg
pBmLnwlNEAFRf5bUtXAfIL/Cmbj/fFMgfdnZDfy5UoRCEp94CA35g8QxAkRCBzLKUHR0WcHP3/rN
iLEXryg3aQXLozhIElOixNOZnRjPsTWyJ6Z/uASZ1TAE9lxoolai13ltwPHEx4V//mCfRqiUCxWA
5xV+V9O0xgGOWY8da/I1rU/RCTQn0Db0QHbsH9eKiXtKy9fdVscaTF5I8IU3XYZTxGnSQYHIRSzV
fu81qYifWSli3p6OYrEy1wKKxMm8c1y4M9M+KUkaH6StxI9B1lnNOJTftbpXvp3xBVhTDmSEzfad
/fFotim1tjG8rOgRDFK+IrJ6mMjy3SsOiBK6fqE3o69rs2kVXHCPgfGItZOjqUIhYpKpRssIfo97
c1hCUtmV688jP8u3IyxSFz77eE71RXvEHkN+WPyIvbVClYLRDn6kZTAVmnPmIE1zaKkCK18ozWu+
wMANlFY9ZHG8W0rjO+WMl7S0yI+GDFxkBuAoMtbhjm3V9ttobEOGz53mjk1P8uZ3tHj6QrGA2gSS
FVFATCrwcj4bBCWWtxdQy6Os9t8V/vqBYLBCLEwnlzXlH4APGJ1UiCX2eVervFGNx6Tq3XnnonWR
U/g+gKWmgvVvw507UVIr60Y9BDZp/cOykcwEzjdCiHN5qJVdXO6UZH3fNBw+UyKGPOdrZ6sdZCY2
4JMYeJWWyImL/+fvKugDLM6q0PMi6A9AoZfk7OJF4x32kzsEwPd6AYdiLFChnBKncIb9CosASO30
KdYxTgmoBbIRW3VKD1oyLKJBz2LHXuTX/gicmd5CQWGqBlNVbsivx1FltqzYA4s9YUNTRgW3TwUj
jssDR7wEf54s5767IqhBDTXohg0a4J7y/ohsNeeBa4FvGvVMFET4H9D4rRAVkX5NQvvh2AeaalV9
GogVgenY7ibfx16TDASheFLh2InXRIQX1wGQTNakHyBQWAzCyZ+KD+gb6QKQv8y7GXHIG6NAhDq4
VEVDTchVyMNhV6BDxIgjVnplzkblwXq+6Z3f0TMI8U9/0M54HHUvDQNSL2P4tq001UI7geqJ6FMA
mbvEGkqleIkbHU2VCsdH2Qg4Vpa9FslSq918oUxmtSlhSFRw0EAWrK7H6SUQKcqku+xY4LKgIvcJ
OUxKkeFScDTmHQNoLHpBAj/m8k+3RtUQqFZ2b+fLg8+4iIHnJGonzbYWwtfhMrgOz+gJ8iU8jZQy
bb2em4fmOLli/W0ssurkdK9BKxQgR8+bAwYw9FNtBykAicbCTrhepJdoqz50OtrhRV/WJr7eu7az
wd9uSw0Q8OVl0EbKnhU35wdd0MgZJbpWWcK9hjXfK663fJRfStLB8JObpwa1rWOGgGqbhbDL+OUG
6Gy9qNSQGPlp/apAij6WInWTMDJJZI6rwyEFXMsIIbRjvgbFmNJ9hv8eb7FJKMVJZh9x72cgkTr+
jPZP0u3narMyiK0q9KiA+XuAaRtLQv10MOJMNouBqFVrcVbq61x+sEkeWFv4sNErK5TdUW0vm7b7
eI0IoXe5qn8gMgsIiXBJ9X54exx9ve4W2/PXeec8PA5O/JmfCDLaQ6SbJwa/ugS2ib6jmK++lIV0
OtHwP/vu6Sul8rgyxFUCDKHVOWyrN07/lUqBGEAYsLPPbMDtwe4xVciTinfJAfz2eB+M7hYotER+
VbsiijmbSp1mMiXRE5fJoDEcQf2YHSKpts6uTfPzpYJZeYZaAtK4gcQVz7DV8vjRtne8TCMpZ3fx
RAjg4msRfYj8t/A9Abroc1I/0vgXSzLzioLnJVzMHcSvVnlRqZjujFP+hOuD6nStBhfPazMm1h8W
lv7nXfndr6SMtAAA2Jds8ca/bbi9ZQdeLuPY/Mfrkyl/izbHn2eEk76rPYMaccSR9R5VP1o2w2F1
xpNVjdb1yRDph+JTMYWFO0yXpJzLcLt47gPjEgAFg0eGiAukZl7A7uXHAF1aO/JnJJPWLGtqw2HI
2PQlNdqqtxIH4bQUyxwiaS+LFw9rRcWAwrEnDPU+M9eW4SclhiGarh83dNGHSbenEZ/kz9UCUz4w
bmPSH0btxMvDBttkHAXhumsNOCEh8OiE5WMFcy7sqnHl+YPSX4ed1af5H+A0lfceD057zz6ZEn5k
kryEk72OkszozlrfhPXOx5q/eYOnIwz7znltd3NYBElHU6BhNxWId1cli1dhx+hGB2jUVNXQ6Wj3
TrWMS+6QuQ1PpttAdQnJFnIVmRFTzgdDJptVMmymp2EjAlLybIt49z+XT5e+dmJXjKDgL/YpQ+i2
DJjPcn4srg4UenbuASXe3RfEh0Ff0/hrsiVXZm2bo1nIvTtVHdbY/utKBX/IU1b5H8pDlng7Cxsx
zWoVNqYLXJsyx+uwp67SgJEDoMEx9Fzh4wA0djaqb6JfspRZRuL4yDgT30a8AHujkBdEYz+C6FWE
Fbo9um+FCkDUKTBNh1scQYwqLdlFU+kV0PpL62IbnOcsH/F/I0ZP8i7wudZH+fF+oSNbokxe5R0R
8D8nGxi1NFIoaSX65sFK+c69SwGnsFJQb6z+QOWzIOcLNTlje8mG+iH2ER7g+yqhHpsUzJJNQJ3v
zi7IVI42GFnU8prCxrV/qn/CLBLkKJFJytiT5bU2DA1BBlp8XwBY8TBA3pv1zpbl0Niy5dKRTf9k
b9jg2gKS++sivYYo1Qy+oXh6Ow+gTrKVb9ZBvFGk/nkqL/NcQFo2CHfYdJku/pMpG9tso4EMU1nS
e60X8YkG2Ef38IBiROOyjzojBHcYGCso1AUrXafQbaSDhlHfBoqrwYGKdT9UR3a8/tPW6GmrgY1/
F0stH3RfeUCjvQsExaEBvzH0SbQhXePmsFlbgcwabxazMSZZfbIU9Yfusch7ubuTNKCCOakHPeAo
LH1MVZZ2DPQaZ8MBZas0FdE662Fc9174Ju8fVWcu7KNdCplwuOO+MPnwi3uNEqGvme/hQzLXl2mJ
bYsUiwvBz85gcT5UXsfkxnNRcmlsjDItgUlZVSd1zbys45DTjohuRs7e/XPs0W50nrWgWxxFTbM8
JJJBlX0k43fnlr2Mh7mOKm06o16i0kXt4vfLaIQUuEoRQNtfgvpHbg0sav0zzDoaYnlB0PIgW6Hd
ZdHGxT02hYIc14oUuc98tf1Cjh5FR7d1XKuON7Td34zPFcMxpZVbahHO/vx5OX3gxHThErjlOlep
tEEgGJs42zCKtrx5QFcW0cwVWxSm5aLxe4hRw1KjpJ613VlpDKm8DKm+AKSpKaWR4jaiIZRON16A
uWIUO4pV9juLNfFkHizDlCqyemGzRHmitjQdy+LVJSGKE/zpJhENvSKKbvqhs21eGShVL9oPkRf+
utcBSGBfc5zdnjDylgsfoHodLXyx4k7yFbHQG7GsVBgoTVa+SODUE9c3eaAhP3PKJBY9XlZYMbuJ
q1184nC1CEcOr8kvu84qp1j0y5sSVToNPSiCs0xF8NGeXlXXhsmQocG31N+ibnPThyAyX5lj9uIL
7JIvSoFS85W9HExwifoNGhlixcanFhEq9uGSIZOWoXsGdea4mjBNv09VLHQ4/nkZKgZRIZu9164j
efHbCUj87bPzU2WBZzdxlnn2z2PaqcQ/4S39GkfPHQN9PzZi7IhpUNMzziqmnJhawemH2ncCx9O+
mOQpZbRAopBAtygiGGPdk0RwSaC6ytqd83asUJbd1mnROkJe/iUTOCYLlsToTYI5J9Axl8EX6qzT
Cg+49/+nv5yrKm0veDW7mp5zE/HLiNtjuZLx9sDXql3daJgQfms0dm45ga3xtW2SZhmzrCC2U1JD
e/POCiBOqCvlXblfvj/fokD/s9kFV5JcmDGyUW75pmNI1A5aYaYgbN0CBYaaRnin4YAaDZ396HA6
wjWPw1z34MSanZ0W4PWn9eXoMrwoAYmndQ7JvQ9W5v2hMK7jLO7l9s58p40hr9R1hLI5tQHV06hZ
/hDNp0emvKCETPlbyHi1P0/+snsFgOPPuzV2/AZmgL68ysFObW95wplJQfnXMPii/ic/Df7yeCiI
+VsbTn0REbb5WUCf/W+9JWw62RhiTSFH21JArJHBer2TNCzrToObLWg6Ehv/5+dZGX8uzFoPn6OT
6b7xqZ0q5FBtL2G4Rcdw/j2zzQ0d89aru1aztpRJgdTi3LvKmNCc2lUBkgRaEWEEDiXnR/ycgCi4
agTBHSRVH8QVupHBHlsK1wfP9cJKrreD57YtQfPF2FXzdmCyKs3jSHAZUuNocOojA7PFdTJq79zI
b5Iqlei3ceSEgJ2ZPJAW91dKWEwhgPP3cMnQekrYf04BuUoLprQY1npxpo4qcUwF3fTdWFbvTefE
VF+LCFbeC9KMBgTll9XCFSp2jx2Q4EiO2TlKFyjP1rj9McgCr1ibJANT2V04hVKmtN/6Nt+YbXZx
hCfIC8QB1nKfwcgn/BcuJ41hj++/DbVTFAWlwWC67jfYN8L88P/ziLA/UEStReITTml3KOKprUXg
LD+TJTHLx533cIMaFe5ZrN2ck8m28sI2BGQBd9w1PqgBzDo6kOimWc8RVBcKGFol1veR6YqcrI38
iTd7yP9cp5sG+9LIhpI/Jfr62JpyCBbPmvaW+SD6nar8EsWw4fd7iR7svOVnOR+yb8kEtAS/C0zB
wpEGc1BZCMuRtTRKzNVqnsAalrdCcF52FLa/4OysFcUjVWj+W+ZsL7dWjRve3it1dYW9JgIruem8
rqRJjNp0Iv33ZHxEI/U3QalWVXoXiQKKge6QTxQPLFiwKD+9iQYnVWo72rUo3sYzebdep+EnHz81
5pfWBD6Sg4lDmrycczoI7LlsvtEi8wuceduipH0hYONAexbkA/mFtB9ouhQ/2mEBcHiHqRoDt1fU
gfZa1/STCIl7MYlXt8Fr48M/d0cwXUoG9VeISr5Qh3s2Ro65mFvIr8FuIvRRmE3ceyeo7bcWDP+t
2O2tVCzkkkx1KOX/1zTgbAcyvZsQTdVeZ6KWSCbyiP4bIku9wmX0BbCt8u3VuZzM6I4Ygkpf1bGX
iRnUpnXHZNTYzWQgd/vcJ0K9sKrVXl1x5LSq1FgHYBV8eG+BJIFbx9vZxRNlJTDBcqmcHEuonJN8
IfbZiGKbxQQ3X+Vbni3hc5AYdUG25Ry7SuW+X0rhtkO9FJsibOKRtkLdm+rcNZEAWDC7DiiNeD0P
b12XFISi8RIPUAojlfbXUccV9ZIS1S9GEwv+z4d1wpMGDd06i/gM9k8keLydPPoE456+cpnMouy7
vxIIv3XdEhvirJKot+3fhe3jzqmrVmSDpiDhD47z/YfMGz5r47MKCIFnzuZRBBHqtPSsyIw5UjJj
udW3IOEc1Oe91uN5zcS99WXHWRvRKef4Js0MS5QjKlgsNOK8weIMnOoDY4WEnTTt4heNET6syox/
mSsz4CoeQgncqpuPdw9T3X4yfL3eAYW/o71hNBqnu0CNZr2qqSOoR3iPrr+Jp4qm0lfg+cI/I3KM
StYmc9pwPI6FazQAmyXCUy/grS7R94zQ4ktxQyo+jyo0x8T6ti4nj9cjf1EVP0wViZg1zRnafg7T
YcdfW4NVayUmbCnJBxNNk8vi/3Ad2f2SMW/CA98hcM9D7wdolC0cTQ4X33ye2xHGbpegGm3OKmHt
DVsrdp5ykHcP+62vLWMDV0wpZny0sm7ib2loDu23LTTVgDVJtSwI8L3jn0oFFR7/ozSqSZ67CyVB
N2ymbgevC3mDLR0RmBq7F1Y5BhsSm5xznhYY20jhRztwEcyWlPXeILNdFwUK8MMLjFVwlVLTayb3
s9H24Ab3x3ieqnoOjBHqe2lBYe92Fp03+KMjRzOseT5GjzPrSANLTMsyaR9F9kTMAZevlgB+gNKr
QSdwR1v0GnX6KdLOWqRviO6L+91jDvud3phsAnsxSp8ISILOtSajXMtPWQ0QkTAzaujfiV7RIwJQ
+bq515KINgvC2plG4c1WMXQfKi3QrGUlj41is3p3JL2+vjcwMk2j3jCK/d5ywwUaSppxf/VDpy73
wA9ed1TtKadNWchysE3pzDiZjX5Azb6JcYe+Oq1pwho1j5PCJrb9NjCquXL2alGgnInYhwQVnSpG
89RhUU0749TXw8x+28lxkWM9X5DPPAbDYgl3+vCz5tiwCX/KyDCFVaSVf/gGbAZXv11zxO9Nflsr
J3l1x5iw1FPxqEYtbvY4LkDZrPUFIlNAifXBJ7vpl214aycjT7dt/3wek+/yjcuy2IDLOOtCqJ6O
FJB2uOAyfnwhmo54bQf3dapHSJDhQsYaWVBKvfrRt3sdPsPUFp/h15ul8T3PdsMVM9k/V5VxmMmS
gMwdG+Z+knaN2Dq02gDjaS0m8cpFLMu4gbkFwoVL4OrrowaqWvuxT63Vhs//q5U+Qu8HyIXKlqr9
zIxCWqmF52g7Nr85xt6Zkv/VEZIxhyOx+9pj/pewxCyTiNnldflMga4lC2wot0RMWHCMYW2v2x7p
PjSR/YQEioL3xoivG2Mc+YxfTrwCXBEZFepexuOAJ6EPulpb7faBuJ+oskvhAvnxvFliNJMKrD6S
Llgjhyby8kBx4SS0hgjz2fuxs3FT4Sztt+92T7KdVv8xTBL/4Z0fbleYk+b4QOcOHoLsXIyd3Fg6
4WT9vIUFx7K8+PBkptDm61xLO9WdnJVp6QJo8y3wpRXuLhM0HkHTx6yoiJQEeehVpSj+bSQ24nT2
1MCZnuK1TfrddvKGeVUzkPIteRx4i+r/XRftchjRBmc0g8jO70eVMoFF/u7VL70xnJjeM6qTeTjj
TkbXp7DO05hZobOW97DXyEo93DJae6v8FVdhFOP9KJQNkwEdgk6/XqvXX9H+/a+eAXRv834CRCES
+N2v/dsgBliu557ZD7/Dj21gb2YIkQkoKwNATjR8HsDWRXbsq0S44e6YMjAlfK1C8Y5nZY7swkMV
7YfXeLbYSxkhLbA232JfLontgIetaRziQYJg6+apP5gVwj7NAdSETZSL/KCu3vlx5cpS/TPQDFWX
jd+jUP7i9a0P74aYEo7O6ejBYRP96j0do8fmrUWnMwYzfivCpJkKATNIe2WPg4qghnNqaAsDWiap
540/kfBxvxd3FPvorI0RZTPOxuOKupX+cmXxy/1YHetjyk12DS6KNdy7NuKcJeZVek2pmjANIDyQ
Y2KzKS2OUT6Svfog/2u2U5OXPeEwqwrg499BpyGCdXm97T4HQbRUNV4J4Z8cVJb10faEUcwjggST
Yy2xC14E4g7SPCzeMTX6ew4L5nf3sqH2539MPk7NASARMHaC79inA5qMplffcYkvCl4d9kZL8Svh
ajgaHl1ZCPHLllljNRHbfOoGuVEH3RD1dcg/G/+KNWYOIfEn8BX+1Igy2mc2M/a6Ktf8yJEA7tVh
PNsTQTvUBGkAf29NiMALDk0AqoBIrMjpawYe4PLRDEF/zDVYn9ailvEDPQkktweTj7fxrF10xY0d
jc3OgewjqOT2xNO1vh8awkKSAg9Xbn3EwqXzbxjFhVRzWQPVCKyIQp1yYgDBmdRW2qMkHK+eVFmD
yYoi+0Dshm9Stmms+/WLQYuSsAFAyi1I6eBYZp5A/7/cq2TmI6nN0Yi7kpfKrhyY4M8R825FKGJX
xVLisBfqgDFvrRoEE9/IJ+Hd359ZsMVz/gbxUCDq2FeADZs82eCT0BS+0xaiytOZjuTP7Wa3GbSv
i57SvDXCEzex5k1L5JB9cVJ8Knoqv/KhRIRRP2RAGfR7tpvv0UR2TR8OT1JwzdeIVwi55nVemH+5
ldXv3jNs/2ASP6OD/ntznhidSlttLOxEVJBpX13z9pUZCZUXPgfy2iWejkk1x822iojqR0ZoDaj9
fnrmlAr4pwsquzZVEe2GNLhzVwTsCE9zdslKph1ttt2tqz2yTAa47DokvmRdXLXoL1ixJ7r9X5BI
cSOUhxSnrNEvSjulcVePopTEL592uJgMVnDvpMOQ04Rp/9VRlIMDNUxJ+TM8nHQ9uX0bdTp89GPb
BPqwu5mP5REMrfIogaLbIniQSdWpKYJHwjOPo029zo4TntmCykllLKeBW1um6JSTiEz/7WGlxY5I
qJxeg849d+i305YNFbMr2v7RY0g1ZizFXdbTtMhd7AWeHsDu64R3rTJx+rb56XCnuixQqOp2A0Mu
W/AO3ndaK5UL2ZeUELmi1Eu0SUF9y1SO9CMjrrPhvYC6oiBPsf/V78yB7NkX+70UActsSWYEayHt
qJ5hsFYGs4DXbFocxPJcrLheuBRDd02XV3UKsEmoQ/yay4EpxTTtlFZL06vlQuN8IB0+9GjhteWT
sgDAvu6GBr+BicUVNph735M2zTcti2A/4GOgu3ldDZT2bRXwHelhyKhBnc9Ju2/qlz3xcc3ZCmSB
B/94l2yRrfvhwOGNyRBOoZnh570vB0rtRNJPSu1LexKnrjvbg+HqeajOC80bZn2e6zosQVCht3kH
DqhMRVoo92IWq7Y/eU8Z4nqzng7XZsoVDWDtRvZavpvPa2y8eSy2xl8L/OZeh6hwyifkEyIf53Yk
r6ci7S8ac46UXA5sRS/RjRvBpObgGjVZHtqmMyvnPBiRyRvRGtmVpKUoCmmZd0VaPgSERYTN16ah
kVXLTzgZTIG5BIpQDVQylHIIoZweoov6u7dbrWY9BxcmPLO7bv/Y7dHGN5OzxtHJ1mj/wotWjiyN
ZhY9af6+4iLd46j1mWid83WqpAvtRFkdgesXlVybwYBvaFqafodozMbJ9FHUwr07auZybwxdT2pq
Rw+Wcdhs3Bi5zeZDrCew4u2qr1xwbXGID9IGqGlrKHIe7bPNO0k3UVzM6dD7bOS/JBm3GZUSPC9m
OiCI1yjkCyVjuGnEv/qEFBTgJxhFXFJ5U9UwsDZaLalw8muRsfFvxwI1Sg9FVnM/z55bEqL5SjbV
U2SV/nft9+DvCD6/WgJFdpPd3JBVqrM20Ll7F41V0z+XrrhTAz0dAyfn5wOFTEoX0tIGW1YYz0ZE
TZMK4coyF8M/pjji305K+B9iquyXGPLo2wYMOsI2Z/rZsh+afJpQ+edcsNTNV0tqZ15RSp++OB7B
ejqPoOT8jsXlmIX5YlElSxW7ukLjTRGgzfBAjXybV88kLvBq6sdfBbwrtE/WBse/9af5gHEX+8Ug
nIpHQpkiIu8w7g2xIKRF06uZenZ/HtGS/kCO+mNw9j4kBkgp2ou3NXiL4s5JxnlhSYJcyB26xLeV
APpPSQN0zhAohuQt8LZW8pJEOd8NeS/Q4tiMWrjDprDcQHB9f2S6ElYAL2vAOe5ClvCGVHfuwAyO
Ri0WMoDTa9Jpd2ZsIhWH97HI77rqAlunjy2vLtbAoiNmgnFi5jfHdxr2hUFXXXvrG8Zfy3/8iHLR
SimOIB4MEFEc5Qnmq8nr51Q0rz0Xhgm4g2MnEgqz/0h7pV8D8hxeSU54W2Pz7zUn3dSUGoMEjnmu
w0jkaQ4U9FcuNv3lIui3Zu/bfqvcN63KeI/Sy7hZkb3LrQiNABei0xq2kREKO/pS6GV1gfUL3pmC
69YGxKZkfV56mew/KYzWsKbgmIHjXSifr1huOA9ayJSuOuwc8QNdeU1xmGgSwzrj/1dcVGinYV1s
IIkVG6dvzPGqDE3sOz5eg5Bjniwdqf7nxMHc2b8pnPIbMl8EgudjQbeSMULFnXjXGjfL+Y5FYFDg
+wx1DvGqDKaspyr0wu3ot4lfHBZBZPeEedScvjjlaVkX7IsPAT/AZithzculj7o6L7K025+eYUin
7vYHO3iZpqoqr/+G30f6bZJCCLv3hzFXmpOjcVZ6d8V/MYKl1NzJ2LwV4cWQ/NW0QhyiZGO9uhOZ
pKUV9UyDlW+7+sCWlAyn83WRSmF50j91cB4acQA8Z0V4JDu0b+9fUDAX0y3Z9PSL0UafVZY4U6YN
rIw8Orr0qRyjsVRwPasyPv/w0vhkzEU1idPNRJmX68AIHIr9LVsB7BWCluOWFkRJwIIHyzSg2X/F
oPn320//cz5q3v5uWw8RbRH8L/I4XbYKkaBgWbCm5OLUQQibDNfzrNviJSoWNIDaH9onrrTj2+6g
7hOX/+6kzYawGLv/FMAviP4ZwCkeJ7fq9mseNe65eOGXtD4g9UzA5q/eWe0sYudL9sa0vrXBm9dG
QWWsfOu+1lZnTLZu//GThqQS0CiSpuAp0Kif5NazotpGwBgEaiO1+P32Fk3ZmylbP8/fkD/T3JW7
Iu542n0C1ngLRcMN1JDAxZfCGurGkfvIpDMhwFuO3lPRakU6Y9gYN2QX9jQ1CW3bGxAJtzhN6vEi
yO0bD9gRNiaqCeVqSqGd3fxmav1N/LALv5SfJ0peK60ceZGYEZckvVwL2qq1EHhRnhscllwi6bgJ
HsWF1ex3WqzrIkYSQjt9VQjQdKrDXYzUyI+QttGGkXkLwsylELv5VZP2vUPqIZvFGDe2WmIIlxI4
kpd9WO6MFNAuzaE9z2bq01RFDHijr69tw/UkEM0XC5V69PgBBFob6ZUpElxESCdjBmuoWrbdhXoW
LJCd+0dqiIorYyLswV9mc0nFmZ6PINYoTrD5pXLChijEC/QYNvV4n1E2jRSlWNurqB7TLJy7mry3
PKfSvCo+DcIOqyc/22AYu48kRgVsd1e7+0Ca7Eb3OvlSLYWUoEk0UwOiRSUiZwcUtDjcLhrbiiVF
vrDgl3VVWbHWGyvny4k2kTcbplvuorNLJ5q5Edt4btRIMUwsyA5hygTBhMZWqF/Z1z3/dPwCUKov
1lVgURKKaxrBB8GQ2qGt9Mgw/2Fm1SvpN+yt1wmmAaRgRKe6c4UYD5j0qUdzNfNB3Tbk1+fneD5f
jgLH4jL1bOOu/5rtzYj3+73+73BUuOEKd1hycwvoCf1+gYEzgTZPmSsKgHn9mNJ7Cr0v06AqdMKz
2wE/5bLm26U3CzUZk/g0qwEhlQsbonFgU7PTLhv7X3JTOi14D+u9VXxUfbYeWfJPJHeJk+rc+1Dn
qSic1OGlL2rqZYHiiRefu+ILBUKfqhLpgkJNwd8aWv8xkSgMb9JlJptzG9TtGOIXrhzb9b9DFBDR
tM8/KbZCGaD5/vU9YL1ln82hyHxCTI2F3Fp4X0BQ0AyORR2g/0UxhPTfigSh9lMRKEeMfgqGqqhq
N5Le3eOtlqMQ9iG1oKYWdf8KntvnKBBz6Zm4VAqRE+kAmzWKuh7dRYKbd/lOlXcgrkZtz07cA5fv
aeQIWSj1WPIn4MNU8h05CQZ8HfaBgO66lZhVGcy7SfaX70qA3VQuXj49tMyC7G5QqhY7xIy0MWLk
hSA2lwxmCtIHs0mXX+VBBI3pqg/ubnHOjEugpYv4GjS0iKwgfmS8OI7c0ZbuV5Ghm20f2ND7Jaoh
oGXU6VbplMystPAGDMa2pi0Xa9ADm84HX2hlx4iA+V6/HThY+2assMSBM1ZPDNW0EWxTvOiQG5jq
7XPcPlVnVBSpbhVSrW+7LmiCoo+/kSa04kqDmDpu2ibPUxQYswTB/bm6AxGlCDjjmJBN0UiiULzb
Xt02rvIpVikvrbHl1PyOKYKXcdttqzH+GUSYZ3zNFfr6v1K/XtSt/2NQnl4X7Q8fe9s93+jBWg+a
TfGtuUOa+okDAUIsMCjMjcFkz7vxOl3q1bUus5RjKFBBGHMg26rHSLatj0QxvJI5tbTdujeZvsYG
6xMyUHxGUzRBlec36X0wZqXAzqRx5GOTPOlo5zzH9XudExiVJoDm5cxuQ+7SG6xlNHH7EHh5AfoE
1YiErUZleboCU55LkvOI2UEukgjScjmyKQOOEtxq0IXVnAze+1y9F48tgAcZKCrAsnar724Bf8AD
A//KXak15zeOIMlMluQiz3er0nBYGNIExHrtQB1YyufcNFoK9n+sp4swMc+vRHnwpGxjVkiYaDFV
nbZWJQVW/a9mb8YGjZY3sUiid+LtWIKXPfVhBNXVoD7C4GKokrNtwhS0sO49I328rDcPYOxk62lo
UgZiWI/jt8vIJxQu1lwjSgav5vNTGZBJXxZLu+eeRp1dVRPdjGVfT8OSaKen47+Cc79H4GJfYGdR
hGmSBCWJtLGlt15fQ7T1b/XFyfv1w4hdSWP3tPhZcuIqSfPAWNPxw5vnmWkYyYkFjwPuOBl0l+o6
+eWSVIjKWhfetuNnafeGjIBXnnzkCV6ju8XBhUamSkMbfiUwtpE9R+b8qfVIcg1/Okema+CoOLBI
CK7EYmzRKxhsAtPE8TCAnKbZuyQbLd1S9hlF+CJzEyLIEmkXk1PFqENOKDihoOGaM0ng1bXe5Tbg
kskGcICRE/oZvXl709rzpmbwW2p+y35EOV5n++BiSEtGNGox/xyav9ogkxXqpPZI/wgkL3sSaFwG
J5420d/1e5zRXmc0tKFOjekTxPRg5pQTDktF7362vcqp1lKnWND3UwMR2dvH03YSpYzlF7fQMwz6
jcc2CzYk6bI8aCBV3vcQLbZ5eYrQFpRx+WbuJPQIf/5sU31oq9aFvQro5MokXzjyuR6YrDtHXhVi
gWh/JG7qr/VfKUFeM6OrTORLG9/yMLo4HC4VQNHhw8t/B3RtSCiX7nnj115tqUVZl511w/XuxrWq
+EByl6xmbmFpVORhw7gh3hmw3FHkkIKovrnAk8iefZNXOjuTR3Hq+e/GGA9mYk/38ybJrs/gdZXb
L/O2CAxv2NRjCB20RyCrZhqwYPz49hqQSBrJ9j/wfwmOApnbaI61kDQxNUixtJ83qH3h9oaHh4Wm
0SsF2ibXmvMmmstn2GY0AKIuojEvbcuwQFxOZSbfiKuXtx1VppcTwqdpYm197j9KiAd7dyoXaF/+
QMLPPxIzFt/U1hV6cvtVLzv9yW26y6rkw1DzfLVegg4adVV0ksEbVt5HVYCVxXCU2mO8K08h2V0L
M1Tj91jcJeSGr86lGi4GuZplTrERrAsSY2J9/cpJ15vmlYQRdFBTk8Kp7NWQTgH5zEUOflpgVDGi
KF55MU53TdLaVp523lu5axX89gsKGs2s/QA376PhK46Sf2/1FeCG/iejRXMXB/ZHvwQMtElxAecA
Fv4Xm3W/P0Uph4Me1z9UoJ/CgoqXkNrI6NeHxiqZwQcThEtQ+dxa4AYx/AsPXQibvX8noglPdXUs
5EZqbnc5fJyyMvS9i81TkTp6FkDx3Gf3h/MNI13PWgdXZQjB9n5XlYOn7O0EhyrcKlRK9KPJ2s2W
EdpRQxLpzj8q5k4yh26cnnxHgqomkCpZc3tCFWzhkT1q3EnA1mGKqUMEoIt1mSHJ1yyI3O56cEuD
UkZoutwwcJRNVMKBf8O5Dsuy4oQJ2T08tayvrX9CKgqGO+kI36FB6iCO3eGioeYYdIyEk+HRSV6h
xoud29jog4tu1o86Km50ZxeEPcHU2ynaq1tPpoToUiD7mzNjPyIGTdSUewqZHyP7l+1kVmKXM7XL
SihLvlB6CyarThLxxS7NMWNnkbzFYYlRoaRzOzAQ6Ypca4BRP7W6Z+KYdyEf7RVb5miXJGXgT6S7
Mj25ucFkcAQV5dF49o2BZupHRUGZdCR1gCEKZB0RauFmZc2sYZP6nTWX1fgsNfI0IKFscW1qOsMX
lYgUdurIMTYHWw/E8KXvfV/Kx6YKjMidjGUYOPLQ4qOTJ5ezC6xREUObra2ZTz9JayGelCk+hUhj
XSv75k6+E9lGGq20D/x1621ZKSjR0dyKdtnKsuow56Xd2cubRCuDMCVKHzu9GJ7W/f1YB4T2jrp7
wXQF5ieOQOJU52vJWnLGeY94NAXBhjc8UmV1bNC6BFpYItjBurJ5kmrINI7ZnJY/uhmKc5Emt53U
8I1GD2HSBSCgcGtSoCAOJ2WjioltpU0u7wmpEcFRZIe/B32d7ZAsfpGqOS3g6Yv1IXZV8ClzSMV9
waqexu/lNdRSikBxdUG8YHx0i7oEpmKKeIqn/i4684MTsnv8IH0duB1dRUoNAkDKP9aGrU+8fEkN
UlZ3kxhWDTEISpQqQHTbGMOmJb8yPuTu9qKcMwYMEpeAartmIPwt8Ppp4Sbr+RcgxqyvFuP/7JCK
ncxbPkC3bJYv56qM2lAi+ihTD3QPTDd0BafYR4Itw3OAGvEzUcW76liHL+rqzohIPiErNAAvFN2g
vP6/TU65ubxxmKzLCVbTNeozYa5hnWCQuauNYsSzTojs+THeDguJc+9XlmzAPJe7HmolF3s7GL3e
rg+g6p0KGefgf8ippHSrBz3KL2+wRuGfXw3Fdg5TXJ+RS/D8B0UNkGSLlv1c+LWvKu3WKVnyDS4C
tTyG5VknxIeH3xoP8WNOV0D9GK6XvP6vMSyfKqzfkGaN8Nlv8AmIJZFk6ru4rOtp8tBwoB6lrT4d
kaVSpN60735BMiMfhF3kHqMhW+VXth8aJqG7w5QAdX/w2CIU8TmJScWkKaqIwZQpxx8p6chKl09t
DbuBxhb5yoW81HY9K/6ATI/JfFszlyMjvHBe5UEcWgSkv7QZJVcAhBwgUJuEVQue8sLIbvqpcSK7
1XkPhsNhk5rEnv6H8p7m4+bHMKfmWOOClZkr7dDvTGlBiDcJ2+MLUNjAHi7u2uZYIzVHC1otnb7K
rg8YwaNu3D9GxZos2SPAd1iOtrJ2VrDVdBQfSYUHTe1mWYMbFBtuitqOPILqmH65EOI4tXI1RHeB
21Ryho0zc4xUNECOISAm5xZu4OZNBBtmyvHMPu19zqeHxSoVURwf8l9ugoUjeBTQksKYFV4IzR6X
9b5mc1/7WprjMbZwSQrQ7Tt4kemjTQuLxM2A1gi+7zeoTfcgc74mK1gDWLRXiFHC3sHANsohmLjt
MSkb7f551B3dO2GRLSK6lqRcb9UEwWXkATLYSP9ayOkoY1VKzNZ/6dgnYAuL2BtN+TTRT04i/SkU
S9Rj6P+lnYiGSp2+rPNcYikinmgIoCeCRrmFfvquCgU/uDkKHCsOuBClhvndxs8jRMB3QPxYJHCH
38DzCsV8tlFG5Kn9dSvFaBgtTcwfT2FaNuLI42yHvdAVcXio9KGdmh6kVdZsjl3QSUml4jAmDpSr
SOjAmAQ2AWg31H51mHY87odmpv0bLMhiFFSPBWxqjgH3gLOa3ZBabGY3pdPE48SmY2q5lJb5Yx8R
bV0ZT1/2A57QnRDs/x58Bykpnd1P2N6FVmvpcwdrs6+XWslgYS778QEa0jlqbsifQu1XEbkeAuOT
N1cxdLihbkn//ZYQjhL4HSmB0z4iU8mjEYnpYksiLYhoWkXI/V1izLWBz1bqCfBYxIl5q57tcS37
ETmE6U2K1T7EciKb2Upauj7LeS/mRakJjwDh7AItAyokRSvpjoFCc3moR5b//wXynnrYD4R7Fn4/
Td66DoMZt8ry8zmboG+kMoUYhs7kMEoiBNz8t1FYF+QaSCkRSLQ7LbXtdvkeQ95uc0qyF4TpHZTW
08GZt7g/3b0FILUOfF5jO9KKHyMATsH8/qXtSWxcVWi4LKDgfZJU6rzuKCsLBaFBCTMHI1YKzAf5
gDJ7tHiACVw3JOkdWHNXa4JxSwcL9vnnx73gU/VP+hzrVgr7ANGjXp9lBnpj0JnMDWgybBMm2A82
wuGbX/i4Z2RPCoe7uScQKv7GfEfoTGt1p+TPwvOHrQZRMm2cEtKaXtbLfYKuOZ1Oj8VYlcmeDOm8
n3GdD8AL0G+8frpyQv1G6Qi079c7ax353J9topvqtQ9Q43NoLZ3hCw58FwahDFeKGs8nHopmVAVE
76pL5kF180YKT5tOorvCw/BO1QU4iGXVsLLt9leRS8vp0/DyrBsPlzGfTMBEPSFH9j3GVQzJDel3
lS+EC5XpiHLcqb4qLrq75va2LBRqwSGQCJdXaZ8AeZMl+eZCplfvUOD3yiSyrh0muuYkwUsbamu+
Kgpafu5js7JWz4FU0xjVBy617bzRhdcqGofzZxfURKj/5IxMz2NnnAOIhNPhFhjH4dxy00swg9km
XDGMbwcuMwF1WUeKGGvKEchO66dYa6JAbfuLxQSkhoQvcSam8lBWnyOEfw7Bse3JSBouzYUQ5nJi
zRNZK82liA4cHYXJwmgqI41UHFEml0uqeuxCvxrynU2+K0IDRTzrAl3yeii0HCFi2303AM9G27tl
otbAoaHgPTH9d6zIkc7GkLEKBlYOsPv4hc4aMFHlwQeCjDKJIyKaORLKIVezY6oQR0jxHc+ZUbsN
WZDkxehoMej7/dKTkid4sZt6Q/9WNOdsJQgiPMH5qFqZ1E1WJTV2h/sGxsRWL7AgC/6ks5uzK2SL
3v9QIyoz4Sed8FGAeuivI6NOBVIhcXfLZjNFkBaMXKhWIdFFNUZhg6VBlJx2RZ6jjd6BOc0uingi
9WZVyRXCajVir7SNk37icbfbMzualMh85v1inAlIcmAr8hetHVQiVv75ycIT+pKsBO6uo8G9kOh6
kgvQJsz5jfJOL+s7AXge0GnrtGT2CNHC52rd0QoAwUDZ9EU19iyQ8pmLwQXHLEnvO73mrHMTPAxv
XoRmu4qa+JQNARipDewxeeSs+lgcvGLLZBYF2MmXokO7v6NC1+DOnIv2bVGy6QIHVBbcnaiILD6k
G54vXYAM6ktOaRR6Q2s4xPe50PzZ7U3DON9Wf9ZUb7s3z4OUz2f5MQfVtToALl/25PAvx9gDXz4r
xhOtsfa44qJedviCyqGk6QOZnEK599ypjL3owBuPhe4h11BeHq3aV6UumVDdwAMH2o18eJg7i8I4
hhXxxxrLgw/G6aAN7qfbwiRmldRJjIwJCBLaZLDkW1yBnZkNwJ04er6OhICikDey1xEJf6QLVYJX
kGc6TRvJsflfb6Ua0L1SIk/3LkXEG6sCBCE9s09/eHCQCtinU/9ybFC+mPzmVWMQ3Wvq9k1IzM59
h0gEeIqmU9XN2DuEogapDzmq22zGZ26pwiglwK8k+unzyi8MjORaGtBYI2N3IGGDUwBzyeLaMdW5
BQ4i8tqVAK/ecq5F8xV1yz8R9tIOqn9SxUVrVipvfIOVz8+ppaCwJcz72dlTt1Ak2b1dxnzUIpsj
Gjz73b2KIK3YVh0FqNZxUV/gDciEjPSngZ2aNlDhvgD6QEll8ax8WWhSixwaduCHx6jd2XyexPrV
iU/xo7rl/hBNA1n+IiuwQreaumEUUgrb1W7h1KHnu+Y08+07V43lrtz6Pzb6Ml1J/wcXS9AAdRGg
1CRn/FmRuHV+Wh/3z4HsNJ18Kb8P8A6erOLUfdi6LEsxWwkp+Dr2geRQLXWMNILtYRQU1OobbS54
8Gi5e3kkrPlQXTPCB339rGrPL8WYY/PEBNi0FyuoBSRvoZKEXXIDkSH9vsTw88YD62SZ2eJYEpP4
ey+YjvIyW5KwN/qkBrZAeFUmyWI16af4pfX2hyFgEhf0PSvq3un1yyyN+2JvlxzvepXxA/UfOPu5
oKXyJGF5lcacjIGOOJZtWaS6cY6mSWdZjY/ITe4f4kmtioEPkPLtmm5qMuDFqJ02dcmc+CpwXazm
OABZDNkU2cLOu/0mQ2ehRrZA7TnOBBqD4W05cKEk4ZF3FVVqE43W5XZqZkLmfnKg4HfJwy5zr5kO
k7G3TzSIp3RT6XqMN6MCBwz824vQDYP3EhzELdkOHQ3wg46nSMoJb35PHwUcTabz+06JpPC/kdE2
3QloQIVyIjr5F1h2oUG9dErxWawwaj7TczheOvgCi3E27YXzFI1scFHpE2PsPddPiDoBbUgNKjGJ
egHQZXYjKaf120wm1EL9NLS0VGEfWGYeTP3JQT/dwefZrSAGRT7bWXWFjDqQK3q77WmuVMOIPwC/
rFoReREibufmR/k2H/3dWzpQX0Dua17F1gzRtIKy5ntV9Vs+WEPjBlKYSvXt6G3tfZwGVZX3p3fK
sYmfSMilWIZMqNXBciP3PFZ1puDiz/xmY5TwONUKr970YBAD/90Z9prvJBywidMETiGylLT1Grl6
D1gz9dQ0jIsSDuscad59w7v2zJhU52Ux8nx2GUFsgnHe2+rZ8R0CZ2elqpLxLDi+8X1meV2/QjRR
QwE96LutIpa0lQ/aYKmliIf8v20TXcu3McJwWee5bTAxJfqLeta/VIAP+NjE/pR+ChCjHEuyz7bL
VjGYIDQEhziP1gAsxefZ9O1Sr6dViN3drtW5n74KjOFrMrw3Hq9Cx8AQmjQHvcaKe0cY2D0Xh0Ca
3vIHxqH3YkAaB8hLsz3DEf78pCbppqbNdipr3BuuQfDdutb90J6QxvNYDJf8kmxfEi+XQSfMYOyk
YWvy0MRf4PMekxFhHX9ZV+IpCYc9mXcKjY98tNP+JiC86kM5VyBLbXqfX9GoGEPR7uJVTUmKvzI4
xyJqBgDfn+41bpfkxcJDjpfxY6Ua1N4YEUoaCtvhbLoL8bAamKMQ2+yzGUNJ8Gt+5Vncr3i/rDdX
U6fxRyYH00vWXHfaUJ8jRyOwsmaSVZElZm+7IVA/DtW6pUG0CkY9N9DctP+f6CQpcaQ/CF6v7glO
3bpc7/0+gNQs++EgTXDoW13kCodcp5TO4/TrjNX1kqiDL9hta3KMSQwxGQDr40Kya8iX+3A91znv
dl/s/0Z5e0+WrCOnTk49wTXjdI7k1m+FQRqJwWYQxIm4j3MFslHtqzo5V5u6bLsOVw74eTuVdBXS
TAMnJijmjac9EQ4qAkl8Ajbvk+rtbeUwoK58DhgJKJYDP0XjjbdU9YQ0BUncjY0yAzUjRt9C5djR
uFEMdOfhHSW8gUKcEEMMLgD0T8VEMsHGwoahDV85rY/k40VPi4fLfVC5GsVZxyUo/eqV06PBdiBW
FHcGt+7D4udQCaVjcohwjsLe87iAUVJaOdVHynU38bQudyiUB+3Q44JCKjUVMtuWFdVBu/bmMap2
5CxWtEGUdDqKOibJAEx/dh24CkgDC7Fv022BiAFD5nOLFHGGz5rGBzjZGwL2MucY9AwstMY8bAa1
SrBTpKlheIOeERlzKLoL/pZtx1i7R0MTGom68oHtlQEUoZ6PvxT397X6/3nosxjxC3UuG+2Hh+3n
RPLl6TnAFLGOB8Cau1zCSyRSIhsJRtdiiHQOYqv+5+syjUS1r30HXmWgAXLUzylhLxJIzl6lNkQ2
gyeHLGmrRqAFQT3BGlcspNproCcFncQs6ZjnRDY1Cw1kO+FEV4B/jYB0NrVEbV0aUtnLqp4SLCfn
hHkQ/e0ugUTj7achYKdOIMs4dbhr1ueCISY3nnUv7q/2u7cJ5iaaiWSldarh54B/HpGwCg6xo9qc
ZbEb1xrF1q8O+zqreFt2Og6um3nY6wqE97iVnyBFSXeCDM+Bi559JB8CNqawcqGih2owOuWJWcWL
enm759ghVx4EJSCJlSDufDUd0U92QLFRiOdl40KDPk4IeO1xNoaO2KwXBIY9w69r7ZVasHoVpx7R
0gLuAT4njtR5g2qI5ARxwMflv6Nh/3FDz3v2Frvdss3LCmTMNUeYmGIrakMFeQmpnLf2HBdO8MZq
ffREepB9nrmvED95OQWhBP0rfdHeakpHMoD9EI1gIcA9IOqoMUU5TtaZIXSuHyPQSey7JmR29Pnu
He1XO6tlOeNCKxv2xHTJLFUmIL5bB844V0TxZMNrbDO5Yj7LLiCKo36R09MZHVvyLYwhVW9r+U2C
UP+/NsVB/wdxA4GerjVbXUTpkT1Tk9JwKQZenLJv7i3L/DGGftkIkW7m99ZrjyO5sWcPsgcoeMhb
ZCJNB8LavwEqz6/3j9igCJzdJlQsQtDf074CXiT+eTcf+AVMKK4L49EI1HNdLW6yybEvx3m0LbFZ
GiDnLsDR9L4bfaJlzBhmrYDvvuNOH9rhfO/4CvzSCGWDZf+WI2CmO9LjhKDHjJ1EjWrqmf68UuU8
GcLvDHDFAFtPFBIGQ3F/F4381clGnRyh2q/mJSoXOx3RS15dChpG63cuwDCtD+frZ5Wab77Z+2S5
eMAioO0TvTqGh+SgHwYpfwBheDcJi1IxborwNTvdH+iHKOR45itRJrl/s7BzBiS0l7BNxCqjTEeq
aXG2lOrM1g6aG9KsOTJ6lEzfAHlllhLOjCMUIiExPEUGQotjTu0ce91lWqpAf6U0AkrBaFrIDiG5
v4WOlpU84mK+gkcuhi4l479k1GiSCNHGAfgdx6BCatwc2iS99nwzGyyLnHpdCR/8h8wxWiFh7HfK
p6tuCpdIbMWd20xc9OLFjcbvSIhAxT3WP+wCPM7icjPcAUqj7NA9Mx2eQMht/ReXmfvaXZn30Bhh
YPUvfWZ9wqj9/8jugxBJvo4RHAEYuBDIKEtzV6DwME3G9j89pm1LDsODV9T3pku1UvFS00d1C85z
mnKWG9XYt/ZWWHXXle1T9kMRRPHw04MzFqGc6zSN56oPGf/9AUlKC7Uo1Bmp2JiXzPbiozXz5ANM
aZ2mDUChxPVK297mz+JJu2PngAaYNkpyo08dGPqVRaZYZBuSvYCm+c9tMjtrdaApzXr6LvsFJqHl
f15tqAm2/3Cen6CEC6MAxmcrZXISeGGWPcGxoY2bwo/JiVJeXVSiBS2o69TpOTFX7elY3Z5ASe6x
8Rl/21kDAlSg0Vb/nEDALaapj66geKOHOl732979/uA/Mf6yd93S0AS9UAjKMdgwOsvGL23GHWxn
y/s0QUR8YTi06a1PpReKK5d4HSY/PggR1/4dOwwqXpjEcOaDQGwJefr0qZBVyK7r3mOTBpCX+Bhs
gLLzmnLpebGu+sIyH00HoQdks9TGqxk5dMeWB5k03pG63ndjkfMMHcQbt70W52zQzXAznxtojULM
D+K/pR7o5Ya4z98vl0zH7CvTRwO1vvCmsGEEYztpX+XID60ENfukF5vbOmR07TYXndgfkH6nsMOy
aBNdzX13ZODu8Yhwp2QobbUYcyGh7ZBOqjCRJanhLvbNqef2g84u0mNtEf3331aakzmXZtIjF7qh
Me/VeRItmZP+s8oioyX6u86R8EwUEB7fNZjSbFIid5zArddazc2XW0k5H2ti0sTBzmJw//Bdx/l+
z/nCeAofbm/TlEf3zU6K4kR0RIpok9oTFietfgA/Cxqmgn8t8yPLVNf23K39a3x9SadUeiPYKu7z
4ZBtwOSNA/vYYBGBWbLXlR5MNqanG7B9etOiR0TiKy4NYNVJ0AlU6qJuLGcNfS4qNzBtHgNreZG0
el2p55111v64xs7M3Ka/jYKKjXRg7xrZxtd6Z/BabZ34s4IAX8U32ka7r8SBSHFZyktxJGvmUezj
J5hwWjxes+f5aYJBvz+ShW7gOaLB/QFcaF0T1Zb/SFwaxmDJ12JGJSyGSXQoKFYjVG3ouUce4ekU
K/1ZWeyE++WcZ4UMmxYGU8o6uYT2FH0lc0OiDZPlmHV45lIdcYZbnZJjQK9wbF3DoWQQd2cRvmbm
Yd1D4iCgsLGFXQFQz4QpvHnJDUUeYPXiEu45ALc6AenjRpTImQ3Le7ErsONcmN5JPcB6j4rOzDLR
LOvtciXuCUnW9L7Uy829uY9gDYrkEvkjvIedklC/pvgkErcIfs+0aaH5+koDXSntt/9A4j4oV3ci
2XzsVq5novDrQg93ceUTM5H1fdyysynqj47zCP843c3HOq7Q+Eu+sAiWGA0n7jcnbiY+/O5LkEFK
XS4IKPjfqvPS3L5+8GdKtTS51qf6VJ/YJbl3RQ8JnMAzSNwY7L4OIaQTHJJ2QR4puaLp+3rtxOAO
Vn+dKOzpy6SC2/VyS5zFtD6XVu6+bPBePiJPVlLNeCLS09PIUGgN8KvH5HiD7xqSAon4SMCMWlOr
si7ABk6JzJ0pF1dw7cdcBeIkXvEs1fJm1MtqDMEHkNNEaAPHq/CXjZWeRHqUGNSlPpxwQcp08Kqp
eEvzT4bRjg0olaU7uu5nAu1vhP4ZL9M9QKLQnuvnHC2cbsHKzPHo2PzwSzKlsFWASAdMxOU5e4v1
fObN0KzpfRmUqRyNpNgjrYWrE8re9+jVZXUw1eINd93vCByWK4Jtz5R9AJAANKXWcZ6/UNn+aUZY
x7eY1lycsW8vw+7m/7Nq4w5h+mDiIpIDgal6D5SfXVowWyHFxaY9Ly5aeoDfeQGW/2hYqEE2jKsC
T9LsZZQ/Pl/qqs0VXC8u+vGdC7+IMHP5x37108Z4Z6n6wx9hLDHqCO7JR/AB1M8g3YUdj9F4z0TZ
GzxqXfSGqEPS9+wKxCrUwqpvnFl8/3HnaDOG9TxzFO54/k8Xeue600VO2PYy51wQcpOadJ3nfJJg
er7BP4WNTJIe+wxJjZ0OJiOIk2yAsW5G2xyCRcqLZJiYsNVgtC6mGFlyGibMbwy4Z4A6EiA7nNlr
CbdW1X7pCGYWntZn1cK+w+eagYrDiZowrcd8BuzM05c1a8oT6yJM4ji3ksLRf6blw3zOxD0CrXfi
KPJPTAdDrbFFfuwTpKsxyPW7iiRJyrYqNQfjzGGcqmOrMW8Nibwcyt3ULmC+aOrkNcb1RLSUIdb5
8kkKou5ioOE6VwmXRLDnJSSJR6puytlY0Wle+b24VHZC08uN+HqT3QFynSBpphFoIdRFFigCvGz3
//M4J/0PWWYSAgPG65/TSItEus7ePhkXst+wdoZDGsG9+eHe29z6zF08KjRIPrfdvSH3MkX1XoCK
c/vmkBru/CRzLvCJqbzLQHLxb8SIUHp9BUbh28kiS9PiO6yYM3CXfnLSh9+GAJrUTTVQKIHpm1wJ
BfgJawtoFjTIuvLY61RmIfPKAJbS9xCpmTgeNAahkP+CuPCwCSM1L4wUUUSeLCUuCpacfH8/0gEL
pWPoPV+gSuap1sj0rWrhId032/YxHJ2qnYezwB+i+GaU3sv3seSTAr5U93kUMbwgl50FCIhmqEnH
407n2fseyWdpOcNf/pbRUysrI0rBocJDZoCt35ZNEVsMDBLu7biBBjU10Xi7ryw4ZYDuatvO/zfq
8QzLzP7PwfJXF/VW82BFv7XN28A1vQ4qPIyNVHXTf3ELQfOy/TveROoBwbwQAMb1MNbvY/Iy5MBO
eKmFYzaXGvCsxXyEvNRNwyMcpptU0KtRn4dmZhd4Y8iGPfGJGdolYgI1RrWMum/B8ZFvxRVQuTy/
XnzQG+8BWnT8k+dmbzEFGZbsBQ/6wCuSM0Fiu3AGPIXy2B6OY8EuRxvl3QnPbVogF8NJB6lo3Pnx
nwSfUMaOxbXWHOYNFEkP66NIgw01AGSGaECN90mRj6e7cNVlpWI3F1PcVkZzyee5sn8WKm7lFpsD
zZUnC5TiSHSiixvUxzMLX8HlhKQVw5tWQl6VlIgIo4r/xk4kSJKMNmPmtLbRRfchoMSH0T8z1cO5
QmhuQ+2RmdtXx7KoL9W82znctoBUYMxY5RfTc1sm8fRBeASOksUczfWvKCJPr3D9SxYF6ctpx9eN
MdVU5WHF36NhEcJc5PDl3h+PDK7UhhBb6wBtWTb7WGXB6FPkW+0DdosTnczMfSsZXG+pF2nUl8vi
CYlY5Ouo0/MongNAhMHmmh13MFWkCk5P/h7pnoWRekHpumAWRp/6mtgiiAu9Lo1npsmmnrWX41mo
1Ca3w93LxXKfibp1i86V0kVSdtp7E6zXYxp3PHx/fWVOGfnM8159UUsRce/iFXzILcs7P2bCjVY0
hbIGfPzneX20grVVem0xf7N+6PiQ0vjnHV6Uo65KnO2gWi6gh1wK6WkQ1iqUk1Mdk26LotF21ijn
4RNxm7iztH1Gk83NmOjnBExELhiPSsEu/mEPtsvY3rBlCr/uhsI9Qt68Hg4zAe7AlGhCO70PGs/O
oArdhb/kRzRrwXZA5X9gjFcgmPc9CG8dLvvO3iiUgNCFrkcsi2wybDiNOB4uYDMTH2twTQ/JvWs9
TtEhI3aJSg5wtS12j1DcdSQGOfuzicKS3qM8CEZe+o1zpC5pSjgZUJNzYd1XAJTUhmsYXFHGs2Mc
MyaOLbb0c2o7A6r9TmHS8FqEW+pXoqA6bL/pPsH6950sfe59EmN5dETgY3Nyi8asOuvoIB2kzzhs
c4TmaAU9sPIwAqr28/jvrHs+p7ZPBpQpfnI5JSOfsPGOmf0sd94kJPRExSVJhr5LovcvDoSlEmEL
5V0I0J8QxFAiuoPKFp5U851p23jjQY4Lj9X+FsToB2A4FK0TXUKdXZorNsKCXLgT5AkIkmh9lSbn
WPxWwtyrzx28KU39MD9IU77TCMuyEwWlJeTU1884A8EifNwsQigvolOhNHphO1+29hjcsQDBZz7d
1Qx9wgVuPWMw18X3RoH1QcU5XB36JZI2s+zqpAnwrLCeFGLJ7of5UFP0NhQdekC1FtE+9jj5Xb0c
5G0Xb8aK0R9/pXKx1H1dg2WBDtSfy3RjF49bN91XWoYOFA8jS4gubcIcMNdBwNd4221MgxElGrDy
8x0FN8H1cPeBz0t6GXNT02Gr3WTqMX81IixDbJoSI+JEB+uvsNAGdNWZsI2iN30mKPh6YTzeqhO7
9UdGQvpPLUNX2L04BN3nN+Tf2INnoVQBtFroi9UxnW0zcMvdxCsu2sYhauJP2QoW6Ltx+Di0O2fJ
XSSKbhHtnKUUJncettgVfx6+ee3hJy9ErhHqRBU+6RymdkM2491j8ZiQ7ryiQ6V6DhCg3Emr1D4C
36q76TbJatk5hnOtAnaaAndHRLjNZaCxTEWv2i7hV3xhnOvCB6NtOh462bFD5R0AvmQAvpxaQNYo
bJ1umNVVO7K+w0baYhZVbwZ+Bk4uKgQsmUzwD+jGFRYQwmOMleB/9WZKXCyUJLRG1MW9loMxTUwg
cN0kaqm9DTJC6DjDj/BNByCDiKKnL3KUdAwr0DrfV64mU0fgaINaVO+5JoWoooAIa9sofsl5xXze
ZilfCNRMVqkngTdshtRnQYV0BPHCGCzwhvl+LT38nsRSJMlJu3G0e4j5q9nCILkyOuHtl5Zh/aLW
KXMRCTOqcYEPbOPZGphFYkji0jxhGItk27812UosZJK5RsB/XM7p1iwLPBd8zDX3wCjesoNwzl2U
YkSskBQsl38dZYtzvlzSTKz71qpYC6hWUlA2BIwL78p9P/cQ0pHBzTi35SXkA6FpBtVSA2rth/+b
w3Pkg2nkM3M3cJNEGwSXwvwRc9A4JN1lxwTVveuiLNqosW6pi0D0vFhC18QkrwW61rTowDd8IBEX
mFti385+Zc5Ws+kV8zG76wMoCLP9MEjMecdoidEtSH+e0Nkkc29wEiX0eEQc7ZCNOKz1wjfBhoAq
fitNFQ5bd9rWXLJtXiGVb2pYtZXvdV0Nt1CuC59OMsBX3H/GC3+ZfAyIr7aFLiPkFf61cO1G0bkm
sp/PQlhRlOF3kvIOrI+4rrEzZAcn4L0AfOGKgo0P6dGF8KhFTYZ6KKPDnLPBFfFMTA4B1YOVwOUV
IHx5mr++hZd9NteeOSX92mc9ySI7+mnEDUPo+mq6jdQXauYVspDdplFQQyKMzB3j2eDtvbnOy2ad
K61lgBWjJAJQUjNSpGcuT/YRvyvMdZ6rV8otGtCOK3kbXT9WgDB9gxdjgNXSulLTjdnSh/g8ea5O
k4U9GC10ay5JYlv3HBZgTo5uyMoWQjSAOJ2qwoK0dJtg/v6nFhmK+ilKn9Rwav9g103gwbVsgeAq
MwvIXCNW3lcFHGxGN1ViO+j6V7VuVDVmiGXSt8Jf+UzUsfnov7qOQawj3DPTgbA4XYKirzsIh67U
ICoVB1jQFLLD0qqnsS2M6nO4nRmNyEoCs2xZtz9vLGDF+GeHB57OSCzN4VJz0r5apAU/GylN3KqU
xD0lIu3P27dpTtNOSe3VYsiRrsEsI5Vtc7DoRFrQ/LxnaDAufgQFOxFkd1iqJmGjPwU+LIctgVDR
mEzJAQpscBBG1P1kbGf9VjnNNvJlfsgZPzLuuah7A9WnDtnIQDihrSd3Jz7Os1ES8+NG9/b39Cwh
T/8YRqrKj5e9yt41+oEh/vjTPPhv+RkEx1X7vulGQm7boA2W8RBi95zZhZ6iyPqZL9qYzwqg0NS4
fzNi+j2FsMmx+Jo7t/htzVWr2hIILUwBg37vwuh4PEbF2HSnj/bzmjXNhm4mEwLjlbKpPVn6hkMQ
Jz1SYabYuCRU+Ncphl36csI+FNUPET7SC2ilb9J7OzMYYhFWbl2mpkLtkgfc/LqHEtQkvhdNpWCG
sXrLQm1EsYz0qwpLGXZ6pNZme0nwF+sf2C9+hKIC2VxaZslBPRwDQkni8fKhI49909UfRWhTxcmF
iuJNQLALo6ZnHUzNRyOL8uc1yF9tQO9/oSbI1iqfcvn9pqjGGnbuGuB3KMfWIaPVCBwnIJeKZvmR
riQcoQZyIffilvyNnpopsuFh2g3k0Z8IcFkj9Xa8GixocAYmhf1nQ4Kz1BVq3YzppoxYm4F6G4IF
t+rfVZSXn/x6GbIR0SiAyRzYLnNTQoZ9YUiR+/XlQ21lIG3XGKojJ2cGWAqdSDEWMyngzWHapjor
S0r5cZ966ImP0CcTyH4JJJduA/f3qOyT/sUq53yjw9T0Vfd1H9HZ6QontqFByRi6IVzdFEtCCvsf
QY5qbCzBtQkARBqLlajfuP9FQ0mMCn9AVrOBZOI7D9LgXvlKakZelTrjWxtVJfkeBz1i6UTupCTm
M4qAYiR4Ff6GAOvPoACjb0XoNfEu6ZAOSGjyiODqSLDXpITkQJ8YdvJ+7JKUQk64ooNw43OT8ZY1
Sf3501rovuow0YjZRWA4a4WI8D5/W13Du8q6Jc/8LzZCjO06Tq0OQrdIvhfpg0P4wCw1ynwHkbJl
L5vbLXSZN6eERcyyLkAcb7zr86nAAl8zlrvVuwyrSKxwSI0jonGRHfjpJrH+m3nCHswAmSWptyC4
nDgB533z8gSFpmz/W70r71lmTnniB3gaCvsCUeSfKFaC6C9RhKJ1IgUe//JxT7ZF5eYaDxSkS8tN
Vdvv80ZNlRwSy6z8rd6K1+rYixlpKQlw1UYVXc7eJd8pB6kyznOHAe+Z2p4pcU5cqRKH1FrWVgf3
Cy7H4LLbNcAIioJuwJZW4Mq+gAonti/KpJguRJKccNN8DNsWWDdw4jXH77D2dRGNMAzJ5RsT5Ipk
QA1htGfiHalb+ajjf9DqOqKmBtJxRb7pU2LkaN1FCFLLdKKlHEPdirEK5JU2jxs0TH4xUTadwqkW
VwtUBJqt22Rja3MmVCpXeuwcm3OhYLAYBe8DwkSo2pVo2mGyq4ayQaRGIA5/N8y/6dAqpEkIREES
rT1C9A03dqhrF2W4QXFLJvOTc7zVRlqcZ7dHv/QSPewO+uZiGL/I9nnKr9exIcJ5nNaYcu4fixoL
4uoDM6j7RwEuy32NwYhKjGlqaq3+0aR5i9eu6RkZwUp2UCO2zYm12AQcNl5qNHG12SBQuvMUIuC1
CCbKMkpoc5RmEK0ebHgThJVj7CXNAj5KQDta2wojifmYfWJbTyqZ6pvJM+TysIGwoK+0g1l/6+6h
FduuVSowfdvzS+UZMlqQHpjMAnsNY/1uFnstbxjlDNa1gEk/gRGoJrI2TJTUhpg519a05abSYsPR
JOmtRlR4K18jh7LLD9FnxYXpc6N+CcDee2rguR3bXpw2jOQjljNHQyt10Fubfn2usw1QNz+2MOpO
R5U8q7PlfNegQ6vNCsQNtFmzbYBDkqm7Hh9XliSTZ3cQ8BLZ3iIcdLH7qN/CdugL23ZAwihJIqmN
pzHTnEij+0i8CgKEth0MEkOSHpa3EnYzHOhM+9B4Tvk46QqzvUJ7pJoEFWWEvodOGsO9ImiWN05h
6ilDgnAMiM0IRQ+yV50OTZrOhdmk37POt+gHYySwu329u37rAzmz7CXTbtdFJD5ShKChBrO+jxmv
Hn9DIclMdd2Uo4JHQlxRSGVH3fKYBzYFuX/oduLxIq0WJclNuzg1pf87DuTRZFpE+DOp2bCM8dft
fVIf93KqhlZQMEM+zRpFtJ5Voxdy7cm4hGgg9yu0JNQl/LimQMvDfdO+Nuu7fq3gXjQbw/3k97mg
HeyRJamb9js4V28/Ilk6p43mWG+Zpfw6LKqgzDh7zDegyigoWAtxpcNxw+ZycWSKBok0cKOHe5LZ
w0IEYV6MpkBdg8ouEqqrLVzh0FIxIQ+05+WTDqR1Vr5nDKbrLdEcrz0B1dT8bS6JNJWCtpwB2VGj
MK73ilDTMLWSZAoNwdc6PFFtVjb0bW2kU8UpbcXkD/OzWJixiB4kWSgYSV1Vr5JVQnjlMrvWgyug
3wN75jQIwXidtOoMfa+sc7OvKL4ZcvApQPNTIIr6601TNN2pG/tI5euz5i+5I5ZfsQ2Od6siWI3o
z5BGhetjgXzt76IEzzO4zSAwps4axv82pYu5+Z5lu3o8xEbhcNItcUN0hTirp5Sxa0zphvw2jp+a
zkdSqB6MUmgcDeoORtqqEx0HQxv2XsI1c1Bwq8mSInvt9bl8l4Lfdws1MtbZG8x7XTuU2Xdo0AZV
s6EA0zHng8n2aDGEZMK4mdf3LKrOc69mQpkgFKzvKD6UMGNv7+INeVDa+ovJa90KRd+DiEbtyy3f
TLHbV8k5xOPRqDEoF3IeqbeUbZWEm119F1/mLak5oe9jcxyPdABQoopwv/j1peKrIGxrw9SU/1zC
Se/slS8Idi1YY0Tf8F4cG4rqekQUiK5FvpB+G6bcidCnP1UPLvYEWHrMvh85H7VldLoEslO2S3Pw
VtmC/Qw5fR6ZWek41qyAINlFe3kVLlYbwRzO1/JnT3NRUuioVHWISG2VVyKYHmjneRmx/I6ebRXD
Dyw16dxOX3KAxf8HoPYrzyM0DfWFVxtaCRnEml7DxuZQEGqUrqFiZdT1XsTph+HaeQclgK5mM9EI
YRnElzIiKRxkWtzhz1QYoggOkMhz3Q9glLC2py3cS6jfPh907NFHGPXDQm8noHF4HhIwJzo2bI4S
bEZdd+0idjLwUP2OTdgazdkT3S+XP+TyZhWAJ3frjJaLDV+zAZHfgaRBrMZtai8jMqoVtGyPkCyh
ZP2YQmnDdQHsb1F+0Smqzzob4wcTaAME7S0XciwJMY9czQm/NJbP868LkT1MSe6uDJxoYyGAremO
7C/XNWZlisRQAU3TVh5oRiKYAbznoRwz0kbIwVyq/fhNz1TMn8dITock8DLeSMx85gEwgwwRCX6T
vVelihiNjcfsd5W4ST0XgTqeNn5kMwGTK5D0HUvQOpdilLIsC8XbMVs0tg8qOVIhKPZGUBu1SZFp
khrOLCfwb3GuqONwUEANp6UBYaXHoFHtGbEoh6Z32/eqbONr7YH0eJLno9idgY9/FiLUzF6+a4tK
ih3ymU1XBDLwW8L/ryzNMf/AVERayz41RqUApAXNZ15PHbuNgoQODVURhLq54h+otftnicsF3FNI
aJIxM0u7ASEjO5oqU5UcqImNppmdqfI8u4rsRrbtD2fUch+VvQXW7vI26ukK069UIEowpsnozqqJ
YGwjKXs738EYeut1SDerk5LDDSF5ulZeBywRx2gzqJg8NRhsMfDkudoF8roIaAcm52d4eJDHtB9B
9TH6rnXWyA2BUctUKqAwvp5lsR4+4qD+p/ZTsHH6tAztBSFLQyrCg2ooT8HTe7ynoMyixvwFjg35
gL7ZcPQAOT+JtdDQ0zYyw15CwskhaY7aqyWS+5aokWjsDYOcaQD87rPz9/W8J49pCwMihGwJgCFH
CnNPswna2HP9/sRYp3MbhOuZixeAf+KJKqUSCpCYx2JoMa+vntMXeT4YZ7Xt1GJD8Xj2KukPv8FN
c/XpRgCXRGKAeJNH4Qa/XMKmY9fVtRrl6yJSvqaSrzmtfaoAMo2depPFWgsya6MCzi2BnQ77lSka
ieF4ES9rIYFYYQ+n6bvR9xOgpa2xXafd9ztdP5CMr9ig8f5AIOEyYVdBPNFamZFUtO122/PeDztH
ZQA9voSnwj1KnhRm2e1c6We4iQjKqEFxrvo7+HZOgqJWMGqRp+HErxYPHaua07VqeS0z65zTduLM
3SZuAvUybXGbFyxdLAbX5HU3fVRDvucrSkSeQXSDvb9Nm/hw0cbfVlnrIFPtSxJpHPsQqw8Wowjx
PyCJ5LRw1eoG4u+3BCT0pL82AiGhVk3YleDn2L5K8A4sgW9pIfHwAg2ExB88fGL9ZOadfqkXxdLS
9+ejCYh+B1gRxjls4E2eH1BlDq1AW2duoBFwGdF6o1w4137OC9PpUd76XxdR2R/wwAs+atnUuGZz
zjnIJtEqk6tnCvuZym3xQSE5+KmWHCMZAnJMQH3fUhTBElzF2NWGAGgnV/6FfMI1sAO+DsL+6R9V
HLcHDabt/fdRWUDIys04tnx3fJbYI49yK7g6jeqnOqXKUa79p1bywvNJTrWKgirv/utoPAzsy8Oz
a36S47CvnhrC1X5gRb2J4cOB8jxZXLEJ+wom13bLHViCXlNu9kvKeyrHMy2YoZbiyOydxBT1iQKN
UE8IiZpd0HNpGmgHHuc8NtZQ0DnxCefAAuQgwaZf6lbGayziGlg49zsr1FAL8+t6Iq4Uhbjr6sX7
AsFwS70Uy9Xcp66h/Z4M7JGiLA/aVC/6Ky31qkxOhpDLK9RxmN20vQekLE3LGt7T3yopACPuVd9i
gPzyN//FkuSd1AF0tKSJDYsXIP8vJbH5w04N+7X3L6EnSzVgEsRAl8WKrrhB/opQhzpb6SmvuYYR
5ddx/0/zmfK8zrR6G1m/tqgJ25Y5taQPDz8ZpLYjz0JPnk78ZRjggQW9n2NywkOUu+JupsNloid/
rKHCNzAC/l4ceIJIGwe5Y1yqVVze/gx8Oj4W2WvQvSrtzd4i1xfPJz7KvmRdH6L7XorbRfo3SmIx
bWdiAn7YG0rRUA1/5lS8x12amZEGVqW21QSCVfulLILbA2+BwRfZA/EAgw2uirt+69x+69njCxAB
fCJ7lhTZ3SDXuSQ3w+GZZr4DtrRnFoAfTof4XP+XX6kTwAbNXKYFn+4/euXO/mbl1uut90etLeKi
WVefdTyhfLJ89GDpqtIN6P4hweq8ZIvF9nkqEd5yqQV10znF8BNix4ioo+7iCJSliScgUEskM9Mb
jq+hBcqhc5EISYyxgAMjUba6HxGNg9H9vdKFRehWZoSls/Lq3PY0EhCntoFJnAicNqYipAD52EWx
2TsxIDi3vt4v/to+BLYT7Piao3d2fPQoUtiNY7zvGaOlBjNB8VkaJ7O0dmPW6oI+ajutE+o4t0or
4D/ozGAaaenYkLdA6LHhCUJKhR2FL0byQXOP4qkY2zE5Yi+JHwx926EvPXjLhSAUN3PuMQrD0Prm
goCtkufw1WWckUQRqZz9UFcbzLAqmK8cfq/0MQ9KeQb8z68siCDzeApDTUyeCS4jTeqsjhzcmDrZ
rzSpu+EMtsNuJL2CxeEqDK6nZTKewSJB9WLJPG1r0vSpIhivbmWnbWoaVzrYpK9AfsYSY1mQcTZU
HNSejySOcQjC5jB+DDtDsrk9I/4OwIdlNKjtANwahvnVvp3N1B2ZrCs5UgMv5dlwLl/esp793nZJ
QrsP9k/C6aJ2ilZEz/m0RRXfFMn0l6gYuYtR+AoGE7jsIQA8+H7a1C5GFX74LSKnypgnGXuB+rmS
CYMRqwn2X9W/Trkb88E8MWlQYOt0FoNEhZCyXpEGkDGoJAOpmI5/G0R96eEy4G9y3OTZHWAECP2J
9Mn6xZhYcUxI2SgVXTwwY1satuxHWZBJ6H6Z5VuOEAQo6pKPpqM8xbQoy2sBD/dD5YP88pT346oX
vNIwoxtAbgYwjBahRpLZwFiqbQpfuyFtWd6KzawJf8ia+4ziEgaxysEPIsq9C+X0X+P9KKa7384+
a/ZhC3NeLlUIK8E9PqC44e54fdWaaOZqpy6YgDL4YhFgGETaEiZEP0Ul8Td0oISkyIESwTcGtDEu
JqFVstXnjBESuhBBNOk9d+7uv98btxtW5TB0/BUZlhgo28AAw4TiL0yisxZtOmvNUwJcSQdT1/M3
TtBPXxSXbcVopzqAuV/fi0ZFnpvdSrQJNmblX9rSa54jNgjmwZhsh+cUQY0bU21NNQ65HrJ3phAn
bgxQD/BfEsQjbYYO8hidql6bXZirKmhrEYJABmiLQ8Lc3YS6oOr3j96/Ps/REr++XLyUX9dmiCPY
0N3CMFnQIlN/0YLQZ7gjQ9f88qeQmAvZa6R3QiopijhUHnnPjw/KCBfhBEnJxzrbgVwRasGroK1u
AqAcBX7Y4xYZlBd4Z2gR0ed9pGThPkGTwwghep4yBxdB9FWpFKnHjnxNMJEPIlPMaTKNxZvoVdqY
8W/Wsge93dzKLDn7KvYTKQCyMd9GgLspdJhTVkzOTYeFIPPyJdZLSvMhz2rviCy1m8IGiq8Y+pv6
Nu/HXf0pD2T7b9jw+WbMF9GYk1vqafGBmrv9IVFP1lu/8ZsjlW9ikRKgjfSU+QZlp5h5w8NUBBa7
BuO17KTiF5972F26TQIP+9Y5sLDA6y/N3SsOh8dUmLu9Q228aSsrIHfvz/IwzqLcYQbPQJpDbSyk
NYXYR3JHYCnEu8uNukCiucYHDC8QZU7h1cM/nknUzCaKKE27z/JSD8ZAyNqaXiBRR1gcNJrYwNDw
Zro0FRtRjJFqHdj82ZNGijR/bnJ/CfTQuT3sSiPCqRLvHzKj5aiNpD1X+BRfJQkEjO6SwN+tEfE6
/u72AsbH1z/veXEwOGzqbgJy6JS5BRqGAkFGKKH1AzsrtbynU0P76wy4Pdr/HlIQeIDbIx0MU6eW
PdETZU6LH730UoIIiAVzi0LxwM5NPKQP4qpS28eSIcarcIRqhswwMTJp3NAma2KjY50v2SkWZuRq
KSiJLSboS2L+L22g6+QEwOrzXCGODx0tsb8HNYfu4cvhWT/rYtrqFyTwnPhCkqIkF0A32DdRnOCN
I4Mj9+p1x1Cd7sbm95lm74RUNSi8dm/pS0ZjZhvjG1U9lfZk+MElauyR6aG980nq7n4LfGRD30zI
TfI0epmeiywEsvsWpVAjLf5fqgxpfa+xG7ZL4Uaj/6lJ3ThZFiy+eYTfuw4Lijme0ONVk/1mOZwi
aiDyJlLuuNCfJIMzsB11RCJ8t1Ui+5nlwUyjMzT8LZ0cLxfBpHvoHnhTQX+iiAbFG/Tyts4L01GN
KOCFvfQNkGAaBdzzv6iaTVPRH4GZ9SXZzdu+wE+zK6LqL8vLnYyREicSs1Z8PAijd93BKla9N6H8
aAxT6+/qHOcK9msTugWgVADPYfk0gaNBb4eg+ZkcUV2xBAiNTTzaSISXgBLVQuRb5MVkLGnkqNeD
VOl1NNxAVCvQFerxwdRbhOS7tVXb3G1l/LM7tdUBtvZjmtvx9qT2o6Yv8GG83qj13S7fG0zPKQp1
pZvxzBDHn6i3vamlAzs7ogt+4H27C1t9lBF4JH3vaqiqZofvb6lyOzw/povzprRWdANycA9lugn0
/d5UEvZOZLk4J6xUHWqbGkQug5+sBkbjUApa6CvR7cO+tS8GewRq1mT4CVEqPuf3y12aDaftVyBf
55B0hA2r36zPclYlN8mkcvm6f7DA2vmquFoEdaxef8bqoNeYx1auWIvCOi5Ug4p5mnm/hxFXcLEc
tXRLub1c5h2sh/dQXPjckSQZhMndJrbF0/LBoC5BCi1M7+BO98qGBt9wVHDEapoDjI0tm5abApCP
N/Y0DqsUXgZ6q7xK6lFthojpIPF7IRckHrVK+S43n3zCczK/4OYbTqhg5g0drEWWfIygYkFI7DNM
bpFQ51z1ax4vSNaVj1xCu1jtleWO1gQipO0n7SEw4eRj8j653V8mqh1La6N9wmnv+gGqr4BGQ+Vw
XOzzgQrX53cAdHh4Sq42GHdR9YMOmF3u/ARXwGf/FQnJ9R/lZPsx0HVADZq9r6y55CKY+6VOLGHz
hm+KJQrcm8jl2BzHbArtB7BVNjv5iTsQGunheEFNFQD4OfLeItygZmj+/uCFbDHCJU2+hYdAay6q
kT/ZWTpHF5VrZUYDqhHi+b2UHp4b+RrM2LXdn2/1/0FkKfTCSrYAE3vYPw8vW73+4kv3Bqbi46+8
XO6XNY8m0by2GYEpo0JH8/y3SWf5QKbcto+eouf8BASWNWyGbmsByZ2zStzNJ82cjcO8SGQsm+KW
DkGAT0iCEiZ0aEIBmiFKS55ymqeR+JaWmAn8EPuOyexOsCUWc0CFBbHT7BwiCTD/lE/zq3PUojlW
bVrskVMEQ1Oi7DD0YUum/XPLew7bNbzblm+pwDHiEF5WEF5zPqulArwellhfto0HXAqp45OuB76M
hwhwtYDll04uwuMe/KpfBA1bQyJLJ/ci33zHqWbHJ4DksxEov46Hn76PGF+nqAyk226D9Pg5WQLn
dn2GC6VVxDjAV0EOM+4Lg1ye7gBmvr+lPtwaMoCZrHLGGTH7lhzSj2zGrd5BkLtRVw1YtS2m32ic
6JZRe4p3mY26QEOH9X2KIew6f69LiA8gHHOH0u9wTmecttS7icI9LxwkdwaoWcjXwiVkjwRqr2h6
cXnyJklPyAOTC+pZw49ENpEUOexBHhqUVoGj3WmTfW2sCf9vW0fnButspaSKCV6qi9cxEs+VMaVi
1uTWQgzNQpccsPzUvb7KozEC5McR0KcMBDH9RRHCgzssme7mPyvAJLGiQoWuFDJvi33Om+JQ9Gh3
dc4nPy7vFz9FeevKlsJt9/Xar7UzXwmRlKkGg4ZUj1P4U5AtaayBHsiibOQfIPDLR0sqNshoTWDW
aimADgPv53D9vuQmhKWAbllcbtnwq/Jzzv5fpm/kvsGOqPgtvy9iSmxHtySQmzDMKerDvjhJrKfn
XYT/Gcm8HvR4S/+dg5DLH1B7Q+lAR8/GlWcGVpjWyAmySvO5C25RK6/kRtQqcq13p2T60VY6fbOF
mL5wBerc3pJ93bt8VhrN40kfplHDKU21My9bsLQ9cXlAKRrhswSF1x9v/n2PRsvijHpDJzHxGKWP
V1n/gu+hTwCVxcb0mFYORCwEJDdnEFqS7guhw3/0y1uvIOIXRVPUUDgA+nxb7AcMi90W6KroEkCF
Ej5YFjiZemANeInNwy/sjWTvzh5UNoXS3X2LBoFv/F66H/cCq4lWmk0U8GLgTQUFUNe6Utwa2zHq
OI03tfFM+rZW6GXh0sSPBlRomNMrSImvb3auQHe0qVHI0Qz4a63VyDQnTf2KFDfngYStgvsI6DV+
xj9b8A1d7BylfInzNjqE0ChaGKf6LJs/BsAJuTFV+NZAHI6efbPpCxlcipAtvqcBuHedooYVRVUS
M908XrWl/LlHmRUMDYwRSmZj4zSy/YA0jSRfYrJGYawml2S3iRjQ1uc1lyI3dapAavvZUpwfLuyL
ynE7cnBySBka+DiMlJfHUd+nSpx/UaI8/owa26y6x9ic9jqYbX+fOqNhkbxAqu8lUbyqn2P5WUyh
BBJsQaXjkY0Xg/Cuxs9zMb7V2S7KcyHETyWqdZAT1AkBLmTk74DM3pyeWhYMtff9ZXK+sT+U6g0U
894LS1P1jAC+dBrKPFuXhaipSpT9HposBV4lzzjvFn70gYIbIwxhsa5JeWTwt0Jm/vaf6bnNzqZ0
Qx2ufRbFQlRZRFGnf12PPE8u/f42pwaZGj6zkCEODa7R0wfR6JjFok62vuIsUhTrPYUNk2BSp8/Q
QIGFZBiESO5SjVEbAEwNM1wrC+P+r9ypLayzNNZ05w+Xv5KkqJsAYS1NKgzv9URGqOhg4mRdsFZV
oFv/4NmHc5/eQPbPrHwJQb5wvkd69XiPiaZVXYTsX55tRhcdSwjk4nTDO5yYSwaA9PktddwLi0of
yYAcf18FoPAS/L3gSF6LazND+ojPgOnHVe/5Rl7ZFll0uuYaqt46RqJhlAI/Y//Fd9suYCBTYZ5b
f7FRiiqHgCvfHPEPx0sg6N0FZ/gyOpDmF8HJUOXcKGQVcYXNmeqIUKTHLTYFSFH/Kbow6oU7CGox
cbv81OfataUoCJut0P2lthAO7rjOtTVfjYGaAhkCoGtBVp43vPB5ZCD5Q9unJYEJ0NqKoi2dOluC
QRtuCowqfI2E2/tU9aVAFGSSpaYccaahBISPlWWWtfd04E9TEDcX9N7UHhtDuIS0Y78K1HZ3gVy6
KGiiphAOyIPDvwAyXHLB5gg0bzkCdbEYNYSc58x1JHCxXEXVCTsw/7kjYOcTCF0ijdYt6B9xGRgi
tRaJAocX+vV8mWLrhS5vLcJvPgEoy+/1bhQyrEfOvL3WCqlDp5dmyFrnbKIFsIccFTW4kpAUQrHa
O4pB+ZlikmrBjijTTnHvjhPcXOHqRdKkmAqeqf07MsC2fCG0waNATldOsUzB8HaTNdoklnjf3xks
DLJxRhgZGVNLKHlP1WL0VGKdfBDqGuup66gUXfhmlml1nIVW00tS+msS5+StgeaiERLtWJbfIGM/
1bCIThjforZmax17i3U8iofL4AIdL68Gqm380mztKM7uYGg44nlnUWyj44ljEc3uN665rq7zQLZa
ibGpdkEYpiaM6rfrTJ6BDJh3yw9B20kkZbXaKFIcbQVHbTjEhB6hTZoENm4/t7I7cp646+ovaSGC
jTCxzntbYurGyy6EeOUNsEy6ab99w0NG8o3pVbcRQjzsMSqMvjAZT/Hqbu09ftJH2yFticMDrakC
oraxMNKfGaNe5i9YdKtyvNo2JS3z/dIl199kV6fZXbK8rtT1OAcmCz88I7KV393j7hqcmf6RFKL/
YqTwy2E9x4bW5gV9Mg2hCKPSMu4nxRv4AhnH/Gx/0nBTy3ozFiYs1ep4nbwia9CnqEOHD0rznP3i
3iSAelUNrqXU6KAMeP7NNrWhAsrcQYyqqOXcEaGxNdqGTaPkq+BncXUhJ7gV8MaRDG4HX4gJ37ua
8IRmt0pcIQLJXlDOW1JKPoRlPRStZuDQbhmkGztUDHyxneCqXazaGia7ZyETFRDLK+fp4UalQwfF
QCekdfksmGltsahNG4RAq9UmAcrF+1a0AqG3pkDgQSRK+QfjV9ZRn+3gkRlEEz6aJ+E1JYRuyHJ/
NgiQnVaK0NKEzn0WFrYpGSPAXDgkLw+ggUIbfHuDD+XGG36MGL+eggPzbmzvUydfBoFVKJxJwEX1
0yrqQ51jEaKDv9MxcZFfvZSm3EZZ+7gQAI4CvpyMwCHgFSxNaaTRO5D3I4tcI3LmwSFRT7JGViKr
RIuZeAe/ji0DXhVdY+Y38TRq/ciBYKVBkIlde2HbEiOHFWYBUK0sPkFP87209KM3dVujg+L+x4AY
R1TVnGDFRepgoCdQnRIJicj5loOqdECf+FZUVSGUwpCK2//ItF1m2PVyv/1e8mVDiUBPUOWQuN05
z616moDlu40waV121yqc7Npev5prbbo+MNdXJLnPQ7nuRh+l1OtQUTJgNUrQBoL8SFGGmpLMTQtW
F9fhFCvDXwH+faT+FmsK/ha8LKJUJ98XvwDa3YuFA5UXuwlmM1Soqpy2vMio2rx2uaMH58NAJeAU
kRU9Ivq59HwWvyBGevATaZFLkBLZUaj+OYO8BE8LCKJyhgpHQ9fTQ9HuTjn4ZLgCkkyVSg5EXJNt
5843k97Y6CsSj88/yMeCGGqPA0ZdYoYpb5eeDbeabHVeA/6OGUVLgaCouSea9vFoqofbqiKKxbCs
IPsGNpMkzTWmSvMZW0CKiN8uLaiihqM6U13n50dIMT2V5+hBUmSKd38YeLa+xpPCDtZ2PkF+xwhm
t8myozJQDPl+ePW7zUV/kmIuLhulSyaBFM3U+scKBSvq3oORCV/RiMacdG6kQPue9aHS9mO+qHNT
6kxrjYgiWr259HOlZEEgWnqopFfnF+zFoPq1fo3KKDJ7VWz2bOaX84WOgP5wkGGEO+mmuNDUqCgz
yiTLKJ/Sop4MxOiaGgwyPh/T/qwaQIl5YjDpgBUIUJLW5nlEQIAuNtKrcAykFDAGAlFJA1P1bKbv
P3XXNT+czaDCv3UehwRgcwJwlhyOrKTIbEPNPc9Cm2LQdvezsT9a/DIaCoMzbRmdiBkEHMKCgN81
jfqyIXfHBRi8thPJnJtXovQ3xHK+B550P0RSFbOo5DBOFhxtu6RBYID923hmmzSWtw2q7dd1aX7w
ry2oCEN38NSwczXjOIeqwsFWU+A6Z04+iiCDPStsTbSGycC1twIxcDlNzyfg/hbxgiJeRTgQSnBk
pIJwdoWxU5XhjlcgQ8JKWKmoKZWYIonGqJHK0uJ9vefl+P+DAQQlmUsyamAWHqmOHYV622ueycrf
EGbYfU3xGxpqjNckIGdTJbNLPTsQghpXxf9o3yTFFTULuLvkVfBZBG/ANPXfwuBNPA+MvB1LfzX8
1VI/kt050QfN1mwlLMeiflfKvH+hHvGXgt5WVvgjyKWDzc0c/R1D5ySGJi0fSyo7bBYGpo/13oH+
5eNRnAKo6AxswKaynOlJIsx7GVanIB21e2z8oxlavbWmcwm6mzncjTeK1P/hpQmYlsn6Pu/qecBd
YpPvKNbH5dDXp2EmrHi7pr1UGTXN42YeSbpkZ6diM4ABFV+cTD+7ladraQ+hwseYAWYHT3sytKxy
YGSgNpkCbht9N0pWYkH+kUTUaq1On7JeISMcO00oOJ2UpKwjN7KejnrE+7iIxqGMQmNRztyAGuCs
1BcuJQpNwpVHSjFLIPYB9fIX2x7x8n5ZECcOhubJpZJ/vEzB8ryZ1cMVES9pQlpDNudpjtwbwjhL
t02ayQjvfxGf/EEn1xCgPmRcnDudGMS3dOgheSUEmgUDqUYhT2vj5w1+g9sToLi3GMiWdmCYJ5ZM
oydCViKzCIM53efvBO3j3IiEObST0AN1HQT8SGzPmcDzU1iCzGdewIq9jjVZpOy8txNc/JykgZvQ
Q85TvWdOxxMHyvUJBGJR384+c43megE47saRStNQExNYzvSaCuUvUaXHuhUpP4Fa2qrDxCLvfXwz
aEcvKPnmEV9IfbGFSMfBUagckA94dA8LA2nySdTAlWfUwcgQzjQ7fHtr5gExjy7sX6Cz4Od8Vpep
ExzIAI+i2mH3Gg8LVE+0gnHjZAVyvlN1L3NG45r1Yht+Ly0lnBZXpahXWMYCMDa2UE/0BGC3AYa2
8yUyiWuFSZnnsCINEVJjrJ0k5Kt0HkLNRpilalBmODQqwqv8nUI9wATWOUzL5GtXCuCTrUtCpi1Y
2ObldSyxf9jC7I8ptKCIQvXXUDc2kr2pJ2HpPUMlcfIly/xbcTLoifvSYNu35ffFo/HShR3WorLt
E7guXv6vYdesSuBqpDMjsforVpfG5xwDQEVpt0wHY2YueanKhKWlNdsPBk8CSSLQSikT4cJ/cQbE
KGqZgfAzhgMABvFsidE8ktxaKci0ytBhYeUFWmH3TPOBJY2Q1LcoYat+GXx6W2O54Q5vGEoNSJsI
rEZ/uON9Hc9hI3zvgw2xsCpizF9QEW0/v9WIw+URKf9Fz+Rn3GXHCJQBdGOj7SiwTuOk1K2b6YrX
2CmVwJwpT5d/BWxu1M30U9BQ3Wa+GkLWLXVUWipUH4xVBMJ4AJmnyWJpD9wKh93FBb9JYqgRh/4l
XEtJ8O7Rsehbos6SSMQIUU3UhM4vUgKdyfQNT4hL7/3fZsG99dE4Sdd22jAftTVsiMeAawTxtnj6
h3T1HCiT4VHV4PbCjwZ1BmvOHsYKxo0HIrMV2J4Zw9GtPZ4ueBCblFiVG/77wBd4RtvtwzV4wYDT
Gv/8WscDr9anrmOsCbbt60qk/+ux4rk08g1C6hBqHLHK8wUKjxX+AxbwCyoTsGR54tcO4aSR5tfr
n/o+jR6yBkrdRGDtK8fLyZ71fv5a9w+dzS0qqIDyUDbSmGf6HvbTXORERTLTuV5vKvLo/6jobrLg
ETrz8I0JFwCho7PlhrveNxx/LJ7mr5/wQrcpcciib+JZOBFw4+76fLdTp/txHbfL2htY7V3NDhw+
pCI4xEyOJybro2LnDYSGiCrlWOkTjhADeB/3NZzLYzamLC9FKRaLfePO5e37RnGJqjYVAPl9T8VO
8t0Ms5cS2Dm4cTj3qD1Jmn432dndP8vEh95haGKx2hXmX5HkujAzjea9hvXGCskq70lny4csl/ld
BiqXtQxTcQoiqRcvfWC5Jn19tvVVQ/cAHHOuo8pkf6TMY2rhDFZ6yOljcCtcAFmumri1Yb8aG3QJ
HcY+VG1/oq69Dw2ErMD1iZlRbar3QKKd8Q9eCUb4aARpCjEfho6RWYvapckFcloAGZV0SpPgEyf+
vv6eTwdTjU4wIwSpU4MTzuxgp+9zYdtRZ2kV6I3SXPCtlhxxOLGiTbX523lZ+LODmf2/7qMasMtt
nbkYq6gfEEt3UYXaO5x8I1S3QaIzvcbp7W7EL+GUxRRbZbAJiV4prHdZgOXaKj3SRrSMQKphOE4L
PiCOFFtk61UxGw8yAyMc43RVxzYbe5CyNXxb8C5+xD2/ed3tZZH1pJJ4JuZO4QDne0VgS0nAAHRF
cgfK5TJW1yNep5/EFd9hVuJjbZllccazmiMvgn7aKmbGs2JO0rrYWm+uUtnzqq5GHtaRZBS7EqzB
+jiyw9RcRRo9OiayQhxIdiENy8TVSM/RE8Cwp8T+ywOSFaXZhEtTGb8R6PNnRo1/qPecz1za5/Ux
xC12NDWUtqDyACQyNfqP42IQG3GC6RmBXCk6xJTtPSWrOjJmYa9JXYUxOo9/pXIduPPOAxeVitZ+
67gz3yeIftPzdqZ8M1IxmG+GKOIQJwtkyuEd5DZ5jgW56O1rOLvQhqzvhdXgcOzHKnkMXrGqLAK4
P/8L5QVmEas//KrHPO5d6IpowTb4/kNmzsX+Icoz0BVwECTYBpHsBEbQVHxbbTrs/mOomBLWR15G
EZpDo53xMamcsTy5hdNHd5OkvP0kKIyoYDXV1PmE1w9zOAS5GTMLNN2ltHQGlfhiqeprPr9ODX6C
d93Ax5nuu464QBMaJVqJ3Plna4TqP2PuWmZN5k/U9hVpvS8nPNI3GRCo1StRsRC8XOHYP/fPJ65F
jBHAC0EUR9d1tuDDjdrnx3EYs0mQEcLzYEeVhHML04pAiN2sDsVYJefYgDomzjOnRBh3/RsvT98D
LK5kUTzBrZTPJSQLYmIj8SyhhhNtTsdaiJzyKdhcUQmwGecoor7v3PZJkGNtmJ/ortJ2APdD6adV
xLC5xtFL+th2YK6u2+zBY/xeW5kB866fxymaUFc2R2pyKmqtfiywCzxPZt+2EOrVHjQM1ygIkbf0
7gt5xrmAl1hmGW/iAbDa2sOq9/kE7vOai9NDH52z/r/csTvlYAfLablycBgNGCG1upVw8nnhfgVU
eg3knSGV9tpyyuiLrruH4J2kyyZQkpWlAuHirDg6Ih9rYspo2nTZe5IDb7Z1nmlJ+NFelozSHTt5
eDvwUFyTa76jJomcbdaOrFGOKYTXHfQGRVRaMYQmonKBJf64LanAPX1iEwjmgrZ6jdvr/pn0WlxT
cHLxZpFiSobZNv0ODh+lp6ypq1psVwGL2IP9J7xyYJZUqVK2E2G+Jhz5frnFm2uhMrYnp/o1J+1C
5aw7hwOu6kcpLlZORvr80GgLh6zny82GJPhG8wdJf4XlHIWcZcRgo4PUcQl2wZLoo7H0KbMEaN89
zwIzH9iE/a3XCLNHnJfm0b1JANskr7nH+8bBaJYt8Vdy5hxOQg0stU1lh9AoJaPz7Kv0RR2iU9k0
EeJqxZI9KdMwtt3y8PwD9ug/ruobrGoFB2DCNFVbhJAsowvdPbr0SuTfQbD75CkRuFGPkK4GG0Tt
RNImamtoiork3WYSd1VqQgG5arpKE2yCA6sTCD+/ijPIJnwNj4xOU+ugp9RznYngJooIJ2WsfjRk
3N1gCiRURNuJqA0mWGdr8b/oEUCLzPDCPjHI/Zxx4lCCOuXoifqJLcGhgU+eKXfYc9XuOf1Yj4B2
v2pcvU3qidfWxcuNCcHpNmJK1zuUVaJMEES1cBa9072zf0pcfzCD3GQbor5vED3v/FedMYo/QhPc
rYEa3wUzyVzNRpTFkH69FC1p7WwRkPqkGWF5yCTfTwLXJjVQo3J2mhYamwKkFkvEUDTuy4kBIcQS
tZyrStSNUAjC3EWe8vr092N3/orVVtnbGR+WIppQjekUuvLZY2c4Q8zE1llr8OhIzXviJ/d73IjD
ErDiOifgaDhRJKoyyGTClJ9SXKF0bOEkAutHweFwjP5B33+za2uGgsJS/k14TNxccFLRkEw7wjmF
uzd4iZg5eRbqo1g/HY6cui7j/ROE0x7RbnFp44KU2FauorPOZHIidI23cNUajC+3DgcFY73VUIwP
xpJ0AtNr0SBIoGw/f/g0Eev1kQ6FeKrc/eoaxGW0e4ti3i44N/cbw5xDfybuqso2SGxNAlWZQc8Q
KHZ22csHFzbUTRKp3VktpovNkU6+v1Feuza1sxGCFvV59a08M/EJRnR7bNI+D45/pvnZh9uhmzPr
F3fcogs+ktBm6RZ2FcnzjzpT1l1mSiDWeY2TfQ1We26eoHCwtqcGc72OqPLz/43N1WPK+z27Hf5b
TE76dSoqXsgC/C66o84yeEjbXo9LQNg1ZtUvKipMhJo9mbwNJuB55RnHNaoSsbyL6DaSxlyFABZS
WZcvZhP04K/xhBy1nCi4898xzfSQp7oXW9Gh34tMoHdhsjySl0qJ5apIG2ENvKwxGbxX5XvQVB7O
ov4UMj2Z0STDZFjfFM8Ro+pxO8SJ42nqd/7dqsLSnvA1EaGdl9Zz9+Tw/ZU+oZd5m9ScSZB6B0z3
l5bmLKL+z9AEjBw1l3kRAlA+ggx0TCCaZAg5hzJ5IxDU0o/8phOhQBw/aiE5mAqv7YhQPnMhjqrV
3oigVbkGiM7RX8RfXVT1CBauM0b9dVJdgLtqA4+VC+pT87plG5F5KYdjDv5puhosexQRCL54mc5E
PPPZ8Hy7XDi/6hrVP/o5GvC/ep9gFIktdyeojV29/wXWik35JFaEN0ky1WusLY69TIrLIgbzW9qR
txx7QANXmp8ZNnhwpzvfq0x14YhKBWnx3NmfDkzNfMUGspsv+rKXT4RWy1sLK/PKe4a9KjHpQkL5
qeLopL8neIJr3jXRKXxrUzbuJldkmmG6nAiIH28L6qkVQYZI+/jBTHfKUOz+wR42uMDXRlErbR7p
vA3/5GqU2OJZJrhkbvwn7caYoScx0qRWnvmpbEuyRdVDpMr4IjpMsPfiENIQrnZu/oQZfvIJ3N7u
W1CoXiZIbMcDiAS90itMvXrSNls6Sbk48OZvU1PCe7NinMxw59sktlYE185DSZIUjj0VMPz3OMNc
49LmIV6eG6eNwrY1fj7cswAjnflM/AnsHr4BLLYGC8MdkM9Trz4gInNewLra2O8kIGvl4IqtpR/u
QUt6Qs+VUtt7E6CK5wolXEEPbg2GQOpVZiY7Pa3LhyE+ynUYICUX7hjKFwBBVy/vYZ7636c2nEJ6
6hxJbgUkkA4O255R0wKX08rXSNfQ23GD/TCNg9Gq1SAOQCCfDyCP6NTSofcFf9rcWUhVDbjjNrDQ
Zlz9hxrO+3p/vrI2xtlGfkGKxZv39f7QlBqm8fIHOyTyd6Dn2LxPL0yAzgdWMvMUH/IjpBog++IZ
UYpaUYQvqEleay5ysfZ3sBNvGvAsEyLyd+QYxEKs8vjgCatunZDkq7iy1JjQrzGvw6vPwqOXGQE5
/YJVoqrYmfG2JUcZqKCmH0gO33h4K7Doxy0/dYh599gbvLaLPcH9cKuxYRojf5swbYFvjapZT71/
C6PBzthicwwS2XgAHoBSPwnRosyMcxu+8CruSW/eRVUtv7zut6PzYX1w1LsjDM2iXdZeyWg33bzK
pb+G1vw9GxPU4ddyYTsy/FB/M7SH/+j8ZQK93G2Afa9+a9Rt+jdlQwpipWLhVY+TwJtLyoz0eziN
xTs9VwFyh5kloM5DxakchKiWnQ9fC1hmtsFTJZYBzGYgsPvrJ+k5PomPLRnftBu+PqOdOgzVosvT
egxki1m1LLsPG2LbnGd910jpPIo8wRf+eHL+zn8rLCLRvYHj7OXJ8afVa+qhoh58sN8AhKyUrBxN
0n7+L0kbHCGF5t2UVye1mqSuaJ/1lrvuSt5g98d7myEqYxy2Y/DcxChLkeHHLuhUaGjM+MktieSF
EvPLyRt1DCf79rFlNLtSGadZOM1NwZGcMAriNQhISQLuDOoSVlNkPnWpxYczeoBJOk6b7PSlTRJH
AJUUQrFT5nqD96ka8o72as8BHu7jDdwO0+QYd7YnAwa03ohyKyJMUJ0XjeUe/Ac+S5YUQW/1lnQl
w2Gq8HWo0UmHZhQXltpqxq/MFmGU7TnEtP+bNgSCdiPCuPuViSHvyrV2aJIvuENHXBHugzyL6fY1
bbf1E3eNUpH3YmLko7Dwg/zOYD/a/e3SsGzo4BrHZEoOH1dyXPRS62U4l73wgz6bCCy1Fw20TV8V
QuAMwbI513UDXLN7/WqSUwXDwxc00si3pBz8QGTIkL5XgevfrwjqEZ1xqQU64x3OswzIvnLBguE2
pr+gxOKWYfjevDVFz6FZOYtiD5z2JGznVSkeGsAtjZtok+yfrWSaB5ppeROE4aQlVUu1a1X+T6jw
ISDSn7YIuvdBtb6r/zUTaeXxWaq1Yf7GdObobh3twfyxsoiThZjNfj0XRBYkOjnMK/d4hHpYggGX
jd95X75T2xO5cA+PCI37uYWbLWSvH1coHCYqfmCo10ei9hrczQ9Pj+mYyQ28Mts0aNhurXkkLp8z
XN5rYMge8wrSEE3WQYIbn4q+Aae6hFpm/UDSEwRXGR+QBj7LxIYGnGqpT4H5krfwJFlsOROUt2CO
ieeaeQ0liRbn54vrfQKNojyYdluGlyeDJWHBgFl2XeyC/s97losTh+s48a3giwdfFBMEa94iKO+x
SKaW+HdGyVViJinUFX57ueyfUExF2XHHgMbwmF5iboNvurH4c4J0OPHylUNSb2fSAuSHD0s2ShLd
o4JIf1w3ZHi0iGtZWP5q9AZd6zPCaa311oKCMZO14hp9IL39oWckA/1cexEHK/5lr31OUZEoqVP6
GPmxWGFg7ZrIOeJcV5TczPpRY6Y6R/QMYdDqKaGCKPQECay+viwR2BX0ztfDXPQxKwVcDvF9YsDw
hEi34v8A5PN4U0LkzJ99dJktFguTzfGsuNW6z+nX0r7AsZtEPGyiPUUzqv4HOetObeDcU2LpEcGL
UOHauW5f1mhV35vbYGAQfSmfukcYSOqvLzlktRyLchauPU4dVguK8Mz4WQL82g43qpS0HP1E9EIx
vo5HRP+2CzewOkawSBm3TjbcbVaLVecxMF6q97bL/c2m7UG8egNProz8KX97mHqEKlrCF9Rncml7
vmQ/Sgrji8HTj1ciL5wGn7qwSXA2l/I/HBSPODD2PkRbmajC9jerYgFIjs4e1pTp4cOD/2INIDDd
i4fvqRH5lLm53hRJ6fXzPE2//zrVD0kbrDd/INdb0wkiik+iBj51zfB1WvuiatiZCXfIMLZZru3B
z4MDfPy3sLdmaIKqz4a8qPkm5FsU/3yeUO/T23uSYUdARX+Pl41uUTTn/8wk/Kv4JIbBX2h2GHZJ
/JHEGWctZ/CbNUzImuviwJ86daAyToqPViHGlxySNdWbpOx0gZ4A+FB3c4/5v2YBNynR+CwyA3A1
n0b6Y8wNgp6AlqD7rO9KPb65ZJaCYb68wxqVS4+6/VUovuGcWYw53EV5MHFU8GwU3AIDcS+yjkrZ
Y79pgx3SE3CYRyHMso2paZp5qLCLuXaXOb8BNiecmOlaJ76BmYOcEFLL1HYcwuelDydk4fRMJNZA
ksK6jb54fAYVWjz4JNS2sdCtVyp3cSXB8cpU8+8sodBU3htJdGWo3tOi/yuXraoWrpg896IVr+IO
sWzfPId6Ed+fHXEm64mTIZh0MTorIf2k48bW7s0vI7byiJSy0+41OdmHP5D0YwCzpQYRfzUflVWG
oGdSFPQbaQ0eIsl/vKA8/bhIMeATW1W+w9m6XC3mWuRYK6yVl2TrE1CIrPq3+0P3PKwRpNW7hpcr
zdaRiiD690fNG0SebRZkCNNUeqleMUVu6e5t6gF5L1QVfSUDZi3fEwY3SooDkapbbB6GRrT6g84w
Iesalp9A1DRkd+wor0ZLmH4VR0wFbbMWRsMJxYHRNei48f8cDM6EQ28w8J+v+VPYJPSjHaaOLIvD
LTG2eOi8sTpddH5K2/0/6hbsf/2uy4jHDmftVulJS/UHb3636qPfQMuwJcWMOd544d2eZubTkOkb
GIV0jqNsY5PBXITromfE2dMgBe92rHrHqqzsoZSABDzpO7e/JMBTlLWh96hSXVhXFDOL7WIPrrHd
RBsXsDg7rN/iFOJ9gnKsH2/EsxOlk5D0384RSE/s5DqJkN7sO7w26uO1ya6cfPTNEEbjjJlhrfqB
bOxP9/pV2k3zcK2TryheqF+OgIAvUhZhqWaJkTJ8JbAgkhlwjOAIcja/aCvo5oM3A/7w2Y7gdVD5
ch/R5kbkduu3Tw9qWXV4+7N5esdAyttxEwjv08fZXybHo7wTLLb4dki9qJczzHdJixCpsjalhZp/
xsAYGA2O/oXnimWrgI9hrkbJZ4aPgcxfU4DTWmvt1GHr9iS0mcEKB0hsXnZB/5yUdn8Dhd5wF4Ja
PgyOtqA2WEcucC0j/3eu/luhuxl94Y8Ke61JvVwzF13X6qNbi19ImiYSZS3m5rjW9b9iKwZfFN31
tk7UwExQ/lwiwYuHeLQTNFZCUG+sfMi24YJ2/qWx42rD3YaZnP+hqTNDQWugkDrVFf+hnXiPc/MR
wQLjuCxPQYgOg3XI1pth+CS7cRyHBeYci81kl4WgN84S9xIUrbZj3CSrzIuma/cn+JvzLlDS6Q6E
irrmAzRWPHCs4C3LzOldJ7IuzaApaJZvScVvUKCD84IkGNyUnDBmWZehyrxzb8PWsxsScgXb10/B
FAQzQicYf7IzaL1deTkykOeEQNhDGhq8Oq4N5nn1Wx0cGpMoBZxT7aV19yElrY+O2EvLAUdJXLR8
8a2bXbBfvzz6KjD62YiYmSeQ++Vqs0nJ0AILoUWkFCKJyDY8j2D+s1WWLFH34J5OHbN8dkK9fnta
vnFd5wSbZivpobR/aYWvUF/SSR5HAQW1hLZ9qrMA1PKClsjglk79emCBrodi4U1HukCr1S007+eu
koUt/+kz0Z7UDsSjF1j7C2oGx/7No/SKTcCU5oxZ9rBehGl4vKPUBAAqiIej9rbBHZgtmoHYSxIr
tC8F/Fk1QzcB3mlTd/Bq9cQhtWqOYZmJThbAlEUTgq3BeXAOhA4qtMYoN/Q1HtJplO9GosHF805Q
ToOxT9jvWLL5kIKKsiEJtV4P/oSVUla4tqds9rEO6XivuLdexxa/X9FybIRY7sneShasO690IIEO
RFPHOuKF3x/6ZZwMEMUbY3UazQ8YTSuqFLn7uLEkPLOofIL6uGVcMKJ9mhJ6wxaPC/zXt+94dLrl
ptgmsUydIrlZGOjJO1am7aMA0N7ucFczjoDnQKvcVr8gnfmZWId1mSiQ2cbVn6SNEKUk0c6+DmKe
RoQRiIKFkI+7p1YjM7cIlsMLBTuxkXQsyycYnyBzbXXUGJncD1Sb9aIXIeZIZzliggFtOyL41La0
v4FF8g5MoxwYsLH/E5OWy6dYiq+MHpOzTkrkcGkgqYDnY01jCUGjQnl6OVqANE3htgyrHMqmnfrB
M9xj1i8gWNP/VIOoOdVH9iByQ/vGNbpNSRYLT2aSykvIIW0rCY8ogopDhyUoGGgL9qFTtoCyl17R
7tx8UuoFoTyFtZnWBxbK5cr8G5Kl1+djyMk5mqcoyRGRHZFX7CLkmNAt1u+fdDftaxfTlreAjbdT
BpNgLdBQoJ9o+9GBw2Vqs0w16g/ckXpg6WoA4JwwiYKhvrpgoych5h1nvvNlyXH5F6Ay56sUGmHW
MIs7P1FwU4ysfSPa5WsS18kbvbPLjml9GxlgGpf2A+eX+ELRF8wecux5bIKeDhizh7UamrBlwQl3
MDf+OsHpu+dRtc5aduStPn6a9/Byuz1GiUaptTWEkTwGeSi/OHV26qpiotd1qbml/cqzTm07FnTn
dxUs5QLwOaz7MU3NH8LjUZ4C3Tapu+w3Z7UoMB+HHruTZv7mWbQDHJZOpxz4XqQhA43EMmkk3gQK
ZwMFVy6NZeoLp3TI69q1HT0G1Oci1ZJvWIPxd4OGsUsuKFCrbGvMcMkOWHDbVNPDBWWvQTghzW16
s2QVsXLOuLxYoziDIkRLjLogwnoq12kqyz7sNU+4PjIUunFATG/BALVWkqzcseJjgF8+DZRXrlBh
DBaQMzlX9I3j8aZQ5lOs/lKFcaYhqZFIQS+R+k+TryVGfiLGG+sFFUKqCM7HOV1u5+fKWVFvQd3p
1JkVWtF3+LEhe1EVMGSOwLLaL+PpVOBMFTCkm91g13Wnx7z2E+TFIX0sUw3xGu26fplctiBvb4ya
qKRP/euRmhFBRXo12n6mHf0y7jzcLtPIjvezvDcnSN0kEi7JRwDr8V8dS9hSEnd8G5dDL0XtSKTy
dBU3mlIzzfNysv3ijATdD48VkjlD5f9kPlQqe2VLe5gxW7ko4AZhV+usLnSzr+1D8w1MLnKDvilu
9f07q4rMVI5E4VLP8CJdRZL7aij4kiKzKxqmE088/KtWJi1BbCg7Y/HZmnXiNJjOHZVs38ER68Cq
9uJqy9VepDUkrvVSUI+XYkDa9moxl3Wy6LZTL+9q2y/tnITJ7dmaVjdo0OQeIEJHsNs7GXmowYZE
wJHVbzbFm9me4szogoTBO4o/Y7Qha1cIeOcreEoivYR8W3D6bV3yUUITHiFsOzx5ASY/cGVbuzP2
7IKHQOXAT19v/YeuHSw935EZ0sgfAQRoPLFRoNWZU45tPpDqn60VXA8FNyzyZKkXcLlCcVWEYbaq
2jU5uCZiVELQel3/wCPnK9mT6zaj6zcTgj+/2k9mcCmWnOgVEJSs3EHPFo9npY1X6+TbECSbIymj
ChVPDRJGyJhEfLqMgnm2jKyhj8f5NUZI5of+mWPmAENfSXVEZ+jbEWEHwtcWQblR4bF//4A/sHAT
GMDQHZBYHeeAUw7zIN780+YoHGbefo0F973sCbw11oy3hGXNImLuWYJt9b0u7cU7S7RguzjBJiHE
X3TbMJxevIJ5v3gVHBXTlKb8So/TEVpE/137k/zULdmCHgfPYpV8r+RUvLOcM1n8BbiohNG8Kqbi
u2SD2sBLfuWLFAfa9fDHdrEM0M/erCevHTxpUyovYszUbcMbGomnBlVb31gEp4dFTnK3kWRLTsZD
I5bnffzCX85ePaegenLe94O3DOiQ4b+3RGJuQD2Lkq2up9aujQOVQLo0LPyGnnUJ1f/Ey2KjraGf
Qx3DDk/OxgUcFBK0gkXEM0fwEd0B8D1sJg7wpfwKcwYK9bx/quKnSWqwe1TgcTUHF5SXzvT4pD4i
zSkzAj/tm+Gmvll3WCEO4b8ZbReYPDHob6bgq4EPUf1QoNzflfUSgmFSkTq99VZ+VZ8BK5ClSdEX
wSDdTMmmVhy45yFabW/7UwlmBAS34Ro8jxEpOMCNYqcNO3soO+sX2L8lm887iwCZivKXd/YO3uQI
yUKe7IbJtAnpVLhK1TmZ/A3kg94dlww97Rmy/F0FXkR0DhCzm7jaleeTAXZAsD4kr46aeNmpG10u
OzgTbUnRx9gH/E7qat8OVIy7OHIKlVFqWcovwXFfNxEUjz7EvsXQUs/d2FqgRr0w5KqzBa2M4dDl
iu/37xZWjskkAzKt9WX7an3Z7G//p21msBO7w05sd+XK7pU89DCH/n0p/l2WDgbVmIZWzqNpkPnq
ovVcTH+fyU0OcXXigmNdbqfKgz73f+IabqwIXcAm2c29aqTQD31StLe/RgWnUSCcrtnLFCOyLpmR
WTVdmWnrh+myjb9nkypYlBgHQkPLkopInImPQdMaWJs5LbLkpmZceMEqFnABcsgr1gC7aBNSLbxm
Pli2DHaOOw/aMwkVR3tb482Z1H0zA8hcU7o/CXGvJcfPtINXOpW61tue3u+d+8SE9a/GSMmZ7MTP
npWEbFmUNqBee5ynd6nHqeSQrYInpTxOxPHm2K63T6PWtiLchX406SDpFcOD5V391/Om7DuLp7lR
xMJTcJgEtLc9XIouzIaCLAztYhE6fjE0tT2TTXUd4prHuK7STkGrXwXIs7RP03AaIuOZW63asreS
VN6ovMn62F1pl6ta4M8WktOAx59zRjgokFKip/T/Rku59T7z92+KOcZ0VtdH6xutT7/Nmo23oPmo
SYHIo9PVTKNOb+2tYiXZR0wd+ZD1h2V3gMd5FAAMjpttSMEfsvc/DfI/ItkDvfi1pmEKaOV67dV2
6TfB6CQbGc134e2m5+g/Bea/Rqt7taTxPnq487JLX/3jf+mV5WHZIQvqOeDtEHHxE+qkY0UeL1il
aqiF8e0iEdI7nW/ImrB0nhUynPGumHexo8MsapzlOxB/JdU8Bs3jeSYAa0dWrMczf5mUdtfdcaef
Yy38a/R9EDCjBY/VJin0A6cEWmbdMn2pX4IH9AwItPgGTDjURKOMldYArhlT9ZTu168h+iHnSPMx
rwodd8MMO7BIclv0B69q9tzh7B/NKpdo44QVBC5FZaJj3hvNQBeKvKCWU/OTW2bQ4NUoUpXvJ23J
qMb1cvhH04QGAjPs+v1hPme8eL8/jvUuangNafgdT+yr36WYZifeaanr2KHgc7roXhBfqXqjFW9/
A++Bxjf5wxpJufjHi3nbdgNhDIC5jkjtVAnxQi69KlFoDAjP9ZeQZi4QsFWbHA3CwJDP75o6ZtW/
/WTLo8g3LFDUQ0oDklDDBU62QdW4y2t3H9UF4NVvEJPgflq4481+nAwGpcV+/PgJlHBGt9p3mzT1
7J8FmbizQD/O//JTMbCT5YyoSv6jjJqMGlcD/dvPdQkPHTDE8Bg0Bor9kFhbIQ9vo4i7kooKUg7Z
FFRduw2drKkhcJHKWiO7lAYePTFI6MdSfZ54HOyaIJgNVg6MWuLFFgbkDuEwtDat8VGMBtQZwW/a
LqW4cJ9GgCtEfheVds/lXQxEAkF2nAQmn546qCym02YlvGv9psHI0mAxt1JcSFaoyUkGuneYumcY
LNxyH4cvXwsltNe8OCYogPmaw8g0cnxeSpUwnyqjPllYJHkbY8hhE1EUkDDeQMEZlU/4tKx1UoJt
/qryz0qhnX6ULmZak6nQXwgQx44H/wdIhKXv5lKOXfH/FAnIzAsx3FX720t+g+jWEazr2BJH4Fpb
7TTXjUxtsN6nWoa9GHFQUMkfMCwlpMBfm5DZ6fS/W7KVoYRNsccBbkkIBYUDW3WsfN6cc5+x+hjA
osbn1j/dPY4vB5fHvKnjSFIN/rHgT5NiPmeD4iz13Jx9mVv+fRQuuwgD0D/DEOqYmIrcYX5tv4cL
ITyMKx7Rf5bRmmsbi+hiLrWINpDkYF7iwPTy2aZOyYr0kdIKoXhwBqZtTTlLeH8SJdYmVjG4hOT9
QJ5j7fD+WNLsRaKurazXoVwpeFpof8fQ73pCMItfYaCiSD/GcRuNVQ4s/s95bd/xq3w1Y9bJg6/P
L1YSXA10ZLfK9mbpUmgKefDHYA+c0IG0pKteoquwWynDfJg0qgg84I/nluJ6n/ch+FEshN5BLbtq
Z1GBKX7IwX9CGyCzHR8cywvHgUGdR21rkdDLNE4ZuA1SJY0rMrEIPCivGCGkBxXCbBwD4oME+H5A
XtbCxZKPweUunQ1yEF6vtZpgRg7u5jugYmmW2ds7/f8E9hEwArNDbvJIof1kcQ7dfPi3sF9YRTE6
jZzaYRZXSv4fIRAYr55pV+CkYhauwHF2S1x5eJBkdRSQ18FLSTCmCmyb/ldqqX7sb7pbBs5XewCn
GH0FGzPPHyTkZgeMpDlhPk49XMOqleqNuH3Vx6oM3Zbu1fEyJGkm0FMXGRWdb0hr20XUTmXeAleC
f9TAlD4OC0wox2Ktejs27mbyzhgCv2PyG/kP/pQcSJCSgF4XnidNxO3MoxkLO5tSdANIvUNYyQu0
T/Rn+eMmXnPY5hTY1vTPvwY7JToo14JBNukUluncv1MSKJYESL5epOO6ulZTxG6ZGyNZry2dhZpg
BIcMO+g1BK7cbi4mNxlBacBOb5eOPPaEK+MWggJXj5vnta9i/tP7VmBfLDo0rG+8Pe809TS5fLO9
EShS5lUwSj0cK8B8B/Bjo4t+T4RCByDQ0GGJM1d2V0Aaonee3vZ8OBwNixQbdXgVzp2YZsjFjx/c
R3ThMfKsYG65JhtsZb0r7LJu9uI8HHfdVqtvXWJmQCECG6+nueraWRlEBjaZ7IutgJwzox01hU+I
pE2Bcrie2TqoS2cKa5B1ZzlRAW0SMjar4yvaRacnQcQh4TGaDbGa6QE650xZZOPh5f9SEvIwBYHP
VyX383GjodqQ8TDcCdPoYyyMlLkh2btlA2p7q6lbiFL+CQGsSv6DCH3rHe+GnsnnlushuTkLuJXo
641cVDF3GEyXGdhMkQ3sgJA+It9ZjOUsgt5uJXiJZ2GWCjvwKukKPStsT54/iHIIqwwtrf7o196z
moTEQr4PAQfrBVGuZi0Ee9l4CTc65L3RQ9hBtg+YAl5Ho8QqkuahMoiJDiA8tnMVC/WdCd28kmV5
W4KN+Q3Y/9LEAF3p07WM/LNAct1Hx0MGKA96/FAP5LC4RkXDoHu0ZG2xY3OJf2szn+8N6IRXleVD
nU5LIGCu7HS0l5u4erAJ8yxxX1rqio3EQjxpjZSglDIEzoQyI7OUioS225eyCaXjlxQXZXhC0A7L
KX/h9vxCzorfOEElUlBtpq8qr25yl4TG2BXo03f/8NxC6eX+6YQ6K2IEW8boVaMYwG34tgDn+ybE
X9Ki/8701s2n1VZMBHMoHAtM9JU5ej30r1Z564VYDw97NNbLkKo5geovR3kfEXHM6EF+FNVecBWw
ph+wq5vxL4hzXmw4mOjoYDedK6TyPorGZI+103iBFhWp+aw3qTlMtliph2fo2C6XqooFanNxcPXr
5nRkw3o5zLbWkw+h6aR8Xh+fix6PDBeC/H4nRgjWmO29HrpqApT6lQkGzIzyx6uzdPMawlYUzfls
Y/paqkp9aFoZ5em4F96CIh7PeGla4D/4GMAfxr9T7QRNYoKZn/11cOCayYUNjEuLt8PJ6zYQ87ZW
O7q1w80yi5qQGqiIJw3Nr294/4Ygjfn910o+yVMuG6XJxw1cVCCXkwPM5N+CQ0Je3yvccEH6dWbd
DwnEioLqhobgegdHXHxYzL0JiK2Dj/tkK7Bz1aIxpmGad4+41G3uYxe87imeIJ5e4pO7hrkUYUQ3
6pDU1rwPJ5fXH66jXolk0EPBk933ijyaS1UUrjXs7CmTlQd6ZGLQuyLMrl2DDOcsYs7/O40/MGi/
qY+uTIMkjpMEhmW1AhUCX7PmgufGJEpjqjsiMHMAnvHbCGjK0WyU9eStn1ixElUypZbIIYaydotc
OqXdjIO4DovbdUAFvaHNfDCluFVjLnOvcO9wmI5+CJXBgdwuFzLpJaID5D+IvMiq/Axqf2uYpqkY
mqNpdi9hFptVhIi454qq7gOZpylG3m8+dGHg9SJq44u8BemPQc7riSOd9lDPjUYfTt92PU/kdvRy
OlQF+cGBZHYzub384LJSEzFxEwcj8hlOBb1Vki4PdnPknt+ogYGf/bvVhb3nXYZYpiQ30l5fnJCM
1SU2UWWm63edr4W3WJVTUCJRNYW3Z5c+1bxHHftu0PIOItUQ0VcHYdtkQLAEesrQdFGF7UqKKv8p
K/6RWOwZ9bhBCsVRRQ/9Ae2drdHsZuRx+RaZ3yk8yItNYVMLCNbHU6SUpKJciLss74B8pwzDp8h9
lm/4iQkXG6CN93xsDlJ46hHx7Kpn2kr1rxqXF7H3xlKVd31sdbsDgYkZy6Yej1C9ZhFmXjoFCGPf
lMlfT+2ERqqhupcS2MshiTmcsHLqyjakDzeIedFS7CTLlcGRHz9xOegBRkQyq+IS8jtcMowVtQy4
3DOBwCaihfokEWbn2xnZsf3raP6WB5RUs7Zsoa9KXUkL3//D1NlnODBtJN8zDY9jSdnC8Vq42upu
wc2wtttsIjqi3gbn5Nj6dQjFYNhaVGweNMNTfTWdvRWgQyNBKOzGefn2n7o0bEyoU0wd5q7Y2gPx
PGPiHHJpymKEd6HE8QbbjZFou4e4jZqwgsQB5yCZuVXdDccEdPYg+z4L/HyxzwHjvYlZrPVhGamX
W3Q+Ungg5bjE2bsX3A9at2NW/a12/3lTUO+KULRSW8RAg3EvfxfFVWAIqpmTOsxTm//2pv9QOhbH
eMArjQELLsOffu98I1HPJ+0xrxAwYpJF4HkNiiz8HCDf3STB8A0VwvkizxIR6FFsZqHOiRpRnf5W
GvSZ0ynzWgwz8yrqaAxX6hMyapu84nTQlNM9FqhT5PZ9CA3+tibRAZB//7HvzuntGVvsh9F1isCd
+Tm+bns+t37tB60/ON3XgDeu6yom1oEy+DDEhii7yTZV7b6/XvDLpaVCd5L7HGmZDaC+ZfMIWzqp
cqZOAakF3vRXivXBiA3T7G2mKFiRrQR2oIqqCVpCA0UwPZiJL4nXuE/J1gv5zXS7smLUan9LV8dx
Cly6vAyOVSmBf6KCjcqQwe+8Onr43PyTAo3KjN60Iy9/usySk4XIJCL9AMnnhJAAsfBR1k0fm26y
0dgk28ip1udVfU7+j+EWSKbyT6HwMfwErqlo2uoaBbvfFSGa2seffJI/C+SV8F1Qgprmon4Xt+Zc
S1F5HFvrrnleA9pUCPh3DZrXofDKrqBhOYaYwc4RdybugdM5CC8TGtQtWwXkeajaf5eNcQp4l/kC
qfnhoabDwqe9lWkdn04THvGnR7I9kEZZcQKDeCcFBluHtmeNH5SEfRL62Tt404U7Zsi+R10+HkXt
VophANNiFFEhdAa78c/SoZA9rdlUoXUFsBaxeU+MUjfk9KU7WvWNxk94iZvgVQJ1D7SiiXO5X4d0
ucGo+LsJOqfP70HP2F+IBGQTI0BGktPnGhzbe1QpNVOAcBxKV81hjQ2+QGh03Ht8ABrngT4xadZP
oaQOOjwn7fsNiW+Q5VRtVBPPsR6CFBFXMXwovhrrHp4SumpPMrK1XxaRNkdWSBxyi58ixGr1Sl1g
EvAsr0u4OMsP94Nvxfd8n/TIYNn50zDel460imUF0pu4pa26n9mqLEqtm2dOuJ5dco+JnE7xFBS2
SqkpnkKp8j2XW6Idc9Owwr13HhMvLcuOviwqNib7BCIP3Bd2tyi1fwiXIHz81n6aNW5hyMJqyMnw
TpqVD6SiVzEOP4eJKGOUGtbFsFMZdtCJnP5m7Pw6kzWlgHdTiQYoXh/SzL4be11BETp/OpOK+oSU
MR7KNWD8reAP3thg9sGI18Rcdm6YKUDPdguq7bXzZk+756+rADLB8or6CJqdTn4yqZOeX9Y56n03
fISrg6Uco7tD+wLGIlm3T2IqpbJofpLa03ukJnZR2+NHwnbR0dyve0XPsKemKHFHjxDcoBuycB6X
jc+3uQN0MzQn55f/JBhEkUZOBxhP+P7PjAKdt5vsC1xrQFPGSw09YZQmvCfEfk63MOxFyO5MbPcL
jLJe2bXLtqIB0xod2G3h4BKcai3aMP+ODpR1sCEVsC+yBZK0Z1X/LcX0L263D+yY1MQzcWAV4t+K
HlARBvORfPUX9xVmfEqJfMt+jFBHHMVx3RFmeidECvLTpn6UqXtnCdCBgJ9r+Oau7WS8h93hHirv
RlYixIX+jGq9eQVUdUFbHyWoHQfnlMGzgeTQtR4rxqM6vCHLz1KTZZ3KnrFZVQtpAHpOGyJvROUR
zVmPleNVM8HFcWftI4S+9X1+PaxaxSxH0uoutfbPqwMh3b/A0Za7rSV0WrnkKZiJVLTqxVpOo4f9
xA2aIc4RBdKPer+THue2ZAt3Gu/P1Wo/P8k2T4IVQU/OH+6wlss/IEmsMzcB9c3b4gu/wLoFYldW
aoG+2bY9XpgYo4aqS+1AXcMAb4AcNAvadqXpt8ha8uffTv1EbRNez4cq/scTXMpXKpnyto5/79/B
w+cjpELC8dP9azM96cpc07Gzh2EiI/kmlBu5CLLZsuSksS3/Bxz7Qpc9PXVBwgiOa3cX1MEJvuuz
ak1sYH+M8+Bq06u0CNY3IcNYu6HDtNJV7hzYrMntt8498gGaQAJvn1n0+ezI63hy5hfH25v7PPFz
BixwMIccTcCrPatBj6SJPMnclsBH1Mtd1l2odP4XRGF6hlO1je+D6JK5cNKyC7XBAjSjqbODGVE3
rd67qbhJtV3B7H7whWfrS88pAE3BC5hvphcoyLfkXvaZJEu5uMbMd5SL/iDSGYHWNYBmLJpq19yu
x6ZqJyREmW1ik/g0Wpuv8zLBjyfnTlnqFNCJ/fLadq713yS+z0khP1NK3RSWXniv8zG3w4svtINS
4YIg1H+RtqHTFLctpdZk8h2jQfHsy05WgzNJKVA2ldF6FqBqQp7mwvMwDO890zYnNZoePVMLkUNs
2iAVF3bestETE/CDP9E+klnjv1fLxlxC7hJ9Doeu3LPmnhJ3HTFFbklamsDDlC4YYAqbXllra8l5
/C2OsOlSC78Spgqsvv5J+Gc0CEy3WZ0KPsquWpeLT+YzC3yN68zA9yqAR02m+2BdCMSHD3E0X+bb
o11AKkGnyvnI2R0z1Hg5Pg4eRNLkSnCU3f9XdNYkXy8uI7urRnhjyyHn4eABXRDA1asavP7eE2Jx
ymbqweEz66JvAupoHVet0gQYhq/r98FWN6J6VWjmWGvsSFjKQJyXVY54wYgb1C56algF/v5R3P1a
ln5rjUS6KgsKw257WKszS8HckiMTQArznXfi4ypsWc4FZJjGxJ9yvXiJt8AlLZawx/fYojwYL2UP
H95SrTiBJ51qTnb8DJvp4niauiRo2h9AhRGaGyPE6in+ljVcNuOnatUj5XT+flro2CyH9B1cln7m
HpEVuE6Gt6rZ43f9Z4HNVjQMDqUyNUji8DixwQyUZuPOrvY4Jf4hsHxAhzAPi5uxnF9wH/4FlN+K
iWrWyvZw1pjYO/99yhax59rWP/0zf90mvuNFCVIzr9SgPFgitc+kH7gUVXQWpugHQbbGCsVX0qwx
4BnrH9YU22hN2ORZWmal0xo7t7rpE7yKByJ5GL5+TysQ2s46bfxYhOL22EcE3n67Mympi/BDzU8V
ppo3NP3uAVIzFrWFr/TTZzYQQehCJBwnKPqIKxKHCIIb4G+Jorf7MM4FgIb5HXKUhl1mLgO4uSvN
BUKuxBaEuEUZqTGbEmJPdjGiuOeTVmItrITgXtCSk3EpGfvRYsx3BOyOYseaOGLGhDUaofNtQkdT
RJm7MpIJSwFoeimUumLnyC7Yq3nnyzYBE2Jjfjp1ALe6J8XyfCgzryBqRFDABl/vnDTuVbfAtB3n
WLXRNDkKw0+oiBknIAmVS6j7VIIl7AGMHsDxoX922zJEvmeu85bbs/Fn4zMGsAiFdfrMEsuc2xO+
ohVBCvv9uI0yblsfS02ARDfu9EgmZBmD1bL+LLyfbto7AuTUM+bU6Jg70Dwe5Mn9JGg0fLmynAnc
V+vGY5j3gH/4KRsf/Kv+coTOS5nhV5YJggwbx+AJs8s2tVuQsqC89ql9h8ZfF5WpzUaoXKs/0WJV
h+ejGIo88pcarXIR+6CqehPx8sDdruH/tqHaMUFAd/KZ/ADvaCq+UoREax0BNdB9ZYmdnprm0h63
b386nliq6fPmkEA/Zd1CHsgyiYm5YC8OC0kBLnBP7AH10sULspTWmg4Mw4v1EyUdGHkkCJppx5+k
6ZVzStRPSmxQ9kP70VHjw42Or/z5G++DutXXzT4BOFpBQkyuZuNlukkVaThuc5BUsw7vj/HlwzR7
Tk6bUNlHhzrtxd54go3JGYI0RBh+Zzh6Tfu23Xmc4bCujWUghQbjEY6J41UN2hl6AsNevjL58jIt
LQx8LQLzJugRTLWogBoF25qviqHCX7Gz/7Lp9lzO1N9+CuGvt1Oj7kkPzv3VbtrSPwUKjiAVeYFi
cHgKRcKBC5Y7k6j+3uvsMLc9qXDRioQsoQr9qo8cA9NZYLl2ABM9TIWQDGF1wwJl45+8Il+72iDo
QkTD8Roqi3b7eBbE2xSzpdVmqHv/prs2+uysPAR5n1f/V37nV6tAZeCmWUfFbNQ2z7bV51JX9HcS
/oynTzgkpO9iw5NkI2YXDgmxZqF4ueYPSW1NW8eL9O+7t9o5CErqdB4FwKkr2s5ajraB0ujlgVqc
jF+PWVdVdzG6Tjmg2wrF/t4zv3t+m/xPmi+YNBrDcNmzD86hQQpN/liqMW8YUt1RfWRP1EsBKxmj
6ZWnG3eiXSEweu9SWSkr7IAE7d3QRCWwrBh1/a7t4P1ioHpfxGliHzDyS1uflGkFKceXQy9f9XWX
HRhqjt44GlYPNtXTRFTbpvg3yA6Xxc/q7HPV224fdXVK/5nI2mp+TlRZQmSOCol6yngxlKmbxrCj
YvK3ZJeSQNvph1FIhpI5JzMU+snWJg4Ng8pMA3kwzbTS5LfIq1v+dPgxu8wQCfit1mt1z6KqzKk7
Ro7avyc1tSJUgk/Bsmn+AzbSCyTGX7JdWbY7mQad6O9IfCVvt5m7dpB0+zeEoXNDRH5YY8VDfD+v
LAkGEKAlWytytbedripLCsONGrATDLYQaowZ07AYwOHYIQK9a+vnm36jhURF9v4fW0bV+QCbfCSd
e7XFSa3HsUq/tEHZ0oXaYhEc5E+0CSpcCKLSuG9VXp4KftbfF7o0GXljrc9yWcF4VyhlVaxsfaGj
adt1p8ZJ/Cpp5NcuyKzWxcwKMEHPY1NIW1uuHKQo+xbCwXevUim6oO2LIi8wj7heYZ5A4Fz0h7rW
IlipzWxb4tBeJiVFX4Lk1eyUzjXGiVYoB8zw84+ZnaipVdPVrxTycjhooPF041a509DM4LoYmCEY
9OITtu8q4KJgfUJjhTgJjy2tccBGDJqCMN0T1LmfId3ejUFtharXMOb/pcU0O3kjuu/O1i8uDYzL
4724SkJhevqRr+/KgrMGcy3UamIsqht7Laiu9g+E+pWrInyMJdNniDoE1bRpN1rgF75Iui+q7Ru+
g8yOtBYheESFQmgeKyjyF9K3lag1LaDGGA9RItWx73qNRZZc8vuId8biqKlUwXZkl/EnUdZUJzdj
RLCkWo1zrZFEUnovKdjwUn9/mDfaVN7ubMrpjnhylkNVPdmpKAACsyjuie7rFTLcVU8ZVqwDE98A
cy/v0OG1/uMwTzJcw1YslW8ULYZp7oUP9MLTbD9pcXXU5LD3MqsRkaceP9GrrUoUgRO4OlrdCDJY
TzAjEtP+NfR/cOg/Dek3HWpCSiQbB0ybU6CwKSALtUuNKu5mh9+wrXFUgMANpTkt9e2Gfj52jm4s
uk7BK3xkrSptiWiVsNispnt1MuGxw6f9PS456asN295/WuyuMKofUsTQ9OVa/wdrq8jVGxFI8H6l
2GR7KP0B2nPFv80ffyNLh86e2sx/h9fGM73zGY4Pc8yBMczPdDGQBFJsgOb/oxf0BB1O12FUmOzn
O5wB+y/E33xzYQVqHdPVS2m9jKJ9X5wvf4/BvU+D8fPAMa9umXIsR3mWpgHuI5X1OEV78eYj5vYW
YijgAmoVFqyPMY24RzK+UpjG4N3wFvCq2Lnl8AeI5H60AR9HnvvlHnS0KkoKGoufz8dENcFhF9pJ
55pCccmN6aKSnd8YUDycEo/vf/QHAkbjjWl6rNVS3+PgXzOvkJk7OcBci4RGVuZkoC0j5fW7BISW
Q7A/C/0lGFzFyVQ6qGAMbxkkaq9ZD3JzIXVEriwxYNupu/hHAj4IpqM+xQzmuReepYKf5/gM4spE
kajPtn1TN/bXL0twwLIxHk+2bqWtka/VRNPVVv1piWCdyRzEkFIwsCnGwv1HzKyG+1/rjqx6RRxD
/pBI/J1lO9nFk3pPPjjSYXasJPOXzfUzFRPR5ic5c6yg67u2jgNB/yu1E/H5rmhSlKVCEurvVYtV
9e/oYzuQ4eM7N93XJrpXdzuKY9olXIK09s9qVZiHMQUFn89TBOPs/pmy7MEkMS4ets/2OHqXWv54
jmcBe16Q/dkPyx2n2K7YEOI6QpdyrHNm3o63hO/XjToqB9UW1eVJwW+ntr0zGeqDsJnvt6DLIILu
Yvq83d1pz4nDrXd4zaaW9FAZwbMe85n2TGJ2H7maL1ZSKiEg3pMxsu3XPdhM3kQdjRpQfUXeYCc/
AjYcUjEn8v89KsSKa3c+WYVkZX6BA6a5rzGofmMDbvpuXUYpPMxLi4C/AO0PH4vUs0DMy/++00C3
Al1Xn6ziJ1DOC3PebjVuY57a5QPlggtFh8pzQdFB306cFKCBT5nZui2PYV79t0U4VzhiK6dbmmv0
nzUsy8qlE8yxjF/KhYO5zIAQ+pmtpOpWPJ8ZWgBciEVa7ZphmxjqloCOTc0o393WJvdNfVFupjIB
Kh+E5ln+vRumh7ovjAmY2Wa8AbzrpxvsHHdvLmE2S/fU5yUM4ObXnhUpiTX0opBE+ukqErTpvRJ2
CszeOb9suWU4WL4fDnJNxya/QDAgaHmJptvUPCIwAtZqZaW/gW7THaS1ELCs6B9Oz9tATtU5i2De
OoD8IxhfC0FR9VLh5QjREnsUlHpTMyx3iGZUBH1V+SsL2YY7mkxtP4xwU/06RtTsezUlQzYwMtdz
mAQ3wY9MZglIxi+u3dWjvo/5qFPvdYiAZE2P/zN6RgWPQPPnxtPOrj19sbEU7VnOwwHOxsLc3bjc
doZQscRcYfOQAmjl+xKUWQ6GRT3pl5pPyWpPFwAnfcGH/BCTvE8sd0F2r6qpCANGgEsbGEwgtHzs
teW+FWXw11xPvHWhyjDGSa7RDJd1p33NUZRMiO3R1jq1WOyraiLSSWuBSkyuDrE10BuK4tEuQS04
YyX1gzew1/cXJ5cTO3/Diq8zZbivfq59B71FcT1cGE6dz1htnwvb3wnmnzFMvv/IpKFzNx8z/v0T
HtEL4mtDNjSZ9begplRJqxakZ7dVptcRBkDq4eY0GGqCdzpHBH+yiUhSltMoBXELUVafehyEsnZe
rCgwn8nmKBqYxzRGKKRUR0tTKAk99CsZc8fdZl7KImMSjY1tJ74/VnAmMT7mAxf3N4mNTCXEyLsh
Jm9KW4ClKzL65cXjiY/i1yMyAlOKz0JBu7CM6Mugj01r0iFiON8f3C1TRx7RWdVB2Gno+7zoXUor
rlm1ybVfUjdr4aCZKwII7CKNfR6Qd9n/0SSwjKNsOMF0HQMdKleGBV+8vYYYpsiYKhkVF8SLcsqV
CPBNTe//3JCf1ZOyz27+PQCrdA9fG4T8oC9UgCuywkf83Vr6lF2/S29DEzKdB4cwJFawbJZMimZa
7/QMOMUwkLjUsF49Fz8DCL6XDfCzukL5iyBovuLTpUKXkPPeIFHwBZ0hB2AWTT7xyuWmVIMe3wuy
K+O70Y6JTnmE4nBP8g0AhdCv+NLv7Ud53mQcKemRyShFN2/3l+YxXUtobOYGC4KewiQh5TvLfwsQ
LkMzQ7xab/oN0XaceoGYjV+CKPxfmM+FAYi0axPVimotgAF4pCN0l3/MoCY95N4uj+NG0bVw2KAs
z9EcIZLW184GCDM1SPwY+e0EADcOoqvrVOzsegpzd7pjOYkWB/2o0FKq0D6QcADdRIuIR6pdG/I7
zgAVXwfeCl7eWvQqJDMhx3RWl/KB3aWLqmrl974KlUcr+eqJCLB1C2CTiJURZ2/d8YsQmc+YGwop
N12neNtoELy3zyLJR992FjPpE7I6+Ez6ANKBRYMB1+Vo0Uj5Qqfk1lmm+uWjyLZV2eMcbp56WZPU
PO3ZcTdjjqZnjr0Skv9uHOgzII/mi6JP89T5Kl0CEuHnQ1GcFGrfQJqX9E34I6IimutuW2h9u6Xw
QdDva2iA4yZdt5Tg2043VwvJXG8kqqtp1EkgIWSmSQ8XZ7wMCcuWJ8YCLzB1dnwjMehgDJDTqXqq
Uo/bse+KzawVXck+1NZhzUlhjYkFs6OsnFYKudESKP2BErGkh+yk24k4Ltu7z5WuVwZECrWsC4QZ
iM5JHa362UN+mHDWlSSLEu6aUG2xG/oWUTMdRqHoTsAF8TDmDBFPD8kkDgs8MMFuSVbcQljf2mjF
VOQvt0opR1TpaEOA/3VRGnCTdie8NpKTcWciaQIBQm2nZgPSrA8ucmKI2kZEqV8QDfy0wOF0h9i3
jObIsn05qXkZqcIxdMxAbz122kw0k/fHWvV8b+G8JXwJPcAW6inKWBef2xvN9Cnv6OqGvQs7UYIH
WHuj3vOvz1PH3/8eDs4g5rYPOXp2Nh4Gihq79UhOeb/haDzl7y0+zqj1mDw2ULPSDhNxTrkmjnhf
7gLqxcJJ1dQwj9y2YiCEU0qK9F+QfcrOlsJELecmlpM4weqp9sywC/hX3Wd4erSJfUX+BOXaopX/
nLhtTKbNpoxvcBaMEULKdc9X24v6a47InGDOITiqTajRvak4pIF69+zU9+zfr6kTu/9SEg33InjW
U3mXxvWTb/u9WJTpElb8VlB8jDljf3QW5tpLLfD/kYqtjXD4MdqxR8rgA16ed7ySyPqwN7e3EJBz
8YpWryISTANo3tDxd4ZKfyoyhJaA7RbqbTWspNhOypJQzJncy79jfnrhVB/uGsedVBXlJpPrNtQW
TKvVIxvn2JW9boHxCpoQhpZDqkOo+Wn8ALwyrBQk8VHdZ8YS3UkzhCWIWhcNTl2qJA2ospd9Hrsk
gdyyoWaRQNiyAEeTSqpPtZms+dDQUuhfYOqACMRdQveCNqQMjgsfBshJ0+dxF9hDJmroDwXa+uLX
AajIzoJ2IeEZB/0sHCSjdqVWGMy970ssgeFJK5F73dkyOrdvAmgdXpwYdv+Cyi/wkXLX/x0x9IuE
5KeD4Wd87HCV8betc1flRvC8s3N8MaIMLeDOsNEePBJQ7CBmKm2iKG7PbfGOxDTfTK3+3P/xYUvJ
ysHsnIXRspuI752h19QpmuP2Zr58luzPCUqpzKw7fPbx7W2HQ8oGGzqCVDMEErzeyfFZwRlFsPwD
z30IlEjMMN/gh/WMCwdLwyfh+Ic0xCcvOlQ96RgawV1xOmEo4jHCPgCK6XhzqE8Njg3xipywqa9a
EUZ4ZIvx40luAio0zu9cYELfNmiqkBbeKvAwUsUFXRvFm1NcH95PISFlmaUIvlKorqmaPjbqM1Jp
7m62SEPv22IouYnjPdHOHra8pHtoGRlLxRyw4B2UE6iatxo3sgMu+sp+jjbQtZa/r4BVu2UXyuDJ
NJMeZSRwPajO43UaBzsSGWIPlFZIkQ8Wy5BqLVu/6mis1It0sWR51TQOgoYLMwv2B9ht44kMcQ4B
GLsgah0HxpZtYpncrbUFn9OqjO0+kp/IQlKRiw5ZXJsTDhz2x8sIOq/iJA6BzSgoNy9LNWz2Yeol
Z2jQaZs/O6+ivW35s0DhYESVwuPi7lo1fzKAdPpVNfKV/qPvFvmznWpEckiQaPLxnF/pgf+L6lDE
HAYG7b2qw9OP93M+r50QVUn+JQ0Gtg2a8xoOCAusNkFsS4WhtyhMYZ5vKoNknm06DCdbeQfrYmq8
k7JEm2KkDzbkOB0c2yTqqtF7o+OcJ8vBhbZh5C4ER6Q7Rb93YiqsIyAg/v4ELI/ilXX2WS/px2Hv
PLW3Ggd/btZSgJw4V4opwrNDS00l+VkE9TFvFEWe0yM8N9kljdRQSUTFvkKqmQaryd0HptjI6PA5
JpOccPF+AswlEFAVhklv0sXrkJbbStvTOWD0gaLoyd+Xfb8hDL3n7/cAO52MR6p3fAyNEViVWcvp
ZgxEEOE45F9UMzRdETjSlQzvRpgbVsQAbEiyT2z7Bq6wmPcHVvIJQTe1cHo+a5cysFO03EocA2UR
t/S29OZzsvzrCoA+sY3JTHbHXfl71uEDhxnIEVqhq/qMV5p0GzHMCgd9Av414TRMzNsPXTDuxQJ4
IRZNtvb2dJpXg3qyF0OU4lxTvplv0D+GK4YCy/S8mv1IPHVKKru1WG1pUK3vV1uON50PNMrtyw3E
fRJvmVEuEHtr005DNuP3qsjoVeUdcg7IEDC20s8Mfc/2uNH05+ERasE0B9VSt2KQBKxgpNLTLbrQ
mqGfuyoU5wty1hD9A7YG5qZLayzm7liVNzEEPXYaDa8fu+10lXG3tm1xZbkhuiSqIvNqEB3UoLX3
xuHlAq2shkyivoOhSZhKQglyO/h+yjtZtMS/n9YGCogWf787lcy5ozftmJe/bXWCgpo+CBkR8yoM
f/FoJqEEwF68s7Qwl20SCF9lz/LIN90OHScvHI/0FhwdrKshQ5hKzINID/ML3I4hW1vQhqY7eR4f
PfGBhrZ9yVv3SCCTLk+tdD+4zutsIyDJ8y6SpB6U23Ylnu2KE3HSk153ZuY9Nr0dxBYKyPYJ6Q9I
W75Ijxj+wlb/3DDPRGftL5fBOcG9C3bB9kznugzjVpCKW9ex/Cn6oIBWkp4TbRaWDW982s8rFQeK
eXA82u4X9FhCU5xTRqje+QBHeivUlJAoFqlWzt6vxTP+JMJRmFEmAFMYPkktBLg93hPAd91owQp4
177yxvO2CbUixtZtnIP3QKTEN7dOwUVAhPXtSoxmGgK4ROdx5QnIS9hOYCSwRIyBzQao20jOLl/a
1IusH/kAsCm+LP94oN3Lgge/I44mQccf9VTD8kN4co5mqdRkf/lO+ANJUgm6i3hcajV0lyRP4zR/
NH6EnGg/ziI8Cs0tVSCyrp8G+I4XD7SmKSSsak3whflOBHEjDHfsD9Kybt9gXM4iodx9yvnDPdJ2
nVPnGQPTGfyD3gGkNa63drVBjfmbLzP1+qoSTKqEYsbWp+9XXtRJN56mV1ISSANw4KDDm73deSSd
g8e5BIl6R5RkBOAtsRKBsy3c59vbPCOe8g54ULZ0lInRiyq9q/EGulocxS+dNyMLKdUz+sW1UdFH
/polCV6ip7ZPCmoUXTXgrbzGUzwmPLSL3ovdl5UPwyFnXJ/Bb9SHo2Af6PR1UYFGHd7J3f4F2NhM
wCbKJa7c2bah/8GnRRyvERJYDracy2Ax8PRtwP9jRn9MNdgDmDGJi3TrxQmq1wOSSax7WVe4mep9
Y6FKmqbEPRMLpzl3yZlQlCu99DqoE2iri13pxX5yiXEwYiD0Agp3DIrDmR1kTIIEWv7exyU9Lfqs
0lMpINOIQeHgFs9XLwV7LgF3jY/pTgz5LYCA9VY3NpFN01Pp6Vk1V51J9u7Uc0vlEz1foN5gHtzU
Nlx4O0UfHldeitIRGUvYSC9fhS7E1F8/We6rOE3GOKMj7UJ0gFsJCFe+NYA+dv6dbj4lij3D1s6K
qim2q9R9U4As/BijbNQRLtMptiESBpAZAJ48sz4yGRUfhYz5vWmV/HeRf0MZemaTcAgyVohuBMFN
rjEqAfbGZNihFEsAj/fiN/gSR3J37DLpgaxd9pjFbvfHs0C6sL68zCb4zunV6hP3+KOWjiIM5Ugq
sHXQ3fJOYJTXk1uTq7tCGywCT/pEInGVZ35xaaqTmZ6NqBXn87j+v3VmNcB87pVWKNKV9ujC4t2M
KFAqFbo4ydACakZ9ZNLovkOg+xrJ8lzYKWUDuueya7PUSnzpWrn0jSTd351zflKEbGNVRr8M8NQI
Oxd3vcYbPkUHoaKOcZEEHsWjHP08XFHqwrzTpWwEplj253braKaWo5XuJ80pe2oTuI+1dehMZp2R
+uKUgThBHPWPhb4ydwPMiYqYhXHwlPVekS6eyw2tM3ymRetxRKiNZryaSVHOYBNlmp+7HZ88kZYh
O4gw1tNnexZdrg8LnDG4ZTBIiAWhRwkE2rM36LQy69+7z/UZMv1ESzTCihLfJZgkq8fPvnpB7z5h
4T2rccQTRrg6l9xFxcVfQzP/jaz1qzN3vlOP2tKcj5zG/k47cTMxeJRcwBjXPiCOc3MjT6D9gZtP
4ye2CMkyBtzCR1q0CssYE8CcAj7guuV7CwMvuieEEQWkXJsI2ucmQq1c9yTAFmPqK9LkShs5f5EA
qA22cbcrRpbzy6crIJ6S1lpJgZ7J8ddoPkUUq8rA6myi6EpAKNczjnClPYfwYHP0erL++ZvkOO/w
SmaBcNS9/q6MWpUt5jxjxTFDM6D5nvUFbRWt1Zk2XTgdmn+vgLBVpUrPmtmcNpsT0F6uBNMliz4w
Onfr1BQmYwN+pMJt6EB6JelsJp0yOBhCjEbmI0rv19dZMtMhyEnSaejG8K2x7JSg3Y+YqS2aLiYR
ILwfNzRKfTjQQSUHhgisrTCEhWIWdwzEIQ210hv30Xz02l/mVp6WfVSV5Kd8fdhhmnusf8gJKMK4
dMKbff53K22wSId8h0HZX+dAt9VMHbjjGSEliGlMHg30snbu8z+pFIUg+jRoorlDEdKW1B5fXNPz
/h1zRWXvM2MbFK2JVpjuP/Y2JniwV63VnepkFhBdJYb/6KxGoEa2C6Ns4Xn0+n0Koh1r1jkzhE1z
kMz1Cw7/j8eLFryhKZnIHNuZQUPSzWeSk8ST0hMCpZf3J7So+qmkpG6bsbAbQ+fdOJ+PkLSeIQLf
skElba5OdpepXpX+A4e43MEGflcFrrAmLN82nUQi7KpiD09B1cSbPpkvQuT4NFfPV2tcTi9Kb0U6
JeuGf7q042vGK7ZbqgcYetfi/97Qto+oltvIZBUXu4+THxjc7fwinyXh64BQrzormVvOF8i118hp
33ND2JQM7qvXcwYmH+osNKNHKQbJh23GRiQBitUyUrjyiY/jjvcbrIvAhqVp6e4q9i0nkHt8ucuu
/E0jSXuY8xUWhLE41gz1BFTYisI+pxhV7ZDoSlXJ2B9eIj5qAF+6pQG5IVnK2eBLS7Bzj4bJqmyr
OCxfuiOG9vHgPjSsMEpt2k8VujIl+ju1hTg16xhHTFspPmy/4N43CNO3G9rZT/DSSd/kt/7/Wj04
n/6c8oZ9CZnkxi+4iVOp9F4BsjK7wUcS2AzMIPlNQ45SurKhja7ydmRxDEWNSvXMbgK6KHOi6AAE
mQyjoi6C5+o3HZtyggV9y6C2+sK2pm6ygIJdBv/zgcx/Hw9yyfcRo8gR7EJsbwi5quONC+TtfJh8
MPtWkIXO3pmmcIFpqKZLqCsRq3cd2Ga2GRq7PsbbI9/Sf0VPtxX/AJQCKNkj0wIh2yxiQsbE0l9E
7Jx0fDYBck6EHjVfnSOn76LELKDLnz4tCJe/e3+rmduEELGu3MmGSxYa0DtHybRrRCG4sLn+PolO
5aEYTo+4wNv2RQkmbTsqTCI0gOoLUBcknGDy+3Csh6vm68f8TZbDsgSXwJAzXbCdyWIirkpn/a8n
Zq16nMKD7ijBhWiezt8uJpd5CxUDb+ugCO78YO/U1M7jIgWoQgvPU2hXUhY40GKfpJHal5bFg140
Sv36gYzVXicHWjtRnpG4wmpUCbLhDwJ5mXABRXIuXettwIoxDUaWHFhoEhcR+UtYRQtp/T+HyF3z
L/z2+uwDDQwGLiOKfq/01AspAruRcZoopFN+4UKQ+CYW876zgeGN3ev7xfJsjYaYshGDuJQjxANR
3IIuZYeO+5Jf+p0DFmmRpZ8cwe2o915rmXH/jJuHCLUA73QVw3NfZoCRBtTLLnA+BEpTRK5YjWNu
XImkLPsN4oTAVeYKDNiRGcKMjTnomBIxqVXz2FDJf237IZzDpr0IIzvL8OrZ+HcxpJY/D+2nLSlK
kIWlRkh9iq+3h+mniUp1+ismf+rSVxOagqgq6H3rhvJk3MKBCH+r8VKEFJIZ+XXB3q6iFyjDrI03
NSufx2xhVyHPTL9wW+PUdQniCy/zoTh6ii7zbKRnVzXPrIcwjQf7BPQmpZU9frnGB+eW11YJPtcj
cS+r3qyFIoALdsSigZ/4GlVtOtIdG+N21jJa8qd93xjbN/b+idZfWWyjiE98aa8tjJ9/0zGxoZhg
tG3v2J5zZgjou2N0Ue+mdvnSBUiyi09uXjWlTOKEZaHFleb5oz1tNV/oTHRHUFl97tgNMw51Vbdd
vXGIX9TcyFIVoaRYxH0iduJ+VbGtxkCD36Nqey9yGS1OExG8RivGv4Ppn7PVXjYoaikOeYvuQxai
p3AfrDSnRxaFTeQFhAXck7HINq4MGrXv9f1awEJq11c9Q/QePT4PmlMzcTHwQ3UbhG4IK9pelMm1
9kYBu/f1VYONsyDP2t9/YiD9/4bsAHAETeVOr0X92A9Ch1TQyV6o36zoFM77Hrl5G09hgCLzE133
5PUpbG4ay9vk0veAa2ZRaxMxYnl+VJwC3X7T/3KRS71pkrOdpS72wEbwiZwlSYE+aT601m0vERJh
CA7KswcvA3NqeApPMvMY9ivuZZvC5tin5zJnn7kLBgLvSP4uXacv44jpJOjvR+K1lsSxLJ6uguWE
3Lch3h2IAnpV8xz3vVuzjYlUSQvbvmYN7a2WA/Ordyn5FyfknCczPjI5i1+33DPb2MS3BQIs9nl4
75VklikUJIvW8E7arfs+lzX6D3xE3BWP7DK/2cDdbPjQpPTbQSy9cAaaChm86rxvydxHpSRnanAW
zfeV2Ngcgyl+9mgfcfPjSxihlM4soPPOJOfIoakh4ewy+na7AbogATOSYTdDoPne8u07a7Wvz/aT
QGM+INYVtV8YGa3xeMHv0m8bkHkiWVR1TgVJ/kmSrUo5EWwEdmngzj7BILo0vPmEFj0rZVVjWBaF
462Y3+jggu/jScC1rtQqv5qs0grW0gXyaD3F7OquHtdyj+ibMlAlDk0P5pia9NTLU2RI9KxIX7Hx
VmRk+394CD3z6gM5/+zIGhU/1EXlnU2qUO1BiKnoxD/mUxGN+skzySYEynzD0A/D+9A09BEODiJK
Ey+C8YLaHpbSoZoD+dG8VNB0iOTWVX9c1vaAJylgLQxS0uS5Qbai+pj6sF0vgoZYBBH6B5wTq/fb
pvoOZyUbDJX4STNfGAjTnfAoyw23avGaexvAcCmtlFeFfkzwR21K2uaHpf6UAEMCapnX/LOX1ej1
8hMGgVRGjowP3b8ib52ieVf5kfzGJamPw3nk5aINvNyBgX8/7LGYhvxamVjUomvTA1NpM3earw7A
0rXc8K+iajXDfV9BealmPhZd1Mm4oBe5jmx44eUsA5RkdqMgLrDhWvBogtH/wk7tR59npMm6FpFT
ZQYe1NMhs9F3NTMniKaRU6HHzCpH1adg+g1+lXpdoagRDaTCTAco5/I0SoOHTZdeg1BnEShkz2qm
KLr+E252LLZE7jUgne1b8r98oDoIYZkLbxxjTnRfdYbJaj7Eh4EOn80xAz4f86mTSrxRkUa9RIdO
PvK/bUfcU/B/TF93GohofdgdsUuRUlLA3uaLew+01osKjCD2cLlR8OTCI8dnl64x5gxQ8dSDx6jN
PfdvO1oNrOmxtXvN6mDYLgDLGJZprJ433YyLYjNUZM2co0hb1zdTEsZAAeaSmNCA9s1DcO6AGwTo
nBE85wtK892TsP5V2pq/Vpf2Kh067D9cXdLpJb+7p09Hn08ax8etEBRR3On0V7x09J+Vw5QOADIp
/3PSlVW0jXQnracRtWEdZn0gnFqq8QjwPYRpI6Ip/QJmD/nMuwMrsjzWh3pXfm4M24LybporMQ0X
wzjfLWQTBlQV7F0w71UW2ddTSmZPnG5F2IorrYKaqhhOljx1wl5V9r60AX9FuXPcyOYJ8OR0j/58
KsgD51uiSa3r+LPyVI92L0Lg1EerXRWrqQeFLcp/PLAoRtwEc+22+JYv3mM6Xq1nV+qUa4l4zIcM
KkrH7gR0MOBuL0Zacr9hcFuNzFlITj6ikM5GuWCwrlylO9TCsdBaY/7OHjNPV+Agnm2CHNdGsOxG
l4AlGyjaLpMBfylqXRk9qWBpF+gQt1CRtfWzq1YrJd6lS+/Bah2wLVgEl/7CtMgaYm3dnfCcEHTp
ArZEUo0e0xWinHRNqFfW1WcSKBHUYMNHcn5DXopt/QbnR91Wg7pXWtWhvjkxctZFBLr3fWzqYcjs
xk0Tlr9q9zqmhBlfTuKx/7k2Wv1aJ6v+tOuec5guNuqUZng9Z6qWbdP75bQ7I+WRFNoej+zR/auQ
e3RE3JvvPd+gaS8pXS5/PwJhu99rym/fU87I42/9VtPCLKT0UWOO/fwK2Z+uFlDe8Icxh4Rs580g
hiq9v4RTEOa1mcXYJZJg2MzbD2gCEU2nZlh0LfuQyZYkuI8MGUtnvJ+tavvJ/LcCVh/mrVGZvfWE
UbPl+ZtbKQbXgEYHyXLItKygPcLlbWxD0ZqWbaYxIGkee/q//bSma7UszlqdHSTZuUhJdX63vf+u
K7yutcgwxXGr08YG1p8dkVmyIha1DEF3AGJDmIJyv/D+0IzMII2ey78+kz+RxCGt0hjBxx/RNFHj
vK50PdS7KUmhoWmV/sTopBVXj+qZ3X8eb7FIynj8hM+Bn/ftQoq9AU9FB/BMJgSmE2JTFHEQzRfN
hEBQKbeQhHzHiO/4Lr9mG+ipBcv6v1KUStnVEf6wn+E4u5y6VpnlOe9oc5FAQ6OgRO3niJdJbNpj
9qMQfhMpOOAlLb5ArJr++0KkaSwQK0I3Dk3UdHgMGy2W305P81QQdg0LjILty9pnLrcbHom4SOqM
k+6MIDsePVf4niMX2GK+mNA4UtjCGoXHaRHezAGm9Ba1Zj6dPZ2kKIXQwZZX5DKj0fuRh7fBKxSY
Xg26C5QCajdfcEBeojhaJxnhpLaUHvcFGt9Y57EpZMpk/0q+1PjcPOtzO1lPR7Z4YaCp/05uaB8b
Wd2H5zddtAXR94XpnzkwgjdMIcSwLfLn6LwM+znDx9cFf1xwxGGgeqGAc5jt2HgVDfSKFZzNTq/l
jD4HjAjpj3n3aBNnLl3K1u8SzmQtZptLexZMRajjWZObiZpsUkd5pp4w0fsAQlNlmMmJSBeGfAy/
NkQv0XEjFrSYrZbVApdApli0B01meCGnNwDEObRjYsAlRJbWhMXJ1sQshgJQqGusF7IWMGFsgEmb
KcfI5ZcQ4C8VY00z3aWHQsJY/nsO4Kgv8JXXF/ayFu/nfK+cE0L9S/QtvVSSFOD3PJKHuwy6AiKN
PZ626w51IpMXthAjJ7NFGsP6r8h/HQSCW4I144Aw3iTXl2K63Cjk9UYqkspTk9buRqqGpqJepQr7
3FKIf3dxciqgFXQdWIZnxoerF6BxIXt8x0Q+E0ylIax0zBXku6wTcUKMn46yPwgmQzpGxE9C5Bt+
i6jpBK+0c2KDtxZSjjdsCNprHp9Gllc7dXUrqdS7y/KPeKakXAC6Brj+VR+M0GjgJ+TtTE4liqIg
RGe+QtYznQ8pV5hACkQEvO+UHJYOR1z6tCIiVmgsB4ZDElekppD4+HnX06L44mzjLMR4d7+RmcFR
QdELJtAPL6YITCOHUvQBz+cXWQ1YKds/H2mAl/1Jn5hjdDlRPzWOphc0oTkBDIg4+xG2P8v+tIwp
DF4MRzr0eYzp7I2zwhT0l8eLWIlzBJckJ+f44tmwiJXT6TubASC1BuhVdW7PX0yMhL7vjEk2qCTh
oZhxSfJnt6mm7YzrwubN8op/S2WRHSLzCW4639XeqsHxgY3gJ0bLmYnmUiHGSrlDYeJKU1A40nk+
mjQKa8ZhB/i3AAkrymRkxH0Eo0+nqYwJ9fGGnzA2mNOXLxZoC8wekzYpPBCnBl2Kbjw3ctKb0lB8
sOfDXNEx3T58MZs/FfUX1aLxRzJzqyLzghuhboO+SK/Q9P9XX1dYh+P61SVObPiVWWa5q8WvShgs
QV82pq8uWMocEZpjNMzipv7SlTgf9+oRpL+SFiSrtnSVuAsNfOSmTt+30b9KDhGIPvSzwGU4pbGj
itvMDpbXv+1TJ19gtt5yEUrenpajCuTmhf/Mvg9CFkFi2IFurpFlxjpKf5K/zI/r/A+2ui0PpNWB
iiwwfyZaQQkkmLQGTHGuwSWUY2eh3rLaYb4aTSjXn08sOKcVB0FNdH1yZJjzruc4DWTzV2UemORj
rGNq/gwGqD8/r+THwA7JF/TVmgzce2eAx8KouDabQFJSU2qM42zCzw5eIJ57PGy3lWzPxjofxfZ7
S8KU+D2eFd78PayIQUuBXJqzYAjNTPGqUDhfhkcnH7TfKCWfScGx1GjyH96Qdg0CCpb//AW5iiYo
nsALh7dWZOa77bulfoQNGDqedEvnZ8hqIBbBeCBu5Zydqd2TO+8/hNHFvIAgIvynDiTUCvp/kZZs
JN3MIjAgWqw2GY2Gvq/xKaY5h8IPWT4kVg41t9BbVo2DV2kYqPnNHn/ghrLi+2v4UQNrOzndITei
hZy4kSAX++B2eaARSl910gN/wfBbxk5phzmNmTRz4PUhJy3cjqRn6ZC4Z6mxOoXiMl/JoEABoQX/
329qnmk2AyclBKzPn1v8JwIceFMsV4ET5FR8qE9Af/fermYsEKyl0YBvFkFssJEabpARpN3zRbPc
3r4w6UMC9amx6eu4GlVmnJZXyfW0FEQBYmgMjTW15Fo50wXZlAim81M/x9edaVe1WraWsFhxqZDC
V8obgG1P9L2rnTr9fox3Kq1+tInbj6OqvhXGsvewRXaO+JulK/beWxJWXPM1KogzbgZ/p1BHRHHh
E8NgO7SbWJQm0klLklQ1pmc0pNQBYwOuzs8ju27fRuHmuh7VsxKECmHB9aLXgLLX3QW1p0gOwM5M
nKk/jhWl3YS+4/9+2kPEc+jVkR45MUYQNjLv7tsLtrWhPjwELhW5Jl4ODIgaq4yBvSHeCG2LjPxv
63xHK0JyoDgSpzMyWIoYL69Ln9QbiHsPbUvh8UxU249/q5woyzpWnPu6MF5rVUtA3jRd83T6wxOy
VI0Kk0fh5kqGCouT6MjR/EQmMA4a6dJRNcS66nnTE1SUfcSnQoKEbTMiY1KFboeVYZlehOD7Kh1N
kILD3N/9vu5km4WY1s3EM+qCLfTI9yjAIVwZDVuWQIPKs6sI7X4ujCBtuvvNr09pJ6aHoZQBj2ze
H84iSNSDYY46RGPgIltCO3RBuB9qq23/IEKhCscLp8R7Ni+Hk/rIcPxy0ASPSxa+JR95NJ6mMs34
jMLOEELKTOjjM2EqkRLpLC7j4Cxy4ddosalgKM6gks09/3bPEww7FbL9lf1W0JYfPUTtuv4W9f5V
lgsiIGET5gzy1TZpqrV/ImOz8sJe2unUmDrFr1xBfjWr26h2Qe5Eg/MNv852/Rs3a89IjMvZ/L50
TG8SLOF8HuVWlYs6BVI0Wowol0N3SvY3eP31Z7vRygkHrOhlht2ELejFa9Ek9Qo77JSqgkACyVIj
NgPo5fb/Pg+QfCdTZa6lfhnt8t2ijcyNydvVVerXmEUMZobOHZOR5FeSTkBLr7776LAnFTfz0vlS
0+TFfJyTPsa/XzfkRUO1NPVV5yV+MR/MNMdmmrF0ZO8uwIFTUWUQ7bWt+dDIRcN+IfTCXIHv+owF
0xc01UVyOPBv+WZfKjAqEEiZBY76uI3Xn/rfJHCMmKjJMMdiFH1mwov3bcaY2/jazYu6vxj6uj8H
ev4VQPiL8lQfJ0GbTFSGM4g0Tu17//cwTDxt3sLFL0GzUvfJGNF2rP0/fXMpIk77kWbLgzz+3btm
EsadUVdToNU70mLn638Wg0kDcfRQcZJnfbtv7kyaFiwhAQq7Z2sAJjqQ+5Hb246pO0iFlUNJkngH
Hs+I2B6WG7PhfDRurcaw5j+JYMAaKHgFVn8TQokKFix0pf7prH+SFpj0eJscKB8rtQy1Ym4OcSjE
/gGfHF8gxyGclgLiWSLzuInHQPEXteIFykiS5OjH7tB44gAOKjR7C6S+wbGC5OZbNXLQLoEBD4I2
kQsOJN7dAue5pgiASbLvcxwFUNIJePNeaNQTKQddZeBUWOoyz0CST0RSsoA8np/q5APfd3IIHTMV
+V5I4aenpioKcssMyMTCtQ2wlco0uOhSZ+mFJkkxwrKU08baJkgbATCADTF1IM5K/qoBYtcIKzTD
0H00R2k1L2V305b6NAkKsfzRyWuV20Gx+PRI3Og3IAWgtFMRFPOWMtezc1lOmQsnoO1+hWddoONu
lau+eBjEaiHbOnix2NW1aA352WnEXFCF3oo9SK7WlcshK+SoS66Up5ueC6m6TIVNn9Z0OCqLD8rk
phO0pzGHJ8HFQlAjZpj8IlWkGt12UIWOAmpytvNDTkCBq5pNJb81/Gl4FTPvnA+jbflrpzp7WFbV
Bog/RNpDIQeJc7o8fTtH95P6+KONhySGDLzIFxQ5dGtSeQsicVYODDSSyQTbXh9Ub8MHyMAVMjPM
T7ja7CrlTnKZNsM3N2bQx8pUmRUHb7vBnP1fApXr5GCYp9FGuqlKzRg8sFBQp99MnkWA80RqwDoA
nNyAgLQEpFkzSlnJfT7OV7R3VZphN2n75J2xCxlo2TuVCiqX2DGcXzLRziIXLnaXINcU3C6BbxWV
vanljz3eJFUDvtMXqGwKwUVS2z/Fs/RD9B9L69uPZdFTWfYhUogUwj8qy7WlC5ozCft1wmTQnB5L
Ho0FoZu4nMtI9NWVvurCKAlhg6rahAnvt+bfVYhv62Qk80MtrBuNtBBF1TSS6mJh/GxN7sv5v7J0
YKjZELUgEQ/iEAGCbheCvATWNZTKOaJeeKyzmekLWf5WldnlNsNyNFwR6v5bpBxKP/sFlMety3XC
i70L33/QYsNqvPEgjV7oqsDSLEEZBoa+ZcdZKJmeszyk6OXjDc1HPl7FsYcPBwM+CUo6Z/NU/4Do
c1nsWbYzOLnPUjlrwEj2YGGoI17KxYXn85akh9Vd4MCcLJ/umbvoNPzVfcvwZEHhAfkiiuZWIsGW
hW5VuudAFdOfn6B4GPkEbyklxLF8TvzHvMubrv8l4EycU9Nvy/zcfN7P8JK6lG4VnPZb0hUIRhTu
OVkm0f386mBTTnu4FPmA85oBUxbCc+zktL/vJ6vXu4WLHdUNA6nCbDF0bjm5zMclm/Dl1f7fbGol
cRvOq5rRRVFV0nnBL9zTzq/o877ikkqC239oBfpCIg2gH3SO/Bfg/W7N2vWu2ZbaH1RlzL0SK6D1
Qk52s87MjGMTZ+cxYjpxNUC75G3oeBM4vGHg9khX9Lz7Vg8j3pnTAkqwMJdbRn/ybSL1VDLLmVSe
qXbnAIzVY1magtFftKwyP0jyFKZ5SCIBHtRisPBxd4DNPCmKMVdlpXiEIKkIi1SRr+d0Nh/MJ8Uo
SdL/o2N1Pv9fEo38pRXTG93AQxbg5IGbvH4+qk44a9nDQk+qKqSlrFVRtHkiCh1JwZTdFs4k+liD
Lzk+5VesirRIa5lcveJq1ePB5ryYInlDRSyFiyBQUuW6y18xyJNgjv7QrfYjSpACRdpqPQcydS54
CIf4Oj1u3DpYbEjdVkE6bEI8UzMOWl7GRFjYI74jn+CDcz7T6ugo7nvtplHe2fEnBaPal49Jrg0F
xhJlf/CCx5NGFhn4rR5c1A4KGmdI3uHJWNZHO07elVzmxHaerdRznwjyj7YlFSoGj9UKUtKrzddg
8MZEyKAaYHgXqlXn/LxftBn7BMjdyMLEwNaAZrcWNl4VElk5mJHddGS/nc8MAJfvz5rZYQ5dFBds
Xn4n1yKnojSfVVx/kwHXZrPYKOZQ5p7mrAEFl3DCCbhHf3HMNU5Fsulk7AbMygkWvkCRmpLrwb3B
iRqpU8CNHR+KipdYfsejwAU6K5lCHXvHT0oAQ4xvz6bPKKM8Wb4RcF8GhBG6kl3qGPPAOQ/DAl24
+Ke8GrRuSI0nKe7QGD8OfVWvXQlcv7uhtThImRRlEpOoJ+RMkbSFScCjtBqlTVzxYr5rc+ks6kGn
a8X+Bd1NeUcKamCeoxs7yXPAbEOwmdiSwcZ0RESuBZH5YiXBaIxw2Ffad2gf7S8i2VYRCnS7HmMP
WuTzUA0Hg9neBw2Opr7KEN8VlLZNgdIcUh0mNidwDGi1qn2jmwWErCfsPFO6Fb99P+jo09xxL+mq
EGIXqE75XpKf0MUNlAviyV7yo9tDq9Szpj+oLOcxq8WnJMOMWwk90Y46TXWxg+jXpixXewT+ylPK
m+GoelDS5rdhoPyHi5yBt4DtelMKnpPXjttMr+bnTSPRy2Z2/TCrkq7WSYaO6XmBWSJs8hnJKC98
sySN+RodMzG3xry2LNcxHiekQfid+SoTiJrrA+95zc9qLfk0xAzYyxKvqCQBoLR4EAMdWbnt5ZSl
4nu1OKM7M33KUIZYOF2W/2NEqF8YCLSnwxnkFJ0foWy6hpeROgs8Lp3HentJ7Pa20Yq2GME9iynU
Uuo4E1OfFl0iIWE8oY/+zqauEOhAU3jbx7+YDl3VSl3rJ67ZrwL8Gtn2d3bRoCA9J13zO1m2N6tn
xSY01Gnko1+/xLNs955/cdnFGB10+b+GIX/JnAYtlF1Vo53/o6AXMlLcIIuVFImsnkx9KK9lHJpA
okpYN7sFU0KNYays+nbx5VeHJCtq5UkGO1/dZJbfWj9pRR77/J7k31DG9ixmU9Pbt2p5b4j9qzMc
/RPHxQPpW3UtO3Xzw16vVsaPl9JxatGRZFl9jjk0CCYq7pvpcqB8qiLS9Ctd+FA3T/CFeD0WqJ4f
Hv+ASNKKm7cMRe500+6Mvgm+sDRIAstSGSn9iomfjw1qIrpeKIuoPqd1X/USPnL9RkXb3r8I41fY
WKTxkbKq0mumcP1zFU5DvjFTZ+79XpMvQGZtMnJaA0rkRcn3D4khkfhIJYNgKkv0zTd0lbfAw9dt
kdgShIEhUCbT70jbcvPDybu0hDeBnFDI6DJLMOLB+nSFs4aggPCK1FK9Fl+Lwdrx3qYqSb55jW+O
OgRNwGxQ8t5NVBvQrmBYmyq87ya2+GbcA7PFcdWD0rhrJqBApoAIAUIAisa9te/SJ1rhrLKXGCDE
WJwgpvm3rYih67/OCc3+GznoLc7ynxsJpWH0EaleIhaf4ARHB+1d72PIAJL/cH9aOHY7+8EI+AsC
ciJjiABbL2ZxUq568jZ+rrBLO/OGL/9rChSmZd6p8mTgKW/yc1A5h14aVNeeiwCRRQj20suMAIAL
zpfj+MK7wjwtE/cfSKqtqiTuBrouoyNSWkS7lCkZwRRW/AxJKTfTHDuy08qnlt7Yk2UeMOw7EL2y
fDhcMkEm8Il1bE4AdOoDvAIMcxSLmgJBuNKSjk7mvT2L3J1cdBADNqzovX4KgfUh+mDt19DWmarK
HGRf6OMO6QxsjwlPFvKQOpaJ6eCYEW3bgPDqVdN16xssfECDbq278GQ2FkVRcWoGO1E3EnMJ9r4K
rCZM6iyvg94Bnqoj32bddXy3FK2DAeUDUOsIalYRqY+ZoWbJGx8fUMtIKHGslVhBWnNBMm4avm/S
W9WqexuWp32x40jCTw24nmV2PMhta3uQyah3mZsPbmlvP3cmtBNqdZt6IVk+dw3JVJt1ZnyeTZQT
2SZ6RzdnXOOlu9cwi4d1hynzZS6DDFlmUzU+WUrMhQf2bKbbKIZSevf+I8pCwkuy2+kAflfPLAbs
zsMsGGsZb4LsIHWHI3XCV/BvW9HfFVu+KTk/YH0Iq1ZCc3/jfah7NUY7e4lo8aR8dlB2Q4yzqqKQ
IviyJVkJxe5wnDoZH0Lf0MBZVAa0Ba4uxYMxORt1/aXqWsGHHMOkmeqBOksjMzauoRA39EwVSmLj
vjeqahR2YLm6s2Obl4of5Qnmj3wyZHjowKkU7SPoPjK5I38rTp8nWJ37bb7O15y9biU7vuCtB465
jIYTkAL+dCSne7mU68RoVMt7Ae8vMROJzPfa68RZRn7XBg7jJDMh+JoewGLrAwat+D4+T9TubTYG
HzZboFG9kItxZGAAGH+VlEOXG2LFbJyuBmSbvwj6v/W8zG0vCvQioug79sAthiARlPSjdoBsoKWv
jSk/uR2QLk9QNHWQXoeONRNqaLqaJqiPWJHpxoVFGr2VZJ8ztJLR0L4DlkUqYJsQjH9Mta/txUV7
iKSmU4IxZAtLS4oH+bgja51sztAWApMJ8hNTo6+ytTwZyQQ7qEYGX+XP7b6sllnDZt8UlMZ9e7gj
Iur1zygWFKlio9vU4FXn00mhIBi2wa4bhRwB+GjcZyOxMlsB9OvTpqTlyXkadtf5mxIm8J8Zyn8I
MQ4S8e4Gy7UiWpSGFTpJgA3JO3ke2Owyx/sbtRXUrPzIp/OECm5fxDIrxbcjlZ9AjXSi6ExlRmaC
jt19wNWZyQYVrr1szPhdQ5viI7KIp2wT4ChOBvmyqpeLETNFS2wDyn0rTOpu20mmy5ZfkVlsJPVR
hDgaFwQsXNJfF0pVoY7qGLbYnk/sVVo8REEpCuUJB3ccQCxEYQbdflKqNzzrku/ua4dVP3QTvCkR
nnYCCBmihEtW3dMp3xQEhaJxtKbME2lxamX3/T2EMShh4C5hRveLNphAfo+nwg6u/UBeh2as70tm
Z83lkuBXaakR1WTuGWvlBpZ5YyrmZSv41K145vsRc/0BHjZLozwt31lWn9bfPGxAW+FzDDiljOnC
kMBxuXRd+cfiaUQxHsRSiPomCOmKKgohTV+coXTF9xxnMnz9DYNSxwSrcXbzLy5jKktbsPGLGmjE
9SDDB8rCrLXxX5xba0FeJNouG/x5UcO+JAL3nqdyqVS9XjE7NouSjn4gpDst6NfJUwKao3O7nSrH
mvwsjB/uUiYzlmQsyrs78Rz70fWOyO/uZEGkdlY5kzSA9mZjX91/M/I6LjyYL7wxbp5GuV23hrOn
i33h7py15fafUNsa+5f3jZqgqXvZSxlzlsFLMwI49PBbFUPAHzEIpzKK1bGtbyKEAcyisZz/Oyme
q3kpZ0R6DKg3z0YXgILpQA+AWJ6Aw4SujtztPvbtohuv7++qzbGpFLJXanAsOEsZxRF62JoxENVN
uUlFnDUes24ggc8ZGcUYqAOqk/HE9zcadu4lLbT0zy2UT1uxti2yXD6XhwXQDH0cL/VdtiW/YFME
4rmGmiBYeRpXKYeu8BrJl8YLqUYzlZP+//Gs16/KdfKebtMGRWSnFgWNfS/2xN1k+AYd3FCcnMAa
ebrugc7RWrqc0uucyNKlmaqAg/8jW2yneWxWONZZpdZ9L6Da2KQs7d0Zlh27gI5KH5los1xQwb+y
nAKM4cguBqMw0qkEgkZB8fdlql6QlQLkKfwRrN25TY1zxpeBenYw5w8hg1sfkynlkJ5t/rbK/x4i
x4uOglJtoYfOfdxo+/hnWA9qy+iQrdELP/1ZT5+w6kZ9l3H9gM4TWKu2JJ/WrOKsy4s+X22mWA/V
lqPWDd0xUvynhRgyxXPc0jgqeHpZtVQfuRGk3B+hAmwbqAgNRXXGmmjYNsypCIoiGQFqaTsBeyB+
H7Ax3e57mxSJH7l9kwuT2xMaYJualuoJ5xCkqqFEbn2p7RMlnYrh+uYPVwAS0Cp5wOkyYOGoLGjd
LTv9RE3CPJwDSH1CVv9YOf92wS5ZDXJnld/M+MLssOBnhuVupURzA/GlW9KDzJ1dj3ium/qQE26R
pUPd68gakwmw65ieMXJJzANTscsqb4wKlNn6mE5HXBSaYdEkbikowYPOdVip5946VBkqv3czshE5
wg0skQ8D4Xcf+VD3HA8w2M1V3gb4N+G8kiE7OY6EG4SrBRjo5sncZt+P/YVtftj96c1rNiM+tp1v
ULRoF+gxZ3N4vutQkasEUqmGvTjGDRwyia2wkh83OYZs8bju4BsdH3NCRMlsXWQ9rZgu9Cdb/1Oe
9+Oyyo05Z5Nu7qTifWXTDD2jGeey6K/MSQS/pihrxqgZmOy7mtVugxr/Gzq9GQfTowszuTzqUMEr
9lZGtzKIYiTMpQyhD6JkdxAkwbb1xL1113C5zfhrOSt/2lU+0okwphHKkffTiNj/Tklfvv+3Ofvn
7xA3hO8MNGWjPNHwonXIcV31zJLDDdJliukppdyaAJLuplTro9n9+RKh9k9J+bfyCTkJXG/+H5m/
YfXnIQamH+CQpoRQVnnD6CxfS7UkNWicYHK2BmIdO1/beubpIt+dV0hqdon48DTHTt38gecNOLz1
yearR4cfW6F5ql+j8fLzVJGYyJzYiUjNQ2D2Nt1NHfd8GhPf9JL8sK0AGXxc1HHuLemhRMF8ASII
n5TEaTAZXtNanaI4HsIS7HL67EgSNmgwMFGVMuF9FK211/bNxTEAhEw3KgSJ4WhRCmLpUf7IWbH2
Wdo+NiO1/fNIpATdrfYwfU9VoY/umknauIObr2jkHmgJmV4GSaEV76VP1i7jg79z2OmeNpQyybEa
fiHinqXYxSjIGEgxFsy/qyYIVoNvgLHLw8nJ88jZrzlSZeBjxYRHKshdOh8mw7ud5/NkNQQTg9dv
7m8b+ffgQSXrBwjOa3mlZdix+3LwsF+zC3I4jHVUwFiY9RDnaydDZRKnyY9FPJCMeCMp9OkI6sd3
s1eUiTSc16RGv1K7KwEBR31w9bfrhBNm1kRt4368CLA/MGlLRSA6Gt56lNGV5zEeys1JdAXstQ3a
Ev/78IykAXd1kkHTtelToTwPHQh2cyGz4K49UwbQHhFJycmAsFPNSzUt6Xjo5PDaayIAVbOOlf2Z
PqV4JKHtkBh08Kz1d+RrlymtZxsH8gjONOJQ1KOwXJgbck1IoxCUHBfoliVEmlhYpdYxv1Jxew5P
JF+1xRpnF/Y3OX1TaP52zst6yi6k4aSS1cQrr7ZGrx4MUfh3Vz5lGZ8Ud/7IU/bTlRhn+6IQCmGF
iStZgE9hiFWA07bVnfJNLN0f1CAU6hxq16r+TUbWl+z9rhqUJ9ZgMk9AwWYN6iVOxQy5l/7TlZHv
1fxMJ84xbFLyQIoGS8rwNawak9EeGsJ8aSrunfle4lgp0jPxcYqDjst/1gaJt9t4t0G3000eaqEP
cr3om1nz4wF5f+voGCp33WrAbTBBRCHETuAiVy6+dNOFm6+hJbwl9GWlBUwt6k6263At6Hovh1Mo
lTf6MmXJZ2QBKp9/W+S4j8YYhOX1adMPpjU/AM2zS+SlwGEe9VvS/yuc1wN2afHWpa3lOiJyScVz
mA9+mrSbT26XJb0B8g7rlbXRK7B+b1f32NHaTonFib58BPC6b6KxXh7V8I93BCEXjAfxWIELbkO2
Jw7D9Hg1Infxo1w8axX4OjkLRkQVwUOAPACo1gTyJ117oDxtWoNSL/8llJ0MZYJzgQtMuq6uZItk
Hm6LCUTNTBKvScKWt+ye0UCJmfpSe/Ng+fHGPtj8YfehO5rx3ROa32n1nFyxO/ysNq04Dkm4XJop
3Blt+kyASuxcThr7RmYl4S2P8Wu5008TXkG+oipVSwQGYBtbFdDCoN5KUgtWZZiEWMrLYXhfCXeF
h7Jllo5pdUflLwfn4LCFNoiWV/Oyiy3OUr9kVhpKU94lqWRJ5PRfuwGSm5FJXOLg7614beXfbKLN
MF4x/vZ77sQjUvve7obxn848v4wZWxh7AMuGNI9ukQpAZhi6rsTnhFusODoxtfBAwZSZTLFp81VZ
mEcQAA+sD/dJcySCryCmOfToBaTPfrzcn8lburyNi8uwkpYDjmYaxigCkYCvXKGxURK54fznGvyT
q0M2feHtrml6YRecyhonofG8KZDUgDm6OE50fZohol0kxLJKyjDa9tYcgwpHiX5egJurRGUTFrRH
oPhe7EagNl4JXSY+aqZulUc79PjwE7afhMHpa7EJJZAaB3h8PoY5bNr2qWJwxVhXKaEZ5iSC41G1
2A1oGYNoruMBytinzRRugHA17WtiNinUc1yZacZiecEUQn/eQGlR9ndfwKALlhyTZ/As+3UZJG+7
cP3LzkJRXLBkghhLn644YetXvym6mSg6ceNQHUKTDKGHHIu0TAXRCphlED3IRe5KShI/KiSrzv81
emK26VbxNITZGzz4KW6kBUXIrcMmObQ3qEO2XKyOBTpj3RXAVXa8IZBq1aZ6IzrGLPfwijMy1UUX
ErqR2SOmXvMQpHuDr00/J4JvgjdrzfU3Q7+qVE5Uv9l4+RV5yL7bCz5m3uMzElsScwfuC2F/Dc2t
ycau8ruzrC+zHTpP4MX4FeT0ySBc6rJ8lID5dGfKY5OQJmdR33q2hRuYpdVPcMwh84djFWCJDWmM
XuxFzhGewEiL9iSi4JYKLJu/xQmIJmIkqI1CGivX3wrH5GzyaolsCnCAdni8QE/k8yBLA25B1uuL
kGWBKUKg7Svxlu5HlbJjZ+94GavaHoWNckkn9O1ttuTxY3SOfCPotWrXNwCnTYFcdHbmzWxLRY8B
5cH0jaJvfWU96tPYvBtauk+h5A1ZTkOiPGT8J4Q6J8/DiFz0blNAAH70/MmRd7MZm2pS6xuT6VCE
lAvQMlZFOU53cZeMV+T3NOiv/HTqQt3I9SCekBx0RDoufnUuoBrn8IEeeLNvxbUpvcozNmq5S5e0
0XGUYyFL2dxsaXl26vSyHL3VCI9ROCrJ4rK/3Ov2utUX5K8cuFb4vH93Ri+LP/q+648UnB+2fIES
sBs+4xErc960iG6QjyyFpm9BNKRVviCQnLymPDTPDuyr3No/+XpzmuPs/DuAFJGTqz1wR/a154Mn
L6zEH/E+sMCPVAgJKcNDF27wWbN83lmST+y3cBtsOqPWRc69rd+yhrJucVKGndyRWy3PVcgoXq3d
Z1luuwv1mjHZStg3MUKCvn8BLT8uOkVbldGmkPN04gB85Wi0dUS+8WWiovlk2MDthJYqIbqlb0/r
sZYxpJZzUyV3Vgm4jfkcYKbXpKKlPaLHVQa8tCNv8z9ZbOoPTza/TzjzbeWLc8l8o4xK+14tAret
2Y1kAinh5a4htZBBM1XvJmjXtHp+G4eoxLN6AO8mwWI0T3LkIal2BPxZF0hsw5qBnQVdqyaY4AuA
IHgOoskhVVWmsyFAjGFim/Z/o3IYHxCQCTafQWX0h2g7IIkjKefwpunhy9/ZLhjxvKb5JlpVyk+p
sD9QHOOLFAlf2ML421DJxtANAfIkXFD6V810xTgqPgopRXVKK4wzftpbsSjePYdZ34ioIeOml3aj
bHVW78n/kcGRVDzpJwluioZXE+BQ3Fup0qHnn/7LNx1K2o8cnnEwQlC0oeWLXM1XNNkK2RyDCrrk
DDZxyPiunN4LwyZX5YqDmdJ4mDh79OrItJGnPVPqqAzUHd8/TtylpGN8tdbntNWiwWAV0+odoH0R
LezV/2hVYq22GxzYC9nl62iNz+H3HM9cfbvbNX1zJg6tns/G6JsTY5crfLtJA05nVjzBjXD3aAJ5
VDFv/+piHF9X5cj85rapL9D1WjeGzXE0mgnD1so9WBdKufMntMrUoBMuU1aDV/3x7r2ty7uYmT10
tcn2twyfpOwK6q2Ls70/sskJOuhbutjkXSWSToDYgvV5eyWrK76nKfPozlnLB0bsvbDA1carkVxz
RPJR8g64cg1PrbqQxFlD6ZOl9goL8UKtI7Ed3uVBi0uXxC8N+hqGR37kSmrH/eanpQXUObcg5QCV
codEBSPqGdxVfsyTBAJAcawJirDYl+HfC03UeA44NxZBnQrjhUUNQAMZZFpqjtSAI78qcLZ5XAIA
75gZMcg/7SJ0GAZKUEj4BGhHtUUYagErpdieI1H7MnwRTPsN5TqEC25zSLGDeyTF4K+UZ8KVkrbn
1CpTro5y0qmQ46cIJaN2CqjRR5esiAB7v4v+ieYL1ILLQnuks/dWjOhmK+JJR9GgCKwmFaOdOtbu
W79636odXWAmOSnioOSZU0+7W0PM3Q4MgJKwGmBDagmX4J8L7JW621OkE0SiIljC0NUqKi5q/I0v
QE47OsLt8xi8HPojutOXOlgqiTSEueMDPy8GxJZL44912SRNxFVorJ8lHkp+zulboeAiQg1JelZH
Jjp0ja+gpAcb9RJzCiX8yL28QMdKdRk79oxOL9cPxFEJTKRlkX9fK5+Rp6RFhGOnFygzNmQMPQqS
xzixXU2Dlyh6MwBtQiP/mY4FyfTlLtw5xvZbCRkrc0wql0Inp0WJ2anVQt7GAONrRduIV9xziPKT
VQzTPSNOjt4eUuXvFsJ9drxLJbOY1nKhLj9ljYECDmFbZhclVNAFQdZVUwj7VSWNoYN4SR9RD5mo
sjDVzYELgijdg4Scpzi5XCNZwkjpNJpnOWVyptklYAZl0R+95unZxXqpC20TZ2+GPZoxOZzKPyp9
hQNcpfMBztW5itd/LW2XD13uukL/HPtKzQR9q5fnlOuSsOFwm9z0uVEi2QSD0llJqjVwY5c0f1JE
ZLt9F3I07ycSNnxvLSW5peQTrq4iBvXYuHlj7013Y0M9RiYKekn8p5huuUjZrD5NLaN1rnpahT0R
3abHiGFsI7qFesK9ElSsLJOx+H2nxDfhNS4HjTIpnY4kmMNfywqpSjNH2YO/cTrzoO2QoyGagdZl
7OrOmEucuwGH26XQ+gLlmxV6xWPHGzUlltJL1jwwk1mwvzhyldgkB1oggGXz1QDmo1oHDaY2O9Fc
6gjxQCgs/w8tlyeIRR0uCHwZOcFUy6eCqizCk5fxi9uQZRb7p498hysbe9vQoBdl0ZcSbo7vExBO
auKRNbQpL+n7fcTY1ZtcwVdUgul/A1Ui9ms9kKQwMTCPaqD3R4tcYR4ATVBHJlvR3zaYC3aPURAl
R9+M4WfjUEIokjvVyPzoJPFJfQPiP1kNTjQeC152gX5UZwbUJHymEg4NZduE9wPg25R5UCI7+luc
YGYxb7VY3jZfUjxmOAaOj7TJH3n7vm8XiDRczCoVprn831QilU94H9B7z5cK0OKHLhBV56WA9lX2
PanoVYqB+P/slDL01531MreahF8SUNQluKEb2vgyzsHC14lZ66dJpKgR8ueQg/stujdcPfhNDyfd
nXE/HHJRHs2b07HcdIzdUjP8zC3zk5glGImE2FzNqTdpDeGVMrJaiB5X0zNsLsXwbA4/wTaKY6tC
f6InBEq4HxUOZ7fcs6iynEZ71XJKideXvcklmjsyFZEX0hvqRehfrta4965HnmQ3ixmv0ETzNkSs
dIH4+yvVTgemCWrouzlyWElgdS8V3NjTpHmbgeMdZGG3Bd7k0JmcoOhowUNQ7P0c/qWQISM9JnsX
/TQPR2RT+Adl+9CIuLnqAEUeojDqZLUBierdhN4E5NGlmjGbG+xCqQvi96I29NlE1g5Jm/c83iJ2
MC3wKa0K0ythee05JfmBpoxRGBrIN0t2QTLRM2q8mKNsNQauv5HnJwSjen2hemkrPqYIJcHsggvK
VHFME0WcZbmNN0GbeZOUq8rUgYEReJWJV6zxFcbUWvxDEVa5n1VaZANLH5Hef0w6sqPzGHQtunKt
ulJSkkJZZ+5BkaLcF9dkJH2TRMPO1pA+J5C90Ht9NWDrk/IxkWmrx1CqQxxuGJxy+eKxiZSxydGG
ltehw/MopJSYgAq/2BhUi4KKSvXUb2NTpWfw0JKXH/zQ+L7INzWXz5dgt9BMc1M/2vsL9FB9A2xl
+M4au+U4yFflMB+K3JtXLuS4SEyqnB3Af8Do9DJCbeXkyUY3AWwCODc3wAmzR+tQ2xE9p88UmDNO
fHK9SMKjU0IWWamb+d7fw2HWnDMWnTJEjKXGZhjNbj5+Zw6FwlZdxAeqkDC0irly5BP6muMkCdbA
q+UGjM8q44jAzno5QVSK39HAuYHLhD+9g6UmfCkpLM8mF9U70CjjgLfWhcEmaJVpDHIBgHvHC00Z
8UzWw0tqP/+QPONi+0ex5hytUKy/XG79fjEC5H2/KWcaPij4f+ztkAJlzhbr7X0MaU8QMIIpAjw6
ZEf6lWr7ZLGkkUy1AoWh7t1suhvOK68VcKwK07XsOJZDRqS5O6fIy1S0tkPUI0aLElFQlXynHY5e
d5mmXpH85KJzJ9fMV2FTp081/wT5zbtUO8LM6w/75XziEb9aW9ryLfWwYXaSAlTcaPj7GCSh8D3t
IUdSnSswROr9czT/Q9EaKTPeYglETevud1p4N5jsgXxSksSGT1YwISr2BJzze96m9BBYa6j+g5ki
g2HmMsrXRb+HQZKQjhHJ9Ym0aNhHAsyJfzLE2Yd2s12Sey6oc5BvKDev8S9vn8rAEXx4KgtSlaVN
g7TZhyb5SunToKtZoXv6dgVk/GB0hp2Trt667o/Lu48/w3K/U06WzIUb70mMEzn2xsQm7q1jkRWl
8UZmQvDhf+zkJ25MFKIkRPLB2iRQBuotQlAGzsJD0zhl80v8J4fYzpRRV3JRaoKGpyAD9ojD+L97
kJC18OxgFZF/JE4lwNHI7TjcyCSMSprLyQIswzyDzNl0ujsHTQHY+6RCA25THlt6svDx2vIqchID
dsYCTDD9+SaaGkapsn1JXHspRaoZ4p18/SGBdX+NbZ8wkH1jmF9V+uJvnM6/ME/lB97OuLNY9zbE
D+HOet0o4K55hsAhGgJKP0DO9+0LhuRxMzYKZfKC5OMbC3YiApFJDaDeGOwf7Wg1kWh2bN9lEdS1
rOgxyADXWE/B8hLkokMcthcXYOSeVjIYRFmDbQEwF4mB4/7tXHT4nmR+xgz3aO6wV4ZztJLENhwU
buBk36N9LVGhykwoCis6PcOR7iDCXAW4YBKFcdjqh7G1bjfVVQMfEA0tgfA6yyQCtVfBJN2VJtn+
UWs18vPRVTt0pyUPz5gODeSu1spuf/02utZhQHCT6PfAyTRQ6yhDtz1Yd55VQtcLKUOAQgs3cves
9XxLF7LXGtUW4vZCz12CeF1YPL7+ZQe3HPJQ04B8RUY/JL5XEZQ46xqgpc744nbsGQ+TI+6fwaWv
tbsYoEnOLC6DjYDzBzjn2Nbv0Hf81N/SPwtVehuTZSqpn366Shab1Zp5IAuxpYNKNNQQxj5jqC6w
/td/Dg5uhXe73o29H2xzSpI6rlmdGqBEeqEC3QOFLwzJaGz4rpGOrTPzrVjr+ZqIYHrdjDv6y/Ns
ZYJr3Xg8A7xJJNF5MZi9+ultYK2EmtJz/+NnTs2Gus00HkhAtrUOVuf3VxX4M34rFwZuc73MbDf5
5rtaXI+HcbM9JBkF/a72zF9uZmYrHDYFC1mYRQ8sgVHhhhJ955nbOUcOgE6mbUkwBXmizk+4CD6Y
tBFv9mpfmVVuht/WGDCAzWvp/2euKEn3IuzBctPFzG02B/f2NTALJEt2LE3boo9duuxo65oIP822
wgRphw2e1PuhsEWt3+HJ8oD2cfaHlEru2TmV/H2DLh9kQaMJrlvrgr1HVYj4EfhY1ceJheAhfjYi
PZNqJXwd7bRfltVx1ZfkvC2kccJISHe2+Hjbw1xPZewVaRLngwgqZ5b427O+bQHReVC4+xp0vr79
BZKTW77QZmJW8dg08vVOpV6A93KGF1IgJmiWIS3v25XAPDUfGfCn5h9dUG5CfV3SSXNVSEBGRyH/
U1/TmvExRAAKRr9l32mhXAsZkHs9kicHONLpfS3EIj3l89CZ0q0oXjhzx58v0K2QPMCVErv63+to
eWNg9kyMK/LPABaG31uFsibEgdj++a/IjY53c2xPBA7zNPdAba1PIP2S95aG919cXVDxere8jlwM
3CoUS6mtfkVjC+VdY+t/L7Kb/MvJbhJ4HC//1D3gYRlqL4kcpzz2cCFDXpslti2IgSuZVN3XC/QR
YV3s6BM+8BVKWz1g4q4+3p9yMxCKFrp+hbFHjXnU8GLE+RpXIKEw8QQyuEiMnwJtYPyTO2m7YK5d
QZrw5+QoBbKlgvZQRycr67/XIh3Vqb9d7HXBEWDlgNJpgL5vPR1v0aF1ulTOJrEb4VNOpqUOa6cq
u8xr20cn+KXzwsLcHleJOQonUaWRS76awzYSrwlPR0FcQIIzaVFXgDkOn1rG8DCvwWpZqb8E/G1A
JONKMogBSVl+A88kbk2Wh4kpeieN2EhMmhn2TU97vv8pLUakB+yETS8WBQvA1qzEKzUkK9Uy3snI
smXc7ipjPN6U87QbitHoDOaHVZB/vbuVN0JG/h6mXgPH9tbqoXYLwsqpKfwS9CsoEWcRaw6Ev6Mr
QhR5oYwCREZA1dkoSVqyKTPw/hgXmq+PYSGmxTxnl2SUju5xYprz4u293IqW5MUB7GSJhjrLkWMt
8D52kXyICzKfQXNF7JJ+UmC/C7Es4kRmineRRhGYeDC5qRS8VoMDcROr01ICeBbqtX0Bf29OsP0d
s8fT/RiG+9TdzOLbf8JRwLpfM+7HsC51I5X9VmgD4sPhTwFOPevOr1CQY56kMtxvqyyqZm5mPDa4
8Cd/KGJhZmbypCePVtOPsjn58CF/7Ia20UQ2lnEIL8uKtlbYmB3DHVscS6c3TIUSdIURErBfB067
Qr13hs5VsIi4PUS4ujAm0vSj+PhgWwjxc2h6Ewayn7hbcQCWKaK0HTcIFDSZdSditoS5i3nA5JLi
DeqkMrMz2nN9AuEk1ytSBtpGnZpt0CH2k4ffTfA7hs+AjD10OsTl2qLbKSDBpios8QUoJUPPfSXe
sWGufixYVZ3zF2JTwlu5YLA3C2q3tU8ywUIQ6KJZr4eBJ/MW9SgRWX440DJ5SyTx9/HX4Xh+jTTz
daerNp+sJGbzt0mXqdG+nMd0smkggCg7tROoxAe9w0McCbvyPbcepugcu/wjDTicklQZ5Q4gY0Al
d1x47Z/+NZfoRly79SWVnERopNdqMOvyL41ivm6KQgJKU2C2d/PPW7c0OcIhl89WRwA7h3tt8tgU
mlRsbx6snT8t73Rg6KGdLGxNV3WUo3jHv+FILtjAVXLE4Psi/bqXmS3DaqBU0XpzDZDRwhBniwNN
m/1R5gL+Aqz1RMbpB21uNoO1D9BuXM1u08KovYpp3NWkMmJiTgJwtuD2jiZ0Uj7fenScsGpWU4gN
LXQrah3pNq/pd4anP9gJWp+rbapAprh4r/YLPJKVGl1GafIVQdvJmM9i+5OxBmmQL0h4fHrxL7Gl
yA5PhV6a9X0UBTuo8tXDQn9zHJZPn5BynX7pa9atuGAwqH6lm7aOmtqkXWn7xZCFtcZeyJOZ6MRK
zJJ36+zK3nJy5HEpp51lH152uNXZyJtytON1UgXcts2qDDMHemiPcQk3AOvteVousyFZ6KOH+KQv
0ijfPWM+0zbUNza2Z+2kjHGWGRV9POG9b7Z3AYXssjVCr3YbgFovqp3VIjwxzD19kvDbWHPGqyDZ
UOHsfFJGkkT6UENA0Ou4Q5qeEK57FwvRx7HhRqFC/5D1Zyc/HlnzrGxPMEMTNx2ZAbfCm3LTab+y
SR/Q6WAGXpxng86m/JO0MqKJqJrPW+qPmnzIsBohDPW9sRNYJzkSZEeUTUyIfevpsyrdgazI61+a
Alo0Btv7dY0zJ/FnFlHSBjppW20NkLXOu8b0T/heMVD1TtLhv1rmOmfmIr6G4MtQ9/5qGzcutvpa
fCr5h7ay1vNGp6yw+NSbB83uTMdTWTTEL+ZJxIF5R+DrlENQYhZgtRx67Fj7zIysH+ySPtXgR4E3
xX11NiBtL8hhWfywXYJ1IGY3niURGNIOwtzXo7fgS3SUqUhYLiXFcysxntA4V7szW5pqMISHIqSG
g8y7bXCgkbonkakjLdJOKP5L+8UCUYDpPeJc2iO8iFhuMlI3pNQrT9kuusM3Q+iZnllyhaqDWNxU
d4wgoULfdL6WR9XHxzArKuZ0pogHHJa1FENMMhDdHHJCNqgBBrBNFnDNVvwB/w5saxUvtNDhCXar
hgk0Zha9UWMz2dZt5hThTtmSki23J0nG3kFIsBPR4d0d+0Mdw1tsB34zS0A2AqOBORE3SZXNGs6o
Z9yfVKZS6NUrjOFVgCFzsxLNVFaCoccXlns2T6K+uGFdQgnxDOLCiWXtKn+8I8W++qhHvnbyFWb3
0gFLq4ag+Tkr5XF+Kqz1UzNGbJUeQPUfe8UXRgTqQ6xirONyg4mKIUXgQwbHtR1u1eizsXBKSeHL
iP9tPV627FQQMo6B74r1p2MGsBAMNnw8w+p/ccB2hU+3mMP6s7YN5K/S6iHzJoYD42TkBCkGyXG2
KNC6gINqfcWza+thu5HmzCtyeXilS7jcQ/6+ikuLqsev7jAq1YU1QFpN86Cm+oZ0C1vztgyldie3
CdoZ0eg5tutktb7z5ajgHtYs3LnFdtyFl1xG5JzbnjmltWkqoqCDdga34wgHiPhlzqCcY9j+hWzL
jUQN2zZnSEvIt0NizBBroaH/L1uTOV20x+zmOoBwy7P+VIhSu4bB78aXpO2bkBGVm/7iY55OfwEz
rXNGmg6yVPC6Dm0uaUeMwQR426JgvqBz/gHb9a5CuiYyls0p/OhFq2ffVk7TElz7EELq8SfeT3iA
v2+W6POp3pyqa8X2VG4aMLSBYoASE3J8Oih4f6v0JKdLClJGKS70Y7xCHyIlMrOETvLE5dvOTpvt
EWuC0WUsuedHeXZWxMjUfDltGdmC4BvCtdSGHhVBY9e34qHM9etQNTYdIjNcZND4+GcO2iApC+Eq
t4UnEcefrrf7wDPqmsshcq+mqsdHs8f9SzUIiwGTNRwR4yt0E+vobYik6uq6POXyfhUaJQckLqe1
6Gjq1uubFIHc8AYi4kUVItpln50/oiJWZX1rkZo3j9RXPLRWhT/mWDYYZJGUBjCktrEUhnWzpSUY
v0sXBY+63uzNjJuemM/b8parN1kv1KYBJwyU6x91oMC5ZHCDkkpe/pfr1WorcaWYvDXOOD91rzwC
RwmULw/oE8tN26T574i8R34wWk0GDguQHze9/JJerCno0pMrJvXMOACyBhWKnchekDfQG5DxeYeM
yHeauOxepDUV7JHwkQY4OyAgb3fxHWxk5Oae5DR8NbfvlVGTsca+IXalSM+Q5aelz0xida71hyp/
Z4AwXVErkELCDbRqshmwKgSgwBfHf+oqn0erwbTnB4yBD8ziVbi/Rn0TUVDX5+NrhoATtYDMzNqK
QEBuzdyYMxje2j28KnfnNQ5y7bBis1m/9s4DvKoR2KWkLSw9cKe47KZlDkW593BDL+8/zyLkQwws
fFEdjTzT+7sYrMlIwacU/tIVwmH9+l6Ad5BlIg1TmSdoE3hGkeSXrzRG5CdWHABOWLa14Ru03Wld
OyX0ve72Xg7vBFuzmfWs5sd6oNxh1bCImkidYYjfJe1XcUXU3YtRsZGB9SY2XvmZt0EAJtLcVEe8
/ONSuaGkWg53zl3t5ECDNOuWL8mDhzH20Yn8CAIrhpV5CPnO/5ZEhRPnJNGokoysi2xHyql8/RWz
mHYEDosh8+nYrv+hthF0+73WS/U5QDaBTsyWXPbNiobCxQBbIl/hr5tVSqP125TX/yuy//Qg0qO0
hzlDWfAwmtDCf86rmGGqseCkXQ0XpG/WYbQ6nLxpLQI2QwmBeDu42ci6qCR3ffrsU9ru2+E/oIhQ
Ton80hmgVmvelmfxT3q/s/WFF4NmOZc824Sg48IcWtkfABRVvE1av2PgUR4QtXLgEVVTEQL8KTHl
l+MWhLDnUhYUgB3JuJYiBCgsCdLEMJhLTKZ7SJIFEdBhhQJOhn1ShBsjmSuDsqEsuBfBt2C2TFn6
pkNuX+uT5bJzM8k8EpP8jO37N24XeOWn2U8bubZ2/JvXQLH9aJB1K/TOnt1O6b+7lgCPaEFuDv1w
NNUoIrCqvH1mveiLN2q+3FqK8X9pXdYlopUBOJGHp3NBiFclNpHOitx0HCqWN3yDjnkUC/872tE3
cLRtUYyK6IAd+ZSYPE0LjCanhdBwAwg3dWYUW8VYxZbvZM/K+3PHuWLEPVf6Es3+BSKUjeUecg/J
jpW85pSffChwKEW4KDWewtbS53DdXa2/pOSCP8mVPSuwpiPxWp5wk8UpqxSc7Uq+zhbcMEzXCSX2
GrT3D9LyD9pwmxCwg8e/bdEBXyy8ihpnMEczjedwDLCdPEnFFHRGgWdjp7YO2h7yRkDyjobD50xj
q5sbTnbpXmxK30LOLWslUsZzm7b0KBLBit5/761VjBw6UwCmbgxL35hdTR35diJ/LL+Bn2PNArPu
QoXCZ8qNQIOUNpI+QVmEBlHAl7KxKi5Egmffph4YiIaoREpg3XhA08Me7EyzxL1sWyilqQG/Eg+v
fYcEiM07OKCJ5qse2bCXlVCWV53EUA3W83gktn470y2lyDCjR5YmY0UmTRmMUfkhoivw5uoTu4Y4
l8vluNVRS6zMztvXy6eQlZIGtYiBKmvhlqE0RIkRqhkEBqU+W3BwaHVjCUjkmMlYkQl6Btz6ZL5C
m09whRCgfg8nN5pJWDbtiujviRRZyJtPig2c9DilifTdy0/KcJOZq8GoKxdRmTrCFmZDlcwky0I5
WWvU8FwCuoM8ClpsKAeatgNsj3TceJh024uxEy3TPh5jaeUjya4uSi3N78uReUevVvonDwOtkSQW
urEd+riHF1qVoa6gPYuD2yHsTmeedZdQh2/uLVpmEFrG0fxQcnmV8TiTJ7wcXJcqNI9sPchPqiNL
am4VfK+YHdV/uYR7g2hcf+vRNmIknL6xKbN2c51tj1IvXX0eXJMUJz1sFn7+68WBkkTcn3m/IjyM
7MOOIWwYFwjd/Gd6FBBbdBSI7ns7b9HhMryNw4ivpsxLHwdF/ISK+9pSHYz+TvZKb9AtGfV6mjze
UqnduCxzHPyaoFoOeM6qbFGZ7EgAaJFCQsxevWhiXgji+sqw5Z/CQ7RTcdHaoPwtpM23RmH0LFV2
Spbnjgicb8Ydqr1ePaTNSGB0MpOegqrJTrxZ9zG7xXDbYTYOifNlmVZMDKKnmwzIebxYq67wO7mC
2mKxaV7YdoPgKlSTSfQ+rAXU9vh5cvfq4jKkjVGOHhgPZb3LKs/vJ7jS6gHJOaxNhP4IQHRWirkB
sdVoHoEFpRffNm7TD059lOwh8DQ3KxQpY7Qds4SF9HAaKDsXAyUDbCgre0kL9QxS3jhfaUE8dUBl
PIggXvMlLTeG4eapFJVZr5Ai2qHDnaw+sqWRiDN0aX/XZd4tZyawfX7dQIvAY7udaDlT4VZ1joTA
BrCbp0zmt0s9Df00uTbkQcFHQlJFMHkV0wVdr6Ay21I3ccRxezYfH4Gxb913BDY6fW/GzqRRMlUT
IpQsUSWm+XJqse/7DZoo19wWAgkTX/axauMC2W3pKgxJSgzQ6KOnLqO/djtTsRvcRi40xuuFJWCN
a7+lT49whsNBcYsN35Y1yoFp8Aw5vpKABBR9m11LrKmpK/tfMi4bL0/WrSyNogJj26SE5Uia7zqY
QeVGVV2EGjrueyCrBB0WjSrT1ffmkpKmWXKOdGPHeuajMn2DwjPaIt1PYqpcRyoAEvEnO4fp0F1m
HTJnOcUsKmPO7rjYw8TJAK/XnAAWQy0xmP9zCYHzPy33B/qNDTwykxCL4tFAg7wewL6NEbgQ+jJu
webWwW3iSCNY+M+C8xVIeQqyrPPr9lOiQBC0QrrdzOo95swYsFt4hOa97fzKKlQxZK3fs/WYz67w
6WYmEhQA3XzOb2ahQN6/Bz+vMTdyyHsfzemJ/6vEiURYL48buFIoJlC/0TwVTxm+oqE8agoMHndX
dGe2Wsz/jHzqu7ZeYpfMQ6CmwUi+Fk6OZiYBqxABI3MPk6Hq5/tExICM5rC3aBslZv1MIZjRtu16
DBWt9hBsYeQ7ZX/NdKMWe2R9fvhj9OPBmrKb5tpUVy9c+TCJ9cnwLSA4oOKNU9zR8JFg17jLsJcC
YrkV1Q8WbEjCqJH6biNAL1Hmwgpc/4DvFPo1WURFswEE2V1MvVDfyjdUDakn+ZQ1/kFjBxm/g+2f
PngevBFmYObvlFKhbB8rpboUL7YJDYU8i3lqs4mzbnJ1xwyPhc5qxJFqj5C9uy6Js8XkR36gy6pD
C3CsgEw3CEOYqVUgAwDTfewhMk2BW9SAAwogRobH1IUGmCWQSNemihbYA4QByZ1HRwBViblpWOvC
P4H6ZxrMEexfOZvc4KtXPZ4fHsT7L+DD7dXDsvuzZVWXLMQVcHv4PaMqv6PMIRAMbQS92B9xMuXw
SJfU8mY+fq4OsZ2hGGm0gZ8QtiChwmT3AhhH5oqT7zmJOd+Kta47lDdZsZlrBWthNT2P1IIym8tw
ZMeZqujqy8q2fbs93QaaQCdKBhLI3xj5+OfxyEEqpZtX5KaRmKIYav7QxZaEygP+DNC9A1BYGc0G
cCbox60lBL1Wyk/oWwCOtiHsh04v1lFVFL3flK/eKJOZmrm/njTiVBRZ12P/ekhQAB4al7Vl1Unu
clz2vX9UWboTiwEGz87ghq/QUU9mBQxfqar9HsAMaq02L3Aed80iSbSsPG+inPJH0d76s6yKiE2K
+10sxR+IymNDHGgPH09tVRi+QPOFpHrtzITt2/vKDagEohopujxCMuzDfE+OS5mrJ9OYZhAPhHpU
R4BJB96uzx2qq3VC1hwfk3JlcLu0oM4+FluuqTHMHz37WwYnMnG+sxJEmKbvKjKJ9EXNg5so8vCM
JTnHNZ+9tAImmpbc365eoiV1q9cHjKh62Xi119F3oQfpoKrKysaUp2nT5mCSfwVPeLTGdVZwFiD0
suC1yx6Y5DkY8JVd6J4e9RUq1WDoW5mB6AqEUIBz4nUdiM/Fjg9btkTn5B3EzIDX0UAQ2JpdvhtJ
A7qwOL+FGmM9Lm4hpwMcobIWGwEOqph8J9MWe8kWYv+NIwYDgh6DvTVfDUmAixxAlhmQaMAn1lw5
yqsnVk7tQG6ibhtCQNqQF2Yz34/7jqyocuuGPgJyb2IUYrO2ba/eBLYE+hccPOk6vp5SfbM7eXaH
L/8Ifg4DVHmyMGKMbM/y53xRsJRn1DPYWN6LKQlLVun380di6y/VMhxYWg9eWdtaXRpnNd7dH6M8
Q9mQNJRm9SkM6QUgcmgvWdkklkREpN8tVse0VwSH1FWJ/mDWrG8HC2uOnAMSwk/lXEhBvuNa07PB
HSP73pfRQ6XrYEDxErm6+3esv2AQV0DBuRpkplt4xFmGcNM7ckHocma1y2RqYieyyHB2Dua+k+Vg
KROIEXgy5c+J6YKhyme2gSAjdhW4u4WDOv0U2iPMqFFd70IPbM678ewukxMrySSeVSsxDSLxZ9ez
Rm3Qu0YXyytJonnX/PxRV1Rc/uzmeV+3tSdq0BKdGaXOAwuq4iqBpoYCBkUO9GF975uofj0/NRK6
hW2Dn+KflE0NekacoUCYf4ZFdh+Jbh0YwTSPXd91hs2SsywGdtSH3K6ER2Z9T1jnY7D0VCGiTMfX
FLULT9N7pYXtXrdCagBe8M9kngzDrghBCe1K5j+oyQ3FOGup33KPoug0u+R/ObDZK5wCRaOoRtGh
xXPpqrDzHB6B1klhQdUx2FThyK5d4yC5qBwnrUirUr6VAuzlIux5pc9dpsKaCZPK09R55IUmTJxG
BB7CunXE/Ez4WYMlySPq0buLBwdY7SH5kmRB3vqx9Wcozp90FuTlJdUh3I8u6SRAVi1es50mSTeb
JKDrdOKC4uPE4ijTsMinuRLnJZ32K/8xLQ0doa71nfS2+5NYk0Xh2LjBRomIEk33xurMev2G2kTk
EMffsg48zUG7y998hVoDjBsZwftKrss6yisk7yyijIrLRROq7GJsjF8m5KPCQlLaEbb8WVq+aD73
fCnFjEh19QaDVPoix4ziHPdnd8RDY/Bo3CRleSQM6vqKon7ELfYmOS2j51QWbtPuL/2D9lvZCdpq
+V1H8GNyv3tf52ilzpRoQ3UJ3qow59S2WvkXTu5N8APfiEPYQCP9LAX0xNpqhjBhSL12Vpnsrj+Q
nsITWR0uBy1jZ1uv/Q1bfpCFeVGwY+hNFbFC4c8N4wa7i/9LDUbOfFpdFAMuKkdNKtxjD7+xbTIW
DkxEAqCST1W/Y5jYJBoUYC/NdsjotnG4KCYj03BU30It1JzC1JWJN5wozASKDJ5xTDD5C4XH0KKL
wpgriuejdipvDzPZmzc+awgPCC8K6BqNG8aUw0eHIFgZrQ1mLl13gzQWxiKx6Svu1Dq6WOT8LKdp
u46ItqCJLtCz4+zeOOLkmTMpGtc4B85sZbFT6+WJpq3iQ0tTodykHhdnjQXgCJuulvUEewUpjLRQ
xHOR1cxxNhBi/gLoyNGKY5FX3QMFCj2+672JlzzfvPwgIqb8HDo9L3Ns2OTF/3j82VkdHKoWLbsn
4EWWWM8LTrOpC3Qtw82nekEedDo5AB9qqyGtBlUPlJwO0XNnYyREyE7AvDROl8P2MgoXLr/hk9cE
XF2k7HdGstBZ7kfZv0FFAZLc/PL2ADPk/h2/yaKaR5Tce1tCwKUxRgC0kZRqndnP7xKZvB+z1zvF
rZUhiwPiUPWyoEMyvkOA49xX4lsIzPiKl+2LUDdo5MzwzERFmaWhnXJfwZ8+7Qp8sKSDurORwkax
5HQ+7pQZ1Q+5yJx9ckr6IrMZ3ZFDo5Efpmj/7MHVfiR1+Xf1SgmHwt+nmLou6Je8jEDCRZi+3IId
rpqeFekvMKshPEQPHcLdGG/WZaVWZaD30yfE8SbpTkHtaYmB1yr1an6kDmD/sA+FzvgsOzeDIekQ
udqbtxusS4aXGkApe6tl6O/xj/VOya3Q70M9SR4UhbfV79Z2C/nIBJ1j4j9BIRjwB4m8qoLadMFY
lFS8tbJcAuhXVCJ1k9i7VFlii8INxEeSL+S58BhA1t/JrPPAiWU+G5gluG1KbOG/pePwD4auncav
/Xssaywgsnuy9o+aNIXjttuwJlONiKyLaqjsHWo5Q6jPEHjKeZt1huhLDqNnhAdWKBoNHEnjUQHG
pCAv5ez0fSm40SIyPRDtqzSCHGcrPCbSuJhyLHRIyoYjUEBl0hoO3Evw62mnTT1cXkw4VlpZOXbT
Da3sKN90E2TIDXRvmPm1uDMD9KwwPABHdjogB5T/T2rbsxap+4zonAy34vTR73HS5tLcjJrsvFcp
8/Xt7kbeH8KMdhdNIC8VVB3a3T6ZTlG3SYPS4O6lzW6ufiAaYdV5l9CFUY0yHjjOCRpVW4419qiH
tSD2Cqp7SEfm89AGfzCM4DKpFMXlr+C8XruE2UmWHWWW/KycM3V55+4eT/kKHmcSpvzht6YUu3pu
0qCDxY5SVZobXrdv18yTP8RZUVy6Ye6HQWJtWGLTDXihCJyYa6hSXnTwt1sffvDjuCUwb0E/KXdy
K1iU19I8+JnWWbvCBVItaB17xLwupXo9z2NcN0wjdFe4Vb8iohtWcMKvmi9zIEKJN3ZmeBaItlSz
URJaY2pr83fQq7JE/ZDYEWPe8yejn4sXiyCCkwtXLkMHL1IoUN9t92D/VhQw2vizYrk9eVBb5Q2d
7CoMIuFexpjbE902Iu4RjjDVbdZpFshNJgVX5fNQ11lkUPVB/p0nbvVUImCGSb+ePZAveBhrb5v5
bOjZukqC8Szie/8KhBO3iUUo9mvQy1rYseLAR7gVmRifEvrVXQBJIZvvRr/6zouHqTxOJEC0ofV0
8PVoMHmtJAwdWi8qlOTrG2EwIG6wls0QxIjF2eYgxIOI5DcF937yOB/SfdkdfE7203PZnmHNdyk3
Ma3dlBJUerGi+mjcXuxhlkYsH1dYk28CeBT/4ZDcjZX958S4nVqyDSLQA8JuCc1uE+8XtQaiBi6+
LddmCl3+U4BfGkr28KjTizfhpPr8XvdR7Lr2FYHIRS0zuswA+Ovvp1YNCDmIrV2hkVa1bWWn1lYq
2YuKT3ZWesCTHsnEiUJnytm3Y1n9VFhglVBkp3oSxY8d/QkjGUwGfoPEYefOYHu2JgGIvXg6OlNT
Gud3nfDw54MZFx9d73BY68Z4c0t1N9iWOQRjRhbmUzjAlNe65x194IQWrfEr8QdjOYtXYu1kAJYb
0IYk1UsXQUs8jChdLOaPZ1hbYCYuavGQJjq38wpV+RlyuWp91IRq6/W196oxrx/36TgtYmfOA80u
v9x079UPw217SMdezHR1XVnWjXwGJ9AWHl32E+PGHYWbMyLct/1yWeiZxA0cXLb5O+iMts2H+J5i
M19RGs543zHLE+REblmHU+MSU+aH1lwArF4oojoDWwOFZ71IUMFpzH8AXG0DdMCPYtesKNWj9Xo5
7/auF0qDF92rAb8qheJoJQtuHaBTlCBnW5jVr00k50lWw+zP+rZtHLCcj1acPQBTfDIPUr8r6pbN
1XiqfdS1J4/xXiCE7j8+wfipzOKNm9QmQkCPz6iIeK9jWcdD9gf9JB8VbmZi2oq57F/SgOTE9IUC
c8Ac+15PFMOykwkC7tka/pcpZ2Unr/ev9QRfYYd/rk+CiKURbsRQZpMWT/C531aAnwcqerkQP7vr
E3cYvHSORyvtr2KPKcX8sN7VGiumvxUDl/OSdU8KVXDLLrwoLwkHAxFR4YICaYXSMS1/o8PmaUCK
Z/UMNwnn+gipZT7MGhqOTwToVb96OQh8U+px2wCKV2HSLDjbf5RV0zJ9zi4q0EI6Pm8DvIKLl+Zr
ftYIspJg5rIde/qY3zkeQeajQ6DhJytd8micZ50nf6NvvNYX+ECYb3bSPrl5f4qBIRft69PTkATV
OFlas2skAG4VXAiA6yQ/H6TTcTa7s9GQjiXD7bSsSf/Neatu4JQJATAy+EOdC+DwAvw1OcazrplM
8HCz/AkBK6wQsb8ihGWu0XFYRYuFcqSIzbsRlPo1uAnOLVH+0mn9BeecshSQgCqsU76Cd4p1YfGE
OSjQgiK8fK6eEIrsAj7dY8xOW2VyAGY4Z5nXVpnH1/uQbYIEP3/xOUKzQ3ha3Ww8XysdF3M2hIe9
KwHs8OmAB9xZcGAliN33jQwiTxHPee06hcCMoIMS8CNo/NelhJWHqq5SqenuVVSO7XoE07Jo5WYU
rzEkyoONQlnW2gjbEDYzSG+xb9KllQJo6DfCc/7/lPgr0VvQLeLI5VnaYYC9DwdF941RT17Vj5VH
OvqFYYN1cgskPH055195lpJeM+LOTOQ8KaFlvYFoRGQeQrjEx2sUDVY5EdWSPZQglk5azNjPQsxL
MX/ZwaogpR24FlU9/mKQIjZ5f9BAVMwiIBykkegwJZshv2vlCWyKwmxx23re+YXDSRHCjoRLmQxx
OetAJvPhM/LhMk/ntBigWrkczUWBDhr6gAsNkD2Mqyfai2np2pW+iwbRmPg8MDZKc/g9GeESnN1W
ss/7U87hXLZJMt0DGmcMPRnOQjgt/7sT0w7Fl+y2a7TY+eMeVneKWB7ioZXsxbD3QxfW057czd08
HxpOWhD2wACTcQM5cRUc0EZtI7aeZO0KHvg8CiiwgwBlEpzczUmd0flCim8PbyaTAUF7it1g7RcH
kkZsH9/WTMabv631aJ9plpG9vusdDQqqR6UHwUFn0/baij1wRXVq6RxhqNg1XN70ahcOw2stT+/U
xkVGNJl6iJv8XTRKIr5bMXUNdFhmDsL/7WMZXnM6V5ShRBQqDusWVCAEWj0j+wPzo2e5mgLndBEP
8fIl7OuI38iPkpsRQ1y2ML26OpnbtKAWy73BT7A1f5E+ysyvpGYpxqOlkezYcxK5ILUpvq0WbfJP
eTYDKxQnl8uphUGWVStQZPJj75YYi8u6uObDTWVwxdLmzW4wmAnRXzwDPG+81bzFeEGhyxemlsnU
D+AmLCV/0SRyUt9QFt+ULj+qrxkhtjP0OCYvMGe1oX7LiJwAeCrkipnr7s4UoDh3hAPQCUVzHkvJ
HgFWzgTineVzNkpoV7Lq3A2sPynNeMtmS4MPHO1IMSy3HZvtBa5lgmbCkUjuimdzOFlrp4bkLpLv
kgwUzqVpFo3+bkywTOK/hF/vNxtudIsPX87CYnB5R4cVuMisjVqOoycjVVO4JGWojC5Zd4BVwFr/
jE4Yz4mMrz0pBllxWe8rkc0igOUw+2AdpuZnMRTzdq6Ou03RhhEwpCmDIFd3PKVygPtgyW5cRSGl
w2b6IuodhF5zwgllhwPcBBikhZHhMA8xFQMNDI5Dq9CLJ9z2K7RY9fOnExeuq4AW+9NPog1TlI4e
b13Mx8AVQOtE5X3g28N5lA1cEtIXDAhpqyylMklUa/nb+aM3g5TqVIl9i6ugj0Gjwi5tCOiq5jKI
4lzmORbEUfvl6fovHcMA68+xHl0OKnDbTDSaFhA3M0AZOIwh9JMHmyv8z/GZv4dr+fP6UaV9GXz0
Xjbe3OE7NZUFwjV2c8bkswEDge89eGyo/q7Pxj1PAe4L5EFetW5UHzJQWwvmceIra3NuQ9/aS22R
4jCYk3Q6ib+saZCM/+M2Jw6W1CQzcYldsOokD8UdouEA/5OMADp2aR9tkFVkKj+tEXGsU1YJHHiF
Hd8nWVFB7W7LHEusSn0VjQkgHi6jzBbIQTb68QtX3E3icTNYfHf2hiwfM5X0vySYQoUNBfS5ck8/
Y5XdfpS02DPZPPPU4CAHoVe+kiWnFBuasjA+RmLHKKcl+NEE/Ldlh7PBVEBIS13Y9me7RZnl3G8u
CTAFipNgbjfns/pd9/BFrQt/5IomY+0iLaZYjVRY9VqCvSiISpdzlQ+Zwczqf0mBu8Ku+sMNzg/c
VtYOW4vKAmjrnAquOElvf7Ng2cPysJGDwR8ugG3NoswFAph2mftnb/0VWYP8kDYwceLaKNpN5gMh
j8bVH0cgipx/YbXGCAhIOujwZPayJ+5ZLmpP2029+LF7f98r8CWKYRJDqbjd/ro2rZjfvhIduyZw
Gnmxy7/RGuFBCnn7WuEufktYb4hjICmJ3bEwxKPAtsf7ulmo7opH9inv21v9LH2bv1ktM+I94tzd
MIBT9xqpSNRBXpvBOet+UW2PmYULCEmkUsTN3Ir9Vn76Dp7dLjkXvz+RLrEf0DBsF6EBGK0qJRxx
MDMaMLqctlJJtKUUgn6yNozXEslsMBS3PT8LdES0pyexBB4zP1cxKjmWfxrHGS5LTbwpiJXS83q8
yWlYjtzKUvMQSkRo4PsDR4dm9W9JYexJj/ARPSCdu9U7MlWDXJq+sEEi69y6K9o5aNgKHZnh3CyG
0sRhHwnZgX665V/3J38F8T+NhTY5wtqn6TPXjuTdsla893sVC3ddV3fJGwHbpmuZknVtNgvKMdqE
9eiNbSBJhWi14TtciJD71F45jSvR6RIGDyfX/TSSM2cJNWdcvSZB9dltFWvcFa5gBQP6ThdXkD4J
cGQuJtlqi/Tst4b0wuJ74f5knq1nhYgSNXnntcqLvkEVWAP/hxfeyiBEXXZFnNTPhIoKnlOIlrL8
81sf5UjMcoWI7FBhH5+x6pO+fAYw5bIygir+fkNkfgMkcWBxTevtV1spC0wvKG4b0gHEChxEy69B
sq/49mZ0tFZi4342ZOsHvRTVfruIisEJaq63qr3HnlRE/wM/oRD+99NsufPrPnekrmjwPtLrD3lr
vq/oZQ8cn0wH+w8hEni1etEDbDT1oA4gRmiSVyc1vQD0aVloTYe0E7zHxibNinHbmCHYQ/wJhb0L
bsrMNgCYIk6DgmUSi4io1kqh8b/UVY0b3j+HxKQ1WA3H1M5g9hzCygc+htCPs2uCi4YEuuvXMbrx
e5b36fyC+RoqaFwoUFMfhvE6xBy0MDp8LRxYWmydku+HvdIRE3QOmCReMPIee471+8snaxEvOiRc
AJEK4tBYj1JkcoUSjgKs/0hzvebzsPBaesSNeDFu90lNVQBLas1VJ9F8Zl3wdfpUrq95fk37KbeN
gl/tElqOHOkLJ5lot1O6TsNdb8XGzKL9lCDZIKPl19ZrDFMv9S8o2floJOkyJHbkY/p17YH4Z0S1
bi+NK+/S57WbTxwx37XzrzDOvQHIqhyE3b+QzJg50ct8iFUh3pyFskiCDYKdmBsm6IGL0BLNlotU
dBQlNml92KF4yb65j/1P9SIeYgbpguymFsrJRDo71/jyXcmhtlvbJD/fSFSGJMjbzZ1hZc2eBdVj
t4K2B1ZVpm7xVTy0KnLn7pX4CPssNqOZYC/mJnoFGs286n4DHmrCgYkvv49C+qMdGRw87/Hn+vMA
dTlTtVw+mL17TaD6/ECbw75ix9tkEg2jWHnsE3QF7lYzM+kY2WrHrIJ7fNExjczs/ljQpo1oOQzm
rmw/ATpI30kPk9WnyUEQE3Z1pMqdAFEvGf5D2Qz6Obd5JMgpv2NoL3Kl9fl9sCTY875o51zM7dfV
UKMY6lXmueCdawYUSoTxVFIi52GyHywSXY/WwLq5CBDDAmZj7n5KZPR9fCiX/KCcyqBcJmj/tbao
OR9INlXQ8TsgebFeS0jvRGGOQyznRqJllxsVe4Kq/HY5fMlwt/awae0Pi3z2tafEv7cs+1Ne1kII
PXKNQFAFCPL6ZIXnwND2KpIECZDegtJzYkjFmYJj1miYgIVXeTZatQ5rrGx4Xtu+6+DDUadN8fII
NTXOJegAlSCiMLt6UJZ3TMm9hgh88e+KcantbwsceJ+hWk9rVnw2q9kNLc+crgeWBtV4SUWm5N7G
bA8z54c3Pz6xAQWX4ce9SoD6r7KYQ7EUubx38QTmc0INGKRcOUq9akkmXe4fWx1xl+pKU+TFitLP
j6AC7sTRXBDONR0RC74t8cb2btrESrLITPDrYyLdQtKKXJZAHbC1ax5Q+qPyXeWItkP02V7njh/q
4LX+iiUPJzQTQSa3ofwYv1UuhPgVqcAzEf8ZoW1y6A/TFMzuwlModJBPQxHJ1852tDecsUP2G1lW
f5Lm7NmNqRZ1KXGOC31jh7d4IymqgLUyBRXORG03ccBkNvaB5FhvytTpDEAMWTtv8MZzWenbAGvd
44fuzYIpOsNMwUaqhdZ/xFxJwb+0evFu5fIns//pLiOSGuQbOFks9XdW1cbCa4jGcCsQ4UlsqIpl
IU0UYtQRXvl6+0vO7neRevlxwM6zkn1S8iEj6noKe1mmK5cWoDdpKkb4Jf3CX2rVbm0fyUzU+bLM
Thkt+qO9lcUT9fEYLJrZ3nWiziTjmLmfO35EgLQdUFgr4g7OaetU5Nu7F6yi7S6ZMgmyN47JB/h/
7KM5+vhnNmg2xSW+01QxaT/APYxYepA7ZYvS3qOwISqFgjrBxOh09LtO4v1/tuEW2U1gcfahcObK
UqOyzyVSWOTTOE4o4JCh+mdWqVpp8zIAdVHPiF+HXGko23axFJZEUj6C/ddBgCWbRZCQ6oXA1yhz
TZcl77k/FjU7CND3p0oHUL530ppAO3GmKQR7mdXLTP1PTc/WcuowrtWx5zU7rbhN4GolNhKGgKAQ
9rQcqxlCurUfig5RbOpIGxsvWslrJZY5z/+kc8LIu2zebzQDgVPflGCg1t5/jeNEdEee8IiMWmIl
aBE9vzWA1rE/dz4UlAAWt1LwEsEGmWQVlZZmPvTm2Dc6kAQaKx5cf2Ria5rBc9hAW/KCtH+El+TT
OKxm2WybyeUXOnWy74WDwUJW7fIael2LbQcPgxOkCM8tX0d3CLWiknfctqq0x6YQJCD1H9ihZ/jB
LCDVZ/CMgC+VMOwVC690ILIB6CmiYNFpS69eIRQOXziYZrAsOFR2hZVDWqAYTPpaBoQCtSMeW+Pb
ZRooCLl4/y4RBb9LzZtA3hqbjxBlSIPhEYwXatpdqE8vmqrMx6svgLziMYRyRQZbWVPlxegWwsvu
5SX7gRQNXPx1IatRY0NUOvjw+rvkkSwgdT1o3uXGjYte+r+Xc9I/v7v8t79N7hTa5qClPxtbESPH
ACNmY/PI2Nh1kxMO2QYfaGhHFGA9TZr15VaB+xML5arUP8vO5kFcsMEqixm90ggvCxSBHxZKf891
P2SX6MOtpbm/c+AYcfm/vFOTDyu7MoJ2ROtH2Z4GQjHwT3/1pwexcMdUy3WyjQ73yiPrtBa36O8+
5U6re9bfZ86GFIBIsgfqCa4see5KaPey7CHuS4aYlPCXZBloa0sTd0Gz6RLs6UaFLSEPzKyS1IgE
iRcFq/V3HwxnV/wV0cGwsGboOqy9T5PSkwoviwUN4cHQxoaqKA4HHFDqQH9ZdSak9kZcjGoVhJc4
ZLi2FFXEPEfh4jIoePefMObKS1a4ZVoYfAFwT756u8bLjgRljq231MNVaoAfQ/4Y1uBcGjhCzRxT
6gGl4PbH+3cG1tH6nPvBAIQ/nh23ZPxX/x5rc9BXinVjKvaJq2kgm26N8OnVDs3Ko/IXI7XuWcqQ
A+Eu44VWiptJ1UXiN8S55xDiveHKIxfuDRx6BxJlAYbY6xFNwDijGgfXQxL+nLQREBVJzJ6SRKP4
YAz2q1c9oYDq4v7ZAf1DwMeJ/pMNsIdBnHcSYtjzbJXD+abnPHOJGB55r3T86eBijOZJgaHdrE0l
YhQqG4SptxIczUm3Db6yq5o9Wa8ttaeB+fS/FqjvWHiOk62ZQQPNUZ2pLFOkFUdRaUb0pRBRlMNA
GGd8GecmgFihs3okUrZxRHS9c0C23AbI09KcoRAmyC00KKPoqhmS4y11OS6cIoIk0fbM1eiipti2
LKqdpnzLKHD/KDLz5s1xe5hdNPEf9uueP8G64hMNbEJ2p6LFAsIODXdZhemZ6o0xwY5jhFSVzqe4
10DaW+DYB9ke4kvtazYWKB07bPmMcYZ2dcP3rudLm1DbM5L+WXPQObbxhqW4+O6reM9/9ZgOSEgN
81EosK25dOCfImYPwjvvh5qAH2O1MgvAbmJhs2Br632SlD7o3C1EtxM8QA3o+s6ntmzTk/5SPekd
ChZBrqg8zhU857j0JGDFvOFUyQrHTqjnuRjmX1KRdlhHYwLRxE2UQj64Z7+OT2vAS9t9OA7B8aOj
eRG127WdyQZjKVD/oUwy0A6U7aGNX/jjRqFhDHX4OdsUS8JYp5Vrlz92aWZIJDfopctvQn2Ym9Fj
ZcjXY7jkVCt0hiiJ4DHghZYYdc9vdVW9wd2moNBSoYyyw+OYbWPOk2R4tNcpKs3Agw4AbEkvbKOF
aXY13NeX4yME27YEYyynkDvT2mSncWVPl1ctyEqx/fMlx0Frms4v7GY5wxm7M2yc9uk6HQWrJFwI
lgGIVdE1fqsNmaAHBy7zcHXDApfH/pphBM1tCG7FMHeTG05y9b1Q+pQR5ONgJyvJe2r/kxsWZn/+
/2BIAe+YQZIoA8ZlLYlzdUewcVZQ5Gd0oDjaIA+98k3vI0nsKnX2kKVJ9CJqDK7TmUE8uqYmK5Sw
S9iGcjbVanKEeZzH8x3ias0hT58FL/r7LPQ0VywQlftcPINLI/oKl9I7O+J8V2t+9tv23UBaEU6M
mau3MEbSqvHODCMko2LRal0jkiBZ9Rx+4L1RUX3XQi/iwg8ztRqEN4ctzVnUV6y9HGQJ/pg5MqZ1
QTaHJwDDKY51fcPEomZqQJvY0wrPHo3Mhp5ZrXRfIrq8HTZ4r4JA/tDaMoCUHSZN9l+bUsBwXJew
Yi3UJwOtqGaoNsALyWOLbdm7oFBbA50jn+22dxnekz037Nfu8iw3Y6C2Db/tv1fEW7sN/Mog7Wz6
Hk1uV86VYPKKgRQIULi50PsWiNDN7So0OMRRmfi2pVJpnGbDLHUjBQocOIt2JAfhf0OGULq8tbXi
A+WJ9FM1gKlYy7LIvdYYeHFKHt5tvR5W0cdk0ntMAe035qIjXpnNDEqZdyiUl8CMTSOiuALoZpZ3
wTfvLoFQD/7phru31lUywC7wBQLKDOA/XkMkbvgXKfjvG5TIvmAcLz49+3TQkfWLq04D/AAUW+AK
zPcoWdyAXMjWLYTfNzyzzKmc/retAAalroqiG8PdrHpFMva/1ku1A2X/fAaWc928ttTxdaeeuDCN
ll1Ri0C2D0w+xHv2FGWn1rujHtb17BdbnGxi5EpWNa7kk2rcg0cUZ2ta534CsU5UG9JtBxTB/fCe
p+epHWkaweMubMT5RW1eJo5NGk9VhFOa5mRsm+pkLrT5rpBi1Zy5ckiJSgNk/M2a+7VaAO+NACmQ
Hy0/nB08ddV/yLCmHUZM2MpbCuYNZD5CLkGyv/YDDnaaoBPih6DEGem0OfWWkLFd30WTWu6QjUZr
VCksNPRqMQnFWf0OHqv16F+yFtgx9DuTjfCdE+1wSIRK5krmyhqGdDfjpVye/HdqnBaHgXZdlLQ/
aIyRa4kgBWVfTPidN/eqPk6WIbEAkBJOQKfw8ANcJPzS4Pl/h4C5DrKwlVPQk33IhtKqdHBhe+tu
Xl3N7ZnnGsWTyQLZ0C1oOa4fwe+6wXdlGed8dJI1C1omoATaWROAOhmTOp3M2vD4kjoWDOeOjWu6
vUHaWMerncnZwGrU2z/49wPCsguT4nLKDxgGAAqLGmFTZTPuDykUtYY+DGr8y80Q+F6ymaKlGmo/
+mQ2Nz6NMjHDnocb8ehU7MXjjbVzffupcnAYfjEUUqAMbwty5wBQHUMt7nlMjRjSULH7S1zEsS1R
4tuEhjS/WQskP1qQYbvT0M8R2U78adaeCEDTcCyawyWNTLGJmivJ+bF8qNjOTPo5RexLTH1N/XNY
aVIskEeHDIJMaKQseTTjd4eoyj4qM6tdEB4N7w00uR+zYR0rJvJiypDo1RKCr47ZpuA45U8Vypey
wR5Gf22AXKqkS1q6NMtOPNxfq/vXlZZDhM3NcxfyOvHK45vaeWuO2RGeBXD7ElCc9gStq6It6RdF
O8/DpBHnmGcLp5/TNRBtz/ninVIst/VZZ5qrlNpor6SifGsPw84FKTblbS54JZC9rpaRJJ366bXn
8jgrksbdcEXkiQbEnZA2fyOH461KrQ/O4IakCR66QVDDJ0scZcWrxxJe0l4cNrU4z5ip+/Ltxc2j
LkewXaY9UqmkSU14he1Xnr0UHJOyRT53P3XQl6CWTRWM1sDDjw/dojbb0kgmSZPtMfjtgOjjVm+B
1aZeEyQ2z8FySgDPr0S/6U5271N1fMSR0xhKkx9hZW8ohZwxtZwjSFzIjH3lTGwba8o3drnq2sWA
0gb1T2U39RqjEm9Vl6t1t06PHtPIrfUkGRAMkh4N+/cnPc6uWqOLuXyv5uJdEvO2kkYf+em0r7t/
XLSeW2SJLOYhD27Ovu/9YvDVYKes1XeN8NHWC5uMkk7AOwOQwXoRawLVKdFE5bxFl1qZDmdO6l3Q
wJTRvSSlQJ63OvrI9lBmq39c7nJrapNz0YeMhx1dkOhJEj0LhV88exbGqW/C3/0eLw/2r6VByHSc
KEgp5NuMPS6cpz+kcIJNSv2y0UmZaSFQf8GCI/8m/t8LLCFiyxBUR2WBoUIZsrGMMzlz/NRgkgTq
ncYq1yTkhzYrsevDuje9PVu5q89dV8Td5eg45vakx+HOYwwtChNkPBFOw6Ip4SwIrbJlISaWZ8in
mTC9i+qyNsugGSfoBTVWXKz2NTjyXj3mFdq1Z4m/JruefTwYyfFUzx+6dY3Zay84RryHZzFswhOu
WtlDITxYrE95KPYHa9i6qzd5AWAYlvjLhFg6FQjjj4LNog4zs0xLonTSjoVVc4k6Nn7MfvWskFzC
noYTTZ347gRXgetW5Z+jJP1VzBVmKQRHhPdi2morDQMSXMnc5Y8ffaoj2Lojm9mX3RSFNuiu0Yvj
eB0+p4Cz542ug0RaPfspbAJHlIZZHAxxm3J7k/57a+fcfudFRLN3pqPrNOEjNJS+LMXLwF3IR8x0
6wrkBS3Nrlge9Ng+XGO8kQbNyPS8ffhGOwN8GQ2/ViLf7a0VQF1uJBXOCEHN3e5rw0R9Poov2cg8
emWYjVXn63F8xGqAHES8mBKFTHDTw/hlOskQWizaq6uMBh0+E054F/AgwMzBJbKgTfKF7Ug/qnmK
Glgt4E55qS1/dEKN/K4n/3hi3MGZ8RNpiOoz8bIo/P70RyT7i9MhVHRc/wvSWENBgFAIyXcYmzA0
P6njCoJdzIHvmbIYkLMc71w36fglrN0SCV14YTSvHyvvIVbbKkPp7UnvfQn6eRWuqlUA3GMexn+r
Us7DEt00RhokoeO46zH88M3eOPt3nK47jgbiTBQJJbZ6S+Rc5yw/WVU65FE8YDIiQBSCS3tDNF9s
+UUfucJAUt2O6SyqOnBfPmTW9UhV/04heINPmHCfZenfqenvRfuYrQ/IrFVjo7uj5I7Nxn4Yro7j
au9tZ2NnyHii5bf3ozEn+BOp0LIzuYWtYYAPWOVODryYwAJ3oZftOkDsWGpSMaas8npLfZMO+ZUL
SAdE/pY3eejRA54PXtE8JtOURf/MfakvOT2RyxejmLS+Z1N2FO10qvk8OEqMI55OoSM+xpRJCmoI
pwKCnwMoGYfGc6nL1IhLASTgVb/6Bbct9Q7UTqWFuMNZSM1kxCyzHdUYSE/9LIXAF9fkvkfNKqhS
GyTnS9maVOdh3kKzlhDwhsWTLgMnKZP1CscR82r3Mub+JTwRFjw43eMGbbDjbAcJi6pYLhjQfHeh
51veWSlTZcMzKNyMItGb6sbH1Fc+qprSk0JwpfvcGUXOF0f4DFLsTJz2ElDMf3zQGNSFknwt6TzT
1rqFKynlgLmYE+fVEL1xG+G28iYuUsXApHXAaiENxkZSUQhvS7m5r2yEmx3XPBZV10HDaMpTvuUH
Z2l8b4hxRH1UXUMZW6Z1uLp68QBR/xoq3kNk94W2B5Hna7rDGIQXlmH8q3gq7GGyPahId62qvlEN
MnpxRX1FAP2yMeICpug1K324EapkPoxnZIW4j5GFTcvpock6i4uQQ3fqeiyf1UALQD3dqV1eB16Y
abixmDSSSGDAoWO2ZQK4o5HZn3ctw5/xNtBxrahDizN0YMe6SAmzzMVSiH/ALz5uuBIcnJCQAOCR
c775JB30qlBMgzylY8NiwBjYTghvvyaDP5HU5siHlVsnn2j1T6WYIc/9wPZ62KWDtAoia3o9SzZN
zm8bD2W0z+pRARc0eZ/P+dNWkmpyB2PAyUX9nEptY7UuNvQrXTt0NQRV0jvXU1cdbmQE6d+DcGkt
IALp3KWV2WTGgVCFj+FBnZ0onN5V0qFP1sME3FFhGQtH7l/dn2kbZLBueZV5ddmXXm7ZmG/T1rfF
2OKU+iFE6PNDU2G0GgTco7eCVGTb/h3RUGMQtH+nNH+DCghxqLpLu51DhQ+LjVNmnyP3NXPyVO9u
eSpHqC4zq+eGWrgJdHWGQ2e+MlTENZr2/STycF+MoYL8r6azmNMhRxepLDuTLGnMTltlG/HEUtCd
MSWFsap9uf0Y50il9Cb47MY3+mwMPatF2Z+PYKzg6BpYUEs5edKr3Y5Zjx5jPRIHQHhMe6fFkdA/
kzewsh38lXsWDsvoNHkfYz2hyUeWExz36f2M7SUstKZDYld5LqN6oU27PeOLW2jfFQMIWGo9wmHn
LIy+wlM58ogHzQaQyJBLBfP4X95LmOOBdL2EArd6oyNj0uWEbx8eUhpsNjRjlWZpB7EuQE4ZIi7h
MmErMoMl49Gg6jtb1LDaE72iDy3ZeGjDwcTnHHRD0fxIq1R1NhQWF3BEDSqWBynNwPG8sa2UvHMM
oIubcAZTXHx7yzN5J04ltyVmU2xA0GCaoaBnAUQJRw/qLPBxpJ1B7WpezHixK6rnjwXFln7nGC83
As5Z4XQaNq6RGljFqztE46bGdD4efnipiYKtvzjjS20iqoabsMXVArZkWBtRxsoNUYleXcdfVc2y
jttB7koyjFiS2tCh1lGqvoI7KtEpRa83hQ5IxpImJcu5uT4Lz89HsKFyjOjQoVwIj+Dc70V5t6th
K+ttayQmZnA1JPDt/FWlZpRbps3S39Obl2s7v45d3/iBFoxnGX9c0PdNs74JqZMQGX/BXu++NQNm
dADp1uVDBVWnvJa43yWOs7FKtV0uOzXAtuBADpU8DY34HKYsQmRiT47WB6yWC15d2nlRY6etq31A
dEqibJDLgbyxosc4Fv4ZLWMeZR7O7Fk1Ew40rNFqotg4l6QXtoBAoml/O8EqFC9k/hSnLPFoMAsI
+qgECAabwJkmCFR2oX+r42qDe5smpT+jwfm7eOt69yNvxwoms5LtbKmXvjKquCkBXtGGkKzM6qiq
vTA+ynRZKW9VA0i3ZI3pETDXWVpmtQtbLUrnNSNY2jmHw6cbof1KzQVYAd9r4VzABZwyeQoMFZjD
HR+Eb5xZemLoTV0q+ECtRPZ7/NMbop3KQPjAi6mvPqbxb40NGaYrFOn1dBY3ydGUw1M/7T2UY3yP
kXLJ2qFq3lmlxTD4CNA50TaPpRaKFckhV3zx7/u5WQ2SBtHMeCMfgwGufeLNL5ohTIvSgZJixsYZ
51SvGhf2SbUA0ZSPm1xek9RN6DMNnWi96D16L4V90LpfValIgCS+VvlkT/z8/JMj3dNWNgKF3fUe
cYHKjn74kXEPhDVaQuCAskSV3FCCLirC8LEaM3vEapOXoFvRrp+u+FUyxMBG75Vo3HuMEdoCA5hF
nwQ+nIC704NEI0TI4TpRN0RhkyPWiliLsag9lGvelMySHGHxzB7mymJbSNUgl8Cgm2Lcrg2mi+e4
A6v1w6zmmdYdmOqNowGFBAcU4GGy/dubD/UYtup8qjBwj+Y/LfUR4WgMECuEonB4GCUg/i9ERCSj
izawSIFBa8s/FHRAe0EOU69y2O/93RjEY5f+QoYFiIYOtkAUXQB0gvElBLVDEIY2aQNKHYVXxp4D
EmmOZiOwc7TApe07SlDOuJgyGlR9g+dGEYMAGvpPDjpD6B9n1mIIr90AXO2K5yb/5ugbhWEJuRgt
iIVzvEvhLvGCcvxrfEvt+oUq6isjiGRfDHKqmZ+pEzMegXQbk4DKjCJdm0+lpOPHiH4wOfAL8ZPC
bPr30WdcWygkH1xoS63ri6is8GwMIMY0li2CLwirR5az72jAa7BDcNEJRA8NezvYfVsGwYociRWn
69M+UunZdCNtYcdY6iiCUjdWL9fGGbG6ibrH6Ex7Na6MKBARcTD8+0efQOHH7KE8uzdMO8DlfL7I
0PW9AYRL9VaEY7fSzQHsU3PlA3gbLRL5cC6oMSuGG0v2/f9mznnsBLQIuNnp0pMyjfCY4kKMRrIB
hqFAo6R1nq3psziEzYNXIaJ/Ha7h0tl7GH2v8VAOSFPhlNREzhCCyuFInI+A5B1wvzHTQGk4MjZI
IWjVny6Yv+9S5NbO/AvELZUQbOdCyqI4m9gWbkcdAB5Vf8jr7eq/J4IzMWvstrVLMBDsxTEeV7Iy
WK01sisUpU8L6FCgofRPdsQ/iYsMbpaCmN3KBp5Xh4zVdVfH0JxT0IRfbUuqpyxYx1Dnw5QIDaym
77MjK2ppNr1hUXx8xIGgh/pf9V3TGruuV1vqM475anqK8vqyHAHjwvCzM8WkOpZORvfE3p9Dbstr
xkZjhT/zL3Eo4wPjnREOXr5aOZF3XO6rW5NHfcLM/kFvHRdXUDsagO7frmaAGC+Wj4Brf7cCAqg+
2dVti5Eq5bwGp/3ZNe1f9jYFBDrGZRZULuTQFr8+bjHU9d9GK24NqGtj/Cz/j6v5pFNpw+6h9XoD
ZOvIxYSGmcloc9NipaXPKsHvcDALZ4iicvg2HUid/qkyldWW/wN3NALiFiz01JMubJf+EknxaanA
LkkiRmM8lWm5kI55CfCHnMIf27nfgjxJ+fAyNq5RROPAHwsMem1MPw4AkHYfffafCHQqVeFheyfu
FXf/2aMR0xxOexoHtqV2h2F77qUUDucglom/8lPihVuaY2P2nlOFcd1oYcvwY54g8JE1UNuJnxjl
SGoSj9ak+2r2HkKpnpMsQI1o4JJ6xfzME8xJdLSWkN6aKM/fNHOdqfWLwU9FSXoMyRhZFIEnLLis
ixbTKExuRLpDqCvRfVfliAt+YkQNb/X0MsGYIcuAQqopXFvfxjQZEKFydbAnMuSm5NJHiigot+ws
NzoIU7WD/6VnmdJu+4Gex/jqre2OUaiLJZLTq6KPEUWPwe7PzbIIzlBWDvEc7xBdl6jRzNKLP4LW
oTaCyQVsc3wRfr98461nK1w/GszuTvZ5N2QOxSpoTfdZnFNmWMXX7AQrSECSH/Oi//qiIKzs5Qwb
LYz8Xkwrs10AcnI+Ay2cQcTO4nG/FKHRb645R7If7rHTi8aUDLFCI8LnSCVNvTG/Zdl+moUUzlm1
BjBqEVfiYFZ7dgXGvfKvsvNsODtvrvya+sNIvagEeU5hb/YyrHsaJkvLdAfPt/lS878lsFzSW466
SdxX9RZecbkEy7EFeXitlEXUfjiast52kTnNhxIf8Wu1eECnWpz1gysmPziLDJETwG27+rhAW5LJ
BitLyPi3bDuEV4tUpS8M9KjsR/zyITMkz2ODp8tJDoWAmsKBDEB3Ie2dtRKis3ez6O0dl2cN7Pfh
Cq+F0LR+jwTm2FAeTWAe4OXyu4fG3rw9zZ36qtnotV6lmbInVmESYOqF62RbKLNcoeRIDGD79zhD
tBX3yf9409udvPkzRx6+iijvcmx2AygD/Cc8ok/1PEpwp7PVNYzEQeTeHsMA6I/H7gd8zNrc7gwl
aiBKyqL0LSS17hq9doCyT6RK3pCqlEkdaQ86E5fa9epguyD+7Noz+V6rWIJ15U+75ge9N6f1psfO
xT3ThsfJ6cOhCP+jifl2dHXjFwN5T3za6lvs+fTCSLgjzNCRVJzKwka/fm5wrbIYb/vzEpAiFtI3
SJwT7xaij5XbYvM/pWBQxfsVzBH6RbyHFnXyi7pR7RG65mS8y2nwJQXHLnAjSSoshHLzJyTZtxAt
Mg0ZetH8IQGObtmwgho9b0/1Y3EwsBjG9VWGuMTbaHspvwGwBS3sjBt4inCCfbz0GZhDs+N5cIsv
15Oz/9t/LicgQhgEdZttpNLzV55SIFRRBtd3G+tNA+77Sg+dj4QWDmXlv0+9IdmZSFLDK4cLKOAz
EJu93Fq+Az+0sRnCzUC0ZXIvK2qdER0ll84iHIsp8BnJk0ZS4GUlLmZbMn7Ef557l4297GDe4PDd
CYOIB75RUlyEtkrH1Cx4mbAv0X/dHMEj5IQNh2vv3pfe2E8P/C3opAQ+7cAOrPS+CLkCDFQN11yW
7G76PDKjVu9rwW6DX6NncpQlKZ6fn1VoADjMZVhBr2nU7MtuSZm6lfi/G9aPvm/cDtnc6AW/krlP
VzVnA8c26PLt5GVV+q41bNktgs7XLnc573MSw63CM27dQTgdt4z9Ef/Oq9xYfm81PdkA19Xdp69L
vWoFyxB6/tsrM/aeePOshJHHe3MmBOaMNYGxVToZPmSgxyirJ25M0YIViE8YajGHvhUTvbapvjYm
vocktC2Dc6Z8XmG1Z9ULm+ExaSZOUrBJpL8bNMsUtYxvwx6Neit3XwvWYytnBBbOGIFf4sDTMgVi
6l2uCFsxnysZIU6Ej/gzxxfUkwkqLrRBpWRyRwr/KyeKzivDp+u3boe0K0/7L+cbkJJn5b+d+XTR
vSSPaqd/W1CljBBojfjKOwaxnv8rMU6zWuu4XbvqY3/0Yd+SKFNg0ZCJvCpv1quttwUrwgC6XFXS
390PlqYc1JWmgwD1rRZECqOg2lwbUBm925fpec8qOWfIpFVoRRGiwb7gq1pIb1mMEW0pjgdBeWP9
RoKWbJQR9EKDtoNay/scRM/OmvllqIOM/9nEtFxFkLG61nHGXlijtuZ45RuvZaa9F9Ekf/EqFN/T
D7hkGNvE3U3g5kwZf7waUbBTgRyskfkCNHgLvtGgORpbs8IGgpupdf2kJ9JfX7oL6TTGSfps7rIV
qe4Ew3NEm82Q8wVuIYYKrk14UxStmyZK+ez8aTxVE3Wg8EGxJdO7QbmQL6UVDgm4BljXN/vsjXy6
fANh2YMN4TKFt42M9tS6mnudCAnK9Gk+iUdBnT8T+EkBCLKPfDAroQP0LK8qnA9DGUYlH8IwKUkP
S5C+S+4OoQFrDzjBxFFBylvgMrfdhOd8qMUe+YEt7RTOlWxQjviprPfb0uIO5wQtI+4fooaYw1+A
q6j8rRLizgRj0hOTkN8qTgx19K6w1faLefRuFcMM6AQEkYGUi2NrzKempXuPdRKMdKSsI7z++JUP
KNVLii5pyoVj4QiFKxMe7AthqTaBpDjTynJnFO3vCVEw73iNtelTwBSt1nWwfekR2DfSOIJlDSJg
9jYwFxNh9V6xvofyyvbNqXUFg061mSDELBB//PIp6zSIjGbkRSmKQ6E0gqhXgkW4dIzh33kq9m+E
Vhuy3GhMJfAhuxeMuznkXICPhudG42FRuqQzAmO8yuGCyzDoZgauw7Lo9BJiqg7fRpWrXX5WTGTg
QoBve74CjAmz3JzlU/5wfgr2/2yCnbzTHahTW0gUWoz7Hy1/wU3kzxly7Gwun5R7A65LQOD1Wefe
rwMy9B2JN+WSNSne7cFhNmj8ro6gh3+Xv0j2DIeGdpaC32rXUwCeX7XixFxySWKFUdp2Xc0VQ4lb
5reldTT6nvolmj46TJhZXgKqHyMMJnuaQhRfjR79nz2yYVRQ8eb9FCfVrJnFgF2zSZ5d0IltG+/H
rzA9NsxHxFAKsQLvyVRK5QTtnrE1yo0TiMnCawR+rDWJsOO2X2d6ZO19HVIjQ5KtMIBcHz9Un07T
3EPLtgBaujdfikZtP/DncbSECL1umJW7zrcvcf1puSxuPor4uy14ziOlbsfEg8Bnea6V8T2QV0/q
zUB4goQ8cfKIFcHUtMuf01IB9Dmja/6GlkB/6Ze2ta/wNbDDhFVCXNv8hvu2HJGemmeB7CPWn1px
bJ6qt810oWTliTCJIpZ02xKgyoOsM/s16+6n5ZuQxD0/TutkY+vTL32Jg8Vm/IwvoMUHcMTuKDqF
e0e44Txf58Dx8JxiSEirwLnlgc4ihbbuZTijFYKvHN+4c4iS/c65D9IQihrORkmmHthvH9ZskU4B
KYrpAknLxRR6IvVnhoeDjyeJa7ZQ5nvabldtkQzgdXqeMzJORCX+TJhqlXAfrOKsJjWVPdNShv5H
YENZOFhJUdyWL1+nar6foXbKqO/iB6z73cUz8ELk+nI9kgAvoQePQ6uCKjmi/z37Q0XCYTO3VdOj
3nYJpWTaKoPewGrsFH6BCFzSYC8ucfrVhKoamjYwFOV7iD+eK9DkER8nVFT8Jhu4RpY45paEjjyy
KVpgv9SZCVfMlBiu0265pCzEYkRn1J41Pw4RJTmR8aV7udB+8GXGzMRTZTkurXYfshdaogiMopdt
H9VrjafFjup+XdSW4yslsN8OrqQL4ceDMjqZvlpUftvN80eEb3FqbexIVb0it6SoQz7IYQt0xbcj
qhSRIVXESzvsxa0h9KiV3BNwydnXuc571pcqAhErtwsyhotHeZK9ljP32/+eCdcygz4X6MLsidSO
0tVT1qchWYYQZIQYPfOm8SwDwealVzKSolUBMI2ONvfHCCbBG1ALtKdaF+NukhsPoXYsMI13wfRh
77gWIaRF6XIKDyuwGrdtnSndjLa3RKPJUvUDfVz5dDmGYKg67L1xV3mljPmFC1po6p9jqwAGoi8v
Dh2gnetRezyisRnBKE7FsPsAXjSzqiQRadRrNLYvaZL4DSxkkk6bCKLavn7UO7W1+2cKYIBNXvLG
wXC4hXC42pp63rI/BORItadQfbE9igmYvF7nk4tz7ZupbdMqC07Tgv3W4dgPsEeFQyAHIPQruch8
MY6LDHK2C7RLbJiYCQrwXJ0kqHS1XQ6LpfJ++gfxC6l8bLDzRizLb7sZJIGwYmM+1XGwv69sBatv
FPTMJE35mgJzx1PCNrso3wmzyXCabZDs9g/GiGhi7fi0uwbND5knk59SyVXtY0ll2U2csv/gd2pW
rxnW9g2fdSnTJRkJaY83yK5qwQJmUm1QKWyJe4OfC8RCrp8T563mGg9VqTC/YGdl5DbuoRAo4sS1
QDIgf1hhy4tFkGXsNxbZgRQnVqZE/gUsrTUrfVRBeTxrVN5jHa4w9f0YCE4rAubQsMEvDzrhreLq
nwrgYCgRhHRkihx4Ywna8LahyeCgjgfKGKMnsIs2dweojJS6ymyUvJJPvcS+Ul+nXB/WfKScDxXn
ppFnfVfq5EwHXo/33KHK2274RlwXe6wqW7dYh2W2Y7t6tbnVybMYUl2jutMaRkOGAOCO60iS5SuH
NjCOcrGUqjM0H2znqnUZ9Kvm4AF76gakH1fv1qfxrC24aLwb0W1evYMaMwkzo3NGS60jfOz8ITa8
OwOKsrckBxs6pqbzgazDeRWrZsWmgF+NsAAv/w6UcZCJGR8TJ4Ec33wt2JZDuJFvlhY4Hu/jmvQb
h9agLaaTwyF3hm+VRty7pJxxOr7q/3Oq3YeOCSRqOEVD3ejlc8hQZD33Al45bONc1SrbAgxuLx2z
RdnAtakuKyWYF7wFDN748TJg/oqeUcsUAXGZGKn4KcSUX24Ri1E4P/LoZtT1s0evP0Y+V7eF8ofH
frUYc+FT84bbth3Sa65tSwnAIdAnnDvW/O66Ue9rIfh5T29y4pOkE9YKCK5UOPuYRHXLM3sy4SsX
CiXeWzJP7TDI3REANEq6GX+e4q62nfRKnLX5ykt+RkTacrQi2mnRoyU4fAf4774MKwp8dU6T7qXj
y4cCudlAajJcv6DP4hfDIyFL/iEiXDhY3m4l2F5g0RxYXUoTXXFXxJCEvvf5q2iGfu+JRwL1IJZ9
dZz/GBE9uJFPvgAlEgmkFxq0udZiBLbtGgNWAdTcXT6KPZ6NqFDXz7s8+LElTOlcKgXKXYmSij2/
me/qwMWmh33N81krnJSp0lkNoqWtg8HdcDyRNQ+jlKo9wx0w4seY6/aMN60lR3V0il4k3Y6B9fEw
dnuTWr0fR8LidXzedmdc39LyP/+2h2jJXdAQuq3j8i4gkTsmVythPVNDIRJFrDRHNQqvC7/WIq+f
vrEwvS0nwjmQiKGc/Skt/IUCEQGWEGxEhhcyeVvKBKq93Mxf/3F9qejgQYl/g7I6wB/peU7e/sIU
weddpGaUxYCr4z7KFgQcLTmUhmZDZmMa2OUq7+JlhzVWilzY4q5vnR9a2a18f/cTCD1aMyksvAZl
EzrPMFIyK5c7I4CcdLJrfoUc2rypczYwxo/jxWr6P2uQcn2s798FRsU8OHQtegV1URVQtF9J04OB
bd5OMzZuiBZjKOTxDLbOsvbjWl/Nl4v9N7D5igm71451JRAcwc0V3awIVXXfQ1fhk5MqHbyzWHrF
6EZZlIKGl09OI0WrIDbJ5ynwpYfPkmvBS/zeXsIOzSiCNPLnPG0Dp7hlcHPQuaIJ4xWb7eROLFFc
FL3QqSTzK/GYNsHfFFk57GOYumDY5jQYlcwtSTPZK3d2o+PfzyId0k4G/ZQD7LG8Uqi4/aywrUVN
w3npWTq9JFvszTHsbiF8A0mCph3P5I+YgDqU35U4jZHW0axc2apLHsn1FLuYB59TK9cZcXRIGLH5
9khBcxYyeYTNWnM5n2WIGV+5c7c9gIIM/74es9AQri5eJkEEaSLC1Uqh/2olhXSXqFC9V09sLAP3
cJKj5bt3v3WeFZE0Pu3m4eOuRn/R3YjQE0N4qKi670aWV2LHQdvC9KbSKPaSV7hDbZOgINbn7KCO
RvkG/Dk1fHHNdE86Qraun1zo0aLwXTTRmvGw74NggN0wrXhBlOrldc5CxqyVQZLmSVSbLy3TzXRj
ECkNrLuY0QlJUxY+dfJyEck+VqdohlHplmsoqCpdYFFmvzyeprOz+QcVTLUlqeC5pZiw+NF8PAxg
u/0upxo1PA36+tOkq+pNb2qyJ4nBwn+NpZsk2wpBAjhgze85AStJuUnuo7jztt8KlVpDsFwevOD/
jkJN2JDO9uH1ftzFfC6Wt8b5K5leqsSwYHxx5Z79gytbBMuPEIqcUJL8bDxSXXBTBYVg6DfBIvo6
8T8pPGkEF5yavae+O2+jefUJ7yo1RDex3RNQ/eGpMyVRHX6Gbzr71Fb/KWK0/NTnWNZnuVMB6xXX
1i+99uDbs0+0yfuQFLb6ftzbkI9UZ/OsTfrvpceEJmbOm2bNASCvnrhVXC+R1/BqVFiZFaO/+YU5
l2zfH4cgYFmDzs16hBvanFxxlfNihbUWZ7HExicpVvWJwZ5mg1Zd6g0iYiPAoOTSd0NR2ubPnFgq
585bHkajtXyVKoiuUQnWI3NkedMWplEaIcY8DDdrWhx22ey6e3/CpBXQH+GBwIukE80PXCv1v1Se
wptJpKWadedDHk02x2lw108IPtDI/7SnvuaEev+n5xMIERQFbcmERg3xAldBbTsRGTSfxICjVm8N
CVpH0Zmjn33BhQzZOKItE1QvRFPD9f4aZwKzDNK6qG2mUkIimS6VClA9Wla3a99FgfXmbE2N8WXY
+EqlQhMEOawRANY3Pr2LNmxUbgtqaK3sxZz4m54Io4MANTUzHZ+ZOB1tEU1M/7jlYxX0Gbfg3sB6
AHicDsS9sP/OU0gZmbPMg1wWbccUwCZs2K0mLnGX18nCjIaBt/A56jC9hzNJ3+TIcmlZmKXOhiws
4dL+C9TfbgdzL5H9PFl+dNk4m7myUOKeBgDjGLL+/3jirv/I62X8qGL6LyhaWPgPdY6C5dOeqt0h
Zo0OeE3TfpoOajfpr6nJVYB4Lr1EQTt1keRyyqs2juaH6708gRuQ0qL8GlMIkuhDVqsYfoeplS0t
o/Qbn2lWncAL0/b1/1C3m5lgyyBZqKwU8tQgtclSOed7sioqCV6NBiZNmeDYwnlRq56VB6oJbV2i
auC+6bwYRGuz8r5OUxwwTiETqqc4DR1WR66Uv/Q/b7Q9ROU6UAU/SKlS8e6dpoxLf/nwNJNKkbW7
hH7tUkqc2COBnNOS51y7by1O2kKs5mjIrsy7D6am4gGdlWUiBdOfptf4mZgx2g4OZPPiQoEGHzYy
sLpvkXs5q6DL2rpzMygCFg/L5ZS9oMjND1r/8gqr0czeVptyzSlzH5sLTGEyCtafHaF1r1p1Fs/A
1CCE1iUZwscURqJ3MXThKr01nyjEGfBJJGwqSri/pEY2djWDDR0GOEuxu3DCl88jAOuDl4OVc4YM
YjT2yJJlIMvEmHgWoKbazzL15yguTvnzUtRB2ukQdtHVBO8w5wkgel+UoycL5iqhkOHgR7BWoAVj
wtsbKLxDOlbaRMcCHwi9FNoukPBa2VF2hcEJjCMAi4VNYE9He9PSWOyPKFqqdAY+jlOZJV/A/JC8
2TqzzbI8FvSFc/Gc7iixDbJ/MTYKpQlFE3lj/glk0Y1Fa603y9brhKLC6//KtOzXZ+FdK1FybZ2r
PsH+Nu/nupU84cG8vl6AnK8y9h9KPqtTVhmK9cMTLyWPgmF5Cl70IoUQ8WQZhsSq5ttpjpsCY1bX
Et85sLE3ntR87v2Zdt3somYWQqky1QYbxOg7W7AZs5UeItcMZnsbLuO1WKto7n/dUVjVXyYYCSqL
QV6zQJHwAhPkiARW4aRorB8iKeqwbLBknEu7da1lPcmnu5kADW6VM5h5IwKVURaBhAcCCAXzP8FO
eMMUavqrUBWKrSBIayYujsCYb2PGMiQd0xzRLE7o3tMMp2E9sdJCRn9SZ5UUqJBSCAENfJTAwKSl
1LPDb8jtYIa7j9VMgvoOXx6Suz9CsYeQK6UL9vBopmEmoeG6sCKmI4mlx4stiuzmgRkKLKDwnfFl
l6SkmzkejnZ+GbxQVlO21HzKSnpeV4kpPBaLstHN5NVKxZlC4xCQt+JUISS6wk7Fd6ttl6G45njq
rrlUZIpFvwNmsoW0yPkPVOBQnNm6SeBTMsCRP1ojKE+J10KiOmcrYxDIkbewPd5/FAyu1EhJi2z7
FZpvJ6Fip5X0HB6NyyhcT7EHpNBtHpMMDf3EwGVtBzMbRa6KKqEnZet2sFRwqOwh3LLgE5CyhvEp
vX5mezUY5d5AQovTOzn+Gym5Oc4cToV7toQtx1QF3J1PMFZzFzcb4q7AuKooQcNPlGFkE+uPhs1+
G30q1RCw4CM0m5EQatC497mPnd20oxowRCkXMdoAFwTXI8bOBXgpUqlVGWfdlFNs7G0sGrGjR0F2
kPV9p3sBRQDiNd1aWn13btc3m6k6WXqmOuMNwsJf9YuZPITyAajbHkbO4ffjL8Ok7q8hPs/qb9wC
+cEkW10l8+BVg0e5/++6OPNMnyAIutm3QKYnm3oIviyuDqS4lv9zjCFoohRhMZV+9Z4o8yPBseZR
XWLk9q9H+A24LnX64Ewb+853ngiULdgZyzBy1IptGuXMc8hYB+MkUWO7zGn+CLWr70TcIe1DbRsJ
egVcZpqoIsjNd8UfJ+etKguyLB5ovFa7e1FdU+4YYL7xJjCaGJDYnZEmdOMubcdvTyJQvQyKJYhM
V1/MQ29zMPRqUEbuuJUKVn1WFBQn0SFodqREb8GXn9vMpVn2qU39OZoSXmGXKLPnjdyw4ES9ipJ8
CmmRPeN2lRhhQwJRDAE9ifoawKkj8a20mZOzdk4bUDWXwuEVJ1A19Izi3N2cABjO2hE0uwuz2afY
HDaYUM+wBaeoWMRbVO/8yuXDFhEGwcvWZ8ZTxxbjGSezdYRYXO5Tj9WyAGf/ouALUgA5jmWbsmEX
iJ79G1xGNutQTr03I0AcTxCY52UpBfaYgzfDovd1nn73MxbM7VupeRffHtl2S5bORea+1vTF57+r
Mhdss5K7g7lgzuRj795SOmy3qeGrfob8znDWG3gNkm4LZGcj5RB4wFwF6YmJ7Y2dZQzkdsKdc3/r
SU6DDgRHHYs8W1PBdd+KHnqd2L4FXs99InM2ibbkZkU55hZlH3VOfscvwCRNa/G/yWJ89vwVKx+R
44Gw2iQVFBO5jrXxnCIjG47BXDdOmsH9GjNNYWwmVgJFx8YKkg2kEcMNJ0eVLT7tdqQABi1YW4b2
t8SC8MLRol4nR2mq0DgG2NYG21UjzjJhy9ZjUjb5fOkDurMMEeeKltj2B/dXOTTdA8a+hyTv5yDS
1M7kTfOTAVrieNJt8WW6MrDI/tLnVUe3EOzOj4AQcLbwJSqiIBgDjTnpJ789hO6Z1n4pjeWvaSeO
2T9zN75tkeHA4mIBW3LyncY5rB02jkEOjNvzC8xguzm5M92UDyUJ8liTPclfbotUIo8ybj4RJX66
Iynu8FE0Z/Mb5FeE6lIb8KNjyn47tRZ7Xdq/2bHUxZDpN8cyBopb0PFslscXLnf7sav3cFh5SrTg
qEsP1VTjftLZlIzdNdpPlNj/4fZWPS7xWxLbWQp/yAkRIfbf3dop7dHiTCZn3W2JFK8kg7H4/9hZ
CFKtoLznf4joUA+IuDIJsRSC/spdYtbEfYBmIxt3R0Ko5o6l/OxPNUSrDSoOntZkUNz0ljfbKUbs
FYijE8EjiVhtp4GlWV3He83/dVxCosyg+YTg1jE+UEUCHu3FMzB29HyI8QlMJmi1wDSv0NvcymnY
alAtJSG5L1N2FPmNJPX09KLtY7rjmyh9+k+KTze9DJzU9Ujsb4K9BQM9aCrAwxB4I7TYyK9G5dxk
bfqFDMkYv8bjDk/RXf8onCikFHtWcq+vCsiexZiT+4278dtjyl6icXh26MDWeEhZ8m4DFPMWKf1F
CaeT9HS7hNPtsPGrr9XldlxyoYVXKHXQd/AlfdzxBPXWNJSE7xvyJXD5+0XIpmD1WomXrP5xuwnc
Ji0lpsseV0QkFrPEPim4mJgmHz8mvdMAu3d9ADmJJMgcNPVCg0uokbizjDLQy6Zhqc+i/hCuowTa
AYPWHKj9x7fCM4h+kAiMVU+scWouG4uLThT16ihXgNSlxrXoo9k7M5/njuRmG2xaBVhcafD1wK+w
1GBMCZOax9DFcmq7jxhXXBP1F13DCMkHU/iULkAeO6qpH5juH3l3toW05DUidQQQLB1+9U5uWbS5
602nHyDL/e6BKlML/DsZ234f6uIzg1051tJo8KJMLCUxiCEnuUyAa6tZmkP2kcgRkXgZH4hrCf/t
znZU2a2+JgfDVqBD6zum/r9GMs8bM+kGJ6ZJVnAATx6z7pHwnJknGMI4h3uVDxDlWp/Viv6Uv8L7
5Iv5RtQAzG9p5BO4pfOPZHgER9Ivnjzcde2V5vmKSJ/pVIbI9v2MGpZKWPv9Pw0x78bsU4N/lp0n
4rIIKfrT3ugYCZnTbOCbwcCyM3ClAmrmEYLDLwX9v2BgFCLIvsIvPN9t+qLxWNd+xYQSeO20xLAb
GDUJRnxw3ZPgzXVBxyumzrGvEIKm3Japrtuo/SyScIt8UES4j0ErTrYYd77B8Y7eyd27U22x3uKj
WbIv9A3KhAhPSSv9/ClkT//vW4LPn60oc9KQ5+CkqFa6NcgcdoucvlBV2lJs8z38CzJPn5XieO9S
2Vs0V21dwfUM2bqwyMwSag9/aFeoUZazs0cKeezqoJ13wviHdtRcGsKhifOPoj+8USHXAtV0MEyy
R8459Yw8D0HTeF8pUC8Z4u8PXbseC6fv4xOw30jj6YLdP5FsyIUbSWdFNihnbDn7G6koCRkP5IEN
Gy4Rkl0zSuSNNGsj97fNjjnnuQtM8qobXAM/oVxMFMQltwvfCK4Z7YjDY4me7smt17dUoco2r9pj
Kl/8AvXaJ7P88WNpS/aHnRPvQ6vSfxGeR7VKd2mVxD2/POeoceh9/rjDmTAmeOndU5ZcSS/ByMtu
PAZVfoS7r3fP3MCihi1rtkEW4zikoh++h9qGo9N/EW+3lr90JO1wC4pYa7owGH9NyBHDr7byWifK
uscciE6+Wd3nQAoBPWGlcxfvtU4P9SWNoY7IIKoIqIt79rH+awiSczACfkm3JgqBPY5+B+kqyz4O
H6HIFl8TRjszdVWHcO6EHvlneSRCpem023aZoOFziIB6ch0bBAXs0UfGweWp2fgLgFo4dSc0WfmO
ABhCmIJ8c7G6L5LIZbdiBXHjfT+98S6pd0uZPDwPiv7t8wiN4P9dvATUrH1PLVCZ3PHnJ6KIkKKI
EmHqFinTXs2ycMWBzv1TtMB3TM5CqazOZwxg5/9hSaSPe9eIV81ehHwOoiygwyNYIn0T1rrTik8A
++yi+YoyPmWuXVFXNnKigrTXhIlm7n35Dfu7KH+WgkttdfYDCSmTZz5Hzb6spjSkv+ExjrHYLurJ
MgTtE8gjWnbBJZVRGlrT2LRlv+1rrPUQB4RcwLb5AHaX64opyiX+sRY6blmLawgO/7CRisMT2uYT
NhHCLS1h/MbvFB09WJsu47qYu5p4opB08O/sbRKT7N0cNRSTrltpNoKF4uflrBPY6+M2jok+dz8s
GVksXVwk5+TX77knB7sdX+rHJaA/m9FRVbvTY67Ay1kstw9mHKIvGUM6LVFGVV61eqCrxXFye4Yf
MF5L7tjuDiTcrMnk7Y7RZnaYOmzo4QZVmKdJqCdMgV81IMA/FsW+JU8i6MWOkX99j935+EdmiULX
HCeToSa8rb6BYCvpHlSVCMuCoKZeVSXDmpAxIGLutIJBplTfRA55qxPwRcUZ0b8p8/HlD6TWoqT8
FtQRzDPtBk7xuifuy0GpH0IobvN5Htv8qUUP6vB4tdnwOH5wk3MeSk77FGvheK1dfOrPi4rnKY5P
8V5A+bgl4N2RQo1c0xmq9/WFMrCL5VVqebT/Pc7cE3+lccvc8XRia+aLSitEgElE/eXgou3iGxNV
aUdHeFLyFyNPZAPyVqzZbQX9+5kjc2hDLPtfK35vxYj9Qssq0n9dY833WWYkwgvO0mEtsyjKdv+u
OshBRhHLHJ3Uyd2eiGlvSELB87H7D/736FvDs5BnBLG8OUEy2ehkaJuX/y8HES1ZGJznhWPPzWmp
vKJdyNVG/j66EOP1fluMG6G5plcYv4f0e4cvGNpMmj38WMoK45MaQzLvCBAEPlLuA7HZCcCjcdBe
Zq1Ch9gXSOw06lvpKCOOFCuRD77GBmzTVX5X/rTUNgS5k/KQMDqYyLWL0C5Q/D7MLOyh+HEfH1sa
yIaz1Qaphd5Jqd6ldJYAkIIlLmjzdb+//uBKXvUs9k1gyN9oW11ar2C+c8uGc9xj9bcSGe5ZTu1T
7+VPDL29tp4Ak3HNCEyubNrdFyJvdkz6nOeU9JCp+2PzIelAuqp1OB86JBHWBizBoI1erkZ0TMgq
dLHi7G+Eetcpxesma7aDhuRtJdAoezRdmIdiDfvgF9N500EfGeDh2MPPHB1vkyF+zggCii9Y2VW3
allEk/f6U2ZBe/DYSruW5Wut3VunumegbS9E71CW6xzYhwrPrmaH4pOmZe7mJM+aeaGCxwXyW2gB
BZUhJS+db/PRwkbkKvP7692ZN3SfwZ6xenfXoyqkGnmguVqdn1ISLRhVmnlAzgxKRDCCBjDH4WHN
2ZS60cYt4Bp71b8pRVX1++sUnoY4PoZwKkX9TCUpYrDoh9Pj6Mgq7xg7AZlbNOexbe8AXSCcXfzi
KGyV+ElMrfiRMlIYWB+4e7SQcSc08Ts+AVkPmb0GYoMSxybOEzRETsCjTqUlUah8yf91mEUnrIeN
4m20JXsLvNRNSY2SLlk1UgwShCR8gE8WOkmTuR22vJb8rpQ52oqC4HJ+hDBMPOWIXzW5pXo7iILU
1d9Em0fxJM1yrLRHfwqj0kzS+UlQKu0+miVP+tOpFXoZJLpEKwhvrtpN7uE4yGYo+qQneAbKjgMn
m3ShQGdRdqUIF6xPkT9eX77FBdzirdBh75XAU6beIub2mXXWZBRREwKhynOkkT/jwcy37m7w7e8m
T/y/ohkbAunGSl52Odv9f33pZZFq5bc2+WoX4zrPNGgmM4fXmdLLJ6ui+UiEXBx4idiELrlbdRH5
A5ybb8JwLVvI017PuNjg4RBT0TgLPRjAT40WoX57dyMJxG+Chz6nLVq9677p5LpdSAlwpvgP9zIm
lyMZNNPFy3ge7nXwlTghvLdP3WLbnTSsB187sIiIrwK+gcC+eyOaxJR05L0he/M9aNHAjtoINtQ8
LGntlJTk/GFvEUE2SA15qTBizajLdDAqWX/Kfx0VtPeGrP88eKN0a9U4h6zSnIMoA9chJRaQNtZA
jXTRwgEYDj5J2/cACySa2mQ0qGddHoeVCV7f9J4SJ+8xuaq89bl0TP8hhDeKkrUAe962IwBmGBZB
3gLj4wYIcNTOeJrpzIMil3QfPjlTuS6yfltUPj6LiXjks7+Z6Qsv81bS8hdaP41omcp+tCuZ9d3a
cLyyjGnQ9j7jSRrHOhawlZa5Iznk/t7Ep2P/s/d+qq39aByBO4Z/Z4gSNQ1P0qY2SJbvw+bPbC4f
6tgm3dVi0OcwPacuwhsGgNcDEqhfXqpnXagESyLMr4xZ3vqTiveTaVoD8bJuRLPbJkV15gbaGZwp
6ylRHRKtRIGV9Ma+XyTrPZc4K8KjNtK00dieTNA4mTKjrECMp57hRVcMpIzeLkIC49iF3jHVfrUd
PSeRKESUGxrFR20kvE0PYekFTudIAhjhsRXkMIbkKvIdwXyLxuBAW3YTeRHCfd1UMzir9DtvNfZ+
LhxJZflrYMRGUK3ohQDaasFh2j1UQR0AawpOnkfePZPWDxOjdY4JS/3nFvQdIoqq6RrdjJqW2ALn
lgvKCCL2bKo2hzeKiOvj1hAxcFfdm3hdv7XqQwB3TY1Qh/Um8yoF2oXuhG8NgTe50JXkRi1yXvzj
PKCrPJmpA8mJjRMTqQoerQseeOFtbAImdQzLYY15qUw/J0lq9fTvgy/y3BR1A5EirRm0wMOHAlBA
6uTaYqv56cYHs1kjK8mvV5xqVT9mb4mCCHD+hSD9cb6mgIG+DIfnhyIA7WaMpDKCPDUqZ3H48l3S
Rb7CeqauTmwRDbnk5gVXD8d7hy9Q97Pv6Pjtn2MZfPlFt4dhwM8ySqZaC7R+RRE1vuXe6W8HjgD0
bcizSMaUL1iJYzbuBGO7lzB0FEybB3pxvTRI0cHwIItZeyOgXAcIdlzhoFiUiGqoRgpg09tSGHmu
iHFw5tykM1LD3LExuZ44Mu8E4bcx2YQNnAx/qYru7FicD4NXyVKovo+u92dOERdUXNNRagi7QA59
XNe2njK2wRiPTWntVMvmw5nZFdTHUaCAMwCH1rp4X7m8Z+8hr6hUc5/edfdMYYIR6Ut12Wfe2JfN
BrLMbwqQgbpDJanSz1uOl85zoQGdRLVUYf9eZbNbqXwJLQDltId928g5n6FfDp2n4KYCj88cNeer
HQdHimBOqI+ivN7VsHXd1Udnkv4vJvbeBxx5y4jGdrn2tisSkU7Bu585+GlGGeaKEWJJWFRILH8/
9Rmn0Z16jzJo8JHaLll60C49KwCKt2Qu7HYI0rOh3RNRb9gxdzNROmZFAzCRhedV+hEw5uDM/Z6c
TMCBSNaAlPgvUyxRin38TZr2r/hquLR3zwws4HEIJ8hBINVSpnJE1WdHhCqnd+2sMadOGPIkAmIS
sqNMH8EBBQefUsRZ/kGyQc3M2gxK2gTjEtAE32D/Zz2+8zgIV98XY9E5AajFJV656fFP9/VpzLmS
G/Er3VymhS+C1FH3fvVoJx61O8IgH553x3N8n6C7FQ9JnV6B0iANHgozCtNeaGF/80RzBasEN1l8
088OUGsxhyayoCgtwnlo2whwkBv7O4HwljIh8eo1B/siUj3V0yfFjvr2SpJUV5VzJ4IVLCQuB3wj
KK4dfhG8miPkefTvel7RQzalIGyyr2SLvFqVjOSiZbzOvHc+xzQCyPkClaCcxguqK/FDipXC/JXp
HIStvGBwZaEWSUjm8qipBbGuafysTJu5lrQYBJrizORw4UnCmkHJarsWgmKOTAo0Gs7mEe+BuFC4
c0eOwnvjYKS/UBu7LYMoBkbCwhXN0nfhY+zFsQgst6JQ02S93G1s/tHMjJBdurJmksqQT/ntOQOb
UbaaP87uSfX4elZSQO6FxgnxbEBksf6amhJZnQgt+muwcRC81AcpcZ3rQgoZqmlJH4iIrRQtw0gh
C/QCa95gEM1Grl3O0cNQmKslggb3b8ve48wgU1/vRm7y/cP2XomC3KZAdpnGWi+Q7WxI/Ho9CzH3
WXO0TAcMWrOGqTqc67cQj9eieTvIwudntZecF1QRuS5bhqyMrstj1KEbvz8sxbUpSPI0HFzvkMEx
JU0jwb4EUrW0K1/Y9/oghVWWkxGPQvUu2Gw7fM/bpD+Z0e/gllu++qYKhrNAmYCSND/TodfnXPha
Z/5FcnVkcQq/oDdjB70DSga0PWvImEENzT8eOlmWCfo/nN5/WIvmmvadANwjlc81/DRcfuyww3Wz
kkLF/dk7L7Th2BDn+Mm+JlG6+FX3tGmedG2/GBeqNblJVxp37bIkUy0y+90JYMOaPXYX3/2eO/Wd
jg+uyhO3l2ArcSRQjmYuEHMcZQfH0ge4tWMjwXlLkzF8ATCaOxh7O9i50zdjAzfY24znLFebDOug
7QSbDtoeIVzOGqATfljH9LUQZZW/lO1Ze4Cennu8HUx8jeRG0WWJRM44+GcfDvdmwCybVSg7rJcZ
zBeg7B9Y3ITMZxnDxod8GgumllCaTfPBaobdEAoE1gTaiBPUf3z9ZSRnmVBEsfJviJaqPUc3PmUA
QNIMqntSUl+hvZIbjXxrzA6EhSe0SzZUyeR3aHFNgUCv4MHuMpxPbA71LFmuboPbbCQMtZ7xJ+ye
uAXr0igaZEG1msEWRCrmkJbWtA8/6UqxBxclrCrnrvFKQbCN/I8Wp2qYDStednp7CChxhzqYvnSj
KaLVsy2Lvo6bTim5VhthrZ9V06X59+RdVc63vL3sCViELjy4qZElZLqgzaJRSMGov5IlQ2SPprlW
7aMtoLUjE6hiSLmZsWfXa8NcE4JYb1uchyOQZNjauDMmxpHPAogGY8SZDqV51oatqEBGyMyeaiXh
QEd/7zQJRo0Ept5hygBviYWoSmXOBKaotj7iYlD0Q0byjdyzZEmufPh9Jzq/9BIRPSM6j7Ydb7Bs
kV4smPNS/TWTAzDGueDi8cG+9jvmKrEsm9j9KtG/2+9QKDhfy8bCBcZOEp6CS/kws2pz8mTjeuYp
LBN7WUDzli3DV4kYdD2JFGrDgdQW/5Vp6KRIvufds0wN+bi/nqDIzO0w81PWQXMbO1DSdb4VW6rf
0DPcRDJvsqz1Q/BnEuPK6e059L8apVXX9IAp7RHeY5BHTM0w5XnQFtLLYLoMytvE7mjkAA22VGQc
PBd07qHv0DQgp6b2w+dD6KKVwCDvkCqAucrwXnfchn3l9ErwGFOqH9RRvBuTaLUVOPxX2eibz9/y
f1bOHlhyTt+ycM54R45c4kNott+Z0BAGYvXApTnawmfWgDw90Nxjq1EYLHH1GC9Mn5KetkLt2Kse
ciic30A658XoKEF5bNb/Kro3I6pygnkb92Zu29YXz4ATRcF5V11IF17exZpcRpHXCTsNHA5R+pBa
FLBB3aKmrFreZL05roOp8pbTL3Dle7e8cwVoYi4UBnvUp1g450a2hc0I3vvgh1tU/3sU19JTIyuT
NKKjEykm8c8+4IKyr5lkjxvFtB8zTbNUlwuKHnpDmt23LseIxflSRvNeIoN3daEC3Bf++E9Yz7OI
P5vdJX98I8X86PLV90h1VAqrMuJjFNqOX/jftikuWYfmOBXbIFwnjxvknhL3MoBP3xNko/bkRMzV
1yDFz/4Mptu5gwQEX+q0dQ7vRrMlP/l26BbYLyLuPkP6KoWTKmqM3c2Z6bW/6Q8+sPdHdHVR7GRh
ZdvT6oLIxe6YgP3KWBKGPhJ1vIezuVnfpAQ8zCSuhOr06I3KHP1DGbLXdZZ1HqYexp05iicYYItW
C297MXpWQ4h9t10W0YRYu4bGeIcpbbgP+F3nh/flVk6RxJs39YpPbEYdchQ1uIa6vYTcRmzO95Uu
13VZZzCRdN8Kol/iTpATMjCSt57ajmJzkZLFaD4RMqxwnoQAaCvTFrgVXn1CPdj3AVE2Wh0kzbgh
ODVdfVMpUvg51r3PkvjlVlUquWTT5JcMtIu/+Y8WEI1bNplypAfbHQVrwwRNbqo5Ujqty9GKvkVI
rfFPH2sG00gKv2eudFaa7HzEToASA/NopkN1sp9dEmjIncxAcZEvgpELhwuvArX/PiKFKJQj0I0P
nT3jWqZ1/zQJO4+IFiBM1OPXDsB4UnXTCPbkpI8d0KeQDC4Y+QzpbZ/3Bc/GvuLOj4qhyP8nQ9Lz
OaVTucVeVefYigJnHqJczE1Afkkur5a6cwuXhX0jZzhQm2Nd83LjrNGU38NYLgGK1H5dghKO2m0R
h9LTtXCXxyWuM+ZmrYaa01AYf0Ul0fdxC/kOuTvw/IVpy1oOzOFb57sJXLegiXM+njWWncdpFmba
c6h1caogI/nsbIqTSKmqxgOfTBLkiBy/aXzfJkUyCmTVsxrZJ1bpt3qNvAIDNssNrZvqiFamHYkY
HDU5MjhygxNV+Xof8At9Jw0ZoPtx9KeXH+l0RYf3U3o7g9afTqmfy+nFp/CKkp/KnBIq06SN+DHt
jbItFuxFM3TW+A61L0H3vV+mRckjmE2EzA3YHtvF9O68ePfE6pekXm9IQpC81PvOzoyiHOOZ9u8k
1l+q/tsr52CfvYc533dz3hCyxpLI9NjyIY0ofEPg9/gJ8iMqe81hyvXlDCxMYb6W4y1txMGrBAYP
PcY+1xQF04H0wAdhi9pa9DlnRSdpJO6j4A24afNuwIJ5CUCDjcLCDGme52DiO6AxSmr1M+v1dXIb
3+x/QsS84Bafctw6evPJkJte+kzUV7JvbZqH7BM7s9JtXthVxiIBtHKVOmXZdMVZIwTKH84ZkNIy
JevF+Pw7qmcFgpNmnwV5SzAUHWszC54CfXuUaeE16t98L8NQrSQ5unNKjoMnd3LOz/2J1vLvLGYb
swx34YonPwYd5uFwO31HQQcKgLhKKzTLuUL8FXxw9oi71UFlGrPti0lkLnAS5ZYefCZ1EH1frH6d
XWCAXnF831Oyl4tYuKd8KQw+jtEq0XmastSBM5LWb1tjmPmqumqBj9h37PIrkTtPGTjC27tO1kT4
azzL7XfCQPj5yqiD6On2W5q4jxJ2WeHJjOgDHdHbHoxQ88ZJ3Sv53TGdOSpC0ijico1JI8jeUwwE
ec1Bol6/QNwXLWECgOFxvqTiiCBKHA9+5zSI2CQvuMWdzxFSBey2X1vLh/iL1kaqxAEQGVtu2+pV
q6yjNXT9mS5UFmCeDXZSHLACZz9q6WsrvwVe2wwRVhdV7jwFAkbZbkAwgpAFDRiVItP1nwoZ5kAE
qad3pFQA1YB1rafqxubi2D2x59OCWPjgZQITjtfZk/csHvH4JAKn4hYSsL8aqCNoiUjz1f87jM7Y
G1VKhJD2CzqjeHjrgEpjtPud6l/MGopHVZur0IUNmdDEBrYBvk14ml6/qz+H1CjkaXm/bHSLMshc
6CKqFpUCsGhSzIIf85WL2mQSjcIW8IypNPKAnJhQ33JRpZE9ujEAO587oAt7tCQ6KDX8H0qWJl//
Xnsjc2GJh6PNJqtpOEiD4U4EGGk9QMR3+RfW15COcTlrshBlbLI+NbU/iUNwjpaStEZmpm9h8Rv4
WoDBU+Ynj7gZ0+a3r7HIH24KNfWnbNMNY60rqGKlVJE9TXsZX/0uXt0DKAc0sllj9RJmq9lvqWhX
gv6+pGhNPpDQQKrrXdtd12TjxDAUm6E90iHX1QPHL3rtIGsyWcOp7imTBQ+4agjK89mfl23rrsow
BpHU3SfR6gl1cX8xvgAQokT1es/jkSwBhRKZ+rRi1jhv4+NaObqWaC0kIvgOyT7JrLzxsGv0oa4G
FLZ6TxQJoBiL6HrXclhOsgRxJBl5h3eS/DPq9Pcoxf/vYhCCTCrhczIhON1RbfU9klIk/kv3Sd8o
qxdJN1467bCiPcblEKJmUY8WXMK+n6CrsKKNBcg3g9riNCLH9QjuQL9326YeMmHs5XEzKWpd1Dra
dvcF3C+BbccYHFrwby2lHeGfnWcyeTir7tnHws6LfL4iMpuFRVAYZ6NNrmZVXKuolN0+++gzQ8Yh
ZRLltQWObFay7Wixj39BTypA6oRvYJeY/JaWKJ2J/ZMeS4f8ip8anTeCDKo3HAyQlVRikalD2IQR
IXHoBcNaQ8mLZb+pIsJgGZbJU3S01Hvrn43AWMi/1l+vqso3rN5TpYeBExSwX3kGnbnAZ+PxckWc
/Ap/VKQauL3y7q3jbsmPRIDL55Vp3rhN9PkxJVCX1gYiNAMVa6+Bf9AJNGsW7RbI6YYmlVUsfuHO
XmVRD4IhgDLd7+/Nifyf8ks0qar4qEc50wGL6Scqv+XCC1RZOLzv6cyN7gHQFLAC5dSMrtRcphTR
evUirkwropK1YW0iZyfB/ijBP28SZWPVIU58p2CGNnsovmsbN6ONmZLqvLLUTPAYHMDMP7d0c5Px
VAnW2MRB8ILq3QCLHKVcc84WS2/0nTnr3+9pqkh6v8Cl1Hj/dyh57LMLvfkCSFi/zencgGyYQ97w
/D0HdqS/SwcihgLdL26nfGtn1k8+Vmh+hQpm/ZE8rY7/3mFLUUQ1l/FKvyaVW/eFmlX4AV+1pRNG
1srQTcps1iiGFMFctKtsyLC/3JHeedag7K2XywdqqdtW103BXCmF8q/HazFsutAGBViltxYy4THy
5WBLNo+eBULajPKKt1i7+vc9jxuN2oNSD8j/P5MIj4b6mJpeYV1ptqc7CN/CNQtgR4Plc6el467N
yEAxlGX3jbr3FFDH4U04U8fL5/8UqKxcXR0ox4Q/Dr0OctWnA+9M2kG1gIFTxt5lgdmCX8KT/+cR
+IsOuVK+6Bx2sRm2ZO0t2IytD6Nu6hOZRn7y0vQ/9UUPJgoPOjTDxAPETAGrAA8qRMqmULB0tteX
nEJ7On33HpiBR1f1rYHcaV89zI0j/eqcRhg6sWNMgm6Zncl7kIBRuQiYttW7snfzNNsj89BqWswe
wU5rAZZz3olKtqjLHNx0gBL4w3rhGpJZnYOKowmeiSPAQL/V2/CK42NYEsE1Ms9qFhaykVLLPEVR
GVbcl9wAJ2ScWt14rrthid3d9WGPK0ayZ+NKTgDiRPTu+C9JzdmQsGpN1NSrAw/Tifoqw8vC54ge
B4E/giCNVzqZuec91EVEYQw/X6PVPTRFSqERpbmcTuLWDbRfMU7NRNCWeqThycwUyS4T+M9s1+2F
QjPb5asiZYXZm5xEuj9E7LJQBDeDFwJEjpkwQwHjyb79orPv48EmVK98OlQ2o96xC8w5xkjz25Qh
MFKsAemLSrgqoJyWr6jLEDP5GPZb4VSaOJxVJT9sxDLBvuUdL5mg/Gvh7zcHRvottKd7uFQ5xWlV
dDe/V1ULt3Peb/2pryMadMZOpojQ++qIILu7mPk4MZJ6qIzRKfluX//m7HC1PaRt+cXJKaTX2LRH
6inR8CtaYFyPJtzGY53DCW4Irder2OXu6yVUax+Gq8K6o2tG+DHYIp6atYRk8h08DwpMeWODe2lW
jEtLnfnokihynoehKyGxmtngIryFy/WVtFnFuqaXL28a93K8FPuscAKVgClWWze1Z474qc7CKxiV
v8aFy290xOOOjS5z0KSFpeXcVADMfAi9yL5YYBHOzdW5G5skQLtQH/8G8IohGt3eyeGFDu7Jdk20
mB0i3Jqjgl3DIpYypUJpjG0T6WfeiyGens0GwBTmd59ygZmdWSDpZOxSNfLtxOtQnCcgjCUq4NHr
K3w0k5VP8XkN18h+S4Jes5vAVaAFgSm5DM9q06ljJmzC8s8ixIXPT/7mpaXw0yrR2os60gtoML1y
wIG1cZedvlLw0C8JFzbdRfnB2tuP3cTr9NxSfhxskBUAjCBZ0gQqAYKRWeikqnyWxqZGOHi36aar
AopUwp1GZDCEveYlFSER1PnypBEl8vWD8SApZzdUpem5tEkvd0Te9GOwUchKX03fF4+wYnbzmWhX
AQWuBOf5XuhdiOsUVY2YlRTPd+WJOuOwaGxPi/WElDKL7ZmzcSeo9B8zEX0Tbh1aJhk8SWCxNzFr
S9KEqJrit9a491ulxltOkTaiATh/JDkskabv990rYyUOeHGRXNUKwA0VTGAz9gw79z8UFwSmw0cZ
JwRyOtLPcjgPgVf8ZG440wPOPENXnePEWv5uBcObEnzENCFEGATNByQCy/ouvM3yRbAeq3T2/Q5P
f1wh6QBhft01r0HjOscXd21QsvOU6czPTf9QUV+o7m6nILvRv1vY2s+eNSJ2oyD9kB1MEI62unbK
p/NpnhsNyCrelLCiwDWS9ZhI3wD8JzOMAmUxnPGPZt8/vcheWKuV01OgFI1ZUwKtKITGkdbXMULB
il7urLqADe2fstpCqudftYRKMEhftoeiCeqBzryqdpfguHxG/gFCSNgxrevPZl3tP/hXdWWRavLs
eT1tpNnZ2C0QCpZaPNTVjFKje/SVrq19ZFriRUuRwzkH9Fkp9To0a3vF2/rXwEfvdDnbfCfMZfzJ
BqOsPbqRxtASz4YMlxHn/G8HVYjdK2atmBgQS88aIwwT+KbKcx46nXv9B7LycxB1eA9j6ZgNmjJ9
MvPzra+Qh6UA/76UdV1xo3c5bvaAcMcX2TQdq7xz5KTZGouEgjxldfeAMquu3VXJf5b1OrjVamgL
7QBDHjVh4WwR/xM/Kh/OBqcLL6gYPWjaKzXaoAkAcjCI7GjADtiwg6LfBKjye6W1Z/bq/QCGGhT9
V/8DYg/FtzNKglSuQGl1Jugb38qhOjefMCH0BcfKzzBWA9/Zyuo3GPYP/UPyzNW9lb+6N1d6ZODv
DKTYZUSXsQzV3+7KXrTnqZWSyzDHgkcXtbfaaA1IsiVvejkmeGv4r/TEa/Yk4gz5tiW26IHU8jPj
x3NT3/Q+wv/9G7ej+LuSB1VVK1KFyN05eOk7aViVpO1rcIbdZ/IYbZNs0F9Cx1ni3g6jKzcGtVyM
HjTjVtZG1gESiBq2aHotarQKMxoCCevZwr+wV5tn1NgwZdDHo3sNPgY/uTKXQSlEzZp0Gp82i1RD
l5fulV0WJaX3jfgrDJilRhjP7mWhA+yWZyZshG51g6ZFcfHpuA0t2E7B4tCD/BQPVhSooLR+6s08
FMw1naBd5pnGhT8LZxzqXZC1VMXbHeE/i5sZ/IUCeFo3zWBIoPSqL4zqPim/8W1YGblNRq8VQspo
9fba0RN5e2c43uPDV+zvJ2MZsPTExMMfkGR13XnIkSIX+nNqHbCQGAOa8HDsTdoOeMyYMnMPKX1G
LMQDrvHXf1rgiLYaVhuxSPNblIG1y0QYJoqksbJ1DMDVPvjzdV+UuwLp1ay3/bsWN5PMP70irgMi
WXdm6fC0Euh/oM+BV6JWu74+fTA6xkvQrM+BNDOjP+VyT27xNMD1chXhccRy2bIWVNqCj3vvL7MP
Q805HSDOSda6Ps4j+UEgbXAWmqkSHdZjpAXPOw+q9USekxf5GbTqzOHlpZTSYolNTnNieZ9IjCHU
yiQCgZHLKIe3pvU5VQSMQ5fthG6ENN/pp4k536Y4NneLBY80881c4EizGtLwxKN+FgYE7MYwEnuJ
9gr3qKiejHqlQsfn8BEi54y7Q0EJDucy8bgGV5Lbv1sH+0q+gyfbmhhzyJpmcHj2Os3SFtk6KXh/
wLyNimk2gwWsTS7IBhFsB4+1Idl7ptoPKkeofDXH0RNflH3+sFzeHvWkiF9+1C3YQGWMkiqC1eTq
BtxSpiGeLwf7PRNDXKNc7Rff3nsxdgPrXi91Idoyuk7r9VQWjz19sHBWUMROMCE6bXQzggo4L9z4
GieXngKjjZ9sTjQia069VUSxxmWC9ftyJ8O9tk+HlnkIUsbslhm0rX0E7+LI9+pzFQFjhrGWcezZ
+YLlRSP0Vnjxz9g+Iv6d5dsLP7ya3NRYwv5RRKwL2QnMYbN4LXgpinknivm+CmQqlakvaPMRa3Ls
5id8XvTVRDC6LxEGR6qJaqMw5+VNi1/HeRrGWIujo2Wnl0GXqmufWaGutUGLQTV3ogICBWWLh0VB
xHRNacmMMepLwe6xCPWi9Yo6JYDO9C7HCx+GpJCE4dCduFiEvEe3MGyvWdBW6R+z4217UI3YCrT/
6F7q7hb9MI+mGhUV2Rcjl/aTWfatjooto7KopVEfh442rRS820Wm+n3trGXDRytIBFeJBzvHGYrq
G5Lsq+ZpKATeSRwOGOxZkT4R/t/3kii3xQgiCoGcH0C/Ju2uDQlWASg/vP4TsxVdMn/jopKUoaPi
69dX4rq2HoexaNxw271HFhsT0gyYo6y7JZgGsGXY8+/3fIaDqn/xexz8df1ZOvuPXXRqEjaxk5OG
9AkXSm/lLVsppG9D41iNpQOzkbdqY25d7YqRmsTrBMPyPilxjGKUihnqmuZ4BIrx67BaOrjpO/wa
rht+T3W64o6c7Mpf1Yvg+HGclQFIrFs68Rc4gfL4ySdXsLf7V4n8m30moWJFQObsLvataIKuVVT5
pdZkAtPD00rEH8/OBTbXzpmBuUC9+7SIu0LJUrfY/AtdRVyqrkWeBi1TNB6h4XcV5RipCo0w4mi6
K1P6Y3mH8vj6sWnlHx8wQb6WPFnDLxuAFsaPCtAeZeQ/Hu3WuIlM2KFhi9qS8P121knP4qHITcdZ
H9DWyoWDrTrP5Dw1KqfTitdDWBR68DpqTZ4dGxT+9MNyOZvunWZS7cJzwT/95HnE4jcy/SoX/C21
O5Zjd51XxKhCEtqdtUhhgDiDnJGfyXr2jrDVuEqvqcLpqIaGMNFcBARV2HioU5e10exCXbizfLIp
2BILMGM+KC5UtSYc3hHZgvUkoQgnmf/QqkYLfWspcKs7Q4ozpEGIbnNWzWS037mISHokOcs4vndx
VjSryFdJe96zSuBdA7CvX+4VoG4zm0WGOnlX4eQh/sFEodALDfoOEijwtKYj0bWwqJbxaoHp4XJ5
xg1nzLhONXCOkHheCtts3NCfWGLEP6yTumnnOVwnEzxfz7gJInZmPZJZl8o+gEF5X2xTgwCv3H8N
ZOtXiPZumc+NNMoNndIt3nJQVOmVV2dbRn5SPxYxrJuzgv7/6l6/lfL0C7DJ/XyEQt4c7MujRoAx
dKQU/BwZ6oH402BJd2MzkSfWDLNng5pFsBlpgkvmkwh502ZR6nJhWOYIjmCYrGdvYCg5qHGw22vK
U5OUZyv2j24CZbzCvR3zxyjVl75Hbxwnxv/cLQg22v3PwHG/c71ySriTZqd4pPkk2glzs1s4VFJY
8XeOxFhH0g5amhivmXqfWvL1WMHM0a/koXvRbqVDNRR9ZNE9tETscXzBxymzKQUV0VXGvquIstXy
ZDe6ckCbdUfRJPjW1u2q2iu3M1DFOvAxBjbtFKyyHNfKEJ0I2/sG4iR4s5kKVeZZ0FMSYcwxGOD/
XXi6MPXeLx5dpvbkCWTY3ytwXsShvlgR+f1NpLdCw4QXS6et079ZO35ut2JGkisaABavxSLEaY0A
qy3RXgDS0vofs8TRQ54pW6PT50b/QJqkjObuSISou92NzdL7bbZpBsqwalvCdVpqqY2WUTHpX9Cm
pgSfMQnAuW0PM5zoc3aKLlTY0zUUcR/Q0xUbuUQu79T6lNw0RdoqlKn+CDpRWFDgwXSc3vyN1XIG
BfGC3+Km4lfwo0B0NKbZc2D5a/I+lqjiFHtbviTQEJ0AX2feJka+2gio8yevi0BwqvIXLHiajerw
Rp1Bv/sADxENddZb4VoF3eqaDmxz/KTbrUW0/b0BX+vRdde3vAglY0FpS8szTsIirkQ5SbPSGHND
Zm3rNNvBJ8hgBzIMUC0WZgaH/N40D01e23jQS5+Tf41StIzEjxJQUPiSI61xp8Nwa90ZsAa82SoQ
WCs0jmCDBqn4zAW6zK32JcOQRR1cGBaKQbWMcwVjGJnPRlt1C2BbbtrtIQL3PqrnemFnK3rprstG
1Y0Z1any5rWSAvQGTm0K2QXqTBbXlKSmHCp/9rdcfQ+7okS0BEQstpHORDamEPl8vrCbk9+ztG0J
87ERHLqjHvupT6K/z7jqiptMdCmm8FSfcWO/d9GUIEjWljmIfqeXKWBVfIaxJXSzWPLExc/RVlO2
Jt0oxTekbaOH39jA8ozdN5T1s3IuFbv1kcU3CbIMqCIe0He5ckUgo53fYsUw8zjIB5322hFDol4p
vTaOY3IBgkTyo7ol/pDZcymaz8zafnjX1GAcl2ihYW/ZOyZG4UbXMCEiUC/dzkRlS9JUQM69Lqnv
d3wE1aYzVZ8kCmMMyWBfn8LhmBbIo3absX22GU2CO2g9tw79igN6DY5dUN686Tbxkn43kwULnZEz
hHke4gMSpAbuz3kqnD8CmfBU3ZhWR/TaQn3Cb9YfvsZk9jDWLjcrUaM84GO0lOWUlMSyqmbec5Rg
L8SpE9K1TfYmbZ7SgnP43reOj64zVUi+LM4/EUyK1cDcmr1//gttCgCmXL5yPjy3711C6fPBb+xT
smssJB8TSqCSsyzBrU006ZqAKjE0HfseHo2UFdnuhu3fjTWIMxg2lkUsRSdIuxmFYTwTWuBBkR3H
1lwOxqhgjMvFbLi/1q437V5Kg3ej7cR+ZaLrjDFghyyiKiYJXHW1MMhKr59UGsr+EOVBBkCF6fEO
R1pVzUjuKb9uhfNaQk1DspzwFwcfXGKj/I1TrMlYslb5OsqjvQvpaf76nOxPbAZY8eDRPwImzejx
pT4UiAgfi55EererN1ONbMQgjOoKCYiSyTf+PXb8hLJtNLIQF3gnSTVf+h6c+faC+Uo4U8ReKkjC
BynTp2r3oMhJffiH9D2TZxKOv2GsvAwj/ephoA+UDiUrIDsCH281au9Ngj1eAS1ZO5ysOxLq/piN
tNrQRT6FGccFazNpnATx/zJpjnM0KkcgQLKE7oW5j1MDEs+o8pB46M3A2lwXS17Q3mkzCQ19+q9q
RHAToue2S6RJuw1l/Xdc9SUBtoL0wiNBvV0b8vp0aP6EkBZMA7kf+RrkRAZTNHnmzxdxWg7E4Quv
EDh7u6uc4BK6sCppYIGTjC2lV9gAgx+f73JqcvObpXG51ETH5WwZwusGxzZjRPhCJtq/88OuJfyA
POOPWmsrUXOZSpoU0puCTSNAghIah7GmFuCB725ABpHM78IkR8TmYBOKERorqu6PVgJyhjd7K9X7
8RUAFiFrOektv91LOUUYGdBBXiR7ArNCBa5I6wDrG/NNOXNuiUL5K1hdreFqmjhnkTcCFCTzQ6Mf
emd++9syW/UeKcY1dutjAYCLYACoLQXuZYOI+20x9+oz7/Oz7beoDiKhE6RXdSSTuj40SoXRQJET
jQQh9H7eSMPL3Ob6yam++8euz6zZBWWyySus13STMh8ZrtC9vbc869UHIv0VPHULx31oPvbXtShW
Tfmftben0wPoEp8iiJoi8ZpBmf1BffIv8YtRX0wnTc4cEahHycp1esZuqHMJ24UCnDAie60QIbWe
5Jpl3xZAXf0QhJwBXN0MKhcE/xYqhglvMjXLFgKOIRrOQ4E2hPrze3cSjY6OQ4rEtRFbEzkHIfYW
EcCLx8t+Tkuy50w0oroV+vze0epWpKhGkHhQV0NOwf5eRwFTwggrUsdzZimIu5U5xC0bB0MsYuMl
b4SNOaAFKPw9gmonDqih63aBCTMTAPshzwqs1nmKkVe65UdIYZuSn9pvRjL5NT7wWlYUPdRnVCiB
pB63n0+7yvKjmnl3PmRjuJ9veqqAcrlc4yvDinzQ+b3/ky6ibU0uhk2JJruBzm0VbQaKakCOEWb6
CjSgNbWNGs2hdBcU4sn3rmfk6nPQHPyhyqUfUdBPvFup9HxltaLyymg8TLzaHmkY/75qn0NFgm0V
yiTLRZSdYiaS5IQjMOsYzjAdH8WZOekRCTjgNS90IH0NcPAN4k9YM/qy02i5JISLggW6F5fkx3GN
jgOWW7iNvBAM79WK36wp1nVitfZMKQUdhZ2almXMnTKZUlZHre02V9uAJ8ZIfl43BnNxAfAzVQ4H
sDBJdaiJnAzLS9iR8nt68nHI87gfqX4QRvK+7d7tG20KwA1e5s0YqI0lxDq2D2sYG8z9QBXRjxyz
R9etvWBHUI7Zwvq2Vwatp0TYMtG25ejjt/SAhmG5PylUtr4m7BT3fhn0TWDAddSKWvMYoHLw1DPq
cxzraEbtUvdNN9fdJ00W70/2aacLWFKSjfkeLB9Qm8/CwOIGQWb5vwjIwrnaJXZBgrn9HxGmN0pg
IS9xRrgRLtG2BbVazyz+s+cIgcwvAESR7zJHv6GHwrBddFY/gG1GXv0TqXvRqiec9HTojHTTFaVP
H3eTrCxRNNHj4ZNH1OCJJnwygGjIAxYsldO2Zc5OkEPHgNt3B9oyfQ4o3I6lu/gupFoP/V97c+Dq
v1gh2shcyV+f0C4Ht+cZjoa5YivgkMIh+uS2ikm+kVmJNR5Wua0tw+jJvw6WsM8lSJnfaFUrQgho
frxYer14qY9V4/DJHR3J9JjFclsIrNG2Ja9SXM1qKxsnZnNG9BdV2tyMjBZnUMv5GM4pDcJQ/z7i
JpWzg+6D9pN73eP3AetoG8EXfz/oBAfzN41PiIw8cfF3BoozmTQBIXaRPvR8ioCMMlVIfrbKsy1U
3Nb7r8djcLugkquAAGqBr7U/v2DiHYsfS55wlXFzg3f3K84hu0jypHW5SlPaLoHWoLrVFkqvW9wY
xFyOlWOc42vXIUe/vxB7lEcDqGxbzXL191p7PaKR+IJkG9S1ODJjcAI5K6eI+dby0HBr4YS8txXY
Iu8nsIaFIfrLIQZdaWlfgpvblQABlvQDJ/G+dRo8wiY1Yla7QtmhtdMOjAEdGHjjBLHySgD15wx+
hVT/exKzZ3WVmVW9FbjhfmyqvRZbAtuaA6IjvkOp06Rv4vEt9fiZUNTBNTot/DqHWfaq0N2DG6RU
nURldrgouESnhnx06bb0hFKElDHgOQNAkcVOk62L0+Qe9O0KhClAhWOx9nX8553QVMC5ZWpoZCED
Fu6ZYNjVlomseqTBSOES9e4AN2Fn2QOMd8D8MvA0OxiWUx7Qe6+qZZGS1j+8Jj0VPG6N2GHMR26a
e8f7WalBPqyUPWGAoRbe7yqF+W1xfVASny7BvHg12STK1lz4nJajPnW7vsKCOiAGAorMcEPgRjce
mAEVef/joM8Z4l16pJ3pbDd25h5dKmo4LOTPRfvr1rRBa0dJUULcM8LoL1LRpgy40X6eJVsWdfJm
K7kpNa/VBp6W8q6efdDX0cod2oIik8cr3QSRiDyVU7I/AaUQwhf60LZ8zQM4AF2P8hMp6wzUR/XI
v5AJmnvjpPZLbfqesz4ePCEbdwvyQrYKa1EZdM2Fl4SY4pCJJnR0aB2OuAzhKEKn9qKDZwZGsJF0
/FIQYZ8nUfrLyZCcnyFQueP8DQryHZWV6y8CswW92WKuEMwgFd10d7bZDRGftEmCBFLh979AF1l8
wFRbbQOGbZkrOZTiaTn68GSVFkRLnkWjbwIkuqAwaWaJy32dn3tNgllzvWTSARX1UEgljyewlsA1
yyZR87OGC7pCNq8mw1PsdBrQAcZ/WtbwxspI72gJBqEjpZDfr4PN2iQFULsg1d6fo2YB90mqjHb5
Dw9i2Rl+L7mvUyIso/SOrYUujAnprs3E2PU/MJ6QngaznLJXSF4CQ45fSp2tdyQFFVNNilm3z4Z+
NpGYi2zQlDKbPVPWb4u2FYvlv/3LhpswIaHGCZDnV+ILtvodMevf+2E9g/pbgxSTF5ENF014LSoi
IwrOe/jS2xTWKm97zldCuVrvszHpcTjrpJQaKx2tTz9qjexkgSQGGQRFsvquEk9mtRI0prN9bfKo
+1l0i1jN+cwCz5YeP2oZsvIz+btMSvqwyC0SnhWwLsuE15xCDpDDBZxUDdoxa510tx1OGmG/AYFO
hwplal5fsR6F8f6PfDtI/p+lAOeUgX22v6XL+djKmjbkeesEeZ4eam8sap0L9qCXtJU7OM/GQUWw
usri15ofaTQSzNHqaKzce80ysi/VIo+JAK0ibCH11Mt05By6pZk+9ncoUoL7qXOBjnODzpEk09Fj
L02dlxW1iz2m2ZSVdshoJFUZ2LQRJsZu07+fYK+Cz0rMu0Sx7PvzaWUbUgzcKfoZGxGKG9d3GyX9
h7CGNS+y+421tcFweyttyhKMab0AMlTZVC/RhJs95jwles19LLXFBmigwNYuCR8DK06CbjP4eaWU
HKUd0wFYI8DUCqgLy9h2V9KOiofAQDkGmoVPWbbOcidOXL324o6MN5K7fvtLQOf+HKefM7dFZ4nC
Hp4sD7jNTSlib+onMIHFfvqvxGyGCNssk3RLSgXdBgtnyb5TjL9+CmW4+IYxNTrz0lB00+aFBG7B
8ET+7lMReiqciCRFWj1pJKYYCm8/dykb5goEUYUcgWjH78eBFckJLGw4AmOiWZr7QmQARoIihBZ5
lngqk1QJIip5Hi9qqd6moT5iuwWNCehM+b/4mMgwtwdTyJzDO9AvjSbeOq93sduAiuppk8qadxhv
fCW1laoLeICetZA5/WiyEw/r80sQGblZGt6JzlKv7H9xJuKBHkiqGHt66DpUTw1xv7G1cK05wIIe
J09FMV7RGyPAFKRqRDtWlUbc7XNpEU6AfJZffvJvj01LTnK15PVtjzJNJ60AdLOkA5Op8oTTJhqY
aUuk9CWf5kToKzsBINImu0JdLehduxziRmvtYAgK7yy1R5iJKdaog/vfjlbpORBetG+J2kAbK9f0
BYOETXI6REXiJw+GfXjITgAm+aMNIR/btZlaXPTZWSViKpUOyG4FEiw73KDKFajAuD3FMD27szKv
xOvS6WzMzvra0bn13zIFZlo0blRHXJAsEvGxgAp+ytE8vgHnKvh1qPNsWrfJsW0tIlk96u8WXMU+
h01jceQvSqO+c3zk/H36/RUAfpmWSXJCndTcR3Ybn57Idl1zaklNYnYc0gcyIEUo/mgkzWvDi/jC
1oTG+mB+PbiAwoMxSDhXCJ/Pc+KxkwjnxaxAHR4HPOn2NPNfcYmdgw1fDiQQTXOgJy/kFPfeHrfu
QQJoFardcaxED6Otmwy522SSeF/Hega5F4YQHXbfBiin4Rv6IAOLVD885uCMtdG+De0nyfj0eaBI
g9VXg7vg9gbWpvmgL9xaLdGteoePYNDTQ+PTq9pjDUutjlQoaL19IdQt+uSRI0lWXSRK7mzUt+CV
eYsbKxzczS2cN0HJhFAAvXmOFfMMNu7tY6pc/ypfRVzsE3be8hXdD27o0nbLMz+/tOwx6cwkG8pJ
0m96Ows8M9VzmP/V3b07f4TtuU3IGkaQMbm2t1CeE2Ef2YOhveVveeSRFTiPkiOWvH9dJ8usxMh1
VOfzKDSQz4FFCSjP+BdxPwKtitF1GKAlCgZyzYkMv7z3E8LSXEcGXEuaZDhy56b00CthoOCHowqf
CEHh5u2KNbZB9x1u3w5utKNDi0mBGT+ZeOF/xGV3PYQmeQEqD2qAX3QlnpwQbLT3Pxgdyc5YkfD2
Q+Jo08AEFKsp9Z9rPWkZ3oH4AWOWT3fkinYTxaqh1WPQQ0RwOY9OTMCfEn3lkM1DSyIzKXY5/cxP
hIpYxiCpUlH0xFiUc/0CayFTshd9RVPnv7UUPB1tFLqmmwQcGBMDmOXJcbexYBjhFdANWPYs/dSc
jtO8SOwTo4okIbFDmBRq/LNgpP9jE3zY/xFOss7jiVcWLbnH+v6a9zrSIX7kH0vYCkh/FZ25BVdf
cMFQmj/BTEcUeVnzvdlDRjdb61epxOeEdDlKFN5BkRFusi8YUPTsmX8CLY4yOdxhcafKCrQshB3Z
/5TCA6s4p/XYug/GXpokiu2uJQj+0mmQr5m01aPN2q0Jby8axWwdbqlNGTaHU6KBaJ/qN3uBWf6I
1YuUDAkoudixNOm3DEGg6iQBdB+Ngw9j4N5kDOyShscJ/J214SHBIP3XGV0sVwBm6N/DkKDoNlnJ
d0BrXHdaWO5wZcmWJYXmLy2Ds7djEpwoWNLRr9jPqKrV1MCLk2GQBNRyXEbALBy7b6MzYKUFRc93
gwywbvSJf1mr1F8Sp3ktN+kZ7NjXGQHjAn4TLifK9b1fmADn7CfuOFoKmP9qh4b+/aEpoERAzsNE
X60VxX2SHGVBD7HLkQ1LpobUa5QsADAWbfX+KFzaMqkVzLZEZcuz5K13/S3YknFP+9xeTdMONFVX
9+EFe9azXVmXFLQ6OqQw4wC9/Q41xGSpzwwdfSz1kaQIFIOVREM9Jp/irFIxAlC8Y81Lf2PloWr5
8TKGWJJEmxWp3zi8jjdX6FF5MDfiGKsLcX0oQx+AInNNGkmSOX1Q3DQXdfvcoccBN5EodhJ7W27u
8PRI/e8xaf2qTAhX3cqdQZktd6qknMOtOhY6H9FcMTcZdj6p2i2ojbL63HkiiY1s/6WofCZSsNbM
UXnofZ5V4AsZF4so2vVA/5zZf+Wvlt6+7Sy5iCapqBY3JbGLXptupq1FxCC0tAhppINl3gNtvMGR
idrRZblxvt3K6qC9wHIOvdnO5KzMvE6EiUfbt4VmJqxK7PIx2N45nU3ZUgPIm4a6Ek0/Y5e1FJ+a
P/DNl19aUcYqc0WLeq2vfrIxwfD2IF132ZgkyQ3/jDiaNHsfZszdl3Q2eOjshYoJa8SgxgxmGNV6
c0m+++rlWp8xx4cJXwUrwLFOvHdUHMcmV/x6I9MBSafKvYAEGZLuGK0OevqFtmAooyHctXT7t6XE
OHHKBCzn8DWfx4voso2SuG3XbFm4J1H54aMFMqYy8xaPo0VFavBDxUJGgW3clPrhR7YhrvkVvWZa
a1pTJaerGUhBe2Q9eYffsyar0v4nVlyO8++VDANLQtfV/+v7VEDwImJd19fEE3r5VuxEGYUizhVn
GhfnlCe2I8+dN2LzANd9ePif0dzB2bxHPmOZsAJKzVHmRShiO47ucTV5wfa9CQ7iTGcf9FwW1Lwj
XLYZWuyP7eu7IWaWj05Z2gf9QGuHm51APcGPWgw3iz59qV+qxLAZA3fdeW5nh8ZhLhywC9Bebc70
AYZ3u6ns18XIuiuf8zGGM8iFmkJj/2d/FtPIP3WO+qFql2wQgmixk4JY6tNOY1q+3nhvzUqo7N4o
pK2gMKLu5ndEs+m9x0LsM7TbHTaPZ9RBOUo5ZFUewSz89UAwjhFK+ydAf8MoWj/ibpArHisPxKNS
6Mv2SAf2ZxfSUhxet5WzAapnBdXY+rZEY3e4qWbyx+JX5E9Z7KsC70Bl28M2kKMCWFlN48U51u1l
wqJkULyxW2BZwNcoSy7M6ROrai8Pdyc+lpXj76TUOa0SnAjw1+PW+2CXG/PRrU/op4z4B3EAsJ0m
MAmqSdN91qNty24VFLTLiQsin7DRD/7YNqHNEQC3jzC5GakGAkDN29F8BzYdXNP0zuOGGJTCg/Bw
j4BBDai3ZfhHg2L8w05QHnWYbpHOmMM+Y4RYcZEPIe/uq7ZAluqJJdIg4ArGdUBjY87E5yzW702a
biPUwGmPulp5lK91cqBJHpNeX5jTYjPTKc+WP5S26tWmhk9rhLG88j3B6VRob5cktRlWbrXMI4jY
mlOjquwS7kLSNeHM9qOG99wdH2Dk0pnfNnnU5z7A8BeJbSEqdtxATO8VQSy2uT7R4eVaTT6mcbjh
0136LWTuyt5d2VdCw4Ocv2ew84xMYcrGgh1UuWwX/H64Ox/Sjt4r5prQWrbVTVMa6/nOCCZBaD+z
+EiZjGRr6mq9K/uFjTkcZqKlAp33UxSmY1MonJMjfrlu/c9FVgS5vrG72guAVuHcZ4++/FRVSZq6
NBh9+xWtSKodViKC1EiPgL4y6aBIaFdCN6KZbSsAH5Hy6MYBGzquPKx8Rq9hY8C9f5Giy+vvhDx6
N8msZ/SJufQuWjcgAnfsYEX07UNF4rHpu2cmrtu8eQWVIkG9pCKgORNn7/JnCV3ekykaMvpqs+3r
kxNIbMZwsZtIlJ/sEAMNMcsXIrlMQyw9C7qm0E1HT+yLRoRKYo7gtNicLlRMpXgz7u++83njpZ/9
w8AO4kXd+Tpfdt7tPt6QCKkezVsAyBfrbopXS5Y4EoO2AUw5eBf39hKCkM6+zaM++KiGlFs6ISHR
oIV/8w0QqZ0Sh1tM4DqeJRa3BwSE7ezOHKQZTCzrblxQJDMi86Re7cB45g4vMpuJHGkk8+WUJAC5
C+tlxDgixTuKwsxqxQD8ThkLs5b3KYoFlf/cp4FkykPuOasHF5hPQhogrGEEaCytRzRo2972FFba
eFyoubBCUz4i49YnlyOSWl3lPtRs+Sh5Cq2WjrrdzJI74BykRS68w6FAYpoETqcUkl59S4F9gH5b
6F0MJBipsylnHT30O795KfzzNtf8Rr36MvSEnYoH6UqqXoqoZGO59QcH71OlkURQV3b31cUyLV40
otalUG+cbMZ36h9+eEomlvpXa+IUKIH+MnQkc75t3L5CWES0ASl34aIL7u1EzTrZk2tFj8JT+y5f
b5kjbyJbalqvDJ4Wu3lRoRVmPDlfhkNo/h7n2uegLOjcaJeqHc8Ew01oEIAbBaYDyzyyUiVo7bnY
dR1fQyCu3iqafPtrOAGMcmdcDqBcpcPo12cKmtrN8/kDhcrd0o9V5an+xHmEqHn94Su9q4PjmI76
fqaGBUnPc7BtZN9srBzFZaR4BdBvy37rye5dP9V2khBMov2XPvNTsxt8IxQwWyIvu05MfX18wH4r
6jJHzDBlnQE50ksgipVcplnnay3L8BD8RiKbA+KzYbw/Ysy7NjiPhHFhRJUxh1IxYC3LGl1jOTIx
oELEkHrlhiCVGPEDJwEL9hLug+RhCbDTKJY5Ami4xUQcMuGRW0mbgto7HDQuzA0yUPiirymZE7CV
cSPBqlgZlTHo7lLcejmBQcnAy9xzToeiAUZLEyHNqux0sOdcqPhnTRCC1y3+L6+nPddua2nyziRH
bsDg0Nkb7LPpk4+bUrI1HwD2035U3DzjZJfZSOCdeVrbTsj6vcnQPIqAT+pSp6BsQYMr8WhOvECV
yhaR93eX6ID/LYoBkqk7epN5emTKeI6tG2j83Q97NgTVxCN044SXbrMObgkequXZtRbEB6SKbNSq
L+Bx4NoT8pS+tjA9y1+mXq1/xkG9nQ5I0NLNWxv4BHEKTXnThivP6OFEXUJMbH80dm8D6fQaiIzR
VhMWz/JrDaCbht4+NR/ah0t1aA71ksP9ppsvpvoJOW+kyd6ljtfypw1N9Xtzn19jOA5AjAQnld8B
EYbSMCDLjOk+evqT0KaI7/P+pdgu1QpLxMB/OHn5HyAfDF3/HxSGZ0CxWaMw7Z6NgmAU5IOBNNlb
npuR7iQ0oV7CzqhxxlEM+ZjZ3oj2LOtP632BV3hlyDsb4S3YY8bjz0QovrVD6y7t6QWqZzmXl5ow
u8xR8lxm/4HFi9/GhFlsiTu6rYx/YMri6hjXmwi3pZt5/GXrtXiVmjlE7Sm6cEWavTibPZAAnAzy
v+82LRtjB5+POz5S9Wja/kbb4wjxxL3W6DkAti0YBuOwjaTqC5yoK8KCbpx2KFmQbBd3MqY1+ued
Ou/6HbuS2hi1TlxnaI+JhkpHru7HmZA6arBVfaVpNTjCo/SBfs3J4gKSVm+IeiAWPOY/rtZdX0bv
YqsBgYiaZCf+e/vy7fwfKDzV/1jRjjAlK93OmBpdJsmVvFaSE2e6VnIHmBxQjz8vJbxHWm8vKqQd
r7IBaytH9u/wtWnLYAlw6zOqgmtXKwqA0cE7MdIYcAY/gI+OGzzt2xt4ETg3I0fLkESRM5FEDSgT
EOYszjkzoDNnNtxzP/jqc/nRm9FFtCSEsgsuIusGMPW0Dj/JmGNQMvbch4yMYazIdZJgRLG9wSx5
MNWxIewocVEzW6rQv3a10ewjpeXp68pRmXqhir3iPW9ZMgNdPYL6fym4l8Y/FEs2h+O63KT3U6Ii
Bm7Jd7Ib0c8dREUKrOsny65kKFm375z5ctQJMsx/J0wJEGJ+p4gw6X4+i8g0f4JlXQGpbJUI8geJ
NeRkIibT31CorrEzVtmMnJoSga08gTrL7qTTpANEN0m4m6f062mqQW8CqIkx1FG0bWLDO+rZC1Ex
b6WpTVLWqRsc9OhSovt/moTnND4H1YXixunGyeB80zwopT4hNQQvQKvNOMSArlCwstYYbf310QJ6
ofqytxEQSg6wGb6F+2cauVECzX/tuQHTwEYNgIxXhtN6hF47gKqFzfr7X0OemJDIrZjcQQYhToun
m+J/NgGQfTAWOf1ECVaqiOCKY17GZRvCVmyCzc9TdLdWb3ej0+fdAeR8lVXqHQ0ydx6QU8EAeF6k
HwQfhI7TswczgbZUbGdkEsLwlluhnst5c3xa7rRfu9/oBLIz6S6ZmhlX3URH7dpZsZQVLQVLV5dJ
Ve1UCz9f6Qko+HHnHkxeQ5xcylDqkQw75cFYMBg0ps1znpsBU1AVXnI9PIDcZkrcnF7BBQpvYaOW
kj+V3IGk7jHIuZ2gd3lw0BWkGuFOg8+Pk1CGh9vdigdOZezEJUL8+cjrQwA/bxfH5Sy6QYHgS2xa
qRx5iTKIK4CCpE3LbGKQdqr4TyhswXxQ2yX//21TpEBVfHF/LpU7NpqQ9OQPLlhw+og0Qby3+XIM
zRMJ9CauoYqlgyeD96bNU29tuCv44iVsQ8p1F9i9WzFjC6lwu1uebw0BqPuNXRxrm4uvxxPrQM/f
Sbe9lFUD/hs6a0+rZRArnW/SF/uCPQ05RNjZD7aP3ZP4yl/AzYhLwtzoWZU24yAuiPzl6AUyGWT5
3bFINeVJK1kvGRDqusFNTA1Hgythexx8pNq5+cRFA6mIxe03y6/8DI3l3pzPvb3vcGlBBHVeat7n
uyoa+3jYzoSbKXqI8YI4H6DABjs4tJBTVuLtmdd/k3WfxsxhBLPBM4sk/rNYJZJh0VRstiVoAuxa
UHE31Wc0qjyErSJdkaYkgtW4UWn98qZKcizuFNqBGvQzqrZwsNHr66nBMdfT23rH4fSNgW6e5GR8
eBMKZkTd+jvuDcAv1x2QFhgpR3vLvSW/D/wBOLJgpK+Ed98KS35fvsNrefh3/scvlJXXNdymPz5c
DyZeITo0HfY/xXNFKA6tb+WeBRPHWrxNp9l+Nw0Xv8lKDOT3kyD0ySj86xqwSWfSpjwcXEwn6m0j
JpZ9RZWJUVH2aiGdBXJCzDyyuoan1q5oHe3EkdvNyJg63+dcnPeXnXPH5aLXfwZhrs0MoOkxVSrz
8I6QF859MmDzIFd6+3wSbYUBu6ZkOQkQkj3P6j5J22aSZnSL3NXDySARwR78BQrYQkVmB4UwGNaW
oWhQYo9rAvCRji7f/10AtuJW92Yv3zIjQMRKfq0XQ167qXdiARp5qMskS8dSVrm9TkkT+zdqxyLh
tFxZxlOmy4NXj+3LSaO8JIHGAHBYaaVw0gT3kHfi4zrZgf8PNYWwyCtp5x+D51nYGKS5gx9pNav1
S8ocAuAf8it9s+WDX8GBpe2nXomYt050uPXuWKP2VdVDDx4m6adRqmDt2YuDg+PNx0Zcs3J7YZO5
7Rx+xqH9Ntz2nAx/Is1o8huXevewuTXo2g8iFHzeirdS8AMTTsopPMOG4niSplpSAzY5aU5Fk1z4
CPHGFEv5/KKTecdRlbANB/5UGCml2oUGyBZTnq8yQ4y+LSpC1/1BOVSLSMHHDe1o2D82VA7A5hRj
mCCU6FQU8bWFkvD+Ms4slLGn3sfchjsWhx159uY6l8uF+ExdteUXYaj4pMV18DBdekblXR4enqJk
+VkE/EFufFjR9Ee8h+pAfjvNtK1F8DkMlw706MmeeAQZbKvCryUzI0fLjYtQRKVVAS5xzCYeaf04
8BDwdzFhcrUPVeXirHKDq4osZqbN/WVFGRFOGM4n700Zt8+fPnjdGo6nfAPTY5LnSxIYXNKT60AT
TEMxu15MnlyfeN3uT/HVaX5qhKAf+J9beOUhd8Ept02g4UcGba5uouQDFdbC2aHZPyzhCYV/M7O5
QteGJ9USOMA0QUcavUJHP8z+S+XOnt8uiRIztdNuf46nEQGvu45bU2RCLQmAjbqBNa+46aYotH8k
ZW6EkSqfN6IUvNvE758c8p52zOmKE3RMwEhcqhyYWqUbnfMiDvefpS/+msn4sD2tgmpPDcAEa5de
LiUBumIsfsizRES6aa+PAjg2XWo3/hGg7GwSD0ooVZlpQ/ML8uWH+uFLa3J2QeREGKa2iGsiuJ20
PXSZAx7kWR2ZL0P3j52/sw6rQTXOwrNgFJqQyJnFROeHQUpmK7sJIkDYOSn0SVXyDYa5fvni57VQ
lMX5S9Bis2tQ794rZ3w/GctLRgMjE8hVhV0dg6koPP5HyqX74rjBLFLgztinBM1LdwyboG9cFK2X
4LWQoVdnbHcA41uWdIZa3aR8bmB0A7L0QoyQ4DzBqUDdDXnavUpPPyV1vOnxXx/5u1K8WgioybE2
2RKhc5FBJ3ctVnc/IJTZ0W/sH6OLO5TH/j97+kQ0D18QZvaa/epcQ+6iC0omgaCXRayD1OeU0b13
uevznfRs7GQmZlrtFL0s2A/qCPiivNQ+Bl6rHbbrBXXoNaJSdqSbCZOel3FJEOT9zBENjX7XB4wD
LJwy/g8rM6XH2IhsEpMYgYA3pRtZJMxgxEHnAOudIJW4FJ+Ajdse54R2BpN5D9zk/LVzAC+Qkjvw
dDifwcPY/pjFWzpsvmxjbPlUjILHBhXX/83ZCr/S8lfuAHcMQw1YGRZJuzWV2Wnb8Y5ijUQ/q667
ayFetc/1tSbnR8DQWIrht4NYUJmorMds6cjRU3nQ0iyFWGZD6Rb6NLgo2KHXWEwUxOEi47G+Oamc
f06dNED6f2cymth6C1wbmSv55fZMOiczhlURNs+IfkyCHfktxMPhxJzLK8BFcVVSN7Hmdj9zt8mq
OrcUFX4TJhSSbBnQ1ojsoyOEfGUC+jK5/WShymfWXqwxUCi/tYz4YwGYbngVh06UhrYIIoDuDDtp
5XBwJ6lZG72amWrJfzjzr214FLnBFQg3xfX5U0fA10UM6yCsgu7zXQHvmHmz2tLshjTzRumaAbRz
cN/cEk8IUMzfSXSCB/Dbtf1+7irKhG9H82JflvlnfA6pRo2CXn2HUomDVC3k06sURa4qGrD8i+nm
CMqDE6wpyOSRssfpOj8O/nSSloUpJIFrRILULRT1wNuPe6rx1hTFRUE2HYmgebML08BZlfiADbWD
4b8eMUhlriE3nsTu8RHh0sPc0e7iV7Mpatt9SAWbJnHwoLJx8+Twj1Xj61R5l/pj51D9jLcpU8aj
pib1pxkM5qGGy6KqcuijVpmjnKXstknSQoAaxT0A6UvFSmlFulFZ40Vv00p1r4+gYZVAOh/2VytK
W6+2bq2TJLkE2wYqJXJ8+bciGjPAoYvoCnqC+iZdNI9juF5eznkua5K2g/uvfAptfFk8h1Ss9/Zs
itTnTdFHai4mgeHyVdHYC/EN73roSauxOfhleKUcu29Udq0qXpP9DvPnO4xUVvzyyRXtp4vDXc08
B7GI9G0of2WgfzSRS3Xi0RN+Gk6XMXFGtwVXXHt193gqVUeHvL67bNfGJso10Pe2a9yRBfXTOyyG
8J+eGlhT1te+ophxN0I1FoNjOfzIh9/9kshZF5OP3oj/bZxxmGTIK9WpKj8C5c0k8dv1WrAhwvnY
ki3snV+LBZPTaX9rVfKkdpcGyERARi1G47ZIbRgv1atQKxI0vhIBqZvJYpOI7R7s25h5yaazvUtj
EPwZlj6jzkMIn0j1b8i4esepkDu0jqCu3rcsKKqO21FRLK+MzJUlNv8FC4BderFYuP18zAhyBI+F
Ea21SR416iVzP2IZWMzBQZD63gjQ4zLv9pEsmlfB35WSmIFMo/imUpdwOoXfAK8i2YduJbmKfGnz
T/bYdLggLBijV8H57lthnxW24MlTb5dmz0Tag+b8j/zzALWLDLjX5gTxZAT4vwwjCE57g7uHzotm
i43uh4vSE1GIvOviJqloceBd5v82k6DZRZvpFlvznpm7zZmJgZk6wdNLT6yojDYUkbglRJqwPCM6
81vkjUxx/ugAXsckXmJKbXIfPNzImEMSTkSpYy5oWJyG7Od3Hdag8ZjuzeCcf/vpepVGM/t+69DM
ptyLBFUvmo6MkArjcyGJwFtu2B9GKfH49/uN/YdUudGWG/YhoqJ9r0EczQ1f1TzI0YyPeaGy0rkD
TnSa5lTti3Vtc82vVu2sIbQUo/dssnuwvXq6cWV2S7S5du+59QmDn+QDqi+oy2I4Icf5NQjCsRZJ
NluvdUCTd8qd5NKf9OTDvCIuXs8ox5kbQDfy9xN7v+0cALcjSw3k8EuNhQob0i6tlrD7bdNs5H6m
GK10KBBBKYeN/4FZwEyqf+/5DyUGKeVpMVTMkd87JJO3QfxfvfIOH6QUkTBF8v+436CBigviIHNb
LnQtJBgUxsv2btY2x/dZXIP8yKQHwaFrp1a0S3H7Yfhh48W3c4sag+oBvMSiClczteJFxXywOxUz
Z8/TqoXYbW298uylgZu6ODiStYDy17v/ox9Ql0ls67Fh4TRtJWwKlv44cuCmZciiAAhekArSDlkR
/oxr2SaUY0CDA8b1+h3fcbKC1UP0KTb89+J2kk/AkNnoSqTmL3C5AAXJSFJMyc63sprx3Ks48rvm
im0lBkNuF+7czrvEsSl95oXRGNEXOk6LHvzjTUV0UXPmZquzsDWeYoVOl9zYlvswlfkHI1iTdA+l
RvZMpAR3wvZYTD57xC86eLqzxvwXiUVMDSagm2JagPR5BSAUlGMj191JunQUSK3lSuswAoXm7A6o
V7HmfdqsBhq2+F19s90/z8McsotEsmwa7BjvTUaxpLGERr1ifWVZEeUpcyqofBizbb77fjgmKWvE
faXOZdjGn/HIFljnMBI0xJg/hX74XvGqXWBF0Via2Vjk2s7NA0OAOaJwh+rLk7dNPraxOdNdjkGY
tweUpAftZ56JbU2FAX4UQb8Rca9wQhYYOBH2k18+yoOPKxjpgh6K0xLadtYIeeTLW7zgRAZZtvkj
8NWxgug3GTA3ql77HlyfsvfSc3GdLkSRCUabnza3vOUL1mCjTNftAhqgV0+4YNqfL3Pl8Y0Z91zt
YZm8S37NbqVEDZFLrFxZ7dts3EwRgueTjgTQgCKiqPZRntjN5qVHQtwW0w9fDmKjDbdPUnkrEIOm
g7iALC4k+opEN2b+EM6qQYe15X1h5TNfkywRDD24V/wMlNzxF2XYSXIWwvmfCJEcvV3DvO+zdsq5
p2wbnBGUSq9CIrYB3ZNMd6XmHXgRFZrRkAL9EaeM/TxUfM8k5pyejkxtm5LTfRdsd+p7A89r6xq6
O7IiEzROKmIGUkbs5yVU41h+HVUESC7JutoB6wx3426iRcnp6nRvVIG0M4iVpkB8Cd62EdSJRcRv
D7sXXDm3nFno8j21R69fgPEq1zm6qqCo4gY1GTXuRQRd7bhtEa+f+E5tWMVkZWYNTxoMy9MNN8NC
d/y36Wyd4sHsVEtKQjit7iOm3GoBrtxnQ+RcwT9ahhPB/c2VVJqSwRqnLZvKdg7Z1xYGSp2sQcp8
Z3PG2m40weK8DJzJixaLi1g1FB6+EyodEnmL/6l0cx97S64lD0KjDqpraw0uc9HGNTl/N4DxIgLw
objI40d321KqHLXOvSwSAj4M1EXSwpXocsk03vYbR+JgQHd61Z1lA3E3NaI+3znyXed/Vcs5LoBP
t7ybDzixL616VvCzYwRQKSB86mu725cQMDFzDQfO/UIi0zpEaOWPN1XcCBugEcOJfHPWDAzVBXpS
A0Uh+23YliqGXYG6eXfwqdlU1gv8xJIaFRAtTMb+9jMJ4GBJLI7IZE/X2Bvi7uh7F50qkK+GUvla
YgQQAV/1n4Aon5tl6cJuDMiJOONuFVFGk5jui8x3HPhYa4ctMphhVJgF9Tzc7tPNT11XVRflHDlA
F57g5fSEyTaMZSC3ALGtn3LWcnERGkOtG5RXT5SVJg3Vugf3iNmNFxaD9fHAYN0X7rRNzIzzvka+
VVavPN18UdAx2L1wSO5Bu1++6ZdirXOAnPxpFD2fbJgMdEjm2IpNKLGY4H+UzGr0/rgG2Vj2QCSU
7yBXu05JBSexKZY2IY8kPBrL5XKBGV1ggjK7G4UnKnIrPgAb1Ji74lso4CDHzZsfu4XlzvF/1f8k
xBGYlz8COChO0jW1uF+2KEqbBg3EZkyN11+p6lkrohCHO3p/uaEvkTIPWq8PS2MAcCv4oJzqB8TX
Nrb2gO3tkjHxktExoQ1rSZtwsOwmgltVhJ8qnxvRuuPinco6DlOn4tgvM0hTF87Z1r+WymqZ5og9
n/pwZeeYWsbu9Uh9ZgotZDp+pe+GVedlMjovAeoMqkuATgRqExAvLHcpn0Z69vpcuR8IUxzidLvY
Mcqx6M7niCdwnA4cmycuPL2Kt/QXGfRmAEl1QVN5GP9XudqV6YGbrPU/QLZsPwyb27VHImtMWUeS
BNAQOr4aI7Al62MC/nTMg/EgLNsjrFjmLmknlXjHoIm/Z6+WZHWokOcBPNRTPGKt0IfnVCOnNjS9
/jikgR7uhW3ajXDLRhNXHKW7zUXMdlWqv//6+OKI37AlAqUyQ5kDjc9VMg1OFXiKI11PHhiczcGb
pWMr+GoC6d/IxATGNDA3MBVnO2irJHaOnh20F/tguhmugpc1yBEmNiTwFtBoskhgBrG5bwG7SXc5
rmPHVah1n6sd5wjjDfr70uH8X+DW1BroREwdYq881+fiTOyV1PkP8mnCZ6ES/wkfrV5Hn7wAWGxh
gGSSKAniPVZ6t3VA+WuoSEf3WlzNp83OGPZiC4HfmhgwHgQF7jenojGnnN9Qv7Jpd4/S6FMhJGTD
yFIr+tRXpBja+WegdUhdQnEzBl9PHIKl7eUwFcZQ+zum/1EaSyCmkwGTNLm9bixfgmIyak+wUN0v
uvlq+PfzsvZbeEIaMOqlfxjsmqrzHdmqHvdKbuGPCB6+POacS7tsv3+g4StAKvSP5l8gDYJk9J/2
A5Z0Ln6JTdLBYZCGZJd4oHlR4R/HbXDJtWkVQbN57QQssK6oG64dahWjj7c/u2lzIvIvb3INWbgJ
s7YkdPyj6wBp57Qie9O1B01KLqtzMIo5FcggfnUzglX5lafhELCJole2HfJMN+dPAqS+/TgXDA5E
qkPhr6bEDqHDrcp95DibRcu+In5lqDxI4AVeK6gBu4APSTtrVW7fN3pt+4ntWfeRqVw2d3lTydpr
oseY6ZWRQ5SJDXRC3qk3I5Lv5whhQQXwg+LZNbDEMZiKTbbw0aeKrYUM9zCSYFXuiNRANh+XLXhF
5kc5NXJLP8iE3Nfis2ZVWnuDk1iv3H6UgmkxPrHS//tEupir9XeXYtcu5Xg9kaLaXGlssV2LVv5Y
5pR03Y3gWPZPf+SLDf/pSB5isgbEYV5bBc7o7miRpUIotQIxsA+I8ZJLt9wtDgr+l9pnD0Z2iUwH
Awn6juZbPI4h8jUdqvaLD8MuXZ1omANuwAWi8gyIduHY4yg1xyniszS61MsGLn0y25rXqJ+V1vMe
PTHcOxBq9Lev1s9EI1Nf9Q5qoYMJupI0eeBDDwT1p0lx1xYrrOEPyp0yu+8axODwxOeaa3SMZ8fk
wtvouoM70lv0AqCEEO07c8C55MwV3GA9zudZ4LGJpiKDgUmFCyCrJYha9UkGrwSDs4wNKX3+aWXw
plBIbmK9q2FqLGasfBbLgc8foDM5zqOfdBY8C7SzDXUa7zyBg86XBAXMXSH4KwthAixqI/dXJlGE
Aripx7bIFpwSiYR0QoNVDq2C7CAVDdQqUBZ7CLg6SKAHohCh7DXnwwzW7mpT6udBbXWmao124PSs
N9E4xjuEWnw7knU32gFfH16hXblmyR9cEb/rTQNj1iTL3CfajbO/HcXMIRey8CYz7p5P+/s3T45x
+nLHTQxlk86VSRHND88q+UcxA7GuotEt6I5eeuG3T+9kyvIaMaS/pXaeZE+Ka6R4cee+FoiAbsGt
MHV5DH0NO3tQNuK6jJjkiId8hllXty74XLoVmjyHyc2hg+xeBcM/V1LhZKAaIkpnBaUpklBfZQYJ
Vqqs0KRlUiD2kf3jcjqFQqibaVTqDWsAD1p/xfE4GaA2Nb98LkC9KnnIrQexKpUljW1JLC8d+ZE3
Eynxl3jq3OOrQkeENi1z11C+fl0pPzavFXCrTpvrcJkP/n/qeWF9Bv/gmZb52BpHpvalRBSPbWkf
2xPMcLqkkrXFYlhLfpzviEhE/4uLLuv8mvRV/A6ewtjQJRIm25pZqCncsj7KXewHYAoccqygb/LG
kd/nwLLdsLjmLOJ2O4/hVN9EaERPFHNyBsYcyKMBBwdHrF/TSA8Q3Cgy9zCoUKeSLviYoHd78eeg
d5Ga78JNqgaQWOM6sXvFEEuyatxdlwdG5vucTcCYnDDMn7VJE/g2usXNsOg1CF8ftR0YfAtdDl9K
o6cgJa9yD6RReArDguXR58xKlxHyEDKK6B1YsE0HWY4rHwbkVPQow9rbfclVXHKW6Q0fUCA6SzCk
YPPSMyd4OZIvdmJdjHAogX5aHDB0xPjWlkd6SvYr2Mss6p8Q4qXY2yLcSHMDmKhpKOg0idE+j4NO
27vcGMj4nwnyjBFCsezQtaJDKGRCoCQJNADt5dTPihX+TbLUuvgUOK7RlM0hTlOrwYZyJQmdj2Fq
JbcfejHkYfz98d5LDDj+vdI1Fnhj9ofiimZBx+55qMrGfCxjAFpMwEDJDvWj0ht7o2bUi+sCoAkD
21puXSQkwN6xMYUlHidPpiRT9iZUWy6TCtqQ8ir2eGui126/spVqsAw/YFFEEQqm7mmVtbT6Bgwh
vRiGxzvxKxNQRX6EVXjFpfcSNKraqabnikUJ2wWt7s/YBg2bl4wmwKhJSDNW+lN1ryjo1xNPLkau
pCHF/P90E7owt1IArd3mIFsHGkmAplSb6AaYOns+kZ7DG3Gt90jvMgfeUN+OcjKHECki37QTV22o
RyiKuClykr6IDMZwgg0oYQrplW6gazuj8gZthIdb9rhrKbNretl9M2IiReGjab/+v7TkZozCQNG1
nY7WyqPgYcJaMFAe055XinFbcQ7Q1JDZTcgcE1iOYwt2AN4Br6S2dYlZx9aoLAIrs7zbzEhqhNFO
NPQ6QWiDRbm/TY60zDioGuMxr6/1vbmBK9x42OFVewDZkmhGTME9o90eFrcwH/vtt0Nc3yDNX4ge
oBXYQdom3DGaUbPHEffGJz3OR6ilNsPb7CzkgC/UXjqFK6RtQEXicCm29TiulGszb/VcXn+VIQS4
G6197Fmj+TyoTDs1SP4ScMtiJeiufn1L9kNWKbwNQOZ4xvlCMmTH0tiOws/Msz+SRP0FNQ9qA3TH
6ainPOwpFsFAzKy7PKyUCFvYrSoPjI2NIw7Sv76fKjn+rpPOzkl0R+OhGOzUD3oLE6zyP5T1povO
mexlnGpRMTWLrVV5CR02ZXZVN/4ivY+ug/+d5uxo1+UgSKaWl0eIFBZnn9/ea8yzme9/WJj8+F85
U3JOt3eao4VWDqgDOsWFHPT8Yq6TjPY2TZD9hSJdtlTdnkbHRDVrw30t0vcpRYMI33KUVjviWfcL
XLXx/YQRBiQ9Smdx00RmDA0qu+iCiBeh4w095ON84p8u0V/gPRTEPgHdRwEa+e3rqjwEWgK9BYz7
LlYiRNaeQExVeEClps4fx8x3xjY/a+AwE5X6ihWBzQ+OS08Padgup1WhOEcmuWyGr7QSHCgpJcex
ccdhbvVL21DaTdyCPUNNCwPcfUh/1cxcxTqjfQGDtt4+urQHINYQGhOosCIAbMgc3wzL15kUe4jF
hyvQ+FIpR+V7473yfxEp6CpQiQGCYwKuU3WknuNp+v2qoJkY9p4RCo7B5dYCewpiC7aMG87wVMXd
Vg95CE51F7vwC3FYcs2J0UEj6gusoxbGMAtH5Su7frLKruwF+qgBGyMngtPa6uibk6ez3joxJY/j
GkjEtIwf9X6prBlmc9hn+e5dZpt0Kf4DJiIyYzqgT7vAmeA7zauHVjCwHguwZe9dGvbEt4/oSwCt
H2PjSwBSJAHRez4b+B7I1hpvpTSTrvWPvP9dQ01EsfhzpYAyfQACs1ng1I5wn6BpgJY9bivgRdX2
UiaKt9pQWt4A94J0w7ARQwGXwGTRn9hPfng/4J3kQ6E/OrcVOGPsqE9DvY01X6n9PfxEVWLDtjMW
+TkdVP3q7C5AwyIbUH0QS/bb/Ote0AAH3DwB8Bg/udnsV4ZQCB76axDwLoNuS9Md1W03bxO39/dC
s0O84iAOh8XMEpDMfuMJaVQcYyHmFxpp8ocNoFWKTrkwquoSv4VfzcU08aKlnZsTQaYrDywdtjvH
Q0AJS7DNrZySo7yAr2d9UxhqLTr+Xxhd2o8DSX0Q1bu9gAPTHJc8s0CkwrLzhvPGkct7WrwGAumP
16TnFtB1XJUOY8Aovczy2iR0u5AbctuB9WJIYOTRb/xtMv4Bg3Baylg9g7O/UBWo6ACx6VvUeUj4
r+gp/zH9aafNTDmDxaxTjYOzxpmQi1tqx0l510Y0b/dZJqS67E2O+jmZCOh5ZGkkW6WX2lzuTJRz
CtDc3XEXJUvPu1MdL/uHHO41mpFc4yoL8pdDjSW4rzOicJPCKGAyKWaHsgl/49+tY5QLvAX57u+M
Bu8vWHzvkBYeXWPKSq7U6SJ64ol2GJLY5y7PiDFXS2K0WpJYcfdY5EBTNEnlAQhEbUlIkkBAnTbW
9NW0oQdXvfy8ZJWhL4AQ4Qoi/vVWBHDBsm2cI2+YBUZMkwNMu4+0Swb9p4bE9Uci7uDztoI2fUBM
0zaTnPjiiKXAFybq/gGdwLaDDoXscBWsh9tS0WjZGkUE5aTlcHdeTug3x7LWp6G9YUrbjgF8UBjW
ozhfQyku59ttqiiT6qsKIrdzfvxCY8WWVw5S0Y84ZE6evkKadc4Ht8PY/G3UokRPb54QalvAv0J1
lbsINoKAvWT0wyqfSrM+7TuKpw0CbciOOCv1Kzy4ZLeF38FriJDPMD/KJ7jexB5pUiLR6s5NhSfk
Zsvdlof1sXUU+0AtLLbaKNUcO+fWfhTr5zhXTly853214+114rvmF09w7fCdYvsUgGHxorbbZrda
e+1tzOzHrUAULi72Dfm5ko3Vz4vF/b94nuGfP3AImuQ8hFtjYddnawxFngdIe8Q0a/4ZUqMA0Wcl
XCM1JeWXZe/b45wcOEDznb3XYAmfQHqv7s/5W6QqOziIKyvC8c9NbsvpgwLy59COGENtZ6qzE9nC
tTJhOVTVhmMm5Y/Vy0XZgb5Q7e4pArFJ3fz/tdcasGoQ64gD+uA8LNNxMLVD9XdCdNPZTd/pIOIi
4Bhz1gswAXZNODx4odhy1nvXagtnXv9Xh3wGW9F2N+nyzco4QFTkjrp9XlCCxMWk6nomK7sXzAlR
Ea3aR7LAnegVAE/i4H9Hc2J4qkjt5CAlmBT87SWxe1J/081MqQOts3+/F857wOYEzkrsQ56t9J8d
W3YcC6s5TpOSsv4cuEQUrASUNQGy8aXbmE+x3PYeYP2FuqVIwRq2RF2a1Lb8vdbNCZAh4jHSAtV1
PSi1PbdBcSOgDcajR3/qXANGB9IOnJvppBbvOkraIWZkNMWuEKDdXOYbazxdEyKSNjvo5id9804+
RsgskcdHqaoexTWD25k9T/jT3SJrl5NvgnT8/ArJzHnjyjOf+CxUXQPF+2NiB36f4SAtFE8IfGBw
9buS7AGpZvnAFpbCnH93W072O7XwtIs+ydTb3JKulL/osUFntTQ2cgph/9bTfsPzwJUSc0GFQmsa
qA26XibS5z5p/7Z/ac6YAjtRKVz5XjXt2f8J7IXR6/CW9fRwSSxpPcKoZWy5r4opSJJItrAdQsCf
1wsIhPapX6QMgfqc9/0gQsNnDEyAoMrZF7WZ0yFbabKihUSmB2qI5jUYS7ZwJ3O+MbOsnhAj+fCe
MJ6IELuG4NqB5VHBoWxdHjXuSMWkRJBxz63OSK48fq0dpU1dOfu+XXZpYTZqV00/BMeJes9KK7c0
SsZgGRbAmKOPjf8DQExDzZjzCzXOi9B6BHqe2AU5aGIRwbRQlXdfYrakluisFlWItDYglS5QMlp+
uHq+3t2fP7nN4ArpZCpNxhv+/gIJAhYDGVxPTgIJSD3yy+AuRBeatWE4zb4XlhB4dY/sCG8bEYNq
i0qIVqrMFlt8JFGjR4UcLFbjo+OHHthGQ92+jYWLH41QhLnMuvta0BS+hAQSA9euLodB/gCGvtvY
/Vc+rXMVcQXovcaIAnYi0HbUkSUUDxPDioRcMP6+x3MZgELqZfJn+wLYHpRY9SwYHHM+UpHOa7+m
VLm7AaXJOh9Tp+pvAF2ljC+aQfOecLkhT5WieyUjWTLwf70HX3UKrBfvzE5IC4z88xtn4W4hjTqR
tX+n2bKofYhDBAKrBfqkLqU4VbHXcWO/GN5Pwn05N5zojHV2Wf6dwp1nHYbP9GQgrxT+NwtN8Hni
uDrsn6wMBiIfqoeTpQwNok3oixdQDrB/czzE2iCVV1zqwL+ASQdE877G/Au/SOBRmaEHKk7Tg923
fzW5rA92rSmM/f2RguTTLsEA5206ACEQ9htURKgqTaqsXxWUeyUt6/L37obAMBMjBnKgNHn7UBzt
y1hDM5pF8ltcVjsU3hDzPBtG5GZj4xV2O1NrQrgGcEXxu5Z+ybAtwEIVGirxBmSyGfyY3skYExua
CUQusdt1kNwbk8j8b4PVJKJfYyhIw+ZJY65IRdP14eHL9vxtuDOwHUdtXIl7eMIieByPo99/LjHV
Fm79niO8g2fo14U1Slm5akPG82UvhvgwSWTYdKY0MTMaZbnyFgFV0FIgEEsHBnHMrqQM7yhGoaZU
Frx68zX1YH2QFUW5k0nWVqYE++9ALX4tUh+kHmUBHNclvXSdH199r/vizC3ddFOSGnq1wOXRGH8Y
AHqqkXMZOBg+BVduqHGo3Ic3VYhUcLAY50a9frNRIpDhwGCKPAk1mSllCeX1pLhEPpfPne/+/gp9
Jv0xmGaoP5SUWMkjR2Sx7XmBLfXEAih14vmm0VieFz17XpueTwWYLsfZHD1x3rsXdd8eQw/S2qQo
d856NA1FWHSPZhGAkBGCjssZli+rNM420NttBoq7MSUm0zhLk23pbzm3fuxzwnGJGjAoqh8+LqpD
lJCD9aEMF6b9VD82b1dWumRAI0xodbXAS+XMr0zNEJfoLJP52TEizT/q1H5blHpYiO5ZukWG0CH1
eypwVJIRwH6OLSoUHOjmloPAmq2o1/RiVvzG3apI/GDNRjy0U2p8Y679ebEiFEsoNtsBcSL1G7Pa
j0MlEwI6QA2ZAtNrxlT4D9I2cBOWma3+iqivHkyFl5cEeTydBLYgXa02Q0iLtaQixspagYXUmBUo
F8MkaozsZXT5yJCqy8Z4zmqP1fOKQkXQPEjjeyEdPLgrrTfvQocQIlls5Pfm+dVEuxWM7xwITw/a
RmjsYPZLEIMUzgyGW1vN/AQJ+3tXqHJAFd6pdia79L3+oKnP1Y7CYWbrdnwNVXBsspBGHkS5MTTb
9vsXDSucJZsck48sy0SybisVNrTJzjwm5xKd28ImImWJH5Eg6R4Q6wS2vX56S1wPpzaB7ylzTXl6
BOclXw1gZKUsm/N24J0QgHK6QKviABCezPWwEgFnuCosklmd1wd2LMQQQPkVHjNQsL1vlUv+K0NB
52ouEvF69pPZM8ORhhUWVK2yCAzL9pkLBIvwPpwnp/oeOCa3dP2MNOv3a132IDtXdnq290kgyYNW
YAPRSFWQzEGFNKpcS5R/T9kZqt0jWzlgTAsZoaqy75NTlwq8SNJ8QwkZyiIv0ax6E7GMYY6Kfa5E
xA1RHAS02oD+hKl78VIbqfxaxQUyvs49wZ4BigGPoH0NFvTbpH+vbllo1jap7a360s8+mRO4amVM
56sinscpIR48hISs6wbJVnFdc6cvCIMsuhBg5vo8ROknVB9fa87zGEYy7yt6fC11j24ilmGSFTON
Ico241iq5TXLWdzgWiFkXYmAUPJIBtdfRyw7YQCikXd3Zfp00vxNbKp65MhIuFpBE0ch/sXLRG4y
ssmJtD618ZSxeY66MKg8/AwGvAM7QEn4MI1mpfGPsUaQfq5HLJcD3WD0+m5sSne6MbHwamG33BSB
ND5q3gYoBp1ZWmpnzg3hL1DfOzF5PPFyo+D8sKF4Epk+cL3Kwkok38ObvkswS8t8YxIKF/12il0O
2GOy4qDG3CAOrWmgCflBMGBUvMtN26xXfk7WW7Irh/cfpo99H6D2eo4gEMRKW8XuFhNuRCiwEv7H
xPnBaUui+gvOa3ybigp7BIa3GXGBE8epQ8Ol5DrO5GoKgXRwoQVY2Q+sgrC2pZKGCdIOWv0sFGIg
qVLoLkuIXAn5gnGRMW1UZKRKyasEE8Bqu7DxxizuFh01ggRJGwmKP5/zXPFtrsEMoDYlPNatq7M8
Z7KczrKISka+kTE7IW5iaqYVK53/VnVmHZbqPZYYACQiugvDHwm0YuY9nh1/AJsEHet+kqHcg6BP
ayxwtV2Dr2mhOpxixaMuHe2XKOE01YkYpTRIOlF+eI9ccmY+qbvCd2nTd2yzibMSugi+EWAhvc6Q
ps7Aa66/AhAftH8teZJFGK0fXFaQgO1LNyFOB8wEPloO5TqPmu1sEJ4upVw+Nno7oIkIUUx2UVEc
TvcWblhRTcyWpAt7ZC72BaCekdHBMMQzHUN97QF8VU5azoT9DIpE1aqgxL/F7Pn/9CSA7NUB/6NW
u9h/+iQmMe0ij2r0WTRa3vgLGK+0hWiWpRpFn+994JBk67e8lRkHT1+FkHRsmHQMWfuckeTiRP5z
IZprxIOLNET/z+i672crH8C6imgHBJwNYQdRfCwrrCXoaT7q5y5ntMrEUwx5hzgo/ukIUO0smLCO
Q55N3yydNopEfym6VXVxu84nL2mDFQ5RXdpWOeBZR/+NRNq+hj4gdzAJpFHjrGXTbdWeIQ0Bsy6X
1lbBnn/Bqvfet/6SaNwCJoeAQTxDdIs8qkDs9PHUMMvTiImFnm+qTDFmbrhC4K5fT7UfOU8IJp/O
tKkdz69SuCzbZbIYv5kjKkmnhzSXCQDK50p6RNYNg1aRTpdoMX5pE/bwyyEDut8OmkCiQJ93SByt
tPrBz0GXZhZm2Brm8JI/vm3Z0gXvAWrwZ87smXp1boXCYmBhHofQbB7/Tr4AA+sIi4q4okfvvhTz
MkA9vkgyY/mWN5WtY1usveXuEBZW9MYlNx+qBVrW9UzXZ4KVWXqE7IFUuHGw0DnY8B6QPkar5QKj
+fTQVvJP9We0YSNFHv+2Pgj5ZgAkSKVzUZZ0A1dAyRuehl9f8SX3hdhRX3ntjVbDE0IXaIDTLRtR
NehD2F9xCc0ldy6XGjQPVO/GtbB9ZsLpSwmo5bpJnTc/0THrJYfTH37/P5I7WUICXRADYvG2Dzcl
drm2zbp3TjhREA9wnO8fIJBRC3sY6pQYNZ0JXOK2M1afDUAe2hLaYdUUFYRpsi1x5DPOzw7FeNri
O4jyiUw5wxbD+IKmVe+BwlBzF0y4wm77Gtr/mwJOwpGBFc2di4YMzTTbuv2pg3d7RC3JSmhVQa2I
ntQ5PL3DgADxhl2OJm5anq+9zScPZJ5PmpYjxsPxtUL0IXfgk5sTmeBV9PvIA/GugOLheZWMUeNb
WuLiif/onuM4kuvofWwyZY8yidrMLug34rIYoIAr8e7ES9BzUfg1V0KS3R8RKMpmaV69c15WjoJo
V/nBF1u4Hp27ds+EVXNeCO1Cj0wphnQLvV5H/+DiomAWr3OLDC7FxcG4SyJrLnXWFOBqAVnc1ZKP
mJBjavLCbNvuglB47yqP9vi00IdCnyp3V1y1yUJ/piHLHi45njRmLBmF2AKFyZ4HRKxXciyGoPIH
9ffZrAT0XXETyBlZUCihZQ9XVDX2UaNOfw3LyTuvfgSjrY30eavlwyOtUgw3nAN+kCsVGZriKL8F
xToETWjfTx9Oacl3v3mkWmrQ0ez78IhdlbPxJXNk6j2LMguW+YaVRv8B47228Ku8hvPu4meikS8h
VoKPgH9xrF/LTvo9yKe3yrm3hS0RyJ5qpYOfM3DfabX8Tu8eZnR0tlWxsLjT9MUFkYjfW/nRaQDf
r5aWE8w+zlbD4zYJaWDQLm1kmpsL7lJEBnPQkkOqs6ndUKPItOsuMCi2ldQ1dwnrBwl7hN0/PRhW
6VpyqB0/19h+jncSdiVDsFFoJxUQ9I7KG0bhjiqCBYQWNINQnXyxsgGPiqETeD7s/3M3RpFedGvH
WsPqtQEO3nziOMCE1psMMNYYtuYKOf1sZDbHQrF9a5E33uYtjf163G1iTno0eJ1BVGYrINnMs3G+
r9Ruqn8VsImAHWiH5jCt7MAS/m9niRJSqgTDjgyzQV94+uHi4tDHXb8pXc4pjRrdXExj/5DD6MvL
9gZlsgzX/ahZ+lbSEMI6RiHYdIbhK8HTP80jodtZU37YWepDiI2X99sQEWae/0L0IGRjFI1ncwVf
deyy6mMjyQpTMwOL4nLfYFd7XGEufek+a1Cv9e1HxwiOvIoqQ3dG1V6uu+nU+sg8aXkk+jNVUi2d
88r3nj8MSkED5GCHEzZKgvFe7wJFR6SX/gaM3gk6dO/CU0o2Pe98LOg5GQ+n4ON5yo4InM5dl90G
OiPF5T5fzF6ps2b3SMOT4C9iQc8AuJsGqg4HnH+d0IlkSR/+8M1k5dTZlrHvXRsVNayfA5nWaE5L
5nr3h75bJ7nJ25zrceYYMMIXHVDkHmG19BNERpjyMDDfVyXXYR7yZY4rKEA5Yi0+hwXg/fvvtndR
15kEGBtVm3L2yEDaMnq41xxiEVakKcwubi3OkDCyAEQOnccS+EQZM9PT5c3ajm6EMJ/WlfRr8a8d
ZYo5LVq3iFy+ng/KM1VJlgdSlr1Bhu6yT02xasIyUtLBFFOo3Zc05u2AwwI9YKSV6L9l4ensm8xZ
G+VBEQWhcnV9xuW7qIo3Eh9urZ12DEgmrv5km6WrKEHntthbXypoT7Q+4WMPuV9FN0rGUSfm0Kqk
+xhHNjaYt/9GKhCMoeBZimcsr/OzYmmEtWpSejRikbM83HpMLML9WK01eJ/NvfKO3V0W4n35IU33
VuRjH3IpW1yvmZohrx8TZli6k/WAUkDTmeIZ6g9zVuRzA2CpYQ46ZRwMIY5rkxXW0OyLdt3Oc04x
xSdc9br0CPON5IDa5VRFFMVbqD3EfRbZehB/ugliVt0TCqqc1Jlnl0mbi0Fewaz96Dh1fYoB2FFl
jln1uSDS6TDjvo+5HjnO9909H/n1BE/k+UcYfiEqMPaRqWeHstdHt7o8FEug+gmCk+W6QR+EUXtZ
N2ctMvT/k68Sio9GmWwksN06CphymWgFH49GLN/X34n8nUDkJJz1sTp+QB3HZmW1i3pHBE50c2m1
e5YEsqySz36jw2XmU+VQQ1o/DAse5mcTT6vTrUBRnQJzhm0p+dmQ8dlyh3wicmPwauRlpqzsoZAY
BxARB8vC+eNIAzyygiGz1G8cJVLa3w/R0hk79mEy0dax2TqF1emvcE04ozp2bLECkh2RNooHwo7R
+08r+R/xRUrdZ6W5vxIs554Hn+AfRyZ0tJJ+wt6dfk5dPJ14fulw/Q1wb5PQZrkU3E921TogdJML
G0+ycgFaIENwui/gDE0KIolHSE/Ex2pSX3Jof7pOC31qnI4qkprIt2iFaTYiiEz+iMyG0qHPpeKF
RS9LzvSM1o0dHAtwXrTaKwyOfbt7z7w+kBD9S3LYkR6mUUSt/FgpBgXJSOrN3GEtfORNjVTu7/gS
eO5TmhTO9Vloz2Grtx4I5+roWNf7rSnA695VshyHUWa/PblwDZnwEJIAlpoMZ8IOUBiXdv8USp6t
jMYbxD01p/ygYbrwPRd4eyiI+uG9rd0yKES9Z73IjboYihyOZQgMjVGNQJrhqzQ/VQOSchVuwYtT
DxPPCYSrv6OUwLgCsaMwIGqR8BXcrbvtKvc4dvP6lIHTMo2gAdObTG6q2LZlpQh2wHVZBo+bVlMK
sZq/vo+Ybu6JkpJXbWFxCf1LySxUoiVoO0GKYtLMlODzW4rizTnNmyJVu8gnb4lmEWTBpmybGTs2
KJMJvDB365iesGdtXEKkto3fwg6v2aIBo48DYorP2g8JG8qUIjSJfdWnY+4AkxBXZM0rCu93OsuF
ZAz+71CoZSQ7GeLcvPUe6+rOXgiagfrWQCoPK/s5vP5hjwCvWYJjfwHHM+e4gSomREIXF0PRdIQy
y/4GnBdHXST40cYUNvaN+D4YFlEKW14kZa4SR0ecqBLQHMdq7NP/GLWXKVevcVri23ZZImS2aTmx
+Cja5MmFvaKJbla73oliTl0BHT/xzJxGqReuI3gBMVVh5N++fmLB47rrWpjrVdR853L1WEcF3tud
9ZbjIrUxrYHAOOqoj9HyrBU4GzTpgKkzB1XBe0SfQaDbgtvTqeIoq4HQWUya/jBQ6N3efuMyEkf6
M8EFodstjV41YMWf0o4NI9tFP36DUuWWhkaOQrmjsC6/nAPNPTZDB7eFeqpkE6/te6OyptjO5+T/
yx4Dn8oCeb8u4kAbCVxm/v0HJUQnc4XZ5SqvxV1p+O+lqmfzyyknw4aKsYrWzGHxn7oxae1To/rI
/UPAEfUQfGmPOsVzLS2wMwhRtq0KFPmOZLc7hR83zARnI+srsuqpDG6YdBUmW5xFKGa8gecCpUEL
g6cXFwVa1uZbunv5WoW2NUGHulbR+QoczUFQjNcxQxiZIHbb710Jo2MTNFw6lanRNnFMFII4shSQ
g5w1XY9SwhkT/KJuP9PP1GUeE8C1V2k5Z3tQk+UPgLqRV7AsLRDxQ3c/BovyLyNgJZuuYneKrc+3
ybwOObH/EUQUsGWLdgpadGX1ANFCCo1f20WoZLRfS8zl9bG5GKYiohI4yMjM8jowzOfsI2UTQiP9
Ymn/+obXlSB8rL+1oq+yn3mN+0R05S9bfxCvrOUToDg8m7abDnTAbZfg0oKlmz/7TO/Jy+qcV1dH
t+LQETTrMNs+4h8YZtWj5u8GiSEM9oprRjIeiIrpuZX8uCFMvLVg65jo8O+Amdb02SdSePVssGuN
jz7PQHAoASP+U29XMtQAT+UmqTKqquQ14UkcsCx512qYTKlRhDKkaIfHNfKinzCx6NIvvufw2rV/
+IBA1sE51oVQu17Mn70t2G33W72PtgqlJ5YgG7zMzExBx/QmC51/Ew+hqSYDLXNiZfRAQUOjc++J
MVIcArPCiVqK+SM7/aTaxnQEjnP4nWl8TaWzSQoAQDzeBU1Z40nNvHJ+rjxcWNoHoasaSZe45/DV
2DC30MlPg2XZTfHlE+j3e2Uy3x3e3UkV3Ssugt688w4FFKm42ojgEi1YPcpj6JzOA/qUiFG8v2RG
qr9+4+LaKssXJ3wCxhCw3ei1Ig1jq4/y5z3B6ZBiejjqdrgAy0vOUyR0RgVLsz634Pf8+IJjzl65
I1I+BPR5AyLsQH1iSMRdtmsFtKourhe8JRTlmMMm5cPnwUgDmqu6DB2FSWNf8rz+KezIUoLMycqv
0tKdwsBPvSlN2bjiZI0cNVBMtCokEr0D6hVsq5U3Bdt80GESxWyV9cc86E2I+zKl8RFTf8qN6HwK
7P38zjFYG3TF9CzPXScNeMQQCqpnOMix1X0mPkMdWkxkJn4T+YGBhPzRbHm3OGV1iUVJU9B2ljjn
fY2Oj1/kYISfC3MbGfPjNMVV1O84IKHWtEOl2JDULP8KG1wGo7dqJOhJdo3hjjJcqGVP5w2tR1hA
LUOX7BJ8iQt85rlucsDSdZ7YgU3FuhWzCghHDI4OXNoOaZxVnl/jQ9IPEI0Y4o1uoCDulNl+hF4n
D1auxrRCK2q9CQx2D4Qt7ogQQgndRF4pzO6EmWCwCSbGqOTXUnA/LiD691DSdFQz99goyb6qCytT
j4F0WIV75YkX/wUxAIe263jEAwbA78610a0wIIeg1+mk7wCY0MkENXR5LmzPO7bEYlR0Q8TuNPwV
BnGEkL2SxKGKQjtEMk16h9aUURBK2KH+PqU5w2fqWjebu9vdJ1e4VpeTWj50V/bA6ut0mFV65D7B
/ebXng0LacAy4c5GHMz9tqTczmLyVH6Pgxeadq23AlI/kNLwXbw4JiRuH5ygVAWduidgwLbFF3Xj
Wzz4jLf5kA5+Rauk6/tFzpbVAxDE/H5e96DP7ytuxvZDezDkrCx/vzcWXcbTiOilKSlqKTzYPqIe
g2rHXDwE7qF3Eune5MIDSzKUr/CTeJ3TUuLhqA8I2Fa/SRwY5WNa6ngL8lJaZgHI3BM90m15LPOD
2W0OCfUQJWlsIfZCjCQwdnCeOblxBsDB0b1DLM42QftogJ4kfZXHhPXyf9cgH+Q+nu45ImPvFnWk
DeSX0Z4tCP2hKn5bV+InjJ2jzCHousJzglw9nh1FWSSMHmpYpNrCQ7kWaro6YxMZ8J7uzG+f4tim
Kncv5fuHNI7dzlDlSargpWtD+yAuJ6h9iHTbF8elMHfLnuAl8X/O0PKGIHfZyznoqrPaRXzGKour
6KNFH4ll6CJTwAdFPf/Kcd2AWp63UrdFqBRNOccCAmrZjDYnLkBO9tk/2pcIjrSBw+/T2CwlgSnx
gNvhpUOTSOv9GnnJWpUJ4tyo+Hb8glbdunizzrKTRoJafJgKpFX69oog029c0d0WI6wNfq+YoJA9
ImGI+upJYEz+WfOl0uyKXg2KLVBcapf5H38EMFh6jNoSJdXOf56ueMuc+r4TtcwPg2V9IjFs75xs
wIrdBtAy3b38WV0DSbQc8IQcPkeAo6O1DxlpRzjxbcqGha7/dLtkHm0etQ7582u3C976jSHaZBqT
5NHzIiIeL+Q5YPrEbVIwdFT3RarpzvbLnx9SwLRYTy1f2dBHOlyLNxJTK9IF1RqoJexiQehT7IdH
ht3S7BDXtQgU5RHjIz4+eX9SqllJt0Igc98NeO0RJDMaZkK8e1EL/T21uPCMiAfeOvxTl3uXcdXq
WcUNw4578fptFaQxU/plkLY1yyg9vjZX9Zdu9Amv0xOZpfGWpObvcNBeDUvTQzi9rZAC2o9HSqNE
TGP+8ubg9NCjIoV9Af3LoGz7J4vDHodlrlpB9yz8A1677oOJFJ9ucRrotKUTNp3ZUF9bHfuLWM2E
tocEEG5w0qDjrKbAHyCz/5NqVItaMwy87wVf7Lfu+y+TrBjNpKu3qXoRbuEKBHDuL6i9EDBwSI4W
No0m56BsvLCcJh4BaBisnnO00FqrLXjfSCWo8Rtu8+xS9g7DVRbRXRg7bS1RkjMmy5E+blst1Yfm
tdMuf4WHBGMefTTakpU7FT2aM+xxkgTVSVyy7onT9qGPWsVKgP3A5MH0fMjLtXxiccGKU81OS3bD
6rX8H3q3ZPR0xEYxGH7USv8rjgLQkO2qbWyLKahAJehuKYc6BDigOYwm7WiIqnU0xkAgFpCpjhIv
Muak9YkMVSoPDjFbvPyYGF/eGtGhZuz+C5EA/CzYc/ajcJdKbKwO7jIG7/eppUtrBrCElDUAS/Vc
GE80xq/ijhZiEuWHYTncQBdspNcHDW0d5F94Pli/rQDH06ozX5wXVVpFu9XTtbu1JKjdgmqrz9AV
svLxifeREh3zhx1kP3qE8QDTviYKK7ykHJ6xxtro4lE1kNjozf5S5xCvG7GrH/imjgwfR+RBFm8x
8sFBU0SbAABdSUIHY36W4BjNCakZjrYqCmn9hsDIcSz7VMwwxCabup28OP7jMtAF+s8S6dAhqji7
fXbFpx+w5lD4n4aEMI3vfSvfwFbm8fy30989SUqI2dmKZ4A457s5xdkLyGv+Rc/WIywsrc12xE4a
hNvz2zF1ksS0oTmOCU/EI1MfRkLHpzyTwBVeggCuL26IumaIlVSmSesP2Ab2iE5C3BhHZ9LoI9G4
HaD/sIwS5hfjDpycA/9Qztn/c0h9C2FA6wptCHMCAaotNhbXAeLyD+5TekLt/4WLhNs4UrjwZzJm
U+FDjnLww50u1fskMhZOGXKtpeQYYGVEa3ftK/41M9IC44Zx02MLmDc/KokoY+97d2J7pawFphe7
rj1MRxv0Gbo1nSViCmLQlQ0oPhf1CZGaVPASjQJqAqho6DwWYEu5SvaVwBQUohFwGzLXMIlSFeb+
UZonLtOzf7eKqqfGuEUgUpqPkvyaFU4tCxkSnzCpBlmsIYAclOUWBT6j0moMVwihZmtoHjwiNNgj
td9Uxb+gUYv9Fm0oAOo6eGmmsp4DDA0/4pyDujQIBa2PQK35EPckl4uBSAuPiw0hJQK/N40gJ9sk
Xb97pqF1jMo2SwVaHPq7blFk2FvJk62RAj0HIe8776iMAK/DOSxbohrdPjz/H5kmna/OqyVYOCXZ
DCgfeK2Z/Z2zmPtBrayd6z7gr59xs3/C10HAJT3mS3zqDrVGhiDd48LqCjSfP2l6JV2bJea/BakU
gzbmVeOlUtQCVZOYHVbdc4tBf349ywQVcXIQSlPHj+K3KW5gHHwYTr5LY2VtrKJ7UhPscNyL8O4K
1CEQ6Oq8dfJf/4EBW/CYg1jTd4mc/jllT6huTLeKPmLpIcjeCFgh2jWsGPMJAP0F4kOB/TYLqt4q
L/2JiHq+v4oW//XceV7lZkASFJ4qHD270B6z9DhmZwn6B5UMy+ofxrF/9TPgg97zYWAlBwqRL8GB
0yjYVIhVc+FPshkLWPZ0VLO1KALTcDHBlKSYNDTiKV2IOcLdRhtNy82ldoHeFbTTA4ZRMbsTzsHj
CloKLy9+PgzcQTQC487EjRXbrfGFbRyDq9o5ef7o3k1M1kxeXd9j5yPjVUz2zMnGoMzoWPQDVIJk
HXriANF8UH9XJJlJNmDqFFYzvL3YvsTWz1/mBt18hbWqhOlhQx7nNLspDKrB+4/pafKpp1ynzI/v
HJJqsSGxQpeoSrzrYqSlYij/VRFtPt6hJP9jlIMOmGqbqx47uCUVI7RHxrdeJpSnghyoQGRmB4LB
i7CEkS58aubq7O3j6bdBnjh65L3cQoqBvjvM2PeOwAU7pqtoqUr/q7dMjMvfdW9WkQJxdUoTew6Z
4Cie7UzuLBnRafeZlc45Bk9HPG8w+0fy7KgmjWC/HrAzwGyr2g16CWBOqrCo1dcHLCgj0ZilQ1Q8
Tghx8R9+FHLpZpk3JAPLHTQPWzKtrkYqxv3aZug3+yqmOZQGHwg/2bBJJN+E5VghsVg92Vd/7iiE
LjikOo7wCPPTTi/xzsX1otlBdU9NNVl8OIsS3an64Ov/KGdmEQCVrgMoxP2dhfCgGZ7EHiKJfL+3
SxhXii7GgP9dzTpwIv5YUCFtBiU+YEakjgMxT+moDtxIF65wNeiCcD2f8NaLWcldVSaYeB5/ArwS
fFA4umm8NnKDahcb+Q+nrqWVPyY6/+4V2logwKSou+yrUmgSe96uG7ommNzVRWpxEdBeanjTyc04
ZNhZMrNS3ytAUDQjER/d42iYi5KWJriaR2t+Om/DX1AwT6IJz1w7gEHaUqI0dMr0Arw0STOAx0Uc
cJJOd1RzN+aErKXQni0Hz+xIsYkcEGQ1Za16nAHxHQuvQn7sC9YI1iqtrw4qrpslhPy+vj1UCRUX
vwAIcbMv3XtAH5KpSVt55ucEl2x7a41VyKUAp3wCs3DeI5b5LPl7d8XALVFgSNwrPEvkn4R3kryn
VD+tk1/XpOOvITd9akGyD9glhGMfbsBeElL37J5sCX3HFvtLZKUsgHMVXMc6gnZzW91BWhg/cHxo
e8jhGg25b5F/fANvr1g4LWBEjyxWBcZOcGnZibTzbXuDffxXcSKnAndVCGsu0cuS7KWT2/W6lwjG
u1AusrS8bPCWh5DDOdhyAQbIrxt6b6U+IZ2fLhoExMNn8gXSrIH59LEXQt4zPGS8rx2PsAPNRSw7
AnYeLHPm9VdgEpL3I9MIA00ivtnHA1iVJnNkB4ESzwE7YqkjPheP2/ihRnEzHMlOdQUWS1ac6S4p
n5tGWTfhzFtYPQyv92FragKw0dQDTKLH5tDIdvRJLcQKfd/KInbXKywbLTv6MMger2BDzosAg+bi
pmOJLr3NBMAxn0x1A6mDrsMPCPVdppJg1uRH91RMw5427YZB9BCXIlF648rbn/qfKBWZfGVT+1YY
whHfJHAe5Z1fyoCLPPepOH+LlmF9ik5alW2ab40ygaV9xNmh9x8NHzRghFOSoxYfkJZbIfJkud07
KnGDvywoDDQ64I70yedrQs2PYwXb8zec/FVuqJqdAo6PrPE3MA8ir4c7g29vCBtPHbjhRhHWaKnC
XhmNHKKa95+XIWmWRXsvBVr3z6mvD8RGjdW6fSi/wuxppaQagrgJxYRWqpEWGlp8olpb/SJYtPmt
3vPUtI2hGUZIt4c9lfvFjb8QZAl1np7/Xew8X9MfA1EnmSh59VgfgqquE6MbcBd57kosNTLhmmMo
FF93/21XC7AtyGClFWJTTeDsC3xEE9YEIwpf/b+3MOgC0HlpXG2uQOvrv8U9/ZEdzXPPS3aMNeIX
KHxPG5j+/cUrNBUmpDwKQ6dKDoEi6eksUzPSx4XaWRUm5VaTLSJBDbWKKwam9CRR5CHbZV+AFZfO
G1HY3k/VeDpaaQE7P93klSfAw8HTE+9DuUw2H0ZDvIposuX0iyc8m+TMFAl8cdmUCB6JXCzEcQ9e
2Q+ZgDx8DY4qy0azgNHCUkhDX6Dvc3B/akWzxXeFrK5UQPLaiQiFjQmYDdfudonxW3g0lVI81pW6
5m2Wh/0ngQxIiX3aVqKHZJZmwty15VXqGzPiJJ8UxqZ/XJ5bfOD6ztZI/VCZM+v+PQOJxqUHiCq6
HtflUpBA/YpPocppEgZhl+n7TBqO8oHcgvcfH7KnaN/iuvPz+vhiHHL4ofZOLD3VlvVG84m15wJa
dpCtS5WahWUlyjIj5CU87IPhNRACk6guJhUGe1yvhDL5Gxbys0SDSnOX1k5xZcpX6MJlbt4luvDv
ORHJZtXHCeQEfkEmnPDBbM5S9iznbdnMew3P7RAoiQ6PsIUPCjQHaUqBAxv+RZ5J57aB+cElCZuq
hPhIp1Uhu/FvTlTOtxC74WEqzGU+v9p22JiBVH6HnFcGs27rdVJH3ryhE1KAyEnQzxPfoLSDkbiK
RWjAO3N1ut8jD7aDnz75MNC6iOeXJzk9qsDpC56Fckz7QLyT9S/wUfJwSVx4XPW9o1kVxWAhnXKT
wzLPzLJ0m/7zAikC5Fwp9uiyIEVFpT3N3KTrmVjNIQKUwD5QzaVPHN9z/Ns249Hh4xlV3OTe5yor
OdJTwO0VvR/V84kbSQmiW0HAHxfkTp3wu29lMFd6yyU4OJ7EHnOluMPnI9kbaGVgRO/aLishZzm4
slqKRoiKdy2Ig2YTVb665KBonIK3O3ERYATHR09d/HR7qp0ONRdqlUoQtzTVPYsjAXeLt+IjsVpp
aX4MbihqqVvM0Vewwa85fqgTmrQpiwKR/74ZRKkxJ3sfwMz9qMeMy9oILGmaVevkq12X3iV0A2oz
sRz7ECG2OJTMLOL2h+ildNKt66I9zwfndvsNNfKefVuV5SbCVeXigu1OcBQHfyeVOjC79y2iyifK
DVE3qPso9yGjALej5SqCqGP4AIh6y77FkhwHLP83jd2RF2nqmQqlWWHF5GTewx/OPQTwrbvoZOEf
wk5upSvEub92SLtc9O8WWw/axo8kklOXAcwa/shewSRmr33yxYtgKgZ/B2AoxfXw8Itte7R6CSAM
TjcCr8RDrW0kS8MjRLMH4Yp4V8TbmYrxdx7kpBHPI9Rqq7cebPbLX7gI7bX4CHn2lB5hjeQ4lvOw
9EPNENyUzHNuz21qNlAE7xErcJ2zDKiBAjwOqBBC4zTrwuQ+6FXo1BM3Qgg0jCSTAhGdOLZru4jv
dtTHMtbllfy0MU2lb1HroiE48EpSRIwn+mjgmAEMjOBCPCLiWO+jdmH1bxUipGIQ2RtwW/X18b/c
fa2t5e07rXDL/q1ENwwaNXaJ17SEd8tuJ4H35LWg+4f+icyi0xiRQpKK8QRZa/iSPX4nSO/e3G27
qb/SN+rR7iw4f1TrKPaAJLm40c8l0Ug1cCoOyXhRB1+KPBdA9LymL0/2sSGDy0ajPBAtBhNHuPdV
R+hMm+M9Y5LZkq8FkgeOK3bG7NQIOvRJiCtihY1IYs5yMEeId4N2vEL+CxZrEGkTqUb6d6TW/3UJ
xTbdfHiLHAGzGYe6jSC98wq46+R2xQfc7z/TvjmqaQXXzBu93LFOkis6BeF+OnvkRQYXW02pBOdk
iNFpGdjhZvxC1ibSkzBQjebcX1R1E4Rm+Kl8K7WNQbgPI03abOgHdUlxoc+YV0ig17jWVLd0KNcx
w7/hN11APgmX/aIU2tSTUvUByTUFpqhaw+p+0SYg2caSFmNRnwLEgbtf3bB806q0oFdMEw7JzkOS
zs06324qy3sfocYawUfiEqDPizsZjc3aAAZfa04Tynma755L0h9wYDv57lS6dHTjdgqfbOJhl9jS
XPJe6S9SXPvJSXscYxyAXlUofeqidVIO5GLmKMh7KDdRBgraoHlqnGnkZ6yf27THveqf2++Yixk6
47mfymOA1N9aTZ6yEL36gHWfaNt/f4fEEJsF/LOe7bM8eAOdu3HXfo251YV7N6CC1sgB1q5PTygW
6nvVay5AubQYCU7LU+Y4DOqvc0tHdT7in8yrUfTJ/nDlcIpWxoj6Nnsy/08lM7/4LPtO/q40g/gR
ScJ4+HHI7cZN7q2zIjqQUxytwucUBxYDSH6OErTdj0AetDKxA/6GeC2BbWJNSrrJEQGCvCg0C8l2
H+RB0s8c6MVpvVGxr/Ak3m+EpVioZXSWZ1yzTYrlOet2GK5jWq8VPz5doFd4Bc80fy9wYZVSV1dJ
AOrk4vW/wgzEDwdKhFSfakkltGQ38w8ruuUs5wD+25ITsbr4zzyGQmWEaX8cEHa5JbVU6Bk3VTMh
iQ6CLlDaFiVX/ffHCt1Ux7ZO8i4ZAPhzEgOj5tYWvJrdlUhrJkZGtD5RUwzpUNySo+H9KAP8zaS8
6VWxfGPfNKICRBhgSnsBAhCaBruXMwlmLj/uUvpTnDgckDZyGdgPuAMvyrZp82RUXtgOVPTjnddV
UBZT2avOimyw4OJbdgThx6YBwk5WGkx9hTWXF3tsRFPeCwk+fGTqBSsQPGOoZZaAPaaKPIWwik0O
w4UyQgKl9HBYY4rmkjp8wYUugcO+imai5t2vLOBLku2wp4o0l7MpexRF9CvYqQYcMgCLieifRGWm
qMt3FxGrWGDDDok5HGEEHOaaCDRbme9RViwrAxXr3SH0ron8Zw2yKV/pNACULisBFhl1W1ZQgnVd
e/UibtRf9KVRHaWmkyRcBJi3CErtWqicTfXcwJsHw2B5F+250uKG8Onlab+A2ZAlkGdttefc17Qq
OdQKsFRwM4sjOBLcuj5nNyo/6h8LwTy1bstRyNSRrorHRA7z/Y7QJj/WOpnt9ZzrAAS7Km4Zu/E2
fyKgyzpXCYQGngD7zsG1bMxivzJSeqRdGDnXMd5uS4yBNdifAdQuq1VrWBzpNLW2+vT5NJYuDiEu
M/zFnaJNbjZ+7zKFqJrmLyz7SyQlJC5yNcdgOftSvwuNH05n6cLJh/D5mAD88IWvv1neUOF9Lz7C
47yNuVxnhVFw2A/FMA5X2vBS5ykmwUyo3bjFx1COwMxFtIF+SL1+scOYlXIXJGEIlxSy7Bh1glLJ
ZjlWUMaINXXQ9KlevXWWfDCrLUVhgWk/cuTrOL6G5YUGPnPR3ezo4Bz2LmwrhyJ5WorjKPRbd/6T
GRSRojCh9domoX7ds2C30WdFlCfXINsX1vQsjolHYDk+iRNVb79cXUsDFDqrZPe4rbbM9UpOAfSE
h3j0X7qtKpp9Pf5KmLujcUdLMo5b5RCIe4uJnFRRce+To40E4DZMO84psu45SifOyA1gNRsan/Uu
gIvi+CFpeMSiqGdV8zVHzBZbd38rwglHSDmK9WIPIW0BUdOmZGyAJWW4yqSyN5I7/RDrIKFCcqrh
weWWa5d+puQg4x9C/+aoNJs7QihKZKqPuMRJ4Q7cGnolbAX3Jv697TU1VzJ76uT434ZXLr3cXhn7
D8F5O9+zastCjJUhA7bVrieQGLJx01fluoDujB0a7mqZl/sUOG9xra1qCvvNxNXa5tGPMU9uKgR/
etuyJcmrVkALZqhIOd4DWjJKRDEAwAmd7DUJJaWprH7iwhpOwLowdGncLgU9lsltEdzPIFQtS0VT
DWXBqQ15x5ZQrmR4SDZCXN9+md5AB7nbTaQyUBqdrjNa3TvrB0vpEvqi5nVT+aeXo0ghL9wwpbuL
RCGpjNu/TxLF6zwJdrH7UTozHyEBFPXqQ92z/DeTHKi4mT0knP5mn9djj2YCMCT8SkqXQpNGkUaP
hbYVXjS4IwQCAeXTpoM3gpDEhTChLGOLSUAgKItWr9UY/rOK/UQkoscr9caeeEqkAz3MYdlt8Q7Q
w5EVSE0DqgTZ+vf+kOgUkQkjaY7yqrbqVdFShU689WgAHs64V5ngl+xjStVVBlHdCSvhxjF9LtVW
pGg17YaXr1rBa9HPh93YDqKTeDcw1z/DoqlzXctIv8TtNihrY35F8iFbWAfp1eIa2egBDJKvSkl4
9303meqlgD28MHngh/5BORqG7T6ykI3k04jYHNtkZsZwJqaC4KfT4muvlMOj4i7DhNf9lU8I24e2
Bp05sl5J8HT3MXW3GJEg4I8iihulVHKJSDihE3dXRBL9WQZoYzD7bk6sPbhuHcVvZpcl4vgrZBoZ
NlkzyBMogJlpo7n0Z15PTXlAJ1Uaj1kAFgryeArpa9j3jvN6KpGIRrm6tf6S6asHVSP1TRzpBPl5
Mtm7rY6ylnRSR+sPBAleK7Ugvi4pu7T0JJv9C3AfrqT/ufdoekPK8+6FvOrhBOU1cDNJlXjx14QG
1PqqRPgGebv6FxCuBC5BRsxsRbiA09VohPBJiCvrsjIK55UfSzlKxHdyLqN/DGLh2mEghFMjxFbU
Zh7jIzSM74haMdD7DVsmoGXo9YS5Yr00reWkQ0rivk4g0a9mD5GgV+HeAJA3Rhb1Qo9eZPJPRLL+
zH5kdc/Iq2b9/mbKcM7H6rwhE4y9SGEwAgYP1YzROBeJQdXmwQnYO6IFr7RW3LwL440e6TQlRq1w
nscMwVkI3svVKUhkY48myugPOfPCs5zNHiiU43l6DuGjFhDxLvgitHxh0SO27gXGLNiBGJJArvQk
WBrn2g5+/o/NYQyLF160X7nAGLlxmM+OzxXJuj35aaojTvOc5lkOEwE/lF3NUNxk5tFNQg8+7DDs
dYXVBAxx9f0RA1Mzne9/31wajq4xu72HigvTn0vUMPZ8N5hr5E50Gsw+FKuj0OSCSFCevEYPC6f9
RAEAQ8vYJlrv5azcKZQbmOkfzobaeL0vUdRN9nyoWxOZ2nisF/Qw4DuaT5G+rzsYBU4Luz8oYWvD
Ng+uO8lGRXLHbKoL2DGDPO9YNb7Dt/DwNWnfeFtQKJdGTE68nlDNHVKv3/z2S8iIuj8CMQ/cY2v7
JAo9K5WbDMbQsvk70EMpYu2jUnUcwcvzbQNfj5ihgtt4aHb4Ri0dqm1Y/y35yfKvWL60vld4X3CI
oBdoa/fjyRqEzNfFF4of3+bsxJCikkKjVDJuU6JUW+O3pbo7hoglmHJc8ACCe0exsPAWMe9aZeWP
9C9oNSlK65U/paMYY/ouu7a+SSS0f8GtS6HdcPsUfO9bvPxmq4yh1BQI1kwgU3t9CS+fHijfmYB6
N5upotoxCl89q1ZYW4YqU8gLBCDNYNifSm49xDrRPquq4l8i2VUYm77tAbTFcWf0h5wT/qBwMHoZ
HodDvYdZKKIcN6EsMwQzIQWdEtNHkrS90ddc0y62PQRGyTFRckeaNbFMpUPEtfBb9fTGDQFTWxgx
9qx2jRR4B5CcPWyF8aiI2aYbyQW+R8WFIE5ht2mDUyoFZBgTGijhEkVSDAILuEjrbqAz8oNuq782
uWQME1N9NOi1kI8ut2pmKFzjB5BIdd2hs8bwYa/STYatqjW/Z5tAbjM4P8irU/NHvktWeRdq225Q
mZOJ3I2a9elnwYbYHbcyCkleq/V38F14OitcAHrUNPt8v9U59eYPhOh/oH4ZQwac0TPtPR8IgmTj
eFuSH9dsEcW1QGZpQo6Vbk96DjypBn5hPUyW/6AlYLpd44YXV65Mq+lZUbmV30aFWim1JaPofAkm
OdbIJT6uIoTGfUWLch/jAiPgiVDjAqvslY4gHzfEnrK3IiAV3oBTI33W4SYp++UcFFka4c3j7CkX
98SVHC5BzYW+OsCLPI/4mVKNHozgfWhfbnZATTdM8qc0FZAVYWO4WoOt+vnreNO6o8izlwHaNcsS
EvXxfZ0uchUQLdUNvEQkNMAXZTNnLzG2KrZcLwXmn0N7VLA6zdNzUF75O6dFmjq6geGfUeSA8zQg
fVXbXEKFV3IQ5VpE9HSocnowEUzsqJHqSHCQBkEtlXKZUJUU2LvgoLTyKBOQTns09W/9ixnL2Csq
H6/y8kBDf+//hzLHxbYyIhPsOqzOsDhlRfZHkzbPi1MWQ+Hphf7KEC6VnRdeZGhmoqkO2oKJt12a
Ul0n01o7XQMwbNEd2hjjLHMCeKfhbmPx8L6rMv8JdXVnsBykqSARDoyrFdQ8wiAYevmnm4CCEY3H
Sh/hP5MTx1je7cCHdCKUpAwZb1p869RGuI6oeYwbTIaVWp6rNobyy1ZWAvbo5488DUYO+GmZmb2M
x0yo/C6CwD8W8nRHDaDK0fpelo8OnXl4dEC5EsmdcP79pc3mGyYHBr2pYFAsXsJ7U2UbSq2ouzJf
2mWOpUs4TXpIzVIPCZIfS3MfXmDlvja7b0VMD9MPngUOxLFAtRjDmtEoOjVaGMRCa2jCH3COthcc
CYprgpyuhw50OKBREO1DxBZ2USSZJfGicc2w3+M4fLKTb71ay1oNvhBL9BttMHq4RQYLUPA8r7vc
8OQz9Xaua2zmFYbF7/5XHUf3/PpfpGIlo7n8t/KszzteE+WQOekN0RN+Hy43ZtD+Pef9P48I9C3+
5D4yxdKX2iO22WbX4z+zeb5VPBTyLB7p3o/CMARLCyAdB+DiSB0rKgp1mef9TO9wgJ27kEFC6QfM
Dxowi05XXY5Wp9efqBQ1MOp/CItMOm3FTCpOQMb1ZBIjyaV6WzhE5EnXdjgeW484TywbBQFChYyC
l7v+Vt5CIjdLWRVorShzuyPusE276vFIeHB9nX0vRmYPEpXT/HQlxabSJk06bt+IjPtYdabWnAGT
k7pIUHV1nRX2r+SWh3Oxp3rsuJvVnW5DrwfoLbzIfHPKvXxd4uxFokVsKCDq2jrx2f8jMqYN1uSo
uhvz9VTMIlWcFTies+C/pYqZo8L95z65A42Sg6k7aFX1hr+MwoCYXrdXulgt9MRQEvxUM+PzmwLD
Cw2ZZg+rs+uilQnuXz/maqNPbJO+J0m/LLfIalVJOJe91nmcEfq5fd/zLlakdq1IZabbtrIfiX7U
d6s9UjxvE7k7lej8G2+au7bQV9ccPpLnDM1/gZtrfy0Vkoe2iKSZgTvqlt3j/q1QNPHwXnfUMBjY
pEvwmL6Qnk+uyaUX01QC0xeKLdJ3vGpcaLHGXW9pC0/ODUjB7VcsECymGqZCXOvoe4H7Umu6k11T
m9PcAKvdE12MF9jPON0ickcQj5czWSN4D3X50E2svUwg2iUmfk4b+jEDlaxG5NO/YooIXseAGrj+
sfD0Co4Nmsb/sohEC7My+dLHZQdIYvjXe0APmE6Fxv+9h8mYVmgHHoKaHyeIXptOO93YXPf8y4Do
DF0ITjT6uVjmjGbzk2z50VNKJDAlFqp7Egyvsa9uEAxUVzs4YYn3JXnbFtQlk4J0ATxmpQh1vAMb
uHwOBU11j1Wy0craW2jBa+TNRJNwijHTyEwxTAkV+K+aFZJI1LkslieYRBcUv5W68mBxirOfIt4p
aepUYYljq2PHa20m6s7I5mulgfRdenyxsUd4bkt6WZG3zl65TEyKc2Q+3n9ifgV+UuCJvMkQf78p
KGdDzDK/u9S5US283yJ0leXBFAhPO8UM4+BilK7WJcm/uuVfpzFRDW5Bdw6XTh5nJtlmqIJRH7Wi
vOaq/ew8K0gWBcHwFMCgRugGXn16YU+Qth64+jGl21QETXUYybh6w2fdzU6pWQ4uaMlFNeIQa1On
PvBIYm4Pp6oh72J1Dhjt4EnclXQW+MybMGUffWizrOw9U2GtAesslfAqgBALwKhYCvgyPeT/RPE+
Lnxu+J4NDp99cIjVYAfx6v4qnnDZDJcLV44lmSIH7mAu8n43jhN2bVqQpX1E3vIRZvREndPaJy8R
HXK/JzwXepSUTeqnWp+lHPwe7XhfGvBpuDMdSkR7SOiXDaWG+LANIYXQwmjYvur6AEry+7t3PT4j
DWhcNzdifolTcjCufqARv7lBMC6FIjVOyYYxkSWBoLYzaRIT/9th+yRt+I7QXmQUGXRBlTokycYU
bpFf8K01qU0/GsdmLLGWk2b47t2eanorxInvhNXrmwviojChgy/1q8hSFI5d5Yp60WiydsuFNAL6
go91RLy6EMytIZ6t8sxkRnmOp+ZWoTqxvnzJXFVMIf+zpmIetNsrbQFxjxPXHBPEeIjrFsGI1YAr
qPiHEcXx4IE4P5DsYeSEvxp49M2M7BnuSbcxXtNmZd+OMmMHLUK7VTh6F1mLpzfIiE6dEAiAJAXp
W6MhmZch5BKIlt17X81eg6l972sUSPLNjHaS82AGmaaz3z4n3FbvQbEJk9PlgWnYCnbwXrtwHbSB
381mwDKeS8LTY4x12F27XCUegCA/eq+kWixsiGhMTF6ZKRfIPEAAQDPChlo21hucOeOKhA7MNg86
sfF9NDzOorlPG7Y8jUjLDkFys69KyTGc4MK5v2UvXmuPcGBn7pKN+nqeevqEh5lZIpZSBu3CauD4
2gnlni06pBVqVU8gwaOmQb4FR4c9jCJxn0EBgavnWAdmgBaoe480KLKf/YYCVIuLcBEM/j96Gi0H
vLh4vSXZw9niL9VVjBqlp7OKI3VQy+NpufqJoI9gjahaTxFlSXRbHu5i6jpvOZY5kJMrrHUaQZ4m
45bx5h5XEd/daCNAbqk1lYlaJyTsH1gIUBX+DusWza+fSCiNobGMIvjH9ouT3xilrezpnLSu231V
WOljgurb7Izm464iLJioYEwcF03aD5bQZM4O/O1dTwk8sDXFjrUul2cRDhiQg0JDqrowvyQx28pj
ORib8Le8BWIUrcmXylja+OGdjAQeAfAQRvbs31+XH7+s9ADksk/IGaTqPOQJqvztcsGIVEhLQU60
g5KwK/vhnXp/m1MWgCN+YfYVfmbBLVvYuyrwtD3vOGmOju7YhdeVg0rj2ln+7G/vUhkH2Xgllypi
pTa0ygyk6istXwuKF/X9dQSQgiJIUhJAj5inFw8+yDPRR5vSsGJ398LFp8Dnt/T2O2rbl5TNc446
RoaY45VnOP7C6Vl35+8HUjPzlRXGcNJ4qIsOHKpDLKLWA1JQgn3sUZnTa78xguIZ4GQ9OnWxg7cy
kYZWzUZypVxe0DUui+eIdiYDHIg/eGe01pUvoj3FaCL7KcrXnbmOsz4cepvrxa8QkVWBzA8KEor2
qp8UivkmZoUFH+wg7uxqTJSbe6CQwOx0KE4JUmfUyLEuME7YbULp7hJNTMhe4AI0Wjoz2UTv+Cdi
vjqF1uj/3OxQXooQHxSfJNtPSwQomc8Odv4NdHCX+TgfWdmy1rQ2PNV3kau9gesCCyPyZhHo5Nrc
vPkbc3lm8pUNJEoexTBB8iXRN5HQ7vVu9OZ/Jo00dBN9haQRIdQs33VR4BZ91fiFlW2+yWx6Rq7J
cY5O3QiifJEv8y4Owo2+wDa830DeI6SuIU4FUpYldSviy82TuR9pi8GL+C+q9bsc2IlHGRKpkbXA
DshvnsWZ85nFkMkH7YoKv0urPUx+MWMirGBIn9pSlP/sk9LHwv7ei+yAOIpvEQl9vlnvfCnUMBe2
iWXDYHvzy26pPpY1S+5IALlTmLBAli/P3To9c0k0cQiNBIQwW4t5zMczud37gXX/GptN2jRCyGgV
8m/OcfkA2sbSmqNEj1HyaTc9l4dpxm7gAvFgkZFXa2NUqgcXrIYPU/2EKlEQkaQbGYG3gNtvcNKY
YxHHHGtIR0L2bYAULLQdHnvD/AYb5KK3OhzdfIJlBk6gW0LR0vDNCj6UnguXymGQfpipuvzMEfoA
Zxiwk1HufIY7dOY8DNUgFzVU1tozziwUoltupWRe9+RyQXRWc8a2cUFNTuXqkQyTIP6I0ISIFuqu
vtSx4f9kAomklMIeBhl2n+steYMx6JY8UZiYPyDoSaFeJFytJfycH+9VW1W3NlW22agGOquzChq0
pFK7du5UTlT1h2NL72zxsRiPFwbW4f1FO4LQ8ZzzMiEhPJgPMGt3XEODXoIpEBSqPnvDOBrSPKqU
uQ38zlt5C70rpX2l5b6i30p/8In2RG9rA0XeL3rGU4zzLP3tfSEDrrXFEZTG8d83scCWsRGnAx9g
KfzIbu80oqWeHgFHHzQ1w8fzwEAKadgkSKVnE/EYLNaUyYTJdSApiLaxKWZlVpyaNEblqyfcWjRU
w6pSxfLIIMDxIDEAf4/eQk8Q/8h7Puz5Z9sp3BoSJUzNo04NTcds2woNpi/9nyrGdmJN5+SDvtr5
vGAvz7w6R/vLgbljzj2YTPIcBRuGrG6ieuDK4Dw5h+VeizNtZnBplQPI/JGe8wXcvsZHkP/BLvwt
i/1lK2A1+VxRLRwNvYAwJkcJaM2tb+j2p7IIpEjPWaYE5RQ2CX0MzxNCfelgTuUT4An2vPNGcjyO
C/wXPhwiPepUGidCzbGC5SD7C5S+RTCRwvJSXDiINPcSyPfFy/tJcshSk5uZ5Tf1f12imVThYUkz
rx5SLycFyy/24tP4z9tM38xxGw4Vv+Fhmhlpj6BIKrPZ8hoyDD/2wRLsKGmqOzR1gi3GWZhq3r0a
72gvIEYIul3dwjfvO+V4vWChhvDO7I8uvReux7jXDOtlnMFbs8nGr6f1Ih5J8/40CJd7IwEOeGZa
qxOy+qoSzU8Kn4F9kJaqFiGXTSyzKKF3lR2cIj8+VQkUZBSIpfI1CwMWRfj9K9e1Vht2CfL/x0RW
mLrVnJQNSrcACwTEvZURne4ZnMZP5h+I6dBZ0nKWmg0Bd6vbijT62Nl0riyHfkZX67hFI17zF8/B
kWCNJHnWYII7NEmr4MSPRDp9qLT7eUx5SAfp+Y90W24FpzDh3V6850HZFQAVKwFnwsVbHQDMzh8K
ZdHJDT1oYOkJSiRSjZvW1TKA3JXudKQ9jCDGnwcnyp30fv5jcxYSJpddax3iSf/WaM5O01bDLHup
6qv9mNkArubLLjYfRb8fyX4O22t8wU3COYLrZjkYS+5FWVTV2S8b3Igq0hMGyQJTvUmmua/tDwXZ
22vrIqg4cO3ppVSzluu3i5PVCqTWduMAWiQHY7OmYQ+NEvi5jKW711yAt//3iW29JcNogykv+cfa
g2RxBLtE6JqpPpK55bHiX2ue5TWbYcARHo4uot38XlgeZ1j0UW5aCiEljE9gg+SMDTAT1IEwNUWE
eMloC9/4m0hSZvsowtP5iaYGFQqXJ9rO45yNcuCIS4B611NztJl4oyTVUIgniHaL/2P9AFSmzaVU
TztROdldqlhTD5pbDzhyMEF22RC9Z1EiXldCW1bgSp+8VA0BDAAoV597/Nxv/arPlmHY4NcOivV7
+A/ZKLkmygRw+YXdD+8rQtf/mPoAzhZ2DKtz1C2az+9j3XUKR6iXBBuNzTPxaQO0SQbQGj4VAF5V
FUWoH0+cIB9/rf4ju89DzgTGUFOcZDJAHeXqJZzAyrJV4ZApF2L6b1G7nS8UzaQWf/f+KAvSfGcM
H0gL/VyhIgNTNefz1diHQ8TJQb+E8jNedJnMreibGF4fuXDWC7YC85k5TmplUPBmQuapYhPvrzZj
4M3IRqZQHURq5TanWm1PA1lOJfoKuoI9K0l/Mi4pTgDrWOaK7GDjf22NvkPxIpWTckNEnTErDS79
L8WAAXsSj+T5Wbs7Cle6cXIW5dgKlrvl22YOte0hgne3fSZz3eGlRSInEvotv+1J84CBlNb5uqeL
dugDtyzBw2NTOPvCYgrqYzMTlUZLIONVGNZ0DKbfoXv174GrUV0DDkoonGb9gyNfJv8U8EeaMaJQ
UyMhOrDOmqFaqG2TyazpJzubtGOgKOuGpBKt1LVGAyAqbTQqi+O8DLRLMVirFiBNQktmMWgF4fzF
HIYuvZvNA0AjUGqkuScEKLDb5XFoofLOyezEMcviOWMoUUn7vOPzWGw2CjtAx4KM1UYTu+YwI6GX
iiWoOUEHYMDPeFV9c5TW5W+chJfya6heJsGdnBMqjPNNedMIWkga6U7VIheQz07pBTZLbZcfLMmn
f6lyEOhf91h8mew2+RuEzlFZG/djw+moSL4bDmAta8VIfqRV/HswB22vOAh0ZA63RCVB6+bD8TuI
pyhFDMFLYoEABgaSeRcYwqKsOWI1iCpBY+JnGfsKpv2PMMP/LdKCkj1L8qbDSG4XVF+sf72649Bn
1bMWV4g99KISBUeBP+UglpOEyDqhVya/iE4CSy6SVhV5wq9ceri4skiHJ5qbmreeiv0pPjvcga9I
b5NdI96lHSdnRMhIpcu1DMpmRJovGkmy/9NTdENH0kken5AOVOzZrTpet+e3e2dwObq3IaEe9vYp
vI0wEQ8ntlWqLlMPlrR58RnJAxR+xNbVoGm4gIZyU2uE/7M+OSyXl+/nLdM55RhaqKD6aKdbyQj1
wPr5Hm2H77Gq78BK1Izzvja19plk/2g5rmI8bvBfNnP+9cq3Pkuc3hbe/gK8GoKsMCVTzgD41icr
sHWuahXlqMuTZjYTYfWcP/28z1x+I3n258h/m0+38/1tJyRwHQ8AdGBffxAguoHyfyGDQQYTP8pq
6/FI7rtSH62tDd7OtNQ9New3CvUaVJQd/OHsji1pAgoENAGQWDp/CLOqgj1liTtOFdQsfc6+pU6J
fnGqcxQm3SPdj17yFQoAYdGZayXRtFAgYF+caUWQRVBOBa+ly+ADdHWVIX7iXBwAj+jbsiLT2D0g
4iEuVkgKXWJztt3DhC2Zd9SM5nvTsIBEKc6KmmRLhDZXVfXWNeGJlIT5rDtb6oq9GXrKf/lbMS1+
dLFgX8Bm8PajFuYIIEA+ZakYy5r23xF2Mx+OD4iZunA7rrQlGaBh/bPd3U1A5RpRfZ3atgc9mTKt
eDj0RQzmJMqexMyS/ceehuArkYaTe5mZfGTzh6PZq50JpkRV80HyQmynoPrfQ//PQ54BSNgHCM7A
xYMbh7mSf8RA5hNNHzdLKk1lmwjK42s5M8PA2sF11ly+2svSetBbzwIY7qBkTBsK2x6/08aSGUZc
vshNpE1rL4T0MXMPjr2TXIxz+vjStKT4g2VfaE5j6fFhQDMW2UnWHOaI1HXXtff5swPQ9F/AV2xu
hAxYK4aN7i9OmD4MwTULaZooHQj50HuLfZdkDpnBCPTawoWebRcLrvCF8JeRaK00qbtBtdHMe+Cs
3HAlGzYFy2WB4NJhobCzLbi99njVbsdbPdytdZRTSfHHZboI/nu+ETG3QDZs5vqS4Z9lSJxdMfcF
cLHiDZitTwnpqi0tkygngRS0Cl2zJDqCdL0cDrQ6MHdWsMHMKBB4EGi2hc5SnNmSadXXiA1nZY9o
oVx5qlgfcL75FtXLPDWOasdAhmKZIhDrGsafTSMROdKobIRTJYsYg51h0xfOP0Ip7rBQ1zgSfSnP
qppTHfy0CfN/mmI44xgrzgmLVvJrnH80fWtpoSgXM0H46F0DztFtQYTL38ZQCyjhuX8sdAHUbKon
Rh2cobPgCEIGV5MjMRR7kFFv91J6v41HngsZYOEIwIxydqMtwZgpQztLCmAzYPLkTRJiSQa+g+FY
jPRg4oRanw2AlTUY3qr+HrW9MLS7vZpTsVUyucp9l2igiMZwNJMPv9El7o1zAdSsE4v9XWzgHd/h
dV88qQXwTXlKM8KLC73oWOqSdrWBrGAU20u6Pp06QIhVyw+ENYuDLh6p+NPGzh2bebw76kXEXXpo
hAVRL1OpU59o0artmq8h2RxK8W6f1v4BE4a11dBK5VErStctYOLyP34EmGi+3iKiNSRhLtVRXdnz
uf0BKuUFPEx7qulHiRtPGQdvzYy+NRrIetAPY3V6rluXMf7TVQ6rAaeSen51LYhETOaRyo3D0mj/
tuf4E7HUIytntmGJ5Z/wqLkYHL6d2p21X8ztJXqJz0meJhllkGgNQ5h+xjuLhqIQkGNmi/Oa1DMf
mDTPY9eyR3Lx0H2lz5+UV/F/Vno9/0UA4t+SFKzaGCJBVmfnXfRVtwAVk/nTRgkaorHiMgKf6PWD
uJEotcvejXCKLjunlLssqddlngYUzkyyNSmJz6nUMaZV0AeftzqjZxprduW94v3+UPGmZY+kg/Bf
CRmYlAf21S6MxRHq+iYU9AZrr5K/CF8PsR9Wg2hu/QPnX+FhIlSNFXCDE8aHVOMNhUX9vN0FNRbF
GyLvI3LLM/NtAqzLhIW/51z3MWnFqmbD12SUGW16onoH5zfZtLlC/sny20/kjFKc3/EFnUSrBkBQ
9J7PriBTkEfL54N1tVQVaPdRxtoHwC2o9EyCyBOeO9hrckkVcD6pAvS/LOONEPlbp0pB1IKsoFPY
mUwRCgvHa2PjPSJ7SEPNHkAsEF5FQqFyya/S7cUJg5ER929yAXZNkWFuNXlvxQjvCTde7Cw/gEbI
DJTGWfEC62I4ZwZbWzssqSKi+PZQ0QSHeZE7mb5XyoHPtD9kxHMfaBcnY8HnwLRTfQBwV8dpHGu1
Ak9W1JnkqgmA+qv/30vV6KAsv2dvaJmM/3CJ/Ln7ImOfOrMFt4hxWBlcTjqAnDkd1Baon4w9q+VK
fFXxEdI0nWwXTCL3D9P3FFB81BUUSqPgrEl6cNQhZd+ZIWFhkBveJ7LRShfVNncf0vCC6CmMtu1A
uQza3PLU1RRGcAKEPPzYrQJv+dN7ZRft9HYfPQDf3tvAqD+vLKKXBP6fzDzpVcRM6SEAQk9Ifhmm
4c2DRjq5C0Sb7wBjRmUufJLG677zag7J6mHAQlUop/pHM5Y6AeE//robs+pLLVkLO2mtn04Rccl2
CRDOT1cSaqPeBYLxMu+7a11D4th+u4UJK0uBLX1BhZObDEFceC8FAAT8uM6o4A1zO81FVderOCJi
oFsCwu/4ltwFyTPO1oq0lU8ZzuRIxWAr3qYVOb8bfUu+xhTzYJ9xnWKmYd2Pu6dE+qqbhkJ+2Vzl
5ICwaV28o7WqeVmHgmeUjMzBEDGMkZ2rp+2s9Sf+nAB1jK4aRFf9Yg9Lfe4eo7W23K/bypib6HcX
zKs0XpY8EJc71IjlBHFSsnd643orXBwMuSXNR3Ej7NoxrQDSta+2uFnE+edTvaWzx7BUqfIs06oL
bz2lB48f5ZgKMtZG+y4boz3wcZL8RgmXaEIB+l5E13T0toTlqCW5LTlKMraht8P+6KUuHKtRtEiZ
Dj0UNzgOHFk5AhjLK9kOUspoJWZBLFkj34vS044KmerSBzTx0+OimrtUEXhiUrxZbWLyCIoMHgmu
ohgTryoSh7pyRAP0sEzESXJB+io6Zl0ECXrpwQg6/6s4STbCg44PmK2GXyaNRChwCimHUdHeonql
fz13JQHPkPbYI/JeM0QZ2po+hjeoenNfdcFnCYHiMLNWfvS/WWOekOTj7rm7sHXHS0s7iU1MY51i
1DwdudWK9dmGVV7Sb3ukJ6+WX/Y5yPziwr0s/xil4IFBcvDOeEyIE+wB/aVRZgXvIqaQfiyfmJXz
jzGSthsumrxtv1cqrCzSNtuRiKrHRrppISI0dCCI7ZCvwM9dWmbwFl1L3VuCVrHiS259V0hk/lKU
ugCwxuDkycbQuCC9fqrLzqUsffkTpzKy7zK8t9z5YK9d/tZ9KsvhPVIiTQ1I4cskNptmoa1u7CZS
xPQTlqhatuT9mR8RAo5tEoEQlJnK9znDKohw94CBuSzw1vkv9YtQeRt0M211asK8oApIe5LfrCKg
BTrI1r4+XI3in+3hKQY5mioT4z65d90GqgcVVOR/qpILll8U2Z0TryboKqdbhV+pbzuAl1Vu5ARC
cOjnjx18nSdcdGP44sJgsvG09Iz3t6mViJiiezcS49/4EzCFJDexUKe7uFNPu3IVZML0Avn13aGj
g7rxDrFCRpaPNfrr4YYGZ2mVUvhaQ/nGogosw4Qn/+xRaEcrTGdMEJx5Jjx3qNA6dSC/TWOXS79H
/TblU6f14DPgUoadgbXE6ULkqDOhwOQhZRvFvHy722ZKcCh6Y5xX7lsTsaNkZOVj7nfPtCfNjaMs
vax57ivPVaVtMusd8hdWmbDKyJOFBFcAxAuu2wAFG4Q8r2qZLnwQFTImUP5/TAoIJwdeKj/5CxnW
M5FgjqBukpFzO70PF7lIhZHWYNaK4t7YFhpwoRMIZUHW4V9nCN2H0cSntd4rQnGZfPsYio8FZRSP
nVsEJfl7Z2ljFtbBufV/aZt7TB298VoApA11tI76CDPT7EzXH4IVyFF+2MQlq3XqB+wYtxkDehQ/
a678xq0Tu5MY2dPHf7r3IipDdbrCloL6PWaX7cl0sWRnllSlYHaXWoeJVMVl44ChfqrlD4vWL/Sv
DBuhiHCPjtvgD0x/x+M9QFT1HBe+a3wdvgSUqM654k2XxUKUw3fxUOQSQRLUt3Ebp31RqAyKD3Qm
frmbeNXgJ40TxMRBPHyAv9a3Zbt4v2nIEVIRzzXupUvIrgcrmX8qkOTJHquhukEk0zEhutQtWvM3
e+52SyghnTpIEt+tmkQlPRPw7ip2DbDqFWsfclT4A4hJhJ6UYSOI7IM0rg/H0XOlL2DATzSggyIs
PuMuqdJy32aqE0qEwimmZMWMuIGFIDkHditvVzLRxYIC6IHfknpgupuhFlIJv6xUckIN/4uW6mtx
XXuH43QvhXxyoJrvmOttgr+3W/mct8hJ3LfhuadR1aiEXQRgNlENtO3nVY6fjMryPPFWba96DmBv
SPTpfrh8rsQetW1gofK8h3qViKlOhwlK2Q2noV1h51zTBKObHpfioiT9RWHXUbBpkU6dgma0t5mU
kE0XJRs4pAeh8Nee8+qP1thHSPJa/e1BSallYEgxV3R+ims6MPoJe8xMZaCVGkrzQ5uGfk8uK9yH
UajNRAm8RtWz4vIR7cfyxjb/8UchHavWk+tLO54JiL0zeI5lHNbW0uL9O2Q1fqo8Mm7aAUBg66hx
epapv4Xekn4NBX/wYayYFKI9+0K2bDpX+2Dl+VN+sSagy3EQgK/agZLhUlkioG9rjAemmNtF2Y2l
hUiWML/4FomRqryzPNf1xqMEoIm1MbOr5JRNBUlCJnjUn/GEvZqwIMl6EO000VUjeOnvsL4HOSDU
x3MmexSOl6UOh+Qr18IxpBWkwLKVPqL90H7y+UyAIZBPn7cC6VCAs9xl2prk9el8C7b7fHDunmr5
Ba9kW8y+/2AZmW4T+JSzj9kE4xHZQwgM1LKRqhiM3ATFe44f5N2SDbZQplL94MUrav8SPVEtd8I2
tbcLdZQJDxjKnVtQegLjbosgt7DbYykvQa57VJx8GLdQHv6kpyAcJJ2FMGyGd9wpu44ydgn5reSu
d041YGB+nBgUQK0fPLtsD1e1EyAKj2Tik+z7zuJaaUaesvXf7o5XssU3LxfdFunSIWd+cC5NrQYS
ttGV9qfJPGISL8BlyrHJ4gVPXeaWeZNjSs2Ni/suGxdIFu0r3+p+Cnhm71uqguN6HTcjwpVbMt9u
fsozUlOxNgrso6lfR4NKUJiJOw9sYGgAv3xZxd5S9bkTu7hOtT3t7VSQcV/RU/vM3ecKx75BTZIU
6Ivo8ZpITelKKd6svNM5hdMvh16OmP9laGqAiW4LfP61KgYei+lsdjm8f7VUwVHU91ZCpPv7C1Do
J6t7J4Dtrnv9AMUJSAwI0/34PGZOqFvfJ/S/62NzqJ3TFCE33111BuOAIBCpNngzy8oExZBnqIMG
kcP+AZ8/8IHixIsL/XlVVA7vO0snVGGNFPlwxsboGJtuUq4zhkcxwExFt26dA3BLN/zTcgWGGE3d
S4zlVTz87jpsUPT9jFMGKxoacsZQtAzwabMavww8ZfJpnH3qIXbQZ5E7TMmH68guwRx8iZGnOklb
zMfIbJjiTMLFpBcOwTccKMn+8hMwhp86+t3Cl5P6PR47Nbj9Yausn3I9rJVPM/8yWU3XDFFzxBSi
+HQfIsjx3q3t1C5NHU3oJr/xEKY8zfYblprp/FzW2D1kCIGfHfD28SPORqaCph2S4iw6xq/HW2lo
ldqEn8rWV0SUDJvClQTNoRIIy26MMuKSBhgoGpkxi0YzjXvK3s+KASfCBi9jvLD9lszXlXmeqw1R
B1G2LiIUrfPFGRdnEUTjRterTfTtgpeGxvcPfrVPQH5axmPjTd1QP4kcHwPPvwFR4W7QpoG9xqXl
Xfp9jnVoeLoouwzRD2KDYAwBspGOCoi8jt9S0sCtp2EV8dvsf6/OHnFjuDrmEuTsJhgDpKdt9nMV
PIfPFa55mFC458j1ZlwEbN455I1ixHthwM//8YTjq2aeWf+Hdbp9pAqbkwpM33lWI++lmDT+AZCk
+Jy/b1o864XJRKZkL1/AIQKKkfzVU6+FzbnGwUQE8+oK6A+aGJZwrYolMw7oBo/4wWL/St3CpAu0
SDQQuo9XGfHzpNOOLAy9DgoO7qeTiGfCM+vC6MOlXn8hM79vQQ/Fx4KrHW3WQ8UKG02/kmGXp8J5
RnVJPr7+T3mg/DQHkE9TWb0LahJzqtF1MUTco4h0OrN5BLkJ33P6hmm7BFLCNEU7X1/p11QwPYys
JGA9jQFFwUX22+jOTzQW7USNRWvhHS5ys7/8hpLtqUZyrUqkgbtujCA1LrpqikHcjap0riUZCyup
GwGzpHTG2FE26vReAFYSZYcBxODln1qkACIUYGVEaZfmJPD44+9aLPSzgRTqMPAhgVucNYysYUBB
IlzkfyJizasgjok2KPv/SnfdRNWnc3AkLrbVh/ekN9ikfagD5w6gTYSdx7IlxRGX2Vjwc9nRpY03
+B2n679UaZDbIILyK2+ljHxo00YvCW4TSFajr+F0QvHhj1+lwco7j5sseCKRAsooEJC/f4iipKx8
9geiP6+0aSe0RTyCyGpPchk5orjWV/LgfefcL+WpSTAOpjSP0Gb2XEnNls/oXml+zNE6rhu8sHUS
88icAPgC8W+9pC2RgyGdbznpkKocZelys5J5WAwjm7qMtcdRhIeZ7DmjrVdcdgYs1sVNGbDFaUnV
rMmrFxzs0sNcmE17gqBy2cBBhrY7iQKMjPtV33aKq6sZrnOiDY4tBw87UuqKxkwlmwn2DLRjeOt7
NS+HLXm3x7nPcH9zdkbNHgcdwxNCUOL6jMKktCTV/o/DfYFWrzD7k5T4yQJpJQRGy/quZaS8Tmyp
nyeCeqIroIaR4B/IywEpZL6nZqhnvreKwZxhQMYB2OU7YugjcXlJlkXUWwsJrdoars8V3rZrKMJd
pyDr/ZdmlaF3UE+2Xu9XxGQLzdwNIJ45EsSVZ+dbH6DjLSSb9r1fim6idkd0jPprXUTB/keDXj88
+6oRC6OPJ1Bn9K4q6CuianOR5d4rhogCgSjEpzWFunWYbequTI/xz0RvGC3xdznouHPiOspe90aC
NXqReIK8dgH15T3Wz9Uko1YNJ0ECs4nLOQRdPVYWrF+h3IdBaS/IG52H1CykBfkEobhD7tuWV1je
wrioLzO0krxkuvIP0UmBMNAkpv4q0kg7H6STocTC/8tkFjHJuJ+umzsZskf0LFWEfmO1ghT6Uc8p
9sa+rVfbN5R/HG4clcTdont1t2kJrQFlvPUVlR01/aAzEPJzVnkO6vp07b+sXJn83ftmY0xylKkP
6A47LesMYrNKTdeSJEEEsJ8mVl3Q7sWR5uVexcNc3hwSglP+xORYu26MIlYcGPYv+eRnv43VXbt5
NYN/tMJ0wKyW1hlNe7TC5xcBDckxkLgE85RKZV3V/73FA4PDkGxg3YO12K0hPg4U8RWKTvCJ1XjO
jEOUqH3OoBONYGKcqpSXUM+7KgRindAhQAEBoqD/BUYQF2RCw4/pBnprtEduiGec/5ESeLKVgz1d
HiYAyI0K6iR7KRXBjyYHDzhjnYov6lA1fkIS3m46ydwXI8NpfWUwc9jEC7LhLQz5k4gPREXejqU9
ucA1wqvd2pS+GOUhxxBf32RFqhjkWEzznR/eupzOxJHags79YPXQWCZCPqXHiwuPClMyZiX6bVIc
pzn5ppc+su3UHbClCTPN1aHWHK+sGqr/MQCUe5ORlPUsaWY6FYdvHlPeI9jb5W4us+peuc+sdzbh
yqyJ3g+Irc48zFVbP2H5VTcIUjl4sgIIjdtsmvRy570UZNeSdsGpfvqrZQoU9sRKEVQPDUG58noJ
kZbfDcJs28lmwIfAL3vQ+6p+5CYR902XYB+96Vm2kL45DdfwdtK7CPGzOzrDWTAauOQqiKEbSw23
Z+lTC0kC9g+gFgnmxGG26kZR3uRTuW6rkv0cER2YfkrZdmRNmNimuJpUrj3Ykl+shLgviV8IMQfL
xfsEd5+NzmLrYRuz1J5aKZ1MOXIWMod6IVytkenb1xoa3EQNMpJGkeRXliiWFoztaFqS8jWPf4Nt
qpkgxP9NwnlA461D4aF6hPDhNz/nAOxMEyLJVaqInl8eMfJrIevDSbyUJotep/MGS1BD5qvDYP08
Knib++WPRciYsx80GUmezbNzUrv6DquJDdE8N8m27vlGqcsicLwC7BI4/Ymh3QrSYOBHu5vVszvT
2WXRKTuGDmzMfjYE+xZscAblZBfYFdUQdN/G4hLGvRACscLsj0evDk9PgWZppeGN9TLYLA76Dkmr
jc9iQL0G1QDfnsB7K1LqnPO4Unsn+d8Zh7nZslQ4gcUVyuTZ/YX0ilZP8EubnuElnbvti1GGFlxZ
Azw9BoCU0dwWJdag+3+L3cD/dsqqfVoejLCW7WKoj8tE4Mj7U64YY9ZInvQablsa0HlgwU0Zgn//
TumZujv7ofnXCSYTCO6fyxSqmgO+YzYYsmNUNLe5eB0zZ5a2tJRU6QvbZamb4cKibP8n6j+ulAuz
7KBpl0IXCodPC41v49G5dFzUOfpbUefTEP0ljrbAdnAZoX0PFuSFVqeZ3eBIwO9Na7sel5mMs0/Z
7c8T2xyQoJgD1nzaPynT1DVgDKKHCELeMWM2QmVg/FC7QtuVMRMmT+rbsLqEeT1jqvoUGXo/2Kbc
FOClZ47pxBw+qvKDlv5uRgjIBhg22QaowLMSJD2HOcRWrZ+8IrjBe1cjIVus+sHWIOYaJqu5vMDQ
/8lIvKBN1ZiVOoli7ea6TYNfhe1S8O9FKKXeYdHHJgCc/0xHIN8j8Pi5wPJ44YmL9MrOBF9EnkHj
qY0xr3s++XvdZSuFJDvCSY21GgnllqJwSx4cCiPxy5DTZsJfYkIytQxPXVf+yqkxyd2t9gLWK7k3
sfK+v2eFWTX82u75ROnYbZPWBSQbpgttBLy+SZijOXk76MBLoHMXEI5ghchg2Y/PP4ekV5tdmwWd
aPSKCMHwHg6i1Je2SMGkNypw8QqNTabqoS96YdSXV4UURGyzzHGEEg6HGgaZErZE2Ptz+1kOkdro
ekntY7vQ7FkZPll9rfrKDLCpSqLtScxLRaBFbwIyidknRJA5J6p84MG7mB86hZ5Kam1FbIHdVMIG
Q6iSMTkg8bATM2r0bx6wR+1HUnpwzrLK6vKolM18ah2fU7HtDR1UuJ962gwtrn8VdwTH7Ld3hM1W
tJngxdCvStsDYVWOAPXUNhA3L4WZ5BSUI6P3+Jqa2Q4qxdUPWOyr4485IGP6ZweeOFdMogQwyIoZ
wAAyEfh+LO12VmxQkrAUwWmirvBTvw0ZIasGqPBtD2cP3wgTj6kkqckSLTJo01oAp5i4mUi5wcfL
z+lMWOlhIacioKqSSF8U3vamCeixmOGiFKIUCPD2Io6u604HT0a+1sKPx5YbHld2K21Yjl65E/f0
5ePg2UXo4Z6cxESnoBa/4jADcYN1cquDDn2/Ui6hA2OLUVo3D3JfEv6u2qs3/sAL5GXwNvhmT3Zy
LAX2lZssPbtpKtYimXHh0loNHjozU0zlvWwqNZOkjsWOQqb2uhJxrSf+hEFXbgrQMi3DLq/Ysics
qkGOWAXJtT9UpHBIboIkXVTSPtMIs3wZpxeEOOWjKEqWQr0k4pClHl3QRkD92D4jRloeblTmOH9E
zpXeMkSo8Id0ZHbngQ1SgEPblDWYDQsCYckxskVMk2vyIJsPBMB9Vg8Az9Wz8kgDz/0/bFuvesNo
RUC9AwtcTR6VZGMMUGLarTRSenhlVrXxT5sqeukGm2Lp3kcXWZ9dUaOcbmy+9R9TlBjxkhy6reXZ
emgXM2BJvr1WM+8eBYhXws090H6ajtvpIfR5Lu0d7o3oE8ds/WxuAjtK5MYDQBckN0cdTgXNiXr5
wYvVgFkA4meQZqSvX9osEghGo6GxQJymF5o3J8xej/QtRudO46iJnWoJpViwCTVdPpK4f0AFW9Mc
PgPpK/MoryRQQLeUqUGA6oOl0v1zo+l8IpPda5Tha1JyYm6UjjWcfXo+PIhvSiDgDZCHB5WiuJAk
fiFjBLMX/YNDHY58aNIifub+L+b/sWAW8f4lDD5EGYCnnWAIcA96PdFttxbjVxIqQRkupbXVJThE
75ARXmTpDV81Njnn+IYQlatpUOYhKHn/doPyBlaJSHTbGgqHTro/7enRRflCKGOwQ5nwNgmBoedT
zIFoRx5hLhQjqdvK1ng7MRwWE9OiwMTDkELEMBXSCQ/MAYtKiO5V4rE38GqI94QZ9LTKxqb7lNxV
5TjM1X23lYZ9RBJqVdt7kFIAFY0NMjJCS0DcoCe8CeU8lsPZxO/v1iq6h9o+SIWEpflYn5gG0yqN
MfVSiRcly2WAO8PGTJ1KI8znHzIh3HvD9Fx/ghC/WAyiInp2Wc6BL2+TrS30SbWhRd1HjVsdyi4s
ArhOq4aIq3wZNb9XyovSc1ZxqRE2mHOjEPzbjlaFTOreJmLzaJPLKJhLV34GKFhfhd0I03Cv97Cc
eUuz/apNTVq3K9I8KaBhJ0zUkHruFowi/Wutm7CHFb5VUjlFbBjY3L3CI/o5t/Qufi6//m5IPDHK
GCEOseGGWJlBNTyXXiO5W4a0zoAgW1XajtU+nUhQKWRV/Yyn5rYJ7DA7Qxu/glhV7eoFwmwcX4ob
y8YBP5cr0GE0giF6KHg2Zc41/r1rUFKi5u+RGmOjZRl/Vjp08JSresyK2MlrelRuIjZ6NZRdyOpq
d0zDl7pV1r4oTOToJ2PsE+ehsULfs83bUvSSpUrhKGiLH64RR6QL+3MCjHUQtqjL2ANaxh0bqRbL
i748zBXHU7+HNA/tEcm0pd0YBPmyaAfw8Ewa9VObKPPjI7vln9wGTDuljyZc+aSqAbfZ8aYNab19
qSuvQmBQaK7+9yih6pMYO80/3Vyi/2z6mtYwU8EpeRF8UV91/bcWuXISlshtlzoUJPnBjTgp6yjT
M+FC2CGvaH/az/mSI6Wdjctxu9b1phdSvAgHWygHdeQtfqcJ11vS9BzbSbyLSc1t26By/wQpAOk3
39wMbK5HxPxBs6YrpdFjJu6cEG705432B9UrLZes6zdl1ie8wyF9P9TpRzW1v69yStOSiLlpa2Tc
DiZ5CbCOBGF7rBJpiUiecBlrpch488WiaNrSjTLdh0iwj8Es1xtC0zKFsVyZ+EDsbzIPozyxjxwk
PmB2L5pvXOjTPUxf44hCL0YoyjcMZ73WKClgXCLE+VGcuqwbBKJvy7Nt+v7NyQpfvL1K4CpEZXk7
YVe1hLAvskLYZ2ZBDOVbLjO9F98sV1vWdzHKwpshf20YRgARTaYIVB8j/svz34kJpXuLJEu5jEgM
lkYuxgMfpTOzGbybHRhEKNSt++FMeIE4XC2B0F2pBaI7qeYsVnQCfHdFzgsxohrIdnmSXxocMhfE
RdHEMQb1uZoevTpeRZGLfnYjBnotHpk5ifciUH23nffFzRzBmG1vWzlWsqjOSQG1wMvM5PUJQt5m
p6TD3O2O4FbIWeus0bdIfaSxeqmZohiNQAuBNKPtjg2x9C9K953KSriRMMmuWnOCJcLwKYw06nfG
24sN0PL0i7YCrc7izOQy4f2gv7SixBkgkHtiHZz8NMjnEUC9g36/ZYiu/NWvBlVorlIAg1WPNPxG
815THEQHx6sK7a+dohqKFZKJB9RSrZHAPZaCD098WJMoF7pLh5X2BEL3h8JmSfpoR7tktycPNV3I
oDayWo7JxjYbGmX1trYEKkL7FPNAsilcjaEJtqEk9F6jYUWmCF8r3ilDaeuUeiM0ooCTZ9iriify
DBlRS+z3tfCflIEiE4PsDY1cLJLRgl0MUsleR1Z8pAe1U1hofdABQP+JLwMbNxrQ1poD2g6x651X
cELvwZFlytwieTXZcURTDDYdVPMKcoeoMwOEfeYf4GlQKMsOZ1938pr7WzHMtisoQvFNqA0W4Slz
aY9X5lcMjLnplvACHhR+G/jmWbjkS0AyGIe5OyeTFir6k839AIUipxRLV3woLc2ZD3UFQ5xP2CzZ
qXhvpVIQo+fOk/p4/c2O05gwL6ARzAs1/IiBUNTEUfGkMdsjvbO+UXu5VUleRtHI9pwHcyJ9x49C
GlLGwOc15Tz4St+jLWCPj8jcHn1Gn8A0u0IXxo6vnuJj3DoOBbFZ8+B5OfuxvF1URS9/YwgAdpy0
pKVyDNw/i0EvAsHjyokkiiQbpLLDVENCo+DNmwMSHwaCJ3R7j18Tu+g3hFx1PRgWzSBNH8UkLk3k
rURlryvf1e2ZNcUJKRYJXTSvER5nTijWaWztTeAvAPwXLxpicdxpZVomgEJynJd+eUVLlKP2qcak
2Zke+nI8s0InOj6S/8FWOg4WHOBMdvvyQZ3B7OdFGCW4rvQ9CKDGpb8IAySv92eM9/I2oTKRgkKu
/YF8u0WMRIbnQveUvAASGqFHRD813Xzey4puoZAg7Klox6hBnZsjmihMlkl+ynaaTtW8JIp7BcUo
XDKNAG8waqEtHxuNTDRn3q0OgnSosE95S+StjMhEMhJ1eT+bll97d1Kesw45O3WsV1K4QN8MoUkr
h5/Kt+gKnsWb/RGH/fywqrrFK8uBNZ3p7zVQ0JX/Z8ZGIqnKXN/l99Ear2fSNI/hbkiIsUFwPda/
SDaxdTqIfmDWJ2RI8VjctETQm27EN0CGvQGfYNf/Mr5SpWNLzENqFnuKSIAzjy/xCgTCBiCYtb6z
nRTxsNMU1DvH+gFvclLzGzqoLwTmj7clW9jHJ07Jwpw4zPMKtregqQPkReBCbgS2Av4GY3W3J52b
DTbaRaMSB3zHXTEllKIjLJbtjrTvJoUruq9qMDQAnCtH3HZJAMLkc7Cf+Gec4iN+IcbPd+J3QAMb
YwYe5nTffd3V7qYAe3ZkDEay/CbBE8VF+OScGBZtJTfnupSfZU/gxqLtAy7s9TYH3EV0ePsp3y9w
cWjFvGQQaf79RC0w7vSeON9cXKvbpcHOljtVifGlFNMpJdcHl/nETppZhS3neKoEOsFoDcCF0BQd
k+NQ/b9Hrh7F1/PnkD4tZX1afuvC87DxBFdMQ5nn1jHo0X/sHQt89aGt3MbWGTwHIC3lZYQYnl+G
QqQ0MVjyTDCIPhAxMK1rx9ub92Scw3m3nnqvUOZoTpiZnfob1ZirGAchsqwVWovGkjOz3eqxxZqH
rKQWCJthgzppuq25inLAyl8brmgN9NEtEZPPIhdRwsi8g6FREJZdcBX25JwcVcOY6bHJXx5pY6xS
Hnfehz7niVpC9PVIqv5Jm8ScW7R7ItSjo1Mfw2KaJPu619nEeNR4vylT5qhYxLaG7IA39R8rWvPz
YuJyWw1B+Kfslc4dNHwy49fLtMl1jymquTmm5WncqCjphVXlQq+6hlhmjWvpCtO2BQM2HEgYriHV
2tJNptqRhBqk3kcYUR1LJLZtkgeBd91cAvM/nJ1V2oFefmr7KxeQS7p1enje3ddSvmAYNkEP7Xsb
ISrF1cANIMFYEByc8ixouTZUkfRLH4ew+cGv3safbR2BSYswb6trYvAgJDFqp3OX6b5BhjV5bZHO
rZTtn7m9vaXXWMAI4C3SfquT3+wPcyme4SB87GNS8jwJ2KGO/y7sxxKspoUz/SG4RcEbg6Bt791v
9XU0MDRlVfYLBneYMTO63IqTij1OQgCu82XDt0GTouae/FK54b6hNLmg7UjWjljs7rQNF9xRe3by
KFUeWX7TMZThYB9NUQJ//474qNLfb/7QKuyPYeK4IlKcwGuts0W4L2tqEMJTaM5wn23Q+fahTrH1
GCYW8rW1PodtEGhaTfIEJLYSHTc4EOdB++8mZFHQ17QzkMJZOqUeFSLRHPNT7f0du+5IJ0Ki5Lur
0fo3y+JvWeoYefmHdKa5UuVBLqIpiXRff054tLE2RqOn4G+tipyyIGWbaGKUE8ponlZc8C8XbP+/
4u10dYp7V3Wj2qQrisGDJr7WboSHsiL4ubodb7R0cqHJo0a0gLIqFX5IuFaVw7yxBVJkLBa4dSUk
IvAGFoHsScLfRSUC8JgF4ZcGnRrp7DL9WT8ky6U8TKYiB0qEIn49Jkq/tz+PNUqWnJUEzjUYmBQ3
ZTAbehDARvBcSg9xa8b6KxSiTw6oHn1W9CuLWjvHUq8XXs08QtVXRd3IhUdvn7f+7UzjXNdRQDGo
M/TBruVwCCkSKugfe0X6qtCcmwALlpYGME2bTTYQEcfPSDeE/L6LV/6GQMYCKsxcrvR8fG/dyJfs
QiHxd2y5/BYVjo0k2JHMNWv3a6dxPu87lox4b8IiGdrOSZt4HUCWHcGTkEyNq5DwqAKLPbf5KdB4
1RfCOsHMg6+/bLGzx1L9V5NfT3Hs1e4Y3hOIppmlLKwzs/Ok0ne6ual4fJHKHV5ClArzYvINUfPd
/jfP4aWQEpTzyLYRNepavgGuQ96Wr3uBvQoix3UYQ5rWK5xVTdkN0wkKyQNFaSbOPRIu+6QoIu2w
ROlDyv8P5URarlCoJt8Nasid+DRPuRjSLoZNHkkle7KXYZy3Ia9430tILiCHEw7NhYgJlyM07kF+
dMjg6KMj8zleocuuaS56tP8Sn3d7Ew/ayQTSNQfNoKIVK+xXdVQf0euvg33Nb2A7OSdul8onTjxI
6ahId1NzTdTnvgxdHdxGwdec2Fhqe31sFINLzsPam2uOI5HohDK2akzYI4ecIzuCKn9sOrWMRte6
zlrYxBR3hgB98jWxyq6WGxVghC56CKo+Jl3aEzNbvkJav2KWZJewupqmHxOXGzWFlio6Ysq8bhB9
YHfbm+818XEfajTl8JDBk7oTeohFAvMZgh08mKTdUWu2M8dCUIM+BTh5jhaAL5I1KhA/Vi3YVa98
W4W3U/CzWDH4HVbHo3csrKSL6nGeRbdvpfHeFn5CU5yo2LJrA3OfaWez0X3gG15RX5W1DuIVYa82
iDNlfyBBy97YEfqPtyZIIcDpnyGoKqq0tm2Snk1ghtUtcOLzPALC4AUUV30gu7SDZPKiMouCA6Wb
hKac+lgdCBQpt2gXG/dEhfKV45hbC3PmUiyTkKW1dhLheOHf+F7NvFYPz7Qy7vg07hQHUrRKgthZ
2fYdSYkCXRcqI3/O32tjvI4wpaV9X8Ot9qmzXT0sc5A34Jr/QUKM8gukc/DRCFJNA3deOcWs+SOQ
kWlQCQQAfLmXXC0QDp+okc6vE0agXN4Ha3yLAL3KfeBKlycfhKMEBTRXAOhCLf7KQwyr/PxPONPH
KYcIstaX+27WPNs/VibzK2M+2cf4CNbUngUqfQCOo7r4DsYvNkY/SldmeIIJZNPmTHb/6g5y3UeC
aL0/EqzT/335qSq1fZET8/8MXwokOE7dUu5l960wle+2bbp7vPpPTL3BV9E4BE/hgH72K5D9JU0H
BLtJxHmnmd2G2mSzlk60ZUj7AxsfCWR+d+95nF7P7yYTTa06b+dbWXyECUQPMLJXzJvsjRzEU/F3
K6dD9fZb88DOhVPRdnXRgTmsV28l1s/1x0GL0zX9rIqJ6QKGj431TvznOw9eiKiIrd52yS6hSami
1e7ylUdQy+EpYJ/MunMIh1Uv+eVIZ0c7sMol8sUbNTxgD6e8bpgwVJaWxR/SfBU3blWOmnyZvtU1
cCpi+bqT+1Q8HHPaCz5V4zAs0lHgilNohakhkrjfzeIGiL1JbIMR7LSerGfF2GEwrQAdCp8tE5N8
CdsW7fmoyMIF3Aqx2ImfF5BQXhKRefTdXvmEo9IGubkAwuPEJlomCuxdD4mGE4MmZpTBJo/6XqsS
7D8UuuZ0sM4kr7F/ZujQZnbGZlhzR/ux0nSfzY5Y+SFm7en/YB+4ixDPPutRGjsNS8jknALqVGle
bw+8Xwq50dbFMFRg0W2JOqoh+w0fw5V6dyhQ5E3+6lW57X4JdDLQ1H+L/qEnRnujJumY3GyFPbGc
rDkEqA5W9KCPewGpM9EnLYmY5I+O5NflPZD/tVRd95Y50uFzN9MldbNG0JNYcFWb507w8DdHjj8i
URjcExT5S9bCFYNg7HdP+I33ndIb1JIabqjKK0Uvly+sO6s9pz/VSsqPvOGXXT445fbDpE0dkJvZ
yHq48UTviNMOQKVeROySMJrqjVf/6TAi0AYnJo0wYsWmc9qwrO8/Ag7my2jGOIgWDjEB59m6ABnb
RHfK+xFVz1tK/nrneq0okMx20hu4WvjVp6yE9yGLww7ylLcbyJKyAKBuSPm2pIYMHznilFp68wG3
ijpKCrix7aGpyJktU7EaIpWIfcHWrxrF9RUL7P3kNwC76ABNOSXijKDbbxuN/vkpqLBvWqeERKH4
AylrfqmEdVeZIG03k5YHwsIkvp4cdA4hdGlqhJ0Ij2EmzbrpsUvMHtpKpS9LG4OXw2wl4teUfUIL
Bm4ygThUN5O22TF31EfpBKk0nmnbd9rAqGfbofw5N64BhyaCxEJJbJIUEjUneZasco8bCDw7U40N
o5XAl1DrslGGvCM/zvyG4TWWoiTYAD9v20Rs6uMAfnVrjdOVLJVs046DxZjvxgN2ebuGq0PFYQbn
aUgRgc+X2d3MMNHm3Wyy+JRQ8rabyxRP2F7MHvZBnQd8B3+z0f9mqob7VbOtZYt/JGNqE76AnGiF
D2SFjc5pHgGp0tdSWjXOEmn1C88ltC7aiOZaEh85QOurtaor/VxdTOOTs/LpvOOVqVAi4FCpBoaH
jLf8uRGQ5hyA0ZoSGStiNHhNm6LCYuhZtnNiwcNcFQHgGyw0Tg8OJp800t5zdhqej6oldOsZJ5TJ
JQnOFhzwtkX7sIS4ko92MpAfQXaJltOi+3O+xk6ji7avxMwCe5Au6nyxzOZUIg8UEl5Yp8KxmVog
ytz7iVw5AkyjQt271ctcEOyPUirHOzWWz91GaZtTwMC0C3HaMAUykMf/kaxFQ6i7Zd0+oRvA8AF0
755PefiWHpIujWg4bKUGMVPoHR619ZJ4Bri9dwscYc1iWfO05fdgt4G6Idm29srKSZnN3AXdtCNh
3qO4ibK9l3yeRlk670Vp2JV93ZDaNlQN+0eQDZvbkmJusgrLEML/M0X1vS3YzOHL5I3X88XGSJev
eZzITwhPbvxT3F0CNcB/RXcOdyQMC6L1cnFNrfYY0OOOm7bTOF44ggTUUwwiexA2cUG1Ga942jgh
bttqx4/FE2O9rZPblvj1lRZcDCaDRGsPR9yTFy5uomyjwh31rXnHaYgYgwolnRnMQGCFeHTom2ZV
Yd/Iw7ALRhSNX1QMCMJPOfLMLJLHp1PiV77bPzr279NnOY93i0IyY6hS7YcI7UeN6XLcTNUE3k8v
CuBv3SCcq4uui3NEg0LXHtjHigGH0TbhKhEZnEEPTd428atvo8GeJvsncGDbQcShVzaucr1M580k
yZnSm3vvRFTYsf9E/0V5KZJtiLmPOU6RIUBaa8idV3XRNnQgg834PuGZuh3vi3XDgQVoteEPUj/X
A2G4ELlQ+PisQ7pgpOa5WUH1IWjcGfW6DC9rXPu1PqLeRs5FmMWPk/0ODUKBO0AwD4js1YzpgW8P
jArZhGq/BHVKh0Bk3heA3WUiluoC2704F6aiw5txu+AaVOP2qXhhfLMfXKR4I7Ngv+exv7hjbiFS
vgh3Vv4LJs1dUohEi5SJ4+UQEwdvuRW1iAB+Xv5bMGFb8o7XuRmn/DCPb2jAOHTGw467QIc+2R1Y
fXkhD7RbxuxLYPGymIBFz6YS2HuWw9FlKghhXK98eowD5+iHzC/ZsGT97AnBcVFr4HYeeu+nnzph
BCEnJ01o/RE1IuAZJQ1+rob04KbG6ssJgVlqEiFLdShZnOfiheFvQAPjVlYitZwvJkCW+t+gzNdb
fEkhrIqB9fMAW2w5zk5PQferaMvjcgsdTxcO6+b/mcBE5XeTqA3voo3sRg/kuL3HElsOXOk/YI/a
n+fXsnnmN7SLVP0h2v/U8xUqZO3FoaMiuIPhpzkBk4MbhNpx3Zg7VvxLAWzwf8R2ApF4iJMEkL5p
AL29P0WqZCmknukT8nfXHnV9039iv804/KvgLj5MCOE+60W2AFGcHv64YDfmMwf2z6vk9ezjLQGP
aszVThlqeTfZlRWFms4z8TBxsJl0W2ckY3vnZwEgcafwH64pqX1j/z8iFGTBr61Ln6kE6dcSa13V
a6KYC7Jl9W2ws97XgqNrcabQZPcQWg3AacXyYJeNcXzKT37seu6ayA1g9oSX3DThLxV42jBOe7tR
zEsCVs0nlczdzKclFzm7Tz7G3AFozZfBQF/E05tFYbj0ArprdnEv0BoLQiyqW5BpaqwZMVJheuWe
VONy4DsDLh1YjpZVcfgjdHjR28uevFxVNnigR3qh68WvhS1fkXEOaZPm46RXo81Y0nzAsfLzemuA
PjpKPLS+gTdzUMePtRaj3auLCcJmTtNvo9q0GkJK5TFnvkPHncy7Bo0il6mP1IEUFMJBTkJEWCko
bXsmp84moEMwgoiELFKUyvlGwL6/zQaFeRF9UvmzKmpkvYEjl5X9FdOrJVXWqIQukEjI31YRpFAk
jZdyBgyynLQMBeHSYw0srRpYlfCS9iS8azQhEkvR8EdhZ8FpkUHWEYDJaBfa1enTq2yCnKSy7vUu
00FyzNKzXPmTtILGe47+An/Djm67XLckEZdhnTtLj8RBXydTimrTW8xz8BXp6tnkmWwpAVrcLYyP
9UbgBqDBBqtWA4Gfon3+5TulISSVUHnCZQp5lEsMY2r44PygqjCVy8mpF9o61L1UWqTtzL/uBGku
PLgR5V1hnnFbLPtGe/WadHfUfYG8sbsnXznDZoAowdD0BUJxydnCNgd04lrUEp5v2AHqU1t3gYLd
uLufdxYmATzfbh8cBEBpIKwBnMalIfRS6CRdKA/dOSZAzBHVPHH3WceyInPatLPXnewJEsfFmqfB
oMlSt2r0A5DNfJ7Ugu4GLbJMFCoc4qLj1Zqw17bztvTV9n8ItyrH2PoqIPcRSBoheCoPqTNWGG9T
a+xy/V73v3+t0hB+FrsRtv+9QVWneodwrQr6yHQrvPRvgeMr1ilPDFTEQC00bhabIst3u+Sdo71R
uYt47iF33f3YjvCjEyAHoIt842kdkGoCy40UdBvm9t95py6l90RyqlMX4MyXjWeE8s+2avIwHxQ8
Em6X4o/sCz/ClBLO5Q2qloS3kH+P79mVuEPN4vtCJjHOt7JE7rhS3ZE8hi+iGnWwO7sLcACSH0W5
VXIpIyh8/AHCLc5WppHF5EFuLFPYgHk5NIaKMZoGLU5arVvOvRRcJZpHq8a6hk5TuYAVLo8e8rCQ
htX8g7xVS5O0a3zIdhbgE7c+WdUIITiYnmN/rzrl1NMsy5dhon3x7TE4rzayvxJ4v95eCk0EWuST
4vtcVvVEmasgAhBU6rtyLhcpeopzz0zzlfYdDOtAR0EwW/XsMfpxT36KkYr8/+uf3qvM/4lNnLf7
wNMA1Rs8XsFv5M4dZTJXKtXH8fnAkXADwaU3eP/6HIj6qin/22Uij5wscBixGt6YntCr4B89PgpP
6tcQ+St9DFg/0iRo1v13xMhrXSB9B/7xM1DBdh1arAD9bMlsVCjkczb3jqvSb9bfHJzbGOFagi6U
hk6a5rUMb9wM9hJADmMxrc/1nDdV/zEROJ3Hb0k+6Mj2RczoozAz8Rz1TQ1+23nRCwTmzGVGJ0Xs
NcjJd7VH0qFHJ4L4WX30VEJq5NEL1agZG4ZawxGy11M8AsOfBJMbRn7lc4+krA7NhrOg549ZdfzQ
ek1CD/su7T50dWpbt8ZyyAw8emgiGKU+zuLqm4RRkHE2mBW9h1DBAsRkK+5wCfqptY+PfBVqi9GF
p64gXxdnBkGrNyNPWCa7KthSBXACEdPxeXWxLx5H7IbtbQcUSlUPmyAnwh8E5YnMDwl0P3HdibWN
3wwxM9UYTXyXYeh5DZpQPIGuINng/RMQKVVxg64yqkdpLSn0QMKjcHZiIUF4kukiOEhntAfHvv1o
1bUeASNLJsBJ4moy3tWEIk9cqbaOHJyqZcPlfPB6UigK+aXB0etrbWwdP4I2yKeaH6j2x+3tQVn7
h0w4cjeV4QVo6SoMyoRgW6V93xXdd6Lycatj4881MYbRIY5pj+bERQ3ja2lXY2odl16dIwqdSxMS
Ytpi87KfssJRmEAOcRgTs6l6hIHe0YqlusaBBzU/0ayjJLBtc+aueI/3T0tXviMhiQS57WRxikbr
/iwWPdStrfyzcXgc2tg7q3rXt6ZpRtfV/DD0UWe2NeAAIKalbyNAWbhX+FJ+6gQA98R4DlQTSuxz
SiOmjubVv25SUw95vNH46TbLsqpIAq9WtjZQ8k5rl36CGFbVjB2v4r+h0WT4eElzijnNn10mmEbQ
XQEn7fAyIq+QrNzv9HwOmgnyfDGPTrAqqYC8h3eWEa02nWuVSn2YKEE5euRiIBovuPIVT7stl5bd
x8nBufE8w/w4GYwM0CLi5s79HF1u/Dqie9SOu+Num91Nuaipz0bS4HZnrXd5hlaJSO5cV51SpQ+L
qPy6Mm11yZmtlea+deJWxG1sTK9BLtusgyZYtdUpZqwj2UEMHn4tZ0yaVXQU+K/WsD7gXa74oKko
Jb3BjPSs5lesJzqrUpxdShHo0+nTdvuLm/vjFzs67kGAesydEl8wUEKAZptYEJuhPpYQS/erPTi5
QAvkn67uUwptqBxHGxQ9iXu7yMPXc5ZiLLkDxf8qP1Dn4Q4t2iQcw4R60X90Mm4lLLf7P/c4Ck9Q
O9LRa1IMM2ZlIRglTmCAbMQlHon+NQGwsOW31LHe4jmn2kw5g2Eh1rhJ8IIA4bIMccPHxH/RMyyj
tQYVE62ti+Vk0RXDWzRwv81DAfilmjjQP1zc8xxEsppbADq29cOjssenXr+/1YSwau0erZS6OeB4
ImJyKMdXuOjzvfYh8RYUPnAO89b268EN5/ws4HK/vWL8gFmBYPppgOZtrvpWPwwLPME1JQqIxipZ
rIxWceJ89qThLs58M9TYYsnupSHyJRK5xKD4k+xrHai+NKyEgFhteBwe/vTMzIyY7rD5JHzbVoSB
Zu5IT/Uukm5eRgSwQW/805zWAao5WnZgUQOxMQjBzYw+g/l6vfE/2yP1oe5atEq2o1vhBzH3neib
BVsUFjltuMssRfJeC7ZBX6DJgn7mx3NkZQfelhw11SR+K8gwdx+Cw/38Ly99Tll4QkEum3UWqXtc
kuvrCpz8I4Fv5oVOsC9zS6awKMuqtNlBfP3BQW6KErxLWYbTIB6YpDC+9ig2kzdIYRitrYPW4k0C
suoCl/d9Cn8Lblde0knwSynsaP5s7JFVXVnKuao2ke+5k7k2Tm1sKuEwtrn38Dd+BcBn6HIoFD/v
1hFwSypJMVux/VbnZ5FrO/4DfZwQ+adWSDJKdx3mDU+i/spoAoC/yOeRoy4NZlHFuKJmh96dvoX5
7uMUbNbCITpOJ5LzNScB3nHo/JfUfpfyfq76qxTMp5BGeuEixjPuwlrikx6gt0gR7eg1rAugoLFF
xG/IZ+XzG5A6p8ZIDQSNyceMKJrH6GgppWMrQKJC+6cu0j2uITty6xMsfv1BWmq8FBVNx3vSvsDl
2X8Cd/lNCwiMEswCxQHD5ec/36w2JtJttCMzSc1OzIR7n6NXsRlCh8l9lMwrXQgKya2UC7+xgf03
oVERBwrvTeffpGINuAnUhlFM0S6hhwwGid1Ch9vDG4I63l6GMgV2xu1CD/WxUt2+IdmHFqwyjuCr
WKnXdqr30tNddBTET8qDSYla1JYmf0Pb200xJ43ql0Z0uxKZRvPizULlBFq9hEr3skc+vKnPmqSa
W+kQ2n70Qo7Al1PFB0Nu4h57G1XsH2LgSuEwu0MAE3tLT/BpD30S/5tZeTVxN4RoHCSaKqqgykgF
6hEnekgjDghZqmbo6FEX4vtb3lmB3P+9d+3QOQ2D0+wDJV0nk8iPY26TrAA2KEfMJ+t3o0lrE6zN
XXD7vpzRXUgkQER3lu1b7pgZY8rpw9DnMJ2dNq03YeITsCY9KqGd4cK64M+OuoFelVmNMqipysfJ
h1XV2AC0Od/zwtmBGS4afnugXPItdYTlpJP6YySXV/O58MnmDjDjafEcQQUcyARTYJZomB4+dwLO
R16vywpmLgPzgbmxzytuOJIsPdz0N8DPpt1hwWqp3QCt6LkQlK1VrrWNVgH3bx7nioKaWL3796NW
0QN5nE7mjbod0jG1KVkOH4hrKedCLUh5QR/RU9FuWO7Ime8Z1AShyZVaSBhJjUZWfZk2mOBy0n/6
rSAGm7mQFTZNxuowjG/t1m7QIZnfClWB8WpYdLK9niIDv2Ag12kdrXm3MRrSJ2opTBQXnRtAeFt2
2P0gt+gJbDIso5KtIsWUgHH2/4/tyavJuce4dPlMFldz+enSR+AQTtdw6wB2K3Qhu2N52AfLcSyS
LEf2+UQkI7KMuFb7RgCbq9bj28IqK1SuQoJt0xB3lbEOE1Cvh/jXD5WY+NJTXVl1h0cFigF8PHJg
kJ7ObXglgRkz1PaW7X7SFnS95qnB1d0ygll5C7TlwD24xbOec7cUJY2TRyI49kyQUhQqtWyX0sMZ
/81fiB5UZ/uyJBnNQahWPsM3UdWonpxuGFSz5qwxiUNV7J2Himc+H9g13Opdqrr6pSDKXrYycLJp
WpP2pUtqQVpm+cDqI29KWAZkFxvLTBDX+z4BZeKtHKfxdbTWmBv6QNq6eU7iQeHbNZgOWVeoeLut
tAgLNcfofPVaEdcH6+F4M/4MQbKLoFYxZI6mY5LMgCb2pElgCisW5leKGY31lFojwTB1GT3xUiv0
qYmgejzJqtoFYl051KG4RA+DINBnDxb9oQZHWTKNN9zgS3C45UuEN3RoiE9XwyDBsUTx/ReEgoOr
90+pN+ykz7agpRcNXJciV5DYlgs/Z8oD0IhpWEinGq8n5KyzSeY+G5Ys8nUlG01kJh1ZMImdFqkw
ebp34QlfPGvErzOiFgFF5OnLxWPaMAM0rP1YLJA56b5vNiaO8m6lhtezjTZQPyaF2kupTiTGbaLi
hsVDCFvTZl0qDeaQPn1fnLiZNhtJJTrNBqHxxdiJ11QKcb4m0ih0FQeDZB2nwENFgCt8vQ+nevbV
r0bPG0IXwYgEfGDDkoUdgvLItrFL0tAiMPcFcqm0FNc2bB+TqlwKksq1Sap3GooIWWtQ5/rOHBqh
PTtan0+UEFnbTOaFh7qqvyamH5ENBAy0APHFpJvQwvA8C4n3kF/T/J/4jsDWUgEpiHZtdfYcDCuF
jD2ECel+ssvuA/doA/NwpkSnQ8s3I6LZK1XTU3gNpfTDMI5tcNLnrkkJEZpyGKEdmO1/gmowH91j
k0FyQWoV9dbSEXOjFdgcDAChBxR1hfkOkeLrvkucQmgqrUGzNZsUVXM8UZsZVCjPL8JPCwr64Zbd
/EipXQ/vcINTcQockqDM6TpmhaUyaP5YuC+d9yiyVIH+1WX1sXLfp+HKst6ZYEX7l1iAlrei3aWl
cZs38+ld2DzqIlLZtu9UgOcmTqwHv1Srg/m4I8gcWp6Dp86m45t5PPJunnxFCeZnnTcyL3bMf0oz
sMblxHt06zMw+PfrDE62dVl9M5/LnTpQJxMpnlChFDMVNah9Bqq73aorz/Fi14WXUChYccDc/xfV
yhHclbjLm/NspOybJKfqpJmR2bEXRoFl46z1s72hIV7cRafQ9Y2KUdgpeoAm6UAPYkDv0Akw2kEt
8VpGDyqS5Jrs6wZC9NNTKYYX6/sRDevkyS8ikAnZgqs9yoIkeQ3QGlPC8Py3CtXYO3PKLXhPkt2B
IhzSIwY1EgkGYHmfSY6ikV+YeaX+Gj4eg4rlm5KuhBnjnxDV1KS5ZddzWzX4u9fMtKWanggxK0cR
lndGzW3l0GPnaB7AkBS1jbpnGGrFpYQcZh6H1TDBvZc/Is8+stsNGfPHQMsg0mMq+hpnX3ru9DQA
BUJdptwnDEQCWNktBbT+5hEaRWYYgX3iW6VgID0IFGIrZMwT0alM+hv4O7ri1ZMTmlG//UISEZ82
mkgOO4QsyUydwTNhZZM9G4PE1R93NBnYkklMsqekI34j6GNShnArg+M2Qeut2Ag4xeVGmo5XzdsE
tnYkiP05Ro3Noc+ilP2BUEvfVogywmNPaUXK53DlIUM6cvmx6T+LM4ngsGHoNJdtrutMnESimU1W
0gEChepvkJAjo3Jw+gcF+N2v4bMDkQT3529FPsW5yXvmRqey5GcyqXuMEjmSGfLoUALKiP5gpDFV
c/aXQPoUteNqjhsTLHXlDLSLsaBkUx5ZwNg9VRgOf1dKPh/mnn1/E2leRy6/x/canZF2q8Azx+RD
DU9r//yfc9xrzErJGrsshw2+uF7PXZiWl02THtvKDixDGCHXGoUVYRCDSvZBHuI8adpspt+zXkhU
ChuJcZvX51zTjnTGRUqgY2g4g9YZ4grsaOMHIyrmSlsxhygx5eD/7ZLAfTXoYJ8FA0BkwEq8K7kJ
/QV17I3+/iLpjgcTFF2rBao/seVKLV1D9gCPwHdkkw/mbaVlVzZBkfrnyM2qkLHPm0IccLMjg6ip
ovz6sCyjINJuYOH4dbWNUAcVaXNbN4N1ri7Zizl0iEVibyiFrPH80g77HupBjVqEl49TXTNh7r54
yaBiKh8lNbTaJq3r0Eg/tVunEr+mYR6SZB+x0AoLSMseMMSJUFDSNezNlZcc1DGDi5urQ/tyKO1f
OjxU8kptD4L6Hk0Myz8e0FhXRgI+00Kprf2jJ407BNyiCo1pW7Ec2rW1S22xsocsJ1yVqtkHxNWq
hb0VNYTDE7UwxqyxCzFkaKRJ55C+3opi4GTCWQfddLP2kCSgbWwEkot6b72WqRpdqfSpgCdLn/dd
ke45B6bLYAVix7iw6RHu3EQvgLERq4Dt/XRFhNlbaWUUHeVdG7gnztfM+MQfqht3FTiB/7ATAngi
Q+Q3ZqrB6C6LEa9h0BMDIPMa4c5T/QYzYVGzTSPvDuxyYPtfH9qo92dSIoWW/gCeIEtGzH0c7z+b
m9996LtXgC25S7jHvkUcdhOUu8zS2jUjpeGJnLz8Kd23RhAs/3po6+0PQW/vr4rhtX4bIcVdnfC4
zuEBVp1ggMxUKgKwRnyLk/P/4nFULh678bVlIfs2iVYnUgnzp9gMZQSrUsSbqIgd95CNvpW7dJyA
gOZ1mbNve4pkJwKeUPkbLorVntfIUWmNM/fXg7Yuw8g3sler+q7k8MJKZbeYmoPpv1yOBe8zpPWQ
+WQvoXb/yVeBWyOqeBbvXXASAn+JmlbkzptklGsCRUCmZjkdDL723VbquTBh1ZqXDIuI+4JqTZ5w
m15iGv8zr7NIlIsRxvbrPXXcDjX4IOyExnjhcOegIrz/QpkrYQYrDbIf88Auhc0/Y6WUbLSVh6Kf
hl9QIon7+aWIDvJwfY6scVnuLdAE92NwTa0wTQ8kgT4GqFULCHTXsl6oqvhxQQM4N1X5FLbmWU0d
+h0UoTKFF1kGLgYOs5Q36PZb0CIlNV5fqYUOoSJJtm4mTK8Z35K0mggMj4FW3uuAcOnhMkTod+Ba
FujS6CN61g6tMWeDjdImVYaWE5bsI7j/3KuPKMCB0K/6kTKb5tU0x3g5xRN17xeP35VlSECraq9a
F9sqTP8ufLjtb8QhN9e+73ACcUaGdhVRt8jtUiGRbU9KDocJviaD0xKoKWXxEV4olxUCqT/9W/dF
h+BQKq4o0AjUnFf/Jm9ueblWcINGHWvl+ueCR18MBjzN8f3yiTfq62XiWAGxNE3Rn/gWXgLr7wRY
+7O44AuAnyw0eW3evzQRdr5vwJuBAib2pOrakSQj0VcrpWmxFXkAxM3yBZVwc4Sqe+i00vRyvgMn
/EXIRuMKxksA3OldBg1cLPYQij/+W4ouLv65Yy0BKpALMC/0IeukVB2at3eH+8jKL9DQS8v4blOD
3Gc/4K1zOXgtA9ECJZX6tDTWKBfHP3rqJ378rHXUX/nj9vSUeeB/4/t7U+EAcms2kxot2gzJYnO/
rCvT+LXX1agX3yDe7Cej01UGxdPzvMY4DQeo1MsvAZPsLjac6ZQMsfzV4JCFgjDQiz4fXOFEWlXi
l4pNxXnWcjN7cauUCQ9CKYQI0moJj4M+HGHrh9ZdETzY/sET+tldTK0XwuBw7amahPNjMpVZueJJ
3f6BjWwNWcfZVjkMeBjzmO6zZKl9QQ5gtwbaPQ6i1yVqfTXqFCKXvPPdxU9DRk+DTKAdcDgNX3tw
SasY+aVDfxWErUhPAZAw9S+PDJRdPkroM/2UMbXxKD/hkb1gG75b5KCtBepQ9tCh5mZrraXEXCM/
ycIA+6++pImyWHjDC0HfoymQro3byGtlwZ39BKFDIraFZb2EJ4OSKcrtVJ1Q7Se0CxAgEuBiiEpu
oEbPfQ/jGDmsMhcUM43mJmvkXsZJUMyrp1dygwg2ZFu/3XccYHGn3ovhfg+FN12/5ieJ687KrXhw
xPv8Gs1clEIAiRYlDbGpbhS/8PhfJH2tLy8/QOaT8Vy6VFpIA9RauPeumuQssZgUeWdji4qvcZDj
SatjR9yDLjTYAGDUOUFrDIfUtyarEHQAncAQ6IiBeJqQ5TacANVvOYTkmHfyoOIGwMmiCt8h9rYk
eyvadPZDLnMUif6efJUii+r0NrbRiTroH3mlu9j3o7ncuGYndenXIPuiJJP5OTFtn6RqJDo75jDk
P6qppgsv94vy6DFZONatNPlIMyRSbGmYtVFA+v/YOj45cbBhgjdwHU7WmIM6BTQtGs4PYmbAAX3q
+UpcZFiyrEAVC1vjU60tf2TIXr2NiI24Te861BSdB8MPyxbdXoOy9gU9vagRrV/9ICon05VlR9nC
nLRBAwML8xcwqowBxz40OTP1rPQhgKWTRzOlj9KJH6CQuCP1bU5cw0vpiRjy8JTB6nqjnDo4J5hG
KpcH4mQdA47gIiHHxzuhp9jxeg7x/fz+/SXR7+rwDsSFJFhNBKK5aS6KZHPzH08dqhawHtNZ3YGR
PnWZ/6xwvRwDaLXvVJyoUMYVj/4aDdoKZddeOm5vNMcX7OaRCqh44Skj9Xq49CmE4LvjG2f4+Bn/
gx5u3JBg/S+VNnEIbNf3FtZasj9IulwsRwIpCDly4MhbM897zMG3RWqZH6/FGqmq99Pz6jixoidp
29mHQrvPVxT0Yhxrnn95NV5mxYCu/XaPNrugGhNrCp0AQLFciE012znhXVfa+Zq2f61uajv6UvZy
frBgrpKp8zXS/Q3LJkZ0RAlzthK5yO0NS2bPEvfu/5j2jNOwtbiZCXi2YEBvMOVBylHyGk/yumkU
Rg6HK69SSMkLpWUbF15rLn1htWO7Idw5GjahNYHoDNSBpWvQtrEf9DgH3nwjpeD01RpvpsNVhGjG
jL01iV04Q4onvYUUqja06w12lQEq3Jup/OyMRGlgA6l/uQJ2yGEQ5pI4iKhJeQULIOI5AwOUAiMB
K3y1mbk+HkJhn1Ha3ciyxlXmYlSGvRNv7YfsAyPlHjfRmjKoiBjeuTKCa9wJ0z+gpA9ZYU6IQwB3
/ipUXA47eRnLDnFPRGSctLS5T/PmIXKLJT0WH2Bpg+5u7nN9oLfoGTVV8mOmWLJ/ju0NxKXBxRG0
EHI8uMuc+fbK7l106E+H31/UR/Qtn7MXrKEWpH3iGnIWUzCl0/AlcNQRX1x+m8ywgi54Potx8TG6
6jFHC7zOBA8BsBASKnLh4t8LAF3DxXi1/YMU4DfGBiZEjeX10ncYugU693EIQayy0nv2Nal3Yiqx
cnpCKZDEYvDSTR5PpR20QPLTVZhn5hdBgSHpJobMV/F78vncSiDQjNLDvIPfWDlzimPhdAdyI+mH
j7Cp5MZGNRv77SnJRl62QRMqNYvc2zL3HrTtzF1xez7epZcdKj9LJlns8CjZLZjf3Bjxm7jnvkOv
IgVCgq6i2oNm1BjL/TS0CwF5YGKTbj1a6ZqgZvxXbvKQyd1g26c+akpE6L96Ry1MyQNupRVFcP8a
mPyqmizAdDwkz3YakkTijdI3jUezoA1fkiPBoqPbuwIk9HCqIU5rudzBpetV3l6GPO+m9/Mcb0Nx
uh2H7Ye6IIeSauXMR14m0F+Vnt1CTw38yrUnCL5jevDLnmw1Lhx8p0o9KzleAfOIJvlh/ssyp7YG
Npa+J63QN8XyRAPxUqmBo0V+VYzBR7J0jSp++c4SBx7BZaZSTfblrlgGvqMCbnQuegKLu8+EnFjI
Zx0HgT4JleYMd9lQH0VEPIvMJrpg8eJIUSQkcjQujyzT36PzxovezXrrdH4vLVST6lniRvIp+gX7
EPHqA7SgD+xt6nbm/0TKQ6zKUIzOTEihyITWR3t7ZeyRenarMcsnACw4GvJceVSxFcpw0ziUO1Zk
ZmjZjFkmmaHUbLNXhHud/yD7VHRrIq7nMDlib4RwAQEjihBwKyB7lqHBLxri0GhuGMjOiyIk7t1o
sXxMDqYjJ181cVyTcNyHtbhPKzJxH9wIAfJuDi293sFlFwrIBk7y1avzM3aukFZYqRARtVZr8TJf
E/HY8V1ylfj3AdQ7MDuoT1Qy4mcs/Zk3ojgyuI1qxNiel7Z2BgtaMa5900ns4DHLHS5SB0Btn71X
wvM0VWcnJQkTCIDOwG0MMmZLRnQKEiiv5J9rrl8NbvZj2nYhaSWioorftEzoAjI9RZwtAlOLpthB
KK7qVESKGYvctofkT8H/WwpShnW5HVcNmbCp2vsY29ieacMPVnm8Vb2IqFFFD4gQnUYee4ee4R+q
aFe8TkcLBJp+RW+JkmaXmZMXtQCMTnS4Nhgmxx95aM/YNhqvhD14DH5/vVnxqCiSKKfXP2IAkN++
qepS713CrfVqcIx8tx/rl68mb7QWy3pCAu2mDnZuphlpmD0MBt/aXPaE5A+i3BG+bvAEPNR6E8x+
ECtWvVFXk18+zPCm4jqA2y6CwioyrXqZYk34Tg5jtqhOqZG093y3N5iNis8GthqDzhBD06Pa9CEK
PB0cf1KAmTpdKEudXkv8Lw12BnGHPcRge6z8X5t01ogGlcMDHE0NgixvlvQwkFSCEIC7UBc7cYbY
x1pT76f3IhIWT7o2t4fgQBUPmcsYjL/0PvNBP75b2KOCUSJ9uBv8kfaxlFPeC/kQah8unOXcob4I
++UbS3LIxBnlNxXC6+zNTadtoVen5t+lTo2LmAXekW6yhazg6ds2S04jNSjA7XdFjETbFau0G5Zi
FlB49lh9qrYQLCiRXtsw1K4lcMP2B0xRcwKVQQfGvsIv642Vekiva42RvMKHs+7B/QtdSFUqY0Xv
OW2V8PzJbVlC8sI62ZRtdOsKK1QnRJu7yurdveXOOneoDVb9GYwAitdhQ+zYTXUJopIXz2xj7Rib
0yNkEBc73xS0joyF0gmpoNzrj1td+ivIeIoSTnMUTrguyp8KnyxPogPu1MrOnkR97HLBFSweVOdx
UbBLWCZNpG45zM0M+MzdPES81PzCO5YhPn1ly1Q2o6fOEQxO9x8Sb7UsvbGjO2i4mk30Aq4hfMxn
3r/+6cKSexvW6LnjURLds2UBDPQvzfPHVMlJndS4Kcg4W3W4WZHel16JUGlixuYkTgQlnM5rmXqK
p2S9uJ8qFNcwymmRldrfzCYC87/sC70uqwOv02q1vWsrLB+MUR4TqD4sCQ0oX1ZR+r/cyFqgFbcG
V/VvzDQP7vqNyVO2j2WhSwGOodISyi9QS/qfOmEqpgv/wDq1aKmpDt4NRZuC1+WUpwOdUmbBmwwZ
8OvpCGDn18LalELQcKnQIndaFy5mn/Yxag0RD553SV3Hvj8pmGdN7ap6HgJ+HljJ2Ox4BviVxWSF
F3NOUZRsJViN3LTj2MPu3M/Q5KqRFIPHYNuowE/19vSCT/N1WAnieA6AwyH/mIzvBgSs1KxxdYTZ
mz/7qTcX3HEUKIXTTX4ds1ELAxdQ4L2KXg0PQ0HeeQ13fG8K1BAEHJHs77k8OXXEd8uoCgiafL0Q
Yv0hCkRQnv/UShrq/qFhGnV8mAuS7N4cPvGk5kuh2WYJBxUvpemF+nOek+iW3pReLM/rETpfXDaL
SdmaFKnXOxpzGXSAAzy0/QDYXfJWS+n0lZTaKE8Gkrjo5NxwEHLzYuQP27yyf5zoNXyivim4fiZB
osVPAbCZw9Mg6s+b/fj8XPS30LbYkSQU3ChzknmuRsRJo3MyxjN/yddV9SER1ANMz+UwYVaQz+O0
Eu6X6dHcquPZ6vGOoqe07AEm8oNHPgr5bmCCJNh6i+8Gjmc/2iYFsQvEPgSXAyi3MZAhwcF+PmlF
J35KAHXBqzwW27Fe4u6IJ13ZRHQNP9/Vefs6DzwAf9ciB/tTIXeTrEqcPhiO0QmCTLCiCiult5HB
gxYRS41c3lMZM4CeniSrvb7v+VWE7UJyPSn3CUnaTm/2Uqsmce4BN9D1dJWc7xddYuikm+h316NT
HuPI7zNgRZjHvckNxH0bOPtTX3OJGsEsR5aHQ+ioeJ1zlmHrzJ3+66WsDsmiO3t5EI0p7ml+Y7q0
lVrwGhecYq9rj/7COA88VNgSjmHtQ/RrzfHoG5g+krRo5Rd9+3JhzqiH/24nh4RgsR70AXOQAyye
6qjOUw1Giyo1moUDAgGu4P9JlnIpUeMeNFOcBtTYFXQ/gJpx4dVQS5K8QK688GzyfOTD2OKPDeNH
DloSL8b9LzshneaamafPGtdG2dia/ltci3BqDpXKNcqmf6jwagSsYD+lwn95U1hCcujYWGNpOt3J
s1Dxj1GzR37ybO9XgmoBsJrTu/qRsYjn9BazxmHMzXwESeBNr5jzuD8w0Xyke5iJeEK+lzo1Hg8C
vjfUzUcIWY7AXQigaLwfXbVBidWMJQ55BRlrG3Nwa7gHYfUZuYw8tYvDXNm8Ri43b1sBFB7BMVo5
qDg9I4g1VB/f6jUv48UeGWCKJ3G4S6DAKSaTY//TROPJutvhWgeiwxhqHcED7Y97tLwosJsUw871
3wNWs9DsO7MpObO//yJsCrstcEbS2GjOO7HfdUTGI9hHW3Zy96R74f/SnQLA3ew9GTfSMLZLG612
hNcktQRFBzs44usjA6E62Fy/3e1Wj5OKjjbOjVVgl+i4+2ju+znHctI71ZS4tQqwSj3P0Rf7FzEb
/znYQ74/womwz9KEUa2cgh1cyWGConzaGufuoXp6aVaqUWXAfHMZgVoGXv+g26ZxMCQekoDZ2s/w
BDElRriJuxcn1dxwLQiMGFyWE88w5dd5OngwO1pACdYru9IxI9KwmgWumK9B5S60aih+fIn4BczU
bfWl5igT4e64lKy9HcRcyzsUo1sjgGMjD0eSCjOl09R41VyUfT0KG5XZF9aqKOFbvW34apTWpOia
Q7gfWFmyFcaeXg6NefnbmI70/b5y9d4l5tS5zr3a98FrCeTp6/mfQZq5xNbRHj8Wg1rjSAibtyPb
JHVFMkzrtfgGpHgqyd3VLeuF3rHb6CF7dWVLIMqOCY+5k66NCrCENYCVnJ27VAROsWbIDNlNVY1c
Tam9NfGYsa4Rz0Umx7nG/wncQ5U8gkUjuVV/pyylCvZtUR6R1KKmGXbCITaJKVmyFOZMilGe2pLi
mANB2pT1c1ed05Ilcev0LjIZBWtwyt4rDuPF9c3LcQ6lyRbFY3itLLJlqyujH6JxBC3IlW6Nc1kQ
RJzuMb5hqhWzCXi9fQN6jqjpun6sY2jey/XSQzlM/SsituKD1VHv6DTJ2zX/NYbN5qcIXCQp56Hu
cCWe6UTcxtwCD3q9cTZJyE+GcnnkNKIi1h8C9UL+qvqheiOV0JGLCe1AmZ59VoRDr6wX39AzgikG
yVF95V8eXngMkfGG5KrtOqeXSFycU3zSNtgpiFmDXoJ+K2kua9D4jdvxiE0hdgHDnlUOda/zvBM2
ZRgU9g5T/Sm2n0VPmVQ/Lt8zEdzu6YNLXRwe1eSeuKoJSS2lA9NrSwuPoA2d8ULk2RXOoNRvLG5A
kyJuePlTYtW0w/tiAPwMzE6hX+b9TAqbgd4FUPIc2x47ePmfUy0KCMfgnzfBu9WVh5T4FQMeyxh+
uKsd6ZDWgPB+FGOBwx2CtLVryImRFTYhEemJHwdyfGjb02eCidjU0LkIQ6RxeNA42q+V9G6ObkgI
+QhpOJizwMKDxvKP/btRPom2bcczNtnqy4Tm6DWM3JSLiog30V9Wg9AuYq9gC2arF2P2rpStWp/m
lhWsfsBDJQ/SPZ+U+KJXwBzW/Oyz8Im5LGBgQwod2Y5DQSF5DE3GoC3dKqHOJSdU1XDnqKnNVuga
/7SPGkKH82Y5/Xj8bdW17scJaDqLcUb+BjtmxX1uJ+OUDmAtUX7VjgHu/yg/j6M+rqeyuSBghrIj
o5OD6w5NNYN/Pk3uCnV3zDGQf+5Z3siUz/2fy64+6HPos0ZrbEE1hicFzEmC3V+6tcIZjLyqxGkS
zEoIpxasPsSaJ5ELwxeMjUXlZGDkRPy9YT7Pz+PY+XE1/mCOQPZpm1ztmdBwHrET27361TnGrBz7
A5hEq7qSC6XzovJ6p2gjfw/lRPOSDWvsNO4LJoRgQ8etODr+OG+sfJOBOcrpK3dSftP1hFHvI6pO
OyW/3StL1ve8kQwWmHZw1hdnTy48HAv0wKs/3/8QTvOaQ/G82QEptLYacF4/X/bz6E7vHIS55de7
FnNsaCru/ZsrVfzic1g7EVYIthR8W15a8glq2sPHPTv/UYa1n3xOttHb8MOLe2NLcSHB+hElvMpw
11UKf3vs8LnIyBOeaNE6IKPIoGC2v785y2VjaPdc/3cnFEb0k1FsgtOnnD2iTNkZ+Rejw4xJfHM5
g/U3uyon7Q2vtI35WQwozwJzqMF9wq3tT/RVZQRut3Qn3tru2aCZwYK7zwcwz/+vugJGojPQydKM
fjuue//VJOI+hpujdKRhkcM4AwIZbHwmtxTNJSo6HbXgMDs3TBjnDOOXaGqN0mYfGeR006R8xBLt
EQzgfkRfFfrBFSp7Yj48ke040fTVLWgtTPQvtMss7TUrzsyJyJ5V2q8thzBhH7In1G4BcDo8Xqvg
JvoWNZvagYtsMWHcv/XOI6lp3CODqmr4RMnfx7czOl7qYBJ6uOtyDsUC+FNv7HoJUuu/q51cpo7g
fJwMlAsqefFqBxfgJtIw/aJrd6jDbrULSreH/g5WPAhmEDlhdD9KpstzWE1F1udnn7Cam/TnF2dI
tOcPIvx5r9285v7b4yQvDnEcH0xkuTDL0HDYIkHCf5Oh1As4K8EnIqLb+q5pfzb4QGWFm7sz+N0K
9Y2m7RPZMdcLKXZedj9gk+tNv3EUrsI4hbIZqkpCixLQ8/QBdMBBG7jJou3hJ4DHw/93Q/1ypmpO
inDAVhnHij2J6MMNC9ss2UgjktmpdtTUvsp8qRxFo/QTdz8v1/hJiAqgkpSZTfK/QJer3JWHqc5E
lozXukR17aOQnyUdvbnmxnorq4n7TG4XC/uNrU8uGK9YyEQcSMZnRt6lJi1RZK60kxQHIVu75xYe
pk3E3iV3dUiJSc7Jm9K1kluiP8hmnl36nxrJ4HXZPtZI8rUiDyUJDvsay2rQQT7KKnF1CBxZgYtO
Edc1QUFw8M2x01NGLgqNZE8No1UzD9PpTphs0HexIeKBSbDyoVIDCaEhCTEX3RwFpytmcDeZnMKq
kuQG1SXVhIFFnYHVL7aV3tsShMzsvJR5vho33fTsBwINFePRIX651u55gAAMyfOcXnmGdcJ+1gDh
VoDXSntOndIaSON17YmICQJq2aQzhJrMDhx/Orut+oGSxXZmZws1nw2BK3HAX3aPhmgRDG4a0jy8
yQEsTbU6Bj5C4/D2Z+3P1xd0ui8JwN6J1gw/EKALhwt/wAYMyqB/IbX6/UiINN/t4Bc1ehUwWqO4
IPl8lNUPtW9WbCanZKx0I5QvfopT1uziDOta/bzIVaINpzXBe2et5GLc+PTaDWOM10T+Lta3vDXB
4V3ZGYRH0k3Ix4ZyTUjdOuf9eIJCFLFSxpsCPiJQssaruVcwuGr62sI2rjOA1kUeg5zV+oTJM/2O
rivll3arOJB1kwt13Xogfl7cJWdcTQvKibwRY0FXPLZ3ug9r0NRpgajsHPXGsZpyZBLmlRUnr3iq
BYO8e7JfFLi28fx/ahHCca0fLVRRg194oY2cgevigWi+PNZNGVTIwFVR+Zf774vwxXCrLwi9ftQl
y8yUrutyx6A2cgVDHDrJmPT6w92+rR6pM3TR0M+0TMz/6EwlP01vh5cRAa4ko1UNXVEPpPQYQA/+
S38GHp+R4erfaIrWE1bDoHvBVaJt7sNwHLygcPC0xoN6KoIZIauV+A6ay1mYMTzbegGmt+FJNDH0
J6T4CrUwkll4MkNLeK9/UUR9I0WdK3rh+8a142BkoG8r3lB4C8BgLRgAiMGIckFFUiSWPrglmIA+
eqh3RycomuhvTYYPYUGwqHBNJO1vqJACaKLkFF6ikLxX1DLt0eIHzDyACULxPpnpbMJRqcppj9AV
lX+YDPI5zifBm7PbcK4tGTGmNuC5jGdyZXU5ZZJD6fewuzhn/oRxPSrDwKbsup3YmHJtkLbcMy3Z
1Yb3HIdxU6rMvuGJY/WkPgjVWbLFHMCTDx9ZckW0uZQyRs+Kc1jxRRPWlq1GZTFNAuTnIyYVqhR9
x1Lq/OkybSLI0LwMSHx+NG5l4gxQekFJ1eye33nzAWTm1iLATPAhtajp7Itd2VCduYOwq/ls0JYh
RB0jqPoVbauAdr3yXXDIjeXzrQY3Vl6bZtBcze+GQV/yOen4ycGhnGLZhW8zw/RNsF1hmpcmw1Bs
RqWUUBUSQDsN1Rfw+hHDKXBLYnXSQqhaGy+5QdPNRlZp6RWo1jsIHv9TCsu2wV29vh+ZANrXiZ1Z
OuqZwDyEXMWUzVdvFKHcrRtMVt1NVhyMadSokYf3gWoEEINiGVFE41EIX3SK9by9uUQjkQXCxPJN
H5qaXs997AxSPwByacM6Q10We9rONWEegU8ctYP9tx+iHSS+YNNmLYjdCpv33r4TCDzhxpdULndh
w0fS3SQ2K93yRFmbrO1a3ERYlC8Uk3l2uQxVSt0guYekZN8GxvyCNz8c2WAoHRnmeWIqmWC4LQjv
vQ22twtHUw8BrqTaLF5Vw3lMiGYLGrJLHP9tBI4LA84bzzUDTOCdkycSsynh9Ykrfmes/3ou5ZQs
+6m42HPRTfY7I8GRbKq0yQUOtmwXV/nm69m9NcrNTepAfL7qhbebZDQWIS5mMm0Aha6TAGXuFBzJ
FD4bjbLTthm5RAeYH/gm9qeQ2ylbtXNmkj8hpaUYUHeDKNA/1IXw6XmmLB0xZs9nJpN2mJwk3Hky
Lnhnz66at5wsgdAxwggVuJqZP9E52aFqjJZ5a37fdAVGbFHUKsFXYsYxWqfEkMEobEoS+hz9lH8i
8W4Q8HjBRuO8EkeWiP/B2Sr2MO6jFPB2tnAnF8+JgNLNpLqYm96hKRlQ5QjtxQRGzYwfDbNh2Ioi
6GtL7xQdnNp0dS4oZOaAG+Veu3pbQ4fJKKLKMTvisfhCowLpsTjjfpkRNI2MeAABBkDMJswU3J7w
Zzl1cwds0WeEQgTkntU82GkJfPGYQEI9BOF6iMCOc4KDyMCTGd1lcDHKycwsacB8thkzBr1+0b8Z
rx+4swPCxdxVAzK2q5YlEaVWJGTquxQuORxCANG8qucX2Fx+RvMH4anqNMG8bks936uRkzPloT18
XSoJ4sUTZ6DBDM1PT5nIstSHQQM9tmB2HJGv9Dt15EW89/reCFwHuY7F0lLgyS+9uLbiXTJzcwO3
HtTENF2YlDUAmwegeEkkd//ojNeMdKSFT7KtBBPf0EzSM56ICtCaY83i8ayNOEHq2J/jpPv+BRh9
kWiHLTsm1sh6Go7Pnse+yVuS4klWPUGMoh9m3raFxPfL1ExU2NPfvl6PPo11/vZysPMiSvuGIHCq
+q99rusgNNje4vdFaZedeyMjTNWHyl9CCFH3sw8g4ytqoHN/gHPAJ20USTzG1nJv6YUR7n5l/iNh
aLj1QbHYvUNiqdRqnHdCqM/1jgkNgh5lKElBW0FunnVMBftGtazjNxtOjNJbVktvvhBFoTxvkY+c
b5vdeblOa3kIkQygNkICUadR7Z0f2yQyrLDq0/yJUxKdZ1Bpw/cD7pGaqwUF6nZ5KXG1ERhF49ea
/zHvi+R6eK2meC3A75PIgXvhZ+hUpWjq5sMkRxY3IH1eSOFz76GZs8EaZaBcLAtUuJlqXIywDwhB
4RAdougXmQFS2qPWogFNrQg/Nf0nw2THR8oMPWxG8eH5QtFUg/lORFbriH2HO/TNR7RtwNJzboed
FzzyPy3IPmMrpzAG5AhhcM9LV/stE9W10yEBx8DNG87KbNeLvrIbrOsJcGimkEiA0YuuECTzaEDw
5bJZSTUK07FC6pYjCB2/v7atugCkurwQyQwlTdqgKsnbuCfyviSgY95JwJoP9SvzXIxTDdOBk5S4
obX/UnbRHw5WDh8boXjUlycr7z+TG/JkmtUFvbnWCM83XIV3QEbw1Xq6EjVepVROZ01xqVwreHa+
zHG1t6eye2jHzE9GIk6b1uLZ6ICU6JSkWJY5JwQgp08iYIOonER6einWdoVeZwRUlbOb7PKEJrNW
D/0+egrorwG4pjmZOQ7G15jTkEL7uKsWOy3Zu6Mn8IsAgpDjnAMRvGQhVNa4LPP7ajstIrgSdkO3
H2g2SLpg9RMdmq/IFDbH4lBoHEUQC07FG7imVu19kG3wf7uf7Rb71t3fHHx7mt68txDaQ5Kt/wtS
AkKvxvXf6oMenY2xyQWN/Ma58SCI0WyfzKHgsafTm372l8tCXG0PBk4fi3RdZrrz80a+Y8RWrnFz
xE8muro7Z1EZebp8hkBLsV6ikHGgrbqM4qr1hVx+2H8PSiKPeeKCIVxYEhPoVPzj+OMPlTukU78N
jmea+GHQIZ2BePHWtwJo3NqTsuQqBOkGn45rVIdL3MgzUbCzZoFxRIff1Ofw4gvGP4a54f3YTRok
HmBm3bAuXErvB2zE2RNk4ItDrauiVljjOit7KRGQ1DdHKUPRjsFqrss353uQnbn4Hj04zyTMNd1m
oCKJb814Fy+WR2F4DtRLlELSlfiSDpZ5YpDtDc8NwRyMCjTuoDZWfpVbas74dBBYrUmwLmnslFg2
4vJwhNURxj/0WKnQ6GnyXFG7zqT8EwBVRal+/68abpnsOcS+h80QtaOQ5ZFq+dI9bKQItrqK46y+
+7eOihwrbYWq5hffkGf/RgeyAa1veAxk6TxFUKhLqTyZlm2ddAdRqHXcNWTUt2EBOzHjdT2vUfn+
lMkWzIq4hiKCFib25IqbPuS4ZjePjb9/Af5S0PDB0gPOdaG0aDtYW8+yt91m2Q6rxxBqosyNInn3
pzQy/tnb62e6QJmNvZRVssPrmF5leVFf8LVS46X5rduGJSoMxVlmdgjqQN0/xuqgysMKQpHyX/Eq
z2743aH/KGl3Yri1vkR0HvP9mOGNxUCmQmZHwOcnp7zFi/RNxLmyz3oWoHuuQZgT+OL6HKfjJNKq
y9EV7XbDJYrHkuqXH4csOmzdM2EtN5VLKfKRnHglw4SdQM6qjgFj+GIKrbXcd6+TTyF5zUO0RlPP
Unv301p2aQ+t8PzExEwVAKtkdKi3jTjdXIBn5nRBM03CbtX9Q3VXvrRHouucJLxP4YkJMweIUp0a
yG/N/fiW3rtRs6k5uVWUqld1/Z5RVnrbnjp9vQqoTEZybu5Q+LLG++4sc8p8BfUW5NffenLWiGAa
3nGbH6cNXLFBp91wxrqLyQF7u1OrkC7DcO7dxyWXr8Qw3unRjY3Ix2t860Ewu+K4B4HFnr8cDQAp
yUMxULeCfYQybIkGqjELp/HCVvydMZiDGb3orvRSw1/HSe7/dTC5xlSNYzksxkYINJLrltE2F0u6
HaatBwKF2o7/j8NS4U5LN2PuqtO3Zs5bTQ/Ogwi1c7+I+jN2LTCr+Q5urNL6E3HBzSfv6PsT4iS1
cxO0uwB+O+JBhcdf5mP0ixgV54nJ8hW2MGIFlvpFoPcDKxCAwPHWy5hmyBJkhME4OY/LVe914hKB
FJv9UUc6oaZvS4lAxK7o5ZUePtxLEtF3cbXnqukKOUVTos753HVYegA0cv/z2AX8KHu+6DqDuw1U
Cx8oXEnoeNoZZLvuL+AQoKqDSQnWrhtPAAEHwffnHsWINgSif0WTNoywpE7HnRDgNnWvc9ELu5xb
x0bD6aIKKzKdQn6QCNL/W0Mpb5sCovaTLte47rVwAfrPg4JA02HEDKq3S7Xkndyj6T1qyj9QXVQ6
uW9uGVRJSoucj22rbozm+WTO69JCxdVoJjmNefv+i/asnmt32OzvacBV4XUaRLm+G4fEvUC2yLH+
7/RGN10t1NsWZleYcaw9jWGHQ0bbiuGSq6OMlKp9Yri+7Lq+sEqj+AkZAvvhAS0V61tQD2LMfYhB
qgZ9Y9C4JwA03JnecN76teS8HN1oV1Mj/jwE/fahYczUpxPpjXSHsj0Ehzq4iv0ARMXh+r3x4Vp7
AA26UsgHnfIf8Ia9p4x1H8Fr921HoJw4hgLQAO5AFh6MJ8GVmOc4XrE/J6BQDc9JF5piM8dw2DbG
SD+KvGjaH99MK0j7b5p8P+iXU2KasoOLTj8IbYcK/1gQdQem7GkwHlN/r1MiH6ZRs/5y272lgp8J
3XQlGvlrJr7sDlEChHIq9FHQ7QbIDxhH2zJ/aIX3c6SdbULRlUYUnerPLYR3ybu16F4+EtiMmk5q
ZYoC1TFo5vqWuTBmfB80TO4o/CM0yBd58XzKhSlqhbhiFNzwTyiL1IIsK99imDmJGsLCWO4zEL0Z
limceYKjCIM657nUWStDpmyQPbzYpzd1n6SmnJ1rpg12MJ0lO3bXB7KasxfSW1OOt7ChGHXRuqY0
paH8fti53gxSXn1NSVER3bU111Fov0oIWqK4BMwyMFdvetHGncWEbQPdJhiJwP80InDOroYroKR/
UPzrI5rZ16h3jLNQ9D8NHUsXP+EKC1YatFH27LHCdqPKQfOQ6owyExXtg+n1A0FcUavUydmzDeDI
JK/hKKHauwyQrc9rcvKC3XfjPoTdzWHH6sTQhVv9T4J7ykaRepYOy11168sm5DPh66iW/5xG998f
wZ2MKj6MMOCN16MnS7Ew51FddWjMLOfBBoYsYlaLi10//v5+pyPjaE/Et+98pwW+ZTTk5OZ/LhrQ
qvVuebT+dTx8TrQjkNTpjeYYSc8rqb6QGEzFCwlFVz8B3S1gosKCbxgu0jNJTE3+OMgNCjycFb+/
jQwTWMHxzYkkT4l68yxxEq6k66vigBdBYglEsmECcMCSDVVaFGfw45rQ5D/gzBmp6xzqSGcgFkhS
Vx9vheifxXo7qJpsFTFVHLX2BcW00Xxe93o9Y7bsiRGyed64SVGDWD1EB9BwY9EJacZ/q7yhkE/i
nuNNRfGgTQHt2TNJSWiwFt7nerjEmBHI+EfcXG/jNY5FERm2qlNnLJ0TGxflE8XzcRLRGaSxbyBn
fjVjtgiwQ1H9fKsCrTxkKPtwI+kMLKp+XzxVj94Tn3bXRuHiiTyXcF/Koox593EBjq6gtxsGtLZu
LoPLu0nfETFPjJqaSQQoTeloGLBMe9XwOr1mgG348AHro6uHH2Cto2o3buC3lReT3tSa5j4zsIYQ
pEAz+xJRXeUXfLESa5ZnIq/dNf/uGbtAbmcEpSmV06+CdOLnxsM/9zPO4NTwBWoj+dxt14K0g9IX
RWG5H3Cq1tM2JgOWO6Amut3uJPTdC2uqELyG+Szw7wlcBOh1UER9ABioN0MsrUmV/tAwGTma3Qw5
8d7Ph8ETBVyZwLmgSRJxJHDdfVZWRf3UfhHSlYKW0YY6miOFuR8g1//TOJ7Ap/T67WsNly7xFyKS
SI0Zg7ohV0wHNPaYHMAwLrzfKhO7DLBkekuRv0f7xf/BMvlXAJPjc+F8mNjau2vji9m+phEHoZsD
jz04eBLEoFg/FuNiX7J311z9Gajv9YUnoo0oXci8okEebyGf4SENR+C5/VNnosDyJsP5Ww/yZzML
GEx8XbZ8X1+vjCvCw18yMzLtZpNqIFVfkjRTz3owNecoERhGg2xBVlwyGFGrW1wpL7EIU73Qic8N
DDYMgAs1YYuWAtg0Rl9Mi/7P4bjHqevqfRSmtQ8XFmKI4+CguOwXeEXUR2eRUSzGbDG9wBOh6Srp
wmhuhPqw+/IfCx+AUK+O3qOj2d3A9j01qzZSgXMS/SiCSjUnJcewuqmgH6wuyfRv3ZtvZpwccBeF
+EtCZ9EfhBvSlFHtZVEZ2C5sIGTgYw85fiiPqZ/QRVn56BzerTEOnse788YuJ/bh4+AFQeUXpQmi
eJR0Z26F5XpEvfI5igHpHg/xc8xO+RDbkbAT0pWkZfzbXlQsN6R14sXEHbZ6lyHn04r/HWApOyf8
cZyL0Y3Qgeno47AkVRxVIamjCTBal/Th4NnXi/8ujGHFJsNEOUruBAHKisWuWwq2rQglCBSA1Xb2
kR/d3ZYkMGv+sRJwGxY2r/7fINXDKYfB7yZSKXHNMzS9L5/B/MpV2ro0KRfgMVxz4l6v6BAoyCaJ
8SIj5LZ2M9SYmo0QnQCbGjUhREnpSI1s6+Bah7idXdBDyvYOepBWifvL7RmVuGCoCVPtNU8GWKJY
2k+9lna3811NQCP1v8qcsVfJ5qQmE43osEg0pIHqn9t4iDnpi8XRIMyQ3upb7Ha6GmJKie/iRof7
m7kM0W7gfqug7th4JOiSNYqaldiIRQmkcDCM2NUC66b12UadDboZdKGXiuXIy2vyrcR5VZdH5F3I
BSloL+Xp611quZgtQuuVWt1TFVFPD19wQAA/DjClrvjLdnEDtW/gJX7MIhrdvV2LL6tE2jgpdgWJ
P9UHaDmuwZMGLiX4MEGicizDatG41+RvzFUZWgDVY5GldSAl8v7nLEn1/XSGfEs8nBp3f6+t2p3l
0qpN+sqUqKQBDHR+mvzTcku5j5CCe3StkBRFuXel4gdGLdLzoHKw/Jm3sFg2xcvkLtHGiVNbutEY
hbulxKR/4OzF1AELlhXl6g49NXYgdwOGtT6MtZclCRdMfDPuxlWPPZbLc7FvOnAdTwOApTQePcMC
gVvk1uh3EVbt9ZwsR3Ab4wxIRTwa0bDtdhjdiNlqvUz7MxVTar6ic9L7mY9lZUClmFYv5/D0s6cp
D4DEss8piQPevqUOhCMZhFKdEGtxLDu7rINwAbKDcNvfvRZJbt+Qp/HbwrLht6YiHbTt4LDf7qKJ
+4bejN0cG66YSFq3vt2dRSr3gMTFZLJSsD9wlUmgbPuL2dCTadQd2bRkALWCSIMTo+nSH2Crhk6e
9jVy/Jc3bwzWcg98+501DJ73Uc2pKJcMU26TlsUDaDbLzua9OOLuRr9AiB5oDqFY+05ZZi0bkitG
IVBLkfdMIe1zOBD8pgWXZZYfI093OKtUAwrHYOeoQrMwZ+TvKyyLkm1NTr1JbfCww4VaIMiH6Gb0
UOnsLXLSNR6YKAYHv6+Xg2ZPup5B9UzY5fjIxmX8nnSyhKR/YzwLTZdMczJdLAip4yKa0kPSYN9j
HWLNgHyoIz3wAUiGrUcLhvWCtyyym/nidp844vgJ2h95Yhi6L9aKpF+pRgrq6C9gn86gmyn/cEAP
MZZTMR2HFbevScN4ZSCmn3oDR3Durb/6P2TyfVh1m1lvWq5PqxpF/vGUu4fr0B9JR1w3tt2AIhpH
M1rh5kicYgINxB4uv+V3OOLc4Qjmd+4P6GgvoD7tg/LnrOVW3PZAnOFODVxmG+I1anwzz2sS2hu6
+doehAjlirqQM+iuwct004bf7jMZGw+duMc6+35a6h5rek3w/EHUb+j73ZU9Ab8iTConh+qvVjwo
xoi7W+uwNhN97phR2i4A930YW00PE77Jb7LaQgD/AgMyiTVe++pdFLrhTWhnKfMx7Yplb/3itAHH
TJAJgtdGpRWKa4V2HTKRfKb5CMlCJxDwj54L8yhtHVtjLKlG/yngQgg/bT+U9UEG5MWwSYFyu7rX
wnnqSkVAXhJfJco8zDqhzP0K6GgJ1Dho914CFRhPNTT4dCbZB9AN4Gd8EDUCr845eTVSkwE/npm9
I5hxFE1ma7ZqEglmsvnYLOK6FEg8v2jyyVapn0bRjiUVqkmA5LAIlC0Cg9k62pXHvfyUWIxJy3aK
2W5qkTRxqeMbR86cHu7fMrvzg+JwRwX5U6t3gKnN4kJ8hfvRrbB99K+o3Egxn0jGY8DLfLbw627i
/AsDpOPdTswlx2HVPvqAWamzICN+6BBcGtDsQd3JYBM6kHwl7UE8qrMblLj3DXfQl9vd+yfmmGnE
+DIS69UDkBJrI3QpHEmxBWH2lEdPQyrk9SMlhlaivVr/ifKIWGASPQfigmwDEQpAzLNkff1j3PSN
ZwfMcCKYDJ/zr+v/cgtILKosw7UGeF1LwNPRsrefQS0lhbfmff9IIbPvvBnRFQj/WxXurTsJ6zmK
AaedtWJmmGOaBZiTu38YdRaBUGWgXOPeI5/vvRCTJWghQyIyLSxBiveUnb0iDhF67mn14gKDytcK
cm0jHWIRkD/8PBANu4S8P7QLiqKWNbuXPIlMTsZTd6OPfQhCFgA3oTHrk55B9JVtvu8ztPZyEX3S
6wxzKMJ9PdU9CL3Dn9nZI2c49eL63+JHa2UeDhlG1xXsBlmrmvaCblNqPdo1k17sAKZkopl2VRT/
NkVhAQbD+4aL+FlnoIW1W2/7/5z1QBtbQCAwZ3INIE2DfDutLAUw44JjVcShUMCa5sk6ejcGhZ2K
66Q2IOsLrquYk4/U1xrEy9AtCfUSe2NNIREo33s3OzQsp51UO0NNuB29wwVrEU8z1gtWQ3jBT/3G
POEJUGyhs3z/Z/+jenUuIAyQOOgZzhsf/DTKWOD6kHM51804PdF2BLMUIprqcdPtAfst9vGENlb0
8qviIMVT2+MFMa2afhDsaZHJrfnCy1TiQ/iVXCngjUov5UVqHJmJfGME3eL26dl3kaGaeURKAuin
cGUdBzyZP6rmTm1D6S6oFOPPsFIGJ4tJgVBk/GnNqROkZGnssOf6z594fLBNdDJ9hAOCZILqUIPs
G2JZP769sRXOLxo5LzEyesyfywqJsr5lpiuHBFhxc65KNzXhYzO5MMnjZc1k1m81oBnMCFZkmHAd
7qe6Ac42Du+KxqQi62aBr7IyFpfgL+wgAvf3gJmW+C1IRMiIwT83Q32uFn9iE6JqLmzMtABRdWWZ
zB4JK1feg6j5Gk6QGpHVZ6KwYgz5w1FCGLX2V0a1S005hjVuePOWqQXg6V9ZeXsTWDS4UnXekVtx
CtdBe4m95+PqlBNXXW4Yx02uRhAKeom21JtTCVEwPvghxfb/y4huYZRNoza/6g3ieM31gNhfYV4R
vh/luAFOD0/m9MwPMWnrgWN8kZPT7T2AUYRwyv6bjSKrgFDVKD9rL/lWGALe+CycnToCJkLJQP8G
bg010YfIQ1v2GoNxGn+k6zMzCpxLUQaB1qPWt/Bn14+1LsHmWhQ11ADkb9qoziREGjES98iEjQQU
b3vdUzwcnFX/FXZ9rBcr+IuDP5rciFTI3ut1Ex5h/8UjksskN3LXaFeOPJeIXCkwvGI6NJznhMB1
FdnaniSSgH5Lf05nsDFfWFyXJv+FFuluZ8ob3Q/m807ELsQEdyOMnKpopGPdnzonSZbHN9uZTbRB
9Ngl+gINMzbDb0r3cSiJ4wWYwAGGlFI0rXP48Cbgp6rvev+4ZtyTDcXdXNNJC7BiO62HnyY2XKwm
kkSDh4lrjed1ylE+ns5wgbVn4AfKYPBjqapaTNPqgKOXulQwgTMovUE/w2+rO8mEJwCBJO5jMf0T
OiHLye4mmMUtXIb4MPMMHf7IMiggRQGGh+3tdGIsKXVOUYPUub59wTKsj/UN9yWepJZd5J2eDMeX
u7RHwKoLPZQ6XWcELEkZMmg9K3cF0tUJ4umhYcS7XrSvZtCfXnJHrcOvI2pNNrTmYTHBd5L3HsyY
EhDJiZCSx71RgxQD4yR4+U0qJq22Q9mxGAYhMnVD7DcZA5mV+/25pxYaBg1KnI6IbR6ICv00c1Ue
DLkFJAVCYX7GNSlllmjPvyJcFnDPRTfW1YZw9HUl3G6SLvOjKkSGQ9HPdJz/oCL8B/H9nSsWU2kK
JvMguNU/7YO1Z8yoI8NwfyFGvHdDbppog4tw/0hXxKbtaAaN8IAHtnpGNvqz/fIoCeMK9KfBVMM2
5OAia8P7+C866CRYgH+bkPJEAK9jGG51+cgcM320tP8ST0ia1pVfsoWgLuC9CYzaT4HkaVJiphZD
K5/rmzVbksIPtFz4BkzvB5/sPgmiSuojySIZV0NYNTsQzVotoM27tz3CZvmhzoHSUK8qeCSAWNaI
mIeLxDO4dckGQBQ4B82kGhjQv2yS59JTB1wd4I7fstNYjH9Bp2pzugw4GIhifMG8OCgzhadUcXer
OgkZbTz19aIYe+TIPFUrnckAhrbUuJ/YBIRYzGVw4m+Yv0TbuweDkt4G3/bShz2qKZmgTS91MgWi
vIqRF0KvG7ajIpIpb7r4680ZQixKcjQ8/cO8c3LI/fX1SoXv1Uii4jnR/zmwpFjt0LASRvM73kXN
hWcEBCvDRBpMnC9ZEFm4Dm8WmuQej3DB/fUvrA0aS+wc0upX0+yXpQACOI5QxEycl3JcDlQcv4On
EPFEzxw8TEnjnFKy5XoPVDxFOWATxxmH4VKJRr933UyPfMRm/ObbGNCPSo0+M6VHxDKE/cdOSG2l
22ShZADaPAKpVYzmZTztwTfrwrvYBj7K0Zh/RN13GF7o4L1u1V79BtHEVnaTuB7x7T4v0I87GLtk
8EJ0Mq/O6OQFS0EBP+1QWuovYhYFBp7VQMQvisAkLWj9Um59jcRzPINdUSql+K7EXBpCOf5OtczZ
rDjulluknpqLm3J2Z9i4jP3CXuDzomxPTocsrVckYpDox5+V8Qe9jfaFMv5ZWPirv/4/TaUFrjun
GKiuu5uq1J3quys5K7hN37R9r8robCk52aS4MRDe/IO7WsSV28lVt1QPP5hvpfHM16vhn4yJ6YKw
V1ALA+Bsjb9DVqkjnl2Q11+/pFuEbzsGnZhd9SHA4kCd7S5ign/ILCKcqvtX2ViV4Fo12xy3Lef8
YEHRxnBJsNYiPBUhFw0Jc3L1AmSNuAnPKBkzdBtCX9WAK0IrIgS+WxH96YdwTsEV4ly3q/QCtETZ
TDQqI2ABW8cBtP9bxr3UgdM61XOKTIPjhk2VbuWako3bmZPvM0BmHEFTOCEqr5dmgutRr4zxcqgH
tNHSPRYrThjKrmO3vM2gHnp/ft3ff4mvWKIKxzOy6ogXWN46hIksxGRyXWWQRpBXnmQp2Gc8YOFj
pVncZhUmpgYZ3MQNqO315AMCqDPZnFs4prIZr21NhvGZvnHyrsF4ewFID22mVOek2JM0YXI5iF6T
zYGQPX6GpI3dUZgh0uy4KisEaYqmuIsluOBxNY27AISZemwFoek7yQlKLchMSZ50QFPiUrbDgzx0
3xU34iZYMEp70cH/qggC8AfiV2WU221l32RAlMkwgkV0OfwkA1u6sHMQdsVl4furaRp5kjcLdUJk
9dJ2ssOLTzdZLBpqaCPQG06n/C+2FEsjVemWOwZqOJg9pkFvxGzj9d9yA6qu/iPodpaNcTUZSKoT
T6KbvXwUQzXg/TFA8qmBC0tv4I+TnBEQvYX00NaxMg8ZGTCgVVlwQ7Tyz7au/lVa5WF3n3Udnlm6
F9NCXcSvfcWYgENlrphTUeXBIHiGq99sxlfqIPWreFWA9TOaADAeSIKjXiSUz02SDiFyFKPSWi8C
FfkJVbQxXK5hV3CD/jRu4u23wklU9slZY8QGnYHkOyIGHQRnN6vPCvia6VpHRJ6X1Aje3chbVMIL
W7YMnCrtFXPfMWSF+eMhTtgGfqZpXtEdUv3ij0TM6slsgjcL4pe/N8K+mW2wGG8pHaXEbfOkfZac
+ZnIBwgt4UYdpYM6ZT1kcd1l6ThP3MAj02/PLbyn33DgJQ9KkwiZlmTYAgBmIk3mxFBYdNuC44ww
ZOH65eXGmnTCw5fqZ8IncUak7dtIqXcRvhxTlqQaHUohXn1nkMdQxfxOxuyDTZ+OF8WN6bu7wK5L
eic6FzDFpXP4EopAL///jlMOXjA4FrnafDktrCNLrmn0gsppB87/ScXlk8TvK0wq4au+IiqgG5P/
7hfDg5s3hhV3bVrZ9aoqvZymwUI59TRMg2jsxQR7w7aHkEPidMHspBMytgsFXWoLovozWqroqy6B
jvEVD7O98SEW8fCoxeos64yUXczl8BXxTzuR2buVhotMvKh6B6zATKu6BlEhga2OUtlFhlQOBkTd
L0rtLL9neBLgb4XSIzCaoMkS4yUlx/XBEMJ4kcrqhdw6FqCtenuUAPUc+zecfG2ObeMz394g1EQP
cFLt3CXllPfXFMW1BY0+k2QgR3GaahxjJRiHAifxcmVEElIhGrxCy6GB6XXX6NJm5+UOaVoNyyTJ
IioqJLJJjJMvQqP0JCj100bUlV+Tj8JaPbwecz3NdMtp8Ts0RQZ2Xe2cal/pLRQhdUFR5UK9e5lX
+rdl+qGNMFmVkMEplEI1XV9GWlRGlOnOnDrZY3+AHMuzZ1s/MiRtL2UbcF2M5Gyh2Yh7tiA80ERO
dAxuIsazI2t3OP6xaPBegiZxCh2oOAfAe2WiOLg701tyx5TzU/84TDLc07JUYC9SumqOIcT9Egcz
63+F3os6LFZGmOOAf0HQB8YHI1Jxu1IlgayeLCgNZldaVVKvTZaol0F4dOcIxIdyp13O3Tb2a/ND
B2pmsO12qeKSw2icQ5PtYwE0lCvcgsFJrXJQl5LNoNTCBz6hvqQHPk5Uk6XwGxnVyLo+F7/sIvnw
+iIWHxE9rgtcN79n6OP4dH/fvLTna4gTxEAIFb8ZKjFI+v8jGn/PV7RgCTrTMs5UDEDgV4LFK2vj
pfFB13mwrwqddOhAUjdIWLVfqxkH4JQWJ84Er3c7xmqFyygTR/Tljj3amnVtOHArqzQqueN2ci8f
mxLibPk4mhJP5GFETRjjSReZ1hEM0raMGvUTjvq/oDUbVYyFvVQ9O0fQTiCFJ1AayJ8p/Oqq9SmE
sbOqrpPaOVqGY3dU9lsiHWUuv91S8wm2fNQlc0XIfOCh0NbEiX2dy1NavRe6jt6fOdyJD8Frq5aN
3dbbvbJcgE0I7It8HpHZqGS48oL+6W7hpqI7uBQYgcu1Ph+5rdUmPFcqWqDOed2+Ly5aOfAllcSd
nQCOfIUMPitrDhdybboGhI+r0AJmb82VBCm7oY9UxmmBWbhDFl7TaSF1BIHszshI2CFaI7JOLK9S
VIOzWxLOMSFDWsBnUFsRhl9q1rXwXavAV86kX3oHlRmuZbOnRI7T5dm9gafTJSzZuw6IlFGqcJly
O8+kgr14PY+Mwd0U3y7+T7XPJVqj+Jbi2WoAMRt8z17F25pRr2OuKLB8I/7XIOCvw6qHre9FX9xH
m7vCFjJZZdT/sSa7Gueej1q/+Sq0nUfGYr/7iFVvy3cpvyRoo43asmm17HspXhTA5lT3lsYaa9kM
pFk+COXAYz3ELVbDWMP10RxNQI7r+rBj4ulbKdGgTzGiz6aFNCpG5JIhnepjDVDDlta+jN4NUBYk
2xg1nwRQHCdyCvtvnSAOeUHP3AzvvcVTiMhmpYiOX3apbyo46czge5z50bQHN/N4h0DfpZi2k/tO
u30BRk1RtWQ6kkgO1GjdD9/2jtx82RSgABYmtWMYo+NjiHiUdQ3f63/eXVh0bVf5XKyJkCGPjNIW
mGh2E49N7+uq6owkJr9vPDGZsKjriTT7yoLs2LQeDHLPVIPRFFKvCyct6By8zFqhb+Agi5KdcV2q
n+9+K29rxI517x8bNeVHnPzzOat4mytv/jI1N4F3g2f6061FBa5UoVfiAAWKlX+fqc/WYF5lsPQS
PKj+bcj2IV8/ZtUcOs9jwHGAZ+CONuTYlhvLbVrB8XSH7Pe+T0EbDm722j3JwuCnmMcTzEdgVfVb
3wd4RvNap7kOHmm1EBGLQKhqDt0QaKpqjvAA+fgN9Y2GfKn0ZlchpbkqwuY75HbQygjOqhq4Cf9s
JIO2cZGfbehzJJVlpcbUux//jEXv7X7kh62Xq8lAfM8J89cQ1H84n5GjDmttwAAKoI4bpGNxCk3D
5IpinPVyfach6lJpc0F3WX5QElL1Aj2IG+lf0mwUGYACuyEkh0SqgNuF0a4Zb/yI8AUEuxW3C3e1
kZcgRwZoza9YynpAwhBWgK/r4su95zDycVJKJX2lGv/0mrCDPSVZ2B/e8fA8A+kq29OnPdhUZWXz
ycm0NDswfBExZQLGLGNBgSD9eTc2Vyhf5BaGrKXOfB072ewj7r9oEFSVZF0Cv/QqIu7yG56l+7mS
iSX7SmbN4LhGTD00DiRfgQwD+++8X9dEPgsJbhZf4ejeqRfT2d66IWaZxYranShFQXeu5V168zHR
ZxUQZpfbi+38nhT2YP2MTBMyLzxyN747yi8x/O7AeM31gt7/cWkiFiP6Xvpu7tzMpLZuGKiwpLXa
CvSsWDCjKAnMCQnK7IkHSHOeCR0kqhMMOgvHm9ywxQmc31CtexMxuqTGb5wZySFoQ7H9GcX8GLQ+
1UcKvOySK9AZzpLVgUPHSXPnRaKl3HnXnnu5ogS1f1tvXP1+ebqkteX52tSaFWMI4Fp+eHXhBOdt
KOPadYdwFHlIOwuj0eVaz+QmIrSLU3b7SBT7GG5NG6WTVK8+uWgIJWuTxq2mVttW6bhcp6aL1k+Q
EtjBWJbhE6dtFhUzQp7ZreN+8aYFkQxHB/hdLw+SkyYO9t3EEca0xMtX3om6O4ZxeU18f1MhfWSl
888AgulRaS9W8/+tSUjSm/oG8yBQVIFdbmPPiN2M6PeUb/C6kY42gKDUUgUJACTusfPPcPX7HnDf
iti7QQP8LlVLYkKX+kqIadE0d+d3fzE3ChLYSKxGZNxsa/qEu82aIzTawlDgBTBCN3dhi7ZfYZtl
lscll3kMCliRWx7x0Il75tPj+bR1jy8+mRXCD+iCHVGtAkJosUaKUry5RdasWW3FfPsjCthAxdvW
E7eM84PLsBqCanLZG/WKzVUwMVSs2FVgNyi5FWYWPqyLB+uNfaDrmoEFB3Dfx7l+WTyZFJf5Ev2y
SmJQnKr6Eh6g0kMsG/HUfw7bKchWJJP8qLxmrXHGeVjvNpMRn+LKnu/7BfZ1PySE4IJFNaPTDMiw
n+/eWpooi19wRy6av3VF8myNhzLNkwkffxZI83cTWjGJQmn+NISDJI40YNpmijzhdUMN5FssE8Gf
6YnGd848jYdh87JWEz2QKBeNiioz3bGygXcQW8M0yfeo9zncb9TXlU1QMjuwSYt5QPCmPLx7LjBh
1fwRqWMIGWrdUasNnnB5eTmiL8YXD8UZFUtslLUTRit10drekbtmfBykalG2d9cryPlRzNDjIvNK
9xB3s1tJ7BHYahh8EB85H9VbxAIHz2eYK07idvS9PQyNYuMjaDNdev1t2qSqrKmje3qi3UchqS7e
l+gN1yls55ZgIM1maN26QQ50vELuC36DQVLjukUaO6FdzcaHRmqoJaZMgMYhu5bwiTO6sZvKubuz
d/a9CXb1KggCDWv7b43DjrDvSD2FG9h1CfvXDLGw0+/rdktGEaBIXebg+FRhAZD7w46bFGGUUWGf
XzYw40BqiP3iM/ZJri9Xlgo7zwxtqwrZUxm/zhUZfk1hJJHm+z7Alo1xRpgTqkOue+IcV6ntHZ2u
PrsVrFzg8uOAaszmn+yi0yJxNT3joS+0/+czOmzrEsYLDsUf3MvQ/i02quzYilVEFHTsaOakzmPL
3F9wmVsIny8xGnE6kRtfTfpfoMAGqvRSmF9++wQ6lv36xF3mw77oZPRjv+Tbh8sCwvDS8wERCtFI
PPJFsdPNIL9TkEam7JXenZRWny5Ghj7VyrEi3w0eAKBHCv+GZ6+DJaIsIPWj3oliK96stQGuD3Nz
5NZaMSzAybHn/HWxkOLuECf7YvL7lgMcbkZV+gSHqaI1UtYsg9wmtNhTbiDFdXB6EVJ8jxG+/AA1
EXI6TS8IQSkxsRrDwDn5t2Ef/xG6AeRS7sPvRqSRZNNgCyUka44OkG0kiwJxBm1hM3Umpuihs8jO
R1S5cq6JHc/vnbPQxxe4uBrHOV1OXMN42FhcEob5iE48Tk3dM+lDsNwNqkI7aINdBWKB+chRAZlq
p+ITsyYTsZjEIuI1ElEmzkCoAMfJEZw1xuRQlx7uReO9eSp2xPyma7moCXtCVTvuzP3ESi4hSB9K
BimHZMWaeBRqM9/mTJf9ocxPhDR5sDQXwTe0oIlkjOGEbYvVcQ6K9B4p3TzVjnznWRXZY1T0KAfW
NIj+ykXQhJTlDkXpf/992FrAxK3L4w69pl/fsU9Qhm2iR13jjt/ukCpLSYAyadpzdadOMBG+h6Iw
VrTH6DLTLgHpOT+0xrJlS1s3ldx0wx/ff8zuV/WwqCF9aWLS9Z7bpYrkM9YwR+o+5mDIh5+bbude
3JGg4tpyI2U/t7qCit0lLGANxC+plMRnSsoM8KtVbwtQuyHhluxOWpzdCJt/czJeCjm24A1t+c/p
BOKraMKNur4WyYtlyUDu/TI5q5cB3yMxBP2erzC51pLQ9t0b9s5uN5DLFisPsRB3QhTxrdL6vHkc
meuS15l2lISkax6veY4cUAt1MxV5t9Q5nuDAkmrhUaT6XwB47+wbqSvb5z8E/hPWJsO1cg4yoqUu
4e/HqELy3RtPUkGaXBDsd2/BS+B7ikV+o3TYU5ZuElvZjwuMlZG60Zclg7/SJtZy2Wlh90m1pHIR
0EGIPLyur2bj9+2SqPnXC24ZWnZM3yxOTJncpEwTvbUnmlDPVGhcCQy4WcaMDiiTalwpcezlXN/n
tr1URmjIWmsar4E1N8D4Yxa/9GVaOXC/uGoz0xFvu14oRYJrAh4RurxweOkJwkiowQM49jTteFuY
bGZxcd3NqHnWFZO4Yb5PSGM2g3mV8uE4GXD3VFTzQEUmOMFZKxXs9Ner0gr1HeQ11YEYkEfu6cDT
fSI0Dhe36ZJL2migySUY5CsL9g66g3ne6Gn1nP+lGh8aOtzdoZSxCj/sVK/umk2/bCP+mfNfjr5n
HpWF1xtiZZtBc+oLgNtysCuvexo/m1gmCHY283T9wxHNa5n2DT1qKjfjpvgJVwByKoASLtEdK/td
hoGFVFY7KlWUGvBDo6Ih0gd9XhdFC9nZGaVyAZeeCFdoQu2c/KSoX2JcKcSo6eEtTNJmuj+R90RD
axLGbEIoyk0qu6BVgTCpl0ggGCqwJ3B8vqHHT/DHW0Qqi9QMoGWQBMsKXig2Uebex88taZlJjt4n
/y/vOIUIlJrFxf2Dp3GgtC3xn/V+H7XXY39Xqmsj13lzNznmALD5QCKuzgdILvS9xTcO9uWHtPvE
XeHI69LL8n21pbfWflN7thb7dVCf6aYpQ4aAp0qQAZBJYJS8uo+rxLrjcWc2PMv9ttPlbZxwhXE4
jqKREtsrPQ7EVlr0HlPs8ivpcBSBg55hfdJp/bFpZHZDbvNTviU3ftnZpeGS01quZ2GQwOXHg2GA
Si+z/49dhEvlna/6Xn39BGqBMPcGsi0OQw2y2OeoI+yiJqUcseyBwka0Uk6P07sA2QHM1YR9Ar99
+UMVDYd3VwmZbfrjfxF+2aBa/i0rm9J+ge5M3f78RI8IBmdEs0Kwgz0WaeUuP66xutmWRaPpI13W
8XaX1KvHjNpL8Htu2l+j4i5u6jepygahBpx/spzysdWxUhcHgaSIgMSW5hyVX7XgGWnm5dxboS7e
bHur1L3yF3vHzNo7Mz01Xm8vUQ3SFXTpbAKemgWk3uODb/LYToAlsHhbinYjFsNZkIvI85RQmaaB
0PRkkLk1ghl1FGGiAUqN5AaEKiwzmXQl+ebhi6oyBlfp0FbR/bbkZTOzKNmNahG70wwAommZfqaa
JHYdKZaD+FJblh6ZwOQJ6Ao4WIH1ebz8KTHSH508uppcYakzUFSgVRcNsIeC6rAfkg15wsSQOa3n
1kOXBCHqXr20i6yl1gMqZfZnHOHhqMYR4Z88bD3Tdg+M1/MqzjRjUPr6Gw1kDbkpD0d1BYZrnwRd
FOG0S9rk0bLCkJF191eZioMtlULHyL3LjGDROQWWwFjB6yBhr/GFnwKdMGMUNqF0+T6f8LOS2yIB
o6NS7Xu/aj2wrOD+5BDbSp9iAQw7/fdvuadOnwBvf0kC0h6N1Y9iT6XSUyMkC7vJy80FKlwP/kns
CP4CvO/074YYUkVPNRgPoslPhScR11ZUed822jM2DZi16EtArkb9PpkkRu4Ayn85ZJcOA6/Bavy2
EYHFNgC6JCgZ8+ytmMSAh3Fe9+HI2dxLueJwMAOrO8U6ikGDc4//zt+BWNg9IzdTwfD+sFzybV4E
BIxksPQUUfflIlDe21u/QqCMOIxDphQCadV+4r+lpOfgMaJyJUMF2KFDvlcfbH9lYzq8AbfFW3GV
uqor5AArY1pQt+nXvgkp4/BuAbR7c4oEZkDrnDMOUywFSMUJaGrxMsJlUWlj9LAyaXtxINpLwS4N
VOuz0S5gTlZwdiaEgGoaDxeNwoIJoRsSz3c0INaAQURo7RDYQeaJC3xRVoc344gk1L6JEVrvkHsC
qEpsvE03CRCJ4SLfxNVAO72JumVMnu97tVvm6NajKfrby8iCeRLRST8NFkLuynXrXQX1XrKDoAhV
ZcMbWNBUM7jm5QcwuJNjQY80w8rJgonsdq6Xqt9mggNHSOHOnX7qqvmggkZ/wCQEWrtt0tIX6M7+
0DPCVNkj4REW6rECHhymcgGaLAhgc9Ocr+qNpSBlwUiz3aw4enHugdP0eul33WhlsF0IlmYnuUav
Gc6txZ6qOMVAYoUvqpDxk5D7ED+Y3slIDE6SG5PtjXedTDSvUxVKPjoIYSm567QrjNjD/fkMd2zC
UqG8bBLnv9Kf7BAfeGWeIdEMTF7R+RYxz0nZ82RUaVsu3F1suT9Bxt0PnWcH/f7SbUL14++72bcS
MiQ9IStxjgQDK09ucB/Lha/mmiqtW9BcNTi63jkQuzrogIplW219Ka4QFRi6PJiJ43QhqeFh+zE9
LiffS95Iwjv4LHCci+Een6Y6222Dd426f7YzGToNuUmqrYtmKIU6/gJxWbr9zyEw0ODS8oqFaaiT
+peklj6/dtA4enDxJrFUY5UyvTO866MHpoFwCBvi9UJVmWSdyrMCVW91vXu7T+GpJn0xH6sDGhTP
F4DR+Zqo4JhjvAUxyjKBTP8MUcqcTpEln0HDhNee0qPJ1G6+eaWGhu8p7t/LO1cy08VcA6xruDkL
78Wu5fyeCuG+Vd+2eVcJ83JxPX3u48YVZ34JqNdOHPGJcOMfIC4q+B5TOKCiJCh9Ci3Dy9FGt4mS
1xDnPpVCqLUHBCvfP+Yn8L3k/udW8SQBOfclnVe+hXim3DHribdPPiYcrbOvYRAOsamCBkP7NUsi
qZUCwQPrnFe0cgnzcxTSwjQH8kE6Wj7YUHfj+m264qprJAvuXDiW4qE7fW6pxK96+dqvzRWSMuic
eYQTeUSlQOJkVc0gwpmy3O+No+RqglAs3Np9ZrILHhK3/TdqYAio7DNp04sfEjfvpOpq4U3b0Ejy
cODIP+ala0U92SrYGv2J+g6H3wJ2cmPoYbzCUYaogaNkmI+pVdnVxVC5LLVHmDUs4vy1Fnz74IEv
6o9V7+GcKuJh/NKTWl2azbHkUc743HFOhGku9fEw19jgzYhvE+x2GLRS2NY13tb71S2gc9VSvYkd
vDVKeCFmIJXEyRHC92pFMxDHlSZNYqV6Qy4Ig0M+8t8VeWmtCmESqGCvvJzwTjmBYayABYRxwhuJ
he6Jl/RkTF/tnhmyWihrPVIFf9afMFNJNc/09GorFn7qJ39hgXVVMr4bNJHP/tPPyB8qY55gw9v1
/BUm6kXaX++7UeuR/XdaxRZVtfzXQL25SWqfsKZpvibO2ILKzpE0ZlbZLt7SXEES5fRBmt641XrV
MREpuFvuQjiPorCzIVECrOrpfGmDKJhWhrs1XKdqT1W+QQKd8EeW6r0Atw6DUIWtgrZBRUdUwSK3
UfYrVTJ00X603lHUmnnWUTyfpj817K/UERIZyv/hjsJTEwofzYKV/zpFAnQd5eedw+kE0WIq/tKP
5ln1rE27uNzpEsU2/Ba8xgmf7851+yUJ+c0qjNm2LpFStGhTNCYRkaiA/I4fB8ia90Nc0MfjSngV
2yP10oXuuJ6iJKpOy+gXquxsIzhU2hQJWwcEYThOe+99ctga97npvGVQG8waWY52VCt3Qta1GLcq
KBhLPJCSV5ogRH4n2sOiNlsZV/m5G1/u85bJ1CLn1LVTQDHAwtaRH7q2JsMLezNQOxSkAevmiuzY
6I1Sh5jxvdcrMeSSewJ2y6kC41KtD0wZ/2mUgX7ME7+PLPmvfhd8llcD9TJ0oAuOfDEUt4wMLBFo
uYYM4afqr5wimZ0pc+MOKI/QhecpKbxiGBxZ609tTW56V0jGs12Tkvej3Ew9PbVZBOE/zobJ+DXz
oIOZscF8R4KrrL/VxcFWNl7PhwPLLROayN1SisiowoSJ528k6DPWpItw82S5h8yy2BjKwJb08dXp
xEPHWVfGl5GD9PDG+UYH0tJAcxjJxVfBs8CsIIEeeL8qin80ApDbVxaFKBXCpWqb87IJUn2uOh4b
wdK4QQEKzKBkL7VbN3dJKgZvBwyAw76vEFIOzQIOWnUBEpzfR7fTVr8IHY/hVgcwFl+4w0oeCEs8
9ZCz1o6emlRFlAR9j7wxpZ0rXOypp0r0e32ZqoKjbJzjHBXZQROo9LT+wrkQ/oq8+EQWodG8StYU
GMGf4RjkYMDWM08wWr0eGOVlvbur9y9SSdOPO0Sh7/e91ZtX62L7lFQQl92indrLYEPpTbDeHACW
/0zSs1shwHJ1llycZTEmOaPHaKN+0kKbE4rhZzs5zGZR6rvFHUqZgO/uC6Ldx7DnfpVILUlQamLy
HQ+dwLOsofcgLDmPFcKRAxMI7M2D+xVmT6IGKfI7AC+Pu/QYFIcOysLvT5s18TeEUuFK/R4bZfTx
eCv0QzcUgzhp9TkR5xW+q05uxrYGq+86TcRf6eR0WPntfym0q6i4Q7ZmWM4NKJBejZb7fRjuOYOs
5GNubGbeCKLMCFfclgxJLPyvvYEG6vbhCa0NOwICX4MzfZDd6UZTxt4VfoyLDF2eB0AcdfjMw4EK
2wDAGHF8VXUbKrh9UQzoS0Pw6EFZQV3lMUYIUt5VNlsNetqHTromTgg4+mSmMIlfdy9wNiD3zfNf
xoMACbS4Lg7YILEAFSwp9X6N2CY1XF0osul1QxeEg77qNIqIYT4r2plxkT3W/jj5PmPvlKMlOfKF
8oBn2lEURB9jf86M8aOqkj5YttoilnMv9SM2qqm2UEt5exyhj3NJSG1B8W/3endVTlP7xAGzdjzc
P9Lt8vv1wr/cw4bCOjnXkC0RDs+k4DDoR/T3l/4gI4OCevGnMtEYAjB5JhTB6a0DNbk3UI7KcChu
pyoXfGdHovbVlU0BbpnYvuLZdzT5Ewj25v5VU1KbwzGBKXdZ2kmXLTXJoYbhRtVZUFE5qE1HpcFz
OMu0YVOIzXwfvruqXbNU8/p+JBtHkNeOm4m6y83I1jV4TyvYEPVgpLZx3nBuqMrEggGvJvlZefDa
25kj6oKmGChDKzwxVe9UEEpyOPSUQBT5HUM4vCgDwQ/hwv540P0iWfwlHHW7THdNmswb7mWW1AZ2
hpqZ04C9YhoMbCSC7AuFABwI3OKEcTMzF/QN5uXkndG9pITU/26vWu+cG1GhNRWCNAsKjHzdEH2z
vWByd/virrZZs9PAk7P/eqosr+IETSYgZQKtednFj1egkLH5jiQv/8FR5H3FrmwuhHtu8PspaaF4
9ybLdfkQX0Z5I/H8LYhbuJ/tmwvdp14NLB0dPJFFRe52CiOO0h3EYj5Gqnb6PIi+5boeRHBj7NtS
ayVGHWc6MJYOuDDn8pl/x6T4fF/m0iP26bd2iCYtMCfsbBS9er6g0M7HApTvGzwAKD+p4rSYQrOq
KM3o234AmstUSEkCzmvOjkouV0Pne9SAB1o7pUINJA0rMYwi6qg7t+qzNRovjoJ7Kdb0Sd5dITar
HtxqpQlMGXbgHIS6VqafjVqzvLvZxL71R2wafYKtRQHYSsn8UL8MpAz817HsFbwL9NBTJ41MYZX1
vscMR9tqEpPZh3udeMOsZ/mCpJjYsAtEKZLk0nusWLQIqnjattD5nTMVtCCZaHug6jET5v/eqnOd
KT2PmFUcEHs8ToTNpavn6LLIol7hjRs10Q06m/AcidqNjIFCl31JUdTgMAnPrMyMK8ab5/LcBV8z
XnyEqTT4wIpr2993T0eYQtKNJRZ9vguDWHZS69zGz8sRs/5hwsgjX5tcyrnh8nY63+Mvt2x4vtdE
5gl0sFSiFKhr9tl3KPEGTBbPl8bN9csE7B0g1Vb66EgHWtruwwyOv6jSeWRy/3O/u4Gf0xTB/IEa
wB9jkbsnyp0QJK5N1JyclwBMpGspc7Q9C+cTrMcS8YE0U9WDmNMr0Pk2vosGOq8p9yYFsSDcLJ8P
xU4usYLjyNeqzxu9yc6EfOMk0dtg75EMUm86qIJeu5iKYhA1OnQU79HcIoJ1h4IyMiSibSmkHHj9
5IB0hbboVwK6AuYxptF8znJ/G4mAZ4MpokKaVQ9IJ59HOztpXauckEPQb3Nm8odNwHKfjBebpSf3
4TSmhFMPJis0RVok5RvDJpOiBDgmb0YS23pzf0ykRTnrnA71kN7zWWfJeX2jT9TDpNdhHaAc7Fzz
3TK0NzDwdFQJOxyGp6LNsCnvD+hg9cIUXl63UYNfDyK7yjeOAhVbXMEEvd8Y69HkhUdxcifbOYTT
Ek/LGr5GhYcJmrBeBZ4YbyvQDi4PoqdcF6PJxyc8Pi4fBUBFJ6PEqddj9gd1O+46acOOYaBkiOM6
X+CjRCfhods2embYzuWSmGFfz0vtrmyZt6z1dLfmotPMxbEfSpaBwQaezLdUlCM6BnTXDO0u/476
BaUUnMjFTkY6s+rgM03O09i1bNvX0YYn1F1DIidOcA7P1W9VvCQc51eEGC1maNPzt8gWH44IpcfH
E9Le6N5A+B9HbLH7ge+CvRa8r+7T6oV7qumVEmOdqrUBMHafG8vDQtprR02lo57MWpB/GsFEvpWT
gK0scFNhRRbT7VqBmLMamnD7TfX48XmDkrLjwMkgN47cwStm7K6T+I+Ij1GRiZlihy/eDeCsW0PI
KhDvQAB6KwIKewoHc1GlPInlrWQCY3LO9TGeo70wMfSA0Vc7Nkt5TNnsgkMjsxBA6JSWUh7cRyfb
RVfGKm3dQT+jguzUtSgGcHDT2WrOu4R+IE2UISQ5i6elMGJmagV6DapZTJfQbxEwqWM/qsO+lF+z
TUpIgzurHrAJkuynlZxluOU1L6wg8g4JmaZPCgZOaStQkJgzqLGiJCY4epREMA54w5pKT7ghwwN8
skIngC8PwiGbNh265PRfyAehAM+smXFhyVtL78/1Vey9qpc8ew8Mn04pKiwPKCbI5mnRdzB9/y6n
o23eiF2CTcFNGazAejFoScmKbJ1NU04xtycGcKGO1a7uhkYV/PtK4HcwGSn4AKpD8DURhqOl9z7Z
St98Pljc1wlvOZfe0/cNi/p6dE5JGiglPFCsu66JEUqi+jhsZikdYTBfY9pHd1LTuDgYtEo67HWl
Z7iG3/D+aikMIwK0uB6zpqZ18JL2BsM6J0Zec3YJVCODlyXVPoVtxupWToFR52R4izEeYxmYnCIH
hiFr7WvIRn2riG5OCHyv4tLRASUw5dwj/9s60pZ6+Pm5eop50oqoNOCwfkxajACv6JgCGOBWDgEc
olIU5j97+yuA6K46IjK6vap3QPzv728WfeojEZ+8FsyRR8RqHRHJc2o2j91aHp7zcE+Xb/+F7XJ8
088hMopcKd6Zsvvbu4GhqBa1ML22t6XcodHhLVy30UFE0EfORwjiEKAHtQEXJpcbCDYST2o3dhiO
rg0pidsUlos/y2i8+jsAAx+tioY0fJR2U4Kd/RXnLgdGXxJxeS8L+12JHD5Qgq2AKhivlDNSBTV8
Jy5A79i2WO6ZOq4wPpFJMJpkJAEwkeMC0Z0DTTcN1XmmTDV2NoktaE6nJQlGnOFN3LAE4EaGmKM5
SF2LMJ7+8ZI+QqcmA4Y6Gy0yMxVVg+ndArnrrLkqFfDXb+RZgf0jupZW0gDI/Q8S5ao55DU9L69C
qo6iFwxnatvz0qeJ3qjgcSkJhvxhr/kJhwu4HuzeO/2NCaSiGoxie5V7Tj95RLIhPxw4mCeke9W+
04U3Td9IQgJzD620tPNWbC/5zrQzetpmrUbzNut+DypcZDsmH+2Q35MB8aeoWt1CIDY29qScMmpt
bVKdtII6eSFIk1fPf/W9+3hY8hxjjI8JaolmZmJup49mSKBbHW5+izqCPcJSWfu9O+9tIw2v/Xvh
+S2Y4gf9HqX3aZlKpk5982E6U50877Eb8/8wvpzGDw71SmFqR7fS06JUoek31oQrFFL0n1ORd7TL
0wdrDU2n5IRRdjit/h7QrjaKMLVaq0gUWr2AGuJ3oWrXhrRxFH9zDq7fvhsKWPU0on75wUEpZa/I
xg3rt9/jw1HpsdwX0lOdahXQrdSsI26RROnHfklZ0KUQLbgGHUK8qulf6yvZ6C5EXurR0wv5AtII
PveQS6npz0VTTsxLRttl1ivg5GBwg19ntFjRDdlc+1By4bttyTkK/8QldbPM1AXSIFNYAi7eDuou
y3cYeoHxkqLZyygXmmNG9NWBBgnI4X7le1oxd92k4bgpIocL28JQLtsccWH7EuDxd5WqeeFe0jRx
OAxMDMdKjryvG/2ksJW82BKKFfBRQ2iXWmwk0WRTJ9z15y1eqFokDLnoUtkRmeLHLpqcn16oJLbZ
/c0VAaU1F6jnMd0FoM4hG3/4P72s+brXZJwcL4JtOgR0ZQEQfa6FPOuZvSeNp8s+yX6x2TgPBrim
Bbfsk27l4TE0Y0pQlemhw97dpPVIc7bzdnOSUyoPCj7Gt79hIaNXsaHvwHbuUogqkwArukKCnTq5
mqARtIwN55bAAaPwPJepcbD4caW9fOrZjuoO2vfY1x39Y4PBJ+Za4ikDjBiHB0qMxkOhXZlrY8pS
h2kLE2FeaRdvzYSxrZjQ16NjRwJSJ5lLFvWGTJ+4Ca8l1H7YpUAC8R03TqtooNZS0eu6KlH8WAWN
lA5ReCIwLhpJGtq8SUPaaB665sPqjEQncyzSaFhGuez3HQvJdawZiQKVg/8H13BihBf4TVUQNmEd
lD6Kc9ubrYcO/yK7CwITotT9va0zIFIJngwkeXsw41F4xcLAIBdC6T9GlIuiIvbAlKUKM5Vkp3BD
yL6LvS6zQArL12hnOTCwMcFaljF4fu0Cr8uKQgwtg0csKsqYXkFXOmHPfkULr/UN31jQOz76e/kP
N+MKY0Om3jmXgawg1e90cTWebOEn06T1x+ni9YUfj3uEtNyJ7VrMoC2EzItHAW+0ltjojzOpO+Y/
dmhzNF2gAk3Y2ZagBIAoW/Ndd37ihYbEAr1V3HyDQk6I3t8rIl5Hjb4oIDn8foWeTsYEAl5Vc/5G
oV6lOfh4VYEG64MkysejJRWrkPWSoUuQhm3DsgxyLbrKKyK/rwSRgRHKyC7cVf74zJ6HSe1U5h6H
uTSVIlbNWAV8oTA9cZyodAZRCdOJ2c1Hssw1Z4DQTfxeALpLJtdcmlBz8JQDOyK7ToKBnG4KsEcj
utlTu2Zrg+MnCpzNjp+5k0AZaMduqMwHV3HbB+lQlsedfKf1PXahe8+LQ7MjuTwv3e/+YuNdPHWg
ewaRGBGMnw2kfHi/xv+u9VqXYV4AG+ih7o7G8VgNkfOg996Q3QUMgIV52jFBA+C/gZ1jBKoH65ca
kcZ6NUstUof/12ur9OI02oYcmRj481AS5pYzJ7XQVp7CxHDW8oilFxChcqTlbXwyKuxqsfWojK8V
pY2YUck4QUf9SlGM2qvQ5kXv6cAbvbfK361EsrjGorTjJ8Iec/24O/gsg/iuE62zaNQCL6TXX5zQ
gL4wzRAg4/7Q1v5wjxg7chpT8jvmHS/h2uLzkgf+bhpkaE5ajPlU4VBcmsWyJVTTiX38D2+e5GZC
HBDMfcFKVIEPNPFPFycFpCjWXmRNmKoEEf9kMpuWQHoiQ8qW7ZxUykzlnIyg97MVhtEq5xUSpp4g
XbBCESWWufqC0yB1POC+HeHn4etsvWRVuDqfHyNeokX8nOtKd2xgqdV5ce5CMtuksuBj79j+e44c
7hk8SZDUXIvf7PMQ2pfLgqz1Zmm9MkVOrWoqnjmAxvVec7gH4ldUtedtCpI6rO2TfG4wXl1sOPhw
s/lIT/VOJXbAu4QLuUyrm0Nj9p/vJ1VAEDXYpcY3shc4JbiZA9ZmKjB49Swjkf+QyrLPjLF3fPim
vopgUvgHwtIQAGrzvcvGxYPY4X4RtyahnmkJJtM0Myei0IrCvqhMpMA86uI9BQ5HNZ/NZeW9UOIE
M1V3IbHpNVqS0zv06ycN8OPAC0ZI9SarzSPySILSH27WmQ5toZNy8INm6e/CYioza5psiLW1WhfS
fg0p23eAPQ3By/pxMDJWMJkNAlbsA16rM07oG4yue8HWIcs4AXTz68i4cqCKAFKmqEONcfv8SC0h
E+gknWrEC5XUhcinETuHWAIUU2aYUQjwo7s5l3sk2ETWCv1J5IzSXwOR1u1Ov0ozlqSHXODzXT+n
pFyHuTOPin/AY7u+L4Rz5ZutwsFPWf+mmYcRN0keY6iimWfwTN8cOc1UXwb97XiHSMoehTZu6Tu3
xCXO+vPmB1R6Kq/VIZH1cwaE/lnxZ7LhDNY3VeZh6CYL7zTcrj0f85bhFrsmW7wN8pw8019OpJ21
Cq/TuDcXzB1r5109RmcwTLA73vRVV5esIhPFXRNpSNS5qnZ4iE0IWUaIrK5dC18a7LX165AbTOup
mzwaKK7/JV5wdhciaLA2BAlGXdb67daD0J7X2FDWgdSPPUeDV3bTD3OLjtIYPAbYo+80bkt3YopK
xqpMfPZ7bGVzsabGA3MzqKGy5yJ8QHUKRHC2jcyU7bLScXkG13SRrd846AV7SRkXaa/oAwdsO6vo
a46QstXHmKphtJ2MPkiZaHJ0tF5DBokvrCUL+jzGeVuONdKGbLcgk+l35V8c2oXTFRu+3QXEY4uW
i0aReFC/uP5DQTLjF/5F9G+/61qoUZ0kqM+dUFwvYqQih/jrpZ1X1duBHBZhcBi1L3wrKa71ZDjT
f98HqYLN8IX+Wi3Jc0Lz1rr5MVotUOyRXUOWOv5PbyUFSx/BT0dumOc2cY5zq4YccArOcVA5qqsw
1rwUUT+QHP6F+njci4zai5IQPUzcyXX7KZDFuHwlxZ3oyMj+1YfOv4U/gXm5/kMa4N7NLULgi1w7
vbl1pB0Ik6URpBgo+QaCgNfxqI8ESRv4NxTf3KY/THFa3tSkBmPP8bF2UD8WsiqHHXMpS1AimIRF
tkYqxPdJMcd1CHie5zVJpkfIjHYPMZQvze/otXvExSjSPmmzs4N0URZWW4s86KDofm/LoSjC3m6p
v+E00/EkjX+6LufGYFNYQ68T9rso5nt8Ku33RNbRIPYPE5mPtyXCmR7LJ17WcjLQuwUM6Gs0xOUg
4Nhoks8desHefBHswQIO8dmL8lV9c3LJ0gOhAz1cY8wNHV8wv4B19a0vi4/WMEbuCG8PUgpeQSjI
uML6D0uMl9CKXnCuZX4mKaju1Kq3B2Y78ZHr78NmjgEeYhq1ys2O8KmB6drz+aIg9RjbISc/iRtc
Vn1jdJJSNFZ4imghMELdeTRXNt9TMGmidf5t9KLNm7yNX3uWO6uGFFfpQ6noLZ4XjqG3CJuo0Zw+
EVqsMth95B4obJ4MATuWQwDHBidZvLAOgGZQ/8anyq8JY2gDAcRBY7faLGUCTWyCc9VWH0btdZpJ
1bplJdvTc8c0OzMVWOAbD8QFQkA3c4amZT4pWIU6htfoYiZthAvJLdiYxAzoWZaos2qmrR4gp3LF
rkyu3dZOtndA9+aScrc7PDpiG+fTZOztBkTUprFAhWPGhw3Ix84e1dio8bEq+sbNDW8Y7ZUv6bth
XcuauaQMieAj/kLyK5nSPc1ffKPapUYSa1OGhKW2gQ1Ri+3DxQv1XL9eEENVRQJMAB51/d9N0/Uw
5oKBhrdyhRW77tR4VpOMxgpf/EcjhvnYVtf0Eu/XV7z559up4CdCVoVNsPTSuKUMZ5wfG/IGpR3j
zihUDaEXzoQJmFlB0xebHvqHBZLp1Qj85xkfznkvajCgopHxchgF66XHydBwNDkPrA9Yg9y9D5tW
BhtxJis6QlOyhDRcUefB3f2kPoNq20fkCPC99JXlGoNxwE34cS6pyRhKV8Ofs1fYxYem+jZgKKEp
FWBJy+KSuFs+y+7OoIbwpM2kEwvnsKqftq+7indyzpQQMbRzangipPWfEpYOpM9ulvOfOgUDo5zi
p6Wdg5T1Or8thbA9qlqHWVxDXsTx1C9ptPNEIFJ6V6woayIZkYbRSsLf9PR25t8949W4na5k2Zg+
+TX0aIwqBdAZI/wcPXw3+4kO2AHLZ/qKJpGleffz4dB8I7YruevvwsgLDaWtN8BCdMK0qvQU57E2
YmhOD3H5jbf3Ta06Fh6A6u0gfMsozfqE5c4Q9+l1pgvWbyCmH0MRIxHsHZfglCJmbO+xHvhpGPJ9
GGXgmKKNn0jpc6xc80HCcWts+tXsAcXEdw8GcNUIkFW2kE1lNcVmorzvPpqXEUiQimYJdV9vJ1tn
yZYUoz4K8UQAWdME5KGwGdzlXnvj9wfBf6g3qpzo1vWqFQx5Ql5kpSlARommKu3Qldvg2sW74EDi
5FsqZiu+JGwLuUVd9eUTd3Tq/5gvFzuTy/IrBg1dB8d5Xvx+CRPLvcxSDFX/5KZ8joy6z0Ex4vlA
tKkJVJ8uzB/hLXTkyHCdiOFyDO76SM4TXzQFAc1HT55RYQWeQwi+nGcL7MizUYyPIVNy7Mv0W5G1
zszmJ1jxst6BwSDs5KGuwfcoo3TBx4QjGWiC7kqp7DXd9fFzovb9OMBwuvtNar1xpQBJrRcGeJ/G
DQgNn4jHiUfRIZKIz/c95oJVBJuxvYMSu+yakD9mXzALR7CYbud1UBwHyUmHUaw46+dUVbZdb12W
Col/7e8SjZxF4noODeV61ogSubEP3bJ402xY4a9NcSqQJIlT/7DR7MFBJcQKeeDLr5GmYClbMXYi
fWrosmf8ZQakwnvZIroQrVx3K01ZPxKx3RmQQEcbvF6wX4RTb5r40SgB/ENM77u/ufplyIiRHZet
CBxR0CF+8e7xarC6/6C789liFVL2jd/2yvTgeqbCmp5sUJH9KYoQfpjlmCduiOFBcatNVy/H4Lsl
tQ8TbrVLgzIjKuhoG7VrJ1qT/EYvknrT2gfLz6wX5a2371goDmR5oDMDEsj/7pkUp9yp6vISwPNO
OUkuzhR/fOAgfWQ9boUx57obCNCtRTGdjkUfoq7ZwiHSToxmdKz1G1Ce/m5zY+q5FX3LqMTjPACM
Jpbw3/MnjhIIu2TBJiwWil4vrjh50DaKJt2w5rLvoHeCkY3XJwWdMY16k+hVrt8QlwSg84cDuZp1
v8uyyywGRdTDHk5orSwnuwpVX0dFX/GiGMWuzLCz5KC5ie6bdmx1B2pJrfuwKJYkQwYgCDdxjm/E
azC0cWqBz7stEDmhFdhh7Tlb6DqYGkDs+7MAUS+Q+An1vBHUipqpJrdsEDcunigQDM4X2/VxPc7m
TgUO2o0KekVkDYSR8He2Z8WW+1hpLOCNzMOrX9g86xNax//2guQzAgp9O6k0C7BBTz94/gPFEguz
ZJznA9r2azP7asI9Fry23PM+pKaDBk1H5NVc9ambBExyy/DBQrb6IFOzoaZHVZ2JFU8P9UwcFOkD
2RLnJhmEvhuGAQ6YkIzB8oA1HgNP/I6LIMVqIbsHVFpNAISZObIRxeer1BYPTHpQoSjULFsEf5R5
N6LVDVTJxxnF1X1NjwAmKGZzScsg9BRE9taFB1GS5aHT024/sumA4WwjJBqkh22LxNOV2D+pAelM
KEK5GO62mBbMzYcSV1ZJSRFjk+JB88bYCblBqO8vWTRk86GTRr6uY2K6amYKJTEUL1UAq5gOXk58
hiYG6Q6Hozsz0JNqtgCELrNLD18+J0KxKoKrFfN0KVlSPIlj/lMfqIAqzXEiILwSfEA5pewTvbBW
Qi0oIblDkyEAH9Ak2DXrQvU7zuBISs6NzRfve/W/clb0zVXa90Xp+JtTEiZsx3PAQYM1Qb3d9fOW
eov6iNXWQColz5SA4NFcRx6VXVgmgui7ELXFsf0SE/pXfhZoBGlNaJ6xZvVwtP99T8EHUEoSu5MQ
vpj7kt1y6LQMr0J1nc/PodmufxEDk0KdtBXDTUXN7sfTyi9rTAXhkUp1y2yvXfawhtUbT1RCBTLl
L5eow3SjvuNgGa+Y2HiAFgfWPTtd+wT6aBw1E15EewWcy3p7OP/otw1hQieAmQ7H7kcghN94z4yL
kH2iRGaKk8MsMWYd6Qnz8gOxV58ZSKvECv5VrMuzTSyKSWUomrnCbsMM4vB5MZo7qss8BRn3Q13e
YADf86TKzjeBzN87Adp9WW4ndsV6aX2UbsKrKZ32qynpClI3PeOh2BN34hGr0X86VF73MkMC1lKo
LVD82/uKYyry3/PTPFW9/ob+O+TupJz4OzRsjgV/tdSxcEXUAt9DoPkWFxEvq7c7B9fmMHw1uGKa
EBvCezP0lFpDTWgl7FGLeD4iRpr2PSg6nf605pGTKm806kYcGrh6Qs0wL/ObCSikZ3rBvQe9a/UZ
Crt2aGZ/lasIp3ij880H0CleuFeJ7Nhpy3UamwkDd8557iJdzMTbj+JEtw30AJTMXdd0z/0YHFFx
7jkEKyiZPtf5quHOY9AZH5IZfpWg6a4LoNfzFr9KlWhS1rJgQvaNL8vI474RfyJgtuSHTJKuSSXB
id/IZ/TEPnoBJ9h1BHgHBN2EDsWoxKb3IjhjvKd31odfoD/ZwptRvk5sAYhMeJCoXtFolrVxWwFN
0chZrwzl+KAQap4j/C2dShR/hrxwK/pA/TZWCKXdBNWRp9I6cDrEgM0eq7q4Xw66T4Qrf+T0w1UQ
k3AQoZ680mhyKvbHXSq/XiCVB/4+Mh/3/kATPXjyIyX80ldlWuIFgpaLTdkhL6uMAdN0LX93u/zv
2H/K35lwZJk2yQ9wGndUWIQVzLSL/u66IRs1K+gU+GZGObe0C3NUXUqyXOSXvKETzcklPEi3dbkP
HjONivMYZci3BhvEMsQ9bi1XIo8H2qjIUjr/Z3LGoz2R6aVp6M9qjqH8aGw34gnqfkREaZCnRw6b
V4zNB/3wzPmgMmwhaXqIzE57/ze6SvmQUl0vw5FFJoKB/VBtliO938nge7xp47Zkuk5t5r9Z5Jl5
EmmUzZjcMVZTP4/8A/izmTaO4w8S2nQrfY3mF9U1iH23/joyXfK2WsKZbr23dFO1iH2CBJZW+fp1
7KSkOcbEDsf5PvF4phDUZq/E1YiKYQo9PSqhTYwCu2rgX9jIWm4rn72t3yu4KsPQ9/MKq5iTJre5
WH9hve9cvk6c4f6NYmYDbIPstlngUV3d35Z/RrCEVBUeEWoPkJEYAomPI1TXQdXvQ6ERqzwybrl+
yelbB9rksqM+Z9tpFrej2krBCEIVXAFQb/HKMY0bbRQFZkJb35/suEAY2EXl/wTdyXt0gLz9S1i/
D1gqVCIv3M8Zf/zYLbwaaL2C6ths/OkF0T//t3/jvluJchQTa0h3Zs8IO3ZDqZqJOu5czNw4bDvS
43I8ZODYnynyLbU5k92MkGUnjrLpwDZeL6Q5mFPvF1E0r5oEu2UmjjsR5xoS/HvJQ6pUsoLZivuj
e6nQBTzFBnRVMp0Lkr/cs78JhLowXJyQiGxgiX/PVxbCngxZ8j5/UiB2zQDkx53qikB8bBtb7SE7
ElA2MdkgHZtzcEQA3VBq4yMBu4y+PXV0QL23vKwEjmlWEQIHaJxBknGLidr9z6r7GA4NXx9L1zxR
BN5Ri7ExjhbZ5TWqnndRYoYtKBLzZA4yPQ3tPfydMc6ZyBeYuCxm6WBF48VNAZW09/khO8MaifgT
hOlhzZlOXMPYY0XCS7m6onJ0DK6eoKvlzyk60RCssqlGiJyNaQc7AZkcgPSUcucVov9Ct8x5Y6EL
otlsC6WwNMhHsqQvyenTCnBr0nYiMsg1wBMjGVPGTSK6PoAt6SsIp8Y7Vq3FupGpVe0f8oJmaaqt
4n8w+cL74n4eR/9nMpBNwKws/tJDlJsD8c2oL8X+a0qi64hCgHEUp4tcA2FLvGvhHgCunDsjw89c
PO7Su1wL2v/7zDmC+11Qn+WZqKBDd+zG+2qiszeA0Z7V7j9TephYxplQtfrRnlcFqXAaWYptT3RS
xc1dg8KK79GbduuAedgbKoNTj80H7ii7sKA7nLKIIOcaege+6W6KC386HWaou4NR8KWP/+Dgq4vz
aspCDgi9MB/HDSPvrx89htx/tjNwfMf1gyumhnv1rj5SOm91d/diD6yNFlkH77tmfDJbi/Z5CdxW
uiyuGs1HPBJ7puxm8HjontWDqNu9KDTtgV7rkjG8fzv7/geBiQveOYa3rTOASY0XK5M/xyUE9akW
vTBwuvIWx+9HyJOYXqygQ1a+Tz7H6K8pI+5UPgztPBsF7wCS+jFem9vYMgv/SqjJL26/lTUKrUz2
WhrDvcuXBN8nKIZrj8t6J1W3cJzu0LgeR4PDm/1qsH7CdWVLfbvVMx8yiGi/A9JXof9fjbTnpiVF
n8ABjxrzFHW7M8EA7D9xBO+b8Vb37biDbjrUz0RlBB0nOrMR3SnSzvPhEWg1oRiGk0ARXh4lQX1o
VXPvpoQBawGSmOgbuST9ogouF3yUqnzDAwNmuqbmIWSaxl4GRt9uH1wsGg8AyZZHA2O1mcAGkh0T
4F8Jov7D78tUwIOsSICt/Ab1/S+FosNva73l714P9q7YUgzAhFc4MIUvLOf2PsUUvdCH7lkHoY1D
yxgVCKhb7lqSOUsYOcpgJFaOP7UA4J7JY1diByKZ5q0h6E9NGvWkgnDL4vvVEAZUvND+o5mxDvcD
BAH3tMNFyk06BBfKauMpiEsNNKkeioj99WDMMb6nYI3bavx8meYGgafzYRtk5Kbzx8pNEKnNLj/y
oVYv1NRVgtwGWY9m7XTZvsXPlgnesayz2VBfKt0umuONTdrZ2fiPqYDdNYlUg1ZDCGcVFTxan3Ee
5/d8fYGbKgXJIMdiNYTfJ6BUcYI/Sz4sD/NRTnj4GSv7bQ4SYiSePu6q286zEceT1e6Y94Gk2Kyx
jE6fcsrNPzzXzmiv992AcP/yi0Ir9memqFQrjYiPDFt6bhcpR2FRTEJgLe7TEAcKI5f4D9y0UUzL
3Wm95yNtUYytxZifqc9j4bfD+MOawB1nwyy5Yh05g6wGdP/0XiMwguQzrxeSaiW4BIttdu8Hxh/F
ROjIPIWbecW7lhjF4QxsJ2Sn0uBEdXYxyut/6KZiGJAhBuC+d2cFy2Lr5bCAz36RD5RWp3J3Uk+k
66XIENa4A1ItLzWdWZWfxb4KtbUlkxXA8UDfG+Sjv+nDyZkQ9eWIuczTfaPbr/ezF+b/wyMu3AiE
qTxRYoVVo/cwqE+YF/kqCc/omsHo5dd1d4akqj1I4xXuQH2sHgLOLfHG0xNEwp2foCbX5jIpeK2i
/V21pMd803PQcs9irE4ru5YmEMywEsrj3rTTR6ArLzVOWx2G9uqvQW4B+Sove4eVd6B4CCJwthUd
AI+xf4AtK9SDbK43oOGZBOWfsyXYNZ1VJ6AC5oRVzdcz0+4VNth3CGdIbaEofPuNA3Zspyh5BAy0
b3jVdNp87ENyQJ50XsAo5A8Ib3TZoFkPrKQGMYQEtQgVq8KeOawF2/2uRkPDiQVi2ZzIRk3Jvcr8
PthA4OCxTpFcQKlOmJI93G0V/3CWcAufBK4uJazJKv8srntfptCfdCVp30Cac7cNmhJRVLbxw3J7
oFC5yQx2nu+GUi8svmaX0UXmNnZX9Qe3aTny1Q6iyAFpQNVJWQQ3AtTRBPy0FzdxVvj8HrWll95Z
w0YMYUPOzkvt3pfR10hJftqV1Lm30aKgnJ6O2C524RtaZFSDfVmTUmDx50JukX24k3QEj60MiCm5
AIxXkX2EMtrHuvwQhqIgE8hM3+LH4nsjyRQyFiD4NMNJW5y/2i64Fsx+obmbNbPrp6Lya0aBPqbs
kWLPGGO9lLPdjzdrGj8Is6kldirH/4C9J+/yY6uCLHeqQDdeGrzSI8WWfMdODS7aYGHG5RFWJGBM
mxxZWCTphlRW9wAGZ7HHijsd2PC8ovxJcumUdLjDLkidq0s0ngMkyhHgvEJ13TANw5VNvp8JR8t2
nwJGx7U9fLx8m71cQY+eGXan3vVkLTHJn8keAH+dmqjmppuw+hcvlzS26KYdKpUKr7xlfjURBJCy
XQXDnyUnDE7/f7810EKc9YhLfNoC5CxhGYIy+7hP4ii4zmvGDGzxyOXaVhuBY9ddQ2PjKrgMiWhF
cbXTsINKVFliBcG5SEYivJwgmMBDVbTXxZBphale9RwKPEJj6xs4OohTcBWKF/JBu9eGWf3YtZ+J
+JXh9eJMAVKWt8IrQIWG48hJ6L/E304Jm1KCIinpbHRf76M1CuHRZuP9+6P/d0BKWnk1aFI8Dqnx
BKLPrLyChuv6KwDzuvBw/8NFEnmNu+OuQWIGNlEeXkFwsCUBS3AJtiVQulC7sx883OoDVK/BtQjN
9OlnMvGC1yRzWoeYZJ+twi57N6PNDXq3QC0PD3gBCTcTgoM3Syf8WLoru03sCLIIo9obcVpnsmET
9V/X7s9F+WX6IDYV3lg1on/xid13I9W2iLY4J9a9nsA6Tpn2ARCtu48awCFsf0s6zotYKA46sP24
2VB0vEX3Q3PnXigmHtjZJgk9PCPAbvePRUCbbCenlwRo6Od/jJOpY7dRDi6yKj0ixJz1hgSEpMfK
LabiCz4Eo989S9KVVi0B4zFUuNJNQuM2JacY+kI80rapnQv2KcVLrNo3NFLB38AvkPNkGnuyqz8D
w9kT4q5JAxyYvecjunsWrKZC6zOc/jOAMN1wVCpOyKQ5MkYpUIgnjdkXNt1KeB5Xg+eUaZDlOXZa
TPpPhf+FQVC1gwgptLKL4lj5LNnNERLJT+9qN2SZZUS3y8QXbBV6YXWEZhDBD4tCg4AmJKzthefS
Zifw1XwFsavCloeVzV2fYtOTWwZHFaLTFbdWWqL5HjnA46IXqxAy0c6kMzDQV69oziZSacG/dydI
OFlyTe5pthAzly1ETUTXx5A/v5Zhb/csjGIN26lK3cL4W/ElKaiheWuwCODN92nUF1a/fLdcWgy3
1R3WslH3f0SRUo/ur18+tbrXIhJOx2dHZrHIMgb66keUk5wOi1lXfVsvkdYX6/YYaJUuCCuBFOdo
PITdO5PrZVEc9VXsC7sumd6mLFG66+Fi3WUODZmCPaEbGEs9XOV4Ili0Y3kjN16iEPQKoTAlWdkt
nnNLfKl/U/v1Wi1n/ldAAq+Bgh9GkRGejVz438CuI8yN0eHtIOyPqC5h4vYS4FWJKVaCtU/0GHOp
fv3/zQ9DRa7SiHIS3UZKUGntUb0jDFC9eQfm84amtkhDMNLUwRUKDnncIBv/+UbbNh7IbZj1mTXT
3hq260degIaeqvE+I4nMv/0/iKnpMLfRULmFKyfJpkB/QCHBcnAMPUkdpKDVvMLlAch5G/1jwJHt
w7UtzDKzlr8H/qzHrB09uvx3r0qnDabDMYtaguqwmzvC7VdDFQuJ+w7chL0Qws8J22x0T/t/c/az
6yPU2lprZbBS9rawNMtbXT6uRuD37tkphtE+6ZEvJfTGoyuQFOxaO7VCd6Yb1EoBX8/iKZ4TFc3b
vMAHlCFgEm8/4VEyM2gKzmVlFqHvKlv9ORDSdQsQoUlN50TiN8M8/9mX5fiaevTzZr5F6ynxRMHB
MxZnC6nNvxZL0RSwB13qC3DLClp6g62gZrq0ZDTr5RGL1PBx1VSMqFcgRja+yfhbQ14RIV+7WMnj
1Sw8StiinSpj4lPuAqxkn6RJ9Nj+cgsgBaTE4VQqupEA4WR82dpcy9V2e0tR0Se9TQJEn7mPX6RJ
BDcs618mqM9wyhpIPtYFMBoi1f/BoS5mVDNljBhlETZXfMP7UIRZdgqUnfqHfEuC8506mxQVXZEo
5RvpChx0IAQXMhoujqyHJo1WGJWRJx/Qg7aroBD3hpJxX71Kw/ClyMVxx/uwRW5NNxHqg+YdZ+Uz
j8oyMUsekM1u2Tay+54B4YeqZY36KpQiQSERL1hM5UR2wNt+br2dVTHxMy9/AuFDa5+sbUT/f/dJ
svsZNmqIBh54pju2go2sSrNp5PXiR5LkkmFwym/hmfR5EUcgXwXWqwAePtnCI60/mZbGPVzb75Hg
V3+kkPvEs9rBFpBvG4Eud3e9fOyE0susr4NnWEyAmqg8xAGvckz0Teh9195qOpd8stLzKrCgRjie
VHRqC+jrS/j/C3MwQpmvYtJaoCcpsipL6T6F3j/siC8VSsGm4rZwLXC04jjV24OS+avKrv9qSYRH
KWZ/pf4VgP8mTeAuCLbl2x3mjr5C4wv7ShuKnXXfP39qXq4sniFPFIMql7phtBUa/5hZgCSvS84d
JjnpzhZC59tuwojINHZVwxzunoRcBP2BDSquCWP0c3RGuEN01J21gF0gpHjuCkiORoxbwAYCV+Sa
m9uDScMWO/smrXtHnt4wlymVzFzz2ijkDPZlqujtCUzcGGgM+a3rFsyfGkXDMuZL06sIflH6wNmz
fEBASegyFsY6puzH2AHkqVkxxwvJjm9UP92oQbWG+Mvwi8S2OIpoEJyXeYN/WtCDPd1PPsSV2b2T
C7GlRgrqjK7OEAasyd0PdGtVqt2XrODaV7mVHiL9hEn3ZI0kAOs77l92nrM0xY2qPTvM7W2cTN2c
KOWVROns0d3IR0pSsOqIXEuxbbbzCtvEKQYQfknLsUa98YJ5IcJC5zFgqCuy05zNQvilew1d646b
zKMdXS/E0PejfrCtfkJtgkCFoaNawYmfckWEntf4cF8BMvmtmJmolN0n+wYq6Q04UpCdjaepxH02
tA3CdlSL6nksiaYsw8fwQBEtxAbnft5QfHo4jN4dV5W/q6twAxLHgdOktHP6lHyvlXCPKV7GsxLk
8qHvtFG2JQ9JtQ2B6KPi/yAr/bZ1XiVBgmw6WEXh8XJonR8MHe5acsCnEFQkDz0k8tUiKf3nvLqt
3BOqhdyLyW/nwIl7JRrkn0wUqQm97t53HzbrtVc7f2iSPSG/Ui0KTQdjoCPwWdgvJbpsomBLrY6w
UphFARI8wbKgXg1Port/PQp5IkxLwZdDs5f/HzEnte+jIilVjbS3X1RhpQqIZiYVyMI6pOgsGG1q
AO/kLUsIkDaQZisVuJT3HK1mqwf9NGRVuCLJqxaLAeRWfZVeUgQgBbDqSKzcJ/O1F7o1KsaVwBEZ
ayRD5reOR7Q7vSlE1qbKniIyvajCW1s0eeODQo4jR2EunoXhiTLVlkfHFNtIsJu+kU1Qm8JmKt15
ZythP7BT7CWtzht2PJxC8x3iFKX9nkz0YYDNmYOLXPDuP6Sxdu5NUvLX6i0nhV0cgroz4yfkV2Ex
IbIOlz43nsKTVbk/4qk9YaBlCuMTF7UoJFZsaQMVbZaiG6qwoht9/UvmuUnCKzx/153AMqPD5o/L
fjDJxzW0+w1HDfTkq2pqunh4pRGwM9lQqfrVnB/x1Y+Jn0VPY4oqWkIoAPfJrcDTcIkFZ45UA0NQ
75Bo2AwlbscgWLJLWeyySO05opcHATLw0E8poTXt2YKg444c0qAJLdcuE1lllhyfroCBievBJjKC
EzFJqP91xaV0gnRDneQ4p1Ocvrf4jXh2WotO3IfQi+3A5xilM4sCYx6pGgqZc+sMEP11JhfMF4NI
5zgS8Kv0TZ0UQe9tlysZh4WNL0+epUZujJIaQHqAH/k/0bYh9P1E/wacvCnElmI0UsmrLsAYxneI
EZvOB3TzKiKG8AuaBvKjERuqSfi8TWSb1YRDePBFq7b3djBL6zhzP9ZP8qXnQtCB0+rqRYu3t04A
sXqZCXfRlka727hwcJq/Iqazv+luBUap21RHmQ14L14WYTHEgFA89/PSjobDrsRMMiiDQBmYZ5VB
mMHweSG9xlKYyKuP/oDkpzauiXm+9Y/uFCL8jXqkggvwgGVWu+cq7hL2730tMBVsh2/S2hjHovGk
o7iFQ4B/sPGEVSZOexwLtwTx4MhGvObSU7hIg4pSFtFQr29489Wfh6Fn3TnYiYJFkE1f2Jsrjsx3
L/k6hb4xqR2jQhu9FbgRbT6EIJ0yyXDCqRm4aCm4VIEpjYYpS5nt3BFt1s8W1HxVkcRpERPI2khK
0U1rQLy3+9DiXXoBp9RPSnTp7k9s3VPU3wgf/08wHn7IjwZ/H+6LMP9pgBbUSJzapgBGFOsx4FEq
qa/H25kiQqiBtfNdg0VsmIC5EX5JNnZDvK5AqRS5fAQBidYJY0K8tCcjtgVpWpt3B46tpInr2Avj
Q6Ey76UV+ezvqt3JuJP+hnhxMmPHyiPNx2SLkNJAT6LYUrtGhQIhFpFOi3jsEJ9A6ZuepnEXc9pK
9fFj70me1gxirkaV3ZBVRIRdvOWH1AWBnSm9kKi2jTmSnf58hZnFeOVmuJ3DFC4vv1hg8Ijkz252
hiCx5Z6dUOp+aCpWLp26rc/rIbl8r1hFbOkGgCzRObbfTTWVrPirkzBNbicTz8JXzvtaumrux0cS
yVkcKVBqtjc0JVK6VThGfzMcMlYWBllkCEBrebPTFdvu0oYWHhbZV/OQWZJFGix2+wqxU9kDEv31
lgB5FQJxl78XFvKjPEFw+qF+jKfMrL3b1U6pbNlElbFv8TT7qlrxZBS1tF9/6jEQ4bcJxcAothWL
HGJ3NnpuNRiLqEY7g0wxbzb1lANKl5ttg8Q5z32QyDhL+Et+vgvDR0P9h31eVcsfpE38LEa03cb3
Yk/e/9l+027TC0/8YJMbUqyxhQaCztrGDd2yttlSdBhU0Km2Ddbtn9M0uwHS/S/rU//V/9CdizOZ
gx4ggJlH9IAMC13SFY4juH+yAHn1ngkczhAHQ0KQt02NhTmpq8ELz3/FmwyXrSAgK/RvjOxpPKlo
rNYTYnCTncY4YruptiEBRtHjfhfN1XXqmQW01NziHf3r2RI89aLIIGUF2RluJPq8CaPTLKva8Wjm
ORXZUltloj8bi7pbntYKNCS7mIlezxEGEMHEgWll4NhRLFPOCh63T6b10Mf4Ny2VIr/2Ii0ILHKI
wtkpY/rkxv57pb2wre19qLHk7HfjqY/FNzksKfBpfgGFx2kQmNSS725nrgB+oDYwCq4G8/nNAmLT
nbRU5PfSmugN3MdQWz7LG44c0vuu7vFXXbETve6pgkKUkhUQrLKrtAqLHQIsKOnllnX9G5qzyofa
HnE3/58z8e6tmdSoEUZapjRUaXiIur2RthRJtQMQTdz79LrbnCFw/kcV2FQms2K28BamClDueZJC
gjiFXERi6pcfcGtmLErjeYFsid8cWVgKO3veb1Dcx/7sKcI5LvivfIwWnr8rnbM+wb9lBW0KdsG7
2eWoA6ONyVlQ7z2seFQUXdbO3J++ooSCBLYyNs49FctwOjLiPpyHInL1BF/7vHimwddJ3sFP7T5z
pXLAjrR0fgmz86M7OT2+oZszS9lY6e5pIe8ybyiLiSSPIO6fS1NMe0E6mS+e+cikCOci1f9AyoKy
5ou/gSwrzTALz1tPBsZYjk2AJKUjtjbV/OuO3AuhTnK7S5gICGwlo6F2mkJKzgMi8mPVDS53pmwf
mU53FsPRBq119KjRb8yed+lFNc4xnJijN3tJvazVFVNNnJMZWuhzJjoRjpUKMnpXqznmpsBNTEMo
4UjlpbpCK1PoBeZgvHxRqdqbu3+Z0Odvk3ThpdzoNhfF0NyAbQV5zxn5G+OiMn9K/wBBhvb8nIq0
i9JkdG2qWMwdX6BPIuxg2gBnMSmhVhFaZnUig/q9EOBGC3dLN3xPYQNM8k40N469tFK60GbBwTQI
2q8LLc6S5KcfxOkGadKBPCh1bQL5cRXgyPVvM0Il2x436JQ+dYRHq8ZuTlD9ZkCo0suCx3m1Xq0s
ajzFbD8h+jV4Kr3MKpC9rbVBVSOkb++7sXp7aKy82akZlARqwNOBmZRe67TgvKy2du2K64HwfdCx
Qw+YEEJNxW4X5VbZS/iJ3k0DVpYpQH2LsN7yKajpA/4Mk2nVHPPuzb8CWxW8cZozM533JzAPo8eO
Bi9srvOg3XX/jq7eyyWTtY03+CrI++1z1dwYnlgJ4DeVKRYRCtwBN7pTbUI1Z47kI4WtTMcYDvQQ
yjbni1KqXzmOwhSYWYp36I/Vp8YdpQ0WI48zMu1MDM+5NSDEX/NCMBncX9LgJuKVRbRZ+Tdr5pVm
rDRTddCuMZ2XuwZqj9wkKMXl2nmptHvLDkS45hC9ouiC+Par3v4H2IJ0MmmKpxqk2qRddjfOhXl/
3v2GqB2LfECMZw/mgI4IhDZsvNk+pY1hLPI6wBq871Z17/Gx7HOkSlvwmacm8zPNlJbp6umlfpVG
jsId1b4QEALMLfPDUoLIHnb9bgcVuPhABYGWpJi9XhVrT/Kp8JRKGcgARxuv3BePjZHHCfUIS5RT
WQc8TksT5bKxjwj7DeVsf3numf0upTfZMcVCmffkXqXQBJCkZ/WNNTRA8VZnyvWISuawNMb8eUEK
aKiFDam/yZpCnPPLG5z1t252+KqzS/n8RkxAO/sDuC+7PVA1shYwlXzXralXx9115lOIkUc0a7cH
gi+IIXDUPQugRyA6XMdk3Ipk3LqBkZ7VpLwT4f3SUSCH3zX+92ThastIXgEmESS6jCLMExsZQh0G
0B1HHN/Ddw/7nDVNlnMBnms4aODal+dJBULMKLMIZ3jSF+Zimz02oTPb/va7SAQzn/Er4jhsy3sx
zVdKe8Do9cVsXDZpjdiLfEF1ZelCCuxJI/bNZc+zCkbzolJqE7dE+c/bf8IZlZR52QE3ljABbcaE
IGpiKA54BSeUeDBgYzHRsgOp85Q0JDd4Nb8tgBkrhbNtC3AcXxAAKu2HtsUEjpb59lUDH4aUWIiK
mflhu92s5tDHE6OO20DYLAMmB4zzwUP04R9hEZstiwwAj8RCFui+yE2y4Qm3dx4qf8U3F0+XwC8D
auJJKTWNLZbdxnlfyBTprHCCaI2GGlNkKsZkRaWF/tV6YlsDyfaDEs43ZUgDbzsNuAg8wtJAlOJi
T0k9Slp6INxb87E7dRaLWWqukCsRYZqNKQmGojDgyT0yrxsEDXxyqni11/NJTEicByUKS43Vpz8n
2dcjX51KwWAE+zOAV/zehhnNW3ltZtr6JBWAplHdEocTQkSOf+fYtJiv18FEjL5OWi7FD/9o3sPZ
msWo+P+tadewJxZ8cBFn/ezbVr9eg+Q8OHChRcaGeQs7huBXFWBLQ2BlP/KBKzm/DELKv0STsOIL
ENKDzJNRnUwwPVJb5WEsdIb5BYIoI0bkupVRogLtK0/Pqz7kJ9ZWJlGc0buNDJQ5mWSIf28LsaRH
xtPCtl5ZyZ79Px3HybSnTOA//mF6LfDzxAr4LLX3YR80y7fcDwJxawBDZktfyK7JYsnVOs5XWIBq
uN9EQC+a7voxo0/E1YArgvre55gNoekJvKMRGeaZo/asCPNAlCEuiD42VVOr2uoTmOdKsbLyUUuH
6MEymH0ZRh9+TPFol85rIagqzH93XhvxUyDK5p17y4bfHWJX3NqOtGzH9+yOzNCHnYiyaMrGEd58
WamgKwXbkoBPzTahpzVY1EvwEnvIcv7ZlW5130UwVmmo7yveMeyuZfdKYlNy0yMtFcepX7B2NOl5
4grUY59tC80SBHcExG3v4/67YaYPB1FxZjFE0eep+iPjRZ1VIxP5WxLIxiJvZ5lm4tj6OmfrT+y/
jcgot1Gg/gItj3ecA66YDn5GUv9BCoL7KZ6p1krmT9NVyz2Fa02MxXGdbv/LqlzyPqPK3iGqlBY0
4nB5AUbd5aDuSjrEI/oHuZAlgd/HH+63n7klP1y3hO0W9kIs06ZcKtnSOugmj1b2YtPeD7fMi+OV
6kG3SoH/XcqC6yu6bhsKrHl4iqN7oHj3CmuoQc5Ejtlr6ASrnAxJHsKGIc9+PJzqgR7yE468cuCK
VjzW01Xjex77qZRTrhVxsrTakySK6Vx5wE6bZYT8m26yhnW7YO7mMax5mVKw49Pj34wFZ/xxPUEs
KtSbJMyPVzlr943R+VliwzqFg20VfOwUjafu/daxtSxLkNeWea9tEaJ2Xud7jvCpHNoc/Hk9BDlR
6cAxlAomwmNqH+G34sOUVAErFbmY5N0V7bM6X+Ahpdv11PJK1njmmKVU3wY8BSNU5xYBOadyIYqF
uWqhlIblPimtNuBhdszEbmMoZLwP7GNAfebzpIIu5QWqqCFGgIhpsuY+1T9UXtPUGPFjznLdNByj
KWf60G0G2qpWvVKkj5gDdwVUEyfAHrIsiMhKnA+A6VuUvKJDc7DQoqIImEueGYkhrxyCRyVRD7ry
VqaHOrkz6CBzqLL1P06ySDEVRtAOviA1+BFAhUP85KohBNJxAudQLPr2vxh3dM0dW7wRo2ACZxPA
yY0r0mYoGvvRkLppoG4epPwb9bkEQa0PHy2egGzMfuXP2LmXEGiJCzLBq0QZzbsB3ZTb4l3mMLYq
Ek31YpJEv/9QrGxZNMiG5bCYXfzMCPoz9vYKJwDtQugXQJc9oqiVFNtI6GJHXxbZQdf/aBFdzjNb
wrHiaP2nwmYFgX/8dxcm4Vf5r7WqW0RhNRiXMzMPOpFW1gPSd9j1Tqw9R6HErTnRXLgj8xS8UZ/g
CSYLok1muc5iC3eS1/MZ9ZHC1TPaNVXvoV0q4vgHNPUtXuFL+RPVYFeLyh3TM1ngDXIAVddb6TY6
oyjQm2qSfil3j7wiz1pgcfzRgMc3YKiOjWSRzbRjF4I1Eq4ofdqiMz1diXyBoSW3C81Pbbpx7/AX
oC5UvpKtJhfMwN4mW/O3YSBC24dAao7nSbO4lZhHAvF6vHvrU5+eoqYip8rNc72yu3UMabrqK0ei
nTqZXwX2Mk3K3wvMXQHiVxSKkGjZi84qiLdfP/fLwHZ6XRzrj7o5TjAWff0i9/yRzxZPvD/58oj9
wRN44a7V2XrZ2IA+HTVVJZF63zY5m5/51NSuOek9F/yAJB7eAPi+bF3iiONvzUaOCOddouCn4QjG
hmwBCx8htru72uWb7db4+24V60bhJr55nuq6Np517/xuo9je3wN71OxEiwzn30UiAmomlCPDoux1
xhtz2ilFb63DNby7Dl++sKtfYHbJrRlRps6jaRnNnaBdBculz/9g/oDCU7vIsFy7a4KBS+Ido59c
gtAEwLaMqAP6iMJ9YITr2IbnpZb8Xf6vsinsyVWx9xelPi4YgDJry54s7UauIRr77Y/YlVMbzDS8
oPh5fgXI/5+xxc6JXUDURcETyrHqJv9lnEYEmvqOOewHLXeod9Il2p6Jucrg5nZ5haIevMBR5p+8
5Uq8P1w1cHFaXTn3TFMX/cR7aaQUkc2iOIt4sTTjoKDiyFkNSuSAr/Wci+A15upPETfv/B9EH9qa
RdxpIvrpGALyGT2lUAXnZRQ8KW9hpbodTInlSvmnLRpkEBfYEt6Ak8TgWCmklQ89LDv2bFyJUTGO
ONtADfrfKZ75LwV00eqOZI7xfXTR89bWwpUietVXixy1yazFfcnju/NDf8ean+hCQeAu4cjqqTI1
YExrkdkqAbO8lAZ5trn8yg35LNdALeU1biYFd70OX6XHzA6hmKjB7eVK4V73uCn7ISB/2iu+ZO96
kPxdUSlRJx2xBfBYiwlP0sNjVHWuHd0RKxlQqnJsNRh7ezs8AgQNnAZ9MW0057PvzIXldV/jBLPp
idIAAHmaxijVO6uGTTM0cEgzvT9G291cA796fEBXVfYcJqyUT8gyFWJ5cohQL5U1glMY4sHkGC4K
//2y6Y4HIIZhRPEeR4mTPeDKh1t8jOLxB/SgLcRapHB5tueDejFJ41/JqqMDVO0TUVRqIsCyWovR
EvzmmoSZdYC5xW7K0hP0vGFD1qfR0JmyfI2zY9gamRY2MUz6/DuUe0x/5TbzqBFjJEDJglB9lhEH
EeMZyZ2pX1FjX/vjf0uNimIOY59FdujMYBlA0CBzhuWaHLPZ5yM/vnyp4fWZd8RcSen1o7C6ZGiU
23G4ejSBV8mralsUt9Gj0Tqsmv+2wDlb3hJthRnFF/THFdbdV13XSUpniPcz/npGwInbUGOI5MXF
5i2p14eeGZogEcS9jDtbqYhjQ1tFBMJDfL60scU8wPx7bGCmDK8LW0C2y9kDyqDhE6ZxIA6cXSbV
Tptb+c38Cp1SPwPhx++dXFpiOS71RYFK5LpbihK02sLxGFaCIYPa2d4VsW5+eYhMshiuQVKbuUJE
mCstg+bFRGGpRt/Ug6stNj0ZXidZxQZAtKwJmjy/P3KT0pqN3WnTIpZrOW+KHZvJulT926L2qXNt
7XL5FFG7ogNnsqIJ2IRqK2Cp52qLRi7pPHnBlG/yVvxPyMKVoeUKlzkpo0Pj9/XB3FqpYMcUYkMD
D5euXEfnIAdfy3fbvEHpHyaXswAbd1OboNC/xdK5zC6WWEmQdMmxki4EwxLrf2czUH155Y4Lh+TM
FTzY+gavOCyrMf6WeJRUNwPknUq3wKZ55Hf5mIkwcrpHmjD8iOmFjN5xkzxFlC7153QZyc4cjit1
MHHCyqLT7AdVZ7GHnej9JaBSQaji/jGkX3gGwx5gMK3WN0s+Os8vC1xnTSvH/0vXZzL0z+aSHbRh
20doicQAY/8fawvewIodE5vs7OOjNCxgC+o+Ve4RiSeOEcIUyCwAN+FAXalkkc4RrU/oU5As50Yl
T6+4kGOoWSn7KcZXnLpoA8wOUhQXcP4cInFkx+X6/o7wUlBiIVJ9jWqp4JdxOx/G2n32QDtRioa7
cVWrJKqxZrRZVDQQ9KkIzSmZdhq+xijSRMmxmAE2F/IvLOd2yAjgpp1KIS2uEQfl88ATV3sqwX0t
hB+qsV+zInPfkEt9wFlDvpnvoHLY1H5J6oaHSe7LUULm0CZi9bspEPF9Bwp/AI4ABWDv1jfWzHMV
Bl+M2Ig6VHoH7XqDvY8BQnAfGN4hFEL34x6D9t45zBz4CKPYZ7evwkOQ6Ab4sDLs9BBsxIRu9JNf
8sSb2LCZPp9yARysTXiGSsWreAs42N8gkQ5QGC6s2dHftHGrNC7/5cxcxwd0HrLn8fOFgl+ONQ0E
oQDfXbiXvQtdLDWMetfBvXBKIFIpD+nsarS6D+sLwoZaecGTvN4F+WzUMZgM7Ta4lyEQY/YRY2e8
auZO9kFQEgP/mSfd3wJQb66S8TJOqZ/QfZea4HK1AaRCTfaUJnldRW9OFqJJZLXKwoqhg6xxN93U
lZRTu032/FqXpvr+iuaNOZNmvpTXLYU6SKdRpoWLzz2QHJxsgXhFhmPwtcfo7yK9hzCJIEoovZRl
DW5wOJTQya1pcj+Fc0JpQTxAgNBFE41H15BQGSMTUzNNy9Y1Mm1Cxf0MRvUOFSKR98kTRYaXpIK8
69xpybeqXACCL/8Qk2nfnl+r+63RSblx9RqohPZrSkFd8cadCwfrXI9GMPLK4GiqLAx0zkxNoQ4v
HP7XCfM+WjA5ej2Mn4JxSAz8zCn7NoIPmZVQzRS7cN9420phxAEV34fOK3XbE6NFkOhjnCkYN+DX
9AhcP8CTf5A4FvPBo/NqsDCp1+vPYQZQeWBhncYPMIkDpTSt96vGErqFi7oubIuQ1075vJU/KEwf
O1tLxUAoV3dNT3nc/Wa1pLNeoUDnqjZv/MVLSYgeJEhrzrCEApQ5sK58tK+cVThIx1H8QbcAuqpp
axrYxSxxAfml/526MJp8nTuOkWsWSArUSdOn6CKqJRmAK3q4yp3l6YRUl9mfxDv6BsNWPIQvuhI/
KxEAAd6K7+eGK9I/Ilsb4c3h/YkgLjovKQIZ8HSElP/ZclC3tLkW7q3BLH2c5ycRVjoMVfUecdHg
HItVHEMhjHJbRLX5+783s14ni9shPaI/LBZSqrm54vXmv7Vll+jp0odTdlhGrw8ms0r513xNX4WR
uif0LVbl6KzEZhDGjgp2RlBWEaDIOeWGq8iyaKxZhNdaOMgnMlXgKFCD2qpV/6lJItAW+tdqLNR4
NA7eeaRSere6ZVGoFSNjS17gBJVOijSl2QDXtqRCnZsEuZxexXJI7GK0S4MtbM7oGmd2zSb/AKgZ
qymD2CaIMC6BWjs1uVZlntx7YY9VDIGYGqzikhWU/ceJxBzS7FwGGFJgLrtgi48Fwz+ijnq1fGWR
80HcicrjDIz9KBL3sRrXNA/SvPI1R7UCXWzfF4hKDgtROFHWNZGFT2c5tWj4p7fBDYobJ7ZoMmVX
EqwNAataN5HZZRPdxhTYGxiJvNfqcnRcl2IZQ8abLK6wQlZmp8zWP0Bzjxv75D6IBeHTN1SGfA1t
ICAfZjlggFFLVAbagmlFrEtXATxZf+XSqJdCWH3Pj87pfJ+dvO1BWBILwsN89LxFv9c6iycaTI/R
6LD2hjcUDOrimRrVq5a8MA081j1CrgNm5mDH1SnHVagB6KcsbdYFFJO4QrcBchAeg2n2tLeUw1yc
YyNHdgxuYK9K+WFc8GxkM4JNT+Qc8YRSJzfyB+UtmM5agHyX43Iabru5hSRvbNmSxWgvcaj5JNzg
+zJYwrRO9Q97aLnnFV+pNPvJv+ap2zEz/ghR5yRx311tuo5WuNKU0dfYU+KJBqbHAHSDRVIxLzoE
pDqEutZGNgLy38t4n4yeVujPn78OsbsTPmpIlHEWz4UIyNjHLjepvJBgfnawMd6DXKzSK4g9OKuH
+4vBt97d5pEuwBYan//1otMIk7zXku1m42vnv+i1tE+o0upoMebhOg/vCU3osEuYuAkJUC1Fyb9H
HD/ZyElMfMH6wbOPwwH09M3yTl9vGvj/gM4QDIKR5ib3TbuvG6q4vGAAm8tymkkYPRgKW9D4FcUd
y8dY+c7aovltA5ZoZ6MmliNttwzBj/Uc6uz9VHrHycl7FI50MMT9HCZJQvpYatBm+lP0JbwVMhKt
hJX1wf5mvWShqv0j/wCj1If27/e4Xcxr8ZhA6l7dht3YSVEldu2B3wOBJdMW5tToibeO1TF9tb5L
Z4LsOsAZ5LReKFL+p8zd2NuZVKWAUjWrSeWlI6H2Nxhz74NDcV/zJwf0DAiQ64JKQP0RRRmbmvpC
GGpICCzpfdT3xdhhvR+NxwLNXwcJctbhdIZO2E7fPI+9CzLGFHxVE/NgR/b/GnCVWVKj3s+dSQlx
8obOM9ZXuAEiaio+gYC4fwJMlrMTopGimzfLpLBChTMxdB/MEL4iy7GOA0e2PwVsRv4DFU0Tta0p
h0YLCFHq7Kt+8i2RsMjT0kgwB2jMkBYcpKMj9RmuZaOkJuQoqKFqhCAAtyFUTWTvrz2LFnBsFx+H
K2mAfX8bBzLKtZS8yYmu1skBF9ht0UsjqjfJ2Rn9rl1oV4T/Rp/swI8RgwLorvQDdjv6oycdPgfr
NKvPxDLlvoMhEdci+y+WFKcAhpxace9lgO5lKDts+dGIfpH4vR3Iyq9zEwB7FrIKcBtCWPdjK5vQ
gX1gPtbagdGtJZl2yPQrAOjqdt7NBdH0QTJ/BbnJ1GjAdgCBqLKsakdzxavVzaAxF4fyj8L4GEDf
gYUjI9lQKX3LW1DWMcT8ZH2Y2cSpuZNjIr7VQ8sxCOJRtZi9Gp/TD2EscolM+ZDWQwA0x2rBHwMW
JGSvx/fYOZXltpUln6s3mZHmaqdbirPuPqqUjtoaOuu7q+aPrJwJoXeub3BSTkDW0go+dHsaBOS/
iw0iu6HQSXfzeaX+/rgAoxlESKVoYG3WpwLjk+Kj1N8LB4TMkgi5ifWlBvDR0OxzhdvUdAJDvfuV
mddE3hnmiWkHLWSjhlkyYvAKrvbb5PD2Q1d6E2Dg2XAni+FHsJ9fbg9hs+OUXqsotAVFJ+r4TeL5
CGgyKYgE1B35kJpMeZ9pBrIveBBuecayylZADUaDFY4aPsEecL4bWQPZ6Pgrtf7+OL9wp03sKJY0
EM+1oKgkeWLWUTxrwPzmoT4sEuTyJSYYlrUrjTtjSKvbzH6uCAcyHnncAaHRRn/8UJt8v9GrCu6b
0j+JnNgP4y1elZ6p+BvcBaViavVCgSEC+P6udDy9j4XngAxP66rBbtx28/Tecal0q1APyR1iLEEI
oeVFXbTr0KSf9L++nT8r9PDutqGJAK6zs++QmaUFkWGrlqROgTtotQRA81Y+ToBThzZu8FSl3fSY
XBA09UKHO/uNappT9KefyfJtFPUCjj/TvQkigzvunuJq25WczKVqAR4L6AFtG74uXW3jE6c6UDI6
HqtKUHOfW96fwATFdqKGTq+LwnbvkibPYAHhhqYkPWlgwaIeFrTgWl5MFhhZf8oycoX5KtuZBTb6
B+JD7lXkUD/OFoeLffgHbDir/shGFrjeHonJdNnB3XVtE6VLYTDQ5VqhruaxXZbruH+CIV2O625H
UBn9EqDwEiMdzgPvxd5x5xPq/UMUL61ydfuBiY6O4a4hipRGGs/Btc+RSUXFgWv5DTG+u8OiH1Bc
nB90RXQEIR1gCwXrYMPN3gSL/wBV0H1n5IhUMfp6HOxSAIR7FPcCi5iP1LEs8hV1I2Zv1TPNN0Nb
e65sWU41Cpy9zUoa46tjbcuUX9h/Rkgi+iUGprzuLNcURoLcMDcBVuPxOdiK44QZCPD5EtA/hg/x
T5zrReKMRtWWdyHe6K0aggmdswZd28M05y4+lkBHJVbGtY3SiQjGFdtFDrliRNbR0WdXrNFYQgP0
zTdxqf913la5IcPd25HhBAhP8UmbfZMKlKeiVkF2FADwmYxa36Nz0UVuhWdPzdlfrzV9sMbh1oF7
SpaDd6mHCObYUASYhCV4pKwPJaZP/ynDOeIeD/8oLVr1887XuH8YA5R4of4a5fPUYL9ot15VPX13
03wlPuFcXlDG4Cm3NlxGeBUaVTiqtK5+E56wzIzRU+fopntrglZFmfCmy3AI1OalrUlneOV8U3bV
2M+HwPE2U5Q/U5lXFAu86V3otDSNtcmwUxeK/Ym8EefPghoWdoMNpg+goILRCxAZFzjoK7v/pc4a
Yx7rqj4FFnx40xSwo7FVFtlL1ZV5Ek9iDvyYO82nXvMapH/kHmOX2ujNoVbFuXujJChQVpNwJG4x
3DpV56FDgtazRUBoLqg/NMwWvwpnU6mcu6oPq6re23tffKPE76He69YNGXoBYH8ad+KlW3g/LsIV
qMREpry7mZzK5pGnZrYTM0to1bvQ6o0mQP4S0kTrxdWzVyg8fNKJYTP7J0WTiUvt0A2Owz1PRTrt
xTE7vyXuxMieJ78u+PCeNKX73PyZTx0m52mDrS1jnvp1cpGQayY/xQD5Z2feJiRgGaJcfbSHcnE6
4rZHHZb8tnWSxHU3Yc/UddPkaUrsLPEpmxKwYXPFaJYoczAL3RlhIpCEpSoKFhw0V2sTCQS7WWG0
5opzJmkJqvu1iKcS2X47TccBembXGZA3TPMwY9pSIgi64rUxbjjco9vt2lRfUDCOE6dGM2tRdgyo
mTyEZEhjQTvHRFqBkojViNqIXiEoNzIJEcqDEgJhpuih1j66Qv7n6u9L0irRCwDmy1ccQOyiMYFl
MNcEoyHPV/jUsE+yWUMpTuYtGBC21Y+uXyneOdjIESCWD8SebKpzc6dVAQTQxp7WrzeYXWaBIG1g
lQ8kfl8C3xXLq14mVvHkzoeORS4LVGopAudcLcXImLa3cawb6bywNH4f0sYTVn0rA8I1yPnloAb5
zyJMFK7KvOzPm6HUiwQ8l5KuP/ctUvijKxX3Yk5VEiHO2tD3IYX0M8hck9k7+958PRPVIIYifzcu
tV+KY8HuoHp5+VEqKezStFlZ85KLR3jFIoU9ctQX9MOwvRX3cqm23rO3oVt/9Ru7/k/rTeaQUuXQ
UnNblWnqIoqGDanUMre1xumFTGgRg8VfJ2W2rD2nZvwf6U+Bp+3cOn0lyNW4XZ3RQrw9tbjCso3S
6o2O2JgXHkfBIv+eKUe2gjYtgGUXN/3bTDWdXwCi/NKFXt2x9nBOMyI5NVOJuIQU3XSfh82Guizo
H+jpmY6tS1i2wzOIfm6a+8SzymZm1uPgWur4oSnrOLoY841u611Xfkrf9zgB7ZUDqlz4nLuBRw+L
15NbrpTjRoecKLVKNt1L9NpWqI+AQflLdY1AdvIN57b2MyVpfBE+E2m1L+dx1QeuBD5YbropuaYM
tYG+B1WVEXCIVYUC0ecp8Tpka9Qn5iO1KU4hsbgPQXcTtR+biEwhgozFSdXBKWtcXPTsuGxuCpxD
ZWY53LBNV9qxH4dn9v8QmJdVxnfZVr9gCVSxbztqpOtTxSjSELUuzstozyu0mGG+DXBmTspnan2P
zioUMDNnT8JjY17nmUagvsjkyPhPtJzfz2MF6gHadbggFkSG11d+kC/lsVIQaIi9Pa8eLCgOCGXH
jXUvwDN8X98V5pcddAt1j6DxpSvqkeDY0XVAjzp6WTWPWSNHfNSngGVQQhAhalVVb0+63jSBuOfh
SFYwxtPoTNSfO1hCuyST8Eq4u62RFO74h3+tJSQt/esiRNd6ZIoCrwSdn4oGPVYWGdFy4J3rf8xI
l8bsO2RxxMT2QjNeQE7vYLBtffIpanSEhwPYslhSAj3VPi2cnt4U5zmFk7fiGMUGy1C6WU8Vgrf4
fYacT6DNKwzx2nmJfTCfdjrCYRLAFhaR1O1XLJe9MPxmZKW70nvJaK9rTPl5OeUEmzun9J38TCJL
NJTEaYPCuwAnqGY7f6roClki7MVCp84NTXeDqMmYpLyIBGGgH+npjkUzhzwaD8YUYCU3bxMknNl7
U1ZVd8cIJrmTbXp/ud/Hd4hJyyEFC/L/xUiaEToXOMIFXS6H7F4FyvvJaZNK2YvnMpxGneTObWU9
yo91gZ2aNvck2cRKuOhSA6euKUCEOi5qYGMRo2DvNH/ETyqcjO+sbk85nFTpe72MoZ1PPUJI27r7
h/Hs1VKp6XNGhtTexO6T/bebggG0HHbTt0TpxmUUimI54JQ9462kS9s9Tn7M9/EGdx0QkpXbjwxI
79zznO85J2z4LVVUZ+PFxcK44SW4a1nSoBSDFK3fDQIkHIwQZDOEkp5UFSDiIiB40ID9Aldysgoe
tHACaziLTtNd332fIzrJFYfVTKCdCqU2tR0VZ+wix/tKVJUoojM20/RUDBXshkzaGGuTu1PizZKL
iXQBuPCj6gntpJQ8pOBQSJziNWFML0xhxCFCmoxT2Pb7XDby0CC9cUGNw6sEduYlLRZGGcvaNMzg
IaLfrjRoXQewiYSbpvPTDxcRNlV63CHhDnzVm0hgVdnmcx2tx4zxJ0/MBqrmCA9sk90RPgNkQmp+
KohrynwArcC9tSUzyys4e/S6dSx7swaTLkKYLSxTBR5/H7+KWOPG4zzPc22Hg5Fjb8Zxqx69HPGX
Ly7Q4wFG9qrxT23rKY+uYF06casNC2aSYwOmyfI/+zI++qlJMcA+MMSxyb2vu5Ocs99qt8Cos9cB
AguYQWx1Y7lP7drIIkDVlDkCpiEN1K+B+txO/019dMvSnvSnn1EMg2MO9mcQ7B1kYV7whVRnlfCB
fNGD2XONB/XyfY629ua9gg63hF9wk1a56PERvg7LV70CQmdA21WB2VsWy0D056y2/GnkWxHFjQXl
4qmf/KuFy9zrShBN9Sx/aqUilk2ruD9rO9BPFvdy0WEbNzyrzxd61eFjYlxriQFkA3k/dBu8p1xW
wI8kbRd80xr5Y61jCTVXq91j4ogMGs84YahmcYm9B70LB4ZQK9M6vUqGlW3x6UNYtwcwhRFmkppQ
nByxCjkKdSkwLrMnFegwGc9H7ZOfCYFn4jxe3ouCShU5n+IzdzQ1vN30eIMFpvwJvEzvCNfBcwo3
PAGWfwjcmfdTvwhdEfmu2AoxDMPiLvT115vlsbQEaGJR07vhy/wugEpA3715uJ0IZblrIaOAMDt4
bttstZyIQj+uReOWyT996tPu7bWRM2Qaz72CfJaE7X5xURX1p5c3ToamczVHTQGPX8akYxaVg1ad
JcKfXAo4PP13JSehOfG7dBXjnZqFl3x6eeZPHDMTmAMcjTeRux6jtU0ahf9r+xMmdm8z2YUjF+7s
awN99MttOsueLJfTTPZ2WuWxhdH3dKxXGm/CEAXFZJJpc34sube4fLNZTKvDYXzF6fSIo95FyOc5
rE4BNeWKFLRHh64vQ9V31DzCWZLOAiAaVykpDZdRTlrjurhVX/yuzBeU4xDKgFjumoUvLA6mPudA
SDt/oB4MHe/0uIZ3O7GZfUwpFviaCOw9pKMadqrVNTE3mx/Lrg/6EVvUQB+ynzBBN+e/yUWZSRMl
PIpY1fwV/pkjcq2TZN4/jcD9WBZ4FzwArEXvn9vzT6Ze8dUmQaq/mgdqEk73V71GM/cmQC1RDa+G
wxkTWQEwafao0b429jwwMjKZXTHBNBG1p9U74/5L8ruUD38wum7i5QquiIa/Bz0d9IQfOKYdNJpw
J8Sf9S5KELlF+SJDu6/BE7A/DlWr0YdLdJAeGNv3x8Mp9Fp4xQCKJwSQBFrhtOalGIslzWvXOGYm
vuf1u4lxd6VFBRrfEeMUuweLKsXsE113YPmMhnsxcwYuvF5KXlkb2akwZamH5TB+gdAFtxFk1V34
poA1TuwU5+SlXcoP130il/PJYwedTyWU5xxyWBJ9YcOKsi0fsSJLSfjTfw+d95bRzIMFlqS8kO8d
OOaGpIaAzIc4+ysKvjvxBfrlCS/o/+1hchiACnl7SCVcKBxw7XAL+0LUNKAf6R3wkm6WJc3OQNEB
C0LfaJdubwZH80SNLKMhrt3ZXk3Kf7yps6lBkBJ0WKKwbVaix/2WkkNkNfoci+R538xJg4OW5hJ3
OLBEwFSRKdg3BmcwxxF5eMbOshpnhVVN2fDvfO7eOzhjHgjZ2vHCTZgz/KnUFPf4fKqlRgaGqYO2
AW5USB5R/e8O96gqmRLQMsCKPOa0eUPqpuAfP8UUZnUcbZFKncSmrU7DSVQrOiNGBIhG4+p6smsB
PTWw09bKMW35W0YuYbQyVwo8ol3e4qOB1kUwLJjzfZgZGqAlUf0nNqMknR+JfWO7P4F50qTXdxE0
Mrhb6rpE14VQKypKFXMnQ5EyV09nGHl6R+bJD8vPPdIpPbhUObxqFwRxsLxtT0pN613UbSOoBmMI
0ty3zfOclCFDQAtZbMzgd1OHI7+izhx3UVMhFyymhxC+quAnhSZs3K8blP5GHmhzO17uybkzsXhf
hc10cMbjIdTVtXDsrEaIsQdCom/+g2S13usllyQg+aurHfM6KjUjLCvzOnJ3m6DqQKMEXsJzHFJo
WYvGuv6fEWj0PKLbCfEDvurG2sa+4jpuVqfV4wa+UAORhs7ZphBlO2rL9aEl0qdgStEV3ycaqOlP
DX7JuEIx9wwMOuoQ/seaV4aej4WfrvgW5l1XsqsdpZS2aAzQnh85lxm6C4EJhDac3457GKyjNhy2
qmWMoxiZv9rpV5ErEtGSipZiPmHR1fNjUPhHyieQLGvzK5oBdcTbHPR8dofXfFVCIxTGvvrZlXAf
psiYrFirastiexjA801d/FEwJa0w0NF0k6kaeScpMAZ1FO8BU22b0sIcT7P0OmiaH/oAe5WFrra7
7wUe/xOqNvXETkjjl3qD7e0ZTal6ULcd/OF/CF8ymaYVni7/9JVUb7/YXjuH98JlOdqgrL8tYmfI
bhueAqWzL33p1G27GZKc+ZFx7VtIxa9VKwSExdUB726u7Zaa5dPcgNZwKgqm9T2O9z1fd3mbNTSB
gCPO+JgV1SAMndmiVphrPBOG+37QAEQ8T0bAq3BZpmtCQcOAy1owMazmVvHB61hDRbqC8bHpKRgd
F2hdB7N3COXQKS+jrf3l7kM9irsV9eF2gGBZV2Rsyv8YIa/4fxRJYHNRosAnYIJNy38GHkTD+QdY
b5u3S0Rdj486xcYxKuqsZVeqpzxb+rAy/alo3f8lBeERPYeJuJ/EAq7aN95lTw08yoHUTFBecf0g
NLFKiXs6brqSb7LwH8Jc8+vAUSgUbmt5sPUJRcV3nmZkalR+gmMz2143ahB0l737yfmUyfBBqn4n
FVv2nwpeFE9dVgIq/Wq30l4MtumT+9jxoAy/QxTbPqbkRRd4fj4tJ8NAHgo/BI84kDie6lrrBSKG
dKd8qdG/Z0xgviL/zCERwFBRj4ZQHy+hpnJT1zU1b8S0pGYgtRZ4i98HhsdLtydc8sZBGwN73QyR
bapk7N8mNXfHxVvSEfT4B+VDRcrzPllxdjeVXXjp3SzbmLbxys3thHEQaBPHN0Dm4nV2ZFd+04aK
IKUQfonQCgvx8rdUi2GnXP3Kq1xcNzCsF+IMKf8Y/4zqBlJKhIUTvDdbAXMs1InJTkHzCW5iKsbQ
lBpuivf8Fq1HpI7B44Lkp8J8pGf24txtG/YEse3VtXQAumtu/1Phkakw3i9v/1mF/KYmlOgYEpQg
JOzPgdOcQa0wLmMqBpHlTeEJMAHN4g+mfECzUiUC9ZKu2+cEFricHOwUcPkdMRDJqUA/4XRdfM58
/LBHsUM/bosa4U6KqDA6CyulDpnCadokNDn71iJvryiDB2Ug5UiMD6hXFp9/5qbfksmEtMpi9SIs
FMOjyQK3uA+a5xC6uanj5T5BTg8u3W8wOTBlUyiYD0ddptr+IcFBl5W2HCqzbI1oCtJ7jO6zHfSr
n1CZBcZYS2RbHuk5NwNIUEtW2+kWBa/iu3bF0Ritfv62E9JVETWELonlFG2pUw6gpJ3LOWbRmPZ4
q3Qd+YkiT3N9GhRfaneS9zH6YhNE91/1EoFevQuYRrM5mafRuBtkV+LJJCRzg17gLAPJfJ8eDW7k
qcl/Sk2h43Ebtf6AUDwiyDU5MuuiPXndZBJyaUIX4/rKFRiv8VlTvMXL5bkEOhS/pTlc79scYbdN
3P800iSoUENBQzL3JlfELEJF+c4wGV8Znow4LR5ztDGhF21XAZQpx3N11CSL697f5pOiZIBKOmKh
UXQbZqChC55EpfPAP6Dq8pEgH1NU6hq2C9J1DbXlob+ZgvFR1b/sQXZ/Hxc3P8wAkqhx2rsghdpa
utS8IKNwJxX+CtJBlxGORa1420eRn3Y0hOKYawnSwpPrNV4Avh7asi47yxr+6VyYxtPAJQ13N3Pb
bR5FsWhf2gUuDEa9wAYVktP2zJzIC2QU70las4SCXUt4PiFp43ur63qFaXV4GsNMCRzl4GiewLwM
3zPRU8sNqxs//hZBSllMl8pn67Ai4dXf7PxKHobc9vKzch7B6EjvlrgDk7ecRv8QbBXWnsLIV1tK
B6u0Wpn43qbAs/moBFQfjovFCLL9v+MWCEWZ27H8eRDUH8ZtKM4v1KyCSl44HbaHzLWWHnpxxd8N
AsGFquH8cuNEjUuoNmbVGMGgGv4lyVpeAjGOJwWm7k/XL3p9Qrlt1FaMfkvWqRaNJepDvlVAQMDo
JKx7lHtmzs9RteCYWnx8Fl2sMeQZ0UMr+D2mypZ7WFYaovyToJSW3V6VqtqzgZSm7t/QeqAAEyT0
aMS3dQgwpZs/3pWevWztpbAyzxKttElV7mp0sACWH0mD2rJWqd7tOW22wj0YxGN70BEZbi7qFgT/
WP1wSTDOlTir7x4mKzmp6sDYtGM7aibYvNIDzoNC9UzR7S9VrDPbW7p8DOxcFbnNEWbsXDoe8HZ0
jl8tJzdJBYiMcXearOgygcqJyTashaG4qSw+IFa8AtML6V0/NjpezqOfTZ7T/vTvUPKE8YNAWcid
3YWUar2rAEYl/t3ZYz7ZOU9DlX544qbcBvaIJ9NwOwsMEhPZPOvU6rHB23KnND7UWLj/EDvKy3O5
cgrLoIJvZc7J/5I7D8eHcwyh9iBCg1cyIv8q3XqsjSe4KOrQh+up3FKTwfK/KAxK4cTZwIvlPKcV
NMoq+dz1P78lHUimYPfy+k+d0eqdGO/d3969dPFf7L3qZjsQeV+NuCrqxeDRQM8JqCbDeknSIC89
3BcMKFAaaC4FipkSZvgOfnatdCDtKNq6SEHS3qJrsvH4BRhfC+ihknSUUI3pWdPbPOs4JqhjXwK4
NVPgOdM0DWdKd2UBnXC6YzT0itsa420gNW8r4ms5KXOR4KlgrF/T1At6hRWNo+HWk3SMhtqUat4Q
7NpfEmOZ079xoFsPq3NkHe6ZLC3gu43BN0dvLfIL/FHkBD3hp9mukiWlJgrYCStC4vK/Zi4+tDIq
m8rz10KAKfNB66Wt2Mg1CCCulhF0IkoB8U3B7T5ht/YKVvnliPSE1sLiHegjYa/Kh4X5Ts7fOwhn
gy6tikShgvMNJ9TYZLIDpilU6wAP8yUYDSlWJOnz6WPtuzM6iZ9dhUCoS9Mz65w04Qnc7SZs7FuU
79W9/VrOuLzN6sgKUoaI5x9Qp/7FcrcEBELWcOHIRufPIsrIJQfVjo2epn3eO6CxKImGo+ejTBEg
/Rj1jgus7ixMeWQdPBzPPGae5SqKq3WxPEQVf2UwOO2cn7nEv7bBf1N7zglK4ayW2xftALX+aduy
Zquq0aafMD7H6foeHCVsjl0Ha6WmgVliboY0rh14T10WjP8F2hLUU1ahfSf6DYvL/BiHkaCG+71Q
6RUrOBdaWGEGzjhgFZ/orA0duMFwQOxclhOZ85rqy4qT6LP6LCMrukTjNneUNEkYu/K6SYzFLbyr
FxAWjzbxkiSgdON5O+JStCXkrnHrYMDgIecrIpQOoZb7lEp5UnbeCmpL/L2W8Ho7/MQJIubk6LVu
1WEei0V8vmCrrAdpqGPI7Z3JEjv7ajGXZ6oKwTXMyxI35nJijOrDbtklffaearHgla5ufAAfwQgA
rsZmBwZC/wuMESxwE/KmowADD1BxHSQuBirhVuQCj8acNean4qCUZ06wIZreNX1DZ2BS2wGWPSbV
dmrgVmWPQTLA/IrUtj96+0Sj1H0V8+6Q+ARtUGkc6Gr9EcITx3PZTYS9g35LuGk5xIjSt+PTsrZa
B5n/Uw5yZ6TpHrGkXFStpvEKRseD5UB9OznVs4X8KCGcgrX7yHGuWl44FjE4bP+dUoVFDwfssGch
Hf/ttbb91rc3cz3DqglTUQ9c3B9IBtuewVOZogO4/VCx0eCoB8MY8gf8i+85P1omMcj9w3UqwJF3
luB/u5QixHnZ9oDskOYAl9ZIA5cxfhk8bzWe70mNyIjWXAjouTyYK6Xw9foKoupt49jaj/QEDKfH
vb2Q7A103PwlNmnMnIIF0KDbRLJASPmpwXYzfS4S5rGXYoRCTaSrvT8wA4iNh0DU7gmBQMXO0DqX
DKN7Eic9fIFN3VnGl5x0TUH2X9H13VrFJ1hEESQhbAPmPyXVIJplK63zRGvjOw/+wr3hUUbhQoZE
EQY6WFeSsos/wTR7zueK15NeVpC3jfCE6WCbZpILcZy2HSDR89sMbjBphVz+fCCW7+FJqXB0VwfG
0AuEeznbx+zoiZz9xh+Pvn2jGkp+zgpiEbGWUp3LZ3E1CUcjYUDafXGxYe9As5pjRyz9kVzUCQjq
ld1Kie+HHiKu7kzQLECkE4bxygAS6kg3CpmMxX7oADOBg+eSIH+m+hNrS+2d7lO7tMtwOG97EdbI
9qroHca7k2d8+0GTR9InEtu/j0hiFnQvfyUPP3eYbG0T9T88d9fAFDc4+Sv2eGVGp0xYezgECKh+
3kw/BepnAjRxxFAlwDWcEsR6OtqfvaPMTajaqFerIyVdZEmAX2nNx/1tEAn456HZbFeO6jnDyg0C
gacGPcn831jecbC7G3WoUD4joG7r0gINAtFwi+0AZqTW0EmQUZH+9bzAXV0P7WRm3xrPDHjMGzKI
WrlvclA/EUdlRl1Q57RT2Etj9q2GJbXtSZNLWIMWT46eWVUGK2HEXYb53uOctAlRIw+p4xQjTNaD
Zj650jEBLqtyu2EFGD5mdBnGQDoWn+S5Sw2guSlj7w5W1tvafRedP3SKM+P6jdv7sM7zb9VexI3S
0xwBmFG8rgFGo+x2Zcx7tfrQcwjGHIGgJYwraT/cd0v1UaATCeVLlLYTKZZg1cc8t0cMRRLGBH5V
nIYarrJw88iFdpKx3w0dhlhxc2oB4dtKvYhP8RZc2cJ74NpGRTelXqIW2s1HOVrtpdAteQ5X5chw
W2V0QOSTp9LPASacuT0QOqbitjQUjTDF1AQnCB31s1l1MAc9zJViRcg4IihO5dhevCAokJmQgdp9
rkX7cDVMisXPUmQtjc64pOMMXamJeTEq7FxTZlaa/TFqZ+UFC7WPJWkdpHR6HCSmaw0u05v7fD7r
AbUblIG8NAIbG7/XkZEy13YEt9ZYt9gCZqvk6A8KM8oZ7+b2jv22Z3MB6B2NLAW/a3abwtZVLsmr
RLb1OKO6L35iginZJ35iZ3jmOazQ0TCu+qZVShfwg/SsEhHG+2BwSnC1Jio+8VroKogaTgZNOsLq
Yd1Qw7exJm+xtu8Nqp358hrJx1PWppUwdi3bwTmCS8LyU0rmDhuehfofu1jRaaNXuODAwcmejXAi
aeKzI6NqUBqGPvsJOqsLP0Kn9D3iG8dvOrz3cJVGcLZLIDzT5WUMD+LAkNzhnyNGdybz96KxPv4P
s8Qhj8Iq7A0Nx5D5PK5ENhejc96ha7UGL4vYq4oHYbFnSWqW8vNIFRF7RZlIf5ljD2ew2+iNuwU+
UwM37ksOpnHimS9SjWOQOvtudDM22ChYbvN2iTwqJ3LHSHga8GzEbeCtrzzA1XoChQcBQgOeZyDI
N/holSIyws/lJHRt3VkkbciLav0H2E4W31A8NTiq5OaLYMDY2fD6YwV6n1gzRQbCijvQnT9Qv9qS
aU7PEaZL6s+hQ9s4gDrFwoxsROClxPbuBoYy+K0VxV4haGzvS9bCJY4woB+KwdKPtmeJd5t7IIHT
8irUcqLRX2IBhc3wW7CKhe9mnDLPk/3F14gTBQ8JLvljnckSFjifjeBBuqtA4/xAjrPO3wM79G1S
NHlb8DHwzrDkwqC3JWA1jfOlBp0xbeeCESbqdrefFmUX3IKt8BTBafYYCq1uucPkya5h2oNVyIFG
r6lcfXeQgj+br91fYkDjoW949B5H1vbWW2h4ru7DZi2da0ttj0/AfLm7xrgUkfo6Zjlwn/V0egLF
HW8nWgmqAcAtde8y4/+A0Uum24ZZ1+8zViAcd8H0DiwB6/oVRFeI18zbhSXtY17LPza8rY/Sv4mW
G97rMBUYdRi4RiukPnt2j0fZgWNoQC0LXWNVtohNLjlxCxn5I5JWlxwG78V/LGflGHSPdLDqRie7
CVtkinxru6gZzJanxd0+seXMvaDqKIS+GK5wTX+PDLXGNZS9dTaOGnIzT+WkUohMbbmVmovlUk+8
jQHuboVXjtzULagLI6Dmjimg7ervH8S1jBGAfK+Lsfa/ggdt+j64c1bN0aarimd4W/ToF09ezbAL
7z4wbxFeO7KbusO6qeBUbs2XEhKucsgTRJujOlzO0eC+apUlw8suN1D1d0GeMm+07iK1wffmrtzl
UtzsWoDF/dNMp8xlRo8QqLPzGK111tQN+rZgtvVYyFap+0et13iASGkMQYRu6LBX8NXLBqex2Atb
kNkXErz4zfnU4Byhl14DWivGL6kwNKGc1b2Eh6SbeQad3zhg5vYgDjJQOLUmcek7sMAh0reRVvFC
XEs/LTe+oL2KaM9AKnhVHQxQfWIw3J7EEdgtMUySf3uPWYAhRwUMZJRrP6+0AE8/7S2s7tO4FvPe
bzhResUw02g+m1aKpz2WU6Sh3/EKF+qIOu9lTlDYse4YC9z9gFU/d23ddUx1WsB2UvpX6HoCi3c+
a81fHQTvuLmEnJvv9oCAi2B0otYJpzoMbldkcTWLl5UfICsL/hBPQaWFELUtY3sB4xbNtqaIQQRM
TyYTJT20rEvfa+kHk9R46Wt2d2sznGvej5Q2jYGE+scNvrj/GWJCAFNEjRj4t1l4mkOmWI5/I263
aeQ52qiuB94o0kOXbi6ct1Ko5YL8wlYrbu+VWPg9/nCPvQgxCExEqFN9of+9jICBpGpCaoB/Gp1w
oyVW0S8iJPVq183KJyCmcBaD2tergHbIqvCt98UDqUNgMOpcWAMbfVtLnPtrz1pF1wgYfvDEdCbX
LyoQsz8Ut2atVLJONxM4vMQQe+I99xMoDwpIB/RPNo8n3QXTrwWLJcMmhlfrCC4PBkQf7k35FwzS
dJ+xfONjIOu+NZmjFrVWaiRWwf5xMhGYUHjSBgcMXb0GKdlwVgZcs4ivu2THES+FCLYFF8OKzzDD
Cq7GQjkGjpNocu8zH2733s4WyvxnspAUHefVnyVKmBrdmVJVZ+BHdaZbhMBHb2rVot6KyZ0WMlYV
ij6Ss7v7EfmLdKNKMn+iQ4jZ/775XWB82LeBNz1/01ykFQOy3EUZI+6wEqWShmQWtoLlA+5Hlf6D
KG7SebaCWYWWDSGDU9gXLQJ9nkmb7f6KfunR3RtHyvyW7ZH9i4k/9oOjYwCfyx9UexXMnTGVKgZV
NydazAfdpV3JoZxDwo1dfEYRBg3k/GyWTpKAgxQSmKWLBie5FW93VhiV9tMXz84TfPqoWGtlPHZs
gHhGmhKzjn/z2WSBlZA9WhA+2VmOu5NVigDbvYOFR1tvbgj0xDEcTXOGfP99hcJWK5PYSCKyKsSf
Ib4cDAEO0JYQVWk9Bb72sivqI2okGKkUb4ENqXwH9GKIkEtosAhQ67YBi7DIKXeprGEJlK9fjEKE
LjWl3CATxJg6QJ9/CQh31HzNOYunjefUq8CB6TtP3LEg9PMNt4RgdZM4x/UvwXenCWQBcD+uQdOa
1rJxK4hBos7mpSwiWFHbeXcXffwuPIq9eKeF1MjxBS9pp4eAWT393yTu9piUGs0iq+bVxce32xIl
Xj4MSYIDUFfVOiLlV2F42KTvevOd8xvBbSeVPt5rFko87lz/c7j0lnRi/jNOLTG+rzjzpzJAOOp6
2UIJIVO9lY4XF5Dg5/p1PwLxIH3PRGUkxiFphebcMgzZCHuCIa2Cp9HO+VVj/wTDel/w9cVy0+7P
HwU9ztGzTahjRCV61UaF+QkOS0om0ztjyNo83p0yvgtGcq33bSuDUfWNSrPa64EilGPZt714SYLy
k45WNd/p9W4FgGsoPPEPqrX/4s+FQk0tC3rDDHPgTLw+WfDZMT5qz7Gi/jEU0KWQzNE/eYbIzrGW
EArtwOaOzh9HPbUZswaTNKF5kgoblWLEj2bbVXvkaZj+R2H9H2IVgYP6iOxfOCHAnv+orXz+5oM4
edP3cN46mohnpzyf2/Hg/h/+Pfkd2BzjhQwtFq6qf5FCrV9SdtLiMfcpyzVy9Lv8I1CzgdIRqqQq
H1qsmSxzcSIAS847/nlaRIZS9SOJaRNYjlpsTVs0pDDpwsFsSJi5x6Y1lh1H7ZE4Tq7+OyHalwzs
7ibeqOjo1Wh2d0Hl+BO9GE397PWn5kNcadCiUX0fOXHH6ZSyZwgiH9J+1Zhn0q/z/cLTU1AN8Esj
ZBf9mWOwq4K3WwOOOiKfeJxxdpTzv6yrb45Gvef1e6Z3TaLKFMVdmJ0uFPZBEYlUL5Fcs2FFtSPR
Rjo+z2mydIUoNmIY7+A4xNscoTApXyNwZzlt/2M0YldqSpjJEW1gayzsttzkFvpbI4dhpv7moKxR
+eJL70OT4NsEzj1yvc+XT53c4xWUMaU9GBlD7IY53/ZmM+boRRvnWMvjk0whnb1mR8KC0h8ogb9E
DL0/1uDUIYX6e93Q9jACUhjhWL7VGl/TETmNPKumEJhNKnGJi73PDjI8J1EJCfvGig7aNOW9Tuyc
vzid5thtEyXWirv2CRAHSiHAoBT4E4oVuuM2FpAwyZHX6DyxhnoRNeJuLSsYVp5e0FpwAPxHC0CV
kDK8PwKkCaDBwzF/IgiXouGhWVeuabrz2lTJ8V5FsSLBpzLhs2/sXTr63Hp3YXqAbYepes86NMcF
8XmTS3gTwl+6sDbOdDNZVGXlmERZkJwlnEfmdyJEP8ykG05h75u2q5/dj5sh1bs3/mjZ97W2Xmmq
SVYhTI9z0Ckvn0LixxI83FCMXp7SuhYA6Vb/OqrERjruEq/L+PHBkqXgs6pi34mJVJ8zelyS0zCt
e1qI+WXiSCpnqUrDjjnlmHRya7WvSXsQcM848+jhwKpM35x8TlBJgDr/vJGLneOTjMgRFaMjjjhy
j/SAnVKluyR9aKB0TqcyEBNIn7QydiQLd3kTciTNiSVz5BXe45GBOlsMfxskcfyhqGNGt2P/RCyS
AtLWhnFnGrbyPB27pEiOrAdidpmFySE6Yjm+DitwdTdefHAKVFFW5m58U0wReGypZnbsaMid26w9
mkopW8SByPxE6GAonW0AQh/6UZc7CDPEjAJWthfSoWEQSZHVeoYrTg8bulzqXEVcbVFcIdOTvP9x
DWaFWvV8LbME5fzpkwCzoJrd2uBwrQG5BqlREfUFp/wccELTk/wjjupNjMGwk3b7mG/jh0Y5aMDH
+SdKtO4pqHSxrUFDNylIPGKMFEZGpoPoFWbTV6LwgFKLgvlb9J7dYh2sDOmAFjCVAynOOR233Dgy
KnlDlqPYEEYgILwHAD1wMaQMYtnCRa3ObUe8iekWfIdwnJZAZhD3YlF8w/12BHRQqUAlY9/YD3dn
c4reTzYmVvl+n00et0z5ws85PcegtrnhusCCSdOnwaFDC/PpQQ3Pj8aCjGGaOeM2dtCxk41jAVMu
pXoBsxe2xuSB+RCEbI/Z2S4ImUCP4scY+draPNGEOljY/5JhV2ueQtdABI3mor9wMLTSpyimAnL+
e4jS9/HxiW5OYAzTtBcf2ZyEgQZUCimdqgQNzen1u6fTKBj8GQMghP/gcbLP8B82Zxc5BafPcxs+
vj+EFEkqtFXXySNI16jREQgEA9Hlq7AJAh1YNDY4m4tEYAO1HK2aLxzcXYRda9y+whhJmTE1Aqxn
NwDL1eT4pjipfR+mvfl8Au3e4QIi5WVnWZsrj19qTVbrfn6+aCNlStZAwghfNGzcLzzsGOS0oUBt
SaWp2pbf+er5onTYLZCa+nGw6ayCHY94lqMY/3y3aoSjB/+EEyJfVlIhHfg2rnm1myYSGjSHM8w+
CKV+dvHheiVkBAcTWdaiQwzcgF0xHZWn1yGFvG1+9xuwWTdAUVROxjU2MMfdF4O2Mb6/eWrPo85K
44qsLv4IcvN1ZpwejvAtMwo5ty3aEaIqtVeEPBkDaHl1gUxEDKdU3yTXY6UP9wg/kXivK6HJqdCl
Nf2BECpN8HpizDDFP5lQATDiNLjThtXUE1uOHWYGCk5tKpDU91ATV5mlRjGE5scBTHIy9yhFntrd
lGoKvPXC+DjcKJ08mXIjGZO8Hm+HfSR9MpvLj3iIL+axL4ajy/BRhbHStPae4JL2g7xGE9yJDVxk
YEuM/RUaWEERsQLIozYz/CQiK9JNKeC2xF+swxd577JSP9Jg17oAcTy2jZ7NE4Y1z/yF2Lhv7jy+
Ehfo1pRrIkGGrwZiq6YADmfSYTelIrmR80Kd6MmZBetCKeUBL89sXEJSsehEVehH8pe7A/j2WJCe
HWEHlDjZx2eLSZI0OjZGZLYz9pJHU8qlUpJ/vlKTcIzB4kg2H/cZQSaMaRnAflVQODVXbvDFYCI8
gVHqk2FLKufQySrS0R6UfpU742OM3eAmo4Bck1fd6dpB5nO5Uyrns1P8e4TCKSRjbTRZ6/G+aK8u
bxlAnbSElWzdliP90X8HaUHxYzodRK4BFcBAACZihZWTnAOP1h6OsBbZKlfdtFHMW+X/fF1f3eLV
ykDq+tnBg8T/egwuG9biUlZn3EnFhpnGN3OXy27b2TNhDs10xDrSkJOLvRW72m7Kp+30k2CfRTLB
GSwPIqodW1hUDfaWqQpPNI7OiQ+uZ6bBsaYyWbPapsjFjzldaMP0v9u6luPVRSCEVEzQnxSzG4aD
jzhSVrDAj0Nd7tvXMGnTQEcUC6ppeKu0C//UPJb44A3xnnaJuj2L8qYGBNHpB6kZRVk4AtVQS9kH
9NO7NSofFXfQCuZN6k3VJmTMRqxvQDdom3km8wV9eeCPG5PCLTW89dekqtraWMvnZhkL+8lYt0/O
Cd6RVsiD+vMjANHBB+L5hosMoaNfw+/H8Z5yAjrXvy3Dhloi/MjFSkX5ySXceXF+dSI/MPkiY+v8
Gpfs9JVunwS78oSZY7i077msAo9lHjgA77eUL+rXGbsnhlV53crfZ/oPI/wwTrS/n80gGoWXPd1c
hY+P9SRsw21EFjiLBY/ApNmtm250eEvGl2vzolhjKiBLD1WO8mtksQ24VICf5lAo+rNP+9oErYf+
GGRmTdcFQUq+GrX+XMLPHgLjwjvNtDamZtD5lUyiJ7+5xmgCIJSofPcFbgI/R0qiZDWFhX/tUPWO
SS8ZejLqttN6TPjPa3QmZweQj2S7b4CevckS84QWaA0WlC5c2MCSX4DYnzpi01xVIjJ8jqN2v8Ue
neg20NpDx4MxwU9580Kwwwh+ouAv7U2LzOze8ita+aBeVovz9HU7XzvD/tuh+G4vDvL5UqwSGWfG
cNhn6v8EuxyEmkZkZWxT7s4xDV1vGRFCOQBwhA60w0QAT8sESfjxnlMM+oSCfuMU4EV8IQK9emD3
UKziLKZ6CdKarUYkSwOGwvoETdFGy++qDoaXgYm9ofB+wlP+ekXyWEBMqX3ScJS7tu4dCkPmtn0z
4uWEQHlOPu4BN7beq8HOg/MAo/cpPKLqL4y6d5BawKiq/H/o1DcfvM4pvOdtPktgdBwFg5RfikrF
eioA2AKHPH11iE1QJwAsHNcZLtzs2b+/jXmgOh/38K3rNkiNfQ8u5O6qyMghVPiA47rIs3mqyeis
Qh6vj0dsc/+9Nph/HNIweu6SagSxOyHqgOO0v38Kix97rdBdhdmOrgrojGM4osqs+6RybE8OwDTU
FbuZf68c/KnwmBHvebHJXgmFsKcunTrwBki0V/okYal1vo7uwgAw2JxZA8SI3Q0B1JnmZG3Dhz5n
iK8LUnJBuMbOnwS4o5PJrsWNgDHWw2omkaniWpGwF/O2gLrtJhlKdw2VrIq3GMcguY/LWaW+qpiV
zjEX08P/fiHfCjbhfWuNdomJiESOywZKm8zUbtNkGb/2TUKXcucu2jfHECNfbzC0lniGbFkrDVX6
pMKggOeOWSojYQEYCIrGdxC6NuPtpruq1yI03lhwuiWvGDPC/YX6JbNb5Vx9ftJmN93ljD/xmVQ0
HY8MYJpOkTUH70BXk46cWzKPbHK0pspJ8indrNVS3ApHX/Lak0NgrIsveqaZE/EEgUgrAxsRYGbR
aGCLRjBoXe7HU0BkUSiiklR+l6yTNgNnVHqkuanwic6UF5VDZ9UJMBA5JTcNVoCYfJNF02suoLZQ
HIbxU2CVIDC2cx7ooZemtoaxLeu6x1vW+/YUJx9nCZpy+sYWn5neHI2PwY6ONrqwhqlhMuS4xMpD
8bcnCXiAixUt+vEHQIPX6zkl0HDyW7YlKcZ6QEMcnMPAl5uZ7Yp03Y7w6UJL5O66CppMpH43v0Uc
rdTPGDGhOmJOQpbgAKDp0FeFpM+z7YySbw68VrUxPapEK6FcgxD//QaDzpqMKf9mFWKuenPwE0Am
JvuoOnmvg917/atuq7gcN5kJQPEsnr97bxzx8iEvgov0uWmIiI+RMNYVWnpWMkYz+hzZE7b5s4PA
acg07QPLRzlRXp2L8VwnryEBi2nKqFon73qPgqb6RD6MYzlgM8pM0PeDB8H4soj1hkOBJ4vPvrd4
LM1FoW1+uqfaTAAE9oqLzYCy3iXzPzD4CgUpmTuZId+pc6lmBC3mFDKANIgtlMqqHNO8cT0oDU+A
Hg99GH56LZ25TL9BCW0RADaCKYp3AflVTqRFD4sh7nmSDhYl2xONh7zckA8PSJgJTF3bgukk0vlZ
shcAjaOaK59JoADfqYAL5IgXfA6gvX9X8KmUhaJltOFUUfWCJNdLCsUYAIyub3BsjOPWj6Iso7+1
b0/MxjH1MVnjL6dUqCrJIy2kTgO5RYtCphVxiIO7fjmtK0IS3Dx4ezpEa3LzVlyF2WpczzO9hbtR
2aYLaiV5FJ5qKRAfgHk6XqNSHyxq+whJ2f5U6zSdsu5A4O+A/oAojYh9XhpNszulY+wDzDewIDMQ
EQOOsCVojNqM8jDighDEEz2XJcXAHpyGwzNWKNyo0bd6GYrEQGDx5G3a5B6hLo0c/cCUW04gb0YX
2gi4IOfxFOgRGyf9w4BHI5WZSCniA8SqxnJFc45ublgfYQ8mZ0/NXUYNb7ReogRy7tFqyYC6MVFs
vz/czQjJ3ISziSor+ok1tY+i6B3gNRNk9WyYTAcleavkRVC3CKllWFpNipfU/w79TehcwGEyhkz8
2KE8V6wafKyM5YuynUxXg61QpJci9PzM6W0sd5KNUYqwjDFrvApI3LNfcjs5h/C5+X1m1KKQ1wpY
Xs85UD95c56LevwIwP7YtyGl3pyNJqPSHYFhqR7Y+knYzM8WFTQVeZ5THS8uIICFCA5hoDJTn3i1
IJMn+Dx+OzxxnsuKflaKx0+L4WY7Nq2qeo3D2svofEBcvNmw2JUuuePBK3MWxAYzMQt7jKUJFAOo
2+unf2GM3j1ObTB7IrOPlXRvcaz8SuTEHfvDK1HY0kPLIpNgY1Wl7izfetdm/74YgS9W5Q3FV8uP
LD9aUQ9Fu6Ksk05JbrEZ/ovBImcRDw32uizPeENnbIWz1gp4T9t++meTODJFzo97wQR+ymMcrWJ0
PwRScRFaryhu+Y0XZO+SedaxUtzzb7MvBnOtUpgYcF36zw8dkxf+MMv6DHzNcrXLOQQE0Ps/FYvh
e5vU07ew00lxsnCnzgt8YJ+rJA2n6AbvRdxUa6voAi2aDUF72XoBWthy8Kot4idFvhjvOib4MPXK
EnjNZleLVtIRMcNrbxjn2JjSlgwkvGl1dMtOIuMuv65Q67jOzCMVI2BcMcuOUz8FKfYvGaOwLZaq
Gt8gIf3pfIeytXmbNtL7q7cMinBMbW5jy2VAYJsaof/SxA0rUC7PArag5pXG7agmo9sIKcStQNTb
cNQfb2TMNl2fena+msVPUlyV/LjX7cLogViZOCyJxHVPUipaLF+hJTy/Zlc1OaUIoFspBD2tF5hU
xXjEQKFpFhsDfk2dCMaMxkT6zmyhz84sAoyR2F9M+KgtEHoRiyxN4VCKHjSZMxCDMOu3YVkHseev
6gvASPWpJUoickLByUvmcr3gZxjRE7XKJBVNgZARxcBh9B/KYVkx5YiNCvbtTQORQb7QsfWE84Ke
xXs2TRx9JMLz9kTwF9BE1p6K9AmrCj+gAOgQ+xYm1CYbehV2JX9RY5YVeSD8b/V0b/acEWcIXCGK
rhHLVGc7vJTtPzePRauDIgL8Joa1zNg3JLIjuQv65M7+dmD1qKMAKk6DyA+JHt+yexghTEoLzP7D
nVzA10zZ4ZV8tnt4b/3oQZs9Ewc+9+iBrfWC9vcXseo12IP2eTNWw8MPix+vWzNzyY5qPZtfuoOV
3LPYTx7OqmjtTlw+vjph4z440QVEANuxGSEEDspgvH5OH3ONYbAaqvC3IwGBo7zLCNf7xQfbQjco
2dhz4EtcouAWPIGAIdNzsepwjq7k+vrGHX/nqOAEZEDXc0y7FqUdHMS6v97YrhQke6Tf0qxgBOWh
btYg+9ojzATHgwXp9XZLxtjbijkfyfqnX1uYrA2caGr3YAe5jmHr5B5dotNdTHT08dJGjF6izT/H
lPWbLQzBN1vMs0KTbQFrXFh94sLzANPI+P9eQK5V5l2BhC/YjmhaFCXW4+9mQbgDeP0zg5E0Hg1C
bMgb+2kysjW8BWX+HN8U3+I31n+1q7XYhGZoJvX+PwzCvnXf4gzJdvuq4532DQBJdipYcvtI+j5t
XCT4fm7a0644cGqYHb57uUEd8/U0flNnoPrM5OXrE/dVzvbD/XmvgmjiWcVMyw7WKEoiyjM5taW1
y8R0T6X6xltPizNBVWk9nXT22q14gxjp6U/a3Rqy8tUaunfdSP4/aRKZ7cAau6fXHano1mCrsUvK
++LKdZqYxLL4w5QgHVOo+48WUhJ7mylUbHyzPz4WquawgiiEru8sMATDGhp41izLqidGpxLiUALC
NJ32z10iF8Dnu0KOcnhqSI03XnmAtzihriQso0s6Ef8CzI6vUI/B8SHQxQQZiMVLSnuYNi5YAZ7+
6eSPvufhRi979s6CVdEtBYlLh6ITptLOQVsdjdYQVM+hwQkuksitnCvysclDKfQ9W5j/TBwbvqBG
C8ze1MIU1lCUgBVqdR9bHjBdDZiJicSRp+vDM8mF0k42/FffLrX4Ech/bOkwPUvOp84y12BFisV9
1ism1mvbqgvUTDemmJQAfmy5S51fr0WZR29LodJvNleydSkfQfO8dD+NLiOT2fRQ9PqFkAvhV7w/
T0T3Z3VDw+XArsswOtUFKKYtNysKqsMq/RofgjkNjU5/3/SlBrZelU9JAJL2ttGxX+XZwtk8qHPG
MfGmVvjeLA12NcDgcfD4XJ31V7VyQzEdUKL5jKzZHwv5aTNrj6K2iv7IcmlMHITNuhcHytMsE2tq
KtHJkyDptGzS5Vc4nAzsuvEF8iZEhY4ubFa5DCpRCszv/qCB1qRvj5acnnhpbRsbgkNQBU+HQdNr
/th+zDDDwTgk+a+iphNq3+X8zB+BpNeQ89w/2rxWMwbm3LSu6dPPjYMkhjCGk1PEJHxYVIs6mcPa
zbxoRq0IlKgQclfsZIV8RIPXb0wektmer6sthiFbMs+IbBY6dLeCVdJNbwoVWsfDZCCfC24Y68EE
bELpjwYKpwvADFu2pAvqlss2dji+vsf/LSLp0L4EHjXA0EVxcOAXlQHdi7AteJi2zVjPY2a19zTF
nLpEuweAUebi1KmjTayzvhVkb9Rkh9sWx6U4PquvyTsr8MegPvzL11NiSIo8F+WnuCy4jKQlHSWj
0Rj+0vND2qBqK8xCvoGmhBolB3einWeePzl8SlG2iwpi1yhf2YYa+GXlEf7JvxtkXio+XIwyIbD7
cTFwihmOWbY+AQuxpLCv0caEG3cPri+Rb31oZztmaye+uIvX36iuF/qoNoworTpuOP/UiHN0MVEd
nSmLNWmU626dEg+l9EnZ1WiqGmBApu3GfzlxG8ev308hYghSb5D6KccDqmqoc8uD9bTx4s2hrwqW
9VGBIfX4MgGUQQvDXeA4OBdAdWH8ru4j0Smn7xEy4OyD6N+HE8l3WTt54vftqRzZZ9bOIOInOXUQ
IkU/7N9Q85duUWsc+E1AN5AcYDyYbDLsSmfHDfu4p77n6LKBpw1UZX6pYaw8RkYc7OMlABHjKkox
uDbofgwkdrgFxu02OyDNcY/3oXO4a6Yj2q3IknFO0gtQZM7+ngKc3YVu+YIcVu3C+9NRGdEUTifi
RNDq4kXaqHLO4hgStBhSDlqeRq++6Ct/3H/K6jrVum6+r6pmNrJL2gSPAOSxyFz5zIITzApg04D0
e2HRQGMl2b5P5MDuO7gfxrL0ifeHzk07rp27NZ5GtjYnQGFl2dSYDWc4UR/3qi+LFt59XFWVDtfF
OK8bi8+Rt2RdE7CHwZw0Ci0W8uPvizxkbQoobE7h+HtN9ufgW4hpYCLFEjZzxt/LF3N3uiDtl9tP
BFcTfLmQfg9nlDJ3FMNZy27HagDfyNGAnzVnuTV5IGTCJ+EaMwhRFD1pcq59xxMDSh9+HJws3ZCG
VTQ4iMVuKG0YXSHRy/IGKDtPI7uD14pisz6j3GXGtt11GGYzC0UGsWn3SCsohVJVXL+n7kmzkLGD
Bdvy+ZGj6KBQHuMCmWzzl419/oV3HOdpE7SvLml/1xa+/OCtstfKJmcY5d9WtvFKDUIPX2Phq/wl
7JmVckoIXWtaxbGLnKI0a9H4GKCqWA1WlxMeOIkWalVUyKtDZ9D5MVbcFZW4KhcYy7HFhT7lAV6Q
vU3LE189OlFzjEgnp8xwHG1GiMp5DWNOMd8kdcE68y2JespNUN6QYNsQC91h96oVD/Cv/By85g6Q
Sih0AJCob4G+hYU0A4pwPZEjFmcyLf5LH8CsSr+fr4iN6B1zq8WcBR2HizvAAzD7bPcRYxzdwPES
Z3RGdocC8+3Oxh03rn4mqXepHG6zvPDVQblfnBetI3a546obmEz4NSy8RkosSlqX4VQ0o0T/tpAk
pxf23CCyBALCowURIRp5fEd494bFp7yf1ZU4amXNImMzlL+4i54qiFG/mcssvJ2+XynWg+Y9vAwI
3E0B5HVNKB1XdWmpEVLWVxoBGWf44xagC9FH3nt2T0QyN0VMwv22nrDCZ0VbTzE60gwK9M6UAQA4
s8IGGQxJTzG9RIM7M00oM0K/e7SmO3UcfOzjDGtRVfQdpG8KG3WydTVNmzSoIICETNjvngokfu59
JSsaYHgrMMN31EZjt/WxpeMPBRvS1VUep1397oPD7FyLJrtvl5LoWA8otVeBXtqUnjgN7Gdl2YX7
1lelodL5VLE3MyXNVrPNpKw5XMCU2dI1+h/TuI4G4/dtqfCkJ0M4/yzixIPsSxFQbSYRj83fooNN
SPJ4GQyYTfIUcI8YgrnHMuhHGQRgbkUYzGqThlyOg7l4JTtpPGHy0Kz+j/cpdQ+uGFkM7vI7yDeG
ZQ2QvotHEXbWLn34Dhk7rnsKg2WVp3I44y5P8QUooAWUdHddYt4pC3PBDEAE7I/T91LMygl9LY0E
8FhukF1vUacQZmJxQl5YodDDtHjF/P0Mr7nTelSN5KUHaUdRZFtU96pVQicUHw7wJohTzLJLWa+w
kOULl2tLl/vbJJtsciudDZGEuNMja+BF/Q9fIhyEtP7QCfPNmKxXKMd08svoDTcMJOScJeYvzfhZ
YqyiN8iAORLSxns2RzGu1+IM0exDWFoMyAiAs7uh7Yxpxk/el2rw5P2j1yUcbTYxuqjpszrjUeuC
UNPg8u3LM3ejoOWZQC8cTYrwgSyXK90pF1s3cRKLyoyd24jwZ5uV+HH1KV10aXjMSl1pte2C8E2f
EJsMlWqDk8jgrG5FOPDgSsJphkypLAo8bL4sD/HSmLCfg6YITAGfjRHfZ89Cf/QINVuSDqXQA2f0
HYpV5YhLEPXJKvgZynI1qPWvtEEExzzuduIsDlS86OHjb9/lRTO+15W+nmtU2oh2hbbz/atOXueP
2kpIUnYDsD+ATX7eFWxqC0dX3c/mIBWVTHjJemW1s1F6mRdBvhCwPc8I/bS+wkE7xhlJYdujO2vy
83+Cr06TDC/I6U967D+LNhm9DHWvXzyBfmmeCvyUDWzdNxTlmnKToXsRmEmrdjhO9tDWS5atUSAT
eHtkfRGid8Z/NqzKMYxc7BWIOTDAjkdt97V/F8ti1mYbhBAnehzHD+hOVM9x4VBBm2+SgApLNZju
VYBu44qy0PrNj5KfSSzlQ78nQEYlLX1CnZbpGeQXWEFCoKYcT13bNWYIZpOs0zGYqEad9tIq8MXp
iXjvrwJ0is29s0G3f/3N6FTDD8RkzL/CzLRJLxnYNay7wg9iKM1IhgsBm9Fgfw8yx/HyTMXBEsFJ
2kn8m07Cx0SUY2v3AmnoYxCHdIOp275l14E12LOakzbq12VyByW+sdg8oQfZcsCxp9gZVo0q2GTj
sfLKG3vBj7BipQQwK5sdiFaYeBjyGPsS3iAhAFY6LuAWGAUY51wkQ7QEyBwmerN4VtgMvWqKF4Dl
t/pYKi/uNuQBwaUZ7fym8Gx6n6x2DBi3JP8Pu1JDInZ6MYQEQ7sFt3YgTuItEFkb8Osp3uPwsyV7
AXcSPLs5/8TkkvLMEaNzH6vciBCldXLNf+tbHUAbzD54oVvpDyga2EhUJtGrsL0pFrNZvrxv4RyN
NQ1dWuazrsAy/BCGzMKAjaub4TckrOSkyVDYPIzctg2PmgDZfWv19RPziQeg4mBRkD52P3CdugdB
UvpLbv2XbK92H8NuPvtu7AJS9ZkZUtZi9hYaacrUhZoibHBpiwwtl5uHKtj/yKYElTcPIZaEeayw
5Af4HZEsBCWVn9wJIhsbaGUOAKzIk7+ZUfhdDRMT250ks0JGT0bMR7kUGRFCnrua+YozDe703U3C
TqfJP7+8J2c42kRhQT/MH3PqusdNfILipQSuQ3+o774Gok+uHrMSviPgR2T98KTqpwDj16GNFbmk
MZwV1IKE3MGZ0yQfG6vUCCSv9qGv+Cf5E2yAdXWHx1mtbCMhaCYNsmL84xVdwgrVyIBcjQhaFAu/
UAOo5OHuAPCisjKg66F+TkZ99JIksNZlqfdy0f04G928wJDrRSTSLuEySf1YRcoLFs2aBJdO1o5p
bY8XIHzuhbYh96z0ClasCVSrzZp6sSiMQlDdnLpcrDw+Y1ks1ybk39WBMG1tuCPkWNzIvQsyPmW3
1c95956tQHau9dRBgCNvOueb2zhHxS8wV42hZKUKMfWKGXp8KQ97bL2yKGcKf2VP7yB3YXq9f3W1
p75BK3euh4AE5QvA1WGacHT+y2RdcHGy1QqfFbw03EyL3MLQzy5U9JFuijN+jPPJ+umnF7EHW37/
afE8cjKGCsE8ovKwNVAXshidK9cGI+IdabXJXA2qAlpqX718dAdwUNviJk3+5hZJuW9gPjqr7hBs
wfi10pj3xqiyyIncNABZPpNi9OYJcllHkKZ/HY9m/9DNh7cxcD7oc4h+j5Vi1wpjWjYOKJgn2Phr
K1VoPEHI390ppYlvbJe/6czaBxhd+jvCWqFZkuewIGsj0fippgcMSsFFJ/5xwEQwWKdpbz0tG9BJ
HUhNGkgsdlLC98PPuDecA1/PVarifNsA8WfdT8kVKm6JN4mqsNtkzezAI+sCRKF7s6/M8/HJD3IG
xxgB4CoFIXvTvR6X4agjr9TNd0lE0GGorJPH1HRQQKHlRgfF/dPwAdrOY75mnRx2Yc0ghbi49KN0
1GwUoQgzNKqTGku3G6UXjnqp0IaIXv3L+zdLTC+NkjYsE8RDh3fGe0a56OpYL/IosdCsW+BPbcif
hcjsZBI3sw31n5kJimbiHZHMvXvyGgYYL+H6HK99vBLHnRrwZ0tLRvmehlp0TiwfQCVwzgFtQM+x
B/ArkULT9hPtLP9YN353oBIg3eDcRuFE9OocakBh11coN2prpPpt1NlnIyRsLyhUioNRfEOHRBaA
QXx7MBXiC2rMhDLqXnkWi32ZWiPkAXi2dcWSChGk8WY3CnCpvOg8mgcul5cPImRBMXK3UPhASTyN
Jd2elZhxSw+MjVJ0uFZBVwWwOfIgZeV19jTIcKgsfwSuNxO7uFvcx85KR/sveGnY6QK3G/rwrzaY
oxz2vXcmrWco5OX3s2W91YmfD0uo8JgAG4iAXS9A+RWFQTmOPHEfXnV4i/kRq0OAWPTCG7IWTYb9
26lTgcJic0ljt0tlyT1s2nnUx5WXrkTM17bEyhNyF4ZXptX8t8pdBsZa0bYjayKImtL8SOp/bEeW
9QTr58H59lwnTLCol4koPh8RnwhMPlcITSDR/JHFBZgbESDWHFieBhu4nNAa9jkAx4uKSLNQRxMn
uLVIXROVkdtzNlwA052qqXafVXHpwhWMr5rUjuGb7ixF2PVRp6glLcSmEe2RXfPjY9tKHwbrgq51
w4+/Y91ZUL6FcoZC6d/oEnER1RoSnsS0BSeEiCfcSRDqpAA4AcK++1DSLZ59QmjklbBCZx1W0tua
lf1YLrnw8Q6AQIvBX9rt7weLzQOb/PFA+pzEU0tdWPLw/xh3Ahlr46aVazEJAeDW/fAaogiN61wV
rkqcVLQduv1mQX5DIJwJHn6aHCPe5mzC6gxZPucDEFY0GMGZnOcE6sTMFk/f0f1vAoZppaMwpcxo
+R2bQUKNAODjTvZ46Vtjh/AIj+ulhz9P6xZU7rqoyel98bYanDU2Ybz0ww+dBmk1ke3CDXEW073f
lHFWdD8mHnJVNJaqxWpukZoctQ628lVYPJOLUr1bwOb5cW/iVibxKwmpXc+rtZ32gv1NM5+iFwhH
hmF6sI04x2ya5YrT/ijJuXAx/Yj2ph9rPICnHO3zJj2QIwf1Y+Aj1VDdp5sg0P+ky/r2gm27ZVkg
XE3XsnWJD/wov0vk1jIMnqwATWZTsfAkGKC/grM7WleHOQDh3ixUmNALWcXBWJO5U6ll54Y26Ep3
cGgnjRAr57RhPMgzHO7jKBKBdyQGSAHYIfRoDxFK9X/VAcM56Ek86v79vL0S1sP1yqPpV0WHK5cc
ge5NydhvwUdQbVZeLtpiXvaLrkVC1u0OY+eh/D9iWwteVmrfT4L70gXGEHW2Rq8vmN9l4yqXZ58L
Y/KwPFFC/SBVj3QgOy3TSOdya+5oPbMA8evOTD9JKZTnWWb+A465U/0ZU8jFV1FhCZWOSGRQFlZd
EUYg2FwruDgUXZXXENl3CPz9c1qhgY+UiIJNQzcbACK1BmN3Z29PMaVLE5XOyTxEY29BP1LgA8Ko
MV2xehsDSORDFzGyWdldscJ/zWOjTAXDXLZ70k7tleorvuxMzs2NADraPL2QNbPKAL9VqgSpJT4d
XhvYPG12GD83qfOGHfMkmpEhgNidOJhG4JlLP5EtHG5NJjA9oA7/uoFE8qu5Mb5qc7lpp9JBCj4Q
Flt4YFgSjn9wFbNdagJ8+fXUGobz97nTjOWkjtqT5JcBfpTHXWte5G8Gs98I06eWZyCqXLNReUKx
qr9z2J9iLZBXB+6lP4YUA3JatUdDz6rdqXVTfe4kFPE3V8ydDuXw4vR90g86fjhc1qzgxlIzjJ7j
R5+scVdom2tabxCFKT6RFLTcwbUuTg51b0ueSeU9pMvP+GsGFAGhCmv8yjaAsGi8o3cKTkEsbbd/
nCh/+Ea3Gpi6dAH0oCmJV9dbvvV1E89K1SQTX0KrVx5EdozJJZeiZElp0leP2aYVQF0nhV5/QzAp
eqlih3UnQnGaP+bYOi3BDFu0x8IFkrHP7M544mKgHB2vYzCI4RziCQVwN0SziXgs0Fj8hOGmgWx8
8YFuvuBMuok2mu2bCM3N4ukBbX7cKRIgAwN2b2+eS28+pA28ysm+2pMKMjBabyCul63SgIIGlcJ2
TqZAlOvZuQuZJE6bztVqakkjx9bv+MJS4fQikhlIoRx7deesG7qaes27vMAli50BdjaBvlmiF2Jo
SAbKtSCVy4LiRYwZtWilGTEXDkIZnSO+Udv2cbaDZMwUNHxxf5okZJhaXMKhSzJSvtm3FaeQJ9ed
yvXVJxThRoCDk5PdcrWS2IauXl4SiZUYtXWVi4rk9K86hca06Wxzf83mf4W3UuCmJeg8MfcNNcCZ
eH4c1AVgjiIKlQ2wSJfZK0o7kqhATHt/Q6JRR1PeHGLkRc/hWkel1mfXAhDuCsNW6+JCl8dtSK8c
Di4za9St1htMZKNsGP7SnuHnmwQzE5WgKyaWp+Mg7kx3GEPWtmFYfB51TErSPWNjgLbIe+z1dE1f
Kmn9QOIGpWwcThwx5P7v8gZ+0iGsIvycmz8ql+jOTGt9S0fR63d9NtOfowTOW7rWO4Az2n4Eypto
yUFmtYbRztpHX5Jp4ag5RY4SYoYIE0GgOc1ztQm6t1ilqeNUelpgKWDJm0cj/dNChF2keWdu3O/O
cIiSJptZrywx5IvVg0/Lo6pR9RPBJ4foGRF1hvPKEfos5pvjKPg9g59sOIyF8Vo9qipSV2L1WgCl
EyJuvM1DywQ/4qaVMFRpfMe/YIlYeOMWM7dHMqthDqJQsoFdlURNfEjOloJ0SFQ73wDsVPDTGknC
FwgxGlJSXUHHmgfs3ZUog/LLXCZ6aFbtVvDFhCvKxIglhulSmR0NhTUmHDPwYhvxa4Lm65QiTcX9
5QCFqtqhPKQQPdI0dMoeY28Le1fbox64eBF1zfvwWQYX2GshKUKzhkQE6/V5s3/WaQFQgPwXoyOX
PGVf/8dBV6HzilBHtTt0ZGodsaLFllDeRd0b+G03XpLOPHyrYpWg3PSzvxTibBfuqm/IYOEtA7IY
ThQ+BvzaD9GJLwKSV/p74+hGbup8JAhCgW5wbRXwViRoPiJAJXvco8InA5zebSUNaavAWg3Ngg4W
qXCUx+/5y1+ACk6bacs7jPCtikf6MjjF+aYeUdvwoQP/RSxdAWbBnrWHbJkQnAuQxGRx1NFCiyVe
Vbcium5THSCCs4MDvWQpReTTMoATKVmKuyqtJIxxvXLhOE6FGQ0laslgXEbPwBrpx+V2gFO3Jpp7
4q7+63wJxqy8cTe6NCzjWr/KpO1i5e5+TUW+mjZ2ycBW/JywO7GyuKkjFmWv20E5ueEK6ooH9k3d
HQ3JQDHVUTOjHfF4gmvwrHugE3xwW+SrNw4GHgNT7VqxRgnZpODiCjygeXFWKqqYPbjzWV0zARZl
cUgYIQABZJnpAjJeF/4dRPJkkDlXIMmbqWhVPe5UpH1PD4R92XDcVU58n06K0ZmXwMCLpPFvgoae
XDk85kMqAgdaAvX6w4JUwWBlKIwduCs3pUUyNcBU3uj70IzZaDqWj7hOMnLNnRtu20LU65njo/YI
CGlZnaiWZrUQCGCFjQLBk3ZnWryjyuRsLKjctyPK/K3gU55ldyvBHBFsSg3M9E6O7hVhPudRsB9A
NREo/i7SoMhiOA8G4vc4umi0nhXwqqo6PMWa6Es8JyDmVQcwXTjOmwhFQyw0aKnwFumgIHLMDmby
mqc0SAggNKML9T6fIs2cno+nwjDHV3acl3lFbw8biiTeqsv2Zpn9LGh+nA4SzD4zdSjrFsmF7xWm
x0UAJI3dT7Nq1OrMBwLtjuCSjECcVIefdEXflxLJBU/zUTBhziDsssDL3577CduC0/4wumY0Qm4g
oUVpRXGe1m914DTPBkvaSktjVlja5fg97CIBYFk/QruDZfPmPlTcZNIogOGAaKz44kC4c8LYhTwm
Dq5OlU3vPi5AFqIJXOjggpKV9qpyQsxidsRPNi0VEs4kjE+22HkIEM4pd5I/x5qCeSNvcFQYk/SR
VM1zGk/ygvBAscKvmHebJ2t/VaGpfSQWtxE7FNK/mlSsm4v7OPasc8gw5pkCvCQcEI9CfLtzdn0P
xJTAi7KPWOm/hHwq32/ZByTOAHViwk55CCjeBU6YVggaTMSoTfR0xUgdjcBGXWSe37kbgB1SB4yM
ljEXV4583jyD1v6ftiIMGihuShp1PAVowCayLX71H325iYZvj/SgoIJ1AdgcR0iWmCjmZpd6og5A
4hogSyaillcHa6n40zC9V85dTv4bUH/b0I+3etL76ebBG22axadlYQVk0oM9zJZogNGB/DOVlfx+
nDDVi0dKuWg/YrPVSFs/V2ccmVU11l1rdPt3/P9/f0h+jIy/8N+P/mct0SGSF9nIvrpVB7xVaeJj
T9yG0hpOQBE7HrsRx1AZfnuG75aFbT0VESrrbKBGZ9yOSk90GpGROgdItLFRlVg9mzeX2UV7EJu/
E02uiCWavnA4dPqEuMeQqKexKkRV1nu1hQAsA/2r4WexeF6+CVkoagekzLQ22F0jix6m+wQZueQA
QpSduseDbE8JL52XUBEQChbZjzLAfcf2bOdwrQf0Ku0mbTGf/3myQdCZCzB+12zxow5wJVwaB2NH
xezbHkpfBN+uNuIDJiVfDdhM4boW4xgQsz8Zac0l/nbbRgSPS2UswdNgrYwEZYESu0LWMAuOodsC
AhUODYVZtSRLKnd7pwgP5gQwHgROB42BxCytI8y5VKpHPRe4wRRSJAhlpFlRWSDqel2LrICcnNSf
3b5c5FSp2QCfpIHqBdnjEt8jocAg1YMJAaU5R0aX/6CPa6EhNGMwFDZWjkjkxRC9wuMKWwbbdRF2
jLdy8YAROuf8aD7OhLWW0y68IlgBIlxyhTKk4vSzyGkdgTpSd/2oJagLzzIgKLx0PsVRkOGh3zSe
Gk4O2Om7XoiMnBl8BZeUhuZA13QkK6MfjYgverCPNnke3A8tpHWz+407TBkVFQIvhKx8OlVLCeWr
NUiEQzvHq2gZIA1QVM/DAM1KIhlMpmx70lDOIvkycy6A8ABjp4VSeYq6rbHxGRKMNarTeGbfg5jm
0aNbJetziElCOTVoZCJPcOJ/s+MpKsR7+aB8vKcXj0G48PnJrjZl6n5u2Mr/t+DkE4uyZnbg6D1D
Ry8tI6zMZD3IGhpG2mEFPkpP4MfFg0nd9O+fXLbKg7k+0QTN43/NUtIEcSky/Ykn/c0uKCgpeLGG
TlVDEjOjeJQba2J6eTOY4bHub+Orc80Lw7XhJOF0ya4Z1/1uS6NhODLKAB5Bj/V30++87d4e51n9
GCSyhp6Dx3IHGNhJNJD9Mpy1L/xlUBYOLkaHWYl36DESVk3K1IXMwX7mTofK2ifsf5+x8Lj3Y0kM
inWWb621D1xaAT0J6wosQkYLTHjWRaO7wFuzp/QGiFSiqejYGwvPfbyEZxaBK+cKyIrCk6Ep1uzV
VWZHmUtD90Tc2+c+x7p5d+18vE6njxWpDInR2rOO9hMBPEKALizlDEAmFk0pZlL/VL/6ZHl0599x
u1pByNYV2HD1iCbqzgdR9nj6QwypjJw1Jl6kcmsnLbwX3mHZMsT720WiCdmkbaazbnPx3kQ1dNXA
bMggL6mwMp3XXjDPzes/WHGTTDAN8qfxuOeoLgchwotdB8fEcM6Tr9NTDHeD3Tegb9Y/wjvYjGNh
smyZ7UQTA9rJSWRX9FwN1y2ELBCl5pX/CQ87xcoVMVLW/aCr2Ur0BybtSnBaZsM9lDF2teQO3VVq
FDRJUpwPzEbMzaoqJGRsyt4PZq+02r/mysWKUJllzDcuqdtyMqZhuM+h7YkeMKtkqvhTgaNFyoam
RKHZX/eEHUqUkzKcw9x9hvcpXC/I2Pr42VV64EJOAhfABEd5F1SLwcFkz5AkK40VN6fcb9nSnX35
SEoPBLbPf0nopnWfqgXDuMPYLpHnjwgFJj/ZCs4959a+tl+PlGDSlPPOL3l2pyXRvwf+751yDv4+
T9M4zXADzewaJ7PwMz6uioRVyJAccGicJrCvdtliHp/D27GXSyWewyBCQPhQO24q0oF3mMv8wI0R
UB9sZ8SYKwQmUHhZ9BDSJLNRsiQw79z/mmJusM0WSNWqFByMJTafdQcn6Z5w3ULr/v8q5DYZiOYm
9EDCZPknMwffsxGn8CFzOOl6I8csd8HxvfSOck1LO22FQFzYZbepb88pKPHsaKv3WF3Xu+6rcea4
CrVfZuJxzRuc11xJ/KV76Ly3DL8E8y96TRUg8m7gVNLdowcfU9Yajs3HqVNTLEHWEz1qg0+b18h5
rfi0f+nb+QV5s6Y1+IQ1nK189EORfL2XQBvpwVC+fJ3c6CHlMrFd+xJtrTcsjC9v6mgys59vCa8y
Xnu3Q7L2CK9mUqb/OFsOEl4g3IRmK5ViBoDYTTUn63gDj+D3jO2Q4QM2kXcb2rAVXVsNEGOap2mJ
09SMoMkYm3Kj7xK1uet+KY0MDCr21d0gcP1E74GwjvzQfpfUI/dVMoPFWqbPZYSEuKB3Cjtm4ZnT
PV+lU9MSAurmeHvpdSzbSyTycs4qZRkcmAeNp+tPSzkX1sedk/MoXvGytzLZmGnQeAYFlu8XWWBR
EIdO02vtdWIfWn2O9cO6bplURo3Nk+K6hr1skNbikSv6TN3W+IejWGTKZsUh339cIY+632rfvOCz
zKNgF7Rc8x5OjXMicChsKozLR+9aY4a2QHSt+n7RuDcS2l5w3lEbmGRNCakpV71Wut7SSQWvJkaU
cuIJHS2ozNJQs9Sm1Gdr2bdmJ95kul+pCpk22hkxrd6W1rUzkr3ODPTRIp7gzmIVW2aWbesK7dhi
22Z04G92760qIQ9h3OY1sF1L5kBXnUsw9rx1DzhvLo0+BDbaTzJZRAel7avHpZ/dIi2ON2Gv8d2z
frK3YlYCdEirvG+Z5+Zb4N/LoKCObSPApF4dvA9RtSOpefdmfWlGJxDRgH4JaIpuLvXVsxGnjf56
VPk1L2t1ay2m4jfAMZIsDOSWrhOv6NlyQYwJHxTKuMJpwyiBA34iwlTapLi7pT9haPbMTF5HFRsu
WhWFs4cxP+YX+FFd5jTrJ4Gh6X4u1zcxX1o4nDMzkReGZxQvgsjmkfWsJYNqR6iJ80/bhxzeAQKt
JEjIKPARGO6dwSFa/s+hJL0W+yeraG1qPUVpeTKU3bs5aQstBOW6HlSxwNSO7ogxZfUnoEc7Ngpv
+8ndcww5Moyy/PKV7ZRHMpfYn9nCk1LQTwXvsnAexOnHZvhDLqZMCbccfMQ9hjKJx4PTarqPDBWI
R6/YmOvPDWnGK1BV6qKt1h5oMRPQXpZ5hcHPegiAZ61BbbYSt0xIyeD9G262h5ldkv6+GwXd797S
1I+Co7zRgPC+QaRFMcfPV4vpdj9817F17TekzMSprdlHMgVmjMevsPEDeXxi6QGq83c29iPap9CV
1qbV/2eUiCHyl+ltkaqIA3e0Ivkbgz8+qoG4K2/7D1mjl0hHlZaOtqZn69L+WdOC5aSlYEdfHIJK
zhD3XKC6ca57ObZ6VSS6rmlgK1NKSpmEa4LddUwLbTJJD9/ld7xQqQYgeMf9FbiQqlnvZZCpbbGJ
MUBs81PV+IcfvS30YVVyyAknylDphAfwF/58cu5WpZym9CcqALJT3HwDkRmqJXCm79bYERfJsrla
xbPps1StMIpdpcKbtC7IsjTelVSlgLCXK8fv+AK65qYDiJARide4VkT7+Eh4ifFbtTymD3mvz89r
Tklzg9hH15TH22gIhp62G/+Oq4WehkToAk5zmfxjUtyJ7t6rEH9rfjXSJsdfUtK/uTR549tsERta
S30d3v4OQhFePjot1+8Qf8ePtuDpAaUrFREoH4zzt9BLkH9WVdaluFpg+UIwUc9EF1B1mJurhlby
szrIVWe8Ch2mTbR7uuQUfC/eYgczTwfnhnKFc1M/MKvy3YO8HfDGsPxZXksuf8f8xWeQZxpmKIsY
bQKQES78cGu49mdnWkIAzF+7CTRRoYogVI11nqOc26/IxOw9jgrmhbl7ihj3vNvDHR7w38gGg0TF
oKthJbzNnBwnJdtE0w3WuvLawxrmTWcn0X7t7pa1mrXuCVw8elQi+tRbHSaLC1c1+IQoxVhIl0+E
sHK0zJuIJjVuEbHFpt9HG0U9ansURq7do4b81SvzgaxcjTOuI6etNWrPVu8pvh3eBPLsFviq/FxD
Ob25DXD4OqQ2Y/21WJr10ai6LGkwJkX0T6AIjKNrnYahZSilD0OhV01L5Syb7n7nlAKWIqWlKjak
SyNemRSMO8ALzmpxnMLcaR0OxeQhZaQySgQFMVRZnzp7x0BTvGHTVu26kWLOpkap6v8gTr0fws8Q
CMrUa/fppx0poBiDh1nQVCLdnMmuGzm5aA1c+vtsNDT6RQdizioPZxAUkEK7VmCAQEUA8RFjN0Ze
rhiU+FzLOwHfKptQmRnNrcaFC07AYV7H7cnqOLl2kACZj9BHF7ZVw8ETH9nyAh52cObKo+Y9KZMH
3PJsAD+B48kvHUGuGA8uA9AmtiGy3KHG0tQJDE2cZCW+CnEv+sRS8nxbtfEH4T7Fjfyv+qm0aLqa
qa0+7CsGcUihQ/8M8i489JaEkMmDqq7uodumBZcy8UQC7DqQk7CTCwYGBW7yEQaS+s+xuf/DBrTP
kcpM7SiVK6f0QkHJQB5YoXYRw+KJp3W7tESFpUsUlZw/+eBfQzrWzmnkyS5vHqz+cnjSx23tpLqY
bZao1PnztDzjnfmJJH8L6gnx1do5tC/nzhGwqYdACfDg5J09SFzJdbzcucLzSfbhyTYH4LRG1IxB
rtYC/BEd+ykowvcb8YwxOy45T4gosoepalnAOEFZ+H+Or0CqNNuScQPDDQIutm8N/be1i/vtEdbS
Zh4kZYnO+3x+L0VCUNUqcjETYpZEaBYZgAJ57b0PKxO/wx748mWjbfX7XWlf/QVwRzdSSUbndOP6
rgSmc0FbARFNJZC5aRuk04vuoMXUboZFmvGNngEDbW3Ai8fz8z1NSH/lOXJ+p06tOT77duzE6EN6
XqhzYsjeUsnxrDG3gQ/uRVvllrKAzu3q4MoYuGxNJuIU9ech8F/BpUVqa5diQrA0xqtu/SqCxec2
3smmONMFfXHqi+WyFpcheh2t06ky/+cLIKRi6JV0Et+XKo4YCR2iBktmG1j1bzync4Bt2DmUKFKs
MFbKXQO/CX2EBNbSDCTZq0z0zuIqhlDvKCk7flosPrc2dwZ9KCU6tukoWtFKIODgpSauMLnzis/H
wnQ/mWPE7dTLexAYdze8tquybRgWP4CDv79oPlakPXz5FVkwP80HDXSSYa3VQbbud59SiUked9MX
P2N6gzih55/blIRynR7Shvzj2n17xTAwmNWbdhSHl9oOwzuXTr/IyS3marORLAah0Onyn11Wge6M
Hy+PJciMGi05zQi48ak6ksYYylURiQ6BTs3yRKom8iVvG6z9ZNQwy3pRrrSx9RGLek45DBhWVH+e
x1RmqQWF6w8OhBfKmFhRYVnNmLifhGlzHXrQrpAVC4yt/1BsNBYaKUcXgKfbjLg3gmBtgKRjnlYf
6BRYnFA0muHRe+EmTuKGXV3Wg7cqLGTHaeiZDmG12iLoQBAXZ8VgvZL5k/vbJP1ExZ2R5nCnEvkD
iHkSq8rlSXLWIVrcFDUExWEhQVIuWGLsDpqSbAh6V4qjUR3ve5KcNP/3zH7uULP5ypldko+GBY1r
TMcyVEQYhYkfdSJQTgTimIB6pp3q70ihBY1o5KcaAOaEF7EjnpEgfoDtNNJtXjt61fKNsNbi/nAn
CbSPb9MwqPIejMxnhVd/fCRAP1xTC7UROzJ8J/A9NpJZUVG0ITZm0zzZ6Ksk4Ppkw2o+kcVIcoHy
cxd9rr1vcbIaBgrvJB0zNPdK9sQpqKrzMQmhAiLSpsgMc72s+qZ4OpKiLb8vvvJiXF3IhSwBckAF
GXy3Nq5dPwOOIGOeevP6coAxD42/NkzzgWuJGKdM6Dhx+/Yr/dy9pZtAxI89KSxO7lrWl/f7m5L4
0vxdZXUCHpCQRVqMi8GBnHsLxuj7nQrb6CuhGmKphkDWAi/dVVFusm/ModDQq0vkJpMBTN0dLsrR
aQoW5Fc/AS4YIAjsgiiSEF+lefDSBezquZWEjSFZE8e3bDoy+PnCNtmovQbFjriaV1MvJv4bJB1e
9W4h29XYr0n7T3tNb3BngsnR1GsPJILGKe8LtQU4Td77o5PpFcJwWO0imq8STnRDUQdhvTfXB2CX
xpabarqayVZCosAZ2cwE6sfr5SdFv7waUQKdU/I6H8T6p0ylfPeA3//HUCw+ppPpymz3FI127B/O
jnl/66QRxlQbKObUV5bH+nRdrBk+MvFlfDULnX4TwWmeSvi/nR2fyzh/FJ1xz6hkug5VsdS2ZBBP
FyMnDAtDij3PccyLnDeJSMcTbmqhQThE71lUARamvZnazxtnSsnEG68pGxf8ZOKTynkeQdl0NGVh
BJGvW1oYR2yms3X2NuBIRX9mwN64ggqRvhBqh+jdxsC76+6FV56RcQZAynA/G0c9uolMjjghzw4C
mElA3ZV1AZRnakVBvEPNILdAxkC797T7M8LYBmkI8L6N1hsMAxgCfBNLk8enI5vPpH6PWM70bRa2
aNXTJvZjrGn1cD49TDCcyquPNxXtFu0uBzglTpCtkTO17cOTmJnklG1IPS70XVoqJeUKjv9oB7om
8AjW/SNlIWqSt/C2qLv/Fyc829G/vj22RQm6z1TFjx9d7Fyxs35mkt3Jh4IwwkyRBqmoxD4A7syP
hvvPRsynPi95WyDM3tQ2FCW45CaiY7uc1lBNdKAJ6sv2o8Kq4yQASgZ2gqkm9Pyv+aHmknYy25Wz
CQ1gEbhqxvvZ4O0soS9RsEilb8mrcObQMFXqyDh+eRPTo9O4t96MEqoBzkmQHBiBZYkS/4tpww4n
nRnOkQdJF3D+uPI6HD8pSO5EJ60GAp3JWB8Mx4C9mQTSKCWtCwdNyqXo1BQPvGPzV3pmuFWgWgKo
uDe21C8JCs8oLrOIOaF1gcijyPkMLHh5Awg4Yw44HhWp+NBkaeEWCKcpSIPT7+axPBY8c/k5ynn/
EjYwz82mIFTtBgEoKy1jgNz2eNka0z8MTZrzwmOR4U6hwds5ADHMf4YZbqYa9qyeNglL6uEON6NA
mM+Sg5N62v5BQrv3FzuOTdst3Cy/ip0z9dWhKrztGVN01PXS3P9qoXkSkDeU0+ahcwWQkji2/QMZ
D3mCG3RBMSq+8FDWui8zBu974ArreANGOHrbMSLM84GXx9v21EI+RBQMUg265XjRA1JdpcB2Ab6N
mfEBQoSgOuPRJW3D0QdIKHWc8kuqqzw6Xa/K52XTM2XnBP3cx226a00H0/ubPD1j5uOADE6tcakT
wZFmaxFyvrqWZ5knJx5BRfxYRyw2G3UfH7UE0ExLzyRCKn2AoWBOtbS/f8vMu+B4LbRbJJt/N/Nb
WVGRE5KMS/3+RZTUfjHelHIJhv68mcQxYXYrYr38ceCZriRWTEXfmuuutfWmya9F9OwgVjoIh3PX
DZtI2tUj5ZScM4PJunOFoO2drkx2O18EhfVGJcr7jneWepghlDFNo+5++kBaonx5Hk5RyS+HNgp/
+1S3NfhNPhp8wNDhXFPxiSZN9GYLMLO5L6AONdOYxJuXvAGDM0Ap38nYx9/NXM6nscOTHKie0PsT
PfyJqDIkfbY5rG48EYhNqbjouGheYQx32qSaJNpdZDdhAWhkP3l458Qg4pL+JJDcNPiehZacb5cd
6askKmk84BXUzI2qqS+93JDExPckYxj0JI7S8Ksm7TWMKiVJIVxvRmAS3zTPaBJP5MfUVZnlTsYx
40HrMRqMFAGgleiew2PQIMl8elI+kYkOF+8dziFaop3aZIMlXxsAhg5LRgQInlAroTxskn9kPw9b
NqQ2BJ9LcZ9VMkH9eGfYooRQbx6IWvPgJqRaXV9seXACQLWhZiHit64yMyz8GRR+ytiVv0rIDtqa
A1MqOzpORzr4wPrOWVWJLZXp3RFoHpY5ETklAFYXnwDifEf/DOo06VTTDpPT3TZOsf2F2ioKFBF/
6BTySK+rLktqiovlf6wNaZZzPzl4Y/a42m3POXKKSOevOakgKhM9VoMbdfNiJhbZabpr7+OrQD9T
ZLCSTq8RAX6CT8nyPoF9/6/AzbGGOkTycf/vr6CUZ+PCklKLWJsNH4RkW+O00UZkAZCNGp2UePHF
tDl2Nfb4+MgxZiv8XizNCeE2iSaQad1YZi2i6Gro2HhtoT3q1+pJNmoPQAdvEjkff2ilRAcD5XcW
mwAurqxWN3Fr7Ra4DqKRK9q8/rOMu2f978ySCnJnylMImY/Ay8KIJA1SBKNoMcqQcrAM9puASSM9
LrzrhmuEXsOA2QI8SZiuJL50CJRue+TqJfC0MC+gSyPjiO7+LhjdA0MoTJrGTlzXwhiPyJZabC+P
D6/eBKbjqhxU1jld/uURjOiQZUEJDu7U/YG/8mPXBOoy1sGuGOfvdja9lXcs72sGX/APVovCE6v8
T8YtTZ6mxXP0Dpg/srMVBMRM6VXCLa4avmL3gipqxigYPA55JaK7S+yAYN/B6wrdfy6FlR+yp31c
9YfYc9aWgtXcq/4h7xX6W5uAycKKLG4Yr9p7hArqxEy41sAwA79WkHei/oh8fBLPvTLGI7hhcete
o+RZzNQIgcOUzEhSoWL8M21pADmC1TsNhIyAHqGDIqf9oi/TJJtQY4i3pyrP+0hm1eHAAMq57QM/
rWGpcarS/1+SXQ9+mGVPF5azut5LzHI1TLkBqn5daeAtAGWXt3+my7X8zj0PhTG3dgO98wj0D/+9
HmrEprsUr8x4XG1QJLbM/gIHIinkKSl7udikVsf0ViuW+T0AIvpPMAhatD4S6kjOEiApApRuBlnT
QnToTssDRfl75Exd+/HnZqCqsyXRj2YBimb0Xix9UmgWGQTQve2Rzi7dm6H90abgDmk79sATXWBs
/m3Xx17HjZYV26XfDtznARIzaGgt12FvKu/CXRxOq0NIB/6xuRI1bGbEMqxU5KRAoFJCgqjGHTAN
boXQGOQ6W9vI/RlA7dgicJZGbv6S6duAwHxw+vwKZ5EiOuIpmNrmweIKeO+JjSIe3oxy8/n6i0WS
zt/mMcbND4U6ftYIYPo8PpRQGMbVLmBm7yoIMZ/a05ltxU5BIj2YFd6iXyvwkm9Ls3bBzYCOTOZz
XhUdgaxn6LTrwtEcik2zvn03HyQq8Y+nvP3yH3ur+gHEZMMkuVd4RqQQJmg+D0lQ4yEbhcaCT/qV
YPRpW8m5QyweNWsTr15L1n6DRti0xQylbuGSBJaZt4EBCUzFuOjnPaptp4uPxD7ayv4vrMdGBYbs
zOFbxKnUuMC2bMbuCGCeBOYi2JuxI81Uxbarqh6XbqGZ02aHj6+iBXoJinHUnepBzjGzt0VmgAl4
ZN4DAoiZU9wMLNr7i0bymJ/wVT9r3XC0ypZpaEgFuz4QhXY4AVw0jqjmi1/I9H3BbNvDG35aUs2u
hRMb0+LB1NgXXDuS2sPI9A5nEA+sKZ3STPu/qPBVxC9BwWxuz9Y0oHaUjKJTImrchYN9/TIfVLCK
BocJQnSllfJYnnbxS01bCW9L2R0d67e6YGzKqk2Ybj9j7Op3jWUlQNjIvUOug9P7aP5FQiprlj97
6VX/o2watNKlhnbWmN0Bgf8l7rw4feEnSv1Q7zCfn91FiuVWya7bIf088q//PswzeLkYDMYicXL9
ZYzNPVzfZ5lnUf0mxQ/sCZZqaQJY8AZWKaQgQ/lRnS3XZieazIjLtDpZC6tmmV9RUQ7KUTST+Rur
NBL0wlvlky6S0en2gPy/II/sSbaref1GKViSycT3j5UoYZGu1khmb0ULQjlfbB4dLkjPATIXeHEe
J7m51VCJMRSkGsJE40noamP+/NwWlosRLJzGXlB3mmmgXwsIs2UafmtwKzY3AyOe
`pragma protect end_protected

// 
