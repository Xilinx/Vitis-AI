`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0INbis6m4LNo5fuoc/7VtaFb6U
0+5fXdMnwe75smPOBFJPEC7G1jJjzTejAYkTl7IUTkgZKL+qPo9QsJV8bWnGHQsxi3gvlQOIaFQc
GeHAIu5kCH4qdG/Rd7Opht+51SV6MCUG+Jzw6T7NCWSvcK1kUSxl+7AIlS+WIYISlJ+EKHtGVS9i
EwJnDml+BfWpTB9xPafHkbwEu3i47lW0rm65AtBA0FQc0g9XjSdqF0izkDx71iLWtwdJ/ACCBQzi
xKAn3O9YWWSM42rUdp7lLnrMrZ9dqlTFLVcDnLb8j2EY862H3wHpOw8iHHqf5xFtZOY8QzpAi8f1
+I34YYGY0m4YOx1cYvkBUwVJemoDRq8p/rkCraDm2HAi3qDHA4rQWnWy1GKi6QMYLW48OO0SUwfm
/Q28Hm6OOnOyBhkPWFCJGNwnXo22Ui6tiO4YKQTmnGJQCP0X0u+Vv84YEzVlre4RdSP96pa90YHV
9DTFcOJ39i9bdmqFxDbMl/PRswwSH6aQ4BluilTlH+2PY/yaDFqL1btxGgwVtm1Isu+Wd6sDjnKb
ntTpmBB81ImfrVaim4josGQ95UtAeU2p1/QdAfIGnpMH1o4ULaIyX1nQZVa8R0OosP9y0KZjaIbl
W5HVkJ3NCG3sgzSUmds5EOUtWLeiZDSqZngpsf8owBjraLlwkS0/wR8H/ahM4p9MmqR+fxPELZiD
7FNBbMku6Te7oVrmuS8L5zl0jeKeLrJnIqgxoDw6ARAocqmXm1KbGgcFW3gEKqRKOP/3L56vbE1/
10QjyQDaiDVqIEFOr79SL9teItqKOve3D6gHbcg6U7CE8oy+IvhYscuW9cYyx2zMHidIyHugbVbC
DZrRBgIIB7RceGw9CsY+Yn14jGCRADcR3pdfb4LEP1OUYjdkBqfxWFiYa0LQR5C1O6uSbx8lMFvZ
cefFgnMcelLIPJzg2OkSzAYkvRC55/poOZbEd0MZfecqWmNatl1Ghjq0cX5t33r1YOBV5ksN8Lnz
ky3brZA7rz/3kTcamZrCb6mPQ65hTyb4xkMnhKBLNCkPZPgswddnYz2ZOpqIPuNgNZpmqKn0jVIy
3Mq5JKy3J7FdJylRCKdreMJcpDltEu1Y/qWvVBLHByCn81xVPzIc/opCQAjJyCJyD7cHXJNBYVLw
SGkGM/p3Za/M+BFxdM6eJSLzOmdz3RPToDWfXwEUpw/YYU5J7YcqvsQ19e09oAIdMhgqTqYTq+kF
w4OhefIuLBA7aYBmaFniW/tbjkVRpYsivR4ARVmYJt8/Ic7VQvP6V5QF35QVCLRmjImfvQriwmCK
iF72q5snos7yVUpYIB2/o05Ke2lBywg9z2pljrBtWGWtvLDIE18AhHw78y1dr6oqHdqTV9DwED7w
4pYgoM+nJiJFZYsgZi66aRFu+PQYiQxvw1Ckqk3kKN9CEIWR6C5QTYqQDgCmEk+LcWOy7SYl0+8T
mDQv9/JrZ4B7WN8PmtQl2FlgioAXsHVhB2M6BMSZCdQjBqCq+e1Mwd+YZqdbMN0IYWsJrVQ+P90v
q4T+XJxzErTvHiFzR1eikS6cEo1qisXZq0I48phGrw9GJyimRwpvTAZ8KhFQqrZYE1wv5y6kzXRy
8nBlhB3aE+txJ8rFbDd7iRTLEL9ASMJ4BU6X0Ko7fy8LDfyvkdjFB821Z8Ha6fh8H9u6QknNVwGr
0Rq1UGGOyJKEgcy/3EKiaW00Hp6nH4xiv+Vt5kXlS3mZigCxnTpNsJQjfmrkOVzh4owwhIsQHvxt
i0+RtFRZRdreIswgsdBlXWvN9TqnMmSzQueOS82DZmiU3rBrWo5hpJakC9TVlz+P2057MkZzLIjA
bjWMR1JZ4gF9jbyNaZSaSAyAg/vAYWDJKXABRAVB8zAOQATOVSC7Npv+Kte8m8j75EcDwLfyrIrk
fuIEJ/M3MeHGEwlM2KSEyS0ZaLBS93sk8elEz8+a5/s74PMi6nNGJJ0x7zYSlTe/a6hPxC6ERMAE
5NdWywehPjJM27LzOfdJailVdKuasPDBx2fhByIjaJ+3+mhoZspXiE5NlBZKrI7snrzquLoF0JmJ
6/+FDCPYwVki3lbHl+uHMxpY/jpIzpR9ep722Bx2tVYl+T3clhunYU1WNio3fdrMHzhHbW3lTDYc
Tcpgcxo3/VjYir6VBUVTokNK57iqQDwyNfZEH/tXxLAKveij0rPR+Lynxn4mG7g8eR1OoW3YTeiS
Inbm999fgzNYxGVC9xFfGBUQLPG4UXHFtKUP+9B8E7FAVi4hENUBkGZKgQHx0wIMNpI1UryH9Sf4
OUyNyjfp1rHqDlCbAVUrgBsvMwdY+cH8r4+G/PZpGGz0nCFagkSBwfQUcyVhkYbJUFoTfuhIua01
TwtX+8CLp/bUxZ2nmRAVtiIzIcs3qjG/YUvMh9EDQleB0/rMTC1t7WCEGhfoeYA4HMkVLHnl+gil
vN+8n7bxPlKOjQGXCxiwXm+C+L136QstYltVfM+v8fWw3Xx4iMsNmgdbHas9pd9yFNcUdyQYm1pO
madzPxhqKSnQ/LTGleeaItrGjVEgFbHiTUxRhYN2B8CC12Zz/4CvVgHQ5jd7c+fKVXfS3P7lxLFY
zSdzEU984EWeDM2KUY6F2Nt9Kz4R+nRb7BSJgLCYe0QXejQxvTpc9sQ0ZAoJHAs4o6kMX/bRtgz0
BAwNQNJi2mWly4L7WncShMPxFtD0EiiTLbytdytDH9wHHRxEHQTeKvVDT+XAsR+C3T8RMJnFwQ5d
rH6UCvOtF/ulstWpW6aBAtiOqQcWVPttPPUxAg1702+UmqV2nHq67ggV4Gv2Z4aQh7OCM9OgOPzL
drY+MCEz/aPgGu8PhCy+kSg9GqEaYrXADB9ssHX2G9zxwvlhziJz8FFEPheVBlZDH95vmEe3T+TC
xYSjL7tyxPfrsa2y8oYk5E82jqONt+CRfG3MVy0fYHtewQVdG++gxGuxjOJIrb/rq2s2HG2NTz4B
921qnQ6nKi12r3NqGdnHQEZGybcxwjDqf00NouuOeIqve9UM/VH+v2NlvIo734XLAzaut2N8aq7x
JHbH93kPheygX/X7TvAbHPrPV19ZmbfgqKZZ9VW24qKDZqmiMiRuy7+V+XzIguQMfumtb2SMT/57
k8sAgbtCJJ6kof872wctQOOZ2nzM3fJi5Y//nsg4RYk6msjwf8JRMW0eq9K1mJHIUGmLwlAkhSGe
X3Ft+UkqS6LXQ/4OTHArQTc35mhafRXo2EbeuNusTKckuKu0QtP4xPoiq9N3s97PMh3RMLqCH5ZE
KqmE4epizD6ihiu9Fi/G9lUWN+g2O5jPLpsEnNyG1BB+VmtIdRaqbQDtTuJA5+4Tr8CqYm1hZhgu
lX4/WCXWq1VQhHDSm/x11PkPjWH/IKx1w0YxV8PnWjZrhMjjRUctmPp1TB8j7/sH/RcRQc3ICSPL
09TVyYng+5Vd7Vc+hXNSP+p70NgXzL6fJFQXXTCEp8GSMcEIJ4bB8wgsLl+UABJsUcVE326X4ZXr
56AXuWklARtO9krrZ66/hEBqT32xLubwPLQsYM4Isb1c6U1534vXU+878wqRtA1WTjDy2oUjOHPp
Ey4GYQdzW5NGqOCTraFoXnzn6xWEa6pAdqW+HigUlsm+oyDFPs7DdjY4LHiRnE4Jv0NeUkv9eZoL
69Nsg4sxmbA6DGDf2ylB+i8zOmH8nyO8tb1zFq+BsP0eYgz/R9vtTgATHFxoUxVWEZ1a1aI8nr7e
xDEDdsc6yziPTV79rUpa4IPLbia/cFLQTF0T7qaC0Bq/pFD10R8GBDgM1lLeHm0My+MFaCChUIBO
d9W0KjHn2anCSYeN31lDwHwpZBBHfthqiUYNz/Tk3leEqR1EYjVKsBVGJV6BQUORM5Zg3U2IWOZg
NP8cfVI1hhLejif36b0TCovMsawo9LwQTrVCFiOwfbhPsR1tLbN5JvNwEGXA2K9XUPTn/SPC8xb3
7M4iPiY/Z/wB0iAVjnYqXas6ghQN0qlGfbNgD55ubYDhcNSDog45xT29LoQrGydqoCAeQuhJmUJz
MAJe6dDd2+ujvz1mfph5WbuGrScMcspVng5VV9oEaEwMUxkR4XOjjOJdqSIIcEWzKUKJbo5i0Rxb
B09EJUsWtYB44ktUw+Dfv6BvL0Zc0UP1xDaMIMZsUg/DmPU2+r4MmOKpkqXQP97OFxT9kGflemwt
JP28DgfcVFRbaW9rjzkYrhcSFkdvg+LiUkwGCAO0dzPLWyfxlvbfCliLdXI2DlQnP4tAucqEcjP/
apImzh7Gd9dhkWTO1WlT4vYLdb7L0dznWEDO30iYdmHyoMpdKddHSsOJOswh+U4HlG1XmDL5dGD2
o4+UdvX+P+iN2Yi/2pdS1kVmjuJW8Hu+jZQVx/FqKNPH//gNqu6NHXcB6Cgx9B5LpB1bCgkieUMb
goTpUBnB2sjEpxaWAnlbYML7KwZkeCnqLt5XLhc5TTcck1KXjNnO0PW5DLZdKljHZY8RGCQVT/Bm
w4N+hqmP8DCgRvWWPbOuOugvk8PZ+qj/eEVebuDDl62aSeeo0rHgwzOH4iKIUnVdEf7/LOdMubU0
yaAGyM7iS8hMjtZUXN2mHPR0EiUIfoLJO+K/9pno59vvbSx1QKtu+5YJhnCl3lRq4sGW3ux9+jbX
Adt29svbbiIU2CaddnA7Qy9yGQYW2Q6DtdPNPKlI6oDE/gpvkcijFk77dVPH3Yc7U0kh5Yj9jcRy
pc5qtfGTpWIIKtTUuYO7LFC79trbX4MEN5lJRreXj+xkoAPVrq17JNZ1pV/AcX8F08zjtht68rvC
eK5DsV8LXvFDuIcpr/exFGrosGtvmGhQkq9OowHde05tynMcQ94qU88xeX4t6Qm+/uSdq1LP8O42
ihmrNed0ERqjRRl2OpMCbEKXgai/HmbGjK/eFeaLW4dAzYRFNH+eEXvVCuzi6LtVHhwLyjpVh/zD
wlrFipVwjtNQ7EZ8MDenc7x6Ss2l4ZPztSXrLW4TgJ4509xVsOYjZ/ElcX42auWQfCgBRWz0YGie
tbAKs6Pyhihhwy0XXqZ+wRXcDmpAZgVpolZ/QHJvgwUS98GlYeZ+7WPICOQxHldTvfIt4PVYyuMU
VGlpwOT5Q9tSCLK6pNyrBZLTD7dQCfr8tg/bePc3AYwVn6XCDetux9Z6yvnO97BDxFrtcbhHvEal
gemPCUYvbHxeaTldo8apmt67sola0h4r8X++j2q/NTiITw+fJ+aDFIvEL44VObluYHVUwjSnhFzn
rHfueQbeQ8ebPjlOQHmfWjB4eifzPcEb4OkeO+B6DAavQiZMx9GDZ82kXf/uykEBOGXOs1cf9jZB
43RDEBEToTSGw21MPEeLgW+zvcSCkP/eMH/JX5C4gajii7sVuj7TuFd50c5zElcvcFX4OlrMNYZW
SGyoHOGTEt+d7r1GAITQ32+vUEBqGZ0G9yXF14N4mihLN6VGvLpP+vYaii5vI0Wh5qFtRGsPg1Fo
MItiLsOgR+5UCEv09FQmcDue4XFt+7UiW7wLQhSmZFj6ByEvpEn0P2U2ilwYYMeRm+UaHy4vQGRZ
nkhmgGcYOY4bmh7OWWu/txXMQy+Ga/MxQdXcgrrBmBGdloIU5UznDw2FZzwPrPLrEb7W2LKcSg4V
zOaNm/jV0DCbj7qpyaCe/mSunXl1lLbueKCqdeS/jt7PQrLtQwhTMkP2VF73SWMu1QbXec5iaZdr
AyTAZtCAUZ2f/1hrNza5RMNv3IJEr/ZkUTGOUxIzDg2cudqfIjsG9CazIz9ooUT6SF6ryXQxB3nQ
W/q1k4DwYXVrVbxsUZLoKZL/k2ztzxeW5tuFYwE7ztLVoqsy2wYx3QM7Ka7HH3tnWJftAthwdEnl
vO9P6R+9yOxDYrWHmPvjOFOiHTjGnXeFETyh8gZZVTbWcIOacGMgcIuye48mwHKDRrlJ/OrCvFKB
trL2NsQ6McXDvXrCuEjr6N4djZstkfyzUlMLHqfV7gkbA8z96ErbuQdLHYf8hCtjm1SU4aaSbcV7
3ptXsgONPArhIdZkj38Hhm0jNMokeWHSNpph3srxDAdnLQSDHt6GU5fqzYhE0XbhEpjfXO+3I2yO
JL5ykywLBMEu6737vfXIKTYUYHy/jJNCxEHaGUAhN84l+O0t4xf3vJzVLkD8y/g2PZI5+1TGxTcH
ivIa39MsSAC3soDlkNE4O9dox0HmpC5xqUa3iHtOhq/l4rAYDLNbfZ1+NEiIjLG+krnViZg2ZuzU
eNorwHst8BnmMFywdO26e4GiHyFC4A5WtWi+qgFP2HbYRWRBQIbOUC+7IbSwtw41XGazu/rXn6N6
QFd9q8d3u0Or8N5NMCSqDjsen/LbdVql6HYM8oY+u5T4Aa9nNv16R0Ajfx0zeHDgW/asp0y6HjWg
jL1cj59KMqLb9bEnQHp/5ZnxnArweWN8q7Jzx36vJEAUJSPV33jr32P5GEAiSam96F3KPS20727h
EZed67qDfACJ3nS15SG6NUFK0n+RvgUZTuGCwS8/Nv81hbIRp5Wavt/LtxY96vxt9kMnJW0X4LWu
7VZWsAswD9sWY7Q9wGg+xQjU+jZ0A3jQRlkS9VHDyQMJBIz9jKt1rqPdCXHHr59H2zFI1kj7+1Ep
Ot9AAUrFvoWKrMScHAbpMkANOPPGeacmZEn4kSCfzbBg5Psmtz3IzQY9+wHPx+/7TX9rkU18OpEp
jrnySMzebwhCBfFq+qk4LN/xfzdQue7cENUuIWmsQ4II5XFZnIY3AZKEZXMsLrjf5R8ywCCc+6mR
hk4oIJ8XXOTYk53xubSJSbtxtaQfNRmJmzGwtU3G24uob068lcy04NoVwrblPKoCAx8tJ48D5OcU
ySRqj01m5fPoNo0UHIFKvsprmcKEyaHQXUYJCvkfgjwUC6zpEBlA2ncZ3QemyhEGb9RoAins4sVp
5yQ0r8vtULjJexeGlVpfvmX0y3PAxZg9xMSD3T35balfp/9ldawC/+vqDsVeEkt3HFo/NiYR/b5J
rbc2KY7AMAclrb3u7LDWda/Ot6pC73XARXHNPH8a96+ZHAvWfLk1choc2r22uKYITH2RxFnW3Lfo
ileZsttgphplwJ199yrqftKQDkYlROj/V6+D4PK5REWrlEaoqJeQJlgVGqO0jsllU7feJosLAqsI
6rIhJu90upJPeoeFvgDt9h3Vg+b3BW9kxHU/0XaPdwKvmXRiuei696Nq2ex0LLl2qwN0vEJOVEaE
w5ZOeMQB77uKgzwOrDXQ6SzykqcM/05zPQ9W322tNh1FaLVAgczvHz7nPoiiqZO5LN0gBIB748Do
QmrG+i5pgmGF7jRVnrljSeQijaIWPPU5SUFiGbeqytu65jev9w6J8H0kAnvI5cghsetlmY/iDwsl
qJycPGbmBjfhu0xmnL+GpPw4w+i95e3NcuhawQXJVAbMd1GpHLoiT7iXPVVgkuYxKemnfYOeBxwG
9NTMJfVNUafTqLHmYFLVgJNPjRJRO4DQki0tZe9I1In3YNcrRbgTtBvQ8usKpYIm6JbUQ/Usc52Z
MGy8UpWxSQGp0pT7urkw9N7c8L7u4rmclb4jbKBkLBFP3VsMk18W8x1Vg41TjgcaRCVZtKoTYQbW
Dn5XxcVowFj88VieniK6DbJrudd7EDOCsvb5rk+97Gx0HpUTpixOwbCx8l+xUZ/GJxTTB4MNYo8E
kQzNPXpP8weuvU1ocorlGCMAPnICrI+5MhwspuBrrvFlI4yF7zemKKwB3e8mkkQD5H8Q3jVS1T3L
t1tOeN9MO9lqNJA0RRYIlHBo7YgtUFVpvsg9mdDCRywgCvlTevkPFCyIw8qxynp+v3f0U0JHXpQT
sbhR08+w5eBZmhcore+xkjCZ/SonsEw5hiiBrL6DZu1csTxv+v8ba5RoxdIc7gYplV2vpk32IIIw
fu3GnOVBZZFAoMwBIyLGREnBUiAIiceu2hMcH2Qq0sgKUpnIZ5pJKMIftqoqzNVVQFikU9WqoRnX
vc4azdpTqbbsvSpHI8f9Pu7hCdVFuHbrH+IN04+x5Qex/3j1zNDbR4ci04/qRClqxiwVFZF07yMq
DuJsNqk0u84hy3p01dpBVq0fjUA8OIwSqRCRyf84tAwBnbPlA2E/v2Ay8uWoPvakf02MIlu0zb56
hvK6uEsnQi4l5Io6Xf4u8O7DYjatMu6gadK02M8goiREmORxOcoXAClr41MHGmkh4NQ6Yr20MmzM
VVEhVB7kZpP+iw7gHpWn2escFI83EKu1DND2z7jnPoW42WsEQxzIEO3qQbagLzJ2rWlIQCYCc8ry
mufqX+N7/2L1O2aYdWrPZpZpulEXT9IT38cs3DdK7kFEIhugdsPJh+KpbVCdGIRVLeFtAPl2jxrF
EH8YyRzhLb243YEgyw5AmJYkHto/EY35nXLTdP7o4lndyw91p+iSNvCAcMYJ4pkY/Akq6B1X8EDm
RZx4YdTuyYDFY3RHZ8eMaYaDC3V57NgpYhfqLvgosj4XvdUE4peGBGlWofyAcLeiWQutcnnIAbD6
poPzywtiO0wI72XPY2jgwiONMaxTlbuVf4gl0i2PIPTAEOst+shhS5QYwh12eCjReI/E3u/DM6TQ
JVpL7AyOP3Q6PgqUpWWRsIhl+VOwcNwPWGysgoxZqbijzmKA3ZC4FzfZWRDG+4kBPGcDfFW7a2KL
ttmgUwZsmcyzRFrNYcdP2HRNqZUKy5olkPQKYIx0JgO2PLWv3epdur+FCmy5N+9hlC4nGDwljuzk
um0jiexk2kxik4UJop6Qh4FoA60LeR/Eg/12Q2mEZX/J00O67ZYv8m8nCP5lBd/8792PbWneBtAi
VXbImTfrr0y87eqeprlVMejcLw7eb9DeqEPAhqjfx5ir3L7KIr1assV4mMOZ8Ig0KBZtBCLdtNbM
7HR8G8jrY1gGJUBSbX48nwXGyxvO/hsskiLpGbiBHeVDG2mDh5dEdVap9DPFyQtKiaCIgQ/JGqmQ
PO+tIljFi6WaZwmAkAo9lsb1bLoZSLPnNgP8Ux/BXfzSAx6KN7NKzpUbp8/t5a4ugTha4tqJHNGp
VLNPI/4TeFyq8cCvWQvntPe7CpV/RE4hySeDFKfCrJ51T8Wekcm37MAgL0BHQWDfHGI7KOhFkHDP
44XIE9bZhW3D3xVb8aa9vtwlJwleCynaDBDeJGclJUBREZPR9mTxT9+iGCwj0OhgAFL8f4P2B7i+
X/nt8ZdVGzIpXRwrtzDq1YLZo7JyiL30918VB5SrBY8jCIOmYYjrBQFunWq0JWxkv2uKlKRE2iVE
+xTdNVovr6a5EIjgshV3jKCgo1ZcwAT6kKWAHbDiI3ER3YzMY2B6ArvrNlCT2Rly77Fsx1LWFa5Y
OgFmlbq3m3rJEe9Gu5qgz9QreB61y8PFX+ArYNpupci4otjpSjpeDCmP6XgSlqc52SS92Lse3MRq
y1xuWhtKXCqA1cCoxLI4gX5JqbF5/7P3P9SeXmEF2DEN4i90l76Q6NcTb41WY72WcC+UYhhbmt6w
nIpvS6pJv34tlS3xbVDrpHIHDh+x7WGQ+RddTkgJFJfraNLRumeS74yyh3rnDyWQH1oMV3C6QR5Y
bnEfqXwJlRKeZkevxfPywRaOnw5KD2b0FUrU8oOYKyvkvZtlhznfcTPGHh47P7I59ow8QcWHwSuP
i0227fMvO3nQGHviTHSxCZ24/CWlpG37freLPBeDTdv7HhPo6ND6piZEZdK/2Nz9XiLwgcHTE2UK
3JIBsPT7LXwy6UxcW488zdE9g8rDYxu03n1FU8F4/446OLLQhqSAaq7T8QXJWXEXaeoZX8+BborT
CyOt6cWVO/x9c0aMU/Q3wNe2skEeA79Ym/zN44cz+RTgnarE42bvvYelKXiNxbwUK5UmFliKe7es
ltFpYgku2QyPAAJgumqqE/GdtRejQkLibRFgnrwJQXMdMbOfJBC8Z6f5NWSkMX7Gi4bn9a9+lGg0
MNPL8xyxXo8SsFkdFIhHOzQ1XHvan8ixTd/e5aQEwad0A5hPhYVuuXwrClxjuM1n+aMtKJfejbV9
VGjhhaBZ6ffzA4zVL9ZSJKcriBabGs531XDvkzrow/llNwnLrWfkHh+rfqfhNvjoonkYS6qgj6mZ
YGE1E0zNWpDykfVqiEpSH8unxL37WqjuN8bArJFHW1W/xGsuBr+20h3iix/N0cEGZO8n8NF72bWb
5dPmBQ8OSa2kR0wO1X7D+0VAlYUSVn9zE06Fmkl0wyGkJv1fG7xxZpWyqpqMChY0E6cbNGgc9d3c
deewWs0lcsKp0qs6Ncjj+dqM4/eUjJLqh/dRo/Vqxg+1wlOnWZyoCHJkASzxZnxeinUu8OKuCDLV
bbgwZ3ZlOZJfwm2NRy1WPWzk5YWeJH7sQXJyNKmzeCVH/A2B/Xs8ylNR58FVCs9ocfJy/CP8JQiE
Fb/t6nulGlJQbTrNYTD34qQZS33sSbPVxv86EwnG/FZhAo8OBKlv22pLisocf8E5Z2nImMBA1CXx
BFZeZCNU0RHOsO/EZ3CwU/kyi8IH0s3hvVIT1/LgDk1UwyqpZjybD1Gl0SeEzkcDXxSjd68rFYyC
BzxiLSZlGflVF0LbC70/tX1lAw4s/RjeIOYHtubsvQ9ItsqyB/1whGr1XKofDHXkCDA6dDassHb0
QyUxM9xUeT8e6exJ0jIBfJFyB2lY8b1yHYCIPNhBjvdJjTkmKopdLkzaobe+Gc0MDfDrQaeMw1Na
Lp9KxXTNHvI3NP2PamQ0cbFoGKhoUNWOs12PzzDF5epQm5KbmEf2jNYhqSJRr8fGlFcvuiOUUAb4
lWUtunwdov4SL4qYdXf1Cce+XxNzXfOyhZHlYWJgd/c2Pfi4Nds/5SvxYiUXXM4AcEKl4ImgzrWt
4qq+1ORVsnO78oGGrInPPKmf3sC9qvU0sxDh3dEO39aATsjvblab6HKbcvkkgTjzszju7PMm7Yas
6mmoDlM2M3lUB0tvHdZ3ilbaWSsct0r17iIx/YOeALnEyD4b3cax7/bc+UlFUjLNMLViMfeFsTj3
ykTDLEH8wXEWZtg8aMWL43qCux2Iiqi91N5DU/PvJHuU9vp+0XU2a58dImNdyoLhA3dGRPYtvpsr
57D6NL1zJ8TOALjsptG1PPaELY5tU1k3uitlfwWymyVahk+7wCo1OCqw8Nq2VQUxbHie3DOlN6MD
f1UIGWmzQaq3e8nAiD5ShTkQGN3XZ+AbtHJxfpGdDrtcshUMl9rvJiPZrGHOMfJbx5TXreRhc1LL
5MYbzIkBLA6l566KcHTGSECWTwe2XNNWzg99oXMINe0Sr98dWpG1udlTDchzQGU3tay9hqJDEYrD
2RnH8yH3TMlIqlgWRaBFPFOAMvXyIWd9ojct1sl/Nmoij6bCINn1EkMHjX7PpY0wJL1y3y5o41Pg
qD7ob9hzheydOJCe/eiqGH9NNiVCoce3sZW0S2fHmbU8tz2n1iglGI1/KnkPnOrWjDXCiss/mxBb
+Y4j88knI5mpAKSoyu2RGKdWkpz27Xxj02D8ssbOl0zcNtpMZQlPZy/53Rfd410Io39NmH61mwTT
tHF4H9soqY+TxqEolSbBLMzYrsqIf4cBqJ967xH1/CZjUJMJpAgvBsUeCFElb+t/ZsP3OIE9Ahgg
9Kr9Y2fr9wIwVGb8pl/vKXI3QloRHkaXeGvqsVseIYa4EPW98m/4LKJT69jbahb0JfRuSBWRoIc9
hUti/dPnwDfbPg1OEXoo22/6zLkXssracnKhtrWPRlzM+WxaMTpu8wNFkOnqqPLmegIFD/dXLeeW
4T7lyhk/4xtpFItiMtCXJZ4koRCD6s37d5O7uReRLy3JMulUO9a427TACGf5vsfI5hw6LCbW8jxu
LNuCl1ushGeq8mIDNA+ohikuXoCGHeBsfiGm+4YcQOmIdxD3rQJGAnthqFpAtTbY+jCOUzAa0Utp
K91ha6rBlRf3NLSJkTNcBv70G/TF6QvA3uNIaaPRdX1k3fqKnBp+3sryR2FlL+Z/jyWs86SZFyZ5
NUNje/MCXXCW5JO+asf3xBvLHwPbv/QWiRiRhPXDFMFvYFr0ojWFVoqfp9NR9RQFowq3vA7XTaBC
2HSg9lsuIBFavAB/FbssSLcEte5JytasG0Usv5yhASiFF2nT2HQa87zYRUG9p+cL0kP+QZ6gQyq0
ZRxeU1wY0KaUK28qVY80XTGoJu49rD6LbzUdIFgnXgkchh2sKprABuC+lGI/6PmFwUtllnRWcE9K
XgCqIpA0kUob14U8sDRufrFlpDxIqRuPxdjh9kURIkqlHKwD2eMNSp7qW0i3uFvBYZkv3hmn5XVG
kkFPbdMZwjJPyl7kN4NKBZqN1h6WgWpS6zJEpjv+lJ/ViT8ZTOQJpVNHgFdBKPtBsZmE+yTuMKuP
46cruwzImlAKfZ/EBus2q/UJTXqC730MO4/o5yTWHluDeHFW5sxm3FtxylQeatCewBsJ4RYW7kvw
bI2n3lkEYwrm/Z7K9oua0+Tm1fcm/S5+QYNRjDoXQ0Per2dlkNJeJErnPJVhizfd3noArpUOz497
X7b+4Xpt8tcZ2FBO1RNOyadWVNqLEZAjSW9OnqJy3wNlqj94DGy/PGFgJ1oVSkT4Ym0DhZW7uvbc
nK4wzk/xxoP2Ao2EQoMrOItupgF3EXwn2tIJ9P4kdB+K93fexphBl6rTglARNlq6dsj4oKbpIHYT
kmNxW3f0FnyarQ71AYfNrl4nyil2E10gXcwcLyfo1cl9R9kwIgx8JrOCLl54OlMNmGCiUtWDTky8
a3YNZVlBA94ToZk78f6CBLz0/OVB0XW/faj3DnZ3TnS4phbsUVUYL9vBfqeEdtuiiU0SLp5P7S1Y
VT1KracA8pLypBBUNe+DAFQM8/DuNRePFC6dhUOhTHGo+L9qC5FHVxI+vlx2D26osCdP8SAbda6T
afDDIjNw1zuMzLHJ2MlXc8KhFG27K5RURC/vgvF5AWvljV4BlwddSzbQ0qkFgQ3kfFzQhp7R9eJj
eovdk2L1E/4uq7kAEMtgbwgl20yp4a1x2lcYuj4nCq3/i5shcuiO2ziW+mCWdVnJFqRBteltpm0l
nrpjqnCnwBFU7aL8TxdnnTbQV8ORAc9X36MD/i4bgceG3cwImc9FaR/LrpMaw+xHfwCwnvlR1YN4
9GghIqtf1egMZLQwK19jxx8RcdM/oe2OO2+xEEO39dBwrPx/7jLxCP7dMWwpBihR2s17uWjRAJ3m
7pZty6kJHwTowa4W1EOzhZjK3XRBXOZsdRNkfyMRYfonRUJdSvoHbA2SO2jA6Z+4D6VVqFJ6avBv
gzmjJ53fqXMYFcwWColu0BbLLadzKMXQatxbskQNvRSdLDRRJPUeZueoeKsIMVg31ZUFTTdgNdt5
hjHc7W7exdA3RnK97jf49MuC06/lch5HcKKjVLz1g+KujvN4MgoReJq81wXYqTdnNgv34pXFMG59
OWrZLKS1z2c2BLvxHRKXiH4O66KtgBdvUcXBC2/LiUxbi0KkmSSK2DfwSluTAFs1qoWmPQ/Do/2y
egeOhwCec4eoVwKUJIH3svF3dy8mjLpE5fpspu/LIaoyAmLIhvvrdhJxsBmLKUybezGwWO5zEwQI
UM4l+x+Z+WP+pel349K+Z/3yZdFJ5QzQjDGG331JmrUAbuZpz45ZnH5+sy0vIGMxRmV1UsLp0XwJ
OktSu3mD5wB32BhHLlKPzAb/y6U5+AFH62/8yNkVQO50vMvhkYuAh8oC0WDQnjl4lUS2KQc+48e+
5MupTp+JzQ2F4s/tjNKxxNvPyAzNtvlsOt78cJGSM9zg81m9+hqmm1ix86q+JiGMhJUyUhHmtHkL
K06tgBBM6BGbQ8OsQXkMzF5bFBCGjTa3/Nja+KT636KUjT3dg5+kyrwW/I5pDyNO5CTbs4ZRs1j/
bEl/Dmp7pc+WgGCnJNtWAI6qyXMZWBmibZ9xp8JNzaPWaviUB7F7XGDUGvE/uO76KAA73GD62Aqu
EJfv5Zl7h8o1nOrkFCfX2CcpD2dr/JvrDnFO91rVxr0jX763QgRv3WGUHbMoUcx8uja8f7TiPbJo
6c/7QyNgrYrzf3tCSfMXybGt6caCA6yRM13lnMvWCDNwPBf2Lrlp0OJYJocDWfjngm058jztY+3l
EkfZ9D1NkH7Gdoxg1YmwKQGQfDtwSFgMGf+b45JRwv/RHIIc2XY3YR945jEJf+n1TvMac0KkADnB
gALS9LBVnmBfxnbggTdmeldAwM/llv5eKZE6nIWyfjob87DtR5zNrK+hOCvCbcV1u3+NWBUc02WV
xWrnJySzZFwC4VwcgJykBLz67ZOvGAJfE1koYxgHnOXj+R+45vTLzdBnYxbbpavXCwOingzMUDGN
lwFKajek3eeIKznliYAx92wedsRWQg6uIFdHgDHixTO87zUTBO48I8NkEeg/VpsWT17GGfTJcHRs
lwXTVE3NA2DzuaiqynJjfe9oauusRTEiLp5YqcsgbRQUebITZuQrk447KWw7sT1YI+5PTYVuQ5ks
1GRl1oI04YRuSdoiKl7/7LREb5UkHqgbEj1AEkyGOwLqw1f+acN3Dkrm5FSEHhC0/N+oKnOGGPPG
6/DIRKP6zDooetMRAZhOsh3H5oGRJtJ0wSFkjNkVrirpCTYRliHmNKvNtNQw+ey+lSSsGQS/w3Ju
CcxL2AAaH4qGnVthkOb72gau5d/WCJTsGqztdRxSM5ylU+JLXFPJwAJ2p3HT/lOzLeOMzLk6lehf
Ji/JmhuTY8bG8Ulz187pDcnC//Sm7FnhR3/DYDsM5Li8pt3IIkVodUjSbTaN4hDE/EfrckqSqSXj
fT7VwVnJSi5zb1LutET0GHgklil5ND4tW8EXPSphlv0Z3VM5NuAv3/YgR+kOkZjxXhv8iP4CtiwS
uZX2DUSrn421d13slpLLYL+pwhFqBI5HI4gIjYQw3tI3T0OIngkb75dmtrtpcPrhwJvTVFlStWCH
vxDI6lch5RdK8qHBYDvGNQF+iz4jjeimMY7qntbBEpSaNg58v4G6CMa6RRiea1Mk7E5eP7Vub17l
0mAiI6+4nsUWFU9es+beS8cTjP0cXE1U4mux9uCiVGuBpE0YRq/0lfU9/x0xxDmgMwGxvUfJmdBz
kpfLnjGDQWOz/Hjj7hLjmgflaHB2Ob/M8esz+peWoW0BW4uENzfxXqIv1aF31gjSP96fSwCmcTox
4vN1jjQ1Q40pr4A3+r5ThgroW2J9+ZJcBIJCOQsyBuzXNLnxm07Zb2gFxBifwN+0K5j+lSYGK3HY
Kx1yiSA8YNpLxI5DY4+hhwLJ0nYD82br8CUDxK49NkDQcmWHdP1v1qx6i5xVh6+R7CjQBNGgAqe8
dN2FMLMSgpRMXjcgTMNhqpnUqaMdZtJ67L4bhgNofLiIRWBNa5LEMJ4ZcXKOTQrokctsw/pUM5X4
6xYpw5SM0515RM8ZJeXJdiiQjpps9tpYIeIrmk6R5lqcYyDbDNMJXs49OQ/aUZrQU7q4hIORbJ7Q
3UnfCGgbhOqkNx0Yu52RSCJh5DvCDNKs4T8GRMw3KimjUkWjL6JJha3p9ksvcstLj+NkRniOs1i2
3nZgq6tqGxe7N+BXv1kRYtvoHKvAabVnQtXqhZ3lsWWn8xqCc+pQDU30MMUYo/B5NmVPSW1xBfsI
QQ7c9J14naNfMna5lfMDpuY2Rb3vHRCcCZWV12Ef/ON+qUQOFKlas+DzaDDaKzD3U58S6IadXv8w
J+lNwoRQ7hRoNUbIF8QqTY0AafHvKqXDkcs4Z1Z6YxRlQ4OP6XEhGZNe528B7HifkfV+atbEWHTi
pwa2jeuf10CWSYA4sHt2KGcZOyYekk5P3NVDwuXzgnfo5toOB8KIuFWDnaNusRkowgBsa6EbPAsU
0TNS6E7qHtF0KC6yzLwzaVIYz9CSUoeGQwknSqRWOP5zb3rISU+OI51beQpFDUi9gcg8mUgUEM3K
Jc9JJFFZxBuNS1+MnyfZt6EwX5Bq989vXDQfL4Dq0r2Lpq4Htb1QMWsf9K8V95vblyfyDri5oWYO
/um6djMjO3aIbq3tc3PrhBL4muwhR588mCxJkm6YP6iXWo9D/gZIRA2oakSaUUDkrxRXRCNJGcIQ
iLyb5/dltLEkTDyynpR45IBXl4iBFwKDct0Y5gVGYIbEwpYePrJKMUJ6qh9gg9tkTi3I7Ujzn2AR
K1QjZBV+KdsxP5HNSLyNS7ptrzrVPipdOt8AY5OVE2zX/128/jgXuA3BGj/0CgMmyUQZh+lsaYPa
cZTzM0SXR7ZKilNeHbP50vMasRXztOnmgcqTjYIsCNRNmFD3/CoKJrfBBgVer3CdBvR8VjqXPEP/
nw0Wr9iCKsLbQm04xSlbq6WcfGHS1t/oJ871EFB6KqTl2GOF8V7QKEhp+I8hgWxcLkgjVIi6mrFe
m7v7ILB/J7raJlqXBrtQgdDR9pulTNxPlJ9RhMCSZdkkg3gfliksP1afa3NYj6YxG1w0MZeMGi5k
HkDb4S1uvlIDyE/l7hZEh8y8cK2oHrn+IGdAsvs3+zWNAg7ENbCkDUb/4ExZDnORJ2kDzjoS0Jzf
rH+i7AtcRdWmC0Bc43USAaefZpbXoJJc00ufindCmvfvB5PgIE9WpA8sAkfafJdmkUQLnkm5zxdI
erbtzFHz8E2a0/Blmn3DN3Dt8kB+bPUJXejBZTBc0EW74Za1Cy+pyy95NVSbUC/3zHjwYc8T+EfR
VjKw8r5mAWxJAClIBfkT6vhtit4njWVPmxwt8Y0qsWDlfMnppfVT8VLhdvhh7HswSas7iL392RO1
PZqmXjIlzS+AJE2Q1erWISosn1pmdJRzyLBOG1PunCO9j3hzZ1FePdj8auxOKNo1Rs2hMzRp9D+R
NnsXqtbWDwp+8VH3zZD4D8y9Jfdhw6nRN4tiZZ9//+nMBEhkFO9HETwJcmEKiF/DvEyd8Zn0jjkA
qciH4e4EVb+3YAG8NWSqEtE1vzh3VyuVqlin9A93il4P7m6k/n6QsEVHqiABbyCx3iwHcQ0vJNYO
8INkvp3PFJ0BveWHxckdIY+gkctVyI0Vpj4Lk+YLyg25ZWXSf9s451U+wYufuaiZJ0IOAY2trtnL
tm/+H7WI1+JA3mBKEeV13N2VKu5pN+nI8s5ustYeb9fF/hPzv/4If8zseHm2WpA7qZ98U1p4ijEt
x/yTSDbM2DpDjC7svnyjJQuDKL17pKeeTklJM/HCmrTgzO5JFaTEEV9LmwLpxcPqLDMdC8t4XRmq
2VaS8ycdmsN1iU5JEAhnwQl6adCJXsXeeU0jEmFc+rKeMJzJ/TDIXKAvcgVhGE+B+BkMJT4n+dGy
lkYADLzoL7uMElQk+eh2FICu9eJIBn7jbRA9IwnCXc211LUC7tCZOoKZV42Fwrbt/sXi3Qgm3i+M
gW1OCVs//TPZ3lsdATylcXEyBtzgNSuBY4kOzIRfn7HOa4OnN7nTqqUhAzYNg2oV8/tzcrt8JuEa
6Esz+1uZZnmRfyKacz4b3Y5RJT1w/zHt6n6KP/v8n74OmwrmLHhcGgo7VgK8i7dXh1PT1QQt+9Ia
ecsoAF2/8179mRlbuWSdyU+5X4M1DbSFlToM5mMmECS+NVhFmEs6S2rKLImu7K3EeAniprRmBaT6
7aJbY0ZGZXWHqH7pv0XEuhjwli7X0xU8l68EmbD3kjzqoYTBmJOO/nQxSb3o9o8a28Qy+zSMD0MH
0auuuuZabG7ttnmIzQyNVtdkrVCu/FPlmvkh1VHqAqPpLFr4sE82LU3Y7Z+9pMOcm6o2H4P4CUb0
rs52gUBo69kEVprl7OkwrVxjvgUNZqDiX7adsdzWgY73FHzUwub3ceFJLKsEXm6QHQvHBRpYmyxn
GaZrmCPaxMk/zWjZwq8Vr0qgukvkOAiJKselqI6WvGFnAN0SBBNtI+J/vbKjwV00oS5W53NsI4I2
tRNQN64SOAr/KpuyD/CdHzqjuhNkxLknxgXlLggBObIKh24tcu5J1WZ3gFdXaYk6yie+vyIJVu90
cCo7y3Ilx2fu5sVST8n8vIOPRH8quajZrYjWJGOnBRrfrg6K1k+rOuGqoREYNySnSYTQPCJPXZ3z
gOYBTlsn+eV7+RVO9uowqhJPZJk3TdW2QqwDbxqK9dqIbwJp+Midahj7aHUM+hUNYvcs1FcsusKE
ktVrdm0KwDxqgAaMEdfeQ75njw3SW9VLl9dSDNjDg5PcQrWjAbvRp0gbJvm6oLkgPSbcwn3ZJnvU
9J5/6HxWflfSnvlcYBbkl63xRXwG7Ep6CqIzk8SNg09xTcPIuzhW5YpSkYurgQ13kMplo2P7TWSD
mJRzhaBHuXAih885QRED02TDsL//QUEyeHZddHkNV1ny3p90tvZKUzC4rWLIhG4EOI8LJK/CUGAI
lFuS16bMCdPg/ciWsDbzcsztGtr2f7uTZTNocIAz08bAy50zcKjpKbjBHz8Rd/OZsSgUt60g2rrr
hRhrWTE9grXljhW+ony/BcMqmB8bhG/suCGl5Dd84Nqexlb6xYMgQZCs37h/vjN5Dl6UMkxuZ23n
yHVWxfq2+vejlXfEN/AGzZGkMKW/qF+ne/OUtBBiJ98C1BbkAEiBrFW4pHlOt7rCTBupPz0ardTG
ljpsZfjJQFoI4rokGH1PaoF4zsRkF2nbHDIVJH4zpPU9Jy+YtY1jZMH0CTkJdNBAFU95cEQRV/i+
5FPvMTgwGjpPkg9a63gJtXtDi8KAq2vsv4vS1khl8mYgSSg/eTEZIM/0MKSU2K1e82KmB3NCmcPd
ubNK2fMFLKX7NwCJm5qeyQvg9qr1fFoCmbySkgdYt9DX1KqL4o2g5t4gLfJLT5V3ft4SDS6vvRoO
AnPmKt2AeTOyuRwRmFmCgexzaaIKlFX2vvj958sahKz9nBVl8r6e/Qrz/uocygnPQbKg8xsF6HjK
t6t/U7S9Z9hKPJXpJQZKAHa8kQRaLvU06H6RPqUAu9nQMOt4AlCv4Ce6RB2svMBdJGlgmLHH7pml
l1Nz1RZtnidCYo276HTbSzkiVzR4UduCcMPSn+iC0kuNAIBRf4l1oPEO0k1Y0nZeQhWzO82p3XkK
2+XvAAFhH0rbDeU3uGsZZq5RSJzJZoMGVGetkzLKMjlrZJ51MBrERml36/oPhxdrgvCmUHtAdW+o
KjCtW2S+uuIwg8k9uHxxqjeTdeafOZpxuEx5oPNLtvtWRiZ9PJvn2Y+MNc/UGJOsq3kw3Qf2o+r9
TjvNslWQ4RJRV6pDHfr0FYGWN3U+W3bCMS6x1fVtxpNPkJFvCK7b38BAsRRb89yrrDhviPXQEv6v
vyFInfTGkWki5ZGJwtd0QlHHtcYyLl9G8KDEbEesCxlpMoDfx5WLcnjWUZTVpU8qgIJVwdktnPLH
bOdiEoMPHMg9MvF+tlnHsTicQfd6BdeU/n/TNo0JeR7wtBldmRNJy2y10SZ0T/4fQplUJk7dVPoe
WxUAwkpvYcCSDGdM33ZtjA8euFdWhgJf9Qj9C4oOditkN8nHy3iCAVu2wX278yu2DxNRhu9xvagc
OtzQLq3yMPH4EGDvJdi5wIsy4eGk6ag9YuXukLmyu3vDPOjHKFjzcx4d6oChZ2Cl9zBvrSKJ3LgM
0kOqz0YrzbxL+XMEolms0OJN9PiHOevd74hs55bOdUOYi44KXyuWKH5/UvO6zHdgA/sn7ey/qAit
t8qvarBCT4/xgTzbCygP0vJN2YdXLyklLo+sDxdLhDagM/5Zyd0Tg74xhMssB6n9BNfosfTs7yyH
T0Gszu98jcUcW+V5aCWyYNphB1MekPXUSFJB9ImlfJbf0pCShR361aRSPUIkHHlqB3qJreZscqLw
Kskv0zR7yVcwFgkWOIH2ya2uOhvX4x4zrgF30sDb1hAKaie3mKC3Dji5BnCNRXl2YnRxCUA/O50y
Jd1wjPOV7770iSbEUlbboLdT1pGSia+i7ijKu6O+4Pfw7t4njFrZi/xlb8Z8HnTJ2azdX01D5qdY
bswO5hzc0bwGqsTD57FqT2xCo/IOhVHDvXuF9ts6VjNnHiRqmfDXsdaTjymY4xMgrP1k7BVim7x0
XhSvjdhWQg3334sXXZCbdRFFxG1wtSLoKXg2Fqv3SH7JQm3Lfi1jnRlvLyAEgwCuLAquAf2FeCU+
MtQ/t6P/h9s9GPFzpHcbhO4sYmMKAnfIx5VxVQXlL45bzP2L6kUQvc1Qo44Zv6jRI6q9ljemLU+z
UP47zTgYcnIzU6lpEz+tVvtm3Ep9vzxcOqA5BW4l387wkrVU06wyrISmE58xbTlVlM0KLUqGCMGK
x6T/h6CuBID59WoOhS2Ko7hmeRUWGUkG2AbZ6BPpGgz7ptvrUO7y2KWN7XyGf5rf7Ri9BfTYSW1z
XSs8oSFuYiBk15wbkFPGyKMbwF6FEoP+RyyHzjZXdGEVFbngUw4himqhVBT+dbm6IBwtE74GUwys
6hn5U9TG2OJnrvB2zvWApmbWVul5/zv39XbFzTdRVgumRR6/7j55BQ6JIxxW99U9xv/RhLSGFIJ/
t7ISD0rJS3rOdmkJyqTb5gmqs82carpA6ogTjS2QaiqPli3lWjI8Gzc6UQz8Qr6b9hfLBdt0H2sB
ymjojDVc0a+Xdyun6XvKRAlgpfzpFmlHluKAdr6xl+fiIbfxziLAHlQb2EI3n/a/SkkXFmVqa124
R4CKePPKfAW3EpzuHMTQV0MtPBi+J83G1C5BsENrQGYyq6Erohi3uaa7U53xLv5T2NsIu7zMUrQk
2a/XBwafgxTGHy5EJDU7FMiScsTINy3rumRfBHJ64uXySAbHbRPGYd5Cs2dmeqgO0Ns+tekJrJJB
XyRRsl7CoC6Gr4lkB8hklwPwr5x5UnXOtqdFDEH7EoTt789bSN5oJuo3+H89FOGeSBj2R2pdwRKL
37NJhycECF9p7akCYJqSA6hYirj75m0OLDGX6DbHG69tXKFkEO34MCJje9QLEWx4IJ3lAElpl4E1
Wueo/wbyIGlDfIADLpIgTX5T5N47FYLlECAwcUuHQkFPv4lFYXFcGIn9/x++A5Uo8Fe02gTB/URi
rzteqIqrXoqb1Z8rFUyn8R9LZqGpM7yhxDdXbJ1PSGUCKCG3vqlHXARe1f8NFVXSZZ0JNdokwmg8
dYws3SdzMGcsbH8eIQ2EkzYsqswY7sNgD75Jn4N9rFXf1zLwS2MxMIYZapRpHjT4CiXn/0QzEXdQ
2zOVcI9vzuW0N7Gm/iDyBkLEsdoxfzbBKo1KsbxJ4CJ4TAaeOeWX/FPsw2P5D7wotHS1ZIVoT+vx
ycT0S6hB9yBDnt2z74+69GM8bJMI/uv+jwqW/slh9/14ndqvFIhom5O07IWxhxylr29maM1zeoFE
YfYkf0WhQT7F8M3rXjV3Z7MnTaUKpIHgscZfE7GZ/Yyvqe1cwTpkvWzivAEJB/X3GINCtnppQrPy
GcjqnA7FbV+2lEK0iLgmL3Ion4b3TPe0NxuaMF6i1bXC2l3fd5Ts6KzArNhOR6xAJDX0agOihNDH
lJwWgFxU/sn/EW43CO4BvzP0FG50/ByhFJQkOlbCTXGjxRowL+djl02SSMtQvnmBFjW8pQmnLSZS
BKOhDwFF2/W5UH6hEM027tGbBEuZ5sMEtzW9IkS4Q4fvYdMjRkaUhCGoCWlVexEVmQouvlZcrP23
XeIjLIRqfacdgCR7nI5z060v+wY531TfSGOFi36lkVyI02WDMwwVJgPVEJ9TjeouFaHuv721gend
X1fjenoznYt+xiN5z6h8T99Uzl2Q+JYeiHEIvs5Ne6rVAusxjkl8BZgULCpbRSzFUmVlClu6zKOd
Nemtp1iJwcfXBBXPLhtn/yeSDLvOIJ8k1dJ/+GZdLfn8xEIhnKj3Ex1JRh5LDYTF+75lpaqO9l3M
0zU8O8x/ebB8MoBAzClXVKG6GrZdrsvEeZLg4LV4fXYkZIg9zpe1YSUC8tMZ0TMeHAIxgEIJz9RC
J+aAKif/y9FwrTDvGGwCsGBa4J1TtWeZ/MUdW87M1L4HV+XLCdHet7rvwND9e7rgNfPV+djCOJlw
Hl6ppKowktKjB2dDxwZi735qdGC72KjeACZVFr5SJffWoP8G3Ue+KIxlJmM0nFwP8ZilCgPPRhTY
oYUy3g9mlDVTElakOq6SLBvIz/17xp9si5Ave/651/mfL5OTnApA/wPpeuBUNpUXZiSdcIH+QFRy
dTEt2+//8U0AAioP7XJRo+p+1KNJcoFQydP//JodMvjfdNXdvPgkDLEmE9T74/Yc+juF7r+Voe/b
LZG4MRXuc/rd6f9/BfkW8EIbBoihAc1LMPTK2kTh93/gSQEmW267hkp7DEuSKhRJDDUv6MJa+46J
g7o4dvLnGOoAnxgfCcbIsihhPpb350T9D/uxInOBavN2vbwYdU6QFI4X7Fr2KK6rKcgA2y472OdP
5QMm9C3ONK8r2/Ux3DKU+GmG7ERpnlPVzwhk97AnqpBfQ4rzrTsrLjas8HUJi4v4U37Zc1/P1BSZ
bAOvmOPUI/M4NmNRKt9CjjVwGaWi58A+5IbgTvaHFFgVsutDtXrueuZPF9z7jjusGk20TkArO6cQ
0jfJzA6hakZjoGN77kTCkMTlNuFrxWPPijobinVXI/V04vTyzN9IeQ85mHZqj57T19HOvZr626TR
hBeXQPNd9/tUFzpIoX5UCK7D4W0ASbz3J3mQGmEDX1lndST3LMOswq0iICyGCrcnlb2uFtkHrsl1
s4yLyVUVEXtE2T6i1n+8Sb7nrPOYXSMO4iU8pe5hN9SGivRD81+Ogtny/+Jgm4Cz0msrZs2W96HI
RSqp1GpNCo9xWbSs4ryelBQvvWLsAsboY4sQ6/RQ7AV2o6O8Zqfb8MJVppcsoZwvHqTtJJcchMNs
xYwXTHgHh374fe0cIiZ3bWU4RkmK6G0CEBxyliwYsoXcdt2PDeDOWw2aVM5h8dctEcjjs5bPcFAu
2CW3hVf3km9ja7uhmUnj9JxUKtNjr00lmuiCY4BEsHYhAwqeUhNCLntbm9lplkgQM+FQsQG3uXiY
rcIf6LTJy9GDUI4UFmpd5rWVUSUDmFlIFTVKpUeV44wrVubK+/UAzE3b/nlM5SFt2kUw9i6sScv8
NGBYWAOrACrTGLMsv1rENuxFpM3RgPwQ65ERlVHUezuIw46uHomomeYyNwWmO2L3T7WkNrR1Nx9Z
erEWR062mgje/IYF6pK3FkRNQ7Qs8S8ZgjhWGnUgTDNPPniEv9ZNb01lTmqn8wU0NDd2Im2SzLWD
WLBkBgTm4a4tujrB28emcp1JJJ6f1z9kL9l9pDPpm7pnm6s8L+xbkjy1IkRu6efI55BWOuXMwoMM
oDgCXy097zQc7fsqAZa7nX44LnUF70esjz8mN01qSVjjcqLGL8x10d409wz1IF5hP1uuj4B60Vo+
b2iswUSHn+C/mzxux4ZAjqHIY0cfuH0wwv7HM9uwcLPB87PMozaeWMhH7PrQXYZrCkzXVRzy677p
lkGr0ut3L/MzR39G68a+/G9E4VBjEl30t7S43a9DrC3sWL8fapPwHaldyNg6aCIau9P2H3V374ZU
ZJEq/UZgdGIaVAXk2950tRGGbowVZ/5+A2rkk5OBnvGBOy1Ii67WwyL8ddPidWduam7aqEYZKFyL
+wgWahYeiMJlb3DkgxEnUIKEStkPgP32b6NoUFS7p63oA9fnmq5eoU9xqDkNlCU/LQRDq01UNTLB
enJSW1agZbPpKoyAczjr/jZtc/pO+JuAaTCWyBExqS0GYDragFAu5RLw9GTVKL4eAcaoFk2UZc6q
BMcxb5O0mIeD/dtrUHdW/iPln/HBUz2h3xXCMCMcRBRbFvk0ewUcYypLpwrvhBu4lK0Kt0kPF33Q
S6DvG+eoRKDE0I0oOM9q5THFxhQj3EMOPh31dhwmGU8UwVvsFAEVkU2fUZKCnE6k5SqalhUKqruA
p+k52uoyGT6mXemmY9Sz3g5rSdYEaylpop3rUuNh0lHxVSwv0I5OpvLOUq87YTDmPgyyrhNgnHoU
+7WF5hT03tRD+Rh7PAjbbeUknYYcnoTpDdCJuq8Pm9XLL/a/0DT/Qn2lsNvdg79CGPy3FIjySvcV
NKPbLEJgHfl6D8XiWSWSjXsllSS75XEdrR5KnjY35X1iKy0m6dE6y2Zr+ZBAQ6jvFQgAZBpOSS6i
ZkWHlqf+7CU3LxnukeRGxlJvifFEAj69n8jDBJFxEWEgOUHv2ryMyV5XfJ9/0pyoy4gmfw23vEK4
7qiNdAFqYAwxQaR3BH3qaUqRXZhnaN69vUdyDsZUIPysfAbwlVbwzPvKKBNPhVX3G5Zu73mAzLjz
tBhvtzio6LxhUwN7lQUGOAg9rLGUQnL+4JxQuXV27vc3zFS5bwDy0IdPAmKOBExQbuV4vGwb6Y2v
ZBkRWv2Kx0h5sDuXpCnnJmoykO3USfJIp2YqsI3PTGXSza3pjAUl0Z5L6Ptro/aStY9qLZY77FD4
KfsinojW94rGalnl9uk1aVnw2y9KNwUf67klguygpMIC1KCxpZwXddCeKJyqjPTWWoh+ZiKih5oi
SpQTCGIq9Zpow1ERk7wR2uYSV+kagOhZmtHE9oTwCpOV/ZbbpO2jezptsT5yuZbeMljogJp+67b4
CT5fwEBC/AQsLZwwCgEcZtT8tHxJgFUzFPZaN0t5zHDKDJWEyj9BUiZja3MqmXf3KP3BW+wvBihU
y4fhvjoKi7FqbGGuocxz+fs5Xxq3S8u0+OwBFDpx0YdKkR5n3NnhEDkC6Ut2tcoG9sj8DuFGICfp
ddtiTjIMq79mUFABPdoPcCLgfZvQI55xtQv05V3zMrf9MZpFqgJ6Br7ysotbxehjtN1iQ9JSE4/3
L7r5MOqc53MzxI2Oj9kIU2Rua2xHXgm+yDsA2DYHzvPT+Asey2ajBPKWlS9VxlTizLQoFQX2GQ4p
dMtAr6wsyWPM/2iccp4kK1cO1mEsKGIubOhUdOTxtlooD/xD2XipCl0YT6xYWpf5W73kYpgBVG+M
IeEchbIVogrb99aqxNaIX5edUj5buO1x5emMmiNR6DGCbNJTbTT91W9/Qb5txW5dSEV67n+EJA8r
Om813FIrUTwqs00mjyr0mTPoWsylS66ICOZR4hPpoh+pr+HJ8xZfjG9JY/IA2ITA0uTY4jMwptxd
qCPqTAICiVMGGXVAb9d+xbFH4vQfVEKPFxhOoqIeIhy0mdBtIYYgrWWHbBLoqMh6jl5GEzgLvED6
1plPOnSvzHpGta/NjXb8EWriuadz2hQzrGGvjsF4IovUjRVYwIxbErqbAMFq6GdBlP55Nryr8eHP
V1jNRH1kDPKh7FmFR8j3vujqmJOGKF5IjKbcyQrN+QaGT3ul+87UXHRFoYaLy00JX8wsQuGhbLVA
+knVeXVuZBW2AfHzHT8i23YMX2JEjj3Q4itrVW16gPAstfmaRD+TBeJGv0QATJclysQ44bPAv9DM
8yQJg0vqR89BsEMUfg2Bj7YpewzULQncpWRafKabDLmTCsdYNxSq6+tuI2wl8Nz3GOfx1V048LPy
3NIumpPuyCB5wEH69q0Tfu09XrYkapDLV1s8FgEH2oESRSDuA7219VfiqPmbJSs4V2kaGtn2mZJT
Rj/2ZuDW4dtKB1AP3xe5/PAqIkoHsofn6m8qaQHI3JWSGyl1SG6uyJBGp7Mqd0pHPznZfMX2G/Li
F4YlgJbeVFoKy8JTj5gL73AmsqxaO/zWwkBJvEcJZVzPFwwAEdj6VaQhCvnRYHE+4fnumGPKqrjr
5SdGCln0cO5ABjvJmEXV+6O02iNyMxGH6iT8cs74eNc8SlC1ky1jB+aqzcDNfOJpeBhlOhM28xtD
EzXPs8Ol12rZBLjUWSuZhHqHRigqA0n9sPz5cfSB3zCjfPoq3IdNq02cwd9K/UEdNt+pAIGYKJmT
H3MtNaXgF0TXBh6CpdMSjLamhEOYUQGlfL21cngKPaHhCDAPFf6dbph5R1I0l8ZbQtK8C9ELDScr
2gDTJVpPuKptA/rNyX4w5E6KfVgsPxZyCEksuMtNn96wC7R7mpOrDkmRxoCugBNypg4lXRXRLUHE
FZzrsE+o22rBTJhUqJuoUDUa4oFYvCqPlVrrqgl6nW+8O6BJLuR5g31dalfTxaoJLRQpPDSXCN78
TmyFF2QR9O/nWQDeljjGKbBflj1rHWQr0m2eoJd0QGQdgzXQXiz1czgnlTCWM1Sl8/S2uND5ie00
6CtjInDaahEhfbNyxKnN855mXbxlvMj+38zeOkeRaqlEtbiPNhpLF0veeB+Lo+d19cgBfEs2lkYN
0+W2rwnk6xNJ1Ka/zSFHEz0VTx02B+GetFMF12dw2PubapMDkpXTu9o2/nR0GbfqaCezan9gGV6X
F8UjfdNUv+iYXw0S3uQ3Ctfhv9vqJAg3lNqLOKxN7YlLKwiRLvs1MXasvpxKc+EbwJXu3ylPko1u
mq0Q14QJj/fE5YZHOFzE7nVLOpUnrqY+guAPXa+PE0o4Hp1OYF/bCNyRQG3XWjmeHDTzvHb4CC6f
Yq156xyhQgiTnmhJb1TK2VftSK5hDWdzGO85M0ImfI4gMNVelCo48kivzR0N+LPXj4lgzkTCqOlm
cKug5Lsn4bbOxKYtRLdGMzjSvoMHfXcOBu2kFFAsI+44SvWcE8lDj0xsOrNqgvux26d8GKweCDXJ
zr88USRq6XrozaBs8F3w+ddVp4/Lc18nFkjeK39MM5ZOkgPW0fNihkKCK5sNJbVbJxFUU0OEc5L0
QJWpZ6S/lq/PeoxV7kRHDRku2/AGdu81ZjFH5MhkRlKfDvxY+8V8J/y9UUkBjG/GPGRhGnAEaOqD
uAFP0G/FH8YzTyJD9H7+Cdfkhsh8LG4DkwJ1Fe86nFx1zE6LKF8rDz8ZSW4KTiquu73OxOyjVJUi
EE761YGm691Gu+6UqkB9CncQk24yPPFPZriXILmYuUFIYtFrAZo2cMXfTZimAMbX+GykTZt8Tr2I
pSY6jkw4+2IaSqOPjEpqhkvfph1DVhlSmXeumV8TcCOrabjzILNxig8+txPsQnU6gCffDjxuds2q
O5mJ86rJY3va0bh/fH91TIrAUakpfux2tGe0F6Nyj4Pgk+LiPPOr0fX6IZ+ERSMhBoUrK4tMZdiE
v6IO9N23Oo5NLtAipGuE2bnfB05cVzu3r7kZIAtS2jljKQ5Llx8HZU5wK82HZ7oawIbDSleOMZ6n
SQlmvQOGvT6elSQMB8vPnXnnvw1j6DwLTINB2FTToNtaeoi91MO7oXpZYwmVz0ewjM61uTp+Vqzo
cxqGzxXoqW6WN4DyFSpLNJeGOyZNTCWflYel4DtB19HKbcfclmnUIxHw7TZKeH71piXd6n5RqSss
3Fxpsu1qbvEzf+UwWQ6xBxXcX3JTjwq1j40SWa61hNIL7ACcix3ngfxf5R9gRUV5NIxSN68vGIvL
ZwgTlmPW64XTdx1ReAArJyznB6j/ajRO8HiRcPZWPwfKheKIw8e/tymZcAziSkFVLrrYSj1m03KO
vTUhr25zHvHiSZwlLKHcDmIWz4jz9ZdMfhHeZE4KJqnuzI3uyYZpkNqxOa3z3ud1GFp7TYZjEWCp
gmA8duCPZF6zQWYxcc5CeSgJ2ydxS4iG3W5TPCtQ9NWaYGTAel/zgtPKke9C5zi3nmPb1U1qJMJH
WYBAsTAU+wIS/7oFhyRAFfCycnPnCCi1CIVmjlokS65f3jUM4cZgpP9NErp64mz6MokXcITS1Lg7
haemhP1anAx+2wg3lts37L3+1FzX/XxjqOqycovoHd3n47/jSWt90ShDQ0GEh715S4h+QSAWvdqE
kjGfYEWV40/eJMNkpRW/Z/DTAdOUaIRDVR71tuZzHtiYmmghM8+k8cM27Ar/51aL7WlBHp4iNXYD
BCWyxr0iMWtD3jPVvvhFI7hzekvOwBSksI4FiMQdVRcnTaV537d+G5E7vQltoTt3eD3I9ZNsCDI8
crUJYyt4NkGpTkm20AolrY3+QcusJe8xZFu74x4+yjcABgvmHKUtMLWQQ5aVKQut9+8oBwzXQWuH
ZuxL1amFQtcxD+S5yKqmY6Kul864vIUZf0I1xNp9syf6UrzQkrq9nMMEnaToD+maA3G0XRZcqQjU
lepf7p+8FNtyfdSieV/9MMZowga8MHo0udsftJui90u/pegleLLBI9VIl4zMUiNLVgqOrz0WyJpB
xavIuAk/d8+CvAV5ybBu6Fvn/yorwfE1Qzpn4yVrTn/kbINHnAeGGEbSHdDfxmuwiNHjAuwhSHte
EjZkU80HPhB69LEefl9STxVC/aC3+u5ebyulTDaci6xBfKOsgHRAtn7/QDI5jLNsZHdGj6NMLsQE
PoCvCNRDhOMhl+BT819/BHBcY8CD/bHDOBg4dJJS2EN6luHsH+Xl07/fT9YByI1UEhCCkbRKp4Gx
O49TRUNgpqcCd4a3wKCB9mVVbLpZV8L9QE9w6iVOLsno1CT1+UtigPDTIsfDLwiFiYPKJDSP+EGf
bz1SKwDOexB8bWGLTFNZQ56n1/MQ4PnqApsGt04zuFl1DKJ8Zud5hGi+t8QxgwsaNC4TwdsNFSVV
pdAnB8/DmCh5yliwGk3LDeiekGlg0aGjQdQq3hD/E9eYQ3yIp4XxMDopF8crkRZGSbPNVOra4h4g
H6+z8Int+0npU2lpOq2ZkDU1VeSRqHacPkCKP92p9AJ1/j5L+Sdf9Ak7U4sjccWiekb3Oxo0qd/I
Qh5m/T8jyRWUd8WQCa4DVzz8x2EnV2L4jZeHqdd1a0d0MeAi8FvLUlhAWM/8qT1QwaqF45PTDM1G
fLcVgokPelfChSbN88BCcegACwsPnfXmz8Z9NBz0LpDkVbiR+TnW3dmPBIkzvIFARhwQoJVLK1zs
LQkKWbDjh8V0w5HfdRJE2fFSqUt9rT7i1Ri+JzWSHCfG8MP9soDbVkUCX32eciCjaMbTMf5jF4Fo
cGWWieYzGnpYgRE/fBqFtnFpj6sBVhXYdsq2Eekr3U2ef5u8hsV1tBbKlKI76w0lhd5SXwONcQzf
3VOOV6LEXYttKj+0JB0mbrAY/IDsBPvdG9Xi983LCnmaDpnq5Q9tXSJoc/1uJmaoV+0rClVsxjPm
S//0+A9ais61RlAFYmM+ir9FB6qz+W5nP+dDy735BbX1vs0rM3KXrsvTehFcJGvWhWEqxTMaf8xq
mQPRXg/mRVTZb6oOtQmemeVAPcHfGUp6/9O6FeMYLusFo0wbBGr6DEOqpdH7GfU4v7ADN9MZplvE
Y8yrvS9lPpCApsP8K1+P0PvFU+1sDMpl7nD7+DYRuH+8r6UfbB5R3HtaoHeMOiSWivDHreBAygD5
KCZ1lDYFft+Q+nqqzhe7JHK/IQUPWVllVL4TYM48nj8MeGXnTWKoXOzdIbUcxyI44NVVxoDe9Dpf
q8RXsktvay455sxW1EoCQa2x2xxOrsBO7FHCCkL5nAgvm8A7FaqGptLRHNRTwM2UEioI7E2E7xD5
3TiPV3z1/M/2rFo1Npa+2cpn2a5qbEStx1e1rivY5kQtu5fltEpV7KeUrSQuTj4znRozS4YU6YxU
P/jJmz8UfB6NC1A1ntNM8HU/bHjShHcUcf88ekAxenb59cVqQzM/vmGsGCAgv63e2RRi+nY9dtFC
7BVDqUoCy+fe9VjUlsxJz3Pj4SHyxDwPvInYWt5XaBndFY/tKW2ugKgzwPDUGRmPgHR/L4GxbqEG
Q3ygBstwBWhTZzLjuQjf6j392qKqpaB6tH2b9UpgIUa69Fp0A6mDnZvx8fBqU2YASdtpeGGFn4NK
nQpag3CtyhzBJ32ZGr6S/rIs7Hub/FCHxG3G7xNbO3KOQH7gm3B9MhfR4v2pc+sNa9kol1t1jYuf
sNhbhDdWV84qGYHceqPOVGZnoyqGcfkIyG1cnKRIsu3HX7tEexkh0lrTgx33BxL0/JuC0Um7FdpE
WeRGQIgMgxIeDnHvM5+8JNd1xqL1rdUegczyt5+CjQjkDHS2dxfNWltCW2BXKXP+oV7fYfHFgJh6
86+M09r446NdsZGN0vnApYwrdGVBQf1OF4NWUH29jfafTXBrqifKCWpW6/8Hz0gKjVRz8gP2shO1
p76STfZtoPNfkN02ORwvF/F/mupVViDqySqnnHDhaMdA2CyD2B3wGKo1HlqUG1Jes6ApRfQ8d8fe
cD7moz5hd19u64gfC60qQVqiPNcrY6dZhaHRowfrYcLhgC1WmLeNFbDOSRpQiiBiidXCo+ZlfFRn
xmDKeOqTqEGcM8TFaUevxteAsqIvKrFmjHlArSlZg/T35wA+N41/v5dJdINj9OeqwmJaC5nU/2e6
QsLHwQN/qnGWRlHgsNWizBrN+OSSeXD/yRLWVRpkU5BFXVF+y9fR4rBUhQj2VtvLsmaL1s3JZRft
emF0PnNb8Do03ZYn6c9uWewNPUqm3hVqD9x2hvcl98Erc8gUy4FnjXTg19CdbX4uCy/LHkH6cfYv
BUPYnC7dpIEQdYrhtJGQBcy4cKz6JN2iwN1VG/N3hLtsKRw+U+vzG+azON/XUjIrBS2xV882LY4a
RH7imsw0H/ww+xukRPnqH18LToH6i6FmxzKdcWZebf0IAgeYUkyrqY6AWkDnzw0dLo/qVyIwFbtf
MzKrQmLDVpMysoOpKMnO3oHXx6ioUv3UVW/Wd3D+NvlLr27in9OwNmNHGZjBmrKIUPIfDHiUjst8
hJv6kzFwDSG5VfnQlbF31v95HEuoOAoptHG0tSL9bYTgomKO5jhY5P8ZWu/fDXDP/VrgU5IuPT0d
KhAXWxP80h67ctjPbnSIlO0j8jXYd5gf4hJ4C19E2Z5UZNn288mqFUMeBLerIyXVlRhl4wrK3wt/
JKK8XhaxQ6frtv13tfHdjFuQPB/CBxuUKYgdVmL025LyXd56RE+mtS5zBsXR2IyHAnVGQljNjtj3
HGhZAG+ds9uN8MuIkxgSYdrly0S2R7A7crVtcPlV1EAkFcyJV4DA3IoSpzFb8k4e0OpGRbLncl0K
1dKuExkU56KjBFj1pglWpXF5T4OO+wy13jUn4jno6GXbNEVAsQXX7E7ZiHtTB1ZWaqnGAEZ7b/EX
isyyXt9ORAZJ8z9IGkjoZ4zUuYDTlFDaJisi5RZf3d7ppSG1Yk64aWqDLI+2rrUKaWRMGAjtzStZ
PHE7wXlM8mz87RQOEN1eh1ZIWMDiIo6C1Prs7MT1kWjKHhJocF97j0pPad0zBzxXw9x7G7ZP114p
DePSnc8G/fiehKsegY7cP+AtrXgg5aNS51/rZpETv0u1TuZ77qWLoan8z8JcwwDUb5eXRU+md98K
inQ6pO5EtG8U8KOpsXIl92UL3nz6NhDqkfyI7tUkLAJeK83n7YPY1UNrnCD55UZIF0cjcCBjQa+X
inqCPhyNv7Y+GkRU02XC0+IQQ2bBUeV6GLrp7lgyUiOnIma25PqZw9QJHwtmPok3EQI8RqLhX1rY
fY2bHtFvTQobFfhOglRyyqZp43n/bhtdeHpWCajLxC37YkagZUg/eV/iZ8F+7B0hAYLAnCmGzWIL
A6/NgoNKY/bJv3xTtTi7qHS0xbG1QKf5i9oU+gJL2u8S1CSzZ7aiuouEOjmvd8No+oW2s9wLRSCw
Mf0hVqwhOWK9FqicsyUmd5rP+Q/DEkSgVR+AjVjHQoc/5gP4B1UG6/9fTo7EoxTFAzd8bz8pr2Yz
RF1pUV8dpxUbAwxpFUPAf99JRqI8Ko9S9mbvnCLC62gu1RoeCKtz5VqmsuDmmBbKCHHLM8uDKLjo
v6zT3QDFoFypZHNA91ru1sqOw349gA2m9XeJ6tCvmXh6X55Gml/+Z36uPU25RUqaKtWNA4TM7oLJ
+/GpaZ3Sw7EBLoaBgfgWq/dr5qM51wflxoc0qpZML/YN+vKiYPl3tfASJgibK2u2TR8BYFvuZsE2
C4gimhAliARXY2Yh92mV5IV8KjydgC4Em5h1TPWqzTFhE+fvZOo2aX5OUoabqXJFdJz1YSbe+CHz
kww7WWA4+gxw/Goecqjrrscgh6XpVUtG/dWj9W+x1QjnNcCDzCPSPIL+DuTG76AXqYjhYEmUx0xh
u7Jvgr97VZUPW+YwfwtIQxSAN+m9b0nkiuG9q783p4akTqvwq9kee4rhk1IByjXMHqoDPPD8aJfi
kpJhFnJ6hDhD0XpehgOtYdpwKcE5fc93u+000KOrV7ufn1bPgGGX7Ckh+8GXBd9GpSwUaS8jIj4e
ixA1qjzchoRL0d0JdXfH6DqUAkK5scQJXKayLh3mJrntSjcDcpehtaKYHLWX3pejc4J6HlCG/BuH
zeZKdK2rlS21sa8Lh8wbwsaWV57c0O5LrKs4N6EU5jt6ujM4eaque7Bte8OLtoMgnbnYySQs/1nO
h7DBGQVyu3zLE3tUBbusQ+gzDlGkgIAbFgPn1uJYezXxmdqM3dQmzSsdImerUzhR+5QF1fUwD9en
9iRiN3+uCRuYpzadZeT6r5pmsdLhznc12c8yLV8uqhRdY8gyvyPChzhXf70NNnv2nPjhBq9s3mt0
7qAEu1iUMYVhZ0lX7ksDTOBl2MQ54FHLXDRSdx3UeMRNxDOkW4qNR5PapyxKmdIhrRrMW128gP2W
bD7yaefh4en3p9fbIzgs2DBFBFgqysjzwXOgFGcoK2gLCIhSS1X5Qs2Fho4bwTB0YbG7AZ2O/ruK
K6yJCqoSnqLWIUJcOTLuS54fFpu/jbmRcKQGiFTtXuvwjxgfl913z5rkLbM+lSpFfEB6MAdmSHj2
gQRp8v6zwX9wH3sYndgEZy4YY7sbLc7zpk1UMEQQjO4OCUG6NkQRoFODeu4DyjpJlvK/qcCPVsnK
dT8hxRot2VNI1AS8t/wRnAOr+aGzCwLDPCPLwDxPGuHeMmFfI2W3JHDWP/8nKXYAwGE6fcIKuNBn
rbtAdjiBuF9Zr7TY+GYxW0A/cEgD8hP/XriVgW07VkloloTbCGaJsDz6VfFfTSVYHTHHR6/sQRBv
25lVci8W6k0jzbYAZrcuvrn+Ti+byLCblabCFI+t+HnbaXRBNvC7LfQkE8z9hM4yk40jU3oqTIgg
l38t5POxl2xpPZlw/aL4YbwfYGRKrujfL9mcIbHbiYuj2q7toesWilL0E08V1eMnSB76uWBvhHT+
dk4/xowWQoLWrK+vyYcVPQnO3XuFs6I18EmxGZS1OROCwe6YR1F2DRfe7ixg29KLvWAIk92ZH9Rr
MpFKsQ9XbYtgQUt7+AxafYmzQ9gTsPK7YDkpDRoevXjVs0pdT6i7SmtCd6Yk9+CkJP+5FlTVSNUs
u0YsXe9cc7A64+Jj1SNYXaEe19zcFAZZU9KLznOSq1GIqpdXsWu5t5WvbocPIhoWm2EHh7TwAbVJ
xIWOs3KgnEK+/1HWWIzhDYFzqdDUVSIOfQjd9lXMmQPvdocJ4d/fL9ZoUXexCRosPfrBlyH+B3+g
cVLEZjddfwSLEYVXXTlb3JmE0zdppXa/hQ0FVGPefmYlcs0W2r5lRsBJF7DoqdL9Tpl84Qim1GQG
k9LwUXrzXFjHt/vai27D6xK/2CCT0IiteGtpKzer80zRZ0voIdDgHTJKpvuPO0aWftVTRO4C+KvL
/I2BKjQQMJSvTAJtZ+NQje4YqE6m9HkcZhobSmF9/7RYl6Hi+3qQy1jh7sjsrrL2MS3DHiNlgrb2
au1wPT1QTD6RgCYN8xjbJea7qoRMFSxFbBSBqZ+ARiDGhCjva6UVsqKPj8/1WQBW55cNPVr8IzA8
zpuDDZc8SPh0DRsToZtVTpWlo4SpIl4DZFiGdIDNYgk02JLBDyn1MZjKDTq2Ax5GDduBrJ9yT/fv
xYfF5OzmDKT2GhAoCejWnA/2nFwqVVq7eyAayR1V2g6/MrPByRkkDWvRBrukniO+k8qQxe8DKM43
Ug0vBVZtF4KcC6alAXk6JPvilsaC8qyllfwX9CYK9Una+OgshQA3AQhwtSEVEHwJGhQpUIsyQceY
brUtcWym5HvEW3lKxjYG83hFwgqG6yGHQS9vorVGN81FQ59KAnre1DWJm4lp5EweWqwKfIs068fP
mV61BezyJi85UtVZkTmj14p8igaGuKR9gENgtl1aAkyKGBbl6GNJVozpMworBXeJZszqcQ3GOt6z
vNMmt/dPMub/gJUM8uHUhJGrJTMsqwuFpuxcr9ooBVvljHFm6JW/baBcmVlS3pc0gD4gI9qcbzGj
JTCdG3BfKAxMyhOwTApbehxg9a040Bm7HQLZScj4fapg1YRf6S80OW1H2PwU1wp1oMumV9Lg3oVA
fH6ooTEs5Wg2iCAGsZbUNHbwuq3ZFXOp3vb33tKCHvfH+SFyUBb77hXSx3Tbgnx7b6ScIYr5t786
YHnP5xmJeqmcl/k7p1o2hCmrUtBC2lCrymSxxmBSJAbFaJ4GvVpwFlWwlGvZExZGq6ov+c66p7xc
soQLJ1xdVhgQf/p+KUBbh/ZGYLaRczA7hdxrjts1gkcomfP7kUfqXR+WmDuqbqds4h4W1ORlL04q
Ah4addi+QUtySXftbYzEY+OgW7Hb2IWrz8/iVseBLxvwOBkiX7vj1zigPQLH16kMIdHR0ieHNpIT
VyNmOeCToXeg4BxnHegJ+vEx9BTp29092STSrZnGwAmYk/MqrknvRKdM8zq1mr1AV4qHLpjz71qU
TeNi0REWEFdRZnDcTJdxaYBjq7/4r9Jwll51DvXWOl16S5qOhgo8x1fnHKEnq6tYAKohttLAtpAF
8aFB2nGa9d/O3/oU6ywz5Ns3r5sQ1Fa0HpGeo8QVhOKmwdY2L6duKyMlwEWIvb7geiq+tbUQAKGm
d2ViT9Sl2/U3aOIqumyzl5oJg1Abj5895PB3wY2yvyUzQxlcPNkqGCFlsz5T2XYu2KaKIfP+oUsS
7n0nM1I18WGUJS/5o/g10mLNUv9idrqhgwk+xJbEY3IO9SSZIDhtyR19ncjSqZBhKuHm3VOkYDWP
7qfz72XGhChjm3ptLqVOowNYwTDFzFbwRAepJjD1rLVKsUd0bFeCWQjvB95TFV/BejjvU7rTtwXw
LmKUY6TlcrAQvxqQpBVx1I47V+cYgRUCeSBfUKi+mvOZOsVUSNziBjw30yPJJzscmBRYhAx9WnFU
YVBy92L8d0g5XjKIMwXwQPZMluYsEXdJTam+6ViLBMGqacwOtYtu+BIoF4IQx4wsOmq98KEOWVK6
xbYl3oJ2JyZvq4KGUxHW8TdPEs4by9WhGsrIlKK5udn5RVk8Uw+vbRUpJawHhZMIq+yiMwS31fis
kUDXE5nvoe2r8YcbCslTYvI6185pBFLyrAaJnAKbraQ/hFS+/eQOCRHyqVWqjTEPXApy8gx4ggMS
vYlfrMT8mJ7edBaR1BInap354eMKWkUuNZL0dHUc02aFq5f3YlV8XNlaWDUUdjydqEhO2Lg+7VI9
gYD+n+kBxuCBqf5HN8+ItIO3jSE7I6MOzBja4szPawroNkZdgxC7BupkIGTOC+RHkGGiOetA4ZrO
ATAxxoMTVucrORSBf7mj5GJA7t1yiCWdqkSJziVUycRxHPBBESMX/ztYDQR3u5liiStwappVwMh5
DlzF1hYOwM98m4GQh5T64X2n/juAw67zVsh9wenF8LToOl6578L7FJgfQYJHSnBwg60gKYERlIaq
zWo0NCVYpysVy4Z39/XUChQWFUXJt24Xr4FkjqsfSvwC0ADbZOpjEjLcA48Ieo1GxzmZwsBX7rGi
2ygCUce78GtwcBjF6PjNhe+z0lPuQ5i8ITWKxjI4zjOFZ0W6R31jLvN1FBz+jsq1dzSxeBoDJrGq
usikc9xmHN8NWgi8iWELOquzB7VZqErZdnjF2KYoGVV5d4G6l5wReFpl0JWYq5FljNvPPz8RIyQi
xuVDo8U2nwuBYythG10kMtffv7x//U28iFSpmTbYGW7KUOP+P8Si1pJeC7Jj3y0wDkoTcHnQfFkG
XDHhmsPqBr6gMTQ4/xaK4T6o9AZTdkPa87/vtFN1g6U0kAfoHWwuyzjLl/VLD9OTIehKVTMajMKb
2VwC4fipwIZfwEyTq2OSixE6Iik7Kncr8RIT5g+EAZk21zAOAmJquCB4LlrCuKY6paRtxWCluiKr
i0YHF5gbjrvmei3C1msAC2oyzKtxQCyZ0UAjLJnJlZSn0EwPQHSfdM/yJ+XFUfziXJ5UIhNTyZg+
dJCffPXa21p7ytFRdpQVqyQofX41M510WiAUP1uO0h1qZMF9gPzZNvZZcThyEBPQPnrUHZpuCz2n
+dsEcVoKrJc74T0dAZfyVBrBD+7mIHt5/CNijfyfXe8ys20w8ALMhesG1FwarT6YG2aXAbQdUSFo
dqJvHAFPTc54d15EILn+ZYedKKUHevuAvnMlsz86jsCDWXVrkgPKSfDtDn4oGbJrp1gS7o01I8H0
AUubEpptcM1t+anUtwwavuw8SO60sbWgdIUfFrHo6cljPXBpHynGU4T9z5lxGw6D/G67aQIPmZE8
hpwZ4bfk+QrOoOpM0BSP0CatD1Scq4S5Ex4Tdw9zcs+buHwmOfE9w5v+gthIPOujEdIvzwWTScqv
gXh/fMQEEKA2j/WN0fxpOmfGZ5T3Gmvg8fFcUkIPoy49+Tra+PY9qciqZpvqfB2qiQvH6QalkrNX
bpZPfBAqOT0ly04cWM4vu6k79rnepaNJ9Rw/qWEyJ9qbGUM3BkqepXO35Tk7O1WED6AkYL2WAZqd
cDAEsyLa01I2ZwmLx6u3eydMkV3+Jqnefcz+ff6MTSiv4zG9RNu5yOFWA0OT06RGqcenbPB5Ibxc
w8/HV0HNl/DW4RcdQm5aLx+JCwtCM9rY07mo8I7nTAb2FUJXFxSblNr7QLgqvH9K6D0R8SbFZjMG
j7u3mZsK7y9Pvl+c16tPzU+vAK5lR2bFq8okEnrk155y4akmv1m7N4YhoISqkr0wlhVQzL5LJQNj
suC0hU7MYSjiEDg8RMBh3WxDn6rpXzONiXz2LG0NuwEvYNbnaFEjQ3tHu7qIOrTOI0Vdj3A6cj8M
tzovraITJuljQWLxnRx7M385F6/TupiVuaIx+KGUT8ivr4OGSOeql6gjmumBSlpYi92eaE6+BL0y
HJxq1AcC5KkF/LH2jJZ7CJeaa5xzhd+nXgvW7Ap8D1nMLWpM85xJloDgs6sldFcaoac20zuAZ5Kg
OMDkMETyJq5P9WEdENaEDd5ke/+ZWUO5jBjhjGH/GzHvodZ8Ny5nt0fipvY6ygIwIy/tz4y5luE+
JSr/UvrR9inP54x9mofomv91rkYLl9zRzG0FJc24TT73OsN+AJKMP+2enTYfkbapuI4eawWvOYl2
Jdv9R+/swDG4fzS9jbnLq7Yy0mjKfOry8kdBozY5hsEOceChuXYBb3+O1fskOpTIEsZTip/juYqn
wIP8cFKgFQfb5QQmKB5LagyPprFfPKOtXP9Vajcu0VxijG8W1OJq1A54tUjBWqDaNLyZ78QtAwAo
BzcNlc+WqBdoxmo+706TOJviVuxAt/7G4v0vA6QXI8+5o7X7blZOXvRiOB00DAIDjIvu8YLTyC85
EP0W7UOCyMVnDF9LQqBV/V8I6KbK1mkl57zrVbCfPc9Mf/cIZmdGMGikiEhIGigTPwBw9sLuDzEq
PCj7Q9mZoPaPYj/0bEzvNFxvfTIpd1mmaBJyuK4r5lryEFVoCe6kjwXWmgWVXVndl5SqHN5ut+Z+
EHoer8QIbmdXX+YCtCh5GCD7U0CcO6I2LNAZWySHeryfX14TFp052RT76SBnplmmEXw1fvgqtdt5
ziZCU+Fe/dECkSeQM/e0me3Hy2N1G0/leiUKkxazP9h3OeXEgxHe0dha7Bh34hlKhEv7bMs/DyPV
fO1GQDDuZXhyH8jWWPTjoaSedlFjZMAkoplgIyj47RlOvAWMIfzuZmMidZ6Xxbrd+8AfdckT6fav
kL/TOkjPz+SagwcB407a262HbO9rYAca5Ifvb0b9kBdz89eWdD0Yg5PTBM81PJk3jhyGXcXureK2
rLqkFE7IFFaqBnlrYnjj/6/ylSnGw8acIVJ6B1Bnx/gIivb38m+6WjpNbs+E1LmWw4lDSd8osbeD
y2qFOoQnP/jcIGxWmoAOZdGLxuK1lNt+/Fej9PPbcE61xwc+2Ihz7pV3Q44/cgjwibHN3IQGVm/x
G1OYerM6pP8fenX2eenLKn5UVFKRUlw0OrCm/YLSXvsOzhmqF2E0z976UMGAQwu8S2KnoRarPPft
rOO3aEYe38GIqUG4RvzuHA5sKRM1mDpKh9GylwBnDXu3rDyEMj0B9Z19cCY99dDe2lxRPKgB8btO
KCoeHtTiYNNa//VhrhT9oHxVgy8vC8cUSH+5ftaZn5Fgfkd6xXbRTAMVL/fTPiDXB5LxkDScKQKC
8ug+nVwtRG/f78DqEb/61Gp5JNvat4vuFMtEZYPiLFXUWe2qVWq00BPLygE4QROyfC8T+m2ENBy5
R12YpuUAlyrym+AqeLazRIoNCY3XJxUbGe5A6m2u0QfuR8qN+8bereT6IfYvUpcMi2/OpXqFVbht
vaS+V91tnUvoSazRDbBRS6i0j0/M5I1yWfWzdGuB5MQ41Klq1QfIzYR5/vW8vELAggteXxb6R4Bc
o0YVM/XrWbEJUb2LbyDA9aJ4GIvlDcBPXpc7rBK85L+xiQWXnVMMzRCh+EXXM0nlFBNp/TCgyHgR
4ccYvAwStjVw+bvbsKOKtUOifLJJJiiTNF/lRHl0Q4PCwA+AETdxZSp0MrhFYNWOlGtHZSMJIhGA
SPp35OHw1ICokL9e4T2bWDdA907h87n6j4K9JSOgPGPtjGqpvdNcZqcfp8JTOp7CRksxH1XsEQHA
ka/AH5/3YwPZmdd1FSs/cfdUkt05Nie2PARC4bXqWab3QU/SCInfMVmlqrUUMK4kR9jsu5C9xKEq
FXSwuYF4y73Zk/KB+3BHHDiR16TycZnfnQ6mAa0eJs3BMU/kvEL/sMEItHOE1akl+9eNPWEdIoH5
5l3FNhxXLCUYd2ZZ3ELdjlQepgu9UmckNxti6UA8MW5fJO1etwZlV4LM7dV3Ec6MhKaXWthKEhGb
sfmhrkXc5Y/g3YisQPJW8sXayAe5w05RPXHvC3M7qhxMdFtTZNJI0/QiMacEgopOkX5l0z2lWEgB
V1qpbZ5UmHaT7GVGgKDh5vfzXCUIWRm+GdQ+6vnZgMzmmF8vK42/pvNfkG9SvQwPKzbd+rv7ED1T
T0DQbMiy/H4ssI1ZeTWxn1T56J5gqgTUsvuTKi2VDyUHt9KQlNNUbho6D0MXnbXopFGXsRmWx3Bg
6gY86QPQ3untPA1ra0Kk+VH6fRycCRFz8mxrU800b/S9aHXC/SPEzCbqs+l1HyGysvQmCpSb5elb
Zk38Bh7ZN+t/ZtBHKvZJqck5SAUyPzAay5UYBeuFGKwsFm63FMz8gVK6eBUTGAGjqENw2X//XqOQ
zeaB82LGQahtLKY7wcdrln0FpGihE0mseVZjN5XOEepNpTwpI3l7gFgnjlJCX+rBZxvEBUTzSkYX
zpKRvUaADHn6yWWpgE1tJxCgk2Y/B0ErBRyLXy6rd0149ANXv2sneGoionn93oKZ3ZJm63DTnelx
M9x06R39XweUYXZGSnTD96iSiEm2fJ3xfGOgk6wvSiKXhUcsKNoEiXo9RJxB8WjKGJjfADQRslJk
xQQ3WY6d4zV4MuBKdD8MM4r1WUkXfGOp2vtc7aAW7jC141AxG9DjMXod9uLDP6mpluZYVt08Soai
YAAaMyKfjU1H3On9IPV0Q2COnwFWan78GnerWk8FKFgHuce6KAkgoT/yOPfkkvb/b0aeBZrkDRaV
2qN1zNbnIbwK2V1gSINBjmjBl84KdCTZD6ECmoc+OPFZw03UGgy/zTafWWIkSJFvHwg8TbEA3XrX
kYxb2de4obzdjZQize3Kl0PLgFx4aUOxmpJ77xZrzen6IQjzfeYcwzlvBO2K2x1Nye/bHpOSV9YK
VBlzMxO8A/cz0Hq2/6B9HB5gTa41FuQIaLGOsfdLzdyWJYpbnizuG8A65ABLpi7mETIo4nK31/V9
6laZOXBvVwGN5gLnYu/QRq6CrjKr3rC3p4/o2qEUrg5U4Q3cu5i5KMgY5LQyAnePkRYkNz0Z65Zi
86WlS7wdw2TG8ZXUfcuciZolAYfhhCjWON7/8H7204S5oqmDzx8tV7bq81E1G5pKm/NX3bX/LiQs
Yqvoauy8HXIlFkFEJnm4gjsbsCPf7+0g+IszciBf2Oi2AazwBybxNBper6l7yRiy369YTlXvkIs+
LiFd0I1zfNZnguae1TyXZxYmSrfwoqGCev7F2bJ1xT5tGmcgo+LGFcyWMCwNnnTyfy6aW4KYfzAk
3wurfBw3FTK81oWm7I4p9T73VUrmGoe6mOWscWy5vNzidCxGKEpYiwNR7M+D2i65b02JvMDTpwpe
VuJYyaItOy4B25EwpRi/mpnY+N/nOCv/hMp/H2BOau8vNf3eN5IPbv7e+VrbCQc9BcYsP62ueTKH
KKWMBgqkWKBzx5pxQvgAwjM1Q5u2au+mQcWThF0+WEv+G7zMyGhs/RDv7lxJ9N5ja74p4bzOILGr
Th774Usx8++UeJTHv32L0NvJZT7GPnnYdVyUjxnSI3vzvDj31kVyu1UFFUSHg7dEGA7zxmnqze+2
3YqY/r/P3F9gDsLu5c+pCeUD3CK//3JNVAq9hhkXi0bU+sbBPwuexr6DQjFl9e/9l8z2sFmYjD7h
UeoqueLJFK/Ob6Kn5xQSVu05JjcRLaubzvtqzk96TaATdN6nCWAOvClFWJqThurfLqBYUnQLMxy0
Y1jOv4OUqDGJ13sYM4E/lWqfYxm13dqXdgbi3rt+ktNRdKKySfjxlCuMyxam7+OzH1Ap1fFmyUVh
XORCDQJn+hlxpy4WqrFyCv/lrcl9BVBtQ6OmQhamkl1nML8wTIMd58Ehw7E1tR9mEjep/0TWPGXi
mj6SsBeIKREGP4ACYrJU3YCNy6n3oBA6BbSDbGeLNiFkKqHjihVekMYwio+pViXeDJA+4B/Zgbe1
liDlnefTVZ4xbdMmckqFVIjb53rMlwR9IE+w8WAWfwlLeJpfz0wBRUQORqCVWd4OykUzREHWtabL
2eCCRnPpvna6166FRpcmrLJJnmL9xjsiJI13SWL+Z4mcbg53/ScsRmo0xGfb1nyWR0aLKrdb5djC
P5K5LRrOp9MAQuQh9JcQQMe2I38ZaIxB0Sw0nFMHgOxSE4IDz7MXWJBSrQVRNufTrCI4lpVFpDQ8
HblmMZ6nE9JCS4R37KiRxFas0yazaRUO8MCm8KX9/CD+3R5qax4kNKb6pAfMDnjOzvJjThixE9jk
Pj/pnkR3bap6svaH+9hOI1wxiYLsUIvcQAHjGWrgMM9FZr7rFNIrPCP9p+k1I94v7N2IZp3LdDsH
Jlowy9sAxjViA7c6Un6kfDXk8L3NLwh88v464Yub4lMEBDdu3Yf7q3ulMb7x5hkB5Kk0J899lwD7
y31saNwU6Ei0fYijdiFXTR7U1eiKi3Pc8inCXMqSGAo8ggp/W5iwR4WVkdKR7ZdnzP/KGzf6PNUv
M7+wR+FkEEqRb+TxcW3j0uiXBO3nQg9So/vfKCQt5YjgOajXtxgfdzfZy8a6WOOB/oq/o2zLLW/P
A3Ne/169GWW5VYTZdOLYfG3AoNSrky8xiuq0CnlcBkKLGHyRwMmAL4KKZbU23M96UhtLq1zkZTjw
MJWlJMuhZ+CG0UfAcXPoVCAuc0aTYV9R7usOUgI8AYGG2Re2SyyLRjEKrtdhYWL7XkOBbaIrbQ51
Vj8Wa4FSN1lOAIOJRvvZf1pKoRsSuufemOViugnSA2aMTpuVN6FzNOFIHtxpAwlQQqvVIyaZ8xj6
FikG5pdsR3rizQRPn4JdRhBgLuK1aLCPg46ODww8K7kms9x5sUvAYVi6nHa/ndCBuFZhhcPca1Vs
uPFdbVSBLrKqLZt4PDZZ9cUFQsS8hwBnNbaUVcm/iz79W4bCtAB6xh6Er2Zrf+DPjkf1nYHHFjI7
SRT6MHYe4GaA6DG+kp+o2MM9wKKUcQUM14ve5+tqKTrMRVV7xZ7+QgyJ8qWQO3d5W1ejxaHCFtQp
lEXQdfZ14R4MtVUBY9gkaBTztbxFymrkFYYU6wKXqBdqEmHbQc2SbuAVoKwapn6Gd2Ai/t36L6Nr
+/IU4Nsg8DRL9HNKCzdj4iWi4RazpFG4BBRrhtIbER+mIYU2+AVokxxRGArSoQqteBFJKtlTdSPo
T0LN9mfs8zLxgmX5KwOQDknJfeS7Ggz5uLhO8OnuHWLsvbjlRUx2ANugPrCyNrq1rPCVZHZtDPr/
oXSGg2ih/h8WfYBabYv9jZ9+eXKvGUBa+oZ6DhU9ekYS2pkeE4vczYT03WLFG/WLg+D556na3CsR
56D1Zlw6DGCEudzFuSlEYPYBkXeN1PKCGw8EyL+JqTaJKo5PFlnK1wMU8p1FPP2MMqkXTdB8Zd/+
IxgXS9cZwthiHWGPYkE9zQ78soKDRhzE0e+ytRJOWw8dkVaiO2w2ASCm5Tyngap0TUY1I3uWXvm0
6bYtdkt6Ce0cZBmNcpQvzXnCzGSjrnnI3jwpptekuLD3UQUxezx4z3dz0OrC8qn0Q/tg47do4LtQ
QFj5yvy+EwxZwzOf5YOlIyyJ67ZSEYNTjmG9FWRfOme+Q2KkfKFuc+yXSNQQJyZJO9oXoRmCqX6A
iKmiHKgrKJvRlIzDSTd2GSbfnB+aOpwGPju82H1Oe9sYvTZvI79yBT6MTr3RdVWBnVdgPOVe3+xQ
Da5n3v5ah1QRjB+VFYXh+QPGfLZAFRWROlVGju2gl9sMiAV84HQtFaqcCw7yZ1P8MwJLLnkZCeLb
R0s4udBCpGxYq/QTc+AYPqAnw79G3TBVY3AWLfupTy6JeLerqWp7P8akCEkH8uDSCZR5egvbQYpb
SiIexx98PCWrNm+hd6BSzlvh53VgPLfjAuw9SDfUdNnXZGDFdH1zwJeGKL9K+EbFlqRBJQCzsyTA
HWwgu2+4NX3rKsEkoUxRH0RAAfmBaYntoCH7vtm3p7YHEOhMSYd5U5kV8KN/51f0Gj5SPecXuOyF
OTdXwyl2WN6aEVhif1fqF+p9xLXwFxjkVOqBwWGQQOXAoWMD0RpF858jKOu9+TWPmDJoAh3znj61
38K5M7FhPt2o6AlqSTVm9UvsZrgiTnDAXWvoNNJuI5/03+3U85XMcvNrgxJJ2EktZ4nKTwSScTFd
wnBtzSgvAjJunfMYreTva2N8uqg9RsZ/6XDYZyt3gmO+ykp1Z6B2JBhxisGqq77+5ZnmOPpVJy1U
D22gDNZpiGGP8vYkWxSt3Lo3wS52wbPzCcdU69ncdJ19B1QtjKbHUHoSf0GHeUJgMA4K2yKg4Qul
ocoWOW6bsIHXTBQ+P5sBzKFE24k1qnMQ5IV2bH3/+95nY4iA6728YnOJzMJzoTEz7UJGljEyXJOT
2du2BjJN+DS+fUB6W1WZWe7kO+NzrVuWvsYsbILIN3JND0u3GTv0+wo2O0hvROK0BgFgjJ5XJoHq
AZEB3akGa/b5zL9026DgeW3+dl7sMypFtwNEYFXvUy2MbDFtSUURPUl7rYmuizaTasadrfvp4vok
/5VamdIv3mGfx0Z9LE8hoUvvU6YZCrtirr3KLrsnkb9HEKl0eAouu9Cy/MZs0XxYojT4kzEkzdJ9
cLeLihMnQBrW2ZwwkESHkyVJRq1hREieFPAsAm4hhJeCdyX9+FtTe5DgmhwC/NHWkPOdciSNjrWN
iYR340bkJ9COimtUEtLagHIcjS0vNjbkrsO2qISGBXS7WwNYNIxpb4g8YapEe2QOWkgcdw4ti7P1
crBY/EOKjt4SepSpaVxrVkU2/uqU5P0IJcQE0GrECoAGeqcdkiMir/KavhsdGbSKScCRaxI44pr+
gcIutlC/TkxQs7Hwm8Fzx97kK7SCEUGc3Xuyuwd71RiivlJd6jDyeYNEWbCKxcFkgUMpq3wv7W+w
dBFubUt+cWmZNLOA+bb60d93kslPNxW2b6KyDLv74wGdi/kx3IdRiaaWs+KH+v0qS6mfAwGq4hV/
G9w40d/52/VvG87wJP7uVScEZfRByon1ghTpJJ/0wrTMOYS3pkyA5odjsPao3Jh0g4DaGvxuoAJm
unEM0uRJklh29nB3hXwJcjdzAuCNZ4iG/ZunchW6N7IwN0Vb4SGpsWFBx2MGNur70a1d3aqO/VfR
NN3aNfSYw610Jt73JnDVChQEaj2ZhsUlMTRIg18IsWiZYAVLSHkMhLErwR2ApOUHZaegDcvkcyLp
qebD3e5XGlTRaVm7YH9kCaJZ8BUt1GzXH6CQX+Y4XMTHLzX7GmEw2nLnMDi89j8sVHGQ+A0X7o3G
e4f5PkC+hENM4Z/Inq8MuGQV6DyuiUVYYT9VGibSytSmsqwL4g73k4tB8DSw7IkKbrpg/n0y2qTo
XJV+sIhUl2sdAhzP8ZW6L0e5uKczpKqyXSDvfeq/EM1avJalnU/8GI5Qdsi8Q7kMKM9Jywd81S+W
zLZzU1d49kzx7CJUrqY6CVBs4vC4dcyaZLaqsInOEMs0COdYhUNunOYr0Eyhv26yYM6SqNLKiZUg
CzmBAjchz6GchB+yjsWT7zX4p1uHNxOUM24lzLJnPp3Q21uSA/sL3vJ06JdEhzzhmqAMycOqowGl
1qtnsPrdxhwYFd/1Ywwq0zcbv3o7Df494jIJLzizjmN1SWcdSxoLcTlCjv+UYDw7KTlu36hg3j2P
LctlhIOWezoCKgefmbDMKBm/fxlH41GOoOPlUwvoK/geGKy3wfT9rRq+tSvYy2Mc6J6+lPSAkwj8
lp7qg9sYR/pH2FGuB3kKSVha6p7jBHuq4KWCgVDij3TzrRv8MM7BmH7gxLZnEJ/dMC76BCckESnD
/Bg032USntPpcqeZHi0cOa83BgwGuB7HwF3qAlFs/XHidAx29f6LgGaYeduH6/nl9C3uAElJyZuR
s2TspTDRVFl04cEmetol1gRNMkWz++p5J1Bu2h6eAv+sG4Ow7cUzPA10yRVrFEsJNQ19OWJqCRln
mkC82NVjaKzjARA5yt6RyP1TaYb4UW/m6OgRimUNPqg2v3x0Zv+zya5Esm2FHnuS0S9yDMOOcSG6
EVvmO5kBJi44zgtWZvujg9gnINsi6vvx0+6CLNRLPgHbXkoCBgTSPV3gipkZpu+zLBjI+aJXjAWk
VMv6umwr7hP3v0VbWtqtS/615ey5zIDYLlY/+VXViG0GS3QSrkCVbtu67QfuD1tO8uJP62Mgv7/e
bBePJH55r4Ch3wXAVNpXmaQUOKjNl73X5GLpEDTDS6zpTLiKfI+3+6T1aw+9i3TT3qDU9HljCXep
njlSvG508KGcxqviKKmfF58CBSarbBuNIRZJz5gUu1Fh0uSTojVZVx4UEtGUdBKd4kH+PyMn73/T
zCtTw8NWftiVIQMtNOZeen+k/SmuVXJEZRPQR98w7WHLc/EJ+LGLLWt25fTSWgZA/n762YAiFZQi
/YX8o0YTxPySr/Yp0iK/nOnnNtZCrgr73UjtU4ju4Q4x+t/wOPGJM9Dhf2AGB/s1bL7jjCgXrD01
qeVmQiSuQvcozcAa/QqYQje8xQBz0L6m1/d34PB++z906uJq/M607cKawt6IQXgQp0Bf1Z6ImZZs
GQE4TGIrVZ4sAiuwiDgNu4BS+G0dJna+xf2IFn3fH1uIboOVXDOqBGsgQYD+GkIEjRX4G25gZr4P
rv+L/Zvw1u2GlejWGx+D7X+8cRoIrMVGeaMYRayVRsoA1EHXC+wNE0yOTTDkp20asB1/19BPjPvt
4SblJfvljnwxtm1JPqBKc3FiIWqmBcLb9AY7oJpb984qrbI1zgExaTkAz8lfFE7pV7ImI+DoHQHj
GwzjX/ujMRBSLpTEfqdS2uPugwvwT/jUuZbJF6Ixcm8mran3ePXJJl6ZeXm84/jkXZ45oiOG1R3y
VZ68hKjmi31ofbIYch5apdVUBvrm6Av6LYGmJGEpwZVR6rCoZH6s6jW89/FIFvmvCbewU/A+xp1s
gOsgE2LxFVU4qbaYC92FuYxR96lGrzb8aOul1NoUMOSMAqryYNgflUZG8f61ySJR5dy1KSZlUvU9
PpmcuXjlXb9NGNmi3iSRwJO3MFB1qX693wEFCT5tS6l/2gy74crdC74JWd0gbF9I1lpAXhvUAZlt
eIcKmREynefYUSiLmHZIh2YLUoUd/lWyRZ3CTSilzG88Soy4Aa6yUy8zc/lsqsZ6/35NjtwtnJn0
V5KN925gHiFMTZx3XwI+PX9piUV0bY4lfTg9jOuUO+pNxZ4JaN/x7Hwe5g9gmm1OwHEEbihKjvG/
E2vZOwuZqRQDOMjsITuvGAcLv6vWHeVrlcnV0mH4tzOq41hOIMtVivnbqRCg1+wMBkpNjxmN0lXW
iR9S5hRW6EW7ls9fDlaG1Syl0+LsVuNqaH2YrbogwErSajc7XA+QnxP4hxzZ/0nv6/7vW34hGB/g
8eWkWu08OIlKqCOQoqbQ5YqDjAjb3mNT/43jIhpipeer2lsrXkN9ZM8E1r2Z8OxLJYvM5PqBnIF1
OfrNiLrrWmD8CbzshZUq7XdwuLYORoIvLEOBVT5GEdFgjPEKHaWH4h+szxjRz+5ZXOIAmpmsLDzw
DSm2uTW0JanB9UdnvtGfmPDnvxk9F4iaJwUQfkEWhNTDR6SxKr16mWZ1oP1GgKhyqqs2xz/6/a6R
3yHVTl/VQ9t9M3s6f6oqdf/aAQZM7MVe/sUf0u0LUsGrgZrqYetJjcym4g5+5Y2W88Rk/MEg7gPi
4UWhOQwcF253kWtMcE3agZN33fZo7wCQnoS/UdeE6Bt2jXzYTpjB2mGLpTZ0r9UFPRmD1hL+aKFg
lq7y0b/no++GO3aD+gE4zeuPSlxEdrZsUycqjUQff7HMT2Ow1O8Z8XDwQQC4YWXNFGvKW+2YpKc4
6hfDQE4mr+6c0Kxqq43U+PPiwR4HDZoZdp094YXHMnrwOgEQ2IOLj58hvS6kDdBsEh4pG8I7w5Q5
w/K01XKCRHviF1wmzQGsqDXU8QMJEPafehQ3wdIfj/qtsB2K+7zewBWCj8uFY5oee8n1thathgPf
+6O0COz10rUfHPFJCKi7Nm1umjWs7s+wGZZeKwvbdtq8qNcSKPKYeklO72nYTgE4yXy8MH1qgER6
XkHazGKR/n5eGxThdUC3/Or84sOxg3XRYY9ofZWH+vhAZ2Dmb5cA2ndhbZ7RRMwNAoy4Vrl3fce+
jJ9maR0MWxMV17EKcAchAB07Lr/5eh1zwIucmd4tH2AJCdzl7Z+yh1vKcfATLIm62lGkTkiV9bxn
/9kfcHzkD+bsJHEDtAYtJByhuldAscAzkQdMULpT64mbkxUE36BUg0nj19gp9LL24HCxEImnOBoO
u5Tlv1+UHeE7mPNs2K0O+7G/URDzArip91tP8BcZKnhI6SFEh5ybOSrHunUCxezQtm3WoUJpoA/j
5a3z3r//hFZb2IT6Ht4xiExXuxPAXgxNxF6adJmlOqbcKCnKV7tDEvFNn/4pmlxNdeM4TywJbQIB
YGPBo6UfCcYzIl4YwH1/3qU91HOy00QY8oCrn+g87nGaXwEUxI3mKlkNjOy1STNyVmf4MIAJv/PF
znenuSzeWcD1yBXfhGzM9Btjr307Mr/vSE93mfccR/xRxT0Smn/OR5Qz3kfq8JZSs4ug5vrP8oBB
Es1K+2F0AlP/hBgKAuoiCaFuHxMMriyxfRQbQyxcqMsgviNR4208dSyEcMgbI80ZE73JGjmdbweo
HZO+ZI6Xj4ta1tsWafztGrq7j1adyl0KoKixvKQBJ2R7pbTcPXotQO5mQPnqNqlqTGMqehDMf1B0
vBsGQzEvs+0N2wWiZCxLG1DtO26TzkGbd+vaoDvGhqDrIEwYUOIO7U3R+I6evCZgVo51OE5Asfhj
CmCJy9hKhpKLMH4gBFl4d5fwCGXKCo7wYbIJJSKRVLAgIfYmA8YShjOCzufdWL0yTeYytAxrxbiT
fKr8eWakaGb2o2Rhm1UpGAPMKxJW0tf4BXuqO7/B6s+baYlVwEGeYaRq7b1vDHGy47AMsxWl8XN6
sZxqrWcniKbOkgUzf+oXkHbbYnu98zvFviuW4WjaKGbWSA7Yvw9x+4HlGCWlfuxTfOn/iiW09w7y
ZuBLbBzkYQE/amWD3+dnveWjEVBkxWyhoRjGC1w44anrXOmDFlT1PaFZsZFxp/cBa2INgHjzL1ov
89Aq4OwasetTPDhXs7RPa8bqorgPsh6l7GbEWeFXb2UYXlLSm3iX2oC7OTcx4DRJLQ6ZfCfzMe7u
HbNwT+XhjLyEdwbQxBGzD11tdye8O3HtkJprAjCARl9hP7jsmK5ZNkIduMdZHKe20hVr13owRez2
qsuI/Oh0M7gP336cQmJoFKb0TIxowtWR8vzk48CLXOVyfvMIWEHB3qDhaaRdhIU1DwbgOMXXyXMr
BrlSlHVPKLODAnI/SkWmaw3u336MP9pzg3ku5QoiwHFA463k9xkntNJBrnXgtNcBvaxiavNqwf3X
DrUXCDJB60Uu2smuo+PSNAkvJtkHkuRVreQUPywt2wePYHqpzYKio2eShH1Sh7muPpxUeFLILJw9
NAdZ7XQsLBeC6UfgwJdLUt8d10ejO5W4jXoCLYCOvZDiurBiosz3WD6pFSYRSoUN2VBsBH5qPmkw
DiZ6AjBem/69rLg5SDsriaicFcbZ0TMTUhLXMgzAFwkGnvM2PmYqC/vEeGCJ9igoKbXKv5FTB2xg
R2AQEdgzCC/AIpj/FkknHQby8rx1VRGTqEg1oitJdHVC8nZp9vbjtXbPPXtS7g17g7ZGv0XquBMs
ebqoPmwzs3x24eQFn1g3z/1OZrbozCSSuZNkZDGL5URcA+SPL1iNR7eu+p8IVIEmHuULzQaD5JRc
edFdvkSK/FKfA0may0M99r92XvDDgSumYMBFxWwOkKbR6C/od7infmas4bfEsdzovE5SUQcawTPU
8PGAp/Bw8/GHgWQh0E5fvQgDfUUsPOGjOAXuvFkx3FE5Ac1OidY4z+XNcXJ+X8me3QvyPIjwMVLP
hCdXKCjoATNNp838SnivPEr+NJkqEGJ7/bvezZPfiiLfrZcQ/UmHEuSoNw18UIqdcLJV+ZO6BKkR
O3f/G33zysp6wHYyerCx0y4W19S5e+nHF6Q9zgwKVLXVmW6TBlRHuy3kPMZtDudtaZVexl2Fxb+l
TkbQgjEpC821IoG/fS2baXEekKlMPyq/pokrZ+Uv1/6KjdvkOViVCJPiUizdp6T5EyJ8womCXYZ1
yg7J375muqi3VIJzfpLyZR42jfYKsbQy9ysUHqvvUYG4Ys+M+JbA4tLjY18F2+RrIspJCNtTqmzz
fHiKU52Rvt1WYAq17KQaMHYISHhs/0UODdZd/qJW0upYlOiPN6w3qaWFK82k9G+wftnIK45+aHzY
cPeQQMAiwMfjXTor2QAwUdJD5ZPPKXxcoYifbX+HiVf08l4xgvjMJEakYnvXScY80nuRGuq/ufag
t26Rgsg2Il9KgnZGBo6Mb6sjTWU86MQp4Z80Zi07EI2HKQ+lnhjnbcM4zQ0tSV/6W0y6U+BejbLQ
19nNkLtBh0L+2j4qNNEBLJro/kJdNczbYuqLa+TPOFIzKPNstML+5mk6hdZr0uNTKGeBSuee/fDg
a5CxIjuFMTRcwiXrp9w3uL6WFltw7ZCI8GJGGpc9PICB6eexwO+1Guu8Vt4Ou56hEqtqUTSZ+WCo
yACn+UtTpQFbalXSL8aJlR2q/FWOljO5bL7hQ+mKgF7UfwfkJkLAzUSf1oSUrvMJg0HNr+PYUyJo
g+iP0/I12SwThnTl6jyBYkbSd6+amKr9ihRbn+yLa9esSsI+nPycDmTO65GJD8TCmeAh8Mpj09Fo
jSd5A3QNPZjfTsBflBz9Lxybs2eT3DX1+qB5Mrw747kjhl/3Slv3grfdx6zj7aN7t5e2tQhUcRx7
R9sQ79oEdMkqW7tWv4+ykTOLZtD3iJ/c0DBa3mYwoA/Ux94eKZNGfDKdwvFYrzDJzdC5Cby4xcF7
9tEYiM6AJ/4aN7xuUGJvQhJ141bU2nZG5jvWBkI5DdcEy0r0NIelgzjwPp/a1oLr0PGk4akUFUCK
22ivJldNcJQXYkfH/kXm2j9TPAWWGhpi/lheJTbuNGqUCw9VACSdRUEzNrvCJFKKmtbgW88chfmq
d2ShvtD4KuJnPX4qeCECuvO1b/kBvBAUQ1FLmXoqNAejXy0UWpX+LVOvD+VLpOLYvVSD0BRqAYSd
tai2uRXOzhCiKw72UP6AgB6FHq+CYbm5LkIWuuABwT1iKTFf9hqv9c27PwoU3uqlOLe/ceYEBV/f
4tkalCXAcb1CX4ZYlSuicSbmmOIsZpm+BUPJ/x3VinIXXiAodUiw2CPTe8WSsSIfhxahVsge7zDd
jRJ8fxMCl69+vyBv3njGGe7REPYQVPhe2HgbMClzbByElHypHycyBV9u2aHgqpipulhwj026mpuq
fDzc7tuASxK8HX9DOGMqiMBVPgr529CtONYqO3Wv1mrE6LXhsBxoTfNQvZzEk+BifmtlpvX0WQi3
mnVYtGIooDOCrmVx2bDDtIfE46IOV7YTs+EicJskEOWpfUjoyeuthynkvc9i/eKiO4G7xl9Jo7WT
3U/GxJVSJoR2EKNu5zRe5EOXRvN2CDBhkktC9rV0tjhKVj3UlvAgXaIOJFPShp2hlhW65xzdRgai
fLvRUokiosSFWvO/GQJZ6f+yI7/koMi4/DzJTIQrPFkLddJNRVEff1VsJ+zByjqF9vjFP7PSXYrR
XMfaLeOdpC0As+mc6VXWrKRis/8hcO8+jGivlFJI0T9etcrIHDWHjyQjua7O8k0Qm9bRHGW7SxVm
P9YFB3EPG+wB8dBK82vFtDzBaqVhaBTbsjThc40eRdSah0OUpmogX6DlOwDY9NMl74hcY0XUQSRH
zdGTXPV/BUpJv0svTXRrW/gyGqMDF15UhXcaQFjSB3trrSrF5dK3WLt3YxASmEqTnxDTT/o7RGAS
k9yzDORY9+G0k28jKGtAJn321JllvmpoHlTikgyfZl4Boq93r1TUw05YO4z9KRtsWrZOVsm7Q3YT
kowUCimuwGuOSDGVmxIP7XXbEXIIZYS8oT64vWbrFOO06NL7mRBH/MoOKToFc0rTyMSxMR5vLUKi
keeAUdmY6JwLASClvZ9z2RZbcU8k0IQanyEA4R5akQh6yEF34dZaip0IpMidoBYP58J0lgJIHAnU
M3pCzpUetTsXOHD8i29IUR1/1QfPIs6gjJRBoDPmLkVyKgRLyxvvVhjACe3S4VQvkr1MiPi/FUzK
Vk1JXSef4aojzW6HGYFaTSLmPnm85AGrcrshmWVwgLYBekc8vHA72ZV/tYIkTd17Elea7Y9PN5+D
P2eEsrlVU2VI74M30hBYJwmmKwlwqPpzUZDyj24JgYWpplBAPxBkbLfKPDC/KGq+FouLgOpaLYyC
V9gMCzqXLbKsL5Lo4dSzUvpJgHok93P3rgtzDQgYhYKgt54QwE4UdnuDjTManUzOQZrAzUW9ymz7
yBoOKCyVaPA65QKZtdikLJcnc64kgPPiwTszsTcDKHhQybE6YLL+AvJvfrHwkY4RyBs0MN/rrooy
0Gxz6tFJdo4HW/oc2RZuXAEt3jjSzLu+11CnIK6nqWm3le8QIWFclwMWnbeY+N18En4jOCIB8taB
8UHEiQP/skAMnIZONuRrJAAv+Vh16nZ0e9aNRb2jog+awpCbstY0gkNljJLsvI4Wxcm0/Wkd5i6J
8xLkRiWILVqp31jTmxZULZfzy3JfJaVhYbV62+Q31/9A1YPdd1korabFveaGT7VFJCwVxtTEys+W
C6avuaTX58hp6GC0ezScoFcKk8h7RmBjgX9XoFgOEuNTwZKyBELJ8F4t/Gl86ehSC7GjfRA/OCCi
rXzkBRaxD0X8cvy5yH+zEQc3snhCRB/jL77v0ZGG0yiZksBmfjlNi00M7NQ4p703P+XQRlRfDwSh
AU14TfdrbaL0GEfzswGD5UDEZ4z8kZpYuGOyTmU89LV9eXCvkHngJHOmEsOKTi+K6+b1opC4Q4Eu
j3y/3DtCjIO0dW1OhP4+0W4FHAGawZ12gbWkXCo+EI/gWb4r0D5MmknB3e1OuCehvTu7IHVcboge
YR46bIqP562d58b6nKi5GT64ghcfePteZG3iBZqCCHFfsC/X2UyDCX4UmajUAdMrlZ6OpLM2Ehcp
W77ay/+RqZWyCU2Zod2KWmCfLkfpenQoPtZwlfdDY+r5qSkQFIQyV5xmRxJVj1n1zzPSV7B/2f8M
2B78Ntd8bO87wDvgCpYsRwGyJS2mlEKHADa44moz3xUIhD0kaBUvV9KO+di9yzDIf0unw/7GLnEe
ma2u9r7Yy6IFvBs4DBYTERsO7HfUh7s47uiNQiD7astyacLPJZBnD8ugad7AbYoK7z4s2sRX6jIO
IkqkhsEaATgDd75Pp8PJxjuUw7V8+Yl6I1UERAF1OHQXRoBeQcslCQUFlFU16khPTf4e2voQFvPN
EYKYfwFeRbI+G4lSngSuR6+L1R6vEOcEFSt325ebHnfN20nrJQhu5/Lu5ASn9sGJhXMW6JoFJEcg
mhciTw374LQT2TwFwRLeCOu8CWBrEWDheZ01NhACUGASJdQIMizmjUIYPGC/EFWsjQUmVLbhUVjf
XE1dSbvQS+j9Oub/5PItzNS7nHT6iQNnHZAWtXZt1Qsm7LNXHIapB68DimJfP2mgakvj9aEGYCZ3
xDj0HMUwTQVHTwntr7qk1Of5U6YPVPNKcjaOxz2xSETftSSXpzqO6ka5ZZWseygmHoO228Z21Cjp
vORNMlVJh6byYJFLMiQebIzHJrdbho0y7gRCmL4F/BmZkKYZovpFMsqJDFqAKDlAoG6wKL5mEFBR
hhiGWFtL8wVxVAQzvzgwH6v1ccP09CkkcGfQjG2Fha/PQneFid0MQiBViDaCLmVhD/aebYTu7RXR
MaXcOo5hyoWgc6FT+yDcHH/BNi00YMuS1oXs49hDoaINuZa4zufFsPeosI1e6Kyh2Dfb5lHevVb3
kKYXnZX4FR6aCkZqo8sDkfI/vn0C8DF81ZlbdEggz/WgDvjxgd9KIF37SNQBXt+YWVeK5GfB2SUR
6FFMUNGLImIF0NdyW/aBJEL64ITrGr8WYS3UwV4PHkMGtv/CZ8PxJnNva9r/TXoyBcfSC5VkWReW
0W7T24TNVb6DvPo47+O+GJKt+bLu4bJF1LGbSASv/BC9vLwIVVCFdwxgCbKyq3ZGH6clQBg9+Lu/
ga+M1RRI5fjOnxkBOdTRd6MuLL5Vt4d0MpdJhvV0qV6dEcQCcRnMedr/Rpi0i3Y96lT3LOOuwviM
eJnqUEAXp552jPa3ajDtOZYfRr8Fcd/Ol2rasto5Lhj8N3MFF+eewZT4VooRzHqrE0siDkFzQ6mo
O3EdAdyev2M/YNz4FX+DZKhFQWDllubs5yhlZcJQWzQU9ZY74GYlgzmWNq7gfkUteECYvy0vgBbQ
d3I5YTm6r6G7TSez+VZ2SzdEcfUzGd+YRNPwAozcMcJr4kL+R0V9SyoMSpYFoogJ10WurapF77VA
hRATwDlHL23QReAwXv1yh40xObzTwrziExSvjy2nf8JWM+SB43u591w2D87lEMXgOuoWU7USffR3
P+2qyQ+k6AX45qT+mY6V0NJxXhoCFEV+MLDQK+VA+HlTFvDPQy/8BydD55736eFwh7XUi2ISdapO
RksYg5C3ZayuPVwQJHdIYN0F3LltOd6zE/uRqRJ8vsaxC7wPmT4X36Eg/NudIjkWZt5CYvQXJ130
5KkYrfv142HxTSrF3YQcB2ILy04+MTThuNuG4kT9W8iTcR/SWWfYke3rkjl9MRWhoF81/H8vpwnJ
tYSjhd2IV9gQuFPIvA8Wiel4v0cGkFWufqqnAH7vdklGCkmjFhcxYtf6B43UFrv3gVMf+gVMmn5r
qLXTDVxEs94kbMPJU7M0JX4432lM3HJF/RKPAiKnmAMy+LytaZRsX2WJ+UGRY0E0GwAHA84Mwrla
NdrU09yBNP7LmoFY4ljwC1KZ/XlySYPLa3Mc2bHD/WJqReDbSmsXIk1kw7xDCUAcehiOU+IP0o34
xhTs07PSLhI1OaVCqPt1NaZp0Q8vyF4ukI9R1ByXRpbaZ2xuPZNkjDaxunStr3WTupLhEA3ZSUW6
rcCDJVr8lzmVikEvK9sVSwPhHUdXCvCXVl621eUWDi8J2uMD0UCuaxEA+4y01HXdithLSqbmdGm+
pGJW106YMDLAQ5EPxarlDsDVRXX3PAbo79AlBK0udh3VtzlgrZrXS+tiUP9qmJOugs9KpaE82Vw7
uysk/c90nZYMKICwl2BfID0rR25EJYsbIIAnuJq+JlrPfHoz02HDcwjMGF86ORDRT/Q4YIt15o8a
KYhJWVeSWlVlxnGmRL4T1ButpXLPRwVSfiwtpsQv/YKhofnLdzZaODkPfLip82v12VMlKrsnkH/7
TTN5P9d5M6uGyGxuDsJccAL3VQR7a2iHDHGS8im6bn+NTXf8yjk0yFJ2w2hnJp0Tprj99OxAABbG
wjiH8vUpDlyUwXf6N9ZAy/JA+8Lf7Tt6UbQEtVXiKJ3mfiw+HHwrOzGN9Jwrm8nG5vZjyQESIje1
bP+UWrxLg0u0DVPSk88aGk0y3cz5yPa5d+wpsX7h2ExJjmDL7EpH2HPO9RiPfmpmrbabIL/+O03b
fgqkZ+pde2txc9xUBotvihjZrFumNQ8P99T3+fqa6v7yoL6sC97OnCsny8ssDygac0cYxpxsR2M9
MAefr2xP5nAgjO+PdaQxdnm/nntoyg9rWPFzu4lwP6A+F/kZsSFWOmjB99DloVCYCOmAua1JJIRI
9o4lA+fMW6+UrmRw0w6+++Sw1LWfo34E9kvVdApPju7GJ+7LB7ZwCMi6Dtmk2OKWXLzNdNqiAQ5U
frmiOrJ+CQz1xRt3/Sf5ykOQXvY+OeI9Fp4YZjVaOIloOVAleWM5Ef47zfjuKV6UX8x8zgyxi2Sg
KADdZ3it6UboXjYpVKdMQJvS+X8UTL/EHIUxyY0SnaqjpxwDLDrvy/NgzUdDE0Bgv76lslbKtTdi
iWvn71I3eZLwFyCCStPRU+2oVmLPGnTBXWCcB9dLNbHEvLasQkfLlZ14+nauRvnhIvB7UibEH5wl
XB3zZkOCxypo17LE+OluYi4SuSeLqHHkoI45TP7eFdfssEeVlE56aIcFNMiQnwjlpugsLQibnYRY
sYxxIoVe8Lbxnm1K2gWFVoilY+I6EMEoUIT7eSuN18tCOeddaOBeqbk031JI/nc+Rhw18+8DGhi+
4FrscqjeBtODV6B1EtpP1cswIJpqPHnhGAKoSF2ZY65CReu/08bonq7AYaVvDqnBKxQC5KlaNfSy
I2VS4pjHZq3lrcdEb1Ppg7kA5XAXlCuxIy1lTEMevpYflr1IKfUn/lo6NGazpvgEZ+/9KMS6HjkB
3ar5Ew16P4C/TI9sDDUPQeCxMj8UP4cO8UX1jn6Txb4ZwCZ2MnMC+HjwfE0jHD/goCQJ3UbOeGqY
3W+W2YBn+DMBde0ZluZkNm7cueAvxf3A2E95p97UtzZsESUwij1jdLrte7hB0x3fnrr6jdWaXiMl
zUTH/aMU0N8OJyx7y3nZh9aE1TbZrdDiCySSXHEYiMmYPQx7JargbMDBN65jz7dLWsDbycJgxDfR
hE9GYOcl8a1ksQ3JXdP8mpgI8RvICiwob7gdb0THlFS+n53nF3LJwlwvaEon7ZrpsU1bqi4BkHbQ
eOERgK64QClZQckO4hEB7rztQAyDBdXqfMRF1HbAOR5ipR6MDKoEaoxSZ73s0As60KM7WchUXxpY
2HUJYzIfU+o7G+8MLpl45rBhtiCJyLvQABR8RPrzPDUkEUv3pa4CUaD3r+k09Dyn16xhxySduXny
ZD2pVXN5guOaRFxw2flAs/QfOTsrWlbxIOKq0Ud8f+0Ba26EyBW+Hz96chnMsuR481aYFh9+HIrp
hpOoRbduWt1t4CeLlEe3jOtTlta3glWKc9fpd8Mp/oxekQHiVlbBe3Ubq/SFUMjxnotez6yD6YMv
tvKXTtBS+5z4OCEBV+GHQVPd3YekZjF0aGRCS6sHppHEvthoH/Z4wV9O4wQKGtYjexoq+IyUqx7Z
Hu3BUsE9IcSr2jEBsCnlo15ofRTCXg5hD4UVfAlYZ8P8wVfM6dWBECII2i1REDwgPEBI42W6aFY3
3aSdIv69BsnUDEbsrKozsA1f8DzTZEFpA5lbrq+vIezA59CayHN6NoW50DxZs1/NL1cOIjeoNAzM
vM0ZaChY/87AfgE8SFHQQK8wHlSUn96X5xWlUUT7fDU0JBOYeHGoR15KBj4wrq4PbcYouzE79Z8C
b7ueiFOS1l18uk1AJdrgzhz3ASXSC2IMtNgo6F7isKXla41hwgegrFYgF4DccfwliglN1BBQDLN+
8E86WS/89ZFdXLDdvm/iMRunmlcboXvIkub9tKhqnQw+yJYszIsP7hLcVTbkuG8NJzyM48YcncO6
7Jlt0KYZlnunugtgwDiPC3F9SLtGJ3lZUsrvhfzANtgiSFZ/4ljQG+PnMHktAKuOfrFTayp0hwEX
dNvCPAF9nSzWPoaZezNl16dxecuAQjysTYYxDe2xlIQC+AydnYdyWxod3ONtMfVtlIUE0pXvSLTZ
tM87fRfxCTl4je6C8kfx42fAUI/3MdXoMl4UxPONXfI/+JjfN4A5UmL1mlG0nlmWkgI7nzCaAiJJ
++Bcq2iTcA83W31i8vVox7+eSKpX2vCAhlDMHMyZpsFvwR5LZ6t37MP+YLIImXDUkd3NgHnRINvn
XUAcnrIBljFDMq5Fg3Z9g3ldxRRO1EHgZCagEBFmLuCp1xyZu4nSqLiVe7Jjghiug9/yrJ8dxZVr
6ALJOSnFW1Z3VKvCMmkASBAo/gSXXSuK6e0xHitcvAw8SEjvfqK/OA4TkRF1VB17GeVJpeSKV1TD
eqVq7cQJ6LHwoY8esQrDfW3+MvYMtB4Tdae+O5P0A78wzXMSrTmQS3Ik/WZsWYGDUeLXRyTYou3a
1wzeTGjgt1PJyxiYBKk4RvPFtERlUPqH9EZz9glxDHovjeGhA2/kNNOTV1zOZzub2BkxMVFqOxC9
BIXe7L5kZC0FYlUcft5obaHapjxR/c4+27dzh7jHP7+lroXoSllyijaFgzfjbLa1L8eoy+oFkO/W
8tL8SgBFJ3i/CeQw164MpltLVqiLBQGG/+7SMKZvOfFdbGX78aGYB1E5khlOCixqFgOpLt1lBc34
VKHT6LCETzArflI8a7UIHWZJaEvZvZ0lj6ffoi46ILJUVFJ7R8t0f1hdsuXma/99dQm+ymHayp+Y
DThtvGthrGzq19SSXrL6hARQGFSlmXJKS4d/PbWm1xaM5i0vJuUeJk/AqZhTonxfkjKnGN3KBXMT
nhF2FhIW0OxysmIS82Tfk/lfMHaxT6wtMolvH46MdM0a29E2dB+f/h6AzhgFo563shBcPBWPm6Xl
BRO5ceKpaY4x9OEATQb3QrcYT3jxE8Xeup2eeDoPOhvi1laIgr6h0mnOfPCWc9U2FldPrNBF6KNL
UwrtEtyNVw27UJgfyQ4EvtCBWWaWrweu1fWVggJPb9f0txoVN4GeSLE+PHv7MNCCZVv0Blb7kExe
D4goLkaGzsqrZOKN7ThoYoxJgHtvqQnbtJBHfK2cp89o6gLP53+11L7SH4DYX9DEGJWD9OQFdO9D
3rcE4zp182AI3ouye6LXp+M9Qz4XTk9Bf4R5G52OEDyULNe231o78e275iSemCZYBlxyoDZ2FIlR
Ca9p/4mL/xqbJVidDvgeUiTMtfWgvBKlqI0DiOl0VFz0nuCYEoBxjlU6V8bEXCtbkX5Ci4Lcmwht
tUR3XFB2P+FJnysjtJup/r4o1uyYEhIyDQ4LZ4klmCotv+16gZPQdSICknzgU64ktM1APWQqVTv1
bclrlIiddB9go9oDlEf5jYya3gLqLIHu9HtubyKfTN2NZ109MTcLS+AwOGwbA3vquRTyfXGaH1wj
Cd5PwBwI80GpoigpCCfzssOrgb5XNakpJ6L4Qik+Bmgq+HMi9quoZ96WC3gBBXxOgp1iccN3myI0
InKZzeV6rHrSTxu2HwR615jte6T8ZqWAAMuvOnYusyzgT4p1HGVU8x8YpnpGq8H5nbu9j4KenhF4
9ZRbFWLNyAsGBVKyiFuD/9O29te7FLHSoCRnmT0hq4YTx2JDY1vmpKZ4IeksNOZRxKTEK73VnEif
XY70Lehf2MXXs6g+G83Fzz+HEAlJ6z7ea6Q1mDTwSvj0QnfTLsfLsXhGN9vzLy/an4F2LvR7Jf+V
Q214/u9Q3HqE8TCu4hPSbHlb2R2/n3TKOTY/lfPyxp32HF+4y6VwVid/y3uScY6CmSWPPZ+lpZa0
NN5pkOk9xCPW2wt8/ApmFr3yAg+WOWLJQtl8YRouO7ffVh+ssa008MMbtKnYu+MxXW7Glw8kwASy
hzI1N85WySjvqoJVsE/kZL0ggMoCe0pusUJUwZmnDlY2ZBotTjB3NYcHRoi1w+kjGJGV0m+8EpMu
jcJTyRNKqWA01iTPyEJ9lwBQ80xs6XOOPMYYhng08hGZrywUSAaAN6yCH+blZd7PB3FSy0+CX3Ys
TeUHKcibeJPKBt7HqgZgAfabAIuIwjUlMfpGLqwT+TNhh3kod1c+Zbg+Fa28OjX/VowwhdwmutGF
Z35d6+4jnKzC+Ib/xTJIVrzHvGO6dkT7PptPpreWyE6BTChxnabi72AuVvMXskVLXFv5Y3WD7OUA
Jsz6QS32jkzAnDhMf6AnNavMf0eTjPdPG3YSWQVleSzE6S9zz2qFw9gEeJTc5g5naBW6Mil4KfdZ
6uZkisCuuOiQYpVuB09DC7zsn0uwm9zWj0CFJpRuIzc+WovNal2V/uFQrE0a04P+SNsZrzLyWpMn
5a1pdKy2BGO+c+QFIPWdpGtLZrILUGCfHaMjNIGoiQD0cvb0ZZ9I4XjItd3hj6OOmDGDweWM5h3U
Q6VWl0AZVNZnNSKLi3QFZ8pqNWfhgR8yZQyM3CCaLagfSQ5qU9gzs5Vi0aFNp//klo1D6qFvFwvf
HWlTwE+wa2ibghdkLcodyvLen5muNxBSfJvrb9FNbHVjeAsVWHIxLMfydngPKOcD0hdueehY6cOu
zTcTf/JH1bcPJumXXwKdYlvX9MRbWlgkcXzOCVoQJt2e+WTB6QWIo0GTvM9MtThcIQbs6DJEhpwT
U2Wz5zA2grf7U4P4sPfVKT7kk+CI5TrHl6+baqTRK4CZHJnSZXu0zoO5nrlKHtndw3V5WTaRmRQz
gSXIew9rI5Sj7H+BO9Vs/lnX2Pz9VtmLlYXRuN26NnegF/DM2Ke0CI8k8+PdJ4xD3hWNxAUVPSoO
tncVLPsup4W5X1QoNxfmZQXzJXmasXERWTAB4Gg3mZ/S332/NH7r1ivf9yEUdNkD0tJbe380ogAU
Pc6aPS8gjy372qLydFnIiKTBeH7G8ryF4g+nvivSH9oQnWMCw37yWCbtD0y9Tm1TF2JkauTMFfLc
hPflmK+lHxazovZYJfplErD1RDiD2lwjaiuuuTYCaKd5wTth7tkS8CNWCgDj8zKRe3TM4RH2Nmz0
VrN268kdLl6jbK9k/bYZkg0nl7Hxy1CLCYk52CbpEEUajBRlChWuhCNq0COAcIAI+MtJVJjIhePk
Wzf7b68t5/y4vfkSnMfopwv8SoVYa3HY25eL2687zrayvpx2hYNLNilSlN4RbF8oy9FG0IKLsntI
GDUpjkl9XtQpd63s5onbVWthUFAcPG0vdCtb+p008iQhS5KNAU0vtE3s5lQk4j77fz4gqkxkcMsP
+7zgghsJMboRBwklwYWAnUjRTKIslG8KpWtZwf1RZfG0NBXtNSVOvHmL/49rS0OjnENKa4LeBtGi
q23mIUcLCXA/v9sYFt72Xf0/SAPXskcW2sZ55tcxa6HbSER8jc0L8mmOFDFrGxva9fDV8TnVeusH
+LH5e0pgrOJHOY1oJwA1uJm1TC9lg9zok4WK5Mn0zEBn1sJLEmBveS+txql4aTfXH2bxPAmdxY8b
AOSBlu2HvJhvVQACsKBJ2m4OslJmonFCaId0/XcipmhvHGOZtLIcd4B9L43M1D5g7UJ76tJ2jSj2
lAtwyf1H4CNCs1Am7xugNtVauSS8F1RpQqM0WCwA1hon8+MgTtlWsWKCkY+Ygcf8pvMjD0pf3lGr
nCM+P6rpX8AutdYAX268yoFoYt0PEPKFo3FP+fP+CCGbDbXx1on4fbV54973CRqjVy3igPoOZGGs
48YkzLLuWOJnKEr9r2LjOxkGh7AmXv+lboa1I9r75ugGW40b4v+jo68cLh5gHgHxva5LGXgU/tJ5
7N3h4eW1rFNJAzc/tbHBUk/b8KfYT3wGRnSMpGA/+MuQ5xEQG7TDhO+0lN2oF+jNgvy8TD85RxhB
mphmnL5BQrQAliDpaiqR2QE4S4aBHU/68F2MdRfn8+2xvfouKq4zAh8ElMxvX3fFuxXyfcLy56EO
8QZQjY10cSvt602iD1wV9wTlLyJOJE0CCmjcQXqzrWhFh4fHM6gh32BuFezsLaWzcKRpriK/vx/B
N1nzf2fe49IRv99/5lOteAEBnffzWhgnL5oFdsTxfIjIYVly3uXawggjbaQIQmtOPlmvkF1n2kc7
lA8NS9rxGTgKl+iQClHycJB01j/IQt5XsP6yv7KpAV/qkD4CnuBwG/fCvl5QkSTu6d1fesQqNCWp
sh2qub2cjJTd55NDojy4welejR74F+0lfcp+9NujgvxtlXRNP1bDAp7xvH7T7B8nq0l0579lrQ4J
4kEq3nNjX1mN12yV5FvuAm5hP9dJHcozPTeAb0+CMjY7kGb6PQgJ0r9cL+ECPxkzO1uUondlRq+Y
N9hvjhrWPIyysca6mtpdNlHZw2l5ka5CH1h8Rm+wjmnzTTHYz0HfxQv/DU5rfxcsRiGCyZvNNt4q
wwP/SlYtctvipvpgsNVDOPCwxB2I6p3gW5qGBu2sNe4+2GamjpaXGWLayIyTFSbwhQ9s2AqFh0rV
RcISMu/6Q3Stcl85BVRBYqdbOd02u/bdm6DAmF3xT4A7UPVUUnYPdk/LgQLZUP0jx8uGd4/0XdVF
tQ5fyuzAumFIrRmlfddNEGfLr8fgOEJCL3HVI6ysnH/P8d1prwoakGz4pGbsAZa65Q0YpTm8rcFF
dS4YaDhtUK1nIG5x2q2aWCQrNh5+aHDlrB80qc7tBuYiMkrMShAJNrR1Kozdj8gz/WsLvOEz1zXO
9s7WZ/J41XRlklSzu96032qhFLXI3Xk+lJpO5kWY5p+HMxT/yS1+QEE9/NyvdOkKtvaVw/g3Z9D4
UY+t9DHj4CNwG7c5idk2KEvSHNB5wMSb/3dbnpUb4DGZGnYqcFn0hGAkTO+EIJ/8wVTXVSBsmtEb
r+V5syuHYXwvxMJQmWiJApYz1uAo94PJFJCQAkWPVv/otHvBiNPP+dHUE1UgkN2TaXo+7QJ/pvQz
HwdRBlNGiGu4WZ6j2Yms1nglBqQIjC6Lu7zzUKM3JLmx/IYrjfS19rDCUD7IjqX5QTwcIKH8R/DO
I1asydrxmQ0gOQuOMjF9YvmN3rGe8wOVV6y/WvP1ZX1Ow/85KTEUEQm7WHIDXKyPlQAnbBf/6aMf
7rnNQkYBB4cs5LE7Ctytg/Z+NPTQqr6lvE6kcdhp5krEINfYm0acb8Z/E5uc9qBkj6UxpxErX/z8
7eh1YJNt3KLHdmo2wM4IAb00nGgOED/EvttJ7yfUjSgttyHevsmtApnH0mjH94az1pcPd9yyb8PO
LQNRgOruTSyDEKjMgtHJ+sJ+7iEcqqKHwCNOrrT282Y4zfKN3k4NS3+MYp1R3IyoP+6fABHMwCxF
2J4DVDUQAfiGSpny0t5uSc7i+H8wn91doaO7d0GdSgYFcBByLm6EtMhuSyRiRRxTjzIfJ6uBjTs8
tvX0GGiKQPwkpjuxsOsHt2mgGp5N6sxaTdBSRMQPhoAKY4D8+71zk8Yceh8yWJxeAtpHpcHhSo9O
i95f3/cEwC2UReFPXHO9oYMaVJUis6sI6DoXdDJvYYYarQgkLefycNKZuJRCmfCKUQ6O0NExhl+9
FEXxbDSLhBfC/74wZU2YZfc3tPpyIk4Bw4PESegDNv8RfYmDV9sq1jokiWVFK7ihL3J/QlRIRu7U
99g3wuUrWXH8S3qZMGf9OzuCWxnA63SigeYtnmId8a5hoe4Y1cpdsGxHJXsxHay1VDo/9hehS0o4
LC+MpWwalrOFC80eZD0iRvVRHXgTzwTzZeVw+/oHQsa9gRpWwhau9Z+2DWRAoyKpbIwLU2dUBxsS
Umcm/QSAjDFJK29iwgLiZ4uzYMvc5RXpsAk48saBaKMs9kp4+KiGE5nDXPIS4hArDGOUM8REaTKS
lEyhJrmN+SvYMwW5yWJOxjn1TV8Twq5pnvnCBzrqrsR93ilXEP4I1XjtdwovtUMUbSveIlSsHcdv
yfvJXh8K1aBVla7/BCKCDLgDD99wwEypShbr/axo0sZTydV6aQfWEQXdwdAs6z7JUWLubSeMnmgW
9vtJnuZzRSX7+4Ta9YCiBjKnu7N6FuANwAzVtFhc5nTwyRS9ukcxBz5s+hEQyLwRnclXd7YMDqeB
yeiJXywNrWb2Gdyfl1Og4uNIbm21iMQcxi26O2ZekzV+/XZBHNhtpKIT2jIxpoKR5XW1KbVudJLa
4Gvh9b1cTRabyq4cjYUYX84A9378RdUDHQ1K3jXKMuQvmFP0bnnPcTE7qYZBHxEubTmt3RnxD5aC
RJFDOyiNIFnvTddEjCA9vMfHtp5JxWAjn19SOa3cZGUz5gnuEnD+frxGT0NhGF26GseNaSZv7A5F
mr1osJRtjjL/X8NbWwbjsPhioCJee2ntoRtnRcxGoOl6w5e5Y5xP6S5y5aOOIaBIUAYXUj36Ad4C
sasYzzWZQSNoF1ubWWL4TX6TRF/OJ+TM5eV6LWIGl6vr8FOyoZ1ulzzU9R6b8jZ6cXzKXw+0JE4d
d39XpMndVJJ2JAafsrXfxuj3YwxbjkF1sEduEX3yYg6qLdPIQEXtKKPzsSXlKO3XPfXIdmtZPMab
DI53/9aTjl4U131q4ZyRJemaMqyV80JoB5AjbVvdOmuffIQHWw0V7QZunsUKPV4jJM2EsldXhrpv
3iDgZfekRw9Cv+W86G7ZvqhAbFX1SlPy4HIoEAaW4ONZNEQZC0nkc8ZggvKjfwRRAoa46Hr966Sr
UrHxrekN7N3UYUCv6ybOnwY4RGWjGbzLpdKnp7r19lUzBt8Q/ghiaXyWvUujMl16YN6VjLk5YpdJ
2C2lmP0ELRrFnZsTpIwdMctCQRrFP9H5lpSjglXEX5px17E0pfXbW0k2FEvTomGcLlxGyXQYwra4
XGsXjMxpx+ckkDxl/HoITtHvDfHVP5GhVlQvsoxTVRLZXUVpgmIQ6qdWoeqr6Qw4e20I8ka5XYbU
5Kr49wfCPma4gPw1yTZHdVSk3WHLGb7VSgs24tkqW6ZQj3wjiqiH2t5utn8ojI7IIxvavkAMlifW
ueZo3RsgMmn3IU7FTJgvCVH3A6v5QNVguyYyUm24/r9GkLo9Z7GUztLpdnurS8XV/QKnwcBnacs1
R5uSvcmTti6h1ocjNEFpNKTtSf1rqZ0Jp+AqP6QNFa98fBnLm275E1+n09fgZJzBqR3FDDXfQAGF
BLjaSf1K5zCmLw8gUFFiolGQcKzSA9BjOVNxG9MAFxjnCgAcpVLlbBb133h5XChWtQ1+H30WPinE
juXPQHnQT8AtiIKHjjFkEB+rlg2Eva7krzOeK2prpkmF9XXM0qhQrSNsacwDbU3fbrD6kEdV0MOo
IvtjJsxCT74EnB1qryfQK/wckNfUbL5csm/5Zi7s4wZ965+gozlukyno0J1hewkY1VBhKx7I1ziM
iK08KZlYtV4kIF9fqoGuzVL4ZU3nxwl2PFBvo4CWKhJay7b1llJl3i5yJM/Jf6Hh580kVQOdJo7J
XpjuKtBALNxB+WqnYNBUzyDwLs8vDhewe3VY/829kUMBxfGMImVuJJVpO0BJlDMcIRFQpxHeLABw
m9ar2kCeMSsSo2ION4u/klxldXLicgJAySKBdg8CtKnZHylkxw97MF+qpZi08IJF4moWi3ik0z/V
z5Z7/qFF2gCzX/j5rYwq9hSUMGP4BqqY64jyrFJPRt5WnWChnCKQw6uvBZeb23BspLf2WOdWd49o
h+2Fq0UG3EiAP/FKGQbIzlA2jgPD4gGphDT20QSH9AR7p8w7JKJEzULb+TAAtacuINHDFSNSUQC4
NIIbwejBn+9gKsPTfbVVp1fc+xnytCNOHs4CQNSR7J4xw+fOhbAe3Miwt7pwR4jKwr9XJ+JupOpA
Uvl42iMx3jf2U2aybfjQ4OH4LkiXGujio9dcuftFzVKxLFKo4DA8xMXWXyXMVXlaBbW22U8L9cU+
CR/ImIx2YoupjBuOqnkaltRjlOJ54FLDR+Rn9DRqxvy1j0RlEK566+7+gd7k2skgQLd8d6+t9rNx
YIdjgLne6XcENQgYgvVOU4YGQdVSSpfOQQ5zDjKVEcp3rf9BAw1kOi1iW5HxvoYxNGGeSZ88TJyx
HiuhPbMxoY2o/0CWt/Gnd2EMdUiEVXb0oZhUzoKdiB640941uxOOBUIDmqlouaXE3QY/iWV0nhB6
+Y6TQr4a07vAk50Rlmpc1+b/IDybgcsSsZd4UQN7zEtg4BSsVm39EaasZ71nZVIDa99sFdP1GVul
YoAcEam9ZveYiPF7ngWhoYqvEQhUFKhP2cxOH7fNgqeQiaF19aAJdRMt8+AGOxILEmONJWTMHer/
0d3QiJ1HNepl3DgUQcveJaAUznVO91ed8s3jHfext563cSc8IzN6brcAmLTi0EcBEUmZI+NlLpbD
seCxc/FFvGE9bFA8qXT0/GtKHJjT/u/T6FC50Sy0cKl11Rle5+jE6DRrObfF0qxfQdpnN/wvTuTu
d4NyZD+TYzQy3uroN8C1w3sbZ6CbC4yey2oqXvmcXro0wQyoGe16KTDcEFdd+0yAz4Em4caP+CEM
teDavunpnMVGLXRukpIdZ4wAU1fTAvtXjp8QFGq6PbqCJTW9BCO8/4kQEDGINF7r+Wv9Rn8xCfPW
l6lTqizoyWLA4TQ7tjqF7unPWwC7kDomHDPIgrJhahq5epmTkapI/jg9ALnD1OI6VXNg9pWtXCGn
W+t0m3KWe7doxYxSqPXvl59HUwtZhuKPIz9LYQHyfmsmjxMpgcat3ipsG+GaT8kWUxWeQR7yGuGN
exhkIYw83ztb9yOZZd8QQOh62GKxy9+8ljD1QopeP9W+58DKMzPdvsfzL6rEE6JaeU9DyVYFXzT4
e2VJlP+mR1oTTtEqlgsNd+3fL5UPWDx9sOR6TDw9dGxfolYNzH5UJotAQLsgWXznozuGFxVzZQCE
9BNQaRAZDGTxvckaHONQEeog5tSKO3C5HTHqoYsfjhWMOi3G1JwHNnSiF5IhHJv/jGJA/CjNCUh7
pdmX72NyDYUupwGTBAVPRqAB+ZeMshmN+re+LKLnUQimRVilgcTwsGK0fZnqyjNLkFhu3/1hsbRW
GyjQwnUsJGcijZXmOLUojamNYK8pdb1ld9AhqPgAkBNqOEgHFigem3zz+/EmiNJR049yMXjj3q4+
OgeRO1UXp0T9+tEqaiIoHPrH+mj57CmTz7263oRTrSAO8aR0KYpFdBn1atOICb8NPNNDqGlcvzD8
Yz0q/68CusgP7fJ2ED/3HQtXb9PyGRI7vHFtr25oUT1Wi5YOcOvuVMqnPqEOQ0eU6QpsPhkMrptM
0MRY7Wsph8Xutj0DRs1VClriVRlF/u6UO8nmA8FifNQqLUR8+2xIRKGrdiNmH0MnFE6NFoky/Ftk
V40MluXSY48z+BCPFFfy8w4BkPLy3Ap7789Z519UzMbXwgdX+/+Ue6EhZhQ4gahUBkoK5L83fdZc
G5t9HUKBmTOEgMBAfARYRmQa0whvAVWKlaQ1Uf2ebVvNx3v/RzMiur/Thb1voZb64Vxx6hJr4yl2
nOxHTJJhCiQd2nzXboDsD7a2GvNrqsQ7AO/oW+IQkaTEog1uxp+qsX+7WKL16mfk5kFXpTyYKP9b
TWPylZHcsHgpK53Bp3TLWZOldypgbjIWDHn3VjFl2n4FMyEUeLf/Hb7UFs83Ik00Y66L5efWU10z
BWnz8IZjsoL6bTgbGYb/3d4D1UoXpIZPQdPHwPoCX02bWuzO+0nY/itUFKYRUVm6sAb1yH9aNYdr
n5L9C3QanQpJM1lzLYGLvF+xCIDsQ1iROyIYou0fzRR5RizHwO76iVEfoSUeCRuGF0V6ShN1sgCn
DfBpyUGQZltbvjIi4ePl4ys2uYNP1xGtX+cZvt3ar5Nx6e1TxfmLAdo6iBJfvhiOA4RDZBf2GHlL
DQt89x5aZy0iLThTaXnbyWrITUcOXyTbykg1xhwl6geCvg6UgcBspvQzvvt+t5Wojfgf8mAMx7K2
haXWRvq/QYAXQL1oQUrFGiwm2ckFMVX0Kmb4bCpHKggsGokogD7Hy3HtIAsJWoPimtMKh+F/fnS+
nGQc4u3eX7TbU5CdiT36piGHA8IN969r6a91gFqBJPNu/mxKa5v5916xEcpYr7oRxcxxy4fi3dow
Jl7+KIYKt5tGOJULlP4f+gaWkCg2T5pzGRPgAy1fa9Aa7YSc2wz6/ZAknhCv9T9b+DjJ1LKHBsrQ
WA0Exp4+G1seeU95fBIgHOTWyWRcOiA5kVeu/0P1660MME69/NN+HvySRKCcTKIxlctKnqX9SfFP
RpSpMRO2S7E1hYNvPBXrBYFvR+PkGfUgi5xeRUx21AZa/RiI/7LuCQ9Tw50u1s9eMJIpElWs7ckE
xLhI3s338R600b2tLLoGjYFaL2Wo2FItryn5cRPsnHAxJ/mwfzW7PrnFINdG+vzmtfw7HSlwV9uc
MfXnF2oqw+bTxa/V92+/Z0S9p2gRVbmY5mzZBZBpxZpyf0Y2okuTZxWU2xdae1UWO66mm+K6gtzq
5RBLvs14g3g2QD1ckh7yS7sH5SkfFeHDdypytfHSobEYYliBU+admtS/uHvoXdYFXpHslbIkFAiH
H2lgkvOXJmNaTf17qktW9pzJarYTBcuR+xe6209QXyu73+unkXRXTyvLyGhQ6WEZJeCLwy6oU1oV
Cezn8DdgJMKPXyOCxA8qrKCAa3aSLtSsx/8hkkAHIJ+SAVqlN3JuVrS3enp7Jkrgb56QXKc6yU0T
gIvQOP8VEVT0YWjcoTc6SVFmQ1hHkFKku8+kh3GdJ3N5XnC1K+pPum/q9YwjRTeDGxGTyq7gd2db
8cxWcvSRNo7IGK7SvSPHmELjCsGRsI2EsmsKnmWgwSIK8WkgkRxPKAsEjRzOP8AOSmrxHbldKThu
4CF3fBgeUluOX2g2DQKIOL7ZVEIW5b+7QwdqVZLl1pceMhATpzXcH9wpEAot9Bvc8ygaYNvTdJO1
I04T8rZsyby6ZUoWR2zMeU+Ggmg+IG/3wSupgO8tqNLcEIVmlAhf9X+hoJg/bphGPBPUH+vMPyWc
5wNYEz1dohdAgHzZH/lDGNDRXX88X9Ua/Z07QJFWAoGlNAy16TJEm8PT4r9DBgSBhNBieUnJYwmZ
E1WOotPYnoBJsWvaH26Aha78HGrfTHB/CZURMQESB8E1U8+SdyfGTBBF/uWVEhG3l6xiAYcWwxat
mSM5njJMZNu4Q7zVDsrHFGyOAmjJ1PXBOeVmBwEqQZJcnxmf8cm06KSkVVKeaE0GwSILPuCr1uJJ
l6Pfjgr74TnGXatopRnlaABSTYxGfsCSQsFYrr665RbxWLlvzClwcNVHLKwu5wtCXCYqdtMO1M3M
0e18nFcJlar0zg4+V7Tcw5hQ6kkuJD9x4N8Aa/iryYJXjUnfVWiulA60pDx1MWr7T5TAjAyQAPCt
T1QC0ZXbD4gYEpPoSe2czFjLKrP+j40bzNFR+Hv7RJhj5uGpGo1vfBOHRx7rKvBqI4VsSmueFP4U
G8qL1CuzXuRCc/VdXDuoqsheMfHBbgTR5ow/MsdX5FG3c+JsgfSDQA71azQQ5bwT/+KolKCn4o4K
QxXqJYxoXkEfFIFqPb9j9yk6I+DLsK31wWyCPC3bkxAZh0JGwFs8lPKuKW2JgMAKy4I3ZsUvphhz
0/F9B5brEQEHak9t0rtGs3x9Sc+LcVtuJG2gbc3p82BYdk+78Wj+1t+DlCJN7qTrXlW0G0v+pbPQ
ZrZDJBoHLSqPLVQrmL0XRi7lFYo1NYP/7TTXe4VbFIizHttBTHIL6hCmZWc3GsMSoDbewnyCAbOv
Oc/LqbER+2059u/dFTcDjoHwfTTIRVBBzsYPwLf+S03QDuOVDeP3kkfcMUkULx8yEAcGymOlTXat
bh8VL8joW3LeS9qxQSE5FeP0OUu+kzvlf9dLHLIZB4n50R3VSC7I5SHUjOG2vXv2AiqvSbK1TDMZ
DmGvZqIq9RDRMgGKQslh7Mw8aFe5b8N3iInzm+9XnIZx3Zunn3CGZyQ1heJY1w8VbF9gZtcVnTC/
JFKEMWnRLOEhjVNJVU+tP3GZMnd1IncEQvZqDctZdCTnJ1H+ERYqKQNW87lZCWJksoWDadkgI4TY
2YkIPXrVuf5pidwRqJTC8c9pGaAGIqY9Bp001k0QIGeQ+YOUiKWaxVmsUezUboRAgjiLr7zBED77
JKMtBO7gIgxH/nopft1YvTJVU8PHoB4mp2wrb7SKlMD+/4kL0lsGzTH++Gwibm6RyNnOkRIm4R2p
I+6mTy0pATz/qzbgws+ldjg6BKIOdZMabS+she89FaSWOSjI4JjX2xSWtU4wNka0dbaiSaHYPNag
EuEmYnP7LYl4YvnytESZ+ppZW4E4aFTnvY4WpcAsqYCk7hTYiFwtxR006u6Nhjg+C1SjAVKDUSjK
rYkPGElF7M5ScIkdfsaDJpgRDyb/+uy5yldxA/yogkKX03y9BKF8GCO4KFIhjaRt9JoyxKVnAtCa
o0qa2PSQyjs+ChcHv5gn0kArzo9In3Rq7xz1ZI1uc5yNnt6n6mpayoVwqv3M2BOsGhbYv4yS5s4v
JOccyO30t5hBbV6M5TihB7mDaRlY4mypKx5qwlPqAvSLKdZoaVv2o3tzmNI5fU+G0y7fnOIUbt6S
SZHOXcKJioy/m3RPAIyQsXuDzhw6ZOSVZZKEilhTlLBcUNM4tZlpoJ9Vh84YUfaHRI/vFepGpjPo
EUfG1uF8v6YYLW4niPcJ/L7YCVFAmEBzt56p1WZ/pvI5PDYyORhzAZOqZN1K82aZK1x8yg5xE7fs
QDeeI/l/RvahgazzEWkUkJqTLwMDg39YXIxiexbjBTLvKFz24zREUumOA+6hO6HpaToYGxZpsXKa
5Y3rhim4rn7Uw/GFs72O1VLPlZlanoEg4h/Ea3jOOniVurvbyEYcML2aRHxHlRKNj+LVYobGy5+I
vSzyUKvS5qV14WpOjuLH+zHKbCCrHZAVpRwbd36xmZnLJiNMv+Qzycb3FBD4nPQ6c0Ys4thyuBQk
Et6kIRonQhW1/2g60rf1doxmjmSsybwD054lEvBA+Milue6IRf53oyDw3r1a9/omH4Dz8R4Z9X2d
JCLV7tuPbhDksHfGX7oQMKwTyfVnnbXpjW+1bzcWQEAor+r/grMsNGJVaxQIwSdpPpcH5sOFD66V
vaQy3YBR1ct9RjrgQZmOTBJyb6kBXsP2TK8aRiZk+noLDYVch3FMWBcKyqKleLkHa7Kw2xruKzjh
FCxNUr0ZUxKXIFXkZVv7lIh5lW6KnqNPb1Xx2frlZ6/pZIlSzT0zuE7mhJpVNdJKdwbldoqYiVzs
F2Y3qzC4JHd1Myc2yK4WrZl5uWbvf0CgLqkrZMo7pPdFPI/jWF8cGN1HALih61+kz8/KR/tRLhv5
Ag7W2T0BeTUVnHkfxU0VyknyHO1FxkaCbqHgc1g2r0axSbeS6U7nXcMA14+GMDphWAC2MPgOlUxP
6JWaSDS/Zcvs6SdjLwFTPRrwmtt0UUq01ValH9xhx43eXiQpPukdsCtcZ187ybLbdzn5qIJSPRMk
JH/iQ1PnySwYYpuLBfkD28YUVTTxdmHJzCtOxPcLDTzHKaHMJg++QFPm8kkR0LbGh86YRL6/F+tr
SP65gmvDnRWcSYLF+oNDWJ1pSAwC7wtfCOq3cUk27WL2mIteiSPnMRj+avOz00/ocRnXF0diJuUl
GOcsqMgFSL3IfetNo5y+QsF9s2QpnAzDFV+nYZ39pA+jkvACL1l8el+zAUW5bPBgvk+CE0aUYur0
i7k+wJvuYXA2/j5+V4En/nK1EfXLVFg/MhLZvNkrE/EQJVCqvEzRy3USag43+KEDB6R5OfOqymn6
Nsa08TOH+8rnNoUTZUcxv8tkXISrMzKAKAHhNowMk/te8scdQ4ZgpAZ9kSESpimULl9iFk3PVfuG
syktzOMG90EypNJeQoYXpTSFjhehJyEhz+ByLtRApOL2D8O0tJ30nEYWs65qkJp1HYjk2kfmped9
zL/DOKLj5hehXimlf8mJZ3E+926dkqGZqavgsDVGBqcIqLsa/lBqs0wjHTL0Bdc+IfGY1PM2k6z4
stBnE78ZPb4MXld1dqAHqF52z9QGhM7h2Ol50SsXkrCJ6/OrEhbGU+0GC8bA+izRDtUbYY6cTw6Q
klVY88cxDFteePOTHaBKEuUV0L5HBDyVB2E0gh+pVJ/Cnl+IFUyc6ZkR7LA8Ahn6rjsxbe6d7DIs
OiOjyu5peW48vtDqRQ8sIWf9cgvyuln8M3xlwHPYwGPqI6aybehF4fcBvQ2BLAhhPzlFBooOCqvK
yfYk1ZGKMWdib5aBsI3Z16jfhqqEjNinFVr+QozwUJxwMwppMyp854gxdmnKk/LefTEsCb+1ZKpu
gVmhA9l0cW9JKGX/drAT+YT630lJ/Q6ifoyg4Z/kfdvjcmaQLFsl+Q+qS3V21P/4o5ApaYWWIfby
7pQUIyBhHuAnep9OG7X24/o7bhL/i82P9dGDDayxc7mbbeouAWeU92GwAlN8gMhs45lkAfX/JHbv
tRt0aOu9zOHVv1CJSko9oF/kTGJgxRvUhY1TeHlwh6t+H8b9GXdFzxvXQWIOsWXvNeHlYTGMJ6Gx
G+Qr9BhTZmHNbzvFGJoVcvz8E0nhIlhwQozqgGRXQijnNEjEKkWsEDHe6LI9E7a7BBws1q0Cl4Eg
NsRWgM9BWM3Z2cagzz/BSlqMXJVIgmuOTSX9Ap63NDub8bEs0uILQX9hxoXzeEmZwtGlFm+xVhcp
6TFjteW3y/8Jmo68srGi4//1cLOGMA5k1nGLhsapHkOejeiniQuFt7fOwbY3hDvD5cY/2SIwnQrZ
6+3ahAbJkgdshDCsjCA7IPhRktg886r3PYmHyxh5Dy0MLmWpGCAA5HwKbJ3lkKSBA4PIUY/CTHYm
Dkxb0MVGBh+QMk1TZQuxvSnsIoSDOy3We4hL5Kv5EUibYwhl8a59oC7EiLyOfaH9WVRcKuSd0Mdl
OJW+yaQ54/cLxFNR857bFirKSBQOet4hzO93NnRcOyZgbR+TWi8xdMpFRXFFt6iRtA57i7FpI2G1
8J6IUGDruL/dVptCrUSHTj9oSoSKGmyI/L6BpLRHrZY/a+aFE/PVvqvlN+NIwJe+plCts6jCasup
xIeuSuykGByh3q6KXBrVG/d2frYE7+nupU9sT4UhdgIQhXiCGU5CUECgvnn12HnjsM0vaCcfKWgI
AkdKhsNQ840e1dmD2XwC2VKDHDCctwIRf5ECTgjRtKE5IzZcgJflRjePEFANJaIM3tQpC/2kCWiW
muyyJTBlfePZHi1c1qoTfn30fpevY9hT0WAbHb91fqdVaDeZxudMAB/091ajWQtx+mP3COHycSYA
o3nj9Bg83LnJ1GUh5XB8pxAVatAq6A7cD0tKwyKFchWrm1PrNYT/ojnCmTJ6JJwcM/lHWCifTtgX
38U8nfE2ofg6CgNEr9tBxBzal6Uo6vEYCoDRCB6kjZ+9F5omJabKgKCzHf6GO4JBv0uBo520puHW
nzufyoWqlgIj4m43zzULQbjYmbrNsKh4E2oG9E/YeCEvg+kDjXtTfV+4a4/E72cgZd386L3FqEjX
KQ76KNZkCmmHpie27Gi8GJH+WuSiiHPSlxoYRnQPEbQO0XnTlHliQKWAXNOn2XL4kif+HwzoHM7Y
KzbN7aH2yQvnq/TMmLERE1hr7y6JnAU2J6gnQzGQtASgQmzCvkTWEc+dCCEVevk/3MiV8I+pS5Eg
3EPvdV3CkSc79hhZwMRC8gWV27Rrj3csB/ZqLgyJJZtYAh8qtAVcaASxEziGNAQfpqxA5W2YRZAY
bqQ7WDbqmVsWyM/STbpfZVYUUwHnBNM/K+r94tR++tdWqgZQrGsPYWbw5bC43WFnMwh6zUN+DC6M
UMsUmhU1k9vuTE85hC4GI8EVtMh/HSDFy35txeMhzQhKG7qBvy/NmvHo2tB4f2HTWn/NfXZHbOpY
HH9HJSva2jBCWROOHvhcJy4f8W3Isep/F1XBLtVBa0+9TTDs/zM5VBjcNUDlOVFsXYQcpj/DvMfD
341Pc0F+4sEsy6HElGph7fiGN4oK/VlK0rB/tQPjHWl/5kHpgBo3STcX/7wJHHK/4lqm6HXMUMiI
piCGX6GTQNtS0yqtyHS5NkD/2fD3vnCfwq4tPZEVIuuG/H9mll+zpkO5kF8pZ4F6guvaj6MK1rau
Nrn3gTJybrnMV/gHqa0DM3tOaqyz0vzCEXYKU5kdKweExHyVfWdrxv9X39N7F9RsOrdL1GfRjDXP
1F2ejgIsz9hLTI8Ig6mmFsv7R2zUHcd4Ch1QKgyk7bhBP4sjMpHjLPNB5BEG5SBdWrhCNFdQ7kg6
iS3Fplto28vD9GLiqkRPBqAzEcscqbqYruy8yE/Q5z+zpzeJHpdskajPqFiNZTQH4m8+V1J/A80h
rkrF+HwbDNedNs4yysGILDrKoVI6dmW6OYxA2TJxd+qJJMXkfDGX5texcb9KL2gR8W6+JbW1cXrq
LmHYUoRaAY4nPFNls40Mu59jlZdNztn4OImQ22g/PhpDNIKO4lVQO5scDeZ8q/F19pcZF0hhzeH8
nT3TagTrkIQdmGpHoxZHCSc4l8FzB1BSHVXN8IjiCUjzg2YHG84rxwz8O4A0lsW0f1/H7OLeiQl9
8EULjwKL2W3ccXyvMm6eCVAofU4fIaYZuFB9mbkiluZRdrUcpZAH3pgs9vgMpAsMylHAgKFkoPch
ZOrVXpdUKN+6E52HSiJn+AoXVDCpinmHXd8/QN4d9h2KA8gIbpHyFKgzSnL+/+2tMgn8swQLopvb
JGR849WByCMNJSBak3De+uC8u7sbCDLyzJjuvrUkNVug6oEjAX5YBKt978kLcqpZeMaPfvR3OaE2
T5gB0xn54XpYq3x7PLxd2NPBpNS+Iq+vLBafiynfhCI4lgdP6MrIZBTJSk9VYbggyUyYMTZ51kBm
5tkMwjKY/bS4Cast0785Avnv2exg6qtE71mLEiF6ILd5HGr8scpXT7ohRt7lCO37PUQk9unuGFB3
PfwdSluOVkFZqPH4eIFt8dW9lQEeVPRcbxeLo4h62C0gQlS0b8Y347g6bejTUJMFwTb+Lk3BTheg
+C91eg9hoOWZd+hTy82BNU7Y0u9OSM25R/WWMnhH2fbpzzKH0rB791RSqTdP4xd4JKGIdVK8br/V
6QW7ddsn/N3Yzo/IuE0xgEo1n9+2ms5jEBtiNJhuVQoUnF5gWAH3aFvxuIMnk00fkAuFCkgoLdG1
IWqNA7TeG690fI362EMi6FyoaO89KAObdOk3B91RTkOio8SlpozJCMwYEmmqyYVdOysdgtEx/4N7
PvSfKDvoOkedCIbX0jM238HGjGjgvlYNZFYlMbMiIPP8FhSPmSVdEqls6CoDEtK5tx25zjlEyClN
w/QyvvCzfy5TP16dqM5GZDsXg2Kqy2ruOZhEOi2Yg4ke4KOYf816ZUu/WH6z0bSDzlqgo6+i6jJI
LJsQM9ctJyJNHnizyqZBtO8n1ewn5P8ZYzL4sy2081nx0mHhsGZ8lbsP05sl
`pragma protect end_protected
