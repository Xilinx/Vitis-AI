`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRnINhl3fztubDVWvJc0C7tRMbp4
9ICsocIfON/bCDzde9/a4p+f6MTC3T6AhxzhQW1gWEpzp4hol5nh8ttUdBhRuCZtSFVZZMyjN/Gh
SpOP+OSVhgkCsFIUan1MkU1GG6PY9e6wEHEvQAuXnVQ7F9LcUEyb17li4yVfCIr8b8xi26PhpV4q
2DAcbThoWqG3NLWh2Y03ESyT4lYO6Oa0joRTyfCH+PZqI/XHsn2S2x6YHeLu+DfZnMWEjGJYz2Q0
5GxCu+ONDmoC5OHIW2z0Z+uYSUdq3fyG5ILasKynUXkfGqCpDPwLT+BrHkUOfHMKOuIsbNejjJRK
M4WgFX0GjZLrWvZWUvJJKD900O01GJ/A2dYbzW5NhPwW+QhCUwYyCsG6ttOj2VTQw5L163Be55an
npXPTS6QG9mwsRIUznJwhUCjYkBBA4FzblmEJLBnVHNPNrSoB++LBjNbNOCmLnK9ubK64WnSne3N
TLaLcamHh+GUju7WQiAT1zUdNmS6Iq3ciQRtNhuDRqrmXRh0uxQoYAzcPyQi6wSfARxAKRvjnm19
i3sbVAZVdlPMYf9e01fEArcGzyBm/Sln6D8L1eVeIs1cYpf/HSVXsxamLVZasep9gGCndRO/c4sZ
8h2vpKt6pZDm6fgW8l5ZKZ/wtqgNxFYrfnxJbDA0xjWlSdEFR/vq4uywXmJW0toqLm681n3nZSyo
8xs8r/TfACbEt0WlhNVYpe2pdGSy2v2waDKpJ3a4g+6j0UbuynK7pIvEYJsyQTYaFloOPHGfwIQ7
seBP/vFdH4bZha+TXAWilQOogviOSUw2IG18jcR4ym8PNuVFNvRrvKdviBQ/rYKfV5kovv1GnsrV
VPRZRFRviVRmSO3LQU80UYYt4WHa7XNDzUsN+4x41YGN6XF+UXzGVO95i8In4LkrkONVMI6+/jL9
2qch2iBzDihC9wUeOUBepbnSf6dZkIqMVvTrdHXdv0tjGihOWsxJPDaxkTif1YiV2UW5vqbmhgCl
qCR5UfQkuMtQ50qa+gVkVhxtXvm8QDGk4LBMvF6z4sO/2rgQCHNHvSUi+eXIwVkv+FL+uxE2mue5
oU3WWoV8FXZsECJYU+CqUoPP6gbr0Ff861uX51GGXgZCg3fYPuoenRLd8zDUtfYmqKi2ML1bhv4i
mSUN+Ase1yKLNt1HUSIYPLHcfwOF1885PH7suNl4q2pG6LMu5nPkKp9s4jnV85GISV/ud8Io42fx
/v6U42VUQ2bIWSbvt4p/gptn9kNC0Wvf73EuET7+1U10S+Tv+bSu5B1kAlHKzuEdJG5dHg3ko5n1
WgNZnxU9hROTQkUOXYDVPkvqAZMPCyhV+Xq+BmpIJ85j7eruBdPnjl7f/eYyV+1JNnrMduZuvL0x
0Oe0ParAVmw/qyVe6hXyJFPZ506DCAhcceNvUDNUMl1hrMxkOqvcfZRQeTtFqOi11RZsDrHHkY5d
TxLHeRawy5Ura980m2r+2gnXdq7AD3e4XlOw7MRv5XqNggbfB2tQkps+3MFwg9rfvc9sLQENqC4P
G6fgM0Tpk0k2TYWdlE/hykuU57agCUzqqTiD4LSue/xZ2Q0o8HayxS9Qd0dXoWIky4Bd07b1qNqs
4sQFr07v6Ax6qV+OUZPtNZNQKr7clCdXjvHUvQaLQpbjkRxOCz9Jm64saZqissjQmsF5xI0dHyBr
s5pNsIWD2z2fie2rta2AdPFhlVPDx15LptwmpO1I9x6k7gPIbdGUL16/p+GPZVyW/3itRlYKDToR
bKCfC11tCSA/tmTjTuXC43bz/JCRNtUKnpnhMJTdFQpfASwbo8T2OLvxlxBk73O2sSG6uOS0HfRe
VgH65Mtmz+FXFETZ7ug29omZ8VqYejrw+iTbkX7FNbSX7iqKjVgMNECrODxuWNs5FfYT+Ryu1DM8
GPCf5h3CfBZjzrMji+quUQDKBq3pf80OEIOkTXpbGWXgJ66Q8HSRJDsGBjiGdIXByQOb8ht3RoWx
VsiMZcRZOsv6ushN29tVvLi8rKmiqhWeNtqjv7ARIqzl2nlLHnll5/gVifA3AS1WOhFVeSAl1FXI
mdjpmk2bSamQAkFwKOBsbInQ7EEj5i0ovIyWEQb7GjpjHnlWIDwJEdQ9KXDwaXU+TNFLx0dxTeU1
IQEBZ2Sc+krJibQjIw3n48HlVFrKlKJMNDorbfAqfz30Ns7b8NFC3d2AL7h9LrATG5FVWlCj0AE+
QGHAfFb8XQ1uQjeSXbDrk/ryWm1f65BXsRXB+iWPvIAwfkxuDO1m63nFq1+35MwRpfGuhM0GuVf2
mogPlB21wVOVVfpy/Mdn8D+oeVPsXeUeMj/CvYxzdwaSzO/zpu3cWEoP24JZmaSG2GU/R+LggecS
qqZZg9+MHaB6HheIAO11YoE2s7qsNFoBarGJTUzcXzlSGCLhbl/HExXKr+XI4KOvvp92/LJSwM/c
0x1lZ+rA6PWw26RTiTPpFpTfT4IvCqmsZ6hi4W092skRMRNMuHssHtkSxig0nItZT9qmffaz9lrB
gqS1xpNBhLFA/cNl4BmC3sw9QqFcDW8HlLtdWA3svhP0QB8lz3qXH+2SGWVfPcKRTiweN77CkGg5
iMFf6wp118ncdvSRvHiczK2b/w8WppVZXrVwAJ1xAB/TeA2O0IVbAd6swbga8YKM+88F6NtcXANe
YbWynd1WoXx/TPnbBhoN8OwqkMPgdm8YeZrQ3IPYeZbx6GJOIaRCJVUMWaLqectFcEqNgg1AZGe2
sJNJkN3gFPRkvbSrViNtF6utKUPRvhyeObqhyGbVxVEsCw/nSeJHvckYwWTfucO8too8Ryiw01Dt
b3hbDsHbm4rA2my8+1ePl8/is5Kd6+HyjxJttVWburj5ym/knvWDWnfC4wQrT7Nz6ZT/jdNoSzu6
vi/K6rMKYaUJwXeaZ/BXaGs0OPztUkrakzoOeQkdiJJgX+q37aGEK4ijWQ1QLmNbKKifUhOE+rs+
WaeEGYpN0Al+qukZ0dWHUr9zLIjXM704IOnSZ84cm0ps7swwg3H7wwlwHORU3ljNwyn/uO0QTTDK
IZKR4oGBGGW9lrFgIbgAR8G8PDtOhYs6rbS+2HyWnkpF0N2WekwWveESLf34T71QEbTScV6qPPz5
dW17eCcgw++Pl8+I8X3mxW4605sCfU/bndolpEorsY/YihuU3SX1R7thFp7xW2ZKFKoAos2+D0aJ
X4fZNWzbQn2aRDhfy6f7z7L44/lw5oyKCoHF+ZOazEp0ST8ryzCpwsHSg0zRKFAeBCZsv1MwIbBm
Bb+x+38S0jFmIzaUutKYXxOjd9F9zg7N5eOYIc6/b+zaSz4Q4H/CGDRe6O2Nlj//Il6Tl03LfVI+
dEslC1HO1OMX9fZzj9CE5qFnDjhdOjN8qxNDNKekABth9Jvy/eS/uslHyatlTPm7Rstrm+dQYAdi
uRamnA5TlQOIkdx1VP/bjNAGIXTgW8mA6jc2Q5z5TbuRdqAkX/oNjHWbasshujxVUG9QxEVFLrGL
MnSn8Ys0CtQZCEDIrcNYNBPGkNmvStZCbgFZ0JJflvjoKtSDFC9z5WU4mb4y/rfbwN1fNy6PGn1e
fpi8v27yvo6VOL09ST8Db9shxVKMWzWGh54gKL6pMtsBK5Q1vTKWMj3KYxXq5ZiBHQmMx+ctYEIb
XF7ZdyBeGqgPSYs0G6dR46FhaUCSqWGZimxceMAKUxLLfGkgZwsG4YmXVCyG/5d8K/YLrWrr0fe8
nv51MGwqLH1wkIlpIW6IBGoVzE2PTTRw6cM6jptCuQyosgUZuZvO5vviwKD1sBnUjyBfyURISY/v
s51aRv9V4hIRQwt0rUZqNXaQiFuB+nPNJQjXjvH6Uy1TNTz3phjcfXCiVO9T0iUL6FIV+PSVSSEM
+ACVNHO4EsKoQDY9lr2nXkJt0bdEMSMIf8MFVanJ+GQesLW3SQGmDusTd5zQhmORQhbzq8tTUrf+
0PMSNFJeSqQ29tjTVTsYihKhX2iGWmHOO4adHjIjEAYvHafpK+mzXfq5CHU1cFczRudDpBddZ16w
UesGmUjFFDb/D3dmMgu4NK9kHcY96uGI5mOEOOk/DjmE+FCNp5VbrsyaMTni0oD7v9MCvQaWh/QG
IHum5VnOh3wzcG7uz5vGpAx3VoIfXPyM7TFTZwe18f24JgchUe1Y9eIKgM+jW+uO+4kHNRX93qlB
c1opITZ/SVVWAfNh+vKdUaLmFnC+utfFHk/dHxAfh/Ss6JT1xa6BmV3r6CBArSzh0ukhq811uZ2a
XhTMf9zynLel65/oSafOSCXRJ4+Vb98lotrYPOTkD315NSDx1viMjDuNeNwSWOkw+IXnWHFLUc9B
CalIcOvQroyMpy8sVCRTEi0xMUUsKvWadfwE8kS0GJqcMFPssaPygRk+fFQ1oTxV/P33yQE4lZnk
+alPvjradVqfalWaZUDRBbY1zy5PORHw4rVF8ePX1v6d9Wsi8nJyUG8OxGkgAMBf32RyMGbb5E9w
4s+4v7JvIF+6tqqM8DxXBKqSqfaBFwbed9CMLyrIGMtIhzXowAxk3HzE+ph3yZUUHqmhMU2VSu6y
+aV08BfasYIWch2HAxGEpIVeOwYW1Ffyh2oRPK1n2hgP3a/MWrPE2daIk0BH72MtNOC7WMLf2dHA
3Q5DzXuDtFGRt24x3hV6nIcFb5NIOc6mwup9TRKiT/Sca2D5LQup3bb24PWoZr5yF4P8+zVVb/fm
nTEcVfr/dd25oX2IsEVVc9VC+OCBljzOE+WKUEfJlSyz/6jOq6BVkaX+scyOWHKqb8ddwnkjp27E
EAeAgHTbiK8Iu3bc+LiC2C+vmqXbqA1jDoEGKBEIIfgUsWsIbwFzYby0x589FYKc2jFBssSRagYB
W1dCwv7bflAQhiRHB/OAUai99q9DJ3iyMbk2MA11PIrpAtaqWP0VoX5pTw6dnrUosZ+GN2EPZd3m
+W2UgRfRNRyQBxkkP796ou3tWWinBLMxqCjMz5Xoqc2nkoATdEbqJpKumS+XxDP83flwurKfr3yJ
M/wTAAu4Gd3ljoZIHBRpg0RxdJIHlFI5cGnkh1dnabh0/EYp/m+YPk7EZFv3Nlq9Wuk7F5lFHL3T
ygh8Ho+ToU15mLNRT+SSDrO7XbiLKYzFZBdUxzokAvfeX7XdKhXIGaFHEvg7Tru5u/hPDPWiGrMt
TFFZO/hEOw8XwYFBhzVmxo3YiTElP12AHHqMd1cKpzxu0XI6darMnNpArQkPdVAOB1Jp0q6USUkD
aZ+F0FuasCPAme7ETvKUmAYMJK12WYPGX7uBa67Qh6uNa/Zi+9T54efPslRz1tdTLIb/Cf0AN2Wm
X17S4r+Iqp/6mJeClTdiIuwBL+BSTR/kg2Oq5GBMznHK+GGPex9BW5gaExdZX614fVWwWFu3biGB
iwf2+m/GBgp9r/5O3FnpK4VoUcLkVPRcCKGAIPPc2VzZ3ES0vSYZD4Xbr76LgoR+PXLIbJ8BD37J
2k4uUgZNPIThCzp8TcLBdXdyI3ws2aWx2MI6j9Bj2XvNCPbVTd4K1MOSdNQ+6o+ZMofKEFg2F8H7
5FFZCPDYvnPSOs4BJctJdaBlPr57gDwSr/hkLClpSpLQibbHncgtpU/wmeQHYsFqfaRFetejGxps
WSmPXjPaeLLR/bwKVWBPSYS+1dfawgmoIPSQZTxMZcBEz2+uj66gYXPUESslqjsGhSeYRcz1nWt9
kjr4TYecWNYra2Dpmgatb98BQ8UeecAUZ5TVEHp579MGFbmfCh+8C/SiBe9MR+TS9neWAjIqvyAI
ozJHBUgmLekfGxPafOJB336wZTY8JGQ8OuM4QhUBIUgHObQQXd0CFipj3Uc5lZ5Cgq4gOKI3xOep
IKiO/Ri4XXyNQL8TC5iABFUjd6afAe9usAIMG5pbATzkSNfYq0iE1nQP6hQh52n4Xjjtaluc8r2r
IHIjutkFBGPBN2O8q4owotX/EwvjtRTH7XywsDbIhWixOzR0WZQoa2u8gtA6xMBDJbePGRH1P2z5
367LZSbvg4cV9NxNja7Z21AtEXWbVFhWi2vlM9F0peFjVBI3pwQZOtTNrfzzKhQPcy7sWMLcvfpf
fMf5OyVZ6CPq98HhmbfDXitYKWNd/hgCrpav9RY96CwwhEYxns/wjC1nER3ljN4skLVYpPESwzSt
eh3PZ4G/h/XmLEOerPojOgwgwdZrDdDb5tso/q0ubF00SdCesYv6YD8xKLvokbtlFJ0cLtxuPhtQ
Sdtm6jcDWLuXVKODfZ/KV3yYazxxrv4PGwI5pGxGM31FOSNCpIqRYC4uvkzjtnekmU4VQ7lo639Y
N8FWvVjSQiWyCOY2p+aR9M+sekXYIw+tZcjkTDAhybTcmmc/klnKHzT7u4qQmnCMOMfVHXukoNlH
5m2nqkurNOWjeMTjhS/qxMDLX2OMh/3bqxF3wFwFvpTLQWnk91MB6rsm2PkS4WccMtW4mSbAnPWO
+PKzJrnEGaJ4G7nAXmZ9nkq9Gxcy1YF3MAV7ly5X0yBXmh2srW5cu6qIRe80wf5micdeDjwn8WfT
LsyI97p2kOgFwdXcq3WZ8gAMYVVsbVfLBp6/ZMjxHoxxg1lsG5DmiIUPLkLwyP+czOdV8+cq1Ama
ber6JxC5rblxN+KSHMAqvxMh0vfRk3TFapQbtBLWdcxXbMJvEpDyjx27vYrwSkyZsLAM2Pojpu6s
P/7065G1jGZxGfUjaddJH5hLhxCVWshkDt9Q2GG4ipFn4g02b9+H/KPggrE2T472spauyREVwCea
qzB9Ww5YyHPdZfL8ql1CjuFBxBNG2Fb+4Ltx64c8qKXFwIRN1IXr1dVelC0ZChwE/4qGGZWccB4w
Pzsi+c0Iyv6pOu5bg+fcpzUQtElMhip+Bl5q3oTEtkmVNY2h3SUWFJNk9fnT/pInCrbjJR+ou7eV
dvcH2fNiVf3ZMFWl93xIvBm4h3JHXl8RwkmpojlhGkhWqrKo2zW8aHEOO/0JIhk/b2iyCW/LVXmp
6MRLmvadhsYWVDzRI/oSDPLjCmAWXJUjr0Tvq8jRGCw1aGiv1xR+yPFG9mCOyoJCjeERHQjohfVA
Gfm1ChXkaMInWa0C5Hj88t5rMRZ3HD1sIuqgPBTpq6GmhV2YVtpTbbLjGEpORHGNkw69/M5bmfLb
lKwqjJKWb36+LWsd5iuEZ+/w5dZ4MbJb5BB8J62oFKikYINaO0y+1I/fP4lv7+uxe8OvqQm0gFR6
QLSrp0kW1zx+1Rp8y8Su1Ed6W0pk9gDbrGa2lyj1fP0Z5Y/D+nXrzBL/X5pJE3VDobZ58iM1+XhY
B6qQ2xJWknL7AMycFka3w3pWU86Sipy4CVG3/MtumPVFBQm1PPvVphyZlr5qJvoW1DowjX3Q+qr+
wtK/yAmObUVLJC1b1GlOy6VgTuZI6RmoOsskTSgVdt43guZLzpHTlvumJf5Ey/KZx3jl5/L8URaa
YjRjJwJD3KQNLDkp3K8ZQ6kX/ZVrbCCpfjCFEvhdFdEKpZnTBc5cHE3S0B84fvN1F1lzEna1jjBL
sHtVlAqp+whBDfYNiOqPbG3hpyl2qADk6mdoExILMOML4K6G37R3ZXUYAEHikP412eq2v1t4vShn
dbayymqZXlfg28zIBXUplfSzDOLIN6v4TT6Mgin/a17BIQBytt51Aih6xvfrfwxdwwN4fOOjQ+pH
6DyQFFtk3FGt5SA2AAm43Q/owpkU3DVZKPaN0W+d2z2hrjY9ruWDL0Hqraa/42CzmJPEZZbAJdr7
68j+COEsnTNStPpwoqjL6CgtbdG2F4Bb2EjYB1pNbRAfyStnIpMUlYkQ+cPlkyo/61Ou+suQFNuv
T1vk6k3DEx4D+2Le08Sg7RPxQcQEQ4w4olG/F0H0XXY/x2OxLjzKREkV91pizLmqvxkBhSn4h0xA
uTbDevj9teQHHo8NdmzfVBY4Qx544V9x83J42DBMFp/KgwXmI74joNrCvWQQ9f9TFDrEHIGXLzYK
hzpt5h3Eulo6yovBTXgfqxYi9s7yxD1KNt2D+fpOoKFnBjSbXssWzl3kEsPu3VeirTOEqIT40Ilg
tNSEAR+QClPx81TfuPhMVQjANdu3tKHoCMbqEw1s1YiRgR+7g4oo7zTdcQKqczLFmsBk9EGn1OTc
6LCpCs766yNHImc6BdKEdXwCezq7B9k4PSD874B//N5jhnlalEIv9sQhkkp9chvqQExOdJ7abEOB
7hJYCzmHJ0ae6tH6r3x9LwrZTVzuRLOOS1yLyUILjjRRLpIOBA2YS9QRFmuFcGVqucZjvx+ltJCg
Zv3MB+0qe6w7+vDFhTlF46r57l7dsHbEABn0EC2P/n7UizZwnf2lCBNGxhYu63ev2ASW8KppfbQ+
UvFWc0TkIFWYeFEHbK58s0MrabWii1FZmxyePL6jClGJdWBIBlFsPbdonmXWiINZene/ZTXD1NvO
LvQgyPtU/nb+DKGfE91wowTQqx6SAjnm5O1sBYNQkcSO291p3woG9Ll/I7OojlizAbYzfmgeuCxQ
dSObTGp8qG/sb0oEmz9EV/XpoTNcPfgd++3DxqR1dNjxuhpthsArJxbZaBW2YInsOKPqyvA9icKR
pPvETHaS7d3xqPkwcJ3TqA1wqIoKmROLuYJmapw8lwx/EWfKh995uxl+IZsRO+11XQV794yVAMJj
7Yk9K3lOCvCIODNoA2MSw7EqTTElEoRrJB9NWiyUEANkH4ftcQwtk3lw3R0BQdC9ZW9sm4n5GD0P
Cf/LzkDlkA49nWLgkTnPtIrf/OnKT1BGg+yGn+6U22AgchUJkeKwm2ZCR7IODJXi4yx2jWVEI09s
8yCU4c9NSUfOhp45SNxulhJFierspLVUMO/GwYZ788MorYm7uaiduquX1QcPmjEfvGZ7EWXWt5Rh
hKlKNGpoWrtOC/Mi7Fdb5iaw2TjCNIViySShHzry7KMYTGYjIk4Tg+seYAtVlmBrCmLRZ+2ERDCq
2CWAjcRqs+/Eo99ndc4uuG5QavvGR5ewlsYy5P01WGj7VlLR2hARdqwr2RZa+i+2SJm3oUcxasyo
cP40zSJPTwjT7uRPQykMiU2njhpTyaxcr9ZZbFGoLJA0p/EOxA2sUaIlMxp/e4J/bTNDHJshUmTA
0NfeL2e5HHigqUqF0L5me0OWlMEAk67r4gVLYDWtN7dujZDdS9ueeC/qE53MjPNTeHrmxQTqMwzB
+igGGhoeY5GVWwKjTiewXJDeT7ijXq6Of/7ydN6sH3AyZTUCCDkLn8rVSgSGdv2LRZkBmwCJBppo
azG6OLdtd02sSH5eZBHxM4dVlJ9q6XicB1LnFE0Rh/oR4p210vJFt33I0vjDZXLI331yclAEh2p9
/2CZ+6V8+teQmW+cb1SOBkTYdjVvWLAzMkrOpxo6wHyCKxqf3j11wCtvLBMhgSyYRIhXBM+l7Xe/
SFEB5R32Y02NqD/DVdbGOaOeBDoJr1ThINYAmoKRf0dBR6ze07tq2iQuTpbh5Uf1yLiVL9xxK6Z5
0uKNPVRjJ8BXZXlCB3/zoiAuHoO3EHcCrl4A7DlB/Dt2UByBLDhNsYM/rRTMncrBlXHJPv0TdZaK
I9Z/NrBxenRNN1UXh3K7mAE+QPqK/rERZAlskkY9wkytZNOOP36ORQTXC8Uzk9/ii1AIpmUa0dIM
2vv3L+lnu0CxnproDo/pWNxED5CQ59oIvJ2an7nMWTHFitEUPp5LnMM0zM1khWL1tLqeYFx8cwHC
yK/qb6BmFunDYF0xSzZWUVvd8xV75EKn07mvFi7QR4NnFbnfoFNtINW6tl8Z9E8rDZSi/EogeECp
hvlFZJE1GcjkAUX3PddeUY4LQpLmTO1AUt0FiuGtBEok04wRPmvgyLhDft6rdzAR4Vrr/4MH//ah
/bRNppbaSlKF54HIAysq6+TjO4AcjFs4fELPKhkimf0t5I2Q67ukXU4+xz31KXye8C3dBsbfrzm7
yxbAgG+hpXFlwzTppqMJbZnobcqGv93X1RTEr4mHCqqNo12OC8gb/w4WszDE8rBW2z/K7E309XMb
G17hESvNqQtOuA8BrvnO8sNbJAhfJABrv2oYBXqTh3UjgqO3qghhFI8UqBeFUxken/g4+iiIkkUe
izBWw7tXb/1qWUzpiSMd3AXpSI3+qHw6o9xLEF8zTgmbKPHKnRrjGKj23MFrpfQipsXB2yT9ia+6
EzPIp3eoshhhl1KPrlk/QY4QE3qEpaWmJdHN5fLprsCcsywIp14v1tQs4g7D7/SijmoKI4Tgmhmi
AMXq14g2D8VymqTnAYt1thvVXvkgONFg9NIr8Rh8KrJDxjZMP3kSE/pb84HvShTNmvouSSKe3uen
StpSm6B+nxp1GV+DRr2OGyWjCQ/c1Ji8d9A7mPQUyql7LcWUk5uGv4pTVGjp33mnNlsw+p3w9FZI
qwh479lwIHy7NzH4LhRAJARqjFFZ8oOXyxGGzYITNkzTnuNpVuG8WRSGM+CMZLucUnr49uM8iZyK
kAfhfNQdzNRnqxYy0NcTVvD1XgwdeKXFdKSgOFPw0dRpYRULpP3ucQ+uZ4D11n+oJHX92mFlP2cj
mB7GrO3Dt6OObO2aBUE++sOiDWE8ESxEXrU8tog5MsJ2+NSpG+DlHOFTUw9u6kCr4umMm2h775wW
wEnHayw0fir0/d1WLfs2XsaWhxYvDrSRD16d0XfXTqS8prvGralRcmD9fseqgw6K2/F/GvkOlHjH
RmVhxM9t33g1TWR221fX5fDDe93XocwA1Ex8RZdqes6u1xnJLauhlnLrg2M14VioRFIItb0gFfNc
l3rRYK8iY4luHvtv8xCfQEAOoftYuSQOnb8Bb4iAsL6leOof4QzvonSVwBaRTMoD21O9V0Hlvk3z
6syKryCcdPUYO6Y3ESvKhdxhwFcReSp7qGQ5zA0NZwbjV5h+EmdOnhKGqarVUvB7XcjA8sZR8urG
s4dds0VIPP9v88kOzRFVg+WOAg/d37etYOMiZuABbHV03dXjUkfBK0EUwUCPqSJRjEBYM/GX3vEz
OeDfw6h2mZ985TW3VMVv+OZzKk/VdOyB+Nn7MTjGN5bD1HA+MaOfSdsBIqqJMo42PZWzWLUYZNX2
x7dXR8lMFq5VK2a8LyBfx+HFaX6GT9ApuMM+fi4BE5iAVq3d2VNFvXGf56jWC9HZ5H2EPCHGMYN+
AyQJ67k0eR+DH5lq7wZNJkT6HGQz8Y8CU0ANqSbJVgvJsq1eojeRwGzcDpx67saEjPuq6H5vUUTH
Cp/A1/hdlJXlBjkcXD2mTzVO0K7t1lzPWzTRIk4o/fI0ijgJlhpJMiX6qH+QTgyQ2TcsfhQGAgJR
zDx0WbF9xn0AvLJaxisbH+Sza3jqsQPuhjSNS6ebBrJwKfEz1j1N4yeAZ/PhX0U1LkW8YmK6gvrV
gTpdeM/bV/LA8+81SRMC2yLgbndQLCKt1Wo6chqKouVPI6BARrk0Nam0brB7v0jIHYY60raz3Ure
cQzTzVpE/IkCmJ8DCuWfBWMCM6mugcBgtUIsPX/SFGUjYmOOaQ1fn4Om1/7xUTgGe08t1XA3SlmM
ECIs5VCTXEgIha2b2P1+eWgOmXWtDDrg9eYSLC/IC+T7Oc8UebtmkZdus48uCUEyfGsWJURkC69T
HAlpCtnY6fI0hyOs+wZFZlzoQ/SPLHbOf6BrzVNFnqmpoKp9oSHMxdjsEjTeITRnTgPTHOkkdeAm
EpS/GH+r1Jg5YzIr6NuO/jsEjE2+toS9ErxdRLKv87PY/poICIYw+hMJXPpoxEvaJa6T/gYWtBfS
CNLDbtCX02y/KpBxw2phAca0j6DALVRFhWj5/GywhHRoplYdl9vkLuYMt46IAFQdYTCzay1/qph0
vQpO4spAthb+bTbapZcJiZ1qFzQqm8t9ly+MT0IQVHFTpOCmcS8nD2kbjBxfaFxEGngZKo/8ig1P
FXRPCnCgv+IIn+h1VenWDCRJMkunnikZJ3gqc2Qih9/8zc/C4CjWePwTTaJ6ip3ed8QHRLGn4+hR
PshFl/WRxKM6X8GcmtE6Yzv2aY9FN525gQO+jY0jJmnvJ/Bcyo2Ui5XIXQybyavbln3ZDkddzRi/
2JGK1SSYWp3zKHmVj4pT3umzFeLfTJl0aAJZ1dLImpTCkNqsa/BHFL1E5rcPktsLXvUcujIRY126
xgGarAxe9bC/N9/+4ErPpIFQq5I4fImzn7GsH1cxnlfkV3jGJQc06K74JSg/y4tTDpW40gRynGxZ
tS8mgaDYs8tcJtWVVjf+JC+6kz7D5wixebprUKBFdEDfK6jlIxRFu12ZrX+fREtXTtciqmyX50Rb
lcH7bpGowhSmTYudRpNGDsMEa8JxIyth8noMhiT8lReQL1xHOVJmr+46DECY7AVFbFmWXgmU4gWC
DqbsePEf4XaUHQd4to2GuQQeY6trJ56jEQW93B7n4MtJvImC5lEQAfh6u+NzjX1cteDS9sxxHNVN
lz1cX+o9eKS3tzhhWLMaWUkrUyC5fzR0OyZmyFWP/S2lqx8dVlGb+3iqoSnT18S+7+do5MC2qVaz
ulFMGFUjtqrjYEuaI1q04LCkS6T4/m45ZZnPzstxF6yurNOY9ZbX6UsG8N6frvaky97GhwY6pcR3
RsQsOGkhHJTOvPy7SoFWzyP5czJiAEqgDk5qifAFhw1FVyv6TSYMu+gNhRJe3Q3VbT4ABLO1Aqn8
gMg01/84YNC2Tv5Rkj8J3yQiF9hIFTNeJF9KfvswdYCHZG22aeBdfY+w6j1Mkm4YC/gzDl5AON5+
YCkkWa7SisU6JDkX93OmcgmS7Yxg8ugYGojyOOe915ACb2fjee9v1e0KbCoMA1Uay+BRddzpg+zD
Uwk7rs/rUW6FxhqEA+aasH7Pb2K7wKl/67WHC/gmNKHgyx1xHiPFHEXneuRWR72Mx5ioyQHRAQPa
joED5asOlnKP4KdOBRRrfZU9qfWJ0o02YYgzhZdH/QJT/RX9e/NlWn5cHRJfUIEl3BV6Y7CeAE64
nFe9Amf3f5RXdrRwuJ/RWGutVCfc7pa0kXkWbCweLD2HmqTI1Nuj5/pmsVd9mQ9ww6cYqljvYYPy
tL3E1qK8qrcsetzd6Q6WhCFJLoigh7u9NqITiayw7dS6XYzPDlTw7kLgPPhjTkehX+9k/Csd+8zT
Av+IMwy7n7YKYqFATjOy6A6L2WQQ4eXs2KkX1cU7359ZwUFGnLJCUtPjzIEUKxOuuSHZ+i4MjiUk
mNt08b4EQvURdUEE3HmQupUm14mFoQu5mPy51EbJVtlJTLADXV/zUEQ69dl0J4CwmHyDWXW/2YCu
mtsiroSP3XWIiVIEz5eXciBUWgdjjRIPV2r9FP40d1/usU1aMm0a/4Z/ig7OWjCQaWNWb3yv67bw
L1FqVxzA190lEAsjSoNaBvNxgipWnRDJOdV/Pa5vLxZU1T2vz7AJt9dvVJDlUSwIuRUurg0d6Hqr
HgID+VF/iH3ZanCL6sLzXiCkSvD9Bh1QpB9poVMKlDIuW8kvN+PQhvvGSyppNgEWRfwkbBQ0ENok
xSfpkfhBg3xeoz1O5r373hUyWFNbjCqhk7uB/ZfnNHWr1877hq52ZHbK1uQBI3hZfTPIn5I1uZHS
9oOZMijyZsCdIKGD+6fiWvZ4Jjnjw0ciepn3u18uG+4sIExWawpchDGZ6cfrfxKof/7/Ji7sv8yo
NgTf96LCREPcPfgkbcgydu/WzfqGQObwOG/ZI1Vkbb1ai0SOMuWf4op7YDMyW1UwqYtdLnwupuym
HtJlJ8bHWFNGc+xl9X70Y1UlucVJI9TXBp4LbaAwEefbkMv+LbPhjC4quGetco0SmEN9Gr6UpCIK
DGcPt2xSPZm7Tx9aWwj0obrsb9vwOqG7wIaV7wfWWooBailwZ1d46BHvY2h9nmQzy8OZyqoa9PvX
fUOqTY6QZ4MvnnCuz/16O7txiwBbWxgyMvd+3HqB+rH42TUUKUgo69reYal5ew3h/QPDHrBGux54
r0cjO5Jy1bBH/ZgE62I9d7C4KrDefYEvtQz5BB1HJ18YAi/Mb6GJMZALk1QdeEOflVIosDGVHCsn
SctQ20c25NXHWc6ORgM8FxMs/Qa16AeqN+cDsmD9mm4cMT5im2dxlCI2NfRaFZGdJHkesdYVqCcL
PvgpQHmq1jRf84klxuxabUnqSFY+5hYTEiC2owH8fOg9E0LjAStriiqrRK7BgEOs/67t0RPCmwJl
sOhGKv7UM+VLg+kSUVtIo5BCMPdrZHa5UtROrQg6tV8mjyUzfODQNs/+Jc2Mw9z5AMvL2kJ9d22D
tPdd+BOTcN6YJW8zU9L9unrsSFbtEVgVCBqYsBkLNpoboUUCDyGOcK8l7e0er6mbFL6ax5nA/ebw
zwO1hCKxpHF/N9dWCYjCcY3jSEZ0VWsTnO9/h7193+v38q8doMZ5c7WCKHr9hp+dZ+fBQHnQTBiM
mIL53DUtfOIvk8/B/XIFHKPerHqy/iBuR6it+OkNaBBQWUbG/xn7BHfeVklsK0sIPPyKM+29gK/+
sWbhwrUmwTCVknxYrqWpXigEPLCN32X7BhI52cZO4ihuXBWk/ZAgz8HQ8L0LgOT/8s9n04noSCcQ
X5Kj47tXKIfSA5fXHOr44DHzis6/H08s2gF8dhSEVqOF2yF7GbIEigDep3TyUOGsCrCoDbO8qtk3
gTQRM4FLASwevHxXRJruU+a+OzytILyDvhPEghLoCiZGzaAyTjr4HYLxX+d0mCjuOh8GmgpC0jpO
aL7Hop/zRtHa0hACWuta5PX3ojrXpp7e7vixu5Jb0G4FYFWgOg9QxF2KU2UnpGEhhtVtEb1gs8xs
/W2NmCsU+GxDWIIyXQ7Ko6K4vqS+IJmtHuCFlihFSn6kdZ2WGpquw3y3v9naZtSxUB9+qMGz8iLY
SO3MTLalRohUUW9m6U8ayaphD2d49gySrzhxVE16TYf6qfecZ4V2NXCMx0hjiZsNclWQ1gRWTY6Q
J7Hv0IMAaF+b5z6w5keh10PIBDGbmYvetk450ZMhJxufovqKfsyEzo8PEaVqVAne1/lbrhu7iAlK
2VI22hcaiwTr86r0PfxxOdpzaryAAJfhB0BEdnCTkckMYLBqvvyI740WDx/SKO31MYKJhTlzCjc5
FLi6FizkrovdBlJMAMtkUDzUSghM3ngFvhCbvGobmpJ0wbvyX7OfxSJvKwz9GqXV4iKzasEYL+lq
BEbAWI4pcnrm0uDuw/99PnX33Wb/V/wFJVgRJkAzURu9c/yCalGwazGt8V6Pmmg9tljGLLnHQBbU
EfcfhR/klY1hsQ/PHpM15MHWDUK9HdTXuI53ArhLsOua8EB74MPT9taZCsS1qSyHvoNxJLgfzcPw
6rDDa1Oy0yVYmJpkL7Y+OhPIdcuVlqUMKZV0iArdW754Q932lqymokoEI4SwSKXjqGBAX55ekDxH
eIs/hYWoLYKeKOp229y9AVXbNY1yI2yocgRlKiY2lKWNyLTBm0/2ZC/cl4y5KRjT59qpQBrF5k8K
Q0NdrqPDEQ47BSQ39uSpl2fKMTMz5cjToLpoIGEyAFs3MG/q5FYIrN8fQBJmVFMO8Zg1KRigXzwc
AiNKEaSHCFIpPZ65UggrfJnO1EvjEm1gy6Ds5FtYzvsPKGztSgVbTq2GQHvvEaVax71RdbJSnpSy
7CWjgDNz4CUquTKTjKXGvHBFTZjxz0lIc4Y6z0A4xHBddHmG/dmn2D8/aaOcneLJHo1l4D3mNFq8
1ggiVgYp9mmpobe8W0gjxg43K2KrzOq6AHd6nFzbgu43JGKumh5r3HbWdYnTe/IfXYm6uNpZCGU7
eLvaXoS/zyzNH9JvqW1FlmSxMB6XpAxRa/BDU6PfIMg28afntpCGvb8eQnAY0vBLvc1IS8uchSGI
krjl+Qckc6JJQ/a+GDIC98X0P3S4F4B8A/sVUgsy5kLbro7JxwA+zqpFa/hlpBBFWC2V9s7pt4rW
XzSMuR/mtUtToqpwJtQw6GcJ2EmlSGSnzzGeByulGlfolQVV6QS/LlwFFMvJm5VmtP5h4ugjJ9kd
vrWDrMGMRBFZ3LVTaXJSCrt7N6N50CpoOyGyJ0KZuc4OE6fHPNHFlJ3gTwpUXdpq1bBdIJhEZ9kz
D6I61E+zEikY5wroLm/O3XOrPJW+G2CV+xX36s+cQrGRPjaCyxyOh/Y3zYicugz1FnIN18nI1rV1
VD3t0qD7TpJVNS7AKGf7uo76XO3anQ6SLznaCzXZGNTL4fNq2BOOyoCummCa5adqVw9uEttmSo4P
pe61IZswMqYGft0i4lE62mgZrmS+CvOQQa/eZivCMYnr39FikyOryB6A/oDwQdxpndEqZCbOyaNG
g/De6xpULXCY0+tFaNBq/rJsvjm826sXjdajYWrNpow48DmR9Effb0/Px0+XL9ld+HuHJqRa2BJ3
LQfKOsMyT+YZsR4p6N4AylMp+UKyjhO65C/OqMH5grKHGBlPhtQ4SVYVdktf79iED8ViEhkoD2QH
VUb7E9wSlzpy20tUu6IZ4YrSnShBvv1Q09LDXrVjVOrhjz/5vphpJmM/V39znBfFlvlFP6HeQtLx
aTKlgSBGVsJow4G7BJi50/CSfHqLtaqWGnmymDgJFzD1/KubcDTqp37F26EKAT4OVtz88qJfTMUv
teNwZePSDVPe5cpDkZpYJLEVA2pflwD1QaIDFeiAy9oWF9Y/W+y2lbVowVrEhzTyXW/9ztglEw9o
kdfZqGdqTDLuN1pVEu/Um0y0RXKjGsQAVt3krh25xISgOx1opjQA6SJoGsiWj6BpzhQZtPZYR9c0
UAVrdaAvQ2qc97CTi6h1H7iA7XCF+MOgutVy6qay8R9RifiJuXX2cmJ2JPi+tMItxCWwByC4CzrI
xGP0a6KwEY0pXd92UVyxVQ4njxu58pE6t211R2zcz2YlhlgYt9cVoCHlu5WFQ0sNT1A+tdtzCkAi
lryDjGNEKiGt9m1nQyuj8/qTbnXcRf9ybJlIQxGmgZZb0InoqZGsGL/NAZEiU38bxxn1kDZExYMJ
aL8bK9yLEqK2+IuJs3zM2pHNlnME6/id18DKnloesaDsIbDgYvLfKvIj6Ts7c7O5zFEIr1LQ+0RE
xQkOJBAkaUKFoAYRtQkTTFh0D9JzJZjUYhsE1PPYEBVA8XZZ5KZ7knmry1erUigrxjMChTTaToB2
QelKkLz260NGUKPs0b3OCnA0zN+fWLTWo4GjJFlO1+PJE0SomAxhAnB6zKKZMfD3AGEULDOLMfEO
Uj2pKGqfVmWA8UPseCIa0M5nIyYczLuLHEq0Op0zgBTdP165BcnpI/hwDIRmHqjD7xa5poBbGZ9w
uCXtjPqOYY8ZZ3hu9pxr61M0ROh0+Wc4sNZUPB0TIdCnwS0PDToNrfLQl9QOXuXXF0xiwN08yWdg
FS2IGIstrWokQ/q1neFIX5VKZNnGEKdevklQJzP/SsSiLGHkybLP7kpF68RwJlu4Tuy4OB+9GR3W
k1J9rZeNT2BNqg7nYKPErF06sx5Q1t886t7yRJsRJa1mwhCENOySKjvpA10XznoZVBS9aehNO1zx
8T4EIL5j0PIdzhXzv3aECdrBlr0OQEzVI7u4s2nH2hDgWFWy1FzNzSmn+yRpA9xrUOuuM5VKTsGb
oN9UidjKzU9e+W3hXO2g77iFWczAx0We6U95dZq1Mo7wdgAsHLtj0CMSfJee2h5Y0+Ma0YBekGGy
+aUz9m8QsEOHWKIql9F2uFDc26YszHrJaUMM4JGPZFkO9gZryZx4KLP0aSM/9wi4jIEI6Y6vHNXE
SPmw1LpGiJAPI3sDtNVeNl0xM+CXuaVsWn4wSX6Mt/3ZVUctrNWAo7aLKQYZY/MhQxF05RGoZxFn
tQ+VUuKMcU8K6xUnkp+PhydoBpT85KepLTrmSpjX6kzF2yfTDNtAejnGDyl3Gnqnmdao/kE42Idf
V57P+3OZosaCnJRLh0qFSjc3Sa4WGF4pfRb1t8xDU+Ednz7xy1bcFzFA3T5L6OHt8ZpIEvncbXDt
SMjICjnr/cRDnhxHWKrqhcruFLiUGpd59MRr1bDYLVzVCLf3nAQQpaGOCaHCg3NC2TLDJFwlYBi9
w2fN77+Ef9AtakGcatFeVIvv/olTREzGm4V1CtsteuYggECSXfa5QHf6qJjJ2toaU+qdbU7pi/m/
7N96fO0yq5SjUgMpBEU1ziMHVc8gnDWLOd4LCtMc/34V2Mi9y5E9WMi5uFSq2dph6DrdxyOXxoAC
Fa0gTI0U1GJmJEzRgHC0jmBnT7OhDgQ4yphZOpfWDdFBCCom9Rcae6aS3D5rTOP9fF5grmU9FsMe
/zyNKEQ0+SE/P+tGmitO71aX36TtUVQ2I8xQW8GKy0UQ0RsMktykkvPmILAGOZ12AgI/di/XDzHT
FaScYsnuaSWZieB2WFiqByrWLcXtCCcW/5cQfbz3DwRUR6fTfZ0yX5I7O3LCWYX/Z/GkwxGS8wmw
W3W3XeARAOhjgBNjLKQjIbWruU9MtzFGt7ePi5ck6r3uNPxSicynYbfsVj2GWtQ5frIL2h5c+ET0
yLmUG+0o7pRpToSFLXx5D568N3biDsZqlaMEAop/MlJFedT055mj6R8ijmgn4FA4mdrhbV8NgbLy
/v0ek1OTInXPK83lStW+R2X/ydaXAeH7+Ix8ie8TcffjIcE2gHL+633dQUBi8tzJgVMkyMhtuXE1
Ywr3dvEBk3p/yuEtiRgA6yY0MGDDFTu8rFtIoTXIoAZR4CDr+jikY7MQWs+tYeCGUgSlIeu8goV9
FFQLkolcu7tP0gKz4d26Upc7gtbBiCafazS5SNWxVLrJ/LAIoVuqc76y8ehyvVDF6rBALCfx1DvQ
TAfhzU+kNthkIlsABryNPgSWRA2TSC0JjAQiNztyNutWbJXptMrC4G+72XtwKyJrScRsI5v2sM8Z
mV6TFy9+oSGch/C6aWWfzJmvydsD9sii8wUZidUjIfL3xNldICs3ceygePLfrcjdV5VziyJEb+he
5FNX5ofzpOsSfPtK3FoItT35c1Kin8v4zaNrE9ucgs5acBfb19VfMzDdGYo457vONtvggAasFVDF
+VESLPeDg3BhT3oV1C4BSDBFf12slUK4ekjxEwqdOolCr5KUVcRrDHCmPkw4bXPKQ5IvVcsKxv64
JuE+xlswLxBHTqbtvN/Fm6qS1AseEUbQKNcfoibBhhHBvTqwslQPT147d36tX6WmUtjPN6c1DnB8
pGsLhYm7I+6F6BH3j1hNsbMuzApW7p/TZUvoF2juW1CRu8ixX1U4mt8AD6gG/muUQOB27o0/A0jm
qetgGYc4KcXGhrokXMOhqEqe7UW2ePjrxOnUpw8CIqcZHvnRMd+/wHfPxmXOaf8IsQ4pzeuGnvTx
t8JpHtmpJqY4ThhqMRZwLguiQHP/KfjYI3T0G8Qdl+00DscCO7ErIhbt1YjOwm92rEizakXOfKsZ
wonYSdKjPMbcw2KITllfp1JNdOysUzlxng+HKHNMKjZ1ZoM68zKsCoE4tXKXhqphme9ft+zAd1qo
ONxTUER3MbbmJiSRhUVlA6HOQyaObCx52amgYfJeoV8bgT7ZwGw82hHlldMPOIQDFJnspk71YyBa
fEmmeEKCuo8Z51ssCQgMTQOZQcCy3sIbK4/4tf6lGid0KvF1C2HNe64awZfUThUrY5kLFnPtLHR3
GMaUdcEyPrzegdL0bOFMluJLxGWh8cbqk1EawvDZfjacTi4FQHXZYynyAfFNIfcLWToiLEN0nWC8
IwcBt2IDLKUZsI4XkMysRbNAG15+ppEP8UtN/hioIGpTCv358FFHC0Qzla8Ex9TJoW0D+pJRe/g/
WLNTzVNHIY1ZDqnvoN10Ci9S7lsc4AHlKttmrvRDmp/687BcxUrLSpyObp3HBnlUcM91pHhCIJY/
JhxdsZQ8keZaoQwgrSO2MHIzFUOCsuohG59peVIMBzdDXATKa1DGHiZSZ4fftz97bQ8OT1tqQJtT
c9K/OxWj0wxbs8Z2LFX322+RoHfH03koOhxU8xQbL0hAZ4i+ulSAOLIsLkJDPDstfLE5B4zVSWTs
IQdPm+/i2IoU9Eboc4ci8OnaAyUhb8sR+ktngjdoMq07CnQnYyqKuS8YC4T/E5kj2NPxiip8ySUm
5eAOrBcr99Y1jE00ryVQVLllG5zMK/6hQzKcoYFLvpgvYn+RwUpyStmbulFJ48MfHcSZt5nsSTfF
tbvbdzCtdIqDg44ktmUfJyQkj53rlYCUWNCg3V5V+NWNQILeiseMLelluQvqT2Py8rIYiCNg17w4
QJMF2U0XF83Y5tvRvLZlBD7D106jhIPcVsF5WvUN4bqEa/3v6noZcxCnqg6ZvJL4RaY9s/VSTucQ
ioIs3Ue5cvnZmNMpPE2NRz4j990HgWoOOykgoJqC1/K62UsHmfA1/r5rhlUG/DcdWisbhkpRmBmE
JBN9T2QsWbX8oJGUHiLijeB1MohTu/2pfEnU1E8Id4yorv4HwYOt40RG9B3x0YyZMDjfJLpwcHkZ
bNflF6hkTLDC207MrCVr+MF7FuW/ZvJIs+9Ou9cRn8U1D+bf898FDLf4Q3okKhbhEOSuCnZFOu/B
nLgpXbS87RHVjFxBMdLXNxmHr+dnzlifLYX6F82iyLHNuGvqiOEPK4YhED8bySX+nlEpSYuYCHbs
B5J/g4w3TIVlM7z7uIqeZC559Gzu3L0FGKWkou4bGsH0TbuyVgHzU6K2CyDXOOAUy2vhXxCFyrqX
U9QK9uKQ58cL6Sizpe4VWxV8jQoQaHxOVdtgQUxFHc1mDr45bp8V/gZ0R6IuoEUUtsRnxR6YMd8y
R4Z2anMlSskcxqJcV3PT35IyoUJAN7jLtkkNPgIKY4JMvlfWNEt0qpfoz5H2yht7H/0CWO+tDOfs
6JgIbT9nmQQrcLWBgn0skfHaKmcr+MWiffS03JlOsw2FKmwjwrTMa6+ZNMNp6jny4y3xawtYQovJ
0H+E8fp5BY2QsOZ34EL8FaPAHQ5qg1UjZfDAzn55r2ARaDOPAYOLGWOArZOga+/HjWmYFMhthIE5
olThCixd4KRl9fpGQufzJnRCmQb4uaD5OLRFJrf9PZYBXj7l1a3J+CPRdt1vQYg3ziEBvtJ6B199
W9XC3WXAWnmEFt4StBbR7fF/WHV8j0pipf+uy2Nrtd1x72CEEyc8bcJxg4f6Ao91PVMAyEJ9KLpA
0h+aB+Hn99uxpDw8T1sToi+zTtKxtbtDZc2UZIgUezHYqO83o2VgSdXWbQJcCm9DbvBAvdEsgta1
L8tH8oyGptQdblZvNle8O9r03dVp9tf/zTepmE2Yxf/5+bTxFxbB938XAnKxXRKAb9elHaAwPRKK
VjXL9NWcH3Wgn0NVmveDT0oBipFOMj368ch00h5bjRK01LYXDEO77cANIWWMuBt7tcE7+NPzNbUC
WcgJSU9ebfD4I20EqS0kTScp6x566sX9BQU07h35SB+PQ99XtBahG/eUx6Bdp9xccQqQZ0dL1y2L
7CNv2/W+vShlasv0DIg1q0ZxnRIAUa/EUiScBe4GPkvX5hmfGLwvPbk67t85T56vJbquPnpFUXKQ
SomWpSAjuxHscB5dIz18DMnPRMTKqRxC4mzsWfIKph0w4MOVjUyM9UbWHK0hlzFP1E/f5JHMMyA5
6h6zVmuaQX5r5s5sDzjyf28Flj+2eXofOWfFUB0iDQ3ulZrK1ydkPn5OZQ0HLHZVgg+jGvQBTLAB
dmadngFUOBYVbR0r6PmVnf10696zfZLSO+lhjUmr67fmsdIvP4DLPuvzywwY5meLodWnYnaIAPV6
xH7by4MzV7/u/ZmRnC+IxHcK84thWdD46Ts0BruR+HEBU9j8rO206rzkkHakN4KbjyjYV09Ea7xd
oYR2g3QYe9JvPyCmGoP6Q74h+UJdM3yVbVP/Netr9R+IzsXxYqVWdm1vb6Xbr2XP6hQEJgXeQJ64
d8+KpGNi64zg0OXhiFfRm5cZPL3DmTYA8XDKRzFMnSjfJDaH4n94cqC1+OtYb+lrQUT3Il2DUzo8
Y7Blt2VLUweOxyR9LfpIOgp456FJcZYTdVRx3XqODtGCer86gHU+/y7pwAfIssAYmtdg67qdN1Yd
B70hPPkq50Ew7YrleFGXyUkUvKr94k/u4ebUJzfiuA88pEJAybCY7z095CFBQL1GIG1/QEXyT3ZU
l0ZZQuE+lKAgOpTYwObZNJ1cyViPrYYdMTJ1LmkfHfmey9hbKmX+aF8kraii7fxpaCcnjgWYMXh/
irJMRvKcdtnX7Cvr+WRPvbDtF+7hENn7jQI9CyK9MktqO4Mt4rmXzwNtkeQdpT3mn7ja5iGokP6L
fYIEGr7dbGKaQM2+TVMHOapOBd0YDvRYXv2JQRnmBUVXOBDiiJUOUvyVegHzW5Wj6cy36arZMIv5
5kOxvNRhBK/HJHRepmEaC+d3qZHFDAqEF++xjdtXDIv5B8UQjJEutjr4fv0olIAflEm9AnHhfjuM
0t5UoUIqS81+63HPO5Kykt4q4JL9WmQRZGyQjPdM4Hy4caX7Nzg2D+7FCDPYvF3RmINsdMWAeBWs
oG6CMPE50FKfzn6uipQILXPbpseL/NeUEJytoM2FX8bNaiK8gqC+NPH5VVl7fpJFiIZPWzvm7bec
v8zfrEuHdRgxa6Jsf3iOM/HQUZc6xLvvxMv7q6QglNUdeh4/FPtEUmuzZxrxu4domFaFt4FSTBsv
HFJhUkREQfs/YdrpULJ5ADkyzWtzR8TCwI6W7oJ8F1APxct4o7RZdEPP9fvPj4BOW+E06bQIILpQ
zJJ5UiGNeEqCwUtBVd+0eRUnnH8xNirt19IYQGgS5z8yDexgl+zypiTTlrq6JBRGlJsIVYMM/dqW
V4ajm8Uxn7sVy1nZnBu1Omd2IJzfrOVnWdUZzYfPrPB2Sr760z0G0IdBaYCS8Lc1vfz0yY8+i/gr
N0/qB6SFw+QSRLddvvwcTbEhTlTALJejLBtqjEAt2BwSLbYG7smT2Kx5RHeUYTZ83rGn2o5GprhC
04m4fq2LeMsGKCivGoWbFcpZ16zKCIcWhR1ZyD8+1oStv9pM5uVT22NSwOFgOqXXYp1b0SctRejy
BZiQC2yjg2moHFeIZTRLer/I4ido2neG0ii2A1p67t9egrEeqoyy8Gg8/nCgebaCwNOaFU6WltOz
jYR6pdEn/b23HkOH66THVanClevdFxSzkk/BqcWosTpJLqo3LL7B/j98RSyCH+AfYbsRYV6ZjTOg
jgDCO47XnBnIlbtD9U+Tp1KnvjaknRriMCQMfgvdgZ3WVQ2PhBKwRERLUrtDHuxTeHZh8OXWp4CU
TEDZqTYNNgF5sQAbez7sAIf/3xYVwtas1Jh6DrF9mEAZMFmTToVHdWI8JsLcfS9+z3JFkMD3rIet
LtZzl96Ki8T+B4+G3njnYqEroR5j4TUpOppZkbfIeDs1I9BeC1K3Y/dOoBtGvdQTAizkHLTLYp6U
O3h50un4sKqyayPWxNkro1cF6jruZS3QAFsUqd07ZSfhnAibqCYeyWXwV1jx3WFib5VrjGVgJ17a
Yzr7MarVD5tfpOzmxSHjD0onu7TE/l02SKNJ01UygvG+6lDQtU+D4R2t64jXFUjENWe/p31ypqe2
eoBJMKKbr+vFjZgYxUUQzcH5FxZDCcLTDm+wY5ksElTjD4j81wFyU569EevVT9sCdRZ1PXa/nyeQ
v0G4nU+t9JHa9IqqchLQZceC9ahm9+ccLaBqzqUWKw3m/L1C4xsdqmwyqgLGKBN+uL61r8TGzUwX
ltWh/1jjVF4Ej4JXVTWFSfGmqYeFKN3VkMfZRZEdd2zVGHo9osxhRCNPUgY2dSnATykfTau8I61X
5H+fAwJDlgWoKIVzJ8qXHt1OVutiHweRWSavWSju31NZIdZCKLKL6asigjzWSswYGGew3nNhgj+3
DsFulnxbKHuMG0ChKYmUeZFnQ9k5CXzlBdIQID12wnjHGspiYSYTDjHf3uFvJYf0r2ilOYd2ryPa
NyjjgWtgHPz7CzkQs4XEOPE7nYidNyt9rOXko+feG1GnYLjR8fJ339P8ZJqPYoo+HGi3INutMgLf
Zb1uwl2E6HFVNZO2kaqipUaE156zF+nV3BdPCq8sKBmNdWyFal0r8L8wxLrEo/pdWxlDff6hNSAL
r8qqviZ4qOAaVNzTMcMRRmhbEs54PoKAY9DqXnVOonaGGel/+KrrkCbGrdaunNhQPFEex8lAVJUi
AQik4orSvMBXJoS4M+RyvHvDt9GkNBIdO7ReRkgd69euC/Q2Xi8PpsGN27f60KHrngCsS1/vZ02u
Z1W7etBqt20+Tb2Vs5PHGfjQoK7BvQR8FsJX7wnGtv0lkarAyMdstHiI6UPZVfa8va+isqKiCoo6
eLBQH+l6kZkbdssl1bVMDO4Iv63fL28NmqmZ12lYm7KSFRotHiitNG6rUXmZLvnHGXjoY0iPH/Rs
IofLtCXZLBBnOZQ/Jp+W7I/mMuHxSjtQqzdjgVqobFiIYWB1A8AlplfwS5Jej4fiYbq2C+Zsadql
Zutr+ew6huCPldm0Ke/geQyG43geRRgkcOmFUhVeCEz7ekKeeWAtMPkLL2K4XcA3P+ATg1CuS+6M
X3Jh7ch4LuhnCuYbdmZwYlk5lsQMCtiyP3GFKi62+HlsIzF94JlUbPT+vT/KQgUVZD/Id9Y+dbTp
0IpC5/GkNluM4cozsZbCyJ9J3DsJ3ftSTAzY0aGRWFlFf1SSjA3bL34oAq+g4c3N3zkCDF8z9Bky
Y2UXvqMXk1P6a2qicrjaguEJFDNS/ar6fkT5WX8Dy/65PO+y56Lw50jk7Ov0rSu0crvcQFXR8aHl
XsUQuoE8PRu/Ud8hpSVnG2glsMQrQp2oCZ/IKp0NAsX3Ncgpfkj6S5q6NjMJ6GOIGxR5q7qvgUr6
3hg4+0WdpfaUrC+HQGJOVTVkls1y6VVPqq10V5SZyTI2EmAu+ewSpT2xGRmIUgDhFG0oJUAiXukt
Kyb0DkSqpy2erbRxVNiRgn6i01ZEn+kO+KRw2IYUnnPHGPVWy6/+ZPZ2Ip879wGZ6qDjxqThUxfs
J5GGVePL9VcIWWIV8nnLr8Q/Sd5x26MqWdrbQNK34l0aN3OGvOBks3C4zZ9M3L7xMU5VRiWEe7Al
L+BZrRUKlBOUnAc29/7FLmMTqeEUc1c8MQ/ynF+M0dModZtiBhrI8MF4JM7tRYA4GR1gp87AIt1Y
K03dGrmFJJPRnZBm20WwaOgOnb2QHrdeHx89VkkUV0j1DJi8135OnixryGgOvCfZC2vRLlNVqWWg
Q+YayWEXHzKIHtl6nKDN7pxzfcAdM/fR2m6SR3mFBa7B7Vc6bKcMvobF/oepfyL//g9zLMm2qfd+
rlpuENCx+c4y3wU6gpXC9KBut06meFsPcqplcI8yiG+2ou3Qt8X2MVZgaPpltcdfLyywxJZwjf8B
R1wY6T45q0aYgwPIFE3/zVdYCkuwvdC6QoS88vsMgraCMtD0nuvmdlebySfxDmXFNSu59OJzvWHR
Ec3x4IOIQYNGL9bwDaimofeDMHqT6d9voJPouRm0RQFUbt58xspBG/kvkqYuwOGdzrl+m4Ie19sh
zrfpnoYC8q2vp+xLlCQYVcY+Yq0Yn2Xhjw2UlrQCJZHbeUX8znCJyJjTbNcg+785A0Y/HV/MEl7k
1vOU5/8EIMFfmfQOkz7vhU5XBMmPFB7MKD5tHhDSfngExJm2S+DzxxFy6hFt2dKeZmheqRn8Ly9R
IKEpht9ohoe1a/2SMfK01Ilhw6tZYL07J/f63JUntu+a1jpBKRZ3WBwnPmF4+ffoBCU43oztPNXL
D16v75u3msm38EQBeK7iOZdjwzuvUQvTierfaDtWnB/3Is+hIcLr0qhEcxQhhVu2YJUMWPQEcVdF
peS02icGw7OjJ66VXxQ9nMxBUx8ZrDn4J/H1V/AyELi54e14uyEhjNpO/SwdkjzaX78ro9f2Vh0y
alUPYCFJI5ty8WRBZJ4VbgwYRQaL+9872FnahAYRhkzkCJJZOj3lrY23fXcTKQcQUW0qaLp8XbLM
wWvpvwD2v3JBTDGASPgA/3N+Kma/J+z59yuXflCizJqEy6I2aJmRkBJhe/IXXVDq44AYv/GGUkbE
Hgv6NI31YpwU+CUI/BXXSAiNFLQGuxO4w0S4JN9daZwjCZykgvKlVsVDPGZQxB4zxk0msGDNwtV0
KyKYbXMQD2+WZNSJQxNF0ssEUPQwj8jKi0uV2IurqX53Vl6eszDuoN5/LqQ/sj21Sw90bXa9uEnR
/YdyC87lfCa7mgBFozaSs5RgUzS9Af5H8VpyU1zxxsOc1/UMyAKpSvO5nynwYujs/d1m816ubgM/
VzUstG+KCm+Wd++eGjG99YENKLMUIaDeaiUws3sWDXNq8st3L9RNZD1mc0+g8sajd5/VmlTr1AN+
bZHxfzgtvTkMpfKMkKEK/pZ2l1OoIsopZUC4xq5b5iutEI0KC9cePAqVmRPhrPk0C1w53baHGpfd
5pyZ9fZIHYrkps4gSRloaSOVMhAjNISsc1z4oKGxwTrKe5NnFBeXM34uTEcF3219D1zwEdpxO/C/
USfAaoX/lgaO6jsr//tzOwzWukP/l8sjlEBAX62hE2OcumgYbzm3q/dhD+90xXG0Y2INr9m7MbaU
h6OHH4kKdCiPK77JicsCjmqy1J4VqyYty6tOW2K/cqH2Fxh3JarJjT8JV/ZymfU+HgUCFfjWgYpN
WUTR8DGwWjuj2RBZyCbjiSbZ41pSpqIImqz+A1H8hRP7DeNxqrUlrmvTIb3p1zSkgqZS5SMj2mew
mVdVMk7A4WacuU2SYbWZ/H5zZ+z6x+36Jgk7UXUXdZ4dIhYGLRF3Pm1HPKrMkBSKLymv79VEE1uJ
iw/VKKo2lBKVmESMOmwYCoaZTHXwh7eC586SbuyYdWXpGpI/B+Ucenir4GTDCo9wUGtSjHRsL5lV
GAP1OOSq3pBD3S2nX+KGjGum5+Yl/x6Qj9NB3oGhQgec+eEgUeqFaFJ9rQYx7xqnhC+EJG2GBK3q
dehG0N+K3CFSHnlBu28JmUVH48V8ND9mNnl4wGfYFq5hzd1o3NIgEu1XTPSSV7DHFwcZ45VlR5iQ
0R0bPS/JXuV4FIPo7fpxbIIB9MXRt6RhmtFphcMbFwLoawLYVLlwg54HcYAFIHTf6sOJ4Xz5z2cj
C2Gosc7r6c1dImBsgarWyXyICx5xt0YXSJnK/i37dtF0BE/j//Nn9MLuq8OqdxPQRSu4xNopYBME
tTK6uT8e7xMZzdKwvd8k7ns7EzS44dyGBRBFPWWxotw1rdZEISDznsVZ7SKniePuCDrqSeHULqXl
r5U1nmu5Hpo5vaSj61NAXcyWepbtaXb2dvRYtOZsb3Eqs4I6ey3Ji/2S4s+BNhhtKonAGFT3VUmK
TSyUkNUUTAcpiW5cfjqs+KwYQPr4nh7RhRTbgoJJl+Z54q423E62S1M9iYqS57Wv1mbd+xFqVU7R
yoZZ43hxhhxiITCKaljfIYaO9Uh6jJk80OHZqZe/h5TGJ2SGwGsOjpcJm9BhbXlFEGYXKa3ZeSJA
Ub3MwGsBuuyD0RlnR6s/KDQuAZ+EoDareVwuV+Yk0fBYlDZ5/QGzG2taJiaoBZiwxTwkVrD0lVSX
RQq5CmNp9QOAaMk3f4oXuRw1GBKgoTnudSx+58bG80N7vUjkTf9nDD14RnCZdd++dXtlSkHtnX3z
NuDIEhtmW6lulOwpev8OJYJ87zbCOzlAAwZa6PqMRTU4kDuoq0mpgEVgtBMAvcpbFkVpjEaVOR6d
GwvqnMnO7JpsmNl/VpdUnQOy5BYnjwYhWMV+/c2sciuNBzIHLj6FDj9DMNwdc+xRGuwWa94hytkA
1b4KMx5O0TnzxLWOyrj2khflZt8hJ6q1Ob2ROwO6IYJ2QC5APRUhTcc6QcAtJDZXiwrtjTyJgWHJ
nlzO6lHtkC6Nonud1L0XDH6t/cU7xMcy0zaWCfuI3ph03yYwUmz/7F1JDtgRDRtL17F+RrnVr8Wl
zBxJmwME4aT7ll6W16JWNN1vZNFhID/RnbVOI2AFW9KxrDlt8YL3Qm9dNBbfMIjHoIr3qsFX3WJd
Jpl6Bm3akNv+/PQixgxQSzRWrXha9HdVC1oCzWJ28p+wmQAJh/Ni/BQkbqRZjn2KCHT3BDkvgmk3
HfyXH70uyZKAC8QerlDe4MTL6DY12tUPm2UmBYPqazZ0hTMd+2ASObtOWLAl0akxVrjIUPa6Skhw
zGWRQbHB5g/CtMfHLBqSZRLEccJHgBvqVSx5BzMD7+nDeSZAPwL/ul2dxQreIbNQBs9Qk7e3b+YO
JXLLre4o6/IOyZZlQ6yuMWTvMXwp81lzAhnJz1fIwlmNTZBQNctR7XJrapoNFCrv5IAgnTfQ561K
Tx67cMtP3RHUMn6MycGMe5VoGGhkRTO15Hcpgd/Nioc46lods/gUfJoHedtaYiO2IsP7zqzLSv4f
1e8EQTEtyi0ZwogwKeRLXcsAP9dJrqF1kwm4Fi7272uH5Wrrsr+ZFOB+s1RXEh8rus36EIhAtQvr
K+1pAQoKQp3C02w7aahskHHmZcF8m22O9cXRvwRFdQHi7GNjpJW0pS6qTmqdCrKs8MlusPL8lvuP
Nphekd3PEo+gzFk7hwMcS269p3PkoLvAxr0j+ra+BHTedUyHI0290gKqz4Z0Q3s+o+Mgzz4oXhBQ
QpT+sQHrADVFF7TGqvvMomzJA1xJQo/mS903sC9vq3kSr6c/rLjYHVWDmW0UIfnKzVGJMftZffY2
Rg8ggaEp6+j1slnttAYCZEbHtu4jlj1lQkt4GUUy9NAfopsg+FsezDAZ+9ep/ly2oGw8FqcHYWwt
rqJ7Zm/+PE2pbY8cGKK2xIzZKyQoVNF6G/XOQOTC//pALjhG9Xm1w+CG44UE8IiVszarjDiusynq
yfRMNtrXj22xF9HbOVDPnq4yqOmWQb8enp1+hyt/stW8sF4CiraJPypWgwcXGvMyg3BlQt1Jw/jL
m6kls8vrNkBHZMqbNoQsm4PmhN7PrJGQRjxtTQUj3VypzE923uQFRV7SKEg+eXrNCd2XIFuND4tG
hQQ9SlbLSFqHHQk8ZjkzQl5N9pYJca+a8brKBZFzkNWz75wWae4WEPB4eO7RtVbfaEIKqnahRR5S
xLXR+61/P6koRjgo2xcCBt9jcR5zowFkUnb4DWjb2dMW8mnuGh2D9iQemtiq3VkFjK4+84UhucQ9
/81VN43ppoMUBhjy5STWiMqbFMUbYEcFeyniskHneSQcNPb5UIE9AX20BPVQnlThBOeTmjSARLAT
ymzqaTeCtm4QGPepJjhkYEM2iSJrKFPYU4g8VPCmMgupyV00UwreRty6/M1qWgoY/gKRH+I/KD6j
Dk6fGrdh+saMJSDuk2Gs1KtPWVE6BHMK5Y6kFYMyj5v6Es3U2VmJq/QB/rsMQsT4PIa6KG7thRi7
y917X58bx2v7Mmy8OnqddcH9+8L0OeMK4wkIHfiRskow3AYPRdzy7sbU6M+WAtwfZWsJvNfNYPCc
QsNsONE4ZcOf9Nv5wGPmvFMG1OZ1wM43UbyjOM0jPiYohwLfF0C5L/l64GKaVTimRDJWerxibNlQ
7b7+2u6aelCkA6k0u96olE80pm4zq8GKudOCL3kKFalax+EYdjAt5fvc7DeaobT7BGuFReHVIHkn
1JNYMkOPXcyqD7cecyGUAv4lla3bcjDvcPWul1QHB/iTXov3owjw8Io9Dxbr+4exfacB/INEgYRB
nXqt5Wa6iDFYIXKqoSCpu4oT7rdL4WM7jOyCYSUeL3NQnSVO1a72Ae9081ixftPdlqvUPIyvdP2t
vNUAY60y8N7Bxe2aXrpYytwVdIA7777hr97ghMouSF3vM9KcWEuAEAHP36zh4E2abuya3PM/mpT4
kpQae6S91gj/IELPe+Be3Ktn1xbEaCpAx4uowzE7Qd5O8TcmXlXCrLbRZwXkgsX9JdcAnAH9rKb8
p16ChrblDxzX3HBmUBgM1VN1g0yOJJfRnw5oUYf+HyOBhgKfxrfeNHDqlKg6iiwb/othqexNkTw+
/07lE9v4ui9JUrCWhtFANpUASz8MRZI3KRP7SxwPh0GHJX4yF8NecfFK4uZInc3kZo2XueX9hjb9
BPzKxPj6SpHAz1HcNcqM1CREF2aazGfV172umJxpjISO1cF+UxCTmJPhbLxulE23Pq47/dksdazi
Hl48l1UbzfiYTIXxL3X4B8pcDox214T9tUXJU5XsTczWz6uf9nb+5OUFq0v0r5megcPZwt5/XrB8
SEtyil2/PG6AdQRtneHpnt4aa4kpoHzmxLQQGNv4SaNxiQV2OaugVLeih2IqjfodeqCn2VEGagQq
t0dsN3S2WG9mmxpXOonJKpwuyLUhomvQ36S6zGIZWQtlXnxNJ2FmgPW9jKG/vNT0PDf5JD8hq3NP
hxWMOihaECwzD29mwqTPVmVhozxh+gGTKY2TC5ch5EBFkNsGiX7rhivaw9rJ8+VHgkBi1TyUg/Gb
XOxfKN4D0WqhVfTpAUtx6pKRb5v4UWxmCPp8yVNcG2GHfQ9pZpXT2R2ZuglfZIShqM+L7yTelGvZ
1SnovGM+k/nJFO30fqLgl6RYkDyOvaOHiYasvENNqRIzIABgvCRRbUv6aX/4urVGJBgu5VW0e/Vm
fZ7O2aRgTjIM6iU+xZYqyMG8OwFFZLQOiBfjQymNSyoxlYyCjmcpcYMBoRrGocCrofiSpU+NU3Dw
wC6PuQkFuTo5tcrfuzKWqGk3glVChL5bSIcldL0AzRZL0Lso8N5WFS940KAWT45a2u8A4LE6OAUk
HYUx14lMpPAT0QEAy6mO82EjC9lpWycbV6CxSgd1VLIpc06XzQoq55wQ/LVEcrki5OamlNYVRCc5
LMvhZQYFPAy76ZtufKSL41WWmB5PhWSRKMoQCatTf57vaJ+bLyaHF/S4OmLGtu7RvzXFx7lVY6Sc
vaicZl03WsnHpSR8U6EpPg/cgfGLdta6tWM9wDD2JgKhS48vimlF6BrjdLbo9lofSzz8XYFaAeK6
TZ5dkWepkmMqLJ/jLu2Cx6sKERijISwWYmNdo0W9/TIYTiWbTwvlyTvDi7zG+T1NcLVH3WsJF8nU
sebCRb+/30hUG3xg6SrOcrunRWLj5HyZ5VRXtu9fzMwZpRue36WH2d4KeFFXt/HwVHEeOYz9MvAZ
2OPzbrfklfaD8Sjj1sRkr3GzTvEuvCLjG3bR6XXSKezH7ptKLtyRkDEW6PABbsIaxXmsjF9wgliJ
L7Wejr+cA5NK+DMljWUvD3JBzeTEz0ZOxErGzcxR2ioJL/hGKAGIa7maud5NB0Ouk4OksllRKdLW
pX+7qAbUrrwK1Drr19HUpyIB2WeFqZowTxbdovMNUK/pJLUKF7p2mBDEt2xB8d0/3/H4RW5s4rsI
aLzHLfMdFZwh+sqYZq20Zu5KjL09A5EemE+9IoX5kFLj1pPN6GO1Z/0KcE5+LJl6IvAFXnb2FWAd
t74ey0OWu8ULhRxhNs2j7kwL2TAE6eG506hL2zJze39dw6xGW9NmhPRtOOhTnVocIvsxDQZD9pDO
mlw3J0UM2ygA7cJqicPW8sO+CnjJ0XMkVHE3LsuEslMw2syJaVbMi3peLxUi7S/Ndrz/dM/x1HtA
MYKFwtV5bgyg124PJP2qrRKRMQ2qcwSsL4UEqExQteMAz0XgsiXdjUywftb6eT+kyDKAw8UGPePr
tJ+0KVWYv6vcEp6NeupndXenM4D83iv9T8oN2hC8puVDy3TKfnSuwzq5YEo7HM5wRoU3Zsx99nwj
JUDxFoNd0ZNQO/WJ0Sye6KOA07NALPsBa6Suco9DZHuEux6vY4Jvl3qUMzhICJ9PHkndbgEJfS6f
2hYmRm+LYM8iWWxPI+2/y7RGejahq/y8C2wXshE780o0/Tsy1xC2nz0Tl8aaMZKEs1h7vJTo61Cm
oamoyuRUYgjSozggRVv38/D9RC7eUUc1TOU2fHnfkWprTq8ao87hwMQ7vfXfLOfTYmH6JIIkOxaV
TtCdnhs+Tg==
`pragma protect end_protected
