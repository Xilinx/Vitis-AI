`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQGDi5+1T0zt/Jw20/MosUf/BG/H
bU1FHIdsAm6uft+7I5naFNkYDFv6fsxdnfu/MX95XWwn1vRNirzvgSpKb5hcd4QOYknPGL4xojGp
sZ/5G0qZehfOcSBTUwqBYwtM4gmLkZgrLiUWeW/+FNXWDn0NY2ltMbohM50vnoaoynLxGMkjWGST
+ShwzZPpZgxAGOV07TAjXi7/AwOrnFMZ42eElNF/pf2qrjpzbro7vBI92w+dAWBMzWukXzhEmwut
jw0Bo+yE8cTug0oIWi2ZBhJrPfH18HxNSFDJmewupZTC7jjCNzL20zFMGBUzKmR88wC53uIA/SYq
Lc+PF0XQS38bIb2OlURVXY5mY1lQRXvyh4IgEdp55Ydci0aqXP/fwvnTNkZahvCMe4C//orCEcUt
8rTHDSfWkzbyrPd/UlyTumWbvWXRBCC9mYfk0CoUaePDtQkgI96GMBDQDIUKhXUU6nI/LFdVqmsW
53aBSvz3ViSiLiviIaw/hQ9ErncRlciverFt/JXtMiXfo2qAAoU6rQl+NBSoAzSp9FV6eQDAU/bZ
Ce3i/R6TbcwKGIk0Ueh7ZGNN72qGQRvO5w1PBhB+T1Yk7qILZnexJHS9J/N6nB+bAyREkAVZOJ9y
yrLY5HcpksLoxxQtp3IKPa0Gwvar+kArsJi/3gK4w/EF7CD3FQj3QIzze/lsyMklDCSK05LLf7vk
AIh2Vd6AN5SgFwTmnCDnw++8lSWF/8A7353kI1qJBQtXU1AEVyC069kggr2cwdpWXrM1NVkjbKhm
dyijKuzmcrARwqvwKQNybhnkLfg99Bqm9wmZeXCLvG6dT3plP0HaDpWVz2c4NiiXpJvYHsntjViR
/OmKmvb6e6oIDxj2WiY7F2r9nXjmXk2C9B+FgdNLSP0MWpzDEuIbu+Q0s0X5VNuhTfLjJTdpso12
DONmdbECXvEGkjQQ157Sgn1W79IJM4Q5wP3Cu2q/CYUFkRUebv61c8W6Z5QcSDTLWmrVUqw0YH7H
Zb5W1p4daPBI9mTGz23wX/5Plyi5JlsLWhrv+RavHO0GBEUxkdEUlP56S2jST/OH6z0jog4numLU
5vWfLddiveHt5KVA4DUY460uGNrJoLYcTIL8yR0eykE/jPq67dbwRpzOc+EAWwdqFc8lMM2ahaN8
/LiYometeCDQXbkORl0Cyc+Wt6KCwNShjYYhAG4QT8nM6MSUD3vxWKyEAGWbjFh2z9VztiXy9sz2
XsjttQiPaz7VA382NPbvcnSuAmwmiijUbeZVIraPiLks96xR/r1AeYuZXBoXA9bKgzHRSXwPZ7/E
6z7yqyVZqN9k8XWgjkTT2hActKRfviPtf+UVXjuhMY6hWQURmA1mtJuephIbaooBGZdbgSsJ2YSO
hWqfZB0ckVk6ecLpUZqTsAZQHzAoRIsj8kk6yly5ihVqRB6Rhu87tnAi0H9w7X+S8GEW/Tc0jLJf
U2KaDwxS72B4Mwd2IgTwPuM4tpcVV5L0Urol7BOgf9v5nbBC4o5emGd3etYgDW2OTWxS0pxfwinM
Mjijg3CEKspPgGF3K000CeBpcBx8mINC94hO9eu/Nxhn5ugALJIzUIb0gbWcu8XpsQxNUO1UytkP
nmDNEle/MT1b/qaedfBa5GdsKaypnC1DZ8aiqB/CFIaCFI5jp0z7D0aIRIRgwjXAr0CglKDx42Th
8BPoRSixpwGR+9MX7B0UbPU4dOAK/fsTAwm39WhKuwszN7X1HhOzQ8zY3ORpTCWNBjQagVv+SBYD
4n0+PISpJ+jvZx+uhX/nqx2pVcNDclwtdEoRwcduyeleXfMmBBGwfkWj7u2bYpqbJO6gIrgcbcXJ
2hhW5axpuqJ150evFXKylIjZTh9m8Whxhw5Gljq6VZ8gPQjAz2zEsVU2N16aVYsHtcPzVkQwgN3O
7luuiZjo6RmK4pIhXI0Zxlzmcpv1HifuU4y206Obd7Zly8qQWIccFZVLAG7XQJzA4C6VFCJjA5iP
cuDsi+WrcP5QsH7hzYsh9HNvogJ72S9BYxiHn+3NUHgR5JLivkT8mRbQdbn7HemRezvMNM3biBB0
aLk0bnIDNqmq6/dDVS1vlPFSAQaArjmaYuAzm3/2rSRcf+eWQq/uDrhx7sGSnwMmd00Ko/HyQZUp
eW+ESLL5dPkgXycpj0bCI0gqJ2E/+csE7lsVuHfcna6XvXNi4umCP8A33+1I0b8047Ae07HZOEye
bEY5G2JvZt9IYU4y8tZcnQagDQQ+BWq88stiKdVwNiMcVu5Pe52fAKUGzqDZu5ddcmT6FKA7lIgz
ZF9IDsLzDkAzkrXqVI0airr71nNXjZkj/CaFBCHbBug5/ki3s5zB6r4kg5L086kf30vvO30J3e1F
eF2w98jfpFsD2Q+OEKgehiyK36HpjOHABGy2/TuMr6ddMKLLT0QtH5FBtVmOIVC9Go0+/+aQOiUq
6LDCbgdU/5hDQqoI9a3vzVKq9Y22A0SXeGjXdwBvV1pHAeG0Ub5T1tg4kiD+hRi8KhDlA/GCanir
2IbtV0OmV+T7TL2leILRAXN+VdlBmRn6LyglzdJ9hZva+xXSCQSxSTfLI96+Aa9wQdZIQ4VLLTmF
kT2kfgm1yYVilox8j35a3mgaB59zrLbM6r58DOxOfDqDBkAAFMoq+00JufEndtxPjI2qpLX0ht/E
2VP4q1QBwm4XMELEgohqkA+LnhWQyo2ynzkqsv4KJYL5CKDMrGY9MKHXQ6G3xH3vmrw9RuqXn1Ab
9Vq/4j1c/b3JucmNcV8YcYzev/WKJnP6Jc7fsHu2WL+z3FdXYNRYlsG3fJ2QHlcTz2DOGhQebL/t
1upLUC8O6d/4/tzfijMYeovMI7QSQyt5QKjoOuO+BEsPc/lYQm6bQ27H39mTuUc+4E70hcUtSf4T
0YZM20ghuC7U8G7VfUIFqtz02bp8BD3lkFjRwGVR0Nyt9dYntbOx9EfLUMLqNdqmrTFp8Hm/1olk
vHl+cDH2y+ZnhLtXxGKQTOjGmBsGlk6JUzF1TaGE2nYuRvu2mwxPpktJebugGq73HhXlo0ulTMP8
1up0lWYX+LCosKJeQ0OnHoMqJf3CdrA0FyLqHfOoI1n3Jdak4P5qzEQ8LnnEE41vMY+XoK0qLVmv
LYTWMGr2W4NTpVoJxU+LCkU7Ur2TfDzWy0MFGopbbv6QpvtGjC4WLSYl+hG2Nk+ONU0Fy//pSUDB
QPXekEVMztKe/wLMx3GzL+rpVepBhfwo4e8PQ9XbSp2CC3VsYNT9E8/EFZwRSbmSNYRyxy8cTa6r
rjyRzRmTn9uFg8LEG/NfE+8HHfAyQO0Rcetubzi4swQWcoICZ3UM0rIwgyAsP98TLge0tg5EpcrX
S4jS90a+6aYrn2gn4tQF4elZJ3KSQhU4c4w2Y/hD1JuTEW3adIoyvAELhRLlMaXDIz0hy96UvgeO
VzW2fEOjufKQ+kl5aPAnMrzZ2Y30vTE/E4loft2H9HCTBsklGJLLJ3N9u/5ogATaGEIHVRSaOcIn
wnWG5EKF4VYqxqHgqZntFngjwGL9w3fmEA0kriFT8hDYMA0TxzMBrofbYs1ctdvDReLNpL6+uD7R
YrfYFvRPJY58KHq1dWuozFIc4Vp0WcR9RfCjz32nfhss2CxGJQiiKkh1oMJyPCDnsPH1WnGS9IiE
m7Z3WmHVlV3aGEP6lBQE4HqBgJcoxCFLYzD10A/yHtNCfUEhrO9TcdTYz1x7j+vResaBII8th6Ie
IciTVRn3WPfFLKKKKpVhWSi+MQm+mWZ+Y/Cc+Fx6tBPDecZXtLmpl2jtj7XsYbQVS8K+FiC8IvU7
HvQzKqkuRe67zrcyT11NfH6s3qbwMtvViNDTEdB4w8i/gfqClXtSXW4P6EzZHAJ1BmfbJz2kzM38
zR2/giRyXTtExkv0lTNt0fNP2cr/WesKGlHY0R8s/+UDOlYVMbHUfNCytM0m6OWCM2ZDDQ/BGm5r
MkAVfPZkCplYkWifR5v8/9vATKz/iIKvJEvR+guqtJzWvTiNOtbgwZ14+NOAjxLDxJ3YlUYmjttH
pFeEEQNnZAt2ZRLoTvojV8VSZyvCnHX+661m2nZqXjRTUJKBKEPxZ8ifCy27aOD3YrzJRj/HuAlh
2kLcEI7zvpn6Y/OYv7EfiI2azCsscKrfCRSjSfCSLbyy0aCRqYlHQbeuVl1m+v8L2/Qv2v8yfonM
NOQnjqp+8voB0GsVwK8KPtdjye70DPDDaoby3vSQFTEiMa+BLjvPRgEPGLt4hiq8KejTE0x2t9if
ECIiq++LOWMdX6U5KJvaiA1QqdYjGKlj82SR3geK/MBb6XTK3ZiTACis6kAbAwOYkvDNhBpFBnjF
Gc12NmnL9JzpPM/0PtuN3V7fUaGlBvlwATGj/SLorOOKeuo0wWFCAjQWoZLugkj1f9XZrjAk5qAo
vM1Kc9qNeo3RDkT/LlUwsLoiz/nsDxliw3WhxFsRoVFdtlL88dkrBU351pHGXV4FDCdaxEYGCvWN
dVQ5jJ2a+EyZS8+Si0JrPVO5WM1Elup/kk4DrKChfiotEgtT4q2G0XO1TNR32Gh2rrWr/JftQBWl
tWYA3ss4Bv+9shX66OcrThjZsAuD2H+CMuqA4fI7w0yaEweKK9aRiA4FWzrgjLb7/cuMHxJmzdy6
Wibh4FsvsYi2WIsYqN4UsepNdOW77/+Q1uIBdGYrs9sTBSOkbsyXDkHL16RRw2FtCcrK3cuowWC1
+Nt2P5vT1K+bf/hoa6/dA7Aw+J3B+L2wcywcZ9hEvnpUSXtKXXK5Gx/TdXXTjc1YVXr6jlgPd3I/
FG4K6WjfWDbyxvl0n3TL3pamBP8kbdUx30cSTcTt6NyzmiSft2eu41Y9IEqNN7PMQtliHPC9iUyX
CCD83v/66rPwvxTb2S2r5ugAPA+O7U/tzs34I4KjeIW5GU7YjIcYETNsq0QZm4WcQAYrbAWs3QCt
mbxidwB5+prWaY36WwjvsjODZkXU7lVqSTZQjwGh2MyRaG5JrJQXYLrHqNG/6rRUkUgX7nnUpjlF
DFYczDolUyYgBFF0kfNyMKFt8hsE2FytHytGkseKZCFzcS0o5HVBTioLOfFp0yZzn3BGa5pHGZ6d
HsnBTRz0ivTJlu0AbiY6R6MEFgBIpZyyOc28GIT1zYKKPlNpdiN3HQbCjZTJvmGVFj/ecVF3qP93
qmpMCJ4n5QyOTPffjcHVnB+pynW6Ey0kUjm4LSG5ZpluBPNlEGlR93+1boFwrwXXLez8md7dx1H1
dQ0Ayslf/ZF5zxuUa3woKNZ3FgRvuaHVWOJfAbkbWjM3nw2VjdAtVKnLXlzCHk7zGdpltFslvBve
PnXMaJD0xfIdR8T9dS1fBCa7yry6THiYACQ1EMRnsoKIwNdJKZzIn4ES1ZL96TwpMwF5WM0AN9I0
LQvUhdXkox/MY2EtRuWLHIuuBnIStuuHHB3SKZ0JqW46O5zLa8Ptol8iWsZniwGytqkSs7g83TnY
3Ts0s0N90JzD3w160xlJYx471TvoYLo/xoW9PG10w7vT4WBJGnt31FrItrzHB20vOtzaw38XO2qL
yWq1EeNRKmhbLJDc+vpRgJedCjblJwAT5kH6o/pXmK6UlQvjDjRdqHTaHD9TqxJdmduzq1x2eTrO
UodlqDLwk65xPoFLNGq0tjBjH5g9UhoY6tzrgeKJJ3zGrTcYKHQeiryGN+8BS1FogWsdyAET4yGV
hBaJDKb5XBjRXlno4FTIt7eR7qVaC/Z3VvuREKUiRmPJvEhrLr3Z2vc/xwPR8zwNaM3APQ096cei
/SL3Qpzf1nIvPlMYXBYniBH6WzAsprMQAIpr9pVyWEF/JgOzhW5NwXNvN0wiIDfXaPjkgavXzNEM
6X82sTQvNUmqtMiybdvLJ5XQkRT7jhvGaphDnv1YWhXgSt1Rz69if+kiwn3Rzi9aQDCXY7Y7wc2z
/uyX7AiH28gsfpg14UgISz3oAqx5cqTcM2Lq80QpxxlK8EnrU3iz8IhPNl9678jf/Yysc/ygXN7a
iHo65oqDCYPYMrL83nehghBcxq6lR38B89+Tf14DY9ULCAhCL5dn1wtddT/AUYoZKQT4iqHsuJGa
YVbAVwo9MAdbUYTFMXcH2ekPK+xyTDmhT7s/lRzBp42pYbcdc/PCcA/Tiv4kbAa8HzsTvz5nmGaf
Wpil03FYauWmYskKCkA/pL1+YtnR6Xp1y5IjaiXfczMhoUmGol00OSsZVD7OkAaukvzy5dt6tFNt
mryjjmkKq9gSgPaxdithcU6CUnbZeEY5oqsnDVZFkiAQFpucC3R3HC0ckQAQmo3A8/P+py97Adr4
gOM306IsXIcNVUru+FVzaT5pwtgYSD0gbDU5Iece595eVqaCFOL9k9SHXQfkDjBCOvIGIT9A/Fof
Zk3O6SO1gmuUdKWqPEMIEYXIMtS3zmjFbo/wx7pYtBHwEBpIQ4M4f+gfBlZHcQXOeuvh83qik1PH
iHM0TfhNMp+129IFc4m8N3/Pnad8HmwUj7IRN6Qqq41P10gbn+COmVwudX3PxOQOMArpL/qDcIgh
WjKLIRLN9iqv8KMh97WdDDkFfaL8UiSN8mMYKfheGvoJIwGSOggz1oTi2Hslvj4pgPENKzD4XxtR
YA+RAE7Cx5noxtOBpspvf60WlA8tqCMmewDPHYbP2KN4+jST8CWmTrh6D+ZAoe8PlG/6GcZND1q0
N7CqWzNNowZ9BL0mIYT7rLKIaqnUHcwnvsdIeJ4ar0ZbcYS0eiVCCRPCcHEBqI5KsURlTFqCYBXa
3OV25v7V/sYJ2el4j+joJ6EI7lz97spjVPq/PeBJ7YQSqviHe8F6qDFtYQ/X2vflEWagq5nJXejN
66zNwRaOxtQ+MDd34u/MQ03JtvoB/V6x2zFdY6jh7JtoBVQTg1Pl4lfiqGWUGiZ0EWRQ6JYN2DrJ
muYfzDaxVwZDK/wG4j0SRU+HzmCTEVTC+tJFHndnGoICSNxxnG+UIXtT6mDxsvZ0VZ8nt+1CZcPX
51l7OZ2n1ttLOsuTFRhu1fTdb/5dBP+YCdqPKteaei9DXCUWO9QjvgyQdkuRUe3n5QP9ToFZMsNQ
6IjMxV/wMpRurBTJTig8sFTo2vbCKxiwCgVxHuaTZT4fIKMu5DDgeKMtT5CDzlgolkikvag3H8HO
da/cPfqlQbwMRMc+Zz7316BZlhiWmU4KWp1qirJbhfmh+f2z34xaKyYA+Oam7K8mwMgS9ttDs3bV
KiMVazHCyDg5vkmbkXZtIzMvKZ4yNQiu7fIAwC1Foco38kUWpdNVjfpAkHc+NX3sKHCVMZjUixnI
4Z5b7fofpSbs6iNcDr2BwWdqgPFwAwpw8/gnZxXi1Ba+SvTho/tF3hUoiUj0aLnuxmWX+x9TaTZM
CFKKBeGPMol74biQJsBdEYtGupKZSwf/veYBpQoEY1NAj/+g4w0ymUKYSgu35CWifFzoi+PDmZYm
+gPWKGqfKXh0DkjMsAYUbV8bOAS8HU3eZm0iqfbWGr5h4c/T9RcG5eBnCQLdchAf/iFmCp9NZZsj
JWU4WV6/9cIcTuxZqEavfHeEODr8+du7XR2cK7tQv8Ge88pvq16jtnaYZiPAJg4c7z4XrxkQwbyb
ir4Hx5RklWse5PGgXmB5XMn1aNwo5btgvGCRUPBROUZBouaGEoUA0sd5l8d1ZhlWpOVyC4N6wtq9
Oelx4OK9S1o4pH90UApKgSqnQNW5hVvOt4lECb2gNXQN0ar0mXM/L2DvqNDj6VbckfIqwTgcCM4B
T9fnHv8Pd/nW9X/cQY6sRFhrO/VgZDeayqwgKhoXhqkyFCzKQ2NG3HxS9y3wJcsoHCg/+TVICgTJ
V+dkEZ6osXTaPVMgKk4hIzA3i6acgsF4XaIHDMo77tqI5GE45lrN8EkTihEb6KaT8w5/a2zrWefU
EORYri2ypuoyK5wer8KQ+BaYjZu53Ik/U7McLzdpzgXFh2SfbqXpkQfzftlTaLlyQ9e1Fq465ItQ
gymPnzqEaCOY/geVdrywgussJtEYj0zR9HeILDakrTUScBm/ZOSXwK/quHrdBJyAdrhoo5A+WKGj
D/L8LTyRsmxve7iHmKSanCo2exR4Igmf2C3I42WGO7rhxG4KDO29UiJRx3m2PnbWSPJdWX7eAZSD
xrJY7umaG/wRJThfnNhFuRAI6at2v5DBzIF6Ab6BlwXdESWw16wcdwaQIeLdMS8OaTIOrZFHpPoj
iby5SXEFs1ORxU9KZ+sQvMUezvYEoYGRpPabRhgRA/My/lyXClR8aoAWrxtgnIkM4gbeMySuQYbm
x6gZC3zjmJPIbkdeFlKUhoE/Zxu4HM9RnQCPBYLRz/zx/XHIzB+7LCA/vsLz1qFiFJvailctiasu
2bGm1K+HAjtLsspFW/DwNodl48JACS31JjimrxcBfUAefWTIwaPfdZSHf1V1PHwsHhZ+ybH0kzhb
Am8leQ/y8GHONAcQbhG6nMZARnbrIvnih0HSs6E3T2wOt9q07pR9sXsC/jUFsJ8KR+3D7Re2uuQ8
rZeHxeU41c9ebSzOIxsazmMcRkYnkTfQZd1JqHW0PMP4FCgFfoJRkR8dmq2eJJU5TIGxeMYVEp/l
Wr/Gw4Jz4x8OgqljbWXsuSXe5IMOlsARQ6VotrYuXcEjFH4xQ2XGCDbCh8Y3q1DFSVEFLg51o9tM
jcV3cBOLkcOKtEhAolbnFRJCfBBp7ZTqgnfz8LVD47OP698i7weu9R+n6W39nl5HtCrpOXPM0T+w
rBM95rPtCYidunp84sKTbBqzcZKLNWnUKKix8VguEHuQsxv+8egOriE8DwyaIlY0+MPWMMAP8LvC
aUjxTZF/BwhVq0yrJ7ABZhPkmKEGqVUhJJcO0J4J1Ztbk3eUdygmYhe0uTSwygSj5T39HWwQKYfm
yrvwhkFdUdrliHsTpGIGM8MjibSDDYnN+hM8z/kE0bibLVDQ7tsZu+yrFbyplPE6rILolQiezDEP
kXvqKmXZg+OOxRrj9KocnqXlx3oi5FBNRlmQ1X8+lgUDdikVjWz0DKMfeyRk+EEW54ZT9hwQOA6h
2NoyzvaB22trtqqFPmtMB43wWYNZ4x4DngwYWJ9eNOSY8WufFTajGYLPFvKqbVSmXZgiTcjQ/nh2
n0cdmsbgWb685Qe+F+DO60OG8qpnJ5pZI6q6/IWtMfol4u70+MhdeQYJkdRidHplkz34P0WId5ti
E3KFriu3NBdqgdVLDalXvey0u1J2DEKVUkSciDnT10BmRHVD/C0RGEL5nR5IzIArnPUWl5CUDt50
drVwoARSNr4fUgBvIARlkYp3tIq9hbz7WEm/MsxiXpd6nZbn3uSJT2Tpz1yx/eAhcNQJIGr57jHn
ZuXXmLothGRk8GOsorFfqb88e3lldeee/9DXU0Rj99SHcRk3z0mXJXLPnMn8vHWCsysbS3WwE162
UERtraqHO2JGmhUX4MnV26//9RC8ENumPJlMlpNzbXS36XJZsUmtAQ3rtcC7dAc8nnLCVJpavlTn
MtTodMtvjAcV28XkBhO7aZQCvnB87HcYujeDcM7q57G/M961JEFTxIILHQgkohrenBOemx8vkV3x
nAdwTELsDZLuNGKW7jWG4Vo0hQMROcPkkBZe7+iDsZESVe6DKp0JEh0qnI7PGlZuUqS7ofFnFJYb
Q/ZEIXihb6Wg4aymQw3MaTepCGIBu9nCwIiMbS+SCcHeNoWlmhT5zkrnzpggE8RhhEHY1a53/0+i
f3pRoAkWuX/l8Xe8h8m1q2ENiFlM72RDkiyA2oJAbCgHhyhJVeVhoI/ylAhbTFCNbYK7780iMie5
q8jB1TwLUlId4wQNAf12UlVtXu5vgDCEZHk/qS/fwRSlAab5HEYclPKfZH7uGICiIrhs83/dX2Ej
dQNVQqUeq8xfh/ojBmuwFq/y71lER9MfSoAH+MUW9qyEuT9OWKCJHzU85XciQxm1DXwEYmjah+Dj
bIJh7VWOgSZJ+RJ///0Ki0+2k7u9MjqGKRwhAFw97zaX1OfsHGP8OJvdTLIPxzgw0yQw150iE73y
C7bsiNSA3zzuTxC3JlgM3/81rImmJqLZKpc5+PFRHjlp2JTMrJvDxVr7WtVWA8SXbJjQKZyNVbm+
MM/MrTnmAlj4T+MR6FIooCJX2YSpfXRIdmxLjigdWxfL++c6zVWJlKknwQdSbKq6Tk+MtdRftKBw
ad9hVHbfgBQZCpY6eoNmTA6iTfJ4Rb9jI5o8f1yKCgiP1e8kunQPxsidxKlLbBDKgz/Pg0ESgYiQ
hKpJ/PUZUy+/0+Q8PL9OHXgFBQvgWdKT1For+kiCrQE23a4/OBZ+nT0K6tZ+bTKIFaViZAhiZ7eX
WZn3kil9SjX3uzp/e3o2GHeo2f2Hu+/9dEIgf3UQpG65czeaB1Vhnkyc7685VA82E//uxkZhHU2Z
dBodXQ74yJIqZHCq57HTvwAU20RFC1jRLlt2ZvQU3R+ZqL98NrAOYPjrJKFDZxMIoNMjJ7TNwcZL
XejU0/0NHD6Llv+hTcQX8x86OxhdUoJ8kEKJu9CMImV6H2EhvdWEkY8EsMwuPJY2wwL5Ud8nxvjW
74EuUVx3bl95QuwI6X8HOGvDcRSbsZQ83FLROVdSnxxYY2t13ecx999rFT0qSu6vufhzAHSxFUJ+
Cdm3IsG3PgqdaB9uVGtkRDB761v/hP2k4mepdnrg24s0o2QhImAZ1614bj3OBaQkQvxXxysBRQE1
/NSmK9+vumVOoifGVh1JsboxAziEcru4fb5klLHXhu8WnpTuXRXQNGPfB0wTRh9cWP45hpBg8uPm
DmcCuLet3kczzC0rciCFqMLq/qhPhLfj8awb6eADkvbUjyDx48KeDMoZA4PmJZHARDy3KrgQR8eI
XjCfFIOj3aIocjyQqBILaBzIlJeXmZhcjT3QAo4WLuVsHVl65sVC7mAjr7zFC4fe+oU3V3lqJSVo
yb/+hjPnVkuqNuCVkTejswmvsfiRST9ALr8+mP644KGjc/JFJvzBQCV01fZb/3xyHDgZVzsEcaDT
Vqq3uI66ZccL3Q8IKKvrEguS+A+2aVYWaOEqHLSFLo972yqW9B0ACub/oiG7JoOIA5F81cyWp+O0
uZABFGPq1OCsRHtmd3AkwzEEOE32rYQW3L+F2PJD8Y22hO2pd9NhXAK9zNVGFgpbsnydYzH7AdZX
9C5Kyj8CT3dqGjo3hYNPISEnEwOdlD+bhkZcAXStL1l4HP3CPPONvnkUclR47eUdX+r4VPgNPtzE
Q/zNxC8QZ1spfpO9Yc6ObQ4hZ+VAdw8vMCTlIzYbD/j8Pr904EJ44r5tB/LZtgLRJgh2AsowZdqf
KJ5BCb9CO930WJiuqZRdhvpFMmgfGn0U/SIg9KigzNtnfLgen5ulcJbGHyxOxCTyfrbczkyRHT4M
+XuE9Xi0kH3mxJkMRlCQ5B//yboMZu2nnknMPBZxlssaT2ZKPwEnaG0t0H/osCYZcxDBEnMhu6ZM
H6bBvJZeKunl05or4j/H/LEdCakunBtjWBmkV32oCteyvbcgqnXl3rIPrrgMS3VbleTxpoRhutXx
vsw/efSrDWzU+qAPRDxnl6FdNX0ILfH4sv+SzpCBK0BT89SEvzSURtLaBIvI9EL0SNzIUO/2qFSI
ofO9SBrpcWRgZIdXqoh3UrfogLLlqcGmlgWIZfolEkwxVtNH6/3CzdONvfU7/RpD4fwHIROG7IjV
WaPwsbozYIod0qSyqvuXmBeZUlkuaTD3iWy+afcmHMqg6Q/tAGY1lJCtTgCCnyRnJjzVEREg+6HE
JbzfEtAj3sXQu7PHjtRJLhJSoPDy1Ty3XB+ZsRknMWbwlMtkJDwBUoAl9hcdQ4dOQixVvCj8mcz7
Zh8tg7e/8heZZb3n0TjcGUzLH55/et5R90XZ7p4F3L7RLf+BRaQc0BLn4dB7qNAtUHZRS9SRXuIA
X6hx3QjGpyIVVB17n2oFuJkuxNf8tRP1VKJIFYorabimfRyx9LHLtYmDJZXswtge1OnkGjakB2Mx
kyKnA2N2jp3eTf1faHytUVoP+hV7pVAba2ckVm7moyoYMG3YqruNo+282+iOSj5kbSjnVq/ulWr0
gCLSo1xJkBxT1VVDqSKWxU21HqjYjX7ZwP/p19jXuaDVDTlJUzQpgWswjXEWvWaitrmDtXzjbmp/
tLH/aqYeufFXEzD3HZu/K/B8S3aQW6LgPpCaeG7o5PPX++5jsfya2tkbDoOwzQdvqso9cGFx/x3O
ObVrbWdG5oDS05UinuoBYxLOspTiGI/bscLGrTbQ5ruhFMn7PFNqUCyq2DAU04I0s82Jf6Lvo826
mHZAzRrJsBpONIDW9oCntMNQZVp0K6smoF9rxYZgp9+pa7ck/x7eTDTL/cY8qJ3IYOZXVmILhFCf
T6tKkhhMrn7xkwjprJ+2b05YNf0jtW3jWFZn+cTYGe1DD0voLF7SwqZ5EUgWf6IVXX6ngj5N68jR
cMuOhs9+1W7C/YWy5IAuixWWUBBqWycbYC/Uwlt0qciZL2B4PqbfXuQr7s+BrgZbJsgsoUtZ3G8I
ljSeDxdO/HqK45A3LG13TRiL5h5BFJ5QSpvXIncizuMGkcgeyOxRXOyZlPQKc0HhMLf0rLHHoq+2
d8nIAaLT7wnYGg+lqqHxn+EqDDpOo6nvbLJ8Jc22t3NdQLTiu516UVxunywu75tkv1jatXjfUMKC
KMHL+S1qgHQNnmxppRTfqV5Y57KNOp+D8DwJqw8P01tiQqnuJLH35Cma25c80yxouevT40S+wAMO
3Suv3o+l87Pg2VxMD4BtWxd45Qiy5aMRupXyfYyQycrowzMBiNjiBFmbV6CtndlKBm6iQUf+3XoX
UJj01h087sRkhJHK+ydu4fjfNx5FsA9G5hVbQOyKX/nC0+uo8WWHyKzAQ7IAutYDsPKBaPe9fiaw
l4d3kBUx7kmeorrZ7yYGuHfri5stPbVM0wrdHunZdmIWtIz/c+r0pFjsMqg56jhK0ZyJr8Y2iTKF
HvT2LDPZiYvi0hFk8nO3QpIovq3VbX5dSrZQQiN1OzruIgcirReS+MA3KtCkBMrTC0kE1hganevw
cPS3Ylov1J5+dPQXTVrPtgkIAhq1B0hgj9UFC9ejVyojOX5NW73MbrK+QbdkjQL5R55M76HBsbbz
gGDLASfpFZCmuGLKK4yeIaZuxd/wVPGG6+PZuuvTL2f1T3YWJ5a2HAULEx8VxKqUX0JXVTmiDBxc
1407AHNxqpkjE4U/5LhArJuuGJwUAN1axA9SZYT5r9yrGnKpuoY/m7a8r/cMxaBTubwHd+TgyDGD
FzepsvtaG6dyfq5MZKuuwwJWkX8afS0Pr2iYDA16s0OROu7aUP8IH/nls3BdCQsbmryLObdBpPRo
nn7+cS/RgVljVPy6o8eEJjYthJE2Km1d2PSKyvMta9A9AJFiyzwZgr9hfxqnfID6IzEK1wUiv6x5
7zZ6ssn1Y8s4u0csrZ80/X7WNb1ta3uS9C3PNcAux6coXziRhxT/++ZRO2PWxuKwjVetdRdP9xSz
B1/5hh3PvkAj9WnVldT9TmrHPwhojqwPiUoO541eSB5OLxAMwAOvKt46omqpXrNNZ4m/TFy9IvkP
+PLSJRis6OXujW82Qb8mkPeN68N9lpRnl5dGaVzYj2DyEIBD+5HH9++PxunARZTxbWxzDIr2LTFo
vIaxuuQbWjW/V6a4nNnw7wby3Tdu7UOqLxCvv0s2eQGkg7miYqYA7KlRiw4dTv9XQIMZ0W91dfCo
6r9jDbcdrfGczuUP7bRfkBVBUJiWMDhV+r2HkL4JNVOFi33MLcXtg/hpBOOYerztUi5J/eQq4ySR
IChhkJZwFNtKGjTwFXOVVmI4/PvtpP1UXa/gdWXDepcKK8beysZayajRhVmgNY2Z9t6x+BEfsY2n
JXP8n5zU+j+BBh1ww/l3Qw1bBWGh+jJunA59u2HK8K7LWD0niExUtzgTzxXO5gCu8hS/ergMz25A
5xCm9CwK6JVQSTZTLkgJh0E//ORgjV/jmnFqacWKgNgaYogB5MtToDGfkitJGW4kJYQ4wV+GeAdW
lCXrNPrn2iBjrLTgEjob30CoVYH7tPsPtGtMoB/v1qAuwGnobPUEkikj5jc2DiljvWEp/NTr6a6w
ejxrKUvhr4jqaXIsou/3e+hewBJIbmsgTr4mWjDvXSilpSiR+iPgoDM+rWFk2oDX/LgGVbxDM1wJ
wNuacsxcOhIB9JEc8/Bbex5l07wwKy5kW1sKoUAF6vYBJbLpmiE5oNhMsDmCA1y4ixrrkaN8ENVQ
/V5YKdm5H3W3VVaohPfV6ytlY9im9KbqkrqLo1WygbBj73GPvlhyjf0BH80tf82PSEIisn/Tane3
z+c+Dws9LtD2UyguViJOBC7h8Q/RwMxrA0D+qHzLYb83Js3Jp460c3a2fGG2kDYKvmwVBzoAJo9D
6u0l2vop6udIRNkgIzG/hl8kppLhaodzezOLbzmhBjsivvjEweznVDeySogpWY0ZjO609XFl2vfB
7m0xAv0GlBTJvQgUBc+KhuQcif0ObyJJilcCHgW1MPYi5wFFl2h8VZm9cq4xNfD+KFQCzyCWK7lF
w8wZs83H7VCOfIo47cPfZGnZRA3HqF0Iia6FiGGuCDyG1snmLStSDCulWSV7Wgyu9Tyc5+HcEZvb
jDCFIwJGYVgd+jX1mdt4rurBhVzzT9B2nBXz5nN23g5HXS41ztVjncXhoxmWqhXsO+axMGs4iZd4
gJONKUdHHeK/5pHpe+XkbJ5nejy3NXUJr3Z0cLrFc0ZHaBWJCCUs8fS82agUP1OjUJU601tbZZE0
0vpGD8ny/B5+pWhqvbqo9qmweCM4OWWBQGos7/vScPuHm8/amublJiMV3CEx9C5bbAlGRgHbEKaN
vOw3SAV+64osEuYN59FBiusqrVsJc99qSgXPfC+AIQFP5cQqHngjPvsMCruXL34krJk4OsPb4+yk
UNnYS+T6XsWLvR07cI6Dm0LiL1CKk0CdA4CNhKAh+5oKSpnU5sHKYeAavMw6uQSsa+5WN+yWFSWA
Whbx6x46e4LiQI3gUAzPJl7FKojrcvPhIUD8nEwwBc4bLuABDLNtlIcKPOsOlqQN3QVpWPFgrI1j
1zcw2gmimMkTWQ45oe02AK/0plXFWdKjjfIQMlifdlWHY7ozlTU9MotkjLGnApqAaiKeK9xyvWP3
B99nh7X0dFnj33JDGcibzBk2q7hjuD/iLdVNNBhoTcjOxu0olbeN32lefH0imP5JC7mpf+3uD1mG
uVB5Yz2/+cSp/hi9ns9lS55WZvARWMIoxH1lnO6bQ/7G5wq7X2HZ7U84c3058Xp84qNPlIINiSQm
JjDGiyk1fCMcXHWog0jprwMfIWSeI/pBdDLiIWq2A0n//MhbbDJ2UrPJb8HBv2s7gXP5NcF1Oq41
UG0ZOnU28ZPUxp6V0bf2KPvdSvW5/PzndT24g51a2ZMvnupi2iXMGS7Bv5CGfv6uGcUF8XfG+cna
837ifVU0dPv+rP27xZi2GommF1QPNjZrFpbDfNi34oMXBkPnc91BB/skPXPUGbbt4PHEKxvL5KnP
F8HfMwBpCL34ZBJ3R3kMr78p8pIUiDLUyBxV1FCL767gQb2paSrNFthGYmhtT0xu5gnlQR1X2+hk
RrV6NpPxAkNMknOfIMppQf2oL4RIjCFFh1SIClg88lPhXPPwy+9FWuS7/b72hi2d/I9L+POsiiPR
xTBXh98WuujQsU3euLFS7W4UnHhG8ZqzrBIE1mxLcSq3vegQj4pghiRYhCTdRkNNQhOZ2BFkvjqj
6tR1WyE9EOcnC9ZqTAFcWgYGflQqoRlFJ/MpwkFzs7imNVO8gTjfd9oU0lYLGYccsYGPP2YPON4x
ZH8Q60KWbCu9+96f+WEBiHwRfGBl1bfvqlBoR1EYGt0sCNRN95cLlHCb1x2JZwlKhdzO5UZnYmaT
T6SU+ya67ejg5jdOGwSh522ONN02A6Vb2KiTztq9df41nWLvK0M8JNPTfheFkS+9U3jNrYLg1+Qw
84O33JhuYHsFNKJ2of/2PQSpbFzoMJq0zmsD0/m79/johdHyShPnyAcWH9lG8JcIMb4Kv4MY3q3Y
0kma0ulFQEAC6Wo7qV+Z76TguXtd0NZz6arPULGoch3jNI1ezXuyNZ0acWUL+z6Lh+C5LNeU3WUK
DxhEXtRsqTMvs/qymQolk3jHyew7AHZfR+8l6K4HCuSQ2EUJ6q/6FjUOuMQYnye5LlMvd8IGceLu
0rVv1DCZkalbQcZL9DI7AuPgwSmkc7cMj7bl3AaHSl53DRYclooxQbjJKysCzX3TGLCUCS3AqDa2
ZFtLbZOJHkVZY/zzHnrlvyP1CEe4h4XZKuuyyB5RP+fn7Pp9id/vctdBPaysuW30qVkiDBTt5Mbd
sqiy0r86yitLqS6Cv32tUwp6eff4sQWdYawSzOphH82nHOsBvDwnDCVHhCNI9LliBFRlpPnPqWUP
Gue7p0BYDTk70e/QRM8U4Fzkd1AZHnvAitjB2rZvzuYdEtyv1E8zutMez9tR0EJOL8dWFl6bQFRY
4qQBr62UesS9M9r1bRKmCf42LbULVr1ofI9fkl48lEFJ66eqyfuLbBISHcwk7XwQLZVoZhPiWdEC
M2LLyIh2Y8dU21bGI5PYXEEzDv7ia3VWsJYTqv9YHDoUSjbNRF+bRBl7kN2n4A8fJJZtlDoYI70R
RgidpOQmP4cd3n7zLwr4547ql3HIecrYHCsreQwXqv5DQGQKxJ4xu1SnKTMqZvdnxBSAxbxrPp+T
55zWyzgV3YrzOHOfMIm64hEUr+0LzJA+KS4vrk4kzfOAc6n13d/wpkln2Pwk/LOmE6F4i7P+/zT9
qAlI6iCrmNrVdzNxXQmKyvbw85RcOpiXc8OK8NYKhyCCa++cTr+eocO8lRqFsy/f6/PLRu4DHNiN
4C7nYU0lZckSexYAYvyW1PN6svapBmT+45onFH2xpM0fbSBTMbw15Xi9oZtasSuXCKy5HemeCUeP
+Sv7B4tRIpzaxLwu7N9OgN/6tF779Zqwf/WdOqcZ6pASVEQsybZyKfeQi4PzFKHGcqfWv4qY4RNb
0O8gGQzC8p8tmWTO9kXIN3I+tJibkEVg/V1lvWN2nZa+Njz4WElbq8VxsaoAnVRGZajLDPmKmfiO
NUBXeodbEi8f91ZfOEOpgpe/82cVYMZxmdxY8kN3ltlVbQZyb/O5LFSLsznfSvvfwHZDgigS8CIs
OKwe99IzdSXJySQ8VG5MO26FWgKUcDMndbY/kOAaRyqELAM7myNKbndvtKMWIjx8JqMwWH+o7kST
fyezYlq8RbKWG5S8x9sSx9K6TICqbnIOYMhVDQWxKMKKZG0EnaqP47BusoNVgakNJlPOHA6U/sGy
iP+xlbAGuwKzD8ljaVUoJqHbqo+aMHkM0o5GmlL52fj6oi3AnhJ6qaF/aYoGaz2bLuzqZXE0VjOE
2hProJTtHOZz0evyniDB9rVoorCLwd09KJfXfrsYgPVvXe2I2cbnpFveHHitnsC0TfWsnjpvju82
kEjVPgHz1p1aTvH5B5/IuXOpEQiOT7QVpdKK80HrwAg1RjcASC0HoheuBjRgjMDG4EVN5QjdGYVf
6/JPqvNSxnVC480Snh68EFFaKvtfp01RUYI9GxLO1q2LJkqvtXkbsqzOMILnBxP9EyrmDGWeN0jA
CmqxpaL3EVB5pdQS+9B1s8pKZhU4dYbDZd0PjRDr98qwP1gQ9pDnaK0F+2xPKiMjxJoP8NuQRD/X
sGYPWFR7U0D5ckYaU0d4iw2T1n9opQ7vu7XVxXo5vuBK/bpzjuCsGK2IsE7TjhIN0jyvLQffEIg5
BqR4GrFJNDWR3BTBMZak3jgpEqEdMBGk6m3L9gSZ3FFCxYMi2fSY1YvmYRq6SulUwgAKa8H+3W8P
yQ9yJOv6oO1sFIosRLFJ5XAyOKtC2IcDj7cSGuEtUwonPpAgZbFRa7hO81NwjbnxwvcLWgTpSv3C
avlBFUlZVobYUnldrjrJbzZ8YAUuIMGyB2XKJ1h/8EygooU5xkNVA/4MUlGVy4lQu/guVyFZTWXK
FQyQArbo53kDXGTEkd6FLVreWCCe/7314MjMFEOIJHFPArg69gaRra6wIhJkvmB8KBPX04kYWTYQ
8QrAwpAPfMToQs69vKlNLDR7ukT+X0TfDcP1i/k5KrXZzj+pxES6+iCRRfqfm5x5izMI1LJWGnFn
j4ChkmbHn/9WIdYTXGCDYyxkBFnyIca2Lud5R7wE9dfEXtx+4gRqHsxKnBa0yP8wCujpTMKh3MU8
78y0Lka4MxfPMCKIXkQkcoEsafFb9FSBlXD1FwKAy5ffcqjqzjlVsG2x+0hAVnmgjak9nEXnNpnU
oO5nAR4upnZ4SaN3m6qWkwmE4/XqhRett4v3WAF8AwStQRUZ8x6NxD3UANybHO+Q04NGyw07RYCm
YsykiUpFdq3CaqBIRDb53WnDFrUfg2HwGmmM4U4fXUMQPIJZGOVioAyPynuy2TtZNqRiUE6NIOJo
YXg2DB/NbXYoWUM/bZRle+xC4sOfQtZ8v7ePtkwnxLswe4Weifa0PkHeKvMvZgX4lAydzKkncZ2q
w2lZ1521g0CuiyqcH/E1vgrQMCviEtA7xGUIpbjOYjseOGgdn9R0hp2JXtX7hY6naQT8y8gLi4jw
YoYIwZ7YibXvsbWWnsfEYzJS1+DMM0M1hXzXTLkVyIADsiU5pLqj23f3LiB+tcocscihfwBroHhJ
EYg/tjjasMA0+b09HLf5JmzyDMtGbHp/aQ82KOXheWqCPIIZAQId92YLdlRtjTyPs784ZnV12Up+
Q8/YbocOdwIMTG+wyAURZPHWHkt4ixWwOMVxRBG33xyUcjVoRGVum/67ocSzdeZL18CeuDOJ6vI8
uC++++3d6a0rHRronHe6zAkAweSTXLr9qVdM90NzNgOam6noMthYHSt92KhCKUitP8TPvoLQ6frr
ZCidRDcvtBay8MMbKGkUFyDDidtZZG3bLG1XsPqMZcoxmPsyrcI8HQnugo6oA2VkeqgZqq568u+7
zb01qPLqTSTXBzwC0kZRwEvwrNdXz0R/ibgJjTIUiEZB1RI9oLJDv56KGVXzrtZQB4yHCF+UsATR
3eTdNodrAFEcDDpU1MvkD2x3gFTUnVczMOP6gP2D25prNkVgZyuoUWNYm4TSxkKN4yKvnLq/oADf
rFXU2B1WFz4S1AzI+1IxckCFhqzMU7UHyhb+Ki/yoHfAM5/517143hdamwwQ1IgsdCLBW92BNOnx
cgadPi5ievZi1JVKHcmRH5mlrG4Wud4akDgdLqQTadHD87aGmOBH+OCo9FgTnAQOmObxZ2sL4OjN
ddoR+9EOgmUj6Zt5ezQAwQSeAxRVmyC9Y5TdKvnQnfO/i2C0pNrBuVscgISi3H7pIhcFv1alHOBV
r1Ie6vweX10eV7q78PUCOrPTAbHwAIfyxH+fUH8pj+l1FxU9GmDLs7K9moKWrwenJwUwgj3XnuGm
EQWrmCdrBoP+ySIeRLHMCzCD3Jno+LOV2NL+n/WAKveXLbsby1YZbg3Gb90Kfm1aPdBG8Pb89orH
yrXpv77WFH/KZM0q4jvQc20Mn9rVYv9kxMVLpQ4/b/BcYTDHHsvTGOoRlgLlINSH9CySWQt2K9yu
BZQeQrkyVoE3fKhNvA1xCaqGXambhPdhPPtDDnhZvFn1Mk3KdfYWOQDIWrmrz5TAhdHXmMKxVZvp
Llhr+nppSphnFaszFJoIb626gKr5AdGtg2vkxoAsT22HRQlew5lw/Rrm8J+NlV4hiBJs2OYv3C2c
gUuUNXB7rk0pQKEluFBOqTBqg0NB1/L/lDXt+S1byKXFH9UgVg4YhIYLo73d0EWNDLEPjQ99HpsA
tBdXlsDiZ3dA4Q9fgG8IylkvJwSFeoGL3/bBYXoItaM7swzb07J0fc35Uk141ANayt7wuXVIClaq
XfpON5sTa2TimnOL0/a4FHAxAdeT0yiOrpWRBiAb0xM6dj76lLi0Iod0+BWHMXdXGw6GBlOiD6jW
4zHKdZcoW39kVGoHB5sw091EompkVabZZtSLUov3nRuXEeqpar8d+nyt8tbtMyCVfnyC3YGkcusZ
cUVE1ro42clqo43+yL2V8XPIcD75qN706fXQ2wKpadgXTIe3TRNNGQNU5oUoSvL+5f93TtxpIxvi
YxEzaibjO/lHQvC6eLZH3GA4lpyy963dwPlqIZO7Ddm10IPhfiPuDu28CdGJCvT+hhTTTAl1zSKA
iO8Yz7vekFlSyxIk3DkcvUcHfKXIoIS3m9Fr5KyBPVX6DDGV3bvHkKET26mz32iZ0fRo4k8RdUnF
unXuiKFCJLFaxv/uPDL29WN5enI71LBuNN7NV+0RHOMR4xtUuAe5OlkV0x/+NpszlBJl80hB9AMi
70yE4dNmOYHZXNjkQEG9OlQ26p453VqsArhndty/Q/rgeeuMF1DD2yuDtvDNoEwstGGOmAmD9FcR
puTlMiG6M/eN4KAter/j
`pragma protect end_protected
