`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47024)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT++8F4PPQq2cD1pLLMTjPTXpVh5mCVTmh7KwU2ZN0/MJ8djRxZ2MAZI3ohxDPoabMhhoKUk
AZEQ8hxqXAacXM7Sj0fRpcRRm5ExpbATJX1+P3Jn0/4wehMIszvxSswLCXgeRtQyCwv2KsmP7NUZ
GJZAAlVYnolFyxpYFvOeD1xcreDEwmzNaVBWYzPOy2HDbxkMLgZkSMdfna5uHO+D70S69yYb+6z8
uVUKcD9c0h7q11tSeyiD7rvwiWANrSoCfE2hNe0CCxjbNhtAYUTFRa64v8hgrFP7Bv4lnKTVX876
5zs0u6L1oO4fe+l6TsK09GV9PmG05sOBJmkSR5ZpiRJPyiPiSbUM8aQ10q0MNmi5KcdIKKnd1GFQ
+iR4gvI7XxAtPkypdcM/5yi1GTtQ3T6oLsjbjs6vGCGdBnKZaNXsIavBojK8Rf0b9mgAzDGyPKqA
+45W1Qw+JyXoq8J7hMbSU/fMrhn20cyUUxolDSbEDD3ZPV71BUiTTrpWnboXneZWMGdkdpNAVssY
PITM7kVGd5EJHPP0DUm6kgBOQ/2zPkF6tdocB6uUZ/xMGITChWl4XOPaCNSy3VCWWeHAdJPUaVaq
0sGqdxq/IOxGc3bT4FPCjX0dwyeIlSJQA0ljWtblryeboyo94rR/moeMS3j5F2EvQflN/0SdRx2D
f7DzZWwUYLqo4dE0eSSMdZ6q5TUoa6CqbXIoB6LDvJHvrMNmGYthOd53Xh6OkeilqG3nXTC+fHXg
KXNlkwGwk1x/8e2jVvLdu5lUSwjH5ro2ZbBmaGXalrHr9ZtuQ2nnu5jlZYndeOAYLGLk329z+9SU
d9LFiyijfbV/Feou1rz+SSYban1RUshTkzwkG2c22nwYhnwYDAWwAeo2kKW7U4cFlzlXe0ZCwmZx
zwUwMaOKTvWPOE4MyU6vmji0uAfVcVvDhNAf4u5+HoMpKg7Oeax59rbpX/8uuaM0w5zlLe58rchf
ZGCfMBtIo4iN6Yz4R1C+5BnV67v5c9AR18AZ88XeAvOCAl+miD0jDG7y61CDZ3b4HRO18n1gmhzt
v/ZmUvgoSftXM+Ez/MiMTrOQz6ouu352N5RcDxuGfup0s4Xa0rrKD+2QfLDSqGdCQeNwX13yJx24
Xxi5+0y7BHlsDvB9SqwySoJ/sOQnUqDzl3JQV16v6pNchArBdWJKaSdknOSbS5jxegH/M5cVVfWe
8DWRZ/xvhHgN8yjSiPXPrho25U4ne1BVD/BOIEC2Jc/uQs2n9smo2cFzQDUSqgtuWM6WrA4W/EIj
dmI3M+YxO1fRCWiL+dU2AeFENyp5vG4+78L6Zh9CTVKQc1h5fk5YL8XJs13N4WiTJJSsNXPRWjej
uRGnMm3+SjKrbgws0csNBYiIaVZniO+whGpJ1hSdf1Bun0KqQy9KjEKautMTZdjHvuRwj4acvr3V
Z+CXq5kP1xJjXY3y9654JzBPa1WoiB/5aWAxPJONQZ1KQnyS5QjS/gtfO1IiD5yr/N07b9lXWJuw
Os5Z0hEAMYLKSA7qTPKLcj3fVHnj1TPuWCHMZJqSiubv4fKuxHwslUBLD4/8hGqvCMkot2m3Ix6C
gid+09E7tqXNRxDIha+f3qw7YwhcaxluIBl6sNQrxjhi66sHhG6AJWi8hKEbDqN16yI88dY8gGBr
RG9oEK+wSj72HDIb3YaBQ47MKxk/lJ+0dttxlazUEYEMm5MMkdOQNt/8U/t5IfBAahCdClqBdPTG
oicTu8DRCxt3jNlV1Vqq5yudjIH07i2M0ijMOjgNm7Tsb/50ykqV4Lj/SnikPlhrZvEPYGxRYpjq
VDm6xNWeahVZSPfvhfVVZtfInW/1LEfGp4hT6FtX0UtE905E101NxzwNAC+x3D2oLrrYOwih5oV8
ocw1tX62MFocyLi99HYBV9AzWA7gbI2wiw8NjSWhuPL37x+YAR1w2p3L5LwAEm8WKqffqZaurdNW
BmpGdIEcjO8/uFrvLLJjhJR10fZzgsEKvp5IplzOBcys+u/FIe9rzGBap94XDSIGUl4x2acVd4wM
V/GYXIBy8aBVW6tSusH//M9qSsNNspxUriXDORptO0VzByp3o4+5EWcVxPPoOr2vHvA8Z9Advvze
3Uxe09OeUUDq3ravwhOFTvIax+IzTni7KG9Dr/2g7565RRuiH5Hw2AaCa3vS7HvBKmzqB8UojRF4
5K6mm1Vxun2JVCNXqdDUu7BIl+YBwhpN5kmqpMDF3KtD3QgTXRq1n3M6xWBcXME1TmsSNyizmwlm
pLmwD74gV3noMvr9Erk/Te9kKXqTOz17RpYabomM1fW3+CtlRG0iyTi2kLyKwyVOOpJfc4XoJ5rG
eZppRBiae4PbPQIMPjAHbi1e7NRjdJNaVSd41fW60rvDwYDtTLkX5GO77N72vIWQHxmsGS1uhL7R
Zmj5y7OLXWTEHRV6lXShTJgKWG2LPDIttavU/5YWGg9Z9gNb3V/qggNCsE6rZg51ukLv7E0GlL1g
20geqY6Ckbf8I4Zg7Dbs/+hkPyOy5CGcRco8DJSfY5H1M54uS13CnzidZExHThNbyhtivKlDy0MM
phRzU7zAVzbb0oDJ92+dMlYc9H3NIVQtI2mMVmkURgbvhGStYlPc2M+lcHo2UkiEfHHp7GjhJWpy
QpOlPaGlKJ71zaRaNqmIUceKe4mPvHcMLjGaWu2I+OBvgPK4Y1hWHPUaITySTqXBt3/zylHIRGjj
SqpWktwU/XF9U/O4DFz++M95XNTq+f1+lvXlh/6+Sbv5wYpaz8qeW/ZyWp9oKGFLF7f6NtjrIdFU
Xmu8ce3xhokbpNHhUPE+gwAa+8pPsC3REGo7yVCSw6Ps9Cof1rgGluyX+5Vo4pzWP7vejnC2d3AB
SOWK61AavJcxuLSzvEeFNA7U66Py6XqT9Vk1NJOw9ZazcsxMlKzOe+Bg/AH3aVgQPb0uiaMSGXpl
9v4WYs7wikyMdXrapark15kJTqkPZhIs6t5DXb6DDzftkhMnSW/1Tr1eElPa1K4tfrZ7OFDdT1r2
30i/i60IISrcLoe/xXIdN7gqkKYfrEaHsyfj6aX/UjhstJ+B7Iv7JMIFb+HuxvPTNYcLtIb3+qvY
3017wXx0SpN22vANnpGAk1AETRQZjidEYLd+tNEV6i6zMdz+8WCFMJiMxVxJJGQzfnkoYESYqP23
hCPU7gdRVBDQbYwLJxpJFyMTtoZFVgMGU48fejLm79MtyssQseCb7RYb1Q631v7mc9SC8CF6HbRQ
R5p6owHDqA7djQv75YWe/HvG5jWjgiW9jgzMjR8oPQ6YoWT/OMoYhDOiuZlm79eHDfY5V0Wu7Rwn
kbBi1haqcHznCAdqliCpENCcYJ2ITspN8AU+T8sjU4059Z0P9vXlu0zpx7Pu3blQiT5HxOMBRpU2
5s8AzH5nCYIHfS538H5TDMFIwAQiXl6sFqWKsnLB+jUDek/XqViiMn3yFOj8qFLTiroR1MiY8QQe
YuzjLC/KvINJaVzJCMUE0lpbaDIXwVFVVCO85vdFlOy1TyshZVEQTwQtaxV83d9YkE5WQ1hggykr
/PiTasVuutEDMDFhzW7n3atDl/eRk471Y6mNpMI/oT4WpIy4p1jf2PAJX3ibaa8/VSCDEsUaovSE
Kof8Yr3zk+I76w7T3lRhfnDlJgwEEwRjmFMfaXJFRjZEFK3qtvhAIjNF09TZnrsi41MERscWPBf3
jt9q/rtYmHStY4mR34BSr3j5n11NGRkC+qFK/iaYi3YfgoBTnyS0croHLoOm2OKotY7/pU2kqQoy
K1Y+OeHaeIqiUC2GdvCtg0xBwMDEZ5RaPQy1w9qt8FGeBh00xOd2xG+XlO+8Kw/hnDfkTDfxdZCs
KD/EjBUz8Q9mhQuMMeGCDEWB6F0RL2CZ+8abSSX+/jg9J+4Pbp+xNJJxwL06tEI5EdTKxvAKiPc1
uJz3iIdjjvzVvwWlaUSRze2B31jkm2aGrJI8XOyyBdsgvzTkfd5rzQ6PEp5Kx59eRmznxnLYk5Gf
qT936HbT56GvHRaGiMTseK10ULE9ukKcjfKEo7iUwghM9bWPq6XDV/+PmhDWll+LNMBjg67FzZbj
MczKx9hNQcqnakfL5VDMBo2Bk4iE1O9xFp6t44STS5Nft9olPHDS/kXIAUlnj9bWEixAjF9fPgyl
0VVWtCgHhh5RQgyBgSnPSo1lOwmr/53ibxWmX1MZYo1gDvwmFAsBd0QuoikTolpMPhs7iDMAR3Vi
ej2av8kLq6v+M36lsnpC/0oG/YzY34KBRzZ7vUtuTQtuGjFan/eiOrBfxX5GQPEHhm2IMFjwdAuh
sEzwWdIMiIgV58vIC+wzR9e58pj12kK4W7Q7vQRQtCZbOav9Ayo9aFoJK0WxUxVt1Uh2qt75syUj
wbG1LuI+bWb4JRpfeRG7Wgp0tsUpsw0XcluNBBdCdbetMWbqqxiA3mRdZfsh9lTAmtqijhsh0Re8
G89FVxtIrTl2CuecZ5hoF5J/FkaWq+tEYqK84lVU4tys7ygklyOOaCGH0BWcfFP73f9G+Ok3VLNT
jrE6WgFxp73mIhCDDnWXSLOeh8AByx0X3oAySJy7EFAtMP3fXiqQBDfjJ1e8P1D/piSwvGseiRJk
7OescUXBTFBMr74KJX0UWVXD/xfu46oI4VmghVkZomeMURrfhUqKDOAqO1KkRpc4tDNq4PNN/Cih
PkP2LIRBJ7gvBCuuhISMVcwhDe5PO6tFNEbzwu62YP5AQOGTeqE6v0bGbzA69IgRBb4sMBuTCfVb
XJ0+qlsI4yxyAf0AKH2SagQCsNQYqewmZrNlrmqfGHLP6Vl7DEjdHzEhT79912Alau1gyoCXbGZw
ex/oPgF8Ir12nyk4PALJHgTAhwXXaytP9jzO3uV2pg83+OUOPw/95tA5OP9RJytLGdSwUfkM2ejO
xxdo9KbddJd+08jwYvbEN5+HxuhPyAM1fk7TNRgwWI/bWkzPyvjo4zNxg5NwQY9qgfbXpepmoRSC
OGUK1wIorVuF6jFpJqBUhcSD/zLgS/3sC1uA1ATFM0TH3A2DMQKHc5fBCykTF/UTnqIvO1K9PKeR
XgmjtLvWHpghelMjea1YW4FYC9D6mox4RbjYQvFssLlCn6THZr9qFErHYSIFHFD6PFOI1o5C2FdG
VeCQxXW5bb+Ld7fYWnsH87aMIfEsY4zVqG49cGdmrp8lgYEumMM6W1dXVbRAalOTtZxJoWWKhkd0
TmlZ3tH9NOxRbvOE6B5ZJvKD28ayOSvfm9JxE7y4gOiYBNnSCI+AoVP/Iskrug9Ll+xVlYiwo0GN
sPv5e0BfYYuND64egNdsi/cirILlM1/Im/Gzaa4CcbMxGRNVq8K6sQ9cmrjx66ng1IO9zN8kBoO9
JmY1S82VFbPxiQKW3pKtRYL9bjxT2lOOPUa/bxgVOBZMLhv6sSAaheC6KryD+GTj+Wg5nsGpvs0B
BzaSanDyX+W9Ut26BBuvvdqyQTcUmWVmBlKJQgcExNsqcU18nfoEqjuApZrB026Rcx74rNwTObaM
CPSEahyOC/QKts4G3mPQ65u3fkLBbByLDEZ/dWOeUTL0cYlOooXQqSAhgnijCMW5uIRvOCLiBzUF
50isxCImw/4Ec14fRgO9KJ2Iaie4FA2sLRrqqHY0o0vnjaSAThDNNddkmJHLwAT/RQZIcL+pwl2g
QIcnYI6Gsc1YfTP9DBife/BlzswMGITNmt2ZRBL/s6NpPdtnEj/LsWfT0nEI8rmSwRLV/maN8K21
0id7mKDS3CFprcwscpazbkP7k1aVa04NMKVvn3h0NFpYWmwxRPJ5h8A2ZMjloamcKaFCdxzW2gho
dBLFVtdo1n3OZ378cT30DQ74gwVqn/Lro+jK1Z+Jv/dmcmGQ6WHazRFAHhur4l1f5aCOsFsFfURY
+PpIDupM5DMUZpqD2dG/i5wTheTL6aKwQMeDeeZFMOR7sH3BImzckpaaeuKkrk55NRoejg/svjr2
9+/z5QwkBh7og3FnEV/smYXR1c1w3gGdVMTq9lvzGaWLab+OZy+1Aswen+r6w9dnn+9ven2CpwiL
M7iJYyoi4tMV3b5TbxDOsGOkM7MmA0L7ak0BAQga2v0NxklUcEQPp3PZZ8tYso46gD2K7hH5f6fk
7dlYqvZ/gLu3JgANlcSMGmoH255YeIONKlU8S7O5EMFIhIE/YlftivUIcuCEzP3OJydwuqXEOVhL
uoUFS2TeT2p3xMxQ78M11huV/A2ydCw2PenCrmL+aFZWkLlDh99A7qSk3sGQzQdIcHj1flxpzwhM
I8iqrKivcHMsGQn4zCBqTypAuWCVYogMfTkbTqsROt5fCtH8qDQbcn+V26iYAtAHKoLfxzArS3PQ
rF55Oiv22y0V4JfNksFMzTwVZLoUSXoDz6WtyblHRuEJlTtQRSBllhTffxj0/yAPLQUm14OpIyvT
/2GEnXeR0FuHHmRE5L1qxLdabu96Ok7n1SGGlDgeZvn2lwLx+n8kYviCd3RvXx+OD6C9MSGKuZTD
rz0ejrmyfd9AiDndA9DPdW0IC4ia8cOyDHdaZoj2Q9c5+a8mgxSBcK9aaljvA7RbREs4mvkh07y/
R2RdW1Qke1bc7DVPHnnRKTiJOQfHnhORxW20QmUK6S//k3YtOV+AZa5Wfnz4IB2pcVVTY1lhOcvs
3GHfF0Uj9wuFqtKHi3eScPQRnn6lvH2W6tKd6mkVHJbRC0vdTgectUs7G6GsjuA3lDrxm8aVB1TD
7yQx4nE7crD3KYBnW/LSaDMoMdqdskoj4uJna98DqIool6r9wlLDGtfCRpGezcxYUDsdTWEb95ch
1cm8h/6GqQI2n9Ww9JbUhbNu5GShro77F2lRYg8zbYVmHxiOKcaYWhytxjGSgP8rJ+vTnu/DbPgJ
v3OKmUxkI0/IIvwuCXO2mrTLt45sn8KKF+B50EsiPqgwk5TK94ArHai9TbFA9YLICK+Bnnw6MPwM
Uo577ipVWq32Y6WQDdjA5rxvVWSw7It6xnL/WWdXh7T7H/Um2fSD6vIbSqlP8fzaliIUVR0kq9YG
O+u13WWbtOPoYnZDrgOrYw2F8aouIsE377FYQSRaxkArx5nnAz87e0vqs5D6p+L/987g2blTFHXT
lBFqVPoRlLeRoRwW4DG5VGGecUTcrOmcC19TGSh8EKGs8/d5mxKuiG+GtS2B3QtfS+zR0DzcsEHf
owL1kChyAp9ucr9hPe28koqP8Fd+cFodm76ADUig19dkpClblKEASsECRV6/F7OBDwObHy3eMqoc
KXsHNOKggJEiD6kB+/iBNrjqt4GQMD1xV5HWIqZ9fEPMye4YqVQR+6Oe9MOy3QkScY167ueF6fhD
b4xOcibicXj5gGhrdeZda2w4wZ8px6mzzFfSuxn2UBGt8guvLOzA0LfhLd2MsI0f+JYzRuzmETTn
vQKfy+9bNISIqySxNUlnnpfjGCN/Q5qFuFDwwi+5dzJWjMiGorY8jsdFonGzCB9x0TUR8zwNHGEY
j6OJAGyzK7Uc5trU8Wew0ZQUTkNxUUIV2MKjA1JnZEi0r1evoxDeHmNZ73D88fd32iMaq/9xa1FT
/C1EzMYQBYAU9MIuJZVZViscCot54jdgcySoTmb7UOf32Uryj0ymgGhuJL6r54rvs0SAJfb/mQMY
UyaRsf6L/nBN4cOcOx+VFwMs72jkYWoYz+THIPqAWq2BWFOnneUPblynScwgWm8GEhh3uIIlgKEb
7vm7IdIBu7oXvh1C7fDJ43i20kbtFvrwVEgzaP4f7ixnYmhixMrdQTbqLMmXC/eNbBptLmZDfRO/
gOs0+kmbh3aLuvh4RcljGxpw04rhhQ57i2yyeJm0xk/MWfCvJVeuZSc6rTRLj3K44ywQMOJsVvo7
5QeHM0+//gWT8k/bYvITzYLa4a8RYxc0xPyvALUdh8ir+ZFj/6g4v+3AMdq5cm+VrPZOK8871nRr
6bDlU0nIW1y2sBmskpHdiXDDlvlXp5DMY/WE7QVY4/pRr8/NfJFfGCj7i9vccgGeKYLrtDH8uNFF
jeIjZjZ4TVSkfqmjcRMZFvThIy/eHAspo4RegRNJBe31n00CyL3gAHzrynrNAmdIYKVji+crji9l
SY0cUELTTjbcephMQuFAgUT0SalF/s3OpQgHqoVge0kVG5xLRfPT8Rp+lzzINPhYNftu8ILjrues
YiQGbOct1wwF80JieLbmwhePdOo8tdx8L7qFbuxVo1PTNDxUE49LmvK2n1QiDVshtFf8aC2/+ggy
tuR6c7+rlJYLP8IWrVsW/HVmw88ZTNsSqJgnWGJ0k1jmV0loga0L9Z7z44lVvntKblK6RwhICztP
PLK7JE2IrCKGp5RmAUjLFcKkvdcJfXys+d3urU3SG05zdesGn2tpA9IKuQ7VfDMrT1OKjr/oQxyP
xnZOPY/PwXCSmhcBiEzUsB9e2XfcdP2B0SBoujlUaeXrTCX0/65RU8YCwE75CBHl8djRsJYXVZHg
oVKjCJ+xuo7bX1crhIGgvpuxKPiRQ3jRreo4IGKZ1GJPKY1qkPAV0xf6WEIWeZK+r1PYM7kvog+I
CHfX+76qCy3fIBfUnQNDmI4q0fBs6U2BujNa/wVjINuYyJoS1ZZgsoViwscxDBO1PAAf4ffaUk0A
fDKrHgx7O0pkMRcAO8oxsKTSE9OzrPv5D+pyj4PcVcdB9zSpKz9UcAhiDoYaY+pyxvKfz5Lea4te
uxkqgQ96oxBNyOnxIrZx+j/WTseWpbtYToSiRHyQAzyRnFfJRG0Z5O5A0Kx3GHL+7TIl5lNtvYYL
AkTh8U9qKYty5GfnULidos1ynE2fYRIhs6PTPKrckmaqEXIRGh9/xUk0dR/brrzG65Hj83lnV5Nr
DXawRc8DQLW6ojCg083+IU54sBdUoqc+//mXpCyxnCPNOzdaWpDs/jfIEYvywXBgWgvbw+ExvLbE
j16k/3NvbwkCuwDrgUEP4swE9Cd+Eck3gQ0bV0pn5Rcv+L/doI7IxA2ai7wg0T2vaTLWwBkRyxlF
tndT+SAGLMUsZwExrgsvSLxvA1+mor8/xpEuPH8mXIi0hxIEP08GSFXCvBewFkutIYeTFKJVAsQW
Y9NpNRqB5GgwnoH04IXi+1J1lFsrMc8kIWia96jseGmAfA3ktjt2RhsgIdxGkjgtghYDxqP5TSK2
Sv8VAfceYIgZAFpPBp7mVR2u+PbqYo0OY/Quj7rZdCNL8tGowdHacmXtivd/EhxqAhaPHE3miWEc
OUXWT03F02q9ykaZVUpr9fs/OBtg0NgIcX/z01aert9OyTChngsRsWKu9aOBQ48C1uMqtwl720/z
7sdmb8EyrOqlpZNxFfE1/NckVk/yMHljvBlz3l3FX7xslJqyz99R2AOZZ1a/98zbpmZ8jeTYIE5G
M/+u4jRXQwr/e4nKzAPdPWAx/TQ+jjo0A4hkyO+q5dIC9Sz0uH9NFtE/3ufwfAPUBZldpIR0XzX2
GlW1+dyLtcSEKF40GX8CeTkILwJz6zdilxk3HhoqL7nlmjqOCLlvGqYH8OwMpX7V/+TEBp5z35nG
NcA3lsoyqHc2WuT/tpYH7Cdq89PL5Ur6OMkxtOyG0tMlkOpPUi7wBv3Vaig2vNJ3M721/MzDBuuS
eRFxHVxX4cDIEpMjp+dRs0s7vW6PCHAuDfcGC7wDfApt2FylOrnELxsYke8xe3JYruHQjlPoKOA3
5NJKaKmVwygj/MNwatGzRlkdRCvFrwM3dXvgkLw2011XWPPNublxbKPPVf9B/FqNxVsng23alANK
Kd8BKbDpZ6bmRUuV4yLCGwOARdJI2e3tgSYxDdQawSWrPMA3TLeDpaCz9RNigB0hmaJElzuGcxWp
/JQkFihTl+5vWArb412iV1QXcMT5zBCV3pG+P4hT+29+NcZAPZEhPGscu2lIQ40kG29nN4zR2JBC
z9Y/gGlnLkA4T/G5lCMq3Ke2pqxQoSCrA1lgYUH+Fx/GU5P/w4Xyjjp8+aJSU7DgC9mAaJ04Laad
hfRDWRvx1D6aFE8TVa51shmGlNBrkSk0b/pK+4UFkoMPXyKreoDhgxf+1fZvlKR9fDH3BRii1uyN
VuJPNILjLXvxu4kBF7W61fgICYgZ1g/bsJRVmGmp5iGhSn/JMjQ+GGecT+ZEXQ6pnmpWx64IJocq
jucX8acDMp9sqcQS9IBGDxGoYiQPAqsPD1H9fZ/z3Z2EJhnrvct1QMElJEGWpNWGXzHjUT09PRXy
ZkRMeybmD6B7G9N1sYnL2i3BllrwxRlp90PaW8eh3J+SEIKYkToCHtSjB5dDYFfb47JgtL6ocqQv
NHsRYIn6p3cBRavALJOQgP3/wwfptkdF1Y2oB7Ea0JPaqdlSbFOLRJ8pVEiBbbpNk7mqHa2yAXT9
elrBcBlpApOwRVOpI4UUeG8aAvuby07PqvP46A4oOdIo0d89yEIh57l3gBa4F1lkygLyRVo5MSp4
9IeVdpAiLTT2zhR0nfpm3KpUrxZUwWKXMi/U1aRrwK9sckX/L5IxT8Z+/n8xtMX02NQyal1GW6+F
gmuVGLImYjqQ0JuzPJy4ODj1nC8OuD+5xX7qzrYOgiPiz1hd1NsPwM95xhDOBxnj4es+DaTLH2+w
nF7cVcvkvj2yQCZrQKY8r/zobYr3pp/eVjAMpvRd8Tjqe7Se73jLZTbgnag85GR36StSh7HOQhLB
xjv8sqLlD7mDjJR4wAbc/IMrHS038LhV81kd4H2o6qygZ+vpt+KDCnK3zo+zYCWBOJmpWy0YgZNe
AGjNvWNL4P0hiCWSAew5y8rP+ZZNt6iISjS+uhipDEqA5J4wf5iBXnNlOajdhz/EieZwwTwkPTO6
Pt3iiu8ybQzy3qIR1Rno/6Pw8Ivct5bU3sX7CqJjWWEX9VrQTs2jLvsB0J/RWkeNGfEPe8K65xu1
Je1B4xUmlNVQZLqYHq7FUXhh+SgJL37XF/Nt/9yusQ6xXIahnSkV9/X5PNnCyRjHBWrWKTJ32q5+
7Om1ebPFM3konZy20n06igeKHMBi2FzfoQmui2DY0F92pD40t3PoOkYbjFa+N7hfuB+al160olJN
tn/jRlt8GN4rQWNc2l7YG+TOVcrGpPBZvPJ9g+k8CEMlOW6AffTck/qzSEDmV2Yue2SoCPMO0kX0
0024pd7yBauKxFZFeIxOgTKZFLoAX5vwx38uvQI4e1fxRiq7RzHVvxsRQDNiKRw9RF7nm5Klj0Tc
nT9rckG+Jv2jGcRuTTpn0raW36iwA8EB51NBMkAygKw/kBu6kW0ADjoxcjdPTBoZsnc0sn7jhKIu
JszAsQ8yNA0lFdgfU8Ywv4K54bQ/HVk8B1fRTZX+ZnMR3GbTqrzxTadN6BGvZ9oes7c070a1Dsls
vcD64fq7Sl0ws/TZ76WltuO0dHVzTxuubSHCSuEszJdtBM6qiys47mRdKyxaCKua4WwtbZa5ROkf
vsl7QiaKPeaDpmy9cFMlSWLfg27ee4xdewJIJMwU69tKFGKa5IFTYYEEp35/YvbkIITXbwYoZR0d
SCPs5Udorn9WLA+O80N8rT7M0Vebb9aevZDFEbMSZ2XASblDIydMto8RWqRGjZw10cNAvPBvhxm6
R4gvd8TGi5tkwXcZb5B5msQ0BEobSaSULSpT+XvjIaheTyWaKLBxYM52kcfKEv34TwkQxNgZu/CI
oWFYopYlyHW836xHXHdys9FqOSLYAbOS93oK7JYq7lVq1JtIIMip3XJ0AzUSzaULqjUrBCut9Xki
+kfHlEgpIeFPa9sAfjytYCExyLB3vTD6NCkmSxnt554YBMFp1JytcuoTfB4CMpLVq+wkpnz7qmSK
r0AaQXjPaG/4lNctG33gPD4QtQhl6Dl7FF7ot8pgljsm9Ks1KJwaAa3M+8tPcnDCxypDV8GoLnTo
2po4W1W6Ixy15xnvn6UL/RVe+TrAgVUm95mUPQGtC2CDJaRxDWDkPJbO/o51Qb6J+4wEXRcSI98+
m8OltadOBwsrQQI20WLEWnMc+Sr1CR0PPMzhSvYhLn+xkkRNXyOGGd6POuMkCRICJD3EAbqmXDOA
dJ7AUZlFCyLsA+QahBd1mOT++5WW7JTHott/MvJCdf4fSwkrRm76AzaETVKNqnS7ZfLwnxhwox6m
B+yuFDAvURGD+ctVFkANr9I1YmX/3HpVVK6QlrRgBVbGzetZV2h3KlbEvHRUOKu4pAoNtLgZNp8j
uyBxW6RB6zk/XpGwwajMiTM0RMTWKi+fMF5GqAPQqku+woSDAjZxXQQUGLQaMeqaTZTRxuY8+4BV
lA6IIOFgbDmQrwPWOVM1btbQP4HpNzBXcnBc7ofHJiETt9/jhXvSrVDn1B2xGqpbJmgPTcTn8TQe
hLh+4CUMTTxek3H19M31WUvfeky6zS+Kc2cuyPRZT8KNJ+4GiTBH+j01im0h/eJeZwwcMuX9dFnj
btEOBCWQ3ZACiUsLvJGohtzlMlnXG/almjnQ4t4DBHLJi54908EVPtbcSRG7k3+3Obp4FIiQxeHz
bgzduT2raHsSMjisoCR1G1o+jAg6igoafVXdLRfkc/cprf6PdjMg19lz7xNUDMuvKxemYTEpYM9y
7C+vg/2N8o9m6mlfm22pKKgo/btWlZUAJn6MvAuUtjbtuGm476lQbTG6dvbJAoU5nLzVUJb+3kXE
dZai22Qbn3BwmxGr0MYMu6d1vTzA9SGOFfl9t1vzZf76DxC3CaS6aKqKojxz78scnkdrLUL/H/lB
luFHCl3waD2sjA169qHsdM9iJCc3aDwNHmOFRdD3zWrV2VYS3Pdn0UCcmVvL82n+JuNVKEX4zIq9
/p80xeuWKfFp86GOX02F/AJUQzEfTTCnwHt7lTXJLxr02ZT94g+ATgYMfRZW9uTdN+XNlDUli4dQ
b29PfSDKNAjnVOqiFP9H1VH7Q0HryHNxLZKtwLctgLvWSvmJJG5Pn7n2YItDjU6v677S0CaPQr2b
4baKJDsA4VFxNA3m/JAB6zxwdlmGaKGS3IDIresN40GmGF3biKnTfd6I8kFhU0Wn4azeqpHMF/rO
3EmQsmwjHNm/DlreNy9dwSVLW5t97Qh69UBzxtgcTrNORtlt3cT3J4IsUlaZGXqoObgEd8ij0kN8
ZctN61JgCzSC/YLy9bTEaRkDzXSnpDCwiERxjZxVubjFADzVmprEE3iOiqFwMXkMkMS8UKT423Tm
RNlCAJm2pdeAw1MbNPIHqrLEqgno18w+JhKZkq1g3dO35pjLK685B1OIReVIsFRY7KDt6jO9RpAB
j5xLaEgdKNbjzyjiG1cJDbScrkKL9i1tuMLOqFQi4t2/jJcIzJOWYicxaoIAbkwdTLYdBrUDKu/L
xQQP2iatMLpve70/WDndDubVBRrs/3+Pr30krdelHvH3iJgcWhdA+/+k58pU1tlSoffhdvS8rZPZ
AdSQxe9/4T740Mdah0fL/muJcaugbH1Bw2sJ4jDtrE6OK0SwCqjXyAIjLlrfICw9Eoj5RMZ6P9Fs
5J/bMbQthNi6s6eKA7fOzyOaEu+BSJ1egftAYkvPCNzRh47LEWDMEFpjYdZEx6gCoe8mITgQxVSd
R//z/jxNHLxto1k+MOlagJCcvOEtRTgPBiD2Kijm7pnaC9SZGi694LYuh8PrBZ4E/j6PLFA2D6JB
yXLDN3YeFuL80KrLrHiskwtLk8/uFMjPgIiirUnZXLjed5Gn+oDmvpG6o149zyZ34NkcOgftNalM
wBhobpHDPOBcMRPNOi27X0vv8Ok8U4Nljb6/JmmCLXN1hjEGSaiZwtgczCtyJr5q/M4u8bOKsHuw
ls1yff/qsIATCHVTsS98RNt5/AiUWVU3ClK7rW8I3cTPlJam+jAvcPhgNU6lqimx5I1XgSVDE+hO
kZQQCVy/A89GzkXuEza1FKNnreVBab/KBVRyaq1Yq74Zv0kUutxKI9rC6y8D6vKpRmKeMbXX7bJv
UdS0XAh1jyv0ZMUMEHod3m4hYkg82qY68UwPKdoqs8x5ae8c/UiiUJfRbDGyYKZNF4UBSSsRB8fN
KPJLX9b5ImdxzzbtJ8o8vzWdXeyQQbzRTiz8dIHJOLmr9eOGCvNZRRzl8ArgmQRnohXy38Fyybli
roh1KIh3yca0QBDPJyRDXGz9W5Qgg0IkXLlZmmFPtziWRbvhfTvKHG9fT2uZ4zgUgpQepDyh2KzJ
qxwol2i+iO2ilQPFF6GWy0V2+XWKijqUyLPtpAihcB498HjfH/cQDY+tuQzQCrTvO9p9ip8mkCCD
UV2/3Ll76VuFenCi3QDoQrE9Z8+DznpwZTkzZUbosrvqeN17M5Dk3WPyMVQJAMkvrAjJiHloHw6s
vewJ4/ReOCyIVVASyz1Pp3FT71mg0yQwXUVuKRXUr7ph3tqwVYuQICMVOesWqgXL+cOSO44w+Zu2
dnZAFzvuhwem15EEywzytSimjXS39ZZfWqTLU/1DFEYMPJZy8UC+qvTZPR/ik5BhtkYXmrKlRdhp
YYOOKmO36tm6h8lqvcN4usCe/NkOuke3VWV2O0hYArMu5ZeXiD1V5BGXH0wT51gTCnVHmW3sumLL
EnODCGnZLsqvD1nwjsgp8pG5Ef/D78jbk/RTagNmFhgAH2QHEsY79lJ4KGGbeI52fHWb7LWhakE3
tIsY3ou1vJR6IXPFesUhDoxU0RFRF7HHjMdwWc+1Afv631+vsFOeaTEVgzDh8TLZum2A/pCooBGx
9o2I+re2Q3KI6eZX9D2GEq7ahgAiOZDkIXEJ9AFc0hYO/bbVXUCthF6otUSZprdeAtW18KKltkfP
qrV9owi0weG6+ETjdTBVZSZpv20fd+wUdWlV/MygwwKh0MpNltdvfxFD9cBOajwNSrM3NeWInlbS
/dKRaRAqc6suby99B/eufBiF1TkMkEtn+UFbTqAht1hWJlut6eUXtYF5K7RosNdSnI1t2oZ8TTlC
qX48tpoqMM4UKVMqzGX3Hf2m5Svt9xpLEi5jZmP1OOFn2dk/qJ55KuUJAqnwT4HVscwpa/7hMhMF
wsv6BntwCPIr2hdA9TzMC9zmyr6vrk1+ZIbMKaOkS65WG3VoApDF8idUypQ72A91Yx83i9BOedrV
JNbpOTiGCS8pc7q3te+iyZOxw1svKVKgeBeVpfEh9MGj3izprH90lOts+OkW3kneDJfP443kx0Kn
ATCaKfarm8pJRwAsulbvz0U67hjO/zqFJojozQDgvnEzhZ79rHf6M0/zlARGy1KGo2Sx5ZAjjIu0
FgyPMhiZHdW76hQcgbP7vU8GCtmvsqO40/rHeu+MSdLMRjf7NKA/4P3FZ08hTj+Fg6jWpq+FdKRx
bEBFeNuBvTWrLl46mcXIxqqG7JGMNitQcL3bLLaSrtAfnvSTQolIveKJXL27veNAs3eZ63Tk5eaT
1q7cZfQDIHCIGB6hjvCYJ3v2K/OdG/ge1l8vuRWsYDnztWpK3+xYIxaRdEKFU4nGmNFCQpQ1m2Uy
/XSEvH7Mn/afaH+LSWR4VTGmwT47WMfHc0V8W4JGatP+E7tkDsDeEpgbKEMCQ3+b6nbo3K6ggymM
mobNk53TIt7zVDN18J0+QHtVTC5zJeOaX/7WbeTS5HpVETJzQWa562OC1myyes2VqWR8eDqZ6x1U
cuQethRFXPbjP+m9NyHuGb1Gi0nzDiXIhsSkbdOs62EbY9QcpiyLBwvXVhfZw6GguZ+vZTc4O2ch
V0GHkPr6vwa3B++RNilO8GE170oztuKgRatt3ITHwoqORGo/HdFBj6pFq8WRl1n9+fIjbFMVf5PV
6TD+KpNZhBE1xlTKVdgFVkD2pSpiXVIgxpXVDzGB0uaf7+mLblWCr5Wz5BS4vm8isQ3K8SNjQvZb
5L1ZxCK7OWpAYxSfp5Yj8eQi9asCktOQ1C1OcVpekTqhuDGhuiYo9lxHpNh5RFfwiPMkz6WGffd/
RjZRh+0xUyDr+h0csDhvUqYSq2P0RGjjyJB4opggPoellt7eAkHy28zdVvruRi9YtlNCxlrV9UZS
1FlkVNK1w6rTvzAG4t97D5tSLCe0dk7apl8FK6oP66gOFvdELo5gi6xy9Ifo39CS2KorO93eXP5E
QP9lYFC7oWMqXfe7JgmWkPWDvRk/q8UlnjuF3UOVwAIe/ftwIYUq4fO0NHkN3VTui1A30LMpRjcb
6GpYImDnq+R2AJpweV+uCDOcNbgQHs+xwLsj1amSD5c+bBawZMQYdYb1AHxp1Xon08FWpQfeSMSl
G4CIaJTzy+ChxTYFBK3GgK1HQc050Kkyj3nDoOGh9ACux7uYqhBiPAjCV93mnIcV818JIDt9XHGg
a0GjgyzXPCBUswOJTzCditqyDt0Cr4up/HmEOCOPw6UEvs2EmV/hSX9fzfObBX10E8PM/omkGohl
v56EytFz5yfNKKzQxNRsZmP5UJdd8YnmIhhehnnl42Pz3OOeLSLu7JwHDpygZCCvFsW6WkKtEmkV
Rutp6SdYtxgswuPb6Kf+E6z/ktRXgvzjY/c9wqy3pue7dUa5sjVwUwkXVDDe4USC8HVmuiWIrZ9o
FLI2ZMAVspCPmMeCaZ2g/QgvVTngViCgjLGxeuBudrBmjxDRbUiXksvK05kwhwF943+L6nlKcfoF
yld5AX5yvwNAaNFpjMh+p40haZabvTFLrCZeFYJ5hImRQdo9QlGBy0QJDZzP0EQontJvV4Q+OiFL
KxhT10IogncC+jq4sKtB/B3GsGVJW1jOs3hB5EVeiHYp4pSRq8SfFzjcDrwO7015Y9Jg9M1yZrU0
upTC9o+sGF2gwTK6FpKYWCXmEu7+uOIiSJe6OXEtMmK5/LkPSIyMOxn6NDgsP7msgQ7AmoDskF1D
g9ryisBmyPCGaqBKrvsKNX3N5BO6j6GLORgV5CO/sTP8ej/qDgtiJdDyOYkjF+Uca74KYivmdu9H
AuoxwVZ5BMJNVq8paf9OAmbBIcQY49uk4Caq6QjTDamsnDWmfsKqeMRiY4s5bUnjskkZAyYX1/8i
dRyVY3gMaW7LnLUvd3FvIKeE4ciSEg+JIMVRX5XI//0may3CsH5AJ44K97X072tYMO+aEMOiKGqx
hBT18knu2ZYuy8XHo8bQzMpf1LqAJeGF53JCSrBgtKWHxi9C+9OJyOO/ZJi4fy414qzzZ47zqGOF
LkCh4nBpjYrj/i9EdZ5AHqQXF/a4aeGP+FhHpmZpOBgQhk3DVFnU6zs04N9lw8WtaN8K6gFCNvss
92xljVk1FdkXoymR2ncz+AZPuSCCaLiCMhwL7SFzbIAnHGytTmhtzaPtRcEQ1UX3LGQ6EuhHf/B6
OW/iypzXUrls8cAKp7mMR0f8p+Dc2G6J7nKAP45MRHmv803u/KfYT+SWBL+TH9xdjhP1UFIiwWTz
/U1BvPh507bJhzoDMfinsCfGg3iRSwUAcji3/Q4TFgYyaPUaiC3twqP3wy3gt90YFdQLfYMOFQWt
nB8JL95l1cx49a1bKqTtlxqAASRqqCZ2YP34+B3HThDUWXObI2EDulXwKCcFdR0PNsgVfIgzMBlL
Pyl/vitQepwm/e41LWbDhf6p9GFKjANFrqETL6e+IzeDbnhbbeIjMQO7+ulA5AnbjJgCeB96mPqZ
967SS3DKS7uIfCvmrFDI9LdIevr31v0DCx2Jk31xK45DObZPQk3Z/j5cjovHVQLCdCLRmbPtddPF
747yFOBgW2vRPiYIs5aQQZLuXDn680OyOSqJ88M+8gyW4Ddl5ylI9u4buGdx7rv6WiJtiexGt2xq
ThZAuIFWE5E+CbR9c71ioxwnrPCyloUObVeNUUwjfU9VXN2gcvAbwh5TIzkZeqZPOIbpmf1t2c8J
LfmCwD/sRSp3gb+rfT9rh/T8EI951Z7f7zAM7Thq0lB7APIDxFnm6jO4OUXtTqcvXUuV9SWnXcC3
rEF5sypKG8ia+jzs/W8m+rK+cbBkWtepGIk8I7CdI95i7YUS+xCB1yn7/P8mx7hRln2HSOv3kdBZ
E5bFml3giOg4gP2UIVRXPP5i8JvYSMLmqhw6lhTxdqp/wlks6Xlp5GSaYOs3HKQGR1ScgsxRPLzX
1BRNmMrFy206kVdKGhN+ay3d1qbOh1aonmzeB5eUYhPF+s0sKOCKLNuqXKrhKPlk8/MoQ9fJbrMW
1x80aXJZuNqnWmGt/1f9pcM+NCN2XvfEdDtInMmCi30REZb5YbPkDyelf9MNWmfCV/o4QtLq76aI
m3zwC5IRDij18TLCKo05PAW6IDatmqrP/NUsBIRf40kpTxr2gC2bpCM1ezNDVyuGh6FzZv6L2jeu
QrtOxwHVJbToyj18BvrTBHycBEcwgQD5TZXn4741uvYQjn2Rpm/Mt7Yp3cyNBIqPBzwN6+zy5LtU
LZuZgqyjocTP/x6jZFJCqv1fbo+vFq1z6HHUaQTLoQ+jXNCi+US5h6Fv+ktmF7g90e1dCVgEYAby
NrPpquuJwOKkV+PstVWLTmCAzsODkIUEc2HKNCFqQ9KXHhvjxFPMWu2rm0NnUseR+cNqrxJx3LFh
eH7Q4PjILD2STmVu1HqZBWCBgzhwkhXWA7iSkzyZaFi2NI1yoCkahfWdxWd/E6xj9sMUYi/jcKLL
HncLtntkL61bqUpdD5hxWldyS/D4Tfz5P906vT/897h2Keiu7/crtfRe/sgHg+ZafMjAptbIzVf2
ARQMjj2UaGTqYauW4xV7wi7O/Jn76bgkQajSyJn30BsJisN65Cg7z/IrkT4m4pQEcnyZ0kqI+cTn
9hZKsV/2yElOqXoAK2gu03sbsWgpcVOxy8klSku1shqvwK0MouN7S7dvDPN96doYsxmXoZnrmFEz
zb0uMzdNyqzLez7N3Nad7uBxe1BzybLvxvKdTKuWYV1jg1yMXpz8z5ibLRHmEqbSyBCCDu1VCHud
t4HANHZN6q6i+BbInArOA5IdmxaqsYidaHYtY9JEs1rFU2coaKhdWqpmjMWz5irK0CAL9hbKcwZa
OL5L9OFg2VKcmu/2WF2xVlM8/pfLEDW6mnRJYVHdK6spxaqtsB/KSMONawFUPzHT5OUQfxmSiPoX
+Phj+c3HxEmFngmr5FHCH2ihkvUsle/OVyxGEVF22mX9IrzlW1oNCgFRMUH8stM7LvG+zaAy24zM
14ZWTMBix5t0ihaJHq0Y9WvEXMy4kN5SpWAEQ/cCXsGJV2KkjRzEuTjfCZuIUR1dqiOQFBjpzDwp
1sZu8GpKnXP6jtz8EBuDc4PdipY0X0QupslpNsnw+ZsxqyYlJqOB0KYbe/Udh9TDAQ+Vde2WhbsV
oec1DfuD2zXe40yRpK4Y13k+CZv4AUiwCVBuTAOY7Rdz/VUmszVAPlB4wZNbvCN9kUmFdrAHisqQ
CRVD0Dn4BRT5rSUk4YsGFvog6kdBT9/0a1nt4GZgXd3ZqIfu1GA94PaMtoIo51hMNCcTg2XvOV+j
CP5buBmqW3RX6ZCTSwA+bPAZDXlyl66zx342LKfh/PiDmQkuJr+GXq3z6+JMipsfNd2bWRxOJh2V
my1kh/O0dM7a3attezgDyRbH9J0iGlCJS5IAYGPxWx6mNHnWRvIL1YVM0zpfrZgJB0CMSVhlvMJG
CYcjg0Y1zxTH66FDxE2luuTX1u9THRGbcKLPwYeNqt9ICurizZPe2EkxKuyNpKgGUM4b//iTxD+w
VSL7WhSjLGUQhrgfHnUm4JMCGQHeLFKNr6W+Bpha4UimawAy+RbAPgnjV7NMd+ZFJYRMteJJebG8
XrZtwXw8fTqfcFf3x7o6BBJMNPXPHCRrNn2K1cTP+dASlbmTUQcr90FTDv7y1mv8l2Owd/dKQYdm
xuTNOmaULpVDNWzKIXOfdzVmeCdWNumxIQS+fktP0j4yk73Yw+Hh4ddZSBZeYF3BQTbuk2gkvx9N
o6lAXvEzEbNKhYOqTinaxRgispE3645NJ+JwORP20WeAeHALdtusQzzNIQ63t32329rdyHI3W058
HUnA1LzoqQd5tuauMGabuoquWww6XfFGJWWXMsIe42ae6uN3+v41GrFfjh5kAG+m2kFYeTw/G7V7
fxIzwLTLet6liYzJLmArZcjpZHGHwkTybDXfBrKi3wJn6f6G4ZNpZkK4OV1TDZwowRcQUq+s9u43
Xmq6aU1/pOqfkCiOwlugnWld4c4cmxzhlgWzl29bMWy+yW90gWqDsWnEnBc9V8uPeK1gK/hcLdAS
Tcfgr5n1yBYuiV3VUyukfzKf8uH5uUf8scGlcviauN8ylQ5hcM3nRU4Z97e+Tf/4r5BVeyxJeqCC
UedeKCRrrC1n5z4khuqXiHj4LsMeDiog8xaCeNBQ/xbE4VP1RoveYkaG+V9M9U1O73kFRkuhE5Yh
xQ5xxcur9d2Voz49O+IRsj9D9zeWEuXAsjLmxwAOAURi3dzEVq50ckDgC54QF9EDa1pDuhLMbuXv
w2WWYDBHy6f3Cx9oFrZOhP/KIUSuvYIt3CUo1AuXO239JtIgg0xTwE8OQ2phZKu5KB6WLZ/rlqx5
yPPHMiKVDbk7WUsLWDAjh0MfyMkurYOu7cii7/OwcJyfUcdOsQ4s5TxpOW+4G9IaYlKDME4O4vEJ
ceOu1iZA8U/pcm+wcSFmweSb19PDhZ13uCAPAzCQrOaC9zmXG+vfAHIXG3OD856OfutI5OeOwqTl
9xNkcSeo3X+Up/x/eesH51kOu6hVbduI9Voi1nRTTDhmgCOIktDbNd4mWf9mqWhvJJnCT0aQwyEC
Y76qqRfQQTrYQ9LqwvyBAhDwsP5asC66q4bT5FBs+aoEtG+XdRdibYEXeBKgEcCKLcP+YV/B7syA
WI/BXv4EyZV5jHBR4QN8zBrKt+l+EkXr1A3SAK3ysyEw5dXxIZbYjUaXLoMrSnR3FVOhbiA/4kmj
PCZWGnoaDRc/wDO0YRYRwqvYgypg+iyGpwUP37J6Jsv8NWGjNMa1+62pUih2PPU8kYOK+uhzh3Sj
1ZPj8bLqRPqpW11grqcRzlp1NOOwhIrvy8EemUs1jtsHZa9WeghEuB8W5R9GggfztAlP1JHJ1K6F
iSeCg987WSkRcx6yaD+BIjnUgdKkOKHY8yYq9z0cV/9hb4xuRhu8o5wWbDAArgKa0KaZeB9DqpfW
bCjbrktACCOYr+9DczF0yWmYeF+XdkQAV0rPYMCfgdY5RecW8opOsnBGGe2VsG/HBveUM23NzFsH
xCY3djWl7dIafXtfnXmGib4PJZ5V8GMezTS8z2Cc+5LptXZJSKdBJBSU3HzpRGtwi+XSF4Z+KCRU
Dne3bjINfFGk/eCsOwYm8Lo8w+KxBSljpA0yHdxomXIotJgRH4hsk8CeCHo0pjnyBf1kEiJbMgOl
bBAmrN7npPOdSCD6oT0OhVPWE6nSFOyQhKHGnubrXuihiZ3qxJsuYdnziXTR9tMoyuInortlm11a
q9Bah6keNHffmc3tsfJK4JXq1uH2wKZptthNgAqiDH3HjFOzqo2y1g6dYdEppcuigYjQGbd6puFh
Ve3/LAcLAKaNNfG37gc+RtAy91IVpaIT7Iylue6S8N9It8p3wc5hXSTossmXk3wx9Ztf0UTTpUSM
2/96Wr1H+WmAqBG4Jn8GDOZBGsQ3B97mPyW4ObME7tLI3lt3og53Zf3VLurXp46i5o2UiE1a2Kv+
NVWC2LOXEx5xZNJZt+YpN5icCo4w9ThV9fVwtwktfSWEcnLEALRGSAO1ByTSjF+OSS+WLqwiwJdq
1t8dz6he/G8WOFjQzdfz5IQM2zBkZ/lVGgu+pxEYZMf9SZGrJVrui+pNWAyYX/2Mc0ubnBvFJarc
S3zAqhEsP9p/sUXBiCp002L6B+6gGLqpXQb1IXtfGY3/Rx60Jk9OJhg5aVlI7zq8ALZvdDno2jok
3R3bQeKeLnXGkpGsEosGfFvVvB7+G/cQYjUa2kWAPKhCj6fsOdF/TRlQJ2mEXuXJZGLSBxxfRNGi
2DfsR5tH2bLzxNKbDrzos0Qu2ojI9E1JuWuUiSfFF8yHFYhO+hUVA2HM59QHR3il7WxOkGm3s/Fi
KGIZMn42sCOnH9NMM85O/sEns8TvoEQmnNJPzQm9o34RTEqNlMuytrphyRIntHjCDh3kMuoggu0S
5gd6CtnSaCLE7p3UlgzKhyWHKi+sJ6ybiPcdqLRkB8poFl1FGTA1im/eFwFPkcTs+2LVNykJUD8a
xW95xTZ8gzef3qBBCSMU3gkDsBaMI95C8X/ez6xAl3IpNZhbbnF3VN12VJEaZsGCSXsJ3zTCr1j4
uAf3Oqkm1LU+ilRfWW+y7rxaawVPAK720lhFoFybs5iqCzEtY6zil46PnyhDSZ4HkOMfiMOYvdAr
C6CnE/63Bk5GVK51QLsKHThQEOwbP8V9Y3oPWB0KZFl68LWzbDKXBvBiJmCIU2p4Ql2a3Mx1MOxV
Tp3Bzz7taD5zSJKii5NthdAfDte/qXtWC0AlrB6Jz2v8SobFhh8nHkUyysKxzDJ5zZJZx8GAtuhq
JkXzDpCX2GRMqWf2znmJHmi0wWPLJbNEqfFdpJ90y1jZOYrX4fs8ZAR6TKnZPKKZQM9i8V0G5Ook
vXcRMZ77uqVTr9nSz4TjxTpDUPC040dpiS9lr4/Pge4blbp0W9dE+2vpDE0ppS/9XYCfJLOzir0O
aThf+ogTlB5jJc+nGBMPK4JZRSVSZhQpJFyZZwm7pdHQgZgUxVtpvLZsAfK+AHU26zwk0nJGkoEe
0uhdvkiIei2di4HfjIQtGUHXXapJcJkva2PqEYSJWQXbi7tg5th6TfaYktj+/1BQeC27RI86nafs
H4eeZ5ugeejXjPfviT4FxN8q15tykeCq3lN2lnpa9MAYxszB8+tNY2iCrU8BQFcECUgeMpyq+Ukp
cBN+mMpX0GDi+0ltAogguiPJ7ViR3AUTkcSe3jLoijM7ntf5NdBBAM+/jFyFmXESQdaSD9Lcr3Hf
68WiQAL9stQv+73uiCXmdf6/jGh2OzGyD28fk1XqnQmAlm0NgtItm3NhmGPNEw35X/Ms85WVGXSG
cZ1AcwEOUkJNc8R9o0Qkj27v+zy/aWcn2pNHT/wQjEeLyVf2SL2dzzY6O35/mTtdpw5fdiUh1164
fy78EBB3cdrSAvmHizhF5LBtrUnukI1ZK8mBlNuwu/zmjmJnw/6fS5g/ih7easMWcAv+SkzCmIpV
vB4Yuoa8xK0ViAoT488ZNPfl3EVNcDjiUB6tWknYgY0CWEAWHq9ZUy3UrwUEOlz8iDsH6FGjBLAc
ejNrqEB2EIKHUTLM8CMNysy8xQHtED9/N2Rco4CdXGh05hE1bnWDWgGSrBIR1s0pkWAf24TZIEZE
ybx0WhOFXsOIUutbnANOipsGsb1DHXB5P1kgmcQJCPs1c+G+kW28T3ez15TCE7aYzj1cXD16Qrf8
z00cGBrgrQPLOjZnFX0T8QTWvTOmUVO6HO7qW/Nkyh4nRxwD8U6rNFMAPs6nyxKvO89xvHiknMhh
w4AVkv6TnFzirSMJzffvAcp6pD3HB7ItRmO1ScBg/hylxJKi5rCOb+3OfemtJYQx8yOFyiOprlsd
ZeIoUjumYPCdX1Qw4rSATqOy/J/fBWv8RCOJ37w9Py+Ej27ewYb6dVJR0fq5quJJrbdJvXm2BpiM
XY/uskNonOkvaN5V4gR4Ry+h+yNWgBPZF+rQIHWwmfGrwqFOP1mhUVEJnk47buR1RBQCLA7lzVUJ
aJhf0yXsHdPMy3NtZcf2T4AudWUklHvG2gJm9peA6al51XKevMt/FXYsFCv2VbjppCMMd6LDdp2W
INUecY7XTsGwKP1UgRKLx1Gi28F+Zv84jtCImBAqT8Z2IhFZY/EByzzamERn4nE0WMXxxUIuLrcI
R8zEzx75/kiC3IKld0hG8oGu69fvQZ3gTdtlwEzNDQPTq9+HWO/XhPinmhLuUIjoOub879m48pwL
drlQTRR8+jPtZJ6YHkyDLuLXYsTbcvRCQSXnWJHEzrqo1PFezMOtX46npFgb4FsJaZOWjTfYAE5B
3oJ1o9cVbokpC2r3JJhy5G1HZOkUH3VEF2z14s+KN8vQGTOjuOvvaPbJgkpGySO4hYjhNaOPDIsy
Yv79UzURLYPY4NltloTA+G9DacQv3uhQllcAXc/qsXQ+tWadwwNSl8DLlthorNkFR4Yl6j1CCW5t
FJoobL0ZsthXYn5lLqGaPHWmeO9o+3+WfBXJKoRoOiBaiRRBygh07Q568D5NiJGjvj6ckbZ3TbXD
8UIedj++mjSsn17a3LuflqCZgy0h9lfyazhing6SAbznJV4EcjQcx9aFPHE/pLr2qiobdeUwWXBe
2OX4b73efAxntButDxn/WgzaKqmzKhcSxkQ5Rk3DB/uzsnJGS2zXRWb1/Jl7fsnsoy0QBU4hFu/D
Lau60ybPfNlNhKtrNuuIRgV70QixZcRTeKWka8s+N5KjdPC9wSthfNdJ1hRH7Zcimx0AG+sgroXC
qwtKUcFhkFNhvMJiXNDjdKUZWHUFCPg6yS0H2uB7kQHiDp4EeJ5YL80jtlIQrYin2z8W2bjk1Yzo
eF8xoL5EbB64/d2PtuWol6ubdnk33zK6RhYzkxxC8pZZ+Se/hUCJ1a4EHee+VxYxQIoCYN20ZvLu
HGpnS+KaThWPd2LOoTmgGE3T00HAN2hK2saQBQ234qwze5/Rkvuiz5GdOvgp6ulANaUQhFZQ8dtq
40Vpe4t9yAoBqNCVZjMMQoXMXPd522nKMwhNq49I1Vw9DCY+U4q64pSopdfck441Kan7DY4NCudX
hEhqLU7jN1+0rVIHZ/MEutHsXHLwC+q/T7tQItSaeGkbHNZCPfog90dTqydfykKcJlHdWafnzNQ9
Hd6unV8XParTJzxsipfNezqf8k5cX/SGn0NeRIex0fhK0a4FAa4TieL8m3E4bkdBQVdZT+wNY5Y5
gv/4JWnC+O0I7bx/U5YHdo+CjqdVnvgGFkJ6Ajo42eA3bKkWhmlCescybw4T3FrRBn0hVgMX7hCc
aao3vC2AOq6ISSujEPkUeZ6/Cidci5itDuBhv9tvy9nMlYjPxLakcYv3yY53sYzc+JZm8tq/Ll7R
DgOHX9T+nZtT65s9SVnYsb8my10mdYhEUu6D49vhC2+PVR/+2tZG4/83kgFlditDu0CPFJPFbXzo
C3LIvtin9+qrC+PFRw7xJpMSSCJH25zkX1TzbvjBmndg9rx75tdp8IiKpQdbgtIxRNzhM8gg+JLp
XXnvFet3rGgezAAcR7w5nIfW/Gww8WVcYfaaOLV8C6TnGA+6AGFe/5GZbY6NSy+biznSkLQ08Lfh
OJLRZp6gr6ICFEXm5rrn/kTiWHgdEFWov8STrH2RSUEoWprG0MpQ03XJlBmbJSu4XyXuSrguTOLI
DO4jId9hiHsU2e+VC8jdypphO6dYGYpQLPfdKfPsbVeB/oX5ZAeDdlFfuKb9gggPgpaKaLu3oMXe
FXMusZ9PKlZgXkg0g86gQgm5khzv4BOj2aF51LIBbA7Rc/EC55xEezSCgudArC0puIX/qip3G4Rr
g7HY2DCkvomY2UTaT4F/bWY7M4VqWw+1/paC+Vp9uZkjuoAi8mR1Hei0fqimxcKrNO6du31laUpB
mRwGZ01Nrs2RBccNrhPXes4ar/L1tAX6va25Ah932G98M0XdPCOn0EtrzrU2qUV/+UO0YJHki5V2
mDzpSFAd2Ldf9NU/leW+gX0t7aB8X7YukRm1RG5XJGFCaaAAzHS1N+UgSVA/8zhzK/Gm9ZXvhT30
hyxI70h/nQKnfEuUuwL96EQ4nKuh/81RD541sH/O+N7sOJ6Y2hjqOlWtbHAax+J9KQVqq3bOBemr
cHjNSpL4Ni1F+lJBWQX/iAsQjbrTIXgdcROY8RIiWNAuxPKDh/ZIjcL9MfFlCRvwmnXr0c9iugra
B7AGxLWA1QJS801W4kq5SbwWMMofE7X0fPp5f+gC3DzPaepj1HZX2UdrfwyJT0JVHH3hDSkJmPqH
7AQ0Jpts5UrVJk/wAr4H7oSupmkuPMWQmjmas4MSqgld8gxpTj9TMYBpFXapctk4VUhykX6VNwdV
BC9k2yg11nOdEY84h8XYNeGcuxSZL/bMoygooG4zR0e7bfjFCuTr0T+aMTrELIiA0iUZqH09mlNG
XC5CyY1Vf2kPtAapWlLqDIY+ZXl0ndt4QJMYLu57TXgbHoqBAWP+UQDCAkeksct3GEGS66tG8EBR
4W/I6mq4s9XtpakAsKPkAJM3XrLYEKWyqXxxUV/+ZXxgpw2Q0eTgEI5Pj2FcWVuzgYaiQ+WNn+fP
hjGqn2hUJCfJT+D/huR5lZ0D5zKlja5RuxtDfce2TnARt9Q2qhO92WDzu0twC4QpIouO/egm4oh5
tLoTYjynnTcsKyDlRKv0mm7sAUpsh2RB7V/3OyabDszARslNJQZ6pJzTQu+CG/C37n6yDbkCxTtJ
1HW+Gwr0Pc7LEm2pcGUvMCNXiPkLgwAK+T5/qkPo81hKgmdbSGLnYXpEwxVuQIwfefgW3NDzgiXj
2Zksw2b/ISGlwsuET4QoN+v9R3s3uv7aM0WiyokD+sg6TlNclQu+vBkzCjVPJ2/lJVeg5bcf9sHl
kzuQsFswXYlrRbN2M7o1jyFJE2eJe1LPdCnaLM8YnCRu33k0Z8mdX3G5omIaP3L1rkKwrqmagIXT
E+/iRXJZosrrwDX/2o9urXogg6Yv+VTDZDPywLFmvb5kzmqMJ5FpZTGRH9UaSvVRrrzGn7+covfM
FVTppDXhbQe3Jh1W//4y6JBAQGw8aIfxD0JtO202rsgznhr6qAQ4APXnNrLroGDOr95kcTKtcWyc
a+OlvEr48domHid9gwJE0qp9J42GhIm9fSswtLwXyfXk6oTt7VVOxH45W6ObSLwVdGxq3jyoD/8y
nStdqzqQ7kxGO1drRWmWazJ9BpgE0Qf1xUUJMhSxDXezz9BVv4OfxfJ1KXc+t9oox9cONjmKieCt
pmOAJF284iUaDSMO4/7HbbszeViCk8xttcQcRr3t6Sl8X9tWcUJEBlbth1ieanJ8sYUN4J/0cE/h
F+8yY50MGr1aR/gPoMvwwBSD4JzwMNlQHw/qsZPUH14ddhLn5CA0TlOSxjSLtC/iQ3ij+hb8eB47
m35XElla+Hah2Z/JjtxaJWEIM3kONXioxloEbVBbTnOFWFrD9yWkPUwI1K+3VMNwPLra9qFXKPRy
i8Q3g12qibsU5Z2g+ktQwvrnChRlolVLiKDxg14NZeB+BmhR+bk9QLGIFUWfzKhwWPCcSQHTg6gp
HXGTjqO+VxrdugU2GU8yJFRcKupkGXm1STjhEfF2GB6teQ0aokSdj7dlstS4GzfDWpNVKnO0VWHw
eYQ5t5vtbbt8YUuqVdZhmgvPTuYfD/4FfHh6X/0Py3+T92uCrTN4nW8+dHHtcEx0RSzwkgGH5lrZ
jWeHcVt33vraIPF74tsVSs3pN9GDXT/NTkmQD7LgrlrrpIVtQszL6+TJn81YVc34ehI5lAj9UaYM
jQh4JhIiMfSIGmiJ3Sh/z36eWtIljNPEzVCnd/xiVsS21871dn/TDlrhmeBfFjEBmi4V86xn4B9u
e79H7oWQlbqdFMqo1t3XBFHlaqKq6wIMWTDWTGFz1tpE6gvhjbJPJPrNP3MTEA4bNvFskal1nQJi
9s7Ela9nEOj3plEL5+Nyr1JHscJLatB18+FPZsUG9o9bleWAe41j2lszPJMxVTTtJKVgmtYdWWWt
qlL7vYrJblk4uLFvMB3SnUb9tejww5kxTk//9R66ewqigEQ9pEcNkaH4NZ+3uQO5Wv3Q63g5inIf
DRvrxH5F5FtOATpYxzeeZsnidb/xptoc+ljXVBxGorK1kHopwMjUeJC9Qnu9f3SbJ37I0pp+0TYy
HIOFpHfgVQlTyyQk+ocfz4erlpKssPJLNvd8ajzPHziIBoojpy4Q33tl2cfQ9+4GqpTlyo4cQFlg
APVoVasnf7qIyr+GA+xywOw2SOdf3RepxNp6lVqBvNSuvQcHdyT17vPXlWc5gNeTgf7WXhM27+G6
h2bi+m5x/OPS6s7I+NjmdQ/vNlRVMjwboz+NK7EiZJ2M6W809PJS5XMbXi83Leuo2lRm4Ar4dJTb
uRNHBG/hpaauQc8SXJJ0/A+FJKQ6K/TZIBJcj22mssTRhKmnJEr+CPz9kEVd0iOo2tdUP8Hq3Aup
F1mCNe2glc1EOmFBLE+epDtopbWD+iirq91mwuGgGME0AE3+Ux5Mcm4CSN1o+5iX74ZuJE/aZBa1
gGKXZlzdNIi2C1PeArPMjLKCAiql+XMX83DaUcGZAkHcdLDL2IUakIuvfPAMxaEjDjDIaWY8uYiz
k2auEj5WYixnkaSuEKR1zPiUaraR+Sa9zPLlR/Rzee54FE2XnmUUPSCNUAtPT0DArf6UyD6o+w9o
pXkNuM+ypOVZh/En/u6AshpUBmv5cNxHVSGpovySFIDzysgO3ECQdXB4OC/qP2h6ZUm0UZ1/UDbe
0R2kcoRR6gogmA5atDJFaUfy6FYqlA7LSH4dhyCg4d1pgfgLStuS8JdrGNSp0H1i72T6mH7zYS2P
ogEEcuhiLyJbLAPsw1kV6+byTN6dYt3JjVgTbIwpQUp7X1DaF4Y3aesEuZG91VOL5O/STEwUZapP
pvKNCDb9GdBLCbX1lJKolxkHV/aCIwdJZ/HIgE+1Kvo1yX2cFUYJvDUjzPU5Y2VXtV8OqCKxw1+w
lFjrbz38yVNupHmnKjNF6Bj9RySP/eQ/ULU3dyEl1Yjwz7hcqVOzgm6wFsq+ofxdWIQlBoOsz11e
eEw5iUfUXykCSxcDW7iDGWtgl3xdP8XFEWyeFyY30sH1eWckc6zWW+SCvRWdePf3SkcXD/G5hRBf
BiKjZ0w88ZiI5WSiigi1CEVH9Ptkq6tAgODQBMSEI+NYgd8idyhONe776ipKlkBfZ38FW0LEwl6i
GkIYaj8jcKW1hx75jGDomnxFlROxDV75uQ9Y5HiMHAqaTtIY3O1bRNKol10BH7EixIbVBgGbCMO2
PskSNhj/Tsk457GQUYvzZLwBycv3zHr6vwmI+qaQ5A/BHwnxUUzDPmEw37nPqJK/DLYYAjvT7xIZ
BTO4kok14+G0Yk3BzbNdRtCFf4Xh0MJTWCvLYMJvN7JiRBumaT+9lIhu84qO9UxE4kgnTl2SF23a
MkbNP6WYgcdixnEDyprOCbjtlc3TERg+MhPxm9fXwLHyhYnSkjz0LTDW3gRkYOqcjG7iVQPqIsIl
/7hQPdhX37iXux4j2pIxQ7gpubv/x/6nS1Hm/px8zFGQkw7/D5kix5RZ4zXyZ/7clMmtMzRL5tq9
9z3imJLufURFeUxhorPjmLCOFCJDBYmK0FmkKMaRdR6sgUyJqRgUYrg0ThlxkfE/MY7JeqrcjYHM
SIbAZcse9iZvLHUFz9MclJ5U4SB06dvskHLUqPJCIx6h6rQI74kaviPz2re2rSvNbg8JsvmjtKJH
Y5BMsfUDNt3dUJ9RH7MH1NOfNOBC8CRs13oVWKv/kgTxY+z7JVE8i89tx8S/KNucUmJPDrHLQBbK
91uh2vVm1IGvxHgz1B/jXrgoLMd4rfmP1TUTTWkS6sD1jDvWjZrwxOJLv6gWTxwtFlHTF+YiK/Xd
extb1EBNtloGGq4kmqOscpxT2O4O50iZlPRu0YT5VletUBC8ZC9/yBnOLVa7iY40RDYdniWjE2UG
JS5iaeIwbG0bSOpFWvIDCn4zS/ifz2g3GLNBTr8InXb+S4e2msUCdp5MBQrDSy0mDXq0+0FCUPDa
d4qqciN/lmj6nl7h9OeoOnSdZviaZv81THX4xwVCpvcJ21Wj5Vq3IASajso8zHuGqD07Z+cLOOZQ
3tHT27fq2VMqcPSp7UEKYKheWNTUI7UWskvkWHE3DQp3hbdjA14t23eumQGQFO3taeUrGLzWmIsA
0zPPMieU8iV0WxewXHWTkfuUy0yY9RAZO+GbAtGelTXz5CCvJcuWH3VpY3wfnX0RYc0ihrE7NSra
3chjAG8UR4wK2K1IXNk+q88szrKSLLj1XcPwt7u/U7zKN38pmEKzs/228aFjN/s5HbFOrfD713x5
0/oLaeNM27IIcmESsdKEMIa54LApknaDA0+Cnsoa/pR/ewkt7ZJFL4vaMhjLNtNXK37ZtqV7qugl
ouuOdS9eadjR/vkTbPs18jpdrlH4TlL6AGafdp26XbFzzqPefvPgxV084pj+Ilieiw/fstPErme/
LsLDNXZCOENLMC4pnTWeMpW7VZ+u9ZggrNUbiJdGvBHT4Og7xdqzng1ALaiv87dyhGhbbLJfChWI
UZNzUzZ0ImCHdrMU51z4OeDZzK1kbZ2v9Y9KaUj1q68KSYOBBeiS5rqbOrlduDuoWzuSNclTOanG
rgsMWYAyKDOM8dhbThhXaBUMUn9gZ8kYBdD0MxzJw3YfUPMXB+28JuMxl3bJJC684y/WM/SmZjPB
ZgT1vkiGYqgDM5SJLHlqJ/QxpV1+6IDlCsFAEo8lC04WYJEjFYdWa/LnJX771mnD3XVfIrLDYOoe
jNwcJ0Qts3UOiwYFsKQpZw76R+/JX55/1//G4mKHKChO6NCTHkJn19tgrhz5Ors6r4lnD+BMi2LX
ZvFIKwd9cyKTwlMAcsUS10TKoZBwdjIB4YUtnqoj+VnYPFlAOZC9IhtRxtkfTqfAwhQHtxm9ssKa
G84TdduS7pmnv6SdqaJcZi9cm8G4GLbd5ZbsfZgCe/dfyZ/wDuy8ULesgcqAHqJeoPCZRt3S7Vcl
TIOOf9GY1PoC2DK6wuSoLUDkxdLqajyUEP9IsoqEK6sKSq3320F9YRa//0QVHhwKiyTubYe9TsPa
sHTjxIhlDdnihmofi2F7uhZoZpQkNM+inifp2tK8kaszMfe9E7Hh3Fv/vyW5qvlrxURX3PTZVa1z
cX48neMv4IvEdpng877hhNwRp6/FKeIgThvGn54fffMTkFhBmg9BMKrXnrPFFRXJvdAhhxdmM6Ao
UrwUN8hgmCZmmBjmvzgO4zUogGts6vLMKiMIqmz9uS/BCliUqPSN4TSxxyxhTWqBBx2IgAS2okcF
wmp6v5nM9i2+7NINt3buqqmvpEJgePTb6ajxVQynWPgh1UXKsbCxVVj6lSUIjWW9qXSfTBWDomD2
qGRCnH0qxpLdCxIJKpVHaJ0KwnZosw/jAS6A1jNaPHBBo6wcJ5h3G8i2ckJuH98jGr3RokZEeFOi
A4jE4ev8r3izAZJRY4eHKaLX1MLpujA2zU0KzsSXJ4RyeLJtigUB9OtSYFPDECRX8CAzZ6AzffLJ
SYXg7QN+ZHTwzHfszR/Np2DwCnxnSGIxtz/Acb0KhW/bx8C+FwmKYBi0jaFszRVnJ+f4y/sU8/0V
oUiE751KK/7mgTzgBFGLozvSTOsimOZBmx2Px+8AfbBVVsWHCWOh4rfm3WI230WCgCXXcKZmafLq
IL5z5TtkEtAepaY/GRNErtlA9kxav8RjPkGEmVXIC5oGXQFWSRchBIdtGACGZyPKrhRbyFnD6VKL
ypTw6X01jv0Tcirm23STRIBaQENDpNOyv5AaHo9KDzeTQ+ATqMNCDAh2hZLRXfhzKpDnTg4cXidw
ChrxKXEO3s1g3BYabEmIPk/c2mCsr1tXy56/DOj+CzpxCPAIV8YnaBJ8ursuuvhOjd5j3LJD5cA0
oYGmfwHv4GIEXTMitBNMSb2xPJuXG+ViOaNpfsBQIDAXxrXDqmYhYVKQs8pF2tjp055marr7Y1/g
5PDQdXi96uidIf1/56lbnwbuboFrLhZ4ICYx7LZkWdOKsEXQz+aPVp/LI9SAbfi4x6sa+kE2Clat
OqCwPVO3BoNZgLuTN/Rn3MJdvRFVQA3D4U7qZfuod6H42G55hr/APze48i8RWYzN/ybiPhDz3Zfa
TTkhCLXhIwujEq8EZe3h6ZZ935aO3bfM7QB0KEG90pKlzXM2IPi7HPh3tE51cfc8e/qF+ntCtVrG
RoV7DdJnZiw1fiw8FsU5p9ajTaUmNp25ObuRNRJbUxvdMK7o5LIW4JC0tphHiLC0+6satlyeq6NO
ZQLAFiM0NvbknpDtF1J334o05et8IfWnROXWF5QoK2+WXFmR2AXZukwfvHcxWhG3JMlwGdDvpf5q
j4WZ23kNvtlfSNPrid5ipuK8NNGxJra0QyW89cgI5Iw7uI4VLXMIuPxP2wvSX2X6PMQBxwtOj755
gpEutLZbkDl/ZQKRtAf088xLmqZTAzuH2nNJqXIBKc6me0TQthVSYLpQn7FZmSlrsBu0c8rcetNp
LYW4eOWKdhK0ER3OWYekue4CCTOlgcaktRehbt6iTwVfDdnylQTxiH7jfH1XX7TThVaoDErPuIYa
4ytoJey+lF8d0DGQZCUhMaoAsX8rGEdqgh1V99+Dv1TVT8OlNnxX9YLEK4drX4xrbwhe+PPYvckx
fecMe/m7LG9iEXJDUu5m3QoOh3mCvZYqQ/Ivj3Y5AuUZ2i9/T/VOP5u1xrO7eGljApQhfvtxIhem
PaRY489aWTQQmeynXxX9fOjQVQ79tlSO1hXi9hkQc1+Q7s1oqdnAPh1xVxXlLWuotJW8uXm6n7z7
2G0JG4/xCTODqVuCE1QQXrq6kMzHCszDk2nWRPPzsgIsFbrwHk5LEFiFouIh4tnYAsi/LdIFl1dU
PXTiDDlINmDyS3RW3OObNQZIQGmub2ki7JxW9+7g/4ARpKeApk3ELOP7xBg2P7IMnUeDjS774A/L
e2GGCaBcXanfVbBhKVaVdsDVejUEqivsbRhDKPQBZxsld8v8zM21PoFBAs8opDxPXTeCUN1V4K0v
jP8gOSaBMi23S+T3Scm2ac1aCeMkjncidCYQ3CSE4e3McAOde28zd9mC4d52/4fVSQr5HerNo0ZE
pe+NbMDrcXMHAjeF6UoZWIKuubUH97MtLfUaWaPv44fbDBJObSR4GDKzqbQhRcErUwntdnXJpRUz
Pm/r6fEBk5fV2qe12fqXK/OAIZu/bxp40WO7Yvo2QW1HPATGe9Awo0n4iv3gdXHW/FC02ZTNgyZh
tqEd8/mYCFOj2zHN8/A9ZzhFo3lz5D3adBqlQBRAhiVhayqjDcsUiGFO+OIZ+4cEuPxHhjQhxN5q
5h+uXLj44SjTR068dLeYCOCG960u9jTfpgu4s5e0aCn1nqgWW+ReLlZVxD+EIJCy4yf8CVNUa0gC
nkutiUQnYFxkmoznR1/Qjx7IuONGCfP7+CqtE+PlMsu6o6xZrOVBbxt4ozIqifr2hzRgorZK52oP
+4muwopuowv4tYWJ634UQuGZkJrNrOuX3p59I9/NmyEAERnWf4YV8kL/Fmbn8vhM+hIp4VgfQsBu
GatugOO9I0GcF1jxaSEJzLOueHbZREJ4WmDrRHdiXVLnyC+gRSAaht09QYyRDY3Z7CxaddZR9aCC
b+nWodWufUv4SahtUotipjLxraIsgsP0zCyJ2FHthpJKPiNTmevc6dI/BmQAi9DgQ3+Qx/dpfhUf
xxu6MSVjo6f+9hVPtBMCfNRV05v38pl+IAOOFT7f2jMDhtGtjYc+AzH1E9GW0/GY7pDbcvils5oU
Q6nXOsl85dxXIhsIerrnlpJ1NJuBFht6Kq1ZVlilpWNlr6Ikio70TEib0LG+5D62I1bOncB73xr0
0Af4wU000Y5pTshzAB1YtSD9i4Gfa8dwh4pJ3vA7r2ZSuwr+MNM4qKSafUEcB9+rNAtn8W2FirYE
giQMA/q674gE59AHOqLJos8T+z+vKZeIQqrqwu1ISNC1oonWRwdo6xMm+6dBawPv0cc/zyHwIRHo
m1UYajZ1t3exnOD8Mq53GwNz6WOvrXVfn15J5UgMsVP9SDRO592a1+btz+ynM7yuXAnxjABaOYKm
73YN9grMI1NGo9l2qj/Xc9WQtTYiNKAaWWEs17pUN27IFRr1H1AiMcMA14+2oywa2VanQDI/gHYR
fYhrToS9XMfo/w3VL+yuULbxr8jE7q8HHl54YwYKG61txx0AlgeKuDmw6JukIOQs6xEXGLJckagB
BY5toe7PKb+ufod5M4+IfOQ8c9Kv79yAJMZIZjsFPN+SG48HekOIeoapPtH0+0rqoZ336IIYj6/J
uwTyK97iQ+wGsV22cMdgmyfkT0YJ/lzJT4Gt5DoTpgvMuG9S9n0y9z6DE3wDCAW8WexBgXYPPQZB
BHKp9vZZ5uBNBp8hY3xH2S+0jzdzV8xil3FNj5fT+4HwGhcUKQaOzuZNNXq58W0raLij0zjYxQI8
cbiXlJAfIGs/RyLYAD3Em1nl99CghqQ+JgsehbXP98X9e7tVcV34+2PYa+eDQLOE+dYQRmw7Z/oT
G0vJoTOLO3GtD4vviwWXD832TnhOlGVNgu4t63rkWsQlU9K9FGkYusKU/w6xbsb9O7Quetj/ysQV
f2Ts+la2T6mSi+4D4S3mGEo3hvTbg/HduoKUjilNEY3wKCMCQOKo5LRk7MZ8HsolHpkxA1G0Ur0W
2tcPb+kc4mDlrB5vqV8rTmNz8kbX8AD0psXbEP/AsSTpbw9nPMGukiVSRUjlPaIGGRPk9I/fUGB0
7IW/Fe0oAF/+ebQltir10PI3xXVeqFQFuOjZ1ThmY+GExeLKG770qZFnQ8ogTSzk6npIDktzwa1v
QzimZdn6Rnh7KwEShwKqKp4vQjr43mIvvwEYwMVjpcsKpz2ItiqzxWhmw45wT0cbNy1UmiAKivek
FA2UjZ+5tZflMzMkzFz6FOrbJVcAT32AvOkP63NG+rL5FuxgTwO4XYQm9xpvkFP+4Y6teLsRyJCm
f8nR4vHlChUCpiTqob8J2s7/felDZv6WVdjBd+jzT278jaz7Sm2mvoilwez36Nfysn31eboRJEaw
NQe+j/39hxKYMOSxPWPt9MIhNSyvGf47wzBNQD+bfaSZbEicWgNKH13yACrxlZo+ejoQpFHzisEc
5E9EPTIx5HMhERwLv2x50bWhm9d3vOI8oP4XWNUXUjMgsTfE7S+mJkmJZdikVo4Am+A/eIW/Nt7q
t5p5FiCS6pIPTaIw7WFXwSdrTQBvZ1BeHlR34qQot/iIzbWQGlK7z2QtT3TVjwpyL5kbVVXd3LCp
GAwAuaHGKTzUwdBVX1vNEE5jmVOzGdxs2nvtLBYPnJLON0o8hT2/0hOFt8WG9DSaJTjX59KxzMw5
Ff8+bE5OpHzHGfb/NHX4cubVZoX1Bv8DlklbpktnnYifZjQpGyKU9BcAgwPfd5hxQDgFgvOKQfKn
im4cy5MnHGlADeGxK6UTO3NQkOkIk84opgPdATLn4ukVfcFyOipFV0F5P9UuExVCMAlwa7CEuKv+
KacG8MhsPRyAT5fRI91wcGOrRGOm9JgHVzV/XM3mY9ISsOpKhpBkRnkyEFYD32AWXlEqyTNBXlkh
idhQHjTx6IDuoZEKLdd/DKx4qAAISd9SPsRo1fUrE8QUIR+/BCuEyBMhCWNKPy6zp7uoBtf+gbev
9UE2iZZCSjtJDM9sxFjY3WL8DEjWHCzQi2pOgKho4npaMAO8jfNm4EX4JUUi3ddl1vYvg/c1RRHt
i7WlhmTf+jFtJG2u0HA5x0TNuQch+o6TXezXEGbE6CZUbhCFNe7+4+VHtK4W0UGeiAFYpDmTmq+J
I8m/ACIfpTyMR5p/bc5T2tOaSKw+eAwemuAlhxrdUcQiz5ym+cw22fbjvUr8jp4KzM6+A3dcL1nR
ZzXRDyyoXmgjXKku12KNgdU6nH2cJZWDigICVsWBYJrgf8ZguPr0W385kti72u6rZliT80m9axsT
no/K1A4ZAY22cvu1eU6bXrcP5QHuPBWIcDZv9aHAuT1qtdbnw5Qozr0NrvySK2/Nhx8fovrJXu2i
XomPLYQ31ts2oSbYvTia/wvwQShx3L6aLpqICij0l+A2UpggQTsXSQBppLf4hv/ZdmSeOxbBRYGF
KEe9hOBka37mjOVnSJPr/Xat8ZN7LPDWwPtunlWc7pTfo3PNTalfkPjfWNZP+TR42/0M9P2gmX1r
XUDP6HJd9awxiBZAdTMsm5nvwFgXAsZ+reRq6XGfnT8Tf7cn9QvRoRjdnt35mLPyvXO4qDGKfGoP
f4hVaMvbbkM9o3ITA3Rs75I3rzL6sqoR11lHSVFJGY2b+fRipre8K6tH0HQ/6/4LtZO+qK0rCQSf
31tJ+RyCrTdmn/uVEQAzL9NJjOQpDLMCrWavoKaCByJQQfe9B4fYeCzCcrZNl0R1yZbKI+7XM7Gw
FY9T9jDNHsk5KcVx8914+P0WIw6KMG2Y8EWUyKFTM64/+WRMT7cbT2u5NWQSQwXrwbndwsgO0X+8
b13xiu8wf7uLz+MM5bbwpxCGWggv6JBt6GFz953YgcTizodFJj8RjkEXho6pi8vhckYEXoeqJuUL
jSPzQdwVngKG81tmv3SEWht7njdle2ul3JwjAqZZMiJPPY8j3rO+Y8RNTN3P61BExUk78J98F9cW
S9EsKA7VVo9oZAXf5grqfaPX2YdPUAepVpuuNJ1Z+B5lpPgja3f2ErYX4/XU4ETT9jNJWAp8Zr9D
TrPoqY/ocI3b+6G/wwck7Psv2hAea/sFCtcBBXkdiY9IuRyfo0p1uS7tuGmsZQUUKpqFSkRDU0wN
f8libkI2T/ViTX6or65wKjqzNUaBz0bLnnteUyoIIbnMdfjP3joGeSR/AYhyzha4KwmX/fs8p8mc
nMQLHzlhsVLH+IND85na7O5cvIvTo7WTMTBNZmvYMCqoR6MYkl9cVmWG/2nxnjzY9tjdTg/ht4Fa
5J2G5ctTAonAAVV5xIPZVsiRHtdpH1pl3c1m6BSAp7gmGsR3tSCCHPDcfUrFM3w00bY0sn25cUGR
+F75mXqckb7fK+uKVzgB6wRhlpBCSjWnvmdLLXVB3TiTSUHJj+jKxs6ZZYE4wcNdLLFLM0AOQqLO
ld7kY2MQTDR8N+NbKNXkX9yP0WXWqjkihlq6AM3AodOahm8XbB2VnoAWK44fW3S3YF+rWS6JNDsv
wdOg35hvlZ1L6qmTacNHK7+u9lKfm1PzGEi6ypLXgDPCYTkP5AvffiAZpQGg+HAFIMUPC8CihOVj
4BtDfA4PXpFLL4AkC29eJmgrfvIa/SyJ3b9cJdUCF7SFkUd37sM9ALNaY0fGXAAp/L2IfpDKRvjk
tYS5dvrZCFeJY4qHevBk1AYKP6Uza6ae/xttDNMG5DIwQ9Z6uioMnLAlYIxwU/dPufqvjamGSC6L
3BUHi2LVMCNq+5+AYTXAalxUDx+ohGtc75RJCa/mb7ejoZx++HR1nkct20pq6En4UhQmAlB1bRnu
0Om9o+nhnH6zWGlIdCU6qGQvoneE2KbGIsaiG+bxsUIP2GsKTCAb1iDQnA/r+3hvxjd7MddUot3u
RnVkkAYtTB0tXVGbp35Lyso1cUIj41G0q6/EFs2uRwIgIhLCOzW8AQfmKewYu0KQiTz2wzmSUkTi
HY5fQll7q+ec6vwUk+kIjGdfJ5Eeh6t9IrlJQEm8nWIzBKvq7MTlKD1qgVBpVpd1bDom/ePiJGQa
rTSCW01TZA09jZpo1p6M0wMvFHpqSlD7CvD1fM/0ddcmaNhWLPtNcudLRYSUmF4HmSlAqNAoKnBk
Y9cqMYDkeOf6fmgJzpkg1weGYUVxTtk9paSd4+ljM8ufRtxxbP4RYYg+URLnDBFX6TP/1s4d787Z
oBMZyTldNzljOP84X2Fm9PNscHBANpM7hWLTIojWNNZtm65gJjovrmd9sHdnE+y6g1UmC0PtQ3jX
JlgZPrhnO4Ts5pvQpHojqwU0ItMurtrRVPpD533vkKPeUDWr4g7UCD20objSj/ZhZNlBVUfslkaQ
50swej/v1IJZsA2hvFvWGFVJKUANPtVf7GX4tovVAVGVwyvpAgVmfMeYMtfixdQP33Myzn9EQjRK
gFIkyMR3bPittVsf1bQ5YFLkAfp+yAuH2yoGI3v4Z1Le3OguEDKUkl5DX0sQLM/HEHbjHbYHL7Cz
0OMcEe1sUuLMQHYSKqTJ7HePL1Q26rS2MxB2RG6VQH2xGQ2NXmUttEVE066uOnlyf+EAY8ulqv2K
/MyJyJISpPthwtgP+92uv+ZM07vaoPNv6aiCZCGQUBpLYtWp+5XoQ8ELvBX1mgfuGwrSwcBsjh79
CXDfvvqOHfx4U8rMKVIE/sA5cdUtGvMJhyN7A69apIvFC672xb2IYNB8p2PVzq7GVEi20mqa+880
YS/5NifMhZzJEUTrbfZfIBzDaJ2npvz8E39JchIsqO7/PjSjvFMDNM8iCvWH725dChYY2U5e7IJ+
iywkRmDSBxe10Thf3GIr8GeC/pOYN6DuhOvtLsq8ScLyrjICZGqa8WjQ26JkhV46EaSLs5ieSarx
NMyY1LNZyWWyK+U2YFPcZg+IDUbsJdyQBm+llmBUHuXQYkjcCzii7gJ0ukkBntvQMqCMXsJmmS/s
oxiGOZ/mdKTGvubGYlXqpI5FBy1Tu4DzrIFrRma28l3I8dMShb0eaT7mqeCRRYIUDuyzkrqiYZVd
gYrMkimN8tz/Ddjyp3MZNtCeEl0cEs+6VdYiO3Rw4Fx/X0vtxhYMrWtXCVjmIB2J7X+XBt3zpDld
VHZJnYWaNsMoWXr6i27JGKbcSq/VyvGeciRtYAV5lhNRGpLef+b7rrX5Cs9J33JzFtzNdtP62DXr
mJjAyCY0lVmuCUrz0PTnN1HXVV/42v5Ua8+AHhS97nTLLJTSwzXiEbOBuudh+eKaEniI1F9K6x18
BfwZw+rF6ybwWqpdhxAH+XxQjjROm6fdYR1tHuFQeU+ay0KLjDUwnhjyzmYfgaFJLPfAyMIHHOCY
pSXa+1KO+lfuVFjrqRLfeGcWxHdBJW67iIuBMm3a6YX/xXmTf6YbBi56hxp86xPPgZbmCMt3csl5
DT+ATWgJFuvEcIK7Sk79H+pad0LQi6kSQvQtl2qxEdbkO4QL16XdjhPHFC9COTKDQS1x1+Safrhk
w/QkMd+Qi5sUQLE1nFeXnFbpUrzr9TSvSZ2iIKuJKkKFaBw7xdf0V7raoASI6vmw+jIRO36h0QKG
8EkKljXgDT1SzZlSBzQPe2Ku37ffQvS8xW5FyTETaNdauK4yRDfUCp2HVFr7W0KMdr1k68Jxyp7h
FeT4Ta8CSi+MlUcHv2QjBHxNMIeXfavrqOTxVnGC15+nowS/6cpjKqwF+KAMLNDc0PMKSz8tGb8Z
if/zbFc7+QwV29VJg/xKzei2EGp9NEpienAgzsyXEUmhVujbu0xo6l+2/nv0gBNIjoSorkaDn1Se
PEbNJnPbxQ85nYReR3LjhVMWa/25J2ZtN/3HKCFw/FMF+sRpYfj9cKGkNIfRxBARk/i9Ss8pFNeL
gl7hwJ7JNNtGKA4GaSFVdxO54j4ifOi+6u0Dp6jbmPBvyXKcNdW8NvSa4BbjJ208a3n/8O9IGF0u
oKhf0aPEbu8HFES+LsmaRbW4H6cSSut+AECtW9H6vHT5VvIih9vrQiQ/Yvl0F3unAw2lG5ZwtXpe
Be1hV78TR5fOX73MT+CKroehWnS07dhoEjVQXbPV05OWcoynJ0J9eGZcyM7lpMJrHCdVPlZ3JIPD
IUS5PZ1DLhD0duBswMGC1411cxsUqBBFowYN8zmPO36qcLQIhMnK2adn/NFZ8lgR2EvJVI5heavC
fwY4fK1tJ0F0Gr54W0bRUmi1vktSaS6wUjDZ1yMhKCnkra8upMnXoPvQrsrLMeOlTqCgSfwEYucr
Q9HHkVn3aFarFd+bavUHyIvpaCuoicmHTURbMwbdkWaMaWqMjT6ST9p+MR7t85jCircmpzYzHOL0
6DR5C+CQzt/f+QC/sDqCfFoUIuTtPj2EAUzBKIarD1pVWlG3xZJu9kngONvL37L7LnDBbi1fZOmd
l6fdDySBJGT4mojQN5RJLcDLDnCDRrINJU/xMrFXNgFm1EqXEfN+aKL0ArVUTQEjpkrg0Gg+3aSl
fBX9Dxy7+hMqdGoiNw3A0xWuHJXkAcXmrKd3K6r+Xg890A0UFfm/OF2/K8CUMM0K6p5BzTsUxCwm
QvGcbvNUBKFHF3ehUXMmmJKNTupnM1jQaiNqfeqAG66ta55i2w0lDKDavWszW2ovQN9kjngqFJkV
Sm/xsfh/H8YSK2k9sgSqpt3ysmXHRkmdlnViNqRMqPCwMdoPu073zvFspR0yzs2F8JiuGWs5wfoh
7uvIqI6E21O9ZMGFiLz+/5nvZPkgWlbwt5qeTkeq16LQ+evPvEu5kiMWVlHG9hGDGaNa7jL4OSSB
1Cl3tF6K0yNvwAg0pBup0aSWvz9eF2DKOqT0iA+Ib1UWD29HH0g4hVizlVTsjzzVosrRl8DuGq5B
rb5+zYjYMgC+B2OA31lsv699rcyqJDfvrBYBEfijJ1hHQBLCjpeOK9JAp1SWKm+HYSKZGssvmXtF
prQBjyn9S5O0H5FhHVgUWZdZIReIgdqyQZKECUcr7auYUXXXmDYboobUL3pijscGtXgOfzGqAJ1s
E/O+z57+lK+XQSWeEZzu0TSdf04IOUxDGGTIFWPTs20k9arrISkwpvuAiFrFeoXE/JPPGAlwpLnE
dHoW6Y+AJke7SInwNGxL6Xp8wkaIJRVgHUsjxJ0t3baFETno9ruyrbQhswz8Nevo8NrQ0jfyK7/k
wP10j2RVF483nVWDQ8HjQ+tlI1UIRvVR9BNOd13+Odq/xz0TVPbOxH2Cz93AjLVlOqpANNhRvclX
UQZgWnXkLcgisa+xV/eVKLhR9/i1oULcQg55fUpDcaPVtD7hMZjuaN1nzZxcFsGlgFNmx0A9a2tm
8Cyc3QhLlSVrp4bOQnthArRwkEzpRSK874NiWjb5VAOYY9vLQaV6MfUNdlyx8Wv5O1LxljZTHVXe
lRn6u+SyS0er1mQDlv1sxjxuoNs6lUrWifdkFijJ0ND+Utvy4pRaTgN5cG7F2JoykLayEQFl2UQ9
gESZIB3E/3Fm3lRCPLbN0PkSSvux4umrd6w1lUB0i0jKu8xLHKERxquCn3oEKCRV3r+7qrLAqwvT
FtS1PAdoDqudi3TlloZYQ+/McDmA3lJnfG268pVgUN0EaZg3B2EYrIDzIXfwP3GE1JnUy3aGY8VK
/MjJo7Z6nDOE/PfxEvp7Qfn9f8fi2IjuAYwsjoMh1yzivTKAejJlrz8+8NGTxaz4Cn0QrwNW3okJ
whBfkNBE1PH4ThJSbgKw9lvAnzX8sXlSpakb8AJHe7FsGTjcWABPpf1QXm7v6KwztPkTbpMslhNn
S/w85Wxk2Z0/RAOBT42otrnrWPKvhbQl2L6UaJXrCy1syb0l9bPaqecWG8lwcn8l8imrwyUdg+2E
V1ZLuQBkU4BQikgjbttpqS4rrVJnPcKF5ZHZ+a1LyRmxyQdiYGNIaqebiOUwuMXUGwkmnLr+pf3z
2ONuSk2mHyI+acBWhSIL+xSZu260cNg00jjf6tcPj6G31cDT6XEoO+3P1p3cVJwyu/WbM+ydfpww
GZsRZhBNXpkDJncPimvL8T09P/vH0yv0VGTB7ZZ9z9KkXXhwgXVnk7OkPPW1BgazmjvrrheWI6GK
n3LPFN3ZeYN+7oCjGWMzs20E4iHx/A7C/cL6ZSwNe5EN6cNeCWVkh/AbnR0/nCgEt4XwFexC7YIS
ToHLuHXjTBm6prMMKpR1CZHYP2+Yf+Cs2UsEi2L6vmkYR2BYPGG2YYhQ+i+fPJ34/4m2mPNhagAh
clhgIdfsNe+qiID3MwKoGIEZc+D7/5w1OSBEmV+ICGUXkt4Xh6+cZxriLOamrmkERmjJMmkw5eWy
3avQD2LEbV2FOcYVxY+kz1Ka/V+liBuGiukYUB2mfdpXQQpI+5x7VkGX17jti6vNnY5GCloCb9YZ
V5SZbMblIIaMBtsZg6W8pnLmYcWjqPJulT4q1qeI4vcnwDIHgRgJwuqpOB3ycTP/q8ZhMdN2DaQT
WGEoHQBKj5eqSLml0UBdFLgH/E+rDZBB4h45grmx+GDhjO1p3MCChF1FWuctVUCBjd/CtcKZ9GQo
fGepmzlKjLBXNVFy9b9vZgCmboXXQkFA1rJyQnIDRZZklaML8FEmaIj7CnYpC27b9F3RzEBm/38O
fUrKQ+vhw2Q80RP5ahPOrsPCuS5VocxynQXz/ds3UzFk9Z0DZtZFJvRzIq5UMIJWfaqrM7xzxPaH
S81efXc+qU/pVtB+iNskj3FC63Il+FijlGp0n3LBGQRf785GLzOBrBla0DI6nGL2q2TABhJlAxv2
331HHwncTt6fatkJP83y9LAw1c4TLeXZ+V9NGCl9IDblSQ1PgSNqynNKj+EHDu/OJrRSdcpenRPX
nGQU441YxEFcnLh1AQNpo7dlKBdwbtEv74L9lglBif2gelfRMdmb0urOj3wlv+gO9jFjKAQBDNet
fqzdfH8TexXezDoM/gQgcIIepHcpeCTsEYweiElREBhABUwo549hrIzWlisd4iD+elJu8a38YXce
CvTeg/Tjwg+rWpyGO2w2JvZcYIaLsnaAlKVWih9OR8Mf0+Vsg0z/n8HL7mIUIHwnzYW6/mSyF2g0
TvRjX/NLfyXX3Yv491rDQwkjdyDFe3nzw750c/98eGkiE3MJW8QKgg882JZqtvrDByK7zQONlZ5P
7Ja/YiElxtlbrTQIJ081AfeajnlexHK+IEtOAi65bpOo0GMdfOXt5WrHioQ5HlAPY1sK3ty2jOpF
3zuU9UCuibArIHQjHWBldnujivDOWeot0KuyMqjiYXFh0u6g6LjuMTo6mdh2Evu74SERKuBUY72x
2JHlAKh7luttdbYUKLbYKFTabhjb3fp1xdsppeqj/58DENIoL4gYaxgcPAzy0Gzhtr9H11swbMIq
JlEVEHsXMafWZNt4srgwzvvaVP+emSt3FdKIMyyIlCWUwUNmaYnElQCTUKDcjqYBZvJkaYjr+8o0
Ujo1hW5UW5aVvdTgzuTNG4tBP1XH+BW9AnqyLzMOTLVwc4G6qB9oYr5r9p2io3ZjZuA8erDcOS/A
hS2XFh7lYLxzkHxTsuLmAnNXh+YWFZwU6LHaJnkW3BKBrHvklTgK7detUaJM/tWOmDK5jQr0QzVO
E2TPnQtvb/To98m3+bVH7eQlkjOzpdDIhb8Hv7H9zwWiMnf7pg+62zpH4I/pTI71xwYHhjz3iZ6X
AcjAF84n7MBfrqQMHbHcRQPO2tB3uUJwJUCsjOOarSNxYjupIGzwA+kuslNwUgDIJyUwuBRXgE/a
TS5sEXBx8FZ2VX6NUCpEdjHR/29VrVb/TIdx5G2OMWJqNmolF/L1STxZVsVZRqToAahH9HjwXRP9
YeK/t9jSDVYiVZpdKLVtMmLMlvF1ULngyQ/aT1eRVypAymqFkw/yNbbyztScw4RMULhV3iP4U6Fb
Z8MeZx2fxoy4AMpKpfOTLWNZTeED5L94aV8UdKD8HjPZ6DmZ0JUBVHkt4UqnmytkMI4m4HFzVtT5
+Na7cQCj7qze3nHUJa6AJCNqLO5T84LttpYaDwKKrXLDhHC1QKnWQqLl3mdGD8Un2o0GQUfPmioi
Hv/h6nfP2cZWwSXERRYZ9SkOO52HLJpgL5PEkF+EQC/BUeqLu6zxVfApdkheTvkJq4GPCRumegd8
bS8zA92U85O9DQVdEeF7n4qqb+mxOxOXbvok+tk85V7R4twvAAgLaSvjQYQ1ufLFzHI2RU5H4O4P
4LJagf1b/xVricpqyRNHm7WxVjm9/NWUxubZJZvztAaCCy8wj/ERtiS6+k9Uu46oXoS79L/8etq2
8DR88WFoFgNhrPF3zNLYIG31UifApeo4GOijMsGockeMPcBzBbeuFtxlwPOHVCujQ88OLw+0d3Wt
DxdG212Hhl0D8+RO6tFjHbDcMr3tv2dttlirr+4LQUcBwFvnvHXJA4jZk0YpDz3TX/aczlE/qDXz
ZAp+y1CK5PexsxM92V0aoHInYNNzOhty5oFa25h4u4QHCLNNtt2kzT5fwGpHqa82bVPDV2h33EQs
LJYtMAoyeJwQ8TxynLdNJoew7UYzNlCmlBcWB3M46o9i41vUaiPuhIYqKAzQ2ZqlmtFu0kU+fudo
Hrbp1GuQB3NJzdlOZZiX7yFC+v6howRXT18/rp8J6CYeZRU6oqmWnWSIzocwDnzo6G1jlmzKE26O
3m9Fu0KrnpGXYK5zvhapW4QAci9nAzfEzUqOpJe8eIu5n77UNedJBIdvkmmpatNptp2xfLBxLcRT
DbkgtwP1Wo7VMMlPMc07YQ+pQCiNgHfRUydGb5+XzsTIx5NOnKH/vxnkJdb1QXhBoVm8RXELk227
oXplWw+Qs6wJfQrOwsh7YbULmVAR7+LI/43bl79X20xj+S+RdxxPuzkNgGSWNMEAIYRAWAMhk55Q
CUyy1ld9bO2cW3njvq1yGgYWxKtDT22dumGBPu4Bma4+q5oKIGu56fjB9S739K7z1dX5NY24rsja
FZKWS84jdDTQXcuu5OImnuWvqJ9W5IExQdbeXCMqOB/VAcCdJo2SH2XYApZShga9GDePDD8/rvec
ipRziF3qgmRAofjeIPVD/GmeXJaP76qRluUl9Tw5O7seUVSYjnwLQUE2+y04XqPcbcQ2rCMfZQc8
DQmBwwcwCdln+a+hWJ3DHHczHWu8pigetHmeKuVHnz5aSyiWHQ0siwhcQOkvbuqGbajg9SNsSRrg
xkg7zkCoLp8zxzT9TcT6GHD8jcfAlg0dyvbayXY/dA3GWLQI+ZME8VG9Hd+2kH0yBEN4LSznkMaw
vhWmiEQ2Jum8Sv741tD0d5VLRNjfNiDIkfkBMpBQoHpWkyQsgO8D3vc0TCpoKVCaacyboPqDpixI
ks08/yUqqvWnReohcbIAX5oeySgJEnY8uNi35naDTm9qcYzUVWkA/rrB188G4mTiseIix5Mbd36c
ungcAWy/yVp8ZU3lVXRuj0yQ51psea5jRCptl3SP7YMX1jcK+gcUZfr93jBCsrLSO3z6MBQWnq42
mVWxuOVQKEJx3om9SEXm3JX+iRyGFhCiREuQdHtK+0IsTTNOe9hynQtFUKSfZReczGclYlDHxZjy
lfuV01oUNsKgMYaM/tjHYNeYQdMKGdYTJ7QXIzSHa6XZSOVVsoOx28o8yZe45t5rv+3zxQ1ar9Fm
8RSxUZdmtFJN9qXtGeUc+sOvCmEDUFLVq/v59GiR1l69TytoPRHR39/IjuEVZ5d1zuf3fFN+z1Ud
uPrma8tDecAFGREpe78B79cGXzhCu/3R+yJhZ7bMMGJ71UF6bsdxX2uvz/HU8q8b3qMBGaGUBrmo
aeHTQA+Z9faJjBkx9PR3ZOYbbsOkqub7PWl7xM8WY22rgsz/ADDLGxmKA4Fs62Rt4pfILrCrx24C
O3Qa6I/fw3AYh0nANgJCfwhAEC/U/xunawZii66FXEsNGUD4Kf1xaqWB1X39x26WCIfO+eq5QMD6
WMlK2+rw4szEqIQXccBhgSIyhjqv2qAXmgfO89NJQzgNXPWUt/KU0tmQVMqE5tww6vsYxH8rjJUC
DIryOZjLx7fn8QAlAc14h1irwnxEq/ENPtY7AiU6G11+kzp6lBEPy8hRo27DklkAhNkmpJTTgckz
HtLmIjq1HaJSZqr8+5Iuh5F0pY65Cy/oQHWUPNVTXPpbYOtSEXzCNrGdT3C2Y+80cYgKfHM007kb
tXVF5wdIpu7S7LbCVRiWdkK/p8bxZ5L/kEqLusNVVpUd29WB9HG6PnIigF0H9yoMda993cROr7Rx
M3N5mqx7oPvH8FWTqygWV4BCsdL631qAAexhsN+LXUWwjk4ocXOMTHAR9KhR4JUEufPtuQaQakeL
PvcotNsTjUoJDAMVqofbnOuy7k4XSczH1Qi5Dl5WlwxkwKtrpRKO1Mauuuy/TIxPUKz5YJqo4Cfk
ARj1VRpSpOY97MQI3jt1HLhBw5MkR+U3vBLaivPYKdF9RxZqH70XH2E6whHoUR856huxjgUUVcEW
csRB60QL+1lzVkoLLsIej5PfBcGKu1zljb0QaA/QP5ErXSQt9rATmlQHaih/4VSAs8Akqrp7yFMh
L5nSdPUjwpQ01oAlBIl88dV0qNPesQwrrpCW3QR1KIOi6yeLI/YQFpacAcngsAmoNXL4qXImammP
ujB5HIHVDj1wjuoSC6xX+tlnfn1xkVfWHDeYKwVFxt/CBs1j/JmvSrEwoT24Cvy/gxVc/5XRvXaV
jBylTsegX7NzK2GmCaJF1JVo+vfcOwQv3+rswW0F2717a3XgDG/m2OkN0qMDyD58+rRfwFgfINwT
vyRXd2CKZvpOAPbPkWMwCy5CE57tSOSh6hpm6VEHQ0voATE42nKWZGggsMp3MpszpKHI1viPfPva
H0w1uFK1JKN91t4v30bJphSUgYc/kDcWq3f7GjK0BVSAchfl4GAqEgaGdlWLLsuaC+XKjm5YSfdL
/pao10YQsHoTavPwGZCds4M43DpNsLomxABRtvTMbtXM2FkvcIlUC35m4FZLXelvqEmUE6skEC4j
q3zL7bqNI6wAPZobMBk4/5fhjKMLISmxv8cri+vAZit7EF1CSSkE9kZG53K5GO4/i9PVbs9CV72a
DPbum4D8yJeBnxbmZwQqZkYZmin2gNe1j4NSyAp/FHCm+B93d09zoSVVX7MTwusf2VtMrWtCIweU
aASkXYRp/CSRgL0ZHJH1qR8stUIvoNc59SWgHstAtRdNpzCd0ApOlnfNpKEdtGepEfUsvQ39Y/RU
4e96Mut7H2OjKxqoQhAV85lXDgTW+MSFxbsj61dLiIXNz8yaJpRR9J7ab9jpwdVnEd7NIB3ywCmZ
hvipWA65xpFhtdTdik/s3q9MQ7qDeYJ6sCfkgWE7miSYiw2cd0MQk65rinx9qeCD9whmmSGvD7og
dTEQeZw604+nJJ1kP4c9wDEXAwMPEV4JltG1pwcV6lqdPOkDEUexoQDc+VqlhyhW//ZICV5hYApI
jTjJoEVd9mFxc3kMDvCQN8Fe/tKQdeqx8lXSaPAF+liTTOMXev3rqKjC3x1tflWbLM1JvopXHDVa
KkINUNt6/bSdz9QnbhSQgEVjNkM4KGDputxmmo4JwdEsAuNbSnzu0O2aylEjqfcARH8Z6sbdH9cB
zyiN0QjIEJDehaTHZjz48e4/78geyKIcTWSlvaCdsb4xs1R1LPCcqF6vOcYHs+JNbKXEHYjjlDvp
CZjVaFQFYrBO8lw+Yt/CfZn2Uicl3EfKcZCF6486FsjUPJy/Iwt9tMh0AlilmyCOXGS63vjllei8
UiDhQNpCfUTEtn58Qqqs1oZHb5BlEzENqeWgqtauvRytsKNd9BLzZ0pX5iPRKTHaURRZEpJF33vp
dZud16jJ+zJjQeu728mw/mVUpdC96cnO04gid/4o7yh/QckQZ9l3zjDtWeFGS7CbHySD81571RKi
uc3u7RbwZuW6kR34Id+aS8t8VJnyzhv60gESEauBor0fo43RNzOfjfnsF6bWodcj48zfixNAzV5o
RqOqHqJ5LgsmoyGG1TvirnyOMqnzF9mly137xVia7yCT+u1EdXspl7qnhu4Mm3DPHjbVECNMT/aF
WHFRMDBlsZx6f+7MfkN8K+Hbq44wum+N4RLGvU2zRuEzqIfgea4eYDTq1NiKvMmGzoZqKind63wk
HSOjFZLGvliSD52Z4qH2+KI1HfhT1lDIcS2MXBzCwmqFKG5CcopM43t9/tbE9vdgIo4ndXv42N3m
9UCl6eieADcVj/zVGn0VaHkvuZ2XnTaRPkeXuQWXAgkmj8ixj/2XrcC8PgoASvtEllPS4oMLBQ87
yyFiFgHWXMNqCxKp4WKRde/Bply7H0fE2jL5+9JYiW0rkMH/OUdtnO4Le2DZ3kNnfpv/rUaayYdZ
zFCmWfk6LSUF2g6Hf1bpyQvo7aOs4SGOVAU4p+64T1hFnBySGl1+1OCzCkOi8/Wn9j32gmvOGjxI
gzdPfxR4YppSgCwQ5fM6CpQCeQl7vT1LIs7fkEF0Ws2agalMXd0yjoZlpz8boNI2AciZ/QZDxtGx
LkVjTVdEtE8nrgNDQNtmpjUTKfbsEvQVqOIw4MTYj/oWoCAPk61UOZnrM1EA5NUV05nxqp/SgQoU
VYuACQPjrfgk7LGH87Cf0HH/xckNzfEUZTKT+jdmrZKBFvk7H8gRBE/14x+rU2mcaZsPyHxjzJNh
3A8ONBt8OtzjNbBd7VxzXU463oBcQfPWUebjqtSMjM4OMZkWIObN0P3pLW66z5RbrzhhhEwUTcWs
9LV0jxPVURk2E0n95rp2Iw+2tR4qzWrxHNg2e8oKgvQHwUUpZ4s8XFp6ZYvGPVdpFN43PS8Ia2KZ
xVD/uAc4Af4gE2V3hNuhRQW+uGuUDrDKiJozQEc8HMFg4yj5k5Zwib0cYzmsS9Hf+AGztXZMdM1I
Yfqtj9H+FG7kRVNeGnX9IfqHIG6hMTX27/GNyOsBgkruE9VZvJR6DqfbiDq8MXpMPpJTqfaPBOam
Hcj+U+0Dw2B2ORUokeeB6sTa9LEBhNgkRh8P2J6XuBO9kjrv8GJ9adQxLVsyI4w4hy/AN1x59rTm
0PZfKassi9FQfKoRc78gu2JiExkBFVuN2uC3o+1tO0jsT6LE9QqJj55fHD83Hlh2AXGWedlJ3LQ5
dLBkQg0MMNXMjxw1tVFnb8V7zIemiKVjYgBRw6VSx+lBD8vy1qP1OJs5519/Hc/BWOivFHBMKQBc
toIa23BhtqxloyaA2+0cWsLqnPgekw6hPlm0+PeqxD56SS671adwoN7o+7GTX1BMcc20S9I2pK7b
JdKVf23A8z9XSOmJjq4CE58NqerShrmTGqAXFxRzzifqW3HbedwD9YFzciwHc2YSQCGSRcFrla+V
P9L29zvT6QSRfjajhVrKPB8F4jbn74ATRmrulG0BJTk4AnHOYcap1FA9wz7ytbwXqR+Dyq9y9GFK
a/+WgmUBqgOYtYh4t4lmJy2NrtIkYMUOEOnCkzT1o1MGHWaT1F3iS8nmsOLOndXlIQBoF7yXpcrt
kywbIHha40g/7gJODFtBpHfETKnv6xOAAcOWseFBNhoBRYy0QjfLyjwl9wXiZzl89ftkaSS/dmCN
hwqBp15+54sgQ4xNfnSRYu4WfDBVHSPsrp0bc7Oc81j8FG7yFWl00+rYF8LRb6I+s5/WZL55SGHl
dlM1Kjp6E+uwFgJFpgSXq+7EaOgznAYwFJfvxeVUw6KeHnAnzb1WlsTtDN/jIB4QnxOdeZ3PiKyy
cHGrRyGCscc7XweQ/VWoXscFpeusOJGwaFEliTjGOM/cuhlmrYbTqNKLtqYUuzMUzfNnRcYLTGG0
aP7FkSKhoeLjHM+hhpVnrKwAvOtZZ+buEU81joTi/u3iBwLo8rhgJTltTapxr7H+F5eiAlcrcIiu
3HZVuQVlxWnFgkExGa+w0v2jsQTsgsGWChA1SpQjyGPtVLW43lp5NQgZUDF1lrsoknjozbphKsW+
R94RqpI1c0DwfrdQDfshVAlkwbIXL0BprFsypt4KcK187dXsFQLQTtCj3W725RGpadosvWLeU6rd
YX4kng4nptB9YrGyINHJ0lV00bcMmCJLNfNzFSPXI8zWimOE/njKqOD1biZKrNNRNM9oKKWKrze9
4ub7VzOwonYheNwNPFZATCXcPK7o5OUwV7WFTwOALXjTjXiI/OUs26LsbtLew0wkegIsVn6Lcz5l
YOogJJtsGmKFItQo1HZ3M/E5sW83/0f4ADmUwluqOzvm4T4Flb1/XxpH3tZknZE1glB1ZZqcUIMX
mZTq6Wm3gud9tvsMLtmWQMYvxRuDyQhcUsinLm9YiRpPGoceJUu0lbAHUwiSeLzVNzAdlF4A83wF
VHx8SDzFlarYST8iyIEU1nqc44dnbHD7VWr/tz+HE2yh2VbHyBhpXsIXKXhWJDmv2p32ciEFrTdd
cJOAhPKmybkHmG0L9MwPrVvfeIppjrC2d6KqBcRuh1qEYDcHxyyz0I2U+asMuPT7w1n1h01KIFHi
4mre5ZnyJEZJbs8RuKR3mgaiWE+bZLHNn2pVcrESalz05EvnVI3pw6CsV33HNo8hohYBQ7zgsRqU
B0TSs6FDFSKqpPJj9L6n+AHUZRMNzE6kDPg2X/BgqXVX18yz0v0zXY0hVDEGgaTXEwhKkK6kJAah
aV6OhH6SMqFDfbBpbTk0x0kYM9RviCdFWZCBT3JT9qkBsunmzG22NE26WS2PlDt/R/bM8J/sY8ge
SFRNYp4e3dxel72UUevkzGEWEKngCjS6Bnypez9QEj+RZllx1imaJJmQr397N9UzFHD+2zacugOZ
dQVh/9WOLPu3SxTOCLzx8l71wLELfpgpDxEVEkdskvSzLG76SMmgVn9Erz4XbZe5z3sQod5pqEEm
zhk6W6/O65O++Sd43poglwkepIP87gbN4PjQbE817IMGNMmmebnZA1rx6yBjFHb99Brw/vO0tEOd
wGVqvP6CZ0a8wH5lFRuT2msIVKc6AaT6Sk/0tjkq6plXyW/1hvuVN2ff9Ym2+lAwKhY1RQW/mMc9
Gg+bUe49QNjOmBzyfkJrRuvsEvPqJlgDcWzSyHYH+Iz/TxL64jZZvmLKfkAbYA8Ks7+1FzZIImtL
zf/hG9NARTWhv5FaN6XEtsQndxUi7uFFHP19hs9eiwJq5BdQWRiOIZb+Jm9JUdvPgLMwyJmTjDeh
1atqDC2dfMHpG5RqnYyLyY8ksixXbsoh0CgE8XLzzc0INGSEljw7eyfYVRT27VBhmFOhZz86fWi4
NP6gKyp55Nm0DqxVU5mjKXISo1Yy8Cazb0EozeqiNb4FNkSnd/NPyHc1XdkENFqMqm/CrUbWu8Je
Lvu5XAauQWlWPjBpjKS/R2lZx6jszdUE4sMUrWBFeX4h1EvaQiexJ3nRsJeNxG20TC0RwDTrYknN
fvvyBoHn/lIrtNCq/XNWiVlNz5jQ7XGyOTwactJJy49Z5HWjhCEwLzJFyR5uRjiP1bLwoWJLOGw+
1u1w8Ri9ifZBVBwRYk5J/LjCzMhFjv7PrUmEf0RZbyU6wrSkFDgn7yp9IBr5kOnou9BwMbBgC2qE
oGbOK2q63fzaPwbp6qpXmxpHieH91nKulMH1ho0mxgFlJLzZzllesPNJZFWQFqRaRlNILTkl7NVl
IGaoclAq52R8bMQGxl+4dW84hM/AMP2oRCMVwp6Einp9c10a0u2VPg+dOfFb0T2Ormy7bOCvhFPQ
V9P0qzmp6rk7tEJlbsXUxn2SnPGMf6dIHN3JF6+W68faPT+E+yHZAIZKdPgG11KgsYjii/TOtwRD
L8Q8z1gMsfaChgvhitIZVjgybQDByrS2NdhkLdyeyil/V8882w3jflBIi4WwVqu8k9waRun3li2i
yb0ChBNpsvs4FMLKVrVx7GV8MeDiOnCjw1uiAyzmpu+Dmn6kt1xlrrOI/9mdqM7W+UVlPhO4cBxX
610KV3bcrL0tXLW3PKk7L1WC3d97+dc8lrDncfeBIukbXd4dqtqnBMi01lr2HZOrnNnON04lAJqx
dN2vHVbe1MsPm8l+v5YiDegAtleZbcl69bHscfH93wDuIymcerYd+9BCxwL7U1JPftq4QM5j059Y
c0YMUtrsOjjKI0ksXxQbLQXwDvcC+N5mZPaAr1X0Y/xt6Xs+mkzd4dFJ39Ys78gZJ2DkxrorYDRn
Ao8KfoXv96eZppFXLjRFmHJVwVVBRQ1krB7JdukKXiHY8VEmEsnIDAopcQw6464Lo0zUJ8U6UjZm
HUIO0CZsjCJ0EPrW5YSWpe23jYUsDiT0ikLZ+UhBdbAaVMraNYG5cpYt5gN6gJzX5CQPyjcs5Lkc
/N5cEmTtki9VDb8l3TcdXzpZVSD8yI0qevllgIVv5Zz2GngYvSEW8JVpV/MEPzbdaMegAHKiHqxH
Yv2Dc3YK/+IilnS4ZT5UqXfWUR2MAZ9iSOmyE+iZae0o9SK2boLfUvdfMRoGwUsAnn2lIJ+AkmjM
/Eq++7e5H0QWG0eYPAYiQ9N4x2kdpphEW7uXLBnhlQWcRIWYHp0hRiHHfRgb0vNKBIr5zE/0eh3F
SKnkqNV+Es5SsDI1vkPRQwlK1EQA77mYQXXAEe0OsgwvW8VGEwsZhX8nEqRvzr7QkoBYHA7IWfxG
n2oAN2jklO74Qdbrv++XBNUjmdXdthnzq8baDCVAI3OuPpcgR0UbVZah9DshRBzPmHx/mOeAKRUP
AiRgL0bT8L92Wnf+30dUn/6C3vRRTZK+i0Y7rbyjmU0wTCuveITC84VMQF55snQRMjcLptux18QE
V2IgRBNmTBn5Gr56KgyJg3Qy1fmZefRU82YUUlVnG3OsQv6LOtt+izL6EfcbsJJba1XxeZREMNCH
hnxBBq+fF3T61rPPWE0qxkrmcqAk7HKGnZeoWqyIAlnvFv7m5m6f+/kHKFTgJslDutFddZLDIru5
z42K20MqdsjyztwgrxIaDVppFT9Wq7sXxOQbbl+M9j03RMQdj2/jyiIetjUTNqUqoHK7wc5VfuhO
znxCunOyFniL0YHS7j17DeHb/+k2Ql+B+gQlukQh0Kzh/jXo3bcrZUBLDrgOoK1xgFzU9JSutkAf
6WiKjuCxeBSr3qJLXVyJfy74GHWNfwyGIg/OatbXh5CXrqC2gEuM/Yqd2v3iAt7LXCGzLQSZtiRL
/ghfYEJgKqxadg3YGH0S6Tfz+XRBjk7Qtjs5ICJdKBqj6D8sLizmLBcnreJg0/gfZUo61Qie8Oii
BfIMdALl6hWV0htkql97pZHHuIL1/msLze2WBcSKvZ0OBM4PKlVr3XpnnqfOszHmAHVFVZJ4QWIl
n+CURBlBrjvLMsJb47JojzyWDBB+sGiGqndkGFDGCRItCEEmVCvyirGVh4/11gyclA6xqULRgzg6
TTWjiL1RhMhOCTIXMj0HYai0KALKSse8/9DjCW9sKnPe73k+FlYkD4tpwVQiF2Lf2Iu+IK9GCf4X
DgWoQIfKeSB5XKn3oFeHbNs/Y2+yIQVhUivkLzn81fiBpsulxaqK6SfgBc3D90L9it6bMJgppybz
Tqs60U8dOtkB6vT3K51gV2dQfyDAQK7SBP78/7ybyzu9xsS4N6Z+CN4r8eG4c4wcvjugW7+wH6No
SpOsuqiKzV2rnD+EEkHNWxWDxjmH5KxWZDZfRwHTmIZ7yCxeIFDfvpsEOQCJol9psBToGWIn6I8e
swTKOLkSj+A7hDNyJyBVgBkrU761FnrDiBQ0bcbSi9fxMPa0uk43ovkmvsRM9Xd9n1YkciPOGoTm
/K+f4tIZKu9sTUpX/dGXaV9p3XNomOJNb+ovXWshj1/hYVztMubQvaXnuu/Yy9zN/3tA8js7AR2h
8J6CDQEJUlSmbR8Rh/dw35FSywLJIJ3pMhy7phVVUJnQCWpbdL2w/a4ZdTJNtQl8+cVKQ5P0qP4p
saugmoWjcMRXlpPfxp3rlEPPPW51ELagfIfEDDYQ1ThiTjf54NBO6XidfwFwdS0qIzXjrLbYxgzl
LbhVFzJ4GYn7k4E+ZCLqwTjh6ZRONHrFjq6DYwjwfkXz/LZzC4QT4jvoh0fJSe9Cg7L6TMso3yNI
ut6Hyfhw3/b1h6Ux8PkYRycbWyA6SYkD7eh2YVRUO1vdZRk5r4jcUEdwa2Rz0N4GJOA5TDoXWJ46
1ZxtIaXnbVceahNAtWXrmWcHEEKh9kEq9Er15T9bDLqe0BGewTTPC/GDKKOI3Hz1O4OfhiMffVLF
N18EOSBQlgW/onTDCzXnpErlxGYBq1AaNM2VMiD4xtgOr460BGz0a0EsRlfydtIT6dLhRSkfWQff
GqMimRwi22kclUefSH0AQB246el0pUGX1C/4dsevHX7AwVzPHrtlQ7yXMYCnSuL+9E3yCbCCHxtE
yS/cEbJKfQ2y2yLsQ4ukU0Yj5Kb4F4RgSNLzvk/4k08Xltmvl9YsUnrUSTcT5mUj+L2+i6roIuVM
JDulfV6Httb0O/7YhAVE0edX3RPVQoNHaxIIRua549MI07BfwqM80iplu2TP0cpc0Drrd2S1wNVp
K/PmnmUJP9CKgEs/ebNAHHqg1yheYCeH7+Pzbfj4dmY10i/+XpOtwxZCkSlNfk1nJHkBkSiNjIlE
T/mi1PVQWpxW09D7PZTWLB0yLINZL2eG+VKDror2/JHWo1uDQIXJLKnMUwRDdp7QcaHnGOyZ/LdT
ZZPbgCh1m4lcATUHqXNFBOYWDryIcXwJDWXNECVI4P/ZgKqBngKnDmhG/vDyMSS6vBjRoxx4Ul93
I9Jss1kVfzNmdozl2MwQSgRWSj9YXmSVqzdfjWtvJ6NrHw60+/YCZ3PixJ16K5SzwfHzkEILCj0E
hKmVWJNpaKap2Kid7+Ze7dWufTmqNftelo0hp/tO2GS17ktkaXE0dDmzmr8KRdY6Isgdb+IGb8Ws
uYxGUDjZm5csEZR4ZIUE/y0qJ+UXrzqMGvtJJCSnv+do5NtzF6Slduc8+WFONjkUnw6FzeJkT6al
RRCDQL/ZqcjXvlkRwXtnEP35tt2XMB+M19wLbfdF2Qmx8e2cPClkwvx+qyDZvKPgZa8kaT3M50CS
6HTPNns+pfJ0aQQ/jYkgt6dVn1+d7LxHu3dFYThFR3wgLwyNwM75wmYsUFtbRhoKAh9yEbtzWFYE
54reeLF9e5L9qq1TyavZk2P4k0XpjpjLSDm0jxU2HyNlks9JMwhxHFe2Btjd3qxN6d+Bf2FRTNnP
acBa1cEtWTNaa7Ns2m82N0m9meBb89h9mClTZWNLVJioE4W4HRXlozFsVGkWsjcacD7sboDlODmb
vHxbDVF4l8SpOihnx7az7s2hmZNugyi/lTzBKZM3FPvaUswyYJaG6VAWqH/BHGLTlEhokTszswT3
0TUpj2HmgnmBhmDPssoAa5MpvGSTdL5E6KY6wvwHmb5tjkRjqaY6VyXN+ugc/nL+494MBYldtskV
fOxoVDAWj9Hpr+H4DYdxiUwH25VR2i3jXcMoYb9Lo91yxERYma/xshB2xSAqILMdBWifu6q6zCHw
xuFSYsgNYWwklRU95ar6wrvcyxHUJ3X2eaEkpz5OikF6jPvGIbpDmEb0nsZH4C2nby8pYREW13R2
5SMFcxYYut+/yPlvYVAyH9guhQKC6kQfvf2iHbHXEyahK9DGMVhBh6Wrccd6I75laABXFEydyx06
aOoFhEalOtsgAvuyaVBnfV8NjljGQx7ZLqQKJMB+YJeOUonbb/XRWcCO5mZX8BDsOBUJDGrXX1YQ
GWgY441RjkNzaYUdEsDr/42PdfdRXlp2agtjhGlPzKhKaLujOPSgYJniJCMRHwjVIwncYT9m0BF8
BtpMMQx3QVMeUmDvCDsa5Dd9fjXLaoLMVE7XXPuvSpB8/3BxMzgCH7+arHi3UyIQEDyZUHmfm1kl
HHEt2/ZCASJHI5iqbMgIi19XSj/IBfqnulgA1c7Mr3iAMnt0W3CX+VJghmq6E2p9UkdWBpzMCTMH
y846R0q4Nl5UbiaZQNqJrY98qXHWNsCBzzF2qR7jMhH4G1DJcNu21T/Nv7uKWvgEvzLnhrAvB7qA
o65Zr4CgGS08nykv8pvjJ+ru1l2dYOa0tt3TUhgEgtuW/XeI7ZeVYjYgUttK0k7NbQ7Y0Tg8UhBT
4/Qaw2qQB5Fpv0YZ7nPT7R3BhHROoGs6kf6XCTGfy3kD6s5BNqTUGxUEPyvVjuetr7tQ8+XrxoQE
WZZ1rNU8Mm/JX6pz8WOCv7eBrZcyDb55nctP78p3AyiHfIx71pnHhBJwGgylgvumDCacaPapWFlS
5vFs3sYmtqQYYSdrVt3LnXWcCkSuoC6dSh12qQWvCRo5a489TBt6G9oOTZ8RSg5Kk39tA7WvEn6q
8z4Mq82Fropj2rHX88cmy2Pmno67BSLQVhtGy0ha5UUPKLHC1Wr5TywilLg2mKNY4G7VlOiWjPAQ
alFy5ROtgiUzCtI3p1x5w5sHoXX+qmgdLkT+LU0bWpU3Cmy2kKlFVfw+EQDjQvsO//ShyF8nUUmM
FB/w1JUhvPhoWkW7l1RU9fWs6eGihoanoXnE0vYc5s25A2Mlm5XR4t05spQsvvqwtF4h5qDcSN70
oCOIFs8zagyMDWt81LCbC/bko5T+WMHgI1eD/zldIPeLgo0T4M5hdPr/JVu0WCBtkJ1vqXzgil59
SL6VQG5G9/bNAg4Mt9HB5YgHakTrkvgYxHH/JRErJwuoocc8T3Cy1SnL22qVX+pxrGfhTPRf1VrJ
et/+AKq0NhcJl7XGwnLCV/jmVmqydOinYRgNAW7tZBWKLD5AfzbbvVQAiNLi2NrhEIW/QhdMLETu
Nf3n166Oui4VvD/rZWJxQm6a7b1aa1Xe0gSnUl09EmKYMX4NB+Oqs7zaqTLvFNCEfYj4+8mZPv/T
J3hC5vYZvbloBA0kqPyPS7DEGCRwMD+qGuak6//CjM/WzVS1cdFEgRyqE1JDEmVW43BLls2wx0zN
k+MnTQXzYQqIQ2wmeAqZRwYhmqCRTMiwU/XIh2V12hbSXRHJvzvMfmlL9lXS/NT4Hoq0bhtBE00O
Z/OY5eqKsN9eL3ofcRjVIuypo9UcaMUEfGoUehmTR6Q8qVApN6ybWAhwFVfdHiRzj2t049kvWvHU
8fjJw/IQ2JsaqK45ALJKHqzh2CoJpY78CP90B8Pl5Wegw2NIHemETJkHbdvDUEIV5fBsdKJ2N8rQ
kYTyjPoam00f3Zs1fGaLpu+a8qE4Q7HnaajpLBNaLGLymWpRFrYwOnizbs6q24J2PQ6KFKOj/XZv
9j2W/GXEonn1IkUGtpuz66uyUJfNKSiGHpSIgv343MkzROhhAvEPmWex2LYhADU1IPNz0c2JhCVY
waGUBmkaNuJ+6/s2UyiLNO7zjklJDc1S+XxK4aZUEEaVi043G3A91j0fcIErWzinO+fBxducFUk9
7/AM9LOp9qLHQHmCULvMZ96I2yneM3Bw/Yybu38E4KjVgZKhWFjc0o7UtHtsiCTE6qO5S53kxZgS
iSdNiqXPCayOaFYIxz1/vB/xxff2XCwKQF0jSS2aQxqMD0rkDiemHseTkDVHFYi8Aw215BApnjCW
y33AqoDB/vvmtzBcwoSap76O0s70mDN4Xwpl2ZVht1OtmJ2WUwEPr1FvozfsXY8eUIXySnp4Esw+
5tId7K3f+65Pyknuxnn2j4HUy7xmkW1239IivzMjrSTAJg94fr1EgSmMyEabdYfsxxAV2Y2QjEwJ
czs6Z+M7Y8zv2pUFPMC4mNNgkUfEQuHCaAr9mfy7/oqpEXG/bqqamf/5PCwffUFuHDDzVR61NtXM
f4td2aThsEGu4dwsuk8jBFqpTrH2l79vk6weJ4GSJcIZIxxUCYFYK/BgJm2a1ETEBrm3lLRI4G9E
QiFOdl20zMJNe1LdsKgmdkRE641Iwk2hNiYdU/0LHDEkAg77OlJSKKObjUWwEexEBTma2atFZeAM
djEWqjGjtbNHFH0Ki/uCKLMOaszyUkTwAkOekuw9MwQ/AjaSbJYnTqZLPKbger0kLlCIBXAo/szq
S83QXlSplYj1pcL2HX7uvDHFgNvn7K3QG8AP6qLJHKoPq+5EAIPiFaiNao3JvsWGQVMW5dGhlWRM
uNyIqdpMYp+dyz+iRCuNqauXAgyE7DWsDEklHx5KL4CRwB6ZRN9318j+AKWT7B65zTFPE+npbwt6
F+fEvoKsnLA+Wdn8aad2TFDzZqWabocMTg/CNMdGRMlwu7kpfP1WK/TGYyD/RxuELnx8Mb+b6zR7
OX1VhufuulYixPJLi4ZWfix6bi410TkjBaY++oItzjkF5JYHL1LM36ToC2et6K9Ooo2Mmf5/QYzl
zAmRy8Bh5EQuTYyGwYvVO8FhUYa9CTOPbPSA6iB/DPbMvT3rqdaAXBpPJFhG2deXfaGlAZiOqPOy
Eyyy1g5/XuDXaQraMvp7J/1Lc3RkpjxzmJzE1AvGzBDNzNmJTYM3YnchMilCBk4QN64649SI0w9L
2O3NcLbsNJ4+ghPFFStksbWPR2ZjwD9/VrauRSrfCaw/I7/0oohZPZC8psH8eFpX7nAKmQ8RUJaD
CctBxhf/dL7LEv6qWQKly7/LPBb8EdCxxsdQ+OBlXVpL1+G5K7Qps/cRpwf+faEzlGiN/BPaz2XV
e8rFjZrKIW0APLUO816t4uu3lW451SrNynEEtPStcwPz/Z6SVERGx6DXy6CmrEvkEw2EB8ttsyRJ
SXIL6tDyITPrIEiTdSoKE3b0od8XgO+xAIFwcIPp8TqOit/aJZ2Baxbd2djzKrSXKyK8s0d3J1xY
qnvod/OW5W4nZUubkNNkCl58qoNWrit+i9IeQ/KKLWDjbtUuy6t7w9rdtIC3yWgATjlPWAtUVSbS
k9+mhfnlaE7mU6ftF189M5n8wAr/xZmQ3xtkM+t+MVydahh0WAyPikWNsfjh/WVPtxyRC+jF66/j
+3x/cCUAiFUlj+LrmI3SAl6ABp+NkbevyRxnTRJB6RyHIouQ3FkpSfOJWZ9IhWwEpUmCaz2aJDdP
tBypQpGyx+lECtxxaMr8ENu2hC4tFNqtScsGW91cdIs4vfimryxLy64na84fnlQ8Ztab7MgJ+pa2
s2raY5Hummxxiu38u/lg3xvkRxJtProPIUQvZX1lEjFNYPBXO0fTXbXFG/j3CH2SxiwyJv7Hre+S
lNKAAbJ60I/ASBSK9X7KMLJrkgiwwrX6pC3VHuFvfpg/7GKuQu+pOUxzcVofca5yQDm14aL2wGHO
Kmwy96od1gN7+auc/n3xmoT3syvWrUPDcauzi1UmNSz2lU4M1gJiB/kpwAfh8GPZnilrn6QANzn8
zDUYV7Bk8PTGPvPTlJXTqBbbgeNdSF+oiDDOd0sasFwOnka8k8beoUJJuFsaz/MpXSDYUjG+k+mx
IeuuYdkezU5oNMYIwvXPh3j4sfqmD12ITB8FwNkHPB2lSDCpXGn0SgUtciT9QOkTkynT+3oqXyyA
MCKGIDAXeEc9UEU/zRQpqErXRAWcdMDQNfLLHZSBVHCw/x3Zc9AmTfnhVUhl0OELwuhy4dZKPuqz
4R19APFdho8D0s8cKTirqGADc4I1pSolkMYUa0DW3pWE+lVBwoiJ88/Ni+FvXUdnLjkXWjDqwrQK
UJiKpNAbzKl/HolwrovQUecsZnxBlLeSEzmSnMv541lOUaHfpAnD8J86EK5ZnxuSG9LxsJHa7JWG
R6PCP+zeQRSqT54VfOta/Cj8ZzppG8SsexGI+MN0Kql5QuSvMxFqzIrcjzODbeFitNiDlnuMYDyK
WinBIrrxGvz8ILi7IcZXsR/K6z8A68UVOeNqB1PydyArQN6UyTLX4ZCb9d1rPspfAGM7kgMCVJl7
ZhSuSzKAhuSjfzIi8SUuc8NxryuGP9F1eMROUYnGE3iFFpAL5kapbAI9W/TaS36fdqLzC24JSWVi
2+nHcPFwc54FqfdKKXFINs3uEn7/p1gE7xRqFs6lwIW1iwmNRLF2VQYMU3wXYO6PYEsHPTILRKF6
FtDreYdKqYqo6VYsanwvuo+9BrSQsZ2d+7RXXbflYn3Zn/UyrAAwB8y/HZQU5K78+bqerz+Se8mT
c3cQE/cveRks7hVvNFlRD5Yqk33ehgShpolv1ggEsJGgcHK+dQ/SWiLsmWc+fm8UXJUn2+YXCwgf
LSsbCNro8ZNi8i7DgreCqZVWufpESE1KTvfjbIIZrntvlmtphTyr/+LzT1N3o804HjiOajBp+K19
LTnXw4WI/L6Pr71xA0UwkL9kGkRAottyFlAP4hmNSpwGYbAsGoatHRTcnyVjlsVFHIjxBHHoGDFB
dhm6RPMrAUbZqu9EGbBcYqd1WObzYxl6iXGHOWbcVadUYmBWgask4RInY/o1tiQz2yAkLbyxKXYa
VEs1kgLX38r5S7VOODujGHU/tLEtlGmKzKaBWNw0J+GlXiKFUYuRjrHNnqiaqs8pYuq9/LRdou+9
Ic6PAH0kQy81EIGInCpKMLNrzKWm6nHEMiIvliuyCbkJr65S5a90vXf4Sl9LSi15gha9HxXYp3oW
65lKGKB1EIJCoOz0CDqrtIzMOlcF/PiZy2yw45a7iWQh1HDAwv8bODkSVrTgOoT47psbPCum2QBv
/Psn8KoDgMJ3Zrp6JKqDdBYty1dR8vSFVY5J0pAhrPwCoAQIRqxwmAdALwt/6R0ETqi6wRAkYhl+
7ZZGozPCW8WYH8vCv+I4YMfy4LonykdtfjcgwqeMmv5R8I7c2famTESETyFj2ZQm75dSUJECdkQT
26T4oBBVXdRu/LF1Xex0E5+QR7wYGRhsfGoOI7j9eN2QooSsfUWHA2M1wEcWGUuyiGd3f2Y/g/3u
C+vxvNjiQwc0oXylfpitfZpV8qcAmNqNLgY8ZCbP0Xjscx3VoDMzcUux56hlEk0t9Lvxwquj2ROJ
g7IRIeYIUXlNsMjRVhq8rB3M9xGmYP3DCMid38CT7rogCSNPk/4kQUS4QYxez2MTgPquhrRNd9Uu
SRI6nmUA5epgDPARDjX77/j98cTEoaZxf1qlWFLToKBpn8+H4E7n5tl9u452ZI9CVbVzo8J0Hrkg
XcZZFeHngzCDPux1HrdlQaUrI+45bVDyI9Y5G/ZymhMms94nLDFHSi1L5oW+JO6Igpv0b6CfWhdr
oe7vDhKMfaiZbD57Fcb1CTUYXZ3j1aKd6mVCnHZIDnmYwGS1JMNYowCqnfvbYxFi+sDBbL07hBdd
1dMc6xuXe0XLWd50ba43u2YN50a7cpFR70t9yy0sa57BYSS1vOUFjYFX35dL1w0FBJcJMgHTDtv/
zMDcIeBT99xvRFbJbmYAmmWSYE4kbv2nlllJHGdLxM9qW4zDLHoeao6Kq774cdhMio/QVZzA6h/J
Ilc1IbyOkfgGPmNFyuwcch0mV6oiI6AFA+Ng9MeWzq0S499HQgulSM/4jBBONEsUX7OMKopDz8e7
RGjXhTP08s9ej7GMpETZnD/48jsoj4CGtClqYHVJ1iRjZdgqYtUylR49ZfjYM3+dWEHNL7eExbQz
7arzN1PrUOPRk8vFNG82f3EEZZy93SyCcptE+ULS0+e9dxzWoZAnZtdoTlsDLc+1qSxJlNNh+eQ6
CiOi/eGPBMdQ6sj5L1lC4p2v8y+eiDB+3PE2FmsCBSU1L9RdT3JeIjm3VIpwxHiaWC9f6L6+DXXC
AE99yJbG4oO2bNHczNtEbuKPSnss7aRnsPyD3q+lyqlCeN8alJRBgLfMBxBXW3XBqF7ClXf4jB+o
D13284og5Q37OL0okNbLzvjEVPwyis5oCR2k0piGzCMd9rdXP9d1ML8khuwWKjj03r83KAlidRhf
kCj9ZSjSgCWjF+BSPz6c2sgfo9AILdyVEhg5TavDMLNU2vdgOQljinmgskeS3QS5ULyaCkru/DHB
RiZothG2h3ytu00HjcAejhKg9huWqdpxU1vKkhEcQpCyFCQGaRnzXDhjbnNH6rQ3Ch9j165t65zK
XIrKi7eCDdn5npeFbKDgXp4YpFRiRSMZUjYnOAcbBxpN5h4JX70pmsq1T3C/QBEDDhYPTD1SwpVA
5ctTUtQPHZr+WOy6qVPjhYpYoIjB/2bpTXWx6qbGnZzbk90aX84H7Tvlxv94zT2xN9kYAVxXsZFI
gIoOS9RzgISZWgA8ElLBNFPmCaHvFDeEg2SdbJJpmjZO3H2vCfKgRRuFWRAYXnmqhd9iZbJUOo8/
45n5oss6+WB3tbQBtMG5lMsVObFn9D8gbL9AsHr5Y3qqMGywvSOFkLq09xyp3FEIyILQ/DqYFFDf
Z8LU8iH3N7aGP5yx0QBGXzPoDO7kxPMmsRiNt1tIeq1A4cq7vai20q+OhPwxSUjPyhTG2Af5ENg1
o1VPZ9Ax76nDXZhNiT1g1QW96D34HhPBhyGBway8OMhtMkIU8UF2Tme8zOpDjO6dqdvHNZFp13sb
B5HhwvFf56mHA5Aq1RgwS+sFZo3mqdkraRkbNA9T8p4q5nNN7iwjdndRBXqj6cRBRFsQ5+NIqq2h
28VIdJNIFhlDNOW5On6uHW4U3XxvE2CGi/NRRkB0pk83OkaAuPkC0ddh/GhmigGV+7C9DBzDsH+7
uZSMFRVMAVMRM00H0ser3zn0Z5FJiFXRIUsF0NriokpQZkjCR6M++68EHAWkdakVxe3fR58bIz4M
w5eFP/QMpzPv7P3MYdjhWJvkc32hx0JGtGnTX3CkJD9sNSx4pYh7JJbegEWKR3Z3VMoogvDE/+4N
qnC9gJTLVir6UmMEv7fsHsLpcZfR4UtL7ikCqiy0NiAQa8KSFIdiQFpzbXLW0/mhx6KBEfD5uTpw
1lc353PCYELDDEBqBxwqa6EceQxSURLZsT8ZMKEw00If5ZTQ4anHRsDXDG8aQkmBMMxaAoib53Bn
R9WaJvSeKTU4IYDr8yRZXfV+pk5mKXshDYVXDJUZxTxKMkvPsqSxVJLWaoWF3DiWhzczXe/9OhI=
`pragma protect end_protected
