`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22432)
`pragma protect data_block
giGA109OWTgnmloyaK8oODsiRC9RZVQFcgf9mR/obyjke8kkfwHUD0rFD2w6Qg5sKJtvAY8b/b0q
V+Sa+ZX24LFU4BuS1vxLWFGohu1WaQVSB9HQcsOWHML849yQr1UuXHS1H7VUn17v0E61+/PqUzk1
X19/pJmyYW1BM5ZHOhJulHdCd99vhdUA5znwgIeL+qkiU0sf11eCHljau90FYmDoD5m6woWzKvoP
6gHK4sfqQrITuaqk25AtWPgKwR1csWbXynMZjHngIasrLf7+j7MenOsVBC5tWag1BnoBGzLC6HYN
Ye4DMn3prRMVDFy9rC5aGgkraDktLLRha0XxXzx156wHa8CnK0BS+sUhVnz7ozoxlQ9B0YG1AJsh
0le0wth/eSyck/S72O1pd6HhMswIMDoh0KbuijwuADOTQslv+ZfG04YPbWWhf5o/Jh9H7dRLJnab
0BY1H8NAcXfYPqXu9n6hj9YHYYhFaRs/0kERlfKQ79DoAQ0lsl+Vm4ztO/JQ82VJGz1zcdZrR832
oOC5pmWUN3PPgHBPAlUS5a+Iyi67iZKY9LmYcj9yuFuDTKmPHgXMT7sPaWIfhXmcGXmpwrwz3k8O
Cpy3BpcBg1VXzMuqfQG370opc+mTQFy/Z59qBpA25yxXOLvy/hH46tW3dSDASYGws+9qFTrKjag9
OWMbg9XEj1DV8SD3mh84UeZnMJ7xiZtO0UIKPvcie8UcW6Nei+6nLwHr4twwtGrtKo0oOUmpGHHg
R5baNwzX6S0gS+wOAWJK1gTBYBcpH62J/CZGUrMt/bRB7ggDs1OjJPmGI2NU/hpibNGAems3NcCU
ckfI+aqHKxHfsyKcZtTpdZ2gkyrM00ZepBA9f56XtrXg3frD2L3CU/248sXUqU4jTV4IASR2K/am
Uc8kYm+ttviNdOcXtyeXwo3W+Zp2179++Q9UWq3FkL0Wqu1KIeJUuqeizS+kw9NtczCTZjidC/s1
L0qUxM4DJ/rjWQaaaJTQiHAa9+cTJWLt2Ts5/QthQgX44m/4Pp9utsc4HGJmNCSN5n1qlAetsBLy
HLVUrCTAKgrXGigcDQNp/1Dxvc0Z1E3fRzPEwcVJD82ml6hm0g1WOF+Lk/eHmot6KSYhzz7mhliK
AUksJ6apco7WgC7PKVy2O1VxSm6qmRiTgfrsetNAxbvmVm90dAXYHp9zX2caW3sFr31GVc6nsoGt
x3lA7Xr7cp7NpjHEMkBfqXgmru1UqUGgyd9jH5WpIug5GPMa/BZ0LU387XsU+bpHxVf6LTbpziTH
kWaTYD3OvPXxhUeyzTiEO38WP2m5lBPzgoOzmd5vLIF22gpQCXEZxZlhzR/VlXZTBMU5y7Fd7Nr+
EvAWqrxpS2DYFv/o6eBO6UUwzkLPEGrMPYCuAK8AzppYe/q0rYwRGDP9FvV3QBhAu7aQhc4poowD
8xZm2IIoqMo7kAD9zQo2+yCw2ctKXf4gduWaE2ST6IgBPKgltabOTS7t8y0vLbbcsbPjVv3KHTa9
L/ZhXtee2lMhCYGBVT47sVwM5Z/bvRY06g34rlOcj80D85uAEVYSopmi3mmNu02AkPCFNEluGcOM
mur9J6sH/J3BlMLQhs1gmPDSWg9IAS4V1lKbSoeJEzhcZcdmqx/nFKYV2Ww+Xu5GnwxHyFNZCX4D
4PPWynFUul606O6Icq9SEBnVYzOsd/H9pGhYsxD4MLhPT6/1a7Ak5t8GU6feHNCsbjardZgoY0eF
9Bq/pEqx0+xAJy88vM+EDJIilY2UtVvzaQHM8UvypdSZRsDkvF6cn4B0BG/KVkSBMTjP/URhNTIG
W+3QibAPB9jQ5YU0dE/B7b/itOCfZ+JM/yX1FVV7kv7Z7ZvKZRyJTRnLZ2KaSI3JDZpI0VWafm+L
miT3C2P3544dAlzArNPGIyLWVr719+Jm3QYyKXhXb94SQEPOIOT6ze1vTh094gWgPKop5WYLc2Ce
z8nQyy5sXt4s2NtgAIOEl7Lqe6C48DbXfmSi23FmlZ2VEGLx/MA2r46cq43lIJQ2eWgwZzlTCcYz
tPAp3OW8Y2fGeyBLL0ONMkL4ZNHe9cMqJEHL7shwfOdgkuPjxl6VkjAs5Tkdz1+NTw55cyOZdFTx
l+Lo2qHRV6JNwmxd9mHzlRb8AJUopA1wJ+rtyQOxEL4jxarTEKLGDN/RQM8GK6MEC/brlQznrW2l
wNaCIJGjBDwqYM36DCxNroN2qGGvn1Tf9j0ietb8u3XOzWcNlR0In5w13tQVmZ9j3fU9LZvPZi92
IHwLUswAXtIS4yX82lidCcZXJDuc3SccBsyLfhmT7hF88bpDUMNpKa1deqX6Oh4+Ic6GCkur8KtR
xnLKCVCtQ4Lzb0MtdPbNLDZ+EtWNp9jkCdZviVRz4vQywySJ7p/ulE+Q2VQ3lOmQcgYdNXdmI+C0
oA6CfIT4y3D2cwjTcX3hpsEavEEuVEO45YNLnpgyjzqrV3CHbKTZJi0ZRNU/UT5TeD0iWzovkS1i
RVNiESBubBz77DLO9KJB1ixDKEkACL5aXi/02fnDA9LbH3tPbM23n05sjvqBPDN3pDfPGDX55zy3
61vvgtHLsqZNE0byRIqFyKBvmIkzrp8LVYuL/Pzupd6HOO7wVztA98m8zzBnInbsqgJJi2f7ZwZd
JEROzDdFqcqgyQZKCxsdUUL6o3kQgIoGRAoTz2Kf2yKmnUIaPtKSLpptW6vYfrkodjnlmgpB0jOF
V548xPFs6H9T4StgEu1aVdUDpNFCydyO4OGyGCdMVke/yZPUZRVsRJYz20WL115AMYUMPh0akQCg
OggdjSW0VD4/y3n7NMV39fpAW4m/imULCNJrjSIuvZB0YZjYZbHmYtbRXqopb1u0ZzjMW+2Or6it
GyotLH3PVF+sSLRajFjTmGG/Aus90GgipdN8p+Fnqw/23zH6Y639rVe2OiWyq3e99Om5A5P6gnQ0
H0WA0twRbp1VHXbyqGZqjiOsMUZRdA7QHNzF2AOP8C8NtEBIBkFJQWz1qM+oz6TPko0K19qLiMkT
6QiFgJGGSh5n4FstPDzAVANSMAaQeLjNUrv/RsHC6CoRALjX7wiKLJUjpoweQbXvpV7EzOGnjYIW
zK2SKAFJjGFAhNc2Akl29Fl+QkozqSfTsL5EIkJhnyA1gSiXKzUToXO/EEbdQx5WGmqAGCLcP0J3
MHOREGPFlsnqt44gtJqGuuVHlYM+qvkg/oWmA4d+F2YLiqan8lV5S0FmrxTY8j/86ulIIodwp+Df
Ir9SXIfUmjZhTWf2gmCyRETDct2Noc6FO7oUifZdB8tb4cLKKIT0fh7xabdpD4jgAhrFypMOz5ur
SmyMUxcUZNqDe+BXul1qKbyIRLvj6wA+KnMzLoo+dsOxhCOk21YyRuqZfCC83kioxLJvwth9Ehdh
ivKn+BW/iGTiXTemKzSJL1nq5OtGqLf9AaXLFv8dJCB2sJj0fb7VWQsWlqpLR+EVgXhwbx9Wq4y6
rreO8JA47Mq1YNJK5VOdpJMdC7RKewGR2wJEu+4Qe6B7nESszK6e3tc2J/v9+Own82FwW5EtjeoQ
7GqVJ1WLbQWOsN7GxCB8/SzpU5LItMK+GQYtcUtLVJsa+unvP+9JY7r0Mb4YyU93m8tMtkvg3q/Q
kDq4M+9unPR1FNStEBDIpOCGiP5rkgpYTNFheg2r2EqBzh32bIXyB5rj4OchoqhT62Bgsoe1MnxT
tPgs2kq+yYLzS2oRC2W8scxW1xPuEOWZMaTggt1gYNqI68CtgNokWjsJuGQ6zaO7gPh4wYwbrg+9
+vXXU9wDGDQBYNlOHoDXLN+KD/2q6j24a5yqpAfrqJCJDEbbtJQp9jYFuMwt9QlTq7pVqBdgE8yL
mx+DMfpoXG8lKhu5DDgMibFCvws2rmkHM2CAQDixUibiq6GvsBBELwpUnSs/RSc73DI5vXl1++hT
wy3RaFdaWqQRQ8P9w6XzTiSipYS0ngMpHEXMizjKR7UPWGmda/jPgPowruodkcqIbBzN2IPBrDBb
TUlw5bgeYr6EJ2XOp9YSQwrTkhvDoggwdKSA1lNJyXhMC/luWj7ua0kEgpVO1qrmIVuYMCYXGXUL
fqA3tBK3P9TjMu83kcUo9CpJg2NWehU0qwmA6GMku/i6a0nTbqaAhIKOpoRE6ig43KELkx41PJaZ
RslPdeKW3Pw+ZxM61Q1kTY4QmcIAodQ+JSWK7/TFm27gjiT6u5X5c7dG7agDItCl0wYR9GT2C+T3
x8OBdkVV0UPtqck13aTezPf+SwZn0RYwKeLdXBYoseZV9SozirfUZGRVu1jS34S0lFRAwz+vuQss
yk1FRl7XyKz29rkKOiAAc9YaUDiJYGl1yyea5cBbpfEo1CQ/JMfmg1czPsAgCm5bGx7Q6xtg4z/z
s1XsUGP8nv/4errkrg25qBU/oadnwkSCCHKdCfyqolq6kFlXFe2Jf/flw91ggsP458sTn+Zq+Ohg
BN9ziIuIH2JLDC9AWsQXEBRvOtL/wTze1ogHmAoD8QZ+UsOwIbkkE8SZHjgMPPc3O672gr6EZsgh
Ip+aI+iWhw5gmpBwWHdAroNI+1bLsrqeAk+RIL2vR+GYdXsjovmCf18jiirg+Y8sYVTH6p5NKD99
suo8FlTqppYo6v4S810zAKKkSZT1Rgu25Fl59MIbyJvY1SDwt1Vj/DgdKS/wNO386FChdhxrLuge
IIokxvlR53eHkJ+fF9YzZwM8DfMLQj+4qO7KW5csZI4GZ7FINN6RBBBFWoJ7gf7oMyapLY8r3xGE
PErGPdHt28LQl+0VFkhD8r+u7d3vIxhUQUlSJJJ4x1xJniNh7uuMrTMzba+66mIwQ2zlvvOh4D52
1RFugviUTWO7Kf/EJ5Pc32kU0tUoYqSeyZqYXtObn7a5XwHTRKxAN6mdjmnxLSqhwaBYU1umaA9M
HxC6DkvkKm8Cav9ks1OjRQEC1oy9/oxfeoN6e3j5/RVHTbHuATRApf90fP2k5+0gIGVH9rswrmdb
FIQB3fhVWRiy9FG9Sy01KUYzpFNYB7yTjfMlxyRL2A5w/TDH3vUhfvSEB21GCJch9C2asekZSECn
OoKDxagp895lD26/ijngMxIkojzpqCBDdQw6CXmrdoSC+3GXd/HBfLQDXpt3aCzy+fABJo0mGCLW
Av6OKlFaDVtziYO6lD5kGgQ7fY6XxfiQmTOIloEitfD9alwQkEniM3uymVtc6vSFwHW5lfxwZtDI
E8RMEWZb4pj62APTkAvAcUZrHC8eyERwJFDtVPWtqHPRHaEOS+t0eMaztHB5EuKzZ9QTX7GumLrl
xo9IBWVWtCBDDzU1NUtzbOloQVyFdQyPWWe0wB8VcVMGX87NsckOZNsDIlDn5dDuJYkEmAB70zyz
sMAoWrB17/jKwaONQkfjUV6+oR2fxQY0nfAyMsSL6mcyy/aQ/ZvcvlpsC6ucMZ7QzdhW1//yS3At
LQ/mUfSV7BFJzID3HM5E7aR2Vi3pjgqYFDtNtsL4ccY8MGYJYEW9axdcVjYodzAgL8LuwD+l90sp
PfDKGAU5+AktgXTCABpj3zznpkVkc77uWv2YjdLupONUppMAuQkF+dH3azRMD4N3tb1D8SFop0Xt
XnL9Jrn8yjtb1OZdz/FAjQpE68Q4pHb1QmCSKZWnIKfbfE+QvnuIxoBVNOV0qEDHiS88mhOjMkH9
lcr/cDEbNEJu29uJ495ec5gT6pDNL22oIYYVWJChrdD9fDVE4aMLxk3yt3trB5Ky05Ak6Km6Z49w
T5k2jOwstUEHG1J7Raa8PFXcSv5ZGPE+JvKSLnEhCbdMhvf22yORfrHKA7wtapHdgb5XgSvI3G6+
6MpkxmC5qr7848vdtKuHR+sXXGNi56BNHcTOZNv2/zWbfA2oH9Fobj7HCwoNOvAV+/BiBsul/3eW
idia1d0rCei0pjA1/T7dKyEwRulitbmEpynhyygEKP1UA8RpoO4QAykyqQ7LbTDQchA8ryEfaHcT
rndzbWmO7OOEZ9ouIefZQCJlnhopa76Q/0ZUiyb1B7QxpdBU7EZi9wSN7gF/JvqWXDhJttk1HakP
EKRSZHjnRww3imnLUK2yP4muXGQgFo6ChIG4PyAaZE7yAyGdxLGgnJMJK2FeEObrq8hUiU7sLiT/
f6qxrdKO9W6t7uPXPXrARqps2YTsLb4TEe/ES/4veYZ7mQMrLHP5GWgIUsf3iNwcfqEydYAwOPdg
yQlhbn4nBrnhyiLyYncevq26BkieLoOtcJ6AxB8SMQRkHejgg7di9ih0BXDoYLPtjbVD57elb2QC
u4ZNpXkLmq6X3kyEi3H2YF5G6LyNxiArLx6KKMSpheIkyrW8t9OisxHBwQBXiQFrgRcHXzj+S/8h
MaJ6P6srwwCJyOQU5hNTD+QWP3CfCVubhlSRY+JMrrwRyF+W/8vfJwh0+zsi8BfRD09Xdbo4nR2Y
9ytVhQLoptQ9UD1hNXgiYNwH8MSSB7wGQyQ3zgnZiy2ePPLNYhLgm3P0NKuCUKDf4pES8Y1acLvk
hEHfogJzmYodxJO0WmQtuddh+srwIZDdyHJFkk70whdR5NAe2QnLSJTktuh39ocbELOmI/KR2YjF
V+YSfGq1OyjUIvAsZD83yVTYyRALmHZl1/nGB3v7tZ7xuid4PN98XmKjspcddbw8t4laB/3UGP/c
TzAOLRnwAP9w18FN6bebbcyKF46Jy1BeZeBNjDzZljEkAoMaH/n5vPQFmfCmTDMrJ4fRs4CNarFj
Ps4A6nKvne6yyD/w1/dX45J2HHVD8NprblrfECwjpNYi/6kSG4Jog7aORufN1tmUQs6ybv53+hDz
I7uzIsxDY6GHIG2pF0ut8B/S8a8U4Z8fiPKmKcG8bL/uS1pzQIt168/mLGENrQwntRYpTEKmbzy1
7RcdBhRCoDclo/EIs+ShpHr9e6JNA+qi29TlwXlxrJpMWn1WfV4SVOgSner+xDxJCKm1Bin+njhg
AJEBTTx/bo1oAqHswsr1n+DYZNsG62GO6TC5ID1Gn7urojj2avLSk1ZBPX+Eqq3bV8mycTPQ0tcW
m1GELaVWH36IA0NcoYWRQW+nYWCsO701Ub0+5+R/G+z358CM+FwMJy1zdE8Nagutr8O99yBSEVbM
aKQ+iEStsvSgdoV0NrPYAEpiFg9vnzBTrDJjuEBbesQH6MIncJpaMKp6Bis6vxWwa5O5vzw2gRB/
9HHSFwaVMSfT/vYC2qJ347wI6EIgXfjthQPPDFQi3RrKybZE9p/vz1w18Gw27Se2kLSTTAwzUKHs
yU3T/guMFdFzNkZLokHWrhV5ykYNL6VG5zm+h7SiesRVrfwArWwagcETdtDwwAb68uAOcY3d0xnG
yzoxGU0pDo2g/tM/JXnzffgct/I/hG/E3T1oQmFoiWDtf+nPvnVhZIPn7mXFclU8iBa4hEqKcegq
FUL6ZODOPKWuUtWReeFV9eFYPUAeg5Prk2BjNCZ+CcQf+vRlkECObqSaxVebrbr4Njkb3bvjisRQ
0fd4s6PsQ+wKy/mL9EPLvDS8WB6DQEKiHU/LBpxIaCHUHZgHRP9Gkn18AWllF4eWBYIL8cqzCUwr
rzbW2tpgGvekcsOjYMy6LgEat68lWRlhljkcP+v/uwXiYbTwsCwa+IPFiOWLmD7HOtFN6/Koa59Q
PnqPa97RKY/vdwq63BNb6P1YOPWqUiSIWXTsvNh36gDPQvDc/ExR3pKckMJ1jRrd3BO156yx6R6k
lDip+pvmhySjuK22atuKXWCqbLINlc1NVkYf9kD0HH0pzArTnlPGomY06AhqKtJQb2drF4RgbYgJ
uPRVuKeKaig2Dy2383g45C4Nij7hGPNXdDbZsr2/CbRehAsA0cm2BH+eW1x+A5v1ZLOLwRCl1Et1
992mSdL94Yqx2rKHkuSovNLx0wAYh5s8BSCi4c09v2KeiQiv5kKc5qFm0gxVcnNAZgDPHCFKbzrV
of/8zX7w4au5KfUvJ+uhsOOghTyRDDZzpdT1IqaeSnVqsYkpYfaylShqJVPuKdTdGT0QKyCGIvPQ
hlMRabF58zVAYaEAZkgZb9BQ5q724rOPxbXTFVlG3sf9z3CDtE9fHpt//v3lxknoacxTToKOQdEj
uKNdlaXuYZWE3IzxlHjqa4qdROuqLAn3fzE9LI0g89L5pjXEaMZ3zgiw4IJpj9cZ1B4XcDgGU27Q
6K54Y+va5hO3bX9WLZNBGAHezDUrB6umZA9tuntk+8zRpfnPu62JFZmqkkGSEY3IE95orC1anIhF
N19O1eR2ZnLeqrFhLIPyOBHp5oIKbBf2B3ROEFmOjt2pbf5dud/c2jqWkjV/wZujmKhqN9aowiPp
Y4ycSZSBBXD+VBLBDPP6QQ1U6BvDjPSBN2e1YvldQlKIQUaDT2+MJl9ZOmtvvxZwR8GUFPg89nfk
gO8/x0m0yX51I5QvP7yFBoCAiM7PJP8Df5A9ripQzc6QxeUOpDqhW2e+56aSQugXFA1okx3QY1hC
pfI5SnUItBp2qJWoN0xUfpOkaqwX3Hri3zTM00bxCakr+J38c7XQZiosp/2vonwVkzm3ewDIg3jh
EKhSZYwUfv88mErrbP3pZFUm7ZpR7qIC8LEgHN3ovKVv/S2tveZ7/KhKDQ11kPoP/AYDSdqDkFXw
p7LEAU7nauz+O6jzr2x7JzZv43b57Ef+SFcyp5ynhbf5Us17mRY28e/+OSbXujWz920RKjtX2M/B
TlKgm+LP7fTEAJsYEZVbsX1c6TWyqn4Pqyu4JitkePl57ysa5CtgfdHrTYf+lCOXZ4VJ659XVrk1
Jkinxwuec0ybIEu+5bWHuOlHPlmGf0E+2B+MACWAXpQGRH7EAtFDv6dcOv2XowCUgBNHgwyX2W0B
at2LVOqz6MTFiNmSk02EW9mCMfmndBLrqThv6ZTqPr7+anxs9fp/zh1nQX6o96j5URUDWWRGY4F+
zbNOMf2fn/cKg+zjpq4hOOyRywWUUT69u2pnTHm7p8A7KQr4UJKbz+Am9seaxL4XLGOHXfAUtlrO
ANDdO9MdMouFEiA4EkwmNEtqdAT5eM5b6HbKZcocOKxAa//zQTmZfp4JnhZ6jDAQK12oyfYQdCUs
iud5+JnCfgmfQXpqHk16u/ckHJNTc82LH0sKeDyYhNrZ/wvyy3YoXmCO3ipMgGf2iIk1s9MymoOU
iztom2h2hG4WIdOLmPHxmcW67QvtCBLACGgM42RRiXRFgvzveMdnyNUiIN9+WFgXFD+PFEPMRFMc
TynlKB/wEf/iw1tw65NyqmLeD7znm+eHWsoDeW6Le4Gi0GO8BTSqzKtnwKnZks0uf62ZYKOlS10b
P3/ntiDqO5xkSrllLwSWo85VrgJJm5J8cAXaMy8AFrDICHBoazi/0z1ToypthrE2rgVn88InstPM
7Hl8Tuw1GCQfV1KRFl5qr+ce8mhrrX2TvgzWk/pxKHUhM6eyyLsilGvVdzmeZl57rAeUgJtUJlLO
edWKkDtmPubd7afgCKLmk4HedmOJfpDK1hI1u0KS8LsJHKRSrGHWF0OO/0aLoz0PUvLrBH8Zyp8s
1aOgXSidnXY1vMhcFg4d+hCDpxSGP97pHZszQ++jPip4Fl6KpIWYNhknBlmQy6dG5pLMy71Nya9q
DN6SDiRYvObLLBqcWHaeAVvZcFNx4/tMLgprkTj0QgvOVcfU8ENY80eaQpReb+Zc42OhOA45oHFV
eUFA0jXOMcsm3rjz+eKsnmhMZzKfVM0ghszDYds1+kUdOrzRpEycFOa2P9371/J/wB9whbY9zpSw
UEfuTqHuuVl7zw07bkDR+sbYTPbf9lcoW4oX4N0GlZuA8FfjDk9S8Q8CnOsQg7i0jkHzG5fxsELm
NjDJtQC4cUr1p3h+o8guwZuCNmdpPrpY3zciazzMKU7eg/SaaKZ25m8qvGAHBhHOvaOeN62C1IR5
4OgdqhQ0T1UdaM8O2S7A/hpIbHIE/0bNw3S1TYcL0qX73l0MYDONodzRHnALxUjUODqsHNZ4t9g/
Xml52FC05lrF7IRa9B/smOJTc3NMLEQh0nQve3sjm3HT7cc7T1rvIeOrMlOULJCKLsx83ek5DH0d
m06QB9omGnYCTXvcjVpevaEzH9WSMkMI/I1YP+GOZYBIcxXVSESfgjO7KaRZQn/PjJJ+4Db/6uP0
VHs4tOEsOKVDJF3PuckFeOgZSyyvTDzLV/P4P4AqF9hXavgV5ZwCd3cs/rDtecJydc2zGBH5Xoee
PCU7kP4jnFGxOnNMWIMJewFAE+YNuhls34rXBJf0jpipWEc1ER5R7PqX3oSMMxdd1GMUjF+EP5uj
9C435L7vrMQfUoh14zg+L7AYtUGPFLH48wqonT/sWGb4vtqzOLmAHrhe7i8Z8va4Ql8giu2fk9yM
aaDxsnSIq9aOdwEC4+tjAW7fH5bmwoSoFpa9RKpvzg9jaCkyJiegG6DXKmG/Oyrbw49Eux1IjOiv
xHAP6SCjY70Ki7sdntGy6Yzrb7LefFO0evjTS0LbKd8tskW61rLeGM1GsrDRIQJ0+oSp+dkXqO0t
SE3CT7+ftuwdqIRxAbMMLtqnB/V5CP0rk3FnudWsX0RBVf29OYVdRVoqqX0Gl4UjNRcX5BCjgUSJ
2TucRGIxzA5VZwfZvBqyDsVMxPnrgBQanmRLNogsZ14TJ8VXJ46zh1wA52ruAi/R0Dp8lKm6WayI
EMm5svTPz7I9Wnv2pSUFVXcknIUnk7D13OryFJfwx5d/5qPVSiwLKD90A/g4GVGzxKJz62V+9a8y
+hGPcGirgv3J3GbrrdptDi+2OEBWPy+6E3rSW/9Mj6W+NDTtqnrrwrpsdWzjYIzOwmEvLAGng2dD
rTu8CvsLpnaYK6m+vw5RTWdqBqZhiq7G+cIkamh1698FY/Cxp4H9XjKAzaH4CCiyrPS8yICs6zgy
Auar7TTf8IzCs6EoJWHuXXcfDwmLoHR9qUFpNE3MwUndK5TJXgCWOtvs0+B+UM+9PBu1q2BABOkp
aspfR+NO5Esq6dnTU82grqLDWn4U9TSY73kGQ+xT/G9eIzBYFpSHT6JaSI9uyTBrNq1tp3Zg1Io7
1imtKSve66C2y5JbsHOyGZPuoZzWGejA3MawPUN4ogOFwftk6IlUYT+C/DmpDtDs8QG0hARKTlVj
NlbGjXkyUPBFGU2qiFJfYgHAMncLi1Vra1SFe9sNgSOJIGi6lNnI6R18dUKdkoYTocmZN1lHnJ1G
xuesKmfPCXA8eqG13oovd3VyoYNiRGl/6HO9Fpb/i0X34q60kISDvchight4GJiUufeE6O89nWvp
wkCEdFVzOjCJCQtd21xYDQe8Mu13TAYQRRf99LfPLSxE35ggjJeCJhoMYtFpwR8M4paQWcLFMHCL
QIao2BD1o1xwFQWMKa+43aE1nAY9XsBbcgoxubVvNnZGA0YoxQ93pNnD2cax1J1zu9azoftGUxNH
4UnT92YKRJ9Dirk8VeUi5lhsHph01QrB2xwJ+aJA0PnUUf2WCjp7z1s7U+CagC+7sUgx3OqVUg3W
nUqQQ7iWuzEEHZkwB/jxUxcI9eap4PnmjLXDOXZKdQ4nrlfo6aFcwMo2V5FtYVaZqiMOo6M73Pje
0ymWuinQzvkJOYFqlkmxVyRZEz27Zo1tuKcsm9bZ+sGHqewOpGLUMZxV6o5i9pKPArA8uSRDtxbx
jLa4jy1MBLG/Kyd/bQ1yfuhvVR2Wxw/qPYxPB7Vcd3OiUhIhUxkxMVkIPDi6heoTDO67VeI8DKD7
VqMuNVOr83oMonuMv417krD1RiHqPzH9yCYK+C9SCawyLysM2hF93/8h3r4y+P6nFK3WO212fxeX
UjJgMUCC7V4nlcnsfLGNtwf4oqPXKrlQBHJYHTWmQisdaWF8Ov310XEsiTgTrNJcVRNt5zo2MANH
fafvtgn6EB8rNne+KaCLIoMr71cgbp2UOZawrEPAmcOwqv4NTalUsGkCM7aeD/Z3ctUY5G1ZjaDC
VIulMQrJf8GKLJGLDeacBvZwO6t/hODmVS7wo/wgosPBrXndMVALueWsxjVxUhq5DjzMnSSEgEAX
wnyk3fhSlL+eXZub+ZW7gW5kpVfx+2o8qTcDCJnMuRaMu5eJk5BEmSRwc7mw4zYFFEso4TFVVXwT
6QNvMIk3aimuBgWdEc9F+UrrHkqyJ0hiJ5UaJQ4HWrzzGOKWGMp6vkmJ13hHsrnGVz0NqyzJPrzy
AtOmBaHkGC+b72jVPSLDhx0zsCMzMlI8KxIct/CjgeSl+Z/coJJGQyQdVlb0BA4sa6XSDIBvPj7V
1lgnZ/U8xV83nhyPq4yo9CliSYaxi4fk8u2xEC/VURoBnZpNQb8jPHRTZvHXywGAeO5Z0m4aPPSu
0t1QQYGiTmRWie0/XOjKOtNZLKjD9pVH8PogrGJOVnjxAHlbIzkaf4R2wVckHsKfHmVZeRHORv/b
j2tf76EXxY1pYyxUI7+PiGsvfF1FrryA7GpUDzGdDbaKqD/7rzKoR8IqKL9geJwkFmUwO/K3DBo+
XDcwBCpkO3Wjsn7RZafOjVeWy5xgcUJXmTx4dFLDMhdaHhsn2uUDiatWfm596jo01GqqV1SSrJ9f
Ys0zyo33OaLnBuG+sYzygYo3WknHKVg+pv9Cl+3KjIOpDR0m12j4lTB/K6wvmwDfgnQoSGnNL4ga
i0VMob0FdwK/L4Vf0geoq0Zu+nnnoVnPevXxpgQQmYNJSM5WHCgsvrmTmHjBWBZhlQ0hyc8ALeqb
M7RZlvdpEJM6S2sn/E7FjX4jnDKlC69lsAbP35aP42ZxLoR2FZlHPmHNCpQg5NBEBwyMW0Kzbe7J
g4VShxoWbW0e9ZNVHf8Dn8s/kAziF1FByi00SayFqB3zoiyXfTgFoBgZonx+c6lOAsztmhTup9SO
CUYmTEE69fBy16fBVJG3//S090jqYQBQw3W+kdbpQCjKIwfqzZjQ0Il+DVjFeEn54FCZRCwIcpwS
XlfrgJylPTzSZ3rTenPoxxHSs+j6AOsPDrmo0FIMB8I+HVMsFXBcchPPhRpbVv3jQf7OfLgeVKkk
oQzfERzYrIcoeY1Hkn0H9qnIdwvH95ERV0Q81Wk16HA14IhlbUb/o3ZuPNrrxfHIyvDXDJTdbc9E
eZCGQiTxgvnIuBSNcV8yUfeX1Aum1UUlSFvGWPk/EPIG5K8ix28PQpFeDr/lkrhie3hv7njv+SEL
beBDckcKLnbedP468TjAWbkuBR2x3bpyo7OCVABLuVgtqkAD/JxjkH/hK0qMDOKzSZq8V4M39AFk
vaeLjCQuZezTXUiaxU1jquAaSAtOp6AmuvMYOGTyFr+l7a/ylWz3aE/cY0oAVpo0sLSk0cszaMwo
9kmG2YGiml7L2Ew8Yoj6icK5fKTh5ZzK0YqGjqlYjIcngCOwFFd+v/wE0VMul4LvBxDJYoacz9y1
ETuSOA8Rt6YQQPGj9XxtlLot2kSNmGCoLXNFySagVFA8HLy+VvFm/rOfnTGkBKFE3Z8SKo11HsXD
OUqLba/PxU3VYT+QZ3aVgq3hAxtLW6cAiOiBAm9B8vEiLFAACPowfpaAY87QGB1RNCgMyKn9RlUU
1C6bnUnVxVkNqCbdViIYrgQyykQY9krDkYxDZ7+z1aHBVjd7UljgcDcpvXWiitDo3KZUk3InYz1G
mjESCyyywUqVZVVSkQLlAiVBSYIBdBpkHML2hJJd2aEJPaC9RkgEu7X18AsHeIfme6iu3q3O3psQ
62TKivbqM2Ooihl14MSkCnO6y90Dbenv7xnFov+pD+KrGJvJ81RFJoUzxXxjNYDfkclpHndeHYK9
uCCtEZnTcKrYbHAVD5zS/eNAe1BA8sdgkC7OHsfg1d7i79WR0QgBTk9Dc0ZOkWVhpt4UUcEIQo2Z
6r9gI+2VNEsRWyU9G0lqHgJXJrblPO7dJ76u5FXdsvdTsLTewax+yWhsJO3CMgVcotFT8YcLDZbu
gw9XJl5KXEQJ1dFmOHIOZJmvlXNoLkJwMM6A8Mbbqk04hT1mj36X68uQxWFtrO4bcTVvoodettII
y3/3kbrhWySaWfw8lzH4bS4/dsb+hiI94qV2ZW6owidkufimlGuJHntQofHHdGBJ3N1bsY9oqCfj
xokKwXQ1lVDjsBqw0yhmN2bDyqywVWdUiSaMCQ676xVw5mnXk3osr64ReISMG6IkGCazteTPRevq
DI2mGlmx70ssB3fH6qBOAzHJNuyOD4qknBBdKHOxuLxUsoZkE+JMi2pQ47gPxqsGj1vTW+x27YK2
pCnXy/cAtD2WntGMjzctUBQbDnvH003pyxvFSuxM/0F2xheZTJMd/8eYfzk7xs2vryyOq/a+LheT
jtH+5lTqkLygPaxMjz0NvlloM1crZIkNAtdiYup2mh/CgywjZm3+JkXsI7UnBDJTzktNnAKFjMyK
EmivQmqTlSp+9diyGZwmbe44pf/en58ff01Xc8+SWnaigw6FFJxC/M2XVzSx7Ppw3GfmvJJwdOAi
92ebem9A0OrbTym0k6WJiDPz08V9PiripLQT4CvF5S781QGOE57+5dbwL6VioXBIGZJinYAIp0gY
+F13h4fxmE8QEuUcpYyERLX3+tbD9RfC3qEgV0xdHMDAIQ5Eaf3udTwxl+8JkLqGsIqFBt2TX5Tj
/5l8/koB82cv1idWpNSlywRg6U7PZlx5994iC2qcIITeWVEsjul/Bjek64QCMO80NCI71dmywuFj
gIWPzrz9V8j0ZJN5SuExEYk0TItjM9zNY4EZqSUSYl+gNawvE2ZjQvcEPb2DMViS0GgfYAXNMftr
tmKzSMr9+eTR256SiZcgRVhRNwEN+UlateG9Wlnh1bh3PlIvYE8HFw2SCcwW4JlsJ0vg4iCqdvP3
xc4qvpmR80rDOJ/NtDaz4W1LsLC8PP0dVmVbkoz/IFxNSikbGpXBmj5HKnLXqMvjYOhYSTQcW0TU
j1K+2t87SzjsukuAvljc3/bZ04x4pr9kU0f/GMglwzaVXlnJ6TnSxFPnxwNyd6qLOoZCqZ4F0MEP
yRy329uYKRyj/9+lZNqP6PzRZ9dAaSGRE2575GvvrAyAc3fsbQIZ7kxhIcwYa4wHNMWQ2w0aMovq
Ecpjz4Qxx6tNQ/MXsnvNLAel8B5BduPZRbfA4VoyF1i1z8Ylv6vLUCr/NkfTLv7IsZBXMU2bg7JR
bvS+xHeO+eVTXlroUQ6WRenLj3IJtBP69IfJP/o8W1HAGjJdFrSvP0P00svTlGDDqSNFrxAIh855
hTgtvrgs88/X+y9yME95c1Pw7NC5VOtLqbRcxSEpUDU5PQ654HtQEBfVV69cMzvZ0Y/BZMnlWUHG
YgHGB1Ie1G9NNdonv777uVXa4iLQNFhRZTFOFnUpNIoypgUNqd0N8ousRQdOLYT8cIGgMCJifxh5
77mRYMlFtsWjtvIcfdgsVl3/u872DKAHfJD7B2svkGu8qGlcKIU/KypEydmmCsTG6K9JGJh7YWim
4Gn/xe1PQ3UpfhMd+VF7mGzvUwfstzIx9qDj+B5QGdAX+9GTInP9NQ9WwUx5IO8YTOXCIiPVs2zT
1xlei/q72faAQTIfuSnrnt0zZBml9FPW1QIEpl9sCZMqJs4MkAMhuI3wKuZJrl+Bp9PaRy73bSJP
J0Tg4b42CKr8Z1Y7d/dcz7oD3n657VSypLzgz8vxvplLijUuZS/DJKk6Zb5jEKOfHmFxPx29Nf3f
eC6YbHzI2/FEug2LHGo9ogcfrYTvNKnGoc8CH3fL73XbRDTLNimwNprzT3191BLlZa91z7T+rWmY
mB3El6lNi2o6hWfK9ZNjkvEn4QrHZYAzayk7hyrZVMl0n4OvXfrgU1ZzrdpLJwohKhTu7FEqsjYq
F018v9dZdDRPfHkm22+w4peuUPRdvSvbOAMsBZuZjDpF5RbSCBfe2JjjZXJH0BYWTRZMNCTTrFno
act3miDhTng3sheZfCiHvBZZ12M/qfp/KZsJHBSSEpIjpnB4fDoF1EJBesMAnoVwcirVDXKyXrd6
B2URG8vtEE/vZhnAk0cUb4lfkjz6AoPEe6uKSSuZB8Ogqh3uoPldV+o8tGbi+Nu/HDGzQdzvFw7H
EQ1Hy9atXDjl0UqwHh7LmDfHIJXaLRz/6af6LqPeQkz/bQl1vIJXuK6hy+2K0w6h5JBZkyKKJn7i
FzBq+WL++fn/QRdvwF48P/Yxeg0VarCjkIhTY3EXeaJdOhPFaRtmSuveA5x7EC1veeHO/Hg63KDK
OBMSmJt+/yWhx1ZJ7yAqO9zkl8vYnjfgVGTwAh87VBG1KCnbN/lpxv51JDfZGozQMOBXLwEyORRZ
62M46K8cLsz01hhkLx0oDierYdyh/UlgKExsCX/zvedf5V1xomJ5xYq/D+yqeIe7ohplRFrWNk1w
GrLjY6i8JkUb/OFYTTaZBK/gUVtMlr20gd273HUWAgxdwU9NRjfHdi2BVg1JJdr7Ee9w7k1PRzUk
4QElu3GR3k8NaDO6QIyQGSsYGhG0Qrp9fXQZDdRuhITxsERs0cgQUAgR1JBFPGcarE+kTUXx5qEp
qLZMRJG6cGB2mZp3A7bnjKFECUNaK/iuhtmzgN3R/wbKi2fw8Fzr5uLRnxQdvB+UTTtgL/szoD/w
NhrYuJsD0oirArrrsPRQxw2cGqAmrXCa1R2CT4XN0AHFSc1sxSrWa5U9h7+XvEbkc151gJA2pKpd
J8rFWpPCxoZNP1W6n5fXtc+3S5nwxtQpF4xV0N8x/9x3lm9w/X/B/qZKSY9990BBiNhmJPA+nja6
dv8OwUz5hR6vV64fyoQbRFR6laaM0Pfm5S7xhkpU4D0A4R1x9kv8hMJbqP+FDYW4rlcKBWGk+eGA
21FLt1uGciC4wpDP0wzAjBtUMnxbgUG53eOKULQejQJxjtPF6EE/OiukL0+BhfZt2PzLQ1ld4CC1
EqcQgzyddO3+x9Ae+VdW32ztBe22jWA6Io8DL5mnoCtzypKTjxYGz19XOy3keybRyId8/8ScHr1z
8rcAFKQHkSv5ssRUA2e6VcS5MyWOK1MVpN43+boDfZ+hqR3BK+tRBh2ESX7qkaMExdsMCQOk9yfe
wt9Z9x3f7UfmWZ/P+bkd8bsmj0cPz9gmcTmHV4PgQEDTh250z4MUVMVBh3IGl58+E431p4xLNOVU
iv5cTJdy5ThtMte38o2OcB7v19GHzMsMCyeWFky+QOsHQN19u+eA6cxOB05SeQJG4o8b4S+eEDmy
FX+e74zx+RYIo9OmKKG6tl/uGA/PrisfujagIJXK1q4rWBQFwfm3utEzWtGGEYrQU6SqHtTMyyDX
sl4YikjoMwwkCNL9Szq+VxgubdI/LpTn/9tUfLCtj3UQCrSHWUBwG+3ba7lBgtmoCCkk9sS+W5KT
Jy5tU2j7cZ0yIH4CIhMJdPXxGsY/ToHOYYRqHS23q8F2jlXAAycRXKz5t0O6b58HYXPHKYrV8j/7
Kn/OKOfYREhvbF/P7OzUHyi7VZ3cT4gk6qdl4JgKjKaHmcTaKRIJdJNPd+NlKVUU/G7VNwNcvRL2
FSR6I4dB6MTEwe578RrLrTN+Vljd7AZP4tHPNILvc+KzRtv99h6XJi5bXIpqFEwpDXYfVY9JxiE1
QTPIj9L0VQYkQXv+SCUR5hQX/Wd8QODdXicgQFi6s+QRG0XOj2Ebb80ZuJhBgQMJxatwZwLBx5SW
iErHHXbNrAaQbsqV29eXZNgI8NPmpdSBG+ZOC1a6CM36BIHHoaiZv6fGokoX3x97NM5StT/AxUkW
C9emxgZU4cbDF1Vs6oGOJmHFFMY1maPYso+LcM8RF/rfH12IcM29zV/SL4lvZJeIuekgfQvdEiOc
81gI+8XS7e34svMaeoGrruDARJGqw39mlWCYmVwEPkyRmaTlQ6SujK9wECC2K12ezV9N2Qto6mAD
N4jf8NyZVkIFq9bcg0mQp1sGM3mlq9wrIi8QKoAdTqZp74y6ZWvbGAbIdmT/CDHt9W1dEvQn6yhu
BhUmog7k0nNWmavzyjtzCxHUfkkBPB0dFPfN56WqiCGG/sQHxhJZEHWbBkvv2ltLHJhAXePSen7t
mZv7inDB/eRBlxZ7SCv3MPUHj2OrygbRVnxLUJ/nFWcTak74j1TEciXayFKTlGyKl/fyDu/VxqqJ
f6cCGyS75CpqHBLAXjRCq3f1pCwvjrQh7x3GsC43XYn1xEeMPblt1CN8P4E3aI2ZLNypK3WFnYy3
AEgOByRtYys3g9aV+mUvg4vidUr2gBdF6hjPTNfLmPWQJCw8c11AuUPdhLPXufsXjamhjFqvqe68
hmJ7ftGue1kHVBio37b9iN9A6y9dIDaSPZubaG7zNHrXNWjcUJRZnALR7hg9mk1SIo3PRnwzwd2w
vy18nSS1elMy32ARJI6o3PG8C/5iJYxvjU9FYKVeMDTjvLubD1PtS5o1g+LmhUR4x3iOqY5fcG36
MYx1NX7Cb/hPB6LoOXZE2fUlzH6A1eDucICOK9cXlce3dRmoln2AkdWDOy6PfL8rdN1PbLG08Jlt
/enVkecLS8zz4+VohIKR5MuerWfxkuMsetJZH1O5XD53YJxzm9R09Uvz/MlnO+9EgJMVy6sBMiGf
xbX3W8mShf4iPNVTEk0DfMoQBczplVTkErjDmsVLWR4G0FmTkFXJGh0V1SsplOZ7eVaOfTifV4tY
3vdYthU853qqZuBc56pZGYfZTufYG7vB0uaiMU1KYJ9uQxn7/L+y+cfeptDMOlROg8Alm8HYrTPl
DG5EYX5M5c9+hTSPb8+B+mCHIjTQd51z2r1KX7VjjY75tING2ancRxVYpZmmkhpSKxZLTnPm+Ej3
sw8bQnzo99x7OXyq5Y1UDrvTB11ZRQXkGfDQFbSPqqPqX1QvCZh4gGxNFDj2l+AB+77XNvtYmsHj
nqMzPzp8urt3NqP1sX6lhmQNSM8elNqODSh9Js3lWPbePy9XXhorS10eI+IIYNa2yQIgwWy81z0/
en9JHWn+P0RxZdsbtkalGY3sIpc1AiBwyFtbtNXacdg1kmgqlwzaICq/Yuf6+PP+DFh/mKuWbp3t
ztwGysNtOgUGowMRyIVIJPo0DOH2x2AjqnlGBPtLhxpabmjzhA5Jv5ugL8OwNyN/stP5Lmi/4mvw
ywktActtHarEV/B9bi/sjPi+J/e5i3VClnAsBEX2NUAqZfyZVPa3fY2lNLGRaToEEUO1or6JO3y4
CGwcY7uWkfFReRCqW+bBcYBCkmk2XBNDUIRXu3qQfd7Vxb5O3S8FoZTOx7jlbOLZQFBkj/hjomXC
6pXEbfuj0XNjE8npOXesQP08TlVUyNGa2uovHwblkQZTWBhbt9y4rb7QWPYJxM8KifkZmE+kMRyv
+Kp/oaNpw6zY54yQoXrpMW1gAB/mJthbO31hyrOcKLxMBX15mxePUBFZ19DQMPk9V06X90L5877e
BZcGX77nfX9XfFSmvHrS37sZ1DtrJ6UE/y3nRjqc73wWxYhHCz2wOBMPOFmklbIKn7VP0XoTHe6t
jUneoiHD9VHveHTvOCVtGy1oD7IQFv7QtrXMjOBFq05ghsRKXBBjTlHb9zCTuL7VjMjHgwfTPZty
1FvsL8xdOcueqMo8bA+uYm+26I/J1UFDu7TxBKDPAw507tcIEI4femqHSekedHyYSsBRZ8B/6G2l
sPMQrAmc2PvBqzKBcIcncyKtVnc4tq4mcW7jptYoo4lR1GKW0e/ljWVbNKEDr6QRcN70UJN95Qzc
y0O8CB+QCiYLkEFFjGfE3zk9oXRnc4gm8sowruAP6PmQPPvyPVckyqpC6hyWi3GtfBde0fgCiRjr
8NfVfZ8j0Ihb2HlBnlFVrVA1Lwk0DFrVJeULjoSpnYKDdH0kL+c9vfi7Dy7chlaEBFA3rN6s5gS+
14Y63GJmrJ6NyjkCsXnOwsFnKxte3F7q0s6QRVAvK5hAC8ZvlwLGBRn/c0D7R9sCYNZL01pu+EC1
qxOuHopxaIFoxTtSp0szTQdVlnEpxKQRXZDPatyHK+nmPiOXz78vJbSxpWg6McU+3zWk/1ZwkBSu
ESb1azAeIagEQ9bjhERHxZ6c9Zzu5qCLl4eRkP6q3b4QgD80vydxUuzUrimd6ZiX3+7Tm9nX9fGx
BSMPO8Ov52VWaCSgTp9e9/Sc1BnNPc+fNil53t+lTsrrz8scyN2N6rJm4nc+z1RYQf1Al1QnGwau
NLwXzuXZE6tuxFp6e+q1ujGKr4XxE0kAaQf0u8QgnPTJyof0zh/tOaEwiEnz8WgF/TYGyIuTYl4x
voF+l0wW9qnUT3YtlKLCgZOcb6l8e0hmsnfXKHLMNxfVxExg1QNa5Alx8FGBotrxDp5tGpQS0mgk
RIO7sy3p1p6e/+/K7i6oOmTWgIUkPERXXabX3Oz8gGYO3yUZ03t5q1enoAnuG1SHhk7TTmGFTFor
c2n1GbHpT3LU1/FOb8n5BAisVxPpVgqqdyOpz4VAmlGoN9EyUpFv7bhrerdWte7FTDmacRi6rmtX
TYN2qqpesmhtc/6YYJXwLv86r2nX8kjjTSFgQhDZUtbXV75QyUL8NamRZy5ehEz0W6SAalyuI9PI
YlcrzKJFjlLomigp6n48vCxmTBL7vMBPux9x91Igxyns6VdySXbeUpfTQDad3w22pLBtEYypnekN
fIzg5mfYEWupvrwVMJiq1B3PvLgNUQSohYxs5SH0aWwvQrbTk4jc0f6gXRFBMbYVM4nPs8dKhenw
Y+YSRNYCRdpAXlT4wwcZ8DV9TUObVld5nQVtKzv3JgACfr/LkuFOJ8TP0GJh8uump9NwR5WZEdWn
OTgVf3pwR8vFO0Y/+3fnjYUOW1fM9MH4Yz3XWFYl/mGnOW5omL5ph15UtwWCXhyXiOkvByF4c3mE
H6VDFeIs0LiLPJPTFrKOeZOwhcZKr6KOHRtGCisqtopuQ6FtSfC+LNv1MTH5q1D3OZSxv/KdRugu
2HL8KYspGtxYV/0HalT0UyP8/SZrM8Ef8bUJWcqDpmvhCvhGBgE4sBX0d6dfHh37Pb2spDkTJ46b
2zxWSWXw5bOt+MOgA5R+HHj0SqI4xWPlSTICWa1r3/AxCfFO7U1v3/GlbKbqxNVOAbkRMMVKN9t5
K68T6L0aUf1e7w4jr/DyhUSYPe/WmryoxHhg7zOZLNMwFFSTZOx4Dm90Fl3uitOlRf9JvFrkC7E6
izd7I+cQh6Cg2DTZu1ODl9+tORx9wWPXelTbHC9sZQD9qC3jbxkKmuGU6AAnSBqmylN2v02TX9JY
wsasbCaqgW/rVOvjasFOPrcHToibTxO/OnPoLb/T+ZmD/opBviurmi2xZMj6l6fp7L8utfnG1BPs
X7sJodaVHQym92WTp59FuZzgywJ7NDdIdwYtxgEvX9iypWPjakuGcFQ23LdmB+hC3CwBiF6EuhTX
eavGAMirWjRsNqLta9oi0h9TBQx+e8UWLTIokgW3mOiSwKOFkJfGqgrnviXsZv2wNJtkg2Wh27Lo
T0GpS+yvZqXIR2qPbLS7dqVBLZ1iAd2o4MJBIRLXoKHjQvclgnmZ2MFKJE+6bX3W9Q3sUlJJZmz0
kzYsAnUQosn6Pn1Eufe4l3uBITxmdHWGXrw6GAB9B41Af6qHEw6LSQnXEP5XSFQ/oyg9/vt6GAWq
ROBCJ9DVT2stpBPlY/b3Cpu0j0vYJQZdChzkS/blpX0LhgD4b0IO+mJ5Zaktdr4TDgNVJodYC1fh
f98r1ULMSTnmb/8SFY8my0WW79AdDnK6aFN64DQ1p5U8URRJi2G0hdmflq4U+Eyj9p5zErJLlj3j
7pNOxn5MqH3FjasUVKQdRYQ4D9OZt6TU9MIkPHt6lyDcqrCjX4ZqepsArIVcaN6AfWo75Bm+Lp2L
NCU+TExbj4hDXijtMoKxSuX5MtP9tfTLCJT+qDWofP7nvBaUKo+tUdXQILUO2+i88524TCtwxk2w
nOWRJlOU0QMNSRywYh8gNQcj5OBQJV/PEpeFlQ5NlnHd0pwOHaCW2OwOTLcUa/9qwipkK0QS0A7L
nm11/pQNXpbP4+c1PYVMbp0T4x5EshS21p/0kMc6UtMwC5UG5Z+7n9g7EyGVVANtOMkZN+NRhPg7
eCYFNEMiG1iAWZOdSZqIkyvcigR3uyr4RmVCDyAnXpP4WT/lTq4OyyQZDFieBm++yGqTZmdF2QPo
HimBWURlps4uL67Dl+Z8Tw1IhpHmXPayewaXpYnA0BHFkRxpKSi9tYzLjrWUYKtrulX2NXmphonk
bnjNK9qmNzxPJ2uguZu6bLCGhr5m59cDlU9fRA6y4idn3pCDbI+OCCNGbzvHFt2RJZfna4m5oCj6
BP/nnZA9Wrbt1y6JOsdfhbu4AhbU9TrxNE1KS9Sd6XkUlAUzqeGnwihal37NAbTNMQ3vitzPdH3c
3Ng18njHr71tbU5xBOZLYpGzYz1DFStz2Y+a6y5SzHyBdoz0gHBfXLSQhcDvawSKSfWtxmC9G0tt
cn+noP6kI3HyvjVnTCXpSUiO0tg8IV+ZWnMMgUI17XSKD+KjOCsRJNfhHygpx+VUIN9vQvidCii6
y9pYxoXEVM/kY8kf59hUt0SKKKR5tmTLQj7TYEzIs6gCdshaCIbxICE94zZXsiUWzn+Kn6CTK2K3
zKk/ewCcyDQuaZC95G1uzaVToyJuEs8gS7InWr2tIpM5j1M92YFs7pDCTq4hNEnsq1UrI0WBhD5K
RgqOPtiEEt4SJK+5i8qXAAQNkVPAy8cW8nuv3OGzIb07qLVZyUL4o873a4NI4y6qnkb09ZF0N3u6
VTZtrWs74zWB1YrbIoQr2GLVvLr64ye/YYLBLrx3qYxnR15mYFhnFvlWrD4wBfxuaDvd86JFPq03
yUFuCWdvlagkhKjVRalG01f1Apt4RD/jo4UHluQy4WobGK+QiyPZfRdBSyz6c7Fyvdpc6YVNMBoc
EMAKj6aKh9Nod5XxzfmKzq9NZ62R4fMF3ePMlyXD0mEpRTtPOePK/UMkwX7j8GZ1398Qw38zJrV7
XekOtQovQNVx96akVnJ+3slrrA6FdWpAiyQzCm7DbglyRLV6zZgY9NlXvp+s80XhWIZNnrm4CP1v
YHG7gCe4ZyGd/kqCe8Hkvg2HosHDHCgTGit0kwitPFfYxOJY43M7WOAqz6qPPNefAFhuh9s4aVdx
cunXxwtw3c8nANtRUEbwJMbUuorI8HGTG937ZMgIK0uee1DKDKWNHp+fmyuerZyevw8BaQKv0Qff
JbDpVDPOs8CmS8hG+bj/DSWrj4QWtBtnQ68FuNM2pZnfG6JAaEAJne+w7jioY2nVhfeafVgW8sy0
Tj6VZ34PiEJvvQnGNmBgfZ7cxzGrlKnumDmoiCNRxMjPC07Kp7Y3Lyym7rSvh86Y32PNWPI9X2X+
3d8QQRloBbEG9vda4EYg2Qqbyt8infIi+Gly7pJVv07hv9vh1O2eqTNSoeYm0Iofe3QxgWdWy7Of
t6idGCpUQ+Z0dN4IE+vX5w/lCN8qAIqSOcnFwOWTYtEjtx7DFt2qoOZGWt5Ins22FLFNDY+GQWQ0
Zw6oa270fQju3TWeTaG98x1S+y/ZwuU8G3+F6eutguE5fKQYyFomUPj/Ed6sZSXPGt+oydsfAIiC
T31Wy6WgYzXDXgDHRHNmdPJEhgAxtNTVMV1cKAX45DzVOPZz+n7vBx4GnSLfgm93IQAy5vZhJlRM
OdohNmeVK/05dLCqUrBac3tZKE7T6umMlGCPt1GCFF2Iv7M10pfD/jKkQ630AmC2kaLZr08DRvxR
vx4C21w6htMA7p66jiKdaj7c30DT+oc301ddbbBHqNGnKdB+GYPLL6IJPqJ9XMV6xYrelBCtbrfM
8fCv2GlW0+Njkq/CFn0qg2M/p2xLY+XqWj1Pe83EVlBuQTAvZdHhqi13iyqa9+s6Ra4AEN4qoi1K
zC0wu1kwf93iSjQ7BtCZIu7MxFqfbUjFUhbJEdA5TZi9dI8CgqbezHhttlKagU9SAD7KibcPlr6l
es1Kw4siH3Dpdqx5XbD5Ah/miAmdAHY5BDNOXNbP3O7SfzxbC5+QgcnZ7U2LjrEZ+PVhHzpkmjev
lRjVDCthhoQ+Y4rm4OaNS1YdzIjVyBvC21IPfq5KofC4+cWXilZnWFW8dpltIPKDHXEBduD8P/9k
sVvXD8YRmU5PZq4wwGpEO6h8VF7L+cVjNDxefTJUlm9mzQE8Z4pyLdxdkhS61Wmrdz5yIIrgctY1
vnMmmnSIYofEkL43tcQn5Q6HnrcgXLrK52SeAGlGS1c1hQD4UvGYWpDbZ07Gj7xNXKWZwNQRktSn
MqVfzA2+7dFy1xGcoZva4grP0vOtuA/YfCbtdrdC5MIwBoVg1c6T92stHB4YzqtvkEz3OfNaKJIM
VxVk8WTQvoDbxqOMKnLrwZiX58C5CyQEFCKpARdXgsM0YPNnsWTn+u38FYgh8vrkGbOMmxbnZqF5
0aR6eRN2HIjq9AT91Ztt21CJkJEtthKDyVonC53ds9fCuXL74jAHdhBr54oTVa9zAas2uLpyco55
4OZza4snNs6XDq+41ptcWUrsTJtKSYrEeqOMuacuShdf/OtZWv1moTEqKzv82ZKGYeLSAdtjTKnb
pXPKHNuXwLkk/0ppfShhcSjeQMSHMKzNpqIO49GL4zqx2WiROQwyN8EuVecoj6TMll75JmN0cDNX
B6GmyKubjLPd40MUUocdXo/w81oTKzIZ7dbC45NZfBZS+gBr/2qLxfSXtt1BTIY0/gatIXaCgxEm
4RU4yb51EDPfGdUMRB5J8HmqC3inKUcrQrlRTfxygFKn9P4+71+yJbv/PHP4TX307c7YR7BrgXeW
cUo63/pbhLoFfCjrZOZY7ii8waJdqnNQJgnVpL+qbiwCUG4YIRyfGRgIBU1CgXGejwrlsJt8BMpS
nfGmCEZZDjMd0ZFqZi8WLGZwHPH3JDD6oyUg39I0WXfLXLkWuXhaRCr6EDwITixDyuW4D8mv9Uw8
U2NL31UpLrKCGvtD8zc/Tmj37lKMpMxLI6k7NGuwTPLtmNJSBXBoQJ5m81MOuM+siK6D1DivsxFT
pA8Wc9fQwwYqdkH7j5Cr4GzTb5CtUaifd3crp6jDvYR7L4MWnDA3FZKWjTPX1sQZp5MmzSv/NS0C
eE7jjom9qjbBu2+qpsNv1YtMwBVsppwZHv7sSaqADLHLvprmbW4SB2fTVrlG1yYGyFbnaaQS+Nap
4AFpGdg3bLm1DDpR794kEI8pV//xXFpUo6DtasWHHEr4XnaI5gHEOZ6u6GIrD0nqpo5euyEBvyQQ
GEbC8yLOc6T6LzatRdPQQaPhBcM+TMAWfAEfZIXRkwi9xkI1AAC3VWP/2vuYBmjjyinycz3B2YG1
dT6I27CTnNOj5mxVRT8X+1ndjcKHGV18juTn+0DO0BkwNsp69pDV7AEXgnNGhKAWkwreSriwp3sG
YS0OT9AZxMuG9YshF8A3csr/7NCG0CCVs5dK4JTQloIoLo0yX0frAKEK6UvsrAid6R5hOWr73jCe
Lbpa52YjP9Ie3/ApXO6Ct4ndBaRVc6B5BT3b88MaWvbRbtfM3ZuYU/dUckbk7czKEx1TBbANYbj/
rhedutCikDiMJLr0pGIkdjqFJRzz8THStWe5P0l9VrmTE/02+t2QQ9+D7IrUhoiFUkn3nPRnyq97
AuPX+mZbLQl9u0ebaaqtEsPfJvnhNlwXjUUFLPvARwnM5rqEUeH8DjF0mkq9IQXjPEYxAYpicXIE
7f/GTfa2251/8B+hvoE5T6fV/bcw5fX3TaAS+TLNo375meRvO41nfr/iV7h19nxptFsiZwhGLsIq
23C6lHf4bpuqXnj1+66JMF93K54XBkg3lX3iC9HOiffuD54nfA9aPFOzmqozmVI7btru3yU3Mxld
144CiBi57g1U9EQYH0VoMfYMnOf30pSVrdqSi53ruV1iTw2G5iHOicKGqjb/ld+A836MgQtPI+0N
/3RJ8cYVJCR+iuBSxcYwJLa73pKJMZaHOZEya+zwiK7T45RvN9Rxj8JTlYITbju9zBeJ7xzfjUwW
zijkAYwdYFf7AftbE1/u2/KTivkt7Nr7M4+R19TneUhDIjq+gni1SL+rwVrVRReN3kKPPtkZRiAu
EwHWDcAGD2h3RJ1ZOBFXj3ZWnu+5e8/Y/oCLBidZ3o8OUJYJZAwIu5+BKEZV6UYHxKRK6wsyNJkv
xpMolDUnuJNLdDX9E4zpbtfdQWSY7Wv/3OkmZ6LSRQG9lsFGJf53sAORA2BGS+YTK50A/GVPTolC
Ft0xvECdQ5C5u8Ct1ZFbSXKr5JT2ErV5nFoHuu1ITZcnK+3XoNzfwXqqMijyyJiEaRx/SSj3nPr8
BzlHul6YgBFK9Kl75hFA8189BhSnHa0Ajq+JqzDnM/aK5ZeZV2YVENtTfc4tCJwNoYi6/R5r8D+Q
XWE7AVnmRJKkJraDqnK6FLK/DoEf1avvtdiK4ttFM4fkPrhVInadkfw25p1iNsP6HVkT+sFfzTYk
E4BE19mF0J76kz4QghI9eCZqzbmRML20c51TCKOmfwa+/rHXfIa3nINw1+rQceBPPccl2qpxvZH2
83QSR2U/a9WIMQfLhenQn9Z9lMRSGBaHyKwB1an4JkZOdcRKDXqORBMLx0oyhlbeu1fY35yaL9JD
Aa+bp4pPXikeJMkSTgOA1sO7ctsmF6YoQEuRmHN4rCZfSjTxurQeFAQuZb6WoHUwOm9aokN45Nx9
UULFoOQXnAxfCY+ocLxXGjBLR3UC4FveGOAVpqNzPzydmLQExiTq3yrMIwNhijk5r3PlrwnmEHAA
03wXM0UDNQvgWeK10tJaVgto2DyPp8aonqQ+5cI+9hWecAq6348SZj7RfaJwpSdZf0wiP/3BVKLG
d3mTY7CX1vDPcXYMtzaezdm7R4E69TpTX+bmSHuLFqBtrM/IkEmzNWGWCQgzEnXZSBsai+Vk0FLN
khm9h1FmPBaBtWlAipi+0quhCF/ezOKi36u1ld3/517Jrxmis8aSL364dr13Vub91JE06DK9v/o2
mlGlzPJcgkc9Mw6qBsnoH5mla3zqrcFnv+APj2+1wq+6R/8qZkkb1sGGRNBs9oEWLrwQKJsZ3ukP
C6UOFTcp0cQewScWLfqQYaRWyBP5jxVzpAK98oi1mDUu1CuT076KDWTopt8oKST7ZSJZjLtajCdg
nUoDjc5wmGaVf9w0dyYjskMLD+JNGSdi+dF37y6LSQVi0OwRlZO3wOseB6MQpHIYmfm/gNYxT7Ba
+HuP1hwAaKff7Nx7fRPisleSSQTtm9uigLkrwMADy4HIYE7NcHIvdE/g9Kz+5L73fE97KjL38gXd
TaGkA8Ri3cde7W+SgSRMDu82khyij5NdLIyk+4+fzDSwQzX9X7XUmvqe4k9WSwswJFWypFKA7uw/
/5ocNVwCRkWPWMvT4uIZECNjPojD1MGcqFDBx3yA1nkok6qp+QHPkaNdh3q9MpxedqmOpmhP/ltt
P6R0bsXcYjA24HatmPJW5qd9klziu2u72kS8EZ0V2m/byeQNNueDZ8GG8OpBxSCdbHlijUjlXzWP
wGpnZ1sqZZoAMMOqznMLmAXvGG2WxNEQC85nwj27qGcrE4Y1wz3z/fyIENNqC5qGmz4OM3w9CvfG
xlHMT+tAAnm8M1yLMi3zAzhyA1eURZBBawCxdxsp5h4knKzeJpQXcfSmrUOm4XQIoDfdy6I2PzXG
W1LiafoJSFc9tKivodCVFekDCh0nONP5xqMQLkrR+IhtWbzELt56pABc2LDtHDV4XPBMGemCbbB8
Pp6w5uMY3Kd0zfBwph28XYZnFTCdz9hZtsPNrHC0me3SAc4e3pZzkcErP3xJfgB8fWU+a3qRBZ3k
Ka7403VquVQ4lVuA3Qpb4hsv2e5XMtFPO+YGp7bDs8++EZzuykl1WtMAEmkQGteMp/r3PDbYnbnW
FkIjJthQdnVA6UoTEaZF+ZPc4vDjsI4YWp69Fgv6rFeKwKcWqnBF6iOxwn2scfwpQ0nw46g1S60X
OlWevyghtGeghc48lZMFMi+mH2nm43cOAd9iHC3mov9iFm9GIdYxo7+eCXAgJzEhgjr+QGlmpf5S
o+p6LUzevETntCnmRhaOZZ6zNWiXXjhuV5su2wunBHiXiCXlgxvW3sKm9x04yJyCjreqJgRtGrme
8EpIGNq/luMRz1KcY4kYdJ91O8eS43Vvs9I8g0clJFGrSyRoe71eBckSxpuo1pqL0MuNGK41b8u3
O/Xqe8uVouj9S27/6O9Qz9uebH26QMsgyEeVFBND8Hz09+H23OnsGmnYm+dZq1Pkgmh72BtR0QwL
W2Q4eOEJYN9g3jFzJdXS5zPHP3ZyEGbDUA8glepws3B98x/QiE7RMKpL3sN+6v3AxC1yx/6JHaZ4
txY2dVwWPfQt+Y7gLHXfQeZ/8IuNYl/vpbmVXDGO/FZsqn6vM4uAkwoZiN+mxEZTp0OZ/uBCTAWc
mKmrRtX2WC/H96qebTz+WAg+VEaAKQ8xSNe4kvaf2y3c28AHF9O72TTl/8LpHu//y+VWHaZlOSGS
pikl3RKMfHeyM/Nvw6LLeCaStL/MLYM0U0K5nMRyPiIBBbxQXA4D2lMfINFmNhL1MsFmY19wTxJh
Lg3P7KwOY+xR3l2OwMYL73Za6O+faJb5csRtz6QuBwPB5/MoNmym952nMJS5Wt818VSK52i+iamy
br4cXCvynxiOY7MDw3WiBCBNsw+LEmpB4ZvT3qFFbch9+8NqEyolDwWnT1jbYcfelgursemUzkDR
UpzXN4dvZC4or0YRJL5+4jywQrR8xDezKwll1J+9+QZGydpmIFFTzNvlX0QfWMh6ApeTlMN8q3Hs
fJ9VzOyMUCr6nU3hgnB1dhUy/de1HKaVMpWbj93EJWlxFmuTMuUocbnTLywJWuV7bkUb35Ch+5a1
ihOUGhmsWpnuWg7yBiqvtmdMRisA+LkUy8QkffZoCuL0X8kZDlUH7QJDLu7RWNYRMghZUayJ1xik
JYRqtkYpM0FMy3MfeiKt+/rXm3IBwJdnCCdVNSfYSN/8y7734jj8VX1wfRaDD2t16DRaRpqnkVv2
/zvF8/DMjPkKVHy6bqLGl37sJ+hN/Z8fz1A8203AF8iZcDUEktEueANCmWPQxJsnx0f/5akQxo99
1zRNeCSpk4D3Uvii5XSSgw6CAj/8ECZeRPYLflke+6Y3QltSLl/nJh5GOmeNdT68tGMAp2yNQ5BX
ZIwnXXPKVQ5LJEjyXbQYRLeo9Fs8iRccZrgACEP4I9520D1CDdf5Ngt92TEQ7WX/3+ZefodKpiDt
8497qNIsnbKOXhshEZ/MFUa4YAH13Mv3I0kKgRLVh+nP0P1x9e4iWpL3sL5aB235GafatB0rao5F
53w3nosY73LL8WY9JuuODgvLHQHzprHTZN8NyeMDQSe7jJwymlB74ImmSAMzzxQkmEmC9AZxgPDw
Ie3acem7QuCXHcs971objnujpCYm4VPk2v6596mpZa4GVWNjtiun+WNtodyHzagJg2eqTeABzvb9
pgr9osWMGF6nFqVWB6o3QOv3deXv7UHg5yZ+IaGmFrY7HA9L/7d78/1pfMVhRP21l9V0OaYdm5gm
neNaARWrpiNPzMJtW59wbCkJTCyE0zAGqxeuwQPS0ny0Z+DH6IKn6fqfr1Tvm/eRKZeCmftEvbqt
ak2h3HTI5LSLCOQKdLmdK0XFGBy4xasOjkTZMGUXA7ZjnU2QwUr2d2eCoPvuPO1nV1h7ufEda22n
nhaABB1ubGNf53JXATZpyn2fy2xpJOmEeqGZ34xyNHYKKV8lwaISHGMEfyCSnYj4/1eGmHr+bLtU
2mb295KfKJ+FrKietDvpRH+o/0ESow8hM0znq1A5ug==
`pragma protect end_protected
