/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbN4ZMpxGVP5KmyP2VwphtR5KHurV1Wek5EFhsJWkA9s4bg6OUdgDRrCa
6b2wUdD/+m06OOGPiLBpXnW/kI7Al2una495pWpbc1x5P9eHcTY1W6K1x4BnbzDqQB3unLWQ9hvl
j2G4fgtvMxJC3AIkPhCHbk2SM55Vfg2yyVWfPMuPZ35DX1EQUq6FXZMawV5uoqnb8a0+TacF4w9O
poTsgQ3QzEh6XXTxOe3Yfc4m6TDJTSQHx0lcQb/sMJwwIyQj3lL3uZ2/yMdHTU0rjNxyVY57CT03
hT4zNOdut1R1i7rim3e9jCc0ojdV4FHdDEZ4/ttEwv1Wwgx+kFfKUVW3eh2xPmBwNuFs/wAhavKB
6lcMz2hU3LF02ApNnjDHxvGzmBGhSDEf6InzFFzCM3UlOf+RKBgefugRzeT9/boxAaTo/nt/+Tzh
0bwI8tis+MYkKbHANP4XLQ8JS7YKNzLloFEfF1c/+uoSIOtjfvz0Qm3CV8atSVPspA5B2olKF40N
lF+HJiQSH0RcJepB7LSqgrqFehpJBb82eeLsdRrwUSjYWDbFs75Ma1cMtz/oXZpWD4PB3wAZy4fB
O2rophpbQeE9vuoWFZmZlQ4bJx2jigw8lVMb8vd6ohlvTOAKfOF/Nh4JhpRJ75Z087G92vOTXWqY
Tlrngv1HOVuclxyoidO11mnrbCfLsD6HOSEXOyBSeeayGdR9xavAmtYkiqFpNDuz741ahZZPUxb+
pyrRGoH99MBxIf9/ypQnh/c2ir61DslVKwtVmuXF9EspT5VJaq4yzddkKT9CsRtEhyJ1mYuHG+CT
KIF1loHiUPZGmdC6svFzYZzxH3Q3XBS89QRutgEY3HUtFxxCh+DVgP1DWrNIZKBZ1qW4W1U4wIyl
v/1LLp/2ohpcmyb92inPvTuTv/yDIYwDMHV2PmZdAw8WUXB+t/RxEoKap9O4sH4wNJdjtJ3advOq
x16F7Eo+rD7PUKEXDcnBoFtAtYEU5LTLqbsGPHHdrjn1XJ1IGGKiRtVc9PlHz9Go4B3Jlh5eph7U
HwHFFHPFtt/Q7cDvKRuljiDZKx2hUW7yk4Q7QuohGUB1yD2wCbs/EGEgv3nUS2krvWEJA7AtTfh3
/+TG6HJwZYX8gnW2nOacytGZjRsOHjyZmHhCj/Ko19wjB7NvvkCvtMmp6QfpCr2AFF3tvIichF0u
SN/oSzh30BaOhqlDEblbkhk1Ax8ezTJgDPlIfeZwVFlvYQ9UiivuxiIpgFrTQk5cnLxw+/MZQC40
AMAJ7/zfsUvS3Vf+/kzBvkv3vaJes+s=
`pragma protect end_protected

// 
