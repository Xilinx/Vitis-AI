/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B60h4NE1NVOoLIyTl7piaoU5hoopR2BKwKi8hCmg2jl5/Nu9/go0tQFwo
WGy/DYmAG9i8hrwX8g3KnOlQLfcHA9LYXiYHLglP91U6iFTcj+D4VO05NN2Jwy6urFouB8rjSKdC
SpnlHmMyvyXMBVBgpVDoDANzdjqhc2gvMkBjo3barngb3Xc3n/0fAVn3cwSjUcAxuLAO/e1/vOq9
ivqbbV3+9/7fDfqSaPmkkVabFWfAzMoHoii/aesx+Q19Kw6BZ90vEdtjSY7/d8wOdBScxhpiKwT2
8gssWPvpDVL38tgWoRv0hya9t2zCQw/ZEVZqqwYPBzYoGgnBBApRSHkipvAPBlXVSksrugPgDsXl
AUyUYzQxKATZZggPAFSr78m1J+uxQNA02HQWKfuShDzCCOEABU9hj4aavw82XJT27isz7bUqWNSI
qED4sxBOLFXNSqogRJlfFHjs5zUxB6v9Rcq4JHydrrIBZKz/1/mbrPFxHsYiTspxrdTOl7ndoetX
fH7t3WvdpSn1Z3X4MCkjRGj64sBalNy0OXdWPIvHNy95XmgdAYIpNiZpZ1f0ubQlY5KHpsXWFDiU
XshSu7DZhyGdUFRExY5YEegiGjQ8ohJRQvRcIDT7gVgHOLHH9vJhZ1/lrmM9i/vTTPK/AyCvvXaQ
dPJDJsvt11VotTY6SNXEIYDAntoViaskuMbSGoZNkG4vrNauVn1N9QbJHFw1MMqzE3uF8HsMv1yD
J323/jmyOIaV9fzIs6k6W0lL7kQGU7Yg6mDsTQXunUmhcGlvEpSsE1icZI3OYlb1Ck3x2yG13s/M
9XZ1kJ2CHTAS6J6JZaGfN+Ve/rQv+TbIz9/16PHUqxG918hIr2z/SkZDnZBPdw8K14MJ8RUgHyiq
51VGAn3sSLHOZ45Rbu54ja4F09YSAqWbpeGFqazu1ZQ2j/4UDIMUa/qHpWuykpCwRF586nzHxC1e
z58pZKAhikVRTjQiAGQcqGtcJ4j+1EECyeaZoNPjWJEB8OsJo0990Enb2EW543Z8g5YgkIQqhaOB
G1Tl9n9m5kZrLnzK/733qBquR3cnGhZKjUwmBqm9BV3wrp42n/b+hR2p4AU6kgRoGJJrBG9WMRzj
LvlYrSS4udAB22L/a5uXP4dRlHhGYORr00LSxi4RbzmKIJ+pKfEsfclV5IseFgbd+lKlUAMt2Pfb
voX27UGIztOrOJwETBxcgFvnJpSU8ZyZM92EABWtGVB2bhqBk5/ZRknvHqenhGSxbNDYVI/HjJwW
FtzrSS7ip9rEvJrEV7A91OjRx0tWNtg=
`pragma protect end_protected

// 
