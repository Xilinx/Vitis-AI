/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2tI+yHFKW6y9jwZuuJw3bkxyJxhnCNy5OoetXWRQwtjZxQiMrBJNRoxM
VqeU4PIe/3kh/VMlKiVGwsGzoF41A1xm4pZo3yGS6JWHycscF56au4hQOBIVK2c19FmNvhE8odqO
D7iqYcWZZVszatWHFBHRRwFU8Bgf9GC7b2fDR4xmK8YFmyjkN18IexTrJg3vRnueB2ZNBcZ7VC/2
lClUyHD5/e4dCnaEx2+JXeRrEyAD6fkU7QB8bULZSuv7iKKCICsWjodawYtvXnSchdrblDQpunpP
olUSuQfVaYlRsTuEaeJiTw0shDDMthoEt9JcDccFldEp9UkQceUxkCEXkduFVJNRzBTSAI2GSSjo
ln5eTrlbXAt8z6hfLlONrHWizdc5rPdIoNXyDJUpioxtmdWZMIoCsQ344WESPDXJz5GTZgenDVMH
G0sr0xhBcsQNyeYbsHw44+hswCpUZudK6SmM1FOg5Vfrf+LfA/VvwblKJznNE08cD9tQ3yaaKEyw
ndcmUTRnf8ZUqvadhKOUERmf0S2g9p8i4iqoD/DS2N0chgPy72b2rH+wr3GEtoIr5wgBVmooiYU2
U++katqk3VNYqNIMlL9tnV3H+/03JMS+tvjCXHcI5VSvh19t/Tf/QmWT9XqdmTEHTiJmVyU8PiiZ
pppnPlDEX2a+wTE3o600nY+VGbSDh8+k6uuXg2kBPGNiLkSz9zHc0adbmGivo72OZbjVrKJeF2Bn
Iiej75g380gFA6CAuEuufm44/+71tORimX18eCFO6DzVJMOk8Co4GMs7kCzgg6dwCJSgxWl8fGjQ
j+jsfAD3Yqke8owPjY3v7ArFUN0iOtYd8d7qrA/1UsNnHn53cmp0yBQloiSddWCgNejoueBDEX1W
G9HK2kRuDoGybN5UcaUHdcUtBEtrZsYVIRafNuEj1jIAQG0JlBsNbYEuLKdzGVrCKiUV8gWKvqjn
QUWOIketNSBB9l8nLA0gRfgSj1CdJ/VpBqGgWXk56jATZw4aHP3yA9V7cO9BWFCpzTAZq3aOLaSt
kl7Xz8Ay2p5OtKzIkVoyfP9hsA8OMdAVuwOekI5MpaquL4NUczSQhI1R/8ZONUW4GQlMDuS4h0zF
2OLGde59TVGuQ52QFQ6d7kKYdbBtRYARIMffKc35MtxKTuZFkR4sgoH5CdpOwWhUBjI9C4Adt5rn
5aD1RjmfGZduux44lGfg/95Rlp/S5N8rLQiwoNkBJ5gJCOs80adDauW7MNPSAdSJhUhixSyx7p7z
G2cteN1Azwpn1Vhp8krEqh8/DboudXs=
`pragma protect end_protected

// 
