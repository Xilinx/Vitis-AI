`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+GzawGdEcIuxfE2xohKZ4YfAgNY
udze0/JpwAsGtIi3JEG+f9Lc7KzDtVo+7e0axUtpWWG2zchF7YBRjZ26kg5u4E7NrejsKmQn4oFZ
2qTRJZGb5SJ+gdQBQzowrZ6DlCm5Ybvng4Y+fKORBe4O+BxCB8HAkjiHJvTxpq0VwrUrB2IS9/yv
BT0mW1nWT9cr5BxcHY80c1SIh2SWvSjyo6t8HbC5zSeDNq/HCBlFXopiOaiYhaqw47uoKfrNcZxV
H0qhWKBZbcORMQm9xN+o1RBYSoXsn8VfCT9g4jPppSBt9myV0dn8DD+i2eYjMXpra9GUttCS3bya
TvIIKA+XHS+9gej/6n2ZHTWhTLL0rGnF0/8a5ZoJ5H37FSl80g50jY1fWnBeKtRcxiITsTi5fspa
efb+Z2JBZFuYz2m5t4cVoJML8RyGrB/PaylHCC7fTYz6H5Q1LLyQt578WtpTWqrTyi08N9GtcHlB
hTUne20xL0qjdfR7ZN7VLM9YJbSpkyVSobJL3d0S4/zQXW6wfOwf072oG0tfWwg2FcC8BFHx8llq
R3PGYe1Kjc+sfNss19AejSO3WVSgiq3Dsj3Si/ECw5gNa0PMmdkoyb/ftqkkdPoOuo6Y0bdWGsNz
48zcBQELYNi8MgT4z+xyuMbNo+EXxd1ldCHRS6lo3lTH1Mexj/kJ+Xr5Dkd3R5foPmPD4Jo4LXxH
VnCks4vL271D34Qf3e+IH2EJFr9Zd9w5jaUHVbJNRrXUdzk99fYWebjgKvbt/hyh9hcwMS+esI/w
XUdzbXttXPavlXBg62mmOaX0PmFOUNVekt9I3InHw9fcWR2SXSbEO1eaFqlB5b22uy2kCUvD05Mg
ZJQ2BAp/S7n32iVxfje1g9ZDmA9Kter7dj2CYeXNPKf4jqySIVd/c+iaDgNpwoiAGyjhK3HkRc07
v3lzxhJfP3byUcEBT28KkRW3Ya2TWTMoDrtJCsXK8Dvov1Vopc/feEDFseCarx1xihLMSU3R5+gw
07G71wGC95rY6Nd2/Ee13vCwngb2Fp1ya21kzSXo83xABGT1p8n5zgGf75sc5V/DWsMwoY0V7sCR
ADBZhVnKI5kXNwadDc8u/uDI1mdhlqROT8IdHWAuqNg5wju1BDXbOsq+jx0gdgGrMi0QFNXIEUNi
cN8scIslEMucRT/fcy9+s9TFPuyMynKko21hZEB3aZrD/to7uLZsv2orXRVeN2y/mnScQ0WeJEJA
VIjm68lVQCkPtfuowh7q61MJ1kcOiDQG6WsKCrSfGMRELhrd/5WqjykvgM4ZvCNu0UimpJj/o/m0
0Zu4qlMmWNr/Iysc0HQYlvZdZwRJoLpgRAzoWDE4ntGoXyzzdzLxZ069qwI+AQVIG4R6RCEXmJf+
R1W/V1LgwI4/GYi2rg7+hRs2wj1T+h7WHDUtgfDLlRksNGDlkvS1MR6WIEqH/hrDuGrLiZzKU2hA
4syQcmbH8rPRjIsRMKiCjanYJ2KPNhFJ8jssLh+O7YWis5sN94ghJ2b1H7MjG4eYX1FCUZ1JCdAd
9B2Leh2s0TK1R7BDU58k/HXxjzyeZlrci/RlFsxPGHmdi0GX4Pz9qR0gbyGW5fqMLXguKt8ACezf
gRoTWhVaFhjjnj9D5FYVvW6jBQw6dXlGKhvWWodMAfh26+3GEYHj0z4yLWx9jL0oGWtcww0aLETV
xVthURy9uFs0jS5mjUXf2KqI9b/TYM2mxvph1c8ekJNcCsBe++5Kv98N/5ma022wBFW+iBplWAQq
s0X0XfUj6snaH29h/Krs4zO5/84RcArF+91CBvk+d5L0N0nAJ08dNu27i9ZWvL9Gzan+fIY6AbAJ
1607KKcct+06QD3m4i4oB8wpZFgaYszziIdsqhgDRNm7knrBWiGrarbt3RqTrRPWd37c/BoylTa2
9I7F5oXR65MoaUKDXFAU6TlR16QJq/KSlBZt9saT4BxgRpeCF4khs/WHauW7m9SM+YtnDxRHVPdn
LQq5tU8+AW8glKnJF2QwEui1LyReU54mJRCH+BwuTg42RMKRMqutMwiZXff6EvcRJ0wo/5laKD6M
LbRphc8gzs7ZiwNRamPzLaSrSCoEcPWrP7Ve3Bt6bOqbpEG2YeabpRDz5E1tNtoURCn+P7ldldQ1
1JV1C24ajRDE24jl/OZX1AQFsquAzVJicavU/En5VtHuhU127bjUthl1VNV0nKbtz25ap6HcaH2b
B+zk9xsDR7XC4RVcfhSuCzN6Itq9Rc3yud5afXGUaDQrHQ7VeWXBpbscvRwkyEG0Sowz7tcgZEMD
l6pjM01pIBqcmJCD2KcxPFRGDsvZU+Nl8VbGJJO40omPDHf7DlRxWMiiX11HZPUzRzVDrhbR6iCS
xuut5yaEerbmfYGZ0Lx6Q2eam15kW8LYKyN9PavCAJ0l/wHLMfg7K9fajL7kgll19VXEjz9i0C4o
5bdcxTSP6j78Tvdoo/SG3PHjrQTf8uGslDZKS4FIR9nl6mfIHfVzqjzpKgHKwiBvqIH5fNpeVEnT
6rxL8spY0iuE+K2/FNkJeZ45Ia6xVXudOUkrwqMfZ/j+hYkkYsiDB2Sigk78V+FmxI+Pm/XfH/7F
h1tdJ+dEOMHeCg3IK0Wxu7XdWjzrRtsZwHHr8RQMNz4faWQybddL1dm0VINvxrPkkuyVr7nn67D1
9nsN7JsRzuTCs9B9hCWBJ6IoQXA61ip5t//lRMzscfo9poVzb2ywSij4PxMG6qoxXlg9pWSIJMSb
KQe2ZBYrs2Tlxx0I2Zqn8ztbw3wfUcq8Jo6fvwaUWwTzgtiqtxFtoB8m9cAy4KG640R6yNBSKbrf
/oQr1P7GMjMNPF1qo6XmWVII+sPgvejpJ+C1N20evwHMX2oObbIsp810r74wPqyuYm2N8s7JqVz7
Gz0y9Whwg2wqZKMj7X3sqIvuZpLUgoa8Y+/Hd80KkKNmqLY4mIXhBYmVvO3JgoBFvgBhZyxYPvvR
IrE/0hmrrPOBvIzLPA9afNN2NvvI392ID7rJmoNMjun1p4XmmX3DwkuYpxbkeVFWXfVzFeasdYob
ggeJOr0jzUjD/vws8TnAxu2fEvMVOkNnPgoITnagMGYtFICdBGwyJOpn42f37HpB6MDp9Am3VxOn
utRCoxzLJPB6P5DqSL6H9G3HV5L5oo2R6cGvel9lBD5DWiM0px06O/qUEXtuUvc/3XPEQfgRSMeR
jTgS+1niE8Nq57M6I1e91PpQNlAExkCs+tkfxUa0nBuWr0WBiuiNIMlVR8TBHUp3llLB/CifUDdQ
xD7TGxLCYM5NcTlWFnS7jvPmjsUYxT2OGcxOYsQzxgFROS0um8QOnsZ62ls65u68i23YHCIsXHqX
P2CpaGJRn/U0T+qt8HCUVatxJFlCtTDfdp4Ejh+9xTvqYv0frQeFJuEHVRAC3hndvLbBGXNYgkgB
0ZFtCmJlYtGagBPUebExoQRF2ieD3IZ6c9CBmshVTPdQQH/taBz5qXIU0h1EZwBitSyhC9A4mout
ZF67lq1t+m3LstQuzLhsl9P/uU/WZ78Ro5Kd5XgZWexSC7AkxFoZP+y0buXtfatOr/JgZwCP2hly
+WJup+6gBfl5W6Md5dF9wlU7g0BuspG99T/zn65HgkG6gtXVVyEz0WyMgFO3oSURKj8+pLzESB47
8v19mzwJfGDRIEE15wPClnMsDx0MeJxt+cbb1w5hweNV5hmp25JzkAmoIvg+MhVgHYC0sQGgUQTY
3ujsH26zatPoGHlkI0hzNpma1LltGHFncCAxoyQWfmPk442JCTp6S1wt90lAMNrLV/9ZN0Ea+vpZ
jU4afPel0YtFB8mKztzXXqIJp7f47Q4TiFQREAYNzUzWLYeVKP2W+ThlGf1+Huy6ZocmouuQP6xY
MlLYuOLG7gaNIwcwqzoxn8/sHMiaiIc/FmABaPk97IWr/P788Vt5aa0esgxVkZ4JgXo9OA5sUhaG
hGh6XSzROincZLcunhnunvSBD/6hKPVzeT0IL8B3IGJQcNJV/3gzhhrPEOiiZhMYkunmoKyXP7t9
vErAp6VCILRAcWF7a8hZf7mN0VvpnfTkKAYy1gyQTurBv/6Bd4gqR25S7ys4KCk5jnOXzq9HvSDJ
BZSO5hlr+gEVin5HdELnBf/YuKg2faY5kjGWV836VUe2B9uNVIgoaV+dNspi8J0WncEma7V4+Plb
4A/Pk36MhxLbgH74rzQjBPkt0OCFaFwaTYmTgB+KZE6glQLtAGyVSKodGEOsQeDFtNQsnvnmV16V
Z1V5QFZkzWW/E3VKP2OnSQbLqRs37YcZZLfC6zBnt759It5CVALDK0X8vr9Vg+4cLIqRS7cqj/Y3
EWaeT6bTkssrkPD+/IfHE4xPT2H0IM86ImXnC9lRna/+kNqpYzB7Y8DCueYhPCdpAyJrw5U7rc08
w88sAlHQ/f8kq7KFCawD8YFcGZl4C8rMRjHKtFcM9KiXWFNxfLycm+Ngi4NCAx8qoD6h1sBoSGho
94Bv06ZRcU6F2NZu9O5XnMXRn8YT1CCy9qCjOcfRAzx6wq/h58GdrRELFbH2AiBgmUenPUolwmhq
eHH4k/lnHjRgLk7b/pg5Wxvj8lGkbsviZ2+g/g3G+/VwEMQ9m6NItY2nPTczzPkrCKTULgQB/638
OkgdFX4pjvffi4wMviAcL0nR+50Lui1EM2ineJ9scVofiaCj+l8npqkWMYtnZe32pNUtz/JbOyQn
1sTg1UTNwdlcmJCMPSPLI4b3xB+a+WOauY1s82EHG/YXV2Tg5YRZjNZ0Lcgl0I96r5uROFixjxwQ
kQtlKCx4YYloHMadCwqK5gNWbrLI5gACvmpeA+9lEq0p7QP/swzfAznPqVZFCw7lpSLf1M3e/p0N
NDMTzYkBkbEIzHW8jtJp9xQI7k+TmCKhomHMi6iAcJCzZ2Qlx/fwYuCfQSl/vU1JB8HQgs53yJtH
oYkDR/M4XqkWUATBwPitMGjj2SddP4Kn+gDPORJe8n07YC54wzeLxHA7O1Sl1EgbzSwRPX/W3kc7
EMKfqWhu+ZPOxtBIW420TOoCJlxHCCS9kJB1xsKoOOQPyUd9ylCBJ0dp5SzTCVKwH1xJu3tVD4Fp
T9rFnGqj4Rx7hnSUZf3SWUijkxY1mMO+wjpA1IJr6oy+1y7BDJN5MuCp/45/yoWFxK9csGxN7hSj
Z0tjzbZBY4XOE4wRuL7gCAe7n5sSKdL13U9IlZwKJDsyos4xRjfJRcKfNsBiFMeEsWY82WXcfZ+G
rMc7BpWwxyrYIiBmyuUY9a1MowZRFw8yls85ILaYbTvHDi0NHtoAMqz9J0Lwe10LROu9KBz1pALi
fr4gzpF/eQ55Ae2uvDjT8Ot+OJ/wC/wNBzqPeOCDuvz51+mSMVtQTPVQe7y7ykD9FYaHX0aifjm5
KgcYNsLukPhiBXrOJDOIbgSWOmWIM/lUCPpw9BjqBuI10RFH08LHFRt4GI0FMC7SH4ROcPALNHxg
ECY4/LD+9l+wG31kAT3cTV/7Oto1sHyUzrHRaao1SYAlKuEXo77TR4YCcaNe/V/l8p/euPYQv7gr
fi4l9F+F05+ACv3ob9sRWYBLGvkwwRocka5TAY8c8Ng4Md6SSf1u+z615aZ3NFAk7TXoqBcH3GEX
BFLeAd+pZ8ZAzpqePzJcVc7szaLiSIvRZ6PvtNEo4HeDTAIWnT6P8Sug1y8xcCUCiyOPk013A5nZ
b9J0YSr52VnOBouQMFjTWXpoLeUmy3WcHkZ4oD9JH5R983LUTxbbM4eZduYywnSLNyWDTbVwzsrU
XoWqdmoqNwuhtRU7M6gxMidIAMSaZT+a1IzH5Oq+uDoI71GMRpP+wcB1+qgbqTT/EW7PzBXd+HOp
883gFbVIdmDCeJK4tzufFOrEQQAnFEqRSOtpY3lYv/NfVPUCmSpHPDxYmPSpZqZ7oUPVsrj4DoY1
5QXyvKQC9gYP8u01/GmGJAIbk6ftFO2xoKQzn8Kj6F7drHwtRxt5uA8XY4xvSyBRsOZV+VDV7/N0
H6Tim8ygZ7G12NhUcIIQHjRGe9m25uatShuXQzvILeT5de8LRvf7XQPVty5+vch/OoQZV8ubS8CL
PI4qQOvcUXTifOYcqKEXN+aFRJSZY+fiRNDEeBrxIPg9qypCKmtu9hY1L8TnCckpE1nxGFlmK70L
YX9z5eDbA4/f7pfgCatuOxXOo/8zQzsXJNRUGwB/iJaJF+zIIYIXEVals6BbbCekx1R8bfkCV40I
yn78zTmn/5R+WEHfvp7gH1BuA67Gs+akLBT13KNEeGPPP8Zm3KZtm2v9EiBzYkYPA9qB6L3T5MxU
oLsIxtP18SPEKt6k4RboSQXX4zlmsTK4lHTc6tiZvm9vtLThUw27fTwXKL8hM8WjYlGQsDrxi1f+
J2p6PWpDT0H1TYiwHkkzGm5IS75fIe0+MfGhoNk90/cN1osZfN7qHijK+ew543CzCd8eAqQxYnYO
EQ1VVaXKRfn/ZQ/nV40oLLskWbw/rM0t6LvAcXSTXX+Pffv80r6bkzjTC4cRBVOaPh6f6UpTHLAZ
V6XirNe9UGLSxFs/NEg2QCBU66RG5DOypkvqrh1Qn9eSIgr1MX7C4NngHrHSz62QdvYHVyH1I+VV
wuRqcJbpVP3i85lWUqRF78F7TjPml35YnWDft8IqIi4/uxd7FHAV3DrXCElFCS2dw9cegFEKhw2M
RJ/ocv/M5o3aVM79nJFgHnxM1cP8xIbNGTy+bOtM62UMe7HQDru4BHqfFtG0EATye4nujqpGNqXh
cRgAFuaFrVKVrvOBErCG9jFeBp23oYpPVS8hZLa0NIgapjbxMY2OpSj6C0VsqwiwqLkxN4w9Tv2g
ViI3RaAW+8TxxzmhvFVJtAmqDoc4b5SkIOEHlDJWZ0ucRPK7Pu2rn4d+knMJM5P159wgga+dEh7W
DK4tHtPwpRinVO/O9mEXf4J483pnirZGrLiBuBusY9JqxVileuBH4RuIdHUsXIvGZgt3fEPhI2RW
1mLdKTuVpv6Bl02aak5x6ClmFNBAAmyET1gxnJsuOhOxqgCGtC/7drPcpout+1EsesoYK2pXdIDn
p8fciVZKMCn0SrtY3yFNMwY/ajH6q4kc0ehbqj7HoqsdEkgELjFgheSFiRohlqG1qTHz2BQoQnIU
pSV4ljZvQmiTe1WOwJ17yuHd5gR//taMzuNolTYsF1SImn7bACB6i9QB8yZBJaHc2orSvG/icA8M
tYwKZYyxhPoS3J2YFg9ZHniIf/7dsYAqwgNuGeTOGKxVnE8id6tpRH8diPlrp7HPGdoDs1LZDK//
2qOJsppJyhfv6PljS4P/nQe7iFAI2kZq9svi77QgyuktaNsmwjz/DXYelVnf0HKr10/LO4KGDn/5
vkStdRPAlVHz6oKJ3b+eyecz1D+ziMHd87uY95UzjGKwsxLj7kRPZ78hCgDCuvCNr9zTaBNzSIB6
CiD4ES9JQDkrseFyzTdBebVSfZ+I9aMmxcq++P6GKZitSlZa3daeGaxLpBG04v3egxLwHX5e+KJv
sgO/KsCFgJzuC/bH+DJTqgPqYju6i37gWCFeBf+CavXAzvdxPjHaCkXhSgSQbZCorrCxvPN7j9os
dlL7cJBaW3ZZAamU/nHXXVi6DRwsBKsTYEi3swBmb1pZPimMGPGKUihmo1F6n9SF/dasN25CLG24
HGJyZkjSniOs6l2d/wt3+sRyDJy+oEj9FMowPeiKOS2NYI8YX4v7Sh9Sz1O5RtyHqMGrPcksfZUx
ysiXdoT0LnD9C0TrC92MHm3DcFSbormjQ3QUSSDNGTlmKtltDm+A7zAjpI8FCJKOPG7IXk5/4w9q
CmLucVaDaXTo5xV/hO5Muoy4X3FFAtxIlToNGznyP4tzNdcvK2hVDlhbNqTe224MmL5ctS/S5D5y
ayW9Y5OnXFfKV98KG3+/AHxGdQC1FIa+cmiY7HJZNViW9yaLLDVY2BFmv53uky9OokxeRmj30ZlY
oYkVgSJtFOpi2fjWh/96Okm+SDnc/tpuzgPI78qpCzdFm+VocNYgQD9rl+clErk7C0euHLvQ9AZW
tcMUWY4chqh1Hre0fcGaxjaqJ7xkAeyBBa9Mwg2kA+Cctnzksv79S2aTIUS6BApbZsu/r5LbW/gX
Am7MpBYuqYBlluCGRJj/ZsLarF4+8IfDYDhsFj3i87PriSQ+B8XdybCU2c72AuZQAlfNP8CNolmI
8bDGdGarE64kWR42g42gmIDjb9iCSXdQnAR5JC3Hq7c57m8TitjG+s2+rubPHRCudPtks8QxjTTj
Dtra3WyT2gS/RiPZDhPxmujU+vPFUDGcObKsXlvrB8bqNMe/vWD2+O+W1Y0ErBl7Yw3Od0NVwY5G
Tup6/wlSDgP8bMkR5G7IUAjSvjPmK2voZySt4J3cwi8wz4v/vdThQZUD/Noi4Rm0MnQxLUfqApHd
AkHwWUVlfKJVlFtRjNYF3yU4hsSMDeKQ4RjYlab/fhZU7oqMjwgiYXK/RqYhPqfAXNNohhFaY6Fg
jBTNXwXPFoU+crDI7n238vyMHeFkJuBxMnL2O3QuJQnNKyaEivvzGPKwIAg+TjvDqHiKOY1okmr6
Y3/owDJj6MyNAiAHzMWHyIA2QhhVtS31dTw9WhR3ywVuc5WOX2M1ys1/pkGCSsfJXoSf9hyH0hnO
Avl4MCYgwxkVzsgPfCl1+hwGCqIEVxux5b+rng9VLc2qo9y+eyO2nH6AeGnnTMc6giz/OYNbNddH
IKpGXy7XfpcysT1xYluLD2bDm67AQXyWNgwZmB/WoaHq8V2TC4MqjpeN3oQd4+FHvjihDU0hTsh9
8sUkZfM9qEOaRYnAdRlZqN1exB3N4LVuXNuwMaNTl+jshM1yyR66Ifr++5x+UxZWkyJvjfIBR+8g
tkh0thhH4dmE3NP4+WQXXeA3j697WlMg9EuAIxNkLQFbuqJrs87+iLn6tqjiOH7+zbKJJwDj7U1j
uUQFuP0KToNODupsVhw5WQlXxqqvUdwGQVbRU3yfALjEkSjUn2F0vF5lIvQKZifxZR3bv/SuUNvg
vN9hHaHTVA2MHR9aSXlhVgA6u18QDb+fD7FotAxXhG+Y3eSsYcGh6WYECCME1nUfoJHlOPQreKEp
+LgMz2+R7VL67Hp/P72zU0NvEyDF9uIE5W0NIppV73LwJKiDDTH+MjoYmS2wIiHvCF1kYpKxP7+u
fOvOulMCUO77V8QAOCdQeet20TUS+9y6g3UU77sfO3+RoGObPDCiwB7bTUWIFZQE/tbWM6/KdpEi
nCtioFl22FAe8M1f9k+7Dg3LmJqyGpL82fBAuA+mFUqR1cLv6/7twTIPFuvUQ1zthyXFn/va38+t
nlc31bwv3/bznz1c2WajWniTNCsL0kS188uXi2CAWebw93nWOrK76wv2jLJWPfYStwVxpm80BRB3
JFz8LpxKzdz/jPKBUydSkGA7N0ULI+pa8fTGLvbdk72muiUh5M1A+UrZEiPtIy7oJsQy0Lp5YoOf
LYkHV6NThAevOL9pLxcsyRCB2sFbQkTpG9GbI++vUCnnWmcAdvww40gUfT73cH1B2I6h28HqJul5
Wlplu1jshbhG0kwo9gm59BIelo4bb4ggvgMAjnDKQKICmyRBRj93POdUBmPkr25yaDXdlnFGpt5P
e+bQc4doH7wGxlVLXP3gXzCJgnJRLetoJrN6Z3/M1FqNshviDXundRsUNFwqQZjoyuUTSmPCuyiQ
klCc8JI7hAO2RRcfwqLRwQimxc0qkgP1Pc0j8I4wjw+V/ZU7hvKk1Nirm0vXXhCnIRaSS8X/1Ki8
bWYHEaL5T8K+brr7+otY1c4v06xz1tUJCvv3T6dA6waB/PHBoH6SKGb1A8UBGHz4Kur36rEvWZ0/
8g+2CytztNLP9xukgOTZw4vD6aVKucHSjJbw4LKG+5YhI/cGUrsuZAckT4UNvEujL+w+R2lfgJ+h
r8m/YzscTWFr+b89MTEUNo4sdSGrrUwVTrG02fdPUHZF5912vMmb58XUebZB62SS6pKjSZHEQ0Ey
Soy7IT/EBTLRyFQ+8oJoOx6hVNv/MmAKqTqANlagWr2yqQlfTiN/HUUmXQCryZN8zej9Xat8PwSP
+fxoGIsRkMrj48dP7fzFXTJxuzkISMu/nBZHTjc08oYeL69YuSQVcoE478aRvKVE0uCtf42kOw5H
LkG20Db45ly7FCWZ7YoWgGDc+HUahhTX5b7P2A0LNlKTTeKYTxIbmH2Fb5LONbxODPeFadEcDpeF
CEW6gRi1D02R01WnIRa7X99CUQ42iXbIiDAyMyvOpyDmfXpQs2drutyZ3FBED5LIDgvILG08p4OY
FaOAfG7F/TfzDAi/w0TF9mLXBvvjSvC+0m8W8GtsGEVOsjBWKAmXSVH+o6aLbe+zMy+oiyrn+T4T
Ljd0bog0r71Bw3DvuKh5BMNFt0XsoAHIDaL/ApuWqSfdW32Ugk8hWcZ6ADpvRVtCYXipctCuAvLM
PMizbqw2BQXzkaPASZ27jIpeYPj7zwYYTcwYXVyr7ZXiiupz2QXSetSrJQRNh8AUtr4BJxStSLkr
ZRMYvGfjb60seaSozGPQYmlwKpJvCcBl38qbXT/iq5sE4qV0hQ3INpshKNJntJLOZgequnW+L9YG
/MtleKVxCb6RYKtcE1eioElZLFU5A5q6vTPxzokCM0MID1oOL4wscVx+JgGN0txe14twJVdfSdxZ
McO00B7WDjiF6P6mDXm8mkEDuAnSoSGcsjr49aZfag/d/8xCADltNv8h1MDaOzxrL49thXGof9Mn
pSdHmBnvVZKErvk9lkqBJL6MV924ueBn+nPENVkzf0hRTuVfuhRPS//VUsqPC8X/YUdiwrBrhq1g
mIZUClE6BUIALd/D8ATQJsOl7CKkiPDSpLPXaZadtFF8tQq8WJtHathCjOsLiflmX3Jik/LuhXXl
m6wAgJ+zCeI0YtutFtQ8JZVzpppu1ajPFFIKdj9zUHXUTjdcuRLcIEheUjGrA6iEixhjcet/xcE5
IXrwBN94uhjNcrWwncbVtb+WPYHT/+Vy/1VTNzqiTbfHxN/yaT2xz7IgXhjTCUICRFE5OOqhq2Px
ArZTLWpmxwxjPMvB7TVOGq0spPKeI9XGtjzMEGSlqiODRMyO8PwK6+3MH4YUbiC6gbW/r+1A9E7E
E4YwXio+ixn/5U+6wGCbvyno/bdlpQY3bxrgfJPklC+lHBu/yJ5cv1VLPM3EeIJJCao0jYjE3VQV
2OhWkjFu4vyNildcIizRNsw76aJJl893yYUN46pMclq95KGQR5J6ZzGC3ve5vtnWXwA6hNG9+0Dj
1Pgn8mBV15qPEhVvPzqir86Em0KIVKOZv3aEzAntZC+gixdnR3C69fUFr1CIg46Efo0bMaRfJz43
ipWg7ATVHq7Fz0EON3Sq6AfKhyV+3K82UCqlZl4ki66UVUk1SeBS9j0pLz+pvUmdaceO2mNz3HRJ
hskF0tFWsyPT8XOysTwgezm4UZt3Hi9af7RcNvq/n2rm/WNgr0LCXf85kaBE/6eb0c/CjD4FgygE
ebrzEHVe0GH2W51/ARSOIfU75000fFpU0bbQWXfXA1GDOorEiUP58V7qGFWpiF24Uljffg1pMn9D
rCJjWqtjSQlM+Xfbg0Hn0FpL2hHvKN1W5ifkcVDMneIxjrqUW3eG1QSbyutGltjtw5Up8igxYtEh
PKCEugw0kUmPQbXFLKM0V2bl1Zk2Tv7SrkUsbQEFG28NHOQohumgVH0bjFlx298SS4BqtQF4ygB5
6FUbHAAW0Ec66DR6rid3ry4CRLy59w5pqRrOJiYTM1KNU4wbp+DUgF7MX3Z4d4hPebpS+K7eJpMQ
i6Z01h/B9O1fRFAsW73X2NYy2vvydh2bkznEIuLJWfwiWQwg9E5oNL+Z+Kxs+KgOJVFRvYb/r9ey
DSB5xoceRwyKhUqiFtkORaTTbhULrDkN3iKYGPY/nKpHiqFLhuGntVfx3anWO+jVdkCH4Ws9e1Ha
I1TLjUmUzSa+KDKJ252WZcevTyjKANtLkfEeIrgRG+h865k8ysN6oAcLEqXgdKYrpXEHXqdNS3ek
6McQ3OfYqvmOslVRfxPZr4tbnegqsKnPzcB9Bv8DNCdJbfzxrlHTG6jSWVBdIe1W6hI+2uBtd/T+
H8Mdu5I49haQdh1tR/qo0H2i43CFl1nGDvR/JDvyN7NnxPXNMqUHC8q6WvOvURcNv8evk3VvL8UN
kD+ta+vs1MvL3SyXjPAWKcvVtFIMxb5STWNXLAtfFp39zmmntzYjxbqpsBqEUPq7UiE564J6HAac
rHmSs0SYPR9mfHRvenJ55SNXwf4jKkmsI6+jKPJ+NMQIQ3oX7yzhHPQvCZjcB9eg6S9IqyRa6jeG
ucaXDqVuKd1zBGKVnyFVvitmI57U4bBuoEA96HaYG/5Q4wCJ+vupkaH9F9Ht0ELcZ4e4Ugli1NtG
xJYJ7836sxekTZNXVhb1I7Btvwy4E/vipYbNEMAQ6Zhyld+JzY5fw6GVhlxn+atPvElr5BXWySbz
IcUV/yfDlpfz2dKWAr05EsVaQg/r/mpq2DD+CWnKAPknRascu19KJDdPcCiYryyl0HtxWf+M+5Up
2vkev0otsiMf3Ag8W+88V28RTBbSa1qF7vkMar0iJeJwGjnnrSiWjYAvu41y9l835MSu1nqoKUKn
kYGx9fkF9+pJQCw35pBHNlfetmenXaCKIM1PdFfC1W/aIDWdbLcYq0Wq34823LpkfjAYD7O7VWi7
/B+oF1nsJQFY8axi3pvj0sJ3b1KcrLcyITP20twiAR97Hv71tSdIp0fPTWVNNKh3F+9eOAN+mMx9
Nw9bQnoGlTfGT3L6QNSvH0p1pyTDONgs8RT++vKZUX0vObSEi6HgpwscMsqfLNR162l9wJWdXEG3
YRifCODChMvDnBBSs25qyShlKjyswjLO8cvrLMkiS9wxr4zYPKOk5GXi+qe6D2JOcbvCub6erhi9
IaaXHx7eHomVF5Hr6TR4Ki8NuQPPUW8RKNTexn95S0XwVAzHsYpuLrLzLeI03pfMla27CTG/7FRN
ko6RH7eQ5C4H6FL/V5QUlDBztRK0CAV6RQ9OT3LDQLId17KdmVkyjEZuDSXkEWLYicTOv4niyAsc
zLYYf9P4/wVfZ1jw9O+lgbQmswflNv3PsM3IMtfjee7BTae40AehxRxookm5LMBeNZQhUz14YqhQ
bqISp/b3Ph/Hka7GpbyuBCcW9feW2WtnSNDlYhI6gTWC/ry7fpi9VJFzTRK+UjYNVotfOIWo+Gc7
OF1ycNebtuIsEbuOOPhWkSf4xs8NQDtcKrrehesTgHiXaxl7VqNV0cnJOmgEqI6X3N9I1GzEoKue
LqDNzKdFEqqCgx/uLSTqZqQXDQ7u3hsuNICVEgtMqMqMnX1WXaR8wDHV3BWYtvpebu/dCScZj51v
A2s/tNA6cdT8j4sILV7sNQo2DtI1BWe0np+h5xjqDC9wT+zi/ruwrxZpmPmgURJQLx4ozKtZcdNn
hTfCKPZWRH0W4J3Ibm5DafgCxT/RGZmqkRWh6tK28yhbP9wuYbSd/YvISJHw6OvFhUShGx9uj6jL
d8P9CGmRXzJt+zMl1iokhnX11+A22Jwb8P570M9BEgXPVOJnBTrizYmyqtQkygDLrYfDHazWHSrb
2kmz1UFrK7ihntWzOrLf272VYt9OpN4WBxL8mFOZUDonmlYuZF95s0d9dBvyI8xI5WZpY1D8esdM
ZLErjeV5c5V/olcvyoOiMpqRao1kHa85E0lJ+KLkKN4y4SMoAhNivtCol/jQnVJUlnQYpL44wJiu
ab1JRbz0CsPfdqJ23XJdmTrSbVs1wh450wzKnYRVdKuAzvQs2sFnXgwzZdvLU0AJDTj43ibzShm2
gkVu+XynX/K7ugnhJFsYLhNdomYtWxPmOTQHfgm4NwzF+r5A6GDwVCsFSP/JgvsamgilUXRDzHFs
6eGagQoq36/WrDbfDZr+4KWdLwyqxo/RV9fT20Ovl7hOUSvqvJ8sKIpM4kuBxSoWo0E4AUUPm897
257wfuifgxGpuwhMYj51vsXaux9v3tP5kqorgK24TD1jh3tXVMYz0KoWcC9hf7Kkvq/kHJ8PQfUs
JVZhx7Z2L70wBLva60fDbI1yppkdoq1lAjY5zBJjQiCCeTY8o4jLxwp8ybL4zJZi9ZtvaMVpXvcW
YN68lFzpQ8wmxjaYzy4MiCWMTFMTbSRS8rB1AVkllaBPKZ+tkskY+k3rJWexfMqD3g0Tw80GVxOu
FDuCLATZ899k/F8N7DyxeIRRAmaKHo9Oj1wsyAy4O7wirE/+WJj1zzGczN1fbizguQDZvwQrjy57
QKkOA2FU4bWCiz8lUgHrPp4daoFC2yTTuDzUDzLR9raTtgrdlO5bsBTwHB+qBYJXE/UlBOnZXJfi
h5qKJg99JjK91k/XvMw5QuMEEkT4cH0A1irDIPHBja0YAUB2ake5hKh7TBJq0ZK9BeqJteKnXa9U
4dtewgcaBwEMxZDFV5gHNCDtPypdJYFbMsk29Z0aJBAkhm7uBg/lrrSipKhxFA4UBeZlq/dLoVez
rRQAI0SphUR/6GT/ps3NG+u1MFUL8agaIaH/xF7p/jihN+/sk9S+huaeg7F6GoL/rKbF0g7hYKkG
XFiIWBcvaQMGrbNHZcPtVL9n4fGiNughfTz9vy7w+mQEy2h6zLDOM7UlxXwc3PF1Z5/oXkYMwNR6
S0mxOLjMjdBDgivW6gJMuXZImF5CIaq4epS4M0q4JRkn+nYr381jVqwnxkFR8eVd7e7XnemhdxhV
4tVsrfstCdsN8hVftfpiqfpzuQA2mw7E+FpedKMdTDZNHyb0QFQoHfGoUL60+5B/f4+nznry+ewK
Ch4IMrV4Qhwwe1obGDKuMTbr8d+GXcPBcfE1K9ndhFIUEyyZrBnW+NhtVBpS6OOjkUPVKgwCrv6h
SZcgZVYDQg0WAUrLfZjgfRnPrGKFuyNLxaLG75H9YX1XfqngEwUaJskjhaaxFCfpVYysgDoPaXnu
S17RQnF2Y4NnMzXcl02aWcujregCzxJz/x5szZQUHsSiOLmH/lsBFd2GziJ/tnuiHVd+35UB+6+1
mcdLmnO51fspHAtQUekYkm1cWtCDrUjiW/Ie8eHc+/XCObIugcSNj0NI4VywnlUMlP4gCp/hlq5z
tMUygzSQPNIuF9tmZpT7Xflo6aSLW0OUywtaPCT2zvgNuRJREHGKP0IXsV61PXhqTVpT0b0Bhu63
Adp+bLAwUE7tihjOdM+yKDG9Ya89pQJECLC9UFQB/h+YE1rPoIg0BKDj04iesWso7Nzy/ERF4pDl
YSkho8D025FG0reP53nGZ/hTO7X65MKr7YlNHn0UvufkwwZBYYp7dzQS+QlriJO12RG3Gl34w8rW
MYWP4cRThWTN1kRnPqWPukJjlPzCzOQrkIIjW5k6YSVGQtgx53+2SpJlFnANb2a+Qe+FIKA+RimY
2mZCZs8j+YBUO3cMCpFLq8GgiO7UsH+SLYOsLVrS5kGdvPdz8nwSBCsoy3z6on0YG975XJYdTo8C
T397huRpXUyeYsAbCsq0R6Cr2qERpGKB9o0X1681nmd8BHnHE1QjU/7q/oqWifB8pSoFgMRe0Mn4
RfVjxXxqBWlf3y2Q8THSq8QnzFV+iwnZyEsgHwECUSl61fXC9YDUzIdYXmbEX4tC8+IjhoJ9Y02o
X69GknCqVSwqsKpZwW1G9BYvil/YAAGww3X1ZYr1CjNyqFIlVcw3gI5qXSvQH2fue726JKyq9L/r
tOo48f6b5CEEIvKFwfZchm++QM+FWDC4X+2B8REG9HQxCo37o7DqQsH/usLUGPxGAW8p+uGIIfwM
zmomaRLKHSbPcZKAwBsamFgpCfzS1d7CcINRdJgQBWYl4VgS0SdXD/o4JFoiWIE9VDuBrDGpyHWg
VHeYT0w1zJ6trhs4BI10ZHfphz539WZI8lY5gVFbfnpP06M0kfm5j/hzoLsOdl3ANk4qvKPn6BCU
xblTbDl5kCbZ+unRQhoFGov1dXdZumZXp+Ej/a2uLKyGe/BoGIBoxaLYqzWoqcH8nErFyzfGVbA9
bHR9IIaApjkVAieRKC5EcVm9SI4+hxGXQjma05LCBoQAj2UfP/4TAII4rOnuh9jtaVdAp2SZPQxy
+dj79NZwLkntpewCaz1+/teVguKQCYHv02CJrbVlk6e8qlfz2ijPqoHZfYkHL8enDe3LUIboEF/W
YH+T9cPws02Vul+YyJGEDLajUS+0lvwODk8wixlCmq4azI5jw+SnkrhnBQ02ej8+cc2lz1VDMGu6
qMxUVcxi0Yw4qwHdlwvtcVyGrOAt9jiVuANQdSKp9OhBvz3FW3u+aKaNXeqNRUiS9BWU6OM+FQLb
5wqXf+M41nEzOuK9ZymmfeZZoqBSxHGRXXHr7mYwhgA06d6/VVU2Cg7SCfnbGJoAej+7oaqDa29Q
ldLLl89x5ZrIxJedatWlzu6PZT0tRq4MH5XV78m9e9WE5i0y2ynOuMGTjQjRZ033SkCmZ9rswpNw
JErn63KBwXYAl2EenNko8bvCEFeZAyrJZiycPXnYIt0rp1TFYa8qBla6Rg0L+cCO2LI3JNmlxKnP
j3YuCuhQecZzmKj24tF9+Z3Moptn1Mx/6nq/aPvrDvCxPqyoA+iP0eJ87HlkKxPzt765e2KK820i
9zznQBlQM07+PURw09zdxLcB+DATXjlGziad27xlvAjP5Eb+nf2gopeEK3hCgJSZglPcjO74V/6T
p71ilCSIvZifuJM3IO0HpyMJYaZHp2Jp6tOGARKjvQRAIng2wYP3lcq0NOU37y/tCCQof9Su/Wk1
B9GWp3cptWrdHnHRfZCFV8n8jUwDhLmx8WujbxCECDDWAdxdRO7/wxl/M8DhCROjBIGPf2R3WFs1
B7nCBFqVPqww4xkL2SLmh0TngCLEEYSokMqOWPhhC7sxQGFzGBhZY5OMqVn2m7ZW2YyKKzDOAaaJ
fUU4clE0sjIOkltZBmnmQpYVFpvYhyX0K5rEydC5EHNC4OiovXqq+gPwHYZjzy/orHye1vg/AOAz
FBGixtfu/LWy+f+4LP7zyahZOeyNwC/GyquiTH2fbjWMe4t+rWtKKf60wSyzpnFfZgZiTPx78Bra
5vMfXJkHJDJGSRW4xzLgTZ6b+ZhtcUhZ+bHaj17XCLDNtwRR+ue8owRJ0yzKkBIc93uGNBIoKe8g
Sl/jY1Sa9QaFw+haFt9i2AaHCX8jIysxcuA/waAPncol/qZodhueb7fUdH/rKuWfLAW12P1EXDEJ
ZpjidmiM940p6flLWjxOEmuAvqhnnBCQM0phjsofna356cFLK6RxYF6/q9gmHqscvu9FFxAj7j+l
XEcijYhd+UDLjfJCnQxnuwa8DJoEaM1CLaavsopziLPlyDR2ekqwfbWO1IfSWkgThWaAieLFVq4k
7Ry/w5D7oU8LwFrKop+YMAOBOwCpy6jkjZWJEtTwuEgYSa9gi8QR20B4665e9LCgt8ijX5pd3ON3
FGWW9qvuR8YfnPNGBai0Ls8xeYCsV6y/j/oAskvYOfy+KMEhptDWTZ8oMKEcgQWx4Mx1lgypvpG+
x3m9ZQQbHCD5vnhTRCKJr5unScQwH+vjMcfgsSG/wSVwVnaEINMUohS4pBiDl8BXLW714LE2dcIH
3Dp2S5ygtHDFyLU6Py17v1xbLuLaM7H8Xt3OeQXOf3Jyu6mHIRawekvXGH8WKFbfpx6v8xI2S8IW
KiIRg1rcVJVnQhAKQR8PP2VYBKSk4hJ87/aOmKS1waZyVGuiwi0bzcRM+kD5U80asOlL6Oooi0jY
7QyR1i/O3g6m5nXtRR6/LDwpb9dj+DbN5+PPEQq+UwDO+hxVKW53hPqD3z8cImA9zC7N2b9ZlZ1/
7es2S7YcPnBoqt1RFLmG3+nnompPItghWp7cJZEthGUnsbVOlfy6Hoj8GHOr1pj9LNC7LNBYRxFr
UE7CM5Bx0cZ0qEaSFbn2FnsgK2FkTsFcKIoEyNqZq9sk6PZAe1lMsyC9fOf7PyjO9HUPclG/zrFn
netqaYctVtaZYHDNAinctELlmNaid0gjUANuz/luHUNgs8bJpw54OvlEc1SV+3PEGbOI51trUBlB
uM0MqPfWiwFKHJUg+u5iYcZ1YS98KPqTdE/EXrakLcNi3Aqa6Ir29ktc99WhE2cJn93V97jtqD7i
JiwHsuz8D4ukx2ysmpZgILRaUOruMfgBm/lS5WDND1qsk7v+L06tQ8+sA+4k/uxD63Cz5j+7zThF
IOW2NDLJflpVhBpfvW8Wrup1Y6djsm+bqGn+Q1bdmDyRC/rdl8W0B09YGKyAKKSNFA8UbKv5b6c5
HU00ccJ6oR8Sq953m4mhu9o9XaMDugK+uIDqeei9V0h/PEVju7DjSyNETQX9yHShTGSTEd/4fYv5
BVycKiNhR0ndQ6Ip5TwqIagmEIJY8/8KQt4YB45PUFm9ily78bWWTMLlNDQIdYLzA5+kBMrqNlWX
xgjyWV6qBLHbkiHLG4g6n87GLn1niSXMAa/30usVIHUIY2ibAS8FWDdccJthS0z5vDrdnEgQfLDr
5iYOXs6TwoIj/VGMYIQdQJWoEnbSmX9StV0b0sNeUIyzroY030C8+G4YN3IiE6sgzY/l6lDOTZnG
wQHQ0L8zeTksSsMIs/ozuEue4xb/5BaGtM87l3TCAmDCGvYayOkS80r0MTAwpC16iRNVBfBzaxK6
NOiBl5PnH3ee7RLCD5AgIjhraKJP5oI0wcUSLbnldU21Z7pIFqb8hWbIvJPJlvMv3Lx3LxiDf7nd
UulEFYkYFsN3X6ks4qnZy9VjlbhtX0WqprwpzVMFbZVWxmFFeo0qKT2Lfsf0/66N7clrr1patl5L
PibWpao9KCvDwKg/mgBoZ2G9c8bTUCtjgp/Rt4ODjf/4snewyQ1V1NHmT0ej6XQW1P0V1WSZO6JG
CBGLxq2b2i4biDcLz4raer0foZQ2T8P23tRGO7bkG0RvU9VGzRa9tEUbHVd6iAHCwxNyqpAgytfm
6v+9lHjgECY+1fCxPZHdT0GQx+8ZkppRVdSP4ERJhgdH/A2/hqdnDdvPINmVPTj3G8jY0Gkmcxu1
mRFIEI/4kKm0zdpXAeyEhE63Nv3jd45VQ5Sw/TLerlg17a98Y5+wEesay3l7yGxDbmidioRDAemT
GdgtO1hz1Nsm33hT6d8IfCLTrxAWM/AS1CdFh1JHjG8nxcMVH3ZNIReiFeLonwAa1W4ikGk43Wk6
Y54avw5TrQXi1qTuHfoBTvIZ6EjbZFMEe56gBBLzBgHtu9JdYuhYexLIcjmVz96FYkA1Ai1KxVqE
sVjAKGhPpbUsah89PS0cN9UNlAzoV6OGlxgWsumDO8PIpWqQBsCDstMTHbPw9ko47b+t6wSFmQ2H
qpj3Ynowi/mOyZkezV31HKQ1/oITA5TALgK3DGDtuNl6pjXbwXotnz3CepDBxmpm0FqSITvxmDWD
B/ND6xtQGR3eppCORifVjAf/7xkife/nUudcDV7G6nzkxleyICJwX8NBI1BqxxmMArsb1HFAK7i9
kOR7jZ1FFw0HIwRnoFLVsRo5pf4r7nnKCGlE9BaJpeVrzRUTOwh0z13EDow/aSfUrFt3rFnHzB/L
lBKXC57ZzOZ2jzrbw2sbgAq19fza8I+Ou3q2sqPjKwbOE1rVflG9WGIC/jbe/7VPF0Y//M03n73d
2ce4DWGiLbVF3LhAOnCA3cBMkxgHbzNSf8Jg93tvnxu5f5FkLSIX8U74bQIzeP76H8WNEDCquOAK
+PxQtlz1JAW2VxEM7IylVa6ctalMshO+PMStaWV3Ly6SJq/8XOQeldP/juUOOtq1jfHHIKTbRDvR
r5Oy1i6xTGQ/yky9uzc/xQ75c+4eWVHGYIJwJJr84qx+mFBdoA/T6ksoIzgPKpU0mTWpCelj/zFM
Ynkg8lnn6s3++hVCk5YXeDwFfOfS3gOLTJZwax0dKi2baxeq6ie9ZguM1XA9FAYEYfbg9YJNvWwp
Dr0hpLCn5rjr9FLSJi5RbiTZs/c5G1YWuRVkEL5zokBWhJoYPWuqdpziViQNm3Kgv4l0BPlW2IFP
ui+8eOPSYIbUsCBmJUetQwmycSg9s6pAVSFSGMr4Fx0QS5Q51MQu+VC0HVfvrg5GxOSdVuwyc9ZO
m0j8idcWodo5wY8HfyV68C5W267igxs1hOvCr/bmJ3nPea/aZNU+SFE87dYNJFi/spAkvcjSUVGh
R4hTuKncwdKyCLbazU3uODSSG7nuhYG7r9rDinXp0vLW38JAQeSH8MjHqHTQl95wAo0QLIu3qkWC
ormoR9mIKLcCDs+lHF92TU8V5HEOW1d06XDlVMxZaGpBBzIcsVQVv/SmUJGGRmieAv7kUCyso0rK
Z7YJayrx+owMclyxep3TH4xmP8BfDTl0/WRwABd3n3pTXxViGM9S5Q1oo2jlZ8BT/5gXR26MtEeg
q+m0BBikf9jD+sOIHAtTkciYcWRiYbUILbs2ztOu9ZeCafBOCeASxdk0rcpxv+8pdWqLjAC3/Xox
tD5OtJoUWFggkcyIBTUIYCmfoePUVMYweTZ/Nz/3IfJxkOMoqV6diEUe3Ypqn6+SS0do/XjWKaSs
ngVIew7Vnbkv5X5HKpwxRl8qvwAEsAfwEljyJlzj48MxV2cWxO9u8Wl7HMlipYoeAPlS/RtrfQ0+
RF3WSc1qy/b5NG1H3nVT7ITxcwCPpiEX5Lj9lEQcss1SsQt/7qrcprWw5J/tfsU41TZWbYQKJbiU
Vuj6s4ltI8QkXAyte150U9mulbRSjCl/gS95mL0fIV6oxlvqH+697IfmQJv9ttLhL6tuX4cYYM4G
2MC3PtBgCih2Uu6Qbc9JS04VcjJPair8pCWhmNvcMmwcDzWeDmUxxfF62D2UdEEsxAwUw1qrt92L
bUei57BvpK69zxkL1TZQ6w7F8AIriWyZlpCVK3zfKa+zicdT5smZ5ZHuZOWmGVptQCHmhJuX+sl4
6nI0BDq2fS3clc7rcNWBih+h3mL4ZvuZLdja469dGZ7HQ5rvuoIk+PLwIOw+w3Nbh72zXhqpc0jx
PF2/ehdYWa8e9p0Don15UMd6uplLeZ4aHoFlL9p8Xjj+HPi5nfyZgIZYQS10RSj+HS1U9IIOmlCC
mUwAfNZwX6fVwNEKpEOjWump+NtFPIqZf9AMEMC1CygSynIHT1AUG+xHFMlDvytIXWBwgsVUTaU9
Jj7kuZvEZhGOMEcHj+nDTGrso1gFAMtAFI3O/PCztpyfYxYSufay7NPDfL7qNrfIzT70Mq9F3sGv
Di74mbvUmu9KlVFGXnp9tKG+i20tKDRqgm+s+BsvIDNdaXYoG7yDyttyzSCaFkuZQ8a8uZr9h+nF
nmSeO66GRb9AZ+Iy2DBNXo0pTy2qviSizZO94Ld638aX7VxXRRBAda2P+t5zAhuj4Z4ngwTJdyfV
mvdbU31LyMBSBp36tLUdClYW/xYUhJYAEYsAuzrtU4tG5LsPgC0vLebmPV1Tm6+g/HMU0i0Y4RVX
vAlu37RcH9i7/tT/Q20BLtvsaMDVWnjRYDY22HP0M3UrKPm0K5xKhyM+HBVPbYYt7gNgj27GhwNv
335fb43/gZqm9TapDoCOxXxiTnPVyzBsBl9efdwGdKbFDrgjj+M5mFJvlIVxb1x80RhDVn6xumqy
BceFDumFo+3Pqc0r2VgxiIPlDdx9MJ0fQ5TTSTgXY/tVC2FRkJsHQ99zFz8H1s9XcUweuojPQyr4
pBOOU8o1jR7lWRmlzCBFEeY8DrywZXdUoT/Cdb46ywRl3J6VdCe+Oxstl0NHBdfj5q7MV7Ln+3gS
lz4h2KkqRDR66AcFMaa6k7G+eJNfvrfXkrMfULRctjYI4ID8io+yQBzRgmeufqxNI9Yv60q+u/Ja
cgMjHCHHiP1osGgHcDLln9x0fbPH/yrJqoKAn+k0AdeVXuIF/0S8kR6lSEVndPEswByNNloiqwxC
n27rknkEbFVd0ucbVtnE6ReqRNqHZlN1lg19VzdLvM6BfCEvGZ9ICGRptWzmU9AEOyG0OcvDom6T
HRMcdyrVm5/TVVB0Iw8eSw66GkeiOFQzyyrhkNO9M4reCqHywS7UMI1HC8qVu8mTUbYu0pyei5Xh
3tEV25C7RPiui/CBU98NIGI0UQiEctO2naQC0Dt7IhK/rqLp1xIg/HoAo/0LIhYKeD7rAPiVbTIU
SktAVpTy4oZp/WMMPhuz9EJ5ngHpUBIfeBWAPLxkErDx3wk2DJOhL9x+no8zinbshBWbXNhBFrFK
GDVmNbMBstmXOI2jp43m7iyaXljVNVv6dBA2xi4L7vV6tGenCwne7tlQOyKz3r+e7JulaqSPdPA2
FP8D6Dit/78nc11QiT5b588UPj2e7aeTchyzMeH1kQnb4v913gW3QBuvPyVhUWif7md8dTEVhOxa
I9B7ETmmkGV1ojGbRU2xSSJjJq23YowXo7lq0wXZg2epclsSpBzKlCaacJd4nZGHZkkW74IhG9rp
7N/mp8jc7iipVySH6rNlZEjvqKuqz+43pj+JRD2qjOBR4nWDWr1iKaTqGRrXYlUxgytQaB4/31II
x2lskKEdjhn5FFfQBDvYIVx4PsmtzfnPihivhh1jVQc18/OLrbTUyMAF32c5E2uSFimygCyFH5gJ
4ysLFu5m0qZVUxGUX/VYN0Qsocme2yFwwxdl2s//fDi8oTv2Hop4FWgFFKc5Xi4lg6Q70a1KevO1
iy0EmxyMbCKSsFT4il6ow86vXht3pubhKM4MnJVED3cTPLjhzQV3/srCiObkTx2AQuLo848ls3tw
px1vksu1uuTbYnDqN8znkSe0cpPy3BC51nBJqHspZU7oxCK8fb6eX8dwwfMV5KTGNEHmve8sXwes
RXYCeEMbfX52/ZrUG+s1s2zA5VJGeS9rAx5zSmjWILrzcUTnEub2hibxQXbYiS3sk1sFVG6773nb
jfaU7pjqJQelKg1lP2zfwKjTOrdcdATtbjp33MuI/885jcuxkLU+tGH3aLuHhZviRUCWjFa5azUt
J3AJ2Uc7GhcdFR11Uc32kFCjOQ5bOeLiUT+KsIGGDO6cDBs/DeqtHpfeQW22fqBO8VE/s0n1MpRe
LBEfn4eNQoFp1Tn8axL70BrXt/6dEVJcPCioNeBelkvohA9Kh4qpDAu3C0SRxItSCTz6J5myl4+b
/rU5ZfFEuCLLIqXgtr45yzXPOrfZmgE3JSE5vKbhG87yb9RrwvgevYdIjGVXYVfdhJleMmLvH161
HD4PfmHSnSvrBynQes7JHpeBHyUWte0f+YGkZ3JE6xuYGRA3lPmbNrt7sEl8zuIX+QnWj9dYa4oZ
uHFcCNZH0tfXOn2316XwUGXeq+JYpGCgk3LcrQm0CLbHl9b8TpeU/63Lk1GbGJnSjH0zcK9DF3wO
0ANjTb/p3arXh+f5W6icZ6gNUP8R0QdBgz+7dCAHNVQVd5jja0aIg9B/ZrOxXisjgj3Jk47KCO2E
BjGVsblyBUnxoqyxNbyBJSGQxFewoYsOaL2i2ddxub00zP3yXjOR43HNRFm/DOQrFD4pmNmqgKr1
xuhJXq8/Tm6vbPBat21u7iVgJSCKsDeDL2L9dwRnfKYndGt2qIIZngKs0Mf/tfzTqhKU4Sb9/Sdz
FORKpT63/AS/tmmlbQktIBq7xgck7Q18n3nBGH/iIv6tdQ+ZcaWeHD3DnQIFx8y3+z/Xxkm/MZvZ
XpmC9OHDsZsCKGXUbuIaHz8fHYjDrnbiLofHcss7LDP7qj1/HNuWno9oZ6EEbTNnu4HZwJWKm5vv
xBpK/SmsOrq+JW3Xo8WcFTSlTDjvtlmcGt6ubvkGaWYVJtlSJZQ8jKR/4PIzIQU5JQi9+AOx6s83
DXSQZ5opkZ1dj/wfW0kiPbTxyWktovJXa9OUIUPh+HuIB+VU1yHhy8OF5rlHcalAHIOWbewDlA1A
zVnMrsCW0RRC3t+eunWVl+ACQv5VMgTBixUxQFrlvTyfeVO1iWg/TXLUlA43b76Vc7tJlQbRHrOq
n8kJd9EKQVooxPtwUwH978I1y8dAOhYUvXrKY/LvdO1Thd6aP6ok03KQTtpvZ6Nq+6YG0TH6ib4r
7r2odqB8wfoCsSlr3vRNmJupInLD7YRFPKCA2CGJbFv+p8JGDozobPj/TJChd1i599VxZwC/5PXd
SLQiJeLsdLlQZiWBi66rOtjhDRbTpa8mwVzBfo99Ohq5g/dD/2Z+16vo6I2gwHmmHwg34T/NMt1s
NxCe0QfLcHSfCOceu3eZPrxzgQTt/+AvRrsnRUtKRrfU7ruJ9rUCx3k2u8WSu8+m5FuYYiD4mdCk
zLOTjwNlOPXNEr1tei6r9hZZ4D3Mr7hr2IibNw18+xI58ioGFD9CaznFh9udZWgktB+0dMQUincP
dRt0VI4vk683Z+CLxlWIN4n398P62iI7VM9MzH0jUX2RBRrJcIbs3OyQOyOxBZkvgI7LWJXibLDz
h6oIryH9VY0fIjdiISDTVlK44nIBNIQVlIvG+uJySM+eqvTRY0k5mVUk0yzHl0YzyNOeL69ZzGCz
yxSvX5k0ZiHfkN6stuERDXkl8VKmzEpKIzf0hbI34SVilmzOuUiZ/Ee9PnbxMkdcD19KNXupQf+d
4jzyVlUh9SH9CFh3oY+nzU88N6Z/te93TfIOGnI57VzhF63FL6rpvcZt7J6OGWqXDuBfVRhLevl7
+2VgGcG3XDKwZqtFKL7BZ1MIghuxV4G3CkE52h9AHyzeoI1mxYKCwTPXtWObEWmdg2tFoSHiTf1i
QUgjOCiwOXHbo4VTuhDgH1eIU/AsjwCZ+AcKhZKkszm5tDkZdzrHEldX2lcAAe8O0SXGy8+NZ66i
KInStJreIFSfchB1yTjycZDTqecMmX20QYEk9pKYm0XC8BnOUvqcTgtiL5R6FqefiRDzFqzBnt76
daUOra5bf7UHSglYE6uAoypOLpm0xSFFTgxJFqflKMwVsYgCUsonrxzvcFRknEuBr7EVdXJsJgdn
zpl3xG6qF5Zdq/1VH1noxuu0B3MUkFQJNPeZpI9LZBvlYE7wMs08RIQyAKiVdETt/zK6CRaZwOVH
fx7RjUcqCRkO5XgihJwSm+1X2jmnk0ffYiW+PGp1u7d9bLsNaGZwzjKowfz3pjoHyu1POKqtExnh
wUsb3xF9OrmoYkI/2MOrRu8hlKx2T5geBctHtZXePszpTHJAMf6ZriYqie6RhGbeylFJXrzvHLAN
FCAofvh2H2EBKD4C/zJQA/EEJDUbYCIvJaJnaKmWZo6p9pNEvv/b97dkhIPfiYinVWs4yvj+BPcj
JN1EcpLQZBd8Vih0NHZKRaKNHqJexIKuChr/6QUatmZAMvroVP+x0VtHf+daL+9XyAxa8Cu2Sse8
BUkeKHHIRs91qnUdoBR2XI5iR5OCq4KjHlwlPXjpkmZkgmwNVGmtPlFQMW6rjTjlCUlqX6ofHoJ8
HtMN3MOvgpPEiPQkDvz2/SqBnuCNbUz1k9jpiJsgxSIsSarIuJECb7y9J85pMTM4AC9/tXKZt8KU
jI5idi0MPnUailhseVPGyZhER8HVT0Bp5XzYq8zSNwf/HMOspQw/sjMUAM/Lb1Re+nABakx3UdrW
mOg/IF+kNukKibsyI0EfTSzS3AlBeYbMokYQD/Gkq/t/No5ZUxwWIeHEphf2BPApTJ9GiF5cCHtj
pl4IhLW0PHUu8qeNq09jnygfHhj7EtULU6mAK5i7SanfL9X4XozZM+m8Lk7O3127/KTSBPLRw9by
ifhRN+1Bi9jg/fC8nrAEoMYUe3oMRo63QTJN5E+Y/9DNuxV+7YL/ie4iJhcdN8C/WMrf6IYhJ7Aa
x7PoFmWjZwg39p7KAJy6U0QGiOn4vwU991yJDAiUywM34bDhcL/OObQpxX4KRvqIwShj7ikVPd0M
D3iLcio7wUL7bs6qWzyuL9HclGee4DF8nKw8goYsg8W9v9zlB5Rd/v7sokEkCYVjt/lQkX8QtGc/
x9snFPr1cEupLOdtQtYg/quEQuP7PmyCO/1c5KMh8qhq0uHsQLTOEN5tgUwmkvDK7QOf8lYO8lxs
rtLeW/OqHuvpPQsDjOwIYep/u2RBRpGNRhPSYEqXNRZvcgVxxbA0Yx8zIMGDnWIB0YsFr3HmnvdA
ro3fJke27r61IONLi3tA0VkMJWCI8p8ykCxn5cv4cfM5oGLHfZLuijhLZayOyjicmL4jVr1yUB4G
xauwF0YCm29UPERu+KVMoXOgHhdJb2K+X87mBmtEIJPqztUzGrJjGqrsvLbcLV00FY35P6Kzknzp
1PKwAFcxHCd4R1EheE9l+UuTSCtczuA1ISYYVS9WwSwlWFPD7DiK6Gv2e/B/6395hhrsc0DNG4QU
VLqCNu2Odsy0LPQNDgbh5tIJmXQ+I0AO1TuMiiBXDEIopYWL41yKrucGZDjfhGbvEFg9869doTAq
Ljc0ovkEjT4X6uZ8ed+Cd04jtYL/9hCgMFEM9ZvxzAD8MjhNVLPeHpx0OULCOkGR0DGkJn52Nl3M
7wr/c+GxULXVC0yIGJF9n5PTl6XBi8bt87TUxvbjIPLJ1x2HWh9o8dO9tYLdCI8wYl/S9MLGbxOj
nVoPHe3AlszDb5mL1JEtk3/W35QSDSpcVfcTbK994xgKOkVIYFOgALKJHoQlUzXw+WUrL/CqG5c+
tldgmjijVhM8ecd3DjgQ3Ey6QCTIuoXOYzGM7H1BsfYDlqccqgw8ANo93LptqOsSRoxuIiW9dtm2
vzIrnjHD94xEdXTu4i0B7vkltI6pP0Wt235Uxc+vMYvPv1a8zHoATesp1TeeJ/VTTz7ms6UNiEMm
Ys2CpmYQ1gxmOqVL0VElc8VAjBAzbC+rDH4StFT69qVLGGgapxPoSaSLFDzTk7OXkr6c5nbG/4VF
UJHjxLfjKNozukOXrDtVS2SdM6NA5yW+sIzmG61L4xMU/6SX1CqIC+i5L1FV0a906y1ohXKUzCRS
4HK67+cN8sKmq1+VlQJZeKnRuyDDwYyIimN8EowAXttB8IPRsTQqcJ+niAjAHRcFmfW2Uu0hPa9Y
4syN9H1VKqIqmGJ7jnlYJuuzmogNkfE/+DzxmAv82621o3kGGIxoPxxFkumQ3T7PGdGR0WPKBqsM
fNQxa7opPRP9gdowyBhDFg2Er/VOFwf0PQZPO+vCIbcCHLL2ewCUqI7KBz54pP02ocvD9evNj8NY
WBscKFg6oCabvM0Kl1p3yCwAXSjbnRYNRKLWn4GmNy69+Dtbg+h5xgZppTGAAdIX21uHTZ+9h9dA
zLY9Fhr9XFba2hNj4THIicV8/jbgTbK4AneVjZT/2kFW6aT9pt2fj2iEJdf5mHFkSs1W2fJ53QeD
+iIzPhSxHEdtCzqJ5Bi1R/9/zVMqOupHVTxO6QUD/i6oV4Ic5stzUMlhXMTGSW+jBp6br5KTf6r3
SmQWx0Pz2F3CrAtXUIivVSGJYqR5dmj6GXw4cxkMhNmoiYTBiJTccN/uu2VpOXk6ueTtZaBU9mst
4/nIYp2wWERQPPGYkK+IEJ9nAsT86Xafc18Bg4ZFAizDG5dZGQnHG4pUVX/EPseW7kiCBraBNDMo
wAHXrU9vDu6mVfJoYll1D4y8TZnZNt+yXF2H9x/X1OkpqCAGvp9mpqVS5KFZCixo7y+ixLTgveRQ
2aTEKnCk0bmkK2qxlbYnqOEM6/X9SSoWnrHqZjY/0fhCw5krBnkZNrtMmSTQopKYAwn3Cz3YuI9U
t4yeW78Zb236gf/R7Th3vhs3t9zKaQmqqEO5120rTgoaFxZZNijo541Zq6XoeQFXnb5BGvC644j3
2mkuJNVC2Zx1Mm7U4VHhuNjx+11HGh9rSZopLOq5IwszAAqW44gGmbkwHG37/eyKQz64Y/91nXOP
CjQhxAmIFhyVSVIV4Dp5a9UCSbmJfq/RVp/JQfNTMZw9PsAtxIsBKti1a2+C9KrvMPbOcuRQQRJo
q3P3W3JxPZfnsSdLCfMLbdEJ7CB0qFk+Xpnxv9et0u0z1wlY2KOblryxYPESmZ+Czn9+mfurkJFI
Ouhhhhpgg6QV38Jy3GTD6HrHeNmBm9QmhBcW315Ede6RNfc/QnPhC72eXLznd/I8mfJJl73kfk9m
njL8ScC+dfselGXxU/Ha/E+b2M+qp2+qhUn431QkTDYrVsaOVeyEkOrdaBLj9WZnmgkjS7Mh1iS6
majgrVYJLu61gODDSgVg+O783rRUtvkIvl9br3Kddo3OZm/SMRCagcsogMGD6VDPlgQB1G9/iKvw
oEmqhWK7ay1/XgD/IZROKiIBKvHRuNznS6E4nylxIOFwOD5+auDVBSjQUfi16J2rnyokF3GZjTd4
6wOeA6Y4l8Zr3QFyywjLRGdZBUQ+64UhcTKVt+EvQjWZcitPtbRVvnx82sC+yT8h/jawY/RkNqbc
XYzgi1kJOzWe6QafS+JX21oYi5aHwuTR2PmUPEsOB2Y2GX975eKROzH6ag7op/PsfEXu28qRntDu
zgYDWT66a1CsETnTiqxYld9E7qf9AMmz7XWhB9BWgnEuct0aCCvBs4OGqrWQUJxGWyChBZK4kBoa
PeopjiAH2mtdVh6/s6ikSzSQOJwF422T4xQ97TLltAI0FB9k91KXaeIyXVYTih6iN17JxSmUsfz8
lRY3QBfHR+ovqj8acJ8wXAd8GyZ26vu5RE5mfwwAyrgpdAwR+qFc4uY6o0k9efqgxf4+wBs9qoec
/PG21ecI8OzM+YblzQo3mqmLpvkgOTppMTePcSqLQL6Och33QoCjZ23CTrxBJpe4vz/nZjkK0m3/
IXZy+CRLzxSVfk6LKqB9lpMjACI+jP2DaUewawZruUty2rdAAbgpZG27zIVFLZXEdo6cCBE6yLZW
FkfD0BaKYnD3UeYqLeaRe2knAuKT71M3caLZgk8MaMqODiTs/Ldl1fk39QHXyAv/HV2ks2Cj9nTR
x4hFLWS3cVSkd0JzVZTIBj6BZ0Ulurk00+eccp2q1pwhHq2mgnCUwac3lKc+RVIpnIdOhK1sb9by
gYlYY0mAJgGir0CsBp4nYpL70uzHFiGP+fRfyCn3FlwpdF72dSZHFXmkvxG9Og7872nqITR5MYsq
CS06eXK+JWb9MDzDbHlLhoNm7LBgprEd3jb8Hvcpk2JqlRrIC5/OpxJQbKVcRw62x/+p4DtTq5es
YWx5L0gGLnEWYoEzo0WcVRM1CCqvd8+qrRUBmMKbrmfrhmXOhman1/X38uMuP5kpUZyauJ/3/ixD
xSYz8XjMbZ/eazO12i2eK90hMQbUA7V9zR+q0Xgak+pObDZmDrEtWboX7+F1uOZBpPnmQutdcgh2
QwGSYi8iai1cu3PM/UxXqnA4fMNNmoW/E1PQZ4ogsmc4XkalPVbPdEmNgIRyitelF2G/yRtGcOvp
u7HVN1U1D4eHiJif7NiZeVM6rTmudAVun0rIzvR9UptMo26LLzvFvcvvl5a624WEzpoNwdEyxtAE
BXU7jKdRoMN4zJWe9fEMAsBrDECNmDh99+DXPZN+7QPw3exwdGTblw+7y0LloEmBxo15n8KLM30R
TJ+ubOtFmQFxL2ER4jGS0KsZa9d7Rcf9aMbCfAtAJdNeOSE/tyHQQcIThyH4dp+WgO0otuCmMZ/o
62wdWj0aXdVNIhnLSubE147pXtSImVAhoaix/GAwRDg9dsM2CjwjirbOgLkIh9dPBOJGd2D/EeLh
Lxa1E4ej7ocHs+/pGNt6mYsLr9Yi/c+kVkpWrit8lvYy7NySoZTcsF96Yb56IP4ULvqBKhVPS4dp
5d5N+XJo6A0iS+RCGLFIugJ8x3BQEF/dNZi6r7rBPqx9BcHd5nmZvqIewEggmWgmnveoNkIH6vUi
Gw5QdrCFOsNKYJaihYCrV3G7dhGMfs4jdJHAoje32hDMS8FCvUpHew0jnUzQrIk5aEzpXY3nqotC
DEhBw2jussTlwHYFg0uX+JNLB+ekrdw5JrkPOV47Lb7Pm3xY2vzT9m3tH/uw0s8F71VkNBko2RSV
VmXFMsN+oKMJyvDFqKJVCqyg9gxNDGGJRCUifmX3v/yDCGqUPgG3DikwIx+mjgxIktovv1TXxtiK
1neBVLaFcyWRjw45lScNyvmVZxHZC0y8gSlqS/hzprH7t3tQ9l0m7ee/3KOCeAdXIC3/Idii88JU
/5EXp0U5MHGAn4CdPP2UrMEt55YKmpPg31IhX4ZM4KM+xVwHrpc2kBYYBkjhys1FmOtRZ79x4CBA
3s/2f+ST57Cak1f8hKra2Vvs7OA3rmZCsSJupjTH0YeGa0BAwEBiHNc1MQpaz6SJ8WZOif+f4IHR
/u/llT0zaKlcgar6Ukz1gckiY/cX7ab70Fd6m0L7zOOp2g9RrvUjLLTLpsvea87L60RWz5V2Tq7O
Yyv9EcVbgBwnBL7l2fiO4vYGdgQENzTeCFxCh6S7qeVGAGEOrJd2xQ0W6ZvKoTWQT8yhXtTIiF3l
8Oi30AB6FsSUPwpXdWkyRxGfTcbOYcRAEuBfYoqV1Z+hiDwhxTxAz9gLbKf1VTgIAG4fA2zGDHgI
wBcXSv+lriI3mLkengIKVNFk/WgJPMMfslXT7jCptv8Ax6NMGnsJj2DiZcjSL177eXAW/43MgwkB
993Q2Iw+Abvh4lQP22bSMpOxcW3Gw8bk56E/2UbjcJYmL4IW3+WuIrGKFKdiWdHhu+z/Hz2MOMiZ
2Mhz5s6c/fFlktTp6MxO5DOE5fggq0UDgl6eHNVUaQNYWzXKebUpucwaQOjjmzIPKeyeRVLTM1xs
rIOm/hQMZBWx86kI2nYMUhiDaA40A8VihpWPuR9FAvONkCxD4ZUoWP2dnhNhvpiHmkiG+ourIW9u
bAPEo+iztp4UtB9+ad6Q7o17IjiS3Eni/y9FYvpH+2fWJrTZo67wyHIJUhKW3QXJdz+Mi04Ccyd3
KtTymJVqyh1CW+vBRCYbnLLTUpUio2IDhRnzdMm49G4PXBsKSqbnNEZB7NJh/HoKnATWjvNWhpjM
j0VkA8GrlecHMjc8wxa5A2NDZSm66RBZyi9hSy3ZGjQnEGaCp2cnYuDxzFzgVZDuqDUt86IzBgqb
R1OrIBR/QtghYXxUo74cq7W42T+50o+9WFmSw+txobxFvCM/chO8usOcBmExDSUgzGksutFSy5Km
3nN7agVbRW13MnukDYqBRbXX6D00Ebu1fze8guWwE5bZzRzpiprzo1KgQ3nlFTK4BuH7ubrkwk8H
FftGaikeBlRzjes7ejUeXewA5J2Cd1suuXtBA7uJ5IuZC01Ou1wtcfXUVHT1UgSSBLVVVTIUHj0o
IrXNuFeHetX5Y8WS6IahjcuhdYSOnDS2LjdK0kDJYzKj4X4tMCZs2UGmPHsGmEBEss2n46KM37fG
0jKdD9TI2ennf28A8ufbQB87QDIMfiNwzIBpaN9Q4IM7Q8KyyVPUkUctEtK4QvAqmC5HHttieK3e
mMdJfgBgm7blVd6W34VOKleJ9SjGSykQie1BsQdCivkSFJ7l+ikepbVefz97f4fR8C+IQs3Nhtvb
QJ/1HWCa8pGWB/8VrzU3OAuDSYEmDQUDLnCMCSMnCSisNMmAoxAgeA41yFFkl5MRuU77d6Z3qx/W
Z0u6jzAeZdMT225nB9bluPvGFo63gxuhX7OcPUYdqjlrlO+HsXgNFHkvhvd091o5n0BvZaalPckB
+z1Hak0TR+/WmIKH/4lrjoy+Tfl0pCy63NaGaYMvZFNWvr93kkkea3QV5sGT4Ps1Sv1wprJaxCmP
Xrk2wUx/zboJDaSk9frPhOIFv4ct0W742IApnC4ft1vtyw0eCG18+vn2YAwxE8i++TuV/9iUkPfC
ig3gHIGTLuyvSsJh6Zg7I1VmvaW4TbCTCER7KuI5PPWdxpWsfjxeKazktYiHO0r/atTLK6hUzj1b
4o3hYP6c+PS7luhu8qusqUwv4In5Yy7aGsEikLREBO7s9KNadNQz/pr9/iVdw/rK/jHiXKt5Vupj
adUy5zmE1EXWIZTpteF6zjwGiE+rRtDrjMdFJnkqX3EVv4aYcOv2l8Q/vuak1sq3mL2ejnCk5Yog
V3rwGH2tvcKoZuq1kasEKVcacDv2TlG7sHC6UqUz7ldMHcyakPmEIDkI7r5U5pjZs1fNrLvjl1i5
NlSDCBw/15thoEiqUgdMATaHQKlCAeU8gGXWl4YVxqIB4a3TkXeGuroH+xZCoSZIaJ5psr4oF4m9
uGoBhjHifsmfMkid0Bszg+rlAk8T3LB23K53VQsunfSGTjohPkXWATyxRzcHhFH3bzSnqXuwMexo
K+fHHx6+FCWHjpXSNxnnZ/gC76F8CGs9KuSVLhLzZ6nLkUXuF7kgbrDqFrvxpEvPgBQ0jmq5Vzch
xGTkAFz2Z7hzVs+vkjyZbG6nFshjsjxcHP9J96XwGOBkK4W36O+VemLLIUdYcCgE4crh/3Ng7GNm
Gfco5oAop1+ErLR2YNgXAWOp0EOY5VDx12Sydc80b1A1vmd1bIB6Uj/A6YZGQnMGyQkgQNSw9W83
Knr6AooQ9ak773u32Gx2+NI1s6hGxLVa9jFQlqrynERp+BVs1jP9jN5CtODhTP+tIPyxgXqxWb9r
Kla8to1j2VXNFJF5U2mzOzJL54ETvsUrGETo//kOVfrIlvIAiJQQwVasDQnp01fV89qJqSSdSgQT
G84HYOkghjPAaqBvo5/xaZvv++P3wb3JccZ7WXw3R/3/GAMolvTZca951D4ITTOQv+PrwiAmHqjR
2iccQ833LdA9p8kHFlSNCyMQtgHo7iMzE7VZpUZvWTKht8/bMrHTgRaHx4SuYWIwHH9+lA4P4qnq
seSBgdaMV+vPIRcysGYHW1KDK7lP6L0By1E8i1em+2BhuazsC9Y7zwnnoYzEfRp4lZfEqsEfyvLi
0BbZfF/78meJREdlso8BkLkh6A1A/E/ALgmXoiIcZ/8hs5Zi4zh5KgPzkvCzYjkEKBLjBeqiIzJZ
oWQ9qPBUI8remReXcVNnXli8B/YEwVwFdW/+l2+stII4/3I+ztZPKjOWj/GR8APXoi3GSP6L+wLO
HAcf9HDhy4B5Uw/uCUYeVHVtMdOsiJILuqXUgeLECRuC75UHCJn2yEd7jLc04YOg8QszxeX+wXpJ
GD2yyPob0uyB0vVCXMV6tKIj52AvV4LHj7dESA5JaRCU4UWMssGYzi1WAbxd0Tf39t/r6Umgr/Wj
E2RifKqrPKl3Hgoxqd4D8I7KYGClDcXBeJMVy+uGS5YcoC/Ci58ZYynm2vyBnsCoeoGxNLYEGUQD
D0r/cRvR7/pJuGg5pUcKVt5s5seqRcE2tbwb2exixkIMBNJislO+DiGxIYa+p9s+JlchcWJCNQaG
ngAr2GRZY0gU2c41Il1R+0mABoj0lxXu8YzR6EXLMRsviPuuyPT/muATNf/eeflsdL9APsBH22Vl
BM0k2jqY+uEcljs8bLk+p6g4YSmhdQzB9LzGtL9G9IJipr3l5fxRFzO13HAMz00ti8NtXaE6IQoL
P5TvWQxlCGIshXm1T/57EHRJ6esmF6qhikqd5DVUGJhUSiLgFZb+FTqzokL9qoQatWHmUPps3EYb
lQ6+x3KaS40L7pWPruZ9Jw74wUZjzLew0JyAc/6wJyuPKkNQo4xAnWohWbo1Y7xGLI6xEKxwbo75
qKCVvACUds6SRaBfnFvm0qPtSL4aUgdZ+kctIhVx4SMXv7wr9Uptr4LRjgDIgvv/cOtDQbeItobW
kPruBNqyNCqLN3ctqb+61oM7q/rabjocr9PxuYIniXsp14h554JsdjaiOLLmlBAreMNp+CITEy2K
69fH9Fuf/Vw9R8Lje9KhTGWCeDMxSU6t+uv2uo3i/HMt2OfBIkO4nUEhpqREidanNZbx8ylvKay4
lMqA1V6FlCFB8hLtCKI8DdHlTjDKORUZqIHBOFsF52psxNZnNVRAD4UWjXoCVVyy+tDvQdC2/vAY
wn5VhjGqCPW0YffpaJadvzVNi8VwmVDmPJ5P7KefhhyO9/WYHIvTj0396u2ACyoS3JT7vF7YLrFq
VQGH2ROHpusChW5O3VMNjx+LFkNp2dxokl3dTOO/9rli1TDTp1RY8nKaAT21miIP7I461abo3IpG
Yd/jcb6bt33DovrZu+1UGpCXpQtBcj1RARp5bvU+26o+I9bko3VuA24LGtlLyMAza6M9Dlvb9yXA
FNU0O/XdzS6+rOz2UWS9kUxdGH15IPCCsGEDzkw+LNPglLSu7PQGoGwf74nyQG1wrOLq+ZZhvKjK
rxQ5Gq8Akq9kujaUXLmKA1vWgvJ5hP5kZ2NibOJyGppCyULyduNK/YcDcyEMrgC0AICOq3iNr/jA
++7rQsPaZ8LShI6d7XDLBZ55XEFxq3CygsR2p0tefywoAQj7pMt44n8wrGWe0LEPxyOyeNP62HIf
dOQEbkfi56iBoIl3BdbnFhywPX+T6OiR+TbHPyW173zjtq3dS+OmNAFfBDHG+FjTq5/PLLzn1WOq
XnmD/A2um9o5opHyKx0VZw4PtABBlcDsixldRrgSyc5DEJPJ+dDo63c1dsNvDNqur5+xr67rfd8W
XKz/t2FUaMi+lt+1KZe+9DLiCeD+II7FXgfXqbvPgOimwlilUbbQ5TiGU/9C29OeIQINfTAy0Gr8
tm5ZnYIu4/fmLRE7Q1ibJuXlgHg5dZOiJoJbyYBbEmW8xRS+RrumEDoScDXJEgACuhIGF6Ggv6Zy
Tuwlc0GbhUWyl3JSMMvFOQ0uV5oDa4FcxV3J5HbUGxvfddQKnGAJrUaknhK5XsV7YnJrjA7vt275
TujmzuLmuVmamOMkZkRozXxQ0s45a1L2hYHIquXqVvyG9x2Mt/EvCkaCxOy6PlD7Azqhl+HzW6Dq
DtyZohGOY+D1oq9A3Yv2dzfCbVjVkqkAVdSqZZTLi0Ua9U48Rt0TIWzxyu2nQ3cC5nbJemI2J6Ic
j43akvva3v+Q/xoLD+bWxHZPiuTOo8UX7LpJGzeSaE2magM4BEy2tPU+2281Chl/yNm7U05l3fSS
cZ8l/bEL4ElZRP3sz4TGzC338gPFjg9exwsQAuNHFEftxFbwBKi5j0+Jc8BxgZnA8ClPzS5b6+D+
oivRNyHUsiBBPaK6EU7pNSjdsmEOV7tLx/0XOSSLg2CsZGrCbHOT76SoiyCOgoHYKbfHxDsRQLd4
DR1Wram2WuxZMq9mFubDfLAvDBZ3OJooIkgMTz4jODXxk7vrSF8xlgRLgXy6FXvyaBe/LPAzxiCK
cuf42jk1s074+a20wV9wX4iRaAahWn07VYIePHF3xl9TvxC1bhks8SDaTVpW1kPfXyc8XYkwyzDm
nY0h87lkZ4ASMXd1TT7cxAhT1WlZqAxg12XUPxjyb8y6qViGCGPsAdAuOPlrQZZsxn7s43coi9hv
dlqOSxSvtCM5W2RCqDqy594P3J63B+aJJVY/mQhltbAiYeYUZxCsf9IdHDWAtCm6L3frf+qsmIBn
upmsyYR0/FBuxUwgya4+W9SlXMOy8BG+LUe/N94tmSvfYpSdl56eJJmKGHeDCTM454fUQreBv53m
85xFxKhxacYVuoOk/NEs18bKRBcSc5vk2FnZqJUnIOmgVFezWkiNdVjvjEix56Ik9Z2egbLM2se/
k/c5g7D8PdyMHZuVwYvIjdtOG/YcWc9drv9DX/D7My6TTq1eAJPaF1Zngt4UwbZz3sgQSgzC/ZTk
pPdg8VbRgxbw+aZOSGOd3xQoDmDu4vJcf8JwKN43Lqo2bH05tVPPZy2/L5DONUw7FJ0BOpzl4ye7
41EUnvNzPIGlH97FDbE8laOceY9xsiAQWm/MQZyRLBgYJlPXiZsfp3r/jpzRpQoQkGeCCwYQCniE
dKAviyQ6UFuyU9rBjXUFIyGITqzI0oVMqGTUF4h2NGXyGq7Sn4cgxZSjDOSj7G6XOaCi+I8YyWi0
pJCOQNTGoh4/PfmflycZ5F2UU1o6hrHy4iRKO2R7X7vFHtHqGED56Uf0V1gQMwUQu2WotI8KkDWy
Qidz9WUumLRFHKgOqqcEsrSs8e5gom7mQyddDbsnYvjNB+BjWLrVD7kp7pVtdwFrvDt8/lzl6jho
2J4SV/fi6wNwZq5TPKJBxfC6rPgeJ+XfSX0UnuDdQBFk9YTcRCliIZFPXoULXGrHswWMKDb0yJ/n
quV5LY0Gie4YySva+hPKit+UN4Z2j2/xdBMQDiZggXEttElHF40IAvAym+7CbJRxkSkRzc4InPTK
RVJasPtB61vJcuZVWbogColKqeuAClZbCZjAuW27WTbDDz94Ezu6LUu7Z70hMiLv1Mt3i77vJcep
ZqdlMQ7Am/4tOPln9z9DPiYXqun4AT3+UbLdSEHhibY8EsHgtO1S9ak1YptsSYGZpnEPZkMbTSe8
05K5iv1SyTSfwTwNjCsSZpeHALSz9JKk8fkESnnNu7B5gH8H7C99s8kJx0VCYae1velGpz8hWCQr
vXkLoXxzi14KiDqeRePW4fQ2KpCb2QSEG0S73jJYKl+9xI5l3Dfib6mkEYo+w3HrYYJT/zKiJs15
OAGoYOjxhV8Woex4zecQAl+GluoA6qswIAp3hZxgbLzv3MQfNSczDly1jyRrEN+21BBTMju1adVe
oJbTRCu7IpIs4+FsgKxLyqDzNE1g51qAXZzhZQdSEquc5AiSchtYl+ad9es9fttGwZEc4LnKALab
wPFRTF8P+dUV6LRbFXTV1O+T01+Oh32PeRFavJZzoXvEgncJCDr9BYZDEf7hNz6s7hQYx4L4QqJq
6YgfJeORCQ21pwomhF7v1s3Y/zPeVAiNDERlmRSgpnitncan0FvOrSjPvGAQ2AIAQuZIG+3LWQOp
tv+QWGMzijebNh5wfASquQVpD+vJ9b/8+LNtGj77X3PigESksHS/Yj0+7GZHmfkqm/cZ57aUeQJ3
x0At43C8OUjVJVXLm0sE5TwMfbPvePhuGBXfalaIUJELHaG9Ku32ZTgVOfttSBX8I9Y6ha7uOlO9
Zd6B/hM3zaZ+os6OfEvTkdSyXVzi5zfcfofgyAUtFwITifRuWtCu2qIMN9unnPczKI6taP6rsYq2
6r8Qu4chb3kbCKrpnaZd/fOEAn6l6XhDwBaV4lAtVIsvomMqcFmM1cViy61IlydeoveCeaMmGEBE
du5iA2YSEcLufMVY7z7Qiaq+3Xp9GQwP/A8p3bs661VqJQCPAG3Zspsr92eNf5EZyBW+I2ZzsRbW
DTWA7OHzMIFtlWY0TngRotXxU+/Ln6kN05kaOzUPlHsQZLbErZDntNENBJSseCD+2pFbJYXSsIPS
oEOeLYTJ8oWpkOQ0iGAh/ncJhQa7+s2gDB9KmCJYLSJMt8r6O/flz5zEUYQmmYCjlJXXR6afERKT
Bas77xLACw1yExt3ZlgVHhJZRwaCnF3ktSSVtQW3bF5Ck0pyVngnT1hF14JLEmELwaU7lvObDzZF
nvWnCUbL+RtlpqDybrKv4MVYxItNRindQIy9BYbjJFrO21QT1IbfOAPN8Se3szpCtvN2MCylDvXZ
AwB91UE6TKo9RTRfbRo2XTZlOWal5EkLIH5+N+y/6DymhCY6/EeXe1fpaooQG/ZbMBxscNX7dUow
0/OuDxHhXV3j4ou303rae7NWpSDbjUSVOuDaPhJLrxSwX/YUdcgnpSJhvtyvsSAOwNQJatwX9bPw
8kobpgC77yvPI2sil/pCUu+DfK5SgPXJjaa7aVDgcsPkzKVXjrDfVu5A7zaPZ/9pTo/EjiPq6z72
/CfqdxCloknMe0E2Ucjc0IeoHmkgbOWcN/p/uT33Sw5xrCxwE3ACXiSE3qCEy2Xquhv/8ny9OYHZ
2JGNiaPDHzheV+Zi+DU9ZwxF7ydvV8bh7DahDL2cStfdbf/zmxpW3mmI6URv5hO0lVQeyVVVuvYB
m45PH/FCv4jwf/dynTKVPqApcTqxC/2Z9b+hdz5acEkTLOtydn18Qanki9tcgqmrJzCMCbCoOsB3
DNB5MIyAepdfbhR6V2HHc0heqyOjV1Na4gSH3/RDmxEQ1jJ6qyJ3J/QMmnwMDMxmmjRcOHUd1vRR
ShGnryQPKh0IdbAvVuDzSnZr2wBSs2jaRFAkdnA4tB8zrZ7iBuuMSUUg5Myg9S1ESvvnViLBTd0T
hAjpP89AOCDI5iVqIXWPWSuePVTQstrn09bA6C/age1roeYsv+IXxwsEz77Yne9tzwHxMHVivHFz
PnuCgAa9NPocq7Ooy9C8DvYm8FF9pRcHlKXVMOWUv+y1DAgzvklwiD8rSDRW3fTR8KDYo3iHSiyc
1uRsGl8aDkK/Q6Ij/KdEoforWv0pfp6pKJHg7if/H67UD9WO8AxlT6vqt/0HTMSd5/zbiPThoMzG
+CvsP5tVLc1YOfSPVlVhNVJwiUelrzyKYSrXt5is+KzePScqeDI3wmGgF6N5+xQpAIVkxoXjstfd
s+zWLns+AvOU0L8cfby6l2ND/LO/c0h7IgqBIhbQI0VoEb13JJqyhv9yNxfPwKNQ+bckYF8ms0VE
nFTL1D011f/AF9FpSmD434MwGlaTVZAnNYxUYFFhD8SgRg8y95n8/fZHsRz7qU97p4WFtKK38ptc
3GtKkgOLllwX+VWhUTCjvpR41TdSf7MBPFEm7/IXOa+w2zBUKpAUEMPKSVXi9frPVidFkQofMLzT
0+RuMIQiJ6i5amDX32kJp6vSwm1JpiR84wJrSMg53VXyt9Y+OGLO38OCzAn77oST1KWULWxC6fVg
DaH1HdTAwDRS4xCJfCghVF8EFqVGK8y66Hozap2Ajc2FXFMb1mv2Nkp6AKWLvIhRGeik8sJ/WBAk
EhX/FBRUs31iyQo1h1Vg4/wSJjs4IY6dRX4ksvl62r1X4pGCatl/3lQMFGnGPKQsBKJCNWUKyqrk
AiwmLqS9LyfQ5MglYB52SE+yFTMjfbajaG8ykyOBaDUun9y8EyOFqBs1eyu/pbjtcX8/Its7jqn4
9XneIUdjl4HyfcGzbYh+5pJ2o4tFEAMAR+evaIiTvzq4ztg6FiLyxzb9BfVPhqZdYtYD0bgV2PCl
0LIXkL6NEaNAIk6vi6PMu02AYlmLCmROJs7Dz4oKxZ1XOdd6SR5iPWLzGa7EPUr5/F7lRv65FlNr
clBA6UDEE05VA9jfWgcZD/dukAsRptjenqtSakDzYwtT02fQHCy53ppLo4r8hYwJG/JwZBgodbP0
b0ZvqMgRxfYI5MP4Q29DiUQ6AvcwSgcmtUVxPcSJGcMmP0b9n4UtF4xhKR0o7aea5bYgb+RpN1+B
YpHZUioShrVKNDXVKzT+RODA43BUn8IAubiIMKwbUKytjoDkbPpkWmOZz37laihamVHXqIVhNUs0
KMo6uctaTwP5c+D7/oEv5RCUYyUou6HlWMh3ZT7blGp405kSIPbcDOQFxfMnSTaseJuDwikUEJtL
J0a/NbNM1ka7/GTA+FlNEohfCIez57kf13FfHg1JRrUj44TW/i+9pcRGsXqYXOaD0VDRRsbhoscn
GXWjy/CPjDZAY6nMKgGQvxNilfLgkdh75ra5/KeobLOkQZUhPwmL8ejDDbq9vrS0vdCXvYvPs3+m
37F1KiWPI92IEPbMU7lD0VgkWimbt8xOmm7ckj8v8fYjG8QN2QDQuqXm/1OKLhEGATNSFkTY5rOE
zDGzrUGafLc9qqqzSlopkhOjD9aHE+zYKLavnPqe1TEu8VLChatpJQ6ec/cwIOKVg10BAQTeVU2Z
hMEWWVvEqlUvMwSVlI3zg8R6bOgeV3ve+MC4EU7XK5Kfus+bR2gxa8caKIPiUGicCLL3UkZ2p7e/
Ty2o6Mc1gbxxRsEhspGihuIqrNdfGi1RKyzB624ppdBz1jejuEG3LnzPr2hr4giFJjfwURQy9uP+
4mcpSgyRYDmf2cJXSIPzDZD0LxA77Y9YwzsfRnSVblfsGh1IEemvHByDCLGDS7FDmhL9I0J2wHNy
MkOS/ygusLnqIYnHH0stWNlT/yPnaQosAE+eB23Ao7lo6gJAyUMZJ5fh/WWC6Mfn2v5EAr5nvdbc
1RaszjsX2hVNcgr6n2Z+a42DpyUqkH139XC0DvYMhnGtVQOixUv1JKVw9lUcARW1Uyn/dDu/SjV9
DNLE3YGqxRRZ9qg6v5ExE9K4XfT4W+6LBQQROnqVi+BINZFMIP+EqfaapDQcseVXhxCf3MDfvlV8
0kaArIDCMehqe3lqKH7Xukh6lCNrXCyrxR2THBwcdyyuOr31JbS3DkE0lShOrMFQYFqT366GR/DB
1TlhEzP6vLAD2borudzYpYIw6ZCFrBqraZXrEhtTMlSFyn2+LAmuCvJo3k/igxq2jOTnSj+LkwWf
L9OD0hYe90qpbPLJKtxpOrbEKmGINhvAxQN37wlVQ4pWdWSdsvvpy6p4ctceq6f/mwXdvf2ppLfg
XREYqCU2rm4XDxYKq0sBBxPqzt7p/V4UHABG2kfzrKRJRFxjxTP+ry4FJIaHrGvj+MsxlZgwmYVL
yRiJTnwOAn40gnehiki0gHHz7GvBxLJCUonSB89FqjOdWn2G2nRX5q3bJAnuSEK9RsOoiofpPtrz
dlX7pzaP3V2EuGN3cgWorUfNdbP+ed3zDP0IEmxh4uehakG+/H9gAKGUg11rQdeB3OhONdQIdfmQ
yI9+itSruEe8LHj51kvWiu5Ov8k/XASZ+Q2tklQiO6VCuljluYifzEF57VMWp5EyQFqmfxen0zx8
qVNEnYGecLy9+OV4kKSdhmAy7UwQ6qWi2vsPEpgpgy5GH//oe9BheTzEgciQSmc/MkfSL8LeCqKZ
7QI6Bd8olddWJ81u+xrbi9N9P7M761zXoZFKuQPo3uuthXG6gs1bBst9agGAb4BmgzqtSLmhj2ut
yiE4CZ9zh3O8D0MzO6TyYDgxMbglmLc6xQETHH8PwvHHh3m3w8EhenqlC2LnSU+ba16cFOPKvM2W
1OpsOkGG8HIEH4F5nTtAJtM9VzW9rRmn7141fzayR+GF+zU7olg2wrj0ZFSLV9ZT3PtE92+hykUs
xFdmjOjSV+xZeEof6qcqr+q8daXKv9N5W8/DqE3+yW0VnnCSk4Y8EISWxOtilU4UW1yX+ULxCAzk
LYprnRUibum8gRpzM9dB/4xMolF/r+p0jXAIRHZogzM+EOnAsPOGgTpYRkkZbPz2QBh2Z3uxtpic
Y7W1iGIG+sm9ZCU6co2WdUpoKisPTGb5oc+K9iTVIE4FcudUKNC20fF44Bmh9rtSyoGVYC24gctA
smEuZm/lyQgdTaGH0vlzzrBCQSdltLyEW6KjBiEznnG+dQIeYN3/4yKfQES3dCHV82f1s4puhZsX
Pwkf20FKb+yLmTJkeqllGt5bsLdmH6wxRFCZL/bGyolA4/yxWFlIg0MsMEim9XtElSUWy6G9lddP
IQOGl7FWyka6zt69LrRPKwW5q/UId3IFSzwFHbs7DCTg4w2Lj3moXWUNP3vyfNoPfwpcL3V5woCu
T6T7qL0mbFvZVi7qGZ2jD7TbG3y+e3Fd2T5hn3ieCixI7hPjh4JOolmeGnRA+S/gHd3fwWLF8QZ8
jO3hPCgGAwmXYRSLmbtAZhGch9806zwR/NSLZBVdfiUg6cAGHZojhqwFSkZOh0u74qF7Z62hGPlL
pMVcpwBtVhBlGmnMp8GrvLxDIudt+tD1nNLibsKvWVoBMVEY6qI1PlS0Kdla9R7JAlD9cPlNYXRO
zNViuLs/N6jw30l44XutTWbQGINfYC4X/QaPHqYuCM/xPV2DhlsOqIEGET3R9md5WIbbIGV9AuTZ
3Rn3Akqs5HExaGTeEbxn/w+wmu3wmxqZ7uV4EYVlDInf3r5I2/dxgjbc4YaRTktkSEUh2a+cAneM
UliWe5OysQ2RmTVHJL1EcYS45ZRNLEu95lu70MHIX1SLvrprWpyIRJuq77RtHYZ4dZlHlhcscaMS
bbSEEbEieKPBEUUsn3+xkGvqtgvBQYkB9Q+MfNA105ETIi+JYuIv0mZQI8tIfMdB7MrUrSlF3REW
c2un0bX7kTfYLmsK9tcYAwbcCeF3CdSezAxeHoM2H28ilCNDqA8kUxttF5IAMxRjTVdSQ6rliszy
2PyEmiJZcuF/LYmb4fFlntQCvXNUvsTZYSzbI12Lgzsy+5FG4uLESi7hCgHDRLysvp03ik1eaVh3
rJrUfbXoV1SjcjTfD3ataXyVy1ic67OXdJnEFr9Dx7Xv/PwgywC6gt+nPkx6G2mU1BLd4pnEuEWg
qSdDpe8n3hb6Ul+LOjkphIG6Xpi2ZRtnswqaTN2KxrIxGcuulEdgszPAzmxbfaLrdKjqEcmvYIsQ
+t4p/i/GkXAcw9nwzx1K7IW9GhboMcs7g6T0Qwu50yrtP8CcPxTeN/2VDvHVeYa85QZTA3Lp6L/g
iN12pwndcyTsNvQUUC+Z1yVE/kmCNpMuczbyYV1eRHrwUrS4GTrb6um/5n6Azp4aV4ZVgOvFshiQ
pO3FtPc11OuF9pBECFJOwW+3Wpg2EpAqEOwaVNZ1U0yElNA0etTpPjXLA6xwtRKYQcJhrGvikBaR
iroMfuN9SmOCvlua7/Dt5N3ksqOsuU8WVV3PHEXIg99Amfg5gneTZ+22ll555ufZ1Y4r9QC7w7sE
MgddSJ0oKZlIVDxyDLB4r+8pOmhXTV8MYIvIS4ardTjtcjqtklIdqBLMm0zEG0u84cFh1RszSk8Y
XgyTACZ15grO+Ni+5jp5wmBCGNqiZGrLmjsaA0XoHgjgNNGdoNZ0YxXYcptVeESfHAAOavKzWJIJ
/GUa83wlHRaLL+9GMmhjGwd8Gee+GYRs96wSKUprcvptY3bzWaYuYNRxXEDp/ZJBjnPMo2gyAZzo
qPSWHidJlV/KYxTXG2N1vxZpHojC+hZ3fVqxcenFcqmHfhGzGT7olVXPNBqCQsYkbgIKbynLMU88
X3L5f52HkkSyEcnQY2/nfoPM6tu7FqQ2EfkhrrFKLioviAwxgYvE49f/vG5cMsAEoixMfkefdYU0
ZexuvrPU0YcMAQdErPHUEHLBxj2hv1Pz+6BXOYbME1agBFqJ/dK0IAJBjYtuk+wVXM0hUdJjN1K/
1nJnXJ7hdXVKVgvWFn/e+RMgyN1uGsKEgzdpQbL4Bl9eRwLWjHJsRoG9klxBdfCY8N4qejkSmp32
cMhj+kURqFpgWFNBHPCtAnveTdEtDzz/t4QJ3CYsk3vQz8ak/SiOgqtdzZXwxiffpuXUbxnva6V/
cuJYh1Q2+XhtDDOQc9FIodi5ofT1FCMMHZUA5rjG6CZZ3gKSKNFEkQTn4omM4OvSbR+9CkPWzFN9
OXFxwDAJ0x2j/YCrOqEsyn+dLVWOaToOwlMOOczomu5ZQMiFEhdBzB37+ANnDhKdcw5EyP424fCh
UgEkzt+sTVjvvj/VShHNeXJokq+IcIVsNDgquqs8JHuWj3TueCv6fzYKoJArhYkl/HMYmHblqs/D
m6SbsJV+f3EzBA7/VpJXwgR7rVvLmUK0rv8tuDaCCFFwZqaHbjc6zx5n3MiR6SqiPMxh4dWVZkbg
q/rZggmn3C4Ho2TBRSpeuu1mXcVQLkUNDUxsYYg0gmJkroWb9rO9zlri/zs//6Gz7+W0cy4q8CDw
VBvwgzBsS3MadZjYqo8ofaccMfLlJAwmnfCCwdGjzrQNEFk9TXnqfSrSt52PLIlRc7dqr9YVbQCu
4OTxbOSFzQHniC6aCis7aKRB6c10dqr9KI4uQ9NKnvIij/Pr5LbLg+y/9GvGM+Wvjb619eZNfUe/
NKaN5TEjUVpOmE0gxzeT9wZQw2ED9e7+5CyhmqxdzUnQkgbTB/NSuhWZ0oKKDZaONgRn2jKZ1QKq
Fad5rIsvGg9n20priTcz2yuuPGwuxXmIUjMp/+mceMs0YSePONBC9IP4YoMBVTtZT3UCZk8Qkz0n
2Ia15T6fKR10DVV3JS+bs8x3RQCzDmV6ffMmu8ohxZVxnjjanBFn1nryGLmIVhrapfc27aFl3E57
YAgv/d5oLGrMO9UI3NQV+3mIR442xaw0Ifl4kLdUkbNTcsfyMKnk/8dsRACUbZIW0F4LBlem6695
ulyqrCCks/T1Cb0QjlZF7m4LugYkT+S8k689oL6+A9ete/7tf5OwFNL9VdarhyGEDT5gz+BJQTmU
ECUswz2Z/NC4JDgiBVcHhqMInSppyVnIp5ZupD9ZjLdRxjKVu4cgpUlaEmyvVP133usMkfP2Y1G6
JHyhHdlKPfCVsEim0r2aAR0gTjk16icrN+p8sOPwB5CkFeSf5SQ+1hXaAiOh6SBUnkGXu6fS68Hp
GOAj5YMYJoeVEVKnLGYrtLBN/GMIZxmbeK/ytb50HnIqtjEGV259UqSDJtFbHDL9R4YwSvMtkoCt
RXSxNOsfTSg4lTzFjHosSLseQB4FBrUXQPwNz6HLhvvIgVq0tjBWrtKvhyB8cYYjcaizd/kNeyyx
mTrZiE8dtpEwBhty2P6FeJFhLZVCsHbqnp4CE7//CY85IqIIrY54nx7NCfDYr7PLkLoBtPdMXd9r
NYX2TgqD6GX/8NDWwVls8geqDbq8IRBi1YSgdMjP6D44fGCHISSyL8KmqJNfMVG8DfCRZJ8xFutf
kAvrOpG0J5b2w3qsJa/zZEEAdnLIIVBZ7DgBA7du0qG+IUpbdsOLkhRADJtp1Y01eSdiHDICLPvD
x2Sj3QNh8sByUNNhZYAnZA4jBUnixyOcqOTUWn5kH9Kcr/eUkAtGd9onb3vmOhIuzrAoumxekKrt
f4RCFxq5Q/iHEflpyNhQtZ/u9k/oqYrUxF0sFE4YGkcmhcAKNO6vu95PNZZfgDH2mbY21GkXoLMz
z6YdKIhUphmzgpSzXS4pzImmskbzaQjFXW18q1I7xtK70qxpaJ8mY2e4H1cAwWhEtKlkRQx09mrh
0JhoV9qTvhhJ8Y33w5grCQAifn2JaC9dzXVDw17fYPrnlUwFP1zfnFknXEI8MnQ9hfzpivmCAKyM
gIfZhbPiu9UcOZ8+lGZnEsl63rGjgmu81Zmt1Qgej/pvB2Vcvi8Mz4oHOdNFqYySD2BZFQGaF3cv
kOf36hJfsc/LX66vMlAzjqzymtIX1NZXGGDw9xoplh4QZZXuPlQBu0XyBicbeZAcsfhrpbac+uHb
GJsKaydJAHbudDgvk5eUXPd518A9E6pV6s/BjV8jHDjazwrvGv6KkXC5x0dGfa0olBPujoQ6ddpL
2OllXySZtz0ZENCC2iugCSWBgLpmptxuetH95xrwa3YFcMeJmJBOORqI9NAAIcYoBEcpM/HCuV1D
apvodKTGKfbjPR1YxsNrrlUpSUg/UayLC5Mg+cVdVcjk8iuAe737UsadeEtRw0WYs6tZ8qtRkval
+uOOAwxYBHbzleqx4lPm63YfsUL2lDd1Zxdgwtg1pMrgKSAoK7tIRI4NSuKNiB3Lzyvp6/PJZZz1
fG9n+zDobHGdQEqQWTsPIg9U9UHpFC2CO39n/6X977chinE1Cjj8eUWzYP5dBHDlV/iIGseSwTq8
s/fZUoXwZNmhSd7z4YXhdwmnGh6h3E+VMDAaFKUn9ov2Ycs7RKu40Bh4EI0JxtKwhEYlYY46Rwle
Rcn6X2dxV+XUDtIVCtoRRnL1KqYZME32aeb+6gRNNVF6ngCnR5hfAS3Z0oc6doXSQDJowa3OWFZQ
sr7H4dRKY81vOFVss1kpLvoh//2s7G3NG8AA84QsySl5wT+ApPdmi7ra4uc69nufta9LoUjhpaz+
E1toHfFUe8eoa2ZkruVy0d5CtLBkZWcRvRQiWeBt2mFHZKO9gwhW8z9yO7lr1EOIklrIma/M2BJj
VrFGdxd0KFkfMhzAkHIGoIn99ddWXVNhH0f/NZrcD6lC7+Ht8M13GsHqA2bC9bXzGrCPgaMQBoqp
ZTjyEOdt/9qVwzB2qmcAJOecllp9BPp+uLViF9khPAVC0La/pYbSCX9BGj64Z1hLPz9PeSTSD1/2
Eidihplo5/1ihmOnLrL0uOv4OyVB/gRhztzogqCcNcfZdqduU2Q4zCWyLgOfd/hdh9Db5kPfiogH
mlO0mJtvq4PqCiiR5jm1LctZdZAKiqcg4ya17ZFNUIkwCQjWmxkdZx+2Zcn+4DA5wIXdAt9Jpvn9
q7oemtnOmPpImfkv0BnGKZJ31QOEjYGKbEnx/jEdFNQQOLfreYi1zOmn8mNZY50+FfTvpf5bWk2o
whkLKlvEEX7fSI880sfM7aurJTMYxenIOBAd0HnD9Fzauk9jQcgJDUvOUUXZWT2UuA6ot9K97rPV
Iv2vMxTSRbUvJdw0mQtiQ533NMt6STDhMgSJb5UjKR3b9DCLahjMQ7ZjEjT2S27qQO/JwVr7/DQk
bOLdMpz9pmH76xnvpPUvekwbAnTenoiKLEPXKrQU87JBFsbGqqHYdzZirSpJO5XmJoQdbeoLdAoa
yCwPI9/97GUNXPmo41EItiA9XlZlgsD8uXGlyf8XxbJqv6zRK9u4avL0nULeepmvwL+kVEqWY+ne
/Dny/IqnSoRobp5eNnQRMIi2InzZPUxNUpMOKizqD7LVRlLtrG1VJJ+f+vPkvX4t+fQIzoFQb2ub
ZnBkUjr4v2SA1FFkQer3ZnVid+yggYaMLtVeKUgHAIzlFrZEh2nIKU1xyiVIoOqAvLD+TdAkoJEt
fjTB3HQBdvu8NnZ/GF7E73VSN2hk47mCE2k3u8wSIMU/oR2WNbJ+XGnqxWZKEc1kToKHbZaVql0g
INMi4f2JvjL1cSaeZ5I4ypd2uYMz5+xJ7EdeEZi1AkUY+Yw4upnb7pUO9+TC5z7qyM1GrwEEf2Tv
vmkjaDW4zov7q5CMWVz/clMzkGeSqOq3l55+Z0dfa85fFNThLPXxWikGCWUTbWgRRosK/lm266DD
U93h04eKTof3OAr50MAv/2DcZGE1Xgqn/9dPdmPPZH828Ok33c0aPp2b/NxE/JyzLHsWm4/yyGhQ
COyPvzvM4QyTef06mV0iEjLS7ZBLHt8vmzu6MpK1lOL4HnwATYs5/2YYjBhxkulmBNZMmqL+zGEk
+QYXEZkNZOr/jL1/D96ZiwHxmMVGlqvcP0SZ3Th+IH8yTcXQYw/4MVADKGFDvi1K2MRIRoBe4Jyt
W0UsFZ1z+kFWIQUM6eniqMW9iXnzyig/tv1CPeY4Vc38rhcWhumagE7xZpGCRbl5gFuQxlwz+XS6
YfNdI+rewlJfW4dfZpJTZbqizYZzsQ/exSu0yNi4IzkJpG8Mr3vWVfVZwpPqW63qua1ZwFIHR9AJ
NtEVKOkkFdLFJY3J9YRcbW99KTGu3oMbix9FXeKVAdjbZr3hUhOmSPXlRKfnXmC2Xm4+a5p/Wbof
Pvr+zTIi6JsEeoMGxhMKoAGrKOzOIYScYVTc6t9R9dUbrF23zWXSSiWRDS5P64GUBvHcs9SqCCYR
dVkGBR7Pv7Bn3zB0cklzQ6zGHCFzBVLO+/jISJOx11/PTpaMmene17oet1z36Y9neVIP6lOact6F
VWwJ0pp3+XlhFGDw8FBZ6y6QvyDsU6M4/K7Yk4SET67zSh4tJzCWfqAFeey4VLnHuvYzk8dLWOqU
EIGam8lBm/aOg8r4nrbp/aEvP/ykk+Soz+GQu4ZCXgz4Dn9wLhXEn6VmShp4uKP+qbK92R6dGZsu
1pTWonasD5V6KXYnErF+ScFr/xCbEAI3vUmKo09/iI8NAiuUphGDZWUyNtr3g+67R/1z0KUov4oY
hwZvx/jHdIoqjG7Cfkkyo7EbJBqIxwd6JwHND9mfU3vUIFK8DPub+v/p/hgTYzoo4+JidlfUB7Wk
lxMu+iDrp5T1M2mHl5ChPVPekazMKCHFjGkS1w230lzxejVhzeOSVsbm2nUVQOnV39vMpDyhxtRP
9ltR6iTTO3Sh/f6QA4BqogwmcHvGDksYfiACuoXJmfYufoNjBRrpTL8o+7ZQD5ahYjJJjeF8jIKo
TBlgKvczUIB+GjOE3qfAeOUjuIiwF7YcOuqem56tMOTLP4iRGgzwgTK8iliphA99UhZTK86eikND
5pWxtp7sEvpVZWhsO2vG61hHV9b3dfE67l+oB+9Ep1oGPbk0SvN5kqLM+5LLmsDnnIWyKjHZTnMB
kxtkz/0Mgz5PxJ2bFd3LoJpbqxV63TjIWvxuIIp8OLOQ26Oko2GH1rPOFNIKlstjNz5dtwlaszlo
yWPU14jm04dR11AwzHwGFLGfAv7BcYWro6hO1FmOv4ubCspqXnqwfKdcqaxIplC7Um2jP+JjgVy5
pwUbowCjkCpI5p4DaDBGr2taOIzEVey30tt1Ol36T27EiNxSk049/yyb5KflfIkRKBMXkp3j+KhB
3sjw5qxaRHlvHvRMEtEzE79YuES1jNDh2VWwutskK55FyfUU1EecBGnAIepg6RpWiKCfG6C2q0Bl
ZgPSvAiH/C6HySc3fDIaMg6AvWtj/qflk+p+jRhhwTrAlWw2Pj38djqH3Tqr6oDQVpXc9H8tfv82
WhAF5wqIJMTVFsZHPV42agAdkhedGWE0JT9DeCBq+BFWoSnT21s3WMIEogo1qkU4eyca8l+Hx3su
FXRh8CcbLjwx5GDjXS9a0RU0GHlLRtAnIv0UcsisjkbO/hQFtf89ilc9oBg/X2LdnxOAUm0F0YIS
4sxH/8HGqsOKytG3VKnQR66v7Jpyy01hsKXOBnHirj+TQ1W/CMxvSM4Z9vUhc3LdtwLwQCiNk8oE
CuXOFf78sETOxezSzLiUMYbCz3e0ufC7jm0OFnZihTNV19jggSnHBfwMtjleG69B5iiLgR4ERbX3
a/xEjlCiq9MNf0U02arX6qJy4CeAogRyIFoLs6IjmLw7g93JgXC15BL1FP814pan7c55bRlWFf1d
5AmJowFBo+huLigiZN1twQLO0/S8I4g0LPqB/Yrv0oAa6dlsfkOGYDqaWVJ9e2OImaHsZgsWKmZD
s5ofZDlME31q1cjjLlkRz2PbThpXhTXzWadv3lfbaL0CVt3W9W/C7Pvf18FJZ/HJflBXUl7HSfI5
2Zxs4V23FMCpsY+uB1+Rf23Q7CzyEqfQF8PNJTXVV/BrN/FnZHit1DFmNyVYrr3Mlus8kPOwlZJk
SSWH8OstHW9ORxSWRbblCQwado4gDi+mFRzY35RTQVBgt0tpJQuTWZ6DXz4Ez2RUHHkMPYgeYvgX
hxYnVSmMm/c1OcgqBa7dXbS2UO2lFYSOy7dF3DrcaRw4gpzFj5Ticri+pAZGWt6+ytZmNONWBTxG
wn1NCJKk21lKn9E/cAmUHQv+yHHOac5QJvhpeA8EByGfjjvgXCm1aqIlnaQHUflY0ZbVuw448mQJ
+H4ZEeadkwLgZYiWXY7012EJtQu9pLp34aeO/AkrZYS+m0t9YN7/+UtFRqT5VdNn3X5u7yTLVO1D
aJCU2AQQAhSryptgnz30NBtDuwgj2jYe7u682ZVxQrwgUqZvLJWyP6LlMr3ksZpp8542MWyvMDtA
lNQb8t8jIJY8Lt1WkoYhsOvPWCMlBfYGBeSyzQuj5yRVlfxsOqct3iEZvkZoEy71NU6CynS+h8Ul
dLsiK1KYT6/wpltequQ88roFJcAWzsxB4fPL8r4K9C7Z0gsfZ5BBrS8jlM0ZXBMouIuzXGywSu1N
9IQTsDxCcTD31h18f5bcx7LnhdDrYi3chr78DbVoF0poerZ0rcXqRY76/BOnlvxutP/tyXkrDAhW
gVAhqM5xxg40EbL402/VhqdWwkOAna4h8Nl/aZn5Yhd1g50hpquCqFY//b2oYpYk0wOh+xFZfok2
oeQV/8AM6DaYIsBiY42qUF/8Va72RfNez5jqNKuTPDpkzvk6t95voCDLNRmWS3uyBl6i7hcB3xxf
vwxoklvWZmbohJ6+5fErlX1Kq2wYGN50sHQ5P2P/gZzmOr0Bc567iqGGW1kPzEWwG8Z3baj+iDP9
NtfIJ2R1IZ5lyscl1QlXoKj+Cbm4lRemojL04GQ/35Sm1BJ1zRvBT9fHyclNyCSmmo/l35ifQyeP
ESIGuExDWfIGsO0DRdYJ7QTywxsFV+0wJJD8/NxB7ae4ocRQoTMZj1fBkSRqzJyHB17br1+nY4ua
Cl1VX8w4YIIqjv3BIiWXhm8/U55ehr97enp+STAZlrzKRe4+aeZHX75XJMh/3NtZ5DXWtKU9J4ns
NBylQz519uch4iLbRo6BiY6a6PxBGwiraaltjDADI+dG1+cjUDkl5zp5W2mxlLmTSiVjHdriAsnG
/mSUZdFIGcKS5/4yEQJ80uwqfS0uJqnII1vWtmugR6sTrYhoDutPQfgyn3zjDGefNFKBxxlWtS5Q
ASQFsDrQsTqK7gk7l3CfoDk82OpwY/4dLlqs74DKlHhERBeFhkU8pO90OToY2Esd3e2iryoCxy4L
08+KjoCnR83WAzEbeQEr+AIS0VTZnJO/55pfEB91U2ayvGLoS+jUUoDTD9FcPNhC5Wcn71pXThOx
hY+LTZwSx5zil4IMb9bC2tVN6GTj6TSj5z+K+Zvp4FlvFfWy6eiQCQIH3wUu9/VviT5EgESEaOik
PkSGArV9EFg7NNEc97PNjNc5Eo7TBISJpl5YiCZOewEQ7kDkNGCWtnsbJQaxoowYk8DA3LgtpJDo
1TD8Yo3bxLkWvvVRqIZJGyFUKHhRA32yjgdfFcLnWM2ERZbduQYTRgsKFuV16KmglzVWi11SowqK
u2tGfvvzkT6TaSSCmMuc6Xwfg7ZdnFUlPet9iwX6y5CvI92RWRShSf47x5zANvnlZlVeDOfJhQMj
jBXRXHg2UbmfEVZjYw0/MTHK9mdnr1/wKqzCEisD4Ke5HWpqNqsAHPNhs3eZ5K8QPBXKyl7rXtx9
+QYBrTSwOkmgZuKrRhSiLIliakydftS5h8C1bcCsVYAFidpSghTYA4/jbDiadq1JczC/OoqwrnP9
AJX1OzalfZLJQp/AOQrLxVld8lEMllhdPrmNjyDRhrRXRT4ui05HfdIIAEw51O9p622owPy0jd+S
RM8mlF2CBka373GPg+Ylm8QNo84w2ca9DttRSg8hTPI0ExcrJ4V2bWQHH8XY/YRsWC0c0Fa4zua2
tULVL7kR16d7r7Ob+iYN3BXD5vcLyrIYBaZIQYEfDeSOwDhUQ2Q3EAmv7bR+zMZBiW8XbnOB4QC4
Sy2u1F5dqSusTh/f8Cn5F6W7qEsAyUNZe+ANMJ6y3Ix6aiStCG8ejhAzlJzkbphFzXtP2wkckdfa
wrXsL41nyFLi9BKEr5lTqzbj8AfTDwhpBBN+eQfhNzuVl+yKiEHaiiX4oS38Q2x6nubKqckMMjWb
TUC6m8KjPxIbNtCzhqCY6FbiNO/Lz8sGJ6MtS30y1GBy55pE/irNu3HSBmXgnMqw+ZsL94ZaShf9
3qQajPg8nfEQdOVLUX/ObfNVlnvXhF0UJK/gUTJZWcW1V9b4NyOwwzKGL5fyO88OrGs4epMlSn4B
v33/a13BJ53vf41Cjx6vrPs+SvDuNVT0gaPJsazCxuMDRqP2WOOv/DCiTAdM7BX1GQWo7t1HQ9SR
QkGXeAJRAFJqoV8UD5zLVqusd+I9IQ6qYednf+F08LO37ex9/kiMGA7XAPsRr2hW5iteziG4qx+H
VOim/AdOgdTZhsQmn3cHP13cI8WkmM81VM1+a9XYUbXCmjc8N3Lgo1XapfILJud79qoaE0Npoj2r
qEBxkKB11KtqqsNSuy6t8Z4vD4z/3YcDiX0hPA3Px1abhHOGOr4aJ5xC6dGo++bebw/JcaF6mudO
FlWfA/Ik1wMaH4H1akHH+dUi1YGaVY84BDwN2OvhsNk2eeOmDmvaXY99HJkbe9x+aqqjeMS2UAYL
E0dLoKJrmFhjS1jzkOSd8U2eQqJvnfQRXcAUSmXghdS7cYbeAWrJUkWlPhBLazWAac/KtclHZIvo
jZurV6YFn2PotBcZvimN6Yq6HN++nMTQoKLEIqCSuvRAF/zGoj6Dr8ZUSuRJ/4i4o0M5VcPBiOEA
RorO2B2IxiELv/5YOzhZ37trFL8H9swcTbt4qRAxUnzYL+M4opKhAtBMGQH75HxGLMWaTkattyYo
RkMnu7Odq7DLhaREPQJCuWBD3jGApPynrcXKXDJW5hBB4hDQIVAMtUY/wHLJbLnDlaCUP591AfrW
4GcP+at8s95ohr3H8zy3AbWHq+n9XEwjghJqO+EGOq1+64kMNsQyU7aJ4HsFCKov54EX2xVZUX6d
BjRHitKrzOJwVkIhz0jytURA13vfIxKMrnXIz0oBAa0sL0hPefJw7sYGMi2417ThdRd5sVktEGsK
A3xKkq41xrLgSTSNjOmm1Y5JEVMZAYY+C8zL2XdHfxUrRX60i7Ov/+mj5AZiFai6JNubegz4phRK
Kj2qYsVXnNPgllPL1up1IwEwuzJsRFnVYa53YJbuhRQvtWYXwsSf2Bm503pkPgvXkehMMjRKoKln
Et/6EOmzCc7YGWpJe0x7NPVxTYANYtK+4gukTFJlKXNZj4f3NcYEkDgiTriWoHJFcEnVy02XvVys
R6XYUGG5XLotCVb5lMbdeCKT/icw+pqg6bZ6xBOMktY0pgHuB5EkP8aG75489FVsZxPKeo/CXByO
WMUvZcse63v2za4aNetHZBjSsQxi/eHBIr73d2sfLa7rYcOr+AQb8ef3zoIe+kv1knMtYD09nvOp
uHuyqo4PAz+dMtd9KavgWascvmL/ZutuGXWh8gXn5AgM9728KyVtniQxtiGwezwd70h+fgcIR8SB
wZu4QJ+dU5DAsqyCbLe4eb9FiXd0T0ZyA16S1f7qZ+LgLplnDARcmEjcCs9tLFDNxgJ78nBbT2pM
1Qi29lzYPFiajaA7WF3SN3EYQRqnQwdDgS0OjAv4mitTIxAgK1WWQRNEN83q+wieboJRbvoLQj/P
7DXOBgfa2i4fqMJ0mRgf5YlqCVv1Fkz07SaS+LDsSDXlcBlXcbghDBr+SlctE2Cwj65u/aEvgMxR
OWR8lnm4hGk/Qmj3kMF8VUnZJQPDsHFC6QK9n3fdQqmqSfFxwRlLVdva+Gtm/r6lP19SNCmOeKo8
iwmNaO4ks0kRuoy0C80S3tucIG0TjlDeIVoq3oqPZ6qgsWo3u3aPZkyNTLO71W6EL952yiEscg6N
Lii3jj6/0bTVtVdFxmBLGUqxQ8/AORj6M6esX49+yW2o+3103/JwtvhUAkTL7CbcZo4d/5zC6haS
T5xcSepcZlGNtw4GRMAyaPOvzSFsISsBs9YW0YWYyofy2u41ksuk72ucVmZbso6Hj0FslYRqHiaD
2Y1m7TtbhbQDQhS4o31j40o+ts0U4s8GF/3ntnyxkGtyHyFuwfvB+QfNQySv0RUAmcQhpRQ7BN6e
cXWRicvZYAhy+Ama6xHfo4HSuZmwd56BoiUs2SltRWqXZyCO1hujBrqJnKDtnSZKGUFxzWT7nlXH
n3QyG9QYksk4TbnlvtXaZ6q+qtiKZVcoUchU1ItQHy4oef7sjaZO6vCJVB94lwyx2K5O1WWr3GyC
ssqGOGi9u3jbaivcRlMxEZLrl1YCf7r/BpXRQiW5Qkj027t4Kg9lczzHQ3RpMp7kG4kPHexrZo8r
KPj7gygIxohKLtnjcimC75d/N+fwaW77iomZoHc7CIKsHwKI17Conx3u6br2lLBjzeeYE4QzOXoc
yLjuiJ87PUJchA0L0DHU1H2tXzYLZUYuV2AtLefvygYHh4i/uk+FHuGqEh/P1iKmlnFHPgjfjJyB
itH5cmke8W9YT+vHKteizG6sxse+n0gmdbuvBXMeXpIUANDCehCHlQHGEkGrQ2v1y6TfFUm7bzuZ
VDz+av5h3FDfreSBJvktRvGoWcrVSxSVeuNTjIwYDs3h9n5a7NG119SM6oG7uDgjaFS7asQGXeDG
VHZEoMR626yA68Zumw7R1puDJGhuMtuX5fzFpR/4Sj6vs285gi+chkQ6Izylkd7YDO5GcGjTCeoN
wUw7Tq0OWnTclpiPDiGo4JqP1hsDCLAL4hai78FD3hRG3WI2oulti4aAlKs3I9zuYIm9TkvEnhjA
3YyXrKZIIsZAJ13EcmtIKYEKpEdR2Vr13UF1FXO+zXdHKAFG0pf7CF5Y7yeIQxlJCJhIIIXKR9pq
8tvqRMNH9lcJPTscaRv8G2MqJYOel4a9Zn0471mk2lquab4ePf7rEgutguN3+1AjWPt6O9LBuKfg
gpqQUW0DxAuQ1kzEWQvsukj95EPf8DuRXqmetmpuvbV1/Y+jicu97YeRC/m+Q++ylRGa4fxO4oo6
DRvvsmMiRkjuTpCEVo59Dj9qQLxmYIZuM7K54oJTKhfSqTokHLhurt0v7VQOaJ52MFnlogKllcdv
qxm+MDX9TwrOjBjSp4cE+aEoEkltvbLd5pYseLNYrjeuiMW/aHzdGQ2KGAXcIdRflb4Ek83SfuQ8
N7G15W+Ws+aBcfPjkZHcOOB+1t1X0T1FvyOMq0nmiQjKCmdEXUglwwvkHxQoMlBHCuJ1kfg7iy4X
4hL7MLEbyzpWJbIha5lQUgXnp9vH33i9pW1AHyz7+qR8OZnP8aDabo++uoWZiF8ikNoJ7ImIXACc
W0WHiRRfkUzSbwcTThXHO/+tNRxjy7I+azKZGThAPukvo0lpep3gQHDu3JsFGa8c4C7K4c4FvEi4
iqa00JYm98QOcfITdl2GFCB7Y3ekqN80ilVSbDHMoXCEVzh+mc6Gl5BZnxA4ko63/J5IX+CbynP+
LJhmq3deNN4JUvYK3VsteM59lyr4gtYHDVhpd8bOvxTlCE5qRkFGmnaRiiWAxwFOtHf5Ju15S4Nn
GHFsmtb4zzsfmg7otL2uvSsT2jq/dAdOqVx07ydLgdyqmAN+xLAFRiaeLt40aXgsujLSfkR4F6Gr
XfbcRqolCMMUl5wyst43c10iFPmeDah+BntUo5Pt37WYXrJSu7MA9si434/IotIUBt5+oYIphu6n
Ca0PfAWILmSmLCUQZiIkobIDuD9zxaMbpXnsFKrntU4B7QjyqZi6SdfQvfsSFQuu81qiITLl8f7A
V9cRC3MUHM4Y4zg+xGL4JmbWLMC4QqZfDsUo6YVYGKGz5LR/I8gFucB2ONdCi21EC5fpL+ONGzbq
io9Ixjy92h9fUHuiPAsUeqnst+S+yfRyeDkfLSPa32XNjIJ2S+YiyApU5F3OJF3r/cHihavDfvmL
IqoS04ZyDYByPJmj+roEtkRZAF55YTRIK3s8tUIor3avzhquuoYiFb74uaTVmCicIrwLHak/d8qi
CzqR5laSVehF4di63K4Fs31Jxti/sSK70PawlDQIzT/QZqMFoDjrlANQ/VDOk5EHTYLf52fdem5q
jKiRzAmpIHeyAxqGAk8X+TDF5SFU+7YdY+GB73Z7cBF0IuhD3Mn7J3/jHPnzRXeh3nU2jqQEP9uQ
HAZw0cAfWKdhIK1WA0f1WnBnIqZUBwF+qQ3zQxwsk9hbN1h76RLJVm7tfDbrcOOJuN/t1S2xw0cO
TpBdlrKy4nAUCGSjPRxj7Xc400Ty5O5CNAp20v/VYQGtEODfZpoP5J73koC3di3+e6J22g3p474k
9Mi56sW8ZPXVJyZfZUKLq4AC25jSkl12/3rA9fEbuOoYSHXbswYFOpad+f4BCIpKoRevpTmAlLqH
qi4ctJBOMuEatTXkHiiAtcLo1mjxUmbErzn6XKS8pmd0/U/2SrSK3XnXgS4+BzhdOrVzOtClAu/j
brCzZJFe8gpHJ9UgOi12xkkQp4FbJMWIROq9p4CUNJH9H8TfinjVEyuNSAOVCUCANcJm34zDxNpe
YVAbPGTqrZch7UfVkVixXHq6LCoJIR3QrrwDBJBn/sMQtezGKvr7QjF2EHLugEXdYzL5gcNc/TQs
0ExiRVC3Rgz/FcEJuaS7EN2RxNsWzFhyLuEVHZZej43aBkbNLv/tdIyE8zbEj8uVn3K3G7+uNW7R
V+8GLCynnScrgmsUejrzSBtwigD8GIrynlSApxEkkfjJ7OddmyCLfMRbZL4lXI2mP0v2c5xX/LmX
d5bGAA+yuJk7o9qYmLl/1T39aTVK3GMS2pAeACt6lBBWNT2Lkws2QEnqW0iXrt+FfoAA940I0mXp
TCOK4+hU79tNVANDQ4RCq3DUWj+gDJzZ3x1ko7sc6RfZquAScUycRNzVTWqiAg3CYTK4EaDro8Si
Uhb1HA8rxOA3y6k9QgSwwPvrfCKGGnD6BNcIoSHsk6hKB4ujt0cQ6onhjBI/Z1EHj50J+xmVsR7x
z7nKin9mbNxLsqKllMLv6W5O0VRk6xSrBQRMcJ41ytDn2+/G9OfnjUK/drOYQqyJ/QSYgUfBD1M9
kK1Etynk/EqjBbMUNpd5jKIgxNSTyGWDaUkgpS4ApzHlwBBkcB7VvMxiGRn6qhJfiu3Moa2lCtKf
MxeC1CYmdTs6TLQzePjrtCSF4xqbA5DTO7pJ1SS12sScKG4KIiBmPZdgZmW9J2Z1VE2/joHU8k3j
OOjvwIjWm1k50f/WSWJK12R5R3pXAuWAeawXR69L1b81ISt2UKsYCgbRQeo95EHKniDfMVJilh7P
+hu199iA3JdTW//QUM/uua5cAVjCQyuO1J8OFn0/hyNY3Dzlh0brA31svpRgGfvMLrTwyBb5GQv5
2fQEURiYxeTKsY6iWOV+C4fZNXvgUGbAd8ZdCqRB4VTIva3EvB5pvKeW85N3FQVBrxwi3OGjfrBr
g3Gz30QmI0GKV/wS/B4MEL0rHi7CDeQor8yw6bUzMd7H8ZgJHENzn+Gak/p2ChtCv3ztsa4Z4XAQ
paSfvRNBDg8DGN2yoGGiOfrOI5JnL77Y8vOjsVSOVt395RTOPjJHNZKuKi0XcBabqqBOPCNPPiAB
ZYX0cUirCt3gGhy73SZpFpjIq17g5QHqqsfeRDSh/F4q6MPea6M2rN9+VfdMJH/sTUCOSdExoUpR
/RWgp1H7XGey10819PL4DpN880IeF4rbR/qt3IU7A1DCxsG/oJMjJWG1iLCOdj7wAQxiE2hF+blT
X9H8GYsJ2J1HtaSX8B+oGP+rP2cn/eSPhpZwcfH0wWYVQO2irb/kfp11mw8GuekfLTBfwixTUycZ
L411dZRyF1o5YLY2EI3WHn2yvi7B9m6MPETCfoS78ignIlVTgKVUqMTEomD1Slh2HyG1+WqXWELu
9Bo6YMsmEJMpTciVv2m+EXKSHSizW9YavLD7UxwzAtGF4HSZCN9g4/+KOC774+qxuF0lzGqTmMLY
vV30uJcpnHlijIKiEb5r534psDOqDTSNwMjLfPvbxkG8wrFRnMVZ1nL1EnVu0fEnF5ClzsW/bwTa
fohBTYe1FJGF93XIPqNrDV/YfUKJoGvNuL8krSaavlQKUg2e6Uwby5JkOaSlY2ObmZWxwC+ShXY3
fDB7Tzctq0sjozByPe8a2Dgz+GNNl3n7YaskLcIyTkVfv44MNBIPm18Ly9pBF9fF1UfDzQxS9GE0
nGoWOfhhU1Zn0hzshuesJq2YjWaK3k3O4dos84RQ5/YVlNrWjrXR4dnIYhf2EMG45bLgx+o/8MG0
kXxUlu1sflyjv24sls9jJprHC+he5K9OjUSz2Aees0zFAfrxx8xg0N3dg8geia892QkNfwz8TdKt
yp7CV2LeUhniv1N59iEVdKtHUUsu44Z195ZwZhrHQ17ODV+I4waEYlIpTxf8bpqGBk5cY5LYPEO7
lo4Q8YXzQjjF9yUJdI0P3wxIVMK+SJ27BQ/mLQQA0o9gshyE8La8Le7v0a35X/2rWGZ8lp7SiVpE
LFeIuncNzQAbccJbG1/zzFQaYt2YTA59RR2voRl5ICgojbsILGWqLTwULDYyMdPaRXfUY9Vfawqm
+HTnUn+57fgOFJDoegAfdltZRZdt5MK0lz1L+tIqoRGhZ7jBp5RWji3DK+Ky1Sk/u013QCdwvyNC
3pPlKpljsjEl/XQBXEL0cwuQ/7Ynq85pieysJhk6RxZ1LJHan2M7j9sMuBDW9nX3qBWq6TaBzwoQ
CktB0JlOLYPzWxsmXg4mn7Otm9qnpYb8sshcp9lT0vXeVFYUV9Q7g0sum4h3HoWzqIqAO88Z3d3w
k4uHIauVX8KuJbeERbsL4XpQIgkJoEDyZLFXavWIngXjgVBrkHPOVrqJcoFJRIzkSgdqNG3YgvZc
EEPc3ZCXxb4Y9ipjVUEK+E2gPfAKZYgDSoO4F/J6Cvx2x1DFG01V1kNEG3d8lgdMdwAWKVzYL70Z
vsMcj1QBDUXSckaIrymbPD2NeYhQe50nxYuQCn9h39WfkesPtpcTYpiskvyoNLJ2mGiyxSm9pHMe
zrNYiiJy/Ta2bRmWKRxWvy2Y5kCd2HclaopUxBHV5TTH7I2EFGvuRopBZGekCMK2TagXjfCbuIr+
lb4s4+reEbssUVkPdNL+Pj/fDGOGMy2nJeJQfAsFMXQ20n/4A5ZphHfxvaWh9l4u+WvJ5/aJYZQZ
chpp84Iz5KDO6nDvVa5KRLD2qHYkSi+WqTZ0c4Y5zoHeD/YqlUxktkCUyfU+giWspyg3AJexzVlF
wGrQDr9Hiaqsc1WAz+00Cby3g1X5CUuQMCJiotFl9gh564Lh1kQQyc5rBRn7f68Of2V89+tK6uga
ccmOqpNYAY84oE1UhfrxwI1gAO3ELHR7UT6M3s7BuS19R2gnfbRR4tlSwUuZfRFPHhHFDF3NnCnW
6oqKjlM0N7x8fNiR9+0AADKB337vvxztA1MvChU6hQTOBQGIKhmURfjkfN9DzMgmRPum+3v1FBzd
5FXlQCzjYz9tKXrF689R+PTug6yDtdQb3j6DLcYxmv5cKmH6uyPj9sgneFJza9iHTaXFpPGbJ8Ok
llkOoXnFmnOzpPocWzdOgkp3v7TOucX/C3pCwcImcw3J4sjhvlux+GYVtSjbtf3kGld58S8etE1o
OR1fSnCLwVND5IrS82bIHlsrrXV6bvWctsICR0e+6fQ4zp1FjeHWlnhl/q+WzQ0ejx1aCjOJGn3x
DrQlBJTDVn9/XbLQ/SM00eg+hM1WzQiEOkNAWuzrkDojevmtP69YbrFdQeqb2aEWVukqhx4lLZBx
ZccUBLUG5HbiH8lmwHY5uP1FTZZNDvNMHulOhMN4Unlv2XB9kHl5bbzNmJrpINzsc+h829fLDBI7
2X+tuRzi0dDfAyhE92I0NhxkkykZBX3haeHuyEgetWRP88AtoGOS+uz7veRO9ACjHBpq2RtcS287
5X0sXfcbwmU5QJMJBPwh7DGuOYhJro3fClffwxffsXR8EsJZ/qbcXYSKB3b/X8XYFwSwZE+ogBs7
q2Z4rRdycajDlF2+edYbc8aPjFEgpy5UlPxrej6Z5QWDulFlb5aHbDfTz6t8h1HoOMWZpx2GcOBw
1NQdxjsGmjaC865QNSXjyjLQqJ826RGkXTXQd2BL8UjbegIREa6ki7vl/BS8PZVE7v86rGQO+2UO
XSolMCWFTxHSNC7ZM0Vd+G5NJE1vUSGhVKHp3VFALvI7BaVgJtXhfPuNyHKyDUfqdrusmd+Qxym/
pr3esLRQjC8SBtO5fnpbSD9e9CA+sFXahySaLdGyBC2scLxxU8DIiCXwPAIsXC2JecV8VekzwuyA
wSXrpnLx/mshel7EOjiOtvexGfN4vD6WKxuULIipngeVBOCNMSe6pbeVlP/GSZ+J6VQpLhPptS5e
rjnLnAA/0zxGtHhe6gw5LKnxK0FOq5DH7ACvdtxRYL++p7UrMVPol8RBxxymL2dCQN+1mBYdqcuU
CocYv5PIcDVQRlwWvr5roS2NiKw9Fhka/j1eW1AKvx9I/8tFzTgeY21Cp3njvRzQZushBx5TCGgJ
+CGKA8vm8WTf+xS6dcmiJI0mQ2/22R3mC7DidgUsXCmgp4S/wTQiUb+od0Uj7PDVgopxm1Xudb8f
qDz5L2PbT6LNvzBBvUyL0iPjjm4SJL1FmlGSnXzqrTW6zQorw57QLxp/oOZdhEdb21HVgBwYOSXT
DpdFp/0Cf4HEcUiZ6qvuM+BIbK58XkfBMMHlKKiznsaHYgSjwJLVBLS0368+k3RsKIz7WDUlk7r6
fMEXa6/ArtFPShzNADvNFvv12SP/HblNt5PS7SGXCVFggKdSIABxhorHTAdQbvFArQ9CGNAToDbN
a+ZjOWA3O/HUctkkpT8zNnPN/LWvQGd02cnDgZN2PIeXi12ycP7svdlu6N8GF0gbsUYZ4gqNVRGo
9zxY2b0/7w8HeKWv7NPl4pB6S7W7Cx2vc2J/gXubgeooYsPbZIsxlapFkueM8NJpFr9uVyapksyx
UuKPRw4wNdpwyWdO0JhcejatjfKOLHFYqxc4iObzkgu/sVgvjT3eE5wVtoDnBRoKww/YDL46aTco
XEBOjkILnsawEtyTs/HKfsNooQvrfZy8PaphV2oLn1hVWU+6zEWD9sSlf5Ou3Pf/Zbj2d0M+HASm
/rAOXaWmAHHcEsbVSqX1icRVCTNrkXHv00qkxLdcE4z52W9SHUudYRUr3zZeb/d4ylsfGoXY2VKO
8u+ArfdBQYrGxqbkeE+ZAnR9RHKh3pABzNC81D5Ay+87OaY2bBADqN+le9PbKnXinmm5eAk4hVqB
rpJbVbIrHj9Iw3ALrRBJqS4amVhSEDtrhFOMmMqf23163Ocr5o1FwQ5gcWCJv5fwVbioksB5/dNh
8vhQiG59CRB7kw6MvYIF8D+Zz+jv8K6JcZRVNtdjEW8M3GO7h4at3Jlej7uC7s0d7oGb+Pzr+i9j
LfkOdsiZmGXHRliyGrr0cSd9YgzYxcZHebFeqpm8cw84hf+bSBeVtS5wsJMPDkTHyHcWZpmDqYuC
u35ALY89mcx6GYkArOArT7GfKh+JHMbsPc3OuprvCmA3nXOcATZl6m8jdQ2sXKZ3YzbDw8NMu6iY
3xiskVhWOjMMjdPxZPeYbqXsbaAJqLp57DbNxJbFMG43wEY6rvSXiGPBBhVjcpe1ZQU36LAmTNzG
jJCaIxW84e6rr2Qng+7WJ0tWPzvf5ldtX3NSQ14MFQooiWP4TllL+AT8YhY/5eV4OpGpf2DsJExB
IvAOb1nsmuU9LuDL7zAnqJmGhwEBaAYa++fNgAcBkTAColQPagU5mOHwlibZWPx/1+JA94J6b/yd
/KBle7YErUG9xMOz7pJ6fXUyiQwoZligmcRFEkegMrSBbYZrtP/FdGXnRAp7xJn5BHmFjfs2HGPA
cMmj+sa8813tDxyuS0CqLsdoM+3NaSRkv4Jy6NAq7m/cSjFQp7nHcbI+P67Z7UTP+ZtGcIfoen7z
ZZabIXMlEwCtJV/3vyYppuCmdYAPDmLPY77m8Htrq13ZNL3QNM3LJhKl8eG6V3gS28MGKHR5F8jY
BYGpzQIc3sUUDMYo05YLPZ7JBBGzIb2CxISrKXWtDp2gOMSTemnT3m3Xon+feAlKh551/Na42jHR
RJKgT5KLjVMJhTEhqaNdaUeUNiFYCxxqNqljBZDglmXmfs39LqGdz1s450g1oK4kuHP8nPwBhaZh
0iyuoiOxu9Y63qvi+gLohKFYh4L46O1wUhSOCXgUmGvq5Lx5lTV78H3lpqYYCyL8ISORF6FWkJMJ
oGxrSun3XInz94Z2CvrVKx68tu4utsZi1mUKW0dMx8FTvOlnh78A04AAbb8jvVfHmN7VG/vrDzfG
xf5BpavR5uvPwyXpx6hcE9INGOpPRdcuINHY1DLLH+XvmV1uuTJtGY1+nAEuvwhB1MtCIlG0KI/p
gLMV1p/mbgUZFF7+rCjX2E4byACLNZ9mkiZIl34BymVjLQRIkWhblQ3txATGp9fIdUFPCDjBq8FM
FHU4n1IYyFw9Zl+368WJyc/V06LZribpljWQu2WqwVRaW40eQModScFOw36M/pg/Fe5Wf0G0m6i/
mKhwLGmL8FjdlncZ692ZToIK4r788XscZ5PydzINaY4fsE3mZiiGWpSTrbkNBKPTYOUCz+C4yqqK
LsODm1w/MMXjib/7NuHM2fz/h30Dl6JZTElXdM6Dl5F/PNef7ECgk9DSZbIJq1aJwWuEUANi3KiG
GkoIzm7wVKtjOFUJ84tH9bsMTEwKyyODp4/tsFFzFBFkWyL2eo7KuI7N0WAGqIfSqERhwRMcso2U
447JRvS2l185Ixd2fwpKFtjS2bJW6qoQk4qf733ncibZRlqh3GaNAReaJvsCAko805KQgp9p+YHb
SFCDqB7rX39ajMsD5xBy7App57YqVjqD/Sp4WfjDqRRJbflz1mgUBZ/C0D9QzWTTu4ItK6YxwSxs
eH5JFPceXi6Lz2aEz6DqzDkO0EVpRvlK7K8trpowE2OSiWwR4WwH5BIDQ8B9IkWSIUCG6EUwFxp9
AX8rAs8b7m4lKcLeRcizAXsfJNSJgof30C4OI1ku3EXtL26ssVp4I6bygbJSqV5M1mCdQVHTiVG3
o0eY5Cy1jyBA1iCgQNAixuyIuNVfK632qhTRWrJTeiQkKG57g2OnhEpDxxhwMeqBFtZTLoOVzEgV
kWRmqLXm7IiUqcc+jwqaIEkkZeGdvrrA1mYGeQR3lhEQP9FKNz8vPiL7dGw9DCPfObHwJ+7ymSOH
htGudQrkqPYxTX6KaAr87GPUjhBJ
`pragma protect end_protected
