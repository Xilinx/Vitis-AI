/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 976)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9duIxhRaZT41b6wj1Ni7Pwg9OTw4eB3A3SLLRgT2y5tJ6sAi67Wlb5oc
bLjLuLqR3ggdW6dqHXouUeE8lM7q8v2s9iksmpSp+70fSgHv/qYzSRUP5kXCcb60BHh+Ng1NP044
IwU26axDNnEz/RfuJfHMfck1KghH4/DqWz7nM9E7bTTkw1FjK73fEMIhl2stwswsFpIeXYRDqZrC
5nXgog53i1y2VjaGbH0uxj7Cviv42TSyLKw9elwDfeRUTd+jmuFc4987qjz1aUN9F1atEqL8L98S
1XoFI5m80ORLJy4umAUn1xtowzRr0qwoHh+Z/HGvhBQASTiqxOfn34s005va+LPdKWXQ9xXUUmBP
DNIAVjqZTNwBTKZQcrNFnuZxn34G1HY05Uf1x122Gwgqet6FtTgsPHbad7G9etI/qGA7rZ62SBJZ
7JiiKPZLYWstlpuPEadekDqUzqEw90QBK367jKDg/Rx2DQYhK4Vs0AGTT485nC5LTYxyGsBcy+PV
awycyhX08zMUID7xy06/UPD57INjGGUMXAe4U+nLvQxQjKrnfk1XL71frZ6Fsh7/zWESFKbxVYrY
TmBmBOS5j13SLer54O/zug6y60SlDYB+WftUMdUVgCLMVoHFRn3SkmF3KsuLFdq22AI3Y8pDrvDv
faLEr9xd92Ty0YUWUUwC+jYNYVoDm1BE/O1pFXn2UknsDOaG3zqW0gwECUhJp4tFUO2LwdropVcB
RAkRibZ5I4PKNkRpIIaGQqR/e1eRzl1O2jBYt5HpzJi8vah33U5f9vPSOqOk+qudGoEc5HV0ApGz
+P6xhIopPXfy5zubtlMWX5CJCVtWSM3luaRTu/7gLPVZKtgrLdTsHndABIkGdLhF2t0g2iO+FcS+
Sl1wSHCbkGjjDz3907fd74a8opmdN6Ltwo37CKbI4fz/xa1ZyqA72mwA9Q8S6ZLhucc4Sk/mepzz
wwWDvQIjyvb/sOLznikr4MpN9Ypy0diuWr2BMAVjHkj7ea0daJeE7NAcJz5/YtnrwHWE55Q6/7Z6
nuevG0qFw2DDn4VzaP0XVWx5tFPYp/7uYO1b+qNDIyOgjYA7B72O6U8ihsF7hQhi8QpT/GQfVfUX
IAiF5AWKqlVP8RSpGxAUwThop2Pvb9wEOgsEFTvZZjBGHmPHd42ECclSlPLqGinygIDj6ELuegZb
OA5Rk12H2OndaFJfmmv7Wdp3AsHb9EV33DIgXDXK5NKXNVbHuLXvcQY9SRBAcmH6a6nJ4NQdRdjO
DCqh6EDUrQ==
`pragma protect end_protected

// 
