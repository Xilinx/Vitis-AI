/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPS0AaAQAxq/IXw8qx9o0tQPmfA/rDkwLQC5gJMTFqhmQFs7ZVFWHODAPG
pWnUgbjoEOJJaS5ds+uUVAsnoL4dPFOHfrckjfC3xNPRs2cyAkEB1BVeeN6CRP1LsO7aRxoI1aDJ
K6uGV5Lc4pb7WIYV8vGun2VC4aB19aHJWRYAxAE1lIvrIQfcThe+K+2gOocoRuhBejwg5/Ot9/n7
AaFHk5+bi65QxX6k3TfG1f9ST995qpxM4MOfWmcQymsSCzm5OxsatpIrQCvtio9YhMIL0D8xPwDt
r9/BQsPB9AMr6KWHIsgOPRrxecqTxM/4dsk2/HegIYKKBmYJB/xwwuHumBv+G/VuTdGzTYjHWByo
7CCDDG2f3Cz5FMa4M4IEtUqWYO0TxDUKCk2ToOV7K1Ui543NXe2VZGjpcgeqkohFl1iDH9YjUvwy
QU7bmStfdcOA9h8vviJOwsK5+YRU/DptZl4qPAtPZsMq1Sob4KhiGE6zUDAXLgNwKaaQtDjipxOW
mY99puwdTnz34NEmo1aS7C/gDznxZNLA0Y/QVsXXAb8sOFrN6J+1Znr3e4yxzaxsbZ4M6MWieWb8
ZcZlNkk+YqT0jip0P7gjf3+QdRBdueI9dOW1cdF75kEnacPyOuCr/yN2f4uxjPoXwh8jIeUe6kYW
b6b/pzg24rYUu0BddmoMhtNAnXj8tCoQkLzXZO9FY/2zFiy/4+hy35Toe0Hq/UAY3IWTFfSoaOIg
rT/bZXZcqwi3cwRBux41VNij/ppVyoh2tugKuqmPclx4yUYYr7yHO9bC44pa5yljCSKHGmCtVXdE
jqUN3a/q6a2nkey0ZXUr/fgDCdlqe6mbIgACqga8hTXV+vsmA4HWFu7DBSAoofFS/1wQLpMTzKFI
U0khbL0YNSOz5HYI6sB5JGSbeFmycrT2tZmb0hQvA1bSqbIUuJc2ryqMj1FGDcGRzmfqlQ4E8Lju
chkH7wxJo4vRU4vnVt3tZQvX0o6RBczQukQjOniEihzOCMyUWMmx9c5mDvAlt4CYAEbVsnzqJ4vD
nyQ2J/gcFhTUW0EyQHpCEwW47oipHwq2c/dv4YuV2DJ98wBOeId33TlFL4/kDsnq8DegcC/bWtRF
3xXACSTSbph7hphVoZ1c7WSLHIM4jV3FlVZZviIMQH+gyt1JaPaX80H3Sf57ieIlwtLC3SDM81lg
MfETCDg9TKv2oISz/qSeOz6oHX5KVUVuG0Hxfa9iV7/kWLC7L6JStH/B3rXWtLkim4Uuk2bbJ/XX
L7rnImEarz3receo5oA52ZYT5xNOcqw=
`pragma protect end_protected

// 
