`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55712)
`pragma protect data_block
giGA109OWTgnmloyaK8oODsiRC9RZVQFcgf9mR/obyjke8kkfwHUD0rFD2w6Qg5sKJtvAY8b/b0q
V+Sa+ZX24LFU4BuS1vxLWFGohu1WaQVSB9HQcsOWHML849yQr1UuXHS1H7VUn17v0E61+/PqUzk1
X19/pJmyYW1BM5ZHOhJulHdCd99vhdUA5znwgIeL+qkiU0sf11eCHljau90FYmDoD5m6woWzKvoP
6gHK4sf+uEu6z5A+3PvW9Z9m55mkt2a/UNoD0i4Gx2DEeOPjplA+7mP3yNFRQa0VErXtpuEnDzdu
mxNQHGYn01YlAL3b2LmmbfdhupYbEh78Y26pBChxvKjb1WIDRSz7ZsN3DM81lanXpKPW7xCVSrZs
EdcgJMnxUcv737gXGgSKQFKI32Ob/mtOBEguo/bSd9IouEw99KI/cH1e+lFIgQXnrA85x7sn8NDi
KpFN/8LX8V2ijsNcHnhiAW7BLfL2zomuEBxqHqB1FHYhE/7Nzj2LV2dQ4ZR+/KWoKB7/dajlfbFx
Mn3SlUUvS3odLmor4IJKJTWNJgn7RJdPUuMMRDiJzjdNG2ooP74eKosnYB8ET1w97sq9J9kBQOs+
w7pDVqGtJSHk+ulJK5NGMXJt212wwHKUTcyT/yQNRKoKKHo+s7Q2THcVoLwnEfA5MEVcngy7xH2L
SNtBAhiuluuFIjilRixC42ntRTfscRMmbzhSiO4S4LCquIgTcxRTr3VrLGRD2wyq/IsA1QIKOj3z
PYUfeeMzy0E/cwtHq9Yc0DktYmXv2hNEA+e+G+mR/TARQJTivP34yz/L2djaUvjbnH2hWT6Gkwsa
diX10zZB+za9GemHh00H7cSPcBOgTQZ/KugldStCgN6LBVx+qjWBCnaSwbrL9NBq2aTTTJPY/ffD
4ZZPC0fzEEpKgDBT932TPzJOKwqN+RGZu5z0Yzg89sZ21yq91P/1DJWOmwA0iPn4n8y8ddLmh2uV
5Ebvhay4IoHrh0T9vKUFP1/GQ05ymPxicE7R3Iz+SG8dlMdB9yW/4YR/o86Y++RW8Jv6KF13jFCz
BSfTRVhGjv6T3If48Ji3LFxQ2Sx47pLljVmHawiFK8LVr9nsqsT+rEO5m+EX2F1HQp52K+yVghcI
4R4i2/c6TWdmVduhYcIY3e3u2bWrvmirP49gL9Aq9VuCjmPvWPz0DCzjM3SHiXn/lNBQXqd+6DQm
OQvJWddLtxUfHvqPyNPGM+7ZafOcsiakrxwt66J7XWJ3dhhiwRVQz6EE0V5L44YhNtWTk9+MYjnm
IAF4K3DLmzK6jq37+sk7o+VKvbslGWvdX3B3OvVL2ivwBMsCUe4FTjIVDc2L5q6zDRGUQtzsuGn9
3F7p2x7j5eUgFD8e4mZcypT8pko5al3mFfyd5auDCeenPfGVlji79eeJsv0UgE3QI5wrMDrQpjYQ
NR/9R0exR0UcpIQ7y1D97XLt9g4VV7Nu1RE7ESAJ0aTkU+xjbJV1RjGBe0uo7DM7nDp3/p3HcfqG
Iq+m4M6Cl+ZMc7n15CU96M437xhcV2yInO1ny6ijuaAt4y1gn0LEojaBEoTtGNrHVTaCOdMlYEWQ
uH2t3Qu+PNlbibqAxjFIGUCd6/Gmgsi0zwCuyhYYzAeqXlFi7SrB6nCgfrbkabVpnw2dHHiyF03o
0W8kqXbH/nV85X12PBEfV0Euo9Qjv5rl0Q30bVP8LY1kLiBcBXtMgLIRRH9KKf42PXR4tNsCLTCS
oBPtFjZfcuSZdHb0MJ5hoUe52pZUuAmghTHRxo7gzFfxWXCrUcpYPcJ1pQc/I1U65rTEjsaPCL0M
cKNh6F556yC3+7UBiKbATHI9AjIBFlCk109ux0MrzahsEQihUAh5M9TqQuMTf85YRtXPnWA66/CG
Fe4dhpBw0d3s/A4mFQkRGVdN3zyGaLEzAVrhQDQrGyef4NVRSPHPl7iFAnYmFnvxRcoVrzd7B+08
e9+Vgle1R4QCk3kSvByI7GcRPNJUSw8XtY0+ECuNnVeDDOct7dVM97FzikCEJkjOC+ZbP8UwIMjR
glEB/By5tIC2lz0Eaauen9xS9i4f8PkzQibL+T30tFgX4g0ke3sJoVpa1aRs3bbYyR7KhEfkirTb
gDIlmymoWnYzktFaMf8+ippx4t2Zyo8zHBMGSi6qYgjCnRpDvQk4m88SEcMwG9WxQKOmUopyJWXI
sSXlyxd3IaqLD26Lx6o7YpH0zmd14jXNTteZT/I+S695G8c/qlOGlkJP9KBEcgI1HwXlEDZgkvXW
KZCkbg+a9uUYAWrvdS7UHIIsnWlY9cF2UPAM6lCkyPJZt1gZpxF70PpRQgvq6A0zYlNMzLRv0Gqs
ea8m4RV8mJYinp05UpoY2Oa/obIBzd+B+jzDeoi2g1Mj5isjOuZEHEfxrB70RGiwsQKTbgHXL/8U
sbzIZzArOP2l6SxnhoAFTbRaLday2V+KS+6Bb0Xj0lDF8i4SfsRkGABSAkeNmOwGRNKHumKrVxKV
1iBUU9LHEuX+FOTvG2S2rEVjEVlD0F+H2jh/mlfif5VC46WuwLAbs0pEYMadezIqokLpwvjnxIhr
SK8EYCiTOqpdJBwnom1DdVyTgC/xbgL8QA9PAksecIPWAqYI3/87vB8r23PlSJo0i7anYZwJIu25
Xxjs90FFFYeIoRyohy/wOgJ30k9cpts1k+3Up4m2aDlAurt4F058TpESwCQP13bAdzZsjwMrRN9L
z0IeVbs3PSmjV4AhHvHyZ4keeGsaQMFqDT759MgYIFnCIp9MwxyFib1IMTTGeCRt6srx5huNuq8j
y6rZi8IPBP05IcFVttOb2/E9OCgTuoFgj3prkFq8tPcFxBD6vWpsvsr734s3a2l1XIg0sM3PNCUx
amGQoBYFnUYPPvhe1F+WKIohsGdJhtMHPKZYL2ZxnoJjiwjtvko5qMzxtY6Qg7aw82NeGTzHwlrS
+NknmI69hSmmvVSqa3UBm3VcjPPj54m6mO1rSRci7ld34bHtqavaefbECQVfX362TA3WgDcIUe0B
PNXyFUxDGI/0xTYxfdWE252buMztPbVmtr2B5cRWeEPqECBzbZIJRaTy0sHEj9TKX63p1bM9PEQm
EXrZHTXZuYGxKeXauaKKkYb6IcGtrKpu74NUpbJ4RWJ15fgVdCDKPgYcIeBqa65KRoBmhB4yC0xM
0+zpis9JeFwbRf94ha5DhhCOVFBobT3DFOiOft8lk7P6GAU1KH23s7WZ9Z9JAAfi8HAmd8+ocp69
n7yIndkFoF/SRQLbqdbpe4FrGoJQsYnODqJXgvbzzqppQycd2dub6WsE/eDfGQJ2GRPgyXfacFUd
YGldhGX4sEjBJWeriTyo54NQKha5iraSn9y3wfsh/52kF93Dy05zyvjggFx97crMWPqNJTvvND81
0FlNUv1eC9R6cburSVDl24B1GkcLy1JiZl70Zmxa7dXdGnEPOIQXq6TdUWW9Tleooa7XQsgyK96T
jxtZWYupJbEQv29A+xqZ9EaUb5T9D9nYEyJ2F+quyqIuImX/3bG0Pz6bfilmODIxLGh16o/1YvYp
5/8Np9z4gXq+ARFSgVixY7y6Ug1qYYTr3UmnraQooQUb1kNIhOZ+6mpkDIAyjAQXy6/SPylaEosB
lhl4zDYvrcBhFEX0wTbizTonykwcvQxCq63/QzfDcMggfHT0nps+pUxc6aNtAn8JwSnnUXyUCWYY
dd4K0m7qne+n40czYxv2nADGwVVrj6qqq7ZfjOVDkydZSeYk01sz2YjkqS8ewaeG4cNazsVqt40y
TUVb92upjyqoB5vK18bhY6as/CbuxI2y+HIWaW2F5rvNPonh0P+EMCIUg4IGceuk6PGnkl+27NZm
9LG7vAgxBjSMjSTRD+5i/sBOMEUgLAM6ZZfayNlm74k4fBSmeb7pnay+ec1y87dKYSTX4/biWJs8
JC9SAZmP29/ELZ2jnfITPOVNW5vSENWDx5TZVxx4KQ4kpZPcFNQTAZT/JSquuZdd0dDCH2FnNHch
XkLa57KZLBN4WxDJqKUKC52C9zyinWxtS/rxxrk69MhXMrIIxWLECJVPs4q5WHPkjkoDFZKGghYZ
kC4QkOR7Zsu3M/OubLuYClWPVFDng1wlihRNHameknktyIaDFpdZndalgC7atJCEoFFdgrJ4B/hO
XWSx7AcaNnAiUlBmXUvXXsFjLPBLqU1hKyQ3KlIJExufVVNuCzCQkJifkWc32N7lHJymYsBWV69J
hjwb9583uaJs6vrS3yslt0pDq+MPQuEcmz5zNx4ZO5qCokzAcuTuMGhwtc9hbWEWUsIehX5Tktdr
gup2lhkB2YiSEXPzHA/nMHw5zfdB+3wU8TcrAKeDZqaZcbJgQ1wJJRcBofTgNs8MCtHoBE3JYLAR
mnk2NijmX2so1U5fk247jjfPvN1pZ3tS59kOY9mjJ3WfhbAy+2VsjN5mWInGgwDGNWib/4IJFMS8
vwxjAQOZ1G0AhqEG02zkAodyH5ymawNa2p43/CV+v/PA1o1dn2tobeXdvMdYkA81QEnWfbj222Qr
An1wHz2CMHNVx2Y5jkzKJ6au1BhnEBwd1sP+VudoF1dca7kOKgeU1lHvczC7hfQyA+QCbfv58YVY
dt+ePpip2cAFCFZmuN4Dd08fF06eSMlt0NtUsdeMuB8kDQ4UEFMow+k4dQh4mM2NNEzrqKH+jM2j
QKdShANM1QWJEt7RXVij8MBHI34zL2w6XQdvQ3MesTTMytOVpWfxMYvN71UdeucF3oQewUMljQNy
nhHjH8rTISiPJxiTVb0/G7fsChP9+eRV//y/oNuVFyIrT+OjWPu6ume3P1BvCCjHTIQqvkZfzRms
GAmQYC1maj0/TIhhPhWH2bhjhRAsHCrhYI/Z8xYZ6uaAqbUpcEj2THg0cq+7rMU7wpRISuBMCYZ6
9gGzaTtB7McPow33zpMe3AJUVLH+bEfyx22m9Jjv8Ul+6uSdG3Ldcspbxgu7XRhCGQUOM+PB0iFA
FGGaJPYK6GciNdQcdOt4khX+RD6LqCfF1gCaMG/U4BZ0+eUxnIH53hfSr1srLRY0LyMP3l0E8qxy
M2ZABQbwjaLHCC2BK5hfu00CubvQIjvkNCkSnsIvHn2mm+rprK73GPMs//0gKQUQ8S3f8pD8rWb0
c/xMGq5CKO7iItU07HrcQFmab9ULnKC1yk1u0loNDsQJsQodHXEn0lgYIPaEtN/FUpPQb7NwaGBM
YxsUuFNDZXGghjt76LZLZ4HBdnylHLaQ084dF6KJdItOV/kOZkDKirjRS2dVuRnHb7UTsVNHambq
j/ews73VOhetRXF83amEzfALILQlmSlOJzbwIxNMF1gXEs0bs2UOt8EfPCvaWSy/gVzx0j6wG43K
eMcd2TRoPbgaGjurNSpMwecJ+txeAk1OqMSoW5QKr+ggqmk4M3/dDtbtx1Ho9MNStjTTYduRA+zB
m4g/+ZPUkuEzHaV3PIl32nkrV9qSK9M9TGqVbL3VYl23mRizr3T/lspH88YZOUXdKSLWLZI0F8Ov
AnqzE3fKM65sFbKcyznVZkQvW3Lx4ROMyqaA3Vf4XRQNc+dgf2QCcGFJYprd/o0cxqgz5G3JYXwl
3Xookky3qTkdE6l7yl8xbWdnHXV/zD5gtq16nSP7KiANt80yDrG8JUNaIbXegO32JahzbcH68z+8
RaxLA2dutbif2wv686qxMz3OjpyJYXUH4EdgpYcLEo+VL44yH0HP4zdT/hmddf/lAtEUzMTl8Mi4
+WelVS+Mqu1qMqfvjsTAAGyVNuGDhiF2oOk+r8GmcLLOxDtpVsatBHSjJjqGcmZBRqzBxu5fX/C3
e84XUDzTXrifGmf0HunY/uz0S/i+VUtL+NHChT0h51T7rDRy1VtIWDWuDyieBeuxDumDQrnEMKHn
gmGp2BX2op5/iayeH3kjlb9RkyF9qwrdZqUC4vglCnD3eySorxYFH1KLhdl/nUDsVewCYiz4DK2g
Xm45gVnp0MExTrzcuDWIuSYlI+31VGHEnfTnhTqR1zH1BvW4PPR/rybyx/q72/TU3wWKeC0HnE8Y
yDEYua4SitEVlwVHOqfTCt7Qukdq0QSOEbcjzEC5rA+XEu+hzFSIQJkzKy1uPQ9dcpAuRy+myC5y
E6lGK/gdGvbFW/2SvEjfPKmLcZMqWTvO8PqsvUr4tu2+I2cC1QZhWRWyLP5WuN/MC585Hot+1A4f
lAWYXGhwHAdWPGCo0IL4PO21q3u9YuQHfgWc6CS5PnTP+C6oBOCUdJKYQaZN+Qe8u8Bd6GBhCGlV
P6mZCBqCRLRGQhiCIopkKMlLkXVoWSO19yC24P7Xm9adbnRNbJxhgDDfmsgrfvd8Tyk7A96S8WNC
NhjvG8eU8pttVDcbKl65rs1cipZw1/w3et5hwa2XFQWSizYzqacd7b+fexERxu3CKWaUKd1p3TnF
FmDeu1FzH0Ow2blC/ZGqfqQDX6GSOV0Su0qFPwydnp/PHZrdrM+PjkKIzX38B/YQ1xM1jsoS9nKm
Ya3aLzbCNReYkClUnvu2Nma8nI6z0GwugyOga09IsyzrWXymSGSCGDchShOHBHaH1eCtie4+OLJK
T3CY3/qMhbeBqSY9M7ZVekUdZ78dZVMwMwKuInN0erb59LTOywGdh4WVJik8FgPrhYhwepYDT25o
kzb27myXvMOMdxuNASm6rqF8Zk/uVK3rDqzYFscYg4TN44EsF4x3mVf35mNGQ1SJgmYnVoQtbc+G
OwCciL7MsWJ41efL1Ev4WnfPYfbfuhIpL9URAaOmS9TYt1ao7cjJ3rlqUMxRtQwcHeHZPYgm+6BN
bfJBwFwlSdf2RcZAnbqVVyNHEAtwr5CsM44rAE69h7viv2gX2vsOsvuPQYvRgMWrxRp3Cvsx39KQ
AcKuAUkvc2tYjEsgs3sbH2d8h6gtZZZHoJhdnupvF9DrwTaxGUK6MQ/8hfebHSS7Cj8FLyhF+5qQ
MGG9wRw4A0l1c2aNAgPc/zs6v9eCLiPP+m9eHrCZG4+gx0+D9dISNSey9dHou2T2FRHriGFeN/bi
/56Dt3I/fznol5O3bLdZlztKXPTf2j2qAtxKBIAU4sb1cU68ESE5cuOLnmcCXe5thYIqVQ7AgTuX
p501AwNrk6gj9Hg0YVJFkblHtg5XlgvTsXnsSfAiPI82uhMpqc1M/e907pk4UStoVWc+0qr0W/Xc
pp2Mtp1/XYiniK2XYi1+SQFoFdDKEY6x+ZBUanUvpa2/vPxbwKGSQ4Qm/DCiBj1wFX8YdgbC2A1D
d3r+0r2pbQjvMoXJnTtrCdi1Y8io/Pj8z9iXUravXOqSlvmC5O4p0QPEJbhco3vMyEvGNu7NaeFn
CpsETX6bVaHYfqf4ObeL9g2fufTXpGx/+rKgevwSCErsE3rqcA/zvGS2A7r9fD80Jt1ZvohpL1RK
puD+HhlASnhKRwi929aqijHkiFQoihn4fpRZF+f1kiP8v+FINHJgRtyQHa0Bu1LF3EhThiYg787V
NXCw0gjyd8GgPNpjHL8QMLgta+cxCHTB0I0guzqdIXmhfzPaibTHByENJbN9tmqdJe1ZvKDXH+Xz
0SDXZTDfTJ1ImXfjM2hQ2ikh12Zn+VVR5ymBASjjRv5ypQMOWTVF4+Tf8MDvteKvS7Vgjg0YT6GC
T89GwvSfCJUPXdE+4uEGIenW09id0FHlOkVaKGM5DZTre3o4VTy8+O+O8jBLhz8lG71YKijZUhEQ
z8nxPUHOEFo7GZs7oPV9fGeXkOxkSTXyf2tVG5mAJWQH8xR9IZxW9+MwR6SzuzaWMlZ6+oa5F9+U
B/o6pR7L+UNfygupTlNzSz4KWl5s9yORLn1RMM+58WWC/Fr6O86cUdPqvAc3udZzs7f0Q+CLNJfC
9lNCK69C76V/HjSXue4yCEpez/FjV0BuMEHX5Ac7ffbLy3cmxl4/7pH1tbWUgQYGnp8zCZgELf1z
WB6jxCwKYDS0jqL+xouyU4cWSdCoqgsd7OrpJw+9s6HaGxPI4jfcV4vAdbi0Uw0q4cgimVscesO3
1NallBl+KU1oMQH0WXNf3qk+dbL6bO1N5QqVRLOjKtjw7npu/Zf+fZFjbmH4jFKeLr/EIZVxYuNJ
9s9pTo8RtU+3wwFP5geslCU0ugnO2Do6Lq7Eh8xZe6ALC6JQZiJ8Ynb6wdWoDAezQGN9+sP5+0RH
mGJM5clMvOLydZsonzAKKsMvuMKBKZOO2nu3gI0F8iDLJhUR2H5RSHWSLNAoPT43VDCRI1OrdxhU
TmfaRv06sevuCe5kRFxo2hgY1t7aQK3jjjhCI71OAsSBw90u7jk3PPCS8W+m5S3vIT08Z/DxN8VG
naBmE5UZVcLVe4Web7S4XhurOWB0cKvf8gPcHLDGiHfwgdweiOhVEEHDOnLjpTh2khmc0maDW+vt
4mDUENfHLkp7ntU3swAYiPAouThG10kNOMmXMf3DhbsXy2wQqU5ZlGyI3qa4jucRosv6DgxH1/yJ
DG1bfIqlALRg4c+J5C3j7vqUIF0rUBwVeGYzab1x655Wvk7NJVAQ3PhPOZhzn5fYzYIvpCWbBf2D
Pu4j+CkWWp200DOTaWtbSZ2jSDaU5LFoogNk80Twxesyuw8t4XFI+fmeIgoTlnm4aPqhCHnHTigE
uRlebnX59O9wtDwfTaujccAIYV1lNi/mXTaz3Zyxi8g6GBI8C6x7u2+2ZvfHHpchXaIU7dbJQCrO
E1RndZwXPTB7+aiYHTGsse55pTX/+jmXbS0JFHgy20hu79qL0/dB08mDr7hxPjQhqUBkj03r04PH
J58AYbFU2us8o4VWrbuFSxGv+cJRpZ8X5qyddF7ls3xkrMxC0wztx1Ha4M6e9HonI27MdBswhEkA
gSFNWIuFq4tSoR4KWItLs84x50Ap6wR+xJt+V9uTu0QUIt/1LKOvViC1ClR3Snk72HCd29KoIt7X
ndUbYOYwvkS5ja91mG5Mz5KRXMfRBjO9ZwzDButRZ1HPbopeCleAiMrs60F5WBeVpajL2OSnruDL
UFkujY/bod5oK1h9XNN9vvXUspGO5K7KcrLFeY283cGv78jG6SeCoq/IL58lmjMqkn5C9n7CuX8E
yLiQAfUewaosotFTO4/RW8iSDiXzpJdb1bQt4QYV9gLbJracM6nnMN+Optp5VSMoWzrA9Ev4VOvT
kkta8dAD3KH9YEzyOOaXpf6FSOflpWIHfE5eM9OjFHyJfzBNHPvQu/8PoNKXiutoD+O0UVgWuFI/
m3Vn5kGB4WXrEYGAmjG24M2ghtcHCH6/W1U37WPa1zdRnf7CFX8AVTP1liSlWvzEXv6vKyQFakzI
xLVaH6EPhPMXkmPvR82t2Pvti/fbMWyVQs0C/fiObn+a18Nq9uMOgmr/kJILoXCysRxYZF46MZo5
P35ishQcKe3foTi69q6jmcJgLik4ku+klYufGr38Dd4WhuCOwPZz4ypWDIZQ0VzDdjmdn8zqB3Q0
mqyTgEWE+pmhpqNk1P42HtOqRsWx42DS7U8Tu6ovbsEwQmOhno3cmlf5Y9ZtS71VjUZ8lSMgEvGz
3UMofwe1RO4t0ZQUBVOS/X2IOHnBYzmpZe1Ga5SSVoEQM3sA+ZA3N7R2Op2adKMczeApHvv85rBQ
PyMS7g4uU2q+wmZRlQQaQY2O/XB+zeMxYz9r+bXadxMFI1cMEY6BL/f4BVfsiYrk39LQGaSSxNyo
pScRztrjb6bpjKkiwrpnVn0V/drsYlxbNyXZUH+npZe+vlg/FPSK8NHqHGZEkQCTm2/STIAhML5a
JdQRPqCVvC/VKP7vrfmocPp4RnrozgM6/brUJV6qP1SryZ7wasl0u99yp6iIY95WdQHKGZHASehx
ZQOhFwvz63uxt/ukOnPDEnQMf7PF0Mg9D0ojj7e10y+xwSt5mi+I0ezyAK2VV2UOEwq1pORaNUoA
JWmkaqLFr2FnTguU4MnOXAWFi4k9mdxxrfqXgt8YXoKjZ1M88lpi1nJ1eFCCEYhXX+XfE+ANNCF2
oA4hwEMQKm2TaIexHWXVourA31bMF9qkVKNE21qGuFVDiH1jt9+abf44VzGCqg0CP6RlVmXYMw5n
aUI3e5JrLfQlm3xfK5yRnlyWFttunF3cWpP30ZXv9UjpY0SIodMiBZ2O3yjpJHTV8/hRdo3V9G0c
SJKEN5VuruvjurYPQVgA/B2kAH31XPCo2l9+zSErO7G3A8GpqRoSmzZy3NdnxgY6w+a9lPMzMjM0
lX5KwelaUc6H4zaS5PDZ4I53nXkGTBoW1UqCbn+gYHOH36PhD5yiHBp8EFBJ3kBLFqhhmeM5cbXu
n6xJ4oZ4nvb/wKdlfsYf0PXLSHvTeh6LoJRn1u2cIVDFK2/eSBrs5THCDzmEFlYOeRkJ5DF0/voJ
kOyMmF15ps+5tNF/NM6EVRGOVCP5PAtwePQ4qF+Le+m1Y4C0LdNxOQ0U6di9/3A5V6M/pSPDLOm2
diGwphAsc5VbRCM0pXj3Q/A3saYKMkRQ6NghF1mRSHGDpMWhpyMfxP7xvOpHtXMl5dqKPvWAa72x
EN87x/zFlQ3o0A9t2ieHJGsAnLYh41IaENyARY8j8uUtkDlRvqU0WqJNcqFxiyP2/aENeL55WwEJ
LiMZ6XEP8WfXDh2GgazoUexB6pRnPg9gBLVk8c8MDe+gw5uAusgwzq0Q6BAiuLndnvO4v5IZJ9rj
s5PwSBM9XNOC+XVeAowDQsWIUDRySsZXgJ3WZDXYzHQ3t5fDdUijV8wZ7xevU5buNPM7PGWfmOTv
bnFDgrivxdWBFxfqcefoRlTesWsSXrpHFt9c4JoIx/mDrCi3vP+pADDB8I5/YRS/9rFxdZSwjgYk
kFoyWp++lpC1LeOYhEhFHjcQH4NwxiBRxsLdlvpjbnvLaHJ6/VzUwQa/f9DPS5PBq2wVYa5SaEN9
flGIZhPgutTtwrGgpoH5dvZDOor5kRD7i7cI9iOp7DOCo6U6lYRW8roI2WCsNHKoeMCR0UQ7EOok
d58llaga+thkHe4R7M2vYo0yZO/Af4+HoHW9erT4iOcYt1T/OEH1RVqFcov3th6VIRb9TdoQ7t+y
ytkJRv+MTYfbtgZFfW7922e7xPEtWRqtX0Ld/dvAXjwQjMOW3jIYHFrTIJRhcNbfJEzEzWXhvhgk
FNn1td1t2dhRyl4BFjbu5DtDpQ8b9Cgws0HnAIEv+hCXPfmYTwTmff+6hUlOSh1i55YmMiO/pxgO
aw/DGXGzwKSAqy/JGjJWabelG7psYkdRffLWibuwTUis9wAAMXC4nY5ipIsKyar/ZgnyknVhu/ES
+nZb4M0uZQr4fw0Te7eeTSa0r/FV9KjiUM4HUEPzdhReDzJgEpO6rNVT1iMmDTH9M2gJZQ3c6l7f
3JK7Si+yGwK0gAoauegP0muwEfbVbaFaRSMQ9Rne1M9ZG73D8y1vPGoDz/AECuNqn6rS7kxOPKWH
PxK869MRvEcYNU3lZWh1rEemjzcdl5z6+NhcTjcI7iaUv4bNY5MfK6ykOsguZKLvf8r29OIwDCkr
8fDBqbrnIbEZIY8gHmVpyTdy/TPYRuqDnOR644i2Myln7XPuRQKu2iZrDM/681tAVaO1Qb8YDGQk
aI+u4IMh9QLcvZiwBpS/tVZlG5ldM74xb3X8uQAEbGoW5ql24RJBXNnrQGH3XU11F5f2MQzoy0c7
JBHCA+8GIWT1IGS6snYyfFJFsOTHJkaKdc4oZj08k4uLFQZO9Um88Ewi27sB94cRiPky/I8o/UYd
b26LPxh0Ovx+XTxMLnXTMlewpLKSumSiqwsBovsc/aVBuJMZQjD4ATE4giqeqUTeRWQZSuvM6gQy
nSZWWsXvi2+IzWwIn7zLGx6P0YIknwuepbxEPe7VqfYEXegd1LTyfZYp0xfrNmFICMotHuYoOtLn
ueO8WJdTuvGwx7K95QfE3ge799ju849U+I7zmenj6qUnGu0SgNBgAUJhLFBLRVXL7ylondvW4W/q
YcKzuXxxve7Zb5hk23wGPDpt7YpfqgwdnOWdQm+YWmT5B841VwhEuov/7xoqH0BG0yZLPPH2i0gZ
zjwkZ7KPKpLS3Y5StpRXkvjbX9ue8gJwszgbZh7PFV9Y6q6QD9LJ2twM741ge50G6jXaurwdGSCg
WXVlQxvvj44c5sBUwEV0o5WrBqk03iPtzInENeH8Kc8bhNOnunekXcnFOw/aj2o38ui0Y1vexUrO
XCM4EvDZZ52ZD55fscCSdtKDQRrOx0CRQu8BqMLI1oHqKE9lagGcX3GjIbxy/nNMPVrtWKpnEk7y
2j+4EUkT4rdZ01XtqIgyqUwuTzn+uJmL7xQYubdmS3bX0u+1i/gSKRT/HRiyDWzNVYOax8NT2Yxt
vjn1maxoeRw89zfz5X0NAE60KhcQ/fdMeS93/EwxmwVl0BDtRJUw8gPzHKLGMpL5iA2vGklPEixv
Z8hN77vOIcF6hXEv9BPXwHcesHKYFf68eCFi3I5/F14RSWndzZBlTpwBN6GN5WGOfQ9PSe+RycSQ
3zH/36OMwEwRzr3NQ8e/VgTUEmfjCwykCA/7stlGhX6fQrZKvG83VgoHcIJAmNFDxXWN4ZPV3NJx
M0Xf4fUGajMtXvlsrwwihmc7bWSLGeCGXzDMwix6+J1I9A+9R9jGEzcjxYgwuJnMk0TVGL10FuND
+HmjUJj/J8gAkcMkAmP1GG7kfw2+TRXEIUqkcvMGqT/eBMyFEyILITahmuQofle5D79z7ARWRg1E
L1jQbqeEzAtrLZ/0w3YW+eqYDvbTCXcQ6sr1ah6gp+VoSLm59G4JIfqqjdarhFvLqLmzhfjOGJsl
jlEza0OAdG1dORbPQPTVKkKZlVum9LyGEMeFsMKRYp06PI7DFUmQZm/m2elghbSkMTLlsZ3tk2ca
mVkV+jmjDjPRKAG6WQONr626aS3lf6S4+O7Bw6+FuRbyrtHo8DbMu+byQrDAjThWz3X8NNArcm2i
ERoLg44wgTKeujBL28lYaDAd7rCGAbFX1o5t0xbdGqvoR0tH/ltHfB3NuCkWG2AznofHu6KL+QDz
4qilvJwcG7mwolMpW/qK8AYpRhq2XylC1kNsu2cwFEC+ZkWpIpYHf4OPe0Q23mgCeoLsQaxz6pkn
JnM27rnp0+SvU3hyp0ijhnM6AHVRY3ESmxpEwlx3XThZKhLQnNcENl9/A5MKT+w/j7J6bBoZHJYB
/UYz2NDDLVxM6wn2FgWexQ1W0YBNYz0etViNHuWnxpJeO9Rng3DMZERknBQ/WwZrj8NC0uYsITOR
OWOs5iOuQCh3KdLqEt4MhWLk1rzcN8tp7qYEZLYMnKkD0h4Bzs3Z0qCXhauQbh5qLXxg35zGOa+j
6VWanp2WiTaGXBM8jaAR2qUVgKs3BD5V4VnMbYpk6LHsBUOExBKca/2Ipjita127W+W6DWRIUxoD
HTcjhQ+9wH4x/XjFmZSAnsrdZOV8azbnXwws4qO/4gYzQKHtr12rXgpEQ38Dc5RUxtDZNASPdQHT
I77Eq/0FV0nNE3aw73a1GwPgkb4H3nX5SjuHZBn9+ElED6TrhqcWbhWCsHWYyqYxG58+lYBPc7tW
BwkhJXT4Bh/znWMaQOGej02RyKDHaVEmxCEpgNXMCUJE1ru+8jXHpmRAFUZLxtTuPDHe0MXWg8ud
0wxkAgIN6pfYPAtOhkpW9gLn3meLIh+SuVv+H4hogJXxHBEVHKcdIMX/IJwdTOrG5Em8erAgRdF6
E95yB3M2muRoiHzAEtx8HVejlEMRgM9DTZvAEMsxGGxAAZy6xsU+C1SoQ7kQxdZue1mfbE5G/p+h
eMxCYkP7ycJz0cE4OGc60uOaBeZIJN6Ay77OGHoTSC7kcrvo45zpHTWvX7yGXu4imuNMsXBY64dE
RxlVAjMSQX4+BNJ2MKyavBfvPeNbG6Luh8tHw3b2GWJjL9UJRekjoM8bHuDKoVYQ6aGSOI6mj1Pk
Y99DITTrO8QcBeHkj0dofe3vaYTmNiM0JzkXD+5vPBDyHFi6Fu3cUriY60QKqPWJgfOfvZFUZgao
3eUbiYXza1iT1jfj5S742aLQWyrcHs43WxfJY0MQn8Xpu0H1MUlCVvrc7moOmaQ53Idn+oqqdWOs
e1RWyMAZurrSyKfvzVIq7VzmRxfGLn+z1n7A5H+uiss6hfaN9FkLBxlJyoFL5vLIpyS33yQhBnaN
0bLOnRwJRNKtaEMOOhFsuCp2OJjYoWj1OHDsv4/BvBexhD6ZMVmxaLBxOrsmQ927vXGTFFPzle9W
wkjqbbXlYe3icGe8JovzTWXai7wh8k5V514B4iWH3trFiqNtwYeYsmPeGSiYx+53d6CHk0jRFiRQ
0MtdUUcBoypMSQoeDlLxUlwiuJLZHyTS0GxeRINT49/IeTk3Dg3O2F0g5W62KV+6LLTZUQbMlvLe
PQWJCanBiQAy4YRZp45mGZvLY67AdJz9yjAy9HuEF77dUB7A4zDOPEgxvJ5N0KXIxw5A4Gx8ecM5
xVSmmJflSNK4ma7AWerURyfIZGvWxNCxOdyrlG5MV9dkOezjB5sgog5yzdRgJMwhMxKaetSJxf9U
05KcRYWx7FqHIPLHLDFXMR9bgWssxgJMz4LmptqvbZQkQV52ygK9RZzH0LETe+aciwS+l9dq+LW/
T1VH7k+om7tsMI87kKtfPv0zh7b8BAI1H3Yd6kAaD2TMhzC3SN5ayVVsGvym9aigP/6bKv65uTU+
XUhHUHEi6rgGoA2QmaLFrQi8p63vEuj+SHR1kovGIvEj9H3mf1BU/AMvXGFeVbsWC13l1uzH3iBo
oreLOaqSP0KxhLNvEXzXs79YFh31nkFaySJcB2XEz2VsShu6s6yv9dE3tv0VZcVqxAqu1OclHagW
fZIDUFSUl+s3zetcw+FJO+38WhzKFmG9VnogXUZqlSMtbijv4zSWOdfKNSAp9cbio17LAgdNxS1O
G9c6NAZMjA9ecvf+uHIopOxN6jVkssxD3Cbq5jgYPVRAdQejSA9Ak5ZLHjK0QwVUaf2kbN/XaeH2
ZOVoQ1k0B92rw1EILQN/W38c2Nnro9rVTbE8Wy44T51vPwAX9FtsvKM/gSLWjhq2VFwc96gbj1DV
S10iOye+zSGV0B9zmVKIDM0RruKEvMJk50rBX/J8glo4Fn9q++/xc+JXwYAdd/+jyKd8jJXtKLoj
fx5xAzQDCoe3zRYver9mwajz051fzOzi/fxtKF50TieVevHtrWm1ad4HoykiMBySVatcZG5ciuyZ
HWbJmYcl8QNpbkJhVN/+ytnFR2IVwrFF2h8EDJZpd2widq5hf7EwYBhKRWbLTB9Pq8tRrJGiZhxC
M9N2Nzo8Cei7ry6OmIEFV7Yjc2WuGxjrhVKic/faqhEWRlngsiXUS1+HTFEgDBF/nz562K43+Hx4
V7C7ya4vj2RNNneNWnKu+4Ac2qJGR939bV45mXGsQFgS/8VY1Ax6zkor2NffYhgeXg2EgEnSLtGj
5awtREZxCiFJi2Cps0Qkjsl2aAseAOYY4yaNYe4F81vh8sYMoIoMHoDTDjZsIZfBEACXEVp6qpIg
Yb/u1l6ndEOQYYEWOPkC8t6njmupois9Iu7Rie51h8rKqfN+7h1B03v9jdOq0ZDGoIug/tDO/XzM
1fMD+6/D97TrNG4Y+RmMwYazyLZWwOFLCBBt2E5tBGXamfN0LiDopn4uxnEkSUH36jmv+L35BGz+
EAfEofcT/55G7n6YxN8e6FkunA+eFtnNSHnrK66QVk4woVvoLDgHR/k8MOz38FsPCoMldnu2C/Id
7IWsZKNbyfz9eTRScpkUosoCmDEtjxqewLRZ0E686YANrworhSqg5K/ydiNYkliNJkk+s3UUEtu+
3xKzdQN2ghe4vEbslyJ7mj2Hmll9+ZIA5AQNSIDxaCHLe5TlzQ6K5o6E8frCshQhZ5FXtWCYnt4b
791jyWmJ0T1fVMnaiOt81j1ottjrHDQimSvHYYvlJgSZb2sucG+MOxF511BRNFCVOYX5Ryo5zFm9
r3u+d/RLLXbCTBzJSAmCt2902orMVxCjh+41lg7hv7mGc5PBEAH1PdJgh/73cIZ8DLlf34wSp3gm
RYv9VKyn14ZVMo2gryK+dhLWQ4oHFU/uzEj2HyLec/zqgpOsFqT/HJmFhN+PXmum+6Ptza8KpVs+
CNHm8c7cE/z+CJy4nKXj+H1zsjhKyAnczSrharLKFZ1yX/FzCeVMseoruqh2zs+7asZAo0Z3HvNO
tqLCv95mBwau0hIGtW6qRCBPZTxyLKWHJmZmA+qhjcGDR5GlvOZM0SrrGciG1F1u3nYHWoZqOmSW
M/lJ89UP0dR3OJ8DbgtahccWhB/FCLXk8nIzL/D6Xuahk+8/otNd8Lxzb2t7hbT4I84P/f1+7xwb
biSaBpFyVLKn0RcAbi7AR3vciGe7Mbd4QsKegTU2sJk8IXWAUex44xtC9qkqsUKSTVWjjh6FRqom
px6SnvYB/0DBQZqx6in7ZRi0PlwyVzzVfRCConGXvLYf4p8/Svad1D8RZew0m2bKebRZ8R2pi/cZ
yZI7h1SjXq8HlkyF4pUTTzIctSSrFRzoUZ2T7ItMT16LfEID/ON4V2ab6byyNguVFfKtNxAyGyGt
Njp0jKTJXBlxSu+ExtK64YuscN6hxWSufmCFNI917uR+fXVSpL0OdLDQrCq+2ziCMKmNELuS53QU
tCkMjC43umWhP9Mb7swYztwY3SIvihkSFXYWPoWDMgM8doz9nzQUTHCz/mXBhQmC+HUwlPaExDxQ
jGTkX8okHkS55KDRXuJWgs/1p7ridcPRXcAG50ZomWR5NL0CJAH+7BEgKarAXIsF2wl30tOq54xm
Bsa7QGXAXd43I7jjfwUAxzX8IARvbPoEclNOEtP1mRBDEE6yJIA69pO43VcQhu2feDQgkc2++L5O
Wp55p+JQnut2FGw3nKdcNsj4uHjdff+3Wj2BFayRI1c6kiVVv7cI48n5ntMEdY0Q24QQhnqoFUwj
5BG+mfowzH31FUg9Tx6Aa062bdlboepKaE2DizIQrVKltw2eGg6ofcuSGPRIFOBsNbJtw6Ob3S9O
s5sGkbXPwBFP3ncUmtbihmBsOfP4xOzA+KO3BamS5wFvfWqTcKFlx5XE9Ix1Qb/Vvb8hA/CXZ89V
z7pSHZlFDIWdvRNgC/z5pn3DMLiulgGRUEfHs/JDmcdbbCYfbwzSXaXvlsc9dfV4fQQEMcGNYgtK
6R1kyzMutnHReW7Sn6qbEiXaQ10lJBz+g119vlelvI2HfEGNmjxriAu6Jic5bYaA1rFap/iwiwvL
wIfsHyvNulqmnnw5mJoImtfFaNw72ZonVFZ1C7mxlItz9kyoTJQkvfTmue8MiPlhrU5IpNYc7PJe
zveEgEBmtDkiAsgjCCbAavKxgPDMGcXE9Crb6ku1L3lvZVf8lsmdzkwJgRY+fKcpNDf1thGCfiIL
SgPEgN6AlGa8jo9ouMlyBpK1VxkhmEdpUXndJcKX2FuHiUtCap3znD55QuJb5tTa/LTatqk4Mfo2
JxI13yvUSY2pKydB6f4KrEE7/GuUY7sO8BUMrfHLd6MxC4Fg4pW+HwRrclb74lbqQ4nw4Wqifsta
QgM2KGhFA0wqktFZO+LyrgDbA4QQnKdr13ocjYIxhSJqSPndKIQu3Whmc+DIm4K2Cz8mG5SKhn5j
9hJvBCS55cOondULiepA/iNixz9Zpj+WFNLEI8eAULkR9GKzj+gdskFXYyoR4rnVsLNKQa/npseB
Z18yrtYk+lZNk1ivbtuAURIlPogEv2B7XMhO0ARi8hp3P/bEFsIwbWMI1wOHzG+nbyZcsgCs5Ive
IGwOn1Iifg0MgDEe9cdltcavrcoxZompYqGR5KXGyRyc1wNFB3pyapvULD9cqqSl2yuXzG37j+aU
eG9mJkTjvQEMhHI2qxd8OYt64rVkMgHZcJCEhPjDmqTJjiY7i7rpIx/oUNymApPrYLlaiWzhIiBm
8rNFNm7K1dNmTkvg23MaADklbRCVE9jspRFBCutgWcSkH0k3GzXCK7r8ybvTLct6cR8qj4qC8nfd
/t6+dCJdREkSqhs5PhjGtUpEsNsjno/Ct/eflADloqljKhcW3oRxUU4+T2Q0wUn9pxzOKEX6VcI2
vJ0wlcySq8lSjWpBStC4goJkp0XiIhaO6rR2Oc9RPI5eQqWdmfhAureQENVzTBDFk/n1Ok+oDCPr
4E9ONiqljHDSeCc3iYZUpHclSXKgJvnN2In+NNINkYMPuYcLtjo02pZNlE9XOAM2Sd+wjdJgeRXA
rUvchjwSk9yya+D7/OTlSglTyYv3iNNMJGJkgT1cdEFqDj5PeL0BD75/1g2OLTXcbYnhYUutYmMO
wUr+eep0+gjBx2kLPSCo2I42M1kKG+foSiOZsiY5BdFuIYTp18ypr7sRxlaveN/WW9Onv6OU2y+x
nGi61fSB9pw6eTpMWFi4M5NbxV9sIV+1/SA+3Vg7OjW3zoBdnyI9uamB/B91ROsPhmK6bpwYvbOv
BcbO8GncRFCV+d6iF3uycMhFHDuDrc0CKG2I9FHCByWMz1eXlrzR6nb6Q/a3Axdv+KpsMgAopw2V
2vFGjITtvTOm1ixbrsAZ7LbuCGSQBKmcWAssjmlP2bl2rY2fzI5uqFcq33appKSPcz41pucW+9nG
LnnvDCXuMzPY5ADtWgO9D24lZWgxlvBAa6Lluyg7TPxM1xPuPcHSEpLwmM+3Qhsdthgdl0N9xXf7
IX39214vJyU1p7nxKHbIwcywb6jhskaxSe4alSpzRYO1zygLpIYYONqjn5fZr/cbja6IcxN0NIxF
PVgOai57qxX8aChD9SwCJoZcH8Xxz7WWxI2hsY2X7exMSPcg8+MvuYkGN1CDWc1FZWYupe9mpSaV
SkxU77BLDN0JqIxB3EPCAKVNaUS3Y8lucLqoMgi9yA+/mTl9GzDTSKljjPUsVvtVYLMvAPTzHQek
cnHpwnDVLN5l9+Li+6j78tHv++kOBX2V+rNwA8bIEbzK6zOxOAMqqFAw47n8KwMHqcI3FmkZxakq
llZk/szrvBaOTWlFLvTkk5xGVQ8r6rtIqXKA7x4/dTunfJXut9HOKKJnhd+foKO/FGYDS/EVIBha
uljR1BAGVWxVSd9Wq4eelYJvoK9N5G0AHMfvcIh8mU3cbVkmHxo83JmwDUuxaznweWf14b+Q+ptG
QCcItqJcPPG/zSD94xoNDpmR5858jz1hT22kgav0GBo62vFPdsCO3jOPNtI2HW4wXpn0h9zD8Vd8
xQ9ecBIRCFYMb1xF5WA2gRfiW8plIyg44r06XTeFS6AFQvtHatHNcGdETRo3oFiUSKUHfqeBcbRS
j3MLy3UgaGRgGymaV2YVkLp0N9S/8ObZZqm1wQBFxNYaW+PyYjJ+y5KOku5GMk15Pj7LL5zqlKUU
M4UhaY1CJU0zWu/kBeMqVkmmxeraUw/vX+76qrFWlLjVwyAx+96+TI3ihoWp7HdqUeSfS6VdGFi4
i4yGKxvlnndSVBX4LYFovk3gnCIXytuHDkJu6jVjgJXMDjh2EuyslxWaxdO+1PTa3I9I1mF3zWMA
9PvMI3cdzFp3qvdbIfEErCIipp//i1midwiIqDUu2oupL2Wd8cqp8TRQWqUb8XV9/m3Y7qmFMtuM
2L7j98g6Or1u/zjOH4j42vBGC6IK0byfA8suUBbfzXTcNgqW6UmBpqINwNpc2Y7e+tKCHGcwWirM
K4f8qUfG2VN/eGk2mXoyuzwiRLPU7CDaPg36UwXQxcCFyIROn8e+ZgffDFQ7Aiolv1UsY6pvWK8t
W0vOO4HV05HGVfALu+0IWOBn+aZRwQSfXHHzHLeZrWUYVgHJ3oi9p7NTu9F1srtIeC94koetG5XK
4j+/j6iBj+ovSiqJqcuNwoOJKS+K/ubhFHoxTMNH8fuKWRXmHXYoYry8pFem6/B3w/m/5OSoqjWH
1iGbtVAgfmzuBhynLoOmvv4yVXw9F+JUfikBliM3cy1/bQB4fYGOMiFG8EaCoYVx5kS2i4pbI159
BoizjiuCtNhJl+4nSBgunLFrYK2OAiK7assYrCEtwMhJViAn1PmF9tl2MlL3mSdGQ3gHO/esWAQ0
2/H8a/geRANcLAOiqHOnPgNgPNKBu0wl9AKZtzzn+SsT8jaDJ7GNNrQE6l2fZ9T/VTXZECqYDrcs
ZiBmyj/xadFGXZ5/Xq8Y+Fx2a9vULST9oVh9Dd6Ago4cBXEZfap3GxJm17T0Iwb1g8/60SkFtcgU
EeDRlL+8FyI7GINzibHfNDKgdBJu5vttw2F4GHgHhrPIdGAqWsqkBQOcBPiikx5dUiIlyhwFP4IS
aGCVCJsuQMpCRlpKbqrdr2OAR37yXejX8hJ3T5wVukDiY0xUydvRzR7c5QJEuN5sIiL2yLQKDdjz
58u1IKbQce8rgPt9vGG3UxqaNMs6iL+2ILSojtzXsuJhNRNvRGAvVK5MgiLR/Jei63kOw6KdZkSH
M4PxQYaHZJCXJy8JNDp2bdKnWy0Wabs4qMfn0xf2z1RfGmOR+iZO2lPuoAjHyRYhRMaJPE9pZWlZ
TdxbCldvqoc+1ba2DN1ubOGpPo/wc8YfiVlE//4c1T+T2sjL5R/D4QUoQuF24DN48EzbehCEnScU
b0EaihAfbY9DUbWU52PT61WdQdxHnnkA0V2qNZsq6aY/7x1prO1OtJFiNm3jMo993ZmqClFCysqZ
YG0ev6VJ3cxl2UMhhzg90d/nA+0txfvCLHTBarb/JTunWWHIcl7uQ/m9kXWCJGdN9ih7yxUdBHWj
LnCBsvNVtXsN/PUyhmOB6VUMs0thpyYmab/1WKIiAtsNDxFGfIVoPRdsg8su6APxd1/uoLnv3Ig8
G+A59D+PvzRD+WfQeYiACrs3/UAY1U6FUFenP/YmUyiiwMytHL66EPQl6C3N+Z7yw0+l1L0r8App
DCF0NFMBgGJVW/hQUXmVVgn3cvCx7TN3w4rsIfUFi6/BBP7JEXYMIBYpmr4NA3ojBPToRdZBBULm
eWZGeagL34au6IVbmwseDzVk/oB6tTSZ7xANjq0STTgwGWM/DpjdUf0m6Qs18KHuq9eT0MVN4wYH
AFfYqKvzqhO0/+7HS7RIjawnNZiUvXM92exCnGDa+2tsbdAT0PwtqOIL9c/qXvWlVuQ4htAFWM5a
qeeZudOeDncWUgHLQKWyPRT3Ihh3/z+EG/mohC17EqP+Q7UH0xyC7wQlXjtT83LjJhm0Dyi7egS8
iMb9S3uMg29GZKlJS/cXjAOxXXza/wunwz3HkS8JXzk1AOgpHARr9uHwpdv2eWZ0CCfuMzm2hz8F
NHL3I2/SRSBtiiwoqxr+g0v9tF+w9GDd+0L2to6WfifBwv+47jdU6VY+6i51PjSXrLzR9OTw6Er4
u/LqFhKnbpz3PaHKMNDucC5Ka+Rgt6Nz+4e8S9jvDG5tulED/deibO2q2mBPgB55TFh0OhrQF1lD
639rRvkxe+iakqUueTzHugUCaOLXgBMvQgWtiOnKDeC+apwDv2zLASiffv6izYG7d92ADMgSsxgo
XUactFf6VL5IZX94Kh/+YBydvPzZaWmuIfkixIE2iw5BjQ0dZhUFL7vacLdVJgAGHx3v19Yet+NW
bQNM/G6WNoEex+MMFRqU1KBwcGf0GG1c4J+E7J6ou/igkVP479ceIui/roIw5iDvbsVw8niUxzEO
eMGytHoeEZ8ZoSLqRebK9UgLxXhAW+izdJGNGXVac1FoeI0S42MtSzjT5jCPYlyGtjtqlM+kEil+
hd2Tae6wx5Jy9tL//wS379GaRvCZfkis/KdPOesGbwuTOE5dpL02FcKVwcyikQLXuZxPNW8b4WkY
4YkRTSdDKAqpegK0DmcoWZJ1WCUhzucMs9keVfX8zTIwBc8qMt91Thzk2g3Mnvz+1gEef06rDlH4
YthSgzoIuBMjcNU9kYNxWXv75juHxdFPzJov9FqlCmQvLVUHA1N9GdY/0TQJ4CHutWiDXVvX6aDo
7IWZq+pUy1DS+WKxyQyaWOYY9wGonmHjn0XlLz8dtm06FJK6izltIxIERbpwsniUmBFOFibvZMQ+
3LYfjfKh6hOfPbgidaCRHHE9JnlEBoE0bun3xMk0Nb9n17duUhfsTc/eTxt7OPqRFUFZHnA70Cn7
9o6tIUyjYPY5CSFpw0ibt+9htQp5R15zShmHzsaE7loSTCW2nw+CCnCgH6TNl5RUVG9ODXCu4+x7
8F3kIEXatItV8+h1FniQ8rxoHcyv7MWIbCwkYvQzqspeesi3BIDXNDy5sBzJ8eDInGCFN0Ot2Nu6
87RbngUq3qvQdfAkNJrKpGvq6E74Uu4SeElrU7y7Nxrou+lcFrkGbQI43CCPko4/fOgrJ8SbpTVH
SZ+kvC7jXN/pXnIBEd6XF8ptwOg5N8LoVyHPjw5DaM4zrfz2HsQ/oyCxc+g6NjHTBnBVY1Sqx1Xq
J/KwDLszJEC53cqSyUCX2R7T9DxtSefSU+N/2kik+7uVNHUck1jux2TcvC5sJQg4F+CslpOMU7C+
bLxPuvvjDy+DGxGCEYRQ2wknSZNHU1ZGv3TD+PC/Bp87y9dTNmAP8V6OeXirzyI2ylDPswOHv7Pa
67RO6NOtwagW+jc8Fbgp/Om5WgSHa2/N1emnt6RT8gggAMnAIrtxasmHPFhV7lJhgLtYUtG6ghye
zLjB6r3vChijhbvSmQ68qQswbKkktWM5iXWcAujkHGeckzX+792A6hGvyItPAJA0PbfuLl63Si8Z
98WDSFzauB4asMX+cBfD4B53IZwXiuYgM7/spdebEYWAHC5GUcamRxb/6z4uweUIYnXFAGI9XUa4
eW0vJkoAtPe/sFIhx18Uy6AlV6oxLH7w+YQo/Vj80H0vc856bPxCs2x7qKzKfB3wgvCcx/28J95u
UXZQc2Wy2AnFIbHyoaWcTpMRw8rDru9ILbfw6LdA5IadAWZ1FPRscQQY3jd6i8fbfYru/YoYPv9u
Qv4I8BkvUt9Lw/lmqGmJH5X0/7L81oPzNXHKWI0Nr2LV8mRHPNB6as5qeJPWgVYTZ/UwHOl+WdFu
5WcDBtV7JzghlLc6WNjfohLHdkw+5kNNu9gDnYl83V2VthzIImX7dd66xMvgV4OZY1exbaL/CWDg
UWE/Kc/wLIemy1z5yzTXvA2QrUYAFOzbDoh/IQ+/Ce3CjKXhFsF+dRbr/jaBO4yVhdqU6B9lGkch
vKGm39jXGmayd0QAm9SrOElJlVIjqb6Rhaf5+HqBbBI8lznkqI8+zLvPuPku8tgjsru270TR18YQ
S1v7YUp77AiOqkYDWELJU+EREFf0DgcOZ7eqx4StABZ0Mt+9s3n9GtbPgUDBPSEonWGznAZug+GD
myWBWB9Rhjbs0W9fQ+isgOuwRrPcA8JWGfqcFy9ikBzLMaRSGC7KxhPxX9y01eyqv9ZdP7ETPvh+
wh65fluqJEDPvnYU90ZHWdJTiY3LOnAnTcMxGxAymKILFZADPuscTF35cCPIJhkkH7BWM3jlUmZ/
S2mynpgjBEixCZ9h2IhGs7NVPkO0gdq2Y/UyTROk+KgpE8uz2bch30L2zoYyK0/4hstoOt4PtE2y
Lk4xg5v+lnsqXV897Qz/RcTUYSbfi0qNpbB3+3l8jtyWWxY7f4fnBkqoQbuqIkruvHvIAfRtWa3s
bnkpuM1Z4NoLK9T3TTc2HLMuWVf/qJMLfx7gGdTuc+RthHm1EoyIl4KmR32Y9NAWCnmoCt6CaW9w
xHjFj+fmUE0Ia8zI/pyLgIhOgBcaiANrRZ4YbBKbDY68tbeIkaCPYzZ2bPwPGqpbbwG4IPlxVabX
5wEsA10b/MJA4+CM+6tyFdLHN110lS++CZX8VlKytEb+PpTQ2weqUmWhnmp3dTmBrT6hOSbxotv+
YIpgMuFakaN+eA51DsJQUKyZs86Gepps1ROsLk4IAXyilb/COMo4CpjaJCsuNVTdk39lw80cPQfG
5YP8n0MGWESunKoEtP39c4GiNU9rcQfrhPC88kfA6vsha6fZG2KJdsDfVR+7ROwI+KpuH8/Mo/0j
RdH+D++70dPUdJyhJVZUdu8CTdbD4dga/rNM8aAwhqUe/puzKQu1gIKXivve8aJgv/Arot2n/DO4
FQyNklm3KyTToz8qtchw8X9y6x+KVH/XYgwSkeT9cjDoa+Os7KtYqMl9L2OeWQz/7Lu2GgZHAyjb
YrtFwh9QMjpy0taEtBHRMV6iU+XCyA2KshLXnPQH37fFyrVP+SYNLRhTnv6/XAKTBI/X/7O9xK5h
930bfuaOlFJdLePcOzhllaK+/ydb7jyNWMe/YA493P3Ngwqx3EfAI16N6PSRka7kFb0u+hRk42Xr
4m3wVI1cvUom2WiQGhpMPS+878nDl77Sw4ewH9hWGonpfZ/88tlwnT4kw9hQOZeexnk0nv9ILF0b
ZpY5DWZT2JPSvrJ+EsYPUYLII07nVc1gBBOEchAuYpSuI11dlKzMug/uPUlwDxkkhrAkxQ6ShVB6
qNBB4gY6CEpwbIfqlJeKtdk4XwbX5V3j6OBD5hEIOi7g5OGFf5lhjO1rD3UZHSVhfok5ah/S3C+3
4sqkfYBgrDkPYxMChtVBOwH5MTsiDYhCQJ35Rly3pltA+zX7g9jYLsBq3rEUUy3j/SpKxdD/Zggm
6ZKdwiZd4068VKiU3oMid8Sg5bliEE42SwycwbH4ek6WkGDT1bPUMXNJcxLBxFHsqDo8weXm1jCM
9HbqUkMRBy4Cu+VVem25KgKIf8TT+Jjw6G1aGVL+EceP9Hiw6aoFFaK3l4ZgueQemSkS4G2IVFfF
iFivD/u6RbNLLJwyTNUbfB6FzU03RajZolVlTp8eCPoUGAuIx7VuU2MDGc7zos5R2ZAbcM/vTXRj
4dxb1l9ATssif5Gzu/NDczkC1e6LAEkq0LwGgl+cjplZPfTVAdarrWa8XG2oGGaqB6CzQ0HfbZpw
g5+Bjebk8QE/ulfBo12vd/Trnszbd+A2EhnXTs059DYGrbWyj+VVDsG3Y2FD1bn/dgI2gVnEQRob
Lvim06IIgVn4li7I9DYDT44wZmQgt6zD9z6NK9EnM0Iv9Y/BYL0ug+Fjlco4YdJzwt5nwF4ZpQUw
q2Ojlk2xLT6Z5n+Sk04xm2TdVkK95pOk1EHYpF3/Fde7u4k1xw11c/X59ooDyRX3Wd/w8a22mWhv
C1MHKf1iCSESTUNJUtIgGFIoQoAliDx7DiPG7pPXiKmhG9XAdRxyfPnEn6zBeZPctQ/OtRO+1SNO
mZInECgl+OlknggH2uXn+tWCYUD71SxAYMThmXB+gQDfl4E4Gf6wNcibz/QI4gw5rGTV2ynP6Hrb
3GmCTOgSayfYKkbOeiZpx8Enh3JMtv0YgTKlHcBd36vL3uY2x7jDs5VY2ueGW2h8sXDIpl2Fm4de
m8zP+y60UfjgqimdI/4cyr9txDVNXPHXa81t/fcV3QB1bLM+aT8KFmTEZjA2LKGXe12tDa5jgrAC
12TjZI0xLuJjJm2+OlNKasa5TXTYseDEn7xdV3aQc6mIQoWuLXn8W7lNG5Ob3lfvmArQ2zEHSBH7
fQ1nq/A3HauwD3sBqy8WfUgJBJ/Zt0au8XFq1O/4eW0EzzDZpEMrnkhYnxYfmKyAa1ZEs4ccZ4+J
N7/54JO/ZI2zQC/gv4wbodgG8XN+yinv5TNETIWAkzOlOh5ik048z3p1URE7U12q4mh7Or9F6vn4
nNdACmTNnkYePY8sOGraoDImeyep0spCHSKjkFC7Qz0VxtTsTiBK0/qYBmdLLlUdyFr/tN4HCXT4
gmQbU2/E/+37+zDjd/EYxSdcgbISNcDFlus4l38AxqtDDBv4rT+ndpmxjnoLo3XlAfXSEeNhST8T
LHIgNIXrvmJ5qVF+zUAVriz7pfiZrPP2SlJoYmh5hs6cAPd27fx7Xwdk4ydqvyI4n6Tk0UHiy3bw
krWLOBEDT+mKqJe7rkyW0JLAPgH1rlyoAotdWztuhV84LEIwV4ZJqTHOce+Jcb6sOlG4uuipnfoh
mXUL77rLdHyD4HKnEgiM3I3IeIqcszsLDTwKbWiHK/krniwP1r+1Mm2cMcOU6SBuMG78z5Mi8xRL
vnfTPwz2bl2yc127iC8P65Ek1BmbAHNLHcLemRbuVOdV6vf//gmf1wAAg3mSYVIAkD2qmASLUhON
aecKcy6txVeZButxgkPH1Gf7l02HnpaUAG9DbCiw38E93LUpV0Mf42QA1m8IYC8/bWNeN/BZC7xy
MzmY5f4khuNt7kCgKqNVwoogNFHVvUxlsI7/0IHPiXUaFqElzauDADPU7zwFIzpL5s0snRcvDh0D
JtQdcwtm1Rw8dv8RTEwP2xldAB9wKUwclOJ6ZzAZ0yEN3XSrTtVIw+AHBh6ecbUblPSSqO7OfWfJ
/GJoFtNLiBJ0suQTmpxebXqPqob4j2NHPLTbrIUxYeopECWc92y3bEr6Q8C58OEpMlsEbKBQL785
jNvO6IC8c5XSZ+wc+rAfUCAjNPL310SEmP1fMWfv1O5NQ6KhE8EowD/K/EWJ8KcyI0NJb16PI1WZ
rc9Tj3yDuq+rBxDzjrq2uDgVWVzJmsFVry0BChGw+nJX+gseUolf3tU0etqwM7juSpri7aE001aK
xhrCexjOLMkgc7o9YAZ/Mk3pdgPyYF+KpCAE3MjGaWR8tTuka52QpUaewOpVFjtbNGJRv+Bde/6m
lDTmDKogbwa9LhmtxEbUqbHKeCYKgbD8NYl7Y1UevmR0YLqR2DjWzEkGTgrDjLE8zw3k6rHdgNdT
A9YdUmIkDMa3ie2I816qqkbNDGuBtxQly0BspGmt9gfV0GkMiSEVkkm6dVUI+W8Ghn1P0n1JWOCR
tjyN3RMEK6ua7ReRXTefoMY3HCpYRdHBZP53RoCU7qm23xNU9N5QjDJieYOS73Cqf9KRSb/1+n9y
3pfk3U4uMZOaaSOIdal6dlMTavENIx/aL/ye/7Q41QN+Q2ShlF1UCQ36zZiN6ROx1itxagPFbCJn
y4e33pwuX7VYDypsjyCybe+2ciq0A199e/73iwXqkk5GDoZHPnYuyOmFBF8GPZWUToEGHKN6+rrN
3NMlke9JoCrJ9x72jjIj565LrQXIsyvvV6C1G5nJDsMQmb8Pv7Ml7qCAFS6tZa7c0yYm2rnd5CO5
VNniTuaaUPfigG1qY+IZLL/Q28XSz0lWC4Lw6FKSC77GmidtF4L7abxhcB0QTk0gN+wfo1Z/RIuU
dkAxufmuRNuj2+g5WZz9YQPA/etnDJUp0K3Ruqp6nZTrUfzTPGGbSRZ+exL4O2+6FGqkSBAs22x3
s5BS2xTnScy+wuD6URRfcUMStBfm5UaA1Z9U8EFbYrOvGobP7S0k1IYEeRrhg3wkhja1pJOyrsFp
yPq6Ciwy6kPRE/MPYtfs/yk9eo528vVgkxYmYFnA95o5FYKH0fRWChPrZ3sYOEeFodi84ZM2csvg
iofNMz6atzvocSi/Wu9AcItBP63eR0IVHHCNIttsWUP0p6l6Exk8hZuo0MyUl2NbSLfDmCO9iUNe
OHYUXowalymvuYbDulfGn8bqTz7aVQDNMsqoV9RsjmafNo4bxtn5pbPKnw0lGbmV7Cjoke7NcHkD
2ziyS3I7ALJfF2UkwsCdaIMgJQO7jDceXDk+Kj7k1SHe8gi13W828LY4fILGY+a2akMuTLJ31Boh
KCYqzPOxgaJiR/E/lFYq2ul60uCgx9aCbh8jEbCAUIVDXMvuhQKiZfYaNrC6N6odabY3qaqI2qsJ
/ONy0EeHPMsi0m8oSzY7SIwXaDVVBzxdu9ItYK/UFs7zmnvpzsQyjEYtbleSJFQqnmHz3IpCB8Yy
dhzFZrWwQJkzYI4NPUKo7az/460IrlE3RWYtaTvd5QQw1F1gtNwXUGlAHA7a/bM/8/3WaSSBLFWq
V0ZcC6ANdg0AO/mIxSOq0ydNZWNT7awAutVA8f9j/OonqwPjITiZKDZqsa0ZP5lnPWedJ8+Ni6+o
u685spjTjprSRRiWFnF28/rwUumDqErIHUIV4+stEnQQkTttjBxa9u+9w88qidcdzoKRn5Kr7d85
iq+GkyQl0KfCDoW8g7rCx2hC2ySCvaQbSq2gMiM07F46ig4kJ6UDY71KZmQSleYzGNK3OCXNAVni
kjdFaqGuBZiWtE8m8d0fKTt3gli6Pw+6J7C8lmSO9jni502WoFCjYYokPydpBazR7YXPWCx7Blrn
C1wnbT3Yc2j9+1R3Jr3pGUDaS6+/DWVv0fcmvCM0b/WlvABxdpyJy0P3KuAm8wPgJkr+jskGtXqf
hC4FJaU5q0eOOvN6dKYS5Arund4UEqeqQb3NacdpAVUJDqHv4jrpkEp0MgiHl7fWdDl+D/7DJidp
D7XtSsDUmmoaKp6oXOtnL2xJJVQH0nbgAOg0uPWYdoq9+GKoUXJ1FpES8ewRRLisr+ptYMRgf1/I
m58tIwPQuqqpVI0YIy4JvM+WdYudL66Q8qU7qpdlfQ11vfsm+LIoPOmDpEp7C7JR7XWQbp5wSFN5
azvYVVWiJ93mvztPVg1/N7v6EeK+zygNXcwSZuWd98mvoDxHuc31LvVQQSfPalRGSTuyjfhFifIJ
Id2D/idMtG63E7WHRGc7jKgUbb9J8cuB9nKqIHLmherKjXdy/lbQS+7ow3kFxdNB2TSv2kjbhY1d
x+GSLkDvmdQELMdf81a/QA8M9uHkpvEe1uLIYSH+pHi16cIfMt5Zl+eHCN0nJZVsUPKky3pmSNZ3
f0o8g16iDHg+Zfnn/pPD9HzsuNOtCCHXZsdmU52MUSZEvR1ME+ws0GgUstnkpy5XGSTLuLPPeYTs
8uygoJ3a0MhfBmFl4qHsyGnFZj1f6Gmk7XrTg6ZRCjeum2hsLv0/aM2U+80mcxpF070I8h2PxDj4
Wvl/s+aS/7QIpp9wak9ED5DFv+u6FJ3+Rx462rEdSzv7MN41szCAIECbpbwE3QrQFjvqyfDtDj3U
zNdt5X+WTngTyDihmcSmqkkj52rhQsFYvd/zSs8V005P05B6ovw1uVMh2hUFkmyiq/o96d6Hxbef
3wNbpDrhxGOQLbXxLZcfN+YhyzgAP4P0Rza3465CIt5j6n+dUPh8vUWvTaqjt21RZHoBc0aNs9RU
5fRmjfASQ/r9kYzDJ4H/4d3JjdnRao11HkrGPO9KNyKhh9G0R6KLpn98ZTa2pRf6vvMjxHln59+B
XwxKkVLSRvsgC6/KCh4Fb/I64/v8G0+wC2EWK8i57F7r6ZpGpLb6Ggvc+VvxDi5hcjg8igiObg5e
lRcKih6PYyIFU7K/HLRYXdC+R9eognlI2zhCxyhFOyE4SUfXw02BTWyDLqyidnA5i+3Ry0jmcWEs
kAxQNlLtLGJo9Xwj2de2nwZ9MrVzWYoydW7XMwJqYO2bVpKAB5qAAtPtFz7Oh0RoVnCkdNsR04jt
jwoyV4nNQk8HkkR/Q9It1f0AmZhWecmG1fZWwJ7WeY2bKpo9E2fCOvzxgUJPwq+06dkJ+y6kWRmg
5bIMHigz6t3aQWnITUDpWWcTLMTcbND3CPRYzRH3svaXrA1iuE03CgUGJRbqFGF9hcyqRkeLA/c/
VSwtvKCgX/OfiuV8qfBgteKT19whdgGTMPx0dAQlxYTxAGvGE+Ma15V3rcceEKE5KorfQro1ft9e
zvISUPeA+1pBPpi6aE3LO9jCBwFNL1tHB9u2JUva3UhUsTTRWzkDZAdcSmobOIq+9xH+N5Gi+Luq
I5WE6AIOjHk5POMNxRiUBFrbddMo/DeJM8KRweS5zm+Ztughq7uyukR28bHL7bB2pFw28UjPnjBO
i6yjNKR3EHFCV+TJvjSgKTQ3lnky/gS+8jai9MIdX0jBNWv2y0xSL2LZwgbwo8RxHo7aTbsT/C2y
dkQ5bwRgwKJrsjOYHv8gbbAGOx8oIVH2hlBtxuslPC8Qhhk+SNfNQYvdRfoN7NC8t+5ZYfddTEqZ
E6qf19JpQRvfuXYHBOIoS/ojanaWgEUSvS+4iKfSsGPQJknIyM+HMUX+BB1/rtaRlFhw5rDxr8fa
G4iAAsqOmafK5s+C/IRynq2qhIgj/tY77no57mpRaN9lDm0yshNmlKu2mpvo9Qbk6qqgYZtNvZs0
hNiDpcMw9BhrykIYl9RSdxsPKe7AWqjIghPS2HkT0HLC+XQ9qWK7uHDzRYSG+KJR7ysr+LhNJO/v
eS13zG/4DwsJVbiDuXeZZrOyXdfm8uXgZ/Ji6BUkuxaZYtnkX1n4fmFyB3N/bQAK3k1bqKOLAARW
DRJGtqe4MHETtePLODswR2A0wZEa54ORi87gsJHBJn09AGp+WLjvBAb2j3Hi5g/eVk9YO4krx65q
xppwPmF7K4UEwdsOKlimXPdJhViRDIZudoSI+LZnDcz21OUSIfIIUMTrmtdeFV28BEXxoTl2M61b
Iv/bemewmDvC04YANPOdGatWmVDE0ltjaoDo12/rvnhohUIMDGUyChI9f9UX9RwIpJnjPAPEA+RH
wfZgJr3TKmd9HbV5PwXqOwk1qwDiAf7lujNHu0AVk2mQmat4hx10GcN8ztK6jbEpdiqX/DohYxv7
VUM973zs/RHKZJxtCSrqnROCbqhRNgbCqDaQh2xJ2D0JuVAcUO9akZ55MqUPz1t9sVg+WsYQQXMD
NlXEKroDD6gQ6pdX9TbTC4/nM8SzpOS5Mtc7bjhRu9ZJiQu4zsnpAK9oRUo1JAtxqSh+6Z1ubGkn
21MiA6SIzQLIpfiNCNmSFrR03XJQz5hVtzquhYKRpkzacOGv2QWPGFVUvT+WPaENzxnFokYYa5Kq
xr7Lrn99F3CQD8rryg6IDCsy4M6LtHYZLPStXxtkpiW6kjYPkp3OISdoP6Rm46eDxvR7iswsEz01
yNL3tGXwy85tYgt+SB/tC1lk48kRlDMLDbmR7roJzsKUcWHwMB+32JiTSYWD8nzfTeue9HQMSTHt
ALQHXbmLQKgSbQjvAU29TJuW2RxdFK0knrnwPYLrNekuk1oBq38QyZl4FV2fuG61Qc+sy+j4pqIn
zwA9Vh2RQdr1TOVrWy2K1oHUHOaShrFvrjApcmmAg2AbcVAk4ZWiZT7acmejlmGL8v5JeZdqrMa8
lDBis+z9w3gOnSU8nI/GQjRaAyUrhUruyhXtvWpjig3NBrHl1f1m9Cqz1KgVWBVBrbaFcXzE7M4N
ITPldB+20WGmuPs4zCwm3SP2bepqS20TMziwrQd/g/jEgKmZpZiAF0eZ1JYmYZwroENyt/XfWK2H
VYU3dyufmMdDWarHHgCNXi/ns1uMdXN0rGEGMxIO6MaXN8UyR4NrXDIVB/SdvHdweCNedQoHDk07
fHg8Ub+4Q0zc4JtV2fsIzsVPsHDpmtGqp/fLnt2PQ/tttdsxOFf/tMGB1I+eSq0nCyGiPbuH9fVP
4i9crI2vxaS64MucK8IO9aac1oFTEGsKpoJQtj3hZDqcfYXxfLTRumqKhKqfOqTyA0QC47+GYRu3
nzk5rsFnZUN/qssm0Ffl08R1G+AoGKpzwHNwHCWh19R3m2HOPEGuWi5gM94DSfvW4nLSCIneOt3R
Zs8A8si37yjmm4pDrKxyfw7Y/B+5h2HpVmFwpqh6wYKdCvFJFtcxsu7lidaCvDs3uDc6bOVPr5QR
pHdJZprS3XpilMjnmckm/U4H05iAe9t0qYnq9txqZgd0hyWds9VH4BWxla1i4ql3MVDAVgJvQaFS
IWAi2JJnrkwSBgLdBEtY9t90zZdBvUuhnw9A9o2VyGICgwSERAvnbydRYWko80IR8mjpGREfAHyh
Q8G5vp67ve95b6beyZGvIO5HTizzS9ayr2NCA+xL++JinOh1RQrdKlnWcSt9JiRJ55m21+/fpdRn
qvAiQ/2es5ebo01Wq5yk4JDdXaRrr709p+JI6Kp25umDMyvsQPdRnYbXA/5ZB3Kyj92TmA9tW96K
wVoGfJiY9bOH6zcJLRzokwvd8WNSc+f2Ux9PvrFjTmg+wMEgFEdNh+dnjW0uw8xJi1qYuNaq0D8j
CqDITJZtOBMgVo0LoQj+RH/13XvORIJbp6QC+fYHBbBZets7NKNCBCKcy7zyAX1nULU43oqunMRj
oC6pYnlvozKSlIxYVYv74Y44fV/Gi7LVO3+rytGlwNvv3ILzT57XvTkTiUJc4obbiRt5BZENgSXH
HOhid2W7VMhbNTik/RBjdRGgMq/kXtcOd2SDijQ161aa9+s1E68lkK4GYMmv1mGjDhYIMEZ1mHtd
oJeiD6Wow4V4QLS3Peo5fJ0o87G5UPZ51W2csJfvT76ex3w+Kp13x+3C0wDddSia4xsJ5Jc3drYL
ruN7A2ae4/cDByswoHCggfSuog2x8ETX9aan5iLdxW8ppX6pILQxauQ0FyhO90ZfoJI9pjxtXzLT
iNI22qTUqdCbJm+Gzh3v6CbFdRwWYhFED1f20Fav1RkgpH+Ll0Y5PTt/LrnVFLhEXa3BBACmUdtW
wDN0mXhj1uDYR+tPQmx8RuS+CN+GgmWDZS2xuTTAWwECyH0Rnvuzx0ik03Q4ovsI2SL1OXOhNPji
W7TNbOtjOz4fiJ3QZnFUiR/ehfB5PRNONaFY+jBCWaUI5UtzQuWxn05r9qvl1oO1xgLZ7RHN7p3+
vOXgYvRb4tfDiZ1D544nLlFTiGTQCyxE2YSk3JUGA6cvWGGiE5kfqdDRJzWnkzWz+xA6VNgfbZ3B
PfJm0wjE68lQVuOQ/j+ncfhrkN4X2Ar8do7c/lwGRT2euL4T/WInFtQTynq4v0h+v0pS8WkT/rY5
HrvJbWTCEYz4r9xgbYg65EX0x6DSBCG5SJx/WJhMj5NYadSL0H9sjGKiz/e73IN7tD50PVjwmQq2
pPPjFUZp10cELA+vg7LOsmFWHcPdf2saMIox8Sgcny/M5Uumtu6Yp8s+rxBCoiNU0ziW5yFUBWVe
KQzxiOIOW8W6Z7vXsA8kHsQxXIy4ePW4ZSm+hdUn4Uoq5J2AU9L/k5rv+THtf+uNS+K6FUm28eDG
iwv2EOQBQCtbsfzENZseVDw1SJqhfK+pLUbYGM4vO3Kcz1pXAKed524ncknWguBJQcmF0xq+WR2w
UAqKfwmgsPBA27sgCxMFbWbkmDCN3HsbfI+ALforqxf4SvWX4g3kIYjsSzQna+FkxScaEwWQYcIs
repUmgDZ/xWBFAcDFw6ESDWLwa6tnCrblIA0oPc4GGES93RmLcEzqL3BJH9CJ2Xs46hmfwtcWbxO
rYhoJwQ6Yh3PEMbpG49iuCyLtcHacSMhYGV0UAkbY8NGgmqXphfZvUQcJD0+qpHKxY1TEatxeoKj
epFm8TQCPSXp0gTwL7XsyNBzJ1g8aDKWGzs9no7riUpxz2MeWG6JfP3g7g42XRXw4zDVVEhNSTUM
sGwMZ+j1eFhLW1+gAv7RLAW/CRPOg0mIk9lS3vbey0UwTy99o5vWVSNqOzQ3BvMrkJ5AFbjk7r65
D22mmMha7XR02RVazWfrn8FAf+mBucvtShBQQhiLL26ZFytdgvarthwfbga6mJ12F+jjLwzyMUi2
Bd09WWzOZVdi3QkwFrhU3642VOljFVjiEKlRfHvi5k4wEWSO1veJBCA5dTBCHfWOISCdJV+xl/83
6nVaMOUfAmqtZrVymuAqQBlzQfVgfkK/kLFL0pmhILH3gziXqnEI1wO+OP+RGYO7HUFi5J6ACH8E
XJjQ1AyBglYrAjo9FaAVCXgFIVXbLviwJkVyzBVkbLeEV4jGwR0zpmNx59qDBCRW6xrRyw27jdu6
lDlXMROYat2yefCxt9N68s5R1Is+Dx0uSlV2QY/2wV4a9hUj5RSnevExP9DlHepnCV9DJCCe+YR5
KBsZaaQlW6LIHGjvPIkJVDSmI+2RMMjJWZEcMpWiIsZ30JAdd5cwzTmbRS8M4OytnI5YF0Mg+3DI
DE126NLtre6O4Q5UmNlBDr4RzbYKR5v5EcjZ1Ter+BSVhtoHoKUGPUGeOr4WQ692Q1hOMSUksZ3Q
Xk7eCQJEp/w/dyubT5fx2sk73MZ5M2D6dYES5Sfk2K9k27As7ZMYUnpPnjKSQyXsKCG+YRkzdVMJ
YQXOPL2rZE+PmEObntJLjCMJqRwdsjbftH3e4vxdfDjCbGvpF9lX2sA7NvtNfRpXunps4cXudIk6
yOOqVW3X+bURZvIF/D0zYKg++jevZ9lv1TRXOHf4TM/Yz1BwqoYYN0bEytrxquFTF1tjtkiw3Xxs
cIN9/QcN6eSwH2q1WiBNiFnigo3rMliBuMSNmjv1efignezo9L/WJUwK/mhYeY5DPd5XZPT61p8n
lxgN6MVw8Xe9/ZaMJnJWZUg90bkmna3Q0hvXDEaPWOCQp45yKGPVicxTrVXp4KKKzA2KtiDQtIZt
fQExIn3puoAHaR0kSWjzKEC6A3CXH2fM8AK3B8vKqoEPSpifaZWQ8TSK4n4qaeel3aa2hPyhsZ0E
GnG6wBkw3JxOiuefacVp2XiYqGuyvakmQ33CyumWbX+07FYfMiWwPzAe0wLHvtOOvssPW8zsBScC
mf5HWGVrk+yXPqTX8cnb3g4kL+8X1ZjZsdl6Ris95+TIxaRVpQVhR/dK9nUa7B2r08uLnVdNKSVC
4d3Qsj9+pKYQnZmYv2Kldz4asjLjyUJnXnsOp7Fco6Bqu127kRYvjrCYD+ubQzd/YaFTs0qyaEI0
jNYPxxE4b9AUgxH/g9nHnYSfjNYCMb13Z22r1eXJ4Z/bdUqA/hlrkWgl/bHxtyr52B17AoE5T1J8
r8uJavXA3WXR7FVSGdjmWvTbI2Txx1iWh25ayN4q+Ray4rO3WRrnV++KEKW4809Sv+3JSu8PmKRq
c/rN3fGZ3Cry5bsNN4a0RqMPrZ8cgMXVN7h5Xybq18L48+6bJbc5oJrT/WvoHXYMjUW6mf7O7vXq
5w5ddkRmVhTRvHlnWlPWM3d7MDY3l+BF+E+VYG5TNEZqykjq7bRCgE4TY3ye4PZbSupyCuD825Gc
sN3g864+YXeN9s8QswINUdV6OW694TpXH77VH1GV6EkLPfUQ3kbT1vvtCwEeXUrXejdk/IChV1TE
T2gKpAUENrFLYKc+Bx6c0J4zV+8c9KVW4IL3ULtjxssxxscUNB1hEqlwwJTZxvcz6bkmzK6s67Hf
zeRpfiKKnOJhDfOBQr5+nudix0/owq8NFc9C4RWeZdIZQY8OA3lUx4UT5uJCpWTH9R/mBrxneTZj
ZwbMns+TZhHRVbmMWnT9GQjVF4Yz4K9eUxBeOMpaKu1UFcxicOEH2lDF1mYpbqkZz1NItI9m6dqO
Li4JcXSBzEGV3k8vGDtFzskDkw5tdPY7Max+GHw6CcJKu7QmcImU5IdCNFOoSrVpMYJIS82uHkxb
NLJ7ksnz5SJiniJLwJj9pVHHrId7+WAzycGrSVUm6Nw16weD2Rk1dmcMtV4PK+GZcGSIHMgFHIFH
UYhqbrQeSglyklvZQf16o7uJDa8NAG+iQQnpiyTdgDN4rHSSKevBRQD38iZoXRyfRQhUHDeizNiK
QCIDnFH9eWjCLj0FugjN1aFZ1rczsjyjPOruE+QoIB5DxP2tvzti0KSy5unLheuSTElKEJzNHhhq
DCqIEpE4R4SdPjqW1UjbYJjnp8ZhJbdA6q+fXTXoMvBG7nd89XvGnTpL3sQjLftVTVEm5+JUPhwZ
oVzDm2aKjOFzXvIa2m5cRHD2TkLszwJECpW73wqM4DH91Ztp+FsM4GTDdxNGa2R380tlXp2G1cI/
fr+EYpw2Iocde3HmLx8rsaoeWGSWUHQZE91CoGtbFmeyy9pQDInY6UCeB1Z8wFnj9uolvIhTZlLa
/DjBmo5KWXwlxKaBaIjGLNMi8o2Vl1+y9rmHi+YKHBm+42sIZ3OgFk38h0G35eaijvHcxmsB/Fb2
Wjo4PF3m6AQOUy4o2GfIDK8aRPiYY+CcIpyinW1DVBz6Y7Gfv+jvAdo1fj9tIuddTwo9Ep4SBSRv
b7bG0SGqBi3YvZg2eP2Ee77fLvzbxwdamerdRanqlQXlsSbAw6LG4XbUkwHR9U6y1yDl9AwEBQ8q
PucP44aztAN5iboere3jrqq+pOLqhazDrS1cTTGAK1E9xoyvrgWyQav/oqnZ1xkTN6FZ0GloHd8G
sV5/2ZnZPq9MZH2bLvJHhCv8kcwLtmxUl8Osf/ACtq+Vc/C3D5MEjwFxiPOxW6Ikjuh0SeOpncea
AwdePfLg6edCYaysL6x6ZUAMncdUjwMmnPmU/chZ5RNzMsgR/cR/FkBXviunWwYFSBK2FArPGSDm
etTjJYxN47+ZAYCZ8Ben+Djl4h4JlQCThX2mR3J0lEOkTltonUf/MXdqrVH6XJZfIH8NsTDDnjps
V5MWeDNoAc0p62rF8djvbjo2rOY//vhsu4LRbU8/sajGeqdGbAyVGYxBVzVJ4cTmecrcBnUH3HpQ
NioNplr0LZwL3MEaMLFY1JTI871AYfFJadXGkSum68p61VAYOmqAqwLeySjncD41/ocVH9M8IUtK
azpT9x2lDDUFS7hMeZMHE8qvC2fvGPpCCmL10wUbAl9Mly1OMiP01v0a4EKzTuXWk82gfdCM1aQk
5PTcU1MoVSQ6lC+HVxzn2w6yzUm8jYt6kLE/hVsy8zMj5Is9h3ltFDk+XmKZoQtr9m4BdyhdmWCb
iYTHFddxSrnlkBqJvh3+fJ90kTmm6tx3+4LZP5DMSZzRLzlkouUT2J6oCEjbst4SLo1lA+QWq64z
5xm2j0A51KE77hZ6UxiRdmRgLAT3NU/+K2GRj1c8DDD3T05Ud8YlcouzjrCeh1nf8Y4COfAc4bla
O73jIcCiN0CscPTrBawhwsFITm72zOYyyNChFKa36TqKTh2/UJHNEz1AU4YDLcqRS/L5NxihqQQu
z6onu0WCkg9uK4ZHc17BEx6Dp2hUAj4prXDFpNNzBEToMAP/jrNVkQYpYcc68DU2XNj/LAqhuk/8
GWhj6ZjwTQkTFQaXpN5w8zdfPXLVAuIFWKTBZFgu8sctNFpm58ROQrkaibQyCOoF3HdAx5IMX80n
O10yGowLG3dlT/SVohb8fLR9TsyZA5KfPUVgmumHG94qrtJrAb/KBjExF6PVp9TlQ+PHJkt5CmIf
w9feMkL5JTCu4yedeSfjU3YaWcNYZS9oPoeSCswihcuE78gxfKWoUK+B0L9yjXNIR9/qDqtEQ4Af
SQ8CIXKdJnNtyTH/0ykzA7WL2DY8ghTfsAF1KK3a6FEdmLHY706/dr0BiV7i+xPMD4u4+jEf4FrB
x8eCTHYBKqlRoDDIl8lUfiESbJ6qK9ngwhrgYwdrq60O3bzkSeE/ig0aqAsCYaiePly44B44D/3u
cX/GX3Kqgr88eOZSstS+c81DanYhZwT1CjLqgkuPFicL8M4hxcXrbV9oTSl1hQ1XdGMo4o38C5C9
OYNLjp6USTMucv9SPyVsltJtstpzV23DcJ5WSG8SZfR299rnzhjMfMVTyeNJNlVL/dtlIH4lSJrL
jNATScnVvSowbNtELkY7qeoum4XgY3aEjwHrw+xJrY7ETMRDti9r/TIIhcdsYAUGIk7UhQkxhNkp
i+Qd+T/FAlIX1mUL4W/R71D31OgaP0Ki+ugEVmtjTNmkdvMbXtrjY0UVXocGP21s9rDFhyAcFHvQ
HqT7eAXbo0xwqTm+LDsilHTKRKk3jsRfr27oOnEJL8uQuDSkhOZhjK1hEFtuKyALz3vkqiS/gXA2
7vi7JeOfrgcB0ISh9Zs71fgdQlW5CGKR21wjXkdskCIB0cx1vNhjBRgB/cJowexnjGUckRG50FKU
QNlCOMbb0bh5E/NzBiZQA5aoskSSTPIivqPn7NtHUdVicSVyhT/JcwH7j6X8Q4iiU5azgZhNiCfY
voe+BpQiun3Zq6cLqidMCoJEMXyIVaQR5n5HbvCNb2E5yR6YS2c3MhYEJgPVwMh4Fb0KzJyY4SAX
6EjP/sA036OlAV7rd168aHlBOidRw7h7uDGUdA3SM8lWh7DUNGRpa/19DuYDkQ8rG8LQtrbN/uu/
Je4L/v40dZRMh6TLCZshaJEWUFK1TlGpmn5mEqJmoQCw0yzthcPmPfK1ze+yAAhyNvc4QFnI3mcG
H8MMhPD0FH/qF3jDY3Phd+W3spFl+35s8kc5p4MMXV4JWcSPo+tEuno3nC5DAng9/nK7CMlsYCTS
ToHoDlAsvwjm38XN2UW3Mj/eCHA1Se/THLzVfNtG/WvLABZtCwtyuJXr4ilMGr99gU5f+hyyef/y
Ec0y0AuOU9YZbXLNXwzR+nTtu95DjUO7uWI7tjXRm5/NecvEsGktyXeZe+g61meQV2vtJpPDFXmv
IQovydcbT4gk/SX/i1jCCdL/cjtarOcKAP91C9RyMtQCQ9C+iUv3bk0/HW+D1QYlQK9T9uc4dCuL
WlQWcbpyUAOmllSn7cHQIO9g186NwAnvqi1j/FGM8Ce7p1alHhHJZi26w9yLVJUKHh643WcVq8GK
tl3rjLQ4hltLJEl6vVAur9wnRPdNzQzk1QddOC39f/T/ri/wE6+tP6e3yjbJtGDS01MSLJTTi9qD
ulwX4k6yIpWzJfoyz5oliX1nID/AIcbd2KVvnLdNcy2+rqPzIb6b7T0JIFE4Bl2BRFpNHfEtxT6U
/JbcLlRgi323czyBWfE/MubU+q3ChNJC2mKmAZ/u8/1JjDv5cqKGRILSE+itIIIMojbrlDZ/KrR+
JVWXko+V6ez2cr+WfTSbZx1CWGCF1woEE3HA8ItuWqm79xi5AAPQu8JGUA06aKWnwWtQz4Vi1SmK
InQ9hRkDWkkSwFACgCoCZ+P57LIAmDwGs9g+mxE5eBJH8H6F3aJWpobjV2ogZibA8haluOLXvCd7
8ntaCaCbDs0Dg4ZiKS59fdzUsMB06G8uCHwdxlgWKVdl0RTdrOkxormxlEivGDouBz6u8EEXii7Z
rCEoK/GdUackDH7pEcW2eQYOMvCabsVKNVAxRNmEUg9vkVpz9zLjb2Oq0UgkB4yVBQqJPq8jnJ8C
JX0fbTkvq2wneBMJds983EQHYL6Pb/qa4cGoeXi1YaKRbEcoqC1kJ0w79E50Vzi6Q5MgLJPuYsfk
uiUsIAxPbF7f2oy9SOpWP12enuRqQ/CwYL6hdj0hXljbEl/DHpqxyrEeYNzYdgciub734Lk8ZwYV
5L0dr4AV4NuRIqN0niQhiKU7+lQGSL82ivaTRP9u2bhU646NitMiHMJo+NI8jI722jptIEa10nK0
7xq531jVl4LdhMsx7mGe58SC7MBXbDICR7tcC2OGL1lzDXa8PuyFc/PXURvr4iRnB5Y6KK65bwEQ
ZraBC8s0EiEEnQ++4Ezl+LrV5I6jqo9uqkYwiJsttIdA8KXUaGdBXo7Q06FgZ3DZQg7dzrsNe9O5
0X37JDvHxEtcwp7CrWrTHuO0FlAy8X7UaKpXnmXVwd/7k2CpW5AKJYPY+a//RYC2zXETqDijbayP
aDvjirt4fHOnISw8srODzNoq29uqaVZq5sT+B3I81Fo3jgymGYRWq/ahCdDsws8SGSrxqV0ubeIx
qoGzPuzVHBaCLx04jO5vYBaS+Jh9l3EqHJwoLQb3RT23skmpeUJXBtj4KEE8t7w0dOXBhwCLm7wW
XPThgfnR6Sc/ADbVa6I9iqBoiKcX0wPawFBd9/j5y4ty8WTyq2abaAnnrrfOdzJfo2aojsQQde1+
wx5Cw59ExctYqWPpW3K3VPwW+JzBG9+fWmXbq0dp9N0fQOutu+Rvvq6sFqdpQgBXvAP9xCLbrqsn
ZIwLZPXjlPnxsZeMLPALiif/e83tzdfG0RPwsTva5n3hY+yHgDiCkxSzWxTfU/9lEyaiSh+ecFE+
dqQm0z2aeof4TkBXT67YhmJyGQoDfrahlIu0pj1Axt8064N+rpuqknCZJfFyxDOO1i5OB2d1THt/
YaABZIJ80/iEy52dTgXa9vDg/cl9QQh4Jcz5WXJOPocogWaLNzivvQhKD2MhHBdwiZSpw4nw+qqo
kPPVmaMiwI3WUT4a0Bf6pE0cHEsTMvS5ak6FqqCLr1CQ2wFtVJtw8/Obe9SHLaQY7Vit7r+A7aqK
+ZoiTrmOi+gBFq9xiPFiWORLGe6sbGGXrP4JyFIeLA1D12uCAh/eH/gqPfoQDjQmvK0TGpKAc61s
NKV0C03d0TgSNVJUKGV9P6+xbsZc4RoplYfO5RvBEGReD5nGZz1gfnqhpYiGcXY3NEOYOt4PIJu1
SqYPTrHFKxodCmssXPjcdKKX4htJjMwew176trZBgHxVvrdUWOIUZ1eTDjKiH+T+W1hdX1QG4E8p
f4PCoy9JBGP9Aew2Qx8fDGmtUhYTpifmEpQNCYQzuthiTFB+w9SRiyFLiszP5+0qpLmU0aq19bnb
eLdcJKzLgYaBQlJ+MXitic5UcN6enbKlvqpSHA3e4oTRVxY1phYaFU9PWXE7WCLkcHkF9ijx3eZU
3KB09V5y+WMWl++QfpMmWK++B3Kmv6ZvnpoK/MXOMRJWoSnkbXKN3GjGOcH9g0bVgr2kxi/i7zS8
ETXICs/Xz3QqFGNv3JSwPUSzVfBncXMDq/PUiYE2hsP8wWvRPrBk9PmEbI8AF7IpMebuDL33bl8m
bMs2MT0pZnGU9at1+5z6JtHVl+eoFOFW1h03Wy0E4PnUbtjmMSmuWBb6ZohLfD2P6XxBs+MkjEAl
VuaFHH2uCneGZ338EVdE47bUOmNrXPwyE5TPAiKqnOfLtJLfRyW1a2DMbI9Xl5cFM1roXyux2ZDl
xAIvnmcINoFnmqfu0uAZH3YgU1Tv6j1hoGi3NuECHfNi2MDyCL36WiojAQflL7raeZk6ec41sDaY
9+93qGmoiDLAIVDhdYwUsfuzw9BqvQRuJgZDrt6z8tVoEdtulR1Ukb0WABqf6vWgOyezMc/o+sKq
Lm6RKAFcKnCFAMYmyTms6yJnilUJ5WQJlhBD0bmdX2YipJxhz5RqTMJJn3Fv+PW1D31pFIGdjve9
JkcLYCz55QS2BAOj8gSm0nwy07MyxvZ0wz2Kc9BMaADLGMeCi5qj6ne3TLHRNzHn6QC7ootG1bE2
fuNBibsIOzYYwiftJBGAOaZ6LwPTtzEsuI+OPPpu13ysTYulHV8cC6iKI2cAKtCg/k3dLzD2O2kj
rX9728oXltTn62LmCA3wZh4E0oMcr7TEP4JvcK5i9lpa1kOxwjaNVQD3xKqbDoE87cFXYlQpYIJN
DwJB/yBdzKppDlgX+8Rj0nypDvAqBq6RoSM1zwHBBYMV5V8W1ARRKPhmZVXdvUTN53lkcYId68Cy
v7uS++e9hnE1IcZ22cXlpWNEamimdmcQvmay2loQnRuJwiatG3qC/IgB3wYNnf2z56MmaoDW8NnL
FpMkmE2ZIUPnDUIVEWA4BQdZrUN8c+EyQpT2iVdY03YJAAe32n1LfgUxwQfYHQqWc5ylVZLACa1T
p9SC9HikvbNn0fuEGg7yvvSECqnkeP/PqnINlVbiSxZ8WEyqdETGBdQKRoMmmAL9+w8PIaJxGU+P
0djatUBrFaXDNGH+g0HQ/W6NTIhImQ6pKLH7a6RMvX2nEFbE4amOl8zoFrTlFbBPbBlFULQLCLtR
b88q569r+4vfS8tz+KxuKry5ma78yL9alOrzgkOB5FGvhbM+wrnJGcNrQw+h8g2uwwe+y5nmRVm6
BdLh/AI2j9rSKqiKn3un7OCfGkIOYXrsLbj1jUYxNnW1RNokwbTPJGf3NcgNOyH+B27bWu3H4pU7
x5DL6AtkKZDhzBu9diT1dstF/MA9W9Xo/qPkBfSJQiO6CfyUoajKWyfy5DHR0CnqS+H1XPFdGVLW
D5WSurXgzWixQGfBuN8ChS52sGsLk4doWAfQKxk4K9dpe6WhUOBWA2aNJJ3ZTZtUy4OpKXbJhwg1
KhF7kiz3OMFgFFQMr1z2fWYZWDnCIqJFsQwoSYGaRzWneIluv5FjevUD4ItXu66RT3OfcquFcIIT
9XTRNtFlVrFSKmGV6J8ONNdwlLk64+6zHCj+NBdqQ+QuB/m6JXpIdKWje6+eloCclz+Cug8oKCH8
KehhjchgjNPpImM9n3GtLueDKMXHWDhZGW0XH0UNe8mLGHL/laKoX9ThLUH2kkTwsUmynqE9SXyc
ZvdJGMVFgorNiPYXsfxcNAY7y6VN9b467+n6utp3ZxkTahtFThtb9FkoWKoz6FsNS4fOsY2XZWlu
WzS/Mri5Xg8j28M47MGpu36g1pguJu9PGXN7DiHT06uRXr+2KytiZ01vMyGbN8wC9PXT8zhT+aZG
G6/lPQoIGpPv34foun9ZsQwiYB714knZJt9MYTjvdwyMAFaoq2eAudDVpBpFl3RTdYoHK37IOSS8
1dgwt+4jkQsa9lh6q+NCQIYy/9qF85mklSnGhu7/HMVyrlUujiHIUPOj+fmO/ilA8P8wd68UzFAb
U+ub4eh5cw04y3tumSxoAOvJgnGHZ/A+hKcWqHMpWwFAlI36FlYK2Ach0atpSSmOsG6uQkfFmchW
r6V+F/sDwhBJMJcptS1aW3rAwhAb8VI1p+6AeI7Z5c5iiUL19NxjSV6Y8TzqfJZ7J9CZkNSYZKFv
ZavfLoUDYmufQjMwqCajseaYqq3k8GA8ZElT8XyhX85GAyR7oBFxrF9SJ98m6oODOaMbb5EQrYZ8
Rf0nYweyEL7tkIuAPZbX4FTiy7ZvcdBo9gHo/vXTXcmYWyaQOPQePbwWkSvNGNs9QKtTw04lzBbb
HSJqI8+hd106J/Dp5z8Bse4RYzER83ROh/vVmrLJdhyBARn2y1RXBlrVneUQvolPkwAKyop1ykmo
TL490w3gnhM8fGx/Ot8cVeHvkfWArXODitY8Tl7dbxWP3dLlChOQuMtDeO+LXsif81Y0/G/OhrdD
Qew0q9je7TZO8C1QDHN+xqGmgvtW4Pv5aS+9jOyZ92jedZb7kdgL/hOBU4ZoS6RqgoD1mf0SMwzo
qJwakEaOWS7FWH+miuC0dprd+Fj5ChIgpmUFOtjFfqfrK+O4dq8+HfUy2uDDRza1HZ7tKWB2RwuO
lN1Z1JQaH3Yym5HRg8Q5wke5VuwMLWtrG25FKVwZ+vTeYeFBpkMf+irs4MebVAKyKZCf2RdNF0gu
AxrPDztjp24EqQRkY+BgVJor7hriFaII8QdXdCRf0Xt7hnWjWc6IT8eqFip+veOxg2nxNCvOngU5
Llb2ANVVBR7f9LADVxJzkpDTeHoZnrsvvniXnQnRMZP7LdBkXGbnOa+6fJKBSHHBwvNGp+nPc8ni
H2St/gLDBe/r+uaGFR+z91yPc48qvhRRweWF+Ul3el5ePeoLl7vqfRWfph6G+LD0y0Kljow50GnU
2UXepfkAnKq54ZSLT15LCXMbW9Lmn7C747qSQkVqC5QP4YHKYI6+B/QMR1/1xbCPKXqB0gsaGLmb
KxQGcwzDq86i+uc1tLEGROXC5RcZ7HjDELLZToXaN16pldVs7lcHRIPi15p6uDCXUdhI8TQ8Byeg
5gUDJ8vFg15mc2ksGXvhXwfLcoiJn05n+kgSn5r9lYr/i7F5+xz0m/B4rIXRkVqUc/J6lAnossEg
nnekCYb1qdA5yceON8rgVVmJJ8Tm5+np1EzF4274J8HYAF0tOEb+9tlOFWaCNLdXi/aaxPCZyCET
3k3uji9kBeMoYPFiYabv3xRwfUIoI288vCd+vCq0l1U69CTS5FHGueBAY80ker7xShzwXGCAcGMS
VBDAAoVdApSpL98cV25oTUv/joov1uQ+vp6Oqm0EuLbNEJmeCy7ihZyoslIA/DPoo7UZL7v3D17H
TRSLR3IrVH5ABvaCLOkjDHHyGPLRD5a2Wv4lfC3jbvinZssaj3cLe8aVGA1KWHV7taMy54SVGW29
2cw0OrJnGq0QiKazSI+IckkSermL8DtwaetszgfurMx2WWWV4DxwRzm95rZx98b0zNuNYIvKdAoH
iU5RhkBrMI9VJzeKknJOLU6YCN6m31fbhHPgytykkoyr76+aKU33uaUFUksiy8OwDQ1z80vPckWb
v7lxD7SGc9oVXtLw8bjZAIuel7PQSCPPF9tYs5mnW38E89sqBp9hgS7avdMMIiRj+VDs1CeA9JuS
rouM0LMpOxuiXppI/RB8KPVzPfwTu+Lvn6z4p3cHolbzIcVoQAYlxsuMTVvlOE4I1hxrAi4ZwJZI
/cneRW5oFe2jXpM69WuJu0s50fB6XqwqVUq2snZ/ElWKVS4LftjhD0c5mdgX0b5r60aaHNBZuB/N
4U2BQUqF0BZ7UU+SqxqcrR5uwjvQRynTamlfaUQ8xbb96xuEzig/l7fSPM06/8yZWTEyjCr36sCM
mGMAyweEjJsVunzfr5kWxoZe7QnoaBhoPhMJraThdXfKG2MadVrWcSY9Y9Nze/dNPb0zAuXXsANd
WBN0khQOhNQHCag7HUXh+24qk5YeMpyQCVaDksPgIr82RK8zUBJ9ophdEOoL/O7+dCZ6nwelGVLJ
2n68T35jXizYTz+8hSSiIEICUIGazeSa8f77kBknMqCHp/1AlhB0K4ZUd4WiMEqGF+uj72nKgGiH
S421wPKBzprqE4LcXXHq8Il28EdBSMprZLK//a0f75Ui1wBBq9TvS5TU7JirBQ/ni8qfWRvCp0vx
JrfspLt4bFFHJX59CeVhECJEY+H27k+ac1EF/wh2qKb6i85jzpCA5wxWzBtFg731oFFiNfI7I+x9
ccC0M6zkkdP5rwRmPTxx1QtQtlxAuFcOhvEsy6316QqSMzR7/YYd/qU7BIB82duIgYcWceeTLZ8K
gsp2xQY2ab1udqwtvBK3EVKwpSRq32IjJkfnsMq+y38Dvkd/L+ymVHP9qHOPNHLcnqTxDL34yEf7
mentpgFxl9tyMoK2lJdVAteUL4xwTGnYWrnza6Ub5Q2p72gIHBTicdDLyDZ9chfRc8IAQjmP5a5X
2pCRcZKj7HhB1wrrJzfYkopJftZJJIrfzF8QaCSNWO+Kk0iG9gUl8RGbK0MyeCBwrYovl9cFtdne
wIKHh5AcabY8RHlCH1AlOL2WUa1Ov3qWyY07rJhmw7Di1ZCxqlGjIhULTRfhPrMMTNWQ8Ue0uC3t
cujLaa4FTXlD61hHk1fk81o2aZVMyNNRQqvFs7veciXD1llpNkLZM1Y25Q3cs91F9c3ljzeoonh5
Bgna/odhxqaSBIpWyuQs6Q6lKWhiqAAyynea8mZLJ3cAt6lu5QIHRyaN7lSZDH9P7VuC8mT+srk8
jTziF3tT4J5hdpaw7Y7kRnuDg6Wzmrc7ZCiYBVAdtiJmSTfGVqoupbbIe3hoKEPa2dR8bluN5Tsd
g1M5yvQOSur08kKOT9dk3sW7KY5ZnadKVN2kfhXC8Za8kE+m3Zdx2Cb8lKxYSGd90VUXzDkA8uoQ
JhbsMOqEhazxsKKpTjxkDfRex9lWZ3YWgd1hgFRMNW9SA0UlSb9Cdiohn/tjQgkv7KnFV6/9WLJw
Gh/L8XTTOe5SqdPCTvcWZQJ7Fbtn/XmNgKWTfi8qrKt+3E6eqhUFJaidYnRqObIwWTiJcPhQ49Vk
m2z+vihPN+f8DCmq+vRBxcPKnyupD0bVzVUeSv9aoaUCIG2cXduAehNeQYO2qqyUNxSzkvKSfLIR
GlaZ0+WEvBvZ5IBBi33XDUsSL/q6/ZPch9jOgbndteNt45c7fqhq0eQapG/DUY3ZIupXczaVlG1b
lrGtjALMOU8xSMfdAIYvpfVmWSrbsqCHVEDVXdzhiZUqkc/kpfqJj0neLaWPTemqPwnZXnuidcnp
qQyAdUF7HBg0UMH+uDB64bAGdJlA4DXQ/RFje6wnlPR80zVR/eilbPcYl8JMzyYBMqICY+ZgXSAW
X6wlxKlL8KBvFkT7ryZfKmy4aMIeyeVVk0uPuqBgQkvB9YNNFHrAe9uNyv7jCeRmQa0ZBhRrbQ3N
hIXO4Xc/8+C7sD41EwOMU8pLx9WWrFyKsr6/WV9E8SqpZS4fkulCR2PQkMUDsayqW9deljSOqNUX
8IjcdQqmj1aXGV7ge/JgduX5sdLbuhWG55DvuQiQguizLiG8eTzdWzP87HacHOkH9M75Rb3E/btT
pZw+FNMdVUrqCSH3fQOus974zXDYbt6hLNbIGGACioSr/6v/jsmBFhwdyW+zsYbcQL4iPF1xt+Bl
oVOar49YFPhp8aRHXEp7xgThoUCOsVdTn9Ey9XXD0ERSyzWBYqxdTruoyeB+lF5DCxjb8QhZmgZj
1byjVf2m6zHb3C+9iHI6on9tRSNJFBDEjujrKR2BnKo3W6bv9AW8z4XCVpNpQKWw78H8oaLZXFD0
gUjfY7jf/0FfxzUZkdxfMwudEXGyIxC7Kof3lcqBRfzhzEzT4ETkQXL6ISYzh7pq7Po8lVRReyav
TYRWhKF/FppiYZNDteHUyTRYgZk8rELv+bTfq/WtgWHTZZsUWOxN4fc8C6ke3B58k79elaPwM4bz
cQsloQl+Qml3DfIQ+T3GnCew6eBMctTV2iINu177CjZqFuXBARMx+vEYXuPu9wgGZa7ZoBhbhilc
3DQabbHwUwjMPDt8Wk5IzKOp2LXv5GC1Y8reXSmX8Ag2fJTogkFJsVOiudRA7V/k7XZ1wWJR+XuR
fRpZG/N7wdBc1o8xiFAdBCyPLF/bXxj6REH9+lOAv+GL1ZiT58annWMucF7lMYxEGQhTLONEigYD
WbFX0UZq/CP65eU5k9zhXwrYG8Ak0vUwYq6t0ilvWNOidIl29An6q1WELEVFx54dyoIol0/xwHLq
/oR33x2SIxM4PWjhWdt4N2IthFCz32j4ALYXXnkItmmwq9flcFuOBOdzlh5b0Fx6I54j8oSYxNh9
LFQZgQGO+I/H4dJr5sBiUVlbO65f9EJMWeuG/rRge/pnQSm1zd3An45viQgHYwnwSjMXh8/pfrqF
VfZi7ma38QwTIrVIviMTnBjLaPwhsPr2b3Q21fmSfjh7bAWAt1SEZ5fqHlvE6u2qIEeW48EQBVLQ
9Sb/6qBskQdZUkz8c74dBleTfNGPa+ZNagl/cZgaO+P45uBOL7fPLKuaD8ypN9h4c6k9xcmcOl+t
ERaa7wKCDf0ChZtNLZsgw8ImuFTpGagenFjTZQ5p0oclEPQyjWQDPyrzzYGjer5u0Hthj5BH0Efw
UJpM+esCFPeEe19oc/lgfZ0RDQY3RRiHQAadG7sw/10eA0Cms1+P5zNU13/qevppt2p/7Bs94jU9
mLXEkv53Is9DxrhcnVnER1tJlZqkh+RPZxKJwf3FEBecv8mOVndb/WVfJD8xk2na7QYfGLwChhG/
X/a5ndk8lMjsLXL/iCW+2u7tTFv1yk1DG/2FA0vibtaav54uC37K/LdTAOGPMOs1jYi8atSh7K9R
Dg0Rzp9htoO1VoxAHXwYqayEUPX0BtZ3ZE5e0dpOAiOK+2D1JHT77v27ddbg4jkTJsjNZP654OgV
iibb5tE3zDTBAgH2sZBTDTOY2ybLRm7Qfo9p8bnUdvHN1AZO0kfhcYVbVFGm1xh5z7jAh8vOoFMj
SI/aSdv+s99mG+9QT84uJb98OtPZpIwcjxyrvCsWjVwHiG9+x49XxfHo8BZloHLY3HTYOLNygfTL
0LgbQVFB3VZVwVqnW9MqGjRKtIJAHGha9QQ9SynHDDu+SuFodec3zU6F3u/c+cj+4KVUZHVgKxWy
DuQSpIfG0+Y0zJl0mzidZW+aq9kH29gQYz1j2GIEMxMGCLVSuMfWOwDhCnyMRosq/L3DdHfkrsA0
UOek4yZNARv8RnvmkYsmb38GAxxpEcIG3qdXgUAFnrjqPgQe/b+79r0fdE3bzFC4lXwkwliw5VXd
OPxp4ud4y97VHDIuTNIJmeb2DeREl3VkQhstkERJbVU7C8M+/QLvfBkQQkWp/UJI24OdYRsTx5Bk
noj7yDdXbT885+pdMeqlplB1s+tn0qGl6RDMpb5BEqMe/T436tG3gEcwoO3jPqn2/Y6urA5CgPY2
5mhOJh15E0rS69jE1Gb0mWrqRp/EuoYnz0BLuqqv0kfuzf3JuTW9toxg6Rr60JhRBIKprdo2ZrkR
B4u3Y1Hdcb9tetdElT0c8gJMyhckjowj1TRoO6mLCQgCdbeqSXRBa0dVzn6JFR6a9ie1xSUvPfDH
7AZx4VmNgk5tz3bnNAJSctySVHyESfHQwGBUOJEe8IAquGPz7gPVc+s/eUA47jxJDyyt77is/5na
NzxAz6PD/ZyNM7CAJi8B/qg9Kf5E21KIaJ/3GH6e3cR1ICSZoGWpQw5xuUZ5STWOp5+EfLVt7ItG
8FrI1KASRB+cBQXBt+U8GHBXltesMsul1GILuidnCWYqFKwVoEenFFTRrkhEFDjVmX5jp0ozEKuM
sXf1G2d1+pp2kKImX2aw/cDSCYVw4mXseYHnebgf0F3MLXIdV7XQPMLSTh+6vh8WJZPOVHDyin3W
rQK0rqrcg/14p8EEKeIcbCvw8U5Y8dOdTiFKZ3LXT/Q7VhtzbFyny9X9GOfwdvEGtAGyHUBv5AHb
ZGkX0KNOzoaZVT88SUIXHYhhDqfAv2V1RQMSpvwybyqxDB7Z4TdhU9HgWvVEEtb0r9GcLCIKmMfR
skqc9/R8AI4Cw719TpLsRqkt0c6TAKvMpEuWUukbw297cTiXoApEfhkfpp3ex6zAVaehuO4BaR8I
OY6scde4pPVVt8XUhhWmMa1vHA4eJhe8kdJZ5f+cY3SjI6BDTP/FRicnuelhgtJY0OjZAGcdiIhk
v9qM1EG+JMup9mCLpwk/wu7Zfab0SHHKgfm/yszBtNSlT4EA6QhgFVk9QKsjTjEAqMGSH3/ccNjn
7t5/9zqHAFtELaJKQL7eOWA8dzRV74AV8PkEpPusLPNoRvjyMqhl2Sb00ofC+iJTkmLpQpySlsnr
52ltdu1GDp7OuSn6qzHt8rXYx05GceldeEzbqE296D+iwSIwDlo7b4cWMWiTzB1ieWWM4ZPtItBo
pnRAHlYs5uHNfUEoftsXeSIZ40w8QA5u27tXfyIaPO+8fsPqbNG6zfHy+JXjnlBL+QUcVjRos6LZ
iCo3kk40a+HcSrhI0p/dzxIS2O4w+MTUWzV5EEzRbqk+n3ebkxWQhkH/VAyvVxCwGSi7N1pyqMOo
AD+8V+ZsWZDPwhO9UKJYY5HMgmQjU0e6TyFu+zdvyBkRZ/dAB7GMZGtEHlIs0pmWWHAb7op5PepL
nMbMT0oO75jCIpzHgaZMRf6WGmOI2coNnbHb7i+mRKJ3vFywFimOeOdFpOLuBQqicVkXtfiiFQxb
5+McUSN32uDQLVDRY82oI06hqx8oxdmpxK1Ymx6U+FeaB7uHpr5cFXspnzIa5q20bLet0skK6xpm
ok4qeBDCr69Teie1AjOYTSUWQhtBnZ438+pASZulDpdCcgkao5ZGds/ImAEcyQPkY8bONXz2XoIl
x2rAkek7sVoUBuEr4/3CqlxTIs/Z3zcjQjZl27uUE6lscuShil7XP3CSiOVIEMst2dP2Qs2Gd00z
CNGLxx6WCsFxVuE8lx4ZCTiqZzJAYswHEudRmp85WSzZ6lgXpqo9jdaCHc1NC8NDFKcxBXOmMnLe
pltcJeSon2598gjSFeeMLe82oKXgeLRc6CbPF17uANljAk/wYwJVWAZGUTy0Bcssdx1JiLntlrAc
JjpBKD8T88TQb9OGd16567Xs4k2mMjLsoS59dBW0rk0eNq2sfTsQSBh9kNaA2DTxzqTZwhj44Q44
0q3tFsOgroJHlIQ8ajGGqhktJCtJUjNbNGoOyXlTYdK3ibKTiwE3pNd/9J3Fq0ZQ8X/Qrm1jnEzA
fn17dRI92k5mUDZCkUFAhucz+XckWbZjIwdVU5N0zbmGthIWRTLZMo3vUroofAnsCRo2nELQ632+
hmrjRyF15ilgc0RCG+sFLhFo0aoVMUMUH6i64qDDLJFnRZCojcdlcIIAyxJ4KorQqTBm+W34woDM
pEQmX95Ioi8fHlaO1h9l34qmP9ODo2WCibhuNVdbT/uRHirl4f9pXr1jzQB8jYGMzCgKPKQBm0h6
EIvVfoDe5reyUIpZFjKkUKqvxRlhXHM8CBEwpS5zALda2R86hswwnRsTqiNPYpJw9M7EyMX2Xo57
qdjOTvF9xTSLRxYYUzNYTOMaTsaA11MsQqfF5BRjt2G1IWCUg/tFhDpcbqjX7NzDt6IcYrgcajb+
+Eay7n2XdbhA4XgsHGapV/VEh+vim83gYXBlih5Zqzr7sdbRV+K5xLoUrhBUBOluavyfElSvJRat
6pLeZHUWDZoGihPG44foqLfnI17KNGdhEByQ6Lp7ARJQw+Y7yLIIVNskMKGlpPmxaW/OaHhYQ/YR
CZiclnpnRgjRDQ7brYyg56DrddiGtHr8uPqqYEL9NMrySFw7cdReijMbgPuENyTkIuNDBdaW+CY4
aAJ/XYQthvtthJDZXmTZTbCVIURDGf0FVMyzVW5jV/FXAs79emuA7zbR3rM1Os/5D48m82QG6q0L
RbhPtt89+osS1Jnf0hM/zWOUfRmBIeVFHgbNEAy8BYY+xjfcyw5DvhSrIRIA3fr+H+UGBro+Iu8E
BNR0q5iQRsSNQgPF+27xwjZDxB/RcXnFtpphNYKkA/MF/Ue6XdDovCKOikDWXMtjwcF1s2tP7uGw
vvDgTdIfPuilyRZixWypT03AErEWfQ2+ceD2DenahhoH8Z9QzbJoexDOOcB8C1rKoqhTq1Olr+Eb
t71IslmNa+h3YuHxNUlxOgzHqrcZnFoKUImXLOWij9E3Ux7/ejB5F/iaFOdqqC+N2+tqMSm1RlJ3
d68TpkjrmnkOa+CwrU7SMF65lNxvqQtYN+DJayZvj2S/I5Gk+ju1Bco6cm1QuoObIsWxLq7m98/t
3m4y4L9LLU1low4HKCex1brCGZcIcGCKG3xJDHQoBuZ1RY1mF2kXHKYXChDZjIC6eXFWzF5XKJDb
n9o1qVQ902hjmG2dpA3ZBqrTSYTidvYLh5vogIaNnHubiB6i/MUOcg6q4gEDXQGg1w36hBmakZOq
7aAZpUEuydf6NEEP/pCRw8aIzlpoPbUIwbBV+83xqIqD8qivqQfdfJY67qXRPkxFeF3+a5Gdp8ZQ
qh/Jv34t+RQStCmepu/NsHeuttFYNyPdWr3Mn2at427xqykUa3Lwn49PgbX29Kc8587JVdXoJx7u
ihfw0gQu6M0B77RNtNS4B/sssawxhvXHguyAaBRHS89GxVlqDKFJNcY/auEmHZx5rsCMyCxBz7CD
Px+Zo1NNuKeTs9m6N+SjMtdiz2XuBO6t1nhZAMBtn8q3352abVHGEQ+M+/Y9veixcWNs9KYBTOZ0
IMBUJwHTcCfg+sB/t26BoMvm1PwLpPDSxi4kkiUB1V9fSjgx5RMue65aLN4LgXNsIextdW6MSvWI
quk/VOEonwu+f44mWqsYBFXZhUNknfBejewqrItTNMc25FgasIBBpVHhAJVReYwlhJOKRaGiJvMQ
lVd8lCYW4NuJIqBprFcekPq5lclmJYONEPIv+ftUu6P9IBl39xO4DjMiuFY0teE6E0RG5kMIqJEN
AnIMTIrJ1afvni8LRz/QT7kgGWtA9Llor17fdcfN1gpB6FSvU5Rwtav03dpUQJmNlKYNgSGn0heS
wYkYja47MEc8tbst3OaMlEJRRO5XnKM98S1rebukkmtMPiQETUKAR9AUi67ueBgHXa8xcLcIwNk+
B+jCpMuIQpLUtwkQmXMHUPezssfbafamVTSJ0bDl3TwCfuYKAJyFNlzgAFtwpqoNoLzWZKsidVEb
JDq/D0K9b/qn3qjPB5Yx5DH0cKpb5EI8zcaNpipAYVUm09Cm2sAgiax31oFkchIvc/239m6VtXuP
aswVQOXlSRvCWaKsoffdouReRYrMDmiYdxUrSfTWuCfdA4G36lWtSpL1DnenGifYqKDs22ANq2ZE
/KpgcSs+WWZBEH3t/lC46W0zQfQ1/4VxFCzfOb6sMIp8ItpwNl9ILwgD8KY4hOoykACPPpF+h2Hb
E8PXBMyIXPqFAzd5wCWWHDFeiXK1x/VKUVlYfXiq9x1wXlCuVZ05E9KEHwOf94pM5zmtRPui2YeF
RI8ua0mGERJYj0PCxZpxoFv/4YqO38AqFSxv2iyqwf4Qt52ZBaQPElhibTiookWgZZUKSgTeJyco
oLScNRJebScxYQLUg6FdKcxw6lqOAASdypNjx1cxfw6HPTE3G3ag7O/IRCqslOyg/qAiglhRjBPH
4oy/ZKZE0eFYVL3mzCS9EjuFtjT2wU87NfEdc4E7mgs25RyvDHSGJSrloaqkBkQeMvSPkpgRT6Af
J+mmhu2qlSjuTvVcZos5mFPTUbo4IdfRgbUNmyZFk1hv9oM++CdFthlXD65CTINealMkSXgQnHmp
QgRsWemlW8KfT71n/0JSc4CWt7hpwmVC3JiSgigPM3e43IS9ZyamonXwiHBMtJBDmxR2p2ciXaWm
Ojvn9vwFNdOebQ9i0MqF4COel5wMrZsywa2tLsqWpoBbGjWS8VdNCsOC764DpgzfuvwjoxWnYtYF
yIqoCRHuS0+yV1OWB11KEYt1a1gKgIIYRjQo1EIL2X2baqiwhDmBOC7WBycuhAdowVawk7aHcooX
EZVMsO8fJLOquUUoLkrRND8zSW3SKuQaR+U18+yEwHWibUi0Lpv8OiwIc6llp3+jJJEXecFURrvQ
cyZiJ49hljDGZa8RJesDascgXLx6HNVH+BpMaRyKyvwfwi0MmtEXSI1z31eN5sTHJfJYroRCjK24
qRRm5Vhf4Ky+h6U7AF6pG13cajebA8SE8/lP1nBTP8OBMWYEzO4F014L6gO6y24kunBxAaAs42Rg
0kez0MyenPvC3ARO1tLxkaVKRQ5E62NO4Or5DYLnhKuIOlDIWPj6tPeah6F2pBfr0yfVGchC+jnL
xYFbWGpsUHnT2iSnZeKbyRcParhqgx2ojMjWmNeqJi7UGvdepXyTPY3tXImE+FZi9KIVDkA2i1ps
aagE8xvgsSBy0j21L2DPdU+YyOxu4leeHWk/18/N28DamdcvOgogLk6sLNadlT4hv6w+1eVaDeU6
UuAMu3rInQTb6uYcVU5NzJza1KO7QLZu0fS5OX0oLJBBT2pZa/UH8qPOfX34V7YNKpAlfD5XR3XM
hQLPUawTQ337iTXCLpHEeSJag/x5jOYN8utc/hpNsSYBu7SILLMzrBh0cYm7cFM0W80zrdo04GmP
AT+rV4n9rUevN0GATIv4YceAULe5lwCAaAocfkUriWuy4O/cnJeP+Y/QjAMDr2ZbgGnZY3BrS2mG
uVPrYDXIsMwK3Jw6UVeWmL/c7nba18NioOoJFjOFkjn4pI/jVfnmnkNylLr+uH1aw+zUHRRo3Qor
EKacWlm2j4VgLQn62OL7buDQhVWi2E/SvNAIJpQAvPUixvBns0CUKPUe2J75pbKp+DJE3G213H+3
hwZzsiGasn7t3ecUoN3e7TSDv+glgSGeFSWKPCn5zEcS5DnFaEF/vZCVBCUmKp/5sdQAaliEGQYd
gml/hGAtFkfe2A2FKQ6OwAqPaUQgAP6XmfzjFAGIlWggSrJj2OPfpe+mxnqgEjaP4brjYA9mL85A
h8Y6V+3bMQTGK4ymznkAjDzMOK3Q0yXQ0o2pz+zVbqXNkcCXEDaCMTmE1XXUYCrkN4qWxC3eKr4K
0uBA8tJ8/2mIx8dt+jqUaI7MU14x5DjjOELGi2jfxzSOSRwoxiJWo++5ZSc0n7B+3Q8c3+XN9xuN
ZHl7uHqosUVeODpqNtNlikdrKLev5KCWlnZsWihMq/TGxGZCCA5Mu6GXq6riOpjbhPCXCYx+ACNm
Y3nwozST1Vu0bKe11wmESTUldQ8ZUoQ6fWCdM9Gzy8jGey9qQQx+IAg5Szk36gr1DO2m7s2NDyKI
PjRx4Rz/QeTkCUV/gNIqDtUxG2K3bkZ0xLWV5agu2YlEv9zld03b6DpxhVrJJvDS2Vt6QZSijiOf
E3unpkxq39+/waFM8fpkhb7lzafCVOCsqUy0ymy+ELHhNCNpmpvd1DGpo53n6Z/1ASjCBnAEXWxY
hWXj2oAYuMOizSMqB/lw00CjGJ276NVjxGw8gnBNc6BCAreniECDJG6JTpHA+iC9PJb1MBPx1U36
8qgcdAsK7fO4Iee/V2htVYFZANJg9Wea5sMm0rtaO4N0crsR2UVhW1nNNm101jz/SL2rtms73NCo
0bj2ibuKnxA7SW4Y7bs9HsrGBRuT6HUSUDT3i6X/vbzGjQFWGqJfqnqHcMWE3GzFN73OvTxnrapA
5YMZWpcIOyCbJmf4rqGegYqtFL+LT92EL/akHasKZ28Uw8DvswZDG1lr46LLClWOvmnCFew6sQUM
7jaFVpKwrjQlEJ5QTeTxk3GzQZ4MXlxnCA+iLvzTvBwtLCf4pXxA4+oygi3mHtyOvJpBkA4M71ny
h6D8l1n+4z7k+yggkwD2fyGQ0VsSQOJHzogZvYV3RzKUsgeKHOBcQT5QDoHnLrS7329mNbUIj5om
xyVnmlE8RW25PmC9ukWW9F1doTa1cSlMI5LOtyJ1EddoDhxvUeenNfROZ42qxxBGvQTu2defEtE+
5tCB6fXDVKb+2jRO6doQcqASs9tDqqZtehF952Dvtmu4Ut2l89Xkyb5SiR1AO75NwSQnUdFA33N4
sx1aM8BMMz22ik/lqhmz5FON1cfTyxafKKoJF0VuGG/NWOhUs6oU8ZPvhu6GqCL+WgjO5CplZ8+J
9biLLHqcz2os9TgWT5ynPQ0TOu6mIHL2S5zKFzUMxYJn6ajZu5oWMGUB37+m5xoeuojUT2JGY/Dv
s8w47ILedmqEWnYk/ufKxeLwjDLLPL5ffzCAYhVZGMSSCX68nD8IrOFmQVlLvn9hxS296Zn3Wg9g
Mwm8xVMC+L1tYu3bjFee2IkeN1+xFyzcBY8goNQVdvFB8RuTV9VV3caZrir4TaX96qt02cIfdQ9I
sAzmQTcGh6fl7PHiU14v30wRr3CYrQqbtr7IGaweyUtUXhwJIi3LgM8tgrlwV2RJbxfCMiCI3tGD
Yv6lep9DMRt52FXdb/Um7iy6HMNR2QjjcUzzDFqXlu6zmbBAMu4NXXHX9N6twZoeFilyJaNSG12E
RjS/IwOV6zNHFP28eGGxcBLUSF1V4ett3s39I9k0b6qu4VpxPvSJIV46oXni/skiHqzwhChb7EPW
UF+r6vobcY+pLXtRs4BwshQaz0LzxPl+WheeFocjVvMKHTUawRq0i3BTWh4yTluUAzXG1N1HMyr+
0jvrQTEMLPLXYfgnZWrUO4cNIZZOXsah3iy0EOafXa8VRJLwnwf+gRTiBYFG08FDoLPERZ/FKulD
EKmsjOLfn7T4/DeiT8mjMT35w+KcEvkyn0baGpd+o1TQaeYNFkykCsPLw5DMRYGzXLnVJvS2aFZv
CP4Z/XRKzgALvvs+G6e4NJD/AQNvkkBhCikpT9Lp6NhO2GZapkQBhHJ1GNKcoLEJ2Eox4imdXdaI
28ShJKQTabReHfgQCXa5jU73Ldb5z2SN2Roz1fIQI2X9MNPE9YNHzP9ESq7Zwc6WO3lBPTbYTu95
xROUODovq0ZWQkGoxIKQMkmUct1mk7/36jyN3N68ASQYGijUOPY5GxF9YYon0Er8750DhgJjH/+F
Hwd/qSOTTcl1+Qit1aDLNJtxMXY5bCL4dJ0ytw3IyeAYKL+zGOwVcBODYD/+O3qANue/1V0u3sMT
C9XbeMf7tqreLsdii1GYv67o1LcsOMWmw6fXrhsbREE+oo1oNc7XXiaoUYSfiNP70po1eVkKfkmz
GE95Vsr5sJ0paGs+pcdNPrGmpu3y06HsusRRY+oRwxn8y5PF4qvy6CL210FChI2yKDDWa0WQdtpj
Fl2Uvp7eOBdrqChQSwbmkjQ6hr0jexEKIMwDJu8tvezUeKmYYFjsvz9vV4JJlADPNLuv9XgJvS5Q
sVG4urnrFONh4u8+t5Debd3LOTA9actzJHgC/YLa6Lv0UzW+BGgB5TwR7eYK2N0BA6dOf33IjD+w
jk3DFaET1FSK/feXd4iKVwwKQw07aolPXMzd+tNevqUxo1QxyA8k0/ANyLp9V72NvsKE+CMR1yod
uw9s/Wa+fEu2noa85RLN8InaAhjFwkwyd0yZ8RGCrkFsd/xF11LZT84GEyl/XKPJ8ruOx2v92Ywk
27z0IA6N1XH0WPGw44VuSCvCYI0bR4jTJ8I3HYlo5aq63f3tMS6frDcG3FQwH9W/A1g0XPYWsQD3
yoPcsU3+BEXPB+7y+7gsWC3zvQBxOZAIO5Rnesdide0HOdmOHnenmlJ4mM6SkKcfmVhXUhjiV18T
lsxreUBXa5nrjYs5xwnxf6PN891PtDcyCgvBqwifwxKnX0zzm6kUu8Y05dN3zaZOJXRhJ3WBaPNL
aFzpIwRStihlLpf5S4nlzg02wyfyjahKe9dCuNDMROmvoG8Ui2siYzxAYf2w2fmAxwgN0zGjcFlk
2QJWMyQoa3cDZ7yM0YoV/YrSOa3NSqckl0ZWy5z7l12FCnpcHd7XaSOXHqvJtXgKixkP+e4vWRwH
WVjTfCrrpfrrBYRtvjJcuf29kPsP6potzs+Q+PZqhhldwDzQLKKrKguGIMQdzTU4yEzvsBN0yuli
kOLRyFBw1Tn57FZ5tGKbA+o7uvVczuYo0vFzls67OP6sCD8IX4UWyVM9BbdTr5jkONZWktT2JVrV
EtwPOCCD5LAO8R9wCcxa4Yqq6EEnppfg8XlXSYMRXD15o8TyJS8wP+NDu0lCsMAM2O0i3QWs/OoG
Wg2mpgoIkNSwn+13VcmueEntQetGxeTo/lWdY401CuTfeSsBcs7B8d1XraDpU8YTYzexHeRT4WNB
b7waBUrqDlZHjYiS/kAVUA01n90L4gVSwf4WyX8geAZTH54NeDRUBKTwm5VTwVObElecSPdrplFR
Pgi83xqLDWRuqdamP3XL8VZDzfuvMRDbQLjUcFhPPbG625kUT0U8C42/VR67NAgsDOG5H61Elsf+
tCR/lPsXcYuxYBgQOqsPcs2dNh2kyvhYZSskNDrWBa1WYvznjEw8kCHzRTe76dhmofjkzgs3GzEM
8AsIA4mclNJud6unvHUnMuuFg7eAAEm2XDDPw8nhNjNVwc+sJ0VtCJwAGDPVsqBuawX1f4oEeHM3
jhBVKdkBsKw2NYOStU6+3oQjp+JPvDIJ+ZGsZX6sw80MHTXbJRu4zzmZBEivNq3ZqGu9N5JzKqeJ
O+GW+sjj4qcplyH/g8VaHhirWHYXpuP0M0aww+4E+8cnp9fjlvysqeaAeSxfmivXI1UrlbG84/Gm
RtYpYr83XeeqP2eq93T6BIzh6Nh0LkXohoZc9V/RG0sPx6/bzYttqRnE5scVpv2xA7ICUHyBOEf6
WW5Ma60h2XVuKuI1qP9YNJj7390iFDPOBrfSNAUkBk56ANM/RtWkZlc6hRTJPtoK68eFTz1cxi1+
g8m9v1L3oQMhCRJD/BODYM/EFSIHla/B1npoWMggNIPzSp0bk9JOFciELL+NezWh4ccoLnQ3ocIO
Kww0t94iSFKelaz+vCNwu6ZCOG+esLPWLyGP1INFAWMX+jjxi1dSXUKb2orao67xeCjOVs1wIhcW
OqYJu8zsj9Um4/RgDiJ83K35SOkFNQDX60wOpSO/kCHMvPpo7tqDe1sJwaU2FI98gWIZib28PR72
jk4nEoX9FyFZmhJmlawI9Y3qEl1HCsgNBgzCzcxk++JpT0pyyOzLrjEApJK+XZc4sxZJaKT1zUQF
bgD2jdD3HO2AM9x1d2Ak7uRPptgHhZ9PkLeMAcNrxKXesrSfwKTlPbgqbD6TEwggblOAKPAAp9ny
PGCV2LvZlTq8aPNPUOYkmqr9zKVxHYhxqJX1b+O+hW2CCo6QXwaIq3+9fUMnPQwxHs+p0ZRQ5RCS
JvUBvXs3ice3bo5wDdAytkulHIMzUeiIIcKXIwVNEtuaLulZhb/nMgy72XwThJgMhvGe/oz4HMAB
yf8Q6SwWekG1R8WI+nj/ZZluFMvdkeCj3r9YVV01ZVEIrhwwXRUDVOoUBzgIVs4wcuG+AN6pQ+Xx
GiaWJfzqER4AnofryQgOiET+1omZUM9HnuIkVhfzdVLw3k9YTx7bncrIIxKBgqUFs6p6kexXXff1
dIQnBlrDUqYDH4JyxDnPhSDdwMob6RnXBph2Pfjwwo5Mr2/k/7yoKDPxj613tqAQYmAKNw+g7JID
kZT29dn2qfAnkAWf9Smqzh5ZA7it4UAugdYWCFwkRVKj4lKiSczSGMU0qfaPiVmJxfBfCyDvqH+e
PeGcAYHRRy/ojizKD6+Xr5+DqYEltHgffez3nRtRKfhxxrl5rMd32pAX8yH73mqlVtGcHaPswIfF
bBITIBVH0fRjxcljTAkdrd+5fyk95KGYANkv+sv0AZ+fMHwqxj4s0HH9z95wPE+VFHwNLhRlVb8t
8ziKt2DVKy1F+PA83+8KiGCiFlUog//HVDi6XZ40OX3Y89PK6Rfc61Mjst+irQVXd/rKFsAwLaWq
FPyOjD1JKydZ9Xwr4F3ec3A4mjsFcQZbpD16fupLOEDBXn/YdkFhub92VTa4OI2k3vppvt/MJ7Ed
7r6XwGK5J1+vlp8wp/LEwyYiyuiSo5Mu8OtmtTa7WK/MYFgmXROvWWNwHIlr+1BzilT1n7T4XSSp
qVkRe52flSfM5ylt/Ar4so7mXodXsnFxRHncEid74G8ZrtyS1Ml2vs6mV9gKMZXlus1Q5BcroMAl
zI9pQah2HQIsOwdaMMy9eDInjT65eCd6OES34izfysgNQzuXqeCBY4/KjlwNburz/yiD/gOUfCQa
gWjDKFiR0/ghcgETehCKHVfDx7vsVbKrHx5bzT5XLcuJp/GYs+dMmoW2G3fB/83WDSJgURFK/hcK
7UrCIpSWbMQi8H8VK141Z7C84Zs0OQjkykdpr9sUX0GdZI5zJaNPvDyJZYx8nPBiubhk94VkEUuy
Y2lE6UbhqHgWperJZjjX7VevDJKcn+zhJ9mXi01vgzGm5aOMG5bgAGbS1vYu0SNYCmara5FmRnBQ
10SBL6+LScla44oCjGkzxn0uf0ERq5zEZfqpYFQdB7N0QFFuEh9S/7b8p+RweIyamPYMDnHORmMm
scH7eP8HWLthdMTLRdj0lccTIAbCfrYrX0HtZ/hUoaAABEw/J/AF4a5GVHJAI5HEsUxdl54V7ncG
qkDbgXwJoY/+RjnjMcX+IIgfO7lZYt+NRupZY9+dzrL6Nl68yvZIJwMwSMgbnnK623In+pq9eV58
l0mqXL6vihqLGlt5ARt593+Tv4xc3V3sn4+WiVi5/lqZFVeaBNgMJHTLUQYG7X+pwtjIpN1eV2x2
Xt3wRFq6YqM9caXfiZ7Y0orcxodyrUgYiBYjpDBAau+5UJim0SduXnBO4lvzBF6uCjSXtd7jFFe3
6OqTxfjwaUMh56XFVv4KRfnTq/lRwR7rXXoqf7nHZoQFdLZMsgiZkpG3m45+ztVTAkYtTSeULj0W
AFVF9GpfUjS3mNUfg9FtFjh3TT/cwLW1nPKKS9akorDe5CmcDQBfEKIW9JDD6TMn+XfQoEAA1AJl
yb3czVcGvlg8C3uSldNDuwKvL2T8b+H/56p/ULU4bu/ZMiR+ULHMsaXcXHVyqqyvG6soltcBNKpA
tmMKoPWRzNUlteQNVkRGHCdgp1UcxEkDu00wN9avPjEo7voj1FXn4u6GR/GUKJr2qAELGHCbRPcT
S3Yn8aFw0ug9G/aXSG1phkYhl5xOziGJOh19g8UGxJR91JPrkYKZhZv+yr0Jeupob1bMyhWdVPX/
XE3EhQwp4TPAzeM3hWnrAciCfGV8xAS0ap/tkYJGlz/MQLsB25DujrK8vnrb3hkZBuKuY3Bc8KRQ
BkcO5NsOtxmYnXZRPYZcpidhE3vICrScYgwONXw99a06rTC8r+zpXmW5xDuZwTZbmyM4K058ULgS
lecct3/TNletEAfgAisjk90Ut7OVEuF6xTOgiiwgILMliUAAQsTEBYDGyS/X53s3EzPXRUM51MUB
axLkO6ECZavzq/fVVmOM16QUSN74BwxvpCwxbCQZbg4MxmdEHIXiy2TRRpVvwY4esl5BCZo2GlAq
qcXHJ0JaVAqrKrFAkRPidCZgKCYvj+i2LYX/DZWEdOU16Z89ZxsLD3r/JXvtViPaFAFAnSuFlYVC
90xGaWQknukZ8kBalnv83brjIspVdXXQx43jJnSO2IMNDd2nWbSKrJLC/V+f/pY5NgSoLoiTSQbv
7iSqi0mTIDA/W5aSFkpMzi4YYShMEyg23ewNHjnTD5NuaN/63xdeNzhpJYJ3dbsN5mE47s4XJ1Rb
BzSil1VxTrj85wR+wVC8ZtoCJOuSLFj9ThnnOHitpQbzHQeudnfsVhTpHg+dIODd6izZESy4RX7j
04U7oI0gW8nh0o5mNcjyqGipRYvm99eGTj37vhxqqAJwMZw3nWjjAhLjdpQ6Lm6x3ctOG2ZW9WuL
FvIEh50RViJsbNw8a9mmSAX6akbqwivoFWXTH0Scm61QQci4pFdLz6AdTO2CBSZlF4sAlE0L5DdT
IdgjZtAhJAIyqeAVs/83q5QEGdNg/7CB40aVJzBEROf9gpUISzHQGVoyMZMP+Xp4PAuW7pPlVJ/t
kdpI6C/RHmMn+NcY7Vck1pBd+daDwwSlJIi0JmMu4XO8KAuLXn/tyKEkLlP28/2KM/fMn4pfE2HC
VgGTzJmOAR7YX4r6/9FJQWNUgaJn6sngI9P7vQ9g3QRC/YUyuI00r76xIgtVvqlvPvOl61FNu1V5
Pdh2vE+L5V7Kh5PHZCxf7RvlzxPXQ1Nuxrel23aaDV0dl9K4I30VOgPmkjY3ymMKPdKjrPh8n/05
lwJc2/pgr7M+hjQP2ZOZdbV0DViyQqjvPzipmK56i9GfLJSbUGr6u9DbFBhszKCUO5PMwdUrAI22
09hxyHqEEvB/SXgMkOLXan72BdRSSA2PJF8Ymx8l8YfWGv5PCDCA6kHbpEi9vpo0B03Zze3cjVZw
xRsjsNGbYHTVvU4FMnCUCSyljkOHkv3kpwzRNTtT4hR9e+xB34Cj5LRx9U9JEKiqeEfHVaA5X7Oi
rJhZ7ncLCFiujCWz/ZtFxegtH/FHTpZpe9ahnzHlLb9Acl5nK0IDy5OcP06TMKEiEGfsJuwp5wyC
2Qo46AUeK+j5c6cduyIXY/zjaFml6kXTNh63al6IxjL6KhOLUtK5pnP4uYdt5BmZqSlRAUoLR+9F
47mKFI2CmXPHEpwhwGwqHYfoUIqeRaAsRSq+qf231c9KwXgg8+UyXZtK919AoMBxAa3JSzxUJ5p3
N9jKBpokb6vfinOnayA7zFcRHYlXeOzNtKiXVN6uFs20/53/OSUtadzbgGStkEABRGHw0HFJ/8d9
B9VVtAai6xLsWPwYaTUIUj3rt75VBF4itjidmOI/i53k92osmNvb0PiH8N+Wb8riBurXMUjeD6iI
EF0gBlJoLYo5e7fVXwX7sU4VxpY+tR/olBsJsVpenBbjt0V2YnG3QJxiwFuTvTr/LG5tutQ3BkcQ
qarxPoTaOgwWwZ0Q0mp1OyQSqT/3XYShywlwfYPks+2oTqTpULFmcydl9EppDPCkjp/oazH9u/Xy
adq7QSr0TsMrwSbKMk02+MQ3EyxGH4GjYUU4fkTvTKb7lvXeHn79e0HuemfekA31yQyWie5s1qoQ
HysLlnVWM7d5Bz1vxV1MWKSfDzk+oV7wMcQ5u3TXVKMcF+p8YI1mxbblh0Uaaf0P06b0PnTtyLpO
K9hjefmk+DtQ5xX3dqY2LMGNPnpmtZtk3yzNRpvPqI2sRUt7bHk+a8/0OLn0+rFiSR1DnjgO3OCX
e1KqUl8qqn0zP0xHasQxhPDNM2LIppgsBQ8wkIYkuBqpTr0NLy/bU7vxeYLH5N8ChbdeH+jeeYfR
kMH1qH9QRv8J+k9tOWx5UL3tlyArjj43ttGqcK2mI5RDNMEMa0H+UB/V+y1KGKXNyLAdYqwltAox
MVDu06ED1jNEtxeuoBg+Pwzao9LwQUUqPXEEaKZ8v5b17fbxbhF/xDV2I/4E+BY12XiWjSEb1Eka
DCdoBTiiTZThJLea7FkfuRxI2aoS3CINCvnb6J7hqo422SiM4GXZJirdYX0W5DqYPC4G+QLULj0O
Ju9xbQ1frT7dcy4vTKs8PIg43P7CQEBDpM+jySI7PFZPcC7ezsluB4utJQ6T/XlvHH+pTAKmR/3m
8lZX5OwscStm2tDJ+9v2Ftsu7jsCoJv8XhtUMqQXOTwVxEgS6NM2Wm7w+dVdi7J1f1RUM12d46+l
Xtr9JbtIHEvtlWfxZ64OOsi6CPvAGuXBC7sxuJJLgDEIuJfAjPYnXLwsUP5gJF1VgRA2yI4WYUKf
hS42cFzCgqBEjPBGy27HExl+U3LeVDBzYyrIEmVtY/WlIRKTbNiou4eZvQbf4qrBg6436G6VmPmk
Xj7R0aFPQiTibzCQRq5j9o8VIwbEIcb7PlfeI4F2SFANF4WweMj9hS9AE2HcAV6EQ70Rryn6n0hi
asu/jjdrAWAgNxgaMxaKkcshBfufpcl2PtBMMXsNdmVgno3EXG8G/FIncsRbUdFgt4vwxP3aWJEY
lVV/TszrePXCuj6tCcpRk1+/LuRuIlUHcUvednTSnZorpkl4e3UZDC+qFgki+l80rdQ/4RYoSGkz
fxI9WU8GmIIre9psHqrZmIPILMUTrvA00sxq26fj+8mRR8ZLKKJ0snz9Tw/XttQKFFBy2outGAMz
sEkgh88AcerJBxRFwcsRsz1npTpPufMJ3gzXChBi8fPVQN7gPvI+8gwXR1vE72Joo3OoG7vglphY
7F/GQBWFaEtCnZCaaryiFUNra318BQQ9HUq5s9dP+vmhuocfbNaPWTzIJ9qVOLEWaP8ZsgxilY4L
XDGJ5j0wmWz0nCU37kE6MRL8AfKqxGJLAOj2gFdUAfWkyoTTGTdB6zRmvP5HE5mvE9OUmxyKt8UZ
fXr8iSo5FvN55xqKrQ2Eo6l9bHSXJgONHK8uJTpvI58c6Myi/R/2M3B4mYTElykMq4vQ7NL3V4K6
RcJzf0sfcFZOLRC29xev3jN5aivRKDaFyXufvYp6CyZPPX/+XTSDikj3VyNG5MMDs9oLTlwOf3v/
A1++hM+pd3p+piYXwUhddTKoqJadUCxvRZoxKz1cxK1G0eDX/owS0bUQgqo5RSrGifiA5TxDqcLY
PFht/wykcNud0K0T66/F4ujjFL5AKSmvfWovn3J/+uC2PKmJYkwpM8sTSEO1QFflJT3YoP4ZX7Uf
JMFhAqwh8pafS3atJV0m9/y0sSBWnZ7uEVU59KfPFPSlNgwFF+heXT5M/nzQ8HFg9s05s5kSmsOJ
/ncNppqeedOjTbb9Ko62uG/2Qg3TX3JaadDnvxI0q4djCVH7OZjqyjijYDVSse2DSbGS0Zwv0wko
BO7R2Nj0WsD7Bt+2ALwBr0tDY7cp9sYsQ+QFo3EhEzwk4hSoGqzrNUaPCjEvjbd6GCst2adGify0
osqwVtylKR6YZxQku/mVnnZOAWACLcKPmA7ejAZI7WIdSQqpvf0liRcUejqVxLNdYMVtxR/ej4QG
YQt2HZCZsny4AB5Bpr+wSn1aRkaRBd4AXW8WaIVShCfV9qysxJjobo3makNLESE+genst+lqEG3Q
UWQjd3Cn9zFaR6Btac22wX+FXyEEbu1QpCZkAJ+WtA3mHsnaUNJ5RK/exyoc7P22WyUjRHR38TkV
9qyU6+Rs69x1V0pWquIpdLYL/NL7s2kuqu3Qa/LddrDrKb/85I/L9vH2Q6MuW6oApSGwttvVeD+m
j5tsuZ2Z85vqXlkjBhEhD7GrlUYovS+GXdUts8/a3H9o5w3jvnG8yDCINn4/NIrJkG6sGwjhXwKN
WtZxUF1FmtbgcYwkIwyVy2fmozixeVcGuiA71GBTnY4FGJyL4PKp3p8GfE85KT7YkQ72Zy7Dy1Kr
wXm54AQWWFDf+aK9gX52/dEdIv/21X+6i/4xELQswq4hXxfeW7UZDM1eOYg+LMEn7BAJKZSoMhiz
rbKT2mfn3wFshwAJ/GK18aZ3rMBeg8YNWvs4g4R9umngkE3n/R3jq8pGjXAQZbrrdbqtW7iRwMmv
VwiD2PNfJEGULDCO0YfUvroCt2dtvJS4ZTKFTEvcVidzJjnj93cjExDJK9Tn9K/s7nEvQH1YWM7y
ZwlQnch5E2oFjvJIb1biORtoXgoy2+/ARPA3J2xh66J+p4uKEvzL4cK/Dvfi1nb0U38IW4JmcETk
RfLljjT3JeNNO7g9zfkEiX/pPyGeGUQlw5DFmgfu60GEVVN7DeLLNdJc5JYHBM6y/2wlkfNdhoQv
FcYUZAaMYveS0usx219oPNsEAQQ1j3u9Z1bBqvb/JPxdRD6QHPtffsxv1KEBfIMOYDnaqRcqH2dB
4HdsqDHD4hNHwdmmEVuWUaZgK6zUHPGWTk26l2ObTP03pAckjjDd0qe64fTQM/wFnlJyPbo9Q7gi
f/Ive1YhbPHmATlSMn+cXXnSLZSvtdPjYXww5GeYCzcbbEB/xf/66DgeqR5DAX9RzI8irLRqXwqy
Jc7nsH2aQ98kLHmqnbZllXjN2K52doCRkNkKPH+weZQkT9EY74l/AE8YCxxedn8vg+E55Ry/KKOD
P7FdfvWHyqfFHLxuI5mbdx8WUnBLR/ohrawY2JWq4NmOC1wDeF2ZANgz6QAapeTvwCr3muZPgfCb
JGqWCn+GcaT8z3H4XS2C/aKxuU4g1+IGPAz5te2Tb7CGs4hHKayXMblWeXsMR/Wjem2/UKRUp+Gw
emi3Oid+hUMjzetUwKZ7HUDwCCgprWgGgOdRvf3HXcMXdkl+fExIvGLWNlGouIHtDl+V4KAPL9Ns
KDc4sbAO7ZrRiys5GXyY4GNlw2UpHEvo+odqYs8IFgjOzydoQgH4DcdHMP8QQWABzDlV5MHrCYz6
IXFtXEPVNrlDBpi5q/mXTQaQ5poV8+xgGT3JN1dt+SLkB5V/s1P4X94MHndMzykLiRibIV1epYkw
4FVpmktqgyLbaIT5gwr0/JLM7GAdYnNudWqGmkgpq/id+QlES5R/8nq8I46gTKGvCRJnLX8ei7To
GQR8u1wBEtczYkiBaFigD4JFKF7GZMgbzOfW39QKs9bL3n1t1x6iCQvNkC4Qs1wcQJ6Pky41Pu9C
vqFMsfDq49jvfg8yVfo14fCPfkWfIqhMK3U9MvLsUi4+YzKO9JWvXZrUYwvr4zq+JHlzeFAAuh1w
NU4fN2HMRrWnMYsDuRtl2Hsqy/EgBlLtUXJHVgr104RbmHRVUzwJ9PG6fGqkry4Xj9DIw4SajmAD
4PnqWGIiEbz3jE+llFzZlQPiFjT2WSn671+NWKlt84jAaGbmAu9CjvDac+4VXNl2fawlMkQRxdeq
oT3qConnL3DbDWR9Y0FpZ2HEoGGJkjQg0Sl17MB1+OapW/XUpXRIrTt5odJfhIyKyA93sI58LM7Y
tEaFRYxP4XTSHqhvgSCnrwEz5htktltQV9Eq0tFJfFLdUcvWzodIVnyulZ3Z3FH7GuvNOCHFGLdJ
QHDB+TomA5pWWONBKN+C1LCpLboa1FXgvgFpC+xElJIZWJ19zze4LuMVZAOyaYV3mo9tkuCou46e
ie+LPXOy4fCTBXVrpKnAn8/02GgDotvxby1I1kjjxSfWlb+Uq2DWKClCFURoJHVwjJpeNW1CunoO
Qc2gpzJRUZojzLPDJhBR5Mhyxn9iZqltssNp9Q6fi6Hv8EgrlGlpzcoiRuBSvEBPUE2HZu1Xe5ul
42eesRqfGZD+ZObDakKTOOkgZWUZ3s3i1QxFmClSe4cBnCeg8oHPIzMOBZxcnwW5WRsP1mqkrVJk
qeHVcQ3ucO5H3XiPX54oAcv7eNydo0NR5nsaNqVmYJb8ilsXJW6Id9BTp0LNNwld6muko0jQvcPV
6KTd67b8xCMUMcbnrN14fi0XB9N/T4pZmuy0tQZXLR7nRYo6wOm7gMGQQtA7GS63r5XGOnJIFbD6
NkqK7Q/wLjO5xI3z0L6TQS0nVAFfGfknPPo11c5Wdd8k1gQkxOX3S1j3tPzD1VieL9tB2gZzt5gi
YiDpNM0WnFprc6Rad8EaQE8eSFF4HnoRyg//Lj6GsOWsFvX27kenVtzYUAHYFkp8N9VpRvWgxjq9
6iuXrtQzl0FHHQG+64Hz81f3rQxXK9HB36uRMcuZO8QuW88bHbHqi8UAtk0BLMbw6XO/v7rkaA1Z
xmnR997pswTS0iXr2YMc5HkhV9RA2qKevPfFlYckkL/Sx4ahgzgL2Y2oj0kodZCbj5zsUzEQ7S4h
OWHsaa5PcDgBDpZOs5+czVwMbMDyLOs8FQy9VCyLhAI84ZR+pZEBLlIucwY0dz7Cpl7lEbLl9EiS
h98eDnF7cmxATaw/BxUXLYY+vKtgLkHF0cSUr2JKJg4AuIRp8sPyiCiigYxA3RXGRsT6lISBdIKa
HyTI+TpD0hBgvAZIr5NEmo0FWKYZpP0DjB8Xnj3eaOJK5FTh7k9RgjCo2YXC83o9fXWRVT6qZYA3
nnO6AI0/nW8OPxXXsnu5X4WvBQsBVdHRjSoIleC1/apK/Bcn3VNhQfP9QMsNawusJmLD6KMbja2b
ef19DeeRJVda0t8FM5u0R91sX1K+sT3Uz43BQbTm+3kwikLN0xM3ghYItS9x+TSRJVG4N6Gn5Ynq
O17CqJVrjgH8DJ6iruUKdvgtIeDCY0ZN+JI8bbK2vaOuXWZffKkSyMLrdCehZ5UQZ2XXz1Ov3zN0
g0p7eywLKmvsj7x6mkixmRC1VM6Z9syiWYQEKQiOoQC9jEByQlqSHxLesfk09Pmv9vw9vQw9niwj
JKDKJe+040IxsNMOndHqkKUzmhGFjnULg+caIMldO5KkLJvJdrwOAyGcFBAN0XwXYdgrgsgtWa+t
4nX+b8YCfHa7R/6uF+6hmEpFkAQS0IIx6w0jYXofa+K0E4v/pFE3xLDy2vrbj5Vghd9Gv0eUBjpO
t0gRNHfSaBmOIFxsmsmIg/Hq9woaWtQLIvVdxelb8NjGWNeJ+QpositK3t2djkwc+fkBdOlnooTY
kEJN7Kxi4+RZ2SfUdEF61XeAg0si8pgqs8o3c+jOGL3S5MQpX2gV7FLcnxcd6G6dFqkKTGIjx3gI
S4ysXu1KMWKEjcr5iTV/Iz0fqat911acMcgY31kt+UV6z1VMyeunMHRGIFvUtYhU6ULgcdmHGbQp
8oILz9CrNSzvmhn/3R66oXBjkxzkfiSRuJCLGg0bsNw3yQ0EsPd8cw8BhzcSkk5vraWAPKtf5J7p
+tgKWlOGJedpANvKjkcljwKLQfS9/hCaQ2RfD1Mp6MxKhTBUTxTjafsdr7FjUtaauZ8a8y8Pvwl4
VbCnxbuyPXupB47TH0L5gufHpqNqtNGGC+aNymLCsvJqNKX6UuDir4yipzF4iWvwvn1NVm7w1qMW
e4aMyRngFVGJOT+vylbeThFjJ9luuDnfWUOloMM09mHRegiAgB+bsDlAi/HsbDYgHQdX9gLeqg8Q
cKnvatNC+1laHCk5ICYa8OVI9eHt8GwgbfcA2B5cUv9782PQh72UVH8ZuGSEEERKrDufkG0ooOuS
S8jLzObcaxEzznj31VqUzTbVa/7W/yuR9oj9nPuVC3P2Fr2uBtVkq8WhJhsc/2zq0QpjuFz6GsnE
BCjVLFqYm4Y1BPdjOQ3njTr4JrUPdOcV5P9LqZhfTYlmkveaBasdUG43TcaccGsP0RikE7nbujL4
CWJIfypeUC+30tXaBbaWKsC1sJEl/c7dbS0p9+xocOktBm8TDfGH8JBOu6b3B2SvEXqL74uWx/DY
ifglzz4qWttQ76YV4f0QxZuyN50ATHz68kCgBQU88Cu0spMK2Hkq71gvFjHo2HYyjXycn6PLmE6X
XZrenmLxrZsDbOSZUPlmV4f+8Wts2fDk82OVWMgwF+CrsSPDKTUcyJvc5cmtWd9O1ux+RnS6yG8K
k0AwdAteK2UdTSo9XNmSqow5L/+8SOJ3A2uVwG6kXOwztVRdmS4vF94rbaMFQu9VxmbNf8ShINqd
t2nId7dmD4x4s8NuRPzvPNyahApzwhZkSNbJrFPEDxHRNehnhz/SFufFyHaXmyS9rSBeezeVeeLq
Eiq2GSBUXTm3CjErP1/lwSKcg80dzis2cVul9sZDzQTiXKnM4CYwNp7MxJBQZ2zTXlAj6f4HmL7C
oP6Bd1TaZrHbOrN5Jmkt/BNDmlRIW0xTekldSyLYa2tMor1JHz3KT09Jm9NSCRKIuZXNHUzUQ+uk
fLelh0j3RnNFeblLAo5l03EkxeZfwvm4HE9aopGimsmZBNFxIBD1xmpFv1c0EdRrNMUoo28iIypR
AWhjJ+QYhf92+Jmt7yfMToT0k6zjA63vbQ4sklF3TewNIIehrVUHQF06K/PnjNQaS5+jXYhOSo5t
B1Wh3d70gRX32Ppit3KId0wGKXFJzn0yDoVP/QzMKUXsn9lE+enXwZ8oGtB0wuz7HLFHiTedYxYn
bGsQG2hQnao/SzAVgveAdP+415Ms7+FIENGGioz5F5ifreNv7mASW7nJiBe/PheIaeXCu4VXJh3Q
/81JAnXDKA+XJ7xtfwHE8VuH3Z8+tRt01V08wJvMNbraOlPX240k9kQX5ODWG5ySwNSyKj4I5YpT
QA7WVTykdI/KXx1H4XBxlgbRT9EK27FT0/qQm/RQCz1NKofklT7i+10sOwAOKCxVuURA9MuTqpTb
UD9bicRpJHmgKAZsPuzkENfesdNKAT6htbm3SfxHhHCoJYD6S3BeUBkbHyX7fLfxrFyW7o8RKXQZ
aBCWzB/0IQPKpQXDWfFzgHqFPrYwEhlsHfmGiQUOvDF5Bog3l5lN9FKYh6i+9HZN2PTKrfbItyFJ
7EE1ddd/yZvxBoS9OhFvorPngv+NSgnZeHKp8sTKXXXaf5uCQYWyr4jK60hSB9IFvs1rp4hii2bd
rYafHbnUYUWUwtGKRZxxbvSEDx4sbtiNBQI8R4XxCugDjJFKKPa3uvKNlxTDlEVmnZ+tZGuFHJ7r
/lo+YlWhhxTdQL3n+nDnETUCHQgXlnf9NWGiPBHVEYahwQbbpCn7Mm67jDpEAKK1cQLwI8QostOe
AZUxymwqsyLctUAkpH2NsC50CcbQAF2eLBizHeHN6PrBuf8uHEMEBPtsW1KwhNe8LiKLi6bhmIzb
r3cGBGNvdOHJJmp9xPjp2wjvKd+QaX+UwLT22CJ12Surh/3C226YkHbQe5CRMZHz9OLeVgW1dH9h
lsOr/I4kKuEHWeZD55WUuiytVmLhe11Yu8L/bND6HbQevUBsHnFeRczr9rWUTqY0bii/lSnID/UJ
j8fP8XIbiJuZVKKMVnSSMKchuk8UmEKVhFcjTTyAFcSic+wtYc2/e0IByM2+8F4pt/2msXWuBjU1
5TpqFxt3v5i1IXNG8amkfHdszL3tgB/zaSWO/Y9QcRP/DjYZG1+lb7q6vUKRdeie7fKWJFt77X5m
Xa/jncRaufnaTcX3WshZFiws3znkBxgQn7BkEtr+79uDFmr44O78xACXuzYbhLauqShobm+GhWUW
TbCDi5q+h+R8K0kMJNLNE2iGoVeOU8L2s4VKPzHkDh1iVyU5pdYnlv2i7Df26BDI8eyhV3kY33hL
TBJalSDcb16vEoQOKhMdk+5/QVxNk2ChOmUZ+MBIbgUz5r6DHtO1a3t3CUdVJqE2Apu9zeU1Apl0
0fJGl5U539yNrYK1AV3pKiOZu319iFDdWNO2PRsMxXmMLkm4ahSQNZupdInl8qk7OuDz5xX+oQqo
bgZBWco6y0lapTs8gM85ImZdse4PtRRS5mXOsIXbprk+6kUQ+vEOpFEzgjTDv4qWJuxcMFS0dVt9
hl/CEXr3FPl0lr+wfu+Cly+Nnb6ZzMRe7z4ToZYltSiFzD8LTRzZGCIrsEQoh3h2UZVJLpNnaSi6
90u8cXntr/KZg6mEJnaNVk7TaWZsFcf7hGrX7yGedXaWYg5m2AMlBDJxJ7XdY63b1yR1VkrVggz8
ftRX+Rbvo2DMbdPIYpAx2NUVVm6vwktRyLLSWRQkQCDlfsg3smpjH1F3pwfA5Tei0O2Y67JVa7xn
V7UgaBpgUFXrxRg4wMmP/2FZIXUQZ5at4hyZlPE5hsMYxTj/RpSK9eGBqwICK1k2di+469mB92YE
xu4wBZDVp4tVs7l6+FiEH1/pPbAkzgRX+vfsxi7Myj5FDTy6+9YYcUfrxBwJg7u4bijRKkZCGuEK
ijZ5ROLPn5x5bxjlQ0uKPq2AHiExRuCTISQ9KFrNOZscIGiKCCrfhVMHzvh+yvEfBLd2Fn5EpScA
TeUkNZxaEkLBZwh0/Ntj+2CjElkr1PwH9OfFkSNxmZtYQQVKyJ80XlSh2Pv9PQSSRinmEadzgBTd
fDTI7bPaXeFvRzUABdPgLLt6n2tc3KssVWKIKOTLQA9kOs548VyhjzG7x7ee4tAV4EFh/FMYrwU5
4keGUJazYpeDiUbagaxVX+onGqlEzIYl3DW9xx+tdi7kNjZRVltoudgFakRapp3bQB9dqJiro8z0
w+XfBpNN1jO5e7SnBbGTg5O5x0Q5BMw9vB6TYDZq7nJmmJOyswv0o/EGPqT7Q4i/5exn1ZxtPLq+
XlNm5ZoXgWX/FbWDd+IYGCYHyVCG90n1aZ+8qm8e/hrWaaIT5UvIikajwvlvHm8l0dpl64Bs5dMA
GHVM/o+sJHn/wIrRJ58wdUDkt54o12qr74KsmJjCtBYhS0Fc+pZ51bZvHYkgV7mx8C6zJf20r95R
hS+88BI7JR1QbOYosIBykmMPrPNz8e1xwZAxuLddIUFDY1eBKPkqiUyTZ68EsbHdrMr/evRWWWZz
W7w6VplAinjuzxidERCN+thHHt5WF4U4EJJe7Urilwt/pAK3+1rgJ4zkZbgbD3OVJHkJuh9QVtAl
S8OyxhZVxjxyWtDJEQTOJRgke2e0U7HUOmo5V8M8i5SEom35Wszh1vloASCS0tsE7X35wKDb0/9O
qkTkMsJ5i3imTLLcVEhgQS8OPRYOUC3d0i1rWwz/6tLN52xMp2DdJbfghRuVsL3VsFZOFOtAqPYJ
wVuVD/VSSo1IuPK7gPGDvD1QCwP0Kk+lEBpDrSPWlI5BFrMd1lBjltcAU3W0RTmZdyI3N5pb4zjM
N83uIBhTjqRrUtbWr5N1LtSO3k/lZfAwAuN125CIk2Ve5Djn02pqfIj3F+MoNdaWe26MLbzImBrJ
vv1UXCbgSECSBqHl7i0HkqNfUunAwA8geOlydYlVBILgcSvbyjA2/dW4TNhxl3O3s4M/4G3imMwn
lYODZZqRpE3U+XdytdxZ4dV9LJz/96h/cQuM4ncbrGLfoxG1IxAbMnZORiXPke/Ov5y9eLfvxMbV
dnj+ZL4d7TPi81r0fLwx09SfV2zz1VZIsaTWXtZht7juwNf0DN8nYFLM1ToWytWspDtVejMm4zDV
yzz6e/ChX7XY72fUs74xEGey1XTvwvs1QJlYMwjYTPwq1//ydZ5121cAbAjZVLQa7SsOelKfrvSa
gNAq3QkKoEgfdcxq4cBNzwurdvWKH8f6gWCfp0x3g2p1yVhlocEegiM/+nVnraX84HR0yEWbU16e
q9U4ueWaPZvlGNZ/XREs+bs7l4yNr4WzfsixZ4mWu9BhNAQJXCXzZEdOhYSxRW0vZVPAnXD6ITX/
AMs6k540zqwbhzb0E52Gik8voEZftFvyM8HJKVujHDPuOex6Vd1dRk/tSmMTkgS4fIQXywEHFAKQ
8nBnOKebj59CLwVkA3+9CqPnDGvwZN/4VcBrVz+eei/hypB4GYRw0fmLse2qBFmT+bVVhFrYa8KB
RIXDvojrjlBRhM5JTPB3+OjXrZVn6obaKnU2f6y++NVcFMR1WMuHhNOlmYYFWu/TRjoZVZ5/JUWu
bi4LBZtlvsw/fh+CHmNIoEtSchy4HyM+RNE/agW9SIH/K1j1uFHa2JbTuX1mkv5sJPFVfvdZKRyl
Q5lbw0ETZbneeLX2zD9vzjbRFS5NHOl+t9rMjXa8U0oiAI+6Car6ztvRhGUvQt5YYFzQew+cUR0n
lEocqaBQbWPLnz6Tf9uL6Kvl0uYeyO67rK2NWpj1Hy9EPo/NFukHGPl97dEswy++M5BW5sHJzlOt
kt1HkxGbNfiUWylOgiIbB8kj/DRd849R7hMzoWJ8Nn/rGfsCrk0RLhziRT6ZFTH27fR15BFtIFuj
AkTmNBLyjlgSnU4HvrxclmeYJN9mY1Zd4oGiKaIIVtqp+whG0afzP26sckXZXe+2vqZxSkxoggoS
kqwQpZtazMnnR4YylbUjPKAf+FbVjV4cOT6QOIPvoXxb6ThPOIUw2GNK+12b6KB+GWseWTeLqUAy
5fVAmm5Uawnb45BParImh82wbYVr1tLzeoHQMaib9vmpfsgXrb1vGxFghBvOpU465C5zMAURthcr
Fpn0mED26jCdAzvqd8t0yVPl0C4qD5/QtWQjIQOAWdjrECCzy4+NR2tZliGwgx38abK/tAkLsrsf
GrGRcLjgE9YscfSfIjM3jAvmBIwtHStB0Yz0FeJXoE2Rq+yb0T8NXBnLj8oc5tlXw/JnHyE3+CIV
P/ytcPZHw+xivW8VTENTBd9Vz9CSlE5JsYKXzke54yuxLvCMWYnXF4oXgKxNmIpYKVZ1D6VdXasT
F2jRb7sJU8de5TrhK/Dr8hRgCnoam1mXphgr/9xZ0Rnjc/vwKUIcOTcdw3bL/bxtbpEUYEl5mRHg
jcbnuiQleklFOkzZjIduqYWbfTxDFnSkieupVmQYzguM9HNT1WGf7bAdsxGFBYm7Mu2AppuH33Wj
WKPX5gK4P9iqnI6uNyygb9drRH8k0AcrYkHyp4bEz6flC0LFCz61GIHRawM4g2clUIJSA9jEBvO0
PG9047iDIY2/jY+Bhx9x3Qbmw9ertgod8lNZCknQeBBJExHIzoQV80jbCM7eY+WjjxTvvchatN5X
H3Y++MejdnWd53l17qeYq07LhJr32OZdz/aGcq4lAk16DkVnio2o3xa20VQb84ETu+YOUw2TCU7j
rTFzMHevPd5uh9tn4jkCRdt1tUWPSOfT/jplBWR6iNCdpb7kIjjKqANPrARsPFdifLcgw7nTsOGW
Ajb2XZRftzdB3reW/qcTi6sUoq8jOt0qoSe0/XAZ3wVc//UE7UcvBW3l2aFsjxyoUfLKZB5VFysc
+RAibRAxhcmJwVaGcFlAU37ZxqqBzuExkIQLtKVb8rmrpJU+tNzkC0DLzGfu6Qf4mbsnqhUDphqY
Pq8FsiFlhl9jYTcNvAUJKY1Q2KUnaGjJU8f1ZxUw3afG8Qqx8QGLV/nGvgazseRS/25AjHsQC2QG
9gDg9w0am5mx5q2gQFyhHH2KQfaLkkd9pvyRvYKg0rsskCzuiJeYLQF8k8ScLJJtXnrs9nvKZd5g
GcCTtYnYOTtL9FZUHr+rPcUILjM8tWNtNV6Ya0aotfKVDh7PJ30dJG8yIUmzmcAo3cj3WU+4Kk/x
JjzIhIStxCPoKfrQrQ18pJixI8oI8eo3rH+gWoIEz9Ri91sA8LA6JypCY0UyRivT+Qkln5eQ3oiS
c9hnaRghN4Iap5RGi3s7lUpHj176qAM+kbsO5JvUWFGQL1/dljlNXVc0Zh3LPrRUpJ34iigB3aEH
sb6Ktul6xlkIhAr3NftEdw/JaGLVvdm+iZRZ/2ldUJnW+c0hwSUnX+Dx56KnI7GPgYVr6/HKviOU
+gi2YeKrsMQFFxO4LI7ArucFoQpNHU2RBjfk2Iy4lFH9wsC6Bb0egjXEx9oscB9op9G47/6U7E3c
CWfgfYL+EMRxN/5KNknV9IsXktGjWs1maHnpqE5D5sErMoTyKLWCRraoAkZl6NoAObeJ9KT5QFCT
EMKD9jOr2e4kzXqq/0qCoPWUnjkpL+u1lDc28qAP1AD3JFrAny1rS5gvLAJDZym8ZMGS/qktVnFD
FgPc1pm5bD0b9VflApe4fYfc8M9OudMNqKQ8xcELDF1M5ZLADQe8HU+jzgtOwkRaGmdlPZtiYPW8
cYbUY7X4vx+V8MB3UUpP9lNmXYsy3cIv5tKgW4t9lp5TT42D11vXxe+TNPMQNGhJc6iLEUeUlrRZ
ukxpC+Fnt+0/DbIsQ6TsyvY6X7Jz9WU=
`pragma protect end_protected
