`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
giGA109OWTgnmloyaK8oOFmqzonheWp9FFhZykD7eqi1+76ImXNhPe3NaQXpcCe3NaHoR27ZRG6y
K2utGZ+Vz/t183AvBWIBVdXB9lgQ99q/pDNA/5GAfxED9O26mvitPUqKCj6YEr5/LsTR6Ty9XSVk
gjBYYnTPOfzjYjNNp1/3Eb+8c3nRxB9YUbTthAZbP3ZaHP3HVDrjyzg1YcQte4JCbYPHkbvz4L5m
KOHclzKOLT4rwxPvIS22ElVT1mDxlQBzfn3BA7wLJwvAFU4ZDhCkFrNUA9/mNwqWxjVJ2jb56gDW
sE4doIw8ZhB3iWVnKpVfT2MLkzpDgqsT/+MA+gyThK+M+g7yCeNjx8TqQXZp+0GvzNzcV/wndXNb
vp4KjG8Jn39XMvfSiO44iKrkWH2RK+OgjmWyg2kz4xummAyITz/MJPj5fi6b2yk7+IRrHCcKxiol
I4cYz4YeKZOxs0B8F1eerEWi2S9xXhmY89eLFSyxoi3IBQxCW/C4srf0iuME8b9PDiNokgun97pK
t23T4max9jOCXfsCt1kcoXpaQF7Kdv3ULUMvQUIIHb9xvzbH+SaMvFYz/6LphKnb+LixOkMJ9WUQ
LDNOi0rc4wWyKYSDVaqej4AFfiR4dXtX4MEthEBgthLPJi5Uiy6XfYWEGWHm947Qb54xsboJ44PL
nel7lNwn7e2zeYcshcPAKL6RqnhqnDpPCur9ZnpEGiJNGZ1l/gmlLkk3KW0qbNCcCkkuCyXetAsJ
6InaE36jWIj2kEXIParMTJmd3Zb5/wE+1RdZOwd4sjF/pKzsFIzYejfALrksG9J8pgy26Eop1KNU
CBd9p2Ck5VlnfQyf+Z49Vy6ZBSIcxr9caSE8wmoW4+Ho1s8AbuDFHxoQj9tqn4xrfxQw+ZYtjflb
HBpTAZ7zumlvwxsA5t/V1qApDtjym1wSZuRaj186IB7CyjWeJLHHthaD8e/crPqJhTxFiwkqeZGF
mTJPcztJTDvRBtAmltFKJplgDPvQSE5Ko58EzRwIVu1SQeXEbn48PWCOZpamA7GyukkQtZ4rphp9
TWQlhA/4zOuOTUy20H+BygItWl8hFHSrskHPi4Gw0zP3VPkWpUEHzySSPD3cwrpK+75uqYPOfzbx
/S1t4SfjNpFOjhosxNQgfKNkjIUrlbtE3UkeDm85l2hrZeYc1TA50+owvDuLaj8i3U+Im2nvbk2u
kdvMFfnedZ+MzITIENfgskT5InOxLBnwDqKpqPsqCYxjn2Lg6jaiZuk2KNPGqnyaWFxs4stOSfED
jdpsH5E0hwmwfntR91++DeMH5wLuP4fdaIhuOY8WIAYjWkB6jL25D6+nOQw9Sh0m1Q5xJyqw6j27
yMzVEvdPl3/+/Wa9EjDedI137Q1SSxu7r4QV71ewtp9fuDA6yZUd2MJKJr3WCGzGUNkDaT86pMDj
UuiJPcEyOMVDsPAfpJuantOMj4AQKXASjdyypSRcgtzwijTXqbd57IabTMbP2VjRfnnm+uMN8aXE
aFMBFsksyE+SenX71+bWkNWiDlhmr2BnOtr44HPilO9WXx2SoXfSg2kuAwvaNTPoo6cuNv9r2uRp
MHFciNQCWTWM6BxhjhP6r/Kstbs5uBHiMDGGm85HXKvhgFZh6Ogh2XBglHmAaxmvNBBRyxebIsUw
AQ/oLKn5fYrKetvUeIHCUUpfJ+61aV+ij9SQA4MfRdOYKvmUrUaT21KYhIUdNsKKocuy2nUnv3x4
5/AzmkgsGDIu5+t73lLdgiSgzdvnuZa1tNe9XfqR95lc6cpIHXDqc8jc91Pnfc4Nti1W/5vy4UEr
CjPCv/O1NqwWFGmU2c8NyQHddt/SO07U6RtOMSsqBdUb8TFjAOVjqL+f3hj3SqoDCVrouFVnxYlr
rCeO7a/nG7uMq1ZQGnuVmaFGNUVKSJ6/E+g9UvY3k2UOIBAfCW09enQsHTSsok4pFQJY376zAjCK
OgpVhJYflLjc4mlckG9NkS2npJ4bjGmRW+x7SdwXwBo0NGMluGZ7dlRPa3s02Yn1wA9AUV7WMg/X
2cYo6TQF+JBTadVmAwO30Nef1Khl/9IF4yxwwi6L7wYXPnksvcGduUa5EiFCauUg8OZYWL2MnWRd
VEHtDs9eFqtT9H20YS2+1oOtmt3/A8NYH3VMytvaFC+L2rRrrCZMDO+K6mxJTA9ItJu94UvJ3zzD
uptmvBGvaeQMjPLuL6+OSjO34z5ZkR/bZugwmJTWknjCTdw/2/vpeRzJg+v2bfhahHeUb8OlbFk1
T43rvNZO1O5uou8L3Wfh/sRI75pbJlLW2Dy2N+5mnAGQPnSIzIQlMwlG5vVKvoPZ0OpZvxUAO+Og
uWdmIoeUKs7E+eDDtKI9CBLq5Xb+g7MzVpl0Rj3QWriG74bJCNN9q/hhm0419cKrisrn3vOfrh0l
cEXWpppI/Fcr1DgImFDrRn6J8TAWdMg+F8WO/LERtZbWlnXzeq3X8nwwdtwQNGe9rIPTp8pOCFfu
gavW243rBAtkJ5RYx7K5SmUNBxV8k7sSdUSbi6a1kkTg7+QHf7vL9XNOMJ95bytOyvnpyihgQAtV
TrZdvB4CT4R8hfK7bF6UvmLmcQvgn26Wsw7yiWFfFlq3qeV9BrvZeo6yDX1YYOhPu5c1wg3G9WtE
JOxVgxXUy61GzXxyRVxv9D1TBh/iRCQxLLo8mEiDdv+CHenslgdOkvigtjkw4dWTlFZwyzMSVeJF
R0ckXr36XrnZwjGCMEE0O5Poh3HvB9nqhcHQlnmTDG0Xum0LUe0285CJuaeCR3wk0UsxVKkHLoMC
X/mM5Vbc/aYFmNQzkDcgnR2mKWaC47k/u1ojagPEkRFl2HNmMfKuA3P7VqJianciHSxX0xySwjLA
mn2d/1ggKhPOUILTsm/7JLas81jfJpoCq5neCKzQbSTmltD1hzCPLgIviDK2XFMSN3ggieZplczJ
19R+548trD5qgjvF2eS4D5bhrkjIYYQTeigkmSfaWt0qvKsqts8rEzDyMtL/RsSk/QsqCltVwHMy
sPnFtn9P5D66Z3M1Kpc6rVvVu9EXS4rcQLdGNVnbBk9w7pHFiSma3lGnZP61b1JiG5q7bmPFLLmH
vEQyiueOheFHtqFvHLMT0ZhqsofFh5EofbP7GfX8QFRs1HNrzW/DEvFFLtPLxBcUyv5oPvYDeB9S
Rc2JjqLVs+3M2kukwfRg82GdXhbWy6CiNSi4KtypmgUwKUt1xToArDVYW7LIAGs7CGa1K1Y04PVQ
2YNMgMogmmXwb12EWQ+m66lbHWW179I1c26cMCDd4WQB5xIxgEa0EtZAyRC4Pdzt7V+WTScej31A
5axT3nJzsEvoAgzEPJkj1752jYe8rceERbq09dZ20RsJRoisZfsMLMdphsn2RbtYaHiS3S6LRr7f
wrgXXp562g0KVbMm/GXAlahOEBXwyKfV5xgKY29wtiRPRrMzk+TLQdDOD1iGcYF9PHNkThzdJ/+n
4tFu//gscmkhiJ7ZZ3qYT6DBLEEJ5dXg4FPKmkAOcPvt38x6qIFleY6Ax5wyIYqK3+oirtV/Z4T3
9qVmFWO99Lh8j/J1Fh5vUDcbNapwcUeu8GRtYA5uhAPlso+6gYGzzKxPyuQ/gFsMbNaEXUdcl4hG
VfFfjXidiN7UoDRVKEesxPD+2wqwP2n3NfR4pmIG9iVYKOqEW11NyaGyaD0auHFixMKVJ9FaAXKF
152cpMxe6ZfKNZTTkitKqzWkzMARBpC3rrUQU4kt9zrqw+ZINUw+sRKdUQ9stB7lDfoSi+GLrmmp
9KcxUTCBl/ICpEfqVYOS/wHp9GR41FMEDL/PEvQvK/Sw5ZGU22CuEf8Wo8FdhlAFpOWu1gbz8Xce
AvC01P/+ula5ffLCkyO94CtXI3+O7dJhD0hR7XJ6l2F3X5a5JCnT5SG3wzSWQGpC0qideJPOiPTA
iaPdjaBIwv0ueYISl0HSF2k7NUKjey6y41exEXVAsUlMFTpmH9O59nSZiAnHF7fB6r/tQXOFIXU1
x/yU2vRzIaRP3VDeJILdErqeUytPZW9mgiLpOy7rvjOiyQi80YkrDIBJoyeZaxKsj9mGMxCaDhM2
6PXGLTuDUxGek4MleyFbFrw8YT9Xkcb0/BrcM4MqBTf6r8PbpRKPGJARF9RkHkoyy0qlurG+JS4q
Cpn3rwooWRqal7bgOHEyYIU9fxaFHGLxNGAKfOBkcuznebqjYpeS+J18ve2p0wYAlfEcowNEqfwn
fzhLlvJw0hLZj6IP340RDwsPqpAO0vJcC+0QBuLkQl98de1HV7MgHvA367eg+cgW9x5GwuntlMvR
72pnV8kKRfzQSgJozbZEjrKNgWaDovX9x6pMlad5yDaleLJQ8+7dJhZ+ocloL1LYkcFyw4TB8cHl
ksqx/iW0YjK852EpTdC4YuiCJrtiRhcpS0XvknMJChraGAodnmXYWw7JGfS6TijwppgzDzQVirHh
seURhWRV3Zgppfgl4fT+NDeqSX78+C1HWqjtGpQwUoTd5F6Y+kiyB5iK6yg2vfrqfhul4l7oDmqZ
snRtWbJp/X9OHomuGQed4xpYh/KvelUMMAe8BirDHC2JTu4wqqcWUtDIBzcIBeQrt030pPRiy+zd
uogS0Y6thW4CF+ml2yNP/Eo3bSEgD0yz8BkTM7FHLZRelVoCuSQUsisauB1d6MDligDxWRcLjPiz
kz0Dbk3Lva+xOBy36axcaoCijMWJhHZatSjDV9HG1Pw/5bKnFrhi1si1w2rcUFuco5z/5wEBG7pt
R1rTfROGnQedDLRIkmE+rX0KvHcAfkuB/nhAu1lGaibZViUhkZ79/UwE3phbbZugB+YsZ9q7c1RP
S+Q2+gDwZhpJtpomlpVWZWyNviDRFGK5gufT3DDd+yJiFNltlFiuVN+oYJNkE2H6sfGYY+Y+YQf4
ASghqGBNu5g8SPcjb5fVp4lQlU2X3EYLcHNQd7Vi94qAcQZBtAriZtnAjCVNV8NfHWyuXfQLgmYT
6ToEsh2d9uLutDff2nUT5Mi7mAYGTWfmPc99mnmYaWkDjaUMEJ5VCZ2DRtGKmXqU7gLLB9zIPdEj
Enaxe6/nStoeHcqiH9gd80XRyhbtMhM5i9mO2CYmvi7dmir1UFb0TYR36ZcLsXeAjce865w1v28d
MC9Noh72eKaSgQVka/c0dVDLAHDdeNulbCHhjvwnagjhtx0wUBKPN/OVqmdRh2IjN60yTyEVp9t7
RpNi8yBi71xa7JUoB5peMdoL++FtCQeQz92wpE6y7VcFfUQ4U2H1JHGnmit9yELx2WSadUx1uj1W
V0YJjJc5dMUBzaZB9GxxDeNrnYMGI4+U7qRVpLjiOIYmN05MwCxiyEPM3hQXaTKHPIOPD/PiCixi
V3jG4xLvJaynZp7pfbG2EnswD58mEumwE3tAa5TgOB5SseV1rI9+kfvlG42309wbOyDnlDI6lh6X
dJES+eWeGxtxRNc66sVgSJr5YRL8KmpRnbV4XjUScxQ1BIFJEyqT1lrkd8jMZZIXRodJXHioG8Pb
I/OWaHxa3LZqednqZagNr79Yl8excSiZXI6hVzYiLXMZ82B25tW8h67ntrK5wKIdYnRnGFTXlA4q
OFB/Rn0dT6CNpWoyBYzdSYo7UO3I0HyNa0pzn2xx4uy2SiMKWn9L+RviRbJaQSKKvb+OBMylmmyK
AVp18h4HmKWk/aA/9+cd9Af0fhEOp2L61pVtW6piBhu8OPskNba+gTeUFRzMYXpWogXUj6Kfx+g0
Ie/3Txn6L6CbTDJ05NGQyWOMS5Jx6nBNwc+qinftBj2sTPJYyKnm+LfKSBcqnMvzqFjZzK9vRL5x
jibiG63+kYr+XntLBputt9ualcIZj0vxhpE0gKiPtb5ACj9rMHGjnvzP330QQRCEj6rdMWHIWYl/
1ZQhKbbpeI3YzavI12Fi1Yrrnh+eraSK9LCnWbmkISWsn1rxhthUKTKUrKzBKg4QCn+KRd+iOGQ8
DEbfxz+O2o/bdmP+INxFD0Ps8Qk50b5EOBm0Yd1wdtaaYn/e9csD0N5cbeDWymhcSZU7fOA9sKtS
kOkGjiToOS/vLCDboldhJQgwOxe+0dRM6Fg4UY4arOOQne93ow7DEChmHEsVVLshnXNN5Y22JWHT
+ADtKkUZBWkEP3grWP+Dk8M0M6J/CJRI7PldQP3jIdr1tH4c+GzRXoK+YJexP8ril9enNybMCwLE
gSB1R3XUd92N27NMXDuDmzFKmZF2dGybihqjzlWtbapTggWGtgJnDxUnpigQ8BiJMErMvEDIWGa8
yUM+IUPIW5rw9rsjJlSbKcBKf5EdgUy4gV9FvtrQCHXWmtHElKcNRUgQhZ6Wy6Kr142g/+BA6UAc
6SyD7ucbVRXqcB+b4AoLEOm7SlolpNZVIPbAPOTgryOgsb2Kb7l+TYcE/KMOIGCHYwvBHfwvI7gk
5sSn9Ma8sGoES5YVzP5Cc0nGoI3Wz82SlcaGeJvzTCM9s0kURDazAUpybwgqS4aSzKraguQIvRYx
ERg8HfwBP69c1QsTMLGXr1MmRCpxDIGt2rfDoxz+qElsGGTcihKXcoTQOCGOoJNqaW4eOTVphfeh
otPLOUzuA9Jd1DRS3M1ZGryAk8nu+VRdv/6kArPSVZvSLhQgsqhi5qPGPp9yH6J4vszf9PvsrVzY
t3noU0fMDFkerVXSbEIuNOvdQ2XIcnzG98uQK2Gemc2RER7AGjRaSz/GATLui83rhy7eAkgcxbBp
peG42oIDeh5qHzxHongJJ745hYo15PYTP+MGMWbJ2VlIL2H1M7L5TU/FFUhmjeQIv7OSCSfrCoc0
wTfxjExEeiSTG0ykfjSok2TXfKvo8qQ3hhOGcvM+pTzVP/eJecwva3NLEDTj/7qXoyUARGo4hkME
xNGTzUobKZ65nQNDhpBrkbIbW52a1wRHmEntvivdChL2fxENKXuJLjWu0s6hToMwJQipoQ6YdauL
s1FekWLGN6zkOqShSHPAPVVEG1kb5D9P37yi786h7hE6udwnYygj5W+/NPykblulxBrgqlfiw/Nr
aPvFUToO3T6mG+8r9SPYlJjapzgyn1nGUFnBxP2nwR2UAWrcmJJc1uD9MEjgKn3VqA7dhXE7TTP+
5qzpwBlg/LVKpV0u8/ntiFwrXL8j05MyJCfEuA47Nd4W2/fBXIyDMNbUl7+FxoETb81AXMovOJhu
knOSRuAXb4tYrK449plj2barXpGaVvKUZN4qqm7xK5r6jIhM2R/robWKrBxjbZ9qNQCZ2k0/jAlD
qn1bVGccZNwWYVPLDrM6uZzirRI6D3AIJxQ2vWO+MK0DSfz2vX5uW4qR0T7zyZbOTWemyyTib1/T
/05rtZBFulee2KhWKT9cmf1WldMvnvCQ56WCcplQHNuTQhawpqASBYMWMdAamRODv+wiDxkhxjDm
VtqlLAs3Il7Ce2biM9vVRPXGHZrxowUrvcgxZ62D+YwIZQQhNljV9pBAw4D5gAX1nrnPzG/Vy8fY
f6mINPA=
`pragma protect end_protected
