`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13936)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vHvH
4U8dDqu02lHqx1v3Agq3S014dUO5JB3io4b7u+E1DXTwTlL/CmbkpmLpeDiwXhGiTlQwaKmxId0h
RQayIrxzA6pyd0kEwRSH9lJ7y1fW9QD+GpNsiJGaXPF1VqApsM0OTSqissRvNtKUc1ejhztfVpz6
w4jjfTf5b4cH/UvAabOK1fpErYan+dQcFJiCgRCA8sjHXizFDKZWr9n//hNNrUgj39Ub8bnDDexg
AdCtToLcQ7bjuDtGloQs1qsppFvEL6+/+6uEscnzyoXmWFW5ChI6/xycx3gkOT4UoqGBCaGvnkct
iMEMWpTNGY74AJTkesj7oEBJYE7znu/EuTC+DTnM4a70BETER1rNiAJEBTrYm10PSgwFpHcCUpj2
75nXZX64zuIeShCtf/7RaruD6B3w0JHB7i8DnNY7GkkqGKaGRoc1Ws8iLvAo+XI3mLmAqGOc/mzO
qY5TTFqy0glZMBJfB8MfuDm8gt/TlL2G/WU9ochDNei4AKS/drI+twQN6AZHztVZ4QiBkJ31+kbE
pTJOtDIHti/xKZrWBqTANq6Eynhzd37Y0rmADy3WQO1FcXy5OeLNbBKmCmw/it1+qxIvu4R1e7aD
S4Zv3wBVtawdA7+awZwSt5d/gC2zkNrd4ccYBBDWuZ8iTa13CmS+Dc5RDSkfRqhmYn6pZqhl+68/
ixFz5mn7nKQeHYGnJdaa5sPDRJCV2NAid+aaf2bU6ICeKgTCTd3WBWOPZfZ/M02gXADvA0cHukYP
BW/La+bvuyOPhbRRdf9EQcx6gUNbTuLWociUVgk9u3bfpTsOQJumG/2FyYbwjr8qadLiwxFVNOgP
0pMs2lJfN7W8EM2H7IPrbzhN7pB36t/+ymWGsBovNrw7gLYuMWNIxplXi8bjYZQZDjYVBBwogckN
oI7elFPPXLiSzfxuX4PKsPo2vgqjmWTv52RHlFoDm4NNbmTrGkho/x+6H/voDMFn06MySj0M/ExK
5vPahEBorI2O7KKYE4lIQIquXhc1Zq2zfmGepurz64LBvgEtIeR7NckS9iwMsYEw0dQyY9XxJOKu
HNff3eNPRpfUMat1y3NunilEbOGz8Z28FXndZ7XKHPdAKZr1ZhC+rPkUHk+z1y/HTIPh5XApx2p3
XFdqsvvfEgJ4qgAqXNWrs0ymfGL7Wd4/BB/h6OwJL0GjfRm8+RcuFeZ4TYN1OQ312WxrvT8aTDBc
Q3sUx9Id1sX1bhK/15mdDM6DMCFkf0Mlc/0MvTZqN9caLQUR82g9bu+LNKaRFjycG61QuSCzytZa
WnoZdzaIPQ62iq5ualfNmg+WLuTsNSiUwmpcKd2L6py+DH2wV3/ttlhrxMwyZocHOjB+BVHDDxj+
ci3geWUCyUokwJvVC8ib1u5w5Fe/FYkEDPncmRKrmo8ErLgMwq8OkgUsZhcEBlP9gYN2qUZofGL4
NJaneQ46OgMjJOs7ivNp2dwamP7sv5eozm+wgayEF6pV/CUML3mCHKMv6dTShfsTdsxGeOOTHMjy
TsNg8UO13tsKANZS2sI8E0WfZ6yZvUemdu4lzIfGVS+09f1dctX6Sr0kFZEL2LsrYI9JcpwtoZvz
1qzQvwh4ihPqLo7c5kzjUDeQhf8yfHRoIJFNNYp9qLwEBHm4O+yjD5W02hLm9QcwJR0d458+Ym3+
9spfQbf+LHDn2ch88DZhyNraL1g2M7oxvTEg5lMXgJYsiYwDIJpUtCfAHkdIHZQ2TNB5DJC+WW83
V1egQIzJeLdXtiKux/yTDRerz7e7e1k3ZtY33rCYEvz2yEGWP1tGBfO0/ZbTwPS6EZ004bA+eyO+
NVa1SyCC6LZC9gbAHT6C+UjC47Y1/QtJP3K8c1vW8WUC7QszmYFpp/JepGPk8z7P8nWiSD2abSxy
9HsE3PFjtQVJYIFKdKL4HjGWzTT1ik8i0YsBpRe3SsiaQ/IgX/IXnIZzxfyk5pHThflnIo1cQdpL
yR18Ytbui7QT+U49HiulBaWeJSyY/oge+3kWoGuz+JQgeZfghpmVowuQ1BOhA8vrUHXWE/eoC+E0
s2e8heIaEMMQT7nEGXMoOoMta7vWbtQ1rX1r5/598UW61IfU0Tozx+c9gJ2zD7z4ludZRcngVVUV
cC2RNyZRhwqKzg3rnPPT8e4gxnoPghM5PrU4zRbYXO+TOBJ/tTrzdbWPpN56qirbH+6bpa1ostEp
ACT+lkQzxd50p8nZoIHl4pLefbYLCjWodA+rprr+fEkYSG/cUEGtuhC2YyNZX17kj6QIB2orKfkS
5uYeVfuj7rXQbftS6PsloE2SruW3UHfOB3vy9HdZGttb6uPUgIaAqvivtBJNrQ1GIonz6OLg4mIT
HI7ns2K4OYSEcTIA8aBgPhAfOVgjljJSjVvA5wuSF2P6oFvVgZw6H9cYsxmLRNk3RiGa/ZnqvvSn
7gSYK8JhzCkgBgDQlV+Ih6BLhhExHwc8uxJ7AQqr20fPRzARRIUftXw8rkzYTzZb6l74W8SAUNRf
vFtSvgaVlm1OZpKHU8zYnAih+2AsXq580ffL0xbavWcXxm44xIRuQ4t+w+JyMl9p7oDJU8HpVnMy
tedQ/mfaZKmGK6CFSaBSkQqBKlaEJnQ/Qz4zcJNHxQeC8T7GFqMF7dJgXMrBky3m+Wzfa3147QY2
SE/JtQxpzpr0DE91ZQcNAUXuTQSzgfVEZ/09bh1EFNvy4MHGx5fNDtAPNd2Dj2Mm6fTOLkeZaykQ
flQWe4xwawSWAQZwFB4wDPx9OrREDfXwZMFXjXh9YhBcDEfgcuf7rwFEA4J0hVmj0XZymQDryhVA
ELmhGu2cJzjOfGt3JjvWGsFuz6hSS9FYcwIrm9hqCMHK7g8sbjyshdiQURWaCZBPEBaAmyC1B1/0
aDiuXOqF2vvrsVjwX7RuP4szUE/2Umx3gz+YpyDWs7B8rBBI4VjRcBeyMyQtX0k/Q80lSFyhQBT/
nW6tfsEsFF+0kGDm8FWQlJrvobb7Ec+HYh57uMW6K5yV1d46NvZ63rFu6J/e1PzRO0TlPGYIS55O
R3ZICtp//QRuF3DuhwvUCR5TsiUCnpzD/2jhNHphavxxrRR+HO+AoaTYzr0gCu/uZ0P6qWYmBEjF
54oDtA1FhJ0KE/Vft+fvw0HrqVC5OLlao/EidGbVAsXtU6S2K2Pjeh4ajnQ7NN0+zFuF89yhuiPT
WgXZf/I7xyZdOxfZR0mhG1iIcHzPPpbdXhPtu2rZ9n/Fc6Pv1nQKk3WIKGsbXBxWfOGRgY4HGdpz
lReOssMld58Iy5t4erRckMZozyWk6cbPNa8sq1HW41kB4SHHSbr2pvIPelrDzLlKSZ9G60pVfZyH
3dR9PQaZeZu6CzZHeclv5YCnIOTlHsSGs8iKU9Uph65ecuuExYnraLt+Ba6RwmYDlsNNhOIIdc5R
ST7E+gONDLaaVzoDkbFDBfz7IP+vXYjBKWsVMbU3OP4msubK3IBmLMki5LpmRmHCUd2guamMGpRW
4HchNIN2qWrknLSJzEvuQocU2CNwQ1DyNNeeHGUbH1Y589bpj4QBjtlaAHGjSYtOhKifO11/5k2E
QNjclR4xGZAY2aRhm4YtCPWMdkdxe9P/us2FWoacMK+nr0UfvQDucrmm9VMcfQVmEymSjZv9D9Nk
MdlKWNaFbuAas9hIrYkGEibjTAqMYVLbf5woS1CcZsU5v4Ir4XHEujuk8+WRQJuMcURiybIf+WPD
ftOElNSwoCcAv2D7OelJaDg43Ro0mBhGnpLvF46ZAFDJ/zhJsH0axXqt9gi7QPHUqHBecK077G4a
cZBvmjp9gRdGOOG7JPJWlyqWawwah6tCZFpl66kyize3JAyDLw93SDJDw7HHImeX5UsJqYNz9IcY
pa33yRf7BvCz/LCPIBtVpLaJjZRD3M0R63eJcjo9HEPwCsG6uAxZRV0fCg/qvRqYZDWFa87y2S4v
soibefPDge+cZ3PlHjnoCJ8qhqUcb5V9KOgqOZ8s49fYESQKsFnaSa57TFyTIQ2RsSqrVOXkLPOk
JYPvqkwAyG1kDki4jivRZK5ansT70BgJlM1LQYbFCLeEtPId8/8LZe728/DZ9EsqJnly7k6I2FOP
q0ZtMDT436/xXz2kflaDGVPMBz/9VAHcBzr7NpDTUocJEa/QuEVR9EABwCPNaz/NLGUc2LX6bXky
962qLuTs1cGH+zRH53dXv8FcExO4fZWadARrHNYPrZZukER8rV74FDm/RU+uduh/Tfut8TK3avy7
/6jbzgngAYzq8q+UFOQ4VQAE5ZDjQHZmlfTlCs5v0suJec3UBWhdSCn9KSy9RArNXoLaA+LRyS3i
W/bzEScbijmbmP5o+A0su9qggp1xevyVbwn32xXoodL436Iml/nPO7ZEdHXwUTe5HLw7Wuv9o0IB
q+uymKqpNDNw0BsFjUPJXL66HaKqC3eOHgQoD60LikkEvF5XouRoVOnCFUhArnxnsYLahWY6Dzvl
lO7ZdsD8JEdOuhOT7tQ81lnNWNTT0yTj1qPfcmy/Ijkm4L/rcFwdmSRgb65Q+ApcT5Rue5Zm4q0p
RQ0qnvB3Cy7dE5aeb13Fvl0uAbD/EkwCfCS8JB/yrWliTdJbF+E+eR8MlslLjflWJk7rHzPkKjbT
aZ6k99tKU6hv09WMC/eD3ox5EeVQhNyzxn/BNrCEWHiGvpgkJ/bL0X97349ZE8vu1Vqb+Nt8KiNQ
fuja+3jxmEvPMsAnPo2RTlLhKtZzlQlQT2NJJFhOGosE1oOQAHP+cmqNncfwqlbt8MwQnFL0VgGQ
+FuJeOaVuqlrXxACmPAE6TmvFQvOdLIO6hLNsOaCir763gUzI5hfkUKFBKHri+0V5qb/sMG00U7c
uNyUTqc/ogpcFxTWo73ePMNLmTDSVtzDu6Zxp9BPiCmIk4bNYQOovhvm56Do1etermMVhOzUz7Tu
uc6hk6RR4qIuO8sOIyJzTm33gm6m5uaJWsp9ijusrFAcSxSwd9vE5gYlFYuhtk1VdBYxynhLZMXI
l5fbmbWmQrpiAxEE9D6MqNdjPPyhg4fM7A0B/mpDfOp0EqNfmaHwbJihQDJ+DWWP6XEla4mo6/O2
SRzwt+wjVi961Z1nsuIdmtnAH9dzHhWJMUq5cWxhdvKXcVBNtTIgzxlw6gWIypuFHuBeCpACSMwp
QrZ0q+dZd2liR5bcUvt7AvV/U1s3ruhJuAOtvJZUSpRBXMZVoWRLLjXMlfBqaOMY04H/ErjBpYbD
LwQmddnqISPO/abigqh0X7Y/u+BnBxwo3WwzFy57YlM4Y9elhRUge16RVDC0B6iW0fP/XMAlyPMI
xvg//2R+ZSCMLBpN1iJDTd4nbNbGEaIPJN/CC1CtRh0B9cAZgrJHAANwOhnLjhjnntxqah0nLrUQ
TghvK6b62jtvtQexvbpVvfWukn1czkhDMQP1rJCk+JXgpxN8KqupFQ7Xw7wDX2+CchRDz3S2wOli
O1CcCayUWrIEBo4wHOKfpNKyI1HMVW3CfeiBD1DkL8+c1UjTXI8Ai54rzXGrmghGI9PD14Xwg2cs
r5yN51NfPT6DELvXJiwYbB3sRkJc3OW/w8trcEkmpOu2cXg+IViimAFiDsleo2ERQH65dRvQYOz1
+7aKF3EFZhuXoZ3DAUFoCNBCuOAimWaNsz+6q/3tTWq65R2iqU/7npZpXWX3ol174EYFnP6AhZfk
gU/l/Pm/r1AEJ/oQ8Q9EObBkGcUr1GFAgqxdCIG8PK8HBp1wVo0qk+s4mFWFXk+WisYz2eWiri0t
QsIK5Km2co2hKrDtlvnXzo41ysCpWv7G0YJBaOtF7SJAQFVK6hEGxP9EpxK20iLPL0VXx9GmSpfe
FlglU5kEflmZisMBOZF4Oc5CC9q5lieZqx+7AfW2WP26TsJh4pwo6aDI2iX+V9ILG2zUGAa5q3YK
cNe+w8Q0+KjzQKNpY5Ucun04goSFuTb6n8VFWMsMOPaprjdub7gZf3r5osKBmTWY5AMo1FoHw1r5
RB4VcXeLhVa2aNMmEUVoGptP2QIwjRDd95joTnlEzM01fFwMPg4jYdjG98SXDO7kHJPs+Prq+dhu
V3w0PzvnMmoQmAB7Bi7o63dQ5F0/s3ZkRNdtRSaXZHPRq3FO7rwcdWv9zTjcenlQIQiCT8pfz+dz
gq8V97glWq4+WAYgRCqRqzHBs6Yri9H/Y7JpMhwdjZr/t0Q2fz0Ud19Oy0XdlMhjDnxfPeExwUCq
8I2DV/5K0lo3LLQy9vKz45gAheO5RVyE9qZTmU86GHSzNAPRWL2YEub017GuqGyHq18d+oa7cWuw
iirmDP/d+9JtlVmwrnpwdM7Ycbdh3jReJlwS/7OxnYIVQnhXFek+lbPJz6axTX5ROPqCqaj4Kta5
vOZGrCZc8jsW37LkEXYoUOgcGVKM1xUvR6cEHU1F770Fz69QiOxUyihdeqZ/5iSokj34tNVNxfna
IwvPscMysAio3lZB4qBhHxPojkW6QJ5EvUJGGXmJ3yrrr5SfVmaZRIxWvfBwBDxBa1aM/EjHKe4D
QtPXPorjaKA3VK1FI+JnvxbQ7JDIjwsvRFi1FhxsZ6oW8oMFaOVvo2ud2DdCn36KMv7FgAKNeqYK
EjgmZliftWkeeCEHjn4XsiNXqcWLdTW6Sf0yQsOUmJjRESJP0jWUk4mVJD5FhI9awlKnnHkwOf04
Xgq9Hek2eqPG8QEguVut6i5W/6DYia9eFPP2c+iFQ0hA8cYyIbZDo7YoNyxXXwV4V8Q2n4B+NbYO
OqSJCLiz8vJoct9Y1HLSuhMSStSuMl8WMdEr1QJ14tTpdOUsEu6J1BjLLBBnNch623HCvBNdiOx+
OAcgeHYjW017uZdox5H1Wz2TUrOQREZJFgSO0NFg5iRD95mZJXhoCcF/rUcuQZhQ1hxiYgk9aLcj
bwxcWqXSoox8GipgoENUTTTRK1ILawAHY/NexRJrQ8234tf6DA54YFetk4dbiYDrxdXjAYeb5P5N
DglZww41dbz+05gDCzyTg4824Z8nf8OTZIpulOODUFVo+R9v8vNIsfucEDJOlmtB7WvIJddrZiYJ
1Ava74gzOzvbhp28vaMlYgz6HbIyzf3j02QJallnfksM8X9NIhSvZHWCjVyK0UyiQoB66oH/qnuC
wMUA1i8OB0v30fhkbacjOSgD9VgLTR9TH7kOWdJDtRE+gJVs2vmgvYnUqLIhtrAfTFidP88dp1dA
Fbjtt8UeE17vGrQFo921AFDrbdEDSt3/F7vBIbspNPa+SvMJ2sKBAOpxfSv7U/o/UV1jmbYPj2MS
w8ie0nGvxePC7V54M7fQll3jmhZXkGO9gqVDvXiQhigcfxZ5Cpbb9XOcg7ILK5fG0haKBRo6JPmJ
YjRxQGl8Y5LuULCoxcmc6iifpbG/nazrT/u9yjhBBkvComtf1g2s1Nde/WUWAURTgo6YgLSd1TmL
HZ5W1XwOSNCHmLhvhbR4VrP0MHhDP7iDP04Y3UBVUZaKkb673xrTCc0qPxHkGiyFO7gW7xJ5WP+J
Gjfzmv3c+B+T0sJQja523seFRw57SWsxz3sQVX2n2URtPxWLyagGs5+Adzhjmu1ouijUgtZVTj7i
+80vW5imKF18C65W9YWygSjP2Ed9Ri2dSviRbPGvrmcV4MQxJ/skE88QHMazap27Ti/bo3NPEWma
C/Ci7AZnnVRxXw5qp4UMEd2gC8bp8PbU+ToLU9eyNmUQK/MfJwS405porDehgcjN7GZHAfHUjHP8
qUN2HpgOLEMhXb3R6o3yte0LH1pa3f9WlNgPrS4J41ZSwwrxhnpiiI81Cu9l7KlKXCNGbzznUiBK
PTDfzypVvwsrFc6X6gr//xg5N/0shCfwYqtITdgGF5nVE9M0kfqRgsa/XRmr5wTH7LEHlKi4jL85
+FtdLup6IaHJ0wY6WAsC03bmNVOcAacSscYgE+qjOrDd/+eKoNmODr3kP3GKTIOCf6iPz2QO+KQC
IuYw5F6ieNxKObSlHsK2CM+v+DuW1DM/wo9Sx4rlLujo5TyWBZIfhyJ8NOLDYc9Vxqspc2K/Xzd3
dfuQ9PWQYq+tL4pAcA2gR0bQ5pIlnn3XE9NInLCzoj6J+EC3k5+pYPWekLXM/T4Iu415O+4N5yQf
Ov/kFKBWZhkXaOX1h4n6X0JXl7pdU0QvIoHye2ZilhiGdLMMPJPhGm4fpAy9t8x2LrdN9D7I4KhR
rXv3dqqEpeS0dPj4agHeknpzVpNO7y6sW+0kX0d/jrxoj2p7eAPj5WoskBhHw+kbm5nFtqWYtmEP
uQG/45KoZHNxe0h2wwgrDrYvuRlUpBcDF2biKEfIbvEnKnwt1RhJjjTNfNuOEkxcy4mRN9Zzc05P
gqL7hN3p03C8NPMLR7oqqwBmAkIF+fTcEYihBnM39s4ADRzy+NFQB1lTAGmFQvFzDjLmcxWlEOps
LFBIXTvkaCS+iuMbFwJs01pV/UvqIuNq46HUcBXprL4z19gXvzh4q/Ma/fdNmFpOq8/uY/bBBxKY
nvep3gIfmdo4RJuIx6aNq0BXuBx2OQXpdZ49mlfiq89hcg65SGaKVbaQetrQBnE5/jsRLnHaq+vQ
qS6lvaVUrtffArtChe7UpiymlkeVEXnryqbRgbqOVGXfegRxWCxbVe07uFxok3rLSlTRac+gt/Fr
Nvw6QBOQKy9GEv5pptiJy0pyvu+pu6i1xGKuEZxXhivQ/y6lGamZ7DEcwdvJwC60E5UwckDJEE0S
x9G4iPEQw5J+aLSChSpRqFJ5Bg5nP7DRTL08v6laJ4kbgL3x93LnxOgjnyR7i6XA0J4OTOkKKpbP
7jwhhC0cyihyi3k9csHQOSeNu7CEBy3d6rNtuMNshHSDIP/RwYj4o1sUoWUTQjWy0Kirtl/SHOFa
sCOvFGib3lagExVL20mXmcqrkMwaxBM5Ba++SMNDmeh7KibTaECKEkR85LMsp/JMrqB4WH4tHFOm
IiAFvEc80FF0DJzWv7AVb65bTqC1zAl03d0Fjv++iqSIXCfWdG62uRhFImiJvPPvuQBKfh/npKL7
4dxjjOSYSaqDc80qlLGtWpOkUKIe4L/TAEyMN/Y3FNIc6TTuvKXjqB3On62k2/ovyDaXY7IyE9U7
LOirz5yIwfHR2OGa0E/XF2mps8sr/+pe+o2BbykqUJldlaoBQXrPUw1Mc25e7p6YOSrCQD9iOPp5
0HcVEGKzeuxBURecaEmgvuJ2FK3sVS5hIAOhGftoNEczN0g626RT7jpDvJ86k0HriKLKPm57Atii
voR75sStxKm8Nw87X12XfdU03q1evDMCVpUmz5sdomJs8qraQTunxOzsPCr9/aTQZCrwmdCsDfx6
1dfVDhZi5ISFHLzyLi+NWUfj2eqScuoOVEjnxHqDQzPs9YWCJZxwl9TSIPkYskNbJVt9ktUxxB2x
m8h0YI/QYaFDLGCXDw0sBdFGi9XWn2CDCTvEuq4szwb8hzQCcWA+vK46CU8oHuRSopc41fzwgCic
hOSUPoA4sPuNDilJHnFhZRcaCcu3JNb0z3505BybQrvQM3G8DbH5RmoFV2YqLvenCw1SJXAFeFd0
QQsAXlVWtYL1Xiprz21MhqKUvkU58NTP++yZgxCxPrJKfomqSsAwYaQAsIuFHIFy1zU8o0k3zNI4
I2wajzpAFjNHWy7gSn4bB2XFes7yr0JZOxaRTXRmrxSueXL/9f4Kkc+6gMwQRsgkKlyOj9ipjceu
Ejs2GenrthHUibwSJZpZOraiC6Q9jHXWBTCrIA0D+8z+LdyAxk6/7+cibOgw3MXqPTXh2VjzDBUy
KdB/OekbxAmciYWHJdpzbaDgf5fDFnmEBEpG4OCKFlcu3DN62fequPrlNlqeKps5P/jj8mrN+zV8
c+jUkLj+8a2cbIpd4KjP04qKEs6Dl7l3fOGmRuCiwBpBUwLIaW2lfKik4jBiJLdq4Wo9Hv+P4icB
+lvTZnj1TYEo+V2kYnLJJT9fGv8xbKvzfBjzcHJ98QqJCeQY7FqURhz1eAKbVS9rZ8Uq3gdB31OK
4iZRTydfv4xhqxUCDsvfdhx/MswvR/laZLsEouUw+pQV4LvdRIo3ORvfZ3Syk81ku6NdyMmbKLLp
LNHvChxdTU3Iml4PkaMakg8qNXRvf6ua2mAu36DqlC2pfIpq12H7ULrnqSUPWZpaRxX9TlkvbKWo
8Hto9D6xklLpMDgmuyoZZ5+tuea6eBlzCw6Qd1M6eQcpEyekY/5k8g2ioNeRG7QNNBdLsriNTl2F
f0FQUpMmb4zsKUYNx6Rkv5iikg7dbUHMTYCqygrIj93a7sd9aXx+v54YIC+MTeK0mERRDH24+HtG
bAOc6OomFlfRMa7FD0JlCtMTZztybX8YXX1DuqA1DMjNok+wy2zzrof0wd/Lzw5ejfdrUzPxHptV
w2rOeVY2nLhXpdM/CAPRVvT6sHDZjZ0pmVx/7CLvWqjsg8dom2uHNJbqZcelXf+aw4X0/sNHaFRX
slgJe4cxuG5LZ6vQYMAU6VeY/35kurGJ1bQvftnwoffv+K5IzCgVMDHi9ph6wvdrXsTKnPMZuEf3
LtJCYWlwQehxZRmHNkTSPvTLwL2fw6BTYXu+hsnZV/ahp7OcmpfEDY0wDIsY/wEu8ZBO0jKMpES1
ahUCuT0gA0MF5dpFjfgW/Bx7lMpO9s90SkWmC9cWVKmYVaDZWsqqZCQKspIw96WnJU+i/RcpsNXu
fYZ00xEyfHtTigZtnqfA0Xr+PL8I04iEmBQckYIPlmHksv/25LDMUUKJKXSwwP5JMzSp1uYQCzVi
L7ctaQ1Al5eJQjyodVrPkQQkkRfUgVrYZOdr+9ar3kExqQvPGSpNoGOKZ+369d1bnGJmYdJDxOFi
Nk7V//YW0jk0RUO3wGeS/FiQuSqCL8Ny4FWtnl6R2AwBMLrrRpmrSAom876b0Ue8RfTf6Tqbg/Mc
pDOzkYA2IqcqX6xPakfbH3YtjlTv6daanDarNeJk68AyRGgH8skzWT9YLaVEk4DFxlYRPf5QH+zB
myEapM10jZy3RK4BHhSanF4uuYsu5HFE6a4ig5hls0nCC2jGT6hee/kPEWMdSu8KWfD6X8wkjtwf
UUs9Z2xVVhjVRTnbYPYqbO4UWORKJb994BS0j+LfthNfTD5tT9SOJlsSL+mx2w5XJmCXKJulGBdz
27xzfk0zpnCPYwhqTH5Ie7R8RAF/26q7JNvl1PgqfzCt5W1xS+8sI3H1xZya4saF49Io2RV2iIHp
uaYodvrXefHSHbZc9s3rFhRJ+bcTidJTV/xjhRFQr0hgM9ywDP+BPtt4T6yEQUUR+toxumgvgCEP
NzsijHAIwQsQkQabowwY5udVenECadEzEnN1zo6+nONYY+/AbEUZARCZtxG9EeU8CBz5008LhoXd
qJhGM3fpKBwd4Hbvtd4U0+IC5R+Y2Ea8+FRT+bp5ju+v70KclL2S41f4gLB5C6LcBBTK7EgWXbY9
702m68br5L8udGMESdLFBBdr7ABCRHcpUloXS6GcBy6CenXkeDneRVGKWtgoOYtl+vr+uMTn1lkT
jS3PMmvyd15B1/HKDS+VKVnu6lleUrIGzi0bCzhJUaXgBtLp3IYgwqD+thYJJq73+f0ZNBJ7IRLX
j2MD8hNbkW8zHP3PpCzWBQMyRRhnfXXe2/C9Xu2xuyBzVtHvTjqByc11B6inYcZrtyoy41uPusLl
Yed+rst7I3zbOJ06qrSKkouHDHqkzmcWGjW/ihKRAUokowIL5TrbmAjMJ18ZHLy7B0CtED3PEYap
fV5bvVnsCJVfA2Gzxc1qWaOG62bOH6KaaAr+4b2ZqdQwiBIEyP7SADDKHBq9ImB7U64yhkIqGKUs
3UGWI7OuCWTSuOuU2o+llIP3xkRKV6Gp5jJe9n+mS0kM1xhfNL/eBe+fgx7IdlACO7Xl15MhBRwK
QCxiLxXZOtPDGkYAHUxq71HkEuuiQt9k1OHR5ClxrOvISFzSV52+A5nRYuAWuOBdB/9ucLQfr0Re
W/qA+YECCkcujAVE2BKwLQByCW7Jcar0Rfw1FpY1IOMQjqcCTn0OmSVIrl2kl7BtmbziSA/BKtYP
bNlSWOglLh4il+fHLqbkaGNNsNKuXDHi+6HfRYUQNmUgqRNm5DD4z7sB0RoyYrW3X2wQGqW/et/K
Hpvif+dK0KjXwOj6g08ffUDbTXC8ZtPbBe155z2ty8vkD/W+pDdPPI4u/KiPL6u0DBdCjJ7dKUJB
/GAZUcNQDwsvalx23QF6n7i88D1NNDAYuthwQidwyRrvaIGjpulDBpb8U3nfviUrV/fqUojQ1rOf
5apvCBo0qkNrUp5nOQMr6qPtnOc1Sw3YFJk4gR/mVbSz1g0g8ZrmXXNKznuqovCk1yjNQGPi9pwh
K56fFSZ5wjbixy4x0pBPTZsFJyyIHuJZBcvslseCkanHX8Y/Dx99y93rsczkdQU7yJESDKxmVrLS
XSFd5b08QFe/7Jp2hJxm59NSA7ffnjEJLQuEjIjA0JO1IM6tf08e+lp28B9lO1Tf5J6gQFWjYdhx
1KM6qh6oMfKnXcL2oa7EwPqv3c0a2TeQ8ZjBPR9ByhHMviR8koCYv8q+xBeV0t19nRsRAlfTUHJu
v0ZkdCwTBTwlHmxVnxfjoGQhQu3Vn/FC2U9byAhlXqEQcKmX8EI+J/7iTHKSxESf8JaZyi4iff1m
mwNekU8pdJI8h89U/rPJfu/O/a9TgHwSg6v6xIZhcsBscvsgIsrnnF8vHu6pf2/m9qnErs8nyLrw
fZ1NVlZSPeMz9+QMlifwe7AMDkNtsm172EzXiwFa6lFwoEMfT+G98q91i+XF8XVNmaDf6WJ1zyn6
eAN0f6kUO+oZBWwR73QLm4IRvMumDE8QXf9ALT/nfiQ5PETlDpqA7DLxlzqNVpOnf1FkcmXkox3g
vWV3WuXrXi4FSmfVwr5RZqnOJID7Zl88II0b4k1x0J+yoz7CtammnxxaDhql38VTrGQVBs67xGkL
Vq0wbw3O7ggWvSZVXri7cFi109bVbApLaUSo42Vdq6IB9SFFoQx+OzDy7JVNMR9GZ0VtiYqEa3DE
l4AaMzH0BiG8h/+9lwfY5tALIEIf+6jnjBG3iJVrLxXJktxTUdxFvJ/LXFIu+ivsU7gUHxQZjIiE
HZ/Y1De645xUjGGhJk1iRFmogPJdH0qfxN/0/u54MlpJxiLSr15cUgvVKFC2YeiWWykA7mJxsWX/
Uh0RwIzuzZ1OGiyZRE9Bd+BFxkweAKgBvRszwMlHLfhUA9Bzse2a6sqaUI86mzyM/LUSMa5KU6Db
ntxYKH/3ngwmHi9+WHpifG21gaX2JPFAn9ovp9zy86TdirlAun2pWwKnFklodJoUaag6bwG6+q/7
XC3Z69ENxj+3VXEzF+zGEelsoJz7RJTHm+8nUGndYzW7oXK/4vivigsJFXj6EUMrLDMYChHXGhdX
adJUF00Oc7R+7ksPiy7CZbmVeQ0WN8NzOZXPKCiMROXDJAkmZH6dDdm1QF7ZLLlIqxWIo7IW6gRR
fhW/CgPpNW7M7DtwOG2BqLPm5d1gVqJeSZnhHHPIITtfQPO/1xE5AYtnQLv7J9XKA8yYk83p8S3k
Dpshh213hN7vssXCFKU3vjEpVhbgW4E4vCnkpGOX+Tz8pz40a6n3m7LmwWM0LTENHB/f2pvj7805
FN6Lp7SLk/+rsqDP2Zw2kasD5KlQyPRuILzSJ7BM7/ThHku/zEResZcQoIaza47a4f05Y7AANpC0
jWzXnT4qA10bfoQO7vREao71CPjMkhdtsAgNrxZMLLl5o7tbXLnVBsHSQLexH9mb6ZIRN7lOVg+Q
2s5L5cKs+LeIcpru8YrIPq29mxZsdae78o80UlDro5N2s236FEyzz5vc2ZbFdWZ+zAS4iAf9EutS
H5MgvuI+l1m7mVbipWe9mHNW4lAA5QSP3BXA4XGxcEPJIGy177wPb57eV+oPY7ZM5bvel9tnXYg1
JfMEq3WKhpSQTitQPqsvG38OEokXIqn46B2RIqIx5smkDNiEZMOIz+okYZ/XPA+h9vtp+rm7EChm
TnZT9BAd+NV3QMqVYMBFJKZ13QnBJNRx8MY+FHG2K8ybye9c97dwCWJwa2mUZON6EpP8dLW5gE2u
YkNT0BRkeDgFJ1ivtdAJ02/qugzXNnRPldFLPao7N2TtkyarJeZIrOwY4NUgXxJ/vF4SwEDn85lN
qiQVdAxjciEWkKpqKQsWPUH/F3/rijqJDtQfEOXuTQ3qU+cJoJbXqGdazFYh+tbXHg9rjO7dk7HL
AsB6qyzwtrN/vpjJjj4KXyRJS5ZBkTdHJXchl6OdySp12ATsKkE18A6uWT+iYuEkm4o6lScSyEYN
FakVIPZwVzmnYB0f+0888OAwfNynesrvvS5/XhUZaz8r1H2Ntmz59YVfLOsAAhwddvpT/bWD+MUT
dap2uBmIlhUPZZTr3Osfph4f/1YxR2zu4Hm6j2ZcrgX8FlB+eSRofXA6OLEkEf8jhwXbplpsVKgY
f8WUzXc7x/tLpTxyqYXPBODvlhEpKCMYJVGdHmf4Uy/tr7WgK2ZXNgZNTq9i1DRR1zm3uhYi6Dhz
wgDRxqLLc/2m+BVe/WdYM8cS5ogN/63dVrO5iptExmnBZSxZi8y9Xn4Q3pFFQMaHVQXrOBEBhnLy
MCsA1x88iaPuOpWbGKMkxrCnPZwxhSRy6UvSJa1Xi7VxhKqOmdrXsPNzj7cpVZPpaAlM9+8GV4rz
pHO7R+wPMUGx3zDlY8032Zoifnt76MxXWB7TcmRCrX42BYD90BTKnGizTo19Gr6qk/krVktDYiq1
E83b04dGXraMK5u2lbTyDkyT0UDqEGQ34z+tOY78bvD/LB7X2iTYjCXt+r+xsU4UMKXgHBZYg/bb
DjHssqeFXy9D71U/7foIJmxEoDUrLW6knZv+dh9BQ9UsGW2cG9+0bqUlXaVScYxyh4qGag/6jRlQ
EI7HyRvMgqYw6q/2vpklACFl3RD7/bfjfRBuDY3jLA+rPH2WpxmkmfzL5zShfq14Z0e62wJxDmhj
+QPRRnhrk+97/T/2w26Z4167tG8Opoo1nGRbHMp/orFjR33aTbiTrZ0RK3s+Htr7GXYHv681SpW4
tZmzUKUZB3tvovX9egfLG1v4s52zfLVCRflRvkUwEo+0k+sPu11jHo10nJJXQpcOobuR6ua+l/vE
mc8pXqnaixIVatIIaSPyzwyZb56VDZIND0+w6pub651vawBJGL0HCsAzIavIpxv+HsKF9ZNTzbDD
j3osXQFRRIugw2sr1ddvbx6Vo4gdZ1OXF4luEbQMFYbp8yrW+vIIuU9nYqre8ME1/s5f6sFAhkrm
ljjv0MbMd/CkL7hcBOkAOd1fxfUa+5TTKeK6Nt/c3U1gq23StcL4lInswKQo/rGGmlkpG7OmBzaI
/sGM9g5KlwMalUC2NhoonKOEm8qOEcV07SLq69Ol403NErHeTsOE0VLrVvnfqAVMM6XxDqb/UPZy
I/wmlp6gijxAaa+Gngv94V1T1lbmIneSn7m6qMIr6pCExygttloXRWT2keqt6AQ/0IqT38soRAP4
7uSvkM/fg+NBGRMZMVOeHjvCtlzMdf2PTRCmqTfUHSL7pq7TSpkoy2RHYrERSZSZTiWMX/M0pCt7
7bwwldkAcugP+NQ/WA9UIiddSC/cEpkfbNz4IOGl56UmMFNZF9rao6VsPiOHspN4cvZzvXuX7ViJ
SKAW3XnsszbtlqrC6kJuJp/21Tkx1MJ0r/XEPNhknLfyr6wk2yRVPTisQ8S2jGtKVcyX5fIyqxT+
IAiPbG9nzxWrF3ASDGWoGkIA/VWW4vyRFMujzku06uKhb4rfyJfqCl2On9tF7inq8UDvXBa+pNlb
6fsp1rEcSNv9Vop8U02AbJDywKDJP45+/6s5zZ/jDtP+EYi1MU1ZW8aNQEbhn2yrhL5zbclEkAgb
OVUWyXKhi34KcKsmF3qoIyqJkRHxY/oAHAYs4nWajNUegCoomoj8MRqliT1/2ioxaRrT9vdrYLuj
A2lz46FX2kqaTOzuMnaJlVNE6QtjrtuR+sY+ZIPvIjLub1+U84aeFToL5t2gitnfr4jGYChbUGzY
Fc4RrbZpR8DifZisB7WTCHb1EIlXkpWAfYYGBoLPpPHAYywe4aFaVJZJpx6P/iEZIWuccqdtJsYS
B6Bw+4pWxNYBFRcLWMJZpFzAZIqXJhJE36jQAtcbTsC3I8WnWciuw18+2B4w+iDdYBxTpyEyp0rq
8pYPZhLfDCvT2f+w1GdMzisuQbiI10ofJb+j4Lzy1sm6JD3Wk5P5rSd7i2+GsSOdJEr4CbY/AJdq
mzGTyJ43LrJyEVn6wu5ZzmCytTTMZKsbQUtqa+hTZvIIqpePy2dyH8ctBko2xK7UCgEVgWZaa6t/
4kwua5rcrwuHlWNG3TJmpkuZ6UFhUL2BzR5oB7a0HSIDgKYQ3kDtGU4bFMugQFY+qiOFhMfYTIMZ
wuf4l9mLcZ5qXwl4faxDPPyfwYHBcQcWH3lOzIjEyri11BTadrPOWjjZBT3900cDUkAviDhJ2UIV
8EYRJMeoLvYegIbtQ8UTkrgkWF5Qjt8xioXy9KeLksZf0qAIYfoPc84Ahn4SqS8QybDcXRQOCl4R
6G/GcwCES0sHrF/ZCFp85iHBWaZshBwRngI1b0aEcOUOfiGF6L3oEJSYY643QUTR0XxdeiBk3rJP
cH/wSYPDMIGo/cQKCoWpVnU+hQbZFJRA7xchQETlIlLQctU22K6Lv95fK4q1wx9sGZNRBCQPINs5
7TJBfhrHu/PUUycop1daOlLBStw8jipS9mlk00hAqdU25K5V/3GyDk63RVeBDkOkc2kW1NDG8hom
Bbxd/0UCTRdrocNoa2JjDaneEZeUTTPRSlZqIN6BfSiLTsH4f4vb+qrO8YTnwYk/LvQ4N4IOrPR8
h9WL7rhwMlM3zDqUANc32QDASyNR7rsxc/2gxZ+Vo840NID6cF1/NNAuzSe6nGj1s+jkUJQnpdTF
iXXSmh14Dck8tiB3bH56Ayshpnk3NT7pqxLHOr9j5+uR7ysfLOF+uo/aAspWN827AV/QHgHpQk5k
LZngmOrGHLIHpuDHH4HHZyCXfM4+vvuAKlLtc6rFdYxF+BhhAqlv3M7oh5SNH+FHb1V3aHVK6J6h
JnbWZCTlbJK3iVtPDYrarK3jzdRIEbYLftHa+uvGp4hhgbc7FO5tNV4QKdQuT7Yvdr7bxC/qyIWl
d7qxW8NkVJW2VWGxFgPyXjD7OQnMsEsM3FRXdFhklnOZjCdlNR//X3BE7OF/ffVdFpe7Vsunh5NY
dKqF9vjxldFqy0D+LuItvRB3J2S/A/+p47rl+adwNFGIH+B0cVJ+YOAHWxkEUCXP5mTH0vYuJKG2
tzMKb4f7UdY7AFc26CerrqGNGQnTtRA+ZO4S4Ww+Ny5aHt0cN1HFJ/J8zQtGn9AlD/sa9nYj+t46
bh93OkGRpeCuYewzaZTX/3orwfVhEO11KTM+wc8Qo4zWX1JnIuIjt5UzbuvIh83IiKA8VL9q95tx
Moof51W5aXcxmcD/I4W/3HUzlsAf1jmQh/TwRfRkMt6xRf6+o2NOiwi6Dadm/v3cdx4sODZfweOw
xjAMOa+0jfICcokXlYhKlqaQ3gEm8gpUQXzbRCRo+/JZBpGgE/emgzAoTGP9AdSWiT3oM/YsDB8v
opOVW4+xgdzRKQqHcwAdiiaxYufpKbV0ucS8EPDUH4ONZ/XuAZ6EmOPmrB0x8Mak+NurXiY1sU+x
YBqRyc3IUk86Y/t5gct5r78nuzb4C6gpyFjSyhrG1A+KXQz++uG0Z3jAdc+mlY6ArPzp43V8bWoC
NBAV48q7vgFQgKIjOToC+7vqkAcZZo3ZeXwt63ObHtgzF4KmTszIaWnddd96STTIk9H+9zlNb1a2
KRYgCGBGcndNiNmVINw6gkzlH9P5xIHn1FgrHxNmzfvwMDpwgPjRxdyyuGvbfdsx6CsS5jccdTKg
jdVX/+m1Dm/FaZP9ofmv1/uAzfRoRqXAdYkFbAgHVrE7BMHs2uGBMSd+ZEkVmJryP8Su0bROTItF
pPg2SPhKSdqxN4B9nu+TI2HTL2sfgrrx51r7QxqbWp11ZP4P0RefjZJzlszDbYN8PL5tUYosmQz0
+xABEjRCyVajdLHaX7rXFKCYPKYitmuCyAOkQ5/ZEQ14o/jK5S6lBkRHoJ/Y/DUYY7xhcQ1+jDSS
fIsLEC0LSwDHwc1dotyduk1iVSS0dNY7Krb0xRgBPqOz75RK/LOwY+FexlftbdotWUyjm+fj13c6
p0ksH1/9jERJKxUcICkKmegyLLHt68lbEiDIPvEuMv1dSPiTa8j/RPfllU/O/Lo+cSc4bp1EzftI
pe7gVleaMzD5SirTNvkxoyAGm5xRX54reaANrw==
`pragma protect end_protected
