/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1136)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHITK8yr3bQv3/nr4uCYkJzUIoyiyUMfZqEsJcwNS/dgRWJz6bRE1GKM1q
JJE6p17D/XPDMoNM2PI1cYxGQTqJ+JmK2XQWD0k8qpp2piNeMMAkdYNLuQD4fLZVGJCRNZO6Ef9Z
RDOpTbXu9LQ5dMezKC8hKXOvGa5I36P1EzXm2k9Gprr7NkoK3LV8aMb32qbwEDLH4sb8+GAAk4qK
rHe+38X+GxV5hV7akx+Bqw3SjO18Xscg/okXQC1fd4A9aE6fhOvSvG/3rCvxA1yMiKsaJjwDPnCC
KsXI+PSZQX93wPmOtyrnNEXImv1XNp+H14F/QBF5nUIowvd0Gyuw/vjm2GrYl7NBQy/mX2bKJRBV
ASklIKTwh2i0jbtbHms19kmyj0s64F4+E+4vfiVKEPC6DYDdtiMMv8MCfKYsyEyRySKkNsowJOVR
d/+ZDUGy4hweH4qNNKEl9S14JzgB1ft9stQGnyU0AQhudIDHTGi2P92wWiPoLgYXqYWyKFRLgu4k
GMLf6uEJ+wITFpvnZAhxG749jYV53sLXk/ynVqwL/pNt92oYh+lDqE5JNv5N6c2hBrKScLTL9num
9CIaXdZLhS3zxbgbOy2YK35kI8t5gUvs9eMTvEMyFobsf556DyGr4we3rZdeP4E2FayUWbdihzcH
ZMMJn1hRWj1yfi6qCI1/i4NNZJQp+AczK53tFFqMUoDo9QIYAgOTclvrq9Ex4Ym64R2VZGwZGkrM
hYiiRI8draZkF6SQUDR2a9F2mFCOGUn0CtEmzCUvtXJKaM3pVmJyru7twu0DQa8fmOI4xOrXIqQY
AGaoLD0+SsFZpqVDT2DrhQ/Cj2g9X0U1V6Sy/dHkWQLosg84gcD01iVkCpw1aaFFaWYXUEpt8wan
sv0MvQbgYUru626vphrFDGAOgp9BfKdzCyoYq/SQQyIRkhtESwXIMGhy06iEOGq5nhfHKCfclwXH
+zGhbHIdssNfv/Y9VU12CmQqtedD2mZgdVgG1v0N9OooamfyyR+qStKZnVdFWhDywVZMrT9SkzkM
81Lzp/1K5Ys3rNOeCGl4uD3ignylIfODjqAKBdUwTrp7QzwaCq5rWVFXzhqsNpEukskaw4OfR1v7
P8RgEx030j0lHqY5LFMyFwVr8DIUVUbQvZrrV+1UHbTxcrTYOgeIe7LV1fUUVPyZzkt9Ydtrylqn
5o5BZI7WtW+yOkVVGZ80vPajyKILW5v+PNobRRUHqNMudcalQ+DPeiGryZUqLr8xa9/rPOR7y3nz
U6Qziq1ltj50mCu6QbMk4lM/YmZ8pSqn8dmharXMw8p1eNhLSRZd+qSxJTw9ZaMdNhdazDsZIGHJ
JrDNT9Fgv2th/lpZ7sL9B+2A/u4vN2cmwfWvvplW4WCE0NAGFwynCxfLqwEb5B6LgBcyn9azw3aO
RgH7qjuosS6Mz6MX+CqYSZkMZYNLQyJLl0VV41A4DIyXSiUYHZ8cLysLTsaJgQBGbIbi75c=
`pragma protect end_protected

// 
