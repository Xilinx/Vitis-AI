`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0INbis6m4LNo5fuoc/7VtaFb6U
0+5fXdMnwe75smPOBFJPEC7G1jJjzTejAYkTl7IUTkgZKL+qPo9QsJV8bWnGHQsxi3gvlQOIaFQc
GeHAIu5kCH4qdG/Rd7Opht+51SV6MCUG+Jzw6T7NCWSvcK1kUSxl+7AIlS+WIYISlJ+EKHtGVS9i
EwJnDml+BfWpTB9xPafHkbwEu3i47lW0rm65AtBA0FQc0g9XjSdqF0izkDx71iLWtwdJ/ACCBQzi
xKCAfO8AybV1FHy18fZZX6JGOYY4nPjIsMWIAxcExkw33RJN92UK0sFJvBRtmb8CnVVgJsTPzqJu
OmUNGCqWgOS4Z4jTkBDRru/Odanrcw8zYExPvUs4l6tYrjts8KjyDGFqQkGbBAtCI83ecpYe/O28
pLkoUxk2NZtwVzGVrVurJFTA4cKDu4dFSHfmxDj/uGVX4WS5jWMY7jieXojAUNZIF1n1Tb/zDwDj
MBDHWdzD3QkeGdDo9C//5HfFk+Lp6mJB1phTs/aDmluMCJk5PAUhKeH8H4eZZ2ehNXZlWe5KWY0/
+S+9zxpYttxs+KwfBiUU5HoO2TMbvFCMRXdePQdiXz/GosD5P/Say5/dtCrGfqBo6QrftVDlFRCr
xt1fnZmy2j0U8RfIF3XP46Er81AgMbNqyiKxKlL1Usgg2GunliKYkQXLJLLHSii+Kohvl1Fnp/2c
C/CS1oQc0cLRu5RdIPQVNMDzjgCNchlv8TvHSNfSIzj6mk069o0kN+VRr0afZULs33TQTQB5eLqV
uYrT9AP12TQ1kNl7nounShVBgskkqYw3yvtisp+Wo2cJj2a/nM8sVNfoOn2ZJUy7Fiaq39p0yUcR
Sqb20CutgoAm3r1FYW15lBVxfp64ivXJ8nICuRi+SSgQwIoCLRigUyz1mfU7dI77jkdb3eENeHpE
GY0+OAblb72w/OOgUm2ktWE4hDHCl24zq9yEvCHUFnLraSeNKilbIxB54Ybl2yYwtFXzgDY+Obt2
GKCvZ+Mk1hJqxvdUa1t4BaVCFFgWHaqsot7O1IW3TbYi5c1umRVT/Ia2tZm2QcKWehLGmFCbbCb3
zLHjb0K8j4y656qiYNAn6En5nYJtfUemqubFN6UdARoK+R932j+MSe6qWeoXrEg70gb+kyCT+yy8
kvnmRJaZB2zs/uaT6Ol40hHBIoBxnAItYqT5RVQTm+dMB6LS37Ju/sSOQE6A4yDKXdc9ixifE2+I
YGXdt51cOjm1VrhEuZ/mS3TwMpifeXE8YgJeVF5EBPxAmCkLL2ai2AFQ+2Y+c0k+E0jZKtnpVjrO
5Xp/cwejIEbYnOkLls7vWbqoOAAykD68FRV/0dKjBuHrdruzq/GHXOjlC4w3pvabNBixJycWnSk+
i7OS9lWQ0evRcgxC+zMKUb+4/dFRlvOxuKVlQxo7ohMtOvdpg930lcGtR4j3RQc97Mn9qE9RJW6D
qKmkKS6CrtSwh96sBXBkCAkX9ZuUW+yGl6qISzmRJesnxZvRAcxzu3OAIEmTUIwXL0kvZaGEcMSw
RetQx2tsq/iO5NsHUA4o4M0GQuxybYj6L0j7vVO4ckegqjhncmWcho2S3eZXokWoW3XYO8Iybaoc
VzmhhlrvwSqVWTkRZR+XAE+JUAGq49gkBjQD3yNSRWm3WMjrss1N6vrODQbPycaLjlId5wi2wGGG
IFc9UiGRjlQGg3Tn4E1jMGG69NBhCGvpYx8TV/vctGZtQZXRDYoCAxasVpr1fQXCMVpjr2gwBfWB
P9u/XyWJKQyKwn6xUmg6hHXNm+QKIA8+lG+pLLFCs/usJhQYbCOpI0WbpuoWnSY2m8+uz/SAozTZ
8KIlcXY9jbztrBlH1aqdrFXLr1hU9YgMhz91NcaDPXZ1FTcj2trtqqnx8gR+pODxC+bVI8+oEdoS
d23Wd3w4kAEWjjI7I9dND5GBO8+53hlycru/kpxnsCztIvt9zkPiIN77D46+UoExLww0fUpLOt95
hiVKEBFSjZacZynYo7lEM4BIxVbnCZ5pubapP526PoVJEfNAPDV5pq3mKrGaTsekx1ufZr70Pzz3
7HbL6cJ6hG3uh1yI/efFFBwwgSpF5fS+FKHSMSSvkOdayHpGNZ4TCy6T0AVyIiSPoGqeBItKIkmz
Gvr22IAfvJ07PYAU4s7HG0AIwyIkN5T5wrn7bxTtNkQEJY0kozfD6NoFKoRVVJ1bNFau/yS99Int
n8vf7Rp+qqfqV9DlOK0RQmZnYDkRsodgZsFIbFbeFNC1S8z3RtlLgF1Cxe2Y+CDbTJu6rGZ+nsYl
Yiu8ks+c49j7h9gIWiQh26xZUR/7Rdg73uQL3kIbs8cHq+F3iHGofxObanreAcbDDanGFOGRZSbG
TpkuRYOtDqnNwhETrjOaWHVxcK5TTLbp0vnbWNJvOdAo8VWKd9sIfedj/LNrFIVS7VaWnZW9gq0F
3dermL7ty3QG2Ad8FYSzdFx4h3rkui/ahZf4T+23IAA0+wYznZ5aLyUJ7Zh9r52XImO6+OX+V4r3
FtmxTMoXZXsgV+O6Nw4hZK/4tKhOCJzQQHHeUg8PpymIAx4k1X8KAeQ6kotClQrgc7CvJNbLJEfD
WELHZX8bXL2WoVJxWWSmgfHpW+XFBhaFBRynz6vXOB3TwLKKEWNbEOASp9Kx+KmKFscvdYGxM/N6
rFPbd+Dit5QjTxnxAFHETCNl9f7XTKfl1MV6VqAwOpO1PMxIMIEOv/L8Lctw6SGXBuv1HiGRlP+p
NDOyWi5sQkrIcGC+qVvUKpC+zqszn/kuPymIVuoAqtp2b3omUHUl1XnqhPaIvXkQiVh28IImmHCn
IDc9ShBKZ9noNSexXpX6xCQfZ3SYSo2qK3j+Eu4AHQ+dpEI3M9jocyEq+H4FNDC/SsQidBqHQqEb
dX8ysr97XFb/O3gU199NQ0eZv1S1IQQrQMxiOomni2ZLh2Ab5InfLQ+/w0trK7xVCWqG+Shl7c3J
wJvDHDAH+Gyd03xFli5ehNX6VtmSXDq5/bJpa58q61AD3vH3SnqHs/TMFSmsiZrHgkIQNklg/xKw
AITtML7eE9wdDpb+2o7Hy6SG90addHm5DsQDF9qqlMdTvXMUNx/am7PFn4DJ0epJnDca449M3Xji
YRQjwT+zev9oGSK8Y6u7K2LfFepLehApnXj7aIeVhqyAz7vq4Eh0UkzcL+nHeFdCoH2WYPPh/Nvv
HeG5fI2icKqc7FqR82ReISBzVcTC6qeXyX46b9B42DqPlx2uYaDynVGO5b1KCcHUsXDFGSwxibY+
W5F2zObbIKI0/mqHgbT2+Jk8Dc/b8O3zWc0daL3BB5a0Ym+/NhNs98XgCrUjgqHypJq3wLsY4o5+
++y1fPIP/NEvrGxXlrqzWyVVUDDQuIKP67ZP9bkGxb5z9Ep/hKcd6kTlbOEfhk5krQX+MWpalGqC
RYOWYzs06fEXtpOW0RkfcPYoEGM0dlEhSZUnLtT4g65DahtiTQAegbYxFQZT30aIn8YKDzNoT7P3
+XwZnPP2CYe8DJFi3E1Zv/0MX0TmKIdJdZzZTH85LOGFkC2hs2Nv56Hm/VSKZ8sv6TP/k44FupC5
ws6YtGmTgsfqnig7MJdYEDhdEb54cgwci/JVAQfzRPXaY3AjKNzcrypNrX20xGNX4r4rUCzR27gh
7swKZ6UdOO7Ekm8gWHDIFXU8ebU81ijb6b1roscX8Kn/OHmOBM+F2h1bC7j93BtCcViSUeMGnrEK
uDZ2ufCm3nDnqzI1W7qMSVjSMRi5xzB5dPUS2IKmMl0JruIzlI4cu4YbqPo0GmWNmrkUM+nhOcPr
IIu7av/YKjlesdKdCCGCf8clxoaYQhSkWiaRyJV25Z5gVcWacdFTtgXGboLyioXf0bYdOeqBZQ8W
HqK26UftW6hCeZfzoCwnbsD2kVY3yCCgGG0z1sVbqF+8mmmBHIv+9eNo1VqmrTrUYOSaH0D0q1Y8
TO+cxaiBbiFYVU1PRsSuR0d8nw8QZfqKuJyQMAN9rNJfgVuBdm3oi6vpTk3YwsRgUDPaBaF4/D7+
psJPKg/naf19qgOWtQGKkLXoezdBzFfxAv+DL1SS1UJXQQsSUwAreHeXnoP5aHG+BEpzRF3Ow3F6
sngEOmxnguiPwD9W49CIPV0Z2VWms77T8UjK8bRPmBUkIp8Q78EHT+uz5xdi9Jwya10n/cxqw6vG
BSmJwRtYZFkP0Dss0BvGT1EJv+YdTKoTbS9a0G98kEt2E35Zbt9enU3Ccj2V1OO+vGJRN0DewcU1
VPeEA2H0SlTQ3brWRZgSrlO6YeV1GIBP7EDJExw56CKyjsmaqlhUWage/YO+/of1BB1xjceyhULr
zTsv7Tt3GT89ZCsmBs4SrvsD+kLo3H7hFkz7os4SbPGZI6SZvQ3/oP+o5GHBq55r5hrSt2+hr0tW
3swshJ/qo08ut3O3liSYRIerF9PmDdpqHvP61j2C8rsiOHU7d8BU8mdVHMA0Z6+7thXXYkPB1Zba
sFtq78bZ0kNaimEzkS60dH5elLDQlspnVTg2jLrMN1zhPw9BUw7xNkYKyMYdgg2/sIwNDR0K7Fhy
MpPBE3MSaf7nBkcU1wMDaBJS1jZETFZQ+GE1AY7SWKBlurKtN8kGL8Api3JojPq+Q2GCg5MeDTKr
932wdfc8FNarH7xmlMwxEgIwwOBx+L9FKFHii1F32eUZrey93uhyCuASUgjQmntfCI/TLNnbKEPt
DExTT+Eg8S2QE22w4jPVu2rKzFD0+hi0xlVzEwOD7aL7sV3v/hQ/NSLUOE4omzzF6vGym+jjc/FW
OJzgW3QV/X5DDgH1Kt4WXEwTd7S6s0pPT7akAYm36iJi4CG+mw5t7faRzWYk0g0jkZMaU7LuyI30
tXm16W6P7OAC1/kovBiC1RGIoTnS9gdMQgG4atwVgHH0I5I5CLA0zrrFWEDPwam3DICI14OgFCoX
Wx/7zb7J5H2hRaEE3o+oujk5QLONsx7bHeVEhw5u3c18MmLAC+D6Vs9vFBPVyIDoWspjGi8/mbvr
9jGdqx3NcVV/NOWeM8mPa66zal7/52tD8T1vvAJLhrHwiw7MmEwKM+3oNkEDN2Byq1WvC+kzlUqq
DywB3GV8ckQanwiMAfBMNYJqTeyb8gSstKFlLaisJ6+sBOQgjnlOwFhihR605BgypHGk9QZem9Ek
m2k6ca7eegzIgGRNEeQO2+9U61tgUkFYOkGkglbZKxDrNbl9v6wRcSMnPuPudI8ZMDlY/KDPOWjO
dl8OBNtun4BBHRjIHQMgrSHzC5cMhtrhh+Cl3JrLeFxb+t9Be9c4wtABjWYhlSN8gG34X/sxi7F+
oKWEXVw2JZCbpXR4WYSlEAFdauCneaR8/yS58VDPuwaBXGvr1WPu8yfvUlxzyzcZZdTu28fXSHAw
VQ2MzxcSRvI8TKzOGrqnBPyhDoF1LbJxNsU+fAwYevplZcumuSGGUGHjN2XbpDYiyx1PpkSHhmfs
WBDqmQ43ly5DncQ42kx5ZOLqLxN0gxyBwHUD8ujmoQMkMu12xFDu9oRDSWeIS87lW1veffVfYUci
//9zA5+JctM1qn3bGl2Uxhc1maVF9FT174mmIjK7IqFGJ4NizDoQwI11uc/GEDB8frlgRir9saEG
MtrWeg3ttpe1Qz/90YDgDfvouBWsC+SDpg+wcUTY46TWMyHfaID3rP0UGTCc2KaOXo6lUes1U+nm
s3p4cALd5i9nBX5LwanpyNVrWmkmHsD0rTjZ6+2JDRJtUi2R8Rne7anBvWSGNrPIyWMcxGxyx2sd
ihIl2V2FRKyGFINjIu2aCP/Kn+z2Q+6Si0DbsAhMzhee3g74ZmzaSLQfH+Fzv4Vwf3affZjcrWiu
Mn23dX6XyxMr3ZZr+bTN32vYO04z+uL/6u59/i6JjkSLqWUNKbl7BYxrWlcD2VxIuUqP2bdYTGCM
b8A94n/Pz6UzcjgonuhT4wTE/ymChek8lPHp2Xw9DY67dLJYpApYBrk13dKARR72VTXRDhesiFGs
HowgXU4ukTwnTj4OUyGMjgkgHnNI/wCJjFZ1z5Ei7O8o2b8F8QGTrN/U2WiEF6uFJVOtixDKR57S
FVKKpeKX+bNY48ind3ZBzhl68VLNAl/F6+VsJcR7RqioXA2PVOuItqnxXf+3RnR7I2kVUCKcI4du
tefr2s9ShsoRf+TE2izl4vMVQ30gbnOPznQzY97wXCiPnEIfQJKkVADScy5Nl9W5TOEJTqDT25Ok
2P9edi/HRwmr4NB+nSnghwj7Ck3fsPYAqM55l/2yv4Q1ZRAj2zaleT64n2ScYzwjdfnEY6wVbSLa
00CT/9CdRl+q2a+Dx44KVzFkfqmZpWfry1dKdxEqZJ4zPs9dBaa9yTC/7cGFWgx1OJhUqZQHdD10
BhQgiifQs+sxxcmPznGQmQns+LpZaKvW6Lu+KgH/5IZbZPwq2gJXdkz8WwKBnaXFFt/V90EiiXid
z7ZMOrNeASPESwWe6mFYUJV7XjEbPl2z2rWFtBjOeDRD6flIC9HD7KUoNFQu/DPAxKjoMGLPzToP
Rx/C5l3B71N5BpjkgPC4dmk9k94rcgHSN1Zz4e8UbaNSZV08g0TIKy8GP5DyA/4uZJ5B/UZDFPiU
BXJYL7v+EbEFYNyX3KplNM+rzgApwMHC/W+iprvpeWR9Y7quxhwyjVRDXOHcp4CTUt3u0/yFtU+T
71t/SKq7Yt4ECqWZn6lFlmnE8go9y/Zg37VBLhvdynIBZZZZpchSH6/vsIlgqh1/G0EO4wh9/Q1L
7SHqURDKpSKSxYp6xBZIiE/gxIZYgWiJnxaN0Ox6ig628e8YanrXUM01kDM4hZ5oVvNuOYkUiEob
5RfWxavatqgHGY1BlqXU4ODSdsppvnedUp4qiuXWlwky7QpYsMNIps9rBm5/pCUeQlo2EjwNb52o
NPOZ2+P1D0LaCnKtu8syZvbBsOoK7OqCWb/Va7xMoKyzWOsTzuO5X8wLIVm8BeSUzCGpov3XaiQt
qKowP2GqUaZxgCinlSVdKzijuLCdSqoH+jCYh3mYrlC2/9U5BscM51htdmpyTWhO1RrJcRSUh2oy
ESPNqHnz3znlBEQD8x30AMqm9gEgNRMTEwAnQ9FA+yFzIwR+DaHwwH6G7bdK0wEblFFf7eS12397
QoNRUFdDTyVuxtVVXCi78C8/PFydqjMgpReg7uazB6urEeGbTHnWlay6VyE2RlX8+9jcbVJRid1z
D5m7sNtGPGGK3CRxRSQmAQaFRbha1e7qTRzKYifDb76LyWA9Rc7S9AtPSi0PqaZc2vyeR+sP3k6R
yyhM/JQwyQDU+u4Qk2hN/+FkuL3z8Ml28TQr4LqHy+FQI6KBAE8VI92bJGOLc/WZ0F8s0IEe8VpP
beeFeWs2BsGfaWGavjlScNGYPmh62HONkm+cDAP144OzaWsJO/TEQGzLrRCT3PO87pZZao2Ql9iZ
9t3qY5owbexoy75U5EelhkJjneBG+ENnuHKtxBM+KPYYseViUJwsQIU9fjMK/Vs7OrWWesqGDfed
lNgysoNjX8wD8VNc85AHnZYhY60+AB1Sodv9SQe3/ndP0ioNRogWewJyYb79sYf55xjKnasPo7YA
ErGdptylB943Ja/7fk8bSgo+Y1MC62N7UeLMyibz4KA4YuSIYG7MNPOAuoTPrmoXlO09I4ndDZ+8
JnhnXq8shdNfx9o+ZXAqNZB2+J/IdymINgUWfCCLxV0PwVQo9SKei3FVLEXt1gTO6QxCaAEqyFzR
/U3j9QCmwbE4nki3MVlt6iNEW5lELK1hnEBSJ+a3Ro3cjdg0yupnQIK3MFP7axwHDPQR5bGZBdwL
b0DM6mjEgcY/D7byISh5X3MfEr9m06A6FhYxIMmN0utWGqQiBZs7SbQaH5rfG/nXq4zfBkqrft9m
2/vgf/86huqF+Hg3AxW+zPWw9DdnETpgHOf1v/8KHEP/nTO116TLg2BdhSQbMZ9Z8EwAfQp/CSmn
Bi9Ck5pClQZKfhnHXBbF6JWknDaYa0SGrdXNwVWCxr+iVjYmDT1eAbbFIE2p72BtNkFNv0vPTmgF
pHc8TF5z1/AIW/R8mh9RbrSUxZiPx+3JWaLapviDQO/+6Swf10iFkizHPncJiLMikldLihE2egqp
qlqK15gD44NNK40A7EM3e2WqeyoYjDvJvm3kPEnwiddJFUIOMrOeTvKf3hhwq3Unm1G8AtaDTQXk
r5WgY/D/CLxgMiVw4qaG6BmYkcI9EqjoXkxXWWz8PLCJrN6PS+sz2aNAamvk8rjfcpLIFmN1yb7o
/JUJHi61Xmm6mWjNSfFOO5NDdGv51rhGFmuOnczjK/hIrzkYKJOHtWyhn6jP04fJqSgbHkCZakFk
CJPHhWhIVlkmDtMfAkerAb0JoJC3GgXqzUV/pNG+2OL9gV+wYiVox0dY+kr74/Jm2PXvHIvbDS2K
jPxXGhvDOtRuOfFNXLkrDCuGX5VqNSdKHdfctelu7B4R1Doq6CcEwWuQML8TjB1g/0/Dtt51hyQI
1cSQ1SU3p8Ql4v0iTkeMzla32q6uYNGoUlNd/vXA8KujIE+cmPiT8YjrFPQp8+CJSBGPY7qoJRHw
fOQT6ArfoIYN6Y5SkpBl/1+nlbT84do/7gt6oEkJICIHWcFUDYI7uKQWcL9JndkpxiQbnCj1bxr5
X8RUTZpXbS0w1neEYvFfeOoh38PEhlFjRqj9zioPPOQR0UaxyCtvRi/4mHvw4OXB31Bv4VXJ+0I0
tyvymfmJIv/V74fqD87Za7+fZ0XRtTqDCpmrWxqtWyAh5Sb0EFFkOoyz1ndsblKyn4K2Lnrx29rC
dmobDBiXjqRx3iQ6g0gNRxDAvX9nsrXvr0cYoHrX6BJqrwvaIXMuxlkASkUHU29eEW3bEnqfcxxH
oEDz/UyjLQswrik0GtRlUnfrpltiIYY0g9oXlid2PN5/ol5fcABawpMB5PagwnbCPOqkbXAu01HX
rLTYcTftqx8kEyOrL7R74fFmf73aY9W5PMCgZWEi23lIla43ReFwt5tAUIe7qExGzR1nZuQj2jPD
/hp2zTzeqx4oxU3fX38P8oEsQgWSXt/X2PSN/AhbIN+lQvx7RYWLsEXV98ZeFXeF8r06jFthTrr4
o+8RU1VfKEUoRip74isAFKY78ndOSnNguK0ro9O0z9fsCgc00e2JTw1nzLyz5PbGWqKbpDvggz+5
+31mgaHOrZ4UZyGiru2c7+uZdttYFfF6dHP/TdW9uG4hrhN8q+7eeeAd05q7D0Kdh+Wz1oL50hp1
P6DhMh93A7ryg48k/Qh9uOpIMyG2awgyj5qFQ/kCjqe8/eWuPnKt7f4ryUVfh50dLaOtLJTNJZ6H
u1GFXusP5eSmdxGHAzQvd5eyB7CWCnPPP7u8qQDljr7X4capYaFpyhF51nJxgBrSEk+imOEslwYY
0knlet386VfPSuTJ/8iiUK/vlEJhFeLLnvTdDIANll2qInLoRSPPu5LFzgPfFa2wC4rXDioWU0Lk
+zlgoLfHDA+9TDoXymSzCJyR0j/drHbgt9+KUB1mNKBOzdK2NsaYJyfq1+tE+XKb2Vevn7agAtu7
iD/H9ZmaJpxx1qU4G11BNNQDW4GCpwF+reRfO69uWOxLrDoZdjne6gqR1S9xSptF/ZSDy4FxbEOm
HAlKeTBeJhFG0o65vVpO8bu6oPXkK8TXu7kmilt7tNGeeqzuk5inOvG9KRkSc52nCFybT2q6wKIy
RmrBSfjP2Cp5g70pzYqiH7KwfuabJnPB4EBWVPE5B7S7ZOf9vLOHIpYQIeWanqUz0K/Rgn4SEkVl
YfztbTDr+EdzYZa3WvMOH3i12RDsBJJS6F4IK7Y4MSXFc8u5AkUG56p+OMb/JmoypXJNf4ld3Csg
Lke9nJiAMkTSviB/RtQLws8+izSGch/7YmDL+3y/fQ4Pa2XXUMojFqK0cNRXhinuM6u+qdsT6AAS
oqYtyqDUq8dfC0yOPICfFtt4NC1YFSkViBsJ+FtwktoaJbeGHv0BkV5CjIoS+DnpbOqKZfb7kb5Y
Ks0VyEFF9TgrusrD9UUxKi9GeWQhzUx3aKcOLU6jazSr8ZOHw4eJIkiiyGyUaFjQiz8LvKhu3u7c
Sw0vpyMFFwT9tAKFTqeMJ30+8Awxo5hmBVGmRYDoiseBnUHGQ0UCkmpxeX+Z8DzVO+QR/Kh7olRY
x/Bgcq6+i4+q7hf7I/zSfLfYpO7hKZEK7Y3TBBODEzCCLIXFuNRRffTtq14/JP2cqOnfV+W+DeB1
dYXmSoVCpgZGhN7H7pGfk73v9tobGennmSyC+YPzHBWNbBYvIroS+5KqGypIzuzTFKq31uaKbc2q
nVt+0md5xJTqGRjDJtEV3fN/TY3+hpEkkIlm+xlSCXhu/VxL0hxfys685Xs6I/WwDSIBRDXITmAC
SzluTCtKK/ak21YQvgwbbsWmEyPsa8Qqyt0Y7WbCYFPwa05jjzE4fwJcrML8lJRgI0JRNwaZBP4U
ztd5qvRIdHrNASzBlAAwmkql/a34sVDEXD4iN5Bu2gGf88E2lljJCe0lnempPdIOHviO+feZ7dGC
YHYo1kIpb1gmCORTY4mtA/qN28jbOHYTpwuh87E8qRL6FCBEtqayjZUGfs4gR2limLb/bJ+Yz06P
n30w+CTePdZoq3tzxyhLj1ds0e0lNETr3hPLP05bbPtdkwf5b/7hikawALyk6kr3ul0ZR9/fKRLU
Bb7eBEgJ8gNSXLYWjdB75ZEYdiwPhcIX1ZnEOvk3vf5BaaNG84m63z4R/w/6chBU7LNn74aguH8a
5tf8jXFwcHA/LYppeqiGT/thJ/wYVeXWoKV556b4FZjF9rr9CCnHk35kSHYjDZEXjCNzJ3xO0LVX
tH3ZiyNjrLbypvTM253v72+t0dQ6CaNOjCjeYwB3Cv55prhVjrT1PEcnQKpeybi5mYTFUbJvsCYG
lwtDTI4MtALeMFAKLxvXPRnw0mX1JT7BrEid4YTqr41qG8+rplgtsEf11EXa5XhDIdlTMZi6yReN
2xS37z4FHmVp2Dkv4Aw3xHMVI0yS2YyRbMr+6fTH2eM1g31RoUf434dOFzqco2lrtcAHfXiIF406
J3FDyq1zsM8H6gkVhuq6TAaNf2d3XsySogD5nDq5i6eYNDFh69dpnOr+l6D+9vW4KQ2r2+4eef0f
vaeTWZwmFOhHca4n0j4pyZ1FdgbErO+zaH2cRKL9EFLXpGVt3kmysK+CgPbJL1YUY9Q1FEb9CJUP
I3v4pXPj83sLHoMkOaG8K27S+Kn0oV07umMPSOONvBCvpEkk2ZehHC9y6J6m3RryyjD57Kiut/WP
Tn7VGR2QHNUYCmRdxIRvQ40shQ8XxHFF8O5T9tZ1rTK6RINrgLRHY0e+piM5aejgAIxrR6Z+W9Qv
eyTVxzFo7wDowO1uJS2iDUXqyjc8JsYQVriRkbJpdyZfzYZxAirGikN8pskkcuoTC2B8XP4UQ7ks
FlwZM9cAnthL3Iy/kLnYVwQ5QTQtyNwezrPExDNcNmt94Ga5F22qZxadZoVmLyBZzTJz2Ec7KiSo
wV797umLUt+BMM5auSnnRGA7AdpFVLua97qu8BOZ/0aba66sGN7gokm0qkr6XA0h3Gy2Bjds4wha
7/rcV8yg/533o0mDZZSgcsfhZpTJKBnpQaFCS6JkQrLQILC2W4cGnp3QSY1RY1dUX1j1OamxTZsY
5UypMyW6r/2+W/upMygJqfJWiYYlbMcLHYxJP52LaFaXtQAsgbfks73JL0LWQxH6+/uKrZ+pJKTv
3G4a7rGL6AgazWZEgK/LXsD0m3t830YtJcT8CkY0tAAn75a3W8maThK6JeM4Ej7E95aZq1QzQFkE
ih6PkulrRmLCD00JHEfq3RlRwh+iHCPH1ez5w2lVGDJguhdnkFhBnB/lPyZK+P161V6KrrvA6nCc
7jF/tUjDbTpIhqkdG2s266/NG7XbsH/v8tIlhFmIdEnnSxeBP83Lyst4geEm1ZYcTHb+na+S4SHL
FmGHbWocOma3nhiPNiCacnjFyqauVvSmqFNfmgghM8hnw/KAE9chY/PVBEqCWzi9QGzaLng+1EXl
taBRmQfBmEXfd/GH3Pi27ohB0BalddxwgFL3bVlSqoXxmkp1BdmWGhcR0pKuf/h3Y1tuNRmUegEx
9wEuG2vS9T4KNZIm+0f7DuXFvOh3uXC8v4JOcu9UC1MgtrULyc8zLMLrTPQ/WjnM2r0g3URdwXNU
r0EkjheHquB4OV4X58V6JbpfmAeHBE17U329LhxxZeR3c/593p56DlZErYAmpmpwW3+ad2xSCbWY
MJ70F5N4ousOXRMWNQnWD8H0RemOoBzFtdEjbjL2Z5r+FRr+8vtLevomYUo5CASj1KIBMtJrQRAI
yeKItxm80QihNDNnHnBLdxY5gZ2iI9QW1g2Vkh0U2YK73Yl2GCmlOdGqRLHP1eUHEf+3eD24v8Nt
P4ZrcEwWbgss4MRRLRT1XjEynEkRTZe8JsVnXdIFe2ORFqPlnk/jcbW2g5228SZPYV66gUxI3fNG
nnzcN6dQnbduGDL7q1ovDecMI95UeCcykb+zgtbo3rKosy6r++DXYIauJw1LZ04yJx20MM9+FTvd
saIpc0VmOEVzaz8qccCCk4hjtZcU0AILCPgsJNG8tNF6mJExHhkrHsTQmg9YomHeceXdvfD1x330
zeh3ptz5rK730irtbJMiSyqrXuTG7kK7CEQe1CKS+ARVJd63uipZWrPEYbRyZOLejSJ38kfsF+zF
s13AwmkHnW0MNJxCYDwFRrWXgAI1ggH+9t6hJoFzVu0MfHkcldUAwIf/4hHemeyn66pQ4AHUvQXQ
B2fBE8VJ82KddlNHLYvsUndGlAugnIi3LJy86JGxitwSiKB270wWmUDYlP2Y4TpH4Y5eMTcGyvju
1/KVjEexSN5hcmvgXNjkVUPrjnT523EufVuDHpt69F1JaYSQ+Ht5e+axb/tgNuhPjUG523BqchpK
k4Ba6tDPXRl3TwmZt41HAqYrTqO5N3HpZd58bjfVezbZ2M43t7vIl2Q80X/YSHxeS6KhiwLmEhhD
nc8gdBu97scQPdGBVkmxG2flAjZo2NVXwVzupQPeyHe2HFeXkyrdHXpa3VOP1Pfle9R8Pj4EM9dK
2PvR/deX+I0nlWYSSqcwlb9ClxXvUd9OGlb646439aEyMHqt7AnstOoFRXmS0VX8DYte20yzEYQh
Na4IFmNIoGlA0ET4/EEYpf80H+9y+RajnICcmHukXdWaUGqQ2VhWd7aCtciBDrN1zxGuTd6UHqQ2
D9zL1PqIvaihl6mpI8I6lG3SzlZ6CeU1Vyvvy7WB6WFx+g/xo3Z9WQs0C09yD+vFcRMaDWl5u+VT
2OIfCuSl+3YbiIg9D/NX9hE94CRDk0H1Ba35daA7iE5vWBXw/ORZdX8bcgOTdV/jEDwVSzsHG11p
KcrIm7RL6+Ih93I+pKaQ0sHJjaDsDAYuljYRHVzjvkO3/nSjJ3HR+lX9wa8xUFXwzgUUlpNvuYON
nZa8IzNAtSJ3B5ITfU0gUzH8Y70UebpTLaReujLYcnuNVfheVGZMaF+z+OL9qDGpjKgkMGLWWV5W
FdN+U6Qh+6Ga1Re3gehXy/NG9+QHJc2LfbUm4bY8df+wU1AD00Y6zDXnsBcQQL3zbkot+UZ35leO
aUW3n5BiBzuOEo+FC7BRJFhFXomkRocdo9MdLNLIzwAUX9Z+XdfEZK6j49twOshviaZ4TijaOLCQ
bs6bTDNjqskWPR27pfTmJncL7R+7ql2/TfTN/8BitUQEkPRcnitrqfUTDLYPrtdFeHHsoJd93xL6
CiYLZUb3OgndkZoh+wAnqZwgn7xOCXR+s7GLDU3Jj1QlfQB2cYOBDG6zqnsviu54DW7BIfbgSgG+
k2jfQMKZofLFMZuRz5H8WNOQh3DwEhQYjVm7Mj2Q1RIfNoqVBY4XQjxnxq0LH6cZ3ycoz9OnS2M1
WiOcys91G5zZIPicTNPI4zk25h0kuZyYEcWM9YmED4wAg8fa/jOJ1rQyv8hYSa9LQ8lgALhZPEpU
w8/Oj8FU5eB0Gwpe2ZX/Q7MQhYyizuyhMcUefZIE7EtjUOrHcz9ejIIOeS+tUuPKN9UUCB261iFr
fVsoT9S0miETsmX2r/9hZ5B2LNSD9ILUQa152jk8lO6fXwNbowGK/NWxda6SvtqlTzUpl3O6TOCR
9YrDyFPo/Ibx49dhMhnHe4UG77nVVjoSzHeoZ4cyihjoHHGQYanDAniUClKUf1pjOQSq0eUH0zS2
KaPzSGs5i14yje81fnP1/MdZQdLfWTfvVsHAkbhAC5fFyWM0+PbegmF7pojRccdXearrY7XszWLR
/95ftqz9i+lt59RC6yZq1wtcT7jYzw2N+DN9lJBK99REc5AdOEXE/lQ2b95dhCDCekyftUPjfPc1
LkfsBmUcC7r8XD783V7csGWlnPqgwzORtXtf33cQxLZu2wpBbSbhqhv1H5Bo68xjyQQstytpRLqD
IZJPTN1Zk1g/MLaYz9+xjiqYweoWIGYjgRh9Ho85jpYSNqQKHNRq/u4+aed7DYLe5bKUmgaDMwkm
27Y7SRQgLKelozClby7t10e7sRrnFOA5lQIy0GEm6Meoa0N+G+J2n/Y2BMDSkYd1MDfdwcg1q9j/
/85HFi8f1MIVEtgCPCk3BNt5vsDbCOHTniwMnikwZpwRPa6JIRvdJ5h6LsMHmMKsMSUaDUyt2T31
4RgBDMOyjQqurSFpz9nWmaqIHToIALL6MHfLMntYl4SWVJmTuCQCUwIz/lGR434TZspaW2SSdeHL
Iu4t2tB3EJQ6O/hbJIIDcf5CHpWNJfBhulWQq7RjM0sadRjl8a2lAlJq+yJIttZAd7xYg7sf8UTN
qQJ7pQZNYnHupbWIvzqC5zOhnuyw2KQrXRZYTvqFlqrbWG9CSyH5P35E0+GRFj9N1Of5/fSPhPKX
xwmbS7c2/HPSRZ1uQsAfQUJpPCe3W6cJ6AhSEmqRESMBVUHThkZEGaopznBsTp71Y/gfyTHN6WdO
69PKBCXMk/tm3iNdC4zgpOw7qRzPFKPH3b/7MoO+ckiHAXhwKoaKwDKo71T0K3PrI1SyYf+qlr1A
bcusvh7nlKxnaw9XziAvrZQAN0qLTf0sT6GgsbFeyGJIV0XXw+pagO2aNAaBCORd7reToKlWjV0f
FwOckcenc6AZ3x7/9kWFMBKtPzXjrdUbaH/sJrz8gQkELTJnzXY1e8Qx9cVB8aoQkL9J3I4NyRio
5FGOz/09d/kKtTXAUr29MTPFZaHbzHIO0sYfmt00wvnscRpQXwpqM0Xxgm9VxPZ9gqoiD08fhsHF
tBm5dadJe/1tIenyhOMxpU2WV86cUQK28i1RPSrlhDMDjDfZ5Epek7+nYWW6/kbCIsrjT+SyuvbO
gGrnb8r0RiPzsjtVmbWElIhlHUiBU2+mJb2U6SBhAu+4P0NvVJTDHVc6v0WGRceoTn6rRmewZcmF
oh3cskBhC1MzSp6xBLvgiY+VhNnEmogh/H9i/mUf7tWqgu20HlQdnCnbdPnfKkDmPFmJt6oECBjg
Rah+nHfAalOhYMPWrqA+TgpyUtEU3XNPSszmu+aH+lfpTKfY0K7eXfBXfUU/T/3yRkKVleP4/PwR
GPiv4kZUocQmUTbTmm7hkYmPyij1/kNtmYyy8T2xZIBUxdXrTqNoMzeJbHycEOOkrrffQCc42RQj
zFE15xkgL5itc9pReGR12GCReypZAml6AeP8hBajd4L+AUfdbRqKcv38lZcW0lvvt7NbNtMPYQxq
QXZrT4Y210pUaGTejpXp1oEy1OBv+cDek+F2XCSI0vOSDzn6lYpCOoGffEIEz16KULom6zRQMmjd
MkXy9Mx/fscDWq6+bkx4svKLxOA+89aMDe/PinPuWJYDxrRPEj60iA61jPmrq4YB5fySAC6fs68V
zKVTDOGVw+kvkIyZFfhAB2/MtD8XvvJDjOpEVIb4Fw5YYS6rUpOoMwxoF70ejOUo/VHyISifFIfj
CgyqC9/BpgrABkRxykzPvQeog9jAFRK1thD6uiG0FFCL41+vaIRMyE8jHORWuoYyFQXI2iqkAwqr
xNPLwsAPYbhFqBBI58TFxPPnJNDOzv9rqpYkP2MjgGouyUHZsud8FAXBo6MtLpibvvN+S004vvhy
bp/3YfiJg1AMDWTEE0o+OOTIDgsZk/RirifUXNfftAAOXdQiWueAjBMNgkACy1Dfj6SpXJ8s5xGY
zf5l0DqCRYeWQnEkzG9zh3cO1hdZ+JZOC7JHIca7ANrEWG4QTwpcJc43KAMGNF6rfsnwd51r0sgL
ZAixl8BFB6ouZQ15Uyoc7KTk1Htj66eKOxjfV6L5E2hKd1sLNf1SUrDxJTVzL04yb869T4xXyV3n
PS45ikNymVItRgKQ5LQAyesiS35OuKFCnz6gdr/EpchhUeuUh3kB5GyzOqJWIQzF0gkpO8qjN5BN
LtTGVkYU4nGxjQ/9z1IvhkkyM6gwzDc+v+ReNAECuoxer/7R1iXnw6yJ9IFY4a06EVVcnDAWS9pD
pyVJ9zkVUEiVu/+4ZcfKN/0h+tqk1jb2ESiBiySDwea2nPfDnRnESaD6d/M7VQ2al3JF1oWwLAws
5k/ZUnFoN6y2JMzpxWt37g9PjUxgWbHFDpz96L3syjj3vxgBlHM+cdBYUQxi0WYlHPIYpjmsK+qP
ebfm4P89VLvQjsFEjWSqaYr+ajyIH7POR5XnyTQdaZZ8s0XFjn3WqS18Uv8AKh5kYvlA1Mn45Y9H
KX9YuQtAMi97Ot/OdrgF/7VClW6wCL80C95KTDiqMQXRdrj266ZVqeo3qQtf0GmzrPfpkvxFjH/s
sxqQnp935HgF4drBwh3ZUCm04+hfWoxFdXxczp8NjLXC0Df/OSeyvOXLXcN1pQcHKywyAOsBIViJ
I1GNpr5a9BQogaJRslcF1r5dbL4Sk83rssUfPn9mfHQOkPmSv+wmrElXAMOZCt1/fQxecfXENZVr
P/36Wq/41KW3900PuNQuiEXlaUGc6G7S6ZBx6qlU5GfNYPYRCe3rDqX3xu5pysFgVpV61FSZgueT
imePdAKlXjZtCTS+PE4EuTYe9xLBjkxH4GeBIHO8wUEIaqjhQ9E6JQCMomD2mfsgjhfwLIZEypZy
HC3pL0O6+vUAfVeF0Xg6+IjjCs6i8mU8Z5q8DmvTBf5va+h7/P7ZAJAibve+oMg7y4uzMaYF9WuV
rqY0N2D/zRSZXOWOuoz0Hu6Ze2H//9oe8kKKJTV5vOoSIPxleEQyJCBSr8A6aK+F1qBxJ6bXR0Se
D2reLFa/VeWGvUSiVNnq+9o10/Yh4Ug6ThF0dOGGaZ13IT0uWv8uA/j8Wth8DlaYXIrpFp9jUskp
C5rux6SrPnn4VaRVHhuML7NQGusK9sxGGjxSMKMms6e1cneFXU3CbfEYyoDpHkc5ezx3q+PyI/kv
Zu4Otj0PyONhQXHiKL3C2UtPGX2GqlXPfgCyzOISATqA38R+6MjEQ6waMXlWHTf+rU9M9zpejjyH
yh6DsamQ3/By27/3je3NtOvldhn3gmW0dLBnC/xmOFg1g2hzPj8nzu0ZqsWFtP0O/nY+JbcAACCN
HKy+H6+dIQIceQnWcMu8s7FQ2HBWOlwKjsNS2poC4cIUrjeJrUkf2WFiN+owtDtAYI9s+8aVdhzJ
zmhkki0AdFQ4DZAo2bhO1yaVQ88OB6FJ5XNT18bbrOFiBZg/bmsCQGmxKt3DhPacyqXpqLuTpzc4
iXDvidP5wgbQupk1s8Rj3coRHXy/vbZoH4jWAsKrp4aFOI2TpgLyDF5iZklij+h8NL2/RoO27Zz9
K/yN0+71QP1God/Ku9AsU48LIqSyLXcbMeKIt6eUHIXMR7djbjcung7A5kloNfqtabioaRhGcueU
+SIYHKJdaUVHJC2ZrU6JKh0jPcCpJWJk0/Ln10uyHNdfAhC/t4efDlRGG9zMdOYRjbtgeJDO72tr
YNEBqZYo0OLhqe0VVntnsZhV/uJQivTdCvTqBmohCZKRD6hfb/9SzgT4Dyc4OhLFuMgiar9seVQF
6Ux4dKwj3J/BuLlvqPOYYRtVXGnimLSrMw+lEWNR8OaQtQThVx/151yAxiFWLRAYGfVoI/FsuGmc
I823yVFyzeSEj6BqR1Uz5bqEqzdGPwFLePyQKR2MIQlB1vk17cPUnbnebUydKwAMSMoZTETS2zaa
CtzdCBNTc88jMXMVXWWUQHwibaV1ZWK5oqkXYv2R8Ai9dYQmn1wstarUzRS+Fi3nSsi1EHsBDU6Z
vRDU7dVYaVj8Hr031ES888eqqcWIQn5Epl3f/bU1y3cODM+uFninDCczQaCf3qzNcIpeDuMu7TGy
4dAg1RkqqJI25gHqW7UNrfrHZufXJ/RWk9rPrJtLWPeK2d3iNm+YPXKFCP3TfLDgJaECZJpGYQc7
FHjhTu7DImzZUznrtKgwYKx3UAe2bhARelVcmSEfOOhHhT15Pa5rdGK7urmX3m516xj8YU/Fkz77
Tob82599DOj8nbk8ii0DPBFqb7JAXRha9LPV9ee8m+CqoNLs5ibnDhN+CI2NkS90z2Ia9ByI9EdJ
tHreelhbN1K3i5GVOdlXUACFOrsV15Sjk2DoYkfLwHwAgikfS86KGLUEaiaXxLfbsdh811us3iOF
gnEo///9Lx3BmjBWp+Ar/facPrkobCddgKIdAsGh96SygfM/J9SzGB1n0jzbrHOqYw7hY+xS3ncA
tKmu+aKfjIl2b1zNZ2vduo8skcCbMQwA+6QEI5aESFt8hAz49C7iqs/tOAdrlh3RDSAgM5sVxmpJ
QcamXDW9lVdmCx4j4BduGKhMGqLlLp46jytjolmFckNjDqMAZj8enJy+U2/ECTWoSeibMxP+lba0
9JzTmpciWdE753PTzPv971jfRzFCitctxkc+ahQm7GPfcpi6L5uRcDHR0JcFC0ZXUtyVAzGMBfDq
1Qn5cKXd++mw170Q6B4a5uYhE+Q5dzJi1tq9o3WE95Sf3G9oN/61t6F11v7Ob5USvCiApj/Uk6Kp
+t/FNIzcfyXT20eY+3Sk3BQUZupdovjfUr4OS5fAeQ2nFC7X3tUzy8UywKds/XGOt5ZCp489XWnu
u5de5QW13ZYQRCMeKAvFj69PZ81DWAIGqjnmLqmPzz3wRWL4NYR4uE6vLDaQRokck11fcNaQelbf
Clee/QceMAf4MHxQdInQcSQ9l7jIyYTgoNjd/ay8LwMPN9d29gK3c2o9iqWmkTBljkKcQqneTP/x
XDQfaWai05utaCRKNWKoOXKe+By4MN2sqPvHKNf36LfKZhk9c+tfQwwWmi1wabsE2TMEEeVjym4a
mRYgcpPfVLOVZsODHSVGfeZ370R6A2HEgM6zcv6icqp+P1VjDQ6UGfKsIUXulwnn8LuMcr7gyKYk
rZUGPTmxoKl/ZlZ3OruuG505XfoQ+rOLL76y1vsVrb+FCLR7yURXep81QKy2VWXhbQKDokX1lmfv
qJ8/9fSAtZYoXdnaVAR/uEgSkRU0rcvdv7rum7Cq962JWWDjLWmdc8yE1g3eV/A8AxGUbjzztwBK
P7jCWsVXQ0wBlI7rE0ZnFUM3X+JE/XAG5sIPlVU81ok4LfkgnrouoXKJ9syI9YnJ3+7qvGlNTOLT
55jbn737R4iR9ERlvv27UzSWVEG8uPLozsnug+kaKmuC5XvtTCl7o9PWnEtT6BPG7OC61ylcLmOX
M+jJKdWVpvHlJ8630rdqo+Aox2nz0+qsGXB1XbPQmRLl3KvexB+Dm7vi2Dt01SGh43FhvAEBD07D
9K36Gp/iAwx6qQuwVf12e82D8Msy2U3kAdLnUjiPU91/Ou/5to2PrP60YJFoF7kVF/7Qn6eiATE1
dOOAjxDcL+c7+00wrLYZ9O6ZwNASrXxJInuX0F1PP02lJOjq4x37haoDuLSwtMF+ujJxXDlY7zcO
AGbGPI/iBCDa9RZq0KNNGJ4bxeIxPv3PreOiSzhaSttnNYN7WwyiDEnLF2G7MagSwUYk7lpOm1/W
tiOAe0jnTL1uVpQ99xVn9LhaUT/k7min9G1CoqOuO50otXmgogIcXGcXQD6OB4DGsjZ5eHuD7GJ4
RKlZRc+lsThST39HywILEBh/HnCkFmq1RLIzrSjCxiSP6H3OAPrb2OCsAlXav4kAMcL4s7TzkBl+
5uuFSRkv+JNdCbRiAYGyFXZ7/O4LHtE9zF3NzdQvevviw5wh92r+lGdLbDD5jJnY+gxQseCe66rv
4+vG+gG/u1iGm4jzZ6KpG+RnLl32MXHXbPLcFSEgOMpxzR6rcYMBv5GOKlaDgCBG5xd46uuyjAs3
XskvlVykm4VcEPXM1oaIVIwIrXQqOfVLg2EB1bWdWkz9L+yZobIyINEIPK8GYayVdXE5ztw58nBH
mA1LcEZ91XzPPr208vmxOdvWeQXEyWnCH0L5XhvCFggjbHGO0d/EsvV+X/TUGXtSytW74QNsegnl
/SM7+d728Er2x16miHFfRtXQYi2hdOejTPRx3Yh1JxMZIOJDFpLm0lRYihVxBgrpIVquuKvad4OM
FO+UBXNX4BwxIfIzACNIiw/AauOf+OoMYuw39i4NvX0zer81VKTAeyUgF4bLYGmr39iAGvS+YuxL
edTlioak/e/B+sjogLsy+Ow8PtuY4KZJseXaEFFHmAo2Qv9gLlp5m1Q2kNLL4ze8a4ylZ7fjYpaJ
Bq4OhXorOJKnVz68lFjelFDAvPNvW+bJmQjCoeYtbaEvTOXn9BeBaNrvhhtJ1P8tRtZQ1irWeci0
D/imOqjN25Gd000kxHSc8iomwURyu++N23qlPJAx7BNlHt1edvEHuPpGKRhlWeqTBzqB3AZgSkUQ
S6VQOoqJA0XTAGwy0/+OFAdGXf8uBGMbdiWvnappOPFy7EA5AQOfChaGDNgt1ihdyomPZvX8/RIT
hwRgsbOFxWKOEHkHOx0ySobTmcAr+xPE+6CVY+DiyiZT4g4jYO7SjBlAOr2wzAhdOY/BpRyzpgJD
VZThQFHbYdmyX+RhD465Olu2L8u/ztgFM7uyi6/kQEHLyv15eyA9k/OxSfTgBkdKVwlBumz02ZJY
EIAK2wqVtVo0kkkFLwZ7VqUCNnCJtRCoDmj8fR2tNZvuTsLLRtabY5E252AbiOVimwSSY0MX2fgq
YwTRnqiX3IxTGNaUKil+SXLsL4mzoZRbQQvVgqHfKNqK0z2W8DVrqmcmiWZ5dTEsnbfyBsyt6YwE
igj5QhgVxGvrDYy0IwMDCuMREiRqtrPvVe/AbD8+qI1nswtjj7+ukqgB4nlDOfzSnhSBupqXAsLk
guJ+osv7HgxI3v9Xkv/CIz5NjvBFOnbYF2j8b1vHG5xQQloowmEYNEofPLBcvOf1ILaUiSFC8BWR
1voJfGzb2ehUhAOrnqYuEPlFjhZwZhuyfeOMxNYtU11UgmpChzJCbuqSJYcneG5g3vQNohllcsXc
kX8QSUngLNIKcvmv74RQFWIru/TV77Y0jv/+bSfPTdikV6LemSUEpOr9XmxtZmJ3WE0/Tqr7m0kl
3q5DgBc2BxbWD0G1IuTk7BDm77OW+jNd6VzAuKTDsjC6CWTPuBqCesRR1SSn9NzRpMR4rII78izK
4mglldg0E9QV7ElFqFqfwp9j8hSPP/oMjlHL7NzgEIvdSyTtuH84Bano4Z+a/9DJhLDKS5e12pYI
aGB1S6DgM5PPds21d05+t09/4bZ8qzZQT9FJLL3T+xOpcvFb1BC3Xsw7eDWo26W4sfx1TLBzDXU7
3HdIDHz3sTHlKjDMoasy5yDVEtAlpteMg6TUcQjIl6QZ0jZPv+gVmh/tUAarGG2FHtdat4JTjmR8
wcUhYblH0S1MY77BHNsjoysH/ynOL0t81ABQVS6cZ1iqn6S3yBH65TnFqZcdD8pzFxi6cT0iq6hy
OtZZzV5L1vhtJhkPuEsBzTpRUG62LeMn/yHegv34Mmz0vBpN2PrX5QTp+poDYmaq+9gV5OBfnEva
7fSlmJ7KfrHSZK4bp2Ab/dSqyOODNfirh2aklVECdb+EoYuwRDtUTopHOLljj0ezaemuI8uuGZY/
ikwZiysU223HbIYeWNeD6Y+mKz4R7ro2Va3hdH/SZoW4O17veoNVmD7xNYOrasD7QCGQTgy2a/uH
knJoty71ci8+kvHa2Qxl3WqGyjRWuk+3D34GZvPo6gmXBUM3mRJvCQGs+20eQ9NlRv2WI/lLscEe
g/tQZg5xE1O0Nw9iyr1Gk+RbeYh9GxWcPXET0al8d/6wjwNiLfqhH+A6lq7L3GKeWGJLpuogtEX9
RNRaqn1BQTyPoiF7xhSeMRH+770XMtpW7tl85FLvE+YpxYZMX/AG9Y5jKsZvZ+uy6YR/aueUnpH/
ITuVb1xUlS3o6kFP3iI2/XxXYqEAGYCvZt2O18WlzCb8WoySEDKvRO5uD+RbuMgsgqFVGed2eUck
+mU5+TKx5l2MuDIPvsIAZLet2Sg9MysEivhhL4lajvoHlSq/iw+cVyTojVj2heDNKBv7S2QPEdnM
gh7G0sNrIh20LLqRxZ8iqhHifjufKxA9Xa6gCiGvGFGfGqwPtfnh8wgbIA0mGw8PqxcLobLgsRqk
3NHP4bbAnhBwpRS6KOra+93q00f33P00ycoyn2zf45t664u1kqoAPfS/PiMLtL6lKc6SSzbO4JXP
E6spt5yj8S8eWKHWjygYnrGTwSOMsfVwgp/YQsuUYbjVdddNWkZo8HFlMOTW7DX8lBjIIxtVtd5n
mDcUzRltnN2u7td1hgZq1SC7v9OrPyzU2uNq2qqxfOOCOTCV/LCrFDTXGsIHIDlRopfjTYlg8B8a
L9qOSbPFxzRXDw6mbXDPcv9CwgnYPEms4+m4hKKDSDtLXu2ANPPd76M6WKh3f2pbph4X+Q1sGJfn
0l7vcH7bhtTrefY/W0af/e5/Qr6Y5MWz8r8bs6FAySRVEpzsfGIqbz+iwqwjkA2ZqsGVGsRuttn6
tWq5QsMyAUt3QlyP4sENIjVW8Er+zFDOI6SpFfhbrry2c+CXomW0GKJc+0ShnEveNAwUKQs/afWe
zidYQk93oEePMYYgNp1Y2B23fKWm1bQYkfgtZ4Umfwed6X0lTeW3YBdBUFHJ6mlCgN/YybyfZFZA
zZGnz35sml2MqR5o978CXsr3Cc4sAERS9sd6YOkJBQXSQuG4WIH4CBtzzKV8hnCdCP/WHIkrV6NH
ZIv3v7Ts9RtlFH6SjTj2hW59TeCTQ25zuQb2QfbRx0s4b0t5p5flivWTgBc2CLclDkBbUuIs4YDt
MvCFVaZOiGEPx04uxpIdhvE5/Kqq2m88HvZmDi12hadFAv0yRiQ+1kpMgF2gZ5LNcrQ03lbDEvqx
n9UOGbqEyLLyO0IPJY0WyTUYBIw/mUIjEuAy/opt6WNFPQ0ayBzMMZSSCibL4yci3iL9XdaIWR2i
OukCmNtHvUm/5fCPhtkHZ0Psmwf43Sa8byiBLjFeuScOqtMXgHeGranDpuY9FbA9FN0V7njmG4bW
ZptKeskN5gSqATSKHXsAzkGKcVjRs0qn5g502f9qTkU5Hbm+3Szuky8jxLJoG9v59oi1eOSInmZT
t/YS3rcNr+Wr2jDa5vcrl1pj92ralLVu9f5JPFGwC8oNiXznmZ2aU9fJWHG6Hbm987pVs9rxC8D3
2u7upUhhhMClxewge458MCVRZV6SKfkykWq1D8HFVhD0woz6uTIuEGGi1WtLPqKsDvv32iYiKNFc
782jrh3kQZ8qPDD8LEJ/FEMFRu8or53rjL61TaCGMSK8k2sqH+lrg3hDriPHRFhygbeyPgtOlVpk
LcH6/VuefpN+kRkX/VZxfrdukvDd0Oef3C8qPWJ43Bd+/WlP9iOfJlInJBixNFXX2vAAWkDUnYY8
OOfGFvxFWKkYvKfElQKvxiIec5OGhYQ0tYL7Ftuy1Gtw6dgRmf2FYPz/1nn/nIncvcTFag8xzm92
9nkPspAcLPTWZTEVz7tgRnqOB7ycwdtXdS1meY2wiL63rmx/+fqbrmE5NdKWyF4v+ghKsPJqmSgL
RdN3RNjPOdcDxnwUnAuA6+AWIml2/yhRIj03wEFNHeA6ypFyDTxlWipc17jrlHFkzzpiv/4Lr1nP
hxYhk39mCeRLiWDlmtErLYt5IwxcqhhighcgWhR8u9ghJkz9vRfvgkmuF0+Y0krF4AYHkDnBU2kV
xSlMmrfeds84WHQAvT/dtKtY6sKD6Xrmb3G3XdmKOmKhcMyZM9IlDYM5um7GAvtjBCEKtDL2B4Kp
cpJkOwqjL/8P7vgSTnOwMb/Oqfh/dWCVZc7wHTP6ahhDnY6xgcV/rLDo5XkztDdHfLjRH6p638pf
5E5TdH0IYb7BQRDSQksPPJ8YNAWWpDOv77Qsb3l3KmclFQxbruzYL5Nd9TOcOv535Fcd8bIzHKK7
YmGkDdZC+zcJQnki89zNsvPNkDtOKKASYYQ2BSDQ6gzaVIImxa98yFvPpfD6/9vOZEvvdouRoHW8
mfghLRt/T468hJQebd3UhOrvYlrCLGErsofjYpRcJ12joOfTiw50+/zuLKwODj8URUid0aux2D2t
aPzhaHQ4ayFOsaPLagm6AbGgSMmKjKRlBwlOfL4cWzLsByzJjrGevF0XlXx3nSUVu1bsQG6Bm6Bz
Un6GppTLrrR+BnZfDf5a6zzLbnYWRUtzajGPHEkx34g7Ti4sF9batyMOSTm6FpMKAGxoAbj8kmXf
GBwh0C5lj09LTW2I1fseakxLZGaoN5PsdEcSahTqfVhudUDjAkzq2XI36IaIhuSRLpBoF0CCg+4N
K4MqgzPf7XIa5jQg0TFRVcHWKk1m0dcgA00BwddzMlrdIGs3ZFBBxTmBA0G99SO6X7gnv4Piy+uQ
da47Z7JMn7NVTG16HV7i0KmOAK0Eih4zhjgUwvEVCWkm9bkOHT2L72HqnsUSAIpAr9WH6S360DtS
KlFY6SIQM3argARNVfXuCAv0Z7BheQXVcPBQUtFm8lc4zsRiKdee0yZwIjv/KNS4N3FOPWbXlT1N
BjhAnvxXSRAuuZoMM3Fiis88lR+HQmwGKo0N0aZfGQd+y/ylKMgBXE0OvUuT3zPupDlNOV5NIRwk
r7G/3Db+LfTMqyVq8KgVQYmqjIG+xVjWhpAWZtIWAEv95cP6JyO0WOC/y0qVjjcpaHFKobETGxTm
Vusy8hB8KXruM/SQk4cFpOsk9hl6lR0eGRN1x2q7VKjXVvLpT0QZxfEnBs3umW4erreVvd6D2srx
mVGrTlMH4xGIs6VShZxKLf+kgEsjxUJRW0LoIdloNluf/1tUjVEghcrv/TG3fctAVY0BTHWS1uwc
FiFuVaUOV0geBD+fUgPR+CufUyy+IycRoEEzht6rxPyj+1hdXE9JOsb+4DWQCaU0GNntSmI9EpZ+
l31TNxoWN68H6zaahj163P+mJavMekkLGeMacE5TDkF6pnobe/9FHaf255ucvcRlIm13tYJzmnnC
rsgPm/hDGSJwsb0fPkTOHkO1mEHm3TODIbEl0KCXRfJn2MmP0MUfFlVk4KDgEYn1XcQdOQpwjOp4
p0qn73ICLqUem+VAhjwb6aqcRzrKV6rJm2SOcMb1SOACkTH4dEhpE4QFFKiLMZA+ZupW5jSZTPss
qWQtf8WAS47hck1FSMCMWhjUOpcwILN2ru5hAVOOwlaVKMQ/84EwdP9Xe0J/8k1ujVFWe75OU3T9
JL1/rVmWzcVlQrmwTLOckeom3WxTOJj3xM+YpmuOmwrWOdFLmRS/YrttGz/vuPzQQTDlFpxxjvla
yflky+vpmJUhygoXfHG4wx6xU8K+tdb3nbwqO0TM2sD1OsLWtOzjM5f9OtCDOCctN4JdvblMUtTI
WEtf3U3ie1blhYiBMGzaRvXLvtHzOoohyjPL2dpWwlP3M0vWCodzss6/4GSKrbryphHStzkUj6df
wnFLdIebL8U42mD6e4vQ4AQBwWv8HXuNa63vjccJf3mQYKjI1aSTJbPgntE0+n6Anwm3ijpYmCmc
NvBnP4/0xsZ476PG+c/npjkV/OIr9mjzWVwFYRTTwSqPA0R5WBtAl21ElYj8u3f7vMEFhbPKo8xr
Q8R1biqirxoyYs3NqJ5ocIArMgIavFTFYow1ewDrjE6X4NwQldJBdNrDsTnGL4ZmNYFy7ZnA1bE4
mZyQ2Rs/SQA6Wozws+ly5t79brlaYiVMOB+G7MGgXL+OVzSfqkGRcKcGXPsKlALXl3CzL0ZXpNAv
/jrxlr88PxzBpmC1k4PL/iq6P17cBhv/aedRaa2n+EaIuLyP7dytcAdplpnqYzu1xDmE8PO781X2
iuN+O8oFSUPgwaa6dM84pDnmOLZpKdD8/p5cWn+ZQ1mynLOC0XTk8Eqj3/QVXbw/3vCxn4szNvqa
wS54mniUBb5pShN9/ZkAAYowSysUQBAhO6QR9azvue8Bu+kLdmgDwofCU7jCgU7+ZJ+XEVZ92AUg
V0P5H7Pbsvs9InxDHOQ7fvrXnS/SNPkSUxcjjx6qgIhPZ48oXVWZ50uMCl6sUKgDs86n14KICN+U
yGaqFCPtO0IidolPd4KyrpuuvMkVMigw8QuBQb+xDn43J3GaQLYpn3Tqg+zRpNtAuuFviwys2zA6
LIOrm+YqQyyCA7bckZgYVI6xteZIo9DGS9DQTKyC8/3pompTQDaJRnMIrPMVRg0m1WsU0J7zof4U
944Rr+1DtMLlihx+7VO9UpYS5ulmFP4Rq1H5VOgK9r0DB2R/IZOpLlEJQKE1ZK2pFw9t6p3oFD/T
1zhd01J9PndXX95jem/iVKeWzQ2qwQJvHfZ31tif8vNjr0ESO34c2bkIMsAN0hNRqwtsLSaK79sD
eTU77KMu9gYKgjCfCkC/hZ2q/M9O48n+OTDKa4DzZFKLafaiz0Xv1LvKXRGxGyLX3tnlweL+dEv2
GvSiWZhi1u+/uYR7OiqGv4p1hWjkkLyrCg62JfunIHPf8KZIhnNKpywLXm6yx7We0Qop3ErslxOj
hX4WHVv3IO5y0zmTxA+OdHkcy2II85SWsdZADZeO97wEAtSvWhLgcNdxAcZLbN2ekkfx+JeTb6r5
4y8BfQ13h/a5m1EDAeier/DZ2ImwcDOZ8Nnd31ZKdLZwaGySkioRvNuHHW39mQrRbAJYxlZQa2YR
CtYOnhymFTKShi14Cvh6/pRnZZw17+sA8CZgJPqv5LQLLLfwfEmeA8DmpH7SdRQG77DqzgfclWXu
H9Y9GtGi4hilUdAJtntWHPSZwrKUlUWzOQ1ihwYhIDbbtGWpRbe9Kb9h6VRqjv+u7m4TvGO4N+Sq
nOMEIPv9ZHk1KusqoTDu2JzRBvm8dLDYSymYiJ3M72BpY8+IfHFNe6q7lyYTIu5EuWnJznP8Z5rH
GulePan8qg7HgMyYX5skNiE0wT1xZFQx/4eqFReMD2mQ/EkGiCWTjMXOXV58fSl6OdJM1zyCWrv6
GJsyElA4EIFmNfWF4XfqBU2tPUjr6BrV2ZHPxbbmZ/19tg1YMy8G2owG0yewZufrae8ljUZ9JAJQ
wJnssqXCigagFWxJythVHG7HccLSGjUKemrOIxMXamph97YUb0AyBv8h+M6zjsLSktkPSXR4UDsz
URWghm1hVKAz8e598C4zrmItPm1xLscGc/SAgG+u8tVFmooRu+kKwVQcZRqY+3WaTd4OWY+tr32u
tlnfOd2gMN4YOLaDsXBF7vMWg/FyQCgZr374UHrWbe1r3cFZ8sgWlYmNaisZELDKEV8BJ9KBtemj
B3JES4tDHyuEmiqYFRanons33UnfnovccjXMpIKZuO+GvOk4u1KgrZqcOb99AviH15I6NQy1t1ji
LN/tn5raYWvk9+UB2zxZUp0RS5uIGq+layLxnQnpViGKef/wXMsQayuPBoXUQAohR4inxLXa713+
AWw761w3VaiF5m+h2P58hDO+wyi0maI4DgMyTzm6Hwg5zgv0lHoKiZ7T7VSiJHq9FoeZOPIi0yeH
4itb6MS1xPrTn+suUJV9kUTl+YvdbbMB0GbCnxDVUIX7ZN+20nPgh/6nbZskffCF/uHedx5gN0Uh
2FZphU/I4RosrJDupxw0VQR42Fz5pOnQLYtuo81kdtYPApFjfkrz4q2XnohVIUGxYj+wITdIIVd2
hSFD8Uzm4Z5O9Bfl358iJLUeJVi7uHCq49yqrwLq4/KckcvVxZCyVhvty2Zen2UblaGkzCau9fSy
dRFKvnAow+iURLTXOPClXp9/DD4QkX6/CvWtNbXTpNYMfI/82Qw5+RzhqrsWgDBQUqOEpjtC5U8m
/vHM3cRpZCcU7uVGgxq3IljrzQ6WP5946mjXZwW2j27Plj0pOMtWMBFlWVna0aARGwJ6QCP8eS9/
XeikHaUl05cc5f5QMLKXRuUKJmaTi9zpvYu29BvGMZK4nbwk8qY2nHqTIKhYdPuURdC7090cBBDx
FmUO306ZvrBjO5tpCmswtpBKCicFx7ahrdkcZqL9/Dw1a7x706SB78Z4/jEewjlWQ/NE1hjvU7wt
f3sxBX/CV5YF+41i5TqGRZxU+V6n5FCOhhy19zno0ETb7H7XST1rdso+CGDTKjJBN36zpnezOkOD
tgerK6x2Zh3i0oxRX+sQbr4TE15YBlo/uNlHyLaCnC3rS08Xv/F07+fGsdBNAeecV83zvsqlVKzQ
nxvfgeenHozHhLcrOKVAtGbhMKB9m8qhUBHDyp6rm+Lhf0NoHWr7sbquuBldokWZOCgBs5E+kgYu
5LDzd2jfUGuaQy3oDe/H3wACvgz7FsRHg5ddTwyngHghqtL+6NS6RhrtFJL7U8KCWEmW8Fv0G+sR
amdhI3byjXcgXAL2fgRqWQQD0gVII5dyv2v2B0CfdKUGFFuDtYWrG23qIuJyUfhXRE59+udB8BTB
3sQokvmQdB9mROWIQflvVdoM4yrzuLqrShzTgbBfO7VVaYbxJfpeVhlX+N5pbJtO7HLZaq3zFzOI
NwjjnPVq0PwvmddtM1Odd8Zpr86NTMdFwRcBCsFirUyp/UrodE70SM7cK21cgdQ41TmYCDyhK9pq
X8/FmyAe/jg+j/3wNfJ6N8syUsdgT7eu3De1vhdbwHNh3qsuinvtw1++E6Vo7zAmr53AOK8AtSdc
KUcbQxo93RiD7jDo0v/L8mEXH0V2AuXUcsi5AVSGYpPd9ZOogS9yORFayr9tLphdCQCi+gG/R+hs
De7176Xj6aiunT4HcBUZYGnY3kfySIWW+xb1729GhMw0b58nUmw9ryiM3sWt+YtpgR1p/RVbTrQO
Cb3/47qKzkKKn3Q1hLOpFDCF3dyR9komX5DwwcnuWNIQ0YDEBiWQASWHG4l1NjwXqlQcMZY+iIcX
DtfNxgKp5UAZMqQaLwv1j/zEZx519hUuDALmATidIWYHbTnUNFU7IPhEY2kq5CPRVXGahQelm+jH
5egc9tMGgJhrmP/PuvZNl8iZuh2Mef/ABLjLoMXyHUVgW1EfDiDL8BW2i9uOONO7Hmv65cigGQkP
qg1g49Fesltj1G3ueV4/cuIxOvVe888IXerWdt4fj5uTIBIM53X1KKfPuMyuGwzf64Hnvgbfl2wT
J0cHeboTrKgJHcbteKHy2d4IKLmkYU5tFbsDjP3M4Fu66Hcj6uYA7+56EbICsSiu5B+Z7VWH41ON
LGaj6rjl2TpDgyD1DZF64Th5bheTcqVSt3s/7FTScVq0i3U5gd8EZD/UOHMqCi/sSc9w2TB4crVq
tog3FtnFg+ibpoc2MIpmxLt1fWPGfwPle0PVNVtuSoRalWeCT96qE3AZLP7n0DXUAcfEr6Fvh1zc
pwyOXTB8O73TRY2f4IKpAZk1piL7TejsT4unRMKuGuujpjmkMeVX7j0/kw4phrCHR2MT0kxwLC7H
zx1UY4lpzFYeayZbVQ5OMSChp297ZQqUG0xJlrOdwviBC8Hw9qWGOWfxQimewgxUg9Zg4MAHmoeD
ufYbhD8DmNmVP+AESIA5T5zmZLZldMVbUlOv8gIoIpxOYD87yQp/STkqBZWNRZUJ8VnjZMZZmgtR
/1/q3Mdu7rOQiZTuCq1XsT1NBysNyTz6f6N57JlYS44AbV7yUaGRozpYc61kn3v/M/ilCnFEJq0W
eDZtfWQ2CqAmhZHfdVVmMpQkswEghbPIJ84wGKRXpvjYD6z9Ilpp1Q0P8OhfY6RZe6nROhASxA2t
VcSiv1LVWps4b1d8mymTfPkeCb1tY0voWAepwJxqL9yOpOhknEeosEdTuoEoOaD31dRGHR8UZdJU
/fdQ8FuKMmyJz64r9NLDlNO6ndqllmNJ8t1QHndd5VAWKSRvuIAgHhmo1es6E6gQwllIxhHk/xB0
gF6Qa5T2dwSUm4nFMEpUKg+14jdPMDzWEFsp101fHwmdoMw2xflHPneeOEolQJUlCFkhsPbjflfv
1W6PAuj6konIDLkFpieH66oZQT9zCsN46tiZMbVpJkk+thHl32SL5F2dAkqauxpqd5l1E+lSYe7p
1OUqUiSw9q4MEio4L844ueKNqJbgeBpMngYaMOoiallch/Pyrg9P/eWVAjasgUInJVABFq/kv3o+
xiMgLzxDcSFVXSGiaVa0EzhvE5647fJJ+OkuH6uQrNUCPGbufvPSx/DHYKzKe4xYXIahvPV5oruw
4M9Ko0pbJ+qL1a0gbjnlgKtGU5CZuNboFwXr9FsWsnsIohaXtVi0NdfmUGSv23+ooLQJYi+37TCb
oS70wrFRJXhwR4kCWskuTa2+JpTjxGW91SDvOvpqPUQLWe9IjC+fiXd6u/JMLPaslH1W6qNGnn5R
3ob3jAXjjjCYsaB/7aaQ64z2jtq3xFk3xlbI1nYGiWYFFN8Ba7tzk9yLXW2wyAwS/vRPyta2wgO2
jnT/UdQhB/BXVrwciRY3f+QmB+BG95H6A+NZkVl0a8QKP+EphL4nfd+gQMFyG9QCNKwwCd3pwDZm
+nSvtivNTYb24cvRK/Wg+lC0OqQoGepjtPIlommiomES/eePJKRQJwxDdzxvc4WCGCNLh/CkUZGD
0ZFt9LZZVELcQo5IbXhR0R37MaKYIXIzUmunHPJU77cDYCmVQAF62JGOyCyrCSdLOWp5PY82GD+5
mtXz+tfBPtlPhnsbLu6ps5YK1uS+vw7CBdILRWCaRMSnSl4Ov3Rh42QuNJSb44RT7P8S15pJU0ai
hLtyc221/HZl1EIHXFHF7YCMki7ezDGEsOc76T+PlnprNoPSsmtmd3IRZSCahkZqLVEfKztCh2kp
WJFjvRiHitHBe8mg9NlygNOlb04jpHaFzvLOzlpZJ2gxkS/gS3fX61d546y1oZV1u5gGbB8VWYTM
KqJ/tJM2A9HZMz8lYz7LbH/GyQ/9othWlqwgnmuTpucqeqY1ffsgLP9EOxnaDU8qLe/gBWvjR+Q3
B7VyxfA+5On4s7g4yAoIK7Lf7QRlF0PaCy0PPNAKWylYQNbfEsOWixySUqJKVybb9EG5OhhO27Yc
vS5CGRMgg6aeM1hvy9B2VSrRRgWb/Gv2DQr2Oi98ymuYh/Kcngkr0zV7VQpL1aRWgiw53UplMvOJ
47z/nPb1sK2rBkYcyzkisiRHBle9amscYwVvGnQ8/O944n7UF2BW69M0/+TUxo/q0uuxVhPZeA0H
0eLvwNXa7Duel0cFJn3DFcxllxC6cJWev9w6+WT4H/79q/s8bis59yX24bJJgBIz9BqMJjf0A9AP
hfZzcwuIyXmzUF/CGhSwZz3zrC+WzJEuU+KeDVU8VykGsn+R98S91li4bjjtFrqzCBU+GoW+IPiT
hrrc7ArUxc5tqtNu6MwP/ZhSabaMapCRMJ8cmzvBGFARJSyw0OsqxuY9mWKY94FSInoLxDj4Ah9a
7opFC3rR3OHXgHss7SFOtftn+K7o2TPByueJ/o0ovCA569IDLIDJQnXQmbVQr4DDgu8AFrnsBT4+
yrhdjyy8+Fpvo3r5hAoio2e+1agxtINRlOL8lkcL1hya+5nAsfxNj7r4y3YR5BME4nIdQRcbfJUx
VvSf7FXjqEZ2X+UNN53fxXooAhrFmCmoVOeBJ14GQCUIvtfUfsjTUBSla1u/9MCizlxs9/DbakmK
QTSor1ZV2VEOhKvA+ZcbwvwgfNYVh3t474UNNXJQL+aE2lbSoTqHl0x4ltns2mmaj01V+q8TU5pr
JkJlrOh97m4JVUsHIJ6Tvk6NGQLqFhq57Bz9eQq2NLx4ktNssi8DnIK7cGjYpu2ZE5hsH1CJRLCL
RcVit2rdXCera4OAKItb3A0IeBeRPqI0tzFScTu9sg0QjxKmUVoCQVcw2QLFn+SCM/fx/9Pm9dry
qOAKoDr36bNs8Eqe1goamG0UB9SEaruOETyjbJ8enrfQzPCskxljtY19+h+7r1YiKPRmN8UUtYOl
PSemcBnd21Xoa1UCik8k7xMKxrQSFjDWegpPq3ULW82ZdhcEoOWyThOw4UpzHsP9SwV++w8+Ow3z
3XLiQP5SxVkbeotyFTkptzpz8PFtSDW+TIOv0//8YeQ7u4JWFM/iQOgEfuHWKIvi53dOx3A3oODv
LuuTCx14GixuhVG1I0/BszFc+xHkJR6vBnLnMIArt9FzkfLxPJkuC8U6W/OYFy6GXZN7rk2BYdiB
siDQ+UL2fL7b4DMqW9mt9YYHisO8qk8TSjVeXT2pttwJk6ZLr7uojJhDOBlxluSuqQARP641QDkH
i9frXSJLd+fP8XsbuC9aZvCEPr62yutIHu2EdZOKSO8/6gJciBVYiD2GxHcETDDHE3vfRg8YTpF2
hbdL3W1JMFl2ovxNGt4q+ifL+69k9/j8mAleEv7NgCLpg8Sjc2KrfKEu3Lcc0AG1AAEzKChZxdND
v+i5Uc1HStOn4KkzYGvw+3rmAvYdQcvqcP3MSCiwxtjeGFSWnJHj0YFOublk6rNeg5EUhPJVXCZY
UlGjhUwOVLDwBQ0EeNQ0YDyydyLSqdweKM/WCmoBJh2BrN81dGH7MvUSZL9MGbC7LohMVIqThEOn
mtVyeUYwVd09xCfJwYxRrPRTJzrIe2yYWkCpejR0bChQHxZChhF1RY6vyJfpj5ZQqCD9uDwlAQGv
g9RNk3QBKjyNY/sWD6hMR1XYGidd+zxBI/stDsTI3+9MrpOi82VFjAuIGH833s5vZArzuW4saJzQ
ppeI7TT63+Hyp8EyqfUSgtV1Z95OsGtTlOSqJbQ+sCxMtnSt1/il7okUufPlYG1MTjqHw2HrYgId
TzvYLnoXFd6JKDNkvDvPQ8nk+LcQBDf9x9rC353qSYodBAUfMCx366N9COGMU4se3aNSKgo56IfL
zE/aJdtmMJ2FKKe7fkmwqtY6P8KfJjFIXI3OPB95AjG0vVhmLcjtPHSlKJ8H+wB9dhr1YyQ8eeHP
nlomCHhm2rbNbUhOhGW0yS4ONLxWAv1SsuRtxNZTfA1qryCSy5LFJraLb/I234HJugiwpPhHjGPJ
MFKWSWKzdtb5zEZmayNzLOj0cP2yVWwzrzg8E3Q3sLTefkzYPJ0nfl07YlpIZVzsWCMrv/kFZ/Ef
ea6/5DiWfgb8ao6x8Kyrtz07PgIBsMvlIDKj+wZ7y7jwxnbtPV0fkS8sPJkyPhQIMrYpNnk67wwa
5fIM9pAM+gsfoq0pvXoQrbTd0C9YkTJ8Wh+aBYGihoaj/se08Qys2+Rzl4HfSuesk13a4EhIdrag
Zjj2A2p+M5bUfqke6EbywdUg8ctgFnuGjtY3KcBbw0ZcERxehnZ/giPv0acw6h0vreF/rT/Qa7ZG
Zw7ODEZxjC/hYpueCm38ztEkokNZCvs1xv+PZewk6jLjJCsFbNXKd5EeW2fOTbwFn6T0WoNTQmze
MT5wwVbGzXVrS30R8BpEPKr+BSJqRlKpHXpmOKmA2D5uLxisVH9gJPmmhlrBvz9ksefewGPa+an3
trKkNo91RZQFrg3kv/K8eqi5TrPD3HDwTKCclzMj027qd3DyetQ0QDs7PJevofTcgkjptKH3iVx2
hfcUX10n28WyG4W89xrX6Pj5Jh2+AG7GgPlZhU/G4rd0E97jdRkard91f1TTskuSDQEtp1rmm6BR
ACkFTpb5TacwY8jYMaSa/eU8Zyu28DEarKYMY9S737LDtjPcoWSUFYraGawkWQEyrqJnuED0evJX
L/yCLSIBNDw0B+Jp+Lrli3vBa9W5CXhG44KLazfqAgjYVPWqyXiow0s365cO0Ci01I8xHCOpgc/k
LvtWi2DMvucHQpImBKtyIVAX+OKF8eJ9w4cdL44kQCHlD2e8o1iV4IAl/AS+CsSaxTcWbG2447ky
OALiJ3vXYPCk/2ridnzTDhiboskLkrQ4PlqWWUuGl73HXEM/Vo9E0Nzjqzu+/HxRdaBoFCHOJOtZ
ODq+mARh7c5Zpots1/6juaXhzxZpP83MqltNhw1AOOjj4Pbayw/CUU1xZQVvfhUQ+dYDTxjjmoWK
vYkIt8lhDTu11lOvonuh0fBMs2Np6IIidCJlnLlykC+jR1nGRZ+GKlTMP9RdvoVj1InUdKTTZll3
V5QUWnGFvInUocPRTEoeKUVwHrTeN2kd02X/MFbELZsrmBnmE33QayC8AxRXhKJhu8hra3hOn1+1
AdsyS0od7BoVQ/sRRiVfyFHZESUpL1pFI1KnZL/rHAomJD8Kgj2bXakUGqRROmT4qJwPwrqFTMf/
OrJ43YWr31lavWQZn3EVqM/HBkcYP0Y02m5EECycL+sE15tSjajUjESzHQvyNdv1mhcAn7J9r4sO
jTrwXFRW7bmXdd1+GW+GRG8f9gzgymWgDyKjfqgzpEw5LIOb0e+oHhR4gc6T/7hg3nhU80KEl8fv
P+GO+ljpNCotY3pPp7u9DOkBXjnlAjDZKWi8o+XvWaBoTf9CP6SwyGQUntYPcGJG+YcHPkJO4yBR
hqqEv/e7E6PdD3mTD3b6OGGQ2INqNT6tqU7v84Yuj2fCneZ3G6AsfGmerJAjbqo/bD407NOiGMYr
hKMZ+gGQiFyObM4Xyzp3oF2YiyuMxPDv11EvRHOIxAbrPOdq80Sigw3Fm33/pRLbhJXAXVKgk/bj
V73HXHqTuEh7MwaeTIuIJdJau+8EojV8vJIiuOVuTGk6/1iRe7Zk/Omcd7+VuUX6JswUxwElsTvJ
CCr0YWiSDBwmTFu2A8tWLzeJNqnR5EorMKRFxzQYMlntB4PAq4zr0YMWzoaFWTBPzqsWSp4MMzI0
NQWJn6Gl0BqnD31eSwRE4WSCGmed9nSbW5SQNNmztlbpumncK+qCr1rnZbeyejY8+ZmWxAqgo7H8
IE3QXNLY0Ah6F01dmiklVZtFtbr67b+mFEaS9J8GB8yEypMWt8OARUC43BJZKjJ3WNpBaslizs9d
zAW2ITdxbqJFITqpCdYBWPAkxp+Zy031VzHb4TvXEs/N2oPFgV0pibGyKaNvzQSVGDND2bdK4Hnp
PWMWdhNg31kis8mad7Fe67DfOWl7bN3xRAZUS3rt+Y//I+DW/E/CmwElhAMrgC1fSzGyDCWLoVsF
KdI7/HNzeyrlXCM6c+bm3dIDaghrdTetZUDH0FpUCczfQoCXKigxrcRWs1sz1p5BigMOrZ6axRl+
6rImYGRxzqVmixVG+RaGDdxvIZHl8UB9iKbTLN2lnMwwzUgNvkSb+84ITbVI2qHJmnca2xzEsioC
F6XgF63uJ/dkCgMqlmDN1y7mkic1gRBW1m/BSP+MtFsBg+iNqGRt5zAKah91M/fo9BjI55NZXBOI
2NUMOdqsS8oVILhDjWON4W2qYU86Zw4mmFhgX5QT2Elqp16k8ymy539jiAq9MpV1fiGidss8Pjk6
ieIgc044CpBmQ9tQ6rNTyjFY07ArfnMcwItSEM3V+3bKsVwlV1yzuOjNypSGK/V2VSSWPUxrLmMK
bBYW8PdKnpFE9HiYpdHsfUbHL0WDUb9HrxCWXwgfXLkkfwgbeV29cSQvWIyCgau8KwbfL7i9Qeo3
CrCdwEK5e9aBjxuEYPp8x+P5LZk/eth6t4LMgiIw7pSfpWO7b4X/Zx5crgYE5/kJuGmNMIxzfZf0
2q4EbTmAotf2W90XBbwkYT81KatvZuJnavdVZjAjRugU4ydkDxCSXRX9C17AVdA7pP4IZRA2b5Pi
nukWi6uLwtyybZWt/T96HPa4ZH+0z2YGHHA1ueD23rPW5kgsFBinqkaZsQZiQSIRBdsxA/NVJymh
PcKqrrcKfMEe5d08bB1i1XYPwuJnY6EDfIecPS26vdq09HuXhBWmMDyuLodlF/0bQJ28ng70cK4J
9Ih4AW2tFZPITi0EZCg6Sq58+P5BfeMNmjh6oBCqc7wS7t8+T1mcoXbrRY4Dt4U1w0x6l1AfuzHO
4vUHchtxI4cVu6JuHqTcY5wWZAtfXbkJOBCZ/AX27E/Fst9eESM9AVWIqHGexguhMv8af408itRY
C55WfviVtXXabBKu9n2grsYoIhO8w8zcE3sUsXS+o+bmLXaSfItYSZhbn6FdFL25t0UCoAwPTVFT
6IkKFFZCgf6nIKWUGmqJSAitHFI5N9fbhDrsk6MfYF/6spk6F8w8aW/YOti7wp1DOnqPthMWcyME
sxd7Iuw+PXwwHDrjLLxewMm9LPxtzqBy5ZDmo/3l22wiSFvkYMrmauXzpvAW4cPTibGp4wWEDg0p
RKinyri8+rSQxfHM86/voKSbtpG4DqdvxCvElLPpFWEC//BWSbyPVVeeXY3wwZro5Bx0FsCaV7kZ
oXwvDQT3ApoKGizY0on/UFXw2Rp6S7VjvGh5Ci4hbBzbmV4J19rcCEASnYgD3+ALfB279/MLM8Lc
8KQu+wd37ui/nupC3Ndd+dS1pCXtaQaztt6Z9Jvfs0rzpDxDhjYSQ4AWmIfcay8lvkaeDf8yWj0A
BUoE4qKmWOUAE0VXOOfow6PqRSbhTOF1UiFEJU08A+9xPvuDzj/nv9WWzsKWqS14HW1iBhN3dx+9
tA/OHD2EymTEoXgTon8EJLev2fe8IBiXzPD8QbmmTLjWovRjvcuPQvu+wXj3TEbzfvs0r0Fw17h/
Jk7pPgyofC4cPFe3WTK2lL+27FsjvPFfavgSFk+WFFUQuk8vgOO74O6Ur3A9bmpLnsosOh/ql10a
66f2U3H3X29B8zzfCEEGUhQ9zmBDovy+yhG/wGAedMU78gNcWPOowUgvJl2W/Fa4aG7o52pbjba2
U7OQAeTbw0yMooBr9Y8YZxTl+o1J3u+Le/32ANfE7XGggXl9Zsu/zJ36DjWZjSCEgqv1EIN11oYA
Axmo76x3PD3f8J80Ctqx+mAtTJ/L8904vO3Xg0FshMtyFxjkMbzB03/o/wGtpExEYU2gXxUGp6cd
OMPEMnuvEKg4PGc1K8PfVtWs7E4rf+PiFgp/78j9wAXdwkwPviS2Z9XE18O5i1bo2KMt9KLMgnPP
2YXM0wCJAdZ7eLDhypLZOXgkoXr1avCb3NklP0hdY3Qk7EIxvFWT89SDbwr7WTi91ZnDJ1Y97HwE
mh/FcSWxiyGKZw+tqXY1PZS+HERUUwf2ziA+p2kYVxo2TCf0YDBhGtFoJYxLmIjDKqX3u0mrFq0a
EAwTw2Xn1cs3262hSJytaqGdrEgmJTVKc4M21rnjDjaTR2zoBBjk9QajxQO1cbAbIy4KNH1mP/pF
WuH1tmWmpDmxtCLICjA14oFQAvR1Q5lhjEFmuDHN9XUYpHGYJ8OlUXILTeKpEmuCndtQptgs/+XZ
B4tyW/XFL//MbqrBYhNE3d2rcVXHacslC5E3wsHO2h6GwVrSP6xa5f2OgHEcBK+hm89Oeyeu9WIO
w3pjaIdUD06r3wNGJckgoGesws6sEMTpujX5gXSuvXfsi0hPDt0UQGlZ3kbV0t1SYtVz3QYHH8R+
MZL1FOfPzG8PD8FHe1Jk7RcSsWNZAkLt1XzGsyMKJhZo7Y7iNnKWwkP0IynRaFa+eJT+4gAICU7I
rHxHcMLc+bxhbdlIPvccUaQTz3MqcnP0QhjRsm6LR0jp7w39E/DW2Ya4eFmlkKZ9xKsX0GCYJs4R
EukD89KxtzlRZvAgBubjAPHkdMFRLegl3FXY+tq+co9E06q4t9HGKieEQi/aEWLWz1X0nqoCAu1Z
rZla+bEcYuh6hwax57olAGKP025RkiJXxcxZ53ERZDaYfXRP5LjjsGnVgNb4F2fbMhevf351UF0k
IX/Zq/dUnfN2Y1YpYmROiFtbKgXAGRDH7zoTCXgVktNx8mx0CvMr0vyFh6aR7ZEQ3XXyQ341gmaB
Cdz8Tk//WKcKdpzE3YmKG+UuzfvMo7/4QKQK8Ozp9TP9UIxTcELTUyPsAsiI1nVXOH6lRBGl6G+U
sxpMbbYFHe0N8ds5/HS8Nxu9gbcnZSJhHQtLM2NdTfy4PPKuE/ujRrHc9MKmF1YLYUP9tWwGQhyD
nT+xhmd4IfhsVA7GfRuVy0w039YLf7v/G+j6a+PWAdvBVwLgZ0QMUzuQzpe9irysPHIi9ZnWSVEY
jYFMlM+OhY1nj+bAmdtW1ljRpWC405+YuePEr2z610ePeXaMwb4YDjpoQTEkw1l1m8CGjqLTgSQX
j48W4YRoTJclxW8sfavnV2+H/+/MI+OYOSp+st9OP/rD7wYtzliYYSgXAmS46To2q03HRrw/Ec0b
g8N6RfCjxHe6YaUu8DNjjQBfcX1+zDCm5EWVtLPua4zDcFco5pldMwRzd3oW0HW4rKKYbUK2ZISs
9aQziipJ0bFLeEixqHUidxMBlgGtkGDSZfDvh3nLU9U7D/6SGHUaK61fcnhNlpvzij2C0IKArF2J
O3lgI4EL1td/DgWGxYF/Wm03AZM5LwgaaQslNdmHHicDIumdJT/mwFFR9Riy6l4SdF4Ju1npJtwY
Wtgp6aMXKQIT9UMYHRu7UqEqQrJcR++IxtHa5uDoHwd078TaX0Qnx0F5kGKowk47LOz/XQu0Izpl
DttjdsTm8jcS/eG5MyCqI2eYIwyMAovr3yrW6mCEHJdjg5TVlUtG+wMOilmE4v5EWo0hwqOyJcp9
fZEXEf+JKe1vNSR6Iz0h4npjBFRTHaDQX69txGlTSHMQr4S1lu96Z+xmmlDR3M1Z9V+FyaxYEU1o
oB6Tmz37HH7SiwcgGnJ4kC2xhl66UUltuOris4QgPItEXdAWefltjjkj0FrASeY9Xj/k18rXo5kh
2ZEiYs+Vcpf/NTkE7sOaD2MlHTHLU3NdvT0oW/g8Ce/BQt3AaAeEyYC5o/Vp8knzuFdnFZrY1Opl
TGKTCuFSo20d/6kLFV04RccSRSiNtzJ+3cMsRoisHbuntQQiRjwRW83y6TXo0jWQGyOQGiwWnQFy
BizPYz3mmaV2T0sGtbhwi8Fu0XWbcG6+nXVWWZEM3MpscIp7yLyIK4VNdTSS58BW07qm04MifEsh
3D06QdN5i5P1WF6uVGLSsmwFNuReA04KHT3O3z/8/e17e9dH6uk8EJaqgCHGFfJDp2voaph4kTUW
4bDJ6dTvHgYEeNDkuM39sMx6C1GsjyMVa3LZL+4AUVBVJLQ/pIJlmkJj95CCSnxvGwsxswY9C4uM
B+ydwavztPxasNRGTryDVVma4/dJbuKPhPJN+8Ype8HxTNJqtUEme9Z0IB13Xg4orTMeFQ0bILDz
32LAjcJy23LHmphQQFckl4ggNEWoCC6rEL/FsJ9vIVvA7uGFBr5NyM1D0UE9WAw4gPATsOn4PF4r
oRWdZQ6pNAP3CGSKXUH3ZJF0COMW64em98H1b+IgTmImz4Km8aCwrBs2AcS9I8+EvGuYfpeo2HEM
XHKZoMVQH5ceP/dGHIGqHpzK+Q2Fhjah9gEJhmCvZEXt3nMR94YGAJ7tok235OD+lGFI1vhi6ZEQ
D5TKSN50d8s/thLhUia0U1s4e24AA1t32hYrKOc5I7IRmkhunZWXMgmjye+X8rufGOM4oS4ylTXg
Tbqsc04zIZ3qDhJ5CdcC6q13cECnSFS8syOgBqZsgbi2oQVmxPteevxrjh1IYs1Bvdv18WCbUFeC
F+/teubVofK+fUHqxsTfIF3O2fTKvN3IZdEtEwmf/7UfhokW6D6AeelL/kH/2G+2D0DumqGSMFWE
FaEQUNk3hmoaMPdQzdaq0zWCURCEsC62l91XkQRpVIpyrPV64rKCzfzv2byYhzeEdNqVik43e0Ps
e5wzNzE4BswEg72Tft8AxQj9G9/w/UjAKG4EqXEEUGs4pha0jMgklDhRuHmTcSCNhqbPl/1uWf9y
j4ozk1ExQlUaGHipUhH5chyWq3rzb+IT6DJqslHCQU1VhKY+xE8prRL0NXviwcAvcdTz/sDxITgv
S2YWt5TyMX5Xxp4FbpHsuiOTTHhF1dbj7Ye66F+K6JH7LX5T0csPMVafCk8XniojaaBIOaG/BMzr
ufY+xJ0yqLRdfy+OncQYQBEfoa4L3Ow/N+2nD833/OCkQPrabRO0o7wlcCae0S8tHR4lUUrBxi+j
VYx6Kf33dqtM+dr9OPk5J1k5Cnh9hZKoXaMkmTFmAE2imC57ZRAOsOoj+aOix392/EGD3YZCAHUd
zBEpOFhkIPtXYKJ8uwwJ9Dfhsjs6IEiT7i9VW4pl2illeFxsYSVrl49ZeJgOJOoTkdgnWomqul/5
gOpoQONFogH5s87q3bryRr8O79iPpCKhYHujMLb9AKH5K25q8ARaiD0ZxBiOwpq1fUjAB9UYUiZE
2jprpwgaIp/Kebq2QB50GS/KH3NFiH+uCbitCw7vZAHxBD36X/pDY7AVahbapcpO6Ki0TdXq4/bf
sHHlslDcVtTVrsnEcS1d3K8EqcEic8erzrt62sNevSslKssyYuiGnro6YQeBvDkJOslkxB7sPu+I
1Ee1n+bFah9D4KSKebh3eg46SylmkvlovdbtzoButmtM3BwStWYO/ls1GWiMO5D7dpti77mdLMHy
6oV62bI+KtsMPAoTRj6GPHMYnLliCdC+0Zul38jz7sX7g0f0bEjjM5lKxZn4Co15X3bKeT4PkGjI
44394WYYWvRo5UiUcseBWzYzuIWMsWomH77kM3lejpZ1Njun2klgZSaOKD68zH+IU1u3puMcAdgj
QJgpIzCVVKSDRRGCPzX9mIluzLP73QjGY+AUm06ISC3/MGND48rl6f2KLFZV/LMzJoOaJuGqEqBH
HGfrlobbjnKYOhckUNeaFLJxXD4WSc8cs8jpdpzjXa/FMQ20lYcKEF2Iqxp9vY2HtjqCuJD4nHKc
4q6fpqOvZIZlJl5W6K82UOBaFX173DS6SD74stqp0Qejon6a8cMNflWj6ZDVPJmeYbbsqr+wD42Q
NJ5Y6+iBE2w+mA07vXVD2ADCztOw8IgXo1J/VMkdsHzrdwa+Pb2P0kfOzqSaWPzsT7YElYJc/Wpd
CMhc0b2QZV4eORgh4RpW45w50akdrK4JUry7od4ImX9HabLz3BoIqxns0cQcnGOP68uyWtC98Vpq
IFKOW8NyHe+3HV2VBf5tA0ojarzNaDSBUa4hnPyw+b3ZEwT/6gkfiBz95JNZaAt5aNaNTKY8sNJl
8RiLpuhQL2tOkZYLvqCvfpQ3xzyA/GP16w0+g5hbzA81p3MsXKUw/KJpUIm6vPzmfm92QQIvnVQJ
hsmuhKk9YC8UZH4ywGNX7yNdEIXDHKY+h2/r/FmPH1M+qU5ir0381gBvZz7q+1ku85yrdFdxMlRl
EzMNt4plQgWpIB7zr0qhWAWKj4IqZfVQCG8Csg7zu9rGnhaw+2BXlLaNpRFB+8c/1ZB836Rwf2Sf
9WoU1mtHrCc1FVIzIU2KjC3RNIPD6vpbiI3nVfBxEI3SLmyeEEblaQIMZexEjOQ7QdNeBxDcTEGv
wNDeK+l4Bgd2iIjNRi40ogVSzOmkvKK87VUG9YTctLNNYjV8sPBruz/Cv8owFZsVtzLncS3I9+p3
fOkxy44tHRelfj+W2PIHA0qlB4pMnPvkacpC7Uf3GR2fyyK7cyKI2A356b4BjBlsarygezxFlwtb
Yf3TdUfrTVfh5iC0azZA4BqV3d1uGnyIUUnmyLPTY1+NLc2ezNC08CSWnfe4IIodLYcm2xyjFxnf
FeUOfjJPeAqtWB2AY59yazR4MAmjt/fIodUNDuYRm9oLojiSs/n7aotYW03MWcIwEh1XlW5orQw5
gPUacnxGRfr3OGVEWBSUAIiqU/mFDVhOhG1tdoxvf/S67PCEUnxFuOl3ytghNdrDuj3ilExAewTC
cR/4V5YVFO7AGaCOQUsDucgRN01j9cc987t/I0kW07SDwLQmPR+wg2jFdAsg+LP+4riWbUPXIZL2
chswq5ch6McThHHoGSxEtmjuITweiU2nCj49t3Vv2SA5tz9mGqqNc8fonydqKAu6aZjkezsAi0C8
o1sTK+jra+ElhJ3msZyTiFQcdJVpnc3wqhH036fUQvtlAGTw9xOt9JPb+Hw3TseeLdhPTvC5IbQz
4ZaoXgr3ofgyqZwancKSFuTPzVCHZOrqoKupuaMjgnQ5pHO7tt+NlJ+iYXmRv0u61cCyrMy+Pr7g
b6GoKANEESBXpI5xarXjkLScSrjMjSC55MYyWsQ4pA75W3Z6z/fNm0Kc20FdN4kAr14Fep4/B6CY
Xwtgvel8oPtevBqdPOmPGgDJzyfm8JRAVlWX6Ptg26ztOjE59sWY8cLhjNsuVe2duYYdIWFiS06m
exw+bddKjGqG02fqgw4iwz3Wp8HD0VIaxK5kOimOzig5Jso35IGeXLd7sOJO9czkh1mA7B42MtuC
1Yt3/V9ycU4evqVFoGslsllWLekgpku47Q8wmcbgTaSIWEEjknPIariqngQQiUyzqOSAW650F21e
aC/4GY3lj439h9mbo2Yhvzghj0yLb0OyKkodmvpzDGdqFZb7ha347Il40YBqBsgsyCRY6Yg8QUQL
EFsIliZEiMuUDxIdSQjCYT7F/TlVOHepeKCslHMgH06sxTU8FJ+yu+cFczQ//UcDoJ+ouwAqgC9d
peWAx35N3neINWxpIuOwdn5FNfM7kya9N6kZcuwOOjoP68TjeHxaOit1rpR9OI+3s6GVfZ0VKWJq
pPeuKOjEiyidJK+Uk2Kkuo0fz8ielfedZ7auCoqbPW/8HpIrLVBcu1+ORgd+Ok0lV93qqIWqb0TJ
6mZ7xuwTE+LHtjkpvPJUwjRFCfhMvKZ26zR2nBlfCKYl1UCHscRoOgG1DP6MDqst+G/NfrsnwPsA
Ks83KVuQhivcXwv5CxiMcyQHkjMtxIh3cYc1Ag3Wzsyhny9tng8SduSRHImdI1tyZIkADF0lkMfJ
SHU9AReq9EXf2wYWw1XDGOKurhMJ5C9OXfY0EqUcGukLvcfEH2Yoq41SD4wdbcaheWp0bpC/4Wh/
9OPctmGt3wv/9O0aaPtaHjJwzrenZ30TmrVWtvhVEDGUzHI4ix9iI+6iNAa3fRpWPvivfH0qce+q
o1qAAWFSJSnfDrvHhbizcoMX4nejp7OXrwCXENks9r/Pc2OAilUVHU/tj+tumHoURNu5qrLqLoal
ZKWDvZ+cEeAdNqhQRCdW5lYlKaYQ5y5lTysDAawAd3lWLhBzQWOOVNJn/Rh/tUULOLyBheywHg67
gla+oCjnLHtf2P57cecF2Zx+k3bfN+mQ2P2PfMF+C+rN4D8slDtW37lWp4y9ZnMNRjvRUKcjQq36
Q9gZFtE4Uskys3Yebb1AqALCCLgy/t/GaDEBF9qOBWgvmrnts+l8GeCSHIW3NDRvW7OkbvCryBTe
1bAxVehrXNXWfm5aLMGhF1QaOlGqNVVIyyNvQ3nCE+MMPS0wwvlvK2UC4PN4MczsoTyKWxKNtLhz
kFkBrWZ+RXdJAXnyPT+b72lLk2Aicgs8VXT8L81jDjn0gdlQKd5oTFHQ05QCXYubzCz9x7wGrBUu
FtpPl/zijrSpdSHfOcfC0pPD76IDEbaRNk97Bwo0+oHU8uPj5wKJfpZ5mOXB8Aw/PDwKLcLXkPVQ
/R8/i0qMyyyiPq90Ss+DzBnMyTrcte0DFXpSv43T07Tr7Y2VGLRNo1dfX2Y0/Gwk+LEDQxvljBcG
bN38BG6U9SLa1NzffD3JIrJBTJiCUXkquPMEc48GSn1Q8Zbn5BM9EkA1PXpstKrnHz14R+9PQsr6
nHOQea/WsbRiOJNpSurH/03RE28ZIJ/0Yv4kcKgW0O2lCwhYEm3KRq3kQlYTMdHIPp7mJPZ5/v2f
ODCkTDxAoWLRPvgQ+WAZ5DsByGwBUDs4wRM9iPcf/WU+3pIMpS45y999BrLkqZO4jydFAZs3hSa3
1w9WuUSLb9mNZj99V+8gRlVEeJ0LTQhroMMdInB1cKqLNjnHcIFOVFxLJ2jSudLggCH9w7W/D/9J
F0VZNBrmAJX0UPvy8n1PshqlX/RPTrbSeOz7unaZHkgzK1SSHd2A45SYq8h+zl87HBRxExSGh5yt
7MVq0s/EBYbUIv2lKDTHplUoeVn+F/K6KzDj1OAKrC2wLvh8qyosAZSngzbKZE8TWz9nmTr8BdMI
sIIxp2FQioIc9FEmANytZkdBurBDTcd4eor5WZqGEYY621kFwe+OF0wa300B9wCSapAQtA9bVQI4
/Gf1d6ix9pMpxQ2nZPp+DgZMUi0GFED5rLiILwrlhGfRvGvpMThNorHTQvv7NahKYyjQ8QQlyTr3
Nl+utAjRJGJCGphNO8zuUWz9zBOjFuwUgI1LrZjyfgI3078yAPjsyG1xPNVpwDrk9hD1chNg297B
QYOzFQ29YIcVgGG/DsPvTazRO/UZfBf/ERGL1VSD4EprhYF2TW0GscR/GeaSWnX/QBg9oieEeUAA
bBAfaVCoev3Gpt1qy/MTBNxg5B3RHLlyWm+ytgVSVteprIxvguMIbyk+qSiZwfAQ7Sv8oyp0K1vQ
l8qot788iGrpeGyeOnMyC0nBM6ziHMcatFLbRbouWH+PBkCWgpNopCwZRG7/ZYTED1DQs2SW0sDV
/GdKSUJFc1yI1CbknHzYoVNICbQdvgS3fGL+4fqTcGi2/pkqzdxzZY8+Rc2eADa6Y7DuD4vUQwtL
oHjvCdseiDfoB1AArYk7qVH0tAFmLLkewG1C6uP8yejyiPDvQ5oncpFUTNjV43CZrKNlCP5PFq02
k28HeTkqXQJHYW4UDEk4wu+XsYq1zHUAjPsIB4EFZ8rWr2CEB3+5FtnsiOs+tFF2Q0/wVb6+Ejxq
PEcFXJCidDkQD+esylGQNaeR9rdvGSbTC+8EOcgyU33Lxh9cCb0LglzYN+jX/z7+G9GYT7G+acV0
MhAnqNmsbi4zQQvhlhMHVcdnBdWfIbIqjdNA3z0EeD0tq8+ZA+4GUIYtLKpvyGTUyrD+WJiUg6Y+
8dBWpOUvPoR5Q13Vx7HsPlwsoonAdQGwcqvHsiGVX9DZRuRZ46JB/c/OL98grveH5ju205DlYhkz
RrljWWofGtTFWNP9xJClkX8BbwVTuH00ZefjgPrJkqu9lD20rVMoVgHWwynvUXJlX/GaFwUhKiOZ
ZfmZxU+1Jt7ntPxZ8pR6Ak4cP8DENfO3p98vmWuLvXPTEEFnID9IWzf5jnItR6Mzgr+3T+b7DiVQ
mAMijjTlHsplb4+qbtbGIfP+QlCzdqS8iukbqNxCbcRK2f83xqgwjEJ41bWL8S+kLQGt9e6Ao9k/
azEEp3tnTsLGPZLaMz9n1UuAJag6uNMtelNtcUfW208NR+WELfGc9cpy0dKqyeYPXHYDEnISFLX6
OEjRdzO5Bjw30w9rmXloDovJsTw+MbGF8ETy441dUCDEXfSbGBYsSrymZGB4ZxNXY5QYEJhPNv/U
YLdpQvgnepWtxID68wi4pNUOltM/mU4liquDpR0/GXEY1nGSsgkjSAJdf9p1tNkdNLJaDuY/IXwO
+Ro6N2gBvsWokvZQIba2U7wqvbuaTp4/8ysC/lkIzcpdSKXiP6Yz0VA+nzvuxmkf2sryJ3GK8oez
KUOyTbuGHruZfCmBDHE39ehG/JkiEAWx9rwFr04kAGJuDOK8NvOnC9rUmIj6NkE5xs6OPKuky4t0
ZWBkTk1lsyi+E3TFUiiDXt2cMB9VfmmCxvgfRQubyNjlZznKtS8XrsLpVfCmsKcoqkNVnkXnWZzI
pfPXaVE9+4KK6Jn0seE2RX62ep9jBteltIIrRcp8gDpXTWR/Tpf+iS/iP5cM/KVAtOQyGdXlUmAR
7efV04/TLUGvwQ9yeSA3U5UAGHg4zz95gnIkPHXgFM4YVXCHlgeSJgrGnB3KTeBgtabvmQBWH7Bc
Bq/DlLQOFbJCV/hN0rLEafK8VuaEH/zq+Y5Oes9ToI7uYBdjV960f21lW1NwN/TQH3WiXJKEdC8O
ZJiAl+hXkqCPZdPcH2HSqCJPKw38viAOBzsjinz7Tpc1ZLWdGmfIwHzFhbHbw+s9fj+s7fWwxcNw
umuJhvQFctxxek7Qh+VzNtcLoUw9WIT2HokmSz1un0yczqjhEF0cm39/1oCNNtVepSao52NbHAd2
IgpTsVP2l2OioCqEUMoWYRAvBW3Cb0PDNkfapNXtU4fQIRTjHEhDN+gb1IHr//TM1YxLUokFUnbt
MtgAAea1HJSaPPel9laMPrhlqTFQTC6F1h6q1PyirNVFqNZLoe6d9MZmhSRTf7x/ashu2o6U0Nml
xWaN0gnDbjSJm1LFQuXjEZdfwYXlNbLy9RIulMWPl/KIg9VhGd77zUTxp6gjoHJZNzxqKpk1BcF/
ur918sYrJKN/NAmDcYUtRRjH/DRk3R0uaK9PAIjNUNLEzbaidSCnLlMVS0N+jGS1KaTmyxpWuAtO
6oWPVJFkdYgc3im9o0KoTI6eb21jQh4OgNvElEkBWmLh1l6TwAijlsfEMnRWFH6v7cmVx0u6cxIq
JFxjW7rgGneWhXlPyUDHLzWoiCwsSFtzNZ78p5NgntJwmIPn6CzusigvNIviyhKLlhUxzYkLfnw8
VoAWmbp3YLttS7zOSXGjnLWA+FsQ2QqvLJUZe89JGTjRdvBMGKi8qyEUXNoB46SCBu1dFHLqzG12
SRmCerS9LEDdn1TIxpkHVQvk4MHRv9YFmkVUja2minEazOjf850hoNd2jL9+jmgx606bQH0KOuim
vG3Ls4VuC7acYpMF/hF5LsGKdZyb7+RjU18juf4rWZjghp2dchVKPuDXkYwO6BpgLS2pkfn8H0vU
5MXn1wIFBD/9h8t6Kn0b0kUjK/pJHixg4he0Mj/0nMkN45qReGefLJyUyG69sv4qpP2J3ZoF0jwl
QUimtPBsZE0l/WYL1NBOWnzTAzThtVpgxRMAf2EpSz+5YmMP1ZQBxfXHDNJno8hr/7PzXQVnmi38
U+XdzNU1X+6tfjNacrAPgCNQN22DX6UL/PlfK963Rc3I5a7Y45CHhnFsr7ta8QqALZ74dSGuLpds
HTeJldmS6XiQG62tL79ZhlAa4uAavKxUYur6ButgxnMo9ixkREEBITNLyA6xeRKjP2uVLfZy0hWW
42uw5IiwtksCpBcKBLHTRmEyxQs1HS4u3bAa3Eu2Z6MV4nZ2RbtIHYDzG18QkVuJfNrGf71x1zuz
KY0sUeRY/Q+d90LZSLVZp4v2qQJw52TkZiy262vXdqFzWui/4oAf0ONZIrsaEzv/OF7nYT4SqWvu
cA7QMamdIiaYpirQxx7nMBTcqhNtnuaSAWFmmsRVH5uU8isots+50h+0Lkmlz9QPwhTB2HgOY6Ao
U/fapsQGUzXIsuPvamPt9RknDogSv11I4Zl1eXSQeR6khPnAFMeB6DQCdV1brawymsJIk4lykhzv
wZvmv6n4kgfAGe8ftm7E20vWpUYFM95hDKtNgUnFJAZwv2EO5frFSSk1d7OL0Z+Zo34VrfuMocP5
11NcRmlZkqoDmAKHZTUmjBNbR3CRJPlX4YfBN42DA8vDfOZ1XZo743c11ysbjuYshMAilHbReW1B
iy2YGHpqgkTXuP9kWVPH6FHauLgnBYCMI5KiAG+OegsGZkm7Ub/zJHzJNdW8krdl7KEC91xkI4zU
UBDE7sMKNcUcXXEvlCrfAfiofH0nnYNqO6uPihhfMr7QMryBLvO2IqhiIP3vkcFOQJi8gDZxkQVf
2MPbTNy6XjhQKtVGidSxaW5HrrXs0jvaPJmVKWYmeMejs8K5XsU6UlmlYegavvYye+47nilT36hl
HX0A7rBGygxdo03kpxi0j/dZiM/Zht2c/tylS5PBGmIFFrkXMtDtJcTC0FZ07Rfk9O1qHhkwWm6V
IFk/ZQLLwStmcwbrhsnqGzpHJARDcs5CplxlmKvyLhnzQ779uXZH7PxIlsNptexEbqnhygurHgbx
cPZgglNPIPSVBhofvMAN1m2buTqRphk9lzUgoMw52vsWAWlMyB3od+tcwlyVf/aww8SLbCZWmFlD
SwtGZHVBHVULX9WSSTbF68I3RjwiVmnNrx5gbJ44gCNqr82vHC9rVa7FkXAkzblM+7Dhq4m0mMYg
wLzc8YFdRbtmEVX5zeLd6+4hoEbTLHEAzQX5Ho/jcB/AAWhNcss1awzT+DZ38joNL/DiYNFL0o8e
/jJzVjwJW/OXNRD8ia0HSOEvl0YyaorqKcu8N38Pe/zuAQnUMw7DK+GnbJzh8VuZXt8BKsGOk63v
e/EsLOkVFXV5ahwHMxQJIpbTP/5uaiqPUlrl2nxRNjgcqd7GckefowxFQoSLGp85x1vPWPZYCX2Y
zf7f8l87W9xFwMyYM232UNVTA+OwgAupP6kPOV44AToDY9yVElrEBL0rMz9UHSlAUomMrl8F3kjv
2MBxMvtzKbfuMdzpGwYirsKcflPxNP7nsV8WQPPUq6RoysQ1nSbAH8BrnL1f68qaCZCAUBz7E1Ad
Ah18O3yN2k/OBEIY61Gu2ezidXyU6/AdtgKgq5dHcv1ddrDZNynP/lRJP2w965BCeSdDajYAZgLr
IS33gYhkXLzb1NrXbl2n5Cj6L2cy9BeTSBoAp5hb4+pxKDjs/QGXGL4Vxal0Wmp9Y36RcdADPEhW
D+9+M6Z2ug09msuOWHMYrBL9FGUYDFOiv3mVAri00Nt9ft+n+NDJlO09OKFvKEQXLRtSr8dDC0h6
NQdbyPSPti+BSF9Z58ZnT0OtwVjEbifW5XOZ9gw0hqECSHhpimmXOyY9B5+Qnj5U8RZpatIViVlg
GCAcWc86nyZtx3OVhcAVSmLidB0VcDNsML9sascovqyRGm19IZjtZl42tz/P0zQtLkeJZvCl+E7Q
MeK576nOjzeeWqgUJnv+KaOJuUiO6oFjLfSmmuBrTBYC//rbVhD91q0wScW7FrsZApQ2HLCGruWf
MA3zgflydzQh/BcD6Vd14E28gFk4WfEq018furw09dGbgay3bjxza0TeiDVfgaaiqptCJ+qN6KvR
VPsd1PCra0RceIPb43ARLfTX1YzFrixggRd4kJPCxMKixKcjWylcyTDHnickwqP7V2YXl+D/frRa
hBWzVR0Xehk2qx+q5mW3qgiT62RAIq6T2foeCzneqJq8IamEvgVtIYg3Ej+QcRnKozYH/vouKuZU
wNtz+m//21zszDUO0utOwV/FIrabNH+RHPfq8SNI1vSRohmMso+o71stc1bBdQSitAZuQ6k7Jrlf
pYBB9c7j4LAwrwqHU2kB2OFA7AyBrsnsgMWZ8Mcxu2OcvAv8+/c/q6hpHnyr14sKvdZJEGDRivsf
9fiqe55Ix6EQZo4HHoYY/06a+VY6xkeowbx4am/Fci4rJNlMKjPA+UhH4ckSBEXxwehQVME5ZRJ+
NQyI/HqK5b4sVTlTWgwMOnjmF7+oN75+eEjqvtHLyV8T62FxogVMi2ch2/9SHg8THoziFb0Ddgre
n5eRw4nKaawWwWCIlcEmKwhTOOjg3stjiPpHLnTNjujuaaEO5y+0nPkHG5USCKOch5YdtGuc10Me
mtd7KinaydnrkmznUVYt0tsnXkTNtsih7MAqKVe7Hnvw4ic664BKNB17txqGZVYbFJb8JRNmtPIc
JE5TmRdCEJavZmETgQr6awJJCrr5ES0gtT3k/OcTOVSWILM4FV+WLxtQyEGVUoPcgEgKqACL51yh
u509qMMNbTGsVumtoCuCOqAlzqslN2pAosCbbGsV3LUxgDDLOjoib33i1kxO5O4s98l4rKg6T6AH
KpEJSjlHivqPeDwPtUixJef3hpKkOrbbTqgJdQDMDj9iznSeX9d7C2NRUwzqF41XX8dLlwXGal4R
Em4iYU6GQlgmKS8xA0U7/n6+qdClL+uDWea79PKQEs4uOaIr2lOsRpO74jEtljaZYIUWKy+YXBlC
pyT69ovxH9NATa8+7ZSv0mRh2Flr1PlRXvsimzbpPW3Le44QZJZZ5fq+5j1UpEeF9EMnvYTZLjrL
5zATtLx4xVHaxijAU2T7KKZUoH0PiZ63xnxw4FQabQFmNbhRMf9RIaPzeV2ZhaFIqvIFLZB46Lz1
qXQNSmlA5+Acu0iyrrAsF3oN/alTn9AMlWkunbtLAk7BIx08IVT9L+aYyVjA0NSk/h+CPu+oziM9
1KATVnoWKup56a4dvtVSmCVEG0+AUQ+G0CIRzEcJpi9mZTLLnfeD8w7pNozNDxwRsrGKAtBPDc30
fS/IaO/7Qk3Jaz1o30KRASMvv56O7H2TegG2oY31K0kOzgMxX9wohSZdFGAPYMxsR058CicCpszb
fG7/eh2BZ5Tru3gmBKmpAS27koNbR7TIrpoJcbZFnXpVcpVvAsvjf9ZPopvmvfH7kWyalSaQYg0S
Vqn/zJT++KxYeosMMa0GPCIHn3DNrsYOAXbKPrlD7FpYlKiAtBLkPOSIscu33VZy67BHhI7NkexF
iNWuazewFMvqCK0qUFFaRUNOx3GO7BCGsUTQseJrz0seNwNeMDh9RWXwKKjBvoPvGAotxy4oXW5o
FWptm/vbOA9e1hhFzxK7uLMj6Wp64anc/9a4UKpW/C8irssfCy5I1oTrrN9132CeijeAvv4FBeVn
UefvyrwrJFP4nov3rVozfZzJ6BYZ6GUJRl5dPnd0S7thHudCK3eboe9BB6UUyxosEvI8ryyCZzN7
CXF+nGj8+mbJlkXgwKm81qzK/yiUXeDoYM+H//XysAifrzGAI4Qz7E6e815EA4s/E0gFri/bRhRS
5gDRw5ztGdDM9AMvuUnou0UDx8F6U4jgFOZdmgfsSns+BWMHlJsaV7fNUZshWDA73v/wdDMbHkFa
eAuIeBy/z6hhhi5FfDb8DBs4VT/CUO1ItqJBDU0id54kx0wfWx1BizLO3vvQ0CAGuQcIjCLWO7HM
LcgGhFWuqZ3jFWeVRwv3Veq0/n7Zv20zzMSCPX8h3NqlsMjjbM9mudXjslUEmRio7mqETULE5aio
NlISF1bwInI8kb6HhKXbQ2Jek0NA6ZKmCilZ//B48sMz30eeCiGUhroNTrXiVFJnXda3LmrJXSzo
b72K9wuXMbJ1vBQt6oaJ2e/0WucI+9GS9XNcQDg48cXc17vmtm7l1kUeZY5iloo9HO2u0NP+KGCI
Sdip/mwOFuiUvfrzxtiJkFnjXWNVJkB54d2jD7CGhrqUm+uuICaQNr+REewRbSD1f2z/9t81TTY6
PTKReZCMtxa4YvzTeK/ZIdY0SHqajjHNxEruUlpQD84ZjPgJ2uD0iu+zHSCW5rmJoykW/xnkLEYB
+uNHPINa868gL1hc8a5rlKiZBJa1lv9nCGLTZ13r0dogVLK0RvwrLa2YGnPXESN97tzGTlVxXLfF
eAMG2JIdvrCxndTaK15JUW64hLYlWwruFceDSDZEll9A5lQ/fX6mZ4pyiLqoPEpcvmp9ztFdAcxW
/Ig9NynvcDYI0oAAYv/+7UlvZijSqSQ9TdX95RVTijy7dLbTBDcGHoSa2Bljps3Ke1qf8g51kHSS
xY9efSYvhzzX4hxzyrJ9LlsdejvIB6X2GO6OygJ1cmLzykq9oh6L8+8P9HFH7GJaauP2rp+anXTp
vJTOwYdS+r59eEH/Gns4vqI+v+WDRKJR+20OeGwXAVl4IviTege6SUqihdWYQOG1/KQLuudiJTwz
Od0apwh63xClWfJe83GCvyNNs9PajaFI+ky1wDbkl1q53Lg4u5DVQnwK5v+5g98HYXhcuD9c40wj
NTbHJCy8ZpS0Zt1QEbVcdpnrsDKYYkxzETNdRwjn6mJ4EsXdney4IflrHSjGT1JitrOndruIXnF9
mYETbEw9BZPjpVs1eBIeWk6lujKIRmD9cjcedhHpx/fFSV4Iw8tLepyyqpBHgrx33oiNEF0yrbZn
Sa8+uzsgLpTc/HBddrtFN+qPU7T87rWBkqn5msVdHZ0hVS8sgdvXYjkNHDT6frzqEerv3ZqgbndR
+w/yNtvqPdtoXI+RQ/KDkmlIJx80C2QJkQfxDGkWu7fQk4JrEzVIsz3yi54RmTfsZky5jcS5LZ3T
aYiZhDAuzJKfKkDPuBszbfGS0zhHINNlasmlXvJ4fgba6MDihhg0P6+dpBt7FEt/MP6dn8Rkdstq
pNN+T1vTzQIPsmEXR8qKBIUVKuAlk7eKVemGT1Scfz/yh39+9R7cJWGwQp78FLdsX2BkTYCjSfaP
dn2S0iCBgvQIO/yO61Y+dXltQ3SU7QEyS2ko8EPX96L2ZN5EqEIv8KyEC/cFp7a9EmnHkDao4ruT
cq8f87TZ2Z380FC3LIjr/FtMpYb7FrxkW6NRPEvhECwbXAuBfj7pPf+PebLpA+y1mRwajeNHbePv
9Nxivr+5Zo3ueSQPhHiMWpG0qXiUxgf3QR4Y9umITj9APopCvMQxidMnaDAEXCXGLgCXkKSQPzXM
AQRlNCYAt5aln5UZ+2EVkOe6L+cuSbYR5Z+Iw3flynHgcCaFnv1XHbhDctmMAqltc1gIqWvl6hYG
0e6lR+B9oQchwyfiFPgbVMssUJodR9U3Mn6GTcny987/7ZptFLV/UEUrC/m12iqL3DR5JZ7mjht2
6Gf4JvdC2w9PXl1piYCcPE7ZWA836J95ImaVSaHYtJWOuWux1RXJfYHRpwq7adqL2wkOc4p8QrYu
Y6Ef8+UUy35nLIcQk+zs7YLM2/wh4o34tYBIwL1gw0qDWfvyieobtehs9nBuKsu7JOznGNtcYKzy
akZOSjVl12lYeuY4++ACX/2r4V/7629cdEwdUAkfBN9mDrnumSgEvKKIpcTpJSPk1HN6esWJDGzF
66ViZGQDAGiZc+AouajtmuVUTcLpYpxnZCsSM/GIILAXChbP+0UWbn1/SW+CKFjt1rRQa0RVybO+
uPsPLzryjZX47CX7c3ZpCZYR1SzVP776I8sPwEvBQVJay3++R01fm2cik1jV1bzOPBWulSNfgnJf
2dXkaOfDF3EXdgZkvXE6iMCQfNylaVFYkmlFXOpIz0DyUz7bbhLWa5EC0NuZohH7kSvKZXuV/roW
I+63UU3yEuSsJeB04ev2WOXAYttGmx05MGWzzaEdy/6oRmpbyr4cfTxHM3mbLNoAwGBCOKXOHRQU
V83hEi1c3v75b3jfCq6A1NQjzNT+o+OOp+BME0vEvBoPrUSVcv4AbyqG7bnxgHNepwNKx3xisF42
t7P+o/QNFMwfTALMTSDqg3NnUsXl8Oaw/3jR05BIfTCvGFR4v6+/qn46HUsewh2QD23WNOa/D809
cgUTe47ErnoQJFb0W35UL7IchZoJ/D/2GRG/TBefgzcJukHlUub/5XljEzaeWq9AogKRL2et79AW
zB8iHmz8Y7rkLojg5XConrhVioijX4cbAyV0KHc8vx0K7xBO0Ds8hfJB6E+OFbKHYfSJpMfCeBUR
a0Qykb4+oBI2Z8Phc2iNsDYU3MBYe66KNJYULz3tE7uS+u4vLJANhPzfipm36O+mDfrp37U+l5vQ
vucZ/vgp8eDq8Ko9jBrUR8nwCl3GgbFQeh/JbIQBjoUsozpxz8vqMdBbdbhNVyEvaNn4jjcd6iik
iWTnS75op1aIMCOXtA9ZQ+TcZC/eRyQtuBPXF3q152B0WlBMK0cqL8gO+ZX4aTcW9YbCKxJ718+R
Mj577A2z220FF5/UHpmkWY/2hcOvXtogAg9pxxy5e3F3f82yKBBfR5zgl4R65kW+6dtTLACsj9/R
K5AZFYoUnoHeOP7mJB00vmnQBNPQNOHNGQCPDdUmgCgd46TJ6vzn/+68Ma/ieiEbuAGqjsCkkxf4
MGUepGmOddyifE3ExmlraDEjrgRl1CMFNtbAVKq0BkWj3S3uo/9Oar4igOEMYXTHWQ00+C7dCUcW
CRJ9YNco2IRuSSQxQ+9XGUPBk9k3G/1HNJp/lD5rc7jni7gk3dUAoEe7vZCSjWfrO6qUg96GbuBo
mnWN4dCuMNS70n4WJ2IQRNuuRv7P96J0srKPYIEnpqrb6pBwwsaAjH2Sd8dBzz7qqZzEL/oHUEek
fPk87zvG3gjx1BglSCYJ1ryoN8sCKePfH5EDadpDNxaVVbMuxtm7y6fC2R62xSDfcM2oWCh6JZaX
FFiehVZslYtK22Unc87zSAccb6vXI4XKIuFwg64BIzDG9X/Nu9TIzQMJIJjJYFfq1AdGUkt56sNi
hhyr9OwP6OTGgtV/nohaamqKht/g8YfqFO6xOPub1koNChF++frOv1zhmL0XV1lB5xods1+ZMr7Y
PNv+12veTRcKTVkGxAKWnvuQ+UGVNLDBEnqbQDNfH56Wr7OWInJ4GPNhSIMs+4eCsYEzMN09JRgF
sU2xJJYeWBn+md2gx4XpW5/GpuktkC9pzgMAa2FPNf9E/rm7ibbJkad1UNx21HMuqf7NI7XolcKE
l1NSc3woZiU1xoZVdJA2NDcXChApDlxp5x/GD1Rpwwq/GhjBKvegegD79t52PjcG0gSV9CUWzTY0
tXu2gyzASq2rKE7GaqSksrN/M2YxZx1EL/XAw3HMmlO2PTAOabjOOctVUTz8gYin36nGRRTb69Ky
wx0cLa3zo5FvMqb7o6Xas2WIY/l+HyqcQjXIqL6vVLSZezkozp/MzLsW9AcDd+zfjlJqh6BIkr4E
4jT/caGwHQDrC45E4d8usgLkjzogUxvPTJJ/s1mtyw7S+rHt/p5++pbJ79rPaFkuCJzdP58pkZDq
xBCoBhrB7ogb+6Vpq/IdNo8yEPYcsU0TlukfUciRah/+4tzuQ0ZKwfP74iKcqWEdS2PU5Qbf4PJe
UBPsBliuBq/Vsdiz24sgzCegiS6oZAmtAlee35X/uBgwFHkPWR0YuNdIO+7m8rNCSkGX7HxHC5+L
8F7Jt535wPMxmU3qQPC1YhvLbmD3X3cSDOGiuOOrlB6wa+vHQiO/Zm5uYjzLdhijTAosBX4BRE83
VqvPh7JKOY6Q3i99lE3hhAsu0eNHDWZ/FzvF9lvBA2uTREVuGB9txPlvXvtcUsbZiYZs5jPX/TRD
gPi+b9PIM662JDkGnIyEAqPMI10Ezo+Vz27ABHztjdLFv++DhtdXAngcisZQRm4YYOM62wp64SAO
1NHFyV3smSphMJrCIDEkbHL2crE01VFS47qr/mtzxmv8WsGBjuQD2/i2thOKyDQStffpl1xqgPp/
hD+Q7kEHYhIEKYWT+JwN7Kyju14E+Xscd7fU+lSg2ejQtVezk6KWm0mb0Efe5VnImuleULD74TCe
pSH1PNQ2ZbK/deyGMgs3HW5A9/ZrMzJxv0ew/O/0ixJytxBrve/SlrI7Qjd2ZZvVYBKKoAFyIcbe
O8B/xcJ3/Onx/0N8yYHXTD5WSKFCdrEFsQNKKwujcU2SKUrsQ/LZpLn31G7ib5UculkEhN3DeiNn
wA03wWqXCdyGt7UxjuBp0WJhmzTGUbtt/I9S+CyXR1ly21OYR5Ey8+0Xqo0nduGNymDQtK4q69ra
bnqosdbabizNZQVLOxSUV+jxv34REYnp99yuESViMdVyUY6AS0H4KSq4ag/6Q7r3UR7Rna40otCf
7wsSOIL8zwbmrux03HdUur5fTShUNywLB0h/7F7VevplbclPxt4lqcgZGHYei444UszCguY+NVRG
uXMt90Ou32I9rCV8VAbxyZJudwLDHvGjoF6es1z9sOAUnCchNiEIwa7Qa2lT5nh9vDAhlu+kS4E+
8MHElKr+hbAblgFiT3oTkh05ONpb8ys/JupgWugRfTuLsfSkTRy4gDb1pvTGAOu3iVPnZhtUrXh+
QdMDlXBe2/XiUwrPiiEnVus2whbordQwxl8XKzm75PZHIgZ00ZnVWv2kT46HdPVJRCcP+9L9xvJE
zFEoF5iK8U4KDRjIkOANAjVya1ZFO76Et4aOFHC0OutfAn+IR5/L5JmBVEUgtUpgaAKLH1jGfUBf
CXLeWZrzK/iRst6PqR8GMt3Zcmt/FvYTFiLmzZmcTO/ofBJsk3agu14S1GwDWb5a13E58DTgkKYe
IP/XOTh9VqcZ+lmK0DEPJHHtEknuvvVLmtubav82yZ+7nfyVnyrzG8nLMXiUFtBorfcermzaeJtd
5p/T07QQd4vXaRWtCT4iIWFoNw6UC5Lszok75AUVlKmcNs3lgNQzryqwLWp0nDr6cea7gtSF3Rza
lXxlBwsY8k7UOxJRmaksKV0o+yprA3Li7K9OunjZTbg8bs4cm3rM1DoJ2NyU1f+xkIMPEidxXvfr
SBW1SQ+FHEnZQDOHbTOefMQY02F/NnDcukRD/ENmRdoglrICgwcErq6R8AGLyEcTHEwnQMB+tnrl
3nZaJRPw3laRqANS9K0XTUkZACo3Nl7ALJ/qV2WzaqsTbGf6Xwq0+4f6sTaib092w0qtE9D4w+FA
NSHvGiPS9gc1NyPct6oT4yPIGEtnBEbzCKnWWeaH811n5oAtUC4a+TCK2ZhdtUVFVVhMzUFsHsSL
SnjL8SLeC/u8UOVXZMqktw1LqfIofN/DoOq2NEQBurS1g/aUqV7cWSGRWWNoa6+blTuwW6hNeOhb
2xzGYVRFq7qzug4JDIGSH2w4RTaoSLF3FUS41N0UgGzeSNtkOOirONv4WQtiC7occRcDst1nrwNl
FvUDbrF06+Ro07UOsIoBco5O5zaG1RQhxiuPWK/0RE3lTdXzZXoWGoAun9qS0E3soOKRYTIQonrG
Kq20OClty44YT43909oSJoNthcoaWgGf8OxRMN+ao85Ll3ShXCi0wTO1EeJuA8pN1FFuaVIyqWKi
Ao3bQJs7x8vLhjDCTM0+aWvTuk2vh3wDjE/ZlbpTnsQp/AvM8zDocOdSVllKTi7/p2gd+AlYQtkr
sW0g2TNz4+kcAKPhSg3/t+WV6+vE5AeTsm25XqVoEySGYvT9SReveo4KfAE+F51ZoQB41C5dTZNA
gbYXTeT9/Q/CxBbHPoiGGukZIvAiOSbpWGiy0mLFiwZUbioETfQqsuAoZy9gUvMNx0QJbapRhliF
CSMqQ1QGYJ/5ymCfQCYxks4DNSDjUnuwYPiyT+VgPuQAE6F0MMnzuI5Vy14/02M5bODHFl/0DYe/
RKx+WdS2BnmR+ncD5tYaucsva9YvYNqm9kXqlsiPfF1N/wrHC7Tg6pkcPL+JxDvrBRLN9ng6icu+
aXERAbbDBrSASMX/62FFxs5vTgnjx5AbhO7pxSBvar+jm5+VwttuobzyWTUHmfRZgZMy0G3h5PIt
phmuXO3oWmmYPFlaBybCN/ccLnkNn6fJzFUpALBV9OLcmnx4hQyVGChlfVCGK/9ZVXiZprK6+OGr
MxhsTM7HvyefmMnlZN59aTdNp907roG5sYbgdbqowM/gDwv+xn1kxXBMKzp5VBt2Zg0B6m/cPJBn
jlIn6jm6mavgoQ8wrPv66tEgLy0M+I8N2/gdeZutFpa1A3EGhUHDS2iBppLDvwo0iYV/vthiM0MX
fD471605mNI8DQM4oGlYfxFUBeKS/kTV+j+jN/XvKk5rM7AdwEnFlZ9gaCYpzQ0hpCOU0VN0piz5
HVNY23+FaeKfYldJ341xpudV7Wsk9dtkEh7r0o+BbTbAe0Zac7zMiOKkoe1EkYSs9J/7OLcVyLNy
NrZeUM0r1z4uJ81SRByHZci9xsIdMTi4wem+dThoH2aP0hsQgY/Yc8u1uJLk+LqUAmm49IbKyz2p
SvobFvfchk04ftMgTF01u/PA63LRfyqHc3YCKgn19/O6FB9nr068R0swmSlwlgzriXgks8c/of7r
ogb9s8+ri6sGSgHJ1nheBHAGFI9MIB/8FzZx5tq2BD1o/RoC6be1pWTeQTW5hhT6VqrxJMvFPa2j
kw0imazNds9yQVO/hz8MZgsfFphRljXSXrPtofqdgZRgcTIa/THebHZF4m8hgfno0yDMcndC59io
HWCBqPCPIik9v4e4EmNyD6QLDq2ANDNsqa1CeTz2gRibzlauYiunnOqq8aDe0/M+Ml1zrjhBYXGQ
euFYSnr/g+mb5we/vF/ZLFrJxgVu53332psIzOgCzSZnob6Qxxx+HcYwoIP/ehcIp2fqxSA2PyhB
ur4Zw2ZrCovCuDdsK5kadQNU7FYfW4zavwGlRUz+POnde2Y45OVxIh0uD6AhIXyqwCLVWze84/Ar
ptVj/5/8hRzcLzDmtpc+HqmlWrax9jeJ90912EBqLoSjNovJIiBRo6zk3VYEZon00c366vgoLNRo
clYrT33MGIHzuW6Q3r8PZebYxDP5Tap0K13CdRKwTqCsvmrfsSUIfXTvyULNyYp2UOyU5ioTOh+0
xEcqGWeW/5R0lYVU8Tuvi9WvkodWIKw02gjz9EW52wbZV9dDcQg254pqFruheWF5p8E3zsLKeU2j
gGfUeQg9eejuZ/gxfqURFu9skUczwkBqK0IgdutJwKRr/NykXhZS/S+qHpuVr3MMo8kfUhcdzYs9
QixHiVJBGFd9zz/1ywaIWwkRjZQSKZ/vcioGSWRxPuQ783r40Go1xF18T61uBddIsbQ9oTqa4QF3
76PoJDx9+LNoI63ZQR99avTOjZfycZGbAwyGcBa7Sm0M62jyUy3YMWmvPly9VlH0jmY1s00BxkYv
D53GBQJM7xag98SwR+ZVpSvgcmo7YBXRHvn8Q10V+UeiaXGNxCbP/Qv6KGL+y6g51uQM06xtZwWQ
p10iAWNs12VuhVGHs/8H3hhEGtEiDlKOs534iYfxz9G5ji3bXLHZ6g9re2JqOX0Rla0ROxf4Gq9D
iIOBgIynTEJQ8steQTOnVZLDBt46m4lMEuY8zRqFD99XldOd/P37CyM0+eKIwewj86Rdtb8KjIew
sytcjvW4kkdFsqt5cp9+nCiiOl/RmqdlA05oe2V/KdlN1Sre/xxFy1Ns5isAzycezRFVXKp7j6YY
yCNOncpeMKmsGpXBtDCqLfceouQjTNHe8cLVL9jstVWWa+QUghBZ/8nMMZN2Fb7UJe/ks7LTcssk
bYzbF9A9hUSEBStu7sQriGq0dGL1MD/Y89+dl1jl4Iee2VlKUEz5MQGAr/8LYvNaJAozs+09EeXM
Cpa644efTkfcMkUnzWdd3iFGBFwEOVFBvWMtu/uNFVyaU1UIiJECGSsQPn0wXHhknilEicwpo8SP
/K0aKnlxl9ssKPHh0lz40mcWYdO09Zq6q2YucGC/FWA5r1pUwfBp/lCsw+PqNSBfncyVQvwb6Zcd
QfgehpgZQYF6xFlBfRgcy7HyRvImNAikX7NsZuhZ7C+0jVsDEPA5acrEFRjTd3Tt2JuCtbQyM3mG
sWGwhJAWDjAcp+hVYqOhl+QYeMEN/mKm2V4okreKn2vuQrW6Si6YRua13cJ7kLF416Me3yEX3uGq
eTmXA/hIaC2tTULnaFdDzO5yEXP5jd26+YFItvy5i5jTceIb6DPc9rFUuACOOSSoK2wzeXMhwt3c
hg7pRJ2cJZu31MqBlI6wm72RVs3St8nGRum7T3lnabZdZ9J+eU7EUO0nf28SshyaEPasRJLC0XOK
wRsTQaZu4BmvKPTLkL57cvTDuXtVOQt1ZMVpYcu0WF5XrzqG9cGdv162xA1JRsaQrpKigfkCoct+
pb721Hiwu9aYi2SgnCz1wpTH2Cy1sLbu3iyT2ud7dniyhgMJSVeZ79rDoDaDXfEiIvuD+H6Z8ibD
cM2Jvj1c8AF8rqmXFM/Yt5fKM1ve9+wSZWCITH5wipORPMi5mcDBzT2CXYkiC/ymx6pvf+JPy1zm
01m7bWAr0T4PU14WsLiuVduMrOcUd3GnDHaS0RtHGZne2GeIYqwGLTeHXMhrqSMAWGuS34gD0ZXX
ITmfFGPbSfW/uTn1Pw+/Gr3ioTeScFJZZpn/WCqsyAmNCSgmLRz8NpVrPE32/ffIqStAPhT8VlZU
PqFJ371/RvARK49r9D6Yc+Of1WPyphDMqyx1HAv7eL7iaUXeYhgtcqqtEY/lwhC5d0VCj1Nv8EJw
08IWjmBCrsSpqcptqSRNUpedM30S2S383lsaPwN17zDDF6LTf7glGeU98WzVI6RuLoTwsf4WreHK
XqfJL33fiiBL3NUR5H8ZlhwSUT5gn0145P2FatXrJKE5bBS3jCGYNDfu9Hecbn0crIoE5xhehm5Y
nYnYVoq/PJ/+QcBIx/pIhKGzs6kDi7+CKWBX5TqQJ7y04tgU2z86pvHmjEUjUcMOI+Up+hcwktYg
IEagJCYbnOV1u5Q+hkxgqG4SXH9zM5nnu+7vboXiLUP3p8jo8mBbJJ0MZd2ns6BQe50U6EDT2p3h
uNNu9YO03Kc1nN3puxh0HA+I1nBLIsZf9Qhg2i1/HylPuBU3U/Ow/Y/8FAJQeI2At2+zp+CjyO1P
G02p2BHpbvWoGGlFGmePNCop5d7Fpr6j5lBqpcllR7NC4GPk8fAr3EXXrow89Y55gPxx6G84HQit
dIA6HAjGm18T5mlZQAjPDoyuez9zuaaKpvVGjec17YAlhbh4PuWCVAUhi6T/ikUvgjJlW0pvtdzy
anKmg9JQWBF5MeyZinrhzEiHjGb4HRTXxTb97ohM04RIOLAMXqfnAGi7KTwahgiLm0WfKRucYF/s
rnoHjM0zkSVWVByX1PtzF2yOnEbDKCystIg2K70fUdTXVB2zh6/YZ2yJSAWo58UtJJHmtCqGatBI
B+N7GE0qqrxZmgDZ82D96UnLSWTJ7Dwhgy0+9ULB+g1QDJnJpF3GQ8j+bqsIZv19mQtDX3cQTMQ7
djfzf9necOANYNhKhQLnw9Svv6JlWd2XMzDyNcCkzBTlkWL+QfbUJiDZ7gM6/Zbq5Kd38aSkO6Vs
yE6g3KHrpJcJo/GAMc8JWhANNJp3Ku12fVMBcR5CXMxwCBrBX8x2n0pm2M8xeijnAYw/iKaBsvc/
phnfxyvoWkZh0gP+Uh4cED5tLvkF9mqX3zyDnGyk/HvTP09MLh+3XXXkEgrZz5cMDafMTcIDRkvs
kFdhPaHnRLNd0efHi6GlXwgs9Dy6B+7GisBm+Xukn7ybkggT7FhMdES7wDgD+sFd4iPAeZlc0ERe
KQ0A6YMyTbUY62sX+j3K+zZUjfkDEBI69IrEZmE96DBmQpA8cOAY0seHepTb/1GgjTUT9OYHhG2q
76JA2F4SomH5Dj1AMQMjYSq2TtNcZCBei+zJLeU0+YYQ+Yv82f/Qvcv3+oU0onkXpDy9zfyIRWGX
8g4Hxb0zuLhrZNoJLRlpisAgDBCptMZy4sSVy6pbyOhEfz3TjEn8O8E/XwdkrW41OzGunctRvEDV
ipzpOuj0xjez49cgw2kARRfa6uwqC7GXfEbv36MIEig+5Qj61xX6q8pzBgUXqPL6AffHxHMKa04Q
cArlyvM2bO1zBN2bQylFCRsfJsPRBVR34rGLGvb4rlMtBkNj5MMdZev/j5ye6WOVPQ0PAqTX5T4B
GpQI52w00yNnxPeDw+RMpUN5cF22MUEofmIiyaPk4dN6fJj1ajLyK0VAY+ziTHnyG6rvWDiUEhve
KLdb7GLVW00sNG6+LcDDjbGojYwpsXJ1xQS2NtzzKQRGEM962ksNCFy+tqqFC+SB/xOY3lkU/Az8
9eQBVkPTHVBn3VaP2Tsy8XEFGs5mV0Rm/SjD5Gc8amy8yjNm1Aq5G+Q9+CrPST1Ynje5e9SZOJf5
eAleEUrwlsVHkaY1pyrubofWuE2W9kOqS+16+MUirjQ+d82AG5wImzFChPZSlxi7Xfg+E8mG4zsm
OpNARpFsJ6dLumHPfJKma6bidQmYym0whZUnR5gTGBx36/NGDIxsFtqdUaEmJ+tugFqZywcnn3xT
AigFv4xkOwSyPRvI58IQYsEnp7dIMF5l+18exZ9LA25Maez5hsQTZmKaZkG32v4LbxDEnkCTUPOx
lcpS1nmKATfDK4rmqLu00grM2ndCmmcbNJek0nCEo5wjHp31JMcym4kKh/kFHcZrWsb+FenjVhQl
xr2I+yaO0tt6aKEUSJl3LDf39g2kIFMzlPMPwJXgcTQ0Uj1XYq4VpjkATSg4KHlFpczXYuCcis1u
67VqDlsfGzfe8Aio02shDjG8DfyHQZa1Vn2aEkq6t4fQVQ6LbDerX5h/JQjdUkTNvTui1+bbpf34
u6m2ocU/AvqpavjleTUBNQZl/viHN2FtfRDLGRw3Zl6Q9F0E05QMMriMvyH9z3AMxKtfbipAzUH6
jnELLQ6M7T8inod23690WW7UJfY/qAYIHusp7d4+jssJWoRsJIDBBmlvvtqRNjtiKg5oSWRaozLc
lVZoWN1+Y8UwWHWI23kWzW066xHl
`pragma protect end_protected
