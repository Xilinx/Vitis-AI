`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk5jwBRWFSkvbWHGfiNuNq0+Y7dg544YR4dDn372hmY9j+L+yzveYCOe3
SZByyr1Kp90wcUEL+uwUxNZiYPiDjcFEtL8yPG/ZeWaaLQEy5u21nK/lyh5C/RBsuE5khshKYdwb
CzJB9+PRkATmTd/vtGCmeI7q0Urz0vPgGOZv96HhKniRVJy+V3AOjqdXML4jsuJvgmweFHMMqvXI
KqByGOJotwn3QtQbtgRUcFsgCzeicqBb14vtCB6t34g3yJk1AJSbajt0at12buUGkElyVPzWYUdV
ybzY6Qra3bokhoQrYz9hEJG9wjqi0C432egcWhK4JE599sVspVxTOcWDkaaeyJYqiLlEj07/UVO6
/3jKeNmJYrQdXv9JGs4soKeRrh7pehU4KruPa2/ghPM1iLQOAl8BD6lp6oKrlRjC9Bi07pKSO0zv
tY10g1nvATtRNlIUwEwkACcIVIBSUUhN75pXZe7xdy+vj7MWv+8LgxDRMKyOVfS/EjbSQyom0U81
hLcfPD8pkcLDmsIQZFQDK1N6GKWr0CUEC5J1Xjv9Gno7XyE2xDn1ryUjl8TynTjRYnQ1MzwImc3F
qzxSX96Hrp2TlgaLTwYi5MTvuMwpDH0RKCN1gHctIPU+WJGqReOnYFwxI4nb+1aGL5q3oX2bNymx
m1LHxw2+8sPIEhIxj38repqkVC3z8splcZRD6NYMcuvjhq7SLdsHH9NJTY0/8K8QwPrxaQOVIrpX
3ZlPgzpgWeIPVK2Gn0jaxtiBBDW0QHYfRre3E3ApF7mC/EaGTu15EIWzgag5Qh7YhmuG27+gmGr1
au3awP7DJaQpo/p8IQzo6Klebp3G7xhXCiL6Ov8Q3kFYSLnx0MvwJHoUXpPxXGKLwfl9sRuChu4e
qstgOebdaIJgI+z2jOS5loD+gM3OKA/9YZHIyBEA+Htoiurhsb/4rl4sABZWHeYHYn/lOgPtTF50
RBCfLZ2OpAZxscr/iCGCEk4YHRMrlQ0qPM0z5XRjlY+X/iolgVcq3WDBurCLUJZwg1Ui1Wo99wwz
UAR1Q+yOeUUeXAze9q5gd2YnblaZdH2jHpYr7Q37YxS0NRL2tRMgjR0s/+58hwcIPk55je2QPo9G
Nq83upun2Mpv1OWKsr60mQcOf7lKK5DQ/uOpbvOsQQ56+bBE7l/uTB1OIhciTIGEvSY5s1wD4akC
w9++qmMPkRTUKLow5Yas2PHe4OHv7ywTsuKkcbtv88uV7La5XVQMbctjleVhrCXCi2SVckyoomVT
0QMdUgyO2fepZk4QKDyQoFfQhm8haDQkZhO7J7Q//knM+KyDwXo+eSu131l9efhxmY3wfMdm6pXG
uDyyMCkozQQUf/VWKO5Sk5kNsz1cn01Q+vtQ3qgzHKD7a1FZH1xh+bdzsKzzcM+nL5JT02OLnwmS
RYsws/2EyYFZtIt83O+2b186yD+WOv9nVb1watCaFW87Lgbz46cxdN8yqWIGrUJFyKyTxLQ6kcEz
45ry778OG06WVx4zy0tAuM3jgC9WBEljP1NvxpmVTIxu/2ZqObKxx4NHs/YTc3bG91kLGDOJJrW1
pQ/FcNf0Pt7638+TDfUBLDVWqcPENlSJVjHyc2DjkOf6BnQspMTjXOhwZnPrv81/vx/tJTsmJLOu
SYTP+KYyRjWWkjLJ3dZm63TVodgmwCjweNH8AafgTmUUGijdOc5/HidKUUvfOkMKZ6PZRDn4AYND
dtC0sgASW8wVqUZfJT3M2Zr4hy2a5SgoT3Ps2fdPwvdIhbA9r605WS6S9kZ8QOrjiaDD6n2yPKtL
i4y+xhvgMHuAPht0GOTNC3YcssbtUjOkos75J4dmihAqAFZ47QA5/8+0WcSZfIbWUBSBx1WfUcQ+
fZqxULyUsdug4QGAE8SnfReVpM92sJ5Ti0HiWGCojgF+tcjKYKUm0eyXvkKwfaCh4Zs3JFKd2RMN
pU0MIGKCNLAcPLMjgaHAbfuCuaGuWftAFg7xhQFl5dmtbkaDcRJyxocnq9kHBaeAfe/CrcLc7f+I
10tGt2JsyJ9MqmXrX38CoHkqcB76gmjK1HQI5sfRxMEp6OA0TFe+1zwOfB61CFCO8S/PGEZUa7kg
c00OjmLNwZqjE/dZeXjsKrI6uMLr7FrL8bYWHwByq23buZ3GzvPHr7EoqEuHok3RaCsPWgOk4C5q
SOyGSujparQm4a4SZlYJuPMCgZEvOdlhZhXFIqoNHs2cyZSyWrB31TxqLX+ISsyKAGDp0F/FYTIN
MvKDYo/cIbuj+KHhd1DcK1ugnJdc57md5rHLhQDuQD7u6ZYkyhOJGndYJHbGBSEgmi1MgbxSIKbK
CpbCssNmjAn0MFpViGBrj7ihTvSlYxpU62QzoxvRwluXjk4yYUZLQ20W+bHOalrusDa6kPYvWkT3
RsDGmLAJySgoDofQIDf5JHxxycpOg3221VZAFzb60N8S1CxO1LKqGNGkPiPFLpj2tYwIGGF7A6uB
XPcKHFjCq4gd8R9PX7vN8u3w9Qih2b8T071MsgqcY14hLVBXJvvL0uTM1J/Um5OWCJV2y5N933zB
pl/IisJrChRwaMi/9NKcn3Hride4l6G5HgSznzNibOtlc8T0+1T7SOZOBKHgtRvjLbqYa1IicDxX
HuNnAK8CBa+VK65fS4z3qYwnExvx0eYKXfadfuCX9rjrsRjPqo0FMgvORYM7xEk6nv+DXk+JTkxk
olRpSfGGA+wdw2yYt3pMBLr2JIFUxXI3uy/gNF0zanuszmn1NL8gDugXOfacSk2Mzl9NLIKkWw+T
kOgNLUOycYEYatnyZkcgRONtvXqhwAdebyiZ9fM/3JDNUUiH8SR9UqFTg7RW6WS9/ovyMVkgc1M1
5ob9aTYyEmmHg2vmvRhtx7r2QV2qvxCTO22W2wfDNAmhe2OiRw8PELMXj8Wou3ALwKFqtKDtODPu
aQSZJ1Q7pOkTupVqIu2rL5B9LYOrrN5diFgYF4KKuiWWqkx2hL5sOE73Z8EZ51IMfVJPxqKBX47/
aGyIoQPCY448rPzpm3A0DHxWFK1xt0XvStODX9zPb8Lg0b1WpIsXNHs/EcuDw9UddjxVpOqKlwzg
5KmhK6CHQEYw/8v+kKKgBJEKqgBOOW5nB9i1Onq8h+ViybRzD83sdjRKc3OABJGG4yCdTEV2xgTl
anQ3QoEHof3VrWOgVl3vIY1+sX0H9X/wdgtI+mkD7mx66rXT2rU00gZjgqm+8OFCJkXKqvVtfN3O
qiQmZLVaScEQqs1UNBs+0Cdpyayj1k6VgODmqM/Vn+Q3OyKqSPNETD2HtenjZf6NgvJRfTn61ftg
sIcDaR3XnMntrU1fCHakPiQ70wq3kDmCiumMN5Tx2FzwsrSllaQXxKhReFpQ1r064+uQUQyOuiJE
sexLWU/gRNEshRhKhRiOip6PMJ1MsN8q5U3xzQtUTZKEBmq1sXhaLm6JXiBniKJSCYs1r+ed+FV1
gaVr5yk3xfNtl9NxiVpNL01GwBFv7IABkKnoqB41XWXShjckZCyPDFhRJtJNglRHwXq0PUpAL7xu
hGPwI+DD8trtPiq48+H1gW+GaUe/d35hFBf0botr21OE96xbmsuDXlvC7H9vJ6KePOYqlzjchxp2
lZAQYt2MFDiZ/gtg0SYTowW+84PUZ95++9Di0EBj+0Y85OnQeUTCy5iI4KCxXNvvv6LSkLcY9gh6
hyXh7ReuWd9lBwOeGQwsNfmicjsEEZNyDiOIerDS0hSZzbs3GwWawd7T/WMMZwlpCb8jmd+KTt1r
ed5Bl6vBaALBBndJ9nPSqYUxl+MTRkmyVCyPNXmrOnZl2y8/2i0vgFTDPYiu4Q8N9KLd5MNL0S9F
bMBdAy6UpPbB1pfuaxrbr5gLh4tHR4/SOC5/eh54Pm/yuzP0b2Cpd+XvfYGg9zik5z9oNO/gDCSD
NEf+nncj/e1wJMIq6o6AQaXA/3w1cq7vVAtyA3f+8JxSpKNpmgRoAWIg006ox0aU3TF+35jqNj94
8bVgZoHaTjfb1jK6IJkOOb62iHQP0K7rVRL8aImVDk0y1/rIhwknpVha8DARcqtoALpTocsEJ60H
k1+y/ic9gfis3cGZCveHuXhh6Ezpq6Dvx2bBo/vGumuB32gqjEZyE93udYzjfcJJqtME+L6tZaAf
aDd9fW+OfR285SusPrdOC7wANNylt024+WHLFuMzk3YqoOThIkW7Dm6m4dNhwmUzciSm7qgIOfZJ
mWLECqF/hXRidgi4tZTBQunvYE1GhY0lye/Hy450M+qM6GhEhBezDyDYtSG2eCKg9/UnhCs1uoLu
Dmrqbv1Kz1cRYUC+VBtSyp+VFzsk5KrcWH6vwWYVIz/XuCXTUcnusSQVi59YvjUqEl4Jorqp29qw
dHnopTg5SOO0AUFUG8sAtH4KRnOt7xGWLUgqEk9/aN2TX5EIY4vCY8ig28kW995NcXGU6YyQRq6d
G8wRR5HZI5zmt8LpOW7u5v8b+rBZbJ+Pipjjg7q1tp5pMJeV0/IyjCKF4oGXzN7VD3JgQeklHm6o
nopvIv+ut6HQ6m1rXxXUAzzmNrSRXlJ1K8kmH4urJ6cOEz7eTeOj4VUzNPNo5VfTYFtvrx7ROjVK
kvQsLZZ+L2ImSTZZrF8G9Qeh24yIcWRswAvvmixuHF7JTXrksjj+TFuH9ULVM44iZDDzHTPCA0ba
0P/9asThm8nhbhJpHtSRyl88BrPPZ4DLosjBDgIUJ7Bach9cWu4g4UIJFqTqmGSQ2JESsWcKux5i
JyurcqgQtB6vm6PTHAQTVesuUZHa7+mzfxbRuKwH8JmNTD0Puhs+xN0A/YUM+UDvwBYPSQLDduon
qajecBm+e5QDiSqwKG2oOAggW3OK3WMmxQ2uJvitOyZKAzVfTQtjLN7eLGjta1ke1A1Pn00pRTQ3
zHNgvo7klV5YJ7X5Ef8L02ZhG2o5R0mwQtnZfFWy8OECY+X6zDiO+amQf3lgymqeM71kKN9QbRWs
/zNhVteKQYJ0eil/vmrMXzgupNYlSNDWWNBzBIR1CALwLjNQOMsT0dhokW6dFlSdsmu4YGQl+bTf
6gsEK8c=
`pragma protect end_protected
