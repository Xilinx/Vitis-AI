`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15440)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPak/iHwVkUKXxdtqF6qlW2P9HJ89gT4zeosXKnzybBKQicNksJJ3BMUpsGYPD9ca9gUeods7
apLQr6Jb2QsIBT4RCOU3nQGexzx1rZU9heTO4NKwVLFMX5LpT+g4SvtDdWTD+FUs2nl1ZUJHQwpd
wOGqmHcIRRa1Ba3IX2snfjhzyafROuaqh2H2nNkxA5nD8yU5+urwr2nsNxYtf5Wojfgc0ih6PNoG
Bu8xN5f5xL/u0wDuzoGASldkA14XGyIr0Gfv0kYXhW0b1fH3pw7E2w8qLZVXJC6015HUuPu0+EpG
SXHHs0C2NYF4axYjyBCupJ3ht0m4i6Oil56m/AUdIctnF/xBUP29sMZlPjRRZh+/NeKtePRmknGM
/YTKnnXejiKV6dSC7cI6rTKh1yAO2QquQJSl299RwZ6xFXYS8h+aYNtDq/btLOkeypZI4Xb+ZaRH
Xzpo21TxnJDmtWrb8dcJ+UFWWHwyCf+ONcKfsZyEkuj5PkqwSZpnfEahnDB6dOVNLJY8JuLnevSn
qBkl783qVOihq4tfJA3fJD2JGeYGlMskZ5d/odsScmc4AnRwkSgP4jnq4GlPcssk1dN8gehcHm5s
GJ2h6EiuISQeymGQDLH4sJZo7+faB5TAqJDp2DvwAdzKu5rq3e3QHzBDXGuTyJPzGD8jS2Zht8V2
1/E2OhXOj3BIFseQrFLsFidQI8hMZyeqlHyntXMRHo2MxFgW3H99MCGZCsxveO0P41icUaV+w/Rk
H6OHvRp5dsFJ1HdBRKU/D2lX3fiSu5gsxtPVVF3n8waTg47cKp9RtmRLMU6T1SeWTx2boF7dp0ag
CvpH4N6rhYPo/zeLf9aeqRTbAyb2H+O2jFWUAW6FDJaSPaNEm5YOvvL1zUTs8htqQy0D1KLRtr77
ZB2twPMQ2KpbUyaA05ddPmA3NPsnvZK+oK/cdY4/Bg2jqzgtJJlSSr/64JTGB7PdYc2QBLRfpOLa
gAQHpm3WzgZCnazVe0OVXz62HL/o2AsV9ImMFllxAQ5CE1syF/aSdUdoh297By/HQ0P+uXJ7JKQI
2nDXzLRo42zdX5xfNxmfUim1s1HorSaKvOG4Yr9IsnTUHXIDVWfikZyjrYfuNo6RF/PHmTbNgRRX
ZSFpleVN5jseJe80nuk0ODuDId1b0t9wKj0PKKt4wcix4SiqhdLc1OJbZIQewmgaxcKuXTYcAkwP
Eq6n5b/d0K+U38uToqXHSNWv+OCA2Mom1IokoQdaUe61Ep2XDtxomosuTZXCUweQZ81T1i0QuNSv
A0w4IEW0NL3JhvKwcY5jlBDg1sVoHgHJuMMglFNibQ+sZFXrTHoiTZ5zNSou0IG/9uA4VcgwpLoK
wPbQSf38xEbfnH+l+gYN4wbiJb0aWXME2Pn2uWe5yRGvUU5FaIVE0+FECL8P1YfBNlnddwdsvJXL
TEIf5GhSWmt2e8q3xp2wi5PHZCXNsl1CHPGeHR6MWy2JecHoRsunXJH38vV/i8BSzVlU19mAa8n6
7pQY3WsKXFbHBuV0aR6SZjd6xDoZX9err/zWu4Asce4oY89+rkQKOLwaOU9TUa9U489Sua6akMNT
L19Q9gjOfKLLZN9Ixn6VhPhuC3DxInhJrcP79jYxwo9xC5c3hr8UvEzKIBLdTSjXjGHMAOsDkjng
zkCqbZb2H8IS+LM9izewy9OITvGe1iHUi5tXlcg6ERpsJdJ+pw4fsXYlyIKuWrhZVq4fgJ27V9ec
vgVPQlxKb76L5CxY5eCbAaFloupS81KUWyZFAlVxn7eJiKRnRnHQPfkTrCvMJy3jI8OfDkLzmj7M
ARTJhV8Sp609mqeJwpOodNrRpK04ghDktW3TgknUh82HCOE/xicY9vmaUj1XeXFlz+hkfQCPd8tM
w+nxVq17+MvicmwHtOlyf6IrgRGQzDnBxRud8GkCxvkEMcH7witBbhTXtI6cJ+K//9TQI/oQTz9l
Y2HjjuRSi2BgipJ4ZNVfkQaxFayVfRp7xzAw8bXkyEoptlIB+i7m3C78WsYInBeLDkFHsTBrI99F
1FL5m+o/5ieSfL2NIdjYRVIGhO4sGMvZ0pAbMdKp8hleQOf7ffTyv7byStteZ+cu9UklRvmyTYEe
7ls1gp8NJnPuH+MdLGmEWPPC3olGGuPGQdrkXdWC42HdS3WoQUDjZlaIslH+JvNVaySHM23k7aYp
WFuvhryatwPT24KCDBxGmekjiWJD88L+2rAbq0zpUTS17iHbmGu/1a0f5bhMrbl2ft4IDblJ4IXZ
GqXg1qw4k85PEEhSKtHk+dNVT0Zhz2VHreKrf0YOf6u8PSE4QMN6f+Fel6/Y2zmqcDYxeVkifCFI
7LAg6bkPzIsSBgHi1DyOCdc35r9okflPkTC5KiYNxaTu+g4+ZNNhY9oSNVJntEJyMRHszV0t+w8o
lmv+X2j7TByCil3AmNtSoi0ipVu2hNsusDZ8RLKjisOgk/+xgQJ8MsB5zSeiif83AorWVDRWb5Uk
lcX/hg2rsaO6eErLYlMIagOc28FcLOyJuHIUCkT+5WnNy0cmp4Ee7OM2gfI4vuthURwisoAdMdyT
KOmanFT4JdVuCBYUVytwJ1XKG+/sbqpJqAjCu13W/NYbbqIm5TMc06gpc4GWWv0cROJHN8R72mB9
kI5eszjZh4AgfZ94JKI1qjYU/rrYuAzUFm8ItEptuP3oMnjvdjsQZD4zm2+FAssqorbtxSP+reE7
c1dWn/nHI/eOqs9zhv3hI/rMoApI2TC83R6abUnQpHEwU3B0769k9JC2FszxcXvVGpbvpacgBc31
1wOgtcmN17BCKeV8Y+ltfMYSnY9JJa15qBuaXWA/IRgnxT9TDUXdJOVXnktZSbJfvqtpXNGgVVqE
5PXlNwk3BUS6iry6acWTAA5xp3aVDqZIrUKHqbesQKWg7hVUVFOaaDmX6FOWHl1fnI75/uoltM5Y
KH9fLsMd3TRphN9l90VIyeUjY0tuw1FFlsAVH9u5Kl+OONuZnlIMDI80pbOtNH1Zmw1+BHLIwi6e
QCSN0jKff+j9VhVekfdK95AvBZR52eW4EUnQ3K6bUpFQZT/ZmQvCsZvG2vORomojuZpyEyibww4Y
yeq8L9CWFCc6ubtRQ1ks/BqlWZS+744BLzf29lU5I0LPJhNd7D/zPl7NEw+SPRkEgLyiI9SqlHF2
rK5etqvVWiH0tmq47qIRSpDZw+HUe3tRkYWTJ4haBq3rlJ6BYZF8JJcP82lFE3F+ANCbHMMKW0hK
TgpRiJsi520b6LsDFB+4jfCI1+iEvYBr4lyGsAyNFjtjITqAFiU/QEoXryjnqVyPjl/5FMxTDyxe
bEE0vAr+BT5nSrmP7xxekyKtyTpfr29H4vtmafXcCXnMtXMNgaeuXIe7GWj3OnVCswWJfR4AzmDC
eQSC18Ml6mWBzIsn9s32QA6/6FxVd4+7s04yqCH86jO1GHm3MncBHt31Q2lwZDlvPSocHFrtGaTf
rKT7j4qvyRvH5wjdGFFliUACH1coPfhlRIAGPTrITvT5+6IP6Cs6FC/NQBa326sOJG2Ke2UwPukz
r1HLh/DQk1Y6kL11pJzgNVn8afs1RNZEF07ZDari8jOBDojVBZ2PADe2QUqVjoEN4aLRAYDFVHXB
7XJPOH1emT1UQ3KysHa0vWr/bKh6reKm25ybQEaPs0NMCBAM1iS68mPF2hy9vkq8jUuEXyUAxD5y
BUBzqi+6ah8LKmogRfxzYCjFYQedbOoTZhvWbKA2ne1vahdXZFCRQbzQLcwFfKVJiCT++sXYzYBI
M7e90qNSRv97xHmrG8gW+grivgxCsyJHcVHPPNy64uaqJEDTWij0FgVSnVOx+lDydNTTBkrz4kfp
EBJYgF5hzLA5jGt+tB/tY31V0FnMfolDv/HjsCJ8L8cbxALq4pIV2rCZNCDm9bPMcatna7Hf2IaN
4/oXyqmnn7Vi+5JCS48VDGWL9dMem7CAtJJH3p84lDgQXRX6anrOKoebSDjCTnVPZYVK+viX9ey/
Pra/RReTSm0JU3FERfT0BffUHcAGg2N+sGZ6Hkgjpa/uwwr+X25WtF9YwwMFPStxd5pQ1/4P/c0C
Tbnm0ThsdYUXwnPFVNhNPIEUGhCitefLL4QthB2d9imEAgW6H5gGISOVsE33lDoxJOT15IOAp7t3
7sibbIXqTq6wC22pOZebEg/oG/6a8TdyMQN/riOXmvNhVu8/zixtUAH5egXzqvEKR922w/nqdt5S
ew+m6LCxTzyHBL/ePAmSCpR9rSp41err1gb+IxgK9nDjGBMP/Kw2Cii1ZO5SvIDKzpWjTjfuB6k4
keTxMv19XZuASYTYIs+CgTgR4micASFMVEsp13/6RHZaxqHvnHkjseEr1oRVYjMX4BOsxBuHd8ru
dW7VDb9H8xF0j8lJKWmHCNukGb+IqOt4wRL1L2EOn5xgzmJwSQx83rB7tX97Z17idjtsbpudKyiP
k7AsXTqnyf6I5JyLX+ILsK5w2FmPD0XwbNxruWyIgXUksSjtJ8syA7RV9FyZVnoBLTWTROSqDrUo
S74odP7/bC4OhBkgiSnvSRoeihw6ip3HPY7ue9Km+sow96Q8R/+OgfNo8xDvySwe20dUjEoVCKtY
IfS/0h1BAw+1DBFc3vpTUvJTh4Q2xJNm6kvMuw+OPw+sXBKjnLeKqeIHrpBOeix8miXNxTdxAByV
Hk1rRs81nmjfysHynMhMFIc7rdVcfoDP/4/nnoyWE7ldQAAdtMCnHD6j4C/G5dkKRrraMEm/yB4D
haz9VRdb6RLquFeCb7cu4LaNhgMU1jX51GGjfDuVkgKF1mYufKiVOytW7u0vTHdIenv3/E1QO5QH
jMqFGgWE08PkvWPgiSHIZK5hRWTmRIQZNplIfgVe8vqztcQjeguDgcAWt/1JnVhjeNHRa3SLGkZB
Cr+hII3E8wRcPZ4hIvYn2bKWtGZJ2Xjd2hqYTInCoecaf2aRBhVcfM10DWm4Y3NHHj2ArXofrg42
JGiZiSfCgcokroeW6r6sE9A6fpWMhIVgP29kgbJMjngiwby81YA2wpYhvqAkXkD0WjirZABwzEHB
nYHuX4l2PDXfCO3QxJpo7cLWeqEkx4okk85fjSOIlywnMfgCzzVMOCXlJ08C7z4Lhjb59sUivKp+
Xz8e5Pb/zvacYMRS9pth4aHXldo8eYjBRtLXfWc2soPC33U3p2HyBAZyDw41Dgzox3DFIYjPd8vh
V5Ny4uxBRZK7NMx0aONIdBLGd0d45TkM3ULytC1/4hdHk1EntyDKwfoFIR5PgelcosHs1nfy70bQ
IhMn2CCMU82+AwfRRp2cEC/e7hHye61Wu2XB/ATiIIXRDN6Hn3DQrvdmmXSfolxemMvP5NNluipC
S94MOVP+0c9ltZo4aLIGkl3xRhy/vhk7yn1HmZw4qEpkgmwLEBEHzOZB0UooXhYhtMNlsrScI4oo
vfNG5ZPbWWvF/D8+0CakErMwYfo3zM5Wvty/Mwl/ZeFnZ8NLrE3wrNDnXKWgpGy2LU4vbjHHL8Vw
qARiIhMVIJeYB2jf+sdjbKuhtPNo6qVIPtBkZ/p8R2e6sIA3doXh2wD9Fn6Nna8mL2BJ78rl3KNz
JTYuTqze/CDtTGFGmnnE3JnoHXZpe5o/N378O0IqihmePxugBO3bkekFf0TvTfGNpUPp4nHhD9OX
DjvL/s6hbOKzNC1Y/mlRkl96jdWpgNlndIPMIxvtP2if6uejknttTjSpJ538+nQDlWJgotXZRt7X
w1Zkxo27csXVIA0DZX+66QG+bBLp6kXSe4M9or9jvA5r18o1hSRE3faqXnAOVS9NGQ/EI2pVsAoK
RFk1FenOu/4f0btGvYmb5ciHZbvDw6aLYIIYTqQt6/ws1Tl68aKQFQe3GS98t3kBzYh5ja50FoNj
JSKLsAqOsuIFacpXLSd793Cy6OrFJWQT4qWARWbKV17CSrfelvyPSip9rrVHeFiIFoX479DKFF1u
UY/pDoT+0WsFzm7pLaGZ77qtLLxFnbWDgni6c+iaK5180Wp+Yvn2BhKbKpyZcCBcWcs+yUw/VGmw
tO7cLFtTswqwtO1iwfgvsSo6yL07o9ggbkTdBkcBrYhSJqFXP7X/K4IPHSoHW/W79YhU05fh3+Lz
t+OADvtWucxadoiWzo2LaIoSh+4hfQ/DaL8UhaT35B9Yz8wnbN77+gXLkEMLsUOVO6j9jM2iF+Xv
C+epfg+daZoQK6c4tIeArnYuBLR35Ucc8276EDWwCBSly6t5R2KN8MQm3uUqGFe3a80z2y4vwT7F
HDoWcgeJnbUy5+lLy9aRK+ycVZrX2ELRvrzMsLD3GDMTED347RbVfG9P/p/fO9x/PdzFhra1fyQl
BfNuzCZi0noX/QUP2GnaPmTPpnBJTmXrHVwVExO/3G3+8/UoJscFZ9xyU5efEmgmZV3ewS+91wEP
B0lh4Qq9zpcudlNIInS8pzPZSuKhntG6jcyiRwRVhOhIyXxhB2vad9taPjjot7LXL5ICIvW3h5V9
qU6lTHMzVXowAbjzvsYKePbWFusN3q6/iEvoVwOL5uYJ9fxZETyRjPT9NTfHrQRMzhz344lAnqOW
599Eu0BPnWGgyvapi9jsiRWZA7j88yGo7yWYeTNNSWdJ4/GUKk9+xpKU/aT0s0RGpCkVyOY6hTRF
bDCGqnRTa9YmmGeXcfoP6FI49hy0qyCIn2eNcTvF17o4J3tfgXmFp9Z5+MtEOMAZoClrI7j5LTNR
Ou5YTqzhUmcHRB5oVeKPpdAsIJMl3bhiV0N4Xy18an0QXsiNZKDL5USE4mNeBPjUR0GwEY2R0vgq
U3pvCq3TMAy3KuZlb+Y0sjROjV8kVSb5iirOnDt8pMrfkmqRDqhbK2dVKKezw6FbveyGM6n8MdI5
SoHD+IiL+z1xiOSNrnIbZJOMx05uTDP0FnEg8N1PA0n7ugcggW0jgQ6vyYJGKNfl2v8T+WxA0x93
u+mF2YZUNX1+F12+CKH6F1YKXL+/yl/1u7htpAY3qIC/7vGnw2++7XTEATIrvKab7obtpMK9dQa6
cxFdLQ+ch4GPc+FPJAQPaGZcowv1Mkhg71i1SYIlJpS1l3vvOvKUMbrMgIKKggO5VJtqcTNEKaoa
3PJoFVePdDF2oYjdATJGDJZ13yynCPZu1IQ/eCR1Q0IiBlfRlexXhBprvAcXgdJphpronIJU72S/
MlCVGBkcBvfaIVg3noV0uzTSZ2SEBXYiUtW71jFKhjeHi+MlnMErIS91FONhFnP5kTy7gMpH2txM
VspDORr8umr1M+nyuWTUPMIw9LflVCAxYLTG8nF8Zf5Hs9DWZEon1FCA39HtpqDvuEpgwAP6nAxG
2svxNQD8qFnEitGUsJBs1kXT3awga5zB0aeduDiDRCFrUe3CG6vFET4TSFDSmJrNzV12ae3VMEeC
oPf7wCpKLbl0RInpp7wz4ZyxT5gTRiOoXPRA9z0sxRe/k0+7XIqD612RUjTjVFYNSrnyFv/XuRYQ
y0wFqYoKP9YjfRWECCcbV3Kizn4LgRfWuISZHdpzBBbAk/uevpIQdQlLc3OPs6WacdodUmI+2pk5
wxtQNQyL2uRaphWE6DQJN4LPE+9VaCZYFx5uvaHT5dYS9vH7u3OIk9Mp9/ABV7yC/pIO3iw4RXk5
2xKFASmFaaNGpltDWCWtihf4hdObrWAuedvlY24WlUFQA9C6QYCE2uYSltDuPUgYTV1pjpGCFcSa
oSP/s1Y+BFwuX+C7ZtOf8+q8lktUUczOpO9rCLGXJnJ5iqYCax8hqHOjFesIMC96d5Snnmx3gcg0
b0Xfa7Bs0LQyqqtrgTzDZuYzcWkaCGfXXWlOjZjiScejEQqsAUrYaKk8+LAwCJa0Ic4cH/hd7s1i
Zmnp8zzVoyJzLB/2g5tNTyDce+o/8nqm1XwEbcOwINwiAnvEdNaubaljVFFy2jFBh1zRlJWzg5Zs
CrwdOifoQ2xDUE9HLnUeJIEC8edHiNGbKoueTkfHLT5d1hI0lWV21db35O2+4c9IQIR4mV8swoYi
uK7NeJZLfVaxzBlXeIL69HEH0pD3XbBuBgHMM7+hoUPgPyv5ltnCiOPYeDfwv7XFS9hwihkq668E
pzCIw8RYjPRbuP1GP/N2EBbnDZZOOVyBpMxw12JuDIlcoMCue+3y/atD1O93oqyaCa9koElpobeU
MJLj4tkcreal69s8jGY7eGRMegp+TUp0G7Yz+LqAk205ToN+V7JVPtKZDerQ4vqSJMZHWdcw/Y0J
I4MSxUtDzSdjJY7eM/ll7de3Zhg0lVZiTG100xag2aeeYziAVs0/N/A8FikRDi32B2gSDTqMH39w
24IDZ5hU6iMGvXLTiZ1Bkwb877bTqTLSxACC41tFQ1i/XZ4Sds1D9AZ/IaFpRk4838Q8maocH7R7
F7K0eEdztbWrRgzW1MFTeqreGNVKm3rFNalycn8+YMv5wqUxsvtMBFR72X1C7qLFyhQ5efcKdHlM
sMJo+8XU7IquFKndq9ee6Sd3LJLDccmSjkmQdE1IohP1GWuiHxv11fqR+8iD+usewqCAVfusr7n4
7ZppRwL3QNn1PRd9RqkogSIRlN6ZPXLzOV83+VAQ4K9/VGP3oYtLUpnJ6Sjk+/uq3Z3+XqCCFfkB
NjFRCBi2TMcebYiG6akGXo33wf614H/oWiuasGkbjhQaPc0SiBhNtOZlD9L9qgKbrBqFMLml6GQv
pZkgCAIAdDmVM033do4RpHX3JBSIU0EMGMkKT0dG3JWHuDeVR50s+WnE+P5iOJ4I9OQ6COLftl9X
/VbU8/u1OUjsSotIG9nH5nG6rC8ThANO2D1xp1IZkYDKKf41DCdcOh1lBxTUNftaJEo6fRTAVWNu
9wJF65neLKENP/S5D4MgogLUybIQbF1ShloBWpUYcMD8VjpdvCM0NH5flsZ/fq8at0sHvb3z1KSG
mfHf225Kn3nTEzI5Y/+3sm+uU5j57veUggdvGrmTJKDKkFotrreG6U+59ppr0MBuoiNQGukVPsIH
6IA3lQj64Cfw+xqhgpusdSoBMluwDQ8GmQxkYLI37RTmmpRfHgEz6RabmAFKfFYkJ5JvbepMweZd
KHuIeo4jUPGtrcSfJVzJngjQfa7JdfdiAaY/ObZ8plJ6E/KGk7fQyWXDrikGABPevk/b+hZlft/g
GuhE25kgfS52TurvOjsJbERQZ+5Knoa8MWJOy0JE+2fb3Xj3f4bJym4SubgcWI+BPY6fY3bhzR8K
c8dDa50l9NDff22mQZCV2uefeujw0f9Z979DPtMmInD6ZiYLusT7H6K3HPO7a0nLRU2Rg1P2CRjX
rGYTd0iSXVKNoMl9AGbrO/FIhzEcQKlExdURRuPCmvYrf0ru6w57cwtkTNvZP/HUFxQ/71scz3CK
xwnvwAlU9j/Zg3R1AmuxAmxTw5ZQ9Yw+vZeY31mY0bl1HNw9aot5H3aK3JD4ggIkbJrxRsJmB3Wr
+lO4+23ov82Rlik58AYxTt2L5r0I+YcOhOST+1/v4uCdAC/9KdLwJpYJ3nKqlI3W73mmPfJj45Yh
Kjh5707iQq4We1TpdYg55bTcxSBSmw95j3AHtsm795PXvaU5ExF1za2M/xMC/Q2S25KIPsUkliN7
JZm47GRjka7cshG14FqVz88wxJFXm6CG4s0ij6PzgyZ2/Zj8gXyDeXZQzbQUq0VfuKvx3zY+1O9S
kAEptntU64JooiSaYDT4JIVAL8N5pTpcEGyjuuXzu2PyNr2Uj1XtzKGosF/3t0xYX3X4e0ktdug9
wVO/GcDwPDPHEoLTFPLpaomPZHssM2O5iTc8AHEbvRq993kQjKMsbPZAgrHWBsgldXbjXvzATC05
PKn8pbd6AMOE8Wdh8mBW5EFrRuxOTlFcn1WTtFCGqME2jpqWc2Fct8MB5mTKnjWSyEeA9m/HJHz5
p2UgsWhYUthfKJkMnWKBnDBE5cC5DaT4Hto2DFHMdYejxm4b5H7ukOmOX1kcw0jdzeyoRxf+gcTg
mVwFiQEA8mMPiT/Nb0KbFXOsh3EFI2ioYyuXW4CjaK5Lx5TGqQo5aaab57uvCaBGCInOZsDuTX4p
o7GbD8ky9Q9r4O0BBC6G06LG3pDYVTa7vEU6Ch1Xb+fzv/2560LSZuWUjLajiCA2ILLKEMypQrD0
W1+f47763p0pMlQPF7DInkuzsr+o51/4ip1snCTBGANY8E7NbhQgf5YJG0oOESHEgu+xMPKvpyFf
MrvDDYrdUiK6kWinxKGt0nEF2DAv6R//FIX1bxfD4ToyVHlO2THNY7dKldhQdo6oLjijYMdrsWYp
HB/xpcWhptfL/ylkxUhWXhHR8M4mO97p0/MPmlNyBsScKlv/htolfP+O2HGvpqiJrp4be0RJLWnP
6QhiLUMLNYto6dBIVQU8CqpPiDOKAVYIlg4AcbdIx3CfyLFUqOhFCcqFNudJI0R0Ehwl6kc/YtXR
rxonCL2q9IHGnvrtmQoVbk7WbgE/yiDsBZ2EfKgkKC/no5iCAkQDEvzG5kc5xVYX4GANYnoFDq9X
AtJAC17BXiDiAVHDozA6N0sPRH0VAIgg8zs2H6+1UV18RCI89e7jdZL35eGVVKF1uLaUkYQIEekj
KsDhZLUaMGkCfE9S54Ftel1NsUsZPeiYKb0UFOBP4Btr4vV9MZex48SoWfp0CKykDsUg9wJotdBN
Dni7uPrNv02N1ttc3oz9H4rzncx8zrBRAFFp5Tx2FlFiHE1SpWkHCSDGVI27Bm+Fr/ouVOEl9Qzq
xMo3sbM2BdMEntxU346r7b2wctcXKHUPDgKbNCzi2muC6sLri32T9FKp7Rpb0N3nPg6tjsozOHnP
pLrfd+Hr2WltI90nSCp3LHPwM6Plu+Ecx5tCY5j2NdKgEDbx9Bia0wZPg6Mtl5Qrd9uigmQfHkSe
o1aL5sZV7LAvABBxdEyxxZVjpCLbFDpD1uH6fZ8T1sPxVHUmfagHnu5aNjcK2Ne3EmIPasW4SlqQ
rN7ZDvKEvJeSt2ylTZ5ExaRjPVQ8F8CYBn9wdFGQ5ykbTRbtM3685EaoO01AapkBgGlYCbSiSgB1
0hmhXFl+ALbZJUe2tB5gNCEM/t3+VFMUmTwuokUN5Ztie5ivHaF5K2lwA8YnP9+AFJymP04o1Ss/
8ewXy7WRZ53Aw9PrgXqo87q5xrJHA7M8rmRpDbfmpgFers8T1zuZhzMUiXSQWK0JCcQOcDDqKZJB
T8ilo1rKRCBgH85QEcZvwdODz4c1eOFHDWltmNNIKGa9fXt44mO1C7IApIaqJCr7Xdm7gN79PQEc
eaYheDWZrEOflVOaWbPgIcUoJLYDW1sU9CN5YHwTtShxCCUjCf+lvDfycZkTNsWqouLac+zrOdVK
IKCHXTWGkwDtqvVfKL+4ntHduCpoIdnSobEc5Dl25EZ/o4ZoJhDcqKx7Spoy8N9s05Qin6IPPMOx
FcRRd1eQZwmZsyiYzUq4jilt6UGwEGBNIjNBKmzNQJFUNpMaE+iFKzch7VpNOPtVZ0CfklLuX9VN
1SJzxDBXLE6vQqXUvJGClxAca0KAlI5sTzL9JOW35l7tLRDaGo77v/FWzojCFE1x51idolQ2f8bU
WBWG7ozgiSvgJ+wqy3t1ItiJQhY8XK++NMuIpk6iYG34EA5XoUmjKUdCioCsmFD+XWzVK5pWekON
e8nJfqLVYIaRFZGchApOg16lo+NxcDmY8e62wqgUJKsySB8uTHBq15T0bePxWW/iK6qI/GE5C67/
2SvtcmxZhp4Q4axF7IfI+lTro6Qkq/6CURjOR+bsRqW9S/N26AHW4oNYh1KJFYp1VyS+lxhtkIhH
hLV7OI41xMdMQB48IQX8yRiui2VHWctQm1vfInbwVNcmupwQwFAbCauZ9kU0AKteKhZPEJrw1oWN
f9Nv7FcH4m7nm+I2bb9pPJ1Pp9fodrNn1hXVqHJ15LpwY9rSHgRXV48+qDdc1qULT5ORbIKn/r2l
LC4zTrmyb3pEEDUqO+j4dBu6tNPqV37tMPHi1ibImk6uTJ3nNnY+7bRHNkhdYwtfaMTykl60oKQa
jQ6YPf0knyVcsOohHpOI/IIk9EX3eH/4GtL8R5kmSP6+to/kWN76U+ANDYuZG2HoTZJKIVsq+lvG
SqgABD5dY6+DJcHBAlk+VOOfO9V8gqvlBQHk9/qP/yvQlY3EONQxyIVGXuOlHGa87zCLex7mkzh7
jlPFotbCkC2/mqws0LUKXOItv7DrKUtQKOJ0qixFkweaprqcXEyO/6gA++O37e1qkjVbvUo6edlR
PicwbhZqlV2hNHRVD/1Mu2v9QOTn4t9N8N4prE4Aqigpr1F7pyL/mBNd9jN0nlldwkykNXBXnXJG
qy31792s9y1zPhNABUpu1j6WfAqGNkFcim6Z48Lx3ISbUauMIKgmJPJZ+IFD4ftiak8EdSK2BYWv
Ns8ulxgySDmOLm31tOv3sTpx1rL0YeXYakqCSsr1a6sQ7B+7j03pf064f8WccHt28Ih4ds35d2xd
Qskd77Dcnk/0wXCyBWspjananTtP1xDoIGTlRgANhgKGxNc2jxKD5UYLWu+rK1bcyqXqcSLDVhAW
cyoozBi3AH92YagjZdaI+2JT6x2oJrmjQcWuzWikLJ1+14eTApLVawTm4BG6YBd38FWS5GrSBAfb
eCMqeiew/RQ4rfIi8EWfL1QGojf+rRKPRuG4ZZutnNuL4hAnVugV8fpYRrXq6DhS1KQanYnnm9V+
rZ6rrBlER/mi9ezn4cm3y++4aQ6VzdXm9pCo7YT9xedvQC31i0eCtnlPlF0gCIE2FqjJNhLZqpxs
vubGb0vn+V4h0koQcU7btOT7LoLgsFmQyOtMYNVMRmJ2CqIzwoxujObT+HpeDinnUD/ZYQlfiP15
dM9qeU0VIHtcT0lqqsuq3hh/OBowkDNu//SPLGa8Pl/TpjxUu2DSQtToj1xc80KC0cI7brWxWvK8
nhGFBWFS83ZL/uwBSPzsOoKUzHpMtYpyIDZe8icbXZsdLwoWTZ0ksTNMnC/IabncOoBi7dG7LGB3
7i9AoPUORtSMqxnmsPby97M5cie+ljGej0xP8o9kQkaAWWlGz1X1C/JDm4XSA/vZrRzyAQmtrwyf
sjgL1tGJjh5MNfelzyQsfZKlBd7aFbfryZmG5TD4buXjHteV2IqenCLIg2G6C7KzKKgIIgpzyJGn
n5gnz51fwzaJ5uo6D5eJgpi/C7lry0gAUUlL76mMx+z9RmSq6Dlj3c+7nvqUoB0Ggr4uBMJe6I9G
/3wQsYBdFKqT9gwVogowzwZGgevzWqS59N1VTYnIrhH+ljSTP39VM/1El0hXf/vUb5gMPh3NtgQs
ijLap/XPRGdS0xHe0hBG/CLD37BxQk8xZh2oTLwPldEWbAYo2arYdHj5qE3LE51p4+f+b1256Xmf
ZdmfdkG6FrlttOoZDHoAqPwqzaJ1A0Y2okJ8YlxG4oWsrCrNVMRhSWfR7410M5qNeba3MSLvcgau
f6MxlTN/VD+FtavpMUJAVnVNOyzBac++HD1UaRLsOMiKtSKy+JxDPJ0S1Jf2u/g+XsEOAasX+Jes
im3HE+IO2gnqMGxL/zMe+1VmzxQ7NtUrpjelC52wAed4qRZZA7ozJwafw3MF4XWIvcQK3jCr+PN/
NnrQFdNLmpXQOC8kU14CFeq9IVmuz6NhLk2rgyZc4YlhQVNZaVHiz32mQbNZJSgNXWWqPtJ2HKDK
mQmd00Jg60H73Mjy4Ukdnl5SIc+IUd6TgcXu77wRW/uh3adEYMSNv/Mib3dTNMPpY7lA88JmYaH2
GKM5u1eGT5rQjkWXzUhLJS+of04jZKBgZg3pt2p5JsBXl4xIXvRoKQ8Iy/NUXlPFU4Koqy9Ltqm8
6y5s4ho8OgTpcPZpkvIraMCUf0+s/barVGsr57FFgu4n/lVk2bdv+iZkFQbXdp3GJqrLJk5qUS+u
RQUd+tktMV28rJfIklw2fXbos/bNK+Ng7nvEAt0xit3UEZ89eG5DMtry77kdjCN3fZ8d1V4OtjZY
MSr+mB7mYOfVrUo+aBMi4lpQj6v7PfE9Si7EOYP9P0/iFahNg83ZTeKu6FhIzbBsV3a5p8TUorvT
23dA60BRleZppGtbdZYpmQ9Wz5UjDI3k4jZOJZsTTsrhaWuTzAQU+gS82K+Q2Lky+69ofugLE4dZ
90dLkfu7JEJ1x984wkHDeTo6bAFzaxgJDrrzsjfxB0HwueTWoV4C5iLIWMn4hItAAPulOBsGzP05
wkpKJLpI53F2j1FOdRIpHmvmiGNm8VOGH7zscw/AegUBexMlXJXLzGkNNomQoEuDChPncMgif8Cu
NQephsyhhZmumEIb7ZVS6mKn4fj/LUFikBQXjKap42F3DX6+0ZHh1DCKbxep7gCzfxyI7rm8/NII
vbufLzb2lW0IHA8ikTjyrweAzEyb9Gij+OssocSCDvyKJkB4JZ8Z6HqSoeJn+gQiBKXGpTY4PExa
5vOj5Tr1k43hEBLYfcRFmir6eISttEcI5xh159+pLNfWqzFaLQP/CuIlxDcxVtuDIhP2ToPS8hM3
kJQzt3GgKepnS6rLtT7EcKL5GHhEQxreoTVivX9yDcqYWbEXJcUeOwaH2M0Z3pFkf6xmFyNvIEaJ
fIP0CbYk0HeqhUUifJ/c6WVZSnUS4f9dgFGtdedp1TkAQInGuJE/dNeFjLurKDtJjwGJOe62yil0
s0rqqki8abO/VivVOsk/i5W/bZaJHwCb8mlkICwKnANWSDu/xmDJC0yeQFhV2ctz50nenSDmQqyp
T+VYlPmtvFI0wyEJKonX8P+czne8TlkEQ5KX0czR2CV7xWFs5/86EnyKc5BZFcPpYqdW4RXPKTh7
5oAPlMz0Hi/YWVuiSAteuyy+2WQcbxkkQYlf9Ys5w6ao4hvbLnqWuzpGiIzZQXfhBhnma8Mr6EMx
bpRKdm01xtrQDOTLIR+N+NoqNsYJdYmwBsTozZzngrdKG8O2YNVArGZmSMlmlf7RBAT6HmHdCJw4
NICRymSt2EkO89CcRjBi0WFWXlc6d9LkVVzyka/0boaC0rhqWGpNy0sWfOKOVP9BzldtqSXlsfoj
PG3YTfDmvqjSaAa8p/htdQh6hZCOOPTxrmpi3mrvn4xaR9MHKFaks+WdCTnahjH/i3E3Un9dpEKa
kt64PFpQh7D3p41pU1TYxZLbGNTjpku697W45EdR7WpVnh9cunuh1uAW5evDwodHi/+qxb7v7MgR
z0mPLLOfC50iEHdgbZ1BTKdruETFUbhwacL9pW6dY77ou4ual98RoT4P2WdDbCB/yp1r3VKIFI15
4YNAeTEzaHmcqZbZz4SSrTmXyax1D461Po+nmvkGtjJ1wLL76Fbrzlw//ymrfvXBSmD+cDehxq7T
lvZ0A6QZUNcqnEKMz/RYQWcKwWvLA2GAAZDa0lK/23MxU65VEIPsaw56BodqPEb+6ygYQfvlPqR3
zF+YpjWKyY5D6h8maKvdkav9VRzouuUOmkhGletXkUPA4zKeG0rwSpufD5GOcxzw35EnRG9U9q21
l8Pg+dXzzhEGaLYzuPZ0Wg3PkM7aI1y27y6LiRAeFCD7scrCFVIttFi7XB6mrEdGHH5+b5cqEEpq
tiyZkZa22BDhEJtoC1aCMypKyQRYO9+q9e6JV+sPYAejhgMhhBWfz6yVjugScoftZb2P99mkoAfb
4R3n5AVa2Di1JuCVX7mYE63JTCkWnHpVVqqYPy9x+ESFZHH+u5Wjknp/a46uclIjRMKXWFP2Q0nt
BJjnuudNETkLJ2lYsfCccQM0oFTqyDPT7UQv20bW3WbHIWwe4XcLV6guZJU5Yt4+IiYCcR+vpHAn
NCXDG8kx1JQuHBlclETph881ovugSdND2ZZE3y5SNzprolgC4yF/HUpFQTvEcB2xyq7QnZw35Tov
zXKXWVYfd3YYlEpyjQtXx4/hSQ6F5XMY10s469wAcjHURFSbqZ+DG5teHxp8Q3dxvQsZyCHvE3vH
ydF9FgLtta1/GvDrJ08/lxkpr+EQRPT9xju01qdoZEc8Lc3X0ypoiJz98NFQWpuHGPzIMvVewWUR
O/2x9XnkjSXDYvObe7w/nGUVgX0EA2YfCVCC1w7RnUpSnluNBJE1s70GMvNQd5S97SqmYYrqUwmx
vuhYULDoVZ0VZDDIKdYQ1vEwXBvusfBdgPNkiu2zIXhxOtfXNmBtmcR0nkADMGWvnHwAiBdVgefT
2ZoqtJC/H7seu50DEhpxYwXFr3l1+EGlaFQ2uVJ7rlT470RO9LbBuVRcLGCidQS++yNTyt/A1MTC
elvFI6zXbn3tAE/Hd+hf0Omm4PqdmVCSPzbX4VcJ2Y2E8UPHO5Ka+070t8BStoTes6QZY0lLmCZu
FaKzgpmfLbh3VsUWYjFmh2ilJJMyrISt3nO/sHuROu0vHD9AAtuTDHWk5QYh9vkTK3wGBXnBQClf
eCGYjJa7FD5Zt+r/TroOdg6PLw8+ENaZ7tJPn0BdcpcZpfZsUyweNnUonVwPGcKo3NC0D5fGBq9B
4GIup/uqX5/Lo4IoWH/jBBfb/h97JdxOx1swVaTTrYOMGIyFt5DZgcYXlS+YI9glJo/fD/QoHysv
GfeYyLba/i4KgnRIpTY3j6k1Y/bVMMgKI5NkTpVEx2biOQgW+77G+fCu81bf3HwZzZ4EbEkXSiiB
s4Iq25Iohp4ftJUxvv6l/Nhk8GTuW1lyvTCIaiZCZ6OmITqzVdlyfECnCfkE62Q50p8RzPjP8mEt
y2azGo4ZPX9MHjBi+FIuUHuQwL2pt3/sRLTRkiUZBfnbSNqs9NySZEO5B0GLIrFaGslcyToN85MD
kigwLPz3oCfNUJLNtxelGZNj6jW9Sx54UHULgsmINUkp+P1xWpWdIsWkWKmx0jql0iILKE5S5/4d
bEeJL0dXuFI1NkHHN6QGaUyrQc8QPJlvk/ejZ/SE0zPjFgOwmoWFIiiOwZPcq5AFBaxDhSWTGKiz
6Jn6IuMIJu7CF1cDHM4njuzdylX6Ia+VYtfl/ikUkWsLWi/819l0DNjxjkHH7nApVek47uA801z5
HjNArVuQJSndD1i8shLMSnEHLx2hywmnd1YJws322kxHWEuwTH+vyfppk6hrT6AQDnarFaaVbgr5
vCtiP56W6Fvu4gpi8iGTEAM4rQkM/DaqQqgyahAjRP/QG0Y81oahXHOsy79gZsRGvY97INXOmDoH
/IbhNdGcSMqr4gixA0NHndfQBmXjQ9tS03YoIBFNqooPCAx1SCsPW6LxSaZaWR1z9PaW9yIoU19Y
nxf6XZt5UVn4XfZvj2tceHUYxu53bxqOyhov/ts1IqM6e7qvNjv5lvXXe7A2TMiZf4H1Ug/S/3oP
MKx/qkkVUbMNyjGaf9pFoD6NdBiJT2AZVhVSag7rnuY+X04HWR+T/D/WRZ5QO7xV1NKsg4moiiyE
EesRj+oM/KXViJBVXVpbZII08pt2b2pPDNubgpbpmrZ0uKNZ4Zn1Z9RIooXJ6BHC308NTPYcE3KD
Fcxoy1u7w1Kgm724/GGFrtcgL3lPwgg8lTO5+0KWkvEV22asRf+RG34HysiprTfqlkLb0Vi0Pa+3
7g7JJ42Va4E3Ytm7j3GXe+T9skho7jE79y91Cx22gBkmFDGxQYBYG1mhWCuAgCrWp+Uu+92qp4+d
vi4TBLlgHGeJA2gpLZXdjq9rJ4NKKnbwnwBxqFeDtAEEL+g2daYaJ7nERGTwuWxnfaAN8vps1Qob
NE6pGcwhXZhG7bBRM6ZX1gQJOCyKvUO2Qyw07NyuJ5xFujS4V65yh1g0TyGezOU+yK/Tci/o6P/w
MWMnwjpgHS5bjyKvSrKqV67+KQ0zA5b4zJfWKzJUD8soquhmM7/jVM+VqqDCFenutzfOCwXCdExl
ElIuO/HzzE9Wv1rCQsZagBc20Qlxy93vZ2FUXHbgejhvaJawoSg61n5pTF8U5wkPVPZ1+VJKB2Tm
TAd6sdFQfYwTOPVVPtptw6GQXnCBGMMZ6xU4RJll7+ChuvNMrdKyuRuR4KLjMzcTz20ki9KKDQKD
MFApu3Er5vj/on13Ok10QemnsWiOdsNOHnP0xXSbauRDBdGm7mB5p3f9WKnIpxS34sOs9re35Q6A
39jA/QXjt3CBWtAT5PcEnfXgNTCE69Dk7OrpRHBiXxIaJXpkZ3sybZs9Yd2/7Iv1qXueN+CGMWt4
4be0TUSzb4OqpH5HniOPEmd1eTqAfm5ZbeHuO4LvZQYEKZM2ONM2JpRubdNYsg29ag6cVyaD+/xN
V8oTIJgEVYbPOiNhPnVeTO2DovXNZceNQmgx8T5zYdZEomiu3cvDDCoCiJPUExyY/52R86aC1d8+
pHUzwJdBQ9SaPZJi6WbtSvNIFKxfzTabhmevwQ0y+sTlkMAkFYOvLwKvCVkLrkq3xPaMED7c+LQk
QLveXhLZkDx+9am2mEWPJTmV3TaF/qfh979KOtTOne+JeR/QUqMguo5vlDAunhKOM3wJMJokBq0t
W6he1CygKi3eZ5b/sTj0/iSzhhhmi3LZBvppZdlNgf0SzPFRkDz5yunMMw64jre2hD/whYVgqNMR
RBDoLDTepdQabWcDNyyIm74hpskL/iNhKYQhGvAMoCXA7najXNlV/bH+Ak4bkdl4kuYZxP8AuqHX
hb8vcI90J0TgsJq9Xvy/xXGD9R2rld6MLKpF7gixBdX1xxR4i3/KLnnxg2XO2TnkhiHt1TSGfZed
FLODgp7skCc27g/6R9bv7ua4GHLh6NELNr13tuJkEizgti0f+u1HIJF36xpgSN/LN1dPRM8M0dRe
xRoIZD7QsfsZ2dHbljLJwQ0EXbaLNkmYYkhkDFdKshbtreQT9A+6dTpksmTtsyrgotnsfQueHT+k
boVom110jHMp+R6t2wF2JgYIXt3XnJhIZPwI6rZet+BCSi3MojrjUI8t/+efCuBTY+1Fn+C2jfTl
5LZruKAYEBNBk41Ss8Yy9RB605URsGfzVd9cQ7opt+Iznj0GfpQCq5zHUST8/jzuotHkslW7ag9d
+NrPNsyBEETn+aGZ8mUNGSAmcdH4u83TlK3QkIgdScg4qzacsjPBowh28E/UEuQaBVtXr+4Ahjjx
PH0oogGdjjtAgFiS4SBgn8EhAl5F21ODdMz7Apl5GN3S/hLFr7XIteNW/91fNWW8eh9axrAaoP5Z
VWXBLWRY87gnutianPFobbxo0O5vx4GBq+ys9RWn35Ey7RMd7tMTS2FCBYJ+4sAsZaQQn1yC+KrO
chJZ9Dd0695bsKsQrzpkhpc+J//D8ou6POD6YPugKceGO8QMDgVMocByhZE5cSYNLgJkLYzaSbyi
R1UNvPeg2ds09FRhdi140PcP1ja6x0XJK4ONxlkRCk2jhkpduMzLUZg+vYGboMceM86eY9AT1Xva
l0u75l1xYss8ZHpm2FJJnUJRHk3oF64aE6U1m9Y9XZa8nmAFrTELq02VzNd1Etl2eYMoxxu0c0HX
PR1cBXTu6JjXjJpnl5owaMmywCUSy5bijfCfPyeDlV/SLOartOm7C6uW+PTqb3i8VtOH59aTRaHZ
ok8yyNvPAkum7QXVQUxmXSAMwdk+5S5COB3C7rqyPsVUC9qowas+pskNun31xGZNOVbxhXnRxiCo
lI0eAZiVbrUKKaePOkdY7CsCx8m/qYrcSFDw51yRn8UvcMo6GI/fASraKFV7Nd7hQanEaGtUYjNL
REbqyHkwuipzqioQvTMiLuD5w062ya1REAxOMCd6mD+GqGA6WzPUucboJiFxssV7tbt8OJhmVweO
Nl9/LNg2xrCiqdNijofMTlJ3a7kq5zxdxNsbb+rzN0IMatLFfiygltsz30hmynKs6Im69PVit8cn
eU0wWI2wur5n5lOatUspG+aHpwFUszo7asdN8fpHcp8ZVDTlnmeOgroHRNU0uwCuXd48kBsdFs5H
fF7njyhImOOnhtB9+7T2ok0nVhPLVM2TDI+v/X8GUAzGlBtF2UQsUsKFBzi2shF1sWoL1CjEKN1L
bVT2J9RSU3KPSSs7DUiMvTEi+qoWPlQU62riBH77l5oWvgRwuuVOWdqBFfjzJ/XaMYVjHFClCmc9
BUvv3UZ7bknDCukkds3FI//0j4vp61uIMgf/gBgS+MFkYpO4ap+QfdNpfd0Nhpqunby6JZ+oEMCY
AHj1tegqrG6e9O279NLvNnzMhnWiSyx7HbLSxErGsIt/gVrJMsAlAJ/5A8+WFmKoYnUulpwTbM7P
4pRnCv4iUybBqHiaoM3T3vFodh7P0Evg/QwqGN+RftN3abu7aRBu32iaiSiL4S6N9Es=
`pragma protect end_protected
