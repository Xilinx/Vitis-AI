`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cpmLTnckjJLm/GJhnEEySb5724
XCmSymMTLlXyajuUkv+nefl4yXy9x2yAhXfBlAkKJiYo+BnqQEh1UNkLqYAA87d8AoAB9ihUb8s1
IgM+IoyPR9o3uY+NiwUbJmA8+WWguyhwiuI5cBoSnntNWESoTGk94tPn9TbimmCK7vJ2fB8ppcY0
dzN/XzQx6rnja2k1n9Vpi5cSISAq+208kK6K/eOIeE3s7kpYpnZ1FcABWMhBsWlFy9vQNq77DLCH
vQTfr5t2/fOK+lVCAVE1F3ghZ/HDrgMng6H2d949ESavHMLEcIAfSvCkJ3naupks8GlL+GMtS0rL
JRcPZJqM74zFjP+xERKiRsZT0gU89d88IDIj4HLpbgHcgBNdosusg5p1YDGWugARAUFCHHIJSzm0
E+V/NLnskNQ4y7r1+JGnfZgeM9dak5q1rfCU07bzEEa+NQg3jdHZ/gSoV6puqkcmbUKKNEfzXdE4
mjSN5mYMHwMtwqS8gM/epnXExMZm9RdksZ6K8SVCqctftG9EXVT6qJdGnALnziFpkJhWVwEYzqIW
XeFoWB8B3qkxzQLRW6ap2ye4yvytMnzvChQMbbTteM78KIEBUtXiseMbhMg/RKDjS+d8Zwc/A/OV
IM79DrPPTzfP34Vvhod9TujdIMSZ9tGtpzwYi1VsG1O0wyy4pSowb7sUWPzZ6/CPBabeFTLccTUx
UzSJhafqTl+ecsulPWedZ/pgv/j3Jsoxs/G5XBywVnJlIM3N/CDDIvEgsSo38+LPjahCl3//5kxX
au8pFm9MvPL47WkbETiUNjG6DAGVmVkQwp9sA+faHBMjVhBDpTA7iCi6q8glNGLNooe9f7Uy62Px
6WhH3nqyhLOzLyInYqprI6PtmW/kqCFY6Tfy6t+3uRxfFVWta4KJjTQZfPk08AHLXO5mdD5F8HTG
XcARm+uQCRP3whgQ46cYuDyCt065gkb17Ek6W5Th7ftg1nObs9bDzjDRRg8FfyHAiegpus06Hm9+
qQZ8TtWMkjyGiYx3BG42xsFi+fZCoRR1YnZ4ouIk7LtV958hlwzgWmcWRn1CzDlebOClPFd0i1Us
imxiJdVUguXLte1GfJY4vW35/S+r56QNy2+5MUADgsJu7LS12w44urZMbUWbnXSaWnd7v3k/ltU8
eSR3QgHPFM0psS2L1vCx4/uB5LKHrqWNzv/fv03fUn0diMh7aeZceifnbhogPME+NbgwngZ7MCeB
aNFsR+ZN4JW7sK26GdZfotqY39MIQmNut1bSK8smHkEbGy7PY9nL1I2kMW9Z0Lm8T14IpZx5D4QX
Fmb5xoMen9yV96v+SaUJje1oA6rUVWb7JE4Feyv/EeFnnhE0qaF8QQ1WX1MgSxCD+PvlTiuy+8sH
LvYMjmsHFb7TyazXqNhUhVlcFxeB83/cVD7irhS+TAejpMr9S+W+n2+n5Qrb7dAhOPhFxhnf8hg4
aSxIZw9qtDtiM3piBwlJDVCi9/xyon/y+vy9g2hgL7/6UzObBSGLQZ6cH1gmIEI1WGCW3m8a+DkL
nc/0ttedZjplnr13j7OnAY8htL+Pa7uTv0rFBh1kB25pQN0x21vG+Vftm0rGMUE/V44Azsrs3JEE
pawbd2QrM/OnrbSFBxyXfgUF9l+B7nvBpnrplr0gM+WAAxJgx+FAaBySK5qsUT1egBlTCSyexvuJ
K8tWM/Q2pEZSe3sh9tCaSKd9Ac4C8cmC45xVfMhCS5RiNNwFBibqGOJI4rs8NppoDGFeJlqTwDuR
KN722Ecx4QQQI3WxlTQ7MO8EubExjzDg44+vhiPj8BKoD9XPlfSg0pslwXb2eWi3Y1xKKzz5RZxx
lg/AWLm3rKnO7jisqlsaSRDQvw0oguPId0lRFz34yJFkGjqcGUvQe0CtiWs5VcQlb6FdaOBE4d4a
PfnJWcaYhHQ2zAOrUN0OGfiynNVeXzDi5bBrdcRVPi8jUOyR+JtzZahSeSWyHC1jgEYjZAW0hIeC
fuRvy1hL7sjxBRyylN03WCiPrHtw4ZCfNjUSsu/FVkwzxORoxT1YMyUhL9yfX+vg/qGWJcHj3Y63
A0v8xqUyOKEHDsGtA53jKJbGQy9aN3xLEahuM+TL4fxkZVbFXKqikseNasirqrdkhR8q/sKGtAGf
/ah8SGFe0ije+q+0Wd97iAzjMcwcqbDXuL91cvNfs7VhvcjQkpY18M8o5hgDLOfiHxgv/T+Q9ysG
r1e54k2UGlOkFcBLFn1qqj+zWSYoMplE1aZOIMylY1NcMBLHtuOfSrEcs+lpr/KQGPhqG0gYRnMD
UYoau2v028ZaaT/TMTruEviOlhGyoXiLj3IBxJnmdEhIaUL5SqZttGJtw1yzHVa7hdbAu2nlAQDO
hkGwu+y5hOCOmQ4Sc8LyauM3z2C89EfznAXlJJOwEKGNR6N4pHLJQSj5robpdwySXJVTZU7oVRA8
/vH7XjRLScwvVYl7lFbXli+WLAtv8E6Mo/ubJeET0G8KBF80Ccb1M9WvQYOX1S7SEaz3n28e5VHy
JYlxI88Yb9Nq2YB2iVjlmjKQIdK7E3HRi65mbFVXVqi30WGAD+f6vO4PLBf5Zvz+cRrRkCi+38yq
IYQN96+xcIfw0r5VMz82HGaIzForI0XKT9hkQpMMTBhDHWEwPNqyVOBEMTFMFdaYE+LbNRrkSkJs
YwAWspVpmAb3NopMgdd1sRZutOAQTrDOZIxA+Tm6XMLnoyZZoLqdssE29K3om0OlLiYD08npsxEw
IwrEjO893lGIhT0gEMktZ1uma71K8bGLrR4RzvqUqlUbOfzsYP9UApNSA+sqBH0nscSroNgc+62g
ftqdMgf9Uh2HB8Q4pxH4LZ/IfJ6wQZdyluaxQbw+Uomk0q9prDsxxs69b6VoETxZsxiVyEmwoKcs
aJRavuJRdiQPihoijKtatmoOtTIqyouT3p9YAYMTscNXyuxinLl2kXvv7ex/dnKTLz9gSRpt4OlZ
f+3pXe0w3yCAZu0zaA9/7sP6ewOv+lkFxQ7gPrOtXb5/jBPrYO6uxPMkwSMuDgDdMdSM+DNIIG+L
iB+qHh2HAEIBTGKZul5c5vqHXIXJpH/Ky5xCFYCgBpO16X1mo6Srn/LfVYS80clEeUGEZzw4fZgg
gNnsuT5EVxgQutn1OoAby4ykF0u1JVHSKV1QNwRWiBcwx54IaDlsA7ztnCKzZLnzqFJ7xh7mE0ZJ
0nktB4xo8uYEUBBcUV1riPt+E4hB1UedSdapFPjJlrS84qWhLPLtzvzhy1QtokXbq9v2XGjuJUu/
ZZrmBdI7gLdlrxf2TI8UMtpgBf9YYlBKcUVPn9VA1N6cbvcxvytZT7t9pHzdfEyuGFOlWA7U3u1v
OSoRTD+IaB+oE8FaAANx0h72sTPx7HnTmzXQSFD/Q1JXpYwmjYj2GFfQeOFEj44habIKXefP9FaZ
zMjZcpgaH83IQVS88hjMN7PZ420iR5wEvaCRJiowxYb7tXhZd9HDMNeuy+95IQAEJOXvgMN1PPki
9fzN5XW9ibptGT7/Y5FLt0fYRzoINkzDrilcQTsDqEJ6rDh3whAzdn0DbKe0Y743rFK7bkGDMCJS
nQGtgXVZA3IzF6N8vzoiNa7V+9DeSQbG18dj4pGO5CC5eMK0SdL/0CTnumG47CW3LSOpposS4cVa
JBzFLSnCifLZ6q2fjKWSwjGh2t7Jb8fPkYunbn+ZJcpNou22CABa9bznCJs+3+A0xHlTK7pxwCoY
usrYyFlalnXOIC2vvBvxZO24bQYxI2/rGcVXL43P5YCgMprwZ58PAwMjMNEqiJhqXVTdKuup6I9l
UuFIAVESRGuYpRuoWsazyMFWp4GgrctA3i5YAufSqOLEswvzvTyBE5xm5HbunW1AkhDni/IjEp7B
MBU2zXFEZNXX4OgWzdtFOgXpVlQYfZGcBIUZBI8MEVtTwz8eSWHmgj3oXd+kvpKWvY5sw165b/RP
JsCrcNNDBCmu7kDT3vH1c7dcxnfElFW9UPM3AEaC3zfoK51jstIb7U1sG6pIH0+/OIcgWyH264lI
WiA73W4GO8S8HqweynKDu0GS5M5weREKnkIqmhFFzVfXUll1MZtsTfzly7lVvgshiSLM2ZBdoexd
N3YqLgRupJGD1XWdxpcizf2HHp627kXot4ybykQ4GLN8cb69RAp4W9FP6f9kMNoFn34yLG+8CSkf
wpMfArmCIPbEw2C4zolhqwBzHoDItlI01TKjbxJcas+B2DXUlvueSMun7Pw91OOW2u0ga2cx/1fp
mVMydqmZtKkxw+cCQ468fLn5P2yo+LiSl3S8prPUTsQ9D5OskU0ILpZXtf6/eVyCtkvMi6W7DRIf
peLuuPJCsn44Veevonjdt5LVhSjiNexHC5IVan/2HWUlYhDHXT5+G4XQy/9SmlgqX9TCyVrtBSQx
odDbIDMa1xR5bLsf/ahiaROx6LSBed3KqwY4HAumWpzJVNJqQQsxwyTGM3e4oVj88BUDl9IRVtz4
h+7U5DYl644RXpPaBUIduBVwLSoOM6dCLOcVZRBBfYwW05HhxIuxnsmOh2uh5U+4wJoO2I/TNsDu
Kiv57HgytQPentKuifvAFYY4wSLJJmDN6d7iGa60WpepS/Z9ip9pf0scSM6CXrlzMG5UawxcCJiO
60cuubBOY+F6BaVEaWagddY7Q/5R2YNwGhewPZr5fab9OII1kBVnnuEHxTDDlmq41VImuF7GrXwt
lAB38QxLsOjI1OfFI7NAtUj6SpemLKZTtwXUVupRJn/UkSZ2bKatH7RwfJij/qeUtsaBbUXsc9Mw
j3x/wcgIkjeqZm9M4FJVMofz3qopZFUVgGPFHwePkWRS3rvuoUx5kBwe4zR2SfRH/fKwVdsglmOS
l3J4Dp7qcJnLi7mPsQiefvRUQL24eRblSJTHlwIAHF8FAIE1YwPWsRuuzz8bxc7UotrWrqvQkxO3
YaraiWqjjMCzLLYrjsvymCLwikb5Fvb79tYi5FC8B5plfKc/4ouYcuoUwgTjPv1/Nmj6BnMB1/9K
tpjvQrDuJxI7CE/D1enhEjfFbJvUW8vLTfx+tlzn+e2jIS6yOCAWXQEWNRUYzCg9YFaN2SvFWMSB
F2RhV2RFQ+iIG5EUxQc0zlEMVphv7VQDHD8lgFZer4XyyNHCStJ7mIv6aw99BC8G8hBiy9PFSU6r
Js3F/JCxQfcU0WxYSA+be4Mizl/COvimdzGvsbg+SEkgg5WlOlihSiK7xoEjK+E7hyV5//jmaO97
xL9oCQiRhm6okytkn6Xq4GvZuTcpKcckIj2UxZ745gJMbQK2Gux5xZ0YVMsUi2VnmN8GVRfJLLQV
PN/zSzdfMchwffzOJqTax4uI/SRx+lcv/XeoDOgWdg0Tr+lCoQFYveh/zynKGBhaNJ9OyaedXfim
I7wBEAS9BXncgRljOD58CAtXw38TO89UjbF602miLj6Dx0XZccDnlpL+3iJb66OBGFaS07HtcZRX
rACWS77zOagi9fmc3O+9rs9KU5dnXu0QbqKA+Z6xgNaPQvVhbAQ27MRatRtHfAv60IQWswinyp/5
kq0KPKETID/ohJ0xx9lKp0902kABEMQhIm20lDmqBBntke38QSvFFX/AxG10KZSiXgJXJgtOBb2H
C4sgzCFx/8pODAjrsSTBaL+b4UQ6y2jwA6EZj+j243sDLvmiL+xurmNt05TOXR954NdYIWn2IzzY
9ZoGpp0OpAg3MQuLGkwFPPmMNET5tP85dvzR4JE+6PbxwOBG/Q97kfyadofkKUv4Kn6UcMct+5wE
oqZK930OMwxecFqw/G2sh9pRcWSAf1IT41pZ+kXdJzhXxLgV/ZUl/vZWtQ7iIHKgK6sX4OI3MVoJ
KJk8e9J1LrEBP9cKno9rnpq/RztqEUY9fvK2+pZQVxMOu3Swzbu87y/+2dIj1+rcbjNl0dT4/Lzf
2GL1l1xukqWARkZc8h6Xo+v9kG384q9v9qXZWOsdTZgTMcqWGoM9z69qdLXRhOCG1M95harAXZDw
jPbJABY7yHZhvzkaW5imBtHqy4A7Tkpsnw6S4Jbt13LHj6fMI8B9PPAjkG2fbv1UEuS4uMNBTme0
bmjaRsOeZAfrNC2SxpMFclXRvpA9/GFNciIdBlv+fbhbZDk3u/JN0j/TMahdicJvQVbqZMswhT0K
mzaUF/Y39SFnWnaIvlo0oK3npr8/7yq47yPbLDoXAGJQDnUNwPlLmZfJLLQz4H7/Y6RxgrOgd4UA
T2wuo/8JRHde/iRIUb3482XA0s4oK++wJ6w9pWkP16zO6J0lzqSuFfnDrCxvZ++auF3MNXmJU2Xq
gc02qvB/zh1MWs6sJgw3ALy0T3uFc/XAVAi1cJ95YZyO8VMWWxpZ6lHqEHE4Zt4Qr7DiyHOgrEKU
FcZz47Znsxsww0oki9tiIfWsZSF1fj/wok+BSEn+tdol+camPHgy+52S0fcc5pzgIEaWssauDj2g
edR/ypL/y1OrkfwX3EOuH33MLSHlrVLu8fYeoMFBsE/4UptwttU4Q27q63hVUUKq202OTfwRuJRu
ACflNz59PBTyhRmmLa8Qd8ZPNUxRVIN2PbHLxj36S63JSk+jfgIKenMSzocL7xKMuYwQcwgNyJnh
63P8Bs423YKpaGG5aQUQZao2DXoMCvOGDEID6XATYD6SNlvInW2dIrlyRRjcIso8hxXrEOEkOJaU
vzOE7OOYdGOb/LhX/PSOQq0iRVgkY9yX6Lz0DYkc+tkL7uL9BWEoZY8CIarMbapobHXjB8f5Z0Zh
M3RCx11tzC+gRfuQMT6oofzTG9nU3f5jdPYhvl+0FKBOYr2p5gPPgtvs9q0ZgYYXbybmD+WBmZJq
F8UGrHUmQ4qaFuEPV2RPYiKZOaiLHCO273XJsE+X5UFp62RMUtUKLuaA8N7G8OqwRQf/2zchlzqy
vvAXWH9pJu8tUhYPjtP3iMacxdojrydblV4hIdDFhRWwKQQwapgBz+MVwvEcDHG/f8J2KXROXttR
69YYYZhhWSnZNO9RpCsi3zcEDRbXRCx5XGZ2sItf/ZjHs4mTxmgO7aezQUslkjvTq3ChueTY8BqR
FXivqi9tNpUch3EYkU7U0Cn/18UjkOZ6eubeZWcdKPOizdXS5wR6XzJKXjVhYGfEf5hjjP4MnJov
DDqGbxhbsWukI254WtSSuBRm8kL+bzsQaxGdZY+f5j06htoPsAqU4UcB2e/KU8mAUJvkYtkcJ+9W
FHqwkAgNYW57+qHJuZT6neLS/1b7dDZAHPlah7xtxN1myDy/TwpqmKYeXMppnGj50J43fEUKEAaB
OeNcyAEVGSrq0vKJBSof3tIrVrc1eQY74tcyRJGt/SUNfQRl3/UniSPd1F2YQ9MN3zDDbual/DF8
Maixq6aSQWYLweTLCdcIm9Ic3g7ue0hroh+mus3jmr0Y0vZ7KJ0xRmbfWOVOVrn5A3HF2VReQIcf
uukewvL0mXVSLSbgbsTNcu9V96QSb1Gm9FnEtUSoZ4/OypfOyttzG2pKHGN5/DZmILnrnJi3FpWx
BePQYZ8F+dj9ftCXcphgbvJXG+1kTeFFZlOk+jO/91L6iycymYZIZmoBbSkaTUqZK5YP3kl8OKs+
zoP3VkiQY9jiloNEotUGwq/+OTNM2Ndk9DHSvW3Fh9wUjxResTZAzV0IvIFa+OQb7kBOSz/djA29
JjjrFRWVXUYryNoH0DnQ4vKp9E8iPkObve3P44MC5LAV0uxXxwxltPDsc1fOcTnCI8sJCYqoNhZC
At727AIuXIct91TFnfTqJcXQkIKoomeNduoxiJU53eX65jPVfrKqKEEtkVF1HdxZsC5N1D/ZOgjq
OEMrxFp6kuDOh9M+8vau2+clazSbaH5Uhi4ATW3X2kKt17qI5bYSeoX4FsWBy1SEgRUAj7LKOTqc
XEjFmdzzKnz7LKvdh55FWUJhcIv8GWBKxCLyVStQpH2kztwGXxpaMfTQomzxB83u7GIFgjtrdFto
dYV79fcp+7Btwt1y+W4oywB/McjAb7PFl55YsSV9hG5dwgBuJARCavC40rMnckcnMTnRZ1Iy5Lfs
h4LI1a2tbUG2ROSdd3vvChh+kt+5XLGXTCo2G3UzIoRcHVr05oe7dqN6tca7eRAdIoMhQ3bh9KyS
EE5nJveyDvzDTVM1i9YLv8OpHst5vxp17z9csBmhxRfNaxvQXlvM40zSgwmw2TzaaIdeO8wXapys
BOclMPwzCI9cvBYsh67DOx/7jgfZTWazou5bXKqKjOqnNXW2silDtWVinLHw3VB41rSqmQLRnQ/j
D0Fe3qn/YBvjIKn4MLEmdJykg2vn1+RHZRvEDC19ZcH2O04ffk+eT0tMQVvMPxjVYh/4uuP/Dr9p
MrKkwbKY4/CBnCtdE9fybTt48FfrEqItUECNkJC55msbBnWABDusnlIuJA0YRxJO1GRaGh+drglF
64PijDLnA90bK2I6ruvNaFIetYNzGvSEOFg/fRAzsZfClHANg4b4cslFvRxnNNWi7Xn0/d8fwtHR
TpBDhcZYwkPvCTfk6bwL4qOeSUvQnMI/J4Tgo8mvJ27JJGGW88ZyYN5vEmcRtgyHwN8lWs89B0R9
HaP+bhIXp3ahKc8OF7HVWk5ZYxkeWqYH2nYGuQACz6GSqXsSHnOJbiU6SSRyr12WSEgzWaEzDOn2
sL6ArB1VCR35JTGmBeuBLQ2e7ffRYiZlJt6IfFiOXE60a/vfNJR8WkGOSHf9AlR/HELcwL9O5TQp
kpInPCZJRcJRONO3ehqbNVCT3gePm24wA6P+zAzogGLDsRgkZdvpMc0lCkm+CpHglaWXqtI5wUOM
28r+rNk3xICFDwrgroEZo3FFV0DYyUB3ZuJzIZf+ZdVp3UeOSmcMPCFIQOY3X+Q5U6iexVF3UAWh
zgAMHCe0uSoeNLnGoERsrghaJvp8qSkezjswD5fBWxgqfElHvQ1E6fs80WkHBPXErxkwcyEpTaNN
2LJk9xPyAuAu92u9XqG2KlUfAfrsFejye4TMU0Q4z0CSt2R4TbncXxO7SStMTW4YayjIPuZAFvQF
zDcTxiDKtS/+Y3T0OnPsIKUZHfyLmSNIQoUaO3tgLJqhtTMPd+5AkPU13civbY4Xgoyr3cWcKsnE
74nrXjdKv+TzauvXpNQY+H1yA8dcuGQIv8uM1wEeZ1hveCoqtK0wyZ3R7OIIihUT4w49WEQjY3UM
bxLx3IRwDGwZ72NZo7IIJX3JI0UTGP2yD/WK4Bscn27Scn8Hq1PJx5HW0XoSxdbxmoG6IDY5w0CO
M329Ja5kzIdFVEbeFgkVu/M6eARmlAEmxUIk2h/u4A4nBAjoZKA3PNvxAuG/jgvJFYVCKb5pSEJv
OIz+fKaOOhqiRh2KbelHIMIxfHGVPgBumS4/ZzAMN1yELP6vOnHviEcKnwr5cstiIMlOPTwnv62l
sAaCz63O9ils/COem1b4z6Kmitg9LUo8gGHnhmaUoyXj2NhCiYywv0iUJMdbpzbQWVcpKQ4NIkXy
dSCJ0M8HxwZtSjU89zsN0qD8bgcaJkrGd2gJbHxhGJmDeFLdtJ2FgNR0CztpLU/0ilnnzKPfuJGx
yrwNhLaD265eUjEdMvtBl+gCrzcDjB1NnQ+RAiuUm4QJMPiuH9CxtETQQYoJmDJFWsvQo5Deh2RP
uQBSl0PmIL8x3wfS2iOi91bF7l8M9WDF8/MjotZ/y9FENYMt0RoCvlby1fQyq7JXP+1tbJWF4PYW
rk8y4Wt8WD4nkBTT22AdTWyalCh4CVMqWi+W9IjK+/WXgmk2/xXKBdYBUCipwbcUhB4vUmCPB+6R
4y0PwVVKii1RE7VG8IXh3Rq5+QM6MV0bfPMVRzwyOkNvSo298RydISUSi5PqcWqVWGELKJRSWi01
m4aBC0aQMYy4So90Cvza2QsngycYwYM3G5MuGd6riwZRi10uL412gtDPzo8Do0OayF9atawEOaUd
Z4GBJJ8wg5noyk4cmHVcaWNoVCIja7aju+anB8oUEAweh+aud7a5dQ9RbV45ngBfMeQn2ILzE/E1
S56+Ggem7R1xcPG32mCBnLaPDgKgE4+htmIOid4+ZxqGva892e7GD0NWdXkO3novuLAA7rkMU7LK
I+hzLhAgEq+gqZt6J8u8AoNDr0zjwZrAf3hA74xhD0OAUM9SKgyc+pM9DzSnj9GErlaG2opSL5BG
EPQnkHPTIUs9pKWFOW3qkBImHt0JLBGpOOydNma9jGCcy+Nqv7PzHPXT7DrY+JACfAZPWlyvEYtk
P0O/SrzY16MF6UeCu66Xql2SQ1/eKhpscVsZjlSTj06JATYuApSv3CzqYxN8wJJtolE3HpiRahq5
MLoEFRiPSYSr+uBRRflmnZmvoZApwAeDz+FzYmtdD7rbqsnJ5HFxbEVWdlIe/SDhdJ1qvN3Y5bnr
Q5rbFOuPPan8AolPcxjx2/yJRbWzHIJGxAHPNhrAqo1tjgUlFU6dNgP76UX72e83KcA2toUAwlUV
/gTRrvItx1x3bFwb6JoVxuHOWaR64EjzVDkb7i1sfMOzQ+JSKJCMZJeobHlXgGx/6yaUsacko1xA
MuoveoU7w1WXBC5wOhkeFgKnQb2djYp3cqijDyw4TRPgFsNvQPxrQFAHYiuWv+s6seL5ETCO+lo3
aAAjSbt4/unzk5YDflqRcXGaM1MPXeyMvDv83/JXwG/Sm+3RIZxZhKDDJ5Y2oDo8zrqxfD3c3MpL
iEv7Xyp7SElil28opAJJ7Zp+y3+uyo67bFba8ga3lK3TK+Td55fCWl/OZxvq4YERI7764Vcgcxyf
R8HSy/oCMEWzcXhidcjdMo0fovzD8C6+B9vkCnkoQsCYGV3LAKr4ZGbLQXqflmk1q6F74L/m36RF
IT8jFgvD05p8BCAWKrd4E71SjyFJfLXdvaZ7fMTLhizhd2tqkQWgZM99cj4UWLsyAsMoLzIvO60V
v/qGDqfQoYWe7M5xb5hxX1E69uyOipiWpELNhl5pc5BSykdEBILKldheBiyNO0BI69xTg3g4CBvo
xlwma+kH+m+7Yn/B8c/bauiq3JiCJqw0C8P2WPdr9tyeLmyLGkQZHx3FhyEbzjl8Y7AGEp6iufXY
4ZPP2IyHkce2T+mKvpTXBL1obZFsnwEDvSrrPwwlLTxEugTuzqeMgH+Wn/Ohbx4DiDxCpqA2ek69
NelEHYMnCw8ltejeiXkJqdJugshR0sOBMhDDl5MBegQgSFRuZMNjiVucyWVDk49cMEQw051twyBU
ym2FNn80I2EwTX3qz2eMdBJUDR9six99UtFwdLnr5/FziVFUPcERUqbcuWLh1pVHev2xmE7AWMJL
0g5k2SQBIwtknd+OVJNweRXyLHvRyqyOZXxUYqWLwO3bg/Scb5cjan0vnROpP494GEyRb0b23R7C
dQjtDSgxiAjVT5OsYdU2BNzUPdwmaxr+70M6/XTRc+lkF94WwrvzW9/lQNgUplzcGoZfSdUDHDYH
QGHMDsj0YaOuhuxSZJWUTcQEKRrqF8esaqL2zd6DyQRnQgZ9xAWlbG/Nf13UjMvu/UKUo6uzkTR+
Rep2+go9hSU2KC4zPPhq1OKHhwbz1jw1sUhT1lK/pmEFiFqev1CK7RBPmuxRDr3sZCrc1KN0Rgj1
KrsF8y+5w/M1xfU0XfmlKDx7gE0/RwgtGWhmYRdCX7Arc/U4wkAmXCsV6PfEFmUkiqMlGnFUihxP
PxCs3yPC5OvzWBJZ2FwxyPL2iVAbO7NaXqYH0Z1EqnVVsk67jl44Qpqrh0S4DoK7QZC8lsC03BYA
xdMoyiCcJPmt3FsDa0M3+z5lsMglq9+JzNyG5r2SQj6j73lae+epReWfPez+CFElDB5MH1DC4VTn
+x99nLR97PawCebhBlWfHQ7N3c+mJCnQLT+bR5dLrapVXyhUJ28T7MUGoDZSvcKfut3shPXHfpda
5qZ1bcnMf4L+gLqhCSnRTa39Ftw3+t1Mef1B8A6cpP/6jWYwl66Z3sOL0VxS4EYsUHh4GAZkHY0x
1ydZ3QW4XwCJIei3TPuBarGvoWySp4XqICj8sMCkUcUB/ulujr2XP+peBn08xlFhwA8IxMSUcRfG
Jlnc/uy5Bvt09Ff12zLsGknYGQUXj2Od8UJRrwhPOuaiF+06wIG12mrCFRtec7WNLulJORDV8CDT
hywDUsWdKk3BdVEklgz0g7iDKXFRTNyI3yS9T49nlaBJPzXCTYklUqmvnXkD3wy/u2p41esCOM5r
kyz3KadU6c/7v+L2NxUxgMay7D2XlB+B87OJg8wVAgIZqNRSaKrXjg7gOW2OHmoMdZoza8n6SUQC
hl5LHzgmxwaGbeoGgMczvtHstxZiFnnIsvIt0WIOZBAMu3uzsolwDyNeYelz/h5emg4uy2wdRc3Z
k21L1VI5ZU3bfAREWBt80CITjnF7llVrpxF5Q1cc4+uyH3ImXEesjEsYanJuSv7o7OWBEMKcrgtL
F58Stu/+DQhcw9TohZ0eMiiK3hBUqVRDJIuECEYYXKp1GthmWzFpnoHdpT56Ujc+ycLKwx2or1Ug
yCJpL+m310I9MKunYZTCqGVmwUVI4gv78CunD59f/Nzc7/4lhXUloXHWktG+j+t9lEipgDRgQ0dr
XlvdfYAK+flyb4RKfiySy5kZPPCAtsF/XvqYGSN1HGORHP6ggmqaeLPwDWL+qJ7v5fhrSrcA9VTz
9TfptKtUkRLprCOajyiTwMXDdQh+7Kng++vMmUzlt/OFXJeRqrwiMbE1Ma6ZwrFMVtr5nSK/11St
lXncTN+PjrBcdrZN8g2CH7WhW1kZxDxn4RlASix59TCiGgsuykpV1/HHAs7uURCDkVhQ3mTEc7yC
mbJw4+ePy5uv73eFdnTnAgJh+7gMy7kOBE5YgcNuIGrWYBuLtScu69w43UM75MhlmpXpZ2fmRzJZ
h5GsySxfOxUGVd7h8t+AxbRNUIQztb7vuhxFqXIgsy4zg0HAyi3Y+yr9Dvp8W2ncc3ODq47EjmbL
C4jq1SIMdwi3JsxBc1aCTnk9fcg7kuBLDU9avDOt05ZfaYuEbxoHEEHPbshi1DA2Vh1N1Bg2CC2U
0UiWfKs86Ni6ANgW8wkbr5wzzXvPYzTQ0kDlG2v6rmqjGx9Q6QVpGicq+6ifVHn4llSFEIJpyKRL
BqaCG8j+c9WRCDkmG3iyXWghpPKBuMClR2aZTRD99/+pEBCOrg2SZbV8GYUAAdcsdBrMZIvdOBfY
qCxplmCbLmfmzEKBBsytCtFxpMEDSF1/25whPNuIu4UYjqWisuVUFKWbgEsBv5ekm1WHLy7dWAAJ
hQTVMeXSQY5YDzgf8++SrzUYH4kPvDvI8DB3zNtvpMBoPZwSW5laB/j3RyZQWAeb29A2EWLHVZi6
RRxofF8GVVhib7VD9nF/9gqF8Ck/a9aMudIzForXZCq7euIh/+Vwd4dasJiYxvL9t+y6R40fLkiR
0ffh5hUL/d0UVEHxD1N7tzXxOCeRul0uEQu6UJHKw5TUEhKzdHm4EXXmFHmMuEZqq5S0AFSnauEo
l7Q1R9QORPp03DUFs2ChHKAWH97UrFsS15cCM6WoQ79ESWcaDCbpG+wqSVVIVfHu2qhTOMTy7IDX
yCZUiVMmWUTo90ICnvc/0KWeFD/bfvjQEbpFZYsN+QcCnHcDz7xrqdOfZ7ljmPgcliQhlcl5JtgE
/tS72asX5Htt3h5hafoV//Z0DfRGq9ZhDqBr6qUbtIV8TqRwXjX3W0eOrCiiuPCHtPRRAIT2lW0M
7+DPBttrktVCHP7Q615/oFxUYK5eP7s2ie3GS0RA3eJP/xGyiR9R7BsTlLOAJT6P+m8KPEnkF2tD
GMScsshtlnPAfMcmQ6qWRiXZQrIZZa4S5k7Nxjdqb753VErwthesB74bvI3B2NuUWeQhP3sc2Ppn
5b+a18JzKsItqfjFowUd6a0CVIAqo6rXloyOyHC5cZAQlujPNojFBDXL9fwaFnkmGRpFLlO7+O45
RhI1LH85zpnjHz3vgQZ7gFLgjpg3avYiBAPro3BjCugoOs74x7ZpnkbTCf7cr87mUneCssNw3KfH
5Py1nHQzC/LiQh7Da2+6Tkfp8R8XPUgF40iAMSwnxXjJ8m7FKToqfErxJAnGEfE4y6mzGvOxVtNk
sf5lQTPpL6/4Bav9qb9q/oCPp5Pq2ccZD0+31MyyWYyIJBR2zX/5xhhyYwXp1dIvYFUkTKbqoAiw
J+7TTQjxc/V7n7E97TxKBfAPDN4bOGj4LYyS5TuXZVywksi6bUtf6Fakq6Jc8rebDiVu1YwEW7Nb
HHVfkxqBivoZhT01g1Fi3ZM2Kr0WqkrfaaJvS5AxqXRDddHYS1WtHWbOAiNnyReYfg51r26QbGHW
vLJVaoMb0HqoVNlo2hOfd0uuhOp5tmQQFwHoEU/z2qkpNoUaO8ACsNwT+yBvm/ksNdSau4zR8az7
K/m/ICYHSWn5ZhV6S06uZT5kJpWdsFHbGwhQ2Sl/04fPpMpfd8I7vAMT34SqZZXmdAahMwEeoUUN
HEE+v/Dhbsnuu+BNKENoXA6uqyHpTRse7h3I8elvYGOhkBD4omH3mdVcmUYuMv486v17bGSE5epB
YN9UHprHkhYEmmcN2xziuuEgisUV0XnkDTQ73CZhpoeMd9QwKT+h0oOL5E3OzsUUzO27mT523uEv
IrnKyybvrnNJ5pwg3vBbnSp8ABLd1gw9zPAA9NBQaP9JaJfzg/soE7gqxYhVxa0r+aw3LRyLWUQP
wRrYUZsBAfJr2a0OQV1lD8ru6dmRki1VexFab/YLsY6zRVl8hLKYDXMNDa+pJ60QJLfdhKBo9Q3p
k0wr7eLj1K8zTJXHNaT66atFDlbIHMumkNcBtatScMfbt33ordVW6WagDxcAqRsqKd+ea0W99i72
0lVIuovDBmdqtqrPcNNCy2EJaoqAmKtKgD1P5HAikijc7o054QqKjtodaSx50iD9XsOTbFFe31Lv
NqdQg3OogpK1GeV9MXQ9OOdPo3+g5gl0MkT75/Zf1Ti+z/uCJviOjGkzN0kILTsfHUftvaR5EoVm
RmF6zHzj4lb87Ea+IxHlaB/OrV5QXOJUFl4IgDcZY4KCY8Es2lFgE32AJUHAi8CO2EqlsVy5Oxyr
6sG/+bOEm06YtRNzC+8ODI8uoWkLOkFqQWBoVmHgVe51amtgiH5QxX2oDmHcNawLbUMh20ZAIf2g
t15OirtAPlauCX2tAVcQb7FwG/jzXNAK7/fbaIZ+Y+TNA944Zi6N2X0+k2c06QnUpx4bj0JRy0gQ
qRUEnPdA0cR5SioSnK59dXHTWzWZH6NpICqb6IripUYNE68//4Hr8UnVS7sj1VxLJbn8E8jSXy3I
6CfDsKROgXK9aMipj8PU3qjMQPhd4TERTIqOOLA7jHvvOjxUTtbiemRAXL3gk1YGELQ1EyOJmoYY
Dh5JiLhetV5dKRROWrNO4uuP9CWkKDJvk+AwIz0CTpSBBODyJCdtXnY6OyjQNzfXs+o7wezpCso6
oVTuxGOUfeJHZBgltOfTrhgnI9ClXb1kK5yoTGeZJyYnKE5rAZ8jFO0RaEeLNm4H3+S6n5EHoLDE
EvxIw186OfFBuBKUYNTxDNa0/eUTiNGUo/eKCDVqbU0NmyqWEe6wUOxSMMSXUN+qG6hTPQifKYbb
R0sx/ayOzkVCimC9TGtE+JRGdvA480CNVQ1a4r/XpoZjTK9r6ILic7+usURnWVtMMF+eMkfrEw1J
HjtzhObxOMPmOrr4V+CP5s1p1GikZpzD+sBpZoh95op8vbIAefit0Zt9EhP2xj5SjbwkXmklwZPl
KSx+B0ORuYbbTfLwqLSE+7Lfu3LOfEIB2YcoT2cv/Orm7W9IOqKEJghKoCT0uGG/MyTgZtZDx3KR
TIZAApn/QDCFwHXLvDMi9082ScJdrVoTTOj6Iuw23kCc8rvgKTIqRk7lJfj/lV7E89VFC2JWqWgN
H/EqTd2fvNwfaIexD7NEJHwSTOZ2K82++Nk6MKZ2tz5Sx06V6b3l1HI83VK1TNNvTAysk+MV0Zi7
0T/g6cjVQGhUQdIyPCAc4xNO8VYbNRFsy6ON4kMwdEDGkgcjyE1Md+q6IzYK5pCpSkNg5Y5Vw0NF
8dl/2ryptMmp+ZgsCAF9asyDZw8Cwu0LFuzGWR3xPHae1nGtYGLtc++2qnjmyIV6PO+5VWnWKEuZ
8TT/nMryW3lM8Hiq4xm7TukIuEqY7t3qlMTrqQKnThiLp795t+pGaicVpOPOX04WAd2fqqx5p60V
v5CFhNiD+pqiZ/nUhcqKB8x0ZswVbmheIUsWkXclSgQkyUZb3QbGlfIro3tXFdgObIalF+sFp24a
ZF2yfiEgBJNokyDUZk3KIhi0Y1mUOwH3cbNYH6hq9b1P2x1B/LdZooJrq1hNSSlYnKwXLvL/5xrn
oYYVaMFRBmwauTKNSw+ezg3ZIJV0O5+LMFrzkvSzSRI3t6ZXyzO21YdynGiL5nAHoopwNC9F6YaK
glTKu4GtGmy8TYVPQ1FiuO5fIci6i0cTBPC1O5zbkWzqpuIo4JR+xHcKwiG5tFOCUwYaoRYkZ2FF
SS8l5jD2U4DyxYhTJPrjTsRJHYsyf0517pH7JggrEJ5VaLV2LTTt3g1AEgHojXDcv9M4ma7SAkuu
rfO00IoLPt1VyspRp705cCVZM3T/qtk7DbT5Ygb/P4EU9JBHb2S1P7MK0hq9KjVOg+AbweXsnt2I
LJFo+91ozmoPhdMoZ2uRvw9MEH0Wb7FknoSYAt7s2C6d7l43qq7dNp1m3aTs8j/PUlQIf4PdCxwX
cdtZhbAHD8nsO7Dx6D1Dt1iPAbynh4aX9Tt354b5mbBlqAIJ0U4ByuhSn4dRHlIEAM5GAPKGHSW+
fLmlfA5lqqAB71rP+NYSDojrHG83VUNaHb3RQ3c2zV2uf2ziZ9b1lN0uUyNqfo+uiBU6fUjXIWTw
Ekxr/totCi7zB+hKaqz1BKGbSYh66Hl6sx0w6OcWtUsNPts2zh5X6F0Y2qU0g7bs/tPUxHaNrKJ5
xR9SI3pIdeDlCKxRI2aT6PkFWOFxjtMBcEdWwhhg1RomLe7+8OvAjaYNI5rju+aTk6Tsv2bG+XRZ
2rWHZYSobUDrcEEqPQeRRcG7tVYJThsMyq0nsdAvh6/RRbug7cjzhshx+y1Ljra13FtaYd0vyAhx
UYvPN97qTTrj1lop4siz8I1ftfSnaf0IQ2/qfMtZSjb/wmMc+re8SmwSK93UVVMiOk/eeBcGS/b4
L8B7ObxfYYIBXdSV5KOl13vO/tS/v2zlSTYeXeZX+SG2AvPheu0LBzIXqMGboSNWT4wSuCDbmkO2
+qtDVJxj1+7/c7o5DsPUgOJvIBVlSamiCQ/GrevSGlgytHm6+SBq5ztGIQ3RFsYO40QzP+4G1mFx
qln6mGPAIo1v6kGYkegSJBnlnbZjuvIUgybIReaOgL1MO4AUmKrUQBdUsW6d/MxwhG77xk8fzOww
QLqRABpsetiR0kmnHJ91yIWFN/43SUU/UzJQ6K1sfw9DimsBLMcI1nNBxW8YNUIysnEmyFCmgx41
rQC+Ph70lqDme0MuZn2RkyaVh1b+sqC4asYhvHhbxbHnG7ZOVnVvJc7xUWguPzrryiLJBCFTpv0o
XOYflXok1MYivvbNrJeyrOpp7yj94Eo/ALnoxaWmm+eWzDfkrIc0T2/SjzMecVzgt3OlphLTVE4D
Fz4tyKziMafwPEp6Mvp03Ub28/g6qeflpOy+aeG0B3zp9nbbCqSVzT99MbtESq4DDOwB1XwBzfjK
6Nsk/IJekGZrJUBC/zrcJdCZcEO2ng+nrrMPMC6sI287n3N7HARBR8bEI5YdlA6Hnvqm0r71OQoy
N/HujlLwBNM3VYG4XhwK/ohJunW5GWF9l8p7xPnHdUgrNocL9CjBO6a1u1ARtq30pJBSLYXf6lVL
OZz2n8BohchBLou+k023p+bDBtWkmbwryEkn1SWCScp3/sZpWeyWYyBcfQXSesrlv62L+eKUrkQu
MohszFCUEAHMwbK67zX4a2HTSMi+MbOKhWA0jr9CN25ng4Wo6H4VQhCp2sEddnPlTtrVCvYFs7yh
Elp4ve+gOdTQN9QGi9HTUH9JKg/bqCSG+vmF8kZoJBwgEqbzBekUdODhCSb8nhbCwK45+vzlhLSY
ocfsC5qBtyYuIFe5RgzUSQlG8bsNTqLzUKw/vnmecU/+F/qfBxD9ExjDysabNbtb3NtkOMHmEVXd
UnP5N/pAZGALgQwsYt8qg8lPSsBqS8CYuVKwWiT23B9jDNAfAGq/wQk2ZDqm5TTQS74m25yHol3Q
I6tjoHDycgbCcehFwtP5pzacmZHbqJOu9U88IB6iyrhy8U1/OCbMUpP8YLYHPf3dFrVckFMS/Y9H
0GYtnYHbKV6jzhWVEnQiBNZvklMgOu9BEcNWt5lZM5K6cMZ5Soaa1I2HVHKNXV4o0ALocXGVjQjC
k8ybnemiWW5n15RoJoPRPRhl2+Uq8UEhTDJR+whPJ/uzmTQhQlfkOEQ0J9BetORTkmlnnqen5Kx0
E1WCpzwbYLuoJjbE0exG/maC76iZ7SQLpyWPT118eOgPRUH9wvUFZvUu4Mz/ZSKM7RcbRxWuhiuW
wJtJhnI5ygE6uw8ouGQ+ZydWE4G8YUpV/6JQjFXa9cT1way+7U9grIzrsaSo2kMTHNNj8KIJUV8g
thhp2vBgCnRIC8p3mQ+khBckX+KZcUYuPp3raNhPdRJff5bnLzXijo34kLzxwJt4qdLk0hxuLNWg
GaHPlo7iKjLmkWN0Fb6u2pDg8muU0izFYmtAddpigtcDKfv2Xv4w63G7EeiC7TdPRmXhJAeSowqh
n8VXKAo4GCGeWaT80FJ+TLO0jjLUblFx7kYGizWbBjwFnb2QHPFU1QBskRbgReJkfV+SfOmSIXHR
d6L4po1MF79sC0Nm/x4bHdCFf0XeRVBugiaRv8CR0ybhoB3JYnunvcPM15tbcAW2k7CInKLQr440
NbXKBrKBIOFY+lLPvyTePOpJv3OnJ6mZRHrLW/jGLZHIJ9AVgjAGmidTef7ef0WtXFnVN88f+230
e4pQ1OfOwcquh7ur9RHpSFAKjsUBTNjKrl/H2s5CbY1B3DGQulOo9y1MwJ1pY6NcwBzKrtU+ZmcE
NKxCh3k09xiJ8xiFqzPVb6QZEhgFnvEANQPjUWcqolfXA1uL4iFrugJBckcpwEHDjiyl+0kG+GwL
1MKcEsAelcYZ8U2njb7kMgw1g0bKrupbYhNVxH0pWP3CsyDU6StTf/NNoQBZFBTV14DE4JgdA98f
vFmxO9czvWWR3tTsF7qklG9M6m8UYvC+m0A8YYRGKgVNLszbtlOaeawtQ67Eu7hPjpsvwzSoN5IV
kwUqKhKFWlMUboA+osnxRJbBW3DCTqiPQFyJiwXf8ztEnBiALhC0kusBV3zE3ktp3Mc4mH6gGtMk
gvIHkCBg4hSG6DXltrgeZleFNMNfTXNNOkIjmYVrfKZUXe65PLzunw09XbXAme22KKbL4eOkKZb3
+9elX1jYpZMV++z6GdZWupvaSMkLGi193jm0A20u0BAFOyKnPoPLSE+uBk9Lw14qTCLYBcWG7zxC
zabSrX2sWF2SdP75mOKTGX51+SZLDsxTVBRvuzjrl8lUSOz9UXijSZPmSmBp1teyg1wBYfJjvaGT
WTR3G2dT2kY5eeN1FwPbiOpQgy5kYvdT9iPL8KDwtDnt9T9223KfBIyP7t4fby6pL54xDcZrEBqv
XtqP8E7ilZ7MpRvgZMYp6vAfHvDFdAAMsIdlWe7B8GzhC1M2Y0KZXPjZ7Ar0nlZSJ04jM+NQbcsr
OQUCWVAPqeIy3o3xg9kWCX+NMfGuX2DqOE7+3D0fqtAlD0jhHsAdutDtxrwJikfB2HntAgygGetu
SA2HqGbPPtSXi2exDIya9+PKOgofZKpRN0Aa2fiZWmfBerqeXoEFxiYOQORpG3/3jU/Cb+sQn/Fo
qqlHKpNoFvT8AHuq3W+Oy/rTeka5A5hAU8x4DlmulRJkI3VbCnrUwHvQPqorWIVN9abg1qGxx7LG
1vGZYVXOFuwFYIWzX7tOfRJ4ABfoOUCPn9CNVbniMPUdCf2YTrs5gDqFwo/HVbrN1DRFPBVgglP/
8SSkktXbTwplFLDkndyPjDKPdJ3f80cjL+Vz8uz5Ve1dhPnxH2uI7eMzwqKtoYNW+i1gGDHNrBuv
SwFg6eeb8UgmylVSgIUw6+pl8uvjN3N2OecloQ+V/NsCeejhBtrn00eXO2ucY8qF1BOGKKzG/Qul
DbGDaKCd5SLrQhxIBIviDxriMsoa3EKnaIi9N1TLnlzrVgY2dr2qNTwA647yTSZjY78DeDsG28Hd
SLdlIKPpNM2+fv2RS3e+4ttGfcmqK2rCRMmu5te0l7ZqI3z/BNfg1+MneHHHSxjkrCRxybTD/N8K
4+S0VbpBDTNZOCxEXPnsdwQntl6aArPs77JKpSi+T99kofaFHT/qhAL74VP4prVPR061tvVuavOs
5vKQiTtKWiR1GAd0Ka2fFeX9Oxy4nQb9EkioL8naUpiSDDyRcNQGrznEkYlenyMK5ANy1sLbbxHI
il1bALoJjHUJNZP/8POuSfgYMe2WcAR1dDmslrJrjptABPRq1mSza38eLwstR4eNc40zKwECzZUc
zuOvoLresWpdzg61tbdxhEIrAqnw+j0kGMlvJASEk0a3vH5YWM3vHfdOd5qjiHamnte/Xy+kKLxC
uDDA1zPdkPRXQj7h6gVw2xWWYhKiGXVElS1tfHni0XLNa3KrZF+uQOk9spsOyVbv99Ho7Vh90vv+
YImjdmn9WSoi7gHPeYtYKCwkdFtdk71DsGK14hCi3Q0Jmswh6aHkNBsCi/lu09aoGpfPXiEtttCe
NbTcSz9H1fC/k9SzMbIwD6EG15chxmdfsReqfXZj1bSdczQq0+oaDIGdsDA3bwgu/32Y4QOWChfB
pcCa52+vTZnUPaoSvIyM4g9usGAo0ECSkEwdKe6IdwwZoKjGKjJZAoD2qXXg4DfIZLyJlPPvdL28
b6jJbeoVqImq+MnmxjB43KjieF9kp2z2ADtizrpDVjhh5AEbW5XsEdfJSwnZclzQpbvm0OcvGLw3
/9rmlO1F1IDeFsvr/ho4tHtpmUz/efGQA2qUSlrKOClcycF/+eJDIWEoVjI8KcMl84uaXMkke+sY
7NUB0eazwJKlDUwxWa4NEQ/l6XYVOWflt4pVRV0gPiM+ok08TOsjdPmz6pkTmejCMfUAeNpAajUa
LC/JWjx2/6RKZSNrIoDma7mzQM6BZHlL6mPYj+unLm4eDyG1QWOSF8IGHyoG9w+72NIlZXaQYVWW
9rxMQLrLYq4MoEKZc786QXyyj3MsIHANe+P1dGfGtZKgH5sjD2rnW8LhB7vWrMo7i7RgCOX9qHSt
1+V3pfAdQgKm12eS/8ZUjBTrwdWGn0MpJTWlO+njXCU6RMdtKBAx0A2oUsIH5owk1m1NdMsyfaRQ
Zt6A02xPq8K9VpxxP1yChL0JvNhsKGDfj+mgawEy05+2s11CGY1UPimm0H6W64rJw/xqxg1MMgWF
PQuIzCdrOK6DhFNMT20PoN3gg/uRdacee7id8tZ4sVAammCf7835uTVzznvPdPNcwaHrHL/Fbe/k
GabUQBY7QbxkaWSwqqmEOElYGQDdGF9XjRXkbNdlZex4Mf9BH6xkXztpfDNnkck7S496lIg5OahE
gA9MCBqy4VeDZnw938CRFbhdCdPKeJ3MDuaByH3BvGNev+OfO32L0NzaRnjrpk4qUHFPfi2Z/fJb
Z6Zqqgv0j15zpNi9xP1FXjEhsgmklkvKeJWP/UD7Lloi0J4AXKmM3bDlKUZ4RZmn+Wj5cw9kLc8u
8dPXJf5zdPnpsRzCV6gyibH2mPjSSwLFMZfLJYd6wcoeHT8LXmpDdEL6fkT0ru7lFxkFQQ6AdUnP
b5UrSzpquOcN6Wbi+0NxLwqXNQZCDOfWWwI11Jg2f3UEOxfEMK+vVgUHVqTpKDN5xY5Tnnv6Or2X
RPtESlMaXuZ512LVGzihaX09/R33fJS/08VWmGKeG74hA9Am1scssT/op/PRdli1GVE/mvbKAi+Y
7AWtPMtwNpnbL4LzxvpvqOPqKr1sxeI7UnhD5sI7ccGFK+M7h2thR2QyO/YVskdzOhzBuSJ42i64
e6SUKWSuaLnYVIoZrs+1wRARic1a+bn69fp+KSzuitITHHllZEnvjYyX39Tif2pQOwOjxONmn4UN
YzUqOxYi7hYQy3Oz5R4H1rUlSsRC/ID5wyYB85j+JXfaZ18B+ajxLE437qWWsASYior6D3hvhM4D
KnusXZKv11ax2k/2yK5vN1ZwKGJhOSR91l9N2ErvhAg7f3NO7hiTJ/x3PuUWZpGYWiKjIQHoFuha
m1CJWLK02nsVoXfOKyb5ZT9c70dyUprtmbAgbqibc0pi7+e+BCyWmkETmLG8QSoWfurBaCIn8uHx
fux1+tCHnbQeXs4zYvvOJgarxUdk8WdrLhqr9jeBeS0q9LK7j/bwa5Pg/1p05ufLGIUAqGJfTiVB
yslpKQ1duVNQWQkhNa/ONKMTwVbyk1fTohIqGzM52Tsfw+FieZtml1438MkZeJdi8PozRSDctC+H
C+auMfYgLqC2yFHbaQnKhgUfOxkhOMpoYWQ08g8TXOPtPdL9ggNXPMhQpspfUsys8mFZX0Hjp1d/
bstDSVTqkT90oo3LTHpOnnlQXVFdoQSok7v4Eq+gCUAIwwX4bb1whw9HoaYGZdjCkrAOtd3s2PdK
sz8Zorb2kqyZQBekrXr2FRVylEYx0UyBco9BJuMGGn6EC7ob1RfdG//MwHZS2KApfPi5QkKzUhvn
PHbe8iDsoOUBDUC1Ph33y0xNlheHvjsdhnwOcfYSFhGQ3KZHtX0Izei41VHFNSfInirLbW2Kq6Pc
KIVR3vV/HBnTt83w3QcWImA9JbHenG56uItQoxXTFRD/eQs0od/7hbZB8k/QYkyheOMm7Q9dMh9b
bex1o0iPh3P2GXB/woe+XuNpFXgCcBWEer7uei9OiOBwNFNlDZqhX/2wenfizEvcm7RN+leCDl4M
7FjYnQ69CCc7l31hwp4GYR0oSOphe7CzRefjbwXLiei4dXWnj2S/WALtsj/TQjDn6t/bYsSdT4xQ
ihzwI0oPN7XgsT77hAcQA1GiXquQbdj88QhH8hBsvgBFpvhzd4wNXEWiWVXdnrkKEqBpQo3ywANd
uWi2umonn5qI9wFGDJoaU57omZqbYIZ8dCZnqso9PmU3aDiK3mXrRqxax1NPk2boTkpanwd5HNZr
fNCXTvMY+JKWeH16qJVqMuc9HBuBce6CRzToIiqrDmwvYA0Oi+tcXEltJyew/jx2ANikqk1e89Je
aFDhcarenSGvFW0LIY8r6fyhtU6nNdUXT/5Ot5mPXHkcy/l/zgtqpdVcuuf1eTJWuvJRVZROmobE
kzC29Tt8J53clceHPi3HH14Ils2wpMvNbtn6Gw5TwigDlfhZ3ZCx5upWDE60UN4ORX0Q/nObk8YR
D42wAj1hL51iciXJCNj3vsb5P30+rAzcRAa0SIK/WCz1lwnWS6zLoSRtNaZ3ysza9/L2Sn3PPKHc
3EJpjdDqD5iXDSaGLHRhaOhrHvpDeM1HS7dqN9B7Bpct3e2wzPjCICVBo54uIP9JvKQWLBbWGmQc
7X7ZWM0+yAojbHEs84HrhIalyBFA0dU+MbDEiVbj71FpPxeru0oYFHCWim4L2UQmSfkUU85qBbfk
kkoHvG+s8J0lVvJP8prlXUcetN9X5INpGtmQ8HMWXvwwaxRhtTp+kkjoSRAXyHkNOTcKrhZmiC4j
qaR+IaoNS+OipCLXR6nS47ib32nVmRt7ShtLJUQIoRP98CLW2VY5K7FNsmu+4vHU2KUmJr007wUL
NLWYv7RCaLO/0Ss5JYBuLjYlAH2xkB3D5XnOcI63tBmGuEaeatU1ayDyZTjyfR1zIsCdpXX+U5lg
3eHKDNRw1atc0jdsl0lYKNdGj9nX3OAxiGUvtLgppHolCr6LHDHr3rMd4aB+4KAl0XbSY/tPBDdm
5rzqi0bAHqwR1yg+0yKQJteRChueKtQ4OrwDl6QuM7ZpfJcYMaofz/U8lqfy6wtoGcYEqB/LSSzj
TZcbkE1dHq0cz7GWYeV7RADWZc4cKO3Gwcqavnubq3Z+OJvek5xacSn6HlvgzshxPSU7kTMMg8we
3sDdv57Q/e/oeCivuDxZljyGWl5H9gfAXB04t6Ow1d4LuQRRZjE1N2MBRPMZUkhOObO3mMlkFpUC
QsYKmElZEhcCStcJJwBbh4mqs32ZGodTEo+UB2V+HYQOw6sIe/PSxvgytbGUjyULNLxoixJ8PRBd
F8Gjg9QbE1lQcRhbsteSeUuDIHisMJ61MADcXdHS1J8MNXzFB6IX4ZFWYgIqiBB2bgkWVtjtvNXv
nUI1I/JLnlLXhaZNzGJ6i+Im3oQZ4TXn2aFmwcZDMk+oyOq4ggw3vG8pX9jQxrBYXLzolLaXBaML
lnnlghCpccLyzJOAZ5hRDWQ5Un5Wiaul+/wGaXXtbT8WzemN4x1JUsHJnv+602z68IVz01oWx4VH
MOW6AgqCbPFpfAGvVV2f4+c56RBaLK1xY8P5Kbk205zXiUPU2Lg/ng9NBkhbQGfQFw1mIULS71GW
x27dU5PvcDvzIyRNSIcydD2X3o9JRdxAJhNL6WmGn+oTKLJb98MAtx/Mcyf3nFZpJVU7JynCDFGB
gvZKysLxFa3BC1RISskpu886c/u8ha3eFT5Hx+XLjA4lOeDiffMDjEr/OgN8DlrnhiEft2wfldGt
jKpoAHu1cP/c+iwAW/sz//fZg8HjkDSIJjWu+nYKVZPpuaCFxEJS22ibQKqDnBxQflonolFAPwIV
GQZqyyGYBn0leRJpFZH6kg5M2j+pZcETwXqVcK/Fgf/aEaIkv8h7Y7HzmKUXCyhdjmtSSDI51eua
qDtwRl6Vijbilv1FHz/m7us/j7OunouFrXIGkUFsT+f931FuaqW4dUqiMV99saOelr39967IJEbB
i4VTKXvCUAbUtLU6Z4qufUaRp/QAsCwBcSdUq08IgOdjkvlJTCA9OtR4jTiMdJ1jkAGYD3mIOFsy
iEm1uqrkuy3fiBe//Gwj7vdxZ+7sam/eqXmNgSlkWGacQB0ALaxe8FzcjDKpY46DXGQgqqmrLnWO
KczPZvYBvRW0Bgk3fvBbnAGujazLRDPI4I9c3hxYHG7m9Eag2uJaZJ0wt6lmDyirhjSXu0Cu6vaP
ylz0oqiuoRhZZp/gW8u3Xv2yyoORnQhPS5oGAyqRXt74IjoTEjWiGRjq9U8Tx+wtlbRCfN1F6M/U
HWMY0NUlJFNGHqQ7K1IaGr49UCJRS14cXzdiFzO5lZLVCTkKJPGnPLY9Y4Uak6jT+6+7Pke3Pnz0
uVWFXyIft192f9xJbCtOw359BaIX6Tjx1T8ckIWFJkVp3oejGqm/+fPZqfihzBRncexSlHu3MJPh
6S/xHxpQDKna7cMJ6DDFf5tC3NE8TmXr3Mk+/pPO3JqXyZL8bACis8B708IwkSiVv7S1T8a8lZSo
tLLodsOoEHK9VI+Y6MPOAdP6xAtX/Kvqb+IHQXfQsJ1daAYKxwJG84zY5V94OuTNZVg/j/FU36DF
F6Tv3lF9vZorL+1PClF1PIUoBjTuJZXQCy6/sei5UsDMo5+ZNLgvP49DeqNSL+g71Bvmc0GymhaC
xN9vZe6LLFBR+qS+dGtQ5HQ3symgUpEn6K5aaOlrDB0gtLB2d7kV4pDfRbwfIZPFca8+lpjqQuWc
1mtC1V8kLb3lAl18vkEv1Sg6dxb5BFIrrMYRF0MfBbjkEB9m3AhRKdmlGUjiYWHS18xg6Kt/1N/8
+L48c26CoZDjYoxcDTr4LuZHkDVDzVnAkUizYl9rGP9WX1xrC8QNAEi1RwzkStlQv46Jyu8P424g
uh0cpeLeX8uS1rB5DsdIuTFu93c/WkIZp1Dh/dBl5vNu4EFptnSYGlyjjyW5Fz1MZboyYbXcIhN9
1h31RKXK/FTQeCipznZAHEufBWThEcCtIMJHww0iouPzc38C7o2wou+JSLI7F9gs6H30FbTXJh5P
1SSD1YVmEd0vQoiRJlP84PlXc9qVzI2pxZtHFxtqyfSbLYf/YUP0lVi2iFRVd7RbsGicvqNSdBL4
S+xyfwgb+rBOFhpcAuO02i+fAg3YkcnilmouZ/T4D948qt+eF3D2QMqQkco1hIykhzdaztMz2m4Z
5Wh46/yrNBw2EfxHPJ5V2f7+HLpXNo21lAopdE4Uut2cbXPupnCseIc8bCo+2wv12fX9tsPqbbYG
JNPgHYctsXREZsI0k6qEpmc3OST2q66uzq0JfxPWmtZk+3xgFHiSyac1fhchdrKNbnXKILqsv0RO
DPehBR8O9IjJRrAL5kBojw6rv5zmaD0qyVsL7x+pRB9wQZ1nod/MZ4ulQPsympOSNOEo8YuHALrv
Ama7cQYfZuiTEwF+yXqD/fXlXjcpuacEMdKeBuNXFzf7/3nO3hfl/aubrWL61U4DiwxtvLD4eZ8a
Hj76tBIFQ2qahGtzwwLn5ANlquWh9bKY8PwNPuh0F5UOzvDG1yoQ+OVaOKnToNayHD07uK+4/OmV
ID4vaSIHQsAro7jzXEVxJ2OM066VyYhYm7IbBL1mQF6u6r5lh91QmOrOdqPmS13JjGdaKP874Ktt
YOtSUeC3hPnPEHDt3WcEy4hlr3Z11LaXvOVUX3UnI9CZbldlK5kTFpJxcRwHNcwJYww/rcNpqFMj
q+JvEhBuSSWKDT2t87T0eXcL8esdlqL88TTFawa2u9pd3Mpto0CzDUFx5YGWrkIMpaKGkp+Uvghv
ZhXsuEebdiAmON/JwEZZ5d8DdOOv91USX2qO9W0yiyegBptI+zd1PIWg7L+tFzqLLiH9inX9xFrO
8F5damLhSSuNvkN204C5MM9L3RObChPvlqVTPFh98Co6VsVWZrl/UGyPp6LWSP/iL7Ikx5SsOF2E
PZWQXaFeDAcSsIMe4/vxJgFFP1H/B3diN3WH/HXtI9W4fC3tNzO32BEYJk0ifIcwTEbAFBLHWF45
4eKGqIKnBihMDtdUYrIwttUXO3hK59lPH18/Rgo6CW+e0miwO35f33XrIFxg7UcWPbqnp2N7YG7/
Z1jJaWkFo3VQwYEXttDmfdsA0oi6eeDfOl1PLbAmX5KgPmOmEFEetgXhYOlD67IR7FKz7fQvvQXo
NMAAG25rmdG5T7Kt2PcA0CM57Fer6xoarFPbZHmo+uyKz/CcY2cW6Q6X/C0kjd+2/+dDohniDotG
GkBqxbMtyvzDSj5rWMYhGKQQVKtWHJdSM7GzeqAKCXEjNq6lgU8SOEaxVyeoZtXcYABBtPwQR8iZ
XyJNZZAcZH/dFaRq2E8hzB7UnKrD01lh4KAq9tmaBBPvUp3r1nJ2EO0tYAct/8Agg7WXOMaDjPJ8
D4tIan5XCvp5PNpNIe9tPW5Bqj0bfwQMcLfOny0JODKwZEgBTHWiUK/Fz16YqVUCH8cJUsOsVQWa
gSW2h8jwacy/d9PG0o8e+mAOPfMOgfPqZ4CIvFKnpCi+kXf09yKMicwHZIiwgEHOb8WYPCzr9c4v
JTLHhKW6y36+UddtyHyhEh36xlponcz1JPo09jpGaIkrPgJJRbHR2fbOjaaKxwg7qE3aRXt53Lnz
ub2noHZ+SbwNqRWuO1vsqqM6Sgc7zfu1rpkS36wpv/4hG5wNWQYmHwCbM8LbwSdvLrNtf9hIhSdP
Sab2ZvqwsnF2b+JXmBYXXkSUwx8Q2E+UyFxqnYKxgAzCn5PBGjP6sjoxZqHSCOggHSI/6pMXppds
rqLCLSiFUWTrQyCwulbB+HV7c41MlPROEH6otk27LUPtdYSvms4aYUkimuSHqwMwD3j2c2mkW5nA
wMOxL7kiSlOq9EYa+kSY6HPKD+/b0cf/cpUAC7J5kK4j8e2iFGBbL0n27LQ0r55yiN/iQY3K6Jmb
hO8nJlELWwFE6R2IQJ/x7dU+JAEB04wAs1pFSK7qWBXs//DuhyIGeRf4lI9AOrhTqzV6xRIQl0dG
hd4zhxWWoD8KXP7LGhu3Ll1PmbdRv6hMpsDfNXoTCDf0hh6ktaVyQQLBZP/vwjjoHo5rh7xRkA3v
67EgMyTSZeqDQDdn7M9W0lKuLbzW+DiJDQgAuq3gVTbpS6Ke6n5+QMvCJbmoyJzadGhOohw+Erq/
HfEwWlS6iabU2w9MVqTgQUJ0nG7l/DTmFkE0FYsTLhZYoJxb3tgpbDMZof5qEVi3eEFpSHAe9xeT
dzLgJyl9UIrQnU+jKYckTtjTh/wVmx68cP2jCYv7ogvLD6R09eT7zIjSl6slw4c6AcL1vMObKaU9
6sItk+p7auzcefv3ckfQLMX0oEE7hxOxBnqaN5TFuBqKAKr6ACe5PaqkxHuff99sj6vx9n0a4XSm
RF8tD+010jQITezb7Hx7gtgmr2gl/AwuPW0iM4Uy1BmoZF1rQEFBHvgectg2HUYDm0CK4Lpmj2S+
HbbgdzJmKahQMcA429rnbFaBh1k3USI+Yx9fPh0RmUt3dTsIOn7YHhKfe83kDnMIxBp/m1VUCLt1
AdLt0WP6/FVrzLOO+LnLXgW/Wy/wSgnzkFH5dXwzXld8dvEqU80j0m4bCpBNk1oj/qEmq2Fm/RvE
2AZcRySmuyxBNTT4xxhX3QI1ADZl5KFXBTyM7kTe5Q483fjKw0Ishte+V5w2msmbA40fb4hEIRGY
/VoV6GRjXHxpNc2wUt4I6AHOKwc1tIr+4Eozg7t/NdXk+0c+LN+EnrBIfb5cqh/gm3MI24hjGGcp
RSOCD+mww0/vRqUmz4ZaKhacRHZsGFQh0UQ0BdppikgCG6O8/BN6+y1F+2D5FE3mQyOary97dzAF
4abboSah7H0FL7owMdeDjXBgje9foKu90vdBzsqxzCuYhJimmdN+KzLcO6Q7ZD7uXnmVrtdWNN32
g3KrDza+DY7RSpzeq+qhdjFfcF/YYm+yJ2/HWx/O+g8fcQHu8+pCDD9mXbr9UfURVhpBaUO6AhAG
f9iSs1RvTrWlYLEKvrhAby/UClt12dkHeiTzXYH8ufPGM5326oHOT31oKuWmv3IyZRC2UdryKVQp
sUsP6RrjhMvx6fwEfsd+Tj0J+OzRTMxWF4XZ6RFcXBcdBi9pbn6X2yGUIdtGdQBij5iL1gmCKkyv
noFFeD7cdt4sIhxzHjvCU+OU/re3AhlYN1U8L6eiZ3A9HrUQYrKUwSUetP/voFKeTkAqzhhz4o2b
OLg73rdSTt8DaXMLHwOdiqND1f/OQZg5l3Q0vAMZ32Qyh9wkmAaTiF9spmgK3/7i3ESDVluAbxdj
6R3XXAQJ8dEvLE2DI7YYVfUKMlX/fJ8FT5QkF7hUSkejefR9X01BJ6F74JUH9aXdzwmx4xLyM9X1
K+uINLUX4/n4qmG5t1NhqqxyoXol/HhhGEnIv5e2bk9J9tNgpS7xi9a11s34Aj8tLZeuGcra0s2J
vHiG0uTmbpUkyMAE5T7p+2MBXD61IeCImL63NUfcfYe9+PfLgZL26FmqiIUPuJvANBoS7mNQfZln
bZ+tYldIvY5fyUNujNUSz2bt++NG1h2hqucbwgcKMcnIw/9V++UtgYYlLbSbsUZGLiFCS5qeHqDL
CJWw+9rUaL1+iE6TNXJ4SZzKtuLb+bBgDCpx1MARKdqhmBZe/ZroXn0wlK7xg4isi5jhZu4F/B8p
FCZQw6UEKulgZ6vVAM27X3X95L5uzk3mWSksVoW7pDLD+wKVvdOoSvomSq7dngIpcX+JOWY0/YnD
MfcKiV2agMWXfsOWnEddCmJobVvQSY9bUF9zRKOTdfw+I3qRN0v0Lr29aIa94c+qozEKkBIkSEUp
Gn2I4dBHXbqc4mbRWwY3AyWI3zQIElF+0xmg407yN3yAxCW2OqGP1T6WMyNOh8JOtPQzDCrbAT87
CR5/DbYlhvJPvKtbbQpVcF3APeOM6apq/Mo5YOPEVtn4C+/4Q+IVceHOO8LnpAL1hs3Xb3sOpLiT
IIZcfw3aDg7DwDwhjnWH9Qq2UVVYkOSzNd/e7sLPb2Bd0g4oiBNEafMFuOqRcyakMQYj25KBLrow
0VHHNnuOx7wJZmBtM2BjkWAcBTuaCtZyfMe1T59N4YixA2qz/umR7hdYMJmWF44kovx2IJn5Iz6p
ha46dIMrpVgnU2sx4DHSTfUwdQoP8o9z+xXofu6972vKbP5E7wyNG8JvcWwkn9J8GFfgEIpP2R2Z
dmdlI8EP4y9ZmXbTE4b5Ix80NkvKL6LF6cd8XtLTdT5LYfzPYsDASlWIexDiHKF4n+YaJLUydAaD
cIRqsTu7/eEZ/TPUz5vbUHwrjKRbqBEQvNhEvOqCey5hknlIDVD6uKcOdnjr3Vez2Ku1Meqdmyu5
YxlUtxIgppxx5hBZRLmrqHRy92+EUtH4uqaU1dVL78yboJkBL6+E/WwR+hdvF7GQAznUm20v/dpk
5a7sWT2jAJiSSvS2MNLY/npP+7ZYdpyn0YtHar9sq2Cmkql82lwYxCdMSDE+1yepwYYwG5TsP5Fb
TWIY3iLtL8YhbHLJ6W8KB9X3uBQNFjDI+9qp9jVq80CshutS9PsTWcjJQ582/aASOrzRowIkXl1b
DaMv23Ga2AX0vJ230oKeY7D0AM7osPoKXuzdWxtub794sBv2DcQIZpz3QtUITUvwo1sokJzhRpwA
ocy9/wEpEieudgYDoDmn9r2p1RF7JL4lnZBs/N8H/0lVxegv2WYmhQgAkT2ShvqyRd2v+SQGnaqd
nVB4OotaRc028ggb0dVVs0qstgTAakWBaE/cjX1sxD8284gDsij4uuI5ZPQ5TJiRId97n8RpOU0z
30C6xQqwg/sivxtRX5Kt3KRIOBXS6u/uec9GTTBJCvPqNidj1HIh0qW6/D84zsnIGWn9In3vHSc4
MU0DZUSTdo0twM4tAhAz3G72Z1qbMA1X8OBPH0EYzh03jIGSj2R/ZIdWZTTdxyg8I2Lfv6XooCgh
65JTaY6SpLXHT83vs3CJQdH/GiODo55UyYJtIhxIR0JrFPBhl3IUTpFZI9dzX0KkULEQMbd7rNwo
CxDBwdOUpG5Pdekmq9eCNNMm6papMh0GcF670Ds4oNesXiahpJ2begLkCGh9wa87z+cdZ2GBkiyb
iHKlmD9yLpenApEbjSAgJG/KEHHZf5Cqm/OR8U9ReGsvAYgvOcEvaaMIHcZ8T3aCoWwl5wbzSb5+
Ma6h/pi1KdU6RU5AeYy9RIjn/1NWY7eAZW8IplXuiZRHaaTSMcm4Csh9K/DKlx46kZIPs66Ct11I
uPEJea7lH4GLj+PTzoeSEWBMKg+uSeVLW79R5KD7N81t4NoYUsmf9yZpSOm+J55v1juqn41ti8bL
WuawqsphsnO1TjM7dxDM+vGYfYpHXXaKBVht31aEg9o1mzU/jiqYsXOcMrxRcJ+UATp4Bp8JSEB4
fi26hOiEnyup/ob9iJjn1X2XbzFgPN3nBCw3o0my64T3nSGQfQW1oXXqitSn26fWqC0kf54I4Kk9
4bS9Sxr6EcwOpwSnM1ERE7LULWWv5U/KQqUNsoINqP4PWMFdYovSjw+4WafQtq3+ThCUZWTjV8/8
EolFQdTjam0pinK69+ml4gRg+XzMfPQFf8wpoMZnMwCfpO60OqhuVGfXsSjxMUHVBr/WpxStKNBd
KjKnmDMiqgHCB1s0uponx7/yD+d4Wy27KCGdCT71mdRjEAA9f5oi37IZaHEZXBPvV6YgfBOk00Gf
mG59b6h/PolyBHyRjKmwnirONThwB3A+ePT4sP1g4c37K3OJFXCAJHNi21cc2SuG8ufmO3ex+WxH
51z52DqaEXLSzvvgoPlmHdnEBdMPwVDe4TTRQ3/fwqdmih8XZKx3Ju/LKPax408AvCD+MozPpojN
DPFx/VYGq+3huljeSYgA++kvDyLx3ORkfptTww41dSDHJsEttHV2JD7pEiYM3nxiXeptjC8Ioj8e
3RdsaeIDnasQYsik7ADz5OAKTCDvloRw/CugRAwOcHf6LnYlPj+0JUQiionB6zfUwmb9n+jPCaRL
8tD6MkRKP7cpCIF9l6UQR4gyZanKig29N41/zISOQ+fHTCsRWuVsD2nvEOBp8TzvFJanLBuyIe0p
VzbhCWZC9iHB5m+OgHLr0Q9uIp/gC+cLTrc74fFBq+8x8nyDqXWAwLMudeyRn+h7tv2SxZtCH87A
UZTN318K9OxKtE7q0EV4KW11Aahi5DEfpRU1HdrAf7rLjPLqU8KdLUyzb3p+bcdhY9pSwNr+WQHx
YTp+7kdPGW9wwmwCT8tv9zKABW8DBEd5rvi1XL4GzoNXIGfxrOpVEg1g1JHvUoMFByvt1abKHyg+
oLxor5N1z1TQTKcpFn0ekjynhipofNBc/sHlafduhj0UQFps/CUsRthwUKG2CeMT5vjX21AI148A
RiisfH8/O83X3asYsHGLjT4JQN3Ik+G7DRNsiwiLhTfUc7hvyPdzy/xykLzmBn0Fm9EXpbCZwy8b
n5NCZghxRyP/Ap0Pqh2asz9HKf9Grn3w/b7vjLpCuSjp8J7yO0p1dD2rIp48WI+8gnmycB5HiDT1
z0Lt3yiQ92G5TPVwnRpnFIZtXlsXhXS+YUp2H20hWCxvTaaT7G0UGN7Z9OwNAeSN0F/eD3rFOqeJ
V0RxSqxqzxqXboNbgtVsBIve8GOw6BRQA0bOrY9fOz3C1saTqOTIrQD20OdL+Ou+kEi95r8aI1QT
o2f8n6yPyAEMjtO3bb7h36ro1G5mpwCdb8B9iC+92aLobcvaBDWNJayXcLwnUNOis/oy4YJITOyN
OB/BxYYGytyyKpGZKZTS0IWzPjFMjb+7WjOHZFLZgKxWtLmUHkgfjMPF00KJAfBAwh6Bu6xOUSeT
+4hnkmoBwc1Td3yTfNJ0htksZXhhrMcdlC054iKzz6vpWdrRHQCF8tIIko5IYwcv53YRS0DOKO2i
kg1CvJlc+ZxthRetaoY0K8siFD2ZCIfCDT/HVOELeNLLGXN+Y0o6LNw2fBzJ/1BxkYOpjAMsYcA5
LQ6DtP8DG14Gj9j5wwsE3NAwKbxY3zjoSXwpCSNHkEBnhGXTm/4jPNkelja6ykXgYflFsIwRkxME
QhoWiAo5uKT0gd9OLNYBmKnzkzhNdrLcFb0sh2p/fNAmVKv7IiYIWii1VmA0Aw6el613tHjr0lEn
QSvHNEB0U+2YoFSvs3XlNh3qVtu5/EyinVPbAbXBn2T+wE9l6mTvvM5LqGhiq835z2zmPRZBjoUW
NF/foOE+iJdPfWByEfJ7CQy+INR2M2ktahaALelUZQ5TxY+UVVchjqLvO1A19epH0QomgyE2+Py2
ptRRmE8hMYrCBItGY/2+i04+xyB1N79UNV1Byj3nqMPIdPE+KrIGJ7C9wSdwzlIMNBGBSQ9w/zwm
DP/eswVRNmyIeqbGm+m8KlFXELBX44QGZ+5dLRZVavmC0BsHXd69LFPecwFJJKjFtYVo/GV1dIrH
7a0DRwN+HLp/eUUR4EvdEOYmYGOi17gKgO15AUS1A5ZAHibb5pLMcKmCwoj8xB2bOIe3BxCyYpy0
TSwTh25TzIu+0W24vfQ1g974mYvwQKPAEu48+sJwK13FFfYJbZ0lT32frTgDEbvo5/clkVfY2p+Z
XQwcC3t2l8y+TORJzDUmUhBeBz/PglQ63qt1Mg81Ax9uLXhCdxenCar+OW9HjzFIXqEozkKVQipV
tsaSCL+1emggwcjG+JjSpIAYYEnAsbO7SPjIy3dN1kdgt0RXIlZeznBvWVGZm5tcQEKGHJB5YTYL
9dEk2dFsHBGfx++UH1evpDcnGXolZj6McbZZfR3ZVvcdf/TLdLy9JGZ3Zm8mdtYlmMnGBfepUGix
3ccU7QDIwL9dy2Zw52dUOorZrol6qP0RxcdziuyY4wtcs8qmWgZ/gA7WGv4+4b3B3b1MBYKkZZd2
AypBHWSSBS5BIOiKWNHOPobsW1hKAq+TEItAxHOdNxR5zKkAVj7FbSjnkRTQrMYjVmZ9Upu/n9go
/tLzJxXXfA2YKSgKkxxEE3yb9vWkjXnriBV5XMyCBwGVHXO4pnbpvInquQCX6CS06va4oaXqnDec
p4R8jUdiKfr7sBQELywdOKFB3gfJKs0TqIOc64YUJYMBVvZ/nk/vZ5pyoyx89iqfvVKBuS3dnvWn
sOCdlYykUVO7WzprLeUxFOiZSLcBoZOdAi/KS1x2IYqfq8MlbQN/w2K618+G3Wom6QtpN4nG6d3b
sq3awvkX5zmEK2FcUSlDVq1qMA1pjYcXUOziaSGSligGfUMjfxsT728Rsge6rJUlgT7FYoQZ+vOP
TLKLpihGuVV/gpAtoQD4uteWLIcLpB1Mkzij2faKBwMvM21ccg7zQN+o7HmQGB3FBT7nUOnGRqfc
m/eVOaobWmavya6b0NDGPefQ5X1HoI6AkYVp9dJcSh9/XZEXlt9TLQH2JNg9n4EC/G8eQ6pY7hjc
fibdaadSUDKHy/SEJVWnaEYj6KM9Pdh1RXom6o1/+XFup9FyICcNXHt3NQQ3OPR2rhj+0aeqZZwd
O92+OG1HSQ5p+/9vNA9R3EWTF1lOUQqAO0aNkNvIqdKv7WfG6ocsgedqvcT56bmW72h5bxEGAnL1
20f8trw64c/hgEAuN9Y7WKgwSYuK5btM6ToRl7DGCM5beu9v6/7JO4bGD89ACaIY5kKhp188lvpK
i91XhQOhKKGModwiPaEnoYOYyDe1EzIaX0IMbNwKadN31nFiwRtqJoUIRIfaDMO3pdvLtbXqyz/O
LxJFFVVTrLrnDhXRe8Ple7wd9h4wXaEhWQ8seC6JXuzjs2tYNiV4uUzDA9bYADqVU/w5e4J9UCCU
wAmPzTnE24q0p1kAF8Fq4nmGyMXZPQztzsQu8ftJ2bApMuG0OUDlQ0BoeKM4hyhtjipwQML9F22G
GGpZ3idcIDICpQyycxcYDcaHfqOWv6nOSQundR55hQ6L5HmhxVmq7xX9ncanZetnU3CQIu7BuW+N
AoityheSk820URh+kCZpXm8/XXqNcjQYrp8mgTfu+rq7Yf0a83+9UcMO6WmWM/tuSCSG2GTx8oWn
lLopW8q0lqVHVmlekkkRyrt9hfijTwoFne5RFnBuLTaVPQNZL+zOHSXlSPQbf2HgCUB5lkvkEmk7
K6AUCO+aX/rSRpbv52RB3m/aH5JC00QUi8T4KK0EEQKRP/SOs+PxzWnxzt9y9O98SoRQWYabE38q
yd9XDQEL6QYlvXYZDrKw3PCIskOW+Xwh3UA16yG4s6oGYWVhzET9yRDyB1kzxz/xBXZTXrLBByIo
NGB7W/9/yD6xH4Tso4/B+D91FO49MBvryfebEjhUXpa4qGQcKQoa4zymnSEB+A3bpOPTSYlwoR15
ytRK+/8VwSvrfbmsvYcIg6m34plidPWZC6yanswIfB0v9bxssjg5pc6E1z+tOn+PJ7MI9KYdqDgI
lM1i4+EvrWbgeYBt2jjoE7v9/ZWyNDdcDAcit5SPC4tLGw5hbmX0SmrRC/R0qA9Qbv5BGm6OL2by
n9kR27EBgUJAypCvdvNDK7LC38fymfDOmof7VsBjzgjsCiHJ95TdmFXY+OIrJbnt8/FPWShxENa2
k3hWfdJ509fOjA/kN5D4MFhnpnQ0wqb1Z/dfBQEqkUiC1fxXV1LlEYka9t9T6hY2cKRLzdlFn+jr
JslB+17UIAgG6BYPX1FggIG6uXFulkhK6IqJ0u4D98IBcgPHaDiJ1/htMxARgnwF1rlMaKH541Hu
M7GD1iNtexJLvz+Qhv2vWDMaecgx2259yUZZu3KHbUmSfFnnGB2u6tMqq0Ef2lEWSs5xo2ddrAha
u8BOaoQNDMsQtvKZVfWNy2ok0+RRnHKrI+xkTGmsbIWvTT/Bfbsfflsum+eSoBtE9xZV2phbz13t
4lmlRDj4UevIMpsFOkUAkaoQeHptXBVOO4AE1pux4S9XIoJ9C7FSQeDR9NJAyI2eaUKD9R0L1eUV
oblE7BYZ7RaItkGbDtZweLLDCkSr1x0KyAeSDtegZ/Mo3TohAG5aBO0jWviiN7L5XkjAL/ZQkX5q
6uxRr4IKe0xeCQmBq08WslcNoS6HqCNpWEAQ0rHoix9MWfVz2EMK5dOCKBi0Po1SPO/hTRyVb13W
0xd+jHpa/MWk3fcPhz3DfAFXXlULjFImqvg+DsfCbu//zLbHY7bH2SRpTR9hwRuUnvMYyRFyYx2f
NlZKqlSoCgfQtwIVjueBOKHkA5un6ONhOwEzWC0uuBm863kPV3PNvK+v92vuMpnKlmRz+9yDvgA7
P0qH3E2kDSIlUrGevWVXfE1qLoErgVbY24rJ8TblZkxT7NkFYy6ADcle18x5QP0Gq6ly2sGSVxxS
w77g2/P9Vmt8/dx8Dmuodsi8d1jiTreaJ5KlLzj/6k2AfMGhxW5gpi/G4kTXX87zVcz6NqUpkPZe
/ayJmG+vmx9hVDv+136qu18b4DTShiFU6Ecg/xG8xujYnCLOY/eicmzIgOtxL7QYiaj2qn/wZou5
ABv7Nd3F5S3bFB7OX6wdsdcmL4w/ktAL84/D+nNeSOiO+e/vuLQg7N0CpHfFn1T73b9hcDe88rGZ
rfCPjFMtPedM5AmuaMrMKNjuCQwJXlzzvK0WZNfdks5y4Cez+8hDC85/FRocRbbBuxXgPOse2qhl
SkLWR8TBEihq9bvVq5+Ob4HIc81zUdyq/+saQSMzQ+ioUGJfVj1yzu9MG6g6vV0m1WoKmlGgqH15
CgSp+HbG7ZOVjHbGLtoTPb437VILLfkXyLNkkXFcdOKICuV3l059ol8DQOzy6TDSArwLspwztEea
vyxTYR7qCZjBEcYXzGKYO6VanntFQ766zAJGb/As10CUukL3O4eS866eUqG/X6Awct5cePebjHtw
uaGBf01/D2xs5yaR5t0H/aSpfMN2c8Yf0mXDqtPCOo2WEKeZ7MBt5RUQKpW0GEeVqrEfFFXWABIc
fqlV7ki4LqjbYwY9BvoXni0ukl9sSb6M3IGyrfFrc2Pbrhrv+Bt/x6iXcMcChgMzlj22xjykCsCn
XzPP2B38B+5LkRQ9a7JYyX4vSSW30bFBv9W9Ioa/cG8MhztKD4z67Gf2imPyo4YZUAU1LMUCI5nM
naadVfBnrJE75pSSCbFW9LLvoSllnIGf62gO/BkDSvlegTVtRSVxjdTOTJnXVLFEUAvPS9m2+ATt
82H3sFmWqefpExJHZIcnf5HeZXiPAEU8Rvi41rQuSJf7CfiYLrzzm168BFHlC9uTLDPDhCWBctWg
s5LJZmr7XQGKDX3jzad9ksPgKjy4wW8ZJ5VsQDca75GjXL4nPlEhHrBolyWVrJbsJUVl6u2Iv4ma
eZmYtG7agjkgiAVCq7JjsYzpU5NwbvL+NAOiKVtT5wemLHFZiNMXNEMmmBtMn/v0aW+994Y5duqX
m9EvIl8zWh1hiHHfBbhrf2I62fuQvokRDOj8wVw1Pd76zj77SL9Uuf9NAtC+EdrsHq4w6zzYyOGN
4pp4zIOB2pkFA2J7n6L5ULiK8zCcMuwFJvo/80SDpemIpxm4bH10dZDHZnHOYRlzJKixvMtX9SyJ
qOwcRQLvTGaYOoW+P5y6s1pXE6/Zpds9d4Gj1H/QD6vicIuOaFDvAL3tRobokT77oRtscKsvdDht
dj5Iunv02Ena6Z3e7Mu6DjMREl2Oz89iqFoi+lYTLhxc49rfWntlepccEztBrp3DxR2GGMsc7z2t
mQ9uzXX3oAVvmJisSOod1CdS38zQMBi1k52pxVvXGbwjmc+pWXPXuQMZTFNUCnmLg3pixcfgigeO
7tLclfTIP8BvqHGfKREohn/BL75mEQz11D7JRKgp8MRyxyngrf+0NSVcCR9JiSTPBfjmhF+AUqjw
XnR4dL9L9YDjbxV3OXdpb64Fgynw1h/wflKdoZvt1sCpPgbOC1smOkMDXYIhKUQ+IDPxTKG1Jryb
t11G2txYDeZc4bRrGtaJMzjWqOu7mAmjw0AiIClbudv+dlKoLK7T0vv7aKnkhy7M4/oqk2svchKE
5ytPk4Qkim6AOWbnRto+7svvWqtrqzfLCSft1SofRGRwQslRbIn5+ut0m4rAhtZj7Ios+iTj1fHa
1P1WiSXvmIJS6oy3I6tacTH22n7SIOuJ5evByAOlIGPCn0KLbpsvmYZv/3wWUwVxWwSREJkjHTpm
38ky7xQ+rEG2jn/FFfWMvJHwkL+H8wS9vzQr7DiBzgZAYR0lv8phyPNtbVSkGUME6UTonVejmFMX
O2Sl0G8BrqiInK8reJfGGRyw2bBlCbni2kUXz3cqXMf5QdL7EXMjwMBh0I79+cWlAZt9bfsbiaEk
HRQTYmfW4mF/J034SFbek/FRAyw2K/kD+HFRoLJOXw5Mv3a+vtPiJJ1OHVZvLVb4DawYmXFSrHzZ
gl0HiBTD2g+umIM4FhDG4KZE4Tsz7lljhGDJCJI9fDuzxEjObtDTO/DAVPa1YOd+4o4dXkY+BCUt
Rq9ODS8wghnae+CgR/Skqs4+gmzwhcERwPNNM+Tb7odCQKPMrwdAxUeGjd7y1PsTLd2v8U5cKVDn
1TymEoL7bTMZ8fU7tOSREztZHOn847lyPBETvvxB7wj/LCcnKkalSgS4HaB99lOcg9fH2+u77qzS
aUGwhjwKmIrk06UTuSFJmQHP8rkVhvcZxp5NVLwonjBQAWVaAldY8ULZVbOpPfzByGg7OHkBuObv
5cDHRnDENREBoWTULfzx5nitrDrxLR92CRZWzk7b7YZo5wSO4ZKC7PzJ7ZGVneyW5xH16M7R5NmM
KWaTZkdzT3jFVL//LgH6kIcDbR9B9pywFfzRn3fmTMNctU9Wqzd6PXRONooS5nwSiKIOVyotV1mh
bfdspD6e4KwI3MlPE2SxcpPGowIYFqHNFHCTFGmYNK+e59+xEkIsXO/rF/IheRoxFZo/uOjbePid
RGQ8SkMghSub2rbF3XHTdAJ1YcKjPq5q0FTvVdLuaG9J+CSEdiUThvIjD+sE0lM7OTyxlQ+nuBBj
uBnHGs9BpzMIgL75AYHOas/qVIAuwX7cE+HAbUY6Wv5loSDDSiZ6rZtGK0pOmjGzDeIh2SDuGc0L
dbvSgJ3IWwFu+uhYFXlrIcqbAcI9VLJ/UWgL8X7ue16bPWIANNPQ3zDQNmR8pTg06UCEj8uh8TmI
I+E85OiJ1/2BwOnG5W3VTcwJWQHtNEqoNQmcLiT47iEQKIjCkvkFHXVZDmZKag6Ovg5Cl1D16U06
U6gGb0B+7JJpFGwmaApKEaePwyWKqSiAzfEIOrtmlTqbj2/YPKPtSTpl5trIQDtJK+nsBUgvm695
aYnGBCD+iUxW7PX9J2ZwPq/SvDR1zB7c+Qg45OcYJaA0WSQ6j5jLbzFYpBWGAKWhU9BLhTrR2iVB
3jScrcETqz890DkZib72GASh/nUs1fVfVL9BSNWeZaxluJy4IWz/CNHRMiWWhOh6967qZcxKMTpc
Sw++b9CsZseSp7LGJUJTPzBA5vbwmfBeoIb5m7hl/uW2fPGNy/H2SMqifbQx46i8EFTUaz47s8tb
fqBzFKYfOwxiDpYp/xTfAR6uyW2+xPvnZw+rgJHYoWPrGWZ5XcbV2DpWqYWlBsN6TZyc+HqaTC4X
9AWdAQcJp22EpNptzKRA0Z1h6O54Z7RLwg/U7kI/IVFOG+8w7EdNyrMlv2p7PkFzG6KjnRMMZe6i
2Heiwm/5OMrUZCkEVwCr0yMsKxY8r0eIj3jSNkENb8Co141N1VrNaN9/0nckvfbjuU/WcFlKnJE/
b3WQ7RDfI2bc2yewrXxg595SHcFNyRNtji4SLpqxxWVza2iWCqOfNeNSP2FZy+4LgbmZGZzKnZ72
yAtDdydq+ANn3TXEMgrTv10yUoVXXYaLl+RIV/ZoGFHJ8sTduwaJcbFVYs1YzzyzYhRsnpJMOZcP
qifEvDmeVSfbYQfss0aa5KRDm4fH6+FKK2aHjyPLJjvyjGvDvLxxUbUr1101A1LSSc3BBXLTmsd1
BmUaxFxgG7hoisp/dz7cEs0hO0WjsX1BxdaFTbriR6jxHS4hWWV1nMQgvJXCEReBHtmJwfKX7xLw
OklTFCtB8DOD1BP5anyFvUDqzyrUI+BE/WXpKjAGftdG1ZXotKrhd/1jg/ZcSat1HgN/+8mk0P/P
MpVDcfHyWE00znt9j+0zR+9elMScZ72Bg3Sm+djNVTTpZ1iBiyGcJEDiHgGI94yrt6uvoY3smrOU
wPx76PCcZxblXyT/7xBXPpEOy5lU/tlXISotf+2exTjDX9Y9Lu5MhOBIGQ6atsieOn4NxjebKh2y
Pvrjeke7BvlIADfqaZ6HAPH4+y1qax3otgNnvbm+/WQ9JehoqnrLC3GfKOqjF7t07TLtKN0g/gWX
5xkYy9T0ZhRmUkBAa0xZCyqJ62qBniyVoK2d/dhyWpJnhlpoNsGJSQfyQ5uLr3RjSOHZf0kCUAq2
lIBsZ2OHpaOpZ7xpUw2yqsqr+zvbOJ6LhvlEEPfazQEm0+f0dopMt6oJrKR522A1VutCVT73BVZN
RKIStLcpLjN6SgZVKbzYcDP6FUj84FudGP52D2OZwQDyFUR7pGhdFYMnSF6fIY76YTssUbSjXM9A
hh/Fh1NiCiA5Q+P0pJtjlRBesfIw4RG5bSU80sY12HyRvG+G594u4TyciZdAtb6Ol5zGdrXFbrj4
wNdYMfZwE0rUUZIQHJCcfRvWkfSoTwiPNL/f0L6GdBeRk3dFRpKpTPXCK39ZcFoh6EqwgUyVTkil
dBwiL8JVxiHgz2rBuPSCwiXWg5D1Voxsv7la30o3pOBONmLnJu8TQAcGdqAfwPAd1A0lYCUgNETS
9des8VNNzHWk7Sg3+pOhaG8Qb3mQByNDGYcvpdBa+JxTQVAX4rkvQVJGEiLmpF0UzfTtG8t4q8Tr
jlficmM64sdSSOyITrUAIIkW7NHVkujX29IrnWt5Jrc5hfRFz4yfSxvGBFnCRVqa56A0lTMjrL8V
2/MgUZAb0lYxTvgU83I67J40cDkbLuAsmhq+EzCY6C0FWu/YP3CAaeyj2/xuE2IWaJarDfI7HHn5
Zxk4KxZ9J9Av1e6+XwAwPiae+u/Z2Bq5Wmf9j69AmXegdD10PjvjZfsk6HkotAgNiTsctuX7ad5y
BLVYLiPCffdtYO4cNsawX2BRETM3hEI7LJ9bvNYlD7H+jMjKGdpI4ps95UBdP6GMWGhGl3WfTr8z
orVb/etFVDtjsTEtHjZX9cyPqB7TjK+ok0zeUtY+vh4dvsIoF76NVAzm+TKb8KAx4xTlG5IjyRi0
ZfbXT7V0KWpIY3GQSjjgS3fHrzlJI4rigog9s/WIZ7ZIp2o/p8iYpMFZHJYNfro79BitS3o+vwLw
XmyjHqYAmm4FxJ9zcBKNf7RGNu0Dfndu46q/qWOVuqsI+1qwlbuskD4ub0cTMq2HilQ6E+2D3U+a
HfBl71zmvR6mtGSPVkBHdgeC1e0Fy7t4B3a9jQbUrloNk/iaYOeu4W7MZTxY39w+ExnruWVtUZdW
oviBJaqO7RAZQqbk35PPDxg9wJfBkXDZ2Xb15cYg0nxDhkNKqK/P4fSq1nHaaYNhPOcPcP/qEbWu
Ww+Kpd0sWqO4ptnD31lhgRvRQudYszlbCeFYl1IaA5GKFCWPIC5jtXMwYfeE/IjwqqdDNg/Qh/rT
Tj6siJZUbfkp2wkzdp0o+y7U8XBWJP9kAm7SDzdYN7hvVnaA57oHMbZMU2NElxgKH7MD5sMa72Qm
Gdk+NIxSuXrqyU4lxx0LuztZMmeE8ozjXSnLRQk3zFxm2FQOUSMxczQXeIQZT8gm+V5nByao5b4r
YKqEbSCtqlZwb6L8jTJ047M0rYxneHmlGPCSWFMV2jRA1p/yMU3nxmMqNrgowbqJFJ7asgd1gtBB
IzsJD5nLTG8YjuTTn60GEvyzvRj/7+fF1zPlWy7uaNzrXyjEshOVgOWL8dJ6cYZOyGZDa+OoWttx
cRv/DGMLTF1ywfy6hU0e2BawIi0ytruZvu9rJqslxproJjSWIuPZZaVZBCOWY6xf9rk9cLD/wDTM
1FdXM4uyj53LXwrSbSM79+H/t7KAFS1X1pGqLYnJV4MtLVA+4GrUt7ab3HHkxZD5kpOs0WqAlPH1
SMbj4Z45AHXhT5FedimqBKw0gYi+kQYtFNkGTwDEaFcT1u2m2pA21FbaWxkw7yoR7ratVYolIPnI
l3hJ80Is+FLqpYpUsWSo3DCeLk54Ig7qDja1B0HbS0uDSludTXeKPIUBNtkC0Gu6qRgaz9ytFQlW
/s7ExoA7RqbJEpuWmSXqgi+C+XsYwzTa/0gsiQUF/TD6Nj8+5WsrbbWaDhLwTPFR3uB/q6jOh1Bv
XCm6NWVsnbSXiHmjjfPYEJispR+CjOo9AQR3mNjSPf5DKJ4d8yswixqWDPcmHRd11b0Tf9f9VLuU
pQPE5umMACdOZ8Y4ZKQTm+x4YfBx+gW9zJa7u736vm3vXxQyKOXNnQwmNaA//5D+4apFGkjHjtPu
sk0uCOekMul0QmSM0D4RhNqHoILaIAwEX3eXmF128izpUX5hALADYF4uX7Rrmi/JPXA+KAqtGy6y
8PUGrslozocWdqcpTaqxvGTq2y7cWDfiXpLFe+Sog84gLLsQdCzJ/G37OqnYZwWAsQS8EvO57qxW
XM+JIITw05XvotFMxqcpRT9/MLvRVIt6AmbqFRc3hW9OWsgqZkHx7RP0UuVvvJaOKiEwccuyymnO
OB8MnRdImgWy7AvfBZ9dJ7q5kG/mE0ozuzRBUEU9IyvzTgFPEoTxzdpej4Ck28BtUej4LpTiPpf3
OQvnBxU7aPR6JoKofMJBO1DBdmWBeI3rLO8SG3XdSg60gB9HY44cu3E95MHUbm58gCdYaVtTF9Iy
IQhMSEwWe6WSLZ6dxZ/TO1df05or0v9jAR9oyWqtE/JsMhHnGg10ohMXsT5V6bhwAVgpT8+zDAx+
xrFHrj+qwCQQCP4jSV4UBeg4HXGAOeacJD80uQdFEQ9hf6uDdCFwNKIgkHd+6nadxM8J3gu3EqPN
tgvLOlSHNfrgsMDiIj2qjH2fPRaHHUrGIsPhUO0nWPQD8oE1I6hqUtlFrfpbxuH1uy0B6A1DOUbr
nty/mRwn5kyo0/ITIqYH/IFfTW2PnigXBSKWeVms1SjO47HTuKU1T0mVxYsKk1qNKgQ55twik1mM
1mBjHQwv3AUYNowSSI/QrwxBp2Fmq0csklJ5G52nYLWQGoIdoKqhE2f3PIqkE/hEpRm79+paKwG3
22pP1emHy1qQ1xO0F4pgQZvV3cl4FatVlX9KOYmx4bwLyrrjYBErdxwqlM7kHT3pdgeE5t6SS04Q
PcyCZlVWDtVW01fC89RAZ1+T7bhYrbJSWkSNcukb0bYFe51PLG7ThNUx5KOxZGXOu14tZI3w/r/L
+ZLNKwVqeYQt56/ypX0cMunHNA+Mj7+mY/QKSfQO+jTJIzQ3ZahpYSWujQHBdoMduOwh4ghPZI+9
/97MAufZFdEwMZQhMBRb9PfHbCVWbPTVkqbAbiGSOZyfCZgW4DBGNFBprUKrEAyCTMAT5OQ8wCj8
1AAKKzUaDR/lXS2hLrCyD4hLu9R0Ekm1hm1VTtot7Sg0x6dg57LvWmQ0ctwMzipp7VrOtLX/0wb/
Kjf1hILR8NGrOCC3x2K+O9OaMQ3J+4/DWLOLt0IfQ2Xw8HVAbGNzaGB7YpJOIQdJCFMXhOTUf30p
vEL2kO2/PLOezVOzsghkDhBFWCspv1QFwKfHZY0eF1ZighZxFwSsqPAimHLhkyx/UBWw2GwUAiUF
yOx2DuKIxpcD1F7Ymdl6HBzpNn6Y3OR1RJjI5u2nzkSu58Snd2XKDtOJ/adJbPsPjvim/kM1QxlX
C+xyyd38t2/jaGwcknUHLYIV4qcRA3nhBdRAO0RVyix8NQs9qtCFGPp6zcx2pTqgbCixjLm92zAd
+7Z4Yp1+Svd2JLGpe0CE+Ih5PG9cqgAoa+nTY1Ya6o2AdxiuqCR/YBOVWkO3XmuIVREXGHuSZyWn
/AntbMFleFTZ05+bAQwM85fwDXe35wEwgBif/OfzGHg2RDM0STahj3zLBYc6IwY/Ro8CdduouK/M
msppcL7sqzrNuZLADxk/djCT5CIkzxlFDDQT0m4tMbIGvUqlbaOeX4NufwGrF86j3FDpWlqKs+nM
eCd3xCkzSfb5wy136K+liEjaSuqIceRmUc3ESk6lSfBT/qToH6CxeCJ5arrisGrR29OK0GkNeSuD
hsWvgFCJsxknR6fxK2IKvKy/OvCzWq4/yH9GgiNtmDrcZl52L4kQ4vnBbc+R+MqDvszSN8pj0WVw
2LtqkUsmYNOjSTlmXuMj+8yEd92nbwGS28MOFmR4QyoR0ZCaKGj4zU9ME6MGdug5N/tkI0cpjAIR
Ty+URp+FoZKM7d3WXAZnXm87v/M0UtdAcjmjCNxlvUpd/Y7l/2P/Hf5Vg+zTxLTeiRUvC/Pi/jRQ
ub+TrVlUn5obuA2wGJuImhHWh5op4aO1w3z/fy8L+n41+E0jbcXvYrKHHnU3+KM59nwh4TNt06y7
fejqEFEQu5ocyeQ/H+WRgtgVLMyww0nYhMv2IyUYs6ODJF26Urjh/HTpaB1pAhkI5fcDf7amAd2P
mtqMgb0AeOAWVKvZVIzn2ihGK2hwB+soxXrZi0ItMupsNU8Cu2Arz4fEVw+LyT63YbmcV95qEml1
zp+jy9/sQYJvMofXpaJqUh2uZ7hDCiCEDsO5wWuQa9M+K4tjSJLhUn1sX6WAp+nrNN/ul6AJNyjK
VY4hI7IDq7l9Y87M6VbrTyLg+TYQWUXrQLMVSr9AsArbbJuvjVOSNtjqU6TOADLpItAwv/+VZ1Ne
7J91jx0EoyfGQt8OuAxpVf908eqS9ZqeMcrxKRXwyTLPaGFAHY3I2MaeQZp1znLQh9UEmIG9wL6Q
fisi9dY/gVjhTTTlqQb/bMvI52EH+n4rNC3D0Q6UNCHsOAahhdTL/zwfmy6paJOndfwLxYYjQKg8
j4cC2gG2+cs1T4Z8wYoB5b80R5MG711lLX4wnXwf70nvXmrAwSE/gNrKAVhCNWXzb8Rx0FKLiHm0
A2cYfKIPD0GVdBW3NuC9Md4m2bEVHIiWsBf8j40Uxg7/Hds6kRF7zJAHJ5MuCJhXbKTus6LNWn4T
EDrQg0NpwjGcM9jsOw6VGs47FjO3JXxy0iQK7wkoIlxDk8rhi3xR1jLMXbB5p0LRn21NcqRvdbLk
W3frxkm7guVCeRRFdFjp63ye4vqicz9NIWmZJnLBog672mqoZ0qxeHQKmh4YMiajFtYtDFinsNam
55WhoDpKatbTvlh1wZmtYnRumKswGlM6DQqx/zoglUBSOl4C849GbWoKS+f6SuI1wysw+YcxToRr
ZOmWhLn7tpfKFErKxhcG1x34+//OtjX1OGHK22gIq4FgFVrMqs4gMNOWG7+ZZlrMY/X1wetRzF/9
oAwQhAzsvc3D4YYd1bkdFAwtDWSmTn0jA8jCSqr4yoALTDkzw+zJPOdhf3BoWQmEOR/Q060XhlrA
uEr38blg5CTr15Mm8kZVXYx2jHuq2JnzyGSTnyoHyFsP+U8j+4+kYOBAx8uz0wdlYTbgHJQYxl6x
BIBkJhezu98RP5A+jY1DFHrSPWqoLmJHcmp/i7b4QsRvWMVaymaGSwEaZgAcrzxiXk8CeIX1lMLL
acqgEtctg/E2GZ1ISZtPEhv1zUgVWhMD6ICbA0EznkacIKQuw9uTyRMuXzrOZHUOeapm1pOQJ5rR
j+CLxaevyolfoEp9rr0pz3hVhJLOFW6XUcHa3JEj0D6dlp+O4FN7/HuJFUJNidyPiStBLaD6YHiE
nu7/xVsTlgv84lkQheKPfKvB10q8URS1ERdo1ZGbJOUp5ICvw1y3L/jFeP19Z7r+J8imLN3u0ow5
E6s+RyrmIr0DeGl5GNF8Qk7xzi7w7U24p+KYhtUqdRJVfNtJt1cihMr0gIzdeEmfoTUiJvrMJFIA
Z4MD6DzV/wcltiZqySoGfy8jIVoicFD0Gas7Edrh1TVQRMaCXnesvKUZymCjmQL9wxyT+xcXxQ9T
oH2oxKmG5FkUArRZBzEe0fThTcWyMg9es9WBZ3MdVe1OitgyofgqbF61hzXX7TGKvateymUEd0uy
pTRk5zLk9hXJHFFo+piIyN/r9/oyjptGdVeGyVOaHzXR16/1krc1/W2x6nhudJbCoJk4xyd3RTSr
F2wJqY+UzCQoDbSd0y+MUWNmYH4gnyYvAJP9NCVDC0YBCD+0he+JgcIG+JgOtuXNdXFoGHWBlm38
jnOKLXGaCX2uKilqZYt7n2Isz7PZG91jfUe0fSPEYFw8appTbGM+LpRb/dlW9lCNG4D1zIzQrZIb
ariO/fJnKnst6qbgGdSZk4NUpsZeh7aM+gJTq2nb7MSz7ON7AVAqH2TCBs+iIhzgx2d43q7APzIS
6EDM7iLcjUPVp5/0GF01+/90KPjFFLZ9YqS7pPEjvDYU82AQkf/mT7CVpkNY/Nv2V02sjU0dCe7d
SAaEaP0oIvAaBGiYmo1Jw9jt4mVENda1bmZ3UWIBls3xj8AKX1544DGgMb9LByzr9TjzPu3gs8bK
dorg2h8B6bFvcWwbd4sH047DuFx3e4gfbbkC+wdNc+CaupeiWNrf1Y3/ZdYZJ3TrQP+SCoOLQAIC
WvgGJ7VsS61EC8QCPcEbwE4QTDwCmWtComLDMuMo1QYgYUBODibOzZBOypWXsEhJLCLEdydxPgk+
9nyniE3Ir67E35Uyzpslv+HedE870uEuEzWtdT5tGlDbDd+PQSURlR/FxufBpkwK+5vbbsLZ5j2e
RjdwsQWPWmBM2Ttjt7YCZAMwY/osdlSsr2DMZvkEdDPOLzeI41BLLRrLl48uwLhTlt5h7pg0TQ1e
vO8sR5sD7+O+1kNuoEUPMrSO9nJAJZLWi6Z9Kup/EARbs7QdiWs5D580o9vy8oI+8hNnVQiviOtp
BX9A7QEPKSvOMPF5sJ+NTxccYXVeJ+Fdv32BfECxCxfAk01evWiQsNvMvYuIbby1K42iujnVxDL7
Dpkv7G1vlAu6Jbidsk+v06IOivT8aldOwu593lpSzFvkSJktLhPQ5R+pQlva3wVncegjFTi2lEK+
yKcUjxQqEm2hqgiEAszEB1Cci4RmyB4M7zWlW6GpNbX3nYGhg1Be8UR3ac6dJwIM5kgekRRDic/5
hQsquixaYT9fsU6tpGnvgDGO0glqbjRtAU75Xhe5GYxaoYgXdrmrT4NlNvoI1PMVXYZ0N2WVlJl5
BMz6Up0EkNg4iYiAoTauncpnugSTzFYVzTGkyTHNi9huIP1RzuflKfQs55x64SbPuwBcLN9RK7hH
nTnjHbKeBsjSmyvhY8d8DneDzkbW1wr+BVUzjR1RcfLD31TGWSyGJ52+7PieTdDq1CkSZVOjLSeV
1fLyvR+Dm5NdwiHFh/Q12xBVcAkc1O7/OOeyEsiWP/g5VnB/bvhNVciWIjlWegP6hyQjtS6VN4Pe
YrQlRJvjRJ/w9BBYkQ8J1+NYHSRu/mAxH1lzj4P0dfAb7SXQBDn5uZgCjB6JJIhvVYlxrcN3tfiq
hQmiO/oly2RySSFGoqqv53DxBZiD44BDlpjvqExL5OWUaspAXMJE62zWuhU6zXgz5nlut/Y9z1h9
ohFLTWX9MYCGAZLv0havpuL61bjpQq98FKb+Zz+74VicSyrHUk2kD4huwSeNiCBW/2hwNl/kK7RD
M6Aj2E7JiNyB8tc2LfiQZdq9Bk/KyTqiLKcn6Wd142AqThxVfKF0kQZYb1LSUQsKnHUENnZMJGGE
rnJL+A3oSOyZsF7819MHfCeerLJ/R66vsuFpwZYwC7ASo/mC9t4gBQxVzkJSHtNcGSNZcMGx7gMN
6L5g2S8bC1q6maHocqp9ShsNufJAJvphyiYwqDMOW9/OWEtG84jwhS+/OY7oCNhS1GCOht9vbVso
Z8wMXcsmxtZlDyi75WAYhfSAFezqlZsImjJkO9iNmo89lkzqKAh1jkf2KOSUFa2agaHm02XbXcTx
m90sa6/VCiUwMSTYVzf9ss9FriMfeSFhxX8ds8zD7c8MUWJhJVqxilnBQYIx+GSNBu03m/yMvThW
ZkT0Qtf0WAQocF1sn89CithKIahhJM9UTDUZuueX83yWSipDVOooKAtsh6kPLQqp37h2SuUFA5jx
UnwoOeXkYyMCMDpH4/P4Wun6/WbHoF+m3i7TdFSsdFOUGAj9JIfFiD4Ud85mLTERVdDwhS8pPGqh
q6P/EEM7ESAPmmLuWmbAPCzejPPoLDG5tZXsHPdeJAOXbTWOWOAtoRTIplVhBJnTtMmQjckdLpFN
mrQaaZTh91OqgoCHZtoc4QsKB8zOTrb9oBFQEFKK1gptN2nk5h9F0SmhWTtN0QiYpC5zJ46XmEvP
4sRADQN8alQoUFvYGcuolT/J3qG4HU7rc3Upg4JS4b8cvvjDSeSAUq3z7k/C2IuRbo5Qnk+bh0h8
TpHoO5zHXNwe1IC55s429wkyLJjrO9gCdzXZ+YEwdOJ3OxJdgcxu/fgCqkfk9YArVmQKUFaX4yyT
W9tm75UQVJyavwfNmUX4e2OZzyLTOgDFlM3EAc16vW3PIFMfJRINCelzP0oFdTdx1fVxZpHVxWzz
QpvmvhZ2fv8OHGunLZYwhhxgBGXQo4GHOrm1hp2u5hPRAb30M6hMeNiLdvRAdOraHlk1eTXTfMu1
cTJGj3WPLx/pBQckk8/Q3UEUbrifhZof6KXgB/5gtzHaLAEFthw8hqKgqFYqYQ2z+KCqkz4gTRl2
c4G5RQs+yLQ7Z54mGZpsEI9BwBMQ/gNjRVqh9KuFrR8MLswWclE6ZwWdUjiaFjpy5m/JE6j9BAaP
Ju4chqU9S0eHsaldVe1L2GlawHif11k/YIYXli0dZf39glqYNrWtPNqdsPQV+h2d52REN/SCzb86
DZs/UlvigpFe2GQ9L4Zo/lrb0Cr6DyqWuyABtJjLqSgyfm0UAGBLKnOw+PHmjUHFyZKfdi/poE6R
9tQLXIkIKu9OWDoJsMUBkvfd5YBH0cR0ZFgiZWvkZmpXAr/w+f7zKcaxCaaADyX+oXxNsuG1aQSX
sd5NdTgq33m1qPjiLehFy4kwvWxwLqKcoI+2DuOgYtYD8bPqzzLRv957PWTGpDEQaBCaaUJJIOwB
OOfMahnrnczevVS6D9zX1Ve3d648LH2PplUvDXp4G8M3qKPwwmXxm5Sla5D9Fw9VDRM+DQe0XOSW
pkr7c1e5/F5nLZBJVmt22Z/f+/gkpsc0cwuCqumACN4J70RMcLjj9LJ6zPONRUnkLWS4jbEA6ban
0gTKfvixlrzOQRIgt+1rQqm7sEGP5VIybymYshqa0T3FN0Y7LX+XQYMyjwaFDKooVOnDh+jZJDkf
S9V1RQkaska4Oon01h/LrViYFyDdWLDDlRO0sxbyFEri4axQ0hYaqNhiHjpTg7Syj86BaUVMnEw7
UvgyTl5usNVKXzwAWKpmPY/QUGrZgxlnmNdnPvL9y0HhhOJxF//tMOo2J2r+LzUlLFvwE9FZIM6I
YIDkkIrGBFq3gBVWIKiMuamtCjpUMhCFM2ot0JVP7+6RugpZwl0QZq8b3xNx/61Dt9w2t3K0JmJv
yrsG6sx6UeFxrzxlp2WijNlFBWHOtmoa/tbxa3G4bw5JOko+2mddQ/d5VQ4JcxSeWFLMQMklLAuk
jydlz6D8pkfqsJTNO036ihpHuQpOhxqMON4DYe3S4+CFRfSEyGA5/nSrYuk+weBlvhYOpZopzxzQ
35n5f32IgGaqZjmlFZfqM0+PRsNuC7iqYInZ8UtnkZWaePaph5LHcQaQy/YgUd8CLEGAu1aBUr+z
nAvIdFdznFUlWzU4e69CVxhyYil8TiWZy8RlVe5yunmpAaR/LvhO+96WAsWW8csDG5/HLxvOqzei
QdPiOlR5ZqwjlBWxK6fXgZeuWgFqFPxuW1KqBAPt55pnC24QjXqnS6EfdxfOcjkLLS8WSGRa7bGk
ytTphTjABfGW4gKioMzW263ayONcXuSbx4BUC/lReRxL7tMWha2XZYhHOP9mjEssP+epj9BaLjRh
c9mae2/8MPxgixdBccX8JHj0TTxczeqZRGasQI3uiLFY8vYINLWpKtgQZnLDdwv95jdvPIA0DpXq
xugMZN9CP5L83RuyIou5mvW1FyZvFV7Wf0mvzl66uiwvHFtMM+02N6EqgJKRRFy15AgHWMDCFddH
VDKtvQZHqwb04ZwjC28kHQyn/dnZUcQaDFT/zKz2kNa/RZP0QznFvyJ386blJSywrMPXco5fkfV+
/PeAXv6PjTn1tUcTBwcSdm6YtsTe+14Nzte1NzJU0e3x+0lgfRN+DKoH7V+5CFaQw2Remt/+kOn2
eQIVGzmjtJtRWgRD1i2mymNIROycy+vUbLPyubSMtrayRU8rM2fRVvscM6uwUr95PJBkRWFB6Szr
TSzfUteQm5BvLfe0fR9/whu+/wJOU66/yb1901/I/1AcJ27xOZZ5/YGagEVmU9SNHN3DtqHomqxT
9A3dcwIEmJIwYWEkQkkjJd0SA7WfqXLOAsfHlwiAzVVOs4kQGOQCzBlWtWjSyv1Vb0qUhu1IT2FW
BRKBYW3r7LJLmACkNyrMydl2BPGmvTMuKsmx60eUY32geu3s4Prx3aCHt7hGK/120icZbjnUUsVy
uzbE7X6lVFG/eGkDOHqLMYVgTXwDTtusMWOKv00q+FsukT09OerY4kQrRADttibOFxc8uDGGZAKU
nFgsNq1SMndTsgBeaME7qkEwxj+miQzxKm/tFW8mgtIurMe88rj908YHYP1k0KxuSQcdYMa/qdAD
xQ+vSlGBaHKbXpmLjYsAImzObn2kVQ6JQZnFNZo6k4NJT95ILNFxcssmdQqUJC7GVnJGmm/9dYTK
EhdB4jrOb4jwwD7zIgGbzY6P47QYFNxDtWlsT3Y2N0ueoQfEepNWp1M1t/LC5bWC+Z4G4aE9lYPD
ALkxQp/nRwgFQOMfDoH+1XpzmT8rffrb0PB3+hcAnAu5W5A12unl9v3QYIoh94oocy2huUhJCb0L
BZrq2xozNVpsi9veEy3+hteGTYnGYw7Zu4/rC+QXdVa7CR1OyMu9lgAI5dnFrl34IGs2QiXbhHMy
yqlJo5+3Vx75sxw6JWMPfUxfvqOiOfPG53/5UmYOhZnxYuCXjIZcN0hwq723VpIr2TtzvD5RI4hQ
vKcdfXOvydhglklWJ7FeLNw//Q/E5rBbWDM6smxHVYDwsq5E17OzRERwSUVm+yt3xCut3fqNlZDH
cd4PtirkWkm017cQ2dP88caIgyg+7HZxXo7Pm7Lj1ohAfePF107CqpniWSUDfwNhK5LWlIEyYO0v
l1nBKPwoFPr7e/ORuHBtSwEI9IjLVgo7YMViiAdcHUiTR7Xa5aTaW9kCdtHOTzHZ9wmzKPNc9MC9
Xj5JGarGm89OmGB7FXowQSM2tRE9nGt0F5aIRbiFt0nenQKUjU2fYzwz4uF02dYyM0PTl1jyFKSg
oP/5Tp+ZPrHACPA4Ys2lKhZaN7uOtepL3FKCq/LKb1I99nFTKlOTUKBdX/uJucEDusuz3lH7v333
wMyfjE7UOIuNHui55ymuCOV7VHSclz0EBXTPzU2VwGVBb/rNmtbITx6LHC9ygRAi+vJcYJ74ni3C
8Esf0AY1xOk6oAQizMb5Bqs/pqkknpFA9XIGUGRcjPJlmMvF00x1oK5ZJICsbxuF5hIsalAhK2PA
U+/LVUFFA5yGWoRinOX27kJMc6JjCSTODnfdFxkblI7sMELM3XE/AotF+vfI/UGeXZunOw4nF+7p
fGov0RNOJtLY3WRe/DDWQN+179x5P4NydhFCT8h+mdWz9uByqJksA6ktmb4ItPYTyIh28KR8vWid
A8/WRzl2uJMwhQBSKju78dfbwo9jOcbiCcPQud5RuhJDMpO9IJ6Qq3o5PPYJX7+4u814Cg55kfhG
q1CuiiasdB0JzZwJ2vvaEvvnN9sXf+ZUDZkJOBF6LgQI4AJonqY1A6BkWW2/rtSpIJVgnShifHez
CBkU0Ej1zoLOtTV1HAdpCjGgVTyo7odXlmUZ7ZGyP5W/QRnyrvrfl9bEy5/JSazI6CjDd+e9gy8+
IClgGT5hheR3WWmLQUHiItCZLxkER5YGd01AvgqGHi1SbhB6SYe82ihkIs5J3vvpVXIkM0B78577
NP7ZxtRatoo/vQVQHzjfVjJxiY0zOc/0e3EG+FFm8ICqDRGFSQgX63/O99KE5aRpaaAQu7lqF0Iy
R0e00KsI5/siCi3CI+LFlCaQ7nytbXr4idH9r3vK2MGkCjsDx6h+ok0NaMwLtc3gl6D7bZrq+8W4
WFEWofeK8/x4KffXNuzmQ0nfv4HsdpK4DBS9f8vUvKlOc80s4oLKoMfQYjYl9Rtx7xUKqNydSH6U
UReIvPDCWeWVofEDw1g9G8kmsJdhir57Gw0UnLQwQoxMxBd7KIGtGtr46wUBvURPD9suYF2Qz+L1
DsdEMDQMPSw0cWmwRy8IiKeHnPltG6W9JmO9YjogqphUAqop3VY8JG1kdeXcBnTLih/k/G3TwJ3O
pHsZUPQc+4M+vkk63kZKU+WLl/faVmE2vz4zWeUBXgsAW8/zPW8Tc8PlX2yAp9dG1gC8G++1TlMo
ZEBAex9Qfe/C5ElaN7iXPCx7GJDwB4PzoX8JyphIFcaykNAoV906CsJyzuXxlAn7R/LRd/Nwmlbd
1T/ABnOqylZLdzp/lQursqrW0CaS7aZzC5Llgl48JdH+IKxj0Qp9JH2zPxJ1a9vGDbHrdK5MBdzT
aA7lSwnRoqodxq1ek51UDGDFqWiacsOKIJ8/E7U8csrcnQvnPnoAP507C1gOB3lqbtJp/Zp2v+c5
mBqIV+oswrJuxhToXgKOCR0ulzyaQwNpWwxSK/L2MzkwtV0E1Lz0qN8ltb2HRWRvqVa6rjDvhbjA
P12hpLpfw+rZizlgRW+XKTTO1dBw3SyT9x69lyIR6lADDPHAtUFiIFiakNxlPuQ/1xXZDc3AUp+A
umYpPFW3RmQNs9Wgff/9wQktyFRfyPr0SleJM2RGshG3/BG3x5zOLfMungcNUVyMFV/WEmKtGQyE
2W/Bp7pnHb9vgR/CszLVZYC7MyG5TX8PaoVvjnKqzxcDAZmW2TIim+d8KEuQ9x8W2qPtcJlcMQGy
4z3t6qp/qOFuiCL95jZb
`pragma protect end_protected
