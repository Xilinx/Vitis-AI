/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9U1pW6nshgzu878GAv8tCKvDS+jodeKAX/6BGZhdnC1fBBUswqyOn5GH
yCM/qdb+7qsTGhmFJubh7E+FuAwTUVVZ7UX3pF8CEyPwZPfaaq0KUfKbnw9NyVPHS0O7qnL9XvW/
yT1dDeMrunwp9u7cGF5cufaqsAmcVQjSCatn4VAK7rN7eAf8y0tZgzPS2+MD5RvN49RKT5EfHQuc
jQ+o256hv4En3oqwv560FWxLxfNsINpRfO7xE09xFz/OQEKouURVoWGcT6KyFe0WaVIQ2i711CxO
iALbdtDYHxO2pNrwQRdrTa8ZLJdBS6pfz9cPOmdJSa6VVxbmU8jbfV8mWQ/eWaFweU+bGRQsBNmo
fGyeGbP8rXnnI/j4CbPBR1P7QwfMkqNCFhzWjUaBCOsa9lNhceYtJeWajEPMm44tO2aZEgMbfaBE
yECRobm9M4GRurexZxnVAEOUITNrWf3c2+5NzqBRzsq6/WEaSeokdPII1ianhrJF8uKiKwiG+50P
WPNjO8zf2GxO4iwi5CLSX1ni78r8U3J8vCUTyinUcjtJEdvx5N45+K8gMy9tWrt46kzokz+4sZl2
D63QGnzxnWthK/xAcx0ie2y1AybP7r3fb3wkgeCgzY0ezYFqlLjAQvCxqDo0Bn7W4gH2iZeikQco
ntmNZTDrOrKMJR5yVPYPrB+GIuZFWAV++6ApgUfHMgVc09jgN1wCUiCPlzn6hZX5VoVhTQoWTY4v
AsNUyIIrMw6qMwiDXy9vJWlNpgSWLh+ggYaTR+47Vt0o62IGcmpVX22/jGZZBkPKwKclosLU4883
i8xSznYh6nRf1KDAUHO7HJuzwPiOrOU5e92e/iBV2OJIf3yvW6/WzBkxr+RrKriEv6y16+TLkl08
fkGGfiRlg2eywTf2N/1vF0kas/wNSAQoqs22jEt2Qi2cWQweAxvfHL1o5lSh50UX16bcTzSd5Pvg
o0SG9XFVFvvsdJooGJUM+yKvPYVertv7azf/J3RnZUdh88+YfezvNIQywVIpOtKz4Gn//guXdeJ1
TXscziGU7vtR6WrbhaZ/IVGckyBCrXPczzl931aSndLYH09bc3j5fCYlud0w+F1DIlGKBbiOp6l1
mknap8L8jFCQCi3zhbUAF0Dg7Bty+/Yc2wbYciVwY/6U25Nv55TmiN7MWxFmUw2fDvcjASypb8by
rdpdkEHn03rLlqEF2IZcGlOYF6ctIjYLP5O8dF2JQlkHO7+jMkCqr+LwXKtbpz7Yr/FsxWcXrun3
VDBRA6Ht2V+TR/TLhFIB1Aynj/zFAI8d5s3UUPGtQA1P1ZtAsVVLeYZGGNRBRFiXfDRploJarE5g
ucnDeGZwP8TZyyykEcxGZ5Fx4NQXXesCID4CVM3sXTRiHhhUmjwqu6rQN7LWmLoRDbp0vlMHRb8r
DEU9mGg=
`pragma protect end_protected

// 
