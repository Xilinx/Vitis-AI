`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRkcajQVnMQxKjPBaLZIaR7/J7zs
kEF1+54ixDuIyNX+QBxUIanAUk7iqIQDed2hUG0kfoXoL3vuow/GsZ8M3G4iHfWrH7YjpZpxAU7u
+39ASljNjmhxyj7sp43zFjND7KB7yDk1EnS5RQNQKgSwY3fvRC0feceeFHyy9eiKM0+E3KW82xi5
RDh2XoenLekPW3PgKxqpPoG+gCC21CBlAB1jyVhu5giqGNu4bAVf/Qoyy4ljAhFmoJLCZWCvKUsi
ICuOJ8aVk9B63NV/fMMZj8xXYg6Tu9XQfx//1S1e1aFKgVKsCqrOQxVqgXUDtON2Y3HoxVf27D51
/MyKlVvp+/wZPJ75oVlGX0sgYKR6T6Ld3fvRLmqrJCTiTr7wttblABbSKmWnFlt2JC93z9nkpXGz
PafzZ2oPBmKaem0aQmwbZi9Jcn3cXMOXD0PByOYYo55Dzt8NZJj+r/9d4TOBE2nYMw73dvdfw57L
URCOKbSSzcfo5LlZBD7eT1rE7GzM+ud91Bb/JD4J0WtAnTz60gITRVNfUEWta/EZEFTiuLBI23Us
w2+6VviY0+xq8+KsfIrD6lFyi3VeIZli253J5PyNyzPVCRe4PvLccZ8DXIk2ds7wrvn3CpgT5Ycr
L1YVrmWItigeBi1j9LFJU0iwAp1uTqOMKEhF8ZiFsGjQvFZ9zo2xV6UyipWpdTsm7qXfSdsP5q8D
yJpr3j/ImVfzBROz3OLfzvsHRu1swDHrobJo9Khf59efzPv0UjBM5X6mRh+GCH13ElE+Q/QT25AJ
V1tf6YqSzZYfdxW8TEOgLU7FT2jVaDRUH2QPduxtX24jbnBAayz8ullB2LnlnrneblbAxAIoRC/B
uQUux1OiXPcj1dGLLIliSvnVko5Zz8lI+9BSpCji4X9oAt9mf5pHpCkLRs5xAYyVbMdQKbIcimv0
4vsr2L+rnwssySDbFxWBmj4ibHjwaB3KOtl6jPOMe+NUhgG8FYEoBMdiHi2qtIVRr4GZJn9invgy
KqJaLOYTo6cRAB8Ip84OeYBi9sDZ/2qcWCUZDm+NYqCeIZheDeZZstjTa0Hq6vkEUwY1YZX5uDiD
BtGgpXRgdSsyUJujvfDVghDLKrWUGufksLilxlJb/n3dcQ/CdXl9MM5kh+k7b2Xgb49t3sSs9u8J
dyXdu4rxSKtx7avU4DvCqeFhbfQ5livdGOSTQMiRroM/CQSLMzJ7k9oAgrD0+rmmpW8haJ7G8J+i
d60qX+NtWkFsoTcaORC3aoCmwwadcQmTpVMBnMM4HsZeo9TvwVhovojPWmG1Ae00AwhQdyPHKgHp
NB+081sVk/xsX+SJ2jc9P3orARivg5aBNv6Mn5Jqx2j8z+nIDtI74DIuHlP3w+qqM6tfvP/vAFz8
Uf5LfTAJwp+hbnS+Y85H4bqu5BDZV9MlZLOivuIyHwKcfChyrZnmUv7zIyXfZaA0nTW5F0Vq6osf
R+lGp8o9Tha/d1DsF9K2izBL+la/c3Yf5XL9uV9EumkLR9ynmcycFyYS8eDxGfPx0fErSo+BDOjs
sxHMsOx3+92PgVbx4NSkuT6usyIiK2nROO0kiHO9kxP/E7YWQnol94OTZ5KtYm45aaJghyJJBOBz
4VxjVn0E38v64R9Ceclpbykfxh0awp6wU2f5h3Y5WW5r85uyNgoj1P8wObG5e2YK8LfihEC58Xyp
iokUf7vanDeFZIflbR1dVpzMHwTXufus5EU3WzBJNt1TTmm2hF2T+6RenZEaswS421Z1/kEJYqJH
Ik030BqoZ9uJOJugzAEf92rqZGTlNA/XVyc6O9byZNUADRY67KRTtSZ0GzpDhPnwNUwoZdyxPEFZ
G/XKy/pt7hE4Dtx9IXENS3ETS9HI9AEVxIHW5P3HZZ3AQs1jg2Dp2QUpd8i2BoIo4RbZvxIg0VBy
Y6J+uFOohkqw7Qxaa0htdk1ugn6ZfD6wncz2reSIWCSQjQs6PDQlo+LvhltdeFvgXO2qG05a87Ct
yF5TFoaqXKeaB+xehmOVWMHVeFdx0pATd0JJWDLVTgT2czwLLqEZZ4wcYH8jjAqyNcJYswxp4o1S
Puo21dXKJ6E1IgIkdaNQEaUBa/lU6ZlGpqhoI/uccVbd/t5WtobIabyZRyleyKdyZpl11FAg29h3
QsY+xTqUU6Y2oihkN+p1Ju0Z+kWJ8eL10INgOrkc0g5MxIYxwiiz+Af0LxtRHFF6jyW5x02ea00F
oEJ4uw6LWvM1WqMvc4R4PKdHMioMRMwayYFicbaAGb320YDM0EPCmi+fuH4p1tyboXYLMUSf3JNr
UKC2S2NFD1D0m0wMtU4gCRmB5CdmswJQaU3n0Ctr+6MVbtr1DO+Ky8rmg01LrUDLwYmBVT8b/4Lr
y1piq1TyeSCJ8O1gSPDVToxDwEr5CrlwO6dUsAakiQTENXp3irUNEVtlA3OxURP9IG0X6gjdxpWq
QSUr7W4kAOoO53QRa6bfrGjVjFzrp1kn7GeVU5UvvGbphoU0NeY/DDsNSkv/Ht0FX4x/cph8zunQ
PXb5uLk3r0wOdbMwIZoI9RioJ9FIDzW6oq7NFwDV51UtbTQk/Mchc4e90EjbwsjQ1v/vSplJuoLq
8nogpKJP3bdnM6n2T0BfR2jxTcBc3MzKY5eua7lm/xMNWqKGv9sOpIOkFmJumoIA67+C2Yi9wClR
/Vanr1ZN5lrtaacmrzRsfBBt0z7o0CTu+Rm9CylbjjsQzOWVIKoeRXPvNyyKTdJVep9X72rKm+Bx
/6KW+9VD1bMRnjHVeO+v2ZfiQ9e1VbYQwInxem7kA9QKyZksoldkRntYR7aq7JCwnKtOgiQvi2Xg
FPU2scfj881mE/oE6482cYD1zQpOkSpjuAlYld6xEd5AVm4ENpzuWLo46JEtl3vDxdLMkIDlyQU2
UTE02FiJbTyGKDML59BvV/wASL8Gay4UDRNndo4GQVJ1AdlGRttL4MviTX7k6NZUrJgOLmhB6VdG
QF3Nt3XnixlDVl5k2yLL+OmfT0PorAjMAcpY1QQnXqr3qnufiY/2+2WYqzm7v00+97phM5QUiHGV
YFvxD/DmkX+zY6cx5z8m1NNjcpT0v2AEWDoxZOBhNyql64pQU/drjFLfju1sIZ7occeL5gWqczF7
tQ4T1Ly/ptQ9FIkxorVSGb0wH8qmRcRCSVnyt99XxjhUXMexzUmc2qEt7YB4+B3yOYeXDhVsp5an
NUqKW/e3Fsd6wKUoHxWY7G3Ib8CMSydpBFGNWeYzPQRs39WbKpK7GTZGHtXHminUS9Phof64AnVT
Z8/t5dJKar3Ac5NwDtGkldimie0eIhKOjI8dw5XFChHs7S9LAh45I1sUsF6F7yROByJqb/Qqa0dR
krbv13NWQuTOfLHZMo24xOhXCS832knu1RTGi4IWVylxy0YlWGPUI/Ruv3DW8N4M8WkXUJ5Y1WSF
M7hhpmnKlruXPR37m5kEiZm+FMSifFEmwHITZ2pS8rY6+vge6W04SVKL0oAyKqwXVe6G2uIj8amO
hT34tRnYTkQCJe6rk7BeaDmYPqfASGgZt0r0xbogXwA/DicbPksyea0s5pXHUaX8FrH0mDrX0h/i
tBNRLVlL0psmyxaNHZ7ASnPPGacZrMmpd3aW+xmVVqtsZHMMN1jmKahu13mRshIpEp2ULIlm/ccZ
BMSEGhEwtfQ+hMdSqggcNAGtfXh6Z0Wh5qAbmH3Im5/0bTcTkPVXUizz+tOTp6Qu/67dvrV6r/kx
txMtl7Ayvieaw5sHmWhIQ61x4X+dni++NTA1hbliqXE+M2XlUSvsPKZiQHSbLoO/CUwSgWlHko87
iTqTU+RcB2rkguV0PDrEYGfgTH/Fo+B6XzsAhxY/TDKCuGr9vOZOAFF3SXa24UYZmIwQ8oDOJcWQ
cW/iWgtNc8gpUH1A5E7Oz8tYOU2tuwE9P0IUKwvD9ut+GvdLkFiAzTnt+8tWmr8zZwXUSJsc00c6
tqIrlVhSihQKuoxRhE+KcbSP8vtJdCclqFv9xXhTwJ+KmjEq3jJow5fX4qqi5dtulRFsdCsTj6QC
MEERA1ZJRdGwI7zmq9W3MI1XIP+BvPotpkwPnn/u1GzjsssKyQHWBBHwZHGa9L6F2LBoOzVadq6h
+XREqHJTfVtsKbB7bXIbQ2O9y6mOe7nCXiliCgNEKyvA2+ZJUBaBjiUViFV/gjgEo9HnVEPfnLJV
hWARZ5D4gKoMrzxfNrOHUxbxW0lAU5G2nJglL7+/H46icQG7IuCR7r34LEkMofOWMBljSLJwHWWS
LCppWQrXAohJ2tGQicXwk9o8tIZgCLPJi6G1ma/1Raw8Hdurg1RDkIlQhX3Jd56qqZCHFbw/aZ8Y
3z9e1kVS/xmfKn+T0841fjhDGjl6FZ+DG/XQxftliyVkCchFJutoNZ37Mij9AUALeqgd+XGh38Gd
tQc1Of62uCz2xJQrDaaTjtDuSZs9YkWHB/3UMOockCSJT5pVFrhrtfiySUkdKV12SdLMnnyNKcGA
+K/QZ2d+HzR3j8Oe2U5gl9JCnv7NQMjolYg1bSbctkW91gty/vcYerk3Rv2dQqI0RWDawn9Kz/74
OrB/qQTQH7xEKnO3f2HwUvKP/MwUjdtmvz7YtcTo6TIi4wy/Ojb72pyuB3TP5p16ISqhwQ4rJNJl
polRXNb+HF2Fm3DTfSgV3q3EGNGZFTnDxJYbeI+Q4NXc1rRbYhMioyc4lX5nQMJDWMtOnSwSsKYH
NYoAQoSA3AVoHRTni/Y2N7wga+bTN5MoTt3+z5pAWCa+P56WStbUW/BfijarlMQHA+I/QkO5BDl/
V+L31re0+8Uv2xA6P83xUsRG7fhZNme6W5UihXDy4OBQxdAS6fCjnVSeaB0XDMyDO4YDNbKTAuqy
x+vQCRCw/XjnYvBr27elKQbvR+3nw27X+YhuxetibJghr+OMmi3aiQQ1pyVRv6kN3H8p4+yqhrNv
Gzo6yvB7TUPLU+79qYSzh4FBxvUa38OOzz1c5u8CtzaJ3SWtPtoY1NfFG1mDT1FzSi6MMtRYCEND
UP3yBvC21E3OgkeLh9lW/vT6nwTB0BGCrJOZ6CD01jROGbDEeA7mc/WNAOis8UHUgeGzYz5XgxIe
YFnKdygKTidtnLtBiyTHnLB++sd9JiOV168i1mDndxN7MXffdS9uVzq79qRK15Ae9QBap7fRmQQi
zhRYVOyW2/bu7xkNpSmUf5y7TOm71eF5DASmpdWLn95pogxz+a7UHHmyS400VqvOeMcKpwkVeUYs
eXoy3JRYfQe8bgtQEVW6LH+7TEqpZMCHLCUD21h8hodUSw7ClTihlDyYGfpctZQQny0bSJoQdEE7
4Ju7uJ+0ijeS7nnK0YyVKTMtsGgo3Hjua0yDeM+T04aoPpuckR2Ja3Mbq2CN/tO5KPqbMSxIGgOz
lqhYvt1AWhqO4KVHKe1BxlCoj/eGNvGJWCb0ZebbN3Aa0RW/5jHZpNsvD4SUM4qveqMSpvLTJcQT
O44fDf5OVjgdWvC1hxSvQpJTyIeBRDSd3s+xKgnCYDS2zycQfg86KpdRXucbIY7F2AVBRa72RNZp
Ru7fM+6M5HvDP7D6oW8jSGLvtVPDcjINTSrVAAoaejqLXcDge3ZF90YPnRoJVxQFJnGlI1Mh0J1g
U1NZ8jANQhf8dQnki0XJYVy+m2rf68vBR8R+UxeRQCE4AUQchnL4+F4rJqcoUER2KGD6XuTLi/i/
0uzaNNZ/wHjR+wFlvFnT4ScccmDiQ9Zbp2J9E/MDaUgCLOHxgwex0Jc7d2uMPymzYIBJFS0fyqjE
Ea4FC2Jp8S2V1ol3ekaWX3opIKbwOyLNwLz1Owp9WOx+V3Wj+mlHaSOb35xqRyjAh8nYbE4w5atr
McvPk7DNeWJUTvcfKBHhpTuKVZ1SDqQ7240TMBTlZDb7MLX/RMy9xaEo30vIdLRkSg6ZPlzdz/oo
w/gDsHYDT79LwFKiRDWnFKn9GfZ4YKkbFa0AZJVm41wVWKHb/jmixUUuUtSOvEI5egbdsXjYtyXj
dP2QuXn8698LwYwdpiW5A2ikLE23TLiQTkvesBbxY6rwu7oo5aaGNM710eut5be4wmi9yZL1zqQj
0N4KDIOjjpyx1+fbCRlBANk30BMSFX1TrUGjweLP/l/Caj+9LXu+SkOYZAC8dgOI4v66ki3jNMmI
aYRC8AzJNckfhyW+9d0VVbkkVbvQSUXmfX2wkoRtr2v4EUsw5v590qb/M4zNrzBXAmyKGMKjKKjG
bqFaPMnvS3ed1q+h9g+yfSXUT3nUt4DjXlt25FV/8dJzufVmv8dXvuUEwDsYjc3yprDkeBJXOn1r
DywPugcaRAX74JUBdMH5d+lKTaF8K6hqDECWMo4Fe6tfYP7UUDwa+kxJPg51tNYSvosz7zcsFAIh
EGrnVz3oSrSRuWtUMFrBtwtARtXQDTeUs5HmDWhVAWenVvUURt7iSXBt9slGsVN+iL45WjEH9Jqo
J41uIGIkAz01Q99udvXBokyrFsSWS/0PBRpLoxH2EG1f16wHwe8S03LNPCI4qvSMo9OgNv+T+rDA
CbB6bJuG255CE/At8tDO15crD0LSGBR6EfUC3t8PLBUHQnZbotvcrDcUPUY8WuOiKF1sikx9xovS
BePgEfQ3lBrFQHyS+6ZW9B2z2FJel88GilZgE9I+JgtfKH/j4U+2Q3HvzgPibKPucAgUbeyzYOQh
IGqBaaPP4ZaUsYnigzU17UjBePaFhhApsIeRUkM75xiEgXDsznpZsbWXaIC0wo1rjIN16WHyPFmK
r94d2jyRMaDMijbDrleakFPGjdwpwvRXgvvdc3quLiFhqTYiyTkwRu4E9X11eg97KRinrLSeSVzX
9CiY2ISaZwrhW2wLh07kQZ0QA6ScultI5FPqm/I9QPBRGupRX5QTe5A7ns5iUZ+a/VwMTOw0IuzP
MGDr9VutMWZffSe0/COdSLOPOOgUfAMRg3c8QkUOepGCmCm1q2pFCLDppv+bx3RgZQGHn6c8ytiL
z3gcPGXjYdm1lMoe/RdGnOt320nLUpN41bCAswy9pp9VvYcMHXtRNnhPVI32xtgXC00DhgjfBTe2
YT7GII4iqzuHQcMQCGz27wQlvYp+K2mG12p3jil50ElGNxo1MLf3/GwiZuk52l3zHWTA1WN+3d89
3Qi232mhgEz0rRcxqfqoCXEG0Itbr1PLDfdLGWN2NhaZdhArBn2Ngz3TLW+v3k5F3uLHV2N4b/rf
LIrEX4gn+f+BbplFXtLQwPl/83PJtcrFYK6K9odBXuPo9skldUHe2y+e/UPorSn3OVPdzXBvFywV
E35UYodMGZVfYc/G5O7ibtTNhaiDSPw+2MRYHc/trXUtf7GY7M87xz1v7+GfusN0cQ5YDbIYvErk
BaATTpUPe/j3P7dv2xlRMgSPQV1IIdjKTT6P0pG67lD7TQNbeoHXIAptYphHwwnxlD7zA8Uls+q1
3N71NxRaAQG4rayWJy8mQtqrkgO5TyrdpBOjzAsUIqLMfvL//+7kS8pbX0ncxLowf1KBkGzhFXGn
C+il11pGOKvwI1xCayvZwAUA+znwDAUjUuEoRVDRMfN1SrQGtkbVa6MgGt22viHGh+kWDwBARKyp
9G4XzK17T1IS/9yTCw0K6e5ge1cwgAuvY3MAuZJTag7oBzgXj5nhtRq4+5cZsS50nY730wnqMorQ
r9tQjPawEg4RciBwv9un1WfE6NKUcbfc+X6VrOiO8zg6khRI+kQHcDlxgeGr0ldkTQ9A1z4vZcfK
fnyx6rqVBE0mUc7NwQ53om7+mW2NnyvB6ANntVVvm2ZxL9rVBbzQNALtyGBnvJCrIMdKpOVJ1UIG
7dAgzJjfim1iatYXowq2PDncj3kcN02eewAhe9+Ol/sxfozlysxWzZMpkl3ZeZ0QoUMoeiSUuIAx
glrOERi3Roh+grVUDGFMSSmmWLa8RHjMSBuYau5GeIAIWoZJUe5Im42WBoWRcQLiwog5zrbveWKt
Qr25Z1yYU4PgsDbJ4o2p6c40k6/grVchb4jbk+dLCpIHwxzFp04shxYMSb1QnsEkdz32uWCyTznN
9/tKTj0rgHmyQ1P0YMpVzbQNr6Mty1Hzrf5ddVmqNGOrpHwQs15igij0tyVIPU1vXvnKwWkFszvr
ANJ8oDyZpUwuQV5sXo1Ll3j6fevSdPVaBh0aMl6AkL7Rc3Zx/chM9iGf//gxpaBTdbisSCvrF9HC
r/swJk742mMg9E/QMRrRomIfDcfpwGWadL71Xj1HWILwiNN3q0sMV0mr6iHSnEC7NJijntxNiSU5
LZaTCrK3Ad2Y+NwdMRVRCX58QL+Gr1JgjmI8GHzXAhivqlirFLYxZyuxhFjaXrJDNYXdBiLhwG/n
w3Z6SwszzxWT9cVfQ9GlxQm2scM85d2LJSm6FvVIa8MVkRJb8c6EAJNtC+tfYfHAOon0d7caJCn+
LYhAZPARSw9KdF6kpNC5UASP2860VnG/lR7W64/3I5hcxgd1Hvs3AC+bu5ow/wbbN/GR1xN23W1H
cOHqGIh4l4oaN2hqhsf/tOyLqSguW71ow5eO+70Smo4NKK4olh8nvonCTfVC5kg5W6jLHKzq8Plw
zdIMqnnGK04Sf5Y8O+YW5ykVjpcIdI7crIeQUZ44zu4siH5m8X//WiN9E3r8+8sOjcddXHfsHKcG
T8xnDho/0UO8GtYjtJjLHbfHnqSvyHzGPKnSw5jytK2l9oCNNLzExs8qqsU63Ol0ZXKznldfRPOi
+2Ik73A0a87nq6CLAjuz0cZ1nEAj7NHAYdLCFUI7JrgtMoD/ceHaKMjWFgqfqg4hnYjh+vG0ihni
Tb7YM3HmbWdRz0iXZZJ0FwhaiJ8lGuYxExYRVtYdDcXLRR445qOUgP65KUUGcRMiTq0SxMxwpW4l
hZvEnBkjWlAb18LNkdphxyl6wQ+9I9w5FvGgLPS/8+Tx4fBz7bQbYFEocF6J2BrTcYmebzKgJAap
tiLCY7TZdqGogxJPRM69KeJkR6vQFRTOoqIjZFqWFCmej5Eg/cfslsSisZy4+5vLzpyDa486CQs5
PcTTkCydnp6VaUXpjkMhotX3pzJ6skguxDCZFRk8NW2o9khnp3vtgpSg/wIvs3ut8u82OwjSqmku
MUgrFalEk/U09WVxl+/Ax+dDnq9QNurTQQ2Iosc5Cc5mmdWz4IR/LObxQ5PzPcCjEBZnbiWZrbRp
zahlSgXdG0uu1Hxmcd9Wkxz95I73XVe5aRVtPXiRw6Oww6BQ1teGI8FNqEfAk7IYlYYm34a1Q6e4
0EG9H2VFt1/4mWrCeAsAInWZA6ONY+W714fax5RXIvJt7jzcxzMAhrP7tc+kiWqehab+UNgvrD/3
KjQg6uqVaSiFd1+YdmjJyPco9TaDS9HLXpczZz5wqQwJ37eqdSF5KwL5cIFvPMsyre8A1HeeZKvH
J5+nH4O8tuD09vRkQ3ZQMFbTXkfby3J/gRANfGUnpFjwcXwEQo06a00faEIqr3IS/FUgP4w5QcEJ
Yt3iL3HXizeJ93iijlonRx22D0JTSGJK9EFSo0du3N/ok4emfFejbp4JBfENQoxAa1NEJZDhIqgd
COH9a41T/EMojTcwRrMEqzsNQEQOtkgfBfIvn47S/xyeMAPMYDOczOnold+jy8c2fR79ByoaG4vO
qrI6LB0Dy3x0+bRgr3/buYOIksRC0ZM79ZZvUAFmMqTbtCNg8lEF3XBs78UkZWhYce35XefspJYx
Rs+CBtnR1UYR+FqPDsAa5LbSuXQR2Vw0E8UYLeFEIWflHnCEoqxfy5VpdFanq6Pg2yF2r0qUb7By
8Tpe3ILHE0MGPJKCBah43Gte/ge707BxiIqo1WJxvSyhaE8PoVin6QCP6GZFEv8ubByzzzGQT+jz
3hoBTYOwL7eWuFdBgidmjkix86XO7Yu+v1XMylIrOI4xUSHSZqpAYhVU7jSY/3Sh4UwcNA1kxJP3
iUeFaoBLuSgIqRT7E1hyVDa/xviaAcvXNKmpuPdCQPHAyE6BDkPWNr2OfEATMPIe3L7rUA4oK6Up
hTRVQTm4csjfIezasVHTczKCNLMIigd69rOF87Js8QZCA7iMZ75XyEitgvmnjdohUx45kBIZ1HMg
nftC17rsivOopsuyjPdNZgk74M3gnJ0j2n9Oj9BSJj+zgsIxFKSjrYoBKnr6Uyi4ZbMI1PU66LNT
FA7EeBRYOkHmKtU9pCs1qD0odQyoXOx+dbrdu0Gw0lTWuy62GgviJqgaNHnzDsd0oMCb/Q3exChn
peUi1LtfcXeGnpafBZayvod5D+3jY7Ak2WMI6xtRjYwZaxQ/fNy+PLwQPqwUk4TL6QRSfGJn+Jhb
cB4Ea0icXs8pU+EJtwci9Tce9ACUkYrW/RNQ2hyt6X0KKAPG1kwwdeZ08YUOdDt5N84mGyeBbCw4
aXGQezJm/jcLH/E34HkGQwvptgStsJNRNQ7b7npYPpgXtl+hS900ZqmCN2Eh3RgSUFs1ENvgj+D8
azEvmJfCDCXWhqblmcPIxSXkD7eK4JoaL4bL6Qoqlrz1FFUrv9GGvjkyvvYT7op3jCCoGGmi5nLu
Uuw91wNjRpfeWvs9myLspUuxECQJAhEtpPNYVjBwYJ8yIF7givk/N1V7DY6tLdQ35IXWJ1LJTYe+
gf3H7m4E8aja1BctN+zuUcRAYWBxtOq9GhaucK+x/hZpttaoPFFSi4PIvJWVEK8dbd3KbBzjHxOK
aBnG9jrbm8g4AAyVtai2/IQrwkaKJjNZqmY+JEA4eEzt295KxYtDNb9bhnbmyHgmE0CNvgtPVBrr
6zOD2Gw5l0M7SBQxMs88JJ4DiOBFM+jly7syMJtZdAy0IiJjMAJe3A8rYMzhJ81GPQot04BnsDuG
twsGlPUqimVBOdMwiASFYKmRK09Xhazev0wgKptbTrCa0M/t0dvCi8K9M1lLB7b7TtK0weHqOPEV
6w1KLYi/YkOSSNR0iWBsfdLha68ZYCJ0inGKCBuCwL13TWaynxNXXcjX+jd/Ol0Be78gqEwhvBtb
ldwO8DZXtNo6c6uvG1+4KkgpkBL9n4x/N6D3mKJeIEkgEziiokjCcZ1YDIJjWfcn7LeI/rvGxNRM
niGrKeI9DSzhmijPU1+A73dOkpbs+W52y7E40E2exSY7WpOpemiqOjGmT7TzJNoI6ZLb3hHFWctN
rMC2q97ahwkZdbPJiLd5SuJEyQj+FJazwOGGGVtEEvzVEOqjXNiunXEsI3tobb6hFgQbi4zKS1gP
XM9WipSt3sSzW4/fDE9nvIy1mqGElCh48Cx6IPmui9FGJmlSkoxEw0XdhAW+iDPUYYL+7TnB9wpI
5hhURlyRnyY9GPUWLQsQ7AjsnXfODSBm1e+TGORTbyGHP1pvp3P4xZ7pjlpvqRt+arzihPNz19jt
2srIbPUAwaDB6A+pTsNeZ6fDdwiRW6rgUFmmKpWcfWVS7WhUvWrgt4VhvgTFR7T3RK4w+05uFLPe
V0I41/2W/iWrRCIyVDvfOA9pkoscmxTmVaL+w/PigdL552b5IiZaOiM+37bbr/KVs1JihXzu7Dy4
CXInzH4HVhvN3a9uXZJNk8aln2EHLm+kDBdcrT1v0OIcZx0JDd8tqNDZ7ia1B9pI4znVkvVO8kVr
+rhzRIaKx8f9G8I9alYy/Z7E5P0phdo9byE/6YGHeDJGt/+oHHU3QeS29e2PYu3rhgAKctwbQo8I
ppQA/q17GSCmjPC+eKlRkR/CPCsAW+mOCKPwzKn3CUbT+iMTJ+DySgApiwdeQxrutQXIb2qSPDI9
Jy0u0F7+Lz20SqfccBfTEVUO/z2WrmUwolSaUE4UIhiTaa1/PWRfJHBv7ti9u9DAk2pFhVwrQI3x
Z09P7BLZo5LJksZRCQHyz5+n5HP9c9S+QlIpIIfGJUu4N+9g1GDqs0VKQXbW0Aa4fn28VCv0KTAc
BpyaV4JspY7vLp34Yro7DHp2G5QDb3ipoeBSqXh2Seurte7XavA9RYnJAiFO8fF7I/pFys6KtEef
syEr60XC8b+r5qnK5wcEzDJjhJ89yhBQQfoYmcVYhM1llOtJXDjBTZkDYTZDfKopY7sJCtWbze74
6gSOqvWU7UKg7FMlysLwu3FGsv1oAv1GxvzsB6C7fjaQs9FFCYR7JinE63prVUlmiEqb0NlOIVi6
YS5ArzagAujsP030XluEKpu4GxjsSVGtny6x8jBERUh+xoLo30qIrSSbnbB9PYhn1MrKqMswuo8P
9jHDC7nDTZI+3jP2/A8rLxWxfOhC4pPgOSKReIFfuwYzCMr1YYKXA15WEpLTHnWnsUfyhRKXDhME
iUiUlM7EAVoELi2O/IDcaofDx0YUKoPl7imW6lnOeecMw0aGCqILVlawJSGFFz5lW8UAeHqHcOuS
a8uU6O1R1lsqCAa66SyBiBfdxUWalzIH0sMQWifEVCdSwgxvfzdno3gOHz2cH646gRoxI3Dk/OLe
LNfTb61ycgrXGDcslP545n42mYoptpgNdhCWqvZEmQbSh+W5+3+2iGt7u96TdeSQajiKiUPNWok7
1QKOy5hUxF0aE4It1TM2KGXEDgc14SrpeByQK0ruoDCWCGBi9wheDbDGr/xTUYddAd20b30fF+t9
MXOF13omC+Y/XPKJh6iGEfj2DkF35FOCuMYB20AGN4F0kDoaU9w25r6Ymp25iePMU1qYxLegNl/V
GUPvwTvruhur0Ij1TH+8EzeYR1AlkMzGdOcmYwZsYYaX7uSfo3i5kmd+UNXKldT6cjd0MjGFqLmZ
UdrQG8RnECOY3YrQNveIXzHhOO2zksIV7WjmaRdsztu28aMCTSS0d9xQvZMkX86ES2bYZoWD/veA
Z5wg3r4D80bJibo5S4EQWa2mTS6xoTC9HEK3D89rmUPe0DA9sQH7Vaorsr1cmQ6Z0g/bEgtfGt5y
6McQu+EGle6lBgRvV+yZvIBLIbrLLrAJ6IGVjeKpWhwH8Lg1c6eUC1HLbQy/mQntcdaV0s+gSsJ5
pH+vvEof43NQf4slnmrbRDwQ17WsI2DSFaznJ71ISzzx9LwRd9bB9lR/4YLOvn8uHvJMs3RFbnQX
0dDr32GF2KJEMl5xSG0bYorloisSQ/n0YnkcIrZKhOD/yezvYmcrI0eIKj78zJzJ2N4vwO/f7l8+
HEo0rxkOl7QInubciIbYa6DaE1cOd/Yt9W/uH00A9GHFfCiA7Lr4d6wSJnWVh7PXhIc3WrxEcHEO
2c9AK3hbIFxh26l5wUeBJF3nQfq7bij+f6SBS29a10JsUaHrdnc3KvMQG+5CIor8ChysVo/Z18m5
SVounBAK0s5nlQbbuEf4pD5gbYgbZiKGqlO6VB+qn7JozUuLMcCJ0hLO3HCpb6a6WOmGsiQbpCY2
uc9Ol8THQzdaVHfy71iPqyvqnzyyKv4jtbIFOw6Wx5aebHRmsSnULH6Mtjterenaa04twTWEiS7a
Rqtxo6KDhaXETQq0YwQ4hGsi4Hri95M7cam/EKhoPimBAzS9vudTVVzFkwk8dhOgPfzxzBdtnatc
nqbQlY0AXy22u1F9XZk8IY2tV+e/Xzq8QYURQVcoZ7VhyuhSy3J9t8cHsLvIOcyZzn4VJuzqrvhj
zqWBnt/wBMvQtIzTnGG0nn8g/gbbRCHKe9cRM+sLCqzj8bQenNgyloS3gSpVCO9zOWqv7779auKZ
fjdYXJSkv6RIgwTqe+3NHnznHQyaGZeSeikKGqYTWaU99idMim9gBHOqTM6FFORJ9OT1tCjTFmZF
ff1Whb2++gI8+7SZ8Cld/aCDf1tZ5HZTwkQ/blxtjL5XWZz1yYTwvbN0Bfdnp/oE3vwLTdBtFVjN
+0lsay165qAq96LUes3O99HKbXRDxms1Z9QIsAsju6EnAxONeNRnvdPiWWsyovedeXmQFZvuqxKz
9gcJa7SPV3DMDuAA9O6aURbFKh7uchBbTQrfN6pvecHYDltahoaMYleYNmTT0N/1p+HGNMQ0tHsj
IOurDpqQcUCMqvt2zM23ml+8AXynkXah6y76JNmtfRcLY5r2YaZfnICWhNuQMybHrr8oDl7lmfUk
YEsBWxnm83fKMMPerE1a+HJDYKLX1zSp6oL+AGQ41zBYcwYzZHm4lN2H9s1gsjgiFsrNyf4e1Vdp
QDn1ifaFhGOo+JBCmEUUhTHwTStlO4h/uQ9ebPMeValm1mKXMrGOLI6oBD0sUOtRZo+dNWq3jgZH
S/izER+tCm/iv5nYSG16aMlSIvmnKvIOV+zpE1j4bth07W+mNeVgmAAQMouyyZQTsjFIZZr7cSxY
+R78ekdUgTdvX1avT6XsZSSAjvhMIBOjc3Bq+iYkk8bJk5zMRFxvXdTXGgZfdZppkfXrYIV5eZZM
w7kiUMSgyf+0zfsliQ8qJqJl9HycnyllfIfuDuRNx9QW/Sw3yV/vQBL25E/FGi+7mx2h5MAfZ7xM
UuvRVsUZ524Pbxbw1KQwjp04/jncxudMOvhadfsxlTDbaZsJAOIxnsBt6ejEKedfyAffehxH0N2D
FJrnfDXZT5hAbdlz3J9smsoTfddBbrds27NZE/Zr+GIHkQ4yUCr4irCbUugPG3E5uMuJs0pSmew8
u704P4JccZ/Y044b11CALIbb9979Trlg0455ziHxnWuGWkOsKXegp6ZoLzJ+Xishn5M9Qv8QqWLN
nCHwS5xF3bD0P9AQ0T9KVkT3SecBj27v8Te1OTZDLsq2OPn8EvK1WgNg3SNtQLjLchJFyBFMXIYr
WREVPoKJs0CcMBnzyHx1X9NNpfyvzEeTVdtV2Unr0tq7HSeQ9x4jSd5eVdPU0K7VSDxirLvSbB7l
SKW1GNLHHRjkqgBSOT8B+HT3bx5vdFcJT5stEHSh5FwvJVoZkxHbY+qxpqu6sqLl8L5u1hOD637M
5YXNEItrzVg/6tTNA315Pax1LQVSBoYukjlE3npJN/CImzdOWkzAI8D1A3XWMkcLO50rUWyOPx6O
mM3uSR2TswMAyyvsoXc1GQQFY1tQ5oUOCaT3Ng57bE6hxEuj3H7ASS2YznUUiR+X+2dUWizz+Z4q
K22Ndh/RTn8A6SV6+B22uIjsXdJeq5fkLCzLXgCv9qYBvuK6Qky2k6XnUEphx+ffIMBjB4o+O3XO
I6IuDBjYNNFWNqX686poJB0EPli6ys3poJN2G/AtX00khgysvDswOrwOCNBZpAmLQPqLCXl0H7ll
dg0QfrFGyyKKswKv+mq5jRJEA0V8QAsmcyQIIZNlyruN+is3AJBZgVYifLP2v2CEePhqgpU8MpEA
HSKGKafEYRj2+LnZJbTnehIEAb1r3cf68bou3mFdIHDyUVmVRV6JP3N3+r67BnN72cLFx+igohKN
Jl7iA/Oe0JziawJlICVNV9GkeSFIJDztFDVbxK+Jdj0r5WsIUI2LjCvMwEUVobqTLRIFHIRCkdtC
pL3BrL8YSFFi5KNnFZHCWizyC76UhSIyLg5FJjnKjTiP9CZs1PrTBlIDJ0Ck511suhuSjPowoCeQ
1cOfcjcfbJth1tKdmduZwLIJLWEeCqbJl8mU4+B5oyKH3ClcopdXwHGRmp4kOmvHkalgE+NjdQE6
ECoMyEfCP7pnhf1n8Q5O5ZxeP2u6KTPL2377JZLvj4UKzdQN+QXQgCZFYkQADZqiEOzNwVZSFSdk
0Xjh931c7MVpOwEnCKOd16SvSqUZDIDcHhirozNC5nhF34upT+Tttv4nzm1xIczCxfLIY2fO6mNp
czLNDEQNd4lgnzGOE/DaKW1CS9jIdsSQqvUrxkehWcHdb1CUYl2mHx7gP5bKncpGutUrJ0lSq4Ep
4fa+OEa1DigF0Mp+9ufP8i7LxK3P01qpFGJi9jeDKMNDk+A3a9rAYejFQ+e4m6fBDW0sTpmj+b0N
59OuBgSbdsKKj5YtdH9w4c+2WpRyazWs3Rui/Y6ceo2rf1Qt+Dpbxp3HodS776JUXbBqsA9gkLV4
Mn4W7S5vPqsaackZLihJgU1GzE9rnC/qKAKMZL6FxZJ5/C2IRePYfG939n82WiVTHX1oBRPybfx0
Eb6chpaHDY+PhXUSdVXU18zgqIjUm7962KO1/JYz/K5uNGp2/wsDTd/eCXJAHKmorUOq9iwabJ5d
wrzPv62tOQT8PuJFGgRXS5hk16n/Lc4OIGqX/11f7yVEMpMba3owfjviRziBKxYDIJmt7gMMMDYi
NqQK20joKtkOS6w1hSvZFjkMyFC5jntdgsMflzn3BLxJzKT8YR3hOVEupQJBgfpyi4H6dBI75eW8
xIAfMVmAupLnuXUX4bKeyAWoIgXDh2kntb4afIMOOz+0ax8Xf6TkQaJiCTxwgyNGheZUU3nk1Ned
uUxaqBWvCPJjxG5EW5ZwYrq1izSg8tXNSSbYZAC7OIGfKcN0ZHehVroXfeOuJHMjep1B7f/8xyzP
yNpOd5eQB8G5li+l9bFG+j4HfwsWK+4rV3rK86At19Fk7t3ZXWU5vhZmbQ7zW1x+d11+Vmd6pY/B
ewJHgXONNEoJ3ZWiGSbPeVVM3QPc7Ry2muAoas5wwWUnrSCqMc8JdiwaL6rQn5f42pMf93VUDLgb
7315OrLjrxhwpTqVciOPAo02ryWBMuC6lmdUyhE0F6Hkt8OyLIt70dcPMtk3cTOu3NgH1Iv59HAX
404wa46gwRIfFF2ZCEQgZ4IG2+8CdiEGdIOe0T5Nm++UB73bFQiFhoMEKz4ZzD6cM8gfX+W1xPoS
C2tUwiVGw2f+yvy13P8F50lRoBevgA9rDl5CTQpZNpM0MFwGtgtf37BOJpHXpQ+oghRE6trTNp4K
pbArHzvqQXKdpJQoy7ID+pXtWP33eEncZ3GY+s2ngv14nceZIkfu6rVMbCmceJA2qaRw79z3pK/2
BWxiok93zJqSSmLh9lWfx2++7DXwpNQR1+5P3WQeTi8h1qArI3DktK7n+DOoK6iRxjQ+db+1KDqv
YGNVh+tukfi0udPDsVUh+QyOzrcPhST0YYRfjCRkyZWIKZA+jYbUVwaEkTCdbyyaj8UqxjnR70TZ
2BGHYvmpYEQ1tudwKZfrPBfHgKXt1H31ZAOtBbaw2OaW8vR2qcPpCno1NI+i3nfhdymkfaGViagf
a98+p8/hz0LR4QKi8Wm2Q7DQjiCiGRUraNWBBuJkiEx4uMZb5yoGehike68GfGlK1syvtbmaey72
bqgIzVd0L6wExct4SD0lPn7gXBiEChEhU2aGfC9lkyzW9pwbsk2Eg4WVrTzDng3zSsJDTMn3hccj
nda9/HPG4q8W73+WXujbNJAKkKL7lgptw77zF9pKbPiVavHexndAPAKZ1Ee+1SbQA0FbLx06+YU8
28oVyTkpkDpu8zqVwoaofeJxgoi57tlULGyV09FzUveYOQ0OqACEouKo/gStV9ENS4p18OOOBNbj
I4+KqlBoKvjUtIWkFniGogk/kSN65NAoVqAfIps5epxUri+CfLMrFA3/FIzG4fAkQC/AKlDhg3F9
cqqw032clzf8HqX+ia1jyR6ufsXuuH/6/VniDWOJZtCBTmYIleJO0GAhxBOXYw8XpKxbylRu1dWt
4Qx7I9i/gGqWfPx3/PF7kN1A++22RtE3TwsmsRjtDwNJ+E7IHefGfAkWA/8jgDKyPvoeDv7WTV8e
odWCDOcOWVZ2s1BYECypaN24C/Iu+Gi1kSF2c1tliiIHTx6TK6+d+qQPyQ7IuisIDxj8PxygD9mn
+N9iIq0yQ1wmTUOhKrR697utM9ttaRsohGJzoMn02EskIzk3HeyJESJ0jDTa1Zwrdh3Pe7FxaCcE
34EiJga5RF8XB0IxLQ7AdE8OM3bg3zvdk0u2GH+gAOQQ6qXctR+Zx51giKhiRx4AZmha7dcGYcy5
vH10dEvVWo2EY65DscGMM0moA9kzXDsiqduK8SEBkRXwsy7KRCiYm/U3Y9vn3Ywey++FIBFy80CI
onheHTctqvrHXNiDlZ+WgVuAbmAc3h779P4Ng55Q2K8RilHVuaRzKYlEKhDrIJ91uokj+3Ej+Rho
sWY5X61POzb1ZYBgTQLQNO7V6h8vSnlm/6uExJAJgUmpG0LHZNxwqcXCKVoodAFzlbUTYS2/xkPt
xmAlWnwZniuZBXr5LA1/mvi5ziIGsryIBIHJv9WMKRlneTghI5f2AUUIUD+3Hd+wt1gjqbglVj9/
ADUPLTQR3Fu35G5dbuWdWHAp/FvCqVQ4CLlkcmxMyxlA6uTiF3rkMZbw+CkZLpgI5mQpM1MfuxTb
Z1IHLjUv5SeQ14Up+CCqCGXBNZgKQGOyAJRl8qEGSYrQLE3DOJliLh4/vj2euKN5VfdtUZOuF0dq
x2+5NI40fF3HonQKsP/ejUmR0IaNCnsj6D5uB6SpGqDxa2l+y2MepTWKFl7y1ApnxDPek/WFU1bc
WBfIHu78wjuO4tiU69bbBEtOt2QULAcc/mdUE0xw2KdxaTjbgMjXdOtTb9qOfyZ44diXnCkTb2j4
7xF1U43k3OudSeB25YCUV8hOk+5lPPW6ERXxTWSwP/g8MpdP5rP+WVRjsL34TG5EW0H1pAQ+E2KV
SGw/5yp0bV6VVX5l8dQ5YOl1ViRWRQ9Ux6r2J4WLb2o0RKNSWH+st0rtmRypvYUMcpF42XbdQp6C
ujq3IANvjlVcEyJbJAdsNPzlS5Oiok+12t4EONGPB/myZN6ZpqN0rYcNAXjT/VxEOmk9n/Ni/Z/G
4p6lwgj5QY34RDSqSpCbNXDYy109vO7w6hLxcQfJwdqFeX39Xe/WfkixJ81yMjHn382v+Mq4KDrV
kRq5/1vsBvt5zty8vCLFbs03t8+js0myC3sbOQSS6aMLahODrvYKKRB6JKr49OQPQUOXuI8ws4q4
fLcmvo6Del7ia/lx3mQ1h27BOdCA8aCyyI8NxRJ5dWTJONXdhAS6a5HpBDr01Nxw4nKJimFpDInM
RKZRV6fGde5vLgRb+s+9WIoNfAW8LYVV4LYBWJb9qBUlACCpU/r+XUaRMp3zG3dTh4JScUEi+yq1
Beneg/rKwaTyrOzyKjzGiLFrrg4esZnSgCffB4Etg3KYSnwWiAUabWPtYBUCbaNrtFTg3gzwd21K
zsLQ57nrDlBZybFXSuFuedpgKgFY8dKFO7AFk0xQhl9NaRhl0rZutqz3pPMm9HhaE++Y8EiQj4bx
UQPLcuT/tlCQx/LgMbcfOUeWeVRbqpwx+vTanLV0Ie7NLePMpQ5+lJg+EKEqiafgGPriiklaz/0n
/D5v6gq3ieDkzj6UYXZTBypJGAoY84MUQxFiZ/GQfvRUqU3kGeLngIbPHSofDTE77l+PokamFwtE
SaqODADCeVAMV1yX0s9XWJiNdcbnqo7ena9CkiLUIY5e7DYe05BOXUpjsrDGFt9jsWLjJJ/NywLH
GiJqtkXc3zx/QC86PBd+NRaSpGxQObEsP513uLvmvpfADeIGBI4r8axlzWXVtABDbdUFKbz88Pfd
CQ1sEVzHFZOVOVb+CDb9jRL5l6P01RZVeV3c8kA0UrPjE+eZAsst5F6I/K5FAnHz2m3xVGy4D2OD
z3Z5am+JIkRJUKQujaYhkCVnrrSHqkU0UpDmhALw5gaTG6oTCJa5nPWZhya9RW13rKeaAAk43FvV
uLR2U5zkqYx/eqlGpteRnDnjehDkt54VQJDMVp52A6/vEol2/vcbRjURme0vel3Askg0UoOJ3iqZ
fcSMXRf+kdmxZS53pJSqBmBF4+Z/E9CTgYU/Ps46wZjwlewz63aDPGo8+TN+VpEjEvgaq9Ukbc9x
9h87OvYqgP7wKX4o42IxRKHSBtKoSKwcBIss5MvzG20Fb1Rg49sKvLLPME9mJ86Gfkg17KGCJLES
RzOZEgFe1Is+jpn/Vui8FNxlaoDTU9ggfH2h5hQ5AezmGQ3mHSun74r0G4ghoqrA2rFXogxx0N3R
MVa4Yqd2LCEC5F5i9EICZb5y08PGHblXoDgL4EFwh8C1yeHz+tlvWOZARJTNS+XLFkfRp6Twr0oe
rDlgUP4qdw2SG6xzI+chGbe5e+AvJ2luDUmOPDA2J56jScDi1b1FCqkSJq774R7rQUIHqgL6YKvg
MwV+mcyD7moS5EI7ntMCrU1NkwQP+l97t6RTkey1pK7RFYCA9BvCK5paUHlBnFoWY1zp8HjZcLhj
5CA/qlpo/6gdhrGbRlz+pnKP6sT4TcHloWeij5kUjyQ9xdTWpEy9hMWGjO+JuJjM9KASbcxNW0L7
7ekgQi5XWhBK5wKw2f/WGWfXj+ZhT1n4eFajCTARyg8a6jiDLAg+gcOO8AJjV9MYjeRTMS7WiUGf
v11jfAbgOIwmFTXYXemQ3pV6E7AWPt6NauJc2O4xvEo4WU/ygkmY+pdouJpBvwjVXc2BwM+U2VLl
T8Z4dBilCRI2B7rgi82RoU1PERSYWnb+2tCrEOI0plVYxcvZtNStEM+lFQeXxxBtiwJWpmM238/f
IouUeynpnCL1QP0d+M+rQFgTZQTbRmCGIa8hA5nqGp4xvStmQwtrps4N6JBsRmnIaZgBdg+ibXta
ztshtTk/BG2wjOdZuKQfulmDEdqnJdLk2mI57bgLO2yPRifl1Tkuowmz9cA0Pczq4H/No3LHcSRU
8smFv3h3g1D2VOOYOjTD0JEeOvumyb8VP1+7tcZUlnY7EpYS39dat/aa2XNvHaiKTRgjes7Pzo9B
Y/5X0FEtmAaP9bU5RE3aHku6zHM+qeAbCxV9GS89vzdd/C/ItvoSIho6vjXpTKI73FNtPOYaZSy3
dl/AiG9d+9prIv/z4LsIoy8gDvkPbFAWdF76TPIQ4W+XlMBKgS1bSMPqwOzBnIsHBTtruxzJa+Li
1gH0twfcttZZ5pn/caSlBXAZcxVhIwGaq2tzW6jU2cjp9jDSz8S5POL0kgzbOKEEpYNcLsq7sm1i
cFlQ5+tZmtiXE8dlgm4F8lg3o68TatnZLK51eF5PvgcRIjYOW0Lz6ghkGWLaW21InMiGRzlAmDf8
dD3s6lZn6c8fwgNwQ2lFVeDgKyeCZVVeseMnDcYlEZoonlcK3O/OIivcMUEawLhPtL1XVNSqLTpk
sNdyizflNCSESue/BiUbCA/sAHd6oZQIMaSss4aviLlQX1lBOakXjmnjv2svGRX3nIiydjpxOjQU
zLKa/aashLNBe4zitWZVIyy8ontQAlFkqfqWuujXMBY2n/pU8uQE3Kz0h4MQxT4avU22PPkCzjIS
2YhCvbFU9GunSBHtxBn3fuDDMS3a3TJ78JSiY5OJ2U4gk9M3/ZSRb2rZsQ5G4I+parMik5y0r1ti
RacLriifBHwy+AEgGidNQyRntESBYB+a8oa055tlfdVmtH027mqpkIi2ejN5hvPAbe9qH2Jq73nd
852+avkKjiake+HOWAdvcJZnvOp1NiPx7JS8mL9cPfa4GiWw/eSsqyoOfq0tbZw23GZOqgxJA3GX
kEpTdJjI1yo1vEbXCYFKtehlNBRWX8lWuu30H0bhRURKKKqVmyEyiYbqqxiNukmYE81uVKrIvOkE
S9IhOG2ctyCnrpzut/9T59NIgdtkOF8eYdMLQxElyiaj8ouGPtrYNZKgVbv9WJtpxx2eXsXzK4Ul
eI2O+K7edYGkJM1jbnUV1dG4Vulha39UXUaI7Js/Ejcv1gNdquVLq7aNcoHkNGZr2m+4n61myg+b
hHnNPjuMaCYSBdp66VsoM/ISHsXQM0CAI+ps/h194/gMvKaX45i8/jKpHx9nAuoKtiJ8PqDSJ6I5
KIZON0Cq0P+6A9QqDexq5Nh5raAaNvpG/VPXkiIlXCuJEEUIY3fLdpZ4l1SANJRacDI8/rRh6k4l
PxCxZx1gix26ZDgTavgA1YUDvXh8MS3Y8F2giL3ZaquymrexWZeyizVoWT3k3g/YqW/sIu+i8lzl
RVTBLKUKabR6eCDCav4yYap/5HNMOptBitZ0UqfmWVTXZ71TS/9F9C3HGanlRIt864BxbVEeUwiR
LKW1o5gAMZ9ztM4IUOy1h2gaJxzxoJxuXBnqbELl0wk8rX+Xsn9t/qni4l4VwZtdJ2ilfeU8Rxx8
rEa86zohxPLLKWcILU2KGITlEeMi0RYUDJsr0MiNAnC1hVd8krNfNUM3vkEIBwbx9jGMvWT/841f
G2wc0T2PPXI1t7omrupLab0xqPjFTZv/LiPfW/LffkSpRf3dbbeBMQMboqakIzsM76Vx9Mx6L8pk
lRVqVjpI1FGjaKGZ11x42DU6nLlfHBZSTQsAV3EMDMYeDMcCLpamlQmfX9Ba4OjD7wXTLGad/qvm
RN4IyO7ZRGDpi1d1VXuL2XlQ+AEwUJCsbHBIpU7UTENFIbaQm4W6tRgtYJziCfygVTQ8EN5o4vIv
jnUKD/4BgHSqSP4bE1i+0bSGSfyAohqsBXu+vrBPpCuSg1byb3XqOZDw5LhnZEZkUbbXB16AOZX4
SPOlOVNlvhd3rOKu5cIAsC2vzgyP+XhTFkZyDy4y09x0saUF7/1LrMXvz3uz5EVgdFMGKIK3VVvg
PD4ZAS19CaX3eBWNbXLMeptW8CCSOPOHwz3vAJ9s1A7aUNzu9VJCqz55cTIdXajUGNVMKk6LMpXw
5wjbxBnc/SCkiCFWbkBDG83Z7/G7hj3dLbg1IEAgCoQ41Ic7iEnynClIoNABcuYpJRMpYjTGlTDz
vwtpCUiM3tSug3A77j1CyhjsJU9SGglzYvje184axM2Jm/PSFKKf4iGUHoHKyYbs5gnc3jbnjsF0
ffAvBr8q0h4bzx1QkB3F/FLaSzmClc4gSv0l7yyIM4vTXh9Jtn7FkZlVj74lj7woELiNcVTvQ6qs
Z6k5CNV+4hiUsn8VmThOXB274uTv0YwzNIktQOm+7rn1GYuPtGHj4eI+NHmMzOO+7ivNmWstl3lw
CiNsiMt8UAzkoV6KkZ6tpJ39UihsSVrxhZx8oEuQ1SnjxCBryZvmkEJeExmGVbOmydjGBTdu8IEP
GPa5PUR+XdkKXmtEMy0xuKnM474d65acMisYc1ZHr0tNqqRWzYgNSnETyGY5T/GYAMF4L/Myquqj
aGiFOw9kjMVZgPhkWp6S/erYRN2zOpMeDsBHRCGslN/+qDlq+YSTINFVizS2D+tj3aMhmyQqDo3j
WhHmNrbH5ssAmAbYUbApMdqklwqifGPLJIE48T9UaqUipreXlfQ3cZn0pQr3n63UOoRrV8F/7Aw6
8G7awP5HtJB5NgnAj05ODAJkNOBH3vD1kzczV3lHWZ+85iV5izi+tFndTI12UULk9FGqSr4zGbt5
PJGFpL80c0fTPdSHFiRSaGLi9734nav6n4CCfKo7CrCNlzheMm01EcmHl3chK0S70fl1x+udXzd+
ZGQtVKUZkMMj5JJgw4vxVNlmKUUcGJiSX+/KOQG6W/fqn0PJ0gGZYBjzpQ4R6p0NUD2V+Ffe4LMI
mwGjZP/dvH1ggVGWzYDk6IB6mKpBO1s35qmRVehYLehO0NEQk5TG3l1QCXv/YWjIOAPe6mkUaHqA
UXdTO+OvE5yVhY1LyM2hY6LjJw72nGpXPRSfgDIhe/ZraY7Zz5qnebIG0iwp5uRLNd4vYRl6pJ5W
C5m/6pmZHGIXFQB3JeYDsEj4T0Lr2ucJz+WeluSmonaDBHEUUha2H39qFY2ucjO5X7rbrAo+rXn7
T9XwxYjLkAnyt/xMPI8F+0RWEg3xW/kbWvfdYUM5iHLxqaV2ImfKyNuuTa2un6sdjsFvrc95CcY2
30TMJIUnPDzGoiVWgakT2Vd3D8MSWx8SrbkhXgjt+3ZJ/UolIEaIdZNz4LdpAgYIZTCowPOKP6ng
W0wq2x1Ii8IcMEcWnH7oDtcsOsPWL9Uv1/PwS8aeG8f8ThEz2rNCoYeX4USVRitbOSlYXddIFonN
kkrh+ckom9sXLxCxmVswua4v7ITYyYMsKxM29Kvb/EcvElcK+ewsV8o6z5BwggbCEkLAzaBJoe6w
dZoRUm70QOVtVYiKbN2pXBwydW8jHyPJd7OhZWPpUAnY0xArlNogNYxZDVNKXjZSuycTqLyQ62m8
km0O5GKIAUIUg88+2CmEL9SAW79lkxqOXlpqKpPGG48OmI2P6dZLSaPv6CbuuJcJcsuKE8+h9OWH
egsOqvAqUKT+gJTtvA96J/zeR3lyOtuLaKcQnkcZh1b84tjxBV6MHKbP7DkqwS94EP15GaC8tEGQ
vzy70uEtzyOBttgW4n6fVV4qQBn+Ds5VLyMgyy1DFKHMbeRWI4pHLW98ybqJGLzrPQ5PUT4WgpOJ
LmbT23htpX6AEvleCTkZ/enmvDKmO30lnl+Xf6vAGTc0iZO829IIM0wlCIKUmyS57pRRO8JxPHuu
k5UugRbHeByYEXe6mf9dNzKwrct1TANh7KI4wsn5B03EggWa0wFqaO1nxEFkeT656hNIDSv9ddt0
ugyRbfBwGovQCxLIDAu16D6bwaGE3c7FY/v3St/QA8Wt1on8Vkyc5NmawskkU1qltboRDYmt7Pz2
/P4h3rV2OkdDpLR6gf1UJOztGC4w20KxtyJDsArWMxE9fgU+vAzo6pEsqNAxgx/DyPnMKiD2c1Q8
1wfYyrend8Wa+VL32v7KvfyWCENGZAkZO0+d/zaJUYdUuyhsRT5S+gBmyKgaoyqAvCot44H5po+K
Zfc0c1KlEF9Ad3cmnTKWp1cOImc3qTH2fxSNAduCI7T++Xjy2sJiInu7bHdxSB4KxE3EiX/Crp3A
ox3lJazdZgpzwl0EbK7rG7jaBUPStofXxl82xSn05jhra3wBRog0V0yvl357PGPCbAJBpnFzp+W4
kXFYYVuvV5H01i7Lfljz0nHwxEASmT/2zUk7FWwR5ovGqEZtE2a7UiQiOYYagIzYSkoTv0eh8wEe
+OxBEgfr1zJJ8m4q952Z/qhY1q0KmuUxTfV+rWd+Vvre7CvvCJg4YHdyjqt5mBpo+t6XMso8be3+
dGI6rYPRYjtcQvaEOV2hekjBCr0Ob2Ds7+CA+r26cu8sM8wahp/0EpTLZTZbmiBBUjpjkGZT83Ka
6oacoZZXEa7SADxpQ6thOh5JTdwpY5BspZm4GixOtd5KVLSOHnV7Btk+aN4ICCwLUupNPOypL7PF
S1XzOaii0WM5FdE+is4a3AmiiwZHnkmNqhE2CazeFNiVaaLqXDy0FbMqbjx0YfWJ4rOR6BLBNPaK
rCqb1btiS/bR0RdHxDe+iLhUxQsLn7xfJSd8k9+GNvSD2yb8NnDDHajL/HZuzk7wl0wQvONxfewK
4x7yuuI8g8Z8vsnkrsoPg00eDJ0aypBtCR9vB5reZKXojLaiT8/BC013Wc6cqPN+KUfa81Iqm4Tw
X+u8nmY+tAnaembImY7mfrAHU0efXxOP8BgF+nFT8xIUFEZFS1nG04d07AhhsFsHTtOL+J9IoJDj
qxQPTeuPIK21BjXab/hvGOJX5KrevnwaVst3J9cKub6NHeAjXXT/BhJfGtl0dsp422/RCYZanK6B
sNQxwepug0slqrTJNz949VEhyzPTxYyoXuf9opOQt3VGjQzSO+Xi7apfGZfdEfgW130/FCzntnwx
nC6MfkXy7AvtrupZyKxC2gXHO2P1yYvLDdfKcKcv6BR+tSDj6dZ+vpEst4a7LaaV+c4l9ABDmVlX
hYaIN60eSnWHsj4TXFCQki3TqjubOkibupl4iCr/3IO91eouzOGq3vquHNMttP18xEHdGo85qFC4
+JHY1RPT8o7DvjcJtGC8Gt95gKQpcP5vBnOzZqG0J8eASm4qtD+NLDioX2gILHVzQvJNXunfq72z
2GtUdG7NRsiZikbntYOeD19mJqAlgHODaMK5GfDHwNV+FR852GRikIpTD8GL32LnPJ8NCowgKVfM
yDAErs0k+Is6JQU5AFPRInRgJ+NECGBLaH92oyP1OiXuHdwbPjSVOKnZX7rjIKGNseeGG9BTXGc2
6z/wqHLrpDFbM54vsJPDHDz/zNt3EUKx1YJ35S/Q6WB1VnDy9oT4+M9MmtPJ0xDzpgMtt/VJopxZ
x0oKchgSE/hWL/7XaeP7O9bej/OFpUr27R7IY9xjAe7OtdNW1YStLwz6+/xx7GmtufkTyyUUXyhr
fsZ7FireNUu8s1VZUjQfVJbh7kSsJiMuo82ivtoFQAS3IVvNMUG6uTdYuBs6ohWjaj9kuSbuLDsm
dA1e7UZnq5E/JNuCgXKEHXqnrrTSW3ZaBYFGdh5AhDlk6tplmIs+R3GiSKLeH/6OnZ+SRaCwzyCU
/Ps3RbO62mc2Os8vAEX4XXojAjdKIkqINFwsNVX/9H3qPriRpm9ESkKW/DbLpuXVUfu6SMuq6mRa
HJExSbjfy2bxRQPtcp/LbwWSMjVYYH4RYomPFjwZB3RcsF9e9gzgJC7jV69ALO6xcpZzx3Xpt4Cg
83pyGNrbJTclw4tM/D3cFW67ujJnV92hscH7R/sd9AQe3qVBHUxzKuKpw8xQO3a80rHYpR5U9tj6
50UP26HYQCfl6R03xdHc1iPtXSfnWXyMFn3X6qVnBgqlfOB4TlujusjmOqxqCRIhu5cu126JNjGk
c1sWPJq8urwjpePgtPncPgPeLNUkEWeDgsVgpjsx/Tr49awoTqDPjQ3eEANwgCJjFqH0gHWYFHU4
x7PTpD/mBokc4bgd8uEBEmA0sGJNusHPpA0V6bfdGiZ4tGWvH1fzzZG5HaTXYfszVFMB3asFoeYD
oaQQFfKaOALiUjvsWFkTbSmXBxjPqY+hi7rknwRTMTnsV4wdkfbZquv4aN8PxrwbCECpsDx3TtHv
ya3QDNjVG1ogTqXogOn/EwWM+0xIU+aMKZeqJaGuuZp1C7mOAW7nnxrbaYx9uccbKGZNIMookvkS
TblwSam2LO7C4oFjqsXsf2vjp+fVxYkLXtv4L2MYiujLEpdfpJqEz+t/V4hrnoDjB0TtbmnGg73U
VRW29NBTIm2l3hEDgyAFNamZOW2pDuZMNSkkZ1p1H4QfCLdtPuTMCe0LqqUcNirCe+0s19SbpQlM
2hUieU7jKJDCwiHRYn0CKBNgheV0a/IVI0T+kI+BJSQflN2gQg2Ar0NAL0oZ/F9a5zI9YLMZvEMV
t+FiPwyScA8SyUwdO0NP9y3HjWXrpOmTv8HbTSgNlDP1NQEiOX5gERmVsEn2BXBC8aNI0f2wqa1d
rVeQZ3Wk5R0sBBCeUOaoNir3Hf0uTr206g7MW+L+leBu/lYg4nHMoAdO6g4JakLHWZRzDhQXpY2T
PhkX443aggS0/sgsh18NsujLRwVqClDAk3wYUGdW2JjWqEYnUF2lWGdI8ulOnIi2XDYhAIBLH7Rx
w8F5LCej8S7v9ijjalHQK+9KitJVLmFTN8aPkA/6LMRVAI5JL8T+TM5vkmh9phBqnXPsD+VRnO2Q
Z8v3W+Slp5czBbpZPvE0wOImSdmWzJZf0bw1vwgGoMGP2uqSFFhkEuO5r2i3QMj6X2lXooSSRYsM
9g+iyVfUbPcPBBXQyYLBgU8MfeTr/TIyzSqq6bqo6ITXo/ZOodoGK7+SB1+xq7bFqYsqiWHRx1BY
87uYBMmhLxyNboU+93w3JuI76i0/hgB8EqMcg5Rk88AKXe8Bkra3MbkP5BLNe8OkhSCy2MRq8lFG
ygsdAfPIZTlI1MmGWWxXu/nSzuU2GmK+7zS3UWXMuvQnScOw7Vc7viPQUeMZUobXESzk0hqpjmuV
EjaVzx84M+WjFmhd2SaZFxuBqYkE/nbUoC94qYxOK1bvR/OcdzEE0cbH6rYEW/76Z22/rq83DmR2
e1AH+j1+fTsKg/xBHb+U5Zo4DGNFuVEBfo8bZ1/u3AkOlqGZOf6NrnyAx4klAFiDL5cIQXEiAZyB
V7LGvPc9XmjvVgpjsSppk700EC1pT6m14oNSSsxX3cKmQJfD4dwR3aE13DWpsDtKoWNkLdDEaF+L
kRZKowpn9PFqXhBDsNT9I9f5zrNpsO44HEKxuxSxb31TZK5oSNkzYGrl0iGN9K7DIVVrC5Jag2NC
J7dWPEgNg4qn8xl1WYjROTXVvjKFoMCk9e+W/JA8RiVq5vqaMjU4Kl8lcxHZhzxJ7gPMm/cFDSb5
GafxCmNeYqwGC0IXl29F21CDa0E/YgztSB4MGe1kO0Sr1aM6LzXztW5dIW48d81Uvarbk6W2Oud7
DdeIBpc1Gu8YdJRQ3y5R/xLtvrdjFRlJZKSRbZNYY36+8YJOnCZW2GNcnBStVke4miLAPQ+yMJh8
vi7yalPRcFMVuIes0SJ375j8fqAqgYhwQRm7PnuJJoAoyOrPWow+2/G/ILlR2/xLQ5trl9C/j7L0
LKRa8je3fjW+YhAh2NvTqXg8DfLgHdIJJXxT3kUMrFgDPB49xpgPaqAMiWQk/mWkvYjWe91pYqhA
34lb5CR+xZOkAZfgKvYXEpJ/Wz7utkZMNxaeWF4qzSnfitVfdsmFgudUQ93TnvYf7OEMXY2iaB44
UF9h+va8hjYjsepx3qMO5AAb/CRamsDvKd5LJOZt+nJ9yV8E/vp2hTS4nhXT2njhWNARzHgJhTgc
mL5jpOnaqZBsHMap3Re0sQq7WU1lDelM6NdfTj3lvsOKVHNB47fGyUO2U7zll6KWUDt9JAJashh1
nnqyicMDD3neBFa5DR/kg+Bzo4nzKWVU5pvm8j91JnXkTDiKijXw8quFYzmVCPJjnaQfcj+8wjA2
fuuw8RiI04eR+nFjgveyNBGUXP5+tHwx3hNeQ/Vm2sEICf5FPl8Cy3Zj83+XfsBECDyXK4N7XWTr
/4i1uc3oimYGGLr4/azbTwwpPtULA2Lz/lOtJJS6KHRlmFW9ghtjT85cHZ2wLMrwtRtdoMqBWFuD
rf3QWrwgCcOlaQdU7vPLb0KnKqii68lN2ZtD0cVD/Yd5BsKSPpt+IvVwDRLggXBaKAILvq9Zpm4E
oWCFIy9iKi3okNKgTkotaEoqbIixQ7a7xPCPqRacMhJcsiqhA52ASFxpwLAwtyrgpCHLwxEQKT6v
5MuRTfl/xBeT9nhzl4EIA8N/plZaKIKPv2ymgPYq1cAMoyqKm9ZtQPGk1Bqa47Gn8qDKRZfJhtcC
g9i4qQhZQc3nHlTbusqVColrz94LuqSNkh+zaplMJBk+pjx2QThFI9S/u62Z3klb2eKUJowoaIig
j3txQSeQs3ucjsFGLSgo4h4AkL069QRtncD33R7tyCRaTfLb55vkBjM+UopnMP6xRaERnqKxivbH
+GP1Xq0FTVs6tzKvYsC21pDSx8rcJODJjJgSSdwUE9JgoEiyL0Ra6u3bxf6XNIPZGn6Dmh3gyTEs
W5KEzEJadX03kBSILP/erzMmUPwvSL+Jy5PwNAgO87TaF85K4KDeiFUnJyTlcFrb1oSqdv+4lYRd
m0KMqPAWhEWiNonFA4bYmnngIp7er3MRpox3uERq9t9IsVan72OrsmXUBOZDiayYXn6i2HfaprSf
mQDUQ4kdmDpvf25nNATfVPwMdilrHpxSnbQ+9UWa0upE7yZcLdxDosodfm9+6YwQ6QlhN/Susv//
Ke0rljByunh4xYCXXcWYoHXfS/OCAdXjsZzZH4oXxoPXKiSFbf5BMydGgzlf4R9dSKrYOzJrGFTw
QJsomxQYLlOrpASQxmMTlllcI19vH3YQw6YkvbwLSxwbkjXueM7rCA9ltyNak4DgFrAckONWCWJp
JsBCbMafPQCvUKAW0X0HAYDlsBOJs+2w7wKDMpkx0uGTG23wjn2CQAEze0mQHBooMZHjNCOlb5TB
ED7Pts55rwWVGNRTQNGQbT/PFOepmvEI2+dMnqb0fX07cwRM8t2Bd0omKlcF/bX+XoH7BkADFFtw
8zizuPVIh5+Py0Zgdas7e2IKiwt4l+Lv91sA3HafyVibF0gJMm5tw+7I6rgs5WlEoxfLMKg=
`pragma protect end_protected
