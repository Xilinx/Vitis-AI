`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrM41f83zxdpq7B9Bxc+63s/ThO5
lR4ebiIUudrMSnsXzTRn4negwrrB4VipTwcqyfoZbX2gIf3gPwkP3q41DFrLyf9opSDFSsyylvuq
0tfuxhMWxI0KvORiuv+DLG15sEi9Zilc4jLqmJBgxaj93813ixDm3VBlIU1BQYAYzQ6XobruGhlp
W7l+H9tAQt0BvNuSDNd6KHRHtkpbBcXPwpTyZJ7RstTWqPbVIiCntrKr2mKrXFSxquvkPLZLq2tJ
HYVxQJnJNff0Cj4DAXbuyauAwQkbGOtfpacCEHBbOoKn71l3DGej87VAqg/NuQTT+sR1Jc9eTKIy
hIMI73mJ4apVRPmItB/MkbCe4DjFMV7lM+AnFD8msIE36fX3yOCJbyPo0m9ABJ4Xz3aXuKp2vrqN
5yxlvKiuDErgESPCYDCW2rwSd7gq5D4Uc12LTb5t1jaDSWW++C0cRq1y+e/HcFaSrGHBU7TxG56K
nZjondC9Xeg1I3hTyA4Iuka1lzZhebVat8G1Gt4Tb6qCHSNcWUiQBbXnnA9GqZ40eAvuRBrMTvvG
xUJz59T4iSVh/WPNOzJQD5VQyXYNz5Un+sRoXQO/pF3fojkG5bbO7BCMXxtIh3OAMAzbxxrNqF6j
RzDCoc4XQWPRbscR4TAKtdA5Imy6M++pnanUipeX+z5kG35GtDX8x9X57Zr4HDdIGw7h7L+S4mUz
r3hPK9hLn/8kbZhP60AkvHiIzrx4JjatwU877jbKl0V4UVNpV+cHaeXb/4uUPFfBDan2kLucyCam
86xXzx6W4foKOPUMnperMrsjR10LE6XLWLoDxBtO4CLTeHPK6nE4Mnd0KKY/s4biaPDGMejJVBgj
Nc/8/7ps+af1BUSqYnPze2Y5DqJSfvCFmv9nsT2s7BZl+5IwXZI+AcTJ4o19CIBjjwuNFto5n9/C
D0sZ5Lfc6E6xTZNY38iYP03bHgROvyPYoTWqa1TQikCAd82uaqxHiTns4VuXp7dNq/+QhPvixF7P
sQxpdMrhuJnWb6f2Hu2/Y1aJa1GrGoxjYEpi8c6EzaKA+eYmuDPGRPe207unfZ+DxMt+1l98zdaL
2PfKlU0dz4eQDi+D3XDyfVh4b0/7akHB1tQK2Wp1PRd6acAwhLtnxOcCRcBD7QRYE4vwLufMwpXN
b/G52C5MjaeDqkLAh6tMmytPnBrLXrDqwL2rqgFRIfGeOte1ggu6GWLBdw6IQkRjuajOJB+b4+Ou
1dl8kGUu2HsZkzJvSJSx84l1MJP+1DP/ktkTOqGGtiuu5rRTcka+IQcFaV5oF5yy9+WeJRDx6b8z
Bh81M+fqCHGbKLrulXtiGHnbDMgdPcFhmEBBFsn8C1j63EiP9GPpqQch/RP4YmhM/lVfnkT1zB9h
6hUdoS/ZXezNMr+XSYnnG1uLwGyD6uzy47fJ28wGWBBEuxfoe7NEXlFDCVaE+SX4oJ/fGj2X9py8
XaU4mSZY2SYjwdPIsQqXrpDjTi4wvURKOPEWt/qDwvb/kz4SYs8+dzwLCjx4smdti5wPzlHgtZIw
+U8LAZCCCYrIvz1AOwwr3RVczrMzuc2uiMF1Jq0nxbYqYkN2qYSQCUz8iBhoejOIWg1n7rlIP3Vb
hquU55AJtnTCpZYcj4iOz8+4ziR3zja62tL7k1F38MMkSHrvLmOxciFgTJQ0WibqtLQqr+Vd6FjT
9mStmVIRWubyS3h9aAtSL3CEgVrm7H+uSFXu11tvhF1t39oJ4l5I4M8r0SVJOob8c2vxlaV1gmPk
BTTwb5HKNjjfqOhbyLwMiIB5m8S4XEjwQAh1oWyHiRvIlaIaTMKVrCVduhbbiMXlXeRZaNRHNpVi
ycZgTuTvQthws2Z+10WwMt+MbHojU69fVNREBPfeRrIte1Hm40lqjya1TNZLZyhBibIR1ATgW/hy
oaE9eO8PeN0cjR5bbSRdCQH2F0lPFr5nCvgiYKUMheKuXOhXfTDCP/cCr1t7JrhELX4NjXusF40l
2pP/5zuH431qm/TtBJJ5Nc0u+l9bNDDmPzbzvzcjMLZ2BWYYI6YiAjGuYC/pcif2bOcff00lFk39
GLk3Ji04p716VHzUiQA60zeV2nNG70xNeybX5hivlxbupn/08B3/ojTPHopaWNvyKvc/Jo6RGhPh
kRXTDJz5611J47jm/Vqxu9ckgINP9vOG0uCbOZtfSmBIP4qyVKBL6fQt6oou2Fuepm+/NMrsfDjt
n+CRG/IUyIAoXtCGWrwRl45hDrqiHj2Nigg5FmqxGDVzRTil2cXT5XxZmH9KUhHRKv9EI3ALcsYo
710ld+47YW3/o7qSxWfjcftM4nY06kuRVc3scDwbV5PMA/W7C6kRBRbppn44Wr4AxU1tfZzULEji
IZ10UEVEGRyLW6Dms4mhFKAThpxS891aTh2fuec7TulJ3NgenmGx57XsiXCWA56BuBq52pXpkz/H
hzJtenIfgJBOKSWm8FZ7Y5xlCajFeaUJRNzWvXsb8xxSTmHw9oqGy5mcNwA06roxxRX26J4d5MN8
aHzbwz+AVfROy+NBxOMuGQ3PvLioIhfD8qmBZQBM4+v4r8UuagdCoYnyeaGgNFrpvEnYblPSUmV2
p6zlar+s5aANT9UMl5fDonJHwh9TyZCeTPycKt1TpI3vJ50vPVvGyo9/bWZVGvPS8Bs/916mxK9p
fk67fS8/G8CwRdJ2lfw+Jx38BR8C/WJPSLZOlo1EnLM/Cohp9HFsYu+QhkAUvbd0gfr0JYgXlaTJ
0LLq0/rEaUx7USyUmV1HS5fvUrFC1WNBXoA0wLWyMaph4S+u8qsqbB6pBZ+BZGDFoBM8pBoRGfwb
iVhS8Zpb0criXWfakYILdmwBEKNT0Sh8lsH2YuAV8f18LYCltAeKIqb0l+rRPRYJr+IkANFgBfEc
1d2a/0N1AEQEqhtj0IUE5n4X/DaKJlTTdkHaQ66tExU+GiA5aTdk8KFyiTALRRFaIoXfL/tl/U8A
uCrSCKm+NNIHK20nJKWQuvv5Q11ZxdWOfN60QvJZWJUNJTBa5t09/a4LdVdFL0aCRHAXPiGzce3c
IL8i4WGYpmM0wb4GRx0i0LVjDg7BQHuY4aznGigkksWhHUvdhyps1B3F0W0bfxjHSnCaj9QHG7v4
p3pdJwPbdE/HGOddSipaxi3+QoYlmZraHtTaV82nLSXEZhSZQxVN2HeuN8TtolQ3/EGa1pX+SSP4
Ovk5nGnkZsdtsSIN/vrFMjEeuQgcOii+umfYfZ5GkZ2s7G0Dmk8d7HtyC/y6T2WVEWd414c9fces
IzESRqNzqDCsSbrHyEY8d5iBt/Sn+nI+qQjigR9UpDpwSF3el6zYV9jnnvTjOQtznZzFUo6Z0gm3
XYJG4MZsbIqcHt7q9FDRl/3/7nq7UtHPF+4518QE70mKiwJP7NSrTjQiSaFoBXPwEEL4fqSsheAA
zUifVn0+bHxrMLeIrGdVpn++cheAvI+cmIESWUEojmXCRaObsJVPM9JxBZtSvBbmNE3vGJOmHJDP
uMqbWkrNEoRVXzycVU32pWzYBZoOqD05XIe/ndEjIsp0qe8adocUZeJjLmStwthVqngX6R0EB0cn
lqxkAgS+BM8Ibe4/DMnzyg4KpX/7LQ5lj2Uo5X6M/rtwVY7Vz3tb4nIrpkW8W1128lItzmsy4nRg
YEQnkGSMn4luAfMzZH6odHUxR9gqGBORJEqPzMc0jYMMqmZLximkrcAhLF407nnQ4bQ/YX1TgWl8
AhhFIdgzJ+Fp19NZNl4jUSkhJ/TtxNO8u70z3DA87HLig+UPKZ7FXxtys49K8oaoKHOZCSG5f8xB
2TvQQAuLHE1rlLEbao+SVG9GU3yfaDBYnE3Zl8sSHLJSjPOXpxMr7Td1nz+WfTNbk10SWVdXPL8x
GjhrZc8jyv5OoHdkfzkqmQag7E1NazeXvaNWwcrYmFoQ89n6PVPSsWrCt7mXwGDzILouSEZbCtFR
JzNQmAizFil0jtWocioK6NEFzjBsHj018GBawPcP8s/Ihta8ogYjZQQhf7uLmhTflEqWOO+w2p6i
NyfNtW2l8HnWE1t6cxOjsfja7RkaHo3fPb6joIjbFjYk7DVh47oaQjSrcyntpbdceQ6wIAOYr9+g
QvopWQ0gaRDF5TIuxwJEiB/fFiXY8emBC6kLfuh6f4vb6SZrlPHUWTT1IfwdaIo7VmL/AaxmYk/0
+FNzZNZh6RGo88jLbx1Kce6Kc0Lo3ZSxwdgPqCwW44a8SSZ3SFjDwdyhHze6bg+gr8+YW8Nfu7JZ
7guBjHxC59iLPYhNcbhNaDAlNILwunoDZvTDiGLQOHPuf1LByaigBdGmZIJ2STOfZTo/AZIlAoJT
CrcRz1aS2QllIdnpQBiqt2neNqH/f00TK+vVrO2yAemrPDgwgku2Nfng3EvTKuJIV9ZpL5Gxo4DD
WIT0/TeJuShGzETvBnn8Z4x8got2wMNOcYahMUx9WzmsNjxJGQpIB3B09Nh9x1nQcVhKGhclT37D
vSh6kqszHgS7XKTKznDKZfMOpMIjOmBiFtUgl4Q+IGzBoSxDK/4yNo+LOwtUktv8+sY9QQryHvJP
p7RZUH1mrq2nSe3gueGed5pgDtqtN0z0WJWvwmytC9S9Sw43eYjrvH/VTk7uaLITtNcQmbO1WtY6
VJ88fa6nJC6DOan7Fx+SH0P3nt543SU7+p9qijq/2v8rJNRB50Y4wfEMwzi5B3zxZOfW8OjpF8bQ
Hj8zYHsklGeWME4Q2jzOExDU8r9Vm68u+9GAJaNU1zvgKfjHYRgNuAvOfSco588zQvEK6ox4FDU3
oAhuCq3MEreaQY4z4JvMP3RBy5+zthn108TXkM9tI39S36o/zVcHd+o8CX9+IYBVO5rRcMDQm5UE
1U2DdNkcJZg+PwPLDqQfnrO7dbf925xcims4QohHdGQiedIxSSfaW8Q7jZlfG3tQN99YofETQGXu
gn4huOfJBr9iFkxnnIK9o+Q9fZqNT+Yt8QjzGKPHjKXQwZkiRg+4Rbx3YPVYdQicEhJVpBIu3CLe
V1ZBGVzOGreR9K1anj2OxPAjMhAiy9sn9w6wYUiwx/49i+M00Fco69UThyMxVm/ugoJuCKNUsMWH
a4tlbefT6HBUAotMSi3dG9EiSybGTCkW4QD4B0THvsF7eN+iKh8OCGZyQkCkcvAoiM8rG3OIQbh1
D6xpJBTjq467iiSmp4R3fbIJH+gE1AQ5Qve18K0pLWhVLHXDIXgHSDk34CW0Qtb72Bog2lnk3nNu
WxhlyLL0kUfbsycabQv4/GKmkXrDdwXYI/xaAxfJlSWYCvDYd18hvWThYzTaasUstuA2KIDH0+/B
eVLoNlSjH3jzwUTi5Y/Mi3gNnUTZ40JD0kUij3x7k4DRtBG2RJnLtS1iXyC0mszw2Usay7yC3PZl
V2NcggbLAFhBWZxZDaH/FPocUfZIhrMgnzMKdK947ms/Dc9v+p9D+/r7T5O2IZwXJpfAbHcyDkzf
zT/2haQiYuQ60Hw4nhJoUuxcZNdXmgfkCiQbVYIIJQ6+sSc7T08LKVDNPxCA9yf8FGhfm2t9tLB0
OI0bp1tgK7rjGsgps0f0Z0G0BUMzVVFzLVZVrlUAIe7HJbJ557JjB450yxr+dN0HsBMucyeajak1
mOCZUR01Woe/DNxzngpcM2tm/yX6L0sc51tD0khE4qIqKR5+CRAtdLeKCwgBD971u/Qz7T05PqzA
XMWRtUNfeZWW918MPbpEd6NXJExmi9POfQAAFSLOjGxh+64zf8njHOirmRpvlRZyOcTb83uZ+xsJ
ZaHUUZ6MtpRNFfVuQHA7GPcec5CxhIJMRcN/WtIRJKoIqOHDdVG9T8zeNAHl3GHKMRmmSHBZ9fVB
0KcL+QWHhZF6tL+wK/4qQXRtfmfD8shu+s3gcTbGHDHT1qmOTKDO0PrasHSiMps3a49eJFcdpUev
twSbiGnONsYwftPEQtU1hXVzp8j6TP1G/la5yb/YQ3Gu6hk6TMhP5/OJ0vxyAw3maeZRWxvvDMpc
Rayd3D/M0nyaaCXZmFQy1HEtbaKHy1MlmS3BftLX87xLDsKfW0TCjli2NlFkDjGVFmSUCu1jkM8q
Y7hAdKNoc/uT8FZcoXAFIxikpP0GYHfetuF8tu1lQE+ol4GVgbU6BhcwiR45UGvqbFyjfTm20hqC
5azQcALwOa4iQyoAr59XdyZRKEzrdLr7D9NdoCvNn7stChWs8Ssosk9MZtaY1p0cndhNTNd7xHHG
m9PfSNIsrsUItZCCmbfVQG0fncCIaX74hTz/tHRygom3R5sw0SLhIPLXZD0mhgRD1HSBCKeF4bR0
16Rx6a8rd6Xkb2Lzcu1wNsAyeAvUbH17PJA9m8paFgjeCKaDZMdIeMVDENEz96OQnPxbo1GVNzoP
Jpk9CN/cYKZKClPv/ArFArpoxecm2ld5Q3xgwvSESOC1TGqNt+d2CcdevIZmS/rlddwUDTNkX+zp
Uae5n742ONNYZ3mCzbIncymBapUfSTb3xqwmVPjE3Q6mVL5I/bn+CmiwF089a1xQU5Vr0QfT+qAe
8muBGWlkxlX2Tx2lyDSDnUSO4e0aL2JZCivAQr9DVyZLvlsSuj+LVSDojUeCagx1dgtI0haTlXKn
i/nbuPIU2L9kJghc7dDIwNPv+h6JPDC4MCdUGRyLeu46KDSsGMFhD/kWUbRmINx7tFqQDS3Y2vdU
Yen7ZD6CFIY7XCVaeybM+CIpROEfSYrScOno0P+xiZzCS0D4F1JuOftIm48Yv0C/NBoVX81J+5w/
gW62HtFfKZm5GZBPoklgMs+e6if5wzEnM7g1+uxbua40erZBXxxwEYpvBPBrLsglpmh5aNRdDHma
yDsc160WOldDBLdDO8+c8u0KVktw4yBBfT4hE7/lzcRYnyCJ9nDBzdzHk+9NpOcoMn/C0e2buZE6
goPtbXRSY/pbB2kvFImhrrOs8t+QGxdHpnyLUW1rO6n163bUlMZ3NdOUss1NfSuVOPCzuAknIwli
e4P2uBybTBwkquaNQE5VdTYaNjoG6ORzuY4HWT4lL7ioTcW6BT7LWTfeLvMEan9xLrL3PSXxkMh4
5pHwIqaqjiCQ4+4uDe1qL07K4CEoac2NkGU4oVHWvKSyc5RQAR5KmvKI5Q0i2ZeYtw7c3YyOOWNl
oRBfCiB+QJ9KFh8wkOX1rrpxgmhcT+5QfUN2VLQyVt/VeldKYCljdRD7laV+O5vrgnitCc4tT/tG
h1n1xSdnvM90gnlxY/rjxO/WERK9HZYAJVisMD/xRD2DMuJmBe+tUdZKF/m0N6h6K2R1PEJNjShU
VCjPbEmpwZ8dcEIsNlQksG44IvigpBEAjib8K5Osi+UvGeP8SpO4KdMCtVoMYggj+Q3+qROf3b/H
C7JtfYbsmVWTaYN9fmw5EF3P3ZTbA67NERgkm6rcGAu27RZ4sfawXcnEYqefmzN1MgN1JOL59tRR
f/d/k1JrUuHnT/FZCO2YI8ZI68cvTxomYp5PqowuufdNuqiQVqgABbP5S4JdOIUQ7mM7IkwLD/uF
FCIx/TNXr+DpmhZKjx49jZnk9plTd4KoEvKegeuCMOYFv8ickj/XyC+YLXPXUOjQfFEwwlEyyWO0
rZinCjOCP07TL7vK5mwwJiECFMid0BSiDTVluYXqC+fPOzK2FEcXukID/EGp9IEIJbljTEXJ6wSG
MJMY76iLKWcIEh6nFE19YpEkrUCoukqn3qFKPIoySOETrsWOutjhiMUeVCHVRtjDz+1rwpI5zuaF
O0g2d1FdvMPikn/2xtBN5Mwiq+F+D0n0fENHwucf7fJrZUrEu4XZzRwCp5Xo+lMLquPK8/a4CxTi
O027jpL0duTxj2sDpjlk/0jC/ZXTRj/POMaIPVzxpJg6OJc6h1YM2ARn96l9QvVoRWvpTzWo7Zwy
dm0zP03c94UONe5f2txJsClKMi85Z7EWNkzWRt2alLqgiQr+3cBNyz6oGVdCwhAl4DmCnbCEt2sa
JHhgWhGMNaByEwi/3M1Nklsx7M2YXGiheRuFpufBU6o7/89aqTgcnSQaSpWRLL/w54Qwkdli69wd
k6AWZ9B1RvWwCE6bLQaItNDfzudKx1uk95juP0gMmvmvrKRi6Crcf4hsK3XVhtpKMbXE9r4TsRil
MOmsF59uriC+gZZyLOv6kmDoGlvzjUBSzPVtilSh5vDcmnN7LzFH21wAqmjTRGiqra26sqqP3+99
55jeJxxwdTFqQKi5pE7BPOaihVGX2AScZUPpNPBxk16bN1c/WK3Npev3C9UzslyXL2FUMDoB1MXh
Qrlss9QPA0CuL2ModkQgWKhn+IW7QShFulDhoQ8iQBpbF/5AGucsSq9GVLWVU8L4KRKjd7sbveCl
X754W6hyvlsNY3jGLFmOoEr65WH+DzQ5/Pgm3p5cJQLyjHF0h48cltGzH2cC+uC6G7qZ/8HwMtBD
VI0PZA7TeA+YbP+HOizgVOua4/UPtaSxNgUwS0Hz7fXsrDjqGBiMt/pEG483KK+byt+F9Dwgg0Ry
mk1GTiGKof/GZ8qlBMvLH9IXk1HHMGEOK96ZwsW4Ys2RJkJWU/59wq0KRl4sYtRyxeLkzjncaAD6
sc2diOSDAulNDilxu+yvcGgppQ6ph64q+AqurvEOGZmGSumuMMkkxNXjB25ZjCUg1NZsmY86+jZl
SG+yVyHNDGVYVDXQudO7aGta6AtpmZe4YdZlE+W6i9S6nQKgT+f506lL5FEmnaMtVkpWxkATrwnc
4wbt9kmEXC7qWu3tqSAJt+PHOIlZOqA3BFQIsqpwPYzVv04qcWmZkRFO9tWdTelc3vt8XNcbHQCw
K1af5Bq+BbmmTY2tB1gv4wl2JGlcTDVNWQbCHZre7tD8lksHMjF9pC/teCC9QZhSi89/y8RH2eHa
0HdSr8qdiNHDYZRjdRxVvSGLg6Wr56cCrV7FvGCwLmecgKhDXTorp7WNcPqA4GgdNYR5mTgIRWXW
CM/zoWvdaSi9isX1vxV9zfC19vzZE2YDH+iRYvbQhSRCnC9QNKCjPN9vbYu2KDplPZmmXsb45am3
KVY2THhhU8GoixlCSPkEulLtnvuV8C3jRYiUph3MH/YAXdEeD2+21xTCrw0lSW3nZ4+J/f49KL69
HOOySVVx2D5p5hQ4qkUWdOy56uBG/OVtsDfFQsY1TznsWe3ChL+pszHS6higWKM29hagCu8AdJQg
T+idBVV5H65CbMk8WTIVEhsuy72oZjaATm4ChiJrFDpoMMSzUB/702TjHqV4Iqizml4i/0mOPCRq
1+T0xx8LtRMP2GX1gVLg8pmjN8c1+j6VP9hrF+A9ndgCSwor5VxxHdAxtJrHklLRkuTPSFS6Zwb/
t9x7aqgKrOW6un7OEQoOLRTPg76YAFA7qKKsz28MmdXz66mAGcAF6RrNAx3a3SXgnIhL38wZ6X2i
cihx2rk+Diu/h3xQhwj7cgHdKrUGQ46w9yJ3bR1Fqxyl+GveS+jOYW/d20OI0KAdk5V/sNECHb+z
1JBl+esGQ05MmJvIkwvxiUOBbclji8MjAi30gPdI4c+WXCW1YpNGxx+Q0owO/SG0ici5W6nyutoj
XnXpPo+9w+LvnXmAiW3i2cgZ95Y98XQ3tLSa9/OcKIIZLQ98mOWv2XXK98MFfchtdciAPNdpLi3m
sTZ6DBKkvxNWW573zeXvnYixP8ZsN6hhsAQzJlcwJxvrs4JIg+Xwkf5XWRd2udLc1JRuSEHpUgu2
EkBxhQt9FZtU8X0dIjwn9hwXh/mcNlU8HMfzORpjSyGg77hcSHkUlPaoPqNFz2wlHuOISQhi/gen
8QxtIVmrf9zYpZnLc++JI0RPbezmhq6glz5IJSSjd5fqdDhSbyo0otck5C8VW8oHlUuYkwMYh9Ae
YNkqXm5X0opwSLejVZ0wExU+78nUApe0+MhKM88+8+n/9T5HPn55qMc+R/kxY1HwWtlTB40LRGGx
LU/+i061T/NFc+c7UsYOGHS75z+8TLFda15BP1diabgP/qNPVZHq/8Od3zTh/fllMB1pDlzDdab+
VII6vnCbrwkz6PAGGxAetW0ytYLFcqPrYQSo0nYNpPtKq1yeebhJjcS+El01Getuvsb8GPfwx3RQ
UWB+H7qVAqS4Xj6pPjYRnCYkwm6lf325EoXANLOrd5A3Z5EzhmJO0bZq8nKG1FF7jZrqYP68YgTG
qOblIVmQ9R8XMxfdzdE23wt9fc9j4Dhl217q5kV7p0SgDVgwUqNNAns+LMTId9OyN2xkH0lsy86b
BkRafFK5tuLwvpVz4i8KM2Pr7h42BDafavGdjorVv0JnBrKcfYF6sRERY3ZAUL30o/I8ibpJMEN0
ysL31LuHw6wi5TFNHvrfWdE2CT5g+gqbWatqR3STOOCiOz06aGlBTHx04GgzJQwZIrxL6mE9v8Sq
fUPxTA+SSkkPx5jTE/vIjiwmuAU0BlWH2PjzexOScYrbtjHsJP7uFL1RPTsE3RBPbWGRfI9a9+90
7BgSWWsmy4LbnpMWdaY+lh4wOa/RwjclLGG5I4MjKkSLMyo/WMOuADND3XILrP/hjv+lnRWsdJMw
bR+kMDoeHS/7tLJGsok/Gte8hSuWDl18805CqLDDNg4jnOKJ5+nTU1iGvMq8U64bmCE3QT3fXGGx
Mw1U9l8UD8se+8UugrC82cW8joCxxHt0/hxTwQVCDSxXEtJyAXvXFwJIy2xs+hg5/J6lzLHPzMIU
3XtNDCWRtNtyebkntOoyTTHe/wEjCDhdFxRFGoYMH1JmiLEB/hcszIKENzZk0xf18+byiwgsDBuH
zrzb70eejEXO9pZ1EyLZh+BF4kcghGtewKxBSZriCN9KnZhozInTHSzfCxW+CJ9uuHd6jZmq2g2R
g0shlwQdSCDaWrSwJFOJWP2Z4IaG1P9DVgWDtiNGN90y2DovWbQ+c+15fqqD1PvYQMWJAFsZWubX
qUCkA3CkjC/sIjgUlHt8Bm3NvXLStfgkGuTbSs0pEQM9MGJ5CTE7jjRueuGaKdMv5h0dCeLmFuOn
zS7NLRNiPMAQFY6PrzluNVEoe4a2JKOKqIjDVCxMdJPZHkslpWGYCp8pVd6m9sM4zryY9k1wLUGR
stzbu2XVGlp6IXjZOWntFt5b0Gt6qmc7n+26fzINls3cQmM8GzOceZ5GK2TtDskZp/qQh++3f2AE
6fPY3Iw/6MEApA3jg/BbSDEdFdhn6LyqCT4w0te/0wr4jmNp1Hz7Czjfe4u5D7n4ruWkSq4SBPL3
Zfvyj7kVzKUXd8DVWEbltSqLTVRLlrzCXUBA0T8SkCGlFbpUxvjLs9YWf/r4rMQOB3eR/iNeM9p+
Ifmn+Z9LKpKCE0O1MQlejaVmmReRNxa8Yz5WsC+ag8Q2YDnLH2GsY5ApCwO1wXSsuY22B8x1iyN5
GW9udErGO/K4iw6+8cVB1SG8AiYk5H7+wVTeLAkM+Tf9fbfj/5zcbnWzsW/7YL9NwjXPzMbSm16j
tBGRvQ5S/XE3Wm2kUnovuGAGswplg/+bByE6YtRCzGUdR9xLyTWbdSL3fS24elOry/TLtc1lyzqW
tZhI/Qi8g/+LadleDqnAOoX+Aq69luXwGnlOGxaRJwersZdT3d1EU/wCSS6aD7hWsqDq5FlwiviS
dJ0A5RG4Yt1lJM/h3Uy3yLYmp7UvEmb4pFA84AvJVtfTtEN4QXJIzRNEmVMYNqMW7i7u8QMCRQrT
4KJmTP+e7YGtOwe5tKIJCmb/KPRkcfl6ndmFTvHNY+t5Vcdplc/Q7hOemm0YkrsEFUSo6+iZ/BTp
dkf0RUIVFHpAqFCApmOToJyNqN6lYU0zHbCzWlpUXqsa5WLPd1tZdV+TTc7p/U2J2t87goEIVTVQ
0y6VBV9iBM8Vvd7vvvsjCqYZT4Ocm49fas22HXLtFISM4MixRpAGN3c507WR1xMbVz4Z7OGAekLJ
m0sW7UnEHOYyay3YN7VEo72YwAVPY17YKJG79327yiA++6Y4GLP8cfOcRSiFcIwT2fF489+c90xP
KO19ZYnbXWcMWla/udJqfQw3FrmyTtyuDEzPkFRHxuOD5w15ZcEArScwP55O9w75N549SQXJxXI8
Ro/RCp5n7lvXjEA5MIOJa/qNDtjJYoZWwDS2FmJLIIhkBeqBjvpAYTEPp2Ldl9N6iqS9pzMYHcgi
vMUGwpkaDBnqQB6c97n8kZu+jFmKc80NtnDL7ji+5AoVmvUtCWWhNPPs0qdwRFr5xzQO7t/YIKoC
Dt8oS5ZyYjcVQq9onhaWoxePbyPAOYtVM3zqY9tWLP3Mk1kYOJuw1IS5c7EcChtZshg+axCl1uGy
KplfFMdzrs3ohcEY46wWANJmkMfHjPcF8wEAkAroVbmYxbCM26BOuTQFD8iw9S7omYfkGcxeMLwS
Fu1iyKM2OdA0ag+L/PQuZHAHPG5aFd5QawZcjhEsf08n5AP+vwTI+0hHh61O58oO/Fwf18x+jkF2
1lUBNXKM0HjH/o4MZEdLpJB/6/OVGVkHalu2Ac3QRj5GkhNOiGJbodC/VnYO0ZaJ2U09DeA42N4L
bdEj/usLzKZ3Hseydl1C1ZVXxXjQ6PW43+GaJyffFqBEJVC2fDxnCj0vpIHlGcDFe+/bF08lwqel
z1//R7LPu3Jllyparz1sqtAcpEk6R4aVIQBj6ATwcx9lr/iZXvevdR1tj4nmlelhc2H8oCpS9cTZ
pcxIeEMJlwZfZMwe6SbsmtUAeRa5sWYWLOU4XbFjovE1jFHxDrU5O0G90bOcZHPRZa9zTaw2OZ2M
G1if/mE3EqmExD+MQyHZnvCrkLdMwE5PpEb6pAaTx0/yoXJQhiD+kwVToqKdWLjFP/TOYS268sm9
DLt+TXcI2mGGne5nE3H01pKSXDj6aMUmRm+PIfU+u+46aHH8sen9bM5g9u6+1GnSURQmdlHtqkB6
F1ShNIqatb0647Y9j2/gIQxW6/RLD1G7TDVJXnKJra/xKvzzhZ42BY5MBJgrb9GTpRFNBWqAycxK
RDR/2uVcOORc3xRxeCJkCuDZlNcqQxhBXAc5B95lBxRWlagwLaZAs28ok9xLeAhIREUp2orWzIUi
KC5X7JwO/4uhoF2lS2G1ocBm1fg6+/fSikfR+OiDmcUnE6MbECDH7mIvcTiIyG0XtN3ADedDD9kv
I0MeNCefPAxCjowmJ1dnMm7zV0RAdrafuOUhfYfCJ18thsHyuiQ5yf1OPE8Ei8D+O/Isbrlv4OKY
VS0+3/r6/eAW6UGAdRfr7XS5YOxZGKgZEb3rudJmFcAFzcpMRi6DqQHnsHoAXF3VXIyUW6fExkDf
9o2mpvRkq080SQoHGaRdM3dgJsWYEoBemLoeFX0v4GnGyZOkDlYOfOcuohdJ0TYhOYf6+rbtxfKl
MttEb+KMpkTwIoy7ZKctiJgPcEDGtoB5RUnz+z99XJJkTpZpwQ3tAp0F+CA18uvmIx4TuKYkBl3K
LfQoK1cKUsRii9ZkdHKzq9wEuIwjnmcXm5/YGVHe/tUdYM93CgvTndS1cZ3gTLn5vCNdtkjWpeSK
bqDlpvQzKORDQHan6SCq1lRN7T7m1q65AzaSpM3kviLZ4+IJGF2cMQ40HPpT/nrviQaYVn74DXbg
KmKf/753qTjP9P0rUNnYSPbUyQWi3midQu0bIqMzqJnFg1XkjMHPwVtz3CiEq7OwIi/g150dDsmm
2k2GM9EXOv3LD3oHbp/VSJpoUH9VdKNRLgwZW6lXt3S1AXrE1h5ZXwYoTZsTsvf+mEH2VxbBZp2x
h8+Nde+0JRWnm2KqiE1A0sQLFuRIbqdV+1yZKo8hKK2uZ05N0x68x9sFEMye8ibtHxop38oVrrKX
J2ceKTsUGh0RVXvSTt0QaY0Mj1q9kk4X+yLoQRtsKGr/MqrU2P4oNu0JMZJszlKiP3SeSLQb0h72
zHzFSeBV/vjovMC2OgDhwXKDZ2CIHhKtysDWiEeMpxlkxekjwOTZg4t1bhW+Xz9mkRika5EE9kJM
Eijcu9Rmwv8FtI+grmoaCKDnj17m04ldg+4a6crkTKhJImojGcJ81QmnKLktFeYEhGmcKl2jRsov
Snhoz0cRu042W8GyWCf881/dsc6Ba7HZEzB9z5l5LpWZsZDkMFsPupKhj9ch4gmWA7WHqWZKhg8j
RJy5wVIzNfbBqpiRHH25Mbcj8gpBgLN3vYBUh/89Y4zf1crV3mfhv22Qzjwx8SQMWBieci6UdfEV
KGK7Rl/+TivSNP9Ch6j/eHg2p5vSJWW6qepsfR+qlyjEl5VeqHYcppa+4kjXNDJs1RfpZdxsA9NV
hMwp2/Gq1FTjJdCxrYUciLoDX0k8wYe2dgDTll9xNtbcKQdTxlVn8hONJv/YZhrHhDB/LNF8GYnR
LqDJQrD9Wi5yJRalI4omAfMUgRk6hPDhMleUSWZ4Tqgc3nS4xpcECRragdeEgnBUFzZPJzXSRh72
qeuBqtzK0gkvkdvxKMrkJQV0B2zH/g4u1/meVnsnFHYTEzgqSlVtYD+jkKgYF1XGufwSZ8ZXAxZl
M/9nbmxruruSvx7S8PfA9afXXjguP+iC/iIGveDGqPIVOdqEthjV5E3tNQi6q5eeQFmusjv1ttX5
QGYU9pnTE7H96yD4/M0qij2VUgEDY2FyIYUTj3LpepyDtxMDijYBTQCoxEpenqaR8A9lmRQnPDQr
tRxRvIPcSV8MydgYsHAsfHvSMvKVDWa5YOD7a8HzSlFTONmmkwyI2LEBjDuOOLm30iRxy6FsOrCo
H7ZTtNkowzVe10aK/oWK9ppRGVfUwaCtAjyVyq8yVkvl+N3ik6AWafAOIvMnG6JtzcGVzOxWHze5
mjeHTxE1cqnc4+OVnutpfvf7yEcTMd8cUHQkAhdXiLXFCdqFl8FUfRW81XHKj9BuwwourVfa95qr
zxfQvwekDWs96rQdxH1bWHeqr3dmB4nxhULx43IBd36SiEIclEEynpjL9WlzdVWbQLPhNV9P7v8z
ma3IvrHoPHGaB5jnaYa0mZSVQWixHsSM8oCOgX3/bCrtch20rST+lx3KQ8v/kMeJS5dbiekzEVYk
y2qresZM0Ji1hjVQuahkWrRuHn47tJQDq0l5jviajoBFo7OKKwFaZbzr23d0QhIptu/18cF7iOJ5
yC/gqcvvZq83e6gF5m+xfk+6CuSXztqb4tcgqX3ob6mx3PEg2AOVmsXTlfE0Mv+az/otrQ1WGIeb
2B3N08JL/NlNnns2MrZotsXGfVxH2LSvkuCL33RkxPTETsXV5SlrMLxDPuNAukqmmy1FHNKx5ITX
5VIhpTNjqT8WIxlej+AtQvSJdUnGwKSpulY1xvwYx+UAs5wCCRcdGmKpr6Jh04+bj0VapS8eds3y
6ICPmEN+CLgzf52qY2ik8IKA3e8+KG3J8/JY4doC5KvwejEI51TLXmow2Gw+GcOSyennO8YMtPSI
sVDq63QtnEHYOXvGKMhnJW/RUXCWLYqYG7W/H3DQGmNzk7hBmsZRanzNS2CvHGdah5vv/FzCoB+j
divbH3OrCFwxd5l+YMm4cS7UBV4jbPIm6iy8yaPF4UUNUGvYLjbKpRQCH0i1bSnzTEiEEDerZs87
gZP1+8h6PVusCMLFGc/9O6YjAnBG3A/2YLBT7+dgD/ziYPny1MWLLJLUmCNXiDMpXRB/AEs0TCbt
0f5DstD4W4V4HwDS/qRFKnNPJkYoZCDctST48OSprlNr00d0pfpC2defPJvCil7X/1NUwezLFrqD
MUVLam6XhRC0klPpoZbriswnmiDZxsbLv1FcEVJKkTVQMe2/XJKIbvjB0IFs866X+G47Q88Cpido
uZlJVaxrd284GQAEP7QXYipLDj320BFRa4zDCL3rUf3q34LHPcWtraLjgANABtsBdjBZwTmsNoSj
DPD7fVetKnz7/2FwKKIVerZ4t3htPKGLnuI1bN/1EEguq6+Ig7pimL+IFPucKxBHpnJjG5OBxmVm
+8ES+sLSNDQzi0iwwjobRRcpxh1K5ZzDpvPn1sRsPfXO3iI1wKqd8g+YbvnvAFTfZV0jFx6C1tEs
pVDpDtYiU1Wu/Bi+/pqGGcY4xKXmQUviVmiaXUE2oMArfbX/hTkpELBJMum7T8y+DlGrNvfy7i7o
yu4jLvlImK2FC00EWEeMk+uSPfFJklx34+PYrJPxk6OMW0h2hUIM4jQUDZEK4zqgAmsPwWtbWwYx
FEHDTe1WPhVEF1RvOiLcaEq4w8pSr4UT1WLzIe5vhHYeBdUQH1/2ZMwpT+OZ5em3cJpWPC38A09t
6kB7zwM5NAXU6vCXzo63mIgttsf/zM9g7loTWUpUKnASe/nsCaD6RvOP3gMUdrWMGtffLNWsmjcf
MQM+z5rTy/bLWT5zXXzDChN0L0xDH+WntaAD11+8nfj0ZJ+3vWvZpCljxIIqxI9/Ab8PCm2cycvo
89vFSf7lljZKSw5kn7nCv2Kdber9nu4T/3MnCFuqbNcXEFToCNk4pIGVAc0mcmGtH1ina0xQoe0x
GM1voolY+AqFwlucoSSuT/NcokStFkwUqVY7+T+PcJxUHSHOw0MZOq8Wz5temA+ExLhUldXQCE3m
ybA1+j732d3hiiD9ETeLq3PWtHGRs5e67i7FA93veSHJFTPf4vXfAeJ9MLa/WpP4DnuJb/RVc++f
nwCQcgc9xiXwxTv37XtJUqPk6R7WFqC3fgMYPRs86x6m5FR2vkB3vGfZQCe9aP3/YHt5CTCZ6T5Q
KvLMGCdQgC3ak7qeDiXzD6ze1wKCIif/mSJDTOnytAONpTyjj3CPfJeRbgiyivmTBR4D5fbHPA7R
VPZN6xCyPuxJ8lMOMUWu0OMiMD+Fn0nTawXTsXGpOAUdFA6pUhPhW4CLyAqyyj7Mw1SwrfWXWO9L
WS6bBIKXRKFvRdkFGmFd4DLZmKEpu+b/RGhDYY9fYVrHEpjQDix9abtQY2zrIEHZeRzEA6PF+fuZ
f71q+r7M+3/Q5wksFhGmL61AwBHcG+W1oM40ajwKESJwTwUDIMykMFqe2cGT30oD8QeR8Pzd9AeP
xdT331tnI6br65T3kfYQ7WHFMfeqGSWW2xzvHtb1wQb956PewvNXRiloXzfVualvr3Q32WQyYfNG
LtwwFH9ef2OTtiWYfKsdCImlAi0mgeNQUuT4ywzgezjsUeip3G35gxxy9IDJwJw7p4QQsgQ/MYOH
Bb7QpwTkn5UVb6IrK7qV4KQTy5rOBqvgeFag55C6Prc5QEau0+CzeN+eM0wJLXNrpuWNCkqrRos5
TvYlxdRTmp2TgcYP7sy0A4O6LvZCxMjZYNNcEgYn6F+ud4MHWDS6wl0wKfEtfvmMxeiMAcDpmNx0
qQe1wVpqz/ahL3rH7lFf1PoyhzlOvJIo8+NpWRoqLeBtd/ISXo267109iLiJn64RknMgfGRmYsdy
pUuxDl4UiSWZp+MTYHeyS7pfphaeDIBpOxRk8/rDEgRbmn793k5pLXaDqXK9UjwZZqbRUy81cRAZ
Ws4BfsrXnZAMHMA9Klxznhg6JczK8PvqvksoR+h3nTlQKpZUHHOuzLpjuaAd1msCYw5e+rJ9K4p4
+3x0evmd9hk/wxfg2LUaXe8L8idPZSY5gZsSDr97Q5cZ5Rbeb0QDPxZXE5jHMRYBkWAVum3DiMhp
/HVRSuur85/MZtqgK/paIZYTxiI36Kb+3p3NGCMM5fYxIVtFtVMh3A9qeec9gB4GO+uJs3TQjBpW
opb5tRjjiWj3A/PnCVVUM8Bg+5CxnkK45DWg8t/1tpS/GkwcUWhwZ9w0LWEb1rF4lRfhJB9caliR
82JIhlkb4RXDTQhF0N1AKAK678NWaHYFUOtEzKAi6UeddUjY/15HNxqKVeYOcZW3JoMNUc1RFF2g
lT9GH8jqU3jy+aIs9xuyZ8KzBMU7ncOEDniq07L+Ar+kFdznAZ9OVnUugUoaPB+zWTThtNRL5Utx
tLJ5acYq0phJRXtgE50wMe00VaLzZp3pEK8akjBIUywqIkeIAZYXeLGRlT3ub4oa9deU4pju2NXH
6cpC/7knIhT1KHRgkERdPWX9kGTji7cxwIHLhMqtAnsuXgIaySgEZGzDSqibZDVrA5+7cknWQ0x8
Tn647MWdq+KRhJNFVo5DlxdzEWhpf2yN0jj0XGV0lcad3UIL2apZpofrbNyHoFi+Y3+y+1Nl1Y/g
pajusle3sMtIHlRGht9LtNkkDB7tf/XT10R19kgVK9hRKjTfF70/CYK7zgPdI6nX9QqXlWFjZTwZ
dhDy12l/xXt/kyQl3tHzXV0ui3/lKCF/3PRxHGwsryLos2V5ncAozyaTdiN+WIwca6mm9Yw2i6jn
9BDXvpZTe6TeMxf7sYsRsG+ozWTbY+5ea+Q0Z01/iIvoxKUNWP2gqdK7xbYFqS3we/03Iy/91WPa
n7LY4yFW2NnUMRWaHbSximm5WlD8UvFaLMBMWRkyp0Cm3BMvcsBR1Hl6x1dGOwtOAhssqlRxn81E
9+8ooRlkHZmGNQNRvdyTM9TpepO6KmRf1cFKGpCdGvR3FNOcrf/+hTekQ1iGfG1qtqAEyrIyb+95
BYdV0h5C2bIeTjQ+ThtTSs3f0YgLqXNvHmLCtfjc81ownwh1eCU7P3ymW9qTBpKPe7rNptoUgrIt
ShWAkfjIBtq2k/wuQTkIu59WFECy0lvEPqbFfiIdZLUJ9ZdAeiGaUfi8ABGx/1H0/05o5G49ute0
wWxdB5RaS4CFYLM17U74zh+Wd5ZgShNdOl3GYZbF/OTPOpSip6DNw8GcdN72D4e2M3i5lNUl9bBu
EjIWpqM0kRiqfh1BhGe/COzTbZDLTawDQp248vv4bWYp26e4EuztC2rJvptUTUNifRazPDFUGpLu
Jh4a0jqlB4KbnDkCVMH6l0HIG6csrwSB+y0tTO8OI4EMG8ddr9I57x22dVWv8Qa+VnMqqVAxmozn
csxNcVb1D4OLBlhlOD4IVQ+OQlV+jBHnKey3ZuUseIYwF18p6tEO3aVIXQaC37yr7WKMI+p4BPzY
/sEyRmgxa1hWxt6yPjc+1Y9vcoADXgXre+pQ/ihmPhlUcL2tonIoNXQpB1dp2pIB5dwcNa7rqq/p
0cebeqKxMIHpILIgWLkkNxxss9I/Wh75ljMCItybnOKXVOr3PriRjE81E9PFvy7VKF/8R7GfA5lI
OgpnbtXsJfklo5pJ7uTXR3UCmNXW4g//YHrdvoGW1rBmr/OnGK3/AQsB2H1M7GCoJ3W7V9C493aY
3n1CAHKCQRk3faCr8ehEs4I3L6g26RnyTFLYCPeaHNk8lEA+c4htDsp0pYGmBuNiyuujgFWwPId+
WQ/rvrEDL4+f6/xIcoACWINGhgLEobnSmgNbz5Mn7NoZhBw/TtyuTbHfNWac2iTX1h7uVNryEehD
bCxqsmhsJMaUDwUkpiLJzh94dDNR0x+/Vxcw7WKlK/TN4wMQH0SdMptzHphzg1AQDsOgYRm0i4h3
VIOGYaY2PC3KFO/OUyuj2FugDxEbkhSfaIsl/XwKwvxToCRdT3tk+055WD1asTSfEBZ2cxF1dFW/
8CY+5AISNma/OEEl8oG0WH8L3FJtm/n2CjKTWKkTefp1GEw1FsVhDCkA7PEBpadW46mh/eWyjdlm
qQvxxdIObtXEyvUs97QJZc6QxSRRIZgbMrr9wryfUDcXmHBG81NsBZ0266XORC8ezAr59y4+Yclv
6ZVlhn1GOLWeCKgf+RYXVUUPgCY1OxGpAked5bsyQopH2l4e6a9kLE3461FvyglDtk8WKS9C73eK
0Dz5hxcBGQXRtQbgyNLm1mAnGqurDTxkoX9SNI/79PCqN0ISB+/r4MAjRTb/NBr55cxy5KkL7CG8
Q61kAkGiNefuV8pZmwKNilEgbjwL2kW+VYWYpHwFQ+pOc/38F6h+a8RbtW/BkSahRATNdTheTstF
I46YnfZ2+xDzElwngnKzJ4uWLQW5RD/bRXx9Ae8rTFVyCCnQEUetrtVXc36MpAObPVmlVd3UV2SY
S48NBRxzJNkRQuYJPKSmeQr/R+macNhsp/Q1LK1kS4ERafZVtdX+RBQ7qap551mOcFs2zEhM0t8X
cv1UmDX1jNSOjQ7oWevKGL85hIzR6iUuR7cF54t6sE9egECfJcvgTG2Cvdszu1meCmGv0DxMtlx7
JNtKbTr5f9MlQnwKVJINAwVHy40zDiwjbckCGHZDKTh9qNXsOcyadcD9ajc7WDJy+JCOucjqcP+x
CHZFxw9HbHKfqjDJVr/PeV6TgFIhthKz29Z/PEQ/HxjeN0xBAVXCRqKnUkzDCmrAAPCIbnh4Spa+
ZHgCF+qqeIK0YyUrfb2mdcuvOO1J2A1PiLlmjlnhd6fe+U46KCwlmmGelqx2ao7QOoScXmPn4F7G
YK5kXe0LBUyxk+656px6TB4MVuOSjkR7eGM0ZN+bLynBLBBjBGhKj2irHLeyBbE7rcSnSuXxDpIU
C7oVXHEYlaiNYEkdebnhkOahUo/6ItXjrAsaB++YDjTUcPhGo4/1T7Mg9Aw6dr6wFAgJyEj+vXjp
M7WkmJSinklFKmKqYrxhb4OpDTyyQ4Dw29y7j29ZyuHSZZv2DfpXHtXQCwvjWVoTmjjIRy0qHJ6t
dIN7+NGRA/erLRcrJWX4QSdzW8DFw8Gn2i8UrYDz+s58Kvv3jiNaFt94N48j3HPIMKauz0mG/CY1
PyBSH73HA0ZcRiL/1N6zk08E+eDPgan+3lakN3GcKBjV7w7ac1wQeKh37l3wPZ3u9kEtfwYEwl5c
32d0LghcUprM1a3sPAnsbW6W83EVaqYaz346zlKntdUEby/MBbpzHRmKSzaOISayQAXIqKSlA8um
lhyiL4rxLgLXI4lyVTSSVTJjvy/S5iwFviTl7J/vQieVMcs0EPppUHAjzYYpga7oo1lpVjDhOKT5
44TXa6+PrgmaJZrxocMI3qHSEOD9QR+OTdgtESs6DOZa1ASKwxZTrU18T6aZBBHVWHaRHhtNryEr
+Pcx5Q06ur3frZM1kLk14phoI8pLNYJ0fCAhBBVOAXbDbxK3BvWPrrJeg56daSYXOplWL62dDDNu
E12u4y+ODAxHNRKWeT6soaOrMUrYKU2zEHBBoM+/SFlOQb8c8jBtUv5FDpXompktTdDBTMgycbYu
DvnDVG03PzDNU8uqU33bquwC5Nwg96A2xTf1gB8I691Fx3blxxhe0Trjhg33mOKle96kYzfc3S35
X1E+Qv+MDMB96eiiqVHDRFmGAvgeV5UTmA2MVgIgdq3zYSZ3/fb12dPrxkgK98oTd84p+y0Y1SjK
ByvflhNE9ZTAfZ3Cyjd3sRq69gxSdORKLZ6Uk9FFLD1mditwEUtYz+fTg3MRMJC17oH5tT8krGqs
J++JvjWZybd/9JVPKaaYPfcRPgHNN51IxP10oOV0AlQ1csgzBxHK5MDHHewmQsAMOveILwz5vyQ6
din9YEvwTSMpbvpghIgW4xIiwS1CR4QrkBTxUVUaqb0+pimBZwcDqIkbcVqAZX/hvSeufK4swU2X
deil7U+dHz4FR8co4cBMyRANf6Xy+xLr3NF9fPrbzExEpI7167FeN2AerU3JmjSosdFwa7b7+yLD
YybM7VkZOLu88+a9KU4JBPMwDkampZ3JxgEGWaWTQ4Y+jyDcneKkQProCS4V2sOn+mcs4TNjYBHe
RiLMZ6fdEb1L3W0GvHh7lUpXvcodd7jeJxAt0Zr9FAHTqMspLlwyBJjKTeCj4GGkbYPWRnCPEqv7
abRh2+a4EtLANem3FAznqPMRu8NMzAdTzruWw0eOHkTsehEFJGnIHIGLY97Y9n3RomkxKWv9W8l6
FVwQOjIKtxyaeaQ2fWL92lXq7BqM9qMG+bhg/qNEnnCQsngIo1r7bNYDQnpYrhyJnjM3auWQdjaf
YIglcV8w1jv/9d5O1D4nx3pQedV95KTMmJQk6IiDXlab/0ryD42D1BNNHOBjssf3kUKOyt2b5yQE
jd04K7Q9AgtsSnevs20q1EucPWTpoYxczmfGv+2L/OtS4RAlNsgH3Y3lNZxmWCwVyOsSjXYFPtBW
P7xGO2vwGPaecb0mPHIhzBoWbQgZj6634dUMkU7JGyb3mklrAV/5GbVonVjPfVbW/bwL1mF3ORCd
W/26ATcv8P9jsGwwz8y/owvcb/a+GrwOqlQROpHtBrQDtcEWs9ivoHSut4SERNbWlB0SOQuPBREX
IHx0YmlS0HHhmd693Crx23R0130n00o7g4x0fVRirnBmuvLu2oApASoWMgHHg7mcm5sT1MXIwHQD
tkmY4UEjyga/FW7mHPR9o504Wg7ARplyt4Bd84wb6lhTgu7DyKsk59xHE8L4ExA2rPQrWIkoV5Nm
kraFhXniITpNID/hatqw1rFk1jFUz/LKH9Z6IgZQtwOgz4ap97H2pe7m41vkIRZrvcyY1OWCViOJ
6vu+zRgv7vkdTtHUf/pSrWlNwA2E3RGzyDaM1LDTEYUXIIR0kD6JJ90TI4K2mywnCQ24yEjtq4Zg
Z1lWJbSeMhSg5HPFrE2aBMqGVzXlTVYbsPCNmp0WJ14MwHjG3iexmDUbNFaGCP0LHRiKZdeFmIOA
rWzhWPy5wk6D+MkKBYk5iODqfiPdmsjtGSWX7OOnfjabr/tcFdhDRdhnJd2yDyzEyG/n4JKBGv3g
ohkzEMiQFnh7AicpZ4mtZLbMlJiBqSn0c9a6BYjpAwF5XbKSqwse7Am1BEjNjGM3br7tohaTcwIt
83Mraxjq3kVpg2fskoe4E7QduOiQjb6RiOZi+hJaWk9XlPWKm+e7XUoPhN4QDnZOMyFdsBKAeCHi
+w7OsRuB6wGZIxJtNZikcYUOLmQqjyvA7dkUyZIrn7144Wvnr5BBwQpO54nT/uYrcq4O+X4D11o2
g0Y3myjtWQ+sg11Hw5Wijp7qk28rAwq+vQe9PoR78pm0tBp4fHfw23FBA8iV/HWK4qFp9N59L8K1
R3ZNHVoraRCSjwttPOg9QDKglAuIjk8872sKZVr6YY8KbSH9LI6WT6hJTAre9idDGRsGnjHLvkXZ
uJSKa+Z5IM7bMCkWz/FOZg6JVhHcIAmFvEwcNWLwrHXqYrT3DV5SKbkaUPEm+r0jBvXdAA3T3pDX
19YgKwrIrZh1acxR5bSRIh7xZnkGWmZiZtl4kOE92Pi3+FFOuiBgEYqj/mNM3KqstfTGOMV2vq/6
steipxkcVCX9ErEXHIsyMH7MgIybqdSAOPIhtXgzlmeJrCOLZvOrqBnHE0sdO9AETDTi+FLir2d5
T7bt8HQXqQOvqNQ1/4kRlOWYD8tQ/65g6hMsbLIWKhIBsIlVJEKFm1YCUPW/g4/Vbck8Eywy/C2Y
lu2dXfp3vTsA8KbZgL0sl2OceZ/CzSBB5TdJ98+CSYipD2zLn5QIUKsE66S+ObpgUfpllpqgbToo
U9+MM71jRjtVUk2FLtqX4Z0MLl5Gpc/v0ZnW0Br3+5PR7IeCmkzUegM5gv4Rcf9YDxUngZOPkw1n
OGXxABuacryNtOsi8KfMgMYxtUYdFTp85eAYERUdsImgws5wh+NVaRQ0X9WGAPiD7QxgvGA0q06o
KXBLK4qFhVhC+XR/VGWxHk75LNxoi2UfIyfgF6hNuPBTEASsXwNQtEYmpCFU4xhUHHgfLPNnDeKV
STqXweETNEzGeScnym/HD04IDI7V5FZ/QNeFCr1gpBHChc1GYgggId1uFvlmFszYXNAvOJhhZ7dX
1ktrzy7bDW6x+ojJqK5Rt++2gvaT4y18MS4KBzcGF+j/+Z1AxLaQz1mCMnhqKEhEydbkkgFX4Tzd
hyS/PPKxpIlWi5TrifhsxgZUj4M6mN3rdpS3OG9E4MXP0oRxN+eDrOSa7dXqo5noEHtocVctTSJT
64ASPAYflu9MK6dzXFbopM72eYKHbhEdUHv73OwUG1lWDn3T55lHMOfiZ8x2icVekNJjSVBtAfge
jzWEdfeoWIsnfC334yHyDHD63/NkXRXOJR7udj51lJqjnijojPJM7zdJDUFEpHrR03VYjhhIIrH0
byD8IYdYLtRhtG93NIv3QPKxCRvbR4ZCHBZLtXb86ZHix4JNsRLLQQGAby/uPO4f4Q4bJy0mp+bm
kTtluamtGZpbq3BFNnqx5hE0Zgl9q+JvGEJ/D64kPldGsCqOYZniUZmuWmPEh8kDvsADyN64PYrw
i2QFbBHHIl6btbIhV2dQLdM4fPsIyoqm1Mag90UvyYQrD9pMO/VgayVH5odXiJEnMlwDMVvTmb9F
B3b80U74bUt0peyQUqXHNjmsTIwZJ46xs/CLPCAF6bxlbMGWQVoyK2BbiRtO2qeNU1KKqbim1fYs
wjzZlo7mClalLd37/vjWisctwN1sFoMcAx8Zr3rRQvWbw9WuGdlDtNbExrGIQmZM7K0bSyb/l+rI
7n2HRPmQAw/GiGeGlpsWbsNunAUXARBKzli0N0DIhYzvl3jDHj2WkidLvyuyku0fWQdytJpjHYOj
FTdcD6JqYotyILVmySZ3FvxUyJzZMoncNucA6kgAdBnsU6Wz3nicf8iwVuyB54QAQ77ZPRtF0cQB
DrKacLk4h92iEti8Dn9K8LwCGKBgWVwO+SgJnS4mbPTtaF4U7u1YmtBCRNA4sKf4elwqmD8CFyTv
n0b8mFEd/7ZgjFbJwHHWz5CXKjp/AzSDwt3minlrpPFKnqb5lvO+IpjVFQEjWQ2fetgs3rqZ//En
SROpvUG4l3bYMgO9zn3sXzOxz6Fgm9uWgw6oODy1IO4Mm5O5my1UUASP7n9t3puhcQ3Uj43yBpw9
dGcyGhJhaYaLUW62CaYLUO+3Qet9IpDyzxNJcHzd46UBnmt6vf6UnMZljSTESec2JXpwmShUt2EC
SkfLZ9gaR4SuJsnbYTBUkU94oaebLV4l6DktuazIM1UHMdxhfWTbhdpG08rlNCgBKXUlbCq5uz4J
wyV5RJKgRO26JYc5DCpQPIoBSg09iAbYORKESM5DeEOtfuOecBhRCyPJh7mY4S+cusROsKvUrJ9A
PYWvZYH3i4Q7nDOjFCmr9CrkEsUKUczXDK8lTLH3UrRZpYJtKWSV55uVgEmAQMOxWDmoA5ORXj5N
C7zZ/eHfduA/8nA574rTM5ExNFEOLBBETa2WaVAHNbj4TmVvUpMTkSC4fC0u9y21d4A5MTji/mXI
h9/jsLdzdoXSFDMWwWvLW8dC5fBzFomyGE+7VqsW0rs01YixpEW7vS5eYpR1BORHRmfBIjPntSs4
2lUl9a59d3eHlJEpUz7n+HYp09TEMhYs7F3u7HFPrncJxOKxZvGGZJTjlUifBzhvXhU6FuvwrvHs
jHFfh0BCpb8SuvNbaqT/fJj6LObF+TCEgFp0yb3041qfiNi5F+K9cqerAtKoB5dkSzZqib2M/SeP
36F8lP7CMiVzaoGIhQdIFnFy6zz7gObZjJ8tDnp+lEumveYYthD/HAAmHyfyAukpI1zDTjamNDtj
AXIEkrBAkrux3vr2GB/1sbOkemY8cnmN3zLH89627G2EJYnOYnhFk872jDq51PaEroXxoCfi8plt
MOog02Xi57N8lGlMzhoPS95lYgd3oJadJC9TtW6LRls5MeiP6wqkThnPfdBljdTGmrm+ar25/+qr
wXMDczg9lmDoBs+iqBNrym1pjmUJXxAqPO48Wlt4oVPaVuC+aYddVhBzPfhwQwHHuGm7KXb28hk+
MADzrfAsVRGvD0/DuAohRwgu/BWnnXmRu9a3p1JP1EM9o63zRAwEpShqEuaWOVjgEonrEsIF+yC4
VHg5AORyiKKqIEbucqhgVOEUSYUL58np9L3dHq7gRz0EelI512J3EiVQICgTe8HSNO4n0WAk48kG
zzldGcaFUkdiY3rJ2moOcNkkyILmUnX5ozl+Jqowe/rA/rMlLKhBdOeNuCPGxQLUU55X9zY4GXsb
1XBu+lp9kFcIPPMPJkzSG9FWKa4eHAVj6+eBSc4gFVTf9cVvdvACLzCPLx+WWSpv4okGUfxEHg4B
H0qh4dLVnWifgIwOzctrS5Al2cRs9uFFBHyox4pPSTsH07Lq6LtW8hldeCG4qYVNE73wRLIJD1Fe
f8naXJ1BRf/scWErc5sW9tzRsqAJuBWZuKfE3j7hz1hIwmax6a1OmsVhLhB9WMrtzwucS8uPsRVX
gpohdvMllfXM3jq0NOo0Y3eDV85id2wqGV9MwQwdSXl8WYByNiSza7htGQuFHKVdZNdbMmCj2Vqy
apC1vuMwo5vgb6TRavrdyXrOfKpsC34CYKe4us1TFCYYXCG3/ChgFAlhfYwOfwuwtogunoVP1hTA
01o8JAOaZRUGobncLvdJ64x79aXzBFV+y3fMZXYUnBSIAe+Fbzs3T+54lJYhh3EBfm+QeUWSE0Ng
UhloKh3zsfStk63o3DLS7l04MM+DLMCOSxMOigIplpGNzs/RrpKxCW2UsmyweI/c1OLD0c68Vz2c
l4VsnQvu2dOc1Ki6MiA4hAOBtNeCkJ60L84g1G9V+Dego2u65ngt/4URrGMfX97bSphH2ePhvXJE
KkiSbLn686ifTf8GzaAYZ0pgpKsWlHl8D9vz5tKda1VY4mFyiigbEjyu6M/rJb+x6nFza2JT2GfM
zR7GL40VzWtbQQobyTmzIOEuhkX7900dArbxZzbXN0qNWA4PJb8UPGurXTbR41mzjYp7aec/XtK+
lVL89107hGXskLXtE4dsvNdhl7dhaoBmJWHEYhbJds70aMp0qHgfexzERNwJxc9oRddgvJFue7MP
lzh05+9ItAnQfjgRh4C9BO4NBhEEJPSPSTxYE7wonfFjiTfG+Z7WuDeKzte0AEHwTVWecyNzw1vq
wRpJWJI8aL8jblPdCZb+tju5PqpsMFa7egf2CDAlLWeoC3i4HhBOsXLksLnafeEoKdwpVUOiU8x+
ClEnYLjvk0GIoBvTopHZho+IwlZgso/di0O1irpttdLE8tPSn4jffgB1X4hktM2BNBcdnWMQ77fn
b3gaawbULjFeSQOUjRjmYCDbnx3pEn5n/8vyamB1jNmeEiBUs1w83nC0fiOr6gK3XFvpYUErfe8G
FekK+ohgibUH4XPah0zTCPMqTpqcDqvmrKBZiL2UD+5RY1XMJDzpBOMC30aE2DRsAVY/b0dTs5Si
TEZ/kRmVBmVIKRfkV/S+nL1qk7xeMGqT+1qAkzb1ncu89cYvBRirkhUIX1syk9k8P/8uVJMHXjtk
YwnUA1s9Vt2wqtrAuKp83k3OgEU+fHmByL/upZF9Z3gtFDynhqm/JhbU/rlb+9nqhhSGTrYsc6wa
VAmu2hpGT1iP2MdEg5mWpb9pKLl3WYH29BNZeETIysgQAXTArcshnCWNlNJSpeA6E9FXw2nw6PyB
hUYrqXBYxG+lJSXgK2xyuFWnSP2OgApT6vDIMHl5LqWTNGU7TzBnN1tS40WD1HMGYOu784HGI6bk
Lci7g3JjEScjw8zT8xggoNNP2yuTqEfDVfvn/UYwWfQhhYWkp50+wEZfk/lAtN6nAjELk3Npbyn7
6ZynCymeZtv6WtoRolZ26SSZT+y3hE654A8ZTFc9SumkwQdBGJ5O7dGj/RRZZ70JMkKDehH96BeZ
NqduOowsTzz9K6+fWkCVYIlmLU1NneEhQpxTWwesDi/5ZUlzl6gPP5Lx+C0dMfGq+kKu0ATZAB5l
dQa66J3WKVn6ZfX59G1DvfYjJcentGDUux7aZL1XQb5iKMr+X+jg/yyPKY50bLDHrO5Wj1FEAu3P
nUUtkLYnHKmQ+ajXZE4ncL0G2MnO2cHBLJY68oDidOyYpF/wMp98LCE3S80S9FzE2f9xBWGUamP1
IkwCSFLQLc/5e0y4dTMstEPXEyAeXDsUXTPk1AjZkJ7rOnNe09qKRfC3SluIjIv8zgulWS0pB7Y7
MKdp5l5l1nOyUdIY5p8hxBt+PYV38eYwPNX8HbZMWR9M0msSKV6LAkLElEBOh2ZIXpUHnOQ3YQpM
OjZoQ3h+pOKQygRXLdRBB7SAqdIqaI3FjOf06i1Rqwz1mcf1F3VnFwi51IrSPAGwmJOjMuxRuRrY
Gz3G/iHi7ObQ4s3mEPX0WFwzeW6p+9FjUMHqsKwP2wn9l/XD22imX/ZFTOdi4441TTSDJOkNlGzb
sFuCkskwyYQCUIKP8z8U4jYXfnhOBG3aSWfB9r7dPodSr+KhML9SSj6a7FaB8XgZzZkSQSVwpDvd
SQTotuQcOqrXBOdRuF7OIjfcnhoOeJY+jrLRaFFiOVLBQAFM31gv6rHe2gg5rOc1yST26TfDkdD2
Fbs+zLpqTOGvT4S/TfSMjn7Hwf997Kh7FKbWfnN0zmP0B0yg5Edc1LLs93/ZWM0caujpyFk+uPI/
igx7GAaJsH/B6chjcSz0ascwFzWIERPlO7KvLAOzoY0TBeIP52BsKvkhRn+hL5tYp/PgbNGOst94
ymNYU/vkUyu764ezOXO3JFHxVdMwxR93Bqm3QppuffPEiq8OS6CmSOEr3bB0a2MmaYp5SyaRrSWc
tZ0wxNWGW138sQFGXuZGzdftOjbUjYzJmo+x7d5EyptKgYRulsgZyofIS5v3GP3tYLyvfNd4vJht
rjLE6nzGBnyhhmOTqGSz4G2EBnQ1J9HdwqcpPc9iOYi5qAZTSBMlQRPQj0tNd7lCmZIhRDRp5QQm
oeilKqvo1Si9ERhzJ3sXy+GITDXk1+eji4LlsUvwBC4hS1C9mFlZVK6Qj8MLRcIhNRu9Gl98DIPy
JmUjRBtWMAryopK5bXWlrlYuoZqKxMZyrCCI0YHMf08bxLve6H6AJvLp9wfp8Zv570t/BfBBv/UP
owGEeKixOvmBTJu55JWuZQbykwjqOEs+tc0A2HL8/18+LJlgiz+e26lYcZ+GyaYUv1yZ8lLo4C/j
SsnlgGgjq8bVA245FGsfQL2TtTrhl2QHUwuCT2d4sYRq9BpU2rfD3v7tj66iE4QOJ9yD9i2ufloO
X+5fiRBtMz4aLsAARsjg4O7rdhfAKD5qSOubl2NNUz68orK8AttfzuWSfLNxUweJlsFmj53xVA14
EX6wbnTAvy6gLsBE7VXXA9Ka7WQ5DHAw/vq0Kb3vt9cgSmsXbP8dy1E5OU8Z7LroNjHCQvobgz72
ovaMTTKfeAMELxiV/vZcybXw3wMXij3+sGfJWJz6VPW9fh6SBnynsnEpDwjUp6XrSSWWqUcqqUOU
/foENwYQbmMiM7jeYzf5YKbUvsKsyIhBQ5/tTBql0CrW+XmAWqxseyV0AcRRwRxLBanwqq3n96Rl
mRuk8Nt7bFIVs4iop/O3s66+aJt3mkkLVIwFU4bHSsIqReoCsTj2ECeNQSz48hzkepjj/lnTSTly
8Z/nIX492BGv196IGMpX3tz5CYmckvfjhRqAiyMqjMO9DQdxNNbYiS9n4D3B2uLsyfg4aA7+tn1J
Zwt9L3MZAPwlU9g30cCMWph/dXqZgxPGIETyerkkqA33CnNNZurPWIiQlq4lHsblZY4cuIK6DRiu
oJF6uhvHfFcBBegote3kxRsqXKJQ9a1wiSwduXCuPC/APHb7tH2mvUMBRa+6Oi3KjAyGcTvcy2xT
4UKy//xKCAuD6+yxnSEfs6Lnph49zAH47NZP0MmII67XU4LUfpAIChFIe0ge18Eyv0+P7chJhm1R
23EE/6+feXHI03jU7oh+rdmZL6xq7c8C+tyKxkq3agy+F+/XgEQhYOfWECtI5TN3ybJZMqZmfm2u
Ig+wnP9PDj8fGReupgzscssKGw0GRsJ04dvb4bkqpZEqjZ3CwyQNzJY5Cb3OUtc4XCngo3wFX1w1
6Z/ZioDUq62HZwmRZWZtxMrq6sMtoAb0Hqqk6DuU5AnW3kXl5PcmErmgvwIB2j88A/CRIB2qq2bc
O2XyglUhxJDOzStV4olzxx7mRTZaP/dYOyM7Yfb0UPtBq98/lvJ+egFpp9owvofKEVUay1CENj8S
V4p7734MfrM6ov7gARN2M1J9CbOWvSUoKK/bU/4WJ2t5rV5qmCf2JELz74I/ay6FZsa/exon1KeS
kSnoGV4LNw+NpBNqm/ZmiQN9EqAqZ3Xht+9bhbU2yq13fb3pUuq5ZVuDfNxljQGYjqJBNvT+XFQ3
I6Gp7RG3glC5QRyn8tGIrVNHQIrZEfV8uP2x1cEIThMMMY/IRS7JhJG2uRby4OcGNDhGqTFqUYGA
xkdxsib20VXSNHiXHIw4hw/4ejDvqpspM9RGHYKy0FlEA/j04V5ZPvYYhPubOkLuuFR+Ikm6wuMC
D9n2y2ybB6n1xaqG/83wWCMLbsbstV3Nu4qwTJAMuirun/VYTXD568dFe+2uC1YkUCSvqKzlYnAH
LTi5qYAYwMGws1L2htfi5TvWDqg7/IUH5WaRiKbuyedb9+mCMJFktzpYhmdynbZPcSEwOFC6V9tk
upS96yJ1Qi4ajEPyBCseZF0aesf7iQTdxy0ibecrUxZs5tQh1WabGE83EMphUO89EeSxQRFq8x55
Mf8hC4bxoEH6Ox1cm0s1s6N3YnPDsI7OZ6m9xaa8U/bi72YmjAjSacdjvtjyglUMJVM0REkjCEo/
OR7mntuNUKrH+DqXS+3GBwLpVf+WESMnXbZJdnFXe6vw0L8WRi24k/McKUz+/Cp6y86IzjgRxroL
YnvNC9s/LvfcN6q3ZmHb3TNqvaOF4h5etMlfHYVhjMKs0t5W8BjUw6IlSVIM7P3QDABf6GTePCHF
TR7gJR+ne/++M5OTB2KV7dL3WzGwydAbd3DATLgioy5F1CvzRpGsm/ypxMyYl0L6cRufQcu0WKG8
CxjKHb/VwYaI2AfhuFSEe6yYEquee1HUE9G2EH3P4ptzfo0FmZiGZBUtKj+bGobVZBWbjhp0qeO0
Aov906r5MSm78qptOYsPSYQB+xpEMNqhwpJ5FLD1Nf8P68gKwEleX8H4UsbLponnSEWUAvwFhmwt
bRmSG5tIh1avFnTT065hBeQ5QZL0iAIwLFfP7aA/Q6SXzbhLKGNehq2sdPSoh/MQVaRDsuZI2101
47Ad7TQkeb21Tzf45H1sYk0PebuL0nmmDX8ts0xnEotjkI/KzEr7yBAtOO8qUvY2aoTt6RWtYOhk
5uycLZsUbWfDWm8trWsWAW5D72CZlCTqEABWfYO/JKAK/lUxI58OQeeztbiXUPOFDs04ZS7y8lCw
vS5UVtPuODAX9t0SC61JXS0q/FUW6XzESoE44I3g/FWNvnd9AU4cQVLGWTnCJMditSvrZf4+UqO8
TAMFBvghvvbSlGvrD0yHmC+A6inuoCm/NwO3JcHQl7Uq/85vdsJHtafp3swR/x7go/tKqAQd7gXD
fb8qfxdCBkE2qbSF1wTEOABQA0aR/gcR6NTYP7ohCTr1f5gI2AnQNYOBo4i+oy0WZ2v34kcdFw7f
i31yyYglNSQl9jRmjq8zjA0g4nPIZm1Z8a7zLjkajjbNRwcR7ghyCPIBcWA7MqgLnUzAzdsa7Y6N
1UNvqVPhW8dHDUeYbmSQnIgMAHIEHmWEsqDDgv0IMvDumn2X9vwsXCX7XE9j6TiC6KtpU6IUQOpK
o2AtNnKHHVQMEDHSUojON+cXX2RMtNGyfaHIPtnBtx/DLkt8iF9kcueJt/WjPXO2SofZNb9twUvD
GEt6XYVKOPUnEpjpwiXlBfqInlOKmcoRBU2iIhQG4xvVOl5F9IGaq5uKIz+Wv+U12LR5d/e3Lleo
87tdVwIAbvl9oCWm2a9XOA33Lp6NpQ5eXNfcLjO6wFc0ZC5vw1NNkAH3zWGlO400JStQiWD8LBV7
UAJaZ1z+2SwX8eluHqdggv0Y4nrh3AE9RT9+KU7rCu82GYoXALpC5DlA5U+HgXb+jDdbIyNzd/RS
mk+42tOVGevxP6gSKlQ/kWFusb9Oe08DRX5z2SZAQF+YBWjCXdmSwL3ZxV5f2i8TbkVigz6wp4e+
mmwUUUywEvYO8wh//1UOguvRQmH9wOewkxuOOFDbqSrcu7rjCFehwht87vI/rWNz/WxDWAJMCWlr
deGSbiRvU800XUo4yqeefOopnEAbKA2VMO34D2SCFmBNQxWPHNTNCcuM/9wDBIG1iT7vD16GP5A+
xf5tQ6KOZolkrJYDkjaO2w/2gFYs4jrjYVzzNoOQqtE1Qzh96g5mThJEyl3KV80FE2BlDhiKVGQ3
+Cucl6F0nsuFKd5/moTOtraDrwkZDa9+S0XOFG4DLAOCGra8DbUFaiirR9qn+IhEXztTcqYSMfpS
D5PneDMedJVMbx+XIwFKWWJaR5pqeafOX8B03PCvQYZrSE6g9agYXfpk7TB8RlYCH06r7XS36deB
u1YzWxKZQYD6hjNx9n9b5YvIVEyuxEjApNPMvnj3lv1bc+pXxEJExhxm4vcqtwUvyv5c8/VOq3Qe
zY56Ml77KIJCmLYRlBUomBLmq5HJhQyIabM43S+woPuFL3TD6GXdCXryJfrE4kqqmcjJuSIuC7tN
aHtD9Drqc2J58h8wJQ+eYk0GQszdOm689UCrhBCJg5DGvdoE6MKRD/HwEYs8FRNAHGojaO2I91yv
N455N21FNE/zxM85CZFYi+wMwu2AhHsPgT95ESdtYx+k6jGhbNnFEe/HiBJHMtNoMz6p6C59ZQ0o
0HfdlKueBHB/j5K7LGETYMk2fknagu4catQHKT7FPYqzMUz73/qq8Ovwky6nfnbFPUkVUiGWoADS
irXpIxCArSq5Z6upH73CrMe8+XW4HaukJI4cGbse6YJeS9CNlM7Vrkfnto3jDf4A6qC+oC+MnYsd
CiVrEeV6j1vCyRnvS02AWVQgkNgznulTn0wtehQgG75tq1948JX16TgnOhednzhgUns10nyqCACy
n44fw4/XjGyvzhEtduuCsJ+Y5pjI63zbe/cGf+kx+00fyGuAlnWAOlqyai8IVQTrMFnS2HPhGAGu
0J8xnPbby1VuQhR0bfvGVWktMzVzAkV1JO8LXxqY0K8GtDGfVrSG6LGMceBlCfpnSDMxSh8qayUH
SkrTAEQ2hjOsm6/vJ0aXQv88qGTol8kSIbR3BcY7Wz73cWlNWGucfXlxVVfZjQqzn7v+s1zLwR0g
EMX7O6fD+vjLWbP9vr9FTOywuLEAGIi6s2x/uXMtBhlwDrO3V4NeLThfQ+X3CeFWj1i97CQQaNop
9gbDd2ozPhPOhf7nZacsG0PXSmT+bBD2n5d1K5F1wzx+2+MGB2qrDvOYL+U9G9NYxHx3fnkcPxaJ
Cp2H5j/Wbnc9GPuZ+zC0fho3sPpHdkUldiZKgnzsJwc7aeDws5JGNH0dGT3CDInNfOOSeqyMTmrW
HOm5Obi0F6kgFcaXMJY9osRSz3laNTFXdBcEXJIomE+rXDCwKwvFmL+kZXlsn3MaGqg29nbtp4F8
Pik9SDd9CZdam6Tq7RZQSq1+s/4J4QynuDujrBzpFVNOs6kTH8PTHYSCQlIlC4Xzfj9Gew7Lz5Ec
GCEW0dNh+jFEu+6WbiVu9mPJuxsNs3ct63hj0fwHgHpClY71ZRQ2xZwE/d6k8Exh++LowT5BNuQk
QFXhO4YZ4AgKBskRg/IXQu7GRWSeY85eh7f8wwrDhJVQn2KQc+dC2l4ZncWQ1jKv2aomfGcPstCa
wzzZ7vFw71pl5Df0uX34k4U4wge8Iv6ARmgxtj8GQD5hfvJ8pVb6z2PHXhMMP3NCX/LrR60Rd6PD
eCHdEuLUNpEFWTxu3HBuueBczE5V9LozSbkNCnMVA7tAlpbtBTKfZjyzbhIkesoBlIn2A0UTYMUs
sE+FdemVkyF9vPDZLrBxNxw6SW8+1ViTGTbV4g/asEz5ArJrc9q1tIyQo3kfAvW+vWfACumfSQBU
s/vO43mTklweLWqCDjILFuuH01HFHKOsqG2Vb76mxLRWcBAgSXgsn4luCk93hznd8sD/auMS/QT8
LwuPHMKRUiJB3aSjNs8NcyTRv/pM+zF7oqbnNYqw/FP7kti3iLtRU4AkJTJ18zydiOSEECUiUKB7
8p+Kedj7Y7e7B4TWGcLnn8qgiFKsb3dVh+7FRk4IhY3p79twtDij3eLkcJI5+Gv6E7Zqgx2NRyUo
sWuUuJSIdDx/s3IiqrAgpTlA88OPhJwSo133dUQTNIQMlvBg2hAayBGXjqgs+Nt8Z4Kz7L7mTO+W
lz/Ygej7g+Gj5fGhkWOD5ggFwYBaBibGV5udng/x0+95Z/63iYV4AX7LBKkVE7P+3UiF/wugmrm2
xotjjgS+7UMZVqxYRCLeuzK2aTr9vmasg6yNYk3suYHeWq/f79Q6miV3LnxjIac6S4zQC19pQZEq
PZJjyklsIgbpgyvSb2TTeEigvbcnCkof4i2s1W5Z8qfVaNTX1Y8pZUOcojyOOi5kFxKI/q9ekS5o
m3Ig+7oYx/u6uxLqRaAEsMagWTKrjBxJX3PpgIPLc7MFnBI83LDNPshGofK661an0hI8izd0lf3w
QMfeusBCUMQL+Qw+WBKneFl6vaE9k8gVI4wdHUEgwMvcY5FdEihfO212XHVBWkx0Mip5zrEkKwF5
wjQrnRQkC2fpL0sUbgudFL6TmVnFNRh1C9eKHvtf6+RG/A0pVBHWlzuQqjk02cWb1EwNiHjj7SBv
4bjTTD2ZCeHVFbXaOIQuzw8XtHPF9vrxZzj5Hm9tkgH4QrgfY9SzWNc6+NqAyMTDZi6AVcj0oPtM
/84ZfO7j2JCYNNqrLMmcbQj+lbcqlukehDQigWI0bsffMphoxcyTTbI/q/II2TfxfvSxQss9XTlG
2rcEgLhDTaMnZSm2i4px3iqjCme/MY3xIeSI1Jvi5TGo1Q+YjF4QslPZGFbXP0J27eyurObO+PEX
6vhdTrmzJIzrBwWMJFCIt9ns0JWES4RB2I+fxdGIW0dxc1zl7oWQI8IZovMIeTGGmSlh5pC7eKhw
ZBR3ZWGZm7DNyOytSUgjovPS2PG+dFeaBkQ0g9N0Fa62ybau95dgDHBED5QVLtxZUtk8ZrI6PpUD
CZePuSq5wdEwI3+b7/K+gpK/s5u42gw7AVI4xvoGgf/R2kCk1B2Xa8yDSqVkdmdjkdVG2IxyHi/M
/4EreC+VrpDybtVArvXfWFkKnlHwuKaJgaIaO4Ex81lX7nUVudbmUAwptgyvn/Iv9QlHACzB0e+l
TLbK/tUcgB0eybuyg2AdOGH8wETFvptsV3pBdlm0gszyVc+ksHFvqUpn8yN/MIEmNZ3NKH3HAZoC
g1lxdsokS5frN1sBSBpBcff6MXy9n0fOOYvq3iSVr84KlssXppasS0WM8hdqNjNBHM9RyUwLkDbs
huikTs4gJdsMMH46Wyr86ZE46vxRNToX8UdoFLZSh/Kz9XenYNqQkgEY7bQj93xf58Gc3aO+OpcD
lB47wrhea3QaI+PXSdckhhUeYwvLSEfLOLgIGnN/08aP2j9gov3Nh45gE+BzD0lt9gGAG1Qre4op
hfJnCyVT7djUfwE9Aii0fWBXNSBkAMJKolrkgJmKNI6mC6LkUn9Le8jhLW/f4Cg8RYMziqSCnUpF
PCkBkSQAtSFQto5EO/R7n+zNt8xCYLCEQERDMAQCQTMj3DR8fWwXnRsLWrAzwu+fli4HFQgD6IbC
zRy2z73LIsZVn5jHMw/VvSU1H9ZU2Qy80aNPMIOgaZWFDCQzOMRz+NqWK5Ugao2mjLs5PjaA1cE7
pxRyv7KkkBTzjVQ6RVbB03Wg0hgMpXzZcu+i756Mopkc5f333bkVzHOSMOVUF8N1SJkMeRyul8a0
DpghNQbg1kRjoqR+cUE7IZR9QRyuhrmhAUt66KoYBKQupwJiVPm3PKyDIC0QZ247uZsbpQusJvIv
tp98kd2TrZLc72+oMytYdcUSle+7Srtsw8YzJ81tSmB0Z4KJxn5yb0BrsFVQIbq2qzKnBUPxPYpD
OIUPbR02wAwzmnP4eFFVrs9JNC6lExXccn1DW7PU1MYEYyN2wIfyS+B4EhzRWwc3ZDXgCWsow99p
XJh8ScBvLg9N0FcOkqzaWpqhXC/8auhiOraVMPz+lyUdG3OKaLn9YryIfdUHPf8hKDPygofQIy/q
zvGCNtQN0qzz2/7h9tA4Xj2uBivu1StuLGgPl9aR3Ld7bDBWcJw/Lv7jq+WwRSvGX5Z37n4UHMAD
s5m6fZIZRi54r1jfzF4kh3ClBwjQ9Gt+VGAxcjn70VEOB6RB+RER7Itaayh2M3Nsp9Uom9SlnNXe
cr/JC0CIUba0Ru7Pq4Gq8QGDJAAozGb/y5nI+aYH2vwbHMppYoCPlmsu21Mkme3/ScFZWdY0xKVG
vjVXREQmRzNF8wXUjjv5b3dLdF+jW/9zm+lzdJvGGfgMF7KsfhLDED/7Co4ESPfAyiA7WbJvc2Y6
TEH4Ougz8foRT784nVyYNC6HAU5pkkGwuTrGQBXORDrPPcbejC/Dkwc15LgGw9HImhjAu1ZJb4Mp
Tbnra+siwWzVyEdWKubi1GisMkgo2KFwrJRcercWnHV/JF1BsBQNQKvjlzOgWoX/ZldNWg5SNBXp
UvlHpVnxgDs3t4WDi/7LBnvkrsOIfUK6YLrUU+v6HEw17y5Hw273976KiYwZLpDzyB0QUqq940Ef
qzj9LzEbJzD01NQOlcp8mkC/Lar//GNzUz4M/b0eatFT2m9HbelMBnfu4uInU1Kkd9zO2NkGVLwS
A+YgdhWp1W97+rXEAmIja2VQDs1xiQM4O7jwP5rUWlyEdJDO/L93IINScALBiGAVn8jKf3eGiQbY
N5CwTnLRe9XiA/OaUBDby5Iz4sClir7H1U53gZm5IXlwzgEWKzP/OsVcwViCEBov5GUICvKWyw5j
QQ1RKMeigbFmC6BgWm2xiFlXDstBqn25QydGVUlZBy5OKKm5GXC7aZ9oKanGnoPmifUafsOMsWge
GikOybQAwzrAqPWY8AGHkBUAGk9uDD20/CxVywEw5+zh2iyC+w/6+XWIHMoQHiokvHRjbuZHvN0Z
rgmsbxibseeBV97WKPwYykmYXkwX7EkggO8AkSiWraV6tVgxlsFRDwzwVQZqjxinICuhZk6bwN46
91618KZ7Q4agr21830y0SV4oHCIqDTpq+JzXdCOAAZOBJD0B8F8q4gyFf8ObyLXRFkREuBITQ2Oy
7/Nt6PBlKQjCL0BehMfRzV5BFzq93qPpDaAogLsuLKBkRcCCRu3h+drB2LK3R3UdWh8UJIRKNLR1
mKX2R7YDI7RGNaQMW/tpExkGLLJ0PQ93nSgWGIBMwgKRegYVgr9ldZ0XZyRw0tFHUuWpJiahxFkq
WXzi5SdMBxdA4JcaXuaPqhz7neTP0CPn4uglp9jDpxqDSmiSUq6dOVZfiktTh/al89sDqK6Lt0F7
L6mojKw16KQ4J2FkGFbpMq5WXiTi6yJwgS6Kb8jY/puTurLknELi9QTLOFodirVlEDznqnCIA3g8
QMAoNQGkMklyjFBoQvHpWS3KLn8pYRe7RMPfDqI8sNVCy+OSyr7UWQJ49qaYUEX5gxMGkN3VmOF3
hT98XjuTavKb16MFn6w1/jK62jWtJn0TnfBZOCLpt5qEbC+Vmf9JWfUuYV+hMoN4PSk7pL8yZnAZ
fQ0Kj5CGKiIqqKSW6rsGSaPXoJJwgk04XxiU9a02B81CbM+tyATNFKisSRslYCtxkNxwr4U3I75S
x8vrsHQJ2Gigib0uQPity1SaadBEq9Y+Q+yU0ebgtnSjj2YvMLb/bceDiHVr4vSUH0U9vX/zsQTP
c0mRbseVOx2B6kAgRGptnbN+kaleCpx+aNAgJIaGMoZavcbX1hEYr4Nh3FkOD+QdWLdGicWpIVjW
UXdpVhrfxq3yb/3/JXhZYCuXOc39kVDf3C9T5eFoYZFe82TgafrI/vtpMuQQhO0g2uDsSrM6qUJb
L8t9ZE6DrKHA+6Dku2OC1NRlmttCsut3C+uHQRmjAIxU839mHe6mWBz3oPr/7jHkR40gCYIHyD8D
pGAC8VI1C+n5L9X40FUrQOPaLUfbJTh28Vo/k88Ev/zVYKUoPlZ4rHobwOodQxBBwawu9almyLcZ
wn1bUIhckXJX+tnRi+w17O3WNqFynXV6NvJRWqBuPQpcB06PTeYD/R4dnOQL/6HOn8U9J6Ox086z
/HuTyl1/jWIx2Z6fZvKBtakf4K1lWjWBymnO88/0EHB7C7YQ5TtvB8yQJjwO9wyZGTHcnMuVJ9st
kIgb0ylKvHQ9oCsdZOSxAs9FtsoGwq/hGX4GbT4UoJrwOQbGodMn3lw6c3sDs2FLwnMYBxdu0SUV
iH8GD23WtWxkR1dhwUVHYj+QrXL9YmO6dEQc3CkYYSzY2IoSlV9283zKwaT40FFBSDtqedNh9yrz
czBcYBxSP9xNt4o3O4ZJlEr0rSqaByxzpYpslo0N69ZFaFhPNpLWPME+aGAKxrFJp6Txs/VaWvTM
bF1fGL36VB5QzAgLCO+xKYAgp2/7pbhFYCYzNs/ZehK18s70xgqEcoZd9xzTXSokVFi0HnAXP3KT
sQIxl38wW5FE43aXjbhvcffGVrTMZV78VrSuxoeXus128UzDoMi64E1SOqDDmhr5zd8i4gw9iWTr
ulA/tF6xklgq/rm9NesvMqkdWezKvOxb3Z+obcQih25C02S0PcVwmCSDBhLLMJNPGFoF8OdpnaKH
VZkpDqHOLndjfKeaZYfJSj4UAaDCn9WNp7tLJ/H8UseT2nPRa0zWlnHL07giRdViks7KcKiIaaqC
/MyMq6Ikbi1WiBbB+j7aAP7TMTF+so7zboO4HGGRyg8/xTggU0SD1Kbu7sLH8PepKv5JQmVewwMt
/I89gB8n1XImxKm9311KvXdMchXdg+wSyETOSEA/lRibsHX+P4tfYRzwzLOFlt4La6Yt15g9vSBQ
W1WFYoaEKhuyfHbuMss2usqh0P1VajAVdgC2sGQeNJzf+vXac5El6wGlFMtSVFlDO/Ev9dYoXV7o
8iXtrdqXDTKIeF8jwH6qra8V4c9EVLGDG90QGQftW+Mrn2EFGILO+oc8Je57mRxaEcLNyln8qQ9t
pP/47zcLLc0A1NX1t5mJj5+KH449ucM2ppQ7pWkrlz6wvbRcq8Wa5I5EqovGPaJGAwI8w2otkw+r
3eyNgPCrk40e6gXSQDYTJYSRNo0AEPX3auWaiMzo0crUJO6c90Euepx0rThxinw+4kAQ7d9OwRng
0+JNj56PXMA8ou3Zo9BNNvh2YaDhNOgQn0sUDc4NpqLXGy23OYYblM9UWiu3oA3tZ5Hhu/uINMGA
8nH4BYSOJM3qD3mcVpJB9cwnvT0kUzU+tDEXKH6nsL8rNlS0AyaLKB0hG0uVlQlelD6czZk41YI8
EzIIN/qwVjiLehKEl+PvnBFlb2irVJv6W1dDIKK8lKia0CVEn+iFDHSPSOphuJiphjQeEyiq3OOO
NAZviRtW9Nb2tGq8g/CtTZde9Wlz5gti4bdTjiH9SB+yaf+HW8uc3L3owk242EwvczaqX6dWf8/B
wgeHr7J62EALNu6+1mPfe+/eqvoZ0b98Q1kx0I1ZAB8TeSUzf8AHoT1y4vTvKv7yxP/dCqybxgOD
FBToOvfLjI6LsFgjQq6egad8T9jHWmluBWQpcLa9o9qHTyDUsOq/KfRGd0LUfAxLwQl+Mhpo46oM
A7RfnyBTuySskBCojYH+Ek5bb2sCqB8+kHNuw/zB108Lppahcwznwn61WhevEdfEQlHCyvgratDd
0dkVWy8xYaVLiU4fFpryj3rMryRlwjHU4oeAT7jYl20yWdwufJWXQknj7ept+q+pLdP1BfamNCFK
TfzfyEhBzn0Ba8WLn7y3DQjLvqbAykYve31Bm55SvklGL1LnQcu7r+A3X5f9CCtT9CPgB0mqklvB
apRwMeMl/H95WRabtc6w91O+/iDNbSYfly/VmoYmwxLOh3uYAI3eSskEFAtxF1tjYLifA6Yubs60
GUXv7D9qeEdRyCt21ddY9gmmy6r5we0ELSy6zD9aOSSaclRJh5wRzRNKRWGW7rC1o0wJXc5yEwUw
8guMCxnqEMEbfhs3oQgCLBx/oIrVt69P1lE4Z/YGNWjc2bLIJCOxvHn3T3rsNmKmn54c2Y5PESYb
gxLPDi0VGa41g63rx6Ww995fj569giU41zdCRw1wPR5/FJ/ScVNe2fTBP8KnlcWb6fRb43aMnHfF
T53GSg6c03Qt50LGQfdYvpcSLvYsmO9Z6RtFSHGnJXhgqU1BRHmQ7oAnIeZCYWqkDYY9n3lk6vMI
1z/Wnb+PkdzIM5eoTlL5XDcaLnug1qP+lMeR1ddXxAhgJAEbOwK42ec5MZOq78ISPFBjJFzLtPLg
srNnOLK7NBDqtETXiRgW9QOL5F1hiGDlQ7RmbW2d7BkzhVYt0xQ2tZmefr2vPylHLvaBjfkou/a3
QTVd2cjY2rzFyhpMnWSsTocCARHwld+MQPE1hUCthfzbG8+eIlPvuBj3rOMl4qFNDOiLtexUj8PD
9rxcEug6f9df9Quc3eSrFlEHlVjbRfqIgS++oGqy4Ds+XzO4YU6WeK4FXQYwY5vUkT26Lr2QYj8h
E0SUN6hoXtjugPu5azYdqhdpsGO55vypW22DPjZ42u2JRMFeUO4Sd9vTM3vGsAoSLYtfYTUy8T1d
y32gUEtJKUpLxauK5yJmKvLSr7SugVngOBd9Lt3sw2mHFRM2rdOGmqH1I3cEouknDSmjp1qe94b+
yYfdEFDtlnC7n4R/R/O8eRTxW6zF4259DDQ7ypWiLI0pBIfOEGKe6dqk9basODuF4TkHIXlN9yR1
k1L81dzJP4XL1+hk+ZDjWCG/JcN4k8fkMqeRxAzmSZRsN5znVd8RIj8STZNBnwaG6kdL8Zl9cqML
1xp6Vxl0OZXx6v2zbzC+BKoDxY3L5ibnmbT+j3IbEpYE39SGuTdjxNz95lhrODNEpAQQ+J4eDTLI
Ee596iCv0COO6rXYmQvvxU5e/ZdiXtBlcwWLH4hK18Vnp1C1TKGUALxYk12ri+CGrputTbnWmxNe
/eOAtpcs3smYGtxADjHeGO8TIbNrqqqmAexJ0cuyJjSOUy6UMyRXiGEX+EQX9zO42j77QaE+tF+S
g+lh+Z6N559+pElTLsFXXm4NEO7IUu8L29ideC3dCJAj/Oilc6g+cavuelGx/IQaPcUnED88EpNl
3MTX+I+OLSmfa0r+ERE8YvF8BXpXlF9Ij7eOsP/7z0k2kjW4Xjjjp3kUa7UDYvPsz+/1PyCV+BUA
s6gpxntXH0O1trfceXmFt7fDn0NoVlaC3Bjs6bRpGdC1yAqOHPmm9mhy7mqloKypeT5q/FyvqG24
3LsNhfJKQid2kWSsDJPy76Yoq0lZnhD//ourmCU0EcivF6SOqVULk0Ha0w+2nWmvMvJJMrT6HsZe
ZrmFHgzlx0Gw1Hrnj8Krz41ZXgyhjZd+9qfIYeS/cxnyUk6OANIMJJcAIRhnfChVtD0M7ESnYHrA
5Xkzl9O1pB6tG0qOqlQ8WhH23ulcOe59xfbWri3FIHZh4nAqjoJauNVZxpvJW6OUiEsc5nJugwlb
dqD/CDI9vy6Bckh4t6TRX5XPTkV5JeExGjTEnKR8WyUwsmyTLPx6HnhbSQfwsJxNJixMaY3x4uIq
jpo7UcpRnD4B6Kuun+KxMUalOAFY/eF5YOwVelz+1dCuUOxbzF3VrLZik3wej3oFDjmc0+pjy7J+
U+/c9BzqH6eRzxK+Pl5iLtLSVVgYxeBicopzT+FIb4pjTKNIhH2Nmh8TH171YEzYY7nUy+AyovEe
TEy9AFw7IOj+CjjT70owsV/avDI4W1c875eEUkOzqN+kVxFve4DOk/eeAdRil8XOkVtLyQTFMZK1
36b6mk7WKPvL7lHRPpIFsbXNtu0/t43NGZgzQ3tvMGGOP37yWfwsBvQJ+IoSOENMyrClxUuhdQQQ
8G5IyrQilPRj72k8WuI9eHEWO4wxefoKd9XHFA8pnqqMtRo6NWc9txEti3BWnmQlRmmYcjNkoAUD
twYfubodrkel273Kd2Tq2UWSvOy1fLzbOPPxyAzCcEYiAAK0q8Ru5uGNijeHhCdlPCcN/fQiSVAN
TlDN2WrfK/FOiiaTvcSlLI3wNJPw2yZApkQ0+IY/QXUn3RYJrm+tSRXn/rDj+2tGRwG1Pt13ohjg
Tzc0i5oU2lPF5itIdiLKCsG3CorVcIR0RQJxHPoAFN9k1odWa8JKIgbcIbUZDszrrN1ua1a7Qlvf
cyOp8umSOHALwweeZV0DoYOkBnBeeFz2N+40DIgpeLwyNHsz4jmC8ehKKVkg/Uqc4WfyDgRZOP4v
5/Cxr+Q4R0mkG6N+/rlb5ffjUs8FYMS3bqJ7fV7YSB3mH9qiz8BdWYbZRampH83AcXi0jb9dggNI
ZJ5a5Hkj3xqqVrxuAJL7Ih/q6eZCunbbMh69bJrS/IsZ4Zqq55JNgqCBX9D72/+f8L4Aqc94LBEO
npg9FI9qqQpIBVtpwVkbr7scfKxt/EdHEG1rif0yL9uCtr8HOVMOhWi5mo8yM/pMwGlVleDm1rTR
a4JGNvuND1xH1JnN2cL48kEWIedl3iCJ3FAWE1skVK/BBuIuMIVvllpJti8ns/4H+TpYHA5KzxEl
ejb7CKCpoOdp+xICQQ7lNl+dj8WTyZ5ko2iiEJ90kjF1+HjEyrAd8DdC3tA4Ta+XJErcVRnGhEeo
1RrseabcuMyyt1WM1YKThfer4enqBDayBe6i3Seiwhu6P59/xTDWayPhVAt3Gf8oGjWq8t08QAn/
DX9nQPOmxmoT27aTZ7HvX+SBHN3S7LUKEt50OJfCGQtR6krVkTNAQrKufVwyyvgLa2lzFxZPL27G
cIJWEXmAsw+BjcKjbyAc7sAwR7imslbKo9be6s0C4UGH/ubIPCowCbKL0cHKMV6heDuWe5DdpwNw
zzgLtGT1rvOk7iRNpRqSG8indPAjFNlGM8A5+hYyjgg9C52F5fsMH07Re7wpqBmQRSuqFZz2nrnE
oLSEjh2jvxL7nGLSpJH6mWRZY88xHRgRmu+md5HawXZnMh27w1BApV673O4dwnEFqKmVOn7mHm3R
TSCbfH/o+yywFGRLRYl/MIfhk+dvM9JVCMdFO4u28XlcsjLgSOUCZu4L4+7plaYLhxMDd3bfz9me
5pe+HhUqg5EST+l8ggmyEOHjYhAKEkIqpq3yCBEcMZ1gr48WPm7Lxfhdc9sq9fL/Pmq2n6jFCZWE
WFBo34q1rtoXnKYL6pDt/wvo75+M1Sxxg9dJmu29D5RR+B/xcDsNzBHm7Q0Xkq76HjEuh4b3vUSn
q+gEcvveuM5ypI+a4cwGuttUCJTX8aKif0Ghz0c2RwyAQQRqC444tI3kh9OIGYCBWiXQFftkW1Du
SPGlLnkQfJ9XF52IW/xFo+8rNoOAWEMS170GEMDq3gvlwFxZ2DTKvbNsriU5nqC14Jhi9XvOWn6x
nvtmipWH7NxvNtw8eQeawOfYl6NQeJ5qRvaFqlQOMzxZ0tl/ufsuraGONurinXKka+KqjLrG1/LW
obpFgN1n21pKROvnEG/maON1B0FaCoBwCucy7GmT/FYpbYibppuETK1dVDH9lZGwtSRhO5nunGLl
fN0I8yHASu2auVxFSbeqtdKW0lb96E+wAUvUO2JBxxaCuUefmbPg4dsTpp6QCeL6oE8fuFmpKkZd
z/s9DyqIIIx0zswRwIlZ7a++rm5p1NyVOi95U9A7DCztLZGLUKcdqij+tCzYsyLmDoJDkOaQnNIt
JnIomxixhxrbvK+wj+5jFhRpZaZwZ/h6jqQ/yX0Cn4Zwt8B54eXD24yW86Q3ew0twZZFpoN+kS5S
ELlUoZ9bIRxKIUYnY9DP02gHn1KApBf/NjBzpAHMRyOwUvBF4mx+FczeBsUmk5Kwwv2Qr+CCkHYJ
qshGgMEc6cLdh2MaA/4FCvZJT9lSP3k4oyEsoEZo9i1kkDfVNRVHOtEq7DZRQDltypCYP3Y0/7Ki
myYfh/0xCTo5q91rWhm4p3MeChY8Q5AznbZybBkI69jslfWi+p2MnRR3wHb+qD59t/uAORDJ3m9z
x4/kY57jZDwqgERnRziHSkTinRrEl4Z9bSlRHe7cVwcTTCzoeurGOSr9wnQq70O22E7MsuScM8Yd
4lzXCHqpkaDrVZQPIpZW18JsVL8A/tF+anoXAExhLnqyA9vA+EstJ2n30T/yG/sLjImPZ+h1G01E
wihAtZoZZzWgkBU4Ksqp5AOcrK9Iy90h4mzLGYtEXJyOxmxmzNelWGa/tTVISOiJjL1sz664/5+2
NqxQq4msF+jgEsk3wgCfHVhcIhsq0il4ECuzJ1+XHF7m3W0lcfVN1D3S58PY+DLi93QcOcgtJ96E
rKVw/T722NCplrJMosVZKJru87NaQ8Uha11OtZOiDc2UxW3jyOpQW3jmhq7PDAnLX+aBOQ9jrDwe
YBCPgcGtvVI5Jkyx6WoNsts9qS0T+i8dCqQpmFDIiDUugMRc5Kelm2rqxgPXo2kTgtTXJ2pubLAK
MWzAwXZ/+TNg+MT06RMMwKccSXsJcjQEOoGePi+cTPBlJYPeKTugN7h/pSStjSSdLIXnj89tfsfb
asnmRqGk8+0bdSPOoR9QvphYWvD2bT+uFZDA7M3RnjXqrMS4gtwEiKCmgNHoxAGgcoM7ee8W4l6j
HANBQT2QJCYL87F1zAnpgWqSJecp5QadQjPpbyKK0s7tDEyeC9Z0f1C5CnWagaF69kuNrZDyUR91
vDBP5yD91RqUPp9lc21CyhaaMac5gq68iZ2myrYSB6ZFl13d9gk9d8BhmeMRpemhOBVPOBJ6tumz
r5NolzWDKyVpalf6sbMWuWtevEL7jJvGhER5EKwAhKs3/8tW3KaBVn130MUTTvbW+6S5W4/wG6N6
npL0cKBowW6x5jWeegXJf/+6/EcO7dzmJkCqUtEjjeC/AlpotBZnW4EQFuBoitr8PtzqAXkuKqDE
ZwrehJalL5m6ixxpVP6Mt0tXY6KEqJxta5uV2TX2ilQfqSmQ9Ub3S7tt4vMFC+BepgnKbqjOIEIr
n8PFr7YHPcPdHw3Ie/Z2BcBE0VPeoswDRjk1ZGS0iAZ3Ggegd1SMLA5eKgWO2hzWqDhey1GB4u3R
AlPsq69bRemEp8+bjITneqYlVFw6yxYu9Tqmi1+ggkqqST4IXnv2AcbMqgEgg1wsUmXkVIPd3XxQ
HbclfhU7A9bs7O6xobdk/bt+zG8cSnTBbo8JXRdlaaOxxbZWCP52YWQHKHRfNamEYEr8r62StScy
yN68eFg5q0Tggxf/6vUr9RiP/KHTRhuImSn5uQFCwzaPk8k/mJtGtc9zY+7ztC++9Za2MOpQXvh8
xEjPYlJe3GcJFz7B/8p2Spu9W4YpJCVjo98zRiTZqqbK3lbCsim8RbKgPbBxZC0TX7+gWUMRaVRO
Ftvt0X0hu7Xtx69Xn/B5APmdenSkyCQmuMaYxRAH19M8x381Vi+j4MAzEgN2xo99T5mDP+vLMz+5
mbkMq2Rsp7M02tgRsxOWG2p2ddaVZdv7Jiww1TcDmA9CTX4ptsr1ctihMDuXouTsnDHMFu09PQzK
WQfTtFudeSIKgPhhmuhZkupcAz0kIDeQ4M8+144lX6GqqX04dqeo1d6+Enrc78jX8gFdWhqcha71
tFCIfjcuBUn/kl4RuNds/lMx2gR9rC52j2Q7sUBL0CE6tZrq5ie2DwrBwzVNoJotzvH19bWCiO9D
t2XzWa4fuYrd16IzkeyIuoNoCBYxbUSmIMBwYFtLjLQtrwvfLac0hm4sWk3YjGgCwNtkUV65Gayp
intMNLY7Qs8zkaC7Gfw7wErkxj5W7zpvUXYeKsnJLSIGaPeyGWi1FkSdLR1fllMT91UQT807XrRS
mJaR6h8pDZhXX43WWHZ11h9dmGlrMJKiy5Oe7wW3Q/VcP622I+6hPN1ZfCwBJMnREyD8XwAlB3s0
fz7bA+mkhTJii4IKtD8ePghdCdlA7yjeerWFOkiQW3rCXindrUc16T4thmbxH8mSq7gy7eg8D6/F
mQ4QAPZGm8a2rWHcmqbFuFBBJx1ZxvzcxXvgPIIeKYNNaCmHrNf1fjiIYQscpRd4Z2ejYFt8sYYy
sPY7p4ByOi10wgmqlgZZt5bTjT6TG36i3fveMJihIH/kZqQIqVGbSw+08RVHypyyVLjhgq/WM7ET
nmJUu/wEXXclB7YCI4DHJnDLA/znXZ/pEf/VwsZFY4e1M7yW3EPCg+ca2uciIbX1Ac9xsEq5swoW
5NMrSpryOXUFjOY5asW0z+Hv7xil8Vu/bkaKbUR68c47dObTrkzHOhmgNwyn64UczXLdDSIUWGMa
qY3a1F6b9J+k/Ys0/+oWYixw69FA3PGLVSd/SUIAkN91JQsUro3HQa1/jnGkQCtWridrs70gze5/
JDT58vsqd+3Zctg6pLlDVXOi4UwZxRi1sMD8Ve0Asktl7SauCCYV2EOD6eZLcaPs8Zd5jR82EGlZ
BuXzZLJUQl6z6f1s6fnbU8xV+MHoNRnDlhzZPTMyKFajZUKQzFeB+Z3QSmC8vx+iEgzsNHXb5VRZ
UVlIzstLevBCE9OnunnrZajP9m3Nv/IlFRd4WugioFJLFqMBWaQ+1S5F0dL8CxdnM4y7b7NAvlQL
xY4MGkImdpcpSvg3IBglSCi0OMVT/9Uxw0X4OzbLkYW1ewt70oeHHcbtuHM08yNRu9B7Gi1vXqQ9
Pr8fytQJkCjWk9dzPLGoKy2/poi23y5NABb2vAimcr+F8GL6Nm7dpfj8402BwDBrVOeWtRs1yLDt
uqBjHUNw5D4Q9Q/Il+PwG3cFtfcosoDGnsMT7LLMLkOaY82s22KHDXBIjYh9moj6dMpOCNeDbTdh
wJ8FQv0KNYcQNpp7Y9gD6/80acuMjkCMtV6MBsJr2SAF6P1I+AdTdnAZjwc2w+H1k6LFSrHt7w2C
bUd7qE7nFRTXuVaDcflIlBFJiDqq8KrdYLDRc0OfAgUN5TU1iecaCA6ylB5+Z8NmC66KlGpghrN+
3GY9IxMvq/oEb36/HqKqElcJc5I9lYVhK1y/aHjAtcGvm9OzfW8mr8hdh42eck9nYoQ1BolIBAe7
UMC2AOUGPO+uJAvygsM+7n185Loj3ZZf/1vdPQdlgJVgGxy2LzqPjw9GW1cFLf/r45Q601kf3FuD
GsF/gKZjCUo2QZPF/Ew1N4C393kOl97C8l4eag+B5argNaenKRhGORWyMMncCIXVlXZc5Hw9CJtz
/zp3m+Zvi5QWGmLCcIcXL2gzFbxdT5TU/YhKluuF6v5eEZjYPAHioQrKLg8KTYZQOcyte8evpcfd
R3pFgGxWgdGjW1eh711munfnPw5D+jB/eB2dFHY7JlfDMI+ayz1uKuUNqRezWsiGgck963MZ2F5W
i1LWmKIxHA0tZEdDJgS83t8tOcxR+fQGtwzbjyAL5YmkMAficZICQiDhZwGxUPrJbrLJ6DpBmv25
jA0iu4FfIlpm1wcuLTUUbflEJGJs+45EydWDU+UixMAGL9zw7nFNlGqHbRUxqSOVqAoXQy4LWGPR
nNou9IShhnJSXES7BJtGbh3kNR10YW5NWWTrh7pLcr5Sw0J8eLAJ5cx3HMeBU7LX5XalOLiDUqP+
9+nXLzKmsAo5DecCqR0HmI1T3GKUmIR+vhz0GgUBu+IVmtwc05RtVBtkQHuSf2WSJdX7bZJtoIPH
2B9XgzyvQXtTJLtnwzgbX0lRpxacKgUp2tFjXW5hiqjVXPXFDhzfEr47eNiDbANzgyrO1A7c5h/x
cj+84tTArofsnMZciodiJXDNEh6jDgWZaQxjkmWm9MAkW+9oOLEGTWBJDpH/fDruYe4ySEhQReJD
IXkojTdmk0Vl7sQn0Yd6qFjtMPinSIW9HdeW8HZJu53GWrJxF2OyECQ2OHbmJlswjwihDOhrSJju
Ujz5fk0otTjPjlYO8QIAYCtPlIHVi4IUPjmJ82ojChqXsCNStEFJGgMyI0CU0nlb+6U6C/WOOt7N
/EseRLP1/07/Bh35vmAMme5nn7cWYBWEvJsWeMBES/QRvYlIIhLB0ZUmotj1WPl6hTK2l+hdSONS
4qcQ3b3GMOhIXj82Z5p0Pjq5p+qYwogqFMSugs/7Vb6JsuSmbUvF3PoqTBx4J1XpEDxZbx7iJDkC
TOb52WW8gpbSEbZ6/t/frf/sFrsfjed4ptbOo767cP4rQqtcylkBQSdGPOVh65DU1wiEmcToYAfa
gzkqnYcHQueze2KKr4VclvFru1w62iZeQJLjf0wmSkutfJJ3vwFgUcW4dklsJlRQhiRlcHyHkrrX
urBkq/6LXWDUyigpRRc1Oz8E+InrfKMIElfdrUNr1E77+CCmxdgaHrsXf2EU1O2QrWxjpyv69z+q
356wdDKy2YnbhucpGxi1fbbPAGk2Ydq0JyQL7KmKTjPR5Nk9XJOhgqxkd1A8g8qgpou80f3rJLf3
efQenVyZ40brjSBy0lmvYQUF65Qhs827gCl6PRA9MnbAGKiAJt87F0dar7Z45sk50RNIQu2WtcJX
sH01mI6wmifJz7C3LCbtqX6+cP2SjQYQyM3IFlJSEMii4WzGmAGL1ioY7O0lbSIXJsv+MA8O++CR
6scH6i2UXR5lYtibVsXOn7PdG4h8DuUSX16INvP90mKDO0YwviDDGbatGpouNIjHWuH2jj0b9K+x
BSlthFIljFzePeAHZwjg7Dz4SaDMvSPPMgg7dtNGUnJIjcyhVe7ALY0r6hrs4iLsBP0VXJXhLl1k
jtovGGvPtB/Ltk3L1qBqlVUn5uP4myz2/MHPqkbCziQexjubBCLOUNWSovQgRe8npFvbHRLUuJ/n
+RcDNcObJQBDD9f5NXyl13Nut5YmEyVEzpv4tkaaQToqfNpVw0MjF2ZD/0iv6IlL7wdx50zxzOgK
UcSQWYp5VX3olgVrH4U7lHc0vnMqNjOdJW4SEfyfnnXiO0JCHueCJhXMYte4/ov5A0YxApSpQ6yG
P2q54D2o1jBC5VFiMHERKpbmqEbMIaDn2/tOHewLEFXg4Anl5J/fO6+CgT60EJnlq4EjUKEsWs1N
wEmDTVcta8515LvnUvnuvQhalefyEbR0AfQFfz+Z0uzJlB9V/33mL3Ws2Xus1cZF17cVyk0cDHKe
kVRQOiCV4fgI8pFZDhUgrqd7/Z8ilV7QK67aKq7g/jBR4fjkKBvsv1i3vz81s3M7nCEF9ZUVHRF1
1H5AXNHg9AEgZG1yoceoU02smEAmyVW/mn6mq/XIif07MWUsFJVMfN0RxR5bAnu/7xct9xvw4JQw
jLxajsMWio5Xub7kohyb2uqzWrzSpp+fRzUG1zisWNX1qY8+Yq7fqAmxCfG2rsgia/5gFpiofB7G
sX6o5g8hCxIoAF3tNq+kcj7aPD+VDXwwp3dTbN3/9/2w1xmBjyYZz4uIR4gDJnmi8i0rkYMD3roy
ApvesCCGoDs6SjrzDnhmgsuoLvL8o7xV8ZwrGV9SkJ5xVesOqCjbV/9qlh7yCfy5S5sl2PUTf/VD
/1rFnjDZfRIQOOg/SuDLZTTff/D/FAlFtN63EAGQWJJph3SExNtMvJyLwrHTZSFNfTYDzobCJXYL
yW0wiqBPYtKexbJ61pPsGbY46t1ZEbnojSbad7YEufsdENJA5hD8mvPQU3zD6i0BHsiuXP0WFPPM
82YVPsZyfdTotiQIn0jl436KEjJ9OPjMQsGmig6qpd7zy+d96J4nGxe986GX/LDtoycu//FDIhPN
9vXAf6jg2j8CIpW58HD3JGOJJdcN9ke7u9auv+cjcGnFjW2stcnIlBrX3dCpYC05GJWtY9VWGOZH
LF1rtWv324pvB8krfCqQXclFm5/BirBwr+LfiP4kTI9nQJQ37paZBYnSWiqRZJsLuh3wAiAP/t4L
iYGnVj2EP45nPxxyYU99FvPtSkvkIC3c1ifZvOcGe4+0vv7KZ+P9WxFxjLQBZm1f8Fy+z2saeRSp
hxxRyLmsKkK1QshV3TbTxBsa8VIdl+pkrHPm07WbWDtS80Rp09mEwECMiwzdZCpilCQMOQSkxVIt
4PQKi9tQfwrrDsMVpvbyfhfyC/oU9T9EibwehOHvj9LikvLuOFSeGTbPHeaywBWEt6xa+Tgv+h+b
RciR7BSEu+DJpM8c/SEjnZnw8JZfAREJBu79tBLCDiwn4n3bm6zYvBxX1XZqlqL0iRRND7kYu0Iu
Kk85TI4fwveXTQCSIc5R2rLq7yWTO78utGy87iQ/HAjXH+EDhg/Ubyj4dUxX7wu4Y5BhmnfpLW6V
jKNPo/+KiOozFOjjSbNYoFj6m4kdpkhEQ16OTl09qqARAR/2WuB5SovL0Jpc5vdh67KmiGJonpEC
MwqVRT179jtS9t4JG1nPpBg8IoHqK2KW0FQKIyZy+0AyW+5xvX19V3iyLRkzMl3p1vX7Z+Ou1lyZ
4k0AVHm9uaEMe4HBxLXampXqtCs4y5hArDgixyJVLAAQ+czr1kpRfMS9yQlDy1I4o7GuIP63B0Aq
xJHo5NXblTux/Fe9HgnO+1Y6MBjupin9J7NT5aJhsYWBUC5WCTh7Lf8XCmsxPNI8ZmCSQKOPxSfO
NlLATDF6pbDrZuZAgxyEfxshy30xlY5ZxL++DbO0ZEJRQe0RvCM7P2V1Fcml+9EgNawN9r18/XcH
Y0vDlxCl2KiPtooBJUe7ThahAugz/YvyoirvbNF2/XlPk82XGJys5fGxpbxvjYPy9a/ZAtV7kxV6
MMmXFA9Zsvu0IBIQaZBWWjK7d+8StU8vssBBRKaMPewBzKA+iyyt3V/GjxdBuYqK1SOLkfuF6MsQ
y6ZQIwO+czzO2KQH9VNXSUhiag+ammwCWxqrrxTf5mk/CVyGFnoyvMIpC93zrt4oBQegEFUIsy4M
QJpL8Cppijre8Dt8gNDZZOcykW76Xjj0hybVwyBWYjivCf39oPlZe1ulh9d/oafPWs6xn9jeuQSO
JJLhBttfS3TRWVvfjyITqtpUyMUwBVtWCW/RASxUecaoDFKZ5dVSE/Qcub7nG+u0xoUZXOKWOgJQ
ZZoRfRtLm0mv7c3YyqaFR6SnRdMuInVrH9gFGKgU1/vgXvBn6sUB3fVc5RFJ0I/67LSogwqTwYvJ
egDNofIQZ1A4l5VB2T7nYxQwvr95Xo6kPRxOuiI6cODM8xKJd6oLeOzSdw/hsc33pirub68Kqg7a
5tqmQSFQfdMtlK5sWS99FH9QJi5MZ6U/2TI4KDR76rHvECOu6GbtcwecOAYEMdqt3VNGKw2H0zCh
wdkyNKOrN7AzjGDPcpKw8uRjPCcGhBJdVzaryGhMY2zRzQIft8vz9cMszqTCcq4ndupC1b5igABL
SzFVEePX2fOikoczSfJnEFA3wOjVhW2Q5/AtDTx1yzHs2Nl+UqlAAtmcj7ClpeDvaPJrMorp3GKz
ms2qt3qI/SDPWDGJ+Jm8K1V5rjVT2Dmz3QMyAgrQeULH/xnrhRvEX7SsgdV+1oWpQlgys3jeIwaU
w0DI9iRXXo4/NIVXJUDgHHz8GI9n/HgZ6WTNMLRl/5DMvrZQ1z2lpAKswgZrIELZjU9HewYuxrfB
//8h9N6q7IjtttB5uP9vnZjEM0Zv0sykxZrAVXmQlTpNrILF8gpo6i5eLOdv50/XWcQJOpE5maUW
myXBek7kUGsTNyizb4buY4bBfTLUNR93go9p0Ty//OoHH+wXXjUPUxaSLCp9nOnlu4OxA3eUToiy
Vd4tCd7nClUS5+ZNrSEBp78e/DfptpDieXxmEwDWb6QKdt53+rLrepHkObAVmmPdeRdPORiZjEP+
WKsTrpetACoKheNZShDHkut7zrh+7SbK+OyZsF2yBytahbVOne3U3VJNsuE/FOA4ks7O/6nGzuXF
+LW7SSSsMAZELFz7lZpJwZi9eqLrOiMzjRy5qT+hZWXy1PZI4pdyH6NcebwU/+eRo/rtvrW+fUjx
1E2Sj9irIIL3pHhjB53rKWX6osurefjokrRNc5jIULzOG4Su9q9BXLoLyFjRYOiEcIy1wH0heVaI
a/p5smm9ytF5G11m3HX8d6+3BqXwkghkr2Pbbk+RNMHMjzGjpKvar+gNKxwTbfrWJo/F7hJ5XVs5
AFhZrey5nzbgRSpvCmvdPs0IEEmX5w5hyXJlXKAQ1sw50zQ4A8PCZ3Qe0WiwS1d75D4uVNIzzZvp
ONI59T4eYCSat8Eb3Jdhsh3lV21QflPzKBhaTZHY1QjpSVTTi8apHOinIyGD/k7at0OL0Q4Og0+j
xNzgF+ce2lGSMteGnAaCL+3hFS7tANVMObpybjCjkI/b4eG+RtHYxmb9N7LEbJiT9FHCkfcUSYfK
9ZkaaZAhS1+ZrS0qL7F+nu0eCVNDsbHJEhxXpGONp31C3/DT5W37IpFLhfnRnzUfIx0Hf5h6dsyC
BSjaeTs+qs7jKT2dH0vWc0iWVW+DQpIuqyhVNJbM+z8UBnKRrR+hZo7po6xkIh8YEBtDhjRbElY2
ujiqthwuM7MoYV3l3ylPd0f9qf8qhb0ysZxpFW9PIbOSgePGDrf0R0xhBqF+3lcjqxF3S1E0E08p
ypxg4ItWGja7MJ6XcqBylUx0/XavOZfo/BDPKE31hSnzQjJjvgJ0USwo6WLIU9SWSriOe0asUl35
J+rASd5nv7wz3Au3UWYzMin9bTbhZbWFGRs25f0q3EPlF3f19cM9Z6+PzgA+T3xnbnORAQhpytrN
G8dshw2bbaIItYVNat1ePfNxdrhjrlFjQ02/mpg67ICb3HR1WGTvqLZGV1lvrpMJ4ewBNM4L4/tI
pgBhgn/cFFrNceOY1KPfXmrSIOrDLNy9VJnI4xOrFA70e6PuxNVHbSXyVHDRY7fTG1RWkqq9McoX
kheySd4qP4/I5VQv4I3S0NlrOThDY3O2949Cofy+0Qt52YHFNJZQ6KyKQLRrhLyuixKuq7UBal2M
mJyeGLBnuXU/sfD01ns0QsDLqN1RquOhtEnFoRNV+MGZTU7btgUXjHs0SoSHLpnsy+AojErLJLBq
RskLmroZnp/Ji3cbUXU+ZUrrkZtOAoYqZDWJCFyxKnRustTK5UwyODghlyEIHLLLuvUJEJ/yeSMM
lNasMX5mMwFd6TyIe96RgtgEYaT9Oavi6HyRHcT0iRG+etciQQUJpL51LmJL0WPL456Zok/YLJg9
I2QQ+GJrAf7fsa7OxBT3zL99Pvd/iAz2bJx1pPrSKNOK4h00ZGHUtzRJqjcgmObcKClIDy0VDAgz
IK1yyBOFv3EJDvWuZ79p6IdDy9ME8qOTVXmgOPikWfXbZCNofOREX/Ty3+mx2knwF6opO2gxDH9H
h9wfj3ZNnJOxjZHP05nh9L546fAM6OxCV5049GE3cdfI9rsePoOv/kFScP+hyJXNMxJAe6Qp6usT
JAVn0iDJwAKWmQzGmZ+KD+wGjxwCOnMVubJ19givxfwDbxfSF1nIFW69rCy5+UnU1o9taoIRA2Mb
VhQEYA7NjQMskNWbM7glKN1LWvNoPprLrmTy1eE4k6klZdvbcKUNM6jmDmddDqyKdVDhkQEaAMHo
/jLIyh4JyEgxZ3GzigxUavXBBVgU6IHsuf3nMTPpuORva3B6U5SMrQiwumvppRuZeASdf9InSGm1
9Sze+iVYvXTuB1OnsHMvp1/32xthcOarSRlfSOLjcjqyW6+rU12Gu3WvBhQvySsaac2vpeyRWZ3+
wYjKY6u63clqiqlozU0eR06tk8W7SlA9ccBGFr5iZnQD39Lr5yaWXNjOEZQH986g3clWkBap43Bh
WVL+uKR/8zB2tx30qH6o+SCflvWafv01yJfwk62MKC+Jw7mfodxqayllr734O7tPNOfDbm2ItlyY
OT0qAL2Lvp2HOIZKG4oAxifPZEh4xrVM9l5t1FvkzZBO9Ze2NhhFF5wirzF6Ni/OWiUb+HA9s9lY
jL9Q1sLe54/nE8VMJ18uxI8kbG21RQBRcJZnNqBozPCBgVzWhf7babs9kUTLTIA3HPmUdaylIgmH
DbBxCOx+yx7jUh0ZbNnDMKq+9FR4383YsS386eD61JjK4jfKcLGqTQv4y8nNgZ4zd9Sct/+HgPOc
9pa+b7lTEtocFLETZaefJk/SyLdm2xSH3Yx+oxKSMwQSsf+WhFaYKI0/ywCH/MHoCxuNk7a0mTgP
zoj818l13Bg2QuNICjCEXRAOX4Bggphlf53w3BNngb0TvTuS+Er1VhsTA4UcwhGaoigD9quBqv/H
4Gmc777FqOvtDljvKRqJejxbuYdgaercus91yumfQBxn6npn//TPaIQZ72csO0/3I02LPKlMp8b7
WtOmB4CZVT72xA7yPihJreZ+D6LF/WtJXkATvnfndpoag+uACxKZpnuptMInbVf+YulDB8XbJKes
j90/faSTZqTPIHvBKNW/J0zlYxcBqmPS/7g+dOOhK3cVTOhGfg3NbgFmWAS75vg98rmVpt0fdlIS
t/9XT0nkeNduEF6yG27WQaSs61/Q+qyGc2aBsIdnceNfrNRKi80iKsiiLDiRfdoMotcUCvMxjbul
q+ceaXZ09qU30458casNcM7acfi9K6toIHYqOL4bm7U5fmy308HqFl0Gw73GfdiJMWNso8uoQECa
B67T0u4+h5xuRSeFQDdyWsLZDtvPX2f33Kdpm+q6FOZsFPLPhqUU0/ah3Gc9F4xYWSPQ1urjllJl
lcgoMmiH01hpoSx3tKIPZYQPwbu7vdyLG89C4dfxrMTpS8lT5kD/pkVdg+BPGUZa4HQBH9rN9M9z
RvlWRCucGSI+IJBb+hFANu/m45QNU0NXtXj6fASm44yYqJ0Z+npg7JYRtTeQABYD2CJDa+9q2YBO
yItXKhE1wYAxdrHvQF/I0fJyrPF3NfnYxPS7n/b53JQ0AtwvXDLPh5/5a7jTq3dFiAuvn0J8XdOM
rpjKBigUWeIvaitz2ZzbdO7NX0xeRwAx1xTw6LYKyPe4obQ1mXtV/8TYsAS198MEfjCnqGnHs/dK
4Ykfp6C1cKqT0xvJ2ZvvSjiZTNERvrgmorp8ZQTTLXzuPIceLrT7ohwd5qU594NebafGy7ZWMHuc
v9wpLcr0amwr/EZzOgcaFTJFp0LLtEGbouekcF3jbBmptjaDHR86LpzcVxioS03qY0+C3x05eS+C
nWxn9S5buk/QZYqgDJlz87vmf76b0P+aSiFJpeM2f3HVA5QqDNfpJjM1tD23oUedD2PlsnSncBpZ
ZDjrwsJKqFRhMbmXSvWz2kTKNhbUXCWaySvUuJjyeszoKL3FcjXiX4KGsO/qncrqDWHL3jU3cLI3
e59GLn0j/IuHoyB3DiaGTGeXXpwniwrUjE8zgX+q9i+PofJle0OH0fRRf+bpggf65DYLItoaPA3/
AevlCT9dJ2GqBKYCHMbodS3T8GiK3ddIxep876PN3JJKqM1FxxYIjmBDtsCBsyuQERzNviEAcJ+a
kVCcwNfCtp+caSzjkNIIPcNELkCOKHqFux0LHyCsupsFQXexj5fS9TfZoGf81JGweVP9TZ+b/XuX
m1G58DxKgycyk7rPVFjnHVQoUOnw0ngxLCCdcW5cML639aLl2h9ORy9FJ9bnxzw7DvZLYT43vJi/
orMwNiHlrCEg1rY8x9YV136oE3Cp4kwLCCZcfUpbhO/CDsNvV+9vB/0NdBqJQ9RIZmdDBpQFJtrr
rqpVjXhqt7uKc8PcuZTaLsFFDzTUsCZbvq0VNLtFAZmzkcn/PhiSP3FZQ8LVjyh9YVKNHBs1rsFJ
QNwVvo+dDik36SLKREytCBo5ZKJ64zI0zjLWguYHGsUUv4XFVEM0UO3lAR5lsIVorkCSkgQMO9CK
/WYmENHOwqBCOwwL7qgB+dBSuv9lrNONFpAz1hPxOHVCP6jEMV6Oe8CGQWw2n8yhOSlRmlZj3lQR
cncuwwRRnMXczaENsENA6076q8zo8jDWMAMIF8zDJmc1MNPhtR9PxCssz/iasYBrdVxRarwjpDqR
onD86z/ctLeVFEk4Q5BsFnFtvkX5IxyyX9xeFxYbmKFsj62Yb1eBpcedH1L/R/5IlklVAlvRQSRp
NLgvY35tZj/31+qUYwk3M7dzU5jKgJ8SJdiUrhuOZ6biv1e81vjESKLqBj7xlzOMpXZd7LK01nGz
NnTy5+u2E9L6GkG2Ol+4IAtUTFXCDIT+mMjw+gZzAHeTDhKarOzrpgr32UQnANxx9ppFWvqpnqEs
+05ZPl2rIVD8Wrnu38de6hGDMTqVLQ3y4kuisHBArxESD5V90lL6K47If7BOTINm5iZiH/pKKT0R
eP8xZ2sATGqkePRCp6FkS7SXx6RETNM/qdCAOUa6GZb7ToLNvWWxHVWC6+RipVCEcdNwvjSR23lb
r3jNUThMWmWlhv71rBssLrLsliUxRfBHYDnVST81sju5E66O7RUWvt69aHg+0ZJ8E5244+mFe438
/W2KG/s4bn1EwUToMUb6VpRq6X9CESMN77Qt8ruBKmk94OalHZ+EtRX3r821foQeIqpSlGb61Lnn
iWqXZJD5OiPjzGUjbBkYGExPbZGVCqD7M7TQjqKlBik4p1mC29TESaCqr19a9cQDIQqug0BNCu7N
9C8vOG2N1h/DWUaNO0mETAvae0pDsuBSPEBmwaDiCIPVLWdOkGwMNHPPqpk56tpqOjc8wCT8Qxft
zhLapp+hVhPHcB4exZHL7JOtyWdHTdR5rtS7dvwgh1cniIRqmtntkHdTyROK6IzJTw1CJE34pLmK
slN8ovxGsPhAGp1e4rX+4S6PW2w0MTHLeIXBv29cNPfofJxd4HQWdoHLEvm4Ry//yJELov28uLRq
lyEKl0vv7dsTUqAg6Iv1qaW8FxzDMiidy8js+k39RWQrqk1HX+s068A5zWoqJ7HJkqGAq5W90dib
YOsbJ6cjfXwYShWqi2/GLUBaM92H/yppsL7/MWu/TFo2JpL3ElrFqnFo1dGBvsjFmcGlibCtVciJ
j2802Dtd7xaf49xWfNUyzljmjXtg5jUERQBH7EiE2CQkA405bkl8+VVnMp63eGVDSvzXlhxFs+FX
S07lJHReDORZuS9uzohRodjD3/26Drm28HMr0BL0oFzsNM5PqaftbkUPfclij+vr85ezSPSpNbcJ
kBG8NYPaVClPpkCbsb3162qPbd9KgTttPgmPBmGqimp4BMbe64LvF9rFef9/7f6oG8ZSb+dWYAkR
UiZWXC2WoTbxrgpTj4dqvM2gVujTLX+KjLWfwwHpq4M5OWM/95sAoh2D+aMKA+zEvHzuU1nz4xLo
a2qc7LG2uJO6WgSKHxTul8RsiLvhY8Of16jKDGU6P4wa2UKU/Py1mnd+cRleWbpIeF4Kpf3cI0Ez
DvVSjnvBxHzj0ziUKJgawEb2AaAh1RrR6J3xZvevDfxL2gzQdlI5/1I5edhyJkdS0y/xzA771ehD
m4fI5RHf6acklUnfRrYYeRjRI7ezlo0uof4OBS+NgKTxntwrPWJkX+6z1ghN5KDiarb0sDoOND9T
Apc1kO11vJnS+B/cNgW5FcPcFm7Bo9JqULrqtYzG72q55ZpaL31n9bkztKTH/b5yXR9RWzysNiu6
SIIezwUMQE9SnrkHmDKquAyFs4MArXiTgtb9nHahWxRRyYVUEVTvWaOW8Hencu08kg6SKg4JnVYl
yR+m2Q4JIn9NJpPntMs/6w9YYtcuyLmrUBBi4SdkmGE+AiP9Lv0/zPJqGq5HWjID8R4SuAGMsis3
MQLtu+JVnN3dM6nRSOxA6eWx1q8SaMAoXh+5flIwo8fsfO8r90IOucQLSDjP+l4DDgFh4o4jpm2y
RaUkmdimNLM7vrb1aFsuemtxZAgtyp+IEwJIXkRxxU1AxtXiQaoRwYtaL8137txQ6jwgUhoYt/ir
p8RFx6bqbj1mqgZZrp8uSDPZfb/Uh6bkoP1Plw4CyFaYNqeMAdF6kMvSNnS/+/WQP0QGn2QM0B5S
NhOJUU7mz80ey1hlo2Kpurw8DlEGPdf1Op//eaQydqC1uUYCtv98WhFFC0C/SMWPFj87q5M2tSoF
5Jc3EDDuuTZ8E8Vh2YNG2iKsOFN/btLL0b01phoPpgQDfs6BjRHfXIkPHyr/Own1+70nkDtMLdET
aKBemGnNIczsYcAQX1RNjuKloOVr0xLoZY2zU0kp1R+ksjDomrQXRM4HUuWVIYlovDfKR4qHQHUL
DCLg54bY7T4IOzSGGytP/dg0Pp2DrRa7xWk06weCxyoLfqTJHO9oSgfuBZpwiOj50fjG788o6BUY
VfhmRyUn0I7VWgXx+P6Daidl4q4fxRUcoo6g5H6f03cqJJ01c7CkufadlM9KlTSnrLScYJvWW0a1
veAhKycPe7MmCNCwoDWTanqsqNsLJ9BnmfvM0hxrSF0k9QEGMs21mC86jMw6c7kKh+BjBXg5TMrs
VPn3TeKKyD9bwv6//qGPxIdQfJPCSCgZcAmzPG1AM0iQC/8jLAq0OM8jP1ZBOZgf4paieqmyWW3q
CGYUPEsJFsP2X6zZq4Wqjf4A2d9pKUKNE6dKh5yD55By2/fgE0IbKkUS6MDzTgf4SsibUmCX9SZO
ZFKMWMQ5EgbmUHN2fk7KcDTqz3PmLiUyMdi4o0eSYIilB/g3ycYumh4JUi/9oyo1Lyh4rVNG56xa
ADvYPndcpxpcAMYB8V8fa1L5dMyeW1OGiYQAxI5n4m/RN6vxIN6MKpkzEvJ4dsAa3pXuqoHx6eVh
U54JllKn/oKrY2PaYrZXQMAZ/EYrIb640EgHUOQyDAlqN6NZiVT0AfHl8PZu12Xdw14i3KwtUdI0
LWDfT9z5l1vfmDhfjT7ofMbPK0VFVu1EL1ELV61p0NS0LfVQcZwzvvx4T3pRjeSNJl6nq4qou7vt
n/+KESN28W2av7qbuQWa2ZB+hs7/a0Znyl7ig2o1Vcag8aw1OJytbJJ1yuBwGauKxNVVcsDEPTC0
ytG635a/pP88JEVnr/8xIQgv+9ydbFq+VCqfAPm9euCPthxmZzp+L4y5PngQdWbI40nzy9ENs2FW
itpjhp42kTg1PlWVT0/l7+uA5RwDkhjWol/TY6rB1Xk33En0y1Tyr0SxK5N3o4V47CMrhYUzevfv
32Cof7+yv96gLRrbUDtWgLqKzB1Q88oQgb2FKXX7d+DiAj7equE9TGgxz9VbvzJiEvbE2R4rjXbD
xX36YMjZa4h76xfrkelbLvdDpt/QHrNHSnTX3tx2EdCYtGdXNlAKfiGhk8XgFQEFrgGiWxuOfQ0e
Sjm2ehPLXCEadL/pt79n+Ib2/N8bHZgwAPqvda9joDktQ9hO1MLly90LX3SuJ78pHZ0vZCJ02xaH
ojENJzie1EsWEnDR9KXGPxlpubclHW7Vl3aRyoRiuTeGq7MZ4/vOfIXHGfW3b6o24mpwMbbAmQYW
4/7nByj8blbTF5oyqtxMgat+K6gsP8HQxRFrnyRtdP+JeeF3AjZrKjkUHuyY8XozfQcFkOXBE7Wd
0Vnl3wEMuAIhoyF9/x0nFnwvx+qZAexw8zdOC082JIGewaPIffLYcqbxBhLZ0wt/zNQHP+yz5shx
3p3WGNErJVezpDK+ffPliblU+adCpLkJ/mRr4UMxVBBImNqDdzHoq+pQHdz3HGynoFa0ZFBxBB3g
F85KofzCYcBi9cza1WIrz+3YR6vQA4jdttlIIMfiNDXcUCLu8waGhSU/wc4lW80cJnnPZOd5eU3s
opc+cdCUayLd+8SbC4O1tl7xLdApMHDanm6ZXmX+qfBprLTv0RPiy4fcuPQE3TkG0lyj6JM8pfPp
Ck8qHnWE/n1/usdW+XlPIEFlzRo6qJt7Fmfhk8udMSnTCyDUQrwY11tr2OhvqMox6A6yVoWUafRZ
EeymEkMQFy8Hokvx9dJYN65mQU95/2ln6QOh8qx8h2qibffAzYHe/ZN0tPb8HKjWwLOJWqMkK4AT
qJqasC1ThfkEbsD0+nvnRMOFftSPzscG68qsA9TiikkaUBQ8mTuU0YLFyV1/QSVhP+eLmCz+O3Y+
VYnEcgrQTqFukTpQ+YMDJ2ul35uw4Pk8ltWvMsLPRUzNiXdhYvQWzhRVbYDXIzRiwXAEYL2k8VwI
BM2ALbvMlvCJmj9OP7oThx9A42BpDDXU1CEdzm6GOyaL5MojIRkE9xsHl0B7DzMeyVwPGrhqnesS
CB9AR1ZZFZ5+a1BZZ2EK4duITNMYJJ3bvP46jsZFe5g2JEEgCZhQpXKgjUc40tBY539b9qtEWE5H
K38SEBTxk8jwZIc3gjvtu5RfDRmCbhNmkawSoQvUzTNFXwKDuJwH5Ko3DSXhgcb5d2jx9c5DH+Rf
owHW8URlV+JqM5rxxo8wfqaV/7eVPUIbHqqhABMdhvUYce5LgnvoYISaVWTQliw/q8CAxWMNyE5r
dcUcv+1yxBqC1O3GNXoWkTQysFX1CL6BFJ7X5EThzo6iX3JI8TrJ4f0UocGaODmqpbYJTMDdzPtI
BkvgIlqtpx9YX2WTSl+p1PrCLCRHfWW+0xSDTM74fDB+bwI3mGr90048kx+a2Cop+531dry7mUc/
YJLrNF1aoPAtVeT+Mf2pkIqTxRjwmw67P4v75zma5vOzAnB+waMLcEkX6q+iNMpbKC8HWN1/0mj7
VkLOI2d0+ako4/B/GaTaFAetzODzNR8gNRu+UZloL6/Tv4giJfiI4rQMMgMAx6lMxQgx+aGd5ZOF
zsnoQ/243BKnvj3Bucpl4qgllreqgaFGOF/b7dhAhU+KXoEslAFn4PIySJkj+xCqB7zHXmWTA1UU
7XYRZOx8YFu7PNU9ZYPeP1iPeMmjPqWE+0714Wrct7hauNfwIP4g+xeb171R4NP8fomubC2GjtCY
E78rPgafEKNLFxvoTwYRQxDdyXmXZmzr8asxV/xfHfZMkpNWeSz+nRyF4QcCamvAHQI3QNYOTbix
E4zgNmZLpcRuVE0np4NdfwkkzRIZ8491CIRZYV5Ono6opv1Q7pK2dt4Uu4J/nuWx0ytkOOECXE7y
ttD4AY80Ca3FyMofiltfp6uxCCLXoVATewoN87dDcQeiBSVse0RAk5k1iulzf8V/84s+okymrurV
AVG8TlCwc9Au3O38v26QUTyVww2Yq4MYsoKIxHVaCS4gmuRZo7+ApljX6dgaGG2h8t3+mDINjHs6
otUx0NQTz+hXZoNIQVPZAktR+uAPalRuWZqJe1CBAvCoAnUc+PxcfjUNgZi20cOtkILbGV/gMUFB
lKuU2o3kMSYr2pL0MQn7zMoe71y2OtTpxEAezxoRoMjVrXuhklYlsaVlQ8/OlIrtiDJlnw+380dq
CRQjhqztBt1TA1hD6yMTq3UEFLCkh2aFkB9GOX4ofW1MYBuUNfgg0cuWqbSisIBquW0/ehRSeX+C
/cKaBeGWjJa03Wuc4bf+RzEVK7UDkj+6uDGs5AyWKpYrDhydwLW1L/gc3/j38MiKScE7+aB1KSFI
aGMwFgGqK6qEv06/Z+VerWsGihuTwWmwVXUf77kLmwFJ38CLJ65mCUI5gXM/xz/GwQeIs/ztRFvM
R5mzN60kMVw/XpKTg7H7vzusYSe7nSkl0nochDregcZZyQRq7uyR1CiMz1WNE7QmW6tuX5g5pQQf
aIKdHRdYqmKzCamRH2WafcuGYXtW0vkqP72pIga6m0voWEavEXk9wpIru96zlhj8uVjQTGmfRCf7
opvZV5nWY5PQuPOq5lKQRQc+vaOhUccVnZDVhqW5MrTZxTfmu4Z6+Rc3U/Xee99bi4rNErDTY/8b
P04r0FAV7C5Jlfjd6mYxXPqStUi45svuWC7EDjSr8IB83i2JJDw86iruKbJ6N+sXN+sFL6x64eYt
HYaI6MQZsV2d4D6Atdwjd+j14tKA/zsOoe9NYM0uLNjAjlJo5yJUbCf+sgzb39rtL1qIXzv3krGL
5K3gRaCw8gyqAru3/BYx9FscDGwWpn/VCVyc43tZkSHwd2F/b2YE/qTGJjmmxr2uVsYa4d+umYvP
DLO9x0vL8DpmmBO6FdxPWPY/YQINaIoWACIZY/plrVVLTE8+JtGcA1Hd3VEWTngRMwMm7sCyJ6ac
6bBCKyZHaE0FxG66j1GbLRCXMGi+GXt7vZftys0/GTGKKwFaEnEc3ivBNq0gJbtz93esKOG4dzFf
Xbz9u4bqtCMoWQI6fKXKo9GOu8hZdSYebciKoAPJb3v/bcZwlqAqiWxIH7r1jz3A749nTqTrJOnH
yOulFbg636dr5rbqCLUHkEnC/wwPKzCSP2TAandx33WUd0VtVDMgMnwGB3HhCaw/ohgiuqTbzKLl
sSPmWKEli9AYgb4Zsk5rh70GFNaZMGr0/fXeUFDVVU39XAH9ngE7gktUD98g+p4YkNFKpG5mNeTw
QSKFQbyTfMetBYEbHn1fTshrWOxZUfEfi1qD2rED1RznPO5CrgCxxCFyV2iPyZZLLIzmkhWqGHRl
ayonAzDP1OxjNNf9xeGMAxcMuhf5j1eZ11KkQVxNU76KIK4kPEAjZJqBypWiZd+/FLu5KvyqSxVi
+M7awqRpKgHxocZWU0fx/10Bd7xucSzVUcwWBqhy9txsY5amaM7kvf4dZxBrvR8Vn2zbNkPRK8np
+jQ49y4It7bOcwus6Z/aemtnTX3fTFb4Q9AksFD1o54IjDUEfNwVZSTQm4vr9nIXVMe+NGNgEor5
oIa1YAjgKo+sQBLOwW7KO2dZpQJm
`pragma protect end_protected
