/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
nMT6e5UPIBvektIu7NIM+Y5oiceipCd1xX1dgDhwm+LJwvCcHTegEVD6rqUUBB0VpPqQLWPK9uFy
O3uKyUHCKG0yFk8S3uPOckhm+hL9nhiKjsQ8WaNlIewjOu1uNypONPgr6zOKwH/MrXnZ7umAyz7w
BhwNBhZnC1q47thiuFn5vcs/BJ+8GEijKWVJAANlJVtUDidlptGDaKePl6H+n7tYj47fu/82nwDU
gMKbmL2uufn0LiuRUv6uZGu56Obw0bd/wIXip4bvQiHyMHO1WPaKLUpRfvEbfGhjsho5Ry7N8w/H
k4EsVF/w/dw/nnuyt46pocXclMYMYfYqq9pL0Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="UHM/MdfZ7WTWUerAIGhpWNxe6fNAbfTR8fR5mPK6k6c="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52512)
`pragma protect data_block
gXfozn8FyMkuR1aLtPtDzAQns7qJFRHHLYXCdFP1tJMAe/FaP100zHT3sma0TgftuZ4kShMplvhT
dqs6CRewcWYnmC5mYV6kFKUeXNWYUQ0nq4K4CmepaX3W+eIi0Rsh5hR8RVARilwl0gKY64qsexW4
iLKJ4OLuTjSA08bjbr3wMPtllQMGx1l/aVik4sutYge1RtWcB2WbrmJ+/ln5umvWdur2gLmiLlrL
K5nIz7aFoZiu3P7CtsdvquWOda1L3ZgRoN7KCqpyDLfqw2dUpeDrKgPdNVRhVxBkK6J7HGStDVBX
TycazOim/7vPzFn88vdzjO8pWzsgIGlZ0hXhZp6x+viJ6fLSyZgeusLoh86tvs8byUnQ2E5xYLGs
RCfPjzVUCxaiNRi8L88Wl15W5m2YWaOv3SJu6FukSJ1GdJKBtRHIyWWHiYUjfWUFZ7ceHAaBldDl
eAzbQLkrviHUw4Lquc9lWJL0IMJ1FMEORgzVLXGLMHllAPwmObA0jmvE3ukJ3kHjkbz8DuPygK9W
pMA5OBO7v+f1Ri/fX6qJF4ZWbVq6ycZR8pzsrTlvkWoRON0Z/4f0aViLshFt9z8YNVIU+JiJBjFK
YM7KNQeR2+ex9+3rTdc1SN6CKGWAZde9xvKBh+zTX+3gDjCP3RcINC1V6rE3Zjf9LKufBee5Dq20
Q7QKupkmhBvsGnPaUeAG9yLhGI0qazEDpj1lN6+XhgNYtSWGBjPQ+HxnS4q+j1EIwMuJ9cg+ATTX
eEt6AlLWsm1XhKEQAitSC95pFlFRLv+qFRFtTqV251YtT4WUHitzS+lFpHFBewL212hl8IPqYBeI
i4u8AmnS+TlaEKX+wSlAsKfQvizrWZizEAyoUK2t5NDLY+k2n0ON4znaBXKCxqyXjw0JH5G4YTFh
wsmdSNmL0Q4IJMLz4YaDSc/T4xWQe+mguwm2yg/EQvrJmt4uyUI2+Dt2+ajBwFOzvrsWYqyzBxb2
zjQnDvFracyGLts852QG9b3137RsQJhxt9IzYNGJ5O+aMS6cS5YqUMpgeeHwwhSBRIGa5Eq8FPQ1
Rkk/NJhGv7+VOzHmSmjTtM6NzTZ8KI9Ng/dKMhJHHdb12VpQ7djAnztFV1vrLIAjwuu9LMcgd/6s
LaQj3E1wIfiwGEjpByh+cfuJqy4X4mlQCRlKIcH5CHJnqHT5Hh6lD7P47EP8GoUs/1TNUF1ZagyT
sOCGfHdyMnVGyvL/NKeV7rytC01nzjknROEwne3tMUuc34Jk1ljAzJVcO1tTPHmx8HiyHNe6KCjr
Y3dGdV/93z/J6k3UT6sPnNbAx9nirg/zEUwHgi6ju6uMoHjaFc6ESk1d4goRKHSk/sf2aEzbMgxi
Hd2xOFy3oLmo2jVce5cCbj8uhNWJSDWxPx351DDcHz/fg6pwQuOz7D4tZoRap/5SNnoQ4y9t2yHy
UyrQe9jdpygtp7swkUlOILq6z/T8IJ4T6X+4ZplY1Wyf6WE9zV0sEm7h3voNQVVbcD7co/9MlbMT
H7sXO2A48rpRs6yjI/Fgm8kyKymoPelA6Jxk0OOkaOsj/UoJWU2w5YLJ+oJInGSC87c7ebkue5V4
4uqFKKOsfULCYOdl7M6/SxL+6rxYYJrVu+iugjlYNB4SR5orhfRVlAia+RdiLlj2neTHpohsmAsc
w8EqfTjO54azJV4XUePR2nys7DUwSF+5SfwyZEKSNlyfu137Pk8RHsonxbWuFBwTFjR+9aHqT9uw
e+X1rUTS2FCwTbfuyyqWwMuceD+xriXnePJdUPEUduN/ilrFwbwonoHJldFBD2Lq0iJ6X/tm2kR7
6lAVWzfWXNkoQtoq4Q6vh2Ahn7x2W+2+iSmlzUC1cpeYb+wgyLzsFnNS3vbUA6mxI7EWJGsuH/NQ
OFcB8RLSSzyl7IGIe7LB86digjPrxX9wMinFuz2HgjNVmkE6qMSOwH24lR5BTkmQ5/0b2stmJihB
eYBAqEgSNUOOHVhNBUgARTKJNCQ20U4qfuLfdP5pC/835Hx/d+SmiSekw3jtlLHolPyEF52JCCyq
XOBls6FwWgX/AVHYbzep9k+7RKEsthrcP3f9xdjHRkRAO/dBZWds6TmjIYymdt+Cd1LordbPZr9w
8YyNdT4HCzjtf45kxt0ThpDaKmwjUh6yrWMKTpv3PfcmeAaXB71JwDCo4co62wxEMkLXNMjlL/dE
IlFL7CQuecRmTLAkOhr8T8TKbQG0aCBfvMWRxkUhYMAXTJzu5ISTpHS8qV/qEuh6l7Zu9MvLqK1q
RF1JFe9NUD+3HZ0pYNKmwUHxLMo0Ruj2kwDbXKRpiZN+mD3Tp/cjekoK/rLL4kD5ky9pH1qrk/wG
IXYt2cSBkHoTAaSle4jgeWTzuqMaSl7U39DKM6Yn9s51+5/nFyy/5HWGezV6Yt/zNtjvs2+Y7N8N
Zn5pxyn24wq4pnrrx2HRKVFApl0/dknryN2s4EqyBvfRJPRloXmP8YavG82tg8WmK9gPcUFLQHPl
EXCgZSziUK0dBCKnavAZDLcPgE81PMFfKwqtM8ymxsnMD/5KfweL5AWp1zxAkRx5b0oX0y+3XJiB
4TW0TW9pFpMuubOMhEdxqPvVodFLphVGzFI5w6Pc4Hw7h6/c550ewrkUJ9H/ZorofReqVFgd87jV
JlMFOKZuPidK3G9JzemfePFfNH2OSIln7umTMiw3b8h+dLsfZv/cngRfv7gWmh2Ra43GI8HeMX79
jw2oZCtmbFomNZKLDR1vGTDJbPDOlocB38ubtxp35ysIl04EdAYSERvgzlJq5diqhMM3YhRTL5bA
EJGbJ3Y0llcayIKpGjnfAH7AGKSlIIpe9l4RGFmorzDeEMv3TNyst4xEqjaCuryXL9YXBVUaNbye
puVak6487pE5xuF6Jt7ZeSnUuekO8qQ1FeUWtqdAmJRwi/+UAW3MfGUvxBvbrFahaoDA4uQV5T2x
aHA3/hJIAThY7X6emciW4B0rUnUVcTJ1GYXPt4xCLweTRhh1gUiPmhpg6rwJdf+0epsYDpoJZ3Sg
QhMwzOJUGox94lpMyQM8pfj2Zl/Id4CWpqcxR59YUe//IKFy/wz3nnTxVFLtB02JOuTrwQzmaW+D
EdojwNHiui7m7UZCve+aX0x1iFTW1/KkNXvZaIYIS56/b466F43cVPq7JhSBO8nQS7/+tiMOWZUn
QOtSAPu461SD4Ktoqk4FH8tKBFAhyS3KLf56y786jX6EVnhpHwP5zO/nKO2DvuQ4zoxHc0cMCAQW
NfNsopnllVOurYrG2W4pOgDJmTU6QhaDVulEcYwnu4/sGdAn4LHW9RjE0KaxdG9Cl2TbzsfGjLRY
mROQ1PRbSaeeJrMNzUYCahY1lpK8mflz+/u6zCwScRge04k+R2F0as/V24sxOJl/H0o+5emycMTO
t3tpl2VCZO70fbi1XiUN7NkPwwjQ6Zpdzr8LoxbgXA/R4p1ZXevM6Luov/8xWHvUfD15/YaQGvOB
oiMhPhulQv+reF6owe1VhqoN92t5hmush/1jfW9rv09iNcwVdc7uqL7vJJx2yyHkxTLC7kC+PfxR
35g3vu4hDdtsWicV6Et3hyTuIkSZ3DQGQKyLKR6mG478oVpCBMrIuj6kfWuc2oJCWMKXdb3LXkE4
wzwAd/pzlzXurfixtGVZzxi6pZhRnftW+LtgkwUch7Fui/1BmCvZgQlQr+k8OWV/cu633lerDYkn
FJLU71kcx3FchSTuLDFMkqbqGILWCR+6icyeh4+UhGyyYdLBspFhakXVe/kgEnKRqvLGoFZoqhSv
B3MP6RS7FT4D4m5v3Z1UJwddu6YLipuFZSdOQnQy3M29r3PghyfCTw4tHrAAy8VrDv03UXXxgRZh
nGSFVK5q4DJCbRcfWejLQfkCZkpAlTD7Km/DBgDO8H59uXlNxqtXoyQt9REvfKAM8G5icO8W2rtL
JbIiRW2eAf/FsHfCcw3lS6bOEcIOeoh7Es6emiD3Tk/V02qHYXdMSM9fG6vCEgLWmghW14sb1Y+w
40d/4QO+7ApWtu8Evm17jMB8zCD4Mj8PRPGFUh8ufOnIXG/c/3bAsmpUtrkAdiVw0aPX32JYh90k
UZZLWmw6N8kHmF4VDKd19I6/ung7VPnDq8yx5PYqo1nPI2aK/3z7cd61JIcYelaYNVIyGRoN32RT
d57AjTLRLuuNNN+k6rm2N4WEOWJbuTZn7aTHmGN3CPp6TIiuKg15wWEL2lb2pGlO+uryPnGxMEh4
7BUKaFlwgKe/WFHAsd2nMYf/kP68eTz1NITYmTsk2LKGpoqVNM3r3eFbFPK9pDW28QSOVUMu+LvX
BF7znUIwWHjiRzT1hNuRRAe2XVYxu3+Fozd9KYEUe8ExT1OrX3Vyyu5tcC7+bzaaT57C0zNLlNd2
Az+94QEWTu4hEvyvhy8zBBOlDLhr5/2aQOL0IHqpzl6/tUuj5cVU6qsk8NMhaEceNfTfvyzaBA4X
ctVFNg4rHi3Kg9ipwOE/QgLppVemOwIZhdBrm4/m8y77IaPG7krX9F5ob+r4kDqmVJHzSNrUjfnH
ZwB162xjLCsqM3YzCJzqUI/97MkjjUTUzvDJg+dQLH4+WZX7+DMGKtNg5KhxFkVZ+4PGzjDnu1lp
X8ffkgpK0Ggv+revUQRs7loA3PimUfizmjkjikDsgmk1RRlskIqQIQIcghElVcxRf90+v9j7f1Io
TaYpNmveuTtukZBtcPyrvs+fMQ0EABnUbwiSYrVwhxRzvjEFHULfICA8dJwksOD+CIYN0bVmZjg5
gQTSPTCR5P8OCEkTgezOpf/qzF+oed8qcK5IJ5mOtnKvmVFeicNRoqyXxpwriBIILwDmSjPdkKhf
TcbSOPHuBl1DJPMP56s/UvIg+srV7kYHDTb09JYz7sgfoBspNxGpH9o0ZSyMU3r7BPRbZpWiAYFx
FaSn5GgQsfAg8JHFrnryDYjBNCpvaLNJB9gRCSS+U1bfdiHUiyiZ4FyPI/ztJhAxz+pUEg521cKG
iyvqjS3DAf6Jj+ZNMXaF7ItejAxZTFHPW+LhGVRRtzz30n5uFRfXFkOEgdFdKQ077ISzu61qY/Xk
0n2CK6ABD6AcK++AxC6jE/sBuJYY/V12mbu2Sj1OaTujoCg5DRLMU/2CsaSh5mgQhDZQRS0JPaR0
0l91uW/ygr5fj1xuBkDWkU7vc1eDwIgXEBZJY2sVuPd/G7sVV1a0fUEejD+YP0KM9iGRs4jPRbHX
0ZLepMBavvFM74ROl1a9BA1w41QaJh4A1/bRmirEHUrd7eY7svI+JizX7UNpuQXdWSd/vq2EulFJ
Yzb1m/uJ9OrAkFoWFrNF3ATMgHiqRIIKlBKUqH7LVY3f+fgnycr/ex8PYx7rkgBX0VdtvoX1LuRS
K4bJY15SWr/G/PGBOiH/nKCAMBxnJx/AhlSnZYRMNYREr5xR/Gln/f3IPFScjQs8X641yvIug45F
AluOt0ZanUIW2uCatN/mXpfGo2x91CnN4UCNtIFCGpG66/girBDftc7KYMfneC8hIBdp3/2Xn6y2
RYDupS/W94pBMGF8IiYqlRkf68vdvfX4LOWjeq99Qd23vL3/z9eSO/McdBxOSDREhMjC8lC8B98a
FeliZtYERT1PgNRett2cfyvohgFTD29EQlzqahtMlgWya8i25jvbqtU4wSMVu8nNhKordUguSDEi
TLzxDCrSu9oGg/xUSQUjHcvY2ExcbFZ2PrufzkbRYOcd2lkdb3aN2uazeluGWiJVhuH7+rjzALI3
arRKLsznG9XYSXGD3mRFI7I+3V7T9pbG0Dlw8WhFhQ3zk13e9NWi2jHdtIbVDwqLj66flLSx5eLw
vyBTdARTXRzgepxLrN56uaQTia7we3P68O5/Qc3DXfooJEmPvko22IbeGKORzL1uXJF0i2h0bWU9
b0BXYXbeKr+Iy9CMi5LCfr4tzwlC3/bFTXInjTBM8TB8tvldZvbrgU2xgTNFjSgz2pCli76ZY15r
ntxsWwFBdWzdwzr2r9iARartyHToY6qVaGBzZrMLE5WQu0ozisf8ZdNn6OkXpOvmscuA2QHRE1TN
77eKDD0kvcaXtE7uID+pl8PTwvwVaLXhxTZkVl0rTJr2x4ZM2NAqGYhpztwY/zlHtGTPgsmMIKBD
ZCuQZQUkkhnidcqgbnUO/+uk6+Yey/Hqcba0nh9AQuA5SVG8JWx1dHDtQuR2dqvY8KYi2CjSYmJI
UrP6cYvJUweskQw6/2HJmdYsuHksfpnEIKo70bAL+AsYF28cZ1/TVAMrYiTUYgxDs8j+jIt6r8wf
q2hHbk4bcuwybtiPoz96I8df9l5lLOOxgofVDqialY1H/viSt8RzFQNNWtBZEWcIf5k0y9XerIaO
DPbXt998gIFJzbV56M+EMevmeAJQfaMNFL9zrubXF6QZlyVyJOn/osUHfWrdob0efCZPSWepBrZS
N/uSVVKbZ30RFyKjlNH+aSIF+S6EoBDGNKPTk8a5ROriZPcftqss65jMAfAJsVH8aBGgLXHP9p/+
2cvdNU/zbG3ecNXMCmpiopCRGIEXoPcfEiauz2zUm774yciCIOrKS7jcEz9j8g7fj7aIC2lreE8K
141JX14qXNGXtyRyTmIrZtc7Xb0m1jRLjh166zNsSqJL1yyuJm5hr1QZve2KKm1xK0qds0/HRrWt
NdtZQ3tTJj+Hb+sorvCcRsckDqv+l0DP+OAx3A6ajLrjuc2EHDL/mu98SIS+FnOXrrMjc8TQcCA1
3iraTQvGLYFjvCIVcfDf7zF2jevkKfxJtfQhCXgnrKjOS3hI6Zw71W/JgUWS2IlD7pnFxUUI5/DX
r/2RvL8Bp9u1032Hvekb8bLlVKgvZ7HpQfBsI6xze39WV5RD5VUcBeAT5UrWWu+IuhuQ90/cZ3KQ
Xk4+7oL9O+he512ume3c/6vGF0qmOONi2TP99nonZjLseqBDtzjfCrj+mD68oKYkZ7wuo5dt6Iaf
EzM3W/L+jtR/R528vlooy1wDzWCGuljv6lmUdzzNrtun4dcf50pvmG0B9S7+fUj8D2fNvUQ+klhe
CTf02g0dbZD7MsEQMGTMaA7VXiXsxa5cXg7TIrsz6IGaLcw4f/O+FCwZypaI+Ca3YW+7kdXDkLad
OI3u2fhQF+cqhi8GTSir2cMYPXz6C8ptd32u8XqKSaF35ogbJVHWApqagCOFVi9/AdEjkchZjK7H
lkNzgJqKKP2cznAcoagq5oQPWXYfyGDeOvVABdxrgw/sRfySsTIZ9TG+ARr7NPL1IKiFYqsrBCBR
IixwAzGB7uysb2BRolPFkYeyxl3kQ7upqDjtyjfTLUTmaJvAIRECIuL4oO4WoQDDnOhZqrZFelDj
cB1AAL65y4I+mQCFuyjWhwnXSk6VYmzMdiv5QzJZ9okCGkt28zyXr4WvkJ1i1EdEESN1ZDstHV9N
cIrAXeDjNlzXKzNmsWwA+z5ZIpJWlThTrHuwaX5KYmt1DCoBdmNqL5sQVPS3cjdE64i1W1aJI3Wd
Th8UpR0ALIPGSV4z7CGfeXD8ETIXExp/RPdrv8kh4fMWimfvd6jlZpz3CZtl5mion7M/bzwmwKkj
2FHN196e+229VYj+Nb8wxrIh3a0wtQ6QWoe7uI5FPqKwEFjcd4exVrvvdG2hCvq2w446Q6tF7U+A
h2vz8IioyXBd5mwX/5AGN5jThMMQRYlBfVTR/wDxJEjP9NmrGc1YLCVcsdrzPhhsZa4ycE4VPvnV
xZi5wa9itdTqNHle8pLku/GRya7PDnRIBVIi21Lrl8z43REbiXb8CUYu+FgDp7mwx/YC7Q+RZ887
sGUVg3PRRLV0jMscXufFNI8YQKbAJN8ywnSo7UZ+ZOQgtmM9FtT3PMsbfs2e70Jdge/KKKDxZqI4
mQTlRmQINkEnu3DF8jO/V403tWm2E8AW3bzPLg1RlLTYM8NyWjEVbHERli5LivKsA7yRqSec9udH
kApolkbxhAUu00eMm2eE+a6kMu8GZkiG7L3jEWr5vJ685aKrVo5zy+uP27VUueP8spMXJc54oaIi
fY1IMeDo8Jqvz0JHlCg9dUZVpU6huz9B2CoSMhSqzyL6B57gtVlDKACMGZSKRHO4pMjOdJYdWxuz
mx/a+wYP6hrGQrLmgg671Y90o+wtv3EyY8yvhrlWOXXsSMIljun5jEi4eyKqQYCxs7WclhZvC3Kb
rBDqxQesZfl4JfIceKAB91ifkjDZ1FuW8wKA2zeIzST3vWIHliboB9jOQZ3r9pLHDqxoYAbd/7fR
r14Lgwq/ceXRrTOwLV/fOels8tzffNs3A+XLuSdkj1rZ1+G+NxVVqvk5N4Fgc/ibn5GMnWutXXTO
Gxxbivyur4FmdEuc1NQWbvNpWIs+u7sZ8WPusBWNkbByKgGy44XwVyVFgpu7Gt/hBf2hwbuSNNT+
mvtfCUybOw7FLyW8h/VRIVVmOwacRu5MwPvK9UQ/seboEXnBFadfI18YodPY/Wzak7d/qN+SPmJi
2gChz/xYWAWvknqyFzBictJ0QM6bovXYE1NE3GY9UM6dGJvrZ8PaE8RJvYIYXYZ+Vq1bakmYLjOA
uGLjHUpAldi84Db2bpGj+xfWgmTP/Na9YgUt5nCFRs9NXIR9TdgAXhIyfxiTvORNONlfsMeVviPc
1JsjRPuBzGwJRy/MS+Yrq5NPcb4MaRK1bHMOK2v7bsinOtVavUmNsoTg4oujb5cuW1hcuyRhM+f/
PwK8Gm++OGjpPeK6a0MkpH/p2BpP2OzjGjPCXsVMnB6WyOJay6Or4GLe6EAQAwjTx1NPSnSUIvYN
5w7Gwm4pTeMnR6m0M8QQDVQw3QrO5fDofY4DAfE0CMk1ykKhPkpZaWny4oB+Lcin/jHH1MVH9jxT
oWoey9uRWh4rGbqI2Gb/T1ULvEEI5t/aCxvVkbY0vGomAO0X7eRr1/TszRBvKFf64gu0drB4uqCu
80HW+aiUwohDk4j9LiZhVgAXXqDLFjT8Skj8o8iWCtlzVc5sI8qwhlDCS9yBGQ3Ro1uH3klk3Psx
RQp6tstEw79vQ5U/potp3QEtcIj/EfHCYsMVJJojh11wQeKnukYy79U6UFEOSZXscMEwHkjpDeXY
TMOGUaYwH9mpJ3gzitrjfecj5pRRgigQVW+PaGQwp7TCMSbyU66ok/4sWpn+TItyK+9n0rb5xNx1
RRRXixZCIfgoB35fVYF/2BcFN9ycOOAgYMCe6xEhQFG/zm7fl6qxO9LUaHFKor5aRI/ROKSXE/tw
7c4MmCFHLTPWkwtlhNi0WYTqjOKnrTGez+pHbypyVcRdfM5lp2GG8wpQdFNb/Q3JFMbG8ot6RHSy
pwMIEA7xXs1yewmV2UctW6ic/BLVxLP2EELIsVC+1rnI1Wgh2Z/qBXv7R4Pj03I1zrDPSa0Bj2AP
j5A4Bc6zmAPL+TuO7D56HYpcCoTrkuN/OhQo+/k+oV7clXu7eLhqZFGI7wdNR9/K6VwgWwZFA3eS
X6rOPdtxOgsWRjDE+FtczxImEqQKSddXh/hOsEt3Z5B8MEWdkILheaqVB0FUpqkRJ2MiXf8EQeaM
011xt7THpszsaB2c5xYwmXrrO9A4rCkwIDvMOS6WKVJj4QPzOPY+SPEz/p9H9ED9NM7h9TYSS+cA
6p/qj+h+xseoH34M1pZMbkNqtYSw5hV3irrJgXhz+Wy3j1ZQ+gevPKmiI3GW8VbSzGJ7ENgclhCs
KgydEGIYE/EXMAxYyd7aO0p4v0nPPYiIFf/D7fqfYQpobVX/3hen4POGEiOGcKTR6PyE+lImh1+3
sShTIotC/746k92/n4yQUD03/y+po/r4iNzyow2E3RrGetom1okPXf1KqLyfB9FMMlk6pkDis7Bw
GPfEKg2NEAORGD3vUx8PCHQK4Pf6QEDIhbMWyD8QNyzHxXjphzXY3ZsgJKfIBbdTWaD+piOh8Rcm
rhi+HHm4KFHRLWDj9KCEoEB5bWK7u0f7jawgRV63St6jy7Di+xaeTm8oKRPEFbKP4nRugm/J9Iq9
C2S7Ooy1Hx4St6RHF4j34m/7LX4YiKKROzB1k+l8yWBSxgojxkuU0XX+6u2x5xluM7UeqfYSDemE
RUJyLroP7tuyhf4yOwiMlMQEKC27AawOHZjWF2VvOBIqYQx0VoJXPJBjrbqDUX00KtnZUoMw/21n
DdoMSdi7cJU+6HOsVMuI30+fTWnq8ola8VM//6K+JWfTjeBE+5g8uQmCJfG/KHoH+6mrvj56TdcP
Y/ewaQVn/l/LfVqxsTRcWy2q0UOi9Z1EFPNPARPMQahkVmsXWn1zx0bP3UdRMik184UZ2NQH3lqX
JdzHzrk4wxVyQjAXJGFHwONQRJKSsAa2bvs3bnbubseug1klKNOhkO6HYyU2OBME263Op7bsajkA
aHv9nFLkLepJxNM5w27MkBYg0CgJ2YXFC+lMakLUmcmtTQUWMnAZKHgHZlm2fP2Ofc/mrzqamgqi
eJrYgtYlg7noI/mUsXxAU8CarLJKsoN8AbdlbIvp9pI5gakzzKVOKjlcQd9kuI+L7m+hHtG+AXip
tqz6HkSDBv2lyrYyyPnvjiDQzJRbBHSEC9QG3WtUmgwVVdqdbhK5sAq/L/h91izeecaI+NQR9CFU
GA+u8oKY6CsBhLLYF9z3rhiJoMU5P5Vlqbf/vOFytAskn4MCEpptIB0NvLhIgB9oqnhYyMdJsLZ6
6rZDRIk4acR7LxOpThd20618yFSjKQ79GnAZdPKY6fagRuuz9UXhnFEDkLlxJkhKe6iZZjd/qrMs
YrzX8Y21tQ40vyhMY1u03RIVOKXt+rr4ZUaSmqoLsZTtTnknAUg/RnYE9b+cCSZsSvTlBoGQT7LV
nvls4ifbm1gjYpMD/Q6LQXLAZbqmRMp4C4FIjWNjvUgKmETGHyQWpoma8e5uhxNLuRgkCyEGFzwg
GcEVQxf5mipN/nWlQYWRK3xiPJlsDtD2IbHCmrXfEQmLXP/AuqjgYKeLmxxyLoqiGdwUpNBMM1ED
ibtG5KMgQUhuVmXeSezJCgtK+mHQB7Sqr0lsIJak0sbcXgrFr/N0e4t1Q2+xCjmKER4KF3AtEHoo
116WUdeUq1udkzfOjqgC2ovoAMgjMJH/xO03X5hWe4kh3/kJT4dl8Mt0JzrjK7T6rcDNEFkKra8N
3s75JzvDgP1tn5saIWSWOKFAgM1GEHtZ8d9i3IwrYQrEnqld45VMly3k8KnBGCu1UdWxMHF5bR9R
u1Tfw+gb2aSYHQ69Ot+NLKPeOChJwzut7F7j9PHWv255edq3dEH4LOKsA1CF9m7zARg6HV/c0lHg
CkM24R6fccGOvD1UGSV4w0c/CTcxc3+NZ6I3JP65bZ8oDOtP6GjMcA1UG73K4PsfnANJiQ6ZlnCk
PeM8aHKfItgJLh84NKAFep1uamRh5S7KCXs9eSEk8Z98eoEqTZ58QNcQoXs7PxOhRTvG8GZatj+o
MwsXoo/WWT9UXEtUKwCLY9DHcApCobUBmcsXU6PO8mj3sJSwks9AUigPukeHyNv1bDrHPn2fzcXT
fJeVyJU8bkDkmpojdv6IWiE1HRrAmsVQ3PBTm7BD2Sg5VN17WPsYrPxybfnOW9m1e0unUV5HXxz9
JN2OwTn9nFuiSZ0X10Xt7qGk8X/uB9ybRiJKYVGKzR9f6hTItk2uHMKkq12RBt8c1qhsT2MiQU/+
S0g073ixAC7Mibq02EVZ5a6dwmQLPNey6umLsMB7OZnbhTJnPZeOt8IDRD63RU8fT+l1JWprvwKI
jubL0laxf9ErxJJP+5vm6aI7YQUray8y01ch0MzzZpGYyDuGqgI4NcQuY7iY9dkuGxBJHf4Hhuyh
EmfbeLnNco27QEDbSeEk52NgNIjOJn91BnjW9P2Uf7IZerlvZrfK/ST+p6v18zOode+ii0vDHU8y
pBaEyDEL1TzMOb+ThRp6nJlgpFsbXkzdCSI9sdiBaFOqmMgCLWZoNsz8/vM5VgWRusTN5R5DLZ2L
X0TzRGeV6l4Jl/BUCPOrF0TLWzFFtOeWeZ13zYYcT+jYCQXDMtDHweZxikgQhJeDWz6BACTI8g1v
O4/wTTfnYbc4cEWe3fauK7USxGuw4B8QGY4YFJjDKGvnd3uwQUvTfrcuMdwfABew5V+B1DC22Hb0
mh7X4MHv2SWzaohFxiLWpv0Px4v4RkUlzXeyULj814RGLeGc5q1YBULO6vpV+FL0CNBhBaMT2JHA
76Dj1RDREppnf5ZFx0LRjD2td685cMYA70hW773LzZfwE06m/ESDTWQC/5e5gCA2rxQ+ukSu6YvZ
Oq0VyUdxfxgCEsFlwCu4svS8fK2oCfGXO/E6BnG4n/9OQ5HuQSo4wfH1HK2kQ2zLjm06FAzDi3/Z
CAm4p2/H8ZBaAXykSGM1Eh7xb2vyRPs7EKBEBYsUpfm62AXePFSKeNad9HRa5CVmF4tmji46Zw48
6dvK2joxT9uZligngbMn0b/+ighd+7uWgsPUNNHL7k2V/syXyES1FIyrAePklMA789McWwN57FTK
oGnDgMmwV85op4uJcmB9gKSX6c3MO7y2Ubpg46hqdOi8UCOzBCx3B4Ng5BZUUKWiZ8nC8r7eXvCg
xoltLMDZLEPX3zFue47uQa/PtsCSAE3xNHEcTX+taW++9xvYNMQ2CxaXaH1yGhzcckpyiDdS6Abq
DlZ85fuEKXE4myJp0LXxqSALzuVPbayCGUemeJsvX/+87TozgkkLIgDfqZxslzFKS7DJPYxlj1pj
R+DjRT40NylTREojzw8ymZHNbgLA1016X/1MUJZyjUpTQsP2Qwfx7thQCS6ZtVfYItN+LPDpOzQY
Q/YMqCRgciOgBa7VG7EV5Ddsxm+WA9gPIrVupyWEX8oOnIl+rQRIJ/FN8VkfYD71bxJ2ZB34mUvl
JAe3v9z9MiX4Vv12ZP7IxKwB9YbZNYR+U6rd7z7zFqq8rEHhGGBZOZYfsfc2YbH0i4hKoQsHGYIc
kQvwHFIjj3xrt0zdT6ZP5rRGRhS7XfdQGuPw1uEHbDlnpEdoEOMyB8Jhfj70fBZQh3XYORddsx/5
Bqj3THwfKHle6N9d0XXO1lv9ch9PzlwRUENpsTFOZ8+QTckZpFniQ7xl2ky/rbTNyPUdNpXo3TeW
AE4+3bHruN6Wt5axjIVOAtKNDQZEozYuGEK2excPFpn6rnLZAIBKQAF7qstTfxU/L3H+Zt9kSPnM
sMfvIwuQv2ychwcbTfcytFYhC/BIVjtqlXo771NYDoYQGCW4dg+riJRur0jpXDxGsf+nluMqm0mU
FMJ1TCVZn/+pWb0fxoWpJkOLhsvtoMWn0f8jREJJ6youo2o1UsIBysMp1STnFr+0Q2Jb2LV6L4MM
EOdisb3zVQKTs5H3TT91VNAo2MgbLmL7Xla45nRYmp5TeEskMzU3rPPQZWVojwBUNo12+i14WZLv
QDjREPHS2xly8bfJK/sl6vgcoghwzprqO2R6ULrRIrlsmmQnez7u/5FYtt1ayR3zXRSBiMP9aAa9
uLzdW1se6nf1qbM7g+UBIrlsdJyI0/tmer/cSTQz7jPo1nsA7ErglA7Lj9JCaMHsvN//xPJVCtCb
+9r929CZx3PpNc28QLo8zW15kslZgHD4KOJooJLSEgaHiumDb/8yQtECi7jpl1LLQj2PvD4Ao2j3
ANIdcx9FHgi+h1K13q7D53Xu2Obq8Zw9mOK+oxV6Y82FwVFupU+x8OtMnMWCPNPaiuhEPQLhIBXa
hlQvZqfVXQDDvG+wf+tsKmDHCWEvEI9uC1alpKIAF0BZKrehhGx0C9H9gzmgK45YcmZZkfXDNIAK
gxlO7KVZkKyrIk94C2hfZCXDuQkuGWKbA2RDPgu2tRLYsFOf2Q6ksWvv3XQ9/bzt1OtgJ+X0Zc8C
WYQXi2M2u0xQhC5KDWaKnUfHBE/UHJZcKk/jIrnERxq87OSmIBM0F4oyAY8dAgPqe83n+7UBxPpZ
5U99/R98E3P0CA3Exwt2Oj7TDh02EZ7asZeQObnUz5S4aaJM9WQVKA1gAnAUXcffT5VjuOXXZkaW
1glPnqJpKawj8H3pYrffCY5iHLAcpbAozCNzMyg6+Mu8E69ZtA47LmJIhrzCRmGS2bwVSLZOfa21
VDfBDcvuX4necDmgyKAuxw3rPomiQvRDC+Ctae96nhRzgISwVgmMyFnh8j8mosoULBtRWUxrF0NB
WbRWvG9B/7NhCsHf3qXqCer8aK2+QIAk+3aNjRg56bGY8Nx4Q+7v3mpCit61GEZjq0AqsTs2sChg
qKyTMGWOGoYI+NoxoIkBei+4mlAT0OQILBXKMArWEbDBGGKtQs0bSGXMnvXVJO9n9FBuCHZp94k1
mNq8eCRAMD9DIxikg22yDo/i73GY0Se3GttMQ6UhGxsRiP8qWNIC0SNIgL7yU9AAYc0kpM2YfqRx
ghjc8twRyx9LPk2U6u6cKPgmAwxtlyoDP3K0UrTdeUSi+m7xIcZzr6zDMeVqeXhO0uRQVSZIexmR
AZf/ZCa4v9Evj2OauI2ZoWjrZ1vQOyrLvbmdp1+wOR0oLO4Bs6nUYE44B+P86+VlkIcdvHz+HVhN
3RAIoUulcMRLYjWZHqPF5NDWSD//tzfxhPBo6hES7VUt5qNjodRbHe008Q1hvaAeAAj+J/OYVUC9
S+LEOQwd6wZO6LFZgOgfbOC65XyhCi2F5A4ZBrmhRSO+YamVbQ0UFkeJ6Pn80t9nykUAuHU1Mwfg
lQC49V+LyKyFuO+ez+R9ifYM7M1khsBBWgC8k7FRbEQhspZO6vWG5NUCUWhhPjJsRhm/oq1Z4ak6
ie4Kh4A6G1VvDE8/dlhyTh/hqfnyhLOKiRTLU+JoBzYP3WsAECThZrZay4vkQto1dyaSQb/7xjlm
LbpqRKHkt6WAf01ZB72fISCU7aB5tqHw+ipYOzYMchhZQX4dhDu/YwNsKCPTPCzkUUV2J/YwOVeM
fiZ9gz/QrnRTCQvVRYag04LXfaUg0m6FLIWP+qKo/nRBg+oAzJ1mEjOmbYtD5smrf3zKB1RkaX0t
9xQvm9koKWasRtjPBwnLikdEbV9uNRI07ZwFJ/r55vdO1akJzKHle3Y+r71JZX+b0DeOpfBChtTc
XWMBN81mOh13U+aPgmapwvXa5QrsHutovcG0TeMrvV85TIDLmxF3KLQ70EoHWL8umQnMyWB3OEmr
tt6T6FWhTohlSyXBfwV2WrRx7yfTGknq7xfH11unDdx+DStbMDcJwaCudDgFzcehLIJwJdw6hWNR
aG8raDMrjA6kICPuQh1el6Kof+YFoI6uVNGkRgEz2gdYWl7PT4VqMY2w0NPcjsa5ELp0LKMyI2U1
4+JeMP//t3XqJ+zBBfkLX3JKSid4IKTAmjf9SfgoopHzynBIPMWtolKfRy07bdAiwOjk2qGuGDnY
18LlBQDPNkxIaPpjvcdpfe+NN30aS6MDS+IjBHBNwothWp1VeRo0DB6EspkBCh1V9GCF802vliEj
gLzDK1DbzjEzovZcV6svrWyfgd+pyUiGnZ8pM7UK5mRXkfgHEsAmic8QoeI5fkMFyVRv4Aok7LAm
VtwDyv4wRsL3qCJErgD8yBtE51xOZGXx0t9SM5XMBoW0C7TCj3wJERYmXV0lu53u90PzMXdUs3SH
oCJzVxGfm9abxizO2BUCZ/pQ2O9ryYycK5nqbgHhf3fXDOKMwtuwD3Ne7IrjgXzxO4BBJQVaoLLA
8FwWt2iw++BIvduqqhQTqWwyLkdbfCqh/dZzcaexgzntvXVyr7a3j2PQA6fqF9Zhwn7gJMWR3Llk
YsilCKhpwtkn0D8JbJmxJ5cOc5vkpN6x7xsdwAkLyDSI4qVNWTjcuMX4Itka34HOQS6A2ClrlYVV
iBL/XU04OL5KH9ly6eGXqXXXwx+pPcw87aOUC8+8/r3hFyKVzQ54iTTS0JSW39vDctvKEIRo5LgH
CfJyW9ldfGB7DkmvFZdWMQKrhskDyyFxkud0dtcLGQlQplD97N1xrsevbrzSe46g93Vr1OSybiDn
l9WqW3xCoi+UG/oiXHHN5hm+AdaLV5BupdTcZMTx/TCrqy8cnZURq6wO+2yIozun368euyqhlEOO
7KdFTShqr6uMiXJ2+m2D+WR8wr6q7Ayv8nhWBFm063WXfvHbDSZFqk7bwwkZ/bU+9n0Kd+98cO4S
4j9jn8EOzMGEGF+A96jQM7vF1XkdyR1M+NgZ+sRjEMFHrOnEQZyo5O6fr98gFqs3ziiR8Cl+Nk1f
xwm2ZTgGnkMHL38SZKV1dxOP1DyPOU30pJSWjyhRJ612Hf98rRCjGIKJw7f2aj5X2GmaHD9BrkcY
8cLbaoFQ5xEqNw9pi5pn0TR/CNd2Rfk4VxutGdOayDP++qYaE8mfssd9u9p/5yKBfHzhwJLRraJP
OFP63YfMlXy5ZYBpe0D445GbgbwfZo39cQEEclJ3pWooJE5mCZbHYK0u98L98FBax+1Dz7+l7fX6
RCajor9bppoBBdumLBRMCC4Wb1SJ9xb611qKkIdH5/uF4tZh823/25v7E1/FIb0/fRSi3Ms7IjMN
eK+uQwLUKGkj5jLAOU24N6HaqoJUyIn9c7zjGH5e3lvdGhomvt2Z+0hxbY94Y1n0BDX2JO6JXmk2
yOM99G5Oq2JYpaoMx8iirTlI8GG0Nx6lAI7gZL5+vxYfmelb1z40IgsqbYZGBt3jwwn/Ec8XhDTF
kb6LTCLX2XlosQIYYOHXu+IAcpFx9FyAERsYB9DeWj+/ND+B7+r2aeK9QFuCk8PC9JNmAa5RHAzb
5pBaYFPvWEED0tUDugwLuTYntY3UD6Tv6WHWMBHzUj4JJuqiAejX3V6HMXOulcA4vjttd8OOqhSW
pmohC8JWmQmubkUQ0RU4ynFWBXHWUJhQEwpueQ5rmbwJcANP8++YXR0ZJ19C87XF/OdeVpPr5rxC
ENCQMn6Vo8ctfKmYU3q435OpbDU7FHSsiYo4BJ8bPVYLOwmTta78S5k25pytFf1pvd4M7xsqnlJT
/NLi7+k/tGVcW4KgnaRFUgaeTlXvNCq1jtSfJga3gJuNW5c7nIqX+fiMtlQmCP55YugwzY2FBmeH
UvioptmdgT0iC9aPATiTrDQcUQZ/sBiGs6PJZgH0oNpIZrTYHu4BhDyArt+2NYaGqNnyxtsT1yZe
hnwX0uhu21bUmv6a499BPdLkiE+kuWZtLqnf2E+xw9aZ8N7CCeaejs1bGXzxeJXmN56EHRbdg6n9
w2jt+zLwmYDUrgUeTnCenQZ83//K+BD1FIk7mfy1/OiNyDPghevFW+x5EeSxXmpaoD5LhHKVNuUH
eNY3Uya/59t9E5NLplvWr5BBuCMisihvJ/aVVk/A5TTRvwM6GEXNn4dJsonj3oJmDYrvzixEPjZN
+A80np3nTjDG83pF6N6Sem0HkLMGTBeyT+HameeO36foyE4k4pAkRNP7Kqvq5dQ5+u+4/mBIbEx1
e6Hg2WF6nmk/5HFot6xPh2weLyc1d8R45tyLQ1cH3J/1WHo+hcN2IGYNJ6I4BdDlJW5vxvPogelU
I5T1ujwEaSSl6hzh2fyd1wr4CNjgTLa4u9qY+mVh8VV5n4ykRytWfcqF5A+7zXj85ViO/5tvEjxa
Tq3dyM3ags0KDjvA16MBudvGgDWziaaNIWzOx/ptOqMikiewMcXyerX7oC5IMYWBU5DBZ/OeiYsL
56EuDci9Vxg1FWlGglggaJMZJO+EyNX5HiMckS6CLfswWk7VGPF1D5C5GHja6eyqcnhjhCOsUkZQ
V+xCiH1YV3mPnKVUSNM5hXAMx86rI80yVUXzOh/ZLTof/btUDx1XLI209IpwvbbP+In5VkZ5kus7
FR+6OcBvpN1lDp3cTvsvt8wgzksZg5QhIaWm5vfHGXO+RWXUdShyJ2Z+wZDawO7zK0P2l9Qd6wln
xMwUBHCumqFv/Ck5gm6RjaVLjZ9EqX2wIQLjePaNMUZtWNTST2mUtnsmNww3wrWiRmk1G2LCxA0V
gRDf2qMEZ9TZ0oYO5VCUOoVwown/6nF2GSSrAASsQNkjbIa+LxDfBxSlhjA0KIlynGevyhtdnmWg
DODGFcZNa3C6QQXHfdPxL/UNLixuI3wbi07BPXqLV8V2RZCfIbGE5SYcVLdp18kKEdT0Qz82IvGx
GAbjgcQPZBS2cKEeNBaVKLroX6HBNL0QxXV6wmSE2pDzlpz8CaIlSf0kc9TQAjFFy6b7psQyyACK
5Ll1QkPBUAmjfdeq7fpXarVrSF8tbzFdfwYItYLDzf0W+WyJi9dtBmMb0fYTFwi8ALKi+b+ccuSk
vplKUBW9Q7jGMyZT2JDD8zG61AyciFWYhQWDTMnXHoDP9gPbzDPDj7IWxZ3traU3alujDC5v1B9b
rKj1O+opsuD6rocjeNjxlRucYADoRnVg7WK80kUyFGG0krCEzAMI/pBcXJW6Sy/0x8/v3Gif9a7P
vEJY921JOOEe7XA84xCmu+vY4r26AIxLqPlvuZv7UGrsruhxdfg2gAQQAi49XY8kD324RT770cLP
CeLg5+/23LRLJRgaw/MDyJWJJ5UdmJAsHvDuLX382HGZf5vyA/CQfqv2eEFkLJxCiRaYbtV78Iim
Z4/vBl9JLq8NOhhEDfuwCI6PSF50km+PD/1ABR7I3GH7OnKYYXl4WrjDykLxQo+z2DRx1cOWmKwr
mbf4vYgsTI/Xazfck6sM16AzF0UfIfA0Kp5NbzXjlXQBI99BKfDqp4a6IdWXKUTxDaWUp9jquukY
pcCcUrC4QxIdJyf1wD8ZToKTCns1Gz+YyFK34D35abe/T+sfRiv9A1sIHJ2BwkB887a2EuJBwYqz
uUBAu3jnj7QqJLd6loHbG8fz+tN62cpI89cHKXColoL2qThYL/AFuPe9GIXZodeteO8E0uZwA5a4
5wooEWf194N6+LMR464DKxggoPvlhQtTdbpRymVXitC6w55QNEreThM9rr7aDMCfAhnO6m4orSrQ
eLeQY+sDCxQ/C6CfQniuZg8XDk9n2NIHwvtfGFHMSrqTHbYhRA31ksUGdmb9rL+mI1JZRCqF5Sz1
cG//tnGlMy/j4wGykS7NJx7KLxwjWgMQkWrpT6ttb7CaQ+GojkRCAqBMHMb+/3VrTUeukJx+cwuO
2FikdrpVbncKpuOSre6aquVsF/dImK3kqTKh6ljPE5lirc56LcMe3GCqzXn0/+BMyT2H20zTBob4
Hp76uW5TVUFjKQwP7g002UqLBdwWAo/SgPVokloCv4F5Xq9FcM+aoxMoB8rDoGOx28TEhbaBI4Sc
JzPctIVrOPbeSHbvHG+V1PiTh+Dk9rH3n+ta5jLYdzU4MudYuOtdK+WXGTxdqhff4AWBeIbYwqVa
FZ/ixbZIBuNVn7CaGw5NRJUZs+iOHuRvAsRYNF+HxRInJuf3O+gMS8oNd+kBLfMzVU/Wx8B4zSXn
ZMPoVZI4Nl20IGtFtVVUN8lOLsOxH3q/CqKKxtTXza4Tr4Ns442CxnJP24K7KsI4AL++OA22/+7U
sWVKPdBapVV7kZ/EFMk+Vu4opqGCSr1TV190YSVjNst6taYa3qbTmlRvUd5sGZZERDe9KnOTsmHC
roOyNhrBGFaihEL3Y3kQGtyDHqUwef8BPUie73+pl3z6KXPnw7mlbF2wLTKh5o5OcCJ7EhRF+HsU
AN19yzLNpGWfTe7VOhlGIiGGanxFmRXGOmCStEGbE8lVrUuu8Jx9kP/7t1hx0PXW/DTrcc51C7dV
iYbjG0YojFBeEK4VEVlq5T61myC0ue0MzCN//gT2d9bftteMwswuYfv1rWaDFkOnYHgQQm187bk1
5lEDFKaE0eIjDv/nRwMPQXqfkH0R3PBgwcwa/HDcN0LNUDMGFqO6nDewU4HlcVTfNEMn4Bb/6czw
whaklyKfEUXU4Z7ROmi6iGGN5xieh5liLF2CjX2VjaRIiyaAzdVPMyODa/tqPlBQ59qIZZlpHjD3
46246KSOXtfuGiXbNx8CVi662Lec66S2RTSi3WgIfrQ2NerhbgxQHBB1y7ot0MzezsWni2Aro3Z1
tVG1OgyFQ/WvLNIGIeCMC31MT6Zl1Ae05F/Mm3wbIKNTDqbF3a0v8Cpqau9pZy73ZbLar0Iv6Y48
7TQK7kjaaCK0a4amr08d5VS0TdD6ghNZqrmG+JWNwGGCbLQQj6OYdl6kXx3y/IKpCAF0A3cGE2CS
VnMp710zqB+cPv0OGPQvEur9ZsBuoHTarsVgSPNmADLbsS+IQLpnEYa7vTD3trVRqpHjh0bKhNZM
eqhhx0PawGyncafP8Q85nZA9GemJCCo+QkfE7DFlNNRFolv8lVqHKtdsz2gLaDD1SnZEL4ytQGiH
rdZdpFC5llnfSTJ0Jnd3ZeqV3sxnwoppaJOpYPWVUuFxmj4zv72SnG0kDlZCiB5HsItqVG1QIwLF
DbuLmKi5OZyHGyWr4k8cgHCfW6gc0yyQNvVYCFy/NB2ZlpW1ItoQkLXWEA1SdEeiVGZixSMU2hmA
PZVuAUlZq+3M6dXnfON6oteah2dzieS1U0BM10VjkZKKKW7MzvXwzVZMhcoIoxTaxKQEKv4HY7AE
Ysm5qUIyn+Uf8oQXyBTZTUZjGGcrG2XIWTJ2GiQ+pIgjrwQnMOgSShHCngyfbDBOWny+d5KqHmWP
LHr1hzNnHvbD3ZIkt1trcjCRZuXcpsu41qmb+HF7LW+dYvcFYemfJhPst2e314orgJp70/fSLfW8
BDnDRA8qLcCIlNo8yHPINhs73ZcFNNwLjqYt4t95DV3MT7TzZRAEzIsgzumqmAgNiYkVV/MrL/1v
JFUfvBqQAlT41pqRrhsrTsRS9qsH4oWqMHjJUmKJnPRczkRW6vl6WEmjK3SqAyXy5MHAXWqyKwmq
zWv97HzgM264vacXxSyLIjZUdZpLs/gwTFF8P9EbE2PD8yloQc9+HoT/BvZ92fvMbJqyW1+PQn5x
JS+faTulQeKz5EAPsRcx0KcOb9rxg+gEzN6vGgXlCbrJwxRT+sOy1Uzl89jCvX19gLyMyDfDlzCX
04SjVystop/khiJxGdYP+XQqYryPmBxB4xrKXqESZUm2q49HZvv35Sooy1leWJi9mq0DEa2WF9hf
OW3931YJ60A3roY/xTRZk/IMJZLaWz1AWRcJEq+e4mine33DNHuRkUBBOzTpmRSorHIG/yMZ4HJU
tlrzyr3xpVas2I6eGag+9IdmHbC5npQxa6EO1EYRZQvqdCkhEhKeyATw51yYMbnRD2YTe5dzQ3tR
xwtIXSC3eQQ/78/mgo8RiEuLbod59hhwUmiU877XKJPXd3QYcJrCC4an84Iy6S8dFkTdgVcYnpdF
nc5M5HpGKf7KQllN5AnvV7ZWd/pC3JXlFKFhSZ3vzF2nEytpljMfF5KpgU5OBB+8KsGWxsD25v1f
Y8kr8cAR5OtK5ZnWwN9sG5JN947mNV3MnfICvvLfD2pUVClwtkZzI4ALJSxYOjtoadG/JfmJtBv6
OKXccisg9+8sg1NN1Rq2ikmp3kfHfvtCs8jH1bfZw++NE68u3/YXzq3zca0SKuSxea2CvNsNq+V1
REoYsBbRn1/2rDLCDdZL+cmqK4SfKTkOI29BC025b11E2h/P+WgljSwZ+v7xqIQks8Wg1WsyxA85
jltippfn6MAkPFYC8tM95DT9Qr5SoVVvIpsMw95VVLdMsm2hxcsbl+CqXOX2Dj2vE9m0I5o9Nn8A
NVHktGlRM3XUyCt1ltTzD3pFWI9JchbZONqzl9Wkr/xXRuX5/gP9oQ07VQGd315x6CAmvjA12N/E
r9zc0ffpTO1rcwd+AqwHVnkD6aI3hfndrCttg1uvzee7l9+YfCowCIByOItJ1yl42QFt6U1SWNpr
581vTPhC0mjHqqxJqhinGf71eceekUSFqz75R2gABa+DbRv36Le66BjROO1UKEKtSZg7tzVjv8uj
3uSYq9iQ1YmXHKoi9/uggiMg/RyjgBgoaCQuxgzruBQ3E3wri9z6iXzJCjG3S9OhrH80miSAP1iF
st0OuKhw1+RTaogtXImIbAjnGsZ4WasKL6o/Os+rZrtSN7nfLh7o6WM4zdxCrDolS7sCFmxtEZbX
HjzTdDrtTO+ZJLklCM4Ua6BvoU/pl7GbykrdwHgnjeOhIN3i5PQgJkDy68Z3UUgTqf1S8KN63lVx
3aLmazrbT5aGQhBn18tiEfhoFrL14sTmGUH/mr3HgjomPakOmD4TX1ox3sMFGyg67SrHhNlNNAkn
bUB4Jq5zkqa6yI9aSCchqUnAPN9owUfSR5kc9FwknwU8rumRQ7zIAGHlonvabpreyVW+fOfXMlsm
SCbXI3ICbFzvmucTKb3XXMAkGGVKMbxFpqfyV1srnxgnkxeOJImh8ySaSEWnUW8qvXExK/JZvXkl
iTAF/SQULC7DePh/XH5CsYQe578cj5J3wije5uOOy59o6qAbGhkzeZVifYlIBqpS0ApNc3k0waSI
aKHSnC0BDJc0m3hExYPXSkSlSn66KJXlVmsSgkyHiaAxwZAPkENPkfIhPqZipn6i1SsFkXdqhMpU
/lFgJc9MPe3zHA4aq5mM3wxdcj/4fdl7hFHHDN7U+7in1Ou0xek64/+aovSwv+RFXMAKanAg1QXv
MS2AXnjSuzLoSqsjEQ7vjL3af1+piCXjdl38ChgRj2tMKwDJvt39j7/61iUs8MRd77nOOJhaddho
TSyG1/MnBR9hGxcwxKWQqjm+rCd6Xq4oNVD6riEVpB248tz9382AYM4qYGe5BhIqmKH30oQOkYTQ
KyG/1h44wrBo3JtM4alMBUjwxCMtCmUmO7Lbj0TyUsyD030QlCvjCHN/iNiXGRKvwaA9/rZBRBAg
DSgYaYiHO03ZXkZT8mOv3s/aODjQOrs9I9xotuBYe4WWknRQonBwt11Sf5Z8tltORmH/svyXo6Li
AmIkABjTVfhUvUltetkTDoiHhhSJSzZ4MjzPgNxqGUGwWovjpy48JBweaNv3tJE62tolcqvC1TJQ
tZvJ4YblJvPx5tBIAZ5prWC6HRimVLEt6GPAEd8BZzAdXiN2Y5gcQwvuJQ/gJ6DfVt740LtCU+7h
UwIcc7/1KtB+29ICaWFJg0vqOq5JYaZ/tQw4H3CRXY9Cp9O+d8HFVf5ItzDzChmUHy3MHAjLCMIP
txQGotji+vg/fY1ZFMa5TQwQRB6E9GBXjFJRvMWh9jJ90Gf5GzqH+WUNPjJyV2a5nk4SUKM5o8qH
3ERqfB3HJUYJSDUxSoNgU33myMms25yxPaWUc0xxXRMU4FN/7kxxYTh7Go+eLV/TKWgFje0po94d
UDIP6cX6vdWD73qXJwQvtKMRbVEEwb/zOUbxQFZYMtUvRfZpU0kjT0Uc3vJM1rHwjk2ebeT0iM1Z
y4Nnhun2mlJPsDC/9wCyaMZPZ0kSzaGPSlWLJLU0ccuoA5rJqY966uLN4j9Jy8D8imJMmvF+C1cE
VkXcYWV+/fbmgFfLxs5g+TeGA3FFYpm9D2dHJweSSbpDkm/FWSKJFjfa2p8KuWRVaebLApmGd07a
ZORyxsq6gQGlLX3AzlWLU3skrnLaEWGqwyjg9wo0tJ5padIO+Ahu1biENn7NMoUs3/YqZx1zAeBm
fXz2zYFHLpgQLMI7feuWdMOapq+6Q18GcahSuG4wLiYhDumj3DGjXBPpRiQfxjmvPrseVPyOwko6
7EwT3UyCi0glw062wMUPlTq9OwUDtvr9ol9dF56fmlw6B+ZIgDsubS6I4VrPs93m89JyRHjjRFtS
HtZqDLBDPlPrlqQNBc20s+TGj5ZI3qW2Xx6OliwpyhR0wfTtcIAvzwDlGWYblL1hejpzm0uVUK+f
4BUIexyLzIv0whFGjyHzbM7jiR05XDgdo3HTxvCFVHsZ/WGmF5Vu6dL448Xt4rH5RgL5nhixQD1r
tWQuZYGEihmRuSD4RVFPPBbdvTSXVV8aablFxM+nOG165EGaCGwYQp5mqBvzR/MxizYPSNKtC1Bq
k5FSX91ZiEleTLVmiqU3xRxLUJ1ABlyCbSwvnminqeuiyV4Eaglo7m3awT1UbRhM2DQUeXuoBKPT
yWsUeP4nhmSC5GspPtPm/qVjfqczNTyxSXGBdiL0ytQ42Ep9Hm5Or2TVNpWAx+/pSn7rb/y4VP9y
WNEsNFEWTdICNDX54rxiK6prgG4nMCUccl2VY4OPHT5yWuEQRSEJmaojeIx9AL9d04XwEcBiWGxt
th4LL+xpez2R/Ym+th2oG4gvEZgBkfVJx7Fu9hS1cuh8+gAzjMHiiKM60NRcu4bunBIZ6NsMxePL
aN66qiOihsuJOqsiAeKmYvNkug2mqKZicMl5GjekXwLO6pKFGb/Rg4Wxt62Z3S5FgnLjp0OVthDq
7bCeqtoUfRJfqYu03RrJQR0Q20pu3MjDojz7mH69PPMcnCjyIuGmxxVTlRzalTpMVysQR6rNyNiz
tTmqaNDUly8EbVMIQmFQXXwzqtQlcM6Es7yyhXDDerF7IyzGrvfprUIgBvqGq0msh7KarV5VX7IB
1hWyqBgEM8jRZBxRqpWoV2shzjxFkaSC6bptDwwimoL0RU19KpvepYOXs93a6h5lzx0KPDU2X7sY
tBl/tf0wvV8lhunI4bAKNq05Qs+4fqWUXA0mVJJNEHXSkmlp1waam0srBmsKqJiYiuUCi7xC6VwH
LAKrDfWgDw+qMlJ1KaxNSCniTTzAGHT0NUJP+xF//iOUqTo+Ma77fLkUq0z7IxVukOQ9t4Vgx7wn
FDDi59/5RZsbANk20DddgeoW8ZlPkg/dNleUwnOEekBW7goy0P0D3PO3YwuIj2cXmTRa3pIkVlG4
vEOvciafauJvKZuPTQypEKcXrsETbwaDN2dVUSsDctJZWJIQvv2q7PjThCjwYy33P+r95roloixm
sYCRsWwvDNEr7T9WBnT2LJ8PLTCYtkTHhchDTpsFVrdfbCAxvO1weYcR/Uj92vE4NH6U1rFLBiGM
TjsPnXEQKM6IYjwEZV4LXNXh806M+CC3cj2Zi3MHhPrL8sHirvrvl+q9t+SWtRblFH8jYgc8JY4E
Vq56u0v5KPua69JEDl42hmuKoep8GmqV1Kt43ccQTeBorYZ7EkxE/ObwT1eg4IfZn+Xw5wUmoGea
pyUG9FNdt5Pla/6KkYqizikapEektxDzOa5A884ctfTH9CGXLenWQxQfCdcvFKtJLbU8yrc3MEO7
m7ildKc4MdV6wcGpBcT0t44pBiO00TpHlhuehYR5jqQetMMXC+iOYDA8A0e021A9hyMXOHE0ZQ8j
pNAGoqNWRB3dY6v/WIZFlhShnrKva+SKXIusXr39QkNS7aKlbN6dSZGfRYW8zkpp3PZYS0ZOJMF/
XpxXeX8V91lNJ4HcTGr2pG9Wd1Qys1lGMs6Dh1Qo/U8F/47QxvsBKhcOSS/Darx/SKK4Z6yBKr2Q
8xnVcK9slxSi+l6n5OSx9sM3YiLG9c1JyX9kn3YaZPhJlqq8K146CNaKViZlUExl+TsxN3CElLa9
oY0zeeUQBrVGoJ67iWG/8aqMhf1SSRhcWDYTyIL0UgZhSZ4BtNSOnT/XyKueEZyojcvVhn6YzQTV
N8lmwJlZV6sU+J8OGyrQgVMCuSgepoCycTfH39bH7weqkZJrJzdIDWI2r+N9gweMdc5NhLWkzWLq
i4g6voEGKNJL55CHZUGrJ42DkdYZpeQoUtxU5zGg5I4TZOUvqhN30WOCMF4K1Vd6GFXJBmEwtNK2
+GUK8ogs9GHkHmVzvBflRQ5QL4y0VmaRhMZLfhmNyMRD7YveTR0zlFCdrjGtuNiHq54U41iRJ8LN
cY7McxQK89oWvYSrUIg5HTbE5DyOh47kRo3AqJ/d4yABy9tkXNAeC/tlRpurA6GHs6YM/xdDq521
Iva+AlkalqNypvyor4IAmJ8Ckzf5/kk+6Ftp55pJn0wYArMPo0no9ywTwHeQMQyqpLJRFdoEua1f
E52omZJI2r9aoVZ60VjuAj4iZ9GPv6PHbhvc9+naC1xWDdxcBIcZDLwTNI+U71DDFCIeSoJPm6kT
jdn9Wr9GEPVBj4RJBUBgHVxD9tJg8u/2BsHIIuv9dUdtB0Cl0JFvsaWrnEqXB/ql+vcvA0KvZy2D
s7Y6UMa0c2mAcpoRtmG8DlGePhcMDWYTiCdzOvJcibFX1Hq7SdMdegQy8SkQgmHJLWTAJ2adpDqb
YLqTt9ylPNCjNMqS5YSWWrWftl6Mo0XxzNEsuyOIupqvVsnHHSapM1PbHimPCQXyIOE6dnV6tnUV
yh04KZCSFXsGLMMsD2ITeo2o0tOCMOcoxHDMT1yjz83TElOF8TIM9YH2sFdLRLYrWG+AGXIHnAEY
k6oSlPcYhN73hAdLiKR4QilHG8zkCa3+dydSSxd5Qb9vwv87FHfRwLSynC+mXr/JjwvFiCYqpyMY
bshMUw9CHbZdFnWUh+o8IyNwQ9PMYiRSzbotLsZSEN0BqQO3iYDUz1LIFa9vxyS2Ix5rvQ1W2Lf2
56tsPi2ow63uDB0NdpRmT3YUx29HNoTOL+FYi3QHgqN0ncpVwTmbsn+4K6yM3ifyCU+DYvYjouK+
5gIfDlYxYP3ijUYt2c5ad6PSwZd03zkP/3luTgJh8AEIboWctR+yC1IB4vjzvXjCSBs1YZBJqAQ8
KPGrsnbMzwn7xA7uUoqCrlNUk78osS7fTE6s5XloUV1DM6rLoRIYkqhE5AMLymUDN2phBlUAboq6
cB9PKSxVKyM/7p8NGiUBHYIgQQ1iREoa3fzOg2KBsN+k/j8YO7qdX0q4JrHa/TWDePtxbw7ywH2R
hlKvs0C84Au3ZekhfqekPMS08gu3sK5Y4F2Jq7Yz1MNdqHaROW8NtXfpuSh28vWFP4/pR+P79PdN
+2jV9TaNpvqOnf28hCfnIpfcly1Hmi5ChlFbPwAkgWa2cST+rnBGH206ZQmTLH9kGkKpNBzKQt67
Dg+l2rRO2yHd11HHlz4yf8RS33l3+ETsfKsj775+vp5Ow38DtlTMUbaUSs1raUFXkRGLk99XfAZz
WsNXJ4dZz0hW+OTzjfiBniyW99P/ZdiPfgQtOmn3MxfTif1zHqXtaaMpj4MTxmHBjsfHwogk5PX0
czlXgC/9dEbgzejib6VRmaf+PSgCley2lRR+qL4HeMb3Vk64I4XmwQnph+MvcRyisZc7B6IjZnqY
TGiyjqDtpdvUsYRSDx3uwJqDnLI66nDEEvXIyitVtbysbzq323sUPrQhRR2cCCJ4BV9EEyweB474
u7Aav2QUzKmGtHL7mVjJCxmXu6Y3a4xuKgiBGxFLOK+13Vs1s7EPCPOJz+F6z7j3frLiUGlathU6
Ereou1rdHVhYdyd/ZnAa0Sl+vnMhDV4IWSptYodjL33c7Jv4s4z+CPa/5FUdDhpdvjvSL47wBn9Q
pf85+9WaijEe2S6Kl1JAwzojZDDdKfaAGvd26lEe98IwvLTGHx3sGckMA7JA5b5g9vqgSVCF5vi4
lrEnqu6YasXg9X3OXA+5e7vBz3AXbIQ1z+z7jJ2fOcemwrhq/i6bC/HLdaWk16b4ZOuTVpejnbIA
ej9Y/hJzfSDUl1R5+8eekuxMNMc5RCdYVamVFkiGcqJSrOafmuuBsq0TT4Is3tIXquDhNXGnw8hJ
kYbCEVCfRiFBzYo1cThLTaIdBcVblqZ/7o5tjQqZAXSi7bPOYQ5vGaxHHQBS9mwKSSjr4yap4zVa
NMVjtgDqAhUjEl0sY8Xdsgwvhu7HAFpSdBNqL9PpZslysmfDcMvBW9w9l7I4pee/AA7yv/0y1tNK
akyq8uO2o4F3GPPl4kJCndqbVXWNYe4vciJMPk+ClSRm5Pbv4gKPfLacbH9NePMdnR2MYwWKD0wM
NLpX887neYMsgSTDB0IAopLlNc3n5XG84Tu83JUoHz7PfVxlx7JG4HdZ+g/x3h9roOA+m8NDGHdk
3wwffBaJsT13MzuUnINlRFam7UWxUg4hPden9945C7+zuCefKtHW1GY7mDzqHWKRD3SVDoUIh2k1
vDGD3GVb23mDykmRelSfGwxMokt48EQMerznmmdCGrk+IkKV6l8D2MzQz+yfVxs8h++dGa5BAwsJ
gcs4g8tKyHU7+oPHaChxdInRLSddr3rE+cp5SSbvtsurLUVh7iYUEHb2JL+fsT6+rx/Ly8/N40v2
nVhdIgVl5lbdsMjaQVsiWekkwUOEjab216uv98DLZ/dENI2GRXdfv/J3qCXfzc4fFNr79/1I6/D+
hQTSexB3/1MMQObX7+Nntr2G2zORTzdDM1DNrYtCJ+7YBry2KIPFYq55e+nB1poL7XJfr5c3Nv11
vVik30aa9RmEQ4rR4qSwKZGiFrffWkFPDSr+PGUBSrErT+Qujzp3kW6rS7vflQx6GAsBBs6/yFuT
X/db3G6FUN7Vvl69+hzrM2M/8RL/lk+xAp5Qx0K78iODR00XjUNZJmV7WQpxII65ahsU+ByDt+vf
j+XEVb1J9dibDuUmWIYRcKOuqrIRW7vSxXpfQn4dsNpyWfFQSDNoSRmM8Q3xVgXA198IR46EFGu+
DixQ/TTw+ME1mZyuwSCYJdEz970UazVYOCtKeH2XI34kthYAYkrwm9UGYKFXiKbmyUNI4T1gTGaG
8nU/ZnFShQX7z/MMeiNw04srvpbA5JuVgaL7HzyWj7IJKQ5baCgC4WfjIWGTt/65ZDHeegcinRR6
rzq51JmWTioWWilNNARvJMqcB2kqACie2fBWskTirM8a3G+66Jzq7WO0pr6e2IZV1OcOjK4dY/n5
o8QcDOucUTK4STBaHjY4AoVZTrilDnPAgQECoHpuTNGnkqny8uRkpkdcTDGO30mBGBTAhwZ0Dwdw
Cab6OtDjhrvENkYN0D6Ti4urzgkcguARniWFN0/9HG4RRLMc0HOKIqRhWRLFqi36aQaM051GjyuN
M+hB5O1x4tRKK+1NrR8G5tXVKQ2hMXhA+8q06lZ/4HRjagWZ96t9vuq95NVtJeFzQ10I8BwnXnqf
f1a4EwEhcoMHibp0lj25uOc3G7IZdaW3PGggzYjTAWiMmLD9g++VVwkUrQzctiSfB1CCecShdDrH
BFhFBMJ71Mjhb1KUNCkUvDsME3GGPzA+ncI9KHNBDmp0zttzoZsXzJkl8ZvjZMXP1s4DLITKSe7T
uio+hVty10ZjaX/XXXf4FPn8oIvVBeBjKpUC5/4nE063ksfViZCOXfM8bXVpJ4ygqnxeVNCYcnew
B1ysG88BcYaS+1sdNJOvmRXHrKEaa3xE6qBJ8/ZflnsN3qZ7gzz+XDWRY556CvNh4sVZ14a0D0R9
glrfbhB+TE1zAPCIkFCEd4+sufbR0d4aCm+GCPRxeuRJNUkgm2UbVxBKVG0G7Pt3MwXF+0d78fMX
chOXigSHTkH5Js8B6wcl2KfzOrk37WI2PVKhxut2gAw4dBe9psSijwkka27dAG/s5tm6nkh+/Wpd
SBRySMRmcQ8uZn5NySban2wV8XqfQ+wXoGHx6OBxRKHMbFg8jc+Aulkq/BXl5o3E8KD98UBKpTXp
amkcQ+vfqsbBqtzDKgpGU5pi7N5jYXwn3BDpXmx6jXXmcDzko+XbYGLBonuSASJ7Uft2hrfJWqrn
fd4zz8P6wgK73G9Fh92UiIHYlqHtbZyFoOPpFHzvAsAaf/UBCmcEeZ2xDP/n7O9aeerTOw3hkWDV
8OkhK9hDjhuJmVD1qntOt4FxBu7mOvikK9E5WSSsNauHYzj7/q6A8EWkkk3wxRijxjT3D68qIo8p
y/eVQvlMBUWCUvbhzLM4uuDsj9gR4ZsVlThnVHORLkJoAczI1ctifXgKH0tj6ztfO3DTE34dKWUC
AiQjbpo7RptM/x9d+Y36Cf9LzsvPvI4uE7rGbFoSF1d1odTq8j9BHGAZEKj3M5a67HQVVE7+hFyA
12cNIzL4XfCAXJg2iXGK20W61NF69K5YfvVGEXr4Y15G2TRyWaD2mNaAPZEsbPyIuaUGIyeS3TDZ
u94d1pWQTfRPrB6pbEjajEYKOEivDxqiI//GIzGxHXyPC1iSjoSGNJl/J0fyzhO8iCq++Xl/YgmC
nOsAr+1gf7LeFwkDE5L7dUJrwhJzY5hKEu0ey5S8hFTh7jsWNbpaWIxVlUPybWjB8QfXqVN4clsg
xJekehlO63n/VmzVFfOUZJ1+23NnicwQ+j+T6MVTqd7NKl6cOwDoWpkTH1unjfrVUykhLnX0NCkI
j59s6RUWs41VFVn561bmV+I7wmAngfrseoW8UqHhXWfXqmL4j5aNic3Q/5zFu2rRVH4kVmktAmWy
KjWcudME7yinwVw0/rdyoSokgWzW0k3eQTspXCGd6YkZvpzdJTs3cDabigO9tWMLZq03wx2/8dqo
mFKjcoi65vB7fISAfzP0yvQ/ucfAUojlFhICyuMZqj8LEA6UlV+OpHTO3hCg7sBoPJMM9x2XGiF+
BIUIR3coyHcRgeXqcT/Ist9kxzl24Lhdc0/7cLb6MbFxDYQTK1913KPH5VOhtoOHU59Nwblq4sdq
4GiHL4avQRAeFi7rIsq52zyNXTB1aSUmX9/W7vmOg44LdXwUAXpuyZ4YGONlqWkbOKPl9JTm1tkl
9WvRZxZ5AuFYUXYusVfwDZoyGhgWOh34Hc1Imo5C0IXWwf6uE1NrW2zTqrCMGFtwLzvddcdg94gh
mgRvmDbWxgUx2qSH7i0mKwVwI7HWwP8SRn/anych43VCnsPvxGOOuYABruC9kMKCiZ1FeC+RiLIa
oDILD2o3zJ2eG61BnyLW+KHIXmWzyh6z8476AM4HB/eyCp3UbIDWI7wA4OX+AyLC3OKf5EsTLHJK
oM2wAiO/bqhMID+Ol8uw/iJ2JP2kBP+NcGWOm+ZSGOdmCFpISF9PZw8mBUi5Em+y01WR/EnJSCNT
RQ91beNAOT2pNKEjEyEh97MNr7PbzMW8QZj/p/Coi6cFnD+2cR3poxwQwc/RFoX85+K/+i1zT6Nr
WXLaaEEIlSwG7Zl0TaRqTVJry04h+IYEbg21AjTgHjszwFafapqTyC/VaEgGUEzfjn38MTjEUGoN
mWvSXw5RGFKSUdYXSxAnyb7vhr8XHZKg7XqRzpyTSfZS9ts9A9VAUK0vfAuLPpFcqhh7lkiZzrUg
YwvGwjkdaS622jjGnaUANSTi9Mwwb90Y1lrzQ2wa8l5/9FUAY186qLSM0+LOMyPSwUesHOTw8YPP
NUUIQ1ksyCO/tcsvXvBy0+EWzdVqgHgY3U8kKWqCVLzTA9jYapPmAd5UJvQLzvAdXVE9HmL+c52y
XunyDeydL0NAjK4UOxRtpSdEFUDT9EsZMh9+KucZVlIfhY/C4a8wLs0pb6AlujpJUlp1/IFU8M37
BZL8zZpi4ZQfJzN6soVhFwng/BfZlwboi02PyitFyUSR1vq6tCMwfDSDd62NkJhsqwHF3tXpY7t9
xqzWrFSfVMtta3tDRpiMrxFfptqNl2x6nEJflWTOPzb4YQK81LXygIXwteVSCx1GVn20KkkTySsT
lqVbkWQ9FeNGoYuQ9wArkpMolteEAfHEQoLixhg4I3/n3FmDAwSBACGXCqMUpOqdw6PaqHmMFhju
R2c5f4UCoy0pemR6SAPji0s/iKGhpJW7AAzrNqaZvmRXve7Ve6XflE262Uo2AsFBJlk7TI+cnKWn
SHELUwicgTfH+U5xbdMBtkKkK06b0RuTVNS7XZ5NhQFUqifvwC1md3/k13X/oye62ZAVbZLp2QQ6
wESE7nVvnnhSAvo4flTBzwFGnd0/zON+dLEWbNz54G+OzmjXLgPLgobj5v8MPJm0okH3jrlDOdaZ
iO3b76IIeObDFeUyGqtrxhVex3Gw4xvoMQ3etbyKG5lpYGcS1Nud1dtHJoSMNzRjL7MyVxkR9vZd
1iKnLXZVmyWpKzm63GgSnjEEYqqByYVkn3g/sHHytruiu1U/SwIohnydro8TDDgCT96romEAwXB3
cZfQJPyPNuONMoNC1zk9o5WE8alvxWGoRSWrkF+G69NyH61GFKsIFI/GINz5JC8HI4RqeEG9Hvse
6jCj1Pcrtw54pN0B/NNKg6byEg3/da1rF7n7aalBYkIHCFmY4quvdyNKY54ctTSTbpkJJvdFON+B
R3k1/Cf4T9hMRf5VJhgT+uPxvRvK8rrOmMLmjVj0wgsIuhCxOEe5LdyQtt3PSxXwMHMiUQRW9Tux
Uy7lhPoXjIp30aQVzO0itLp6vj8kT10AaXlHvYrltaq6Nb88XvBKLKPQhtywsQ64a/tkhm4dnHkn
CuUxuClnnlaskgkDZfoh5/XQibIFlqzHAsgpO7om3VDMwmVIsOstv1pRMBlmsqLWf+DqRR08RgN1
d7ppB1tAXEbuUkQZJasYZkIs5RbXq3c9RLek4HDnHuoGtQtYTINkIlrQp5qliX6zBB+hlCM4E845
4frBnLhccqodZbctW4LcvRmH+kLNrSiwBeVa/RKJnU1B7kHZ5XoRFEoOCeHwmyspLFwFbTQxBSXp
sNF3srmEkJPes2JBpJzgqL1XuahOfYWqdxXTkIcVf5936KNbPNYlAeefmWrWyhEAaQJfbd3uU2mP
n5plASbIxWO1hTsnnFljOEsA44NmGfEn3EXRFb0f2fN0yldzSDcjPkFyU2x2xAcnTHe16qGMqMcx
7g54NDml/QGyzdHW5b6Xy9w3fD8AdL1srp/yO8x3Udw8f+d2k7f1CYmCJjzExQAb7P80A8z/5khK
gme4FAtlpPDURhAQ/8q5rtRCPrWcGTD4PWJeo11lQJeWbSTm8fRRddgCuL7zUb2ZxFzBpbCA5Wge
F++QM8Fu3CVXw7Jfl4x5qmX9MHrfegHCiIVWKs/5jg5Vi9uIKFlay8XWdQcxcYvXEe9qA0LJzdFi
oqIPCd5hdv5pTiZ/KFs3DnIygXYGVuPsKQzOkRql+GmWUapKpDEI0wsTCEXpavIi/nrE3w/mwpaM
VCcoxkdSWfdo18+6y5EF++WTUil0kdF2seIDhA4On20LAQ0gZmLAnafcusWEOHoW9T+l9LHk1mdf
6LCs3JTfoFO/rvCajNzuR80wgMGH3XdPOM/VfZzz6CIRGJdYmJPLywUOMRxlhy1T30rQov3CCsJr
WremzCGmGMVQL1OApKV2QtpgKCzEQ7114drnP1iT/Fhbrhm5m/0GqZDFMBWNgAP9biY1FHelS3WA
bSQWOz518GfT3gcC6k4OscycI7jqX0dQmNsSjbGU5+anyPEB8YUu1tEVWQDCkjJxn8p2GbCpqwvQ
4BxJI5FCvVqnuwisdcp8irqR+ejCr71BYvGZv2R1ahymQXA4FoNvsvMZd7Rjf3J/HBdLimwKYqlq
/z0J9kr/4eCM/SQLul/Y4F8dB6TEbUtkpyCQVr07FR1PDkAAYCNMv8hdxWwU1+W2waj4J5TgZG+x
jP3vsM7vAW9SNrqFAPXwAJzYUSxbseyfkt/c09mRzkID6GJwR/z75SaOS4kgohF+BetC0be9Bs5K
Gvb2b6+u/OcTkGcYC6HzdwONb277fVzr646I1LcsUgfjF/1tQk6D7UqUZZdiGtsc6xCYfPisRXu7
yoxuekXvtuSslI3WQe4aGSG+br4eLPMnPERfXEvBjhDf9kViHJjkIrQqkA2re4ohQi2T1gMNU1dP
mOfh7/NnW7u4f5pJ/jSPfI3YSa7leYD94meZ3y2jEDKGATisUFZNHBwkhuW31oVZillmg6Q2X9Py
uLJ+e9dBY0BHQWBbiLxan4vKRHkIJhyPepMWIcZxLMJYebzlrGM4AaF41LjnIH7K7pw285kbZ+fk
IOmIBoruiTaWH5rxa/W3YaoVy8dRMNcJFnPLsv9P/IL4V6ImHMOBUZ/TbO9zFDMSgUj1Sxu3xnSr
aWWlu3oNErQSIa01v53DisgOEHSJfVR65u2NFF9O3R6xlEr7F9zCUEvCFrbtL4eAkKgiSvtiLOHY
TXCqyFT1QLlT0Uorvft/RzYxDN+Cdy7n63aOVK+w4a6pd/k+eLRBzfcc6ZKLVSqLYH9jLO1f1+/U
TQM9oQD9Y1WkryFeoHCq2uBtIEYa1Qn/UBYgO4ZOniaTRWg1ld1/FXMCamT1WOXQQ+sbYb4EgsjV
8jUNsNyyI2mPj9xCJ4m1+/d/TE8tCQ/voqI1lSMCHOmWSIZme1WzaKWsEnTrJF8TdONx1tLff/t9
R047Rz+KSsI6GTB2ZIusY39DiqO6TnJ2wlLxViuZfA4inWJ6e7Qh5hpegegTvr5kJLb59Tm2r7aE
zlib57mmoOR/N2v3AsAVcvcxEH8W0NTv2rRHqDYml/Rc4aqboTg+XVyZ7Xv9ZnoEVwEIr8Lbhz/P
pawd6ovjQMKdm5lJMdhv+uioeC++BY3TvYCT3CyOxSe4HlCANxruqxtKuQBh9N0IfGc25bxSF53y
ID9YdJNQgWzNmimcmVIt86WsKbWPU/zmlF8fYInOaD2lzWilfnDvPYRoPYhqOqPD39ru+oPC8t0s
OjcwnAdAlZv1Mni/YjDKfd91rLJ29X40Uv+YViZsLreWUO2ysX+3jepISp6lm8Wfi/XFWEalCOEY
VbgnqbewNZOzJy9WBsnZziGXGBctd+7QoSaZsml+zXe71apsiU1z8ozNw81Q/eITVLDBBGJEb/VN
HwMTAaMuxT7bY+bs015DtXPfKmNrYa6ePNU4OtsOKOtBKSvzwFklX9YFDy8u1aI8p1b5zXwfLLTh
A/RKnWOfCh1gsC5OiS5uEkQCJjAL5qNBYCS5rmjF742RbUwOg/qwND1or++Vm9QzQ8HbPkh1/gKC
SxUseQ45xeqIJwqU3alppImKhxRLovpkcNBlJrXio/TDQaAimEq+hNraNIWLiKI1L6eu6kyaLtkZ
FK0U4jMcOYYoSjrfA8X6ejWu3UBNmDWm2jvLZ6NF2NsDYq52tMG2h5FDwjl/O1SNHpf40fS9O0yr
mDRqIxINjty8CqGkaLFQdzerpupybM8CBAUZCDUFG2SFbVrMHYNCbFIMskSRn/7Jp3q7yuwokn3U
GoaK4/Dtc/SZAW0qbelWMU/u4TpdQxm4DYw4Svsy6IJSkEzsiVkDTGrE9OaikjWiuhhaHVfzDaEF
mkFaziWkReplhClgTOrVAaou1V7SMsHnPTn4uM7q4b34YtkHHDikpa3axYZsDLOLHsAsfVfL51/q
oEaZ9o/LONWfXwVFZX5vbKG5v14i/X2QfbczVPYK6jhye0vCgNC613VfwIdUEK1rt72Mev7mcTpY
yK6ik05qSZfMTdsLVbJtEtW4u2QfACWVYfzihA07FYHZuzZE0Opqw5+qGHcSnUB/b1XOJMixUiRx
EydUOSY2wJzM6dIv0YB9hGCrpDUwIyrF4KuJVakmz3rXOdg/XQxS5BToJX/bAspy96Bu2gd051h3
hi+9O1rz3AHi6SQzOMmKXi4czmY3yhEua/fDgH/8aOJgp/IPeh9b8mtTxPzagCTxz1TCTMn5/L6T
e5Woqh0r7lurDTo4FvJuzfqdLE+orZ5uwtjF4pBFCU4pGdgDwsMZbmCCZwBoQWhFU6wt9UVP1Sr+
Ac8uETSQ/XAAIwr7mFzDID7cH8GrtyF81O9zzsRVvGyMiGRlWhznNGzuovm8LpdjVE3traup4qLe
OoKmYPqh49AIUWFUvdlBunden1vPDP9QI4x1icS9VXKQyYsaOoQ9UxtfDMILAIBjtmLY2x/akYnq
IMzrC/MeJbpJJSbNaE7vTbuq/kITGIYKCjaIsqqDUO3aMbUeWPZittM8l2DUS3K5ZBn70BpbkLAL
XXKPkGo+EiVSD2Q7FgA0eTVbjoqgm9ih9ke27OVpxJaED7kZEWs4PZTfoeIuCFzO4lthx0WwJ9Sw
AaW0I7kDamc5xqveAZkbqrOMBqXmcshfBC6GQWUHBypvez4ffWi33d5Pj+S2yAkZCNpUdcAFo01x
gz7DCPUac6Ku3is4sTrjoflvhxYONtO02l4fYojnNJG63XHBgZGIxV9Ow5wUMkwAtHqBdOuy36Xp
QBOcEOqei9V6A/BuyA3WX03EqJvxaeKT2JtryUsEFF55Fb+bxInl+CCmef3mP4EE/N5wjaOd9+Dv
49DiatUlVlsW0CKhAtNAB5LigP/HJEY4h38Hv4nqTP6bzctj8Wk/EaFbDK3HDMldei26DLx+h/Y7
kZE9+sc0UtBH7BlbyXR102XfJ2jXvBbxe6xrnfpdig6Gz3Ge8mxU328aPiFtS/nsOXq9ikNFEXYO
Wbz/K7cQ5sRrLHmZBDdNkvcPK9XMd4K/GWS55WVG3oWnO+19gqVnulP6UEKzePobFb1nk6v914I/
0MUqJVI5ztEcNO9XmbsPQ120NZH4ZN5fkbEMN++zj+Y6I+6UKjzfwvduXoWdyVedLGPNsZDVp/NW
eGPAUKTCL20uk/uHQk/Ol5NEZAgNKiBfzc9NRS0pzwa+0q3X6DFErdbBWBNp0B/QVN5iGpLEntPW
uygfiX22dQ4HWzfNqH1Sc5vvM4xJRCntnz8xLxUx/WeYANRzbXax4OHPYLO9q+rxbhDjcfjR1gKG
oN9TFYK3jb0OiGpWljfUj3EngBZcF5RQrAdVXb6GJlNLUKQVgB/Tx/PkSp8GsCsG0NJeyW1JiOB0
1BzaMedl5M8ikLkkZW9Ze9aW8Y4BEQbi6oH6Z83zBz3q9MehQPfM35qqSnNhRbSTnkMnJx/2Zwl0
QnTh8ZlL2C4wAz8xZ2/JN724A00iyWSM6yv+lCrLnypJtfTXGfOV3qQ0YgtVGLtt6i++OUdj7pxG
0aH5I6wuJu/6k+JkJ+ptmqJeSgJ7Osczq4QtNImJlaUgCKYv1auSsRV49un1il+WsxJe3uCJ3hQZ
SfyvEdGu7UlHuALL0RWUNByeH+rlfxv4VWjgFVQPXU0xsBKv/Axc5ucVGqLVzgLXfNr3RI1rt5sL
rDSuOmxe3VtVR8dJAVG4LssWDSP4a+q7+HsQCHZWp0837on+NA2bwe2MSgrbaH9DlyYEKOBHGvxH
7me2XfGPF7aaUrSMSNsRfkz5ZLcfdFq76kpmAgmSb6rhJiZeUS1QroLyX85RRJNSk4fDVXNZr/b2
TaEw3h/F8HHJSdG2IzmDscjQNJEp9kblGYuzXHs/iIUuE61amKAy1byoJZFnHJTo+lJ1Xd82iJni
cNyk6A0Eip5S+y0EkgDQiaOhM8eO9hyxjHaLx4VhnTiZzyqJw9bj/yPjfR0C3I/a+bYR/05/3bGO
4ijJlY/Evs5uJm1Tac1Pt+IhonLWj/45qmNIuipDFZ5FHgClH/oKA15Xmkb324XQMj4HT4IxH2ks
Lhn5xQNNGHR2+qOsLzQ0vr+Q8Fne6LBKLxYtIXnMUK0sS7BRGkcY5YTr85WkLdSouskfJydI5jRm
p33lLiQX3HZOykbhfUkbf+G+Dwt+lkE7XAPBHrJ9r0F5xIRs/b9Z6o6C5ZMjhSSutktERVH7Dtji
nikc48K7m0XXxaHVYhaZ/m70PwPc0cYsDIYw7OmuaKg/lqNXPXojY1EpancrCWfa6AZYSSn3iJPe
WiQpQ5sLR/2uw3VtZQUe/uXppAxEDfbBVbvUT9vQoyjT2GLZpPVa2mtTz1y9HDzxD6npswWLWWuX
xrxPPOlb6RCME8RkfdQrLB7ssT2PN4Hra3N85kv3YNMefTxaGry0zCOv7JaX+Iz4cRoNgEHyqZQ3
ZLtBO12I4sWp3vzEvoQgN5fWi3+NWlEbTch0ZbrjFLoyHwIK6G6m/f78LDyR6aS7MB5mLwchD+w9
oF5oNhiX0P0/Ykgisi9vEi+aLWyDwPaibqQKOhAweFSxZQE7zZo++GqX40CTX++m+KjE7OJE1UwC
CW/1cp8wGP9EqExVm7Sqhly3umJOZ2yyCTQFyd8mgMIlmcm2BHY839rlsl5eKYAcjTzuZM75tiMo
VqmLyVI0Y9feiARj2Ph00AN9q17YVCG+b+9p6rMBf0cb9MUBlRD0knXCthiOgP6XkEbUs/BHZhhE
RLjGEWPNdiDORYb/b9TV8Vf1URmYgC7kNynzQ3Gu9baWJL9jlcMcWU1IWR17xfNn/ZO3ZKTlWCFg
GqlibVL5zjSPc3ENPYAsmJF4suRcwrvFr4FpGOobhW0JyuphVHcvWp2q1AZUjB3mOp27Hwjn5Owy
NCdzQOnOeIicdrMFhG/X0bnrnl9vTxTcY7GbETifdTiPeHxehwV6+wFzYgvzJ+Ze6f7LVi753AEQ
pVUOOh6pOzci9en0g+Vfs1mz/YpL4m7GyVGQWiBcFICkqJsRmxp5LEh5ReDJQ8W2RCGGaJ9rjh1z
FVqGBCwCoiI8HVnEUxdlvbNq+TSd5I4puu6typt7bDSh17GuzEOV0ze4Fqa5M0ZvYSqUtXKCxGum
f2JnHbIGWp32cMqJx9X5g7k21dKmP8965+8as88umfNC84mf20enN3tEpRf3Jmmyk1V9QlB/MBxp
tAHvyO2i0GlJDP7Rx74GkbJxnRrecFLT94HQpXWnBzER/NmJ9ImN3w7bg1g/BNmqGUPbOJcAA1HX
ujAyxA21yPfAACdJRY77DfgO/jiNThp0r7k1N1UwWHvqw8Ey4VNo4QuEXI2WonP2Gb+QjYAJTcqr
j81q4aFd3BD6tGSuCBfiRxyZVKM4RD5JAzK59P8ChkE+2VfY24+xTUctntvnvPWUaH7yNYk5XItw
P+cNOzlsAGGF+7mSr8g5ApDZxieVOuYetTYlGD2lYP0zc4VVi4gOyuChI+EDMbbIxtft49RsUj+J
9tAJw734lxG/McoJcL1OAyJNZPNBpI+pjf9Dycr9gTLSlfoKeddhMtJU/S3f9NTTOf6iIJzDV3GP
YwZUFABnkge8X2B2Ky1fg145U38NEOrkEeHVEMk/Ifl4MkKQnxobCEtyjT9lch0xVZhRQcSjo8vb
lhoTGibI4PXpnBNbd4gPcNbwUQZ//gnS5AdheAi9fmJRS7NX6GI4KtpxXgHhd0I67rgarNcNVmOC
AlGeKT9iyg9oZ0Tk65ZDu28Z9LVCkUMT5rF7uTP9aOae4YVivSoBqJv41nPXjKPOJ5KhgE8mCqaF
zSFvSA8XfNJr4rpLw6zB4IgZmeX9DOhnczwxiKUzh75J/e7/E6VLl7etYUgjgRVyBxG52eRGJ9KO
j/Y72SIl3iamCJasO8NLMk3V5zBAKfjzaTsockJUZrKp8Cei0U4Ay7dpkCxmxNVom1sr8dgzHzVf
C46Wu2TQZWwizkFA9keVZnWf4/F7xlwXssnr580BzEfczA1eqRkdWTJF0CVhQDtsil/cZ3B2Qt/m
HtNt6QujSxdKXXIGg1T5onV02eqfxIAvwEbMGD2lIKlN2lgiIRydSXRy8sGif4EqiGrHVxoD7ymL
UtlzxmdU9qpYC7kpB8fBN7HhYXR3GtXuThN7FULhSrgZNiC533SGvoTPtor4mb6KVWrd/+2R7/Lo
8S8el/WKH33ODpRjkwja6iI4jxw1APIL81sBET2Sl/3p28KeybCxUFlsTWlbgQblEu/AulWKtMbt
9qdMkyMiCr6j9pRMZXxmVWWYRrcEEejt9MSo5pAToNsoV8nmGNadwvqsftV+QiXf2NyhjxnLg3tx
RRxD56NPVJ5CxE5cud6YVucbgY+x6OKzxgezyKPryOvuEE636v1JaggDApo9aBItwWJXwZfNPv7L
sLXa5KZOZ2CzZtPHx4Q/G1F+w2P2f8pu0m7ImD8BVLqF1V5KUApBMAfb/rq8Ae8p4/KL5xdkJtCN
f71IibgoolpVVbXk68JZm9/AO3lFBu0Ujkqv0SzuZiUZAfwPtan1EYbLVhMjCHbwvnjEafGnxkZG
XMHJ3KbYJxPiEUrPMWkOG2FiQDrPIlIBP5B4d2GcPXC+NJJKwqo8x2l0CU0uQ1cG8L3DaSoHS1cK
rlXC/z9Gz/b+9kuqS8N/5SADMMwz/QutDp+Sv4UIekmewjVMsEaJQ8hA7fweSIJquVJ7F4rJWaH0
eowL3O+NEI9WMymzycRWvUlrzSXwpiCwrf5aQSzuo0Hd+QHFi0+Btcm7y75eUEpmiYW0gTFfp4ps
rzmD7brqv2vfd78S1CiNaJpudhHieAZFBowtWTZ6wj57dnVPA4xj1nKnnVqtrNO9a6RrBN1r3BJZ
DGoQXJjrlF9Mwuz1OWq2F+S5IooMdqnofZPjNHjJfUxpQ4KpeMIvjDklnTA3tlWDCC+abfwQNLBI
+Yvi0+q628ryfAfYtF8z94WrNH6Ez21R3MotzzHrOMc/4A+xyuBv8HxamjKlUo5bOpdgAX5/UFKv
91k9CtyYeInqyJfBuuDVjTFFxEjvoBsW5nJ7/gPwI/UeDpv/O7//fzxC4ao62BPQAXSOGN24UXgJ
W3zq1FV/kHGr0FBzHWbPvGgLjFfupZI3uYy1vBE5v4ToMEGPtoz/7Gyjm2/845JdT81zb23gRO7m
bStcVX3/N3c6slzSqKgFOkSA4D26Ju9o7XSJVgXPNhDvbOUxfHMd/clfXGZQwixfEyT2uzExj0Ss
1wFEifFQW0/6mNZqQFlcQtnC8XD9x2b1madMLN7L7Zh89d10eXk/1DxNEGKXvHmubhuobZKlbeW8
29Ilfiy1QS3652UMtki8Mzql+1MaFzLFQ6QDqV6SGxOMVE9v9YxtCwG8IEYctJez0N0rqoWp3Tzu
3DfaaSY1AvgeWDmplA2YhcgyQQbRcLnD6xdg3bUNCMec3bRgkceDcMMDTZK+evdmozU8QiLer8fO
c+FPo5IB73DQGzvhLszyLuIeLu0KiZopET2rsIySt+ek4viInOI4aG8lt1YmqoOO6xATgBq1pm5b
s6sYX3WGnY66kNiM+YRInm+j3zzW39po8UgyaGCxZEXsWnx014YSAyLxABXN8pPat+UO1e8WSvIe
EAhcxkoMeuaEKHoZULBpHKnPf1lnIfikiKCr7DUk5ztIdyviT8cO40a4urIdYFeFFwrgADUySRly
AO5ngypY91VqC4RXW/V1S9dPukiWajtLMx/cj7+smQHNYO5V5o0cxyC7yCj4w9z4SxJY4qomjsl8
c/dunPNGNK2I1tyHX/7OtpORq3xfepLNdYSjCqQdNcn0W7snECrPmS+zClbhcFIbujBMVQL0H2+6
sEornAh87ArHz7FigYbbm5R5SxjzAA++gGVRMoj1pqJ6yKNCPi1ms9G2KtjZk4l9Qa2LdbmCdoVX
tS5W1MpoycmuAG+TO9Ln0ue94tPoo91THwWqEmOQn1PKkSWQlutEgP1tEW7Q0wPVWXeYeNB2sVwq
upFqp9eL5cEt4ut72RxNUDnRNZ+K/HSJ7qQTn6jjQYkipqs7Gd0lfSeFxibNkPRPa8RncA73ec+A
eAWfEQFHBYBsA6V33yq6uJok1A1APh8jtz7rrj0G6U9aRWsjGCPWYjb+10e8hBUmZzuztcJXCbdZ
TuY0KShNAIUINTWgMcbxQJuCf2/ZQRfzEsXLL3ocEJruffE/4Aok/FjXBuR+qNCqqPWijAqLjxOA
47kDkemp5JzlUApKul1n9lYpUvO9ZTIAdRMMuK0AzW23h714gehpu7XojkTs0wdCFs6GcKgE5cGt
Ko4haO/YXUS2bajoIhtVQ9xNbzZ4dBVyy9gDJ2FMtozp38xZ1d07Y2pRhFBJO0QsFYevmXkn7TkD
GB00r0MN5jCJmsePPjUsI0PC7MJKSu1zP9cFmsNSoo3GeE1BZDNP4C3/PjmVSF0y2DGCwdhF8cq+
1IT3bE069s6MFaY9u5PTesPva0igtFtE1R9Lrrpo598FGVEqHPQ0ziUVBeeDlea8qspBKn5iXQ4p
yxdIcplCUGPkweM027XuG+Tg+WREPFRP0nX93R6xko9Bxi4TXIkAVML+olozXbnt4UXRlhfoRBw9
OLjYf1nbrVa5e0K3HJeAgJuzj+5ISoMz8LP7Hr+FAgCwEhh+yBgSPIglNXHA8VrWQhOw7goxoXgY
nMmy4kpYkeOeF4Mla66tu+mgprY1YDMb2EG5EHAaRnF/S5hNAo6f9FAPd+PT5ug1NggC6VtUKJXd
YV4/T/5W2byPJLKzRgTffNIzzkYLVurLCgyl8c48C254RDaKGDfjxrDnCfi/tyuLQaQs/gkxsKM6
8A27rQoZIIDBS5AEyeAWckkU8ef1yvYPXZYRwQ6j1qQ/N426yEzDOiexst/hUNpuosU+rttodnGj
pEBrNVs+ZnydEKCvFkrovrP5TnZhyd3R3xqexclxG9woC+KuB6U5qJNb8R4W2atACTl3y0tsfrGR
v7C1NALr9sXhrGEvo8P16F+XENiOL0Ie81ISTvl2Bn7xzCT5aWS3piWjGDEMEjO8t7qRS4kIcEAk
7Hpo25CwrrkyO6eb2HXOb6sDLiAtwaCPquSkzM55EMvihQSCcM9C0DZO78bwv0TyjqYMl7qIcbXc
boMUtT59oKsyCORb1Pnk3XcFEwo/Zfi4i8VGLSSFK43KnXaX/h/QCfkUD8bptwTwNuMma0PmfPgV
Oehd2RIzqo7k6vWIRzhGyY3sv3rtkFioe+F+i/Bv0ntsG7DSb6Kgv8o30qBqEpg6TwjGMGTBYHpg
uKpUTZuM+kMc+arlsgqJsNxa3bkZKzg2cEeXNs4Bei4XYD9TW3rxoyWi5kEg+TSo75J3/4sucnkd
siCQ8CzKffw9ZD4TOVedgCgNZYzK8QqBw0h90mTtnx48O9YwRxDALUMzLTTSHB2lKVLT+imDUuDr
bWgzRST+S/raI6hQksbKkI9/9HLMvCSffj5/qZLuDWZ1uqf7DlbuXroXN5ntvfTtpYHA4pTlbSHf
qzKXf46PQoRi9yMaFfRVonzfDB7wdzNqYkjyZdH1GsRxLKbdgBk22vs+Wj/Ky82AclHVMjSvyrt+
90lY34j1ZVeZim5GJFsB9TiIzQsGoeND4Vzm1CBNWch5/wQmwgL9TCnW2/c3UYlwl95fUhNAWcJ+
GCGVDrwiS9KPztVqkcQlqIa+DICJRmYwzPv1x5eWqjOk5qHTyfywe54ov2Mlrpvy3SvI4o/Wd7S5
PUqn6PpUOqAb43+Mt/i7KsFep8pKNm8PRnTCt5O1DCcIh1xr01q9e7pv86rea0OfpiM/s0+jXvPw
F0cX+O8MkfiKsSCeTaYJ0Cy735Vnr7V7tZzqmROHCF5aI5FlTQH592gs3QKbC8QigQX6/OQJfzX+
LOF8Ax3GnsixW7X0YREvMwqpXzyyBxw709eS8wH9wdEUDP/IMJZrCRJNk0OWGRBfjjlP/1tVQqL3
HrTfMF/Zy0zH2L98r6EydrcKS9UK2aWKODHcAQ4xBNtef0RHHas0ClslQ3NirWFpdjF/w36xqBU4
oiaDWX/PrqFixSWqXjXi9e91cIkVaXcXNHgIJ9CVpz2XBCuEfHoocyFGFeKcimVPYw4lXbctImjF
hDiak4sVUG/2ENEWsKeGxU4Q9R+XGmxlv/aTrE5RvRlpRrBeld19wGFBJaQ9qKsK8EGvRhEgcoVK
cLKt46ueAeUYYzNLAfcSE78cRUZXIwfTFxLJos5h8Y4gRmcqWRjs/ZRF4Jr6rkYXQY4DiwvK1SRT
IDla8yl+V0M/CTaGsDPfkfNAa62OBOtUTSbelZSNAGvs5Ybfx5CJBPjUzgpWe468tdmcWqCBc+l/
dtzAlNwdQ9PnouZwjowgw2xkkRoHGIG8qs1nM7OYu6/jPVjn2LO/goFqwfdDP0qOJvWyLmMCp6wq
KT8YLgKPTjukhKH5/QHfIKhyORKhh3JyjyqcXzDAW/V5yt87jDOYRjKF2g8nC24pi7pJSU0VnxwN
POJ4333y8DOUalxsxfMvtogsxMRqpgFQCpZP8cPU4ABcg/Mf5OjwjiQ855PbAzpukyWA7g19WjFo
pg/DfCg6KERgSjXXOcugncEM7SI70P1+5n6g952Ak7QBnefTuQBSpav5dYFOypR64Unb67qTrWrZ
Wp3eSlJsBI4yghbAa6LI9BYilhZ/+JjNgxPjWWuYP/sveunXz9hODUCIBHjgfU9Tb8FtJHiWLkk6
usF3nszSIUSQ8piu5oap4JKqKMw9n7NoFBD58WYllCuku4DV8m7MKr8MYz8SGbi0y+vu3ue2vJU3
biHU9e22yGz1QYrDbkT+ZbVjXpDsj7rtTuVzG6buSMm3PtL6l20Tk6saLzMF+4zfUkX53igZ7CAm
hJt9caIoK1ymNd5Z9q/JP0htu1c45HyvkSAlDMqYJv2rMRvCCFCVpAd99gIJLtukK8q3BaSrNykT
/4GHt88e4tah1VevyBt7uTLS+jpV1Ig4jAOp0uN27dESM4NUqsGMuG9NBWj9ujQnxgoCee3N+viN
vWqpVzqI7GftagG/+VdbvgdH7OU5qdz8vSyuQtzOYJnx+JqHGBqK8jQOyx6juNUPsNYvjxQZbiHc
iSDfkdeStmgRO6wlIPCen6+G34KvP+wHtq2aQY0LUoex3psNNRgGIu9P1gsJb/Qq3ABWGc5K+Q8V
P421iGUsbo0Hw9mlRp3Et8h8ROtn2erOVo/Sgt0daabLGMGucKcXVkEZgZHoNmPwe0Mq29XsGkH1
qV8JAfvoSxS/oKXHFwyZfR/HX5tyAxwkjjTgMbZsvWxxE8RA705oSnQvFlyfVtEZZe+Auj5vfhHO
ZcM5Z2rpGuZAcepQ54lFd/5eFGkBNu96y/a7lyDTiZKA2IFSs5iO0gQ+Apgnqk24yHNUz2z/QFff
zvhg5R7tyrKmNBvEm5tm1TA9+D3lztcGAbtC0zD2gnR8+4dWdv2queT3xhYB17of2EOHU5bAupmF
YQCbctffC/r/0tZl+OZcHYjISFFHHLb7zgue02epDoYFH0GkWJ687BpQ62snMrQ1z2G7LoR61LRs
zbdUIjndsV61D46DPqSYhlSqgjruOmhfvhnzbCskfrmM/G2wX3TydsvK6CL4wry/bCiC/XN7VxTS
waIoUwVEycxI0e3TX/2ajyB+J8NYRYViHcU9YpYZfySh5Ch/sQ775UZdJuVQzJgfBNqwvOsJeXZI
lhd+O04msblN8oLMXdSn68UuW75AKSg8aeHsOYqTfcXvy7z0GEgZQSBU/8gU711Lt7adj4b3mYlZ
QYiOwXjzItbhlMBPNTc4HX6cCxuODOTaUgvL1Dr6ZOw5ZXCLmVvEuDrPZCSmRiUmOoc/1eU+xKI9
W5PPPYft6foL5nGv1iUODa7eObMfw/BEw7z+Sgl7llKNuFGEqL4e9W1pKbIlzusDApWkopTYiEeg
CJ5nMw3O5w9/YQbvVJV++uGXA3oHXuwwjBS7n39nsZiLossgxKlJ367ncRhoqhM9kw9LCno132Bw
9SMGMB6o2ctxsCE6UhKLGSTncm2l7R5t4HgmeNUfvVFZ8O0+8j0ra9aoh0vFiUCFCffiAe5nfhGo
CclaWJuordDBD0WNujzc47C/vNqD3Evbt6GvhbBR5EisOmjdfORAfBOFdl5a0stJoonHWeuNxelH
JgBGBYyK0uKAq9ell1B0JmD2esmJjUYND05xb9ERb+sVebFRn02HMGsoFu5TEXhC++iSV1xE23Xt
Jo85XgHGXa5cXVXvKCSF7aQ711RVkzpwk+00+h6w5m2r6mh10VYfrNcc8DP10N0I8uICi6Cfcn6i
9szcy8XPRpZpR4e4PB6TotA8/W768OBd6yG0R28xZriHd51CazVQ5LGKBfYkhsU0useSVcd1ydLB
Fu6mjudtLCe7YuavyGW0JBaffOS8CPNdSYvrENo+ahjw222G7lkWsXegG8GmpL50kWe0mkzDpxc+
FzvRgQHagognE9GPFof5aMvZyHDmcRRgaMrFGhI8I8MocwGhIGJ475CfZzw3g8KFvAVxJ6/Pp5ff
MvPTIeXVFYWPoeFbTwwNWcPv5b0pwk8DKRxNQvTQ8PCVpLYWEGYrspjJYgdoJ3HjFnAydl772xaX
dT3WSNrw0WAhQrduvKSvpPSg6LNDr0Zq2g4bgB+wglGffwgaZyKsRx6J4TdnQs7Hd6PcSkai4AqB
XXFCamzm7nbzbRv5WvvwM08qtXQLgoMC2yS2vloRLnOAr67xCv7vETNIJtXWCo6qMes1OSH6y1wO
tjS16RRGkNbNyFfgakH/fQX2PocQukj9+K7aDu7dMztl9oCDDC1DQYwPtzqkXEiyUoPvkg5uih4V
mDERogy/Rd6ePkK+1GKA9Lem53FcKDrInF6QTtv7CqJqGh5OVxCsfnGeRT2oOYzjo248ilr50Ojx
1XDhfGOW3MlmXB59LsWejf/3BHXc268fCQye9kZphjb1ljQoMOw/K7SYKavsf007rreQpB9voq2U
V6AjQwIrnaFs4zwO4e94Qrm3McMAaUz20t1a8wIntXmB0xM+sUcfFUDoiaoJhre26tHI4v+Sz83V
/kK/ZhYxdzrXG8pj9/RJS0D9SziTpKoGszz0d0wbNdgC+Im3vTHMq1EdWbmMmELezQjU1d3L39lS
gvW5tUa64+gZUzU5NvOfi2wGa/QGk8XwcLh727Cxcv1cnLBFlXmRbZxIZINs7bL4Wso77XDIOP4i
MSTZtrNu9OUCRsM33Ui5/J9sx6H9WrxGDAsU6QeJg6IiO66NwXawWPTrYmofO8r3VLT7C4mQ8uRw
V7Q9aTlnKgEJm36Y9uNFKR+fvtNoT5Sz8LLK663iKC+KIqKNnsUf7vELED2UoNAchCjIt43Ea196
T3WssaEXKmnjuIwoZDmTOzBuH3W/4B4iQ+7Pf+8soK97lndYwW8QJy91cWLfSk8SvqK0YOt97MlI
cDiJw/3i7UFMsV+Erx2G5H80Emv/4d/9URAhi0PCrELllJYmyFOhhmwd0lQPMZGLuzDfg7bitTx3
RfrIYlXqsLF6+EutSvrefROkeqn26jDLUNytD5TXFi/RSw/zj76z6ywoE/D1vb3PSah0T1jfDTmz
pH3S4VnA6ESdHCp3nOgAijZiLCTgfyDWZr5ISUXNO0EVHePNnPFCyR77ICG71AJAeyoAaUIqxWyS
WzOncQQKASGPZGgDBDM5uxknUlzErV6hCr65EiPzCTqMVEkKyBeTglWij4U+x9UcpIWsuhihUvsA
Ls+pfzqXanaXqYbWt54uXfyuEeWB3aRN5EOsZn4AZdL/zWACQfMXOsu6IKfrVn0OBFffham7jt/F
ECMt8Becmgx4/hpCfIorUOJPC2CZtZaFtYSIPg/5zxuyVJJuCWnz+dgizlxgsPr8ay6+pZWw6/UJ
5RWnORMF9e1R2J2PQOLASD0y7B0Pk5ISMiI6vGh5R+bwfq97rdR0pVERWU0zN52d3RjmPp3eo92p
TjKEWxMq6sfSSwDNJ8Qq/GNAOwzCKSbGQ+DjnGS0HLl8E2IKNsaYgLNro2FwzNPAYKxyJWOvZgTs
iPZcfTcK4N/RwcaAV/OWggCqQqezZNJi49Enn9H+ohLf+L0YoL300Hcr/mf6ZUswMhUdlrixzcjA
DkYUEoYTDXDcjJzp402i8pwotfpFUwY4lU1nQttgpJpFYDiR85BFF100HZnZqSzhoBvkZwQmoBXV
ANe1plpoptaiX+yU9xXFAglTA9emXE8N9FlLnH2b6M2Mc1qPirfrSd92WhW+0YWzJyTnfs1Syh4W
UDsbMix3koB71V4dERa3G/Akv8LgKZNr4tOlUZevunULrmj1VrT2Tlw/q5VWAUFlNyyKbCIPSHq5
eOji8Dnte9Ehz6Zus9slyoYqQvmujj0pmBPrEhlcmyfWsObTc9SwR3kYj30FzOVermWE8dETBAjr
ZSuBU4RdCE3Z5Zy3kt1ANmFM9uNDHNfDSuvD6TDbzVoFwDyU0FYoCKrV2cXPPV4zD1zC9PK9CQal
5cdYzCtdfzeLg543COIFY+MkVhkIHychHkBZH/XQrvQd8LTJ/5hTJEmtTlVhcEELwZuo9R5NIkrq
wsmSzkJgaPi/GeAN1Yu+v61J4sp6KxLjob/mwmf0DyC0jWFW/aJjnuJeD1mP32UwrOazlqqR+XFp
2o8FlTRLGcAIdf9ZcQ5upreaVNTvdhs4TU+of1Vmm0z4OTE/wAkQ166eOoptx2N26XJPU26YRJd/
vDT0ctaIED+KGbKncoOlXAy0BftmOu8z+Fo3K2MuN1DW1n4wLqWneQoskbBs+Uz/VazbU+NMIV1w
DNNIxxLNYNJGHjFTg+vFXNawCRR0sKAK2nN2m2BVArlsdbjHPfSybqvi+wh8unuNzgGzJhqPNKNL
Iab+W6C6v7PWNgo2LAd0NS3xluxwKZxe+09LHa5YIPjpEqOt5Fn3nuzXg5Yn5Vfa7ivMr46+CprA
0Y1XpQTnFlOtUqphmcwYXew0fIXRo9vMmXGOgN7VAN81Au5+wUgJmdIIQhs4wHEX6SBXh9KXIxFP
gsFqrA+onUwp3gWJlIv0+uIBsVJ/9iEBsos6vfDeLZW333jwqf8LnSH00HUlQr5BbIUCHqhJuu/k
4J4B7Cla2nt8/1Wa4RpbHHkoIO0NwxBGDcqc+WGeeQltp4oxv+w46x+veS1I3PJypoZPT8Fs6d/S
uvKOT/zCt41G7v1t7rPGAAj24WDxr6y0PSQZ5L5tvJvHlbWQEXNT3zsLRNXShV4Gi5hfCo3grYVp
J/Oab0s2NWyKS4FAZxo/Qy4rbCoIKh9LDszHaYZtX9IbRndguz4CH5fCR7LEcouvMD1vZ8AhqYbg
CfC9uDhM00YyhEEhd9T7AEyZIQTp8XgZJLfrzRUkVhuDKOHa+ruevYUvwlXKysFEeMtCa/1WwMKa
PtvI9k2FqHWCZpwulOg6Ddm5PywAsYPxMYwBsIyJY5C7bbeGUgHJ88ZNj6hXrcQvfc02Rab6tJNz
6mg8G7K4obEzUUvwL1MZT+UB9eZnIqNutaPK5TykaHYET/Zuyl8iZB/wUn1eQ3+f1jVUvLJfuGRK
mFagBS1S0GNOIZ0gQyuDH6xIEDAOf7vvcRQtLeLOHR66uDMPfYzhxD5tGRimCkl0D4wO0TqPwrt+
3u04o8DX6diM/Gtj4hlq/eHWvMzZCtBn2p7Ubz2iKZV/rszFyLJdp76m41vR2f8dxYyv0ElQJ90D
UA/OHj1vPjhN/cx9u0m1g3rO4F/I1+IjMZJVrrjAUjarI/GW31ZLs4kTz0vFO/YGWCQoE6C00VCR
Bg1CUv1w82qqZ/UcKPDeeW0ndim026NbPk5mpOaNhGFoNWsuwQDeKP2bIZBBLtVLM8zfP2s2TYAU
ewTi37gStzMQLKndkpclXZT+85ogaa9yF2snzGZfwP1UvAfUurjiUI/cf10LKKli+F09HfuV7sda
ry4lvIv8p6bhmOAWDQlcM/JV6cEeaeMYO1iuwxfUbm2z2Ns+QqvHoGXEmt4a2I7cts7TY7QPZpTK
lnKF+xmZhiOjOEUHl1LkeHA7sqnD7aOp9KiOfuVhgfd0AwEz2RAb68Yn5zNLIhL2WajG/kgctTXZ
Q4PRI/CiMm6/zS29XxHD5K4IDcduKo4WSQ92O8Ia0Q1EBJwooUt3DemaqsyPKwHMB2I3D/Dmz4o8
LFhhpJLtLHf51KF8V7yvQfBdcHzNKnyMvNciMVo0tHNqntaXiads2btoDlYKPYjTC02DOYL9sWdz
Rn10UzUrruDleSgJJRliIF/Hbf2PbBEid0e8JB2sCS5x6hCjsXvRIqymvfi/EqRA1Xw59jR/BcYS
RCS378HNk9Nwnt5NV09vyUFjK1tjkHYjGyh4DwbugPZ27z5Njf5WbejeC/Qi44v/9Zu8DfT86Xqx
Z++UY9xSN9xHDCPWHoqs3/X9Uwor0dMnCzIkO5hxcAiahThMxDVku8ygVsDIJeKJhxSh90XhVTFP
BtN16eQRXv3tFChXINSkpKsL/eQie8vsBAZqc8391vEXIqW9ZX+zsYM91sZmnl/flWmoAg8zZsSP
LF6oJZwwmS8xP111hzt4j2fukbllN7VLZFjuWdKNCWa5rJ3pDxx6V1J714dpzBeiuWICdH0b6B+T
Xr8oUdIR/ufe4K7vMHFhxUVfA+hZEMBHxbtjKc5hGI36R6SmNwRAr6cuj/qvp6AyOdG2HN09FtmQ
m9PNyzCj2U61UM8vBS0xEHT/CbfU1l1h2dwAD0OMvO17SipHtIqWhyHhRN1utMCcelzfAbPZEE5n
+GFC8hZY6lnuLaxYXhNYaPAlIGakTXzljjreTbgVUdgaMgAXnULLVn2LiRQoB8UN2ICN9VDrfNm6
iiJ63BtJYjJCKb7+phrVDm6yiwhClAUYd/UIDtEB1BiTyPDHeOD3KYewVi5v8kEGfrzmqjxFo6Ky
SB8JA+0LjWeA5SwTpVPsp3oJ8FgEsTF4f5Hl+IzspkMAP9V+NFeo1O5Vb/w16A17CkgmvL9GD3mK
wP4JZL5jMmwvk4n9+4wHKw1L+roAn1uw28QhMK6ng3I/Mi2CaR3y0yosJKm950WhTvQycXfRCZW0
ql2+etX1xl6srivSThrLD/AngY7HoPq5miV4Y+fzVboZFQIFUPLG1oVtEYCQXlw2DZLx2VwEUFrj
+m+D703BGzFpY68cni0Hblpe6yxQsjsysvKK5VobnHTxPkOdRhkYjbJKbMufZFKBM98wa+wd8pOU
54lh6aYvQl9FOAfNtb+ZLUaXXvYzqurBqLmzGRmPpmCrSyFWE32FjdIagjgPPTR6Hag8aeWxvtzs
lu0liq+m2Ka2tK0VmYWfz0sKawj51t46OuJd+WzwOTxcQw73406IuE37gUrEob2RWZh66h8JB8V9
8fw68cK67ssgZJWzPznV7F5Nq1G0sPva71hwM/xvvJWnmyYZM4XcC9+BV2uW9LxO0jK+2vgC947I
g4P5miqgIF0VcPWFabHPSYETeunIi9Reh5FQC+p9vzta4+YXgz6s/KrlmbTa/c3fS3mGb7SpUjT3
l+r7z5pyUSOjp2BTrKg66y8QxqYiJAtfFLmap5i870h8uruP0qus2mZ2i1jsHu/J2+uXt/gaoSPG
8FN6W/B6hvzOCSIO3JrzkwmQpd2G0EdZn1dZGr12R879jBNZoos93yzID/CTocE0PUOuObZAzo58
0Wv/0RMsEAYBUT3QveM3R4gayC4cYxpMRdnEGHcdcq4tIHKS5hAbwcvT2s11Xi+tNpgia1xFjy0q
sBwNoGbsZYCjaUDBCZXb2FKpM88N7vYtri0zuR5V5bUxE1KihCOYhlyNKFTD0LLaJSIYdYRoekgb
A0oHOiyPo8jqXpP1kzkZ5Tn5wjulwJCM7/WZ0sCC6q5DjSuAeLXsPpjojit+Ux3RzyxdiINxO3ID
WTlnBanx3L+m7oyDfEq0tFN5maThMhdPrrbY0wEwmjyMWOSEm77QUzfiCVUblAonmR8B5FJEXFhK
3qrgTr8klSaVNyR8ciROevdFRM+yBRpx38T1u+/HCyY/1PbIOlYcmmQKlJZzzAi9oE2glglouohO
Ms0Pzx4HK7sMjOSAHMdYDAdK57i5xQsmVWlApoKe+IHQQPtNhtsKmjqEU43pNUF8oxIKsA98nOJF
XJmvK3afOKr+YiTtaugg4EwBAY/kCXlZLb05f1xT0Cd5nCqBDr2F9qDSONbWN8zw+s0+FiEJU7ts
ILGyYN2b/tmh8jVHTyQdj1HoXek3CAzG7skV0EeiD+gpmnShwMsovEzio/k85aCEGZkEmSJx36Sn
wlUBSOysfUJEzr1paJ6eovKGyPzNfN25PTqWPJVplI86PeAt1PKO5qDXpc5o1SEsZuR5oclkEa/0
4J02u9qI3bRWFCo+5To/YN69Q+vZrBdfUa7BjNstsZYvcj44lg/rEKRvfAaLaTKzrcPFG5xshXYI
qpX4bZqcux+jJi9Pno/VuEiHluggQ+3CSiI+LAZ+mUxXRhCaWgJgEBL/D4cKRigY0woW/68Qu509
zj1pH3TkX9AlKcvKKpvHz9EiwcB2beM92RW8YWbDVkta+sqSjb+rqgC0c9CN1oghC4RqvcgbVfxu
W0K71oH2Q3jpvkKXC6NpXHmc1pEUq3UyZrokbzrv8rEyTNyVYa/EA+ncpzwpgUNS4polguKsoJ76
loXriO10v0ptVEWTL4mRhbt/QtEUI6Y7m5zvm5W5IEkXFCpKrGWrK/FQaKuoXfKRCVxAgh3ZF05p
lIrR4r2MH6bAGaArc3sj41II2d+vPyd/uMDYZ236r3kkM1XUkmGSwApHqGISnnbSY0fOrsYWSmO1
CJN7Wp3bzFzS5A8rV4KkiaewOoGtApRoCfGo5bBplT3Dms2dODeav0e3fMchbZ4Sa4PZvWBLcm5K
1mycJWyNQMUNSHKMH4nXNx0G/pqYEyamaTRJ1Fgpz/N09teLetAfdR0jTg521f/s4itUJ8/xiP8r
+JCJ6WLXdT7Nd4eHPGzZP09I2/UeH/TYh24avBMlFLtEyqccMVXemODAdPxievQjh07FrMoer5oD
c+TyADJRQfCjvJC0T/wFao9E8YATU5RS4GmPD3yzFLCRkAeRQ0t/34EdWuppcspFdHrBvqIhUax/
UDQJkwqeWUbEF+NV4d1R4VNQWo2ye9c9F+2WAhLqBxe+5O5khjGHkZJ/1mMTvJosBMefne5gy+JG
CmI6GeR80Bdmzsp198gymfhDN5H5XEL/GL75r8OZLNght39hy5jqSqzqvA08VZ6crTl+rSwmVQ5c
UMImIhrGcwTixgO6CIAr6sg88qdMde2wBO94USo/Ipi4DUpV/8kLeWyUqXTzL/7A4q397IJVfty0
tF8AppC1al2Fna4AVgfEggh0wCmRzQXUF9sCxZG5CBntIqU8fswsX+pre+WosSlT1P0DYMylWJeJ
TdlCqU2k3PdR6aAOhfUdP1YRQb/Zf/jNvRVgb2vQNf/E67XbR/Cnvnnj/ksiAOGfNVQZdVO49yNE
E+q0g5icYBvz/V6/j4tmOqyYWPzl9ELa6It8Wscmzi546f7nY2hx1z+apqxDxMozaKMIfpHWohnZ
qzj96KFO/Eixbh8i18soq32QmFg+Rewp+3CxR2ApY6RyRE0jV4QBi45btE2epxv7y0rujsY/eP8m
oQHPGRRMh4Jb1NtC8ZWzq4HcFy0bNSbSgquNoNUKp41kY+G7chg+5Br5NFK9+88tKRz3wKovAX82
nywx+Cq2RYviJZ2mMTlUGop0E1Zqyb1bw2UXjfOKWaWax1u2skGT4O1LI17FrU0018Y+DEgVH3ua
tOkJezzBT2/gD5y8xvX0efPXMWSt1AHmAa2BbvhyVduLhtoANEFl/V5NZ13+Jb6vamOH+aCE2On1
vGvDPz9gm/dz4ZIP8EInQgLLfDe9Bq+LXJW1iwGK8t1PLiwcX0w8BWvIr7BbW6az1d1R1x1730EW
rbJ9hU8Egj/r+PIL4/2QPYWGKrmJC4eQK4x398OgfQR4NZxybC4IUNgwWBn8oiWE+z+D9gsv0rCX
gBroF6B3Ft8cc/e3yKVCvE7JAKhT6QmQJFnMhGuMOdgYDiBC6ef9x4tSEkycz7u+oGVtpEMdI6AB
uNrUFuUYcVU8+gEFiVMb4w/oTVyANsTnVGRfJq1a/SlgCimN0FJLPy5fa242V4kMcRJDMT0hR/su
U7qEw+y6ArkyW2/PT03Id9TxLEWV2v/UK5fd+Dr1T+56V+G/UZqZtvJMWNmvEUwOZFs6TOy8z4Wk
IyvXWnZ2QwVT+uYuBTqkaGuYEuHxj8gZaEeN4KxuTCoSwu1j9oRkwPG9bB6FUgq0QyqJXwlzwS2e
ahE5QHmoeKnLurAUrdW9pXxkDmnZIMiFAmyyI6cdK1yRZ241jxedh800a/pPk4fwaxdph4lhnbq/
0BabbgYQXbAfiAXoXIcjbw2pFVfJR497X+u8Bs3AZMw/H2TlebqWYdnHlEHY/ROeM7X9Cn3/IE8e
CMwwEOn14b8JLu9XnKcSk8vuIREsF6Xz48Nhe3eG4msyqAmezPRAe1cjEoLFfGejPPzb8ByEoAEL
TidI/gM5LanMQvosGh1uUc84lI4A4rcUHfPVLD74aysaFomhSP+EV5pjQOUrlekHEfJyZL9ehP11
IyyFXFtwjX4IbboY5PJ7v8BV+5/v6KtXpwzRY2m2MkHqOJpEpXPDy1344j0wdkp0rnNlznQz13mz
q/snFg+0L6wi5VSw3+6gbAMNu+3vDT2NCowagNLXNtX7863ICAdMueOftLoywlrBCPeS3JKLyZKB
1ZT7SNJJ8L7Yas0zeknYHDNLBYExj7buBNZTZdHxn2UJqQWws1U3Kmt950/UkHQVC0mz7PPwfb4l
Kib/jJ0mZ8NvPHmVSURnuX4L7t+SW1NSdgCOGt3IHkTQ9Xr7hmXGwoVq2bS39MceWzDaWPj2bERG
ShHxIka++B95y/zfS1WU0Nyv3We46ZhCfD0Z34vZ7OuKOD4KUqzEabOMZoJXH9eatx0gNUh4bAR9
Cw8j9//stKNsW/CfCDflXVZSiKBezqxqAtyDyPTpvbI6Seao1ogOrnxS2ZJ9wtf34k/y11aQnikN
/hXybUPc+8iJoQgaWfjYoQkkO0R0A1HkjXbz7CRbOcAwihZQru0U8FOgtS9a9XvijhqN2At1XfvS
zHKWsUK6pwcU+SJFiOtv+IlhKbwE1V8QMgKQpAnRbFXOvy4jehdPMbB6s2tjQ3ly7+AWi5ThdGH9
BC5G2XClDUMy8rdB21bRQQxCnORRfv4nTQSdf5IE0Dv94tameA++LuyncpLwLj7vfqUg3KSIsEXZ
sG0NKBa8IxUNuNGE5QpcUlGfTr2vZwgS90KJzspBnbRh+J1yRf804uKFuab8non28UEs3ttktGfH
RwXKkXKZdBMbw9cPJ/mCTDA08K5CIcwMwp4mP522gIb/7sRskgd931+bDcxB+yyoIgbNHQeU1IWT
Up+7KO3S7roNJAWlgJH/WcRv80gBKEdhJfVaP7TWsOUQVL9nNb5jn5Chjop0sF8pKWiPLAaDwfQ6
sN6dRnHDsmJEModHdVt5VADyL6xjexVrK13ex/Xd4iVRBbqUChL5hFgY+FbzD2CXcjilY/pxHOVE
xdWhiAj8VdxOl8GYVKNWzoKUR4V35lgXH+mdAEIlf/kR7G3wSG756dMAURjHOdKdh0KEJE2jMo31
6JTUATC/09U1u19z9d2T1pUEpDpWUj9hR8xQV1g4m/2D7uGNEV+ZzlYUHnMGzoch9ht5sVl+qamK
T5Ezumm2YKeMSmEcyljfxV/3d0F10lcjmjDNfx4cBahYozHIR0zm04d+SehsQT7pwWwuOW67PPU3
17zUr/hWeE5CXBmcaXWGkLiorl/dY7Px5Eb/ioSICPL3pe1x5HYHZoX3pWwHiSq78jqsGlMmLMVi
KU4qbstacI9eKGsAPxVKfMueGhX02+E94qHhHt4mxpLp/vMdJ8mLUZ0tRo8t1FWMaNY4Yi0ZpGPc
sdN6ODT6AceRt9iLQKz+KGtNIFAr3cE76m3a04dGmkP5fkXdr+kin7r05zelytJJUuDND0FU/0N5
Q/U0MuIvjy2kEpAO3efJX4AOHKW6X0YvJ9DGuY49/o8lN6PJaa722ipoC2zHBMfZMLbtgbH9IZcZ
7NjLreD0v1W4L8l8wLq0xc+Og1/rTgGVIanLjBcRV+bNcr9X4lRYB9o2he3w7RvMw6GmPtJE/Q0h
X294wplpRvL9wSSzgrlVZk/H6hWm2AyNOziUvYnufb7qz3Gy7u77+ZjQlkMpoTsIyKM5GOu2KDCO
Z3A0QKUm0Xi+qeLFuF5DMuYnab7wPna1Qw0mVuGL1bvItdbYYc1E60DX2BH5kQ7DmIZxQcZNGv8b
rA4ZbBxKppkuI5cnDvyDPI2e4kmTGHkBIIievvSo73UisGmJebeczDBAOUFn72TNrPYY82SNvA/m
jupXe4VXY019JBBZflrir5ImYOz57yL26GAg04GE8a1f7N7U9V/Em2j5L/9M2i9oOYbgWq8rAgjN
LsPVV40bRJf601v5yeXnJvlDysDFV1pF4doPU6PK57VkIS7+t7iIhfguU2ZerzMYyEDNaJqlloUj
w5x28CUGdCPs4ziOcd3toBPPs9Xvog90vW5aXfhNQmBWg+63V33GdHFP10pDG4gTy4SFqebLyO7W
s8jVQFBBlVo67GfW1KjZAZKOXGYOGQpT529muaCFL6bYr7ctE+k7TgwhSyMc3y+oLd76pYcezChx
+bwppbxQAN+Zj9xwNslYW/pEX+K2hvogsaR8/N8JZYp90wIADPW3/zbL3XADqyosqly4OUKoXewJ
QaHQ0Eqefhb+OJS7N5KaMZfpUHxqjEYjD/2k9LDfJm/Tac6c9i6i9smzku7xhKs/DrU4Aagsorpi
Dj7+B4LKM0teedhrslWpaQ0o8nKHZEZJ3YOslmqV6o61LacidxlaYY2I83hMc9SQXEri4sJWeDv6
SiKJBXUKfnU6/tfTdPdN24emmaDIaTAhSmVkwcDM9TkEaynY1R62o6KIJg0f+lfV48gbWzKMkhf/
LM+4keYY4TR2Pq7utOsJP+VO84Mup4SE5ZC74SapF6C2Ya3njs3Br7/7r25DSQLYhcpVIhZIDuu+
sp/fS5kOVD0DcAOWuePqjvzNHKSFPA+rl/1GM67bOKr5PZc0Fxd6kcqqHbJ7FjcN6h5RHOAgPNLJ
Io4AgUiMejUhcYH1jBUwYeM/pDObe1Whx3936aFhwQyvOPIEZV9VZBHNlpsjpETZX/YeLGTBm47G
YRrQbR9NrgUcD4VFwt02xv5lks1Q6qGVyDWGw7JPmihPhtq7+Hnom3T5ZNlbJjh6HkG2VphWR0Mn
eHiZjU17puwgUX7lbmmAXTZeGqoG72x4woWT3NOxdpc3ePf47ROGuZqmCigMfy7cskWJYAIcqh+t
SajmJ1VW9daDaiTu2tUFWSeVk2BW9ZsvIkYbnvmQLnJtXt961B4OlbNSG4VNbTdlEssswFj7Bb1Y
UoIjMzvDQaJMj1nAGNFiSFw7smdf3T8jP2/LAP0BGyDad1i0obd1XD+zCDbUC9DqWmFHtd8Otnus
4IbkGqK6uINIDOM5hCFlGybNaanZj8iX8FdpEm1CZ/TYq5eae7nBQ88/ObLYiAGixGeuPu+rpFTp
VHl8oOObk0mX7vUl9GnCTwfjJfxqiwKbKPviGWYo6FNk+vGUmmqKQuwm4aijkjZPwvHlPlxTAM3P
l1+MjoS3UKFDS0s9yQtOQpkyPEjP8lATEiqFNVljyqv5jtPqBJ+cr15Dle1b6/qdsVnH0dd0W6HL
7NTEJeGXk52d2T5PytHXgT3NTroEYv1g7Z4NJ3XG3Dn9ZeBd3K0/4yjKI6pDCC/3EmWMpLDbQlXe
p98NqBpbm6Jh34Sif/KTiFN+ypw4V2d09t0sUxihSQ+RRYkwryJU8PTnJO0LmHS6a5VLjERmFsDP
Bu6i+BCiMvoQ+7bNBSPNCZb80pecqko1SUiPmuLlSyvd8WxqK+jOceNcZarjLNkGyCPBfoyVvlwm
u2tUY6Yp4X9Bg6mMSyzZeoWyeY7GXdSH0B3hjF+4vuM5SuIaNrGykmIqiTxsNIT+WJVvwb1aXOXT
7yB2Lzym4iy/Ccppstns5qlj/gDUxbiRIs2a+0yrG7UgYGOJkGorZYmt5OiBGUbmZAOZTOIPqhyd
p3buXWAQ29yq0vc40ZgPIpbFd77fhVTK5EOmleYAibsF3CKhNDZEs16JWneCQLN4FyBPN2ywmMWv
7dKyVOx0xwgl0/EBY1PEHVNI3fajT/PsXBJ1oj7pCxMIwqdn1M04we+u72nz17GNjXTsOTgBxHRS
C6cnzizQjxygpA5VsdXuNP8yNIZEQY78KePXxOU9+EDedb5O8o/swaQnw5xq2TAj5EWJ8hEulD1x
EJHFz9E+EVHZrgZ5Ddu8pb/zZpY3ONL/rs1NFCbwa8q/oFpT+/z/wnJi1obZdScC8Lg6RpRKTryu
biU7ccUBUwjXMh1aTZsk4zN5eEm7P3AZyef35ac1h5+Bic3e+v9KXySpyfDGnLSut3BPHNNxBYIq
dDq6Gqar86bAyQJkvhsKYjc9hJoPyXTCtAk2cTkFCAqfI4XiNN2d/vG4c6P7fs6+EbSRdix38RB2
E9DEGZ2715O/CxfgV3nrqAIkLdJfhJsxpyKQ2X2Tnek6L+fhMNyxLqqIK4wq/zzMBFhaVWCV7CoX
+GrH5bxr3WjSc/j2cR64tTH2gs/FKkRu/R+GyuCFZraCDOydiGL5GN5HvU3Y+2/OHX20uSnpx2Q9
H2nOpoBHhtw+U3Q2r52bJAmaDH4KtUJWlrcZs0Y1hLqdINNtttZfyoKpfTyat354NuL1C7DJutzZ
ry4QBZMsqoVdp+YyuvV1PhbKO7DkdYZ0zx8hFqT4krKzbigZbV36hfE8ttJ1LdWwvGVzVdHgdaqJ
kTjWBjhC5WuhTfZ544uPCROWBlvK6FMZN15kdRuXL4wSlfBQ4vZd1+kHRTe/tl/BkGqB25IVoWIN
k8Ot/l2CG/L8U1lYrHiQ+Bs7HtPW7cb5V9gSi+qZcy+LmyUT6irKjIMhWj9570yRVP/+FWASbs7S
UZqaaOveUVwhcYMijDoxmFQW+CWPlylwiSfbv/GIQ0E+W0+oIgAVeSfD68l7iZvPxzod0dq7VmNq
ZZjp9J4YSQqlTbjWDh183vfFb3/XnwScHWWhlYzaqSJ4q4u8aBWRUxN/3pGdKoRsqdozb7xpWp2x
7rs90ogxYBMBMHrEiTgQLOla3r59CI7cOvTiJfC9khpf6luxVylBX+9fVtBu1DEQeUB1ASSVsYqu
v/7/RkZqf5wwpfateErvEsW8+0LC7CA36FOgvr2lY/xIxyLLiWvwpmbuNSaW/ajAAgUv7/C9HCdJ
zc6cxXCjHEVS8P5krOOiIP0dYOcTeorgBsO2DoT4eZqmIBsQzsjt/MztMFUhjslPGyH7W9iIj7bw
tEN6uG+Gft5Zg324o8uWGNGbqRih1rUUAs/xMWL1nvFEVpBXiHWJ/M0MjVyZ7v11JxNNpkSIAUCL
mSSb0nfE/y4Zzzy48JruCXbiZhi1oYxp8pqXLs1gQB9KSacPxs53HqjxeB8VBrL2a9Hqtb9drkQ1
Kq+kEjPhO8nMGUARylQwMc9C8mUnSotb0uQtX5DbAKNnt91nAsPQZWZC583UbS4dEy51u4GHthaw
q26zSVm6eHJaDno7FNHJz5LVFgDlq6pfvW/evE/vv5lJUTyTskeoRVchzt3ubnwPCuahN8UJ0LHC
ZrU4v0F4YJdLwVkUUHN/fB+ByiTZuQxaBV2284Kmr5CMUucFa6uw2Amx3UK23vDd/CSncLtXP5Nt
h7r7iRd6/cSH5Da5jhTYi+Gkn/0EsCwXhdt5SQfBr2T+rKpXFctSa+Lec8WmeUuVYduzogteURv4
NT4j5CbW4yglv+0C4ehsadlZ0hTApMjGMJPWiEZQyOv4T0UlA8Wv/nowjutvvqNt22KyxVZDtLWB
TMEYd0jVDP2rdOsafpCzpwMP0tpYuCwj4SoPCp1wITJctMFbeY518GX09DwxkF7KUfzkGJG4W0XF
v4l5IoRJm/9rrcHnzabM8iikAZxLYdIAErZvjYzOZ671b/gbqAz2nm4ZHUB6vT6nF4ITad6Otjo+
Sa7vP2BB4Dq0TSYGiaGVxzoM7DhXLrQ5IIY+p8nUSZOuSAiJFPwKza+BYEch4slqBynagK1nics0
ubdzY7cOg2yio3eW8O5SJgkFuT8TF7cimT14H/B17WEB74m5j+LQMb43Jmolzas+a1FF3Lfn/GgQ
pZFkUp0RMOfJzm48/SnITljwVMUaB7TXGI9etH+WYsKTSDmGRPejL7lr0uBDVtlO58I6ZaOdvoz4
54fM4vEHeuOlo9tpchQtQfRZ1jC24dadKLRLIPIJJ3Eyo4XFCTJE60Pe9c4aDSIypY4JxDukrKOr
U+g2g9MSKegX63y6FzkDjmM6Tawlh0H4VF14Ec6MdVIODVUmAHSzh7zJhQx6JvOryG25EkFr+jj7
D+jGPQUcazzB2tQVa33eR8q/WDRI09rTYb7PYB5Ze4gcCIUAS2tBjr3veSMcLp1BONz9zeUGS39Q
c16jD4UQSQycaENUkVFSzBA5XG57PXuV1M41PKQoaJqQ9iUcEC5eeqnN1S7T5HIhQa/NrJHZduoF
J+oYVetuQhbVB743luqwPfik7/q2Rway4KtRY4TYTNH+kILuAggH49b08spGYpBzE9Atgv7ynwiY
5flU3n+Hf/Xr6CHCX6fOSmB8a+eCDg+QhdtRZlNX+Id+2w4XFyhkcO3bNRMaR48xSZ467yOjBBkF
OQJUgZ8gr3sP46P5UCuWepdHWfFU1024oCYAQXYrkv2YE2UkeJwYdt88uqoPCx9gJWuk6AGusAfz
e73jegDwojuq7t4GHHNHvW0qfMRgKYtKBQaBRpAhO/m7PiDt4Wqn9G5GNHMhnpwy0lchJ3u4Iqf5
MTnLcY0r89Fo+4JYSlV0VI5N2As0ygygl24YzAmjKfREwKttHvVdExoVQ6K6MKQUQSzjURJ3lDTR
Xh6jQqL09UtZFsBC9mYQzu63MZOxGrqgfecQLeWjcY8hrHYSHzTiXx6TFYNwT6Z36xotRCDJsSXC
3Hbj0+seOxb6Itm8pISbxbhFG91eXdGqgsrOU594fJc+wYTUYgHWDIXXbg/nY62ey6sbnw9i6B8j
ZDwYT8htSna5seF5F8N6VsGJkAOIGkif7q7V7WygvzDz2cm/WIBD1kaz8ED/57cefjp2qII70rBA
IWiTPQC6G2pK3BsA07U87VSO6a1dYdtChkTs3HNGox4WQ1t7BRtwqf73uphbR+LWs0WxX6R/9KgI
gfAJiXXydtVNC109Q5MrI6TBZOLL1uomK6P9WcfrBa646OMI5oCLv481rJ6jKnDfLp+m69fabAnV
MC4o7ro7rOh1beXDK6kPJ9ObS/XDke7R/g0q0U/gWXjtqXqVZwXOAsSGvEL0VniEe3yQpmVC7mm5
Bw+/aaWcDNtgnK53NclssUayxx9CIEUpdGytVi/g/8InZmRkgqYTvDD0KqhoL5RPs5Gxw5TzFfxt
fyE8Dgk9+U1J0gbek9OvfTxwGqgqOhELPybEHL/8lGpjX0e5FOc6OzCDAga1DG5bmAenVCMDIyht
MEbNpOSFrLoRbmck9C+2dqLxgCnUuU9khJT8OwRCRJMhTOX0Vxr4gRC6KeESbM8R7BkV31CphjlR
zDR7EI7mV7jaUWhB521nkzx6l80Gx+iIHdIszonv+7NTpifTa8BkQi6D+Cxgzqj8C0oj9Jvy/EuB
Y8HJYvlC9m2eAQML80Cx4jCNcfLjTdalU/TfMbPIPYS+OsdGVY3Ep3Ws+S26FOEkIqj6l046wOnT
wTngnnCzEAzlsJrOlgKdhL2lvMix9Cw9BPkgNXGaxPHRGp7fE4yToqUX46NXauYlermz0f6gj/r8
YjwBgnzb2tis9bnDcaCTg/ZrI+yxtdM4Y0wCAi1iibuWL5Eah5TJ2GubrV0qJSlb5BGquzqYyYUl
NEPc8LQ1RDRpjdfq5B/oq5DrReMByU2CkRKdElxLJ/PJaM1E7ExuOa2VP3IIOSxf/hPJn2dAfN+w
19E3mrt2r/TM0Fn2LoU0uODo9hcRlfeWH7DQ8vqAKX/efytUNLwRwHmWY3Bry36YEsRZf8xIllS3
v/H6z1xnp7D1y1XYJLFvh+ioy7zJyDIpLPlQZhauje5kuj+cuVKwRoAOcnIFfsp9Gefnm9ejyqU8
CP84Gs3nglsKv3kEctEs8P5NZCV4H/JALpI0FO1BDiVyH43ird43i5pw1m2asIAmm/GVW/NTy8Pu
gpfrCfR/tGlJy042M2+3z2WSIws/QlD6ghu0TRp2xn7gHV0cb2i8yd+BtB0/W6ja5o84c4e78iQX
YAMKV4B7oXSh8Tq+KHvQYKG7s7jDIdb1V3nd4hIYjMqoHg7tWPzLBkpk9FnD1/0LDWbi6nXbzFKd
d64YcXL/VJXGGOrwT8WCiIiThYDr0mEByz6yu2JmwxkkVxw+WZDKIzAOyCTX9AeAnnNhyhbOBYSu
+gAb5F6oXK+w9ZEGx49gjyYPv/5wICIHgak0NFMT1HXgqhjXSv+LKaoSNXvvqzv08u1QostidyZI
dUeCxE7sDip+VFXQhRg41p6ETJAHXOnxNYtwFgOrv/Kaap87KHqf2xsRHFCR1RytJkyzg1JQG0gc
rEYW5sAMlL9B3YsIStclHgXg9O3w5FJSQWvO/0ANcPfRe1+JW3d2xTDTWwrbloFug6OANK4Sdp9W
n4GBGw7PinS16NudYvdB6i+o5NmbAVC437C60KxCjUwiahS9PN58RqIEv4Xhw0ABZrv6YIWx7UM+
xXLdEFw/O3P+t/Hl8b7WedmNzsRuDU9e/9LtULtHSTtw7tN8oXEvrZAzepMU0UoDl0i6GHNRoYA3
//T3d5WkXYFSJUmsJNTjaUFvxn2ZjVEW5fQarZB3bwp+jLYXkcUE1ExijMG18Ul8DFO73BgzJchn
sYiILNqH0QfpcCHjYKsqOK0ileR6RbhurxfSIdt+jBk9+Wzsh/6dhty2nec5EBjcKR61S34Mzx1Y
g1VJS597yKZgs1ey/QPoBqEv8oFvw4FOhTsk2It4wOh45y2artLi95/1XMCV3GVA4VOsSXoGw3VV
yS9eDV75dGMdyJ/NngtdJXXZ3VeU/WaLlz99nayhY4F66MtEaoka5VVpSV/ueQLe8Zq2GC5OExwU
ISrbt5meBz7deQ5fRJ++DWlRXQ5lcmFb+qswalYbjQ5+w9J7/XBUf+VVUmJjxfBK5Z5knE1IbPys
h+EczxvzpmsD+x8h8qm5XPRlBgEM8gF44rpxdH2XUbG5MO3ccgjNNi+c1DN5WBv9Vyz88Q5EGjmU
N12M3POO82wbzIonnipnmJVWRX+IWszIYwTRRUGTtQN6HR8cQ043GIlRhqcqJibDm1rWf0LfFc8b
e2NV0wuvVrTatiOpVRyG0pmAzMdWYvYWVfq5PrYhFZDcbAcQWhyEkpqiL9Mc7OCGSN0sIKETQTsI
0Mge47bsS0fJG92dMbphXW5jy7Q8WZNWXhLwKe7royoudFe0p3Jh9ikoDBdfXU+SJnEvGjprz8hZ
yOlELeibUdovmTpdWJc1aj3P6MOt6L2N5vfqZVitgoKU0wSX5AaSiOyU+Z6lh1Plb+WMYKKeehLc
G6RIa+8WhFqqteeu7Bln4i+O4njNJGsy10/l8HlN+gfDntU2vFka7aRQIdfdFXu5q6FOgzzCbit9
+WgPoz3Ry66ktkywZQU1PSFQ4XBYFfZDD1ZCWfvsHh+ZUvnNhgL8cuk5h1XqAzMIGF7WxeSpiCRs
sEiuzmAQ+paRuyGcHk8nZy1XrfJZX5mNmm1i+hCpJKiRr/iYtggh1ANIUXxrV8eFMCXb/RZlTUVI
4rOA0fbA677OTWMzwhZkicaBV4cGAwty0Fn51vGH3/ggGnTDp5Aumq4pU/pvxAHdp2+14660ywb7
cdOI4n6yRck7Ml7Q1ijw4yIYXBJj+559rX16HjtPn6LdcRq5jt+rXR/DpEX5sXTlZc++nOJgmUui
VQW3M2Y9dbkqqBS08KMAzkh7xxBHItHaOYmPmH3Hw+EI8UbklmXEg0fJsk32inFwNygwl928Qu0C
F0hrxEDr7l+c9IQRXEnANL1FJsrqE99woS+NS/8PBmCIztqKtxThjQxkUIaDVfegPcmNBx7X4kQh
+eSwizMWvuxwJAZcMBH+fMMhwDkUz8aIchQmF4CNGj1jwYI2v/SXMtj33riKnPLUnQDwgBLjtsXO
MnvBeD7hCmmAdKUOu9iBEy26ov9ZX8JvDEeunJUaI6tL5lvEVQTzTu3IuKmH4LBj1l3pWroJcscj
nI1QEdbnlCXrawReikl9P8qGVE990x39MwsQdb069VVTcaXa9U2VkV/3n840TdtZfS8TTJT4uwVL
zt9uWODbi2zIYy+3UjyY8VmzwM86jFLb5fxGWiU9q0ha6/BN8GsV35U4u+irMyhcjTeJyenUAe1S
FqPNYWhU9Ra8vThTwX5lYMYqdimSASneCfackHBeanplvmZ8jalFLx4o/hfpduR2m3Iwmr4WjJfF
a/GUxYKLeSqD76cD/3OldcM6Yh+tsG2MyY/VG8yntKOBFEjJj875UyI5Omh3kaeI6VVjPsEjfpwx
uTwno99Yiig9db/whzl/xU7ODBioDx9OrHNmuop3PY5PZkjRTjOa4r2+iXgxcZhcQSHeuyoidcwL
etXiO+/+Hy+r/ANAMQqVyeoubYOpJ1uEn//IDuXA5JY76yIuwwQBfwM3WM9KHFJNSMWVJOokcyLf
foZDePHL2v9ODf2+b/PMftMI6woocwQxexh6IQRc6PTS2KnwtNwa8UW7b4f9IDzN1mXtGFiiztzu
qwOraMdLkzQMdOznJgMI88l0DbDv5J68IxN4YZff+yCmMny8lm7HL/adrNzaeo6NW1yNl7upiBrT
OOVGyNP3hX08DpOFAtsGtTF6ybJLiMZuDxudhEoNf7bhim1/n+T86nqXIl3bEUqpEnIhfNTpe/B0
/mjfJWgY3G72rckZI4xWWtzP20AMFkypxIPGqNxaOWQMbYE0xbsuWWUjj/xvu/dDvAzW2KkXY61a
DufrALMq9fmFOGTjOpKxbW3dIx15k3s7abLLDmKPJZVmn4fKNLByKoMAO1gVkYk7/wPVdAd3lLeu
I/PMP2TY3CDr1XSfKBqn6WwcxmoKO0sZXB+TXt1xH7gDSZzcpcw+wR/SpFgvsmilMWcTy0uYCQ1t
U66cmYcuiSdQUur+B/2l8XnLXhU+LYb4IazHVc6SkTLhXqCUby8LZK83htU6nNzjLO/vFkaqJDqV
HObO8fsxb9onIYCV/zpkbJddEGgcyf2fxVbABaSVIwAOBUqOm3aBCJEnbuz2sY05+QdvXWTz8X2a
Xga5JBPkrlDyk3bCC7mDI+fD6caqp+J1brxsUBnnEFNdPYqToenLVZAyNFTz4oTkxobme2J/gm/3
KoANwtlhp33/kYLPN9utiKi83AEEzeZ/eJ5+XNXSOs4g1Tf03kLK4WG7SCvikKiyHw1jyi0DXe19
0t5njlIPR5ejfOIItgPkkP/XRhEC531ZmOWOD0OjiWHyb1MfIlhDghXQimontXjOe4FoVH9fPrPr
rfhHPIa92QqZEUr74bCicxFHDvN3nw70K1ZdYQbRhVgVSFrIy6BzDfsQrs/q4xw23454eRL0meAw
lifLkWjK2DapiK8xFkEwni30HqNK2TcpUuouyGoG465roYZJ43U4RHzwneraGcR6MGqgXDpib6ju
KLLqdOtuCQeRxqGBbm7sLtjyu5OT84vs9eYA78xp/Mnj+TUIbJ8PuVHN/SnJWodYCw9l2zRpOVoA
eVvCh1KCAiiL/6u32Ni12J7RgXzByOxq4Fti1hKficB7Tw9jBxqcsI1howvmIqQAgk994I1sKrXA
p64mP9Q+VIBJZTwEozAyJlANuULj0MyLgwGbyH30yfnLOvMdAgiwXrrb3ssM17Z9Gsvw2k6eYeIJ
6bhOzB9mVJPbiwHf+bh7YYyRqiTtsBro3QYtcqojvH+CpE+YzV0ujSzSsjNxFb+rSPwgPDIbGoCX
pVdb5FJFHPgZEuTVcWhm0xkBoBuwoP0PnhtOW4ibZIjAK/FOtugzEmRgpUp0fv13r5uu1IWZQA9+
Frsp6n7KrbPeIqOXgSXDaWvcnZhfzwJ6JfG4iXfyuy0cOrjJGHE0BeFLhTLM0OajVkCvnTQQSuzJ
/mhKV7Ip/nty+af/IZPD0IqIfVv+rzDyEEEVIbonAR1eArra1g7CNYx1/0gR7UyVVo/MeAkZaL/N
+aKLUnrjzZnLEZl2xWCpOodU9DY6E0K8MZz0c1w4y2rKsU4ho9dVwesTMV5SZ8FaiOQskYh/hznj
nHm+GyMd+pppDiL0OpICzOpzPLzZSGxPeHSGFjAHC0AV+2CiROE72BVp7B2mxoFpXGXsYLQ4TZu2
fomIYDQPx4IFQIFDsfgbXIc6Imy9w3QZUM31CZE9/pMyzuC3kLqP4oalGTuQ2be49O8S3d1Px0uf
Ax01SgOAyO+1YFsePy6SqxmZdZlTMERKV+JBRDx1QTePcj1J/X3CgW+SWu2bikd+ZL2UMZvRZ9Vo
wXWHshb3rWgGlc19LkACJRRIQv3t5m5RlZOVt+CqqA3975I1TEcaIpPeR1hF5t4xgSTMp4Ul1luj
lSyfgIH+4x+GEn82WyUGNxJtk/4Wd0UdFGHM2ODMO4AjQjZsM49gFeeKnzE8lDpOgXFzlm33/m88
cMdWCSrkaClmJ/TmGKmnO1rloAwB5tcDtmGNhXp8FF9hxZPyuk7ZVZpWfB6AEp2FAFRhBRn04Oib
8/X/oe9i1qyEAYcRY+3hW3Hczni5XrOEV3XIP0fagxv0/TWbaM8xk20afJuH5E7hqTjU2uXzIoZe
YO2JMKK5eBKvWGcMODXG124cBExUCC2tkvLGf8kDaYt8KARcJ0lYC+oTVhzA+UiYLjOfET4X9D/t
FnTpHZ/RtzLtKXXzY/mCwMa9wRRJ9zEScc0ho0oVokpEEtX3hWXrSLzlsEl8boeJ8Jwjx872K91G
bsxDztLS1IsUVx+kASPIsufG8Xxk1CRSMcN3P6C/4Z1NUeB71tM1HS6AN4gUpQ3H2o4lGlf9q5KH
v72K6rGkjrVOVEuFNGmpS4UDkr58W+GzvGj4qpr+K2PS9s6mN20R80C6GfQcaZ+2T8R01TIkVPdh
H7uXlLMYB+amM6FZa8BxDMk00JyfrVxzZDJcrBcV4QXwTJiCCJ5TjfcNx6/YMcPqWi3/aNFLkAHV
0Sagv6AcASJS0mLQO7//oj5AFIeq9oOVBgYJf4rQMHzg0AWE4aPos9RY0/NCD7Js7H3Z4Q5Ecfh7
ySdJeV9Wjrh30iZf2mtbmT73NTk2imZOg6/ijNpKGLidQddRN9drB72TprJLpoLqtLcr9sF9Sukw
BL2mXijyA6I5xQDikZF13VgBgfrlHeBb07xlrk4xCkoTk8ZknUGrrVMxT3bZc/zsQ8Fl8Q/kNVhb
df8a+JOADb3sgwKQFxdEbYoeZwJYQBba0biQAnvl6ETrckM8avLHa6JDxAiYQM5rs+iZ8QCevhjd
fYOoMbqmHzpTKcIC7nlf6DV1nOItlu3AAar99Z+CVFqURxM9ejx6skTjLLZ/SAe5XX8iniaQlCfj
McDpuQ9njv5dPV8EFJ6gSO8rqotBnxpKFG6iaozoMwMHZGUIeJ7d84c05wWW4L9zko0A69l8R5ia
fRrYio+bTViOSeiHz5wDKbTQKOh410gH+JlbdgwAbJYkddh8Keu7VdG2KPgMirpYqxzuVfgy5lqo
eez6llt3eMCvlgSVVL9E70UYD9OVOqjQlqJrKehkmf7lTptEC74/i84DiywrLV/FgNYEZIJa+fBF
wAouFZqdy3839l/YWRdUIpOCIBtq6yk+3QNyp5/fVoxrMctKnx51I5hVTaDA0xeYG4moWYxcKKWb
LKY234NUNMCWnUx02tvsxBTI8BITaw4L7/r84QJuk/HTSJzocgHeaG6sC6GngHxbqAEXUFNwfFTt
8WFWUkPreqXhP2vGOsNUu79lSgKMUZwvP+9DlVkLCOl0z7WGWY9FGWtuzGG+HQ22+FcQcDzLUWJ8
XpUxC5m2pq4px/eZGR/ZQsXLP4Ff8ngRqkICIfEQrip8hfIzXLlKWPvpLo/33I/gFPzeK1pYLw5F
mFiXK/pA+G4cNcgTqX52JaQB8kEQp3a0cR46MTbr5chv9MCEeAcZAgDOcGon+t+EE79gSDOhE9lU
9+lJUNb7Ed/MLllGDliGNWPQpvz30ZhYlFd4Qa/j0cj0SM6ptcMHFLMcMTfsWgGLHpdk5mWKcTVK
e9TalqFPN5m6cPX+76iJKC4NHFH6JRqODlNypvex5JFeADN2mfMzmJWdxGfyxd8q3NzB7LeGJAre
jWxqLpN2V6HXYXhdhdl0LeOrx7FkFMT/tDZAH77yx9fsk35x7q1nN34yt50Pz0aakLcUQ0/t+swp
xJRbGaztKI3X5FO23C2CyWljc3tDJzKwVGAHPlLajCNsRb1VDKtFgipP9wYo6APxOR+pp5fD5Vi0
KIvrasU0OeY5MqxhfwTqTgc0oPyumKIFG2FA4ZhaZLSZt1xpF465FXKannJlbJWRMuXj7BV5iuZS
k92MUrS0XjCXUjYEmRsYZVrTesL0S1XcLmeSvbAWQ185xeJc+P3SlxxlIhvV5cmwgJCk8fhX35CG
Zz19yvVJ0t3rUV4xF5YZ1me7mfcG7WTR7jUuFxJFcEPKKVrdPcft+D+28XiKPsmf/NxJ1WRnwwjZ
dzBXFSgRqpHnwtBhQE6T8ZndsqjsIncAWc1Bxuy8O7HQDEefsYkB4JsY+Aw4EBDVTzBYN6oGK9yC
8sYusp8d2W09e1V99bAOT7adlIY2SsiTWxafXl97kpR4YfAKwxjNNBsAQj7Cgb2CM+923l/EEANR
9eleNfCZERWbRKOlrDap8Uk1AAd2F+A5unZ7fKgnvX/5edawN5WD2EhecT+BeYXZPkKdQSWXNNuI
RTOLaUatE4siFp0JwjnICLikH2/+rkgQ3RoMCEVMRG3qTxq8TMyOclI5g7d0b4pVWazluvHGTVuk
tZ+tcejMtbAdD8xIcXo0WTQho4V+HmCvjyOrs3gkWHT5ANmCFMMZ0Oa9ie6mvi0TOvHHoDFgVuvU
0cy0p4yihBwT86AUdWHZEh8RIh7m3MHCouZfIWIoV5kMtHh5f+fj/foxGBDqjIWhVWXQY8TSvY6L
OVDaP6eM7S06MzZXJVbyGr5eZS4YhobIi/daH/hqrlDmrH440MhUmCdSUNlfkfbF2hMQYndqqOc/
6XO9bvccSIit1/69rhU6MYwsRwxpOvl/FuKwi0mthb3kVHkSvAdzFwsm6sqg2swvi80v3QJWesVN
4skmpahZZeKQcYu3zJdyFGb8fjOPDAe7dfW77bQ/MONGVMGutukXPukASiYcxyg2P1+v0+bHrvSf
rz4MwIz44CNp5BhvOanr9YGhiq+3ZjYPp5Fw5vFxT38cAqDNoDoAdSMfTtgfA98Q/yzQy/HamV+h
a5+kUEObHCiK8y6FUHY6zbsPWv2fKgWgIUsFZHXoxnGPDba9JJd5tgJ7qrvxYird8/NC8KP6jNc/
/t0I5BycjNR0RK2zFkjDs0or7UmRYIKPzExtZRy4P6lIJyduKShUtJxuqRuFXrG8iHAgpxpIVcq9
78HzZmMqWTSKxO9orEcNPVBzTA+HFiAgwZPwqsFHJnjawAGc7DjuEorijLe8YzoT+PhB9jjkVdjb
jAxNNxSYQvb2nHT1C0dqrxUkwHLA5RXul7DTS1+tSavwC1yYeG41fujFiCqqynwV/dYFxCy/8GZR
XQN82e8pssVNBbcdRPPgndip5AWS6RYuc2a+3U8TK/+iwz6D3HPw4aKt147+xlm5ebpjE+mf35PN
oUg2xB8cN+fmiOOVUVFiS7wOpvnHOy5InHJc5+f5KtxDw3gPJ3AbwaI4s/LV0mJs5jrhCyaFYPnf
Q2IYqh0YI7Ere/tXlRDstJE3RnvBKAwId5mELHCN1WMPOZdktYEuzapCfNGinq/wfrXnnQmAiR0J
LL3CfWQ+3qbZK7vwGpub5dnCKjGCSG8AflX+QaKAq18AqMvMEUzoxawZEcSBGl+cMTSKLsIui+CE
dnuEoAKPwluNjlAfCxZ6k8vhdsyQ6qQOuLGmoqx0YNOX9GdFhyr+MIXYxLFR/4oU2g5F+noJcxKC
9rPKmRJ5YrQpDjhVFQrsx2zBIJkQvu+wt/AHIxbfKZ78fnvccFOxcN54Ub/iUdb3vakeTJc1oXVt
BwjJusqVIPUb8e9dUVQJIWTqoezcFZkk6cqq7EKmjcSpxBx0w9xWgHdwJLLUWAJqVqQHMi+BAs8E
xI6SCd0qGhNM+LRw84t5McZSjgGYoGJFFDsiymuFzkhNgAwDGr0+WkrwS2XpRdIJ/XaR2VLQnD4o
aR5XIsprmG7nFXEh5pX3OVveXEktmkfjy/iB0jGElgvHCiarD/mlHu6sKur5tGM5wmwVkSUh0CsX
Q6S1Cng9ktAK5Q9X1muo
`pragma protect end_protected

// 
