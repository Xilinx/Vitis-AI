/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5920)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9RAxj/UjM6l7dkAv5h35yjN0zrqOvJLjtj1Glv982n3uIQIuwIKWxVnh
3hh2UtthEJRYikcnuiV0K2t+bD/6pOC7xRpWOeowX07hyyJAbepIlRUkbHxarP0aZKrYP18i6Ens
UjH40z+I8TsNFKenjsDPD+zc8qaEH+dbugratd0fSD7M3a88GB3L1JU7IBtMS5Rb7p41cXAI+kLn
MWHeyffWIvLR7Hx8ldCLpI1fdMGUGuYF4+W/rRZdpY8YWXHBIvrQJ+vPP8PgV8MHb+S5Z37NKBjb
CLbs+0HHaUz0hbs9HmrdNOppLa+K01sP5+4M78qZsv/tqjbaXj3QwROodxIqWFFEIxBT+IwSDax6
iYUmPOmGbc16DICeqWxHAXjfn1di0kHIVWvhYqbCSjCqSGW1R1Gcs3dGouy1Yw2vT3fLQXbOn8Fw
om9L1nGz8gHZ6pHMAq5SZQKHU8wD6DKZawNFmhNsFI1KjR3L/3/GZe1BNVm/J8akeTcfMT1OBAVh
1OvkyutGeGpuKg4UX50FEPLx2wqGxQVqbuY146dqfKyOV2tYcr/gvYDvoV5pDaVtWNddqa5FWZlB
IUtHvvDn1dSf9mVJ1hQ823Ym05NS5JyPqQXpWWxEiha6y67LTLn17kGd9jph6hQBZdumbm6zxgKn
51vhZ1spnDe1gZy9zd/U/uz/zQm5l6HnWTiR7KZRNJJPKwdeYvhCOOd0Icth46+rswY8wWqpHb9J
b6PFGQVUfeHOf5JI5o+LEbA8UDsMWPbkdHF7ZlvRlrO/UvqqvGVBi5rx/hHxjs8vFKdJrJeGaa5L
gcSdzGB1yTnZdJqJs6G2e10pD8u0vC6OGD6ycekQqWu4v41WdJ5BzqohtZpORcoq7h19iOGuIXZx
fpCDDM1iJa4UemCeSvwPGH+XpOrfFwA4e4JQjs1EucDBncTI3SvPy/dhz/6XkpTT74GkNfbBBpys
SI5NSrEq/o58N814wXVdS3rJ4nRXVNGb5n0LEFmLZmTdaSo+K9vpBoohQbvGoipc0tmooA76bJxb
JUisUMkp7uh/VtJbpjg5b4qLjEfxH6uBny6Q5m31cehljodquX2F9Zfo8S5ObywrFhea3f8JIDJc
UTnSL+ohzd2Gw/96d6u9w7EJZOdhaJDfuEOlJk5bXXkkO5gxb+03Th9bHW3WqrKlhrzHWhSy7fHb
sR/qYrFO+7XJOpInB7ZwmYawBCWTCl0CxYKZ7gtJHO+/vYIbOYMQT/yLguH8cVJdaDSraQZF0DGe
vTjNPLlCRW7BUkbLq9exM4MiieTxftq1+mRXBPvZ8otarcxtUxMmJ9pfYyB2tMQ79SvOYjc/WSyI
t3mnzrjfXVIfqt3LY2xJQL/Bfbo1yj+2gZgMQ6SYQvd8solNy0TZTYaKa9Glvs5yuQkgJ36TMC2l
Ix9oA4obxBrJeU//HbAqGKJeVvF8+SNygXl6Z3w3Ui6XeDn9+qSFMGMVHehJApJZQxFSCoJzlww6
8K7oeyfvd1VOlhShQaO9o28GhYU1hM+BOyuRobj3xrXRd8Otzk1vP510Og+MJSScoJKIWaiC8nBZ
fejSXK5TZDMklyTcz3dUehtP5LEHQ8zek8nwV8aIMKYquy2hxvie8G/oDhCXIrHnhGlIYC+HEcUk
4cNcpZR0HkUbz6QzlaYPH8xYhCBMxs34L5b0nm8lCObIewX6VoFlVnoEP+6BuEJ11vnGucH2Dp3x
GVX5YaWRKTecx/denC7tnEHjyB1JvLfL6Euls/sS8wFrNDuEXz/PKifjid8Z5Fo0MpJo5rmHxpz9
6Asci7/8ReZXwFEgm+SFI5g7lHgQsYuzGA6oO26zkHGxEVor1I09+PG/eQ8LWnIN2IPacDbtplpD
ebKYDMPV/1xJ4Y3ASWx/z3vsHlBv/Izep7yrflzGvKMB3lwTdnERNWJ4wu0oMGxjMldq0lENeOEN
PLIjdlvw4F+CKjXjE8aqdjYhdY3APlwrFwNODaTKHyKxBNC3u9ut6/PqFdVbjbChVNYxyHB31Gbn
BPVU78z5Y3yEC+8icbR2fIUA2HnSUtPgRs/I9l8vUZ+W8dEuo5cMXZAnExCDYIgNBq8xNmo1msuZ
rZHZvOG0pJz5gPsXVHP18RHEtXcfuw38WJYsAfAgG50KwHL7G9MSwn6WCqwCXGlRQdfwB7KSxbDZ
92MWc/JVx03droKBNkAy52ZkCfEH6jJLgbASfW9ScAkaNYoCy2jfH0yI9Co6e/4lxiirYKZa28+V
VEE8YBjUA5SPvRcvIhiAuyYaxgg/eHhmtntisrsE/DvNhTo/0Pqm89judmS57JEe3AZAE/VJr5B+
QOvAuIX6oTCst6F0TGprReAbJ03VkISZpshposNsrb/3WWxF4JZOX3rS9uFAdEAUKQdcWRSXkBNY
ivpnfERDZKf+XjWckHk7AkGDuTwFsUrNn7uQQYgnZkS2r8zvul7oZcisaeBn8CmTT4ZYVukCUdpr
/qy0u8GkM+z4QqPAkfXTk+7PwlynwFJUcKyBuiXIBXk/4RTIlUP3e3Wgfy5XDTOOuL+HymVy8UQV
6ifBYMxSySye+G+Y1t9BUs499+4rjF27obF5nuN1eJdZp5MFxzhYV2uzC7jluwa/oEp5BLYa2rbs
mhupESsqmuFRPvPYnfdI4Ln7UW4GYSbDQq1mKlajMh6VAGBcvrkjXYo22HyKV7RTRbEV+sL9M6cB
03YHulK5l1/G3zO6plZ/hE4yoBfY4O5OIjqrVhMTZPZuZGfuJou5GUk86YRmTb6ISaW+cAoySZEs
+dKQE93/3HSIvhPZvV5uEWAK04+xoMpGJpNz2y1Pp5NGDT2mwJXsqKmvmjq1Zkm+eqfSp2rwiMKM
F9FQ0z83LSBXgbbirDMOJ4gBAN15ToVDdJ8jW1kXnMK2CnsKfrWoAn1w+iR0RqzngYNGUgwU+LP7
L5+3M+NDn/bUzwWTAtRwPpkegn7X27UaD/CQGy4+Aw+vufT+LF3PDyOu0GDbsiXdqZEvkC4YiNzW
o0hgjYCj6yI8PAt4L9f+ON7eb2abIS2IvbAtQwe9F4BDd5iRaQBeqTvWeX9MAon/J5BTmh9e4lfo
YXeB8NLnkMeGEM31a8KWSk4I4IYaUiYlC7mHC9XpDuaCk2jJPLBZ+XRVNENjpshIwxV6zFBl6LVG
5/EpMaeaA198ABJN3FjiQsyH4x2uHEXrWxuFTJqDk0FG2tcLCFRY1X53lZOcFcHZlbDx+HbOmdek
5ptxcQ0tTs9Jn9EQkA9JBCf8NDUH2kfsb70Xk/ZEe8XAZ0Rg7mYTJcsdzKqGxN5nWKDYA4dqiQBC
LagEupKfiBYmuGImvRXko1BWBaIXvVEZLtIv0mH3RMkbXvEkA6p5IKKkYzSism+sfGYZ3Ppi/cCp
w8BX2YyQy8ZCUUDf6wsu9QI9ROE6hTEfN3xOkMdUA9QBjyd5sVLEukdZaz5LGg9O9eQ6OhkiRHWD
44N8CJqG25EZpnYi60/yRGHjJ5DLw3HTrAmZUwJcElKq1vRVp/3EdXlQDvgHFgGG8yaLG2SPqkM5
xD6XXzu6Rsf7Jav8it0bIqAlC+lfZnb+ybBD6qUgUsotnsode3HYGjq1RU8a3UHo3eqt8Ja6feln
k3Mm2/rb7/jtjTVGQOrit3fRPNVegap/2mzFXTYg8/h5bJpmt71Xfy1VAahACaKDzi3UiFvdWXvV
56L5rMX/jI8RVqw48IaPScNbIOCPo2x+fUqZ/MXt0NzNjCVVc4tMW2H+Zh6Wtrrl1Q15D9dDNosi
vaI7EBhdIT3B5sVXxGey11RgFva2JNuwg2zEioAna/4Exaq7RY1FGfuqJpZJzwtCch1oxxg4PTJp
Ulal6eS+GUULu2jmiqt5H/MicGipYln1v3GQY9Kc/VagcwAZI146UhNdz4W73oO06szuenbtk1VM
+pg/x1GeJO34ghRJtZcNt9evEF/Id16CuF6tItyEANI0hU6QLiHWAWrbKl4qn+HWu6I4peJNQhVs
Wv5Z4ZXBc+8gtGPqbNZiynBkxhWl0gfLGEL32Ru1nPATtJn61+Sxw4AaHcKna9XkR8RA+6Zak3h6
JpSUxwbwjLHSFAe7SltMrHoworn67ulHZLG6zxRoKCWCcep99Iat82pw054iPcHMW580MTRz17Oj
kka2qHxHHQK4YGRmTuQUasy5Is+2VwollhdGZk17PGMHMsj1SlDiRy+3sI9WqkqzGmr612pRL07M
2ogMRqKk4G/gSpCYtJATfWzTUCE2ULaVAz1oRKPXaD0XHJsdV2NAccjb3Dt/r7uIduucwW/HEmH5
cr52tQOBbyS11j0Pss5loZUFenP5tiGSnEAB0egEuJ5HZHek49O5Wj2JyPrhq3mYw0a2T8/yLFto
umB+lNUUioZXbdgTVs8U7runPYayrTiSEktiCkQqqwmhiQCOUabVQ6zozfVICVvlg8MLsurA+Wrl
QCZfBwyEs4fFNblY2tq4vMsxg0GiwKDRPoNgUCA1euM3t1F+IvenAAuEo91XKOHxRAGPnL2m0RXr
HZATZwl1XxyOgfKV7Brux0VLputuGeR9lQxEEGg8a0eiaYyeCDIbI9mfvgSZ++gc9fO0NcVnyisW
Zxb/UGIwBf16gIkgtbqpeaTl1Hanpeb0zQOQr8MWVjaP1sS6EsHOhqDr3JfUPtc307PS8MEBEV1E
K2udPuF6eI+dXbIMl4aYAWizTM2k5D8/JfowJoGYwwPoQjMgIUDGb1+GZ3RWN3lvTeGM9oNLVT8v
q7GHsTv4jZpNtGyLiBlzaisM3xUqQevXAvOcnGfZmhPGCmwieYT/Ws9lS/O8hauvCRCfSlHw/O3Z
7lYYf+7P3cWaWcQAKAnmXG4TynuW3a4SItRwVLxdQE8OsKVW/7TXIIScwvFg/XoyD3pjpp60GW87
KvVcmnohmstS5F+D9vpqg/yoeRf+NTirlyDhxzNVLF5hrpJI1KbZTU5m1aD5pPnQ51o6tW+qj9ex
5Y1t2v70ECKwb4viISiEzSQUoRDj1JJPkL36ZwiwYCqcvxmwJijIvGv43kL+hAYZXceHT7FsJeBT
aaTYctgcRtml3nPpxGQGyhv/74cfxPKRhTnN3et44LsSoGdi6G+D2/kQJxL85w4RfMZdXaKjCCEb
eLAc94Fa9UJBhNtY2P3l4mV9/f9xaOLfLDqOAKC48BK1u8u2WqpDjBMZPxXH14w7iaxJRTe7Ec8q
2bdgI20dWLEEhsL7LWW+W5UaQpgAPU25y3Ad8tfo9WGDlPHhZSfoiaseoLNnRrKnKPW7L6mrpSAj
aQ+1f1b2/s1zjE4AGTNm2dTLw4nCQ0/28jWillOdlwVPlNTrYq2bjrmVQtHBFBW8q19pW1r208WI
AUDzSrk5GVU7Oujft8mTvDPDA/plbWKVWFrQw4synwrkIyydW/OINc7rwVVctoyGFKnzk+JNJVaf
CZhehjp/kD8yRXsWiDVRJpdnq+0dZAQ9PwJBd1OMjF98wWaoh+lyEQ8e36VBAOMWv+XrJjf4CKTa
TNSchFbOxRmqKWW/n2WqgvRxiBKAWDNG0gyJRcWV2ihskxBy2ZHuYWn1bYcA/J4fl39pWcayTPru
8KoHUn8V5HfcDs7rVuTzYR/E3k4yV+sG7gLxwSygvX9LCjuZGkC79d/2LbGXfxrMmdHzzQU7ZSxW
KDg+XjyydzSdFU9k5w0mADSVA+Px/MUWcaltGcfYr6cw26hT8KiB7eM8bKQUU0NGnXfQxrLX9hsI
jv21kejSy8oyHav4DIdOazkSOoM18twPiuk+zPhusO2N8T4PB5VNrMyptGI0Z/O8Vd1+QbO9KXZh
JoLeOq66JsZcz2etiyik8yZg8msCOaA7kEOuMooQvLh0nfuSAN/7BcbLfJ8NWwcGbBoXiLjislkW
TF22Qw9+BH5iEiRt7VU2gukbHoGBD9Lg3Pn5glEGYA6i7Pxwy0NwEI4DJc+aUcPpOEWvTFzXza5+
uZhjLOETYtZQxnChyqmDFPAUW09sX+aX11SVywC99FAGFfICR9svlKUsXbsw3lk9kfFFlQicyGNV
nkgtipC2laf1dMGh/5AhYmG7iJ3iDXE5mKQZb+sJq0GQ2VA45N1PU5mDV9JdFft8DA6oFUaslhlm
yKOTaHQkUpb+wCusgOSe5iAEH7QBP0D/pHZZz6E71fzhzWtTlOkQ9+M6hZgt6t29rt/7d3p+6e+z
a8LUi9yArS+KTozMlnw6n7vEcxnpSnRApChtEIum4VPGqc3V0l9/Cu0Lw8LWh8SaIG4DAewkEaAy
XA8uy8y8mAiaWSNkGoZvpikukAkENFl6gOPUSZJU1zwJAMECINIwZQX8jiZhTd0q92ztFcuFkbwn
AVqWYKsp9MBaXuX5Gn0d6trLLdLkhUztBLyiOC2YNmaMn8EwImZ1BB9iCTXC71B+Zz+a+/q8pmpT
S5/hDnRXdPtjMKblEZXP8XV+eGHPgJILaRwiPAPbOtfRWkUUDUz1Kl5AmgNh6hTKQhU/qPDEwfA3
pthUQ5v3cEYtGwlU/aC1e53KM2jhlQXjdd2eKxuYRI41fJsLIGVLUa3sXLJ6QVBzZAWw67pgulEe
jDeVNcMOmpXJKmATqYzJ2bC52nX41fUP10sJXUSIshjbYXpVT8Luo97NR9LSpwSFXjnVXSeg01bK
yeK24S2TYj71fQE1QUrwEcV0ln6v6I2/CuaDEHoPIccI/+CRGTW1jOqrqe5P090N8r2Fi0c+qzXP
ZUIyKkqQQh7zkmXWU6ZQbxZ78Y3yt1gvIzlCvllXbFu5XLHix9AonLHRNhtKimH1JUtYEZXST4jO
5QrL3OueaFqmuOMwJLT1HlgNx6OXn20r9H5TsSkOEykPKNmHRR8fF1gKpW1oNNCo8obAeWF06VRL
FzYD5Dx95Zkr6bK8I6SvVDRpKVOBi4Nq1YCYNJ3FYdjK1w6qB+gsR+m4oOiNsCgeER+rjXYOZPni
3q7ythXsBcIrFwbOadAaG+DOaUY6HhKnjlYl8qoio69SVKEKpnd4lrm8yb3IgIEeuw56Cwi9P8yD
Xm/38dKz5er7otsEcFUrognKqEjScvdL4Vk7ZDs5juCjg0u2PDeDRRu6ayOjG11k5PY0CEhVAJMO
cXbWw2W1xWt4kmHeWq66N+5rAWgaW1jyBg3kF3DuWTDocBt3gkwMCJw4/xbAOiYrnnaRr4J5N3Tq
BHcoNJpvul+71ov6C6/ejeDCjeAuNcyJlDVauVzHHGHV2BGDvyQ5aqlTKXlux8ZK1EbMvbROXvB7
RB21qvvfV7FTYJiODk8x+nAfJwJz8ngvBz7pEl7aRmeQkbFHJzTR89JD8XxSfOI7QvzFuzFRjF2D
FVgzyGw7khXBRJnrdhCCQbJLUGvp4W4AJeuVosZyK6U8lvEp6BablgVwZkcms+oGi+rzx3roq7Ra
UGMoJmPuZerU0bMYTmfJWZxmn6ZcHcDXxjGN/MaJ6zx/MFrAzA511iX5R7TF0HlDs0Eag/7KatDO
MHvI5tmkCPRznFRhcwAujfvCCWSNAkO84kwxEEC4z7IVmxxPqkPmeEPe3AqcvWYpdHLujsiqLm2Y
fNZ/9pHWG2CFJ98NwCFgIgybkEVusIJ30bX7eOWCpZtBLkgTjtQuY2TsUrr3RsK0YauwLgSvRpVs
B0pgJzs3N7+FAoffmWOgRgbVrd1teYcBp2sGkY62wBo1Y/XHyUbCwnghTP3V3NU2LraoPH5PwKnB
sC4Bm7Kq8CJGPoXYvutSXRNWAza+O30Jxc4lTVI2uJJy8XF6hj8mx8ShFU7imELShG7gKt62oPpy
8h2O+cE3B+/jhUuQrxnmbcjnZkWF4dxv3mYNM255RQ1q4A9LZryP0wZ10ZmW4EWtDQ==
`pragma protect end_protected

// 
