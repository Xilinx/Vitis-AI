`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cCVCNgEi4GU52auCtlFiSuPUQZ
vSFGXE67wEUFdW4WipeikQ1dGNIjntP1EQVjP/Yoj5cHBOaVEFYFpH109lY1viXaSxUucQYThFaI
uOo1Tk+oEOx+nddJ3dr/t6DhWUCq2u7BrLpdzfvspJFCrcAZ8xZsNZbFCu07DhDEX1xUQQrqbyFA
t5723VgmB8eTkPUZi1BfqMQdGq86Cf9AHPUjr7SwjnoIchZgagXbn6NslunGZzMyqx4lQf6RhAqt
NgoDFrGyl9rChT0BvHOxtGrvvVOnoYg0UMBLe7SiLKLWvzfJBbrWjayRcg90JCiW7HAKP8JPkiYA
eDpCyKNGxIisPrn66lb4gvW7Z+Z3krGPHuB951ki6jiAem1pGSChHA+U7VCaOX9kBorR32D+ixFe
Fkdrs9Adns3aJQcLZRpUZ7fnLLEdoao1IX521Q5hdKCa4X7m5diZnBO26d/6cGYY4qRqBOfLDbM5
xn4XHJ3TStmcZ8jLfsUhaePweAbK5gTMc42eIKcyPNlidZ8B+Ugq5MRHpr2mFnGDMJOuvCDsipll
KTE91DdaU/DRWytlBE69f1bO5yI5TnT+A0gMBFXCcS5ZzIvrtQ5+8ABH+2LCzFZgvivt8G11PQpj
zd+vckKK2lK3vOOwA8bWlvtTAY6sZFqv/BIof8Ftu1bI7qHIrmXUJvOBPT6tx8Zrvbi5vDgDDfvN
h0ABUN/xcFAHGmDn9EJHiFapLHJsw453iUn7CQjOB0T5HVsHmIlSx09McG7oCdTlQUKksHu+gmNS
900uxyNgMVfmgSDK3oTDhTVkslCwWdMCZ09uHzjiUUVo0gMAwMmnFEiAVeW/PTiVc5Jjk5GsMtNu
CRPFwFq1JJYuw3gKiarc16WaBsDsIsJ912sQaJETO5L2dxcl8IRHvfNde7/k2xlvPDw9JYB5e9yx
o4l3mlbDELf/hFUe+gF064KmkuXv+ITu5vKTHGb9CAQ3MSk/u5Wz+tAqbTn1oikGU/eeHtW7aUVw
gViaAtpFWG+a9TRqLIWRXu3iq9Elkk+VVb8QG7oNFzFQCUymP0IxeIjEkrzPTQBzsbLH8HwNMx5N
YS0J/RK8AL09fZq0hXd9TwK7GWpEXqx32X3TnHlSrfi8f89Igw5BhBJGap5wEvqdwdZF/ii1iM+O
8dVe4flEprqXAJaSSnCoC5BlIkdfBZnoX8GToCkfdwWEAzRiymWlALG+3q5FRMQ3TsBA2sZFwC17
bm1jyXzKsettPUlv1HxiRRca3bcNKeQfVPRbJymGMzI547mcu5lndX0rknupCjTvn35bG1xZKvY2
iEHohBfuT74kCv6rOfTXIYfIdJrPbpr07kIpPKMaqXMto2BCs5/si2cU7Zxg/p9dOxQJrld/hyXk
d8b1UIh8r0W1+qdblrumT/vERDRd6i6y8jXygMANujCC2grCCXutwExUZpkN0HzNjwDAi+SD7e8/
7u3JCfTy7GBnu6mwPRRd/T7a4YjMqe30GA26/RxBva5+u21d8SnYmF33LK7xa2T6b8Vghy9pEt3O
sBnMOKVLWrqDA2SDVKNoSu5RvNG/y+vavBOfalYyTI2reoXc9/xDOOocbaic+46Mxc2Eh0cxqWNk
VzWh/BVaVWb4Vd0JSoxJW8kI7sgjZZe66X5l5Us8IBpFcRDElfs+HoRDQ5ASMEfZNjDB2LFZXLHM
HBlWM/e+C/2r9Pg9ij27ZR74EPw+XwB7+N7QoQG8T7i9bRBY4h9zUuUdNCov4TKV+SAi9OD95AZr
krTnS2STRKLky0OA7h5xDVoiTE3T2XqmwJTQGzadr8E8/Gpv55mkkEBIByXlOM3/D2X/iiCJKFTS
ptVWisxOD5XCMcn8I4t6lZusj3TwLEYfPQGrPBSrY9GMeGjW6LcQguiz+ny1pl5H6X0IiaNroapH
zodYS9Xfm354z70EGKyN+bzNxdUDx9jbRTeXFTTfcbFsT5IzWxqzfPvrJ3hvtHfMEYxAFHaJ62d6
imhJ1KXq4pmPWPilTQFPYN0ZsJj3Z7L7JGZLt4fmjpJY27MX1FsBMkX149zazuHBRke78r3+KsGl
v9q+L3jdarabAkdpkS9TVc495VUHDinTb9oPhvNmmn3ONJ64aXsPokYiUL+WxEi7OzW5gP2UCSHl
UDKH88KHuu2myWKhfVs8krnefJ2rBmseG3b8az+58InMb/gMWLNhgwupvlgjitFPyLyGjMy9Nljt
Uh+1P5PD5FSW8Riet4wm7mDb8VGfyg/xdpGSQdb30r+xCmy6xv8CDF06Kf14TOzubC/0IBZVro/b
MziR882lfaiDldpuk3HCDFwsRzlqaCuMR/0BMbeKHzS3GCnF4o48vR66i1h57mS2JC+AiuSTU/bA
3jbVgkpY6WQMkNBngq1lx6KQcL2uiS9/R1g0w6Qol2mVsVk2CMHWokQw2+d2bw9tLiMYAIzpvVBs
rxF/FM2WdD2ZZ1u+CNCYoC2lHg3gEjY9tjOZG1fNfHdoVlH9wgpbAi1Gs1akf0zw8EU7tAm46/jz
nnKAraPPvxiCH5PcAnnzPGyDLUpQDrV2o782HxrCuw6ej6UMDHU7g0mzBJAXoBhl/efk+pKJ9dyc
ZFXvXPi/VjvnttoCr+9xW/Xh2mGZ7gkgOa5xy5XKTrf9ujB30MAGXSUymLIavXyP+qClJQG1A47d
1puCTXEDw2xJcJnWjqyhZePjPfDdyutMWykjVikSGSAwqqHWjw0xCOz6LtEo0bXRFws2f2Uhyfll
tkGY4YcSlwkawIL9c23/mCGnHt767tPZWVvR/4MRdIzPXYQMSEKcmUjPwCsgqPFaUJKWkYDivqmn
qQXfE4LKPUkm++xXjqBkQ3ejcNVRwJ20hRn7rXxydMA+EkSKvlqBAzMG0JaCBrcIsqcmG50CWUWV
nFShMNL/b+F0a/6xEpmVDfehYQu0WMQA2iYyU58qrAa41GhNurjRTlWleVsw03cnlS7+xuwg9gZc
q6WDPxDVo4xh5oAo9SPHnu21XtLQrw8y4AzXQMAStKB9RVxl2tB8htEXon09AwgVexQZ1WblCdKy
Q701Oji5dXSLaalPI9oCAz1f/pNXnrY5vgi5iR553cwPclyQwEE34BFRoAh/E1zG1yXcaMWaWEnM
bOhrspDz0cbEbFS2MWa7sBm8sjVBwCa+28scD+s6A7hXRGOnRaE9RCKcXrpxCUWRHhifi4YYtVE9
q2dF/wh/Dk5Ojl/1WuhCzliS54jqRycSL/X9ETsMApr4dPoKjjJ0jfjuKLQe5nJ5ps6JLHCfuqPd
lY4amEpRmTqyy7RPOmMTsnBESIuw/vP66OewsO0qBMgqOJ6dyWQUbCwn5rPSjwun4Iur2kM1W5Qo
2LWqy3I1Fnv9ZYg91gDctUfXmlgSHcVJpvh35Dz8+cS1nrJkjInSzMFZWucUa8tgWp5e7cqwzFpk
eWa/zAwKbJXffVwGBtbOUUWKFHZaM83KLWUyNBynGmUDVTSA2XFYiEzGPtskKb/0LjC1rSgxvxtu
pUltqdNZ+GrV2xbL0/eiAbXkFC5BnkoouHBPd7xPvNfj670b1xgcRB89EgQ4SxdY4XKxUUpyUdGn
BnpM5hYb3CYqA0K+XonRz/A3bThFMVQefiQ25eP5d8MZGtSRl6EMHSs8XSf9Nf7QuG15Tp52V3sb
/aJ+m6jkaYPkogjfvUMxXlL/TGdH0mZ/kjmXne154qgVth3UT41mJdzWvVEUUPoksp7lWS/akN4W
iGj/D+hFUuvQHqk7ftJQ8cnYDNyBy89PVesM8OoGSynaxbGuInKKGolqNGNLri1psqO7ABWDj7Q0
ex6zNDFkX8uiTRTdkR+aF/eFZEQFKEnaDJZzK5akuGdJ2+TeiI/vLmp/E2ctQEQfpMO5dpsIf19Z
DE+/bdssfzZ8T45RNsHdXy8XMF/8m8LaQzRvgRXX8Kl5qxZ/lUeDIhpmiW+SKuYw5264zGohMcMH
/AM6z5UoTSv5TZpnGqUPXXFxexSjDrGuemx2szVo+pB/Z7ukgQj/EpEnrq2uTIJqr/YHnFxjqu9J
fOuzvVe2e7+1zDy/eqHDoTTWmCL8KBCCkuX7IBGRPerviCqwGiR1tAo41+aj20BgtgVPwJeV0u10
ifJ4gk6yrOND5QTRboeu+E2lgLBg+h68ZDlDEkWn3WiXKHGY7matrOrotalMIjbPGFVRGsAjmJV1
vAu1OPoMg3trsULNXyZv5oStpvKiC9xLbFysfGh9ANnWnOfcSfo8TvMCpD7cmQ9akgsCGMisk5vm
iRmdRgGz4enhvWaNNDLlsDcOpapJWaVhmHpGUg99pTCUdkhcAvNR8k1fa0btUovvmIDu44hy6QoX
YjSbTYdN4StW/5gmlX2J6TVz9dVbsfc3Es8d4/hI0PEbOmSHN8Oo+heZuxRDU6U1gn5RlYyCe6Os
2U2Z9t/84jP+E86ltJUFUOsN6lE0tvFV/j1voye7bKRLC9X1zqAdWvNp8znOBT3o29hfLH90MtrQ
iHDYfonhOBMEy3PoYAVt1rRPmeuB/TqK359z2sWsSydGjX8UNo+Jm+Vev8U1T2L4wCZNPjYRCfYX
hlTukKoHC63Ugz+H8kkRy8UsO11VyxOdoCYIaHbOm8YAQzAxTdZFzrHW23vtbeX/wimteDVB7Dv/
oI7UhMkCDFpV6VuM7jsl1doK0nYzIdUss7h+s0d0kHo14/fFkMyzHr7gPA6EiKT0anCijjO2W0vl
FvJnRbvHyuSTgjLkfA2P2OoEoMssTYbMvLr20vOR0CQLXzPDzGDnmuxX1hadHbhHXKAhHk4JCdyP
c3M/VW56+CXH+DshyiAwN306b2kC+bZ5FcNjKbHzznWMtkMGZ6mCvnhkdykePvgu903ik4pk0Hdv
jhSvbilQ9PYkJj/+WpSUCCPaGyNCTIKIOMaq4aMR7AanbCXHPcpVFTpvNy1VmikjcUQhsfJmQjcl
YLQ7ADw6HexOBgSPyy3mpSRumdukFYP83xJlsgwqax81LNy6kkmEyrN3td6ZWiuKjSpmFhaxx9kn
j6XF7rEswquh8nBJ/VbqD9gpQXeXENd05oPgr0Cqd/HCCjpTTbr22AGiMSWHXeNa3VGtJ+m+0ebH
3Rlzr9TQ5HoQzsqvl+T2LfjcTxHICc5LTmiGUXhgBglk6GQ92GdP45GCeWsPMG8e4sxSILplgQd3
aTVh+kEXSxKOqcZkb1pjJAPIhSC73JQp0b9cp5zhoW7y90WKRpeq5iI6JkDtxuUomBHPHb/LsInp
GDa8QJQYg5JzyOpr/7XwtdHFdEWm4EBlSGqkehYw9EJ4eBkD0OrXpijlnCksR8JRQ3tMafgc2wt7
y0d2T7WpjoSl2oNHGOpY/V1RLm67XX8mhPlQcdNQR7Qr4nFpljePjzCQoT6ddkItjNSjjbzKfT5N
aixT/9vbfopMcbAu8FkV9RhOWxSKNB3VeJuIkbcWGucMW0ABBpqo2DScZu5AtHI3b8ZoXn/7jEdY
6J5JVkF5yAo1B8IAcr/GLi7kleDBKih7jnBEiyTk3T8SgytNCmXHOeUuVac64jzO6axk9oPKNdY6
XNfu+JfMFT5UU/9b/NeLLNG8upaaxEjgJ+IMkpxCbNy42Sg5r6C1in3FF0UUKkf94J91vfevGlY0
SpdPa439lVlC73ZEi+SNGGJS3ke/nt5zYMOOFAgu+7Ldz785nUDLGJ5EOfH+3CIJBMz+l4BlbuvS
kkECDHnEzDzJQohEJiCzq9ofnh8sqtKIR5OLgVjYFZc/FhQ3Jt8rGlQGLWjjddK4fSEB5nFeIx58
V371KxXSq48yUGfiD768wkN2q+lqnAgQknGrmZrMwVdTLfgaELHgwRtIt7ZchuIQZBwZhel5iKMm
coFTdw+JwbbiCSZruC59apjEU7XW05iACnSqiwfmA7RSFW1uzmsL42co8wBh2Sq5OOVR+o9s+8oJ
AJ8F61LQxqKUNZKAAD6DFBawNaVUtJcxAJYJAxO2/aruAcsJYoayre7TK+jp096fzucLNgCjA5iu
ha6GdjpbKODScHpfJs06oDwyzuiBEgsXfOaNGrw1ksQX8vkZWvX+XZgeLu+KwTGgl3YJfPPQznAf
wq6BzELTh/aE4yWooWlzgTL/HMsU8ZiAXWFukrS31eX+7DppONvAlOFmicxrzNfbeadrRZ82zHG4
jEmHtsSc0hTMwGh1nWshbBgFoUNCaAJ+B38Ehbmt6ez6Um4pIOz3RsAsGXgMQSF5yoO6684R06Fd
C3gZUamZLVm0pqzhvU8HK9XzPcdbR4iwI8qCvQUZxr2AO2onadlvGYxCvxqP5vgkr4WzBTMhu86+
o1MYZyFhoilVvjVLbSynvcjVwxZeDrbkS+BA1iQve0JSFS2ZXbTaMJ9Gq9WJAYdgCvs1/7tavRTg
JgwhndJex0uuZnHApBjbW6tazr6DiABSGa5vu2EM2RgAMdmjIcHo0fysQ0t2davTqB+B3udO5fqM
gKdrRJ28Eg8aHUJovpZZXwhtG6Z1yZCBZUxCQmdWllTuqmgVqZA6DC1vZM+m7Fm40cjG4244s+cT
FVffiujAaUaLn3NZMiF/aJ8Ur3ef81eDAfs2bcEwtO1nVriQhWN/61W9hJnGA7e272zyNY7Cffxn
jy6NyUqaNvecwV0flSvbH7Z2Jo097r+NeDXxOEmaKjrJ0dOYGK1MlwaIb62P5DMlbYzmFPD0vmRi
jUuY0IJx8/MG3PpiRvwGR5uA3JDMf1ROr8r3UGbEgwEFXpr1HKxW48K6qcqKYHH1znjXW8mYo0hQ
OJkEMeQr17j3ISgZ0S33y3UJs8553w/R0NPi00pgqQK/XVLMKAg5FLp3SNu5VEApGuJWREBShQXg
XNo8jTzJZg80XlR4DWy9lQXL20BPQoSbc93oi7hDScId7pEKLPt/p7eU98zZPO1/mzF1yrs8jH34
W25x5SHbdNu6cp/tlS9DYujIE+lVKSasf5tNgLmOb4Xi6wPVsi4828z2Gpc0oWFE341Fu/+S91UL
FRva4pPjvaQ8mRmEciONIJ/1RYihGQz4J7JD37jceApKu0FX1xsA8YOqQb4hzpGxKysAxRKMWQEt
/reWzdNHcv4vk9QYixQJ5HTR124bVQgtUYITIlvXH50CqgY1bBpUKhhTZzhPziow8cZc+qyN/Pke
4YptH6ZGvY/0V9ypK3bJafSVcSWqZDfDt4fy/QmJScu/0f00rXtx6ao3ipxJdRGVC+pUJUzhbGNd
Ea44KTgTLxolLq63dqrlpBY1DUSxThWEVVKGbpgtBWrqk5p5O7tanLviAsrwUyZfcYFK/Nu/1eEp
K8dZYSIM0V4hAlVSb+t1VJKTNKaeD81hMc9s9clFiGo0F9sIixbDRq6HbhEOq4O9kV4CttEjKFlI
tPLwzQVxp8XbinObXxS2WR+bCP3lw/MI0ieHueN89Zob5MGosk4GRaPkyvvgpVZ7I1JwN9jvcvbZ
aPSQwZ4polqUrInPNYhNj0TXL0csERQDInp4DlWRqtR/PioazvZoUvkkVlzlCf0rBBZ9Cjx0tP46
3Zen5BTffbqshk7JE5TZjoWmyV4Y9DdOxxsKKP5dmIL+AEydIlrDyYryWbNg1i70ROdG7YUlh5DI
X8jgivB65ZuwUxhm4/ehydsdTzPo5tItAQeilWz0N4VV0R5Jm9yCsgwa2Bnxs1HZTIk9zUHwKUMN
zAWNVsXX1C3wkE+XRD2BfiNTO7ZDAJiliH1Fg04xG+sn6mDdfFzcKqUi9e/n5qaAHNuf46ic93sH
3x1yDSMFpzyApKJv2A1w7E7N+tlkg+Zg8nDxb7ea/HBMJi8VUaNK2nemKyirVVwR61BfdsjCos7W
GZPdDrM7DPTqRMX2zFD42fYei7DMUsEVM4T2PLg+SUJ1FbpSa45oncwSR7P3UZsmJzFe9xMpqLbb
bp0mou6SpAwajjokJ30o1aQ7RvPterSaodMR06xZsI1sGbRHLDJhmWRIxYMXyEoGXE4dDZCn+pwy
frrn/ToDH6/utkVILBlzwLv1d7OdumYhDEusB+lt6xdmcF1jSQj5HHmO2/v2lbQNVDTmmu9CBclP
tQPzbe14EtZEkNxd47B0+TieArcOQjTXTnv1kY0slvPnrOR8qLAPeRjswK6YKss35MNitK0LT7Mg
J/PZrVa0FG3pbdS6KZXDU4up5cTNrVFfsnzeC5nUDEKHRVR+DADPROjQxY2ierRuZJRHUXCQAH3f
sieGE+q+xNTwS2Oa1lsgCcpV52zPZkDs41Fl7zbTI1SaNg/T5YwoaGYU11Kw0ZzR35Ay4T7Lo6UT
Z7OpgRAsVzQlwsd8+oojl6GD92Aa2Ok7CsJWojY/FVcZgh+bSCoM9p7hSfehwbAEzqkU6AlfoaKW
tSTtMLoHmCbCyoJXYT12uISQQtJl535TGQC/6T0adU4aAAo9GMojsx8AA0R/TI/rAN6HjUse6hWl
khArI2kE5KzCB/TynJrj5E8QgU6x7KzWXEyTa52XHVSCEtgkZNgV9P8lEXuC/Qi5fVaOB6mLYEag
LIj0hHKRuXOMdepm1I2MXXTR7H5ReXZsu8laMGoIaSN33fXo21tahzegj/7ymENYDU3pmTuyBkWU
QTt7zoplC0suqZpCWJdx2uayxL0eQpS40f6Br30ovEwVDvrmNtxrMgRnDUaUTXeQocWFM+gAnpEL
mPBbktNBG9ufUpz64QxTIL+Bw1aEN/qKwN8c+cWBpDV+fDM+PoOQy4VVu+zDeVr+iHG1aVBERy0A
TcceTwQMcmxbcvSl21Tm7efXcC8LiDwFegbd6m6vLfvmODEeoEnws/JUqHDnzVJE2jc7ga+eiyUx
JgPzYwfLWGL1LwTBebRyAtZf/D9qixzDJDyvN7du3GpKWqd2KkukB/ei7rs9Ehu8F533O0FrriIS
sKH6KLXi/7IS61Jz+926ALH3aZJXumnFLw5g/lgFo1Dh3b45vqj8kKXh4S66OcaXiN36/qZMB3A1
zdew6vM3v5NKmEtLE/2tfCDZ63GCqsPnEcqLzffk0wvq+iaaIcLrJjD4u270/OLgN5k3nCAF8KS4
qU6HIZVl0Qulo4VNXFqoOqQV/6W3KP4zEKwehovOAAjfyDVMKry5qYQqKppKdhBggV2WXiS9WjOc
PiSDFKG82H0PA34yiq+++z7SxwzVY0sD6yBwKADBw7NI80riCDd2F1Z3rrmLePYLVelAB8ZEKIah
+5NH2A70x9mfuX042dFPkRb1eIdAf7uREb9rUPGcgkw6hXbFrh+GYQ/KPK5y14oiLydeB+D5z7M2
lT5oM0HmEQSHTH5Ci1PUxwqFfA62qfVsaPfB0NIVYHzrk9/qGIBZiO0EnsfPP+4GQcxjWB1B3SDG
3a/x3xzV3udjDJed/w1pjKR+X7k3RVHCkn/2V2M5ZlGJZrcBJZMoTwwp3UjjAO6eiub9lbkmfu9C
kW/xuRMS4jfl+W8acou/lN+q+usvKZ1cA6Ileah6asErhnufldbeM1UUp9Z0XL/xf5gKxJbXx1iO
8o2kXN9hgshAe0O3H/00FTDhqMUxkHS8dGBZ8/zF/5lrRSfV1EnI/D/jSRfEM2dBjhGx+BcLlOY6
mEXBdyt4M/RYJ8wjbXjeWegm9IGiAVNUYnfdTIAyMxjXTutK4/WNv/FXywpb8g9ZnNL0P9jMVdwS
tVYzOzMQjVHOztZcBbCCq465s0Jz+VBfeN/JAvE/x40U754lI48poyvqzgSVBqHpo8pUxk81dWQB
0To7FDj0ES07NXkXOR01+67aHWa5Y1ogOFJNHYVhVYRtJrUM405khLeoZ9oRLtO9iPzc5c91khmX
YqjLv6G9U13fjPnsJmXQfB8kt6g5/4hPx/iunsF3rKnv0on/vRIGQ9XwGXXRwsBC5f2CAeon2cQn
7iEOrP6fHzIUVEMlWoKyzlDxydcq66jdEWchouVw+R+kwF5UoBDTg8OPp04wZVHwZqqYY+coDPUo
sTgfT9FCo/PKVqLM6CnUTWmg7d2tLe5kn1/KoZHXBpO8fPu091AB218Z1ieXkarsFLnZID7I1pY8
ofDdvyAsxKK/fbzDiOONgE4cmSOXa55qHnStUuAdfHmMuhivvbQaOdYyTIwhMhDeQVLSkptSHWqX
0uD4zDJMkp0Vm657+h2B3rb6XEOfl6zv0p3j/sNXlk6SirwCajsybOCEHuHZqFaULamo6ZTJcNKH
cydVjNmK3bmOyqkwoq/giRGrILFuKWsrNPqoS8d55y7GVmGqqXcmw6uOsOX0bZiG1sKfND1zHWPC
KS4KtBC0h4SEediWYZenRLSbBUIO2pSai3MCeVSRuODR4j09NezaU3MoFjvSpmkxOpayGq1YVA27
ejMAU8a5UW0+HfpEmxgrVWM/Pm+uYhZ0Dnt+PzgE9Nz9dlP5LZq+D1yB/Ruxv5uu8Xjn1klPWUKM
0Y+jRVLNtaJ5DfqVNIJRfq5gRvj9y4gdNcorCN3x6H3cJ5P6YyAylXTvAGK6vG0/v8i9SBlZ9weQ
6J8BK5Dt3LaoUdc568DKslMHVdpqcg5ajShopuacBuyrm3YJwwBnBQM1B6C93De9vgWdK6HKrtWP
KGyPhh5ojyW8A+Hp8Zobt8qiRwr4rvq5l3AdztO6PYi+oYo4NgjzSBOTUuR0EzZfeywBCpOiraYD
qcK3KpLKnU8JvY8apLMTMYoyhV2Lz0VNkTlhTirfVlxr0SMP7K49TSfxDI1CwnIBWbo/9cOyMNEE
ljrVsOgJjASPkv6Qec0O1T+DEqWqz3dOnvherxccqZgfaN5sDBy8hdskaE1/B9V8gHnhC7YVPFNm
sm4NLmdV9dFAvs9YpV15m4yW3JEArdV99BdfUsobbMJg45QYNwhrufH83uqhnNkYFsqyfD81PJws
GT1zaQSdaO+R5TvCe5vZtIMGjZiUO7oid6WxVNsbEhVxwTYlbdcQSwUZGtB5RU5TiR91JN4ZXgCK
CTFTsbw9qMvdJKDQImAxLMKRZHujHyF9dDqASpyb7s3lyJeXh40WmLbNJZukNiYlW46ImACflwmI
Xus9OI7l7p1mc+kAob8esw/VFe8w11F+VTB0sjhTZ1RpgQy/UBbeMtNBJfd6KqtF9c5GzPqMLM8f
AKXVRM38IT32XOU56Ckn92p/qpEHayDP5iuMWjO2R7Q/4Ll/kfvxS9lR7k6u6TEiis/gD44Zpegu
6KwdCpvICPC37gRggMXL4M9e2vqpJwDWrMgyyjxEHuzNkICWgIjtRxUBM7Ehs33eLZAS8kKMB/nX
Ikm9HCvUbtvx/9axgic/cunJnMfuQQmbj1ETgn7f9IyxPqhGLRnQ3QNPvtKEUHar/a06tMMl46UE
di2IvB43QCIZIFmdx3WfS1v4AxGqiwZD1FOpcV3Yj6qN+54KENb5vS/QQXug4nfsUGHumwlYSZcs
TV6ZKgo3PT/SAeCG2+JdzjhP6fazo1vf9t8+r5FVipiGc9kxNLanbxr73QZFMOH3BQgDLg+8S9qN
SFM/s6bM7XhZ7iOEqOpBTKScSB1puHMtIejltevK7dfb9c1JiutZ+8oe2Vw4YWejXHGt+y+fsCUn
/5VjAG8vCOHUEswApf4HwRa4218iuCVRM+SSh34rl+vGkbnlzFdazchIMQWwlRjsBoRDvYK4dpHJ
U5nIV8od2zf8IqriVBiF68BYaMxqHLMkeNZ1BBp2I3hh+Bhu+H1YAVEwjYSiUxTANhnnqzcnT08c
rZllzlNpE+GhGqB+dVibvgiELb9QVzKQpiSdiT1pqYGzO2/KC1MH9BnzaSOh6yd4Fwkz6/v6dbXH
SDLs8HCBV/F7BVU9dq5f68ngGvtWDJFUqUbtuu8Ja6/xMnOet5Y2OIzfwaaJ3wIda4Sp6fcT7/UU
dl2CavMv1fagKWpPQCK8gnBmv72YF9JeDKQvbCgUycOZeIT9UfZG8AihqGwi3WAXT1Xoj08HUaAE
GPJK5GWf1u/NlJKWQfpqpS5eauOA0E+4f2Xthp2oOuMCYhf9zgkEf86sXm5+qs9TpmATH1XMSiWk
3SpUjXP5eoBQf6V+bBz+lBT9H6ifXf/dp/3sTJYHl6QetmNeug7XuGkPCHDcB28ns0M8yqmBPjoJ
DukpgFeRFapOytzAaWuLyMgM8lgNqeLYVC8rEKAmXiUlbF+CBdeUmTpHt/9kM1kpUHKT9HuwxxqW
85z6JTCo+xtPZHb654jIFake9wKqlgVXtN0+/2IN1pPH4R1Uy+RRZk9oaySLeIgG24TU8C+JxozX
HRIjrQUbs463dRFdENxuG8gkV0fvqShxEIb/mnRNRJ5xwEVgH56jGgi4VsD7Okbhk5Cu7ZOnZiLn
rdV1WWdxsgd1BaPgyqneWaok2QDcxTC3Irk6CNa/oKGNvqnukKVUqZ/yAw0JwXvEhRhl4IJuwl5f
QzFG/TaJX3V/OkTqgc2X4fERJM3ulgtXNJusX0PH214IIFvMvv70Z7ZTFCcwRckZcsfJYoWTSgUj
86w7EBA2Nu/LpVkNc4l2Q7x02SkYVUA257MU6mRkopQZj41vyq2TwUJjgqfHISvgkdaa85rzGjbm
AwX+Pgs/BI+RDJEQyzuEVzdsSdrqaqbJs28fLmOXNnP07p6ojZ6aMo4NoGu2ZOpgKGnrLHFjW6BC
UB439avaoBfGvsWSVLfTFWoa+E0j09xUHuXpx1y3CgNLlUXk5l8TjYFOGAoRi63ZKOF8l/cMll2j
HMBMLO3oH63RuHboAP0z7R/bm6w7sYQaFBsyf1MsSlY6YWdxg1PCq22nfRTREwfwZIWBmAPB455a
4mMY5zd1PIFijNR1swVNjCrv8C9Ib9tD0Zh9PrdntB1T3tGIMvSKanyUQ5dM31MiGQnUpe9209Io
1xg51MhC55zc96/98jzoLEs9jVaj1zYf+QV8T2qmPD/YfaDkcByFDjRlze7Loeo2ghlwNH6Q/+h0
3lCSsb0hJBu2PSfwJerq3LoVB7EFs3+T9M7EsdQuRt5FEeqDpNaFYsB+uhVzv24NgvWRZxdGYb8G
KzGMjzPXiA3Dw/oagjN5Q1xnNjnkJTwf3ngP0BB/8R4F/EEGdcpcFrtvaJ6sZ6xoqrFX/evH8rPj
1EQFtc7B4pygsnXabt0J5PSRbpbw6mDHuJfGspvdPF5e9dk61c3KyESO+pfV+EP9+1vITCmHcfTA
fY7u1RvI69zCSMLY8K3eNrJ9UnQIkuRs7v4KHEoZaby9z835U12U5q7br5DJd9kpBw5sR4UJrLPs
4kNiNlh+FKocvcTNkCQEWA4UjQ37WZ6HMJOpbd7Svp8Hq0erUsnjNhVNP061t/Y7LffKMeVogyzW
X2YPNmdWh1xyv4EsmJOcG8QzWzkZDysqbQCfKoMk9Ci9PUvyKDUUvZGOCN/AHALnaIYUsCXoqayt
sFI7XgZ+ojE/RTHCW9aoxMIUF2NWrp/7H2boFh8QVKPftor+GgirsTqGvSwH4meJQPzCBhvassn1
S8GPsBjoRqI/BbdLi/ab7Il5CVfD1fPZYD7YNPyUtt3lrmPNyGeNhGNieqXajDQuvKWh1lRIihGb
Iy7g1PDwOu4m4ODjN4tRrMHAjZZl4g/cRstRa7Kvyok/7MoKmuDqC5MVNzouatFZFbbpUqVwoKDH
amQr2E3Q1w/PhDIw+36OgrioxQkrMZjDPvGGRjh30VaeOocOweTfg43bKKLgBRJGuqSZdIUt2uHl
PCB48zu1paCU1h0kXWTkemFDhYrFww7g/dLwjoCKg5HO0DW6YHmljljab8i129qAj1RKMEA1fU1F
5EMkPDMnhcCyxitCeiTGISKg826uT6u6B6iQjl14zKFXP7iGty9a5KYZs6MEo8Q6A0zkFVZOM4w2
GmE04EDWoM/tAoxWFFi9qoXeIS3NTzIx7ilnHF5Ooc2g3i3kvl449KZtS9zIK1JeUVFpmCIlyLH7
gaP6cSN/cS5UIdTLfV/63BXTbd3gjXCP2Lh/h3zm21YNqHRg0rHiaFt2mb5hqbGYFeV4Q0BMI5xm
mfzGFcZ14/VO5/tK55ut6FkCCqZ6tMHMOCtn8mZV11anC7JLCVyDA9NmQ3q9s2rWssbYk1pPaQSN
adiALuV3i3DbpJTLg2OVpPq7ryDS24UGq6MeBEYxUgvpdjxOjx9QQLMZMhr7IAA8fulwktbFLmdd
dTIgfLm2hhDqIBeYYMO1DtX4q9vGZXvHSEmSS1I/yIuUjlwWdjYbUOakz/Ves7WFZ0TaZ9/z+pAR
NQVORtlHSM8sA9Us9wfXLadUFBOE7z4/AHic7JkGOv1ikyFuELXMdpx+jzWlxGI9h6SGBBXfXilA
HjliXfBdh9T0hiERCjvwDoKrxsWET6thCyLq9jC3dwnx1Y3ge0JRbhgjeS7hFWVJ9r2jWkYA4eHL
fMdoOU1B+YG6vQ/chFePSLsk7fwk0U94PddL0hdH2dWCfvbQOSCRqGhOW0/ha8tTvLAAyUTLUQuH
lUAPZ2tF3dQsc7NurFWU9GWcJxtu51jdZDSkFuiZG2sE+orb92tyYQsSU05iyHzMKeaUgVUlEbGI
cmlVscISh6AFj7sHYKGNpTz9U3B+QkznTATK+vpQQyH1sUvZlYlxcdHW329m58zbRpfD/Uts8TN8
10BY0U6/pHpDTiyfXWMUpbEiSjqYqhGNj9vPCXHNccHDyvVeLeeFoRjJa8dNV8syFhcxtRwqiobI
pGowsqfh4BLFYi3LerFOLZA0hlSV4uz0uYjZtxcWDOl44cf3QGz2W5Zq0NcaNDqO59gkcGAcLnd7
fBMprskxtYKO5Rg60h7P+4dFtWWNy1fx/rxxY0Cllpl47mBRVGrQSkp5rv6d1qJWjRTn4AqACYmR
XGNMUN2RkFor5TIdMC3xo7p4akCNhnq9s4FflCohlEVt4ikT/uaToajDiK653DGhKJE52x2JRbwi
KBFaqzW1kdGsGS9ciR/sPhFEaslFe46AssPB1LoQqA0aRsOzOeT17I+UIPtvPbtoa4nM9QAbLEUT
x+axXmwIRYiZNT1drC5L9R6lqy23aoWbcGqq4nJJLopf22TUAlnrDw2I4jra7tF5Ax0ymLEegjjJ
j3gPPDZtQxZQIGQCNG8A83xfSV1ZODDS5mO0b/9mTg9/lsb3KkZ5qn90hGFEhyxPGgo3pXI+sjre
LgiIoigDdkwVnWptTljdzur5+mBezSNdNikO5nEuK9/JC9nzM8a3OIS7DvTc249bdq5nnoSSHFUA
gvubs4iZYm4bUB7GXg4wdBNVfg0yZkNB8r9YxaUP07nKHavgcH8UVKprieXEiLBirk4TdLiDiA6p
UgApZTNHo5Paokr2cbbIcQhKA+JFLr8ePPWLXk9mDyTsKTNBcwpNhnDYdJ4Q3RSEwdC6DNvogdQ1
PrNZk0ea0HI/MzWSwz0XLF1kOvAxkS+P3U8C81WrJ098XpXgJb9fmmVkaVKaAjsvQLsQOuHPgXm2
EMVjERLtwLsscRZslmpaJ87uhW+Ec3OKKHXIYIJUYtAK+V23ohocTprizBjykcoETA8O03qfZnKX
CBxMr3hd3iBKi/Cqua14nP370gTnxe2JA1GK6eR4mDckWaYzFejkBIMPvGuRYTbyBf4A34cq3fW4
Nv18V8XelG4/wxUsvSYoVti9pQ/l+7fqqBwsKKScrR31tKJj1A6AAPWf/TvD/RKxsjxp71FPXsG7
N3olP3o16/VtRWdteaDnd8mdEgEdwN6HuXukByiwfAXf3Ut/3KaMWDauGEc1J956eKRkxPoKqU3w
LedNS3PfuBu/HicIrMumrQawJdl7HHloCFwTBqyriHXOkjoMIWtMdyPaknyde6ca5VwAnXAw+V9r
LbXV/z1+E7J3wyYTjLbLk03n+iLZ3J7zIBbJQrOc7PUgxLLeLHGIOXIIIyzLIc7nlglAcERw7K1o
maA6lX6upG+YXUN84n5N0zj6t5QbsOS3Koqk1bxLpxYCowW5He6K1MNOwVSsWsXDJxCHuS5TWWQx
IUoJ8ghbF4UnUSCmwPnWHf31OpR4i28BnGH+V2w2EoGpaaP7sFbGH+TCjQ/RASVmUTA8UC4Ahp5f
dh4c/d2rGblysJyyTk9HYao9QO+/hvs6xWxaW/8cZxMLOQJnbbJv23AtmKn/4xLszVOHIrbnY0r2
xLQH3zCJZvqCeOQZQRnM9ZuvH4I3wYLQuj5x74A0X/o8i2x8ck6tHBoxPUKnxlqMfYuT2lde5Wlf
+OwGrymQ/6qI3X5ifk1DMz3loyJuGlM2n2US1GPX0L8Oq3F8cNJ9Jq8cxn3nQOo5s3pEFxz6LyD2
suA8Ex8TvtrM0SVlQp7La6eoEPTvNydvWSrUyQxy4lexhVepyiIkjiUyqlgD44gEAnmiWEA4UqHV
EXNiBogd7raMz4Mxe7a7S/BZ+SbXKI32XAG6l0utxG88IHBab4Ao+8XP5gMMYAO39O+ZhKalJ6HL
hqGRaAVHc3rJ0BzyWg123HRLTwldvocnk8yoSxO2B2+3iTfjYVE4ItyrP4zioX47Rbn0iRh7BMxL
tePKaJK6/q68IJYbnw5n35D2X68atI1AspuAOdPnlzxhDlYdZM8Cnjpg7/gfP9GA3SLyhyfbPlTw
6ngoP+QVFbQMJuDjnfib7ZQsdKJzkjtODndmyn5IsAEWRVPzmRZi7F0xx7PEOUSLAK222/cPGh7t
V14ntZXl8CnXHpMHE75uLq0O21aQjbtARtw7j2hSaZTDS299CYzRcF00KufL9lyqMe4UJO2jkow6
dxD5ZoNK0oI3SnCdAacALFA6lMjzQJOn1ec06JZvMKX+/1PcKpzynPSs1A+nuq1uWjNlbXGa1PLI
QlFuw4f5bbUMJDcaOf8/JjpmaX1KhNz9pKJls/WC9LGFqaaVKxeNrfS4q+sRX2WbcbCUptkdQdku
auG3iyZXQE0cQAXFe4Lm/pk5/SjBnBC4MD3jjfRZqpoP92920JkwkFRu+Jf7UPiVy0q3EPWjrd6K
V/2dZeiNL5y2O4NfY4YnRfnOs+6uAd9NaXg7JTkI9D74ZPMMgeR1t56TcC4bzah9T6HuPXxhF1Ja
o9+m2mgtRde73EidiwaGlMPj6uBxQW6tzUU3wlDfbZyjhPxWtlyq5UvSNtNu8EiG2zrfbqtE1xFw
qE/VC9w58hIW6W276AVR0oPgfX6+czCSgr8sB8HAq3YGm4laxFOUNS0veHlwRgI6Obou6F0dR8kz
EB0yf9N5GOvAIbibbJ4zJd53xiGzYg6vLGM6oZiAJ6KahzrQOJE43f6hoy6DjXakrhHAsA4zt77t
QZI2hVPwGAfu2D3KvCvQop4XcGuMFK8A1Yha4+MH96ozxRdI/RyigZgvQKyj0H+JJqiC7Dp3gpJy
/5D8/Gpk3vQFRwPOL+kgUfaN1y+7X771J/M9aNrt16S6ZpMeXINgYduYNF6WhjDK28AEr2pYCA1Z
u6wLd7BJCUmA+eBFHUFdMD8lI6EqWK9mc3Ju3ph52SqR/Wi6gWApRH3ohpW5upC+MBLeDk8EBAyP
pZQ8zonIuJa6ByWmnmadlcLRFObw5x1mdjY5+/nRuPI71rd+gA61L7vqu0xEsfAFBBuBaMZuIiAH
w0606+2f/x2l1XNT9ZpKzNfCzpBjGD75uTxksm+7JoK5Qqy0XnHvgR5Os2zJtE9yePQ30MHGN/TZ
RAu1BaHZ3LYkHamxXjkeVs0O8V0g8gpp6U7qWwlhc1IyxP7Qg6SDzRjSasXHIcweiqCoT1d8lH5R
uoFmtBbiCZYQztztM/+yCCJ/OV8OopMl9yS/RngkW6uQ94whsUlwHYeymr2UijvzuJfooJ/vpyzM
JYV20Dz6hSkOx2iKElvz5hAl+lUQdSdGIPiTiH1liS3nUyDoCOdk1CyNDiC29Wqs1onxkcSj9Ztm
nWAXMhvYYbxI97K+DCl0cFFEeBgovsFlTUiMYDch9jqkpMl0Yo+JauWPQPsoIov34vckx8dCL1HI
5a2R2nP0Ud2jPIrFIu3f2FpLhQdQFg7gkcD5VO7eJCAPT3aSbRaXwf2hwKYaSg1chHx+I2EkvEV3
+n6utV5Kqbxa0ZjivzU9b9Xuv6OyxwmVfngL0Kbo8JBAdIq5s3xT+ORj157KelfAviosZlFz6Ti6
mut4OTfd0yKWwGUAhUj7H8tPWumiZMk6p+XZLZAiCk/shb4W7HR9Ffc7lQDH0ReE4Sgwm0Boi/32
qClUz/unK1+6+xqZQI+jMAtORv3lwDIl0kwg46rfBC+FnBJjPLfLa282aEFOeljmDzyaJhjOgvMq
d/WygLKIJtzO0gu+omDOvphd6s4l2qg+oBicc9GqzrPhHvBANAnRIdDs6B5SNXk6PIWyE7x5t7t+
2E/gP9th+X8zHtVdmLoDtHbbYYODYrEZ7LhgeR8iqqAPLxpkqD/vD/ghtAuhywU8Y0kB3GcDWSlY
U/khGGVQQNa40jKdBe4Cmob9lJsxJQMGfUtA/GvsgVW78xoQG1uTdvpfSnAh/bOQnaa6jnvVjYfF
WxT93dehGiZD9vHmy2E4RqKDvnLEKoGGEPrnmu8oPa+wIlBMw0K6aaRi5vWlRFmJbynOlHqKfdqS
VbuYbE3qsKZL1h3c5vsfrPyW8GDvowiueTFweTFP7ct/HQBek1mAKzZI5fZYUWkgXP6jD/KSVtAh
tmP9dSyVzFRcjFQdxebnigKijZsu5djLw+D3yvkheKi06FsFAT5ZV7oNPeGPXWe4yCaXs9KgIZ5c
z2PKv/2EMrsqHY9xsey5ydyUaFGHJHuw1QtKM7tj7foGolsMUc6NY2Z32JOayFr54c8SxZUB2k/G
2iCEju6ET6QnZ5/O0GhfIx5knMfUAJc1NgAuZaPYKeFBsDageFKBSe3XRjlbpWLw3CzZhCB9RHV3
rLNXAxM6hu7gAfEXw1di5l9FNSmAIvHg92GlOVBbvukJXf+G7TUG5wYqOjRhB/2bw2SFIsnHsArB
cFtg/zSq055vt3Tn91q4cYZm1hmpXsdd/lPo/MbvdrOwdkH9f8nNNW8RpAM7m8Rz1eL90GhyS4lr
q7kjWQXyjWxJ+I4x4Sk0oynm5ZeaccE7lZK5kwsJRI1dM8Thd7wWVlVwEzb+KIR5ei2rvxC5EoBg
xisfyRHzW5ZeMf6vsePkuDrX93lCeb40s4oAjMDK0BwHTWImaJ7jUdhqxiAlwZXYD5QAFi5uOFYX
6ZAUvu4pulTLBYGfUA9kDth7ccmSk0xLk6uLJHqPLj+bvm19u3CRS0Hass6L5owWk/pg4B06aLTo
jny8+eArlwc9p/wlobLDTQ25tPL6kenMAxcsBhKw9sJjMtQ09DNnCZUcCc0TKICLET6S8QvFw4wb
z9eyfp/WY5O0uzdrd96WkzyH4bQikTffe6bFo5k6WY2mjFX76X2PGwXfVCXhFhfEu3WLY9p1VMEC
ni/Keav7Lxqpy0PjMGJ+rtw+zAOoBaSPfj4rTXcDHmNx4MFbf+e/cszFmnT8CzZ/2qzbzPALOvC8
7V1y7Zh5+eXTtq9Aku/os8xFGlzpJJbmKytRFMKmM7A6rXxiON9VC8pht550qqejTRIP5ynpNn1q
fEKV2HEcF3PoIOxVQJugo6rXkhFtm0p/szuLr7UzfZkLT/gVCDlQOSs+cAsa9NuIgJkWJRi9LveP
AAwtZQIw9NqW5VvIvZRYeT6mYPheyL0FB4Md81N2hxQ2jXVUkxYcFkCw7kjZiJjjDcpZuadNdr/x
YwcJytGFs5EZRFa63dH1jpnuf7q+qfbeI4S14oN2pjHr3NRfbZ6VgZNHaFB0denS5T/JJg3Cvhnn
4puKLUcAdswrnNwgwjLfkrkagwDPah36m8qygazxSzrsZB4W9sChgX16ypZG2pK+SAtvHV5ncR+D
Ozns+3Nmyb2cHFk2Lcu9bcz34mg416tFE9Zse8+86dCKTQA0kbBl8xNblfEuqOy/PF0LwKQSHakz
MD4qTSHNUr9Tyob+aVdlpSnHr0IfRQB1QIaGpW23HtBsObg6OMfrlSYS5hjCXSb3e3UNFYIsIE9H
8w+ZXkwtRNAq0YMMXGmUI9utiFuorw4x6grC8hl3UUa3fDVK6KudNM8nOzMQLw8J0iUQxMXGu7/X
luwia8UUNfmqGfE2YvE5Xmc6LqFV2k2gtd1NHlrBleFGng6jNGEnVCCoT0docOnxyeeLtS0yOd79
d1W9qbxcyf6n0rBHKWzmlWeTfOhjFMRK3TfJ0V4jM2dqK5p9VTA5nOcS6MAmdjK16v9X6tvFPApM
vML25GpSnRp4tRC78ajpg7DWRaBAUZwFOFkr4DuaWNdFX1S/uQbDBXHp4ursllCiz11EZwcUsN65
ZG7xGN+2GZcMxVaa5+yosaCQ/Cob0K+Dk4Rds5b/Tt8zpyMYgZFrHiwIF5SqqPGWtHTIzrv2J4P9
f2F9oaWYpImg0KJFELi5dGpSa+ux/6Js/xWGtkEpJm5xnYFV5un9yspOdpaRccJhLFFXiR/VHYtT
/hNj7Mj2k9HP5x6/g1x5WgaBL23f2Z168hNJgt7INyTk5Q5Ggiig98qW/Zc4jsLvdxpH4pKXBUQs
vs1FMSyQ+qJd1FogHquI+Ghj9KcJk2N3cF9iGrclBJE7L+G8nnSjOoI68d+Qw+LKAFi3YzIYDd2O
7xSNHizTbImiIlBaxFnhy7KEJWtl503rW1tiYfmFjWe7QoZotmWY4BwE3I0KsKkO5L1mjdr3lBGi
EKIE1i1X6PEQeeDljcT0mv13dQUKb+MXYxNgoH2EOZVHHCJF7DSs1C+XiBvh2l7KyH/uQePPNyex
lwGpHvOTpdgOCfOa8yav5x10/ZrK6WGGToQ33LqJkVOo72fkprab98CEdOKC0d55p2fvv1D4vbA5
TSoi3MeRu1MK45o3fR/bfrz9ZnrIvvJtTTdhmF/tqWxIwe1sjYX4Zyxgei53E+pk+hplG98OFnDQ
Hl2184nEtRUkjToPpz5P5jrBe7cIoSzl5mxeduTEvj5n+Tym14fHq2XJEV9PBoXzMDhYjuorGtOU
FpoH9KlZK+Uye6PSNlD5Yy9ETmIPEAAI999M5DeJfCml5SUMnJCtpypHj0qaqVWZiqRZuKIjN5Ae
6qqOKhuIgA4KaLs68gcPGtUcIPnjFQ88UnIuTboaUmOUjDJ2w12QAZR/D4q6NrOdn9hHsd6Xx2tL
6I0slwrjzTLTVjphp6AsvDXTQpd8ht+S8rCfZvwdXHCRJBDtB7c6APPJzkKxQTQIQDmGfdv69Q76
5OzQygrXmHJ3zE8/Q5QkTame5A/s6PPDgeUK5TDOf97P0xzKAoSfR+OngQIMDTsQj2IR+2O12B9I
lKvhk1v3x9pOWPTyD5tUFD2tlVISdJCCbngqBdmrE7CNyjihwzfDuuTiEr+OyurnRInquf2NoG/r
wl3pFc3IzBNgB4CidmhKenfNllegVyBkUfzDpm9XGTbOqoCovsUUgtwWqoBEGi2anqG0Sje1YatX
GGB6ul6SSPjmAceqSjTfDhodvhtiFeQosjdgC2TNUj3BWConZdVYKBiTUBezpmZE9DxfAjIvsYIp
xtQ4WYiH/5+443jKJNFchx7yijv+QSwc7Isetwtbtcr8611VnnbDbx8SXubOfWim9O0P9y+v60vc
asJsjAgkh/7YW8h2z062lfMaeuhCp/GlsIBUObb2kHnCDQFRlkCVxUzuC+pi1p+jMlaKlppSF7hY
OQXKWumAg2/5GGq1ll2Yorsln8swIySnj4SPL1WBHAnlM/loSauLkCmyLDNktgQ8SQ5hDDwKMolW
jLAbg8aPKtpQiRPopwD4xV4gznu+64+F1VbyaztnprvEYrd4dIXd10Y96OqO3u5n+TF8WHhvESEc
ZSytIrJYDW+35Ae4hR1l1S8MwCqR5/mUCzLnw3EmGiNQAKA6wxERTs5TetuP3vm7OCu9YMw++bCA
mrjSadaeUU2t338dMm1CpiMPpOEWngOceamj4wyy/1CLmefUzICeVQKeRfk98RLODJeXl+jqh4Cq
GU8/upPYAxW1oseTQZtN9fFQjbfF5/gukuc0L6AJyMtpSKJUK3Ok5dI4s/ztvY0KuiFhCLO55Ydg
titEIvSStfnrFaLAT7efyEZdA0zdktv0e7ZcS4+7+fWFZ9Zf8Pfb7WupIA9HesyIuQLm/gCE+QS1
ayfn4+CdrQrRAyx61Mk9AX1UoZOYGs7HIs2L72iqQOUHow2/2bmi112376gEnK2QjC59tBtkGJRW
35QL0c/y9fgnLpFrPuSdsLs14Dq8375d2nRcuLRx/4ws3Rc8lVkt/1NMt2qVe+/f9WKEgVq6rUtP
uYXQyNRIF/USogrAR546uOg0AzyDwPt7zyM1S6glfdWKlLJWGz7VQZKx3WpjemSJKlI9qrKKq7D/
IJPGIpotGf7j0PtN/Q3xhKmJwPw68CjxiFBLFbtS60kq6V6Q2BFOEOg7pJbGnPyf/40JgY8rr6S4
EgyYfOs/GdvEZ0B3ExoW7hyrmAQAT4XxhklZnGAZFe8jCTsZx0iZ+GF4NtVef698bPW6zq5RYcCu
NbmRR4aZcb8hRoJE7s5gYEcAsf28x0m/RSSrh3p/g+6AQkkzyOI+BvDRqm61aD+U7PTZ6PLP9O/t
Q2B2ZEz/ws8xOHsz7O1BgrnHdPZJCeIPsDbHi2CeSritTtLQVRRvd8MnoAZcGaz2g6j5lxckHMXv
+KfKougME7R9oplz3LxOR1dboiEhggjkOKTZmHX89HFnoPyS7397Ul/Gs7VW0v2wVnUAsbnw2kD1
nBdU+lEmZy/PF5vWjjAuqQBVYCCuLc3iE/W4DqdlxYDdHkan21Nw9n9b+SfeHouh1lBNOJWD6x6L
mr4+OmjFUkRZIz6LB5WlOfJUs7zA5N60lAhDZ60w8fAn5JgOfdCAGUXkVGRdDhIJddZ48LRSZMYL
VFc32m26hwpSaSV2jbeq6RB494NHhpeZW67tOa5R7wt845ZTKwA/aoBdwabtRTAVEM60/1qOopF1
jDrDA+O1SHpMavmrJhLQZcpq64WeXK5o9iUTA6pNHexrOUC7XsaJt/ZGsq2aB92nXTICQW8Yshxr
oN1+jOXhe9I2DSCZ2pAVqFoWgUGYyuG1eJsH7WSwtsknwVaixyFoSof5ce5BGb0FxLfMGSDbpY84
ebmsUyZkNi9xLskIeIdkclep6voQqniJMf9Fn1a/+BuwfZQ3YzeMtAm0Ht4lJvOYjxDCsQD8l6Gn
jliI2Ab/n8Sp3785GPWcQLjjqKoBnuH6mwrfQmCclyzT6UNzUczjkNOuvhf3gdcnUp90lc7y1d/q
dDtjb51qJsLBsuAlka8ibQo0NiobUW8/9NfOg5Q3Ol1GTD31EfLvgn/mqRMfNqwsS5spcWPqEQUl
2MhmoxACV/1YzV/Wn76WFrJ9H75mHzNnfUvHmbF5Q6OO4oKdUEWMdFYivsfh/Mmvue76xbjCQCu9
sF8onrGuT6+7LZ/kTE8gAM1mmXw+Xcm1Ya3UULGJXx02flRSYhy8WQpuo+v0K/2F3Xiy41iJmwm0
3Hy+ALxmxP3/1csLFqIQuritV3nTfJcgb+uolYC1eqkfcfMJYuzYyeK3BDZbi0sLRFGIrIstxEaO
7dg9sGum6pcRHLZG1wzfYeXbhUDiO4jXXWNRUNYZ6G7dt/N8M2XF4zyUbEcACwXv9ihoKRiH12pR
7EHJ79rnzKObLU2ojZBjVvHME7akRYxONawc03fxH7BJpKOESXbghpN57dObf1AU9jVBwwNmXXUy
01aqyZDjoXZOwDC8Bx9BsyO3QcYKcG6WsqwS971tS/R+9YPz31jbSd1wQytxrEKJL7FA+PKVyWxh
8jpszibSxR/O7G+cNHUwplUEl8pE48YYuJqBOyykxL2ddxwYjo4vpsPAoRex5V75CHsJ5ucA8G+/
NN0G6HmD78x/zyjzylI0VD6Iu8B7DDNEHC5wJP8ZZU1be+NgjthGkFi2ZzaiMzHoZh7fQqhSVQgy
7pRiqtQnF1Rpim6zf1vHRB9/QnPSbkLmbEELByddud/6ijzb/DKBmfJu6SAdcjOJ7aJgqf4ApXZj
vxD+VmZdF1F6KsIYhpMy3Lqkf65m2bX0vQYa2NO65mwtUTeT9MUVIWkbV/Mwu9N97SoM4hi3TWS+
C19pAoX0kTz0zCymxKAmbIFahRLKXanyLLCvMPR/Y/nOvBiAaHDFUDo0R5V+6F/fIxCD4vfg+EvR
DZXqsDtTCa7+dqSDOkVa82X7MDtF0r7n/pCMPw7sGW0A1CbtUGAncKn9cwYvX3AZNAX8pZqdCPJk
qcMUoAq+JvR0ItJclhxxskDpbSK0Guf1mAkSe5qNh4AcSmd9wbuS4H72tIkrfIeikCfO2SXV+4Xv
jP3oRZa7cAAw6XyQVWuOGPC3sd2xATVZ4C+lwvMDXaEVhn5HiiRVPRyESMAWs7oh5GNaaTvxlu7Z
7VGKxgcoTQHX0eR9CRHDPch+35hp6io9QCXQklQaeU5k4Zq8cO2Tufy8kQOGPBycSWAtfV5A0717
Xg4AT8XizMJy2K114F7/TCTdgXgKd1bACoUzl3672IwSVcQJi7B1sk2fVyc6ed0FOO27Im/KjvwN
+WIt0CUcG3iGKEuvhAYV+Xf+y47mIvkgf9qKeDVfsLSttnh7YRTsMaCU+Eauiloz39GV9iPqVL5y
synxtVhiG7tcf4hzVjQTPEEDdb0Z2kCvKkJsrYwhQrcTuDf5mBJ5WIPC3YTz6C5mYBU+gQMtGFc5
hO9kC4VyNoVNDT8o9+fonpYWgBke/kx3gKsTOhiCzAUzYSz4Gp+s5BOBNpYNOWGGV4K7A8GWhScN
TxjOC01fio02/SZINfJKXSOkHqu25896WDXtKPj/MqmPxzeNsA6n9Ihf4AmI3b4augali5nck6EY
NpTF0VIbIMuBfNG6y00UT1tRfE3je2tA94JL5wSONVbXLzT3/7bkePMncxYwrp2mnMrVn9yiwVdg
7HaZZN3Fe6kwfv221BGvcGIKlKdHhX8Ck0sfI0cqBzGRO8BcIfMow5VDAbCaqCme1kjaSvM1YIcR
+4u/Ezw4bd6ryySy9tIccS4DPT/Tp8Z0NqWdzs9qWjGKKB1PYdCWB1v2nfE1zvUcOmtOpdW3tz0q
gl1nQd2YvhRIRZt37jRGtoEoDX8/wwJz78/8fuzAKoGrS1yCJ4xdObFTnrWd8yAzo6UNGAZdnsB6
V4J3fal4FsN8Bq9wLfS0TLQ36tsxvELuYaMZF3dAzx9eijKvXH9eP9s7S7pBHohheRw5zaVvH4k2
5oXNZ0TAb8VkBxnw6N5iux0B6y1Ek6uk5hqx4SIv5A4mjzRc5KXeAdqdAyRKnP0kLCPN+j9Sq7C4
g+IpxOeoHRdF5MaiDrem1Vy0SOFIMUimYBm8mEI2V8Cw+9XZ0ByFG3kt2X/pXpQ7JDn1D7xx3XTN
LRkabjDeMe7Wp4UQ7jSXcRPYTDMCfArJosp80I+GmMJTgc4lXY/i3BLePIcFJ3H4YcAY7NrFQhkn
uFOap6V513v4ior3Weo1weBYbAdKoCIP4Gm3CE4n43pbPXmAOHA0SlojYHJIeVdGqlO8L2JGgCzt
XQvbzNNkT6CuhbwQ7AqTkEcOwaEIrVn5wEvloQkAThyKibvfM5CUZ/Q9fmEuOzpfofLNXxxqMWa2
EP06xOvZRE0Y/kqS7rYdQ+AJpKaGmEkcUt7lRpZ8TOidRdHdsMnXNxvLG24YCqfEYtDIWpLcFIln
5+MMewlLoMTBwkWkd87S+NyOVeT3Jpx1xYn5QpqOgIsN4S3pcLZUR4LSyvIIe8zZO0xeSZBan6BW
RPqioIPIy+LmsNkqHvH7OEzyJhBnTG2trRayEWiNmgdSkU84HWj2qgWJyCTspOup5s1CviZnsVzW
3FXVjZOIySMlBxJCqxpHSmM8Nc4/EKussIcPLn3g11LS1Y2o7CYvbuWDu1+C6IQKCMhLMwdu8QfR
gcKEhyMAl7ZOJ2fnv6Fp5BUyb5M1j1onff/QBx3AH3iMXiS3UKAVTojbS+iH8S49Xl4PKK/AiftS
y7zN+yH3dTKcKveLRygJtwWf1ZxNwZnHM23tF4+Q/L9c68WtMEycVJ1YQo6woFw7264ujt1A6jpD
yVg5KapITZDbtbg0fX4qmz/yoSfcBJL5TobPkTu74BJ32Fnu07a6d4gXJ3AKzVShTNvsuN5FmhRN
Uggwl9GS2wWWkOqvXQUu/7lY6nDfQoEZeqY5ysqiZQPdk2nxB/BGYgPzwTWV59V0I9cqdgCXj7iO
4XiE9uFCZJjd2bxxExGkjKgXoll0siB1kQzcI6rPN548hQiXP3T/iSNvXZzPDPuiItd3EQxs6F00
AXvuLtWO+nP8OWbFHsZ9lfqYRmyjCYeqyimIw91frSe7AqpkACBuqq3+ibjxRXKjHAc0f78nJaAL
Bm9P8cwdGky1iTQY9wfoyOE+synCdlWPopASYrdXNcWlv4dN3p/Sv/B94iX71kEHzmCIu4DCuB4G
44RQh3ExB7sbo5leVGwZcd4Fj+TmDhUBqjou1CxAKAPoHjLTXX2TwvNdsNhriBOSnC5lHy1QZrxA
tBPQ6au7pZO2fkGC5ysvTd5zkOSeQ320D3pFsOPjrLsGYgbwGy5PxypQKBdCg3ukXuFPdjFmwBbl
w12MYSzQrSH1dWAn5xZiEKGXpKp7nq5iA/90LJh3RZXW9Yg3EmQuG3j/tQqI00SllEAydBgeqd8D
4AwxfF6S4/L6MBKiAtlls9kDNAUdIg3/1+/GrrQuZAP+fJMpvH7n6Akoq5zF8t+GxdkIHGwx5om5
1W3x/5MyCKRhNZ7hJlx6HLfdyGkwCUCBFY84CZz49XlWpv57u9n4cNb1Whc9GX8d5jZ1Kv8neJhp
eUh54P20//ER7JvjQk6P3xgusRFDw3u6rMWEOQnSaUqp8332dJfw/qx7g0/F7Ovaa+1Swr1+kVsl
ytnY+e7No2T10ZiIJ7Ixe3ZrRhEQfULWunCd7JNvZHqdG/3T9X1/850vBCLFahQHsZM4HIN2k/WE
7bQX4ds/eEvfr+WEZs6DV6U6zrV19Qs2wiz/bstdh/zQxd+81bMtUUxzAIJK8JcvvVz9vxt6qOrA
97KyvDg4V43NJ3tLpVM673jt2BcC8ODhVjGIz4Ln6LNgKbirr6Ygr+pBoKBOGZXiILJRBbr1v650
shAgbpXZW41jV7U6U7OiP8B8MgD6c2/Mdo18JTYk4kf+Ity4M2NmJwu4xmVUmus+GzVJWUmCshXM
D7w3vjsXQ2sfMAfBN4LvJxosg1Fgndpif9/30YTNnoUupRodhplFmMvoI32BimmF21zSCpLsOcEu
2R1tQEslKOzCBpFBGZyFAkdF7AJfJJZSXRO0dnrTQyE0ZMB4xRlEbHy7xkKoTkIfbbhiSs+/67mu
cKEqjIRWe9BjJO2xNqBcc2UtE6J8eY5GYvgkDUJlTc8aMtGN/yHF6kL+KhoiAwRG2VpvtP/MaCM3
TvU34TZPwABG5Kf/ae88jgHcth42Z0I1XEUnlNL2S1pl75P8gac97aNf/3oNJgtxP05QhG9Wy4eG
+Y1h/Sa5UJT9likujzsXv33YDLqH1EUw2PMIyxgaiuHM7sKf7QfjyzYYWq9X5lNFs2KhWcl0KtlH
2hB03+jatcMn5eQqub1WW7i7dtX6Iyogu1jWtsQxoQJVUQ68zi0LJ5K3haPdGv6xsPzGOcl55N0n
nRjNke4qBfWSNKxQ1RFJocWVPNDTZLS00CDnI2CBaz5foxD3MEdkxepHOY6VU6DPV0RRA/OQWEDm
ycRM53YoJUyzxSN9PjixnJzWtK+ZjgXltAR1QrYzRZxTDnGQn/MG9ycllozyUwZFKZrahAPhvkLV
9ulNaWvNk+rvRqyCBTCZcwwlH9gExZ82rbQ++CvVG1EXyxv9nPk4WeCoDi/MTa6CVJ8CmS6p5gCR
rxa8uKjx3qi4eSDHVfhVsNfXQEXNWhcTnBEqeu572CR4rBo83Pn5watJ0u+WiQlB/IrSQe1/inqs
tJKKei0aPUjavf4RYT2K4u98ImnZ91ZR8kH7qClOrxc418GBi2/uk/Oi1bcR+41QkrO/ltPh4MrH
sV7853YayYra0jUiL7WZ/rgFZEHP3W4RKQTKluwLAjJQQEI4DoBtSD0kBceGlx/NuQx/ZMrIbJoJ
3LvHG2JXFt2tJcK1qPRjAacCOGdcJ7rpXvRpd82Ayd4EojAlEDP5vv/yYa26F+TuNO7rmIGlEVx6
ViZxwyDB/GwbpjPZjJHu9qT+LaD8PBsvJeMYykGU3G/wzAEm9HnwDxC/YKfD9d8rO6xWhguJ3u5W
nZNv2bYV2etTCeQOPihCB2lVpbKCCRpGtbUv94iI4bnuAo1/f1r/Nv2ID9TOH7FqaeIheWFFuvBK
P+QE6S3b2no14lpTximH0LeTVeNkZoKwBSngphLVRkckaO4NHLuQrXxNkQSALWsEnO/s5JArhe4k
pbaF2jmLCsiOa5wj+IBesD/MP0mNOG2bCSYHDnTf3pigb6dumzV94dDoFi/8jEU5po/ba9HFp7aK
TmdPrN6d/gFtlTOG0knaRaXBI5GPhZQw0CxahDFQMlCeNIO7sv1MBmkkWQtWwBT8B4cVDoSqX2Jm
LRyN2DHzMxdLruifaRDTwAQays/9HsgFExKySshqb8Nq8ubieTNYPqFwDajpvlVNJxH8cfu3wedT
Hbbd8aXuAlCzV2362oAIvMGobQVpBcdNU6gfZVzN65r4Rq7QEg1zSKatlR5bFtTICkU8Q150qAVO
0GprXcCp9DrBlMOEj2k12ikH+mdDmDuUcTiz5Hv/yEHGyTm0ZS11+TOVbkFFQ4rjHembBP0JIsCQ
kV+qe8Lzm7sGk9BfTLIutbdJABEvXAGXJjOUrLu3alcrdosNTbbsGuzXGgpjxjEcCqnvrynpIFoe
okclhNL44W4s4E1Gc/9SEL8VIJbHSvLe9ehuv4a1Gdm/ybaf7Xs4FikQ3zTShiJbF8zeOzWowLN3
ZMJ6VbIc8CT+bfVfFwm0Elqnn3DAciz4QTNF8QI2wmjnkNaJMdM6p2wjUo+xnyog9aPRbG4axval
msWZLWBIJV1OjCY1ZEOgW3k7cnsQbFgHKE06tZpvNocxL3ket414drRL2Sqhc+hG2dl79Gnoy0Pk
ZhxCETkil5ZCPvcI5htkoHJFuC4ya6mlLuGS7SPzb89pvCxqt6GlqqHaNf9xRcTEcuWi7636tGd6
ZAL6PFGZ+5rfGrMSU1b2ltrXD7GlrkpjgGtjPADgS4SwYkbFeOfC/gweef+tkoBCLynqawOUQQAz
MUjzcqCBrdcsnmS5SBMsKt0uthMmdCeb0dxxQoxEHBDoTu8iaXmVtUPp5Nxaw2FNjCbGwHJ9BVbL
J4vLbr4k1nHsQa9/ebC2JuuHCXR3GV3UAM/pQ4NQ/cqzFPH5dTWFAAMZiRi8Md1Iu5cs4RtVOXpY
H48kmKaUl6QTdDXNhKZcKD8Ke8Y4ULGJ4Q7CWl/Jul9ajPOSJM+UeF/f1KtnqdOIw9qRhpacEqgE
qb22OaRmYJPQAiERN8GshSigJL7UWTIrCY7KGyupfKOSqz/E5N2GJnDehYoa8B5RlS1DMjdBZ7Cz
Yq3WIxAgtwwuJ2PcC+1bCuoE0Fkkr6q3KqUgmKpFnxwQO1Uax1LnOo560CwbcI03bWd8gN3onGrU
6DDxTREXX3iirrCrfwkcCITp7TNpFFbz0libAJ6bKizl8LFWPQ5MobhQg5y7tcYiAQ3Rs39jRb6L
pUYCXzrs3JTvHz6CNtVdMQ8dhTX/QqsqLhg9AyGei16OO+au7YEqzGkOlrR7hX8uUaRlcXraw0oY
HFIerWXzSs7H1OOUkTw7YUHlEKoevBN7tK8vRjJdm2XGlpzDto3uX43hSu2KTOLrrzs9f1pSd487
m/Ky4tB2PbgC44eqXLXFWoXCGO5rDHZxZ3w2tOVMWfYl5BH9om5U0cCNZtPelXYGqNFn7qHYPlmR
ceCOYaXMI3kAfY8vz6BhR11c2Ql1hFXmb+x7BrLydl+I4xjlPyeFdjONLS9OpcAS63NrYbBXh5eR
v/gtsiQtZzbvPUymTBN/bYBfr2gn0Xo5DRU6Lny6UoCiDy59QpQSlj3m3ShmQjNPglglOkK5xzx9
XpMMuQcYhkyepaQX3alrjYBbEfAoENw/igbixiJFm0RlMoW12gk15JQNUvrgVnBmz0nM672VCU5v
WzWgyjhdJaQ98Iw9xD/2p+oEMUx6Es2C59/5NSH2xATtmPTllbE/JO61DpzPLGvUczvI2ON301UG
O36yUevJzboCmNkYysu7BYuOjVXsVgiIECij/CC/VjoDs+R3VXCyWs3wSb1iZdIKa9tySnPyqohv
J+y1lQTo8joyQ28TkbH70W/QLszhwWMPNhDM3HoaIFG8The74u3EHb3JxUG8C2pSb7THd5AfM86a
DS7KbInDGHLT7XnSeXqbZsKIab7qseLjKtlVbAm1q/59tN5bDjwl/2UejTDeXS1IMXlGMWaty8F/
rI6Z1F+5h4IddRuGhXBXqdoK2pwIImZafmI9QA7HWWAv/V9WoDdf/lMUikc7PZzcprXbpfPQvV9n
Cm3MJYTsym1UVEkdO7PBu+5hgFO8qha1NIZ+KZJl1WBcx9xrHBw2Q2PTJ4Qwtj33vxbHDVkfH17O
XBJGbi13tOK7sLf91RZdo9ITquQe+BM+2CGsJwZFHZPxsow1sRQ7wGvvZWFY2ddrdV8mUVphfj/R
gQ1m4rxebxgZQnN+d5EeLawTgZvABOFegIIihkHBGVyBSqzenzGFQ/aE41LuD0LukmGDgkbxNDVp
m7HYLfY1VdatIwBtvvHr/y/Ql5Yum6CtsgH97eVQQ6aegBS2Wrv0JdZ7NwfykDcJ4RhuFajGVqiD
5DKCt2/RNb/uvP265ZNEu6UXcwk+U8s+wrOJPl11HDuRRhP16/tkSU1D77A4JazYCu1u0VetrvcR
2OQf+DTSvMSkwneLN60rc6PUx4f/uSwGSDpYldMFYGfUr456Yu+TzeOlyMvLx5K6e3dAXRt1WNxi
Hh8ux7zorOT6NjVZk89OJ3uZFgPufTtglrozc43CP9bvYBJKkxDUjLVLv9lkxVgp6vpe1JTX5/ug
Vqkv7fv8ZpIgUqY3oboCnL32cM4oBnNZTHYYv4nbqPtwVCVlaeW1C/m2iPywrE1N0CzwcdYi6WVb
UjHpP6N7ZHJZNDsGHAhun5fqu9tZjx0mf8uu9picwOCXG2zzrA3zr+XFym+zXbfNlVUluwx+Fipa
4EQs2Gq0jB827tV9FxcrNVqcDe3qwu22GQb8saGc97xMHOWbAhuUS6A28k08nE59+mwyIyclKszE
56Pngs5bYtGP3eeFIE1KgzpYF/4XGAk0PhzYhv/pCH93mBhdjIfpD+Ewm11NKL5RVvRu9f+5LiME
K9wch+8JlCD2deMAciHR/BUf5mR9dQx9PIVVh3UrzQaoHo3LkvohRBBJkb/7zSWy6CGAkGwBgjtr
+Qt8mplX6llMLuAy95IggA7rxyVJdzVNj3H/ZEwxvP1XP4deunMqp2o9c1v6Vw5vevNb8HoVghWK
OImDfhP7O0tSMMaOERuHIT2T74TAj3btfWVHAulwyA5pjy/AkKbTKglDA2keuY5X7I5DLXpgzELw
U7w57IYet/lCbkJwtKk9smBdedAdCeV4M1JpK5F075MLPs596gCSQ8TdI3w/wHMgh3V5aVCf/oiq
186rPpVd7Y7AjCH6tDokSSlc0XnHxnnS18FswF8EYXpMt8lO8/xYnAVas7WuhePbarxCSG6Q1qOH
Cno9EmV00Da0TbemYHJuQqCR8giIL3KIbMPv+62PUM2l2e+F9w5yDEqRF653f3jTix24p3wSM1QW
S35MhOsu8iEz9S2tloUNKdjE9OvIrVox8dZfT+YE9hNPjU45q9K9Bm/94bDcpWwqXeZdgjQe+v1e
thv/QLBbYdHOgxn06+lve464dvB5NKCB3EC2Td3xw8gO5tddAt5fZ7JVO57jDMLyZfh42IUtm1/1
uoeTUw0KXfEVDciTyakep02VsTqLCwxYtchZVDsIFUK1sqCw96XsG3tn2Tb8DodZ9DEM8WqC3upT
liwg48N0kQ==
`pragma protect end_protected
