/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1264)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHIeWT/W5v/8QbpO2byUSiHrOk0XuMRlTFFsz6Hxpw3IdoAbrSFJ+Wp67s
4FYoNw39/09gD6KiLvCjuMPeia0wq0npIDhCmXIACmJ3dDPynxTwrPGFZgU5E3IFrofcgonZmqpu
IHv/nbqD3vtOPzghg96fdQyJTUzqiqYWE2eeYuQI/uc8ZCnEniB8kNh3H9qwvgCeZWa/t0r9Alrn
L9pQJTct2hJtEZzzvsKdqTOwLa0Uo7HGT66EZY8E9VeH3aatMpGBM2a1DRujG6NMGJrnLzpV3k2t
lsHsfyY82X5RspsE9kLkMBpMa5NNPve5ncl5QELUL1RtHkEC4ZErsImUDSKpNN0AKPwCEbQHLD6f
Rm+rSjq88xAdbm52o/aXrB2BDX2YUdG1ifSpHX1+MD3EbZDwFYf+wf7zNTwW/7TmXx5x8pekdoqV
IPTyURl65TcHp1EjGQ9V5WyCOtJ7t6v/CgvB47b9mE6GSSiXjMWysBrWDYDuWuMWNOrD0P70rDNB
d9QdrOEqn6StBRapsgq9GJiAnnO5vDAMGkhyvhDO9TgI6DLISWkWjGeTz4o6lj3llWJaLxvn3DM8
uTsmLSzabMtfQMMGcIw6S9lOBOcfvD/xhEuk5tgCQ/K4MthSbQWcMEjAkeyAguKSy1qO1rBcRACo
mZOVz1sHuDKW3jge+5IbrOtl5KxCrAn38Sbx9ZqD2wtBwq++A0IqC2c0yHDu9AQ0AtJ4X0q1SzuG
tc1Ih8aWWYUXsJxRXQa8G1mjA1aIwR4wZlar5AwsAwBKwWikYlgRREeHBl0R96UmhRSJqC+GIr2D
IL9t1Tz6vwlJrf1+9OYRMfSy2XjwT96AkaAyo52ovQERqOFVUypn5rUAdGk/msoFHOzjJuMaHx9/
dswJnNyUe8V8lx7x2PhmVsILYPGZw+ClMBiE4aVCS88tfQ3pJQ6Ml/yG49jqFCEKlUylMnpdxYjV
KvLDS1kHfWB1L0s61zuwb66AFkT2aRNqyY6Nksw8TeES2sLneFPbYXvXfMOh0LRM/YHOfW9VOxoa
ZPiM4Xif/h+LKlNTLZcLCVKXSK9oHVU3rFpQkgK+9RQuqbivHsCoi2EIh5LLZT3q8TyKibj/hQuG
6LLYFzbTftW/g+zubKSEAGtCPAPeHfnpQWE6CgGQuqVIbAPqdkzRV1XKVZt1Kez2u9QlMU1TjzKK
s/uskgBZzPZncjPesw3pRxXKC9R9f+VN8Wh4bQRs3Zln3GtPwubWLOzT973tkIC/LWMtFXC2HtRP
d1u5+81VTGlod/S2ZHtzHMkK3Gj56bYHHdkaLWrYfZrzSnAn4gSwuTrOSUpsPNZ8kEth3FJ0ymUD
LiqmVcEo68kgpnFJLEPPz7D0gd94ankMvsMDYnshwx3+FwnFBOL76L9tCMoHh93VsjnGyYKRb9gy
PVf/KkTDHMg+vewQcLs9kR+xr5+JGUkYWqSfLk+sqYJd57X2CUXV0Tp2iVMJEAlKmegrMe7KewDc
2y3JBZycCxnB9AamWjaghpgk8Nk9EhoMpwzg8LaXzD5s9hYXjXFekH4diEWkCKhVIqSDp3ONHmm/
82z+BjRhMzV4VvS/KldqIrRkvUvKPqjf5Fa5+eEhbhfvOPeRZOJSV4AYwSyCH4ZJA18s2Z10AIuF
EcI10NnNzHnPBQ==
`pragma protect end_protected

// 
