`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXWCY1Bx+m8ih111jhQHe+j2fAyaBsjyjcHKwYRLDGRI7bqy1n3yCrbO7
1zUje4pef19laXmBYISbYsfnsAmqCivO+zbCmVw9D1A76j/CaOJ1WHMJxXcGvYItozWvaD1WX55N
9NfuLklGYVvVdNI3R1kDwv+rKdRqJD41NyOwWNdtSUndAVH05v1Xk1eKHSABNIQsei5UkGe9oKbE
ffNamzafQbsgFLGCrMknRty7N+10QvI34v6Q3MSmQFgYXT/B5CD610okJ+BhblwYcvKJA8ASgI9w
u79w+wk6QXJkPlIQvOiz8zA3pDflvRwosASn9m0JmRW8p0FRm+vk700uTj3puLNJRLdolab00Phb
vHcp1U0tnfxvIplVkTg3iTW79bg8JQVQ/xlPMVrAKgyl+GuaecA2rJDZwoJJAsIamUnczC+LWPZm
vV1AxGkiMwQAJuoVy7P3x0qbnELghfpiS4ccfjkDiZqBJWxKh4ZI1a3pSB5+0tD3Wba4/Ml2jvuE
GolB/qVFuu8tty2HlgAZomK6oob8Kt6a7BQt3XcU8lYQjSa1rrv7YBl3em2JAaDTzbcWjmNM2/Lh
FLp40m6uYidLiqt+aYvhJ3utO3ADgPrdWt18kOTeWfzBx7Ihiid7mpyZQ/C8fnX9Dj0XnYHPJNQy
8bfGnpFO5uUQ7PUQ7u1g3/EhzJezHykuEiKeKCAnqW6/HsX0JTqX6yr+Mb6Nz5EOmphX862HLpJK
tfgOAmLEIKczifw5v7fqKMe29rGYJClTsJjKi0+JzLNNF61Ee/cpmLTnckjJLm/GJhnEEySb5724
XCmSymMTLlXyajuUkv+nefl4yXy9x2yAhXfBlAkKJiYo+BnqQEh1UNkLqYAA87d8AoAB9ihUb8s1
IgM+IoyPR9o3uY+NiwUbJmA8+WWguyhwiuI5cBoSnntNWESoTGk94tPn9TbimmCK7vJ2fB8ppcY0
dzN/XzQx6rnja2k1n9Vpi5cSISAq+208kK6KhLcxARN1Di+/5T8WUJbGsQIEAp1zBaKpFTX5V0rm
Ql2yMw9+OvgJAxGyvSLkasl2J41ecDsQfJu5XANyEZFSlHjJkZXjOHjgmmwKtfFMzI9zoswai+Ys
KR3wYYFcF3umYf1/CQnnBqdGfLLzijDrJzGGRJgGGaWe8g2EMoDSlbPP6/VtEIvk7f4hVT9aqbMv
X+Y+0mIISZckunInlgx7Y7MCXT/+bv1FTVOpRCxFuheLqFRrGkeqA87+Hv1L7Hkz/sCfuCPCa1dA
O5YApp9fAx2FBbiTy6hhMlhXzopsd6hc5uJZFpeW+/as9kegjY5O8sY4Pz7zlf3H8dkTrpv1cE2f
aQrW1aZlGicEdshgCtF5U2aWC7Kn6Ze/VdGsBfb5rsUTEPqTcAZMoNO/RxpYWLHZJELUgmtbdLi1
Kzp0bvlpdkIqyYhbAcfGrB3xe3O8CRJhVNsDS1sv36LhcMP8MMmoaYpddaeZ7yhryhf4Oag1D40j
RjuxUWLWaOnBw3EMkhU5We+z+1aJKld9td9kqZXtHOod4aESr1cqQ48zxCIXwxHwNV4RyT+ilsnt
E05Q5qYRK0y/i2lIJpkeKCpQnSDHk3EzQq5aAkdRlSJiUfeCkpxvnd6NwJe0FY9GZphDYCjvBP9v
sEF0ox+LJiqvG7U5W7MZ+abOIfehUGA45ALFxJRO9OQvRt2ZYL6srx7vIFDvmsGj9yYMNFR1FwwY
CIWFf0S1e2EdGt4eQYDm+CVtNDcjQT+gXDGVC7om3kd0s/SYRGZM2ctB0oH7qgGJuiE49rTAmMh+
BQIk5x6IhTnJlM7Rkn48A9uFJjflcvmDo86k4QPTjHl+p80OIZD4xXJFBe+UYHZ2V4RfNhpg9Nle
4wo46URzVw/WzSsKHqw0hLGiVCTvFOYhbNOsxAn8sff2XrVzPnnN2xPUAsXV5g6JTNv1lYldO7JW
7JfljX/lZDfW8vXg+CFNOakHHxAakLStufxjf6MbC7QkACOymnvRK07Yy3NRy1baA5MU1c8IGgn7
/Gc+Pk2x7+aykNrgnGzIw0ce/WiTWE6ww7UyT77pURbf+gS9QD77ALNU/50I40c3CF6J0WjOftyj
fEIf91j3yuq2baF8SH12rTLKBuDxdNcMXkjvJSY1PkCAggeYjjaCQ6Qnnh9qk5KUcW85dnZu+EKa
9IDb1T0q7Vxi98fa7v/AVC9xvNvF0cgXBTEDt5tVcs/LyluQ0UUd5VeOilAkccxwcHUd6zW+SZUn
5+hhhtVJBd47BgZ4jwY76ksxb6HhkzVkLpoJCfK9fSkvjUVszVJLKu3q3PlbtdTAuKQkw1IlIfUm
Ls5IJW9N7YlFfsc4tNtNJN740A8WTn2t1alBhCq0oBBdkdbrFvMjuVTGd6ErP5ZPr6XeREw1jaS5
6fUF4WbQUW2asDbn2EfiMWCnZp3Eo2pYz3PTG0liJ1347E/S4YDW2RWn5O13FJu6l7zJ7yjHfbXY
1cvr6yDiU23YGMykVQ9KAdE4VFpjzBm5mifqIJC66dXJOEncO3nG+9k4vgExD34xLEDN1q0BWhfj
eW78j4JWjeqEE84yQKgQLWIrZ7vje/IxplAWftXv0yc9xHFgWgNcD7JCJXYMo2NV5qTZDGqAmPkn
vU+GxHJJouEDDVC4xWcUchiHJMfRG5tJEXRqgHM1lFX/86CIv5v0GTARq/T+83B6PDTRgj3zfoT1
nHOQbFPSV6URdgob2OzR42GTkcfO43ufbrcU5v3gD2KMa0Vbf+jFTJqhPx7h6D1hb3WVkmtS4sr4
BOClKknWLlcI2Y76CKGrRmTmZ3Fl5rsveGAnYS2YMg8xwrXWot5L3csAOEMq4O8tl4lzlwfomZ37
7PhkYOo8wc///q1T8om02W8dUI/nh4zadm75am+ik8GLLOp5m+L4k/6lpJUefQ9ODpH0KbVkCn43
VxD1fqIYmWTv4yBkn55jwimXIs9Yr0Dsdrxz56yfaGQFVVNZPK13NrGXJ4SR4NaytOK5Ilo0LwwO
7F1wD6HuzaY6wymS/zTGT176cVHTH5QCoNjOzsiy/amLfcJNBrVCgREe9LKRdl7SueUJdGfQJ44F
81b4q51IlMxcpwcs2r776VYXSJUFyupD/GzNGKxtSPLJ4djzgkyhCRWG+mBkJYMJWoWRypXO/1bK
orlXPXvisfgls2LkAswXTYUAq5QgAUSwGG/NipusVSjjRNCB2BDU0LgeH8TfLxKnzPre9zxIa2kx
6Sl4OdXF/wJ9bp8UUKHzF9xDks5agIAuID1z1LPZca04E+OSjdrRqI5sdKbXwu4A+Pcvsq9+1hA5
GVEjzfnxChImJ3gGplsMwEm8H4MktDCiAww//cR+kOCIpFN3A3kI4HHss+DH3nIxILGbX/TY/WmM
f4FmE01TOYWQn+WcCaVG2ql8a/V9JLca2K+nCVGQzAiUOJmEAxf58IxRT665VsFrJ3K2UHyRL8Ma
xDbBMsGgJuzpHLfUKncf7O/AEs3PfYKTNR9S5IDvtT9gQLw7PYtIb/sM9kf9v2OhJndj77At60JU
JwRcjzO6wnU6oMLdGsLcmX+wbYz5kbO6gks4P4IBeENkDmMc6EVI+RXDwDrv8J1ZGGOfNHSsp9xU
3lXbFw5t72HlVTd13wMjz9CSzTPPKb89F/ojpi9G6dDnaCVAPrH/IS3KceKN39/feEJvGp90R8Fd
Sqduq/kmpGrc+VR4QktKfkVd8gNzv/PdVz+U5+CT9p7Bya9mZKJIsrNvj1GNQT7n7NDB7ZO103Kh
C7FN2L7C4WMTc1vbCloHFcSvFyhvBjeVvifYkTlp9OdRfWn0CBMzf11qCUdgngk1iBV8fyojCml6
wVtUPCvpQzXgHr2Y7pijF2FTqJV2BTjMawBnpJg+c0bsVlN9S7FE2KsvR3/nNAJdGZnLuZxIoJbt
XbH/qkeerc1358C3ysFspMMkgATqbMWR4RD/idJGCgiEIChplX7vlaZzOpTKJ2gRu5agmOo36lt1
MpqpA9/HBnu2cYoL93s+JNmdSuaaZAhOzvb12wx/iPD2nabeqP9SgNuEPajpR9FYZx4tqkJA4tXq
pUlvg4wMDhiVALrMHqc8xaA2neZnAryAZk78sQMqQOXPzMi4Oea83djUbh5FZL/VenXZXKF5my9C
7acgtQ8kTqTeIPYNDRyHpDAPBFUOEeAp1GblZjxgKpsGvX49S1asR1j47PQvNKl4kUuijzQxNsBm
gC2+6tgaXKD+mLbcrQvRlVOFcBJzO0SwvfyRa9TZYrioO1fAj57GsIcxwdGcULMLEi7ZjrKdOP8w
2E+wepRCkaOkEA8tq9Yt6/I4NP6vu3VrXhb5Jn3g7IEozD/IPI4vbETMkB0oJhnoPzU9xt+M5N8N
Wu82sxZB70mRUQ3+W50Y47rvxjiDrwn6mCzijcUBiFRdSxf9QJ61jmUR/b6tc4E2zvpCXNnErJlN
+oZl1Sz9dwY8b6mXqRqeeU4YHGwGXXe84rYJmk1J/hd3iMVtJ8mZruoK0CfE0wsr3+W2yEA7gkOW
K+gD5CLICAsM5HfQUOX0ab+PCVL1wPfA09rqZQ6NT/tc+6kOugY8tew2aybdeLUgf8/PMkz7pVFu
87KvJX6zsWFqiJnWR1vQW1JY9tkE7jzSEkMutQ5gA/vnKwQ9y1EDgaW1vuD3AOnNk0kyVyK3WtvP
QA/e+4XiVDwadbhvL9wVw2+XrNP7iTSNCiT2TKTyXp1eQHbM9iy1o8HdnQl0UAsLFMcuV2GdsfKn
GsKVdIqW+UNnWKTMvm9bNq888Mc+yUPZXQw0fBPuhEBX6pNE0z6U7Ry2ejdWwC+trlFp55sw6PLb
fGsn0a6xJuO71JDTGJ8vi0NwLCkJPHUcgSdFD+TahmnxtSglguHX6HFj3PbDc0nevkKm4IGK2Nh4
5CUHtf8Q9iId0RU+ZRIGqOtAJVrBcaxYISfHzjlVEXCE4Om70uVpM8Ccg7/ywAFLJv6IynU0o9v/
S2LxO4CcO4jgOjoPc39j+NKW32paqNDHYGVGL9Du9iVR5To4n6idKFwjfeXdYt7O0DIOOv6dC60H
x12ysfy3kTYl1hHW64oT0xePnBvNkiI30YI3KoYuMmGA5pjS/PmKNaCbx0P2afF51+e1e7E+2Cc2
0N5fdckvUokdv2izvO7c1wdrSLWyGZHIJEDG+NeZSUDBo2F20rSvwW7m89UpFl3LiHiYuGkPVfft
hH3wIPv2AmQFZOeao2UyQT4raoGntcKhM4ty8DPB+lwFS4nQO3qeRrmQB414xQ/J2ZBKigj2CuYu
c9zAwbYsDQA/jbI3QL1rEcBhtToCOkXdR3VdEwkLq+LGGh37hTxXAnv420gs3jY5UKvhYsUB03oq
E1NzZD6s7lOJYLLp2CuiMN7maiaJXCW7c7PVy6JxuZCIzKs5+KbGxy3IxZ/jHBqO+nA/w4Is7TTT
7f1cuIVJM/eUKE/WVbbgR1spN8GaH6zbjgHkmN3Py6WDQS2Ctmf+KPd5JaypaHuIdQSH/l1ipFG9
oafhUM8QjjVLiK0iMgGIARpUjAsAwgD11k5M+o845xlvNq/LgborzPd7XR9CQuN1tvNs8n3+GOTE
D62tWu2Xucv+H5azCCC59D6HHpmVLS/tlkPbR3eNGdG8DEiVgwtaSC1SPlT8hEoNV3ifQ8kNxBnP
J0ZpmhOtGFeaZnA5V39qxcX7N6PJO0lqJkl1Gd0JOtPevLqO2OPajcVF2lgMEQK3MCSVe+mnSJ3N
QQc9qNjQN0E8Hh7SDFNQ3a7sJFPeOOk4hwUWE6Bs1Uc1niMTeGpjDVs0cE/F6GzVFdM4fJzRhw9c
8de9WKr9j9TLcUvqqmDcn5SUQJZwvoiQ5PDOi6OFdziB/yp3qrzsSGM89q+w6gV2RKVMu1EDy2qN
0pnjv/ZF9eC+Y90HeCfNvQVunRJEK8bXUDhEfSIyKce1T8k6b060Y2qlC6lkYudCgztKlasATJKm
SDFi8NsttYDQr8H+/UnFRCU4KlsX9HQPfq0VShdCyq7WIHe0TTNLFB9Or66oFc1OLgQcYar9+pcR
PJB0vPU266z4/w9kRqjaXt+uwPnyfuSuG2GMUXjiGkMPvN/o331ZzN4tNFMPr+ZFYEaQMWEb7X3g
CzOY7MqxgA7rBVFfkjpkFqPB/YnDteQRlsffb3k+ODsdm9V06g+ZOfkW7HNhTPOQF8O5MFCe1j7g
qs8TAU43cEswOtj78UQnVBr4upu+PCwfm+XWPVehoipaOZ7Ur3RWtWiya4dK7LBnvGbLh6WVioDI
+O0Dr1FqCBalFrJVaS3pUS69SKZFdFg9InXPsLqFrxPEu3mpiY9/yjh4kpu6zPZ0LpdcsFRNE2CK
5ChPu6L1zR3pobWv0LQBTkCftHouLRQtKNIo+SMSetc6cNiGoYJgv32Nl7WjfDyzoMPohHIW4/FU
bvxPXBS3emoQl/5foYF6M0xCzxSxyOr76WkGhCpEwP6CV4Pc3WwQIpYZKISpz6QlgYCZHanA75aA
SKStprMYumKQCugDsd0/TAt4Z9RYhnj1fSKibL0mGNEp8ILzcAiqohjn8FYbaNbF55B8DgzB8gyl
kMqrti03Si4/0apR4v6yFhrPl8a1IImucOLxrs7icJSrHd8sojo83G3bP3EV4/gG0PaQ3HsSP6bh
zhufBsrfoyXVJYFaSUU4UYklSiGgO02jmJtV/ZGFdnKGnkt2iNIhry1/4uoisRfX8JwnT8j/y9+w
infyJSrQBgy78rOhHMAi6qzCAt++eFfq+Vwi3NOSF5f0/NzrkTeq/3UjSUh1IT8+B6V5RKdtDsuP
6kG8/jFUn68gSywobHZs96hhNHG9LkKTscodxTZamKNllhropTKzs3IvIv3SzGRnnBwByLRrwzXi
Q9nwB7ucFyP0dzPonGWfcNWV67xzNqyw1ZdCZ2q8NLJvLHI7+X83Ds7MpQtz4Eu3hv04HPZefKNO
Y8jeZVGcqq/DjQ8VuV6wCOogIZvKfJGIlryoi1WYrKClrGqFiAIyi3sHgu+skaGER3MiGv9PaJBZ
zan4XApom02G+uw5/WkRO53UrTEbzsJ6rEJI3w3+rwZmHvmfsHE9Xb18yiDTlS2/8eOfA+sdBwr2
Ryk+WLyto888E4Gd8+7RYNkqkow9D1KzwR6htWZzCvw+yVRfVKCwhikLZIcFCGaEt284L7Qhw7c+
TGpcw1PjrQvbArV5xFN9yBgDMoKPqtmX/ksqMvTR3SeIfYjTIDWK5+mpkq7Uf1SKP/QtoMV0mawZ
bTVK2EF+svwc4hZqvvTVZRptetJHsq1BPdPMW6C+A7T520Oq7nLjhq2zITeoyHdetQHvHuE+w889
mcC87+LiFrCGsf3od8lSMu2Z/NKH35Lxlpo7c2iOsaWNDWZoTHqNVFg1Yg2B4T7+dP4euaQ1068c
MBwBMguaWxSXV/rfhjGd+xtjzbOuQ3Q7pESFrSfqFpHLcTPmVEHjUcpqjd5gYFtPSTB5RLsghO3l
Yuo6S6NNqDgKKbk+6gTG8ayfl46Fp3M7zDC059t+fGcPWRF4x2oXhj63mD2BAKtj0zN45SWCNu6p
h3DYxAaPFe7Xp9pOlpGNT/ytvX3Md6k9GV5C8maOCRO2+nEU6MsyOZa8FsbzLjKoX2JGsKEKW1Hr
vFSVY5Mjt7V8p6e0p+Ph6B2VcH9oRgKm26e1jWKjDNLpV2g3Aa1A3TNAdhIEVBTCQwVUafh3kbmF
0KlLnlpqnyq/u+T+Gxm8HkCnYHjW1SwrOir4UNg0ZtSic8XtCudeZIozrxxYM4xiHlglqR+xQjio
idaw9+A6Nii/jb53KiVRnK7xuXngACX/GEbw+C/MmKxvKjGHmIID8sWMQ3M43sEI7pZNRVBdWlk/
/JxTQHy15yswWk7GWe5if5wGBKX43cX7YXrRHJE4eFq5GIkUGEejyzcgjTNPDTo81T47wH0YMIOz
bbPVQ29tPLALfQ9juFz4O8sIJJ+jLPXGoq5OZY3vfvJTxi4zf+MqZ79e9k7gdiWWQNuzOKqeOZPv
2kj3l6MxT+ZEeDqCaJDpPyiA+RjE5eIDgav0VgDBsT9MsSdsMtqDtg5XCSfKFg03ytOkUJzEmAEB
LY7FFkhBMc/FVJ3+7liwLSyjBKirUrQwHdv46g0OU7kNwB6WkRikbldP4/oplb7jUNfL6av98tg2
0qT2DlQXRy1/PPeSnaIfO1cUo7FSeHuSneObtlXHMC61F7GSSe6+POD64M9WKYCE/LQvC0gHZbwq
91omCjZB84wsUalfAsgWMHeEWVUhnAf9KuS/2UR0qG2OuSsW4oN9j+8SoCJatmyFiRmg7x3ZCqUd
4YY9JbyPIwgDlnMvcgiSuMkrnl885oBT+spL/E1xvZWHEnkmqg4csPFC9/VCIhbdRylsXR7mx9vF
MFkJVq8pWTFIc/V5gqUc9M6MGwUaLLaF2oZCu22QmL3MyjSBgb7y5OorFbW9wAD58zRugExTy40c
wa+5sIkmvaLwNLgJtETYtPRt8cWpZ6vFfQC/xkHw2dHRKV96kKD3b2K2Qghjk3zRSvsDmaOEtsSI
wUn6HNvxjJ5v/R+ICcxcWHWYJYaBkpzjmRrBOep+Fglom4PXS/MZn4iXCs9r8eN7Nst2gawHFcFI
PHHa+jL3tROMpJU4ia6m99KZkuOGehRryf/3n5075hQPfrZ8pYJHFrugLxRzxk8CRcsfWbne+wiZ
QE9cnNsebxWID4tcJKP7aTuST+vRx8NORnv1WoP9mUeKTXXlANq6EszkZWtVQ8XaJzkvj0A78mtU
u3gv7ElzqpcmMtnrjMZ2XE2fyIAP1HMsFNdAF7JEutw8F1Gws6lgzHnEDOHprXrIvNoDvYH04wIK
Eykc+uOKIkf15lJiDMVTsDP0+TsBcmnBp7Um42V4wN5+JVYiK6BglcAhyg+6g3JpP6uXctTrovdx
sWOxb0vpkrCWrd5MgVz+17YmNJfjLqeRyTiBd4/Zot4XN0/gaTccqA2iciGYRnJWGFJmEy9gH273
Xjq8ubG+s/RvqdDce99JnXnJQ5BIsXd+fsG5lQVaua/DGr0Myf/TICVKv2AIOC4WZakIXutKfs40
Ddnk/o8bKwTl7pUK+nlgRmTVYwC++l4iQ4mmPYblJ2gmI5VPkJvcnrbI6kwZUwrg+5PXCLIHo8GQ
yfVJC/jlz+y6RVjd49IVzXztJCgSrMjB+K9EYGSCmUP8jg5GniHIo8VYTTAxIZm8hbPBdpCzZf7S
A1Q5WAkYgbbXuVA15rfW3XMXXeRLm8e57RdFl5nAwdqllJHfwmkGokp+fdHj6vCAH5qzECNbiOWP
5tKrGBYu+ptxiSUa9Tg4z3W2r1Ibn8M7kfTFzjLG2pAkygJ4bg7/muC3dirm8lS2XR+9VLZH50GO
Fli0Wt5Db3cFfX8SibrOB4V78EPldOCaeTNf3HcIA89aVad5cNb2BZ1xxHEUG7e80Tacub9vJCzs
9NYhLW/yXTW/k052s9CByB6wP6JpnDfzd4RCRFzk7PgrtuObuUNVTuunk4bfU2/QwCkFpPrE19wr
J3sxqzA8XLqQhSZ7q77nCsWHLPSwhporZgw6JMBXf9dKbGGH2QCllm4RfXRtcS9x/WiFY9YUxl1X
fOmYeMDboIiAGfzFCBQiQ9w8l3vF9ylEFgZIsqqvmUv/1XpQElcekO32lUDCtCJUzWryT3yTDnjp
MTpuUEHp39XvhdSRBYCWUmH555MqCcW56sLu7XqJRQeuz4NYZhT94Ro1Cz1WZd9PET26mz9u0WKw
GkkrEGdlwT1t42uyc53z910+rlHM7nC5KA71crteRKfkUdoyOs4djMHQ2lzgHK8oEDVcbAsjZixx
oJY9QhPA/Z2L9eIon6+MTo8DFgbdVukLrsNtn49YwZoZXMVAWtVQCHpIGfKYxIcYOPawCF5flqZI
dfrHd5ZQgIocOirBtHmHBIS7wUdv9rt7N2KlL+ihg8a7J2ToA+yP0tdAokqfkk17H2gpjI4OJpV6
lS9WrdWFSmjblJbFwkn/S5bQLtzWfnD59Vhaa+lM4KsoG5nabc36ZOmqrMazEyY8BskY1czFP/ky
4gIyh+G1esJHM3qom6RYF0VNPhkVTXBuFV34C6DMhvN8SkYM2KAf+9mWTbYPuK6WC72Etm/iTwTt
Lria60o17pbHk/Nr7jIxFDygLLgNQ1imZQ2twthGM1Z0S/uMMfdIX3uGEufbY9ZCwm097gE/mkBI
lzH2z0Av9Ty0PaUsX/xahA0ELYtc4M/UrDcOBYoam6jx7eMKDi0P0krmTNgMgoyzDs026SKf9vg7
Vbbee7m68q36ZYiMzOS7TOq1FMDF7GpshpM95JseftTyfzJ/Dn/J10HeClg8Jf6tmPS1q2yhX9WF
yt3YKoj0ngHWPEB5D7/M+eo4UTpmXV66E7wlBx5aBRoU7l+6N4jvBm9Ly5VhvjJI+p38iiJFqR8t
XkDVhxLT0Pw1082r1bEpkytNBGGxDNkFBvFpfHZfQskpGWbPzSiABt0F9ML3G4oFb487E45PsrOW
QRhRCw9xoFV6otsoXgQSxqFKGzQNn7CcjmYjQh6DUMdemowhuydMzMkM0DYpr/ej29ee56UVQ/vC
R+PUuwcuabxaGGYQNyk24XGiEq3odHXvT1EBYLhuxvWFU93U9U1BplSYc2zSVTPAix2MnqEX2Ylu
zKzqoH8/qkJIYbAzgcrszP3SdKTwYG4/W2IDZSRFwtifioywdYFBXR7UzcrQMHEKpicWvUdRAWzL
ehjyj4BpIBMVKREjKpubgFtJ5cS4tHeKPfLYWG2Y3Z0E6pXGaYcTuq38zWdhNsj042EP6G+stdkb
YZMeMcvFlUHCtVmqV2Om1eJuZgT/KtUytHaBoawkIKVlj2fkpfMnRSnBnlJE6UhSRIeqVI499Lh1
zXncFKypMLRl9giQN8jQ7jzcibht15jmubKPXpetMJ4EmVWgQwkk9ljlMbbHPVblxHQHwRhuSfa+
5Jha2OWFpRhgGyvIRzA3zULip3rLPQdn8010eW4msHSdCyVtFuCd7pMQuVTmcUOII9jkdvmZd4vc
S+7tB3bZk+nh9imSw1otTaqBPMfdqVRlf39BcEpmBn+KqS6bxxVlAG6oqmzJGL1vWPJGqt5M84Wb
Mcs5JWmtafU3tvBpdGH5/UBpEkmWH/6NEwVwbU80ibICPf9AY0ZU3oEcRa1jjVZWNhqkFG49H38X
Z5fdgZvkvmS6RS85iUU0ihtgRtYZqz2Fxn8C3785NjXqInhOVpuac/vliU90urt6OXeNNetIZMLB
PfTpXyr7WpaNToAfdvzJONQYpknPoJPGutX6HcIP8xoOqzo9/0kqGt0Urjeo5k/mWAYDSHzflFsD
YGMGejbSjgE39SnLfde7o6T8G8NMr2UOJyjoO2y3KqgNfJOWBnbJhsIYhxyL/0q2iiSujh/5lb2u
xgre6n5NVnRaPxJ7qkwCdQhJ3zLyQLEPXfiqfwVZa6gA/9kLFExB4bQ1dk9Qpev1qcKAbxuKMDft
lF3xN9R9CqJ9PFJ+ZbI2zLLzfl4yCXlkFu5LvL2tur5y8APL2JJAhWyEyOK91jpkeaxMHQNQEUAm
siOGvwKVGhNUltzMguKFs7x6WKoogI8KK/lmwOBG6rYE9VQpRtyDtZdMXA27bG4LjWOisyUlOe9H
ih2j2Bz0gw+jFIdtzr+jTvUAKNCcUoET+wV0ikCbBI1Xrit8rjnKibBEiBmOOqKNhEqn/1VittgH
1VlKNiTsdbs/UO3/KoS9MAFzXr/GLKml/VV8GklDnDpgEp959CE8qi1qQ6hUc4ksF/8bAWY7cFrg
rf+3IUqrj/5TMJjw0ivuD066BsNRJYLVkh2/I4GP1sl2vhQHcGu8l4oGP2u5CRurx5+Yp9PUUlCK
Sm4Z9kdxcngyJWUZmTWOlQDc2v2P37VR8CSoEvGISXvjmOH1VmA1sbeMMBlX1/eU8rcbS2ehtjyj
vjIFZdX/yy4V2W+6AI4u9iR/cUEsTZPWppFXUs2VukCxy2a0FbJk0P4/yuAyAnO6cr8+dRC3yEXm
/5g2onMbPZCQu8SixoEkt965KVTvmyRFyvbHigGKA42DmmtyoWX1BZNT74+WQKgfmyk5wjxNIcf1
KnVooh9uNxt6Ja0UBIbdbhsYk/gK82ngwlO24l25C4MebWwJ/e34Ps93cYR6S33tPKrNEGKpPHW8
IjqZBY9A+P3Xc9iNConS0yCAaimDeQt8HDxtlvOgm2nyAmuLb+1aE9GImuaMGCvI94cnaPEv867/
uzzLSeVjYAvPY7PQl7AhCwEcYZN8B+0+mzKqwZPUeOp0RBJY/IuUKpqJVyg4tFpFtajnIF1kBiSN
50icfiiF6yo+N6H9zQ+FSCnmZR2+ztkqDXG6f/QK2vieFVWyPn3NhZSkfBYnO015PwZ1KhEuOgk0
TIylHvNZmJ4tNGaFcgWQdJm8us/l+moMznibnNJ3DvHc7NChWAELXnina69LBKdM8kqhKR3W8IMb
NqR5R6ZV16gX9qHnOCl2sM8vpl4YTZ0PvEn5Fu/ZwuY5Woa7Uh/dNPlyMX/BlUCm0bvyysV0Wm+E
Sk0UzMa/9wpu85DeotZwK1WTZbT+5bpm7ldKCiyw4wquvTVy+4d+g8KfUVqPLKL3hFfvvs/eeEaa
1QDE3qynxfS8RjGnTDZiayrQ+Hk5nr8jkoZx3RAZJFsQMXORd4xM6Ami/70q5jArzj2agbndn4dG
HY3HCCqoHY8x8KnfIRBNkuyQLkQYWAMtr43GyLkKG7r8RQjQPQi1J39QRZuek2GOq4A8nejEBIgx
bODG0JzDJVd3SfCwcXRGo9USyFxqR6IbKdf6+WddFERk8POTXnkePnYEA9dLHT0MSwTj9J8ythxu
YrJBvI7EDZAO6u3ENJDrz4t1jGNiHU+t5W/oTOY6xpDlsIPFU6JzO+SyM0zcsq6HY5jfV+2jEL0z
M3tUHlkyZJ2YBuMStb1gn3IIZMn/vlpQ5m3DRXTg18kH0TlqHaDuxQ5wVZIovQpLp7cvFiQzO3B/
StbRgc3uEbSWrup8DGl30g3PUfIM6VNMw+nK90GegkJ8UocQk+3cOEI+KhvydYA5I19rJ+qpMu4P
xp8stFautVRoe10nj3dg2Ew9kRikf0wcv/+gZNPD04ColQVtURzrff6D5OvwJ9CMRsTJLYD57go1
zhFMFpIXRf4YbtjJdARGO5AiymErIRRuJ3Of8EDkLB/DCN/uE1zhIokI1qfuyRMnuKm79NOevi/W
iyrvpL7/Jtw5TrXaCoOTiS20v0paUwF8dnICNNczZLPv4gfdipQ5+gtlBvOx9UdTR+jWHU46y8Ny
ABGyZwCtkjkuTT/kgl369S6rmp1i6mEdn6uD/y4io8Hrasek6cePjdwsjpdd2Nskt/elguHmQFIc
Splv0hZMcv2g4/iRHEi55VGlwzDBzPlJRMPQcXI5CALEmV4GZJnprAbt790g8+HpxD+B+1w55EK5
q2A2Uo8PVLOrbBaY9XaQH0nYCER+O8zzW1R3w1HRWk28mMVYYnL4SrhqQCYHnT3kEHc2GCj9N+qH
r2L8aAZlSOddwaTnpjPFvIlBzpgA3wG9lIHA3+fKUehvHzYbGPTh77lnmqW7e9uYTZjUCi2P7auk
hfNotNk7KPCMNwkS8Yw7gW76BWh4bzlSGTNx0lUSsUQF1UYpF0CxG6KjFaRNeJ+9PuRvyV7FDYEQ
fFk1yM687NgUFNByfMCQjvMrQH7mZsjJ3cwTS3X7sKcvmIXi0Wk2PgeNCvURJj6+X5a9w/GhlG4e
oesFF4mHoh9EN98lBfte6hIX1hbMN7bXaJO1x4bJdtSpL8dMOFkDkP+Pl+Ddd97fPZrYpl3stVYz
X3/HmkFYZS69p8f6+HDUEpRIBT8Iri2Nw2/+058Zz9Dz5VqZ5Mk7U+tVbuuA/iYqgi2SCjjTa0gB
sn6FkSPZtBHYiRRldM4ALb9JQnq8wg2n1jpB75ouV0vqyRKjODQJhEwQ5uc2G6RIKsTucN0IdRZC
SemKVxPBPX1x6/OwHAsUA8U/+H1WV5dwM5i3l2fhMNjREGPAxwG9EHIacGxNmSwOJAasEW7W/Jt9
0veMOa1pXPoAjoWF3WkA1oHy/Rjhyn4Al/eYsVr/Ymdos+yOuK6N9y9e2F6LMxxOJ1aFTsF97owi
YEDYFweYN7Ja1S+osrDc1phks5uO3A+thLTbhob52OBFPTpVRo8RMeDQSODfQiFXNfiXszhlcobD
LDDQhHwqzBec6ociO04HTwkteqTPbqCO7WT4PG/3s175Ff1tofSr730p5NVoKeGPGCBx+womenFo
oTLknrPKZK3WZDfYhAKp8JMYtXksIdGqd/JxrJx5t8q0hBC0yL7eCA04bOFyIfrLFxYzy4xXHFzb
GUU8OGNg5YqKgsFvhhj4f+KKQaaWM056uWyoxwsKEChrjAXEH2OzCbKU//9SH1S89mkOptVXmtqs
fr/hyLUKxH/T8frNMBz2zANjDE/6MXt+tUKT2n+kawctYnEI9CEGnIQCdSfYAhjK9uow5ZtLvMWb
ZWXiNpEiRhsST2HgoRe36STnWoSJyn3Q3tw4ofFDAYIzRWlqc+o7P8EhxZKzJw2ov/0qmgUf4nql
ggDyROP948j6I4ZGKz/kGV1r6lz0v3iciPVlvGFhlaUKzv+PL0NH872UOkbB7FlSDS1xOYhG/A8c
HuO/wgPDEEZUTgaGh72Pocx8mXIiu5ZlG2fvJszBrU28f/sDTPrfxsD2PV91B6Lj7TMqKWF7gvYj
bhou0mdQ/flnUTFEcFMjwubEBU+Qgib3MtnCPC+MXdn/mIylnE2XUET848UWvUw2OAwZi0Z/aFF6
tYJDhtulTlgLEcETJ60KFkq7bACbL1eo90GV6WXfHqycgJC/T1+shRWlvcMDHAWM79+Rdnn4FKmQ
UGPyEHDNs7QSblfMHtesF1caC3rr/x7YtVsjzyfKFMld/s1tsnLVdsWhnzo4FUGc097yjn2sA/7H
JA5ZbDUjt97qEuHvS0lUNN30S6U0RFibBZwMUg/IOLlytHOFC0PEjaO1Tm/LVYswVqaIHlAvRRmI
8q3N9TnLb3iF+oikLt1pqtVmjiydt4yjVjuAlmrc/gT0KwI6J4K8P2kgS84OUwF76eexvQjcuaiG
s8VMMspBijY7/tOGaTPe7EHPTACH5kqd9wnfFopiY3BFhE0UJIClZJMlZhRA1PU45Jr5j60G6ayv
+oo0/S2Apivlgtx3s6ZZj8HGnADTC6XWF494u39wNpOy4klZJh0CpxqQHnMMVcBl+crMWT+yrNp6
2BsES0hwWtGaxBLHeVTxjO6UCne8oHRfumZnDbuL4+CUaETAdQRhIoaoUFjw97yV6I/vmFfasZIi
M/CzZkIvpfKjb6h1Ef3rYzQ3JmjunZZbX4FyZcB/1ouUIO/QMTFsBM5/AtAeB6fExU0dgIVW9agr
ZzGOSu0fila1T3PDpXZwPjBTCAN0qqt46KtGjsHr4EfhDGl0l2lnAk8rC6jqK7B/o7lPH5b6i70A
QXPI6/XJuzAd7r3xnnotu3Lq8rbMa7ZS4HKa/6ExDYTejCvTtbj0399m4t6nkD5V7v0czOf5uAGV
vAelUHWEiOHlj6fLQnbmTWm0250HDNOvLXa1T9aCZvI1BMaiG2Ixp4ixaU1Oie48P3pXbTTJy9ip
LXjcMnvSFYyUzC4OY+ckrqc5KtEVyqBvdEPTPUjXx9ZWrEm65yo9i+XOBmFNHb2brhuISo4AECsd
Gl0gvGQoDQ6XtP8GDkOXCmhny044QPJnDXl3j+lr7lPotJRx2NqpGNj4Hp8ic0X1eLBRVOXT9DRY
iN0udIyry3VP4+iGskSPGcY+V5r4mIrpv3f94wy+2D5tEmMyupCfeNpJsbiB1bg3seX2U15VG/2Y
Dh1RXtIb5cPFhBnXHKAGdAyvjC4iNcJXGhdFKwM0u3hAWpAGk1YKhb7H41aMKuF1LZ6iY34mFbYt
aiJk6HGUUSo/h2lp/PJjhD6s9VSEyOZGucOBo/XeExZZZe2v61GIHLfD7ItedadxhD3owkRXnMZN
nSwrLetOYqTf1DRVrK+8y4tU/MDQsxkJyuNs2G1uY+i7GNanAFlfZyhBbw0S0OY1JWj29nielPX5
RDzf+cLLZDC5GwrcohBZ7E187F5cP2e6lg9pOAvuuLJFYC+5VWOQ73pptSw/l6izURb7KTxaJ9Q4
6eehhImBeO5NJtbrhs7bgPKHWF1b3lx5lj61imRnQZEVPfM6NtXjPxQBw1b+rr/GeKt5Dj5wYXKd
s5ZHHkftDTnYH0TcYbJe/R4CDAAsm1OMWPNQARqjkkOqVGTVVvfWaGCcfdRv7HBHGw59A5VLv9l8
uGmZkWF+Ys0aIGTEhX2aZuduRuw80aJlJKhpCS/hNzeLijLut0y4jJ0sY0XCPuB3zVQ/Fc/kEC7/
lMDvpUuwUAeSROJ9+NFdi5uABlwj8UiRmtR6rAsUb+bFyCvhY9/Jy1FuU2HXlCBtvXs+AySS60+p
GBxTgOceEIP+txznS3c2LYhBHnzq0GXTW8922CxmJMx94Ok5sKW6Ef7m6i/D+Wv2ovv0S/ZsmSPM
yiJxPkrQuhVAJtA0qZcXE5fqj4uiMHnPl9o93V+6T28SgiI23xsZvuZZ1m9uH7aGRptJrEknI9+W
ODRTUGf2XtrH0xXqPGma+svqj5Jt4//UkmyaFCbkQ/uyjaeXZ2bytSmBsyNiQ54fiZF8BSzSgmdh
r9kjaKamMkWraeF7+GfXp1JC+xq6F2PgCBxhBQhV/cuxu4NeGK4FF/POvZpW12w6Mei/sbfymVRd
lU3sJKcb8PcL8kD6SkfUeYEfYYTyPttQeSIrcmlR8JFGyilVF1+QM0Q4xIXW+9QUFrtZSmgszJ2r
n6wNcBcLbs4GYXwBWml3iZG+4tfxOWTHZJmNhDHtzgL3rgo26mKZMw8cXeevy1k+hyg8l0XspZW+
a/QXZ5JD/z9d8DALHJEZu47qnGqr7g+ootH306QDDJxtDp1lzaVEiSxK0qjKFEXS1CCM9HQqsnG/
O8wmVQ4KnsxreUHJLPN2eRHxUqkSs2cJl6IChQqxvGzxNUmBjNRbOxxgETyQB0/tPNIwxbCg0WG3
wpOwk2azh3IZOJHlSqqFErPDu3wVAFqYjsUAZ6JzWxrY/j04rsb5HqV4s27HK47j7xsX70ZfDs1t
RRhPuoQ8ngTxbOCtsfXT/fzklgBJJfYhYXGPYuLHvD7wGszh0Eizd/9efUtB8VlALC9eQ8n3Yq9b
2kXITBEBX7RbOdopk60itVVx99NDcbk+borJhwvEiRVqzFsLjgRBPvXgwaclRcJ3KIXTf1KPQ4w/
Uege1cvX9bigD++NVTUIPtRRNi5j8y6xPVL3bL/7NvV6Bs5qHORx/5JrjEOBeI4nIsnIy9ow5Wzl
YQnOXB1JCsuM49jS7sgP5U1XXz42Hpp8Qq3SvFgnWu9IfwnuvnAD1CGTJIzEKCcyHxNasUE4f9lr
H36rlRdM2YjndbY65XKIt2EDk4xg2+Cp9OWhnUUH6AvFIu7Zg2jCpFENtqft7xFtLBmN3SDympKJ
ZcH9MRZtRCzowLVbqAXyDHyZzEJ+S8QAB/sk9dlVXHqzgJO+aJUVcSDM5Hm+nZnfbcBJH8Lj4XvO
TKZns6tt+HTonTVNVAU0fm8eW60OxPRpizmSUcEEFv0a/oV+zeDjxSF+OEq/PsvBApPHPgN/IDpJ
sGcul2+52hkAwwQhPIRL94BXrmGU1WQM+BYBdLieVr3gl1u7M5AfP5PyB1giugie9JiAQL3NHGy2
0jukdCFBN9b1ZH8rDg9ZEu6af/gbnOiiRN8CNhpJ7llEWvCOazw72iYelj0HXvkjWSBXl/cF+w0y
6xH9FTqi2B/GOC+ryJ0NacyZseBrA+mDJRZ49Yx/SnruXL2KN3asTNTOPbNQDZEvMqE6hrstSFNU
hPeWvPMjqlRGW/rvLwX3yPFnYr/mgetbw7zCv4Zyz88fc2a2UO8mvbsBpG+QT2U4YVQ0JUMEQY/H
eXKPbB1E7xzoeZJxbUPPthvpnvIetYRCZT+/mTxMNTpxbIwWyM39d4kjObrnMBmtKtDaLdlh60AF
Y0GtaXfzKBb/ed9rxilw3ynV4uFdaMjPz/D5nVSUC9uZ171r61P1s7Mxr+z6OHSx0Cwm4TbxmsyL
8bskEzoSQaKLNC4LqDePJl66DwceeV1F9fr30+nY+Qd72GY8kmr6CUqwZyJjKPtNvF3/QWBiPDOF
9YvupdlQPKuWeYEzZhlYOS1x++o61skzwhk2crDITuc5clDc9MVoKLSmoq7O6WSH4E/DxJxUBxZh
AoqCRAKmewNL3ee/AtP9NN+xsywOWkwqVMB85ZJg/y8VLcp9mpGRrmDmcB3u0aoqGk/9ZU4FW0X0
OZzv4qMmH4AoE6QRfvBYHc8O+NF+1FWnO8qKqQ0fmgRmKHvd2oxdJ0S3HPZP73mzonslwkossAY5
Txc+CFvPy9G7k8q5xgkjBak25Pn7nUcOEIDjrqWJfnk/I0wVN5c3/zWk1PYD284tMRoyjgvRjItF
fQ6C4LMTmZNjaaYdcWTUpHMrbofbfacYGVJ/rWnwoH6qhwOfJSHZPS2pUKJCRlP0Ys+l5zsRP8nz
RyqeTHiwQidSLv0s4tNdt4suAb3zh37fY2Zg35GnI9DSNLbgkjmoObHPt5huHnIxUEtjj2Dmz0SD
mCWtIHl+ol5uoDkW1Bw2KkavS4BcvE2NnDGmPCgUwi9edig8k9oVcQ9218ndKHpOhmyMmM3fDpFO
3yF7ZmpTtQDxXm5CCRgjneLtHnKp1vQ3W/cnSc6fsF9VyLGB+x1JW+dEV7wdN3Tr1fldLSz/BVRU
pbFlO2DB7gOElHCtZxdpwVZBeDFUeOrR0uIKeq3lN9eoEjXx8uUdmckKkstdrvxZPuwJ5nQU1Iw6
S+mO6c8e7dRjBheEidvJTm5aBQckvS8iY0T6BQm+62o6g03nvNdhCIV6g5fKZJx4Fz7QUmcRSh+E
PCNZwQnPUDcBrvEtT2iB0gWbTOcCN0erjYettaTYS42Oiv55rlQNyRzRBfKeOBZTacIEwgkCiTC9
by1yKUVAWydSGZmAh6oFfUxuLZ2locfiiqCt5nm0I1AYCFAGu7G5wThyR/GRAkArr0dS4Uf12XpB
/9XSfV/ZzRn1ZxFJX2KdFKp2lo5kKBn8ie8DVCPaFV/yTWAi/bwp0Q/Rk9zOek6HzKKBV4agcbSF
a0iunDPPxluhQ8L0NXpC/Uio7nGh0j1zPo0G8w2kp9e14WiIeCjlRBNT5lFf0IR9TwYwNrVVCmXh
3ssnHW430rkFZJcwFIiErnA3zEICti251EQazCPSPDd8kORHYNCONx29UgGyNXzpJL/Wj6Rr4hO+
GYJpuMXFSbhMKRHKp+FEwh7/15jbMFU8tdSh8Y1kkOTGYhGpc4ibphwB1zM6v5sQ505pxQRN0V2u
hAJKMy5Hg35tj9lTm7hO0lHPriJODE8qt0r9/s20QrnDaqHnwrStdH90jTWvz/JmNn2oXH8HmTdP
w9sK0E4EN4FWWAsPmZys+6PBd5wxKFL5vYk0E2KSmD/6AXzQmxB91Qf8AHRE5NEv1W/H/uEiVZB+
kMFgJJpeJIm6hHlR8RQa3Gr846mh/53wSD0Z0h/dLL6SC4zE4tr0NsrB0ajefdEQ2hCCVYUw+nQf
7okyvERp2X/gCaWZMD5hKxjcTv6DAszLqgJGnMTRbxzqu1sGANI9acrAEeNRTZ6hP7BrzZ91LxwB
oxUPEQ2WGrYetW/Yl+81pcetLa6pHPzsfUzad6J87zGnoC/9tIJPX3nsdL4raJohNIm+TU+oGl1D
n1vmNZUOe2BZwrzmlyeN2AapI6A6DltJy51gAJfYrFSFGxxsnSkfAtNR6nBtq5LbvOE/G5PTM68W
DyF44vylHsOR2DOs34OmShLFIIFhuXYh1vZPJALRdMBo91AqaDgLsT5NbEuuhGv60tC+bE5awLhq
yg9rT1yztyjpWSj2oyThzZmpGqCgd5Sd/BKKnapEc/slAtepg5Q6lMT1yb5dM9NUZwZvnM73PyqA
2AVh4l015ZvbEiSizePAlVlL/fRAAt8MziPsRQqJC3mQ5SmaZBOyAmOjhcHV6XoX8AbSy1bPVZwt
SibgdQCIMRl/eoJYc+37JO7bKRdmZwWQ6LE8VpItgAdvbwxZIxxjYkajR0TVUy9/EE9EESKcAKxk
OPiK+M5MkMrIr7zb2atDlDCe84QNRrkIDaJDHBtkvhD4OeXbxKJS9ynAwiIdRjYWVkHkeLY/CYEn
1fgNe8Z/Cb8koI5xlhDw5aymlgo7JRgHlG7MH1ZD9O9vSayXQezC8RHo7255WXbJj98td+uVd1Dx
QshRoxM+jo5W9J/ekjfcPFC28tcnqCjzs9B44JgJdhn1tU6ihz/jou63dcE017PV6MSxzGf2oye1
UdWm6ry3gzAFJuJCeLwvj5R99DOYE78EfTwHtv8CStrMxh153IZM4A91MfpaSC9xRQsSwY0Io7nI
cSONbgyxCJBHU9dpETGVuMETvxW0VR2ePdfIclsqURr4J7vqvMQt752NXzAdETMPWzqyQNCASPS7
FLiKJsjsBc5Wv5gDgmqHikqltNUIDdq56uCqORUnDtx6Q9arT5Di+M6ifmNnVlzAm2e5Iwh2wFRV
MCsuOWkTVzkfjcmOXzRk+/PeA1kI9paq2aUzQXNsGbXcaB3m/EKEFep2SXPfwgTflmtznGndr3g1
5AeMbr0wA0Vi2UBOrxzHOmwA23tU+f3NjblmaBsCcizhK7o+4W4YJJHb8IbrbOSeVYS9IcY82n/Q
ALm4xSXD/Ii3oLErcLZ7vzAUIAne2jN3TulHF9bPHtin/FVzztiAae8JsJMylX6POVunbewuEje4
R2soQnYQh76VoSLPgmF/RnozyCDxtSfpU7neALkSVvDDTuPv5MDVorwS1eRVaZtOERBLEYbP0yxO
5+kvgHk7CgwfhkpOBdsFzdMm/m3HAlKLb+S9oL2LUNXoaRrjk0eCYHLPTvL1byRFUpV+DsB8/KVC
sS/G2a2GNG6bPscxewtM8y4EWpihRlTtMy0nHvmZnfb6ovYsFPy6OMndj3EuraYNk1WebYFLbhaR
ambD43IBWK1rIInEZO9Wd4d70Pw3yDnO6v3vPb6rVjL3Oa4mAafUswZPjrpSE2J7sOz3jUbtdMBY
E+z4LHcIwMfXRkkzINivlBx0aAjiXm2InkiiOriedC9Uc5289PNIXmdGdtCuqhulxVG5dyXI43hU
t/HwipfLOVZP80yfYT5RVAhdV0/5TjMWh22ESfzgAz9CVsJ9wHSmJ/jrEGOw9isPuuWbnvyqft27
14Lo8R1viInhEfmS+VsMWqF9h2D7PvGA+5deX3jpri5R4BRNzvBoEmupMoBZ0738t30dFBvfy3s5
Z6oFIdwZ8C3fstT2rbrWLc/AzZvnPdu7cq6IvqZwFsPTNQjq3a0goHM7vEwqhBtcyrkpzssrytHH
ELva5ZxPLJMkHeXzQVcRgmQzvraf0c4W8s5Ygt9k+Kv6EzwFdcKI7v3O8k88q5X2ofEXHLlF+oeK
Ovox2oM6jK3FXAG4W+39cx1X4Y11CDtH+qCy8jWlF/IMKQAuLZtgFpTGPi/+4HiL8UfwV2D8U4Zn
4ljLBH4k7OPzd+rKFNCuAQLHwQwBc746/5V3eB7B3NFhKu9yq4qOVQS/hiaBsViriXTmv4gIOO3A
wp6b3CZyW0g12oZRhA0fpYS4GvrfWBWFXP72E3SYzsMOcEyW25hELWhqkNhnwxDWNyd+ryIBToH/
gD3oGjIRfCflyWTKwLtmdVWn1S5dz1R2R0GRNDR936As4lUXBx8BsprGr9cbL3lYa/AiXT5l0/0j
hB1oB9HeGeUjDMBmuXiS67bLnxaoaVrbP677T3RKMWzm+zWOBx6BqPQwXhY2oZgz3jiR+HHCwRbe
zzU88hPgBiB2rGd5nqHqKZHnOO9wiRkFeUUIpZaYOHR7Olnf+AYymnDd869RPd27NrXgH33wi//N
qCHLTnPUPzaTFmW0Fy1y6nDvwpGW/EnTrHZSccXn6B0mhPeegQr8voff0tofHumssB9xDhNf0qg9
yBMoVZjpDxS+vT58RsKcR2jLQYNRMV625gPKRtQPDYnrWjrU4PvMgsS0d3pzreCTCrAB81yMuHFV
uqbooCav6BpBUhzE6qwVFtupNfcHmsLULr4rQY2gBthlcXsfGanyiSO5kDkVEApCf2igslHFzVQF
XKVEox2sfpCXI55qRn4SI4gRpO+QFKU6dyZ+YdyVgrxa60LTx9Cn+Cd9QRTFN20niA2WqE5Vy3xo
iu6ucDhMQZwAv90URfVmYQ+RYS06jt0HJm2CD+Ux4xY2tJSyUGjgDgcjfJYlgHtcpEJCap9lTf8n
vzRGR+RagtLoAjOskYt3Oi/av/3tW6HHaEvCf3gjaCh921pD5Tq6LnZJ7JU7GT1JedYIxRakU8Cx
I3hqQknWksccZ6KYeoomU7PasQu8w9l1yclX2isJxv+1hVCtKVAL6tZZimMnQved9DueEQOJAIgO
MNc4X4leJ/o1XFsP3Clku/0DMtHNLflSBLawFNJwfEJRK9QTKFAGYcARMOc8vs/2TJmEKGb7knH9
tckg8aG8GcIa3M9Dq52MxUH9UGmAfr3+AAkjs6N+mGtWiQ1cOlf+VBVnGY7BLmEkbudhdcV12qu7
/1KrXhaZPmAeSk/HmNwrAKplIWwbjYolXLIcYSZHEuD0+DpdKGWkfMd95ZYtSeJxb1Gy4augUdZE
aNNuFmqVU95htBERV4rbOXEh6frr2x1nH5oY/s5BIRQGo19Gztpq04bWRHtuFoX4Va+6vBzw+C6j
q2J48Q0HLvaRS30glQ6IvaS6DHTaBocwnNXMr+Qw+zP6NK2qSgLSjKidbRCJtJ4wR16P/l/rYJsT
029x/6LtucKSnxTeFvBR21J6f4u0j4/5LHpY5FCO8F1HZYqwz6NyACwSr8rokXARNAHOau1+O0ji
66RJ16S4ePgYT5gxMoJKX8WxpBIvoZ78D4O96QF+yTjRpWT1L7yrroOJrexcvt9WAsZyhu5nVsYE
KP2eUF9Pqb/Jd3/+JxyrMMqGfWGbtVrMtzam56GD0C+vWJKvacvftXUhmsSpVLx+ZNhBtMxLHTSO
rxpNLYBOrGPfmSvLzVFevWCrNO/VpgA4tQ06RJvJIx6VdlzNLLDs6sEhWswlVAXLv73XbwEESlV/
TcqBh00m0kjH4315iGQESO65nt4Dhvgl0ev/WjRv5L8fl4ba/dPoD4aUeLbCmQj7HIXesRLQ8Ies
pzaHgCHVyws8yHJplUwOU6KdAeDNhRkTL9Yp4QJpIlp1g9AqvsRGgnvXzQ6dATpVJDZLFP4dGFou
Bw7+CyXbcQWb+s0W+BOOBjdAWXAeWjP3Rjc0eMUqbANhQa/5PxjJMK5zDnsdTfBiK8VV6Dvn1h+I
jY6jdbWPPnTMoNgjwDqFk7vZumzC0z/5HZ4oOypBDeXjENJc4vW5XjLNAXh04oQgqxpbri3Jtv5Z
dtk1S8xnUHvDo6FhMxKWID/ERxOnPaM5v4M1uuz2bLm2mA2JUVrJMZris35a9uuYewxfHC7vFW34
csSfcw6l5xGs87brtRyQP8esyV3scXECeqxRQE8hFpxeaVKZvFxBPzV3s9GlToM5B4XQjoqaGbVx
ErcpUTXNaEJUyO/Zmt0SDMOYe8iX6B2F/ekCLT3PLXiRDJZrK9eufa5MilhrHV5cI70Ay+8nlBgg
T4rhveE02tI0DqP2dpk0d3V8f29ghBCJY74FXxTJgnp+l+RFLB2PvOY+wFYGcpLdL4PO/+7YzWyW
rhakOvH3Qsi45Al/If8GViGh6cS936cvJBeoBVq1vqySFE8JGYNab9Jjl17BI1mETsOYL9Ew+bDj
xbf4nAKqPPnDc9Xq+gCIr5cbzkJdSXJ/cqHlG+ewMEnjX7a6Me1xq8eyhHrK7btQx+m8zuDh4pEz
bOHXTzi4ZaHZja3X0Athq0fe9A0nlfy8Gextf9wG6Nz0erU0jQRxt5QBIVnMgvHdQYuxyELco7Bj
qDkAqW34fpNDiMcNIsL8ijAye65lxKOYxhipu6dK0CSBXHYkeSSbQHB3puZkw3/oaClcjOoQ7xSH
HqmPBXv8eHMBWjFO09il3v+9xVTT2vB1lZBwPxTVdHLvyM7NleaHOD5HtcCvRmd/FP7Obyl/w9WH
/Q7UTE9wUkMm+wkWtwiIA1d/78zLPuMQzap0D1fkGBV48SO4idtggZhBE0c+DXU0UMHSKzONon4i
PXiLCJn/Km30DwWOb1gchMBdARZSPwRAP2CYdcpND0pI0Z3QhRHgUYenK4gfwhqLtsJQDbMZy4me
aX1U5UhifXZdq/k4QgKo7xET5bS0ugCStI/fFafb3cQ/EE+OqX/oyBXOYwpNdCEQC5O4sq2IuXxM
FmWvePzV3LaMfcp4aSIcA+E1WCI2S9t5EQvLUAYRorDAgIYLXJ+bd6nptsG6X3b4ExoBjo0OWvKR
c78ywHFJd7kSG4qjDvmMyudADFLNT4vXSLFggdXEyRuFP/VSGtFG4DUG11IFFxeNyCu54Yl75o6f
oKBw+x0f++uzWQV16Ji7tnXuzXSZ7F7+sgJzaL+BS64lDHxZt3/rqwqpu0+NyIu+GZudZg4mTgod
Z9857AAewkSmQjwgThivKEHDTRm+4gr5CslmWz9XGVdDwNQ0QavtLrf5y1iJ6PHnrwCqopI1eSIg
YEpKOb7pbX8DsCH9VtF/31GwvBO7dxgPCyrRWRkXWoroFIrQIInR4StE2rd4wVUR57iU92dT/13T
mZss7AozK+xY3iWslHIxk1cwRl/fwGPNNsPZjHZmoLIkFud1/Xx1RW6c38qVY1uZU8zFxlhF4er1
lojMyHdxReeRRmkkKoNwIFd54MlYSfNVW1mPdxniZ4HD2mLxm1+hjE/bRiL6toQzkAr5Y+blz/T0
JOoQ4YvPDZ125Xev/31uKjBjSpI6/pL417rxF7GD6r2Ckdl9Sc0ZMEhT+a8KsRj9s5+sxRyCybtm
kNsJbCzkW6hNItncId9sFDRK1MHlWSmlcTdvpjuEO62tFfhJuIa7/o2dcCA5sB4lJ/LdW6tRrn2X
5S0t+cmXUvpJmVz9bJ97rSq2KGWZriC60Cl2JLDcQF94ABR7K2o+yhud0ilm0JT2qk7q0PZtGt9T
/OuhDcTmodLWz3CQgzDJLOGFjgess8EROv7Pz9pK0AsVIT2GGr0qUoys/4arIROYo0NVwafuoShC
8bkkNXCBz+p8CNDR1a0HocEbVvMSRZ+X/j9erJXELfzspXR6r+NywOf+XOdrZvnwBXKaiQwqb7fy
yguw+koCeP+HhsiBrUWEizgN0Uv2N4IhIwCXctWHrYhEbbMOpEB0XcuKsi+e/jf5U+n0lu6cL7Sn
MWgu376wblGEgnHi+KrpZnqap39zwd2y6l2/oO95+O6AjdWk4Z18ngBibmXF2lFhvIADl+hWBzI3
HY1XPSnNJTzkv2npdKBTxXTrLJHdX6C6FM2Z96Jk5TLzetlwsoGi0UsdNWtFvuf+NngMSJ4bc5Sm
GKE0+hMbEbEcyWF+igX+whXJpbXNH5yiSBQyhttHCoH3EN05fh7PbSzOyFyNXgt0g+iLqo0UoZ1j
wuSuIqKfUsADoDa8PSRAxd5YU8BPNiSHqciG3ZJPSBUng/I6ajzkKEx+VMZMmp7+mXdu3XIzsATw
YsyDyuyIEbb4q+0tkERtgwbstbGvIK7KS5Sw3Ug3ns9XnpELpBU1ZJsqezaBPOcgRTgLBxuOrd6d
qis/Ac6JxWj9z72vmF+LRq/Ntbvy8l4QP6DQUwLHhQWQgQFcH95sSWv4NbZeCdV9OnDFpQ72aoAz
D4M9FwlbYk6IEiEH/e7xA89bhuszEFIG0fgFbl6atxQQh25SpyGffXrv0CcXqxa7bQF/UBNVb0y8
2QFhNsPi+WEtgoJo3JPHisKoFjebAcMkZieJh3Ui4v6aL3QcikR76cvAvZNUvNnRMAJvnC9et3oM
OVEOz5JTomaon1/HvxXj58vXFCAgFcIoCaGEfgOFvVhvJQ2F7pYMkVu5rOpWs/RUIzDBvrNhou7s
8b9TXeqBA7Z0ihC7QjpdsfyONbOGGWk3E8krz4n86isYaq63CE+ALZ+XtsaJetkYga7hjUOj56z7
6cW5YXOlyOj26kr3rFoxEXIEb47krYbVkFDhLrIhdG56Vr6jW+/Al0heMXQJ76WQ3BRNGbWTagQA
BnmPAf3MEECXtxVDGBkFt96lQ9IUFbh5dK273ZfR3xDkDpu4UV3q7q9vSxSmZ5H2JLeE23CT9Xvm
PXS+I72a4o/Lk+9H3N1ZKdq0OZbWst3XSlI1O2PAHyEOLVQZGJvjUVeLaODw2TsV4uzFzEaND38K
J58ZaUbB+MPaHSfMeM6I3jgvzNKy4qIu69SdCeV0/NMpe0+Z5NZDGFk7izExGnnEKjOIXsHqx6bY
//A/djp80Oe3mJIF3nKJY2vcf0pcqPx6Sg+BHvyp+0EwF8kIxUowy2At5lDTY1bdU8pa6y9ccY3o
XJYi0EzKH3kSCXkEqrkhKGfBLzwXmcrRGY0BMdKbX7F9iGVdtlyTRRzhalwiwg3HwNaqMfAL+84O
VvEUQ2iqocwPVsdRYtC9Cn69ZK5sYIRGRoGLZRXnB7j239xHAuAsHFGJCL6oah4EmIqwPfP32noR
KZL2E+FbFBpAxf79HLdjKVCOHboODMuFADD8LCTKEcPk69GQFx2RmyCT4a4Y2Q3W9U9Jpno2r+4O
zS9aPgVUcqm0WI9mllbYX6dKn9AgB0ePYOfoz1qD3ozCSD1TbvALvpoxwSjMA4nanDzR4vWeTRCm
ndEUzugETz7BjlTaB55LERLI1JV4XL5nLRRpnwNg8Zy0e8SBgYasWD9tINBQagh2vRAsTY6YtjXH
K1kwYmOV6CkUM9ENl28Fb0deQYc5m9LYTEfLJpKj+GbLsb3/JPvhwN7C+7OLzB1TWZ6hfGrMX8wM
GXUK5CGsj5tcm38tuQ8/KGqHvYDoKzV6Lbi2TbKEIiB5/7uujhoF27autTfgv/Vb7g6TjPkipZiI
f7e0h2yYUJLq6sixxZFHnRSl2M66L8ETGXEb1RwseE/kie1yXPdRiVHnwndWN3E1fkYpCTLp3VDf
i6CMX1janvTGNQfFuFKTJb687JdRNUu6j1MaSGPCPL4uUdj9FBxjdstJSIsK9iRyeLSGtQNF4U4H
tn//LKAJtgs8/N3KMplu0EOZrJQT15c+qff7Cp8ilFqSD9zQwkYOK64j1uk4Ehh0XytmULfitvAI
DsX2xzQ1srlDldF9r7p1BLLdpvsZsUR4cC8EFYBboF3D8d1IMwQ8gpUnTRkvk6nx9KfXIWB+O7D3
dIiF6xPPDRY8zfvnTJ/cBuUZ6wFdYyEG1Be/iEJ/+oOr101cm3yYMpqLIZaNyTazY5WbRDIgGcFQ
s1ItHzQfMJ32MH1kCRzBENNgv4vaYKUMJh/QFDJcHth0O+sbI9YpzTP0bXw8NWifW80D8OOvcjIU
2SylFBjGX5jmX2DNgDfG1tfOwVMc9p/+98/WL8lr6OzIo37Cg+uuoo3ZdTGmzIREx3wQW4n1gnJU
GTD4sasS0Nae5TPIn7xwgWlLQMCIOwakKw5KYGmZ/InRk+WeepGK8LUX/u/VBDXtHUwwZ2Upgtyo
ibdpUmtsSJq5CiU9OXldyMw5dTB5e6qm4RIKm3gc+RIAv0SozKTc5wKZO6I4VK9vugLhxvZTT9Za
UNiVUHXjz/nFofp4jSf5XYpt47XtFCl1JXdjogimYMrIvwjXQBnUYhmUWLaeX86ClOXBYN6rrsca
gWpAaSXYGy+jykX8AARskJRHUKXIN8UIYE2hBq4PfC51xS4WtHi/Bmx8AWR0axfeTsPymp3Zkvnn
cfBYJw8jG0+WQ2ZDzuzSRPRqJOMkv3IaIkmduIVlBFp95Zmw+60+/YRnjtUU8LgCyJgWtUjW9dtQ
qraHhIJoshijLb1cBgbUKg/Oi3maGty+xtkHZeLSZsNGuSs+PnPyIUb1aBA2NSWbmLFxioc1N/QX
yc1Vnlbj6a0akqUklkDC+NWEDVQAQ8gx3NqAzBBa++oe80cwtD+G0g8fAWcSKtGrEkPTtFqvHTV+
SQ6xO68c+dEZsjDcrw1FiRyF3bCGSTwcYBReAFRMkJ+zwGXpT3LOjo/vyd2RxWpAxwOecfL0u1nP
9xj/pCqcIm6bwEFGOJQmLNsgFZUjdrhW21+TCOXCXLT9iVEaRw6JjlRr8vnVe0bkJ+7NBx5/xvU5
ViNzYoVWSZIqypiQNPx1MEtH94Yqkl8QYxdcaNBlaeJeAfKgTonldWM830vuCk52O4IqKkn6G0sJ
tAja8Lw14J0S2zIviUIGfaM5/Ij30KqFO2i7tKG2fmaNJJ739FvCLO7XpN5/fFYDAenWt/uVt9oO
VSInjq0QByjFOX8xocEwXW9q9XDKcOGwEJImfjp3A2K5IzxpSzkKr3upbfKYN/SKu5FyTaXoiHiU
IgZAO6uN6IqkT7oQ6IgiGlz7KTYDyfzeeUQzbKJUJ2XljJKMjIeZ3+JoGycY/+XV8F2BKzUMQApC
l1kGIRFjCeevkXXX9fjxOYFGxNyAZjwgs/JZ9/E4RXs3zAyJ92AmGRZdv2DFv8b6YTS95pRYxxAK
iR1Cu4VMdVPC5d6RcvRvxPTGTpXEtARLZKHVLCg/h1/BCCik7wYNYgIIetIU+9DQZ3XIQ5Hs0Num
5wBpNA5gIkiuMFc68O3gi40wbXWwC4ztxtlTvVRPqGdj9FQHkPvb8KTvsIcV6yWYyn5vTj5j/LXx
CB0gaAQVHRVx6hKZ3zkotIFYacJHyqLRPpQoulEd0szIwPXxVCanuatFDuPISItd9GphAme441nN
uwdz2+sjykyS+RWl8WZy3OcsfTJyoBQ62TRT8nkviTu1lgg41U23TpA5dpJ2cPWk3HCureG26cMi
S+g9SJwpp7hdO5cmf/F+ZJvyliapqjkG44Vouf4GTpS9gaYT4xdEm4lu658b/7PDVeOmmGZpMeAN
Vn2hsr6uH9IM5DGhuSnMwC2G+2wsY7CeeiADBe9yyguMgtgvs9fbSTdP9JCa3FKWd70GENx/Sf0d
KId8F/7FKXXY+rNdFp6I2s58hDtiWzHVrb8yyZAMs9WXC4AtL41i7HFgAl9ewcJEd5Wfa5FnDjej
tbUF/DDeMFjvxBrIgNU8jJK5b+Do0NKaEgVzzxr+FYxHp0k2enacInR2Nx7ghMQBEjz11NyOedQG
2hK9LhahDkmyPElUdABn13hH1xnm+KbwWAKeQ/EhaC7k0FVLGAREhoMylj0Ef6LaFcZiWmWno88O
5pZabWfjZWFybPgu+jyrPFf9ZCWPy5gKj0IqagyQqADDRpQIQJjUQFe3UGv2SY8TFud/qZCGAmV9
WPO+b930MskpkSBzhkCGX60+ikUtJEdaSf3PXxLy86jntvgt4LFpzQVX6Uj2tPeC/TPxFpjiXe3C
W3V656fxX+0Ok2EcF845YjPm4S/h6JaF2aCvvPTiV1fYyU8rpaNS3tiiA/tHVON8OWCTA6w/MeSc
FWBR6Q/TVcCDaOgBiW11WPfNVfX+UxDDlWTGDzyCIzctXjRoHQ4MZF5Jz9h8liQvMcF6Qw4Or4+8
3R0qR51gGkWxqeW3LVAgIQRl/xoGfNWRxfCz34DadFwUo/AqwWEZ+NsJ7HLsowaAbDCaFYcb7g/8
Y8Xv0Frs8Qm94YG40Kf3+tNgLZkFoM1e/5NnJTyovMI3AL6DMYwsg+RThv3Ez/C7uBMwHMvhfqLH
znb+rRNrfs8VhwQOyrsoXXo0qts9YUivPTqlgTlbK1ss0hKYqsN/z1SwJ5qMDIC4PQvbnXNMfm17
uyrdUg8ZqE47NS6uoXKlmvjR9E6j1SB+nFJRgM5vcY1OGvrsGFgfU55BWJ5ytTtNuxmFXr2YGa3u
mmpXk+bX3JcifWHj9JfUowIG8U5xgDgftx7HniFWqyxzSXwlwd7EqzR3PWhcxW5InsiAswZw1yhU
6mLtCUxGK5wbn1kQ+P9LHw5hg7lArotU4Q5tW8DqN4PACSklCTCvPe9ztgmSR4JV2g/jAastDrcl
PyNqvZkOBDq+ZyPudYXukCpsrH5voAaNPUb9YPGdRDUAIbNL1bHgKMdzvz6nQkgc5/sLTD+w4drC
a05jRPqV3Ully2AUE0raAHlvEkvHiVp7IkzQUzXg/jP8bV4VW1JtBdzvXLx+uFNKvS5DsXL0pGxN
fJW9IyPdx8kPZHgilmeVFHabphA2lfa9yxPteqmeufI/pVP3PA0FDHRlUDAS1N/iEZZn54eDLwR8
bSkjA3d2WjqqEV/FcXkP6DVej//fQbUWy6GHF1KicyK4/dZGRSXnY8VE6OEMRFD5FXsNVJgi/8gZ
pegK1csSJgMZsDbyiKC203M3e0bragfH7wnm4/Rg5o8V/e7OfTA0z28msYCXeE9tJqhzwtias9dP
Dvtgd+HLi6/xZsFPB/VzkRegugP83vtMP8BI0rbpeYWXXn49wmYrB9w4bW/HxHJCI2/TGYk=
`pragma protect end_protected
