/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/y8t7h+x+Jglo7rP2r7/SH1cr4Knakp1jFPyXfngFbBlYpsZvUNNHL4T
KIdfbYhRBjnkzFS9q43SIkh3l1200DW/3W/fbbgSm3OjcnILJ6+H9GXQh6lB7Ok5mrm7nc6JJo9b
nmX5GqqChrdPN3P9pKDDPuwQ8FES/1SwuUfFQm70V2NTxyEZ1CBN0qJlj3eQtMWuNylZ1efV+BYc
P6WQZ1+HqW9nX+9b64tSWZX0obb7aOBEalk5H+a3VUapQfZNqqFlKTu8BsE+o/8y7jqA/SqqcYSu
Ur9qlWaz1NsUGtqkjGAvfak3ynp5xdPVQn9sdAkYjTU45iGFmwyhGEsnIt1FhIbqI0v+o8TXAI91
fPHT6bPF2RXEgttlO+gCFyhdKwV4SCcNfpnobuHLW1tqSnm3A/R9zeX0sg7PCkGv1BArrCpbdOMz
PUB2k4pAcz5knn/TABa6hAnztHLsJoKtw59/O47+QHNg6nZCclCce8q/gkBn3U7O4uNyeGiH54zE
Y0gebMuKdF/ZRHEzDNEwDOP1cFhEx2IJlG3MW8jbuL/a0Rqis8M0V+c3N8BT0WYZr1lMP4ihvw2B
4vvlir4hZeISYcHp22LeUkXIPqmBbyHpXJQdcOHzY0VGPIaEcx+y9FQh8qw2xh8qUjrKPiAABicr
FYSrGrUvonpIwN1l6KbDyw03PYCIZAbvyjkL8RNPAmJQXxU0KQTxmcmgFhH1B/leQfIcrJKYhVfk
Po2fJjXh9ESnfV1FKBVTx3x9FGmPADbRzduL4py4ONOKI/BF7i0I4D8vTDD0dsB2dGrSi4uWPoUp
BjeOfTel2wOMASodm4VDETVenZWOlXhgjKhY1SF9S4FZmvbB0co21dk6xLOrBOlB+NQBU+sHrIUD
3tA4HjkwlakXlutxJph/JiMJPX4Fvzidb7bqrihR8eLG86wH2ti8S8YgRX8LSaZ9ypucPrmP8G6L
0KTDGkMlsYdDyO4xAI+zgpHvx0nz26ddIY3rLeM5NqF0A9FDfNih+BGmymIbR8ie3GCu4OFURcgK
hbG3eJzA/jjEIQhmMECpLGYjcetYP6E3KyMXHR8SsCR5QbWd79kFMDhcqgnwkxl3wgN7s/fGxXKg
eIv4IVDgPvu4orFENU2rexy0xn61uk8/z/80ttW6yDG2NEDxr5JTvuKuyEaFtao1DV3zoNFiDG/X
ZTkhnCFYx5v630k92tyAW4NicVxZCKEE5zRzrRA4Uu45+APU07Z70ORJCD8nHM4TXzFTRapIN/AO
xGjW9oxEKv+o7goWpzds99Ae7/D0RVg=
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
