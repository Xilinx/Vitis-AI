/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 301456)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLALC2JsJjFocyaVPIBk7fAMHdIuJsgvqr9FQ07+F3u14b7XQbcibIKtNG
3frss4J5UT2Cl4zYyIMuw1+DRnYAZLl6WEz4yhzN/UYe4lr0UfYE+DzaaKuM2nlxWArvLafGLwyZ
W0xsJMJPEhzW7IcHi/bLtor3dXJ0/gMsP12iQqisw3muHuMXnKWJFv9I35Z7i1DH21EBqbiVRtuD
Mewy2ssJCIcaPV1Zl/YivqOcyYdM5TkwALKmDq95eigzx9Az07BFb5u+WsNZ35lQiBefGJc7oqXn
iRVtKjtYJpRS4usmkz3oOiElDkKulpWugv2F/4cErAWb48uimvXsYkrAxBBIRtVxCpwOPB/CcgBo
gMtBsbg2J9hKwMRjEd7ri8je1tjeN8pVczALjHI9d7aBJ2n63vzTO5plPIIqOrp/ucRpJScxvEFI
R9roziamLmZQ4cr95hoh95umk2uaxWIGX/jcSe88ttjF7OCbAPIJZDStlF9HXkzOs6n8Gcs6LERb
lsRo2WoNQA+MwCrJ03aMf3h9eK9T0VaM9pX3k2v2j2pgch65rZN/PNc6vbj2bemFMvFEDNRbCrU4
hRKgxlS/EXnRw9AaHane3qGmvu5UqV7VIB2mh0mM2QhM6wIalfYt2h3TNaoADd74tzo5evHL5t11
4H/Utf3BBBY4FlvS9Yp9z87YAEysXlrEPkkZgMbqm0HBt3WrbeQQnM5SkVoSVapHNhX4PUHuZtxv
oofeJ9FSbGf/hgj1WLFnGjsAFglPrhcWD2PZC8tr4FFMz6RaljHpR2XcRbFillgg/Qdn/N8paFgM
PlmJKZDP8vcwxxDdcsKhiB+8bmRI4CnSY6HBX4667LWehW8ybNEavRtKW/ZVMI23+iY90TMqUDfT
49xcNbLmmI/tm6plw1MPWCMO+3Gp8lYIFgtvcAiNoBVmbNKEZYlPUkYxOA4mdkrhNzM2R3YORThe
bMzj68XOAYTAW1m64M8vKMzRIsvQq35B30XmyEKMzIcXIoiCdtiTv3DwO5K7VBueK9l8oL4woq41
8Gh3l4zA+UH6PL6t7IxOOjY74xICV7o8UW7AaX5UCCgZ9sS3ZLiN4h44HWB4fsoMo6JF7P2/U3Ok
POqNLbXI/+kVW4DcAR+CQ+LdHBYTTl3PkMq9114ZI9+oVdK9gtVzqYGeYuHv3HiDbdkT2dPHmpvo
60SEkzdKu8Z7bJ7VUQCut9i5XWJYQTy8782A11nCvNxXLA/S+kckwjTfCFFBpzRgBQBV7AJTsCV5
J7gBaHAG58x+rzouvvrjPzKbjCPe8LE+3cGEmK8eudrf/iykfnX13q7QMoYq4K7zD+PlDyExcChH
vefQVEAZCnLJZBqrW8GD1N1JYYqlouT9nmy8rrHTqQq9G8bN2zXH0cqvtoaNTiIO923ioTZjnK7C
O9PbmN+1gSULitZzSJQvGTDTKuCQLNJjkWQDLoDwju+G3xYjHI0vtcIso9x+yrwba8sUZFk4mgU8
1tWglDffHXmYxvBV6JdkGreh680TSpAsbWc7jaUZOnHHoQI3XfTN2vw2mpvTPw3c3RLO3t14+omz
0RpUSpVAOOz+6wqIJGCImZ4vchSm1ezy4cwL7xguRt99GP9DblWQAI6i3uKv85CQHuq5sNIFfPuc
c5H7YSz64CoQmmQH8cgZX7Ad4azWhQ2typRYBcKcMkZ/A509E0YeC1qhRfujkogohOBLeZV4fqkA
I6NDkcHW+Tk3M7g/ljKbz01n/+cEpx7arz2q2rnW15ZMXpYXoWtNBzA2M1EAuyA6O4aSRrqpZlIm
uBvK+ZTmoW+eodhIBkZoJbdurUs8IO8Vs6hCIychWT6LDqxeNFVmjX8nRLndLDyEFNbyeHRQyscC
w1AvLlCZVCJ17OBv+rY0TtBT1ipcZcZjKPsPsTCyYrdpVUQBXtVk02CUvuWu/uPCkoeOk3e3fLlr
yYDFvcw09UWw0gFGWbcGCz2HY5eunmuEDLZm27wYS7GXu4mEfn3HWRiQCqCFqjqn8DNRUm/z95QM
flFF6H+u2Owgvv0ygZ/h/NOOC4Wm41+TnN/nROkfMdNFzsa2N59FjzDTNDI+pah0DR30b4LXNMFg
BdOU27Dd6wjvCzHEcPaUmIS1uCJRpQJd22gYVrPAWWYt07OzJZmP4+zrFfenFL17Ivdcq9VX357Z
I4Xt0SziipbU4W6Zwat2aqTcXBgXQ3JwQRXGc0Gmd7BrbLLCUIxEPXE4t2xV7ZJB/SeFbYEJxex/
wIYdd3YxX3MWJIWmoXNEKFPQ0wO59UrFpo0mB68KoVUiGVlefFdtK0j8w2QGGMk1MLuMU4wazRGN
7MhzvGMgH6EXEjAau8yL87LnA6JPXDfB04rxdy0wHZlZkoLRTRlthPrUi30xWOaSiCJKBAHkR/Dp
66l3i6F0eVWvDsxBSz/FnG5EBprB0P8ZxB1DzFjorcO0DqB7bq6k8gXqxCJ32Exv9ArO59866ehb
SiAQzEVMVsGeX87Yj0uYT1a3WjH7HJfMiYSpcZKt6NF0SAkFUpFbE+mMCJSWbbcSAOjy/Ejt2iJq
R2ArqO8BFFUjzUHfEdZB4R8f8SYhBEjNxLMGR7Ft97V8p+HkghAN7B5y1bbVuVrkEygB5zySHa5g
gG19h1j4cHewxiDUbCLX079bxJR7d5w5vVnzJBqn1N9mz5lpkP721XfJS9WBnYA3avVl2QAvDgnR
XTuCMMP0Stxw8Taf8mtYvHcGoXyzn3tFmRHnwf5VD2Q96Rz84Ar3EfZ0pzjBqBtdxQccBehFkA7l
N7uyzc4Hc3VgGUdM+QsNnV5TotoWX5lgbbf8PjYV4p+9rL4AaktflNx6ZOUKehY9zG2+O/qY0Tl6
wkCZYejfblq1LzI0ULX+Kh15rfzYZuH++TizLxZFSEgWI/w+TaGhZarPQgostJJ13EH4Pbt1wWCM
7XXxEjPSE6MAdd4YhTG4Bfe20iNR8S9tEPu8aW4homb9HeYDjMj/CLGsW0r1oKiaNZtTjbZEyBo/
ChhafbvIPwr8OW1BgTwhoFGO/KIvucPW4h6XPje86cN5oqLxmrdMOkzbrREhuQfgZoFQIP7s27+V
2regc3+MTNSKsyKbmGNS97+rmOMnt4LLclcRSUwGMiQxHI/1bZP/Ej3Y/wbrqXSaUZEGIPHQBCcC
9E+Rv/FlI2J+Jb+FoFulvbMXNmJWqoJMSiLrbRIr1Bt7EClYEHrVcWo8GFmCsnCU1OMKenoNKR7/
zbieGfeMOJJCu73UHobNx6YY9Sb/bOu62VlY4sIaGFjgj8tFsSi8XWuz9U6EC4AFXFq/VV8fF7r5
tjgQHFnmfbla1viRBwf6aHRZYO+iq5K2BBqnqutazl5hbXOiRFWEUrANqp9wk4GGEpU0jtMuOUfb
Qr/jtHejBzg2NxkUd91JxwiqtTBXI2LIYAE73SKED/UM+5SjnN5U4w1+XLNhYEJoy49CFYQ8Rtjw
ti+6qNkLC9vSZxiEeQEXKZ5DtbZW+zpmTBWebnG8ZR+9y2jDepaMdtzD6ZEGfrQ56SjQQ39gTKFM
c/HjgZfr9Cw77GsFetVNPaYJlGXvUC/oEXs7pTO87blKk+gYEi3avreMxIU2yHvLmsYhYek67PGJ
uo415VPgzFGye7i87IKv52pbrRSDKAsmYxxgK8EJmrsJ2rQTEI86cBwZaU0RF0deJWVFnd8BAWfn
bUB1oU4DKefDKLy9gFMO+2Wwb/L0SBUuHU0DzrX8196ZSiapMjJ6atIyt/xxylLnbmpLpk4iB88g
RV7lIoH6d+kDVtPO3IiCmD3hvJwPf2eHEooed+Ne59d29sRUw268jkraufjdVyHlZRYSBCkiJ1mz
JGdqx5ZbwrvYWtl4y/jk7vNx1jHYaPslD/4EeCHg7GK9AAs6eCZSidgipG2BEX2QvgSABtioonEn
69acWk8dBKLL5yUOuLewWvuYGbELUvEQWmciGZqGbXRUfzPhU1vhtzZi73umlgQKRmM4dhIgUfbd
PqUUCOsT8AvO7FZR21A1TxvfxC+yediZlnwCmPxVzCwxt12P+3KKZCyBnipCGWrBIKfbjLHrgWCB
HAuITgN4NwoKxpNUiJSKNnYzY+mMDbW9vGs9L61dLN1Rh7PCQNwWcNlCt3AxWKkecPmc/30c4ayk
HwL1rljbFPI+cuYA9i369WT1xgyBWC7AX4YnWLqlrAzfyWqK+YvZrJlq8Nfx6X+q/20uiPQrH+gd
MgjznOXUqMSBgAUEkR5cMNZBrSDJv9SzKWJP4Yi6Cu/jxxtA+a54LFfg8cnh5FGIZpMBoI8WeZD2
GMAK4AWHaw8XEVShoZBl+8yhI5kEvxzB1NEPA8Vnn6TeZWIe5V20ODtT+42TuuVEPlA+LnkMK1xe
2lyUBxg34llF7Cy6bTsPp89GdCWKj34hbJ6UYmcnUk5qkUJhsxAWogX3vEEoDkgOlSVlarFQOEgf
NIqfpeT2l6GQ57IGy3Q8ZGkjD99VUEjNS2CRzBHnvyOFCLxkFURAz2hqvQbFddAF7jg3/ydarOc0
oD//LY4jfq5sg1luat/jc7Ps74nkvhESPfMWNBU75PvjnS866ltuqGzd/HN/JbVzGMPsrkg86QtB
YInos5f9d07Fdo4Ht3BqLQNG/5TU2BkMqXPpchNKi/DsoS3jk8QDKq5OLc72yBQ26J1jdEaTieA/
GhRM9YXslv1ISn3EwmWZgcaTtiBa2zAe5/p9XbIEs2kOFq9jM57p8yJXsP7hyFyX3cwvcO3/e6yn
2QST+sdLcVxNvCuR1GQmmbILFXn3TFAVxEAY78m3JEwrbLEQ41roQAQE84W5pNzizx+046UiF8+U
FrBJRvPKcJVOWdpCXSbMG7l7cGy9Vg5YggMLnVJjMTgQ1d8yuKA0qESywYVvMfc5Bxu5vz0uxEFq
AmFTJH9o4Sjabh01QfM+MoQ+4554/TPqyWf7eQXu4ZRBT62MB7v3Ti5Zx16o4LzeCNRtkG6WE9o8
aNvk9rUFFeX79o76PDd1UlPpPxtQv0+i9COxLVF/5DeO5+nL77DITRtXI3CUS2s2+ctCI7qRjMdI
PRlvUr74gwWcuiDg1udj/U9bnS1/WfbPauq/dBWLSogmOLIaOZTFhjvkEetsVbU56lz9HODdf8Uc
vqH0y2FEtIMZixraEPyRcz8K+HJ+Z1+4a0NPkXFZ998Nbl8xD5uKJELiXa9TYDHvviy8l1fur7w9
xW9gBhS9krMbK+BbOoypElS/3gz27iH6fmaZHBy+bFLfnzi6KQrPGLHUHJtmoS2Oe+Hy2U74tPdv
D1gSV1dK5R8mibSINaoReGBXagvHD9iTyvwGhNIJMVEEgkW/dDySd7nc73qRubdWVtEFhONxOvXO
ZzC1+hCuQ09fLFUx1vtXsxnwWxfHjFbmiIUNIxhCbsCTkBZ+N4FJyHKkMRJBgMqXTJHZnVVbsXic
ZgGQJFUgxQBj9wCrKfickfxImPHSTZ7PdQyx0PO4l6E4rFqgJcVRy6lPXe0AtOqTiBetPBYWtK3Y
m4IvLwCoCnyPcketZ8SiyV06g0/iskP94sCZYDTn0kINjwCExNt8okziWuMv2SW5y6NVcYMBdV6e
eJ1Gem5+FPoUkMB939Qz91EiZOzTEv00B3tCtCRYv3elvhwQketEemjC67ec4GC8GUo6bJD1Yt78
r5Dm8ifr+MPc8MO6JeTjhOFjcu2W8Sa5rjrjTHwLFqIZadOCk+dW5YCRSFSbFOVncxvdxSmUC+VL
Lfdoc+kgwbo2wQLnfnidyhFCZsoRyI9sZ0TmqI8B/qXbPbaHLnOXLk5D3yuHxyBoGRWSA94Quesk
Ts+AMNWvWquYp1c4Vg47bJ1+lyDQdxrSpAX1cqzcSIMKVyh9B1IQyScwvKP+hU5WQ8vCJDIAvXON
DI2mkJn/5RA7SEpdI7iv0kh7e/sOEwl9iKfRnmuvZ0kHbYqVl+4P7AhyM2IyhosR6oBK7SX+24Lx
OTJgPKq8YgSGwJwqiKgY89+cy4ta9dBP5X9SyLfEE8oZo5ogWpTbkH0vHgdsVmJZ6IRwOQdMF1Au
ga1i6orAqNa2uwZfZ5T5tuqty0OAJrM6gTA053HxUSI+WZM/shRus6rGF4cCYLXba6Eae42ZhWit
G/1UBG2fteDg7qMb6E+z6O1jhaWXv/RdF1dqWpOvQo1C6YSlWLw1BUMf2sNpJ+oRo9uEqI23aRwr
Py39ioDrIPJELpjwSIlys+kYlom+rZcur2Xs8rE3sg00C97/s5Y0IonD/Qp5kcyUcBcy9+DO9SGA
qVHJNB1hySaT2xCo5yrOTbwOvnAThcRHOcJDWELG/bOOgX8lD/FUl7q8CAf6kD/b7Q+GYQkkAN2H
9Hq/Jx0NyV7pFr4ipi8vUKpJo9Cz7xZnl3KUpSAlcSmQ3GVIulBEvE3c9Ia/P2n8BgK8sgRC9mOs
QFPjf+HfoydTwmEMtop7KfFMVUlq/Iyd2LQjna+2NN8nVIslV4dQrez4Ybz36jLCeSzdkVQlIQOK
GY/RMgEi2HLRZMUgji4XGpxZnySHcJ09ihNT0BbaUjbRFnxQGw+iymwlCDdvrU/ka8AVBCA4jOpe
DpJFTMBTTDL3bO9cxfSo59G5M3dnJK4UNkwOELsA+rS39ZqbsI9TePUIITApKZc+ZgfwSiLYqBFY
r0hQ5rXU3x1V4uFCHG7MaqOdscv+HHss482+6cxngEoM+xx31VX9ZfZJMGIRyW7Bt9t+WRT9K1lO
Q9QVkIIw31kJ7EucSjD2L5DEqizOT5mVi+RXN0pb7MLkaJrQbqcwUFRLcbu505EsFI1893ZZIp2g
1qPo4dDQ8kq9pSALhH6BSaUotEp9KS7BppOp+uXbZfwXMUlt3lipAXQx/IzH6pCRYTGyD49CmUnl
tXobrd15QHiBh4rG2y8fZ0WLg4bs9KkQPv0e26J+d9+VZ3c5yymftk4v1EY6ot2wc4wauXSZqDsX
wiyWoLrZ0FLoPafI6RpTZvkkFqE7AThOFqvAr8ZpF3+mNofWyOO6WLvkfxBr8XCXskr0H976zAMX
7TTwh4g0urEy3XpXNAb/KbMcbYaIHZce2A+v1l8orisL2AXqoX1ELObRTbH/BOEBpFXHdgBLCqOB
cCapUgzFQZOWGzLLiZhv2IDjeJKWH/6pqiKXa40bOnS5fyKTTWS7+GCfC5MtBR55l2ezu8/pYJz9
3VCqrIwOUrpV3Dpdy3bpbBmS2DLElP0U4tHGTJnZhzq9hGwz4VwZFlXMPa4eIi3EmJOrdtWXJCRs
QjiAG8hYYjD97RBleFCsozAZ+v2xX0bME7rKLmF7K+jAoZE37OcM27KtqZ2nHjoOew/sW6Z8pdYb
yfiyxdo23oKgPG2g37eIPpD6p23u58uTl2a/8FVvE8f8hfp4QQs4ekbjl9Oj/BZik8OFkX6u6dfj
aJRIuQPumY+wuIGbOS9iOo+lKuJSmB4goVH6YSGbwUkoE51LSne4RItZX0LDySGiMAo5XpAExP2f
KwyAp1+WzA050pOURAl4i2lAxCSXp1CmvMi1ZXFA3DBml+SQCmvnfL9egtN8zoU8YmtSp+OHcum5
npL6EyaeJFSWmCoRjw2SmZVvOUEe75PxS1bCDxxiyJmfsgPAKBRq2Zufu7QEhAozp+M9ziXQ6rym
WPLIhI+MZSp7YWu+WmAboFe8IJVGL4TgX9oPJRu6N2K6jRsxxea+QpZGCmtMMbTPDJsRXRNU8ihF
SrEC+hhpJ7Yhm9a1za5P1haDyHc5k6imyX+8vLk2Q0blDk6rJH+EskBIOHSrH8rpxLe1qBu8xHg3
/QZNkNH8L3gGtcJiw7O7u+qBGU2n9YwdR048Y3b8wLrwJp0bJj03jtDAudLqgxAlEyqK5Xl2kIGi
DfqFfj8ep7sRGkTWEHLs9vMT3lcemAOZyed4TwHNIUj4Q2wiL2D0PHTp4QphgFrh87a3oHxGyT1Z
2IqBFV4e/Y+iU7sI0wv+Eqqn2ihAP16YQ4ICDzlQ+Lekh54hGwPbqq8GkfNrbvGuknE6RjnkKpma
8D6SbBFpMQA2pjXVP83il9SSaI6TOJva+nO9HiQw8qv8tRbQYTKs4xNFj8AqnRsiOl67thjwrqsF
BQSpw616yHHGDlt1tFoHIIOLH2xfnE9tYBF80mu/g4dXlv41QQ2ROg/NfkSXSmPc/E7LL7OO1R5u
11A1KzrJ3QgGb4+yfOssQ2d98GPugCpVXKFN1Bc8rhS6zthBeNTMfJlcfi4UHw14zdnzKRMZvJE5
n5lhOW4vNbOmNZppu9+QZSSYOzxH2sBaGdsHyKYtTGZnezuY4K7WWeCx4OLL29UrvbxCdJdqIw2X
+/38KEvVkadDqxYFISTY5xNX1dx0w0BctI+3pw1LM15K23PjrUiGT6P6IAsm8Vq4qgtof5KDZGT+
nlV+Xu+znaJ9K68ieOZnJXAWiWKkZ/oNOCs/SEn3YP1uAIR4Vm+QDw5OF/cBFvu+nIoS24unxEzL
DO8OaCe9+X01KijQyzqqwtM/F7dd/01qtTFXpMycFVpMEQedW3E7QAj/23BBXDhhNdgQK4Dpwwfm
9xW5Tlw8oPqSIQRSehyNR4CfS3t67lZOrDdhfuJ+KZ8O3BvKt9Je4wsGwswe+fk4DWZpoXkJz6Cl
gZWvFeoWaRve88TdAhtiLPIffXzoswR9gaGi+5C04+6KqkUgi26g8mnJ0np2TSfUf78/f+w15N91
00+cYrpGs4aNRauwLjnf0Y4JHRLQF72ohTlWocaDUqZFA7uibhgsaDVnJFKdi2aOx5sEsfuKwyCz
3KnV081ECuD8A9O9e440uvfvrGq2UlWoyg/74jcmOIalEDp+Szkyl8y4z9RhzO5WtFbPPySAbfJ8
aCq33dgHVFeCxUStbTnBg4M8Z3W4h9j/ETzyct2dwPorm+/F/dFqaDBDvUXk6txHUaWIwcVGX/kp
xLNLq17r9ULkRFLTQHGBEO9Ob20ZuF/lpBSrMoehwzsoF7MMChWF5P2MRLV30dmxUR2HobheIKCM
TGVGnZE7chJ3gDX7KOIyUHNf7whULMbXDfEyNh0k6mwJiN2Vz6RcivqgLu5pcuHhUQUWoH3/C5q9
nHlg4JXJY9CQuvlVHGWJGGbLtrwNSZ5I4VewreeoP2pE8VsuU+GBxSzdU2vZtHQIAgAsLuEfOqkS
IcjVIsYekKH9Ca6M3dN2muKqgX/k+ddvZsDE4TCJJN8OzGeFiqHCCQDZUZ6RqNI482liDqwJ88TB
6jOhQc0qT1aFZ9cuejEHvvW0eV7z22vlSpzk78cF8sEMFMw3YV/4H/VNXt30XtbC8WRHpqU/vS+E
WpN0/K5jA+hLo+gGgcJdsFKPhm8NDhZNrmEza6O5lJkETGRg6fPUInG90mpgsYRzE8wQvGBDMkhV
aL9Jbt+5iz1aiZAFEz6HTgm1j0x3ge772X/GLVFzY/Sd1vW8s3ZzyBzHc8IykBDN7P/Av1RyjfJJ
3t4udhWJzth2Cqb5Ew7Aq2FneruQYtmkocbOwLDqr1SnYkwakHSDbNAB80gNZRlRLoFT2BFMoiBa
+casr+fWzSBXDoigNVeccK4g3jfrlfoygTiGb+LiG3K4QLnezhBVPhBYrWmeC8JGC/9koRJjC3/M
lztwOHjEPaLouGidYV1YOWl0XdhKqTwGFuxbnH+ro8YQOJ6jOXbXQV0C6ALinuEOIBeoUi0LEtz+
VCQb4bq8S+YH/Yrt9Tm5K/5iD1alLm/wRQi2zeUWdUjFNfK1opbD6gNPy7PrS/hWqpKO6LM7EP5i
XuNZHrkoxTUxu/ixw4FLizmercJJJVx5tzn2M2ipHKHO9v7EmbJnEAHxQULXlpDYpmm6nZLeeiqj
aku001v0JG0wmrxK3lBSHRnVV9MwDQfAXCMgZdJlFrvaA4a8vELPWhpF/Jqj6QZ+JxcUHiSghb1P
CuMip5acy5uoaBd9bbeaaWhl/iQRiPxHBL5gl/TlHsGy49USiqXUFJFski+q7ro+C/1fDRHZZdwJ
cKzkI+a8XPZEXSfD+m6bPsIBEmWJL6IMKbJ+0NnZcHKiwjwcXeE9eqj3F9yWExpwFW835+avD33N
lAwimEi2VW1xOCCc6NqYrHbH8XUQR8B8ubuF+hqfLaQRd0JYzCGpukIo2iid2+IxIYhPaxfA+QNO
KmFzc/NWmQOS3z/QicPH1USNYnqaaWIdTJBgnVvYD/zA30UNdR4XGIBvfeDp+Ddcg7s6zAlD9T/6
/DA9adH2cYNS8+c6hKLvWL8JKIBleIjwi1dkVXuIZxSRA0XV/eU5MxMwrAtA5c50rJ62TxNKwRWn
BPciquIjKgXSzOmWsPedDPvR+sc7lGq1aChBq+XyflK1iJVA4N3bfcZzP4CwvfcCpDEPr1RkBir2
JX2oG6a6O/h1I/jDFY6+DLO7+SX9toovPuADheIv8/gIHBoRJHlkghk1oCt69kSBNDiHpDPEj41f
fOW2IUyC7HXUTzEocIGWMMw/vXjbHfC4xwHMdrq9vsfqJTd51hNguPBEqYqsuCZ18bJbDPguijqg
27U93g4NwPd0wMa+Q3jFLx0t8nElJxf+nb9tEUmDAwoftCcaKiLhxNHTbkXjPnCm8w4aV3fP9SD9
PeVFOEBCdf9pYOukjGAnbus9D5Gw3HLUCQiRr5Rd0DpV7FWMDs7kN2HcbQH1fCGuigiIM/DGdxJk
VhZpwp1VCx+eHQ6n9JFlRCIeOS1lfn3aQdSofchzuKCQR3UTOrKqfNIy0spMTicRa4XPNgzyVYHo
ALd9EnVSudMrhm0Y21jEQyQASzRYNSDFELjZ7ssTuzlEpF08Yx0jOuFQH+j56sHPqQ/aH/Xi1lCQ
ZLVScbhFe0s4IOHv0/Mo9OesQ0ArBPCpZ4YQdsLnUeLoUleHSVga3yHA5CKDCnOcCkcqREpNF2Fw
ERuX7I5zP14HhubRaVonqQL5POCty6XNmtLfMq5KwrNNJSdfd2JICcCgwGvMfZtYQdTAYs8Rd6/6
qCBYl3y+nxZmZ9Odt6SuzHNGhbq1kA6EPBdAIuv+5qxzsEJJLfnRsB48xzUSSKsSgx9XyG0+JXJX
5bC/H6UbToGfdNoYfIQii7+kZx9zqQQZFzQZx81QBrggDaW4y0YEtL52OSIba99fT/mFU2SIxsfN
bD0evClCaIRT59oU0uOqrj/X0KHRFce7jPhHLQ7/xtATYc9dOx5x8Ef5KJw5cUgh+oLhsZv0tc9G
oPLWbYve67qQ7F2sTUn2hXoHnapVtbtfeGH3Y7k5U3aRyPQi5FU1h36VtNzb7wksXN70HB0SRl56
FB4H2d+Aiu1juXiUs1LnXEXL9qrFjOKCJ9/se2Nf2tkQH9PN9kPPUE1mW5IpUdR6qLXjcfQyLo2l
E0jx0t3EYHoTjy6hdMHp5AwR6WK8NExQy4Vql/rBqGem/7QKvgD2j1xNnHdrCdw4Ty9epn7HCywD
aT2Eu6SqMO8C2n635sMkbYPScFQzr1QcXAQPEAAV4l2Xi0R2boRp3wzpn0Tac7S9ifSnNCeytIhG
z2wmvCJMEW7K21zV77Z4eTlqprohFptYfafC1Wv4jxlVHRO1iGavt2ajmgLa4tFCnazRJ0/k3J12
DwzOsu4kzZNi+mUC+DnGWiVurHlWf2eDTwCOukMyZVSn32suHm49EuWCnX1vK2QV2D+NfftMiCmN
qzFu4l618dGO9QFp1b69AurYtf+wPOkKkHi7DYn9RSzAA+GzBGxTFbAsA8CPiDpPeAP5wrDtm7t5
KXoktxxMFCoMBnpUfXN62+AJrtvDfXUBfTIAJjT5iKapLZc+UCQ1dTN/xUfexSPMAX3yd1ZC+Yeh
8qAt/RC4f8pCtjWtlGiMi1pzhAYJ+pI10rCD2YWrnQN30zNoSP+s3dyV38qNrVURGSx/e0cQTDT6
ZrxRpXb7MSrpNStxZrIB7YdGjZSmKlLCCrmoYmzN+ph6LlTqkw1nuPWOrdggoinv7poPtIELv8GS
D2elKH4peecuxioccLwwa/dVyluXbtN2vld51tUJL4RnbaXmnGoxnnmGX5PKA2llKYFRn/kdt9zc
IZLW745X2tvU9cQXQQ3zbFxEJ8CpNe8r1j8/VMsbKscnNq3BKK02Zs4oZ9lQaruCikNqhzqZooJN
7oOIjFr6yb47ALPNnnhLs6v3Ny8oTgjef9Pr04rkIK6EIqgjkYfxe3GRK975c4HXuba6J6ciE9Et
58REZk/Zzm6qn859gG4gShiT2J2cwi3sBOjnx4YXvA03QsfKJqQjcd1W3mE4GwuyHU+gHflckcto
WViZN2YL4gvUZtLb8RTzXX7XdcSDi1fgBmal2L12IrfNV7Sa/mNZMS7PfM25UxA5rH24C/pwor9U
eUtJf81KYmlpvGGwUFVNadbJp3bV7ExwCHOKUMqu99Sj+PKSbGAQ5H8cMSUjqKArrt4htfywTu+T
2FviCL4AOd+GscGsViY4Kgwv94r2KRge0B/AUdHn/jQuN5Us5L8cAuSmO1l53UfU+Gq111tRE3rz
/uOESJ0BKtPyKN1qbw2Vgx8CL+go0VmMiklIFdGa5jqEVqESalnMvmiVT1fH5eMUJps/8aw1QXzi
5aSzxmHp2LCBehwWO1Eqp1FKSgT6NpeIJpeXZWX4UlTSRnlB8onqVEtk7woatWP+FZuzQnf4nnZr
HTrduns71H4oTDF3UhQizTRHXP0PxFIBvhVxaoAElzDKGxkege+uan1yaq/hGgYbWo0UaMpBumWd
jmCA6wurRl3Di7ch8pXcNqIdd00CfBed2+SsLLkxqtW/uaId5dXnlDCK92fIXPr9LZinq4Kpm3Ui
c3f4vLd/iOBXrLXUxcX4WVCYIL3159G7SJhLuxZjnq0Cvu5B7T2zg7T6LLoL1ArSWzhpx6bZUY7t
my16X6MC/y1Yq8AkYgEoFniHwFVKQPFLJWM0BGMXanUrRzWtezU+In6Bqdf8Qxd/60AuwomVtURb
W6RUC+RFRzJOBvLezXztcpZ6kYgazIMoHD2IlN1cqDLj3tnos6cXR/CwwH70zcd/CPJEEfwe+hfp
HYtn55hdX0eZ3KZ73U4BASAnTK+dt2XG+4EGJ09d2MtzL14tmtyDxZsDD/PL6IB8oDUPOLoC5X54
jv8GBR+tDoYJjp1jj2cAFXI9/I14CylvRDUvOaMfIyyLC3BZBlB59jkJ2pGMbDIQlepCGQ6gGLBG
qRnKQrGbVwOvjXwllJXP/8iHB2hRNPAJ1fwnRm0rUzvFgu4HbNXxo8neYOE1yv8TchEHkMpQAPpD
50DLeKyWmmBvEpLnCvbhtJB6g0N0amLMKObAlp+TQBCn5YbUqJ7hJVmS0sTPt5OBk/VB23AGVHBv
ZbqzP7Lrm8Qg1d4h7Xvt5JJsJW+3Uw+ZDRXGQ0vjU3a4xyxSlqICwiy3SOMXXD3y++7ZVFSn0Fnb
kEM4cWaVMn3CUVRTgc9muyrghFrYWXixm0HRnz3kUE5kw0U/kT5Aa4YbEX2BvKfI1g2mujZ73Ap3
qw1mUjNJxo3MCw1ySonhEcejxZQUPWXc15i2SacxAVjR/AUtvSY0dEfelu6720cFj437dX9KKl0N
rT4v8NX7dBsves9vf15IWnSE1VFNX5y8jgc+XiiYFsUE7kumppMdv0oSgILeKFXMXkrimVQtehnR
1v2bmQTNn6L4jFGUpj7tm8dSw/r9I1sDAcTpcYXVpOAxeI9Sq5Yffo7RksQURoG7qHENo/a9FMKV
5O9OvNgkQ8sXh2twGy0eCguJX8LBVfHDVCOqYhqW/yu5DOJrxmDWNz9KVWUEVtO88bwu+e5xGyIF
5tkEbU+yxAADO+1Hml2s9f4KqUB1vNQmDJmjfUCZKJUxydrwZr8Eo6IFlyJGixu0R2OXNBKSRk3m
9JeNi8uevksprmr3vyU//75XTUBq2aRYi4K+fUCEyFlfYv6XSzkZFiqu6jLlqdz4j1sc5u07lx8+
18vQi6RKBP0trBrzK10B4JRXhs+mUXjPPFo8rGjO5mnZxDLLCUSFQM69t8K87tXZqaiHyVyufR1I
XBSr46oj4PaG3k470B75yXVpIWnH2BkGrO1q98hFrNJNDnUg9R7D753fTwk5Mn+ae6MFK3hX8TM+
ZuueUkq7Q1UCRFAicyzxIScze7l9KWwifcG8VRpTdDRoV3FXZQL5KWuwSYmLuBQmxp4cYsJpT55m
FYLZOs4dtpwBx8bHg1SVKWmiQN/BFg9lA/JZnbig1dL5oumJ3aWPL/Xadn0/O39gBbAONQqKKeIB
gH+b4iyW/LxPLqKFbuDBBkNTHo/8m23BDe2UpWKWfW2bIIzWBCPveBA25e5kUpa/JwfupJ8bJVD6
McDwOxqKOiy3uU+7Xe2WmV2EosbsnLN975oYE5W02kIK259RzGgZNcFeqK8EBCgAnFZo0CFNKD9H
r4PRf+69NGBLP0za52k3MBc5C4/ga95yUavUUxCphZUK1WJd2eZ7pQCWI5nL3jxX13zNHjlne+a8
l/GYYwd6x8zq24U04LJ4QUF9eBphVWl4TnYEuM1F5EFPv0giZpflNg3S0pLeTv1EwbOPwteGqRJJ
i6GCSjZJ7wEd2yOLJxsDo5sPTXnkDK8xY/X3KPUaJBsNYpss24BSxS92m4UH3aM0/ift3V6CFGAg
ziV3BYYnPFEDrqPjhNMfRDKOOWBHnEcWqa4FeHmNk93lts1cA+3FaiX/tBS6PYH+G2nOy0P9yRTH
hsgD+MiQbiOTK3dO5odpNucCgqDID9InoQ5ebxIvyfb2va7J7aGF1F6DfoQio5Ae3lGJ5zFodfe4
BWj03Prxn01v38ZSn82E40TmGgX0EpiVNySgapHc3AJFQVRnruDVOnYonXh2yaCkGChNgwP3j1MZ
f77bayNINf4qVq+pXLwnQufdl6fP4yTSaEu5OvIjcy7sjmBBoK4Y8uajwdpVcgQiRp34xHXHvqjv
IKParBUQRxwHKHYTZnWvILqfebQneGpiFaPr9SkGdWnH+opYmLCi86CXeQQIc2Jcuzwz8jRqxmpO
gZbS47Qbk7ai/RSrojP0I/4rR3Y01Sz4bBhyTAMojPTp9mt61LHb20jXGSaxw10GU4Q9GaENFaOV
CWLsob2Yrh329j/ZmgFqSAa4yy21HhVTSGOKJUa//zqA+71g0+2lgG+2Ewuz/H8nByEN5coR7yEe
7vWIvN5fx0aq/CIS/uGPHhPizkEqQduZ16QTUmGhmNsNT3oJD7PRhyTPtlbbFk10j2QF6PZoeCnw
lbXehG1yKNpvMNZ5gqzNEy1lg/pRCgESQi3ePnRGXU7LBj8vRtaVXV05/H5vJP1HEdAeLsBXpH9C
mKda7+tEqfLW2ligCRrpAA0cWKY3+Zaw5W4Szkk7h2p6gyiWlyVcK8VQ6t4uLlLdlasWOd5tf9Ey
AYjd205C+7MdO96P/SG1QpxcLHRb58cAeB4SJXruFvltCgU0sEZfpJjO2IVyOqCtiIWx0VkwKoOP
dnUJS0Ek5eijNjV6EeimUrHSfLGBHiZD0H2fRCgVuQDHGbV79an41SO5jLDSORX+ns/1Bfz2/Xn8
qMhOhU9ZifTHnV1bk/nAJ8n0IEA7gxcDfnr43+rMNdn9kXEHPCAVAA7XvHSsw9m6ku7KUIYZ2hfk
avkjNxeMHFyYcla93OZlEfMbcGHpwpMpqHU/CMlSkEi7f2gCNJ83n8bxIcPvt3mYE+IzeONXF+Ts
+Jxe/4wTlI93fwGmM8QJyG/SpfVuhi6fbrCtf2Q1UTeuiDXq0Um3kwhjWi7x2Kiefc9TuYGKGxDu
eVCzSAy34ob7t4XdKhFz/arfGjRmL5nxhMXjUJ+nAFZ82Y4aO4KjL9gWop9As2Wibxi4cXdDcUdx
W+aCVTQqPHPxef1SI0ETZyfWdL2oGB0wH76zY9YhBgl0aIUcfCy9UsXBZrpcuzhxIO32DqYEJ7q8
4j+5F7jzqfy61qTJxFzBR/CwmXRvKeGsODyVn5h4nTQwLKPvuYEr4Ji8CbdVeGKRGJqhMLPMo7WM
xVnzaospZ4mFFlv2eTqPSwYX37Z6W42e6H7P9CQ+SEKsdJAKZlhoOsmtPggZTlqa1+4gSu+Zu90n
bc+hB3HnekOiYsmGSixPE0V+Ffesqom2yhOWdTaF1b2HbCIC2Prs9hO7OeOrTT0Akv8Ygu6XXEIk
at2OxDEz9/ZtmG3NCHaQjIxHLQt5ugAAUHymJok2J8vQkIWBeXYjvYmyXFhxKCvEUY9f1q992UTa
8SYSts9gztioEUCHg/Nv3l8hWNu5GfxWxBAKqo0Gp+fP36+sUN1S+3XyCTDZBFmXNEs33o9UrbU7
vB7vKLQFhHUnCJuYfgUgUv8bFl6o/gtkz2wScmmYhIIrM3mX/xd/qSghNLbHC75Itamkey6gTz6e
wtBtm2kCDojoEC3aymwz7LqS0gaHbG5EVgYtZyG526LBlwItd8w3WwwPQr9zNfLBuuShYA75TwGI
zHgTM9wnRvPyKYihJxyGddP9Th/ix2/uTTI7gbbSggfwxG8hwQ+Pp+BUFdNicuQD87rdS19zR3Ry
cF3Ye3O09UrVPIBPYca8Oq48A5Q62KOw4wdVAko3lDS0z9JRod+VtENCf/9chE3x82EgiSXKYujh
GUDde2L1/UrqcpYQptW5bWAQORtUD8NLLwqD9kSgXS5EuN/kmeV4g7O6PkTQeuVtpeylFneraml5
BU9LfTtDZqweNY1GLVWvG4mImO/c1a5yJsZdo2noQ0IweDz5gTEmheCw1hoKaQYNBvEsn9A3CDVa
hGApVdzPxUkAoWKY1ekO8fYDEUqyPuolk0ZUOviGZx43IMcbr0e7Im5Bh4TbalSY0C3xkTiwKlBk
5CEKTbR2e296LUiERfD4VLz+2ku37UtPJzDoxcuI1XQ2LjvqxHvTA3YBrGdQHWNBak6z69rSkljF
XIUn3IhDjM+sWtDE33EIt7AxdsOPj/FbznXrchJLDRVOraO9O3Ta3Q1vp+lYOQy0LHAN3MxcJ0UT
N3fSn3e2Z5ZZlvpEZyNXi488K+LbZTJipXJ57E7clg6i+M1N4bsQOq7cWJZv6WDm0MFWUc9Scyfo
B5qD/7RRGYxMisaC/aPI4NhOK6LBdJEafJVV/fgjUR6WAkFlU1NhK7KMbAo7iILnwgZedX2FSRG6
2yHQH7HmXo1g4AIGIpn/h++gtZJ5wby9/j+FMWVWMvnvXBwBHB7O/bf1QbrC/guz7mK4+zvhe1fl
EjxWxAwxo5wncNC4ceuW8p3GLNxcOd9PO/NQPfbiMDMsXuwJcsTBSjlj0dbL7kQ4oqjfbRMXJokQ
noWz1iGIz13VOpMvP924U1iDVe5/GR8a0tmU8RezloxVIntz4x93pkKFsKO2iv1+oklCqWVvO4iu
iuwTuFN/rA1b6qgSvyDitZZvNp6h+MsuqgP/id00m8qD+OatT9olmjj0PAdWn1ggzJ1Knc1BwAg0
1GnoaIdTqNmRPZeGrIxyeuOtQzCKGsbqfDwBeH4Jpy7CUa7NH4g6sShVWWX5EmpCn774s3LGbrJn
c/3DPcy3AiaYRjJXVMFI+dq/yxHfdmGYObQzhRAK/XdTS1u/EWeGI8E2eUZ9PCR/RnzYFG2Ux2mf
qKUNkg3SOE024vBBilrwih9zj/OoIF2WJ/vHHzmGT3gLHK/n+zGZLiuku7Qal/dqsqcP4pjktLDl
+MXdudI0MPJOnNguSzeoSaNS/xso8Aq/L1FojOb8fPXwTBa67lRQk71umiIUPO4tW6ctqcglyMjc
dCgyiYE9ekX1ohCfUluiTiTTBA48Pak4R9/e6cBbIfk9zT/0qyEMVOkW3dmwVTK5jQjbLOM7RJwc
ZAXwKCC9erqernu+yCEFi40rnuCxliwkrmsOorLuhxUath5lLQ4SUctk8Rqn/hiboEgXzzCVpdRC
1EpCcZEMV3gh1zzL35bK1ByMnjUHRqyeUjRqZQghzMxJWMRbG561/3nxYEMs5BR6QUqEWK1rNQKa
ufcvI+U02p1xY5AVq32WyEABR4VCeAhaH0BTU8F/lFBCgj8cKaI+9IJB66VNGd53b/5ksDWeODTA
ebUgTiULM8J5bGOiox0cXkpBFee/UXSFxToR5yXKcpArpKnO2GZ/G3kWtoBHjcjfdnSTbcyM8RA5
M+13J5nHPuXUgCpeUZQtiaNyGsSK91xf6v/5vrGEeVbUJvhYzS90Ueggx8YKA2S1omsCwTri5wuD
xBiYv4szwfZTT/bdzA+TO+qc5YiU/QgzyqYLvcrzNBoB5plV/S+3HEisv88V6xXpwujDa7/Zt/Tx
UofpRofJNGgfYj0veZOjI0yOq5AsyeQ8PUeYPCRBHBcnwxURoxyoGQqKs6U/f+6eqLBEvwVXPkba
B6c4qMEMEGXNOms5eI5jqwbxW/q/zzjB57tcit9uGzjXbDb6pjGq6Kwq5DMMAS6ANMIOhR60kwtT
+UUVx3xZyI9mIlroSP6Y9w8dj/t47iQP7skO6yca1fZCfD5u3MJxGqYqUPrrb/rD+i+TUUhSIEsz
uZ2/iHaBwcL7tp74+WFozqRLWN1JHjHMSa1Hc9pjsNp1VbodxBYgLX+MHsn9wPNz2ld50a5aSLkQ
OQBpwVeeL4hzIUScXNvgPjw5nXZGmzmaQKBgHsOVkYNzL1wGJpUAUuA4GF8BFZl5ynyU1X9JLV0x
fzg7BUmEUmXdk/uOTS6viAu7RxQMKd0HMee+PTW0SriYNIu+dPa63+wkN0C0T8iJwkrsMRNklx0F
JeYHceMO8wSYceZV69qWAhrKmTxZov6D2rZqGiGPJ81FgJVb64C5nJIqEXw8Ty4zuilUauNm9x7u
7ppK2TlqFdJowmaoe2bzFVx8DKgokyl5awamxdyKhst+1oGZQ62FuDD5DJxW1TPqBmlhaScwACjU
zUFJvnthNmcx/9ZRk7SUUOx1udOwiFuxfCQf+p7uR7/3H9SakYiUPjwCSMPdxYkQB+wOPPt+ne5J
xeOvMSiA6Tb+W/2MiLKUieH9ljEs9QMGN9F28bLkdXt3dIe5ezC7Mlgkz8K7f6LWsKY6r24HSySn
xpGddtOkc+8Ai/39Gj1A0pplCHSKkkU004yP5k3dTJKbK40fBurBy2v7rNBE0Z8Rn9knm6ebaNJa
aibuCBenGDRPD1HxTMrMcDeWmY+Ccf9nyfeAkGO3spoLntE95Bv13qY+erFhAy67hWFEyXOyr2c5
BYlzu7PhlG4uyu6GnvdRutuK43TtGiELV6N1RB1ICeINmCIYxsMYvYDvb/iasHR5Cc4/H9D1fTRB
teJwmqYkActXM3Zim554gHGz+8qeRzwCTP1MG/m0T1iOgjou6Hs57JKIUM2cDS7cnOEwi/qFpsd1
fkkK6RAGQVDmt+83w4lY4fpUWGmX/lfxYyhD0Sr4q7n5bs4X5hU12XreLcIjqiiG3h1HX3ZeUCdE
mAApK0WqYTitoU330nN3meYPaAVx7DwQpFoh6mi/BhIsmWddkJnbS/EhDkv1von5GR1F51gqaU96
GLqDdONMW90eLgVek0Dix8D7aw/N1t6lOsXpDqWVm4ksIfgCMddpPuxWdUZc5atIGypiYRgGY8ia
yU1WwLIljBuBqkCiv8v88cZ5C9pbnrNIDIaAdCWNHEAUGLVaZYtiSAiOy1rtZw0Mrz9W0W/yumAM
9eX6q6ay1ta/IPOdvdrCj23BPo2Znr5bwbN+7OAQ4QJd26A0ZxpccijIkYj6P989nXy3Eja6pEvo
TuN2gA5cIImeuWf0yZHAxaKx4yYK74qVGVFCnjBhuryro7lsDw08a1XVedmmuPmQuIrfGIkNo9Es
PF3HV9/N+c4mxMQq2P9pPuxQuNOfmpdl3s7Mwgr+b3uTCqEcXt7n21CExRYEcElbSSbXokBB/IEH
NoXYH9gMwbl7rogtCr6Z0cuIztIU+Z/K0DvYzqrDg2Xt+OBVoEPGUqLJGjGjok/nUjs7zU4cr2oF
EIE1QkJLYHJrBcErZsFIau//HrgS9M+4dvESq2qFckmGc4pXAKvaFllAQNO7EUq3+jwvRoksa/H6
iOamrJnmlrNmQVhaVcOBl0n9zBIaA1FB+ctDRVpCIhzk0OgNI9UB4bfPGE7gaxaEjfxIA+5GfZ3n
4q/VEoAtJGaf3p3VSa93SzxLsh6lZ2e8uygaw8XHu5oOPdX6wPsBCmCRD/Hl8VfpHeHM8Hf3KUGg
S2YCp/hk8Ui7LX6DYwXLXogchcLtycPhzix3ZIx2FWooTcWC7+3buK7eOLMnXmeaB/v/s/ObYc/M
dAD5uZ82uw/1ZriaYq+I9Pwx7vz50S2IsfOGDD9kQbOqxXQ10qPirzkPULLW/GGZAyChiGINF7L0
cVbXTs6esjHQ/OJOofG+SVsTDofyLYNHUxXXGe0wzN3DQ14zryNW9MyxiJjoCCaNuzLzjRoZQPav
5J3Obj/YYNw2a0XfLznsX8aTul40Tdt3f7WDVfAUvJaLAFsBblPP/tGx6UJZv47dBvooKwHsqasp
9OgVNcuHZ40Nupd6Ayf+yEbQlQEkIXUp7CFBPe6WI73vHp6V1nB4B0ZDnXCWxrBgZ9sqK9CBbCLu
lc3FqeTipUYQVgjY1wbvznU1JQILaHp0IVGa794tELI9CG1+fiIZqEn4+C10N9CODsmJuziK9lcT
7AU8OQAPjfNF5hBLzfKa3X7diLPo2v1YGV3x5XZELYHIIykqVpb4y2dJDkW4PQvtkCOl+4EBr/SN
mPAuIxpREd+dHKqxBZ5ail6XhZ1RxTgqZb39xFW/Oujp3OTDfBso9KjBMZ/iZOt65YIuEdltwIQ+
bPIf8csLPsm5UKpRSW18tMpdn1gIQB6DAc0Zvp5ItCrH3NcHRI6WJSY0CafG88xfwLZ5I2KPAAxS
WnBI7TU8Xf/v/8Jmw3CYAmCqMYucH1fJTUaZPhhrtyMswB4kmNx1dRbzzV39hhszmovTpjfG0AA9
hyDotUMVexTagkoIRoSfWgQ2Zm2ci48XO9RMb2WWli0om/JFp+G72Yb37afooo4/tQmC5ZxeeN0x
keZczqQFYhYAxyi4Nm7lT6SjMfb4uvHRDL3UA8NsJ7hcj8bw+xENgbIGV/jUyo1kI+ZTruO0zd6Z
LPALzyh9nAFKje9bGHu52fFc9aHoJFSTuD8ajScqTum9bmXlNYnqnmQT+c4ZTEIUi1Ow3q+POrSF
rcMEhYyomUoyz0VXDVIXellsAXx6Tg+p19FZkvpguw3nsj92F4Rs38OBN0PFFSdwpQheEA+PmKJl
XPki3sqhOGQDNdyeqk0NYRLdTE5nUrgv66YtNQqaNyRDhOPAUnjO6/mlny/kJXtZ0/aJ7rowtKsy
eKhegFkzopf1lrFMXVqW3NifnOcb13rbs8fc10BiiuLptcu2b+gKzyVAk+M0sQX3GKwi9W+ris1J
yF0j/w6LGRM0AF0Dbwwrjjuvc3V925cKgb39aGduWNvg/s6lKkfTMcxCuvWEiCk/GnTSCmcjhWud
GDp8G1la2+kMTqrbu4anPqfdG7RUFNAnoKBdwOrFpyOeLh1qA3uP+4+5qV4VTxB0+xXIJFYEyhEV
qwq7aPCeJGptqm43KB1U8ntZNB4VQE58XoteCZyRvPpX453EQPfI9Kh4RwkyCLxvnt5GqM3+bfO4
fXMtGh245pmiVvcr1r1UsKVXVvzl4P3IWL0dyEjlTJ1MbY/mkAG+aGre79cltb1H0Z/v3sk3sKVu
j7m2zTnA63rjHD7lRI+YXfWlQ7hsVXBo8FKhvSiwyM18nQME4e5O516RLXDxJS1lf34y8VYhkj0S
8YR/M8OnV9f+hBRACsXBJUub1P3fp+4Gq4ESdXe17G0DNnaYBpu6A3aDD/eoZHeSNMkPImTKymRa
uAd/l4Tt6ayKJgjz1Q5gqZ5J368YfjY8YRGdd5wCXHs1sPmM3WQqDXaail7Z3A0eBQsqO57umIdF
retWSylvJ1fouCxRfuYGnAJYq2eOE13CK4iH8mNpZw+JxdCZOKHRNjkMCHD6xOIdEt22w+SVy12i
Hp5QJtItTOkGYJURi39uOZPvwC4nOSIu0bLznJRx8GzNKBzemWi+rU8aBTljOktImS4/nZvQ1PBv
TTgnt9tgJkrKSuzv5UtrqmPaDKYu1rwrsE/yZuzmCct03Wqcnu3gT/XIYZK8J1YY5Fn/yWo7WgXw
OD7vfjEgkpB9bZRh3LrQe3OSoG6DGXmr/ZwCcsCB3EkfjEJmQP5yE3XgFRZVMUwUQjVVAUN8EhLF
99Phy/bjPJe3EdRNGQb70oNEgbIRhiQyqEwF12jJXxhT3ETdnUDftxKmo4LpVaDVBhWN3RWWfMc+
GFEcCklCNHEs0+PyWivTZWfr/kzOYIw5UgMcmhqMp9u29CU+8Hs/CgRveWanRE/I9L1opREiY74O
8cqztei5PeLHtasF3VGpMJjD+1bMZrqfb27mdZBMXys+kP8RhMC1Qg5CJsz79LUOgNLGLyngjwyk
8vl5OwhBEdvPcH9DOfeU60crpyY0HR1GiyP23+Dw1SHGcUy5GD8AZ14Lz5AB8AdMQfK9R8zDR2AG
nGxm6q6vL1rU2FyX5GvPG7WUfRH7WFRrrj+Zpf7iNHKyFsyXlhhHgghvOX03idC91o1nL2rumaXq
3V/GJUgfAGzLhy4OPcol1CTixVKX7bZU7VBfd7AYtpiDaVbNaUGl8U0+ElBZVFDN8kkD9SMfPCgQ
qparNJ7fMkcK2NLNuL2gdUTL1MXBWx++KVpg6T0MLzXMcnjkcnm/dFvvaSPy/X/lo4dcFNncYRYE
O9FTOuHY1ikLWZTM/Y5l/jMCjYbDZJ+BTCL/v9jvMFwyhTxMcaB/vyONd3X5al4u3OLwUJPdDgse
WOR799B3SiDA9hzI0W2PVJRysfrfwCjUF4cEil2AJbfXBeSrbmynfsTs+1GDC5YY/ssa/qoo8X00
h6+hsjYm6IKrjmQrOK9B2vGjrMEUiyxMVklPC7vyihgXnZPI62vPUJ59Cbm4W/wUuQVGapxxXOvg
7/mDPTs1sEyKc4NUfhL3wt4AzH4rx/l2l6gFV7Qjl4jC8qzw7aTRKyBmvzX+0I0Q5SYwcmDMxodb
M5m76X+tEdXj8kD/GNP8t/vJdZ4tz7iwOIOJRVdSPjZ9OkkKQHV0KqPJ95kDakxFVxjXGbuC90mH
o6FBDaMrsGDnq/ZkAxrPhtSSfN6aXNEPJuMvtB9SP1r2QASilENB0tXkp+OJjXQnnx+aBNvqBslY
7BEOPTcA8n4rBVCPS2KPgDaRfBMpXX+uyR+jcGTudHHDxflmaAWER270yYJ0CyZ0OgKSVhostyaw
Eu0SzP4oW3z+FOntlru7w2sPeFcmHsjgsJSHlHO2aGwtyb+tn1sJY6BJlAdZwheqKOJ46MIAj5UI
tajqAOb8kaPbLVDR6eYDIRAujK0bNhimY+jkfJGlIVVh7prEdIFd83auofB2uhUCyFBSuzKbKNJy
4vgwicmvTA2Uc6VQK8aEu1kreN4JdSYWaZgoRa4jcqK42vx19xcRG/wh+8FzaCyxu0q0KqHPg28q
U473tdxeeXc2Dk3h1anuWJhpDH3IoV0jfCbNLv5K5h2yXbz/s4a3eG9qUV1Dk3Vd6QDGZENLSCug
AyMCrKUQtaR4Y9M0bfDYh0AfL0XsKBoWNgwB8K4B2epxQJ+gi3F98lcfdHAB/hpH+DjjMXQQ+Vit
8uCCuhExbmAkTzOV2XzylZhjl7sF1Ber7pI+5o3XkIUnYhib4M4+DWubi8ZIidb3BQbuOBrpuKvR
KTIM9TnMjeINo0rLAmHJOgXHg+98SSXinRyxjlGwCdxSD7U8T9etD114EqI0x7yVdxxhu1GcAp0f
oPMbkW9M3afOOoIR5TgNYWU0iyKWixpM7UzXAjHk4s2BFK2woh44J86gNPNeWEFhwG8em+6lwT23
vD2+779qzbQReF/U0mjlhgMla2kZ//fWZFtNcXmBjcuiHn2zJIxSdjj4nFrU6bpgQIOOylqw+OTc
ZO7HNGZjoVXrOiIEtkYJUcv7OcbYOfjGcD6JZeOhG+2thd1uF8mNeGA42JHMyj+YZopA5n9eiHBB
sqicpzGPv3SjVtTdrUTGxtr9UUZmFuiIJBPobPH14tWOEH4ShZZJKCLcGMUe3/4nuzKmMTOv6UAj
rKuKxRIfrjLvOXuc79SX45LXjjN5auN3A1/3jzBGLqjlBf6nz7IUurW/0U9MdD2oEa/jw6e/1Qn5
6VYhTkhUM/WHtIZ+za818zdXfiLaChcvUbP9f8Xmycl9FXDaBCxcW4O7TcFOrEGliqWIrOCpa85i
J0DzP3YwQPPZa6xGeoITCs5oPLxoty97iyrF4L5sA9mAkDX6sBF8cMSmFodgX5rAkz3rOHnq7XHt
hoeMWc4cSqrHUBF8fgZ8PhojOKnJXyvgS+AUzD0hceAYcK58iyltaH6v1mwTq6qL24eK/sHWRC/N
+wDPtDGbQ/54Hcjf+9J8ZCric2ZXJcZFwPzqEOBu1O6sRXFinUtW9VQuHtgGUQgiJ0orfnLSVt7a
1brO3bv5phudVxpPgfQGyW9jgL84I2wpS891MPgTMBJoRzAalCpc7Q+k7PH12lRr/eMWMIVqtCHB
GOcgLlbOBt8R3YQmDkrhphG7TtF1+YTSYP2lMBH2k/XWBMsKYZcFHmyli3Cx4ZcTWrmyyKRDVX+X
2+tpxs/ELiDVvKSRQH3AHWp9KjpMJPav1yqvQ4dL/oRNBcJsVo5IhUKigEmPRwKRp6p73uXUz5Xn
lZohUktMP9bsMqX67k9G31gJ9jtiNNf9HAy2T6og3jIvvnaiNim+lPrjX96cgxAr1sgxBie9FPiA
pd9T1gf3pjqa2MyxnPYoVbvznkSLNmMwBSxi1JxkpfNqavttsZnQlPtrIFkuJuRj6HHStx+LF24T
vSrwYlHgUfDz+vpvlxcpeoEisjnt4COkT8jQ4/6bwninjkUgaqSdosSqeBdnw0ITWD/ajUq3rjds
jiD5HULmq0Zz7dHzmN7vX1k7HUIkEnkxqnWiA/JsaQitjYl9d9dNlG/ZgRXJ0MbSBowRfU8N+va8
/eN3pXjd8zXnCQAxOjOdgoE4Ex/Gtw7t9ivtvwGRhbKgjYrBTFZ+LLMhkJj817ovXcN8C+KpNkXr
2Aw6B/cUMsfMsjO85cg6JLj8gRj51QVXoDzzdebZpg0ohw7X33dPlpH9QFiwluLmfSQOFg9YknR6
YrNU+UHgMI8kOGegbuoil1CE/3USTxypa9DQexvcKPzp0QvxOJjL0N+f2ZeYVvaLVWLXQkW74gmW
/euKbnwQDVxDzSsINAMrqOFJNRnJ3tin9ncWmnFRp8Fs3sK18eKHoNahag1jV7SuO4Z//TUgQY5D
y7hTM1qb+Sa5FnmJwOhOzNjujuYKxf7+Z438A30P2GZ1kX51y7dcYCRpitxP3Y/RpomFMp7GqpzC
gu9tzxRu0cKcT9+BHxxT1YqImHKtBgGYfR2pjlwHcY1PAdgNs/1udyUhJxjljLbd/Cmt+gw0odoP
L1G+Yd0Ngb+TsLy0IEt8QZTk2Nrm85fB6r/gTu/w82TnAisM6SH3ZaLagkYFehWIKKDz7J8ZnzSj
W+/empDOchZdfRQ9ao2GHbBxzGjmG3LIKteK3o2+8AP5w0CgmSM9a7T927hDN0LK5YY6uYe6+Vfz
5fSdE2n2JGjvXIaUoiRXThm59vivnSyI60A4TlZj+3uOGjzVHmRDFCGCUQw1ctN6ikBrxYgzTr8z
f24+BVcrcgiZWvJO1EecIKGaArTJOfLLTMezOBDF4Q5V5xhsqWFZRojq3GJJdiA/p7dsWr+Dr3Tn
PB6vElFdCLbsEzV0Ptoq50RRSo6CrNWfQbfqUk06MrdBNRqEcogbzyc0gfejXBPWJDCS9Zs9e7uS
PmAYcZtMvrQQS6+HdzYin9G4Ysfg8SboUgpIXSrWomw1Kfm5gzsBGQjzTFu19hn0JyfAzwGOPG6g
iTEvNshCxmCZwKk1o3Z7h8rF1hy2/Jl4gFeEFQwP36zsj4x/xPrs/6TfB+e+ePqDbhF4OXPkX2mf
nlsr71BOAZ/DkdQWYtMcfvEsPRX9PQskc34gGkIAYoo+LvHThhIfmsPQ2kyOTIYR9Jf7aOP5Cmww
SB5Gu+EgSwLqPiknNDlYxA0mSxs5q1lOsTnYlO9q87UuAbvUJfX7qwZI59VrFHgQnCERqQ/0zTNL
zPhcg7DsxrAArRNgqOK+2HVA5DP48kMJ2/Cm3ItRQJfQbI2Q4Fex8eL2Tk89Ei8RYZ5+1v6Ug8D4
B3Xwkj2HT6/nN1xaWtMdDwmIZhC7DtI8hie6yv2m7eVWud0qu/uN8Ek5/S2pgaHCOcH2LdHaZFf1
wQiGbquomRJefaChBpqEj0TEicx7jKvs02mwx8AhGRZfLSpNeTix8UTS4Sf9j8NqdbnBfB/oCGvc
VpSHMMfkSpsXRnheX6iFjOYJ59HfVzHG53X9DBR0SLQoHrzYrOAPHZ/HWoJMcOODDBhFw6lBr3xj
pm4Q4TRhpy2CKK70+yn684pH4f/rKKbXkYkrKZprzxOLtcm225HpbkmfDVdBtssLra6auDvGf0RU
8zxN9UlHiYed3SnYEUmEW2fbxX55ZbF3Z8RtIPbQpTkaNomIFuNtCUrNmyPY04nSKIggg9HBpYW6
SolmOHEihNPzmOg+j8+u43H0JgRFaMyNYPYtuEnZ+XnhYkipkwVYeUmWoNcYiXaEuyixd3b2p0/D
Mu2XcmjcZHcbi91xTArhA+3D67/bZ0mx+6LSSlBAvZkZ7XuFnBf4pkcltE2XaMWwrjrE1pcYnSa/
HUEnVGk/QJxAwK/7K/VIJV+w/8j4IIyjoRfEiJyQQ83jqicuY81EBA8jb97O2QLs3w1QprL7i0R7
qnP70P2N2+/G5wXkY6EqXEBmQ39XnBRkWQeuei52xPPgrJRLbQdCtm4ImvJj6QIv2ttbWNct7VOU
euKJNHsBW0Zt0Zz38f8iv0r41TecuwJ0wQsNjL9T+u7BLS4VJfXjwtCuIWXd9GmxyJlglo530yWt
PNuVAQFobj4fBcCYByr1SFLaKMh1x234sEVfCmJR/+zlKRXPHJICuHCGg/F2QD1JzSXnl/Ti0HMd
q7tk/ECaFiI7vAvPpQjUdKA7+XsP2uOG8bNqIsT1aNbvK6RDEv1TCQ0CJ5PEBYG2+T8GJSdeh2e0
W6APez4E9APWzv/AUVyAmsoAtoW2ZDvEuO2Xi7nz3fZxicxaD5KYNdkr1JfGM5mKsWyaTRwIoFRb
eGXH8oTa0qbcczP5x0zV6qYhhhGgigMa1V/KF0Jmh2zoHkMHg7gm7UfVIE3pIcPXa5QnPFxwS6gg
69Xe4VTeLdx73zCpa99x2C/kEK7R4YgL+ikD+G7D+s69CSWemzIukeVGSqlaG2xOKH09v0D+lt7m
CMxfZeLxFdi61R2qxGVWlocFX+moKtqfa6FKed4Qca14ePQO+Xkkmc0X3I27ZstCENgPvU3L4Dw4
+zRAEXrezFFEcYEJLUMyxHPSk4s/5dmLHyQzKLYCkMBUTsgwA2QUeT08guSSoMcpyB3okF9TbgSb
PkoEewZKmmFj27irw8KAlocoFLip0bQ7Ygb7ZltSi7b8+pQQecFsr8RLUn961a2BAdM6K+WJ122T
d7lkUaaAr/UjXF4KghsJxFDweFxgqQ66W3qOpqVY0MB8GL5WgGj1NiVRSZhPW/yfuW3CbL5UOKBi
sfoULHUhb1yuDu+cEkpNhY7PTm3GWyIPn+WCgLOfHGmBzJgVnSWrsJfSiokVheSJ8FCS9yAyNVTl
9z7FLWbKlV+TIyM07x0DDhptIe9QYe4xxc28nDAtyYb4wT8BKlfGpyg5SJULfUTy9HQwEqCmRAXT
FwZ+SRBsrR08hEGY+77Ts9nuhnjhuktVHLobvguPRZKyByIfrZh+yZEvOIeDHx5jxfvesEvZUIm5
/tGyzZIRwcmt46SFFCxqXFljTA25M9G7J08soVeN8Q6URYcipR8c5cGolD+qaIMGy0zg8YS8Cuw8
owjGjjzH+s8SycDPuvHSfPja2j/yfkLTdMUZ0Cy8a9B9OQE6UY/N5x8kZJFVqqpisB4xb/kZCyJp
DlnN/VCi2BiNd2Ud/tgCuWb3GUlcRWn5NxfeXt2xNSnlBVDt1323fzBqTA9+np4doRGDqD1tMerk
569u6lZXXPMxVdOvXDhjRdjhf5uB5m9t2TtickHtvfMT6GK8jMscYNkEV9wTUOUBRD9bTKiBMep4
85M/fO78vi85Iafdsh3njzdu1fAZncwUGpfoTRTKUvnW6u1E1tJmvMqMcKSqxC1onpU6SIRrme5V
CoolychVyHzNvG7iIETHykZS+qgzCMBt5DcmrXTRtP4bqIocLTq7nkZqPN7ZlQ7SYpg9ql6h560v
R2dL9FCcacd7PCJQ5PTSl9sAO77hhnkLNdgZYUymQEn7IlufkdZ4lGPKJPB1JmlJEJ5H3RrZUOXj
oXd34zbclCN6idEfRiMlx8JEhGqdarPEFjHGAb5XUPrPRhaepsaPPWqyyVQuvAAzDkl4/ZCTeCV4
7RXeLdM8RQ8gA4puMfc5aFO4ED9VhQbFpASp3IY9L5U6jChQaa9vV5crtizlNHs+9ghov2gwvN2i
PyrLOaPOziaqyS1yx+oCZWhk7BAaYnS6HwsnmAHEGZqMOsEvX5eheYd+1s08KatYkhs96qf5hDaf
YjlJfgvehNfA86xK7MtvytT1D/BGNoUQslHSXWeR4LeBREOeeoYGCNbFMIU/aE90+j6AlntvtHU3
msj79tiW+oAbcNU5eiMHw1wm1Ifu1+Vj65yjFjcka1O1EIO3JzNy16yWPVd7LDeYZR+u+kBH666c
XVRbJgOJlgpFNfjaw/rJYt5WmFZbtg3Q0ikLAFdz/PS9V8ZlnsBvmQqLN0IO7wWrae0MgvCaMWRW
3j1BIW79M3XSOOQ1hptH5ZyTIEOtG867RwRMDsqlaMb1kkoJWGkfUK4hLKy+JJnUgNmkxWCsBGFA
Yls6xvgkJlzsZ+2rp2JN9csk3bMhWgPo82VSSH6BN3YzRxo6k/meM4KeJhA+DmC13VTB8KRUgIgV
SbJuj0TkSYsseMvB/kyhHMtoAo9oTOMTMkHrh4rCaVMWVQDpt03z94J61asOcY8qAaCtgAmzCsXG
L6OHZOxgFktbD0/SBloE079vSBkTK6lQsuHIIYUJb/HTM+oHXI8EcQhB/gS6Qjaeu5oZFi86Kt0h
533iw9W8NGrl8ozGEx/pQEN9+MP2OXI1dNjNaZWGN+wI/MGFiuGAJEEBwsXcTswJDhbMYyWFQRbF
wmomt/zFoyrb1VmqyORfPOLlzopkLStY1qGL27iYK79ommCT5ggjGdQbrTk6A24DaQvjro0soIYl
SkbABFgMB/r036XU3fo3Ow5F9MFZDnEdmBFIxcifECbD3tCNMyArv4k/kkFavOT6ABubk3qkH0Uc
DvcqXfjWeXONgg80VFjozjHITftic5AZ4rArVsrAsRYUCp9EMtLBzXdiQrt9nzptZZKNxei9scDO
UXrM9TjjeRFUOCTz8v1pZxbBDMIQANopz3R7RXwPQw/O/o4kSzbZrYLYZ7D5MVHlYf+VWBQzup7R
6t7nL0E72uu4r7g/KakzvGpqGPmwdIaimJD15GYaYkgGeXDjyoxwOXpL7xHGqikxmEujEdrecIae
FiJVdtHJd9vRxxP9VofpteA5N5rSrS7YgrRqYdlnuRdgw3nK/wrLYpFedY+Pl4+H56nyUCWeV85O
lF0hLxA9HmydYqRSMngX1xZnWWsouBp5jqj2HY8+BjmawwGA90mtKSGPWcJTssEYkC59yMlsuH9Z
MKArgEH/fYYvxiOXphD1bULyjYZR82pYqNyvcf9gZiaxCyG5RVmU+uQs0xIuo2MDUNBTRx5dYJZT
zhhtnmI8VukpSLllxQfq8dbjm+NNidU4m3qKQGNuv/VtE9QVWV8WWK0DUbYRnvcHXqkvKtmGPiJg
B+WwXQmdiwtHiXcBYkKsEI8tr2fG96ukL15VBk0+QCae3L60Iw47Rutkn5NyX8aYZQBCRpnxwHSa
3nSqEruE1qErnE3SNKtZPz1PVqKGaWvrzA1bApXd8vtwzcNkJmVeUj6odA6fAOxnxSE4g+Y7xA2Z
Lhjx1FS7nMIrP/YLpqAdIrWcTywsyTohHVBF5gdDMN9fgtidV3HNgx+CZl9jC39oq4YPGGaV24kl
Ud/rWsi3z48o9Axca3TDAo1Th84zKwMEgEIYQMGHDE2kngy3Co4bOAHM5w8wB5ElvGkLMNNlZYxY
Jf6Llp4LKwSuw5Tb87KpDC5LMuwBLt4fDOSkY6StwvmSkuVolfZovCS6Zj+5x8nhoIlsOSnanfKz
dDz9rbRxXJC5kcRKT955+4JTYIY1KzNnLI9JikFyKje20bTH5hIEyYaVvrCNgsnDoUPKqCZV8wvl
TbiSCJKOQPIi4j4WjtoxDs30ZHTilBd+bkm1m6QDbK31ebq32eXsltBeQoAjp09gHAJ5kOowhtpI
h54ce+l6B64jbmaSCYCGbuWYJrFLnHPTq8xafGzuqxmsdMmQ5/KEVAE50FlPlG64A6uHTDvnBly4
hV45fEerr36GVTRLASr9aDY9trKujdU5ab4Zc8YHva5Fx4nqtOExFKSpwajhYCTov5Ujgy9tXVQj
lx0KVH65t724GqKo5gbKPeNN/bVmcEdXrS2eKz53OWqKkWGDIV/pPUNzCzEzV9QwvkSk5y4giiFD
Mj+SMgf1ck/4+0WjbUJy7BMV8TdQSLoT/KLSEkz0/eYQsgDJQThdGRBdtjebz8eCEsT6PiKH2FcV
i1vuEFYHKaxlZxBnHFVdUuZpfpLk+8aVUFFTQ2QwaR8yDfjble+l75gei/CAVhATa9stwzuKvOC9
SMfjJjgtKKg4N9sRFJz/R+clHzYjBuytzotsUE1UZPs7vcJyXpyyjhkDy5MwLsF3Rj/xxoAUIdYl
/MeMn3JjPLk5Fyq88Er2+SP/pWlCJk3vWUOwQo77T2HW+1uFm4b8/myMLUOaJpEIb+UKjVL/Tnd1
eJ8Px8VEDGhMPyW7CakzodVTom764EZTddvNMcihRfZCNLw6/8FvkBvkecVAIWYxpx5zNtioUdyh
QasQ+0tmkaHDOLAF4/GMwOE1VT2kBMvCYBlR3GU3jKXe5Dox6lZ4073vQeuQy0tBTGfOUDTaJVv9
mhaeJR3rKAth7U3DRY/n4J+Ll1Slrfl/S3ie8k5To0x9nI/MoZyfSYUnFH89HAWE/vu4cs7zoyBF
f+ELLaqY/SXraZCx1c4LuYBsAmutmKSW2u1w+5zkcewcyTzybhulJvQ2oFIqWpnvzTcofgkrNLYX
Ai6lOw6HIRkuzjYBv2On7HRr44qfU1xqWAdIdkNneItrCre1aBslvO1YPKc6lsp6Mc/DmMWVhOy3
jKD9rl2KFOfAeq0vHyBXWWnP4fdQmr7RrMvgK6OesriqDXh2gDRRvDFPhKKapHRIoCrZT09Kus0B
ury45BUHDkFgT1LlJiyge/5WChWJegqpHAFNzWr9xha7cSmzH04lRi9OHO2IgyzvxHzVmbOzA3Z0
vP+5hLntyQjKihiHJOUdETAKjvqdF7BZ5p66yIue/hqPkFLsqbXxc8TzIv2oJPeL8QT9qd/MMfqW
W0KCshdsjM09zMz7d+ut8xjL6TE/0oHMTzygQlKB6XiRPt2XnYzSvYeC5LGBJIsXP6ChEDS1T6J+
/HlXubwevft5Brd+UqDiwT5vym365W+n998I3xhqyDjdVzjXLetyo7SEVK6Oc8ogjtXkpvNdVZun
SOCwdwAAlBFChB1TGg/qF4Z35jzH8mzD/VYlPHTauc4DymXDHfS+C1vLAoCzqQ/1daQ4zSFNopG0
TNhG0rdtgC/wf2VO49D5y+65gXDKqIf2HXgYfXTg1k+ZxSzMQTXos0XYirCA+hDNdVWqilY+BhIg
DWopp/qIgETtJZQ8ZtFmvv86FYgduu5B+BB4SwkeNtGy8CYggEnlaXojKdwMJwTqpXRZ5tUtP+w1
36VcBQ5vMAkWnTzmFmLpezMg21glfOoiUtj7TtGOPflUCYA+kZTW5VQ/mp2yoskH0fZcPpFwjG4A
KSjg7W55sUdnwfZ3Jbs6srOuTOp81TdVqXln2SwtbyindBYOoas2hzM/X0m/kGyOkCJWnd6bocUt
9vwfJlrE3fwFQpsVYeAM0yXi9LDEn7IWBD3JDWU+Mr1cxocu0aCmrumHP3ijcPF5N001j9HPZPNz
sdiyldL4DANKsJTpVr1BhUYUryTwfJEfsBuOqZcZ4eheWIro7jdnEVEgKC/rG/0rghkU3x2hHl/S
CKq+5SN7e2RmdALhDu9/m5tB+UlKg13Jj19yPmLDhIjMoR5gQnsbyMecpIws4v8Mk6ke64jjC0ir
Cr2sm2al47B5cs6bKYy2jx9FI9TIk9k85dyKgW0j+cWwhT6gBtifhZv7buZJFmVi7QNR89xUEbCJ
rWtROERl7oKIMNRUJUMTikauNsBu63maOcIHJVKF0oAM2f343sAqtqa3ka6gpleAxMKpFZ2w19wX
dXdhvhApMBjrI0zvchJ7sINgHesF09uctg+1Cu9431UkYq/ADU18yCh36isaUbeDHtaTchkcCrgR
OO69dZLq0wjrm0tweUVS0ISQ989kpK0GwpdA7LTX5aTfXtDNCzdXcNXLprxjF77bz5wKt+KPbTtG
bwKhVqW1J7AjYKBxqqzPY2Y4x1JlLJ/oBUOzYqyqEgjyDJW9gbbBwL1QbncEBsK7nZk8uL6zX143
hBtRMVXwsrRfChLz6Em6gqXdAlihonmHZosxcKJZcZShjA6k8ahLieJFbRuvfNBfJBmrNcZEbAom
INn9uRrV7t7aee9l0D2oHE9VjDwvA1hdrUN2+H8fAK0ao8jVlwlEvkc4QNqOfrAr41qni2gF/5j0
XVKh/5iYj+LSex6hGB0jLxAqThgmt6y2dI5Pi9HgR5nZF7Q+mtnwEL0rppPiBleMDVmDPQyoMpRz
5PS9UO5zdnIpHvQMwczQZZulSil15IG55BwF81K/F/nDh2rBO69lLd/o/JvVNq0mARi9S+MNwqgU
4wa+jPt98LJfJMPYvPVq/fRaMjnBAmtlNr34GyHVkJ6EWUkSlwt8I+ErmFERYPvJIX6NBjFbJ6Tt
A0kpYhwwiczL99CRlcCYbvej3DYJllDPZG8L726IKLf50SDEuSj2neUoxeYZm/SqpIlGJS+PUmbK
I0GII6N7is6GxwWQJqg/vDnBn7mDxOua9Be8akO145W2spTMtqlpm6VmcJXu82uEmmQ7+1fr/JmZ
P0AxXEo5U72MnfSQtLnxQURrVlw3vWU5BajkRsztmZowLn/aYcQMM2djfgxxx7iQki8up0upFIPe
9Qvm51TYWRQCK2Zl5SX7ts8khhIck7JTHBJHIj9I2fOioT8o1vhEpGIEVJH//+qVoEniIZul1Hds
X/2MHDdU5fiyZDIqb/DA725Q9Q+xXSjn1WKqcvU7jQn/fHt1bktgDh6px4Xs2XcF9OFsslap6+Et
HxWWGsSarDOfqiPKear60uDIGP9Q7baCthpvHkRkFgNsnsJCHRaem64Y8N4WPMV46zoPWBctrw/o
QHhQwweVJ+nqK3NMT7JmSJcE0u4IXpfgz3qbYIyAdgfR0FFji/PRQQISwQ3VTaFoPUeocaNZyWwz
IHk7XLSL0BwdK4VMSiSbj/KZyenZxXfy1pO6zQBqsB9nVmYZVUFvqNXqSS5TwTWF50aH8LWBE2lP
vHrkOyHCWx+ssRf1X9m+rPD56Mx2BeZfCyGwPBp4lQqgfKg3A/qgzmkQO09iNcH+AFrNuBMeNT9m
3P87oNnDJ8O9ymdvyfrUyA1yyTRmGezsHiA6E/JmYZD3qdRBRalCkGzNuhRguvtyLnN7VNRsZ9JR
svGznAGthQs7kum9bbll9I2T9X82KlwOqqlpnXamHmIPZLc0f7MPzI11p9cKOKNZp/Emc6k7qzSk
ei4eX6gN9Toh6EOp57GviIpSY4d+8QNk92bn1gseLwrSZB+3uawK2UtLfgEeuZAuxwXYxXQuF26+
MJV1Z2bWrxmlpcQuiRBheUYJwX8vxl0FertDcpDBVCTfHCRvlGyM3JjwX7JmZAhqcdR/NRpEcQ1u
w7mPhw5vIKo5kFWw6bBtT+VDK3KWOnBOstVBJziR5tuzyAX8KGkuXLS1C19sVpztsoXy678P3jua
miqtngQFWtgRdXDpEZZjIsZyTI41fjaHZtS+NpbWsd9E6r0Ehe1NMhZ/2/zfoBhxxg8DEQ1RoVa8
RNtqhri6hGE6BYIaHHHmaLWJoYXU7TNgPBYw6CXJbiLH/xKH/4ShpI4PqapZ7eAA3yVGdw+y6Vfj
sfMdX4DK7gS9eahMcRQfjTwVlZ8buuH7gr2DHuYteji5+8DC39O2dtjPhAHsbH8BphMJiuXtTKir
T9tHj7KvQ41dmZprVkHtIhAEAJN9a9GwDZGk1nni6qrKnygh5n+I3tcpHe7LeDVCWqBYnEPaYbzk
t0CemIyyaqYKj/ZtaNdrU6ugrzWsp4q9yP2rTAUUzxsjBlywBbpcOh1K3vUH49wn79h9NnK9eyO4
sPzUP8xMLFgdwc3aBtv8C2PLwBNs66HH1UOP14OxXTszIBDNOulO0XD8zp7lenIlHbAFCLyAZga3
JytSnnlsMLx9Wm/vrStD/vB/WmpyFcbCYksKU/pRM0sWRkSzBkCF8BxAmQhEaM2MGgg3RKgXoc+y
9TXaUhppqHvWs6uvzNmtcKIRMzyayM9oq5TOlxRwGh9WOY41t3uMNzueyOysE6EjMM8Q/1OXYF0J
rvHmdEO25xpY1vGZwWGO2ARcJPqMHYNBwEgw+i659UNDNSnDYx6Xk3xQzIfCFh780A/4MwX6SU3P
rXsAMty7HL9JfInm+Resn6Qgrjvp5I2SjkW6k0QFUDkG277rjUQoUri7Q8y+DL+SAw8CzlSvglXb
AAWqtj4GOLtEND7u+l+dhDIMzm+xzEgO3N2VNiwJX8LiQ6jVRWsoxgdZUyHsTk4sqA45iqPi/M0w
TmaPfKudhfEcaM9slKnSHlYTEtFusZkFIclm+UaLwmJjpplV/zDiDXeLijnA4Pwb2Pm/nlHNr8WF
EwHIR+AbAJULbJyB5HOFl+YPbLaq6BoUnYCpayDMdRZAS/8k5r/MLOoZmtTI0HdVigt9DHurfIYB
evL/hxMEYXK8e4NoLpzdFm8zZTEIcJj/fBWm61tXCWynzk6YpJ5mtTbkl1g1ZGZLgYX07glm4KUH
2Vk6oZvsDi5UFUzB+rg1mi7PZdHUwtGxz89nYN3v+SZmQr5OpcuSVOAjcF0BIWFEcK2o0YqBt3AV
VB47woswMOgWzpbGUHFqvWpuatZf4+mmJXRFgQx4deyRSmrrsclVA57KtPITaXI1hafOd9c+4pvw
N0nSSM1It/Lp884GqrXHyxCu+SQjIgNp0b6ckxqfzLJzr03j+bYeUJKGwnP2bvboaLQm4aJkvuse
De1hoC5e1fxAU9f3swizz9aHGXoEmBpU7AAScEYItBYa9HgIgTKUoKGKt8EpDJXc4k5fNP2Y5ovN
q3lqVprLYkNzI/vTbUzPgZIl4Jxu+d1HYOJpwbakzlnsel6KgVLtKl/qAO8pck+EK+q6QkFn+OM0
sr9+gPPhu5iS8aYNMVwmJKVkA7p+QUboiqyhre3EhQHyk0iUqlRs2XhC1rtYICmuuSFv3MtcXObm
Dpe2s2VQKdmgAmPtCv0UNunB9KUy0nxh02mjhthRwNNBWCNlJbALay9r4d0cjnaNsNf2yWe4FOxC
/Goqh5vzG70XnU/yIiaxuCrcdn4jycQmBYI1x8PGe08n66EGOqwoQhsyXkj7vhklYYKpLUKlrf0U
4t3qqFJtdDVS3WXn3iNBKq+duApAczxlgj0TcCb11I6mz+jN4D/CsnxLpgQNU5nL+O5Oohvdb2y3
ciDirbRiZFhT40LjoYpeLWJ/at6uZrz9C5Ag4jLjaJNiKqwEMUc3zqWkZcsg13790qo8zZa42wK9
vWKqvEiipPXlgkDHGLJ7/5Ol1Ev20aSLuuscYoJEwjrMgFRoGQCRzCZvn5cxfQwN5qhn2swWFqdu
CfBhTrPfbKomH97E+vzMd6ommfkHx0r12IJCtiIcXuSVDMQiosXEWCwwBoFZciuKWtAvdiMIufRe
/zLrenfCrpDpaB1sG5KAnMMona92QDum5ZHjpatWT0UjFabcihfgT0w1ivMUBqxHLz+NHIqq/ZFo
AFQGueiN7/3muRUWtgaPIDfcBVEJsTkbrYLjpM+XJgyIqtCRdntF6KMrdZ0I0NUzar/L9+VK6W+P
pfGurAzE83Boh7snlezyAqXSv6yanmAVSD+hrdPfPqtDUK5eXywYezvcWg2A7rUZ6CHClISHFd1k
ExRH0JtLScVWG0rh15tvCQ+MHZ1Qg+LApinCKCuxf84ezycQwLFjGp80Rou8uDNQWriqBc7gRXfV
OKRFHzYAalkrwGl416aU7JGYwiyjccrnmpjrylhZJYbmAibt4derOtfdZQIR9QMoVUYGf6HGbhhc
1CdU0wEyvU002qFw79+0zh+ghjrwWsiHOYTtwk8xUVAFNHNLK5mKBTtqFc4oW+PuTVisMgsunJ4c
/6JVYTVihttqTC7HOWcLGCr1kDl/qmOmAD+W8x1Ey7jSylzdVKYCbkQqd1nqhnKuJdcxxjUZH7DS
cwqWpZM2gFpdaArlfjkhF4fiYULeLj9tW0awZFxJqyCJn3gwvimrUCYxfW1kOBWgC4E8A5VRECJj
LC+jcKrkutZXfCZzrM1r9xAFj8xWawn/rZvLSddDL1cJ2ERiI9OVJBuOQvtI5UnopZC32EjqpFWK
3rNkQoWTq6AHwGsMNlEsUvQMkyaS/AaGlxo4TaLIwk2HhlBGFgWNpCWPo3UBQLifXszuzfIshQi9
fvvGlQmIJ3ubceCrtCUyHCtf6qSrn3lAzX4ilYNkjnhFV2QbFAQwdP2qqpgnjMVmMN0uN1wLfnrt
7pCI6XZRoFoZf8KXQy1lIuM7Xsrg94LhlrJgnIW9cEdQ1G9U1JGfN5BsmI2JIK3plvAorUVJhwuP
QnMKb83PWfqZRQ9KVtvwBWRnLx04XB6lest41AdrWg2kjOqsqhoMNL3oK5Q9iIjX9qYVVXItJtQG
72JRwIAyw/EI7rkF9UPitnhaR5L4OxrrNJpxrTOXjTsskC6p9COuBlWAvInj1IVqtWqGgIzXaK7K
26LLzjgLTwGttiSUcVBWsAdgGmpsm13vuCcXokMqfWjzG+VIiTk5VRyW+WeDaFfdYJ8BA7nzgLkx
PMCX15aHk8IgSXlUxsrAwUKsBrv1Lc7d2Y5QFMET1B4Oad85jZki0LbIQNfMHcyr24Syx1w86aAh
Qfrglv+clfulAT3YkgDguHXtAPBU6X+bOPgqvPjB67GK5lKIiiMV+nAtO0ZhyUtGcT5g1gGy/iex
WX43Dvu8SB99IZ9DtX2+ThM6LxE9wIHPx1/3CZpEGWJXCNqOdpRFZFVrmbc4BVuuQJs4/mzf1O/s
G3y+h+jT1fFTP5orEaXMGxQLsViakmnP7OfuWLAV5Gc+901zO0QjFgKEEnAOLm8uWfBlweYz2GB6
g3vnguNU2hGLBqnrSZYh8dNTUkedMmxdu96fAb8Sw5DiOeJFWKoAuCK1XLySexo0sIj903YEpjbK
TUdHVh1AK9CDN4SXNXNjHbPt/n2GLaLzwPU/vp5RDtcKtvKS3AFjh5KT3gDt8CZV2im/FDdvRPim
fJz3+tFfXopEBPNB6x8xgVEDHtEYmWugv9teAWBfK5Zw86j/HEGRODWJhg1ODxKprmipFlLtBsvd
3iGrzh6EIKFQisd5ch1T4fm69jx68NOr60n/nHvSCciltcDU2fFzCPRPCjDhRD8fy1W0OGrnAdVN
vsg0YiWXTTWCmZJtgz0TDZ5tj6PfCbfcXpNiOwtjEdLh+FG28u4Ae6tKGn2Fp2pqt722E2SopfSJ
FuK+maeZelawxM++6ThWTFbAtiVAQDREKX369v4Foy6z6tUOvua3lU32FQzecqNPt5ksDwGhKJah
YvL7bK4dvhEIKhGWqpRG454yjCQYZfmAqB6RQz9iIIT3yJKvq18qpm4mhkGxlRhMxFQEtFqXqsqX
P68l7XHKNIxjkwAKp6P/zZfGd6+SjpP7BWcfpvWGW0EkCy0kelzDfA3MGp4dYLQX0IODj9K92Jpt
2ewRB3/c2uYTDjeePGZwn1KQFcPZbDHgCpoHwl1rrRI/m/dxXGau+sGEtagZ5xb5ER5xFajncJA6
mZZp68RBxR4bLsOG69j5Fh1GwpSlmoXeXf9lcrDSXV9pya40B0I+6jNlrGzKzQbWx818tyJf9q4y
lPdTPbo/TKn9elukniCk8leQnBTDHXMHl8Vt3f7p2Q8nq+nUlzRKd+ZtxHE7R6JJRGqrlMV+XZhr
bys5GHdYmcU8SOOGrg7my3Bh7oFmknGSKOX0fCSVzUsuGwOga5+iBu8CfEcWzdeEkEYaMKdj8/+g
S3Ioq9+ToY2IPzQuAV8MB0qwaN22algaw+Qoh3n0bGNy2F3zOCs781fewgAvmjxNEi85PT21l1g3
T5qNhuX+/HTO6UomArdoPb+5zWDTSpjCAyYf/+1F7QQCVf8fHRH8tDdfEpHQluAE5WhEnrESqz/d
A8pcA18LihNMShi7enPC3ZFrmBPQBSfYFGHTNbUZx+uEG2ddPFsY0X1qUwSJSrwU31krp9TT/OBi
sCU+/VD+0T+0yG0xSZ4JfyKPdUm9MXIYLctXiB7phWOQFglMRlIZe/N1zS2ybIEAzkOIscfNf+eF
96rxdmNoiTdMbIhxOEquFd/3SIIg0kb2vKAx4rdGDUg15nZu2kfKcpjIN1dkM1RsN7Cj13i+TKHc
ovp4dFgYJHCfeh/Igev8vP4aiw4CA8tTCJFnqSjPU6goR8xsMUkS99DiHD/qSMclCUp5rojPXdev
mLOzbjTlB4PPiNy++idqRmAUsh4U9Cjh/9U73axc0yOlOjUbM6pLA8BJAO+Zh8frfBUTjhBTIo6J
fV3SQjWhhuvHsqGkjDf2NWC3q3W/n68Jt/0qCcppTWTaHBzJUVY23S8jamCt80zGo3EGWHQY3UnV
d2VzDGWGHqAYjf77El0CpagGc7OA9mZ3hJgfmHb8qhuP0e6WRxBG6vKj5bt9HAg1ZsiJC2hL9nig
ob3EYpnIKas/sShlckZGzPS1tGmsDEReG8Jcc4fGFLkf2VwZ03vjBa4qaxbN1ZJbOz7D2jPbHB2y
3KRnH1a0GVq1PeS3jwzYw2zjrOE4Tl4EPobVKpFKujpGSqASexzUGRtuK9bmoPyr+fKOVuMU8dmd
bvtPXtvy1uG9EshraEZGSKx1Lebgd0KWtpKjn5WpsyRna88qNkH5RGDiruxTeBVGEgV/GAoguBQZ
VtI+sNkEBDHVRvGY83h4Mv4/XJ4U4NrS0V0Q0L33Fe8LbVYyE+snBeCbmdpkD1MJEx1MhV9Pmkun
HVnf5FRKr7hSf+UqNCHGEbT+DfTd1DBFUmSDUIcSWR0XciERj6ks7avr63qp1oFQt4Z7PyF7+QtB
bgt6UdZPRpqvCxRUVRxjN94EZbQBP2lHuaJN+HqUi9xKTrn3r6cgP23Tnxo5azquTJf6efX6OOOg
c0+F+NL3JVo3tR45SMOgAFXG5AVTNFEGB827WPEPdttW6R0qopvrM4h8HcGZ4ZnBDjVr/B9R3eqx
QNmFywULNnYiNQNJrQvoSTAS67cz5ioHSz0olOZw+9bXdZt4ITdKMkzO8GXeTshb0tERBAK3SSaY
2G5HvoS0szQHbH1PqwTy2vRadtv5TwgOrIq7msWWjj10OlBSI0vxj4VuC4XS+/Nm4UQ94SJXqVFu
6tXs2joajZ4/nHQDO1AN00cDeZ2Io4Z1VLyckh+K6ddTslUQTU3Ii3uWuGf5yU07/J2Rr81kbmFC
1XFn3MCvJHHXFwSMWIhuLoCuxeztcf8UPIdvx7pqAbTtefySduILXd5UbwLGrvTIBMRaW6cteOPc
DkKPb5OI8G9IaTWXf90iNiRSjQmJoyYjV2AHiz5cvvBhiHiVe0FiL3v88hqV9GAP+CMIOASXoKdD
uyImXjdl4PS6l80CQcBxSpOdE8//3xPsP+bdwGta3P4O2X2e9YQ7tnPVfn+2WurlExNWQpm1lglw
93zUTsQL5PcTOG6EZtrAdzrqe113QJQK8exLhoaXkG1sVTHRtdTLeWYsQfkkS0/mrODypBROb/Qt
T5WNkQGGu7jZ9feBrAkFBxaTeVkojKOxp5TdbZz1Lu5y16PQz7tyu7AO2gkJbNKEZL6sg2gpjUlU
nzYCytX8Ai65JxiG3dBHSm6mjzY0Z4I/0d2B5l16yddmVsP2XM4K51NnAzUxceRxITvMuprScc6J
F4hkXWqMk6riB/PeQ3FV8oFp+PEr8vwPYlW7X9TvNgIp1ECLoXiUALEFwQn3EcaFCAUIehZnnNP9
oiKxU6gCM3VnvEVLg60uYEXre0FfpfvXLWp6wRd6ufouWwCdA87uZ+IGuaAatMTdc8jQpazdLEmK
jR96FbMqpiaQLu24v+puBWplvxpHxE3fQNwXTQMiJwIJ3EaM2bJWOYGQa9AMDmlK+g1mMCjlMdDr
Xtj+f6NSrcr07dzaQSHoQHzJ8To2VIrRwLwFOooEZ/FntR80fwXxotYXkdMu9H0RC0D8huZT5djL
e1ngJZr7ED0tXRv5T4yEjaavVVcL6LgsogfVE+wMelbni8SYfh631A4pJ6UO/3j1XxttbT81bQBW
p1SLpG6a1MfbDUmcJxT9GVIG5wU6CQMYKXuQ7TiMZWPTpY/j5Iww7OMAUXucmI/Z9ugLSCN74j/P
wStN+vMDbLG+Lc6YACjq5g/fTyKaNe8U1J45s1AaQXCVXpVXILdhH+YXO50vyODFhXIJG5LYwLC+
b6hZrl8DBFRva2VKRw6s3LFYR3zDLA0fS43L9Lbiv5k0gzZ0xZ1g4AYiitkbNOS/CWd4TCVIXcpL
70jqg0Yd+Yyc70zHlA4rps/9QaaPYZKvkeLDXWc0acTR1RMul+UxY9C83ZgkW3WH7iFmOCaTpYzn
2vXEa04wSpgbNi50uUDdRW6EkYz/Nnwp/yfK6/E/Ux2/QItliiAyBTgPGb7vKkGh3J3GFR7lmsTk
9Wc18Xf0Ng+5R0k/tgqz7hYufAeLtXuKUanFbR540ZzIhyQWOCaiDmmDrMA4GfUmynzGMuwgDMAt
CRObHNh0asHTJzar+Xz4AKMDRKHKgRaxRpBVlRq8jPIVYn4DoYshr0xlT05zpEUTLwzKmZ5vC6Hu
sOWpiDDJ/kh/lYsNuv9BBLMLfYAv9+MLLhr84U6zuJpmLlcPMnoYKNSTlQ7JT+sPmuTN6JulEdBy
sV3IBWaof2DIljwClVBeO+J6xBVoRI8+1yCwxfY/HmbnmcoGdnfvJ0/+i5F17/gbgpxIOmqvgOuN
gcIgw61axtqwbIYiCDLEYxrqsuBf6w3mhknnPWD1rSdURK9SgnMZcO6RG0YcENh8GiT01sKli9EO
FSuypqoorGsTjjTwGaRQjzXu0Kq+NUXWe/22uBkmwf+5oPa2vFhK7LDUM1hAArzHGCCc4QbICMLo
uTy+d1yfwEHSk4ebnhxMA+b16KjxW6GhnQOXAXUIlxx9E0eXGiIlr723PBWxoSmseVYtZN9CzQme
uTZ9CCmYxQNkn9vtY5wbQgwwcCWMOF4wG4okVzMzFFnHDX96ILQrO6iVAEBSlKkNLWHknqXQP7fR
x69THpJD1sBU5x6YYqcJ/dCD+sPGNdDACxs4t5ZwCJMK9uElrR2QnTlbObvskqBOgeHhDhRCZmMk
HUeJmeptT4RcvfRnDIdUHjwBltu9TSY2ahrF6bBGzKYP3/91uLYKNfuzTFcg6Q3XIqKlJR4cvG0O
FPVdhLu4IIqiqGG9X7zgwbHDUiCI8gd0jR0x1Rsy0ITSrqxE8+JOFu4sexpxsKHtI1HILK7O0cLG
Uafhqsd3rugvIYP9sI8Qp58AFTNWIpd0IqnumjQ7FFOPBJ/KK0N/GLd/yOtL0qdKDxSrXspy9nlN
YCpDzsLhX7dTSRYK294773IvBPMP5HGGvCudctoHaNbTbl+RsPha5YEk46ChrNrvMQ379I3udrXx
yobR4iVq9ll+/1KvAwa7cpYwW/d7h/R5dmIE03qkLDwERk5W28YU1irAK63loS5J/7etl+JCDZRE
kMMpamRdREWImYfIi3kIedKLkSIlaKcHkRG1QdGwoA6Gnd2+MBnUJpPOxPFg4acVX7WIh3ajepLN
eyt1VVgIEXd4CQbrrvZd6pUn5yIAgyUMR2RXEVs658piIBWgaurm/07egBiBIXfRDxSKFGo35mIW
SEjku2f15MCeQIg+wFrdV5SJLk5NQXVXzHUR5ibwxYLWHGfBWH/Q0VsvTXzt9UpDSAGJ94KkO1dV
sRVpm5L+kkbnciiepi5KMw4G8sEjlCKLa4IEFcO1Ezio4zsw2Rjq0mawqbrfLd+iXnxu4k3h3bV2
Xn6lZnWyr4dagpiE3UqDuqcS2h69sBazAct+sWKC3+LIkX938wsKBJdbIjUxz5MTUwtPseELjQ6J
zgmk978GCd4ETxr0QiaMpMzy74dLUeDKVVjD4Kx490f2Ac3ZVRTHkCKTrskaRGUPgIyA9C1UCank
CX8a2d/2QL/dNUd0Q3YYK0iABbU78Z10rwcBzcYV8k7gCOX7vXr0JMQRtt3HL9oHWVZRAod5yC6y
Axlh2v66JAFDL6I7/5mPBCmCZPGVEhLvbyubq0OAmnuBf7KyArEEP8/8IA6iycR9++TYdfghQEm0
4hMKmtaRPMkEGcwtgohgRhufFS21cf2cAaIL7LOlYU/9KpAAeNHfzz1s2L/hAWSpv+C9UlH93XST
F4U2Bx6sJL/e+kXwedPVjMKwbbJNFh2SxhiUkSsQWp4sNSu/AR6pOikv0IhM0cP2vFUtXm12TEZm
eROAs+48mMKff7FKQxX34h3UM97Sjs85zupqO93hI1JenlwT5g3aHEzEYRVolPxwVwgu3NX5T4YY
LYAWhHVnnNXMLA280IYw/46l4XejNe9hVV4plbXDx9uo0PJPjEyE2v3unSIzmKB9Xa84u+n4jXSA
Mq0Nr8a62cxPLiaMxUkIeM8ilMjo1g+FDth655pUqawUJatwmKtsdPIvwZuNGjGs215aX+QIb6kA
QuE39/LhKyfHSixFcVV7wTJfoX9UBqTsNCEUdAwAS9wP1nQjLaAqt0YMmy75od6DUP5s2Go15fWn
/DdxVaW5tEw2+/fyNHG+gwrIsjZuxwkLxEYrqQZzkM+0xqXwA6Lgx+J+hGvG0Xp6LA7i/tjXV/yU
4xjiLlIA80XFlmzVGtPQzg8gLr2MeN0Jh0mj3SHmc75oeRmjIRJlmnbWqwejvJU0Z7LZ8aJICZLb
H+C9uOXosyNDwEl17K//Ave7Vrs69nsddYGnm0LD+EexYEdxUJ7tuj2TnvXVT670S/6kQo95XUbP
j1xJxY5R7l6ppPfnqWc9nLmIhW+kcFmDvAHbxaJhn9IJ0bpGS1NvYtXQXlpTYwI062ulReAE52xs
lIl0in2CLUkR8qUEk51fUI5JiTw+T+VsKygz4tTjSgRA/BHg3Da7ZFhGHEN7b0vEHYf00dB77KO5
/apsPM2v0E2/zEP5IWfT98MwDWJBAXrsRC/OF3V+UoAXLqkjG+mFyvefBEeGz81OKO7lmC233Q+L
OnLeEe7E6zyMY2UVy8GD9uicQZgl1wtbOe6fkv/FYVA75icMEq+c1lI/YGobkQuCStFAyMLGs/+l
XLwJBmOIf2jI9Eugu8V8BB+zV7bda+Dc3B3PMzoODdBOalNLbMqq8tlaBO6w7PBp+ewGb6CqgY0T
IKs1Yt0vpl5gOXPsOUDiNGKd29Kh+v9wF024NcQR2sa6jkXFnQEwT+IW3X+IwZckIyUEUK8/k0et
16rQkHQ1/DEcl0e5oSWu+5dN9PV7pasiQrfin2noXCdQUu0kNECmV1s6aTpXVtF57AVdt33nmJ7g
5pOy7OXd7wOAesfJzWHV50KOcUfZ+TacDI4Uu9v8Mk9KbjWWK1msCwUNSikPmfZeBWs1cSpE68gm
1FG0u37xj3fIhiuY1G/v2ECdXGWMTmgHGQfVGXZMxvP0n5ia2LU1m786sbYSycr8UnVYe83w180X
ldUmD27+aqvOurfwojcbLRDwyVhXATcyaac1Do8aaovtEeSvkQDYhXaqcgV7rnjSNSKWD2XzwjOZ
0qOoUVkYZIlVOxHEci+S3DB18OXhnLsMrwfyXQdZaChLxePC7xLZSzANAeDJr2PolDbL30XpS/ko
tdYia/9jWqYa9axDyCZ6Fyv3VbgZ4soSD9iIZvU/b+tZaC4zCpYTRhhEclCHL0CYooNt3scKVJAF
MbECmOuIKmMzxyMq6Xr/Lwg7nLoPwtAUf2DZjfO+AYAB8c++ub4oJ6lWleMvvKnr+9yHv9rKrchy
1Eh0NCAKHOe6AcEKmmS3cKyS7ilkgwrYAoZ4Yu7G4bY/tZlL881wGV4zaKYsT8Y08CA+/ydk7TUa
ufOz7rNTbU4UDjtMpro+TB+ODyI8SaD1RZRLWm/PnFOFbhPc3kJ9313y0ZGqb5la1drfsF4smR2L
Ut8qMdt3z2EtnJlJt4J+FkkvG70Q7m9KHTyvFsskZG+Z7sTb2tdif3GJGGDeN/DEIMICGFQXBOrI
4uNz1ui62euRvq/XV6gwQ0zfm2IpMBqQLlMP+QUFRZhFtIDbwxXXOEnRxJw6oS5H7gxH8c4wOcGd
LObixUA9c4DjyZAO+yxeL8dSZOyOkqMfj5LtiufhO1JgGGX4aqwFCO/zK/lBiEfPGApv4exncHMK
4OHH/2ILk5xcwVA5KQabjX6rkPfH3DSzGH+bXH1k5UMaSLQSIxlmdUlElkVGD4wYkEqaLG62xJcF
B8jjougX7WrIFEGGUlV2cc+GD3hR0jM4mZOz8spB9GmSrOm6nK2lPHYdBT1LqBcjTm2ZMs1c/3lF
mzQ9Ft4fFTLQXj1HSFMnCUWWzEr+rNCZ3mWp408Y2IRrkuqvkthFnkGx+LHWv6eKUIwpcbnmQKzg
kwfEHooGFyMqnX0TuUsNJ85DD1te8n9MD3EimMy7mZYQIHjSE4mmDrs75QQGkodtRNjj1m6MKiGq
wNATZGTopB/wtF8Rg6guWfW5bYfVWeWshkgSf483b8kV58Nbq+g7ppG8xoNIOEbAdaCOYpdNO+XF
0wmopL0NmGMREzH9OYGoNTJrFiAOo4R/g0Z5NOYCJV3RvquizSHTF+JpmyAIXkukSyVbxU4EAbz9
UZcT6UD152H/7UpmiLgQhiAUCRoL+BIBhLPZjw+Y1//8H9lH+sZ6l/QtETJbFeaA423hwrKXCSLr
oqbS2XcuYPyXynGDdxPPIPLztFtGxfUwHMCdK5J2RO6GQkVXBhqMn8g0DVG/9bDd8FvllrOYsq/G
SS/riRQyo/n35zg8mXStA22BiTL1nU1sjl0WTGrmMHB/armd8ocixKSInmpIIKmWht2/BcaD9LXu
EnByM0YBB71Pvc7xiKf/zRtgFPTQdHeSXqqGBP9kJyhjOlTabqqrn+AR9YNNzjnYTrZqplp/7LYI
UgLCxUxEdLL4ZHoeW3WJSzul7VdmJhjsIadwC8eyA+KP2w76cSv0qiqZMmJ3RiCd9YwXFeZyfHKL
L2STtkWXmEO8CsCdFKe7Vxw0uNOoy7ryOEDW207AK5oI32M8u3yPKEiH2Ab0jB80t/JfpeLVgwWo
OZqJVuKvuPdKwbN49A8EDtbO5ssbqnwUOcd1lTeGLTB3TDxlyfiaK8HqXG0dFu2Pbb3SijbHNXq4
6309TPi+v80VUfcJvkUl9ChxRFh7Rz0bTMkr7AslmGZMlSS629xVVizPvyIjLvuQk+OKTd8WyowP
W8fpSb0ogx+4XccloHwsSOR7n8dxtYxgKRRCPMf31a+UYoFsd8M+UaeOJO5tToBnd2xTpMKZb9l+
OIMBDmxwKUPKcXwbn370VueP+GMr/3xpZrtkPCEfQf7khd29TGJl6YWjRTyjYC2txc01OTSJryGd
bFJmEVKYCTMzT8E6mqgKrZiA0aTQrI5QjtCIc4p0Ogc8mu+X/Tzy2xN6fthwgcqZJyMWZcvK6MRZ
aIWdYD1YZ2ejp8yEwdNSilg0DwSiKoMAWm2qeeS7e8zlS3gR0CYHJsz6k588p6pCRsg8JUwnoJQA
/boXxSJaO9nTP3VgVR0KEu2hTeQTiIw+Hhf5VG1ylll3LtmbwDG34XQ5RM55qUUaWeT7fzkbrJKx
1y9HnETmovfN//w4D1fpODfQ7khmKtxSb1NW+UI0goHk3/LnU4O5hndi5S4MHq//1g0ehrVEyKXd
rsu0yF0jcJEgpEEAH+qCJXcOtLPCeopc89sBmHMuPQwt33JytY4VNXFzKMu6+Hi7ck/8iC5g/mEW
w60xCpBbkhCAGqiBx8ScIuttNA99mOk/rwZm462g1diAZOgod1H6DUl01fOtVafZ8qREyi6d8NLw
9dysPSpwsejvHIwU0GNRB0Tmo+JGUR34Xq5v0074mtAaZf9k/HxzOQch9KFri4sP4A+H8kf3TsMZ
BGDBdJxYPEBx7eGEdRd8TRGj01NhdzG+t5c3BpuTwDZZ2/Q+oEBamyoyNRadJTELKXj8+VaFNv+Y
ZzdkGusZIWeENx0GimZ1uX+gI5P+kA8dZGB1aetEEuRvJlUxCDoJKz7nVKH94JKD2Ryo+iu6kla9
9bv/setUMK0ct3DmUbS3E9rSxivlTDAO3cWF1fPJuFvBrfuEHRfAy9yHzUvVdrqrKBclSm1IdFu9
3ymPUB/tBfsrVqMgLSZ/62hdhJhbyglpLSHvQmOZFNnCnou8TaxYzmWOOkQQLcfCaQDsAXVUqWMD
AxzDsu13uwpEsrRQ0EskTG+rQNUmMOn9e8Cex3KYudOX8/3PSKrlMYGvmK2CFKjDBDc1ZYlM2zLS
shhOG9zaCHsJ3AmIn3iTPeUCGu520Ddcm7GvLkBdTh4A7rbgZ7VRdnRXZ0QNfH2JSvJ+T42CIP1i
Zc7NQvHDRfEkDQVlL9DNtNPspiOxi4XkufohGTNZp213G1Zq4nfZ0HNVit8ysPfMJ8a2pMOHIxZi
meRpFA8CoDoNyJl3lF42b2QluzaD5nK4YpOHBTJKPnpfGcbQZYgWpF4NPJrEsn9mcHOL6Nzi+p2c
wT6fWXexeeXg6qc6feCYqi5ZX4qQwq4bcUlC2o8LfkmX6hB1zugBySP2cCakcLQl4PTpkt9BGvte
FZpStpclQvBrUwGc89/GzTiYeQfU+5RU7sHHlYDMLODZR7P/Beey0sxsmxIuCHlXawZCIgx0PSgM
A6H4ySvAplgSG9eEEmuKnqcq6XsPaYvPpfQcptWBV6u1VTS0+t2A+xuUX70P+HvyFQtCrT51nEi4
NsIXxKFPKL2TtmCnrJiKXqKszHjPgMH61Ktl/cB1QrQf8/zAYww6mMhppyvtDceXJoQkpNNee/RV
nL2CUi7C14B3YEXOMvKmNJvoogtROjdVF4gyUwi3wOYfIfOIGw7vZjaI1ibfUi2X4a3Cy96PQkMF
09lr3aAOSeCyEdsevN8T23/6+ZZRVtA9pUTZvbXhCKj5d6Io4OFQ5oRerwGoIlLC+QteBExj/gA7
xdpgvXJXgOGhn7K99X4UgGVbH7ijKkVTco0yZcT5dMufpo9EoEaGbYbh9A10SjxsOO/Bbr2F2Lv2
fNsDqTqnecGMWFXDnNG98Sf57ZsWeRK5L0lBMhvWnXtqU4fBcgg/yLAaDiP4xnAukc319th1avJb
syW8Sip9M2n+F5RcBA74w5qHdp6sv0Ek3qbVCMe58QtONVIKjF4+JM3rwxXH4bNhuv4SK0yT7kNB
9wbi9uXqVe6DRy87iza/UfiG+f/aVKQtQHrdQ1v8GWowbgtpcWDPZZKRB8daT8JgFJPuMoKFS+iO
a3KTrbg8S1ff2JQ03w9iepjsemAM3n9rMLJgy/P5JWYai2x1j+HbE44OYlf0J/EP3R+GTSO4wsqx
QbhGJ6Cl4il+DZXjVsC4/jHCH0rhRdugZPWMboPS/DffgzVDMuY9d7N0Be1jPiarWGBUGvwCEqmR
U00zBA9wUjhczhvRPpG880AmnXE7kS9igquUtbXutgV/YDnLjaylxE8Z+yMKsXuGHdDD2+vW2Del
kMnWfy/U3ipkM0eO6x3zwF1dlQZG0WHetjQ8UB88eCjcPC/H2LVvBkBdqM9oEWg82vD3mIY0K706
Cwv+EB6RqPzbJLbOowVcLtXHKqfWO5TkUC8gkJJ3wpzn0Kpp3ZeNNeC4aC49U6ZMZNtn+mtYb3H0
fRqZhdHiV0dn6nOsPzLg2EZnNwTVuJHLyWXcYO/7/QLervKxODKzCt80M8GN+k4uMF04zVOowzco
dyhoLNgg7Iu7tDConLxY7sx1xY9j1yFYbtBqHNoZIcoD31l78XaEFdbN/Tw/gggKVyz92gUXoZM9
AtQtuvRp/tMzFq4BJhdc/s7SDFoB1fgXSNzcBaBYUGyZLNSBA5xr/TuJSjnyo6mDy9KP8EjPasCh
ByqRXJPwFsuO/6ipxnTGtaUv8wSseEhy27xZ9SLgHeIS65EI3DL6i66odg/QMnUdja2E8BrplCzQ
D/6RukCvyPYgBpXKVliRxG9dimY6WVs8o+9QCaEuKM9KAvhynrSl2vIbekubk4ld5JeoOm5xpZNh
UNlaZ0VWKWZmBft2Wd1l/sY6ywA+ezloJsBsiXJZtCing6kdpIzfFbOqCTCp4bMoh0Y4+CYRB9lo
f/oCBKW13E+8VBmPFjDgOXp/4DgRviMTmGkWvv7WqV134S8rhnG8KDTRDl62oUI0CoZx0K95wF7O
tE5/1KICJzAh1VngC7c4oXKDtkNr8JZku8uVLpagDCp2Nf7xt9imC+MrXqQ36l+qJpm4xJNy3Wme
mcfWzh7yAbInUOmv/Fx+LCmsZjb8+kXJwKMWP/m/4kJB8czvdBZ8dRHZgAuz2G8xV06dqVuzXelC
/ptHRoBH7snTTwNEZOQqG+AxO1yDahY1xP0cZPIpN4ZJr8zs9hkASsf9uXuBliF5ySvuxoggXxJn
NM6oZ2BYCz188BjCsNAJa//+EVQi6BPTG2UeesrQFN6b2tEV3SpiSMkfouPM+BdCZ3JY+NyFIrL2
QzUExulH4nrnVQGNis6cOb2Y7FHs0mKWg/deCt/8GzWeouykHUM0kTxr12bROKgKkrdbdik4K5J7
Ih1aLtLmd0Occs7/wWrf/xvXxpOS28q1opEVh3o8TnFuYsmxZayALttSUAjLhkdeQQNKhNozqX/6
b2YaPvcIEtAR75H7gh627vJBV09oXg5UCTLa6HuNh/brf4jGJJ/E4GRh3mCaqDUiU1HG55Fyx4Qi
KjeqTFOqlrykBHXRyV3/Q6Va9MWVY1/kfe93tYiizmXAvZj0rfg0aBF3N9/4zA0wYqs+ZBuWX1A/
ZnX62vLJwjSB8MkJzmluMMl9gNksSmhJuUgYWfkccOvcHZJcUh6bKX1ydD1kWLqvPqKpHVJ6Eyh8
IlcJZ2qPL9TJZkG8jMfzdxmD03TpIek73w7+oPlkjK8GsR7il38PhFtxgUHbYy/8N7jWvfr5koOr
G9h8PqhtZguSuwi12PzbatspdnbVwHYuncyyMr+S3D17glt6pnAK5q4lI9eqBJGXnpmHfQ0Tl/gB
munzPilwq4evpaBD1Slmqpd+vF5IhlUUzdO46AjNbx+yHZ6H248sB9TAQWpgiQd4bbO/qFrQlddV
VWSreUXaG4Xp2yJcqiv/S6WHI3EfH+ZdbHiil2kmcdCOfZMkB7SN1Ihl6o+AE9V5YMOcn40+2Tms
MgR9GUTuXh0DjCr+Kbi813UgjKXi8umQ26lsYZ/XDJCnHVc9HLO6oL1LWMzQt4heWirOtGuLWTiQ
cPAhdtnrFfXMry0UFSTTwheTQtfq+idqoFtO9xCijZIGh0SI+xL06iCu5CJoFCOTi85tb1H1h/5d
XP50SAkilUfSYj6OS/1iyDFvQnC9ewE5bPLK41N1eoVCOaxKQxBGGdHVlkAoYjrCe5BZokn9sYmd
aJreFdNsasvJUtsA9gG4q1YSF3JkQKwWgBSvnXB+bsN+TLbo+/gBlwrLf9TLkJ/Idti5v59RjwKS
/Wp+ELbtR/xit78qNieiHtNBAnme2i79+17GZUjXYQtLnamy/9B2SHzAvrCDBqOMF6AMSxeJWkGF
qXDQEbEtUeXY5n4GmJL0r+mWiW8a9w+21X38uFUU9HQo1eQ0sONI6ldHwIL66uv+R43EPSqI6c4g
vMqnqGzOXPmKDnZXUU0javIU/2PVHhicqfR9idVts6u6PELb+hzHT7/I3pPyYD9K2xruof1m5l3a
RCHG77idmcMbNKyJtZy1rpEJhvER1OKuagpq3G4tYVh1GDwmFhHz/SloabrY3ulwUkIIsefou+Ob
tMs0tvtJDM8T6Ze80Ggf74xN+1Ml+kBxEbPB2Arb8TV3si+1815YAdpbJAPcQwKXjM8xkg/4QTV4
7IDrDkhStHxREm15234LxED7VQ+ReT11KV5f/qr6qnMXTjXP8jQx9cTJ4n4YMQbOHqu79tiJMyWm
EcgEV+0N6RfwCgsMrPHxYsdoVi1UHjZmGgqh0L26wWPyJ/z3OqIWvmRAJbKFuDZbDtX58NAAxA8h
GhviY3zSKqKYXjKpmtM7VPG4tlqMfFMTKParzfyUuHUD3tj6buaFOqRBE/azxPGcWGkJMsdh4jmd
kKGf0W/7U+EmGQiSIwXUtuGuXMcb9tN4CQe7BMxAeAgvaCNO0hv+Yb48l5pHTpsvATHrRvvQmJV/
zsur5PekmH7klw4s+e0ralhfWNb0SOgdrCKe35PX3Tp1HWxwworAz3VC9arX97gM7iFcqYejHpzm
4hN5LJqJJJtATeEXBXetPNZp6JFSYz3v8SPFDuLiYNUL6GVNSCnM5syjyspUMx5wIacw8kLwBZnm
uo8nl1naT6zj/OZFwe//siwZq7TypLlwTK2cqP2YxN9cn45dwSM1YhGpvPDrwTa+bynvYX6VeDXt
mlC2KXOlPZghpNru0ed/wgv77GQGGv4T93u/Z7/+PV8VUaScwUW9PpLWJvlo0g1mh81Zj45GoCG9
nzfFGtw1VEqaU6QccUcKdllCgspaeRh1MCns5x2ImpsMcU6USDQoThFbdunga7/C7bjVmuCYhgSX
VOZ07/Cf+QMKGDSVY0UCJW6S/H4JqApVUoBJAQnd0xoHhRV30HWxmDAV8Y4hxvFmEZa4o/AFGfld
e3ahd78NAxu9D+MQv+pNnB1I3sADGV7j48tu+hWDJ+PvodRnMOwHxzA0+3Vp7pVz7q3qShZQO6AP
k2WpUQfMUcUQux3TJ2hNRY4nXGbJNGScFw7s3RV0T1SCN/hPgSK7kKhp6ddt6B1SXpNSWRX3sLXt
oxlzKVfxJIIxS+ZT1RyGBbTYfMglMwNl/GrKA+179p8nm1sve7KEinLuIGT+ijZthkdMKOgKSvVX
qtCLQfo2nJyeGXeAnK477vDogkB6bd5z9JV3i/1ltm9sXPMVS7BXp/8JMaOL5dkdy1SNyo5qGhOp
/T4VnMmKFdwPRekLCQm4MdR/LJxfXd0S2mjF2LOtg5+stN73h1aoc9Md74++AIperVGpulfemTf4
irhNe66cJrX6ClBl+jLWrSRBtl0Nhk53WA6P/TcMoQi+tJObLgS1YM9SdLaJ22RUCdiY1tWmlL8y
VzzF2nsJXQhi8dn32mvOiD66hTIeooNPRO32YaOdbnYA1EuvsPYCPGLnk4rpiVPyDpWHt7dDeRJc
fZkOCIaZtBIqYoD2e5SHSEzqQBp3fXQrHegYzT5f4U6qD0NVr+n/UmHlbaOJnffrdVp21p86dDOc
eeDpxXnhBLaaIXNwgvg32WeKJHDAKj/7NyDf7Ffu2gWZHLfai9BHNU2b7EadiLe+zERimxINwikG
TwH5M80+2w+/eVNaSq+cyV2JJRJ2K4znE5ZDZG7afbd5UuTGzMwt1qCnxamZUGNU/blxW573O0Zi
G2bX1EFSDETw0WqHzW74KVztPH6xrD+a1oBOh0jGfDSRApMJKsz7Yr3RSKXp88FI+Vh4PQmlqCYg
43XgxcC7i+5SaZ9/MG8OBXVa5h0RqakWBaZFnkuGGSsSvZQ8Gd5eakPv2KoFKgDcA1rYZDTYVEBV
PM+XQAqCn8/Bj9aPf4cJ1pJhya3QtZCe59emzPmakAmK49aw9DwKOv7LvqWxWuj4RWiVrhd2rq25
D/QcCI3nVUEW1MiTYj533sE/Et15EgUpPeSx7DZwPn8bjzYd9o1QBRBjAEsTF6wgOtWhllxXSa9D
2hyHUuu5XaFbHQtUIbRlo8bA35Lh0FWOjDOHQu2Dhu7tyoPV+fDD4X02nxc45W5AyepffDiIKKxE
d8C+g+lUpYHBd6PEfjMeXZoFBUjSHiL2xjXv1Y1CfOcaR9XkrjLBBKaFVILnp8lr+CHUsDvGL+S0
y9uM0Yr//kOAIrDx750/fUmjh0I0F5UyVwk/xPrAWlTsLL/oAxqOlvWrch1fQLI++JAmqvw/Yn3H
6S/Teg+bTAnHSpiiH3KdELBhHsjN1vB9gENkkWLcSZ/CabIaTQTFieHDARglsDmQTOaiOu8O5/HH
QyI+jGXqGePZVFaqEdo6lA9JTEc7ID4SF+sA1Q1qQO45KK/WDUdMUVbsXeLb7uBuazWZuDgNIIFz
T02S2mimCd73BYO5p42//EUYHhpj8PZ3pyVajq/PAwcIYQRFNSwRz3KG+1osZR0iVl/dRVfTn3OL
Cw4aBEvp9M0Wy95kWTeKmhRTXOIqc6FNngxqHm2rtCDNYTN7qS5mSlLh1u81eCFwu5cfhmRVXMvl
mLEmfSH/xjiYcXs6/QdYL7OLJz3uBlitlrtDohizAKLl29X2PEbpxIjVvkZcZYYxPlVYGcBIkaQ/
Iebh+Jtf2f6SiaQLWwK/lM3VGlUulKvHObs3YGP+RWQMEGkfXF3eLiMApn6u6vaqCcCNIQVUAmpi
WRBHDfcAIHR6AgEEPHL+RELmoOa6o1++G2orhF6NUBl+scVIEAuKitEPpGpP095OPl5Kz3NVhJrR
NAHxaHw3S92rZgfQ4cVUekOPilWG0AzWGvlVaGTVTCxktY1AAlLiVXERxY+efWIGGKcT6cIVC6uz
uunJ+gfql2TK8TH9LjHgKNnPW0Vv6X+F5vA1BJ1RDJ4xKN4wcGA8qOuR9tag01NbwhO2Qjw4/bUX
JEf/S202QePXJ7/1UB31IwfaDxjva+WaYQFsQsd6qHFqo9TIbch6FfAJTtykWOd7/qZiiZZt8UrI
EBOVscYnRoC286kDvNcbyjBnL+bUKXFpIdp076CaGaJqwnik3RJfLf2+kNCu7T2D4VwGTo7HY4kt
afOxqi0Wmj10Q/AG1ri2oX8iH2ma/7hhVphzPzWpjfrPlnFVMNJA1NfrAXh8pGM5onHjcH5sGWpZ
sbl2ZgLj22TyasVuOCVzpflJuJ5mVfYR2CDuL2DRiL0XUzGJ6xsU5Ghv0cIx5oWcjRpj1yMk9pUx
2WUpA49PQfU/5PK2/1VCkYwNx4cO9RJPJzmyiMsfeoNOycxBG43UEUhLzkZK813hyRDeYAVC4PcJ
kW9CxFPDvbF/eNjzaCIA7RVe9vbjD/X709h8EZDivDnnG1W0SHJb4lxMdlN5JB48jEmUCRA8VMvw
3Y8K1NLeBe8NQQv49JYVNfmLzO89xCVeZqIGA9Dx1vLXmuqObsFx1WXR4JSvvZLLkyxbLHQjTCON
7FzFb30IsMleeV2BcmTHLXkdaY5gheUw0FvIPbiS7qhlHvBvdJ5GV+AUdq3DQpPd0Y91ARN1boTy
hDQlTUwVB0zxQZKOKcbjWOrXSzkFYsOx9/+aV1E5XbzRT0l7vP1VWwR6ZNFpiSJNMGhLiXUvhCTN
pCabG2OiI0DK9TUd7EDp9RB3vt6gXBrgcrw+I/Wj+VkrNiv469wwrx1oV2T38BpMnkth0xJsOjI/
Pmh/+9DAeAYlKgLyf15ixvabgcL8L8GslclklGXcol5SQrveYe0vcmsX9dULn6xuTvSh6hJOFtKo
0wPgcYH2Kt2yPz5WmXpUzHT4Glf95fHNZ7Lv0M6GFaUOSjtW+p1F18CqMzMlhk1wcgfv5ECFOsW7
1SG+oALsKNdjbrCEO3OH0EUHmxri552OiZQEvd958TeiPFhHChRCsU98cxgAcS3bm+KKZt2QQ5c2
LHdOutYopXvhKAxdLaN9mq0HB6s9NLoAfk+CRsxsdUmV60qemHmgPGf3qLSWzzo3zW0WLE2Jfgus
Wu5OJSmUvHDbNMiCbavIL5Q4w/m6uW16B4BSw6g+iZE6g8FwSwX+plWWJ2BcnYLKbXHx5ZGG0Y5y
cUiisYubLLrvJPu3ldhreO5EJSkCU3JCz2iHAtrxEiVorajI9MUjITtAzrsHZY0x47xTSIQwP7XH
hTN6ifk61d257Y/G53f6ztomHG+78HY7eX5JVJxA3ydC4xFbSI1fgWBDKzzK/mri6BfKYcGu33pI
8+tYT27sMLXJMHkMfpjcdKWCRbukjkZwbdZYkhXRS84OzDatawPpeMMQVN69ur5Z+joJayLbf4mf
ukUcNCmYPQfT30ejUIVSPAe88kBVXjg/PM00tlQrI+2cj6klEsrArJviCNLXwV03RZMFOrzSeh+V
Zfr4I5dYO5mEd5DafSmt4XzHbTGuUIdZAvItgjb4KjrFqnRY42ta6UObS1s2O65BFDqeCxuUmst5
kZ2sQ8TG+sF7hdH7x5upfPE3dd7wMZtt5LQijpFffJL4JfdpYnzbCPHct3jLm/PCRFp5PHp9Itp8
LVVBFq0rgR6okT/5PASTYagp6gesBv0kpiKsezs3emuLtQ431dFE7XyChfFlkKK3QAIccJ2+Astl
M3ypgEZ/qPY0u3Mp/OONg00wycDHwfCmVNEJI1pDNjjInJHz4MhwR6PtD+U3OiEsRx4Wx2fBzF1k
LZChe/BmP/EhwrbU4gQbz89HeKj+MFIxcq7cegFMgGDyCpzTRe28SmYPUkv+o+VeTe8RKWdtZEJb
1KRjtwRSmzPTUHZQCAwEnT/HGBv2KIxm/hXYPAdefR9ZwnMUrnoEfSh9FkUQns1DPIew6uWo5Xx4
gLpQs7rh4adCrpBcVvChPpoRL6CGwmmAiin6ynvt1gsuI+9BNjT/vqVZw8YVIuQLxEjzrxBprGmH
Qu2H9NdxaLfHOu3Z8zBbELkiytGl3cRaHqifvsFoXrJCBChvOaoJQcXmhQDp1gYrIfKRISr9QEtB
ogxMXNhe3AO6tiDxdwbAr2F3OzSFMNwOp+l3ph+OnhS3OnB1WBRDOg9GtugmmlYkMCe/nBvvH13f
oD5Gu5ZBnJNx85ztNlDrEVfVJLYaRmuP1b/sKEjPu3+qBaWjjMXQGlMRQIoibxUsIcCKm7aMdWm/
KzUqAuU5mUiPGvU5I5nFcdfG3aGXMax7sMPPM5TVKS0sd+0S628Uc7V2lDQ9/EhI+7s0H5M/u0es
mFTWIXSQ4Di5wCcVna1E87fQkuFVJjTmb9r6QZ29CB3ZithuYPhJusLg6lMwcUrl4n2HO8Ak7/cA
JChxQE7pnvnGcl0n+oh8BA3tatS75F1e2jQBuiOYGeCzgOeiMFGzmTsW0RXVmkgpty6ih+xebJyo
67K+2rMiauwbSf+8x+rcpfgDTTjemkfXveKnA183PJVkIxxwsMvgOh7sgkBGeET37L1FYBlJL4V3
seElDSaZti0QVzC6Rwu4Z2/hAnKXnM/nPD4lVEWS2Ok+fdQvezvNgSDZdrFyNvZ5j1x1tTTCCx15
cdf621hYf965gXmG79H4WAVXMqED4pzGnuK3o+ZTt9jH8BE+nDnMrBWb7hRoGRwDLaMBp3/LvquU
rFCKZ/pLBR25xaucUsH5//NdFihFpYBCRllwLcLfSZNdqho2j33Vg6JgaTEvUXcWOxciM1olsjLw
9yVkdcdvGphE/2MnAHmMzEHV+Lx3vRI4Ac/WyaIS0F9sA3BBFAeNSn0OJverE6CsNLA4pYJv14d/
NP2+Oqv3fttqBS58ezaKYW2RHdI7PTr27gqOY9t3fcNiTjXN4dimVpiXug3Nd5v6r0r+JXHuEmCr
JO7+VwvvxxD5bzdMzneZ28d7UV5hJuK91p7ct+0dvomlHFJU940nFDaooSGv+e64BS8aPsZcyHe+
IF7zOBcYnQv/GHXpqTVKfZHsdxaZmEBEFV2fr/mrnAhxV0YdifPoeYPMu2EvYLMOPYAit2GnhSFR
uDDWd2N0NV0Ajp0vGsnIoljzLtQvCL7LiDXRnW7y9ZQML4OEsgjNShH74AsXX7p9We9U0znQBGCQ
Xa9cF4a3HPejUqWGPcLhkuCu/yhUxpe26Enk0KPitGwM8yR4zm3DsBkVyWCeGPmJAlrWRQ8jFwX3
3bKE+f3AqmPK+YWhougX2vfzWT1RXdjzOGseDSJopB+E7EWUFkXuOX5JgwP79g6MKAixA9U/X2Vn
vGEIC9D73hBV7cbF9r1K88ystWbpht1xZvlARvqqbX1L0YPfU1aqfL4ABZRcEOTzcnJ3WtyJllqp
DtlhESMe/gfc6xAkBPYb+51Bcc+3jcQQidnQx7fGqBYFWbw35fCKOWtLlNx4yP0bYHJlrtEBg/yO
KURMDp1Z/9TACN6yA0XFZDFRZhG6igv0WVjCgUFhPnzCf8K449Hu6Ob2UdKOwUnpI0JRvfCPacmC
tsl22euTE8Kkgp3cfBIm7K97ZqneQYcrzwd/O8LURXHTDHhabf4XPvVGZEF/xpPYYNfFVpwq6g2y
/bTuLG75xyCuVxPX+Cz9EEcjIs3DmAK4hwVf7DyNu/4X9dqO3BhvOClClIBxLRcK4bfrQYi2NTUM
qD02cCC8hXzAAgoaSsKEP+a+02aC7plFeBlEnZMT78yzXrleQitWrqV5lDz1i+ozfHOjLJ6/1N8j
sfI9h3uA7w5Dk4cuiwx1QQAHVOn/ic0bQ3MGftZfEwTfkmd610UtUSkjwo6IYkBRt7GRQ9vcuXhu
BkJFRWTeWMoLj6jETD3YGOetQRUQZSurInJOyjM/jyc4q3muhSV6oArN2IU9HsMlYLl0fDAyMLRO
KroFAy7i0CMIWw4elYBk3sU05vDzaX4FRANEm5A+iX5mlx0mptMuHZqd3BqosheLuwu9BruFat8p
OlgbSuUUySu7Z8TPc79GlBBOaqhPf6n9MEOx+76/jZIkkzZ7Z8EXG1EnsFt7oax9EdHzHL+u705Z
neLjfHAgGtpT1bwqJjDQOMq/3yqc6TqHd+X+zZu1a6uwg9kYgSDNlmYK9/rCXlBzvAWkZgWJ/9XH
8d3Qrb5IATNY48uhXtTq8MYdKnYC1Cb3brGCoY4OaOM1B38yFNdVop+J1btF4oMpukk/svc5n1Ck
ERV9crhWsn3jJw/XI8wq07wRvZgp2ytbnU77vgBRUBYypn3wmm6fPJ4ImBPAKYPyz7o4S9A+QDUB
zT6mqFiTp7rwjQFBhGbDHNaCe3c/VtzxT85jiQ+/9qjjClkkcil4eOQKtuK3jP31MsldG0p2P5u/
sOyRJ+ecVB+AAmZQs3mHkC2M85g0GaufHrDyhKBvxjWX2fQgvWL4+YrIDnqSTrqXhdLMQMBhSmgc
ZllA738ziEpKbhnOIO2iNA0Ehnd4l3cIqYFufQdG+Xj7Z1xWr+xqOTwZT6n2lHcthJTJrxWyZOPA
dM/++tjQt0ix7VcBZRCplRKXEp3CMqAp/MJThiDNLUCYaKNqWIrlCz7yhMzNBr1c3v99rcwrvRIA
+UR59INd4NMFN9OpL6mbrh2jUkw1E1eYMu1V82Ew+EqFkAPhaJSP4pk7CP6n/3lYPtFSZm9NwV06
7zCZvmbLLVBDfnZ2VNfM888nirIaZ5bwblFGIKCeUEZteL4EYS7vh3naa4LOQ5NxvHiPCuN5bquf
CB3dlI1ul8Smi6x2GnWXxHm5uFfHGw3dzPpvw4/cOsBBOhuX2xpHNb/Ll1J8kzUD3hb8YxZx1xlf
riTbSE32PtpU/LfXjV+s/7aPG+lVE8CgMp8v1ENFgYVcZ/7aq3KtQU72sDppxDqlpK6b3LchFHZ7
BWtVwLOLpAy2MqEYfTrZ9KmvnEfqKC439tWq7XJakfBuVfMaMQkXS/I8tpnHwF6WkdmGggAQ5BBV
/Mt+D6yVT0BKlzjO+CqMbZXe5EuHo03EEU1vvfx2ccwNpeDYke9OdX6DcUO9gpiEuVvcen9SwV5J
LKGGODtdSc0HZ9kf73rem4Y4AN0v+nGOZ3fg0B+4s7N+t+/Gp8sNqy8vpWYi+IrP4cHC4E7P2dr4
KvMSZznSnlNvbjnAGld4lKVgGsMzpfwB867O3ghMyb+7WFxzxvnDb7WtWlkRO3p4SNP3gGcT4bfJ
Z0MUxOL/J6TsyZ2mFl1m0odkvsrburMpthjOOydIX+cRd7bSNX2WZ/pN2UJYz0cNkTO2/BmOeGhy
aEe/y4RJzpRv4VyYAVlx/quHDNLnc4H7agw4RkvBErAyAMkTnAAHjxsSpsUGYGiAjxVAi0gOTJSo
aBDyB3CW4m0hEe/mnCKEHj/rndKduGEwakghnXsc3pfoMThBFkA2lQZsZATitSOUMTkmyhFCLexS
0H3KABGRdhi3gTYlzrgCn2On/NOCg8RZ9ClwCSn+HkpTKkkPasHWPcXuOoWRU4QssPiWJ7jiiiAk
PuYlh665ZjF4wjP1gh990IIJCtVm0z7WEnE2+RPHloKTE4K8Xl0azkDMeY9pcQyDxOj5bbFXK4+I
dE93/9zLVUDRN1y9so7mj4VLCs8cZ1/1aBOT4PG3wI+xQTkuRdogGFsdRZtThHsxMB7ImDkoALxr
wTEBhXQVnnQwsMbC+VTA/dgmZvHuUY6IUvF9xx7G1gMgtHtS57JrtOekNApYtx3SwTAod3Z+plZB
8VSs1vGLMpqAl9qy4MXwS4YqzDn1pKKIWAhf3DmP4I/9EjPZVnvLDGHQFXhdgIw9qpFgeo8+tMDM
p+om7bS8ScyHsgA2ZTbKRfbR6ZQn31gHj6lvWHdHCK63WXyw9QXy0t5g4dJidlC4AMI9n+EFgxWt
aDJozTQXhV8MMPtUU1Iwcg2ljKZt3ufseO1sbyn6jR0/P03cUST73aUAj3u2/RLvP5zSp6dhQCsr
gPl6kGNNyqoXbcqHrvH29tdmaJ36QF96aY+jyC8GQHF7u8Mk62e9TG55SR1zwwYov+IvmG50G6+v
kDmou/NOFJYs8yWcydWF6/LQ8iPsLBlSMogB+cK27bRi4cEoGSGCjDXw7AzTY94ToOBcCYN39XLx
phh6GZsCDeDbtx9Z9l/kzPLmu4GZyIdeT/X2iWdJfaUNQ3ywmSBJE9K10KiXsLJmkIlVMh/Xs20x
a5MZU2Y0ho+FHzeP+oTVwzpJ//ej4P5pwycz/0tC/VpvPbrcq2HP0w8ar2+ycvccylgpmGmmzZiz
7IJ/R9NeXo4X06r6WyI1VlAUjnwWLA2UMPRcxMW3gzVLjfTFH8Kq9XfnV4esFp1KW4v6KMVQUKpI
xYZxC+B6sRHqoF9lthMCT3PyMY5gIba0o3MI8/OKINR9KjMZZ0c6HLRzdLrMLGoLrJGs7mkh4bmw
wR7KX5V/Xl9Rx2Rli/k5qCZHspXcjTiLfMjaHF/jRdr+cHqQfj9OyFfTuyOOA31G8duKYnkL1JBE
paG0UMunD/1ywVdz6pl98jqh95K2Ufhrl43/80oo+tO1HI8ktkcGabF8pHmR/v3mOEeOCKabYT/k
RAcIJzfZNELR/yiwPk01dMXZDTcrwV/eylsXgdGzMXzhqzkIQ/wbwij1mUqEj9fbn2xlPaHqkOQm
0AqCqA3eSHUAJJEp1Np+mrlER+aGxcN5sVngcF1HO4yb7UJlbOwTVkao6DkCfZ8nVwLpxEoT76xD
Y7vQVHFH5EadD8NWN8sesNI9aHNJkoEAGRGAaG9b9Xk4gpIc7pw6uc9PqOzkZhwNrZyhkL9Hy7kA
fbd4C2aywelVMgm/6i+kkXfhwnRPFNi3GPAYgqjNVnvcPnlgRnEQz/Q1YbVYLDRtkIFyoZzwiuJP
sj86hUFiy9k61/TnrPRnh3g1ExGSY1AhHMxVSZAylt/7V5DassD54ujTFjTlFDFklWyWqGitTqe2
Oi8QbIC2/Pm7FK9oksnK719KDx1WB4ozvyFyOKPOV+t/V7ykT34ZvAsdNgdARm6vUVEw/0pI5zpN
svkQXLkZRESmVWDZ7W156gergFCDBOd16QbI4RoD+QnNB+3QG0UeJM3PBw1gwuGgWW8KtTb4V2Rn
kIsv/wyoXSNr9o8vWfMEZPXQXz3K08//ReNCwbpMfUKEZJAJUkANXcf0hEOpVW9gwwCpTzKYYc5U
8z6oHpqiZG1B4EXP53WFBoAroh1seJFnpU0YLSZTk39Pp/8qsFb/YIXQY0qq5hLWofZpLGuRzTPi
KLC4fSy9aYlQdvyS9LoTIXEgDOnGn5HDE8pbPo8pSj8wGld+h6TKb01+yJToZVjoGubb744yTslB
BgGjUfDGt5ij4QsX8yYVmSqTynWJ9zIvMnI+XDiFZv2W2uuYcf0JjEQJhNQzdeRw/lnpRwv72rqw
eM6X81iquielyQIwIjfeqB25N7yjVQwN4jCCgzqB+wR7qggqEC6qhIl1omRDIKzZcZ7Jh65qp5Ln
J3e76ftUCy0l0+EPGYb0LdqUa646uSOVJWibo183L6LpXBci18ooU820dP1mJjSVCbbYO0rV2k89
Y6+ON+ncfK/KT9rakoHABgimJ6FempWI3aUkpXFZwdcWaaEM4nxHJ6p/CdRYDG8i9J5DwzK/cFZb
3YEvVvkgWhlImV/8S9DkWwrZuFXA7iyZir9btfGxTz8H3aIXz751gloQM3xqgP7IOLcGj+SFTeEH
Lm0Eg4bIPmRvMhbw7OYYKN399cUoVQOqGmvQCxOd2RB0HGP/dWFo8W4xwHVLubPjnqAaoXQh1Ot6
z7ZoWixHWGOGTtHquU18e6tIVWeuHOjlWVh2ZO9ppKjWHC2cYyZvwYdyo26UXdcTS7pqHDV0LxEG
QywYXBUdSW6AFcn5fH223GSsnXoVnmgCNdvusGdzXGInGEg5jk3y4gizyaQbAIG1UmVhF6nrtlzk
TYsEIxZTyOj1KihEnC2nXIxVr7WimrUVtgvUf38wxKdKf/zLWHQEEIxWhAmkH9IsvlTWcxTarXPn
0G13NXiB+81ujPNs/2E/21qyjEAZ3g5LG1bPCbbzT9usoVo4OyuPaP248Tr+RHfEn1nWZ8XeL3xJ
XzKbqAgmaIGVWvFTxOXXoIuC/8gReskQsE6ILE20gqnUzPBZ0fZPPixX7fyeBhBQBLF54shXCJsq
Zzfc7IuovNT2H53bQqpcpfalsGajnBdTH2YDc3JRzzfVJd+b/gHuusdVbixs2nM6Zyn7c0m0un4L
2hZT0HZptlmzOl/EC1v+rJToIw57htW0JePTIjH0/TV189rUqAS2Ik5MwE0BdXHgyLhG4gVvPWrJ
ngG6z6HpFMpkARrhT+sGTl3yCnIhbdEDHiaBxkjvrI51zjzrXHzs6HcueXhe33OzDjYNbZk/peJf
nSkj0H5s+aUnJo7bnwkjhMWZZUaB0RMtGcC4GmvaXlHIR6B28WLudqvNeRmTzXUfDmn2y5n1ywcM
iQvYRd9HbvZ2I0INFE/byMaIhsN+D5sNzjsTTVAtzRlHk8q4K5vd9/JO/Cvjouul3+WSw2/JzbI9
gj0+P/T7kH+DtWu6AX3rDUm1wiszLmuW3GkfI/acL51F7yeLdJ5gal1VkCB6fcRejnTu1MI4u/c8
rWqp2Lk4LI4wWYJKgoZ1tdf3qw+n0nQyiFoPAlNF6BUq75ajTjgSdEthTeOkmdnktn17YgVST3Wb
Cu6LKgK8QwrqLMcQ3tLL5c04SFTXE+q1bIZ+ihXiKRSkAtPXPayI6eIdmtjgvw0D8tyXQxSEAZfw
1xgRvMpfKcU/E+4WuoY1OBbiso1ZDYyZeJTP0NtWO5zpGKy5vkLzlntUJINBKVGtMGD2lAY//OtG
EHz+ys7abmDY+t/69jE8q06ehkdZb9rZ/hFTndwX8fKM7erzj8nTmwG8XuVBzHkhcKKU6Bg6/9z/
hFdxL75GRIiPlClJWVl3tiIB8LNsw15qrb97Qd/HCVFG8A8hjMUN6JfxhC7cbNGqJI4bk8eCqRI0
ZyickNC12bluusg+xAmRQVAdmyT7Lv2eJOwFX+3KpFoe+FL7wlUjK16ExGhDuD1V08ypYkOnpqmE
OQwaNvoB8wBOxREjE4or70ui7qwDPKWl2u6VI6TDxYQ+vCI/akktQxO7r0AVJUXdHab7DiPY0gNH
d24U0oYi5v8uzzMpdUoccSQC2vniSl/+uFbGNhGkrS++V0Ko1hMTQNSlTnsTdeqJUXL2GN7Ogyfq
t6XwbcCiVwwNFFKQPEmbPimIcbFNaAw/vPkWiGnx0/ozCP4Litwfrm1efGHevImrEipBLSVd6L4d
5OIqT25uHgUSJjeyPSRmwmsbiYD+b+GWCbfrWpn1M+sZeZ+Jp+u9KYJcc7+NKbfi8E01GvxRAp59
p3w30se9aZojX1v2tS7bOaBqf3kj9PRYL+kB7J50zYcBTjxS3/zAQ3PQp+6GE86Er8q8WIJBbgC5
RzzcF/EcQU5QEf4kcBwtsEiodcagvLFtv1y0ZQn2uetVAp3jMr8k48FfL3ruXWNLuy9Cp+lbbMBx
YoNriAoGL3E7+lO96ibxdg8l8bhHEQSZcVNEJNZB+qDUylQeUm3USEK7sRIcZ8HhemcngYJCUMFU
Py0rPzdN7kkp7WnzMFhJYZ3zJNcf8ha5iNqb4XAdof6MiN4d2tsV3UDhI+Yx/I+lQppgNewwoVlp
KUYoeKmI2L5eI2NGkYuXcrfFwp8jhB5f79IUnsx6kKtxRrK3kXfRFEzzghyZj87GNh2IotJ1KJNw
v5mhqip/PKwgx2WwXWwJucrk1XFRa+Zrbgm88Zti6O0Z5FISeNm2RpLWWM7pncF17ZTE+ovLpUsf
wCDoZb8UhXQ3libIdUsjxttMR5ngDoQzuFaXch2m6Kb18aHu7sOgVCKHJWUm0l/KL1H8N7Yis5oS
tpJffueU+P8F70YWxMj3J6RCtungscerQp0sJ6p0aVSpIzJT3Cq6Cl0++3Jdy+i8PUBceWQAIeff
wsoVoSrGYWvhRAyssi2VKmDfRnO3BCMk1eTxsQ7eEZ6ZOFZ+tWljdmaf5QNVjsmRCFTHE1/59wLo
U7Fl0uifOMVW8fdDFOALxDJK8ZkCNBLvZUZPJPL+5kx/68q3igmDNp/kDApMMYsVhJS8G9DMJrtF
6DdHVf4FuncVSNa1FZO5jXeMHHMOgtagIF2vRUnZrJx9UCl8PjtGP4Aol8Vvj4d+1hR1M3+qh53v
d6gklHodWEA55Xi6zs97yluvs+SrGM7XE0k3R0LFqliTwHJTKOIMe9r4BDc7CLdsw6ZyynbF+0qp
P+KiVnpzScyQwyn7owaLkS4XV2vLnPqwTaudU7/euHdYk1edhpzY57aWTQm8ziQtxwAnpKCpvFVt
W9yF3ny7o3gnjwmLjgGf8L+CXTiUWv8p+Nfu9wLk6yWqeh7UJQn55xMu2/ja5SDoFndtLUb2huL5
EBMgm4z4UjFVJqIo7M2OhewBceHCLWa34JF6x3jiuKzqLr8f1ce8sJu7APV4JHW1w572QwjxF2sC
AiQ626wa6+3fiJLDgHDEQEeP6g4ZsWi2CV8K24vM0noAw7NEyJtcuu81JxVrrx64pckZy3y8YSY7
ejBaWrXefHIXU9NKf2ubkKpjy3345tKeKjBulqo06rWgrSpHit2m1eEfidFTNsVwtb95giPZI3MX
RFuyHi+IYNn26lG6VcHbEfSgYlTjyT0Xg7PjgfzbtnSxVHqE4ISw30VhA0+RJaxmMRCJUdxdjFMB
ct6LQUWpwGlpIrTC2ojIBfxvt6WLF/E3npN8X+JAgAV42JXa/bKGKdkOmyhOWKoQSX+w0ap8+1yL
dJmJ4BQXoD98m2Zjt2e+UIshxJaDglHiJteq3lrYs7HO2InMFtBbE+HeRwoV9ZGpyZ+b4Y0gVFCd
KgEjjazStMvZyMZWHGzck0DsHjkRnMchPG/ads4KdlEJV3OspN7W6lGcEXsOWnJAgfqgGp4V34EK
zBW6F4BOcBxYIdwmgd+2Vhn6BikipSelB0MjJ+2qovcy0+4cpL9SqhX6gmiomHjhpOfxbqdCvGDz
rpSbpBe611IFlQKvyeEwGNRhzbhHKtGjOhcl8Msc6apenxXunWG45WrQEMwyrsxmZtqSqs60PrcX
1Wm0cK9qPimSg32Yom6C2RXoelBXpdvhd4liLIgpD3F90ieIN3Fptk9ydq66unEI1MEiai+5kMgh
+VB3SbDPM81BIzRPTYdiU0yyvwpbD6Vt30q+xQulMXRKZE5rLU62zoT0/yfw710ZOlIMVoc3ZU4i
JkOpFrlVQReiTtnebeSCTWWlGo2FGbB6ZygpifDDvfjgsSYOs07p5tTzdEpzrIIGyXNW/+Lfv1Bx
lYc4wQC99XLgyyYhoFyEiXwk8Kpudu1xt+3wezyiGpgWKgYKyC+8t8oyc6UCLDiOeb/oBmh7+IQ2
O7Vsd21Yt+/8zntJt6tNv7eej48xd8eHoTFDYSA8rcGDBYYY4B+HVEeb+FQTMQbAhopQ5EFwzIgC
e/RXly292IXjXiJx9WncwmPrjCUG0zwv30IAYbXHjLQPKAnOON+ElubU9443M314JZSDY0UdHYlg
7VQDimsY6ht1VcWXxdbfxTtgzmBLWXEjlG5AEtHbthNwaliN9NRasMrqcVUBRltRvPu/AkXu6s+Q
0gKaxEzpOxUh2RaEPNAzNMBns9Ex64fCalOdDp/ZEGNrrbfatp9BSU+EhWNWLlv2T8l4SFTDOd0+
p1Mx0EAicBucr1r4s02t3TaTV5fkD9ox+iem1gE0qigHgLTyxwWMboyzJ1nO8Xe9O38AQtXzczVO
bFd/dIIJqH6WDnn9Qo4CJ7XoduHGlFWWpJSCjlZoeXeZsou4pOjC7P27MvBFNEupRWF2cCODgh9T
JMK5pMAO0Gsr81oRMjrQQpi3RJdZ+M64XadzIGATZmBBYKHwvB+ed6mTTqz9CKaTIvHkEgGEwxzb
NlbAKCFiYrYjr3BU8ooBw0Qqw4TK0SXKCrYfSymlnazW3Ea4YrBJeyCU9vz5gGbfltFDrJgiJAEU
CdCD0MmHHzO9lyqwrecv9P/HJzLFYRM90OdqHa0TVviU7dilypKDuiopce8TEOekdu6Uj485X62M
xQfGAngSiDvUc9n2u+vPDEQ0111R8y5MTntPRSNN3FYM0PFONmA7pLVdHQlVjJUp58UZcEDT8W12
TnLZPLlXjPF/hBtEzuUxge/mp4HakgfwXKf9yEibOGaQCDv/Vr729BTDYndkWmdxYyO+XGqcc+QD
WnOOZeG5ml/mL1TV4/andrj45bU/98siFFS9tCQqoKtYifryf+M/s6snjfbUlFVRjlKxHv7nZDkY
USF7MLiGQkTQ2ceuiuDWEkbo1I0sOaWU7l2XWfMtpsarM2hWVkugYW1eM9+Gt4PqoD8b/IgKKXZa
fvzHp0uVdLZdrXZLgBaQr9c3B1DhV6RvfwdiYgQXPmM01VDjHT9N+IIN8wq8w+5e8v5As5/0rgyk
oNwDJcUqzjhR9TcTgfnFVP7jHmW5eITDJc7xYiMkOJgD2pj4EsVhAA0f8UVMGLF00lMaMdvTc1pp
/JVlaKnXSeAtJxpKosn8+7rzuNoiTSf7SeAewpond7N+NDl4oMuYsKYKukOdTjNUuX6zLbANxvcV
XrdlBd0ralj+bsR6t/Zo/h4a86KnF+RotkOWMpOwsqFG+B769D0CEvr2uHlGFNZPqcMghh9h9R3Q
381zKlyEfqNdWo0c+lftdYESyfPe31QA7yPKSdoB+0m4CLJ+wChuGi5ZcNmL1Wm+vUXl5ofnekEw
wlgCEVvnn/x/hBz483nvweL37smFo7yCXUllZWhAlGC4UP8BGo0Knqihe9PeRKCOMgqpZXLl4wO2
eVRuJzCn9yaGocCliAhI6KghDGXAZavbjKZR0rj+BCR70Cq7V+wR2NZSUmgsUHHSF5vhkql3SWmZ
AOm2bGDN16AwV2Nch7BnYEzwajT9xONL/z5PuTaaRYK9R1Ti3kqwYUPFXoiDCPzeH2gZMUrM5m7o
ewO4BU+ztS1fhwqc5uTKaAcEa0MOccuTAcf6mkzuHGHk3wFKknyEZslZtK5ohCLHqVhUFuKH/QOn
NSY9eAxYs54MDTOdETmf3/+VFrLOLi0z0tSxa5QpG2hWLqsuZkOgHLleJHAqdRCDndhm0x2C+7+0
tfBzKmQ2X3nRPYJbHQum+hl83hEXV9OdVQ6wyUnKD7i4EuNNUXYsyZbrcAYZQI5RGaCApeI00FSF
Badvn0IkvyxZbFiwGXHk0avcAkrAoFmVT3a45MTgeUIoqm30ykecIq1DEKHoVviV3bXmDPxVHOlW
ohM7IRjJaa79Roqdh6zGvqtDnG2gNXOuURObw7StbCsX5tABBC/vmfEgdKFXlHSPi+UFW8fMuGUb
euHkYQ73pTpfHRwS5DfCdJuhw4T4M0RarDC0vim6HyFuCV1oJPvW0j4FkUW+PPdDTNExe9YNS/5z
zlMrQIeV7fTR328E5MzOI6hYeTArLZybP/1fF6DvI0JdRAzqEOIL/PSmpecSAz4upnkzS0mpTQB5
uDha5p/5X1FhGZLhIE6lYfOgx98qMjJ3Ovwr37cM3//YxZnQ7uoZag/fssu8xw3BsIW0qkUepFXt
GDDOGEcdn2YqpDrroJM7Xwr5Ca9/ctNpmdDQOjOp28n4daZSIJos/OI+d2OtzKKnt7X4huR2+N5Y
IRFLz0O+o8ijU4YJZ7xhg9G++NKOyopqQn8O9OXDL1vxj8NDr8svxv+vWNHaHYfD2FtN+0N9s4sX
1HlP1A6eU1FNw3h2dTsWtO43ZXXtq5IdZw7y1t3ivxFX7ibjukBKMMLeVvZExEDn1BdNn8uLaQdj
DzfKq3Do3iDDY4k8zExVGkHeNpPgLADI3xKdk7jsjkqtGDXnrUgY7+uA5oQJKgBhcWGeiN+daMmc
lPWWMsi7EVk8FV1ofRIDu0Y7CL8Ed91VKwHHIjHggLHyyy1nqb+MZxKu/03YAh5iXjJxeWJqC3iw
7BcWHS3hObLriethYJ1DLBZpg1wky2/Yg8wntBbpv2VuVnTxhWOdZxwRLVE7Wf/3CqWPpXIS9ah1
Fh73DFuAXOPy0KkQfqoZNQJureZ699zfwtuRYcYWLB2Nf9mz1o4Yujslfqnws3zSg8MchQJ1WFnJ
F7vHLGK6T1MQlAHocEj7lgVMhwuGZMI27ukYAIVSmXrCGCAYivqxTa8JwVvwVE/jVuN+zxP5qMe2
ITakUaGxOEWoA4Jj83Of+zCmjZoHdyatrGhmfHOfDYIqRYozDOlveC8hdEGsgUFtuGWXDNHczhYo
Kc71SHqBeXdZyo5uJocMda48keOtY4xjJN1mcp37oiTjk5KuOR0KB/Z0DB+3RWzdOVD8BhR37Niz
g9hKCekjNuJFNUooyI7U5Rcem3YHRX60D6wOJaJ3Iqwjex9I+hIGWeWjbuI1NeRysGNvOkpMPP8p
UTQfA/aXXcacGRfzUJw7jm8LweiUHYyIQHZWK3thYG3lRcwnUSc8l/FNEVif0pCX0tVuiag3Qjma
Pcg5o5WyPr3oCV4BE1hdganZy2W2VsUrtxtPjwgg9CYwv/QunwGncV0CPMb5F0hJGKhP4T/GPyRp
YJ3ghUsF52iI/vSAxWN7LKOXBw7LX7RUbdQ9KHd9ctbD2rMdzC0jd/laY3MqRmPdOPM6sZJAUHip
bevYuG4p1Wc3CVbyVLe8yWT/xc4s6cn4D4btAQbvGC6JAaqtHPU3ChS3AbMy6GOzkKmda7JJYHGi
+zBtqU57KCgine3MRzlGNNfkj2n1I9adwuORGZqaYz0XiQQmlpd6Up1UQTG2/SG48C2bQJfQmeOt
Q425mClxsPQsln73azizjUfGjTQKh2pMRjSJQ/0XrL3wB85dTRk8Z5xzusjLbvbWEe7nZXSEd/Yx
9jAu4YH49Cb3rMiDV9m6INkAFo41NRsjheSCZpNymK7Y3UgJl/m6+CL3R27gEcNG7JUYkN479aKx
yYlp4DqxTmJdSxc95BKQw93eODtD+eZwbh9DbxgTja8JKiRVYMN7D9V8PK2dh1r59FPoSBA9jmGr
katicEG9RXn076vq65u553N77ocpOcN1yiRfRby4H0fUnBZwd4wUwxp28PrVU0Wo/+zKE9NyGD01
8KU292+NbbQfGQVMALT1V63oHxccy/XheX+q/FvXJ1HxtICZS/wLn1lX0R1ZmfAH/w7hH8Yr0fjo
AO3u5qaWlBT+Uu10cm6DWK3DlP7cCULWRqdmhbOOxk4wKwn0gXAGoZjqlNPn4iOYD+znt8TotVR0
ZYaPHtNntxFj/eIol90Jrdo5FvZngdZOMmf5bIlqzYvzIsHRMsvd5IeK+DjKbr08CL3UofKcOaeJ
1yDLjRumxGKIMVfDYRTPYxWMwaOhJyzMUDdnyKpCCr4+4eCCs6T5WjcrbRryt1hSGudswHInetKf
X+4LFcag1rQQ2GfQexifrIwEYffI3Nu+bidTv/qYggPXOh4Kz6vyQNuTC4IlcJJltW8wNbhJgsdd
wuJsWDGBLRVQl1qiEG34/b3tYqG6sMpBbMYApW0M5Ekm52TELMFB32/0OsUQecmgieNohREi/D1F
LfiuAszbqMl/umoTU9Ty8SPUiqCBg8YrW43fhVVD5g2vAx4KPk4ZD1bUTwTC+K5v65kQ1xsXj9/M
DinZaOTtV4tFsFKFcRX1TySWk9fHxrZLx7poL/Qoelcob0bQJ/B7r78dg9r9NQ1u3YjKN7a3gICA
8QptgbemwgPnlTTijvGw/z+A9KgxjQL6pored+1u0/9RNg2ssxTCOaPXGxD8aiW77HyAw4XHqpb6
Sh7gVdCGus871cN8WT/rlOoEIj1Z5tO4JyQWvi+He6PeBwvejk/MDkUx7RmKzxhAuHl/yKxbI2o2
sCbMBFKExxjqYsXNJlVNp3PXttOr5BYoPKGStDidRc05iqhITPlAK0kEjHi1u6mCTLGWRj8XJQWr
FzOAqTP80faRFGzS243PlsZrryqBW9Vu8QTM0OAOT9XyXAYmzJzfADoC0CjSS+w1ZD6YBOTBT6Pv
3mPWNsdtovPGkalHR/BcMwDRb7rS/KWYvTaVixT2Kyy9YPP25a/QQWXJqfR5jra4w85tyh5DNY5u
9NGrAUAEPUh6OfKSbedEP9MB3xh/dlilYm/AiXT6Ep5YqEl8JYk5+FYhKiKATul0WTtt9kvgPrCS
TCaL4qfOBgdC9B6sIzvS3FXxayhKJGjIISwycnSt6JjCV+K6WvQXtLJGN/SK3Ds9k2ma4guiFSPC
WshfkU+3Y8Vl7qJpiW06QOY/Tst3JCyf5kta0eEQQ14TO4AzUNk1nV84IVCJEcBj79yDNM904Ip5
AC9ObCpuqfqo+KvbbTbG1iKynEJFckJNpBbrz5cTinX59uwm/8Dj8Lwrrd/BTN5kiilaMFXdeJYw
KDW2kun241zFICPiBUeYZodC6fnOQQl0apBT1DMTXmBWYK28RUBdm14f3R3cvhj/i5Q6fo/o7lAM
4I7FZ0rQucLcJWYtE7/6NXZhfTP9o52LjELuxjVewkc7lROO82wGkUzKyvlk2ZUxO+v9VsXnuT2K
xhcFOBgL+kFXZy1kTx8Jt22NhFWwczXTa9ddEcIZKVcnDAS9z2UD97DxOxrZXFkeNWpkiRPvSDby
cxIE3wrWGSU9WQYo4i9BfH7mSt3qAvSPg84cXxzLXh4M+iiqYDFSbFmJEZUi6NAZXqhi+pcnG/xf
PQwBVCh94gs0+/58GyPHWZHTWKUQJlhROx9b5MfjovAy8zQ3XtX2MyqipPXFepfI3mK5VkiNI3uq
cNFTpXfOF4wsaO3eUi1fcxY4AFxzBDATle/hv1FHQfkPRlSjDOw6rDfL/DqtiMYikliJn9a25jnB
J68lQKMm0gQ+RTS9QXGyFdEy6rgb1gZ8XS5OLVqWd61mqnnV6UAEBeF0MKuGyohkq0sZbhu+hF8D
ap+NGu9LQT0y9rc+jNr7cZfVw3OivPz02zlxJL56qiXicv4yQoICuBvwPhEE3VlsCPFzp4iz3Dbd
MwmvVv2YoKEcBKbjqKjrOU7vJO5dk1ScRpf0+9dJyw6MJauM0iO4PVPVVvCconvDYSrFkxVpkz84
0mdEtU8v5T7KKVFSavBOt0bEiwyOlbOiqgVFunDHkWD6R65XKNRlBC+zrxIzu5teFF20WZToeqA3
Re+dwa4hJ45HDjjwNyyd62zWytD+pEflsMv2qRWhOQcCd1Lx7XE8qGH0EEnD2T4imDSxMPvEQDvt
D1FQTfE0V4r4kZNPe4sKbA6neNftwFVKq891x5InkuCvIaNFv3H9wjQJd7Lz1YJwuzeMf/miiYN3
cuOr+RWKtobkwO7ZMGnPfivuHBT7c2Ht/Cdpj2o7B9swyWRolRz/0brPFw4t9AbqCw/XMM4e57Nx
huuU3a22eflPUfG29RJeXRet10awAywcrpPM9Bw+r6Vx1LedKYsXyiZweCr/qqrXn1N1EHjY6q+h
VQg4uTnMBckFr0XP/rNIzS/nkWz771RbF2DrHOJW5oZsATe04PvLk2goVCONpbEyRuXHSHiMs1bQ
+zGLZ9ZpI9aGy2Nl4rfcQyTB67DqOcjDlzjSkZM+dWFVOXaumQDrKKHFf7gzslkPUPsQlX/BZkhE
lMj9MtyP8tDan/40TjrdjBrq2SKAVb8ULY1qUCLUWN3Urtj787jiX2tz9WBLXnSiJd/f1a4x0q8K
ES8/aWIr5I1ScaEGDsiheHqA9y3byFdwodOSCVYVp+v3+NgrkH6z9dKaV8IdjDvcyPS9O0nmUcAv
KH9L1NQ2tDZZNq1PtGHatRP9n+c3DxdasZ0OfcG9wRNxZHIysVt+6KT4WaEGWk4qCKT8qbwL/s+B
XhLz7XkwEjCmaJiV8T0tObilY5OA97/CMUaoNxvevyrlNZfL0+RfLJ/8rArl+5kedQLSmgZjSuXX
bNYSZduYB/1kp29BJ2O9XA4FvgKqijM6KPMs3EXEddXwJPHvzJAk5HeAJRRTZWHo5F7TOvqaT740
L2efDu/48weUNPO39WmBChQnucVTgto6wCNBuxC6poZQkWT2DUGBVMqU2bgRrAXmoCfhq12eG++S
6COrVTGEeIXHHb4xZCYqG5Zp7u5aDLb4gCWjDQ+iQYUvrOa/7uaFJqikK5ydCa0P1VXf/3p5fCy0
2+k1pVGFlVqmFgZxhyhClzmbWVzvQBlTrmTvPnH6nN1rskJ/hmaNEKs3xyX6wW+QHyLi/4/yNHjD
iZgyhEWhi1qCz8dsvebEnBLoDREv3gu0rxbvXk8cOPMcQCDuiNcez8c0wolcBarPj2oB8pxG61+7
eQJVLDJc4Z7jDVW4CQFkCQ64tT6zph0O5uRF46ujVhJynWEMeU9d+x84STLZk6336GbnhoS5067Z
2idLoA6JmNaszmI5zPR56cZMDxKFmw1rnNedWksQ8kEcep5hBHRDqbH1XWgEk/U9sQqFpAbc7ja0
RbHvdbSgiKZoni0nzkJbF2UX2pAt6w9bHvjXkefXYccwhQ0K9t8miIE3keeQGt1UlvCiPtzVsmYP
iU+wWp6cYTM9p3ncZ6Wln+f2ul7lPsY5IjXJ3YgQyCpB2ivgsD5ukycD1o+ny73gOnXRnxsVqOeA
krgbMZQHvaEMtpT0Z0NJ6Fzw1uEnLY8lEWA5bxqER1wbfd5jjchUuKo97GeGTLreyemWmasd5Vbv
nOY3RTRwdw/aUQtjf6N5npoRGoH/Fz0Wfe6cWvK5EI/V2IlsrbGinEp5KbX7Bb12cPmUCovUbOAp
CCvvYOezBkwe8nDt21G5lqYW7VqH1lNAWh+YcHd59BXHUm3xpnQfzVAJoJuzc5c2XztBG5L78Xza
vu8RPkCHjx8xnTfGsFgjKlluhJkR9dee+CI1J3Q+6Oy5ZiqE2TYRaIvcSy7HiDCcH4z5t8acJSyH
PSDzOOYoiexjmayx5RIa7gnhaoIwPqZyodkcfknIi69GTHzuHvqS3qKb+S0k2v09ZQBhkEhci7O7
tE+A9ROmYodOortdZSfNbmK8O3hE4Bc/QiP7wG0dm/AwPrGRG6SY4cxtC0qayjVjzS5lYaUejuWh
JszBSxUZNWpbvjk4FnqDSNuo5A55v98877QO8Orp7t/92s+TXOHt+Pgt4TqXcdW9jy5bhY6ip52b
+Z0aU8PMz9FcZlnVNwC/pnuWLk26FD+/ZNQ747io4NO2GoyHJA9zTIV0RxcoLspnZHA32r+a8cja
G6KsWH0CBtYlB+11+LDytAy3GSMsMOeWbrmXnU6VDrC1lYW++gmBLblvAOZBM0FHHfr7enhkRO/5
8Ex6V+9YIFM7jizpuEyF9JpsyTSVv6kRUp3rNgQhO3m2eypFQlmazLENTInrDWsHbHZBy8Fx1OUM
uAYahnO25W9hznBb5YcL7fTXSTB+8QkirfHKFoPY4nk4eHxQyO7rZiPmCxZlbc0gU/bdcPTd5hFg
T+Sg6GrUylnIeCweaxGTj+xGYIYa4t1ZW3FZy1KSLmsmWI1YkoY8OR3eFdctZPmFBZ8glemT4ALf
7aOqV25OQe6Rc7HFM/pUA3FmTpDb/hvfh/WVFueQ/tAj5N6R2z5lHOfP5Mr3aAntc1fvQNVX/vBi
xTgJt1pHFDth143sG8EMrpH7GIGaUtj5q+3Q/JPhnasw4i53P+c142qiuwzQprXyFA+8q0MPQPzP
WOgSxCuEB5AYFm7JY2sxsPif3eiWolqv1fW5OrjrhIHGTFrrT1pOgDPA/h/TYs6K7Y6NWOdd3fLG
iX2fSO8eYQU0vx2Y6oReAuBxvlBMIDWCui1E/7qw9iMo9C/A+O5bkkDIlZmkj4uOIc4QgTPVv5y2
4FmUG38QXvt7T/cwg/KBRB6RYOeFrQH7Bt8sjS6I//n4/TBDb+fm8jz6BomePxg7cmo8klBLSO6r
ikpda64809kBtRjAjb4fkarj+p0UZb/q6BOvp1KYMULMkJGRiaQFEHu/iYNHmNOCzh6hyXmkklM4
G2hB6x2f6AziWI7rDUQsFT4GbJsY+Hltl+VwYDo/hw6WcDYfSku6nHjzOHxw2WezMHBvlkbf5sD4
sDpQGROorksGGW8NOkbA9J4KMOkWHN3U5OELYMAdTLLkY3wugw3/DRQQ7PVeSXjlrewK/xNdI9bA
R8avigCiSQpbzRX3k5T5h5M7e0EgXBODVqMMUFJb5Plo2EYhSjepBKV3j2sMraNAUtHnjDKdd9AR
akZJMwHsB8sc1pnL7eHcT/dUyG0+OES2dzJ5XrEuCpUCLaFHrd2I5zLzchfnL3X4106Ggyh3OnfF
vsJtOZXxIyDJ9JLm5mulH1s/qQQBHBEHG4FaqOCPE97taUkjoaueEE+WeOynzZPFEwRN8AdWV1ge
Z7B5vGxJLC9quPuTE+BrZk7Nds0aJxctJXfgzYTFNEsnLBdBm2AkXydJ+9Gdba1s0zcfwtQDIiq5
ogRqkKin++BKtO8cufDuANMnZpouC5Gs0SYcfGPt/PKrQSvFc6uF+mJtwsyhCUTf7ULIr41JxuWi
Irftvq23/N5G06nEYnn5qjInJaTdvQMUWc2pHyf9Fx27YYde91AKhjA68WCGR9OEtu39/u2/2Fb3
OdnbOt2oyQdgP6DowfEterCvuhdW3CQiF66Oj3IOAHX7zcpNq4XEGoiFD8LvzkwsQgFVBD8Dl6QE
BVr9LxaAQobwxAUhWtk9dZNn941rXCLb4ow09/qPCg8IC63mXFRsD+K20huMhXCiEIdGReGOQrMN
/BRl8+7bCuJcCrdiDr6hbmludEf0ebWPP2ntiJU8pPYgURhbPJdHGQV5wrGcKgcNI/ePWOagnIpz
EKnUAOIkhtlHue2rUhSivuwAREB8UAJItpGW0lMT75H2Jd2ElPg7kK3K9px0wzYg8h9qNLpJDkuK
48GZtiKXqLbUVK+pFycb7J9PRd5JqR5UV3/Ip0WpfWMfvt+xZ8cb3FlsSxzgPt1E68t5CBzHj/4O
5zbOrcarJCHqRlb/wUc3415Hw/prDDmPWcWjHc2Hau9PQ4hQcZt76lH8QoIzRabbe0jathPHsKG8
2HWS0N4opuCOA++wmRtKNPzizi0G8Npj2BvnY+/KZ/pUzvwx5qvESrjMYlmOFj5GzjpMN3VidDHr
htfZzOpSkARNwJDLtQVAjvY5mel4lHFFMT8XGVTCA9D6eJk0x+8WlV+pswj/9cWqRoMggbrU7KXf
nQ+LWFdJw+rws91/wDapOaH+wAB87itfY3q6RmGX/0QGUw8LDDfjVpz4IxlR1gnPMtW0IyAdcNTj
feK9q/kE/nr3SoXYk//v+gd+hAw4mYQS/RbO6BwHKSfrSXOQiowS09vJWtQExJQSg4D9zbgsqzk5
mXLAY2HycY1wCExD+ixHcG+cwATlEY2hByRk7NMFKT5v6uNAltnKjKW8xFai6PO+g2u3o+76b1eK
1FZ93Isn8ZSBNk/Mi7LSL4sM7mcWTxDJALPkO01gFQ5X72s2u3i40WPOtNN9XMCC6EFuUzMylWx+
qqin3qYnvyb5/o4kJDmj4WSGJ1bIGnlMIPPoEQ76AoKrfBJjEEyPSFFclnll+Rs8NsMWThK/ZIEN
DepOu/IRoY85/PYzfeigy4hTZufoKo82/eJEA/N5rVEqNocMCXgcoREmV+DTCxPgcDZ8sUoBVSV7
6EgI71E45kUKwYot0mGYNGvdnzqc4CjD/wNzpp6Z1sZXaPS/EMWXEv0Q0z2ei5IE9vL63QIddFc6
8LgDgqKMnpFvvrKyBwT16MEJjqw58ER9c/5DQ5yVlZOVxk5mOWzatMzjx9HlO1g4c5LDaXdqsAhM
DgRn1/EJ0LYcCAqM+bFkKcJEyS1gYNLcfDsZ6lgqy7rMDouRnhLopyUmTcCfK5vBkmyOZWKZPe2V
F6emFzBpQNLFuvJ8xh26idEIfTHVYcGQufcU0roJXssnaP+vbJj1F6F4nzuQiU5MPMGOvrYyjIco
RpeTvnml40rTWBW/x5VRNiZ+NvxZZ7ynSZazoi+1fEs41uDetUCJjc70L8k9qRr5eLGW57N/73r7
HmTZ6beAyxWGPav+EZyX3hVFGT5gC1AyETOprUUDQQQOUmyYtZHLViuCrztePkmWHRRTr3GUDqpz
1Ve3xT27+L7SRl5i+ZcN88OqLL2oKT5gos8QFHPRd+6tUglUboMy/SxqYq4JtRd+dgxlPphrTUSV
dTy50rn2uZTJ2zcpGTINJZpzHghXpW+WQyZ1kjfdDD2Odxz/wMEnl9qxzWOaegx8QB6nC0M7z8Ek
7pu5Ca1Ul6mEVnFu2OwCxlwWqJFCzAYgEAIQINu7hLwUbBiGgz67qMJJ3q3J/bzRc+bcSKNDHXtE
xdQ6SAaA+a8wGoxR8VTa5ovTFgGVrNJYCrPm8bp+OIr/MDGMLV2ltPH+Rl30E7XRmCwCYYaBBNRL
NXkfFDhS1hLSQgBRe3EkxGEcedwaR9Arv8d/f5BpAr6LysFh9PTR5ZJx09SrdhvO2HydvoU27SJc
IjanZu2V4dORovwcYTcWBqHB3SWJlP4JedOiNQbQhflvV5/bl9dGUvMkBogJr4uWwcNPkFYOTe0z
SW7eKiQTI+uJPd8izpVAzaadrpc2+j5luLYaJ/G+wBorZqjBOFd6l/BfphGpp9zZiZDyPLbB1srz
7oFOr/1KYYzG/Atmdlw6ev4H51x4wqeODPZzDOOWNelWxnRoyR/5GaOr0PTdGUKu0gkizbjBa8A0
yRkt9SgEXnbX0JHBGFz5sDZ9xKGi3Goi0rWg0FBzxcx4C67o3fupyStxuFwrfVfmW1OnPWayQqat
YWhKq0UllS45hdrh62zcDCe4sO3VCP1wIqNRWpnEKi3ALg6zmsJ+zFzKki3dzDob/XOsb+x+QNvT
oGZ/R4ZlTCpegZZiwl/xp7wJ4bxY+4Ym5MMBhp5RvtTCltnbAFcna0aEq2SLckYsXiWp2v/0vuwN
xohFvsY1fHqHq/6yI0JEeiIB5TZZPHf/aYAEz9e8WOKaADT0Pd5k16pIwjupW9FkTAXiMPpqAG8h
8/IvkRa8X2xTNOjqSydajkn9TRJ9tdXp8yXzxLPOreo2Bm4qdP89Z8mtaixoFCmwxrJzIAi4Bsxz
n6srM3Zxhbf7L3IZWH+ol4b07mhSBepIz2L/KzHCdDC6ZSJ+VQVB4680ojQZFZTpYeNqDQr8z9od
dOb2gZ4Wo055Zmv8yRm3WuOpp4sPzSKsL7V4cg/oIsE3binSVw7siW9GPuw5AVYGW8acD1OM0fOq
6iOoxjHCBVuyAit6fWpa4CO61z1pvOqLeDQw0mJdD3vup6t8QH4yBZqD/doAHVPEuE5yzgYkFT5h
9RL2ZaEI2X6j1uA/5tv4t6nX+ABMSTElpDV42CJ0jYqju5VwPLLGVvyssAtcho0s6D5ZeN4mZYB5
+xknSHepIHU+8yzAcN3rfs2jj/Uu7NKw+dAxgjMQMJry/IGkLgo1oxmocwGJoSDHwhY9QprdG4PX
R0gBdDJvbcUqwJTBG5WaYipNR9vRHGT9r+uhFqkL6TKbNZ3YQbOWvj7FbJR8RfEE1AwMCyZjapzd
ESGw/bzWekLP38S8Zi7el/TVK6I/Vytt/Oc2avRCSaPEJZVjaftE+2vzcfuobb1tsMNQDqGvcHor
V+8Ws3cC9CAf/iPJcW11UpkEvJoMpgj/EAaYj9Av2iHoo4086SXRvtYweF4vAb5PyoLmiijZwiSp
yd7fdJ7YItXAjLCMtj1ZWMVrbUEVjWDimI43UCedZ40HzWNo1ljXkYg8xRX3EdlLb3kqLFFknhJg
7ekc4j/20q8a0e5P7J1l6IhvrECIXh8hgQkKBeXzXE/4a33qc4AuAgyDeVwOwtRwARgtuGtKZMfH
rQtw+rxfbq4ta1pwiFZo4gie+Q68jHxc3vIplo+0SmPU33yUV6cHEBFPetceUiZ2zJJSoKEXW0ZL
u0+706ELAjwVzAF8eGQKAd5e/omSD+l80LTC2HuDlbQ7BRtDtujVt66ajj4O7J6TrLphF+khk1xj
aCpI31b5P+29611P6p+to3uljWilMyRd9VAkaQUN8z02JgZXdkMKg5omTT/J5NDBykyKCaZ2tiwc
7iuY/2CvAIMCejXRr+503zNpuOFYDX78vzMb5RHOFdj4Uua1srD2I5Nso/HR5lVdfXxZcKMiq9R5
V3xcfnZwqIh8dXRTVX8Xyri+EOJHoyIFvOoNd3/aSeK7Ek2gicNuWuGbzqkSmcrRwamAasw9wzbd
kGwBi9yzlpGjr6LYaVLTAFA/GXPDz7fbHL5B3pA/iMPtV2Abo24YYuvND0qvDVyFKk8T2Plzm2EH
u/CLbeJ4YIVqg+CsMPyxwo71CP6naqqLzxEzdh2BgK8IbfZHOqbOickMlxhxoZ1ms8j/0DZXo2bn
nQrpHqQCwxHGst6mjWoCQfFB+gNk2zPZ98V2p3tPeCTbLlcBVTuq5UtKfuSnaR4wovupWSBMkf/F
6c4S5UEWv2ZmEgF6S6HEJyrqMPAsroIojd3BOO0wTdgL6ZgeDn8mbZP6POGbtmYaN9A67m+wHrwM
9UhInKTDwEpO7FCc4h9IUEPd73FPldiYqtc3Bq1n/ETm4JrckhxKTzHjFlVNNlmpm07v/LEDkwPk
LV28X9mES1iupVc3xl2RYCaoZzLi1pieh7A3dZpgQ7cPfRGpFywBnVvncsnbP/VO26a1XW2cd5Po
qXIgY571nbpM/6UHVZVqP8y3DgkuqTpM/kk/UHiWmhcSRdAEJVW+NhikGT4RENrq6QAmNH0qapug
PoE8OXiwAT62muh/PnZTjm1kKo4YLJtOLzahqe4Q+8r9LAw+2vP7cOxRZTHpG+r0tYrV9/0oMZMq
TxuMV4Xf/CUXkWVv9otoMH8XGvwf9wvfE4kINz3wuLdV+iSponw+D9bhQdqySqrj42qo+UHTb/ZX
HujEpie3pHuJHkqsLAEM8AJbxRc/i72i3jdCERgVzOeiPmQMkPUjCXQeN0wOIWSAKVl3FXnoE75d
H6AEg56Qw2+vOcTu/2/ix+OhgPsWJRUfwrPTyVk1fP4REPyy2jVv/QDca01rmcO/HAd0JChDq+uX
MT7PHQB2fbCfeSMR0bDpU0Yy6C4ckNyMfvKbDK5zCg5I5GqC4+HV6LvnXDIp7j0JmHFRvUHSg42T
v5fH/1vURIx1DVbQX6kEbbhMNeEYY2H6M1uw/tZ+W1DXRgbgoqQQFalqbz+ZEgFi/95s9b+KeRGO
T2YLYzP71Gnrt1jjvXBKBsXyz+7z44NKZqRZixTnwuqCQUzkji/xbwXxTQcrGJSCDxj8dqIQ4/bD
VgG+wDbTxlzx/hkVkZilE6qIQhN6EUMRtksiOemg27hzRCVMVY9mDOr9UoLfL9i5K461gZWbgcrh
QIk2MRlH+8pX8kCBiEXrL6VOItmyhJq3aHUWx58a4t+wx6dk3n/ZQ7vgHEXw6nqmLuDVdk5coikY
mBuU7PQV1EJjx+ialgFcgXqDrBfr8Wb3QLNVz9wLt8OJlJPnCaGYOvY9taXFEPun3l1+z15WjbZN
4EclFHrMm5CRyXOHZGaYYTK9AwoxdMOmA9E5/5G0XQGOAMgcItIQCShgJ6j6Y0FFeOJRwCqKTltv
AclZFrV1afUadDOCi9gUQ4azhjETq5xvGwySwnPmstVN/boPxqazwkAyQsWYWs7EoqUWnItacvop
P9u9YP1BCXb8CNn2TXFFBxGyDFTM4GKjpETfQzIAiNN9Upphei4zCFyrYdao2aIaa839PVAe/Y63
w72jIcrC/VrLT7obyoPr1uTt+CTJVdB4ucNLXhEGmXZuKH7IdoQbPnvO0DrUVuJ2uEB+Gud3Yk7U
UFTpBuZda7NwOeLSfA1OewMdOBqutWHpihYGg6h8OcY20tSUWu8ne6q0q5thx+qzFAndDsCGRVPp
8lrJnjlLtVPC4IC+3fZ+++15A+P3XYY82LphBmEl3wzBQTaI+USUL+SGrnq6scD6/WBse78x3qeS
tV+r9Cv2uFAZo1KGgf7pEVjyi3lyjVbxIJcfQg8Ar1L2n399iZIq9sQ3M0NQ9YwxbuKtoowaU8sq
P9uiykeuDo9bSFZsBqkjMW5pLvsxtUFAx6+XIZ9/5tIi2jFvTyYdCA+IQmWFFRFRrLyVPnyUBRwn
aBx2TUDY+bZopQ0T2xzramq8WiZ9UQzqt6xXsuRmhO0lHpjU5OY25BEZSDOeE6m+owbUd8rj85iM
R415dIU9cEG31JUMsdJDnAvbIfFmB951uBvDjT5p7mXdGAnt5PJTA1q4sd0CQjH/e3hJE5PT7417
r3FvESxnPQsSqgs2C8tb0+HnLgOeP/bVo6wfXLRslQ4z8KpElwmXstGUU7UROFiOqxRYik/R9FuG
8HHsNDuY+rUnx1/4DI5ZlX5RLcJTuYRmwROdc1Bnb/qyw8ZY/7QEIvdIqx0DL8n7zNjkNWmJQRn1
ViejtuoqBHInfaPiMjQGzqZLBjop1QIRdcRi6O7YYIQB+oyVPKCGypYU0iS4olgnCYxKHOHtHj0R
1cHiYc+Td2AVdEkCaQC7TI6aEbbGsdH4DlpoQJ5sXTMSOZ8D0puVbtDY/qR1ChlwYw85mQnM0ROq
6qLHDyYLD17yxejpZcC1szrA9fMxcdQWIJ+bjDMD2r34qty5aFyGig9GRtsbkhW8EWTaNMx72ypk
DZI7WlDaGNLIvJDcPGuIa5C+RnfFE9iDboSVlbrK0oYxr8urqX06WW/4aw/bCof4++2i4ZNWxttD
PF+B4mxXw7vVjjx5gxaB/5vneY/K7FmJ7lcVBVb75rZC7TUSu0q97jsvKfh+rRKDBUB0XnUkI6G/
Jn5kKmJBQEeQnJWI7/qBAx3+UbOeEp8pLuORNP1vKafVAZcsMJWK+SZIsMN0aUCeHKrLxRpLFLEU
1wtW+mpfaLUQT5SIKiXFDxiKKIR9BqFHGBBPReiJvwIBUbEGWAop06aGBYr3nh7Y5zfB9afZWyLL
9+Yq3y4lwEphu6pb+eXBcjHjyucgIaQMVuLnp7+pPSSUmmnVA+K/qWeib0etmZv/dEakW63T0FEx
lYIILZ2gtIoGXFlUVmQQL2SiKkmDARaEZBwSSh5Hge82IyAZbn+oBFrmiScdlUJQRZfB4u0wGEc4
/nnz2QTMGHWExb423tLaiWlap8GHUgSazvAUgwpX82abLxW8nqss2Pf5AoECuKzXVtnEWHOJiS+Y
+W/PWEdDdZQk8z9D5Gru/zYD0VL9lTckOdrdoONL2Bhb8ZAQ43dyeZwlv4455LIGK/5ZGU/k3Q5y
ab1aRmkQAn24ypADml7I8bXg8A2WZcNzjTey8HM2Ll8TCETtE7UuaUN+W3SDK2zaNCpSakXBUpVt
BFCkTX9uCi7NkL3oVtFg2y1Vq2AuKAQSSEIHCgx0OLYwZxoP0lL+G08i3Mr4FpxB4pFeuASJvYWc
Szb3LL0IvJVY4k1ihsMG0NnrVgI34vqIatGfu0v48AK/BR4MYz+mDLR9GznLptB9Ajefz1HjsMRJ
qZ0oRVE68Ymr2qQcE8uqtioVqLyJzC4xNunZ4ItS8bPRBVyvInpGFmwfGPJinNTenM+3W4eAdCA8
wfdga+gAikxZRAhAEevs4C8n4SBoZEFG7piG4xG2VEEoezKzEXE7ZwYYFgQEKOUsSutLSeHqsjsI
XHdLlozXQnfykCj8PwUSeLgplW1N2BAe0S8ZLNqtkk3ySxgPXnf7HzKzUdngJENkVj5JjTcSYWBU
S/pX1JTs4BqgfI3ZmYsp/Z44qR/Db1zV1w3oIMkR3usAYl+hLIOUtSPOCsg2xfQm3qt/c1+exeap
zl2bg3HnWNIRfdvQZ3pz+HeK8jddjJ4Jblyk8CZgd4+ZtJ/2SxT4y5xzD1tHRg+O18xJp2ZA9QQp
9+qx+6MJS4WnRGeUbujY7w2bGLqVvl57ZwccCXiDYJZLwVemW0uYO878XNjrNx1eMa5/fVZuZ6eV
EQbmwkaPqf8z+GJt3RIoDLzgAny/y5DEAicbAOIK0cKUjUh/ZIuCgwyVL+zsIChg2sBnpdvDEZDS
k9BC/lvn9bKDkBYVhKEobRs+wOSzjWJ6+PcviF1uTn3MhFYkicDnflCTU0qBEVmS+FYgPFPgs2l6
Y6+ouxnyXD6Qk7xFEJ1hxU6dgiM26krlj6Evf4h7byhUO5mtBsnhaRM74iI3nSmf+SndDYCHAIj4
iZgKWEjfgyBOSRqEt6S+46JCjUF2aJuQVhBUp20pt+t7hs2dTvacAmgb9vrGcYB4UR17oVJ6Rn5I
QdEmXT7rSiWbJyoBrm07exgNDy2PKhbmcve2h1u24FntY1aVWU0671cNfXV5K/uuzpzfFUKge/5f
s7++29i/N5Qqg12RTGAyakX4fri8Oj0KjGNxZSFYlu+1DEhN/ihAtjKntupBpjs902P53Ao4Komb
2MxbJiFz2dnnMPjb/xXHM9Qk31JYCnHWahNDf3RU0t86icH23tBLVKSWFlXahHy7GsqssjnTNAPh
AzslkauoEWUNf0tA/50GGBoNUX2ZSGhTj9DVeM+XMvwo2lNfDZBU7SZ97n906bVWfu5D7hnNy55z
cC+liGmV+A/j3xHIv1yLcDpOsLq/RQ8H8WFwqV5lQdSi99VusXcQGyjg4kA5+NuTm9yoS9704sIL
52l1V/WowZfNM+3l9fKUoKK2LSor/q61az11FMMf3VPXDkojVZm7RCO8DoVvalwrJ/ZuB+ZtkLO7
8fJHKYNENeW49TjBJDNzOHvK8OmxEHi6WiQltKXcSknQgLdkOejNc43lft7h+gAhU6g7G1DOQzfc
6aZVfUtpOiNiawBfeAueARTRBDD+DSNYl8+Dh2Y/EkFvibokRznFhMO0SNFQyimZzoUmyEzTIUDM
VI19ZtBJmSvn/prE+cZHEHx75enVE+0g9veYCwtd2I+QLZV5zMKHz05KxGP6SlrwEadz9FDAAFDR
z1M2cz9M2Jd7xYWZ7Bnz8zXybDqC0rhz0inirMTcDcbUW5pvke4A08WGc7Tct/NrT3cCvfPtKYGi
FSzbT4+5k5kHOHzN4F306j0qNz+Ul/4bzEMQNWGbhhPuJUEROK9VL45VTDXwCE1SAGeLEs4fOWX7
8qu4UiZCFdMa8C0kEJaL4ETuyfk/9DyXgG+3HLatEnpBaT4AQsWqJMYigUt3QqKWVkTJ3WM8nQtZ
MjOR+hph80AmoyOQ/QR1LAoKeluDcXV6FSV3VNM/nCBicJNZ+OLu+KMvUStqTPp1KFUEWXOS7POw
T3v+KD6eGkdMW7snrOYiH61Id7fe7Uad6jqknLP6S29IAjDkG5H+t5pSHMq2KiCsFjRn35m+rsJb
i5E51x6YED9IJ07WjkvNRbvsyHJzPwI4Oh0aMBSAwcu+sSDMMa8xilEN3WiMKpzZ/5RlPf+vISmO
wfcgX2cKljzJyPr/udrMM+2CBSRDjid61P6wY8ktfjnETZshFJnImhPje+2AtnxywbgN3UOZjLRz
59XZGbmhYyC6hbO89X9gXPUanhBxkWRDKHUUzQINWXV1zQi9YRPkaP8OLz2Y4wik65xY17bmim2e
oI4vlhdSO3gOI4QsQ5Nb5xhUtnXJB3EUg1dRNwDDR5GRJJC+sXOjnsQOWKF53OH1rfD4P1+xru39
bzp+CXBnl7BU495bq+t3BJDRsUtdQISpQaZUyvK09nq+KULZvZp/9NM01coDqstlzCD5BB7S3y77
GcWIArkzw4tljo6cf+89798O+tHmFtlpkCW0RNiAim2RXoKqyjdlYb0MMtGhHozezQhox6kX8Gw3
03+aD5Rt1LxkuPSJKW0M6bPLjDzO7C8SFv4h7QgaCYa6AP0W0iKXFmR7/fXqcQmXVcq5l07L2v5D
U/zozPr3M6iZXYre5v8tOBiDnwv8qkf7boiePAzfmFxT05wHEVTlQMjKnQ1MtViLi/MfeTm2x7yM
TlFwXbryn4si1K80rek4UCJNXK5TLDALIKb0T+eCcSE3GtJUALXv0PY0dEzrUC48J8haTZ3ZLKBI
9/XQV5VsFvh8zC9nq2PMRyTa+IINVswu1qQUStEQ1K0vC6/z68LTrpx7JSMNECXUHXLjBn/C6cZS
YuQaC3ICzlvwNCZuoTRYwIxgLIUDuZNmH7tdT7b4wR/QSNxgVVM2+ckAtT0LGaJq7GmkqKy4eB9v
xKb6kxXJGkt2H9IxlEK+7Kz2iSvhHwSSzzt2wTr5Urlx65m72xeWHj+Ls/0WzeowujtJ1xUG8xo1
e4JdP2oMgr+l+8tcOW0EHTsc9Mf0Ex3cc0TFd9+M1OY4D97eAFnrFYLGR8HrUms+Fain7FcuoP8m
am4rZ7YmbDbkKe2RRZxsXAx2ZJiJOsULfcO3JDNjeZxAeA6X8y4cpOjH5GEygMg9Ml4icJSMzS6u
YSEQsjhERARl8PGWvs3/gn8nh6uu83oVoV6d7FSVkWi+MS+wazxT5jLKkh1PmCmlrDF0YXL/MUXc
tG8nKzoNlliJD97z0bHdGjHgTsCaxUIa0hAaG2rvdpsnuEW7o42LJL1bUTqwnM92nOCWAIofOMOA
SntJDWXiSlhKKyAbB+Gdn+MGK+ms64jfvq3XwviTpNNk/QQh921lDWiyIrW3BvpYVhPdVXnH3yoV
B5hiw1hwGsT65O2rvU4YWRUCOnza7HLxGaPm8lcgcA1WB5qmtHDoS2oWsOYNg/xd7ixm1z1qVHTo
c/VXOLEinn+muevRgYoy1BnQYPey2WgC6eqY7KV2TpWFjkT2KUnKag7iwsBfWlYKhN/G8g3+wy6v
hpCp5X/9FjE+cUoVJvIffQ3ZvAixPQjsHkF28iHD+dVr2t+0/9n07I3yMYotRal8++88HwlCJERc
Die+5RjDCgm7WNmj24g0wSdXeLxzQ2WgSooYajU+YZ3PPBEjwxcbAE8/e3Yhw0Ob/7WYNIkLBeIz
QnkFrFLtJebKj36POO7D/ZtBNnLD5vPRgtbgc8Ta2FSFKMc6SGJaQ7/lJweMfKVLcJ0IiQvwb+w7
nu4cFiwomWaMrmF8aiJcMTV7DeV++NmJuIwFdiHzgtW31APZzjIPefHtSoOmwe/UDwHwpR55/GUW
36JjqA1is6glS7Z8BrxvtMd+p+fPmcG8iAlZgugWrGwYIA+H3dc14o0hZD91EoWWf5ngycj4YYEK
ZEljhywqXgA5QVEk9tyBYMsmznNkmWF2Ewn23pULj5QRbcwNQgGU7OSysuYUYCdLPm/50dukXV8S
RbDxa331MxiG1zb5fct6cQOKwWs5pYgrRstw3cbnRyc0ahkxLSN/FfVvlyMjYJk2IX2q9NnlQI0r
QCsTAC8i5L3LguliMWhWFZIS6SgbPL5A41zAI6xiBUPmOLycS4OR0WKRWMJfUZkLi3dS+p28Nr/C
F6JARZudygY2+yYgCZ3HVLP59zbzLaT23KL+YQbcumMYaVWb2Y21xOhzwaONiYWODpyukH+YdRG7
6XVSs31lqqkgRP/yZizsiqUwznjSlvp9NZoqDGMIdJltBPeEsGCqny4G60/UIVfn7yWujBlly3q9
pB5hsBTp+jxinzoIxEPz9pqsQ8sMbqsd3GXtVifTi9+uKi0SInF4TGQd5CEQTK2KTS76ixqY7xSD
8Oot0OIdjYiDg/LAyDKGpHgMNo4klQFdVu5BuwFe662dq34Bghe4LpDTrakMGYofYPkg2NJE3wmt
kSgUHo0kh+XP1gYMvyEVNGuwH2rvEf8KS1Vxo9ecrZMOZT2uFYkLosOKx/VwBAqT2UfBwVsRm8PF
GSdD7e7Bv+FcwrBsXFWhGtay8xhozH6ZoVJYfpZlrvIdvFk9fjnU82Ux6TEZcxZ6LQQeVtVSdfXd
r363o1VHMtnmNWo823JQTGe6MoJABlu+fFhzaK/YOkaVP5mWYZaPYhwSN/i01qHeWpUEzYJTPRnR
j+OLj91D77f9aTIR6b1lxXspqiISF9LxTafuvc3MpJ+acg4e44d6Gt6MiIzwmG25LL1XGEZjLWPc
Znfn99aUPJnOmmnj0XM6rFymaF5DqnNukfmjMqJgLPfBQOU7hOSLINXpfRFFiB7Kkduz2WbFWJTi
2tA+vbV8iicI2O5UymuDXRrqSgfkRCw9anOg6IK9GGzVGZDHOFgE45deqAoz5F//kbYveGjrkE39
uOkAkkr4rQXWoVFoX6JlHbA9AGvOFf0aHTG09uWMo6F8c7lGWYPjUtXZlqy86R7WPzv1qwEUcPp0
LCScStOEmIGoGlQza4/C7DarjfeWoIN7DhFfd3WGrIVh109veNbTIdKT29ACjSwcmZOCOVPqmEww
ogjn+UEZWedma1yxq2rjrhVnUJLVXtOKhMqjVBPk+goGTHFWNr7lgT4Z+ed8joqgJP1O6I8R64vz
ZSahNUsxpMrSK1y/tJDmIlvznRS95PujsXx5ZQqaHFzjfoK+dmz/Ddo1cdA5GnwZl8r4NVMsx8+t
cpCNYH1A/7kSR2FivMQSEz4NuIa12guo2lNYAp7hdIWpZUMnXtyvKz/MuOp/yG4wAaX4huieP9ic
0/nNRAxxZ6pKFLLQ+9dy3v+vTuRGoW1huuRhv7s7JB8JDX+RFjK7QtVOrUuqwsgsPuienHaR5byB
DewJ1WKO7wA60R4ZQ65ShcG8MZ0q8Mnz1BHUpg5QlE6MBSum8ATXjP3PJeuwNyK9LjDXJCBRegJy
gG03A94aHhwsB3ArSwatf3rgMgvoW1BcqNwETeCdUgee2WXJ2d5ZOm337FLs+kCULdTB4cifGzq8
bc27mpz0CUBUcnlaZFyWQO+to33uE+QudWrua+iWmUZORBwa3WP3Sp0euY3leMIE7mwpqyXqwfpW
C9BEHNjGKc+10LQ2yhQLUkk3rBbQtO6cFRBwEfp11M2uX+iWZOtSdebOFrhgyynJ8XqKEy020hUl
3H8I8TD26HOt3y6HmpKYRcxoFzAAMzW1M1P9bjy33O9+G/e6AezyfO84SWAqtrrJtGHSx4w+n8sW
ETaEHFtuSYz/Fsxm/2QCckzri9DBcJnurobm9nvulCzdoSvsxq1a4G6awHwgowbSEknbZK4gMJvg
Rxoo/loJ4v6hzCSXD+ApGCqawd6pGULI7FWwsFuK4rkpGZqCQ8Q3bjBf3L9Pc+w3/zXBFYmXO3nY
k5u/LS//VHjCVLv0uiQQHJnHcjZHStRXuPQ/1fO8OVczeiPflbKQHjUzTfHhZjjDxvkwarr17TAq
WszTRvP70/PQrO8e4vGWCysFIJ6IJnu00WkbUI2TTCLYFiJW8F2WzQ7B2iRYr4xPF4QrXt0v+M1A
bnY8sBDTiP45of9y/vh4pQAfTua+fp45wOCtVyFBG7d++z6152AE/GOIK6ewG6daSXGVCgD69m7A
LDen2w6Hz4RvIRFg67yrWKSCjZ4Gvtv3aoI33RcLxqOSAysILOKKOirQsvJpkIJN3e563IMIef1K
AEMB8T55Mmhfeftw3TYMfc13qMWGA030CRhYx89JBFcQYQvFr9TPDenaejlG3usNAnN+woCss5JK
jj7vIGPo8/6QQCE9KcAdR4KSz+ukltmSUR2Wm/ntvnM6j4Y5j0p8KkOlNW99vNicO8cjqgvMiyGJ
2hZ9KhK6KkwdA99Vi+ixMqikF/SrWFIut77WZv70AvZRlxZ+UCtYMyLyVuQTFTYmIhJUigMAmnp3
gK4haRjk5E9Xy4r6L/aC8U2sFZ3gtA9ocZD5o7uho2bpkm7y7FR73F8EAkxPdO3vJoIYDURS+unU
fPfdi+3/7DHC+zyJEpU8HDUKladsucrN5OCz0AKDhs4Udpee3ApbwSroPA4BBUbb7roeDEVJLEBJ
PoMGpW/+M7BnPWE/+Xk+iWZmguScflixtds3KOilmuCnIo1rj3IwAxSXNtHrM6Yxg7edL9Rt1yo+
n8OlgYys0vEmjxopsEVb8mB9eRqO1eIZvrnn3dIAWiZimHJWgmpnDAbEs/jGcmDn1Kvr1uabH+uf
bOaTArCqrsdBuTIoCZgDlBtS8xsVCeUQsUcyX8sp9HR1whSb330f+qOZo3BDzFK+eZCf4JDWqfGh
eHNq/0djon4aBoa3VOU2LvcIis9hRdKZPU5qf+5acHVfi9rCvTg9jnaXk9s6Q7nQgs0ZfDE4KC99
FJtiYetdf6F+YPId+47s5/jhyX11fMNnvPyoJRGVlNhe2TJq3+RRaVzYkaGT6XPhBojKxKUhJ0Dw
HO17GZka0isKigcs8NxHwH1qP9itT8ZJFOkZK3oJLBR9uNkfEWD35OONxiQrrC5QzW0enyoLEuH4
LaVss64aUpyTBbGAyJPEvrawRJmzsjNdYWbPNle7F3VVeOPczWVabTyLTyV2UqhnoE/FNRmb0uvM
6sBh5SLFzYMby2GCPX9KgtYdiVzbNCP1YdhfbgflWlhip9En4LeXh1V2UpdYqYp1WtIZdCCNpEXz
pgqDufxrksJ+n1/OQfb0fvSKb9likl6xX51LeUjtUA6J2J6zXHvu3dchwuRF45Z4dCeE5D6casNP
0XsQh8y4uQfDB122XuVe4DYYkdqZGshj6i3JIb4ayR6Q0eFnTa2b1QHiUS77prqSATRg7iKuUjtP
mZaQRuAGZXEsIcXNRd7TCH8XmF0FGtocgCc6HcQ1wFZSn3R/dGORpNTzhunBPPUgxnq0FGMqYcGj
xZw+VCmnG3wCkvjXVRupKgU5gM5gLgwaer+vBItfxKDWMyS2G9nIa2+cBblUabPuPZCr+1b2IAA6
iIt+eMZAdTfFfWlzHurcqTt+pO7FajzD6LHtAb9vGMEUj8xQTLq8YC+rK/ydLAgPq8Dw8y0yduHk
AAOsB1fbDmuN+sMd1k4/uBxf29yguf+Qg7ww1ICGO64z/DR9QHSJ62UK9IZekRFHvJRGi4+6tP21
uKcC8O5spGIs0wMQKuPc6KszgfY+U5YokIwroQwR/GQMrrhDeEc2xtlgjWey3NAJJo3u8HbAIPMb
z5dmS7iXwHSG+ivP9+rsN/K96yuyEtarF9ZmtV+4+XYxXQFRgsDmKDguh2ew/9gUOZx9kKIRNnR8
SejoEivqempmrvBTzi3bpoPYlKqXnrwdy2xDLIjOrtiXrBxIAmM1xcICnW1lQklDTgvF4wRY2nLJ
kID2cwkrer5r+Umhek8OdQSq7tSc1TYc95YKYgbZq5o0KZRfH4sS2yH4oHQjjVeuU0qvxOUprrv5
yOXy79iCLWoLn+74qQAzTlgRJq4M2eBP9QYeB1oY/uRxgfifVRjriIif36fk7rYiJaRXdt5NXo7g
sziHYu5hD5FMD+Kg/Soi0KA345Fa/L4vhsyJD5fiEAJplEm/xs5Oy92KIm+1E+r7J/SPCRNGT7c5
LbZJwvvoAOo45udNoGdnLuuIJkZ95fJVokQHMauekPXlCM3QYY9EyRAyx6ysGYWK4jzFiuLPSxcH
i/5JKlFpssR12tg5sw16AP67AlydEIgy1qFxwmAY9xgERX3AcTuOyCPLg4pREZyx6LOtHSctGIno
8NJ4Ap0equU090D/drbIqaQjku+W8/syvhqTeNqH1pyMsanymTd9mN5SItJ75YnHnPjQGvZwEBeq
K+Gmn2XeWvQQgGT3F6WabhNy4ObgWS0r5grwF/9/Rt64Va++tihH5Ku58sKkbldHVV7OhVSZn//F
OoUW1hdG9mnWmlMtOarUWkBANRbrZis3wcMT4hfZ7gizYCfT3TdHVkMBIdtHea1gov/LoEMBnMf2
gE9NMI+gde6Z42zeCZ7owWx1PTlckaOk8/vKvvgLTIa3G0EA0Fvx/RkpsatnCnFbzIg/DdYAWMDr
qubKMiq3T1qOqmzMtSaF1no2dyy6UFQFry3fW+RcMSNPFDSkNbZxiQ+S4UnCWZgYheRLSWiYqg3K
+HhW5S2i4gY1nfjndf84kZ3nzb6efeCP5ZTIslCDQhyC09rqhx66la/JuBzIrjJrm0VrLRe9ClKA
wTQBy52QT1NwgJLUvUhDvzhIhwcvWWGAZ7yRXaC3zYaxmAzSg8rdn2auSmRzwVXULFC8VXOlfHzf
JQ+xwSfuaZY0Cayj4zUkjyGa/UeWRUlUK8owCcTCZhwZzqe6UHbConRw8WIuR8jbblHDn+r3sXx0
zpJhwm4NDc4/Krm4QaEDhTMhnC5nKYfzcw1N5FyTQWEu+fR8yb6VTgUMcdc0teNlWxmsjzPmL03p
rxwzNWyWjy1n/p50BEueLv9RxZ+BEBkFZlFqVC54RxuXs9kSgTr5NfpsZHmYS6PDC1If5gYviID5
fqXFATT32iMANk4EHisauuIJZyAB49ycGHDWdZQcavvP50yMKcotpkTeAWkFZ30b8Cex6LE35iwP
aKxLof6YAs4uD+PuOM/d2tGzQr7qHdekF42Pbj2+e5G59Ayz13I+MjyMnjSR5RqMRPnqaJz/+/m8
TDoYa650rklsftPAJ3NnXDOv/+Euwi0fCPtgf8xVvO6j/r+FdbzGqyOnzeKRBT32ldRWQX64UNlv
fzpy9MjAdbzIvmrMpq+leDI7dAuSY5HBNY25/kvL4zYVjtW259oE8Roq95O59HBs46TzX1W4Fcvm
6h8mKUsqX5MT07bnHe6SQm8yG1CjQaS2aI2i4aFCGaN40JdwrwB9sOs8dni5PJdVAdExTvhzlfQf
+4yrC5ksU66yZVKE+ZW4JxHOErjC89BNaaCXWYg6W8UoNkBomw+qxXC9SM0qWSPemyoRu/o238Lg
sHTmQUKfrHLnOx7RMXU2UF2ZcXsefz/RazoyOR//Vvhb0JYvfg7LOHwVRHeVbM3VF8chiuAakdhW
zIkMtqLMxJPXRn+UEAbYqYmenioCzbToA4ZOAizSfX2VbeSiIIjv+Aq0II0iOJfkCe5PPcSDgToZ
dmBSIe5rfnNLiV1waZbR1ocfS04AS7NGs1VnZeJZdIsjt3+hfnH7ELTuL6h5weOmVWMqH+0eg0MI
DRsZBCJVXttdWFosIWSUGyRlv49NKn08Ca4etBo8h8d6ok/RYA2Lt4UNx8lRu31Lsb35AlR8MRsZ
IC5wcwb2WZHOKsHCUeepnxSG/bfbt4u048MQWJUwOjskOteX8OiDIeBbCB0gf6MATUhOp7ou0C3p
jEWmCs+CO6c5ru6YV1vgHxm/a3lAqjzsFK3B2vZABIXgQv4BBk3eJ0qg80rVMOk/98uJUA4PzyDQ
EbnFoGjusfHWJN7u/0xOKsttvj9hAGtNJp4OWn65/uUt1XnSTuu+SYr/b5OmLnHZCeMPDhFNOGtE
ncL8ZlEp0qf96j/jvhdtI6GreTarwQ0EZQ1l1RcWCoY3bJtefq0tQ45R/DCY4sFDHHwnl/0iuUiE
UeSq7xpSe5BTzTtz3J9Ez5TY9bmE+SfjUB8XD8BllNJIvLI16gvYa82L/0++iCdN5FfBxDP4F6U7
iqc97dVVs+zJztdTWCGxKU76Bpcj8iGsUZFyzTZAIhQl+RW6urKbhKN+MJD0Mf0OXOAd75FiWec1
wh8Ca1P1GXWollTvpFgt+joNt2hmx2/GPXxQn+5XPj0pl753tzlnDQDW7fetmJ2X1RUgYpK/0o/g
MgdiNZpyhgY5+RheRKH0s/VWPteHYSi4xhBkID9OJkOJbR39/IPooK7RpfwXpDkNM3dgFesIzPPK
TvhTpxhhwAsBzcWIFjBeqLEAh6pTiUgYY5W6+xOk4BlkwbfleTaB3qfQR8If4gWvAPWvoLmtb3UE
WuIAkYDlaAfuEMfDWdePgDH9hXBdgaIQ9Rue893jE/rgamFgp8CIYlvFmsc/zta2WAxlVGJEIyig
G5KHTeKrh2OOM7SjnuDdrIr7U8KEPrnkveeOR+zmHPue/iDxA29bCtK/Ee0rd7L8wBSabC7EI8NQ
GIPtXnNtXFn0iiZ+QVJKMDpsmwkmxxIrq3NcKFa9fiw6P1dkb5PuwabmvPcIcBpMKlTUhStY4zvL
60iqhN0PqZZcN/iFR/OxAofrOiiRIyYd4+7B4ZxatUz8WaRiTt0SHDrfYWixe07cqTVrHu4scXn7
Y4uWvhhWQ104QPSMxriJo7Fw+5Ca4tJ4TXwow2QEtBhYg8HUPdE0YQM39TcZtt8dCzumUW/oPfKa
3DuV/ftmGvC5qMAG+Igpc61DETh+t0XE+BeAtNXUC28rl8YRzmTlfBnFoV5jd9Ozs66MieJsndft
E5Zb/iaOApnKJ9E6v6nXbfPlkT38nayCvJ9/kqww7A6OrOK/LXUd9RohTDyxFZk6PrrPQCaoYHoC
XxmQkZX2PuVC9F1fp25q2qfChc6ipEv15TRTT5iKzXi6+qJrN8MJkwCPYxtRsfygYkP7CGwj8lBx
hQOFnOPCqPAnzhYMRTp/VNm78IlIJ8LsurgxPt5KFsHR3h3X7Ll+yz+rXeblyzI9TDmk00HQjt2H
uvHkhXEJHFiXI3vzp1+yCGvlhvkKiwGY5J+MaxiejlTTzyrzAY8h1WB0hb5j4lQmucSZpYdB6hyV
6FxILqhbNr4V+97KzW+pmm2rFZETvYksiAZpi2KK5PlLaOOABJJ1PDn8rF52zPmIRgKICVDxjiTA
ZzdLg2pHFvLP6j+qbNQK5mIGeGpafeaIc+f3+uC7u5PuXcdW5Db0FSfr/Po4Mrjvx3N8Mg1OScIl
OHAX5Txs9u+6Pv622HZRznCZEqSAFbrCiKxIzHzpZSVNhrlJSlI+8SkWLpgOa1dZEYD2MEpTMJj/
HH7guBzcCfXg1SMhWCqusXIDeV8IlIqsGOB77ECpL+aBjtjDfQVU90WyOx249AtR3UxL8zx2eZkt
UWwmO2CtbR+2kKPtk7VW8eesHmGfl30lKiVPPxKsnax2l++RDxgay8mJbbdyOglXJkxI8srAO2Qu
i+4bp59w4cZUmv/dy14Z5c5ehVxOQbquZCxAvXNO5Eyw8nxLfdyL17HCDngOTkf2ZV0cRvb5RU4t
QonTX50BWRb9iv5De/F7kA0RGj7ADAXWmTMjBwOSCCaZMoZJQdJkXj9ua8f8t0XjEgVRZhi8MIfr
VTLNvvhYJpsilp/LgtNTU4pKNDrZvR2SututgLgjUNyvbP2XWCX7ckIXbv8IlC/GJfEQKmda3HBb
zYAufQlTl2OP4o30mmclOSojOTSEf9iwr1/y+g7bskFZXLwaWYwjUKBl+rU5cK2b3CYzZ71Pp9Yb
+xODlwpUUlO7avxeefRMiUoxFP8VOmusW3COtWIC4ihfWz/W/klL2zRoQkT/vDoPHWhp/fgKljlG
kT+8irW0PeX3VFR8KlvEsoc9oHaMSjN6Lv3U7EwKFTJOXojnzBXMDfYKIvh9UO+ABX/iOFq1Kd/P
wJr98F0VDbGjgDkkc1MDC0NCXhYeZA372vCvI6C/PsprnRwxVBZHJyaIdHb5ytAPxQUgum3iLPL7
+ebXJYRaxdatxanb3Bd7KiBb04qEzgD2eBP+PcJAlEyCIyJpmh1WVjHBAB8onL7HAqpL9B0qbXbG
+UVx6mXskG0YrepPKa1B5Bzn2jTVpfdELvhpuDHkqN2XtWTCsUEoQgcSQB+VEcuYSVaGznknaOiE
RN4gDrNmQ1xnfoSKXXSe1kgzOmyr2pOi9P3ED67STMjyIXpHGOrv/e6Zdf5Mx01t93NilnlV7koK
54DwACZeo6muE4cuW8V2nrwBMk+GV6K1M4BQ831S5exBVIIk5n2IkU0pRxgv9PyK3PW/BkLx8Dp6
pIo02+QQEFJZaUNSqnC5jrk72GY53kW1NaqtUx7N4P6mCy2ToeQ6QqQFIT+amRb9cGwR2NkBUZ6C
JOL67hofg3N1wXYuuAOQrrSvifpjXoJ/OdFTBFn9iFGiIMufrXvGNQmEzJXpxaFcAnaKlSXLMJX3
bQ8/s+iN9I1b8hjFzTTJ3L369j2AflcDUIM/GbaShj55OhdX5F6/WsJSrZhEe+hltojjRT1kX47T
y/FZ/YYNZ9acShrutHtco1ccBxzcDOgDFdemQ2r033oVeonolbT5TwXPuaJR00cF2cRPd8FDvVio
aJhwrunJqRuFjDDrrNPJfVxEVy5XFlYs1HgN50i7zmIhp7pbp1azKCCFJHtq8V2EzubwtIGjACZH
On4OxIiA77/noxMGQIMR7dCLDWW9uws/jNLjbEoblyh3qcD5e8PbisNvk1lLHqkBWNzUssQO+7o8
FfpennMXUn/TeV0o58+p3Y85DibT1rhZoGhHxJAtruqVLSrBjkBZG5CFYTdQkubAuMC2Uef797xT
n3HkbPQrzPC2vNAL3BHw2rL7uv+2v1xS0OrN7rkNQjHAhEwuk1dhRep3lz6m1m5U9vuzhZ7/PrxS
UZWjVKBV8ljGY/1wTa8go2g71IVJnSIBvN8MBofz/YMP/X9klmvnBGgvXYNcz7NqdduHH7DSAIsc
KJYCh9gb28PtPLFW3mqXkMg2EjtGVVsuqBhFWzQNdGp7lfiuS0XkMqmJX3nbT+h+oxmnEL3codAy
V4J24em2s9b6Uf1a6roFLVBxjlR3ndjz9XQMPjohXcIHJB+qVmRGwJ97NX/L487KqXtlx5yoy148
hE8PX267kGzmcfiOSwoqEnstuB5FaZrfyrk9NxtnzoYOCtpW7wUIHhtSMPVfMEdiaebm9RELVxeE
/l6mtTN9hGVXrpE8ohr02o4cpfqQMt3ec06gN54cwNixqWHMUNHpT8OshZVs9DF3N6II4Oe5uU/1
A96mqbVrnhdTTFqpt5GEHmX2ELjK6Ri8Zkx6AP55o8GUzZ5TSQOQzii1wxl05KlH0NScSVlR5Mu+
CGwURx7oa1j+RJsQOrmkEPHTO0gjNyElFjmVxcmfU1A/Ppq7z7Jjn0tik2hGVHD/8792tV/Ocafc
zcMClw2XMRkEDsLRoapZvu5bzfmnSjr57ZOd9JDcmC6Roi8BJ+yylFEiYdgrY1aLC9xYV1MdrMQx
BdIsPanpzWkJl/xenlJd9/l84hkLw8dmxGvxUF023Mj/zJwC1J3+fRAqc9wB1NOwOfmLpSWAIbEN
5/dOrRAcCs0M/2CvAt7U1+CGVzV6Zky4tPjvePiOZmbBAVVod0SBuozZGAMf+ej2r8lXdiAqad31
gdpCaKVFR2XES1jMqwlJfpGyyf9hntXJyfiHKL56LfqatBBrnA0/tmov8DwIQqrBA4HXKmk/6XKY
ijZb8SOM071QaMAR7GTVyPovz5NTdQNSGR9WgDVOdGrl5KJTwz9LDDdz8j9zjM7Y/tQnYsay358k
wgCY84/WdtdFDmp7B4Sjhdsy2MAZo3jmR1q0jL+fy2HsH9+p+U1iHhMilNQLA9+/GUvkzTECHab0
RvlC+CMA9aMhZBuEY2Wfp67QoKnnyB4E0/RSQuCMDYQdevgGzMgsIzdaLGuDRiQ9eJXVxLiz3KjX
krgxO1YNRGzCIXs+1CVEa+bLPoxuhHfj+ZG0C6FXIz3zlkRRlNIVJq6STO+K4fqFrnLf3fwV7xEx
GFkuOQnMbxqlC8zL8AHAqh91ScU4blojyTulV1AZVvvQPWY0odYEJPDaMlAAnkrtKo+12Vr19Wg6
3O7N9KZEF0rbF0Tle84m/GDWQWBZQ9QP5+FuTRAhWyrkS1pdTqAABw91+o0zaLnjQZsLTvjsUNEH
lQiZQz+KF4E/9sTtBOhgRVv2rOxf4+IZ/Xj6Ty1M8/kdnl4u98aIVYn1/xvKkFKbnUAd6XcAa4os
e2mtaA2tdFYq0DojOu0XxrfQnjZKOxbXgLhjimch/1ORMVm/tdLg8Xzf6GEJoaWA52UG13GA8Pcy
6XPmgtj3iRZEOGnwIZZp5lrN3h76Do4jJrDRAy2+Vy6wm9N1y0vnlzRArU6Fh1gigFHL3CEbqxAM
QD4JopB318h30DGDJMct1nqGxoP84egxMS1YtzdRu7axajyZ6yqhZ35EPAoDvNmC8kwKTEgdW9qq
gx32jOsX/p57cVtHCxvLobeuRXOElQnH3ZJNZtISyrnEUwlidwD1fZ7reK9ISMJK7Ld2O/1RhplE
rVLBhbyoyV2a6B8PYuucWAzb+p7gPkiJuxpQjklifjSHf3R23WKZ32zH1+uwR5SSJ7KaF6ehN6fL
dH657hw/YecxgyAAUYKgF4X48NcQgXdFpen+zTYj00csTfn22X+VPyXt+zUZz44zsv8qg3OV1kxO
aDtzesrwtecMmikTdR6xSJorzwA5bjM/LvCn/5Mk7FpbbhVt2W/1CLlio0RYLvOxbtT/mpW0S6kV
kOndpXVeDZJpCQsLSFMLoOhydJMQyCpGZmJUZV4IFXpDF2MWtq6XFBkebrO/cLYCNqi+oskRBMku
m/Dp+OAO1Fv6VTUkfNF30umowF5YshU08+hveJbvt9NSiavhJ1VTzRENu9DwQPxbSRzrYsmm5h+m
M1SZB/t3C0SncIr4J3tk6nai2dd0hSEPz891fJZNnTIYsDKgXWSyx9KHa4lTo/wfBWPMHWkT1VK/
NWTHgWrMVIwYaBoWh4N6crDdopCcVuYdStXpXDOD0bo7XdOL+Si+f0UKHV02ToscyHMyzuu2uKKw
JB/FWcJmw7EHIcnK+TzPkdTz6TvhuxbqU7irQC7YEAli65AvMkpAmaLDBII4Lucj5y30xHweLnW9
d5g0EvXJrA8TZoOML+Eh/oQjuZN5Sejp3ovAERihzunu+BxDeaHDYeWk/sbUxFLJXfgZzi/+iIWD
NQQ4Y+QHEGqWT6n2IJM5lag/dIadQyZwTtevkfFawxfQ7NOXOtP7CDX3ysBqLYDe3KGaITL0QZlo
5r+4ObRJtHDL7dDGdq9YZqHpZGIi7YRztwo+dO7p8/t0rzBuYZs1B41cBFtYDbyhyRvP9QBztNpy
TU8F0bGRhlccuVbY/Y2UsJ/vaQRSrG/xsM353OU7v0zuq4QF4CzaFVjB3gsWtVx+5fwUv5iOs3mx
RGXYnGXspSulirafOhiOlpqJ4VegjqR5yvBJYAk2EraHPla0qUDsbdH7X7hecWBzYeyBi7ikN6yq
TrU+52AC8mk8DqykCuURjkvICWFuiUlQSbkyu5t9wVz7B2thqyhQ2t2PMVykShfhh0XCn/TniNLR
ws8oBn7jr7HCiy2BcjfI+3h6sJOnVVbuxv5qMtNyBdWaI90/Xzyg58BbJtlbB635npL4Bt0Yz4Nb
mhxGtKpli7/r45BC8lmWoBFD/czLmi3wZY8f0rJ7a2Yls8s3L2EBT86+pUbnCWjkQopprnhPXhME
S7o7lP+d4QbXIWWIYkEZzUGrdt5H30DRHug0QdWKAB8YkLfpo0styuoYnzrl75SqD9D8Hk5w6tdW
Q1JBI23prgQqpsMK3zv56HFLpqaDWpQGqkeo2gXM/L3iYxsMFz6V4ZBWEWAEUhjZ9NyFJ/Pk5h/C
2s2gkzftAV/1k2nEBSnZWDn0pfGZ7FJ4Elt2ja+Zjl1oJuLuB0UL+MTJZbdjxuwhm7bRUW0k4JIm
FufICw/tN7vQD3KxcHqobOrFCZIbtL6Wco5YalMko96FX9tjT23tA0dGYHhbyEDVK8c2XE1SwVSG
W1GxgLP5UalQOb3T8bie9rqCyWSJ1fH7KaUQFMeK4JIPfeQ7tbDGhOL108ehjlEwys5/8YVv390q
fS/o6BI86q/r+V6peCyOIBqv5L4zGbQe7hTMgjkC3I1XZGqe0E2SpP6JdKzA8uebzJ9Genq0L/n2
qsiJErA8SJDxZhPOtagmW7cIw6qEQ0/o7KOcyrrMEwNDEyeDJOt/Iyu0xgPpBN0IVOrcpU3D3z7Q
ipZNkCjSfjqp3tzwZnivseIW3ZYOu571f5GSj+4P8q/uEjP/BSSgRVkSz0IEvqO6pWAyzIoPkI9+
SoohIlKDrK4DgP6YribyykM4kjAN99np4qidto8B0iE5H0qy0RMjgc/1wwmJ5MSdxuBuLGCHrvgV
QSrXb7PwHNSAU2MO26FKlgCa387BYob9HLIL61Lgy5eo0udJVC8BComBcc5MlxX05cljieWm1AFL
jfT4cSr/hM8rEWFKaf9lYFUKuhVBWtHF1K2q2OxIpmkEYCaV4KoRPOkSu29+AD0n5hJJw9qonvBM
bY2T1Y/nscu/CTGTffwReyH8GBAQDW/TNhqUXjze2f0RCF/fkCWOqFsIkNOoHLeb63yThwjfVhsX
QTl4jhhe0gfdhM/AHOXr64PCHDX3oLtI00G82WD+HVsCoJxff+7nCaslNStQ1xApiy8T90RhcvuJ
I69Mo59fNPDlkqQgRhQiYp5/pUqGjZacEg0BGqUCmAaBVvGUmLT92dX2WHYBJ8giAhElQdulHlK3
5dcrjsj/XxbeQREHevXL142MfFMeyFT9E9S2P5hrkvXladSpOt7U2jswvpoy0wGbbKj0MDMZhQ1p
ls0lj1RNS1nKqtU4ZzkCUNNVACdCTWBdddfjmZrH4TBq3JlJ3AqvaBe38tHYDUiG2xsEBdVu9gBD
hjZ2mlZ8xl26BsFkUeSugETEc3mVMN3fhAaDs1IGzj498mkg8O1Nzah24soPOAYYvHfPHLAAvcQL
BlNCDUsHURZeYm1L92A7i3o2cl6idE88uJwS5nUsHjfAMmYIavWkXxKRtGR6plqfMlyg9kblryqz
FLITI9ebYzLws2FkrV+dJG2ZvpEDbTLOo/9drwCJLMjZX4TkJ2oeCQh1EYL7nQT3k8GvECeOZScr
8gGCW92+RayP4Ick3visW2zs1rsLUHTu+INIaWw8spgBvK01T9o3annx1jVsoYGnhXKDdF7AiWZQ
7VTbHMP3fdgBYF2yh/InY0Y5cX++mN1/hNK5khfoSEfaV0/t7DBq/eB3M91yC+KXci2Q2PWQ3j7c
qDLBmro+ScVKiYsIaE57f5D+GjmMv0sclYKcHKml4lsngdhXeL/g/A0JU//WaBGSZdL6VBRaVHEI
NVW1AjHAC/5uRfhiwHRIQcThP+9vSegMkugUGRoZfzyxRCno3m+bM+H4sCfeLd3LLA2nIZPamVsu
H/zggYcDMeQjFwl9RPrEJLpchGokF+A1nIjAEK+BGC+Ib7fztIbyLxfGlUpUzf3V71ib7yu1HVgk
8kTpClrWCijGQCwpCGBstbRzH8JyFrM33XzxB5ibhJg1kccdnRwazDSIhuTj3MLAG7yqNER6Us/K
2WhFiHF3Alma3EzalTGjCYFaXQvV7t4PX0OHwZH4/agxQYm8SCwKD5ESoUBqAHOf+GgDpmAHXmHU
eSHvyMN1DQ4AZHAkx7ZE+71sI5179y7zLpHmcd/pWFAQ2mgWjwgJ/m0Dcb9bhA1XsTnXoYBhZpVt
9KXIf3ET4WsHzHrE2u2Dp20YdgT4wkbuC4zYYKBavgtRQqBgNtuC6u2T++9ECYGy0VJEjaYdOas0
H/wdnWOT1uRxs7+u3vlmM8ymo6uPnR83VmaEDhjV+MOBJ4fv7BKztQvBg+MGEvNDn5xN3vTotieC
IA1pEiX0j69np/k6kSlZuu3EQXIEOowqwFUA1npQljnInJ1nx8q9obv95SO3Gp0hg32VmFbftvVs
9j5Bua+LJl52J2ndXvOgQoQ7rnZ5QHlZDqTPOm8Lcs5jiG8nMArOXSX3M3r3b4EHvipt+W3N21sS
1Ggfow0ffRzg1ngeci/3BZScKvmZavTbT0l3PyHvDvyAIEnwNeSDubP4IlJXQUvvFRN9o5AbrTA0
a3vNCOBeJfIx8lDNZqSnvOFZFmhTY6zx75VdK+X/9KsMzsMJXlCZbyCL4x7hr/tKp2jQheZhL0iL
uB6Los1guEZQD1W8poRQizNSDePVbOxdZ8wn8xi6RoPYBNU4yuET/KYb+6rLp4ARAJI3L/+fkAC8
6C3FB2AQTHO/8Qo8OoqcGOrfLkcgRDxN811Z+HQWcG3KBfFM9EmZ7ICdXFdomZMg8IDQmIQ7wLDw
V5oFfD0VpAA2pRAqC+uqCWfHkbcP1XYfynoLvYD2isw0vwdHlG+2dZg29x7E15B+DNCCMUriwVWX
OLg04e1Z7EQ3TApNP0j4hxzrhBKF2NOAXOvLisgDSRTF0jKPFi5vv65LZIUF0jfBPYiobAjPpwni
4P3z7uBC+qhQTDwdYXxrRt1wKtO7n/3wWa1gMR/i6RuSX/5Zh+FpHTGNpGI6HqtAsfs5JvsTI+Dl
s53hU14REwv7UiGVKbYA9yreLXY29gqXR1UHNNkhk53bvCtQTchQV6MyyXaZ6ibPskkcp2zFYLov
wqEs5UqUvE69ckvi4HQZOdS9mrjWgKcuSIqVaF6+amdlSzOgNg/Pa/DzFix7HKoWNx2iwpkfLTkJ
b2dn20EDLgLtu+KHmwCeulLYxDghhFU4Oo6cdwaU19Od8KXwyGTD42ZW7EKouJFpiRuiTOTFoMp6
jk9Wy3hqMIF/07nZwHwfyhjeCYSqaTtMhM+/eRlcuCheprIiWEAqKLhKg7TZNsi6EOuqkkht5EN5
PQ+9FKrV0zIF1BBGjdjJBmwfg3TgxARhoURhMsH3jfi5bXoNeOGucRUE8+z3Jfxvd6MJ/tTMTj48
NFM5roz84v0Cuih68Brp1KW9/zUdiK5DLsvFkz8d5nc4WrB93b9JqyA8qRBb1w2eymlIfnaAXTxf
diXmOsZIdfTTjqcqzEgvFPlFc1nmStXr/xSF1lpnOgZWmcXGUR5sJ9J26yFYk60ojZJ8PcEwjNjU
vA9v9RuSD0y3l5ZnD/FRgYG1ZAybFmKtRDTSFmogohb9INGMekbfW4Gww2zoVUQyJPedszp7kSrW
8v++tex6EIDtCB2b/j2atJxvmdSUfccDPkDluStHrXjPuINm7V7TkTRNHeHyBh0nTCa7fEHMWAGC
V8J2OQjsvUZwbY1ygNMYL4/l2eQVrwPywcGA8TXlGKkn2C9GZTbLe96pg8sMWt6jhpcbHvSge89Z
aiHuCd3wNCV9jVhCW4oSjexzj/nO4yTpVTkA3Xq+WsYS66e/FkuSjSx+qdPG1jzWsXXmfLqTx3hQ
3MSdRSR5QF0+ZjsH8uklTFYmhLFYqb3bCAqb2WKIBXVD26HKSnbppkTW4GusbyXt19zWzrgZTdr2
c2Dcgezk08dDTROTT6hF5NpMuogkw88+sgQDONzaJcup9rF28WME+Yf9x4X8QiSo9M3+dlcJA6k2
s/yW8C3QNelbiOamRBMhjzw2jW82I3dc+cik98iQ2WQ5jXxeVTFdZqPDHg/cDokuLwBhYzn1zjNQ
MdXP/r3Yr8LMQ3ZULrlVa7yNLdkObemvcDY3/0nfHyDpQySEGB9JYQwMfmGBp9d/oEOisOVy3rEI
248ztB/lUjtMybdyxV/qJfAL2ucCpx0qL4ZtyvErPXL4RaZdD+KXuSGenXO0XgmBDIh8A3mQOZsO
lCLiGFAvit6qDl76bY3tF3hWx1rLZRNgx+qvS6TPpzPKovJ5P33NAMqS3SyREaydZiaerLYx+D34
WVNFbSMOVN0gMzQLVL/ptN6NwHYlIpsvv3QAe1j57aEErZPWhyNmEhtOL3ArhM4406vlNbzIUO2t
T5orSq4ChgNtJXJ2Xssklu1Eag8v0+TPS23T9ob+B84voHna3O99n58wVqrw89ZqW6orfXlNNjPA
h+o6C0lvep2LhIkzjmIsnEzFn/8VajbyA/Cr1+DHRdN8pwM1BAZX4kVMNVkr5BkZH7kdyzAHysOS
ZMSZk8dUwXJuqdEU6yS0oVaIs8ce6fiXQkurNci492DhGisB1o2xw1mYjLPLwjcWcjcHrZK8QPWe
dlU1A0LwX5mC/Bh6sz1aNTMjGHe5QqMoxxbx8QRnxRJJWbKGa/GViQhSpwq6EIPIjlz61Xezj5vD
tQjwB43PxonalIqFeCtkg3/RIef3JkTJgltkrTxVdjO08/bzNajzz7F3izvoPEk8AOsWqCZgCYpR
KYrFGxSSmb4K1Lx1GtP5MsRtUGLeVAWFxwI6Q06KCAoNPP4b+TUOLtXEn64igpCs50f0whtRIkyK
GrPVSG0w4chfHFS53arRUWY2C4x89T6zqfLExVun0AtQ5ibKQy8Ih6XHcBbOev0MHeEMNK8d7xJ2
Uo5hOjmUcU5fbHu2PKzM/VMH/oLRHhSXkWPXNEAukhIk9MFYOCHjYQLu9nnqWZ07m2ePjs3HskRx
1HTwfzOuiPIXIXY1Wqp1Gh/lI0le9Jq8asHiEWtHEBAF/+F4ACgkPyfDjKU4voXq1grUQNqxNh4Y
/FaI1z/0EfdI33epYHoMALEZXvdRd3WqEAWXuyX3GUEHfgdwVxjszbaF2bzM03qDxovjwCQR/CjZ
huUFN/AFXrNlhZzzyWypblpFKXceNqGyKLcTc8HafZub58pwcztJbc/4m8I/7Et6GKxtm5FjF1no
IppapbNh6IRWUCle01ZV3skFA3pmG4JRliCyh37f0mMiwqR7qNq1p1Q9neQFbGVJlAGxGiYIu4JE
gZxsWjwFwwWTExHtiukugNpUOh/nZFR/GiYwK3Y3BDhi6hhmI6BjNXxIj+KNavg1+EPUcwCHQrQT
XelL2AJxYYTU+ryqPTjT5eu6hJ2uwspm4zKpvs/I+dInblW5ETgGIdSLwcDo8RI+ulMHtWgcewXk
NvySVlo0bmFQHQBB18noRrTNmCIYpbakRM7hd2nHdGBN9oKeIY6fi1g3b33kJ1Gxu/MWQEKFMGUf
4OXBmjn3Lrhj/JdJyzNlfwMSv9XlD34QLJNBdkfmKaBzNEIyVlUubPjEz86KdFtYd9lMEkvLOOii
QUcDpJJTDX6edxi18oiQlAzD0jeKXJsbwcL8LqseZ6BRO9v2QWUBdycY16oLdsBRJGJgJysofByy
x3u2GnWhJKstX6jBLE7jIbpbK6+BlJb2jmMOUpBvpVsQ3E8yFK+lEdTvIErfUJtKlRb1KljPnulU
Frkju8vryBujKsCOLAOSAgy0OOjjfyNthcuDJUaChREw2yFzte+aW60zM+AmywafDQDkvx3qHRaT
OIgvsbrYIqvD6RrCKudlaxe69mcLfyxTEEjmnqYZTlvY1tPkLyFmldF5MOWKg/0urPQ5iYmZ/QdK
p5iy5wTFkbGw/vdumX7aYzVxoKo2VcBiorhGxAAO4G3HUa2CEfvM7+mDWgfCGKd/3n0wvC5opo71
H6He3pxiJ819nLpfjVKtKiujsNL0Y60Nb+xVHeXg/jS4QEGNhksIIENOzMMgXdtVpyTK2iuvqKvu
bNZ8x01UbhYMSihrur6/DgwV71/ocSLljcJs3PgmlrIl8ohz62OOBnWsOwP7Fv95/Nf21L6l48eW
ixDk2oewt+SbStKtAHsJQTzUbIe/+tE7IAioPR5Re9eX7mDQsMZskct++pwkm7YIkfaxTMGMUESr
qBQNGxJIn+rIc9p0mjnumbk1WCKpH7EJzsBH0fk+zYeh+Jlm9+Lw0CC5SQEfCAkMgYko7yMDURTX
cI+6XT4BAKAmgXvidyuOjOuLTDm745WcSXXCJwSpIV4ceV4mj6sjmWzbCD6oNhUOjS4boQQFyLsz
XcOhzDQLAqjnBXTh6fbnIsF/KTMTntsXIWsDW4S3+996Wo/xLmki+xHaIBW7kGORh0QF6WZfbOaD
gPwzcKSL/3B4o6aHosdid4PfjxF0tDpZFNL9NCW696gqlmJpxJ729yZboW+zZyyYDVZbZzd7+dy2
D61syfrPkn/SPNvP627ZWcgQzDvIviyWqH1pZSnmmtY5YNx6vPIWCC3ZpP0OubyOW0WsCDuSKKZE
006MbcFrc6ciEIuWqdlyCsHSvs7osGEyXlPeEsQcO8ExsChrvNpnLo/JxO8Hyx2KbYi9BxZMuwYX
CA2iqtWUSSmEKGelPjFdB5iGtjbM3SPZWNN+jsLT4UQjLZVeKLFe7ZFq2mNSJZb1Lphwwbzjtudl
jZ9nY5zWf8M6Us0wpMSB8yvHGmCBYajIzPUgPtxmc4xSBy8YfpdwXeStFSD1WCejo67A5FXdEDgo
1n57xh6cbFTMVCMZCyvYEjIbCgTDYq07+06FA1rgS+SJqBvq6Le9YMtzqVOmPmVgJ/9QfvkKmy46
+lFCMWE0uUoWKWCV+CIRVGLqCAs4pUCELd7zK7xlaBCLO66MFBd/syxSKReVT0E69m5HzlxeF/az
OTLc/MGHZTsXICCQ12lEF1E+RGWt9kOZuBMOP/iG2Ga9qdW3JmKSSfctP+o0wT9ZWTHz9rhbWkaI
rYoT9BnHHx0xMRnNjIQcFjoznERmwMaIyNu4QrYDoKkMn48XTTZuS7oYePWXMw4x26CLC9qczHoi
/cvYKsObh1e81Qpc6dKe6CRdSuFdbG4DvQcABcWjwniJbC++KZyi3QZwj9wx6LoG/H5LO93CRvu3
3AizFa9r6RR6ccCJ7UT258j7mEctozc39/ddk1ZDwXOvD9NJMQWzkIbuPwDtO8kZ7SnF4rbLYdpd
yeUhqmq78AnsujhMopj84R8/+d2ga2ZRh6eDJW1fQcEfHsThsH3STKJxHNEb61z470vaNjsO4RLx
kCBYLKwJYL8muEMBFpFk+SFiOoept6EK6u3I2Ifx3tpyEhGcQ7onHJVSH4ki+sLXoXOvJCN/+9i8
dV9X3tXlNkuLSPuMM7BTFF1JxfiLAtysDcTajx/d0lkX25e0NfTNfThaPfCundKxyEzNR4PI6+hF
gR9FPA9+iMFb4Cvp4HNRdyITYMopUeDZqfJh3O6b/Zmam6de2C+eJtKm3cHbvGgUrbilsAxv18yi
+H+sTUR1KzZW3TnS70vl/nhJ2XGnH3MJFdhSxfNsM+llYltX2q0ltHYqxqsbIwu9nNG6L8Dg+L5F
5TkFWLHvrSB4f+DUO2bGf0fKOKOWOW+6YGV//Ey5wIWWI0Dga9jnfla3LUTw6bRnoNJwg++YqRFx
MJa4xrzPeKTPDDWaZITHyZ1igF3umNpEbvRNNi+1TUxt3Pu+3OhkRGfTJht3COD9R6X5ipPN9ZYn
L0EyJtpTMZt6236aPUTiwn03FgXNlYN05AKRLdiVnZpkIUz9P4q7lWuoy9dFoVJrMWc9AHsdo3xI
RUULWmXfpAeypGTb9hapy59WD5BC1aJ/EfpmSIIBJJcAgHbKTQDZre/+Iwb5dCeaNLu5xhnXsUTr
yLJvRxvlYjWroRnMXQ98jnsX3HoAyXUszsrH374he6n5cZ6BGZGjZ1gYCdXm8G+ysOd1kAutQ9Z3
mIJy1Rn7RcKn1Gy0VFaWb7oiOuT7WO2NwdpH0AZhsp1gSKpXy/3S0GNt+FKCsN/zm0A9MKAPd29M
gxsH6bBbHJkGpQBXXS84xMzkGtpB2z60Bhq+a9G7b9zuFX15GGanGkIhND2+OcM53sCyBbEftyUk
AnXa6yA4C6LFBmWMT6E+J4WRc8PVdZuKm+zoNIUojOTxCsHwmKlK7lV5UGY8zhsKKz0WsDqjHS+y
FhOxuVnpyuaFhcJvYZhfHTdhgkqfJKVZlMpO7qzKIJIL1kFxeRJfeyKYCCyy2B627HTbJNfydoy6
B1yoPSijpLVa3l8gn8lz96tttJgbyd/QZjkKyYWd/NDRgrn6V9eFi27sBmfWVMfEyE+YICTzgYaJ
kofRmilomrhL9gyMm2CZMilin//pI3zNwcj2gVIcv6fy0rEGm4VkcXjWhN/Q/Kqd0cq3f5chLCLb
BBdr8ZzPoic19GSNbDg/CUYIWwCNgFBPSTtO8utwqh3ZTD5kdPc3K5ak/SxN8/PSiyAyUuDcosJD
onXGvZIgXqFmJI+X4fS8vkvdLaqcruIndn3CC+eDcq5zdlednEIhyqjBijn7nA2TBHpXHjxRZHJT
slQhumj/nd8JnmW/x9FqC38i55kzI0EVKO1j6hkOqg94xSCTDLfI6ehhBj/0NF+lVgAl8r7oLH5S
tjmjZai388o45hwG0EMoFXx4qM+7SpPHyYw3ev6K8pRQYDb5U/E40jByVB82RZp313VDBg6XnE5A
Kr2kK3y1laDH8WpoPOHAmLJJDIBUeBdWB45qrcTfKHdmXLHHWAqRyr5Dg80ViW+rApD/JlPzwKzJ
exuXd/nbOSdKEAxDTb2vt2BfhnOumTp3VgWUVwIRO1o92TF43vC7NcEOyDDdHYZ2fyl+KNP7uuAj
lM53xSSwEyf5439Sk49ALNinWOTMsPnqO9zQI3MZYwKkoB0GoULyISqpPOf2pfUakQxkio19kJCZ
7qcQ1gKYqExxdSjSY7awsmXt0joSl5zpIM9B8Rhz+FZwgSzVloahIKsSY1IzQpJeQ9HwHXIww51M
zQQX5ZvUHVzuR421vlEuxnZEIeWILuJpi5FRLaxFkGddSTh/jD3ppqQFURvHbTL3VMFkYTsKgEC3
sd8asS+KGot+TkRr2/l0oh6GZ70pAUoy+LCOYWxcrT+gA69LHl2oB5bxpbdspYWVPLIjRRvMKlFX
VoaNvMtRPBq7Ewk7SPxxDQjtNSS9olHu2uB7MEn3Gj/I7KwYa5JKS4zMf1Zt16RAlUh1LWFT5DlB
T+Y224zySUpytxaSRENNzHEEVKkPSEDmahgJAdZppfLyaAQ61Jz6Wblf9Ca2C76XmTqPLysnejX8
F4H8HHjh0gtdByT6l68wkx3sZKMDWLtm2Dyg9zJO5u7Zuv8KzmjtbPUAEYY7BjwafLcMq7kwmUH5
V7AXwqWePwtFz9Wa8tyD8qTmyGe1PR6grfBeaIisgykZmvhz6KO4P1H4r11GzSypRROHorvhmD9C
+CUfXMHvugyaRFoUToWa5JIpHYk/A/MWICk5N3d3bOjrXM4P5gAJqoG7wd7giv8liN8P7QiXnx9s
xWDJoXJj48PM90SU+QtLr+ZtYH6Ka92UnQUbqAh2OCS+g3j0EJJ26VrBPZbBwkfkDX9gxvYv1vbU
h85TGcijDclf5sCk9707UBSldOn8H4HEZj/WUmtjrPEqItw7ocUbagDz2C6lwrxeM/PjzP7tz+Hj
WSFEo6H3RfsyEI3wpZICrLdhWVhuQIJOsRzOPd/w3OvFAuEDuF0jSxgUc5taMhjV3ifnu8bAPKOM
eJbQ/L1Tz+vX1RL+gBnKVH+ox8GJ/dUW0hCtCNloSTIMxdvd04og198akK+qk2DSWS9HJ7j4qFEa
X2IzkepfKEUVt1ZoV9i4jLf7UgL/4BTZva4M/OCI3o24oZTedPcJsXAyh+3tkKd5X05lWS7rtKVu
y8XiQr9Ra8uGsidnWCX+i7+ksDH1qFrb9Ocwby3OoBP9aYF0srnz9fmeQcgXHPBch9Jk0JFK9A+e
x3SkKyjB4A6kYeTZpIHmqvtMvjTAMU7MGKk31rQJPeX3R3JHZXe/fOUT9Glag+C13OxLAntnIkg4
MdooVGcV0RssW9dbBnnogHEw7bmS245/1zdDG6+4h7xCNOYhD6Fl5pJwHigmVhmenmL+5XeTZ2MJ
c0F0ONjxose/AHJEfOTfnLEzJtyeHOH8mb2u80O6CS2ajzCLnBuwXdejLPoHEju2vKBoswCJ4HtX
JFwhKlzZx8f/3ZXXUi0UjEKr7MxqBDhOhOhUYtWNqSVrU4FfKk7+DyDmdyDCF1ngk36lh+96pmPH
cWGoJCX7c9mgqZAeo0L11DqKHmG2Xj5iuQnwtULDoKx7m6HKi72xh894TmTvcK4XULbiVH61rp78
n/X8WbACNXYGNUXfqTujlg5okb+3K0nT/mZzX38Ka8uKY27hZ7Z7UaL2TBF4ewAHdUJJW8rwGNGq
xbs15/8VzI+uY+4lH73ULtKndbMgagMIDSQEkbrdc1uuKd+645MAbVIyrvTTDEnPY+vbFpDE0/zu
p2Q4paCPEA3M6IVwrfe0bOTQhmaaNOWXORL8Y1s0n6LMQhJeiajOIMLi07i1/Jtm0p5o3u1L7G8M
JXH9ZPuaixZ7d5bgcZyd8O7NqLVKe1VAjgSMtWHyXKiJqVhmYRTiDolMN7Txkral6PRarkw5aSWt
rrKhenEprUTrAsa2cg0B9hLLQUcQBQFv4+LVE/rgKWXUigMb1gjVFvZ1i24t0xj8MT8KKJ3D3tmI
I38TIplMj+U+u9ei5rsDSNWOaFnMcAz8QiRoKKBJ3avP1A1dKv/kdqz32Yy3+JgCSMFlPY7pT66x
p5y/CKRHeq/xkRVn0gfZbiwBZVLav2Rcc0fPRwgYWGaT46tcyuG2cwQnUsV+Noq9BzQ+E/dB7OKt
vsWp7lX836z+tAMUceyrfEcRXUKBsLLZIzEFscM45HDNcP7r+L5QfNcaS+lw7bjVdO3vUmSMG7na
LIi5xjx2GeJ12vWOabjrWJPY1OqxiZQgDm24tK23NTq0/Hj2Tw2P7wQQXe4scYJ2yRDKJoXPetue
uKteVSRgtprCksFPct3FrhmTRXiU5j19nW+p6Z8LYM7fC3l+R1nuoYuf5rfemDEG5/UpPnLmV24c
IYjMxDtzyXgx6Ci+E4dSQNfQyOMwkT+QLtNXK+bxWOE4cXbJWlJew+ojnGbJXa6+QL6p3HG4ZlWc
nYzdgAzzn8be4Pzv+FnnSranFORHibzUT3TZwWGzZQpn9g91G6izeo7UGwl9S18LHHHqgRnGKPln
ED6LoG5gCTtkz8A8jW4W1Ka9t7HLV3yEGk1bPy683NZmiN8mUaMzblieH7jEJsROK6DKYGsAiqsR
G1Hu7uPN93kvpG3EY70hijeYXDtjw4FYkrqnS70r5u0JVuCiR3qUpFaV6cXGW6B9bQ+vbbtp74SR
RmfLKegjFlv4qsra/KAHYa5AE6wcxA2AkGMvbzXBe8XK5hcUTebZXxz5f3Gv/29/ZuPfy+yf70+L
1lekFuML5GNkg9nQka2WIfqTTcbOe2DsQqHI/MpgUWXuHy+Vs+F0yticMsI3pIz3lP5/uGLg63dt
cOvO0pTyF8MVMXglB9WmEEpXPvJiVIh+2wUVltBhfqQR8HjR08A8qmnqTAYapW+tohtLIVWIBDt2
iaIB3bxtnzeiF6Zycx/5OP/qhDXVUHipHFVZvl4G3oBHIC16X1Vx4JrhmBCr+W6cx4exSV/AMfMz
wJyvrbC2E/QhS7hsHJKUB5hJbmscKC8YKi9aRoszI94BVWfIsw4ZTXfqHGLRtD6NI+jjTRxn2HB1
lbIb/g1YiAH+dxtw8GmlVo0Mj5KOwVsKeaZGmP8xzeFJ/FhycfnswKH5um9xVVm3YeTpnhjw4PLo
cZHkqNv9kmH8rdOrAckUHPmEPwHrl+2iM+tzyYVP7nuFabFkb05vlxZOVu5v5NOyPFObwv3wnFYf
k4PatIU/U9+bs87jURo+fKEJgrqVHPdBxnsmqaQJSHZy4oMCIMq9pNL+uOayKdF6fJnEa78WIXvn
vS4bnDM3vVzR6SFMnmdk8SQy3XgFByME0EJF12xVU6sIoGRA2y5rMRJFucJCMcZP3IyeZW5i89mJ
uYQnKcJSzod/IIt/rq3pi2pwxMh0V90hER5/iA+u92SzRAsJFJjA1mMyW2exBP7zpWSmFQg+XY2X
iOXlBGyxFETC+tCTj5ZXAlPd+4VxobgMDgMs1eUOuhI4VBi5XzUfYyh8MB3kFwhtGWBUrQqnsSsg
4h4uDWdiPOIjo9w7Pwp43x0UZpPWkGmlPPJAEMkuYDHKTCQj0bhMtSOLeHsO15Eu0CrhRLJYJTPr
p0+GjM2u3WHHvmaXprISNj2C/potAMKCcbnYmAhxzX4KSdalvchTF7bmzOXybT/VAKLzM7GYYjiz
Tfolcn3GD0Zou2ZE0n7g+qS/ojn+L/laeDrJUnSzU8UYB02pFxbJ+xnb6EytnG2Y1gjXO2Cf5I6s
h/5iMk97raMa1tFXwf+3l4RStd+O8KWzHeFMNwiFH6uSBlCNlymk6ph5PQ+hdl/Aw08jkMUshkvH
CYxJz662MbHe7iEihwFgcxO3KIl0TX71leDRMrzyf5FMfC41Vx5k0t41Hj2p1uinEjQ+ggAyS5ax
WViHjBZk80/u6xJh/LaY7vUHqgVDJRrUwvh6Wwvk29DZ0FBV6CNw8nAmBEJ1oc2JhJzO1oIvAKZb
q5OMEa2MKWp3DOsIJ7V34Vf92UhehjHbyFSTtA4Vq/Hg4KGzVwJsCRgp4uhHwLzf7CqYMAQb0E6n
iVsh0YAk5TNFPjJEYix16x+PMWqwIy7dOpHI2344w6CIsYLQjORwG2U1OzTlltrfTsM9vbUBa+Kb
PSXdJxkB+85NahAEuBxskmGsQKD3ILQUXc7qXR8+qUz7+jR8uwCLKkrwAh6SqSkLH1W6JNSAqqc3
YSC7MOUZtV9lJw9AnCtO81LV6CtGdoUpTWWs9TZBfayRrxU2wY4mHrDGraKbokQNvx9GhRI6HB98
EEjKz18PpaYJGLQEryU73jJWwR4IGRBPr944Ou2YCErnGYrmK+cdPXK6Vy0AvfXM9FWEVpF2Jy4x
i76asz7REcHqgohlFEQY1RwCYt+YcFaXl6vuEoBG137JMfQ9su+ALsZThqaLyI1Hs295G72ELDuQ
WN2GDNv2mjkUe1f1OVjJJijyvGvOMs/kNnmhXVBzZLbmm0shGwL41RmzQLZVaUoeGAFTQK8sr6or
1jAt+cw6BDxG3zLHh9hgyOt0cRmYG8FRLGFPYVdTXmWWnMd0xDIGLXWteboFSB7gLy684PVjQvbU
Sc+k7Sz0Y4E+NUOXjgNK0SLCIvqE2x1VkNNG3UR53/lrfmY+IUTtbKN6kanKYdHnoLAUKCF0WSVv
vAeJ4mIqI3PLmXaGY5QlPgWSNPsUfaR7YgGVSTfb9XyP4pcJPPYrXOqpW1PgRn4SAOBmyTJC6tuy
dnx+zHq9j/DWqP2NJfMWcFzHuPsHTXi8y3cHRxL/Laede+wv/aktYdMBBetKiORkI5ylEkRyTCla
6679OLMk4FsfKeTWJGySFv7MSo3kTYWBc8/JfUqLqJsIJBDf8n7XfmXb7ndLicQeV/Nl7ZARCcW9
bi9P7UvFHU23C0xI46GowoZf/3lzfTGp283Ug5orof/TIyvVnDX82scRFTrwJIVAhY0Ijnvi4bNl
HdL7WX6M8XR3O/8oplWNcKblVy42CZSNlgOLtaTE8BlpumKd9+lUl+5GspzX4XXS+x659yLOU4we
JaRjKhLkOU/1/i1GmAIkIdJGpcC1vhFgysdD2BpAUbVAZK0N6xsx3EqZdsBFKfUx/CmPeNRdIv24
dHRWF8oZjE/dN+mA7k6vKkHh5R6oez73Bc3rh8kNSKfbV5LShQIFo5NO4W763S6ggaGYhd41io64
8RwV+K5+MMsYdOoQVQLKioZd3hZIT6qBW0kf2slgzPOLA8q7fACVS5ARhQO/S5Ka92TdJTsxGH61
i7rfo9A0+WP02YRcS+iW+IMx8uF9ZHImGU7XJJr+9JwPQoPYHs2CA1bUI1YWkEoaFOnGOwRX4890
pYOxtp6R9OYU2OL1Z8II5kexRfeYrHHmthxISQbz9ipSCLeVE278AsWz+znnEs9MFfhX3DFg1fr5
YScC6YlMPA9I3kyQzw9udBpHPMYeVz9zZ7DR5HvEAm8V9K4rQCz/LogDYI3AFIMWiCc9DzmRFxp/
lM36oZsZyxwHzemoetHgJ/26k3z9Ja0S0xTn+KGQddFthiQVkh8MhUiyiTIHbEofL/G34O3tgUp2
Cal/e8P/JAUKuFFU9cqEZj9JEMgyYE5sCHm7ptCJAhP979ks9KhwxnBoXHVbuRpXZ1JQBDMlrjP+
cyQUCciarKA8+LVbFHJsvyqgT1dWC2kj9Jpu9Y1cTU32Jp7vsg4BF5/8dFi2qcj/NVb8GTsx9Twb
tDe0EEUXL1UlcbCL9yfRCn5QoQD/gka+A5y/u6+4yOdR5I0P6fZjMKN4Y351fazxehD3rLFXZdWl
s5cOipGXBqU2ma3v82KtWmLRv21h/EidlA4JMPZ5YH47Lxx7E7iiZwD958Uufq5m55GQt3MTDSMv
Ed6B1emcHsosVgjlKJBibV0tLpvtagnfAYIflr7eEKzn6KXsXlnrm5GGER0VX8L1wcS8p1ySWiBa
BSzQBVtiEnZtek8g3pq13XE+KJpftS/jkTzBuTHFuauZhNKURaGTa55JzYPzPm15G7M+G8SBLq1t
oUsG53V+5olODVCfDABiOZstUHe6gEcqHvdmyMnWNxo4/V4vtVO3Zj7rhll+DOS1zRI1eqO3Q7Zl
oufa2CgkxQfiGM7I7TjhphtAxH/ordJjLp36xxEQhPTD6C2mVM6LJp3LmzknOaKWzf1A0AuJyylP
9blEJVzfvPHW43gW2m183W2JxAuBe5V67waRoZHDcWD3XBYmENO5M2yymIigYSCR9Ig82ybpUf2w
YBLszKny6cpttDCCvRK4tNDFCz4s3PKApN6zuin4cvVAtHdnbTZqU2FBy3jiS7z/EgSuCiv/OOXM
4J2uNoZBg5fy0JxVWP+B5Nf2C6HnuHKoQwZd1AmlZJ8gtccus7wlQfRZ3Cj3ZITu91ou4Z8cqpdo
ExtjUQij62lMD+slY10oLRgbZa9v6YlDFE+DB/aUI+LPuEiTtDpc92KQSsew6tEyMfFtZ/s8p7eo
ujuy0lXAHkbSyhLrlb/+B/Xyh/qtLqgJUqeBqz7ar2vKzkS9kALsFOa4vVC3vJGOGf300VFNuDmX
Px9MoTY6gFVGqw6+WVbaxMwGFaS+nRXKMwZG9Cm/6YJ4j3cqrXOHxHrwTCObJHc8l0RcKab/DtRD
pn6OPNwbvnfjgS7dHNH6cTcwK7V7gEuKCWfyct3PPRs8NFW3BivM4+ar32LXXgMYfv76C3KY6GIL
bbnvNMAeweriGg3qPx+ybuW3pt+Nh0GveKUmT2W4LBYeNaGbE+uNpEZUCrvodVRWWJuVMYSBtPNx
TH/MIt17KIUUPRf4tTFPbnCk5Rjvab5We80lxk5WtVjPkFm24ek3zu7pYrASSw0T2y1kCGKHzXxL
YZq0VHz11y75IRyWOIYK+SLOJS7L+H1ann9oL85ryoADVb7cmjfhkWj7R6hVuqkUkz0bMS3f75Tu
AfV4/jRmeBq1JsRXBEHiIemb0EMBPRL2EpIoJb4YDYYt1bx+I/+cz9Cq/jmW3AMp+BJZ/NLgM+hX
EqycEova7F5ShTHSwXhkjQtgxUaEX/AwwD6tbxOMz724l8JV/XnwFOvVThY7BLoBnj7VcYOY+50B
tGR/D01eQU2qyxIRoYr3BVCFL8rOryhx6fSW/5hb5GR4/smsqPX4I28r5S2P8hgLBXgrSd4xoUkr
aAmW2/ZJINFcloKXL9ehkU8hduN5LXZ17mweL4HSaIvZgzPBwsp9cU6mHAfMHH63xwU7Myn0R+4G
pJyDi9OqioCEm3rzHqAnGie4k6Y8uj9Bt1Tgt0PMlHJNuMVe4J8tMRBZ0CMa9kxuCDVMbuKWg9vX
PzJ5qdpus7rY3cN9rwA4GAro9YnC4/j8gxcfR/govVaH59wCayebNvtlSxkZ86QD7X/vCmjOx8EC
cAOvGipI0ySEWIE/wtyp5wwtp18xb3ZGHG4cnXiFosY4GIfgvtpij7IqI/vDppZSXfizuidYK1LB
afzbM3qT8TQmDR0NmruF/R23T4i+bwOM8xfZ/huQWlYrcj7BQVHiNapxcx+qzeyiZDpsBSeagWl5
14WcGMwoj5HZCB9881HD0K8ejo0zemXrQ/uReyl+2GX5IgIaX8GCIXIXpyeuFkrvjrHtkJmI6FLd
V6mhBfFgdMpKIHzywdok30bLDAibdkrT39AoFD8Q+N6TB0ubn/9waG31RoCTClSa+FcoN700Czal
9lqi4H4/odNtMEQQOAW9g+xtwsP4GYtcN9py0oq7B0SuUfrzvRD7dumcw74nS8158+9JlHXdZ7Gi
GQ3fre683lUZH7THlTL5Uhdktug3k6s1Vmrg1Tlt7kQPmgzn9xUWeBZ/rZEGD1mQj1PiMNZG3IEK
6hXEIAg9g6pyjii5If4T8GDV7q7JTe5LjHFuMbT7jCCZcVJApnv93wq5CgtL4FAUfu52DJ3qpml/
vHXmUIQZbzmETeA7BLFKYE7NmLjPxvKK2mn9NB6pt03DZV6fr7HN2FJ7s14c0aKNJKcJKjvWaStC
WdhcNkZKNFrCVnCUObCdPQxH7LcaR+AxpixfzBR9JccWsyyIG8wKNZdFpPHJHKK58eCXYlTtrecm
dL1NzLsFNB45n4kRbpmza6JWGQqkcPPWr4nONn8iS8JXF/zrAoOtD/hlAORHp536Dpapj8LJEqYi
b9JhASzeiGwoOlyGi09hCNc+RvIOfhlu/nez9PnhltSrrsFMwKpgU8MbJdKGo+tygUerJJ0ew6mr
vMVE5a8QncfXjZcoRorX5QxuZcd2kDCXNfhUscEi88ZMv1/6xlMtdIxpSDyO/ULehrccx6TvgKBn
bcaXK3My5pqwA7jqCPxqHdgr9bL8YW91K6ncxA3MvZTdJ5ZLmq3QJZX9eemRbwBhGWLLhRDkfr/b
RblQjTXa7KTK2xFijVjQd/poKnIaq+nEXSWm6YXCfuUXqPvLxZw7qKR6rM8KaM+BnFElz+/lZGL1
DPhjQ3ofHQm64Z4S8o8srqZpzyv3zgI6dtaVBoXahZEdygD7+c/Kc8RvjQEMTda+0zEQS059IRgQ
qKfc1GgRxltsYQsdWoppmQ9T4+xcIZIGGAxL8Po9lA48wRqjayv+bSUXwHhG0oEnb40lASojd5iF
wdkuQ52bFKJJLqeArM+M1NTuibs3PGwyzAhq9HUNY0VEMSifVhC5vl4FoeFFOhufNAduenKG9p1m
OjcwSy/i7XSoCxHPANUKJ5ZLKs7gAjrlzNnBEplfDxxLgSMDRCFp85Bi6zzi/B0n5O2mXj1XA+Og
zK1h5AOIJZW59KdXiyWC3qRHZnVVLtfKc907RyKIj9UOgzp4fFz5nAqyP8VWCaopSOd4Y0iHZUCR
kq2OksYPhFQS3Brf3mS7e0DkccS5WE6uOMYRmr7LdPiD5GPPIgxA5Nclm2kuL0pEGxYehFxZxOVk
PxSynJ2nF2mvH7yNWxfyRQo8zjrC96doRQlI6H3AqboqtBvSAOUAJYxXPjeWm236bIvsmLE5iS37
IRFpd6SC0TiwORSVqgE8ysL1poVxYcT6HV/m+QjpQUOuB9ugZDEhFXsNgqNEvvU2tljxuNz1WpkJ
t1vbnW9Oy3Ws9QYKchd78KzjC5icYsJGCpxjTumYsZZlyfnZ9s3I7XCvHGHocOOEEIto1NWXp/jF
sy2IpYVyvwjwlzBJ+t/KZFwBAvhRS3D6tgUOubbteUqS9vh7ad9V7oQi4Klx7IntaGscNoYLBJtF
EA8OAcWf45DSZsO+Ng/FpfeHsVTtTEgjXhape692D0qo1Nu7bb0SfkGU8PbU8dRnKRWs8mtNpmsZ
o9TPv04MrHCVPNYcEne6mXXRiWoq5qdLNSMjeu4B4BzlNhJWUCZrz5zTbwjd4wFSf81rcUSeSeVj
3lZ+xDrfl4fs/gQqQIVtfPaATUB9RipHIowJ+MKv+vhl4gjUxpv0iTrKnqc4hDv1al0BZOpifCOd
c0vD7qtHMMtLdGg0Njw4ix3fQ5Dlg3uzdcIx9dAzfQAs4khKv+qpd1MLo/wxdMornAly6EZ9GsI+
vRLc6uScxOsfCcGXgoeMMq4ZDmOObQ38x+oZFco9uimTzpRJWnVSYGwK4Dr6BOARWsPmphiO89l9
c2Qv+J9fC+5jm2t8KHuww5wMpZPgrqgUxUn/Duhoy5dQEka4hRVUe9zH6Crh0jUgg0xDk1PVhs30
slWW1M3LhBgnNIRwTESPA5QBWNYHEnj9G0yryUJuUpVaZevy+6OhtfX8G5iylnOGv3GB4sH4WEmQ
pJpRZ3DRZgeoiM8AM4DZTRhfa25UsRqhuBxTewGuENjBsBzqCmp8XPfhPSW05t9MihtVsPzSGjcX
9x0zB9LLIodQnVYaMM7IQ5IuyVBHq3JRnrCoCkgard9Xtkasrvj/kCxPtRKYo+Zijjc+lHeEGeD1
s4fiZDXXZYn3Ub9hW5KVEUwp9gwxjz8yhtCVv1oB8hDnCTZs0ZRFzJN4CBAL7IRzeeiyNzAobuCc
9X4qYcuXWG0d8Uvy6t2+d42LiPZWhpgqfdVbqqwtkGdBTahzbtdXacnQ1wzLT9kPfVPwlGNgoQ49
7WtQqiHj1vK1JI2OsNvoXwpJspdyh4lw4wO3NJ8v666t+OPE9Q/iq3jxzC+hA/MwoiP2pB3NWd+L
0PfTtZTM9WNIk0f63vWSYlv5dbijx77lWGmWJklzgMgitkmOyx31XFKrJJtnITELTANmU7S/W6eJ
vme9YO+Xi2f5tYD5LPMoxfDrdvhIuFtucw9FI/23GmVi5RLJTf6pnxa49cs4UNJy+ddy9hC5mDjl
L3qVBH/Y/DducpTAmG7cKVUBaYfWebC/aTygpmtnspKrTLP65mkfm28kwMYWhqrtfQM7WFU+khSr
b7iZAkNotkg1AocZvAxpluug5g0xx5eQjEqyjguTh0/hPo5OnOcbZK3w4rTv2G58M+JZrXO1eAx1
sWDbKDTTfyy0mR/mZ532wVnaLViEUbQpgAOusJ9G9pIyFRa10EakpuOBCnvp+K2IrkPTOf7Jxbnx
7KnLJmuq8Dxf3yEKJoz8eLaxbKH7cGzjY58rb+jOmeNG880cz6VJJSFJ+4BJs4dgScJq/XFmlIHu
/5kbPAOrNFPeIsSrOVgTXQLfkvKqvT1VHiSFAAzWvrvkfLrFDT6tSRYdTh9/tK87YnB1DdhWigbV
fOZqhfGEfs7DKLNMY647S8L8jGQF7gx3RRF7JHKToaXSfgVXe2NcW5OhE+4o4Gs32mfAABIZKqLf
rW7Fbz5O2NqG9adIuBahgK1m5XPGrwyHOXHf5/pp840bnSBaPSFM1WHWAkuAenKsPyQgafL2L3nc
id3ONnuBIh06r8pxTnUNQz8TSB3n12gTCP9MGi8wKgQyciW+ddNIlCj7uMTw1I8l7zKcaXw+TE4m
tXQ6rB2lchYnstbwooT4RB+BISAjHipoR/GSRVmTHbjdQWOyysvW/IVLGt52YFB1qbPeltXEkWYB
jEjFvZ4nqzsMqctTRDy9dLxYrBhjZTNIYqHHU58pXtsOrGV4qiwraGRo1nRVi7CS1f1pFCniIoAx
Wpx6bwSBa62Jc7gzs3EUAnrXAiIMnkcgfleuXyU6mGCCIjX/kxYW/tuI4RY5+F7Cg+eaJw4WuzsN
Kuj9TLqRud/CBcyKmKFVO/XpEvrTpJ0yLS+2nTBHoVwxNAQTbXp+4UTq+Jty7ErZhn+MPU0hBtA2
71WNrX7dpAKoHPorZuAaOuZuEREPF6hF/1rIUXooE5l0iCOiWhazTWnDR/IuxaKJMpjQ+8/wroo6
D4hh3Rdm3OVVCF6s5HiW4i6pj5vJ8G/TJjeJ2sRcXV3uIib1v7WBzlT0uTFzBagh+lIvyGNrn95o
crgIQMQIxhVYDTZe5jfnEMBV28JnoA3P9ItXAg4R05fNyTjuqUulAZ6egESfeGXXBMkVU5n5HRKU
XeshmERf8/M060aK98RveHm7Bb5ewUw1hCZXYsjz5MDqvFkP/1bM+62TMZlrF8rjFYStO9YMLzZX
R3q26iJshNC37uBaYU+WwnRVXQEmdKgKYGldd2b5HlpJYRHzoOgOUoxlbaaufv7zdcIEnGKLj/0K
xC8SIhvtI9RBuygCltOpjog55S3p9UF3hc7wj4jenutkAZlSdDGjDOKbl6SVIj+wNDQPGfrNvo0v
tKNMrX6FyYHCcGS76PQuedJy0B0kb6I6f8uqFvEmjqLPSg5NYfUBhIv8FgZKVcZV3q+1J6FiJJ7/
uQWTxiLPP4eRcMM8nJnTw7NyZC+KUdgegdWW8K+to3wRaj2ahKlj3AXwvf7MVIw7O5LbiqI5xJQn
i2KmaBByccmiiEOXfwwMl4ssvnr+GKCz0gi4388nrmFM5Mhk+GdthfAm9tPwUyOFGNn4mbIqcPAh
J+EyehYH5wu4B8pfCAktvLKgNzZzSxmM6Kg0afngdTYZjbSzMmnMkbMsdmRCfFe24qQw76HqPf6i
5V1N48dXRtOZ/LhSNUfbkG5f7tq5P1ct2w26jZGLwTIBXNwFeBAIsmiv1c7FLo43BehJMCgDyYYi
DMbeYfOJUc02KzBzahOBVW0cTbwOuMaVQ4Cm1Mqqj85ff2TdukxmomRTDKmFCBh4vuj1C+FDFv1S
F9xO5nVVCceSGGktHLhdFO5mHpq5I+lTKU9jDeFORMV5AbjSvfDmplS64MsqFGSimBC1dvxs2Bop
U1n/QPIU41QElwm6M20v8rHi+tuLT875Jx98vyuV4CAAfkJVERkKB9yOYHhH8SdIBvHiBwJhHRB8
KlT9LKCPzcjUlSxjmTg/5q95U6g2Ge1SGXrsVPdZDPESMCshXfCzToeRhQwJ2OYW/YKyHpqiBSxH
sRlCUzzwF3Hk1AJmnIsxidBsDjRfBOSeiBPB5Tuwdf7kcbgwfJAgypHa0lauUWsI4Nr9pelUfmMW
mN5RyydUue7PVcDChstT3H2ywpuKiE63IY1sTUFlm2Qlu5jCGtl0iTI6jWvwQR+DIQywJlDWeCrf
IokdZDJq6THxR7kcHwd+/05c8yovsASEcvP5NqvTBMTlhGDw/mAQv21mdobvSV18jm61HrroL2k+
YQfZxgYjEBzImauH9P457/iJGKrINzmdmra6XLz5MvUejzI+xYSD8j1CjVMgJ88FzvSRwGm/WOwx
VKifbrmIslPBMOhW9/jI4xuaULbkQC71cQ9pP/NI76a4K9imdVAmJvpi4S9sOELqwDABxXvcfz1r
iLwJGDIxHPeA7uuLovZbxmpRLBw6ZRPVjLXbAKEvoHlSCYB5plyOGnO9fPRzB+A7M603i2SYRLIO
QUH2QTJOr2s+Lz+YoIeQFi+qw+9U390N8DR6Dyj3J6hT561wrmRfVZKCb20OLRMHZ66+7OFS3u6y
5U7KlAKbZAu6MrAkbPqUP8P0x9ClKdYdiRtRNas7jkf7KKL8qUuCoYo/Kdm1KKFI4HOS9/z4ySON
D9OjlEI4RY/B8IlCnES/6aoYwHR77QEnBJ/rBbtpELGf7grB+eb6yr0ZWPcF5uYcpiRCGSydKXY/
IvKGPkyfhVyaOuf8vT0/+Vi2KOS3y2grXaCj0qvAUn4dDII1IpePW8e1Rt9RZk18s4UPPnuqoPdW
/l335TuWreKP3PA4W9Zdm3EUCCrG6EAYlWM87p67J76ihGnSfvkzpZWqBJt4QRD1+bzj8IoiteVb
ccIGP0mO4aL2jCOZeraII+IoI5lQIs3BhKKPsD3IQNP3Sb5lFGc8aIkdCxumff4yE7B7iYDHoyVj
30IeKcfXj7PGoGctOPGIyCTP3dgcNQLN6TvHxGVCLE2+dubZB9jJ1DQtkR/F4zSgSOANux/lAXeV
4UI6WTpyJze/552B73M7RHyUHBQBDC0/3seVyb6xqryNjxtcRHuYktNno2hmlsccjr8O+ylbvp2l
MtqOewevSNqi/rCmUP7aN/TqJxDChgvnuYGkG0Nv9ki+h35kDaVCLNpGN32a6u8Y2a5wdvBWWAv9
d4w7denfxp1GLlHKp1om9cJqF0AOYjLnROWnJvTAvN++Pcbf2U2FrkTP1cLFqoLGLyJKL2dBFzSp
gEZINTbaYqNa6fz4oOYgJe1AGpiz6mpIIBCn6iPKsyOHhys0uuI27jVWBfm+2u+JRN1luDMtRuPd
+NLPHDVqybwromhVAoSs3LmvZBCFfQtNBnAUBZDXQP8dg++KXIS4//Vw0aqCJwF6LLMFG+pAoqk1
QLabOPy3gjFQ+gDbPqUlYCYStZmsYUct98zc0nCQb41vRSAkSLAZfk5m9OTWaI6EmsV3/xJnmnm6
tBo5ofbZtCXp/t4+P9QDfthZ5kK1ZrAO1lmXHRY98FQ/8QuOMbduHZEETwYHZf5vnb1myE6D6KBe
niQDvp4cSPWhF2hkcBQ+GoyA0NfwhhtjJ/5FWEXjBoyMMJ5usnrI2xoV6CJmXqbEyCYLDHmRVfQG
7Eq6nuLfGcHrcTx7c9sdqBFKGbhPyAeMg08PM449wxA9VkziW0+PuZpJzv7wdT0Ua2ZAy2RLvqHY
IaXEeiaf7ammt9ltKdsr8+qQV6bZPnlPPa00Qp+BnmH4faVBws3x2UL7f0w1V+dxhTzxBC8+VnIU
6WorOA/Z1L8kpJs6GdunrYANVZE3RnobBGC3OjYpNbdWxF44zPCOfpobDHqgaBu9eQuzjj4+tW5G
yjAaMvYZfHVaOK9EyCP4NHHg8Xs6WBJxVURWqfFxCb9yHB56AnjXHorEtBVYA9yfUP5FPh2yFy1V
iuqdhZoWJaTEVhzi08LSuQgF31ffmVY2nnGzMcT/DLSJVnWLe7Kwt+kY4cOjy0XgbOmAADoVRmOr
EXEr6p3vtLqUUZTz/5isJPJ4wEG+TGR+rZr6sNY4PTKOF7wkJkt6oMw2aBh0y4YGB4ZCl3KbuW8p
lZDDTNA8KK4o6yE7BqdiaGYq6fbG9BwHUDCEY1Wph4q/lhTR1nXRwFUEf5DNq/Nzybn9KuC5T/RD
i4XvHZoirXxweF1MpjWVsvbJUwYOvpzI7sfNT88CB7QQ7VUKGu2bUvmB95e54wQWX7DH7id8VyId
ql4wCza8jCKbG1nT8xZ6Wb14MT5u2i6FS831XWMbpRIaGBBRNQaBqV8basoiM9ksPMUt91v5mJsa
OUI/EAunkicespEUYi1N0rTawCVUqxcuDJsCQNXftiZFx4R3J210NPWJNbE5gTtPHuQlcEl+Ai4B
JMK5nkHT7cJ8uJ4PrFV3Vg4m3CkmYMRFHXovSBYcV6L11OuGsrEAxrDNjjCq1yI3AY+Af5MOAJfO
0sjM1/JuEyhutwnaH09ahorP7IRWBqcduFiM8tSV26cWu4vZ5SHPp2V+/LcrZnIbh0glApbd2C8q
MwC6ymm6Cs63OryiIkeaTHLAG7HGdz8FgxQemVUhIxwZ2j/5KHTIB7oEPcHhT7yIiqpTjRtkC7B4
lT1h9XCAO+El24364OaM6ii82fwPY1jL7OVTsmmWvtT8jazW7bJJezRk/T+cho14nmAp5Dx3++eE
VMH8HY6J1QCWSF1l7ikioy5o7UtwVjTUFfeO5WAS5RFAHUdu/wEDH0KtXdrkQapNMbc0ZwJr3d5D
6ExMdIIBQccQXZfWl6tjfbXIkWetN01XVQNkoXiD88mRjZPIsW7FEgcSt184CPoRwuGy68mwYBi8
oaDbXAF04v5nYhLzL0kW6UdflXfoVtj6W6h8q4hzCk8hNf5tF+GqKyaDLrfYz3GHkR6xaVBjbRe9
zVcmH2nTkxhHqu/Az12Rhot1HycoB0420VXmsjvKYByvz5gFO268Qhpsko/V6C00nnfc1pz7b2tv
v62fHvxz3pIIcw5GMvIPqc7yBFagy9LLxXRJm3hNXIq2hVvMcEurjDCmqvGt58GRrItKtqTLZbcL
BhgRsi9eITutDRwYXX4mmnFVdMJI3PVrFoxSor5Q3nCVWe2N12qqjPCl/OIO9XKGMekjxX6993CS
J6PoLciNABP2Lnr5nmiY0aZxYR9/8r581whLU1tT+owjTQi6mfEWGYlnYUMSn8MT/GnIzMfCT3dG
N7Pz2WsJl/eI3RKRDJ01UqhBPNQw9IctKXAUG2vi7ufOhBx3dIB6AUKOMTiiNNFIEidnoHHCJZRR
My4kWu3whX0LOarnmwGDF4FRn4qxmaX0IL/vyfw/HniRaYfphDO9rKYjSXEX5yhTSTnqV1zkxJUg
UXBFhJe/eqlv4fkTGox82DSuZGichjl1eYq+Nl83DzZ6qVuDcVqnRhYNZMDZev2vP/Z/pJN+A/t5
ruWJDdZKhhJ8WlR+2I2OPKK5fJtWOxfU/XNLPaUorOSn/FYPekSnkwu/CWuGwXEqgEzp43MtvsvC
1pHFI4p5t4BQSXqIZuVG9QS8L0tcvm6tWBJ3wEj7C5cNkfnVZ/IJADjPtfN25dzmi7Vb/a22YTPR
EfYSDhse1dEPOp7PA8TX7utFmxerPUXbf6nCCpWHjoo1Fda7t5cBi9nXo9FaiY6uRJeIsPhgGK0E
EzO/LIWj3Cq8CFYq0CFoWp176v4T+VabbN/aaDpntp3Rh90N65b2rqwDUwEbreU61byVmaQbi2FH
DyYiankvFH/mjnw8Unj6RbkJR/zIKvordm2iMKwQGQbUphXeoYRM5H47d2DkWcsTrzso3z2RLYLr
tbK7P/JSS4tRHwcS7bkbxBBZnebPH3dOtCdHdHHLrQXxshRDTq3de5eUrPPcRpJz6n2sNiVya80O
d0o1X2O/jORZVz6zLGj6USPeu0NXM9ApR0tjYQ/q3IcLtH2s7ZKsWCs5yiVRUmWNBZPlRhbswXAc
n/5LpHJJ4Nx9yFN7MDr37Bk9DdSeb+kfjsYh+TRTO8d1BHPejUAyX24T/PIS+8ab+dUUKcTVRnbR
BxbFaVABCOteK51Q+blX4EQ6LTGa5xxzWcIIMxMX6fPKbwID1CCXvDEeXXFxK7s2xldgDD354N+x
6n+h+3cPUiPYuw6tgB/d1pouHA9EHFcpd7gHyM5k3Y3DtHE49maEGDfqSZQgHeH5Zg2O9JgBQnuL
5D+oqP08RF51t4PGblQj/4GXho7TL4n7stT35RoekmmyTblpyGiqans5a0KJZVKkqx48HzJ/C6jN
RPptP9Z746lJf1CCvsfIoQBqmuA3Uec69G3TV1kmZm02/BFZl1i6yU1B3yFg4CrRPs0k0mMDLLwb
46Sb8iqp8drnZVmhOBfiqMh1V5WrV1z04du4uTz1RGtW9Wal4aCzNbvSYwICMUmW11Cf2JSSjsSb
lei6Heyay7qkrrd/LewXF7vO+i96WvyfSx0LssBexuWDliOXSLCb0pwul3VgZoLsejTUgHpUumPx
MZN7ulX5oEY2Bmz/61PmbcQLltkctZVh2xvBsEpnYi3XqeGayIuFRGVO2B/OgmOFyrgzTlM+/IGH
Ej5u3NapT+jSA5hI55/T8CyD6Qm51hCwu4Oyn3gmM0dXtoBLq7j0zPc3PBJjEyGRnemUITTL07SL
P2wJsmn8DXknqdzWKw0RChK9MmKt4gcp4MllFMN5XPIIXTrQva1iQflC5g1ZzX3cUhB7AWoUNzaH
9JDllbmvSICIf48j8NESxuLj9zkllc69YEwLLzrGobe8WzgR6Dg6Euyjbg5AGfSop8CNXFhL49cw
FojLUDc3UURVppLhOEqiOwIA+/vKyhQRCUkbevPbXnPtXSfUW+YwB8F81HHuo3XB8sb4vq6PM3VU
K/m70c44aFgplzkBgwufYXzaK8m0hsQ2Z2qtDahLsT5iFpilzAY8x86O3Z2HYArc73qUsggzz5lg
KvLzHFqokruvP4ecVgz0uAFca/92nn9bSmxqkU93GTVapz0nEal7FqIvln1kawH70NWc9OBV2f3B
+Ua00gBaue402cZHedRhEhnd5g7FKRhZ7RogUFF81j5ctObWe96fd1d7HisrIzH5Rd1bediD5uys
vihR3KzhQuQ1VfRJfyPZJbRuiKX97VIk7ECDpLFLGSj5V3A4EfCjU0MzO4PZ+xNBB204ezkwnJJ4
8mJXgz3W/IS6YoS60vnW3znYGe5u/NE0PH2P39Ay1KDSC254o6n/J9s0maqT1Jc1Dru6/+abnapZ
xGndyHtWu0uAs1OomAarNAdodTN1IsV8Jvp5PU9Yu8YCJninFaGRdC+LvFZCzBiorgLAW6Wrid42
C8gfkej//KOSUR3x6udfKQm3TiiQreUpgj7p77Y63dJexDGw1TQBdHj32skFvstw+7JQvKOkIXHE
7zHvwcb0gbaI4x8gWptVvOU5v2VAqGqQELHwL5Tly3GQMWLbYGPinlpdUoPKNCo6dDDIbk6ctDFy
+B94Ak3xEN3bwtMGQLPp6GedrV6caBJ22FSphELLZjjZDQ7r31aWYNiPJxqx5wPjkuxCX5zxBAw9
i4W5WYTyDDDEwhFMOWQqQq4ADKSRjO/uLzzKmZ+tQolGYoCwNvoPurKdjs6/Nll3J63T4J+obptV
v5a2otNzyhcf6+f7tRJuIUNkLPOzv2SGJzk6IVVvb31ti7hxb0lKnzqS8Cg+uR3wSJixg16t137L
+401ZTY3lDUQcVP565upZqGKYVd5YjhHiQtBRWZholieBcdwbzybC3D/KxIGaRTLX70QXsAQzxt3
p3Ljp6wkcmE93/C0gszc+mWebatqL0F6Wq1Pt52WqQlZ+Z723i2uwnF9R5q2kz0Xa4z53dLBVBAS
L6zTTxz+fjpKl/Utsr8qj+uQGx88BIPQLZlMhTdxjOUc8lZzetgTGsi6a16CcQY9ip25XJ42fCCl
WWxsfHvIKvFV1vvBbeIwxLbX5RTpcx+fyAnY9l4C4UH/J/yAYQD+rjokJfu/36zotbTYbFR0zf5Q
Zeeu5Ao65+5ecfNzsSO6mMxSpMZRePIGvqoRJaVQQXMkBSdZlWhyUsY4HZiqRTKeFF7VKSO9Wvg4
hrNRaGIbLpzeTU8cHJpYApRjEZJRk5NkiOJQJFAX6sQPbqNcg/dPg0SdsBdGf/uwVYGjRNy9oTAP
ghyvqyA6DsQS4S4/DHEMWDQVvuYUekANSUH4Soosqi1uGFAIH0W1N0zDJxqddjTrcwTSH+D1vifN
7zqcwqufcZ8QdpTcNcObASl09qV6OPSt0O1mjhYvTJGilWQ4K8sFLgsws9MKZyEA6S+CMz+Wde7w
/zke7ISL5HI79I9RBGwsivLIMzqNoqII+rIFkBwJL5u/G4o/xfWYIKGOfiOAzUFylsIKNZjoBl6v
06AH1by0O7HAYDu/GxLfMOa7PggaJ33aw7OfIerqTW0qrmUlKY87XSEUzUmCsczVASNSfoJW4ocz
rH9g3YpxzlFBg90PJyeO0cK28Z636Ivai9QQb57oIg+mt0i3VK559FEw6uCOSpCkKj97zg9kBmCQ
Cn3QgyLgSfT3VvLOtX5/5lZRVLczOcI51ubFUR1Mi66L8iN44Jv5+n9f2b0P6X7mXNy3oA3EBhR1
RfvqJ9NtzodkgZsq96m/w6VRAR20dFK0LE6/mIEhV7276yty8zF9tjbRkl9isYwDIrxcxvkYvyIb
6KXspHzt2CNcPFMsY20uw3yvwHiJg7Qfuk9t8au4fLyEK9abQ+xhHt+PKKeNLq74JL9UNG3+cUDV
dI/RAs0bPuu7fe2MsNdsHqtGW8hqVXmGIg26FqGKcyTnwIkuXfF01S/oopzN5fGOdALY5JlDZnSr
ABYTCw3otxf7/788lRdnw+zjg2c2Tc4Uh/8TcbBaBcElWo107xD0MRxagQHPBVut1K8xXNYDaRPc
DnUq1/AcN+I4Xzu7wS9dEnkc919a2pQhGdsdUz0TGQ7pBsPzylEJQQ/nUX7E88ZTWy/NA+5W2nMy
hQuzVTbm5U6N5dleqYo1bDhnnNnXIBXASPAteg5hSNxM57vQ6vJMsrTcwQhvvE3RCoPvA5jenkNU
/7JnStomED56Y0511U666odzqJIqM9llmCHWVq7Io2e/PZe27nDT6Q0m+87pyNAEfzf/3sTvZeeo
5jSDT8tgkWVrZpql/o01suVOPG5hQvfPeekHcpX7XbogSDcOhA47iOXWQWS129YWYis5MmdSWol6
+P0qf0BPskHVPObRTbvN8MDIwW2z5sVuf121wpLBhksG3SXKgT98lspORER6t+iILr0gutnFBVV9
ea69TpIyp62B8UmZ10ao8bpthKx43+enLxXFbmn1G3/Ph4/k3bJTths09kj8hnSBwv+AA3zP8CSp
GhowvhpNhrSth+/zptBxIjpqoh7Qt6JJiQtKrk//JfbRX1LrA5lE0ahTPy6KxgzKSp1uJdCGBKCM
4/n0T+WvNPc8eJsG3t+u8OoDy4kWX8mPI/SbgxZcGzml3nFiLnsF3rfmC5vJa2LezfzI0nM0R8G+
DAGJBTfVTl/K1tI/eVYE2kQHAoDqprtjbFR81apVQ+jOd37DuCCLhGwP5DkAXgBTvqhojDRrQUkl
g1ASO59BOzZNkkwvcQYcR3SEO7UewkdwlhlCr23BQbDlj9e6JxVtvutFU/GSwH5O8BD0L/D6oRRw
TpaTc5Kc29Eok2Yi0HyrdiiXHtFUsZlYUrMJtrtB7vEOSAIQKc6uhD6VLvO2nbnl8YWI8WfDtE9M
dK2TlNoaCFE+yRVI3/7tGCfqW8dSMpW892YXcIBdWFjw4NwuhKJ6DqkL+BxnWZriDy+mBsn1F+Wr
JGXXa/EpG/sgKILbcCnjZ7k2fxMQnFf9kxahR1lDOUH35vTYLT1TZKib9iV0H+mXoH/B6u9qpHoj
gFURd+rMAHpX1ywkcSsrJw+oD9aq9tYRLWSOZyAmeDNxvqbKH2ZYA4jXeuAVz9gjCO3NbW2/JtBi
VzdhKKmK9O9kvpLlroEtmDEZosvd0t0ohO2HnHga+c1sIAk0aSKQslbNa4qNSFKLAp/+KuSb6qtu
y0Tod669phGx3eSeTM9Zk/I1W1p2PNetfDUynkMbGpWgHOm6r5wStSrL010ucrVuFlaKo3LvhiYJ
XxkBTL6ZN3euDTOFUntEPJDMzQ+DC+aDCC6QrORpW9aZ0375D3yOmj8qQ8cuLBXU2WHyP9H/GDol
pBa+e2m4iz3q9WjBZyYOG/IlivYQRc0RbLfVMobDMA5l13yLZkBgKIS+rA1fzLqL+kfi3Wute87d
IdhScrPM+ay+F1AFlvPwV9WhTCS0QV2CYvnGzfp5yC5h7T6/rt/zFiNAM2JEz3Nq96Xo1w1joWQ8
nM/0DuVrjROSqVjCvOaZT0G5S1WIvN2yRZxtEUIW/xyk7ACmH+Dr3w287ZiA0dnnhSjNnbsjrn63
OOfsbPcSdw040YowEgWgMCOc9/+5MdnyIbg8rElB/GYGlIzlm3DzC1zy+LKmX4EYIyHqKLEhZytb
+A7kQq9L+GLVfwYsXu8bdSWnqo9cZ1D2gMGfMF8AzbC+ieHN/XzHRchQG7T8YttOFbRe51zfVNOI
I+Q8Xfa9rZqGv8YQbdcSH3Zxkpcpsd+CcmS7tAyny57d+OSOtaRx+Qb7/gZpz5/4PehR9PK0sAsY
LvjVMZIUQs23EVBZwyWMJYguQTh9uV+Ah6RaX5RvTG7KlE17pUeTcBkI1G0tK3xtAHlOTcaOO4lw
YK3CbKdS15j7hYjdXIqzwRxRIVah5HfSKHprY3/Wxp/lzbKczxH5qM699OsRMJNsquYmZoancFhD
femMD/KIIvtw+lfbrRrCVnZmWFMXVn9QX1rmoINu/OQhuKqEVThZzsy4yWnwF3c+AAPclst4UVNO
t/3sdsgIDxhVxKer/AuQsHY8cybLAJz33+DLsZ1aZ4a7lQHuIBG39CCdiTVU+SFpaackNdtQbgn0
/TjaIVGjglci584FbZ52Azk15nY+OBiSWZIWXy6mS3B5bA+MKAJeRaeyoxPvm5TayY/6zl5u59ot
qFkZ97agF9dFwAvaAI+Rbm7ZrCcatt7oWUeh16asfeL1aiGnrecOLiTpbRRPsbH5c/3/IDoGT8qW
shS2i5gYsclsO+pvp7V2BCAzmrudEo9Fyb2foCLNncNFfdkhz7j7jFYEDAlnkBMH33lxD+OVl6wX
ZsuSvsxeVIjYnwDd7xsoiFlqABx3llbkPAdhDrn4gvl1EUMDOTgWSP0pkw0jPFwwX+NlRcEQdD9E
zfcuUd3jruQOoRxoe+YQ2sPN7CgcOaFwQJH33mEedrg4JxtixC72JRvUUdCcRf/f//Lpeb4kBT+Z
od0/iSB+4jtbVYnfDMMW0E1LxwCTJUhgrdeI4PAj072/WtvGzlEFL+sBvKuqErPqU72Ve97laKIP
phUhWM+1a5jrvcmwWYH3KdJzY0/WyRFzO30MKWT6QPK1AuAQ71JQ7rqCaATkIQinr5vjlbKtjvxV
q/c/yZmBVFPmAjOYef0XAZl8HVCSGCbUdMcJd0XxavrsIxgxcnPVpODSgX/qvLYORxRBfMLQG6Lh
Xn6xQ2ssvrTfzDabiOHjRGNmBJrbCTljm1+xfBnVaK3EgFshOdJrv5d87Au5KweZJH45rPODhX14
5M07KGfuY1T2dRr1HGYRXwnCnq8SikljZCPXqbQUpEUHErPOEzSuPcneycxTGvDNz7+PLo8wyHUU
G9kMGAfOrV7eR/oZ1ql8Dq7ubkbPkGsoFOMerbiV9hhTdXzWJ0XBvujT1aU6y7mbLU+TFKJNFVx5
OzfUR6qnLq7y/DLzOdynBoDQFLyxJejO5DS8si20M1tQBWz1sInkCXmJmREkDU8TigQAH+Qmb4MQ
WtE2KDoZsS/qMRSA5E0oNvgieY+KOkQ19Xs+a/W+Nq/Y+Aw7Y6Vu1XE3k7NpV0NMgKVTAMwTyQ0U
6SsbLTPTDXgOqq9bapVhca2IcCVSrM94fHeUvyQ+E8WAquG7/fqW108+yoqI04b2gdaeO8R29yKj
OZguFTFoW+XHcSoblPGJVNj1yR3tTG3sMPYrPdpYlYWoMfKxKD8w0pYnxY/VUCzzxf/eySoZ0GK0
hgCaW9VXSJ7D6Cq8G9yGDw6JlaPrMx32Wk++LAf1IRdaIDUT3ubRvchUQPgU7ww/lntcz98e2shy
Lb63fwlkbd+atyGz92DAC+us8fKAcm60AEuFKpwbGK/g2HFkkXvkHWRJjmhzMyIJFxocbSDukM3X
64DCvt10cHIa4hi4NPz6EggvusPlSU4FGmFmBj0399E6XqbFPjg4vq1mLRms26T5AqRd7Cu0XfT7
sBW71f9I8WbzdOjlbF0ojDLcp9pPXchR1ovJ71Ll3tBe9eki7Y1ol9TDc3pt2gNxE1NIvUuiPBk4
vAuYxkyMGBYSUOjwYaNUvckwNwDITgJYIHK6mArkh3HdZocWs0v4/1AaS9kIDbMWDpXUiuEVWg+a
Qz5IquAII6uB7NCk+IYC2hvoXqUhqKfHMcGesxdU5zFfJ+VFKdoTliJcW2FaHJQ+cgJz8Jf19PQS
8ROpp6bm2xBujE8MU/8wRjLUAHpI+8VOwhiwGILUxQ15QjlAKP848vhpt0zESKNOCrMJNJG0e6iH
ysdCXbz0fh97mJDFfoJ20e0ZGIE4/h9DPnXXhNBYLxRJiumbnS6jJ8spFfaIQJl25YV1dcpHCZ9O
uJkHC1B8LLjy1WyEPeZbSK4omWgoR/1tCil+BRj/xHYy1zIN7S2F7FBmNBBmCNaICWmyCKvD+aXH
OlpnEuAm3vquaXkjYMlkIWOQioq2pmH9oyCDVh2qP0Wh10WKZgyW2yDh3UsnGyroVXscMTsdiaG+
UT+qoRUCwjjftUcZsF1lM6izywCorl67TGHFJTQfnB3CDpWudzTVq6GhYUQn4JrqYKQ2Xuhj58py
oS1SQb6+Uqs0Rk+MkjmUeFsijzpOu5UvI082Dwv+MSstE1If0HmqPx8S4sIm31z5rvw/hxgMV353
0cLVk0ijv7UAuTyDucwJWWVvjQtBtp9p20QL16g0NKqajiBex6AD3guhUb0EX8+6bYZtcdklHqqE
eGt/151shzdiILls3y/2sM32Q9AKLVz5UWkRtG8A5XDdmAHHgTrdUdbWOA6kx5VILcA1NmL0xiQL
O40xShh0s5ii8XnDVFMRnWHzSQhyONOvG3AkIHX7QEoYvifMxmw07hm8VvD5WCcEL0MJSVJiLzvQ
0xcpdgofK7jUmyQDx5PUqpqI2rhl5RsdK1VFqQ1fgnuPbHWble1LXPVFSHFGi/5UvUULOo8TQWMC
QckDVjRVqD6C/yIbc2TB9kXoM8RTKWmA5YZ3QJwDztULuyvp+BPirnR7SRs0KqJRWG5OGdAMgcwH
Amsc5pxDk3dmjIaV0uGOI2D9R3vQLOt5rN9GH2W+GeZ6/DIQc6AFVqH2g8t75g4YwAEOYAB2bUys
+Bm7GFYoW3annxYjvS0wm1hF/ULLEaf4FJe0yOnySOqu0h4zQXDc/TmRxw2hRgejJWs4byjs2MtF
9B5iGTpCx8wvOXKHnQBdBJgXNeUM/DAUo51VdoKmuKIQ/Z5UcWLIg9hcw7PKr8P/m0iwt3+UjdZ/
GV7sP24NtlJ1CmClCbu5MBC7goJDRgrUe9h3NCJ0hH+ZEkMqA5W9fIFHFSsECZEaXAoh0/6kyY70
e3ibJ1NcaqB7vsf4EPjLE+Y0pjZPy6EPzPvYgc5M/F7K1BiI41eO2qhcmobdHBZqh1HTNRY1TYVT
e7RMhGDsyd8wOA5+VGc3EAVnw24GjYOXeGWN0KtkoY7Qi+MtbbNvQhZUKitdSJ2A6La+JJXlJqZA
KK/DvuwYLa2QumCxiUdxMTiJzHLLGqraWe58cIfm3q24UiWJiv2EIWxfPwVbTl5qGhLbVNZbMC8y
0FlNI6+kTSZzGzDrwjBSkysVU9NliTpQvLNPMBu3rLCTne0hPwLDaNQCpgivNcK5KEpZLbhIGeIR
tKVdIKwmT3xWn2RaiEpqKuSz4QFVAlkrMNbCi9LqsxHUuQ7VMje5v3iKljQMRnH1B49Qdvhvxe8z
z/OmFWnpffgsrdZS8v7/U8ZEVQ9jBX5l86EQ88sTtvzVrpsSMOzgStR2FE7totqdW83vT9AJB6Zm
V2rkd7/WACMwNYmDNSMCW1AzbP+2nNTB/2/nRNMdKz7VtRaeaRtlGDgl6voqEz010HLOWvB69Jdr
0xATCgxJ0ZgsVG2Fu7zK0+EuxQEIX9T0jjG/P3BjrJYNNn2jNuxdF/4RkqtuYG/F4XH6QxkGeEwX
5N1JbmRXq7azB1C1VRPVFmLwXftU535dP/4V5vBn+k7GzsOgIb0+7hMfd9sioCkPitGWYX6ziLRl
OALU9aaXPGQjnjQkFci96myI4C3mZqSu/Dr9tdB1N4lkvpsBvH/IH8zU7LXVt9xfPjU8Fjtznq3d
7bN6b00mOdi7QHSwY0QgZ/rv5vEQqAh8230WHYqYjpIAlVRGnrpv5Ky9FKlU9PjhbsDA9FQZg9HF
zdcWKrwKWw0olr7w4gYFaIhMQZOsqp/rGvIjce/R5WBllFieZv6j6XbohoFEIRGs0zoDfO7KKp8K
F7dz3534S/FmpGudkFuyts6ZHwZbTLhnCoocZJrBU1k27VLku337SiTjg0sjahV1pQs/1fKG82yA
1wiQgyBiGQvIX1h26g2+rSnCVnOPDFFm4QVUZM3Uza4X0rdfFFxzm4bGt5scc5DNgFJaYnHohHsf
uz7Jpn2tfkxhKuZPMIrRRxDNehfMkhnoxwFRZOVKeoGkGiTXc7qhsp5YYDBspy4juvGh8x2DGNU2
xJFR1TGDgUQIgpUrZDiliNvcGOeg6EXxn8auOfys+PxOhpzu0r2QV4AHHB0JmNy8hfv7/G22fJsy
z2sNjsUOiCX4Dp/W10o4uGvRjLOdK1NGNlpXSN0iSlWp8LA0Q2ThVGQkvMMQfl87Dkp01tUAhby+
/K7JINEtz5e/reWLJn1ZX7d8EwjvSv6Zr/2/WxHtH/8x82kAJUAdEAu6Q+3eWT7LqNpIHPB9/VnO
VX6sKZv6ZyuZnMkvH/AKX4Uh4pmFuktKwWSOEBqQL5NiUiipRc43dtT2V/4iVsq85PH0Dr14N/TT
UhpCKejHt68a5GvAbRKE+6Ibp0x8ipetxmEk1h1nUMLj6sWqPM5cUB1da92q2AQYTkJzbQG7akZP
6QBCFPt59a+eSs0e4ZLkHD7zEUF1nx0VZ6D6hwyXyaoNw0yqn4SY2WvZRq5UyObdlFqQ7np6ufLz
u/bLmo+IhAgmc6Mwia8/cn43OOTFLwZdW0Sa6Wc9sfIT07C9JqoZq+AGN95SvGEs21Euf5MmeI/6
/pRXMqFoFvk5N5O4sJzVaUd7T/3cTX+bVADfQ3ExK6f9i+rDd5AKgI7+rNFFu0AB7IxGBUv/p3Bs
t5zLOqfY/lqWOiem72pPr13T95hyIMV5lcEQzlu1KM865pxhT+e/X5l15j4t+dJJP5tSIy42r7tO
hPL7Xj9C6rW3XcKMJx46Z/3XCiRUt2wGnZk5cKsZIR9A+Ks2ADmv475lb0PFZXzSmaJDrdmqObZj
9/cZixswg/ONUq95xcFxj7dv1/dS2pcJTkXLYT3brzUjpcgQyaPZlFO/uRnN5fTWz3rJwfuhsZ1r
9tQmr3KINuH2Plm2U32fJ2UU0iLz8+cuaMzbe6vT0ED+y2tzUKfus1a4AyPQiySRWkVi4pO7vEj1
JFKarDgXpp7BQpcE3kWTA+r2auuOFqZb+7WJvt+pv8+YO2Xhx+VYJpg6hYccplY2CuPdj8ZVXvLO
scBpWEL4BWf2sQhk6Kcb5JjYX0bd5CmVASP6tgl7sEXb4/Bvc1YcTmyCIPEHEXNooJ81rhcI2P6O
9F9bl6PDOH4la2d1v/oeFEPWHFWUr/ZYr99QyhpKHe35iGfJQacSp9b4nmRrZ+sQ+VHF0SdS+Mvu
+1syDFwAfFzBfN5Gzp42/sDnEyZ1mCrebJ31d79aVjTge8YHYC/FT0YIHzQyNKf6ogFEblV+k0W4
2wpRCn8LGCivZxsxkkY4xhRaJXdZSwLJ2hvQKYezt4InpuVIK66TIY26/a7xmf4X7tldUUaByR/J
+mkc9VWHLj40D8kLHq3JfyThmb9djFOUlGdW8XKHjYezDxvCQGCO7/vviTZDikXINUnizvnda++v
ya+mkijOjib/nnNzwO+XRD0n4YypPQ8vPoq5bOZ9LyDSLBCW259/RSa/5Rk8QoYElmJ/Q5wAMQiX
CH69f11q1Dm9fnJC7LwSCXJ3XlmBki+juwXJy240vUv3hWstmWGFL2ZaJhIfpKDsY+0Mso0s0DPI
bsshr6JlSOkTu7MEADZGB1cvAzkI7fvSfAXuRupuuTQ1mwOgCx0qP4UnXWgtg7iTCm5XL3Kw8gVu
EK82kBOF1yhILZZFXRGzMhwLUMgqUvSlDVU24k0Ia97uF6j7t01PUWChRE4uz6VoSgW0iOfiGiGu
NSUeBzU7/Ds/gxVYLptXpFq3eZKxihxDlIY3WMxUc6Yf9aOz/XYB0nuu8L9vO36Q1B1Xi0qHrEFR
ZFd6iE2NauKyZsvXB+YToDfZAjlalpjCAdwx81fMN110f0GC3ORiJThKArSUgcUfxE73C4Fh6Fuf
b1s/dSld4vSpYry2kIP2VLFlkabUNrDy9MZt+IFmauWS2djd0GXWSRA77BT3IEDrJdRO8YK+rpwD
IoRone/qj8+UqsIZebITeND4QKZS93HLUh2y6Fg+vzo8pKh+G9e7YM+U2vXP8iyv5IfyMU3WpMnr
SX8kRJjXHqRz1PhHEzZaVDLOSn0Y+oi7nQtHOIED/gUDcCtsTThRuAf0vKXGo71bb2lEMGMCh8b0
7K5/M08Y2ncS1lFxKtB48rwWQJYwQ/2cJ5xXNMgDSU6HBOtEf2SrlPcGeYlF+3VcMnqO5HBJgtoS
DwQt8D0ZNZ2L6t/Ik7n09I0VfZ4ey6WTGT5RU05HJI0BucI9yEK3dgtRhOf2Ah+Y+U3rYDnFNXL3
hLuh171+w8QtTUK0OWe28bziczOZI0xnIZpyfBAGDQ1EiuK2/jtrslEg/ICOaIE4CICeGf6S6iSB
GhDbjpQd6Th0UT7rBVC9DjQwc+pKjl9TS5D2qFdMWn/2FmcLYlfUsooKXpsTb6mzlVZZP17vNkF4
segc1TorniOt6xmgnKzXhKUJm4KHt0Oos0r42De7uYWdhqyze6qjUBrU0dqbX0v+gYsCiMVJPig/
89+Q3QvOUWViVfGCQ+Js8tv+82aMLSiKCnIG7Qso6FyatGgJHrTcISnyJJ4F62Quf6LVWVU1wUmf
ah3YdHIBAi/qmIzKDhduW549nmpA/Ugb15I/ke4TM6D0gA8fdHCUA2ucDSdydOhKWRdj1CPlO+k5
LciDLn6T+wye4hcVPMIARRqIPtpHkA2Ydw2tFkhujWA/lu36YxpmQGg9KNSdMU2/EdOpX5lJbSc8
Lk1jZZCzIlQzF3an4iQzdJL2t1NYbZop+OVKNKAtFX8IcVVSQutWQWM5xX/ZJEB7E5Cb5RBnWRlR
iOsLpDxT5kRfQWYzQclB+W7a9gbXkQSm5d571X1pi9YlXDpi0d3PZ/IJfzTAJOqw5Yg9Q7iCV4P3
IFvsfSRDgn3fw7ta6lJxtQHwPFa+xorVKjaUtsF6qbrP6D22BZ2/71v+4Pqh8g3aOSix35UCqvfK
JrGv8QJkW43IUM+3ftODMn1p9GAf9HFVy6n5TvHhcOHV6m1y2StzkzSaOxfpSZBe45AGtIOOURyR
6ESUFsdQyKVk47yHEzWSA2un9AfK/VBtW6K3W8ECu8Mer1K7BVieZdPcYbIk5EwrLpxS5/rUmA+p
KZPWzFM2foh/M2kczXecu2bwcEZX6CehGA0nOR4qPTKhtPbk/+ExwszzPdZ6X+HrkQvKvMxxJyi0
0xCBRmtIziq+E1iM9gPRCr5PO6VyQ/5Rh41M64vWR08Mrzo+l5vNFYmyGoTm3KFwd3XNlNNuUS74
5luYF9uXzgXAefuH9Zvvo8Xqj4X29tWik5TMDW/O8BaWNeQdk6TpPVi3Uft4iDIw2jKJg6TNMMWx
AOaCS7KavHaOMnB5m+9WEI2XEESMoEQtFe3zwJKITkgDwyrOBOx6uuAYHdpg2nzNK+wEoUoYzDcb
cah3OoGBXsPcAlZ5BIddyq4sGUbrjl3B+eDa9rRvJL8VfDNJI4X1BkQqxmHV/LxRlHoKjqXLm7cG
31WMp33OGiqajtastupr2J53dJf/FyKEezNJt6HqiIZ0S0rrfkl8SyErLaSRJqbCUtQbZUzLiDcR
PfWff3hyejvwY6Lp2i/P7VFlCfXhuPKyky4pSqJltvbeo0nrLsSOkGvNjaHCe2hgfn5Y6mch8r0Q
Z4Qa6FaJTc4QADPSro7legp+PAdgEM/s9WSYfbpJDV2eNzseoXT4gJTndZATonWGUIXALJ8fJ8vj
hPQRHdXJJoxv8olPVLa7qtz/MECNHvza39nAW8zRG0ejPR8OhldVN9zqcrXOJI+OIAisre+KlJoX
8i1gBW255qFxxAB34lGPnwd6P8TiQi4OBuCIVXU0ID5qLaoi2OJcFm3welhIo7XPjEEO4rRAz0M2
w0TfWbRXm0rrpducxxBQQ+HCCE8el8+p1Ohc9oj+J4EsiQP9RK6iTMjzu0QIeYXCXhNzh7c0N7Q5
pyF5sB9el/Rnahc5YakjKpnU9oUVXXCcH41f34uHU728Q8Sg2ZB1WmeqA8eWVecISA2SnphUhNiV
mlAZM5hk1tlg64qatVb1yKn9vV5LZvsekMN1GKoWStXk5keM0EK+KQ8Xw8v96fyQzaJ5OwktAuBF
9czOVbqxEbwt8IiTV6hE+0PqeQ7NP+vIjLIa1isrHCNNANRziTDXnngxdwCdTiB+HKRRk2WH+AO1
7cUCVvUFt7iAR1688jcK+O4T5Z3y6KlojtSTzYE1k/4YDVT6k4y4MALloThyMseqy3lA5/MT3xA6
s1FTu0EiiV3QI8ZeouSUXmFhxGZNHwrKN+S4TZjWEcm7U4wb/5XFOX6gEIoZBGf3nQsOqCdkhwEh
hiXLmqyzlG8pYxZQbsHNSfTvl9MICYkCyExya3Heu3RIyM4UM+OH/QhCU/r3FoCrCeEzo1dnAUYy
qNHw3nzGLi9bsuKMRWkeCgoL1Bc8SZg2RC41tTlSDBc+W+22M7ILwKYyTG8Ox2wZJKizbA55/csA
Jz2cdXhppdWhH7zpcyT4/JQ+928PkfZr+nDH+util6bGVwI9wzlCfCQMcBYyWZvOvZObw49ayMp+
eMZoLIuQEsqOOoESbk2mGMsPkfrVkdHEG/w1C2Nxi5AAi5gzIZ2CpXe3JgSAUJ9t/+jd/Kd8P64m
m9yXN/077oH/S4EFckgMHHkcdX2DhUoBAUoa03PcyOGY1vLGyrfNM/0ZG7Cj8GCXJouyXsdYajbl
TbBQl4M6NZnRyGMzLgbhLTVfkribWAPVwLdfTbVax94ikXI4/wd4M23Spkp7QoK8LsitdHFwDd++
9ei/7ry1rtmO0kZ5CxIRnqcpkOtR6Wn2MJqde+CiPwdnAYlzMJfQOmFkrMKHKnAuxcQdLQTNv3FW
UgPFZMS2yWou0VjFDSnhcUYcKSBAmrS69vIeXWixgEtYOup0qGD1hiqZEm1oM1IYXexuajQ0PdbJ
75Ye5cOIGs0bmkU2uS5OVIs9CanngpKYeLQFJfaufIQsiaTXcCWsCi0Nn+gYLzGQUPQI1fjEasPW
HGo8lE9IL1svGZwBS+I5OtFgBWynN74MreYLlIElU2/viNaoFqp4Y06n8zx615gAmIVZmP6D3GoJ
r7SEjATRMPipNydSHBZkAwpdyu3NEmoC88+KvCk4j1nttvmIIoNqzEsNuXjU75bfRCaZNaKm83gj
9kLpOwgNKN07w1BJbobsiULOZ9CqbGWzC4Ex91yIWakLqn3IKpU5fN9WjMKpbU4PD9AZWWK9/125
Rp7aKdm3xOAMb9Dv+2Ys7EkLgCV3YLTl2gPjBdwaGjjD0ILGVGJ2szOzWol3faqcMfWhl8Ad4Wfl
9L1HI7KfkGo24v7rBlzAEDV0+gHKSixxeWdzM3/ZP3bbOlEtvZW1pEvWeojcpCOK0n4P1E4pQext
mY9qZBDNKXCAo6xMUCstejWGZU/Joq+waUZLsI4pU25q7N5dg3FZiYfJT0Cxi3QGmXTeF+MDrnRU
INcHczDMMLFokN6aAMBZpRdWnbFwJfQK7Ajk4idzvuz6g/5V8Ru2mG/CRK/5RSJdXmYRRyWfjXB9
aU9xsJQEouu3R5yIz5YOuMgQxUL/IbN0VxMxrWGgLH7DuJJi6woBqvXqqxX4BzFihGKBhJyDpscW
J8z1WjKv+4icHOoAKMrlp3u/8LzJHwbDABrUYoiALaXkZkEHbJKCyiP/k4dSSf7KfV5zhN1GFW4t
+vRO22IPujYQ4FnBtgLahlqYwL0+9RAoMR61dwC8igz78t/YA4AEGrsmV4/LnblXuUFF7DNeUmjs
LHdMffaYJ0TbAGDOG8yS4/O8rKkLZ6qNVYQTqT9SGlvI5E019CnyLBtxFPR9A9njOopq0aLeiH0W
OJX33haa8Q9B2vrPMzWzfShXVy0itp7sFp8mWuWqCyzHzZpPj4n2Vc9EpvCTbpHk09/iMKuS/gi2
Y+28njKGpCH537eU9TcKW0zsoyoJ1gzFPVu+TssStoXUnCVqPnIm5AQvABE4NFZn+MzdX0+WKy5O
hNt37SKFCrzfww2G/57bRohri3A5RIRYpSlCCUCL9N3+wfFYtj9Y9SZ5OT8xpUlLCQ59C7+EpBLF
yBZGV4DVsvPIt5C2wRNAr+IZcm8dtSIaVLNxweXO9WjYfpA3VlEU/RkmOa2cf0rh61bJ0MHeibh2
4uxEkvYY69CYmyyuRPK9SC3A3PK0WyFnv1NIDhjpkbbTtE1NqPNvZT+luxPwtZoRa9LpPKa0nOKk
fNaZqP29V2k9s9DAhYSqrqcVIJGpFBhOJSvA9p0ELWMBs9jQGo1AiP8UUs8wKs9yOAIVAughbBDx
0gwN6MOED/wUrAf90pRJ6TUILAs/QSjb6x6Gd6fc4FG8swdQ/pJ9Zdz96DzZBNK0cQ7FUFER1qjG
Q+xAT3q5yjrOqBD0LzZ7nivOLZVnqgHaJ9Zq5HsB3ZMdhwZjLNBtPH+0px/egQIX6izMuobHTb6z
5aCkMYL9nzrCKLfoE7fERXBs2zfwlDa2W1THd6N8BXWqkQ5b12E81o1sbldP3mYiBDmgqMntWKXA
d3PjoheZnr8UhbajL8zQz3k58O1gT6V6l59zzj6QLaMcO4Gru6swx9cRb5ZYvph/QOGedsBPzzju
x1Sn5zVR4R0i/XzPgMCCJm105UjIR/TAZNnPQ4fyJ2eQ8161g+7f2xHjWVNdnZkUtQMC9m59Q+R/
Id5R41MjRy9DgoAJOUmlpvcM706uvdwlEgCgHg6JXMWG3HkQNcvcUBR3AreUHQU5Bbwg9JYPukz5
JJAW338YyRAv2ftcMs6Ebw507+xIhfu4OjGJKynZT/SYBIBZfUalBSBld6EvS0npSImmUpKe8vzU
ubpXo+3CF3Hon2SUcMpvmtAHLl1uTytYmpV/svlVTaigXxYLqgm7uBJMzmWzMsdC5CZXqsC1x1ir
+lX0ErgT0Dua4IyN+cEYu3N7p/5eYVp/yedTcL2sUBu+z4ZrC1AjENHqGnWCPTMkgVhf8+cwRO6u
bFEJl03ML4E6oHLb7BPT1GcLFYYRdN225i5sLugfYSAI9e//38/ieDsS+bMTUKn0Me84xKsWkfsJ
nr/M5tj+Cv9bY4VwN1FRij0XJH2KX4RfF2c3GIgWt8EJIzkcaHcQAIbp09099cP7cFOdvO6GPZEd
WzbxMxG03yNIhmJM+VZHl75m3+BjFKgtI7d8JNiGCgefPwXPapipVjqe83t6411gJxPKxIVZ2cKY
i+v7AYmQHkiApQzYXuYVNWUkfk0I2C4kYaIk13fujzPVv0uU9nd8XPjDiil0wyIEgfBysjvjU4pT
ZydBlNxZ8deRfOoTU5XZvuZUYw5x/RKCAGb3ECjOfg+FtZBVpUEl5jYlqpJXO0DkXIXLsp37KgB5
NfZ/2dS3OfB2OlFsKNJpgp17d/3dwXZitjNCkZ/XDWeGyuTCRkIDt3tK56cdmzoakgQo5VIVY2Z4
YhnzURlxYuLjALiHSNd0rfRTvTYr7QGmR1DHGTY/nUEcMv/zMWD6qfwsbxZ1a4P2ajwRi/w6yIdF
i0hf0kFNQN9cQOksDTmzQSuPUiGaVZPePXdSXymRTqQLpNmfsVRTPmjV10VfVGOjBIJnU74M9/Ox
chxDUhQXh3xu5nfvTP4PgYxBixX2OyybwUkAASJcdpbP0y1soMy3Vve3lmV8VrsGfkx0o13jax47
lcgIeMMA9oxvfYm5ai9sGc6UbwlnWmfcCgXS5Wa5vkBq8AGpBvxyFlnRNfwU9re9Iqi49Pv2zlOJ
PEjGriuOpf+wVIwz8GTnnxxAcqGNKRy/AaA+Jf2Jj3JbbBJ0YP5dz1ORSiJmuB7X1oP6Bm3HKYgj
qtDw2Ojjb8DW8BTKAwxX/ZaPmEdQMBFuQjMfo4IfLDQXi4WLY1B7VaeVGGEj30WlmkXWyHMEUHAO
OMh7cWofiZRjX9gn2mKACOSkl5kr3+U4t582AOvVGx/4iRG83fIpCBkAsJfKPV5afY1zFTuFLDNC
WSgs/zBc5Z/JlErE7gk3IjTMx2c4ZqlJPMNON8Mbeg0KGAa/AZ6RAHJg/8OyM4imrOUrWZPL2TzJ
+cT12HwDNi3Qi7y3RttzmldhuKX1VZusG+dcCsr/8TSzdBC0lG7QIGqTn8TiUVzqXV1UU5iy76NF
UHacR0FrWucrT4PqMU4M+isdNqke5glXFcy7oDGhLRAlbxiOhz+Sk8kaIwdj9XkjgYV7Kw8LpTuD
CMhaf4kS52BSUkGJ0jhSg5kjEkR8Ya4rR2KSL2lEYK2LGXuKgds2Qjs3j3NzkMio5VgXOHb6l3RG
o3rBp2BEhPu+AylpSYYKvtIWeU2M9tPGz0SHN8Y51NK+S9YNxaLWoCtRVrl/w+rWefgJUu9u8AGq
5zuVuqd9FDykTfO9LmitlpiM95tguF1VeA0kP0RzzOllRL04h3VQ0yG/SYAl1k2MeWqjiaXDNV4y
cSKjJ1/cOKY0MKbVawomOY0gaZ/l8uvDrOGctWwwltcfxINfMo851VbO0nYTS1w3iTvhByh+j8RF
U1J6bzzhETPB3c4HAdjH+0fN+Gs8CwJfWx2O79ARkKXgvP4n3PpQnfvkM1QGVHqz1KtRLxvdoVWY
8cj4CSZdsIDA70eqouLdbhAr7/MHrIXjY+fUWF1HuyDW4Hp0MFaUBRRlfElyOAhja/eQ9uNn6HMo
t+9M44kuy+FO2hyVORP8zI3Jpq8lwFU5/0SkdxOb7ZXAeM99bngV0oVOOVBfxDbHnmojmgYHrGE6
yt4gP4wzr3llQo3tOB/FYKa/CUfW0uRsH+oZaZzo0F3ErfCypdYSTLtSVObMvwaki0dxsTa0FJ4F
xdCOylTGDH5R9CMXDi6607QDets7SaN3LYIC6pWPlpvbZ1LJmsJEqi7rfqIsJ91EWDPmpLvKIccC
r52F1VfisDNVJx7YYQBwMJoygbDlQoZ0L4gCYZS0sBJjXK0A7wC+VTakJDjma7M7z3xNkVl75EB3
NdoZSyjBxqUNiAmxyvvyOMNAs9xNxX4MmTpcG1y60Xt3Sj3CY3sjmCw+ZoS6u6CNSvIuQvf4tuQI
nIVqI/Q/EDShMWYW7KWg21pgZV9zwRb5WSmu6ddi2XjznVH4EwCpJ24nIfSPXlmmEx63MxMi002v
PgU2+MEOQNNCZ/C1ZuXiA9BowTHfGM+1X/m5RdD1KvMh1Tn93Ossny8Mhib6q6Hcet2L+caxLi2Z
M7CB85To8OPeTvRJMMeOZF8HBBW3z7eNCfXp6+rKMFgurGt+4zifVHOhRSQIsQb0YXxrflrraFwQ
ikNwKlJEcu0TWomi8gSVZ3OA4rIrmASYB/K6PsQVTGulUM14NXY147M4+M3Yj2mf/nEMsDKDZTHH
Fvcj5eePPPGEp5mVHlm3PS0o+yZW2WG9+3JsrPWRxX6+sKrg2eNLz1Ln78xXPqEIpUPvRDkxKcXN
BUFsKG1katXuLJD5Te22O5kL9TS3UW+ceqzrWiz9Ob3sVvJH5zYw73LV4XLc9Yxbm0Nsjbsh3kKB
7MOWIx57NBS6Ldo5EwnbksL7na5OGy9r98clWiz9bJOzIWanwCubOJfS3v3MIvgeSuEPZ73qWyLT
ZeYp8L4lV7+ZwPVh9bIK2A3mUykysuEhNh3KlZrAGWnqdp4VKjlEA65id5DiHymtcAXziBuAZvz2
+xJK0j61KthGm37A8Gc13FjKji3RI3XYj1N5478/fAYB64MtMob/Cma3Rk4yJ8iHoJjZGyCfGvOH
9VRuENo/pRG1lpCN81S2SmdqEOJQm+AC4nuG/tUlkStDBT/DVjNPk6Ek9vXGBpaIUq13iEih/6H8
HEHfG1X8GKd9WHHWEzj7LbIgTq7WYs1KtwZqOZznsmxkwCOUdLV1ANpsiUtpGFaVzvdMmL38nMB7
aMmoSG7QzOFSUw4yaL9hpFsR2ZE8mx3rG5mzRpNv+LdhIwrNiXEp2bF8Ycsj3rRtZNSWCAKfvL8w
mNbDSiLkroFqPzTt+ONkpShXCg9oZE8ynoG7GqoNXHxzo3Ct/UITSpNSSY+xNsV7Ws1iUpk0QOip
3TzI+enUlv0rcB7N0FtEszi9hjmG5vXrdVNfb6QiEyCaE+Wegq/wsA5PxwFM2wQqVlvXwSBp8btN
M0+n3s5nRvze3c37sJXq5V+oO8m/WkuH12uGf6sQ7BCinIKE+TS2ogtygyGgW8g3E+lpDzT9423T
tVPOXZ23yo7PbIrFrkTAVMuUkTiZHRNbQvfRz6M3N9YahOxzT5Xo331zIDMvG84bESSPpL7dYMAO
oLO431DPa8zrooqli4iT62Wm3W96I60mGlNWZMhpqvY5Yng2gTB4jkgYLeCVkdAqZvIaJrPeNZ0X
cqBjN6jZJApKfe88KIy8SlEsWg+dHIwiKbNv7AGr1Xrt2Nqa8LaLDz7oTrqLFBrN3jytFv1bNJ44
vqcaW9kz4a6JB4cYwRTgUkaErjZY9tOCAWaWKrh1fCweozesbxcrPGiX26Xb/3NdTwlR8had9vTP
oOuOUlOA08kxA2k10kFQLyC1CZDFlvM9Bu2M7lXkXtDFgCrWFAf+bZFxkuIsc8m4zQpaPF4utPhK
AP8kwlJ1PIawgXfvat2nJDmadIeFWwWFYIyipJ7+ZafpWGiRLXY74ReaqEB6yza2693k3b/zmFg3
pceXTKa9ORPeLD4U0uzkKqMeL8SNTpV8fztOKnEGvDr2W+xFz/pRKJzqYAtF5EOFhWK5ZnzLZD2F
uZ5WDLE+KabAN1czxp5B+SLmpX6vCJHiG6hYUHP6lXYrEUzxdY22QrXxiosVojaFwA2awV4NVaWr
1fvgyaoe8AuIoQU7qEQ/ODZ+abHI9VWlG16iBTLrB+E4BipYC8dn9U41IJlY6YiHaVHenn+ulq8L
tXDbg0cf//Jf/+uy3w7oVq/9lJ8+ttIZ/8DIyHgbdgYX2QvYgNlt0dbGjAN5O8G0qyioI7zl3Com
kYevGrfHMfJeYC5SNefUkXLURbLocVml7HgbOgghQb04fgREheH8HZFDK9+dGVsbLrp/ejbmo+ha
90YqBERANkp7DrT7zThfiWCCn8xCJkBXKJi3FrML4+YQJcVqCJXcql9WpQon5hKukfuGXKXsBxL/
+yAiiYhCuMUUQ8P1j1kQ7Br2hr4JA2WHVjddoK0rhTtBGzZ+Ib70OvRwRSjnZLR7b0f2AQOPRdtP
p7n2QJrAJ3+GKsSw89ShnyCz60yYMkoLgicgPGNFeiieLs5wCZHpWe/WfvVktgo+M6brub6hNNrw
+KwvOLqCO7fa9tiS2saKdVTCJK4kDl35ybyzbr7V4q3K8rvx9svbiKThPuughN/AkosYaS2nn+Ob
lHiUdniBl8E/FYIf2Gtv2f7LfjQLPW7CCNFLL0xM49DBzzprRggvQnxXeNIpdXzEoabuTU6bi1u9
NQv6c1C69HwTf645wb6sPWQd7XjG7f5sDlPPmo1osPuM6r53bY2tx3od4DBvSjMzGsKmW2qfcUxR
Lm0HTzNt8G+ept5SeP10zX1T00nEEHAUialIZuCRV8xnwqMCAQi0U8rsQqPQvLnNhgoKiat03bph
XWuvzC9Oo2UsyiwkPyE+1UeJEdYngib3tEFcq1vlx7D5yNBQ2TMyFBB1p+f1LDHDzsqqwlRhsxy5
PrnmSnZspdQaFvyBdYrqveIPUVHQtN2e1MvjK5n06UiCUt7WVmZ6qXGcGsv8QuEHnFlfMP9by3AF
ISRIsMVZK1BKv2inZJMCo0otX4jzhmnAcMOFqZ4btRY2KZJSznJmRFNt1bPMNwMavDlC1RV2AyVB
MKM2JAI3h9X9zGzx5CJOoiKf1VSr/or7vjvKqJbfh1+p/FZNkjy0D7cejhuflVa+hqV+lFydDGwG
3tvaXfQowvzj0vU6cBDSkLgNevLMYzcWGviKN2QpYddp40uhpEMh34CLSX4+MgfkyBwnm0vmPoUR
Vy02rWM2fPHsSRyXZ0oiWrOWjBPemV1wjq1Vi4d9UUYD2SWoJuRRFdeB7Uuj3u+Ygt7EbPpYX67u
q6I3H7kNpcphgXPTzBAqlz03DnltXafmpvwq8tP636qZUA/N9PF55F9R/hI5m54H3noWiOieW3Gr
DkRlRM6ensC4B0XdGV7326sCnmDB1jaTy6C8s3WzQZ3qB5qKk9auYYDuE3nAoKhrpmLcBjeu0ri0
JMe0jRL3OvUcoMV8qqeqBS/DlUagG9PXTP9RPGRhJi6NnyVXfTLGnVKfe8WPBzHRa1ZpX94mMRk0
RsooCpT+KnJXStQB1AoNd5KbdAXdUt7ci/mP8JByHe3bWDP8ZyCBol1Fpo3vR8F7mHRaiOLkyvQj
I/kqvB4HSe17gBjIiNR35eYKFHw1AVSwnT78MizjVQn2l+HS2MVanSJFcxkR7zAS0ZdygIxyw8Ty
NKbg/mdMkyFnAjWtitGZsAOgvigxidfHQh7ybSHOyt84Dd055Af6/WMInirdovphZV8LMo+3YWvH
mApvoU7NObfW/cw4l9E7ipvfp04WwcEnMcb3bCo8btPxE0LDb2CsMW9Zi/nYspWjK1xTsK7E3f6N
1dVhicKwN5oVKnqPw3ZoYSLrbkR22cuBZd+dDLdP6YkAsGDf/w9UyZOioJ3V17xtB8D7QMVTkpll
oyWqRAcWAaNaJYdwzlY3oTeYgwqr6p0PBtu3wT9cUpVyCWQLlju/GHB3c8sO3JIXma54P5ndijjq
MmNs5++T1kSH/76XuE/dDhbfxi9LOJnTZitOMTTCVr6zVmHdT9ZZIuz0ObHgGGX6spPF/Jyu6lRe
V4qQsG6uKS0Dq9KuoqeB5hVy1JZ5uvRO64MPkB/qOmnviJfaHaS5gNyiEWFFOSFjTTYF641G1SdM
RkkeIisM3Ox+WPvQ0r6P68KNty61+KJBX86NCu2RJUMtflwQxWhRkx0Oj+X46UyJ0mSBPb/OA0+V
V56cRtfrrXFSQ+vYicKc5JGs1R+Nsho+ZrLd8L1w3KM5XXOhyM04rDRbkv19gNVKrf5HQU7T3TLF
PpHy6Ej9tFqrJ75/aR+QHyS6hBEB8AIJ1qIS1pzpNfs2Sf5ZYZH7HgKPTOZBgvDy5PoEOOx8fQ9V
2wE3dOKpB5e4P/IPiV3gcq8d+0KXuhUrtbGPstYzm/DE+OQ5o3YzwPqIL8AA2F0hKynMEg18+Puz
XEZ8X1sw71csEs/uWCe1k/rWMCNXG3EDgTIWTTeN4fm59vwdUsLvJAET2Z0O2tKbRU4Ux+K9bUgo
i+zTr3ilpMct/hvTpYVf/DQE12/QvFrpLDuyXrbFG2nECjSSKMlBQU1tz2Lu6RTjtSe96cDPcDgj
K7VUHy4gvqkxHk327d8CHocXEMM+EcCdafmac00rxkROLCDA7PGXr+PYGISHZ3O6bRFlPtwhkoxz
hbQD/jLDpkKshQoIwyit4HOkOlTPMAgC5NjZLYe7i1PjWTvjYRzVhrogzxwlZnGiuKsi03e2rPN4
c99PBgZPkImY1xqt9ClBJuRvHba/vM29UFNyYBXVEKcPbgvNWZ9iMBSU7UjttkL57G0kooFKRfMq
TvDQqBCqXjHAY9UxkS4fgwahUcddl/zYn1myR+rTFg931oZ6lJ8xJ4ss2lV5t4foTIZTO/iL1QAH
p8lrsHHD8yaCdy5ju2MDs4dsoGHmWiGFfdT+Q8FbnQ0gZ/aUh2QmmEf6OT+F0+zC12I+MXZWilKU
3vmSmkSiZooL9bpMnED5lXWdq1tJGg+Q5UQ1iGrAbNxO9BF6K4jiRbNsBZ2Neg7JgHkVh5RoWJPZ
vlH2qWLZw99qd1lavPHEklCS1MIzRMS3V6Cidf3dCjf3jCq3l5ilU6/0g+6Ou5nQRMoqQ1aRha5v
kQser1wpOj86EjGmLPJwCb4miz4IMsBdtASklcNioUBjTBiP//FFDpMabpXwjd/GpIKbzyrajAZh
9lgX2DXtwDDya9JsNWffXSBM2IAPvL0a+qoz/+sQ0sNBGO2HB4VkieA2TNckTDO5rAZslmE8q8X7
GvD7OfRVzTF70c7MhT6OgfBC5cPaqOBJuj9r9n8/OLKHZJqktse6xaaJT15uAbNajGtMxFn71mf3
k692Z/DoCr/kJggoZrJAAz8ffZaZ6aae6wO/jiB8LDdygztTTedfCyWPaIYHqfoLjWrWzJBIpQSd
XR3GLW5GWS9YgHrkdz88S3JcQqGM6Q/1MdbhmXAzkL82FjxMol/Cyt71EYjpsxn7B42fu5Wlbtc+
2hmV1GmbzoHew/JBZ+psoN8Ud1/nVC0EqjLg0fl+gEwuOE8Li1RLRVbaXFxsBw0kz8CwBGJB457O
SEOwIBIcGG1jCLLEFfYu9KCSDCEeMLj2vpUS/Wv4yeMo1Wu3BqC9J2dRH0R3GBhiV87Jsvzw3rOO
h5V+K5/ioo/o4U67tZ043LkBB0UXyvXJ3n01nzVBh+ZdYrOVNu1vLLCqv0cshNcyjCxyL2lQOj6r
ECVjODcgw5Shu3s8T1IEkkaMmTwKjDH+nLsUAAK7Edm5++ODRLa0e6GrHpGHxCsAx5oCVdCLnthO
Llt/RY6K/Z/dqlTqB2FlKf3jrJIiGeRSy6XN02WlATjrFwuW3eruR5bsJo6bf8mDjUvkg7r5UXp0
PieliL1AOdk2WylSo1VdQlzHiykA6m4LXghJILvC+bhiv4Yf+jTP2/iltYlKKP9in+07tg0L9zr6
PxTdm4g3tc3WIdcJ8Ns/x4PnztGN7DUS6DMHvNy34U9vFrkifcxUoN8aQqTw1WGZg0DFJBMBUW3D
c9/DTcC33JIf5e6itS1ptWgPKI4Be5pUNSJgawyb1GkyZfZepy1Hf8nUFO3+yFM5PEb2NnjRKaKQ
a/8zN/ATvs/gHr+bqSPgqfAy9UOWhwg4kIcP8iuE6yfjz82po2ih0fwpR7XldAjPQMIMDjoj22qq
NxkhJj/8WX/mdA35m1MHoEvv6EUYAitfBnzlYEsA4xXKT+HXUXO59nqe1PYxFqUH6F9Gv6fo8jNl
R/P36On1dMesUDBhII8cyQtCFIBGWQKhEIO9YU6LTx2w34Gbbxr9M3xzUHH4sB0G4UYMa9IwvMOA
fQkSCs+f2DZ5X9/cQF2TOOZtQ9dNdvwj5UdeGa3+cuPlvnbBx7fh/CM9iCHWpmI979kNztQNl2YP
7fqAdPLL7ytmDOW4HPUPk2YuYNQpjvhgiBb4LgvUXlMPtB18wO3xCq09WqR99uM4pF0MSvwCDZgO
p7vrcMa5mriOQXJHUldmUrSPBYd4l2vVl7/DESJGmGczpPXKCySc7B4jrhUdiYMMJtVXZarnxSwt
X4AUDr5hbFzMP18GyUdcKsT8eVJJvKE2VjHklrirLq7yUPBngih9Hc9i1MMge3KVYfqdiPVzA4aq
3aN/8PDDrwaXqcAT/xMGBtpdK38V9bJLdKSmuwxAg+JD0UkVUDslZqpffWFG6QdrL4qq4OEWnonS
KgYopcNXgntDXutma3pftUkoKWC4ivlEL5opa32VhdnZebMVNkHXldvsxar9iTBBZN5Jp2HZt+Uv
diI9HGy+Q+UXPQnaJsmECZziaMTUhgYUSt+/ZkB5bmpoq9Ztx7XxIACh1UygfCo3IYj4L68NOYfB
9H84dTD1WQD4Aa8ZqBU2JIeV4TfTFx8eKQspwvgIEgSeGlkHwTfgf1284Yj3UNOvRwpSsq/xkf3M
QqjHQcikILaokh/Z4EP96jVKS8knxfwJwLKesylTHLUm9I9X8AhS6vVyBFh7wMRWJqGsjHQblrf3
6YVsmr60EgkuJH8zqRns4q+CyB+TS5YP9Li4Kjw+4T3Jup/MHxYxtRxDKJs/ObWV5ugD4TrDWLLV
gNsWmPH443cfQasMGWyVtxjNpV1Su8jjdzJqfj1aHt3w7iLh9mZi6JVDh9rIGOzsc5cIhByTlDzr
12p2KcjiMszi91B/cowCyWqWdMZSaeTEkO4NXOU+/kph/3AqDMB2UfljurEyxNOXpYfZHeBPx63p
GvSr17jJXmSCITvnm92WRZFFmqxZE37898x2a6zpijRMmC8ndWdIZnETE0o1Ua4+aDCklrvhpkPl
wm5cB63Mhd158XOsY7Xz3Gt6YcmJUxZRFErGq/PpH/d9zAgjPb3U992kcKWF2YG7zfbxaCV+pei9
UC2J91oGuNpouG0n+QFvNmUU6RwsMYLrmGGnaG52aoTgBDJixA8OkfuLSnUDuv7xb3JDK7PQFb/3
+yKBxM+/Szop0RTkpVA2utFeH/Jm19nxmt93I6WTrOzHAt4TtWdrTtXybdm0OLdDrQJlm1KBiNYB
kHF+TRSSk1NeaIodiLrul/pfegg1QG6JEE9cxGky0laSRl+KNsfDmdd36VZ4I2QzEE8t6zbBgCVG
/pPztckr3lSO3o4eoEcjuQudOysi4ePazSITXb4M9SEZYDvbZS3tUe8jNTcIjcYbSUY8XG6acBm/
9HE5F7AsFaMZ9MoT6PLUwU5g+8ZZCnvTst55jYW1KvTunQ2xh0QOHPgyyvAylwPVV1hq/czBxKB5
eMdhBD+E+5n3Q+igOnTKmpqMwSjR6RSRvPnC5m7b6xKfpwI92zDrw0jtL57DLX/OJMc/AnnEbYRM
SQq4Ca6F1ZPm1GpkgTxQFVFHVaHvzp2Int0Lo+TzSPAZbWPYeW8pTVa/Pn8+ftnWybrpT8EJK+86
9gcFvgcJV2Voc/ZNFHAxjYab3Q930bWrOUPdJob5SuxldWV08xn/MdvglblXnjNRi0ZgOROOnxJa
uBH0f1a7DlW+0sR4W20qx4k92Lo3JCq6BDoCCjkqMCquUT2O4mBGQd1udsjP8P+t+rcukogTrGt+
Sy6qBxcYzu02D+hfVQt95NvRw7lhVzeD5UYbLBOFG4YRIbDSjk4Ds0OuOYk0ns4mOQfLmWLTgQ8z
GOjYdeNToC0EZPDgjZL9vI+HJqSAMSM6asb1XjbPUtCAnzzyPdpoDr0iRip6O/p5M5EcCCH6yHhK
Ll0Q/ldS/pkamqFQ6kzulXz230CjmZxss9j9R4YZ+Urug2Gs8dZGkdyZ3P+usfslLsIXIyjiC4FU
9wzcNiYj9uy8ONcuCfoW5dq1x8SHEy5kdZqulj73bXXBNkKdfVaPNImYurhfKwxLJXB7J02iSMpe
iRJ4iuw5AteJe+BGQJttXxc19MihfQU7L/vqGTN6grz4+xLcMcQ8PE8YcmJrp+UV5qLfLzTlPm0Q
l+bSUFXFu4+cxp0kg7+0g4Os8AyvzKQQtm8noGcLIWfNFLZ6FFlfjQ4dJ9wPGikl4EUT3isqkcMw
OtBMdxz2DDmjJgLzPrbZPoigzcJvvvuQqGNS/xvXfL922LBzlQFed6EHpIYlKEoZnVLaB3j88+t0
chnbSm/ToLOMmKYArGNKuZrXadXgVOtDGgoMAldVl+3poIjogzSfFnRe1HbG1rCJZ368zyjDwQtC
ezjKHzhwNfkASbhvxGy9izDuDJHvesTRZym/MoTagV2qFDbVgfIyQDkX8exXb/CEIlhICnrBHGkh
KX9uNNEOJNooBPCwZRO7z+EdnyVjRtv/rvy96omLXg0ctRUi0WxErP+REkMNx+5/Rr4r9wqdHf4A
Q1hDf6ZD2oeZAoC8QlFkn8NYY18QmsQcE5wnYxCuthMD7r3Wzcvu38rTHBGTVSkLNCXcL16fDUiN
lWy+foyFKodEs33D/M8b6sRVbcfFMHP6H3UDmCEA/2I61zcbxa7Vd5ihwwBIBNULHOcXI5Ygb5xl
1zL62O7sFoGB/xJUz3ZjP5q1JQjPDD7yKju8+ENEXj9JmZQAVQI9TtSrMuwWvfY0DqHHcne3hqzb
ZR8pbwnaWgAth0JT8kFlFKF5frgEmDGhtJtWiuwLj2ZZOdLz1Be48kMAzS4ZCbBt5A3M9Ksteck6
Y6+1apJXQ8J9kCDmjOsRhAKbmfsOAQe8Dbt19GGrvRY6tVScmckBmqGlAlUqYET6QUDkfeDVz5sN
v3lIOHG/EHkagHeFtqJhaJT+7IgKZOUagfoMM2OINAunIz6wHwkGGAPxyWg8q43nQyTUvxnK2fhH
+KdjJRDzSt4GCNoZpHsZmt4fgXMJKf9W++bV9VtDREt1hlqj/tFYa+CPZk39+YWdL9e/GN0h506+
9HiEBV3Axv1KJShtazdqX7KPNm9/KRUsPSBq+5/QZ2lrB2wy0o45g2elEMfgW+ezM7z70R9LBEBo
T2AU9tOy9WbltIdCcaSkxUaXnrNzcvUMe/GF69dfiZg7zgW0QnfR4LUiTQdJu4G1AknapCsBh83/
jHBM7jq6ZfP/M8xHltUKtOSS3QPG5+fD1zVF1/2SZfa+cwe3kYPnjRw38b7WixdB8BWvLWj/9EGw
WT/i79iiluAAdNIc1IFYHQbcu+asgRqWem6bkQPVgGARakzweSf8v6H+JINY3YIsRRuJP8DvbMpx
vVlDM6Jqw/lzHg5E2groxQSwCh4mVuBN6C7iKHN5l1z9zi2M0eu1gpc3auzm66qb3NCxOqS/0KKT
Wth5meiGFqtEiJCm/m/S4RYE8OcmXrXA41pRKRcSJqP0rV+ZRiNJla90SGjEsq1NapCJG4y7mUA7
PKblI7oIYoHzsOZwJnvppdURdgPZL4QjkWO/J1ralUK3j+tNLlVJCHLaYW58xkbQgmKNRtF30nYw
RYZGXw/CrztHgtlVjK1CnnjT7Z3n3MtxFBmxzW8q2GD4Xr0udYlf9X7gJ+ZgXPWjj5B7xjYU8tT5
ea7UdnANOgUIPSG9J1IBuVnK5c1t50Ikx+oNkKbyy3WAzZng+qzRb2p1akVzwg6mNgcZAnsYRBy3
evZY5hS88W0nexn24JdIH41bJukRWtpx7MjT+JY29YPhk87vGJvJcTMc/4oneAFkC5G26pvNvfRw
WePMGsXf83t9WHLW44jXnwsUHQH1e/Um/1DCkoJDN9qoBVqxqjoy//zDv3miK7G5S5jG1dzCnbX2
DPNqkiEg3YsHUYpF4U27IUKOnIlZ6n6+0uC8mTEE5o/ifBqC1W2Gk3oKr2PwXm/kclNa9NyRvTpV
6agZ1NSezEQ1wF3fqCs+RB34m6R0p3byjExW+LqOqXeTGAi/70q8nn+Beh1asMhNy04UiTwT15C9
zoQ52HBcWVBiEM913uqR4nEvBsFLf9KgsdaeSpw+G3GEuOVWN9hF5oyKwX9gjKNt3QEBA9O6pS2W
LGGH/QAOpt4ITTVI8OiDiSrE6F+q0/2IT33k1snDu4rkP0Fko0ZOR9WoteOtSIKguRvWayTBc5UF
Q5lGmKqdaDtsGt8+cBavEe7LfrBIB5Jw4quvVMBL8BuogBTtUUupHvF95p57TUdGzQbqTqGDh6V0
ZgmDJqUHaJ4PDO86T6xWJ0CVCW3MyEA6HLI/oLMN7mNi8E8kqtMdjrPX/3qUHFnpflZDtv0u7cu6
K7XS6kX8n4JyJworO9aprCLkX6CZM5DYoeDOw4N1nf1gMWpI++FISkCjmQmnURGwxAtpebxlAP3G
aEObDJbnfiINqneRx/cc+lPbwWQMW+r9XcWcV1BrlvwpksJR1TvCxHKI4EqUAO1ZAilP+vce5RLu
JEiRQZdoqL1Ya1yauIDeVWJlhJqoX4JDJjZU9IPDxbqv58odUUf+HXQM5nxh0M+iEm8uC4WHaFeG
9D4bZP32BQmWzpB2IeG6Am29UJoQiP54tUcWqd3H65ccA+7B+L2MHHWTychcZknfHrJQbXAUwDRa
XUqnIZDkQKKwUhVuGRF6vayhAMDb8fyyLu5e0rPFU2X3ayNOraYgLKVA9uhcVRZRwmQdO6xUus/I
jxbK2Cc84wswPl9V4W3NQFHNg2Bud8tew1td1ZPLBW1GtHrF2JRXyd1yYyfHlVBqLhgs/KSPaQVU
BMzOq1stFCJqCAPh3CAwYlxZg4i+gbpTaBcG5RoyOk7K3vcjw9PwaXguh1tfWiyq3fH+3SnBdCDn
yXzxLqPMn7Ek5fzAs1F1AlPZqMEBB3POK3OYvIm5eMfiLFZif4zoENmqjxNzeB4esVoz4kyhf7Ik
utZj5JsHuawdXiaKYe0xe+WYcCsVc5ATXUEnv/83TFPYnuxB9mUce88MxPoQHJwhQ11ocTdo7q9/
GHUpPLIZa0kU0xQO1km4Z/qt/WLyttjk5CmuEIHfW8gTqOteNkzmrYjbIQhxvykAr39JcnShczZN
fLEQg7E9UkDZ88Jay6fVu4aIJWoqCc1Cnm4H5USwUd1t1VatYpVWyMuVGwr0IdawCvBdH2mvd5eG
i+WxrYa8Vya+zj8KwEJb7LmutVxM/Rwepl12SWMr0IeJR6FlbinmPtI1fM7CtnnOitJbjF+xi6uU
e7Q1TXzKyMpaT9jx+UlvGBevVwuFZRDTNcKbeBEwODITAXBs/DJEb3v0Qg1PLePLvDilGxP2TNjs
p9THS+rzswcn1yYVJC+FkHjzPjkhn6WWJhB7bl7O1ZkM5nZdAJbL09GUZxwA0S7I+Ca94Xe7ToUY
NYAOg1cZJ4gn5VtI61pkSAri5NaAGPrxrYhQafymGk5Ycq/tRSsCsnZ4SmrG8pDAVktnK5Fc9Nx8
Xqvm/V+6AhabgYdXpv/GcIiJwqr9dGhu+bPyvpT9UWjQRhInB4ascn4JwLxrYkCJ1uHiKzWWEwpR
nLZZ5AAHM6dXg+aLwFDLTlEassN++xzYmr5STIrN+EPoCt9ykuAdi0GwSpLRzqC+wNx4QHrPLe+m
bcppfSYRbSKsRgpkgOiRZWkAZ9mpvR8s+h2jzWFiIh3zDM0pPYKE379R0D2Uv8BLXpP5XlbSXILV
M0kGgKBN0EMXqosOm1yWFbIhiTBAdLkSVtfisfFrZm9gbDzgjmV2E79gmHAlRirbfmkqQaxcAqcW
o4qmDq5EsB3Kk+34M7gDoaHD7rEVEDorCeFl+jalTLMfBGMiJ4EusYGo6MVu6HUAg+f07Usm6eDd
Bm1gUep2i7tW9ujqqk1G3k+AXn6HjQ9UGnhNFET4UWXENxcnNZhzSQap2rN79hxW0UPjPb+6p48B
eKHpuRNBBIzbyFc66Zu45EnKkjCLCrjcjd/SeM+3dgABFLGPdFU5JQhHAeiFI6aIv6Wn9jaQpABQ
ZNU2iKETkRG6Hy3nTr+DXtfcJy93PXU0a9wOY1Gh0Nd+EqkGAxsTsDdOWy/kPkcCqOp6VQ2z+zmp
BDG0qCAaynyNQGGl4jr6AR05MMVc+0d5pVvc+Z9b33hkJKZQfYZdMSkVsP8f63VVgypvqMHAJmI3
1SKWi3xU+90TYPYPAr3Hsig7b/QYgICxfcs40L13SK4PULwPVdzap2/YvdCA3+lCN/cai4ObeUGo
bBuMJm/JlMZcdol2leeNvhqgRbltUppyeqZnGTeeVZsLou0jQKr0649AiUX/WMv/zG6Bu9ynP1A7
r0pkE0IkbxacTdrhl08KLQHE2To1Wh62cfgLCECv4p92VmZU3aszdrmydyjE9+hb6fWL0FdymhrG
egY3s3nLYj0nn1JfFQzkNSiaRrTyEXFd68qZdU4p9xGsqxQNRJTcHQ7vJqIsYC/Sk5fHkCi6Hoz8
5Im59pK/vfZhSa0ZE1ZQ2MYzSmA7VbLOH5jMs40KFE7QOk4brwkoJvFwVpph/BAIMttcCqqrIkXl
kGHKe2VnxP8RmzuTunoiUbvUiFhDYJ6nFcWEIt63GI7mEPIcMwN5w17pBGz/CoxNGIuLAtrsfMqN
ymvZ/szsquRuhDxZpuw+R4ba2/cIZ//BtmRnoILotcQ9buAFLbuQHGPYaJQQSScy4kovwrUWkBEG
E2hC2RDdobFAGzJyDf2NjDNrL8+J34EWzS7hPg3o6LkUF0fcpcPfYFL8qyCjEDruSpyKwaDIdNV6
9zXZ8mf9LKlsX1vWTkk8//WezPde4CisY6xQJhI93sfm9bbpnxNAtP51zIFuasdK3XBI8uq31jj5
70++XVTqHz1fS5I4lKgnbNPH6Ak4SWr5DhyHdHkR3Lq2jcBpZe4OiNJkotPhe50XkO6zisdwhQy3
x7Zr0GcRaytGHasGG9F7qXkNc2093RvATO5SbFlhI/wt9oMPvlEtvdxyQgK7HNas6Cd2ZiCsrShI
DekhKf26iZ4pv+6Veoo1PgIShlViKl65aJvq+R0ZMM290ws8fNSgSzsUCBH6MIDnv6A+wEmGBQN9
muXR3p9bdtmzgwtzKhFQ7HexVd/RBbizI9ELpE2GMhFG/EZziD7c8lviYco+zuv1q1edUHpi/m3E
i72oNjvZ12cI5h/IcOM6ij9nwlUrVQcKIVnU4EpGmiYNpVSwFkvKrEV693fnYzgI1vgpeH6LZJPv
pNjgbMNP+9ghwKd2deNArjDyWNxAAysfInho9YNL6bpWxxFYb9N5Bk3wClLCP8M33Xqvfl281OPN
IHH6VPcKzSNekdA8963QN3e9bPRq2gko37BqvCVhVd1D9iuqRMUDngLf08ygXFpjnP9mNVxzLoQg
e+y38J0zbvaWjGZQh7RPfjRw+GI7nuefV96SvW9w5TpeMWN1+wCAJ5eDBPEzhm4ZHBkWGO6l4Wj2
sV5ewhaF1PPAL200DfTSdptLibCGD+SBrje49eHKeVCOR6jc6adR5rXd27/DHkCRPOuzNiT7XnUQ
gWDOAN04spB5oRLROz4JpQaaTDoVSwg8LBmSA7X/Mf/SOHnrKtQeuF4FPxJEsFzxVPajguaQhwmx
Nkv6l0QNCk61MrZ6gFhJ1Lfl6vOoaPRByvsPhZPfR2wI4+X3NJk0PCpa36MU3Ll38xwft2DnSGf/
DZslCX28Z4EB+AyZifGJ3pZLSbl5TM0pi/W8md5TSQyoLdMHv823+lhJZ+uzccMJ8giL8DES9YQX
wNsHrZ0tgWRxyaY6k4mpOAepe9iSg9D33PZ1seFKHLIKd5yRK4IukgKqGiRRrWZPoe+tIf0OI3Gy
kZnX5v9nTVNVcaPYe9zNPxAUgr23WU1UfDgNGtte1b9COt8/KhOHqNk5EdLD2TyuPpbtyuekbN30
8i0J/C06xjMSttEhSqwy/EQQrRxN0EbNZx8M+iOuYpHtuape+PwgEQYKtyL3LCFcnn9maCjaepbc
M+ejpiNHmJZKw8WrQ1zfp9Lum11i7gAGAtMekcvXDD0BXHP1a+ZiYm5XdQU5GeDf7b9qvZ/iV6Qa
m43yVIzTFMuorWnf2emy0qsgM+cBjwd9u8B6rBYQNvN8CWStBOOsbAnxBjhExa1Fp5DVxrcNGJ6x
9a6GBRHAvH9thLYndSJrcgC3wEGESJm1HBolxDrL6tUgHICj+tKUGiC02RfCkWdO/jMEyvq5y+T3
AWKkXxvxQim1mOLa92gZe4UCMemywvTpVzurLJ+/zCrV8HpfQ1EkaUrXJAY0uksuhTaOH7o3YbeI
0SXTLBB2LT4bvDxcycPcSEUq9vqUAjZzZIX3dvJqiogDwcZ9pS0tFuKZSdNYQbD2P+5wafHBE3IN
fE6wi2ZEa3sqfDmRIL0x+SPHbdj2ZVKIBnalcsf5B7tLgDqPXZ66s0lM11CaIBntcA0Qg7L76PBC
AQkATdRpLM7NiZ2IFQeml0RWGonxCeUkOr/uPxfUGQQXIs8wD8C2cmY1kkEYX9sR+486RQ+q5xSE
dENjh3hDAXlJyIs597QOjFifPGdEBBYPw+GX/fIQZu5CZW6U8vWqhTaC75+yIw2RismcVgaLtHUd
4wnogEbRLf7TMHuDzVJT5W4NZRfHlOIbaU6KPaG1v6FTDNWq93A2JTFWiuw5LAbe4r4yOXT5pQ0T
l/t0fm334unu5tlaUPWxLxRt3y5STn6bXpaMJJ0B9U0EZb/jv2OHU+agiBkHoRVJ2v/RS619ECpp
OSxMWVJQ/p8eWknQHO6XbK2/k2T05ANmLKyb9AfdrqoA46Mor4zyuEKZdD1bVQTBwL3vG15OVeqT
kYIdfkgP/h3beRf10HClupQuG50jFuCmqQyVQKfJdtRUHke7zpy/5TjYJ6CKPW9tyF1jPvOFK7kT
KhxbN2yOSl6xmNJK7PZX7QoxR9iv5cdc8EOqSf95UmBZHo4afcTPyW1LgXhX0Sl2bKJsp8oQm9Vl
Y5lY/KsEX/bCD6p4D54Lg/M18gbhgNXlDjODbe/NIPbhWaDNhxxcf/LqYMygVPvNaU7a1FQgpKYM
IeXfESDTSLefPGYHsSwA4sHGYPfQ/fkTD7XKZSRcrhuJaF0tM5QVnuyuOyUCkMSP6VdKIjoodbxj
mtTpSSi7phjt6mMuv38nvcxaFgwDzHDxuM1bauEiLayE6KlmEprrLlCNEtFHDeqe7L3fFZXGqxXA
3id0V3n+pPzQ/Mbb3BIqrkHCvJQHW9CisvgksjUNWggr5yO+jhER/6FPzSIr1x12f6V6a97a9FNu
z7SX4vdaC+yOpLXFsw2e/XfM3IPJPFd6BfoRaAisUTUeqogo1BtYPc3cZvAg8/wTONJDqYhz8Vir
dg+2lM+TIGLfxQQAzMxz/RgB16lCW2M9SIS24z2SQxl1EwLvE7g/qjKg8/OGl1mVAYHZnyHvyDBo
Mqh81reG08I+ozdL+G8jVoFhBCkOZ2g9Yc3nquYIjaXTHUzoR6rQ6gwNabOX2cHYxeplFgSygxt0
J1T2O71hdzNl2SFGe//AklPlEkAvJjp4cD9KBEmS2u2GX05cwddTxiMWgqBm06vFdytr/I+F7cA0
iH63qbqC56CYz8ZtaKbUsLN2cAhMg9D+cjAjvA1j5umzOkn7E2Iryrh20VOhZWxAZNLrALADV3eB
2AXzY+0Z05sxEUbojyc5bufDoL42tOVOYs9lNxELB+Gl5RttKSW9OOjz2sf04vbGj3/mD/aEWBLD
JWnwuJSMbDNCfl0YKOj0fWwVVkXmrbxSNNS0c6zSwYDPW25zgTwJnAM0WOT+SQtHYDOXw/W8hydt
eM1v14uGJZp5B1j4tmstWNKrAkjP6hsNIH4N1gGckDJm4HPlwStyh1uHRxtdMJkWK4Jiqpv42n1Z
RLN//4kfJZYW7NjGxSjsiXn3OxbCFJwk5cA5UpJY/wFNGhKlH/LrtOr82r3ALeZi8xzKwhb92x74
RuxijRUV7dU+gC7l1CFgnOpjb5+Etds7fvrTp5ZYIuaPN3rrHaeedNdtyfMEmZsg/cmAsWpdrYy3
f4bRT59uFOnGbk31OdHXSa0mtJ/OzX6moDtpLzeUvHNhFwLIMLqLlihr8EJQ6rl7sYcwNdbMrlyi
NVkpcmQgpY+M5mpTNPE23Cd2jHPjlKcaYP5joOVUDBG7GhpN8vRE22R5FaK/w9TsrjtOc9I+ZadE
v9OdWghEKuU0cn7J4oclMpQ0GR+xspj8cdfy0L/9g2tteiGB61bZf8bXPN5WqbSLcLS7VAX3kWrV
MdI+wi0mRIfxwHLLriLCGor27G8omf0skf+xEWQwqJFiuTD+Ibl+Tp5h/7dXzln8K6gS7UCgWHf+
LMQjnamyYXorh87m6/E4UNXsGDUoCn8OH9AiTcf8CVqws3ifxACKhaTFzSg6n4QgjHo6+cMXGmQd
XuNeGO2flGn3sNmrdZjeRVsUb2lA+qjir5XILhGUi7PrveCvqv5TAX/1y1UqW6/Xpv3gpe17yz3k
UJuT7Vo6UFHXrDSw2gpXnLrxPolzCeq5ep3IP2/dzQF03HdRX82YwkmzbL+a7gDus5oUQw3/r1/L
bknprE6rh4pJq3azAVsAkZ7mXwhF9xidbfTCv72Qy4PGTIauMKDvl7FLNPNZ3eXVMCdA5Vs5kAlQ
OZFv0y/2ZOR6h80M0BsU8Hfk5nruHQnLbBk4WQU+JjUDgE4NnYpa/50OiY6PYaR60eYDQEBmPB1o
lZUYSSEknzZY2l5GQMKBKHo1foVe4FrPg9luzkpeDzpcDqLg/5BsxvKlbCCiHW3kjauODuLcca+Z
y/ov/mUlaPMha4HiIzoeuGG2HPF4midLhuBbZPBjth/+ej1uU2sWmu0J/cJFWbrTvqJo6mvNSpsq
fs1Kf/ytRQBSk4uxvVUyVaSiYIAMBRDlpHixJ0scEoWoMTUevC1vk0E9FTVVOPKP2omzt+FzQvuN
IZ4zSCNTO7Jm9IbpBlr5lb7bBLu1DaoZTLO3aFwTlYkD1XTM46lsn2U0kRyBmIiIMZEdnH57VeLL
iK4WOp35VWbxY8hp052R/WzHXyKx6J/t1OFj3bY8oKqSMvyMB5YnQ4i6iO8vcZ695BU7atLTyy/A
wNFGWuCIaWLLg7iYgvSDLIaOjc+o7mtovVVPgoBr3TDHjWFJGu6IbjqViCJje5kNbA8sem081zSz
xbPXVbIOib0VXJnIaLceUSPHXS2C4hsT2VPjoLh/0a4BS4Q4yfsQMUCDPvfxaHv6imFDvwDjweIP
uk2TgPuqobvNG4K+Rl3XuQArZb3/+/k3/Aqh7cSXv3H4j/V+vIIj1fFHaCsZ4Tu0yriSFW2TyhvS
T8VCxh0khQoaS0O76rHaeo7fzRfCydik8+1Z6QF6iBj0JpHCpQKj5hvLgkOIy8ggKYMTHE5ianzI
pEm6t6HhIvWEkbieHKRyOSR6CFYyelcSwhBLo6etbYp2SmWVaOwdYaTMz67QRqFy44BSX7Uk19St
O+hz7stQZIFiL2QpONKEbRfqEb8h1T3O4zWkzzaJ3oKbT4Xd5XPJUo1iWBavy6lUGGE2XoqN3/hl
TSD8VnIS8ZW5jDDcFFKLab7j3hQxlNsRUvZyWDVvtm/aodAtzaJHMqGwwv9V1Wr9dx12KMDCQMiW
wtFNcYVsdtAxY5acQbSxCyb+aa9w6zg1CKKaeL8pSjLn1LapQ1/QQ75ARBVO5/FYItsFfRkOusAo
899W3gSj7z2TSFuflxZGqdLG7OKqbNjn6ZpkGDUMRcM+mDKfGeqHkwScyTtdTyxx0NxEjj3bwPtA
BLNr8gkhlw+/P0h5RuGI20bjo9P4FRSMFVnP9NJK93YQ0VlBD7vK4AwmfYgXGfVhZTfSTtC7yes/
koyAnmhwtlt7KnOrtHwkQZ+hY2VjZ4CWmDu/ef35To9sZX9aJSxdzlcYqcglGmocJiZNPf4jyxEs
cgIzvde6oGHiHd5iGMalhjBGe1Spg9tpsrZKuOtKyz3qAcDfRl16hjI/CUHUWq8i+M9FnNunHVhd
ukovLIuw2gJ+mWcuU+aMckELDMpeZ/IRP7f599a4iz5FOfu4TZ3Nke0zjSTKOIUzS4dKsKQfgKKK
gdYddFJyfPqpo+5xLajtz9hQXboHpiR1mx7GlEbD3tTJIjI4n1tQq0Eix4u7oiJCrJDebxROF8Aw
3SJm2VtJ7ZXJOV73otTBH0yHppTWYCX1Hxg46LiCrD1s5g3xU9OkdwMJKc0KlnYCik5SiODIulYd
r3N/RuMn+M6DQ505buQ3d6RdQIWy0ZK65AWfN0GAD6h3qnGyi6UcRIIduI/8Bnwnjrxd9IWJrcL0
7ZkXM1tsxqLLRGXdk/fQAWCnGFpfrS7fROhMp9vhRN60fsF3nUVnxnS6pyJMlQRsRdn7fRKMKEb7
j1Vgf+M6EFtRhZfUpzgwuUGCvluuau8WLFrQvjbn/P87Aqyi52mpaw9T80CprQX6P0Y6UHbbuUUD
/fvzy+FqSfYdZNO2T+1mwu7i9ISL5KZDlGImO4wJSGTAkDdMs2oV+U7T93SPK/Ttt/J94NVykY9t
iHptDWFdVGw7H99ECnrVHpIxc0pYNQbpnxw3jEGbKSzYmJojJwO6IYKJgAEVFxKglh8Rcag1/0vd
D/BeBqO1LR49Mlls3q6LpM7zZTF0hGclGmUGSsREIm6B+bSQF1jI9ES8vRYf5pEdjaO6MKcHxZBw
cX2Ks+ZZpH8q7bHdwUO+EE5RamUpkauYvLky02cefY93jgnXror2WaHWcBVBkVKt5Qr+QMIQ/3O8
v/70LsCrUD6q0l/O4wst2/EIk8ibDcopwG4fDKv9E5G4J0Lq5weEv5qYVP0eEbOB/5QAUhSIyhD1
Zibfuk2cunDb4rqCCDvUlYsCU1Q1Pzu1tP34OMAy0Fe0iMb2ddTwtbsAEKLNwkbb9goQ3Cbwshuo
2bqjbkFuDZs7uKCMsNjzHE5gULy5vTfynReQ7ePGiBAgTeOgTf8ZmZPOV26tj7Ku0Qn6ZVy/hY8t
tvgXyZEVLap2EkyMMmd2tvWZActVd9abPbAMu31DL14TCabe/6p5g3Uq5FBLDEcQVSJmO58Tuc0A
+TK/88P6J037tbba5QJiEhiKKq7+iq9SRkwQHWnvA1NDU2aDh8d8hJXgOz5rEzTDmI7WY11ayBPo
gfOdxLffCMN5II/rwEvSeDJ+NlP2P+UpCrcUy8SV9J93Qd/dEQ/7LtFSVGfFBE+vmm/fSS6h3Ot+
UpbJCbneu+NO08tIrbZkMg1S62DOS8N1cWLsHk0Nm9hNKYDtDlmzBQ5wWoHiiRFqirgWS5jLIDOg
OSgDbDb4v2K88TJjlrTkW8JBqNz+U9wTGYKagSIbQJy6cXPHe6TANEs1n7LBvPoPKEUuSAB3liMI
4er+MiqGRdd8UHKNiJvnopcoip7eCjz6/9QoorufjfYq5zjqRjEC+hesfIdarOpLiZjLnOJLXx5m
ag4XQJkkJEhuTdrsr6NwbbJGDecXfwcSHKcvxcs9JV5tNg8yC19/ECct5e5YAJ7aRpEGlFq+1BpY
CCGpwmerh/vvekAt2Upm05/umS9BgVJWMApeeAksL2BU/M6wNzsNRYZF6hJTA6g7JiKppvKsTNnd
py6/vqjExeBiqHhyRm9gW1Wt9UZ7b1ISf3kk6S12usM8kpkI6SFJ93wfPiUmuMrOzgaCfbcDsi+u
rabulMtf3Uv5F5/nvhz9x/IkGR/9h2h/zl8YcYf8bw/JchMRg9dA8Z7+k/0XwA2yJFLGMQ+V9Apq
zN03pBznjy6wpAzHRvdcibA2us+gvETW3/gq0wflS8W/4/5cXYIgjG9dt2V73B6nGImXWnlT+QFo
ndpLjEz9Af4jXIgLeL0JtOgaZpDbvVBaHYUEvSVL2Vgn2Lb2+4eepxZFggaEzPoNkyRyMc/zzkmD
iy3pNVTswXkbgklRPF2O9O5pZ1VpEUVdSvkhIUoxYgb9v4OrfWYO/qv4ASm68/FFlG9L+4zo6OFg
XMsBu+SYoxR4WvYWYUSSudBDKw5jEgLsow6vf+E6G2CmUL2nHNjGwz0mh3fdkUyRlroO4nyWs3yA
M9id6Nrk1sFXrwo/HnZXu3xXU80pVw6SUWOcozXuSke48p3zZVa3EpN84Jchu2J8BuuMcybiHNQs
GirgckqTCOvU/6Xn0ZLrY6FJw7kxfnWCqshdy+4GwHmJUJberEyWji0IFMwXrKbHQdxTkqJKtVR4
uSAfyF0nJA91GX1G3PBnocYruXwCypDfACpCzzzSmoVYgbafV5KHdj5tT6kDiBzyF/etC+XPWwLQ
UljEu8NViN2Vcu7+eGtfv2zsdP+m+ZtHYmzS7ILKoXePYPBnw0TPU2GKBHe91LgVgon3P/lOR9in
StvNLzIPYOaWgbFTNIRFBZs3TTOVYSfKr+rODYchC/dPRSq12/EDmrN2XuHTUH/JBkeoSp/mLH5A
I8cQ+eg747O46x/Z5DFZJd1qG4ktrTNk2Qg1mMjsC+J7l0fk/+CFprw0le/3ozsr59lrnNi7lv9j
uVQuorBsdcEb8cMWUl2DeaTeSZ1dPs9zL26zpPEFnppVi0ZKrCNqbybES2GYK+Coz/y0u8NA8hob
jlFsOjvpARwWRpzrjIimJVoMgpBNTl441h6Ri5QCElY5cfd3FbI445HKfDKdxBANSR3J14KE/HT+
NkO7vA7ZZBpIWo/XpxXI7iFAg1ktMI2FtXcGu1iLM3sEODeVc1ny0VL3ZkxPZ8utFllZx+dQKubd
CRKSrlKpDqk5eVStjJK0Ju/3Lvb1iaeSY/n4VEQYqlVF9ZTguRg/g8Ra//ZRvq8aOgtklW64+dGz
FVg3SAOpf6gBQUUhvVbBIfn6bRNPr2CkpK5/flCIQfSAK6OvZzXnDmDGLTjgu4F7N3LLYCxYsmSA
sQ7OFlNu7HFXOtqYMkv/V4302AZnmcCEjfLLZd8F0jQnT4W6kmAzBUbTAA31fNXhP+KHUiMt9Wkr
Yx6K9EMyeOkd0NkdyfN/radvxdqU8nhkCB+fPrMEPV8KoBEVrQ15W8ABfPFEyv9Kp2/j5/ie3i8B
SaktopEXPrGoYpfmAj3/FidHnnHgU83nPXXCXP/OzUyHIdThU2+EbfsewpFWIOebDmChu+QN6JDV
cBVgmHfvxY2YmyRcnqe4FBuYT34j/DGSGlESHmh9hfLiW4WwQTQRLkNCZfLGJMPgJhXRbA+g+xbb
E9PfE+cR+pu6xVAlwrurCbgaIPs9TtjHKM5AVZ85b9ImsdKYZCTTsoHFghRZYT8O9zgC/0m2zNkR
hzPe+rEV9fxbfCha6dxV+dtlbEpu5vyLtQNinREdg8U2Z/KvH1ufT/QrcNRAkEonEJiEfKzbc9pD
wu2DarmZaZuMl8dmKnc9MtmovuRD0VSbOvhuaaPL+ckbYoGXff+RocQGSRNkJSDclnFS1/188L0u
40vZ1NJGh3c0+rdipzCAdspQwhHHYmPrwWiCOn7IqevTBdzgWuK7nMnzeT4CY/AKU5lyh7LPL69N
jdcRby6B3+DTE/SoOWViTR8RaeceVXzXqWM4T3Z+r+iikZhuUJTde7OycIgmJHAbnt+fI7MeY/Xc
whp0vr37hXF3csH3r+/Ze2VRasOl09xBWjoSpCHZPmHXAaI/Ua71jo3cV9dMY4w+Gl9oq5pGOD6/
KKMZO/racRD4PC/eXPsy+2SpkPGSKLDmnlkFa31F/9iQ1xjXVQqKQtnjRZYA96Vj3VFWv0OHuIFO
oZ3M5xUTfIbUDK/Q4vNy3yk2xiQbv6c4Pe/edNhlnuGsNnKkH8qq2LZPN47ssgaqsj8/ul7oY/TP
1Q2+lo3gyt7k4xZQRMz85tkCUSLifdUFfkh1h+DCNC65OBxLq8n1h9KixUg2kaGdwn135uZwXpzr
FbgxQWulnWvUBgyKDJ750ne4sgwPJCbRjKC0p75klc0CDhg/CCd6oEAS5AndL3Em6cfRk8hvnWtI
1x30C6BHjY3H7P0KAmfyTUj8ng9epqXmg13KZ2jDiMxncS+lM0ngHQiuyVUtEVDRYAngUB8qp6RU
j1c+vNnhQTgBCjMlVGNtJUxXw3dVY2vlfTRDxs5qNLpuwmlU1pPh+mOpZTonYYPuX3Ml9F2HZkNA
DxpJWJSXEktnR1YKcJXP/uaTbu5YhYrVg0U8x4TlrAcvgeInjrtie8m+9a1ubBPkE7pLUURDahAo
YVYZDiYlRFfQFoLRxY17JoHv1jBKg6gq4C+Gh7tacRXST33LgPmUgnX577r2tEPblaCtW4qBkTRM
7iBzw3RNwcxlgrGqMT0HI0L+8yRYmeBELL6qCHwgDhINCA5Rw5cDLM9ya6npN6RnXnKVxmza/GRh
c+r8gmQLYaO/EJWwswgAVTjqVL/5r6HYJR57U4J4hMDi/5qnDwXuODybHZx+Tyy0gEjBRtdrsV2R
3lP2mNM+h4uDM5fZo6aL8kKmwdKPMSPxD3JACbqkFkOkmblI8xwPa7F3c0uL6AVZahroqIyoZ5bQ
+q7Q/o4WvQVY/zO1LvyCcOjpEKT52uQ3PT9LtsGZs4a+yCVEfBedfXvI5HY9m1scE55rGI3ntupZ
X1Gb7E7qTG8CjmfMjVuw5mJokvjP+1DKqd8kDcDaAH3dzTWP3ZFNL9tAkVft0LT1pzpVCGOqTfBd
g1fGO2hoih8Ggm5ynwRIh8rVZjam3EvszXKuHgS2nNvFu71gJkHQNWnPshtttPhqFi+KZBph4uRj
+nZlRSk4szRW8NJ6DogDpkVCF6kL3eaJO7qiF7obyrHZBvpS5JKh7YFTegRb70u/5L0V6MgJlmWC
y8M2wp804TiH2+TFSZYi3r8weddIL55Utu26lPNJ0ANDWCYcxbI3Moruci1qfYusye7n68/E3n30
nJUzUDPQe/NUCsgpZIrvDSsh1PK+jnWdwviOuG03pcz7geps+sSbJ100ME8K1OfpQ+0FyTu1ytX5
KyoCMtRu6NsnBmx9pNxQZ5XVXlGqMZ64BfdIyx1w9D/Ggwk5bOhXTPFYsgr/BVZ9R46D4aZ8HDf5
2NYA2UZAO2MsLvjdXcK2pcfvj03Lr/P2dhJAHdkg7fyRyXtAgUH5lOVh48mlbe1kfM2TsC9ctnZR
twbI4wNSkppRckXKzXF3s642KOrSJlwROgDY7SSSJkkF0LSfsBiofyTl8aYmICywEJpXTYgoyfEA
OaUMoQnauZzxh5lMrcBB2Loiwk8niMCYq7jE/omWK0bTKzLAjCVhwCQYzUxawrvw/lvK5oAJvCdQ
vOsviO6sjL1xTLOmfbue/pN9ahamXFbdJNHn8k4JJeXXycQ7E+m5JkeLJ8YMVoEKbIBGYHH1wYgh
Tf7rk9omC6ewH+l6qShJiNmVtpnl/4ySw56HZ8Ti31XD2gL+agwurgYAcFjxYDCGPlc9rEWwvT6I
oefJvcwWBzX0svN4ltuK7VzKQOptOxx5Z0Cy3zJMehXz7up4aIUp3u1b41a2+8QCYyvpgzoUlFIr
L6+fePCrRzbWoQhxONaEzkzds7WXBfGLzleNTCUOzsB2l4MmJ5QErTe+xe/DpngMpa99u7CtGLRX
FJv+fszwO127D0DtAp8Yi+bbbp03nhzxdwNEReyeCOul8tl6VEIwm98HVFrQDV5hF1OpgyLtD4tZ
MvFbG1qZMa9el84jLsj+io9CxwDXEAi+z56jXwh0WNJuZg72OrqSrr0OjgEZCtOYwFDsaQVSS28H
knQJ/+rRxV7P3dVi1+d8Zd7zSk87QQ3KyafBkJ6vcnSnCAdkapAEYh4uZnVopQ8/p5Hj74TN2GPc
aRQhYJbKM6CNmmISS5co3QuIog/rJCZ1rejrGSl3ux+rZ+dK9eWlqHW7emIOgmeixmu5dz89PvLf
i7X3IE1vV0LsKPTct/NfmhzcBBuQsh2YIjf/mxVG2zfXGqF9qLVjWROp8V2ZIjCSW4VlQQWnLUPE
a4QbgUmZKHPkl2eMkFlTfNJmhiEhLHSQ0JRK+hh99Nvegy+csHF6GsuvIzTXWbmCln2DTUfR/z7H
lJLmCl8jEWQY1qHikBUKN3M4VcBIIMtoslPVZEspWIcazhr/KzBiHMDzYCd+kakV+mCVQha+BB5n
gyquWPRq8inFkri4SQqmjD6WenTebR8jMFUkE3FZCARQb3G3dKtFqloJfRnSXJFJ6ssIUs7PBPzI
Mg86GT0p5znwcZvux7WK+iRnn7CaAlzsIm4cx4/b/2fv5WAig67CEePFMnr268J19lvIiC7oNBAc
hwcS8tkLk52NYmbi8S5YB5w4XSvj4+BHB7onSX1o/I6R2gFai1lzsTBpDMgmU6qnrDt8b4HXslsH
WJTtgWp/PkeyMB6vv0UQpAjxGM7hcdzA0ZRYzzjBEMTiqcNfjWrD72GsXhc8HGQ6nfP8Ve4H45lB
Nmjdvve7S6qld7bX0pHNrKBd4UpMdbg7VC4usaZC+PElnUv3KWwpKD2jWdJxzCgJP3KkP/Fc0h26
GawXjlMexXQt9Qyc7jM9qLpt8hNnUlQEkRv5esuxdF2Q+7XsiI7Ci6L7E8MdQIRQtNbxJskn+k1t
HfLCMsV0shEUs9SrzvlgNoqPLIjn9ooBZOLfu0l0Qfcxs6/qew+3kTQITRmLkVObHWNChTxtSgHV
mEfOleSzJSW8y3zqoM85/c5YZ643NDTWbtCLv8q6vy82NtB3xg6Ff9kVfQ7XyJPYOcPbuv2SFAZe
oRAzQPyuOhlj2nSsTqtQ2QE8FVbN9lGAw3lcajSiraVqLsIY2VxVnP/eDB1fuTFX1EDvM00PU5Xd
lap2cGXPJL0zbz/JSouOYywumIthR47QkzkpZXR6Fl0UqLhDzZubpAe7b2La2XaV08tF6QpsnYar
YDNHwAdaucGrwE/hRNuaVH186NwsQ0N+2shB0qDomLx71D/UXZ11/NsKCbQZCnz2nUXvk+TmPb11
l1SQQhyXnsc3ZuQPZVVNfAVphNR/Szj57rrInjdMFFlFG5HJUukTzqRFQoymHGVW2RNrj7rjpm3W
80+SCaALkfT3ANQVOjWuo8jFOmMEHu4q6gd08DBQUxh0tjJncaTRhJqv6efF1tdEipcXHj3o+8/V
6LPgNZZ3FA0DeB6zUABM/ZXQ5ts0TmrLF1kYEJpRv5pJayE6mubFsZUBGg9XB1Jq+0K7LThXWpKk
MZaJ/qB3OF+kKuA9szbtexe29PmZGs/TJp2BkgqFigWjU56aHiuZdupcbAkEwYW9W1pKjkCFaW5a
9pkxm4sKU8O8r8qsWmCEVAQr/kc214aTdPV3/1qhb88xGpFL67VMa+3I/aK2KJrEBj8qkWyNlklc
qAzFZ5MT1C4fSasRaxQssl6NGpW3Fv+s5uy0lkCp8adFKFthOEzmKSUwhBo9qiJP8z9D4QdsZatH
dLYU/GWD0wG5wCn7SznLAKBU1OuUc8k3hE0y3/oiR3sV4tw3M9kUxUtv9dg0C1IIL6u+ckcyhR9K
naIuzZstvBdQ7HPjuuw3TF8pdzTMpig9nEHIqNHhkR775EXuskrZVKae2qMS1qbJ3gsM6c+lPAGI
1Osf+cssg1xvI5hIp2ZyJldU9s82uEgko2yQtii6+573tgtbxf9b9wCbO6pDt/3Fd+LhYoIhqxHF
ML4/yOw3mobP9LqUqDcliCotsbEuCOax4DMyvtfSQXDHqaveeJxcAAzBibCY6/qjQFn0eMHrKBW4
sNDnHzVpqt+x/P0Pt2QivHuMAP78efR/iaDCiT+7Kbow51jRNeyB79tCAqswfXwZtC2vDfb8KWR4
cj2V1v//n91qc751JYQi4MbZOfjO1OTDLI9xfqTdDM7NnkJ6Vpg/VjjTiyCL7SMj6MLOG+glM+hT
T/fyAm4IxMF+DWap8SAsMaS0z7pRjTfdK5uHyvP/B+ooaBK9Cs+icbfnEhSCvQxsQH0dohhCNRYf
waXImWOl1zHcdY6K+4hmjZGCjlply6n8WMJhHrTUIIRXk0XTptGbzbin4qjp13Mt3USDEkgCkjf4
S/AIIDMbzhIJPIGdODEEToLrjdpyJF7kPKeKUBGLDwle+ht0GH04FD6OkNkQ0k96p7ZQVnhIgWAy
TRMUlyzl626G6MojRQ8zY91yEoLRVzb5lb+eRJv835AuCaLCja+2oolHUdFVxsnoqFfx66gd3A7S
ovyLQ/8EUMMYJuBknMyrNqt5BzBGbw9+jOOvgBCRqPwxywruqT34j3cT5OIJ7vRoP9QsAk4GTnap
7OoL9GHy0QTfAywG8vnL8x7GyR62k0ch6RsbxJdEkoLlvwa/qq0EvOPeRKezdf8Muzf1SwjwDqP3
bbRfjhcIIWt0U1E79UDd+YtBL45kLGbKGteUsfUNG/Z1J0dx3G7oJqqGsvcDq8pmfTddDGB3eHiE
bR+Fb8wDVvDiv1jctXHm1t+3MrCq4A85xx/5T/rN0mZEUoRwbBSeAI/MpVfNiG9jABrf9xb5dnQ5
NOO56RO9d0s0jzLEM7lUSm0Xq6V72+l6reDNbGtBZOlhCJG5IG1mqSWB235vZFBCc099TkkwoQua
bzpUeloZYaAtdo63sfa1WVA6AE/U44Omos+ggCE2vQGlAF+Lchi28eJWlTaRU2RJNkcEBLCFj6bq
phRVIjjRbNkWhL680YrsprFZfXc2XGM2ejRgVddNQXxAKn8LmE0TEkyf7Paas0X6Iaf5oE89g5Yt
Pg3QnElV0SOt6OfBiT71nVbR+e/jUJ7T17f6wdczmVQOctSYKHDRQf5nYbwfnduk7EPfOrvCvHvv
J21Cy43TF7Lc6qXU5c7WjF2QSrQqyIvqB6wzNxB/DtFlPt5Kl2jjBvRCqbY1s4OdMFiBbfRFyCss
5pbn/P9zV/4b9gWFvVudfhhxfU0Ox2hBjT00OyZYEPpKAaFQVbG30/HP9UYGgHjSQr99b1d/WoMi
e3pguRagt7s2V7aQ35aYUhxbWgKzZL62thNidHrVjI/0oEQVpecbGr89x3rhJ/9axjjfNMSfcAn2
32Sx3zv+iDibUW8BMh72C1bxd9+iym8IVgI9dStGJJ4kfX4MJxtywDn7wFgHhYqkLJVyn6yBU173
gFcVWWoofEy/UP4NRMF4ZwBqAGJ8yB1Dzw8oWWVtEdCiGf12FJ6IJr4e+SEy0kvHRx1mJ/oZ+4NK
aLRDZhNzOaJCtofZGBayFizvH33D48vEBIFOOZVDVJqRZYgWUFdPSprRFN3xuFHdCx/tkiC1XTLe
wgh1lGcJoXVPS/3fpAQexIIdbu9j/LvJvFXQBa4cTo0h9xPxGKjFehyR7KfdH7s2isaoif9+VYqH
YBRiKz95Fhr+xm8y3Ca4AALCSwO8btPUdZ2mmABMQHUsq9je9i3b5EWPMyo7HwjlcKYFTYTD/RmN
0oGBvmNuzdb2QZ7jC+dRhB1qb6qokBKJkndo3aPEG2RYNY7oWA0lQeLY8yK047eSasQUj6c52okK
cVF8SksuQQbCYlxu2CL0V2ixeunM9cuiz+iT/W874g/WAbc/SlNm56VIAdUHfsveobWY5j6E65Oh
0FwPDzlKr6nOnqygsBMzK1Jz8Oq4dQgIu8ytIOLXTtXO2StVUOTtLk0GkiYUyVx6Ddw3TQPTrOFl
nCAn9GfodxtNNHB4yPPNvFWAZHeWPUHHCyH3dcr7xAhbC59I3ODHRPulO2oQpruU/XQIokq1/5z8
n5CSxblMCWW2Uiq2YTtW74WFY6TLXjRVkCDRPRFlqY5uPkkUi9yxW9GtBLJqw9wvoVCho1AdDfBj
WJVYH7W7uV+Wz8wv8ujgqOK+lT3e+IZYZlPjln9U4FwQPliWR20gFVHazKpuS1ZaT0r2WhRbXeM4
MmI/1uaCIpmYwz6jF/fE5gIuDXwxilojCSqJRynNP+sHsBGz++/l9QT3yWVaO+81cw/DYCfvXsuZ
Fhf7ODhi3doIU9OR2Pg9yrnEw0sXKgUSRFQ2p2G8a+ayHKzlYKuF4cQslIB4gPYcYMq6Iu18EphJ
p8Nvtop6i0lFOszGFQI+XJdnK2LF2mJPPN08w67Vj/B9Sai2BTaydJ9ukpvRecSC5QtUExJL8KbF
M+Vbuthwy3xBfF/sSeA/91ib66rcTQO2IHIKqc3Zzc0G87Yo2RPAZ4+COwV7D6TUDv2G8/6gcmem
99GbJlulLEdv1iJ5IU9hRFo11npzhNRx/xo8iLQVu0Kh73H9AtVTb0lmJ95YRxINbi7tXU3IV2z9
LSGaYQQsk25ih0AOySORtbS0aSLGsqI/QP3UK7OF89W6MyRdXayBPBqHDUbbXGg6htmBjwI0pweU
RH6jm1Sp30FhDjTmnZSXlzsxeWpAeC1ykspuZdEMxff7COS8n0hvd546IRl7vBgEVx58CGoTgwbi
mtOIhgpZ6wllXD1sO5vp05mEGce6JLYH+UhMAYMIIr3gzu3sNGDImk9pXrf2wG2GD+OAwSYy7TBK
tns8wv2zvrYXAjDiGS+LTOhannOTQi09Qis4ayZ/42fmBpHWeO+thEYvhAuwAOLBxFS9tCZqK7rg
raSNJ6uBu4YWWUvgeis09pcXnb5lK2ezYxZxUHjX2UWIjcpxjWHfhb7w+KmfqHV3+D67p0tunCkT
KXP/7lF6Zued0d1UiJ+76ch8tcK+ffk/6rYGXgrDtklNcG9hl36d04UJouQRkyXskhUtYgKVrVXW
qmaFMUmnAPLNrGq+KtSXQrkhX/744JrwZjxry8P37PYNN9X6pJkNjCyLShPScU+6Mk0uKTuzvoQR
mMsag2ev7gOHw0iw56O142broAF0+sk+N061H+nPZE3fPKyeqjF82/AcJEZhjrEvavFiWfwEky8g
Z7hqEgdCZvsw27SvEFLdKSUEW3fddkValNJrePKV3vVCGpBt0wuAA4Pb37ISYHIY+bvdff+CpU+f
AH+DFYtW/TW6VW3n8iVHXZCbGbwVhJKAc0imcwlz2wnQMybNTwyLV58wqEugTosYSwY0uuRjkPbn
p71xcm3f/QEinK3pqFsm+MuAKOo7KRF7nz+RdgDAXPfBP9vnQFI5nPQWQJkeyuOIHqSx8i4cvgeq
jnjBbyxa6PPS2C6oEeUvFDoN3z9H+Om8UuFMgJFmGfsa5nkgFPFoy8Xi7fjZC9qYMdKhS9HyKE9+
onZXIfEsClNqE1Tf1FZLzxHaT3HjZgrvi4sIZPHwTurkH9epbHW+2j5FcX92YGjiDih2Hgc9D4R8
aG+KBWnb6WfS2UzKrdO8k+33U5nf8x+AE+Nrx6oKynAYOdaUbzpgCUSp7DJEWG4l+ooXe0ycChMJ
DvwlEHoPiRJRCS8EAKWGKwWRn7/HueFiXpiwiW1GHlxPe/O/NMQj5HkYHUhiy4z60nbTnzYnVKDW
lRmWgCl5K5iN8FeT/HuvOFQH0i65+2nOc6oujUiaoOEKSsdwyZ0GPmus9UcjGxXfFDytWy2eZsnm
3BxTL6Ket+sPc3bRRQlH5ZiDwe2fpH+PSU8QCZ4+OoEjcdo/MPojC+KYl6T98XcG1JLBeXuhotF1
wlW91hgltEEzIrtpy0f3TnS9UJuV03mQ1ZwDL7Zrh6eVCnVpoCObPEqUtUiLcA7XUmkpi31A1b0j
5lcggSFSf8erEf/2LZMj4Z1VLog2DidGYyCbAB5TcqwBKvjB691mmc1lHQGlYl3KC/FS22dRWGTm
+1RhqvUbes0yizLlLnoMkdv2R2p1MBfq41R3smYaZ9jMnS8f9dKMQVPglLPiW/pPaBrcwYO3Hqhs
9KmbPQzK7hKu7S3FPpGG8mxNQODIhfjuDWz33Nk78Dm4pfw8lfOF3YFIHo6mCdmgDI2OzYuNT9LS
oml9g34krCS/6bEHskRqjbF6kWzqTExLOV/pH5Q9VpeNXO91DauV9pJOpSJEwhpRv+4YxUNkWcw9
JOCqQsF2tXiycDoMaqf1XxNfigzwCmplAuejw1f8WkdAKCA7k8ey5ydHSqdgVD9WHsnIJ7ArxXq6
aILxl6wnswoKCkeR87lhSSdaP/ixjP4TKewxmrTNY8QyGhGvYHgdVlhyktzCHw4LJS6HpHrYJ/pZ
rnky4QE2/Hjcug3W83oN1r9Fe9ENRFqYJfOXXwznw9zrHZDF098+mfnNPdByVtNkZ3dLSFP7ySme
CvDuQZ2G+4IhtgkdL8tW9/WznH/pAbvbwEhZAxcQuNJK52D05a42hboJvIQix2caSNG3hM8COPOR
V37XVs39akGBhDPZ51kJPhKM9CZd8gVfSHmPvJQq0K45qpBA5P4FN+gSLBrjrRBnhg/w8HRlhTw1
B/9lv5+mgyCnolnjxb8jAenooYVKuiZkkgRG2PtxGv1qZ5PKUvw4d7XMFw04VO6j+OqUymVJ8pyi
FudjCxTlX1xwRBnmalcPuKbaNrz7WIR4W9gTNW658yNagt51aAFLZs7csoCwEOgbZJ7tHYmxpD+M
i4PqUL3F+TYrjRTlZXIqhkeDK39b/N6e+0CK0AX8uTHZ3Jf849Ve7l41/WEv5BRuhLxGs9uNJ/gN
HEeLHr33j9rCgaM+9L/faAPeK+ISV/eZHyEnXhbgdwZF6ubmJJ+Ugc8P+2RJy51QGPz+9BwIBQgc
tsRen+lFaxsC5iFKGRk/19zRIk2p4adwnXgRULdBzizGiIQM1I9hS87zbvcaPZElrm1aQqmhpd8X
KLzcgYer2R4SUi7368XBvvQZQknejqsFOm96WFTbaR527dx9vu6F9/jDQqvbrGI2kCZntBEgz+Ab
wTilue0SoEN3BlLiMUY9+j6MjbF9verusoQYQzKztwnFgKcja9ecdajzqLWKghHaqvyGcOaqM5YR
EJD2PJVeaE2focXC/NQuLc7bj8jWejfwFQ+RHGj7ywmAhWR3N6pc9R6q0ymHpwVt9VIBjZPc9dhT
RAKbFdYyEa3kfVd/OfK2BB4o4CzCN35sp612ng9KJ8OthXkTudP9TWqGh7RomKg4LNKREjFeJfbO
E+AdmZpSPhkXRB/iEArDi9/b0cjzO/L49wqaTNltFMt6lyIa31hF1R3DFPPGWcv4+08llHmmETdv
PXYxbxdmx8okkwms3oJpzJOchA3s2BxyMiM10hrnK5f6OQIDgk1mPg7bQkQzYkj+p7k9kNYjcfxK
+KhMBaG+g8gGASarSVV6IdMoDvsLJlrbCrVMWyDPsrc8a75ZgZos3ez/gsGCiBleko9BLpQKVxe2
oszBnvmZrecYmot2c/7mCWmC4Ox3Thaxh186j7BUY4X3PiJabPu1A41MbsRP9pRl7H8NBnuYgoWg
MBiKRm6BJ3jtb0/MJ2UNld72wSxdAwb4nHhvYpiXe2W6y+nHkKkAYZw/X2865ToaqNT3Rp4kK2I7
wXbsGICO+e2aS1uCGWWzHWKt/1u07jVfzqsHUhPT7mY0CufuQPYqm+fYIKyK0ZyRiHCaB3G76Rxh
eHjGPrZ3Aqknr35Pr9Phaex4DCjX5v/uHI+oJUyG3Ylxi6nvngEF1y17cPOH610tJ/OfyCUr4j6Z
JblJLtChuluMuxTvhJLnnR6d3NtkMel7cX/1+LBGFGKt2YLgHqMW5SSxJJZLB4Y4TPdTR99k1Xh6
lsPo9rjNsJiQ2gaCoYSSVvh167Wp75eLhX427cX/DOLeohoarURf38i2Vu925eou4G75QVtpvTtn
yeMV6XgsRL1bS2NOsw3KY6ZqkeUvdT8Gxc9Y4C+9lqmA3C0xgO8gl0GBqvBwGGzYkCRHBq+CCbba
Ub1FMgAbtF1VER9h7F6jjES7Oqh8SXfRGQyQDaugKGm0Y1RicASrShaguPM7inTV4dMPLsL0z5Mc
taIe53etIDuYqqGMO5XtgcUi6VgpvwkhsLfYKdmyiSV8X/EM9DBQJk44b/Tiu5eu75X4rv1nBy9R
Lf0i7L7joVi9WxfELb/jbOijIkLqbGL01EbXkGvdR5ytZ0ph9CPO+m6TyP9WSbASzet0ISLcBBXE
09WhYpUCicV9OtgsbgGJLUe9cUHe6HUeLd5O2XDIkCh/FqlMk2GldYAfdt93nDX10tQJaGCttCqK
LfbizSA9SxDAIKH7QaOQRWr1StOIjlGZiIoI3fRQqLnXM6ILo6zt+NjB9DKlt4ko+LDTv5Cs/SXs
jy3TprDGZcMJPpsev5nQHmHs67XabaNGBYJ92jzNjHTOxQBzXpZ+/kpKKl/ziMcOm0AaHf8fnicL
yfDSAqnyovAM1mMEuYDmcuI0FETGpFx79YfXAsmVEtDviNfkdwSHZrX8lsLgf5t2vhumtXsax8Sm
qw7UETI66l7n3FY07vbhojkcBVlYCborUaVIC0MGwHrsD6eN0V3elm2SfOjE2xYRzAT1ATWMNpGO
Qx9GtU/nDLOjoJItk6cCxf8bTWX/QpJHNge+iSPPtXSt6/jFKVC87tgccJNvI8+uU0ehCyKnlbCQ
X10lbrRnQ6u9NhXl9YrRWAGsiUJoYJUkaLIXnRLZsLk4geUsF3XVPpCUVx+Ls9j+JDjszKzbf5mb
nSgCAGfJpLzNYS7DwSOpRghII3cd6qszajtTQESHvAE2I9rkJv+QOzYkcqLYA+fzMdvPQ8q6t83K
CyGXFILTqndqyMjg6fQWgNpRphxXuquCYpJeY/cDmEAbG0rmuw8dtIazZDzUXy+TLLhMRIKmNyuZ
D/nmgrJLLiASVF5ozWteYYyH+9HUYZAKUdvO6dsFJpahZi0BIsIy8DXEmmXuUtNDfovUIBbz84/R
7yJiVCJFsAIw8Oc82RYrb3zAhvigqd+VHBRxhe4c6DAMJHSYv6qNwihOMS2fx5EfmC0KhJSqcxYx
kN7fIdaN5sY7B5YPp7Qjm5O6kpkiRI6YRkRAEZsYYQixwkEdecm6pnJbMsDNjTLYvxhvjeRaPix4
PRTzntOYer34wrSdsRJeZrEqg/2btsV7SzhZaPw94EDzcIs3+lJZyNj/+5LTDvU6zWkp3Db4g5fj
UtJjeAd/ffGdUbKpGSPUXYelGL+ONZ3oZcXvKobvZTvNJ/C95aCSSZXvPcEf74pXbl2luJBWQmuf
cekFycGB5gwWRu3dTwC9ZAgVmfy1BpqYL7Zvcm2BCJZ+ruK/XlD89DZuc4l2FnQiAVxEaWFeZCrF
xONjLgkcIJSw9sw+lCmks9AtxNsDrE6mEFYD5MFhzXfueFUcHKv+bAyQlHkVbYdNocI8EIUnEdj/
ZCFXCvASX2g+XccajsPFN8TybkWSV52IaM+gwi2rVzaj/EZG0qB6Vn5ize8MvgYH2fKd10QfZrDJ
bN+v80b/wKrg+1MebZSLEZ0Cx91AsmR2RO7H050s5GrABEttR0DxKwwqzBRjU9zr5yKso07YCX93
DszDwfh+Uc2CODH/woBln9FYzdStAhGlfhGgYkwusg4iPdr0J9mIGptiGdHs5ZPZszyZJCc6ukjw
m2lK7TQjEjdeLi4Ka/JP+SlKWI4h2AEhhZgrCxWYiW8N8N9ijhZI2KnHBmFffN/2tX5shvHXHOP0
KVmLx+wRnDK8Vgs+zPPOWI4rLW4Fg5tVw9qZof5bnjg71A26sLs1aiddH3uL3JV6PZ9b+GXzbyV5
gaaZyIXwepl13p+cyyzb9ITLifwb3oCrPbYV+FL6Ihad+jDxQ5axaRs8BlxxaXFLrTQU+yeBPvIS
PhBSU1cwc/G6ggNqI7ZShQ5vDcbiLgKnDYlrJOSQiW8mu+dY1Jz5Kqc95ejp6GHO3C+47/UPY+37
2coxUET8W29JFRmn3OkV2P8WBxeqHPAArrw0hMTOW4CGbHPERfhei7eW0eXKIh8DjpebiVgKcHhA
ETeUelg5YWJoCnHxTqCAtXTys5h1P+B+Mc3UzbG8KyiQ0pynsny599N68kkRCP1BhI5poKG8+Ziu
8EKJWBCBlIGtjRrhczPY3GWElyRmHoXW+PV7TJCsfMsr+xTIP5wsUxmUWQ4uM+dSgZ1LsChj1GDj
DYXRobd/iIDcMDLbk3fge7MbyJc9yKFFHQt9rFXK5ayumZEyG0SdELhoIDbvw38foim49OPuHFVj
F0c5yliT3NM/TiYFdnt4MND3z5vc+gNPYLOufny1nZpbh8FTUhlKg1cZBvHINRDfXi+OI3Yve1fm
XBEUAToGGaxh4hm8AvDjqSSXWLl9aIKujw8eJbt/VL1qk1Dm8opqlPV7TqEHdjQYYcvZnk4UeTAb
RONT4iMzBJ2powjClAIrSwua/KHOmAlb3ecPylolTcWDxoEQAuTSyqlztfuvoTzFvgHI4ASDS67Q
3LhoOA9YDJmbEq2dNHQ3Vz8Aex6SIcvx7gm0poeLJikZbulczXmMzPCwJkdy/7F2PZQpLM09EgM2
4H1H6M4t0HQ+xzPEJHQny/4CLgzSG+SmNeZyYg0pS51TiRXCeEAatakzgAObFoTGvWm+th0B1Ms3
TG2T9AW+Q0+c6PhrAG/5dDmN1C3CxwAbhBzabSDlUE62petLNLBYgRRaJKTXH/rUR7Su+6vpcl6P
SqsbxhTr1AnLsT/juyeisAbiTMzpZqdmqxclzDujqj9+Jekg/1/yl48dqu/3QS61cAZ24kPy8DRh
OJKkIftzpX+2jqEy8elcVHv0n1tun2jBPEFj7WlKQ77D+4vEtI2fFqtGCwluUdAToMar00UWjW3P
/qmyd4zrgnGckz9sNgiLiHEy9KEbZiOItpk/9NI6vxzBTu+QanpNrI2iLU7LoqXHMI1k+cDvnkzu
U4U97qKhi+VpUkDXWhFOX/jajA8ObztS+RKe7HU9TOvZjEpWif6XQgKo4hna1Xjg4ot8l9TPbn1v
wwdSIqLPRo9IZmL7cjJeh/MDlXm+Pama3ajY7SHRyrZHukxG6CJgBrG/OPy5tR66Y45n7psPEzVo
B1q0O3TG5brc2V4XgAIh35e/5P8k+gD2Cvsh3bZhmUt8TfkyaGx0e0QzWgfs/SSPqOa3q+DQx8Wf
eOITSwPxXxr9yI+8U2ic3johnkAok37nW/EnXYD8kkOXqs76Y8JJ7PthENa25/q0B+CJJ/JZaKaM
B1pES8mG3d5V2P3FoHZVz+t/7+FiInvo0MiDsIeBRgZDxersP0rMkUFDbKllz+z12mtaiBmoTB5n
Is/DIgy4PpHwLBZWrYKudNOnybCSbVoBnKx48obb/r07kwTt5+b8GZgKMHyVhDjtFhjiW6UBV+Q+
gkPOgmORuZK0VFkxdJZFwIzDQtcTwZG9F17V0BPSxlIZzdc1WcCd8vEuA1ESFTyp4gdNSn6zS22A
UmLhtw3qT3Eq7k5kmU6M1DUunbSebtdn6cSd/nijr19HKpueGeppG72YAXpbFolV81ys3/v78EF/
xBZmid2y0uXM/LctIY3I1udZyGFnxDd/BwgACydJnk5aC9f548P3+d3549avmxppc73Jlzsh15Yc
UYsvmbYB0gUfJvYnIxv9hAiu8y/BD+NlRItS5d8svAhIHXGT3ok0ufiwhQwNyEK0JU7QWEChDmwq
/NW+9fKegzB6sBxXUrIjItmHgwiCzq4T2Vy8hYZ9/tjAjl8tUwiLDsoV51EscJsLqSK/Gz7EiniK
tPaYV6TsjBd9iCzH+MtzuEQl2GbKZW3jeOsLiNKgbR++cLHrtoXvAnqge63++UZevuFjOib7fY0s
EDFiCD7PnX2zMgBkEFvwiwck8d8tw6E0XbJh6tjOgD7YujrcTebhufFkMLvL+XEl+PVdgHF+X7MS
M31fhlPioEu/5nA2LjAjJQyx9d8F5n6v3UUgw7Y5kj8ppOUussIfc3pnqCHDhz0jrohT88N9OWqE
B6lLwrr0nxo+rjPq+yS9qchFs8Lj2rntoBZh9bpQKAa6tkjCIuFriR2T1dYHdhpI2ImH0/4V2gOl
PTr9Ive43O3qU1k5zYWbpv+NUh6HSaDpgJOooR60IWfLL6XqFv2gWezh5+RuQokRxiA1XkwFHUBh
aSFgXwPa0CsyQAw+1D06UcsFH6TD+cSFKyAg85xRx9/GEXjHGBG478S6xvYLpsSS+9dX5alsQLtp
419FHGi08bDQik0caM7mzfn7DbKJug7TLzayhoajU485PwFVE/9eUTpPARYVMaauOvMxMYfj32Pi
NmHvqttDPzvUymMRty9uspMD59FAijCP/sn/Ln5jEgvvbL5Q98GCHT3OauNfq9vZpCyR1qtijfUI
XOWOBXOQLntx1h6Ox+rouIN99CBhTjivBb26M8RDKvBBOc9zB5t9VtrjZ2D4/7Zgu73QfWeRiUVr
BzQWDXxy4ia47qwuPAj1qqD8gz8OXweC+gt9jnGx7gWPH+Femhl2o2y99oY08HVibIPFZ5QPLZbg
u7gNA/hHdltn5IhF8i5E9mo2rMHwtbhjxsHyFvUvSh0/xabSfODsKR5eetrwo31ZsWPzOut7Pea+
+evFxelRgfvELc57UkYhNwE2I0r41wqXMyYU1nfg7vs7DMBN/ioDySP7Y7vxUt9B77BM4W2LAjLg
9AWJLun35E61blUnWQ9A1KGfSnXTAOypw9PEo4Klblzw3CI4sPCepHO7U168HkoS62kKF2d4Lhp4
qH4rJTNIoOiC8X3SYCs8EfLW/7odQ/dFgAy8rGV+3aCGdb9h+4O6BdkvBMe5V3zOm+63iEX5scKM
LL2/9jGVOUPMli5GI5nSSRTVl5r/v2q5CbEBZeWTxZ7hQIw4JVqiz+i1s61lCbVpx1u1phzG/FDF
CAmdxwObtzzhhprg8FwYF7+zJLKP7clNt110BfTqHFbkckCGGUm+4N8kM2okdKW/Tve6XKoOAFpD
uvwBi7x7r1HtUtf8ikvLbYgvpnHrMi9tguI/M7R08qOEo8JX+aROZI0dhecPJ/lVQXBJLsi2iE+H
HGTDNo/aCRj5/WutiZLQspqLZn975aUG8t7bq0puYblzoDd+3fpIe0FeWCzE0wgNwcfeC3hD9vwN
JnjSck6A/okPcDOhlH1Uy6IoJTS+iGHzp0E3CwpfPs7QiRUsouW60edLt9jCr9CFE4V7oKcWlWyq
HWq0BVal2Dhg9/rZc2bU7VNzHSx1vcClT9ODp6apVZse+Pjsx/sgL82zcpxndk5ELmFkyxkH7O5t
MdhxoGrxdtoHW2xZDzwcF/YUWRrP+/KpEkK9L9CpNaw522IUYjDVi4DGuawt+aq9kmAeDnsiABAR
XL0JAhY9euTO0tKg5vME1XjZTpg0ZxeMUMLEvcxOTjbXIqwnbsv091+MSmURR1SPez5mBI4Il04h
NecDBN5jPZXfeohbmpCn+/WQRLBVJ0t7sUQs/vN6/l+/pI63VTTCNOdHxtPDd5DW9UJsWRMXaPpn
M1XpPWpAyz8z1Z4uI9Rvt4nL478mZwmN44IowxGJD9h8b/dS0zNBOa6uqa7TeBrbWjlnPxk3dN0W
tbi0z/bw9okHPrf0E+Cce48uKvg2sjo2etBMKGKrbm77mDrdPiJeuNuGd5mnbAm0eCt/v2ldLowM
imINbqfIR34vdGdqcW6Nm6ELkVmf0GbWQClgZlplL5aAtoLhhj7ADtTNui3Qv4O7Ghu94Qe+NNvt
D7NFG8z3y9JZ7z+/8m/wF5fLkMSV/crXgq4G4kpuSoTubcEZ3g90PNkgw+q+gz8YEMlFSR+0cKrr
96wV2xNJ2aGd7TO/3zycM3lLGfRTf2jmHT5x+KFcysFZI/oJhpfLVfFn3EK0e8xpLiqzQSN+D9S0
0FtqmOytk5ZAbxA600LC+8omWbR5L6K7bYPwES9aFSYhbYx2H37PE2CzNFiRddA6oIpRBkTBi07B
txyXjccXTgtAWbZYQ3Hvoc8vJX8QIaP9I1vjkQ7jXewjPLsGGdkXaNdY8iSE9+XyXJZ93exCGpyl
ztqt8dgDqttisGr3nNBzGqdHldUySZYDeJF/NyQgeU/MEr3VON4zsnrraJxyU4coe2SSVDhC0c3u
V57kG4isYdwnu4gL3ibtqBa1oNd+dt0ruXP8tQwC8wXPrLyYjCmpBEu6yx54Rs/NAVdsoowiuPSO
OxHir/HbImtmY4zuxFMGr0GLrNGNgh683W8NYMZ4rXxwkPARTOcbynT7jIi+BwBt3Y2IQ7KSwzla
T5ectAVzul1JM5TAwcbv41YevjXn8Qkio8MJc+26hrl9/lZ0VTe4Aa6yJpKs9S/QkEHJjAB5MMDJ
BW6JMwwJHlW8Lj1wGw764TGKaUFS8w3PN4aBecvSwdq40TJbWnju5Af4jtE4rl2p0fPY/dZqfb3Z
Q64NHOYWl94JLnP5qQI2e8S1mP9SrtBsF/5jCAlPXt4cOsJxvzHRBC8fS0a4TJhNwheurEvcyeb8
BcQmSkupnJ1UCHvQ19MgsSyhsMnk+b7oyq0icK4QvIqnkFv2ZEqrFqqBWKdJnoXU/F4GWGsnB0KR
WPfyIu//RF8jC39sydZxWnAow3zfKWrjENZwESwkDfbnDgkEgOUQENUM3isiNLvFQFYHumDbqVKx
CgfdMDl8vkB18OznxYbdl7c/PX5XiGwI/0JusHQXQxQKK/5hC4FsuVomOjjmPufGU5tw68sPRCJD
Js3KWzqccxnsI6tbSZHv63d71I1heMUAv/XstgD5jIe3ZzL+FazEJAAqCv7bGaTV03e2rrE41Vok
1hxjk9PD5lgk+eIJLmpvWsX0TYo3oeZC4ow3jFP/X60OMhSNDbhdtIIeelURdwf0n82etY9/5GPP
vHBC7J9VnVyFspGmMqRq5DQ681gAWPeOVDLkjjbH/B1xXN+q4cleWO5e3bJVv1j8IYvTGlXSBuVT
Trw2meE2xVS0OkqhIl+01nQM/1YMe0ON5RG17JL5jcbfJLDIpHU1Fzu6y+9LELrUBc4GdIad//HD
fJl+lEE2ZtQFkii/CRMSZu8JhyQshTJexlvvcGAma5rPx84j1/5vrCFyc6VfWT/nD6bHwqrIJu6C
FlRFwd7eNvGLYtDOD2F7v/v9ronbZO4B52ekz46NBrDNSrR27yZ28MoV2HbwEa70RVgyDYgc+/1I
GwFQSFqDyQB+2QhgZVhuCm0Me9sjgu/2hpmDwUwKbQBu0k/u1mU/4Tl/d45n4sOYvkQNBBir3N5b
VeINEvUmyRhguAEQVaqQbp0mHzJTFI4CQUDMh2Os8wDWb/1If5lN2ysy3tWSR8TEnfXYorUWjA2F
l5dpeTRwCPAld0wKq6Z3wrlP+hYxVGfTHamrF6Ph8sRX0udBwp7KJe758GQ1b2qm8ig+WhrvZ+D4
DzbQQayaYRFIuM/OX8UUUtZl9suSPhqKFdkwFy2nMWoRYFxA5kkd1mjOe2ejO/VaLjwMXl38uU9B
XtD5ygKJNmp9v0lihFX3BVSs5IqUadz6c1Po5Bacbkva1rieCK6qDW71e06l/G2zQqvJ/gGbG34P
0nnaaQXozr9jjqIUfrzK+BLH+/wpii+zoKhm7vjpCufuHgSf1SMtbVzU8RxveKvjC32YZVu5q2Fj
zXPtKqko9BECYg6YdZISF5i+MDLjwbbj76RvFS9SkASgrjcrkq4yE8hV2EqMYHQKvyj05PEjD2PV
4NnqfmG5/q3jy7FdVGO9o1ZUaE/PiWSCMsPOfwzvEZr8Uxqk4g785JsQavd4HYhrUbt6xuIryXVk
fN4o/BMcA/E3HJ//DoWodcqmkf+5ReAdtuhOxfFbAheLtJAWW8AjRC+SQF/9dYN1UNvbvWa4n8X1
Qe/P2tpchdN307MljxKnCnN3dQJ/9IpNStlb/u5dKq4xEaKaUOCaJZF4dKYJcWWQc2dufHVjMl5T
Sy1Hud5nP1/+F3wJYrnRf0wQVKd/Vo93tG7fYwbzU4jzndWg8fij4Pqa598kcw7Nem/Buw8M0mlf
KjusPMcQQPeG3zaV+eBNb10fS6Vj75kUGKM0y4cB8JOLXi4gLFl0cu3qDj34Bx4dXH0y4GxYskC+
yzWBDmfwfesQJWK+ZFKBcpD5Svl8Z6mQVYlHdKmDOPhTuBQFN/lWGje5xP7Hs9yjQCxCXWP3AdH/
y/A9xFzflCnbRk8oBef2lDUeA32ZicH+z+V2qyF24hcg91bSmL5HixmXPrT21B4F8yhSg2zGrkTE
XZDHMvnXo0cBAU5M2+5ag7pyxoVt13nKE0VHCYcxRvGQlsl3IZAnvowY+ZBSySv+k6Sob6Xco13Z
eap9oQaTBdAi0mPVCO9566kBHLvulqoa3nvcFI2JR9teTrldTgN8diers6ygWdiKLXzCgJ62zVdm
5/8dC8v7Ts0uv7PRNejMXj2Vb3d8SkwpvFUN59NLQRdxxtrQbL29LBnRzT0U/CszsJJjV6q0GmOM
KquA+IDMpRrteWyqmP6bmqtMV6whLzLB+72UPAvDovYnyWH/slsB7AWbvywmJNxfDhJNmNkoeZWm
kCZkGgMqpAtn3A59PaC8WUJ8lgQsL3kmAxd6ABKCKm5lVyXIm+p/tEsogZw7+W7vZtphhjrZvuY6
K+w0TBLvdTcYyZbnZh6/vvEYYgJiazFU99zAYbSLhWPNd4FH8NQ597D1G/X+o/8D15yPHYj8qo+0
ib7B5boYuqDM7cBhezsPGSIXCN9qNrJwHMIBAf2fSpmI04Z1zYo/MYLmjTKp9Vg9Y4+dxZPLjISC
aqrvRxrNU9KydDdQ1TLpP9/OAZg9eNLJHFyG6VkigIrGGdcVuZgw1v5tuUxxxdICATdQ0yQRsSP9
j5oprX295QHWj54Rq1y0BDOJCyRmliDqKpmBJibyOmyOluFZQDVulOkznMQtDdpIK11nurt7ygvk
gEv4JMBRkKSbB+SXJjHkvb9ebUfLLwmTS4OsAOZpsEx82w3l2xOo44pblkquDLzZ21lnYWvL519c
n5dg3mQffhcGfIyjx0Qu5K5OhR2cJpAFVgR4pV+yJf99Ajy/aC/+4nDGMF/QVl5kSTDJYulWmfgQ
p3pr2ELjF24EqLN3YrxlwEDXeVN74woxrvrxg+F2SI0aVbMkbjyX43ZBLIuDfMr/HOhvufusTaLt
FFB2osiQ9v+zhCmVTX1DHoRK1AjNp5a+QHgIpKQLuAX+4wiS2c1QPughtI+CCmJHwnzF+uivQWxF
ydmdrVT3uzQtAlU3k0kRB8FdiRgjNMlvWZKJNf55HekIkek90UuQ75X7HDwkkJLuIcn8zl6Tt+DK
odABPSpuBb/hB2wCtlb27zgSc7Jw5DtccH+nGS27nRy4zdXpcmdUhrT3aRAKBttcpmPS1rjhEBkT
l4PSZA4in87fYIvzRzUB76TojjGrZWX0mjoP1Ksr+uGgXJXTrDyaKHEYn9zBk+zeDM0QcLH2NDEV
gjmJV9maMSDcnDNnHjjg27g7jVENsSC+J0FbWMb++ZBnj77QEAcW3aWgeZa/jH4uQbotg6l3+U+K
iOyTaBaA6USMwNrpxgzEPmVArYwzfU6ic3/SvoLjycsOSk9ES+5RFMdvqBbbsAGTzp0iptI/eSjW
vvozaLLwQM5Kjsgtf7dlCl3rJzgSnBTk6s7shZsRJFVMocVbNKdJBqqk13pB4AetDh5BH4Ebff9B
CEi26jAjkcsCFCZ1h9/Ge6xp42vfisrQcty8uB04U8wyrRufuKz4huEZV1DhmwsXg5rAqw1oWDBx
kO/aUWGpaHXWq5QI6TvBHtVJeBiIFXn/zBCI8eqL9yD8z8V3HBFty24Zbc4we4UKKOGtECykArNA
s7yRJ0EllphBrmjHL6Kp/+G1AUam5bBLGaIHWqVAGv1gKV0tFfZ/q8U2cS7Gu7h7orULl4BX40el
eSA2SutV9NFdj+Zsc0/lOYLMp7LkdEE/Qqp3sKx5tdx0nYBwtPCWQQ7JrJXACbKhZq0SqIdw5YJi
rW4IQ3gBrNQC7s/EPhJECTOwBo1XPA3fhDKYKbrxoIflHmYqIk7tC/FMYE1d3wmq79gxJy2jJC5B
g+1y1RxX5pNYk1yqyBSUevps90YY37jNhEOCPzlGzaD46OBt/OXF4UMiAm+QfrGB91tHE/tCojyI
d+OoVIORxMI49lNnZZ2JF6iYJCZo5Yc3sn641vH7phD9siupHkmM1IAVkwHkJIrPKQxJ9Lh2/zWg
ZHmrN91Lc5oZvwBF4q4SakIUccC5PGLGYfK7NykCtzlx4Mb+Ew2cFzk6zQgyMEJlatTykAfB8FzB
lXG2ZEmfnvt+9j25vz4Lpt6J7H69nffcZ3RLfB18XRifWZeT/gO/gI+ST41P3z8rVgPvn4o7caTr
59A4oPjSueJHKuP/JfQFcUb+PXUPC8hW6JXHfLaYiPVjhZ1/x8G0IqaGkYyxvDQ6B+UxkZ5smQNM
/4YYZ+AAuZ9XPQZ2VLh18SI12NhLcD+8RJhHe4or3BmNZNjYhqZi4ndvyKH4I+L3uJDI8X1N3Zpk
4oEvIYh1CFeDrqsajxAicWr4iCcRSIRslWHeNf67+2cqNr/exqrvty7dqRl0PE9D+dLty8SjssAv
f+NhJdysxgrsXEarR6YOCXDBevPICUGsYytBAE7bI/7Wiv8SZkk75v6HiWdVzTvK0bOlGpjwhKuW
OATZIvdZY60m8RSuEJUCUDY2GmrAO9wAh8KMHWsd6mqS5aSvIiKeisHovpx6E+K36pO6id+INZzg
mesVDSEjeONfRyQC2AYCvXth9atK9DHUZ6lzpKdeAVh9hgNfwSJzgHMyOveD4GpHd7vrkUlxSuKK
QafbFsTxcxZKi79nKCpYvfFJdnX9rnekzz/iuMa/sJhHjZaHVraYFZ+OkBQK6O+RnEUHVjAEu2EE
aKc6Xmc5txcs51F3K1uOQZlyiWZXSCJsquhUbqJbSLDQQUeuOMU1kfVhzUCov/dfYIjQsaEZ+ppB
c6Rpj0f69b30lcDUa1/7hWOkw5rOZIoXithr5bq3mOfvoIAqhmAufcdg6YLBNg63DpDhWHsWYHJq
VDJguDrd5SvqhLaxdepV+pvNTSwIHRtPNVV0EZ8vPoW/SuwH9+75werOd3ArDLdmP6AJV2Y9Kl1N
j7POe0vZ1jOA639N0x934gg/+MvUS+rVTZOJPpkDSw6fEPp+/gTC8gJQe/Asy8Yp3J6PxlqDc8RE
u4Jlv2BQyc04jd0ye7oPbr2RYNNFwIFChlPuf6Vj5W+FCxICa6ADWYpHzc5EPjYU8NTYv4crIzuA
QYdmm0Qah0sCWKYtnBkz42AmgJ/LhEcxTwGeG4t2C9K2kNeCJbEpDbFPrznDt/KDXY9OLxl1lrXJ
z0erRdwlBgyOsOB9WnSD2bNoPjUSkaPe5EWOSxnhlTRTFERHcGt95LUgA82lLoh7j+FtleNKDR2R
SnyRilg8AU3YdMPvwD+MIqf8ADjugzFC6KZbqT8prb0nfLFMTIei1fIqd+xJokNswC/k6UPC83U8
NlxMeo+imf9uc+sCGUE64CiHI2xdPkPmpNpTOKg6CycK6apdv4bZ8oHY+S1egdviHCAoWHhlP4GX
Dy1awC3egyEtEMd5XovjsM7NC8/eGBe+sPLOUuwvoiOd6zc0zai4adVydRWGMDUlpXXSHMTYKLX9
63nPW+weLPukjQtWubCanQe2d71g5g9tzvxqD0vfkix33CG0Qu8EtYUtqO9GnPZiyzAwrjZtKQ/z
C0HmB0wMnqZsHRUUhnDFd45eYxqE6KQlv+xV3ADGBkB4RWaP0WFK4FwokGYdVchmuryIMEYoCA6q
bpgHMOmoZQimrd8G35tuOlGjtmiHdNj8Tjhb9dyPZuN3XVkHDD6pRg40BJM8Cam3uzZilVESUleJ
fl7QO6avmIc1sfo0f1Hozuckln9RUxvuscqiuqVMXJ+lwq08d7kHOam3p3FFItPuLdIfky1t7MKj
Xz6r25pEGFLPRaXpu/dsx8UTHg/Adp9GeSeNmBJ7BJvjUWUbPUlbe8lASn4tPTENzhRXE1sB3G+m
MAN0v3+cZ6oDhzIyU39Zug77wEH9yGF0kGfOkn9K9i3WREg/Wdp0eZvVIBVRqmdcps+m9U/VehWE
R+RQXdBJsDNyUl1KLu56viHjwCOrEkQnJ8DfmUdjLR5Z4VUGSP6ir6j/+RJcxZkb4g05OE330UEC
xF2dTQnfPMn2thVNDysU6QaAjLXxV/QA299tK6854X3S691GomZD08An9DCQG2FjRM/mCxHXgZs0
sp8WwdPvAj4xssM6GufoLh8x402Yq/E2elO++PAEadIdjhvxIpGQUWtT9QdUbU97B8o+GOhxizwT
kaO9qawFcPkgYBsZuytBBKGDeZgPUuDy6Yd4rdxcu08RmOwqqXCi70APW8k/EBZcuX1ZegHi/jav
Fxy7nEYE+Uuec0kxjX6VpPcAN7urDa9BjQpiNjLTTtDmbVwo45hFySW6iGMdoE3ZsXrfRmU/ydHw
oZCTHQDVPPTkhqTU33nNW5SAsFG67wU7nNJRCYDnfMas6/RwG6klk/V9ZwPzINgFHyN4ZbGE7pBZ
ghomCBQ2uzTeLhT1Z1ozfjJG9hAm3+U6sc+pzpKs+dhDuUq0O6fGxr0Mn/1OO9yOqG9+JosQEeP4
ivooeaUcfzaPHHxyXWANpyMG/sWyzUvReCmlQHdzyZnD1MiI40WzRivW1M7BtZ+ifIYa518fgdR1
C6Hxcn8VT/6rvfWIdLWFWCJXs4OZLRR7eF7cKl4K1ONo8pxTy0EX5zr1PCWknbDikHXtvb/tBXwC
kpuoyN+P1ATZiORFfdKaZEgp3bMLuqRLZpgtOir/gjf83IMHofYfhN2CL/WG5zjrp5kfbAV72TCA
n/LsXfwhomZbkmCP921qvX4OwEpn9wMTovM5mbQ97nHQEtH1afUx7xvJxQ4/qgpfpM1wTiyElcyL
Hucp8LEbgCRHuJ9zSL+l7MfZ5SoETVIDYf6KtYvT6oMXuoVp4efrTvGBBE/Egw7Cw+1J918G7JB6
gvnBIR7J43hPXGP3O5URwPPIYtEPVfmIDkH/BsAoLMENIg1O7PPaVROq14GjqxUOAn+DhZRXTuA+
4jGbR7tufDHg7DHs2UTT44dWsuBINgo2jn9MUt5vJAp+GHwxtb45eSl5kcL8n6+XcCKvoCQ35FSi
kjiSOOXI/O5WdDuYhRbOCIyWFrftmK9ZSkpyQw+JZwgPWINnP1riMkJJm/w/tkaO5PqjUd8Jq7Eb
+o1m5Hb/Ydfu2cKVYMZAhfan4kDNvQ+nkUQuWAKoQM/pPk237n0Cat+Htqpfg6yz+XWaETFcutPb
3U31lvsPZszAssFH9KIrYIchca/W/0FMYT6BlFUXTgkmhTNDToQm/+u52moKz5GVmghnetd1d71w
SLUZzd43kIaEhH569BoItduSzth0IDzy9n8Sq5QTySpeJZ488FBwHPZHmFJWogWyCmvjm9HU/fto
NkHxgvXY0KszIDMJpz5JHKf+j07b3Ih/VHvi/So86KXt1szx8me/syoESRHupMqCjF2skBppErjP
I+5ymTuinrD6ZeVWhGuP9n2xSEwG5uMpVxPch7SNO/OfcKr6STCDFsKZWj/1Gi6Se/d3oryFgdpN
CIpyHlf1pGggYjgHUQbol3lwCSyo3FnunRNC8zlDW/rMbENIkIEGJZziub93k0ajorl3cXgJvK+2
fye6b+/65OYVjRd4NR9ruRfN10ZUemMXiTlaDEWzoCnirP8b3QMVvoJbD/bR50l0sTpMfS0OKBWH
akuQpBPrxPbA13PYAJCWxxyErfsJ1vZIVAR4UTni4qJrGft30xq3Xhqx+th1775DbQpheK48OMJv
x/kGXQ/MN5sKDXmtimsBvRD1cyphEPqEX5ZcLhAMGi5Jtg3zs94eYfK3GFd7rBQZODc2tEgtdD0r
9hCR5CNY0ttS6pNSXL4Nnv+CT29zYr4NP2UipDts36E+cdJJ1J45iX+si+xe1I+N32pzqq8Ui0lk
gK/wM/s4rz/j3oC7n621eYTnKfQpdJwwvBrlgl9IQr5+Z4D4BHiRjFNCchdBgZKyrefLQ7rv97DW
OV/dEc3qKuyX+Q3jia1cvgjgL1vB4PNt6cp5jlaHjDiQslCx3KQFEwAzXlzylSJV4NACRK9jUXwf
GIXiB6zrPOvR8KKXLfBAjRaggQhAdnt4z1OUFp3M3fUqQ9Dg2k8V1+G6PEg/K4MWSQjnbzpelbpA
+8oCzaWeI4Z1pm4qAqxh0YeS7PCgdy5P0tOvjDnxU7Q4EWaVLdjTcg7ncpFrBwG9cPMSFK4Srcaa
62WootgVEieoSdvknlXkqzWOvyJ6v+I1T4qGMWSKGxGLGSFwhN9Fm2aS5i74UVd5/OHe/HOoWZVT
K1bEsD9vKktX7C8ePZfnITHzMuC0xqdNllzFCqgx67uvn18MGslRswkhYalgoZoo3qLOjvlvosQf
K4Mf0OwA7dM3gKohVbpza/I9vuckL4qztXaJf2dgzManF/dRwAqFukuethBy2fdAT4sp+afSt+LV
l8IIY588VPrYzTT356R7MLCPu9tKx2L+FXJTMMmi/cXqqqhwRl+zhSBvWQxIpHOYW5XzZt2ewaH6
duCgcLQLNfwTWjdd5eP2kIO/dLbznjBIs1sYhDCcI/BQ4QmD6Mxq0IeIwCkCRy0+8FSGbvnKmpkm
lLnvowPx5Xwtx8lHQtJKssU34U322d86f98mKP2DuUPku2F37Rxv0iovaK/U1++hJWbTl7NjhsOb
UUeB/LTSJUy7GE+Qm7L7p5qI/q9IKDcWm1/6z4umfkHY8ghcyliCuewrAdyLZHpTsiI59HjISwUH
ZJGvwa0Bq4I+OZq+jeADI4qDf3G9gIjg/PI+tKR3fAI1DEfu4l98QZWtiAjFC6kmyme4/yMOdPQI
fLm6IKofK00GvEjSA8xCZOnP7oYz8IILuS24+2Xln4VkOyIlfRM7L7PwPjBoR6aLXZPU0rYWOn4n
gZxN3NJNK9Qah9JwBuIo5hXldKe2zY7IoElqW09WzST0RZb4JPVzESyZTjucZHMEnfaaNGcDfJV7
T2hStdV0pdRXQN803eiyJmLI5ci0SCIBJThBCV9+SeWL8Vj9EIBBw4sNGPKC+jexRZY01tYst5/w
RpKiBubHiCEJMKrpEhAfqwqPJ/5ixpkXI1SgaqjXtjopfeE1mzk2fLzh9YY7i64WfdzIy8/Ejqy2
YlKHBmD4jLhcwyfyFpRnWL8enMD7M0Mq3NiUhONSXm2dAD/qM3MZPlGn4z/ePBEc0fHSOYZEVwRh
mK0reFkRPlf5yTZCHMxUPg0TwwVntJXM4REYf1m6sQA071/3PHPwRTdtfedMjHtJL2MiRB4JSx1F
9D6lvdPMc609+KEs6LraTNJhbF38KS1Vv8Wc4o0y2MTEj5e5JF78Mx7S/bQZhtsE1HeNdlQY3FFZ
QuDaEITd1AZb4Z6VGZT43qAZoxsxtJs2xaKIoKPs3Lpx3XtOP4/atWv9zgwy74PO+Py4CIL2o1g8
6YxJ68Rn4XXS0r2wms0IIrGheYNa8JcNN61dQzx7ND/VfAC4B+j9DSRz6Scl+45gf5jyBwyhT70h
kModamhv5iFnEtw0OzBoF1UrGW63glZOeMckY0cprQu0RoZvZrhKGQoMvkaNimagBVdxWa1prWLE
XTEM3VNTjiIUVnuviiGzYtEyQQC9m9LFkk9mUMlJBDKsWYX9jGRokO8TWTbScobnZkLfKEcYWQKp
XOP+1hwoP6Nb0ZoR9ZSW7XikTUxXVhBQEjFNSVd+Rv0MlxMbpVY08n5RPYNGv756qNLj2mdUTX2t
GtWnpTQAf54L6p/HmVzoZnjNkmTO5MHCxnk4psnyg+dxFok1dAu+w0b3zZsfnhAKG4HYn0LKSyrN
20WVrFsi9ORTEDjNcrt5fJ+pF8gXSp32FTyDZWA2gLcvfnugYK+f2iwbaTBbzn7oaENLn5aHjnIV
d6iH0SEA47AaQQC/KefwZKFfNi0beWt+GRWaaxJNXEfxklJ0V/Mw/gjYhSnjkJ08OyyfpolWOCNN
SMY20kWIga6RIpHr3zaWsUlmzxDGklQjE75FQPjQ6OazTp8LQE367Uio0lhV4Q63TWHx/T9yrte4
sfw9maglQeyVsShX0pwRNA9hiTBXWUgo47kunvUTxwT0f+TAXYOL2AZ2tCoXAy+EQh8CraP3an+6
GbJk0VGNaABQ1TYi9RVMZ00JAZwRD/ar6CqnYdq14F2PQD0XcNld3z1a6FBHLPVb21jK5UBdqyGw
fjHy8nh5M3HPkptIXJz8caiJOgjdgh5VJanLFpwCp5dfxJksExyMDdMrJnM0QmNQch3HPoBtACci
pjsRZJrDA961hrLFbSQtT6vzuPbQYioVMBRF+pYmWBNkGNS5ZVflH0jcSS2eBYch8TesOmrsICgE
4cei3VGM9sX1pbdSdJj+0MD8juFNi9vkNZEk8OUa+T4fEe5m+F6e5CJ6zEsJgPjcls04x2cDTThD
ybpjwW+39zUpq+QPHK5xd18VWRcKOXFS/lrcM1JLYvqLpRYqUhwFuxa+igc7UbokJ8CDoUexaPdn
uJ3qmsBbzXK6FRi5n41TX7wn/zLs64dRt2YKfamteQ1xwj12NuIkekTvJ3a5/y5x8UIq0pyvZkH6
xsBBfaoms3gVDoNg9sIoKf3CSF75WcFzgnbwe9iYEPJk7wEwfXrzxyGYgHtsEBfpZKGrRLy1L3Ez
TZ6WSn+hSe4wfx+EcEXWb+Mxha5IY+P9fVJFNdIlWERXAma+bue7uB1Wlxn7ENw9HtRsoDfmQPpe
3udFveFUUFtqZqA2A8b+LD9U37Sn0GlOLHXc7ka0LmD3QlkkY6fr/6YEB+uCMDA7VleYN2vdp5Pm
KorIIKv8lcbV7dr2qJphSRr+D4oOu1786K6BF+8cPBQTOp6NglljoL2CGojUhlzGGhSsMmwom4zs
7hNB/FCztBw+ENpAqt/MO3ILnMIA6XbQNFEL7FX8YQUuiziCZJ38Xn+yjunnUvtrkGq+WNY5ZRme
zW29e+vxW+tmu+4JNWpMEPFvH2/YtZiPXMF7kSVDp9QN9LizXC+HN1BaPwjGMNr4rtGSOE/wlXXA
m9efXTlpVnZo2sNXtDqCUdo/LWuWGnZ0iwSjoLaJPiIhp58CPlBbDMOSL6nb8WlpVx6u0T7VfbA0
PDSnX6n+NXm0bDjRfjFRiS+L0ozdHrar6uaGDRW7M9FdSFASPQXU4ZWVvPqVYMbuzqa/KYg4azgl
mLaLoHrv/OtOuFA8ZQqvnrvSP94yxkHsBPm2f3LCiIL0tFnFQ6rlTW3jZlZM4zZ3CH9qbLOY3OyS
4i5p7WPxlOq9n87F6UL0UCjfW0j+nLGVOgfOpdgm870fhU/MaQOI7mRJSdts2LvKjjWo77K8fiYD
/qT5taSVxXt/PX3CkKgrJp/TZWgvl76iEk6puIRq1k1gHu2YmWzUNoGM1HlydKRAGPbu/gHQcrlz
NFe8YuuECnzQArlW6tNXn967Uy5kIQz808fHYtLoDd9Rn0FWN1iuMHtZlmhXebj3ik1QuARSxwJ5
15oAsN+W9+oPsms6xZjzxKRvfHICiP2w+W84BTbP0ZaBlOVbzSGgfd/+trd5B0ig2KDUNXOcCjfV
x7MUqnuIUw6Je1MGPlHwdsfAXNbplVS+1fz4hpYA5qfmYhZiqvphpVZASsqCRqyYKcR7z6Iw6Z2w
S8HujRk/7A6gnBy1AYpokEQPZD6zSjpwVaA90KFk5Un3a6wIpq15UDTlOfxStSYoSV6XxaCO/Kwt
dPzSFfeaHUarmkcwpMnenzieJuxGB/ZfPS5FUBO9Vprhf9uRwwMl79z9ELOY+b/0gOLop+q2bYyl
UGJ2YswUJoAuTGaY7IgEtxaS48Z10dFkbT+wbsYbb4+hFHc84EJUZFUYGjU2ikgivznhHHppMTDZ
BfFzohp2WOHaqThuIrtg5N2F0zBd88RKeQBMh5OmLh5S6loxZfjKIRtY7DCvWSGLbMlS4q/ga17G
ynVsjp1b+Xt/fNxJewOnVhLZlaSIqD+dq/xexbm0x0Gmynm9VKHQnQupj+ST91na2JHVy8hvdkhk
DGGfDXyWzqrzrIbW7zf7aB3j8mpjStP7/hEkB/+a6hJlW7fPA5LJm6k762WHU0kTCsFBRqmnR19+
vIm5G9DopRfskPlZ+pFUGJjFKoybB8wQCguooNcL31+y9BH0Be0mEaAjurztv/nsD/lfUg2bT6Rq
RnqP3pgaoJ9PioAzz2CiIypVaalhJBbfxnopZ8cxkopB20aWuUDKC6YYGUnptR9zXweK/N6s8XoQ
iyYOk+QcTBTSsUSDaKJ1bDipsJjowVFbfyPx+Gd5cHvIo2zcLfUbP5eejCAIKuj7LKFynkaock9x
2XL/GwFDVfVhwsM2/OQSG5l+sFzE2F1zjSOXmelZP3PLUHfYh+5yglScov5xTeixcuTNNYoLuTwV
waIzSS8Vppxu+Y9DP4K/rZmwhhFzWDxTCj+MPKKaWboMSUzd3DSFHI3fedUvChfKDbmC7c15zaBF
wKn0xrLB9bt8/eP3VlQE1WN23jCHRzAmL35ShdTSBJ3xOPdE3J607PMwY0c5YDT9Wn/QG/jZAhnP
i0VTxsN7mNE2M7LzYBx/eTiPbf7UKGRj48Mha/uyWVshGuSMfaBaG9bPGXgiV9PPUJCOBqWCggsa
0nSYnY+c4NOwGNZr87um2vGAwSwl6VOw4G3EsshKsCTINuhEEexPVkPSJriMeJrvpjuT9io/iqhH
lU3iCPw1O1Kv8fam0piUhvJAXZtP+AEwP2EWtJOsGuYjctFLU9gAZ0xmkMPXasEEoaATXYfemeTv
BFgHyI/Qe7rXAp3PUUZ+JbhsAjiVgU/lgESlwwJCiWnS/a7DFO1Gn5qlUrBafGQmV/HAUVV66kQH
UsWo7NtOa0mJRUe2iasjwviiW8m7Q/6buAUDBklepCEBwAfQ0teDyBVCnGUOZLc7axjS1jqHagnI
4EtOaa/tNXqn57Vt4RpZCt/09ivl2X30u5uqcxCaQOiGt2s6lVCpjzyfTkaIz4VmdKWcfOfPLvTV
GElyRBW91VkCbiyzTVD1ghSmjsfcyG/RsCe9hdkU8x0OzPivbKAqQAHHz+PyjrJUatvzZwvkz9/0
f/1PnVSrxvKCmRW1esIL0c6zqgEHJCd0Qm0NSsVZquS7EvLyIi+icYi8Utyw18EWQ0irOV1LWlpT
VD/1gr7xDA1diXuFNGsetfnjGrZ7spxPwnw3DqwHvzPPH2RITkz9FHtLDCmRTVWQ4dKmz/bQDdJ3
sioH9o9p8cqhtMcoomzVexLy6b7yhGm+62bK44BqTbIhuNRnuYhhfujP2APJhQkxrql9R8dO+p7s
4lUd946DoQ4r1p4vsZiIKcr4diVFT5cWq1RhAu43DKpvB+SapInl9od+9hUfWEJfnTS80j+dO28o
P5ke9CPOutHh6aiMpt/xda4rHvYLcY8uJkVr4UT3hk/WuIUocmiCf0J3fhXMynGkl4HW7U8perS9
WWtRNJiSqvjDDmdHXXFy2Tumzn+fXOmK57THR/M1IUAdKL5+W5VvIyk4fA+xt0mo+mWBVVhTvqhm
0x10dO9k870fnDQDfQ/jKrEiD6m7cbzZ1vZxTAb5/nzY/Is7L9zI0KU6kCWjhYiqhgYxlN1ofzQE
bfw3g2S2nGemoUB0c/quRz3FD2ETFPa7CyqIAA56RN8Pgd+d8N/Jib6wP8C0w5BsdSizgf5uNJ/d
YpaTxdvS0/VQJNu1Kgg5KrsQyl34KApQp6rARidVInddcaEKYZfdsBAFlSZzR/XSmszfLa3x9/bK
VAQuKxMBB2l0WwEeCHs/1pT59fy1WqWYPOzBhy2GGw998bLgvSBazB8y7A4wc+It+iUMlZ7XyJVD
3nuCAB7DkaFrFpaK09bV7Wmf8Jr3VJltq1LX2gloEwTj87xiOfJXfsmWDqkWhLJ5wR50YSI41tdP
ZOlNuvyM/iP7vUrF06CU61WOiZvTXEKji+saguWzalwISzzijbBn403lEsT5cEhwH10qDDGj/FsO
gxRbxF7PC7PxtsQtPMA9obDPJ7UjYtHlrJTJh2dBoM4QmrTjkGgd9tK3CJnYQH3KHJ69KGTmk6p1
Qv2kSQsOX/0gJVCTXdiatC8tgVKLv7f+erE23bZ51nRCsv9tPdQLTjs60Flkc58j4zathPpEwFQ/
cM414hgu87BwqqbWXWS6HG4TVHq53/CXlK/Zv/lhmGZML6GI3JmbWemrJXsZ816lTi1dvSZI7Qhd
6vSNtvvsAZ3fgOQE0egabUoraJS2MTIbcwPsyXZ2KJDTerJgERswf5oTTPXHn/9p/mHMH6LkvGQe
RHpxplzNXVVTJSlilYsWLomyMJ8DFNa89q4LY76LtMQd139h7QOkT92755u+rMCXOuAM7Qh2/WYr
Xmp1qSdtvxAYCSYE2sO5mG3L/3CBtmYAVfnhotCX5fY2vLFGqM5Wm2iPNAtf8KFbvVisAIYcBAC2
wP0VV0dcTL/n2rAYi/v0SZpaQVP0J/UshsuF0dxJ5nSWoTTV/D5dbu8SxWlaVHolhqK84gJUmYDX
lVpcTPEECSxhgHCWE4En1a6ewWQGe+RXS9HZxlX7vo2YmhpwtH9AJHiXdacQjB0jCnCiEJIvQ1z0
U/hb6lyVQ3D8sVsNPjJUcOwCsUi9C6YAN7nwBIFluRDk7Cm+EgzbzCxCJ8MD/0gOgkUsflhAptzE
mXETVqfTwDsAqfSyETGj4AKL/VHVgmMp7+O9gFBH+5NkKQdAAN0XM0iujMlmHH1lzpMyyVFrHgNM
m3OlAYtUUHlp4BmbHRZwU8yyMjG9/jTVOSFiAsAr9Efvpw+T96zDVfwLqku3fSUoQSART3VS/C6M
8a870WNqowGoXG8uXL276Eyz4MIqujCJBQXW4d5bCDzgcUMixH/zpEbyXashXsY2C8Z+sVYqa4iN
33kICOsCHt4o3jP9gaB0lATIc2VqYMBdfMA4voVvTQ8WZ3bVb9x4s0fBQqJkAVbZA+uLWOLyfdNh
LZU/XDuACpJxEAS1O2LioeQwPMvtl3LNPFu+hhJCi7ZdCEI+3/S8br8nEorlJBPk/MbBuhZEnf+y
P7N4J+wQSbywGWb9oh8F3hEeuidDpG6zSY3Nh1esqRci1x+8p/Gk375LZOcCG49d4SkGJgSF1QLe
VyHIlSREF7yaLAJnG1j+BRJKU7lhS2KI0e4WVo6DA9t1EI0BJLKqrreDafm8b6QAzZdFYxJFstgA
71henKb2Qu33VkAP/xA8Hc0RXM+YCbRBeSkA16/BcfDHuviQsUYle6gKEz2AMhKQj1lIzx8SlH9h
LIn6XuKQ1onsFvNXu8/nnB8IjXnkGryGTkXbkqIbDqKM6RGkMxNL0KcMufi29O7oSzyVqNucjMKK
2Hc+xj+IAPma6wTr2DKqU8OWYSSOCZXU28yYQzokdxgclbE4pLIvibSQk3V/fo9/kJfunKF45Ifu
9uUkLEFWhmWuDj/r7C0nyPWrER+/tUyzbObZL4j/Ivt73fRWKOARH5hxKDlPDRSn0ESsDUOPpZEz
9NEyQLNEJFoNPKFw387Z1nul3+ERNvOAxTx0IGh0058koZJHXpS/Rfu4O3WhNaXkABrUjMHQoSxp
mg6iEm3zOPMwy4xyAuw8Xtjy5+odbG4O+vme8X1t56TGfVfvEhOyLCpuDoDszedBw3M83LsJeevJ
+BNq1bAFMDtDKeDOTjlcbYzYqU97lVUzYs+tjdNS/UlA/gOWCvk29O94k8N61yhOR+NtIxI8x/yv
WxplZtcAJKzm2zKX2uS1fEKxXqs60ZKhY5alXqkAVqcqtpBzTu/KFP3B+fxMkQZ7Feq/IcD5WTIG
62e/ya4ufIB4KN51360Q2d0UedY6Yw1Wn4zaxfW4zesYuq2/M9SgGGaxXRcZjTT9D5vBUQOqeXZb
J6LmbwGVk/eo9Qw3aY+whyv+NLiUNx+wvQWFieUpJ2ILfktVVh+yW194R2bJhSSf3Lr82CzOVRVg
9L6Y5O0Ut89Vp9iKF/jlopfbfr5y+ORAyT6ZbRnd8yOr5U50Wa84oNudHi01eQwsoFBS1EPe034t
o1mBuoEpvkd7V4JLJRaeji4eYvGMy89MPNpe4VK4/nCVnaImjKENPCW1IAmuSqAyDtWzGtMDdl56
GqQbUF4wau4gHGHKwYsYldT0TVgJVd3l4HuMQ/Z/LNgiKgBD3TNDLgj4OGmiAu1uR/e7Xx4bQYx7
s2QhY7JB5C5hubv81bYy/GzBXcIMyWVP5mW2BWRrR8oFQQ75l14cI7e6vJpxflpgflcpKswzrHOk
4Ysh2qe+5BIY0fGcQIyLXCb3BeofIevSX/kgeaBgw2oGpn3J/1QpL7aZR4dmi259auxxVr9gudU6
9ZhHwSeSuHlUU6DgmxxOPgEc3y3pjYpj9uW5NwTpKLCEtvl+ZwdvY4wGAuvfFISVgHg3l+4XnN0U
rfcJShzO7jq5SrEaRt5AQLAMXcuGP4LIYtqjV7kK9l08H9mm08G8WEvC3j9kiGx+43325dzUp0wE
hUX8phwht12JRWKp8eWZItfBF78wxN0Dp6KwG+5bgzFLBDQQ4RlmLYmZyD3bnCMTfLt2boJnRoq0
0kKvToKZgwCU5XGclHhhDp82DgKsZXUtdQUqsZmuGByK38QLFLPt//IW6tx1gddgUGMfZF4dVmo/
eowxHsIxhd5H+/cnUswtvqlabrERc/qrfMG9GDbLCkUn4Cx/Yq1vr6By7g15WKqRMtWraLISlS65
sAyXq9CK+o3ZavELE7SGLNHBoz7fzbSiRAhgtoNF84c/uNXE1ybvunKf2CbRRj2d51j56gnUHV1W
DbeifqtXtVw1qSv4g+wn0X7jo/IsTBtYtSphyjhgJr+iWDdcytBpY6Aq81nDeOzyt0COsgnE1XZ6
NtUml/Oae9YZF+9WCuNVpcqw3wW9DV+XwCEVhgbJK7X81nCTd/SYyPk9cr4BGlHsYl8J2JXEIB5T
5KYU+7rS2iIiFSxj+fd7Ou3U+bnY5tY/e2vCfGwujprr8Z9qOjGy5xkXDs1XfFuUdEL5FOVPVSrd
dQqZJLTVZikmowINgYlLJP0/UWSuVnrvyQ7iwW1wbjImatODKWbs2bJ2UARyd7gC7sSVXOoDLuyI
6UTvyS/yMvV2vxHU4hZPb+Hf1hTGPJlBucydJxCRfgPMZKA3/8odly1k0gRYi2+W5/BndjFcK9g9
c1LeRYwjVt/NvS5VGOlL+Mnwb4ROCTDuSstUcbuvAXxCTXQdhMKI1CHNkl/OBCWFCkKxhn+cu5tN
akW4RSDOYcD5dh726QuvdEewAy2GfQKdpRcVei7YdDpYP9plSv6DTp9QliAV1bB0UNmyVEMazLXH
EMl5/032JZciS4X3+vwZaZ0qL8h9hQURz6Gmcw1z74lg+yQ8JTJnwBzgvzCo8oH1neA6MdziRR/g
btrmL0nb4mxcjzDou44UGdyjgR3KufEakAR8JT3ML1kA5ByzCjn+uyWUQdJkTt+6XCVJz8QOTgA5
xEddI80M7k5XZGVewn6HNqMltrnF3837UF2xP0bjstVIGovWWdVxXrkSF/m2Z5HMHNaPqSXiJAE/
Iy+EA3TGd7PKueNMnrMVLsi9Q8oRco5X4okD8lUOLko9UphgiTs1qgztfRBaCdsrBFCe1q0TvWoW
6qrWuaFNJmsEyFV5wSGm5p0SZfrK2kqWj0SsIXU48XUnGKPB8WZRXmo5GxAr+VJIFPvfWiG1j6vz
/jnh/Q3ghWPhRJC1edaUTPWmq+SCkGzhGnRFQ5ek8woJV8+PVFL4mgbAiNnQkX2mHwzGH6c6kBP+
cYqhJBO620Zs+mI6DCeqqmSrjBYzGma4+Pc0OQ5WbWILx807fwpTL42iGOgfUWd1qsPNKGuOcQgC
lY167rhrjvJph/mNS7v88bmL0D+V91Gx4ZOKtmR9t2x2NRLGpqu/YJxhXdbClaKoVgGO/7LVMSgr
eU8XHjNsiAKWGxGwI74Po4xTSjTvQBgUnGWJhaHq2oWvMj7Oanz0KSd9un+bRSR+MFwSo3nB3XIj
7iui/4vfJz1xTPDYsusFV2nPiHsuU7Ap1WjbDW5ZzM7KeCxm6+LS4ICwsF6MkciNvTJP0BYceJhb
nTbPdnVwEUPx+3WilTGPUVZgKcZEvZO1oQNIysYrlmIzTCMGrefhbd5+/ZRnnTpkExss45lWnCnX
QQDRO+S3zBl+7MDjBkSX1+ZodskO99zoVxcSmGS6CWF8ob7GG5vf47yDgK4e0xx1eOhbpvKC+5Hh
cIfgLE5S8C4ee7UEspBaeV5GUIfeVlF51atNUYAFe7lTq4YoMf2yWR2+oACBYo0CIZAAiJG0rjh0
GJ0lRwU42EAxle5wvHX8xaqe9H/60SMwBad6BieaNYt3BWjOLGhQCgKltyHCh8LtIKHrjpmM9B4j
wbEWSRDBmmEZep07lM/4yLZqoieSB+HdQ9LBV/suwrcN5lvp3f9H0drkTXomWkob5ou6IEWc4s+T
Tp4698O30HCzYRJNCi7K9wTPTzqORlLl4H2mi/xe/quPDB0yxFYdM+08+vuf42kJdQzQsp5+Fet4
uFc8BzLyvdt9Fc1lDtq93LYDTAzjVIt+qjFclOt11mScZvdl59oOqlP0AEcHgA6sh8Jpvl3LL7pN
Z1IFLLYnvfAXCabP7+k8c5kOuSL+lSRtD1pMxjQkQuLSx6ZxB+2NEIZjb3Xqr8zdvuIbV3X4xuIv
P4xOaT2oqQ5tkxDD9L9S4U4DQeuLEfQruYKjlaaVo6dA0nCbZYkQsZPEqa5b1oGPYz1CadZMV2I0
vd8H6woZ8dPRY3OPYKl/WpjkG0uxgqAkMa0BYcWbbliclN6Wx0lpeZBZAPcNU9UZ5FrEtrq5SstC
qg+P0QYtnn4YBxaFe050RsEPXf/8e31L9raD6Ee1zsbKAjMj4c3w/lwqUvHIQsVwhVN/8dGOPUQ8
WsGYMeW0Bmi9jECWvmwPo3CeLVQmKVLaF4+x3+Q06s/AXDxjzipKEyJ6DYOi+YjU+cL8KuyO5usC
bTgx+vLQSlK0oDQDRElI1vdqQOdHlzhNaw5QqkIqq4R9KhXioezK7/uyT70dKU8wsTD9w+Yfde9X
VHfXNhR8xtnZmp9QBCBqbOLTkaTN469U9KrkHn2MJ+OV7HMNdqekOKEpYqkTgj8M8RAIzHaJJg85
HkCSy0K1YTvg0QAbNdQ309Gn1AIvYC/poUYR5+12H1cUYS16kWtbTi81WP5vmpzr1p9jCBx81FQR
33GoYIlB+7nElgW5FMd4eXzdP0T6lHM1gSIi6cZR3fCcxIQABXOADMWeuSz1asEV+d8jk0Ii3GTW
Yp8SUcG1eCtsxbtChCzNkIgwEoS9Zrg7yQRgeEOCjlBn5MZtjJwBgW2j/B1UJiBZyDtWtt/hZoh2
su+T264aA6eM1blUbhNTY/aNKqh3gF+rT+030UxhoFWC5zKocfBUpw2T+Q4O4A8S2Hjh8sC2h/rq
Hd1vTUsj8S+d6no39PqhHJveeSXJIWrSf2Y5BOiILpfHrVRLBjScqpEaEHBk8mKLr5WuUDYhh6uE
JsZJhMmKGX8//H4lTsqEKvCbDPWlRbOkkAKoeNshFlYynzh0vGVbVymcRQ2Bf9NdswPUtsWcGQBT
h5Av9mAZHKfFYUEZIj23KTj/h2vdTgsIbpY08P5+3Wt5F8qijKjmXIEDaPHxoEf156dR1BLINIOe
EH6ZySyhP30xSO+2oWgu9Wp96MxBFdngP3HA6+5iMWE+YtvODBNLLz+3UiyHqUti8DxyHdhaEG+A
vx1fMOQc6q1+Axn9NH177VuQazhOLr0JZ8gw5fdAixc2Y7SbJ4C++u0ygpGTZbLlunRFRicTgoqy
qjNEBr9bFDSBZtRRmhArtX4MOoBMRdRKQMCtcd+F9Rkt+iGS9PGRX9kNMFOjXvifgqMxmqnwVBpS
JF73e+/SdB5NPUJdof9IwVe9Hg/Arn+XzpD8ajX0NwKpSlM1Qo5zKvANLZufPLnOd+jF44fOTUKg
ka+p1lRh8/t4AiX4F4E09lBSk2ufKUbPkDuYbfKFeVLqrC6AK7luU+ujXAIf2ZaBdPBfhkAg6sCg
X971HQaJrfMUoTp0vnYl5qXksTRJ4hEoULC/yRMXKO9dC2WuTGd2uK11a4hRvv8hqmD2s5DEVYRN
uWBu0z5EqwUmiSemQkiO+1otr67qBWDyeQJiPLI/fBzOdws9mZXn6fplX+HgAGo8IPlNcqxye8qT
Oqr6IqlruZKt6caHQE3d1DnL6wT8Q5da6bJarj9LADwBIbYNeToQLle46PvS49Eo8S6iwg4xHiN7
yiDTdMotdmxyWUaryQYFyqqcm8/clb3WWZcITMmSg+MJkpweQhotoBr0sbphsxhFB4XAPlx24Ifl
82U+f2RNfyTKWpX/Kwbw5MsvlfH9MPA6qve8HmFsQnR+kkhzS7RVaZHwrebekmMGOnqI/YcFXHjs
dE1DEmzlZRgxJE1Q4uEj0bIAkFSxY28J2f4cJk3+6x7IyInkYNtn5sKs9KUOha/+3ulDYE9JUUqs
9OuTN1FvlhzuA+iNMQb6NEylehuWtn6i0+NQq6HcoVrVf9EY1Jvbb/J55Y6AY+Mv0gXBDR1JFnBG
lI+pZLukcb245apFoVDcW0yxoGGJulSuFJE7rbD/wxOkONfaGVCcCsFdHMkR+EoQALskCWJcOV+U
Up6OIwAfmnbyyMUpus3aKpvFAudoXxYiYdhIr/6NnYbU1VgfoAphDOko8ULon2xmOOMl59ugcaOV
jIRfQOp+bx6q/1JvaqpsALBWmchDDN0fElrVlxtRePSwGXjYVCEykhV+XZ+Gt3SCziGMblzYPR/L
oCp9I3p15qtxLc5MXFC9/Ae5fo+h3oN2lw/DAsfnrSfVu42RGJGDklqCUApx0lKWe4C7KryjRutb
HU/zwG+S4XtyEb6FLN4oUmNZekohYfrBq8sYdKTtNzvjubovgHYGLOhZXnlEZwedb+AflK489o7k
XAUk74cauoToWuYkH9jtTZy+hSMcqjFBYjLtYDCflVdGh4YSCxqbSpfnvuuKKYKaJtZUc14lVGqt
+KALgXWuVGsQO6DA5mRiKtq+f/4vYUccSilcrADsD6KIfpCaX9pmcA4R6Rm3HtExguvDMnSpSR9q
VI/71jk5T+bbQbhL5R+sUSE8BByYmGFLEFadeMHV2Tdq/vBD2giKlcJlK+R9VLHmiq8FYbgtxkTO
qi6aoteGwUoLOFfeAaO84hNGr6AQzE5Q/X+KM7dgUuCxHHTbf7onnp6gCMJ1I1TgxA8+utwIwZJ0
wV0nmZ9ut2BWtWvN8Y4Fr1drfopocCZ63NK3XM3J/3ByzzIf+bn1tTkFHlCe3bLRci/gvvPLUskT
c2qAdSlMAAH1oQpEyw2Dt1Xf5bdd3T8SXRgUOqaZXUUT+UD9VCCwEvoTFmhJj46rzd25JxHIF9d8
VhBGmtxmFQsLUtuvaP1WAg7fQ5zrMLqO7/Iup3UvNujrqhlFVs8/WBUyMbjpRG4tA7Rb+rECUpHK
8YSEuw3qaln7kXR0aYf/dYVsSCdiXpiPjYBtRSjRv0KWgMxJr9UwCv7TNNJR35BVfai2mXi0jV9J
oUMAcGFOpy5qnCTRYhp7Z0dxQVqQMwllDBHrirNH+vjxsZACvbWfLEPreWSsnodceoXaa7yCfbOi
9DhBrVgdyfecwYFGST+KZfzeegnuhQ/QaEipvDjBD3uPxTa+PJrfh+yQeWKWIkURz7/lq3ruY+eH
RSGB2bVZOdT+3Ml9Cc7fdnuNcuQU03zcLl6OBNpR6pl1YrvtOVXt2uQl6nD8fcEMRLHZ4XaeKI7r
9TWGVyyk/MvM/6j+RFXDQz6rxJCN91vVV+FZhamuRTbkrVno0fpZkqYTERuwpYHDtyfgnClgnQIT
3DXtP8R57hJVpE70A4w7786D9hyaUUyeZT8NAm212riB9ry7IX3BIoePlb1hXWkyBunto0VCpdoX
6CnyeIzDz3m7r+3GL1np8r/l8dQZXtUp9O9ikkYpDzFb4I9Fl+C6fv0C9HIEhUZI1L3WRVV+3kIW
twGJI+QAMh1XWfNfdc+IK8jduL/FKNf0tcntfbU+UQiXx1SWxpbkn3XkIFYY/AYwQrhfqPQN0yzP
2sWXytbMacs3+MI39onrOI+GaezJ6NZqqvsbeY9zLHM2UcwhMspxCSUdOEyFtfzninbNCJIaVaYT
at3TJZtu1If2RGsPMtAL+GDmUwcVyivxwb6NFrKJqtuTKvpe+pY2+E6cfUMJ+rPFW4hl5DfAa5JA
XKSJfESKz13JQwLj7aeV3cI1jIIMBkV0gVK2tgjRjcoZDmNw5cLIExeDNgANUDAluaVeQq+FCzNf
YeqMNHtMQRQT/nz8u0br5Swq2CnYwQNF3a0GALW3Oyga9qOuke+QRcdSS1vo5kMTjjGDauSua+np
86reFM3/InfJK3s3N3KenhACbR1YiJOKYd2LcWPL1ftZQJwl4Bl4KnSfMr8Biw6BYWmicw+kKbtG
0YsPhOF4bRN7Kmzq1EXy1wendruyi+m5Sze8pCslAGdtEkt+VO6kLwGCGSI4SJAKd7IGoNmiiYyA
OFlLH2D7cau1hBBplGhrYp1JlcMWW3lxBNHxsrs4Jd0nfOlhflEu4gr5i2Fze3MVehqqyHuulVVV
ODHDDTHaRPP+1eM6oUgW8ysHFoNAaNUlbjPzM47pRUKDAPWOKhzuwSZAJsQWavh/BlTY5Efo+G6k
TagaPmL1TwIQYFUT7How0adDaYNbV6/4SkbhbI1GBDMFHoIHb4bX6/J/RW7DRVgjWpmo0lEWm9IV
7zaADyuXLKB0aSdTX066oK/BMZ7hN9SANc9Bf2pRyDwqNh8zvlHCUQ8RUnFwn/ohoFgXuZFj6XAO
Xia2EMjrDXI13N6P8ZYHocd6800969tLy27gFhx3DZKsa4u5t+vl3MGlILy1fveHngRqa0KUj1y5
raxBP1YxaoaAyUNgl6Esl3PcFuFNUL5Yg3poSKKzXV4BwfMHJf4OesWnP5sGqwS14ecnb+Ij7g79
Mmr6mr+1+lYp2KDb2LXSMfB9ztSGavcciawmKwci1ezzNkPFYgn2XliQkdm54xSw/lYfhleUN6VW
3mFVHAlTEjlX6CU6Sa4EQfgVor0FeGEH5p2sWfLgh9871GokraYa5brZJ8f8i+BzW5hOte2Ve0mI
oQ0/RPZ3D6EE4Gw9Xefj+ly5MfW/EgtsQd0+I5EyKa/jTDT1P6oLiV+gLDrXMedmylk1LLq+uwr3
fu3zRt0TKP1oG4gDbXl24WY2OhmvuQlLCeKPkUZuI7wWjaPUrNFsnEYZoI6uKzBMmmbz6iMrKdY3
M6jNWc8GCfgQcq2pzvaZhQSHvvuu86JewQoOLDOFXIozPShhN1GrjDxgPdzpmNsuYUttx6JjhaMf
vTD6pX9ia8KKncDVcnwM9rYzcav+uJZ3d8gIcTPH8qcHaQFCTOFX/HiPiQhbpu/lixaaOBTtFc4N
HAiJHZO8FggAdV5jJfMZKIC4mKJC99QVlpFgOVrazqVwY72WO2mWOQk1LF4NYFnszngejWyGD2mc
/kUBNYVRZLsQQQLAMx64oiz+T0NZ9tu3bWgT60Dp9szhiLO34eCGZZ/aCnOxj10Kv+rRuCt5QGdC
ceFBZFx+D3C4+FBR7uNf7C8ya/0ArphgqcN/g8ihu3OAHu9kkyj308UI4PWxZ/YNXOpMuVgNVx/O
N6U9MYSY5HQsuJ6g0Frn/NRE9nrcWKi9TWIz9KxZAERVLzifn/fZEL2ORwlhY3K9n0oR7//cv29K
GroOuqf/3QNWeF1T0Vg81z4EAIW8j+9fr7UxcCAOQscyJEsWGPshU5o2u4y4IBc0MBBp6+wSzKGr
GcCAGGGpy8tyVOvjgpnkXO4TXytsFP/tmbZIaG47A2H1hyo5J2Wr/uJo6j4N/HVe2x1xQbW54am6
7QlI4GTNamrKpIGy2pLmchSvgXXMxk+isnmu58EYiewkDyGDJElrE00eIHHvdyyi/28NHk6JQjgD
lG28Y3nM6R8Fuh4TqZVjRG68FvdqeamNak8Q5E9PXHTENpFKGwg4zP3hyKRONjx0Ejy9bD+ulUOn
Zlp5MpqH+m6wam2ybfPDxIFPnIbMr6cBWniUqzI345TJvW5l8Eg40dwGAa+Di03M+Nb56Gj1vqpT
fMFWsPSc+IJ35BKB1uNrkDBeORRbDlsBQ3CrU1LhWblcquhM/kaBoYjvxozcmRgJDUxTI3XiQPMy
BsZiaD7XZFbwGcSe79MLVnGfqxtEpH3Ggps4RDBWXbjeviuvs8hnoQnD5TGhVXS0t79nsPgdSfQF
Dhir3efSHv64wI7G/rpz3Ofo1qUFRm8EQOaLgxN4YKmUiQc7vlZUI5JUQOUaxjPeMOsXwkHFfrdi
yUZzYvhbt7ymefRJ8OduXazglVxb7Mis3nWEpTOONjvhGSYvzlqlc9yeVhCCBlVP7XupIsB8fYhY
/fI58+Q2bVREMvqxn2w3Xqfi5w52r75wgzH3/UXdzVyNa7NtMhbDNEKT7upXXHauhXvS1WEK1d8z
t6mWrvjfgkAYgR2G5SxT72YNQ5LaJctRFZbBK06/bc9XhBhyZjmfj6LfnyFUwTK+Ncp9EBSw36vd
m3ZCyLb/GoZtbmCQ9mE9kcp3fRd/3w6d2mSVgh1U1m5q8lnPZzTFA3niU3qfoxVQ9qmSpL6rVl4C
n1tF8uBkftb+wktgOV57KSURsBmhudcGG7CEZ3LbJjBiJ5lQqpvft7NrePfV2UaaoVAyoszxKR6a
zqZPCdmsbe0FBugeSBE1X9V/YCqLwsfiErkZvSLLyy6OPQJkfVxXSDsNQIDadLtCblSJS3FLom9p
pTrWNGT9aOBcMq+g6Eha3GAoWShxfXgKxmiQheIC3AbNqk+ZTs8OExEiakY3ruQKYfQi36ePXShm
3VD2psX1/0lFAPRpubCyFdWJBm24s11zr7PysCwcH4ivfhkmIOpnI3CqdsxYnxI5mrvfTEd3lWA4
L8fWT9tQa3yvR3JGIIG++Eijqq7cbtr1jBYl4LEyDroLa6kpEYmjYJ4xuDKoF0woOpSL+ebye+W7
+Sv2rUZoLsSD7OeY73OJhjwzv+/OK9QRP1q0+9SvanA3Sv0rzSkbFIgXjXd1WmjsPKZ/h1qrE9f6
+r4WW6w/12+JCq8B2XrAOD33+L2uiV9WPS0K88D9znt40hcy1fzo6S/yGof99FJdSH7aIy0Z5cth
70kMDrCgZGeFseRCaFwguh6NGrsjKCgOvzP+ayVCLnWu8uyFseZWymZA6Akn3p4F6vu6I5BZhEIw
pc2x4NkxwBa85vT5voooA4AWDatULwQL12usyY9bEvbnSckBntslxVF/Ziy4F4znZQUtauZNe6g8
xM0VchUBbgkacsRFzt63cBSAMmfnIw8Zq1m6Z7RdCLBEF+a/tQwuZsPsAgvVeP89NBbjdiDHgTYR
IyAwhktTP4GvpnQ8XJ7V0PZ6mWdreB02VCbwBn1TvvMq2v2XnacyQPuQsWQzRaypmR9PSYv6TBLq
n1iqNeRmLt9NNxfwpmzzuJe8lWUB5XOWZTrHbqLlHTZIn1XTbW2A1mp7gLiR/aHOe70+QZ+qdInF
1PrPC2jgLT0KsKwL9MJxuFLKFISBn72pwevPXpp+wf3HJCZ90Zqojjgg4fzajzCQMymyKazmkh3+
jHn3CaDTDRrxaQM3iRIYJ/jfvSHPx0JVI0PTaWQ1DcreMEjw4Qz4kyIn/wagHY/GUvDcD+ivqWn6
cD1JzzerFW3b9UHD1dXkhPUzrYTajyRefDvsW0W7qyEN42loOTPkQ663ijOFyQURy2QmAonpLlT1
Xn/qHpShC37UTZIrmB3Pn5RWXk4M5LYiMdqVxnRS3Z9/RHCybsqEfBhJoi2B9IIMtoS2rx5CciGZ
1efY3lYLjg42cwJj1UbGZvzBO0MvM53wRcqfdvpTX3seLQVXwjeM2VisZy2VI6Mn6wqBFXo771Ts
Ruh7giEb0p4YJGvgLxDJ8IRUzdZhJAzyDZuxzd7jhHcG/XqMVTeUrxgpmYS9sGwpFa0HVd8OFUy/
rH4FB0gGwWcCXr/QQaETFVQz5bznG4cAhOUmuz/4fibmww7MbwpDOXDjMRmMrBCjqeDtpezlZqp9
E7qY2zak1xr8/Kpkk3sUhS5karwy7JoB/5kMbBMXjOIXR43AqMRXt2kblxf2mwJVE81Jy6DyUtB/
1Yh9rNYugBfQt6T5eCen12BzdLOc2c5ctNEpAIh+mwvs3TMLq9j2YBWX8SVGi20VYRhm7p4ZaXB7
fyGwk9+WRj9ZbxBmufxXxn+D66a7IMJ1mFxCgeuugOEkZ55QvsruflySPyjhfBsxi6ONuRJ+s7gm
O8z2Hr2En3PpBaeLbSmAFXhl3b98ix5xgKvDtH4eryO7AshKwnV/+Z439R2MTRQ/xUG5v0dGW6GL
jiEw3vzJlyjQipJAAS28/DTWPrtqfOU3AnIt+mJsyF9Mpu7dZ8dIgg8fsoyP2h+GolhOxVxY7SXj
loCREzaZlzxfNxyEVwH8h1yHNrtwHMZYuVR5AUvgHZbOjfGbkylkjI2IrSa9Vvlx0v+fdVPNtJii
zfG7wzF1QwjGMmu40Q2Na6ulVl7RvGTXniOYEo9uBSz+fc3VWffGnCzaDhdvLs8ydfSOnm9bL/fz
NokRQ031SmbXGFHkCFMODmhRAOlVxeloDL1Gkt7vJ64kbtXIkwhyXXkIvBqlSJli+g9oCzjOqjkT
bD1kI7u5Xk0vEfRaICgyXicBVim0ZowpY1LlAgjEwIqZc+4gm54g0IZnlE8JlYGMKONHCZpBJQI3
txg4Sfh2mBxuvhilmemlyrZgGZDU7VnsZXAX/5eACZcEX+NRJ8faDwT8mzdj1Hto4iVRsm7z4mpE
e6ivuAafnRewn0It0tC/ZnImOLkdDvWoZeUGV36C0BHGsTdn4prxrkPuTLACRpYFKou9ckOQbKY3
1RHg912lOtgWTWE8pvxOSbJRru5j2gMvq+i7gW2Ioxp7Y/WXFE0hgdQQ3xybkJU6LBNlZESJs0kD
EGfqUQXkPJqMgFoTxXitrMbFUMpSnY21oWGEGIx8QClTPiA1BEvVCEmj7h5aqhLgkBpV1fhwJ/QM
qJtw9tmg4nLGa6b/C6FfEGDlX5jDAUGUfFc26SFvl+HL6jQBimARmy51LlL9URMmYRD8dhUJdiuY
1CUR8DhgKKTUlts2nkhmxkdWfQliyMHdemAOaeGrhKtn31RvwtNNxJ9ScFxSCON/Vke6QKpz19IL
e4NHrIUJIOePgklb5fP3votjo6b4uZJxa9KnMHdR22/f2ts+ST9/AHxXH7Y89fJZ35ahumHpLnp4
8KUfwYdm7MU81EuO2JOfO6U2CZ10hsW1La6amXdaQLhuZ9Jujjc6Dg6Akc+68lbJfF1M+6q6V3QA
2xx3vrtVQBBPVwezNARzSg2wJafQT/z9CO3i4/0PGMxoNTPGQKixttjmvL21riOaCREaOgHWG+XU
IacVf56L7sTki5Gc4bEUHUsTuxoQ3dofmC4cdcYWMd1k1eYJeAvLksSkYRXjeP31uBO7JheJqecV
scBW0cX1nBA/uruACYmI4DSxOxqdYkn5Dn2wQNYfYeu/4dJfjywu/8aowrDKQpS+pZUUrPxyu/Vo
z02q7oe5UOlBJh8LCS4hMsgXgthMi1pecQv+tui405izVtL0sqPmC4/oHVVPHqPeBMHeDaIfiW2O
drWTWYtTg4EZeoSazx1pe6GILmFlR4g+UqPfnj1VZWnkl6Io5xjd2Kn3np6mYfVX/DfV/PqI3fMm
Zk18+wS/xcat8wkyDw1aWE1O6aGDWMVpJUQk57p5Qd9tCooRctuVf52N8YAE6LGwpLFM7kDHW3Qx
z+3bi0kXGw1PtTQMvsXCInw/QvsQEeNgYyqfEz265m8saO/1dOsLxJRHS9NDXiXxO1eV8cLyj3lk
oCm49yCiYaPpf8iJljRnBOPOmprgZq47HVVRoQXCe7NRjR7YZj2asIbHTU00aRccdM/ZL/yIuT4v
7J1mb24A6TixvKLD5eViCB+fIZjdJugCsdtHF3uAl1/bpgMzyKluKaug3A8q8wQvUzuCi/PhhYhu
xVHknPAwwF6K4TZs9ux0Ysig7XSCy9g/yZJDERr5pUIdIsYQAJAkxnCGfZJSZDqgys0Cpp4n0nTC
ECFmGsYEoJzKLBkuMQMGa8hVE/NNXr2ZVjuuTCtW8vloltzrNfR3DbA7HMM6MLFXw/LUtj6InAtn
0eCNaBhtXFvSGXpOKTLv5WIkOQJjbG8sWzjaOoJ71F+0cssfYZOM/KvndQi06swokneYj2wrtF8a
i6/7JFfZUBwh+KHIBOZ8+PZw/asl2v7QOl428UKc0cEByF6hZd/uMFluqR6dQTZnq+XXAQP0HCOb
1TWWXnk77VYN/zd/Ap9pvuf4d+q6Otg+kaxfNBhI/sdaIw7cyCoJZFkxqTNwzIXCLLxOzKnLUP4G
Znb2FRnwe3JkFQjbF1Sq6/Qr2OKuXFAZPcAVS3u4bXhkM+dUeQYxOrXYEZXKQI3j+42ziGosqqGX
FTIcQ0SygLqEGcXWABhcnF3VxLLJDslpdGTfEGv1cwiGWMqhEVR7UUe+8PNExUgWOWwmsOcCfnNZ
CXUbfYmoGAYH0Rj14IJ0orezUZYxeo6KQzovvkByWxpx/AKGRWSQl8ps3NPtSqU9pJp7q6tfueHp
8K0fOTBermYw3dfeVSVr3ODYTk2lCUUlS+GEQJmcqDfmTiFwr63sFCFfl1DMckaozNUp8rKcB3P+
MlSAr2ZjVTzDVUk/MiAALY0qrWcPfmv9+EdUxR44c5qu+YMqWDyjdwKHeBG1l1GfPYfkFaiPRnFV
Ahw5Gz+WMcqIp0qnDko+/GGq3kZZbrP7aQZ3kQIc9lSC0vu/6mb4o338i4quShXcTu48hicdn6E5
soARQUKedGRgyxS7I9rrCTbmL+twU7+DE6wvaZxw+LQX/AoILqs3ELG7CAOAvTuBzbI6EQoh1AuN
Rmd/oQP2WpdrF0xSqHngg1cnuZ2KydsJfa8sQOXV8sQcdLxoBTB2PjMD03yB+qpLjtQ5WLxbW0jr
WErZqKSU/LBs/63ba1hT4xttLjsSRPHy4lqYamoPTApKBBBY0ztphV1dU90eOk4oDFy/XRefQpV5
2ASm8GHs4ZriixvpQWVbQBBQVU2ILeaHv59uWhJgoj/9m4WXM8Op334k+kbdiGqLxNyHuIm2x7Qo
uuUpx+b+HL6gMr4v39Avrkl7pLaXlJd/Q8kGZfbBvyhWpfODzW70QFrOcTFH8KeTJ2LvbLIuwOS2
MlONGpjIJThTIImdHcITQMXF4m2s0lU/XOLOezZDNLap4Ys++yGNRvxGe5MkS1gaoNQE2JpQThx5
/LQhHq1TX6EYMKes0tZB31a5Bx3INZYYa0BarSY9pINERyW4xMN0xs7z8kAy64/B/srgmN3nP344
r4IQcJMfPReDdLPns404l7WB+Qy89h5g96q77HUrnQPdgMEqpaQGRocPJRnyXrLYGM//ZIORA7Da
hnmH0WS/sUEb2dIZ9nrmGoZWKXUXVNjaiboCXiz46nObsc85/8EjDAJiRnOARRWb94dPJrHRCMAG
j+Dk7BdQcLTPSSZ+BNa+vyYR8aplpiL1SNOHBEqWFJZ0svZVHuPP/Wm8y8SNZCiU177F100N413Y
STzkWGntjMeHokgDmzS9IX3PLNeFdq8H8vvmyuV2qKIze38eRNpt0AjP5FpPpb9i/A+QqTGTPm8X
s9YyOPFYbx4l80byuXoSLMtg/CzU11JfvJC16G6qo2f4z0hEBqxPmNqMerhVa2UJCUEv92lGY3yn
8FyAnGIWMKLAQKkstigl/A+dpoegQVxn20n9v1U9v/GWaJ1lBd/MN+RCu2OG9woT88JOJe1fZNcD
gvBycYcr02Um17dAvrSFYF1Xqj0ZAtB/uS1A+wTpme8AFXSEkc6BVWpYSKYW3plvlHwSZEb8tAyz
GTLGyBKoIUfomNbj8KvAPHUTVrmx7gPVrFQRE9EDXfSf5AX4ThO29GluqRm7GqURC8ddYtQ7WMLx
56B40QwFOwu4UKPRdHa3hsQthaufNg0GH7x7dDNP1GsszxhpjigGp18KaNKkRJUS3+mcVHXKQYqR
1tGAYktcAFAGlfnOHeqEgCesi/7ZV4h/jfUCIWFBb6IRNtOd1g1RyQBntnBxHFsMADa3usiVMXUF
6b+gCo6BdWxezRJh/FI9fxnMvyO0ZEhkDplqHAPqPLHW/FgFpfSq5r5+SXIt6mMtlVpfwM2luWZ4
vcJDXx9M5gyNaCaCFHBZHFhSH8XBEiUs5RR1qeg7olonifnoTpxeP4Pdacl3YySNpQDpg3O2of6T
q4DyHLCZNNR78ooe3cWGe9wIX3PCdTjBSCis3tkxwDl1DttIZP5byldVwEhZxsS+8er2XVsMqt9l
LlmV+eyES3weAhCvxY3gdrUU1i0qn6I1hdbVT9d2gGxXkU9w9JNV8V9dtU2Gh56WQczA3XhTC7YG
MSDo6TiomQChD5iRwItDC+fzxPsTjdwmT1B5+ZqRHdPtO3sg4jHzse1ercG4JzqD5mbXW6hqZcdR
F019Q+WE0PgNSX+EHbXH4VKrS66vPqfBMfZ4tMcdSvPF6BxmZ8vYB/1NXFzZdhMZI97F0y4kp3yJ
BMyLysbLAIZcKIXGo30Pmo9RvN3ghw+JavrhgKHprvvDEDzTyP0rKH1ItlvNfkmTdlJIsjFJpL/h
k0Xa1R3DfIuz4qsfcohQ3xPG1WSZ4lTJslrt8Y0aG6pe5GgpRfTolnYF3BZtroZMRAuh4GWiKgot
bGMnLrrAbK0WvOMEPW6b0EWpxSHFfA0B+R5p6Ei/YGklLbj112QO5ogUR20QRNPLk7rgj5xSo6lk
txFn5bys/23dMO/Uo/htRRMiHEUUsB7SSwBaTeC/uTAzbE4YASnqQkfd26TTx9Yh9I4aMo+RLTd9
uoJl+18huPhhE1JRuYJ/10Y+RbOE+f5g77y5bQZcuLBuTHs0Yt/I9PKCHXsPmV8pGYvUY2F+fmca
uxKPttKBtITFhnNw9w2dKtOKpkaxUGta+EVCQsQYy+EvXVRekjtseCuTAm+RVTPb1oRz1ILrW2WV
fiupMXgjGXl4mx5mCSFKRvg4Dcj6xb6/j+4XzXlhAYdCmOInCfMiiliZ7UEBRSY33dJ4q05L9PFo
zNNWvOY7igsp3bBmYMFGtWdc028A2Al2saeo3g6rK79f+ZH3u0/S3ZX3s9t84H6ghrHytVdXwb7a
1lCPIx9cS26gb8A0gjhmGd0PtLeGgpdpkzqD6dWN6/dgexGobE8zTF4GnxFrLDZlewQvoK06qP0G
1cjfTn9BKmm+YGzaGiwcDNB+FHr9ZbUV73pdLd5y7Sw8TEY4vIQE1N68tgXQnms5P/hm+4qkfoZQ
Su0t3l0+wWcSXJMwJMvRuz00/AKtOf44flNYZA8QzzLx1QEM/6OJaYFh9OLlUXuWNq1pmgOaSpIy
0aHUAf+zDf2FiGksjm8V5U7uNOfjs8NL+znWMDth3Wmp/En0+49gvXDkd8ormgnNksRN/lFD3ULJ
L/K2akPl9UfJ6XGrvc/VsImFsb0WQxf0jdjqa58JHVMV6NDVSpHNweTSb1C546uSKdIP/r/+7eyP
t3P54XIdDa5KX2tJqtzTbJKaamWr31cuSpm0txfzXPyJ8lvSUUucBJdFGiOhcP+f4cA1S3tGBh8o
3g5AiMVcq4M/awrm/csywwJv7K3Bn9aGaXNeQZyQHqNM+v5SPkVJctsQLnPuewicviMmacEurS/G
jOaJ08gmWsghiIt9pCUvS3gqGFm+ofKqiChi/3odn7rLyrk0AiRat6tdhZEtdDQXYSwnilfPRdmn
P2Vn87fFGr+sUfXSbtkB+rw7obmY9KTL57b/OO272Smzicr7uzh6czzu5JEOMjP+h+h1voljXyQx
mSoCKgb/af+87hyWhTnWPPqSKwHD0BlHTML/bWIGEG5sVN5cnTahMnzPFRPyV4bwg4ZbBr0U1Zr5
5gzvIzet+0HN5K7kTqP+ap7Y137g+anoM7fMr3Op6g25BRk3JcpWCpLhzCC5+5FHrNyFAwKTQBIy
lCRA50JPqpHGWupZcR938eOCgSSmQqg9ZgscAlCT7GFfyVWnvpUcAZqAanC9+HbPKxLK6smAe03c
5p0PEQX+Xd+0JWzW+2iFMzg2QMOooI+0pi20N8JhR3NVbKxS5G0BrfMcGJ18Md+e/m/nuhwaUfbr
Ih3bh8BOU8dJ6HVpVefY5AkOZI9s2yhfBD1l7wUKZRJBQLoXCHFMkJTG2wshCFuzGPa0yrLCImVD
cSJK/QOgI/C4gknY7N3rQ3djTktAT/UVmrx3Onyva8A1ycggJSH2+3oj8h/39MDKtIVEAGqMZeVW
3gNpkfV0rI7X02YvY73EJUQ9zbGgzUDKDE+Aw+27Z7hr3/94WUfcWLtFSvDrzkQilcSua4wP6VG6
CfR2ofTw8bkL8HVeVVp8ZG+/l0htziKTjcj+HcDiuBQM0QCR4aET5dha2FlLWAx3ftUQW7nd9oZG
oLIJrCRcw2IiQbkuSsbP4e8uOjotg6blvsdJOk2wYA5MBo/NpKJep7Wlr24CANuum4Da/1WxUSI0
7v77XSz6mX4LGmnRffEuV+h8i7zAY0DQAYRIDPDICfb2AAz4EFs4+8R4VzE0ZOk5LAgKkDfLS4Jt
3W2r+bYk8ug0+cg2+0i0dBBvdfYe7WOdITl9lRyHhvaPyrSYvfAu9zRDIdtp/QTXaSMdLYkGQaAW
qkm0ODHaJZr9VbqPJqwVgBQygAXQrH4/D8ncz7sJqzJ2l8xPwt1wu4Xp4LBGssJwiBeYm9skpPax
lNVG4jxnTPqVZob7fLaZy9OQAu8vKZdvKIgjLLu8abboa3VoCoWNzxPlSbNGEK/1Bz/Hf/SmHFec
Pzf8TP934YSWnvlChqPLqvqhzHC7+kjcuoSTxBUF5f9EN/k9UynmzMQHLwmr3DFPlev5Tp/iLqfL
UK84ELkmLTRzGt30GFx02n5WNT1k6Df12xFdMta9DCqbIWzcTyp+aesWqLm5lNuosHe+jTPx6bad
4nZEEF2loeUkNfmArVvCOq3+ZtN43Cyi+LtwrU5b+QVhkCuxM08vqUY7g6kMIe2XTucucVR2u3b/
EzedOFjDwBCY8EryA22eqBv34tmoEfMScyNTMkVT0WoVqZQodziU0SpK7ojghEj+AWilaXiAveIG
E3FMQCy+qDHFehFJ4qSpm9ZAGfz0JTGo7Zr19v66u1755G0jcPvUxOlFLUfJkA/VJebkqOblmsrB
+ZAm9j3Nk/n/Yf64Hq9uznu11X347eJmKweWLOw9ymGaahxGNW44yCX0eYuJjZax5m0PAJxRLoft
i/OT8oqWDfOINzibxsQ0L8Kk3x6Od4a8GlYLPH4HP0yYjueXQAZUC6ovnEIKotHnH71r06tCur1f
0Li7ugb7iS8FaF+tS1rdzdE5XabeQowT07dzpF510aFYXguwzMS7M2noWRj73GDOicX4YAT1lkW6
/GxSA6j/norYX+q3Wc02caxulhIKAYcDInZ4ZMaKvPKn+tosJy2Kw6wp/A3O4O4OsgBRqCjJtVh4
3TuySqKPe4QMdG+XqySedfrK0+w9vzkB18VfOPh6HRw6CIO+VNTy4hS9ULnMrO5KCeGOGsnmkxJ/
snyVA0t4b7WdWr4VYVVY5twMuIcilYCzgb/lWTIXqXVu1e48+44zmZCG74huzhbeoITF1vYA6kD1
zJz4kX+/m4swVh1AzDkBYgDiec4drKnU7fOGW5/KZuIUkmeHMc2EAy/Fpm0nuyK5NWGV8cJV+r7k
WdVs1Qs5lKDxZS05NKc9Lh2h9i1fluONeUcSCdxTZ7qUXuQ4mfRyCyCx11nluYCwVbqCuneEgJ4U
YOPX1rQnrz+ofhM5LdA3YhCj3m+p0lAk0NYLjBXb9Z3/puh6DYhTC6Mt1KNtDJck/z5m/bx2Qb4w
bJ0SaSV+D2sjfccFpgmdgXrSVS0HLuO+EPG9XvJomyYonDMf5KHDHwiJF3tTzkII4yTFoXlZebso
YTXxv0Ns6X1pxM6e1tOQLVAzFvpL+6QJYBztIR/Im9qDNcYhKMWWd2jtxboftqJAHosVVveKsvQ2
it5JuRfqZaQxZ39bMWqZtoY8eITKSWvYjMcXl3YL5M4EgLNe435Tg2MOf5Alpw6OZjI51uw/IX0k
096jNnuhch4k1OAM0gv5NbA0v65Sw0luacYZnF4c2ZrMQg9DwjaF1NHLedoOwUF7Cll9ABolG2Fc
xVKbBYymY1zuliJsANwU/zWYaegOaBn1mFk8DVGPhU7Oc+h3wqG2ZKy5mSJsRKBFqcWqo3Bga2Di
BjZebl7GK6YjmvmY/09EeSxUPOF0lLFZ8tuc3ALMSKDcYLLMx1imNPIwgmKmr40xq1tqXckHCeVK
Vurk7NEsLf7AQx+t7evntHwE3c4BZxPM7mHtI/66BjdgAbZBERQWsbmOL7r05hecyOlBINfM24QU
9WshdZMhPKeOhT64i1f1tNQxsqjLYBmcFt+ECDhPel6MrA1uH7MXZ1CAw225sXvDsAG7EWqfocPQ
cBcsy09YUNL5r5/qN2XTzMT7n7Vez+RvSxPDdIZOY2f06VzLBaCRfhqIGbPzusSAEnjDrqhDtDTB
bHoq9wTl9+mLpp6Kpp8KC477lFyDaZIdHvzykNkLMgkvRgx2U/T0jfmRp/683PVhqOAqs83NfGi5
5/b6CLfolJKUW0+Mbz6ioA96bnE0qu8b9ny3Oe1GUKJD+bGauRAAkGuFhEhtyDWOJps4Nit32+jg
R3/l34jRRC1jEozmV8HUdUGusKNl0OvzBlAJb8ov+NcBBDg+MnR1iq+kh4qYA+QXDFdwxdhg8ST3
wlXxaAVX5wn4B3HJasp4ey8SPu8qdlJLMnLo5AamscwnlJggaWJoPipn/YEBvNckDBPHM72XoL3O
W099yZZLBtlAcS27+54J6RLeRDbqWa+QtY6mgpyUTyGZ7hOeiUQ34G88K4foWkIGsSNJg62kxamh
seAPR6C2y5k0noOJNN+zKYthjTd0oPhKnFb4nuEx5j19/FgcUXLRXJgwSjccVxeTvb5Sfg0W7KCF
fd2+JJyMM7568BgvugmlfcW1Z9SOieGL7hF8mFAYHpO+NDh+wfXjT/Cu8uX6kb2Mv3x3RwI6bN+8
i3CW2D05okcAXNoJIe6zRHp5qh+sM4ZQ+VXD+vcsDAR1eHGPLw/AMDfm05c9oabiXTGhbT0m1zJh
9G0toZOxVIb5yuv4rjehLDdw6ubhmGM2QK5aL+oM9ukzWayZHFPoFL/VBmy9cFbFuc9H6w7l+Y1+
SKUtB23xkaCRJ5KyAWW9tslpQ0pLIcGRFYa76Wtiq41PHtUM5ufdIjIJBNFiTgjWECZpr0gvmgbz
bjuy4uE8wM9Sp8nKZBhCfm1fPtqKjkSgJiKSqKRcFfUwGj1t27vW1ywAvqL/x34A0UFIHF5wCsPg
e/yGS3k4xCBoXkTwczpIO4XICalEjLwwgWXLaERUEWiI8YPbitBabgB1xBIML/UV2cFcBHKsHAnD
PveLras4yvM4VDsQ8WREFyhtjLJh87o3wRtUfXSmEGptg02oDI0s5fKxpVGkeqXTr6Bud+U/hICj
91WscPQITJbjXnbhfZOfeml+FsvCn1Lxq8yDhcUEc0a1GLnzYpvLyI5z2BQ4FJXCmyGWPBeJEKm4
t3N1rIjMubs+ekZFRuSJE89Iu18Dkilx2oR12+NCv0+inGBZU9p6iIZ18ufoxr+7i3KFS55lD9tS
7Sun1fCrXVaWJ2x0eiUHG+3nJhRtFTKZZlbQgHlwnZRASAYCKkOmGeNxTgQ7Exs0Ju5EglRoCCYj
BOcJJIS9C0Lpg/FIbenjKlvNLMOO6u9yOIuCmfVxaxcYzORc8oTOnKRmmuPdgF9v5mgy3z8iYWks
5hA91A2nggSMcVsAwnsKSjsrWHhVQWTqpcBkZVSIsOiYPAjPbrxcPKgktg+U2RixcQlElNrS6wlx
AXpdJC5kLbyc5bdR5rn548aCn1IK6rm/d9n/UxmcASP2I42Sos7QUq1YG3eRNJsCuKeNI4wE3jFh
IvXewiaT7QiVkseTrQkdJoBOrrXOhFGmZms22CngWlnRuOkThFSeXmycMKuLI6VnL5nmwOW4/Kbv
2cVOlO+KUC8eYh/GUjNlH7yfB1DyRWt6RkrcvBh7EYDfc16quIUFq4zjfBqOyr/dooS5thWufOkF
/l5KcMIzrS9+iO3Plllf1CZlkflYD+7wgA5bYUe9y3+/FcnvsEt93DWwXd2475wo5Qa8ZDUSyQrD
QSCmF/ro5BcoZ65L07MnUAbNnh86FDgfwGMcJ7EuIabdTp1oyJDcmROGXJOJlZlYu7bm3YD9S5S3
rqTC+ty1EtyEhPq0RUqUqxjGSWqig/X/cNzwsOskuxhZJaO9KstdoQw0gMSXSvgBltDFQQr7BSr8
MLg35SEBWbVmy0Ut628qm+T94Qd986i8MZJ5JdkwtxK7WtRDyA50RcdAM11y7yiTPXofGYGAhCg8
P/xX/spa0uUQU8//4lTNR2kJtf5lWcL7WdN9fISK/HnRLmI4Hu0YD4KcOtQt9g1HXHme2bHj9VRv
0GuG22pf3U+jgMJBmKzpWe4yTpxqoLZE2RfmJOhyhpL9gQeHRnXP+4liZTxSJUgz9ca5PtrMGMro
YlTIWvXN/rj2CT/jqSRsiPESxC/nXwmgy05XU3P6sJVuIOUnQttENCHswq/Qkcf6H0TzYNReLl5p
QWAvhyRZCxvSnLY2+jWc/SuwsOS2T7ZCNb4KYaUVhbN8Zyh7HOn7do5iz2pOefdFJEP+fZPzNhMb
PzeiAo1oXN5sAfYoZEV3ILLXSpAcD6f9gaEjLZGIOaDYsFtx2H1SL3Xevcxdjd+sDvGN84zxHygk
45LJatZJImR2w4T8h1LY8MualA0w3k6jk08Fsl4SePLSzyLwP7BBBj1zZdQU2MBDlLWXPP+XM9VF
tk4VCUoJVFgAqbInVi7vjX2nx1gn8+MvefnazeWIHsimj57S2+4Zc1/tw3HAr0GjoSbvyrx3ZNWi
eHH9LFKOyz198KwuR7i4DfL2ttwv8tkn4IQVgjqRkExpGxOMuMhJKekQDsueBHxLODTvM6e2B62A
uDpxWvMorsObE272Pcqx3jO8aEm8fkP4ByTdcxlznZRC9Wceh+etd8XjiywOfyQgWP66Sb14g4FW
C+kJR/maMuzCk5fJ1RrTGZ83yu6jU208R28lTrtBz/fwBZGih35H4MG6M6gbjnGMnRAXneNaXldQ
GX8nX38KCENGWdZUilJ3k8aM1ye+IWwUb1jQPcfi5t06mlhUiSnJn2xeYS86hGkn20LVMVI4AyFq
YYCEKH/iF6uFqE5JE351StNw/uBKhAQJazG9J7wbwqwKc/EZ7vCkWRI6FTiRDCUnlOp4f5EB9+eP
v0DkNy7JMZpvapQCC6yDDv3R8O/ZC9c1f3LEE07Pze8YgGQnRMUT+NermJ/5qdKCswF7j/nQb7WN
3NULGVWkokVXwsPb+cuO5yZCdfl4AdDs7UQYfzwZ/9LGhlzaa76Ztvm92q9tuue4PaMoIMcptsO8
0BiRCHYHlpi5hxAPDm66pR1uuyB271+ddOTzYF2WFwQeMXk/cXdZjDBObrh6fJSFZ6wiE9iLUT/6
50I+F6RJrFzeG01O//VVp4ZPmPE+9gG9pPJqyC82wJdBhmahAmoGlRPrVwiY8mcntq5UmaNj/kWm
1a6+nZ539+nrUikSk/h20bXLkPAHEwwPKxrIJ2xKLAnwGtbZV/AaBeVHgYGBuPAR9VUqGQQz4iNT
IjpDRrTR1AqBXWf10OeEMSq13B32S5rqc32qf0wCi73h/on24SanoI5kryG+4BkiFuX+xURBpONw
m5oXz761OvjWfNioLiUwo62NBD9wR86W7gst7SufvX21QpKtkptkJquSZScuwwbzJ89jymacE7lx
aEM2wfoFF4vYzo0U2pGecTLHOhUCGJCJNmolQYvRLmMMlr2SRp10NxopN1TSdC0QnHc43AWqxf7H
3OwK3okdnDjO+Omdt57kujDJnQI+AKZa4pjfD61+twCD/KxC40pog3FeUONGtbyldLnUF7Pk07d9
NYkVlJieWUEYq5+VPa6xkiBCipTAjMnUVgL8cZyqSqimWHD7WER8kzYhMltiGDE5HLVRLGTVz2Gg
BZcNjsch1gZO18itP75ubzlcll9OJ1qqv2GQbXdSEPo6De0uKBikZUf2hWEfFLI7YfpcCddsjhY6
kYK9RUYqyHEpelbrasfuq0Xvr8vMJsBi4ZPvhan4jjzRDyPVj7SL4tTu1vpQtCTdPv4GjV81F+yZ
b/92wX8a01fwUZrrCoXGxRiEHh3yV6X7HXC8EaHtYFMfjQenjRWpC2j2Tmgk9h3dNyzjN+IIwHf9
re1zkQaNr0eFrqE6XRw7zQFAzi4wBJ2nk3t2PQml1KODyoltKMzkvn2yV/9sOteIcEaAX6Sq52gf
f2+TrhYQWV7kcm8Z0oOwuIQ+dbbSWJIeWny7eMD8YFhPHClj8sLKX9e8jNeYoTr1jcnP8mIjzj4Y
GGyUZbqVCFqyJ6/KsjOzD7b9FaHSmuGYUfF+KQE1L0SGqAw2CfLYVFf2iBR/Ep0w3m0Mti53fdB3
EeAurQDwSh0EIMNDWa479I/z/N00tdvHa3VDi2JV8toQn+mWWrua3HdIoB7HKBjbcfN7W6MlpUFq
86CL1lUfFJznrWf9B1tD47duet8deYbr6upmq6dvpQJKiHiOpzZ+Ngxm/y/3nDReIx7MGmVR+ULv
Tu5Hk5No2cwVLvEY+789iIUE9m1s1qrkjuVenZAIuaqMA/T3MSW+iUv9mo5oV4YyEmpJmK3zpS++
milaLiZxTkl5T9so2B5Vcr9YCYfV5tYut4A1xPH5GX2LpMIQEcac40rkVfVbkuGlBkOLSfQYWI06
QuI6uV7yMZTTCGcZTxgRjBM5Y6jmammu+QD+Nl0Ak3jodmxJDwPs6kuv4U+hjcBuTabkdj2q78vG
Gpml7DEDjkkr6AZ1JWCchBb864aOw57RLX8HU2vFzX9X7Ow/eng5e2UkeU5vn5hKXm0YW+LtY88/
/8TyGDZg9H4j8ly7sEJ7vxC6EhHWnl5EG3/NdLaLB3+tS81hpafxBzcbNnhUJ+tjQ8AtPshUraEX
tFHhPDNxeNw8n4u4at+Azp2ujgSb1cckZiwRdHlP7w08BF4dmVq5ywJfds2G7AMMUEX9/Dpnkt9D
p6Ma2rY96YCo7a2oUEjKa8FxJXbFGrAgPET2j3qf4VkH7YWa2stjU4kBoPire+OACWk8Bc5t2mCR
YboR1SOdOMkd3mr4oeTuRF6KC4Cjbtw2iyRzzzBpYM0atp8Azgmw68R/homdAklBOVWViUdCUdBk
jTAMKnISlHhDwN7Hr1/sny3nk2f/ztRwGfBl0R2fZ86o2RIb2y4tSJAvmHf3uAC5PaA5wvgjj2V9
PJiGBfxdZ3EpUlqEpKpZXHhKoYko8GeLIpDMkMo68Awheg7FklE6+FL6a0+ziCsQNJnpnBuOSfQX
468LppcwVU/3E0o5UOQddX2gT5J4dLyJQbHNPZGgM7Fpj7t3zpNBe1BAzO7uekNlZDSAjR0w72mL
2+PB1PkTjMHnWRdzjLR6au65l4FL3v+QQr/uY3+vL8ufF30OZ+EdYc5ifXMB8DA3W83UTuQ5WdYu
KJW+bG/mRLK1Iwt/iesR8DLlCdkl4mhkfQWhi+hDTHslYQ+BIR4qWPz/TzMaVmBx9GgMjtM8J8ib
e2OYD2Aba88XnxPwpHVzEA3EJrckZ/5vgG7tJZnjR8E3UN9m7wg3FHppmrJFgyBFSvYAZHugLUhY
En4kzfbofkMJ9nW3N4QHH30IIm73mSu/SZRqFdQmgA9YOG7TYi87qsCoLQFnr9kv8SA+1bZ7pXZd
Pngp+ran5jWeP6SOf7hrSQ4BcYJbSNtlJnYEmPvjuxSEc7fbNcG7iOKtbIGNcusiJ3szdSkYAmbG
VbGcSZAgpCk7py7/g6KISYNvMeUj+keZoqjRIzKLVkdLbFRPCEAvk0cYlLSN005lrwsCxv7F64qp
2hHGWs4DxWQeKtAiw2JVUUsB3WlKz4HmvgH26g67zeHHDet8B/x5jCyxhkfAWAAzL3C/fD7i2h+s
ZYXU+J9Ah/FwZSSN2Ul++wnE6J59ssVevwFYM/f1SligAWt2m+mPKQ18WIo7HbsowV9RZNr9rY44
1NcwFVwTv++yrg06WMhcmnwyspuqkl9y72AFkLnNbxeNLmYguZ9zSfU3lbivh8a57QpMsbNfAx9/
mYcf/1LQrVEm7Bb6Iqifr3g4OlNrULTLaZI88D0LaBto6+smn57DxS6FBPPBs+c9AJ4SH4/GZHWz
3ypWFOLQDq2Xgs9FbHxEmkGx3e3JZ1/H5F2fgWz3SGAVmbcI/l2xL2hjCt4Hh+sbumQ3Yv08Q+N1
1IVGPwl9RpFe+ewfxuYDwz16t6FoKex6qLKVBgEbz3PfXEDVeiEeaq0Z2dBe+8tOg7duMROhYlRE
hqNv1xgKecHXaxMHryVGFHRtVAkFfIwy+4Mpbo29xxY6KLjx0LTTaCKjpZrjEQp6euA5LrPTB2m1
CMjlMwyRDfa595sT9CYHA58+0k74+cAqXzDC9cvEuUzzS1lOjQhGEj3BxMPRKcRluc2+caJY1ByA
tD/HUapMZ/VgQB+e5esCkVl/y7BtqzU25zm7C5BE1CcC5YwMKqeIDa7t7IdNUcgvO1IUaqJco8re
FbewE5pBmhFjgH+Ng0fMoStsYtZcx1SYAiZKtK33sXezGAH/UA/XWmymvod/wv7FKkdL+q7D6GS7
ar/5S98BRUUSP1ka2DE09zNPUygfRSvOZbTINXa5fTimQCyZ0UTiB90Xxp91PMw6aLhp0J3GMzcK
sISpN70cBOzUSwb7kSA3hVZ3aHskB5UYUTQTI3u69dSgZZ3J5EqD9y1rhOFH+yLnrsMIUhn/wNG5
avwEQAz0pSUEFF6CXtgBv3FW/jFsWDgYkc7jMj0ygmIjVExC/gbhBvXmjny3X/VDZuVQ54spTX3X
ASF7Oo+L3eU7ifs1pknvRR1UOEcCQaK9D2IN+scyEx2d8UYmAzGQPujdLjv2EaFIyiLdAyNsiYV+
H21DKc7sJEFN+TLfWyHpzHIf+OfSS9LcEx9lBd4xV2Dq5iNPflsUomOtPlKb23elBN4sFLnnbx+O
LroVB8yUHT7NKSRY5IVS6ED2rv1MHduc6oF7Q21zPh5FGoP81QYsnyv99W0skdvBec6p+jOK6N2D
dXuzujLk9jkhwn5iGNIjqtWjBCIiNbRLbQcessRS8CJPuHHI6ZgNCYhwgUXvYymVCUzVgdX0M5X+
WugjJsOEZn6mlGv2airRF74Uc5lPX/D89ug/T4/u0HD3qAc+ASyoV2imH4kYBFz5dXajeymaO3hL
VrkzwXnV3jiQSjt9qPeGc+2d2EPNFXupcoFkJfvR1IgToKnoPTxCeyDgBjgauAzk95FVrK14OECR
OdEOxWWkSwnPgGGguB5PR+fvEknz8kTJbvQqvWgrzXEclntKHj7qc5PQp/9XEgviwxKnwOilGAlK
ZoiPeBoANUDgjjkYEnMrE6CM7ZH7jq6d2YmqFPTrKYwI0ij23N4dXZV5segDioz5Myc3pdyiisEu
+6ne1vuvTK8M7aQUbvFuET3K767Fr71JVCkQHDjDTGUtoGDYlyDvEs9+2NGqsWv5/EpM5WxX3Hsj
wDGt5542eBi2K0LxSw6aMrWbVBoWECZyMxXjpxciapWOkKO7Wi41ceAm8OJrLKHPkqle0OxqY6q/
IjqcGhqZeMpKsuIf4I8hoWsPg8ghO3xYihlYiMLtXSTzxgQTNWXCGdHl3TFesr5osNXCZegwsKnO
81J09/6lq8H92NQq+Z2kHEg7y93+KASEk+0tZP5QiyNOYmhFskWMmYADyCad+Do1bTBkmVmLqSHl
MIc6quhG1ZfZO2XVxi4Xdkh+hZPe23sxmf5hteL8C1u6v9ZFY8nHEoY3tm0jDgkwrikmodL9uj9e
0VQBc15tC75rA7GeA8i8cnLRz0ka30ZU2IsLoUf21qkQS2PzFayDviZ254hnMj4ntFdPGUgQ/sHf
Pj3M8s2Uc0TkH+LTjvdlqJyV0Ln8oMeEAxogbgtU9UNK+mHkDSrAjC3SJrFZjUOL3hsN6uxhWbbZ
NhJlKiRsw15yXQMW1D1b0Oq12omrf9+yMrRaYCM/GJ/lH5ejhw+SNwc3eJk6hKZ0ilpAPcuPjqbr
y7Tk8wV7tkz8RA7oI3iGKPA8fflROHYDCNlhfgimDIMHlFSc5TjSccBckIc+rY6A64PN/+ozAjtM
jgxuwiMMyuLbu0412MvW6u+ATE32s/6I20dei33bPX8PRCTlyQ70ad7OGHYSFLcJ/9vQt2VPWkN/
liqkLEman2pd/hqsDTRs98ZMC9c4yXwyGfHYk5WLssHrAcG1f63zGL7b3rwCnz6AFwaGLIdR9dte
P++mjSAfmcl76IeJsc3o2nbgLPIsJKtSXTRRcCFdZn0+dJ45MagSLiRGKFYDEI3kPoYIkleRIt54
hCf8yQ6vYJt4Frnp+QU+DGIdXpoxJ20EoEZ5kqPhx5PczhmHJE/xzu5Th8odEyBSw01O79VStNgC
kXDwt2LfoU3S2jCYxz8Ycf3TSvYSkEyRwTYFuBv2+1rO+++2Hg19vaaForTAHCpvtzajwnBdEH5C
5h9kcsdZPgly2IJ2RxMvcwJSHyYYcJ575/IfXMbHLONjtP5klTVSzdTMoLCMMJS/qp2pP3KKfk6T
Ik2YzGcbVhIsH0Oq+17rYfZcVtrENhXxURt4Vp79bKY2eAonoWTZW2RuHiuHcGWSVyT4Cm9L51I7
Kyn1+QMBl+EK4TbowPrsj2rie4JeZcTxineblx42fm3NjvvWj1X5wlLCzb3zpSEHhssEYLqljaQo
MAQ92fjNhvMXVnTnWSjpY1+XYGkmccurI59k84UzmU9jzXe4CX1EJMaOtPvYRRA4JC4usMLm3ZgB
Pu9+zYW3leIj46do0tUaTUDgP4SOglAdSDso30e4rdAkspZt+ZVvjkYIaanqhXJzvtwA2S/bHx/T
UdhkVr4EFBDd6gWii2pXj3y89oB6o7vi2iWa6qBwGCWnhwc2/NYKCgv4/uBqi3Jbt3dRk26Fnf4c
oAJUleknK8ARAKd+ePzUKNvzEWLzDfWJd3tACy/GILXegkGhCBYCIlGA0bRVmw/PUxSRmNTN122V
Bgzyz8mPKTkMPE8CdZZMx7iDb3VNX48wxZDa6y1uQXGC/9WqXOIt3/+cy+xOYg6av3XaLRkcfLB9
usstz/z+Wwd6JcHS3Sijv3dclwdGURTkSNm8Z59yMfp3wlP17bQJGy6wHYrwfUJyDRX53cRO8XkO
5v98Ywl9w3Di98XaWSurEyQvQfUpeXnSIPzo0qq4fRB551xOKsie5lGCKvnbUtfVeeApm4hdSVQg
6tJhek/x1//lXFRD7HfY+x4uN6/28U9f8UH64lH41akCEVJJVyIP/Lp8cBvtCcxaLr1yhjJ+g3ba
tbBdpy5o4GE4bgRnCK4OB7VpU/RVeYwWxw9yMTA+ppnHehVhm2TzsBG/bc2NATW6RvnAXKuS9dy/
Magu1KHPno/MEFjMmxmGG8uPtXAVMcKs3ST5yMILNm6XvgQHTBe3FNylp6ycjG/CYVyH2STNiUu/
q5IpEpdfJOzRaggbNAaKgBrKE//5LBTieXIjUopa0ETK7M221XrLuWaxeL/fyJSXPzsUlsN4TVd/
IjDobOIq+2e1wYJSKxXWL+ewwcKTibrKBYbnLr3PflB5Ms02FmMHoVjv23PfGJs+RNsS7z/M81Pb
8eaebippM9tpaLeox92l8crme6VlpDDjqByon+y4XoJcCf3DucqCMTePYWG42H4ifMcj8HSiQd+D
UUl23yyJxEYD/f7j6gWjIfx7BkadTyBX78pJDHRKPikJF6KdCgt/g7yHgP4/fi88rV4hDT7KKaTE
Fb2fDC/N+Zn+g9gDBiRIX8ALw1oAfNbfnQPeg8cy2CML4LuS3Dcvd41XTaouct3LHY6SGh8+7Vn4
+CCDuHVdTEfzm9dQtufG2lhwThWv9CR8ywnrdX2/djxt5bMVtl3U2lePOqaKudZU4NfdDjV2Qdvd
t0CojEBFxi9YP4aBULDdNnqeZLzAUWYa6DpcgrQDRKnivOKMYbFvoKVAMhkE7/oY2XbEhZ42T5iW
okSRCQSqRA9Nvrd9qmlu603/ycYhXEZt0uyWyxDysUgVqkeILFpSl5WExYt7COI2CzsLv66wdGpZ
+MBc6RTwyjHPTS0/y9aAfSvRE69HAXdv4oYvzl/wGFnXVk6E+W64yCLHo4s26aSqm3Oi7Uz+F63O
n4SIsIrJn1FPCZ3x/yIF2uffVc2Tc/OvNe9zUcaxO+lBXVbVk2QUy4bmFsQXPn2FeO353iqRDckh
hLdRiQhNvYBx5RniJ0uSzsP0bfZSOHulKt+rPcHT2O6jp36+pizK0StIc3tjU3YzQGu1nvdsLpEM
UIRbTzJVHrJ7gury9+Tc5cgl/yDR4pv6HKWQ6+Ki+FI4Q2rRCUeKyv3wfTqMF56SqtW5pq37Wj5R
DKY3hOdgDg3LE/jRvpz18tUAEEBebmECjNBMQ2P9GkODOqh/kTCT+KWm7XvB9xSD1Qs5yojBedIe
Xmu+cOvElx51ZgALlPB+P0xzxIM7+ootyvT6D23UrpEFReDEnC9C/EBAmuTiHNj6luKN+2rpFazJ
luOGHSOyYAAXYFH84H5Z+oSj7553Bf95GleLxP2kvgHMbAad8UuzqrLlPl/G66RvUMPIUvnMJ5v1
YpWFeGLpdjw/2zfZknRMnmAbDOiXNojulB/6xHWhxVR9CBScQclYFXKYMLk+nQZ4B8f1/ctuX9z/
aLcd8ONey9LTxWlosiO9+PvuDMTu1CpnpC8v41UK38ozUr2xaP1QNJKMFkCYf99Mytx99WS7O2IT
rS8QXaHAQJfv/tIIQQj0C7UAhmE+qIxgGAswQCh0rWBrzKL1KmKcqw32gEjcwBZQZUt7KmhY7pmw
pG4PzJPXkOKDSEHsHCcwfEZ97tkaqFisR/vNETSPZx8UqPefWikZUCvrl5i/+Lb5LezfpCl6O7fB
Rt6natYr2jUM1uG4yEpeABCoO+7R7MZw6QxInsmf7i4gjiote+u6IOJbyi2ybQaxRXUFr7xRk2bE
l6v69kurziFxbJyR7Kaa5U/y7qVv1Zmf8E+Iro5ZexrWrz+4lalP2XQxCcvoc1pxPajMuYFYHigZ
9bjQVS2b15mO9Yij9Ah+wvUSuEVjLgq6HTsS/o9eII6qgGoBRnLR4kRSUiXXYVhYMsgvL1V3AntF
mgblkI/0UOjjdQHUVU5L8iVzBVD4M7+51ld4wOcrNCCYPNp7zyCGOEBzjQpWySXp8SAD9TQp4WKZ
CBNfuL1QfZNFgFejS7S0vHDhv/90O0FSTSqXGeKyhotkxI519+/yr3OUIYTvc1uDtEkbYnrwZgxf
w/KtynRza9/xe2b2FTA5pW5jH1h4Zxp65DSVt39q8Ayr04SJgzcf7C4eEQ6fYdd1aSpz6iq56j1V
6B/1OLmMe2oH1AQXV8ScyIVN5StuYjxi1i01y2c5j1LpQwrmmOh/zGOzKm5SeFAISGECKphpgNxC
zOVOD0QQQDqQNn14QLPYgbB2TR/PXvj/UpJiHsgAwCTDlWkjrcidGTyexJOriy18G0uCK4KTimD0
Ms6cXQyHN8T1XuRYbM1XmBmy5kscO/gBa7djK9otwgBNLKJrfv1mGfnQlrDytHkGWGLlkV0yZ3vn
O/nu662Aj7R9xEtiifdYfba61kMx4tAo4qDcfQoqEAov7751438t0KYo33ME/KGZm/Az3b2ZGpZj
UAA1HDRSH1kgXf/meBvNjhgIn0bmM+N4vM1KhGqXEyAgJZ2CC7yEYnZJhVdqWldJsHoiOGec4v82
r7JM3dCDkQ91CBUZJjfjFnunFRQhhErrvdc0rqHi9AiRghiZpMpKBAFMF33UaeNQk8gM5BYOxwD4
8TXaqOpufbtkSHcyk+wXzAH/UcyjsYW969UFHx712E7AsLcavLv6JRtba4zlp31K4wsoTq02dyLH
PNUm9lfMfVUPzI+0QACaO1tplILe6q+5QB81ITqAruONz9chcGsQHvStGtzlFBbx898gSMvxMW00
ZEBLii/rAshmeI8Ttw12KnJ0YgphYoigZXb0XJyTj29Obhw/50QDnL4coKB2e4jGqBo9xTsYXLxV
PeXImfJ4uKhBdE7HWM2kUM/ZAySa8yBgqSu6kwj+7kWHqMuHbof4GCZ2uPULY7KADQu7oU0pHUBT
0QjkZ8zmh7BsKPxwAqIEk/mrbHYGnTRtzLGAdvgHLjWEwVZJxMn6ipxjKsSpr8z6dnR4s07WWoDj
v46Gn90VEqxJ18KMMD6HhQEgdn21Ud5fJpu8CVlpGTxMMJcsulyau7xx1ZVdprvyPYbEPpZAvR0s
MRldyQP2q2+lkFOyiOfC6TqpyWF/89rxOsRt8HftMB8LuCK/bSnzC4nci0wtkvHHm8y66PPQtkh7
S+RRtPzNzJ6LvTE7Z2ZYvYwpcQrD8p7sfzdF7RODvbS5eJKoxD+lF08MkYnkV+Y8mR+qZTibIjhG
Nl8chvqzGz4mva8wZh0u2cD6OrATJiMcUWlRmPv4TvOYx7ts8sVgssS1Z2qPhiZBVzX/eV4jDaVs
mSeaf3ZhMY48Hhttsbqa92c9FC+a//62pf3dd6Y+sRLkZ5xi1qtiVI/+cCaoQXp0rlfk+3I5g33r
kZZfEs03FYC44rQrZ+QuMwrht/1HDIp+XnIAJnsYO2aT57QBCWjKZ08N3ve6IS5cW1GUfCwuqFbA
sS52jxAkiVcWbCZP8idwCrw/+HqBDfV8faoL76bi4VJPUlqnq2iMso0+Z7QXpshiD9Qzq8D+Olu7
ocPn9uU15KdnB8/3DEJBESRbKNSx1IZb8e5s9tUykFyV5dCNVCTmeSXlbW35QbmlovCYT3zgfgip
tuqifAbgAjUEDwqM785U3vpkv+o2GYltMuK99BJLGcVKFFwT+yHG9C6s+TzsN0hBb1pn5cCzmf81
aH/I2D0bxWh6LfrwyDJSLcGouS72yAgt57zDG+dXcB62ilMv5ASfBFiyQPn2mJ6dqHf0NEFqWB05
SqDDyeZ58JZpPhERUBWZI599UIS5/OPNxzMW+YldiiizT3nGKtjqO20b2BEGpeYXQuHF5bridKNU
i6wd1XmOMHb8Gv2GQ+H+QMDjwp1lX9bcXqHE1eYHgUTNWoTXQaE8QAFgSBZR0v1UPnkZDs78Ic2P
oi7RQ1FzCWch6XbZEM9JnTCSI4EiqHY4BDMVkpTsHccQeA2KTyKEC5ZNeR0QpjVI2ccTgsHCErif
24p+a48+TsC3HxcY+kmYa1lzMWTO/IkUSeVKON/CR9XUIQsZcgNlRAi8xoNw7VoX98HlWzF3R32E
pHZwShdcs55Nct1hViaol3VLzPfPpxMMLBRuYSMK8WrpOX/Z2mDrone6fgEfCDC+PdevVQcSK1gc
A7tdpv3Q31N3MzsRyAAJ4aoJN9A1defhmGDRzsaWC5uN4zaNHsIWUj5C2l87NTPATzjnnwRi/j+R
jwAwgOCUxI35HiRNyCyMAk1fGAGsw/uAzshETnDfCppefwLXDucoFJdGR1dC4fFKzAjGzM6yaF2Y
FEb7SwWJno+pzsUkGNrLUxR3jQgkN1litCA3XAz6H70pBTcK/Em7fOAVvH5jAuI4lPpW44YgCMI8
bX3eCnA2HlToAhxRJZxgVQNyUsEOKWiVRjAH9IijvlrkBAgBe3xI1zWOiNCl9t1oXPbyNTzEWEhc
Byx9tu2P4ZXMU64Hsu1QASLff1n4NvLmNnRvKZ2sWnJeHrIbB6AzC2D+3+CxbobgbftF/QYAFbFx
+IcviEs37+gWb/eWs8rziwS3N6WoTCgV/tcrQTiQ+50SEA+dGLbAs5NGjG8ECpRl76oOaifeoMtf
DPW3bzsck1pH3nE76J19UCd5tPlcwwHnikx96Afe/efX22e0VCbnN07T85pB0wrIg/9rKNEARUgj
MNXP8z7lcmxXRyvpck94FwCkZ5qwOrLV8FvjvhcOCieEjF7OSIKYybIv7aWepbAJniGV+5cEVRjb
STIVEw0zUGIOLQO1l1e3K9yoLHABLrPoyScju2FecOp9hBFQeKs4Fr5exgM7olcS/WIjhfv/PVVr
0xzc3lJ8kzRz6n2OOECWgupbW2OrJM7NHsEAPJlhgh1V/8I9nVsYHK+oK9hMt5+BQ5Vw3GjeN/sF
UjLkjUxDnWoLFCwtYkAnY9IkuEfPKSZ83jlHgL8ZSQ2+QRdtiSoHTeEx+Bd5RyVOirnWxLLM8VW/
JH3F4OSmdTSC2aEZopd1eD3DDzWdCH3HvyrzKbepSWYZFhL4FkIUOdPFifCIz1JGs7L/M0ggtqeJ
hZBlIVT87InoYgUccIcZoBL2ZLeo1WLG15W3zJN57roPlYztFMqQHsMFenVZyLbo2QmJTlel+PR4
nSC8LgGkrziQ0pZ7VY179idBUK0gnsv+E/0WP8NhZ8m72COoXR2ODsBK37I4nUZs1JiC6FMn4XZg
eOVXZJjQ2/CnVhE0JO+YtNy4fVl/9RRwX0moRs8cgWAf+3xRoNtxkCJcpG9IvdIaL25OJrlTZVQl
hdkogK43pYYhl0FUT3T4BuRUOEEMag6NE2fOFaGMlY9OITu791V0GcH4zJhdnzTPAJKtJbSRcJ7W
0q6gah9V8/gWJE/KrtnuCkfHQV5RVJE5LUnWZdtLO1ofRdGwo4TiW9eIminQTeCPJDHeP2G0eveK
ab2Gmu+hsZdVLuyZv7VzrA+G9erpJOsAZTOGFvnCsNA72HZTlNB/d+MOPCjH7EL2euaN9Rf1cY2h
RlY4pi2uBMjbEOVM9hs3BzVebc9Ben+ksUN6XV9lShw6yMOypQfYn/4ywdNL1wdQqC5LkUBKrA4P
Wp2d4nJpIWAjDUmnVW6H7kl7t/c4K08tbuWND/Q80O7OHYKq8NVU8LTWvnvcmGOtAZ+o1l40951O
KPIfwpTCA2dmLDx8gMpo2angoj23ttcYOdEYgHi2fJpbFHyffh6c5APcDvG9qtrVe3kSdrzCO0S8
bM0eqDpziqRMWQ4rnq/D5czUYByejawoeIw7HWaCfc16xi+iaZbgLTAfV9bB6egTCDFZtTPpvMq+
TAb74uhBFWyLYXGqZ+moikDAWxU0yPsoRnMULbHQpRxw9NK3uIYE2Y86jexHoQXNO71CCkTCRKa/
u8PbkLuRMpkL7pmznbZd4N/xDc+imhkzFA409xcvArdqr67PmqLmWw8GB2X/ASEKRDokz4Lnf1W6
LBWHtgfftQbL2zehG3UG1H4dla4yrmBpYHg/q6qQdaU5/sVS0MvJBCx5d+wpP0Y+cFXoR6eZQW22
gUH26Z3EPGwHGbRRsW8pmj4RJm2lHXVOVuwv0dHf+YdVjaA/NDK4xse3f3yTZkSNTHDRQi/U2s/s
+anCtBpfO+yJMzSn6UgcKXV1WivR40lHyV1m9+6VrRTOssH8zZFfvYRpemb8PlHZmmP2uyrhDYyB
0Pr2FvgE40ihgZlE3NdFYpI7z/9VYx7qhOXHxVIuE7yjnlOihn6MUQBnxsXi8highuEZZFSkUkmQ
vHKB2q3o/te3voSYQcoZ3kTMv6FVTN1VB6UODoebKyjxbbUZi5cHphjk4FDOSSdgMzAoNwygOElX
yNtgV9SRywdelw12mq2YvnYol1Nh7TkmubuNkxdQAWlVUw+9OCOQEKvOE7iK4CLu7rHJMz0Mzqyd
q5P6r+F+hguKOowzZoZuu3fhtqi6Go9tfFNrIK8iZ9OnDkRY30BUrQfrMbejLhIxjWzI2G2zNvCS
sY5q98TJ92jPdLu95g4l1C19IeyUiR8Ts5yjiXKbFsjZ2pXZOLXxReICyAhxuRXq404adEEmDmGH
BQWX3YhlDUSF6WGQii9etmklconq1XYs0iLfTgocKcWEwLkZ+UPb/wufQvj8ULZyIWZu/hcsVUd0
Jkk4lMDUgatp5vyYUVHEXp99KDE9F4NMmikiIpfFUYfFssBggGPBEylpj1yZuEA2I/J5154QHF+a
Y0763X9LqbVm2YVC+WCCzU/Lv71WTL0+YQNp5meaOG24SJNGXpqUAW+6cdA5STgk0fjzRx3d0rw4
AtsZ3IZeDjfJJJy3BD5yFPkFzYGHs8ZSA+FSane4l7Y9i8cvFP9chx9RfbUTcNcwNMSmp9T6Am0r
of0+QGf7mK6D943EryPaRn+pehdQDn0hEpU2cJh4qAx1YdOId2EhIb4K47cFzbGvh1+r7lspjsKt
RZyOcq0BLYgajK90ulxCnH+vJVGP+P0YTGS5YTCa+m+RVUjEixepUJYqOQv0bKVmlgHVbgNn+eJN
SrNEnACV1BPNNIgE88Urb9zXm+je4r2DHN3TC8DAtHqMxMIcDfIuuX8aejN+y3K02nubEcQVftj9
BARS5xNoU1CL9BYZ4VTLNQOvcMsdHJ2JeMvNqmd1plRi+ZLeMvRg6H6iQWfUTcAOWkMMa6Reh5Ml
V8MKKA3U4rBnEembRPZAYoMsKPIk+gkNT3IiSAgkwQALIm9gVXaoYFElNPGZi+JBvvi2jh3iaDS+
MucPlQvKfrF7eO9QxUgsWLZEmGmTiIWjzZxrXRK4Ey91O1OASJiQ/4R6JAvpsHnxong8ZhBYOBSn
2UvleqtEBWkKol9ZUkhhf0prcbhXvTaKEFIl4x8b8jEwSaLezOxZ/butU5N7AWEajcH3aO+biWTe
OD61ydAi+NQSRxmmteUumJstIwess2qAfdobg1NucGZeBcJMDS0KcR33rBqGWQLO/jR3apkazptv
s5on9ulfXhu3tLJu7tcvhQJfogPMTL5RbNzDvJO9CvY6ZKaxinRHB6JfJFjnv/e8sllzmNqRn1co
jtgxODho6Q2niUDf7a3pUJYXMd6AazfN5cihiuoPFoidQmgQyUVUa+Pdun3JN+0Cc66Y1OD+FA5E
dM6b2zsz9MrMMW/OYSXggfMao+pxJlT1eVSDL8MSUVDliYx5nBs5AEvwekgq8U0Djt1c0gA378ah
2/Xd5iCv+z5aF4iDw87RBKbthhWLFb5pmI8h8jNh0RmoWEQma9k2lNFCltXhhM9CUdytEcijd8kv
9G6cZ8cu1CBvzsaZEWTB/gKdMNdicnGHGE0AIi42F9I+meDoarQMLRyjB7D+Eo02N6oRkdiLPZIS
4As1s6erYdMCdg2V4WgfYYTLeRxpbP7kZMQYf+NkVPiTPZGDaE73TiqEKhEct1i5JqzceskwnY/F
SCpOE7TwXgPkKCM9D2NuYMxp02I+kbGPw8z64uEBja3UbfS6D/1yEAuRQWuwsov9j32YIuVIVHPz
druAtTLc5NnquByjRn5Rp/gRuXCR+GgZugp2rkFfurWDCLyHbcs3ax1v3FvT7+9JK3To6lzD67i4
mh2bNxQtQ/maZgwHvGsltRAs/BYY03UgmuLg62si466iVMiW4Hrix/6Qppb83wea5ADYzCw9m6+o
Mit5ItP2nHKXGAtBZIEnjQux6Ty/cdH1X1Ws5zOGU278Ex+oPIat36cZ4kXsM6w8XCu5l2VDc0U1
gmA59mMW6AvpWR+XaTg1DwM2u7OWca8oEdWD9ZromkLfTr99NDYRiR1HsIGIP2MXAFMKf18MEt9V
OhCXKcv+ewQRIaRDKNjm+H5rj7zWmKUlGW4oCF73hWT0nC0FCnOBt4BoEOBB2uhn6/98GlnZULiA
GeoQMG7kcfNtcIKddS535WzPVnfcoD6ZaWusKL4Dv9nXkw/QscsK+yLFgiRdSU9qnJNhWLxZH+LZ
ZjuxwNlFYQWuopnwKc/02KYDY3mpii76ZtP/A6Y96qNlPc+lvo7TI1Bwmh0RNDGCoQ5KNc+LTrSJ
Y1ddqgWmDwqgvbA9NbQayfIL4h/NS4a2eShzoGmn5itvDfEVpOOwn0/FdgMU3rZ6HNVoUO+TAxNH
tMS/AA7YAd/Efjh59q5cKJyIdCxz9JiHHUGNocYJXIFWGcM0pf+7Kj9Zu8UeDGEpcc4JzuaabYkW
BUVRQJWNU3SzVovr5yzCPZZ7827pFrn+aCocYIT2ZpKkDHIH4XX/dV2E40yPbZgVpZPpNiStmoXg
0AzYWsWGI+pTkXwDNEU5B57hE991bH2eL99erowjRJIM64I3999cNI6Cz9xbH/XtpoM8q5PwFe+/
AGyLoTJ2pbmoCVU5eW6pdahgdcOgdzTp6WS51MMdWBUZMTOJqR3ZASfXAscOxnMI1F4VpBi1z2Te
P+PuHXA2P0WJlci3eHgVrILffxNmqP5IAZjSNP9gFyX9lbnrCQBVUJYtJZqoOIWcLFq4EqnU0nMT
Od4KOyE94xufizqlA8Z4gE6Srx0LC3elJnB3kiKL5d4IXZG/npXfCBzRBiw71+z1YJVMGPpUNmjJ
pWnlOR/wm2qb0GCt21ZPgF90kldKurR1gDP60voRSO96u6tx4y11+ec5hQ5vewOyErgocF/3Y9Ct
b6uSb5JJRUHq5jG1PFmG3Dw+T88PVKSByDoiz6LILv0ugHeSRKqn3g/KxuBCXvOzDW6KuwMROJWR
g3Sa9bIL7mmXj8bW2dvAnh3wnLTEQTO2RVgrzOr2dOMfiPgSy98QTWG/d2uMqOfy7nTCyQZe+VWO
/fi7DxJLceWkzvewoCwxtTa1SiE2BiOEdQTXrepS4nyPS+OI8qBIdMMtK898NxlFi1bh0AtC7cuI
fzZ2oMlNtQFDTFYIJUz2SLQDedDUyWwicDqdyjD/RgAB6X5KReAX2Ab0IXyKhOXCS+jiEeKpiK3g
W3+WtZ+DfVoWWKVw4aq+cfp6BOgsUfzNkJ/BwcA3qh/sYPiNfhakBZYZ5c5KOukxHuiBZulJ9hYl
eu9B3K3s39+b21JvW1+GAlkln9M/jAQYCSJgjVZul7i86BxTxHHnXZYgP1OJNZR+GSD7KUhaCZba
GnCLZh2xJRWXM8zt55gAdzpn18mrsq+5D45jLCqMtL7p+K7HaLmT3WWKtgC7Y3j0gOfqeBlwHwfo
MlT9U3IsK7EB8NWjihP/hYBTqOrMMmhi86EtfSQUlJofp0BSfmH8F2GbG3dQBZ7gl/iga4gmvH6c
FaZ07uMdhZcJnqWPQgvg3InEuSbaDkZ/Oqbx1rAjCkqbQeTn85R67v2OhEABdziTg/lDU4H+PxXK
V0cufNVa1ZMT8aXdRCWYQMT+8/yOUQubxqiUC9CYM+Dw9l8gW6TiZ6NfOgpzAgnaRZQ4zeuDzUGs
mPIZkHy/RSY+wvpbzSt3SlE+oaxuMK2228xjMtJYb/uZM/CLH8yX8up0PlJbb8n/gGxl6QrmvwAG
HhYZ+geN7aRZMu++J8UU2qVEJFZ1aqPPdpePOskkt0PBLWZOe7u2WVObV0tNhGsQQOgT9XhU4b0x
2SGfkEmNYZ3SYuPaOr6kOK6XVXbkqv8IT23vBYUUw/63UByf266HpUtpfJBZ/ZQgt/6I+iF75Pqc
XaPs+MDWXsQcRzD7Rx/H8Qg185arB/x2sH7YsONqQYytT1r34rDkel+YsKcUUalYmJ93m7lDWQDl
egx6EMRPMelfopTpmT06tLbN0Dq4QF+JhATJjr1e14QU6yXxxRBTYz+uK18yq50l/OTs9ikOrIs4
ptvWehdVnOwiF4C7sR1f1wgtHfbRm9YhN7YpQQjB37NqkTavNg9bjtthCQAc9w0E8wNIwiAkNxb3
TVXY3Ksx1p3exK38ICdg6jwgqJulYh+II+kWRB+a4/tYFwAXkNk79itLAbq3MyVfxT35uXZ6jGTD
MhMJ7Oli4OO/H72oX4Vh8CZDP+bsR1bTEqlfGnWD3sI8ovwDWrFGm/1IN9RKQIHleVk1GBrOlPuP
vx0VwlonFnCz5EPNucBeAwe2LnMZzbGnFfFk0rZdgiww2skyUeCSz86fuEUkRR29r3Y9ez5VA+6g
JkDqtJB92LRi2vkeFjOAo9vI1RzTQLJ1IObwRbse4S95u/B8L5NonRY7fkkfoXnVCUP6dPSMSpVO
bHYL4biSFuGJPajTFz5E5huvhmKadZ10Qf1nNrz0lhyibbOCrdsY3x9zLgFsx5tOHc86qCrVM8sP
z6XKuN2fF2SCeoQ5/0sOCDLHFACxfbcyKSxoRJGeGnxQYv/PuQNywYQi6LooL5MTh/XVCNGIn97W
+vK7qC0yb1xghTdoghFCC/JQXjfbFNVSkmjAEm0KksTLSICEkPnCk3pOGJkPs24O/EVuKiJY7zd/
4EE7+QXtxekxK0PIRR5+4q481V4u7yUYg/rZhvfy1lGjl80CAu6+aotdHN/GObGH0S3F0NvaX/ow
hjtS/KED2B2sIVlWw3A3XyeGpA5OKitEUiW1oXOpIKwrzsJxEdSeXdTe4dHBqS5gFdF7J1EOuc+X
Lejhge8GOfEHk7qyV/qk2xWGXJ8bmGDe08v8J4HUmq+ihO8oPvQlk9BrcM9s6usvRuBAclHOgw13
Kiqclq9klEtfceEHjIAOFUiTApd71qycxWqI7yH+z9JS5dKeruLiyFaeVYtMp+x06MzGCkDNORAn
Ae+zSToMQ7jd65bq8pUubOyc375rJN9nrgfnI1Or8jxhdvPP11Hm1dDDSIiWGkgz0npP21oGytyc
/Y9MTd3cEeeqRysdW+Q/y50tfiLzqiSszVOPd6iP9FfJzySyfs+qjuG4fz/pI2NCDyKA/Dn+i3af
bD4UM9bYkVOu6HtgIPJMVmFFcrJwr1u7LaApUoyeOlXy+73HWMFiy74cIPSx8JVFfdCI5ShaeWwa
UjlHOJboMDbPQy+ufixXPCFY6KID+MieU2A4slyQQOZVxDvePjkFNfY11HSgDsTHJj2ciEVW0Oz6
oZ1lzvBMIxubGMtvaqLptlOCdp+E33EQ/TMTdIKs6wIB5pEexolrc+W3ZPmD4eLmypCdbNDF1GPY
oBoas/IsOSzrhhC4MO/+vVa/+vVLXxD0RHOtIwsQU6EW8PPzJjvCqvEmFXk1UPImzAanChTwBjQ5
wlOoFz7Vnk/cNfaZR9M/4f6bF9eI0Fm5vdUEguodAbt52yAP+vmhzRlw7//+6y1/U4PZbg0UjZEn
0f47UfU/fe+SOfqDQu+4mLNDltjt3gFqjygvrMR65KX8ItFbgebwcoxzv5HsJWbMRtosoCCAQZJp
RvbXxovrLU1rrRjJwFUSgQzah2UpbBNG0yrwRVE3f3hlTDFLK2mjWHPZES3xHthzPQB1BaS0GcE3
MnJ3IOolZMQ1wcOVnXn2vgVMSd5naIlyB0qiPaRxVw2H3uUDffo9+/rBXVz0i5MekXjXZgmvHS9j
SdelX66a2R/i5eUIBQRXoCBsqab5HJ5DotjmE6j1wyMl05KXyKKtcTSeFI+dSLZ4Ieb1TJlLN+rE
vU7zB3cIkODE+NZUaLNCYGzHH6/yxIVuu78Sb+N1qXzZcukuaWYqacMi4PC1adtr34ueKzU6SJ3A
Cqpn9ljz2lHibjVhAcMLOLIzHemS0ZSkTEZbcPMuMHWTZtkTfhX5XyXOcZ+fvB0iAlAL35+6Q33p
/n/QEue+sgG+/6Q4n2CRREl1EV8U6c1s0xID2f9uHcKV4/hOS1Q5LuK1KHyjiBPuQtz4UNh7ZVmb
2olCYQQevLk4wsTagSqY3o5EWn6u6vY+TZwj37bdDzy0/4hMkCQlsiaZ9QwD3xbNI7FH2bVybCxe
bZbdSsV4Oo7FQHdxlR/ZjVB7VTcLQT0+NqvnVNfvL33X9sLTW1GKI5lD7OmCKL1xDXMUPuajBejE
nrgL8mtnFNWUQa8WvcQ33lc+Ab974BDc4ewxjBP6OPXeq7egRCH8v996Wmp1i6Stp/XR8/reX7vG
9eEHVl607v7y8kZlSvIsEQw1osRf/huGklJMiuBLWRkpt9tdHGO7F0zbyBs3DeyAs7DbutZWlysX
w3OhkBUDiwpx6o9E1AgTFNklGYvrn2/ab2tamjfvSo6zg1HwclR+kwfq0mQD74P59SX6kvzQ+G1F
NPe4Uo/rp9j9LspjfFpOwUBJwDlkXWdXJxGahuPdisy1F4G2VpFGKkQoN3J4NvzKout8IHOeiTrj
bxl7aUtcZNMfNQ6ngtYuHiw03XoEoWjQOjM9I3FcIlRftsymKd/r0AFm624Q8NR9MK/dOH82Lgpj
3hqlUBG2iSUCr4MorbijVpr0Ub9OMM/CvcA5tUsBBXmyQ6lG4jo0qCDT7rFXbO2ZBVju9Bu7qKSA
kpCqvzl4yice2IUYsW7rc8sqLcFs/HtOmOGzRNX+638Hy7vFB3cGwRR4AgNyhqDZlDXjjM4e7kn8
XdEuoqsVIMArilw/IPXtlbSRdOQ7i7dQlVPqPEv9eRSu4nVlkkWGrwNKTjNmzRWxoGuQWe5j/YOg
xdvfmet9+YBvBER9r/Ugqg8+FibQoTWoWxZCDAqwyL8ckdqCUaJo+b6VWZf+Reh3RsojFsHF3yqb
+Z2lN4FDpG+GpepgtcpwLX2KIUEHP/vFlaCA2JnNF+BYRdW2wMaS+gZRns7GB4ceD5baefiOcLEX
fRVVd/vJD+tyMsXBQXin714gYIeQnZWCyRfMebevgEcJWWomUHZbQGUQSihdDVGMmxvOtIMYe4xn
DN+G7EAK+pTcUtYaupFTV6ddEXkiuGLNEIjYZ1n9CkaCFVLwcjQB0GljCA87LxRuxRWy+kWkJMtS
ifCvoeN+MO5ZqtKEmixv35LRZ+LMIJmuUwCDk5Bme2bVnkjFX6PJbWOnkrjZpKi4Gv22tV17wrE6
Tp5R8Jb9Or5DwbL3rqO26OhgIUtSt7Ih1TsPeuPcdJmSt87SxvqckN5iNWrlSVD+9108yzyVKxdT
mFcPsYU2BenpaYVoF6E4UDgCBxNVWrZqGgl1Ge4hlAvfPGCkUH3Ci99s9h0l77xCl3fVMSG/VzSw
YzSWQq4czohXtnoXCXxtzjO5jqD+PylXBOXsZtv4Du9bD3b8JlRkGDakJXPR9741UgQDhC0zUqc5
nzxlectF1jWE81+GLMOow/Ryd6yPP/sAhs3J+rUAoXS5TqZdSo0AO/+6ipsnVcokKJxsNHtv230H
v2cUMgIqH3dx/ttq/tmZ/CN2nEa8doEFJ9oZf13TVKvzbCmqtJ8QEQDGGXscZNodP80jbS5nK+9Z
pQ7Q4olCnaj1amq3gYKPlreoFuwcOimYIJWGVrh0g1Ssfd0yM9PTK2bgyPT9i9MN7jo757Kd2Mwp
PXN6DWEeNdlywasX0rEYAG7atSMoj4UujDnlYd/fAyS7C5tyaBR3d10Wj0+pSN2HobosTlC8N2wX
peUqaYIuUDyFUjZ0iCDSCYjqoNhdFyOngwA450LE7bNrn/RA+OvyLlSPoargHocE9WIIT/EhiB6T
yCkgUrrAowjphXcRJ0pi4unwbib3zTKJkkJ1bfjBvONUEVfnrZbqb47KpfBIg1jM5MrBA4l/JpYf
sjFRex6kvOFOEwHoGJdeWOuUS+LZqfJ0XN+WtNNfHqkEqlnyJAQb2GfS5mBynBehMpYsbewCvtgY
Ip32W9u+bfP7I5I/cfzSwBKEJW/5PHj9Y+HljDScbrT0m8UHuSWzfdo5dl5gyT4HSiIYTy8aJOaG
eY/LR8gFBuwVrvnZIZAmNr0cwyYavsHHt6n5ZNaz98wHSfMhagD5RamVgnyQR3qQ3caZuJDXuRgx
muPyaLxFTIMWwS+ybkoIQBNhyPH5oCmggQa1C5YmEMNLAsug8XcOeoWE3288UK3QKXqj/YyPNJty
khnv0cboAZUmnYVDhGyrxasq5QKV0KJhbHc5IYWdJ2VmbSsNOLGsJ40geohXJBwnIv1OqGIeLgU/
319GqxLXiQJbwOg7veBVI4vnoWeh8CCQxPnvZWj+kpztdU8VYJK2vAMnfpfkfCRft8PLul8b7Gbv
Qq6azdZW0op+IjD4oXcFOIgakQkIVthHUiik1IP/3U2tGcJibm6ajO4SALxzCbn+RNsYgiDY6oCl
aT/j7cuJfcwf4h5860TO/OB7WBzt/PgDRW5qSVonsLEmcErvs2oAUnJAdVm3e+FH7nI6EhRUHAM4
vpXSU6f1brYxbpI+aV01pZjvnLTWKDtnAUpJqlAYsLPjHRnBwghyh/L1y02GVALDspkGO8o80D+z
rR7g6HUSHm7U+3tCPvG48tCC28m1Uisj8rvp7duWsQJ9YtdwDR0y616LT7rtlMGltj9tEW3xUKMT
dd3OfRC/mb8lWitUz0FaXGMC8H4+uA8+5XxBCg6ARbiCJTjhl8CF3H+rgdHT6qmZ7PWUcI+JNlx2
9iomIZ0j7sv6MQ7zhAZYjz126k3c7ZwSJlLzPUKbLOAbfF760jAjQRA9Uw+U7w+ovlrHzRjmzqbE
cuIzgh9G0YdpuE5HbptXdF9Q9/0XFSIJSxw2xMka0nS2hoFvhwzEHlxHSVfyhtN3eqCpIU9QRg43
jVwyciK0gcVa9UwaaXwu8Qu0eeqGRDIANmb/1Feewyr75/XTPztf0Gb+w3s5Oo5ZmqXjMaukOly3
bB2M18/nqaeMFz6E4CgzFWwDWSdyQmzOmGptkGAswt4f1cjjrzEHEpjU7A1fzulT07kw8NaFA6fo
7sN/JPTBkGYDjSPrD7zq4Dtpe7Laegv9kNiOphGUX3A5JMysWtcIXKh8MwEwjUXBatsWAevMUDKd
/48KKbnI9lmcmob3iAUJn2G6sWsAfL+oJgS07KrUuCSE45FjipYqKXIyfOLh/Vepmte2ShE0FQxO
7CgKKuf0YaVud7WuSbNp9ggoPd5kVv5Dw25hQmgU2X1XE2aMLQ8xo8uFkkuxuKY2ZYY4/Ck+U/jq
S/paW2pSGPFWJrDz45OAVrkDdPW6M8OiVlp2vv7yUl/+OaKk7w7tCiFCMzjJVPYjEKJAKh3Pt505
UPLOp1T3J0GLAJqCCNohNQGixOX9GT3ulkdE+R2niE8h4NemN1ZpC18twUsJ550bZcqpf6vbSCVp
5uWicDwGdqU/1TsR8q8GdSYRXjvCCxciYAW+aRiJTiMokvLhclciIZbrm/PZ0tXkwg+FiuMODh2g
Ehzcrix6jxZurKzFI//nPIcVzY9COgh/3vOeqy3ALjcK52MuzvD1FhZcVAuDBS64PoeO+oIc6a7t
vybkOR1Tz6e+IjfffIVAxzcTH4YSpgYZdyLfyoIx1nifiF5nXYtlPXpcISYzYukg/sRiSd/I08iG
p/IhIHSGYDr3oDSjzfxxhEqFw+6ZL691g+9hFqeS6YokaTFuLTcct0EOdlIOv2tvFSbDNCFUio2C
EndHoCrjFxeZ/4xE3RmfdXUZawgOFD7kj/dUwKXtyptZCdAw907RNd0KNxRnnYkuIBKFUv10p8Ix
wCEj2r+mlQVIFEibRNiWr1MpNI1OGg++KF619FAW8PFXrY/hBhxt7OIJVtiIzcvuAsR3ScGPJ3aY
9GcC5KiMg7R/yG7bcVp9IVcJff6tK91kkpC5rNdeQgCO3OLAsGzXJOVeKCNwQde9jN5BbYETbJRc
I8wTuz/nhiwXGLJhxJTrStBz9E0gfTx94hAXTn4ddHJ19EfWHE/X+NhrltbCXvixRYzJdhn05W5c
D+jN5JgwcRehOZ+Qv5Y6fyuiHFLU/PVsrtZ8GB/M46YdYDsjib2YorY4fewVSDHI1LisbRRVC7qU
W5oL3CNfl2lKgiTHFzYdyjsbDjEO43Blx5sLMAFRHiFAn91dtUsyv16mkLzQ9OGvT+D3OHsR1tml
9tl78O22Iu6kUkxApFQt5cwI4gbQcnHNuLh51FCjqNEmlAoj4mHW1kvccOscO44mIFP2VhclDB3u
BMtrEphjKDMWKWgMp8CPtD3Ek2NnhpclhalPrM9+XcanoF8IlGsdJSCj+1AJfQcekdemm9tB2all
OiuC6NcLR9KTBvOzrEhHXfpl/FTPf5SVY1dBCnJ+XreiwqHyqOzCix7WqM8qsEyo2JzqL6Y/f8cM
nRWcdVavL6xScg8DJgI2bVpl7hQV1wjDgqyWRYC+SWB6zqR1M9XbfDRqBskce/5dk+jbWQoHL4ki
9oWV6VnOUKwuiUbpyFCdggHPxz6pbDvXO2yBQnGjEgcDxMU7LtfCNEDDptSO+EAi2XYY/Z+uVf76
uJlfi2cpDxs0F2OJK4ofzalrCJdk92ljwdScVzL0yyD36ggyDnS67LTyIRavWLXpT2ZUixigBk+/
Km50UW9Zk6m1FHyVyAIBVqTGe4vVFA9wiXYo4Hu3JZU54e7J7Boglt0Sd00Y2IM9TjbjrPYxg9YI
nTYP3S2vRiBmbyawWQ5d1+BeLvf7Yiov3XXW1wMwFKkLC2o7O8+gZhH+zQMYW9z6njrsjNfub0Xk
t28jY+G3YtqI2Ty3vWE9f25W0lvHbALgrOnLO7cQAFt7SHozqU+139SPQ1SSMMMQZGgUVOFedago
FmLvGBxmVTJoXcObhGc1+2IrwTZo/YxJvucQ7SZI670CYWwCw1M4lO+1NxrzaJYdKs3g5bJSpxXd
XO96mXHFiok57wSWshRt2e8i58o2pAtzb5mV7gn44lIBPebKHPWfMEPh5oCPu+vYCwDhsYb4cdkL
7jL2KdHM2MyZPtxwE1tCalnaJDClyjrbvjJmclVXzPWDiVLtKBlL1IpNWwTjbxL5rsI3pt1tzIL4
s9f+2oI92fuRZ6J/EfNTkJar5jQcCQynPYYNeksuaRbLuE7p1poNd0S/Il7rJU2mAztGoVEHXO/P
ey4Iq+RKBh6z//cZD4PNo7tFvsaBPpaHPg9P2BGQzCmPs9/FFICNeuMS+MTJXXhbc7fL9h+P1FSW
wTNlsyqJbYe1goJmKCj2hosSl0QioqyRXctCYE0ydrZ0jeHsKGe2zJa9tzHAm5Pm3sFDsAi5RKE4
P23FMVg2ZzrtjLH/kM+6kn3d3INpSBJjpp8VhUC4sAxUKY40KvcJA0irsUuxx77z6XSwK97hiQVL
mBrmKANscDMsdZeyS9yTd0bjqqhRazOVCCn8wNk9D4DEZDkHIHtMtUEz9A++6oCHfSJiP6D1ZhKU
qMKOdNMW8ICkweADqp+5Ce8zA+/V/OgV7lHay9ecZKvvK6plqC4n455adsBnNkU7RsjBDS5YcM+F
NAUZm3fP8OmnB/OvYQS/JiGkAgkXsdpuvQs0io+4mO4P0FWIusERCKM26/f97gvjx+4pvUE1Xvn0
87SL4ZFMblUDRZ9M7IZEfcF9vZpkDDe1BzB8V9kUB5dqiSOliLVlBZCCmbeEzkOcGhJua2EUIuud
88O3BroyB/OuXpHOD3fCRTPvhkwqnsXD1nd/IC3xtjRAnKkl5Jh96sWYl8yE84B1ZSesXxcV4R0g
jY+vxK3UIxOLnH0qJg/XArcBRpPL+g7g9HJQFGSInugIAZDitaAmFzk0KtGJvjbeRDLI9wMnBije
N7DROO5F8MoEXWD0cgoocxuHHWLZB831WjpSbAO0ReHiXuAXxASOBuHqvnwQlDlNP5CLlqzTPXWQ
V0OGvqNqspCVl6saXKMT2qAr7YoOi9BqyonOOIJzoaeL/Nkd79vYxanoH0VGKmWTJ7/Pqc26sQM7
lpbGN6UCVKHGujxOM+NGjPxgO60v7VVnJBDuYszumvh3O5sN4ewg7c61FV1NkU2atA8YVlEbX279
We62UyWE7MRfBdXeYOWjQnzvdCSIOY6HjDoeiAMOTEqIb7svhDr41kHkreihJoDLLbn1eYF25kfV
YbitU3HbW00oWEg20Ti7qgRiUkPw2+lUBMp9Twy9r7fVxUAoMEaYzVOW8eAQwux7meDxOV8XUr2d
W56fUZTzinl4at7W1g6Zv70TgsHBSGPE+fHnTeqAuO8lM7LUivN3TDQWWysVzpJ9kC1AAK7ANR9S
A8UzbhldRJshT2iNPfAwasX//FcErdo5bw8yGkkYqXQoHQTIdjtXvXwP3i1CokspDM1qKXII1Fpp
0LKp8wdy5NN5aaLN5g1dOdO6i2nlU8gdk/CDOW72wmgIMA9+Bgqg63BDFlOvyEUV8KiCux54RzBR
cdvA99W321VheQ3UIQMMmlBWN7X+o5i/VrTbH5iY6LVrLHggPFvBjSS98EmRXTMn+nGVCtRuFylx
cRzfqXY20kTyUN/XhCG1wAyvX6rdDoyfTrqh8nXuNHId2IbrXn31JEzmBUuUmI5eB/7gLksVyr57
TXac2XQKbX7x86VMAUd7Ozpa4CpWahgIzfxlop1FgFsDvrMRI5J5quYD+i3YlWfVoHFsOT5Ld1Fc
PxmzSgxq46EvjsDJjBgD83K16VZ45nMZKy/iRS8ELpqaUG1dN50nrK5QZHxArWZrbD0gJudQ4A4L
td9Q7mDNgGP4wmGQaeg1DOPpoc81w5Y21+8X2ITI9aqa+xq1yYtl/imMAq0knScRiUb3kF5q/P2X
zHbDbzEF9jAwLG+GG1HJ2lt/jF+ZdOIcmsuBWfB/1K9F8QF3Vf/dxVT6Pc1lQppRGuyf+xUo4YBp
kaG8TyjHYnx24eCAn9Fapl8hYwL+52FqBEC2x71UShKLBRjo3OaXpHVh7LsF7rVeTjl4xU+G7Amf
km9Sa7l6s9ERrcaqIyCCYLK/p+Nl7jGFe1dpw/U7ZaoXAnfobJtvuXMoIfa16S9KQS6lvAy71ed1
NCGiwo4jWuFI1eIodaofHx/1PTTRu27s3/9geRwaqmUooHu8UEoMLxPLx4LWpGt1GN97jzgz8gsz
OP3NdOMQMzpk9fAbYMnc1G425W/6z2x215hPJenYxmVXlQWbhcLTXRdH8pQSkPycysnESKyexF5i
htLv6mlnFB2LqytdejoH2qQ2N4/5C0ot/BVxQkcFYiCZCdkQCloO/B2DDVz7THxrQ1Us3e0OXZuW
6b1p1ehJyIP7DZ6Y5jsEG7ucP7N1MC4IYLJIGb3BtSNF5CW13VAT0UXlqOP7mx/fvgOwj0DYUmY1
jdqBj5/HP3lKfBR3VplT2bmn1Cxa8NnmOgWjELnYqyVrM2SGtMq53C50g2KBpMaeSJrA4Kp4eSr3
ca7Zx5w3fdvRGswbPh2nEiRKQ24HP46gQClydDYO69lNPnZIJqIOcQQvAfKeqgboHiGwHDw3uEEg
b33Nxf5cmGQd2k9f3pTIQd6U4xXSK/BPSVpS6TH/+v6s8OaZtr/GZC/pstSo2JAkpjm6rrXU/+Hk
a8VVjsjZ445pk+qtyCW/gP6gr8pRnecykg2OJnvSZ3aIumYoiUKfjgbSyCwZDqudAjWKwo7EuxK1
rgyk+tL/mm6qzOolZzG1C4U8FEa9HEZvCHpsn9ndW8aLJx+l58sGSweiagZQ5UB7cihZK00SyCPP
3sR8HwGZwaVfjAl/qofnKhW5nXq5lzpNJa7w8nmouOgoZvFeS4hiqPGa7QfZfZUXzFa2BN3YJS84
RRjdEec2vpmzihVr7CtNBn/0Xch5ZGCFA/7hg/LtJKK8U7DUa/Ofd05zt9rT+lyEpHX/OEphVIIe
npQIR8kqTZccsaBx1nwxPLNhrYlMC/pIDFlscrzXMsMIDrR2AcZ4nIq7dAJs1XyERp10QiprULwC
H+IsJcwjBN/aalFclv2Wy74hywByEdZc2fWgqTB61A3JcvxiIuMa1ljHZvZ5OEobEpVUL+P5ON9E
2sAT3uTeoKU+l4KJnqTQ030sdRH3KYwlg3n7zQdhi/QRb3Zq/VedxGfAdzSaXj6qGP7/0mc/N2OM
y8RKu+P6fsMxAvGg2FRw/NdwDE043ZLa6bhoEdo3fayPxyqMeJbfYfMCoBXNga9w9eX/PxmQ3Fpt
i8IHSzoJLFXjc1AVGHvB0ZjMWzMJaUpFpDJQZ1B2ld/OytDRKpwHlex/3cedAOSteFH5vfW8ZcDc
nvNr1qHrfAn/i+NJ7+KnMTfAI1SMVUsK9JMUDGZcK23yVzp5Xm6djnU/bzhFjxGD6wS7numxnghd
NkjefFXemTzODxXZHoXyxu3k/uVm4w1cAiF/OtVcbeDQc+GIdPIPNb5YJNm/DU1e0z4DZVsdoxrb
LCEJ7A8VEB6PQNTj57FjVPpMTYrBZ1v0mCzJ3bPLjCAEVgvWknwKoqCxEqnqc253vpyK4kUE/FXg
kJO5ej0JdFBroJyMKrulzb2ilDCYX3X3ubDJZTNTGZQyze/XI1ONSEQz9RryYe7YtZqbjeSgDPwx
/dxJk/YBwgbXHoZhXOEgwUuWBBVe/JBigBHrQwz8xeDuaZs9jSi9gZ8Quoa4zZFbcCpeG2N7X2mx
yqPiULEoaLLrNC4NFiMzaDx7zs+0aiOE++4/KjspNumBIZ32V3OA1VSJZ+IvW5gICNKp2FgT9mvr
z46FKpz5fzhoXIxuiBfdqIPNz8I6c4wm/nCTqvqbjfvBhHxjWAqwAXIzYUzLgzDK4sF1/zL+7ZqS
9ALhE7S7clMKSdHsOVVqjHbHx5KqXiAyRt4wq5sIHTXAChTirWmpySKjUj0zC8w4XITbdCTKLKiA
7pdPHUPKjLkowJyHpQeOEZ9J91bDaRybylmaZ8fXtMNVzJGp6e/qwXwbxU0HA+QkwAOCbI0xZ4OV
8m2HTEUdjwRQoZEWTMRJMC42HA0Cy43f+KBQWZGZ+7KrXvN3AKKDhMHV1NRJDADy5iY47X7/tOc+
PC9MVsaKObr5DsPWGQeLaH5hYaGHxsgmHzGyS08eYARhyBNWP694cFT5DARBazVbpPZfzzgELRjY
kYCFCBnj5DcXCJyhTitwyg3cFD5EPEhH+Tmh0CIzxkxqdxRErdLrHo4R7Pqygd9mVBVAY5yxmp45
bBSVQfTd00D6JNrkWLq/Ivz2F34MvsArlpe8tSwJRUYjX93S4hxz3C74ZPV2XgSYpSrqAu4GbQ89
Mpt80V3PQr0xo2CFE94PrL4JqvXlHcdEDszmRSjcbCEHwlDAX1NsXq2WXnPU1FBNYC+CX9YlHnuY
v+NSKywYmPh7yAsQqljcBC/IMMO8S9l7pIW0c9eSkOSKVapymdrICsxybM9YW4lqERFrnrjH72Dh
Yi/XwK863tyWxjxalj2HdJg1P+Wn/3rLB/rGBHW61SAil26dTEt0OdSTHxzgvBmkws0DgAbMrqLz
e/uQDrBRr3a+fZO430Z2qhFm3dxulrL6Q4Dl6hgeTO/A3C3Vnn0MKxDyfBFRHL6mwxTSHWkzFUWE
W8vBR0z+nfBHzxObSNky2Lz0kou9jrSKXKRMpRR9mNhFHU+IB58Wa8aw6/00CmCJ0HqIg5bOs2Rx
AeaHwQxooat3so5bYPoxCvvc0mGbU8TQOZR9E4Jvj5P+vJas5nxbhAVpQw2HZ7fhk81X5QXVLSMp
lIOdYsOwaoWBMqo3jomwvBMuG7TApoBDgUyJ3Tjs5onTTj3E8qBvJ7g9JbQsJA2yUaaUCbyGzROp
cpuYEheKVHovMZFdUHw2jSnN0PNGgszLfVdZDTsy5Uu51uuKeGTrvIW0i2nn84ItgYhHLO9aOOCa
pIRQ+FlmIfXFHad3kZLTMY8+kM4bRX8VW1vJncDtIRzgJLJSyH+ikieRoGlGQ6+QYohF1imAjvAa
z69ot8Ma6gBIeANX5mqOBwTpbFpdHs1htWvlk7SIxRuiujvIuIoW3KuXrAQ+WEkBQHDg18J3sjYj
rkRFMOuCHcU7FSccxQbXwSPSbGdB1d0m9WMPACtIB0H0y8htarejhMS11KDHJtpq64DpyOd26J2D
68c7/zl/62SL5/jw1+lvhQC5OVTk9G/78fo62oVExNcgM+sKW7aJrOrygDRY9xjxtmHEtvD5w9me
zPckZFiL3FehgRvOjq/LGCTF0dxOc3g2BbcA6szVJK7xFvGYCAR1YGWvmsuqUzIhr9XL29tpbGeI
3ZMlNiagDADNEe1EX6AkXQvfYQ5Tdm2s8aO1A5HwIJN762HToY3G4SvB31nudzqLiNDzH5kqJD7D
22rWO41LmMNR/xK+rzuo0Fyz6NxUdxARo1/s51winWJoI0AvzPQQLJJrCsxVmg1yRyY1mcUc+rEz
G3Nh8Ei1fgEHFhGnvNpI2HbBp6S9jGWzmTxt8mCnm55rJBi7kbD1c0Dc/pxNRPphIhvOce53TxL8
aTtYwGzShxCNDG67NheQ50f37+qDTfrc3YY2XIDiNdagCk8YDKBzmyCsVFnjv/3G6NXIcUgEvrI9
grcnoHnwU7kvB+ABRMC4K/5MuayqY5g6Oi+iwMY19Xx7zIuuoAkyMGX6zI10EqWlejDnT5nCeuKM
LbM6F9RV+tAm4PIW1LBfeBLKTHXaNzVFYeNTkSyq1cuEzYWOkDHFzSA2HIfliIA1JUFrOdwbwDd3
YeRzwgygI2KqRCswBpnOqQn2icAJu04pBJpmn39JGzdcxthiR8awXWIWxmGRqsJir2A6wMK0wBJM
9pDb0pT0R/sCsFL+bfUeY9CaLukM8xaT8mc/TMtL6z2c9mRzw7cEzG4xtvdn+5gMOv44rRpRL8J0
v+ukLCZW69qEFDM3h6fjjyuzcAdYMUTJflnxzSFWhkqnJ0H7DHcY8QfoxyEaGfJkxndCWO9YbFZF
/Nevyd2uo+gWOvm2dCAVyQv5h0fTIn+tjVpAgP1pQJ2OStz6nmY8ratGUYpI6NTrpSWoE59iShW2
FX6GvKig4nexgcj2pk9z1Of0Rc3r9BPBwRZWSYpTAJK0mJj3hoWvbgCRaxjOyF4rUIed7QjsOpy9
i0dNyYUtXenBMomIBbQjEr9JxTMwhQ6KzsMsESHojUiVxanAqWzmGOX1OQXPgfnO/NkCm0CIEaku
JSaX7ouaYjJ1CjcvQPnwYOiUgK7PNozeGwmyb5vqf3zVcvS4850n9f+j+C41KJA/3KRG+IzweTqw
IlQsGQNJCygVK3IHBk1e+Flg7uC62H/RNKVhYFevgYl50K4TDHBHbLzLRDKJiktCmHoTGWwh1+wo
DjgMEw+ojzDZ/VLeLOYxgfGEF6vQ4FgUiG0Utl3aVSez83pHcBqtBD/pWR3MoziNcSPp8NwO03IF
D6ycncRVF9zKFC+IWYn/JlqOLBRPNyljrV8LHbeOgLeQka9CR97CcG7KQjvCP218++3QRVhxrZ+5
Vd0f3DbgbN8Yzskj5ZZ52cX9M75eIxTQ2PgLgrQfmPmrEJmfZL8pIAyrddMBQMvUxaZdh2uvAciC
0Q01AudfIBoRAxUWiMrDfq2nOrGvlcgsLhKTC6C7fBdqZYetdzCpRsMI1wc2kkDK7na3t7TPYcde
dvPZ9RaX5EBRPooqQzot4Df1FO3UjYuIiZXvtgc2JwgGypmhVaivH9tq/oYNVPuzSU6mbbt8ZzqZ
E+jQkimSkrCDaMFj9FtYj0ZogGrcZxJmRb6G9FV+uC7cQxAdXyEO9aX6rhrrNzQf3IDbgkjE+sgD
cnDWpuhdVKX1PDfAybfD4o20jHjPjU3Qozu3nj7yBg3KY4ENhQWEzBo9PGU6su0MH5gaz1WtZedZ
4kf9v98sSKjkgLSAJozncsewWzXTGGp+rDq6J3SRGyfHetryxmZ135oLnvTmi6haGOf7LURuJYxm
vg4EdqUkMHoHHD+5VxyNxOygiqGy1NP2GNHxTKjKMcE5mzxvNNFiLbne7XpCsDxMG53ABT7DqCaH
ybE2wRYIzPiZBmNp6mh3XK5KqqJOHC+C76Wug88KBxVbTVkJyoPAe9aXN0Um2/NQJRzX2eDguPI+
XMOB+y2fBzo2WGj7JIhTaw2yp9iNweJdXYiAC3BbUVnmVzwjS0YuwaHE65GjDbymGo0cUUhMsX6F
6bb/W4NuH5iiryNSJ1f+FrJdLfSOB7hVOXifUYegqfYLH1KrG7bVodEBZjwac3TUXVcoB/lpxvXm
1jnVJDN3EgiOPYgSvYYCXNkmhV6h6tWmOnUE7y18JtENz1PedmJUdElpPwkiU28j66PSjljfJaCr
J8LJI1aB7fphipXK8g7BH7O8zhd0IHY0Nzz05T0DIGzDxIw8Jk9HsCIohbeXdSAk1SY6huaUJr2z
agQyIADyBerreIImIEnCN9/W/dMznRN6nfu+6YXBXzFGMwWVFUNbLmZclacov2L5vEsDjxXUUJEL
hA6ejjKoSF2qSTzPLjf3aR/Rfolr1NoW8O1rfiBhgN/WBGfSYqX5PGfaFw0mSmFzM1mPiFY3eb2W
BktWK+8i6I8lbgHs+bnrt7PyfmGMbd3OW0t8DDLiuzPoh96Qx+8YNqhx/ptd6pOZnn0GrLSvvcth
ejyLDzMTK4S52dAOWT72dDxFlbOSqRPdrwHo22eB84ATOCh1OVYtaTCjiLw4Wnu0VcPTT9IBgwiK
vTgW9RVxLRbUsVP/qHDb1agSjbj05C3ebXWddttjYQqkk4s/7jNudSHzHUSEEbytmnuVhTZK7HUi
7i39nJI8txpDYjGOAPoAkxmt+VX+HPe5gwAzckZwTWpSCMA8RM/WEdvoxQMgBdaQJDYyP3dcNOpl
DY0y9XdAcj41m+z9C4bdcsryrB3/JCBWUPLplgz3yHgBKqcN+03O93Ob8ouOmher7UOi23IEyvvG
qlFYOmJUqhbKk0nI6CpwatDU35rKFPIlp8PgqpqNplxyabB/NiSh1Luo2kNr0fpog4GBNkwH/NVM
WsHWPIKAsoI1/oDk4Y5ZPXfjdrJjxIsck7lvNz98PyGcYwHei0VLDkZ/LIL3CCkf70JG4v3iaKVf
ij4Z5ctwer+52H5XhRG87gEiAXPkN7KKfPGclkLlIp/eQ1HkpYZpXBZgPoKGWSYCQ/58QLKKtvtD
A9LrBNYAJHmSkRAbq476TuQInGvIX3/nLh5TkHWFw3m51nD2dazX4eR69FYxmyXDrRkPs5ado3WN
VwHxOgZakmzx+3oOj6YLkWCuwA2KHDAr9LBcdyq/n4QxaCc2Fkauhrx/mvNsYZNEtO6+BUyBvDiV
b1GEJU7l20NsSn3GVSCFTB+pldm5BfNlt8o+MAjJa6mgt8r2mHAvGv+viNYj5gixDjmvQS7+ORMA
bINug+Tr8e4Zd5mAhLuv9/ILFy9hmyMgTDJDnz/iPhHF0v8ay8/DkItPAUwVNFF140GpeirbZu0K
+cb2EmZWDF71UhIRjd9ulUmfFpIjLQIQvSBcTiWPDHekQUFLGUP5ICiZRrFORHw9qMwzP9I6EENQ
H9n5lGKRX0IEtEAGLsp3ujKly4vpYSPT7mOOxBBd9/GMVYXIGacPBlETOmilzbKzqtFuMTubINew
qpN+YkJeDdNzHKe1tGW4m3C++JJyYulcDAJ784JnPqtgBG7ZDpsYaWzUTRtTQVOw4YiStqUD2zj4
0xW2P5AOJR89qVNNNx3SdaEvv8sPpxS15SFwYr5J4povCaPLyDXNcAiTtCD9as8285B41lvzqpDz
BO8eH7aahIFa0nc+G/iN1om0+NJ5jPRIC3SZW3hcF8reaF0dImnSmM3UCFJSHQI3hFK7OTQe08ra
etllCvO2ioqhSj29EbGNNV1Lm24WUe0ziN7iSJnbJHrGvHp05iouA9girXOVvrF6ff+LUowzH/V1
ORG5RzJAWF4R/yOILWxWaY/Q7RHeszI1AT086UVl+HD250y62IIN0wpWDh/7CbJj5EZXg5CC2zxw
2PQjvywuhVF5Q29iYdpPbxCjg5+4Vr6bRO9jvMan2naBZDsk74HB51XucfFT8VTkAF4w2VJflKZB
Fg3/QtmNGXXJS18iZ8BjRpV2dFQ9BpdS0Xls901Ew2aEj7HY9rB6ODZYEz7/f1DEgarLI9JcYIcK
9TDKnNGL8gRx+5imb7ALF9mMIDoRobL8r6yEEa1iJ5m0ID3Qcrb88fSeQZSgT4Zov1rn5sQLJDkz
bThZXOCNLq/DoejmZgOjRg/p66qAXrBwNLQJtAxWA6OFn7HRxYCfxCCTl8IsIm6PIhCEsc+Rf3vr
VM7zNKMJS4Zoc+9EjrdX6JejO0xPrAbrxLDmyNOxKGw8RVmBF/+E8OLm68wICc220qZJe59VmrB9
UGYrssS5LnAiu+kHj0RB/RomVcYr1H5H1EbMkdC02g07eyI72KjfW76iGOLmjm5xmNoO8xL7OuGE
DlBT627gUf01nNpkYDPWD/Fg+y7Y/v/Yu3TdtbyGMdJyGD64TpuvqslLCoQmP4yYwpq89wsognWp
/YS7iabrzj5AorTfPiYuFkgPuKA+jQ3xZm2Kyjl2hGs6rXfHlWPlkqOSsOYTKISL4ZsghFltJdHs
lz8sHELFFjaECjjh262TZozfVSRD9cbQb0XsuwuYVed+0Rv6vyubR7w/68Zt8hdQEvn8/8YRGpSF
mu1RbgAwEEvvrlIVy3GYRFplZTUlJZk3rpq+J1sHsDRCJRIR+Ekk/kwyEWVaJiOieNLp/FKpKVi6
CmZOEO2vg/Ilfz/5evK89rlWyFKkCVUBcBGEIO2FYiU99aXbPerKv+LViGYYouyd47b30nV3r6jL
3Sv/932bG4lXQZh+VlG3i33LWA3OjyuFTv+SKolhSUiyfLEPX51wfS6tWrad+8hIzEZX6N3PIT0k
NxwM/iwNDLWQ2Fy0KhBzRskVsL+XHv5fsfbPDqanTb1RJfx3p9cAMvGMsbwYzcNsDvAofunkgt2k
zOMDazyq9dTXTDCOGBD1NAcORKQjnAEYZHLcuovcJwnFBbUf9jW5OmY9+i7j2RvfJ912yX/+fWNy
nDip+49T6qiOw5+O5JHG71D36zWA8qb06EWp/2q+5msdmQrQ6Xl4Nae1+kLvQeMRHH8+QHP1yTeu
pS3MkYHJH55ti60rKfJS20eezvICctexeYWSPMVQ0pzp/NZgOpejhjFcj0nMFKawzRF8oV6tdJP4
wOAJsKvl7kMGzHTAVl4YPuaorsKLLcnbIUxWBrc4DsIxCzOGQ+SddVGknhT2jeTe2B/ifbWlOjjg
tn2JHq1MbqAcBZX3Zftmjib7vHofSJShZSoW9zeOIGJHgStfuFTEhl07QqlluLOtJYUUdrGFZhaq
i9HKogNIBrZGua2+b1KpBF0VaxIyIPAGKB3OB3l3f/pfoZmMRqOcJJ0NUMi0mIlh4I4baaKUyIlq
VgQ6+vQrBPUu83Aeoev2FoDZA2RvH1ySuQEXHRH6tSzVNIXKEU61JiCxTdyjmImdibKCO3H8PbGp
PlYREuO6srZqkt0YQ62SirbZdTTdx4c8XEiEaCQfZBXR4ek0I58QqoWZEOMppMDBwutcDFdePUor
WmdQefoEO5rBB9ulZeNpYFWA4rHoNSljMy22Qq0/qDKSwhQuQGwyewV1JpjVTrp6lZ1wKf3SNOfc
bFRMI1zZdj1KWEjd9UdT+nTwRlaxcE5Idx+5Ik/daIqDpnp+8Hg/6QHTMbtffET5GPJOOlpjOb81
oUYPrU+Bt6pj+RnJr5KzfYFKLC6LJQMbZXRpTtOyelG8FBqK/lWLAie/3LBBgmN4egW/k4GO4olB
j3Sg0MLkjlgVUqNYbuzqihUjRF2tlHdoA3vcUtB+2Ij/X1LSYvykeFXQwM+nwe19TZUTioJy6E6W
IGiKHBbNIuwSn/UiZQtA2WBj5HXZWvgTIbQD1yGX4iqvqSSaumBBsfJoNe29C0aJKbWjpQLHudxL
V+2paCzgMzZfMskybskj7rJFN9HoaakheNMVgOneveiX5+VrD8lQEhswYCfNgOyf0gqoSXma1WlG
pegS6Wg02S19Cme6XAADxB/Qgioi8sjtNtfuC2pwwO+t8FffgFA5yqsOOwW9GwLUA6hbxKgAGnoJ
BpzooVIft5yie7xZXmqJz+lHgCVuph6kKFliXVYvDJjCArjREKacT1iYnx/2AKdRQqLc6STsJbvW
27idecADLDOkM6nHszqw5WtvT/t+SOwX8CAmwm4O3w/acS1BdID4+17gtPbJufYn/+xrk3S5DYtM
W0lxDQ8ijTyMbhatZr6kVQMxm4jTKelwz8M4+piTGIOaXecnV/wJ0wWWF09/kJbtJMXSgYAhZ+7c
en3A2+w9zIQcmPHek1x1ERC1wpILVhG2RgTyDbg6bdataCDGd1mPk8mWcmP3zDcijE8hQGo8zdo/
RLYHmgWeEhr4TxNjbr4exnQZ2/21Z9jgYyqXlfTb3hXpzRhr5/EMDpRkacxLd76p3FUnNaMQGJV+
DCWV5z7R7g0modq8V8WDWuTn/rO7dwk0G5A7Zaye19183U178Zds5jFZruI3H84jkR5BU4SN9JtH
zWw05cngg7qbsFgd5LhmOEsCPaZBAr2G9M7k7DZQpG+Qzvz79KdeIUKFt/SFSVRH8/YcbOOprHro
cTRyS4D/uooSN9AOJuNnDJOZD5XuTRg9g3nmmBj48aWU6It9TxvF8fRA9Ot78GqnYdxI/pGd10TZ
JlIt1550nVybpEWCI6n8VXMVTVeAfTfsV/0Y11YiTTCs8zwB27G2hnLDG4DqxEggjBH+h6UUpuXs
+dAyJ6CJ6GgYtsOpLi2UXLJggTN5pLUy3d/Quzv1ImgnthzDd4+ETUEXBKvokrSmkF5XtNAva3RN
nHO2DEHfy2I/20qCmPWppcolF30GwcPNW/HLVZOs7d3nx5UgLmhWifgJNQs7UojhRiglXsGwL5Az
vwoYcVSuI/8APZZwIjvDADEDNzLl1iwZDs01cKab1O+vw5Y1Aoe3zzAm5u/PYngnIiVW/r+ZtQ2f
9JTFWt96OofveaWMnkJROv+m3ZkvyaoRMo+hz8aWCBrOzwH88s7Evo21bczA5iuYiSiC2HBW7EP4
bNXCBYD8kl8y6B5yYFujxHhJ1gbgzxR54zM2oslyCX4aMRq44pjGTZTbWTpTRoCa7j5hL1+EUGpq
SXgvt5Zqfn+qZ2HiNGKchVuUHTW/yp1PoNmKnQv3gF0NEGXEbRzd7hgxQUAi+QuJ6uyIWhWaSINB
XsPbB/hyfrC1YhSH7RF/wJnkhq5ygs8TAFdXeLwC8Jkeh+xOAm21izGqn3rC4o74VTQIrwD6MPHs
9HswQ46T8rGxDK0orDo+KmmiJBuUvLfzWXd/RtXi5kFF5M3eO8rPIOypkKfdaqtB1BgYlKNnkbOB
v6vOAU8mp3LwLsqJx1E1qaw6aUqVLA1oMGsenL1SSC/jRTRxcW6jxNyhlSNM1WVUWmpbW9HL2/6v
kNks2qADLfbh3XafzOIt6EVjYKeS8hLgJTyR+uEZoQ7InWDcG0B8YdlMwyVZ5JWPrRZ5trOce3N5
s03QGlkkmZdHabDyPI5bRF7xH3rm7dPPszvhWRFbKv9N4WhpYNvYzYv0TDMyZRu3e0Ba93onsZuo
TNjxJrZpY16rVXM2SHAHKw3DnpVT4Uaqlr/vPc45KQu1A+JrZ/WfsgtirDsnHrPWdE/iNMany8GE
aQHqSE9DyKPQNHrXI6kx2RIIWUa8Ql6SbD8LSBaZP7JwIiyy2u9orZVx4f6Y30csO1k0fJSGk7pc
Bx+WjygIzPlZ9kEILDM+hq7yR0+hSTZqbu58sysffsDEMor0yGfUFpIUiwFng9gHj5Gnb5Z5LMSX
6bUOzEVLwsJTuEfyoezDxhUp8HvqwyEVBz2zCfU51hlAK6p8CvN+Z3BRG0tCrYEI8FdAnKbmQXkh
W7zzfHXez7VatjuHxu/pztFzngKvyYZ36W82cba04aE27QX0nXJq+zfdfu9JBnn6qT+HP3NGD3xK
n5TNxsV343/dC4neQDs/TEsJC2l/dHYsKuNgMrli+eN+TqflWZJGc+LFX5sZ6GiEi3S977rH08aj
pHasMkQo/ydF/xTlII0xQRnnLy6yxrmBJNOFKJnEXIuZotsuGBE3/PjqPLFCfbUd+EUWMeX0d+4t
DMPdfQTujhvz//EADM7YGObiFHqb0W+myWaS8RqtNCv7XQbsdrcOMucjG2l2/ynPOG7PULzNhIgj
fAuNpZne0FQor9FdLWy3uJygGjvJpS4GhREz63/cQwjxlbBfcEmJ67fLZDUrW4KE384tYlEiUaem
ecjGn1XdkXg4m6I/3vyUVTdx3m4KoebPbeakI00unT23GBb3xxSW0TIiOpkTRw2uoMUEXT0CU1qd
UhP8QRTuT9OLdzhHp+vZaKOYO5KGcnMgUygl6bc/tyP+ROSdTwF3rvH7BlZRMqFs6mQs+lLHvPzl
EWacURLv5g0zc+TyX8xHeQt8ZmzU+WIYpH47fPDJ/iKhToMKyvph7FwXh7mA8fUgNw8pabVLY2E5
gz1+ZoOVW1+0QoCeR37xyK+V7tEgzBg9u7mpdopbOAK2fe7UPGgjHTsYVDCNOsbLk9VCXAjHsaCf
RzisMZ1YLwTuXpgfGVPFU4ZQP2UZSfUCAUOWnlRSI3pWStvK6NUP3xmAbrn1A8iVlRByfw4wOOBI
14UbBRSZRvbjQO0aGvoc6w/U4sAva5HMaeIIfo1E2lFiB1FLhqlbvAwshJZD0Hh2Tza+ugdMeqId
4QAgyvVnA8TK3rei1nyCxo/YWwvMDpiAqJ/OUL56mhXCUYvswTGyOQ7dI2GgTsOJEiOe6h49nVuR
Il30lsxGzoYgk0lb1tuSrbjfD5eJhxdFqwQoLDE8dSe7DtoiBt+qhcgOa+/EfO+CKF2HxUJZf3pq
Jp9l9VpcZ1CCKIQcp6W6f/Qcb5uSdWiCCfcAq8uMh1ei2q8ZInVxKEzwZwFWuQgGl602PWZ5LGmg
/Exh3ZmP1pOvXZITQtlvn9Uz0HKzzQLkBgD4TceHmyn5NTpyq5RUoPR7n8TtwXGBRcEkLYrFE1Ws
sYFkiEunV09wZ0oiflhmPQNymSxpKxB86Ii1mEUlsVNiDSSlgnYxBHmPtcOXvpo9GmieJID7Se93
85+ZLSLhqdfcZNSj1jmivV/FDIBorDprjTE3P+7Qy2LPQ0+29eCzEeSbTH4fsAsJ+JYyBysohM8F
cxZjVwmIH5vqKwEjvoiQCjaim0sBcQuW/hSOMscUYplnCrcMUOZl0BivoKl/hOk4gD+FXX+WA+50
r5UlzyFPdMhFSIv5EY9ZjAiJY510JFdAKSItA0RH07gERaXlaOdi/io3lcgMdyEhkGRYVifcc0cz
+rwa34Vn4+j4neRmPGsblbf7beRl/0hDg+Cq4BYrSPrI7BAW3hyunW2Oxyy9uZIY3Qhr0G+XJx0X
f0zOPofJj2WwVAVbDjUMUl5lEDRVeZnuAwgGW/5Ig1rI3WoNAalnl7nfVJZgzo738a+Ctqge0NFa
cwI+Tz9Cx9TVJc1KEm5RvCcsDD8aMk2UizveHe/c61WEp9xvH6ml5ekDjzHaFinFfaJc2v8A9Fc/
0nNmUtifnzGARaSpIhso0u/o4+JrWphELykCghVrq8yf9e04agrrs8VK9S/rz6tE7ZSG7qXaWCH6
f9kRD/6npt8CL0h6olcs392RMZB5ryW42UT7MWCb/Nj9lYCqTPXzAp5YlX41gkkV/aOC5dgrOmLj
eX4yEuqOGW3NEy61o03FPDzcBr6DJr7p7dOSKpnxyXO/1P6t2YbLQjM5jtjbqSKbYjzP5UPRAfI1
Msxm99aEP/oMdrvCxSVnPBCp2wkIpIOw5O9tWvnFeVnI30WrIFDbSzDP6f8NbAuanc3EH5sNTkQW
0yMC5V3qa/L1+n3QTCTRP2A9esnqeqxb4G58aEBxWbwTDB2Ruel/BazyPMWlIPGwaNcf1b4RYXC7
bQQp8HZDrMOaQnsv7pubJ2afPryOg/IuUVHYT3LTi9U/HDnIxU2v4AgQkylHAMpjLTt7E1pg81ja
0FH16qW5fkHtLbS7jcDYpCbf7+f5KM+59ZKHEB9begVMLdSZHzgbL2LdXnZQe8qLfxrke1jIEk1a
uEABJlYw+dXHv/3rxXf35wPmHT5Iluq6yVSOWgfsfplkZPntMIkr53TVXk5ZnbNF514IcXRlETZb
MkFcKmT7/O8am6yZ4XqwRWMWWkWzyeMCIh3EVTcyvTd4GnEC4VHV/d7p0rqnuhGVBgtc1+vd8OSj
sY1GG82/MBYp/GxH9irIdNLMqA5jtaBHpOpK/qo4i3U+UjvOikYir6tvhxRTr/Lh091VA7pmme4/
FLbgE7+coTcANeCKeYpJh15wzIRgoKI0xC92cJidpXjgejfig617KxKFrsLvRWWoQl58a+pUhAK3
qFBhZ9fTL7/ZcElz3PES5TeaLx4yj+R2iRNbf7F7kNEUjlFsoZ6KCKU37oaDUfuvy4aw42lqUuH9
e9C3wH79V8Qd3kSOTPieff+67B78RDpReJsUe0ChWS4xQAg2FAPoNDrBUdXAc82yutf/FFzfpuLY
tQ+RrECX3XL0uWtnuiSdRN9XjVniZrnWCQFegMFZhf/xeoS27YFs2kud0pz6q5fWFRsz4dUh3xud
VlkL/0+e3vp7gxhl3zaapS1L/cE3TiRx7Mz8pjVTmv2sEzDuerixw3Q3M7AzNgheEWwJDduOVpzd
Ezdcqv/EAixZctO/Hq5oXt9xn1/bphTrdI5XLKJESdpXQBrYqaAXLkuJsy6+JAflsIiJwYkwAzjY
TxPybl9AgrMtX/cB+Eo7FYt2S14168GYMmi5lEswBQrXyJMALZu7N/i3VYt2cXsonNT0WCicO9rm
trSMPCEvNKYpWpG46CO1vjYZ+pA4noRQLvgCu4Bau1pvxDAuPl4SU4qfylonUiqb/enmO0RrwiWh
7rrZaqDti6iixrCQnnXxz9JC8cZ2s/mowL/zT15om69XaFQHjy0dS1m0dt/pbr13Oz61P/LoNhNF
2Y1W7NbgcIbfv6mVcU3KqM7Ekj42Iz/20cSHpA73TFCnYYq8CICLz69eHojefC8RcrMWLibYeo2m
r46X14gJb2LY4YoOyjTiOM2VP8qdrR631Gu3Afg4AXgvlHxyltGOA4z9UADqRqj306jUilEJzwcZ
n2ChsTQXD8Pwz842jlc0MKblk8weNlsy6R2Y0j+J44ihBP73xQtQqVw61LOB6ngxAYqMtYEiW4U9
a46nr1Uq9/QUWdRD78leUedRzYn9Hp/QNrL79e/bjBMhCixndrnMpDVLIklDz5mqJUUUICxAzcqk
ecFdZuhY5WeHQmud7ahfkRpMRh2wClt9QhuTNSfJ2ewDNVWFZ5YM4/s7ND7zUJz2DDiEJngl2zW7
hZmzob1WreAARB2avcCCiCZgZHJnnIv8HPwwmbsxvBd1GLEoYC9TeDc5ZpoIgIvKb0Yi1ohEMriW
VO9NbndY8TDiz6rULg2h3RxEPJa93zbhBGOO7bFG28KUD7EVoxNWM98NS/2y6yDDsGsPn3omOvrQ
6lwv2k282uwZ+TR77T0bHPwhEMaJLuuRH9J7ln+xiiXHhvJtvsZZK5DmTAei7gtiDtQb8WMP2Leq
XL2Hw1w7B4fGhj6v/623DUO2O8EmLjieLSwyF/sQb15nXZlGRoFCeDScfnjLQYz838mKf+IXzC9F
pTp2a9kRz7e/i7Pk1EXwTBH0t0mQz8rCGxkkQFAvanUF/2gQ7HlCKYggYxLpb3g5lk/1EGfyklCO
XrXBLWxtP2NebWB3qT1Eniy/ZXOfXQKGgQcRoNzwZr5EoP2PAsfRexD9uiKUIXiUSztMBFzbMfrs
tH5ya+gPx5wgqT6A5TazPaQhqXVpW+UDGVUfCIoKQGaNL+0iwaRksaKWnwRfjinJV7P/KOgjMMiT
aZ5OXqJBKGuWPethAStVZXI9XOyWicT9OS9FP3Ggnw1XPU3gqeULAsbXRNLU7ogdPEkKBctGyZgi
eGKLyKv4alJfDhnDBQ+24giuM8uRXw/t34ssnpukGaf6qDG5Foskn3bLeCJbk0GJZtA/LnykN/gU
hAqLzsrxoQLr5ZFRyih1+vjpxO9191M3X76B8mVno/LVgrgT0ThN7RYyRiLpwfC/QeZF/o0i1SyD
hpC+6+DEdTk2XuQo92LeCK6WPJ/EF/Tng4nJ0tM8ZCmGrV8xeU8sQt1ZeVVMr+L3ph1QXbE95Grg
xvLBIWHEcjKQ+HVZaw+c+HD4+pE6mawu001BitO7IOzF1v7DdvFLanl1fYyIWMbzUIUxIG4/rbqK
EhP3nzl94xhFOKrwS/WSRQIa85qUjBgrSuoRN6nbPd6lh96lTlJGZ5yu/KQNAFYnW+7Yze7bjUFP
MuwJpWcmJortu5J3t+hhmmntsjstNwyKOWYxOwMybssma3dviQ6OzmWiFBWvS4iWCLaj8T3gEDXy
QtDMCOapXfw/KuDyU8nuWN9e/HkhecAD7g2TsXM47O8VjGC3rCrA15ZSWxfjtYqG4uqRSd2oJYkz
Xs4e77Dieln28fgDdpyqZ0/ahYShzPcT3T3sg0tqm35xoLKxhUoAePw1+tRWzLwIfLBj2e+v1xVL
foQoutxbCHN4WRrwnLlNadls3SAh3nzE284dRJ6Ak6g1HaH0rOMBXOoOVheLBCIrofsT0SQqKlqW
Gr/UIfX4KyfbXyf3xdoeZItBcPuNn/5Y3yOq6ooiCofgaqAo1IH6azmFIsWc6YFWcNRwU2mj4+Of
Ic/YbYwN39pc3CP1F67QJk3QJFU8Tove+80SYDnSiFbo7/itT6p68u5sZmeD+My4gWhu2j1LujQr
qTYn1SE9NIWB5VnZ7wwG4MPbP5n+iwF+x3yguhJsGXOXaWWc+iJYniS7xZf0uV3qGadIi+++LttR
E+TFYB2xkjK3UdnGyWXnNcJK69yrRuBe3PZvKHsr471Qgil3ubxhwCpw7ZRZqvnj/3IN8xBAGFSM
oxFBvhRpZWRlIYuq2PfPIGvGYZxPrdXLgDHpvdcovZnunIVEqH3rEk/DBccX1rb5vGBmnwW3onZ2
6vJW4Lto5o7QQNlhe8pfDW1/Eo3tjOi+LNlj5GttAp802pqlbeA64o7S22RZ/ivqzTNU16yb/Dq0
sRAnvvM9EtYeo+o/2PgXPYUSXa+1RdmAEqF+1xSO4Xa6Bpjaidwq5hRqOLZLey6zM2Te5FqC+c+n
yxF5xyTbzCMjtXpix3E0y9+loxroVMYM30wuv3DCgSF+I9kV5XnvqCCErqJ5jyo+IGRYBhHtMNgg
aAyooFN+W3R+HhTWsKaeSoaHreXILVMJhoSRBHjSAX5J+emxAqCdyauKY9HF/eZuwCAddG00cEf7
Yo6isIH8MWm2IWj7SwGeV8f/7P7S05DAfFNGd8TSxtr03/i27w+EY5rxH0VmGIBb3iuk4b9g4EIJ
zbfjc0d+nnkNqPmtw/uaMLjTBFi2XhtPn0rxlIrDZX9n3xYSm3VP5PyGMFeU5yoXCZKZYPdIgSL2
SCM93NnD/GLEYHSAecdYRPwmN2m2gaP0ii56fQggdBxuvD7dxJ6T0v4iL2nXnq1e3Fz6+jxb5+ZS
nNULvinYAnEjauA02GDMYy8WZGYpazKGXSPWL0COse0HNcysrQwjUtX8IFS3E6H8hh3C5rk9YJsd
dg2GqhROq/AHhaRV5bbgBm1aXa8iG3RD0YXhOQZuGhFH8W6Bdftt2pnsZUAf0Hh0R9BJ3B0cUXap
8jDnrNHlsmsE6CgOJ/w7E42J5VN6Ztuw2UuKLl9zZrvUyVjTonjkulAG6AuuU0UaofW/X281dE69
C+/fDRlDhohBXt32YPdsj/pVG8uLOtkMMSF2OuGFrXcShUDfBWXBFwiAYi8CRKi+zfyXJmdQec8J
9Q8GUgWjtOHvVYhBx4Wb/VCR//KmhbtblAKb3lWBqf/5ePFGu5FFKyeTx5TILw+usiXsKeoAAnis
gV5g5fq1JPmYYSux40LLRrsyWQEkwYn9oaVeEAskg7jNaCdihP2T1HkULIhoVs7heugNga55ZPJ7
9K0FOx8g3L9HdiAXkgk59NYbHgjPmGtm0LSlttN66BvBby/nMgaFGjBG1LS6XC2KaJohFEnPOnAU
2R2z9pA2yX0WiOGGlqVf2LcUuZUe3qfXcWpYBP8NCwt5eRDxJdrtkZoWR7R4VgvPCGqtfaWCTnV6
uTgdtG+lorc6XOBoUnn9uXVbkin5p8GA1dHRhkcUGYPqLr6l4PIKG+ybbzsZYAU1OIzVTueOLkft
cEkw7N32SeDeMJYMBsJPpqSKoNBduaxSiPozZn85ubD5TQbU6HbuU0BzhljYb5Shsmno9FjClj8N
os/BpugcnuG1Q1cVZlNiQbvJbkvbNoMY5/X+Mo9/kPKRjmFJHwbNPuWfm4PY+NNNCgBJqSfP6OvT
9gTsgoo5nZDkvh2piAKN6s28WzfgZlJfTVwSSLuL4jUqG0eTgPBa5uBU0KC9FhhDhtpJa9Z8BvmW
nEBw8O6Jeio4o3npOPOiTTaD5Tc4ygqyYQL4bQsUcZ5GblkXqbOZcCCQrjkGS7P87PvK44SDC3Cy
PpBnCKLr2vpXRslTBWiDtKb22bMhSo/WKj+Rwp7PUz7puDqQLyH+Bu60BKsx7pLB3W1f3chBJzbi
/k9i0on+wYNL1Yzb8UugP53y9y6mvU7g+1V6tO4ARWsYtiSO3xeyHTSwH2D1u0xG0tvSqOCqlx2m
GkzTZ0XGboavZII63A3/lDxZv6N6RqTbs3qhhyTwXYBaLKB1kfTuTVLTQL4K2BcpR8u+D6iUMCAz
hnwBPvqIG/kXiCTSFZY+NjP1WSCiMuUG1THElXP5QnMHMTPg1ZEFR1/DuV2YQUif4YwBxdiCgq5s
KejZGe//zYIgJtUT45CpGUICkzxTRvxYyN1geXoVtwYL90p6r451XxR6Tm9/EIzJM/VgNoI2TbO0
71udLJ1rr6PyEF3f8IihNKngjMUx8jno3tzW0p4kd9Wak5JQ3snk79p5r1gxT99EtJrnjowTAvvq
Rs9nDdLoiwWWZ7Fn3VcGTedrw0YaJ2Yg9vuM9cD/ln1K0cAPJlI9Aq4Cw19CEseual5/uMiK6jAA
nijm8Cu5gU4gnY2rTTxO8M2Chz3zWFLNCuw8RVgwV3utmRo8rRVXZpw0GlMWw3pFgfdNpuW8wab3
yWYcx/mXkOo7lGJnWzTt+IUWYWKFYXQkXPwJYfnMZheAqfOcK9ZCCcj0/3uGPmV2krh0IuHskVw5
4DiGWhr/hHcaniRff0YEz9QsqVmxRuzdntSCIpkBQbQX3NF2CQt+woNnyVSXNMKiIzbq/E5RHFfK
90YR3PdXHfrQQFuBCyq5lNdpCEoEiC2WhbZpQTPUG5w74CMqMa3tOHBBnvht7J4YWyxO9tGPkXj3
tw3Q51R3Eaf39KYrtleXrOBdigBMMXLYmUQGOxZbMJdnabzePRTlr8nBkUkc3r7teekydJegAqOx
XMh3FcXPl4Z/WIBf7+ah3E/HR2YH47jkr2lyVGKBQEPAWEsgPetIOellLlGL/IrGszL4xh9PchkZ
GdSRHJNNi2747zdobZh8WbcehB3R1JfPipBUEjg4mRB76wOdDPdSop3W5OD/XAyCu6eRA9S8GDve
xClnmtQ3k1CTsIvU8/+i3D93va6sbbmoVkSyr+ep4WDW0S6YH1EX05ngbKZ54nHwPcjCUsxEjAxi
5vB6KVLAzcOIpgAk0Nuy2n6b/27CQDZHmL74kO+g0oD8ULFZCejJOfiLAE+dW7RQfyh7ZmLoYyJA
0H5cpbMViWe5EPxqThaaFN+kXwLodhJgXrxl7dtj8dqhYhqLvwhBoC/fZPgE1nvZNN5crQOL2ExO
58KUI/XwMpktmgttTzBjFhx/Begi3waw1yFBLCeNf7FHUcQgb/QttIrFnFBApoldkRELWSq2+wAC
Nvsic390kDHIIQ59Ud82fOC0hTSEpGMcjI76oB4eyRKrKCfgl0Knrt39vVSK6DNuTJb/cyMTaMZa
SX7zVkgvaiKW6aMmH4s7vjq8n5hHmAYaqGZ/yLU5gmOtTK/rBNHiAjcYuujbXrGFwWYL5dg6EAsR
rDdAKR58E9gMZX98L51jGI+JqTv/Fjkq6FnzFSluW4aKTPlii5ShLJh/Rp3BQIHIf9pce9zuvi6L
uDlxM1I6QE1ilCLJ55ydDvs74NkX/Yu4UJsHPIaljHwh5XUw8JYzgkhJJM3xj3eV5nhXDEmTiXJH
U2jruu7iJiJB9dN/UlLLRvDK2FR3Xn0TJaxw8teZ6ULANBaiOy1pPyhUXgYEHuZL8O4J9qdFZMG2
06Cft2zu0LfX825Wp0hP2J0vCRaieRVJhywr0qO+UFfDfjfaOKO0LcPeWSKSj9q4/DcBGNKvpD/V
x+gyymL4Zl8zWl0UXvpehY6BT3b6G7pSba0CMQ99hKrEswLepbk4SAsCp/uZLkhfN1BE4GpBNBIh
j10k5qAjdwyO+TMthQDvZRDao7QSJ+GeHI/4ISZvzYoCF286L8R5qJ++37t1WJs1qrk/S1dpOlaw
hEgy0y2vQTg0fDDz+VK22e23HADmFArKbScsw+GJZRF6Rj+AqEO5yiELEtpPUt9wh9HKNWvYQTcu
c76glgfnFPrmKpOWtySYlgy66x490/2LE48BSkJKavncTYxP64LjhTXazqBiwttg1OIR6devsPrk
uPCWjHe5eFMpMJG4gO+VWCV1c417G7Q1/R7PMNzB6ktQzKsLB27Hw1BpJ4hmq/tLRpXc364gO4+q
5iAyFwxYQbeNqVFLyWu3BcJXG/k/UolgnM7y0HW/GWok1ijNv2XIe5mjpmVnowQs0r8R69TLw7VQ
uwWciL1TZ3rr/4LKHNZbXnIvarNDvuEcQkNR80S7pzJSkVSvs9UuvoG4CwdfdVH/xYE966aYcOKQ
EdGxS4BowEMRhXLw+h2Sjv0AjVPLcf0x4sb2UxIyK40lxhMM0XZ3HXWZtNUWNpFdP7fcBmg8ePyi
tMiqROhPSUKsQzw/GknZxO7zN76qufkrUitY2fMrZO9oF1S8ebhudt+cnoux+GhA+tdCZuq7gWfE
ak60KzgIviTo3Pi3Cv6cnhK/9ZHCzyB2ibmUzDyNafj/oiz3oL5Ol5PeJhPwkJ5H3iBz/6zG7Ig8
Z4EU/6a6bihPVXbIvpKAZ3hiQRqv6rHjScZ3pBQboJfUdb6WynLs+IzQz+VNkv3j17XSc7UZ0L3Y
mKrXMF6qYP0Mmq8dvrNIYakOzfPSbOgcTAgbseiN6DNHUS+vsUT35RjIYnwkhqDeuae0Sbrm+IIh
kIDXiXMmyeFvhlzuPreiBvbLAXR7LHKF3dpFWQCCCenZqJeLTR/onFTJuWmmmYMX+kmeqjdIQ4B+
tY2A1+UHSRbu/5tnHJIurNDI5G10iyJAZysPo9xZxiJ4G/4PtHc3EmH4I1PU0SJfk8aJXcb7+Vv1
G5OpugktMBmzgHzsw4xJGx7HzD3B/PccCJxpaQ5PBr9rHgdpYZVU+FbQAFVCFX6RZ0q0FpfXaRdv
pfpa9n1IBMMdCFRRmt91nzxpR8XCmF8nu3ctwfIbdEhyrkvbsAO/g7B3CSSKkacEabSS536vAn4c
97Y5MDmRHIyXUSU9bk++8oAsgmYXlu0DkTZmZ5ldK5xuRO4wNHBhRsutGZmIVKBftN4gOFjbfdZq
NulMtKTa1gn5wnAMNHEh5/ckeFWVO9/sUAVBPBTOgRGO7x29kCjr6J3aydo8P4dxAkm/4RysSn7v
/xLcH8joLh3UbreCXVV+qwBMYQtEABtrEGkcTd5xLxq4S1t4JLPvvDr09jr5njt+uRNN4FFSwV9g
noc/Y8/bjXpgyHxsUd7BVyk1Z3RjOk0LwSPQ77NbEwqkWC93TRvdGrSKF7X+UdwC8eyx5h0gbDdW
ZzoEl2FyDQCiurizqqcnDmr7DTGhFMS5FVB6DNdVwAKlT3svU0GnqqDP51ga8thlhKdVwlXgExKm
kPqjiywyHbH3nYlySOCIknmpsmF+4WT/zC0cwJFfBxqbKTyWY5fdO+S3XW/mYg9MlkFZ7OBOajv6
c12/xLFg07/1LJ1lqsTlCnfg4xsCWIqodBKZpfB84c9qmtReHO+WAFzqjzMzohY+eboAlteYY9O+
c8xNPlKAsOCmQmZHn1d0B+ka0ryXVL/9+HTqe3umY8u+NBVImbf+Cg3NkBfhsuJAFaFVP83wa2FR
DJQ7U2V3gRatfOOrIzD723sGinZ4s7+x4hWjxfZlgIO0w1ZKpxfW6Ct9RqTtJ0NNhKdDFwr3Nj5W
Ollz0pCPU0A+mqA9XKgwvmkclDaLO/VjtEblsqWCdalDSiFj36VkNMZZL/Q/csvzN9GGxTgrAi2s
9D5wcEmWV1OwmBjAwI90HA9z2tM47cBgjsZt6BJiAP7ghhWRIAO4YcEs8hNSG4cC06irc1B6F8hM
NpxmTfaxcaMRH1IoqXXyS75fVaWfPUmXa0XsmibSuxXIa4fqU+SuS9WYaUng0oCMKgvgQFN8peu/
lwTTJ1kCAlIHswVZ5SA9/3rrZjt/AJBkKS/tiowLKlx9O6Tc0ih8hvcOzx659T72VCJEku5nFPt5
QePGAqD4pe6OkWPKTkmjcn0IUqBaUFv/hGqCbINry3ywQ2i0a+ZcNdDbbQW6lJnw3opm00PH4NYX
a8XD1x3Zd00DgQmV7hfdz6oR1u0eEtxU4toquEk6CRGSCJkoPZKx2QMMLlwLzejyEyI4kM0W6DCq
I9W3NkxrQdDBjQA8rN+L7+r6CdLO42/Y7+yV9JUQvO3tKTr7zT54sH31LOMSBQFkMMuH58KsUfW9
Ma66+6Um4x95E90gKNJJg9MF4CWyOyaIfA6bVz7v2DxOubU2jkXIfd2Ttd8HUday82KpsGx+qLYL
vN2qKjDEPNMfQ7osHGvx8I+OrlNU26TWwiy2viBbhHiEduUNH6Seoii24dab6HZHDTWGVlyqqX0Q
D9NwbwO89MMluQ123YshGOVHsCfGNujoBRssqa5dA+6CndNv++y4WZsxHql3Tz/VMKun93W0ZXlx
yZ1CHhm6+FpjimOsKS92bJn4sBpxmApNevMZI33/mmdlF3OBrkDbN8qh22rQvTSCgF01qbWozn71
sqLWilnh4M7fY/cWI2T0yoxhPs3Mv8y1zyc0wG9IEDi1FFc/3DFiZ1zuwgQNqhQwxvzF4JfT8P9A
WADOoTKTYTClzVN6ENxARL0ayUs2QXU8DM/zBeF7P8PJIxPt20HTJhA9mu0NSGy6TyakPZUvD11t
MVTFUPaAcBlbuA3ZLjMcRXK6uMNccjNLNGlJ72dZrMkKUyZX43dFxQ9SEILz/7ufwbkbgXcPlFCm
GFis0euJIwHiJSXBe42wJGkiwoPOzoKYZJcOL59i/lwTkkO+CtuF5GCqO0xrrWnumplbH8BxXAeO
Qak+AOS/njyq8OEreEQ6M909dS3RZYDUBSlga6eFa2qYuFSIMihXcjTAexDbgtFhaZ0df2xvalQB
5gECJCFwd5pDf8eezSQGP1JNqo2ZUe1wAVpflwoPbOrOidCbKWLn2O99icyZdBT9V6Rn/59cllrR
Q5gHiBBDk0CXy/fxIbeHkn3bi8c25OIlVFAWWKsnHttBnAgmZbbVxIwNRg1lAU0en9LLoWCOGfZi
9U3tq2vDTfwM/wLAf0EOPFQ6U1wVysvoaMMFqnJtYP/YF0714Thfeq+RhLLbtM7NxMLGhmCTQ7xC
ZM3FHd9dKViwhdQnVk9BfSBbb17VzDKqg3Z2tkuUZghwrU7s5yEQEHFUOrCuTj1ImuqjWVsVuVLU
X3dAQBQjW0kBc5uFE0CQ5JfsFavEyUITVM78xedX48MUGRetWe2Qvmah28DI5ONfWx0fm6EczBZd
O1Gw/wo/8k26F44Wz8Wk42ANPzxU0f+KwZzwCwMm0ctRBtVFPk8wcX3e1HgsnKn5mcTryDXCBHZk
CdITLvQ6FrzwxTc0aCixRHgs7oiEUxmsrPMq1eju+gaGDvEJUXE6zI/1V99HXlQBmj1CMk2+71wr
1NWqaHh4v+XBm4j6FHjLaPVJ/hjcZGLaVyZ0LdiFU1dbyPH7P7UKiaDm0i9UvNCpKwOcysU/H520
6JRp2v0MAdancXqDnEp/fX7cwonmm/7sfNoiUhvLneZAu7nCwPHJsaf8tt/II4sIv39RiYSfkrt9
eIxUH1CmQUuxJUEPZz2sWRmW3xBrsYemb6NzjpHmk6WZpRlu2qo6lbOjGW0oTa7VhQC2RpQy8NGv
yfCqMGvs4gcCaemkgLj1nFYSvLnwznKTEpS+DSMCnkVfkYBbcMBrsrHeLnGkwYUPc8xNTy9b4RYi
FOXAb97+y9UJVL/P2sI4SQgRmJ4Lls/4cpL3k2Dh8OObR6XTygE2LV7GurdrcyATsx7KzElsaaAF
Hg/dhxk7ZJnGtrX5JsYyK0iB0AMxt12TJZWX7VFKLG9ARt4gaj35fiOJS/o62ochyLfOfgKS5Bdf
Y+ahWDUMLg4J949BxlsbcErMv0MWhUvwqkzMJ84YuVm9Bn0WRruLfoU4Ou5wYnQ5tKQzjhaXLkI4
2SMufTbbZ793rHCvn7RJCrSpMgXjKC8MKF7GgsSFFbVL/sfpNR7llACAu4SKH6XfTpyOxArVngcv
r8BHCCY2TzyvcEJwaKEKCtvHCvVWNKZZgOykwtTubJGzqSmwcAZN+T4wm9CHS8cPRi5KU99LBtm5
alFPM6OuIOzrOyCwK9lkj3MMjAwol25yCZucIgjCrdy9MoFFolEOOrhrbDEi0Iu9BmXviwELCAyl
vZeP63kL1AhIUmdjAi6TsCShvsQFcltN98DrpFCHQdkGYGYeLbVMIYUyHhKz3QPsumcLk/cu3GMK
wd9rQ1MO8my8LJpJa15EtvXZLcb4WF2llWejgniZ8km4RiWj9YGZIigRz0tAqp6FZOounz3lEXmw
iqdkpmpjrCbcxYQZjH6TnYJKi0OM/eHVF5fkqOO6TLsTfQGNzA8XjypGq/x4bcK8lbma4nJ8hIuW
eNXFY7ZDsRhsEsk8+EpaNXN3KjdDUh7/8JRQcSb0Dunj62h6wsUm8RrHHrL9Y8QILYPyeZTAvDCi
ce9dWwcyD11PWyZpugiAhh+G6RwujzQ+HJck1SNMB+usseCxMrvp5SRy0scfXmSVg8ToOMPZFD0H
VgM+8PxVC5kJKVCf+ix9sfFHHX4ercQMPuB9W/Zcr+acIkkurmwso20wDLgMKElrur3QgL6Kxyhs
oqZDxcdbyPgsJB4EOtKlp6GGbkNuINOG1t7n13sVt6JFnwqI+Xl6Fcv2g0/MwGcA4d1GY8UnhfLp
zfK7tdr95cVN9irFqXVfWeuKlYGWvQ/s7CniTlTP6JxCgkFYd1U2aGLyIrCglImJ1HHz0gDaOL+g
8zmpqUKZcC9n8PKECA00oCn2+oazERrUorrRdCESxuM4xrPHc+WLSWxNBRKtd8CTu0UEzwhUD0Cp
DJQfk3ZgJdUJX1dB5lFTPVvZuWuJPkOw4h8wiCkxsy1ZWUoYmWqyk5AvV2KRnviQpdug81H0Pojh
sK4JTKC+eWfGtaTSiQpPDgKB02+7qeK6t2b31LzLt1WdqEmOdahO++ljUv0P00rhj1YYqX/Htoz1
U3AQHdjxfmGPEB9LD5cSX/v+p4oqQNXB8UwPglfvmXyac/SeFqpeQJCgH+kSj3oKZnM2XmlzefdM
d+Vyp0NZdgo4XbmD+cnC6j9bZspbUoat3N4actC/+X4y4iD8ncEKIVTZgrLCjHmna6+JjJqmvoTo
NgXQ7hyWA9CmNunK5ZDbb9Kq70ycZfVgtay0MwC2NiadBVdh4JKwVmkZ7VLjvUDx5GEhVeLgxNAJ
zGcwmQwjs17/P6SlTmh8RScZAPth0678N0d5Q9kxBPWjWMvAj7v7Q22XlYTLS8VOO561hQ5uK7/j
7QOn5t4+x+jAVnLbqDDfWsA0VdA5OWbA/iyv9ZQ9uANs8kctw2w4KfovsgN+h1CQ8wSjyFdqso5R
AnOFvRpvdBoT1G12HEz/+w8a36PiVFSRGCQS9y4Ft1DiQpGFk2+PNJzKCgnsJvNQGUQC8Pg+jFWZ
PMl55EZf3skxapAb0f0g4ZrCbuA5NouTq7W2PB1P0D4qUvMWZUZbiv2N8osGZjMiNFnCPl6qc6tl
LSOgqYDFERqj2QNoCvwbign7PHeBbgMLRK1gLPB+VZv8s1ZSrfi5HVbnJHuXiMkWzg/GX0kIfVZT
C/7QQLrRfuGpOv4iWDTi75jTw8ldlzFF6Y1zDsDi1hfpJDo4d7uBiZ9FVKp7YTdOppMo9xqER53g
w/JCNOpLbFvzSb1mmwRQZPGXT9U08+orT/fkwWGdWJKCz3Lz853qTUFKYXHu8Wg5nhVFAMrtnhkE
3sHyz+rpaVVJLjSAEg4CkkxIMfq/Mhpse9xKzDBajo88TfjI4PYUEUIEAL4MlUR4yY/lvoyexXnU
YEsoCVmpvL9ft/MckEt1e17WLJUXx0byuCI3fD0GC3XTRe+5Rk3rsXiD7JhY+4pKGO5Ht/wGu6Ng
rYsZdtQ25/YnKHmiWUhZtpoK22LQkhJx1NFrSkwRhGGPWsT65K1egpKCxEJQKzi/3XISftEQAjop
2bUcZVQ/6UEl4mA0teeuP0Nx/MrhmPVd/70pKmJvNA+hgXyMfogJqtqPctBA3zVeD8vbPEIMkc2z
cdl3qoGBUp11UaJlqOM/by2XGx49sCOu0RqvJtGqhaaXJnodo7zL3Kcr9xlqocqmGAMw3Xu+gjGS
EMTPI0djz5HXf+xIqPniLugEDFpdbOgIqlv5xxynjceQXKwOGhmImb6toQsY0SEJpF/eZecEGPlp
Rc7ikyt3IaNdgwWXtt4FMqu/PkYRZY3yuJmPuSsETBLIvmHYzUJuuYXuCCFHG3de4bXRs3feZUq/
MoNa7y7Z7w7D/J3Kv7r7IX3hGVupQ5wba+lLstXPl5U642HfY/p8rMDtvvQO4rEZJRskR8DaZls8
bPuQfyiO16OQYjgCP+VGcdDTaLaTjwwP2OVni0KZ5aaulQ7ehEYfS+MLT29XzlviWXfEO98cpHQQ
QjMuvDhWV+ZUvW5W/kMdN7dD23J0mV9sxyXnzcuBHUTDemar1lTYDi8QrmcygrBTxYZEKTF9AMLh
SZY1Kikenru8fVfmnLWTIchpTMgQv1DsM3BkSrcmO6qP5JvTEuCp/cF+Oqcvbu3ijsHW8Kgdbg/j
pvG+VdyVIqlrCEKXLdUVGtCEUyiZJKg2wqlcYEjkaAKgxE+Bnbo5cOjg7qPDNvLzUzoinDfjFFgx
vshlfwWzhJSyQT44NC7d6lFbejA7Bg+sySkdiz49HrYmY/yrOr+MxqYMeGi8NkGh6DFzYbxTEaE6
iRYVnoSCnci02bpoUGeYU/M0oADCRmZ/fApR+tAwm5qmaUrD6c6xU4B0rWSoLWuTooIgSPjTqrDj
/edcT/cEnP6ZOXVHBNzdt0ksfH6nLWXRbqz6L+K7FvTnMy5gaYfiUUjvlhLv/2lvHgrORHMN/juS
wAXJq94EVBEdZhW2FcUiKOQeTn5T3vcAXUglB+JIGugW1uLYxeOCaCS0UwiFCrduzfLYQqDHuAOQ
xEcS5iEedsZ/ef23FYbs811Jn0JM217b/xBKnb/o9q81iOS/IVFGHe9eoSw8oNU7G/FKgx4QvFxZ
huGLUjKr+H+aFuHSpVnxv058MbbxlfjbVaFR1QzmHmw0ZKWE2I6H2lmaaiFiF/GDQ1SsWX+yysOf
Fgm4/lRUul+7/vaLLnYYA7IJd25QgBjN8wIvME/LkBmrWGXGWJRjf2PJt3UAaMgnpUImnRIUA9Nw
W+K4fqIjJlFDTP5ucBsy+IQUaVW3hkn8zc4M18eqh3q6SXorMqL6FOj61SYU89mNEwuNvg8B7Th4
an8fIEr0qGU2fBYFzpWxaFVTLmbOUIV1iW2/0mrbLv4bCDCLCelXTECze3b7NVzSzzrlJ3Yx7YqK
NmJTH8CYT46zGb7FknZaxSVT/KDbV2j1w2YYIFAm+o4p389VQJ85+KcgjfxsT+OE7B7ecVoTB0dz
LtYyhQua2NDBWVdwljQkv4I/3F2WKW4gScvpqW8iY4Sw7RF+8ZhIYsCou0EyFroITvbDfeo8dCaf
UkT8onMT7+YzUtYO1AdS5G9SP5srS3Lgyzt21t8rV1XjEO4ysfblcF3W7a36ZVC0ewmzc9dFUqMr
GEErm6a0BtRkj4z8ZYOgpFzQ4LSq55vJA6VKfvCQQ1+jrKqZjNc2ktcT7FI/c2a5pQUe77AK/2qF
lhtqrb1MkohguvjgYyrKeKMTFnQR0F1tdwk3J2d1POWGv99GW5qZ/fHA7z85htwG8IkTrB1Nf/9t
6cDOemKjEvnAwpVhL7izEM5NQhQ8BAbRNZnlrweNAAtBXJ53kdNx8nh+nUvFK8XH9D0AvEih0Xq0
XYOjx0aHGjyUSXKBkd/MqSpMlHt2cJKvSYE8qsABdlFhGs6OVaJcaAkZbRELCeUtBkWoe2Y5NGpw
Ly+iJFzychFHMctKk8r8L++Va41v+t7BrqAY19N0aojadhM1hblZmBhgc7ru/H6VvJ/iNUCEGh+/
U/3c0Px6z1BpsG+/0Bh13lV85N3DM1OAvCNjYxPPKO5ZEC6d7Mvpa9ju8CBzv6sMmC625oy8jsZ3
O83aBR7eo88uoWzJfUL52B10neqAyoHBnzL1JdJLnjbjSqt3HtGA+Ko2iaR1GSLe/m+pnEjHYc7S
opE8BQWb+XzX9fj3LMM+LqLqfxCTLZsnaGtv406WEGtFt7ham8xAQI6k8aLpleoM0n5wAn0yjN3D
mJjGpuIDGHcGec7sZ4lQA61Ov8Ss9IBv5rTmNXIWh72dF98Lj8Ikipuq4Jr2CAFh7Bt/tg7/Eth2
Vgo75TP64neHZp/xuTNZSpFcBgutccWmDZj0RU1kPRdcLzS496um1eLyD0wbqAbtUYVyvrRjM0t5
DZ8T8AXLHIWXgShdmPijCxiSGmNMPN0Knuh08SfcvUwKTv7qmB8DfWdkmsZhrKSUaAzGCnOEKLh1
FVxmjTBJ9RwtdFNpyBN/tcPLt1W0mlgTETN5hvzdBsNqJmol2BEo7ekl7kAlYhMiKRiEaPg6yS6J
5DnJb4a5oKyQE90s88Y5QT+desTIn449s1m7YCtXJ0Zy17Bip78raMbAMUJP+Nzf2BsYeH/w3KT2
nXDnLoyYtQikZ/GXH/ltEE+YsLczEXiBDtp1FGT8eEsIwVZGKFjpgNtKHOTAny4xC3gS9EY8Ly1p
SA7Ajtqneeis03z8c9EGHcOCPtDkkrbIcB8l7f5oXgcjjHiDnKOr6nFhmmLz2mUhQymQxyEaXDt3
6WTFlFuihyAnN+6UIWHT/v8k79Y+H7C6cUPVk2ITaDHe16mTA+sHc1vDnqf7Q9BoJW0zgLJAQpRl
uBBnZTwdLdpkvCJB7GSIQUXCkkHkHuMDKImSWnsQjqvP2sxVKFt0hEgQHD3oIEgIzt7Lyu5byGlP
5IRLOzQWit7fz9KMIAzkKEBGLYe+G2Wdkxzptj3GQpxOQKFlHDvf9pFggTJlPX2hAfjVhbG9mMgj
dgS4qGPEPCSmI8u+mHPKF3Umihhxku3qpGdWEl9O8Exw3flGMUzGmc5PU5v6I3kgaW6knirPHU1Z
cJiBI4X/QNXkBzAfqBFwCekVp6s9C/Ib+iXGE/J1rXXCivSyijM3VrMWWrMmP50CMKDFSD5ThBvq
AEuv8oWvnfvsRwmZYwilPEOJ3i7QoM7VoFfA/ZiIbKFtoYscLPjqQimLZn2YrI8Byem1EhvgVzwg
NRKgFBHJI0em05JavAhrBcOk2sI+GRJUC72XhuFCX2Xd0Ws0P97ISNZeOZBIpFlzo+khM5Wj/Do2
v/zhPSE1oezHZAWGXgnlZfjnqRtu+TSdOdNNqabN7u0JN43qk/35ieRp1Yr7dQARtB/CwqILDVzr
bwxhuvo78xZOyZ+yMsDRS1tSPPdFiQBPr19TgDeDpcxFTtRREBCa8+QqYM6q8jTJFxJ7cQzG3k2x
QRF5kDPAATqDwvA6DBZdfNrdFqBWZnpGYBl29qIIC7ZyB7cCVlsloonxSObFWM1vaXDSwrwt2Se+
LysXW+HrOGJ40lKPCeY1NqyiUwb2MZ1CnPkBqBi/hGvjauroLzEgdMr1KYE5Bebw7iB46hhN+RT1
3a+KpoL0VYenMh+PGu/xbrDBabFKqXYcGdyXthpgAjovRcP6SYGArxCdgqHKPv81lqMWKAy4Ud7e
NmUYsHoM41VsmWbIWtoJhalWDLSgRxw2y3gc1ECZZZznoaIhTJzpkLpZbYj4mVuF0O9OGZy0qH3K
joS0FdzVqjNTFwQMhJe3KxlbAfpRBDmqVU43MLpYRXnCSyEZc5fgPKZOeqrvMmeQnCrDGZcNo5rj
jsy55kIsXX6ChGvoHRc47XhoQ31S0YBe7zcppa0kDr6JoSBYKpYlCq3AlxkMIRn3yaxpAeMcGAi1
8CIw5LhBt+Rl3jldOoCM1LwEh0tYDkDlvDy15tZdVKKOhiwW0DApPq3p1wCssZU+zJ+aMhJdKkIR
S7mI5eKYUV48OkJRjletZUGD/BQ0qSwZ2pE/qY5e9LlFyA010XaNbpYwwRREAeW+KalWkZ1J2GGu
oBhiXBtAI3I9929ZDzeC4tZzrpRIALEOOSGuTMFC8pdIrmOy+1Z41kjQgXJsOBD5gON7VFnRLT9h
5UJncZRcJnuYNoQ/gvBRFOKfSErgoXylW32QmqED6yIPRntH9Fcowu334AmpJV/qz53cUPELpwlH
a5dqghybo4IbVgKdFO1L/g8jjY7C1eaLGqwygzhQ3JKJOvzg8oN4Ej0oBWpjeDezo62EmAvgijLJ
Z7JlhtBX4FZt8uhqoNK1AVwZwwct2Qj1F+YeZUOfQOK7gHnAxAHBNHn7xQzKpIv7aZLZgp2d9jPf
OJX1nkqc7AYSGsCrulKzEHloHKcx0plPzIof/9EJH3KSRKvTz/8YNNQu2Zmfrx6jtLqOoBidxGQH
AwyB5h36OZx8bCFdeQxL7BbY4LOCUWhMjcgtdKF3s19MVsV+UPgU9t4E1R1yxekk55/aix5IuY5E
64NUXifygs8RZuYmGhLSnZftYxS51pMraTsMs+w/ZyCRdKc+ZFWerDUu22jZ/xLOuyTna2WcXFrF
tuBdZ2a/GfyjIsdBUNQ3Q9slxwdDEdJObpPsrlATfvCvGQTmCGWvNFSlxL0LinCiPpXpv3O5w/GZ
H0PjS3Z0UCmEGvX7bPh9V7zGqP/BjAki6dksSq0Om6NrwGZ3jmHhvJWlMzTeEWuJ6k8pHu20++MX
+N0bHhI23TbxU9KQiPCUgeoaoJ2bF8A0Qsm+E3wXcAGyeBkoLL9OisHlvHiKSEHdZSV7w4DiOO+N
YukLFxL8cBUHphBkAK0d1LXtSepHUQwy4DxeKSpmJfhM4iBdH1wyCBTELjyk9XcauyHVw5auCWMj
f6EbZMU9CzsiKSCYHPRszbJIl/Ii0mrfeScl+Cos0+Yg+wbjZbtFqKX4AccjGjlXV4NYUNqibZrq
sbYfpyMcEUMrx1tVyeXHoRpdBEnWTNlogZieZb4NKCnTJARA+uz3xDmdj065chQOs7zFnh+X7iaq
kfdr4A1lGynsbnp5Z2XanMLoKntU1/lDlf5m5dA/6kYZScp5GYO9wPBts7K0ScnHShiw2qPah/IF
r/ylAmxg+wYyl5Mx6F92wKgwTNZcI9mgwi3gqqMvm6c6ogoAazYG0L8bdBKkIE2RkbUJSS8iof+k
ceoiBpuTHFJfECjSV5Sz3uc1VlxLBBXp8LSQ2EK/A5Z/5R4s7LTSxmTE4zqou1CiaN9VmCpG8jLE
xdlBKatbU1FwbApqGQc+7Q4wS7rVIEXOU/AX5gjXXraizi5dYtZJHXFkpuAAJw1Be945EbcQwv4A
NyGcpUwSaWvlMLwbmJkPUZ+S1M8hcMF/IpaCUkAjlD3/cIWyQlBRV0/zeW/eZO1frsB38NiAEOp/
4Ajut3yxXPN1qnK69mSGtUghFDSH78YfbsYNDqhzwbO6x/SXhRfm4upeIQcZxTbT81ue3LWCuZUE
aQ89Tv8tbt+z2iVVKJOOMgyLLqKKFLfE4QlEUGv9jkr8zfiaXDGYsDxdwG57xCLRULh3ChzA3MRI
9Q3daCYxDf74gtRX51oYqwtYyY13rmuxux69QowBoKmzJ9PD9aC7Ol9fIqrrhehvJvonE19aX4H+
luKcuEox6emGQHgYJwykzAsyizO/8Sv17Ja11sNWhEf5dIEEdh187I7fCiYdmVn1KJqGnrusqdyu
OSrOJNKay2xpn71C2XasG8UfFxg7lUf7Gz6HLadDuMXo8WfS6MHjz1XF9SWUQcjARRvzKYEnuz1+
bdTO2t9KPClEeJhB/YKwPQmyj38BzpcExD3Z8GpNk75kPITXT2yppXZrL5MsP0J3YEkMmiMl4dka
o7EsKfaGl9mN9MtHrKfAvTzGk186tR3l+Yp7SHasl9xj92i9lUlSDoZ7iR6wADV9ueI1b/pyalOZ
N8KuIVZuQLlShn5DYpzw0OuTyI7TE4kkF03tu8B+05lVvYdWVjt3mUQhUSstDojhSYsAKNc1Y7sm
YAHLjnfSTsN3jhp4IbhVrTIOwuZss/5DnmdRvyKinn/vu4tHG6QB1iRqMCFabKDyJOqwxEuPxJS0
156uaKFapnMjrmL+AbSzaV8YY1Y5JCg84UdfYZUaotCej16zO51J+gkgcWV5GlIxlDXaXR4F916H
o4nO9gol0ubUq5Y0Q2XOCEXXvy4kpWQMy2qsnsBbP4Bs++oFW2jRac5zU3W5rIfmXISteR6zPmF6
37/tyGdNMHhCPLstRxi+CXL/CRofFaOVXAEHkjLd9guh+pRnWQByqa6aqayT//aTDAGvB5XQat4v
bRV3dtkkem5oGPSaWrrCtWmXKQHC/C/sbVj7pv5DUL1Kf7GAaq3K1kWiketkJM6wWthGFBqqOrCs
Yiu4xGn9nnc8kLrrRZRB4j/R6M0nDXU3z8ZDlast8oGmPcAKoKmJBheOrhgZND71NpeXBmcm69d8
TdqYB8bRk+rAgKDa9idSbxblPpW8Vfq7xR/gkgm/foW0MVD2k5VVAQJepo6fTmB+POdsvA0Kqhg/
KjMfM11fhX9bJAODQoyOFJSyQdwcvQ3U/LBrkDnqo1/1UKBYoVuvv/TsjSWokgjnQh+0tppN8Tf1
TvZhjkY6q48f1PJbEx9G71OhLtsr5zsV42H5ZClDIZBlhF9HV0wuEJdqLM7SFo0Xi66YaItpLzwl
bnCc+0tWJZoWvLhkl4mcXkKIIeHAYzO/aMu3GKKAU353uIjWznZOI+ogQetseW2ITSiqVRrVSDRh
GI6/tjw8IZ32wUWONka09wya1kjec9qqTybkHDXIVkj3uBYUVINjC7bVTMkAcLGn9s4BVRlqQZgO
jHQNDMkbZAEdzAMrg7rpvpQ0GIv7pDgZFPX7zpm8fXvo6jydpgP5I2AnrUSih7iEqA2Afrcn+Xv5
EI4lPNRvLPoCCQmg6GH/afL705H0zUCoUZvdeQxdwhv8x6zMdg3of/oGj8q5107iqhjK1Ezme2lF
Mf5PCumHRVhoZAnQbk1K431rHIwVfSGdvI5ntz5y3KiVAwNTmf+FacOrdM/ZkvAUxImrBdBh62sD
JxUl7wH2IWSyd4Ak7ILarIHesiTdKizZo9bDdW4IBXYI3jfVjpkiI2gUF3mBvTXEqErLy+4SY4ut
H+vrbhmC0/O7fVyfEJz1Z2WsVF0aeYsr1j63Fcc+sdzuBmm/iXWT0N/StGOyLjnZd3BsmF82RhQn
yXagBres7PjWTNDyleO1F1e3sqGmKXdyEfz9NHNkXUXBP5S6ex2+ggZi/rFl/Sq3u85ktiFOm0Gm
J1er2arEQuDSsW6O1jHGc75JvkDyhyi71Oc9QZI7Jf7rjwvT78rrJ0HLzIArBP05bX2To0wWGfch
b4U1SBugjsi3d++uSdhvAUQTAJZ8T+pOgSXo7tF/zaPKHPdMiw2uPv05x+wkF8GWtMyv5ZeVlrk/
KQwwVb8vCtArJ9qmREQY58XZbQGzqLOwjlg5Qxn4hYcIUH0RjKHqCE9KE79IDBr3zMiuSjsE5lO+
N3U0yxHBp42okooPNilauNs30f3Im+Hc8+H+Ql0zI+Rq3xHmxxncZT2eqIaC1LPL/y93YARuEMyY
BzPydJgWxfU1mKk972a5pOjPZ0c+1DCDRD3ewBKm4mflAmSarP6h43gJdfUtW48ag1z5DYr1x1EJ
axJdObCRi8A+6shvb7i/ytzAvdjK3M1G4CMTUj1cWBx/LkYJXnEBlIWfL86SKElxdxwNZRsPEHW9
wsqYf44F2XmatMBYQtIbQNzQdNRglKHWSPGrUKmhj7QlVCe3IMFNcnPabhs2x/sf7PiX7FLnqEag
hNZMmc+3nDl2QbMupVFlJoG+9V8qd4hh1SaRqsr1ahF4VZSQHxauCUHV8IkPwnBOsLAlJPwXOJaI
VJFm5L7QIkXS+IntOVacpNh890HMrRfo7Ycr8gCfm7oA+kQqw8KbySq6Y9mW1FUX+fwsUaZ950P1
JvadRyd3EPLbYO3S3UCwFqzvJIiQBMlDZWyTd3qHyIIe90vKS2Oe4BelRvuL4PEoNL+tsX63RJ/i
1hFNXjDK1xh+zoZj5OwNIfvv3yVWyMXqnhigAoxx0m1a0M+jYnUNgfTncX+6E10KKkD9UYaA+B8J
FX0Mc08pT9U4Sz48nhcOxpsfMfaAiyDK16sApwjFKRIgOaHqntzvog06jWoC/KDQX0/UzS2ywZNR
kx5YxVcg/NwLkYxosDCjHprEQcQKS/BoUJW1JF813Wn3AqAwjI9+7tnzJkQ3GZk/uTG2YbKqW9TX
voiRfKNWQ5okwfZRW7FbcAmrEB0PMja1A6spfc7TdAPKIf8kWeDt/qVf4G7pjLe6Kqa8Hh5HUF0V
E7GjY2tLM+ptYqtAPnM4/aySB4N6oj/o5NPQDySTY1pN6YJ03NBfwut3SCdtSpx5xSZU1rRrOEjp
zvi1IotBxNjx40Sn2AxQ6Bwwz/q+j5IXWvusoDqJ8L8ubriWt3juNistQjupwQIDv+sTYJ9BP3EM
u1AAaw9i657grlU6NuMOWDBJe02sVONYV24Aj0o4GRaOguG3lDXjQd+5/BKJSf5DJhE7hJSxBqtm
90VpEc1Oivho50V5N7xakLmUk+V5u0mx3tK19aORa/j+ocn87hbw57xy/6pCGSoBszUtXFiBM+PH
Q58+SI2pjWyx3CR2pbKqzjE50dxXtyFiVkunAfK5sBsIuPB7K9Awo8f/95B515Ta/JRhYP7Uf9Qz
yTXFKc+++icOs/w/VUUYKCSGCarFA3YmVhTfpdOBW4/PCP3aegrl2GWgUGRvbd4YS5ZNSoiPBIvU
g//51H4FUv8HvladjLkSlglieHNQjcke4jCTCTmIB0pReNFkt4A+3cLLLrHKHwVblSeABiuhXMsa
XWUEJlVQnFY9YbSHBJIaGJB7MvYgszXZTOlVTveHkHrwJzqrPf4Qo5mEEZU+QhSSUngANNeIykPg
2wkpqEaXVy05QIb2bQM2RGbXcGcm6ZNq/uxkp37St2H/ohZH07kNZVMMb0BP1EWDGsvxS0RvaZ/c
v+2fIHQKD/zonUKzlK9UPkmeXa4j5rg5avscO3Qx4UAlDBEM59NBFWju/P+P2kzBybIHHY+UquB7
/lmto7JUZjj6a+8mlNmyqpvtNPeKyXC/8pYTOU0k5CtWC3W5Lv7NoGPUyEv8woIlfNfqkLcAmKtf
hAo8dAK8QseSNzHDhtYQVnnniDWrk9lv36ar3gtlzf1zVFxdo948Tm3vsasmh5BA6nDRVqd9gi/l
z/NQNVdZrTrq4vB3/mcUNmyQYQfXPXeR1aBhB1w3MbKR6gvXlGnelxRoDnzh3WkD+xP1XU8dN1MH
EqSM52qD2/j9wIiy1hy/Weh5pAGafsyVg0RzDWSBHILy3H9hVp2gB+HG8Gxm0uui2thE3Q3jGo7U
Zx1OL6wZmyak6VjM7zrnmDHUyoFKSHEDuOLR5wqE7Oure8u0CW0hHeUKKGdotvTEUzYMS6qjStkd
vp+7CCFQeAm/BXyVKzxaAxceMdpbSfK0npMxpZ8tgSExE+RQL0DNG305GLK2Q+5x0bv0yJZnd9Gh
GFokWjCz5+0MPH6MnudDdwX+rG46w5gCDZu11voL6KpQ184HzPSRMSevTShc+OPNjbDWTtgXP0qa
bpRJnmLHHTcEG2vh3jNt3FfKAkBK+jmJt6N2LvoPRuAiLbuoAv6+ELTcb9SFkLF4IPesyJzD7jL+
85RSLkamg69Lt5g4Qf1DyQZI3YxeIV0X340Gwf1AkgMwRgCJO/cszdMsYgkHmNAAetky7dxkhOWO
zdJz6cDl0RJO6H8eo+fgrSoNI3dAdVTfXtZr5I1NV2s4sPPHj/3yzMUjfuGPDiWogQzcLpU1OaB9
XYsMZw7d6TQ3cXPggvOmjR1i7CVAgT2VtH3ossLEppMCh1rn2C+KVrkWUBrRUk74cpfD4MNN2eGF
Vkqee5t01xvr/gJXlBD/hSvKM4h74a/ZsCURPEj0W+yhrlwtkDg7oEoBC3qawDi4Ck1hd1p6UOao
5vft6cLyRUX2I1+usalylRZC5sJ+3fgBPVPAgDR6aZvfF4Zdr8sy9ZeGOAdGWpjXnLFOPpdwlFfT
63zo3CF6ITKiP5SVTpo9Mpd5Y7f6jOVvmYxUhEohChOr3+5WE4re1VFLOHwn7iJ2rD73VQdGit03
ug2XRVhRiQY53ct9ObvjmDj3ALcSgkqfMrY3oBjt6hfHzj/yjNZNsEktx3aaY5iS6+ENCyDCU1OM
UNXUyGC92mzT242gp0+vmRjK4NJ1WUf0/ikBJGXsizHb+856VgutRAgPtsen3Jq7BlzAEWEm4ueP
swdZ+53xooLopVBjm5a5OQyzLYTNlhDjAVV54ti3um6GvJftVFtpK16y1KZ9DBEJV63XMzOG00hp
DLco6z7ZiT3w1J/48LLnCuatfrgrgMfico5M/znSYIp1QynaKq90EYytMxsLFKHaralw0R5x9kgR
yvgLIDVQvKIMDE5w8d40nFfSDZU8gkL2sTXCRGnNvApZTzTrJqKj9yxJVPxDyZJvqFc9H0zpS8KI
HgjDOZCcMQqJCc1mxMQAkFm36+Z4M85lryXAZjqAWPuzjdCUGyCYGV1pSaHnWcd6U28HnHGCFy9p
jRtsQc8NAuCfaMHdahX7NxKGduRq15HASOezHLN2J46K5dM7p+20UvU0TcPBWb0zBXk3wjlU3zE1
Eegy7WjrCrGIfK+Min+JbjFkeE+cTBrOcCy0Xu/t3yaV0qYMEz2CJznf+GkHh1nbRkKuKZFwMMBf
YInKKcN8+fPRCrchB6O3jz+HOlauTKZrU1KutM0Bom6uTI1SHi85Vn5K7Ips6fgVCC2aVfb1uBEi
w18TP2oFfPyyky4foNVvRI5cRG35igm6keIZJFfcY4Z4XOIjd8DuhCy7KPBarVYME/5bg804UZiE
bBJ52nwsbffQLLf2ZkMYzUKsdSgzWkdTaiqb3weApHt5z76rfBViS7z7KRxJlX+wEhvKpDMc+j/q
aiUF/BQ9Vi1MzZ14A5TcQjuvuDcD0u0svU8Zfpc1BELT3x26TiQbwn1lVScWWzlMWr8vlFUA3l5k
Zw1Oru++hOOQQQvE0tFKkcmKNeBYFnSe3sPRS/UrxK6qXMp+XJ4tPX0lSb7KJbqGvmK98p+ci9Cu
q2k4BsVsXvUAAr7pVnJjY/gXhwpIYpoF/2+78JaKac+KGQxlF0jzHCUxgq9yVscmUmMnLi9V+iYd
WEZHyDO6zBjBT+le4p5DO+Xa2VMv3mjSWCD3fY4mJl8Qzj+uh5foJj3Gg1a8w+D0OCygG19R/RmD
LL3QtqbwsVLJrdheWlJ9WsTGaHjb3a3QVBFFdVyTdFN5/jaGnk8OTzT4N1BPCDp4KrqBCJSncBQQ
9ZXa62w1BHwd1ziLLHaDDRpz3nZmh7o2VBxIjQmQz+TWwyjjV9Sw8v8ms/elZA+EEJOjmH50Iebi
ASn+6RlrQDVbXHPcFSjYweHYL+9+ZJzWMbKEVhTQAjHjD4vJ0ZV9gpXcXHJPHm+QjWKeAbMPE+36
xlsyFDGWwVo0Kf+ZfYkxqU+rEjCM2TO0QWi65+iL4Ud6NQV7oAqWVytQCQ8lM+MQwM/eMtHA/d1F
od2vxMKXbtPxdD9NnbMR3fLDdoCu4O1qp8lVv6UnGbakqh5kOcGMAFxCLHaHBIlCNUiUqCS0+v/L
is12ebwPoCKBcB7+kAqKsbbZy+6XqGTYg+AagiCBZfmOUwFBUE8fBbB7O40U5fzE34SXseToWNEU
dBsx4m5eKP+zToIJJ5WhCoRHH0BAXXaVrW0yqb5uRkqpJZF+Py6m3mw9nLvzQlwHVE6G2+xV+HFk
GlsfWVkJnDcEN7iJe7QkPF86KEDaG5Ff/cJZ/T6CDCBbIIrpQ7FgvOBUcEU6HU2V21YvDjLzJTBR
tzNZBc0l4wHw0Z2kkmhLzloMT5jqdbfvFxD6uLMU9zmJ070REF7h3ihuJXNECUaLDzafBhacqhP6
wHy91/qzDry2QMq/kArjgt2uxyXX07Eb+sLtPe0fEJt2JdAOr/dh80YslsOhQa1ujB4A+YQeYSz/
3B5G6OOoM4H88Skd/0NTVKumApj1MgYtlxeWjPhlaA0ssH0zdXsbT2R6val9XAlChp7E3uorHJxo
XPQiDfJqbvUg9co1y+7Z17fUm2+jWCJL4chLX3DKlB/+Q+uSMLI7vqnhRXwaE1dxMi7z8K581ZvM
M6Tnlvc9qfH1KdWNAKWMSEoSwSXFF/8kYbA+cCbbFBZ9HxHiJR9vgnjRk1CidEgOe4GfqwhKxZCt
43yqYPklfjMaKptzO1GPiWox1Tzz1S8IvmhR5pJBxG6FKanqzvP70q1GHqjSavMDhi4Fn0tsRl56
+UbYtjbAafXmEK4BwN99ZknqneVfmq1KiEKbDLdLSIav94HPgjY5bvrNv0YrSvLfrzfFM5D2yJ0j
Q0h4zy/Xm/fH2qitItpdCAgHC7ICJ4l1XVDIo3kgo0BUdoZF3eT+LjjH9ffSgrjXXy9Dt7I23Jv4
d9U+AEq2K8KD9EhowuRfTnm3DM0vozaY/xFr5Ll7LBEooxzSkBWjn4oJAS0eTceXzUufBWRANTvh
LC2trnxIkQz9YMKDWcg+umIo6Xgbhj9w0s7h/KIlME904HRYCwYRsWGMaz/Dwj/flnEbXkJy4TEX
XWuXgv28ww1bvdYp0EZg0ASqnxsAchmobp0qGSYXbH26v0X2dHHZL0rYn7x8m7NqJGFE8tOtqlaN
AK55+UyM+DLtMYndLTWbYXPvbfuLGmpXNOnWNkoQWDO8Ke/Z5HStsJqb6Oe59+AZd29JVFbaX+Dm
ehic3uxnScs6uHxeC2Ci9ReuVl7/yqg4ToTsfLtQuhzy7bbgjqD5x97ePcoTzLPaez4adiU3Xwzz
RVqDK0SdpJ8229oRvQIEiqFTeNUKCzrFmEHQswjtS9jKO699ZKMcPZIEQwKHyb48D+w+Eag/pT+g
3dDu2fNzN8xru++kQzCYRjzFT8b5rvjhGpHT2xd9BZ7Net+kc5uotd2VJSvLVDUMPxhOpfpgHdtR
5XFBmvuFD9nErrXfMBnbQW6ECnaKeiYTkKzTVg3bVPlkSS4H5T/ieeOGXMEQ/1IM21H+WvuF+KdN
pIYGc5AbjO+jpegdUAMmuioHryOyqTFA6VIDVMTAFK/CKwGDlwEcNSou+PCF9Ffiid4+sYfd+cZi
EHa7b3J8RNAe4oE7JoHSHHV/+t/I4Fhfez6qavgwwMIrtu4YF5lfiWwOhqO+/DKB31LUfEwRePWU
OdDUC/FHybsKRGJ06AdB/xRobUfqrTGS669nIF7q+pnNYvl25aJ8fLsMkCVuIoOLeMfmMcbRKfzj
aO8Sx+KH0KOqvu38MhtocnZUUxZ72hxnYQLk1r1SfupdQNXTQzcxoTrDCciTTpwZHH2FcflMLAu/
J6iRT7TMOCpUExIK0S9sWTf+iDinVUm6N1DT9gn8yJCFo5e8ap0WUDYyWIvzTbATreABkQQnzXHs
oltUt/CvZCbELxxUJtDTLZMmXBRAEBBgCcBk/5oALFyJcMznpCGX/wgqbQO/VUEICjLuFTrNHEi6
rdDj/jBoYnlVaFEM4e5/l25g/1S4ntSSqjl6jcKxLEkVrogSMNRyYEhB2jXAVQZrfEtIBo1tfV6E
Ql6HMi8INyvsiD6IpTRJXtpJlIkoCr/b/LvdKFpCOyb8wt2n4JJbfqU9b7ZZ9Ha1CkiWgUGM/sds
rTF12qQ4+Hw3ghYT18gwdjEwnv1NOCXyU7jhUp/xTXzUfrKgzZmTYWA5YeUHjiomDtX1NmxCUs5x
aPKfF6vVx5wKyP0rZxX+kdt+ADxVbrAVpQERF/Uf95YXW736yf9NOy9VzMoIVPMGEd+R+VRYfOTA
JOXwHMSQL+ztJFJpkO3HQ6UQw74ubnOP1RQ49GexUjNvOQtsFmiBSTMFxRjxx2ntFxx3KEZ/r9o/
2zLYvGb6HvooKgNO2rMNfAw41FWvLghtNmagcr0J+G1favwRONdticNo/4TiOkCv0P1kfxatBfws
e4zRQq1ajBZHybiv7jLCXuGzGSabF5IOuScfHwr5w2IZKMNWdMY5/KwQHG04BGS+qQCn/UCeTAHO
mXH2qvTP+MJFtWD1mTt+M/otf98atPhnxgrlJ4d7Ee/7dDXLP7AKhdmB4BVqNaFeJ36umGsK4PaV
4jC5J6poWpVMb9/k4B1GTBo96yl+yF9f/1aBF2O+CqJVeDwtK/oq9XRGG9sHTwJgCFeK0amhA0rr
KKAYzSma2VpCZ7coF+QQASOv7lHtHaW9yDJTuv45lqbAa6/2qRz0q223KV5solHQivLE/Y6Glj/w
5D0xi1Zwxfs1KFOHZehjfl4/YB3Sma1gsY+Xtw2mqzLeckuw9hHpdGtt78YJVW6tptxVs1+vnjmP
gJ9FxZyuvvQLSWhe6p8FgMTnFRxigYJ9f7U/G/g+zPQTdpo+2F5vSiigH8oc0Nt1oyx34TFm6wm/
cQTcTt5bEjBsyIxvlgmx9fDp5fHQqvUtLz6HXczuMUwoENAYVEgsw8jpK2650A28Fr1nJSkthSJA
xYVar16riq3cEsngf1Xz2g7Ox1DBlXBbL1Exlnz0OG/zizGaMe8IGxQwHJWGYUoQ1jMQ601DYyZf
yVwPZYUpxCFVyvKYrirtXFLV5ICzNVxLdyTaoHujJ2Trb1UkzowxrZ5LlixPD0v+1XbCF3J8rp35
OXxlPDHdSnIlbt6Re3neTV6QvMXOt0ec3i5HQtUGXWPsobH+tI201CGOUYUIKpmcjzE+goFeveyN
21MT/WGd8clhkolMFjeVDJ2M092RdRb8tzh5qr7PF5DIKfr2WRa9RVLKOqEgl7OhZAHVYSC5r9Rv
n0kRaBvvHQ6yJeAAkN737rCqJ7dgM5OJPtJb5V0GoIZBq2oWYxBJu7RB6rch2No0LtVjlCXyQuYQ
6HX+0XpyeA06rbshiFvKgPqdTJWMbJM5J9XQbEBLsmDm2ap6+wu7dUq1Nd2GymDCwMdUQgWFT4AN
HaaIFm7yrjiun+udYRRZLkZLe6neE9dQwK9+n/eOAC55I/D6//s3XzRdILgF/kdl0vzUhJHUffNI
ESFPHGmpmmfIBZGex6m3Iv3MDul+OTPVa03MLlvVBQmks1Hh29GBcSNM6pA0/h8rrLUo47g75OYo
ltnBhiNi/dVZ8jBBczTaE/rSEh2atmRx/tVnYlBSrHYNwa1QfYxjJ6P2Tj35XGiYv/3yRcKsibRX
n8EnME1vom2GBvI5CpyHhCvgv9OMWlWAjbCy70LtNRD5PAHuT6Qzn73qr2a3ZkUIDJc/QfAS96J9
4IwqIGUPEQuz+oFi/a3ERokzbqANFOuXN/ipPZuvvtYewgc20s79zoFEd63qNWRuSU2GLpY7BSg9
uJjWxOSp5NZkz+RNX92rAqBk9udNtJfqzxROY7rI73w1D9tQZosMxOacpzJ9rHs+jFvQlHhbRJOq
UW0mAlgdoPYsqpzvc0BVIQ5QCwHOMuUThrMhzUze1HXSpx34on6HHKknTN7KXgADpvCDxWurAjj+
a1uGhXC4ckGczfJSIVd8n5FjOptz1Op2Z6uv+RtYe2wBgv7wSJwVFw5E3a7anPu/yuZTdjAGyslp
1nmb1EvEVguEkp4HO5dUzxK6PkLAh2pThLHUNvHURZNR/sYb0EDLqadLLnMwxh632xsBeyAfQxIx
O7eMHsMcLNT6Tif/VT8I5dWjIKObhUJ6ASwJJhpUeGQf88mtLxsAtXmJp4qiYvilQcLD07H3x+KS
e69/+cOwSR0v4rnOTf7UHwtu55JWBveM4WexsQA7TELxs0f3yUoM6VMEwjruRS77hh2PFcYrq+Uj
XZX5mSW1HqvZOY6Q+MR2X/fsl96nZy21Ougaaj4PB0zCbGn5tgTo4kK+KPMa4Kh1tREi6QvxfU2O
45jn5wN1Fbc+avXVF70hcv3IA+gqyyi7zx/srb9nWx5SI263Zh5laHA6UU+GifeTuS8t7yfySWZc
LIJGPuqc60jNwjJkxKC3UPw3Mg0+so6N63kcK2OLBdrGZ5fnrDmSzrFETuV/A6J4sCUYgoxYNfqq
T33hK/oQ6zns/c0zO7i8ABZ5E1YiiYMT9X7jW6rZDFIdqIU1EtqT7QnZRr3+E5asfGNTC21m1Gzm
pDyLqLqGHgfwm/oHsLU3xwhsx+9omd21yjVAtxpFjfU8uzkPgty7TipdqMnsHLZzVCm1obfzQazL
Efu0eoBVgQQCbWIX7vHbCREvXYDPn5Cpf0vC5PcJLwy0jonTfeXbBTEL61f6eel36dKImEiWP9sB
Utp+iJAmBvAgFTV7uYHIx6qNoiIpCFV3w/6trQkBiqoKuTlPL6RuYNot9yR37UCCua6OBTC4A8zR
qkZUe/ZarKm/tl23kWT7KG4gwUwzN3cn6OE4gvIAGGR5QNmh51//l8yLARqMVBfNSsUfSrIpcnOC
eiBmhldzeW+EykaDfDqJuqUB5+upgNgOMS5MwtkWbVav2lpU9dr48/1/DQTDIz+vuwaPmn5e3ihc
8KtnwtDoOKIOPG7zuMbnFNH2iw+HPwsXF46uBCNRR0/cjOWChbZ1BVzNtvu42N2HGZbEU9CF+mcT
dujyqXu1AjnsrqFf577cwN1U5fpGgWh8pajx87YbBOEGUYbzty43ztR1jbdee/vm8mtzu6PfPkae
gjCVF+Cxv5A7+4Ju+ll0ipxJ93HBlDPx8bGrtwSCwr0OGKg8flVjLAvH91dIjSEaO2Zx0V91lE7U
Lvxzr2Ad5mN1J11EgoDABDlHWOxFMNAu7tJnp2tCf+5vgSflIFKWzOel2GBypOL9o2BF7BFcVX4n
Lm9m0YyFMeAT9ujPPeq380K6qMspwpqUu9x7cWCBeYYt8GJkWkzFkbrRbCjEwQB1pYd8C4nrvi/a
wjXz1VUZKLFTjhOfJ6jG4bfVQqNq3TYDEWiqnt2xQlRXckK9J2F4/dxGh5CATKdEKWQIq7BMLdwW
e4n3AepWuYdHOgvmn22XnOCEk8uv5SN7bKGcZQuUYZ4u7AWdUsbVjCs+YYrBJK3cVaIj7JYfFJZ5
PE4B3otWLVaG9U1jycFrq2ktb4poJh6VjWEasv3vYic1mDyk/IZoPYHHDN2F3K9IgcVT9aEvi89l
oLS6yyoyYACXpFNIyGR9hjiPF69DMOnrdAXdXRfaBO+XqOCOnsCyOFtwQIqnCUai23ozA29Aknum
3O1nkQmG6sBEGUCpLgV/CJ0d+ihzrJVWt+Qw/TOdIDbcZIq3KSTsd4ZneRTMaiZm08HTYBvjMU9p
paeWjUxwN2eAtX9Srkm30Go2b5BHoWAZ5UXoPr1Es+VL/x0AcnfnafHZtLUkGfhb6t7n2YLcCs9V
a93klR244uds7cZp8/VAbcF1WZiLsNvVVdvElk4KjCEwGLQrAPEQU227JD6MokCVAJIFn6voZ+lV
nZrxQONMhCaBmvK0lkKHBOYODczNDcg4QZolIYx1NkDfxu+SmkMON/8acvgELDx/NwbOf7QMAmKC
ogTNVxfvb7Df9tulVYofN5+0OUyTmawuBSu9Lypz/DWHkivEGPeV/aumKwhvlb8AoY5Q6KgdYctc
LnhdH5+AR7zyTXH6gC+JieKmf8g6fnuIsU69jt2czZawp+lrsduSOE/3Ovncdw2MAuThWnVM1s5g
xOroGyo7CQ2bbZZQiy6A5LRytuBmbnQ3FDoCj/MhNHi3qoKDvG6F4GQo3+XwD9v0pgPY39B3QWMz
rWSwfooT2uXH2ab5TEqju9c7dTYS76FJVm+RLeJcr3DT2rb9K6CzTveiFPxftmfAwHV/UdL4cYIN
AGzhDgpcpcsiAs0KDDRndMovP0KGkBKucGHqGlm9MJSvrpj4ukT9+P543p+ysguG1C2rjgnXVseB
bBCiR0DYzLBxJNbo1ECvBr3u1PCSxQvcyDajol1zFNpl8v/+dsR7TedZO6LwX50Eu9LvcGalU9Zu
Ay0oIamkKgjPeQcFsSYibFnPMpb9Z0Lxu/gVlNyS5AEMttt4R8X4v0V8LBsBgjV3Na8Yov0tYrUT
Y0veLMYDH7qMu5KAAPF86Rc1guXZiDDE82MEJsRr35RZ4nqsMuGbSduXA1W8A1gEUST7keUZn5Gs
EEL4l1cPsXy/SmC18LlmYjjfUmCmCCNf42/7FUu8OBFGP8ZhSP8gykGC+xaG4dqWpJXC+OCxG9Rn
qv0TfIvHg/tKEVLVW9nnJ/GAccuBlrO2+2Vtw34iVgYtFm7WYFBJqDf7G2RwGsXp7NLQCOWkV9RC
uowV0utULI/HLwNtvqBbfWSwc+PoZ+qFZ0C5DDFQXq7+mw/rGCP+t7SF9vnG4zVYlX/H9GBRHqBE
B1Az+rCoR7WMpNJvZnK4/6v/SzsEtkPx7+HQjM9eLJsyFD9ZGuSK4wFVTLvT8fbW7ggadEvUfC1L
9SFWcnXuhqLEALVN6i5crfyQTTQrIihMGempvpKv9KZGKKKsppMvV1gGHR7+B4S0Pe2aKaENWlCY
LBiGbkNdiQEAembACl/B9UlB15LGpmVtBE4VJYXoZmrTSrrduiFunPVME8WbYKSmuAN6YJnBOi3F
dSg3dDHPf3yFFxUHd+FBa6IKZf3KkFqWVmJyMHdyUnn2x9XOPpMYHzjLJJXCOuvM74pfwOWibhhM
rYu2ORn9t4xTbVZv2WNMprhZpuwnTxshHd1ZNXS8LGQHrDwEibHM+bGK1WwnmqAsTLMayfngDbNX
+/KsVoDRi6Y3EajHQ+SUPKKPAtFLciutD2pPovkNg2tNtHcgnLt8rMZ6jEZcGBr6MCkDXN6gXDF3
yZeUYmIRepL0zZoV7ccb3ecL+TpaT13FgWlBd5LD2SMamcsWIrJ4IojdaC1/GF9l3k20CxNmJoEU
d0Ofgxpo00WrtugJIrg/QDqqejnr3qbvRe4/mSsbZChfGW1MaewDvaNdakBrFqzY8jJUSVWq4arh
AeRqZs9MqrWGyxDBnnJ6v58V2/jmILrxl4jrQCryGUItNtLnexgGZt6tx8ABIeme3+wXyGe3+hg+
6nllR2i6iurQB8UgMtpM4ujNr3EVYUmoyX4QVbU7eMtD74OuBsQ1Y+N+oIqiQODIENCsJYY5a58q
ZM4QKzHNsUFjwyVrKt3cE1gNbyrtlFN7/3v68qlWoGZOIqkRLnq3hIquCTQ36yDiU2TTa/O9LBdw
hjouUgOEHoo9qlStoI340CHtMRsscdb1KJocV+GZSDhBrBtfgsu0RsqWTegtj1ZnMafyOJwo6P9e
df5InPGYofvSDnTIoHw+p3Y6lWiTlpM0XHCaH2TgbWtrYcunrEj2bBITHnbtsUHyV3MXqsHhBdhP
6m60NfmMaRd8tm2fymM72/zjO2rGrY0VlTqp4Dw46psIiluD8iRDMoCNWCfmKO9NlrPQRa6FuTzl
qlCMsw7rplxBjd9nEiL3G4iuYSnKyMvPw0qsW7cvpVF05vlE0v0IUZyoe2v1uoZKIPV/e66YyxsM
CWMDE7kQCPZSX0Yzc5FHLBh65EQRSMvgQc2N8+4B4xTk5TlOrEZj818hz6liGqkg9ys/g+PFIn18
CjLliFnTz+OOlEkGd/xQA72PWzpupdIgcbn0mH0OBu0TNhosl0K1dUOYjYunAzi8g9+H1aNwUSnQ
bxepWJZRdQRuE95x0/OKq1Inq35HvsLqZx83Qb0/8vxL87NR3RmaNjCc0BLLBvhZ/mIUgq3GchDM
L4kj62ij7zTpsL0DdujEY3QW1Gt55TPoqKIDaUfFxysY4Iy5MafStVcJ/jO4qlvPIZliz0k+LNiD
StKhUddF0VtyC84K1hprVd9ARUja48Ct+Z3DW86/MCh4awTbh1AMIdr1NHRtOgDlUGFa+mWhy6Xz
MyJesn1j1Hdeujq3h9p0p1RVFUHX2bibaFIbVM1UHkqOGL+NbF/EhWEVf7jQf8gz4Dmroa2Mil+1
OYpS/xpqIFN3ykbJTep0v5cCpNPQaWkWBUfhcwCDg6cC8fPHrblK141vGfScOfH9XVNccw59Ggxd
8naq16inshYNs/+vgwJGh41Pz5eQqqxoVNMZegjflsS4mHFJ0Ibg5wT4aAE6DHC2Z9g1US1BCEva
wQBfGGv2tEtz1xjzf1z0pusR+tZmCiBoXbf1dEfCOWedEKmvoEDO3GbtAwM2r6te+g7ReBaII828
W1fj8d92tR1WFiDtwrRsDaN9cpl0tbNBJBA0b7KYc/HCzCuzmLyugmQ+nHZWKV2smSQcJanjjACr
dj64OnV37Okb1fzvgsTaliolaiaLS0Xg9tnWS6Q3+4i+vwhJ3eB9CXTXdCwipZw9ntzeN0vvCa5Y
LfQVdGylj7qMx3Me/l7UkzuAaJ4gJa7tfd0lVxBTW/4bvqiVdhG8+MEmKM7ewkTekgybH5pkZuEw
RQa6cpqB+Qwc33tsK63dPC9V6sCoTgOv0lMKddGVKWmjhQM3k18mN1uPuIx/oJCaY2X9UdC14bRK
e82UKGgAkvhVb9B4L8xkfqiKvUupqeTsWBHiISNv3BgwySwkHfDO9mRyB/wrOIbPSd4ZSrupZvNd
5vd1AyDP/fjplB83lyRAgZICAQsYu21alXCC/ri2n+FKUjlD8Eb3QluoXgUjIPt0qYVlwLa25y1+
dgSxf5+MC6END3wFmAshDkWC94qJbLABQ9V6UDAXl/t/x5aMXo0vNy1qsYTxFSChgG3sweGiYjy5
dY5gpmeNgU7LEKJdiF3gP3k5h6Kivh2ZpDw6hAKd62CfDzVzEmuzzVBAlL+ToDERiZKLRJys5y1p
WO0XjTRDRy58bcYqngDwy2yQPJqF/9ImYV48M3K+4LvabmfcoWMnsB6ysZCzh8udNujMNUJzbcdW
9WF+18K+wZN00SkdRLhkHZSyXSGiM5o6xsuiEhD4wzUuD5pzDQ+nJAK5eKPZ556falrKNggQGKi4
u0NNv7p5gwpbMjdDuQRAa2CIbdXK8F6tkkbOAZMcQRCfAdG8eKsxOs1BfydAftuflEVEJqczmHnK
izE1L5JHNXA3fh86LKDfrwFjp14/MVPM69cBaDZDK8QyqQ2fOSolaREZ4OHLjII0FzgYzQgfqTyg
BT9OailTOJq6meKGEmtvDnXfZrrIQtnCwNGZAQijK3J89GAe5j7eGPhe29SbtaNq/U46Asy5yvSe
90SAf0fbMpfP472++/duGZjLmBp20ZxPdhk6RbSsIZw0kpfQISol5ay0NaPP4J9gmHAQ/p7cZE1S
iksf+WMK+5/elVRNWuSOs/xbnlnc5dfCtLxGmxB0ZbLt/KOxiads3XBfz/Tv7qmZTtBue4bVdnie
dnEgBfF2i6GQagB30dvfrfoHpYUKXuHyzzu3O9ucdVrh2HQx/906FPFlrwmHRnnf3c7JczPsf9SO
S+qroausJHXbexmTezbz4TTj4d9pIrs09FbvLt2lDS9H9PDxnUERM78+EeqjABE/x70nJaDTbBt+
lQfyiE6SYrZocfQe7VMnbthTYseiYtBQ2U63iKDvvUXklbjE8l3s3pIMTUrN2LE9AldeB0VXNdY7
c9E6y63q/azf3dtl1KXE31jsxlpfvJsYFklroJ+zDt14yio2jLraTHMAlCpVBditBPqlbvO2CM2s
8qm9/ZhdXzDHM25tZ+I9q7FVsdcMAnTYy9yzuz4nSxMGjr/37lG8OET3M+O8uhST668VOOGSYvgs
DWx7Nd8DSIbftaFHvnN0kS/evvsAzMP7bwo3/k3vCUDk7m/i//ygexWBv8uZAt2LqZLRW2JtA+Zi
1LQH+24z28TGQpewxGahMbqIoiwx2leXrC8XED0Nh8ft1EpWEk0eNwE0XMOo+z+hdprZDqFXMw67
8Zg3CelPWeQmXsR+fk0oi7oJy6H9ERdpONi+LgYYDa8P9jRzbWNntLh5YB4wZ758QeZ/MtM2cV5v
qf+X1ewpMDlSEDvbhI/SDolPFfBY4Z1s9UDv2DFMl1oSgM9KpzTE57KgDjlgsn01NKXokM87zmOD
SOmn4+NXNCrz/PVVg3DOZrdjc6cfC1d3tfiljjTHbg2f7V9KlxxV3ejkXot2QDsaNsLcyR9l9xmr
TwJHrXUKMOPxAzGwEvT6Ho3a49qJyRQBwmNbSsfm5JFUu8HvsWdqgQR6NoCTQBOXBRbKV+5wlFoq
QrRKbL1YsBAOO1d9Jyf9497gfTHLEHG8/L5xYqascovuCikc+qSw6riiQ6GsBSD3A7sdwL+RJ1cV
Mlsr7lCFFgo3rYMfcfLrfV5PA5X+RD4Z4Gew623ENHvJ/9nR1BLK3k106PFMHHj0bBhp2UEap0dl
MrjuamdzW7aQpBY+EZb/ZMgCuyjN1VjKjy7BKIFvi8xbsYuscrkLPkpHo8ECCBVTzVaS+O9BtKZQ
4Kp2AeyR7lX3qZrDJr/8Ec9GGf4n/xcIU+zy2LC02V3OTV5NTJKw/4lseqSGAYcouPjnw6B/Gjq6
ieKY5pgv+5zBGbDETzqYor21DODcGeqGl2CAJ4D7I72IimXFILe3qR2J9DTOi8ffE9No1kdFSmch
SP3Mq+fkSlmn+tL2DKKYevLoaGbxEfQeMs2LPNmVdVYRgcN9nkxPI7f+3twdmGyVA/8jkfAhiPS/
X1vQHTXeASTo/QI1i2UAE79Tt6ik63fadoDmtVU5Zml4CzLbc9rB9SlYDuZcP9fYkz2kOPauqfM2
H78LJ5LqFweHARKEefDBg4FlAI3TepAHZdnrgNkLMgfMS1uSXb5O0TIRNnIAPkRu3NM9nxjMrLdb
hGXowNXcEGzY49h11ReMC8UYPFjuqZOYnJu6O2yOtvC1mewqjAiCpZJHxh8JGHuuU6Tj+e4OQKYn
3xhFJY2Z3SO6wXOcSnrkr1pJ/0CVWQFsfl99Bp022rETFgJd0w235l0WOvk/5Be04lA6K4YA6/2t
vQkhdT4XqMY0vne75x3Xt5Ut4sIuW0y9oe1511lHmjhBE8lE8tcGAsrNcizxHX01wSnBbNT033Tt
HEO7Lf5qSg84Dac3gVM0fOx6Ut1pPy8OKKxWkAJCjJ+txPEKAWfGyIP9KAvFt5lCjuYxR9OSPeZc
+OzqoKqYzcGZ0U3kE6655w08LXlj1GFxxER1C4X/lXZ60kmtN75aE9vbG+HecuYRgh2k/sdgktoK
tmr3XuCPMCJqFtKqO8Do1zXHCSxFWp8p0r4FNxSSQtoix9WiMf8a77Q6hjTDA4AdA+dZhkius2n4
0rGo4E0bLJWEl2xHtFUhKq/X9hqP9H7xU1TzpMCLepb55xUlsFv1C34yvg7rAYYCbHD2xa7skImJ
Xhe5MPUR7ml0VTOhZ0YUoJ7si8IHmbymLQGZAzn8KuAB36TqIpU7J0jB6JEop7OxF2nu/HYGP40p
Co13T1xubtG1povgxpVdx9ZXk2AQetHRNtJwRrfcTTbotWPPIer8O6GGmT3XNA1tiMXi5JzN7Dw0
P+pIYO7Pdil3Vex0OE5vMtI6UNI+AmiFBs/7Mnmr5FBAf6SCVpVTw1px4N8Pfgd6WjDp4UsQGvp/
p75Gd/2CKfkI9tUNPP+UtoPaY+8cYIiuPG8OXhSkKUy92/a23Ts3975neMmnIW1l8eWpn2EklnWZ
GllilvIt2DOa/7ssDvPUznm+z/idB023nu6GYHSSgO9C2T3HA6e2a8gkb73T8Zk2KAsDAJRWZGpf
tE3I5qKHuL6+bsCyB9IeVi/zZ+TbYUzC9TpuPBeJXybadYkVEv9/DID9J50s1kO1LCJb0+5YqbOH
19FD+NPN8q2HgyGhD2s6S3UdtmxODJNvsDPRLsGfI6gRGU7Em4/IamuY0+KJzHVfk0BShS6/9oWW
eyE+eIBm0aNEoozwPi9tVmB1Mo22FAZ6lTNL6CIzl/LshniGU0MFyKkzmV7fLW+dfnOKOCMN4vFk
ISjo9gatEO+Hy/t1IQlbpQ49IncVaO5HE0H8v9y68/PU4bXjJaMZnj/JnQqd+be8fih/itFAHWuG
VKgEGG13Y802JzhGEqNYdNvAeRaRw7YeQWNrCfmrFEYIScCcpVxiINJ4kCJ2Hk+ins26I6Usr+E/
hWZw2oIX9LimOZw2tLeV5IAxb2IBp6nXT1tHAikCAvX6k79XJp/tnw6h8vkluTeOqs+c4d8OaOyU
pBytTQAyBRs7ivUnpqBQwy3XRZlfeFz7TIDFIwVixZZfDD0yFILdne/BQTGdIVeHO0vELYX5tf1R
KBxlzSeBCQKh5li7OkW58FAsABc8roDhzqXjyAN+5eUQJCCvHhZp7tTFITxsgCVcCYU/JZZgL9/y
qXJRAQUrM8A9TaO37Zh6YloqOQxRW5+t8JWTRDuDSvEgIkMRPwTDS4vHv6/20x9Kjhw2x9gNcHDB
AQJp4/rRwF/Epy2/0W9cheQUzjWncl3zrykNVS6kFjb0MkChNjapVrz+++aKEyr8peKHKnsd7xT4
MDxj/JxOfw3qso5kZbZjdM0t9f1sivfAsoKzTp8ztwxmpelPffycw81aP+2QO/6Y1TgtqmBXso62
JgpkipDMTRAKzYMcpXEmRNMMJLT3V8CZ1vSCZCz/sLRTj+xxHs/cBixvV5yunDHMCnZ9sWg7puE4
b3XZoKnIacYGCk05aFBeyIixLr6JZLm924nP4gS1MpvBEn/6yuO+cgts8+TLwLSpGO9qIOottcG6
bcOzA4nub4khRGPKVqNOpyZAxog1YCTLKl4dMPS5LN0Lp+hedjkJi1EacqX4Us9qWZnsCdheKYtH
yaNiO4VsWG9rq8j9uK1HiszjE5NGenhDZRrh6m7A+SC+pAZoN2qdcCgAi+mIILMWw06rc0npo1bu
E55etivdVXJZyMuZVFPiJMQLDFnyUtrFNYx2KoI8Qgm+wDipoa12vOVZz0QE44g4Nw+lb5j9Me2E
cJlfqaCp4kVe5C5f2oo2ZeeN2yezD6xap+4Ysq1OojeeowMT9YFZKZDbsmyqWrX2IirElCQlpNet
j5xtIKh8B+6aWlpQBh3b3rC/7i9bikoA9w4AvjinphhVKwdJ+dYWJ1nEv4zhk5G4xVRXfl2tWW+B
v8x7dmIfUcciCC+YEwd1qUmfPcFcf/izpuKHKvccNLhm6R1r98/XJmkSCo9SHXZaR/SixsBX+hVF
hFAnKaaot0oOtHBhgJ1ZlR6nS+ZIyQHZs05+MnGaSaS078K3ClcD6R9O6yglLUuLQCgMTcst5Ug5
EATcgFc1U35ZTEiQblCERcbdXQ4dhYW7KVXI2RrBBlEcHUXW/5Kz8k57c2ciq1fNEdKi3JvI+KTh
90eSmpiMT232fVLTGqVQ9DCMQHdaVMbr7kC5KWvHwoE/pgiXu0wetUBMqZFYIAYF3YLBV4t7p0C+
KOfh4ttvKqtqa+A50VBNABhxLaSC4QVfWTf5fxt0PfGU2xc6iOrBkfJNxxpI5GYlrkSIHPGA4BTD
uecWjG5ZQzHRhJkRDc9wrQjJhITa7cs06qWh7ef9SxdlCwPU74fJc7mKnl0uUo+MnIv2dItwlG9k
Az0AiTD9PsuzywPrvcP6RnVmt6u+pJBdXpo8tK3oLsegfeXaozDIwCCybnrO7ukPDuEVAJxlx8xQ
u/GG7+T6pFxAfEXy3vtbNL7cueZ38HD7rVGYBxm7GUKHwxKSv6aITYxl6R5lDwHeSEqmWpC185PR
sxlz5Q24SCfdtOEY0AY8n9QhOAmsVTCODZbb+tWL5VpUMyPflfNVHxd8EHNUoUhBqO6o3RDh/DnJ
JtrojXP5hUzO0jKyBwTbWiCiapEJrEoXfVc149lWquJojsoTbIS73UEg5YC+hf+ftUXFo9/u7aXX
THLDHXLWp40KS2z/l9M/gfUaTo0LZZTgiVwZnusVno4fkgHFLFuZHKtEC3Yf/ga0W8xMpwD19lNr
4nIOOSCjeyWl8n2uZ2yhIXuCywN7pTk6LBoeVgM4Cm+fC3nORtAAN+NaUQTAb3nV5cCXr0pOqMbd
WywHqlG1V+Pk++o+jb4rO43lGhTUm/byf+YYh3eO0cxa/IGC4Wpsdui6gp/03qbuNy+Px4+6GzxF
lo0sqdQbuCFDTsVkNcCeOt8xz9FQdYM8V7okBEkrha9gnKzK3rU0NMiW2gK9/udOV7/M/dL5lY5H
nW2xHAiSk4dcPSqRrz5hYB486ijM97BwtAgaiWPHwdX3DLTqGtna8iCYemVHjVeHPVuYjbvh3jWR
Al8qNWzMGG+OW4Yg704vFrh4KeALbjMWkMm3nEbJZakZ4PyQPRZhWDVvtyGz9XmJTCKro/OupJn6
jj/yK+/seKqUnnjhJbqdL/gc8ke9MitOX8bjPKWvu/1w/dVpgdMJpGzQFRbqAQQzA8uZE/K/P+rj
JFPToUX53jYod+i/SPhgXc6LhtX/zeSu9jsTYd4/hsmpJas5HMkbwmu1Beq+SYCJXbX29S6v3nQI
pPXQr1NAeJgRbS87PqPWXsB7TepoHrG8AvfijxPmkbEusRfLEOGpkQb8jEVvjlCaA+tO9a3cz5f3
os0l9obkKoibXvv/JzmgJtrcaiQT/rVkUoyVWSpAUjL+Hj8RIPP1FSrqJceN+nFaJhfUQfNs7kZ6
YtYAHw1GJ6Jf/OdMWZ4LxgIz37i9tGw5JJGBJo292us2qC8x/W6BxVGW5u2yRVfyZ9xBezzd6Czl
4RdQb5KFqhXd6OQtTFeAp0cxreDRZGunK6Mbnu5BRQPGI4P0Z66yBWVj0CgSorjeDVtz3AR6NUAa
dD6X94rzZPkwO4rGNisGYypsHlmmctqKsbPVXTAnP8KPT5EjduXMrDJz220aTvK1pBv8kK8ruOTx
b/rwJzpn+X5LR6BQ+UNh3SNKeQBdH5t1kRTJ+pfV4FzkhFxz7kOysNnF1JJb0VO7pvKwZbPMAAOM
2GbKXlR6HXAWJsUHIWF0cyoay0NIXrwfTUAS1TKeLU+/T6nQTLmaw8Li4V4suQ0HEjIptc1/MryG
7ATZ5f2adYUzzUu+cejNpWyEQ4BvfNi2NNqw7B3IAZkmkej/6Y6qLxhSKVCOPuDNKogGSZt+hCCS
z4GUE1E9MIZU4Ej/iS9XNXe72yhUDydXhr8XRHQTzjdqRMN+VhphTM/5JmZ2E8Sf7a38qci3kn7H
HJJFjcZd8Bd+tDEtMQ8dxnjSWOkG9biTk9j8FB4umKPb9k+unX6skz6hT1pTOfqPRLIPRVGo/63X
Bu5YVzHA4hX5yRQ4fJtYqzhv6iLB8cb8IDAqki5ow1DDvUUGBhCDiMAubcLhzvaK3KpUnOoeaxRL
WNsSjfhhDzuhnTP4U9zUfxu/VZvRCJPs55wOH6CZ2RMl51sTqtYiDtyyVoXjokOK7qGwBID4BLKJ
JmF25HmQ8oEYa2bOz7sBiDDUFtFhEn7kbdK3A8FpcSNwogmI77Wumcx502Zg2903Jjz2tiQHQa+R
ueoKCqMucmZAhtF6/Xy9PMSw3VlJxxmdGmbmtDKioOX5r9tnW3BVFjFKRUjhMfoD1Kvz1eXnJJqL
7zhJ93Dhnocx/aD41pjuZBY60EbTSPUFYf0nWGyuCQfzH5mXNO7Ffyn0ZlHC1kmZqcSef+L/A9TL
LlkK4A5rMRS3EUpaM2K2JpB+BfNokQOwX2wVtlxIt5ktlIpiIojj/ksZYFCvM2xTv88TQ5WGwiV7
2L9sMQ0aeIkJ2uUByKiVnCm5IelCK/8F1qULqNp6DWUinv1loOjvbv2FgqENg0OekwdSbrjtcAcz
TKABnz97kU6UdotkNF+DB9R7heN3S8Tu151LAheMcfI3SCkouZlyWt9Ovr3Pd83YW+OsoePLATOu
qH/I4H6Ezc4i0+7dixm6+r7hvtnCwdra3QVLfPBmQFO44V7Vv1+AswkAR+iBWbdIhfeMfMNfSk4j
FGtP+YZH5R+6N680F+BKBJ0Lg10Zt/k3y6qEJEblEg6MtRbq2koETMEVvohF5o1Lwy7nbCsU2Gs4
z81MBeue5cg4RTvIQ5Mxl4oCPmsWLcBbywRM08VBQt6siRxn3JntwuvjHb7hja9CxNz/ijKXYeLt
64cLqTRGIMS4vMJXpimF9A9RUjdpgHdk5/L79/hAp/pRqbBLqZnV30N8sMwinqWWV97mj3huHkVF
HA3hfp2Yhkl/uW4t7fgyiS0A2ly8COoR8O645CxN+XXg0v7ARoF+cWgZaUmyRbDSgKyepkulB73T
OIzjRXt4tPr0i4DrUYhQrEa2Lo7Yp99r8HcNg1RUAlxKkPZNf3rzpXFMiST+B+Iv/qRyQ5Orod6N
ba/YSWM+4gL8XfR3YnV7xPAiS5T6tGVv1Z+CoxoGdM3erHtpIWNkJZz0egtdSGLSWVER6u4GW/Fs
B1ORpbntngTy3zOfl08tO2Ml3ONh4rxTEDZ3wLeVBg9KY0X47rXtmyy6Af2zvNYnzoT2+kqFgqtp
3WF9Pqma4kOrRRr6mxNUnbpWOzOeqnP8knveirCCTsoEWGgBviDFx1Jgkn2oWhpAObFt1OEkNasX
Ql3DEfibGAFM1DgItUOgR2Y6/UHLygEv37x92jyAfrpptBaKu5gtjWbB8Z/MrpaNSmuQXFSZNEJG
nRNdUNu29I53n5CoaDdErBvkxEzT7FVugzyjQ2pog5I1Sb8za/LuCnxGjN9YizVvAliO576RFME5
W4FcffZgZR2M4lwez3X/UeNofz4hJiyzPCeizoRi0vLgD59UymCe4EjVZK+BSSRGRGGq2nYqcOAt
bmXIE/HhPVZY9YrdspjJrtNEVgsOYiMED+lBD8EqKt5tktwhf4b5jMcYK/gVo1y2rDJbXe7KfJTH
mAQPGfsaYC/GkKzCtj+MK9FXpxlMZQuA5/E8wWU4lwyYth39VlFiBXDl5TCGMW8xIj5PA/5nYX5M
rcqlczxuFWOijQFuPBi0BWeXk1NSJmUjRihrLaS4hRphtEhmR6+nT3XN6yYYSukyIolKDYiNUJcL
LZFZkOSzGIL35eSOp8PPZbRZeQcL75BMeYHTT0kTDAxSJmcxqicRiMZubQ0h3hvIZeVQwCGRF3t+
dQrF48q4ERMYWj52cnsDfbbx3OqOPt96ANe4Ut7Bx3wW1KuFakJ9MWcg4QdXENuNZl9D8i0mWCRC
BENXdG7XdT9SxrsWejEkQkGQ3g41D1dm50RKPwqpo/EYYwaHBFV/SGw9UadQdp//BHYfh7wubbv7
OlE9PcmEV/5tiyMH7XRCHRl1+wA6nXFzjXaR6uwBC3EGdVNKMnkJYn3juvtj2+GuT2ydKaOOhn8X
rpCIuf0QNvgx+2IAkRQWnEAJhOBQHWcKscis4K1SOMJ/K+Q5rmeUxeyYcVlo1x+Sd7YztLlb7+l6
qlW8Pq4BgDDkRhIGidRXBmvO6lTHq4vV0qvc8xRn0qCmbiHWwD0MrRZO5hm/UAT8QkN2avklMSvH
BztxDJoM6Gqbioh3qlPQylCwfIpePOCiPB+xCS0ocFwQ5S66PvYs5eOyxi3UHlIZgm8nSKmeWnvS
xqHfJXwYwIg8ZUf3sgMyioqdum8IZweTDtQLPfzk9xjxRtqpeokqW8SZbfXWQI1Jh69zWn84SkPv
rCfas/E06mbEhimCd+2GseN79h9fzgMf5yB2a3KI+6LaDXQSNOAaS0xSc35n/QiL8uPJqVupQHm6
qvXH/pFkbobzw/a39dbgHQX0wInjsmUb6VRAEOJaaVZXYyq6X24gRQhhzfyc6i3g5NusO9p54GFf
iFGY1XG/gV+fR1ujTubd0a395BkXwCXwGoqMBfJnbZALcpD+i+TfXrqhjMJSaGqAFDlPcfeWAROw
0yRipMqg3R8czIxBeIKS1POleC7vD+/1dobs/6mN02KkZtP5222jCqZB84iJZEf3lIntf0fdjg3p
AyGuCMp5iAA5EMyrMwXeQPH9/DN9VCR5oyS5iQsbVQOoviRQXZ/62pX/Jz7W+fQ5ep3laZkDRIZh
szkc9vPFH+KqxSGOlfYrujVVgEFY+BQ1+CPH2+x0S3B3nS3ZusC4egfBjIh3P2kXSIgz1AJroqXG
FJ81RelzWNMrBmb5RUaLmvWQXzF2NW7SiXt0XaFb1FairS1/COOSABp00gwalY1Mxa1VWE9F9PTa
hzlEqnYXUj+tbM3bO6uCycNvZm17/9KDNVLmFYT7xbxqq+J9pYlaxmgiLSBu5z5caznkWGkLACSB
MuqdUfeWE3f+sTyXSRG496NOv0REtT/JvyG48xzuRLqq8KjVzZWJzEgr84uI18KR1gy6AOEGPwHl
mOO/t9j0btSvAMHTXBJskfE+u12868Q4E1uKIqjjGfovFxbi1xgJujEHjSobJy/npSPdNtcmtXA5
w5ugJm6+np9UYAmGkQHAgEaVoL0lQStGZiXgUjuVYsGJ20noLXOLmzP9VpZ7vbW3o8vKMBhzpNo6
+TIbqluBIj+vzY+8DbFAWXjl12K2lOftKOfj9O8vdtqNAzdxU9WQztDisNG0/ua2B4RRhS+hQ4Ws
pFnm3Hqjjh8oesvc5t+ho+/3e7dE5TqHpTboJclh2/KTvc2bUkAsiQra1BgAe6pBIvgeL/OHh1h+
dEtFEWXKTl9GdI9ZsGQ33L8mqPOx6FEqVU0GuNpPGmcP+EN6czJ0uH9oGFrPAMWIaXygNWxxzPBJ
sQwOrKj0GBXT3DRKJDaBuVLpX9bB0KpXE6DRu4koD2JvPKfTiX5wBCllaHFG3MrJkquy8dOqxgCt
t+Ufsja4yZz0vQeAj+Nce3SrtdXWCTedI4shgMESywWPAASVl5RYCk8eizUp9dSn6mrnEEGfexMV
GaiQjq0x4B04d6x2PDo20YtCUqh1hgzhl/sDyFWN0YV1XnmO3lIy8vMwFN4Uj0tV8gc1Z9dgnrKV
KDeLdID01+NVK6XMWYggJbtl7a5K7QfzhvjzYZxkwuD0GiaikeTnorMBGEAM2QPv0mIa0hvEGCs8
ut/3APZvGx1Lt1p125scN8knVu8Ks9j39TzM2ejlp9aFcuXs6ti7e3oQfX6xcCyUUOj3vnrt7lxe
5CJT8DdViQuMUIAoExGF7aoGlCOoztn3z0g+vrkKWmw23RgGyXtVptN8hq3sXxTd1d2JKBpZmSK4
IQX+JqoXGdJVibYLIUDxXuobnwYxBpy3sAIkqMGucOWSEE64+9DiZISxqX5mRa1rfmYhjVzaB/l4
k89ryQhnavGwrTVAodvVmzwV9N84WQDsHosJSnC2EBnE9lcCphEBrZHyXkejbmtHW0DGqUpJd2Lk
anUeEwndgnsi37fSfYN6IxSGqDlWeGoC6zYQV2Wwidn8lTOIO6rOhlJkqDqXTmbVALeosWFC3p9E
UwOK7Pp92Y6eFud1UAb1B8J1twe8iYgsJ6PGCIRtRiafQ3sHGqHaM0+N4EKRPaLHwWOQ1pJFsiqU
N8xoFNe0d1HAlkEdTHKhaSYCU3WzrOCb4jLhkyBLESVguC29dMQj1dMrFfIpTr5mJNEBNqrSaUjK
QQYBmRe6i78K6/JqyBT2Z9csDFn3Va3iu6LwJ98X+OL4zgOw6Zwt59FCjaqSfsignq0HElbPMrrC
9TDpwya3n86LteSyoAnrDOWKpMU/IYX5uIuNQF8LjbTU65GLLL+dcyJ5Y2zt8dDi0Gn6DXFWLU6R
0CMIHj+OmekxE5zV83l3pBzyEvnQd3+d8GLK2Fc9yxvDUuViyK3d9V8QyCoWrAlMuW4tlxoKhtN3
yjammmPx9hcZhG0pzGlih+PFUC/RSepjvsXWBP6a4C5a5OGneNvAvZCV+y49SxmL0tLOpgo2opGH
SmwAvWiZs6Qhx8q03S4xZ0MrBhLf1T13qBbq9ksnL8A7dp717dOL9dSrHZEUAfmeQ4pNKW4MbZvk
xkrZd7S2FN4Qf289sH2qMedGw18cwg1Da9ImSUFHLjeznGZj2p6MgoOVSiUGzbGNq90b93uQtmhn
xJw6lBty4bM/yXZ9PRMdmYbhFvgT1abTPzD6M2Mp+UszZi8+f6R8XNbNU5DthwFvmUcDe9+mXZE4
/oMMSOMtufKIJ/op0YKejymjM+DX1EMqbOTCZwc75RLSEXMFptj9wXMzDi5BbQfmjEmzGZlhsUnB
qiRHiL+EwbgBGdmlBFu9+IuaDPKDb7I/X7SyeOqnd9pmP+y1lzz+tE4fTC+YJKENPLFfCPCgUIPg
Y2i1e5/qqVIlvX2RGqJfe3tw7Wl+aGkFJwPlemh/miWRzg411kOltOKHs+mp4niZxLYfqXnienPC
FGSTXnm5w11F0PSVB22PXZyu5G4PjIFxwctpP6mlBtEssLNmQZ3jWbNkSl56fiDI06aWtxv8ioVb
m34SoeFy34rzKIWcnphcdILYTAPru9j28asDZcCXjHEjV2Ugs+/If9XAKVG2Gg5Mrgty6pM4aEsA
AAPcF9aoDy0lNHLkXvHg8qLKGQ1+TiQO0TONCuGEmqJtVX5Ur6nf+P24pnueV4OyVQpGADDD9rhS
vVA9aDDJm7FW6nKL3oDRkrLjFyGhhDu5vBWo6lxibVDdVwG4PIHkrE5/7cFrFzViE2f5gv/Ope2z
pQI1e04NeYmI6iaMHlkun+o8is8sdja9RfobHNup2VzH15sIR9MU2bbP34ArOHF2uB8FItGh93fB
37E4o/zfDi/BBcczifsZvMou/pd4AiWeI3OXtmygwiFeXv8XobToC/c5/c6z4iRw/uhgGedoEDIl
e9Aij7G+OZIaGOi2xullXWvDe7SqIUt/fXQeSXUYCxqGPk9whCiOQ/85eJ86bDfK+Oo6tLZYk3c8
VaU2Lfm1sKA8TPCS71q60EtHgKdLp5WZFEKj8mcqEt7VaowDyoYzCHfs99e0hNYPeanI7IumqCtU
BsN4gJ/JqrCsHoOoDQigBfkaplnc6Vdu2pKvb/v8h+rxp/72B12bKiaQXGU47wAm1OhU2MVFYa/Y
BBqqNnS1fpyBWB5Y4RqBwnHFoe7m6VW3y65tgrLXHceSnsn6JZHt+pGc9C7abaCRocvZxkWuLHKe
fI7dDqDlUwYr8me4GE8cruSGtExA3z9mmYztibE5JjNXvTqJrbvtdoUbR2XNXI5N98mrE7DAVeYa
va5b1ebfgQfKqazykFhyFFTBfp5xds8bRvmrE5VnHYxCFwQdn+xOs3hCVHkbh10TGgUKtvIkc3C6
QkTmpxEjGiEDZQXAsHZFN6IyLoflaq5eUzoxQa2QtlBS63L8eify1pjmtU1szClylddqWXTRBkqT
hWadWiXIbRzyknzgfC9Mnf79kDR2WqC/ANKVGKOZWwV3kwb9k3Vl63QtzD3DUiFWyxWwzrNaeZm6
Q2BCFsYMaRgHdE9mytfzz4ubYKLTTpbJdoTf64zVUqLzreJnO7WtQsIcTU3/dql81QVm/yfv2bzi
x2TaZmhC0vpOZwVHKObj48nunvYdRPkf7ux9Dn/dn7g1oxXbLgfobvQAAwqvNprNt1NPcPob2FIa
H0xdDIC0FWSezDHY6ovHD2enUhCQx+L/ZuJDW1FOIUOAcFq8BoYRInupHOBmZYNaqCg/GZuVpGZP
9fKcsaycTmcc0DYOXelYoXEBdJ/v1TSdxiUdFl/3ICOxE1/pxBO0MWVrPt+rUCCO4mW5S1PTZ7Iy
30XoU+HBbIjreR6qlFAb3LJFGOboQTizbLM5KtjqiLrARYT+6YZRBbY5gBN4QdkFqbynloDk9o5w
+3sKJNfoE5iYG8yGL71LINiCXFVqAOkBVO/DI32i7aQOzHRRWxkdUzFzGNhBi1x3p8H6rP4Ixt6b
rtXbDEDkNTDGW3JRQdtZZbMzUMMg5QjAFwpk+7kqz6hj5jal67b/IX1673reptvaVwUkf4yt3woF
KGOT47x3TFebF3xGfJDbegi751FymwMeU9CdHPzNqKMqMJ+f6sGKX/47/rfz3vVHTYkErkUv+1Ck
EOnIlcTf4oUZ7CSSWfKQM8X1aSNsMDGbALNSaQ1MyfqaGDvj6YdOvt8bh/gKFwoiFQjN7w8iXY9C
/CzThU1da0AUHeZtZ6llNu5FNWXFADnc0m+SO0ewz52JDh7sAphf1g3OToaKqzoSXKx3BbsvR5VZ
tL8Vvs4o4o5xPe6FUbIA0m35+o/LiDOMzVbRY4bQ42URnGrwzB/qMpUQmmql/puYzC4Cl4VOXzvg
u66fYGQte3bkJmgaLNG76IeK4W2rd1nTkmvjSBlQEQqJN6dC2OBwCMOc/iMvATK4FMR0Gm2aJD3p
PoPh1bCVSNw3fmxjorzx81a/SVNc85AczDt3dCwNg17X2d9jNQwljILsA3rR1AAZaYLix9hIyVoM
ZMmpvm6sqRqVFhkCwgJLprGum9nsJg7QeoqyqDbzHZ52oOuzF1aALA2X4V9Vn9dpo7+x91xWzwTs
hNhTOUsB1dYtVIOmg8sgPhkpEcrezk4H3HAiqmEgJ7eEY94iiamu+lVHHzpzTqkeym60Oa8mG6CB
6zXhTJ/uIEkjVbO6qknGAqjyM8svHtqAdp6Yp9E7sYn7B1PCZ6g0szltlOXQY+9iaO9Iz21Z1qAC
fgaL8y84R8H/lBbKey1oob0j0G8hajxLtNMPgt4h0rVVgvQHMNptf+URIawNiyRr8z6ExJoYpcIN
pR6g4c0+tS2eaQ5Jy7c4XU+Aee9ZZHAT5m+hW+2wXpTHrBPOgRR0UkOHafvn4/LC7OuO5eL10k/u
1+wplNjS4j2/MSPs9hhuXc2yn6KpCc4ac3LcXB7UTGe6RaYp2jLjcnP4IzBfhba6Vb8JzeiT4aX9
uPyqZA+ureFP/GTwO3r3jmuPQqflq1ENZx+55fjTpFmxQ0Qb+wJDNgRJ5e2u+UGCJRuNxrxT9o3U
dz5q6ObkqZZVjlTzZ6C7QjYzUaVNakX0KMIupw3dqo3e7SuP0CY9pcCfZJehlgL/5DxujBb7Kmsb
k4iPQkNzniOFtrHyIkiA6NMCeiGRlOYSFikGvo4jwPorBReDkroqsespWXLRtxSAUYlX+NsXE2vl
UkUVLQnd61QHmhFdKTlgamC9IT65zGltxjzSAjLhFDnHyckyF1s450JiR8fUKYkuhce1iFRqGb76
IOjaeWMG0mBKqyYIPrI029pz5ivAoT1+lCUi/1I6aAFJOg8LzzuKoFPi+gMVwZW9E3TVRXqmATvd
CAiRNLOzW4IQQbzYWZnbZEQzYPZvP62JMMggazpbNWFnlW69THJjXJftpkQAs2S/qYgCadCRJxmA
K6mDoqVUHwlVUYgMf4qHzRb627Lx8y+eTJP6agDHq5L5BAdwF+ucERVEbLKy9lvxr9bvGbvgU9de
m7LHJlMJpjdm3xqtorpQkIzoSB4pJdWu2HCnxiicQahkfmZlhFSF1toqz6HoQcICh8SXnSOMonM2
J4jdKvAFvKpBtiwvs9O2ppJj2CjD6eRNFhXe6fV37/n0feWpmRWYOptB8tnZQXubqV90GK9cE0eZ
4NeEfkfD8Zel/gvTdNLf1k1j8IQDXtvfbp0bxTROxuNJeXB4X9lpDeHhk54YLU/YAWCzz9khQcGJ
W6nSt32I5JRu1p14cZNxybhWnZ6Y844y09c0WUajDKs4ZUyde6SVd4+uer/9N3aN2iNT7fLpvPaN
rON6BeYyZkj7dHlgRmYM97PmbnTrwhsHV+fr07IIVSdHMx9mGnbB1gs22wWoQdqk2Qjq0ofe4U7E
wJsVKLq7Gr6Tmnpxf80PpNfm1Q99XYrmVerKOXYolydvwJZfLQPLaIcj9b01fdG1e11ayrTgPo0N
VZsXJY3EVnalb6Kj2iFgvaubBsuIeTTHl/hFfnxZXhLLBvuAHnPVqf1VulRZL/p3XB7Gxa7cT8V5
I01VLCuArzir2S1zqdA9fyLxJEsrOq5zNnuJlOHooBSU1u0RUYYnbW9pRdYx+xr4430FO5e6a1UQ
CKUmymazZOGE6uZP/dWd0sqOAeJ+vm+tFSyndV3/dsFzIorKKvekarFvT0PyzApAWjkB4p2wa2ri
nu/fs/zLCWTg5J63BzcjuTSx3wWMGUVQu4gYCwPfaFH5u7RVUJA8qsKoINWZWY5JghbOUyhN/tjc
DRRIbtytmyrYFupvs8xnmfMY6UV88YKbI08MOdvZ6s4+pn+T10e3VOKDVDqAVbgCD404eIbZOxx8
WVxDphv3yyDoFoBSpkBvMXzWgrz0JICGgh9Dax5nnNj+1vdT/0SmYbUiSiETIJUy8WrguLXRIJal
RSY2uFHuwYoB6ngCNek2qBY249GNxFOcRDb+B67T48Kp6T98FVv8WRvSt1FweCh+qbJLtSwhW/HD
NjvMjAkHBXUrZUniBlv267hRFjRMOugumF6Kegyh4ihCb44ZuFgU6zpO73VIXs/Yws6hFI0fIGaU
SHBK3kG7957wttM+u3ThfEc8Sk+OQ3Z2QwY1kORq9lS6uZb5AOjZ1hK/TTor16WTLmn7tw4pxPDo
ySBxXcFtZAZztpM+g4EilsjPs+b/ZGRNMMk1kBBsf6Cm3DjzfcRuvzxmts0I7gFvL4tXJnpw/Rjg
B/pKgmf15V1dtK4CCo8QgUuOLWRddZVwuRi//TVplDR/4mUF4f4MN88/lb12ecn/DfUZq+MbK3Ns
oDckQw78fVmnL0/MxYLPrWqCHhVjYhbBN9LwQ/wAlMSEd3DbNpLFTZs3/nDrCvNWGwBwl/tLIa8t
6M/Zw916/6SqCg76QhQ+Ve0r8ROSf4VDmRa9FhnEKdpH9tP3xf1X/Woz5bVOnzU6Lh+oEM4AWF6T
QiOUJJ35Ud6GNXqMvR3+nQ0v2xa8dmoJxJmXQRoP4OCh1rqvhf1ljqJrUIE+Apb5o7IkzdG3zP3c
5TXtMckphCWhNzxlzwl+eOiy2ftyxyhg0Y+Pmj4fLVeDX1JMCbV8b0XzKK6VKara7705Jr2tNHkC
pSQQKcKxMP7ISmnJlUPh6tG4JqvgezL6fgECrhiy6yOXYb6WRctDvNJjiYZTRVTW4CEGCD+Lqh70
B/VY6k9IghQabN5rCtOEs4LWagKPc01bAO5uq0S/WOWbqLKodcIz5Tc6Ky8CPjmh55NZ07q7CMG3
U4wQTKgLYjVHbTmDStGCFp4psy87nEDzpwW0ePBls1Tl90mI1rT7T/4/tbXhW81k16UDWeORprk6
7TEQ0AQyXgzno8X4ogCG6N0zLwltfBvq/g/Y72OKTTQTj9bjv6IDEON0VNLlnuvsTpNZpAVeXY3t
YRlVd5/1OHn+Q5nqerb8v8Ufuzib0luuSdSLbd0O1UoVrcYPqhVorjsPVOybCQOXMySZmPLQwQjH
mDk8kSuP9ZLX/apu+89GeJO+KqNDSwpEjElOr1ShazehcfUfwlWhUECgl/YdFeSizYMF6KVKbYF0
AT8ZvrP1ULgaCF9fYMLfd921VKA2bnCX6WVGoXHehBLG/ZZb7HYU5IoejLuTxEE5dDP/obUgYjrb
DbMlaWkWFmPJJ4DxfoiUIgskiXynitz2PDj1sqfvDLH1+2O1d2nBDiWrMpDgybdRl9G9laB9mSW5
D6PsdcW028TOmJ7tAN5E/sS5M+aiCSrhObJqf8T/5TqFq5YMtES1Zpp+kIPi/+zPguBFifqZ1U7Y
7/6xOJ3IxGoqohoJx0RzlZ3wtYn753D0u7vKVKVzNGzGAHWVQS6Ku1bPgqH+gxnKravpP8Gk5VFE
NvqMUj7OLLIvFPogPiRs9hjLCzXgKQxB7AmK4yQ6wU3klKxj+zQ8izPYWrn87yw0E4n9SFKjG957
Rot0qoWZ7JNg2ZIgSG6W2lJv9S7JdzUOeWyMED/8GPsvtUoBFeH9A6/TdHi01p02kQgClRX7kQJ9
dg5l9MQbYc2dMDj2GmwiZBpB8RM8myKZJwAfI33jjm//24cd6aOnRkGq+3k5YCG7h6Serz9Zckx1
j/RjbtdP4vBQohGpZDWuiNMBF9h67LU2C67XftR/RzTaCpukXJe1OkcwWtKM9Lnd5MYzWp1Lg+Vz
JNGH01fSR66XQC0axLLj05+7Grfz0X8mIpn/jvcO+8XjaNZUc9xXNjrBLAwjGHVlk6lIj9eRi+GQ
skpouDqrOOsba8Pho7F6G1kK4Gshxf1kHt9eYRRKhPm8q8KYARkmbFs73oQUlLc3ZLBxVzeI3Rm3
oe5VKyMhTbz9K+aQwR+AHaZee+F3hDZXg8VG64TmYnADkYbRoOzwnhX71mtVVPiIGvUnAW5pHFhm
RsEXpXMgbtAsgs8Dr0596WvXda6A9IXfzYtgNQJQj1aGNfbGIMZIVfrbhumfHld7IG8PfeECDqGG
YDjGJ0PxTBFpaK3IDVbxvRivUdJ5qkDURVKyCr7De3KS/9evBJL344UeaPmXEcpDK+gpKmBUoqe5
pNnbPtm6kfB/0p0yMCrsi9XzvRiXiMo6aOxjmEEkJpNDfVnYZEnYY0uW8Uf7C7vuprIOg1MIVcU4
TB2BA4PF28+nlVodlnIz7x5Y0EG7VeBcJS64vWitCPt2otk4I8lABrELmY16ba+ISqUd0teiJWSF
MkqCw1Iq8vLgoAUzpjVo2oyR7683dMkLk5C6BEwN3pUTGMkaXYd/b3ja1mcgw6aSN4GdBqMEf0tm
mZBXhSutLhp6L5bIun1skDRcekYodydAMDlCgmp8WPGjDw5TtfaJJpBT1QTvAa4su467h0uDW+Fy
2IPZsluHhcjIYuohZ2YLrLjvfOYhPmZALjmPkDXhcxMr50rNrFLKq3J9dnbf2Y08MQiMgsoXFNqN
EFCrEX8I3cnVh2rpyqVNXgDWv1MEyUKCirp4wSK+RXSgxLxoOxeR/8dAXanHtnk4+AsUoqZC911j
8+Oa74LVyRVhaBAmKB39WGzm/bvwr3dm04GFbHK2c7XvVVmSmTAiU94VuLMyyDjp8MeLYIkkjp9k
njzqNL42qsqRj4vUWAh9scnJuZ4ALcmX/IXH/5s3gUrnu+everALTmkBAtHeBxcSIw3ACiPxKrPG
pTa4PKthCFxxmDdyIkGGN4TWenxsBRE0NtWVl3YWQZ2PH1PV1oZjt7aGkUrp/plsi9dwEmbMRrrl
tLMtyK2cDm4RgQGvG274ASgM4GDOC5uC3pOqMI8MPI1xvjUbRS5j1n2aXT3N2k1OQO2lR/IPPiA5
Dxou9tjH17oklnZMCdjBvYTIR5tHuDbLpp2hEWFxQDt1g70e5v+jrlDoPtNztlWJ/yDsVv0NBkch
RTv9iNGuaah/0D5CXPrygEc3h0wt7VGtdgY+tRBdSmxfwt/hzpbCOt2HDEyFbQXQi00xi0Rqlt7F
HQB7671NiN4nHK/VCRbFIQgaSx3rsEUCwo7yqWuj6v2vOp3vrWupSteoJUqAjGoAmGR+Tm8hBHF+
84M2ub57o6biwJwF25hqiScKUxvUi7AUCG0I3Y0TJJtHKg84Rql2520sjwGTnTXJ3I3w3YkLuOca
rcFMpfz8IjIqcPwmOOe/UNK4YQRmcqLyD2rjbhv8u2LMpdo+VMfv2TznJRzJAmIFInj/3hQuucan
WXq1L+vsrH3AzURbmJ049YlbCXkYsqlStfZfxG/8JVYXFCQoz/mD2DpNaQrw2nu/wVSv32RyEp+O
b8vEnvybmlTFijJ9VhrLtrUHHQuoeaO+MxKWgC66xEt3bjZ8NgwVhKZ/eZibGmB91V+kqH3egFLK
Xcz3Y0SowuImn0ZkX9IG7EUM+mQN2U0vlAyU7GCV72z1Vsatr8seJROPXbP7pNny/LnDYt0i4/O2
obKM7HFCxelbiS/ewOlNePvpjfVSmJKdu7bQmp80BXQ0TFejb0iG2cUcEZm9uhHjqSSX1l1Mqns+
KhZcDD1YqaTb4qQTVBwdCbxTkg1FjF+NgfeOZAfiR/DE/n/+y+vJNUOWL4/uETsXopVK8rh3U0+Z
W819pfRHjS/77jPQ+qf7arZZlM0ZjbZZothtYT3UXGC9fB57WPe1HX6owM+Vr9VUKZDlQntB9r0Q
4zk979FZpUcxxcyxTnw1mNwJsAT/7LP7L+R2L2NqAVIYua+9CBvHSRtst0X1NfOi+0vBJLtkU41p
6Y7JZpT8cjJy+czGDS18yiD7Ifq8Vob31C3cLtzzYqCsdIQm1CTgzMak5pMrxkaFB4xfAZV5NWgS
/omfdMBrFnipkAUH4Ix75gm0+U73EMzhNELgAfzt32OuGgs9OBaXPDwm1VQ1ZwhcLYZnmvI/G55n
z7VmTuXwmVDRCCwHCRRw2ZVt/z7qHPVMHpgYGyWtzZFee7AkF0S+31Wy7xg2w2ID9sgriheIqJ1x
CmBphv24BpBiWsfhA58haLU5rRzy2MAavTeWXllzBU6uCQx/QB0phovJpeCN3TGdJxmqD/sDHjYX
9zzjcmhFO7JUEVxjnwbct44CNB7vICY0DvywWqRJb21Xp9rTRiZVNthXqqseSQIL6fxj+O3vXnp4
ilqgCn/+6d9XlLTZoivBxyJYfTXes11OSmdVL91NTWgb8fMR1+PYFiC5teaazgELYnwGYwSVr6Lk
dlBUihVKsZhMAWqQxAdR9KZIUyc5xreXZsC5RQX1UFEB7RfAHXD9t5GVTg/NtCvjU8at27++lefU
iDyxhv9SFcwAHDdBm1FlUl1RoeTaeflq39O7m27PuPrYDoznaaeb25BhfIXIFAXJODOpKnoS88t+
fPlM4Nef8KZ95WEWNJ8AcezAGeZRlee+gmMYqTP54sEYc7I/jvZi30DKW0bXTiYbOshl4jgC6tTB
VbtbAYQ5Zb4ZDuVEyWbi9I6A4NCH1alakaD1Xe0zMvh1UFVoXTCacKJ/VqpTxMKYajCRntGjs6AK
iKY4hFHl1T44s/X8v2whUb3VIPmmo5ks2i/jM5i5TycnxO93KUiY//Cr4t6G5it/7ub6D9Cgzr58
Z4Nwp8pTfdl2tFclNEsMgZuCPixGO9RhB9aUwblEbhNlGSe/w7VtLmhxxqbI4peB1UI3bJHOVCwP
JE8dzow2yvEpsFr2qnPIs7r5D3XapchRyCkDtANt+iYLHB0cfZ8A066tRwDg6LPr0vuZVg/Cqoml
DGSIitltNBHXz/bF47sOjTFMy74f5byNbLc49VOFKFe1MawqJmp9X7pnuFNbOyqOLkiYUjQWmxLk
vApedI+g28Tio/vx+OCYFDekzmalkCrr3p8w9IPNxt9eHOEM1G8RkfQ3KyOPnpoQUa7UOBEGikKb
yBAcFpTI1ed3vymaR0Abp80DzApvfY6+PGFd2U8R73YGYlpow2Jv/zq+G8yN7QlEPk+UZ76JlRko
UC6VJDTB/Y8cbQ3fhEyGFxGb5SiOiYCKsWuQVwVCKUEkmPXp0rYMR1nAeXtiC7vZvPex43ny3Cu0
9wjzZedk6c24x7Xb+jVcAjDc5QZ7dPp0Ne13blYU8PJL+TTMSmTllQnkve1mI3fdC1FjDsuWPbIv
Cs2h+aSIFoI0j2PyCcYomuHLucIOkAwTL7b9CCENPkiOXpFKq1KDjGMKudNGk8tsYBvZ5aOR4z+Q
0Ybemm8tVdru2oZmPcATYjawoEdPXQ4eldrM9IX0lk+PCLsZNdDvWQD6+Gtr0R6PfdF74w+3+oda
v0GRLp7W306koouhZQVizccTNxWCaSn1VkrKDXl9y4O8R/PQPyzN5HeNtf4wwIGRVkwbxKobxHva
+E+omE6AEfXpCvVPJDgToeZT7FWDa/67XCeQ8m0pLrq1zyBHz7EEgeGgmYDklpogQB/vuAwPTkVz
vNmmpm46Vtp+2s78zT2JNJlYcm8dQanIwbRO1yEC0YLl1yjce7Sxbz+ogHAMpoJFHUWXF1O9BRxW
s4bn5LunoGoIiaYsnNb7HL0c/GheubRxi/gvJvlRU0yN/i3kq0hT8yKnrEYUA4FwHUs+ymHXork3
6AOTtuMcdmYlg92IsnqYl6xhrmpHQ6iJsGkrs29CgXEuY+zhVki5XUgeWExuD+LwL3k8wW3AedCM
yqxy1EkI1JUhXLHtlwsBMmqGxSGgqOohbjvlO5gvkqpoOHVsGB/4VLURKIyNvHHum9R83PWcKYbQ
DTbRYV5RsgFkxigTTB7hHq5WvVhgtSWZapMZJ5Iu8U7drKBVNSQn47sibj20vuM5+krADnYHDSu+
su7axJqpko/shkwI/w3s8L2Ueef/nU0eWQ8oJRCV5jptisiGLsGOt5Tess3fGVGmknEZiCCB3DOA
acXAbtOx4mNnVg0Bf3A6mBzzVeArL27T7ZAZdChqX+0o/FvF4HNMiTj24GHDLMmy5wzcdevvFe8o
Zlb6MN0CngWk3Vg27DqX0Jd3ZIaqY5YHcSz2hqPdVLlviN0lM79VV9GnVmmyKQ0hal3A9S2S4l4F
nfnOP+YadXTtOKNWtSuToYoQe6rCQMBsNasGKBd7sr8rXCnn6nzpUAPCd+n+RjtVvdFpb8KrzxL8
5uc80auy8aWio/w+ZxjZAytlvn+kpIO9bregRX0qH2q7wYvFQQ2T+btlaYpdLHH3JT0cmcu3LvYG
DcgoOeWqS2KymlBHwzFg4rthY7S/1J17cmaF5rTIjDopPIZfVjG7uwU7dZynTbTwbeSd8elhuoJg
XNuSEnH+ydaJjIxFIGGnj+gOFwMI9AlN9cP6kjSNUuDaTe+2eAFMyP00/Q1SFFhnrLshtK0S6sPS
t4HMaRQ0f4ZImaIdzOlqu1Dp8XyyIbD4ga9NswBmqKcQSdS+urIVqwGVx8thOS2m9xCFkYABG9ki
Shq5GfcmonedxaoubbLgS/9nZmOb51S2ypbDjqXmeernr9Vt9WB8ArtpDSoAG8lqBHh0fzOX/tB5
0J+dpvduQSwqv/tH1KDrylNe2li1eFl2NFpYShjcy2XE/MDHdtp0u0DmY0kB5ky7LeeRmPvop9vS
KKDJ0OPQfuP6z3y+8mycGZ55nN9vnPipG/ORh8BDbXaZ9G1wi+0sFoapaW2c8ZelZg2u6c7sGYk9
iJgNc6x8T2Qir38VyLlYpXae8WcoTuR7iXpVzMEhVeruHf+jGw08GMULoQZiaLGfiLp/bzJT+xUf
qttbWTp6zGiTUASf40wFeAsftinJ+AHJ+YI4GboDgAJ7dREYKpTphQZyczrjS1ERMlk4QlO71d4p
HruYOxGggBkkq1h1DTFX71SsReBDTU+PvqbDp7PhVJlIDWnWc2DVylpfzAMh7pIAlz8WuPxsw51x
Xk75uIgg7XAByIn30bYmC4htUvz1xcrIHQNlJXCkPJIGLSLoo/CiehcZUXh/NjzxMjY4oobKcrKK
RI61ikE7yLnUtF8aMnbjyb8NUjRhmB+v4gpt8msIoRRZ2ZHm2zoXgzrkF3COWpSCaxypJ+GYAwF1
+4pSYvD0HDeh4OrCDTV0khITlBu2WmDFkTcElS9fl+Atis9EdkzME6YuPSDCgs2FHtnyLSY8sFDy
n4lJEBFn7tCyDtnKX0yMZuB98EDHijC9Lhzwmam/7Sz7XdQpAQzRIyYCVWpwien/wk3S40Xyy+mO
dL+NZc3oy72i3SiOrzQ1rYU4Q3mIRjiNyuDYDXrCxmuYsj3v+SdKkn87GV5iZKZXSZy8Maqi9toH
GwCF+VRvzVvNddYuosBK01q4krTR3KHpkeplh/xvkArL2DygqW/kUgMRrL8sFgek0x0g/tGczcJS
0O26LpLbn0h4VgpV11sG5xgZsxCZzVruozp/prvyWb+pxNBuOGWSkgr6Wg+9EMc7iyq724g8q1bx
xa0d1HCMVcEHa63yTw1JpMeQjiGuZJjXFIYVHIBcp70FYcFN3PJ6ltk3XkyMCcT6dldJWaolCGQa
1infSvPkT4vb4JyTS/4fTu4gpO3C0yUHkrPkoJOzogv73JEpltyN/UY2vMDAz0DQhReA4hWM6VWI
46NtZn1gdwvs0CLbsGtZc9iLCwjvxQbUc0RG/Y9gkpP3lL4MqpnmaYBIiyo+iWivzXd527g6MU67
PAgfkEhPZkQjsnPizec3cdkE1NTuS1p6w47qdAEOaP3i8xFJ2ZT7jfkZcwGhW1Vg8uqY8VWwnAdf
ha7c/5UNpbe12n+LyNBMCT4VJmueKGY2us+W2XiKwlior+dGZeuKwPxG5ZKB2FTviIZilT4tasAv
VYOyuj80gDmPAGR5jNLUAP37aVmgojiH6J3pXLBOGceQeTLF+oS6R9tuuc/NIAafj4SyKgf9Qi0D
27Rjer2BgCmLuh/jiI5NhNg2mfmWIJ1rIuVjK8Bu/OMjGETN9/JwTjEbpDj5/tjhtgtje6Y6GSfB
8csO+QoVebiVVB3TXk/YRbW9z5Bd1fZU67uOKdCCGZISRu2X79pRKUAmz8vFm7fIGOqrGQbOofGm
OQqCgq+ZAMtN08SNHIAzJhpPHrYoCUOsbODoNWMMGJA/GDWM8WwmonFnDaEvWWvlQAfoRBoSyJ1p
yBDqOGXQ4OMKkOE3uittxag3oJ4E/9ViZ/NwhHsRbtwFKX/t06WdScpjgJ1vgsu5D+6PMAXeGMTr
Lx0rvVMCWasgvHh5odPgg+wiVRD8e+LOMVAupGrm1vNoR/IwZjEdT49aOxnlgdh0RNxM4T6TP7tr
VMh36L4lGqpMuPWezMGgappmDlLsKotHe634hVxMdiRrT6J/XItX0dSS9rU4WOsxZWujf2MZASOC
ypB+fil4IFdtlu+7m5U6AMo/qCnNkq/kJG2pgi7mCeqqqzITn0o8OJvn8XdnAQH/01nBklnHc0cr
loqNc1Qh88C05PBLLzlJlXMzYUF7egy5kSczcECrs1XjpDakf4IkoJVZatDJtBh6BfEgQFjtejld
RaniKsNKoCG8aqqLR9UFdv+ebafsGsXKZOTsmREabAZl3VyIZLItCZFLLYNHPLE8MkzQfBOYSgmb
fII71MGoudzxs3ykqT4oshWowx6Xh6sNW01FhOOF/WLXF+MajLROcpl3MotKpqWq7+3DJMqQWYS1
Mw7mHYgcwaGNkvBlWcQg5ojFET2lprybPuNEfbn1y3ob/TWihQIBbBzPpAZDcWqtaoiZMfrYSO6d
r80g6SZq9rxZG0/GC6Bk/oWlwgoH0Dgvzs6fq15L+wPBaYjtbjSUk2qjYLDCYY52bSdm37wCCzsS
kqixx0MHvKNR5ogmtYUN8VI89F02hS2R62RLDqQyGvMMw+RvBM3eGK5kl5UkXhpIBnlYA5TyMxDq
SH8q74HgbU3W5do7Jl1qeJMYwpa+xDTHQB42q+IygZY9mlXQcjrjR4ei/mfJHEg73k3WANFMl2tL
m2FNnsuIOPDXlAFiuZqNdRhxY7porOTafDNrmEv+UZsxMXp46hAWLc/DY5eSyNqrxoC/jgz31ZkM
GMjNDpgYRh58sB4ZWM9OwPNhn8W+oYHSGqqcoHDZclNZBLlaNp/8vlmBjFJ7XmS0OAQ5tbRPLwKB
QorpseXBwN+N4EJibNpLcRHP73tGG19MjEkTHidruRDyUTxavaT6jLIkZbaN/M0cGOks3tY97TDM
aghYb/z7/MjU/a0i2i2SQw/In89Ymz2o2MKsuIOZ7icVahj5lsZgbGHNzdAuTO0HdGWt+g3yAEQq
W8xG1Saa+nfG3dQFs7liAharnFsEYURNIWKwx6diOgRm9HiovQ9cXkMMBC9pXHqOhvy5cNir+7ad
KKZ8SALTJLW+gY1+BLJKIEkr49PEryERuPt/qVg+iCR6IcdKil7a3prS/zRQZpzbSlhC27an1ygz
lJXZvcYkWB/yJdP8AVkVZB8YTVTub7cUV4xgm+esMhCkeQvb1wlpYz+IZ3Kfo2Ofize4icVIU6kX
wg92b/1yr6o5r2kEk4jBz7XIhVCAX2TNRjZKllZMuJZUiyhjIV69ZWo7hLVmjicVXLS5JxKzQCxt
aiqNxnKhX78mruWhzmZTIka6LfOqFlPe5pylOwYl4DiLfWOWNZMl5XK8C0BnREbgZ3uWHAaPqgTo
vChDK2Nb8FaEoZzMVtdSpKcQZXuDmUbZO54cgvzh1jyDEJw6Er+GVhAxoMFoGDvlQ12cgZNjo/Ff
eSHugO2TB+mSqvEc46fUHLfeS+i4KCdwibvFYgG/im3mM1sE/RREP8babGlgS7fSwAuSo9MOph/A
NDDg+GknZC5FqMGeSCpbjlbGy9mZKBWnJZgmeuH+G4PwHlaUqG1Rc/EkKt+D02HzKmEPsNR5sle1
0/Wpo/1dHqS+WGDbGAaL6yTJ6NjlJhS4x17jiZVcG1JNGVAzsztzrtMj5nR2eu484ozqYvc6CyHY
n9AeuS3ZOhyGcaWXXdbm8aVRdMU4fQR3HgCNrAV6X3zfPrYO5u9joK7NfkvV7PU9MTmoQVtvdmyh
0tHQoxhSIwVP58ORwzwC9Frkw5ZpFQ/ie7q4z39PXfpSU2uj7SzdkHLUUqhMOHi+xP8AoyrZd2So
0Ae9I9MIH8HNQxzu5625ZazQPMdpjqDMUXF1W3xg49Se4WQLrAgy0hF88ldyQEbpwsNihUnbPa+A
YbO6cx8pqLap8rczkt2UYtT8Djusc7ZGIqU/CgLc+Vv4993WEmgneimmlE5zo9h003LJ+C6QQajr
Ej0wmG7QoADfUqNIyZnkb8FpLff4cD7aoxq+CXnBSrA7BqRC/wElZrt7h+qQz0eca7mdBdAGMi5S
9LJA5sM1bL9eTmMhAb8RX58ATWR3rs//kITjMkwhi8usN/TKcA6C5aE0iaDAi+Dk2yo4x1BKkIt1
APH5PHVng7ukO4GqCVrZrR/iJTrn+z0fStFpzJ99a1bM3VoWkFFnR7i5H7dqT944kxV1/5L8ZbLH
RmPhAcpU7Jk3FLiRR+GHtYHLflJGtJ8ERtPKi+jln9ft4nWlCfhUuGYaInS5JncFaGbBIx3zw1at
yiYQgQO/ayzq32cY5/zEApPldBI9O4ZPigo+Q7VOEiurnSq0XVdYD4gZz4K2Ej+h14AJfKiCKaNz
y24u4B0RtxDRs8ftlf32O8VqOfuVXhBFyrSs0snlxuEea5miaddNmpStOJBQf9ULK4g8xngWpi5X
8bfU+RRboZind68nUVOBPW1yuyewQiQY2lOFp2IFTrCtFd7cTINdeEiC3PCqMnuKNEqmf/j44yql
YqwmFWSOI4419PI8SkOuipONhiqrlI1cdzwBkmO1Vsrfsn3LAdKCiutlyTLSrQzI71DTh59g785W
FYLjU5QFCnmlfh7v79HkkYP2pLj2U3g8agaUsBZNBJGSdo2eYBBxPIO/1a31H+YcAPc2ea0HNFAr
3CyvgJcOqkyfE7sxpsO6+ZFOFIWr1tfB4gHw/UFonRoKx/mHnKKWdBGvAlnl0Ty4wLSGYCuOLAHd
9OnPBOPEZleDdIYORjMHLhohX9TDBzEFqFwKBuUhoE30C7WvKfAc/IeJ8VfIAqP7AEjGqDL8V4Bv
OdBaroL0TmgcPgTt0mLPkikd96s3U45SlUqej3nOY9oKQgehv+fzNVMglgHqjPtExq6S8l6i8ict
8pVM6CayqhqrIIZ59b027SYCV20Gi0ReSNBQV7Lemv8lUIxScXqDLyqukjoM8wJNzptmUlDNmNcy
v4YU2E3GlB+2Cb+SZNpMV194S+bmZywmCDqGcEhpi74pPPnhOYu7XcjAX50VgX/s5uQDDDU96jiK
QFyj7GUEdVsulckxI7CRxVzadE+bYqYqgxRsldyIQt9wg4BFZS8lHNjTI51x3McOhWWHNfD3G7j5
NNXoMPBunBp7T2a2hof94Mt7BJF22tJgAeqsWpdl5BXAMa6beFbMscGcKRSMy5eWoPJQJuHGp37T
/pgU7cvbJmL7Do3YPWhU2RFaipweKqM3dlKz84teATc31qRRBB7JPK5Lk2FlEJOS4waozm3h1Jud
jvcyCc2H9GEG8NeBBPnxNRkNZ+HZ+ZqG4uTSubKhWiEw71MGqCHeK9qUivNUSO7QK0LbOyi35KOI
uwwvOHfpoKJvFj9T4phZ6NkjfSpkhUE+bPmBxFTDODDh32ZMvWbCbGZpQDUqV0EtGlClDQtORiaE
SJwyJcZfoEdYDX/canFcF+hhChhoDp24jsI1SvY+ekUcjOc9pHkO5fNFIWEc3FmggvjF3LxYeG56
NOB1murwTWB3QRs+sNlXKuaoZVKOLkMIgZBiaVap7zTb6k1S/kEr2kH6EP+PQxt+axu6xJ9RGS47
CkWXaZ3DI2sb1OYgw4yexv9Cp9TsqxXU/0uK3SHG9PME2XQ2ER4WQ3kyWn7BgxQPStOeP/D9UVZN
3+jRJESl290UnUXtbHYTYyhTFKjHmDGAXmurg1TrB23RtKxBiDDpGSTYaUnqSQ0S3CnqeBvkS2MV
cDVyXA16Lq622RZSuRZp7KHVzL5Ddtm+PvR15DML7O8yIW7YW+iJc84Ox3QEjZnruqjgmCA7a+uh
x7Rg27XBgYbA3V6rd3zJFV7qmk9j8IPLQ7u1p/yKMOx1G7Wi0FjiJek3usD4eOZygwDfjqaDUI+G
ZPBUwupFn6D4RKdwn4iOqzEiEJBuSs1/foTtVTwdXznymuO11pUUj4Seev1I3F2UF/HzkDhdrVIu
X7lXS3FfbSlw3+TttP+vb9/n3z2R7sesQJB5fp5DwxgLbEW93703v+BI1hT0+9OOBumhieAh6QLT
3F+aAEhEWjGOq8gt/1mi6V2OC+bsX3B0ZqVilZ5etmT/pAWPjlfaT7I7VOG3dCuDVS7h3TjzSjD1
FFlITm5n14U2pvwNVWMdDHBI0qkDdnSkp4Df0eT7fYY1UeQT0JJjUyu0gWdpQGyLNP+y5MbThK0F
a3il5ioksyDo0e74Hq9fKRvi+vQ/174d0v2UjxkG1q3nuK7l2JvwY30xLQDvebJthY/bSUqgL4oC
xsxa/ctISParBVfH6YyldHQzNqRxfUd0ZsiKLYCcdgGOlhUxx2teXxlg/t8LtTuU6HLGpF+d+nYo
+joNXglpc5fMeceMdawd4DJP+JVgV9rjMfKFBMPXCGUaaKKvdE+yLmiKfI7OpeAsWoA93gGkuo+W
3U21W49DuC/cFWBBAU+llMCyYgoUvNUtMY5bACArFFgu9mvcdFtFabGfXLu++MnXe6ynuJQSSDbV
LcHMrbjJVUze/Nq1K2lWdXHQw0b38f0YlwEIntBqMcxubQ70uGE0HjOeDowjPtvlDMQEY/23RxSx
cG8hczad7bjCDlxSRD3aa05WwtpH+xv7sVGDtdFV2z30ovCIRhTXECbws6X2Fbt7dzmiSMxC/2AU
4ZN/f94MaJVQi6GW4V42bk9T4/yHgtQJTc1QdMnR4lc+RW85us9RMZ9JouDVBZrBe0I1dnCXKtNA
H/gbHtE6/2rL1+skOjo2U+l0qYK4kY9JDNjnBedAVPS3PBrtrimJcs7bqB3923xRW6ODuJ0qIXSi
HslZRd6tdD3sBBc9r6B1eATAmg12mu57rN2yIwxxib700ciXGqnoJZAg5ok7NnQ5qVqLRBtSTjqz
tYwRXFdqFpVwCRT3d7tD6uxsE/hYkiKVBT+Yxp8fycACEHSJiRyqQ/STYUBhfF76Lrjs9p75vKtJ
caqo01QhzpdWK6wy6pkHZ+gO961CJXHjitgaW8My00fKPtJwbz2ONwXLgbb7crXNHtqm1swwI9Ug
QwaWaJiMc4HIqGAI2d4i2tznZoxdizTAj99UY8vQb7jS96BGQLZrw+U3WKi9z5zwKX5PTvvDd87F
d7DHSh+pFcPs4hfN7KreUrN0gu/TRbdIgz5/xyj2aA5O/hXCIbmLhwEPMe4n1a5dusjfLpuakdgc
eMb+ZhrTGK5ZuJCBBkETDzvMLxR1Op5RFvmfLGT0htu4+3YS+GOam3T+eOmirhZVjc8h/3Bf7A6A
sjeqYHt3bRhK34GCpkEIXUL1TxUR08sqdwhad6R87RtDNvkQSe2NAMKadKNKeaJJJLR5m9oDfLLY
NFEJ7Y9BbkAGrbQaXq7ustw3nwhfwHTIJWdcvyDYS1s+xF54lp41t0KcMHepLq/51nJbHgm8Ckkw
CSN8BnrewiTL1AJAzBPpuWREpfVDqvULyevT1UG6cZdtZkG/qeXHabTptBFqfTiUURbowviBXiwV
D8I1hTYcseOqE022LEWgdwNLnCTih0xI/8ZS4hBH9D6kFBykBb7hJOdFR8sakLXVQRMwUMbicy3X
8svxRSZK26bQN+tAvoj+uU8gwIIgl/NPQIYSp02Cay0wN+UZlIKQ37HxHP01xwXFBctT9EU5ogT/
wr8aoUqmtGh79DT4LZLYb/YyldEV6hxu458GdkpYrFvhExkcTVdCMEQHgINKW7MhTr0HqgSjUKCM
p8DBB45wo8x9XFJVMG6/0nNePMIWIDf1XL4XvGbvh9Y95l1lX47VFT1I5wB2BUXntkL5mas9k0EE
LbGoLn/4UfbtDdD2ZcTcRwZECgRLMGWyBXn9BR4W99dAO4IIlMlvYK2JPq0LcGQBWT6NKKtwnjc/
lz0PGtTFFoHCXOvsOCfC0pbr6Lixw47wVFwtYAzTRYIO/lG8vkgKqlna1sVogYsfLH18+Ll/hP/X
JGe8KqiA5yuffOMkB8JXVHHF/ncQZwTe8iVH4zK3p/j5VIEI4PFGkkQ1bBqo/eMB+ufR24mVpwaa
CI6eyTY2pS9s/Z7EdC5FiYefk6pI4NW2GJbFA9YudCmibrZUHNs+e3gnokt5gAGMXeEZDTOg2uGD
Xb+SgiysfIyaFT7KiF62Ot8yjIhGe2E6p/CMnowtMAJ6HHD5XPhfSzC8g0Gky6fQJBMbb+NNNLH1
XWZjsOdfAojAYrkevR15BSynJvyNAHQtB59NyO+phzJQLA0jOreJQvq7CPNpvGZmw9gqM4WuDYkS
Zn3n9NST/3Z+E2AikN5mHNjSm+2ikzls8ZEyigXDrJokMoPNq+q7l0jJh1YIp8H6slGUBO1tBTs7
35ibshAeBAoX0LV/1zJzummshFLHp275T8GRCcEg7F4EmqmZU15qEi3f1UVAEqLH4B5eq3D5UqJo
pqQUnRoMWmXSYRHnuKaaz42jtRG4QC9MX5edYr4W0KZupdT1im/NH3Md+0C4VW2MSrJQJQbcVgb3
ypGZcf8ICnlmgipOQsd8W8IKCeAsnn46EmNZRMvcuuxHg3pY1JjXmnWlZeX4lBWSf19IGel6W7xR
3JfUqxtIbl3GJzrLo664wS+oEDOZ8lRTSKmfQahbI8hLxZbzpJvKD5duGU5bmeElMoLvhpDU8K7L
Rw3h6ALzkkV4S+i8G44OfpoDOe4HH7XR5RB/dlovgvpNezSQWrwjSd+TYKBg2Buo16xj5fCXWzJF
PSz9z9TVeXs7Bp6W7RxmjhZcZcBppsffgWQ3UXiUXDPFIJJFP3bsymcT24yxxYPaNceqPtb0mHfa
YunklTiH8dN/902TKVfECdtfrhY0ncqgthIPKPU+DhKSkbzbxR4IbiBi+PEn/NEDxQb5K5HiqyXU
5geIHUKfvlbjtfocxTYw8nfqOzB9JDlo6imzzIyJcITiKAMw6iWtWbAbUrTNvPmgzf4IAMFNjXyr
fANtPY0LZvkORr+/CGFWtPJl0wkPeX51joYQWR3kKIBtzlTypFaZRyN8BeYbIi+06Ei+my3HJzBY
qLX5W6fYvWAu1mVmiUvedl7kJXn+IcvoUXwlZO4gFhCufghDb8J3xxCbcVbg7hSzqpvi8Kkhw+n5
DutqShkNRB0PHNNHVneXmVef3ZFytaua4WWC6Xw3HDbY22WO2CnQzIyEddWPS59QwZHyfaOrNQLY
eWrikeIcVGfA0SSXV84hxEdFe4b1Y49ZaECV50X0UXt/7rz4B0Vz4FmtAJlUSeRDZ1DrXAiZZ6bT
QlcR/GGc58StgbyYBWf8CGXob8Rc993FcJRMIG8drErzSLR3siU37CsAstptMvxnNcXt0L8RRZCW
lH1tu6IAgoT5c91NmVPExjD8k6bmoIW6yfwB7NSLgDQoY7k/5pIH/dpUX5L594ek85yUlj+qlNjB
Rfg4jCrDD9nHmluH60dxgu2cw+OpZOXoogtvAiieJj0CLD2UXXywMJ9QdEhZvqQgDAv35JpaShze
CdVbkHECyNzTCSEFu9F75rdgncmwcECIHfBadPiUTstRh0ABxpq4SQtJo0+nFIdboJYi8DHuuMWw
PksIxR0OK5OZWrWiIv3CWsswpJOBfbnLvOQfpVK1xJ+MuOyKUzgKKSIvt+CVCFvvSv4qgR2aI6Zs
QB745YkQ4HFDb9teUwTNElaidgEuU3oaGl3ekfn7LwSJKWbOSw0oYn73d+xBc3+BdlNPrdZy0DGw
yaJvXs/aohU9ZURK+A89kRYY64KqtfuMwX7JMnVpi3VWSrlMiakefkodSY4OA/w8io8NFFlALOkD
ZGpkYwqPpKNeR4LuTYWwUBrx1hk63PVYFC24Jud+yfKYyXttxc2swFWzXoAs27YE5l9f/fZmyCoo
lx5pqDk4Hyr0CvSxNs90lXeSh9XfiFlV6MEkkif66t2lYgcGTIMCE34vTlYFbs61kOXtGc8lXPNU
ynKRHrLDdFXyfdMY4U7j5nbC33zDgI5oOASZ/3xQgKHzy5yCh9/0nHEVKyeD8W3jOqP1OqYxmABF
BSE+c791p5QqUHcwEhb8DviFpNaShN8Mlja3xrPCJX8NlgQxBsdqyW+8fxb7GpguB2n71Z8gWHx5
dYjxIeGrxofZ2p0+uHCTvXreRj3tpXJw74ReQjU3n2lgovFr2xDmdno9/FWOGYLE5IrxXStF54yj
2j/hO2PArWtrUMAEbr3uDzRX4rKMUH6eFwy87F+qEOvwS7wLY38nAPoPhEvXrVxFMVjwKS98RlEj
OIpxDJTk/Cy6Yh6vXTVjkvS/45s2hUxjA+2YlT0hQaSNJ2jlySq3Gi88RuahvLl65+0o8dOydGvh
pSTBRU2ZOBhtRN7e4AQeXXPXlXsH4eQ3l6oAzCyMUUV4liJhYxRiVhBZpTIg5egjf84JyMAFFqYw
pJ+5MTFGMk1Lz+C39SzRCW7JJ2rea3aWrWqNMfEkMjlFlQPq0eUiuPvWJgIrJjgXDdgrxgHukJDU
y83MFSSe+nNMXBArjkIzvFLc7n1O0K2IPf5tmgdR3+AApvoCMQXt//p8ZazaWWDBYJElOWY0zH3t
fohxj7iqVVmtJBgFiF7oLk4Ik9moaOFZ2hRTlU2iTxQGpR63U/3vEMlyMqOCDDN/V3upFR1vcha9
g+R1QcpZX2CoTc5anIuLPcix6YKpLRBIbWwE0uBcuZvS2VZ8f3Q2ygKvzZBnQ/oVDiLa7shq5euX
4OuLNAJ5Xy9nT76/lsV/zqjBEWjnuhwr5zALU/mfaP0aGZuThK8D/hWICrP7hv8KxJ9XTrwG0fpa
35U2ief8eGRggdaqy4Ri7zr9HT6qGxdYiTxisiqwDrjkrWP3ZJPoGxnLcvTMhcHTYQ1/3UT7jRqp
/YM1d+CC+9Dao14NKES3cmaLiEGEexcDJMgi4D7jBrMJ/REU9GZwe1za/uXFLLojlEFlKoWeMXbg
Qknxb1NOiustznZGy0YUTTunu46s+FIaoYp4BIgTren6HLgbXAs6WkEXmAeYx1T52nIPiG3PCKHD
SKY/2hIuquAsmg6q85+9bryXR+yprxIkUKhku3Q261d8RgaKvVb68Co0G7JBRSTh0mDB0facgnDr
betyf6UEMALfd1cYB2I0+kWC7Ab5+r8bW5PeSVwSU9zawLRT+6i9MTxCp0eU0Mu9fPJtLIPejOQx
UFunRCRagFjNQZ8hpaFYpcGa5SIvdleCiYMXVZiTDHcEHqqFDWzF4zud/xJTY3oSm9Jz62/k5jCK
adRg1XG6XMwCA1mq+JFFZF3ds/hNgJfC616vu2n9FEfpnPs05BbwO94sLyx4V7XA3bOFXs7FGmS0
MC93wgjZDz8/ieMIKRRiKWFSTqbeEAwGXZUM8Knxddh0EPb6YKzuixnRNxOh2r82Wu42qCzfv8yI
ci3VGTIbnPm5HFjtksZ99Ycp8SzX3RuBoLdEzJWZS6B640G60842/6qI8FDwEcsKIBH43yJRd+1e
BEzYwa0JOyDgDK3kJ1CEZEzoxQzFqhQ6wlMSqGykK4clUdrn/chnUu06tEDUWor8kiCZgOgbo1Sl
/6/54qG/Bub+Qjm3DSYxWivggTyJUM51RzaawJN9JFw6recBw9N1VwsIACXs6fiBN8eT6gZJhQ2q
8pOMpJ0x2LOSuD8JeTSegN/e1one8hy9EUpzyHHema9Nhl6xBX5jFeEY08zSqy5lU+0m2y/xfDDq
5G1NB5nTVlmpWVo8m9G3tEPCZYna+Avb1UaUM4FcvbLRuE5QtNw7AID+iD2U5tDTABfWNN8waZIg
Soevbs1hCyqxrx+vFHlX4+mk5TZ2/WI0Ex0ml8BOXFon7eN+rCH2dYQHfNbBb19IExKGFznmb9+J
AW5rdwXM7KQlG4dmSnI1Onn420bmRQtm2Rhj/n7HVAxtzGDyv1JAIpFk275J/hlCTyr/GCriZvxn
hYZIo115sEzKioLsNm7fi87xJtMEwOk+LC5bETMQry57jbPBI8qZyLpapsTg6zkt7ewGNqqlswxM
PVdKBmupbiPY7goLo9VwegOQHSvGVtKDu+eE/x0FSnGnqsym7L02zljOmvMD1p1DHZLVZBGA5YxS
2bDs4sdc3ZWYIrCSOZY+GPnd6kP27PSlrxCgvOakppPyP7OZPudSu/18Ab5jeRwC8FrGPI1926NZ
4l79LgN8DuVq7K+u+STfxjiS9bWIWKNob77iHokHVvj6Z1rEF5chFrmnWxQ5s7XnX6euwNS5L5vj
eAlLHV5lQVe46oBlp7sn4sCuan3bZ6wW4E5M44DW6wtUkC0OnSthn7EO9PtKyX4buOcm6W+GdKcZ
O8Q+3Rsx5opNY+teoBFel4oZXobjZdZiYu2SxctBwGGcOy0kkVxvfMgxcmLNx4j8fD7LGwPJiayc
r6Z+TzN1RS9ja4wg4bWpANc1yG2ZM1tUQZMrZ2U6JbQ+dRHjksKFHNeSbLeHkCH6xYQI45jezPLf
KwVinieQcUihdgjDj/UIasysVedo0vr+/H/bkEDj72EIyezZNnBF2V5NY61b39yefDKL1XUkmisJ
ohUxOk0r+Gn/p11zRz0dgbGu9m0cbeA9J+PjsIaGs0PPuz7HdN0BxxBUXQncX+5EqRDmtO7BghME
KCZIZQXwDffUwDJKULRNbIRVq101+b2b6Z7ntN4TfW6lHyCULO0flR5C81w0pHEExnAVNf+JiNFP
rM8RiXwujKINzclQmueldnON8P/JHJSXyyGkYnsO20Ua3ZgNSYxymrRmF2DTSsERoOkRjQOIhdOB
DJ2a8zbhsApjskcLnsx7mfzt+/IoDcAxT9x7EdC9QLwOVD7C5SQA61jQujUUbEplyqRDZmT4wrxG
lLJXIvoZArBS7PNSIIZtX62bEnF2yECQku844Zzx0Pizr4xLSV270pMA1w51XII27t4TStMV2TSJ
kwTK/5adDhfxUKA8RPDe4nQZSrQcKeHZdWJamieYXYxj5YoINbVtG3IctjxduaEz02xtYK2GRXU5
Z3poKRT3tK15cRdIvedVxI+d04LgtHLGDgWa6zma06M6+J3o7Ifrd1BOwNlqkFuZojnRTh5g8CGk
06L1amPwen3wmInCqzC+7TDldxSgKe7K4ZeWtpYUAsyAX+3N5dgG5YOyRBFiT+uzNTpmQGLhn+bP
7UrJIfNj2aZaVI9yWyXuzdYhzCOMBuMUPC9kIO4GQTEcbZ4agxrCKjWLvtAZ3XyCgh/NF1uL/Rb8
WkeE33lJmXgUAgJYx1Bpqozl2/2dL2lhtTZVFeBuXOrlHp49eYhnAmu2Jy0TNNxmbKYR6sJHaZ7U
FVruM1jBQy3ulO6OAgaa50hjWrG/BLUhELK+MopU8wVdbeEZAh+9iHFmHIDZVU9k3jr/Fbrbr81p
GsC88xPlsEuCToCLYRIBi9YvFiC5lpgWfHjhYOrbh7ay3KPrGrxusKZx0q6sUAhOKkaq0TOIt7Zc
Ofj+NSB1AUzdBSncSWbo53BQ0bnhXtg0WYVK7TKbweS5h1HIZObrpt+jq3+Y7tRLA/1xc5PfAmDo
x/BMDwdL+szX7ZVEKXE6hBgnXIvgioW0lcBHIAl3bEaKoRJMiycV6+oPYR1/qD636BU17+HDVrPu
gPBH8bmXPdloWiOaKjeonMey5lrGnZMpQUFNg0T0zdA8mZ0r+QJoRST0Ck+KyRErc5Ek7hMKLSuX
bFgiQ4msHwjZ+F5YwG6VhzxBBKqMsIoUQB+SZQR7pPxXM3jPAfV87QizERVbyrx6vuqoyncqgwgj
ak6AZuf9/6O0n7OcIMArmnXFbSw1im3EvMVmf2lCYlj52ZnloIMRWtB9L7BjqbuvjXb+bq5vubmM
08ypZf8ldSwsuGod9tMEKJ2pbM1cgiCntC/MPrQsUhpZEMb9+myiQN5JL0zrOzW2EaDRYVFjsBvG
CjCpM16d5x9jG/w0cX5//hJq0RlITacHKyfLJxJS3U3tcHHW4TvUzDnJF7s+jdqQapIJDRSBM2/z
yZKdqCwd6o+0enPVmm4R1hvdC0CyKBVEs50jI7jgS5/GenlsHIkZhdwlF4dLTPdw4lvNxZIqcHHG
OPByBTwQlXIiOOf1B34b3xEhQh0e2YJauyPz3AwltH036wcv7bAFNoTKOwYvkPb5p8bLOKQ4phoR
Xf19oxALfno9kprK2dE52mRpKnyPjgcs715mZpB/Z4VAvTqFVN0BrGIMWI6JQfbfNPS0tX9gvJaJ
aUW/eBAuMU7vV9uFBI3KzkzBbg4iIq0wSbQVXRy+coroZDfBziHqyTkhHNjNmXLk1E9/LW6QUxg3
7unbTbDgR5W7tcajaKpPs1RS197CtHiV0NvJCgCWk1YZuILy8EVV+Gx/HQpTGSeI6mKfk9i4TU/o
2aKMNVIYyI1UbDjJnpWwp88sf9IjthsokOfxpQNFqpqG0kIEQn1mSUfV0vh4WPagvE6/UVE3XV9J
5lfiwr61jwMqsT70igwTwK8c1zUV9+AOvBam/TIYKMy8LmzyJYlFh9Fj5Y0Z05vqJK271QttXw45
QEQ89JYdbSjZ3mbL836YbTtqdUvBDPLgpPMui3twR8sc1x6i74EEWpPeLKXchtGv65ZBkHSnUdt1
1aWjT+XWqVs1NKcw0zXMW8XFpLfMdw1mfffrvNfZT7JueOFAyzPOaNP91v2YWdSRQnjF7a0wdPxA
L20zUi/Pe8qWvMyHT129jw1H26fZ8Kf6/hx9mc+iLuJspjHVfPk7/0mDjJFkv24ITm5vT/45psgL
gSloXbCvV0Y/iTHcgXDvwQP1W+QucJb/Oo8bcD/GpZxkZTUHP2X+A18XMtVE58F/TPctZEHFO2yE
DFayo4HP+Aalfffh5diyaDfF256sVckPEo0+ucmoRQsVkrS6veag2xrrJ4GUDWb9fnpaRLeIKJkL
FP7vJxGM59i4o7KNgsbgLC7kIgqy6fw/0dtoD0lcOmw0Lz394V2scypZVKdFiuzc2OTgQEA5Da/n
n4Yoa2WFtif5dZo+3vY63BQJemWvFPW5fEQMAZwSJiB+A5d7I47IOC2HFfknFYqIL+mxCQF9Nwmf
P0kW+2ZQ7LlbRn6SVBqW53pC7UIoV+UBD5q8iI/AmaRIdRwYNHnE17fei+4RGzlAFCL04Fb9zyI7
ckENnfsoviMy/KkkqxQb7ZEZPpfzRWIUw+7LqE/4nmsFNBXM26EwkZzApw86+NZkasggFZJ7Kb65
z30lJ4SUp9THIageWCZN2dfxiwJKe6D5chkt918gjXRsO53fxAHFROXkxbJQ2IOus5iIck4ddgiz
H3OpkGX92InxWsyWgfj6x7SVyNHZj1Kz9+DKBSPJkz9rwHXN2KN1noY/NGQ4LXD72Ln+fgqJ/OaC
CTNZ/I4JQuq0Z8HJ1bAZBeZwEr+TvLx17uu8/xcbX8oIguoqaPVI5zYUCUesO1kLstf/3Sjf8lgt
LwuawcGrBFEzr6lFYCnZ0U952rg9MUaF6Bc3+6qqh+ZKGrrM+013pZn+do5hovNBpy13cgdhY+2T
VYmqQjIQQ8XFuWY8Wvui9ESfu5FGKL7LddFu+frAYEzqWI9c7qDbwLUcmwGx7shQmwTy3RgPY+kH
4GRTC+W0B4RyD2L9qP+70GyKNnzQXlKFC4zFniSyI8FT8fGEverenuTmNWaP6y7WRLkz/BVWmnF6
8xuMh9Ws4NMcThvSRtxMpFf/rHoZo+lqfteuWyothXL2tCC0NjF5x4iWy/ljJHCJQRtn+dF1g0Nq
azdkSdckqiRusPIvhCaipuFoP0pvpUshdjPq7pGIKxulkdHV8IFu6VgeBVerPHrEYwx/fIafuYnC
oDrFtXxf5naKYkgz8qjkELVJB1G9uFeEHMDLWKkA4X5JodjvQaVymeUvtFpe38CTLZQyel1Am8NJ
qz6+uAl5GFrSXmRoCzGoI3YtZgdJjMXyu6fqgmJXGekia2e/jNgPGSs/rD4xItMnqoYhZ7mIlXtW
eZnBx/ehNoYIHdvCKGIpyetCt8F2BJE+g/5dVOWDBO4O5CtmXSDHvyBmRPv8ZahiTfWm4E11zKi+
RWrxJU3lzUY8uMM/XIHDG/lPeMexOoZCfQLgmAGWA6ArundhG73Mgjw8B/L0py1YAy983HUYawst
5zILzoJ7jVsRKkKB+sO1bsiSxNOZjU87c5y/IzN49aT8OXaYlPk9sAg0PFf5xHRPA5gP3zLz9uZv
Uf0kSj8dCx4MgLOekT+Mafkoa9KVylDvQUYHfnVPFmlv51A/L0Quz8ck6cLCPaZhiRptPACsgPij
yh4HL9ti1Bq/b+kzabNi69s6Rci6GPdpPKZAmaViZfFjka+798pbLjTzeD9mh8s9h77+G9aYAZ4T
8yrZQlrK6VywwWbNdYwXusEkAmM63aixbgW6UmJJQskuwQ5Co5c4O0cNhZdojDZ9xarV04734Op0
F24ETnWmfygIFcxycmPARuPFHMVUuhINMPSSiIIVGwvmc3Ltntlh7WVSIbpbjuFqc0J027VFwebW
+sapCwN21y4v3m4vQei5YKRSGa9wEuPAJqiiHDichiiu4aq7ac3a4bpkf9GQhlFT2PDA2FBtirur
tRqisEZY/y4ksHZx7VhwPj8fIVpT40jJ0wi0eEKsotamPvm/yKaFnm15vAEmiTVcFFnQ5RRLiS7S
dFxHxHF1ClzRc3ti8q8ZY/Oy3xK25guKU1BRPgkYFUyEsuQTbapaZkqcR6QqBeoJ2qMnXYJMdNzj
/dmGr1PaFXqYtlx70OfZWxZJE3CRxsPxDuatTguLaOvwZ+uP535+OqieerlPKm/Gd5mjeV8/WVsk
cBxAhEx02BTAzdH68o7yZXA0QRxHbh0/ZeQIpVD0LAmEgHkhIrfuT3YFdF5FEri4Ey9ObYcr/ysd
N8/yt9VYtbtbIPV/dqCI6RxOTTf88f4ppHdQTkTtSEL9ZzMiHWJ3mD4fo4UvoBAGgPEq/U6eBw8h
PW+xypsT0FjB/Gh4eWZioZpVhFV1MRbhsYRQ7RdeZkI/KGNTdKglZBD50IFNgc1dfFNdlVjQlimw
hCmF3Vc+tYxAMx3853qCKcopGRrcA2IyvmaPMdzdGTPJWqcKmucKUGwHgWKdaa3xqbHJwV7fDaL9
sB8lwQWbQRqmRgQ3ng6Yo8kZTxDPROBL+lUgnB2CuZGXf44ahJ8qQ/h8SQKtI0doylaTLyv1pSFx
QoXv+DR7H4VIHEKfR80yLY0wlGxn3mcsO4+PHg/AThB/eVsiWc/zam5ClMZJiQjDO42eKt9AOyx0
I15nL5Oa9/VkvK8ABHX0/jpoyKT6Y1SOGmkEl7APU/XhWaMX1eANHfkYA6kLMAH5RbG3aOt+9T+U
bD9J6pYMZcryi1VjRSfzyFucrkn19TiXkelxr3ZrmDz1RP+JWuCVLq7SyY4d/xK3D/MRa5MrihNt
kCS0lZvm8oIGXc/FRI0/K2nwUp9tQ12gJdnw1roqjdn19eDnjiQDfyKdhVLTyJxtsVkxkA61gJ7U
XC2EDpYMh3ZJ/BujAA2EmmfApRsQSbX8fWid33HhslT30qdSw/45Hfn1PXAXZZxZGB+6112aKmas
uEEplacjLKXj6xbNrlHjFzu2KPZE4jRzFBiuDVJ6prcizWd1FI+7MvmcoTxn2X3pLjGW6urse4en
g8YFueMBVLxHi0BwXA1iWKGL2plOYrZ5r9hMQCuz577LReXE+XwCcynioCQyGBZ2XlIi3eLrmRdw
Q7x9Fbw4+H19bH9qdZJAYf3FV5GAdURG78a42p5nCMNr7f+q7q0k+y3H4gVdDEG6vXzU26Db/AOl
9JEOAVaBW87qxnzwNXnv5RzvJT91I2Sn0s+T7iboDGK0NdnHAhK0FHER0iopHdjLWYELDpfyHRbI
IYALWvfoLpDfTykkdxiAeOt4RqgzK7rG1VU2zUoM8r3ZMs9Qg00HEO3sh2QH0raCG2FU4RQywTKB
Gjj/QFLmFwVGVKfuuum0+C+dz+U/dY/aovFu/Vko1lukjtueW4iz4RxvZ1mYw2pQjwBxJyNuvk8b
K/YAxnF3UBT6P+42xW/ppUn7sqfE6MYMaQ+whBOORMGwO6KSSRenm8c6jR+I9hIe3Ksz9G6ncFSc
hweCpOaJWLjQvvGK+9/MtCAe8Ii5m7nvWc3Lzgxc14pd3UpzT0AV9uy5JDor/mKaL4jC/+EU97js
SX08jt4GpPeMu481qgdWKIl8OGsKZHU2Dq5s3RTkBTMHmN/Bcao6Pfm4q8n3goV2QIbrHjxhqwlm
scxsm8t2PHNikQnv1M81w/i4aAHDCbFw8lURd73sX/wnWb3fshc+y2b05wuSFgCCFwEv2mojXfCe
lOyOczmLaycOxz1xJhFxdlUTN25uo2Ex1QPJF8bxPswL8nZ7BDm93FBEpDH2pfiQSf/chrWWTSmz
TSbA6Spi42xpHygoiGzPOqAWaJVzDT38Tg1FtUMnImU8nwQidejBkZ2huTzv6VfCuh+4G3yLkwmg
DTSzgdw03lF4OrxluELV+/u/AjQikqU9FOpq2elxXY7ix6bmC8mgVGBcinLSzQaxKgHFtxQ+1ett
dri6ElFi+M2YZTPWGywBZQZsyd+arWH1oByVSPglZ/JoW2fpiqHPOjzTfudrOwEdAd4bjzQAr22k
Pg33MTpy9pjJtJr6AwUIpA1UYYwK+u6yxjkGeWblRc0csu1aPziXWJdLxZq+85USogEX6n+pXMIQ
ur3BZ7ByPaPrW0cBbbF3ObUDwevXv4FnRuQslBg3Fxe/Z6FQaoX2PQTFndR1y9VuwAIlhDhhSl8O
1aHKoJsRBJLn/OYe+HfW3DEtpHh7y6M1Xf+0pYlHCojeh4K66+DBAXZUrLfLOueCW5QZC6jx93Uw
o8TGjxLC6O0bBixMbwhyk6CSS4u3IuB0ZhykyUuN3KB41dLD1SrqRC5BES+CEoGvC0Cz7AHPawvN
dqf9N0VQeTDJapv2wtQZ7fkNstKNgHbH0/UkdBlmUjrvVYG/saHX35TBPnv7/oAvMuZP949XMNI2
XmGF3n0Ygop8XEVcO7HPNtB268Ct88CR4bsCc2CoY0LSFn4EUo5HXNmO+HFAW0xU802HInz500kH
svQBsuz/N1GbO/uNIyNAUp5zpp4ULlp3OMr9UV0ZIoA6Hs7lxVD2fnHgtIx+u5dVZYtJhlSlRg+w
S9QA8qLqgvBjN0cLhAfkbpMEGrq0xlq3nRYbpObFl498ESAdyuVS034UgmgO4JUSs1JplsuzEDaB
rItJmTcp7G9E1UL/FUu9cizL3hdkQY9TQPcaJHJFvJA3PVW5iHFaZU9hxte15W1vZcxTzw3eNttt
D2i9TohcFhk19bOOso6htx9Lc4O5OMChfjxuVgerIUuMsIvcfxWLlH+LgDGzQThcXkXnYB9wvSUi
x99f+hyO7FjqP58kCbtB4oeJwMFPvnOIQVOMSmIvy5ZRLt6WX2i6RECN9+fbMF+KRuU0Npu9LQMO
ckGSqx6yvfJRGWgzeO/Um+BRq60RwQH7FTc1gcXKlYVqUBUPaXtLO6SsubQXGOSMDwV0KgQviy6G
K4N4w/HF0pNS5AbFbRvK4oDyOSC3Mmqysgw5VUrvt579b9K4lVxNagOygHE8ElC7KSglhjdxuBR0
APGWQmSxXUpbU/5x8sto+NStWeZ9abGSxaJIO7L4bFi8KK1YfvjLyZMfRGgKasS++I7IxHgAKo6j
bWUbt0pHkuaGI+3r2sy88f1GAb2UINwKdePwJS7xx/B9iN60zOSwkT6QSZFukaD1/xnhDkOcSBus
XZFEhl/wmAg7Nt6TQQoeqmb760fYOlkFXInIx0GnZ6v5s/uXI6c8YmzXFY5waM3G4jalm2w06b/c
uxM0cHSRaKauftGm1dfOmUqYHa9OWrQ8zX5T3D0a0kqXZwpxiAxqR0vwcYZxxY7Bf3WPH6siMdIN
S3C1KnwM2nOUZibquKCceYBYbKRTeNqEpeGoao1V4l6v5YGqkLmZhlGOCyIZb0TTqeLrNHsYf70N
B4hAX/3AFcQqCaNZKfYpiZtZ+BKCyNJ1sP+s8n4nM0wqnIpi4mFwa7bCLAwpfetUssEsdwCFAnze
c5cab+cWmTZnZBvyC9T1hYCmgoHEUs4nNquxNf8AFLTQLcktsijJWHOKdS1rUFEr2zARQJE2nfPF
1romBAL1QisGJqxH9EY5Affv7s9ojkPPTPexJZ/MTDtQ72uQU302pqfn16OM9byDgnISMQsQ3mO6
K/0CwsV9u9uQQ6JhMGjN2/jeo/McUGXYZQigkEppAH1TxKQPkhzwX+O79prlFpXO7eQ0JxK/MUfk
RTspMII57l+ct+5ktQKOZ0ptttqn/ohUoEGgEda2BasycRmOtkZ0+KQrLCs+c2j2BxtYtufpiphP
GCyj/owBzxq3l6nkJS2M1trDZhQwBheG8y17QwwUQAW6watSNcgDWNEb4yqYUn2mx2k7PFad6BrQ
kJbYZMKSff6wG/T7+1U4VQj+Qv+ILFAMvLbQ1qFlrbYGLcy6BLhC1p/9dXfGKwhx8UMak7V2EZyC
1nXKKhAx/odHWKjZoKLgP6JQxglYMIbpzOr+lvYFx1E+Gy7rmdAQcUI6BhdBrguBU988ZIJfZAEp
njLNF/L1983UhF1a1UiBF3bxSHnjFMcauaQ5HSb7OdBx6xMfIa6TZQ+Y86u6me9CmMr0xxuJwQYd
n0MneNboN9N/2Gev5Joc1d8ZQ1Glkq/ZwhkeaXMNqbnuK/SSFP9F4nbOki85e4PlsuXfbqWH0X+N
1sAbFz5bGZs6MsQsNbibBohGnQ73UrKk2Xoigis2FTxHpha8nA52S0rXGrsyLRAHX/u1XpiwRwj4
tPTj4rsmlIGN11V+vcEYhOUvEs9kNnccXPHZkARDgHMytD/zYN1eDx3/GDGTTsIiWR+ZVGLJP+iU
InyXu8jWop/Bs7RPqOu32XWvfR1PeGfq88MDtbjg4bKlgtWCNj/P0HNsHeWlWl7QFrjSiS0ZA0w3
VgILDeq1lIrS88P3p+Yp8x2rhx/QQr8uxPOONROoMOKOmly1w75+lyUSDb1gtCZz3DbBvgdz4iNQ
TmWUex5x3Uol7fU3NCTtKCb2pkGxqB0iY1cU1RNk2oNZmKI4e+OIUe5hdL8IuFGey9AL7b8zzjyF
OPFSwJJ6q+w+KtK+c1zEphnHpjAskOTy78jJur8byKDfl6v8FA/zw0A9WV0jI/v4iiw4uJYfzQRo
1I9gIEgTKv76SoVXW1bEfdlXrO+5ORLMgmriEk5sSv7Q7FRwrWj+HLfDGWIlbhNtYTXFSPUdcZFy
c95xnoa7W3sBKnGh75qOfQFlhNJYPkVwqZWCu5uPgw+aFkiL/JHxQ5DUvpdEONBsNA+kUtm0PDP7
nthoC51pqkBbkHPnqADZTZzZpFUp+hYfluMUaN2p2FwanATyIeql8TPK6WMLD/IvEf2Cmh54rQQR
1spRHy7b4+DPcThON/eyJIiBmWvbgwiKjRH3h6R27VRCNqFumWgNkbcvi2oJ99xgXhyAq5CvxQrF
tQ6P9bObY6BVhbXSEhEoEhEE7avkFaDO8/XgG8MzIY+7PYnemJfH+r7qDwsBfxbpjXBVoDooDRTc
Y2iz+nSQ1B/X9h1xocb466ObAiiY+QvkqHSIVt/dsxagsh7eET09KQALr1lc7go45UGzMkiipvkc
ZIHKsztH35Y1/j3X1H4MYPyZKVcDpQ0o8PgCNAVqzcHCzuJwlSDLb16vdi/n/GbI3LirQ5vAby6G
CdnDlGYC+PlkMFwp6XmKpNG+3wFzWA+ZI77di4Gxog0VpgyUi3WTw1Ltydmvifd0bClzEZ+vinOd
B1McjNYOH/6lF/Bw/Xx7KSyH306KHvoQcDmybt/q8QNQa959oq54XViOTK0GDxr2OGTDmAYNB1lp
9DQFU5SXu4wKKvFZ/lK5/f5RrkibWPJ/9faaAVx+x/kwM6XBNfImwBCsgZzvVVo04ybHH5MNzT1k
z0ryLycujhtO0sOQ330BlPR9duUbM4ZtvBO9h7vfNhEzQ52jU0p24LyKfGx0lIsK8UhCO5PcuR8F
L1U0gNlVDzUKYrJ4P+FFhtK+WE4tk6OGTEz5FQil39O1Log+tvtj+5ZR29vf72unG6mBiGyQyINL
tdEio6qierHTFui+KiNmCljE7neXUHFHRD5Wqt0H4vEp2LRfAm1RgvBMOplPNoax2EO9N7byVjbA
ocjUjT3GeXDSRxIqFo493XHASEmEZJn37LyKz/thYgiHPRhb3kcIorp+xzi517yQJt9FlcXR++1a
LOY7s8l0W7Ktv7B9IpYhQljNSDMFIKY0E1XmgRCA51M5vbue51w+ET7+i3R8uxgfV+Wj9a+fWooH
W1QHfVpCjdYMQlOoGW1StAx4aDf+tg9PyR3jHtoWhnN7FRhmlBbotpySzwnlsFdCvAyHIyfyWmup
SMoGLN9Npj8BSrSG2T/McDxtxbHwwTiawu9hykyhUTQrOK4XCxksGVhh1JFLS0Frnjp31icFQBn8
aGJC5sMcrtn3whPI5jCc8H251Eid3WEJXuqp53HSMqkJdzaTg/npbsPdVFkCV46ALpo52pxnJNLZ
A89q0CDZLzFVARGqppXIKx5JsCPG5IEqushKjtYVPY7Z0YFF0GQ9n3b7NRNcxPb3OTSKEoLCkUNb
1K1rd4rPDRQMJbvwjInoM8KIvzzZFenIr1YkuiB6d0Gw3V5TjPgiP9/yVRLPCFtl5VxyMoPvZCRy
I5hWXGd25mCWU6bLYEeJL4It8n2m36x78UYMq6ef5hNizW9spw+IIB905HZMV2zI6Rat74NTqQlg
f86mr9Ikhq2k5NdnwS0zn8d58IRAUXZoJF/iOy8ZNm4m9lHtcvklwndSYgByH0lHa6wpqa+YMDFI
XzRHtJdAqfK9d/nBJKB896BFt/y4dKX9YYa1pkQeiqYZrX1PY6mQlN+wpT6FhTNf2dNc+vCcCWac
dOQ1zLUkqn5xQKniiRYoLOYQ0jWwQecziM7tDjd25J8Lazqcd5dT1J29RMNgoQnqWuErkpzj5N3s
on/iJ+FQoG/GcJm9l29PionJIrgyMgQE4JohizM//h7TP2GQ7IGEISwVcjvlDXqFrbxeZ7aFG4nz
s0pYO6s5BYDU13gXB3urSD04ntiYtroxG+O41wwojYts3Ui17cErlrNAMgnbBxFziSpHdTReNAFC
H6cIXuAB48EwWv7ddr0U+hTDSGqvQu3iQn2BIgMMcik7MVyVZodfWRP2kFsgc+thEiBKsGI2HiXL
6iO/wY1q2hyse3d97RcdPFi/hDlIhsYZGguCw4WdTZDU/yuKXOFFjXKiAWUE+B2tonJdfTwSVM9F
d7C5WlLE0LxqcuTHJsRz/wltd6iPmFUU6Y+DKIhPwzpaVuoWAbozI7ng3VzDnnHtamOA+VuFi0kC
WP5VCLQa0PwlxlVeObzNjvbw3mu/+/o6qjYqrxYDG/zeneyYtfjnOa5P3T90W0J0Xoh89F1UMk5S
+nA1r/MelcaAwBEbOJ5/qIOcXuWynCu/amXtxECiAGXZcxy9l4elQZv4jlHjxWuUoXRstXM68hc4
IEjW43dhmcxPiDt8i1uEiK/t88qBAh34xm8KYSZNzCIbevHuDwhRRMUJ7GlQoS1U7msHc2jb6X0/
9/RpU3WwEiz7pFM2O/WVMBLKw+fZcb0uXqWgz/NinOnKTlEtp1nSlmud8DI2n3Gl8ygobr2MJc6r
7eA4E64ld5rU3E7xFuN0Rb6RoZO8MQ0qnzkCHFbQ0Wds7riKWrba9ijI3Z+T2McfTDcsRJsA4EUn
WKzs2nwR3/oAM9oBizhfXr7DbQBp9Wm7h/iv6oJz5vg2P4+105y27oG0Ennfb8Al4KGFeT3yMcyT
f+DvSv46qm6tB7/lWTLerqrApBvMCXOuB/v97hGFdbj2SVHe0Vr9pRzbgIQQGasV/cJ5KA+hQHru
Qo1Y0xvC139wwGTRCDPtq/JCItllwJwTuAdqzC0rkXHb6Od3GTW8fsKwTPmhmKuWvuuymO5emab7
thbO2Iuxqml9n9Hnr1yxjZqevTRpxLCWqy1bH0stIqj6tgMLx0OlMnntOWmoQ7CAOmA2YlVSF5T6
KzZLQmyGkE+iAhMqIK86p6yxuh579j50ZpxDg5Jrn5/DiC3MOXzjtaFgDIpy0GedKrEQiEb3L63d
sxLYhbJi47JL8eLrlcHASyPW3OmIpBVGD7JGt9hSxQ4CkMYjP93AS82/mFRueYh5XVfKj09Nv4q2
tETJ7LVnBvGMaCChzlWasrjHLXbEBcaJoFTmeEKR02Fgs8qatiGzJVOCn5aT04ts1zBpa4T6kL4s
Qt9AZP85O7zDl9F9SuniCiNgGy4SItJ8acaMwZbl3sHpALI9JBRyJeFS5971fMawXEVUczV5O08N
EoFr6QsFid86jeqreHuGRmzQQUdYdMWjxbn8Lb/hLHeoX9eGvdtbVHiW/8+J1bhlWp/2aFYsYgjz
L+ycrJiEFZySju0EbCxgJipjl8D275uxpQVN2BPdKvqySAZBpbzq8ohz4nwk1GyCeedZM68xyhLS
Ir/iTcgr3OZpiLQWDQGzzxFqTIO7/wsaZ9HOt3iWEq9wk+SBbpoVLsIKIP4OJoVkLXcMOY9EaxtO
ME+n7Ce3Yq4AKpSlpLlUtWyZOJQNnZmG0hQ4NqeLXY3edv1OaYLUvW+Sotj6ReeQrG45EE4wx5oH
U3QVpUsjoG08FraOefXjkBE6PcZq0ef1htGwG3S1x40fyFZwrZULpYuIEcLC7rs0MtSfCziPfWrr
WIMXmSDNNC58vSPcsmJ0OItfaeiwbk7eq57yZ9B5v5GineI5dcXDNyALScTVgoaUiSIquHDQ0Hwx
ZY0QpWkU8wLVfoE88WJ/H1d5RT3wQYEDbkoQ8gx/thhQnWTF8vNh/pWQ+VwHGolwmd5X83gwpAcV
x+lLo98f+tn30SPgoNLGM+VUhQkFSyYwg0p20lrT+Z4G0q/k3YW7F8JQkKmip6dTA7M2FJaQh2qW
69I9mN36Xm8NeBA7AdxPvAujAyoAcocYJiAtydTj87tvniSX42frD7wK8biBkhhtEn2l1kgMCZvO
SdGvOjYad0Z3ePDl4odSawAVnV0037YXe8jqYYHqrNfzdq1iegWiU+LFu1kRML+i40xMkcno0ToA
cdQRLjOLHt+fkIo9fbQdNljn27ZiHe1SPmOSa/GBNLK+CAjltb77OZwwBZ5q6gY3coBIWG2FqDPx
rir9Rt5VX2aQSqLKm6Wlck23afKTLPqj132ShXiIwFZZx+msJSyuCm3MsloNlRS1BXaZ/UpZilEW
ysOt5z+o0xFIhU5obIGGh8AgxUzX7Jsd9SgzFly0CPAJ0l3vADXRRiYSP8JxoCUgnSVb62clWPFk
jp4GQil3Z1N5Jsug92XuKNCYrqnRWSKY0JFdQTT2Mimd5HUGGvFtQLirXW2oiDQw2ClqUj8iRPIS
DeIzl5042F2vixyHmh4eTkoUUpVEIgoGLjqvzIEepZozdg+5u18J4ybt6Q/c+j1OZhCtsgE4EfXp
IOS/N1QqQmFFH++BbhcRVoEC5ZeVMLGoI/n4SunmYHGSwUIMf1qDaGIbelVygQm3Q0+7Z0974zo+
oCiuIXYU+75ON4aIoF6AisdQNIK5Rh/F/PtTcFwqZi9Ewb4ltjP9UmfZi8Flr/pno2z9Xx/cMSX9
nOTOC7ZnkIpBayFadR2uFu643ZQF1FJzkKIVRMRb2yt4kmACyiZooCTb4xHBpzcrUPThVHy315Fy
dFbsUUrF4lavuo0Wt3d8kEjD11ERKMnnonv3Dug0ABWndd4bOiop1boeDEb9WBYpAH4kKZAve8Vi
iWnntEkyby5E6ZaR+MZe1DGRtSihbHoryF5+5rJBHySQiXmdIEk47OAAcGsYvD9CEL8VhuFExKEK
HTT1o/7Q6UVuk+K0waXq5Fnkc2cv1EdVTPWPrqyS5ZmL6wj6kGd2VarPSbE/WRFYXrr9cvPz+IWj
37QOeKvtVyu0tnZ2IyF5IPVGX25EHt+rdbNkgB8RJhJecuNiOdDk1Yq1r/HfeUnJDtA7G/+NBM6t
htcnxTAqysp6QX8hzEYuM4GbIird9sfAz30arGP1ChHfqvaAyRrODOS186w/iU/IQJ96E67wlT4p
SXUU1FN3iPdEKgEdudbSdIADqPEujHZX/YmKAJjfFjyn6kGml671Ub6NYvpz07Tu3DrUBfJYARl+
IdoUI/Xroqqnm6DTx8nczXG4Fy/gpneL5qPgWUrR5Npd4AIdQ5cTp99tgUIWcmS4pqhDSWFynw5m
sO2o7PBWXj1ueOG8mUziKMYQDOdk+mVYVeOx7yxCcWkJnO93ri4wsA0OU80UpZswUgD24hcw81Bw
SHhnTJfy5XDdQN+zsZLesEGc6dCkKdC5AxSOWOmMeWWdO5LiBVDrau4C6YQY9NuSqU0JLny+174Q
4ysl+RY/QwSgFYG7U8fD+xUZe24QdSUhFwnqEpRobbbSvZwjbSKiHn9lmYhq7NQFX0eRwDkH5dya
T11UPdKBCGJZDg1ANQRVTIPKKaE0z0xgMpqpphu3gunTXpKYu+XevJiYjRyuTvSD3kBmSm+jNJJs
vKGUy+H0EotfvmJVjKk1O4dXp1E3i0pAGHhXZbCgJcltqfJWdQJab5XB5II/0dGbUCFf16ucNlMT
G3yxo9ad0smc5PgX5O4P299ncQe+V2zN0RqMJslIlgeH1BRbSYWLXnEWW6GV6hZQpeq7gk35JY0T
+vusfKnIDDzwF3nJRMg33JfL3shBZxJrKsoLSYzIyM+rG2DPX3ng1pBy8mvwPZ6bdMeh3oev/+Vf
CJ4SilDUvvGgq4XSXHwWjbj+FZXvgKMkqVRPX5en/jrOVXL/GUDo9MlWuUaQQrgdfhth+ojVBvyb
Se3j34PpOYvvW+sfMFS4R46NcwB6B9GGns5unCElLZSNkxty+DF4FR1ufwPA2QbL7a+abMpWFkOk
wjEdVEl7kvXbwDCAxphbh+6qnHx4LH7oI6O9iFdqjSwX2OVCcOL18blXoebHM+OKNJz6pp4LrhbQ
sXnweDrYij0EdjlBANuZiv4M0rPFt1LTjOKT/nbmwbOQkoW1krSuGbdZCFC8oxvsfLFBhXHd+916
cMraDl0EB0mfETVDwGFpZf8YtjBfWLAp/QAhfl3Ej05YDWXlP0PHkuBpkfWA5IZeinwDEbEUuX3W
0Jj3Y+OvaQIdDg6X45qQWbg5TZGOXyIw1Aed1+mUy5FIJicIikeyH/9361yzlRerQv+/DOzvQnS2
5wi35Np4gE7S1jEIL7r4wKA/ZIVERBqx4p2MhBQDHhVW3VW2ac6WbMWznYcebQJMKcV2toaxnRQe
C45xoaWQH8zvlsGHiDOkOL+z7Q6WJdn+26+cUKoPgsqs15v0yYO+KjflglkDQ+cGeZn0j/9cpWtB
nTaf8a9RQuH0AbMaPExPMQGQq1arXv6RRerjeYHvGzbTRks6Uh8SId5c0JQzS0XX9Xr0AqyYBMEZ
5tDY79mZ6GNjcG4XLcCZvX4QlrIIMWzuG29lHrnzMJdN83Tvlo0J6KAmM7EcXBvzWycn3taGbUr1
hzpJ3+zwhbhuIxGBXFAWvJeDYDYlbx/H38Z+kBhR+VggetIg3UO/UXONqEs+POGcFXFsbKJA2+vA
iieyy0NC3K2oZ7kx4ei3V5p8yC3ZgW3Y+01uU5kfWQhkeTJh0VtX+6G7nS+IcduuxujiYJoeAJfs
82z0QVEZrnnauKRk+e92JYeREgAKrCLmdu+1Woq3IEwMsavvkzw6BNeUS9ErW6HC88bZXKx6FsZM
7a48ow/RuiivAbnLajtGDKit93jp3eZZXoSFmYlDv/U+s3QdRUz6F28n+lynMGjlAfTwBlqi12Ek
v3KkbsY/q8gUcVees21UBNKGr3IurZe215kLEtRybmjZzGVxU1s33eR6nLbJ3V/1Q+UjlkeFV3is
qUBYT8x2ebeN3mBdRgZdDZU85Laxuz68WUUHbCnWwgsK1V0HfwJnPaYXrXZJXEBlnmlvlEaDr59u
QE+c2tnZKrhwvKtuPgngHdOpqv9PBSsMQ8Leh6coL+EH5Xv+H2pykY0+02r9WvANnff7GiM+9tou
swg382Dyf+rvEBMujj9hAKEsmIndUQjCd9UNQuKbbBdE+c4dj3Lm3//4aEz0y+hzz8dp9KPwiM06
u4/kaSXhYAnSpRbNSqAMTPpt4ZC3ieLsAZNpFpvDCnkNURnfhqeMEOQRKSD0lSxxD96e/44Ug7G1
m3LWR7DyL6hg5ps2/aaSlWhDLkdCxa6BXkk+/rK29wDgzY/0aPM4d5Q5CMzSnZefcvOgfa676y4J
CRRYifqpsskuAw3o5ZaLdPu/Hr/hfHdZfNT0Ob8PtWYvWFwR6wYaYc2LN2HyDP+mchjQ0raYmr42
IjilQsQ3XEFT5YAlBgW6HICX+vugecbNMmDHf88dQraiouHlIj3UT7Un/pOo1Eso5Bp61xUVeGKr
GMRw9dbLDjiJOOLEPj45CZwDZdnHXscN56HVabrLZuAS5BXNHXN4BaQJ0xxYJPehXwORig5WxmNa
9TJ/faAaeoARx3uGAJO64sA21qHpCxlqu+5wMj+rGs2lLBkiYo1vFo1fo9rQtrwikAUTwrmE50Ro
D6SmruoGCAtuWdlOnLLBwg+TUgb54FxluZntlZlfCyl1Kh5sXwCeNAzFWj0UtleIPXzMUg029oWr
w9sX8qElCqZZBYhNbVla7L6wZO4XXyBwB5ZBuyee0+BSmzwZZyHMxDfsgrJin4K28q8pcEkGiWBO
hBiUBKWB+KZMm3DnqH9WfMeaeVZDB5fEPm//Zf0O5D0/kMgGxjd3R08WvcDMLOci/Z12h+B4Y/PS
KYskMYBf14jL6aY+NO5PYLtZcGcvnGhCZVE6oUruPYQEbRmaGM/7b9xrX8nBsy8rtZLhB7UQejcv
UYYyUMEPHLRwpI2gFj7o63Kd9NJlJNlhW8IxUGVe5ZWDgtKjdYlILjuTHASLXG2mhgCT2zqwlhUX
twQnOgKrRQfjQ+CRuX1vKZTAQZ2rr455GLsuSvWinVvYRNLG1HFxOR62XgJZqgSlmqCZDmFseogN
OJqiY/QtymA9GBD/rryovHqvnCyDjYurki0ZHteqWL7y/6pw8ZxXsCcu3LNcm3RGenZ/ZN8oKKMp
GYEN70L/kj0WLeMKLIMNe0dR2doMP7Bn4GJUZbemTZIrFcx05gdzruLM2vw+IBdYVbV33mDVKGE/
LkXNbDoqqie8j8I1F31YOpAeNU1namuIKSDAt5/C2ZVIsWRRnIRCieD4zDLE4Vqara9oAuKPZQTg
0+FvzDXfkyL2GVu9VDf53hQWdUPek7CeZeX3kBtLO4ZDfmSsjrVSzFB5ed8ECeX0kNtrv5Odgs49
lO/Hwz1RUz4KUYwo3NnYBHTuhlPetwKDqOVOk+O62W1b5LmefNju7KNPo6OZ3gFBbuFazwJi92Hw
hVc36/Aq+gk6KOojeVQF6RjKjVrwdcXj/g9RdOu4/lu2LRhS/UXRyBnLhictccXPJ2ypHHTbnPM8
sZBb74e4YmaIFi7VQToIaK4RQsA1obmmS8tHJVs1FsnJvS0bhn7OejCdewoltY5KrhnzMoRETE85
RX+vSe4Fshtse4t0BlKbZHkNp8oI6f0whmYhxurI6CvpB0U+b58etKzP9ZmF+z8YVyindPuiuXTy
tDbuE+RRNcYkG2a5e5VpZHthsIkJ685Xfj4nDo0f6sXv2G4Z0+gDjyJQzMZ9PuCv9DUb5A3KBf/I
9k9fkQyibUAOyOauV6SitOwy6nVqOolxM7alXidm/l6PIBY3Lnk47zf/sp6+9F9jOqCwgGm7Xxl0
Hq12ekGvnS2umO1XgJupNsMO6A5g5/uNbbfwPqD0HzRxxOTGY6SyLeVOqgt7Vq6Ime30QgMSfZg2
iMTiwLic5VZ7Ws3fCWZYiMKAGSL7SWTj3tUonSVNtlS5UdVt4+sN2BM6r1frcezDF0N6CcpOaMOz
Rsl+vYeDbOlmJICiJUOHxw+C2I6PryPBBKABwslKObXgxggf1Ueqw46UCfOqylHI+sh/5GUlIDAi
fsoxDJ6AsSTrLDLWuVk14NlQsFxuiuZThMqkTz92LpaHSTZ+L7NeYH+tswM/PZ4vkEOyFad86HUR
QSJMS93LODgwziA73dy0/4bncb5eQjY6jMQJA5MtZhr0+k2PV0eTYETTHsLdXIPUrYOH8GRuTA8k
y0+v6IX+6bKvmFZ5UNYJFY9vO9diIGwqrYNJ1f7uYVOnfsF0oMJ4UIX1ct/MkWJmSLos8SqGHUDr
8RIkNU85okOqy7hPoDMZ09hoLMU/4djig3vao9rE5WnT4G0ygcCDw1o8opPdhC0agZz/YjCDLXHt
NPR6Q2JdESzNHhnkkGC386OsNa4b9iat/Bx7xovtkaPyqjrDtrnO5L5Jh8UytEkfmbhXOdjaef63
YcC6MQ+8raLxzafr6MfeJSuCy6P8+ixG1VDeVAx1bTU1vvyZtf/NY/A4nUQYk7+39Lb+hRWqFNDe
rGKO73JvBnASu5vRB3LG3ubbnTTEePD9eQTm+P2ZLQ2251L+H4f5x3jZt8mnTsf/BSx0ShEWbFV7
wGB2krny1j5rvILxw1VUe8kCLxhFSgZruJy4yrZzf5bx6MmiuCpMl38U8hoT7ssFzPdWa5Yx+3f+
hR+8i/Lsqz1DvRDiinUXT8s2N11CdIIeDtDjJuoTC3XRVPqJ60OaMRd9IHdmVqoKBnBepBEtzfUj
cuKVqlfiIO2sK16Mkh3/HPQsabthXqdQyhDdz5lQFlGE5jh3v3YeqEmmq88597eIKVao3mByjZAG
HSzY+GU1Mm5TzdoYpOVI4hidtYJPiosaeCKfAYdAotJnEOAQUg2IU94NtUV7rSVIgC+0ATe77eSi
PWHcnhF4GOL2fO1UEkxrvk9w6XQW/qUYLFuhcn68n/pjJZQkyTbVaFAdyYuoisotC4ZiFpm/jbZw
hEM9Q5lIyXtKXtrCCrhemEtKElwt5cjhbiBYMikKUYuWEcRYtCGTS5ZpBeChoHXtzXQ+ClbLQDdE
FyqyzFxtiDe26VTBPIonWLLUxC5V0zJ/IXM59FiSfdnUJ11cRoLrC08z+6Z52Bi6LqZPoRNj/FYn
CUXIvicJKDKFOww5hgcG0EJIb7T3wYO2No5PdDPsRlhoNa35i9a58TVQt7XlXY/xNqLz7sMHSDvW
2OZHwlyk3uskrNZsAZNWiTSoinWkysFJ9HIcGw0AfwIx146cIL912ulkU2mmpgWSEQ/ggD0lLrYB
34hVD9TR1Chagw3533swKuZ59W+tn3QTWLL4pRcreVpmQ5LcEwq0L+GIhsYJ4Q8uec0gAWHUa46h
36YxqiXKJ+AuWDE9HjRiqBTqMAWINLfGq2H++3GTsfxnxvzjK323I4OIJSIAw63svNVi+qDhwknK
8HvKlaEwAi7Yf/7rtWZ4ykDq/+piadynu/bDXJUIu1Y365PsLe8/NjLQcrWeGPea4HEtc+jQSdv1
Wn+efXqNv1GvM8cCc9QtFzNxZbvNq3occhQs6Wbx/Tj/eS/OMOj717CBWF3Ru7I/FL7I0ESt5pwz
9QQtFFJI+qZnKHaqzndj3ouzvP/6+4sUTCeSOWFiVVrRsuRBg3BHwzhoZ8/88UO0sc8CRgvPwFsM
hrcroQoxl880n59hWSJSPN/GNBHG+zR2iR8q4C4mFtf9FfKNTlKSxbTVecG2w3Y/ZY+D8UsM31ai
IF1cr6Eyn4al88SPPtlQZxwqcFn0QaT5D7pGF72C6/VQpkk0bEDQvC5VMm7nTl84nCqO4HL51krB
aZlh2VTfOebrsd415yqWZ1KaJ6BcOajASLf3sM8x9Tg+d08SbPa8WJFJYLtoIzIrdfx/3G+cxasY
TGATiVsJ3CJGp4hEBcn6+SPtVbbQGwFSqXHMyLqLtspxbc/ZWEWSinEHFbFTOKneC5UWKHJQxqdV
vCJcgmcOsYVXEn3Iz5d8XqSuISZ38rAixxSAre4pYoz0lkhyd2psE2F4bFN4cqj1KUX013icEac8
WECBIcF5UImg6BXZM1lUj7w98qkz+9FbilIjLlX3K8qUq4GYoA3RDPBOTyTWQXnNRjIcS26BYDJ6
sgXJbQwKHBi5n7fGSTBocOXVUF1sXlKIiy3gAeFGKoKNZViSaM+5aojOdlIfhJSpSRVxsp/xvifv
kmr8ic5OY6ZJ9x6fxEYJf/3LtrQNlY/PXOUDjKcPuZNtMtxcFtmMaUwOnIhnjSdaXOYewV2tcjUm
x7JdgEOKTsA8mpcd3+DvECWPamjzUcQ3yrlVyrKmami66Myuzv0k7uc9jEkWYYoalITVzO76MUml
CTdRPrMxf32FZWLYvcXIeOkQ+EoOTI/sfiH8dfYYQTh2+vfH5WgZpV+bAi2Z2ijkHISYiYT6kpPn
Wyy6GeCzmhVU7qdEwFnphlaws5tPHONhgj/BhJF+/JEkrw6qsleSxpcgEIps3EiVNcjTM+2f6IMu
1dwoNr1hJX2imgFMaQXDpEI0BfLGprlDHKjVSVVs/baMBAdjDODG2wD4XymQNgBTNJpn67PKFbMK
YxWTm65T2skwMb+P2+XYAhT4fedox7+jFqRxIwhB+a36lgpS5riMf0aCWP1UHZz1PFlXCnZHhWx/
dFsP9t+fQ3D6xVkGyzDlV4pdmEftdS2kncICxpbnTaCb5ULZAIcmr4DUxi4RDhCzfCKp5ZpCjivJ
GiUb0aUyBsD4gTMCfnK2mU+DO3W2gSK1eeAxSVkl2DHzCKBN0VvBZHTxA9KAEKlfefP0VtLZa+2w
3L2kduJsFUq/dKHVq0TTaN3y+3Ng1RAoILx5dysKmW745kQqJgjvI9PrcsiTNaXcuuNAnODxVCBf
p9Ibq+FhPZJhxK6+lXp68fFw4LlTy4Q8wP2RRCdmH+/seGxM0sWJ6xn69JQcZ4vPD2kGB2aXhy5T
EuGHXAtNoKUt4MYGLe9A4j99KNa94V2wmPQOHDRItXlBLoZcGPvCUgJtHOZs9EOYclcd9ltDyBwI
HPI7yokxlXJr7InGxE4rZDkfph0ewosgWphkR63CnNwd2AZzYKM5olBvMqgJqsOfJOqG0+4qG2a1
vJsmk4T5CsT+RZj8kQJt9D+cMbVEx57WodIDToDHW5bc5Rg/VVauqse56D/zCqnEAvobiN0TkNz8
yEf7/nByFdiRfH+OxTIWDT7XA44N30i+wN/pMHfF41NKE4NbC/+kBVYySKOp3j2rdLK4IcWMPZPD
6c8Wqur0ePwZwVhA83KX+WHMkLNMLg9XYEXxc9aloSaDxYX+xHsfwkzHeP9idYPTRUBfVjjLSUOG
zH3Molu5vXAdeA0V/HyN7HLOmYvbZ9w4F5ZbnQUH2p+OBuyZXwspyXSJx4ZB+fPMhuKUwHgPPB21
k1/+P1rz/Ok+Y5aRLsnGJDlbMlikchymWEpF/jevVl062mDRjwT3yADQIUOlsljg0DCYqTFOnoH0
BRjKETvDsSQ22aU5c3eSG8CaSDC4/7OvdVINiBvYxcQmfGVSi6IfO7oQfs56w4qXH7mnh7RaAoEP
Wkmito7VNUMtKkT2QdoKgvMIP+4c8XPmWJqQbjupWB8ZDGB4yEcogg46+RIQjZaR/La7C7krytbZ
Ft4ngwPiLbHOMwARX8xvrOp0JtI1yEROutIeoXA76UQsU4RJ4uW7K9MSQTEc2iyZu6Hsd1AN7U1I
KzYGr6g1g3ClqZqG3fdadhqoak2b7Bv4po9ZzNK8iF9qYnERXZgd49mHvzMsg0PEZcC47UuR8A0v
O6PsQI4inLNUPk5D0qARnpgfXP9dXm1n80RuosRQh47FBBmQoPhPVZFN/my5lSjhiOn0h9RfZ7fV
ppx6M+g8951osKNHrUuTUh/Atus/b2/mejSxq6mJ9keoCEHFVxcKbj/2q/e8hKpMI59aC2C5FA/W
l9KUQ2kCZUb1D72VaCCQfwlnLHZx+ZplaXNhTUj2P4iPu8bmJ0QkMTQ6hOKCW6Y1KStTh4vQO6RT
mFPmrCWOMjW490EkeYE7DyoaZW0Z3+65ctx9RPKEq2P3nWEB1xrtpBwMGvhrxsMCW5yjFdn4QLrh
5E5GR1000xjvMpGOq9Yxu+Qk+TnE/RU6ny5HN/CSp25EfkXNBB7M3xlGQoE6vqJo3kaS5FgKG+bN
unDjVTQ6FILWsGQCutZjdmnBZxhZCOnPYCVts3AbS4S/cEaz/qQ5Y35g86sZM1mLQ8bWnwv1TxCr
i85cGzyBl2ZJFvcJZ53w9j4/st+JQgJPB4qjJcJSFCNLMzfZJ1ZganTcJsADB/qiKSq8f8jfB2Yo
Nyx+ARNxkdnbV9PnMr+IOMUf5c7Q6LjiODevpGdc2yCH3CzMv34f9IpcPwgLjNQlJH3RyYwSXzn/
xguC393P1QQPWY6Vh5WqOHGeFeiiDPTF4R26KHj+ic6o3fjwzWxj7UpELlueCAOrpQzIUS1Qb/mQ
N6zPtY1TzMJoXiiFZvM82O4O8ISHOCPN4Du4gxm2uEDJIam/SAO3q1ilUyJ9RgUqnuJL+Ns4kvZ2
SMeZMnaybNNDfmNRiwNGsvgLYGIPysuAaM328TeJe/MIdaozScOrrsFk3BsvCpzfY/PSTw2IoASv
IbmfaijBssKsk48Kuhh6gA7X+tDjxJBS8mHATnWy8hVpZdyIf+IUs7u254NYzdSUlFQvt6rTsxEc
1hRYb8DjA+JFPsn0RY2upfFM9rd3k4u/0tpwkKqdJarH3loVaPp5lR9pdd+sTAVxqYxzHpHgXcly
+SCnQAD1IDF0EinvbnTW8dwTHDdUDCWEVjIeSNsKF45G7mHuXN15k+0UWAghnBNXCtkW3LtjXbdX
OXJVk5muNy8O3F2Mw/LpJahXZZQjilj+pFfVZz148czTbCDnxv3Cpe2/R5FTPB4Z9c0mC9nQXX1P
xRSXKa4nOhS1+DGN3vBASfLVqCICjh2yTqYwVFhq1QreIXvQSyMIz0lBD3hsDH0PPA5ULTy8okT7
sT1MAtPYgkwPjv1VCnWFMLziK7HgvrWmStfIgsi71zoMoUMieUi004SdiWa4259McxNPH9ykwcwx
dNtrjFwPaGIh+4c+EPpjyZk7D2AL1xcON7VrYxHmAwK0IvHC2SJ/CTEM+5mpLjsweBRnUGaPtNbk
6C3GfPf79oVyJe3M6XqQmYJEQFiMSpF/UcsrKq+RnGfVW/kJCI9WzTkjZNgb8HH4cM4HbLHlAxe6
5HASVwegWTNiDZ+QstPINtT7M3wHJImk7OZ51AKRJHVR/CrJRA4qr2sr/xS6LIivsChu+PSq/y4U
bnl6NNhCx84jaiA4n5eGLmJlK/emREO1TIR8ppVjy9vf24ROOZZl5EO0+DiOWfROZZEzHU/dA6Rv
iLottueEagpTCzExdZKrkPwRPAaTrk4FeZVeD7SNGZK/4he2khNkQBlW6PWc1foeWXiOcmQYMonQ
aiD01vAYYhmZ1uj7vWGp+KpS2hZ3mYNqymSTDhhl4ZRbslrdmNVYm79mdHp07z7CcIgqbpfsfcS+
szwcmIIXBLS57YJndBOgoWTyn6hYMQeVInM1YTv3scTx77bevquTzvw7YAobqfBR9UqvFv+BhjeY
1gpzJ3AdhyI7veG2dOYpUOv1P2sP5jmVtyYKRUuYO/qqUfWJrO0d1hhzkhEcpKlD+HtN34Pb9YH+
azi3PMElC8/iO+1nlNrYAaSMgnAOxeIPtWpKzxwXCr3yb2XBpDj4FS7K7LoaUl6gPUYg/BMjcOmT
FA8SlZB50IhpBAb6yjfpXOBq7O90xPM/e8ZVFVo0bgeqWTo7WMn3ITtSlvi8K6oR2NIw4GUPT910
fIGIu+3CRzYGGwZ4G5ZKPAd1N4HZlJf5MpVeOYbut3Uj8pxlMMlUZ+4zqmaygceeEX5HZw9eemLx
Qyf5sdh36E39Qz7akeXneIvd3SuIj8wGULgXtI8/+eXxXUjWNR/epsoynBU2rsDUGv1M/EPqkNdT
EWfDPT5W6lbECIBsw/KPohI4CpxxzsYazQFefv5UXy0z1MALnKAawGUR/sX5A/DLyHO4IisSJIkZ
5wjBdPf0XrM8mPN181qHouTJad6rp1QJBslCbTAzBbKBvQWfGoJQSwFYzWkRsoG5I/fWYwsVwTZs
WPwis3xpBWIdoOfJvsWRpPD3/z7Govx9vxC4l0rr1HPvDOyeliLDSWKFSnzeVEfBesdX1ZsNqyD4
NpVs5F4CgA/5b+LcbNu/Gc6Sxs1yh3ypv4V0Ilo1TjzfIgdWpf2XIo85/8fYbK/PUJzPGoeVXtor
xZ14nCK0+C+PPEypmpdDmZut5DDzIjAUALM/sF4vkmd0vzUOQMh5YUWUV898K0Wpp2EkIaFUjwOv
99tep0gk1OGlsvbXPtEZxNA8+nJ9ql+apueQRje55vU35ud0GabF9+M46EhIAtWmo4BxRoC8qioZ
M6Zx+l0EVwBS0Di6p+eC6Wh7ULzHkXsyORHs0hzMBqVrkZiik9qpGR70hfzWDywQbYc6mRXBJKzG
8FPYF5hPswOXI5BCnywo+vzp6UeRrkdWE/M0qGqEXOnGihVGhsnIPsvOk41xDyIdwlP4wW6J7umG
cM7CgSts8Gb39WmEuNqZvOT7EMDi0ZFLLd6M7n+Jb5bw10lf57CgeI1pQdYKHU1UiqstVMBIeFwC
GsIvN7zWjMzr4UbVwwhTE0rqsBbduYFt/BG3TX+2wuxeJAolRvJSHgVOCp4DZhxmumWl0BT3PFe4
1YI+6rmLyPoENyke9dmGgIUTVJAAjouUwIs09qxeYK98WZJJcYlGofjadz/HsAcf/chqz6gnePw2
MQmpycrK94QMnYE7N9MYeakW0yDuQ/E7Ux4LLvbbNICsGXpHR0tmg1o8NMprii70CbOUuCc8wDPU
0SPJfBy3qhV/w7+xEBgt9IeIn0eleASOtmNEF1qYxilYuEieU5I9bvUwjvmWZhlArjmpdqEey9Fc
G/ci9m7Ajtu3VkS8hk5jpAPeOjkdr1G9E4aM1Qx7o0Ml4X5UeHsAwme5n3TG8qnxwXFEa42wUYzU
gEq8P17O0jPRSCbi7Xg3bN0yflkm6jHVPPkcPMbLk+mwOQc0qv7Qben/jOynu9LI03RIulZwX5/s
YuuzDzgO7oYTtH7JoQYp/w7B9sap9QwAONuVJKgPljPzhl6aoEv3dviXOljwxoFDKOSFaQPQnxNV
UndRvPkvM9uln83Ba4WZxQgaT8QXcWEcwHk9E1kbrLVobGVhiNvLhVcVcLhV4gvHTAYKOngmQSMt
JicmylAcTzFvg+yXfRoQnNergYPv6TfKTBVB0sgWLbC7OWrgmNuulpn7NfkGJuMvg4f0KP6uIHpO
KnPGMekmfQ78SjsQVBJ83Flhm4hQ+yb/uS954HbKvQa8IaicdrHgdA2AJRhLWBvFpRrTLiBxzTg/
fhV4kB5kZ7aOtDltJ4y4VvfpTyVjJyjd7Bbykm0xFoptVKdEDBVB0ScpnwRSU7g/wodZVjn2hxj+
DbhZy0dKZWDWr3g2cUtwHycgDPhJnDiN7nr1H8L3lZlVS51LZIiKPstTr1In1h5COX+VQ4S28/hP
0nDjYDjyYnyHQI1gmnRJicwwySXXrJo40PGdv3OKTWwKJLz/kNL6Thkg3UUPbWPDGUl/zEv8rcRT
UFWSkY8mR08HWJHmw9Kg1aFu80LGs9IJlteHqUAaBfYByFF+2osM/AjvltVgpxZtQBCJ/pvh6kjY
z6YIhlEtmhMLPrQpRYuxnTSN8Pq859ut+AVIHAOQnxMvIjzORjIuEDwiU30CiNgyNYnO+oxui4b3
7kjstuTmHWcloXJhXQwET3aqLY3q3QxiGaZn6iCxJ6GPaPyIdeiNDPUR6TAccdKefudWq2Tevnfd
bDq1xlmwW03NmV63cKCgslbQD2yLT8m+2Nm4y+XeiVTB+9uPbjdy12SRUX8MnXZ54VGuVydba3LP
x1p0SyGZsjliPcpQ4mdzLDrcf0DmRkcf/wi9+fSK2QVciFH5K+8DBoYggaQl22LPJyQryXc5D6je
idbtPXSjhcZfN0dgP7ruSH3eHCLJYFSe4fUvaJyR0cgGXjk6QVVBuGf8tajQAM1Vwmif3w79m7ma
p9lYX8uNcDquofiFXFegeptlV3hNn9xsqrhy/PtqwADOu84eNcT9/J//ajiKwswXhn5QNdu4oXpM
HT+VGCtEcOxoeijqAFb21gQqXDf76FRhm83/Lvdb3VFKMk9Yq3Cs5xpUgBChp3RJzmE8GetHoEPo
kVU8wvzKwLs2KOGSsvqobhAkG27rTB4OWedqDZrIOEuO5d96FnrNKyKoLJiVxGxj+fTjGzIReQdj
yZvqzW/xgzOS12bEx2vltaIqyEfBZ/kZJxcx4wEH9CCAyrPyLe41BzRzvAOict5PfFs5BCSzTKDj
vQlVww5JD09WbO7B9SdvmZ53FClP575VjU3JzhWOyViLWMtvvACb//kHzGRD6+xSGqM6Aw3POlfO
9rDVNyUAF3jfjHuLuWYBnCnxaqff+i7neUzdC8oB81ZE/fmwckTgfnPNdLqVNShi6iKlVeRHPJDc
40kNzUlCoEomy1YaqfhH2ppQNgUDcXX0yCC8wrB41SvotVOUy9cKiYpjVbhKf4/MdLes6uuLR1lF
W0v+e9L+nJhiWfCSTByYYTbRsGZQ9RJ0EJddx9E6gm+MeSfHVgCDtSR3Te45xHzZKRMHhUhhsVnq
0Xfs8oEIcqiIuSSq0M4xe/+bbQ/boXhIsbBi/1qsxsVCM1aWPLrgCS+GQlub+J4yYmH6jkV0BWEd
BveOjvTl4EkNgjy+1LSBaxWsT7gRjTPLcyX0mH37kUy7BCmYQqqLk6r2HtzR88YrleX8OJQsvLfy
ue0P20nwKLKh9/fZNCq3YDYOeh6ZHivSydNoahNoprkXQZ7aNP7SCQwMjJJ+HpTVYEDT26GqmMmD
+FnnE7KRSspyDNaWCuHZXrG5Uf4ewjUvtLPCzDk2cB4qm2J+oC5KgajKNJ09I58vQK1n2vnwvmsI
Lyy5Nv086Qhrk7Wd9US6p2uFz/XN/DtFXTCOikRHlBXmutlm5gafGICWxDL4pzsgLijS4orREkqh
OtQ9R0z0qeWLjOwFA88QUo9uHr6q7vRES0fEW2DX8z8NQenaBB+AlhxoN1NhikcN2tt7kbC3uLNx
SVuK/77swBwtnKjTmyplDUjb0Gm0KYGCfzOi7hpkICWhPIFOJPFZwFF3ULehoFP7VB7mtAzTfhSs
0pIRlUtvLdvyijd/0chlXfYpHGXvJO+tzucNL8HTLnGcHQzKG3Xl1s90rgjk1DZYPu49x0X/ixoF
yQFZ3Rh2GtdeTRw2uJsqfuP2lLpASeHfgpW7yRisKgYGc1JxPoDeXNVD2/Q3cykzQwW/p9hTy9Lm
I/xOnwUV10b5JvGCthxX5BCpsvAqcrXcrwtrQInphURt7jKsbWk5FgoRKVi2N9jo0Nj3tIzKDpwL
I15fIXYRe4G3khM1va8XnjK5R/WrYqqk51A3z52BJXpd80IOvwZmHfd24+Z/xpymXDn065SFehua
FFD5CDoe4B8tVuwZPTW2YBn/CZROy6BbxkHukhLPEjGg/k0SnTTulN4/t/JesIE2jAGQ+2OxnRcd
0i6Sp9E3R7c5mNZSH/d/oYcv8KKhfrNSbYD/KNMAj7STro7u+FLuaMGxVpHTKy/jwEmhOae2X2vq
Y+Ne3cCy3HFpuWNLtMwdJllu2vlLpw6wx0ksMJtOhIholYLgHAhc44EtYBLXXAD8F+0x1L3oZ8yL
qk6HM1UHjreER6zsm2AvrG1RHuJvm3TVPvv84QFuBdw9OK1PyRFNwrmkUPHnNl+nh4JmiYbm6d1X
pMw7B0nReDrwJHd0TdyZo+cpUNEnF2jRj6F2gy86me1vdwFh1gAYvDQuPnmtFWndKJ3pPlhuf9lM
nfU0WaESNuEUWjh88yKF7Bp6LAKXYW7O8XZMsmZljJeqsCTDLX2JvWMd+RHjrfhImb+3ymZ2kgG4
w3JW4mKXN6t+4V0HkG0wq+RyK7+tEg2/dAStvaa7uKSB9qWmRwjFF3BXxDqE74Jj3a+0UDKSMKCn
by8UNgIhAh7js0H5qZHEmN6z2WmOKh23GkcX3PXEOSQie4mKLzPN1QC2Rd7cbMEAXynGJ4A7T8iN
Y2hGKDFglB0D//V5SKQYPXJRXM/+SkTw2dvQrxr+P9xz0gLveSgqQt4SNRcM7Zf34RHwgZSE10eE
HkaCs9fRxIQ9Aq1Zk+qIZwVOJpHauV83BXQfu+OciDTNCXSIJSzz+XV0HId5JgSKx7vZNuM2xhH1
/6iNIxPCxQ9IrW4SA9FI5++YF/dRv17+zVQLUh3yBsIM7Yx1iR40pFLLHOu7KJNyGb7OoABXDvtE
PIERT2AFL9b0bUbIWYDMnRvlZhuEkhjghWNflrhkHMBkdF7rb2PasiLQ5JPPpEAVYMhCquWbodm+
KKe3sQLe91eT47lecQdWTuL1dJgieeLW/PjQblsSQqLn6HsP/NW4Ub1exz1mfrD5TVh/zByCfaUB
N6hPJn0qb8kxGrrsjeq5inMgMoTx0Lx6bKWeVKSmSyrFNOtPY3rI93ah9fqAIQDKtZ8LTC+ahoGk
Wvq+9Wroj0pO1oANa7Iu1x1lJsWB3FCJa4qgA82FoMsaO0oe7rhef2IjyCRfHf3UE5PqQyp8YfcG
2JtkxZhl+kmU8I+RkcA0zsuZ6WmWVXA422L1PcxNWUDMneTC4kzqTHphoLT3g85HlNTw3VH5D7sP
Fu+fAFfS26INceWL0tDwsW5EwPdosqmdM4sVSVROB8QReSPxAOS5sm3MulbjWf26u3DEBsLH9/UE
uzDtkZJWySVJfYMM136PiPFmikJCSsKVLMQrXf5qWYvuAHcBVPsfBeBeZum4CBTy20jaPpQnV40A
y5GOfRGlmExKEYLR9CLtrcTsB8bC/2gqHDor0pQhHUClpyubbGIFzZSqLDEWeV6pmtArAAEWaBL6
JdwmSg8Hr+pU+Z2dSCUTN0U3XUlZ9qVT5a5poW0kINYKZfJChlPcpoKLvPQx9LwM41UP7c3GffSW
eJSkRr5/zK/0qFMlepFJcPlCV06HlOZM54vbSjLf6NvmKgAsxiXjqOBIpP9F3wEJIYRZvmiL1UA4
pBuZUOMNToMWFr5cCDnXHJaFO280ema/rUgRSxZvG4FLHR4Veke2VL+VpBWHHAH/i918uH12RokD
Epk4x7l2vuNZs0nu4bipiV5M1IkOiCxW5b52Mk4vLR7X9C7H8jsefMmZ+DdTF1CgpGF/Pv0ydBaM
b0h+msrlwAuLBXA+coXtxVSsR48d7Le7O92HgTzYwf2T+45+fddsIt3B1VDfXcATNb1qKRtwg7Xt
0IoLgl4tl8alsiZU97JFSb94AxZuY1BxfRuq9S/DQFPPfmCS2CzGX4hJYsjox6FzvPreRfdTklt0
yw4QDeYU3oAt1PYy9NBx52SHAql/OCY6NAsqo0472decPHyCZE6Kb8lP2WHyJ7PknjLG0NVA6dCp
06vjXD190z7aIRLbc8Vo1FsDzZv28Y9tDvJnqEeY2wWxGjsuDPgc7AiDtTIn0CW7giuc1wHt4eS6
CepinqyevnLoPDFB+MGZbxfx28jx8IBGr/2bkc9for+EqaL+Xg38IhcgKW1p2RmRzxKKjujNeMX6
AOunBwYr/Y+YLilANUCnQz/NiiEpyn2hD7wmMaDE1zOXvex88+l63q+J/OoK3eE8Z8lgltCPaF5g
E4EElhHJcXA8bTw5IfCXKDSfap9Pm0PeI/k4lE8QE4izRERqB+ZRI5yIitrn7BttoMwI0Ohndwxe
1vD/ResLgk22ndogKUR1L5pth6dki33Jf69Q3X7YYxOn8WYGIgMPq3qPUwH5iHLiO7qkssue7MSw
R9axPQBeFQgxQCFoNTdxbdTBu3gjfBazS6keH/yTyHCHnvX8aE1qlACL2b8X2F4TNHFf683+N9au
rcD4GUQ0+Ln++KteOGPeeJFZiQtF8/yXVKmFr2AFUmu774MvMQeUi818RTMDmNCYZ2TZW3OswrzI
D22LhpwbDtZCCl5ip8zW3WbIk+WLZgcgLT3/1q2uDc/XEYzz23qiJBL7K6Pbr1JtgPG26jP4USUd
W9yd0sz1Y+r3peQQW9hNyvAKdiMMl5y6okgn5Yrmy1ZsVN3zdDHOm9xGqdjOQ38fm12t5R20kYtZ
coMQ0maXlrau0+ph0mejzqcLwcPvLBPUjASJ6SjKAFRL5GjzTi7rLd7AMrfNkPFRtLFwrCqAcg+X
XSwaS0ShCojfL80z7eMGl4O1q5MBY+EtaZDLiO2ebtQe4gjVKAzRJ4nrwMERz2B5rrMCKGUlVmnE
Cl5E9Ih2KHLEryj6Koitje1Ct+o9vMIiOLeMs98g5d2muYhqeM4Th9lIEj9TizNaMWXODARwWIdO
Wz4dwhxksn9LcdfsXdhtI+t/s9eLrCcyxAsmAue1jG7b3cx1/sf46v/SfEHXS0r/ss2ZQGZS8zik
50EFPXvvRfmODTh+yDz00Ayvj2ZiCDzSiUvyG5ZxfO1WsT/R0lpr5fDMRd/HRLgJVflFKwgqPGqy
0RF+IfgVYMQcbgqQd7McF66aTtujWgA+bWCqCkS3PC8Q7/hcQfN1kXyEQCUOhcvawu1Nmbc4B0k7
O4Eb1+QbaE4GYdJXvxUqScJtU13GcbG6UbysLQqELqVto5/KItFu7BeLUUJBr140LM3y70gFZI1z
K+5qXzme+EILRNcuUQVhDnxpVHIw+h0OCyp6c7in1W1FtTyXXEdjKs0MDit0G2MIKVr/6mlqUCFo
xPhZYoVVCuHPwmUGxDwUFX44lAA7rliKJ+CFrVQI/Dv8uXKdrgGly9D1zr+pLBkTIfNEzYZv1nk/
xULURDeNPPaPbYfF7B/6hqMaFPNEkXPOfpzRZRL4coRLKwnnSs2RmjDCDYgNXFpx7xjldx/E9Ji/
CYbiKLWbQeTnJ7F6GySPd/2qrP9gUdvLT0sG7CSMXKFb5K5JFL7pu7U6vWlqlTu1bB8g1Lm51HcU
OHNsGeldd2I/FzRriw6h6OYM0/Rh2XMrWWbANyy4wfYmMp9yK1DUkz54wliZuov2AtrYnqD8C2Ul
zlasf6IPwzjRsv2KsCb+v0WvoJhXUZLYfmJZswuKveH+CuMsMbHDwtok2uemoHmv6e0n8myeMZYG
q9xiOCUebqCcts9O8eeSeQazAgD5HSAWUGV6q2TAgCzKl4BpoZ0u65WKD1uN68ahUu2oyDwc3fjE
aElqA6fxFAKhpUu+rCkVddpShElXMNTy5GtmmzyeC80K9IA6vK3XCGhN95zScsmirZvr0BsAyvi6
bJLF49bgkXEQ26ybz/s6A25zOAb2RM64u/72qb7WiUyxftUR7EAFJL9ffMxa0J91qkoVgitsxiOS
zQ3vRcHtTcidkxcHhmsop56hyAcU5pJMgENHRMOjYrbRHq9NJoSyK2S5Xk1jtPqYPGiMPQ5DNLZI
fuT7VgH88pohE7CU49ZGnrJVw+WVCj7+6sHWWnzgX2H356kJbrmGomoSQ55vqmr976zqRa/SBG96
4tc/g2OTXbuBH5LwIk77I86PvZa70rSQE2OqBxXbLBwvAyTEVXIdx7NfVL9Eb5sOfNkqIWUA+Cl7
g34bQ08gLKrdDW42MtknrQTWqltXtO3Z6loQj+atTV+oqtULxrwF1BlErqfdOgV3cjtMKLYd0ljo
7gnFSk2pJgotoWQwUI//e20/SqKhBBXb/BFIkwSSonhD82Pb4Q/wXVe4tU83INorIp2R4OLFsrIG
wNhKyWMBV14Rkz00YQWFfbwvCBJjSjJvXESq3ciSlEwn75iFmEy4t45tpWFoq92ygMxpPkumd6aT
Xc1+P8k2ane9crxvs1UEuzh2IeuW9M5mhTgX/qkkdiGZ8NRCsYtB46lxbXrN6bUyIPkG1rme1kge
FwL9CbLqfZ1wfGBEIoQ80K6maJSxfyjHpzr0rBy/m7yJuZaDoguWKsDQxrtwc6d+lDIsiOzSygDU
zBa909c5Z2r+8Oz453JojytNRUvVEtnFU3tcPHMllp19hXSR9KdT/uAthS/aAdgrAGzWWACtfVky
PmuqNmWLhb4yYMCVDb33TEwEcjfcJjuSD3vHG43txBfJOqseG4R4QLgDRZaazz0CXAdbjK5O9W8k
25BXD6+UO5ZWa1x8Hrinbv4ewZlrXDGcudUyd0HXionA9RPtLP+lqWlZfiAfv8D1TtENr7y0Ebzt
hffW0LaFKeBKTDXY6BtOXsfEyVRbS46klok/9JeBLUOpj6z03O3o1ZCadjydwM7if7l4A7u96AAw
JSAmAyWBWlR3cYri03QWnpoc0ZzQvPyhWDmu2g+AFOkSV2N36X+/1NzssLuveen9ynXN0Ow/KMyE
4aGjdCXM5iT5vtIXQSpsn4+oc90L8YgMV6X3IW7y83O2BHQcvNPKc2B2qorAGjo+9dX+BJazpYz2
3N9Ok+h4mKLcONf2OGhIOMQhzrIOLkvBneNSwTZ4osL7+FkXs7lH01hhR16CJI3+0J9RSUCNYMpJ
ztG3D73av3fuJibolVBiUCWyIzumhxxKKdbdTvMG1jQAUzLn3WynzYvf1AR6BKNr+xgfC1+bAj+X
nbU5Dv4IMMJuKbWN2e0P+7PoHVrh980yJdDppJ24lNZ0boCjoPhJ+ww+SBMxogSvCByJWICL1xN8
72VogXI/co5pA5kkhbCFALl8g/BXNkmO3W3Qk2yqGHjXe9kS1vOxr1zeaJauz6QVvyDFmBQ0LTM3
wz7fGL48UkaqzBmk8z9Ex1JA+oFQPkLGPFTBLbyjpEurdiaB550466MY5tXETs2JdkLStSOeyodn
r7Sedc8ot5N9uXmCIYS0TxAfquAo+ayNOTKQBk8Y3z89x7rOXaZkVcnnP26aVuZ5F0vtOQS2pd9i
BMSqpLhhYFNm2rALGcro+5DziMS8f0ZRBv51EHXI+4Wk7aehbpO/VjPLNIbG2R7cX5iTBUZc5tet
mmmzaspXSi4Sl16u16rtam1GkOjwf5kJuz7KpT3Z3GKs4P5RAS5oR6OEVeKXaxAaR7HMPfpLgoEM
ftfNONS/u0lFee1sljiqkpRj4u0LN422+PMt5esor0zT9MfFWGDAGK9Ou/ulZDUNUxR/MQ2ymqjI
LZ45/yXzHn6+i+YuuSSLeLTG/Yo78PHQchUr0CoCRGQId4xeNoRW6EJHk/ckgnh7Ibf/KNlEHIp+
0Ryh/EeVErTAZp9xe0zKuAx74CZZIIQnQBrSVo+pvTLQC1/2f12LLK/gceK8r9Pw727VCQZ/jI4g
nNVNCMhV2XjQwSEK8EQ/rnSn8KJMOnLM31UIoxRKzd1be73hG33R6mMDbr+Iqq1OkB7F/2HHtQSy
nPtk2412rBRvIsF+pqgZjx9QqfqZoqolD/5y04QI5xdJzaoCwFLlvmiX+PwsRyiT4gtOKQIYARmH
6qkDYssappr+Mqg0nGY7QkaF0lvN+wWiJNY84Fu1vrn/gkFD1Pyk9eDkwYVMor1+LWa8U/pklulO
A8lmdKCQC+t6OnSPeAG1jsxzAg2Eu0pM1gwuurwzrbRIy6fLUfAO408+Cp+UxtNDHKX+ajvJCg5A
1Jz9xy04adXJEpD/CnXHW1nb6IpVliPhT9/288C5SkGJ6ZfPyTC0Lsbai20lplk47uhajPHPoQ8A
7IIYGkfbzDdfAiz/xz26nXf333iWkkmnBN4XA6HTDKXjUGMKjZP9bAE7gFN8H3lz5MHxYAY+cHYR
sdtflZ09UFEYZQV5h4PLHE57iGa00RDG9b4pAgSy32D4KjZ7LLzFiKly6hEuN+jJkeRgP+XfmG1r
gK8/mBBnM7uIaBJtB4/dA7vMw5i9oykA0yG1l14/NgLq26Oztm2vmIFV/E/AOLKQZDVCYr9NKyX+
d5lDcn38IPGKDxaRovL+7ZAJ+2cz7tm7CI12Ru7lbEVCK1qJv+vl5NbohiDKs5Tsn58RHp5WIQd2
jmmDsead6VobUpMijB+ZICtBkpKZjMqAAMBID9wtG7hNNjs5mWoTDDgGa/ex0GEIK5KTAAMwBGff
W7KEvGEzd/o9gDgu+giZJiwg9CN3fSOVM/v0ZqaKLNVX8B5bKSdQ4/DP5iJrjRtpHz712NJNRVAm
EJgAwhR4Z80ETR0UDgfM24+6uK/kk+5cKHc+3s6Fn7hH+UxboVGNlBNw0yNqNKyR25ZtaeWbL/8V
26eDbcbD8vdDnTcTV48Kbt1c1dYDoauZURkNXBZbnG3TaNYlNZxUlznCkbYZ0XMwsigDVQc4iOmJ
P+paLrp1lWZBuDmuyp0Cwgp8uyZSRxVq5Pfh+vBrFTSlHdm14Y1FGqvraMF8jr69AuIVozCnpvay
isAZGkRJCE0WqYZHFN28zPnumaauiMIVGIQBGI6TwU7mseQSS7QQYNnv/9wRrtV5hZA1VTvyDT4j
ljBd0Cy9xzURoOCsdoYqFMS5BvIPM3N23anR/Mr4lM6welcDIMn05jGX7Hk0C69tKp5yhe2zRqwm
RwUonJrOER0xn3QW4yrVlG3FPhwv3hJgem29MPPYkhFzX0p0mMnTt56gBw0mRDWZnS2BfMAtEgkF
3ZgtV5LD17Oq1sGECivNCIlbPfdGh3kdmPlxdvL88cgVA6BJ7jV63ze/BkNhwwHTBo5WJcIcPSTb
emVjQibNEYpPjKd9+VTu1p1WsbYaPc++3Qy12Vg1rOHeMbwzkzc3vNrlS3WLWe+cgS5aK8KOotFQ
mqUqOCMnLVA27xD/KJMBREA0gBnd2wbm9wxPSQCTUfd+9KwwDWtXwuKcMtFuyw5QmoXFqNwBfpLM
HMcywRxyiQqsbLfCZHgdia0v8lU3uBxlfNcQ4QifaKTc7u0DSnvraB6hw9rsOEgMsErt0hbafvD3
rK6jzqrIXypIKZNTLeIq3u8oh25vsdygOzgp2dK8X6bDgVcvP9BvOYHNnGERw/vH5Hf529yP5PWx
W7H6jZm9ouQKueIJSC5++JnGI2LO6tV0rfqyIz1W0O7TpPyn2ikHeAPoMVAHIB022Z1bnhf3K/W7
R3xmhPFqM1L6X40hBiGb30w8AoyMzT8GXm8aM++TqJyaGEF+2co3O5qW75OD0OdxMksDW0rduew7
d8xcmzV33Fw3ysm989375pZ63n/9dkpLLoyd8QxzWzqS7BQSbAYmGvzOOebd3jph3poUIckHkx+D
HKE7HYc4F6vMo71yRqUv09XlxvlDnEVX2cGeiyssBM7E4bTBt4+5R7nfuF9+Ubl/3bzQua4RKyFc
2/P8a+i45K8lHBEqIxtuX2cePaWovwN2Wj8s5nF8Rjk2f6YvPjZJKYJgyubgWeDyi3CXsKjsrmDh
PDA3Frq8qGHuLPFR9jkHZ9WAF4l4ZwKIqAu+klgkjY1xYhgEdwdTZS5RF7MDACOLJLI3A0+S1Apm
lGHBdUsnzWf4EwjFLgqkhMzUfguaraBdTIu2qhkbPvPT6S5YxmVKb10NBf09pcjKe78R9M3H4YKx
degYQhuKcry1DQe7FrANFF/T29cmr7akbAQVu+skaQ1ZCWsb0eili2JoRBVSvD8boZKIhWVZLupp
ij37CB0mNTSfOu/VEMrPknclUzhoYcR/sA/dRCl18E+RCFeZX+exCM6NV3zaESyxlcUDf9DU2UNy
gqSxnLTuscsaTn3X1/nDxtGwCz2QK6G2YyBm9puJ94VmiSxNPmaWnE4REg2GSF+vL1w6yg/+QdUk
NDk0cbeyXEdyABQiD8MBr4WAsqLItF+upNj4e/ZAfQtzGewr0TEMkeZrR+5Thpjz0WNSeTpEbT+p
noB14Q0I28WsLlFsG0ncJFr+KtBxmeUoSK//Br1SIg3rdjf+eZnS1ppFPPwzzqTl3GaZwndCH4Mb
PNuTm31mb6EiyqUsMNcv043zdMDa4TQmWiU7MgymVTnGfIH7ecfAgBd/2IvBpgHVlqEB98+PH1MS
QcvcYOeKSlFMu7PU+9aYOXQXxvMtReAnV5JMF3hSjQ/OsB7OaW5a6hverf3dSo2+b3TRpAOG6IEK
Gst9Rbt8CgjwvgQnUUBA+/HC/zsUqYDcmg4MEwGPBo16anmHRfHOxw2ao9vlco6t2pEeha0uGcVb
yCSevkBM9CiDxSjbbzD8H9qkUHmUSS0H8XWd2y/sHBPzuhdJ4HHLZpOx3pBMkW2ORUcHjEyuyyAX
XyOt37rDOv8WQdCWj2vGtf2FcLscNo5eoYOngqwDClFBEpANq2yLlhML638lGwBiGHpxJi345Z8d
EekH+NBtf8XRgUGwe2GJ/Wc/II6dCaCY0/hx8lCNqa7/bS3oyMs93OVIx3VFXrddY3AVsoveaNl1
gDEkX8DZ2ByBgtPKVwEx4Oe8yU3M1cAxKZRETDJUfgbK1OhvOV96RUAuHlQ2aujspwOBwdITJ561
dLNHpSFSp8AVoRYWoCVayd/bkeU995hMTgk4HNJDB519FiXjx7jY7/2/i59+3RVqBnaGJv/Uqz1+
IPd/QNrlO27sxTyedbREwzoXvimCEnvRyMmrS+sOxH9KL5ZWRmNOaBMu9HrV1/6av257aS33Yv/F
iXVB38IUkquaEYU0lOCqhfKXlGWyNpHFdtyv/fa109urvR1P41fT6eiYB4dd8YaI4J/FnZ0rXNnI
x2MfMKWZLOfyfz0hutv8635EkOySEFDWnwjmrP9kBfBWXRks0vYez5vwFnWgvQ8FxrjqLw22rCum
0Zv2VP7RGZ/76jpriLXNEqwrXod1Z1TjcxZGqP/Hv/ArZMkbQCUMFm2pZb3XARGRDbXk76IuDCbg
/a/twNcfzMIhRCnzrTbihLruvX8ESBQO0zom+HthXHkBI006DjPw/1YGkC1mYDwvV4dSSO5qSG0B
QJUDezj7jUEAO1YXkMGy9n2ZrDJAUjIpPe3ev886j/rfIDkJtdHOP6VZl9UZifWRoDI3o60tbZkD
hIYrC/tGEcGaYoGbjHS2smqz78ZpXIjkdovcsOiiMNZdOlAI5jsztS6Be5+X2EdJ8cMrVr3U7FOz
RuzWq9WeDNWqBK5GKOlD/IfBikdWtTQF/RyUmEtMkq9i1qB5mwUWVQOG+vDdfMFwRbwGepE/16B3
vzFYjUGUfxg4RY6bi06VYfRsmAT3MUFURq0sr5YMNHAyCy2DQcQj0Nlwbic0AoeqSHPyL0TITIic
a/dotS1l7KzKK5fTjAu5x0qp6PcwyTIxbdxfIuipyFSZK97QWn/bqxxn4gK/59/U6EMAposygSmd
uxV9eIswcIa/OE+mK8aIPtMhTAl4p9ZXOcqS5i9s8noMuOF5yyN2HuKS7zfIzBeVRowz8mMomxPY
ybHkTx0O47hepmcBL12oBx9e4AZ+PTWAqkKuDx4PlcZoK1+XfDs9c9iFYEIIYxPSiuU04dk4Mpnh
cqtjPR+pk5PlgDvkduazWjcjOoNJy0ibtIsvAfHEkWE8rifN20iUTFjHtA91au0PL96MuoAbblP8
xBWlDPQcApd9z8CzvnulrNqUg4p0ypdQteiuDvodkfiZ68zskPsjmzMqGCuML+YfWiMt6Ajgg6Di
QFnu44Ks6TiLiMNSlyrzGSiP034IxeZWaGeHohbOnwojSss/O9u5B8Hnv+Ai+1aMiiygE27rMI+M
msJbtIEsz7wMMwlCR2rJZG0UxinZUsyYNXMWUwn603AnxDxJbPUUaUb4o/bVrimL2LCc5tiLV4pX
YRG5MRVjJGZiWQS2SBfBHEhd3j2my1jFy+TwtlEx8dhSiM+MNN1NHaiY8H/rq5WCDjhkuvhtHqr5
fJh6CIC8rXSTRWh4AlgomB2MoxgLpCTorlwx4cdWg/wQXV3WvnQ+vCp3B51rehuqiM60NkZPDUCQ
4RmNNZEk3bQYuj2Dt9yyGvWHCwpp1XNs+AkoqqiwROA2q+GaOFHi+xYocTV48JTEYakBpk6bEBSi
kHAZtxG+g+YHVZn0hxpsWk+YT21LZxTqvRyB1STMrhszZLH52hKirN1cTO/Ikcr5+wY4A2aYwQaA
Bkbsx7fwjsj4/nvlxeBpyt6k6WsH7TXrz7r9BSM+G3whQC2nl6IxWMkqmIM8+8xlgjU9uCTXRfnf
b+pi/AKOlrZXTNwh93LIIoICNzddzAuUKIKNVDfwBS06adqJCMMrnlILD3h3OcFvk0gd+y68cQ6K
/NzFIoadlXvsq2g4gPdHpSb0rNav9eCmUW5jK4ZA1XshaCIUuzBt6p0zUH8k9OjztGvE9ME63dNY
wNtXbL1OMosbnRdO2+4jMvh2YajYFg1P0x0FGQcuUB/Cj2zwaU1HcDegaGurgpENVBmgr6mdumz3
qyWcwvksOIRxE1vXwKlmINiUAaC13DX8y/kHwwF6ARXq06384UY6L1cYN80sWrtpDdCOAJfNIJ2n
+JMJd2ZSQ9RaEzBHIruKTbihhwY8lZuF0h1WVpBWP6JExKkj0qp7JYF8W9UI99D6IX3ZgCH53O4V
E1kK89KkrRp6vhpVbWUIhJCeUmcYmNMM6CK5UMYcfxum1tc6fjHpf0tlrrLkIWVnv/Fn89saQaCW
zYVyx87gVYxP7xdspXcm8MVTEbyMgde1F0pEyEqBwDSN1Joe/jf6/ZLqI3wtFmTC9I3qXjuTU1pV
X1djzyckBqI4UVtSidjxIsc49DSbIb1AvzoSOw5iQeoyGOHqY1dX4hbDeJZvTiPdRaitQGA4Hzav
q5mQouASteRW9Ey5HRhHxoOH3UgqbCi0U3WOW36wtYoUP8ATCZNps+0UJIhOrCH3EkHIxd8xK0jA
ZLZ67laM3W38t4xmSRTn7GX/mRwymkHfkOJIYYImyugHYqScob4Uxg6rb+05NBrXdR+AlXyb+vhs
a3fLxO3cbRMLZr8fR9SpCH6PEkBK03lNKQjG7dnUYFCFS1UXJNMNtb5NMrzZOHpvFAqGvycw0I2q
LThnBeN/bBMV5vEQ0I5RuCI3PEMTUTFtqfIfjlLHELstuLPixxq1PSF9meMIuoj1ZaTCPJwLTdiX
tI1MMswfsDvAgi5rRDevdBnz0xDWwAwdJFngZ89RjGHiqy8CKiRXSo5dH6orCngPaC8tD9EMtY/Q
VviGcqOKFshmAyph3q93YkcVgS7HurXBD4r5TFGhxOJ40mA3D2PG/nS7EfCeq0BhEcxkc52HdiX9
Dhnn8ps2twS/dF73xjwaKI3H7Bs+tS5mqroGnhPJDLcqi/BipJI5Pc61P7MzwaU7z/BzjouxOz3v
SHRjuaxW/gfWL14B3hpskC8TXSxg2swW3gFcmgyv1nVtJUaCWiKWb4XqeQCScG03MfFeL06rPqHS
IACXqwceP7v6LdTf2EOZ3QfugWENYdfm/6KP13w8bi3qArtUKf1/XrIPRCLS7XnD9W/6dMlkIGaS
n9Pi+je0N7JtFd67RnIEopM4hgWMUZuGsiIfoJWctT9sQ9G2UVo8oEukNn0EZvQ75Wt/+i+N5ElC
Sz0KOFGw7mIM+EvRaEzeKLA/MgMNZSA/rfLjEcbNVGN3/sBEAXAVan1Go6shXJaK4s5YoFnJI9oB
m5afklQkTm9nruZD8La9H4Yt0iLWcYi9RgoyVxbCbOZnps+RoARJOrARb0Usj0+3XX+AzbqTKN0x
wKfcjH81Gr+/mz9AVc0Jq+ez9Onsrn7AeBfx7ufOeHD47j/Yc4PhzNoP1nHstPRID1EV5DBNVGdN
eSTyDgCKvJZrfG9CAVmzY3mNrEBYbmvNwzixGAf6A4uP2nC0486EnCgIk3WqQgOssB9OImLbUCFa
Cc6YTCaWEwBZQGT/vH4EO1nZlEEwvtzsM8SXcZfO0DHRsPyf07jZuSwx9B/DIkffBer2moem5RbT
LkdFAXiTpvEMaF/aRwhEAAl9SocwQHuR6es6Ks55TUOSCBCJj/awyj0ZIbyDmWK4ts5G3a+PwiHM
lJ9HxK5XUmCRqX0f7Fi21Qz/4u1aMxtFwZZv3zIgi60lkGR6ephKoypJsIjhNCQ2Lw8YHzDzitZ4
ecspXWRh+FGSQBdmPBTmIQpNTHlUJ2WppuM3EDi6EGXPsSrHkgHRAoaEzd6MsfTk4I1Er/r7UMV+
Lp+Mg4LCXvwq66qs9+ZXPFurT4e7U5siHm12WkVS4zJn+UXP+BiBxWL04X+GJGwUvMj/h9G5hs9c
1CZiRVm7iC15h2YY32sH69nAjWo5+vYonmOZ+X3blba/kKn2paZePJ74gCyshjqwnGuak7Gaq6t2
ostD9W3jZhXRFdGxJ6PLHqCKd92Ya+Sc9f/cUd0EJxl6gRig9uJXqtLnDf87HLZeNPivGjRhR2xq
gyGO9xiCrQHafQC0Ut4WXZQIAvr126zo5RnamFz+Mc3EX8mK1jvhC5pV3BhoWoVdmqNix/sOg/Xs
RJVODZ0wHNvM+aJ/QVl7VBLmQSZQWinV412/mNVZ6Q1IpSB1ZybpOwOYjRw0dNlncl/bReUGJ3sj
K4PekZbHWPttvsUaRLzSLXuhGBlU79Yd3OP8KpFN3BMAfjDp+/2KCDSdtaGql+kq8akmpXg5nv4E
ibBOBfNkKsLRA25UKDfpAt0e0zWz0/A4xJDFeB/hqfUoIw35dGNc5BbvpFO1NOChx5+vUlRa9qQf
u17GzG+FdvMbZCKL/BIP6FKK34CSuHrrh+n6YRTTkmqYVzKY67GEN/tchVoWKgil8MhGB8T2TNud
1PcUkHM+TnvNqZajExVTu9v+DsYfbh1HI73lUfhCrnfM1Fo04xItJZ0bWyBZRFzZ9mhfYGyvx6K2
Rs4siAYih3YW9arCNQSbpOMQpgfQ8owt3VAHdhoAHjHGRxREuaFvyrM1Adp15rlQLLKO5kpG/2bZ
AkvfforAm06bHaq/mmmAz0Ap01fs8lmO20uEQdNElmR4GW97gOJMnH9DunmSZtKPu5tWJV5fJ9bJ
FAKd1NCHaVCUE5Z5LzB8HVVhtMoTp+5n5kFLKQSn0EVZYgq42ZhFLWxLo/CZdiDxbLVo6lUCPDZR
OEawLk6MAGBGiJTsSfGtCdoVPWbtoySw+5ISt7au88a/CDphMhRrvW/sHUjnuUyPoOCM01Z6BUMg
/1M/p3AKBUgA671tspuovp1606e4RrTd52LODJLusAU7FLpTHUyrWUY6Hcd5hRK3QDYUKHFEH4Kg
TthzCDlom0rDXLat54ZYtR6K8R84ifBxx1sW7zzRoXMLrlTcs3UZL+MCf88ZdLxXfSw4xYJAsbaT
cqxDc1MQ5pAmhqshX/dVoSZIZqDd7BakjKS38q1L0EsKGAfdtG9OOHiayAuTE5WJR0g1kFsPPWzY
VkMZURa1k213vCz3ALrYmjb8pUFHwYrqplrdGgh9UbSCvUQnS4uk1d4hKKkcu4uqzDBxVht/ogYC
B8sMqvZHsJavvahZr1PtNGXgRUj+c8y0hTlAMUtTysC9TvBgk5VeECatS1Ees7iLCYGtW99SDq4H
HEUVH9V56svW0OKdE2+eUeDs1nNBRu3pLbazQPsbIhYX/pULjYNmnFdx4Lyu5zxLuTZySCYSyVIB
MF0RQlaop+rRqKVnncWrtJnhmYHupfdsLhD6gT5vepuoH2aZW1xI4T5yK0sT2yFVcV5FiQvJYaMI
fMMZKbrNGDtw29q0bFQrzr4l5V90fnayHRoCc8AvkQQgXpEyrYSaDF6D1/4ZwILFzGH2f3gmvYur
kmmkjVKqn4MFI16hx96z/Zy3tjx07nFp1YG9pdgiKQcWv3eZECocVD7IBXll6zRgDXq1z2lLAHWq
4hev+8bsdPjy8L5ABF0oAc2JoJ4JTUVS7DDjHl4a/rwcF8LCy8AD8iM9cGBVm8xvpPHUhBA58QK6
yM3CB2CB3keF69jWfVH1LCA4iuQsxPxg9nfE5Tlhu4xPDFZRhetkTGltIge2Naqpra0BcYVgrvFB
3OMSfbpjxF5KOClgAqZicH9nJ3lDClkhqjvJDbnP1JpSjypEJTz/9s2Jx7f9yClv2BvtHh4kTWva
x9NFXo8qK/TEoz94YHMMAp32iiEnqfjJBtFGYbeUqyfhQ4PNCTnEwgHj39n9AKgQWPK0xDxX0nJP
B+9mQjuxuFE1ko7Q67TNsxjHGPzvZ5gxRzBo0VjxQ9kEG7R/8V31NKdfPwCb1b0vwktX4B94mWSs
KWJYFmMWqYWuwT7S8TCUnVBZ7xuB0GZ7dLf0edBevse5SjWEr+U8gmaxnFlz7/rplAjKNdKGGRiQ
Jka4WCN/FzooCVKmtmN2UZL8vRrP5XwScFwWmoI+pDBmHLNUQvlzbUM6F6KZaz5fP8hKXMRd9BlH
dbvCqH0XPI+SpJC4cKm94DX/8BaahWhyQ2VZGSIzsqlw5ceglsg1uAPf4fa07hvKl3Ea75HqXPz2
ZTZKJ5cjOyuC/9cbqMFCuKnAcraIfTDmFpcxMTuws7pUS7YGOXroq5JixqLWKFbxyxL4gXd2129O
nzwonJvBpNdCZbmGtvTcoNenQ6f5q2Ixr9v7AO7UxqiS5U6jAn2b9Sqllwl+63BVlfriqxLPtM6G
zn+v3RiYPf64cwW9RErsidLoWE/wwaFdg8oNrbJHqUqKQFFmm/33Ilm9fuYd25FkrzgT9Hbmq3S2
gnEIBkfUOCKo3sdkBKS/3UDKrLjbunV4V2faYOVTQETmnWltIdaX7dnJcxhduemitiool4QeKc+u
vmlLW9TgqdxQ8BSsEAJjLNFadS+5MVx4lIyg6ex0zGtOM66m8/Bd2GqeFxKy51Bw+SYCpO9zOcES
6Sn33+ukZJyLfk5IRrxCutlLbhbB3mtot9cwIp7Lb6PGxmZluh/6nLgU7hbgAz4qGIDRt9zehjw4
Slmf9MX5T8SwTIxkOR/CkGCR6diUmbD1Uq+NuGFsoZTdkDGmzLeXyZacZZwXicBoLmxBiRG++M6K
aMIt8q83zWKO8NXM00IzeGLkIWfuzaFBXw2p//R4i/eFwNamBX3sLL/or2QNXS+sVuDfXGobZ+w6
/7EVCL0qxDXELafuiesei4gxg7LmdlIaGqvJMcdRiqIfcB20qSXOq1zuIWhBqclC+uVbwQ74kk1Q
CZ56AmBHlWw3ct++AUYKPmNA0WUMSQSZNRYxiajGTsyHvWxyzdUFU6JaxBEs3pXjTQ3e1Cpy1pM6
rywTz94UYo9yeFMKbN4anCrR10wfPInS4FdJrkAzifVfpHNcO/L3pxx1U6tZzj/t0STQj8Jfj7zj
1RnYa5flt2m3TfT9L9ak0d0V1QLvA6VksFD8xm+rOxt6wGH3uT6NIhWsQ7w7wQJIdj1NLpPmcxy+
b6MpDtWeiwhiFKjXTF2YyXhJBb3YnPJP+dLfei43bKggfzSwmRY5ckvhXXE5SCqNmSmltVV6Yu5V
i9aMJpexwnXhV6f3VlvMPc6ShL4XdT17gztc+tsfZljyel5hPNMc6ZwFvCHSVVhIdTDhklfYRq4Q
ehg0E2bSFNNNALMOr0PyAUYBVnRDhQ3hT6bq55wprcWBe3a4nM+OJlJyzj7P504e5SMIOK2xz+fx
tZB7036WRKl3/E8w4SHy+R3GuVeJW+55U9xOmgsvyN3XtKelfyUyP8PSpZEUtrghOgrEnK6so+rh
UcbTqAMwfJN6p2Dr6L7yCugVQiwMnY2oYSKuN5ZRFJRXx3hXTDdlxSKItkEsNQXyMlPWIWHF3DCI
BJfp2gD7nw4LejLJoADX2lQKidn1DFDlnRhMwyjy9E2JhDW267hkfNIlQEysdUo7qC88eLr4tL/y
dsnmex8haq649hGufSYwD5OiPUg4w0rD4ZvL3QqSbFm0V0+p/lsLKQdQHjSbWimh+tpn5czucaOY
Zr/yVju+pxDS5J6PexIMD/PWsUdM+dHr0zqXEFUEJfdWB/MwNxguT1IpznM/L66521VMQLzdUn9m
FDs07CbHRJgW9yzXPJ2DI7eoCfMMoP30rqeTjMZYBE19Vj8s69tchFBtZX2BV9Y8DEtdscrBXjmw
DW0Og0oA8wga/McsZWNPJceuLgIAnHyZABs5YyCanHUfS4NVaPuDGln3WNcIbnuo2P/tFPqLbNra
aA2lns4A3cUamb005eOrFp2C5OKSoCsJsW+0p5Cz0qohWNY3ffPqBGJRNXW5yTg/iEwhqFwD1ezG
wdFtXmxJDMPnmE5tUaBD5N9jx+jZ38WRzu/Aj5CjPVhZYZY5LniaQgg62jlWkMyvuyyE/Uajk3BI
yILen96jqkwUfHcpRCWZQR8l1VoQLJ+/DK0GKgxlF4V91eG504u5hkjKCJLSTjLai8u8RwFv0MWF
1bbDIgOCRqn8+g75R6cXRyhgp1o2Z5bpJAZ1m5SLBC3Sa5uYpjoc0H1ehe66cstbvtIAjgCGrfmi
tQkeKzk8WUTfOX6/u5bs8KMHWvpv4RZqkAxQQkG/Vkcw3QaZktGL8x4nPzLlc8bPS1E2o3udKuXx
svU3Ay1ZirATZpAQQA5qn5VZLVRJOWLO88gVMjK8207p5ncJBzhXiZlzR5lGNAlTDcN92uIx3Vyt
W0IErUHiHHQ7sYjyQvrEY/3rpiBl66TLa/3W6C7P1Jam0Edy2RDab93uYEHqMVi5FGfkNNGHLufp
oFqdC/fkM4VVFnVPgN9z08G8G1aWWwUOLocesjdpj/ifGtmlOCM8udkugTD5k07o8kF9d43XTxch
EEZG/Tnz0B/lpnZh9hp/D9aqYCQDSniIUeXMwveXbFRyuU3oSVxHb9F7PG8NLNI1VXQduTQuZSXG
k0B6f44Q8qYWsajPQb/SDnwxB2cfhSodUGeiX72EOsGYgUiTf4/OYVReqwL4u9VjlDSiaPX/hH/Y
a2tZ4gp53tchJqgk90QeSA1F5cQ7TP+hh3lPiMMy9sJPVbnHS7n4edFeJcBpage5K+4Q0FhEoVvB
i2vWp07Gqw+CPaifbrMxk6N65wAk8WEQvBW4Lwb1o60VgRK/JiWS/vLZ+apwF02P3tSeGYsykoVr
h7/AxAMnB7DroDDmdWOzVBniSMJC+8FobdPCVGt+OHTwX175kOW25IuLz6roX7M+9KcBpbEcYGx9
nhRuY8IX6Oq0714/140w1DBp9qf2VfAG8qjXixpeZrZTKwFJgJlFTDK6wzK5oSRAzLWhQBf64Xbh
AdGXsC76gBXG668K2rmjxddefXNAOD16WE8XnrzyOA9ookyZQHfWnt0vvOE6yCIjOC5IIr7pRgFO
1++cd+RXaqu+q/K8xEnZmCc8Sa1x5r7IjW4Wpnb12eY9pI5ATduNImCM9l4DICgsVl78LhdSQsSK
BVopEzNY61bKO1gqoK+8wDD2Uk5kEKOC9g6HMA2oy9nHTb1g48Krdr5o+9gkyEraudtemSM0eigu
8dg2lUd+gEkfqwbRMGu29ghhAHyogYbhFacVk3vcL+Yq/PCXJDSj3upOozt3SmaE/NHHakiZwYOe
Kt4ax3nz1OKW5HrHvg8kP6B26cHk010mh6/Jctu9aK+YORhfrf9MP4IzVg3UQC2s0zSqzJVlZFj4
P0eum0VNHpiD3qBh60Utk6RR3/jrmzG2NBe5lyscdfHRO33nwoB5OVDVodpVTdqIc2I8NkwKMNKT
/dsyffVKDghS6OegU3Ig9/1urZmSRdFB+L/qL2JEWbX2sQ6IjGflq0ehgjYz+0uKAHtexY9C6QSC
rZF2lNGnUfYxyridQgDNwcY6/BwBOqhNyGr8iOIKG5ugPGdHFw7hK9GoChJGzr0JQH1nArkEa6p2
w3Nt5Umh741AD8aRROStJvSw3N0W4jW2j0W3N8pTZyZivmc7otlQgN0SYK2WvvqBluTqff5u4J1+
+ZN50TTyGwckaGgB8CFQ0hvj4edy10wf9h1JntMiu+ArqaOfSSRZudo1jpCOl8UW3GCrVIvBS317
9rS1+dLFdqnMEBKzrA42W/d7d5TApQr8UvRiY8ptqsyPvmEPch0RFrxdptTlSV8fmUSLaQon2iKp
ZyiCylGt1myZIMQBUMG36pmtB7ibxQDIYHrbWj/Rn3DOy43C7UgNpsFlqf6kwc/WmGTaMbAO74kQ
fnB1A0HSmeM0rlA53lNiGhcsbk8PQn9aYIjBQ1nDNTY9YDXmGsDMqr8xL7gi7H0uFk5sNxruoWbJ
qbim3elZS2rDWNNdSstRrVRse7uv7HG2sDl1U29KzdQpiluaMTW9FrqtBYW9/HbewLSsg204NC4s
8jrhf/m8gk+vOzgpPOyarsGSwhb7AMYhvRriZZSx2zRtAsjc0d+3pHUzz5GdxhP/NBkZJhvuHdxv
UTNGwYg84dM4wlOWua7xkddu+WGktq0BsF7Wan7H/Fo+E57UAHWg/esy9OygOXHtkRRyUGOXstX3
ay/AIGB01FM+KwxD4oPU0iJaA7bja6PhYHSaXoDoyh3UDY1tMtA/wQhi3WO9u2EecjGt6uGwsulo
oAPK2lIIEMkkz6ScivQOhhykniqIpgidAx39ylopwWLVlftygBRzIRsyNcgKDmj4y2wuwBH9jX0a
e7muOtR/dqlx8nX3ngaGaa8fBtZs2AB+T7p5+02NtWt4DHNBSTOI/frZdELuS3XASSGNEfg5HcRw
H1Rn/bfSK0rnzE6X1VBKIXBbWw7zuFHUTRdViiqewwkdFATJQ6dNQzNURIF/jFpODkWRAllcl+b0
xWPmxFnCwQEJ4oSbdiARatXHj3MxWdONTQIPoEQggrvo9dKAqVXnjGzLYd9k35ZeciRgQr1EmBuT
2Jzxz8nJcZRTaGC1mujJYSLmjD5Uvy7a8YKm1JPxUJlgsG0SwSDBtUY2hPZ+gZPHDShRynWo6Is9
za368ZbD8zDvzEEhPH03nAoL60FZIMQ+HdY/l+9gUfyvdmgc7FrmSVX3KRZ75ufPqiw5LauuvDlF
8SiB1LLUGac659uQ1dLXxmPifSWSumJeRNz2srwUmNpyi3CSnnTPbPQC6DOz/VZxc7MIGFNhbKA3
ObhgGZuWqLoHv2+xRvXeh3toDwoHVRUfCNIajuM2hxW8Hpu4Av9f4A4wrGvkVqvGYLwXyu1iqjjj
u8WboE8V7jTYX1pVISkX7U3aXlg99wabujgpeRxC4EVJSs3TUVpsUOHY+KUot65vMkSS3dnUI/KD
RKyE3WJ5h21kM8o1Sz3X3YmujPPHCKX23opxJjcBanCq0lj2355KZcGFGX6umfUtpS+kueFW1gVZ
h9K+KK4PmkkLIi2AXfImTtlS9nHsFmxpPbAphNhvpmJ/XPrRDcOIzxL8T7ER0EZj6n3u92IJk64h
qqNtgnwoWEismnFYKLjuX8cUM8spBAipmCTB9g4xbtdul2mF67JNPvwmcGsjr/SR/3Z9f2vHsVTW
y8JTaqdXlZ6N7mZ0mHZRR+96xKwCs9pHZe2ZK/W7yRAyGbh7xvTMSK1lmQt2ByB5chH1zoyRTsdj
oxMV2LiDLfIz3YkZKT/YKebk5z5XA/wdTZV1uWLsII67ALdx0diWBBaFDN21HD+ERzWm8AYU2dx0
bZzkArk+b4TsYiQZFC7rOmaSh54HDX6rd1dSANU5/cL91yFFCxTkdPJ9xQ0D6jKRx4GwFt/KU2bG
nttrO+vD4noCmNpASdq7hd/g7HoNY7P0JzT/R06es88SFDb737YcP/2ZjQSC/Xv+zSzyHZetK4WV
5N5gS8ZscMqIagGgmcddsb3XgVjqzLw6NjDXKEmcCKubEcpz1Pp55wKdk401khqbVdJ5n1ndkDNE
z/f2bpc68109hoJKCS7HHPi66oWUpdP/fovx+6HtI3rRHEK4c9N6K9IMT+UUqxwEyzVdjCADlC8l
0Rb1EtQLGw4KFpH8A/3aqRKjHxbmjA/T++VJsp13JQD7O2O6IdnZRS9bbGPI9zWwC8EfmhiTi3pp
Ie4aPRXTbmDsCkkNYtMeAcycThEaL+Svj3Vh0hRBztwEKxppVawyOUFKahNziVGz/4SsCfBDEiEe
hCcttU6x/kn55RDIwd5o86It1fAKOObaxRUbedZFyZj6tcyhYhsJR0III4/a3rbNi0FXUEldicov
mE23w9ZrruBbZO4C/kjtiCE4Hg/jIND1gSVlLIoswlEF5fQyU9r9H2iC7yffCECTL3gvpxUBrBFu
9oQQceThDZHOfuKDuA1LrYDcmU1SN4kf23RTmTRQfdUOBgJbneAEbHoocBHD3t6A/v7QZnL5c8Jb
jjVQO1uV5cfc5aI3/+n2J9ayN2LVUUQh399xsH8dhWyRDKBCVkuLewEBpSKMhTa0B1/0/HkofQqY
jwqElR1Qmmt5lTgt4STCe7nuAqmK/PVN8vJ2FHbRI3vE1I0k0hKSHczWNWx+rmrfpQevE75Bej+h
QwCzW2OdItnRH091M70fCi0UQJWRnMzhnnChNaiu+NyIdxL8xFzKZli4CNDgr+7bBEny+g4Z+iG1
vcR6R1UcULzZe9BEESTStvwxvXdj5UqaMcPZH1nMJZ0IwItm63yfeMHFigc/U8XAja6MD4R08FyL
knTZ/cRFA8wisa/AP3vY6p+CFYEVwoXpj+wdvqWE+GcmhduFN8AVWCpLC41VZ9Sm7WJkPn7/77uD
XT0AEqKHj7yWoE9PBIvjXuCZttdq3LABlUjCP7DVJOP3yo14I4ng8ELNIxi4JcdeKbjuBfeBXo4A
C1dcMAs/5UM+k8Fpj1zlXIORPvlU5/NOvJFrjbIKBAiG4+b7WthsoDlamBRdqyfSTbMPyrC3HWvx
obcg0OdNtXDl3PC5xj5RefSiJ86q2LveyANpQYyvUwIulZSh8buOkPe64YgOro2yDaQ/2M1DYdHG
yA787GYYS0Q/Jtf0PJZiD/BfruLjTXQzL76GuIvus/TSV4gQMa0a+Foz69Fk9HHEqFPV3HqWOMbV
BmQSgM88bl5FTmo74CJ0BV3Ye/x1CqpCxGtSCMjJG7T8RN2PQ3IjBsaf612BFjK3agCVIfk1DLLN
mjK9xEYtAjXNW4I3uGVH88lZutE3RnuuVIEGUCdmUj9z4Wbzh65jku3HMyacPo+LTG6rRrhhbohX
xVryt2+QjMdrHaBuGDyk1lLXLfE0pw9wn3RBb8EP7csQ9QOsCSTbQ+JcIb+R4YU9DyUabO5xL8nx
O1w/QAsrB5ZoWVCHfO0ORc751Kg3fGkHwm+PtPCIg4lg+rcxmb2osiflxygays4iGHTsQtnOCfs5
4TmyuKtrTUXiwdfV7roeXA71B1I6QSyDpjRsUbBcgowK92RzQGqQ1vkL7mJie3xCpFaMf7Gqw7+P
8wpHV8cRchkBbCp8Q62gmqj06Q7lHhI1U636UICfD1opaZDTjmYnEbC5rcYj9FZPbOPJSyzkFKdP
QQQr9otMgszRUpRzRD04DVJ0g1oQ3BBQY7ooxrMoEQr5mvEAyQGzU++e9KNNPH6RfICnT1+G4Kx4
k1mA4a1Z1fPm4JHcy2Noc9uPOF63dKNmE9UiQ+AmD9aBCwtR/OtlC41o/OQv8Hb7KCDCCKGWruLq
0OOTqjfjvncOBpuT4zAxGGCRaUZUE7Elowaon+5W6I2tuuRry5FtdvbwJjCDIwgL/qDyv3UZhRTm
RJNk3kBw6HsDgCSyGJnr4+8ciGuCKwjsdr0asnzYWeXJ7Nhwh/iM/cnDWyCskw61lCdQw4xqVXuk
dcLSXuD2bFKSxKPo8fpHlvO94fhgOSMhl7nrv0FhqeN20bBG/sANmA6pc0REQj+qdh95Pxd6FHt3
zpJ4xY587/VgdHVTZGoXsk0tOFbixioK1rBdk3gSQCK3OC+3pNrOYxscl45xAxM99F9egMW9rFdE
XrKFJkAQfMLBJXUMNTaPI0QPLM7aIabrLYSPvlQkYnEPR4WjyId1j+xySwz7+Wb0e6urVn/kaLSS
/v88wO4uLYm/M8ol0PR7mkICdfMNO9AjcipNqPjSS1C2Jvgtya16EcxG6zEOK72BFMpSSLugowng
Tw00dENObA6aXRF6tOo6uuEeQosRkVArgvQL6sx45GuWYJYn4pBnbOVtV75oEqC6n/QWJZjGq2cW
sJx5STm9rVqgzgxbrP/edmYKhxIB6/6w3ft6kZ8q9iuLjti4InBHhtwQOFBQOfJQM72NZ/pbP/VZ
5+ImHKLE95z0xXMacljZ3ORmSkRYALjXxNzJZY/wNBR1jZNuIV/NavgxjfGGvBbroaRUxHs7mr9v
mXLvpy+QHjRiYwTucU3J66e+RiZuokFqNOTdEyl26etjXJdmc54Qv0l7fBi+Wv6mB4iMEoGSDaHa
miumtln6X00f4DsKXclEo2O2DtTJtxD6XOyniiuR6DEswtcmRI0ML3GXw+BlG5kLS97nl/mjHgYg
TF7NIPLUibrxEeYPOJ1KPfQLQ6DrTUdtr3wAYfwOyaj2q546aH99GFkt0EIvQwI7hz4p7yrPBKFP
dLDNnwhmWFn6R3sWvavNJ9xU2whO9jSDTK2g+KMKOpPpFq/M3N6HXnbiXXUH+ZeHCh35dV0lIZme
vDFakEA0KGjC/h0ixBWMeFhxuXArTh8wZBMjyHMeVnHvix6GAYso7F1Uulyy79XMfxdSrzRtTNsW
O1CI7m/hCKkfwjv8Wbs0NckCiCBcTZeerAHmelABMlERt8BoW6GebKYOeL4gd8YQkQAWQ63SKDKu
de/XRqZtyf56B9zfMJwU+Y23APOOyqNDoBg8NM/G8bvFQpJchjj1AlFJYrIS1KSPIaRu0iyLVfwq
r0UEw68DT4PrXFFUpKk2bFkofCn4iT2vaFLemTYb3orJEAiWqNtrCRsChkQfNkEK7LYHfxia9UE3
HhblzwJNcrWuMKNpWa/KNZ2e+Bu+pNCg5QLurabkqys0OtqV9y0b24G1fGZpAJsmBXHbDFr+G1t1
bCG9YrqvKDYSFYDxP93qqV86HEPbo8t8LCxJu9lMEGnaq+Nll8pr+7PccOi7EX41TFIeyYoTDZNd
vRinOZ5hIGOwJdKvNvBXPZZmaUd7dBl91TJIpms+23YyvNU1WsEYHAX2KeNOtBi6IOOCpDmL37E6
z4eRDtrD6LekKOuGtce6lVHpK/wXnNYO8YcnpRCpjqrplHoZHe6LfXGsiKpMr+cxZZ4CUHY/aIle
wrUFwAsqZgQPzOTt0fkYYcb564hggH+IuiJCZJrFbDsWdlM9NrsmwPBTVhv6HBJD7cIzqV94NXxS
tfQM83dD7D+cN0zUGbrhIhv2uQ7vfnlJjIXXFQAEOTQNbs8+9L8j6hY+Vr/MCNQroc2E9/WNKy9r
6mcfPnuIhYZSe8xL5jvNHff+R8A5WUPKxES2UrsbCaaBXsbQo0I34JpgcTAQdjrS/x11n22wD8fq
GtPPkjrSuUipmDdErj09kIkuFwtxy8fv1zDtm4dJL8Bm03nQHzn4xqoI8dfwYkUjg3VmPDMPvhQa
9dfjmfV5SPXpCrtZEDwZkHlmN4EtfVo4nzkH27brvNz5WU+PF2OaDAM/Q6c6ApNv2ckGdD0NQUeU
K6P2+x4UrIwIWMDv44gHc8g02HfNp+cTpe/2PM5zwGZqiuj1Is9ck+XfZdHg6NwXVjiA/Dge3ifn
PgeDpKb2PT2uXKOJBEMushnYaRYsnHXowtdVM7l/3MgS9nLUZlLKwlKzTh7XG0JheLaKPXnlHe2I
NzlsHp6GWEpemmPis+HkECLm8bdKA+zdnX45RaS+nRAlygGqXhuv1U3UgLb7WtWQVM2JNw++ceni
Xoi7heD9XHuobyn5FJKvyrEcz+YQhv7n3s4AROlyDyZ0LGGeqEoKsDHe9RzSYXBl+7bdw4WED3e8
6Wkkt7xIHHvOZvzYXDmIID+PpXix76DhqXuHsuhrllMDCi+d6+Zt1/77klRaGVblDfvPCrL/HOxA
hmrr0/LtxERRO+OQyLI01N7qx9e5ZZWsjUpCESx7og9ybL0FrAVnbO6A2Bv1IaQzZWQcIrujk7Xq
gVh71YcSQogma32RO0iXQw0p7v5UsGhclcoz/Lm+tIv26KFp7XRO+NAZ8f1HwNUCxkSX6Awyclsx
3J8/RzsGb9VkKDa+sZYlhwYDkfNgUqJICRpXsCH9zzjBb2k2Vie2RcqDrbFp0WyqxvvXHrGTWB2X
nqvahomeet5tFQ6XmdQ05pUYFgWXAWuk6kCOgA2Y4HyV8C/EhVYJKMACl2hmzqdcJlOUm8BUvAXI
P5fTlNtiai+v1HbC/8TovzAAWErSwWFE5ZrpJEg/Am1Scsf3WU9hEK82rjYHyERMQqcWr8/zz6KK
AFQvbKO4nEFAR/ccOuCIsv1zdP1TNoR7mFn28UTBZyvTcXD7WVwqgMGr7rqazZiZ6+wmEb61QkIc
t+wpd8E2qG3Ks1g0iW0Ma8oSYTM0gE27HkCNCvfw35g122PdECKx8OWgYyACXIEPPB0CUyzYJJoJ
H4H2TOwq5pR0P3Z4C76mpG7VAjQe32w/mVc0aB2C+qfnxgtWQ0g4jLJ0U8o75rFoXdzIRJ/JjjuZ
66iu/f66lnRE2SQMMEiDPd9ODPRdWoRXbHhyX4dLd2n7iz5S2SU3zgyD+XGmuUJL8t7tGbAjbSnR
8+z0aA5oN/v5qYqdOiy/E8A8jXQbcxQmSaWUJHFGr4l6ErqefXIl+nEAvYtE+A29IFIipNKCbZ9V
LSFoqTtnR0YY1oVMKwk2UH0ThqvX18YSjlZjMxWJ7Ew4+ViAn7ZXfJ1FuteM3Pl1XMTfh1SYsXeV
aQocmm7ZYaPW6U8PdgDkeTkn9xggWBesS/e6na5qEQ6usTw+2VMkBt35wJ5AZgf4n7ZUVxSas5dc
nT1K5nG5NBnWXDZq9VUEFlLsfRnQDtwnYu1jR6c91jwjSmvWN48N+Yc/bke40knIoK1PKJUmijvJ
y8wfx0oAZrLN3F4Ja2RYJvCy6RPX633GGwCpO6Mo6RgQ67q7umgWk6Lwz8wWTaXqeZTljP23sH9j
9MdJfDqUr04DCVgG+S7wr1SzPWaOuZxk5RJgJc342oZa7/8sG4nUF7T1bZdkdrNIX6aNXSjkvFOw
YneXjplxAFwmpHrDCLzLaVwOmW6rkKHp2K3KXoy+VZ2tR+g67ZdrEzL+ovu6fkICg2ek/s8US3kb
lEUV8lFk30YpdDX2cnFwgbZwFo2UW72KgQqm7impQ6/3celD/mQEKmqPrvy+wGwgX1fKtV+s4d1I
lwkUNnMeIS9aqqsbqTcf5oW+hOgDUJXqGPoLOLrEafSnDza1hS5HklFMUv3Lruo4WT9oB1oB1KvZ
ZsXWsQPpVqPrW4RFEcXVBzibnM/E+0bo/vjcRl2lPYqcVagJTEgWKPAoaX4CWxkLAYDfUAyrGkfd
YDOqzko/C3Ss8/o3DBOhaeSZu8ctfM2J1EeAWKaihFpXXoaAM3p6FQtwLk+anH7d6+5OCyF1/nEa
SGiH9C6axNXC5o9BnRMxlIBFUvFH1Jv+fspJ0J9RZLjI26at88GnL15osT517jF2TJUEUbhMtKA0
hSlRn4eCGwQ5FtfuvwDFnDC5zRTvBLBfZg9seWFxNQq8dUkcolUrxnbpEkh+5oQJVR9KJboy+QQn
9F1NmIgFfckIIU/qcQPw8IgIiXEE4lIPVusl8WWgGrLCjxZeAccxhC/GLWTAPcRSgZMIVuc4Mb/4
k/thoBgx3JD/ylF1pcblZ20O5BeVeEwl7ZAQjYJnL6p4VGgblZhha4pRfcD34Tmo8ng+zeqwNJ0v
NDeEUbvFr65cXgvEeAneejxI3AXB29EywTBQFbFcYgCic8ALgMvvKxrouc7RhqfDztJTrSgt5zua
bVIwdQV8cqfz7fap7ECqXYd3IfV/s0lBzW4asSz/Iy8HM5A1STVoNQ2njv9+3B2Iu55zg/hS0l0P
G4SGNS2U6kVrhnzJyBLeruah6axwQpk4Yv+lCfKFHyxKjMuaKPzeul9uSrRJZCkK0j32UFVHXfcD
enw0YDpjMiiZMEY80Niy0wq2sJJOQKgCGBZzAVMNBG1BTUcXqfRaivOLwzqXUosdpRSNc3VeGbXs
FMnU5zM2RE8f8z0HoMoXTW1VIzDDFg8cSaV7p+8xbWmhhdMy5tvGAZdwx45y/MB+cg5mgWdDSzWm
XC7KRofpFeLCsT4bu6Yk1d0I3Fa2zEWaYBHU89xK6o8+SUcZlIqIYYfHB4W8bz+/yl4XC5PL1DSE
idyR6rdmqswIZi+wOatBtX500PemMrNq2n0F3AEZo4VukUz3wf2byjlzTj2knCwlT6StMLja4q6I
io6E1bemJgHJJ2MM8qE73EU2izperrVHImW3XlEjsEzF8MMJm7WT1bD/0Ip9ErYE440bgpq+2455
c0/gJlD1Z8FIJO043/t2gvhRiAifr/5fhQglGB5ODjLVsJZKeyHeky7LQgnjmZJjBeBZOG7Deiay
C92moCT89r1wj1TLncMOVtPQBOZjCNvzIPl/UovBXWzBLAltrWre3iXs6HGZvoDDqMpMEA/AqzJ7
lPOlVMuhAqk4gcPbIlKrSoSkJ3zcN4i3yGLj+9oRg7EQwN/iKKInA2PF9xfWSlKMi0rPeHJuvv4i
LLp2/DGt70+L/w03IEDwjvv6PKUatjQsK+GSi6qGXdliSJ9sImKGSDR4UkG/nchOB1YZ0CQNdNbJ
DTXdFjB9BF92BsDNRmDPzdTlEorc+2OMBMX/L+VFKvKrzcGTw+HHoUECAVQdaj84wQbP++cbYTLE
URnWhp7KbRHHKXmXmMGHmDdwLTzn+I9+P5bFOPLNbbLdgI4FHdCQyttRKokM/CEmlvBD1jxmNwB/
k86gtU+Dnmg5hlI7sb8LaTJmCI+ihMoBMggWmZCch+/PObs00CunKv+rlcn5VgaDIqvX+AKQ2epX
Oz/FhW8lNYF06D/Xo7nYMYHoI7m+4x6fTTOw4hBw78EPeFPRy8Kt7U6DLVTmHfh09CLyp6kUxqhl
zemdnduG6cAaPGqq1CcfbUjum6vpl6mo8gV38Kfa4goyoAv72OOdAkQApvxYuOMlBfZY9HDUrs/R
Nnyzygn0uK05jFfXcLHkIQe2K6AAcLLQVrBfUPE7lGMYumkMPKF3yUESduFheYlHVZAYyqOsR1uJ
YqZjjG5fMxgOo1U3JLPQr+bOV5IoJsx4TKZHt1710MtWKzr4gJ12Js7eINSWYqjvcIKIUADk2+mA
J5axOxYyWfDGPRV/xTovNYt3+2MtaQsENr2oIzq2dtdftqB6PAQsns3DcgUa3PZsugd+IbNrj54M
1yyHSAgGJ7gAtC85o90oA6e/nT9OZ1c+fJ31hqD7vUFeXyH1TacQHbZTRGZiQP2R/kIfnW0F1b7L
Wb8dxLXtUhHimdiCHn9h/M+6GOyLv5ue2ta2SzzNPOvt3Js5mMvm3oYRnPiegcjSr3Wu+RoEY+BB
j4tbo3Sx9K713sCkx1nVzUS5ZoDQpZB0c+KenPrnqzlr5wfrGyNqc4JYRMbkeupSP9reNejuoCgM
IkDos5FCdv+CFA6XqIkGy8bukUbfD6CkMqpIoHRoquabTKe+MMDMloRl4wd6qksaDxfVrk/CVCMq
4HiYmgXJZ+a/YFUwZ37rp20USHjfhtlKQie5wpFtvZkSCPdUdKo24BYMhpdxu96aZ8A26vVHp6s1
4p+LyKDkNI9+slQgM+x2x8bJUfVH342mQ4JwL6+87GqPOI4DIih3jFBWYimNuRQ0l7CJc8CO4E6p
qP1G9sJAd8XyGPytvIQsDAVojYIiNH1OnGAHRAKNkQ7rP0NjG3K5d4SQGyA/W2YN8LtM5792FSgm
9l8KIkcjxBssE7qRs+q/cWJUyUfpO4XqowTANoR86+xQhkUC8viJ+s1Zq6T6oRplLZLgo0BwM5lG
ZF60h54DPltgrtBE+ejP9zJu+cR3bv2odr73Xu9bhgJVum+x//u3HfcCHg8rspQ1ZGU36qSK9QmQ
667ZR3XKYLAnUJdIe6cPMdDAlnlSKD8HEOppU+gr6OBOvS+oljBC5LlD7y3CqryO3oc9QDNageFK
GZvlBP/+CgPUjEbJkv0W/hTol5+bpM1O7AI0rpYN4wceWK2TJ3PoXuq8B8HPqbxq78biFGzuawfS
yQs8RtHEYnG93vWn5368qFu+RyaaeZQP5wDvulOgAjUeJ0TK0NAYXja+1ZK+fUeMnY4cfVAwydRD
3zzXa1Eepwy1jWQpgYvfuA3TmL2007DzHUg7JcIzRk54QF9XUzkhou3m2ga2btgYtEJclFodGp/c
kmYbxfB0hYu5SWwl/QC1/5aInuXn6PfCHp4bNrBZmlk9j4Kfd5klZ86SBkDNPZWgns9PtuiNctGv
FR6TM6Zf0VNzMSFHLzAEXcXaGvu8qVZl+WX+f1buBFmewPnlSiS+KzuaGM2N1JbituYEjVTy/d4L
QQCNq1mEFHjGUOOFTUwmmgWwmal6NoMs9gs8drd+Y7AJzaFjzZS9O7Xgb0m49tWKfEUpgxJFmWlg
5PiN79EcYiSnlQTie6E38hEzOtp1iQu0uZa5Nar2FJ0zV+s5vfWCM4Bc1Lbql1M5Xzke1HrqWlx7
808iT0jUP9lFkI7h/xX8ZC7qjaLAQQWCupfPfhR9hRhaNd4JavZPQkYVL22PYhP/cXngljX40R+C
V2iY/1kfZqr95tejlhl2UVPhCj8d32CFgeKYapTyp48jwK2B6d3dIZHAVIhMWjTwPbGduieV3jue
dTtxX79zRhcIt2Fev7WVJm2h0ynowNeYXh6c4qxBWRJDgnAbSoCcxzLxtdEBUNibCVo1gimeWH/O
gl6Xu/aydr2Zos9ua9L/a6y4cgbC6+gIIjxeD7PrSgF3j8pgdGqVQvLZM4Ygi1+6+Ayf09Sl7yUX
1BvyMM8OPkeieHkmTmHRMbu6w6xDs4D48Ur6lzrmCqhJjqQ0VgpKh8zWF+SVHswA+FQRXXF32uDb
f1qcD9avSFXTL09y3SFp7SOt3IbvTdsemaO/ayGhtq9slMNgdEnlpy03rzFgMSAyOpoYuLhsd2+f
U2771aSaJl+0YWN5zbmh4ktp99fKrn02gPqMawUHB9S25nE/vUqWKVpUTdDt1ofEewnmd0OAh4AS
x5p1dUR4toIj8FONoPB8spBYFM0M0lihGlPBb91/ROAoGH3Q4Db8l8zh0avkYoaAX6ZkMb72mWpp
+Lvg9gsnJA7vb+mihjGah9Fm61z9ycNBUym9vT87EDBYbZmQ2oW48fELlCPOSjolw245ULpM8Ojw
OdvN4/OvMaZjLdov2babUkHHHyJqL8lAMmQgbe21G0xwE9esBQqm+XNRh/NHoKF1fuSxGdDaxaEg
zGi9jJpZCmvzybGRkrWykpVYuvOZJUUupp1GIt0R2Z8d5fbyKJ5E0x2mNnqmEaHLOstiMgxGgybL
SuqfE0j0ccAjkIEal6TdiAvOkGTJNbDJnrLe/pwBrKBj+EIkSiNr3rYwNFke4YzTfbw3C+8TgHKx
99aA4k5Cr+kIg0M+7L4n8QzLuZ8hSPTvEw6RGrW2Qepb1CDKeTu3GBdoRdjwQPqYbx36I2yh5rcv
BdJgjuFRcXEe7q3BAW9IovVbWSUaZeVru2Ey6+c8jM41+vPS6MdPzcWQFqiTN7dTa8MqBmGBX3IQ
3EnKMKP9N9/1AGkNmD33hh2Uh6IuCRVfLFlJqciGo+4WjbZE4x3jG+H+BVPqepIWX0HYpE0FSKvk
uQTyq+7UO2tfY5k3cI0+0gtBl+u7EfyeVQt9AcOCsSEDT9wloTHoe1MV92lxVk68ojG5nwsTbEO6
OBNzEaLONb/Ob1Hmf2x7o4FYvCTQdnawNCi+s4GYvg5OXuwbD1zWcBGNvkiTwUvNu+AdmC12FSkv
tVryGgS5LBdSSksNCjp6RKsY+Ln5DdVB7eueoDdI/mMsTZdRm30Tsn/1Oqp7g86/b5bcevVfjDmA
7l3GJ7LCA5evcDmrMqO5Y62g0mpCneZNk9J/hd7glZ9dxhTEwMrJYWtsklBB+X0IjGK31GX8GT8E
vB+i4442HZNnWP85z68zFQ50KkcmC0mFcRh+G5D9pCLiZnIIY93yfNA9eeWFMI/iy1jyPRLZeecD
adQUfqSSzqOdbdxGkEbMjAey9+/flRzTu4uNo2l6NeIvjOLs2FxGWD2F1IL3vIDCdJJC7rPYy5K4
maN1b8cCwE5auAYMo/s7azQVaTPYTlusRD2jYPw1Qjjky+rW2/0ZcE2UaZOM069kFlNtH1a5UENt
9re9gfET1V9wzENgMswz5GvH0p2AsfE/vhKfulYqZB9UQ1XDfW9r/RtVWhHQvlOGbXya+fvJ9QRo
hcPLaubsIzIPORNk6pbFgJzt8fKH+unR7rL+cvgRoPNjmFwBrUuba46M+FcWMQxVeK7ATU3fYo/8
6lkcy8QSnMSl4Ws/fHsm4LjzS+59o7bjUKfOnaKvMgkKa2ibOSQ/Q6vWcGStL5IlnHyTH899IX5V
Q5izOg9mnh6vHCG69GoyO7Lwp+LjWhqu8A1Jv1Rf9Nb9KLTEIe56v9EQreHg8o+W3ISpCMySNe+0
SwQr99znc2fAWtnv//kDMpux7sYxSiAXoqZH0YbcVC3K+UKWgnwuFaSSW2vwQQawuUmAzheKyxx8
nAxn4JweUR52ALE6MBQbMZULOXeFSMHX59kDcJWo6cZX07TBtJ099TLz6SKdcNYRmoKa9djEczVK
5vwNidJIyUj2RyRzRrrHJh3cmiPJbLWxwfFt5tpGQ5EHDGraa3+6NQtsF608I/IFT9aA0LwiBmzM
UMemOyVe6dibA8265NVsNAN+Xvx6T15+ipd0izgPP3r/nE2d2jpS5sA497QlivhtY4cn5kiGbe9W
9a8F6j/JMsCsh9L1b3H+uw3+nwVHW6tSVTXvrtxraKIaVrbgjiTytjLDuMir/8kD8Sw9puKM30QO
zpoPHepOQpQh4C/un8r/1p/KHm/TN0vOFoc5AucpeypVHO8GiDUgBW4g5CMeohCIhJggRw+AhFKd
P55lOoCNwMnA033WzRSZPtVR+c3xkSyYI1Oh1O8zlhhuEYGd6hxLDULfh56wwfn/wZLps/uZpZyO
E1UxOC8oH0N4wfoaV4GnIR1g6WahQf+TG6j2219q/no0xF84xa5uijmh6p0bGy46EO+oQjjGZgK7
CkNBh96sKerHBgAMQKkvx4NTUD/rYFtydM0tEwhZcPM0BI8toVWq0VjN+kxJH1HZ552Vvi8yCz5P
2PDZqR1dFxX1ASeNoDHTzEZFPE58JJPZUQ7pmygSoxOTuidBT0sPfZrqfHZKsGMTTbJIhYaoZCyg
jKVc4A0k+B7ogFeAjZKvE5BXw6+EjFgsUOxjv2GKbBe8YWPB8wH5LLHu9GxhRaxJh/4mpBI+W86Z
ZQt7uLbB2S9eMrkaT/xBiW9c8GzQduc8n0mucuZl1kOmdBTVJqPOxola55RHZifmsZ9LzMf/phLc
4Ck+baNi/WfrYK3kahiisyDAqbWgf+hN0498HWOukkS9l/LPpTsUsM7GhumOvFf+W0BaNBk2SDM+
cwPYZwgNuYF3mzo0+mIpsXtZMj3fji68st2zlxEkSDsmY5AdCcKfylMwT3Sd+KQNb1KGMftw42LG
dTSSK8XM+tuBoArisW9DxcalWXujuoKk/sOGSzbXmMVlutiXXG471jqGD+ayo5uxbeHFHIviyTCb
BzmAVsFQRegFOPET5/WcOJihEAvpwm02GUAnufy6wbyFcmo0Llb8OVCILYvSsttUMDxYvqUX1//O
8CtZ6ymfBCgLIlP8CMzXn3y/LZnVjWRzLODn8Ubtw2HVJkjfXO5X6kmf9PLEqUaRlwqj76BzJdye
9YeB2fH+k7NRKFWCMNwQAq1zxbcps4+yiSb6vCV9VDWQS67F9HgOgzOFriqFUlM5mDA+U6K1QQzE
9FlmvMp1MvBuGJvzzogDQd31WJkHeHlySRtqcHXgGG5OSnlxfXpMUW/wS816CsjCmayVXez2ujV/
pMcAR4UAKe6m6qTCqts5lE6YqKQc0iDIu7VMzMXI8Hl4dVDNZ0HV4bGXXpKhzLx47cNUyefdUUrB
xJleiiEF7MAfcCQ1SMwL6k/qtJ9jgHQYsCfBUaYA/WYlHp5WD9FHQdC+omwe4ShZy4vVjFEALZUS
Dlc3NoLEP8mErOCChzSirfGi3CT0n8HOREMaqe9mf3upgLuxo8+RYGW2zmCiFf/H7sSwHLs5aV1t
/60bjDf0jDBpOMDBHAj/Zl4uismfg0q86/wGbGn+5A4xKFqzaBrzx1v/r/RrJqIJkKzZwVBiSKu3
bKIqlhpyKaU9tsU2whsgD2v3znT9lZtKjlysv3CO4SK02rb72m4w7JhuU8JzNGEkRwHK+h3xWnzO
2BYMuSKPiw+X8uyhcCH+HAiVUrR32NdsI7tGY0UtwKT/OxW6gJ6WwyVsERd/otrRujKs3VWR61Uc
4Oy0CRj+dIdxD8MRQGbtNEQ57ThcbxDwS8WRE7r7WvjS+JlgxjC5oYKDhiwozSFRZOhUlmU7RgFQ
a1WTyR1mNUw70jUy2PAnLmjqyBwTH9nR762uu6vcFa2IiOwOnvrcisSMlrLo74vZJMpA+KTSr3fq
uyBWnMAgXZwCeG8xFDZmovfCEaOORSfwLxRsGaUZlxvLibcRf29cTXA4HCJdgQ514eK3Yb8mWKBT
dQTBb7c4bCboOeKtlyQtXbVzQfXXYRW9kzhhnNUoBUFQ/2Y3JDwr6SQ6XiwJ1iD4Ege702ybGBLk
QSycP9uh8tBITsYFDqsPuHiaOVZmfDz+eAYY7fzKYK43V+LbFIRX7RXWr7Sgg+t+curiV5yvO8DZ
O1MeFsU8Jw2qthvNv8ZhjBWTP/EtXr4m3TROdaXmLXCk+VVlvszv9PyxPH2t/ZVfkZkeyglTQmOk
ki11JkWs+nyc2nED2A4hPkQk1wPUxflpQ07Mi3uQUwdbicamFbei7PR6pgbkl5PRdhWddoiFOBpF
1MHPjE3ic5xG8zgwm1AtQz7A0ZkFw/WxQ/8Vxi2kmT4Z5k/gSt6w8CeS+RNXEuMP+qYIawm0u2Mk
Ejjk/wLBeURnekHp4mzUSLtuMd5CT47m5OvFaJR4aQiS5u7mcMiL/HieEYzQqraQO1jBLIryAAEX
jj7ni2HgKx4SPgrEM8sYWwOIQUpkjHU8SIKx39phhTrOfs50EFi68ZrPSnzQh5143sF35H+Ye9X+
C4Nxkuf/uWrsD1jklApvNqWiY/xET0PEiCMGZA5ekVefHAPk9DaOksF9V2EnErX9oJycZCjEVRs6
4v7RazfDhRoTVjy7dWIbI8f9s0G6P0Pd6Rj5DIMDbV3UnZ/pGbZ4BLH4CuAsvki7IiGLI6D0Eaxn
gkVbckfTjGr8cXoPqPnqCYtVHA2jDZ2FomiSctY39RCksuRGMZvDmfL8xthnrAPPSVT8RSmv5p8R
aaYdg5Y4TdOmpNgSTCt+YmnpOOyfirYLXZXBPIrtV9UI6+e1oiIWqN6NMP5tRV+fc8OdE5p/epge
gH0cs22pmoWTftik0FSqNrwdze5P5k+K4yqo0tg0XlTQ2r+U0nCCBsu3WeFA/ugZk3C5oYfHL1gb
sSwn3VAcNC93DIdYUNt+zeca4Lwogz3Jjvc2SnAOnOLAaPxViJVZa9c8OuMOpvxlzjZKDujFop4G
8Yc1JcJ0q669yQqBmaWMw+TG2p7xCYj9ZvTHNjl+7ENiRPq8T1Zyq8c2hdmlgIyh1jglJKg0RXff
0cscAinF0NucqgoUcsCQodq2q5pEQc/bF/EZSgn+xAYOXHuw1wIDpvOBXDMQzlWtwtiGkMiMj/N6
aBd4Qae0136rsT/x/cry3++8ztWAmjs5cn2PE/laA8/7blrMQHVdeoneQDZJysZPcwTs6tXXkQG1
cq1/R0/3XqDB9dscPLbRQhL4qLljO6Sw1tWM06RuRSz+6HwcdOZ1hhWCZj/7bAElx9QsPoXBP7lL
Jwv7WKv/RfZ5gT4pQ/HMsHDVGbRSp1agq3faRXh5iwYoMIl43uQL9v5sHVzKB6C9v6DMDdAyLkAR
KWGpHc7mJr6tkQxG1aRd9y61pH7N6F0bXOuULHQR33reaDdV8zFtejo/DrslFy+/K2MIVM4mkEyK
Lr3OnKUkKyzX3ja0ZlsfN2YNMfEHsIn3ZoFHyRF6UABvstcNdKxGwtwxejfdXP5BBq1sNEvRv+mW
qZm66XbYPZOAM4y4OrQN075SJ/653LXpCkz3oEAtcdeChbfYkkBBNF90xbZr0BVkVCQpC36BE8oO
OXMM7wBwbKViM8+kd6ijVygXYLF1KCbUvBASM2DKrf6E8HdQyMR2iZy8s4VDJvEPlRlOGVdBoTY0
+n9tX/WKcaAEjQa7Iww1+nFqSLh7NSlzbjEUXjELiAHcg77CPUWQoSx20nCUFayJYeoKWIvHV6Hn
TrMpeE3geGqFayYHQ+KEIDSuTyZv/1fNqpw0gDfQ+T62dFkScJ6kRlaf8hbpXHgqhv9CZ8upZU/6
B4eka0rc350JzW0S9+4Fb50gRg/xYTn97GSnERbbTBS0ze1ecehiWFEVFOxTrJycQzbQo/o4Gz/P
ZD8ey7ZfNm+YayQD/cNFpYkygKrF5Wh7oB/I9jZ43gkoYq+SxCN4sSTHwBgSjgGY5UpHryGp3fi7
5ZkqrSxYrKwsW/u96sY7X1OhMSYVz8azF+IwBAxbMFN3ezJ6BMMGXgAXl4te1z+PL/s03rHjiG6Z
bUdweujVZ6ISJKPB4Ri8Un6EePedza9GLf2Yw2pZFCviILFcgLKG06lqLwKo48aR0x57UvTy3PAE
xBuwwI6U05bYZh+B7dpNDVq1RftuhvzfcA0WAocGGw7+e+0b/nhW59ZnEyBuXNmhyeSqsqbLXPRT
WUn2HYQ8DZXjJkHKo7q5aAdEfW5RMsAs06zRRPRdxqkmsY9kErUjDHcdcOoq5n4bQxxRZRLC3RaJ
4ijSwmSYap5yycbwBlaCcX5Tw2PwQF4nf9ZpuBvXyx2HBO9ONvwGj3Ti9rt/z0kGA+K1uhOUC/27
xurSZtd6DgL4Aqpa7l2NDCSKH6LAKxWaqIJztojXlbXhQvjzc7rYWoWJJhdwDsKyGLdySMCS0iVM
kf42gNBKBwuAPgQn36yOXBsKtfXk8GXjUwTGZ4wUekBzbRP2WDhlKA/Ax2EbDH38JIQXx2/dKi92
u5+6/ZPPp/strQnOyCWkV9dxFkfGl1hge3c7YmfdImp+/KOcCE+5K9VedWbGFwbAnhWNBag0ghwZ
r7/c5rrrEuIckPwwDvGmMUVMxjO5PREB5+XYtUOWWb8DEkSQd4V57IX+5uEcdBuV3U1xdEYldsWR
emsLZEkKs41/lL25qb2rXI9Nbppu/370+BOni6i29Bv2usBvWH0iYe9Ekaa3vBls7kRkqu+U3K4a
qeKrD9GTTxgAcYPLCCqz4423jjPhWwE/5ZLA5bKtdNvi3u8pwn7LWHWoKYKPQ7XBYdfs2TqR0TTO
Rh+lNw3p5QCVzh+pvEvfGZvaEScQbI7ogIybE96p+AyRxHXfI+XmvsL3yoMIutMY8LqV+fcFViq0
PWuajJJ8CyCy3XyJ7ZjmoBGsReg1puiXZNzw6c8wTLAEApVtYtGk43Sqip/UxM2H3SidsPi15U+5
nfsvJlGGJIKVCSbnWBPC12+ljb58ZVEkz7Ud/vJqVRiPb5EXdrydrvnVPvryyECA3hRpLVHqHizU
BtEaOmU+SEiohYVIw0HT1JIuVZWRUMX9lbMb3ujvUmEZdZNUaCmb3TRoHIYh6vAKbn1/9rN0tjjM
m/om1I3+UUBtgFjQQsbRh8vF9pUbKrVmirOcwleUpndOBN0WC75EUT/aS1Kfc593SLP4JedSHQNp
6iNYE7HdN3uXuJef1LOpPT5CZb0+WG4uHETrq3SuQV4GNnfXcrqSmmPZjRX1GpySU998P5Ijyc33
bWst257S5Cl/8zAyfs9AscB0h7kZhPBm6zk8wNI4kPrG76g8idhcjcFs6q+t+HlN+lpWYgqkqY7A
gOygHlbdFXYS7sSndkWmM2ME9gLnJ+T7r405p7lvUz5Dn0oHoRK3GWnBNWb1WzUGNGbNw2lagtw3
5ekKmRKRIFdGCA6TrX7oC5PKLzMy+i+MZRphFJLENmQhJ/JzKu/CBM6hPam4ikOE/mEyTpvFuQyW
IDyv/vxfKugDQssWRp1R4bRA7ETCILzSNd4o0zYa5kuOXDN/sbkoFVmevlWIt0yeYIfO74HTxgJ9
2EyAxFUaTEN0/GQLorVAlALMqRiooyKktsJgmNSocB0bk10Y58fEm355VYvg6ws+7zsZ5YGzaPeL
dnRKWhqsc3wpVRhiHhb2/BJY8G6DTOV4Gh87lmvpSoUeK1Io2OJahUDL9dCqZQ15lhMdS8J2+UxU
ap5whkBvWc3woHseg1GiZl+hoOZSlSRYNXkknwTWVbgoqT2fTgnQSApNCNsRBwohQERUyjLDiwJp
kULVq2U5zV9yrP5FCyFijs8LXKTUV2Ov32s8cQ3WfGd6PIAGv/6ubHECFCdGQBOiVwW5xybHN9Eq
X2g/ADU4e4P59o0w0rrEjWeyJ3vJMFcotusOUbZHmD3FgB5JDE0myFjGhzLryVBorDkqJ8tvN/G7
i/CbtZkhlq0rJWRZJEWGdm3eGaHnOFsvijaRawsMSAhH4sUfFGrD1qGrOuyuaNPj5Lc+YOE8QKKN
JPLKPxRn7XZQmfYgXD/wmEMSYDXo4xw94+dqqIQ1PowDZYM6vHfkNHcpsBsUAYhlLm/EixBBTjh8
TcsQNLFDNgwZc20yJ9P2u04FunN6Lznl6ZV5kwr4SBGKGaiFWL/jLGzSItyK0zhBjcyQgZrxQPpp
c7R17byJEjIePoB5WcjLeHcC2IyAFRk1Ke8LRCUvCgu5D1XfIqQZQE4D8nAaFAAf8txXKMIS6tDM
i2P7hrExdGkzFXLUgE8bAbH62iL+D6BYliXmrz8SDkz7oona0J1YIyXJEKLAGBPlmgJ5jdV2R6+P
tHdagAqj3Wq9iVD24oMfXxjWksx84QLZGlb6Tb1KRJiUMlu9fUs7llh5YB/Pc1r3XBTGciqVBwDM
9JCZAl2tVwMvWhbs8xtOV0aEJGpo7ITBt/Za/a/DRm5unEAopqEmy1AOrYHaHqIts/Ry8ToETe5w
HAtNhTzK/tc0WxsO+Kfs8KZHPv8h72YHK5FkZA7q/JRCJievbHPU3MiQb0sHA+ljACBRg1mxH9Cp
MTx0NEdVPNGHK0oIuiQcQivX/me+F2C/MuAJoYB96omn4v93BdLQCA2N7yenFF0gL0Pl+VkheHKX
RRpTFtrwMDP1kkec6WA2YdF0oSkizv6X3AR7u+XRuW2mn4foRHUel0TFXffAKywQ3a3vobX4eX2W
yVHu0LFQ76G0RLbAxctA009gjJPW4braFkam/8jvcddeR0gxd8VhP6hder0hM+MsgVvIgyi7uQft
CSAftkbHQ3kNe5J8pu4ZeRxD8TVHtOc5/Bxtk3MksVi96hEnOlCxrzFbv6Mr8E/MPdkLf/z949Iw
XUH5HPjHHp2T3FZHFKlk4hALNmEqyBR6xTslU6TDc9FA5e+2EBMi8lkbV5+aY0/KAVG29AWJQ/P5
txUONjFVxV7plWgCATyduMhsGoftbrBv8D/+09VfkepPLEdihzLjyIfm+JQg6Gv0lzpJQ1rGw6st
o3QhMsbOIKRI6QjLbF+IA1pUenXKUvMTxLnAKBXmeLmFbtdRox2lrSCg6H3gITmD6GKIkSmcWqXq
xjmrIpoGS66mat1iPKoaCGXNZcz4ZHW6B9xAlk8TTiG+gKYePARg2uMp95Hwdk/CTav5dWMxDLzG
Lne1L3/upsoVOmzp+YC2etBE9F0tNjacunb0CNlm5B51yVpEynZeQcP5NsD+QzIfL2nfuMUOEveI
zWCx6J6B026cfXvzxqdKLcmMJheV1mJBse0OoJoprTXhHaz6QNYLk6yppjmDyY73QK14xloCxz3H
s3HS05Y7eIAHT1VAkYq94c2KpPxAl1IGyqal/WUMLbJZpp9TeHy1zzDMZe96lYE8AyaZriSBAO/p
+d9yL/hkyRZU+mSs8PpMcHUVsUcOQ3oPQh8bx7UfkJy7ZsIwYe4cxW9/xKxwWU7mfT5JY72/7/TD
fiFxnggCsDlZGxVlyQ+UA2lcz+0IFx6Dy69oNK5Pyvqa4lRdG+eJ5scQ4B7JPhi6tbSP42Y+DyN/
TwNEFDeBAJ2O2i4s6e9fL6Sg00RH7k0MMgrKEpJs2xAHPat21nNoRc+iM1r/SjmfB7qkJMrQixv9
uLeyQLjiV3chfnh/xooCfhJOR7x80n5bWBchRHEvjcZizc5Y0KLTQbLXSmIwlCfBqsiRtkcm4Ez+
AD69IrTEa3dIAnyTUvRtsozPMFal0JGeIPs6BDRa5rVWcV5vPMF6mtF8HVBh2Y/vf7X+lYlJr7KP
DwcFp7wB5FyIlfIjfS5fjALRItLHTG1yhX5K7ZQjTa8heTvmwzUtO9+1A6YB7JWBzR2d1FDrk0hw
tfVkzv0uUWj/5EcTSsnTRTq1S5pzy9tioWTSG4IqdaSe0C/T7J2RtJNnUd95emqZOXUHFCag5+GQ
51iDcxlB4sKZvahmR7648l6t2TKQQE0BW9kUaDmnPq46GsntPe4+L1V5IbSRE4zXjQoPPP2d29Sa
6H1X/MT7mTwGc7sgSY83lmNnsyGPOFA9uniLacknoZXeOhQ9DeR5vEjtVJcxz9oYg2Y5FgnJ2hmh
XSYxJCJd9OYXQ0omJRO1Dr6eeCZ/a7AY9u1AbXxtEcPhYcV1w/4W1UUo8ztvd+uCBFidbxj2iN67
P9ZBZz+BjzpO2ym9O01yrlNMlZlwNpojObPkGyNRz2uh973GGNDtzaZohx78aKHNWAU5pVcJ2WtT
BU3FRIJQUsmMF/soecClKD1ytwOH5acqi7yGDokgOZ3cGw5JFCul+z055QA7HSBwlgamebpsu1f3
BLae1xVuMdTkYbQGey5BuX0/of0YRtMOffWOoqEMLVzGTZwI0Vdf5+sJm4eUfiCH7SrQqRvM22xe
okQkZLfoP/PZaCEK3EmtUggdQF2dYgf3kJSacEcueUBtbCZlBQEcEmMnL5SUrvd1PxXlrOzCbk+K
RjclgZ4BoxskHQ+WW/MCJMIhly8BRvRPYpl8lLiWzR6G/tTN2qUxjna3FE/WgMlT5LAUf5YD+bnA
0At4e9NAb0sb+rnRyHfsLYQ7XcfTbxnUtiUuEpdJx/UtkuLb3EBztWPJMs1dnihOb4E9lV7RiquY
abcX5g/UDzNsq7sFxjtBGEqMbpd4jRvzPo/+P02KrBuAPLd3nAxQoXvhUlf4G+8NMoQpxWs2SnqZ
7YEQDUypqLqmjXDPIyHqDINEaMB1LCvKuTC+pRTGdQr3orCYj6Le+yEToPsOFglKQ8mHof8H/REu
6wIH71U8S/05GtqDUWtjjnYOpmEukMDhhZ1ro0gibwU4O63EnnYNQTA6iBE+CVq5ljZNFiWw3zeZ
VRiWPBP847k+w8haqmHkO+7aBmi6Opw6OTCtIxCZc4eXNzUFJGYwBrmwwYVl/CSDL8ZXRHzHJzFh
KFoQL1DUTUSlFJDGdG3Qum74wArc+VjkJna3EmrWb3iVnDrvK9JpAbrv7PGnVOaMm3WENV/l/CoS
5MRcDZ4KSb+XQCkQvvBDonXVpF62/ewxDW4ofuGgEiE6UDP05zu6YkQ0bCvy9fH601ZC/DtHQu2i
HFSFPqST8rGqqbXZE679YGXHr7NzrsU4u8R5XO4PXk8zfAgbyheqnxjGt0LXmlmVo6Wmu8Khh9JM
SfHTDi7ByCPVw/TAiGk9T7BnCc5o1FIcVSX3GER1c7K9IM0Z2oYqyJJxHzF41Ycf7teGujwWGyAV
Xvlv1+BJfVOTYRbgztcLEGD92jQ2OMK+4Fr+jFEPxMcIdWrQop4L0OwGUmu4mqivTGB1OYgDi9HU
nnsT159ztyflWRyL5IiAUDtixeoUi+x2CiBBL70ZL/b9NRBCGwUii7K1UZ94oZ4CUoNsFz3B2M73
pf9YJe2hvFPlqTCQiAglolnh69GYvz//sdUiNN9NhgE8q/VOWPDQx+nhg93dj++89RJ8a0O5NNWm
jNkPLQm+zX/5uLn6c9rvs2RPOtXZpl225nxCjf26VtDDPd3CpFztISEis7QhNO0CE4misB0KWtoj
QJfoBxFO7V37hAF1x60CgjBh5cBGL9Vd/mgMONzMjHcaQsCZo0bU/wPkFkXY/QgFm0OHRDXvzfQD
3Gc30XQLnHNh8v0X27QStb5Q4y41QXcEdzQS1TgnEOI60wdy3IDnlLabuc88ic0tA/BJyp5rVBDy
YF2eApkVQ2ljtVsqBVuyVTWpD7/vldTj17Cgi7GwFJMPG0x+FfEqjl8ohTW2fsNXEzVgDcAiz08S
GeQSarLqRVXgBSk4QlekdEQp2JKIkNb0DHR8PhHy3HNALLPfL70NJkwKOdtorJfbocXbpsUCSDIT
Ct36u2NtLH8TaFt0KxyGigW7z6fCEfF0QBjK9/urxT8/zpajoOkcplB+dO4/fECT7Kez5z5sQTrM
Qc1wbbrg+hZ68NobZxTkfSvLmQ2dn+HkRdz7hSxPY5IuPeikjzaxkFePrVI3ltlSSHNH28acG6Sn
5rz5JC3v+PdoedogH3WRRemalq+8jbCpOLcRaCG/OIeo++8JCLMbOIFz9czCxUlDfyfgsDBKpLcE
h68uYwvq8LoViNBmBlDXeCLR/+02mHbqgL3h9qsNkYCUG27sFCZAhZLk0FBDhZZPY5J85sHt4RfF
1il8TlYaG9ZLf9Mzai0bG9W/fMDbuNTLmSeUGGYgo8HzbOlLWTsHmN4CH/zlBvJ9nSX5+MTmZzmO
pVRhZ2PCn4Kh7fcSEX0UuhCVzroCr0NawPKrjg7bO9FDMFCoghi47OyDlGJsw0ZQOhcyWUyqGofU
9lM9+HFODzyz3aMOH88dEMr7hwAxtBdM9MyV3zgs91HqSK/CvF/wTg3hETQroS6wV0SgOhir1hmY
un0uBPRzCRuujUTkzTqPwAi4GYOfJ/oXyltxk8Cv1zv2jCgnrZTxmiWI+3oTdu/PLTihMZyFYDG6
+6alLYcAvo71JaFqDndSQvMd69ddd+dO5mQGhbKIZJg39xjy+W0zwtJ0INgI4X3ebFc8aCLcZUsS
ahPQwsVXNi81ugvovAvfGDohTnF1VM0drl8xb9jRvDEB3Qxemvle3HXP+gfbLV8f3KrK34R/5NnT
az0tdNGIP+UA6MyHaDakaM6K4MezS9Y4dbbtsgLJTZOPP7DeWRTX7JdKR1f7S3DVY/cYVnP9riOL
2PmklQOv9K9Q7lKn34KF7IdKGC+NwddXiqwjCrA7CwoMGyY7cPfpGtOv60+VqzGnAicqEPvbakfw
sYdvo/l2aMdM3HN/w8R9ufvup1sQuIf1rGe0Qw8tIbD0XHU83g6UOSuune9CB70HMIYUxRxlta7B
vnhBfbHAFpVD/pmk7vnQeDNOWJknenEqooXOLuEuPNQB0c7mRLNUtUNYCvBXdgjK6QbUYe8aRQkd
+gdTeat2+Ub9gK5YWPuhlAghKjsifRaBdM0LVRJvm0neeOBLABkknxyYLyav1JIie+SPdv9dwSvJ
ppkBLmfozrv/pGJHI0pplKAgbXI05sbuO4EqBtjlUoEC12uioEhEyWRk3les8tJQlZ8gCRNQ5bis
IE72qHu+b6CgSr5b8UG3Q62iQag6vI5HIyiyuoSaVGJ6ykqgKWVnDjisgW/r7whuitdBr0eJa8rI
o3BJB01f+zeMBxdGrGRdSDmwiOBf3mw6Q9teGtmHh81ccnhcGvm2NpVZm5ov6vYewr/Ni/BzLRmh
bB1xJ1QdlsIhQEJpHvi7+kWHsXipT3so+eNvF7SCh/ZpWZ4v+TddG6WZPWmzoYZk535Hc7s6mC/L
ey6Hz+MUYtCtTjSYXzZjWjQV5cbJj/Tn0KKGP45xBqAcmchZPj+uOW8qRgpj8/kICe73ThZLQ9kj
uhhkFMkmZO1KfjXtLi5PjTz4acz7plZUnmMhAgoxNtv9+w20hqJGaH0HDw464NAMscmK9DlkxHSk
+2KF7k8dK8GEBQ78+Ejm66GZiKRDbVNdwuJhJbA1MHeJoF1HCpSwD2pvJpEENNGtagVDQ+IoRVNb
JF3GQuL3t9qYpUavu0g6BkDxCaX77UvH0odt+U0jL4/hhqXUEZQc0p9lurMgay4r7y2JPIKPDYQA
gkAzDwa/1JblAdRWaKA4vG0u2hbFd5LH++jit4Lh8MgO3AijzO52yCvXAuNcPy8PQuOZ+/pyyE2O
NDpu4azqfhAJziBfmaezGTZjADfkVCo3uEy9ONGaTfgVxGCD+oz/jRvbhZCvXS7jxiz8oSDN3w54
fesIKx7SZ8UyiSN24Ny6jD95+5FhN6cTJmW+l3ZnPTgDz6ONkKsuB+qb9MW2R/tJWU6szbfVNSaX
AyGiqGtits4HN4/3WAyATCeRz8XzNPv62GPR87jqJee6WPLkF2ei8IR04G/qhbDf+ODUloVXsUsj
BPWNbzOeEvuD5jyn0b2FPwO2ZPSviBRmaHdr9UHQr7RAz2ySjoYpLUpqZ33thNZMi0AwGHxb9AQQ
Y1+dO0krbG0GjnAbdx1Bdm0VUV2t/dtJgsJhNqKAhxuTqY3GfZCnyIuiAMpnvrBMubDfURwdiUks
LJFhxekHN3kR18l89OwpKjisOJOnmGdt1fQ38fezjjGddMGRYmqFD+ex+PLnRfFWNw4qF+HQ5C7D
/3a+sFzEtOroSCzWA90YAFo4kxoEQl8lWblC3jJoxrirlyh+BbKgusnZ+r9KwhfUOZ0EyZGaXbkH
DUntUCvJhwnCmdQgAgS4U6koA56t28mC1xZULqR8lkDAeP3cUCM1hmXeH1/SkW33I61TcTW22LgK
VnRjbBeMEq4s77rR9gmFA+e9OXKIdz4x3aRTyabLPW6BXZ4vf7+deU0CCHwpEyikmhVkyvKHRijJ
KEKTdLOjVyB7ylZHYdWW66YCa8d62TWOKGO07nxKVSoR2v/BHH14Wf6qGqrM/xYoat62x+EQNepF
sOLw13ajt8KlJ7g+XJqKM7scAIgtySK44/GnqCbV1GHW6XGjV8TRXISA7q1rVALH1vbBOF8OBENG
8V4yjofd1S6Pqd5HnAC3MnD2BLt2/02CPBmlFED4sFXCKP3zyS8kH9QLg1IgZgPpUXVBfrmC6jZy
327/1IpxzDY2Fuh1ZQ3uA4vSmgQjxzhMUq+dyQlu+/iHoXguqdZgCImKNmQAYKnRg70xQbUBC3rP
4by1Vgbw54zfTFTyTLxoYUwJfDwzaOFIU6o1e0lcLE46WJsGn5/0IwlZR2IWxmbWabjetxoI8Pcs
OsqS6Fm/HBISjmdkAk/aNXlWwsRaCHGRi6Pn3Y66zOMBjgpB6i4VooF7c8ZnEguVR02zKdWJa0MY
xXe1z+tmZBVaKL4CaObjzcWl5k5zUuy3hDalm9m2nyu31RW28O15nlAm/xnXdxA1BfpNyjNsLiAR
7E5x3LgutoC7u2mw4tAl5Wbqea7p7Ay9dl8q9QSJ8zJqm+zrkvgH3I2DhyW1EzX+oEOD+eBY3580
HNCqN/d8ezpM5RCSF4RYjPGeqXUJFdG9htm2L5Zrw3R2r5Ob6iEG1DKmzuQJErL/sdqu/GYJpuAD
gaKfrr1hbkjiovi4k7Xs3qggGF7f0WvairpjsPZZ/0XNmZvEIJoCNQ73QqfaVeGOmoOIZmKMPLT1
OhILMWaxbNy2+o+U3P7LftO3y+umLyoDGhpp7x6A1Xzv2spsxoN1iDUiXpll5akkt376G/Gi88w8
JuUEnXbUu3hzuIEwzurN0Zy+Yt+iAgWufPACGqhnTW9tHTMLNArkHVOLcakd1L6nnSad9qFPuU3B
tbQHunotfHdVjfiQ4Z7C/9tNQMTJo2fXr6Vsd6Bc+1yKiK+vPFLSCpMxJBz7x1UtzaCPhLhLfpbO
c4fZ5cSYrNVsmO2RXWtd6j4i0UlrvLAh/ZsnEC4j8QnZlWUz6VKZ/x1lUfgPlSXpEtLH6XSOTGzG
h4tPrKg7vQQgC/QRlXJYt+pTmqLpg7ct39TY5qNVKPTx910DQRuQQgqNB2auO9vZnw8A/f2h11/Q
unciytXaaYD9i5UWUAWflvorIfIavq4e1KLYw7dWRY7cw9gHzWKYgPAk/pFGnuTinvc8ks1+SzDQ
KWsi3K0hen8cAqyZlwpEHal5GjHk3+R8kU8GjcDEs9XXHo89AGc6U0fdi7mnxYjDxU++Y1GyvFKT
+QLTN1NWRev+kj2BLV9r4142D6IpkaBpi+zk0htblR6EgCFnohW2CjLDdxbvvNCfzmmdZG1pgqh0
w5/H+rDnMOAQk2wgZ4HvFcyYCg2cUSmq4VnojYLYFAfFrlh5ffYSub6x3+ifID/yzHIcfqFQQMo+
aCz5jWUhiWxKnfj2o82QefIbUavmkjrVj3ZrKH0TCi2K7Wnv5SiIFBD2NLnYA/Yerh0wd6ZhQxpH
rKcKI7AIdsp4jj0PqsLZi5lEZAZwdviCY4ybSZeu9ltfg8ds8FxfNPvBIozR/bVSXHheRK52PDT6
JnYxovUqbmyDwfCHYKXiGkLnEqZ4jijDySH2GhCq0uydH0zy3mygSSxCb2+fjVM+D3czmUbBSTsh
Rg9nLUDnGeMQy22YinNU0OuKuKK33Cfytm+wExvBxfWNzUcAkg6u4AJzcb/o+6MGBIT5pSfrGT25
h7b3gsoft/p/K247vD+OV6ocLfsRYXCTEbbaHxBcVAv/M/dn61f6GfZ0mL483IC8cg06vXlntudj
jWpo/A1NU3y9x1v6A8GwWTeWorhFnsgLSdMbVtfjocwLA7VLnMJ8MwKukMLQRRahnFwGbaoZvq6o
zEBjfp0kxzs1G2BaF/Do1GGT1UBlJDsp5LI7rS19CbFuXlIG27AoGG/eh6jQPft+MCxJfXA3Is5E
5mgVSL3zLpgac2+r2Ex//q2TKbHnOAVUhidFiQI2hMDHN6EmOiOGhw2cBEUTxp8bSn4nwXhbe0Rl
rNVbuhPrUdfABtINNTq5K4hEQA9RX28oEJ/XiZQAIHgPJFYI78aYX3E0s+AYBZlKAk+bWrJuNoCF
zI8PGb+WK8nshyEsEYX3QCtae6RLoFvvUqBKMMelwc5S6E1RypSQR+ZebWpX3IlYPesFd6UBwM3T
l+2V9/g5tKdiuN3s1kYKjGpe3wcPWt8pIzmmYd16F+1MSk5W75O9h1h/3C1ERA6FRHVA3iQIRQBa
f4JGmNXlI8+QQvsULZc937COVRcXK0NBgyfbE8lwZcYLnibEW/9YWN6h/9lrbHlNORrUv0Ilq+Gg
YNTWfPt0aVpj5clUX9A9yN5/ppYk1wYd66ldIp0o93PdLPVft/Sl+CuyMMrKYl94vIDP0hF7okha
w4Ro1zC9Uu7ErbzHNNDNUal6Ir/YcOIQRFaRSij6duBUNsPMfxpEtuWWPfArJRuWu6nBdYoQPnpO
pqDSe1zWo7E40vgsv7TMrXhJ7LpS2HIs8kN5vG8n5pt5k55Wke4lih2IlVkD+xeF0dDgbdTcmzjN
tyF/KwlqlezoVh0vkaDYkCci5vj+C9uO7xfiljIAMszv+Na5/Ndx+/XCGrTSzjz3p2B0ix+x4nN0
wpoKnsqf3+r23RSjbpuO0cABLrzCo3ag0GODs7dIxPcmrULBfONRl1hFWpKqPGOAYScssc9n6y87
lTBbmoZJNoOZCT3OzhSHj5e1cAG1RAbeCUU8I7GFa1KBTBaCuL9XIFC+6KmfUrFQdkDTMCzQpmpQ
kbHA7GVs50/FdxFYBbMKIuLJByiIOvG/BsgVIJSDr2EhGyBaFH/hgf1OkHmf8ZzuKrmIExXWLEpb
oS7VQQumTj2ZRVEddbSQiMsEGgu7dM1VLZcB1t+l+Dob4sg+5LMVg5S35XzBXEs12KHBLUQgzsOO
qkUa9hiNI2tJvphZR7aJUcYGXQqhd2Ze08trZPHokAiW1z6xE+kbsJ3+g3f/nNpH1ziLHPUSQ5i0
q77r565Ne+EuS1QGMf0uDmV6gayYc3pMxmwmbuXemrqyoyxt1VHSYBs2tLqsEMBmhg9TWERyx/tB
rrKXevIYvnS3tPijc3XtdimEkSJ7aqaHJzs1Rjd3NYeTWqS7ThdKzzKZsGUpSkLVV0se6ffKk0tE
CMbflObs2mF4Ed26pvlo8R46wd8Gr5GnwY698XC/dg6SGitBvlgpisuBAg5W4LjRFJR9Wmq3B5Wv
SfhqbkaTLNYn+E6ZF5HNJrkuhoWRCW0hlScQMc4Dx30N07Fk0EVMNhIOkmZhsg9NiLdjIqdhn9mX
aaGYZaC1bSCBPdf3oldrMdECRayPRI4S9sgGMh2Qjb4SAIjth14VZnerknsrs1gDv2/NTUetZbz/
yAbiLf+LPl2bCUhYs6I4KRJYMxZuzblGcVhcXJtQDvJaXXu8DtFP1MJ6o6MPKBvzJ/NLOJziHuGh
2Z35kA5GP60gK4NbnC17QBO+qZO1jSbm1fhJg1e2fCVRPaq+FECUBvM8SQvyFfqFRq7dHTHueZKx
SVqny1try6Tqc1wNscjt5bLS3ARYMn7860ubvPp+AWYHuzDAEtZBvGxja/YDtJNn4fcBjhpbidRt
lYGVpd9sZzLm3ynVs6mDpbgsj5HFLu144oCFfcMww9s6N4I4DUMKhCNd5pLRQTeYyWPK72YItMNq
GtJRKnmLm+rBJeRLa4tAOsMppf3wOWUc8CTsJ2QlOMAQ/KFjiBMKt5lBalmNsMU+5svb9ITYx4nV
JiEDRuXQIfMoRDIdmFAJMzon4La+rqIYYV81WxxxH71N5bTFp2dbD1nU09jvQ+IZj5cWao33GzEJ
KJpIHUsZ8AU+4GM4RpC3Yp6HRj5YPOQ6Ur6GLrXw+p0Ficie1TOe5OCObUbKXgB8m+K74KZ9w3BV
JWOtNY1HgJgruO85l/FRVFrS7lyA/y5zrKzU/g2DSXIZbYp4MV1qga6r5dmFxgvp5eWtbuAtSjEu
ry+s+sQWunacebMomeJkGPxvIqEX+WY1gVw0nVpVXYeuEESpmIqSWTJ+QgiDwcNA2x4WEEyZMJpV
904CNwx/ybVtkgXEeO53IY5qmvVZVGTkLWb+/n9oMBfTcDRbRox5C/QctWRSR4GVsiv8I4/37XtC
cSXNE/NoJHbpGMCbyFT5H1N1hq7dycGhhqAPVpbrZZ/4QtuCvU694gzCkvhiQBqZqLBqZPHMZJpd
8hZ+z3p9xNcOdlvU93Y38ZGuqtX1E+oUeJXDaFJaXm1sTpjAWvT79974ly/oJJM92ILppZnbTmzt
yO08mxMj5wAH9u+YpjzdSxvpA6GHcJkZA+U0C1+b9TbUC5W5eQVc0E53w2FUHuG3FmnX8+0Ua1K/
8LD1VPZCh9l/SduvqKPGrNf+gldXdugz2zcZu3CQlpHRTpTyc6BuAeNYPB3lbSe8p8KIOaFe4JVP
2bUxuqCHr5LPnBf0Da9L+m/I8l5fqAhpuUj++MTV+V2Qfid6W3WNuUwnvi+LmdJP+as9y/JxlWcQ
A9KydqvYVAWOCeNrnBLbCMGq6XY/Y/RgVL8sYV5q692OtwfPyDAhtrRHLN2XZdzRdaJDY1acxKk/
b6CYMx97C+EH3ruPGTx70Bi3e+lfmBvxUd91NdEfZjw0JAvRnB1n4K1V6sgxS28We3wJi2SaVAKJ
99rWngEqugSNnqokJVYaugoOGqBdSMh13cZo3RKKW/NuSz2HtekeKfEcYqkbKeiTBdlXYYD+zvVK
tMJszElPw07iXj3z3Spx+HpKjJG4yP41fEpeLEXpJCfQ0jYtV2dRfqphQngAzctOYPQk84+2/qoR
kQqdaBtRYl4j6mcwtrpvp0K5LO7+kLZDsAYX3WFNIFbUhNGlbR+gz8S9wThpopStOGKZ1bRMlnpo
BF2QwWemGBZ91km9fjwK/5+AJRIlINkuA/YRRdmm2geUSuhLyvxNoJSrQ7Hc/q3wQJO4Y7tQRfON
pilquefF2PhfHCyjMOrdQZYrrnrp1G+ZkZmROZ2KeVDKHdhgY2NuO1PuWBkG0eZ2dmBTDfaplHUD
OZuq4AEi8XUhRzrbxr7V+rKIMquoAjx+REpbIAhz+GA4GkuSjT3wH1lqIp/rN1ZzEvL9GJT5nsb0
UgJqa69Qg/6aelZSdpUwSRi/VAwJz7MhyN1sbojNaehp7PbVvwCGkiJQSBkh7/gi3cq75UbFW8M6
Cq8RkNnngowNRT+FIkUW2GdNIuE4ey2K4z1Xm3SstLMrLXRgKChtCxbxpONurX9cVbnmBK6r9cTy
RTNT2+c/1l+OSXTDXPIXJ5p9DE7tX99bco6xFJsCrXtrk754L1yENmMzyx9R8sPUNRrAj/FhFbeZ
ZEuFelxCT3xBMlxM4T17RCoavmyV2x2fZSzA9cenn1sC70fyMO1sM0AaEVVOWHD8IRy9BOjzaqLd
CHACReWrbDT0D+Ghy6NhhZrPrUuvmGqz55tun0MBERFzPNd/kUOJ5XYt0vt1cA0I1n3RJjRNq4v0
mbdYMInvHUsR9v8jXT3biqrFqaoodVYFeO5PwtWwsN2s2HlX5LbZb3hoRrX9Dr5+NiSGbRmg32CV
4+GDRvaC0R79qp2YpU4LqQuoFV8BcZ8ebv0Hw8IA27GZCVKf3k2efU12bjcBbm2NSURI+ckTqpyK
IVZYaXIEI97EwiuNLmK6JnWoKL5dIX6usE9fpapZGEu565TwPL5VUpGd4gjVwSZbmfW/RCvuzqUE
4TnSiahIDSqDk4AqfrOWwhoW7/8jBRSb7nZPnt9vIphM5/WIVsVnaZfvLUjjWZFN5LYbLdcyT5An
m/6YYBbqHd/2DpBTqyxOyWJsijhtuIgCYgaIUL9KsTac3m7qMza0Q5wLBB+qRKtTdDu67h17AQmo
wM+V6T+LFgta9lWgaM3uFwvH4fgVoigXe7T8nDLEQU1cO1gJyvvjoMiBGgi0z2N5Jq3C5mMe8L2h
3zjxp3MOpdPvDHWLdaWx601YgEms5h9b0omDZ384Nvtek7B6O3zWjWu/FTipOE1GgJ6annePweOM
S6PWaab2kvv5hr4WHuXp7p8ckCjZ+fcKU75w611QD9g8f6rVQCFwvZ1zljD3WwR0iyza2DfFSUfQ
cjjQiWwCLidTs9eIWNw/2kjs3+Ody3IKaqFBpxVGP43ncSPgQv05/ZsKEQ6pTpIKfWUkrrQUw+wk
AdsGjy7nfGOdn1wVjLUyvPUuDi8pi8VxqIb6f9WLVcA2JMa1bXYI9KBqFPVLoPiVdoy6eiqbVwhE
l+GTh3nmmSLuWfBlZrvpWA0t1qf2E81CfJhr+PpgrBl2pdc8hO2G/kg2j0UIBY/sCOdipmyLpdzz
y/Pvdn+As3mJnW9t0fkGOZP4yZVT5d2u3IQXNCKb0YISiQFK/DCl18eznQnTbHnvXhWvHvjPxF6+
/TaNI//Sx2k03kTWBHUkSpph72oBqtqg5r39YMUqGSVieJw+55a8EievxIVKc1j/6dttboXDobJC
HmfnVj6xmv3eD7D+uxjhdtZ4sriXe1aOdTjg8UB72PFtKeFw0wsSLohRRJCwk81bG+R330dTdHav
diAnH4MTbktPUlWgiSYyb4TPPb2ERpixyPm6dgodgyB+jt2eBo2KURhwi9L5+8FuH92HDWFgoBhw
UwXUMsh5n1q4MAOoWT6Xd3kQg4R8MZCVxiu7sqRhA6Kz44au8VOIAl9o63731TtFV2aa5pABgPox
QnG5FkspCrA4hSxhYHNW126uVVmA1vYpPfSc0Q9uj8GDeWrqNzpkRW1ux7IcgjJEvJqz1dYk88x4
muSLA2dCi0YfoarHRAH9szKy5ilYkclpjWNt8pUmK+n7gtmar0fofIxUwW63dP0TGvQfHsDrtCyb
ZaLRgg4UfC7nactrAWO/1WV7NgJdF8r2oNZE3XWfdO9WKxVQKFfmysa5oayW7iN8kvd6+yesMcov
cZ1QCl1oCfdS44bWksKo3p1AVw3ma9+KKiddHx/nLhjmyRjgXKvt++IlYVI21F9IhTYcgod6wqx0
v23a5o/prr+gP0LL/AKrvo6zkYXsT3g+SYSdsR/IYPzFU2p5Jo2xkc97LfW2KOLVULUOHQgbA1xU
1+JgMCd8Jvw1P1332vVvSyBHfAUK0DDavWmxky1jkajZUI5FTy9C1CFBIxFNLAy2B0bXVKDtHx3e
ul+LhoHNmScURhEor2zUT0viMDbCgveIgGHQE+Sm9iQGNDNI+RyimBIbJnB1TL8YPzEQo1FvFs5f
Y658luiKAchSNQkYt8HdoiXwYjUmx3V0ycKbDJ8e770LOmj9M2FWeG4GoOJOgCGEECpBlqqM5+uu
JVP9R45YN6TFCZsv8ZTBFuR+rhF2QVRla+yFQPqms1PptZmSitHgvL2f80nLbaUo7DIzV2Amh9Q+
oNJO89245z+hXJrVWL2UZ6zdQOnYbkUaoCpekxd8/Sl9sBERuYGUh/6Tx0SITUMYFTVHiGJ5EhKk
n2wxjnH2oiD2pi94AlF6Y2I5n9Zzg3rWU3P7ZTRX9pP+XTRmovXzCxCniBbDPoGmH2pKUtw6c1VT
SmOR5mgiqsWsk+P3FLNcNwCaUQ5k3y3934rvMQsN9sIdt9HhxO8ah+wxRQ1ehjDrRAX91vXf2PYz
kcN+eegvsI2YpnVIUy328aCDwG8CKqyTxmlEDpOaHGq5o4c6QAxm6NmMGarVnpGlkm0jY5cTtvy9
12961QYqL1nLjVUMXlMm9MSIY2td8AMW9Vh7+PapSOK06UXACpNi/zU+4gTCfxXY7x+4ROr1PQdf
bjMPnghZuXpzsqsooGVS/tan083bcgEM24UOjKpujCXSSkg8jfT1xH6cMP8Cwd69FSWaz0Na+WUU
vQZLE0b03JaFXAYOYgbqjJAyB94+aSMdCQaFxuUHbwOhJPpsbJ8hUMSj36C5COeIkTSYrroAJv8W
gswKMZlmQ0k9ZhSA55ZLgPca2kCzv/cpz/gYR5ZBau3Kl5jRKDU6nrRx3tSIcP4D1lEddjC6RQhb
x44d3JOffOLhdps225lYLbKPq3qV2iOY+ezS4iTI7S0LfVatX1GDKkuNEdsQW6g+hNZibBcVcR+K
t0YNPYREBoo7n1Q1m6jVjCC/D7doViWP6yLHBuhWO/n5WVNa2K2SyCF0uDe55XhDLEn/7h/qK3cl
ouboXDmNDP+0MZR7REoCYbr383I3gek8btiuJBCOhT044PQNPPK+Xgfnt/FSpy7nGSb7Ee8SBboj
8z9PtaYCf7Nde9S+AkDmK9pAg63KX5td9mfuMsntq+TTtx4Lr86GOgF05GPTnNJiCyWeWccH7biT
q716a5rvB6Dsjm+hQng71fEnh88PtDEA9ZZQCT1i8SQwRsVwS1J2fjIIrq7cI1Xv4d6BOFwYDngO
todVz1bqhtRUR6Op3wNbzDWgz5/BCTyHqs8JrxsSO+Z5VhPG9rDv8/QsPMKTO8vrHt1ND4R0QpCd
cJRE1nJ2exbSfyvfHrcvgn+u4dqrnQXvQ1Cvwh5FG33ItitmJqPiFfrDATpCgRnwKR0JODJoJAiB
f+WApuNgRzIl0aRuRIZZn0AORvHLKjasiOdFirywy8KO7SSwiBxwXgndUmwwMVOFEpeqeHSbeP0t
untZlwrjxeLwjNV4pCyaxWW00g+J5Os6Xl7vqQfjbqNG3tyXXDSP+rcGUb33TlGElYnCqbtG9k1s
Az/9em3RbR2QcdwNllY+tNq6M9XQowyNKoPl13ojON7IXpNNkTb81XBbX1iCVcaLq1P00podzpYO
osHqPabMhcg84Ar18Sfb0BzlVuErdQjLgcSF/AzMwpw+QFS7Zmku7OJ/Dx/jQamnS4P3ZPRYxTJ3
sdG2pcnNo67lRqnD3HkocLjt5+bXkhgmqUhvF85gzKZLeXLpMDx0sZMtMWKb7enDgTEaKflyqL1i
USHhE8zPY6QYNCaLUwB6kQx1sTbyzMqS683Hpk2xh3wF7mPh6vtc0iYV1ZxtDDQDhtgUdWM7CKm/
YuYZaASknYMJFwW0iXfXyE9zDVIIilq6XusqAlr9gvLGdTNSCi+wB/C/vtjYT9mLfU5VnGOtUPLQ
Jp50lgu7ckHmaijCyAWSfm+/st7T0SUFPUSqSwG75R6OGTVtHewcH7sqI9Z2E0F2yTYU5UB/Tj/H
GeHweloMNV0v1mb3UXEtzlVIuntnnDdhO44sppdYb7JLQtm+Rk4Fa0GtwgHiwQipDyjHY4NC0fNw
wuiSsc0xvumARHiUK0gZjDFZLcuflnyHvrmRvBa1Nq7SgmdKeluaAv2u1Vlx1oxoWwc28g0wLgIw
ntF1Q8HuWMlUf0hGsRcjlozPkDGCJWiwzsIzve5KopNJuMfq56VI90i5LaPAq+SDJvYfE4Riawsm
btps06/3wqtzU1SzBOhdIWa1AT1W5FD+TsiMzakkFAkqCAFMNhSj0vN4uxNwC5v4s0VIdV3MsA8+
eGAk0ED1E2GjTyaPMsEBHSVZ+TA+8OPgrW5OgdTUVcoWapB/1ZWvP8alQHb8bT1lXPTo+pIQx8Uy
4KnksTaVmUfJ0LWLxs+dcDg9WxDZpAjMZ0CV56T60eXb110tEzfJwLKFrnET/umn+yWwQxQkpRnS
i+u8FRyQKIFXo3sTNny3dkbm66ZKS8FsxB4u+XUVJAnnSyyIi0y7aKvtojKr6XSbVvLOpw309Lxw
UqAa8cOtRo19oCu6lQGfdD/Fa1CYY+QUhdfaciGXHz85GAKxECL/Wq7AHSlKQCPT2qUwi2/QPi26
hlBevqjRLMRE/M+zDv1Fy18QOeYeB+sWEtcjGRKgPGjB6luoAaV5+Bzp82dbYhLSzVIKUt8Dq5hz
ZEM5UytZ0CekE/x5IBzoBMi3cHJYSD9ZltEnKdW1czxX7tdDxRaX62mD33DKB0+RDbMU73rGn5bC
65cGw7rfgar/c/rdSp2Q7ex4DCsZtsiXrtQayJwycQ5r36VcdeH92jtscfjPGcEIPzrpI2k4X8Kv
fRd8b52o/ZZgBbB9sEdRpQfa1IvRfY70LX8TtIYZb21bJaWFsarB33IuXMMa8kzugS6NfAHroHA2
K0amHbA88oGDP2CUpwgK3Q/CWb0hck/xM7BXyAOWXp0hw9vR8jbEB8TRO7YbZv/YTWHz5sfMbPgE
zIkgwH87P/bNZyDq35Oxd2ZcnO/xsOzBim4VYGBfdf3hHaCO9V72VmZEclTxCV/NqeYZr533Bz0Y
PHjQFF+SYggpd+DYbtKVet/F+DcAOlgtGjeHx9k2NUFSNlS35R6hbxYI9mE8ZWH0CiBbZ/2a+Yt2
tDm+nleQH13lEgjlgzuuTdnk6rHup0OSOQ9MfMT8osQckzVALUBhfOfjU6Krno7WLzyFYA7y3EzW
6a5k1jUEAQAo4KCVBL0DO6+MjeQEZ17IRMFE1RoR/TeBnpiZJYxgjS8Rq/wZzIhFlJNfwty6Nics
FNVVCRQzpFF/jq5nTzB/6T+165X1GWDCliRddO/17+GJnBglKz6QrrdAlDo9wPsd0I0VAuNAqeZO
l7IzMafNaTCGQXTPB2SY1/4mejjusJYJNg/egiPksuhuF4C24s0bdzmPhZ7FPXxlpigT5F+eB27r
vemdRJA15q3R9ja9pblmcEQNzrHIXiA5Wxxagd52ihcskgeib2rRSdJ4mXalQqBS99yzAebT5H2b
2H590VJeq3d3yzsPAkawXAoWuM5CuDvZh0duqUkzJhAEukVF8/qJq1vpvQ6MvWSMBD3WxltMOarl
5qGI9PXTMRlJdC3XqzY8ymqLJEz24w0wopIaH1KXw2L/XUPrTT6hLg==
`pragma protect end_protected

// 
