/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbEJ1XVpuWmqpjnbJNvQMUK8+AJyFO5gGidGyA5iKLZ3IeJN+3FPx8DFs
XiHqdTTb3cOblPfmmTVNbjVCFENrLFEp/MiQf3eIfV5cA5oxGidSOyX8pO4zjhZCzmlJH9crLyvk
g2yFsg45VNmOHlKz8LQ3CZoux1Tcj9BaJrntSYFgBmXhNz/8jEvkcqr18BH4+EqJGTb8JWFLdsHL
pDyUT5kUxSrrgSSB3lvFIACltGz5Y4JmAvcXGYOQm+cVUYxnPN9aKbdClTiCu+3t2tgEQyUmfLg2
VhYeFrFS432Q4hKA8Fr6o/wcIg1C8y8VFupaCZygxUceFQP3AFDGNsB+hFaPW2O7A/Lg34URIVCs
B4nBX+vutOqgYHC6hzNLaa2pxSjB/ob0n4Ismzw5lfhHtz2DZQ5mr38o8LwumKmhfkc82jlOnxxd
BuF1VsE2VHqrVxlBuTu0yEydefDlAHLhogp14ubLh780I4nCBHxlDqRAdONrGWr+QHwLtwmsVVS3
4kgN9If0QQ9hYFmo/sn5+Zvbp6psFlYp7NuLiEDNYWkO2vFDQRDC7SP37w8Uxuz86+2wE+PGIn4K
BN58ztNToD8bwwtG3ESTmrCj2OEifuzQDHyouz7Z4kJsBQlXOoXH+y6fMT4razvvd4njXSqBq32T
Iu+3xvE9MPiJ1wutii4PIljDOyCjg/DCMrY+wxGB7Yx3RINcRURf4SRIGik2uMjq6BkXBOuqX7Es
qjpqTapbLRRGGpJ3VO8sKUAm0Y5xrWSUl3Vo/dP4WAyE7TTGzRtE6FEebrpO96l+IHP3Bzbn9wTX
lfFv+V5zdsXIvzbmKzQ0AWX3w7TIp1dlk25Gt0buiirbdlNtmgsaMDkuFi92BoFAFp4KoV78aOBt
WjW+Hy48wr1RoFqcsGM9nqZjyLafVa7P3F+dDV5H0Z0rMdxOobqhx/Q45XSaoYYodx21PwJsBkP4
k4plXTtkIM9NniWuuvd4mLkoJICqhL+iIZ2iWdr3rICswGczjU/7BdL+kOEVD3tycRBkS++6TyNJ
hckZYVrRxDGP+a+fsj/XYlSItwrE7eYaggn0HqKL/xiknRdVJ7+M3DAk+rCZmspbvIzvH1GfTQld
Gruc5mSlh+gjvS/FjIQElJ9nWzKgJz1srfNXOfXo+3G2BhoT8Gr75qTeRMSnjnIr2HcPUhIAEy8k
AVK1APa8sO5XlnXXnBC7HturL44Y6sFCiTy6R1TL13/o8WIsoi8VmNZIupT/pqFtwq84Bb6tim1l
6Dz0qfyTFGqA6XFsAQIj6flsZ/nui0Qbgspjo+LuVxPuwnisL1GZc1nxtu6r5NWJbXgKP208QtLR
0r1r7KpqL/8uBirtAuT46795ITYtSJ6eiqxjUKk7O+wkIv53TRyLAY+CPv//659Go6tKN134RpQV
PKfZtGNjIc0m4J1e9jd0bfPRudUPJfHHiXtolDiXop1b45cROTlsCOsDrY3L0Yvygv2KErGIy+/f
YY97hQOnC02uMC8xstPDbzhc9TR56XETr31a2rSs1bWHE3zf7l0xi+txIM0K3x2Ix8SGmFLOs9Nd
JYkPFRHl0RT1RltdToAS6323Xx3Vwkp08duvO/1tS1xHXP1JuC27D2JvThFJywDnSLEeF89RVS7P
OhLuPGzRyjZVpQntp7hBOgGSxu6IFb+JXKkP+9pr3KMqtHzEfSNnMkp7d9Og22AgJv/ZlTMvnnyv
BuDqe6OsRUUpIhXL3t6z6f+4r5aV7q0NPbvIvygyl09ks8uLWphSOKamZy6m9kTEW41Zqq+DJlnK
V2jEQc2eqlhZujU5Cw480TYuCeCSc0kKSxTUkg36fEBHrQzltVLY5hegAKPW8/9DvgsQ/94Fo+jg
fW0POyTXYmWLTlBr7i4jcx/vco9Pg4XJh0CfUjPmfMypZOH/oewW/Psb3IptwundxRRSo8du+UwS
mSYwVVAIaVa73TW9TaRPyGbkBctF7cnO9mIpBr2egDj18ObawwULsrSFhimTKTAy9rO0bW2xQfwr
XHcFxUaK8b1kR6oOm0gu5XuhwfGyZ7SQL7PFEYV1Tt5was0Kh+ruDTTkzPgmjiN3WZh782P9Nor9
h+tMaLIdPRSmkaO40VUfd/mbYeGrqgI+u5+Kr4FCdcXLpCScG2VTT/nd71j1/N4xpzoADBWcDplt
6k3UOHHIJ7Esf5PVu18zAckl9sPPqKxBt2MtLXXNo3OCTPB9kf4F71mKNEzUVyfaPacT/df2iZNO
eiAoIiLfl7TmKhJ1WZgPOzvM4XxYEBUbf+PvhqBqKwbU4925ptPyXlD/AiFbiY0XWWxq3xKZgxtt
1eUIQR5+5nfsF/ObMsxurcVWAOB3FN+xJi20NLMm0dmNSkmrpA9mZBjZ63jEg/Rwmt17AwIQ9MYx
oYEopMdQ4dncUPOLMbjoD8JQ06bhBdHVifpeaIfL/JzoTHhMhia+1XO2ClLP9YjbvrjZUiQvg2og
fGzWD63wZw8V1Mb2XAAlKMH4rUDMbhcy6PgbI3UjKnUKv/a7RIBBigY7/qheP88Ei/N0cDJ44sfL
0yROpPNDih52pBwvvFpVTLZelpudWA4LLtEU/eZBKu7zScPUVrf+odCGp/7FQWRid5msvT1HOmh9
TPNbse4LhXsgB4w0dSw3hUUEw+zciQSFn/OTJxPgalfx2LnpJaOaZ3+aDJlrRO1UY68vU9zPYFIP
pSTncLr17D929en/0X5AoorRKp0OoPJOsuO2wmuvxv+6GxFDvHTdzNCVNszpvYguyOF9bIFU41UN
1+wDsI1cauvkA6+hFGjm7FziN7r7VGF7b56ijska/HH7KcwzSANQEKxESmJ+jiheqyQAyPv77pLN
PtHDa5mIW21yNh12iGc8VjSCnZU3dE0/Q+LqjpT51WprI2zSnB60FpOV9OVAQCkpmgxgltRu8BmC
bHa1BLthnWG0ZoS6oQEu0g36H7ZE6VU/6mxRvN6GwQF9+yGNPYRJnQFkqYhVc3fe/8YXd+BS79md
1O6uHRH03GR9cx31WzI9aUH8NlTfwTtu1J4cIpdcDe4ZdMrjKH1SCTlWaidw2m5oHpdGoRFvI4KT
zXp0lQ7ZRyv2RBS3CeQt
`pragma protect end_protected

// 
