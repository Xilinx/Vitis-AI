/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1040)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPSzP41JMNuYnf6REKvs3Q2S6fyNZD46ajSZterAVqAPMpJn+AepeJpMOs
lOCiCMdeIiRybsKm9PVRzdxju5Aj1WkjBJcaOHeRtqOkhN5GgyYfXQPmUCzP2gXYfJkNxNa2gsdK
RAJJLAAWDwRe5Lt7iBffzZN7JJb5MjQ4dYWxsmVTUqegaLhGnAuVlcx/XMbb5W9RHPaccz4qFO7G
zGe1z1fJJyz8syAdyLC8Cjk6m4SV8AHCtsGhuBSVUJHvGW7a/Yymi46KHMaZAN7i5SSFEolKwFZV
bQTKzXFotkUy5nCeb2rTsIlLr7mdg3AeB+a8NVULWnwm8F7feAiMNQdFxIooLMFwXflMM32lSIFK
kJRdxd1heP49u5bEc8jx5ouGiR9jxQ4CS45StsPO7dZLCI18BpScs6yhawPJQhCB03dPlFvL7GYF
JX5bK2YlG3/CA6AEmVjKr+aGa674OSLa7cykRp4FZiR/rM8E0w8oRPD5zmpQGBrPW4R7giZI20Zf
ZRLhEykH0YHZaYpOKWzcYWlMY5VxFz8GaEKECiFwi7MBdJwCa+5b1tIkUy7+kt7gPvoMUDab4m45
psEThZe6eKbwLTSjD2B91OkisWVVuRCJlxSAyeQDVCzM7rrQ6wie9vmJnL4KA3lPx/my5tNBZHCg
PebUKSaAPHL3Nk6hknPRO53T1FfleKYEqbmF+j6kxZtO2995i+THHwYsAw6SG3ZEAUXbY/wRKAQB
oS/xqwT8/pQ0QfjBE6OOuKbLYsIPPQKshZ/FAumBhn009OHBb7zJie6tZPBfXHA0+iXikCzsSF8x
bH/FPCmfW/K92+0oJhMgtO+c4Qgopj0DFLrq6TBw884L0J/tgnu+FVuqhjjkBRvHiamWVYgzJn/D
zcOLF7Rmnq7ZiArrKrNND/89aubHp6f2JK1lGRkF/OpVAWhdVB7DwrSEQM3l+mIGnUHkA2ShGrJ5
P04O6ZUOGEUYpAeznj6a6QnZrnT9o6keYwL8sKbUaegQeW6PHNEYq+jc1Q4nLnbtRlHza0r4RpI6
V5XYJI/ejoWY0j33c9+BiysjF1jjnS1jBjYvhI+lGriBS5E0thjJk85p6XIGs4JQ0u64MsT+qrL7
c+Q7eRAVJtd903LFRmEMd3pz4J3AN8oqkOr+MGaFStCtZR2DBIsQrQACyoJEkC+Anl7FunBHcnMj
qsmsb6A0pBjv4pVjL1OR11fNmhqmCydSh6Z0ysyP/z1acRTg+Fnb70GJggUplfP1RAqf1w5ht8FG
yZCoufEbT+HEj9XvWSArocLatQfCH9vecxFFOjtxYFIQaHG49ylO+tk7nCfv7jGsLSyE2GIo2Rgp
giVEQXdw26CS9rILApM=
`pragma protect end_protected

// 
