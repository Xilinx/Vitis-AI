/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2mCpHp9D7qetJD3SkQXLNdz/T6lVtmZ7z1+wGRULTMAOIE1kaIyfl1FU
MAvEH+9JeyWXnx96+QYFVoFBT7SRlPOOVk9bjVTFav2lKqNEzItjt05JpFv/EnTcmIifpdY8ZWXI
c4ybjge81DJ0U61/gE2N4vG85FYzN7gQrmMnHH4Xd7XwvBAxU/swN8ODFiCcpcJnVDPSPaYWGAE+
qRo/CKbiWbsfdIOEytqSZI0Lb1iZUdW0GsF0qkYvY/ymkejuuCuHPgeTure5P8VNFDaqnb3Ts4bJ
3txGtgf8Nl+I4RkUBqOe3arCVQUYIIxHnGMbdYTEsFbNsoD9EA8AkLjGJ6ax4hH3ZWXc2p7OQ6mK
4QN0kP+6FFMVfc0pX6zHrKWneAhxytc1nLZfm0uRN3dbquaaia8jias6En6UIEaGja1hwQM6QZ1C
rM8YmY7lu2YEatTaQplVMQnJ8k8D9hyX0rPP+UjCHNcfPvKuH+39NYmEZ4BzM8LHeRnjtGSlmEvq
SHzEUyaq38jgyxGDrmv42Jv52Ee94QhjIQTAwI482KbIIYQfwRu81HC81BkaO+W1ceQYuS/moxR6
zuDMeaPUpqRCet1s5Ih5o7zZuJdSKff8Xin2np2uYOgPHcP3+z06ngwLVOhFiWLbSmeTaZBdJ4oL
78a1AQjzjeTTpAJnlhH8Pr6fsi0ebynzPzU9VpIIGtq1l5+XaRDfGtxvfazsIvK9K9GiNSa44gF9
wfx6EkupRLezUjYdy721NSmXHMFycxcqOflp5dEnWCsenfwLiRUHOQGBheMkL7qakQG+LxRV+4/W
eY6erVkUX1I3K2gFz4Gdhrg3+bI51KQyXUxVGtbQe5WqdbpoTcEwqCRZrN+NhOpr2dwXiHBNTMu6
ixd/nz3qwvhci3wpS38ow10nBG22N/q+15mqza3QlF4+sebuLiMRr05xDlOOAApzCEveu+KvSQrl
HWJIH+fN7mb/eeF2iHeBrSYMJ82LKKMJBvdfk4baymWXTclxvO6N5OOE446HgpKqJj3tLGlbb6Wh
rHvjd2FAZ5sKNB8hgT+jwUwCfIiGh2bOQNXOx4CBjyB9qRKiTuM2ByCFK8AaVHZ/AA8w21NDj08t
YYgOVPDdT4Kfr6MOV0SVued2IUUE3+Pnuijxc4ioGGQqwWpyQIZNe0jw/Fvx6hbKx92bxR5L/2OR
jYxTNMoVetRi/Ufbst+az8z2oF+bG53iNXwvzc2Yo6deGT/2C7CeAOdug+x6gv8v9eXkiUvQ3k+p
IqyA18ks0NDeF4OyRf6wOr/nYn6E9LhphU9J8iUKQCkvophmfAkmIROee8rCJbNgS6JX7o/cnQcP
r4JwCrD5hSm3+BmnZiludHYlV8Z8PgKc2nBAH7AB3mSJaKqTqz3+KOvRDQ7vfJEc+6A+7kD+EzKk
eS2wnOpBqNx//acA1DROIEIlJf0XQOdfMIt8S8LNn1QU7XFh2IAbDls7iIviBdy+oIuUqsRqOOVD
AQL8HBGxrw0Bm8aaShgBoEDY1jwoWLNhYTPKCQODHLvQmQ7DWlNeQ4ybA60bOfcwtxfMxs7F5+Yx
ypGwOTzpzILwiVgnxMM1KmTl5KpLDTBJ+WNqIJ9Xk4rriAl+whAGxsWPtwc6Y93ajGAVW68r/gIN
FY7gJAuW867TG+CN1bUuMnDgxK59nnz6BSuxE8SR2p9dow0WBJCOGs6MOX4MK6jBTw+ZNBjRyc5V
IOa93N3kmpAp/LyASXt5+zh3+UjhNVtlY5NzrrBmY1IVymfYj6/Ii+0KhojPSI4Ktrp3Cu/HELTA
VYRv3xi9VaN5TkjKHAgkITBvREruZKMVjYpVOOi9c22I2XN9aGm5YuQTm5mZolTHm1fqh6s5pzlt
mdipXUrf6Q0iz66BOSERbTcGTt243i9iEaT1Ga0/UwrM01wxLAAJtzTrd7dvNBoBTuggL2Q/gqp6
NGi6rjYb1kEQI5ut373RvYPp3KW9e1eRxJNvBsG8hbbWtRPJmy+ut5eh03tR7VCz7lb2P6ItL+28
2o6rMZBWPDbxnB88mVwzZXVMDaTOE7VnHWrvwxMaVsn5cND7Xu47JS2C5Bpt6I+OCYCOJg+LVCw+
tNwbx1rvhdjoIqlOvWq68WcnTOHD9fmaBFdk5Zcz02auGYHp0nzuK9tRvGOiAx8l5HSASmCXi7R6
E3lZ6LrB8hC+C32r0OX0l8UTA1Y/rf7Xcpwg+lPFcHNvYd5UbCgTLyCGWodZYeQDtSTwafCRByS7
o0Ks0Nki4z9cj+quobgeEGB1rpEOfPI0BQHsCSFUpGyTKepgw7Ef79Q+5pWZ12a2bVKJykR34fxC
7w7rVb313CeB1UuAA957XQEgGLXxbT2Na9NnXseHG9b+iroSsdVY1Tl5m5AhNQ8345VXd0Gp1LQm
88TUVoh8yRlwJSaHHB6/jnniZCUhrknFFD/yGNUAZb4Xh2XAufN3285jJrbLIGIbOyr8Zrey+6Q0
uUsgmrMV+Mht6axlv+fEaIEavWx++XvgXGse6JomsHaDeqrKwOkBZqKFO4CxRxB7qQJ4PZvNT0hn
FZrf+3T96b062u5n8GHiYG4z7WVhhZL5+OMCCiEsdKPIfzSffeZyiDGMXwlUUF4s7BfdDaYgl+Ah
87Cj8vVdDdrAHQkMbryKmEfx5Ti9zDxHfPOcAF5gLH0a9yGy2wyMDQD5kw7OZKh3azXTDvi2Jhdf
ImOzkLesHLyw8yUnf5PVO06ae+PSFIzNXOWYMbH4wvRodHAlq2KwFHjX8hhph1u52XP+ewYNuhJP
ys+aooh38c/DpB0g7U7Xg6AM2akXqLlm29ky0bJ4hj1UEfXtCOw82T/SGDGsdw7QMIQl6mozLt7+
wsqF80CVtW1eggqVH3GcR5sMPR8uWP/apguXH7Ol160HVi8hv8bvrhLo6tRqYXoGtsnl3LqS1x7A
6APBefR+/+iYlF5wLp1aapTj0g7S+UtSen6a9QGZWrie/6UWrCt+PCfXAbiPBzYP7yM9IACkmTc9
5V3+ovTPBdRu8B5PG9c1g6fgoQ8V3jtJ0mj+pkhWjDEjsKbTM2pjo0BcwF/Pa4vG6iqneYpfXNZZ
YTalaI5GhdhmTJwW9Fs7
`pragma protect end_protected

// 
