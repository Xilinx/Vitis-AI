`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22064)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPak/iHwVkUKXxdtqF6qlW2P9HJ89gT4zeosXKnzybBKQialRE7ur2A+8kSh4RLXhMpjk4PSF
wuVi3EhccpgeSY0nh2L1fj2IxO1gkt7rPYXKExhEw05T1zqKQwsESNr7u0KJnHXBGJeIwnaXrP85
EloNbh98kjIuZL9kACQTly+za15Z7uOxzuWSYJyJXayUfLzRZsvZTlUnnZX8e19MoNjdpKHW20yN
OQFdn3pQf+QnEIef/4ZgFIHF5o5UHieylEfeSBJvQdGYXs+9fIj3UG9DmIs/qLoKVZjXX/MyoX1W
nEagwxyKf8q0dFKN5XY+N3PhBtKjCFQHZ58Rcts9L0uvqJA86HMmJnCzNobTSfNphsAqAIJXYCX+
DX7V8n3xu5GkS70v3NPukfzgLqGzopnS1nE8Yky8imYqHggnDzjF/qyCf+OSPhZgqbUjMLEMPHSZ
WRWhRhDCzv7dfD0DDzNRgjp4Ql1ueTpxN9Ca0QLRfplQu4ETyZRib8vdQZy3Wk4PJMPpKpMiySwM
eYa/TxLYGNJlYpMAIITGbzjEv0AUzpLV1u3RS8qeDeUWx1vfxJOMsSgKOodk23vxjeiBSH/zr2FH
d94nmW4mB8AwXSck+aYSNkBE4ajMXBYGrYyPWBkZnOc4Pn9mcP8Kf0DmMC9+mwmfUlXGywrEI5m5
I0YqdI93DSnSjkeR33OnAXRB+WGkYzXip+lM3wWByxFJecvwHb543tSqshwbZ/c2MzlJQ5LRXr4x
9YYuj5tGU4CsLJu/YFE+Nsprf+o08xIyXcZfwVEUmdgMHBl3LJcckE+SpGXaiKbRPp5KnnQxr194
QLCMXO283xAB4AmXf3GHZAKZza933nJlBLkIwo/P2s+aisG5POTL691/2uz0yvTjCH/rEbyj0H45
1VZMmS4qRHfqm1jj6MUw+hOdUTgCz1unk5Pix0UMDc378uaNwYEv8GdG/5Pbw6rHVoJc3RRZHoBH
lswdBc+S9nOgyk1qLCS20EXS20uOHGhbOlvDINWOknVmUQETYNZK96spUNXjDv/d1ceEqyXfDkHO
ZxMNS7TWqhYu71wLwi0t4edXyQcvkT1hQVn0pbPi6bK+hGnq5ahA4H8IqbpV/nhzrELeXvqPs4p1
3wI14m1Vybd6KsLQmLAWtyFJB8ea/7HK0cZfXzFxd4T9Dr579oHlEHjiIOFUz++/YXo+f+OLHNZL
UrKF1aBgpz7MH3wuutWmUCRBnh3/AvufabKy5WOghySm3rrfMCn5TnetMjvNFv2p+lNqSsO8fgmH
lJTElPndop/9EXUHhBxB4vUPlEcqVopQ9ULDlW1Bkra3rWzNLNlFwpUfUaUNFA0vIwlL9LNe39jl
tN0ut/GnzatbONNWH8eE1S1ZwEeuMIZMLzNKTIp5Mzd1/9G7CoH5MVhlcJk/qT1gBKcBxEnzVdbt
eNWYl30TwFBM6V5RUI8a6i44/rsO8YBODfBZTf0c7qCwrhkzAL/yajgYg5WxJw1Is1vmETfO1gGa
kvmWasoMRTWbKTNCBcbJcTxtnGEykBWVWI2fedmDeCThPipUSsqO4Ze05TE84VTECuuvXiPs2RfG
jz6ojUC7Dql8LemOxq6q6jkg30hPtN2P9LESfv4DfETA4wp/YhZpd40YNoZhvN+eza/B6Mkq8uCl
KoZHN2s58Sgq9YB0l2H/WrGDyR/G8eAdNvXK+v72p4IpCX8SbQvCMzhMHeZ8FbfGArLdU11Nqhxr
Y+abHAaWFvKKy7OlaBr0tbaCMz+TO+eEpjpGNBa4MSSLL7lE4pmsxt+d23j34VBIVZTiZH6xxpYE
hd0T22fv2N8E9o7braiV2JvK54vCfgd3DDvbGiSXrRzH+t5929cEltq1+b7c54we5G1GbU8+4r5f
PWdpGI52mpCkwagFwT2FNJTRNsVJJ6f7n6OIOA2YoERbPpre1XiU9Fr2rz98iAA6y7IhfjiJIzvu
Qfe7f+AhcrRnTQqfQVqVdsuMzdzRt1khKZf+w7sopdqKGi6tNEY50yN5pQ+EuEVt9HDHREOrFr1p
Fr0bzEtXurp2/rvyU4eCwa5uuEbCRGj7CtCB5jjh9IT/sNL8YB56uiYt88WP5tQaibq630WWhgXS
qeKI0qDAfR7DvQo+Tvh2fEUaavjybFBENgpvy/NGdgHpOama++p1GuoI3JSAaGhB4g+1sCU7Lxjn
mLnrZ5YNWUM9VU8DBk9b3UG2h0MYtmYNn0ONimws/ndgY7Rh2oFkjRBlKtGx3/C9TTWVFjmOAsTv
KFH7lYniaheqqiJoySqymeH87B5OkfSsdp+Pl+HenPToIlotIDbiNQp1xQOYM01ybcdgKrtgIh9A
wQRL/WSObxff2qn+Ze5cYusaf6gawsEoBYYnC2VS1OJ7HZ2YSAirX89l2fUntLKQtVtxP/JUL5wN
gxo9ztu5FEOlHLX/a5LaDJX6beaygmJV3T1ussPG+otx3kS23VgRw9BefZHTfgkEaV3f4ghoPyj9
RDY3KUBAjYsPeoxqLYCHu8TAjN3yWt+ZO47E9q8SFqgnGNbbEmxJafUCDChskPzY38NdnnXUNFmi
WTr6jifBE/f0Va9WS24nwaHPI83+loD6/Q6N3waDDsIhtLVynrPs0veG4CNZKfSOSQkbEtuWxIp2
ugCY8TaRQX5ubjkJEZ5N6d2X/a5kta7H/ieydHvUhcqp2Olj5RUBVoZs7Rv2cLJbAzAkZZjdlI7c
Up6iy2+SMpZPCjdxr2q9VVDcgALtUcJ2+Rnt+ON5Hi1kapFclhNxz3LGLu3chjZiOW7xZjDIhjfE
dPKtEGDJdJwpLQciwAhcdMkmTZSfjZVCSLB8nOWgjJjWCP6WE4C6OeMdpgiNP1e2Dk2XwLhfuPxA
ad0NUPcZwWFqIDzHX5ImKA0u+7LF/fTFaHSE+kDJZcSnYYP2P/4pmMSm4IpJJGU5JEUVhwZXXPto
cxhvIK67Igd8YnNWWRmoaSyLoKYwuvDtA/hOg3LSWbePgbQBgUDONomGPwR5SaG3xG7AM+pDAWuD
DmZRTczRcYTvlSQrzCSRCaMwARP1/gCe1+31uvJJtH5jWc24STtPgmKc+vv/KDMMNQK6dRJ+shwl
OfQv/TNPTtfpKe/sL2snFvHsSZyH6wSP+Z4W62RdCROqa18w9+1rt5hTd7BeGohYXHy/eO/lYxJd
tOVkiMm55chEdKRsmpqXRT74vuZ7Hxwr+/4NMPGp53XhFfx4kPEyzOofDuem2+Zh2my4ePc/NSeH
VO25b9IDg4dP7x0odchfhQqw07wIXlH0+Gh2wzs12sVC44zuKC5bZ8U7KdpQp4do18fvm3tSZMw8
lOIc8f8mK+uHGbiQJIg1peKsn3IAN/6AUKrIMJYrf3/NN6n7/W26zaZS54ZFB8cEUM5VFzSyRTk4
hpStGuE83IiapQyprGeiORIjUjejedFlOmYnHmSaH+sZWFw329AIcs3BTxngXd5k1Fjisyw9o7pd
UpNiBK7sgQnVQA0k6Fhe8n3H3Wa+imAFdpCBGZWKDokmPjLXYp09N/iusEbKeyrYCqu7xAxNn7Aq
7OvTmCeJ1hDv2fYQDEC7WVBNnTrGMaqkj+kjoL5lX6L4S8axFY6IrBn9tkMCPgjWBTJUDDzPReFW
V4xyi7sIIMJcx7sRQIGNvPxLI+e+M7t7drPdiFoSVk8bToK6tf9DjtnQYCwwDz+386OOc2VdReW3
iNvMRk7GS0RANqqNvFCBNFugvqJfz3SrsPtyegOj275oPcrVHdCAu6dRmPU1Gp/FYTZo+bSd6s7g
8fQowsrVCyNFeqIVkK2FuRgU4c4a18sy1IEdl+6tU0WGf4r4+Es7KoAIjsDdeJDHdDXBNJShsMMg
Vv//4Vyo6InoDqQV+rJYMzBndQ6ZV93v19sdWrMO4nuuaW7mbtgEDdG/25rytNwdg+jKFZt2xpa9
nQu69F1zlQ2s8j6H80WX+ExEbwkpsF8KxlzP+FJ9R+b/IQeV3DhUcM3q1YtJngC4gdjdgsmKButJ
VDaFjA02R9qUDT+D2KQrPbOyE2+UvnFjb4VhQG7mU1sPT4mcvYddMoZ/jUXjz2OLvLns/GJwo84b
YOVW3vb0CKBzkC9gdcuz47Ysw6IgWYpShSkE4aRLibkmsewSSJyD1E1YhKnuj6nsRDpP4UwGdlQX
+L/rdY/7Kn6wnvh6/PgivkDNebErQQV0GS7Ja/Gs7hLMBqtkOp14uIMir17on0QwLWRG/IT1QwIl
Y8vi5x39OIk1d+qAlYfRXGIPJKCNpXkH9amk2e4CGs70a5QKrio3pgvv0DZLtkdaxNyngabZ823w
F3SDR9KXZwdoooif7I0CwGgvZy6wUp1LZBNM73evpPgDRvAIwQHy/xoNxNorrqYUl2bUlB50FP0a
l5zRiVHBmZtPKSpbf2KwO8EwaM4cjqfsgnftBasK306JAVo3+MlkTeKuojNzTUHt6/X2qmsP4cx/
9I8eN7nrtJDYSVyEwRlfhWTedYMWc2VMCnVFPEzHgthPS4yGj5grUNzFKKZH1AI8U5Y5Wu4Jgx0G
ZvXvYmaXlyr2huIKztytUQaS2qC0xzhlj3YVLJc0qz9SwcYzqMp703hf+WdGnBc63kCHsRN3hT9a
D4I3Ai0ekH00+qqjkz6cW/ktD/UJGocANKjrZ3cNUHmTtXPrPwtcUGlm3gkD+8pw2txcX6qq/V5V
PeBpejfODfGelWQs1Y3IZ+gKZGZNl/O2TWpqFTrb0rG2JpsDHq/JyRLUNHx/dRwyIz1E1YRCZBkg
Z+8ttbYoZeQuvHYpU7PMon67gzCMQ60blRI5gB52o7qcHxQjvxz+3eRFYtZ/kQNYtvUQpjbxXcKt
6nWEfwzJkTVtdxQNg1ouNclmy5NStr+golo/SstZS75cWgvhp8hioNQofb+bWlGN8pooh1kaFVBO
NNyfuSjlZo4/fV9dhgRpjFyEHxcmD61aqzOqA8ZRIqVOaVbYOlOX6UnyyyX2JjxM3GxAtFkDKrdr
soDycNUVo4ZMN+fd3O9kRpa3nuvaAVP2rpmu2vtRGsEguXAT+kx8y2ZV8VgtqpyfH7YVhmmppnWq
L4E3a30noiIAYJoNYvmIbPKjdnDc+wzv2D7+3vD+lxDc/F1b9kcCa97JZ9vTnz3EuFlnOM2o4Lir
moC7c/N1M1o412SOBoyAs6WQhkcwWfWvCyxYsCtR2zlq4aPDlxHmp3TR7HUVdOl0NNxxr3wPsdtb
osLe8f//XOCXmQ26GLDdNuffgBOz/aq3v7LdKtH5wD+nS5Usv/ZXDoetkteZXTro5akajIcydhfR
9bqOAGejXsUQsmj7Jd6GEZBVEtZPnR0Tm228Y3z5uXEelVMN2zCf5Z42jwfWhbsXYrP88KyHqr3e
xWMiTHRiaViYQp2psVbnfNfrcFb0h7PbNyoPUL4qp/Xtu4NAch09JlcaSFNpv/+zCQXVOMx1Q6nj
Hd87r8ID6NXqcYn+t+e7JlOWb87g3t+TyneuNHifKitYw9huNwEfLwrhbMA0RZA657LPPVpX9J3H
ArfJZabKXMRxqsuL0yqbbKzBEULs01ZTqDpUddIZ4nDxI4RUIZikOUqwZqeNv32DAu6jB4sRyf92
4vbHdrsRZi3m3EsNg7yFtVfTuKkMju+0afdvEkPPrNaI/+BaAhkq9aLggv+q3BD272ExNvJiPVD4
SBfwjfRBkhhAAyj7UHcBVRprwTw1LJRer5aS/goUFMi513c/U3G7b2wW29RVdDF/txMgERGO79LH
+jX6rqSb8GNYVhYR/iNhgCTsCVqOi+t+flpsw1Y/H6ln5OQ3WolF+cXBkNRVPP+jxJixvhu16J0k
qvWXXx2eJPp2dPf4jnWHVy9w8gTBJtQczlPrX9YQ/cMvv+yOJt7VedQS6VCrgcCpXi2a4mKEcW51
KmLvmR9lJHSVQ6FEWFHMsBR1ODoop+XRrsqMv0OvJnQHBwgaNiBS5hROvrj0jDJo/0zrF+9QvcZH
UBmNUmeWBktM3ByCr/ajDuX3ED46SJLGlpH06ZjZs2rIwLoG1nWd6G+i4t4/oJE2FsJrH9zoLHbW
r6D1PP8/9XH3ZatPvyCYCk1SgTrxPBUIN0bdp2LHpig4c9OaTHRscII0xf0xQGKBPsckkyZHLprs
7nvSxAxJ8MURm7usQVjD+DkySeBi8zeHr3XS75aGrTsyHRgXmQo5yHwY45SahtN98iWjI1v+iQAH
mcTfQ+un8aC1xpJU/INWnhrNEXeCPLSDI0bs2hGb9X/c4IDQ2FMf1iYHu4IK829dwNdjvAjQhcHb
6W8KpztvLnC29gVZohn38sSyYk33DlsUYnlgzA8ps+vFgig2Bro9/ideX0YyDkHL1F04jR+YUtmY
3+L8OaZDNjSxEwA/wm26tcV1IcUvoicAjPg48ww0tw1PXrMQ1hx1SWrpCJ1QzlaW0qprb0V8C0qt
P8TbTqx8u4Y3ATTiSp9Zsu1IfOlAQiWgT0OkxpA5SMmcUOtlcJIwViJEXSyg6QZu2Ws7fJDDXXZf
2jK9yzh/Inf+HX/Xh2ksugymgTgrp3dMVkC1ZJdEhFSYf3JxUp93LcaQpdJkL/z1P2o8/PbfQ7M4
zUwsI+hDWn0LPArr3f10J4L6r8wFJoyXC7uKvZ5hMKlpws7KH/C/YXw3M44sh5qW1hGGr7MzezXz
p/iE4Tzs/TdRAb+nO59/24qoMm3NfE27jfLbuYkAhQeSZPp5qDB7ILt2pIbDOZcCZ1GZWjfu5SST
ksRuY3xNimgYRBAZI01gaMOuCwYuA2MvOLg1G01YADA54xRhTptjLjDP/u0nS9T4t+nxP4qUB+qn
DWZv8bq5OTwA54IJcQpceM7MJzNOhjW7tI1vwMiKrCvWOzcNAVxlzZdIm74nmla0p7i5Siz3wj0h
u8GenXuYW/Su0qrnfJBz2xmBGjyPxycgRI8X2fzmwYg/lNExYlUoUyk2BI+EaKvwZk8s4Ycr+X0g
Ijo2S3XZkNsk1P1c4OUAnGYrkgwq+nuCjHNdN0iDs86gbTZdYYXtwFbiA92mD+eTkhzH7pg2rjTL
s8MdBK0Ad771NUSNJMs4YbakEKUUZboeLmq/Hy2aM8CNiSzNwTadA8Tr2fzLZohz3GhX95flmW3f
0hEnZjMyIknb29PJrTKjNBLRPBpnjaEbSGnOb578j2Bb3/ExTp2m+NltGEOcllbEai2YB5IA0go0
XcsBwtkvZF8q869DIyJEQRKzEVhVM8P1TA8TwnR6Ls9qtCo7zsyK3rzv4Feq+OOU3DDr95s+9dP0
JNi0HxxESN/ftRh1npM/HwDpUE1qfQDlLqlWls2FL8M+8YbYrDkUV2jwnFsmn7gfpsHrnxA3Enpd
GmLm9QZBR259dzDVSTkLhoZjcqyuuvQqLrRATdFIfZGIcK/4nt8BPQ5AGJqjnZG1F4cdZ3LiZEAT
lPyUqXUUecBEJCNWw/e+Ijm8kOqtWjlf4WLptwBzaZLgSYTVF5O+9tk1/0GYgFKkVzmXaucqLbns
ahkCLtiBp1mFjty2KUqPxELUIaXa31Tc6+D0N1CN9xfVytsgiJ6SwIexUHbDq/CtLW5SODJ1SdaA
uLTmVzI7H+hiZOEqdnQTEiaU8AjVLoNGN9YYH/XfQFZ1uPQRt9Id0InNE37Np8u477NwM4PndrVi
XjPukw8cIcdEBq9JAqjkgoX9VWlHWTvsLmIXEP7UpiMN5+ybW8tghRpabpPk1/j6idK/0zbNGHDi
KTxxAEjWuXQCL0uZL64fnPmqIUVecBWfHvpHZCUKl/uzXGjMSMnx/asvA5uCAu6eHAc2zRTFqZZ/
13Xjx+kflMkWbVT5OcFfpI/y9kiSUnht967Fn+5ZOP9VkNuB0AS8kEA98qAdG+72GK5NiBl+ZKEW
ZlrR1UYdG600ylLPJXIiRgFC85X+cjZ/LzZqVOz7hx7CXIjfqCegHmVSt5ilB7J41cAfPExiFDez
2paTzz4Eo5DZrdAY2Xj5zzjObV4c05LSoJ8XUyQGPp/CknCmv3CxDSzYLqQSE/NF/qJb7ZONV/7h
IwSSF9k7D3UEvHqig/EX2jVHT/0qGLRbwf5n/3rNe7ckxfHfljT6Vj3hqdFKW7wscLPhsAtrn39n
7HhvfEKvztMVgHwe+8/XzUOeyePRDEe+7qFWynos5N9K64X4P7PgFq321poz3NH1jvbYHJ+IxTNU
j7mXpX4AegDNGRST0fVMn6jCHonQ2mdPvPAFRpP2BckGnhqmZw0vLdV1CAblaaZgDNMkifSEH3Dq
wS7/5QplX6W2VzV85rLAtwpSza5ue+6mwjGozAz4XiqeRLGQXTt1F8M8fjPKEVd0HoALj9pfn6rR
PHlVRLwlNWvQ0/7nIykUYzB4lbK7MGmN8j3SElx4aFpP+l4Ke7DKwu29cN6Om3365oFDigxUF9en
dXc5BS1+YYpTbgDHYptHroif5MR+vN7e9xWkO4G6eBDsxKh2iDyK/+yXqGR3ACLRUFlgrSuYVzW6
WMFyEpV00jvhTXOC60MUe3zwcLG0d9PRze2Y4Dyiucd994+DxBq1494xUWF1tNFBz6QKcU638yt6
/VKVMR1IdHbN8rFcBi8yuWpKK05oEXQ5rV2P+rRTMko7vqKwfvBFIi0zAMMYfVKlycrIjYKySF0t
AEZnNQPuj/0qMtbcQUHxvewDzh1gimVVCElwQNtygY4TiWpgLl9DQynAnDrYKjRyrSYRO2ow6BRb
B6/biPAXnMftLlOefnyrl5xWuNp6SIqpujDvJfJwCt70rs9DVW4dCsYtz97vsUFa+Fszs37DC+xL
k9sRDHgNM90Ser3Xg66ApjpA+vO/C1nkAJqu8jCLAF/Lm8+m5BDGC158EKUCdlVOwOVPWi1YSaJR
kk11M7L6iCSkcmRbpweJwEDNIWH5HOefsUHKNq1++Q8Jp5XNnJ7z+aRAf688jqJtgRUOCDu4h9Qk
UZTx6Ela6Tb6TLGSsz/NSQm5zOzSn+cQi6w7c2sErD440d2M4iNDIlYBQbuEKCVjAIGbJ84K9vaE
3+ZadIKyORd20TE2F1AoOwrQGrpk+NBNDdJF+kOJmMTFreM7rvivTxTi7HzctCDmNlw+baUlW3WU
1tYFmEW3MmzIvo+4X1Fi/xutKjAdWf/OKTNFzI9a3hep8H3XtNzvJw6XwoB9D49nBLUKvAYd3Uan
u3qYnpdDCCuhANRvOJU/3Uo/8fkiXAuX62Lhn2WyR3KrIx8fcxiTqBbRTO9QjlVUucKbBku5nZBv
TXKKhdGBkhqytmO0TuqKi6vaU00olEyDK0Vq2rF6dnqGwz2f/MQfuvIsXo0Mzfm+2mrOQE3+k5Qj
h6Zp/dFz4n5Ni/oW9gG04OuGm/WVdp+G565kN//WZ7ZZrla4Nqv8ZpDF/sEz/D7w0IqwlxM+W4gv
Xkg84teqLTv+/RNmDhsqnjF9q7dijwS0Triohry6pE5RUW0llu5yTdyjYs0D3d6N0/hyW8pkm/lN
qtYWpQLSwHz3JKYOtGESqutc9o1+y3/YIKGOwoAmE3+dyuCQFOrqd0O9jbpag06a+gG/JOl0cvPz
0FiZCO1JaeEjLrZYDA3QaAvR7/NzEVsfnwukLVFcenx4q4IU9FNoomRxsQJEgCmPHZrMUZpi0hr5
V5CIBPl9rG2eONcXIfNXmk2qNJQg0xKYStKpnCZStz6lz9fSUEFs2HBIevKizWXH/jRVBcqxNWpa
i/vu+RXobf5xe/Fjo17zNsSjTr7UxvGS+gSTIN4YU6yLYYu/kKRaPcdv571vggkzDAZ42e/oqwFD
QmvbsoHzF0ZrS6Wvus9gNvNtLWf1kJu1/Vu71ow0NZzjjZj0kzaNipgAs0VciMxRPZdH62wg2wA1
jJaXEwCY6x1IdSuPl6d1tIPJJyPCwqCp21IbAMYd8oazvZD0pFHJW7+MH2fW6L9g0sW/IV0tbIaO
7hFpOlAoDiDA2pZfcAa/CSNZ8vpXEtDkb3xbAVCgfabb1SP5PrH7w7l1vFOp8VoEjIFufgHzGLE/
5LwnGvHBnyln18Ba16YyiPttcmI1QgkPN+tLrfcDAemwK98WGcs6of8Zrily9SsFVdihVKVFbjrt
KaNXYYaq/j4j3oktPhU5k1wKupNnnxO+btvgbJGi2T8ZNfebDx3OpML9I4NTRNkTlhFLZ7NJDygQ
NRBmV3EOZl8T0I+bUO0ES/MaSiEiP8rAkVTwa/3BcBmYud+YRB6WFPUPjdGbk8qfMbTcMAFXp5EK
J7zL2G1c2YXmrytIQlPTLoD0vFhUGiRIbZBS86hpmLWTM718yh3hAAGQ+zJzWbtcR1tPXN0KjamQ
ipBAeYBwe8unZ+WLWfSoOVVbVCoaSbACgXMoz6jVjGSbTPxdsnTeUlKM+5Ql14y6yglpx95An+k+
/7V/8oSV4bqlvqKjOaQjj4lg/p2s2eFgyRfDgWNRmTkAqC4p77rj9fFW8s/DzmmUsIO9rtA5ZUf0
h3p4sBSZ68FiaLRAtplt2MTaVfN+vr0vjVMnUF50bHyklQ32zkA9iVkycs3WBRrjoUvvtH/IBUNg
AbQoXX6EPUkUcYkwXOX8Y/J3KJBHsSIGuNLl88altJ9JxrChvarwU+P2tz+bVL8qajZ90fbGF4Ul
pZs4/nlRV12VH8R2HSZCa+er7mgZrnkEYGS+UazecdRJZrLSm/+NUuoR4e9uHosqxCwaxPGkxM89
PFn1CVkVQ8D4fJ8ZamhS+2e7K8+kiMCXNkIO7dZU8PuBtPB2/U6W/Vja+9Ir5BcfrTLVDNlrKOmw
VCFHSTsqQrPH0tOs3Jr0RLSXLuELiFbw21yIYyCJAqS4gY+MQxkQfVj6fkqkhuPa4zNH4pBUK5jW
xvnLko7Z1MkQd+AQ3uvMnwa5sppN0DsiPDYcVM/T6IEk4AyEEcLHDyjLgePDfQneA5qOx0H/C9z6
8xPY6/PBaHmPjtg3zecHDGa84sCWE5QjKQOPb55DSHvn9ANhuCRpYRS6oNRxxdOO6e8dAaha7A73
4GNQtsnYvJ55VuC93lSfbVtod4w4XEY2SQ/dfhsFGVyIe4YepXl0TWQdEDzW+c3acTuCTBa2AT3g
+ADDf68kV3pe1ZBXzRQ/TpHpp1AL6YzfVyYTjw3UJ1uig2/N0B6gEKMS8u1odG5sKoTvmpuaGkgb
A2dSQ5sv1wrSNzZf8YqBVCXkHn65n1eo7cuqt7EiJSyC8g2pzqW1Vh62Au86+aJuwDces4AGyWgZ
b0u3pAmnyP2WxqxpPoqyT2pf/Ov+QqPUIIhx8X7O3KywXUdtJigsNoQfcyT3vmZfAsAAmc7Mse0/
RBwZ9LJnYR5e6LzS04NRukkX/1UC+4cwrEc738RXeTyF4RXfPBo2hVydOCwDH+tLbgHeQdrE/Av9
84pnyBTUtTcQcoxWXijbq0NPofKXUc6YVOYy4HBKLi60nFbASxRjulythamKD3Bf/oDC2mH19I0T
miVDciyix1RUJ+HCd3XtoPyL2HFVBdrVEfrWW8bzRKdLGti39kSuZmLOhGot27OuWIXXrZ1AYwWV
M5zQiBUZXOlo1bdKuRulkK1mO+tiEIapYsyFeWhHLmqyxs60kcuIUaCSOSmZWj+wE7a1BuxOQvJq
eqBfSaJQn6LMRkimLabc+hJ0Q7GPNuSgdTQW+04TJBCRjkOL+trOmLHblPX3apGwaEi+w06IMRNx
0V32OsDvrg/dKsG8kKnrTdBSOoJTS7zF1wYr4/jBX+wV2+zOVr+BPSf7Jnlf4e2tHX9P4/W0fUtD
+MrtLrYw8HeaQYysGrucvNfpz1wojvtsrLUN8F/MrmRy3SqT8Opj9aLnMuqndulkyyD7Ur2OtyUQ
Gd62ZdGmhJXSHEpYWFYmF3MA5Vyj7KJa/C+7Y6ZVwjPSOLEFL3E8VjUNmKKQUhwEAb3s2O7q7gzo
IU4oeR36G3eOErPYYtU729mUPdVf9WQRQAXoNdJpx4udP9NgCeoK9UQi8Xp1yiYjOFDEbtKA7Hmu
Nw10gBtZGF0Zl435+JzpkjZkI4Kn0von+JF1C9mUlo+PmpfWfer6bdMKlQUnJAezsPpxnc64hZVq
u6fug8s8js6PtmdUOXTKzGgkWPqGCoH15uNnUzmgIJzBdNqJEWzG1O/YF5ox6MlTcQZzdFHC2AHm
YOGr6CjdeFdpLd+s4bSv+uSoWQPD6HTadz1AnNdCOQ9WExQUDoABlnQVB3Go1f4REvRIqH5U4bbQ
/cGUm9iJzs8XUeywuXTvFYkXkQRchWC/dEvAWFB72c5XqdgOXAt7lvoPNeoKmM00VbNOxENF/Ap0
0qm6Qr7W0sXD4k9DXR1sHKzbJ48Sp04HWVBbb4pDgRoLnUJCThV1TvrmkVg/ybBRgvp+7uDKWuMe
TO/yxbmKFNXQI+HRyM6R1yjSCZQisjCIkVt1xOBLYRb0/Aq6GNxeGqYJ936lUjVNMtcyRZCnBb4A
qfZzRrSZYG5QR6PRl9VxXg3f9CEK9Mnl3oOgAFZRtiw4Tf8bmYdRVoFHkZGDRmkJ62cair0ETfyk
bKr1Xxjjnk31qZFHBmOE9nF+u42TDTadh+JFNE4KjIZuWG9bHn4JQcS1Lf25QXeXn59ynRwLHSTl
xdL8Jq2PB0NpNF94q3H/zLtFMEtOcr7tZtW5Frh5jMSkbRwruXU5JCN6M/Z8lXZFc8coArbk1vXZ
xK6RnkZN/XXqoP5m3GNRNd7bImdqJg+7vR4STY1JqOxj3beXX8RgP508ncgS2yjmFyBfgfXFYY1d
td0+AnEA72+ixtBqQTLSbBriHMBvht05A9pTYuHlnsAcqUo+Id4YJl0hTStJabb0CDfpKIpjo4Jp
ZCT8owi0kQDqBNd2zrJgNl2/wx29WcPlTweo5i71OwT664JycDNf+Q5Cb694DSmvGZ8O1Kg0jrst
jYxtWQI0BAkpaAav9FZDyCBVwG2aMu42xfXpCAGRBD/sj5rnn61Lm9LauBammm/Ix9UHQ0UefjIm
cHPUCrYB5Xo9bMQNo+xPrx4m6IWlE+ppgB0nKgTj96tijxawTRp66Qvs65gl+RQvVSQ3LkjA7VhJ
eBLuGWcOYQBh7sM4Bb3z9HXegPsKgI7Xn6+d7NHWglkdqxPECSsI2iaU37iAybrlf2/fnzC8jKVx
j7CWNVRhb1s0Rpm8XcMlYQ+t4kP8nytN8KgsvtGzXix7HUQKT2OQX/PGzDLtkruJmSYeeUiUU+mG
itRvCw4ZlmmhLDQvao2oPNC3UX4ZLBHb0kcr4kiMWJlIsoJ0ParnQuTjiUZkw9oh6ZqcNtAs/H9p
eerbgKPn+79/3VwsWSGxFRDBMyX6NQtprYFQfsrAbEFkAfL6d3TYZviDbiF1SqjIN7NtxI5B9ly4
nVNDHN7guUck4Puq9rngtJc089P9MD7t4t67AO9x5eTqx7wLkwGgB6iUEHOFZcZc4lgbof94z6+r
hUsVVzdXxkWaFCwZHba2TB6kc0jZPtYZjJNDe8zUMKFVOB/wX0PcsJLfO7inXsHf7xZdtzvVMxPP
byte2EkGZ7+RKjoZZcqs1LFbNKyEGAFuSzLmrZkmDvI2Pb5Sk8sBjC8DWWRMZopBJbnk44MiD+9S
WH+65+i/8EV8rTkG9adnY7SUxcOam4hLtPNPBvVoUUnXCsi5LAEmYdOM6Ta/pKLldoc+u4bS831k
38Qg94HcEKZMrPGG2Zhi70aNg42O0+wtAz0UUn/K+/I5sZNr5SGW6Fl0JKIqtZ2Xwla/2sdZnG9A
bivNVpdpOT7JEgauLf0XFLxP97Kc3HTQ+coO/75cvsvTxS0lnOnCQEgdcYzTB80ceCpq33cx8V/X
I7WAWED2Rl9gGDX7PqgyLxz7GIha3wLSPg6tyNDu/h90Qv6XDSf5Y0IOkrGwooaKpvUMXoSkescr
KibZFy7eu8fu0DC980RIZjbis0qZMadGNRbln4D1rClH1y/kxsmb2flbaDTig0dtJYjPlan3tvRD
YMxBsjjqz9Z5xDJEIXIkqaDvq1OskQ4Ru0nOh58DIjD1uUCPQHs9nGDtO+B2/ybNxTzJmWRl9Lld
pbf6O9A0wEsqTiIxMgg5QgZ5xRkOpipuegKdVXS7z9f4qdFEvSI3OchvEEPX8Nnu26fwtgWtLXE+
twxLxK9vu9E/yVOky9I0fgAiEr5YigeXiknP/AKbtF5rc20a3F87BOx8W0J4xJquCsbHSYvIT6sj
S7NDwDrtJgpwaXiWMZi92iJU9C5Nyi67FlDwkZQGCIAbMK8Z1yN3bEH4JBCl7FQz0LwRM9+aoCV3
uXTmHYU5dzaD+yHP5YylZxsrcUqhsgQpgHsdymfn2bIjSqsDbS71wAAivNh3JHidWWQRrDX9wcFn
vJEVn8dx6fGWfN5ZM1uPEhMdtwIBRg52B7O/ag87mfdqXkUj6GyUIJA0iJ1EsiVnLOgWaNDk1hXh
BS9KRUbR98I13uG07+XfSX9RmnWgEH5K4Lu5rBqjJqI/ssFBVS/CxPthXNxAT2z/sWs9dXyhK5RG
VmRInezYXO3h6Q6sMUnjvvLZN5J5yGaeQhjYaLZ/cg4DnavB8PpTqsukAdk6viV808I86FyWQ24v
XcuUrxZSYhj1+0jqdC4xoquO6dVX04K/1xumGRUpBLSPkrBMqR3gnAgwTolGKAwGk1hEbjhJjFpo
G/vMDoQTb3tuK0E0EaZTk8lI4vLKp9XM2dsac+IXZeNPccbw18bkjfsiJMxmCzUa6zxuGXpvC6Zp
T1qEizp5hwc5DerlfLa2/E8HG4wkkRaKpfKvxfkvvjmcttCWdRlopOwsQZNwi/HiHrOGDz54KHws
fItIodv9C0oyGLxGuIjiRznb4dD2lzQiU/WaoTTBAVBnRmcWfJ8Nl6X2ha6e1+rljHpANdimYJbt
RbFiUJZU3pgAMIv61mGAPG69l6RAfeT8ZYM5zmoZEL87o+vXKW3AcuBzP8WRD+O8cX2VUzxOWAxx
pygklCCtS+QohT6ruzYIfyoDQ0DZ2S/9bSPB/ugmD7z+rtHs9I0EYMsJAtpvemHLMSkhVK3xggQL
k0Wut502ZZ85X0qiY5j59zTJ7Y3E8e7xKX8tZwPvvx9xg9vwADV0STTdv6q1jEpIck1CO81ufxyn
Nqf93A/2pR8dbUWy4B3431ncrH4Y8N6NShziSxQiDuVhQ1sGeoIYdHEb1b3SYWsxtAmNhzHwrRy3
/ds8kL4CYSpIoZBtzR4mo3s+n1UDpHB6sWJXLLJ3D+x49c14w4Mkw71C9QLzFBwQZIwGdMwqjCIl
8PqapIBC5FGQS6oabldxMiFCbnbkpO9Xrjj+Xyj408W3KD6g0jkXD8qmoqN5vnceDU4uQghbbCG4
AFqp8XoonEzIMdzhTrWvl/wa3fXMbKzvClXoIBLb0UUdvvlDBW2fp3g9ZkjbhxVs/UfMmfx742Q8
no2dUk/VdLgTKPyz9v8vlADtkGzIZR3ZQulzbd/H9B1LzJH+VJVLMGO8O1yzaG9M2QtbGoxtMk1p
46g6DXmS2eJ6zEmmlYXsDYqjPpEp8LLfM6ZLfs9fInDTentRJKAeQ6EYc5mAt0AAsYoC4XQCy9xb
7gb35JmzpD3GEMsG6lrgFlllvmunQd3wsWKiLBqrf9ia2KwDSpn3esxrKGjpPgEORQ59nfoCCjbD
nd6Op435p4t1wQPSRE96gmNB4NgZUCGyiFQLy7M4+6QUzODBafOMc3whIwU7qRfivygqUUxUrv7R
kkApqrSLjflpZPGzA5WC4sGSd0VRPV0WTklIHu4MdGtRZyt6F7LOg3PT0ETsui+B+/zCV6U1VVXe
SYD6znNlyLid4XJSq3T54xPgHwKGZIx8X1ea+zQpX9F86GQmsHUDzvhOhBVkP0aqtzKwx4XB+jAa
r5qPiQsmt+HKmseO9sIvJV1diyUXoj0JzQl6LQhNdrd2sqsJc/HC+EF1EuX9CfQQbRQk7Zi8o+WK
tDw/XNTrLSNSZuHkX7DtQlgP6iGKBqQLjHdKAIiYVj0DaeGo5vzMHybbT4g5Yrp81cWz89qkjjim
rkHJlPGZBSussvF8lZGD9rjoVnHC6h3IxtNDMwQAGad3uqZGGLFJkdkDq0sSLM9iL0RvUbN6yryR
yzJoytsi7htz2w2yh3WyDWC8sylzorh/h+VQgJEmBd6mArjiLmMP/0GI3GLBzTNR4BfH3jJKSfUl
ZmL+YyniA0bMNQE/ouDaqQQ3gKMIMmIxSzjE4CBOSah0Z8sXjS21N93pqSXBTvoUsv1JSSy2Jczr
G1mUPCNeAjOVpSCTKAib7K1y7oIC2rRS4ptk3zKO+3v9yVmklqzrkHVeusg0Th2jaelLdpjqiZdT
xGvlSKZ1DiFAByb+lAAZXEKFxBVhEmY4NfoKAENB5I/9H+nHLk0g9REL+u5AySA/vAg0ec/5m6ez
fVsaXMNF0nVT7E6fcOu/hVw9Th6699dd8XSr9m44uWn9iLo4laAAvZI/mlBX3yGpZ8xlbgDKZiXI
0aL0ktcvq3ojoPGeReRfJXgwRSeK1k+NvWLlKjMOR8M48p7t5WxbwNCsyYUhS+bjcZ2ZSytVa5zD
X7y+cZQbsXVg2PaZonbnl1iFrmBMFTxR0XzgVPhb9suBdlJLUOH77Wjqqt4C/f7f9YV2IOFWcT+O
Q/BWMXwUsXtqNQt75mkzbUyyz0CSbAV3sJ5u8YR1McG6+/iQBvrgyATmNbsHciTy2B8leHp0JMH2
GM+D7JzTnPKCwiRDb4ZAYWXeD+ATKZJrfkxsDvm/zY4zID2cBiyx9K3+PPaE+0I5X/lD69FHsm7/
eo1L+EuzHjScBIKvPeRpSexHxkzaCAcfcEqNQCV5LgbZiLC3vjgxyCoq1w3IP58bOrgcLt0A/iPJ
JVtPHucWL8cDHAeeMjFz8RQJwI56KbwTHJCWPOjBXOn385akJSxj0m3uUYiFWGYR1dWw5vPrH6IJ
mSKq/HQWiwYKzHkruLSxzbvgQ3Dph1/UGE/VX1ux6rYClKMT2dIvK61hTXHMXM2s+Fy6FMedjYXU
lYQfbKdzqqgdkCQI8dr86UHRBqQGH5+TfJ3QTEj6dwIEV6pGof7rWng2uhpdDRWDoSAmvzGwmD4X
Xg9HtfHPvdL8AtI5OFQinkSQ7HiCVZe05wDuxiqc0HEUTob0czY2EMp8JYvqpOY996hHsqyKsA8Z
NjWwzZ12F7Z4xYHhkzr7/yFTOySY61/07AKFcgoHFifsen4W7D+/wyqsEsDb1qcadMxblSGXR3wi
Vkb5yLHMNU4uRvcph/jPM6QotyV3XVEU6UosmxBcNKBxWX3Gu2AUR57MPJfgU+7YD/UuC99xnQDi
G06MdZi8MEpQut3fMZKp0859wdjSf9jRMiuIH/pqy1s0SW4BjE5kuaHdi+fPqPo6MwZLiUHvYVhw
yOpEypsR2b2XyTxg0tBZK8gYThfcvTz5+9P5A4Ru1WHbbd2wCARh1n71g13JcW41WY6I2Lt4DpnA
jaixvnsAc7zIUIX4r1NcQ5xWl8qBylLVsey2ApWu/XkHV97RAPThd8qiFk30tAl4dOsECFDAkUol
YqJQqt+gqH1YvnyKzOH7xuwZ2cf3Ayzo/BEUvA4xHy5mSMOaeMRwbgLYhZXhrt93kQDo/xnGlzVt
9HQCs71B3W1aRDKtL0LixWFGkkctwMdfQY0Y7ItoUSUCcMfi5l7lDdjzPxnQuVioo4Jg9dVgBcHG
NmmZt1jVt48ZyIAwM2akNPjNuNNYPFzzlfi6CXnjBYOoPEJGQ3+5n7Bhro0BRRXbgwMcu2vxszK4
4qSvX6erenw/ohZ+Ej8aogznKm2CQxVWXSXOjsmw0K802/u1ZePL6sRMLNJveUUZhTmmTfLzveDa
kAOA29X5IbwgvrRRa6gpG7iO3FU1tlk4lw2/HCwZMR5JiRiruBdlUAoVRfYS8sz+7ht62GlFRbhu
wdhAtyRAp//cyinPNQcOKrO0RAfzWMTmzRLlpOycewYbN2XjY71ocOjvqG3zH414PKGrjPCWP+7a
+WY2KK/OOs1AJsCzsCYsvQmaRFdH1a1sLZrOU2Ugc32Tuyi600mhuqrdG8wgwc8PbJcZ3JfwfyJs
0IASMIKc5iC1gaef/K9x/NZxa3LKaP3OkmUUlVFiUznDi+n6EXVQeZhLh3sj0wpMAXHGi6dH3Cw3
ruaFwij9W8nCb/5MScUOak9ay+mvM41ozgTCpFertOqkw+Q7KTg3/Hd5ZSzErbKdJnHqd3YaCnFS
TS4PnMYTi46z1BZUf4YK3KZYZUTdL9t2VOuatCOXUlS27ifSb42SPhy0CeZKUCeMn/yd8Rb5Mnah
DJzHSJSojfcdOAY1OHQEFMn6uiHfbGpv7kYWGfMq9z8tKlZM9NSlcxHvnuuFGRb7TcfqYQwVAZNw
sGVRIkFiLPNy1+68SGivc4WqU8UCHBjO0hj8FwqegxeZydMj/mP3nVG36aKKVppqNBexzTZ+Ns2I
AHTcy3d4MZE4/bF0mGSHzi64q3BG/oQT3HBAcQv+LEHvIWNJqL+/qTbMtJm+rx5L/ERwP2ugDf7H
9QIqknsSWXRT2cs1T17XZrXUlYStf+Ywrxqx5tmsc4hi7jEklwhN8NgCOnjB0at48rsLFRRA6lH5
RNtEPz78yoMG4GTLVfp+GUWNgZK0ac4lse2CU10IEXMx54HHXff+45+QEHslhm5p0rCh6lFNhChi
HaKtCgPduF36mE0yL4/jKSEVpDaZNWEWjkrCA3pwMXKfRIEPzhKZ3/CuG3wQOE+GaeoU4CP/LnuS
j2JRgHFmth6ElxsecaUXxeL6pMIWmTef82IeN8Bt42oSfmnMbNhUSpd0VIQlRIxR8PMzoFp6XZ3j
k/VAgEUREh9wWesmXFN4LNn5tc4RTzD+2wb9u3pgXHITYqaR0X5CZv/JTEzifQf1f+lukKzKdbiY
jI6KXhqr7Ie1CCKj4U2E2b4fvUMQuxV3iDyryTOjbfUnzuF03L29/fw2sx5NV7PSE88dUo2M/hZY
lEjlXOevlpsPYX+9lIXJcMac8Ts2+co0Ag9Sf28E1L2Y//Cp3vMuoDneyFkuMT61X6JQQ8tce4NO
TNPloqoocz5ZCj+xOR+jFkq8AYU3bwwqpElx0YenC3c1N8byKPZaEQEvCLFMk+gatrYrREtxiL6f
MJoypQ1KPm5WmVfaqQn7dIYTzW4abqxNWfmXEogO5jw0x5ieGj2q+AVWVb5eiZMaOL9CeobHPWkI
dipmwzY0hDq0jfptF+PMHC5Xv3ngDpqH5e4079WyG+lhq8J50VQcFtWzQVF02seP3mN788iwLX8q
4MDeqhbb8JAsajZjdiM3z0hwRYg50iX0RtqO6UbB6wGG9iC2OuluOZM1oc4VCJ71C+qDWXwcaq26
8Yuz07g4EmwwrAtl2oLJ4ASV9UeHozqVmcokWwAwgXWHUrqnz8JJkHWjIux0RShc/F47IAE+bCCX
yHRR4usZvs6kPI0JkVBuMGuHrvtVW5xXnI8r07h9vwxxJ/YYVCh0Y0E/Le2Gv36sYHAFj1leV6Cq
fMwShObF0vb/sc4RGAnNDLxbFgV1aEP6mdQoPjqtHH5cMtDPA7C02YIE8ifPHlyf4OSCSa8mm2pO
ZuI3NKJ+/QpVHJ2Jb7oSX18H2hjqzmM95f9Z2e/QdkkqCx/g4a2c7fKybqz4DeTgrUoiWo6WYzO8
QKf12PM7fjQ5J8GVbGEl4r4oaiM7+XUIPooblXSyPu5CITw46h3fPCso7/0cNbKIVrPEOoJ8lPk0
Xp74CIebhG2TzcMqHwyF7U2APuWnm/D0LuQg/Fw1lptUCEMDDGEL+FXA9P5CAflz/I/EdsqpiVpi
iNbdqPjCMUaocK5ugFfW9bBmSWv4BQuV2o/OsfNrkoGu24sCxb1KTMT9Rze5Guj1NsGC1NbAFj6d
rZduAvtnba57aKzpijCXRzjuzIehpaJJ887+gTgJyAIB/tVdvaabFMXXod758ro7K7bUUMEMp5pe
CBCfSfQI4BW8EAD0jyXXGsOq7zF9xSSq8Gf1K/wQncj6X9F1Pey65kOS0hHQiJpNYRRspWHLRbcF
cNXXAMu9oBvJ3Pz/p9+/TRq3Hp7Y7o5jmae6sxM+9f3BaNg2g1R+D6xhWDS3VvB+EWtflnLPRblE
lX9hPmLmlCWW/Z/2PU1zrkDmUqdi5AHj/0LIeOvlL1DLadNbic4ApIezkW7aFJrcBlJxfHNYP8YF
YyW94q8I3apRwCYHKFeZ/VO//zPu9GRbO3Dn0IhsRD49dQiAjsoYKiIcqG2r6W6ShIWJ2EU6GrtK
N4Wt35V+WigHHexG+c2/DN3PtBV0m2ddVeDkhhGddISMb8QbHf2guU31UfYqjIdHHIlhQN9II3XQ
n7qHeD1IuHF89HYOF6qwhqo4KlU81xbYpfmTBV9DKtvdDysjLKN2jWHIcnjcKVKHBFE6170cnb/C
kMASC4HAK7QS4dHeg2UsMcKDD4x+MrE3e4Hsd6Bow9cJ88TcYthfR9KSdr9FqUku+5AENKF7RdI1
n/tC4RFQC99by9TRaydVuV1dPNrlinJwVZb+vkRdyR/rFszSVg4LUP8VWkNkhbOBAmi0GFbec7E1
jO/E71kwWfJ9XWnckbfdS1tbCxzpoTH1Q2luvlLaVD1SLxtL/Y8K4FCvQU/O6OVrZaTFfizioDqC
0W7u+PkuTzgnb1iMMJBA4GgZtGkFKUSvhRGV/OQdJwSZskSxfCmSm+eq6dKRS+2GmzHU8yRtDH/f
YwR2zy3oy71WqyztBu5ygbA/QSnOxZV8jJQZ7Mqp6xVg8QJUmiSB1tEU92L1CklwitQhELh/hnLE
tk0HX7Z3IwSoqelrTu2TpaYe8fmK2viBvktO64x5iWMzKH0S/JmkSHT8TCT5BIRI5RRI3aVlppay
n1AU94Vhy1p4vSw4jo4604WIGa6uEypDy+99iJ8WwnSQROY7ezki0IjV7R1p5je26IWmoKWwJkF/
oig/IROmoRQm6ZOspzHs5pGSUPZ4j+VsdF80lmNqfticFTsa8qU33sUGjMsUB99isrmNhbvEGV8u
cyvkHrZwny6O7bmGVYP0rWL+LPwL2inVUdVYB7pYb31/jjucWT0wOarixfACVnIdFR3JZ7qPaTZH
tbU/gTc9HG+dO163mrkJiDw5Qu8gH77cs6cnzzFlmx6FzjfT/PbbuHZcqveJ0aPZz/yuEsO7Zm7H
ch6GTPWxUtngXaBgDDo01Qro+CYUjEoa8mbDXgFN/9vV3i7/ABukn0ZdEePOADXroKvBtCVDCy0E
3/sOU9IKJvbSAuQpISJoiAqEgm0tFCH0qyVU/2iAzeqQX8PeVwQDKeYURL96VaGbV71Xhe49tyIS
I232NtLFINI7cFkp3sHwU8rATIRN5qu1pfvTrDh3ggMllILpazjXHWlhb5Ip4OgzIcqouvWfW6p0
jceEDjH6G9vBq6tejJXEEuhgRZTNgY70sNBkr/UcpwGp37uw2xl6NjiN/teu237fc81l1pLbEk1v
FQ2+dZd263vhuNzf4+oTxHhu1N7vlqNAxxT7xxgbAXCOi8fwwvGx3ia/k1eclZSYFnDVQBEP6gTy
192fu2eTW+9PdZnwazTvL9RqW7uKq9eA+sMIxqwRIxFpePHya+0XxjwS/NHZIGK/k589Wm4/FRTY
L79LhsqlTUzx8LyNDlmReY4soaadLrfxYquG27HYaiJL/oSiiwsVo8PwPR7/m3twOkaUNLXbVqZf
NnaghnsJzpfpziVknHljwlWx+3D8+bCJ7CoFIbO1EZrAfOsJw61bbuHG4caoXzMy/omYWIlDDG5N
o/8Rb6mGYTieARQ8UrR0j8eGem+heklLsWYu8H3K5NGY1BL5ULe+fQoDI92DpswQMtUpv0JBRT1L
mqgOypabYmkDojYmNFlSgo26IE9LM4dvfS4W49y9zNAeuLJW2IiG92TOAssfVkfLaS2UYAZcpjbh
3jVjj2EPuh9DJ31pfbRdV0qsTn3TmKn7e1mTn8wxzdivPTDQr3IVMq9Wqnq0AXCF4O+sRwG/2deg
ZFRAUptRCZ7LnrPbL+LlDK1F5Y285K4vt/doXEXQl5BwUhhEVwnI/u9PYDpBFIN0El6UgsnOi1Uc
uwiWAKTFtnRUxg+Pyev3ogqC50jHwlTD+l7UpS9EA46EN7SRhBzpTRcy7+Cjrp1/C/DqMyjp2qTA
9iADvAdmssdVxNzRUPTGDHm2AW+6k/4i3qHV6Ic+rzXcAajvANjZPMzQtBzE9dNMNWNHqU78FZGM
yj0FeTkHQ26Kd1jj40LnHTUuu4J8wSS3d5NJJMMZv3MW9k/xz9gB3QrpS4z2OwJ/g53RtQCaO8yI
RNMFxZA4wS506FFrT1ocizTU+EcxMiYU/+3VWXF72ITlC/Ngda3qUxDXCgdienKGLWXb5Vwp/dXH
7s/Y/AKOQyS93eLgpWPX1Pc32CCpFK10lNRBwdisB75gbqooDUjXWerxHCTGzU6XWMq25AGKPJSd
HXr0GONg0HzL6L9q9Lj6qIuk8+PMoG09sP/fEa2RP1JF0Gc+SMWj4Iff3aZ+06yM1HVdxETyv2N9
hYt21scPpsroFC0H8H9o68MY5DJNO94aKLYkuTsHrmW6lCVPQX7BSA3jY8hqnoHlU43uXNU5aXpu
3cEyXjYuwJ0kt/GQwLwxuQFulOJ0s9d9By0MjX4ObRVyYOAVGEpQaXSLMIgq0b8rbrAQNvxS5Dso
oQGUJOOU4+d/0rTG9cefhXRYC9IaC/UHQ1W70RCUovKxFAXLyE4C+YwG/gSQfnJ+1eV5jB07YUgr
Kcz8CggnWj0YmIMpZ1B1rwsDrG2hEi7BKaQHzQt23B3eMnzPJuLn86sWI2mts726CRz2tMeKrH+z
ZLz+cxYPn2j9vDW2W3aSH7yHUUJnEOC8+pEPQZ11jMbPtRTwOAH8G8MCfeWp5XAczFeuvYu71rl2
4xjNE3NmkEVt8OTPBdqRdEtVDtw+SbcpWamNM/MSmCJUwIfCnXztAkKPJXM3aKJezexnVgNjN1UL
8NN8ZO87m6NhH7rc3Ik4rdSAwMKnadBT7DefNjqY+ftOqN1g6iGyVp4WHe+HdKAxPngNaNWWbmE+
0dvGGAhFy9bMJchIC+jjBXhgOxCANLm96PWuBjMEPKwnKB8vPGUIqnH80HftGtNNMoAeEdsoMy4q
s0B9phOYoEcJMjVQ0Y2JMBNUUetwk3iqymQL+kt1ki1AWsDUeSvGEaEMOqbq4jcuc4k58xM1WUwe
6dhYUExYmax5zxTnL0VJ4wEo+eopwZYgfvseIFFHj+gdT/VXn/B1CmrZ6b0ziVZ4tWyWYPlaUWQa
HbQN3+QhZ/t87mC+jdFNYXdKjyQp0p1SxaAMvMQ/m50vM/ZK9vrPb7irfrDssdPOiWwiQNeCajWG
TMb2bNPPFe41G3rL3jruiW8QJEsTrtMQ3d0gtd3R4doOhHeb9t4Jdjk6WFAljp6P2C2hDLhCMhEJ
fKAgLN6C+YOsMxnZBhFsr4XqITls96GEnpfVx6OQdY46keYQhR7GXPPBjlXj2YchWBkACv88dvdP
NtSUhWufE8YYNv+8cdHsNeAvIpaxXekKOliqZG1V9vEU6TxxAkyEwTXmzrjipylVK72QY7Oq+Usw
r53BwxxOH5dqLdEl+hy/tFjrL1VoTOGY6tKnplTnnojvtRIFz6WI4rHizWe2sHsFdHjELfPgdaV8
CwOYU4Pnh5btZLJvy6bjnjIAfNh+/IFPcEZqDHWHEGUUkOMg2b/KWDgr6gzHMb3xXNv4h3kkT+Pv
lH+MHd9zHVjZSjoYy2NWRYfoPslZzFM/FS2soQyYtDMDTmczy1KjMGudMl3rAc6BdJEArEI4LP7k
s6dTHBA93MmusHWIIXZNpSFN3RCYQzvjCdkXc9VqaoAib+FPMGt4uxLInW+FF/kSP+jRDx7FDNoj
b5mE0Hfbvpsm8Xh/kkLtYzvSsqC4Gq8J5Z+IcxyXQeDcmdBM6A+YYh7HAeMto7Gp3qDz9qDDS2wU
KRlAxoFnUksk850YYuOf2m7FAfLKCbSqoMP6dt4BQyiSy/FBwHr7IjOdqyZ4OsvAZ7JBqbGpLiIJ
1hx+kaF6cNHG/bxuPDQCKHoD1VtGvAVfLSLoPh/O5tIfNet8Os+DlLIZDGHnlOujNjkEiwtymJGP
biQoManVlSeFO5XeqHl3ZjHNuVGOnFBSISITCYh2mD6wVA3llWelAdpdP8HDI2df2oYWnyZn1kBb
wZWioFslgjMSMaNRLmHxdslg9btskwamRNkb0cMk4yL+UoAFoMszIjyZZV0E0FMaZbJqfqTJ0fUL
jdi8U2YqHL4CElSH+/xfE3heeKBuDYHom7WAlCvbvbAP1U9oz7M/6vq/mOMiOrOGyIjBLLMhL008
2XaEjaZTiiCqVzfbrlRWUWlPY/Wp4BNVIzhrIghDdeVEABMHilgV26SrlCqDNkRQ7wMI3sWeUj/p
ALZOb67hmxCITag4OIN0BCsi6+s4HzzwP5EI3rpq04dov5QPKkgo+gTLY0AtjH5EFVnyuPyQSGqj
ClYWDnvPUDC6xiqhLTM5z6qAGHoj+0sbvSPvStO1/JZusr1Mo7I49AUssIYBvq1RjoCwfgevYMFK
YCpxG7jKsNWof/XgbDBvGuQthIaU8uT6c02mGdKJMiBuUjTQ1zXA2rvQloayjjBXhirXBg5xGpuo
2i4Q2Ae6jWT4w25f1jCcyq4/dumsZ3V979bk8XkjGB3gjDDFdS/vwxc2pIjEDlAShzqHjkkQTq+h
l0Rs9mOCCY59g10Y1kZUiu2FkoI7vwY79SMFZgVjXs3WWpdce0bG/5zukbNS4BNbrsFHI9kkKhn4
jjTt0e3vTw1bvPo4o3GLdtj9Gtvn+tLfgCGrTLZU4Z3IvDgVQ5HJEXxGKzEpJFVAswtn/I5z2LoJ
dqngJ7oZ9IxCv7PDyZD26o4QGPBbSzBoD8M3Q/I8t8iIC6C00zQpW5AHQz6HRf4vJUjFJkcgjCji
gvPPMVQ9w5/BgtpW2si1ZNHyinAC6u4XraRnOaGwg8bOif6pnsdNCJCG3K+IEDqQo2ytulYoBhkB
KkJv6DCWvVfHmuZ5rKJSTM2dc95G89jinwyW+PNjbhTVa13EMeDJSb226Modw9nSARD1LMFKpOgn
HQfoE4EDlPfenoxXiwZGnKz3SH2q//+/nbN3TgF9TpTJIHdmByDqbRZZ0lcSN4691wM4wil5TD0o
FbjLWIVNC7lwB7l+Ui13UCMieYh1XPKZjwI00WSPMhGcRZQmi8MluOmYK2uVlZ5AhNIty77IzjH6
oDt7tv69klLEOtCb9R+BJeAoVzk14pgriRRrBkLsYYH0/ojv3jEdPDCZY6zVyM4JpiMfPw8cPxQH
JFP/K34gP1BljT1/TykG02aUVds5riC1V20pk71gGQCbEVcz3E4GHRoEmUwrOQ0eNBh7J0jr30/F
1Oom9vUPAgyoBM5Ocon9iKZ4x7+NJY4g1jFJJ42DM8PNV/EL5sXYgRwu2084hRl/jXn07hIEDsmj
AbxoH53fsD6/1fo7WaP2CV2GDDuIdjleqs0P9Z+g0K6CEi8tz/yj8NqSDTgc7ZE0ZSXJlOBpEynz
7uCEV/qnHqhPuws9G2ceGA2CH7XTneTe29p5PmtYETY0oMNJPq2QDllWMEOBuT/peA+1R2PrsIYd
rHolx17Fp20yF4eWTLRe+2Ujjf8I6jvc0b/7I3W/2m1xfHnwOM6Bw3WVc1b0fML2Z3d261QsyVn+
ktV+Ij4gpWG2DEtUVUCmlwBA5crVAX3uInj661I0Z876+814KI+7iRuS0eqxSUk0RimKtw5AemCB
4BG3BTnVxn7WkOqN+szcs9pEswk/f1SuB5FCL8mbMlkXQYWA7RDWysHQZibrWJO4sFqqFRuVsD4s
a9enaoRWd6dXyLVc5GHZMEOztNbD2z2rbfq5oUE1uhgWZdTAXYzv4T+kcK9f6Li9nDcaCReg4pq5
z8As/myJBEADmICrDREv6lVLDiMcUMRq44iUbHYiboBgr3wCUp8/2lkseACOnqSl9dli91xeGRrb
EkXRNLHywS1BiW95O5BROrscCIH2m6RfOGrlsvSSWZSJh2Ga/j7BqYnH8VbPNGEvE1L11iL/uhs+
7qEMx/c0m7tpGmBWlZrFBfTNV5MNlBVa4QoAv6B27jMGDG8R+6iKIvpJomL7suGb/orNneq5XsB1
CFejKF0uIo5VseBWbFlof+7pqyFttVxwq85Te7Q1qWnSM31Mltnzm15OtgE5zt3fwnPYfBfEd6ne
+SRYS7shNfC/WB4JA4f1+9T+miALfwaujulwi/lraTN1f7kLNsDwxgGtqXVMmvnwYH10NdSsywjR
3bsxSYnXxwtDRK+8WQCnCi2DGG6ajtXvIV4Z5j76RFP5Ofi4j66/wMhfDjdCKkBvb1RJ3xi6kQ1G
xstbPCfo1WdEY+fHFI5cyl3MSJtsHzWePIGNb64SH6MFXTD+Fh837AdHdnLG+m3RFJKlbVGdR9Bf
i4gxF7Lk3jvW129olExiNz+qAujllnii3z2afIjolWou3DJQ5Uy2QvSVpq6w+XqLPsrNJiN9I4+t
xNinBzhWuWgTilfYd3/vzbRoNzitFVWQBTCH8A9IZ+64Tujj7udQw3cDE5cKN6TRPeDTzIqQR/X7
48otJ+tMelccaL0iQOfcCAnrP2fJDsDYtO/pGL7BshrQf7q/pF1CbJ4AyXQ5RydXml4SGtPHNA7s
wlfYfOCrdseDg+e1kIpbXezObztJ+yNmKh6ht/OUvkWuto2uOe4KKkddxWEValv2mWBg2DzCaBQl
nkFh0c4pyeJD1Td0qN+10Wx1YjODL+6G9VVO9wZgd1L6YbFXUqwqiI2dPJOmXGienuZ1KiPTe5l+
7ChseRTRlWvGE1qDMAnnKtaQ6Yv23y96I4B9Tit/nxixGFUBXdY4ydABHpcJ6ks9dQZyAlyvNK+v
n2NahQ2zuzVjjF/95Ex6X8iimcw/KmcA8CjKujUreHiKgoGqUK0//QNDLoWPNA7nhsbpirxZgYiH
Kpo33lE+QDYDuzaAxaQzT8swKfFOI4eF62VZkyCP2CzGS9dyBvD5xAV0GmZj6WLuEqegfBe1cvgQ
QreXn2N8kb2rPvc0NAklXw8IEpKMephF9uyHyV+2bbdv9U6eYvF/jpv+/MkcL3HgKERoPOvgquj/
YevTMXttr5VAlhsBXvkfvrs8hFJB0wOCBZQPNhwx5Eh5HhHyRTTwV0a7+lw7FplZC4AnXfJ1bMjL
09BTd9JBvI0tYa+ueiL2Wju3mbx6DcVBz+nO28oCNyr6kqiBpxUJ5cgnATD0kZHRocF6JqXvMh/r
S29Rpatmk+Y7Mf4pe4qI+jfWsrsfShf/JOiVcK7RPSAYF+dg4Ju/w3b1ymLpCKcGAp/hs4gMNg0q
jDF6ICW2HWUlTKJEBmeyKPvwPNgVRb+ywXHHz5cBF3z0Qio1+eEwXmBxCBB9yvR93pSPftqXB4v5
WcJ1XOySSfxcFr0LlRDpx7ZWi5+yYDvlEY5EJRR4dY19k5CncRSOZzUyf82dHDYytHYaxPyZLndG
cVdp3MtJJ3QSEPQvZl5RyaBOzPZ3CAQmxUcHueoOKlbof2xqfJPi38U4VjEU4aC0UzSV+tRAyBC9
MJInro6kzbHx3VrEyDnfuIv0Bahsac6mGepcfalXr+LZMHJwhiTWdCgxOSt5nNYaaKvDj0GCNNEJ
lISGysMNpcaiCD/Cl0+jpPCTNOT5vbkIPxP/H83uoUdre0m5zitkkp8lBDc23UMrDIkGHzH2JTXa
5syFPKcUdt0E/9+etqD8Utohk2X4DtIKX5fy6m5mdMLaPyjTp6oANf3bo3/kSfjMcgjYRBSMeMQG
EMUkmvLxFsM1UuNIxNafeqY3nEOU/Vau0hVqlsA8vfrF0s6ZQ0F/C64rvt76I6x7PtE70FsGWnNu
pWJ/krGVlJjgpsbMMGlb8dd5Y5LTUUds18sBSdbNnUw/S0V3BYnvTU4gnZBQ4+e28hWWFrDqj70o
KlQNpLUH+tqc8kMd+IDJTwHjkSBhB7aVsM60acsAyck4ME24ukViCR5EGDjDuoohZCsOqA7Dfh5+
XHcbxvs7/4l7DlWBxeFvsljUADM9onKiaaM57IbSHHG8IzCUKTvKwCy8MIFt6V30T1R18196Maps
UDElM7V7HsKBramgqliGnifABC6QuNY49QrlH/9se1h7GrIsjgOkkMWcFrtge6ElUSWOFYNAlUMZ
WkQGxqNlpK+cGoEhk7TPKluRFK5RNh2zEoqUbxwqsYHsmopeZWTf0J/jZQotwa8HLtPDpArOZLx+
33Uo6wswfWdFig2YRWY8Ff2LIvjDVkQy6rsIwsnYzVRVIMmzoKiAwNhgIpGEN+7W3DpR+YY0hSD9
5uZbSrUCJxOcUvRRJSTxpkJYjZd6sNaD+5NfGHr7P2PsvkUk/anXR3puZVrwaCL+dduTz6NvDQ1K
8wkYlx0RJGFN4THIXOgkXFxGpNnGuTrEGCOn30H3YoVrHc7R2Sq5chITD4zjTwfCys8Hk1N10Ngy
sWxebMSM8SotaZzmyiIhLj1uFyxlRMXZHX3W9O9tB78u7wkE4ukZDJizsS8eZ0seUCc20KdZGCPB
viuCc0So8Ekv0VWAfp4qy6pVUEf806zFQ8UymKeBqLgL9Ort93ijr6s1Kc+t7NInI6Fzk99R8xJg
7e58F7/749WtwTskrLUmauEPLtxYWldziESSQ/BmqqvSizGqqiAOm4PgZR0mZe9xIvtwUBKj4H1b
Z8y/cKGuwBfuKujb4/pGRAsFSCz7L5vC38vtVApnWsNIFiORl36pSodid7bYxpR8ijsCYyfSqpj5
ejTtn8s0xd10MOQU/HbiN21A1B0cv6lrRuUWPIrUEn8p6S/gHpx9vGdxQpCxxk2VZxRENHrxzuDD
xuxskdVh0iikTcvTcXlknmKyv5o5iiT8mkNWMAs1ocqfMiciQFrqYnxOhORwVQ5lV3bhPihhtcW0
n3w9hfV+SUQRFHoU68Dks+FGGVZxpjqJ8Q5oPTgMWiRF2zx3VtEXDvPzap5EPdX7dtkbUd5OsA7M
8siFZ9rDUNQuWsdKqSnFLupXSo2Gvzazo25jWMQzNGOBtzLPB1DkQt4SBwYPIlbaNiJ8WbHskAPx
PSvbJUk=
`pragma protect end_protected
