/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
qcbaMgJvo60Pq5oCDZjXn+/e0dQgF1WAh32xcrhEgLZKJwMnlajQmiCtMaOHEDzfn2csJPlCZoZN
OkVWHeMdR2vTURKFO6Y6KnkwGHJHlqDpOXI0XkQM8erB53Q7lzNqL9oGZcah66tGkEIAHpDaQemS
Fr11EMuWwImHBUzBTc7LxdcA5GgY3SgNcVfdUyXSoaZ/lGiyOyesJdiSKEmJ+/2TcLJ5mJbDl8f9
xHA2xY1MY21PtbagMRDYWgM462GICZLFQ43QfF7RrtvSoFj1g0MOGg5S2d54mMrzpry4G54KBN7T
9ihV0UwMjUgYLLpQIcYu9465/MXeXPVYBuGPfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="sm0IVXHFawobgJlJbl86XgtoBn10LEFi5PF+jINV8yY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1264)
`pragma protect data_block
75IwcHdBz4P6xhMfY0Yd9S5e6j0T5wY6OlD7PdhgWTIXWrcGaSQZOGXaetpukg7vdSHW7W7cdBYR
5hKcaYhNJSxSfMP9eJScLaCagpbotPHsQz50aLATre4pAtHIp1HqjEsDvIUAM1cYeBpMlKpCAidU
ASAXao1QvzwQ8WsWsStWS46/VIRo3Vlq23vLqhWOyTKqRHy6Ie6TAKmxLWRxhjHnpRyyP4+sQQk/
IwyDRnNKJsSkz2A3ESk2y3rahFS2S/k1gHR8ZoYyb9gg3kDrGR9y22SetyGAza9QGuLouU8cG6Eu
8zr3OKBwLHqJoFOdJcLiIc7O9ahyFuCb85K+naQ7OuroON5+UzHt2clGb+3o+zt2ujNpOJRn4GgY
/Z6BmQWT16SU3BqGVdD/1MiulovbYWKuX2Vza1cNiOId2+xnJbjtsDK1aWe+ZE+i7iv4kYBFF3YY
LWwt9oJu+M/4ZqGbDFsQpVLmLMLy8yZjrh855Pe2y29rMZ5j9axp8RhdoyjYdDCjw1EIbl5zJGGE
wp+cFPqA8/BfuFthl3ouEZZpv+WC20wtCLgbDY3y49inTm8dAKgsHqLSf9GMM20pgsHJrL/SaMWu
vMGM79kI/SGDm2UQfG7q7qqi4NPEKe4NdfE1rxIr6d7rASsdGC+5R4/I6m7D1hpWGjVtLq3xMpgR
eO+853QnrLLKKABCdgpGFg1I6sdv4gTnKJcKSdLnKptZx1uKwZSETlNV2XBtZKoZHLzBMZcekWU6
l2nWsxKaUuVuk52dilzPSXJ+qlEciF+tgVwnuEpf21Xx4aA2EpVDiFK2ieXpGv/UKjJXQq3SDDSr
uU8geP33VbECQeD0wCWP+xwzfqKIHwrPiWPcZyqJBT1+aaPVNFRUNzlmQbs/zCcqGbZotfpdP7nx
2HeLbZy/74+xmWhkU1gOMINGqjHBZWLEtgQgD4cIz2fmyP3CrFayuxTM5y7iB1j4y1WMysmHasIU
bu6+0dUykj4KYYC/PwhU0oaGVLEHioSWR2tOAodwGyQoZm/grStBs7D6HlahKQ1uK02hHHHB4nf4
XCrYpFG+0OGPKsm/+UYFX658o2t6LgoyY13deoC9ey+2x6KRcCUG1XknPafuCX96ukpFE5zOTxCG
ATWvUu8TAPB+4MIKkJ7rQ9/WnWTyXqI2JqM6PtoXcOTnLehoPXWE8IF38xK5pRZiZhSqig9HvZLc
7piOZmx1BRZ78upyBWg1pwU3P4cJJzITRRk429XSOi3J2nIgJT5feoDXk4zyuvuuZBWxjnaBsUoo
CzdaKKtgr/fQMH02JTUBhiHeknyrLuqZjyD9Syv0TEw4xEg6F4DQ8pX8fU5tRVYV0Bveh4YKtrXP
m/cacdekgFdjvHsJSQK0BTlZNsVHQhvB/gue11K4V/VgWA8wOeiMZ0q2szxfs0Hped56Eh+kfHRf
QNQJ4U6Ii2rm1rw2tXfm80IAHAuLcj6m60kaWzf+upXFTF3YLokqlKJCTorMrpzsMkYUy2udfQPh
gL9vzvf0b7sI9LDqmyl5JnSaBcdphqaHnVtZyD/VAAOvEidIEgIv1esdTuup59vSSfVafcjRYIxe
2wqhERZqn9qZIQcvvQwRxT9MOouCKR5IKl4uSCsB0FiPPgFVLMg8CpRgUNWvGe1VpARwDsy9hrlR
UQRGTZclevgC+g==
`pragma protect end_protected

// 
