`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TTpFicC9+wJbhghD7UOcmGgqSC8TwSNojXM9T51vv7IVTPY0NL4jpFwgOuqzxlmVeit7066mR9z0
ySfWB51Q58TpW1oJ6Vh6yCJrrmnYeFNVx8FLRAW8/prCNfTJX4FogTh/ZNmlbGyoPZEc5eur6xKh
3F593yhnCpJKTs8t+23wdX2VG9qVASbAPCVCSzRgKWFpWsjYfaU7duorpkNryJNeZnZeiK1IwpdG
jYcP5RoLkDBYBUB51iL1LiD8btGihLmaZQZMckqVVBN/ZVXNSH6EBhP2cBkafecmqvqnN6QlCSfh
CFV1WuUhGO8oePThpzRm5zULqFC3hLuPEk28Hw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="bp3ou5+8ebIJskwOPYlTEoxoB4tP2eoER+X7Ckh/Q74="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
pVzI0I2MU3zVLki7YfJWXSNe51ELstt0y+owk/Lo7QEhp5L+R7Dj0yJ+UEcVeuKe3REvYirkhAtp
fPeHcI2LgM5nyv+6e1DZ1ILoM55JEtYHTFIvX9ETb8N+i3a/W5ChQThYSLqiGlOJxb2RwyIItivD
obVeUkj8ESKi8TWpJ5bXTnna2Azr6c8Gu72LWMMuBZn+Ash+p8tqiKxH8MMlGSBECChgnHgV7DiP
l8wk1AuuoZ+6tIFtihilUhvazrnVSV1KEpM80GrVnAs+Gpssl0dbzWJAD/8b+XpCDII0f2FPoDf6
QxPScgm/BSvuvcxRz3/knAeKWOb5NnBL+c7SvGuDevGZ74vUnZk5fZXE3FhL0dRb7JT6KkoIIsIo
3oikfh2NaAcGghfllekowUAe+bXZm9VPJlgf8bLvCJOLPfypDfq10306JMYzFUbiCiXGttlEHJbo
Jd9GUrLj8oO8EmmqDBzo6uz8a3Pb5WQPTUj83vpRnVtxzEJNMsvw1b/w++D+n0gpiXCkUNLh1+0+
9p1yw/lb5e2WF6VN3w9OfGq9dczfIhjqOjTvRrqYrskFFJ2xLOTsWTIaO5D5HrSjuemPw0ZICV2n
+RG3twoITTrt1QAE5MCrQyCz29Yiz2TZi177UUro5dwCJxI1o3alapYF3Jo3jvHwJFyNpgMzPymw
oqNMCPqtx0/cbqaEOmHoaT9tN1412m9eBYiTdzlgGu+jSVKrxI6FpEyB5gsjswyx8Nj6NbfxpAJa
bQaPFK60qJcnTrgQTYbcnieJM8aXIZXCZkJA74v6136Ln+O3H+XuziZZ1fwGx07nwswgP0W2w4+9
LaBZxYSiHASAuZvTqag6qZUzIFJnONSMnQlP8YQozQ5cBkhvWX4SVKAeYu2PBtmptGx82OFqsJ1X
lFQWQiZuSR418I2iJJC1wZiJNs/dT2krcH665BBbuhFpsdVgeYZWzQmrTkP5aZ44qp9sh6xCscts
bq/IzYYKqIexYz5vqMGbNd+SbyQ4KNWCCRMpacL+x0RaJPzElr1OyiACHfCs0ZPyPGiwkPSRPitG
eNaFwJt1cROzy56eOs6qP26FsPFz8L6+E12XiK4JAs/D7RETm/N/6GNDMeo41nq7dcnK2KD+amC8
tsf4Eq72t/n9XRHFoRZsSidsFeilSwNk0j6zGTgIJe7f48hAqO0tbxtbxqng1S+b5/En3vni80fn
lSbrSuRam85/QxQOW6H2ItwDEMb2x8W+G26MzQRDcTKJuBOrumYol90xaCLZwvhsg4E1zPqkqIsd
QHxnHFox3gsm52yl4MX6p62WXcr92Wg+q4dnzUEHbueJbi2UaeSnUJWbz/XOJFprmnBhmQw5ByGS
CBJeZRgAaJa3n/3oUkcL4KEF3crjIAk7LjwowMlgBBlAzMfzj6EKxn9JpJHPJomgBwPIMhPIg4ne
T2nRKnoL7hdmSp2enHB5HNXfqqyN+NKWGjdYKW1+9ZHpMRKycuVUykHL16OcHnwd8U+nhk1wz2nx
g/+U/AudrP/un8k2Pjmkwwwborb5LiG//keiGqPqVn5FsChobOZUekrHU53zB6zQ+OUtT1VnMZbY
LVTjMyfMh20R4FUS3SnuQRaiY8mYBPTeFZIodrNCo+0lGCxmDrc1u1t2N27zI+UBlcfSMw8gVJE4
+OMAe4fUMGRFAUADkW2UU864pgwrfU5PwW8lChp+QB1ER4CKNrKI0Jmsi02u0m/vtA1uxVqiivYJ
49+VwN34UFnZ8jmLlvfKCkvuAkUmy/lAZyzlP+mDGai37GsvTrNkPKZZjO+g1V1Ip0MyPbtElPJL
ti67+rh0iSiJCYNhIpgG6V21JYyVW+u7HwT60EfbnYd+cWPRO39as3vmjH7dGu2b6wmwRP1YFPEG
FrvPsq6be77myMuOOX9pecjYEBn0jaalVB1lD6yzeRWKkb3fFT4EU4X7HxPPVpXSiph9PDabw9AQ
MlQT3lbz8W5BdCMGZXUoLD8qjs4Fu2250c1gDBHhzNRWp66f3ejnyorG9r6iTfjELTsXo/jCTQhs
93ep0HEyFAzSXG2G6CsA86wi9ioCZ2B6hywwxxMRipzdC94cXMo62BukY8ufTrI4XfeENbUwNy+V
v4T4uZTLUjM/J5aPqwPyPfvTTrEJsEojqjfYMVbT+XaI5oXORd3kTjyjpeDCeVqPAiapZq1/T3GE
B2EqASsIFto29D0UeKfMnLGZf+N4vxX5jKWxC0W4HUbqTO293wJKfkgHOgctByTzPl3mNW9XOUU5
RBX5wZlQQaYqt9Nm+v7ZCiCMhDNvTdKjDzcna+/DusskxpRGU/VV7Tm9B2BhGg5uXzsAa+8UXUQa
ulGfLUyojvaul9J4Sa7HHgBYU/+oDx4+HUqPCp2PLFPvdxHOcaAwR5J5V0M6f3IUx4B940jjozH3
VcKy2HCPQIrrvgJKkbbPzxOFsIud+ycmLHc4S4lmzBhcM5dYlhP3sTuuXV9t2NlQhR7xVQnhh6bZ
9aoBxtZGExNxuUZZj0UsJ+6t007HuLrpP0zgi9+WiZWnZLyjO75ZR4tfpFmjxaTwjlvLd3UUOMX0
tCKdiqSfOIsZDy/iOqpwVjssij0EAK65KbWKotH/5MiMlmXv83Ovgfiuy9mGagPlmMMLsb3q3x7g
sSGL8moiinlwx15xwouLLsO/A4e7rVbELMR8FPbKl6O14NN2/wDHgmEvU7t4lstSUBxn6MReNAaE
TNKokpoODKR9yZDdTy42f47HPioc/SluRsvZwmoR4a8eVu9qKJ78eHMXxU+wYuqtSfRbdxELeuGm
UMfJCjzfsYm3hC+Dl6GSmeKAvvqeXNwHEhnqKFedA9q9BhIyguSUx+6ql5p0TyV4tLmPe1Usnxep
qac/rYeNLiyxUwE3lxoquI6CWw4AcMdq5sYOnJzwE0La5W4f/Pqr13BGuwjc/i5NMYe9kvDjljs4
eeGAzt4nZP99N+dLJLXYBDjS7GCW+RhmHzkwx+zFHa0SMqFL9dFq1grVYXllX53fHtxgoD0l/DIB
P1P2gW0PcH0BhUC/jePVivSylqGR7/MShyZXgf8GD7x/7CdUKhSx8pNaiUAw1/wvdRdZnkfDHM6d
g81h1zBYHM6ZxFEosE6HKfhWVaR/1Zwdb7JLnuz3TD5F3vaV5bGIg1O98k/0YNK7HS0qSArXHdlD
VCREhyoDgM6fplgA9AXidI8kXyBCImcPdbnAnE4p2fmlASqcRWduvbUhlWRsQpJiyPtZF5Gab1yH
ORVJiaqhBgRP7Lfg1mTpfyif7R9VUO+o8HnyfZquDb4oNUEenm4EeWD49jfUGQrTb0lkBvPeACnN
J4nT1MTZmhMI8/vazdgxc+B/Fiv7jQtm5FLEUL5E1BeOaD5DAizp0RP4F4bO21b/gVCok6qyINtw
Q+UgJfM5C3bO0SLt9c6GeqoUNYEFELd9nhpkpcWtdAzrNxmSI0ubqTxeMwai6uXk9sL9NaIRMAmH
jMyAtHaHz0Bo3WfOFOY6cK/ZPNsxQlH7M74mUUxC2/9j7Ha6oQoEFzF/13yQDijnYIYHrDgUOwy3
PYfnmaTc1LCyapgiGb2t62hO2sokO3jL7ToM8YTKmrNqL/Lp8HXx2XAGb42dW5WNDwXgu/aHaAlx
Ot0jazU9ilWvMapFRK4HGNCqMVXVEV9UiJCe6Ge6Qq9U7GQBmGwRtEZd4Q4NaCMpJNJkSvzs7PBH
iFCwsbzuFavFicoLAh+wAAzdx5X0dqaInNXrzdVbHiBkStT4LHJxxmm+aCQCrZ9m3MJqt19eFihE
RcLXSc97Fga5RSx8nJ6FA6Rh6YSyZDjqInn0tyNTQsMD/MGr9lmBL7sCPyZsxJSyJ4QcJqLc7wQb
3kRAwzXVPHmoMCEsbgcGWOULLq5xmU2eHBUIxUpX4Rgm92yDaw2c3CRQdMzlsLE1wZMi+L4PioFq
IDVkKvmEXNhHPQRBDZjYhit4GO3k9ATv2gh+uBULc+P5HZZbWRTyQvbXfbdwzfyjL4GWKiyp9mc2
klPHsE4g4FsuLqmkolvi3dDR4n7KUp4uM3F4yKq1OgouBNRJyInrERmRBaaxVAyd5ojKuPlktlfk
pLXxppDe+pC8glda4KxPs/yyacIxfOdhWQnMS9XAezHpRbKthJcfTQHctT7hYv8uKDJOaRYr3GTu
8xdTaXgxXV3bRw7ht47L+twSN/OnYBPMFidob2Hi/e0LY0FoX8ASpJh6GskwiHBOPq6zRYhu6ysN
st9xxvqKVNsBWy+AlEzbbC5F94cjur58OioqI0fPe5OBmLTc+M2FNWrhJGj9I5ARIOggX+P76O43
BJI5uLBfVKQRbI+XIa6S6543hz9ZPTLDepdJo3mpSydQvpQqwG9dAefEk70RDRbZuqORJwq73Zjo
JLAuyOXGhZoS/rkgAhQgOIt3FZYqG+5BHRYzaKJPZSYytK9PoEbNLGjgy0rrFPj4js4QT1nuKuo4
jtCsmuSCvxlL0aPxDgHBHHRTcQmqvRXO32aHT31/3ktERuUnzDneCPAK3fEErieBAEEJLCQ5msZ1
40/c8j10xsM78mWOKFcCjC1MqMJxE8KWbNgulwm3plXbOAr1ZD0z3nr4OBwD6LxbnkleoV9smwrH
MwvdWkIhTu4ygXHBfrhCKQd4NqLgJEQf05/KO+pcr1I2gNV3dSp/Oigr91+92w+SqXcxdPwrwtcP
IIwcWdnrzkjyav6Mk+H3iL3cfNF3CIPHJXnsbLrThCqing9jRk0vls0+6SdGunk9YqfjCTF2hZnR
gUIIiVq8dAwQg+ZeG1ItDO/zm6wA9x1jofHh4GUFNMk6ImGPLAOPGbewXxoLi+tuCC5pYQ/7LtEy
qJzyWrkuQF5/uX8oYI0xf2qSU6xB0sIsNvGLlI37WHhy8RbQFGJU0z/su1+mMtFAIZPDDdHJC30E
4vO/Z2TZpLgyEbJJ08UdFwIN9ns+VCWt4JwKfNh+PMRXC4kAzdfdpPEM3h5j+eebEuVIwo+v1t95
ty8cZeliCglgqGgPBTFsED0/pORdAXpIq6/bS2nPAh2abRQGRXaA5wqdMSeMtGXYukFo46S4igoP
3WRN6CZrCoiMJ3X8trFgQYldtGfNsYxLvFzquFBCMdHv9MDIB5tuB6pM/ypBrYLCwvfMHynPEjy8
AQu62rlRtsXhY4g5vWe6nsH0JM477Cvimg/zPvqmGbnmjG4xfDqapbaFXysecCLvHDHB2Ybb/Ax3
O7v7oBCAF+amVIjdt1qX1vMk6b5w/9ouA7gDjQ/gsiB1gi3KOQLgC5EtF5V5WbWhqIoPv3kzsxJJ
f9TjzNbUjXz1mawKpADUPhHVNVYXr4z7yaNt3PJtAkOjFPvl+gEKcHnGgrrtfhTVcNG5+1yjMJWh
RIT5VxZoRe1K8N5+U/QwRzbIT1yxHDxbrQCUf3dKdc0HFWhmpTxpX5Gu6L4ZtqqcT+KpDBdWWT7z
oBbvHZ9H4Dw5YUM8wOWNwxtI4reY9VtAXn5ms0UhBNWMWU1IiEe5ket0+LmJPC+YmsRFk06S60Ij
CaxW7Xij9pxjN+tYnRadspujYTcPQ0OgwmYXafPs+xyYs9WnBZ6Gu9qtGFHddv1o5665rbYDyGl/
WeUL/H4Oh1mxaFfZlX2Gf0OijObD1JHmyB+w4Zkcy5eGrTfQjz+KAveV3BvLua0I5kLZDDPKKzge
/mFmEsHQwXkfDSiamm+mUp9QHYEH/AYZPqc+ZHCpUjofXE1HlpAKsdelfS4dZH2M6GmBnlwsYlW0
O8oKrtaJ6fhwkZ4YvkGltwvEuMUkdmkee+S4L4HqCTKKeRCVU3qW2eHpPEtVVv/0RRRY76BDak0b
VmP4jrmJapQcv+pnFVOCI5Q9KDNmlTP6rFGUjVydUCg4tjYF327vONEh9m7ovTQv14NNoPanHdNB
THOD36Z4dIlZxazIsQCjZuIiyFK00QTg4X30Ipv1TIcXCmREzIV595Ez+tpJ1/Z1/NPAcTtLvWgy
2EDlplVsxfr83c1YlumgalcomYH2rNzUtycWhTJRFXcVT6zSFgJ8As+gJbAbzML3IXojH6Zu3WPX
W48M9Cl95z8o1h0mfWwp2WYJ9w2wXTstHbf9pMZPbp3YA61nT5czuWDYF2BJdp6hun5M/+vV1x5S
35XJpIU2C7rc7gL9xWMZ5sZZB3NV9DS1a+uwPkKPYE2OvU6Sao7kadiDt/bYxAlOR0WCbQFRNJiC
xA0JgXBiekr6vd0ZMx17QfwppOP3kDCnzR8TwN9n1XcgNMQ3YoZeuvDdhagR0iOFs3FWe/9HpgxV
X1PELpQ6BiKcJ/AiOJH/T/QSJH9V2VWTM+n0H1cSr5Yynjt4s3y6sQuhm8I24wd1VjPfyaZ8n5F8
c+s7d/41xl3Bv6t68HSwezkTZIaXGAHhrnE1oBzWFasCl8/le1P54CqMGKk17zS0N2M3ulZrtItj
r8bqCu39507J7FB6SJlDJYi+UDQm6LZIcy0DyiNs+Hs65PkUgJShFLBcRhqeUXhonDwU6KSDbr5T
FJgpIyemcA0qLYwZB7e7vamHp8xlrmHn1CFlGqWlaatCtOQo/WdwKsWTg0TrGrnnUbpZs5cTV5Ja
HI9SlZa52s1BgM6Nyo6eQv/vMXOvYC81o6ZVNZCx7PjfyJYLCD+YHzhgW+P1LivWrKOIcHTqOmfE
MJlpwQE/BhqIuInUwEsCHBHmjl1dpw2ok+n0bYbbr3558mvPNKJGoHfRbDwJpWxybKrmQXh1AO3o
ULqmfz5Ygi32g5hlp/Xw3HiJNT+EXqga/tEsJ3fYBVLF1Jzn42eALqyI9Pr9eMw59QWUzSZ8M1Q+
5Un2rWzdGjyRSJDgwq0MdZfHKZvZve6fXhgKV+jE86TnJQK1XwwYkeFWlXiKyUFt1y72OB9pD6+S
kCYPNSlC/zJ+AkFHlrM6MSMrQZktu0TC5FGGuFYuXP220SIvwKt5zIV0TNaj3Dgrs8f8Scb/dI2B
5H+nwy3UH+gdgg/W6+U1Xivq2enuXBdmttnt5s9/Hfvsy0m5bPMpJYqeKGclBxuihxDDnGc/aKPS
tIbC3mlAMzbOoSCGs+9Uv93aaBnYeDCKbUI+rGXSQpjCuJqospvvCX0B9LBegpFbMOeMZEIktlui
gVa+vOC/+mwNX6cNFSH20+4bSjxNDsWhlXkbMQr7HcL1TTflkQxPoYbXEXBSBRXd7I+ijVQOnFNX
5oUiUEYOqWUq4DFKd0Mp7mclfqTzF54xev6Wh55qWhV/JlpgzH193cssyOEw1RzpuuVmweKq8OHW
6CDQS0gibttPi4Q8laNNYkqpbU9e6BPhIqDrTHgRVTbgWp/06H+vy1U2pbJTJ2+2qcxRHGNBlFrP
Wby/fgmBC1mBhOEPNtntUYWB8h9PQxXEc4EYFfiDlsJn4eKM9X5Dl1QsVIZLOl5LBEv7Y+90SGCK
wKnW+WPIjJ2E8zyMmwyBrf1Y/5o+6151Dj+uGmMm9NFJ/pN9N4K4mboU0vnC9/d4Nl/0ktNhUbUb
gQDm+I0=
`pragma protect end_protected
