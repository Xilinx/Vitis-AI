`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrM41f83zxdpq7B9Bxc+63s/ThO5
lR4ebiIUudrMSnsXzTRn4negwrrB4VipTwcqyfoZbX2gIf3gPwkP3q41DFrLyf9opSDFSsyylvuq
0tfuxhMWxI0KvORiuv+DLG15sEi9Zilc4jLqmJBgxaj93813ixDm3VBlIU1BQYAYzQ6XobruGhlp
W7l+H9tAQt0BvNuSDNd6KHRHtkpbBcXPwpTyA+6hMW6u6Ccsl4qsUag/gM7FTpREXGWubujKpgQY
rp+R3/RbOFiTkF+9XB3PcW6M4vfJf7FuItJ+TUqq32GpP2JaBAt8HeQVKtrTXfObKsVLCMwP4E1R
tyAVw6rO686N8A0sNSdMyE3pASDfGpvlX9QqICqK85Ft0LJIfsOMiI5tZ7dP1zCt2f3oWdfDg3EP
3lItKyP1gfL1kyFw7e99tktlJvFsQSrXdzh2gyciLJbFm3k4DyOeX7bxSb3YW8qj4NfuSDIOhHtG
6sVeBYqFfL3gXy3NQAT5ANAP+18upDCmKmlSgu0+qu14vgUrzLQXvMeMCAmemGAy4r1LBuoEn6lV
jv7oGBg9rDLP534Uwv/DomELrr9KD3/QyoGNVW03A4SWoOwoQpODoxVqTv0ZQ1PMc5tOj1KNf7Gi
9QcFqUL2T8FC+7DgLFohEhJ6D28PPzwOC9oneoSTxGcSMXxJBnoLEV9bWjeZqNvtWYtND+AznsAO
EJEHTOW/vJBU24zurIg0oIjT5EYuu+IP5uO/QVUAKhxZx+bl/+cRBfSttM8utJRIPX2QtywFYRz0
TR0iyd/DikZ6nD0uTI0Do1JsteVsggJYg2dTm2Z4Br0Tqm8lyulsVA3WXo2kBuI/0AllhZEPIRU7
HcFX8lTKCvp1CDnOZyZi8uQqQfZcNpyRKLN1wV5VojfU5wxF/BePgtPFytaRZAvz246rAXl/kMqG
LsLuhzoqZadl4RZ8LPX5I0fYebkJJLKUQdhYQYujimaqq9dJbpmMY2/wYEXzS7ieJuPEW5XPsesy
874i4AAbY/4NXmA3J2x/BNYt1QsDYDugsU7981NIJ7PAhHlvo45f5McSAH9Jzrr/4ya6z5j+6K3u
yHpk4FbJvp+5CJ2rzdtx8A3nykJMT75OJ5Lb41ln54kEoPUjds+SK2jyv6kkBaKPUwF4Ue3qbB8C
aOYuOXvAd7h4428zfrF0Fm0WuKbJcOmBu/mOIZBkh5LifzQNnbhNT4Kfs7+sKPOmTjbLBT1fXR+W
RtM+JZBt3edbBO/oDf1iiN7QqJfvMWYbJiOIQxQhulgvFyWxI7AcF+XK3MMPO4GLJ5ImZiv2ldRP
UEzRJbI3hbMwZtJLou7z2a8FzfS/hgaEkXyzksEnRlzDdLbKVIN+HUrBrYMAmXRk3oeunSS7PmUh
dNBstgFzrjuP+JRfM8PvrqKf2NRU07qGRAjN/pSb1Qprt+1eYF/z/s1veAgcYDq2IxTIYvNK+bPh
OSNWLFiNLTJomLKcBCo8cccz0D28mkskdFjShLYOSdaSJjSvNZwcbCPx2n47PZAEnpdAKG8/ueSN
aQM2k9O66LCdtjvfEgn0/zEYEQbDAk3pEUYECHy+Y69VolX2djv7r0eN2tIJq0gz/1D8m1O/aYrA
7Ld11FCHQKRVFy0JGi47fF7MvBet2gaGgQmUS4iIFnVGk0M6nEUymoO66PLObZhcI4OvqaAC8nHq
pHasYvYkwn+msJUCv6oau2OgiC6RxP81Ko7dw4Ire4xIsBuqrl7TKW+/Hf2Ul80IcT+M8r5J2NRj
87YHs6qqjC6Q87IbKA5fxePUhQlx/r4F7rkfnvOP6wtQ5FK0QlwJAvbeAG1v1Q6x6q0IIuBeCDjt
BurCsgo4UossZzlYOH5lp/X16/PDUAs/fzvleRl+qiTDl7zKVsmnYKTAGWdP6SjKwr3VSIIsbJPn
MH7xxbxOGCFXny8h1yJyinBVrGCHzyBUJpsVA2B5wnup/QcQ9CKpvmnfGzJdXv56uc4rTyZp9M76
wG7eaOrm+yX0y/huken3b7iGcu/i1Xev4cXCIQSOdxf349WzM9e+CDustcL4XhWmJWCW4dmO+/T/
zJuGZrk3CT58Leio+x4gOWEVT9Vs/OV4hkjIOE7RTK4fh+qsoNMnZ1hqhG8qwS97LBdlERccZheA
jpu7aUvr+yY4eAJ9ReoAIJl3nSzmMGNfCNczN/A+Pc+6IFVIcKIoLZ+SKzCHRVn9ntBaTR41cIaX
QVNXeFdpZF9pD5WEZyOgxif4EQ3g/YpX3MIOxlcHaz9KBda4qpOseETt45Jvsao0ahCIdjipStjw
utrttgoCtaPpBLMlLlgBDqN5Iu686pf80eTzPgBoiCTOtoyFcEg3dMCabBLK05ymhIqw7Fg2xW1q
V2ELUquJOcfkXkJEI6efDeEXxPMUVdXYEfxq3fo/+IQ19fGNmVzsgaT23yccyOJQ6+9DwiNsQnR2
43W9j4cDEmqZ0zMNb1v9AXtfSu1WAb3RfXy+SUygZl2CjUZ+bANHYTwKg5zic+r5GsWFcsu/xldw
hLQswJMAh/Syr91XJUr4b7BalZG0Izr/xdSmHR/Ms0EoxBuemMnBNL0x6oOS5ZK3XovqnrWMGjVm
rsTQaxajRhGnLq/f/cM5gxQUuQhcyhIUkC/25JFhDo0X+lmQmX6T2rOxf7HLaTYJHpQl/O8LwlaJ
/9ThhxpuQtRf5aJC00YVAwKGqzmRvg3jfbkGNV93qLXTy2u6OJj9PSiFRVLymdlbXTnNLLnkask1
5IKD5MUR7bZKC3G+kDlQ5II8F1mTnoAwPQHxPXKiL7Kog2YD+j2rU9GO3h76SEkUCCjlynYUA6t7
QSK3Xpkq0BOeZdLDqoIP09m9S+dVgYzlKw76Q2hj8voOB+7iAML2cGwDV8cRjksvpkBvPGt83E8N
1/k5HyTCVZp7f9QLIY5hEoJvhkdKN044irtchF8xv8yM2PbAbfmLB0FnCvCBlAhZPK3m2ZVI420R
mVN0814n1yUmigyeXC32eazte6nlvGcqxkL+3cfE64t6sOAVxJnQK7kL9dgzk2F/IRJSxYhGWGZf
0yeUgO5000MyOujY/maWfLIJ/bDBg4TBWDGf6/tZfNJlgSaYLC3iaDWn1VsCAAJJq5iFTBGLgMve
kK36KTQHCKIbc8hC51ps7Lhzyx1hxM4DUCIDCTDlSYLO311BCrTSCHG+S/IYqHi249cQ1w9owTCK
opnwDw5HOd5+PxzlmALKkwSO/59fBt1TnY7APe+WH5CA/hg9ok3TcVGqrphe5QU4yc3OWJL6aATK
knl3I2KdIgSux03svE53mt+mrF4P72OgtVy9tW7EOJtocP6efaELWM/tkQV7dxPnx3GbnlKK0kKy
aWduaMNk/tt4XqqGSe1/vdCE8yO3ABqQ3G7ST+UdXIKXNBDt/lSDL4X9hpC2XJjM/ydklRhRSHUN
luikCASOkFzGpAduWyQRT3e4XZFkYgwCIuSgWddO1P/KjnPUSTaA0ibSSE9gBuq7sNpk2hF8JqJR
Uaguc5VssWE/XLpn5DbrSwMAkSsyb6AZOgR6ouY1bvUhINEusgGJzCF99nB2oh0fTb0MMSaMh6Vb
uqBOKnedUfD2XvIxrpLJo9HAqleZRiXq0i2XaBEIzCf/nQZbzYKgDJZcdGuBZanhBz3CIuxBOTFr
cWnyZpJgYmgGuAqAugDd1SKDSGxJGjB1ds9QtMWa1cJF8y2q6zEokCCfQO1B9F+uQGIRfwWdI/Xw
pVSOZY4c5dBKnhK3D/Ro7d823OLyQFmnnuZddTDGPQGC668wiUgNdc/I4xszRd8gxwt4CIkZf221
tKZNvYbm1oKZ7giOpiLAH4R3tXsomNT53h/E1fHF7rEI1zoP4GoO1ZEUUjQH94DlgHIaERDp6yxn
Z2SXXtElRVvSs21AnqVd4wfNyZXG3ad60CvwZHB4nSLSoC0tSFblwXtLyyvDbWk9RHm+8FmWepO2
XLsEZNyWqV5Dak8Nc1G8Zwun0Nbo480IViW97v65v1mEOEvKNGw3PxYX5f/aThExO1xYhKXcBLM7
CsW8C2LIPi20UL8V3SkVvU2wSgnhH2+WJKUVhcZiq96lj8M6WCfGyB+lr92WHr4VPwAVw9SN/FCO
x69bZ3zA0VVlWL4MGser6gqzqkgLoRnVXO/NDxr+PeYEVY/hhF40eJQ7zCi40N2Sc5YZgGQ7ucXK
PSgrkNUb2VNOHhrxu4H2ARoG3cic+5V7hdn9nhlC9SWbUbP7y5PaoYx+fylJkE+qZvTKUE/gaSNG
lhne1OIXqzkhTanj2fhddcD8tUrdiYBANwC9Y4u72B7ED/5458BZlOR4Thtid3KhpP3/K8VCPwfI
c6Ijrg1ZmIzBwFcmfv9vk29iojex0mPWsaJLYclMj54ChG2STVH9Ai3zK+qygyVOFKZk258LEDnl
KSEumQMiwRLvHrkgwa4p+hgz9fnOpSLuw4P2i0ubmxGbWp3R3s5ZO0w683fenTyRbjorBADdZSjA
aCTcwTz9+hbgAkVof+zASRXSa9MFbUEatWb4uQXmKadmNa7KnRYjNCRVjdB8Y3jFqL0emVAoQcFh
l2Duod133jzpsmCSa1ty/udVTXwO4yFcCh7WJ+3YPgMySAtTPUFTRMGRqDhSl+S9fAwUQz17lwCG
euYuzGpaaPNEJ/0hxBOv+B+hPWi6LIilOuzCi+0y9o/+lDb1qm5wUTlkKgXKcs8WuRJCbqTpyHJf
MRZKXv9S/a50iV00xe4I/z00NhIFuXSkiVYUIxWqXhEjhs/AV7kZ4C/yl/ewTGWyQZcsCB/Kaja4
/fdQaFi0xMat50zrv4dkjJKcq1KW0O1GgYAQgHBmGY6ny63pc+EzfnTEhqDtC2LFnLbQaFVzWwfQ
PC6+rbVq/UCb4xgDq9vFBXiVtoJGmYUS/SpJg6qomfjrJBFyQRduSDRa1O7VMdWxD2o63JeqorPR
HaoYltA7wjfSq6ESB9IgnB8h/FC/hm+QknKkDVtvDh4BJhEvG26sfrvuBt2mx8GqUpaCLGgbv/Wp
VaXFGWPaQI4W7ghhcmlIIvNe6ZegSBmYqr0YBBiLoidwOKpIoqypkk3AznY39XAa+Y4HnErrDafF
4tyIpItZNTjWsZynNhOLvMqEiCluU2wFMwsIWH2v498jjLLfzdy0Pepwr6m+lkPF1n12s0nIEysK
Xrr0ff8KhoSItIe3bF6UOETpyFh0eP3rXVJElwFwfODBFa1qzlAiYeE/qz+zEoXVtaRlDG3MuBbk
FjzcAKoeW5tgbeuuK8c36dOW/VkUW/xKMYo+IBZAB2rEd7Czu47iiFAfxLe7pvi50kVfjsjCfE+k
9AaFr40i3EsXzkKIiMxPgc5oSOJ47JuDm0ayF/CvRw7bKZvyXf9F8cW7Zmvq0HSF5kfmaT6eeoku
zKrbOw/k74ZisDhQsRS1t9jb2RU/yvasY/Ist7UdE/gq03oTejCHv04ly7X/4EpxyziHUp5kury5
roFiang4rHXE496BRsI4/vpj+PzD4FN6yDAP8B4ebHijKu60DA7HYmV/1B8Cli9Ke1NnFwgcSNfI
mzr4jR14IJNcX7IAZIxRVVLGIAupk9NfZANSbUFbqdWY1VL+7wmY1wP+smK8NDax4EwIJSpfeBYg
mp8bA1/Ticht9yVDOepWZDhc7ekn/7Ko8ZjO9Q8+s186ZG5N3CSmc6M5pY6E7ZEczUy0flxqt9sm
iZBMed3/IvWyzqvSlhGSRSiTXs9UKL4pSLPLLPAGHFLKKrDh5NDj1gNsB5lizo50al9IcBeTiecK
G6CcZ41xTYzpGgB5oWPzWyrYJMLeKTaoqoYoV2hlXlFqTWGbCKSgVlcvPob0mHwJdch9Jrih9AWt
yCJGIbKIAOm34VpREwy3EK8g+/Ze6TRrzszVwZsPS/6E1a2yPk7s/lBY0zwr1ZDtXaOGpUMnEYom
rIRLmWvtd9IwqKdu3lofrRv66gUsc7zjwdvurzlJjO/Vd06PnFFJvcvz4dxXeY0wiPHrIBdcToiY
vsuN09yRLnt4mSV9U51wZ0WuPSEzKQ1Hwjf46BRQFvc3IPcX6jUro6GlvrmwmRAKZZohqlk8mWG6
eVPsnjscHVxuEVU0dT+EKP8iHPQBQjsjPfnC/P5+XfWfWZtgN1xs3VV5X1tR8ozIRYaKgTT0mVfs
X8friXeiT5VDOKuhYdmgXGiXqjqTYtMq3S748znAVtfNGVb5cKBZtq4FFSUGaIRaGsXg8HO5TSsz
5hAH7F+JYYbl6Jj39f8tTDqhzU+oOTuJnQcyil8sPC/UyW7/lvC5sZjk3LBJrme9aXdcGJG4ccAO
IjZY2k/OfkvONsL5l9gYGl4E+W+ycW7nyezh9gBa4a+nNbFFrPT/1tB34Fd+QOMMbdG9Q4AiHkMj
E1EBiG0Jl/9iCeV+43wP90eaSNhfuLgnmTlQtnfjAa3GF9jyPB9N1Rf107SBMcqTUCrtzk1ne7X6
hPDmah4fcwP4pePXl5X73cPXKRE5p4bgUVoCKq7Z2+o+cGWn4W8zYT49d5FJwzJexNqvbZNixOYe
j3DlJjqXS0PGY+9M+CDQLJ6CvlnGgBbs8ua+5YFQjrVY5t++Fm5mk5rB6+SR3+4bjxqCRmOrBwlf
9zU02l8URHQgFBLF04EkHvU4nphrbUN3yUeY3kVfVEaSgp9QSh3MJZJBLOzIWhgkgAIsb3npk93w
R26z+mJNadHWaoX/erAJO0LbJOMlb8pByaAxxNs91CG1Xvi8CBwh6Yw3+gocROEJ0hI/3A3GfVUG
M/pYSIEkjyOMe7m3Z237bXVHXqa+TecevneD+KQe6Gv4iw34gC+BrfbrAS/iTjcm0eAEFV3S2JWp
hfoa0lywkTr2g8CKMwkkoNdn3WTpi7HDK4hym3cqCwn8HGxncCdTngvFgNC5XYbgyH0AAuak9+/P
XToXFVyBlLrwD27sYuiU+WlUKE5gtYQuvquCr6BlPMKmgZSK+PhoYWKPrsfbNROmc4eVTz0TgErH
5aauDi8Rud5fL/T9kEP62jEqWf6ryH4KMtQyIjhiwNolIEcH59ICFdWS3TvUMHM4SbExNZ2CaNhb
PaaH5AGVBV7Ga0KvrsFC4UYYRlmAXBXGEb40jOPttxbJreuf+8cRGb4JpBDAwyvNPt7e12zXQndl
VFIbYCRXAwfGULuKrdMITf8XDNZGdgUQD31DkfEbgf7xrnYWfkLtlGCEgneibNwmjIZjtbRhAH7r
6lEIm1/1+BwJuOiDxKBTiGqnGa3ErEHB35sCuw+91ED6ytepvHTwDI9X8x9RDt9mLUBerCbECAsH
si9eAOTm5Gh8AK/VE0e7R31rkKQJ3BT5sjym1ZSvWMmHWIqj/f46bGjTZw9lATYbkCOjyaqzw1FT
a1XS2EY+o9H0NFncSg32fbMIfxmrbrh/J9B3SCzUVRZU65tEgTH99mV+yMRmDUXEpYAFTgsL0guh
acWTMdFEkjfrzGhJlm9/tSwVFL9PCF92hle4hnnJOkAZA4DcZa41IJ5ptDDzSG6rnfgCy91ARBKd
jV5scZLdHgYnXYFFS/+SBjBghMGvz6lCU+ZNTLo/pIIGf7O2o0RiqUOsYXPqJdd3pE/Ehc68hPC8
UISH5Hw8YAYhlVkVF9OfUSDvjQ+sMEfegSYwNUnuYC23OkTreTlY0lNusexVyPabzZZHQW04c+iK
FZ5z8DRia0XDWZqcoxCKysYiqYI6dNSARxdiK1kZB+Dgig6Y9K9xyD1pkVthBx7Y12pStc8rGwrL
Sj1cChrMKAkj4e0c04HZK678AE/uEkG/sp6gnvljLOoK4J3vjtjTJvuAq8FWg1flKF5AhVun/wN1
QL+bfW7EpRfmbM8DPaJayaHYKXLKxswZpi6iR7aZZKmlnYAcil55Kgidhd92iAoBtFqtutXAfRJa
CJKQiYZ+7btfbNBUiLQoC+jXu07fN50Mv3+2jNXsDawFUuMmGfbGCou4w53AW7bywm6MZtL7+Smi
8aizV60cG1Hq4kSF6f+sTckZ815kwuFT3Z9wZSuo6N97yw61dWKPRNgwB6K+h0FeBmEhSjg1O4HC
1tvkJ/menbM3m0I5gCKe0erD+Njljq/AzR6EHaZMdD3at5baS4JJORPRxPRNOuZKOOhjmOYs/kUw
hXSrx3UUW73zzL2SqaPU+ovhQetYdlIDARRs1H54kAJFKHve7IRS3HdD4TPxzc2WiGa80O4PHJvM
Y0ZNjIW4Mv0P8/JxS5gM+OFQN4k5MRf6ZxIL8LZVdn+t3zcGxgHYlCdlWkLlUrXDISDJoQnH7U6S
SjxFTfJLt+W4nKHtJ1rpqifdIx/smRs98DgWZt9kpONOaTRJhH+EmcxM+O1vSn88v/5y6YROppMt
fZi1phqgaKuwjwFbAEa2xWVzHsaK/KC/VwjqaVOgxxvjrkDKQdpXhwuw6y7HU3vyI7z2d/iMNCQj
wzlSTRPDHzyNbt5B1JJi3ziXoHTKzvWEku+ThQfGoU0FQzEtUjk7ptHhVvmfBsKFL/pKWehvLg4T
C4LIxcP8h/fgzY3q2cEesYO8Py5ohqfSrcXv+1zm1MjJLd+7eBGcz/l5/J8QBd96M5UUoQKlyor4
eh6Vtr17L8Ifd+xP1Tdr4GThTzCIAKD/kg2cRrUXW82QEm1BIQfNjj/o+hJZlhsfKEfDuJnfSvvb
7kQtP3qxnKjm5d0e2sRh8tozsWquBS95r6LReOZf4fLJUkEXlh8JuD4m3maN2UNCKgSAvMvGF8aU
JpZUJOmNcqHQcU7J88YjRNGLldcRDrBYyiCh/fbQbmzdeOd7BW6UgMT3sF1JVf8vyk4brjkqLwvF
124UgJjzUE0jK1ppLUajza1SYVkNKAENyLv638508o678COuwzf1hOB+tWk7ppP/PbqaWQ4eqVDE
ivYJ8K0c+Qm2/pGXnrFrcdh0MZt8SPJ6wHVQmaBYlbv/zEqkSdFoBFVMto3tY9RedB3G0j89D+Oc
qViFl2wB4sYXWfmaKONHK+oBDooFbCuiAwyWBchOKe90/WLj4E/bE/E++YTCVP/BKXKCMqlfqcX4
8dQul5wzFM9L9MON80ofVl/nJEGGgI3Yo7v1/Ne5iI+ftc41hU5CQI3jpPXsYTbpi6s7ub3i38pm
fJ1tyn0vFRXza/3rKDY0FPGneNFWGfM3dKj8b9dvsEraKyzjOpL7a+xXqlP6PlKuOP59TBlgiKZi
JLbIPfFLhnbnpYJuia1/iPl+lPdHTR8yKYwtEvKO7+GYLVvnFvvFVwP/aPE5rN1UFHz/1uYjlwco
fP3GMkLH7vTxaACVMfOYeqHwYaLOy4maD+OF2M7COoT9nTKpv9T6qnUHr9LxH1NGF2m9b/4chJ9m
DEGyMBBuLsRAfr3wzaKQXzVhL7H9I0WYWrZKv30K2sEXSP0CLd2lAZxVR6hcVLwGOIlse6L7ueF8
c2O22PIR/HUWeoIEvVix6rYXQtlGavxMoh9sx+nfXJmnCS3beEYLDG3MYk2BRYiKs5DAR5pWy9y8
hsXtcwzQWMPER8v0DJCu4ApUB5IJ8TrPMssaXVLLIKxOLu8hM91fBPOL8d7LnYavCrGhadsGtt18
/IRyHgj5cu5Tvc0R0x+3k9hML5NtOTLfHJsWn17xfjc2hHrpKEX3kEaDErwqJJM4FosHnziGhe6v
WZjLSxWmNOyg+/TsR8rtpX7stjBdSlli5fQvIe47KjJ7g7M/FCPYNgf8buaFJa3WTtF0adSJduvl
RLb/557sHlGBlrGS3ASX80007bb2ncz+d4eI3mj3vhfZcDCuLeDSQ/ABopNchOs2ru3ZN4n4/dCK
TvoPq9ZP0erL/pcX9QuxwS6U0OywhM6HnigI3LhYbhqAc+MTV0feSUbLU/m90ncmffb0ll16Cfwv
UvF1WPmtiqusW2xfz8puprnFgCZypyEa2e0ua7RRYDAunPFS5SqbLG/9c91wl9Pa6FX7TpKcXWDa
Vbx8x33lJCN+F2tsUDTqT6jbbQPF2c31wVFjAOFJlYN7CAKknCUZt8rY7N7NXgGCuSzePNHF3w/s
/ThqHuqK1o7Gf1oicVk3mlruDaSSSCrPw9NNkuhZnFczCh40eVQ7bFxGBDKcmJKkOavug5FCGcsV
jb40Q7Uoc1veUeYiGg1pugmNDFiX8S+W1yt/yVA7k84hU3gHcjTSKJJT1GIlMT89HcajMAN9iqE8
WOnQndjHN721iGRQuDwnH7J2yoXuZVqsdzEFTqvaGNW8EWpktLqh3sVnpHGoCwkNFZtzkvW2dzJ0
s62DDzi2GT2XO+fhm0CNCCmxNS4kAHIPSFRfEiNNeQEB5prqyjCa/N0eWuSY3+XvpVO/j0jMT7d3
zbSFlyphfMhn7WxGp7BSWiRTZTVm9aYzWUWucvOD8J6WKrRBcnwkSHcLwq2ifnCHjp7qdJ+pplDb
6HozkHl99ZcaDj+D9WWanVLl50+6mS6DandldP6J9mBxkLD7jiyDeNyS7yyFAwdtmq4nYWKzaJCa
IUAoMg9dpKuqPcDN6+0Qmxhfi2UvwfadXkJ5EXyC5IlX0ha/paVHdA4MLI8JoG9P0PZ9xmEzU+G6
+j027xPrQsbvDzK72YyVTLpiWzIINZU7dVJQrl/tdxF5HX0QW94r/egbbce0HxZk34g0JM9OjCHK
l3hPk5XoMdqFMy0ni7gausFL+ekyUlj8AK4XOwfQLjGmx2XQwClwdRUnfu0aBYed4vXRbyDsGKNB
tVnZabKEuVZPOjYxozGZN7Epzj+uFOz9mTswmpHkQ+WPAMbR6Ke5TShjCG7aW+eEryu7hhlmPcTY
Qth4TPt8QWPej7AQtlOMAnrCKLB4cYMKNoG0o/TUObd+Iho6NtK8Bm/fWrQmsMo2mA5DWLEAONyY
8ObpG7X15cUn21S7exF0zvtLNqBC2iF2Urv2TuPLP6+EbyhXaIqnPTbQiadGhYpJ3JkObwz4zp69
ODx17wXu7tBf/L/qPdgZYL06LsY84yjn7I1aVCSxlcDmnFC0KFgTmpEbSuhfjj81mb6aaA+aOIud
UexRoVYEY1wZgAs0JwgFfhMc4YoOPZL3kjk6H6SpziaAPg12vB17CATreqfUQNAFNxTZmIlbSJ7k
IYbaIqFRrs0kXjqvIbgaCVDJJJmd3J5wOf7JYrzImREC0bSUYT+yS+kn/dGLcADTzyufxog+fKKw
tB9QxNcx6/fdR/RWFLSwsMH8WQZkoGOeT8dKYwAnK2gtuKl7bSt+pPjUWF8iuewVHqHgaC/VaWPV
cdn9GtuEqWtAkfY0BKXYZ/3fuJQnT20d8dTZ9Ijsiv3ofYYxB6fYnT+n2dnkbWqcbKVPeJqq7t+8
yrrGgUDpSYi9IAQy9PhDOfSr1HZMlTwSrZcP/KaCxq6Wu5YoEKdxE4+ubWvwUIfyer/UYOaERPCI
8r1dQcQY//ysRE1kPcXpRO9BfeIhcRebkIvs6Hn80BzC/REUB1wl1K4I3yPwlcoyd/NdyZ7HdyaW
vFjrJ1zDzInJJnZAVH7Mk7DgKdzZ584F6udXQ/UjGu9lLtH0PMpDmyNYkXm8OiOUm/7mxghjvo7z
KqQe36/hRBtjveKy4mAhXLEOW/JCXuTUMG5tPbwjDDCnRcHKSS56heX2EJy/Nza5vNI98AQ0TVS6
HZbR74TlFKFZ/6OLg936dpjBIK/q/17tKw4qN+LcvX9lk1buFq8pd8Hkve7mWnhm9rcaY7ci5H6u
1wCGfPKyb2HvR8JdpcNJUTjCoO8gx1nyk9P15wKFxcL7DvIlmeTXkrdTD2KuUpUZ69xiFM+0jDaF
U3MXDmL7SCVRc1o5C0qzx6RDc8BVHEzXKxdOoYk0W+G7RkRi3k0eDPZXXhXCCRldwzyDEIdKB1tp
I7Au3Tlf67XSJ5Nhnbdp54mbwKWDhhZGHuZ5xY0NqSRnTtY4/UoWGh1JE4nYrMFIDL74kPSuGUlC
ug9sDeOKjF7Qe7YaVuPuou9RmtP+WHXDXstW8k21D2I5A/ty+dC6hmRQ54yxNNP6HuDNL/MC95oK
8JsUUJqfZStnmQXCzLexB1UxqK54zaDNS3uePeCJ6xb1SGFK6QWc0NBjwaGLfrKWY/5UrPmlQK0h
kF5VmmIPLA60RsZ5YHFmWB4WB4s3ag1uJkiMz+ujrEoQYYLQXya9ndDCxlhyf4gUdaGEJ6taWiqR
gWfX/nLGU/uUU+bxUVm9jAPw174nd5llfUuwe2hOXLJriT0B+JGhKDvFhvE1cXEP68JmDyhdxT5G
C/HeLpx8lahT+n5/Tb+iNl+usy3rdeMXdTy5/FNQY6lJnAbIiI9Nk3Ue7MsApGT9x23kLUjwHaMJ
lIztuVsotjVfhMpjf2F18P7db9Kav9RuVGk0vxevZNuwA1OKninsPgCxAWrqDlYlixajB73EoxcW
sPyC8KIEe4LMzKSfBrq6u1KyAsVXaPGF+n1L9GADYCDcqh6pCc4rdbmmybYpE1MgWi0gNjj/kXKb
dMR0szs/jamvpw+CFR5bLdssKZ9H9/t6ub6BO8ZhOg+BpflrGhjTwaI44CXgntpIiMkoz4T0I737
MW4QI/oMRFshRYEIfFYLGXBuLqOZRHycux/zOQNtfoxIcNMkwKZxvXGgW7xtD2FWr7WuOeUeCwfQ
5CAxAhplNeDN8ewn6ATO6/x31caM1b/24mSTZIkqp8qMlwahl7J8J4yymacLV9mXmokQRdV5et4y
9vSQvuqP8glDWL1OHQ+bP+dCBd8VIOgLFae3Sx/Cb28CYW5N+QrlJCTMeUOgckBTq0fuboV38lJT
rEQtdfOMkiaOeXcs13qnS+TjuCQRzZV2GZvwox3bXFNPNglDkzLKnmCVVa9bDJsuqLIGzN86ntRf
sQ/cHHHmvT9oJAne9zn54eftG5V7fzuArBVfcrIsv1vC5LQZOiO6DWtoJqANjw3novIAJV2qWJBr
xUeLy63AngCzT/DZdFhcAJRODwKy8B7hKWCGPgD2xxqNOIj9LeJz3vcC1CZpvAxKs62n4F83jgS2
G/8Bhb8T5uG6A2Ix9wJn9I8E7pjBHVs+34GeVRDz7l9HGFzQgGXbyHz2MeLUNfTLOeEX1tY+rEDW
L5Mml3nrthcQYuknCe4813PmR1LBUBD/NVYgJgNCBqXLP6fSdt+tkFLIyOPCB5qIozXrBQyxY2bK
+fgW6lkq4nnsEU3DHSZBTYG9IA8tdoLrmgRv41V1OdEhV9mc3+zvKzHEebUsAtOJspzeUieTuOwd
BHqKcg4+4t7XxmnSMrIQF8m0sVzgr2tJKmY45XV2bmcVDq4gx5tsmbaU5eeSmZkRakmH1yeIsuZ1
Z5yp+VMDs1hxYUneFQJTKes3oINKc+zNmo+NtLivRYuuF7dc+lE/bF5j+GHyrPrR4NN2jZw5eGRd
JQZk2TwpcG89YWILpKRn41VM0kzqvvorQHntoXbxuN1GjuMHEbgWplbU4wl7NuN2MGaSkjr48vfh
d07ue+cRTtkrtSPjpfDbNyxyqF9O5nAL0/yZlrlgfNH1HIRcuiIb4+EtFNE4QkMDBSSR5TOzUnZk
FRe7d2dLMY671/bTMCJBcOhklOjmfi5i3APq/QoKG5ovCS/K9dS8nmERZiKagY7q3twGhNUAXn5E
t7psJa9Xs32ayf68uso3fw/mhS+W/8aIaCj0KeblnCSMEK6bmvXdVc3YL4c6ibkIFQ1wlHp3Th6X
t98mBfOU2lY4UuLjtEolQJ26y3WwGGCVwNFdthkAh7YuEVH2hwsyWEicO4aejXVzoocaD+P3acuA
IcjMgocxKr4vuWJjW22S+crfMc1lPbgwA6LK45qbqXSJBiAEyxnrEZdgcPS0hIlnMpH4TEDjIPOW
Fd3uM2tfr3T5aHNSp1GEB6NONXucfy9W0XwfV8fOcYcwC2CXsVe6scOB/kkzyAdv/43PBBQxo+i8
kCCpZv9dScR4qtMQPdWs8Ww7c+kC6xouCvUofojw6knzoZ1iyT3vFi02wT+q9KI62FnmXQHzplEc
RGzOGkROtdujd45B6yZYrU0YQ0TMIeYQRGgdoyZp15KhJf8O82m2QmVS6425bdptpoicTJvPqTmo
l0QQ/7EvQ7h4Hxk2kfMLs5sJoWMG4dkc8luF7Xz9N3EXj8dKjx4hXBIeotUx4rFOnG9m3YUVipBB
k+8OgNzVu3Pb7YvS/ZBM6CaiMfE9K/HY39LQnyzQS5U1vhNhzb6d8mgtsj8umiCPwza1sHhdq2q1
gRLWyag9p8vxkv5hrOCV8dkfWnO2lw1Cj1AoiJg0msfNwhdrBm+KUk3OReDBJIrin9AY4x/bNFjt
3ar+sO1MtzbPddVsUfhruRHkTZJavLjcxTTkSGDm2H189MMs76fDF9kE1WjOqKG0hXeRABTC/pI7
4cDhZGBc82ROW1Yu6KydQUHUBX8C5AAwQerW7RWIKSWNVQiDg2YiYTHXr/L80n/Q5emwCrLCpLDS
wqzptJ32XSkwp4aMpvwHmeopG4+q0rrY+w7ohAlF70Vp0B1vGyhcQeOMCfeiAWG4lNO1fFZvTbXD
+B8TcFe5557eBLLj0zN8KnYGcM+qChN7EinPCtGXeGQBuFjJlDgSxdE4fu1u7alK0vyuqVJIvNvi
/l/PGiL3FqUXMfo4q6RNjFvD9Vz1UNqxMe08Wqm5W3t+n9fDk8LffyK40mIv5J9bT0ccJtiuUvFC
LeeQsdyfJpJDWX6pwwQeCBG+HjLVoVNBbT52ZnbZFNV9dcqikrkfkzq+i7SrnFsZBTOIfw2+1zLn
vLsnnUCmDl4FHCdpYldSoqW4YgWPjC88yFcqtaspfbFBzdpQq1ce57we+8qzh+qDwMD95gUO7g1I
7Hu2Gv01TW283inkhdlFMfiIj/iXNvTYl/lVRf53E8Kgw5ppUgmYynjnoejPBHR69Vi3lOqwBXEA
jhvpP/pURBvpNWE3CWG5ghqUG5mMbSE7Aolcd4mLJ3ncgcPlYvSBUAolpY7RwEOls8AfrPF6sROQ
/FIirWFpMepQcTIp4QTThqKAKAqKhzLBAsR1maWZh61A9wVzyQorZDTHYeLjJlS+ZZ+YS4htMyr3
17GAZqOzHuEdgydxKlnm5yTDu6BfM/MdBOLYoJ1hnm3kzIxnkqPIt1pmJQrPsHUFp3DOjR+VJ1O0
3CtIKsJO14eBNfJrKkTfY/2oq5geNPqB0gBX5jbMDLDSRztM5iWp1tYLzUYYdvnNplzNQ1tboo5X
4D2ZLydlOoqAU5yrEpKvGy9vTC2HCOoKg0e3ITXUPioqJcJOk69IyyVwnDD0H+z+zLp3IyMjUzeE
Lu0q7WcuWN+x6liReazYf+taTjgEXu8XacMkC1cfosRaR+7794pQZI+Tl3W/zCYNZ/pkVo/oIKUZ
YD5c7EgcJbtQSFU9n5iAqucASvgVpa7JfUc1o0NpyOVkCvnkoemITcJ/Q4FDPJGFijxhUHL+OwkR
1CSac3x7GPUNrMEnDsOZHt2Pu8ta4HATOHdH58KttI8Y7D4tlg5IVRXrj7Jk8MryBwRjXSg/jPxi
j7vY/N30QGq9Z1N6eWWZv+SeBMJQhGxAoVw13CWYwE8qVZpAQT/NTnYBsb5BoHjzSkePJKqBm80k
bJFMz01DNHjtZL5XXiArgoSloEKzXrNimCtX/vac7cHTZ3Oc7U3YfC06WWgPygk7BiGJmTgp+MU4
vICXt7iH23b/9PWYenDmCDCkJjt7GJRuxgcUEAVXimmpCgWIr06MIkntKRu5l3YX1Ji0/lAPctta
AHyFXoDc28GVJqg7aYZZ9NCXw8HAGGmbVObvafl0P23IkXBRVxMWHXOK5571ZJklwso03VjZLJz4
VXDMZajI5Jyob0lFXv7XeoXhxmlJyS1XIv8hk2XfYB1FKJYVHV0QRsX9g+EjXlK1R6OSMx28eM0t
Oggao2vZ/uAZ9rcXvGf5fNROLDYecbUyNXhV2c5uD0c5tLReLvhlOaCY3RsYtL3tOZFb4InICP36
415uCdRMv2nSEL5xHzdEJDsmzovO1FUNJv4g719KY0oNy4HjiOjdPLoopxg1wmBtYCpkI92apUZG
ctQFCTsZW5sd7pSA2BGV3+hhVc4jKjqM37iE1xNxakhvE8aXG/T5H0OVQeivP9p6lkRNtC5HyZZY
4uaiGmWJNoz3ICi1+Zin32imsaEtzUInuWcQGbbOY5AoZGFBGB0ZWEBTIq/wjeu8FWDJGfVwl2Dc
mYh+/T/VaDtoYTASXvYWl7DZI9ENsDWpMWqDvKbjbkoqjXVX4FEe0TX1ONVynFfFXNbeUVtK/8zg
FJO01gU6XaU0QxJ7I7EPzYM8+CUTvRM3Px+inn4GmBqayYczndbeNul9M+o7m2mXxPN+Y+mmIUVH
4N5xSX/2qXWozace7LMHnCe9Im0JBPoJxxgBQIpaL1lEZHHpZNYYSsEw7fuIXAYTU6YKkyL6pCKR
CxmAd73AUkMvzPPFkObsgfqBrRMb8ZGeNig16glr3uNrd7j3WpIxpGw0U86Sz+clGRgkAIDooAf8
Z3z/kJcYF5IjV080Lye6CdOKjhwmzi3zx05HL/qramOoT6ItfbmOPXx4c1XARxruzczIre5GBfEz
62gx187Fbhnz/0JQSkOgK8cTHuTCjQZFK5Bli5YlYWMEvNnpaMZrVypwhm8iegLeOstWL5PzHdYH
mRwF1Zut9hyMil8cSnU08gVXPRJtJhGqJGhyb7bwNTGq5xxGiYNI5mG+YC1JMGW/UsaE64S9hoxJ
bijLSR8EQiJ/yRbzs0svjruhhqqnmxsvfL6WdMRVdYnIuJ0P5tbDGerTtG/mUtQUFlaWd58eFHLH
qcbG6QyibAAnEfC47csowGlq+F5FwmArPhmfEs/McncydOgfbUsEg9DJ3tivkgvDo2jn3OiZggCd
jNKLgruMyxUn3zWbgyO+Iy+terXuOH0Vl3/AOs1YQQVWg/PU9RCjk0FgTSslQLeRLSaWpn0dwuNE
iGLvH+KRA/amyR2k6hG3e41EVEFCbhKY95BKEM8BPPdxQPE6tmAMZERGakqxi52fEvXqxuIYARpa
lGFnzj+Fxd7CsVLnUKjOU3neHHUNSntiGtyf1qFbqYENkeynzGQ2eMIL48eBTYviVZWXiWLG8wGK
A0+Fg3gw5sZ9g/VtfU9/noxv0bJLJlTSx77tj3FhqFvfht7WL4/AhCUURDfUPxBm2Ta5VUR5eWuB
RJOJLhUh0Y1yGJY2JK3p8B1VRUuCIaeIc/t7C/vTIoRdGSDjZxU6lrNrWd0c+Ltij+23pe0S//UU
0HhCczBxMt6mnjx+9cfqWe30+awyHtyOMS6wImI/8z7StHCcRqiGO+nFnTRj72BYnCZeEag0/AjD
YXI4u2wXPZYsd/y1olLY7ATacFlOjIzywq5pk3h5CaieN0MfovKPJlFTIBKdBcnIXc+JMD+aiuH8
t58vCZuA5yQ858WZlIGqdwxqX43cGKZwPQe52J/8xgZeLRDcqD7urhWJyOMmF+7eAuHF9bkMQlal
j7uOkY1tf/EwunrnYw4w/T5XGNy4hoVitWT8nJprN22Aj7XZKwrvLobMFQF6Rgn7IZMOdcyjJDhN
BYU9HGPNj5XJlygN4erLNAqquqLxWgYUViJtONt35niaCTwJm2iCz/G6L7OVRoahjgFs8fMku6++
jUvGqW43WWuCVXZngIgTTckzWeofGcbxBTRXXhIsyVPaMEz++VZ/pbYkMO10HgzHzoYs8GaxJOS/
8t2Jf6tj7EcXgqDRdQ24XF/oMxyKncd9WApP6+uZG/bVAt7hjoqlZl4vLyeWtXsWbvQrrNUL96KI
FAasF2U2Sr9mNDDhfMNMfvQuL7T7vsjOox12a8A2KkFZsiTJiq8q0pDMlJOVKNPzDZ6X10tsauTH
9jJMR1E4wFHP7/CR0FWIZkiIzsl7XLN660UEIZp2JNUZI0GXTfoEX+XOTSZCDQa9i4rKyFvOhX4T
T/FQnhpM4FzMI04vT/G5k1aiTEOliLnp6H0Y2ik9RnKL/it9KK8O7BET39FHvvUcQcO1TeKJ9jVb
AxsLOxxB9ujT4p2gTwqMDws4IbNmbbuxceUybW29RZk2dA9YAZe9j5nSvVnMVlfpELSO8gFnt1w8
7cRU2s2vE6bSlImdGBEwLR7xjq194DVA1RtQTo1gSZ0czLFKZ0YZutmD1EUmfXr5A3yetizj4mSV
MftIwUoDVpkzeJrqL6s3sMEZwO9YLJYvYZhCCSlbDgFBCGHnN5n53HrjnJKuEUWiJF5K1OYkiFuf
eBxPrMtSjvuPhbvPPktYXORu9RKmGk0mBRucMR+ZbNHn6UrLj6V1r6gtWeAI2LVJPdqwbwS0SeJe
gHbwHqpnGBLsZI1vj+r7LfX/p9GXfcGDvTbrAmF5W/HHDzr1DLmC6MRsP/ZRS4S2YUUcKj0nWLRP
cSlpb8fDWeUwSJ8gv3oCQKzSIOVKfibLWHpol27Xk7PdwpOultHWex/6suBcpmSWy3z3dONxLRYI
JS7MuULFqPKJzh3qHY8pDpWc3TZPO7sVwz0enNiWJrgojgH9x5+liAs4BnLwnwHkqjAECJskQSPo
MygdYl/Ip23/6pfrS4AICnhnMPps+lQFy25YwZ0ITXX9BzErUY9AZr+OkAUa9PnM4a50QxJf4Yzm
qKOQsWj83lZfwPKlPvqtmanjqxlaPQMP3ymdW+bry1grNWOJkNAg/asMnn4IllNS9XWD6l04tbAJ
DK+rmAMdxt1QmS8vcplktrVgq/ocx4QVx8qiNb1ZPyqqQLYkhG+90NIi9fzBoNnC/ydA126UGpaz
q6ukcnCpWtpb78uwbVfLomytSK+ZP1GPXgND5QQrT32YNvbejDOfiO8/euyfVU3ugAOSJSrAEhF4
09uS8qIVKlPjOs/MT9+fkktFKafF3Qx0L4qvnXFA0oC3bH470/qAtlL+r/UPPcRmQPnpXhOENdll
y3cO+qa1YwIq+DsLyH52ljG31VumNLIaDXa7LAr3c9LUt/3SdoGQseVpkk84Vntg3+FZsSjGDVEq
1QEzXeMkCXpDTSt54ZFIo8Y0qv94xGAIFWBSZ922twqBIVQsGN2iTpmtY9S83TtGnXYpvQ9ErKop
zyOdTtmghdDDRZKPgYZIS2OLlKHWYnj+uakC3M14w4r9C0mnlyUQu40l6SrP2zVYGn50NFuLdOrH
QmfZ8Kw/HNGskCRnhJzgGXgz6d6j/Nb3dZ0HNGkEey1OV/QjPXNdupZETKvHmEYjSQyFvqcZy66Y
6KfUHbdpsQMPQN+kJhDiO8qiYwhPQ4dHbLGSvh7oNT9k4YNUUIZdy16mhGiRHP7JDB74DQUwFrGv
aZBYc/tsiGUe8P8aG8OD4uakjiCPoXW9HwTfZl780lSGJwAPaqXogZRSzv4xiYXXuORrTwBLI8+a
tN4bLqiffRwSMWqpstz65Gl4xkxXQif4DzRNeAuRg6nZjRoESs9hmIOHss+0fU43Aucy0LeUGz06
RgN/B+tKCzThWl/RBCvm9ARfb35DttkyDtce+or61wLtyJdLHKJqYHc1eOye+qXsGZVNxkdR60dq
4gwx61dvFHUwVXGp/bOj6MfiX5azfwndoZh147ty4kRPPXavcbNTR1ARhXh7Pp+FeZVcJXWFoO+6
DawPgRLM4fTFLfRLT/9WHM1VZZolWPiY6BUj/FIcshZqQ1OecmZeAJfCZD8i6g/s84sdSKQOJefB
CakrmosfJHDdOTQb4arouy5MvlIB+5q+8Rt0Fg9NvohxphjujfmO7NRZlWGItT6SfQgTU5lY/mb6
gQ5f19FvKCcroVZM9wDo9v65T77V3YzNVnrp8g/UsdrA1nQBFWQ4gblL2dj8WZAPGz5i9BpjaYQd
UisZQ+yhYxNTZuxoddFPimYu8X9L5A3wgkaWY62759+HmXfSjcrg0UyTIuTB2AOl0kSkMYHxDGNp
3nqhikYslgui2tMZJkwhf62T2BTya5dtBeoo65rnN6am/mLcpWVvJiv4O/kdL1oIgix3mi5Sf92C
2JxO2ayLfwRPEAamSVnpo1YbXV/nLmFft8C5ZgyJPii007MktVGMvNNalxabY9PKGF6BmYge6mFX
vdsnXM5UL1t3Fa6vpU6v/Kei6ZS6cWl41bFzMpbsbBieo0HQbAl/oGQKIKlNsJ1pOYsQdIoMVhe1
iXpKEbo2tnE7XjM7SO504fv8v1kFjmbMRaMdF7GPpzG5nCcq53N2lMD4Lkh8raqrAblOOyW8bwmg
wIiev7w6MMwb7q8gOeL4Es+ibnOs5sF59G55Dd202yGsqwZAPH3liUVKZLYNacFmbNiEIjGGt8vs
4dt7fIYWLJ/eLVQFU6to+q14IbhYFPM3eBt17/hu3FRj5WL8ISSgbdZ63ex1yrOoHpOcVaqMD34m
enXNbuP+kOP3pbN39JiovcAX8b85fMnVNCXwt6DhwmHJATdwR79W0FR38ObIJeDOOx4pXCqkZWTV
gbFScgrrYwBsUiD7Gnnj6eIA5gqWMUkvKDROUkJuCup6mZ61NkENG1uqRKQahgJpIiYaDu0kolPw
Xyu/K+f9+KALyoSkPFHNhHYYUsPT46vMxu6+3XbMYc1s2sBDEJlm42Jjdfn0jzsaNd6elV8vhiAO
mt0EhD+sfUNuzgfH9ObzeSKjZD93nTEMcW6/cainyC5JZLZ+jwXjBtt03p+O2FtzeEJS0Yx0jeYT
OGZo/ZXVbcrqkC9Yv2DislH2F74H0ujPIuMvjrI/NL6bTpNCdNm4p6WYTRiBDz5dS/U5+Z9E5omw
XBb4CFoa5iFssYq8Kc0JOjLL5rgd97vxPoIzzkAvhPHUUuhc0/ZDyal5DjotXvqE3BjPX+gnkgD/
FiGbpObmbFC5B9Y/guDBGlSJz3c0Ejn1DBbADb559HU148YBTQikf8+botqwyFhPp295OKDBaZP0
mczi6wJrHx6RlcQxPcJOh32cXQW8Pm358aVeVYFanoxrLIizfFeUIeKAEypRELmG9p3/2HdUTnhE
Sh7ykB1qV0lTfOSWUhDnMsyyYZ0PlVLB/khiDUCl4Eh/3UAeBDNm6P1hxg/DKol17i8SkyLqW91z
0EbBh9PS1YFBNmc5ayDJtA1ff7/52sPaq/OnXK2+DBK6R4FyAZY2YSHMQaL7pwRT+0FN0Khu+wai
cwNwZ9/KFsBLH6RMzNzco5jC1Bc9ArTPh4JHBbfpOqUhLeqI5UG0zNttphmKpk1M57u3kzsvQ4df
NgtxGhgzInQ5/SOGgg8XCZJagkTxQV8t2kQLIg7k4RqQDXFjIADCtvsmuIbM1n10lR9ssF41pM76
MRME0ATBu8O9BmPc+SU6RnmV5tOeTraWojKkdj3b7wXqq0TPW4DaMm42eOJ1jmzuWeiIyldPaELj
vUCrUmCfoq8N0FeR9n8zVY/PEdOMIvynzVJ6+DFV7fvtcO3RXRboD3zKrxow11OvOCvPvptyfYy0
3u8BEBPWuvdyj0ZVpzE/jEQS5jtZwurSRlH3R46Q+tn80fr2p/EnNCAwdDRoV+J9qMOqfjZ4ELtG
e1DAQqTocqRulWUUTVviGV4NffB5xse9QZxiiebaJDuUb5prEeSEIK99XWmyuFpRrUUuhMD5QvMM
1P79QbF3ojurOs+BeJGtK//Q3ZcagBfkncqBxVfJujrf1s8ZxqYyo8Zp4TXKH6Lp2+rHwJr1jq0b
AIS2g0zPqQwMJ0m5WTyEi4muN8ByZSiDVZAFOSV7G1XX66Rhceu2LfohgqUQbBZUQj8bv7t/n/5T
Lm697TbhBtJhRY6hFL0StK6gZrviPb8NoAyW6+54dxaBthAxLdJ6Je5fIQxKG8IPBsVoo8xpJpyW
OxYHx/l+0ZCCyjuYwEF84p/zHiqwQhqpvM5Y/dpqrUz0QuoVrGylh2UxUCGWtwrFfYP+WSp7E/X5
zubADUXGiu+xqdJ5MtP2TaD7y5QkmxnIBZFasrp3pRHF3BpiKA4OHdxcMmvQPSKThP2lcVP2RLT8
eQAQxHA3nGo93m6Aq7b3K1GCtyBVtYNBe3o0aGsnzcaIQc+5T80HRr+NXMpvfSmLmy7eAmIQapMD
VfRzyPCOjr9HzwEixVNjLpP4sk27rnWM8UTXHTdWVvohqFPBnjmRD5n8NFt96T3hHb9HCkG3oHUc
Efw1KZGTgUbu1ZmOJrLY++lRY7VcCu26pXixCh9vF+mFnJUYie/nlQ3/Du/yi/2HL+ZIiWuoQ04j
Vrf8DrYy03jRLmqd9QWkXYreF7HA47yQ30uTcyOVRlAMEKziJ25S3V9vHBZwx0lCeQbcYwhmU3Zg
AbE7/VfNMGLHPJIw6EP2/QXrcUysSLXO4oLmrMXL1hlRduPFZv7uUja6+lMz4Xj/If+P+ULqpv9A
OkrJJp439BOOOAHSqsRH7o4IIiwmrFHEy9P/bS+Ws7JLyBgzDEvNwrybPaEHSyeMJ28U/NahKhLI
9y4zML19VAt+sMqRdeKDEoLyLGoKtuo9XCuO3Gy7OMBXHT7BtBVJVVjlAhPBSPCAe+Lc1jre2q6J
igRHpLhFVt0oezOroQij0pL2scVqQnZeYf0MtbA9OgA894kXO/LyMoEcAQ0uEIolDylvVGEVH8OP
GXs8MjCwOqMDyfYuugPneBOxevCqYPCL6i5cYtOdPzHrpYu15sVtRePYd+FYBfK5GHi6huO1XhU3
FyGdGXSNrsUAo/ctH2eIAIc3TksuV1MU/2Rdpw378iTcovmEDOlMEMf+mgUTxwMoNO978M7diYYA
Kdq+fiGw8CNiMzdz2qvmugovSSQd8TRou4EnbMu64OwEHyKcqMA8XkJizZ6smr6qgFLX+ydmcMYc
IOmSAEwKBJHMPmSeMSHhyfxnhKxdv8z82ybqRZM4NUn97DnJmEJ+3A2INZOwE+iYVT5+edBFIwyq
pQ4mbTwOHbxuQtTUScU6+JEHtFVlHpKS2mAj7NoJIFCGvi9q1cllRONuJp4+gvq9o0qGfNg4S8H+
8Aspc6o9PGzkB9P4UdHZPMeGywRjNVlbZ/LFpG563zcihZ0AfGRvnkD9VO5hHGfKEMxciy7uR5CP
lu0/OlykPnsglftZ+d5oFZIPkRedPc97C/Js8phVTaDIbNjSDX2uUyXClgLMPMRV0r8VXlJl3aDf
h7ync3fxGZM8aJccRoFi7x4DokrbUhel1ZNBsScELqSa+DLOU5xlvJe0J4rkKb41xLBhpRqSBsLw
s/x+PCs3vk2QahaNr3NDEekF8zF+OtijKNn6chJVycKaCm+MxRG8a8ouyihoFcb8BAzWfT0qXWDw
XtDDF+nYR36M2fBnkQR9XDrK7860OYMUFnfhpvAAO6vneHk4X8CLDcRjKW/jS7GRUmrp6G/QPrP2
RHgB8WZnIiySMb2GiB0lihVAyxDaFhzkL95EOeOK7TMgO/PgbGsQFGbEco7pOpxUPbjiyKajYMmN
527iXT+liME8iFjaj01ZadZguauGH3lHxEuy+JosUumqNv+aWFNS9/1XKh0vNZH7GuM2FFLhHnnP
5g1WI4KbxyRmkv9214mDBRA9IQyY60HDKUUxwUFo+0qV6tXt4Ei3o5EUMOAWznzeIfKKJokr0QEj
ZOujf5MMEfPz8jRajDrhxFZtqtbp6Tg9V6m2pPhj9O5vJk7Mf2wH5mX1kea+RmLYrMrHN5tlMBj3
7K2ovbNB6wq3gZghI/mprrUlVRrDoOsuJaM1CjqHWhQngL8CptQueJQM8vD4jSnmSI5+AwFhq7m8
1h97BIiu3PJsXt//uSEWaUaTYq7IOXRaE2W4j5lM4Zpe7sSvnAu2qtgW464OO09LOIN2OeSdVinm
Ob3uIwBjEdLEI4LqI1TuEcsqhFlVAYnVd659T1+M7hWWQjP5drohe9ue2B8TjH1kJ0ZawBiphUOr
zMMQtmzcrGOGWrrt6J98GxAstr12bAinMagN3DWg48I+DEt7/NBEGn3qkl70GndWG3cJQfwiJMx/
EuhwgkYT9EGv5rSoM1RPL00+xeEsdrdXfDMcEEbHp8BZ94OEHrmq0IyD78e1H8KVEOO4youI0Uv2
h4DlDgBXuEyiXrw4zzn5K8JkfLq9NoTQNS5Pqg9QbSifQb/t2WqabeULswenTGWZv3tHkuB2W4yS
UHjenE6QYmfV654OxhDu+Bhc7YernNA2FC8S1vvWHY05Kh7gKMDPxMwMcojqA967dZYXaK/SqP8y
I1LIgJnnj1LbjmTMOi+7VjyM4Kipq8ypM1BORpF23DN6UVShx1PAYpIyOgYSu8k8o8EvDKfREsCi
TFr2J2dr8+/BsTEPmqpszONqDfJQNcAJiiONoLciUjOKpOXhT9BlCiY1LG1+AU8y6KVvtGZCbIge
50qn+j4cnnvkTg7OCAffWU5nKdivj9te4MfhzLhEEDVh5jVcG1DNZ6kx88lD98SqGcUbzOYy5cNc
RwGuWLGkkQjwYkd3v6v63INlNO20zxyPus2mnm8LVJzbLnyk4gGxQdEBnR5MNbZWACBf/xdsUh1R
nKcIeduvLbjAeKRInLwlD7tqNscTIGgfamaMLV+ih6FHPsJ1Ike6KKCcZSCnncnjKE1EuPDc5YeQ
TXJzmHnutTvPXiTmEqQzoROrLC7WxCmFVu/5F4WzmLwDr0xR7SmEkQC8Slgy3XRmAEc+nzqK1okD
tl3bKyV9ImdN0DPIQevSv6KMP/ews7NDD4Ys4fnvRWvJwXsXJB8RqbNBdPKTr6MnZB4FJvBA0vHY
4F17o4QFCaZ9UhXDMEWMpyDdZtDygBNl8xq+B1LnzomchFQB0YV87+ja8IBk2AslTvBKrDnMiHM/
WOj5sKXnlKUMvXkDFqodvt/uhqE80e4cAMHHtUDCiy7bgxrI5/O313v935eUPs8LceLLF5ppdbXM
CzJCfuJggZ/0SzLhG3FaiJAc7KokMiwAQLhQrUdsvNSG1UqzxihDgQrOrZwcv+Smis27l2c15o6k
C1dNejMPoGWwb5SRwpzoL10+hJJ7zwpMhYJKSLTgISPjhVQkvQiDXk+JXW9LRygwvBC8oXuV8diQ
dCPZRvLPxtG3BxVNuWhKDtqGHntN0qPe+KnlwQaJ/zNt3K+3W3dWqGBaAXPKyxwwtbJ70cmj90hR
Unr8BNw/Y+FbJo1xjtItNAdM7qfe1QVbCiSyQHfvs9HQdCQ3PHObd+2SZiyaYDR08CoRSFqbvCxV
cJrRPZnmfyhDcmLAVHX3OFRTxJkEAelk3njhs6BpGKfuXh2KGjlMLlOkVgJX0Ug9x8tWANqMtTfu
zqRwvK4i/Lq664fxXRUDVgZKIvT7Nj75GlNlq+3w4f/BIwZSBx4q4QAfpkxebf4yH+mXJmQYJ9sf
K9P03jo8+Gh9y7Y7mk5f19nQaEDaZMzR6CnKBjh+3Qg3IWWnn62jCEO5zSvtCNKwM8GzDNBObzIc
X7DMC5UNNARB+gDuHQRgNnY0ptXIzVeFvxGs51NHaeQUj+WHlq2EbV2qaD1k+Bu3XH7wHsP/Lemr
tQ3iAWdr9Y4AArETVDdf3McTlIS5gdMImSZJmcr1Von5JaJnTKoKmwcH+7zu20UEuSe8233qnVgh
yS3/5Zs1OTPyjs/l2jcg8aNQ1CDw30s7wJ8zeedU/nB9UD1aiuFNKW6sFFOTSbl7ywkctC0rB3Dl
ljRClxckjMDGfQNNTSnaSO2bfU0paZgrNuZTIrDK9Qna0m4pFcDNV2Id+cO4RToCHG19MjX4pWIm
E5dBT5saZu8URsXsQjHYrAdzwHJaCCg1s6ORPE6Y9MqXo5/XArtvJxbJuP7jPiOcc0nKqTSpHu50
IR+nQiuADQqYENKtqHHZxDgquCe1xEQktlUmpTT4kzoml36HPP7QGpxP+hHJ0eSHwH/61tmRBMbz
QvVc73I0FMKZ8O6AdF33nD60Qw9VTgugWYm2UhA9f6mMgNqCaavYzVunOMA67kM3vmLwATVCw8Z7
cYv0scyyjLr442QdbSNgT4Ajh4GNgHPtDyfgF2QExRiHT+ZyYirj4OT9v7YvoYtRB9BhGpbZwqiC
N1X8LuOeIN7b4k9YEEH0oawXY0efDsxrNjk7fJdCHlq+CpwE1QNNdqAinOmTfWHo7C4bNAg1p4so
B9NGAWIPaRwV36bbtGJJsvR9C0LF4Ix4vYWITlDXIdZ5WBGtn+ZG4NrR2TWj/H9XpHUDfVifbVo/
rxrCOtMN/ddLixJa9fYB0OYw13KqF6Pttpllufh7AWLPUljGfwbLrZkAWp/phaBTFEd2ZH4hD0/x
hedy8FpzmccbHdekoap2zOsIivsIbYUbgY9mWUR5O6KzqS2w0uVeH1RQ9z6wkf+mJ2fuvug6ISRM
Y6O9W7vSYsD7JyfxZgeLi4KPFLKWPei0PpUJjsLqS5D8FBWpR4kywdDtzq+CgQ9Cv/MO7ocgbz1L
/+tu4/IGQ2NPsTmNF+3hY3Anfh1lnM/VtgpkSOrVHNkQHtJpcBv6ayd/XBjerg96D6etm2xNJesD
RzvThT4ENANQGCgqYrO3Bk9Lh4ObcHcndQ5dc6rPCk28f0tEffXCFxZ0+iCV/FjN8KF0Rx4+HcEc
DAWXLxFS0KwmNC3VSpTVt/2OnpJXLB8i02pq913ka/sx4Ph/Tam/5bXjDFYYRCjHVNUeFNupndue
mkJQGPWL/yOn81MOadeOeZcZknLB9RVnAcKkNLguW687WbBdQPzkVcd3u1Twzy8yqNFKxBLfDh8n
7N/J5zMh0tjFsoS4nfEiWLIwc2IWBhGREzJJaco/VFeDhZHuTgJ6j6A04904D2QpcbtUfYL1DJfz
bapzrhUPz5tfp0w875sB0umfQe3DCrEJpOA4cT7twvlkbmRp99DQesUTMtEjnnYJFuZMUugyGeJY
E+wL2qYiJ1R19AHWPUDgHCeLs7kIO+HHojHX4gfiGeFyU6lWEisJCs5m4DOXSgn6yopaYB/+k0Me
jY0eRt4v2orioRB3JibP3gX3bI6eyIdVdiNeritLDB1muCFIMrnQgxVpZkYOE3MWmD5FoTLFl6Ep
Hyx/ftoS9k2mmsAYLNWh2CtuT/X83zBGbh4x+DZ2LxZm6YEiszKDS5vHmj3DWgI0zCHtjPTU/jOK
TIFc0qKFNnOpVo9XxlQw1dIIzB3rWgeqa0UE7+SF0NBd8HMng1BgvyN8VjKJT2BDr3uN4kPZH/TH
o8cejETGAnsKJzKFVXfS+YT/0sLwVOt4dFx9BGmws3SXaY8UY8fWmr36PYsyN2kCne9ey9AbB/y6
30ADBsn5AQ59Vs0t3TkMviOUVgiM7Hr1LrExY5K59qdnIEXZVys0dXDCYr0bY1VsS9KmnSKwqph9
7ka4yyJ4i0CV3j0YvCOCcQuOD68Cc30yjv+K+FcxwxRF1aWJJb5CMgw2kpKAgNwb8HIRT8P6KxZP
iLi0lqLk2gKRiu/kRoweZD/d65Us7+cLXKoUgzPs8rarN7qHZ1Z/0d6U26WFzPBd8X+ZcxrlCUCk
VLXdQgLonVXMoox6LuD6O6n6dpJp8dq5w52fir3tNHmFYHJzfhoyEIjL9cvmUmgTRZVlgKOqQh5s
19ffcWBDPKu/XE5JYOmJUn3vlS+K1A4XlHde6vFxBl2L9EhU4Tv808yAqRWZhbp2JZ1S3Jio57xF
JhRUfLD9TmkwTrc2Rc0OICJcktnKg6b5yTZeunSbDNrvOLMigtB2AT719+dsqUtK0U4lGw8WvQpF
Jx/peRLndXhi/A9idJ7LfybJKle8ylLd1IDDV3Y8Xd1ogBJoABIj+wkQ8Usit0ZkLgEId4VDrssv
0QnNR9KkkC9wJJCrC+pnWaeP+/MPhod9BFCWzSVC9XGQV/OpsWHT3C6wzAAlJi1yqEznADwNHWK3
jseL34umyqPBY3FNzcIlPQcoqqCp3faI0R8Su8Elg5BRXQVD7+5REjDxpbX2akmXMoUhUDuzRy9P
K26h5MBTm/JtxuoR2NU09ci9mBrhUO0qTc/dV65zJf1qko2qEqgqEFsGhOCACf4sMvBs8NHXLFOV
V3eS7wKNfTayX5pCsbiXDY/ZcY+QUIK0AUCM8V3dXA0uckPIs9KBVo5l0PoxvMYww5KDTxignR6F
57ZtitkhSNHwPuNmV1NOJ1BpPu4nU9sPzUOkgpF6+hfLp4EfGnxV6meSTAMUFY++84pfq+mviEZJ
rTEn9yWNrmtXik3R6I0sfXl2R1vIUeKqKwqvX034tn+IfDSfDF5nLhM18qccmTRG9I85A9xZnrRa
nHaH8AMoCkTuAXw10scI74s8/G/+PEXi5t+zvOyUx3+Ar0b61CsrGT+uQv+emkZfgTq4uy409Hto
RmYfGPu/KAV34uR6UL0NJh0bzs/s2oCatTtdy/Blx0yONl8tzj5V/lpJJOz5qNN+iVvjEH0Wm/GI
UnHHZVB03TQxGwHgU3XfUAi6rSeicuUjCh8CsXu0FEPo+NH6PHtORWNIRtBCOfnb22vW4HdCWs/v
1MGYEGyQ6FB6K1BiAeaFmysNmv7p+e29E5I9KWaQXBhyZSVfHcQ+nfy1GXQCKu4VffYsRHr8DFKP
IAmfBFaHoxRfVC0aRTaPNg83p9+2oKG7hklOSCV+18jTFDvU7M3PZ7NPWHhvy+6H02A03I3+57Mc
qdl6SbzsP3yPFujUmmtiULU91D6foJL0gkQYVXjsv92TmZ2WeuVpnHQXG26LIAvkfcFdL2RhJoIM
zh1m5yPrD6+VQBz5d77ptU8KpNDbQiRNdFeXLCrHax9603DTABEO9BN5JggnAc5pkb5wS049+DVV
oNSBxeHhyopUulKGRniCULsHO+CkNgo1NtLnP1io1RJ0Ts5mdyeuUVvdDWCOruUM9MI04wa4Q1wQ
2li5lCU/IeoWmZZB5l+mgpulxUy6pffX5UviY33ctcXs46jptkJnO2xhMCMKqvOTdt9jfF/wzGIy
dGVkfXh+Euvkh0J+g5juZLAgRQIK/uI2nqh43U+O+tfWoEZDGnmFenEXEaDui2oLkWVLo0rYDLw5
46gkOVTam20fyNW94DYUjk7Xy2g6FCgrVoWKp86UQpmttPzv+cZPiAyOSxh2KV17JWWwXUC8y04k
9lRdt+4TRN0XaNw/dJ79pYdDcsFPLrGfJZYsQq8hhGKsjv2AWPtFfyatUAMDDrzPxV8B+QW05+O4
imw/YK3MpMfUmXg4nN66xZUmEWM+HIA6grb6i24vqBYmoP48s7wgyIhHtSK/6F2OCGDp+n9iDloH
5XDycA7432xKQrecvLDlb9nZuUf9YHFq79zpstI19+HNe5ffDLGQUJS19uMGXOPuhl4TEtHRgtvn
BT640qgwq6Tx0gK/fYveMJg7bmA8lCd8HAK22KTvlWLLXBwmPEm4keDz04NTJTmAf1vnMnUquKzW
Q5Zo9m/IFPtUYzJUfwcEQNfY8MVFeyYufvEeHfB+HTy4QJFaMlAZQ+H1cX9bARjYWaUZxEj7mt5n
e42nYE2YG0E1yxLGVK7SZPLU08khkT5ob7T/0e4kYv7HojLuLHQh3+e0KQRNOCAsctZX7LzTdkEQ
V/Z9ppKzGa8RjDIyWDveztf+j/8peIXENcAbpZBJjKsyq75lHpO8y7iUiSCryk5Q8mzTmCC0YvsD
G5OZmRhtQ1xBjKVQR/4fSd37qP+nXHRJEi6P+OhnxG5Tx47D62nUmOzEhqBljQFuDvVpRt8Etm1i
rh+wH+gJtbbQsH7BjJBAju9ynLZXDOqPBPXroGNAKF5yQZUvLuOBdU3boDC7WHIL+x1KDvbbWTAb
YwackbuxCJkTgfBEQOZeQAiCbr7QVbQVyxwsdds09vuBIR0/BDXOnsoEUQdDcPszAJrKT/TQFV9U
E1Icozk1Hz3liD5zsilEPnb/mxhtrKfYIx2D1K5Xg4flLKSBvTu2sV63pvOnC0n60Xj2kA4=
`pragma protect end_protected
