/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3296)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvlx4PpMs/gLV21ib0v1qxxgtigNuFKTPIft5aWUn41a0jnm8x1Aoc10XK
2XE1OYaGVxnYNVP7d6PNBL9C8md0Uxl8FXudYQPB3aD/x4steUwu7u3z+HEhA0ErrNMYNAQMAJgQ
t29r+xvhF7ns+be4NtmTqAvb4jTUNKzPCQweC4J2xJCcIP3+tDi4HN77K5g9C+FYjPAXmZbgwtYc
ABfXKA1oj46uK6YGSR4Qdx2qM+qPYi3DZMy7CAEuPvHiREi7TNcNukjO5M3MI6tlWIvqNUHjGuQV
7a2LvJLvUhYrQbiIusb88d3/qV10jqEkgS4A+Kbb5iyJn8ByCnplhe1objzr0FZKnnrRnCiycQuz
AxkwnHLbWWeSlwC6JAFf+q/sM1O/2H0CklLqKxA9xmYZmM1FggT66NNyzhy7xtNhUo7TrJiNzAb3
5HRiogj7nL2u72QYRSgNGU1GVkMgnc6EeVCylWnh/ZW1kPcQ9zsGnmrT7Jj9VtsreQc0ZnA0rtaV
kYu4sTD2J56KQB7r2Lo0QF/jGoc1ewHlGupC38fMFMrTyld8UPQbU3Skz4K2WXL982hqcuIRM5ZG
9LFBIWQBkPlLCmfayFaQXjgKrgZlZDj9G1oxxzlmgRA/Znoc51iZHPdmkLQosUvbuhne/d1P9jjy
/1gida5n4Zw+QibIDXXdvdud1mBgwVVBcuyM1pfMuRNNmhZJY1iITqHRTm4FJLU5lOnDoJznCGwQ
kweAdsEcbR2ALOzJaHC5ux/pIRwi4rGDQNsC/nupOHhK70a25lPh2REwIFcr2Gk33gAdrXduKqIC
i631szVl7TV5nF11Dxl8Mo8JVY7ttREuJ+cUcfjQAmZq9Z4fVW3B6UZVx5hgAzWoHudHWVZaWk04
ZuGQQAs1ATmNRLP3h8N5jmPaB9qdNgrE69qHQveJ5drSJYV1riBJP/Bnd3GUN7lmdvSPpkbJ3EiW
PZYA5Y3V573ot5JuDywTqCn+4DvhwrwwVxDF0F/oy7x0tJFk5DFk2LFfi9k8zZgfxE1PV/MhXuA1
6yue1UzhclC83cZRRRlxxGMoPMDRfCMIzMOsSIjYLQiqooCUukqZHjgdJt2Yp27qfySUby7qUFzi
aK+QozOZsROda595eLEE3X1tHCtdEdqpyaqNmkpB3u+zgjA2m07189sT7q+/F53X8sZ2oUZs8+LJ
2X5uEvr5oIywx+PKki3SZyrXekJoiteZGPF5zzokH+F1Yf/HVF2MtZaBnrso0MDgVShiofn+ITYH
DF1i6NCAfL9kthuX/Ac1J2DRJfwUOqe5VXFH9Rr8vmYb6XrJN8/wszjvEFjwR9fnanrFqCNHT9Gu
s+VX/NhwnGrOrpeYUFH8y7cN9ndnhFzCpZ5lKhSN7Nkxqs9Ll2KYHK51QUAs+su0+ZAwe8phfDKZ
z2rUE+w6+KyScMA+5nv+xOVnKvtvbTD2uKZxhYn2NpDYvywAZ0m6/00iX/2zndOzoh718vAm0qiC
WOUmIbfK7G3Kd+5zyjWkNlVfyh3M6+oK6JusMfGFNfnPxO7Wtmnn3s10REeER2cIxcfJllI/euX+
SiHbWlkXvz/az195AkVpRPxU4TeF+J4F/MnXr0KdJfOrKJOE3Mg3rsR4SDVgOL9rzq5GLrbkfRxr
MkoFqIeaqkY/jXveD7AppaKm6LuF/lYvvqY8XuyH5eBELJxP2Z8DhPudZQ6eXMCcngCvhCduMxD3
FeHoInSKkfgEWT68LxsHYux0GBb2pWuqV+nL+TdrqUUSwE4bsURGkNspBhWaAeYTNZJ8B4GbfxK3
EXZDLfbP5HXlL7QleGQMRI5dL0N6aGxylwcsvXuafLhFvRlZpPL5aIZ5CQSo1M4Ctjl2WmMn8f3p
yMFKe5jFRpe/NZg0CjxFfGaNw1i8h2RUVk9EM2ux74uSVnC8jdPwci2cLaQgTshDMOeeJbh1B7ug
Y3uaaMuOHDglPuSR+rwPmyQNihZm3RAbw0qPsfvvU4JOf1mu5XWJ9SuAJAT/8ni8JJMY0vGcMq/4
wuJgjU4PZ6fj7aIHoCdJoym9MMTYCLBDD+0Wpz2uLMXeHsWFVJN6y5dsYzhnQF84S2rIG6CBVPYP
eM1WhIBgoqZ+z30O2uobOmHtdKMDpSeizeTjGX6APkElNtjMMizSL5NLtbjHzmGhVrweciePYAT2
uKu90cHme48SzapJtq1WwtBm4g5gDS+qf4KySEbjYQPiNE6Qg8tbE9m88z1pmAIZ7BtT4bITYMRs
1/aTXQN/nlZs6d/yPrFlCsCQIiWgAWgPLANsIOxDPperPEi9V6EbGBhOYSDMlKHQHIYSFeGTL210
y7Bbz/OmlQPsDy3FrvsbNh8t3Qgx+oX3jmMHN1s3dax5OzsfTYe2A9A8X1Ez+ysciNAn9YYK9EpZ
EMGBxIRms/qattK0kAU+/Tluv2jjTHsHi84xL74MIQLTAByxj9cBybB2LWgUk7QEid7GFYDHujUd
da9Q1LWA3qpjBsuzqdIrrYTnFGW39yRIRhet7mDHFYKAMQ9fGTkR5a/0j7RdqyDTP87f9spUbUSv
meb575DoTHvXYr2yVoIdAMyp7FFcBMy7p2pDR2MMt01x5fkkjyFXqMjBeOQQsRpSigNHyjC2h7sd
+gO7Q4aZwatHHC9sX0TB4an3DeEozi1Jv/wjTcZf6ywARYWa11M90eXIfbBZDfLRynTan3RfedUe
JMezQ6Elk9CR/mpQpmiJxJ95OEFaWG25jWAfII77dhry5Pz4vdkHJAl+GRBDSbev12O+e2TRmOXx
5r5Sd5s1spm6BjxzjHJMS6nwyKUifNAI+fi4Gymvxh9d8t028os3ZdULFjXRvDOGNUcff/Mynz6X
1zfnTXti3FM3WRN1W1cjNMKNrVJhtoqQAoXRE4G2Sk5nC1qN6kRf4v64/zhE7by7WtPwMnxhhud9
9Q2u5peolNgDFsJk5pvf+CxLtwWpHe5Qbz0BvhsBGUocraTeHnY8m5ijGiAqo218PMY+Frlrc1LV
5ZKTx5Mi26h17tgWdxGV6o1jMswn+3Vgch3whUp7zGO1KggVcVAnx5UR/qtM10gRGS9jKPsDpUXl
VGfqukSBqVsrUsGqLqoayRN2UbtnI+MWOq+7v2e86u22x7kvZz/YYXqo6oWk6nU1oUCgP6Dk2fRr
9evEPKC8renn4dCs0ydvmhYL3E1ZA7ydRhgdjebD1ozC0bRmb8/FGgwWRiwLGQl006DBFKE2R1vU
s3x3Drjt9fVXkYUKCiM96lvKPgr8Hzey7Z951lpYS3DQHElMwO5lsk1nSl/xX5FDrsUYYJybGMP2
rTDXGcJuorSSE04apMGO6J7tX082bpn1Wwy5hK8JQdMLQSFX/NeYXvWvpQJpmjjZDDXtjRq6pJxE
LgdarONAdHX/AfA85ea1XVMoDfjHo4n2xBFBM5i7WkQREO1Fbp9CGiu6oY4yVaSqpoqGW1DaigzY
sMuYFP1R8ZzibH+B7HhDkQd8uyYjRRfKjQnFxHAmHclAS7UbjJm9ccbkmv6eV6xcqTZyizLSl4hg
HAhKOM1GjlgMNk3RMaMBpHZ7eOS637pE2hPiQfKsW26aloXUhZGewQ+KwmH9+tOE5ufa8u7QR5WT
9strSrmFoeHk/PaBruBdKz9+7FA+kAvX2ghfumq5CrZApsy1av1SS+E/3cj0cHj4EdPj+Y4CU9MC
3INC9gyooIj7EWG2sxkw2lrdqebFpMuNRRYO7aKub8A3lLCfGgx37RNkyHdFDueRBewUmqTeeMey
Vu7Z7k85nSxq84vUNtiHsHwgxpQNpKK76kYn9gytK/0onhhtgiAtMUvCm0QKzqKt7TSeCELqKuzX
V3LzcqOxMWAI01bAmKU1nJpN9CPVZwoUReUNYrg9duxOpzWYtvVEJHIdQzUzVApeER3XyzOjbe4k
K+Gat9XVdW83GF9d8cu4uojfEZ9trBguuIvzx4+l73Aqcq61c5w+dXpDOP+k1XjmoBoLx9Zjoeq1
GgTiQveaGw3OzoHyuNly0gTdPkzjXtjVcz+Qv+TPxBTlv14B3fN1meJXT/6H1LLcG9ENNiQdwJZw
Q+cfQUbiopD8dGKhmBtVbLGywL01DOKsgeaoMRV/uFESzRFqYSLCgnp+jWwH0lyJ0q5VpSj7chNX
0S1jLok3g8dVZFIkN57ZLtUdpxdHSAccAMiX37NJx0rPYK21BIA6fj6zs6qXbDXpStYRXS3yvGcD
lpgrsnS5mBIEVN57OZKwR+OR2ouczvglFUqRSfosHk8rNfLlKFrJCPihnUHExwVws+p+iEXYYLiy
XGbtwINAmg3HsUVc9L6YFo/HzaSsml5TOhbl+i83RO+1kY84vZtVMwUVruHR9zs=
`pragma protect end_protected

// 
