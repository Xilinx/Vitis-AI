`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+GzawGdEcIuxfE2xohKZ4YfAgNY
udze0/JpwAsGtIi3JEG+f9Lc7KzDtVo+7e0axUtpWWG2zchF7YBRjZ26kg5u4E7NrejsKmQn4oFZ
2qTRJZGb5SJ+gdQBQzowrZ6DlCm5Ybvng4Y+fKORBe4O+BxCB8HAkjiHJvTxpq0VwrUrB2IS9/yv
BT0mW1nWT9cr5BxcHY80c1SIh2SWvSjyo6t8/Uu8goqodOeiB13w7hFPS0GPtfT7TgJBs7CKLsW8
/uckee4oJ4wGpwWVllo5zGtXYtybvAkQuljhLL1WVVO7DUOzC1K6BMV5MUhkawsVtSIUI1uopE0+
XdwuMcILcg+ooqdfyok1IJEco0IMvb6IaruZgQASyyLjD2hGN84yqszX4+Vy3hlHCOYrpAsafd03
CrxsjL/cJ3sllMpg25SVUfnKro1rWCtVcekrwX3pI9JuZxjm0BtVCfM+fLsDltG1tHUMvP0ZBUt+
+eKbTtAjO4hvQbsGbW1A2OmIiRqnDMgEbCBC3CRGwcaahfTlGG3yYVSffP3Oy3716LlsjUbttkym
TO/y3o122T3+ewWwdzcbnE8Mo6ycZG8vhVM+ETU2Tz9i8hCMMDXUQ6I9JX/ayLIpQ2HvHX0YCoeS
zn5eaDdSfmojCL+kV+lPW7SZjlG0Ev4gkpRmSJPheKjSa8QLZxJOEoDyK9TXJ3cpXf6Nj180lcZt
e8EW9dxUv/iaDjOSr3uzhXW7ZzRR0bNnoBuq3gMgVIfLdGv8Mqm9ZvJOTv6tTHKnHdy4jreWvYZV
SN67O4NPI91ApRZ9AvD/aDbF69xe3HahhH+fLgqn4e4xKe/srHErfk0xWH9MJIQqmfJ9+MEFN770
mHRebfLNNYUe47cCCrW189/ycaezOyGY8fJ2MiQ0JoEe6GlfuGnSJMtmIzMnu3VepcmHX1aYfHzO
XbRULxfEYKbT2fe2kYHpJSN5VBzg4hyENv9EC0iygH/bCaffE7xqPPrMSDabmR1xq8JhbhPT4Pn3
89FXqwiFv+7AhilKlgbJ1urwN92E6PtjyX1VgOevCbEVVJVr+9YJ6qzl7RoqE3xPZi9lNNCU0BJ7
X8iFIFjyqzrZG4vyaKRtf9r69aqK4bZ+kGR6S3+VT5Cqg0OA3f9djIrMrt+YsqYh7aGgfdzXfLDd
ifIMO2aLnTBgCUgMqYBW96D8hn5Mz/k7Gwkpyot15mS2MSF7rVBtkn8ejQO/shsq0eeypgc/PZbq
1TbYwYTyDdMrGHTXm2ePU/7+ltaW22upQZRWksmXtAcqb7JX7BspsfOJKE3JmM/XpTZBTAC+wHEH
cVngEi3FvaIXWg233AIOwPlPnMclWJB2fBEkacFdyUGoYgr2Tc+7kCDrdFNLAgurZ7JNcjSe/pvZ
YgfHFDECYahFOl1I5rFof9UppWXyLVpnHgFZByGBzdtEVQxyFEowx1L+u7rofWtuNqR9elw2X8sZ
5t5FteRtmUpJeZ+gwvzABWhlpT5WupJvhow8dCrquLKdptzW/f18W4i+oRJCYl8aluCEI9X7N/OG
cvwQz+Gc8O5SKLKQ03pH7kg9oKg6pZrlp2Ndk22ptK+Q32En8xsZ3QIbHk0Fi4LWgaWkMYn/NftB
4tjBjhZ26/l9RrF1yULhsplYmolrFNXynJMdbUgH7vWBmv+eUYp0z27b3xyTqCoT+JnlLxZfPjwP
0EpkzG2/RwwvwUxo/8dOjloxabdL8lF2Yx3wL2SWOwLoxbkYXtn8XDl9PUAJTkRK7DMYkszi0wZj
Dp3AqD+DEPx8LDvb+dqMpipRSUiZEpOViqYuAI0+k+bDhxYqnwba2prafkA8V8sooLz27hTT5kfB
aeI8GFCko7hQXO3CMyskes9q8lmbqu81rA+N7L0qTogZiwl9L300aq5S1GcX7FNrs/czoBSnMN1i
yymGWigWnECRiHmXpXLbRBmctX3itB5Dwzb+KQan6UZcYqzhe2i/IRwK6k7htBy7ky5Txoa0hsQZ
snTpWBYvzCe2MJn+iZ5pmLJkkRPqCtpk4Jja4ax3cNzwqheuZ0sV9sXcZ4KdXgoUrGP/y1GWSaLd
Rz7T6962dqlW1bTCcyum7CuqAi+AByLthclPOynJ5dsTGd7EYqD7Ck+3tKD+fTRbvoC9JwiLauYm
yuOmB6+SbytE/3KkM8MTh8WIYDrahA6qRyyO48PfnlD5EbeeMJTN7GnqTPOL7SRchGz4/AGZxAvR
7r2jU7IESoVZ4ejyJ60E403xsJZfbJC58OHbF+9DBWLfJegaWl6yAsmaPb/gmERI/aSp1OD4HY2B
vjpA6Go38hDAqRlNntclDTTqqwVHYH9MDGtuKucErBw5D/70MzyTbPjrWpJD6uETbxdTToBBUAJG
Th0aFdsWDgLq4958B4sXDzc+aiKpt2yrutnp/xrWHfScd/BJJ8bw6bA74PTc10ovwbz6X8SB00Fb
ovTqbXbAkYve7hH6S5ijRfenrWsMl2M9vHaooOy9pIDM383A2QJgsVqE730kXMZCFL1P99iUZo/L
A3sVBZnsZMXH6RoDuzIBzjNy3F5IDl9588zUGgQqICiVh9WZee9kjzcQt1iBzilhMAHm8FI4Iqcu
P0bsg21L/tUBHHL71Z9gb8B63BbLdQpxB4/TC44cNXg+1HboqmYZPuUVi34eRDN9mc0gZB2xOTfX
vNX4eyHexVLUkJoeS0rf23Okm6XHI4hPojKsk9Lm2JEt2X8/G02fOJxTNUwPPkDnyLTeRgb867ty
DJ9LuRvFCL4E97BGzL28L7HWcSW46xwpQf0wBuV/86n1ZsLnP/DIYlJUnZSzs2t07uNjuOVuKdcM
fE38sbmcOoeUj2GBAoSXE/1Toqd4NUAVRlyPBYvY3DPQSPpQ5MbkljXmej+UUttKBe/1nCwQD8qz
JGcxcKh8P/YKSEEQ6icw4j94EbPIYDCZJRWwVzK64UvHbc79i+FbUfQr9nO6u37SSE/FU3YNIS1O
oI5U+tWAoVVKJXADL7/HZ5pKEAYPkvZ3kppa8Pl51M3IL9QWeuSaOFdqUMDaDL8csa8kJnmfzLD/
AlVFPmO2QgGqBA3MP93WLNN4lOXmsyZ874vG9gMZF2QgxY/bDNLjmw1cof711OPjMyZz0hV+vdOP
AR43pi37/B9K+MuniSTocPjfJQ33HK0Bf1AEqbyGRTtpzCKt5OukQJGABmWGwPFzVrRnFQwWPIXR
j41zzIdrnHVAFTUelbPcrtYPeuxcYZPH8mOeyqbSLb+MBsjwtL5GUAsalmBMf7ifReqX52vA1nPe
pLP5ZqACMSGmQuf7u5ZG272/TIVNalbb22m2oeUCpwz3uflVsONpTCCLdUY3Wbin38NMfwejgo5A
GkH0W4dRAVUWet80IXN24z3aaseBb7xb/FPqav/9K0TdF1h6B0XdroIjDNoRZqc4HwVszjyMTlqx
LHSq8AdUMdN0ZDdD0JnDFfYu9E6SIoWJLS6IJ1EJRflIOTc3AKmG3mA/OecWwVf5jLozogPCHUj/
sBFSjXsCLUS5rK0VlG1YuCwRGz7kWUT13J7ubNSBdGHy+eHTN9ml84KpFoB0MGiLfECoYvRNk1ih
TXqv0vWWXmdAUrb96QsLDvD6Esrq7IR8eiMjkbvsOV8OyUmWnER9fblQLeXg+bk43OjRWR5PSO2Q
WpqMnG5Sk2x6exEpnQMPI/LfE4eVq2zhY4IMajM8FX2L/Ge/N0fs64KwKSdAHeee3hEMKT14CwnO
WEABLkqb2gtj19fMjr029xR05BCzeK9Fi9LUbYuf8dq2Nz1I5bhXV8gp/gFNzEVvZVerZwOkq0jW
akwyEzjphoNzaU1KfqTRrXN7RSUed7rVsQisx2qrsUa4SKDwQxf6dbsS4ekIRKRfW+jXXjMxo2FF
mCyh1pQDAZxEQS4qaeJeqsxmlLoM6L3oQgvXRs6u2sYWeHifMGj6NlTGjRoFcxLPmC6zDl+LjVlM
0mQjPJBLxZObzNI7i3CUlJ9EJK92Rpx2qbz4r8lipCivUNdxLUHBTW6IKXnHgyIeL47grgBNsngB
VhjXC8HPPnwoH7UYp5qVjNcVdIf3ScqOmL5ovcsIYb98qBOoow0XDPRuSSSDKGtINGnxzJtja60b
vhjpjkO5htwGDSr5swbL4qVUWCD/xVqKRhgm6roNcegQkEYnvfxpepAlLr20I1ib91XZ80LcXg8g
BwRwdOUrDuu3sTPVBbT4cLSEem7ZI3RuJyCJU6g8ZnrZgidiHkLe7Gur7fH+iGL1mmnlIi7mpINv
YUXK7pBRh6Ld7uDj47Be0Eb+URd+YP3JEBsXc8FpO08ibv1r/r89LLfnbbyUZuMyBDogmi+yBXzZ
3+tDRM3qqvm2s27YKyYGDIrSBjhQJTvXbJeFnbjkB75brCb8a9fJtYNLrD1quWCIQvbKAWe3K2OI
+yyogNCi1vPQL0N30+Ck/WVNBmj3NwAJ/mpMOBnuveB0qhdIqmYQDp8KI+12uGcsS01uDyXFYvcs
OgsvWm/0UQn/aui2qFyy63s4k/lhQqUrdVtULlp2wI17mEHD3yJJfeR8CrCG2cSVBn8FGpQzyH01
Crp+O6KWRgPIp5PT2WEtgcUkIYap2b8CVy5jB2QGzM+mjICGKFQGILO01LUgo8JsJAIMncal5Tik
agBIXPOnch7bhkQRMo8nlKtO1wuly21n/4ZcbPgaDw6ggqcEbpijOYiYBB7Sk5O6OMfWfc3nePfq
Y5DTjO5Yd4uCNv9xH8wCOHPI6Hah0mP1bC7Qc7xfSQ1xfZSU7ZMOcUp5gG6ubyriHirv+Ls6p6DI
ULEMGviWW7+SnZAS4nFTZRzea8nJPuOlfn/xzMjo7k6EZDoTJmayZKQmt9XOo/Cgfw9+8g9Pfu0z
Ul8iTg435OuyATSKF5VHWDqg17j1gDJwYaL1fZrnPyTMYfFnZmG0g7auCW07tP/PDuf/OxDeHr20
GbxWwbCrVQeo0/8JhHpPA7SYGMwXMhQi2h5sGrRUAI3d3//1/GawRLPAGfNiDPjJ4bKAto44GNJl
0T6gVk90x4J9223CGno1WFd7pslXE4M/qDI+X+46nouAOQroFM0DaK/RRsCdXIC7HhMxd2XcCj8d
FdTY33U2gdMT5ELYUJKyYI6iQbmk8SvhkHsk8HYrgswyCRFaQmdpD+e/LnQJ8D9JPTLL/CAHkn+Q
7ba7oEShjIcdKZiDxecgEhVLjD1NZ0HUXo38ZPni48pJ5++ZyHma5laSDBF+Efr7HTIqEBzYYthc
h5AglwZ42wJ8Bq+PknUnx5Al3vOvFRAB+WehyemvkWB+wTkNRnOWiitUtayR33ux9MSIdCaizPcY
b8hu+/4KKRTmuSvdGsLUyui69uL0dPm68BwO7YEonDF2QeCM6u0myn/eMRnjU0WCq/iMKyrarlaQ
wkNqVtGtxVcSlqCDBXd/P0xE+5s/ed+rpIeHJj1VPDiV/Z7DfQ/EweUVHxw0Zg0i33TJwGshcNIJ
CZDwRBB6RmV5OLz2tmdfwU3Ak0sL5SWXEqT3mRYSFPOTbfYzsvNtf2M0/4riRrVFDyV7QvTzvF3o
QU2YdBGpMMIfG9m+v8dt3Wj2JPsBL7T97oq3G0iVGB3CR7qyQQE28BVCVI98GJYUPcUE6WObKO7i
osc6P415c6NfCd+OKvaMh6KWEM2yyhoVQAPzQMCYrqURi0117r1W74f+AIO503a2R8IaMz17KV/6
ADrPxDqKkPxso2eSj0ceF5hg3tw7Ka+wSYMFmpIK1atneiGZb6JPGGalnDl8uVtUgItdDXOybhln
1Y9twc499aOEYtuZUtS0RrX3HSw/Nu55f9vGXOk6m6/sI8Z6zX+riCe+75oSSLMtgEMJwi6OA+0i
ElsAlK3kInsVN/8cofj5X/lGn1/t0bupBFAUXcLUSlb94pPg2IP6lPsCrR7EXbPhKaANCUhRu09m
NvoKRq5baPx0BORiuW8S5Ga+08kiCTpxxuZa3NWAp2tuHnbDS2DVNx7LHvJ2ikrlYfzF8jCgkp1f
BMZmdhHcrYReCkYNhtIAznze3K/xhi2dxvMCPHxMbPiGfbIoFmhE84YYUdNy/ytWSarg2AxxfY7V
WdrhjUdcL+Usg2vYssaCQ04BV2FS+Fd8aNUv01SR9kruxYoQi2QxkG2+o7Zq9SYBRNM1Wp8IwHPC
k3tzwlQix5xsqnMNdIWnrtlALM+K8KAAm+LS6wwpt/qdDmVRe9LG8O80Xb4T1p+KHGHJpx6KGJl6
7zfKNpRKof3xoO5brQPCvlhjJCovgzJSTV1bUbOaQnUXkLTaAxIzGGxokygWbCl1hjoD5V8uvsEe
539L+tA8F3NM1cq8Q+d3MldLeZrDQ7wHax+XkmCTwgKXEkBDGaXU01GoaBCcyD+LoESvg21vImf5
Lz0TFgApJLKKNtx+jfSO7g8VYZR9kTr4aWCFXamFSDI5dQG6aU5A+tx8vSlFspSyDljT15nsvvoN
sHzlnZsWYqTPXx3x8/xKPrxRjqP4PZRvK88ewQi0lAf5phHGjs2yEmACW16M/tte8nZ17sEZxsPx
8XBn+Ob5HUWZ8K7g2S8DVtcRMFyo/c2ebHMzfWDiQTxEx4ytcxRkvfpPpODGbcNEoy+xqRY47tL7
+7SCTknkXFb96JHqtS1uEVwxCNJR1Knpgs2SzXLYeOmGO50r70p1BTC8W3P+A8MD4cNITIeF7gk/
TAWt/EGzGGe3sJnS7YeyFgPT/semOZGUnW0y2nAn4giluOdKpntcOM71kCWTToHXqB79OZXNbe9M
M+hTS/sBcAOyoAJjI+6Z4QRMym4HZlBoPwsUwhxNV2BgmJXCswRQfjTD2YDFSTlc9QhF5rYT5Cj/
D6EqhYWbFR4V//EuAzLlHA9rWWUnda6WUw4/wUBTN4hGmmu1LTr5WyFha4iMTvzqWlHXIYkJZ/jk
quL1uE9m46VYKp4jLjTfuuYeUHzZToCQwuAWCHKToW+BtON3Fh92VHdrRfVv5AkPGnOdVnEKby80
wCqaZPXJM4wXQQbHxzI6JLAr9z6kdUlvN2psasA5pHTUginRdhREM5tcoTAp0TDUWflBPU19ANwa
qwsYtVBHYpS+LvLgqTcAmPeVJM3jnmwb7zbI3MHilib/Ddx5E7mXLIziDZehaVC4X8Fh+kGb8urX
EgspoC7f/4I/1aL96zMDVnWMZzoS0ORQEjwVNYXawjAAicvH6gEMxH4Bx3zOTLzSrWrAlC97nhYO
+EWgjW3LTbjBghbG34q6NQ9Nfwr4rAu5H0brlp7oDuFkCBdFocvyK+0cX78GrXtdmx5Ht8UdHMwK
9KWv8eOEq0vC5+vGdHMbYNlr0GxK3U0FWlJJ3TcrGGejPzbT/od1yEvqCHf8mtA0Z3iTnwvssSEV
gxtZlw78ICEaO9ar1WGFFen9c4mMVllr1wkMH1Ixhh86qDaH72XOkNv2qai03Tkfyh+mvSJEhSlu
0bSUV4CdgWMUiBgaidpS4yhhqWejJK8dbfdVjvHHmg/TJM57aP1Skjzeu3LBxAu2cfni5jXnc2G2
QUkQOfvKoRA9xjNld2/jiUjkM2gHn20+9oyGc4QhODnmB7+U+N8Xd0S0x5wmo0tkSuXHbsQhIL0A
Nj2wH1HEGIULAdixXpDerDDR4+4VcUECu+S9/q8osLzJj1Wm4e5nUzAZBoVyYAXvu4qaMV0xK5Gc
t7cF3Uvrf4f/OqypRO3A+LrjIM4e7rvTNsgNlkFhyGN6zu+mkifX1zAciaUw4/thiNROjcH8npf/
xOIpyfXj7MdFSMOiYJ0NPdYlejWRsDNqmU/8Tcjp2DJe5oio2KK2yIu1sG/dTtxBF0QBzj4CqfJQ
1KSeWp8Id+EptySpr6V/87WX3CBSlUu2aghfE/qujJTmflg6/PLXYLR63INP5Bw0+KyUgs9Enk81
YqWCeXLxwOwwDH6ug1OyyZc9fzXaA23mb8cP5nnHjnDtzigYykKXqYVBy2S5h+K5mE9DVb2FVM+A
FqUK/afzeZMtcoqSJaP6grDfI/wedW8b7Fh9flnymt7sa0VlHJuWlKR3g+wnVgUMxrrtUVc1OAF9
LAW33Hz9hRwt+wtFDMRXOmkbzJF07VoCJ7dqdCNRqY8/8MLzwHJHh9llvfIye/lCoTYJhaHnHjNx
b5JwUsNXrwFiwuY8q7l6+mXcRpt+HVvG0tXzEJwZMLBNe90lUhah4wq4FhNx16H/DtIi3MTrAzLD
SfZQREMfKrzUqvGGer05msXkGoRYw8p+HfUfKKqGkTTKcoSIxxwkt5V4O1IkF7UAahYczo9eW5cY
DPKuPzWE3plbLuZdx5LaV7YzH1bqIB3tePilGozc+ltqs0zKCa6JgyTDM8w8i9GuwlUDOCfwhaZL
76YzoFyAY8VCHTOBEi0Ft5kSKKzzFOZLnstGz1Gg/pN9A8duxvMlxyRCmhYjOYBImXwVWKRzMyrk
HbqTvWpj2vZdK03qsW/fRpgcS9NYfqSmDVvZ1vbZuEC2EA3ET9ouOC7Hx0xhxVJeu2M5Vjcq9+HW
M2DFXTRgiPZ4il9m6uXnO0V/KZZ0TRK/03S3ghIT41TLPam2J7CJTIszfHPJ5RTf45+viDIMQ+e5
aR9W910+a+3cNYxWAW+U0tZnaLCgetl2HWW7q9lJWm/xWvC8ZitCdsPHH8Tcr/U64hrX5SNxuOkg
+RpvXND7dFEuWSEy5qsoPbmYUBLSmcaGYJV1i1PMO1oyyzgwF84Cdts4mRGUDVNjm/blXkk0itt1
nn8yY7CA7XVMNzgLANz2RUCuDniZoDzYVZ/+t71+5YSAEZFBkWMEJ464/U6RSJkHYhPkWoDpdXb6
e4aiwaptELu4emn+k/wqcZq1sR3FETrpK8ODjthapeLJFpSWVjCxdhbGcOYsQavaPto/oqfOUEky
0pEbPO+rTEekhwM9gbnefG3T1oKN22Mq2sbST87IhClyqRi9bP7sUwiW5EKgz+CJTUG9kSLPfLGI
Xloyj0uVOuMHV7eVIX/10cL5XXwm/zfNJXmostGWe+EX/GkRzDZiwYhqX4NrZc8Qq4nEHqKqo8Nj
cZ6u/Fu9eOJddq80OlFNH11shejCgCeOFX2tel8G6wxQLUUm3Zr+5t+nqMnM8K+SL0nHXXBftZG7
GCxjAe7yArsaSqH1iPTqWysDjQx+itMFZ32jUrClCXr6QFreRP5GNhY9t8Ug/YSUCuZK0RuObBhn
xkBnVXXz9PSflS0XcR3TWU29aSNQjx3X3cDvvRjYVMoEXE0RQOtN66/O3Owd5HfUNA3nm6QYSx1k
MuM7Ol3xGU51orndcBJWSUiOWJKnEsKuZmhrslDkfSnYf4oZgz1ckKNztrnKERj8Vz1Y758e2dEP
TULFq+nnQsW2+KIIqjjj9SF8jg/tKMG81GC5z92ehEMVmEAC9vQvgQO4U+OxyXRhJtIQbbd6uTfs
X7aO2T8w9N+axcju1sv7Y98DzWZT1pMtiYblume7jTnflEwIXg1E1ntEnKrIYA+rlJCCBPSgO8uK
B3HyY6Wk8rX9pLDAEfN9RYNN3D5yfAnPjw0125bVxKRtDfnlWH3rtPf/9esefXzGahnqH4UNcTuE
d+3WcLAKMwh3IlrIVJP/VUBqoOwF5b74ro9Gb6HoOiWWAxHs8/+8H11BZ0IgP1mpy6lng/LdtME6
2LyIWkwYbrpueQBT5I2NaMhfPSn/rfqMaer0gDz+670V51rCAotgJSB+/Hw6j6L5M+GgD3z/7n55
NaPxuTs6gA50JddUdPrj4LhZ7UzD1c75uGI9qrgB16/93CLrbXvcuqQHrzIZx3gxqWmf7I+N4ltu
I6xm/SNwoynZcvDwdjdyUH6VktXES9QNnUAQsnn0Nb9d8c0hnX47iErMvhkHUOtH7ZLnRll2UIGw
0M9PP3SRk+hFask+gxFrG2AbMoaFyBYsysY38qSlmxpmpjdCUNUK2apdOr+qaN90G445tInXIEAj
d+xfZ84WuJ2aUSuG9zdxczepHHXnzcIMDjfyUtXqYzBT1sVxcwI4NJ7dmVgi1ylScpoZwvByQsJx
0t8O9VQJJQ2EtIB2tmQO+YhrKJTvchjVPLgg6P+k0ds3Q3a9kfntSHR4jYG7gpk9vnVvjo+GM/YJ
8c2uY7CruFoPPY/mb4+Ic7rw+130ZXNh4VeGkYaMlQa5nsN9G5ZX4je2o9qsNlblefSjzCWM/62s
7NyDwoo1SPc7vtV5MbCQVQsb57xSPS2ZhufkU3Iyxz9FujZhckZ5Pb2IGswwMDXMeaJIaNdPeKiC
GdHGOpOvSspCobpKY2RToKCI9Q1uQR8FdCOTgtiQSMTcCghRqKc+XsEVIkjs46OK6qi3+qSbgBA1
teiDwxumXaBbHecDFkmGvkQ/KkzB43N6Nxd9mWqVBJu/gOTNDicFRS5KXFktoYhtoG1dtyyCBxLj
wQ5yAqA10imJ+ti8Tf3raX1q17JzZZFaBaOHCCSstkFbaeJnz2OUUD0+yteQtZnryztzdeQCJF5L
ycvFakXL7oQmDa7m8AWvSvEU/Tl1MdfAW5A2QjADh544BZ3Yi4yqiA4Ivv8g2KuUA62P+1wauaph
pTTk6mmw0dYQky15KBb5D8/wptpAOFJO4OmF/6mhZ1Q+Twp02YB62rl9CuxmSsypk1XBjhlxZ179
HAZO8IOmjIHDjf+xKT1NE959ev90Y1mVTFjixHSMOK6EysBkIxKs1t/dP566UnvPLafX/WR/MCea
qCVM9l36F+ShMdXQRv1kH9QF86UdS2apM0Lf2wzq0i40P4YuHmeVARkOtz8cFZSUM9h9rSK/LZD8
dLKN5ucEAZslui9T04xyPimVRnWh8JGnvuvzwQMOFvTT64iQ1JJPXn5+dzvs0OQLVS74vPJfru+H
ZcAKw02MfUzy9TzlAud9OpM4thvOF279Oq08UT+4ZKfCZsOfNdiZquJ9PCQqgzYTGbCm0ft/1aFL
+6r7txUEA515mcHsiqoRsTjqDgzKqb6414C5zG42g/ZPM+VJaVZG16H9zIu6fcmYmmpnVvcp7fba
YECJ1WwMKaTno13OYk6iWbdjai+/q4P3YO3JyLAuhMZYBhAoa0nQDKUfBh6i2rt/OGMxOxV7kfmZ
uwerTVCxcEgSsUtAmWHngSuYt3szsnxmuE8vE/TirNqRQx2Z6mqF6vfHk6lN4c9XHsWrhVrBq15v
yKgHTBbQSTtUHQ3RsWDdXL4EbGf5P1pOY+EMZ7mgbkVT1oZNeJ1KBqe0f+OOrEQSWVOk58bFwAz+
MmUmFuzy2ebEZAtnjqGXN+CMABhSeSdghCN5k77EZPkeE/8PtdKSuFete0dnt5FK0oI6wnrU0nW9
f1ttF2xyacuAOIauZMLMtQXXeJY8hhBwH+5G1X63Dar1osfWyPQa+SNPZqvGTUszoXhJ4F2PzlXb
TXTQFr9mgWrSAR1o1LMLJU/QzbmslhRvhJ92/PYSH/rBRNJGp6Nj9SSSVM1ee6G4AMrKq+V0fE0h
1YtxzNmPuE9lQ8o/HQgeo9lM0kGbtQERorXbi25IEp0hi2qXS0MUVHk2SACxxUu6BbAYGflaYQtG
AK+4cHlmqxHXtRL6I4pM+tFq2k3IT/W2sHTD3bQp9nY6QCS+1ZQ+xK2nsWw7FAqrVNCUR2vSao3A
PeD04Qs/QNbE3Ecku4zB0jmsIYh9wOHfq+0ZBjbHtQ9sGjeRgMsiKjjJ8CnbpoK/fig8lh+b95KT
7VSIVmuJnuxCHDD39NzL0OrMYfFUe2UO9gqb3K5DR/vMV4acYFjjmvy2GkX0tW07pEcXJOYoocwV
1qy4miOBmHC8LnXa9Cn1+2queVmddkvGX9vu7oPSQHqKlh8qn3nXO6I1zkimAhptsACWd5N3biDe
Opv/KB+vUaK3JBINFu6tKL8vckOnLghCWSqfOaCKd81LkbK+odE1bS9GfCkwLoscdRoMkIRVvanD
kQpHg63cu/0ZOGryBeEN+cAVefCBjxHQhc+Z6pi7KUsHzN0mq20Xz8B32QBF1ozoocDCkgo/zCtJ
ktlkwyDSVkS3MdWB1XpUSFQV+MWAMBwuxk8mQzewPOQ2Z2ZljFFDXb5EnWdiRebeeXrhOUGaPaGX
rTJnF4l8oDipcguXjM8XH9K8hVO2FOmpBCYlQrXCKZwL0wJm19cmaBZZeFjncEanDvyHzEIQc+GH
tl99S0+NBvE3H+7Un72arhTo8q0Xj4zy2vUYBY07MBvcrMJ4k3j6988cOUkI54d+j8YJDwTBWtgc
a7uGcIjtgIqlRK3rw6qfD7Cz6h61jrpUitxmljpmoPtS34c+BSgp3t/N+mG6CZPCMMTsJ6KBsyAv
aNsXKnkOurnQ7ZCbshwlJX9Obx2hI26ZELstIssn9QWWHIUo5xZT+P9RDxFT6JuDlL4jTwPz7piM
Pdc350Lcu/fMHRIvPmh55971Q9ihCIy58/8MnZXWvPM0REJQoTJ5Ty/GY1ipkpzrdlY+nShafRjg
i/xuGdg6GPUxwoDct3RS4HfbbFkY1h67Ny0eSNQjXuG38JMUYCSdMVD3ZvI+cK2mWYchWQp6Js+Y
bYQtyLEFBdYkkhQ+SXl3uGeIC+yleB298UpRT/5eMmF3lHuYBEkfFGrkdFFbv1wO/q7n33BBiUjX
TPIJ0JZVV21lA5+z6KHPp3rkQ9VLv0Sa9zWG3R8SxuK/24R8uWljc/b8A6ootJcHPYke2DHA8me/
n0nuji3nxFcsSP3D8zCsDliqoZknAZHL/DXAG9GOmPrVwDnIzKltrAJYT9QTzMLaP4cRkkbLvbvQ
lBegoUcbAtUijkGZMslsaV90skPr0LQbrz9lMpgbrBG3lYuHcVvpMMuvbNxZE9e9HgnWHF7akGS0
zqoJ30yei4eJylqG5sULyeuPLjWhVPX0qwuMWWtNT8YG/fEhOpEvUn++fYWm/zlGGwfV7XBPxXG1
mkQZyGMEBvNaRhtpUicUBd+ZMPz4byF3MLgKnB1QaBVRD279M+lb5/OswKOH/r3FWIn9mH6PIJut
rbKtdzmlCuPnXB1OVdo8osTEmJkxu0r4soG6POCRGJFddbjLr4hqKGia9VL6B2Q8TDvsBREqm3gR
VwqjyoaFL5gITRWCUc/hnGjXLXv62opyERlRCE6slEvXHPl6A9KrrmVaF2SPSk7qopV5OxQ80sbc
/oVzyuKq8iNi8eQmv+mYyT+uSxu3iRb/FIEi0u6Q/aRyByXVOL3fQ3zhtxXgWAmH727Fw13iYXHm
WuXbFuxi/zNq/DvUwldUWDz08gMclxiODRnYb85KEUQMC/4g4qEWljdo1+46uP+HVESR44hhQWVa
IpQeLDJAGLozwTWOvcsIz6XgH5hBXXmIRKM/Q4rFgR8iZYR4yxz1w5Z5Xkob5ygGhs7JCB1BfvHH
fdEqi5Mc1rV2ozviJZWGvFG8YtgH798PPX8fQ9Ur1tJgDGGYrccWGqHK8pgrQYLno75Ic35BLgTj
GqoIxQv6MAoywrTOoeJKlJSs1TKnq/iZcvvySfRJ+ZJrSldvAADr8Cr4FzUh6Gw0/fbwoMbNr6c9
JP1cERZkg2DvfZVtP8CzWeiEg2rKAn11xGqtqP+vXmo2k/Gryu/lVWAnOVYuZevtbTdYIekIdge+
AoE8SX/qVM32QUU2FOGjE0/Rdwfg3CCqQqGUv1p9Pxupqan4HZBVORfIoL90QwiVJbwrdOPc7FPS
2xMHV0n4K0J3AVgfpjDh9L/QFahQoZcQ7UYS2virrEoCALGivay1gLD+2GRcDZikOk+a2vddhxv6
/cGIAQ3ukQgPmVIMZOLC4R+ocC/nVLKU4NOA53rAW3k93iDrspmBIQknx4ZrsyjDhdoI1we6t8V3
YMIvOFFsGZf8f4poGusa19W9504CuLhKBNRdANJsU2xTRVVcDkRHIXc9vN+S8fgp15UPlukNCcKB
c6nES51WY7yZdCbwxwa1WkGQ4vT3LZd60CflagonhnLcKHe4f0O14ci0+Z/THpkh91J83ehaLBVc
+B8cBmaFdMPwrWfWVAmL+xNeyIKpD9PPZJTzG/N62aaGvdv4CDcOza8MVjaQvhkgsTny4y0SoUZZ
WUmuG2J6/JRYgWzfJLT7omELWtOSnGzxfNgVAeEecsIyzV9PJZGe6Pe1bQxh66gibrg0UQHIWYbT
m9EQ60kHzOAWw8gP1mf5zEULF7tbYTJ86YI+Z6SJxDpOyR0Y70XFbf8rPUX9n0o1dFgw9vzD/pAW
xHbzS6SkkQQulbYbk5SEXfm70fohKcsB/ZuGgpiqD6Kv7oCGG+m2Bt2eksH03DP7mAoZ+UkXVQ+O
dF6MEOVjh9AnggokpRmG07CMhBLnL58NjLIV6Q1I0kyLrLyQ2VClkzVAJZTJjy08Jq+E+r/+I/+x
6MimQmCo/l+wtisoMm6fN5v0FfAGmvS8+zKK26TB5buhTp9Q4l+y0HdwCvwfvxt4ubeHMCllPEs3
rkoxmNSKHf2+932kigpXsIU9fbHNWuCg5XGDJ7w03UulmIJU0sCLpLsPz2ANU4t/VeAJ0BuLz3ze
sxohfULMGsCaLqtFOCBUgN9DWxrP/OKz41pbJmN0xx6MV/WF99XPJpffSL5HxO4WgwbHBvIjLKoV
Oi28EIkp/eNH1Sk1g4rri+kXZZ9WfSSNrer24LB2WiJq0PeH0HcgETddiXeHKaYv702tjZ7tC01r
dk9MqoYbTUKmhTrlLlwEBqle1W3IGbc/b1iPd+wB0z86wjeCUmtXiKqu2NfnFY8fi1EOgh5jLRR3
0GDK6NyGy/Yxlqb+KJIbehuHpM8FQZ5QuC29MHbhvZXf0KnPdn7LUQe98GWUdlYMLCzBl0sRAYTP
wn7hlcDlm2n/QuX+8u+D+tQ9CWyOsfqHic1IOHk17aJhDxV7vA69wvmsISk2ZwptOwZzK2dftJda
ObjZ6s+b+l273WJhTXW9EPyuov87e2JqrEoX2CGrOg+AnP6bg/j6Pt9PEyd6WKg8o6bUGo1kLvUo
gM0Lx3YsD02j0LsO1LAPirL7MrA/F77A/HaocsKFHG1R+4Bz3syJvRlkiIZi+r90tWP++8tQU5y/
53OfoFgZYV6TAxGIz0ZwSxa5y5KIUdz03XoFynHEghe6gonc9Br4G8qp55Edh2glSUu5J9Hp9oVn
uvGVLCr76NHLs2viIPUVsgQ7AVRS+Ao69jd+Ak/LjXdtAJjGryLNXxTrGQavtIYR6Bi6MDOyGGqM
vaAgARG3uDfu43CC9HZux+40uT9mZ1vktjd3SEwSSc1hYuir7MJsIpSnQj7twrxhTwicHabLWORv
JJxe4vl3GTu+6xmQ4FQmaIxbEFCW1QieE4Zn6udz3DqhjpnT4BzYkuFoTrE/KzADky73mH9nBmjs
+fA7AIek0CCqQNMnxF1Q17cgmhO/oO1WDOLuG+t6hRrzAgUOw7KS2wHdmfWwNVCxj1ZYiuRewWJo
iJpgwf1MZ1YljyTd5RGuRiu/n6MnH3oBLfC1T1VFDutQWwbiNnr7vT12vjgC45yTKanzQ77bBBBb
1P0/Xr7QHvPcXIu3XED8eG3shN86DpVOJydCgaNuOODeDWObByWPWnAnEIKk0mqmEk32GIcXk/d6
cStRnJlM8dSXLpl6GsEy2/S4fShuwmxvnC4k1uETsTAdl17groJTlQHt/fyFjLIVlyAWUEc+7WRu
lzecYJRmFuKsOLNYAk+PsK/lDDnteTeRFqApWoE/qz+22+KzZF1ZBwxUJ/ZKEfvenR0SOPSOBxR3
54v1qx0y7fmO3TdYeZ4mCY3mLSlnPX/q9wfgebzoCcENpBsQVP4mzs+spswbN1ppHMtoOdLaREcv
+i2r9xDdLoF/HfIwzvnGJxB7X3QRM0dwIlmSeKxUwCfD8AXDC4UGBKWAc0EDUhzsqELOt84B/WjP
jLtOq5UNN7diJcHNONjr3RSV952JMrW2qPgMP36tHXv1By1r4QkzwIMTRklurMhlWWC294anDX2V
f8c/MFS0Uy1VrV3iTOP5iq8kfml/osjo9Zpssvg6vY+DpnFEVZE7lC45pnCg/RsIN2qH5kU2NPq0
2SC3BuSUEFLsfWr4Rj5AKwc88gKIt8oS92axb7Zi1chLthfl/VXxLrNVIgeIc3/oS5mGSiCt4Id/
SIJcLKvEo/uQR6zLonpE4TWzhuDFVLoI17FUfYvEtucjqsSTE2aiPbnY9kj1/W8PRvi5aL5NBWPG
wHDpxtGdsZ1KXKuh/c/wfhb/w+GrW4YHiviKvDaApcqcOdZ43DoWHvxITbumMXK39/f/E1rBE5Hp
S2QW6U6Wgd7emzQijcXiaLdqUiut2rJY30nmX4ebwtwHcmwrRHplm0jfMWHQAAg1in+m9nE0uTva
xgDAmSUrGDRxUFGN4mBoxYtS4ICyKQn86zuBxYpfS+jT6x8mHbog9zzz7X/li58V0Gz4ioqkVCDN
d0oAW+tgNuVY9rmbZF1U3dplDIQFqCtY9x5736PxXNKbGv+oC7JSQvLqhufky+tnCCH3w7nzAgR1
5nLcv9JMu/qXhv7VlB9CP8zeKb4O/X2hVIEKiF3BWl/ghOGjB5QUI+sooIiDQVNt4dlQ4xYTBqMe
vC82oc/m8kbsqSQAeghj/2nSRMvRfSdB3+SIZO15lv6M6ffE87Dm5QvBNYVOmB6SCjsY9XUWj9JR
/M232kKFoRkItUWOoScU2TR/rugRKk/qVtJm6/GZPUHSj+b8aor9/B3+ovd/jqGTPGV1lCVMlV4I
IxEWySzJtOSxtpoAwx4lnd+NQkHw3vMLFyCvcVs/4FHiwilL+KrlDyrV7Eee0pXqPXUxNaMRMYca
OkH1Eol/SaHMoA+jmfdyMxENHP8/Rz/2S5U/IWxasRPlzVNftz4ql+m+gAo8N9gVhGihHFJ2gs2B
s7qiWFQ9d9w3ZfVSvbsSBzoSn+CgmxpafJCZRiErpkoAFhlMm6UQAL5jzHGB4jwo+tm7Pf/noAdx
7XBFNkMALAN6VOJcoNtqCAEICFMdx35EK2MciyeN5KSRgH022Yff4zFgzUaILrn6LwCCrqLs8q+Q
MOahOUL9fiPpR07Ont9/1pnOWYdN2kitfA6TcZuA1f25XCMn69kd844RwylVSLldefVwEWeTCle9
mbULJAJic7NtiN37Fn/mojsOoi0D0CE+lMPI0lXw7yfMd9v+1VQodYojSUTQDUdUzjxAQnomfLdi
8ZaOWXtmoJhso57uKPot9MIVIEKrk+xQqEB5D0sdGaM3ewYdcrVHGK3ouZpSTkyps6ZqrFXljfGL
JM+F8WDOr+e2RWDwq1z6yTt/PBCqJmZtPk/Yuz+9m58NH5SWmdpS/yaibIwVvFT45FcNAev7UOP+
kN15VPn8kqmVP7Le3STvOgxkMiszQY/qIvgdqXCnUdmNxKY+FyJ2StM3ImO/fFrkPctvs0JD+gK/
Rc+obDKgl+ZEYk3iPf/SHVX4zvlUEkB+Q2qY2Zu36ql25oZMKnkWQng20Svacj4sdoOxvToauzOD
dDNfoBVIoJmPH+GAUbubQ4B28cdPBNb0HsOJ/SfttiuZ5ImR4DdKHeDmpC/bXnAQ8v+sPOIzlU4b
npx2BPby/f6tJyNoapoR2zwL1a4zWGInq+0l6cAGEB8v1OyL3eZlJxUn2sIyoPoT2s+gZW7GAH54
rID6Eht48hwtOfcCk8tnucP0fWrqZ5u4iEarcSbLROhAhUYWGkIOlDg9/+TRCsRhVSsxMdx8Zulp
XP5Gig0HSCLbjkZ56R7Uj+N1p2KdrAxaXdBC7yUWmPzgJza+PHX4TJ2isZX0BC5Ju1hQF7dJ9m3y
AtME0nHb/EO+nsCV5DBkInbWFo7MsAiiScYpNePunRuve8P52rkt7AzMFNkqJ0bWSeXaYOVgBtqM
aJnAjloFP+RR20513/mkblBTwhGGmbBrXKimkEOzGrJcU1RxRJ5afWDvn1HCLSv7Kss4go0Hc94B
m4/H2hDTe3haxn4b6NEC392HWz8kI/nM1fTark6mJN7QElYjpDeZxxRvR7HzigoxVGoMzyyIeCmZ
cojZOTaNd316jOx+Ba8RiIUBPj7IvpH0e8+kjj8sLyx9O7ge9dJgMehF6dmds/aSeFxLwVxtCDCx
IzB8SDn+QMFPw4YfY0bK+mgUGR4IOKGBIB8Zqjtj5mdFM8mtb/ubUdzhjwOL4OtPNgXt6nfYDOcu
thiIBKo/bJgRi+HuaZ/B2DAiWQs7+1RKK4sSjXtDOB/8/R3Giu7iqqRqBCSbHioqgOYlr6nUX+nn
B8uKH1LEA0g1XUs/EQfIC6jqFIwtvuNQ9byXuo04O0G3fXUq65eMu3MDSwGnRHBbtGfECvdWswwZ
fvB2FrF8gm/IuHBLrf4Iubus1x1SN/k0pZHJ2IkNNLuoP5kKY7cBwEewjaTfL+U5B8kLpI/2O2mr
tK3uHis5UYPbSQj64a0htleuf5U0jNQ0gVWPgutMkV2Ee7aF322s+4BYSKGZpZNoaDOsss6VCcHz
R52LgfGi8TY+YK2SU8J8iyrZKqRpXM8FSBNY1JxMiqNMuWL9LV7iVKGcpBSYsXAFhfckeXrOMlSx
QZAd+hkolxGUIQgWRDSIACIbyD96Sxgg72fy1GVMPSQqowmNGYLN5sOsALDeQFuQmup2mGssc2yy
Bbg7sxyFvSvgXYEVYUi49/eDpcDJd7QpyxdbBVECCM5/xntd7RizMtPd3gAJJ7zRCtY4p/6i6cUH
Rbcw+lbT4/MR2ayThuueO2BMQVuWG4dG3I9B6zugMG1c9SdPWczSnIoz/NcQ5ewsjB7dKZgYrN3k
vMtUkhpeqLtf0AeQOQJjAKW1KTLIyO6exMi9+vmYlm/KEhE6rxqzmrjZE3LNiPZPPzLf+R/BFyha
EqEsZ6bPC4t9YouqVxgHnRoqvlvdmlhnDu+IfQg2E16/3gAR2A+2GVyWnA4fEiwTqIupgNMZE63l
YXOzrFpVwUP5pc5gPVwHyaki1E+IJ3SMqVyzePq4Jv/6HyNlKgMrrJnuV77/833Sy+yEWyCoth5d
ZCz2QYypIdHsa4hb2nD3LKGQ8eDiEkmolR5FDWkTb1AQ7YgXWX7vr8nw34EtEAdeYE56jukgFkno
+jstPzRte1H3v+LTKabDAJXd7M83vU5psZYQ1gF7ikRmvrImageYxeFBoKmmV0pqq72dBSZr3kr5
FG93NGBE2194rMg9KncubKTQSZOc7icqh2m7S7XTyHHXU30zIkjh2YpX0aMjt93bjfSlV7XdRfLe
wANFbzChqqqx/fwCx0JbOG33tjvG+WEP34NZ6Uw9L6YjUXsqLetXFWqpr+6DWYr3MfjL54N9ZbNr
g2GgwnKwg6wcIOFTIwYLDirw9r/9MThPmzuHeoBh1i6B3pRJYHvEyLAYB+wMNtFnxknv95cqZ84+
ppaLEk6jguJkPqVlrIwvYm70U4RUcBC7vitwyLj6Mx5LOwsf8vhaWS+3VJMJyj6sckSKd6E/jLQP
XPVkYQ7KjFsQ0gHX4U8r2/2+zlfJ8+STO7r1OUmTmXEgNWiKWqajI/leNiIjeAiRIOmR66Te+0R1
1nnLr48Sn0kPQ/dkbVJf2gKA6dea+7Ii+2rF+nXoTvg7qmD8WrQSXrFwWnCmNfvhMnoiIFQZ+wgO
Mg/4bPnQU/Vl77qcY4b6SxytTEZ5xGezCt+x9wp2H4nGgUjgeuY7mtdIWWQAinVpvZIqaJFHeGL/
Xd73bFM186QyHxjdRIw6Fvpa8/YC4fxzc9C8AioAzigEzzgUwafys/7iqZPY+g07kwAiFzIu51Jh
RqVSamCX66RC5vRxGcCd5TIuDSEFXGrveWRxvBPpLsAEZ/wL2xgTyzcAr0UyDzWFM6O1/v1Gf1yT
uq/ez1xvF+gRpo3ycUwShZI7csnBX8a/P52n72ZXBbmf8VbtPN4buHZ+bUGBlg8ZVQ7LSnKEeQLC
X0CQ0QDJ8jbLg/JEjigCLrJbcZBCEd1rFRRMlfeAOGZV4nkaIn7HExwh0FEQ6lUKuownDhKWjiRF
PmP9Usy5KXw0qh617UZAvmwMcxJJiDVEuwHxOgHoG7V1kIgvpOwMg49rx3ZbCxOMSdTOg1iCuZ0A
5hAOaoKd8s12mf+EpAQp5cVthvtZaIHyrUx6lRR4/5TIDlb8iGnejFXnLVQHTlpfYW91KiESa8ev
ftFnwn99zRU5NiTQVHREhdXUNlQ/5oA+xKjMhXsKNzKti6IswbJXDrpXDhV9vnIAyIBvG0+bVUXS
UhetCydKD/d2y82b9xP2dfYklApf5FbfbeMNRm+qwPD1f37cpNdXMRA+ttZqHNmA2ljA5dFcUxTa
J3sElNuxXE6yIxjG/usqBJ6ZUF8IKnykejb2RuvmiMIu3NIDN18EvpWVq82tr/vn1BoM5uKn2D5U
U2vtMxfEYhZ9F7BQvOSGbM3HsMVfU0zu78v/5MMOmeSp3tSKcSHF2158HoTh3r3TPPKin17lTDSX
ssPZ8di9FGe0S7cMsuLA9Z1jci8mIjnTptwA3iNKxtmPINt4Y8ItUKXVmpkMJOX+SKSFRWrYbGzl
WPbLtN81czoLrU529YzBzF8jaAGkuKq73T3i6Bud+oAnLDysXliow5kDWErrPdypZPaTju2czGeg
WxXCa8ceOU5DJ0YuI+xvoI1+Q+fzoJ4Gi4koZv9mmynONwZwKIfaYrccI/fB6BpULn5PRQQ0BakA
uBHSXfETE/MrxZc6dXSp2y3VDguqV0WnNmrefxkfYHFWYFV7Iugxhf61Lc8oBjPIXQOqtf4apSw+
TR7qTRtsl7I9OecQfjHjVnuIRdAONciiMqRm5h6XJgM5571qGrdwy8vy1Sxz0ob/jW+UEIGn0kHO
ebDboXf/revXJS8OuMzA6DEyqWYoDvDowRTj4KEJcUifuEdALbjxGeLM7eOuBLh1nOdfcM/W1ajx
lC8uv7dMF+xka/92nKRbk73ObMszUmH7NPd4eHxB6lyn9rBEskm/rWb8HHWClWTFe74+fDAwcgBf
iy2Xwk7hU0yjSs+TwTHp5g+bba3P22QpzcaG5DAAvekEBYjl2E0BMht5YGAPkLnLZBYVIrJLZBD3
9dNu/oron8IITFMsl+ngOIyV3BChGry55zOMF9zc1QbnLpW5Jo7iv4M2Znr5+Yh9WUe84tvvgIt6
zg7Nx0WqAj8SpjRKcckBIHEPMtY+za217YfrDbVq+T4ntoI86NfSnb/Nq5jgiJWhiUjlcGyJCkEh
lHXPzZU1dl+mQTibzhzzeHsOovbnSJLrr23TLUqV5IQNLOgf/810D6nzDU5thu872dNIIw1MRMqZ
IlLbCsUdnSA82/pA9Wu10IyizgQ1yRDyaMtIFZpIoE5fSW8O+TlJ0z+Hx2y7UJntbM0k8WOjSnXE
7FyiySiA29JgCPhiHww4E0x+PR5M42Du1iiREvj0HUiIxr0V3N9JJDKoCQZbeXDzQIs4rP36bQpw
FkpAi+1RArLu8omwhPeszWv8JGCFQ6Kt1Tfh2vAemw88jDrm/tZyXt/ppKhkUi+KGh62t7nPCn0h
rSLUfXXkFvf4oNz8fuXuR04lUPD3utj94wjRtldBkhHrt9k/a7JFKJPLAQW5Ipc9YJpDO9mOaYPn
W9Hi+LDldcw/gRkoGfU8Er4ToxUpIuZyINqVH+2PsL3mrw1pqsFT0ha3uQ6aoWKMmRF1xvIA+VC2
rYLunUfVCBe06yBN/j2EoiEntJGcCJBvdGQTtsdX2qaJoLuWi0mw8Eh4rGYkwQbiS0EjFasRzaZo
6N0PgUHv1+NIO0pPXBndKbY4vfDJf3+adLnF4+Oj/Ntdi55FDtrBs8pkdUAQoJVcTVC62mUYy8CC
Iur0wbAERwoI5WSaEdaXADAb6udXdf52sVXR5i6xZj76+1HxTOtz2XolheMdHkKrxkhzZAZgfrLP
o1bjlYaghIPGoYB6DU+89KKcXtStVmaOFCvXY9LPQ9arI+UFMpXCkAXnd42hzkDwh5UziUZZgisl
7GGBqkvieoDf9reIlzojbLhz6MNiEQMyoCdBqzzq0oPHDFUdPFbVbZ6uRT8SCFZC5w5pu32fPqUF
sA4Gl+O2kJFhn9e7VroOpJv+Up0FcLcWA6qgBP7zjHNnKXdCJTfujYPAc6YApCqHpTeHat6f+WkB
uKn6KHMC7i5KwhEwWlWXjl8Cd2KLjHygWraY/xI13KaecleN9HXn0xA9Ar88MDBYWhOv0pS5Zztb
wtgoOqFI0w0rHVoDzCJiBfYyhVnJSnqiIqRbt0/tltjBZCH4WKLn8c50Nsktez/t0T5IMc3DwPgh
rKk0qigjLBTFO+nAGxEFB9c5YGdMkEvR5BQodI2YU61StR76RLckhZgWOxkvPNAdsGMrTNsWcalI
L9x66XChgoNl8rT+xGXHCcUM0mbTLbx5sb7uRCSK/bY7byvbqqNG4kzxf/RBpHEA1kfaImtYLYzG
cHEtPAIOGl5hGYa9ZiDEGi9qt29++PZoh3tHSUBTJmCLSCIdJZWbl4d2yOyQZ3dfOMCPBGkDSOI7
z/VjVROG5Fg90o6Gt9C+axRkJEbtuxRlz/ZlotHEdidqb+fiUoQDZDsVs/jri5mkXcg3l8epNWd0
uJ/wAiNOL9nw4de1xU+8HNHLzvdd4grPxTNA7RiuYys/FgoPa87dbHIEsL3zoWWT+zEfBEm4EXxm
nNBMkSBR9vdQ9AY2X82+vV1Yixl4ckymSELDRlykqrGHv6A1kgSas85y4h5QVoGhuOqRScbkXVlA
1rYFW/pfe6AyJAYx4XBLBvixHndr3Y9LkO2crgP92UtipgyFwTWky1i3M01N9lWl/A7nm14Kfh3h
dTJA8CiMaYFumDdifByX5k5l5nmmW72Evd7DnzNFWkOljZ89lp3XskcI/N+qMNNZQqDebRmFCB33
gOzSBAMLhMmC/zQmdCk8Eibgek/F/Avtf+0KZmN9TWMdBlvUnLmEH/WgTyX0SsaN6yCijToDoFOt
uJRecbEK+A78R3Siq2nMsProF+c1XBlfJwYXzX08B/dnQjlaIjUoRpjX+SvFb2HP3qsYDRIZc/pz
W/U9kRa3n8bdsXOaKbYOM8mUSl96WntEwGN/6k7o2YlFEJRmlH47MqrFB90n4V2RPdbTildL10WE
FfVoZjep7LM8kO96GoWNVaITwnOdgr6IIjhCXtYJK0TkOKvT0XvLNhniIwmNDuDk631FMtGO9oIl
CfApGV+B2PyNi+riJZSyfXk+FRA6BD2APCKwJD540Jp7lXmHgJELv0oggZXk6f+7V9hMl6e7SFNF
J6X63LQXzxuMd9+5dL1mOMkNwWXFe6zPu9VnYGZTzj/tUiO8+De+Ri0CI2HlY4/alI2FJ+MWTWBT
Lk7dNvf9xrWhWxRvGKKIktJXsMbqE8YDjmnyTFeARw6xaMCYRIVN5X+2IcM1WG2R27AJ+RwMNcGT
Ygz5/gVpjcPFMdvvPXYxg1siZFkljhDOMaJIOZaGzPbbqsqfqnoGn+WTF5Utf6A5/Bx9/u5KM8aa
hEh0Gfy5aqEaqAqc9End9nZ/KMrlnj70tAgk/wQ/WIZBr7ZG0yC98Ec8T1iDQPnE9HV/GU0/722f
XOSiSOVgesgyGUPxc/j1OBtPZJpypBvApmuojn1cNGzWZ5+nGio+CtKZE80kjNdntWxKMI+KnVBu
64vZh6XGBioS23zjLvciRvgV/X1mBDneKURdMUA8TjEO/8SGteqgJZISyKLRNTg1umEdNri+YwYB
HoIQ8OFoqVQ/AzX/UYK9MXvQfbZ0CULLzFCERicmvSfiRVCqTEi75PNglIWs+hRDXTE/p4T35ltq
WrEQz8RVFeuYs26CNID4GD8e9Cqgmd8kozgSvcVltjgEllt/msdK1feUJWrLE7y+ys5DbLyuYaz7
/OQWkdiclKpgIH8jYXT3cy3YlQiae8kK/GtXC8IpX40+TGTFkKuqd1An0WPD4HzFtHlZMdKsFPTr
nUDtTf1QUjrKA4E5dxcCJYcNwESa+PDxx6fdfxrMTDiIQAZIE5ZKziGdT5oUUzuqxX3hhhIXa07d
QEGb3ik8h51eHrS0KXZQyVtdZ6B6jFGgbH4Oe78DcyZWb8WIqo4NmsVn9w9wDeq83VrmPagKAoT3
xCxevMoB3ZbExdK9LAiBRTtVk3imW6puB3y0MfzRErdauLjR5ZUFiwwVUey7gx9VkM1ekojWyTQA
slfvFIDT/kwzZ7p2TBInpZanLyWfYwM8chQcWRa+F9AmxpypOrUEva7KH3BKVJf5bp5/znJZUveM
Ob73g4uhuV+JZUeuAhbLOAkJrHG9q9DzCIuskPIx4+x3/nOs8fXok10o8vqIZva11anMS9FeTlLK
c9wHzn1Uf0rbPvpHdhUhRLsfthyoTGCjZgkr6PeqNpmHCiDJ/k42/EIcCbD8tUpIJNfMmi4stVbV
zAodluFcnxdPuJDAmfKK+djq4dz09B3mFRz1xJvpuKMRzadrGLHEdYqSpFXHQf0keZ90lPSBvvJf
d6P2W/ALgGtI5Pf1i90igj1bHEjhjTL49jPWkGo3hWzXQxoxhP2poGgIpPyI7SAbomZfOCLw9ILP
zm4WAQPvhb1v4267G+c+OIhIxiIqS6Xtvixom/4M/gzgsE2Fr8/2NoHqomSZSN/RFCWUqxxy99pS
aVlOj+y0DFSmONlXofbP525l/MZP+oHvT6T+M3YJYdtG6j7xYS0qslaDPwigLIRdVLcqzH5K7dKe
hcbOIXwIWenTJ/UVBhlNNK4mWbK7rB5v7SfCjDSXw3u/L/Z2cKf1X3ZKPK6hF5CLCNuQGEbUnfda
SodO+Du1hQt0jr4zcNTIzPSdwWAYWMt8u1DyMr/rRcrQaxVHITAJQuN7NMyiquYDM/GwsI8SC36n
D05dpGcGyD2rsAAwPpPAPmqdGYMifNtknbZKS0DrtzXalp6OHEnieP5bCoxugAIDcsYCkiqjN8+8
aIP37NK85UsS7mtHI5o+DyKBIYkeqR/LkHw4jXmZrs6lAzkiac8fnqnuwhwVhjLmKNN8LKKFgYlT
ST+2QanNYFD304i0/70A7vhrtqgpzfOsJMGethWwSplh0vif4BD2FxU+fdct36FjLYy2kGa7Y1Fn
7yiXzc7aqd8+w+efjXdy2kSiLVrQX7/Z18z1OXqFAcnvaKH6wtx+fUFJL646Oz6hklVnU9EMeO7o
OlC/kU4eWfdl0QwobpB9HqXct9mW8KXppECzCdDdOh7zmh9uTAhCe0mt3q9ZaCnHMHj/R1hDD88W
arc0potq7hFYMzr4mib+fsbHH8QvNZOUppDK7KlLhKYsB0ZwvrWYgJW8pTHgG6JXKtmkKwuB+7J0
/oVyc2RXwMlqW07wBC1EhGZnYGHqsNWzOjrlV2XlCgYIR6ruPylJLemRqL8Hcit2adLzK/Cw45ls
wfEn6pxXuWC6A/CM6xO1ZwVF5wypgtNXQr3j03b1NLEHWxR/lKXNGYXhICgudnFoH8RU1dt0HxHS
Rg1zcitsaeK8gMlthpzlM6eD0IZhsLyVuHFZN5heYlGn+5E4tolMYLZWnv4NbZu7VwY5LS9Z1ZVn
cQ3Ml/d1oM/9uaD1x/RsYimdva7UTrEBRrjoU4+MxnxNPvdZ5nEG6ONguVLBVVtSu5R2lEaMvwkg
zhuT+jSsRlBwAhzo1fOboEcrj2e537R55jFc66cR6ydIqH2CkIxICzLEd5Nx72hM0WXt0judekPb
YCA5fEWn4GCPH6o++dJpTb1rQklpQzUolb8GHPTEJ0hQ9ku8S727qf++mXHoXXqkM0D3IVIAR1Q+
fEGzgfMa+4w6tzSqjlcuanuBu2fDOMy3sLagsYNVdIiYc/8R0u3m//cMVO7pgvtvwRB5tGrm52Jv
b/mvRZ0ivQKfdH8+QIwlpkC5/c7tbD0xkmkIpReH9IRJZn8LKU+jbcnGgo16NF82ML9pI8IKe315
Y1YGddmMbQTiULyS0+q8gxn5B6nE07eBlGC5SjcQ9yAuIOizaCzNO53mCFzOrGWSXSF8x3bg4Js7
j0CqmQZ7XxHZVOeNFsnfXEG7Mwy5c2WkV9qp6arddiYqu0txjZpkhu6NHL0ue/aIvwUnjVbOozy/
0O9pETCpDTnTOAbE2KIyUXTPzb34k6LX0kz08bkP9uVGEsBDvoD8G5N6VpnlC/Eb7IobPnBrBgq/
FO7qfKYDXnA505Xp1mraM5wh+aRYjkzypqW29T0R/jejUNaq1VA2nJKCu8Wi2O/RA5k0YgvMLLZw
Rb6y1K3nJcXytqJb0qPidEIU5cikW9Z7pB59I3g4acuXl88VkTaABwoutRZO1M3ioywnQgRw5F08
DLiIyxoRGXFYwrNVGWS4L7Yr+8z1gOk9O+X9N7Z5+S7WuT3otENfGs3F3e6GPCCbAOlrKEXl/Db3
CYnrEhh/poNdxaV8OStUd9t6psWhz6WHPz35SPaRFVEnB0gsxLhEsD2XS9Ra82IZMfzOEqbuc67f
X9Zih3o5lzjOjhqoDDvXmCknGOyd/o2qYC2Ip+Lp7QH+jQNVNkhDZ8YGDaoAVrFRx6zPvP9otvCl
+1rJybJ63jcb7Mw82797wItA8o17emM1IdxbghqNwv24DnHeMnGqj1ybRfL5ePoBNlcDvZNDv35h
iOelUgucShnhhTIsz+nOYTir5NhI14pjktIkTXREnxEWOPpTuIVhZxfj/3vybvCmWYHjo4nEZhXJ
T1FP66FojXD9gIAWmJ76F+s07/y73RH/mn3F4RUIwm6Bg0cdTIIwBSUuvAl1ONFPKWefTfvaYrA3
IUd70mRZQ8irmrMFH/CKIog+xNou1UqKFDCUrSW6RJDvbtYvGY3yTuOrRY+3b3x6yaQnQl5EZsJ/
dES2EB5k4JoqGyxJVp/91bqy684DuYrolreuNEHxyBKCOGM9JCoOTNLVm7ZeXCDho1w8v6VAEji1
9MjKor2L3tefJSbaoLtDiD30e/zJ24Bp4c+wLHM23Triw1E3La0Sb4NRbQO5ru1ubE679pYJghya
oH2GodOi2oxaxHkmftDqpi0Ot4amQb07289qr6TZoaGY2kJuNdtzt2S5dS2yCZ844AvMryBbo8gq
NNCbcmkVAlyjgr8DAHX7HOTnvm1Byu6+eDzvlccxZuDxKipMMVLSub/m+rl14f+7Npf/xg+VMptE
5QC3fDKl+qY7eTMyXKy6NnKcbbDHVGecE/Lx5Gfe1ypvxk2UOn9FU7ukk/7XIlO0hyj4sl3ewOu/
7+BKyyFOYCZgZyzPODynIqWXBXaEH36eJssUJt1ZaCFR7tg3Cqc+yLd36aouWgnKYiPDFEczqpVl
cWztENtrBz9axmot93/TlTobmqe07vlfnbiPnYphRxmUwu7b3oK6M7Imwup/lrnvdPN5+urpITEA
6cHn0craeuHzEcEe+/MoDx+QuBe2MIL7B4dY3r4FA0r6wUHvzWsgE4TeAS6DueeEat9cxERQM9or
GoFC62sEVB202lC2udOlMhFKUJOgLzPAHkV9hv5EYZfDo3SHmZaKpGf+xzX2MESwfZRaR48jovDp
Q3oP8vGHH6yCq3K5Dl3/iG+3U6pNKjcBTlCNTu6BEH2XU4ekjMNLaukzpbwpvEmw0sh4KAo/EHxO
UiJvaPare5oOWj0G3JiOmZl47m02No1VgMW0SErHywevEg0IfEC3c1ozjSjF8ADEkMBjoBPJXpIW
khuJgTMuf4yGICCsGnwzsp0em2dyxcFTwkfEo8/w5QYM6JYn56vd8tP+yLMUi2bpk0ijRqRk7DD+
ntykbPIjHTZBJzQpOpuia5+VjmUqR7nMcJxtPUg0gs/Q/X31m5illMILSg4ZNJRlBeqgUvYjzmIs
7WY7eHDcFyNOvBJB9NcxvatTb3876U2nBC7UNsW/O+vtcT3oucsuV1Wc4eDpIt8s1vtsRnaOFNav
CP0QN6//ykhMwnR3EdDE/+2Wic1JUf9TxoVX0ESombUEr2d3zn0EDzuBU6/gaLsOxjwIkxtTFxqK
+NhcjZecumEWupTlEc/HX+pTYK80twiLw9hynKaGJo14cqFEAV7HZ5sCTqHtx7wYRPlcpdOANRSl
cxqz0dHzuU8IY2E2Lg0tpA4RdUJ5siwjMTcwj6u4NMM1mk8X2TudyV4TgfhT7PB5B634BYmBMU8o
jsPoFVCzN3DDUCSdHYNVWXgQPF6ExMGMdwRvkjT0zUxs1dl2i+xiOQ0vX3NkAtYZn8WbhqcKlNtJ
cRa+8kVzHgJFFcX5nYq6bB9QBr2ywPlxmvb6Kie55E01xW2ruwVAX74qqAK4Zoj5Xd39uiBJthzI
krHaEnfWZNHxKTq2QavFYfSnRalxhobjgFyKLWmmxh8oSJ3qZpoR60NwYDpaIfJ+s6uPVWtItA0k
voxpGElEdaVZb51Dt9H/ZAEPDViHNrOdHcp8VPk1pdtUbx1QZZ1WZJnbOXlpoiFA8SW+v80Xi7IS
it5Z6W1KX/kviHobnVSUCDqYiMndMAzWNDvrfdspMNuu79u2k554iSIBqHszKSIXhlK2+4FAkxmH
t/ZSWrpa9cLwfPnwvOvIx2fm17v8nWQvvjF7CznRyLch1f7OnKRhjqKtgQhHS/R0vJCq2wwTZazZ
B68Rfxnq7hnKpjFUwHzSejB+ZudNfFHh6Pr7Q+6uBU9rEsDhGpAHwT2UAF0P1lSkRAhFvG5G1OYL
ki9zZDK/4b7TtMNvW5Ci0ClkMBGrZxwDDxve2bjMv27uGtqxhqo8w1gwNaNflHGtUr/qM5tyOcz3
eRZBBUl1wCMtvV4JSicUud9hQtcxU3jpLyrdefh6UnTlP8Pq1gbNRS3kUZjiDid5iXfCbUUXQITU
hdW8HGkwhonmTfNpYFsjLtnbD0wFF6/PQeh1llCiK2H8B/2wD+Oy8VBevTZkMCIGvt8qh6m+iLwI
MAYOiMf3PRU8WgoNsWyiIAqvnGIQfOJ/mSJ5cU0EPhjlat/lj1wlOB3wil4iV35hj4LLgyFr33jf
aEhpMWZZI4QMgZC5Cej59i3a0Ya5x58rrOsc/pMob/y77h1I8LDPoWdzPVaacZHBbeUx2qBPwbYG
vu4lXw4DCw2SaaU9SRmGwnEnVSDFKlbFMo80rLy7UCDcLGyJCpmOSipsAlRZLIiQCu5n/k3KeJzk
UvTaNvCnt69BxXSFDv96vWaKeNOBTwZPzBnrby1HDwP3BvIvNs0TEhzQQuTwnxHvFRq3dvrv4Rhl
Z8NUyDfAZvm+Mjqn8e3fvCHnVYq47AtXTWmhU28DE213AWd3sYNQlWT7JU22ir5Ct40cTbO+0ErG
GOF/zdxK3LtnN4Bce2h7rnQyy/VOuldg3qVGJk0++4m1zIBuFCiBfiNjfK7pp0Oi+RPbnwAa5U+u
1HipMbxU9BzPJqCZ3gCuQ3Gk9W1KjFNXnSgeFNoThDBgw1upghphxkLzXCGMVS4j2WOI9MCuS3VA
V1SwyiNZCrChEp2PrfBvfjm0aRNlBlMyTDU54rIHxIXbgJwdlyieq2qgrsN81AWVBELSTlAoyIDY
/Sz6OoEN6uMoMspbSsrTKSpDg6H4xQO9DQQ7wDhCh9oRYNXrBq/Z8FACp5NrZoFChfIok3L5vIuH
1KlJu//0+d8fJXZQ8BfoXt84FqwvMiwS0yFxTMV/umelWyaKHFQja2ODEKo1cgplmLXWwIgcewUO
ofoZPTByw5AOQVCCyCvUlb5NOgQIyQYaOqdFb40tAE+cxK3DVwkdxN2hAulBVSMw11GHkRRvNT6A
H4j7eSO9IUmm2b3iXYhuFaWjLRn3LNRwIB1TKOPzNAK2PcyVeg238BffKmvQxDvbktedeF+QM8BX
WJPImuxx9rOiEprnGcC1EjYNTl3dHo+FwNCRJFrfSWJ4WAakb/oiBsTrDwcz+FY1dla72/o=
`pragma protect end_protected
