`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24096)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeybhskZA9S9tlfU9OcWLp2F3xQfV3HkcbFFKuniPHJk9WUS0c/JSGmLpuy
zibMaJ0wqurW4BmskEDM6CFKgFDEY7egXvWHVRBpY7eGNJ5t0t74Sefa/OsWk2MEW/H2nxNxfHGf
3EvKDP1QqQHjPODzWvkHH8CkfLuqJFhJk32a+WKLTTC4WUv5um2a0CTINTd+2vfs/22GcijSY1NO
h4UeRBxq4rjQs+EsKNiTPaK7zt7tkS4L140F2CFgw5YCzf6C7taZKmWpBqhI6YgZEbl40xszslf8
uSDr+s4PpVyQWRSVeUoPjoY2vcS5TyjaXiF2g5LTOGMVANZXAUAM8azmUlCvarxz5lzjOOO1orEf
rusMqw3wO52JIjGZfoO/PDxF1crBSw5eqdikTGZ9aIhowakNtIZjbFgaQeCl5GWjx0FA9R6xcx9E
F4AJGOIp6qqT4J2AuqXIvlcjJfh/EtCzN7ryH7nrnJYTSXZP+w0oprCDmNSAAe4HdRS3LZALmn/e
VdcTCLtSRQ9XhhlYP4n27VRxRSlhuDEgTdVD/gUwAHovHvyFIFbUP+FYSSDuozqzc9IdwEZO8ysG
qV3+y38nvYBdP/0/GhioVPfZcDnUHaUd7MO1FgPzpX6suB7VUgLcFmxcLIgdKIJOP4w2gMiWt//L
vnUJxsEYiOsAnDJ7d05oXold9CP3qK9Y1pZPXB2HXXGdOo5lacc5MDfYUwrCMxXs6c03/iJomgN6
c3JlhYigyrP1EAgDNKyrhEKr/0nNL+TbD9TFGueNnnyc1clPJ7gRQDP+EsjeKuuQmoKRRtcsUX6h
yExWTugsO2ZJC9ercUmJ+bYl5uMjq7pSF0Bo/9lXiPAcHPZh/xbqWTvBdmJlYpApFCG3mWXRtklc
GZIWlpxAPXUepjTq/3Iv8fvqTRv0OBFL0aLami3+kWjlnJ5bknBhtqsEt+eaInBSdLm6bPlP/ofV
DrVvAGXYcIqro0UtKoY2NzvcWtF2Ij8LCN54XhI1cLo9RNjfPcvgDx9aVbt2LojKqr8QRowl3X89
mUG/AXRg27Wd9vzrdX1YYf1+cYbPfpqs+1bRcgDCEskYQ1fnAMaZjbXTeOBlbZyTwTRYTk9KXTTD
cofVU18oJHQD429X1iwJpfchzZKxv1jIs21b93oImV2y6NtdIe+Hd2rGxymmnV1+Alclyv4Bw2iy
j05C44dk2ifc2VWXe7iEosljZWFDxzDnNujmL9p7vfAY86WGi+C5bKkgjMRnOTMsGAbSp5XnQBgg
ggkIR6ocgFn00wq7wlSjUNgO7/A1IVN9wYpAdPxH+kQUYZ82qSvdsqg7Lm12qxKRXR1gCxpaG7w4
/NLtb2XSTrYaKDU3HsD0wSIRDJziuLpWSqMtAmo47tnf4/NLyT1D99uBxH3bCd1PNDU0frvoj45b
7e+nfvYMkdmAqfStlcpoinP4pXbVMhBgz5Fqf/Dw2rK0cg9G0/V/yxtS3s4Md1DdRttv4mIWpBcP
46mi31JRVQN3b9khbisajuFmpK7fZ2h0fsS7pA46LnUQ+kxY2NZeKVnVVXQ8vCeIwP8UxpRnT7ag
lWlu0HXQSW1G28mQm51qRqBbiSeuscs7wsJyLmFoXVsQmLy5dmA1++5PG6BWQIzLMh8GPl2Q+UQu
tTs7UJ3nq1O285offVvpW7Om4+S+4CWo4PMWelGH4bN+6/MWIP1SDD/OX4TTjvubbVgG6NmYCHZq
MDW6ABg9K3BArQtu0MY9qrnjsDpyHyiyHgDsA1V7yWevZMBIPhiFtZ1YKO0byEOj/gPioBSo9A5k
W/50BOfEBMv9Up8mJmNAW720cXLSdIZFTaIu6wl52gjZrEJsyr84QtH5bMa/16lrsG+B9lVKg+KR
5u4tgSwE2c7WIz6ZdwkOJbRxXMNRhtugdvRR25iaeYgBfaa3X//q6Wg2pZKK5BuGzn05MqngdqKm
jIL7zX8w/4V9pFlnBQCAYrARWyzEw+h33yuQfo8x5Aj9sIqKcSg9LdQmKXBQg6PDIfoKhwINDnQF
yS0eheXoALHpl9IE+OamePQ4RfQO46MA66JAJ+PW2vaxjA7BgrsRVmvg/GmVvvxNJKUSTsqhkrMf
AHc+uTS7dVIeYOwTJSRHBuJfL9PaVQAZckGDikoJ8XV65/lBcsqSKyafrxRWYspPXT0vwVASnVcm
UJ3KUQJykhZZEVdrcgAhyQjz3hcnlLIz9O5f0QCyM7Bmh8ohV63QpqrZUo+9HSDI9ehrdBsIlIr7
oxScbfGflnaX0+broYDpvHBKiwx7i66UWuQK1WbG3FOgMGCcamWLaEvnF+XbowMbkeWVA6O6bxw/
bqMp8uERspxCWodOmcARWDUT0YV+AUWQOTGv655BTuNDb4/P7ExmlTKXxVYLGqQC7bMonG5QgBAg
oBbRpCMfcOqWyjtH3vn5UjMZZLEUMeQhIUlMv2PPS4+9S2XP4FNHSJxQPps9W2MeZI4daNM6Wu/J
ZskJFD9KrjzYp4XRfSy5MecBOqJ/aOE7wM4XiRlX9/7xFO9vZh2mBkxVxgLTkRJFt0rvT7h0EaI7
/tUUcJ3GuFi5ogxD/UusxkqZmQ1EoXgD0DG/d30iaq+1pTGmljdMqi+ttLMYNHo/sigpw9aeMILJ
OVaj8MrO1uXNG15XUh3XIUnJaiOb/Iqtsn/SgBFHjb6vmfYAgNSynMHukH806PtIEepWKgpWJeKL
aKSwJMriRouBSGBNsMZ5iJHRPw9//2+ydMcxsIRq760ZqxoXiIfZKq8S6eWTDktYB0Ugoqav/9LJ
VhF76QRwDWu4iHOU66lLs2wkDkUIRVfZF1Hy1/bd08ewSGfE0Bpy+0hHZRMtuPFP/ULYYQR1igm2
md6wdF4D+nV4aAbHVA2jJsK0Vc7wYrX0rr2x4e1ofsOExmZDWwNO0/hZtliC4LZCp6w/foUIUBpj
RrTuJz6ptqEi/6bOz9mDsAivFiUFvd7dUEAk9usw1DV+z+dnfCymOwnY+RIPr2XXT8CageKtu4q9
4t9CgeRjM+h+jBzCCqOZlLFFXPPfVbdStV87PHB2Kma/7a743Bvps6pxVTwUIQp/9gMdLe5qqFz3
XjE59JtZ14dPqNcQheKRg4aXdWxHfzknaf/ya1lS8PdlgBUF0sr96ew/zvt0GBDeJu1cC+MyFtQq
c5a4Nx64GFob28RuarckNrzT6te+OJQXZgddQ2FVyfJDqNPP2qMdB7T4uLuA3d0CFw3sJc8eQnZx
NirZf9m0WcR/nG84z+QMmlLhSMDwge9bFByUtKxhXitNmcyasLZ7NWK/+7vs5BvHsbDuPMxuW0Jl
XR5lF7Ia/PKH5A0+WIjs1oRTLhBrn71DCFRl5yGQlT6djblaDQ80GSEBZkzC4qPrz1QSNPEv0zKk
bf7NiUDa2C9pOi6Sdr489gPbScxcc6yPE2LxMQGknXJBOZIyaFB68JUe5A9E2EYKFOxjJVJE+oGW
7sDvNlafa2Jkj46iXZRzNwnYgvCGDiRr+9kYuhuhsTXnR/THF9225JcpkCguTSzuHQaACxXerH5e
hZusUyiTBfbN2R0yRNokAB1NwzKnqz7gUML6tRZdyLUYHxKIT8r0UpcXZIfgy0u87SQaRtUM+5bA
JhDB/8cCvLWX2OQfULApQda23UW7RqPTuT6z9DN3GIOIL5CSVblvF5QbkH4Kpc8FZAR6h2ERFC4V
Qe/Vz3MqWpgdBBy/0suaFj2m6QBg7d7ShzmGqFtnz0s8PJ1NiXPTA3y2J6lkP6k4d+wbo0TIN+3O
9Ke/HZnA5+dk/553MezQGdYFJWO6LD+ZVEnA0CYBCtURTw7755hapnxdM40KLIC+JFWzsP5Yzxtj
zOgN9DZUghhzIvgkN/0Bf3l4VVchbz5CSD9w1RVKGEY1Uxkk58BP2wptUxNtepU5FfY78CXnG6Q5
B6W3jwvt1N7r/XJfj1bZwWupbk8Dgb3uthQf1BIoIW9BxGI1mJFokFjZIJED6wA+FeyYVC0jpbXF
fz7r2FjEA1xMRxtGZycrMcJ2x90cLdka2BduoyJeheM8nf/6EovDiR8vbhzg0IDjLt2gIhkAWpZv
6RVIZy/RBZTIJNSVT+6y8vUBOqUmm3mZzEmyrWILncYMIO41w7GqFHvc8NKy1SKTudmC9UtobB52
A8zgvsXQgc6DvoZHW5ndPxgdr1XR44WvSXmp5+dVSJc2TYUEIQdBl2gkOFmpuoqacRCiKuJfXES8
DXGK+axtzT8LNzqtZ9nFtQSQAo8Z6Ce23fjYxhBPTX2Y/DEVIOiwYBLbODyhbkIdp2HgbeZGpGd3
L5SrFLV2U45UKbAuWyLNhXZVS/WnIXC02Gvu1kgveXOL3b+SBB82iRr9G8XdhfxA/7/ZUDbwT5cS
IZztLz2K3gRzQAJ3E1E6ElOr14vsceS1O/cEX9Df47oO8N7KQUTZQA9oRTRsPJc9gvcyUIhQVeqW
salA0d8tDefMnbQRkk4CJ9s750e2TJI8Jsows6aJNlILTQ4k4UquvvY0s1DmpEnY1CmxaSvukdqT
PFUe/yM18NHJ3nJZi72WFFbjeFiRmNruS/0PmKVCRHWkS+aw3tf0zsv1jgOFQQYPG9cHL9zxyV5a
6oyRlFPzaO//wUwjT7fvK4a4Jq/hp8WIhtQo3VLOOFsoUPdeta6e3tpJn8QObHrlbu4DUPdMp4DQ
8LPD+bH5/UmSDS+83xmAWIRoXmt5j87pu/TX8McMWDmTB3M/O8QUTB2VdxO/jUJB6UdX2EoRWzWR
XsCtwjBBOMuur0PTvF8hLSY2ppqs3sXnB8wUUvh5C8QwgtvZPlT3hv/q6jvJnEskoxT592Vdlcj6
ykPAmG0PNe0TH7MJFGwpx7qnxAGr0FkUd0EGtAozat2+AMgM6PhitQ7YtjORmVVHgV0vdvQxOBzg
vIge7Am+PBFg+rN0TzgOMe00k8je4Z4A4bKEFVN5fSNB+Nj5GUj5W6HJile+6+ruGDyKKrZLDzGO
lfHGWVAv3vOWS5rqdP3sUC41C5W67pXaJrsid7FwWVBKPQe8TDnmRGPUM9DFh/fIRGWWGlcOMft3
VPNsgLninx+m1Kr5ZgiwB3V9KV/ErGTp4xssKhvvJm4YI4xsrBwX3h1pt6N+gPv58sjjMmefpvTM
u6l/FKVI28YeDPZcRt/md8+8TvbywTZ+KDBevIEy/SSiKOxjz8pokIErz4B/vqg2JQG0pys7iJj9
SJLw7sfnvktY90EA2NLWqPhCWIZeyBzzaSSF/VEyjqnZXjLIBYutkNeBp3hj5CQ0xC8WClqSRNru
ZymYDLZTrry5ZgiP0LA8BbNXoTndcPaA2MX/+sW9YqZpbYRSM6so7Ko42fQRayFeXcaf+xv4bUaT
vfukjbZAzlF/QBj48qdlao2xdLgVSo1p8EHgmmeVdE24CzMw+LONBjVpzy9RQledec0weuOPKMVr
Gu0wHzlvV9kIJjUAdOYRKmPln4/84Yp+mqa22B+2zS6RmImrPdA67zzFpMqlfTj31nXGTxuGoc9+
19Xc3X0sYxj3aTPseeMIfePNu7Dbi8+fd3g8ZgdQpv/Wivko9bl7qc9ygWzv1PQ9IGILrpSVhG/J
Dth0vx76i1sPtmiLN0V02CdwPDa9JoXe+NWwFi0yi1sgU6GeGTrcRoqoJ4WSh3XqJ7wK0NQtfPMu
xv0m3EtvG8UGHYWdHcBpXv4St03V6ztuZ2m4NtTebTEnQs5wEGeAb9adQtgTj1DkQLc98+XqVlxs
QO2nkTZiTwwEjSJVWt9bnj2Urdia11zxO1yJ31w1Wo9vQCTtTEqNOloIPCEyZkya6+tmrPHD0exh
qW63p6wKW1xdDAyT/o3KTuyoIUu0NFgJKGkDwjG2FuRv6G2AT5MhyMbAUlwnp4JR6mPDni8DjeDU
YAhIlKjpKcLwWXMs5iQuszp7TWjc8t+HmnimKdY7js6Dm06DQ8n6fOayu4u1Yh2eJRE3OF1GMNZs
7l5v8tOgAzuF4JQFCQe2QUERipJpCjWLQTKHf7AFgB17bwds4WLoPavwicRwO5/BH/Qx2zE5oxCP
YpFk8cmkUDhrQVZb65BjTtEzQVy4dNGq9zkjdSVO0lqaTx8pu9E9MKXGJRrziVx7cpKq0aQrzYQV
GIWyzeGxbk2qHSKreX60hJXasxdAxgN9FQ3NYzPdHeWo5R8RVymn4UOmz5A2bpcI0BWiTJtf/Rv7
OdX6xbH96qKCccToZBC7xmyyN7C1SuxiSaby4EktjoXKn+lLQUtm0PCBxIbJT86l8xCds9wTwNy3
FmIXRcGGVFAk14ejnHl+02n679c0P7fT9dZqMf5cXd7SvN0e2zuhEAhWoKD60WYfTC+XqXoB/G4v
JlRH58Uqp/qCOHyjtz948idBtzdR8f6UQD2OZnbKYpcM6fKwYJwEyq1wIcmnZw5bKlimjywMeUhj
wesxGrrAOwRxGsPNuFCUr4FoUufnGKSHy4ai5G7EtdaySo3DsX2Gqswa6GQ8xfGsuA8tFGeMvxKY
wf9oNQUHvssQPd0t+SHBa7PheyzqtfRk4gXpMJIDQfhKmRj0sJVwl6iesCh7ri5stmT8ObA1hNB8
dgSRnOBie4Y9JWhkdNzcpALP86Ebfc9rrOODpaghwkaPD1fWbvA2DE/wp9etgRcT5NrLH5zkoyZM
+chZJ5SjPEuKnL8kGtBi54ElzK4SuzcNg2649zq6u9BMMMAAvzWclshrk3pu2YLM2exTY7Lzy+3Z
/nShYkye8De/JdMRls6rbm0yBmBfCBGcg2oHwPIv4F4NtDOeZSKBYfyHIZ58I9gm7i1NsI6f4xOa
PsFqEdYFc7YPOLfKcIJtJp52xmaHgOGfadyROWu4jIYyoBdo/2ZcCbJmnJBKHQhTUNCPxb130qmS
ByaKrpB8/neFF9wIxTcy9hNRaG8HuLr3KpoUrGrPFMejSSRsnOP4DV69sgprjNmcss7/d6QBUxcX
5Ta5ybdSrWrV375p50CFSb+JxUjGBTQqP3NSVysI2vj/W5GWAYg86hEkKDPRLwAOSbo2i59q7SAV
94OgP2ZvoxGaCb6N/rWyNPIfnr0yflnxpQGopF+QqzpjceAcSmIHNwCU3/vJ4+QwIDzJh8AD6mqg
EMRfoFnBT5CDfo2Dv9uT+hQADoM0t3OLEfhypdW4whlvxHcazeKZ1Yn0pLGINjySFcs07qBr7LFU
ppxDRRtBtcC+XCRjIG4FCIzeJ2VozDAESi8XqpY9yrojlVlwNj1Ok6wZKVAfvJ0O6TXrvvrgW0hW
Sj3NJtUCu1UCkBCQD0lT3tWoeFK/8NBb0khCt1z4bp6j/UYLHNDQailzjJdGOAqSpUvP9Slba/Ke
r2RmKRLjn6M1Miq6Dp90iqKyJkFZYJqtwSlpRP/5KcBn1NmVztYoCeVZ7yz9JZebVPc+oHlXWIVJ
8wiWcoHGXIxSGvygjlut1aDeYu5I7UNCuQf3Eybb+TDyREo+UziNelhj2THMwdOojNPR9dSRwwWu
gtNjcdNlDWlDARHiYNRviveEHVRgoiA6y6CmOlIixrm6aMI4nuxsLfclycDsadI3l986fliSvcX2
dfufTD+EJQXeKn4PKovMm4YK6tTsVuGDB3wymt442R52tPClTL6HPDf1pkepyt0q2mOBMhYNpY9j
YKNDD29bYBTKaYokr+6QjakjYGMxFHlazyXbGd6wMGBfR64SGhVK10Vq7LSGzYfHSpLL1oMEd5WX
3LiylEb2D7uprzB9RE4ltsnXp+/GVdfokucx4UDYPPgOTsMnfiwIKZJW1VLH5Id/ibwkz3SRaoIf
nQyBu4HSG1xvRzZ4TUJwEVI50NQMtFU5iduPImlupzMOuI+PiLMbNYhuaZZW8SuiVANyngVDj3Ft
/I799Bp3LhjleG6Z8Rn4u+g/btKwiKLSja2sk6qpqHCL2Lyuzc4GgdqVa3ZWKmbpVYvlGfAueEUJ
HLdXXbtSGLJ6XAoNEGrTidYUYSx69F4aahW5kvK7x/ZVYmrbmqAh6FYmZZr8/N7D1qGe/2kPFoHJ
Fp6qB5aYTEnMIq4piqzljSobimepC/Usq+aPyw2vP9hmDpy56x6B/DlYUWq7eCSX0MXz5qhafYYq
bDFzAF17DN0VuCD37A3Yd02bsLhxOeLhr1liYE1tBVH7CLzZtun+AirEcgqe8BydSDUt1/Q71CyK
t1rtPwiJ1diEy6c+FaQMy8jTmBBPf8aAermDVKRyAz6RIVAI2vFUdZCt4A823dGBRDk/iygjBUXY
3pm3mpqknJ7eDyG9Rqwr7o23QKqP290VzVtdiuONRNENBibYDR3vmWEE0RWv3kJ/er6qippVdtpC
xYPQ1SnZ9X4xU98slY04D0Pz5Vfty5xpSf5F5MZtqvfZSm3hZJKgrCM0sjW+GEZWOhIiWFKEB2g4
D1gi0S3+D8W5kEi52Fv2DaQ2w1eTSVg4E7rC7X+BTtB4mx9JpUyo6jNfSZIJIAg8q1xC0Kg/9jeb
g1pfI9xKh/C/ykiPbN6qkNS0aHsnIC7+wWqMrmKaWDbJrjXRlrdtoLAV/vQeKLHo+RBnM8UYtxDU
UulJh7tk1ms4G1SStExFlouGU46F68wIEIEkWs0NhFxSujcgiC/JfWqlB2W6aPCqO1h8PCuA5clF
4cs9lsgYjQBr1STJ19pm5QrZsB0d2f3TmEnyA8HrLCjUApmJNR7UzvLFTJZIZRM8HwVb4RcWde9H
+22POTxq5JN+ruAmwYbRf3Zlkva7Apn4YkZaWSz6sguQzjkWgOdTcb/ZsVfQG+JJVYiYKjrttrqk
jcpFqFcnChv2uuhZPv0YBlo+riE8RXbShmoS/Q12qfBAnK4jmjX+fRzceGo8INZO9aWPzavnNmke
fFBnN22Pa1MweEKm57fKrY55ygqh2guu3QhLGcrXpIFOeSoP3ZGrSuZ7B9GlB7xSYfeBNeby9L8U
1Hn0XtKoNfZfa9iuUU8Kpyn2uOvhSZqFvA94pcapnoCtRzPt6G61ou59MKIvr15NCg8tSzPW/ZWO
N5+RfnJYRT06qtzdCiCB1xbdeHGp0FDNGQBRVnVojYTEXzeukF+mD51UEvjJn8p0k/El5HShriWf
R4PFiEQ4ai/17vJSCPDPu4tISvPPzHOUYjiuZvf+Hi7QGWtpw8agxkbF5PEPJokqTAR9tBJmzqa8
ZmARtAoPz2Y2oXE58kpsVo1XSUjdxeKHhctdzFtYf+tmzrVIBdGgFVyFfkeJkcaFTkLeBulJsEgv
7CqgSFaTzJQZRLxQEdebpfxbvAYag2u8ZGNXpNaoYe5oyKCLH+tEe5RgRSshoO6XRK/mOivEzEZd
1YK4nh+qGZ5SaQsjMGrA1G0tqMF4zodaVHdgK90lnCeLh9nl2p3jtFFCsOsh4aPFrQ2C6hXN5loe
AUGbCEgT6orzwGrIYEE1jB45f/r0hBffjAHW+I82/q5BGZq7WvLUlFwDdSdM81x9A359rg6wfKU5
gpZda+KLuVNhJDl39+D8qECmAZ44IHMxbhDq1dlw5pgXraL6YyeLFB1ZI03xsD3VMgoAXr2sqmPI
xI9ZKsESXWnPNrUHwPTa/CsqYu8ddXo5QlZIetaYEq7dDazZTQSqLV8hSLKGHx13BflPBNg1cAUX
VXL9HzR9yVxgdg7pVv+w6hFMWBNVdqKDDM3bStZ2Osbwg8OU/aUcSW6mpfxRskDqzwT5Ds/tZluD
+kF/Q3uSmFKe6XB3vK9KcBNafNSSB8519dRseZeAmZ9PEiTmTuqdypzavFZTOPZMHHvkeP8pxPj1
AvB4uVp4K6O4hLA2KAlETx6CLAA7jCMvgZgJGthf7LUJIm3aVbqEZ77//N04N1M8NWu6j/x1hKVE
pvqxcGTaRXPqACNVhJLtyoKc8gkzTh3iR6QyVRwZf/N8b/a0EGIxT1MmQLskI+8MFLf2wMkzF7mP
AzRLCrME21CxEQm3jOCrJYJiGqZE0iZLmh8zGPa3SH8sSfKdfnEIkBTznFZpQSglTKoLUzeSuvwY
737045+U2jMhkI/soBcFtsQwJY3AMSs3jy1fBo3L2vKQw4lcxgl9Xov1uQcOTzFc2dy3lUd+FzWY
Wn0oEmw+QyTOyGBxDGDss9wubPPyJZR4ahPrp2P4W43Uj8iTTxM6LnYu5cQgTJ5+UAK7vPjyyvob
p08hfauRAmtYQPIkgVFm6fiax0SK+ooxKk682+3hfX3pubPkMhrq3Bn6vKYvCNyRNA/YqDN+M0vu
ku1eu15N59CZZ1N1vnrqAtPU6ZNfas2LqA3/UHdgqbwSb5Fjk+Ysr7CxZdhrNjKHVJK1b3OhxYi0
WGrvmOVXPSoNSGPaugxDlVLt13GRwexOEuzG2Dd64LMalqJy2/m1Ib63pWAbfxUbsenKOB9XAxg/
TCy0GIVyeGDEgs+tnoJvqkeBj3OphhMcV3pwD7HQRu20/CDl6EKJfh2eizgvHMS7mrZfInPyoJOU
g+Rxv3YxIrP6RFErXYPYXvUAYWvUIf4Qfkz4kXwhr/dnx+Z0OElfVewjnrTs+gOpIJk6xMq/nE19
vWWXgaPopkR+ViqVQsiBP5yOS909A2HcVK8K/THC8YYzjeU3YAyS3Cl+sJIRZHgEqFq8wMvYrwpq
e62YUpPjGbENnZEhhajVy2+4yGpOcsEmBsTzqMai9+J8xAkmHZksaZd7y+G3DOc1/CLndKEworqp
y+Ec1hVLtaMSr7YRkGrsG+MjZ/6rku7kWp+ScRiN3YdkeSVNa7Dzr7H5SzajZvrYHWHoXRNrnXJt
gRaWdrxu0QrJilpoNqELvyEo7gCMtpMpe0Rc5S8yhPrigKBD7JTaXGWOn9HRY3FZVDxRaxh1JdU2
qtXpLn2JO+GBSsKj6umP22Qzr58c4OAWaw8Y3DrazI2hLt7Bosct8583C6rFmMJQj8LmZT5IbEku
5b7Z3sFwHrAPCCmLUF0X/WugQIYF0CGAKf0BZHE4XKcYNHuI9X0La+0ust/Gi10eqIG0/YJjlvKD
kt64AKmiVXv5kQyLO4IFRCM+chbFRE0ZHAoabdCw6mJOKfmPDTKjKmYCBDlgU9Z/q5MhWNVzTUg0
ER7wCt/8ZkszOkxP9MD6GiVotKaV7H+YExGkXGcKgpN7Hv8zDc7h4hksM7+u1K9yayozda0+DESy
WFO4wmRXZHKNeuoK9KtogmnDkiP/LG7rBX89FoSL1AlMgDbIZHdloHXpwrxX9cbNvjV/uLQ+jIfF
Jq3ArxCmGc/7WkNqtVol0I3bUhznEr+EkiIY3oVOtF3X6H1yxcNXFfXR4scrrWmEyLo047ULqtIM
+Y1OXeVmHZyie3f5Aj4XhijFrkjHTmEnrnvVSJtZa6xp1XLgmQ+WFBlUL/AtkLcI5aEJsPhhk3sl
2mgOSWLHXQ9s8QcjDBJQOEy8lrTFCbYCDmlt0jRNjDXl4nGlnVazjBFcgD8J1g7kq+JyZrOGtE5F
FpKUnWSkmh4b/Xd7ePURWhX0FIOYJN+I4PEXw5GTGZmu7ZrKtTC4n/HPQ1KESWC+/NUWlUYY+U/Q
d59nhzbMEdICW8SNfYN6ShshGZYUTBbsqYfrvUX7Wz1yfZRKTQ+0E9TQTlmqcnxYdzvc/AZc8kjI
toYXPbOWPVwOkJMVjNPp7nlVHq8uCoDYR6ZDUL5nw0YJKK1M49war8JmAYC9Mx4/ovqs7i4UGswb
fZXfuHTRpfD9t5Iqfi1czZDo75CtWylZipM9r3q7cX5qg7nnk3/neAWEbrfzaFhwfCeXQcRCP0HO
/ckI02MzfRjoRwH945LaH7OZ2cOvETmmoJT2b2nFf+BloSq8cCk36t9KBwEVr8cbJRCUeJrKDqf3
vHP5/aVSjD34DSiX89nfpYyf4xmmttjQz2y3pWbcL50XF8JyViD8IIkE/g+DmUSMo7bVZnpR3xP4
3o81TUooYsaJiwirsEQNdXhi5ANwLC3i9jli7qhl2Yace9ajElkgvD2hMKVLVWGytdQ0xJFNylsj
SIiL+Vzq57AjbPN1HjkEA74wBXYg7mJ1BFziOAi8q9gm9Y8KOi7kiEkHdGzZsgdL+3FKBxW+LuME
FD/KVDs7rclcI80wjE9ne4Dznby70pJV6cDRI8g3l1ZQmMT+0i19cMAK/z4Z96KgS/Ok8p6qOH9M
LnoKUDCovwmDPnojt2xBn12XUQUBwLbJ45DOS66r8KCXIUg5pQkznMUf/zZ97856pVHsXz8jpEd4
WBg5uux67+iTFcSEfmVqzk1F8oF5KTeTj+u0TZ46vq5eKMCHbSFyNoLj83O91CLlOXeNZ2ksLJvh
w2ICWIQDPvQe5NV6rbHn7WFmRmCVF3zxlxHGWuN3QLsxnR2oeVqmAs4hEK1/XH/J+2HUgDCp852D
5BqCy/+RaA5Z0QkLfsTRKnQSYcGAtYPQJw37ypWw5xS/2z0ODIITrkGcDo/xqoyccHHodzgtZjhu
TN7a6NpshJBEHadDMs2BsgHhcKha3M3ya1yUMPuI6JVx5aI2vjRyBOa4JtZzIRlKn56TaXjjV+GF
WjMlj6TNfbKVKisz9gp6E2KogS1AL4sXE4j6EkD4NRIHf9D5477E0nqSZGexQqzi/3Hyw+0H6xsR
m1da7a1VsO1yEZ2m+AU15MAvVTD9c6h9K1dK2vRZwhM8TkZBIO5pief9Czm8kS2QnHhNFvo95Ue5
Z2Nqc6TE9/qtfinBu3hfkWGeKA3c2cBsqgq3XkVnBY5OE1T9fmD/8apVAvpXYQSzAcms7mXCwaw1
i+/GXNQ+/A0uP7Y6//YSYhRV0n2muWk3NYs8Atd0ShseRPXwF0mUDGwuPY/9m104Ei2kvkYApLsN
DwNXnX8PxUyFka2rum0TKNHxOMrGiJohCtdBAR5D3OpLfQQpCcHYFoGZIyKG69/mojkIrS7aSd1M
a0Ke2fhP9r1wq7ELV0n3jvilWIy79V+A/GppAz+MJSf13JGV/NJFCtp01o9q9gqcOlLn0IKqMjdr
YUcUG3qZZkrbzdGU3UBCyrrKxi8J+BS34+1KTMtkZs/spawKquJ/wR7wBJ1ff0ggKcQXi8b5pLVr
eWgWgZJAd3K/xO7FEoUg8LpTW0Zvw2yCKsj/KUpDxGCp/oPVJ++ye8rFBy5n0VpwJQ/yBfyhqBTl
8KcvtZrHSXJiG23qJQDl1d7lNAybcWs3k/PyQ3r/cJ7CiDWrRDG9KjDJKjMuFB4iQ5SDTxcun+m7
0hPxICDukvcXfTr8ms+YU3zx7VtUo4d90BLPhyOPJI/UkZpqXcsuS0nBOTogzq56kpxlkJ4Do1tK
lLxqyaDOBpP4RvyIoWl72jSRrydYJrk7stejV/tj5fxHPh6Nyus5VbxBntZSjYblIMLrO63YkGh3
AqY2PkjjcsgtJgpwxWMegjrEg4B/60mc+u4v83mNbkdPJI4kq7Xd8RVYDCSxJ8HQN9tIeAKh0aMH
ixgi/fDC+kgEQvf+iyZsvhvS3LhuTVsTOKp3hXKbwVMo03szKBOFDk8Ji90QTA/jK2w0osWjs0u/
s0yUl5fOevCAANw8gg7d08ACs3YbNgkkaoIcnEETrlhkbSm/XVj5O5WXU9gQ8Y9sHXGSOQSX40dC
jczq/zhiBhLjnDQ+0aFYz4Ts0rp21A/Pa49ADLRRB5Aw0ox4K9hyzMDplTekt+SByDKaEjfEWjj5
hcjbDLoc3EtvcD5fh2uKfnWrjBEUu1D2YTugscl6euwZjhGLMVXSvIpYwdnvIAxHgDD1hP+D7cST
I3Oak4MC4H+8xeq+PKtsUrXoKAjN0OyJc6vR5s6OxZBp7gP1FjnDVhkr/4KccbEZgkfyjNj970TA
mi7rSiugKnvjL2S7EFF9Jblt+joGyuvWPBUvpxtUAr50R0sfdg6HBHQx5pMpufOHgb5rb81wEqEZ
HDEXVc6ZY287NThiLV4xjycBdZkuhjMLqXbqQoFStl/1OYAEXKnUQH2gR2xlOqnJot9eIthtovyO
h8tJNOtHsI21FVmbUDEpWddAP6KWaOeU6Q28qJ7MyTWKM7U3V3yAFnLgwtqvxV+fSksbf26EuUE8
NN6r24/iTD+E2tQwPo3FXuAXR7lRtl96ny1GBQAjSQxD56tx8PEKg+/ZL74Xr7FhEO1x4mO2jauB
eRMqs09vOlrGF/MYYgykkl7VxX4lpgYlJUetrJpMxOqgGNfMBW/tOjUdUlge6IN2ZxQ/mty386j1
9ARFsCtQLuB34UaHvhmCTdqvWER4TeOcrX5hcQmZhidxuA8Bze2/2XBBL2KDwNMpDyfy4+Gg+pFO
vsOgr+5zfnSiso1uCK+06K8ivfxyIMP5xsBH8fx8eq1VNG7dLn4L++KpPUQQNidGtcFWDux5PWle
zZAzl1mrF7eEpL1Nc1ngbjlkRN6IxzX+SZ1ETuK+9+WD/By95ZSak8evhYtiQ4CKpBwa4D8DcZLW
eUZ6aprmdjhL1daDU5umMFURzcKqJVGTaxOYYbnctR1Er0KVyPsMO31g2MOqGCTbpjOndD+UPwo5
IKAfcGyW+6Fr7z90dEnI4CDPmQUaFFrNRWLWcnM9GvBXWiqX9SZQTZvnvJdCAF/5KkwhYLu+aGfD
N9M9f4aAZe+km+PyEZVsp0EiX2LmdCQ3bZHemgO121y3Meek2pxcErvR+U9I4Oum8F/vxVyS7Kq6
A25v2soQEIpTCwaRfC46wzmCkVuP86x5/PLy0JQ1d0aGYpSneXsKOJkEAtokEhjiZFXMw6xz4DX+
cJSTSN00KxQdd8BUT5epdDriQm01QWcyg7hMAX6SjEJfKntSspHePWEE032mLo52vxsrsGMBmQrm
4oFWyCwqNsAL4CjFUJ0i4R7gzCabR7tHb6830EdcHu9od1aKbwJhJ0Fi7Y4V1eL0ZqXQhIRQKzoK
qeR3zc8qA9YlS14Vg2x1WUDC0LZKHJKgOOv6zGFFRQ9G1NiFHZvO5LKXKD19gioktsbqSTrZ72yy
pPP0bkhqhOP2bBtmWh2KlzQczS8ho8ce2UiPJOhsSeIbyYeDKKj6wZMY70HIKxSoRP/61ujnbXNB
tMrlDhVjerRvCH75txP576wM7XcxZC/R0yVluvtqYjMnzF5Mmw2Zrv4E439L08Ev9v9rXmW1CucX
HJ+p6qnQFzqg7l+5zjz5nnoaazz+6ugFaqdbao3qN3RPYVmCgVR4+sgEz+Zri5I65mYIkeV+fOxr
GAxnPW12ob6d3lExZiX0/dRfP7RAf5QNGQwliqU3M73b0AWmQr0noXyzjsi81iKqtlHEymdMHnf/
Gaw5jI/tzmHsi3lCVgpjVLRf0P67IW1RZik2fNTiRCe2rsg+OnYGKu2x0rrkGcAJIjlMjSY5nquf
KKpZ/hehmxZ4P5JfOvV1Pd7bl/ML7nFFMrSKSD/pEfPFUjOh1tYeCtralkzAq6e8unhMLTcpw7bs
gUOAWVDWojsmlK+ZBT/d1vIoLxlng83WED3lpVemRBpsmOdq2XAR+/BaCCll8g5roZOZG9w+H8ev
ipczene1e4LcuU9zNE5ZEnAV5Mp9ur1Be8VU8WxTnRMJPkao3ao4AMWMH71jE2MFdWYMj1rCyFZo
ccGYAChq8yOLeyja2JqSi9Phax8+Dbp8WFuLqSIDAC2TulTR1A/1vHztbI9GftxQa9rdkKIgwjZa
yi7KrQ6m+HWMEF20VjhoosQwh/sjpAqRwi6w46ix2OVGPYQp0uZp2vBnf1OGCirSsDo13zDKdGbW
ICOCa6F3+2GKFRq2uooTmaAtCV9tYNDAMeeesda7qe3a65r1yFnWVDoSLpA4LrZMcqNIifoYfMrr
CyZ3Yu/Am046hlPdRRlKrkbl9lel2Kh40YhqqhPBV/rqijg/dygBzrHsR5HLjv/Hg8ao5GTiMfjF
wRKkf7IVTxqxaWpizaSiZyGnU8Ydw+Sw6wsrUVyI3wn8ea1qmCgHX9SV+JU1iMPY19xLdTxK+FFt
DGQShRc9huvV03nhTliqTx0N9Y3QlgAZIjLYTzBWjWYLc9htOaCZxxshGcsTZVqStFcNx4okLXfy
dIHHUvKeEcxuGHaDi/zH0agbbQ/3hJN35Ldi+hj9vs7ZUjQc7Dhu2SENEqLeMJeIDDANJx3EH2F7
nzWQloWkkWDtE/8Ht2lUOctc72Ce6PQ4hJ2dKSABFx5AFyCVm9UoDzXcmVncU1mkaenR80Wv/vEy
qtOBqv5kfmpIZLzY3ACI9dzyeugqZH5SZYQRKSvl78dhM7lc+sL3EMPA28DnfW/fSbWR3byMS7dl
TGBP+UoTCeLq6I5MR0lPErjUSJCQh9sJuPLHCmfRgpRt7SfcQIgu+wHQDUpAr59qi8p+M/EWu6gR
v1p+juuOA8xgUVaxyLgqH1Pjg3dWSUchwxcDAgkvEl3kdom0E8ie2CriftZU8CSCojcsX44KD9Sb
jLv9IiK0kYiJhAIKl67Ku/ZH+AXO197cD7dj+KdEb5V0gn6jExgLPUB7ZmwJwwIKcuMGQvrM59Gs
7VStofOjM0UXwCAEFBJ3ZvhAssptvyEIvO+28Kha2vI4w/n/QEafHuar97rjKYDyBs0gbMNSoxDe
Ah/7ZhvKZ6D3JhdOrdOuabkEeBL6l4LcNIl15hIXaKSBkUAD+ztmUxmf2cwQGUVPyJtBJe8Mf2+5
Aqws+UYrP7UN8wObLw9OV7MJYmu4GCk/2PIgsd5sonsQvei8PEzIy3THNPlZgsC7g9VGxIx3yTjT
7YmByG/NxJ2EDN++DXHN6Na1ktzsHQc3w79QtGvIYrrup5QEwb3tWFVALIzqNIVZCdD3EXwGWyDX
ZeaSqmHY2af7lFXhdk2+0kRTVPVHkgCpuD+h1Y6tMXwQcnphPQ1tmI3IrjRT5icTj3d3Tmmr2S3B
So6Jq+zaXkEvA3WfKWkvNFPc/eH9JnLpi5UaA7AturnDRFbb9Se2cV9E/0z5SxkCd6iCXJ12yM1G
31lts7tMCQVYHLJ+tBgpdEWGIADXVg/uMQ9mq7LqMP1DtqYQj0Y+V4xIg96rInRgPLvfN6lxeNeO
xbrBQMM7clBqn6erBQaUMo9YWdRXs3pjrmVLpxSGA78PZiEfDRlaEz0XNTkpGRQrx2rWNWuZcPCA
RJ/0ztYEuEGbw6nG14bQRa2AkMbkaym9G6Qtg57C0G7q9pioT17z0EAtTtAVwQHhMpSRb0eWnH8s
BmN6FaHVVJE2rqbpw7sYQPT5FFPSdTSyS9EmcNGAslT1BvPi+VIy3OeHg0EK8Xg3yPN4MzCIBkyK
N0QepS+Y6fvw4GM/2xi9eIU2yRmOCTcVc6xX83Xe666pEBpWsHKuulJR30E7NSHmhHwGbiP6iAh0
DiurMm8pFGZ+2bn22V9k8qSpHbFb/eBZXEUpxCmmgxMotSkQuikufndz2PXyN4ze+6SvFzeS9ItU
75lhfEDP5m2o5ZxrWkoLPyue6UWum+Q6x0SytNEyxHrKAbwCXWgRC6dyJcG9zEqgi6+esX/5LzSP
6GQmycGOjkEXq7QJbmanOr3pmGDYevboyTt5f5FgtUeSJkw1S/I32j4AIlAlunCLJnVWrvjXFrNY
yltlYtGvapVnSyjRwKNSbiW8fRJ7J8OTWo3o61HbWUlM84q7/MsgIZN6gP62fSELfUnxapAaTZiH
JCHL0q63b9dZeysyhkIfnQ4IvOygQJG8qcF4ZiM3cA1TlpzWdWiDnHDQ9UEgCgDo+GJ3t3KqAZv+
a0J5nucqjS8cy4qbkOcu7BQqCUPgcD5E1dDQE0WOuk2DmJffTx0DEJst1uf+j97KYU/ElLpbjdk1
cndum0yuZJ5+qurqAT/knOl2OTQFd4Nw5JLEp/DR/+cpRLlxXROwGxuiJRun4DwvwTqAck8W+moI
qLpQV+82T3no2Wi2cMechfiyq8V6Hc/I2LArHybjzFXdpJNQr5y/4kIPRkS3AOjGEtl7uRaSuVFW
TW0WTiMFoIcDv2qV7yikBMaSxP7aMCYmf9TBzVbVX+D8nbKb6RuvLgN2RUMj2PE32SBvhgMJKDp9
pQPqf21MOiWjFjFuy1WUydPasLWWde0OSL3zqaiEFuhkCUIs6tJgRsscYEVwZsEsR1v7vxez9U+2
o2cUn1AGfmhtCZtzLFvZRU13O737CkLLzDVC+Ie76JvXHbcbZRAA7fJs6hZ39bO68lMtAkh7qU5s
MruZZFbBLcO9T0Xdg5XCmM0MSX1khPX6IMb12yTY60gGSAH1rBRw6ORXvO49Rkyf4Xvpiy/04nfD
e181sDrHOzsvwctInPntQoFFhXxO1aBv4ZrZAm4Hi9ZNugo5rFSsXx95MffOo0JxE6lxczfHyyx0
u+mqQ7CByxKjjSFpSnI9pmQIU7Vt6vjfRMBJjRgiGlGiif5x/6SfKCGNJbfUlnVxhGsFByU9tzRF
ynHZXkja+YhhjScGaiw30GT3WWbUozidz0EAXH+UKZSFUVHWe2BFx8CCMV1Ldg3h/bm/gAMmCQwM
09n1o9ZzotvwRFtLVt9+6GpRqRGCaXwA3Aa7VgfL4Vp6iRets5/SSuZyxMMCRzSfis/GFcCdwEd/
manTsl6oIUi9Vt+NgsTRDPJSzjIsGxXhrHFhS0xGEv4iGx3eoBTwHflwk4Kw4sdc4+/3hUtMcdqm
ENYR1vAKRbMmBrqST7LQT2efaBc17NUh9ZzSj6SDNYdmCGqW3pPHFsHQh4snTqtaEygpvvz444jC
iKvTYSZlDK0ium+xhllc3QKi3KhF2qHI9fSRd8Phv+GjbitTqqNjle46NOnGHBKhTh4Ky0l19pVF
kBuyRxcODYbLJxHb9JNgFdKqKjOsxkfDYpfr2AAJAeHdkKyNTe253I6Crk99OUokEDFSaNE7TscX
Ju6lKVObIcP71T93Kp3Qkzd9xSbhjGiwcEiKwAkquFQYKlbUITL+c0sZF5e9YLW6adzDDok76sN2
9VpXo25f1zFdAZGL5Jd6RRfGGb8/7IZlQ0hEqoawMQajh7dvEGBV7zYAYLL+7Cdy/ve+IjC2HhuP
+G2L7RY6w9BzD/FApRboJ4Rqgo/xdfPwp/56tPWE2A7OtjEa1DcQUAnkXkEqGjbR0CFVuFFFmluJ
sOopBtfvd0Ya/EG9zsUOjSBLlmcw6tnhxlt3KGJMubmzriRXDh3QvQCOkrj51+ZRzREMMWXtWpEL
iWV8e9DgeRM+F23YGBdGpm76+MxbIjmzXAuCS0LGkmLi+ty6PlI3JLmWPrSApx0+thpHH1PBlgyq
tGEtJz6hKyuVLh4Qt2wJRPgib5qBC8D+SCVp0ag5Kp6SKUXxEBcpHP4GdUJsDWTp7COmlkEz8Xeo
Srq40UetR0prdRSF1fNzBUS1sTemVDIoMNh77MA4HuLNkuz1JJ0m+SjmWG9JCc5CD9AduAGjo72G
IZ5GD5KxkcT2qcW1qQkzoLOyQMWptr4n3QC2c5XkUzpgrmHlvcHP2oCn66oaSWtKl3ghKLOgxa+6
sXS5RTi3dx1IH4esHulO69pWGJnhn9O6RMC+/J04vahg+0LyY3KQX07uq2zExV30vzT0eev0SmBo
N2zuePncDHcE0U6lqMvrFfe9S1RM1aT0bTcgRH6b5VvSyfd5G92RIpiNwCgvnHmlq9jnoyVpOB1t
iUC44ETOcs3XOkzg697kqZfDdccBC5fmepUNHOtMAPUNw3bMlHd37jl5v/v85ykp4zGBXPk1qElq
n55dHN11TppMY5wFgpH76hc1jxiOzOUJnWvZBo0gkpfm/fsgDvO0tQtq3d09YXInmcMblizGJpBu
fKuFZoTJ3MVe1mkXZAX6CRo2pxwMLRB6OWUerBeb1bS5OWtGB9fFbTEjBogES2V64Pa3BzFqvpu5
wK4otVLK4vZFcH8cqJiZMjejKFcTFcvw3lYW99yU0oM4ihO8DJKgRXgxOCFjo9iVIRFph3V/Rxma
iL0XTOvKE70V5ekMJgG6LQHDvn7pbUMhI0qbvXp4bV8My7nuIBJz2iCexwblDhGGpQyxOfsWDxq1
6rUZt1tB6qdd0SnUbskmMSF/E4I8SequTlHTJ1ThpFm9SqxR1bqFsiGS0mGyuC1N7b13lwCPOlzW
LfQO4AcYAhUsH3SoScWALHmhKuE8oak7lpOpnByHajwZRkOTr0oApJ96GvMGIRL+OjvdCkyt3XUS
0aazZ77qAW+ygS63ij0KDjaih0Zvvtni2imtC1DP4RpKGEeHg/Wi+JseOsVGujX7f44OfJW/1Dz1
awLEAfRoNIhrkZ4awuSByJpcQ6YrvO+T1+GbAvMnfq4f61k12hZsR4MD7uKGGZ4EJC9598gxRR9z
8KtU8lT3f/8us4VXR9EzyIDxdbxE/FoL+kIYaSgKC4G+V6vAWva6LR1BZwB5NEPxssMIaIIFBvdN
dPF/odZCEM01z1aDKLKNb13E9u1H/MaBpm/yWhAQg/OFDyckK9Vy7G6Q4Al8mSHvlEP65T+RZe8b
HKmM83LIZrRgP8IDKauDFeZERQ6Q5L9UDMQs3WE34ytdrP0dKFFArD1/399VwJnLay4kmQ8Xkq57
n9pWTmoXHrSW1UKjqVfmhf4LXF54sM/PfkedEZNhKyxZgLl2GlLPesxcNAAa+slvN92WYwA0qSg7
YpzftAsWI39ZDNX+Oz+lDe9pTxjFacWYQ10176itU4/wHob67igOfkZXmh/YIT6OGtYMAHkTaxJ4
luhKJkBpIEgfM/d3CaRn84oCjgweib7UNGFtPvuSBFykaIXz0eduazeSD1ps4NC8sUk3Sbh/HCN3
W6HHjFi9aEUgWP56LBl0qswTnAf3GGloESiHeEkG0Dqyi2qq7+b/ERjALjTUigB+U+FqtZ698CUc
amZQKXeK32BtgYTSe34JRPf/VZS6oqptBRfXFbefrIDoBX6cGkjO+f1FMXHStRG/unton0RWRLHy
2eh89hbywq5BtO1tnYl4BOnMQJMbb3kafInmf7PaIciYJE89OFyzDq0amoBYYgQLV+8up5fKpKup
tDyWjPR26vhFN8BFl0TmBqM6GGOEK+yMqmh4jcsaHmUx0/xOE4PCzEKodfBtwzbG5iJMB1m3Bse5
PM9GDtJACQY02qEck0JCLyU9ubiIsi8sQHnAf5Y8Kd4xzviAS0Pm4ma5sj6//XvmeHXmCJoYiH8o
bYkGbSnY7bWI31EoAaxD1f+BnViqfye3A8EP+7QP0nidJad9qaxxgXTDkpTZHW46ExCUHLpvS3cA
S3HnnHP6CYHNuWDcZDF0Y5VrMZfPW+ldgcsARFzk0TmklfZcW2WVIq0zOJYpeJe1/otZh0K6O83I
T3o6sDdoEsdMEQLqduSGyqCIJ/7vdynE5lN7hAh2b3VvFQ5jhKiJpZGBblzi2r8ULcgcBs1ul/2b
9k8uxTzwfxJL4XC6Wc10JTFuvrvFfzkUik3C6GVOl4BUtgWxss4wjiqQYy8naFGaqvYZD0JIVCsP
Py4t/eKos1bX1HD+3QXPUN5tYuFiiZAF2futxx6T8nwQd86ZOddTFsUi6Db+2qYZ6LoMqSXkPWpL
wp/lnF0C4hp/WghKuO3///AupFp9IOW7BuXZZDu88IjOdel+t75r5I/z9C6kcxRu9gcjqg/zXriN
p7QEBFf7nCOOcBmRC7Dc7Bec/s20cDyZFsq4vNR2DkM1Ur4gQ/XDdUtHLTN1TfYA8s+iwZgjAmeq
KnZ1bgGKuKrwp8AmjhM7KhkDu9HAimSiHEJJSSDUNUODSRPsjrIQZHmbNTeTdMWmiwptrCwflUTx
coWAYZW4ZN6yO7mAqjcJtgxSJ5sRw9qeQMPMJX4Plbr0UZA5qvoMuZr17tGgC1opK8IQFMlX2i6h
0VN1qproIOqy3U487I66pLvnDRipa2Y2d+Itut9/FVMDEI3587GuOB6DOVC3gYJV2HZk02pGd+h/
1mWAtd63hrK3aoyrgaaVUzrpeHztPvBHwNEGQMq4Z5hQX6uS2vXchSK1QPXItQVuoPnatDFn/1YT
kJbgEmzT0saFpvf+1K0hmH+SoC08K2XkW5psiitLFRurgHxrDtkPeM04oYafE9lbSU+fgUhKyV51
lYGhKY3eCMr04RgCz+Neh8v1ORO+cOQii6+ZGY1dI7qM31/dCq7whAUjNP5V1KpiDa8lzbVBeDwj
B1AnfpmaMn+ocCLPnnIorZUG1kTtuo0p6/9U+dj4VGRblBcZU1TbZMUsOZMHP+S0QuR3CTRDpFiM
1xmJxR6LCdXP5fM8BjDbuAha1pSAMS2CZL0J6ehgp3IknLYgIRrslMWDMENHIf1U4JkmXlyNDY17
K8lBce3D6sUDmkRdFcmz5KNZAIE/MxciD7G0+SKs3uuA7KlCVNDvNWSYND2adjbQiblOe3VJvcfi
SsCeecdukpAv5EM4D4nScotd8o1rkEWBxrW/5uzVfT7Nf6r/teTBRWs93dP4/t27oM8LGQ/68EQC
yA1e/yf73ltFaySDfW0yMuImR1p4tioRvHaOTVUrw2aQHQhEN/WmWYLfapv2FrF/mJhaH1MHAuvy
PTWvnRGReF8CLpO2Z5ZrkXWnKVqCFHd3o/jPc2utJFT+1jIbVHJ8xnBAoWWEklcbYX3qDl7lw5Q7
RXloWUAY1BFWU3AeilylMvO/f+icvHaXsKI5GcWUlHd8L6/D4rGjjr6yzaaD11csGShW9ZYWRix3
75Tl4NbrLBTEbwxcpSUK+exj1QmaDdz10qmzhw/ltGaU8pNGKNu37DTToc7//FjuwkmAETUNDOus
1HaPEmhO6wRC+2P5IVzsdnXAOYYSpr/YF8d6lEZR2gHZA74Cos2d1x2j9Z2ORl8c5E4zrHzcMmgC
dAEUerXrjW1QAbDQG2HGyDi/zbakUdVgLZWbI2RqPgnbj9dZtGWPSaQmC35miyYvTLVMmrwQpBLe
aeS7ifwde7Ymat2TTKFAKMnanXvQ/4gxhJd0eO5pT03Q4SMD/JoOC+fEOvEkXhwxrclqyPVjUY7m
xvPoQPSkD6rPgAM06ZeiA5SvkgPjR3IdHFLCoTWh+HBX3SDogGrY9A+1F45IBY4CMuYcURlde/SA
E0HDJMjwZ5zP2YxZIzDCGYvaUmsSFRVf4HP6ZmSW+2qi6f2eFxm4UsSKA5y6EdMY6EBYIsd6skud
dPbD3D4yuAGCdPfLIoXl8hpt0fNED7/AziLCYdI7b932pmDhxBy3CpPPwbh2LiKV0bPnXev+T9kn
4WYbpa1lOoAFJTMKb0K+4XiI5YIK5NSLzZeBwjV2BJsLyPWz4yIJxYGCDyaw+CdrR9dGrPRjVvmM
Owzjm9g0lcjffxEyqW9pS7py6LQewri2rolA8DSr1s64PuV4f0ABPy/Oea3nR1VHI/ixpcdvkFgR
PTdJ/9NYvl/5rJnhg9DXZxaiXZOoILXuGhHeHeCi2++3IFbHkgflSedfIDIMLD7sxcF/aS+3lmir
AvwW0y9fIvMpaKHv4EReKVLTOrRe3j5MPOwfpgCijxKBbjNKMSqxTnBkqwRtuII461KayGeyzbB9
ZD2VPgLdh5qGazkxm4JaiklsEr9We8XywkhxRtYCTWFf5/Q974K/7AnwtvGfDhT+DdAnavzwtIw0
wvtljX7LT6cYI+D2g41DbZqJGyi5V53mKM0wTTKhSsziC2dXrLiFrNEingRegaiccFE/KzXc+iqB
tcM6iyVxECM/pk+QjxQysckUvd6VfmztjveMb/qPi0KhXrAiOQ/eoWIMApkLAPuU81fT264rIIS2
yLm1QRQcX0So/oJLAAvy+wjYlskt9jYxnkW+xdRu0L5kHyqH8hSUNsnfeDFNjPACWcCRYSAFg0Zm
1FKRMaK4hW1H/5dvmVtRH26txWW+LJtP5pAmFfC0w0POXKS8eTVwnn/qrG1GFZ6ALWRhq8lwvJd7
0/EmIPSC89cSE/1pYf2z+5graoyMyQ07mMypB66ZU2SHYre9n2QBoSAhmcMtONo4uAvf5RdaYBha
sX4wdXZDcOdLnqzgKiiqbPHQ9PY/eI4A/T6bKY/pCNMEoF5+CSKkXF8n+v18wFn+em4/wSauQEL4
UosBAgHXprTyliN0pO+m9lazrfzesO/Bx8P8xafBQDDpM/CI+66WoLPYxBq6faDppviVBAFBV0EA
5scKT1SJO73r7RWJuftjINHPM9VIF9mQ9jeoJWWTy1hkii1pLRGc94ceGvtkSLeUmzmu3Q0RKj4v
YU/O4+JGJpAeZpiHVdIfdTwlZjb/pWMYDdUD4aWirFcfMsFHqBj+mLyBpY+Wjfzvsqb9DQmezFNM
qsJ+SX/w9wrSSCVGzdXJEuqpq/1hKJPPkZfkDudLs2+/k2SMM/0XAwMgu2jOEP8Ev5i0UGYinQrz
AkVhIxU1DTlAPvcQFjKsjQy5/QnOnTTFVHDuZVcKiHQy0Lmu82m2JXmBiAhnkCqg+4UU6PRufL/c
fmwXCk2rIjyL24fF51bnCxKbH3oLnz+46p/5vQhMo0ZuRbrYls5VPnDaIy4wwvEBQSgmf4eFTcbD
txto0Q2cQImkg7V+P8F/g1M1I0KnUnsZTo2QUm+6KyGfQaNXwZzF6sOtk539OI1+yHg6gDfBzUvz
eb1uSZjb8omiZLgpI9yFJvCGDBrMlk/nSwfowh85xyjFpBN37OWD13iI96c5LYxFYZD1dVGgTA+d
nbyYWO5Je+gDTIvG64seX16z7iJ7KhiGcHO57zU8OHfGPa5yZHYEEOwpRiFjTGbYzbZaEugshjH+
9DAV0t4E2X/bPI0atzx5jfYszf9Xcq796GSy6CRcqJLpkprLkEYqzabNS4Sam2RnfRSqtTOZ5SLj
fP4Q8UMLPbE2UhiUXl6Ny8hPwlTf1TDCYr0HKEpahKe6y7l1fspjvxlv7ZpdWF/sKaFKmri33pEc
enXR5bx+pI0LoryvOLD3js1wi35Pm8KujqGHiyT+yDbYXWKhkTlF/bqrgJ346NAPerHwpu5IP9x4
KzWmCYBIL4OGcV14y5rA2VqVeeMNa7vdNIgebNLz9cpo7tfiREBMZGpSi3YNclO11xjYucYd5kXZ
TY70+y+Ttmdmv9heBAjeE18uwV1FCDQN1xncCHl+7QBlUgTrCLsqX/M3BEZ8DwVB7Oqx+4G2ftJV
ZvAajxTi0HeVeY92leFPNUgqZ6OZODzYf1q2L2COVbWh60Vn++pFjrUNA6C9MDhq32m5lUA+3Jcq
spWk51FmxwcSbR7qpbMMiTDGYkOIJb0Nszji0Ve+y3UT43g/EnrGfAZ4l5BWEBezFROvmvF+FRfX
ygsmXKnMjf5/HLdXiXOg0hgWRAt4kptzaKObfKzirJ3bq69Xzqey4JtA9WKJ7210wE0PFE5thtc2
T8udg2z5WVLE+abCZEcVRRap0aLKnMNB9vK3uF6eAqNx+0bRNvQna8gn0v/8QxEyDNcV7VnYxJZP
Jtf0su0WFY+93UZzB49H5kAiDXbd8XNqCfMF/FZkwOEmbccGz1sBi1VUjSyznW9LTS1jJPNwcJ+2
I25QPA3xiJ5pdngiTAzw8GX/ksAxFxWyochUux/oCz1lMKGcCeHlACiQrkd+j07jUxGBnGmaEdaE
Dc69k5T2G2YMyaaLb1/jSLoWHyITUOaL/GpgR4otpRQOu37jL7hKTry5nrmevYDsLmjQpbDc/9CD
Czl/AM28a/+6jRBWQEL1DkeLBYVlcxHfCwUUxMgTAmSYjy9QbCrmMv/t4hn7Hszvo+6NlsV8YKKa
9VXhpocmFBXQkfMXKZL2EkBBdwMoFT4hW0qUAkgokfpU7VCNByqoDPXckahtZFjwQpXypYDdXwG4
se0biGyKX/d/r0ol6F6ZNBKi7jDWpMKmgaxrBz8h6dsKIkkFz/tG3F9MVkF4k0zBPmHeXqrSlYkW
ljSrZs3gjzfBWpScYXlnpW8oha1cfCtHR/EBqeUcDd/d9oBcoEf5ugf3FJ6/mJmBjy6oElG/FnoR
kBjkAhBXRNm6DXNCT3Agzz2ZWdeXQm+FcGuAA4xaXkR5Xid3Dt2Ephgab3znLoOgDb7BPsQ+y0n0
AmautzOGAHThWVxeJrIARuZo+ni5z9/zMtUV+gFDioS32hU2SR8JTpFvDY2uzCCn2dj1XxcTMk1L
PqItG2C0s/nMOuuFqsvaJAWdP9vnlAJ4SkGFpeHwMwHpCcG7r0ki8q3I2s7nWDHGtZwa0QM+juEB
gDy6M3H/pRfi4ileuqs44y0ETnZD1u7d7ik/Mrih2JUQKKu4gM0D6LenSmnBdVKhpBaM3EGMxm7/
DoZBYEez0Ce1M+Ccsfhh/kfUepq3gdq2cpeW7TVEA56lg9ikM1JzUgduqLPiafON0rD9yBsvx7Z7
zjAUumBb5fbhzCg8LF+bvEjXZWveibdELFSl6g/yRaERm1EmJEJ7yUb80clMGM6NfZf9cHBNMEUg
oNlK74RFdqm5ony76yNtUY+tvqUcHNxJ3ssxqEux0MXv19Tyy+V6/5bfpYg7n6gBC/Gr2JFoaPuc
Za4Kpod+5/scj91euNGZziy5VafXbX5N1gIJGG/9rxk9JFMhLByeyDKvtZhNJuXQhCSLTN+1aYVJ
JtcrWPs5idt7AVmiWX3mAABAk7l5wz+zjs5vaqHNx3k66t9AbEaw1NRYtd1wmrpGyobx3GWMV3p/
K+7qAwUystT6a2gH55o1KRqVOUmygqjCNI8479WyH5FFwn8zJ5F5PwOWKPYtMqj75CWCE4Zbehcz
LkYNcwTK2Z3B5ABxdsQrZf2RRks4spq0FsUC7F30b8s3pgP0EPXvLCnYBVZ4TueGsdFDHvqJinF7
j7QX6VS3rsjoAmKGM2iUt4WOyMHkogGbKBrSUEYlllAhd2fzuFO4pXOOowdcY2zBA/Bdg6AGGpZW
05AN0B4Z5aIEwQ4ChC6m9IwOWnyF3s6zmOYhqEhWVGXBR39CUnbWIeFdQbqn5UPyPvIZi4zZNgjf
MQ9F5TWn+3EXFDm7FPsoeBn3e//HQUvwMeyx99WfYUcuysoBB+V79aWUpN8hl98tqy8NXOnXxBUV
pmb1Ip1F8VOYFSwme1OOqr8tPS2HNKqu7BY9LmJ5aVYw9n30SgRDHd3faazk4itJMv+3QHpn6tfE
CUG9kqYyIBVEGvD0pUAXbTN7kMQEBuHhZF/muNa0nrzoia4hEdPvmWojwstVvQrqK98aGWZVsbci
1xCLDsPfJu3pB7U7lqTYjWPu8Hl1Rld893nY4f2q9EqaEGL2YsiLHSLcjD8z+QcUIRk4vvXcJMk5
Zt2BlG3tl7pXG2PV3oOlJc4Pt7BbBBIiU+Tphu2uxeUANNjTgEPYAm5pN7oG/QnhQvasauE5Wx5t
gAT+Cxef64Dbtuz1oSH8B5rApeq3V+Zjy1JS00ggmy+8coRnPhpOrASVsN7Z17MOE/TyMURpcc8q
DE0535GYt5JQr4JaKZkNN1AlN81y4UELAvHyEbCSs+FbwugdxLm5LsvSxxWTm/z0Kr2ve8+XBglB
zYYSQIszWARvtzCyfIYDUAWhjxv6+soSPTMYWjGTVdhkodNcFtAHU1y80KlmjW/8LOrxQ4YWij3y
54gIQjI+cfhBVQ8t/RgELYtS0bOs1gq8LJEQrZE2+1cYj6CMfUCtCO7AFACmuC8hQuiw3uVSVc5V
gtnHMfEo0tL6iBtch7XJDVbKxKorj1n+k6aP8P2LaBjmfS14aWxOZgexaDsxgF1xFIP48k57Z6Zl
XOyUhRcrmwZIof7YUPQ616lBvYyffLgF/OxunHv81v/hH3yYJ/4ejzM7gv3axitg0gxnxn6+DCTV
zcRW2eR1g9O85AQsnka9j/qj4VWVoSScjULpZ7VPyaN1hBYnZR3V6/9FolW0BXKYYU08FtX5dYy9
bbuwj5EtngokSmbImN6KGYkfQBkK8+e1JsrgT3lHAt2VE32JAef/bIPj9HDwEaaIGE5vHuYOKlJB
heCzaHzpp4ghwSmLXZz7fwbPZiQJ3X27TTb+B2O4nv1C/54RcW3M4LDAUaJrdxxC5I4niaB3miWT
y3Ee3j9qBkF3cykDInPwj/VxZC/EOAAlSfI+ktPn2nCIf43zw0Dp6XvX+IsWVlOraStI9Of0IfTX
Z4uswRQ33fUWl/Vsd0OG2EmvzULi1KGMhJBSeH7JM+6xG2+eA3j2McLOL3qrTmMgCDdukNt7RWu2
YXGOoxroDH6p5G9A1F2FzosLcT6TtSuxtgv5i4gWechQ5HtIW1l+EKe6WFLAnB9TX8WlHvsf274L
nbSjrN3IpB3lhkY/Q+4hceJOWK/U0fiy+yET7KP4azieDr97JrQUTh8rCv258hTb2d+o4c5/0dQj
ATrHTrw7hv8SDuKCJT0z6ikrfUzalahz1kn2zXRU1/iZ6T7iohwn9lvZrag3mA6j9tTE0/LUhwiZ
VHMjcDdt46NU1Wrr1THzA/xlOt6gp5EHbuc4Otw+xzKiq8q+fIvRsLOTLnhNgGZf78+da0QdUXKd
UtYeadgGwm2oA/gfnNU2QuRJ2X+7Js13TlBN9EKoKPTeLh5bDfpc4NR16+/Ao/u2NV85ShWfS2MP
cDKWoskPybU859CZM5i7/uuwM61f4CUbtQCg8m+llTB0qs+15HJUfv9+Lz+wF5OALw2tErimaqUS
QJ3C6b5ojgNrSf8h8xGbsiNPlkyAo2c63a5IDdPjfvQ+Iju2cnOzLbuyiBXp8pNyRnMEcw3VRgww
BOqe5RkWLrucua/5AueQSsuDfzNH0maBNToNUCZPpXamghEGJ3FZSt0CyHkUHQELKSTqF6sXxO/K
7DhrhvZzhH6YZ8tW/p1X82LQku40GOsQqi7sQlsUpPkWl4FMQQps1arjJWG/ePSBssbh1OTTZiHj
iZsvUdTwChn7ir4dn6vpJxMbAxc+4l6a+Smi35PchD6+g5HqibgbGzPV3tGFE7jVmMfSL/0+gHWn
KQjmNypsISfNB/7Tn26OC4FkIx0OGLkGVVZH0rgV46e8tZfGf8uA31fk8eR9aRVJl45Fib/MybnI
qryCxcdH735gjxlpS/S12fIBd5phwqgMFYo97tNrFsG4HndqhHy8dkWgbqrEyyW8uu4EZyzykHdT
GgPb+Z9ax98G86s08ZZ73VyW3+yRtlxpsTanGi1QPV/9fyvCCEOBCK6+cbLmBZ5ddaUFaLZ9Y5+G
W3+ZKuowNu6B5DYQ2Wua9fbVppRQ5FB0JTM8DZFqgpavNY8uUPTFjfC+NcgOGOCLFXz1CqXjZJd9
G/H1ov44WmH9IWOcQ/pUYimIuBwCmH/OChcHWuUJ7dphjaCtdtLXe1Bn2eDH6NHSmszoOCcRnC++
dKdDANnl2UHGAXXUDJWERjFjD3/TZQza808urzh4sOrObaAaH3TTuphTfbn++4NJlTA6IspUxfEj
KY6K+7mmQoNvIAIxNWl7/YrHmnAVTTE7XOKis2YTPLgTzM0KrtrJNrK75RpYeJJu0WNo9GonF4qQ
dj926xuvYVA8cC0MHhQ7CDb3FJZCYGwbCaqsxEROBJQIlQuZwvvwtO9TL/IZmpDJ8EJTI0Zkk/mk
8oIycbaksvURw498yvhZKG/Y6vdNj9ONS5CFwohsE5lxC3bV2zt7MzqC0e+UpisgmUpplBG68uWM
Wt3RKCBW6qjtoh3oho3WJZN6+FADgBeoKEbIOKvL3O+jevPpSmuzHTRdvWfQ8kFt0UFUI+7RPD4i
om0hc8QVUBprxDDbhDXYljjdn1k189KWYW2edsCTIdZmVu+6r3yfvkubvS4jMDHAlbgqMtOHN7TE
P/9Rb/A4J2P5QLnqPi1y/2+EHCOkcMoZmSk4T0HRMtTwFZwxiizp2OghSutP1tms2MPHaRcNbKBx
Mo4OtQHVSl2O66TL40rupcY6kXEFK6hcehmZ6ul8TG2r+u2dBGLGnLg/fsPZRF84IUnAmaG/RKk2
+DIuOYXKzLGZ7Dk2KSFpsRYd5GeNLolZmYDTic5oCdjFPP+eDX05xqgMnCGPiSGM1DhA7WsG94TA
7JVAiTOIrCirHP8WuQ/L/C40bV05oStMj+oqhGPAW55zf+9uA5oKsgWTb37YB2Sv5KnZF/dHg7cO
egI+pFDeXQfCQvPG4dX3WkAposb7Q2Je7D/svIbrrOeXR8bno2t5sLXal97N2Bs0EeinqI4uciM/
sIhyBZxbOU1om1wzG+gkSxstffrfIBlTaa69386dBDV68Jb6nGzE7ZykXFGoKVRcsJjuKtf4WiHE
QAPa0Qb79RAi39yKVhW0vEIyFfesz8V6/vWQfGj6UhYeVYQwzL7O3BqTbrSVF0pxYTwN150F9tjM
lnKUpIqqFoz9zfrKjzcrNaWZjmF/OuNgYlf5MOPVzgg7R0KvN++8kC0ea7fdPU29I/1Egi9MpFmO
8Yf0RkH/X07emBofcBBsPWTxzQHmRwewTlxEVTGuWv3i3a+ZKaqq88VYlKcGCl5fdQaSrGDk6QjD
58DyziGKW+wcCZt2i/CLkzS8SQo8izuNWPU2L3IPvH8ISa82zrWpa1/6GkcOdcEmu23l7F+2yWf4
kisB6ZSrCVfh4mRq3ZkOvrJlqCwILT65sCyz8tq35j1fML+nJYvex/XAX1o+vS/bpxRjaC5GdQJf
hSSSGlG6XkMk8iZ5DwjF+GlBCqrLNMuvlfGq+c/zVzrfBTrWaSOn+IMXdYg4NQla1txZpbU/6a3k
m1Y2iQSGeVUOE8XeKZ/VVHzMHOrrIJaJ7mJFFXpNdgZZ5jpTylrJKPvwDNx6EnwlgVF436oMqyu3
G5UsDFjwK+gEmWhVgVsQrS746zhF+lBoUSypUlVPrCH7D4krfFZTTr6y50NWKzrhNFPz+QpFAgi5
vC1FfY5HHNag/2iyXpeatXva7K7IuHFhM0P4pbxfiFbCi5NsXB1S1iNkaju74zmuhGyu8irU4EeG
76mLoWeYVd5Ceea+2VHMnNH0lr2uuV+VTXI59MRMlsavoNrSXGDTLXpcn6ys1owq7bLdIjWgEaZk
Hwcfc/b9ucg8oZMcEnpgmzA3JQhLsoDRs3poeJ6IamHYxfHwLWCjPE/IIZ1VV4e2BruWeG8Wnao7
bu/bwYra9TJMEinfjn8h3rHmNUNbW+qjVshd7hvczaNzbkjr1PhEXS/XniaLxDrXkUJRjfW5guAc
HSjT5yYRUw2acgZYib4WK9JcYh0OZJzsvy9l9bK5YjifLhWRjv8bwjLkux4TpcJstcdBjdFi+2uP
4Vvtu5qyEXtYU+VfCXuSW00WaCJpOjqmc7NrDDQtD7LJuHH6hJEcJgwW3Tj5dehTIqtOvWd9pLPz
CyQyQxhs2ZKLWhPfXy8OS7L12VI8W/sWjUH14NJhdU2mOS3SmIF7uty4zi8irtJPIWcReIt80CdR
PIu40XX0F6mnyrzSKFjkeduhazAPgG0i7+YIDyalIjaeie9jcMzTR+iq5qMbFXOGHsaDIWlXuM20
nDW8LcrYAzJPO/S7TeI/kofoprSGsid+2ZGugAgA4HHzJfllUtq2+Pw6s7v5Z7vUGiB3L+ElDz+i
Gk8NiX0WLP6KX9iB/XaOv0SyorfcZfQQWQUFpoehusSVNP5QoMbwCfv55n1jGlgVcviIMotXWui+
LsU+36zHCoR3P+2HOpI5/mwJ6ZnsBEBIY9BaDEMcoFBFymRxXA06fcbOlCWI+Wviph1j7T2h8yvu
vJu4qKGyW5qbkWloYgADMgI3U+3+env353YQhTQ/JDx8yO775Dps5I974w0kiZgzn5SLT27xKUmp
4+s3BvlkTzROIdsacqP/i9zkhoAcXyiCCt7BLgv/KivuJJAQCZDYb4mwgBa+353lNwLFe4xhQJI0
pj7te8oR6VGJrMkO5vHRdvkA6aY8EX20j6AoHv0Kn3qsPYmrt4+ZCpPcC6LXMLrU47j6E6HsqbaP
U3rAwuj++Z4Tt0wRwoCT5kW238UmpgEGvLjXIsnZ1ArrrW4nYvN7ahlXDk2tpALZ89t9uEoUpysQ
z4R2OlsZ9I+Euaj24wiATdYqdH3jzH583DrIB2Hwf9sP620UeWaRqRaG5TNQs+XUrayNhrEbn/GC
lMFGmRmjx9G6uJfOSoyhe16SY9cI5DDxgxlL9gTDv3hDGJEkHRXJTw1iUOmDGcEnMdsPrWI1W94X
XGfKIsQP1PU5hJBG5PB5260+5YLlfstYv7PghSwymCWg7MHY46ienssn
`pragma protect end_protected
