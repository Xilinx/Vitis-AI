`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vMl/F3Jn+bbJeZ6oONZAAPbmUyI8nO8pr+MpG6WMo4k8R34R6Ht3+nsl7K6UiWLjHiebbv6o6faP
VQSztkQsK3vfiz0mgF/c23PD8JWj7ETGP0YG7/BLFgTUnU0R5WStJbAfmyrJhPmvdd04Mn9jKgBW
zCiKn5dL/r82xVP0N3o5klZK/09H83hQFuU8KdEGdErKKJ5cwaFBicXxaQ+7qVLR9xqZt7WMrEMW
iBX/ZB8YJWcFZVHDielKlp3r1agEYaQ67LllAdiQBVI25+YX7YvopU6k3gtuHSZ6C65gIjDGiurO
TD57ihw0CDtYs1WbGFVXBvOMB1YDT/8fLpxv+g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H6JCs5wBp0QM993fMUtscOIxGEygcaiMQd6LzQYXmdRksszDiTXRFjkGdbzmkkYxrO09AXJIxJmv
OHYpPb+SCGDumIiT0ikq+4EwqFo5wpo7ZKS6iZW8uYULSyV+llzOEGjDiml8a1NyNGqtpXe8jicc
5hQvCsrJWdjqyD1Z4fG6LEr7l3cCowu65JYSdTLqGrOzQO0MBd8oZ3E54fgDZ4bDuRGb9AJFuNp1
G4+VeqpQNWxsrYseXTtdNdbVmc1PDnPFt3ghvfdXTUaZXaBfGuGAp9B42u8/ZnLh0JvYpU/0U3VG
73M89IkwSVikAv128djRBwrqNg3qmkZOQBBALA==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TlpXcKQUZk8r/Frltm1DjMB/QV34UgKJSVDkIWGmf4WGGchWGcrXI3uGxgffn4k2Hlk0dxVVmKZT
gBx8b+BtVjKvtakrclKcKceHvmtCTXr6fYowtGMegkF+DjmEjKTCBoc307lnXWu2l8ngz9ezOz73
wEYpyR68qSsMZfDvwV/x9I/bL8fxwTxFuL7fGoG0doxRn3jwmYM1W97BqrXwDLYe9FXk3u2sSqMj
qseCIHy6sXtgFbMwg0vMEDN+1XVBcncCHvtJQwmgfnlxiYpE9/nZCRWFZQq/CnlWiQgrW6XXH6rl
BzMx+eCNMz9Rk93sbAO7Z82H8PvpP6dvygmXsQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 864)
`pragma protect data_block
BclYlr2aGa66uztbYnsMeT5EPNIPpvdvpi8Oodx8YVU1UDk9yVObHI5FXeMKLkynmUS9Oayx6Ruz
pVOlqEtfYnEIadD/2A7U8hyVbp9Kw4Aauhus1ycqWBgdrqjaFpMPoa3GJwaZQL7RpqnsdtWiuI+J
Gude/W1KLi0/BXvSlO0o2+gv0H4QmBU8evG7TBi5TgPjSIWI6qFSS7pHb2u8vHZleQz9jbaaqhCA
hiGPyZi6+N/oTapKDkxXMaX7CGyfRVH2LG/K0+k51wum7ltCsStWYmtuW8pgytjdwX5uzffuTxkN
VV9Nc8DSSgkBXzxcrr1cl1ik2pTr9KkHhwF0DGnhVoNrbaSFit4yt0Pu/4ps+Dg+ejrc1zEZQ816
GCnB3WX66bgkN9lK1fCB85iB2hB7zIttNTsTJX3zldONvIg2tOJGvgoOfUqEbBW2sZhsWe0aLoBv
nobEeb3EWujXVoGQshHsO5iLH7MBMzckX3yCASWbkIEFbJeMxLGbBgTf6yzx+Ma4vkaCkt7hhTeU
neMfvsKBCFhlhibzvee510PojyF1eJ4jOn3k1TSEiRq7G6/gsfidW+mCXTJq9iTZPKtneRWcgwPc
eb0juxQGi3dcNG5tvSdtDHMLto1uvP7hhRd0UWhVbZe5j4CE3qUp1KPd1dB236aoT47K3Gl6aGxr
0qoehAKG+y+M+bADtlcV4FqXz9cl5DBldYF0ddmWv7/+fQX9SWCrQZmKHCZQfzFertNIO5GvXGsS
5PxXBegtgShTwxqsUcZbau4/JlTaFc7n1MvEkG1jyEmofeMVQFFx1KQno7oaXex3ygsaPIwkPKq9
9PaHXHLjJJ2bZuyjAgiCOiE0q8oANioJvkDZfnzfgQ3HviqcJQi3rdB44Ht+pazky6+u5vT8BLAh
DJYknhHAJU3DrFlvby4DTk4I2SYCQKbfmClIb1OCnKXFolbnzbvYbaEwE8BkMc5LMjhA8dIAAFZU
qXoakIxaPgdzJ+jmZsi/GOcDLXRKZnZqHN2crppvgH6xJZBDgbVtHKXQWBpXwkqKoo4lchPQcL6i
PnjO9bAbkahm85drBR9Kl9rR9QLTqq7TiwhyxfGwlaLmBfUqkfL0H7+wQvDprXjj7JWMTeGRG8Kr
0IhjjxDZSlFe
`pragma protect end_protected
