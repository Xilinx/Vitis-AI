`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhedE81KxtA9xXdNnI5GE1hZLIBUrDtSvHxPXYdxW+I8di6Hea1hWaKdVE
mLeFVggHoBkNBbER9FrvAxORBWa5psFkN6uxNsySt3aoN+GFf6biOwQ5fqwCPqq9J8wLfwa5Jsst
n8jHLw54O/4wcCXiO5Xt8H2TTxVH9Dnf50BrWjyHMK5O5qC//7IDYaXWEC/NGZgiq2i94r44+3/J
MSqPrXP8HeXbaQ11gInWE1KTX9nc50bC8KaMva6fM5Ij6Lr4HvZxx6QNvFdNP9/e0HhZbMMuPUVc
WsJhwX3LQNVlIsOzvjbL8oy8blilQgREvgiYE08l+5JCGSPrjz20VNGA3s4EYvfTu1CQGx0uFuqq
iM/BIq4HOie/ULwlE4mpwF6ydNxP000LPs8qTh6eDAfMo6fuxbefH6VOBiPeCe0Q7lDdNRnZHsW9
ewFFv1fwh4tk1lJzsjTAptBC8bKwoGejd/yVKNSxi6CsATAUT/DNBhMJOTxoYc+EVUwVUw/F6zGp
h8epFuvViDB+z7ERQzB89biuF1T2vGOoSM3zqiiVYi8hvFuCJnubYV/suEJ/6SZD2Ywjnkoep6EK
iBwqIuewrgPJaVvsngluBnqszwejVCXE+VsZM3peWDOlpHgGtUVE5VV9oS0MyJA/XhqnCI17G/TV
OTWqZvaem2sijiuGmLmuKdmqWY77/i+rESJBc5MBj4dQ3aC3PfC7jFm1hm0bL86OIejUTZLco2R6
NHpVbJWPUDOHmk4IFkGocJRw6UR9xbiZl3wTb64EEhGAST+30tkbhg1gfmmsWP2oy51s0fp0PPFZ
Bih7J4h+e1jXQy/Qsltiy1qhiaIJ9uZqL23fOildaodbXboQ7XLNwlq5NTIIlXbIBUtuiuPzwfN/
99d7ayYVK/U/eX3vFjDiQpFpRitI/PKBxhcdN8+88BzzTQ/eXd+xiPx6vD96+Vc0j3mxpGZolpij
DC8u/Bc2f8m48xKdZdnG92avhH1FUWibFsOJVoe+exuARznnIoEAM1tj0iqm5Y9BpQO84sG4yQoG
G4T1LWWCOI9zmVXX16dEjkMBDSjOpCI1a01rT0Nun/BZprUMfUFgIMg56gsngD5FiaqSRH+dm/EY
wEdEFOW7Csb5WV1NSGQUDdzB2218DPgUCr48eHq960o+5J6D6NxPlSVXVlpvXH7oeqnmcIfl0aAP
dxz4fQgG7yqQNtU3K+u/v52JHYwt6nplYDv/Ew2v9t2fPwMe2FJtXDwo9BswzT8zVt0lEjQy9W5X
ruZ9rzUiCOvm7Q7QHrEdwE+RZNI9tcHuygOzgSdg3Xk+bpsxd0VQe6Swi31BdSPi+5eXjeAX9zZC
O6TIlbfaBqdx4u5dG9qDxTG4h6CcnzWuw0V2AxX+3z6voCP3sjQcZp3oUKSxYF0YdHAlkWAiCE3Y
UQ9jd5Ir2WF+33sOFNJxH9oTVSJLPZ4KitL+2omN/xHDMN7Fdwfpsb6lVyDtFzDKUVdiESamNEsi
aaLbfclfqze77N3PjGYmvL3bn857mYu11egpQmIg78zTHj0H1cV9eGqRvbIUG8+VE8oycrt7XHr7
j/bM5Nfy6HEDEEjKxZ23nV/xojrJRJCqyOmBdgQ4Uvuxy5zc5ouDJSoQqe/BNIafJlcAjG+dfmMs
d5b4hAHFsOxODY9ZOyEjved4x8rjqg3+u3OAp74CzSyutaoBSWWwWQeJeizpSeQ2XFNl7lpJB5xx
CqGX3RHNNj9+3BX67CiuvazKKCQJk8K8az35JKfQVSK1cf7PiwDhGakJWGj7p4d+9/KbqJ4h31xc
miaA2KL/OzXvan7KLM/ZHQaNOxXcPE8t8o08BgpH/ahGwvQXSX05HvleKpHMawbSuSwuHklrV/MM
GQyDChw+Epyx1OqpaWOaepQwh4Lld2h4iL4PIVZatC2FIjICWHIlZKeHTR2OrcYuKrAdQ0fQpH2L
BZBjXdMv70j3WxAHBlcZEYsdrv9nJXaCEKRtcvG69ZiIvVmrgAAttMvj1uNkhsLd34TOzL7EuJfJ
xuroEYtld6T8eD1x14+FVp8T9JpBW7gbKupQOoRxZESyPXeRYtQmiQwmqdg01BTlAyvnu6dU0UP/
rWX91uSQFEV3t+OuWpdzWSv8U4ma5qawTlyvitXb8FT8sSDW8OcUBZ6pnkJIs5bJkiBiwt7CcGwh
cO2Qqx/qpdUReTTvKlPc0FcPw07GGHp7gO0bs8COmCfz/qMDqP0/aBTrxmi7AAWk8VOofmGJCEK+
vgnSC8a9wLm39pGCiXQqlu5hYQW7ZG2gFi/WN52t2tmZQmonLH2V8yO9o/Z5p1z9TBtoFajcUL/L
lGaYQnSf7jgYg1UjjUOvc+GKt5+fFa1WWX4VjyI96RFD5WnGND4ifEApybU742ovFCZcHbJtByoB
bQdIr1c6/YBALKU7aFFUxX9bXsAZigYNW2hZJmk7vEJEwV0ipOnd7XjixyydFYUz4BzmbSSwHnlp
4cucSaL8uMA02AyyXUBowrLMjmJcOV8vzoUKmCM8ezDJvL3GPckV89HdnkX5zVRp1i8p92y5u6tn
La1vNbR5FCi3T7J/h8QaLhLAQesEI25i+gl0XLj9Ukwskwsjy0DtrkT4NJm98IPZkihQlPXuIW4M
jiyYmUi8WG8HWWVzrmmd/Cj637sEmSTmWdKM6fK/blpEQj1t7T4yGAebi3M7HWNr7bZitec+f4mr
qU5peCzArHoBIpFncypNS7KgsFWm/RkClfElO2ANhZPEty1iocVvywlbuq0q6JJRZ/RksrYnLPmc
XwCCbHz/qCMG4aH0hSmLN/tCJaNenWMUX5FonznbfphXxQvOCTfQ+wTO2nx+xzAx89vfWtKiNSZn
1sSVUXhTXgYdp1oDuowd+6jg0o8IgsvqJSpkTKKbSPqUhYRf09tkWdK4e6KUg3Xrwvrus2ZcKB7i
2gdILQWm0QeX7MqSsRzi20ghXtWKkAIfJtnel9NqTvlSV92kfjdSnY/BAQvbIx4xZ5Kj6DRqFldh
98Bunu2zPxx3geUoobTcqPxkF9yJHzJGyvkXebqGJ6lBOnwQamwaZd/bjCaW85tyE40FMZPIhKjk
FePL4cKTrcyK8BStcKsrvS+D/cuMRON7veUxRViklBNKsr2PFsw4VvvPB+QTClM2ItB4YGeFGIb7
rESyoVjb2pYTNW3o0MW28mNWcgIKmQlyWr1Wk6AGJZyh70U0yLBMfja2qYwEHrt5mg2WomrUeW2+
9O7Ih22kZ8yHr0eKcUeXSAXEtZQcB5/zVp3PHFcsP2sDSBjCXSL2sj8lw50VJcHRp4HMX16f//WF
y8Pwn2QoJrRun3Fi/qlqFqBAitcB6ITJmZo7XTkZBNxtUkpy6I+G+nc5ZjeJjtiEcPJQViqlqvMc
NW6PKCiQwtYfgYJlT08KUBUabol7Uy4BZmpbwwoFbKIGG6Tz6PuECdO8AMHGVoQFlb4j8G8kxfjl
lyTGBUOpJ/vS5BHfR+cXNiuaJzghJqicgWG/gwFUyTTyVhXUVz/vvxVjwo1BEyhuciM24Oqh4auJ
7nhEB7rPbsdaUkSUxDmhYQZEvDlNppl+okP8LF8opGRY9uf4ejyoiHZKpHvUnUd376hLP94120g1
wPFwGqZ+D1YAhGNo6DARseurbRW+JiOKxttcr3+h6gMnh5oCsQ3n1AKss+xnvUG7eIPndNW05GR3
zZgLFRPmZOLZOJL68wQ3kzg7P2swbz3zZpJ1BT7RH+aTQF8Ld14ybZ99IgJO9s39MosXmZlYIC2d
unbZByR4myCDCmkKUbIZHqyWVYkkAvsEFshZWdVIZqcfn/erJrWOWr9ZRo23Gs6byEo4PLK3JW8r
cUx9RDYVzgskjab0aZ67tODQEspP0yEINeIqIbLfvl5TRccK+05C0vKhL/hSeLmvT4wP9GeBoOP7
uOgj7ddUkJZOusrvK7vbIgvyb2RNn+l7tJ0o1cmGS+M+yJcWJhu55IBb78AaUs1E4Tjt9rqoyd15
c2xTE//L1PK7n1Qzg/6LsQu4KQt4wSTXPEd4MyMGCSSBK1VZHpIFHu1jZxuTMV8yldhwkIrQT0Rm
XuzX1AnrGxNrGgcGQxmMY/4ETFXFdC+x0G9WL6UEC6ogymcV/4PGsrOPzbndBliTdAnk8lYPzvXT
C+fT0BdtEieW4nm/Vp5zj61m/MtHVuJw0UXzQb7dTae3UbXxqWkxfQwnVaQBK1EDvO4tEAcFVX4J
scYvQhUXQ1PTTPBaeF9odEXzJno/ec0Cuo0G2DeGikKsXmnnZcqfHGqRakNVsdwa8+vQF3NgnbfK
01rB8YkLFTIFk/xvPcXRyzapHZ7TStkJK4RSH79Cq7eYTLNeGWzRAGWLcLTD2g7O9d48MMV7j9wK
a4GSuau/U+BN608gvcGbwHzFq2iRFq5mAqlYVr343bDQIZK2x2wr9brrSdE0VDglcOMbAxgej4en
4RMOnCFh06W6ShDkcZ1ZwuJlNhbPHWnDmn8KzZB58Z67DIMiOLASFi6QZ9gATchfF/43cFX2qS4/
eJS6rg9XQmeDkqbAyj3dz7vr2Gg5DoXSzPetcAibni2enpd4B+XhsnnEdckrkMmQop68c7lusrsx
Xzi54SwwdJ05J78FdVkk16TslKEPhJGrN0NihhhPhSYpytuv/NOyls492i0wFOPdRleCguVyIK2a
lxmMidF7rFcfDvSTE+dGQ1rlozAteapfDbL81N2pILus9aqZixfzf1YyUGkUuPn5Xh3xVrJPK8ig
Q3JdUeA/T5NTDi7v/iKGjJOFRWv7aX0r9Ue/cQdiBcu17kmIQHlz9cOYrCTUjwsTzOkKThJyUNkv
PASBN01lxXQEJZM+ZmrzXR81VTvlqtcfIPLkImsGg7zsMgkjmdPV9bZAzjgSB0O4diCUyUyos7jE
Rjun9K4tIApUqkQvbzYExvUczdCzx0leLunWMGIExgZTZSoQhPh4DoU6OqYSu5IFdAO+i/949E3S
npMQ3RJ7n4cxdknOA/VU6pFGGyPtNajyiDQKqYsX7QHEiK2VVSCuzZ/f2G4t2cfqj7vBg1snalov
RrMu4TE=
`pragma protect end_protected
