`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrM41f83zxdpq7B9Bxc+63s/ThO5
lR4ebiIUudrMSnsXzTRn4negwrrB4VipTwcqyfoZbX2gIf3gPwkP3q41DFrLyf9opSDFSsyylvuq
0tfuxhMWxI0KvORiuv+DLG15sEi9Zilc4jLqmJBgxaj93813ixDm3VBlIU1BQYAYzQ6XobruGhlp
W7l+H9tAQt0BvNuSDNd6KHRHtkpbBcXPwpTyZJ7RstTWqPbVIiCntrKr2mKrXFSxquvkPLZLq2tJ
HYWpvRFENhYb+owwD02aaTtegiWhzVX3slkMrIWj2KVjzVejsUmxLEN20l+AmBdfoqRUVfD0hPkk
Gn2HZt1Y8LgSlHZ8b8u3uZl1v8mlUEAqWmfk6Nm0kSbt7Uo5tM403SNpcniXKtxBK3m66f1qTV65
32RLR2euavz+BgcADS6174GeB8+F3OW/FkyahBv+EZsET873uEl6gUplps8f6eOkldEgxQbPh8iS
9TlAwAZGT+v4TsS/7FtjCK6KFZe+iUOWGytqN5v5BTkGziWo5TgMfyJnCbVAvN3OfNgUJF/66yE2
9sY3l6u5V/FlHGUylukZelb+ZBqHP8UwhU3gYNXk9MGjdzKFPB1ZknfM/HKdkD4bg6iqXwVitRoJ
UqWSwp+EWppkbXw1GV+onpAzyc+nGVRoWH2Rgd6iLjVxY4BFIqU0ZQhnKsUVNz7pIABMCqN2pDfx
r4QxWCVZmMr0E8lRRJSeKgnpd7rTU1/YecO/2T2oZmhIczMbtrggkZ2Tag7z1BlwZp8UAcj+JtaQ
KjpMQElhFM4kkRLaix/E7J0GFkyi9aC7+pvi5uVAjSne3IphMKMmGVJqaRPx6h8KHmpVmOBcYJPC
lx77WoIi0CfPNjRmT8oa7dZLzsyt3i/nfchqgFWU7sB3iu9lta6iVIgkCjZGn3KjOfuHujEhG7P7
G2n+8BJ8z+rQH9QGVSIX2tfArEYdIpubY4WnK8DwTJAnMwcr0fH+gThtl8/3tFTZb7nmAuAgfk+C
UIYMYbB7+lfABket3vzTZqNIEr6BOR5GmxuXgrQA0OpeSWGIW2zunqHbhye962qipRao3mZO/od9
ADo2fYLz7lpzbwsKHwFTVZU/Rl0V1IxnGWXlESxg2/HHfcSolmTIsjZ5tUu8CQWb/jHG/lBvKXxG
xqmu4LIlJCroZ9KQgUv5ZvE5TWFssmV6VgFvQw0aEBj69sxTCsiLNdEmirbggmspzKW9wgtOb7Wp
DfZeloRqLFRK8lVQ/w6e4aXamWouE68fe1gSDce/eOykhEecKB4MpFXTxTJHKFm1DehsJDyHWMTr
S6V1qHCV3YQw+AC9cdVhz6aZqN5xKsdZXW0SPWVTizJE+sPwepA6okSEwv23s1fi6dL4r+hBZmUq
tl5Z7QEM+pAmQiVklowZRprAFi+WOCkvOPe5fNocvjeky2+pAdZLLEMtM6rqndqMU+2VvF5meBtM
1xQNAX8UzEE0rck5q/7IWOMvJHEzr1ccytYtjyr36HD9pE1c2VPHFsLUV+B7QCw0kxA1FT+LfG99
o7cpCd/LsTyyd1jtN4R765SkE4TyVxxVS07IyjOMXsFierg/DMxF91bG7o7WBLshDSwvAwluaYaf
xvadv5pdrBM+tvdOEHrFKacVHmRAZhKniOnGe3VvxL53mm2LleyzQLEStEofDmK2uAlQPIPRXs8V
A34eZF40hzS90QXVLRO8NL5eMfsdaTZjkhZCHEj3LZJo8OPSlrNzKcScuaodxF/iLolag1f9dSmM
0hS0m7s4Hl1tOu3meoZpH5uIr9JqVVko4oMhrVMDNbf813IC4Z5PjGTlnskJttwFi0BhuRN3XTyN
UNRRkXvlWbZLSNYPW+S0fQUvFiG6OrOWZGKzcwlHhKiVJ01qvOeJOvn+K0gb8CyRQz0XPnMaKDRu
xWSFistK1IhzXWx+Vgt3SRdsG1k8EHRh/V25AnsuBhZ43MEDbLEzgsDeQYNDOtGW5d3cLn76HL15
ymKyb24Z2+gSkt7Z8MPIHJflySKYvstzAA3NFqih6PhUdtlWrBL+PvTUfT7AwUrLTsy3Ip6veuO6
O9lAGH0NiD+l6JJTuQpJ6J7QOLdE5bCPgRopccHE8NHFa4Tphj86+T2ny8Xbnu5HSCbNRGYHRfP7
R/s+Huo/1Qyw5N5342dJO5ka4wr8tsHk9SDMFtB/PbYaYNW1u97LIctUw7faue3ywvcX0TazqUjf
hAyYVQypV847CeZIkfncss0jGS4mKWWz4vW5tXshm5Vo/qqjq2lLuZ/2AcOBUEE6XXCAzuKGQyrE
6IiKxs2xcx7tgVQAj/I3AKwSjgfBZjAFJP9ktHCxtuX59MIgGg30epMabFzqF4KHVJmmI2actxZB
Mog+lqfBYx9TU0riS7CZEeT8fsm+lzdVF60DBGcueMriHZSB4L8ffn6nPUWjq4XOgn7v0j++Wsl1
5VY6PNNKxg6AKTiFkFgSR0sVetUAmtgh1v0l1pryAJJAAMgyssQxuqyH2q0VLgIh5syfNQ/fKZ44
45kTrIpr5w8+dAXF1gQA1YMI5Na+dT3UFv4+WW56z9HEDWZY8Nzu+nTp067Np37GnU29AZ+0x0Xm
6KCKEjZVGLMlMnONSV1qoLjXR6niJUxKJB0BtlQfyVST9r2wppOLSmwOCcuLn1BNABRDakONydId
yOsTMd1HRatfSO/p3Dr26bYJjxCE2pt5JmYkJZmOER5uyMTeolqqqW7DOLwQur2n8l5Ch7DpdmKW
ahfaBthDcB/oXl8IV9uAhGiYLoQ0jEDXkGZcPqUh2El3IZfvkucvo00XFObUydN3ozNe4InAVaJn
NNi1uoqloQ9X0WwhZusOqWVwQcy1poqOEvpM+xASBt3a5hScDU7nBEqxgs2WYxC7pbmGkKv7984k
/8sg4jv7KK/PNUlJXY8LwQ+hXONzpFGH3szzEclNDNiZCe7XhoxASMpVZPEOr4jQkeb9UW8SX3gT
0KJt8au+FLBgui7nTAD+d1Axba+wX+CgTMRSd877nqLnMaNX0Avx7gyolBfRWovHY6bBb3Dix/yQ
59QtN4lxR5Mj1BGGL85WCpWu3IfWIYA7BUxucDFY6JO3LDlfER+5A2VZ8cZFEaSjQ7gvs68BNFxI
b6yqLMIrdIciE7a1zaeA8FVWdlqB+QOwJSa08pDYjjr7ATHZQwy4xkr3t8SNwamBxS+R7qetDxxe
TYsyQtS8potIUhoEX/s0X7DbrCcB7n2QmUr8dq7bMWb0pNxzTFN4aM8s+Hfk7ysJF/zXc/k8kD1M
WNQTN1QVeCTLUK1wdqr5TUJxRz2yyhqRaJnw3K84m8hZsIgeATZey6rbnQcwRkxpediBpxGiipTX
sy1/VNNPkLlgpnbO88+y6Hue8WvQQVBLEG4PIiKMQLCSnAFeWAZluvaYvdCT/r2wFrIhSrormoWn
JL/IPfa4xr5S2UErDxUP6ZlU0ib9dkZwHTBc0G8zulD0GS3uuU4cl3Zh4zPWj3/6hrzXPCB82A7Y
SMIZJQq2+LiCB2E5lNFXcXy4hZxd+Da78X2k8r51LAIQ2joS2T6v8yDrx2Jau4tvCUBUtz3rTkO1
soSeAa5OOvhqmLGe4NNL/Tj7RWci8B2FCRyk3xRBk1Q7zx2CPfJ9wS/GMq3vKVTFmTyBf50DVhHE
ZCLjwwq6c576yEZiLt7h4loUP8JNd7s48WM4WezkwbCsJKwj31FHSLoDZ2JC31SVMTrux5HjccXU
DGLKibPIRzcJOipiOTJyqyQ7ZYFd/P/5UGtCnki6AgDpS+m2x9ID0VQXag+eNBK3YxZKqVFVF/Le
k5YpFMhekHh2aetF5t3N/ltypEWVaYFD8Lpyhu+rdhRnG/jbMM58qiGsRiFaJVFq8FRwsjeTJsYY
thxoG+iQTGEMQjTeVF8Z+qnmraLBjpxFxo4oBA5bXQd+OJlXvXRkF8C8pt4J27i2EWwDi5kVgIGU
Tfp6ewbJ3JZvQPADuMfr7A6RKjBOfERym1Msb2FlYAko6siUVzC3hz/l6Qn+lg/DYUC00gqemwXV
h5enGqnSwl7XZc3njQowO/Yitank8VsRF+iiHEJQE84SqWW594ri9BOKLGHrzprTFsbYn2oeO4jo
YDGlb6XbXVVZaT97KW6hVtfLERPuFi2mCmjcLMgWS0zGU/Fj8J6mlEBHKTFiijuVgEDaik1EISUa
6vMhj6OIqFoIrYFQo+nO1+UO2wXpwcyUGAF2Xln/nbenWcoBYGx0Z+JsCOAaN+q5wzO/V/ISH59t
d28rjDNq/hwsVku4rXce/ZE/yKxwZ1iA8o1oH3HboVwvkSghiYhx2AHhNnp9Hh7e4yZRNfMPyhVw
hKasBC4WqbyL4ZTX09DhgQWPa7CYWcqidxrsRyGiuyMWMoms/qUHDW8Rr9yDzHZ3lwcotz+/R0og
kcBqDqH8NvTgyE/8kFEgwhs/bXzIEcrz5jB4dVOj1cMknB2WNSQbYmO4tF0xAKBIQ7XPuZ2BVB3M
0PuGm0xnw/P9/ea0ZrmILTYilE2wSgo81N+hkQpZubNd+5hb3kETwlPwM5u1xZ8PLC5RM6ijFo5O
oKOiT9kOI1dRaV8yXzAdafeIYs6EDwL7d2fp74mOspaoiJheKmQKC5HI3C/xJOkP2vY8Y+GffDNO
tVAjZZXP5HALiaAEmIKiASfox4JjzYobpJuM285dkwhzw9lhIEQGfTqm/af7a+b+ykTIVQ+1/Ubr
2TUMXAGXobEd5zLkRHQELoxfatplQ9Zr6TiRR7sqlbxLuyiZgpgpv89MueibDEPNK4Xm6FHfBDrc
ShqWPL5VgkdwJofDgtkA+gNAlqV2VJYDNmEsyAkqJVkJjaBY9JCIEkN6CnjOFwCTdVsaC/NEEcQ+
r855qCRa5QZJDngP4C0ik8lTl4b/BRBI085naOf3k0HykTrNaVpVGMaq+haZsKW9GUdZSTT2jKrk
m5c61WKZ78qLJf7PZpHKrFe68ucOqo2ZS65x7MabsGvHQanDRO7qid0u6oKAe5C4FbI6CIsvbGni
a/U+92GXABYh6ZV5gLRD5d39RRQ6IR04qF5jX5JIoR3zCLcJeKHykS0TerkIuj0D0Q/Q0NhBhcwJ
iiSZPJaVPNv31I78rL6sGcuMS0YQTuaAQ+1GxvA7sbw0ucYRbMOpql/CRtMEDn0p2m7CLpUBfFDG
leOjxFfnHlBS58uZbbXlZ9P/GDu08Nl3tvqINVJOSPpZxVsGFaMjGFcULpBpGSkuldkbOCPPXwEs
9gzRDRx4HHLv+/lsVGjvEKndaW6qfWKjlBLGmCqI+gNB9NPkSqk1+sGHh09vtt3ZQ1vtJ8w4c/ZN
VVyw9jrtqgKUMQg9rBiVGq+isfF9S+EuUmf814juYjjj88MEgwHnaGJKEIydBBq6fnjDHNdhzc6u
oqVWWJGIG0HecCuexB/Uh0SmxYiF9zNkmLg3JdmXSVn8Iq/alEAZ0NZiEhDn4BKvditEpKA5SCYz
7XEzefyuZ+mqNF1Ll4oVltITTzG6xbH4iGuzYQ9CyaTRQaH6vNfouESYKR7X/7KG41OTKlPUmRAb
AJB8tiekb3vwIoTSKsybPfnzn3VDIK6ugOzimDCAdwk6WJLsBhbtCmUTHuVEyBIdKDZoK+BY88jP
m7JRazSbPOMm22glP2+oJloZG4ifMOJm21pT60eHFX7gUpQ6k8Emc3pF6ezHHiLk5GzaG5LOaT96
K/bxu3uRuspVIFVMKpxh7onHNucabCFbqFsDCNnV6rD3EG/ZiL8lUP9JcBx72oS5RwhURdnRGX1g
bZaikiTGRzeywq/vay/2GdfnpU9wInasEb2dTF+O3FgNGYAsnYYIdzkwoKVYuSGdOD7Po6YgGSsV
6RlOfNOcEQGD7zSGO9svgCTfg8ZyBRrmlmVUG/mMOyhi/896rHRkbToBlDb4uduR6i39POYbFUSC
f2n6Bg0TDRCtdIhWtBw38uAr3OUX82ybfhAT1qbokOnicjDxy8ieGAFMIFR9vB9cnEBof7dN6Rve
Qh8+Cd/FXf8biPD0w/UkX7A+/WdUjQX6igCNR+c0unITMb7k/u6ks4Yevu0kAcozmIp7jgkqglYa
Y/tTEZemC8HPWpVwmk8EHKbA0qLLcxglaojwLrNRoScBcy8PsVsAqKn1XBr/PqzHTQSc2zAo5+hn
14cTPNgiSrcNMQRoKPphlLiiWSfH6nA6NXTqLfWIgmP0XMtuz41naKJdzUZW+qcj8m2FtKP6jV1+
ves+oydAwKNTPLmMSlSpDy6LKHMxVK/qDSxOJT5J4bus3V3nniW72xPl1kRr6nrkEOzS7agc7etH
8PKw6HkpoXjXRf7W0jVcnMZeZhNk07HcJjTdvGWwNYH7f8EvXtHSh0GhQoWr+CI6gzdtIEUkIfmY
bKDHejscXG8ZLmckDRHnvQE+kmWdatMRV8tk3MODXLUGsrKNNs9Emz6DKS9NA6pXYx27A9k2xrxx
pVnUt+Y/9QwEHkai9E74Mg7P0L6sf2QgQhY1C3ishatuI0E2Hu+gjE5EjMFIbiaHFvgF4m5p2kla
saEeCfX5jTL6QhRxg18AvdmQZWySdzmVtdcCoWkk2G6KKMd7S/YYqUBjwg0OQggf1ebV1fYii/Wf
j6gpAzRL2jDw3B57jrq6D19SbfWozYUQ8i5dI8WLiKaOiCDaPSkNDSOOtWU4B4xHdMrvrm4mf13Z
mnFmTHFhMQ+ticJePAjumpI7hPq+359qtOA16QiODnjpJf0hk2b+d56r8Bw5rBncv5J2XhF2I8xW
jSGiFIaNDSppN82xZG27WsJg4ADoNXqDSOXc3sRGYptMuTZcFXV6FCCF4CuQCRIkbjyM6UmVptdu
rpPHxq++xY0apomIzEgIIGFhpcbZrRKihb71a4tqfbwYZ5O+ihQyWOe63Z1CUc0vE/o69Io8+OTA
GzBkWQa4i283fWQyO8rcbCsOR/bnMuicYMUdjWIPF6QrHDqyrvUBj7PTiA96sjtSfxywXFhOo1Z5
A5oU3h6yR9vdf2xA+58DDH7zlDHx7yNUjmHrzQqV72YM022wxuyGsjEEfO20tU0cJuK468D0i634
3mrPYMcgZDXSXl5LdygwvQLRf/yNbV/IOcVtVNL6t6A5V/G/pBj1QuH99l3gm+j/IWhS6UbJIqiQ
yE0DkGGfyUWdCOHiEKPcrr0WbiQHuBCRV6JO2dO/aKFjWJUCpLtFiYNkP40eit8DN/EfBF3s6lBb
ecFeVGxS9a/Q2eo+rRcjcDeyp9yn5Tj3ztujilI8DU7T6MxBuwuBtZ/weVs7ZPw/LT5kVbA7EQ/3
qJgf4sIuSJZOfCGstWkQ8ZHgvqpr9ZPQ79Y65ge6cqlkpq9r4JuBVsH0q94Y7YSAm8ZlZY0LhjLA
JUsO+/Vh9PjWpeWyUKO/fus/pxAUCyf/6oMUlsjJT824lzvsD/3vvW7lnnbaLFKFLjDxXbUruWp9
tDlCTHic3rVflyDKLY65BFo83yYk+62Hs+OKjMEGXbNvi6c86gc6pEbPLx/UttM6/36pSIn/qy+F
2vOBrBibySpBVCJ4kLSUwapfvtUjKeElwt1ecpsrGPqyFecMg9xRn3cjYPtWw3yQ9VagLiiFa74k
tTrNfJ6Ga7LF7ZfV1YOeoPIZ19i8/nPS5Rq72fP4ekXpYsGCuckEM3yZjPImMErJbMIsJ+WqxXvc
tw8DCmqKwv7XJSU5+35ENXAyQOyDa8nmtQjjDGQZjHKw/NSCsfFGOJg4q2rdEbW63G+V/6S1/g+4
TNSZZ/DtLESkmcnGqRzxoDjOjxqXUZSVZKp8c38RwW2SJEQn1BIJnCXkzGkDA9nVVFdcq4EILqMm
cGSJo0GzwfLMK4M/3SjZClnPg4rXFuPc7uhPwQumOmab39UciIOXaqJJTbfsEcEjzJIpuv0w1ET2
yU/B9mccTqj1e72iKWVC2SxdZ3p4JOD82PwYfdVo5Jzd31Ehv2XjNtBJITrcbr0p6cM15NMYADLh
KBo8YkMyOzK/asUP+aMMhwZu3/97KAyVwtxGHhjXQkWGEoN64IgI/6zpg6YnKc3NRK0KqqChMDCN
8VA210PlXv4dlisvvhuzP4OsvRW3BF1SNUcuZFbqBMECZiPbOlWWCYM3X3dOoNIB327x3m4ZLyD9
xRoplEHvO4hr0Xff5rWlTLxCd570M8VmGLKRYd/kVxUOY0jWCPM3QnONEUNQfWcJzozS5hzSzXbO
damSnd2ijKBCPXK4gOthZX922qs01+NJ2feETY8GeOjdwZFDMjFj110US7V8AjJW60YVIf4iGhht
QFkhDR36xTOAMzetjOnyJiX6M4Jw6d6Too0EbLnXvEN8SEdobfIbfrJnir9HH7D1m7vkAsiznwB2
aN1DdN7Y7POatXFiIrd9msMsVk8uoR3Np5RAYk1lQ/jUgGTcpr4F6iWGbitmbpXDtW5eXpFr5n30
8kPD4/AD8UJ1BPoEcFQB4twcXImupVHIWtMGKsvEtvqwtMpspbUdJC9gMhjs2phLD+ABJ3yecpOy
A9n0PjBJ3NeIfbZi+uZduFiX7zEmXfECqce4UO9RKsF33LFkZB0MlDAU1u/LVd8+5XpuR41FQOOJ
9DtK+CynH2T8qkVZQA+8DRk6gO+LyiSeWa9qKIFfrxkl6vvPYDQEtnkQAUSlfVshGCwIBbeBz4CZ
4TWSZLjy0HyhCFYxI/kdYMpWf/CWvdJfb1zXEQ69tM4a+lHVNBJglJtRowtyjVmt/Pv9zWIp2HOE
v7uvWFKBmqkG9CSBXRLXaSlANiPVUgNfi6GM9Rz4oLtl4SFyyJUrLPXMBTRtnBbDoxEX3IhN9cWk
x455FQrKpupDq0JRuln67ffAiqpmkVzEERVOHVoogREusoS5ArSWCk1cZNQLfggH9BNWIqSv56p4
4vJt0W2XE5FDkyyrb3V4rwMbuUud01XC0PzA8geZ/2eirhN6Zv/P4vWI8i14JK0QnJLuLOvPE4Y9
hHBCkcn0tVgwNjPQy4TnEkD9+bKOhJhrQGfEkMBBgxRIoqNDopLAnOhOEEk32gQyDTZluBxGCRIO
FwshrRAK5//rRZlIr7oQET81S937myvBvf3WjmVm9UJUu9And4/K9vdAGHySYnQhxjd++5f+y+A5
triz0w9kzGphUNilmKWI+bA+9Ts/qS+zqKmKZzp3Gc9dhXKv9I4Sf9PJUUhT308HxmY9H5TtfsHV
UKrW+nz6ooMiFcgYl9kN+U1+ZxcZIpgn2KCuAa2c7nBiOKYO+l3yX2rsrRMnTE2sXt1qsf8RpWCC
DjmQG4p5e38qIQiiPeGOxKNTcqB3H969xntXAGEFueaF6U8ZDFNIjuQEC8PvVObcidV70vPdgBlU
UrQhWgn/q3rV5agjwS4JuE8ZtU8IwiKiYRzC54I0/aE/7D13wH8+WTdI8JzAVqtmaIVYvGm6b1JU
KIQTPW7rTdsMFinrcdsiQZEzIu/i0grSBeevqlkV+EBBbE5TFVlXc6KOVh2aPw9PmbeHJ8YfCBVm
2Qkz59X91xrvAUJ39CcdWBopDz+S/UWMSsppt81Vx7cYiXhO3iTtbi41zN+wOxuSwdEk10QoJJ4P
FNxbIOgEsCeUP8w2s/wXTP4JapeLrDxdJOZq4SpR3XxQgJFg2vuiIBfLTw1w6dMLzIXhCQ8HBkFm
f/rFdjZCz20yOrKcU+Yj+BllSF3fLx2kReeaAGhu2DQd6tgh0cTkM7yJvckJjyeRONAuFQIdrtFu
s1cAz8OrCLcswG/FONmLS1lhQa5tvSwGC/ehPMajqOE5Au71zd6q6wO44B5yWi/DrO/ldOJEa0eb
Gra7a6Pa7VZAhNNg+6AVynvzT+e7rb9kJt711IvH1/8ErSGwnrcoQyY5Vp3iJbEHurR0CA6H18lf
tzClbwZTADeUFLccOfeiOlF5SoDvkeQZ8MyY5ge3DGhBD4V+J2J87Bj1wR6spu9mwlfjfD11gqis
nxz0EFGmSB0jcENRs4U4btnzFOOFIqXT5SjUOhaqpKijtXPTfz9iwpyLn5rcqQ7BImr6r8Sf4U5t
42ifVz1Y5bSFM07oVAgltBsnIe8zWtY2rNUO0Im7pkuD1omCOEAcVt1M+nAuOp3nu/2JO1qtRoam
hpS2vi/8yDgw8pLtQto4yrizoqWKUd5zGDWpqCNkyZWKARM5ukhw4wpaXOFAgPgaGEGW8m5CvyrD
fcUe0LnJ567x/5x3lmmN/BJn/e/2Uq5g/njxZDNDqe/vF6iZzDja13JAXdIPqFabT+DrFyhO2YpC
VqLEBxUwVNHcSFhxXTPanIun6iG8CxwbyA75DPNlxSOchhWS+3X6mCYST6dabKj6UVCXbQKLON83
oqxm9uLABDn0nrkqjGC81qjBeMeJjyzXzO805JkgmsB1Y4A6sXiPtKg/mzDxnNp7dBw30vgHcAE8
6wM2xGeUuw9WKIaTcDCgjLtG3Exn90lQuZP8E2VpsZIMjWIbr+n8U3yEx4BQkY02WuG/0KCzINUT
SlMrWGOVfz0W3RdkvU/7W00Y+4RQbhtIUFX+ueKQRgFEmVq9QT64N9JywOY1uQlua+Az2OzFz2CS
2DN1Tzdu5HW4LDepHhLtKwLy9iLkoA9Zydfg1lkYupPmwg3Uw/Gb9ynC+CtEU/lPhAwfNVyc0yMt
3y9V/iWTtjDM+aIc8a5tAetTOVRDIQqDrdw5tqNmPcFohOC1wZhaC0eDhFJaZkgaLSYLi3HKJm+A
jtI9jegOMSeNtxR0c+5/kMLTl/QyHBn244xwUg4pkjWsPbcnUWGANfy9UnSL7X2rHbLzFtmCrrnx
K4ax+hr7YHCooky3Qj8vNqvuGyHufgKYsW/qceVX1YJ/TFkguZjy2mkQQybTl1Pj+MTcVaIqVvNM
Q6Fc+dYPjRvM/Gtq5Rl3fSZk+wqwv59d4bPTeta78HqumRIjIxb2UpHataloXKFmKZM3fMMdTsSb
oXmyOIzpA4U88EqI4ElNHNB813C/Puvc+/VhxnbCLJKXl9XjAQ0fp90gEysmS8FK6TdcCXEVnc+v
0h34B6AQuCLXZI9fH45VKWoaeNAeUGeh/UJLHgRo6MUFWKGWJJ4oogupsFLlu/63IUMww+7R4BgD
eCv2Bcsz9FGycAN4N6ry4ugtx4PwfrCMWh3u9NGZWY880jq4B77xdO+lnNeOGyjGmYXF8MMaEAai
CjpcpQBdUFna9neqM4Lvx2m4Oyn9vZeylQy5Edzi5G1fg6RVRQOHJ8CyM4sleUAdCZ0osoyidwzl
3JDdujU/TC7GcpH7icmEfqHbyVW7KiYDOUvHoFRsBHQq+4rm6ncnyaoG3xNvJr3Eo/mGk+F1ax2U
BaYhE9JXJagGg3l/YEwhGZftAg9Ose4DY7tCGTqvgUV3oVmKWgOVVhoH/t915D1jA5Rt4ZaxOOxp
Z4mb4FGR3w4UaKrcUmb4B/v4eeK+GvUGLttBxPHTyyU16XhUPThHbs7tSc4hgwGSbhKwPbwZ6Wl1
L4pagmfEdtGqe7XJkT1fqEBoWlmKYZGOWa8+KxJprTKRxmxsw5ieEVRssiwNitrKdLLhYcSe0o4G
WN8VVNdB9B89GoMu6vXEqXdYE+kyO/A5pEHwjer02ZaWjWXdeLyPCynoJx4FsXHE8HeOYTtbOFdS
hn6O728oNC90h8BCcn9krDuPxawCBvSKXpg5x/H8hEijodN6vqerEdIdmNPSjueHSNhSNgmPHY5Y
mvchM3LMSvdUa73573YqmqtNeZHA6SmDdBuWy+tXn4LI+NeJCvBn8+oQk5CAu3v6/x3iT4yxemHk
xJNGRgc2TTB9lyyRNX/7XGb7hadss3ru+m3WnsOMZ1AZAP9wRR87hj9Gv+/f51x3RSQGQyuxybob
5/SES5gwCsZh2rKGIPhN+0bAWTl13FglLcpWRG17URyLveB+ZwYU4eYFNf4+BJwRDWLk9rnUIIdx
JsQU9jCeMQCkezASvb+SGhwXJ3us+ZCrcozHjLjyMHzkOUNyxAga55Ami6JKx42LtWsLPx7Kv/+D
wEuybgVL0SYklmotXLg4L3wM//HPqrRMz/zMRbPHUmOmPl+Sl4CSRa8wtXsxCPuK9f4PFSAeKZNe
PQ8kCqhWDBD7BznZ0bjZlRZUmV7gS9Z/RFIsmuZK6YcHnC16PRxAisOmDxB5+nObPerDYAlemmdb
D4waA2wk14sWxk7bT3R2uul+WKmVDbDSQ0iJFXalrhz+sYP49e+u3bFbugPIT6ZwKaGyAXQnuG1N
WEPPmHPGOn/jfyazZ+pn6abPDohWFrZhifM9ywKwbdEHZOglfmaQIIYwXrCqtydp1NGGoXaIoT8o
553Yi6D4y/qooQ+dGsg0/wij/Tu0BsAlOX7IvTD8XDccCMqJ9w9jfjguJvXQo5P9CpkyRGS6csl3
c++n9gsM5BVOvgELoWxoaSGgKyDLl0/gWB6SpUfKws9q7JnobtAex2I9My/2Kg6zc+AIA7OPzQDv
2FZiWH1nvR1CNhuoIlGUz54/l6ghQ6MYMH1gXO0yawcJjn8EhmsgaCydbcOvtQ6bqJ5xD8KBQwNQ
A755KkcFBSZBdn9i7M6YehdSaKFe9KnITHEezNgYbff3CAzxnEg8CtuVcfTjl8dwW5WbKcwTuHCO
d2jvdZ7Jr+GAO8qx22qWRiKvfcoqm92Oo9d59+mhJZ/VUGazswKaDJiXhvzwTi3oKP9atpnfmNXP
XKP4vFW8Cc4CMnFIRob6stLy3jO4igC8mDAPc34vwpzsQxaGsPoQskyTZcE59rUBGGzSeCuWCbTc
uGsMtdpo7nLQe1pvFSO5ipenuSbNyK3lYS/3cYIBmGXVG77/mh+x2/y6/7KZsWW3/01OUUV/K4Oa
D0/i/lykFmLk/j0AZZMHLXQVswlTEae9JQbMpPviadQcbOFrZwoJISdG//2JPkgkb5tQOz0HgkTW
Gkcv6W/SG9oiA0+ELk1QbUCQnIotNQx8m6B4f+HWS3AIhCpVBCBhUGWmIQn3JJzASD6pCNXn4+Oi
dY4IC6C5abyoaMJMznrWy4vJ+LbDfvYFv2KdzWQ2oWb8UdtximZV5BTuN4Vl/UqrrIioq4C+MhdR
w7q3BAxDxDjjHfianlUnVV0WFd50yPexjcg0ir3GAam/KLs1xBc2GWZI53SllXnnZ8PZmrNsJvNx
8x/iycFsv+vNBWPBJuuyILfDwVla9wDpU0zJ1mznSEJKLATCqvW7ItT/INpXEGf/3hIIjlt4IQ3E
3DL/3HVK+Oc9z1L/sCsyGi37blAPzLL2xlflhNh0wdHEf0P6JgQiz2phqabGyDHXjH2DNcBWEvtW
NSB5r8YYKpRqeUUcsQwF59ASup6a21WSQq+mjGRrCs6QkGMzIerYr+z1LPhfDPpRNvY1V8fmyK+4
YS/utMGjTlOlx5hD7lBam7NhN482hqN2nHDb08qPFjCcQJdT63Tt0Z7PEYl0Qt4e1FhIc4+WM4l3
hBMRjuCwquRZ1dkk0bdYaNWdvq/I4IMnIIXfsvPMw3+fUIpfXznGufxCd/7o1Yziv6VYAH6zw2FV
FPhkF53XYZJrIykefyYTiBnqTWN5HFzwu/2niZ+k4o2vdoOMsboAFUqMBC41uyezRMBs7ts6l54Q
uenY8KYrAvF5rDra4P7OC0z3i1aTVkX0/7A9xTJjIxsKQFJPTwRm36mceVlSjNDwp/x9nZlohVjQ
ptWKd0bpQ4soianTJhidoLLWOHAuzoqTNbyhteCZYQownqOfdmRMhf2sODFDg2I2KPY7EaAv+mMc
/uGCGtioSvTK8yPUb0uXcZh23gdVNlYSaKX6+7kunGUXd0EhdtUCjgfNTqTgPFPAMgnN/0Gf74PN
hWpqqQa8ZBmLrkoQqkj6HHgawMAtwZV9y9q4vCJjI7WZbOldSy9tb6t4jkueFYtk6kz0kFUOKhMc
YQ2wsKhpLUkbyJd0nDNZU8ze714vi3TK9qXj8grnHxD14nsxQ/wgQnqgniweF31pTnpOcWrCd55X
WXcKom14ny2hhImBDasf2rmzO9Y2fKu0lG+IZmga4JjFm2Ire9A8ckt1Pb2kPXzPpKp6IahRYgru
NF/q6DvSO7sHLcNH7dHKgS60+f7XGBlxUi3iO1W+Sz2L6sKYGpYFJB5LJypbHUjlpImX/5fiqsJY
M2vlqO1krkqJB0UAemDP4Fb3bZbTe0gVynxfnAJRj9L1LYLoMkCvi12qGgwguPxzU8UCOTgtHvSP
Qo7Z7t0vWSpgKts0NxzWwMx8BXHsiBPjMGM5TKQiFCwgpeGb4UjRYcHFOj4TKNEQCzAMV1OZcRnz
89grQI8hrn15nLEdVBDZy7M4BayTHeQRbO7LpSMexg0r6DIYhwCgKXe2cxca3FYuN2uGzw/o5YX2
zOZ0jKgEG9TNkJH/vGJH44aiqrjr8JuA+pqP1VbQylg7bNGHhDKCyPWWqNSlH1PBmO+8KcZH2vfr
47zqFc9B+HKc8+UlU//VS7kR/5yYpUfS5EcrLv6DZE0VeiuAhQP+hSzzkt3Xm/il37gJU8SaavK3
Q6HXhywlZIR0HdoUxkZgRHGA51pfGP9PSbuwM5RatneOrZ5z0nSb0y4EmCWnJmiZwqi+LaAwB6ru
3NN0KPvEi6Z4//24B1907rx5zGcoFLFhbHnihpCezgAIlWq7Mbwn7JPYWLG334vnrVMpcZpYpkRC
fJUnpq1WGhLEp/a47/nCP5f4XBW6QiLnIE4xzIXAHXipd75KGwDDZRXxpM737ApCxP6i6Ml5/ynz
Pl7XZUnCGNSh8JOdY8Nv2yjV9jMaMF4WE9w+tW4CIcNzOhUdowWrULHNlUHKbV/EHZliB+/RkCHg
XCst/MGFB8w8QyawmY3Xpk2c2MLfgyNpRIX0Smftb9/4leaun4sv26n/OGLA7yRoVNQpIuAY7Uqh
Nri2UMa6+byDUNea0oCikfES0nyfNV0feB18kHlvhgg2MrA59aIfcRZPy9d0+TXOBtWbIdGjjvfT
6xIgwkLSF4DkuINktpYNTQYZZpeA/hev7Q5MqcZjoeJ4M5Ii7OcjwcuUfmonfR4G+hXHXNE1zBZ3
e/gPqGEmuM3HnBCj86lavVN0tt8bHnNy7hqlM19WgGC5Qq/yFPfMLYKLFuAlljl3uE/lZnwe7MOh
3qKLUL3fjMD2aC6kpw2gsrQ6Jgj4DhkZvnmYQsxJRQwqr4gi2goSPMkmxmyPf49ztUxSb5dajIx7
V5e5Y0lBj1pLFK2HkN3YH0hS5N8bkQoOZ4su99XD4P0AO0mMVkrmXOjlKGQ+GPltmhLwhhAHyPKP
3Kw9w79JyRExKaIvgSkXOIHXrRYbA7xPUDxg/1F9SLPTv72SEGkeu9Ggu4mJPGclK5yO/8JNKy2s
s7j1OVT29a0ASUUUPytIUMKstjKSSHdag6eV5PWIPlbY4DKBwX2zlZvItU90o/nfBmaMEZplmO/+
Vih21SbhLENoGz4FZwrMJMeTZz2WhLpOfxUbIl9ac+xH8hSNzgNYggTT03jwTreC9xiBEUCFy9Db
/xOaaF587OOEs67vxCbfBWfEOKkqih3CJxcJynsS7m7pz9nrlFp/NnCi2+qO5N2+NJm3paedGavr
rFMcll4ZR2oDZTQYpl0sx0PnrsVoxYgE6th6g6YPEnExz5AZt8j87MKoSO0Rie8KlGuiOosC4DmU
LGVHcXVuVZh/udCS8tfXlPzTD47l8nr1ng8SJ8PpMcVMSP1aNaIe8S29Kf1Vy5LEJ5x/voyY3uaJ
/eoUwLf5U34f8oH0wKIPFQ+nki/9z4vCeClI85+ZsQj6FcFya54rtunRjsC2Dy95SdB7OEjEdhdh
z7suJ/VrUngnUSpq0rb2V0QvNs7QO0b7rt/N3tT+0OIi+cGLA+eOiAx4+F1ixscPsx9+lKQz2jPh
ItQ0MlnpYv28cqdlDZdfWsTKKO13stmjxj2dvBXlPeklBoU52ls7Oj87jJawmiFTD/t10zJAcv1D
wcj+zXQrO3nRLHBBKkeFo5ObDo1bThrjmz8S+G0UvzGc5bdyIoXZJ2AobKJGwU00d0qHczrrhRmm
wLmlY6uVte2OVr+9RtHljXc+URPjmQOyXXp16x+yLFPKSTi/ic8u1yH0Fpl8lx2XGTtLo96iktp3
9zxQk9MXjl3KmDngBapgVJseEfTDdPNe6Z1gPRitp9GjhPnxAVoRMrszQ+griCZV49hd41dN59K0
lqwmmVsLevazDCFprxnEICllYgArdiZIGulD14SF7xfhm1wk77hwgxeZz6sFZl1k8YgtGM1sGman
jD0sdOKA2PIQgZvyEwsdN7kCPjOYLIhGjUnbGfJKfu/2qNX5VtwE9IXC+mNPOrQH3IDDaZdeV+K5
ZHSwEI6RT0K7ELspAlfiSKfsFj95EmfwZnJY2iRO4hIouOear33WIAmBxMy3IWnkG6pPXGuxrk8h
o8y64R80cSE11VPrhCymIz0v1hpc2MAapZ5fnUqgqB6MKjO9dg/1jp2mczQiHiRcZ9Eva5VzQC7c
kJYETYy/b8oY5d9rsLiZqhAi3VaaZzAU1rGUHQEwV5QsqUMpb/4ZgdycGeKs69495rtPvryFpf0x
cnWYnqFbSn8RUqR/0x2egH49pHWxGZ8l1KbfZH7ifCRuLF4I1vf8LhKrJmh0toKo+89V4TCVXUzl
cw7blJtVDz9NhrctV28M2H9Q9T5yzs5f9KxO1kFYGQd2ZAZHrkQTZRy793ybEVLzto6GKNKjZ+Vs
1sYrDt98Jo2IpaY5RJkYnq49aM74jKux/5G9Xc/LWp5n1308W8XGJwo2vH2f4YmcnBsU1Qywzd6A
3jXAV9n9M3A9dwblYeko5kkFfHs/n/K3k2VY9iTJlZLizV4rhA6OMbHyR5yQ1YctX+TpsDIvhwRX
v68qQICdrZH7n32VZzvSVkReS07j0NWp9q9H+lS3+dGyaLY3peiz9RDNkvgTCgf9KHDZSP7+Ofs9
r5MYDJFaHfMCea7kPLhzBQ2tUI+x1k6ysRQqwefW1ws3qiVeyUSPZ6k4wKW4eKnRDrQvdXtwnABq
pJu9VAa3rtsrt3TC5ruHof+eCaeVjfpg4xA93T/unbUjLttTOWZ7g58a9/51qL6Ck9F6RJ2/EbBP
egVbpQJd6USdo2e9loVib0EzbFzyW2Lis+xoPFePRSFOfuVctGRQdtsnYLFlsNGYLbb6yfn3crK2
UVD4Yf42nF3xeHvqZ/pdJIhTsjhCmAzocX9nZN7VWC1eDERLCHtkyey3zXuRda1FwbgSypL3CyeK
T8O3Xl3lDEe099KgO2wtdiAQVIGwfls8jDjwSLwZmDX+gG9fQQTJmYmXxTe1BWf5So1IaPn5nHNP
t/KQ7z24XiCmV/kRG6cnJlACbyVRUvYXsZeyhYtOSxbDrAgjGcxhV5CYj4tNmHsePYWzqKojO4sU
WmG5NnXrA+5rTBRv4SlmQauHgahIZ4r2iy3aYhuDTEZWRgNpRZlvLLfIbdurlZLVcgu410nqISPi
Cd16pbDWhKxlfWsMsIe3tHCUl11phDfG8luxyIG9QsfFtw9x9wki+7BYBpm6fYoi5qLZ+3ZuFPHR
DezPnnDRHIgyl9U+V3tzGVKEUzKox1k7HW8wel2Wr4mFnKE+KsTJoZuJtD8It03xKX0uZ+Qque6x
y+yfHgbiK1wDwIqUsp88gJUhEMkC0Nc1j15BbA/El7htP+y2CQRChYm3z2bI6SbrzM4januRJWyr
D7V03S/Qw6lgYAvWx7rXDAd5kBqVKwWZUvaDlfN7dZuKBYM2cBNw4AuJlsM3n1IoSpBKCtGAD7+T
mmatK68AD1RB9osGatHP0cf4JBoP65vu4jZBd4UN5cdE4RD/+/fTx2YrZXfzyq7nzcIxD7a4C61u
Vm5rtEoiO+5Xwj9brPR12KaB5RLFR/bU/p84ALNw5rBu2h+AibAzEhTtGJkBRoCt/F/hmaIRD1S6
4eGNngW4e+smDSnUQY8RWOw+GjJHFgWqdJCEW/CjQWpAg9ufHmlibT8SpjpqEcrlY8iB+cdnmc/h
pJ2aNjsaNfwYTM+8nZUHy3aAq2z1fQ3BuqqAuiBa1Oln+fcKvom2ozILOzUpyzc9UBSmn6X6w0ec
ukW6laSa14chYo7I+dpiPtH513THF70YAWevRwBPY3BZqKi421gjyvoUf5RhFTJ/pYOhJRM6+K5X
zV1KTvDBDCTPJEEnA2fVzW5DxQ5a2/fxLTrPEw903jC8tKsvoQKXcV6cvwHJMBSk8ihb/JJfzGXx
JmtJ7KBLi/bamwvQzzBK+4dbNxnsCfxqxfuaeAz2BmdZsSKJHogc00hROCqI/sRg06KHqHwcK0LL
1Fkq7jcZjnbfOosReqRTxzxnd3i8xQARH8FzulLB2up5xR8uybxBmq0mazPtcVPDemEtxFXmZpYS
1YoQQCgmPEIO+YUisCVWW2ZDoYK9RaXVRAewdh5EO+btZpX12Ur+nMrjrXAF45HpnytMlIaYhuSM
SMoUYVoGBSHpxbcVKJmqNvHLC1rsoanHV6Um8YIZmFkGhdA5l0pfaEHQ1Q6FtODlarO7QpuXq/xM
npub9Ja0Ok7naPUzmnENV46apOfzbi4UZzG06NB8SVYHkYVDS2RL9vKdtUEJ04wmVcsX2MOUkrZY
a6UaZrroL9zEgUmURM49u+Ez1R4Ap5AT2O0IWy+0i3J5h4m/wbND4R0xubfVsPLywsAdi/nSPcyE
rszCP9NT0F+QtiNwVa9Qr7auDYiYsaU+t4O19td3H8nnfIv3WF0M8bUYhq072k9PnRqwRZBdHYS+
I1NDPTuTsLjJzeOurB+0eljEvfo/KrkRURlOqstIPsNArR5PJpiDIvHQZi82JU9dIU4Lcif0+gS9
l6zj+E/gM2AbCnfExdZif79VKdLfHQ0/p9TiYTjfXHR8xpl5wb6YGXH6nvc4eBPQEsyrVzgGIuFX
4/1qD1OY1Ey+yahCwuSx3sIsH45qPZmcOnYlAK2k7qdJDD35wo0cZvIlRFoti/iWKN+Yqz9whJST
f5eLkSS+vJ6p8E3YveAxBvy5LCV2hkcYpqw+oK/Sca+oRQZNkloLi81GZV4JJFApGl+Wz+nrxDRU
VNE6Dd89EmLqZ4aWEEVX7rKKGMVd09aZP8z0AVK4eRHJliYVTmRJN6rSyRmtgWDz8SCrgBKqbRfZ
EZDAjKDDjMGU+/j5G1XlWzs127M5eA/4EQqwk1j8/H549W6EjSsPuBRN7fCFzEKAOGSBKtfPliaB
Gv01RDv9Sh4rDTUWe8r4NwRvn4uMko21jrVvlhOivfD8B1w0AX1Raj5Pl8PVZdn4eIKGSektSPw4
OLxg99aLl9N2AQsrySz2V8xgjcYwnmuKGWepZPMjzymLw2J4Pn3k5+kKkcTWh9memuMOA67IQtCE
h8HcYXUiCUg/unUkKlqdVHOK4f8tfr/AmejULXDnezUf/J0949ZpbWbJxQ8ipr+6L2+Csitc/k4g
t3wZ9KHCmgzDGVgpNDct0WRloPjHNOrG7OKjbGcJRlTfNELy7n056fOB+N/3PvPlBorbLyZ4m00I
/OdaOeRpWGAmDKPPO6AmhGWBTZ5q+POYEWXYAe4LXiX1QMUZuvp9c5dk13Y3DSbi/Z8lJSInGMhM
2cSWzOko3gqBBgEZ46TzN4O+q8yB71oGzsck3eT1jRNB6LMG79ZX3mjsJTrbV7JcjfuZ0ZmE+NJf
Jc1kCL+EmpaIyebHTyF/FTCp0jajOA0q1n7hnv5qHe/Wz7YJqlBrl13W8ZBB1U/A2nI1LWpjHEUT
E+ENtXiCnkF2SphEKoftCwcN0L6REeKburgJyM5kMBlpOtYFAyZuCUs4435c/Q6pNg+DXMHyb8dN
rTufCKP443yiIg5QJK2j8pJwiki7t+F1ncYM6iz84GgV8x9Fi8ay1Ubt9XeBCrX3Fda3XRd1BWq3
y8uo39AI+JShscdyEPGU7EBNefOnoKpO2V3NR4ZS6F0waJFfBcsLXZ1LP+MnZ5X2Tfy+0sKDW8XY
z4J/G91s+2/Cllx3tg4egcvhEMo2DTDQsfZn74zq5aIGXS5TY8YjrXEWvNRxShc4vkk/1KcmED4M
ExtZRoDzL487L63OK8GqjGDU682dVpXaEOT6UK9xv4wordyWwAoSaR402M9LIrh8sb9shM3FCQqe
YACrril8SovUqALRMx+VV7925IHnZob9b6bg1vhNWdIWkxHm51GtVXWqasSHi5GaC11EAhyIGW6/
zs1GCn9xwSwI6mTxbSV3EDY9ln/cT9LfkhGAIZJ43kHxMsSzT5tP3dV0HgKEdNldeDa53dtRAjYe
qR5ev0Wvd24QzQ3kgx6DdKLEt3LZtYV/5Un29wnI2Q1eNFJEQOx9w2Wd+U8EEAtsJqNsyUF1y9G/
87tyHY+7/z8gF1jw0D1wdwJqMr7GpW1tZO82YyXDRKb87Qkhy0LL6qvJEJMte8WF+YopjykxeWsb
tRrXgfUWilZxk/TNqgv0QoTf7GNwDcuhSZvu5qtQDkpSYdzGs0CSmaG3H4djyf41bRfCxIYMB6/0
u+LJif8cfMNEfj2bfwXabrvQUb23x5AEgVS9+2eviFYjqs6Gqo0vyVjG0tndiRIJ6Axmr11XWNo7
XEpaTfj+GRT3efe8aeMaPYLvoOcNwrUb8trhyU/fNtYxjo/owN3Uj50CqGHSqFYGPyaTwG1mS0hP
8h6HjzMZVw2iHi/OcN4HWIvXYvw3xZspFBa+8mNIFqYXzWY+8nx3PzFLC1NlHuQGu2h8FAmCjjx4
1j4Pk9Zw0sDyKgEaTPMGpUsM4n/vNYTvqkvaNzCaDMq2Mj0iebQCOT/ugJh+6n8/UBB9j/MpMgLV
N3RR9M4BJACaFz+bls7+cyWIHl6b1xjCw8aQhNfOE7KqZCABbvJzDuTrTGo/GLg83+FEaw3p7ggv
YC12+RyaH9YgyCRlgLbNshUBQhC6tomkgBXyReNlJZ3JkkRND3oJCZxNzhr5Cv3sxXkZKSwqgvhC
OZZDsQwv4ZepAZ28QsXuJpIQvt8kI9rA7QrOe1UzqgRLyGtFxhF+4Rdnyyzl7KZyV0HPCzUDbBPZ
IHI+Lpc6CZoy7dUl4k+vnMiR6Bj1xtVe+QY6vNDZ0ixVyf1qOckGWzd89FAY+bHJBiyDfkv3I+CO
6Cgg8Ktxi32MG/4BRWwwZT2QW75UAqq3RadXvlkOg77FLn7I9v3FEI4gOmG1FYjOt9u3Si/zSqwe
MKWdlNjp4DCZq0LwGGMG0+wNA16lU9muU/X5otcJ6VgTrs4KflyuhqqTHhq0X84ukTkEeNQC2+EY
QkpAktFlidqU0oSNE5KYRWv+hVlTNs1JFq+UBDDHWQdFHxEsl0hkZ4Z9a84cebScZ1N00lkHz2kV
qi1K3BjAmunAqIMess+BCmYyyoZGRNWxordmzU3tvucYF1yMcJW5lsjohxnFSN3OpK2NpK5yIj8K
hX9L9YA4E15N6I9o4kvCY6rQD1MedXfKl7IumDphySMWUBEwfUMvaSzXV9JfZ1+4HaKyLw6k4Pff
V5Ye9y0MWU+RvJOKf5EcZ3OeF2oMxwy29tqiFMyhWF4HuMUwXnSY3dqa3mRR49QTyxgMbtxFGhle
8RqDENckpJJcwOaQ6Eyrc0r+1hrGaKN4wfk5GCgWGMCUAOELCRTmzZ/iPEfcXNpKDMRZCtUVCZJ0
ZEcjFL9dsQiaj2SnQmOQzowjceIRrc9C28oJjT3lxecw+HV6FNGDWQ0QfFwUala/kUGZr+Vocvl+
PpraXtgUoKXWQbOr4iYpI5WV1slFn5Oyp8UgpEoKDB7P3tAV66a30PNT8UGXGHh4atVcRll+L5Ej
+0M7TVCY+TU2f76syRAxKa2/bPGhOL8ah7/PX46qrGIr65eIaHUcCwNdy6VsLPDdWrU+bZDGnSeP
A/Fqj091woNxATXnqwnOwg2W2nxDWHUBwA4J+3rEGiLhXQTXqKjQnkQ1rtBRhYw7mZFlv46n+eyT
xMp8PcxkKe2m4hRkVDMA9/k/DJ3QAz5d1Vf6o7GiFBfakB6IgsvVDy3Rd2gZ4w9WRdnPiuVXd79z
as4FEpEgF7e3o/P9TLeh9QyHmGhFMjCJj5x7socve2KDdrgzKs5F8hODeoP+o9kzBM2jr7DNKYtt
CF5r8C2drGyTiSH0p25Hw8eqxcxebKZxqr6j2cDmKzmLGItgDJTJpXAOdb9kMjAC/JN1KgKjFcr4
ktJhYLNCapeaw+xhu3SmCbOHVrIOzYxS2LKtKTfxX1gB6Ais6a962R+hz/7zXQWcb6ZmZg23rPoO
aJTnEwYCxLFcAJl2/y476VnHNx6dFNDh4PDnX472GTue0VVgxS4l1cktTXgzHbySg6rehVOfUdep
6FQsEP8gLrkaIHl1N9GZndIaSHeK8v0CqZFf3w+WepGLhvxRWDeobNj3mRnjnahmeNO4od8QyI6K
m0CaP7cI3OnD1MeUbAU3ZuZ/+kzrxVo+XppUEqKeviwf1Et8clyAyUtk2xelAeKs90mZNAdm1NcU
IEI1CUEGcJnwmVapbEiaMYZdq/1ogn0VXkIwIJ5dRw4Gi5q8AUo0eHY3JA3R3CyBir6OXpjWqUTA
RzIbSHi8qzFEA3gWOrZK6UXnCISM3HzrrGa9QMRutgUTYtaolvnTHnQSc2p0MCklEOwkbmO4Qk2H
pVwWHGD9sGhuT/pXbkXDQxA9hyIQKwoJiw3bxd6n0t3WsIipBir5kUCm/BJ27XwS6SGbGfztFC1p
HVWJ9/PpnwAG7ai74nXWUsOJKWg9CJ/y4EAqjnrxomxgpgOIpfOg2GpNUSJkkEd/TFgkfS2beh0H
6grrMO4zidOvfa6K0r2t15WOQV8r8cJe1Flh56rUA2OTZG2Bxy+pgkuTYFin/xQDf7dDC5vgQEJ8
yfI9ld+6iwWx2JORMiyLYK1eCtw1P4ySF/3U1uNAlBpIcHjmziW282YL8KTFa1/q0rNgDkD+OAnb
lvHEoOpQZF+trzEzpl6cZTj+askrgiJt+BgoogYXE8aE7RY/jESucexvqT2AvZfGPR6gvEJZosRP
mXTC9y3IJzxaawWXgEL23TYKJ/BRDJrnJFXOM0kjqsvG7IP5mgLg6rrhYYf1Ze5/amwnt10hrdcr
tdE4iw5VojXObjmLBWV47BPEOnMF+8/GrQCsUbDVAo2IqMah3Oc/cdqJ46EHezt9AZbvPBLVtabE
0NBqDaAa5x76rdbBuQ5g3XCnESV/3lHGoOobw5aycOf1vx+Z7ZmCj0hsp7Nc0yRR5FGvrDTkNkbb
X9YcCJmjRPUw13ZEyjTjQR9kd/OccAJc9V5CHsYMbJ4xX3eJIKAFa5qunIU3zIBxtlFA/n9mXJMN
sQHH/g5B28Lq5INK2O0PZ38Py1CHbnz71VL8FTCPh27+5b/LW0KDX0R2G57IYfXosOJjU+bryCKu
z+CZ/171eRqi/k0P9UEI2f4bGMez/ol7hCaPj+l+TPsXTbYeS/jz8MxLPkESpJFedDRIZf1W9ZCq
t5T66HiwJvD4inleRKWRJk0WcA6P+wKCFMhJ3nA2RZoRe5jzdQAjyiZ19TXu7xxHLMsf79LKxWhJ
CSJPldnsXoKB2AQzs5H1oaCgCNm/YIwknRgz3NDcFMXfc6QA7QWuL+8oO0ugHFEZ4mHJPPrJJneF
seH+XJUMLadpuSNlZsCOO5tC1pxkp9NESERieDYgWJTo6igGvOWmxyJaaLYA83faQnT3BULfoBRS
gdIJa6Ji9dZgk2RAJYSLE1OnwQM8UeqTH/z0XOeJLKFW7fJa2TuIUaHzj9jNtXmTC9IiXuC5F6Bf
RE+zl0HwHEHNT/YB2/qZCyPX9cqI2vGZhnMMsAQJfYbhzNuLU1vYynOVf+oiF1mSIivQaNpy9R8m
usfaEMNeefnZXbfpzaWwjX3RbEjzShzXCFFox+MMDsRXuApYYnr/wLusaG8SIlF3f2epXptzDDfd
1HhCSWFFwy3JORE2Yb50plowaGbZnaceiziNuF6OzOcqw4bqheq2Q7y4Jv0rR/MzwNyapz92bzK+
1l0BgNnXhZsVZM2t0kZQZOXf+QzIrRCJ73rEbnc+7O+UggwsMf5IC+Y3sbxLelc7TiJ3SkCd2VxY
viTCeZQMlhtvlW7Hgob3jfdc9FHnmzVWnX1TnpIStUuJQApQ8ebYJOFbvfaOTo2SluH0sElv+u6L
lfuo3m5tMUkrl/F78sdDSvhzIBmosKm1RUhgtWdz7j6IqNXY70Bb79dp56wupI3D+SX9PjTDzqKc
25usw9fyAwxNKNoCiuKe4mgjjF9Y/imgs8kjNJHAR3bozVyCRLzfdhDiAKHAQdLtJo3/sE/ZwFoq
5IoYEUwxpcUe4xxpFZC6KIdFXhwPCIVjF8L6LXe2oSnru7q5oB9numBEK9hGG0j37Pah6MtREZ2j
6NtcpF0JORGcN/QkZ8E8ZAJSBSdOrpK+TrN7O/B5/d5fNhW6zFkMLdGfKjSjADuaLRaw3/mxx4kf
sFcmoqWutnuCb6kAieJwn+28GwoNpXCM6CvY7fisHJCmEW0FN4gde13ZtlnbaV4re24YHFMczhz3
eUz3T5YmrOk3eRxyu2q2QWiUzvLGC/o+Rz0ZkiNcxA/zv9I7DYg2AMUV1tRvXdqdcM5JOsElbO8P
Agb9QCUqqSTleCejfuMLckBbnb23KdckOlQLffQa0sZzrLF94MssfsWumR/speZfakjoMb2KSpuW
SbGOJqNbS7vLPIfDUEypZ8RCEpx0sRfNRJxpkaGFFuAIcEQWKN9P4gKvGBsBW23a+nW6jlmHz57b
gYDuErdXhHD4uw7ImL5putFqkEYcbe3k36Vcn8DtruFQdlOSgIuqDzoHRyboTZvYYfXDRv9MkJoi
PP74QS4Xiy6eAdPa2ClNM/j0CHabk526JtvGyYFaqS+P8gQ29PWZ/iYpITtGg+AHIYQ5Xfvbmu0W
4j3Xqg5GRDjeFVXu49OBilgkqBdlvRhVUtd4SxEhHwd869F87337OWlG3zMwRkSmgAY2OvNy0Sw+
8iyN9X7C7iJ9k8eYkuSqvE1cA1JIz6SELHJTbMQ1IMTPzxTv2fJ1+1PhwTdMO9V0hUQBw4VUNN+H
zGmiUH/xM8JmWtNeMTrrRc8QVQER9FahbRoTT0awvk/lVPxCIgsxgqXXh46sMC5Fs05ms9crocN3
Nv05jxrrcHJqV24tqRNUVlmiWeAe2s7m3lfdPz2rcd/8HC9Y2/vP0C8sG+w0poKFbNxyEOYCCaY7
xVUbVJCNP8WwggBhwdib778L134ejbtciUGIZtex/V1YPktF1PmHL+zMFn4KSij7j25zq3XW6snZ
x8cXhTL+iENTK8r32TVS6dVZ++MY38rET6dzzNgv7GwMfQPOutxzs3BBV6FpY5BpnNZzJfLM2lHm
oXXhe96gZ2rat+FAPQb0HeYucDj3kuBv0QPhQRjRGYTXPBu0H9KkjELCozrUlamYDwmwpguHxNvl
RISVlTwh29RmtcBnqyhkvA3hCgZzIRHIz3ICeQ/qZUcPIAaYfTX46L9tBuekZwqHjHJsGxmXCv1F
iD4m1cS+kJ1Coxoouj1+HDW4s8WfqmvVzObwx7XIDfuNigHAq3BCFhlsP8Kq5SZTazQciLZ0ZPJX
EYJaBQ6aJn29VGwqJhOLyAy0JYVIYF/MD9lnywXnjIC5XHIsz230KD3qpI7MPFgfHFjp3qqnf8bD
Smy37SRBCXZgo0bycg/SW7/hps87gN5cljBwtPio/aAFISF85pAFJG8S3tfqrbIFgpmWmDH8k/yz
rviNGPs9293Bdt8R8O0uTggsobo/pj4drTR+18KVl7OYC9WyjrVC7WaL9FLtgsE8EB/M6MLfy6Cg
9BTOpHMQW8cdCT1GVyONUtz9DjcJv213qbIcNlgpx8rjL6OE1HsgXPhqYiruf5TBXRzre3MVCESE
Jr4SkBki9EyUA/d/FBCsCr56xP6rjl+SDrbKpka+JEfk/nxWmuVNwNyh+qJs5s/xsIuKhFs4cfZ8
9Ky1aUIa2lAMI1hKgEAlJ122FekV2tb73z/cNCovQSw8+35P3Wg+x2ImIhKhmKtqUte4wDz/hZFe
DeaJ/4+p53UPx+kT5NdTSjD+wfyX0gvA9WvQiy/TrgdI2GmdR2dEZELxHSm1Mz8uXqs/K5KL1U7e
XT1kD56yU0K+fHyaeJIq8uySe+FUrtu5S0Vq/ZekWzAY/DbZw6DWhWuFQySsi9Xq8CWHMN0knFnI
9tKnQQab33hRU96ymciOyQx89YPK01DlCxSvTFR6GvybYB4jKkTauWaHwwgejMpxk6ZTaS/N0WVO
xvKfzItVDLkC5M9R9EgoS/64xsBHQ1MNu6VHe9AC3HgDTICXyDV1kNbQws5LQysUKAD/XhXVRIC1
OW/RfhcGV5HSiqkSLL1BCrCAVPnKzX8HSI8comHFM5qh5bjCrVyvxHdIJTYtUpf3pomvJ4k8Rkub
0J1QWLy1NGEchOuZ0fuuyqrgGehdRcFHqZMv+1XFJtDushhCc0soQyve4vVDgeh5Ttw8Yp0S2A+d
hUZnEoFBEiRnmRSsa8sWbk4PhLr4+KVg8OTQmsjz8g4xLp8h27P11zHP+x9OemtvLYczvWF+J454
D5AAcFezvQF779sy2ec8582EDTGGOQn1x7S/PMel2+ZcadbkNNMf2lW/Kd9RmQvfYEmcIV0A/Q/A
IAWJQlZKldiIE+Y1ZZdki4KZ0hIuSamwylJYtZqGpY6qgmPdBgHSA9p79YLucmhBgctTWR/1UJAZ
Nzvtefk0GKs0iJC0w472SisV6p/rdc6Q8YIGuI6P6gpDq8rBhVur8Bk4GqlMD6AVjqUMH1JU28xW
uXXl6RJfNkC4f+qsYAlPfwcwCrCda3asEOHSkR8nibvLfzbgxMfY0Bpb95aC3VnWpk9uXh4TCWvi
g1eY0i/yviTRDKo49HF4Zr6efTHTQNenRwbG7Tpfw6HMbREdEYEDlwlSuoXX1Dmdy2Bb2V5azJvL
VcHQIrZ/ZOaQ4ieLm129y8KgpE9sQJZpMAA/JFjZWoHK5f7LjCHtNqUP72smVH0X6BKcRAy2tmx5
UTqaRSS9zEFXk3gU3KpqFxCxWBDP2TDPddv02xeRWHrpiR4x8G6c+JyjDAYlKvWfu08VzTEWMfTB
wDQ2yJ0hv7yFJznPGxDDiZ6ZTYs8Jb4xylb1G1UQf/h7GJ0+Ah8HeWE6fyydwN3NHuQlNt835I4N
DzUCy/lVu0zVxivmVgdXrCHY5zata2L44OPh9NheVDbYaWe2b53FTr3ipuPJyzAEcdeJlirkTM2c
Z36K3HFnfrn1d6J4Q+td2zD7633ct46mw+Tud/fyJOhYj8JsoWFXxlnOZePfbypyTmw/OtUA2QlO
utZ6cqx23CDbX0xzMl+fiMEYypgJSjT4mqssKLfA2fkDGuprB7pdLKe5MBkI2S11oWyODIWsSM8I
FDw2AJV9zmfvJftpN3AfxhA4vJNlbnNedUU12PpC4P7jhpu+G+co4o4iSgPywmOabpos2Yrqrte8
eMG+igTf/OuLke1whNUMRI4hLGdJSW/pCWSFMPWq6zqWwfjQcMqGAxLj5BeOnKCeVlf4db/jZ1l+
/FUsHX0VWZ3hkndZy5NniGF8a6s77UMEVGLKPVPqUAeR3lbqeaK17LvWu/q/35xF7A5IQ2DpTSyH
H6XYL/tnsavGs92zjyI/iWuSbYvxOQ7WZD3o8X0veNiX+WvPW+yiB3W4kgOfjN2e4N/SxoWgWuQS
9Hs/S6upMvKtvQsapy4l7FZafnzHmDuTwnRRuTulBE8QQRPew4GSjSjeqomcpik/A+8SAyvOcaFP
icM+BQRVBU+cZpMGaVnvhQSyZtxyBvd2ctGj1wGr+P3eyse8N8Wyy0MDq2UCxlBavZLWqoI6XALm
TVrJpSOGN+En/UzgY3NTAfUk4EqpjawZLsgtO6IiYLDqVud4TzSRQeMpSw19g+RdwKGKdVYGujsX
A9teqRdJxkYFIvOCiJtHvaOS2ycZ/MCcIvHAzi9HAYwYTVu+XEfdzHPhHxjEOGNM1ly8kCgar0zZ
NS0pYkQzlTNeUT00aUjWNSWc2c15CAINffSas8I5IF+zMPU4+0fZTwacQOeoU85G4Qn5s+cj2udG
m6N+5GlFCjJkoILN91EXvJZZJmxcI8mu1c2fCpACyDa/9RfzBKw8Gm5q+9SbAoyDbjV/EBOmb23H
cCG2Rl/iFe/8Bdp448jFkodqMfyjLbImXviBtUVR7bOmS4OLXtkpSu4VUAAgRConWL4nB8keTYVe
Y/bI1wHtqx1GMxsZIulmG1K+nReMJGAu2GMGW3/zvosJNb6ZbHAIW4Ni0TArEV7gCcHjKBHcEJL6
rNRoeJbohBr0DIfnupq978bbUkv8efk2+qnEud/1/iHyy4P/HmUNY0iWe7kesqmGFZx4NTWSPdq+
FeLBcBP0s/MctERtDWD1CE4YHyy+G9T37tHtAkdYngtYu2OXLsv5CpjuPO4gb6rOnz8zSVEX8BZq
SV822rrT3Otw0svBKcnusGKzbilbqkABCEHlJfrMK0hyha9Vs8CPpyS33rxQfwpwxGTp/vDONPMe
OgsK9ja6Kuw+TtfmgrRa1OP1LstVRT6+qKjBv/YuJMyRkO7mM3wqWKNwRSW/Y4k/+m3jSoX/Tv2z
hq73UayEq7wTlxJSWw7WTpOsxZAgGci32sacN1xmu2jt/1J5XPll6i1JyGp4RsZoJE9dTSp2N3J5
lzkOH2yVkC8zjI/0plvdjnfqJlgTq+xplwUBAkT2rjn9M/dqaT5SNOMeo8szS7LJWi3qKg6xwLAV
at88GGRynlZ4uahDsX6KiIUhBRNyWQ3Y7AgcLpAJcKgwwUQcIDpUcNinAuIY0d9TPf3pGyPfRMWq
d7biAi3d5JfJ1UQ2FKXcbzjLjXRm/Dm8Lz8jr4nb47cjJh/Lgh6/cHjg1AOwxePnW9bMAcTcrqxK
IQHA7t/pqpvYwZNJygIXbBEO/CCv0GJUpFzj+PCcsEJfAirNlIHEydWz2BIGSE7l4BeKL8kstGhs
gvx4aqxDAj469G78EIMCehqxXqIRNS3FPtlbF5pWA69qcIt4nJQ2Rxk3PS80mr5iwfSLh8JiMReh
T/aAspxXrWzMk7UlcSrM+DPos8AcTgNaDQm3cQojBIHghe0hL7DzfvmL7ZikYNnarCEAG6tDzsbA
MSHcMv5igIc7eQMppt8GCH8WRArTq/doUpeGUpbRTN0ImFtr8sq7IzkvLLiChGDnHlIU3dMYK+Rt
qUhzfqnBuZB4gzq67KS2OR+j615cO/8+zKkHPhRLAjfGWDR/AcQW5AWa4yup9QOAMFEA9/+hJ/aA
OzCJyTqbgZzx/KdSHwPR0ZAilQZFRrPHkm6NdtkLQ6W+TWXKI8j7cIxT0VwM534biBlEWTeF9efE
H9/hbDZJpxjbqEwT4NK94qNDYyWqJKYT2QcQDlUkM/ZuGrlGQ7plRNEiU9d3QrUeZiGeVhYy2WjM
Fvy7RKORvhtMZvqwjcv5qR7678qymy3E37smE8zlI47qXEcgc1LgQEz5aKe/uqVH/N66rEboYvMF
ypZBQS22ZovmydWlM/Yfs8R5CNQAtIK7ciSjnNlhHvUe3QTqntnMSMqFPoriTU303OH9h5wBHNqi
hNKI2LY+XXIlfV8OACPi5flLczcIA/dKYxd8Yx9v6JF7Tgu1JFaJyD+pNaEa5DtRRhpMRZmpKl9y
7Dt6vLgUONj/wIE9k+wHWrsmmXqTkXdQ0oTJPebauYgi3WKrw3ITpmjPDkmNO7wndJWm02OWnLMh
9cA/U6zxml0WEwotUAzCxYJyMBdHj/4MfCM94F78pnHbjgue8RkqswzJhNmOrEEedGoAl71jHcXi
bmFeJTk+bI6ND3E8gKXuImyqlFL0UsLksTdf/hRwJ4BW789rhPVpIEpFi4pBNHC7FqAa36w26XHP
VPZsFfbmbuQN+Ib0bPX0F0hZUSvNfcSTYS0Eb9eSeMEQn1v9uC6hyVrH0vt2BoGEq5+H6HgJMmH/
RS5Z5wvRayTaQWqg3XgA9u5WW8wFCddIz18kMLvL7qNbrsHebkgsQK93GOSpaqXvEZpoRoGMuR/Y
emU4H9EiEt19DpSDIeJsvA043ZW0cMxEt64aJ/WbWgSxLOHvfLVM+TYytob5tAu6ZOZVb+4Bd/Ea
NlJ2zlRnXwjeeuRC9qXcuAIdq6Bt++XJtWvoTFEW9Yp1wXW176A8RRRE0nQ/EMMG7vbFGUnOHjQD
5F5KA3/hNpNzdNg7XgiVduwMrl8J7G3tg5Db0DTLFsxmLSIZg30eKYfJ0whp0P03pV5edlhez5qU
n7B48roq78r5mo14GUU+L+QUILIjXd51nu7wBhIazmRr9/vVj4hdHcaFqrTwjD47n1ZFdy4CEl5J
y0hJjMNcDd4czJGmF2SxJx6d3rGTQPZulYAuDch39a94wevHYgG0wFojVL4NaBNBnm/JvmhAVtlB
I8zmGSWc1sS6qNdPpHVT8JqQ6Q1G5q9cGTnxMTqTbqcve1pgpn65iIt8pmrONJKpLxIQxYuUwHMQ
JZ3cfO1ryP9Eii84XZS/CDyvctMrtloQzys2z1V823WFo+FQN8X2BPT3OE820Ql+gRsinU5oA+H9
klyJp+fnpPvYDmezlnoIGAklOdUNaujRg+edsXOCvVjJ1uhK2UgEo82tXK/mW/7zUzqZAPuYWXIk
iOsQaNrYjY+5QzZ9MLogWDC9NlVlN29t0ai+qUWDVfHW50hKuLOv1vii4Si+Qxk4p6+Bm1GJxPXu
/GPCg7NH/43p+947vFDx0wdG+07OahJjHiEioTzSa/sAOYGcqLO19qRMdJBzFA7wVa9VGv7gh0Jl
jFAsoAECFbKmkOr4Gdg84Pa9Slfjc+JjnNDgSKFijxeltUTuuV0TqsWu0uj0rZGRi/TtdyJzYisU
wxGNZddcy1TT8qdO3/Q6Cni5oXFociLkCATYjhY0X3HJubCKd4qkoCELjxStP7Byf/FiluYGhppS
hTiFrvQ0C6O4iDVW89muipXm1IcqsGDX03Hvr6dSradkLW6GJMIXvEhAj3xq75IRrIX5380HOBH+
5eZwG9rltFGQA8N9q9gZSZ3eWooKGkF86D6Yqjl3TGgQUvVWo4bApDX7T9UCZ7HXY8hzG30JkaUE
rrmNW8Z0x0N/Nbmx3uReVvshtywJq5jqU2OgyuCjl9N8hC5U6pMuvRFltWNxkgqUIBN0ow0I/Xoe
nqRTaYSkVlZ0/QE8MD3eK92dUZes7tljU4vZZbDsE0fUYCbVaRUVg9xJHUnbFwyms9nU9Z4QJ7K0
bUNRbtwVOFkMxi+HB0Xk7e4Edp/+pYJvzVSoxjwjINWno330oBQ/MtIJFoK8kQKFiKvBdrH5Pt1Z
4ZMIPiWVbAhsZ2t+8cACwG3rHo+g5UzllsDk7BrmrDSasr3iV+lx8WbmhIwEEUZAHIzUEuvFFoCI
lHWEDRlaByojc5VyJgVSu/VX3+IsGMPKwzZCP70EJtMOnKh67AwozA0Q1nZExC4kN+dJf5WNfRo5
tWa8vC22QZv5xPnhHASSANbk/+yzNwgx8NRRzFtU2nMcd8POLkkhg5cmyu7i3lqkuXZXxiZUTqC+
R5MmGuvImVL5jYYRx1FKNJb8s3I4QzBBbIdr6DIHkeKv6CZWPYlw09Y/ZuGeESNplYOxKQNpk/RI
xXGcSOJwD0MDGoyyeLceXiVCj6aMSMvjj4nLiekmx0UzwpzNKGElfbNrFaeUD4SMTE0lf0j8MRIv
Pq4lRdmdq8PMmqqxmQC21M4DZi0YWhjWuUxdLRHhBMxMi3acLBtlMD22Z115qgYSn6hzetEDiqyr
cbwUJ/+fM7QdfaZJefMVMA/BcDnKFBv0vhCe5ZqUNir3ceJJngQSWtAPTlRuSn82BeZDFOAFSzD/
r1+fo+TrT24NrS2tHVpSASANrXAm0byYzubThLw7tYurvXbOj8z2/xVemi2JR/tS+YyDjVycQmT5
v4TT//5IrCaEDHDBlE2d2/Z35vso7lN/SYDIXXpveRq1VE4B3MAYJgW6NgxZMDCHce6BxQgzJa85
Fm+YE5OL0rPgglzq3gMErPoqgkrWsR8yhkapllOsYu4pBOFlE1817uQhblP9/tiW/aI4+94Y5W4o
3iev0J3/Eog1ZbOmxrjWtx1h7fMn3LwlrZOgoIKYigXvlCWlm8JquyK/ogQHarhRVT5vhW9D3B11
kPuBvwcFWSoz5FHmoRdKQh7kuSou/ST6eCq3TTo2oUUeafSli/dkNtNDHliOuXByv+QjOSmR+T8v
EWkf8ysI635hxOe3DyUKhlxHcWoWqFqhLWp38Cfu2Qvklsi1L3gUBRo8WR7uXztvZOtJqXDmSJLV
8Z1FIxnCzfEogE8lJhEtp2NGo4HtFbmzRMKlsU9OK7b7PB2hCr4Xafn5yl2Ng/24T2j80aYVAb+Z
XHx5Js93RyLvQ8jMV6spUAqulncPoT8VOEyEeOKYfUMx9nTOp6iCFGtbBcd4rupJqx88DGry/pBg
Pmfs11eEb2ehBjo9A2/rnaxaP/0/Hu9yZ4N7M0CTBdr97Be77s+bEDhLTDwPhnceYUbpTIGm1FVr
K28IUEPKxe0NxHAKlIlaQRZekoYmjHpJyCPT7y8aNK90gjz6W75SPFgbNJ7cSrsK5iUZrRPPG1MG
oZOkeALUNLm7tdiHR3T4m+l29I6m9jTRhJClWjVez84yN2Jr5z9eLjtycC8/nJQt645HAi7kKEm/
29jogQ3wk8drvuI0zm3H+SkARHG4yopmQWfYoemloo/WJJLEX+xnRUQb8ZXlRSrece5h3qgPm0kE
Oq2OfBHd+x5Gd5lh9KZZEQbmQ6tR9+AilmxUjt74e2E8+ZpfHu1W5Bkinu2KrjrspQO4P/xzVsTh
GPWG9V8o0JCGrEGFWiOfCj3NxFGzf745E3XNEqxrhgScjYxHAyhuzWv7SaeofbqmggF/sGVuuPty
cwxkx5z6djTHgNL0+rGyBh7THZ47Cn5INPMCbrEs4cI4EVkb7uWVmyMmkh7vZviYAdcDr956nr+v
9Lj12vRKDuhv9eis0OxgCno1evnWb24lL1ta7l5GP/iWY7NiBgoZvydirbODYdWIHcRnxjIuXtY2
OSrDiQyL7Bhn0Hxrc3bkznXIvFl3GeJ3t4MZ7diIIDn1uQdKMebMP3W54OIJhlTmO8kjo8uKdCkp
jCcit3eZJl5YukwT5j4NOO+6c2pJsSKCCSpRDkdQIcATuTXYD5nvtWDskZ7TJ8i6Fie1eq8egG7t
3IMcpYSSQmXsvdowQwpVG31FwINwR4FXJ51nkwstYoyrNl4qEPPymKxiUx15zP+AfPDbjMEuCBpR
5YxiK3RuccxcT+3e2yqvIn5nxAvbcOdiWuAb0xN7P4/Mc0qxF6i8uUGeF/JpzPwnPbV6UaTmkGR+
PjmSwjgXr34g+DF1Yg+Krq9ilNdFiMTDvFVJXkH1pC+G/e00WdB7a45BP8bd9IswJCyGw/3VdXd+
UE3mryAtMEddjJdEh3P3p2kKP459klBWlZs/Wxsj99QZ9PfEjm/CIxbG7HefK4r6UA3sEKcH8pDW
WuwDKD3qk2m5XCucG2ENCryaKSRzs+v92xH0FBQiMCb4GxVmDuY+MWJG7ZNe5HnB5MtUxUHuqHfu
+46kDFAKLTyvjBExi0+e/tnEqmSv7glrbYkSrcD12maLfr7+qVozALpfCvlwHa+jAXNAFquUkMN6
8Lqg3X/nzN80R9l614ESUey3LQ88Hf725RC7SHlr0Ay+dJ/Y3ep2D8JaEiCIBLQ/tZO0D3UENrGW
bPc1bwnMGOnL1ktUmfzHfiFrc5sF12jY/giEikbM+OOwma5kKcGgtrO3phySD3JoDsKhkaCM5Rpm
gCfDEehstbZEIPfdkMIwCCk+KCAkV0AdobHTo0/uk5nPs8mqUz6pYVneG1WNHJnesCfVVDoZlVCY
UEYZiQp87OK1LH3a9ob2p7sgKjKx/UC4VumNqS6U3TJx7cIdF2K+vI0Up6Dk/yf8i5W6Qd067k69
jVRbxltGe/iQA+KcVvFDZ3sm0uFPbaxXm8V/ZZ5lAUsTsy7IM6QpD4WGWIvw1SOvRM1DoBI7dC3I
SSy+7E/pN5Mju6/BSUrxMJ5B+n9pt9wlKI/E7NVen1cHLT7VYPGU2IpKauAvLyfJcD0f+6oKVVtP
l4CqlWb8p6+qogcwYlUNbY5mAGsa/gDJVZqBuxP7cO7Q/ls1eJV/O+zyLrOK1oT6dzEX33kfClix
MdrYLmaYz/PX6JEJXApiKA1tNfIwB7EL+SPCHlu3ASgSTpggInkvF8FHB+NnzqzXc+6M3EH6Oh1g
bG7jchx9rgDIBumr3DYq7K3ewB+NExU0uG92Rs/czVzk0ccdaCuAxUYXnnwsJXhMDXRdozO7PYBs
512vsJNMQ1AkEgJ3Uzf7DiEK5o1VfBTvyrYt0YGM56SZosRBAC9vXOnEczKQnQTd5YkWM7B0lLFQ
yuC6h+9CDHABuwtJkRG23I9I4WMSpdE59c4ugvKXHdcl7p+AEiS3Pksi056mJN2oU2JNzchXsyLh
0vO9wVZxQnXqtcipj4RntycHHzo/gIayPDMFLFEIzBoViP8S7HzCTInYsHMUbkhnp1GGY27cwB+r
dxr/ASHTTmDL6ctf3I+oLXVMn9zfpXVlvz/xoBlOf3U7dADo5RDJ7QPGXYQXczIygSzzwStTtJll
0QKKXAQZEWMO29g4r6M10g6UNRACjM4H0gsspm+BKnuVw68wUxXo3Vyffnq+Z1yJKmfHDcQCF98I
vBmewIDQOMOvGHpEJi0JH58CSMQwXAiA8b+lo4ywey8uWX5Tog2cFJSlEs9tCK2HnVPAQSw5/vwd
g9H+n5nX7DxCUROWBG2bSqJS/f4oMYh3n7UzJs1eOmjwMSf2Eg0SyoSEUj9BFvSsQWzA56PyszEK
fYpSPk7YgTseOn/0N1VBxutq0yrG54FptQGV0mbYkS1ZiUjhBwLnQihKqeI3bzqgbtF3dzbDQRI1
AtXsRpF3v1N3Q11mqRCHd0oU4vlZSU+DsTHqoJwWTwuHJclOGL0hAEBSDp9aYq/G2hIvxYbBeAzT
fCpgE736Iy/i32gT/4z9g6il82US6UWdMLEzY03Qk7stxcKRyijjM0JUlMuK+toT6UhAibGSd1GI
H+d9Jp+ij3nraCyZjk5n6jLinnEjDdBF3U5yVbWbZbgvjgWU+3LQ4j2UHDudvjBIHoQgiLDmwd7X
2CCsqWQ2vJyS+AVfL2i+fYvDAUElKbWT1fsBM+qse/m1nkgEgdq+9TU3x70HetSZnZBhrHzV90pX
Eis+adyedf1FWUrNryvCKhCuwWMsStmHlCq9TVFB2H9+/3ptH+kJRhsfxxusElnxxMvpoPgwgpIQ
bah9CV3UFdgptwvbZ8/iQrhI8shbAnkMBLpJI4hj0YDoDgfI83RpIngHsIhFwiWiwtukMRNER2PI
zEYofWrP7VAI0uLDpoV/zFcueSerFe92sTc3PgCUeZsQ1TaTPRsXf0na7zFc11mBvI5eR7hAYduJ
Piwwwoj4hBpo+xmJBlLCqt9hzupzdvVQliViqKDJ51tACwtDBThOvUO7HrdaE81M2AOnBr0SrgRc
+aBekKsGfI6mzsf2SsSR7gHCLHWhNOJVjfrfl2BnJ0sLoJxcXhjQGPutIzq8gfJmGL4Be+i+i8sk
3pj5xGfjaQOn1MqIAIo0ECdPGVtSP3oxGRXbsV261FrD1tordPWmZY3HmPC+NSbXOuIDIMH24Xda
sUyvGnjJKoO4QoTr0aYMkxWuSsIBXeWoM/zQr/+FYMHmbUpWvO3W0Z1D35am0n1aYrZeSNrBNjZ/
gSVt6g/Fwowk2NoAmZq49K9KK+o5NCk1PRlE20egbe1S0jDubHZxdehMP/9S+pDvfzepmpKDw9a2
WKnqrZixEYOaY6e+3YIelTjsh7SKoVKkM4f9p7se7C6j4twZ1+P//VVc2x3gDMNJhZSSYI5fTTya
sjkHs2+wS+GISxq2+GM6+B8MQr4+ml6zlf0Hq3PoVfXpIMxRT70oRSaxb/PyRLLaq3N/duWLzJeI
IYj5CxjRNgc0V8Jio7+qP0xul4d3Y3mEQpAdGUHv5hW3rMlDweJMFaZfvZ6TMkpRnYfy/iH9AmJm
/WppgpAiSMbt13VNMIezM/XfvptCm+pQFu7fk81o3PKCGbW4fID3spdAUCaULqmWNzxACqvwCa5z
uisHCRKGo+zVnU006xOadRlhuPoRfe8iRXhodIgvEq09zZ3vEIpP6c7c65+VyGvhecZNLEW4y4Fm
1BEJa1214KiwS6u/8fYm2+wpHDt2Fl9/4c305x4uD2eAHBtVl57s0pGdTebsRjiI6I3eTfmiD11X
yiWvb8Ox8kycteqh0OZWJp9y5UknIwN8tFPCBM4Sl5O3sy+5Orl1PxoxW7XEbhfOlzFJ4u8XZNkW
kOJfebJa8dLHSicpTa+wM0Wle/m1Y5nEpG8z9Nj82hj4jmR/NX6xcDF4Y3MMyjEF2CJ5Raazfc7G
XfkoKIGqLtl7pWDM9iAeqsX5B4HEopdxbyiWmQHPKtlT3kWepIU13CzBRcVHkOSuaOaBQpGtMbb6
enVjSmSJ+GPn+j6dauDb7FjWSOzq8d9J2ayXLLBTRNee/6ud1008BsHHsuEJjsx1+F12SQB3KlIn
wHLarAnEJZuKge5BVBmn4wGpJGOS9JxLvtZInmTRQK7QBL1Vkm9qK0ag06q5AsLH+rz7tNPEzIya
Y4KQcqF7HutR4yShYl6AqtrHVN3uT06rXQLztqyjta+eNaGcbe6sI5Vv5YW/y6O7xdGqd3z0HLLu
Hh1s8e68eWWRqDMUrUAVP6OlFqBNqFYXJdP5OGRyNCIHsNb90LKWYWWVyqYvBDt0omUt3hoM8SGw
mCtOk7q0SX1WwvD9vZ5CvlKaFA8nHG6GVmX/JkB/1nuHrR1dkk2OCxDV8++HbZRdG3oJPYreZNCy
I0KTKJIx3vx4lgpuULP8fOM3lkCiF4jgrAqI2J8F7ek6KBj6sT3nmbYly1fSAbaUXANI7wCCIxoF
AeZNzPDNkp+JJXD1hZpv99RigT2ytwemH/hfddhPw8+MMOaxaFbYzNoGk7QKchSwfu4sp3mplP0S
bWBoDc09zWryl4lBaWUw/2I3Jy53kvuVb3IcO4AVioGP2xZLSPTOyaQJzL3/ErucsyAr25vrmKhf
KJ3o+J7mdJHG5661vRpFcop/JalnDemq861sjhmiFjzE4m41ZGYajFnTq4SJ+fOMiQSM7yaYOPcB
5fly+0mndEUQQ+68qScA+8jagt4FENWFz2RiSZuqHnOG5HgwdPn0uPe01+iB2uqq/501Lzm2voel
F+L06IlhVYFskOCG/LzSrNfnC8Ve7Xy+kZ4HEOhRmQ3TwOMvmsef0CDsCHUXUfnZFhPkjc+JElPl
yF7thatzjZW+u9Dv7959xtG47Mrsm/55dvxR2wh8tdOd0Vr166YxfXRQMj1KBS9JCtmgYXy6hejZ
MMM36kSpE2RwJbxF8nAYmG7KvU/csVG+1GNdogzeElSoZrg+9OoiNcn5EIUNVInV76v0QKaIQtjC
ebP4lLnJR1KYrp7SO6B4c7R5b968fSdHMBb+UU8YoV6Qv+AjGk6W9s8+de2QgS7h2OYKCtS5aDxk
609/a5ZiFhWxexlRoteiGwNi39oipm9bzyxUZFkpArKn+EUgMkj3HQAY4yuMrQSZBJCrRgXd7WYT
YxlTH/FrOm3h02fGbEC66GqbWvdvZamtWRursnweG1bVWx4Dk44ki1icuqrPiTreOJVMKTcZkF26
liQms7YLc2nl5dzygB2Ws8DGWYXscwU6e2QybkNb/w8ZFnA4dW0xTcNQ6g94VEw+TH2g+JLfXdk1
SZw+6V2/1p9DveBlfwUxBWe5uQ6/PqWmkxg6z3WzA0jQeFXdNj77ikwCJkWTiU87wQ1abAOyAS8W
wIo3wcOOq4B1G4aMdY1fWZb7iRAr59ns3t9vvj0BjweJncdN5e9wfCnDjMn7r5J/VhBL7E4nmeAZ
g6WY8o3VGExW+pSvvNX3ccp20C7OBmzjNC/gb7andKG4yR/gpQDlHO1NU5bxAesSztzgEdiwps0u
6Xw8y1dBzZ+9zz0qeyu7ln1GiOxd4Sl9LhDWzFgZEehgv7JJHHgapZCCklPPpRDZtEc592zBtKj4
nV4pGzH79sBZRD9cJXnrIipKcYjnpUNOP3Arhm/lIvcpDFU2js0eHALdiofK9yvn+V+tg/QONWX5
//Df0TrZzhPSVVq6FEmh9G1D3LN1UeMQ+hXOO0nQSHSElqaP1DBMl3DrblzjkTCuFVGmBeooVI0V
vq8Eqf17ryOuYHK1YwbeJs8gR/63iKtDFRHhKAtGUndfAhR0SNudlni6PBKnTX2HcAqknvWSX8qb
OvZnntenQjplflw40i5DQtUkVb3c7JsdduS6uEjxvttJMBzigHMWsd+G2HGsvfDGVUEF+fBon8vP
RTy55YYeUlrLHudR31eaoHKY8vFcJoBOqxfdAMK3/OJwFSuJR7hhcbjvd9Q+6/xcRY2Ks26fiHsA
Q8aYQGoaMggr9Nln/9FXUR1tuaJHmKRhaBtXAg+gRmfIQoQ/NYkEtQzB8YfSZFy5w1Qo/35X7P2F
xRyj3qencof2pR4JZCt7gWosnHnBha+e535d3O4Jy8ZYjyeCmxOaDbkpXpdE/kjza96p7JHNS08s
YktZ7VyBzcrzXjaB5K/NR7JrykmAQeORLsRVs1UzzZv7zi8FA92PLIjdKorsDVe1yUCDMgQZ5P1Y
EWrdTsf6OFc2mMsYBL4Fm3qa0H94H44nVe90/utn7E8jfmJn8aMUNaNX2DP3cGRoVld4VaHsld/s
y/yJBFO+3T6bBTMwjb/JP+E9oxRUiunxuS7XVBfcTEBEWkj1Jz31NsBI1ro2suFKj6NejcK+Xi/v
LG5sHZcIyFc0f1Pptw1tE7EQoE/VrCwNlwZosUxnNOSqwraEXYkMt+ZypRfqV9/VcQBGy3N68QZq
OyYkM7Ws4PMNVsbRa31VaA5UK11mhF5sBzLqo40sokAVKnuqwIJO8wWW1Rv0aRiE4KjImx6PpEzb
T36KxN0Xm21r+8P/UG15Q/VHUrG9Kz5NH+462rVS6S2VHZpIBF1kxhefyDtAIdZQddGWO9yiYzG2
Vyhjdo1Ja6eq22vUJY82CNOcI0CSxYICNmjH9dt7SzmkXTjVRsRFqDFXKFQKLNQoP5xYnKLVWtUv
EolfxZnbAeLQzBbRtRzBc9brv/H80YEpPb8pJAmtZaAZ/9EipfQgrFsKNWPMzjulbnaCWXqMDBx8
iZDmtQA60Vb9kek7kn0otOmd6L1CYdJASroL4e/SIiSJSdE2bccAlcDrFHl+VN9jBpWUndCd7Nyz
T5j1lQ6nUJn4IDaFFkp+M/qnGBpd44UiCnNRKoOJ+KHVItUlf7xfpcX99+peOUsNTIloeWnlTRzH
Bu7UaJ3fc61Ppyef7Xlwt7YO6//WGPpAPdG41Q+Pa0SjzD7WwAWhSlGRJp0dlqcXkdOyvRoptivY
IiCgo0/i4HUewsxmNw68ZCIx0tmMeZXDAEQDBz4OE0RIhr+v071FzIe36/+zN1k5vC/Di0saE9fC
GhwVXF5qyPjAv0o3O9WimQKohkx9+pJskK1XaY2c9JIcJ0R6+2ZiDDacUeswNiFF5+apwdTAmpgj
m3VeKT0POI5vpdEiDJY85gT5zw5ic2T01palF5TD7c2T2EkMmZ5LquY0kvemj0yzbhiyVHjhW8CV
KfzufJl+7QKKZ2HKpPhaBIgIkrqrsy5T1TatOz+0gEmkKDb2Z34YHztkNH9OkkpZ9EqowEZNkmUM
cbi3o62keBsErxEURrVMHbDh9POhHvapotROd7MX+XiHWVNWZVUJrg7UaTIY/fifscUt1+PJHod/
Gu/tyAwfjWuqsCLthg5EecwqFfNrpCjEhgA6a4LFcBZ+3LN3LydmUsESoiA6lpS+8pDIv2bQxXaq
uGKVq2VNz7jCnCq/+aQVsBE+GgmkekYH1MiDHYDE7cHLlZ4n3KCchKi3UcqBEZ/AqiNuwWL/VPKz
JmNLrDbn7uAb8kl0Dg9X72pAH7XTW8ksKxbmOpVoHnf3H4i++Y0DY1/YivrXzzIwiUBrzRQQxZvq
8wQaBX/brcol+wgl/UlDZeyuKvTN5eUzlq3d33z3pITetOfrhSxeqQ5CvNq9lh1kjVf5xRwc4j7r
RIv5dHksc5L647MgQGLqopFAMzhDEj5ebnr7pdR6dOJu+5IXZ54V+APvertRhXy7PYIiAFalGMgL
mIDVYB295UvYlnT0GPhQefW56wS9Y38/2gybQMF03djuw9CBPCS6NC8FoEs+a0cFGVZhCJ9kcCYF
nOpPaQxTiI2kFOlGRi91KCa8s/UnoB9+uM33yKeLuNIGFCRWfSFnh7XXeDLVjFoBumd2LW5Jd46d
g0ewIcsIbanVU9wECTVo0AdDpqhbuqNJgWTcMl7JV5lKJHFoA0mb/Dyix8BiA5R7WUtTcc99Ugx2
nvRxyFNQxUiJPVf6HmVaVQQF9DmoApW97Ef/sE6TIUPGq/utx/wosTGlTB0Wp5yqI/Rdgt1P8Vc/
r+mboGL/MqE6gAxlOk6DZ+CR2MveU/twnMd6qwgUf5qOHwfG1MoSX+oqXvvll0E5+uxL76GTWLPb
JBG8PR7bnFjp4Xt5HJ6Wp7LrT1ph2aueSXEjVMLvTRQa8omgRsAELXKJpjodDLnfSwiWOAJ/Nr1y
KulprjHFAzk5yFxC+vNGRwqVp5jeuayXcRMu8DThGjMHgiH7ub2Qo0iyfks8RWp38NwdfFO/BiXM
HZu0bUoFWHRhs4QxJN8J6fYowsBjJrD3pVFEQmpDeM01rxZGhnLw5U5YwhH1hrmU5JmvH4ItGslO
b8bB2ljatFXDhQ7uLrp5oa7brnd+JMrIvpIK+yQKOGPGYLWnR28cPm6/DIw6Q2qeSREv2wuq09E2
XbYEPVj41fua84NHEq1H62Boe3/LldtzTY/hPMftnd3U/w7oEnbnZKbYvoA9Z4X3J+a28e9oMi1Z
nCwvmkjHJEXLHleO7RdEq8t04SBeXnIfAaljEpIRQW00//jDn5k3YQBDc4AudYTXxLRs5YFPEPEa
tDRz8GWSNt86JJ4WIrtHG66ziIrOAsCVawZYwWQimd2ADhxmWGuoHPUad37RZ4HyBshCBATpGiTb
6kz0Hd/RLr8m6W0RPmEqeIUtBldX9NNAFbadrBfTHsJkEtZmwcC+TRX8Lsg8ZdhlCxre5DucOSP2
NAD96VdxSyRUhiW5H4vN8iHq7ZFpbAr81y270xCn7qDwwVOPoTwv/FabEF/f0+ZtxKtRtqLGgbgK
cQeL7L+rfZ4fcTS9Q+uf51OY9vLqogdIaHA0brVYuqiP7+AdCVVJsxe2LsEihIKa/3QFhC/NonE8
Uf6bcKKPd4eOtEkbIVHZnM0XYPSe9MJcSt08J3JR5JBvvilQ54etVPXu7xJL2ZyAUvrMz60XfeSu
+zjbb4G83WAQ8RM5a+3BJ6+3x/8e2gSPKAJz2zUDVun12dqoO7ll7UFNKoqY+5Uer4cAq8QzG4xS
thdYnpQ6+lD1n8GwYpxJ0shc0Ss4dUH893S9m1TQRaWyUH2y5qq4o7G+7uWBDKdRTje+M60AF/dJ
X8+EGW6Z72DT9qLfgv/XmoQlZxHulGqcKfYTkylzbDYGfXaHi9G3ZuLXTiULfgQ/F4JsUozdWn/T
zfJ+vTZIlxMB5xA7EMZYUe3G3nQ+RoT3B0bvElW8xR3NAXKEVWHdWCR9zVcx8Dt0FEnQavex8DqC
XNKYfjGP5dwqGP4rXPpNYBEmJp8KRrcksPjwzRUEKIoYQLXONGzgqqrf/MCkAIXFSpVlGGvmpYie
l743fz/yCHgqiXsRB61S6D7LbeJ10FOrEhtIffhkVGG+HnsdDkp9MaV0Q00VTCiY/hYbbNKTA6Mt
3r+jvndFt5MeDRmxWZeKdvu0K2kIH8hZOy6hEJUvM/rmIOHOKd1UvEGVzm3VPb7ZcCZrEoFzCyZg
tUgEYuvPq10ADcm3plJuQ1ij1KEpz/fjXJsjU3CA+eXLC+OwDASMbUz/dTlFDv5PBcShzlhRlpTd
Rwy0PdcYqZTfr+O9nFCwCQYMN3C5C0b3IKATx+oI5nJF0w9A7a3ebomgvnJixcug3m/RnJZrl7O3
Q6O1LHxgjQDA5DtktZPHW9y+wOLKdaLx2/qIIDtxwetawxKYmyW9Xwc+gpeoQpXG5GVmFVgI2fDi
yCzraLoZR5On8YpsicLuq7dpuW5gjRxirJw4jX6YiYvhL+q/Nj67PFSRyqkO5VxzkG/2PImybCEv
EEHjAqYAITAxyl4TMDuSrpfEyf8LUgNiXx54riEJ9hsfS49DC2cF94jlOUTw/gYEO/uAVqkr4mh9
jk/qwNRERvXgyCtOAysTa9r+UVTcVJ8XTeBubKVVX20GvMFYcpddw1CLqdp5a724hTblmeJ39Lpk
cOvlSWILhMoQHWXrnRSQF7a9zj5mMzr8HsbFaLllPHhN5bJB/cVK2dE2TCOQcjTrcVtstqQeVcyT
V8dM9Nh7kdRl5fgcJHHKo4RbaN5Yjfs2KJKiHg8B3VUe4uEPIRSAXTLJu55c+OYVLa7yp2AJ2H4T
FGIHMNcNXDab4SQ1nnjIi0/Zoh8QRmTq/QLczSYCZ+Mh7DkaHn/Bl1GNG9N86ptsqDSwJqtT3NNs
b9b+mJ9NHkLejuUeCZJL/rNT33qJB+XYDsiN9DZSAqrzD5P30LYsSp2ucQNarqtXIVLRjkI3jiHZ
+55dSVy92BUE3Ifxyuf8G13CUOW9UT42uImlccef4R/BqPmmrrx47X/6bXU+drmhl5LCkKtKRomg
2YIXtcwGApOM/j0UIHCEJfxqBtuH4XL8jJ5zMQj7n4pp19qtSeBYPtiAfRHaRXTEp3xZWNqpoZK0
OWz33V46tmnSOtuIhlxY2YE12BeoIMPfZ8PEhgxSTPNdwMkOlIUHrPNj9tpNUawsxlcIXlL1vDXA
gD7D3IHweHeA7WvlHvJFv2jI00yA/0nTYucHRSi1Ne0rzNl/Cf6LwOBzSV7ykT8zhUF3ylzhhQel
NW1wQVdEk4zBdTEweKSIHkfYRu1PnIPOeZ+nMhjt+ka6R5op5QaIxCg4oK6wCZ6tGMpLfoHd8IhC
ZVj+hEjg5Osjq5XV/movEH/meV+tZh3x3APadGH+Q9BLDngzSEYP3kIegyBYBkeQKnfqGCB7OV0P
yZbJ83Oa5QBVqnWHl318Z0zozNSCxb+zljgIiQ93ZJtGrwCri55+V6b3lgX55fd3K+wg5UmiW1Ch
E45YoneACVdpKt5W1g7gU08jKL4gW0S5KPT9MNOXGrhMQx6CJKlfuDsuonR4NrrDBgZCKpz7cXXL
CGFTkbolyWyXSHtPl4YV1AcQORToAOiMtbU2XoU/VlOtKBKc6a5M8jRV2Z8aZ8zMroTXB3xnBHmW
nIhqNiBz/qK6hndubpbSVMIJfBXj31hsl+TTy0ka5tTWeiTq7FFf7F4AifvyB5P4mX7eNwt82ZDv
Ykki8Wpr+Sg3cuSDMxTePm+Wbiw66jspLpzbgeXGPZUAKlRcq1VijxbYH0hlxxjn09iiOHoqeWo4
CTpG1DeCCN+AkEuF3QVvNJqIWi9vawdKeW9H/o7v9l8awj1hcs5B4HwkqpFAOw4Me8tq1x0tZeXf
vopKFeK0bA9ajWVKIdApsEtg5fZYQ76GFQ4mDaQubP41mQxOP2x0KTUgUQvXep1qSY3zUE548SUH
la0j62a4NuegQaOb4RsifN0xZ+SlpC5msCM54++ps3pnXxXkgEdZv4PxVRgAw4apelEkHqpC/E+6
XJrxSSlJlBzQJL2w73FD5T3sD+VZxUWXKQ8QKTRaQlLC9jfL0igmemq5Gd5DLngBtEdJcF6ZjLqZ
ckIqKkkpKIQTNCAr3QoKnfrQSB42jdjnROEWOvDxakfmzD8t/ZsitU2/0iCFWEmY6EJPSZ+8zvXb
R7ow01MM+2JcNTSUBj2Ax5E3lc7RADKqN/Ay2j+9mD3xZsCQsgdVX13BYlpVmFTSWsfsZWQLebiu
Nv/LU6ep1eESTuxMUIMYBcymK47dwFXKwnfNKxY4xBLbXSRenCSP1/zqb82f+cXDksmhBhP45ruL
8NpKiY8XzXCa4i5XBJYGwqyR4z/yT3idd60E8InHOoOWsV/2Snp909w6la5MkQ6QwuCLEpEoGx0l
OEnByWjbqR3++nSfj9iHjV3Dppvdurhj6UEXKlH5cOoyI7NDPV3ApdS6BBRMYWYBtTMO5UMETwBW
AFsgTrjPm4onpdHgMn1I2nmY/WnLDYOrsXJH4h3Jcebc1JSYKb/FwkFkwDm6NPsWnn1yV/Eu7XuW
rZn9WrI7tgtxZ4sC2nFLGXH67nca2wX6uLMqcUA8pIan7SxlFGIwXRJ/qsgGIWBb+vS9SJIbv5TD
6+XpxhwCRP0Jd2rxVfv5ALXPShpQMB/gco8fH+xae4dgvXS3x7yLJhuTfalA7b0XmEWX05/5j4zT
b1OaTxfnhBss8BJ84rdoFBpFb1/MwcNiUkPDY84FcdpK6K2YNynK9/KUliWPjFKlnTScU0YCcGuV
4T0pOOAJSzM37g6powJRP0MoZz/s6L5TPbUs4gixEFj25Liam+2NOZBfgEsGniGaNixGSDDa0mO4
ev4fIEAHi75NFf2Zfddu3tH3FgtbbznCKXi3aRJqR0/rboGbPf/zdnDrf2noXL3uRWpLxPTHujgn
RUjiHx1cmPx21GPqcZhVgpEfUyrcNy/jSOMPkyaPc8y9NsOSueuSKW3Se/ptfby6mzPHEth2qUrf
WWFJoIL5813pII6Qk3IWNLHxZcVIbFZVviL9S3GsYrmyYlIhouK0VACoWpRMpYXUV3FFYpM6Irli
TwCajfT/jyD4KuYDZ8CiQRIeAIQm3k0CgreFFhM1H9wEc0S0uHK7tCDI2KWQZABAGQ4JQX7wSumq
e5Yg++JOO90dXxGSyDiAYCkrBbPBbUecFzK6CPAY6MZ0VVSwud6628pmxkvkgcCz5sANXLDzQxpR
itH1MDGarX+k90MW7YdcALpm58O/bzN8gAAMCQVdJyQDZCmxaCQeMo1QR0No+6pGtKHcHIhkyBud
ZEvxVEmq+8Bd2i3Qpbjp+acKf64YuvbFtHkOpuN7xZ+rz05RcBKc+8LwqXbOMVfUgWf6E499CxDI
k+GLcnDmeqYfeDdJcJOBYkKJ/9+OyEAak0rxJzavGzV3fWNtlH2jVc511rU4xCKJsZhCUxuXnePh
XQ0uX9y1SUlbbfriEcbyxi0kp5gxX9EgVq4ZURCaLMf9JbWj46aaKmyuxSexR/G9wo8MohnepVVa
rqlnV1p20b1myePdHu6A3JH18QrWtx9RJHqdjyHXppOzGkITbauWe0tdEydIK1FZNf3unZOz9+PP
ekB7LuhtrDM5Q5PxqJQYcG91iLIJheUg5JYcs5zTsqydjmWhB1cu9ZgnZzeN1roqOyOEJghcvOtn
uL2GDSElZqAzgo76XqGzaydRjRdNJOiK1iUnFCLKdi9jG3mmrYCxjDyGXJiPfPwQeAp/13KCj5tM
TNxOmK7H2TnB9IZyHFaPHq53toSR/5gaVJjEUaC4CwWR1V5rmrqAQAvM/kThaPV6obdnuzJcw9Gi
6b0+Kdbmh8KSOkjHaAzEpS/LJx1JsEogvdUdoMpVKPfjnSyTZf3B+4X1Q52EGgALkZmmIPXkJVfF
it7ghiv2Q7N1rzkZxYcMOfBm4HEMVrPCN/vwwvKgBMar7W6dHPMXRNhJO4lMQXzTBaWFXn2K0uuM
S+CUDy6TZxqLFu4qrJa5dNl3hrrazpFnACW3UyJKZWQDtGu7GSlQipxZaGWCq2eOjEE2DZIRPrU8
DURGkglu/CPhi0r1CmCju0mhSc+9AdMP7wVjJ8qQS+NopxVWQ5x48RKA+cagJNM7ab/EEmQx3glj
ji1SYMqfMTYMCKmON1zRRVSHrkGY2uZN8EN4i3lkMduQhZFpgVD0z35Ge+Ib+X/jgQYFL595y/Wx
MEOkkip7EhvlV6kTeh2njsJhzSOP6SNtP+Qvh6ktanzOt1m7+bGrWWSwg6lGES1Jt2blXIWay5R2
nx3atNXgigPFFcsNqG5NOlvL2h0IKJdpvuFd+xnvic9AUVtLFrNxd+toHyeY/9YA2WVWg1vVw8Bf
taIvw1CeQqXsysmi/YExPToySSuSdGR/9sLWjVf1WnfYK2wodUz3vUbWgu5NMeEyhEC73izOrj5r
bhL2hppnGp0F+g00CVKzHO0G3MypmIbqx4VBNUxUu91au8sn6aWRbrPfF3ogvTKsZEffq7ANt5Wz
U2J8zqf1JP8EXOVJOCV8AvtAye3MXdEmzsnTeu3Z5q0Jv6M2S6BD3Ol2yAQce1rrTG+qge3UINOh
R0s7Tl/KHP7oL2viA5nyv10qy84v0vCDzHVvQjtZHtfKrIjjOzcY5VHlO3nI5fgQkkFl1kff19pR
2JUE9Qr0ttTqAq5ig2hocAZ2gQdlZzj51t7y5osukugup8OG6/sKD27MMXDzl7BuYMHyHUbLP19O
obh4Z41Pfi63kTqcO/k3aj/GBfKCemq0YID+MhhO8suDlh2a2FFy1sb+J4r17yqgAYhejhj1EWg+
2g9axb3VItUyx0OhHDA0Nf9sczOVXfewqAmlAxuuk1l0/h1tW5Eld+2xVqLhO1QEX7jYzQEOf+9l
hkYAfLydGRJy39BBzgqrksZQl0XKmfLHVkAEXpbDeN6zh7ATf66AHAQAvKByoEEr+iNcn1UdJGHi
nHvqyH5TULt8t/rCayoEzlOxdXbW1pI1fZDZ5pZJLlsvSg+nM0FO84IL8RZltxFCa6LbmwrZDmIB
lLONpdh4eRPWSCe5EsJUXkB6rHS6O05mBK9R6v/XECMgQtAeNiz+OfyV7QVYQqZYQDh/cHPE6X+v
VgVEVvdozT2KMsTg5GhCLLuP1l+yzrloQNutODFgYo8LCGmScK3fkqfqaaWBqeyWwIW57N24DbKJ
r6jzfPlqsFnYzaZDupnJxplR8SlcBlQd1iHuPqcUNMNXp7z4gR0iYdRdIRRln/Y2GDSDeigaWZyP
RWI5JJh2H5E7ZsWYsQ6bK8Yq/tkHR+7bf7AbkDq+z6VEFTa7KS3HTPoTU4SZRMZU+bhDjX0jUDWP
ECeGacRwMTjP/sms3uTAwao7we4DKkIXJWp57mSdZiRHe4dfl5T9h+6ng3nMtYsZxzu6lZFY+hu2
gs6obN5iNl7EFUmNqqfbl2P5UJdprl6qTdtc1sIOlNQ9bxc8EtYjbhqKFiK1Z4N11AmeSuogt4G7
WPfYR1+Ib3Oxjlt8M5uMAQ7r+iNcrFBa+IpVSmBf3VrUqj+7+orTCJUEsb6n5RVNAobHrNVlgyAd
FLqpLuFg+HD4BktKwf67vuG8ezU0a/s3K4qhZnD6bdyCI/ypJ6SKJKB39JkfiG8Ccdf6oAtfAQV4
KNZuKMWp0Iy0ldyfv6iD2suoD4zKj1ph4tXT5KQDj+TPRIRauTcHr6NafdvUZVXO/QeeHch78J3y
xxwNIL27PlRTSTQVTJtWYCRwEnF+7w+HrU+l/v0fctOIXHcmZwU50YLdlcTpNzEfSH5TyWhAHiAX
fqCWcJizkfRPliV/YQr4eu5ODrDdFxcG4omyZX7mFNXkQtO6THJTIj/uqwa87WplQDs/8wRkOiCC
Z1c3RKj5E1cz2m6E0SEkJmXxfyZGyO6rQ6RZPWya/8dm1DYr6y3x1V7u40eeKskpcAtLLhdzkzQd
wBilg1kkAioO0XL1efV2JEtmDgY7b3PjjYl0fPFTWiikU7bdDOQvo2kk1juzckINZ0PPQD2NB6yY
6zywsbbFi7oT2FnEDFp0bJXITsjoh430artsEJdOQhd1Mq4mi4LJCZAWbzxVN529CaJlzhL3wLUw
ex2tHHoZKFiXHy4+kwuWFJgUKIJ2GTn3NUm2ldd0EHz+r7wOl5O3B1PuAQaf1v8cvwebhOKLtCwa
PLiir+uw8+82zVa2qwSVPtJS4cN3hfrREPfymb6R58wdFr92VI5Uxjz+l1yyPThMzhciqNIAce0y
xB6JbHsBtzUVTWHnhUn95xrfSSrJfo0ntXJFrymPpFF0vm3GzDWiKWpoqcMfCH4w1t6VALs2NYfx
HiUfl3q8L91yYMyTi/gkIKHmDTAdzPTos47CU913LbWtuAX5u7JpSO3FTsrbEayOZr1eXXnoZNpG
3c7fzhjWCK/3GhfK7tN6pV3+vW9ZGr+uwMmBKAjl8Ct0ZeoBr9z6hLzyY4oQVOy02n3E0sq3ITWj
8MFeo6UFA3e5y85D5knN+FD5VyxGCJxf5SueBB0mpLsj2dOEGK/1lgHH6M+dfj89VdASwm41naU4
PyXu/+P3DQjaIuwwffbLWCA6ukOLPGzWnuzpcaJaVp8Bl4JjCE4cpjJ7MX4dMUzBweQWH8AaL/kf
jPvZaxY6IIG9bPOVTgbPujrkiUP5VevmszqaEB5v7KZ2pZleEzgtETy0ffPHtz4EsXSPlYA6XP5p
tTbco0MxiNfiHZuWjncSK4KrwWLIZGwGIUzD3sFHbGMYWe1yxYBsiuWCmyDq6OoF6dPYNgL04QAO
MZJX9IGOIeLZmaJMbzCaJALXrj5dMgd0V0me0aJizKmqXctR5I7oVu4pAJ/5J3dcBqpgvCbJeZgA
6Ncz+4SvI6nFIIZrCuXQfWjbT5g9waTunxeHpvseMeECIY9aqphns8HUC64l2PywH30qUI50Ydsm
BJssyl1IiimytcnJQ6FlmQoDctZLWkdBT9/hzLIVGDep0RgxjQ72QHMDu5u8dkV4Px4QuM1pnTC+
cW5gtxbEWPPQ+8Hlz3zUBPk1ObxeDzGZr/FO9oMqLxbcMPvx3zzihHJTbWBXgLWkh0/cBl2drZHd
2INxgPSXBXMdHEci8OTvlf31H6HPtnA8SoqnsvC+s4mq0PW+e3ZrUqcLS89vST5lMuC5HvUkFhUp
/hZi7oMUsjcpaW6wq56Bb3jTk5eucRSPDpqBdOI33x5AZBJV7RLV9rv50s+YYTRFSjhLRqrt/OVc
MS1W72uRbVUCxFNAaOvgWaskAHq2I4Mf/4JUv2Rd2F0oTZ4RRtZom3ANcGMH8twp6flhTn2gHWKM
KXSB0F98aZZqdOdE1S9wfJyTyQBN9Y1saiwaFaDM3tACcIg321PQm1yFLarIn/SZRCSvV0L4D02F
C0rC4KIcsUVuuN8EDCvMBdvrAoGJjnegh7nefc9qn5KJyiq359QXIQ980cE0ROHrtEMxcFIIZKA6
Ws+CLZ+ygI7cU1radk/7MZUFfbZ77RcJOxh/qJb6uEF4QC7iB2HjmRV8PS9tU1yoSqZUfw1aXc/Z
QYmoc7yowlyxQaMZ75rmO8RKlknjz5XD7UOf8ql7Lj/iG6DnXNAyS6ezWNYUqKtGjijSaC4fIylQ
h1qhrabMw5fbAdfak7eAPuxlmoTbVUFy/MzBco/afa91RE7Q2K9tKxsl2l3+rZMeyw9+SVSuYxBN
eBMco51v0XBahTi/hQuwusulZkarDSGEBDYEO5gv8hS7mxtmdPLadDnhW5UiwhEOWiWJQ2yv7xq2
T0DaQbTS/3QE1ciMVQoVfp5EolLbxpXXNYK5btXJmngg4JUJCX0VsB6psKQbhqOTq7Xjlk5BhpP0
+qM2WIq97GPbVUa8H6tNfjWr9RBry+4zLSY888CKcDcLTENQ1EjkifCtPZ+ZRRQqL6XR76aUWa34
GnkCERgk3wfhDGrAAW2kHxPg93t9BJgS4KaK4wjWW2wTA8EOayQKWArP/awzgNcMaIS21n8yieCx
YsAojryxlN7yvJPCwFGuQ4xA+8BEiFeNPrApSfdZRNDpM4rm0/JUdMRLJO1RWrxLOEhuaaWduWDD
SgamFwLg0bMVx0e7QmlHDfNb+K+6nYpEpMME+gVctfYgtbLZBjuQg/Qpuv3JGFjzfYl6QSVNQQP/
9N/DFi0H27UDVLiwS0/5jIQlbQUEHOPevAtB6etHT0z1LxsAoSzTIcG695jnTVhaT2X0XwP1eDF1
EtG0UGd7r65gkeMUZVqaDqHf2vnnktqivzAtjoNqAP4H1yxhlLd6e04sVNATxGZ/8NdeU+Gukr90
JW0qA5T9JBgpdz3PJi8jswgskExmty1V8v73RlwwiRI6d+K8qN4YlZyUnRICRZwrFvYFZNoFPNoB
ulqiDNMBVCodSit73hqNxRUhy4rGDocvhKUmVX5MkJRBvCNMckKhxXg1GdPz1D7TkCroTCmR9SSc
ve3XKcaZd8Z320S0hZ0xZQcNdMKwcdyND99aXOspU60ZIKf6Lm5laWvzzb70vehtMJ9trq02tjkT
s3HBKt2upCNkIpFzVoawWHAJjWtAilH5Zv3DHqC9aOPg6kJRv84waOLy8fRBcoR3Xw0mg9ahN9WT
IoB+3mHnDqEw2lt9T1Xy5FkMf54IFHFoEyEj7kjBcAZOrOBq62+hb9Ou3nCTfFs5xiCSqAdOBi1b
cu2A67CXjIuCGnouWvldGKR9UEOJ7wTHe9S7Pf9qrz0t1qzqp8pXMkZAbUdBZxC4e7jIUEfsJ3nM
NKQl5yF7sPjD7StGp36c2omdxTAOxnlONBIGIWQ6uODo9YJLkT/Y1csEMMrRku8Vm0zrH97GHOGK
4oVWRuEtFXQoNpjkBnh19wXSvHkr0tFuAYqjZwY9Pi91UBGb56H37WMtNSQ1OCgD1IW/7Pay521i
05mNCEaXBYC/4mAs9o+Hkx0CwlbpZ556ENQvWTzwQYSH9jERnIN9JJsRDwszcc10riVuzowcvB8f
fVntbIT51JoNqMtuYh4mkanIGaOvYybMbs2o/4l/Pri8LAy2Ztlb01u+1YGeZkLVH89k8DHTpeK7
7lzLCNEswIT6XJFidzNKRwU0+F4x/PF2IOsJ6rqVilC/V5VAmXmevpGsG+qRL2e7AErI9/d8LNMf
MUpqPH+pivw25yjam8XnuRUgmY/MTvq2VOy6TvT62KjN2J2kSYCOAVuXcrS1pLmOUC/YXWVD/5SV
PddbGJcoX/KVAHlI6BmQpJwB7TmOxPMC8XqcY/B4DyhPw4AAs4CPK5fzl/JP4EbCbJrAlxK1XvqW
1X7Bh9Qw/5ecBOZvWXnyvcng4epf3SaDaAWL9w4MBRZMFYLwvgf14fjhbTSptF81aJdI7nHVclTK
/2tzpCbqpE8Z2eqZY8gtpE39BSCV//GX688kkMIFU9U1uTbAOd+Xxmpk+33dmBYYE1N0CJb4DqRa
MOV1x8SDx1JpofcUc3Cn6Lo6zMayAeIYIO3ZasTX8cbTJtPlE58ElSVW5DLKDy1PMuap+102BMdM
nMC7W8C+A0NDUxsP8vx6pi3pVII6JXQ8kcLratIfzVvXp+USILqxvBVU6ZWGFV+j2zfmSufWNGYe
zCa4T8brMCEfK706zvQKubUWNeKhO5RwPV+5ULXZBNH/Q5Vod9e5BtXFEk7htp3aZ7s5hEGgIMx3
xiFPtP5/VaIr3RVvKd/RIuthQBZNx9q9KOMc6+qf8/C4UUYrxoXHy3lS0Yz2k0sG/n8DiWV5y/KT
+6hyeCivQIPdoWmR2ffHVc5xPtgYgRS0jBjhDUjw9QZo3GGwnUZNu8KGw0Dz9q6ac3glprSzqR7m
54wKnZjA3NdwyFPesYe+HVHkBUxcFp6ACqfeRuxSINPEMBuc938F23ZdX8/q+FUMkmfaoer8/FCF
XnE55Rt6nuMYrnNi8zoZ1+UuwdRJuMOQHai8eHQ1zmkH2VZSgRTvxeQtyeVnIc6QQdK/zYXEyybJ
DwSVYXwFE5oqOZg6KT35/JoxhUiZvwKDCEJRtH9FsamojS/Pn1uzBOO6HgKQib2Bi/a1/pz48pQR
qq1jbKHchb8Mm2krNZbhTA+lVML8qcXh67BsEdbUaUe60VZ6rNF8Nnvdj4CFAUKYPe93vSM2f6a/
OzpuEldaF+5xMImt/HyPLDU2Wa78E6yofMI7sQ46ggeMv026MFTh4cBWMypGrX+Gw9G+FOLWk+o2
py9/PbW3+xDB7Pnng91L62Ma63Y/P4iCc+EYQM4+DJ+uArUxomLS3BFl/kwL9V2kjC6e8PX3s0Z/
5DEB76TqRyqBBvgc/KpC89NrEpgN8UICtffnvFUhMEGgLUyNdJUGjVtOvw2+4L1mQaqdmpCMNWJQ
Reuy4m9vrroIiG1Bhv1kDM67BRpxjugKQ4+6weslxpeGOWWvtoHjmkacQofyj4oQszUaFsvel9SP
tIdcFbmfSMBa5euB3z6ak35Mu5IhYD6807Bql3gjW5C1myfPW/Fsc6RoP3SwZqCnKo3XRnlYrlfy
8gKVr/DKYPD0zdxytRkV1i5QytSlR9T6j3Y/VxZPFITYQgI91EkiHl6paH/193GioRlpTKyZNUNz
APsWaAUsMqLmkovoHpFTbjh+fabkLm3hMiXU9KVuqa2ncLci99TrBAlv7GgOBNJmhYCrlBYsPUka
+/wA+/jS9PBfw30a88nEHAFv2E3+0o9EKhLRP/QcYngfTCPiqitNm5t5kIvkeWbSs6kMz98Xrqkr
69b/JPfEa5BwxiaENeWyOZ2rYs/HneGKj/ERCSaJNVMkEXGpRPAlYRzyHdySpl9xBoRw/a9t1EGY
ay5d43RKrXs7T04Lbw8u0Sw96wLgIdu4pdCa3APMQdS0gqYb5UVhaxlyGa59w8rwP6nLw2/0yLLb
N1lNsQm+YK+qZt57EHHSE/KPO7whPzHBT1ydJFOhBv44Huv0To1sS6kkPI4qnjsAUUqZvD5w7Tc2
OtXG8p6I2QmTLB1fEQ2g348t3bdZQkNFuWch/gdKPqWF8ORO+xBR7BqHRIxexvd90N27VTzQ3uGL
DKRWo/wAXVcAZYVUNpqfIaSShjNWuVpHpsl07Vs6/K2Fl1sO9uET8wtvEN9l61fQJyphPTJ1IoZL
g6ZsHEgQMadpdiZwJzkIeHe/ksuDJX48x17bpjsM1JcHWi3krl7c6Xx/ou5XbD+/SzNsqEjVAE+P
7pEUBHeZhzjdGmscD+fdkP1eRPwmmTxUdca8X+7UHzVtZEdvI4UfiJx3+54aAcU4uMgsPbCQD4DE
m3gQpwvpOMDVW3PQHeTj6g/sBIWAc+SrDYYTrnNkcr3J2EdDYUqurjkLtbLF8+Dk937ziv1WzhwF
rzVw/Sh9fl6SOnFqbDWgzV1DsPBIbEp5wYNagIH63CGg5ssl91aMRQTPJd4LRa7j4x6IjGF7Klbg
MUMBWsNkmjZeGu9l0LCA
`pragma protect end_protected
