/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAAtVI5aZCFGLkw0koOIuztzkqcaTRkNinDkbTFdxxvHc82X7sqCC8S/f
eGLYewQMgMq1XcqtZ5QKV1OntT87kZXdTHmDOalhi5+ZeDETbafYVpuiVoaNJC39jIrjgX/vzveT
/1aHfXtFu6ZBEwO0oxeHkFQEclufqWkP67tm0fuq7wquPwgjNBflwtzuBPvuKnTZmf/wHAI4cZ+J
xU6Q2/Pe3iLsuEiI935YMX3oGp3DNLC4lYnX7tOpDhFEARL3kKwQ2kP6pkNsm9AowVfBcONvUhDl
31EgeKud2Co2/UDx4uCVljHpTmrozMMH7vt0xC+MaE4/gaukOEwavTAttKn7GA+MCZ/JsztD5d3u
AW25ppV5XMJAT+bnxT3mzFe2N/ORBA2qQb+YmN3KKSmvD620pH+tEsg4igOVMdUwdjuzqwRaQgPe
Gb7CR66bMEm4NW5KM9WF7QGt2MkYQQq8qcob0VRAU2XDnRoNOUMWjkjbiA40JHeLI/B6F1Ecayip
7uN8muesdO0f8YNHvwVELsi9V5fnKbBgQ8CXxQyGQpUHix6JDgTnCWgpRcVSG3WQAEpgYn8demMc
rVzM2VkbwdfsgnklflW4F5Ak/6+bc54BZOR0Z0+xY+Q0GZMKMA/QUBx1lIzNMVsctNpm+A/id6LG
VHrNzMhjmDYksAX5bK7cQSB4tB3LDG0GS0d+kuXvSrRKOuOdQDlaZYuGuieO9mgkNgUabpLoimrV
SJ6T67JM+w/2GKAlLjVIGA+JqT03Mh/mMNup3O1OsZrLFhLg6aOFTe8mgKuihalFa5CtvfPRYdsJ
58dafNdSohCs+lVad4Twp98W056izB42t6swEWTIaQAJ7amGoeA45lqTm0/sPzfYBrLI3O6fQYpf
iaoCnTDY71kB8jPnPsD3FWcyIxZWnKy9KmSmyUyYVklOnRq4TFcYtEMQA0UbvDMNvgLi5qhQo1+v
Cv0zSjBplgaVhMJTHeMFcdfiLtX7UEBWDg9GOMIEIHzgRHF3jXPudCyMfqS84BBEazzJAvD7hQP5
x6E/saHBBtTB2ZGWo3YjBmkHmS7MqaGLgEYD/1FnzAN1NEdaZaifUnr2JqlGjCwCezUjjJbINMNf
KzEczte7hftJv+3q7nUGWRqNkSU1ftdxFzSsYvYcuC7uY4xrntIvy1nqxt2f0uMsCXMH2CiGv6EE
o+2xnFi9evdbzaXjeHGoXIiiDYoJAjQKaCFvCLBwS2yy79HZ9Xlo3111Q4bA4AStU+wvJ8USxRgp
b8qX7HfBfvxbuPs4i46Xzj4mr2zERc8=
`pragma protect end_protected

// 
