/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5744)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHIcQmcLVzx+N5v4ymSgOgCQGG0v5++ZTJzvrbGtX47FhVKMu2DxBguJPY
M/zA5DottnuQBreui+6jXyJC/Y16bFcS299HRr4n/kqclnFyJoxGUGhyAJKpecjXqCrjJyZ1lZkM
M0dP5HMW2MSSuL9PFq0CBL/qNWlK99UR7MrBIx9n4877zkUIMb6kyx7MZfcUxxmq/CvgjGw5g3sU
6fWBVZrRViMS/wygpecTAIKa75l4fQRd6mbb1+jtgfKTL2qokm4vetjIsEq/G+Vjn35Yh2cEiX7I
oOSESWIpS8kAJmaeZXSobok7ZQ6H0QnEs5Ura/EPF4pk+z9ciZdNHR94I/c3pS+QFRtyKy11JB7s
vpiKZsPv8rGeb5D8RPgDUR/vAVgLig13ivLA/0fasM3/BA1K/QHJmt9wt9JA4E5HhWf/e17Rm5JF
+RSBZHCqgnkcrrGhDZbIbhhakgjPrxX18ie0tWRzOjP9E/QtipTJ2B2Oz+B6KF2cUEfWczZti7ph
6pe8g3tSytsg3eRCmSMuWqllGwSPuit0A0yWiDcXX1/t6it3AkKhX/dRnYCQN3LWUv/A7grScEzx
9R/LliBnXl00Shn5zcC2je2ph76kaO1mKvJbWLqwXk4hi7/WtBzHfkVD1m2wy4AWPePy15MhkhPg
H1qRR5CoVknO5d9uUELXFnmyIl2PjVFD+AgROamC904h9xBCSC2Z0r3rDL+EahKU/R0yWoySceFG
hQGy+fxjiKu4yZNVlWfLjtEuj9EcLu6ak3dniHvIooPF+vs4Yiqxrx/oRWoDwhJo2F5iYbi1XK/D
jICWoZnGIrUOzN46mpD54LxTjmINaeBX5dCZ6X8LPZIiq4LLyNcXFErtJsYznvIkBq+3ub1uZqKf
IeQunC3YieEKsQjHK4KZTa09RZBbx2pj6TejtD37wY77IBpW28zr5EIjA0Eszwm/WrhcCLewKYwI
Ib8ir/V7fyAK19K2UTI87c3kv0ECx1Kc3SCNDwc0XK8/b+J4hzdVwqzlwsr/rKcsweBiZeRLp8fG
Oad5jUXqw/tB480IGpcUPERGwvbuljtchKkQXAfyRPC8oP5pHOg0Yd3fnQkaYLzh71v2G4GZ4YYe
YYY0RJVLFLUTBqqTYYXyV3K6WmL3t7OYePl2JvctiucZ8pCddQ8RyJuS+QGkfrr70Eq5TyNAFhxK
DhCtbbm+xJKNX0MemlOEKQY9Ejvf+/o5dEVsbkYlm4TzSbFXd61h/YsUV+6LwYIbiMUKZmVYgNJN
EbCQkrRh/JQ6pKSZ5F0nff2W62cks+/B30QXrL5gdiAsi1S7Fku5Qv5/+3wWI+onjk+CKTF3zuET
yx6SHmalf62WhcmClX8eXGqNNnURUjSe59i8zN8DzuCVeuENS2oQR1A/nNFow4YxaHHKKWH3KTlF
CNf7mme9ntOU1xEpEJWWPqCcy3fgTX+A2cPcI63ONHkU3opKrZr1ofXF7+Szt6xSvOuTNujR6WyB
CGkkjGoz2d6uc32/oKNJwxMeuXzizxQdSmqMslr5qpVhtuuVJIDIPVKo5+Ddz5yPv4QdLDBLjXkL
GnKC0DY/ifdpIOWjQGuXMe3wj5POxaNtWvg2ngx6UAre9gJTbji6/miAN2uqDhNXRLmzD4Z502P/
HrOPk8q2serWRs3NWG/2RBx/1mYqeFX97BJMjOlrwpprVUIAOVzwign37NzTEXGotOH+H1RGGOU0
+r/gvjwL/CBJqc7umYDuBtstt4aPZatx2wGStvzqfokDMISkXL1vuBCN7FsWWVQ8laCE0qHjMPhq
oYlkpX3QKXaxvHK3CjKNZscnGq+0xOMMrN3oOa/JEDUlDBp7iNOt1bwHMmEzNM9D5DzNH6eqOCnC
IadzsomKaRLTJRK9VrN7Ycuuias1y7NJF/l58oFVfTEefnavXPfpC1SwrkC8m61/BpHiNWEiC84l
EvzQXqh381gAP6FB/cy+bJ8cNuk5n0SVjwxchzIdUQMGsyZf4P87dxZFY8LnApDqe575nhqlIIe0
Xd+M3OTUaS8NTRaHW8APhIby4ChMr/+tPfwI1FxzxdkGsdoiMdIKxYhfSAF6Xk0srpM31mJg2Ede
LeKpT6f4mew4/xX2PYdSpP7SQ9T09Q4E/RCQ/AWT6OUgliTEhrP6W4ov0NEcxcPKB+4GSxL3d53w
vvF/kov/nBL5tOagOMvHS9JMZZY42lANFcbcCZUIxu3KQbn1SeZurx4lTxNfdI2z8p7yjP2ma87x
xYbWgRU+BGSzDMh9UCeOTkrfID7vH3hGI9bmhwAmn6nrqxDVnb7Mw+bUbjN5iUNVWyiWnDxBRQZ4
pXJpFM/6HzSXa+DeK0M3IFjVS/RaCcz/aPJXUbw8ti7SHklLxQ5lWbDs67dhLA0vvSzKemRIb7iy
FdjnF9KVZxGPXbmFwOmz6KYJWjzYq8xREs57bLKwEgTnbS7kNvdjjet2Y7KtjQipMkyOlnZwgwqc
BwVuBzAoYNXb5JoW2CCGKUCr/02s5rtBfZTTRMvDmT3cZARSWjCfkfbfzVtwHA2guIlSMP+i9Szw
IGNrvKU2k6NxVYk4hpv7rFaGFiOUYpSie6LNwZFGDcb4OBCk25S8jw7HHf3SzTnraAULYUUTVXH+
P3iiosHdkosmLBuX2cXQlS0D44/Yyv7CHukFaHHS79yRO/GVZwRI+tsIZIfKlgpVCIUYGTT3XPS/
oKxnu8655qaWUeV3bDxfJ8sGGf8gLro0kbqb7hjqffOWCBjctMSD6KzHtV9r1d44hO9aeD8FIDm/
w9obhIXBdGdK/Lf9p2qPVWdUUzSC9kCt9Vsp+ZYLnaZNm3NNMDRktWcTczk1VJNZqiHA6kBTF2/w
1xmjHGeQTyyaADcOAcMAVTY4TPc4Cwszybes3kUWL7JZDUicdKUwHdlbTqbm2bTcoNZ2YHd3JKFM
i8hx/tWuWjd1znNy8CVCR3Y0qA1Fyjug8R37Q/Sra1XSAK8KfzY8RrqKaS6IToPNnTMfAkiTBcPB
LOtJfeT/MIlXVJAcuatmC5xT0HysDUf61VZirO4DRGTSZDUyM3eACwKT/PZjbbvrzjSsUrWxj1v0
RJU1ocL/GTJ57VwR7y3Ba/jMnNSeqMzyh4Em1rEc/nJJYQxx6aFpvB9uF17Yhtv4piI4ohPhTS8+
Tr9eeAmwIKLUEWH/WJhHkOkSebjpTsX2/kgn5BiD5H4chRF85nHL/oFSyO1BIeUxVj5JSQi/XR4a
301BBYRRCLEss94g84NB6v4swZLcsV9KhQq00GDBpj7z45mba8zxQVqVYz8tJb1GaRCSVmrZ9gLF
VPIZoQpv2M8CY7ElYufXz1NW6JLH4n/sgbYaPjmN9Fm9qY7Fr50htLYawAXgeanlTp4bzsx3PZ5O
jVTHROvxTF+IkbiSr1X+X4h5CyJ7wfRqeyNtHEkjb/L4nM9c7GdkWB3j4bC3yuw89Rb2jvowVwLX
lYbZ6uZuJbbvDnUCPwR9Dwi0XiPIp828Lrtj9Zzr3edTUuT4nor52qtXfLI0jM9Mn1MQr59XEJbY
NFXhUhuyY2pHDRxziH6sPjRCSdpLxIuuKzynKKrhi4LW9TTYgd2CTZJ0G9a5mahTsOSj4q1Dk1yh
u4L5ONjBYbwpjgcWjQ0zes9IjcwuBDSz2lDfxA+DNhUtG2Bq0cdWVGFHOndvHtpwg+B7SMcxtHgS
OYavVoZzNuprGojGzKWPml+4J8lh1sYqyFbNqY/NwJc6L+3KVWW2K076sPLGAsWE4BHFazAten6i
Yv8cxDXLbGc8sjAuOH4pvqtUeVe14tUFAIc6kWNP2RGSNVJSDisJlWZBvtaMThVmcRZdNnD/zRuu
R5XBPcWcfI61tTNUFFEry/dWli8d18IoNBTznIyt+oq1xOu9x+p+NmjDxL6SmbDKwADp8w/pPXOr
gNXtzgB23uMYPYREnVxMYZ7l7fjqHUdGQUI4ibxbOlVdqi6fACAe0OAER4fITzTyJw2tUbngRZMC
hOhJzFG5DoPq1qL1j2Te1/EKuvUIfIEoAUdZ6V8H3c+TS1qpFanJoJpbpG5578vEuAzcOlC7vOBj
8Zut8XvIo/z9wPVrCmKxCE2YCWRR8S5/TaYNJB5KH3vcEbH8b8cGk0sKLc0OvdkGX5subZos4zal
NxbftNXFqD0xQC7KmRTuk69cFgiRngrKndqrBg8ubv1B0vyjbefuJmNW5iyT7fZhDkA3d98itDz+
xfcGJjLuTP84njJpgzoiwWN3X6ufYaGQfNi8yCiQ1pYb3Ax8ElM0uRfxbAJ55IKgFbwWlv/kVXgh
6A32sw+sBpkm+xj1iOquX5BN6NY2jDe/jW7xLBpdi2nkS9bzIESTCL7wJiaSfgWIQz/2TV+Y5BrA
OaLgSHbCJ3bRSBWnq4rQhXjwinQJkCkDLPwwSFOoFx6UaDv7mC2NymitvfCOWNHGXS9LlyTzcK4E
mZAn4gOrH2c6K72+/ymGlO03sDdoGyh4WF/r+shNPe28Za4r/tKQ4VWq7FAiZQo40aLvdsBUvNIE
HEgZG8sIDnyiewrkZximV0UMTBtDCXtKkiQL07FHUXkLlR7p1bROYwJjp4iwdCfLNlow9izPcYpN
Hn2nGLVazfehfTJ1hJA8q3OId9lxKdSf/50S3f+O3lGyrhDPOwORQ65FzHF0NGHJPeXyoi/H6IAR
Ct/vFB4l7i8rQPfV8Y3n0PdXJciA+E/HawVo8qNZPhEhpyfpx4ajejUS/yRTfdNyHR9HrFsP5pkS
eP811LXKiErVhSuUdwPqt75CTttBLmV2UsDwqZY5nX6QgbNovzgzLP7uPr0w1CdwAF7v+4/d6Iu5
oBbyO+W65fDvxrO63leKpWlKGXJeLjuMJtvhEmZFZgMRbJkFoTDvEdCm5ZXaQOnewGfi2jKQXOPh
S897OZIfJr0iL+NIj9Xa6Rn09J8kWm/P+k7eeedmlLfi6/SA9uyrGceCK9nahThLsjIWyIQCqJlT
0y0W8tUbG8HeKS9KUyG8JqXXN6fGRFu+SD5Mx8JlbVlZHfPAyCTqbw2ru+ACkxjJJzLVmXJ+k1Wn
JTznnu8SqrrT54rXpIfB7m8ZSlWDIVh7BNPPgsFURmSke+V6GuxwJCWauX3STF9i9v3W4u/55xPr
toQ4qd14vDr9SV3Vs6jfekNPnJWECH+p/zYt9iSAolTP746QfJ7JxurG+T63qbmdexJcvDNGTnml
FcoOzsBwCV5A84d+wABVXlIPQRr5wLpolT+D4St/v63X5E5u03mtpSVtcfdkKxjBSZJZvvcAqRWq
w/e2JGlPPSDXr/RteDS3sLwCyIOYmb0jL63+zpCRZgtU1Nz/Qnj/cYkOUU42NJ7gxe186MuUhxOG
yz+P53xXhbqe2Tr0KQHD/vQ8btzItjMa5+1nvhhiv4CGj4qAIyCnnop+gA8Aw4Ob8nLnEb6Zt380
S/NXCwrtDIGHx8nL8ogp3E0mOy/QpHsuhXTiTWYPllcBfWYN4c5QLf5gsXbZ1HeYeGatwJKlUlE5
Muo6asEbJCV9a/oMRio4B1Aqhu7JiQTF/ybIldstMtzpi9XAXILYgXOxaqGndOHb6KVsp6VjI2bF
NHQSVJgv3PzqrAVWGNsu2D91YWnDYoWEcJNbfzS55u3HCzwsXoIVagUZwNnenwTFG0yRGTNN9cbS
jDtH2bJV6/yRKF7PwvtdPHvWzGigaJD/BrG5Prv+lLYvxsFpi92MowbJUNOGosj6KsIlskXNbCVO
+WaIYsqfRrc5ongqF+kcaWQymYOJetGMKabJJLu9b4jqRPKlt/vv5295df8xt904pFNXvPKieNes
aCKrRXcuUfIFoD5nELHgaVwxyjBUBfY2h5Xf6A0Z/eWx7t2qJnFg0RCRnjdR8g4IPtxaXu48G6s6
yueueDktMUQmkLKN4dwYNz42MDbJd3G9J9KbRquE5yB8TeStEH7gmxAoutyoO3+0HAgO2+SQ01vo
XHG8YTKmn6LgA7C5TmUKagK2FZn2yOAjqA7uN/GlW7RoWsE9nUXHu6616GrSGmW5u+HINpW5D4C0
EnTrmoI8u+klH11USeANI2kykYQ0fzO7aElshf1aBUfcs4r1xvXJZZxgAHRo3eUVwC4vv/mhkTid
rskK5sIHKOzk0lCHZN0YiGS6qudrhYkq2pdYAKDS12bOsFxqyGUYnwzgJpp98JAScoBCpTIuHXV/
QXeE8Cp0CIe3wj2iaV41yuKSSYf1erIIERJA798GBRMNz072s7HzyMCuVLFzYkPJCNb0UWvAoOSA
jUEKDvYbYRiX1YRAsnaXfXpTsLxpuxok6Ln9AQfCKtY/XBEyzV7bzoRKIGDIzOTPoz3B9E2YMP+D
qe5fJ0FYuzXJ1qRvllUeFmWZrgdjxSnve14zfpOn/TBBrtN4Q74IzapnpsCMNsuhM6PS/o4CEw++
7CBSv2Jz97LpCX7p1tGNoa9EH2mVAJZywiohGKyJWoxpJ8ZzmR9fD3IFbfB9RalzmMMp1jvF8jct
+9vOIuS0/NnSrybJEqIN/KMsZOPpcvX/uLrgTkdAiFqk+q2eqDSxF2FaeKVD6Bhdz+So97E2ih6V
vzTuVIrix1s3eRb2hKz8nxEvS90A4LMjd6DKOQToNoLqDvZnliQ2IZ1Cb4FDk9/IsZgBHtebd+dz
1FlRWyv+EOEo6KaDEtXGwq0lllj0Z2rxZ/uPIdvPG8qTvM1lONTDWjUdY2n9PfTzmZiAfzhoPT6P
6qyDFkBVIy9WmEA1PBnrG3rtMsE/YX66lQ0dvk1IwWfNvti8jfrwwuejeURSEWBxxLgBqqBFBKbx
uxJnv67/ukmvv4sJ/Ia/LdP2EVsrXgiCpW+0msYcVjtj2R6srefY4WaeIOa9uG5beabVkPBOVZsj
hQ2ZUENsd2/BDqsxQUcbQ7uvxsKhxLDPNEKdCRa7PeE10C3rWhIaCsDn0VUWNpUghQKPdgS6BqYj
m9w3GP31WUgz5pkDjdUQpDgGjRZur59xDnPjj56DKoqBmW9EutT8DROxyWjZl9hKbKxgtgkh6R7c
GOTwV0ao/wLClSKDS8OIjfFt2dA+k6uMfv70KBW12yKhnIYnZyQ9cL9dTLhKrRaL3m9efqZxC9sI
gTGnLdaOrSeQMlooEMo161T5ZpKQIr4AxS5Mtg35A8Kfmq/qUUxzpwgbHgm2VwIynkMW7CUpFqi+
eFfkg5+1x0Mz16oUtnxI2I/YB0/aNACW314AS0eLY+V9bl+XAV/7cffMHscFmm1gaFXEwOoHirbg
4AAOi5bZP+eOTFomGaK5sdVAV3ERACuWeGh8MActTo/U6A+AHkW5OgbYi8lIGSitPhYiEzLtzSn+
1yaPOWmp3Z2jCNOpSUW6FT/nexgJ/wwjZwCGv/zvSoZesKY/yTZ/GUhYIXw0XXodaw6u0ZLDvBfL
LLqow0BRPjvyj4d0hyMm7Z4Aw1NjGvnsd99FbJkylSguR5yHDAXwKXnqBtsVLF6mk1P5sMThxKGq
hQ7dBlTsJnxNU8e3FRkdzz3EpcXJpLO5MXdTatz8B8miW1IEyewRx64FgUs7zlM0CWdbDMTrSPbS
o6+bDx1GoEpc/ecbIY3/WiyVm03PtTR4rE6/Cyv2otbEICnM2t1ypaVDjgo=
`pragma protect end_protected

// 
