/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52400)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHIdJJrGVFHax7CPaoJSyMptORLTqt/RjnlaD1cXog3149w5oNYYsj/TO9
smLU/dRH1FTe5mUG8MXpUDTu/jRRY2xcUrJPMBwjyyBvSuc4Sp+oniJz+PX8IhbdcqjwBCtwfS2q
kxkDcPy2ThjVEdl4JI1GIBLAj+yPkDDgCI8Ml/6a0zr7f0TRb+QnPv3vF0akOSHiKrZ9rCOiNwEU
ql9iduSb/5qCY+x3PLTVDIgZwCWXjbJ9iu7v+OYSLn6a7XnyRTa5lQN61knxmp8Q4zlfDqPxnLQl
dh3sWtlNd+K6GWFvQX69cgNs0MMQhdB9mBEPWqHW9v/x8XenLYDH5K8PPFN3BEy/sRmWmrA2twig
P7GWzLvw9T2RycI8bRyjPX8rmrksIP0nbMSaEk2qYypUIAakZrNq6y19BDrWBTPoHJoEPFU9F+Qv
DG9K3iqhgzgxP4laPQ5QoQv/uAPHqiRUpUigLKdfCYVmxL5lISU75lOlM8Rgs9UXGfJunB1b9cY8
3LU+UoRHLcjyW82zvqUMZuCBzZZ/IHAXX2LdZDLf98WfK+au8+e8iEZ1RNV9Gi5X90K6ckmrMS+E
3enD2iQqWl5JYxjlOKBAz7a7Mkq/qUPMRWEiIWrxdjyvrZvsb/SwvwR1xSIdVJg+i9jhAQk3j4kG
CNR07wKa3BPapNlPY4qYhzhZkder+Gu4BXpEQMW4IBbkQ60K/49gMwt/LRvuhd+NDVXcgsrbUhLE
N9VOB14Kdc8nOv9zhmBxPD1G/HdFV0oTIyXKrXwu9m3WgerzWxFQz3D5vkrWc2jQD01BUg+pbnyP
uQW6EkPe3yM5oOBTiFEBU23mSq7MKKL7tsLpjtRprRU2Z5JMd5Q5UZHzHIcfj8EQQv9wfQ3n6tEE
RzXSLz4nW66bErCbqPDBPSzGI7xfgcVP0tl7qrR0d6X/cxbcqmB4VEbsPbXghsz1NcuvukoMdz6/
Hml2O7fAgbXwtzZtPVGNg1YcL6vkKe4FrDtZz1CECpz+2S0XVP2ZkfcS0h+oi2Uz1rTJdDBqkSg2
9dgs5R3cnV9+mSmtpAyWKBwEc6gvCqC/3aPqQgHBKxiRf4R20U60UazmIgKfmxjykBF2aHbg2SAu
k1nNY3pGjU2J7oM3u/wWKTExac0Gjm8/9Prb/d0h41vhNsRP691TzU+GGA8hR4UZ3oPRXy1bo4vY
S1vkphPuxW4P5wZH2K+v7qjHpPjpUM1yfYcRYPL17LG9D1j54xvK8dcoTVhGsZDOBr+ENghZW+La
KSxPQWkg2/AlLv9gwNLsRAGqexzOxPc44c/bWYw3dzPs55QWve3QEAWOBaRkEfz/KgNHcDxsByrz
PRIAkfjuaQm/+QO5Qs091CM+BZ94dtFUzd+X1gTZhgdA9Bf5g5G5NHAoQvzq49XSNBsyn+fATN0U
xicCrBxgTTQSMi4vuJGJmdo4GFOBdg3SpK8SSYypS1TuKha0UDoDUdeK8glRMiDtP54TChYTCmet
6RtO4ATvYe6YSCNAq9d7McW1hgdRHyJ656x+6aOWdvXuyIYFPmideKUvpnCnf0hnU2pPf9QYAzUH
5MuN2g/s0SCxp8tswNz7YdhfQII/zxfFb2ltczmZblZ9rOw2RXRZTZbANVFQ4mRqAWpE3lTSgeTi
OTEOJPImtsxmbwXuC3V4pq3x8NLuUbvsWjnUORsJzVSEThZ9+5bo+vjNavco9WlSGSKzm6qsVXUD
jV0BFWIX79RxtkBzC++unTs7m6Y/1ZdBKy2oDlHxJDQCm0uMLDWGnhY78AEWkO5bBJ4qonlMSl0j
+JTfjBj/jaPgVv4fSAEefLxFVE60SXz60Fm7HV1J3+3LoWh5uXgZ+rrMNiX1C22bR4eEBuA5h31e
FWolvnMlVoO4DeJ7VimC30Jz3GIAB4SoWX1iJj1HwpYqozz/MN81R2zgHNXxXIUmcnHonvAfyu1q
33VGSolBhemr3ms0Z5rdpnWbFaQ48vWrVo8/cCINrtYQbvWsUnlPdUBPUVnqcpERWsn3W210kQNp
O6lglILCzwni2r++mTqQIXoupQ3Ufyh4n5Gd16HFj107YW/wh8jmFsqMPZCo+VL6M9/ySYi3HsFI
AVpugI1U9VEt6j5wm+lDbHxjSKlnuiSuFYhbuc/rcCH6XWlq3Qi/UAxRd4KUnqtaLATv+akWe82v
0ywZ/msKD6/kaFS6wHYKjyN7AAr4aM+/84gWyq9pg/Y2q3clVSFkJaSRpc/OsH1KrCFgtTAWMqNG
/J3FMcjM/osoi7IzQE5RRL6YEQ7Uqd3eYujvBetADHCNjGBKNmgpE56FqFhLEVwEJbAdiwQqg8qq
MD1lucmMG6+1Ii7lyrTjv3EkRO09yvIhCa4mQJKcApRmlSbkjRWClpjunvBaYbPaZqhbBXTMqijb
rT+PhEaVh5AEwMziDR7CP2djgNgXEgjSc8HmBQVExYGRAvl2sl4GXJGtmKdUEal1PadUE+nhcBgg
DIro920wq8L0et3fdHs3cjCiFJR0XyofYsyUnmbdq11Yy40jZjIuW4CnbStc69CHP6qbAeHRwyzQ
lKw7wHen8cU1TGS9kRGLF3caioxCmjw0m4EyHS3rGt0wGXiu8oE88oGcg4srGpALuvgeQVRFkg2k
pgOmbMLs8Jo3Xh0k06IPoIb27ZjQ8ldAF9mnMpmrBVNnOKdE2Z3+c2Q81J9G7dek2+6AdzN8Itm4
jMKPVXscR4ilvs9jpAR3QUH7xHnNDdNLuCXj3Sjln6X2DZKEobeCqcYaXlTL9MtdQnCYFaE/7jor
S0nKYAZktxih3bJCIbeMsYsbEd1c47RVkbCvvfZ7rL7lrWkXHxWnilHy8brmEVssXn+ibojIrU0A
BS7wpY+Vrkvpl1vDjfa2SYdtzwqSU6tEXlEslZKDzseMMV45dqVFbwTT6hPOKSOIRg1F3oApo4UQ
Ip90Y4KsBx/hP2AFy/1BcSvUJq1sDuVIkghuaXba7y763tWJIrm6Zevrnl5B8TsHVrxFUWW1VJHP
Wo9rXUDQBDAk+ybfDnD1D+ValcdMjxDvwvc/wZtl8KH/zRq/cRsS2k433hp77amcFattohLLUwvj
hzQCtz4jF1FFYeOw0SZE1eJkj+DLkc2LS3LSpUUG26anWsswBj99Ya8VpHS1di5bM5P6ApNRk+C5
lqSM2vjy4Ay3z8W29AEaYfebiFsXoHlSlt2HAewvNhDpE8Myz15lMHEa9czwIyi2wPkjqiXz1aVu
CPzwWRp9FhMieytBN+k2Hji64X6UDpPxVhDRB6VPEcD9k3Itfu3Dz5UfG1A2iD5C8S4ZGwliwaPv
FCNhIbWf0I0Lxmve07ELJ/4/8A4Jx8Gw7zVYSxjf8NI4KAo7qUYzoJusQI0cgNjhJDQWRCwxGWFJ
NHzeR7G9E4h70GD67WERMF/7e6CKwsNra/RqWbvFhFP2rkUomioR5Bhk9KYlz0YtteDhohJh3AR3
Xx0rat0Yl1KNF/fI7Rlpva5BugI1ZJkpgAx7DjOHNkaUjUIHJf9yY/bg5hag7XbipEftwZHBjQ1/
jdV7lD1sR1u697Axsb6710mVDsKxNm2mjFaNOLdB2ro0eVqd+A3RIpW912zYOO2AyGTJBi3MjxLH
xF2mfAHmKqidfSFZmt+67BJZNANfEc73Yh8QRZb2A+apFvm8CosxkOnXXKo3wTc32ClOSnJUC1Bi
PEJ+rBVNpy3nbpTOT6yd5YPMZNYTzkCnWXQJAdz1ny54f006pIgGLnTsnCMg+9BB5R39Lb5wJo4e
0MTFww6cXrpGlnwOBjFG96Q1Lp5KWCzRXOjeoG5LLbB+1zlUgmesNcaLEhqQK9JODqdZ1nKWo2ee
bWirWdRQ7fc9um+nCyV5UW6socP2gpzSRmSAuJE1K2sEsJEPLqy+nsOM1F7yhic0jrXgt4XdBVH6
SZmpukkzZhqj24g4/ZUX0vDKxKykynGK+Mus5jw5vZPj+QaQVc3T6J7u7v7VhEkwpzpO+PpKjQ00
dhMAlxdP+EtM+MnjY+HUhJWZ+FMH9elli1pDCtxR2dvwf4ZP6wqvY/Tlj/WDCr2wDxUuitSOwRGi
6DDFrymoOEwEGZkbh4Rum0/JQsOP1IrxLYY/zcFIH48EdB4fgA4h1Y+G9kqGROmQ6/wDqAVqcAlh
ROFVaWKyjp2O9UDPQlp22AQhyJGmJO5BRD5+z4j+//yjYncusSW5R0KxbvjRfjz4QB9p3IbqKgFX
/8idO/hU1uAu5MvJpKvqI2vMR6bvBUDG6pvq5/UfjqXpBgG3CteUQtlA3uyMu9rjG2k4FNB2KeTR
Ldq7soFT8qe/bgN2OY9lWs5MOtXImU8j7nyhIfypjZ8MBbO8RV1haUE12bpZJHcfgUJZA61pgCDX
bFKrZtYf19LF+0d30P4T8gL3WN4a2R9FCYMCfFGXiF0TY7NoXy1SIUPD+6MzxQM/39FP8HOjgpZI
Zsn8f2gqsPlj8au1NIhwTk7TRTF5PFSmJ9/WBezMGQiWrx5LCI06lq+Czskd9KJVN2PfuKCNTBPE
oXpWeyhKVgSE2IvHnIyHnbRfq6rK3nowjC3nZUQ2jKEThihKRLKKS5Nh8UOuZ9Ri+CZucdgdMyh0
y3ejVIiMbUeaE5xHiDB1izwDcTZr7cCzhTGDkxCoENA9dZra2CXG6I3QKIDtLA/GS53qvJ/mJMoN
YieU2Kg9XORWuL+dlGIR3YsqGOiCxVBMhO6dal3RG6yy6y9wCuYOD4v0l8KW8K7w7RAYksruDb/c
gj5WJu2afhRiWbJsv8M5ACo46i66yS+RJ3+9tjG0Cd6DZ1jhH1Prkr+VNF4k12WanjuGi40y09AQ
zK0rzqg3ddxgW2TBQpy4dV5nptQZC1WQo1ZnIbP+kmNS5XuX3IvI1eEX42jkVK8TAJTH/3Lu+tml
3NQA675TZtArWverpafUW86c1NcXKcE0GozSXox8IXZXhpLZe3res4q15D22p1m59MxZ2xQhTa0H
fp7gbA5+DnM2I5jnhLwW+AqPX0mDvbBYfmK9aGgOk0LplZ84WYDessPYzKdCUSo8DasIVdYWMtkj
EN5S32FpPgdpJMccutPcBY2nY+xyRkRak9Vf6qr4FVn3ot92IvMsTHQirbAUfJek7CfUj4/EYmdL
e++7E0ikzBvzcjIeoOaJy+rwyt/VPjYZxb0y2YJ0GNDj/b/N419I3VwyjiPRUDR8avW41X5Nw+zj
qQZlSQPU3Fs9vdRuBmNf0WeHpLMiOnYTABHsVbB01DNStRyamUjmzm9sBC7vIekAw+YoSz4oQtza
J5zRRDGqKDNiBDwVnkxI1kl1v7j0FsiwmFdC8rPaCea2pgM7QNc9RcPFr/x5fD/DGemMFj6W5KN7
q7db4vQy7xV6mUzsGJbx3daMrq6ubYMBPB7afb5i/J5Lu9tIaD0RINKVhrhR9khnbGX8IqvdqEe/
xzENqWiHDYErfh8a7hqY7n6I0YtAp7BWCoGezcM3YgzbmLUCYQ+Apbt+3Nj/6qDgL03QTqlxNpc1
LpYv4rRIcdgOeun9inrtIxeLUye0YuCf6xP3B7yZMaq3x6lr4NhdD0HHJtoIKu4b0quGeUIWt1ZU
pi9Dy52hGuzaVI0W0dwtuNgRY4F0v0uqF4g626qPm3wS34ptcRiq4mYIK36tNTGHtg8i9HTjbDE6
+prIkmIfuD9hFISDWp/IWohjSFXqYq9NnyaFEIhYDnhJ2DHhSbmAW48HlkgXM6sys8UkAPECnmtV
mP2Q7zJqJ8VCuwIkDtfTtnE/7v8amOSHaMvj4G9HYw77NCjriBgErmagLgaNgesBHagdNUJFcIpy
LINa1XSlWVccwKLxFkq8ptPpYWztiBLViz0D655gLCd25DD3mDAQporm3ldFuEDlRAHdnvtrfSr8
ekbvLSvrM7dvnlpTiMDluDXECasJY55oqImALZmn1Yf9e5jSItnzFGavyJCv1DCrSET+sEeTntqf
YiJTa8VK849rk1+W+Gx7aP2XdxQKnzDjc4LKnVAwO+o/taltheq6LzYSfnMZpJlzIy+tIsh9mvUd
JgJ5n7Ahn9PgbjP/aKFXmLhdWiVI/EVDgj4DQAGNDEp2XkHXQEgQpOHHbXGEnst/ZR6Oge7WlbAo
SHgiu249YtqSXgjaPWnb6gJcnIsKkr0VWuBzlOpvlw9eEec6f5cvJ94hPTPuTF4dE8Xm18XEfSxl
JC2FPkeWYHexgsBsB1BxW2kbsFrdU6Y5viUQzt6NJ3DwpHdsluUpR1+5sD79O2CB0ykoj1nB6jXO
caVdM6Ldr7Xf9gBZv9OsFcpTd0DLSt31aJjyjRiknL5KgQ22eKNL88D+KDQivKd1KUrtpgfKIEUx
vK1ew/IsYTWroPSt+Iu9kB2oChdA39wtJmdigSAaCsEinf27acda+hUvlgZFeEqS7y0HoK/FwmOW
MMYgkVJvhvDXLMIaCzx/gXZuiLmKbN/JBI6IK5nAF4Yp/h/qgWvWuZf/iBw9IYg+I5nAMylG3m2q
eZLhZtKK4yl6DdQ5wJvLKOQZVALX+EWVJ1j0HXVzq3pHyuqk4mWlYOTNBEMQXP77D6a4xjTUv+ll
jexoluD3LHsn4dE2BpRLMGAqR7VrBIUGWdsTxwVmju5d1cyR6rFTeoW+Enmi7NTwFyDmPr5149Ih
0Md/+11jvIWP0AR058FPcxjXeIJOObWjhtCVp8M7fd4HRSHSNbLPag/1wIkcXzhl+xFc5/4ESM+i
e2gI/IksSw/298nouePtxd3mTeG0N7voniNOeITLDBG/IqXAamyHpoHFiHRtKaxFmG3QCvPND6DE
VYdozSfdoI4oK+wDm8RSr+5TXf0/obQbuN/swhi3lftHtEa65Cfb9xA3upkbK2Ua+bb0He6gkGUI
mg9DM+WdGq7BHESoapzO5ktKy6BfxUPckciYkFK1fqGZzG8lrHb/fyikGqHwCQffBfRuxNOPPq2k
hmwrpMryedDIHQ/9BEs21ZqNBWK4jhkUvDlcilqNLRQuJoTMFDqPjSByB7jZMaVjLSuoLVHiHUjT
NSmCVylaZufMbdxJRcwU6MSqw4LUR8JNcaHYTrsPd6eBaZSI+s8ImKfMlSKrSKz+h9MOxOlbNNeE
8NO60PSncdf/zaStZiOCXagTkqcM9fCg01AED8Bk122S9x+9uZBQubi8jlLi6xBg3keZ1nRV81A1
rpqQuMGSfue8a3sOwXJCclR2sCPNef9ImsxfVB2naFlEXBUHCwHfP8AazA5fTc9OXC5GW/Mb3uK9
ywplCwLV3rzbI24Abj0Lz7bPr8CnMnQx/9tNnNj3rVKOzJ75dTVo7tYIr7pBj4hlUX1zWvPRjk8a
FKwM5ojhNMEp3UH+u5jlg+gzNHrkxjiYsJl0HapfOeugeRTckdkx4OMBRpSUz1WIKiSgv8ZF/k9L
jRGrUbEWVv6iOyuX2S2QFqksY4A5Iud9gFLLKUL8hOoN7gjKpocjD5LyZ2RowdMGtl/kw15yyMPU
7saXa4LmJkxwl/66LDhYdkybeRGKEuyTRQBSTdo5ChCYyAqwtiBQjpdGgSeeF0LkzBjKyieTBL0V
ET0f+a1pW8loF+Wld4dkPZ3nGKFSgVw8ew6XMOjhzhzYlgqaEZksW0J091EYPp4oEUVoIbU05BBL
cHGvuC7A5VwuqbpMVx4D93sEaUjvyLI2q/pwf4dsTEw7OkfNb7+Ssbb0DrtBAAWZUTev3YXpzcIy
7LIABrSI0vRcMH0/bfgo//bE1si7Gg0fRNQxFgherwQNoSIVXtVzvv/Q7j1hZNu/0g5FzHoezQf6
WsDeReKpq2KiUYeCfziUBsJQsTvcXVgG/6WUI7fwewH1ZDE/aYjL2KD2x35DTLxJxw9n/MAT2XkN
KDhnDYfBNx8IaKdG9ci59WMwN2uIC9VcQVsRLdZJUqR/jyNAoh+JZteH2f3MXJnBJQXni1jFVEcg
+/BAkUvp3eYAZGphHRFflYeJ38IOTUeTNX2r5f2I/q2fg0sLLPhC6EmSP+pRe1BcsrnJefpLWevS
gWwhYLiZoJVA59b8N3pmAeWlcyj8pP0IjBeOsQ8cbL51WwcgJiUjtoY+nGHk4tk0Tiz0ZU+bckre
qBi4yQ8nb/FBvPPyp9jn0/5u3VvsE35qhRiNhQXPE5L3LutaSTQ/paa/oeCcSOEM5vqieqW16Yg8
TF6Za4K43ioA0ijL0FqY1VLsMRiloBkf+cjtkFensWx8B7MktQFqQLOg5fuVNEKYAGoCPAE3NK6c
tZEpjYiCF11UvaMd1cF4aSkQdZ5ZI84tcO0VeUw8l3Sc3KtANj9X6OPXnPzQcA1KN08Tp8OoE7xg
g9D0ZSWNzqMNy79sqIrdf/czLbyrrGJopujEEVEtU90HpdHPzap94zw41Ftn5G4FWjvD36UDiew0
uWiG/D5UmwIDN2DDIclrmnO3G0VPZFXCKSFM3sJygf4dbdwaA1nxfuH5OwNpDUWBlZDteoUAabXP
xh8L0fCUkKu6SATt7ElwxYeWyuEJN2dPW6EHwz29BECKVB6HbbUaAHBpXe1XeC8c1WcehbGl3Anh
EJp6DyxKzPQx/TP5xbtuz7/BqOI6OTLnauWrKCKJMmZBcL+Bo77Mow91DOFmWiegS2YVZ2C3QT9d
MG4WYxTZu1pKfqiaSff4qZkHcvP+F5dLU7g9XnoKtrfJwaFRNSHRth9/EwdBkRg/0XIEjwVfP8WG
L8xOaNSZplvPjayhuw5Bm8p3PivrUzJd733Kgi2i/QKCA9gp3ytXCPuu5jCmxHlEUF9d7hku/DEO
DdpCTpXlNTqRRQbkIlHBu+Rpi6B1UV5G7G6e/QGYt9DKMKgGwPTgYNjXYZIoNZwjRhsSprLIwD6j
RyWfYIgYb4YwbO/ga3gQe3JXUrpfMAe6o9k1t+BiVmxeC6twAmf0d4paOIwph9y1+VtTpsCiiSVb
YxUDGENsMfkNySDYK+utPVcLIhDw63k8puQDW8bsKW5e1td0wTZtOiOieosZSmGwpLhSgHWF1sZe
Y1fS/5x87Lm2+usia/QrL0F64ynJtc0uVViT0T3+yFYCX7+/5QOqFLTPyYu5EXYdOB6/FAVWqBYB
Y0gEub83nSjTXVUOUBR2radORAfILQCQ7uJ0zXcPd8UTkQl4+60yqpsoDRRUgk0lkx/W9CdKklnI
AB4Nvsz48jb2Jq1jO1XBL3bbGUlgtPlGzNfNI0dVxfcqRc0PYQvKorFPwc8UYHjQLsFDlAB3pzcZ
iGmV6aA5EoQiMAw+/a4rlh93abkX19k6/P6vKtwskcR4BX4fIrVCFJErsl1uCpzYcE2L/PWHPwv5
qq5J2Z1HaCEK7UjyGyE1qNJb0gDxmQUuCN3AxT38lGgkV3xr2q5DEpTZJ61F3nfuPlMcLfAA3m+s
iLcGSL2hZezOA1TNVci7MUbWnd79xrCMLFQGxHLsMoN4XcVOZHEaBqO2VBjmsQZKmBBiKadjLJNG
3e3l5kXC0B1YSgLgkCW3uRSrLd/8cu7hGWre3E66blJaURdY/I01uMaGjIK95DSSXwhOG3VRg6Wx
pobK7FaQeF2/HlkaNSrORZDLvdgiWKewA1cyq+Pu7QG2VSgJisYCRWWgOi6GuK5RcwvWq18gSXDP
pFswmeTlcpTkNrKPRfIHuOlJMJ4MpNQVZW1rEAtVYY4BQV78Zw3Wfcn3JDKS16ctMJ9rURntPU6s
GIYyIgQSE+9NEodZSS4JB5EbCMl7ZU3dzLcesDidsyVh35RBq09WqmMeAX5vrg/ScjRxDAnmOFnD
HVXqzFZk5gVUKf/pdxuUMU/tlNgK7l3SRr02V7W5Pvh/AzqRBkxbJPyDaYLUJ80Vm/GrPsckO8zv
bf4zvvcObbi7uy6ixw9VvSdolWq+8QMLLsvQSYjuqFkJJxtTXIQhnz+fDFwLtsnSEmkXpR7giXNl
VJTJRut3RWgLPUJkMhY88ln8wOvpkiTZCQXQoqiKJ5gLps2KDRJzVQ9X5/+mo/7kERHnS6Y0GvUv
Ct2UqG7E0UYd3YU//Q1caILsp35UIn5+DwhakpgCu33wypgviK2CtbfiK/Vt0QLv6I0e1yyMBk1S
tknoWe/kNfS0O2ASFu3ViS8J2ILMPpc/2/TMp50W8ycFi+J1F/gfcDD21qAIieGSOunnckzE/UY/
6hXnvS+FW8IfBtvS4XZQMwBu4XGv+aLGcdANH7euqCEGMhcSDTGJmMehh1g1mWhT/abfaGc/yPbu
P2bhSFJUZPJoEbEsYofhdXvCEY4Sw2vxhRWH6xSKpG4IXwmN/jLAD0Ml19bC1ZPggtndlP49P9Kz
9GuHnNsb3AjCAreryYtUPay1vOkjmZ8F5LNyekKEZr7D6IkwzUAZZgRgzNiyfhss/7yUbeeTL/eJ
Hn6CLQNYnq6+HBICVchU8o9lsSltmr38TQrpTMoS6exiQYqKxgeSYCxSpI4BQW53Q+C1YEMqCyyu
m9txNEJtVBhOE5EznBt765vhbzYEXw24qeJ7NBAV9tvS6en2oGJKGaQjBGuJSukdlrv5URdgnm//
fud4LsJSxv5rvH6oOi6UWMYb7KusyCTnxfrUKggvdWLupo3Ki3ATMNMGIWSoOHxA3e7iAwvxtzll
SV0vOgX4cZJ/jHbzPXFSqAjS5TPy/53MNmyZ68QPlt5hGvC48CQVvEupzMs8YgJD9JYVUJxhwbrR
KRCGr9tgZEKnrayexeNaqfxF3PP7aibp6dyO9ACpotwg+DJRgsXW8q4jFMWYmhiUIWE0h+bnTNwe
24oq4WvJbRyN15ElP5r1FTn1ip+KOQKCf2Oc8fajfWM5ItpzfjF83iVXhM7/xB5O9p3sr4ZALHCS
Ps0c3gLJhBA5KmlHc1DSw02P/NOFuv++og/l/yDMxm/hmkBDWeVNMdadAtCFdHCycjBvIIwU4HjR
ZPv7jq2FwUB7YAEE3g2dbxR/M4APPN3s6dQaLYs6IqwDXrpZIeyVpxaqG/FpkcpVPdL7e/ewsfAP
hPwBsoUHXaQSpn46/Pc0egnQkTqTPIUnzgiiAfTS4R1W+PY7EXBiLndFR3agE8wSny0EJbRbBvoB
CXL5ObgAQFHc6wdz08Cc6euxrK86SoQjZo2rNRj7etNQCjP5T4SUfZLpUxz/05cqT6r0vsEOsW5c
MhsbagZElZOoJogCh1raPrzjhB+yHZkfeeEpfKvPrrE7WxqFifmhytN2iiN2cPRbFgewev12s73F
10vCwZjp7376+QT3Isnybcu42B+IgqnfVS+5SardHPHufE3jhSccD4+qO/C3/JBl2gkA6M8RJsVK
4mAjqQM7FWz7k8vKR7BeZQ52K6qH0j3DRVy8ZPng54QFGRzKR5LChpprCEuQ5sKh/LdHAj+4LefY
YwHoPycZJbQX61vcclBo+xWpBtgtIGc+kIHHGwreCzVe8FT+gYCDxXbDdmC33fAtvJnC9UryCTKk
Um4R63a7d5C6AmtyzMolGJn1alKmAl7+g7IYr08chsdXw5Ls8QbeP7onudLNjobEZFoDdRvts2Jj
JupDCsHJ/gyneyVNy9Nv2b4F4h/sZUzjaf/2ylqhMtH8FgtF60uDCohVxzoNZqQf6CHkIJHUkxHt
75KyVeFEu5X5pJH7DTlwLDuVIy2g5+xD86yd6+G6f0BVqPVyvOtvR5u4D+tpvWiuvynQNWNLUyZF
C2IdxXGxyOs7SnzTWKhPjLsvY+xy3re6/btS0IgCtAb9PR/vb447BxWxx0f3QNb6/YLwh0S79gQy
oQybqNazk12bFhTED+x0Wvst4IsKnuXb2+SNVTSGsAY1pGgZ7X6/630ytuSZGXOzWFgnRR+UkPz0
hejy+jC+OwYPF0iagC8YBgtGEsbsOxpXSoc1paabpsVCQ+JTzAZ4Kg+NRjHxOG+MfZ25VIfP75mZ
5TYx9XTuJuGEeVI9KtjnWOBGYlIJb/6/wKvRi9h8BuHlamu+sEocLoFug4ZlEF37pCXo5bhVWrbs
DimqpI5qZjvnvWKXDdKpE1N++4rHrLVoMiMIzD33SyYx6IWkynC+j+vSS75j+938li60FOv6g6Yx
NIUjO3zqF8eHOhnZGFNT7vuBce7W8ECfWjsxEvLM4VMR81bcbKWz4Pf/MN2+MgWlGLtiDow2zwhp
DUEcr11jaNnAdqlLuJmiBGlQ5LN1l9XZ4IGbGLYEIfI5U+fDqeGdQj/JpFvSiRiUN0yLSa6IzoQy
3eQ23Xghe3xxzWTVNQAAUe93lDkCLpwh21hu/pYcy0+wdyMDkjBkCU6hq/6tDSEr8TetD0iThmSD
c85LZgBZ15AaKKYpbTpIsoOwzqeT9sMnclr14v/W80c6zc1qmssGGuA9HE/mufDe0uGOKwMEZdnu
3f2GJhmxmjotCO8n6lVn2ohRwOt6qTCLhthWeHnyYqorPDs1eNoI38IA88YAw850dkUCDLuBZLlp
XpH1c4MPeb4iqICBepiY2PRJl7pTHgCsBP8xS3adG8lgXz1ikg9dObOFJb++VkBNwQb1wSyuOdFu
rvf95GcUpe+UGm6dEOI/Ih6eWWMFDrUUmAaboq2OreHU5u6YVAggy0l0F5IDr4n3mf6OFLrmKKLF
QnHkByG5R/QR6Am1eG7BdsoS5T3GnRiCdxrRfvGP/8K0qTSyz28wyWaDUxX1wmXqvR6aKSK4kMaS
qPqAPGLDyxVjG/ImNlszLvrC8nj2E2bGTtID49YHEWxOKhPGSd/M7+s98rT8lSPdygV6tQWyh0FU
igT+hquBD4IGo+eje/4JkNwkwAem0PgTh/Pl3NluW2d5l9Eckj6HluQaFzHMKEOk0ho5MGJAFEvA
Jbd7tWNzVTZbPkQQS1UgRhRKJkBO3ruUHuB6Hc5JC8MA/PPrzv9/o+IgzIsI9JIemRvnJGzOLq2g
/uIe1JXnfLuVh/IxGNawg+lEpVpCkLi2WKR1J0zuq6knDmvgTsClMGLYLrbl8SMafsqlcmSmtqju
AiV29uSIzxmGCQ+9ki5xtJpbz5ce2a2YnDiHOBAUZy6ueqxUjVtJL6dSdDpFT8Ngv6qmVgmlnnfe
oFPxJ8ul7y3nLJHT93aWmcRmVELYSzxu50jSapKgSODHvSuTQx98Wba8S/adArTslocEj6KOYK/3
p9KXEB+7+qNA0BVY/vviA4E3KB+OwCDwVHUsK1R9BbmSNFfyDpnEzjerNWf6z8PlbpHAfAmH1W74
OZGBoLRxZWqBYlqaxc3uPHBX8ZbR1v6CCQQynchhi5P+HLXB/J3dsumxEs9jbo9gPILhoyaLHBxf
0PTZy/9L6GgoroXR2ghv5mRxSVolnCLolHg0noVhOKcMMN88bMUQLiQleSBbNegWmYoZcWWAUobg
G9lVzVyv/Q0ftD2uFSmcQ7zFSDNQn1QCPyzE+j8mLfTB5Vg28xCE5EnfpQfVIm7UYZnWWwoodK4W
3/4p9aggcWDB81Ib+RMMwQezZjjKUhtvotYoPcr8m0lzemaC5PjiD2cyrmy77nOBphaibN29poLn
5d1PMipL23HefOI8ysulS9lujqb+geivuV+JPOzz2GbZqoKoYQQ3o95ErTCPRI7+5Hw2fsQcqxDr
Oq55/ftOK+OkUR8tV/HzAabDuzz/0NlEjkcM2Ke2XVAF2a/IVbLC78lG7da9KhYN0ezUvtbRHnRw
FvedVW6nilLhzCe0ja3qsvIkgX+/FGTsZHDGr68hYsTOkw3JgxOpHM+4TpK6UQlFRs2TGiOo09nf
RFzxx9unWIa4Dao73QypdTpJR0VOut83b3efxsZkqhg/BrFceiOAFhr1sRSb+5/DXMht/MTUuHOm
31s102QfuhbxAAHbL8KgYIRs/G4H7ZkLQ7cSHBGV6msH8C2xqO9LsBiMdI99dKxQJncZ+cW6qNJ3
Wuj1fBTuNdw+2DkxrgNFniSh+/1PVIOf0bRniGpkEnJNTSkmaHyqF0RBUgTrQBznK6xgfIhKWkQE
y/+xmVZ/yyNwv1OZdI/vhb22jKlLQW1vsQ3r/oG0HPpbdBCpxfSXiOzHY87Z3SVwJGe54RdqlMo5
S2w4IAobx2qId2Jrz+2xP7B2qgkSxaOSrLn2TUpaeOjo3jDaoZL2aoJAk6idiFtoWkSiUoGrFZ5d
/FQPfUl7bw/RxDuntkqywgYmWWset9JB7GAdFGp/qpAcD+VSxvWecZJWo8ZlKZnYIZaZQ9xYuN1f
MaiGj2A1xraZ6N6HvUvvRuByGVHtEjrBnlCsDbcOLZP0nfx1r/LKylWGXsI1A+t6X5Ba18yyxIiZ
2jfJA4Rh1WoaWPCSNOJvgyUPDbzkm1Dz+lM96Spi0wOzNQ7wwVNSfg/QOUOoAxxVit7qu6hhmqEv
P4UmjqE5WcUxhpZVowtjEBILrwbeIZVCUFVk+OzKyDZXyAKUbfij85XVy+KODMA2eFbuya9C5nqQ
gI96WqQl83Mxd1bwqnPIlFiEU4yzzIl+Iq46OZC3/nDvOHOaWG1cqHpKesqdAqi3MqcwpF1K2BxA
FuJZzCh6rJrwo5uBw3YNV6nLBhgX6W5PgqBLXVQ+/VgQQ0wwItVvO2uu5GFwrAMzlOP8gzoTbKjs
1dmQmoTf+sfJ9KLf0Zm7U6IabMXu3b0AlaaOHWyThWkmmZ3H33NjQ1vlAiT3OPtHMdd4YIvbc7O7
lD0uHSej9B/EEhPRWw6zhdflTqCloXcSJnhsxw4sWBHWw5Y4U6bgjYgJJH0ICAQehbX/aLRJ9QHg
asE9+hw0E875z2D91OQgnDq/h0otjnDRiCVBgPTVggE2RGnAi+W0BLlMfDMEUU05dfobdDMD0JyN
bTaX5DC4dz7yH5C9VIi7baNPA1eEjzmhcqG3MVHErXUf0uLKEpzQvF0GOvWZQey4dw8U8+19lGPV
+py9Bsx/nHT7yTKywKOwp+idcg80Of4fpRZQ+Z3zZcQ1t9K9zKaAibd6agtxyZ/Eq1EqS/XCP9WI
h59Cf7AqX0/aY4PdYnyfJMCY+witu4KboZor7crcITRPK0Wqy0Q6VmKTAaaR677uwjgVGEPX7YsA
x+iO66cQeJnX1ZHeeMU78DCOsg+10fCSSuWSKHTjM58/nrPgiLx4yUSnOLrykM0M5gYiUWREqNQU
T/uXO35AwJmYcfKXyBTkf0583PQpWOnHIMyuEBCwgYgtq9Nj3NvffqhViSx+P1fHHNz3kUji9AUy
aKaLphmnbu/Zr0DqnoIf+5UIavKiG14hSyvZQ5brGYWrNQQ1w9FqHuoc7SZF+TxFK0MHL170G1ii
LaTSCFcko32CttP73JGJAiNR9s4HBDMJ6KPcpSrPBIBq0trK6gjq0gWOW3bXK2d+oGR1I63J/Kr4
1SXuDLC9annOJHrkOKraBH8bfslPe+d3srB3Btd8JMFiStF9zW28enJ8n5HnadOfvT+9DNxkwnMN
DBe/l/JzfI9gn8Cp2ZlNKtxrD0eIkZo7x3vkyEwpfHpeElUY8s+FaYEY0HeYsJVSVwtWwb7yAfrL
1JiTKZDx5EWI0loRXorb4oXOwDZUtnuzk6kJplkpN3ny9MMUtd6izNz0bIFbdN2zkl0vzAHsZOFo
jZ5PIyUGiAWGb+pR3riOmDfdH0RK6oJ2NL26LIV2irrMqyGjRCJZIb8XC8W02EgjiS98Lmfx+mXO
QdODxWx0ynlLNaDKUg1pKJeUM6L5oxVnL5+wFfTCe//jy/o+5fi/bik0vLx6jbRkIGpLGp9XsdcT
npUoxrqv6mg5m2CssL0veUUo6BOw8PzkWB1zB51/oHRjF03ZRGV4AFcO+5H8bfNew2aBYs6uqgh7
UGEj+m4LKa0/pBr5PEoqFBtZHneOThTEwA24h1t/vf4JSJfu2ManzH1Mtvy+DhSbB+jr1pQcdeHc
VBHiSpRd85uiokM0w5OdRH8Pxi8f2r0+IdekpHQlmP0MlhrS13UW0Nr8AlhlCVB7vkY177jTQWur
NCN/rqWNvxngaPyrm6w49K+V0fdwnNGaIqqhimgfI6dWAkh1JuD7V7BtsSqHzngGVG3reYV90+00
H3atTSKowRqBs/wwRldRTUTPZO+5vkD+oXhZbOG9n2OYEzZ8FnXzJKz1l0VCqCxQeQ/zwYPmVH0Z
4cIK83EF+fJkug3nDy6wYZ3z6+DfBHG8IjuER8SAA5zGGqbOgbU+C4fItK+tm+kJpfzt2NnG7qHA
KXGyG5GN0mgnpH1GoZLtGjGQKmd7hIOxAoE8tbr+6MetXgoVjjlW0ZKiGBXlmo7nYiyDPeCQdfLt
f1DyN6ahZboV1D+3oYbnyYf0WhgixCJ51Hpi5cqB9IBv0w8NODao1JyAqL6kVn9m7JQv2ZjoQqmY
7rzisFhkmnapE0JMtAwc0zE3NNoq9nKL4voHaONT4pzB116Y5uWeLevZG9BPB6R0ffiHpRfjNSPY
5PpqbiLeq2QN8V5lYtI25i1prcTD/nLSlBdAF9h1Ev5+bOrBoZw4mgddOpU7MrNgDDSzaeqN7n2t
DNAO06jrafkD4KjmFJcmc4B2Z2Q5JoUoNY7ShbxN7vO8mFIYhB+dbWUq+fseiX4CGiKeYFQ3diZn
99xN6cobqFzMlb0I07dyZ4oPZ/j6LsKAzMx9znOMhJjIQyOZWu5v9vY2rN+Zn4Mc7gip9iNC090L
3+9gtrpBj1rVcOMHdzttR8E+UZT+yUWoh76wy6BGE3Y7xw8YkcDZ7Nb/ssYO2rltV8Svh3UEduy2
1aKDONJy/0j2NRBIRmHP2uyTAZxUZL/LR+S7Qb4OWpoRvE6ZdHcTu1d3Luc3fba8gP5yZh6MHUrn
QGQGKq0jAc0LEGqobWFKe9ZhF/LxDVDJCvwcOi0pdrfTI7+OWEHMklb9MhLURskpyKohn7NGD07S
wsa79M4T+QkVm6RunoRFzKYd5MX/EM7FwKw7vQhIxqHrF911DEmPQPlpa1BVe/OTYb99YhwaYf6K
BRCUgEKyVoB1ZJB8juKTAwgQL+LqOglR660oLYeu12qkktF2S4B0CiV7aB62qJn5UuAqeLBGgNP/
+ryCAZuCwWOnAOlij1dM2etl8elwnoyrt9CajfmHOlH2OEn9iwUm1ayxqq45F3t3EbqnECnUDXTp
8biKIFFhvVdGna/DevuUUF10q40NUKvA03PHpWVUPLi/TaKCSEEHHf2SY84KdDDoAcR0zGvbh9Lc
ufL4Hw0SixwpHv0J1xjRvjZ8Y40TuhnpjWOiXbg6f0xJBjEGvhoDnU6IteSTDRxmZsVBlP+YNLMy
4wwTNCnyY8YOWcsl3WqIQvBc7a1pTBB4RKxE7FlBYCI9Q1BGdnCMMYW8472R4olxl/nRfPNJI1Ao
AoXzzVuUAgpF4QAKTLmHiWzWgjfPNP7/h2CvQurXmCkX3i7xfbU8OmX004eE8s2dUW+4yQsEuyp6
R6iGmdazbo1TSQz33in62jg0/ZISOg06UW26rMX9Cejy+Yk39mD8IY7i0NdSxefRjbWcGyRNS6eV
X1Ql3pjMHyTqHTSZ5p9kkXNiExut0gL4kNXzrZ+5vyphzwrl0cfmfEMwIKF+tL3xGfRQNUqCQTJ8
lu5FmMVzO39NT4PEBgUlJqpMl3MWFqM7IRD8b2Tdj/jVruaF+Pa0JjAiUvVXPJg3sPHatADBr1SH
SU2jI72PDxjtQ+rsQMB5ICHnBO5xz9iyIP/QXgMvfzcbDshNGsyWFSFFtH3ZbJgRKD0TfsqkVDs/
vIG9S4iQhuupQRBJj7lHyZWHxPM6HYHoCbzhFmBG3iMjkup24gqyceSZfkagjkYS7s4yJy98NINT
84Pnfdzsme8QDggnm0IIiI65Bfn8Yah3hGzKd44Ioxds6B+glx1zLe22/vzhA7vuns3w4ovz7Kxg
XhjnVvArdDjJxw6WCkzOMNcz69Vp8AJS2187E0t8kJ1QRkqpZeGf4f085mwqwW6dHlq30gC4hJGi
SMbkzj2MtSJgLIyLe3nOy92O5yLGN02ur/0y/HyRI+zOLi1sUXn7EC/a+MU0wR4gGQ85xitEDVh1
iXUKlj9Ru6JkrDcPC5gwQGXq+9ZQww1D7qRhj9ZfsNjew4uCjWAjoegIMwsRhHjAHNxPjJMkK77Y
Ji3jbO90dszuhMfLBWATVzG7y/Tol1ndRi7Hl873B+YChwKRERmuOFlfrD7y2J3tXk/J1ckV81PR
J5H5/7U2OH8sfgUGWZyATuMH5fmVW5hFzCtTf6H2OqU6hBMtJMFWVZwn1GZY4xSj2poaWOGJQELK
sO9BKDUDn/6ukUFlOeYrXuMvcQ/5MJ7z+q4x1e8VNB+XkA+Ow3qh/iprR97Lv03HRzBylknKli6n
OR232bc0on9W79dtIfudbB+28AnANcEZEbT2mb250Bbuuq3QFrknaHFpnhPr6Oro179kwQrAT9jE
9jdoestEahGLUUa7xhPriGdArHAOa3vzS4rldpGSzV80nEgKg6hge7C4aLXijxcF0H6RjBM0sHI1
8RXBm/q03CR6atIeWmTwPxQ6d9U9omAoCnqaofgHQEeuiPGwb/P2cynIZDo9iQ47F7s6GXqJZaHP
d3IwBdz2yrTpCkjsfMb5CAwBnmlXrT/tGbuMur1dovBpA84yMDbRNmRuaZFw09+TgrkkEzvmJ5g4
0zWHaMMZXXlUUnxvljB30KYoO7ak3iXIGlSZuHL82aG4AkANUXoRoZt3nma79u/eOPwLIODmF8SW
aNwBnB9+nZGdpsrrAgIhmxefyYlv0gHA/daGaXOaOCfUQ1YY2G1i22VR8H7Jdy8kHoYtMuVvmaSD
trq1vH+/W6cdOGZhltWaZ5k+Jaej+0RROI5hI4vYWk7zCCwz4vBegYpQvgc2wA7Qtv0yjenOTJg2
HeqwvPbglwsaBVJUwDty38QDbV8ul5U/5ZtOfdfjQKhN814JvzGEL62gekB8eyjUX9DopbCo/QuT
YF0LxoZp1tlY/CooRjocjoXF743AkuyJ5cDjQK3dccoorVccmRqLgv8+TeF9WOCfuHNP34ts5ogb
bwT+E99gkzgT/Enfq9sf82TCzRUt9mr3+VFEOVMm6Q+lR3SgBJi1+cbBBFXbb+soUnNjm/rtaBu6
/S8LJtEbHesOLYyloT9x8TCnK1d14GejNNFUVL6Uu9AKh7pxZI+/Ub48ZuqEBzjhRUO0PDpwmtYO
Z1lK6Za7XpFSTeL3t3+7besMuz99XIEVI2/ega3iFG5HmXlg1V6eMmrnQRcyyB1jPxRAtsZU/8Mc
QEcPiGSaMspx7rCofaoAAQf+MAfqQf9Ytw3NJBCQLVXanNeuAqMryXgfn6TeZW3cBx9O6J+sgVt8
5qutwE2HssR4ZRekHanWJCxxR3SAnmMGuJo/UjvoF08Cegup9nuDuHTV/WUIAQNU4eGCm5BRkLby
fmBe8RO1C1wAvK1PE00Qt+8Fa8iUiPFUq5hZ7zrtGYrpVKm6ciAyxLTfrG+n/fUtyi0/l2+jL3DK
oeoNiUPXyi6/CYUUEZ1jJJOSR6CQwbfIz9UjNYybfKjQ0+d4i69qgIPZ77tx3xHOmMvFO47Luu7X
MFMVUl+ViZcjS/tNso5JQ0mr8Kz0b5bvzPE7PQOl4DhsMr1qh4hdxIOwAZaRQ7T+4qfQYst84ftj
1K/oTkvRjLCo9ODrkUTWjluIP8OzRz1T2o+08kfqSwQIqYsagep/NGQ6GItLlvIRH7y5OT8zLj/C
qAX0pJbg9ey4fUAmsLBeKgPdXS10tH1CehBnY7hyCCJZDPWi+BNq9HtTzekw0j8h/TVYBTxqigsN
sc/AhGhhH+qfL5vs2n8rP3cTJ94YIjD9T0uLKNiLBbpxP7Z8qV3md4I5GvqAkBqzXZU+fEoE81Jx
oktArv2aLSu6XdgZJ2U/FmRWzDB7YbNVyIaQBxNfzYdS6h7L1RnX308vGhbro/nt1aMEYl5QMA/u
IRMsKKMeAYb1H5XtWP4jdApbor8Y28DidfduGi9Gpr1+ixq1erT7/HfKmqRZa8VLAezNW57tfyzn
ELx9DF6P1hBdBs8A63Du1PR4HDtz5RH/mJLneBFw98iJ6SSlaZ9o7lS81tF5jG0aGwyBNcQkDrLU
hn4zpVQBShUfgX/e1/L00rCtWKqVlWstwl6+XzmuS6y6VhRdTZxuzuZJb/bMRJm715MuKPbYj21k
O/y6X+M1S8AHo1Bf5cVw79UYyX7RACDueFXl89la1iZ9wNdYQr0PUCTqCsHnCgkbiI0/DXKkdoI4
jaIBFosGiTpx1iJ+b4NMTRT0EBQxHT+Y6y07VzEh+GnhDNsF5bFOF8y7u2XgvbH7ejIVGyH/7/Ru
Eml/WPahPaU6ExGotdz8xb/Zt4I7XfS5drLzZ20xbm9tOznHJmFBkjelzR5TVHul4gj6GXHUiWVt
Hql1ZrdOITf9Vt3ggE1sqMAYLT23svodkRHdXEqL5tOO96qiGKlNVMhXMaiAQaiFdRFD97uHSnrI
FyX3G2ibbZ5K9ggjEzBUaJsXFIQCIvlfr8+ggS4mUDG+0/WnJWBEXVMJptqajUvTYL4hvlSxzDu+
WaoblQaV62FFw/SMIioHVG3hrBygQ1G9NO03QfdooXY6kpCbK6hEKFnpC4VDT53lzGQbjWh4UoO6
0HHfrg7Sl9mm0knXhfdawU81FG+SOBbU6yr3vQgdtRmG2eDW344nBKqEPQeveve0RNIarhXGmzXB
zGFCpp9BJGQ12lFOpYl4Jeq1l55W6dOobYuzi7gkh39vvgDoJnH2oUQdk5Nqmn3DWSAjBdC/bNWm
iOFGoHZzDOjysxBabdBm3MzSNg+24ynr0OhsNvy8EYIo5jwEYZF/Lgpi8R4B6rxqew1jiCWo4d2Q
+FCG6JAyUpw/xHwPcCsTI+gtbnfUoSeKj71QUvn0n4ePHnEgn8bcG4zlQFiSCqa2jCv+Ni9UbjHT
wthuk0fBNBw3UvbT//+P/KWRofDK/7pKBjctnYhx/3OcJ5FxC2/7THgpm0YK1nTiAZ6Z1JG866g+
CeAbjxCeNnLLs05kAJGSD28m9WtITmTmGgEwP6l7x4sa8hv1zXDBxJqGNSMXzXQK3unfweJVtybR
D882i/MIE9Wxt3bfbSVnJ7NVc0LnniO1lfPaFaEsw007FFKPvIEm+TWwNcbqn9nMEzas1qEyTQ6b
vkoLxffMDaRTJRwTHNqnYSrUTVVx/0Bfs05RR8yhD5uNICuTxFxy7qrbckBRh0Z8COInOULn4h28
QTlHwmdMVzXLCBF1MvsfWqk8Ty1O75TeYJ7++J+G7QxDJ91hf5eu2k4rL76j5CDSacJQdGTj8Pbo
b00TW4lPlsfuASADJKTlLpzSJS0SQ7/8IX3eH6vDafkRwiUO0+KNjVx7h39Ph/Zv81BCZeRxdsdG
ObAAMvSf7sJhbNOFqYB34cUomcZkb57yOLDnCePnZRyk9zX5bpx/2MhCA6gXxuR4Wz5PRws+XYBV
f3x3dtuzkY/V5YBwWTzhDWIPrvoAZR+0lsNTgPkACtznnp1u04TdGvZAvgRc+iPgcwZUpn/j02Aa
iHSTi0wr3WEQrKPUqAh1J5CsLuB8oGeuHU06NLpNJouKmgti80bsobIEXD0tBR9GJ7DO2rGoTxwg
j/MnD9GU7glGhIu8LrCBq4pxXkB7jUn9UAEOe/TTygYKNIh30Mw2NUr6e3nfSpIB8A8Bzn4vnaWc
zYALJJAhSt6d3f+XQClqLp5+c9716FQe8SEzyR6fT+xWfhWaECl7bv67/uG+he+XNMQ7zNnkr64o
juXeZUBVAoUo26gjB0fSomn/85Sv2B7E0piHiwJ1G1K/AG43bQvkdI/DiN1lPMoBbFEVFDOqbQhI
I8vyzMDADzAMaRf1GDpDUXkyQg2ZlUQEMzew2XHXQdyS2um82BVi8muo6NSJ9YauEpCUsFdbsI5r
d/9keELZpcUCldk+5kCsT2LEblK6vK4SzdDPuvAWdGV6xodhgr/nJIzzgTFRDIFQa3vgMh6z3/Pu
nP2AxQGODnDxyg5oTBjPF1o2+mUuT040OKjb+YVXMJy/U9wKI09uYiRsPqKpZPwB8IQB64a0APQM
jXhFxNXbJvVJbbkjdjwjeDnCjmPBszytb6DTaFnScTHeyEc8zO8woWVCb4O82pcXspn1KX/DQzCB
joDW7JcqLDtjGo2ePqCpmxG1IYiIYRC04k4EsPwBDr1ZCZYRhvVRVukOufArQL/pRV6FNqVBjtib
boFPrEmsWXqO9LfHP8UjI8sUEvNk38x1epyu+2Zy5AeAqsEF+wju0K/tkyH29w2Emss+hNhP3+ij
KadTV9JgKkkh6Kd/dfBg0cOPHUwZTNHn6D8/Eyva3Pjv7TMh995xjyYsEPfcuCezlvtg+1g8YG0Y
NVmEqh0Vppt3IDUCH2DpWYHd3CsC7lm7VzXOKW4cTcoXjLEomostp0e6YNkEj8XZjRisi6y4pGBS
ZYCzpY3UyKIuIZvSXPQczlriyDskYHzrwWSYZRkqWg0krRJuuh70SE7uNo791qDw3Avqh434EEMS
wuIXxNhBlX+4dUot5CtwMT0brqnrinpfIv5OICNw5Ei1Bh7GqL1yZczd9NiUpTVeY1dvDNUEoUgt
BG4OuMAXT5/EXWXF/lpBOjlWXJml299x1wtcxES/hG6L+q4aeso88m0h5+1zsV+tWv9OYjyd4LdS
47AXKDYEwf+P4y70sSmUfMDsC2Weenmh8AyfP7rpeg9QtajCMY2L0TZ6gLgt/snxSM7fI3oYDzeW
BFpYJGv9RqQZEkVZTh0cN8DXHFQUK2S/VoXIQhtgKrynZQNufmRjzB2b390jnXpwiS/sVMRoOZbA
jdM9gY4ifUYGQndI03ZPZ2LuCU/uYSElMNctSyKSzlQlEuQTnIB4h0o8ApsTtYI/qwmm7xc+Oo/G
8Mj2C6MCiyekJR3sXqjfmCQ3QihM/uNd5Xl0lmBS2nipFMyvbedZY7mUhMMli7/rtJ4GFaCI5hHq
3TZIS0jyOPPhYir3GC1cCruMbc+guLakquFx0BVybpU2RnHAmZp97VG7Cjkw4Rd+BJcOpbuxNRcf
aT2+1gwMwgNtMowFzduTke5GMwLgl5OGVb9XF4/mlHbpTgdgSYO4NPVcy0mGMIqcTenodnXhgpzZ
ey5Cw0m8e9+lLpaifS3tCZCqlPeKKMreu9Kvyc8/BYtX+UlSPedKlHCDcvStp70cEz4kTLJHXtPN
K42P3ktoLLRLx76/k1gmmqIRNTY5mLHDLvcjHFLiKEIKIh+cBWjKdBLxrdKf4js8E/xSfUvopnow
Tzg4v1pt81L5jENeEsY9x/Rd6T1dDMDUODZarcSVvQB8Cj22ySLWzv6rXiWVcavju0IpY2U8cRIp
kI+RyGJy63oH0ztKOVltrYxH+G7yfryGXrDewLBN4WKEp6dwSjnE8RWZhSSz01D4dig2MwDohfzD
b1hnPyyX673MNSu0i9CZKVPExL5ZAeZVYx3SzTZxmYCUWs8eHFuh58//qlCCC1lnJvwa0RFPOnPb
kdzauBnu11NDGaSn8QnaZgOKK2s0WoKttVW0Sg4hitWZ3JpYg600cDah+FyYB2ZlJPDsAIV4WiiO
UbCI3QnaLQYmGLBxEze6UC24nJ3qzYY1H+kpN/EKoaADI5AGqQvGmU9oEHCWm/8z48LYZz2cNe1M
tdDuP+isjp0retj1QHBvez5itmSPe9Oc2+sLd137yKudXpsXeFqkOA/tq2YDRHbrjhKcvGw2h9So
nTyl0PKNvafiL+5XPNri5c82K+E9GfOuoXlTpVtqDoE1g5OsyeFI9Izgm/eXzNsVWJJKOqqrdHCR
F2qRe3Bss67t0go3sWnFRp62FzKmtlx22gWJ8ZKN0snY4nSABW8Uvod/8yT0Rfj8AzrrYeLsOim3
2PJs34XWcQsyp/JHDSkHZlUc+kyKeXo75S0ytPUxy7XwPb1vITT2CaZJhNjahTJRAfwK4z9Iw95d
U3gaAc/idndF6PXGb84awR6FKf+xmjyRPZ4fg2se5C7TT2q0C02yoMCzi+rQ35qidMfJOlJIeFhD
bKb68r+HcBCG7SYnpyKY0XSR/HVRFY+g4j+edgNpEWNnnpSluqpYZ8Kaz9vqaC3Ke3S27tbiZpgT
o1+xpwAPxmFuq7nEN3dFlGPxeJGeAQeNlWiS7ERFQX80wyAzYsfJHcq7TtL1cW2dTwskGCYE+mwF
8LR9EDEaYZsBAfy5+Em1FI2xUCGdDBNsJmSWLwF1Gmvjj/iacFtTJfRIw4jxWrTCdeVwcmc/ZIJR
D6Fc0LpLmyUFwRGxAm3+jPxE38d0Yw7V/b8SyvYfGPXb2EaEksOPF/5NTx3PB/KisFGSd1v+gTef
ArJVdPsWyABZlamt6OChqQeeg3tUlfUr6JSclmgDV0KOCXhNya+Ecg2ZBBaKqJTjewhDW3VO9ZYJ
mKz0NS6LfnJB4twSrjjeBhDbazC0KwAhYeds5+7ypVCJ8C/zUwppxl3wtu72L8O9puI9Q1hn/Gvi
LJ974vflSwWWNUofU06tEJIPf4nOq5V6Butd2izBepLU9DekD0SannIre/EAO0rXjo+ZnEGgxFxv
cBaERhInnJ+4r/I2NyNCm09PV67BJY3uterDT/0Arv4nOlv1m2sj8aPvOmKklZTcW1l6OG1zBPjq
UBMcLF5NkiMrHCj25j2rR4s3g+NAupeZKrGBqzvmo04QcFT6W86RndKbiI7g/yFAXIub0wbZLlV4
MF4wCoCjueQSzEQHmVkz+jzYLBFwS3PYhhAReFctUW23AFQ6jR99j1/bjg4ewapniWDj+ycojhhq
KuFWbgmDPRcj6eTl6C59KjXAZKP/tGcFdNc69jeOJwzssvefrLa6i/jl+hbi8uiAx1l3BwEF1dtn
zXW7iVQ8fOT9b6D49CvrVLz4gPUufMRubBVdThsBfRD6WKfYmkSZlCs8A/gkRcPSy+BviMWp0ZrM
9XH+bO0Efjnxmyli5zKJiK8Bd47TOxBXO4cKZW3YqjVeUBK67UHUvik6m3+z3vSEEaxYWsmfHgRA
V1IXhACTZlZunn1akFyWN2lLhtvvEd6YPTHE11GKMSlobUSiBPOPwvrIa6VCkGoyJIIA3HI9hzRI
CtDGFzzKgIuJJCjjvi7pRphUyWf+jOhIZkG6uXZfwRlAKrgg8wu8rcWvIPdc6vBT3hmOq6/8hcH9
+xMqy/+kgAL99FBMYRiNubpUqIVMw1BRNdha+EVPEsTg4n0p3kOL0kZO8RbvrLEpbyKGPyCsZSzd
sECNTG/xLUS39eMPrPiiezWpVk+/guUVvQ6u4Zied9rwPRt0dmx5qUMkr7e/3WftAkCYoPtJtVLY
0SUnLbgq5OqjzmNege7BD88JPSTpzSNZ4loE6WxIPwQ/3suI+vqLaroIgWASNOMzhS8cNz47gGuE
w8J7dWe0JXQLUW4qdt7GnQBR0IWDhWkTd4g1BlaszcpZRFLkMwYmiA6s/PTKIeypj8Y8RMgIN0ru
bEos/C+Ch8SfFpmjKw75XiwQyJooEhpbMM3/waDslQjYFgVJQbvPDGAogOeiMuqRxk5jVyU9+V0y
L41psc1rDdR5weJku6zeIgD4Knu3Qp7Dp3fm1u3797pYADLheMYtj9AXLe3EDCLSGZYItNKcZod9
hQdtiA9OHvLMuQ6OsnKvzndCZhmIRH/ZsRcefzAkLq2ojHifUoBD3nu70WdAw0vR9Ec6vcUEZoqE
ZK7zXo4Exc0YGWfiFK+qEtcj8o95KyFqAIEQRH6T4c29tvwsCSvcWSAGVRqEHzus6284Nttfj064
Ivhci0+sgI9KGvgh5qraSpdek3kfP+/LTa/8/0TS5YmZuSpTBGqBhv/T1vpGxjMwx0gIC65fVuZC
apA/1Q3kK9HIBbjmmdZemUhGQ6daViveIu/BOddEH3coVpCY2AGQ8CcrphPdJsGR2wkGlZTFgyDk
6pRVMqJtwhtWDQ2w8OpUmPGSX6HgsoBqwYLGASR4gJQMiCcGTzd7oLaCfsGzRpEmepIwzGn/ahmo
KNOLSAy21DZQuMIhb3NaXwIoTc/tSAS0p9Mcj06cY3gsUKNogAFLXq2hCTvZ3K3tjocrQzcCDX13
sYssIuUyt4RmKA5KLvmX558kV5udlvQwDnVjiYW7DJXuk4CkU2rR2nFi1aWYkAm6Ax+KM0EwNwP3
+bKsAANSDnxOqbiRZYPS9MfTXhWNYUk2qXf33++bW1IDM9f7B5j86wfyMkslRobicNGEiH5ehxoS
ICh/tymm7Q2FiDnEeRcDAaD4BznSrsiwuBWGfX1kct07lGlugld0+idnis4d7mwi3kbttZL3POoO
aVbfKzCJyvRFo/uiUcQ8639i6MlNX2YnYTE23cyEPpeBVTGY+58UfHIXnmYClvck1ksXb4WEbf9i
RAcR+dsfZnoTg16MCR1iR4Q23AbwY9ZbJyDfaOKTAEz3N2nWx//C/5EJUWKUcc+sL/tfGikndcsl
fBXTkdOwP71ZCAroshay7JAWTonjvdp7sqplQ2r4fXINg2JamxT5G7tCPxqHOs66YjM7cB2GdnIa
o2SzI4FxOEmwQmqHC88zthsl0Wo5TFrrdoNHh3Xid9hiqLeEWn2jnGzHIqwBTPpGyrDQDOaCNwP2
5dtdAjJMAC2cmzBlLuM9FsajJ3DaaPgGV7Ut3xOkaTdwca1z9pChPlDYAfCmPZsZ3/DlAjYgoO9o
X8wnkkGPyPZEjeHIGeL11Tc3gLM73u70KEqIR0NeRgs/dqlPAJ7w1eqOtN0R8CPG3NsgzWh8lT4+
APK0MG+kJ1OIU0yws4gI1PWgf3eq4easgFGxfTiRIkSBkTUd3dbaSrbDh1dxVKCzwBRqui/cWgsI
/piJzrklmlBvyI4u2ggvgL3023qWBB4+q3rvoVfonEuMlEF6/rAtg4S3YetwZ4zCAkhhoSsTE1o1
ZsCg4+nfdJKG/EUxZ6UXrzQqxbIKONoALwFRWq5AbiAvWX0OhbVFpabX4hAna40a9Nwpo1lJyGdm
n7FzSrZvCkiOSIbohd0BltN1wo5Lrp3kdlhohBIDh9F2fk/TrpuJ56Gz+V4h1Do95+VD4sIjU6cu
wY5lUCilIfL1sQt08Jq8hHMcimyrqrrG1ELRSFSesrTNFZ9/cFUOjd3pFBQNRsh2mojS5o1XxhKJ
qI1SBU80v0vvxdArVlQyGaRrBLmEOqULc92cdS+Q9HfvNiYPVYaykae6Io/wHSWlNYEvxvKU1+KB
2hsL6vw7NWnMcQqqWRUrYTEU8T6rBzTHMHFSo0vqGZdqFHCN9m3uf8BI1shmXRZ3zlPTjEYVY3WR
C4EdhOSiK5FY2NDd224A49OpoPX6sWTc+1vWZCEc1LQcVb0/8GyyBbrYURMDoSSgcmUAmLXQIuKW
YA0aUjgEKnTFDWdfBH9FUP1zeyoY31fl4U2vvVPGI9dZ3MGB2jMd/csaEDEQPxomqU5R3SmZBGnw
efT4q/H7+sHlXE6KK64ySsSIpVcs7eNuTH3yefi3wty7N/YE5gW3vMqI8gsTNpBas5RB85BeIABF
D+J63xr//w8Ht20b64Ot/m3t6ys6h5XuEAp5djvhgYNac2T//6lGj3WekXpFWB8uKCye/m3KwvMA
Ae0HD4VHFGD62ElXVM4FW8ybJDs4sKPVoQzHicsNqjuwcvFf+wJIfOJ01A0ACZOs6c5++GcH8JR/
tNIlsuY8LDxBgZHLXySfMRHVLP3sadNSIQnvinaBeJLGsxK54QOcKBmb5ojJJvS2bhbGh8q7Q+wX
9faiNMlqN0ZaQx7sZVkwXkF38yX669HjH9W2b7DyykgXZ6qSxZ6cmH0n3XhIELwtJbu6Eta8kSxt
BuTTtqseX5Q6Lq85+mvfxTBVZn8fmgGP2nyw5IUu2gA50W6m/E/fBsHtbn8sVOGTDiMm2S2CkAtS
jWKCZEANrlkMh6kL9mCt6GYwN49M57fpKyVfN08YVXpDaZ7U/cwJJ8RhK7kGVQGRkC0dNbeJxLfz
kecQoBtCsbHnlCrRPsgkWShLeaodTctKahgHb5UNXXJuPep7FnpU10Aio5C5X6xDHZ/LOsxzQbX/
iVpXDxouv/48qYLOCgZ8oksfQmtI2YMH6RvivxaBs6+MkIcjBDI7VzjsUxhCEBgekyaff18CcT76
FfMoPv1ebOfLvvLszELggJ7SUbx6vbRHdwLgVa7espXtZ/6UPPCby3yieCN0KDrg0vc3Wqoj28BY
JDeV5Sdj16LDfIn6xGoIPoVVkIRp4sLOXlJPCpNAyp264eenj71rWoJ+xI+OwxOPpwdYB3CuO1jH
bDg1oIjaT4cHkI3TfeEmGypHVz1lijor1uvoPpyf5K4SdQMcNegVXGQcoJLAeRAurzbuZPiyEOkB
pj/tR0XDmbafVv9H+VSHQLnOQ+I4kNIwZmlAReiIqKjskpA4H1QPrljWdBLZu+LEkjHo8J3wMO7Y
Un2kQJpKhyiJOKmKDMfgS71pQiJCq1tYVKgI3ohg5ELChhzAwjL5UcAYesMv5kmyZoqAKbtNWiB9
mzB6U/oC6HZIvv9LRh9ezc9WOX874o7CgpfZ9K4E4WHINJ+E+jPOYfuoof52U9oC5JCuh9Vv6zSg
i0D4cAgDHnOJjUIUPhLlbiEvMQ8BHKLnmkj77rF6v3S9ARbKk8pKfwMqEgWSjOFSJnj1FzcWU7Vt
KthIL2SVCZ0RfTy8pX24IPZbVczUa6bYdddqX2sLafw0CJxYM/sehy78V2CT0RIKwtj5cUjXTnId
KYiYSE9MtdqYYe+pmNp0Et/j74hssnWULyer27yZsZwoEvAeA338z0P/aZHc1WmGaXECNLpzH+eX
pJODmRqq1Idb12NExs86up1WYeGAEF+oJmoZvW60SELOyMwPFj1ODZlvlMLcpYUIQ8t9j+JAb3aA
2wtLU3tzr2VGv+issEUdUj4pfTMpo5U9ClgBA63aI5zCIrZe0NJf8OxgVVGgVOTI5mON05xb+JYn
SJLsH9nf4efKV4iaPSFtKjSEKVNIxeJ7KtlwoFrkoscZ8IPf3LLNFti33jwSWPWC03HICaKCz7Fy
B74mZ8h3A4xVzh+J2Rp7BMq2w6dh3KiMFYeRZ2lXBC44t6FSFn5Doi9N9ULn2sWBQa5IzQWPgVpp
HU5Q3WgQCPu9zyPDpaZosl7//ORFDYxS/UO5Z7EkRKEaDnkAL7WSwQ/EqFabEjYbc+6AVlSmzVjk
WEepqVxwRpcrhgNiaqFadLYBTnukbTlpk+P6TLgiQ4JGqsbf4Hs8W4TETT+B6SxzqISe81Iwov3o
o1Zj+3jIGvEj0OHHs0K20A26NYARpS5YStCDl81gQQHvx9IcdeYPfH6CYtOs0HA/lGoirjEndBBe
9SKRFFn9LcI1dUYsuKCdlVIoLn86bALBF4Xx2+SI+UDQ1HI2s7BFyUIsYXgdiuYyJ7yZo3N5vqGe
SmIsq5H7QoCX+dqZvG565of44Q4POz/uMhaJRJJRRZmWT+iJGqB2u9vP4w6g5frmyZLoeaxT4rbC
2aA8dqOQ6H8COAHcRipieNF77HoQ18l8Rr50vIjMWmpI1/LmNara4t8dfIHA4NptpSb0tn/iNdi3
yi/5bnW2IB56woxSK5pxwNje7ESTVErDmou0GWES7Ujm5LR4iOe9+y9TAhxD+0uKEHgQ/DgKo63b
m5M5Oo0Nvf0nqtnZl7iTft1R1nXPfTgoigwFxqyM+HxgUgd1W+gN/0pR/QW4yw0g2MTfTXyENX1N
XOQUni7KIXQZbT7pe2mMyq6G8WbO7g9VG7OZjBaXKJqGRCgX8NoPVHj/c7pCmn8BzkOu7GlSFANr
HNEdM3FW8KcEGGfsho+UXYblgyt8djedgJdpreqVkHKA3b42AqJ6d2nWEezwsHIDgb/k4fxncsxh
wYXoKO/I9XZJV1b+vEO/WhFbby9u0LMSi4nHrtxmwe3KcLzDYKuePiTUezI2Gwvy9tJRuSiIjzA4
/aQzjIR97kA0dlJL7eU4NcyyTYLmSMT92lnIKi5et8wAqgzw6ila3LwCay9A7wXkpmaJVLWP/9An
it3ulMviB+UBhvYX1mqnUjEc88Bd+tzpeOd/zL25v5/z5nnHKthMUWZT13C2liAWoPRArMqtkcn7
M6lhlVJPdfGCNa2hxHDVoReaZL2GPKZlDdvPh8BhpcvyXlCnaHMfKOj9W+HKXtkoOEQztMH3NJHZ
wB72E8bwSVuOvCt3pwDSBhMKC7o7cCZbQZNPfaN1lR0KGQ3enHWJVKUEshFGpFwrXYgVWl/DK0CR
tcJC6O5WXsRGu0DUTCyZ91dd6FcFbjkOyDVJng23quSPpRWW5RQKG/hntzGAfXIfE6i3GJJKIpUQ
jCe4W9niNfwX/rrr/D6WIvVYy18gKe4DJQDsQ4FMTYykvCBCriytnle4ZlRP4PQdf2slbZnP6M2z
tRqtKsV4AOMr6bGnB9Z+0uPjl8Ao9dIDyLRIbYVX1ed0q9psl5C6QrVZN8jSzs12UHMN0bQPaAI1
eOmFI00MzsBDMZe5HK73G7S77KP9KsBSh+FawqbPLUfkSOb2TWRWB+zSMhpSU6YbMeSSBOrnlo3O
jGOIt6DTW+buUhJ6NMe0cquko+PnYNEXbiPN6V0gNoFROM48KQFEwnlrOpUsQbRtg1OuP76SwLFj
vXRqzCbNXsUJMLh3/4DMRi4GVfrUTEMmDTEzf8+Z2BbiUXRutnxRBUzYcu/zoFYxR8w/d4JiWWzd
gAfGlm5J6kE4oQeh2vqg57bNiX4d5mS7nNdD6EhHgiaCGtSCBKFigi1r6H34++I4dsJemSPN5Ht0
16v4wSxdf6pgU3Tig86H8scLw3OfPyCZKfZoTvwVAUE0fAZUynKS7l3QnpbRKOCG1aRbLuFdc7Gk
HuGK26SwOZ9iNahKMSFFoxVTM9JR7W/FJ9y0HkgTuM3kwgwYZNBaepbwaq+syDEuHxrwYRdbbDGr
kS+uNAEujkGLCGId4BFwd2m9lXBezk7azizH43L3qhP3K/vlObB27SsHhgiEHa53xxxkPv53l/+y
IyfrruWiFCnBN+SqEVv5qRw32YnhDDz8fHANJcAt+bYUg1CRmMe9AIurkpPGGwdEI2vXjFlgYTuP
HZhYeaAVr4pNPG1JtquTxGu/gtZkalMJOPwvoMIlsEb8Punpn4LBOpXzBlM9Ns2QjE5sak5Gr205
wM1SCMdFqnlo7I9qc3MURBGcnCRxmY/845gzxbsx6M6H8CglgmfjxuGN08K8kxUebS6Oxv1tWlht
+jnTYx3H1AzoKPQiFFKF7Gg8+hZEEZkesLkF13dfyxD15Gmkc+cQ3GCAfQ6NmG6ACP5SvpcpPlb0
EXE/Dzs8ZWRneu6fsrFX0C3H8op/5hvLAdvAtAug/RT2ePReBR894Ak0npaQWbDhhJvcB2S3oYx7
z2pi+jhgu+ve9ukUaDrD9JX1+YiFCvVouVFzSzRnaqygp5CP1UDD7ozMecdZgVm+LD2vizSP4k04
KMTW5vXkNoDca54SHmRdZS307pm3yC72dQpoQMleCSY8cKgozAFfxPiRgCF5O7CqxsuokYPJbg0o
FGhbbGVbtPX/DJP8k0zSBHYNWskR9yChbqSM0x72stZarB1+x8uFKPkg6KTqPtgv+L20WAllsNXP
MBcZ7tMiNod3hppUboNx/rF7BAFRxNnP5Y9Dq6O5/XXqSTOyYMYs2UYbkXKUJKlc3AQW9Msee5/I
d4Aq6U9xfhKnY/3PYT3gVwCYe6mKtw5LeYJaeQYzUKU+5lOVLLsSVUkVXXXpzKsNMcGSk72y0uov
yFpCk3a9TlnNIUxwDhVX3AJ/qgbaWQOfn0X2WVCLe2Q6jM48yuce2CJqt1TqDxYcB7Bi65MBrolB
SKU1PQlcHYvd6HXn4CCbNNWPFSIxbRiWNNAC7zFAnd5KpXD1tM3ZmFLy69pXnM+VYg8hZmw1YyMs
YUsmiIhhBdLj1eR0ma++o6KRRdH/C4pzUCCPeq8ICkHYSDVlSEmVSpzzcsqcv5c++ehdgnJiyO/B
xtHRS+smk+/aU0ZdID8GerVYMGHndp5g1K8n7YRIzGCqCW+WaBiEQyhIf5Eq+6nJAmnVvhEK+OZL
sRh+MXajoHmvv9tc/z0BP2GN3etTy7SmYj2ae//llJy4zKS+Ie3LToIh8LF8muWivL1WJuxNZ0eo
A83cN5YiA16MrIRzUh1+je2xf+MH71f9pk2Cbp9SxW8d+XM2wdkRIA0iJbGcmzrGRRbOcH2dAFlj
4WJV4bhqx6aAWMRGz58+Fgi293bAGIzOzVcrPOdVvNaIjp4QbuIPBQtCcyA23Byt8wCh23yEFzTJ
f4Z2mh07PcwArEz5JhcXBVd7+eSnEph6MYKQVJcyni+jatmNYJDP59PbGLd9/OIFpAhmkxUGCzOV
a0wAB5kiOTIiojD/Hcn9iI7r808okFW5Ig+Z70gqdoC/iSOKNYaRNQkbvBtLjbvWMvTpB03KgHwy
TddICs8DEGv59/9A8m0/MnMsQxFF3lzE1PMjEpKQmEggf66wDkXMsYH53anDXH1QE5AZ9FBdp4k8
joEkWeEXOAz/W71fJ8y2tIuU72PofXFOAhB2jPiLiRXeJGhQG6YeYomgtAaafQxQ8/4xU0jgEPjA
45u/enjgHt5FEHrUJdXfVNa6yqriXXimxxV1tKjxzBeTFk2IV6XE2HOo0P5msZD5xNQ17zAoiQDl
3Y1dEpOmIVIpHbcM9ZT3EY/mkuiraIyk76U+jYGmqa51RA5oDloUBnTI/Fky8HiTfMdSMJC/9ssP
0pSM2J4LB9bhb2dmwBpU9o+aBy2A3JIdG/pMQwZj4RSO44krPsS6c3R94bwsVMIVEqIw0OR6CVrF
IYEE/e+iLW6vS20fTlaWrEJYy6vY+ZHkNOFYv7FbMHlrL9LducqNt6em00Ir72fZcV4vlbSnmJ+3
sOVi1D2GeO80xpdnnNU67NsrgYlHzm6GHMoL6mj227ne+wPWbgprx5j97cdL1nG+AC5UamSrOLF/
yP7EYAypmhw4/bXe1WIFFMwDiVcjmkOPSc1u8mkGr8D4yJ0KbrVWLfV7dQdtnG9ammtxOiWhUYK3
CwBAM7GstNXYUZqGxoFMzoOtpRAevv4f3HZ6NiPC412eyu7rXgjYvm0U1LNw0RFBrkZ81OyhYgma
6IP/iplbmz7VsNBF9mxSxjTJsf9Lx0KzjP4Y6FXtf+sNpXu3WQnb0K5d2grA7JQmCYstXJHi4Vgb
H9myamCs6hmlPNNel+or6ZB9APtznLBDA6ZnEq+TleC44i0k6M281LNtc06VnPgT+1PkH8t1/kYi
TYPozkEmCePsQ6cnLOeAIiqkJYniK2Du1x70WB8Bz81gdjPqNjjyttkEgxQ0tpTnbSMgd2S9cTzr
HEeQNPzvRV/Olp5vnOoMmTAwmm1rDePYe6F7pPiCx/LWV7UG25ZGIsiHK3aE8NMimEvrA8N224eK
b8n0Kkh/2ODpFHK8pyE2NnId7VHmA4YDgbT0qNOFCNWcNsurlLHcelgcw61tQjcchtslvGr+UmDC
jufsGBpRCmrHR0nj+edvYCTKT9XeVQD19LnJ/CD67SAhd7bw0PQoTDA/Vmq6rFwe0QoI/ZSBxFDw
5pWWnK5Z2MAsh7cNKNY/+TnKNDHsgXvV+wXedRNwgnj3EDblQ+wFa+FIgPwlKTLeX0xab+zcEmrc
mYxZIcoAsbcjSEH4+hUM+0UvTQFGMG+yZ8AyjUEsO3JGaLgHMGvAjXTnLjie3V3WP+BU1aApkY57
nHYR/Vf0GDPeV9xEp2MsNZ3UzS6K6zpnwClNeJOzDH+6wTFdHKF9wf9flNgk0pjJe72t2HGiaeNT
J34OpYFpzauUqhNSDr4uOOmhBKwFAzeg9rqXR1ldPHZHe429cwTc4WFjx3IuE2IeIRkpZXNZnGAS
cWQcMOSdYZwS1S3LQlFgLOptJTxkm9BI6FV1ZAXtSzSEWRURVJWxERTMp3ck1KyFS0IoKnLZ3rF7
ABWL+NVO6+KrsSuUqW+OJoE15VhCfFG71cQbfBCY3OR3kv5LMqj3diLH8JcJoYyFfJ8L/+JJSmlj
qI458K9F1Isv9+S9ux/Qtm6pqSmIrqZGPXNKPYygOPNouoJK6vV8akl4/JO6T9v248E8/aCzNd7L
EIKcmeuIeHOz8qAw0YfzU7s33JqtC8AmpG0WDw71/lUthozU3wllaKy8KdihmMg0dhGqg5dLIT/u
uxCPqPUvvCV9Ojgl2mXKlPU+Rtdz7IJaMMH05a40DeYunpem+0Ja+AmjMfTkmE7C85G4MvoOhGWP
MfODX1Ss0DNmBfxBbPnh3pMdmoQxzRRv19A+6vBRzTdbXv9T6tyo4tKfRY3GPBh3C7mZKLqfHmF+
OjASbD/ZNfSxhxLOvovY+YOiXmicWBb/jr7FY/5hxoCzJZ/rijN9My3TlbkL5yOt+b6TbRulKam2
myDB5Mu0vrqkH4sFSAbm2+NGFm4Zo8qReeHAHdf5YzqpWTSHT+2mLG0FEgCqsTi1h35hcBVdtmOA
q3BAfEyI+rTxK8IdK2Ck4Yt9xfjskl6IwVCp2cIBWyZHy3TWUxVLY+MGxBWkxan73NTJXIjKQU0n
lIZ8jV7Mms3CTLd190yGaWdEG6SrPvmGAQLKdFIBlxWYhySjPkW3BPmMUCiq/g83gKDg5ZLnFMA3
T4p5DmVOsqZs2tYy9bu8N2lrFeNpnSA6Zvi+ZTASZcektYZxsxq1V73A7031emjX24AYsBa6TWfj
LyCoUgAuvlGSV/weT2Ow//PZKTlDVOrXKCAlJKTTpe+GwuzqkMmVtS486tm+1d3kQPjy/7+QDOMR
ri5I+T5Zw8oVAY4ta8sd5BzZJKm+40AvCzMRHb91q23XPxWoYpzn2JjlywVhTGUiIhraK6F0GlRQ
oohX/bI4s09n8y7/MGnRPZ3eCmjrOus2gPtINnlTuMdVwy/DTC6U4oNkgu1bKgi3CU8aqrJ605fa
O10LbaOCmk9WCeuOt8J1oTEF6w2v53tqGu/ZxxE4xa5+ckXKaY18+Is3cOk42+cxl84fFkn4BwNg
jlGn4/LqA+XvpJLNZz7+/zkaFP+zZX6o86H3oyOp4pL64LU3K0EORsW5cDoKirCTruUk0KBvXC64
1n426nyENnTK70OXJY1cuvz2YnbbA/3uNYZclAPiO1R3oUQe8vPfKSey66Jo23Roc4b/9YOXZywV
2afQlpAA92Mc2bTQlG2InBcl8gOEs/BlgOQHzcF4TbgQIz4h8iUs6TL6sYbT0dLCDOigSgi2UqfU
9hTmrOQMpO3AYb94QnhACCw1fhIBi0dQKyKiuS7Jk60SLYJlH0kGBrLIJmUIcEJWdZGlimJpQhmG
7SeDiW11aDoQQKuXlIb0GvnpYntzU5SlEltG4e7knps2X1Emyf/JKIE6RdHHL7tJRsmt9Vo5wFw3
KwYsBMQUgqDnZPR4uxjddzycX0Yue4Hi8yRbqr/8ZlUO6HgBckPAbO8vFuCAn1b7LJ85zYh4dGh9
NQrAylMJzJUao0b+3IXbqlUAJwP86oX9ehF3tPD9BhT7t7K6IGYGdE9yQyMwx6ksCeEvliPI83v5
EZKP+fvh1cNYuDmLzfd9Kmp9OsQnT+6jadTZdmcxIWpP4oJqKxPvXI/8g4Ty+95rq5koNucqUJpX
2QgEqZiqdgsX2sRrfiTjzXt02iumWzhWDfMAf+x7C3HYWlrxD921K4rjy7kDK4cAyJ6XEwJcV8SB
iEKcD/hADdrjh9pbsCVp/ygtOAKcsdDOjFTwUeRYkrPxmLdHq1WgXx9A3+k8MQpEf1gQ9wAcFtxf
uQbuvcAmjusPvFsb4l1DAXoqDhTdKD5MSzJMYIhTpSmi9LfNngLRq7DST3oMtxdCo0XE8q9jhqSh
gTOg6BLpg1SaKGQ5FIkv36XAXPgSttdbyuRdIsDZGOmEYxoM49pJqBOJAMbe93xrsiwFJmmzFS42
eoc/SlX4aL6YtUhzoBydLAqiUeuZS2bgbHl5/Qnjf0tfBgMWNyT5Cu0QtE5scQkZ3pVWn3SrJoGd
3dHZe+a1mFxnaAnnWBZ2lS/VpOpU29UGt46C5rYioUZvn/ySq5eVZPE8sw+0IkgMQx06NuK4k7qP
+ZXlTS8G8f6+2qoseSbQ7/sPH81qPNf1zaF1KeyU4P3NqcQ8PTztK/pHaEeUzEf1bxDmYYchZGpW
lI6WAbkowDjCvxEaXkj4MfoMq6ElmsoWE3+QGoalwp2dnHnhsnMZv0yhtCJYGUyhQda91sEGEItt
U6UgmHF2G2Ql31nN68tP8xMIOMGqNfusFbnzyj8J2KgWPOQkgZU81U9m8WIOKhNSq67LbZtSY0c8
GVafOe+RPRfzhFiv40gc/AmmugcE8sr0HO6y/IGu7STEcas+y7GcP+VXn7Ow9vM6r6nsRJeHbtlc
KG4CHKN/PrOVtYenZJzGhctYR1mf7D46dc3ee6ANxiEbfO5twEdWrQmrhwB+3RchmeZfiwy61XWk
dndHcGo+4wxGF0W6DoBChqLM9NK+H5xg15r6Ui8d+kBHwNhHDCdL3DzjS1Be0nmw/4ptnZKNWV0Y
8x0i/cFFqtFVov1Axyqp8jtUqWl2VgZvqYYoNtrOmxO12DimhuGMV8uZHC9fKkYKihfHOFt94jKI
VLVn8v0RM+SDK+TKXgq6vgdfcqkNiIPzOtIukO54TFhYEyeWK/0BmkxYN565YZZMhBhFxcfYumZM
F3wNN9rjstikVhchqSK8RmXjuQA0I1Dkve9rO4Is3iFedFHKb8xjPgwuPDo/TwclhUYCD9q+9N1B
Qe9vTlhOqCb30Y0nJ2lgM7T46zqgFSBkEhRawqExOeXKv1X0NmhG/vNeyApP+JC3bNWroy5CFbm5
4DDzfBs3S5VOw1nHLf3neSN6SSvYtcxhP7mMhaBSk48C1taICTWH1wyH+0xeZlKIxX3D/DfQxKfB
Nz7jD/KCaMPykwbVmvn4yEKOFn1of0M+EL0bAuhLOjV4aWBsj5WT6r5Sy0Puns/9bd0vIWDJMtSs
cTaUjXWhSIl1OOh+JNQTYX5ERGU/jZDgRrXI27Uq9kfIn9+rpXHgz5//DIjBxL0hyJprLaPU/2sq
G0P4Lh18/1J6K4VIE3PcMIEHJSdrr533mS+ndQ/3yOyo0HxY/Q5OqMlQJVjVkG6TZ5UgwzoQSp+B
a2dmH5jwrqCvUNDpauEMJ0T8fMuULfzpa17mdw4WQcMTsj+u8wpInCC8eqGbAVAC4dZ/xvgtKh7y
qnzrs5jGX+KShEO5SSMXyQ8+O6nyhM3EE/nexQoDbNFBiIkwBFt3pYf5UJSXXNQI4jSOAeWn10bh
dV6g4IEJwUEBNHSxXXtv87pV/5cavoDjLXlPwBYC+99e2T4rXsS1dTO27z1WRPBY4tsvd7jL6g3Q
of5pndVKcRaDujr2towLiiefis31OYk+JjVE5ZHDGxtKM38uTkW0c5VrrtOvuh2UNQwE9SJ2jQea
gY02tdFzJWBZiEq3o1iIuqftTAW1hQplOzMJ1C5QbvyC7v5NkDPTcYjsbtEfOLLjJk1HOvQR5rf1
i2rIhoBZ128zNHj313jx7/x5wh3b+73WsyUm5VDj2dHCPGtrZJwXBNqhP0dzXld0678EOIGCJ4h5
4QY6fEtOwRM3peu1cN+ANuTj1LQTdufErORvPky/3yO33pAVx7Qu233VhYVuRm1k5XiCAPO2zoua
LSkE1vVMUwNlZYKtzwZQgxaWmm3C7aNRhBTCbblzdfbp3NzLiYcHC/fZIjgtdsn2IrbTyQY6t8qE
K9W/z4NdHlOcfpwOFXwTKgQ1If7PtMMCaJXTdYc/RVmYvSTdjXovOPFq57U8jDMlyPSyNtDILF41
PyZ8/MVbIkHlqBOk/3unvLBZ5Q7Cx1SDxT1l8ltFfctKfl02NoNOBMTQWrgdCU/suAk+Xe381MuW
Kk9XP/fE5KONIy5NDYj9Mj2sPUEiUbiXla2+3sBwu2MRQD5O5YG6m/LIa1BT9zEqRpBvlzLI6LPe
DrHF+NIwplzAShiGx5Zcd67fe5PjY+zBFkqMkDTj04T23BwSZwERkIx+EtC5F7PmIZxWfwlpscSI
7wGfurzY1oSPJpHkPp0caUFv0CkcaPugxATtSgQ5dt2ZV0zzGeinkyoEKTA79cjFyv6W8dfn99rL
cNMrd5ln5gJVyMZd8yMXODvLc5KXzHHTcMAdc+86r8BXRBdiChdyn/y3MHQLkrh66XhizfMBPdyc
frt04BWtWOdQQ/9m53vW7hvA1WBan9CBp+cWPg3kWsE9svWo4hYnZv8uwuh5JBYctNDj2wn6xjy9
xrwWdnYKH74bnNNq3V1zZKcbGg621UEVRWf0+jjPKfMv6C7GSBboqPbLO1ePKHnxG4x1/VXySBmH
UznSVZFMkZzicnLbaZ3CuvR0VgVfXUkTyk/PFpUkrEcPIkaN/lBd+6+EuNDM7EQf4Nt+9wk+HdF6
1fR/ZWkn4IGzOMuy21C8EKzfBkqM7Hghc9hh4oW4m84a64l8iOyrmODe/idxxVSr59CyZKyoaZ/Q
KD0iam5qKx0NQ8yGaJwFh/QtamjMROU5VDsoK8aG6Y4A3DmWAzQ5gmjoffUOD7GEq3F/s5ODhaCK
bLYkMR0Ly+1Tyn85l7t4zusQMqDXlW0ZWbplNyI8L//f7OrCN0RPDHSRmmitB7HyhybIO1LF2W5b
x3uCQV4XSvJpofZ2TCFIfOJuw6lkK418HH1/E/JLWqrKQW/uFQFA4e1QzIYTHX3Jg9q0r8zKfrBm
ngsFTfZDmmB65Emli9hxv9tohl6gMPeFBoik8eJcBNnr1vUHW7K/94fMSVWHn6wFfGRs+k1xt+Pb
Npt3Ad8JwGg3nTlt3NI/4NNdwCq0W+3IEyw1q9T4NEMbkdUQpQJvSDs2ts0OysF5D0AWcMgb2llP
p8elpNaf9gni4Xwo3l/WNR+MYVilZZ2PP24t2yqnaelaxEJeS0sCLnvBPi8egmD+N3Uo4VcNo+WX
ecyqWY4CJl/gX/TGBBt6VyUNgqXO/ZBwdMJbAXKzjzYcUyoKgApOsNBC04rJLnTDBsYGc1cNI3Cc
SDIIPAZcF/KB2tiKxzWoiti3BrzajjZZ9XjYim4hFKAbIZDttxUSUMQNkfjVwlqW2r5oS1FyzRdM
dW1QtngC3ewRddv/7Z1128YysvhuUuFZ24XCCN08pzLXqa0eSuplTuiRSjkA+8YtsZ+0n8OtAJI2
NGBXEPLQxs4Lx92x5CExZVNMz9aU1eC+4bO7UCFJmd4Ohk69qoKztqhU8ADsjX8m6CBqFeVim0ra
FnPOCFWW5cF96H4vcbeG3azICHaI1jV6D0py/SeCBEQ17bHR7DnFzW9eRRW1ufmj8AdXUDOssnrc
GyCkvd9yPXglczU0rUPUaEqNbMAbiZrHxoZhC+gH+kSyKyELZHg4cwQiC+kZPYuJJCrMVVuX76ST
x/jBE2XO1i+nFrv/xTKClZJIFP9hJA44sC3Amn+GsfCOHzSTJ1YqvMJ+8kWhJAPGf1I7ck1wXMq4
X/Tqrm5k7HnL5Hy/4Fb8CZaEGPb0xNT0G1Hf3JGm347ds+dPNaBByaSO4XC/mnInOQ3nTauNFjFR
CllsfAyM5k+NqX2R4RfZaNvxAQMzoPaMsc3kSMwXce7PC6y8hxvZLHtCRL0UKl7M09uTLBY1l8DJ
nYjtYtE8+Y2UvX8P9XFbgI13xBMzMOJQySNh2ynJVc9dFOIyLewq5bq4IwMJL483PMBHsQ6GgO6q
BYTNWIxEpEpSNfiRlcR2n0OXqAhp9vUTKKFHalCzcvEFDVMig7xysaI0OcDaAJF2nmZOQWu+II3f
StYdZ0HDnAEpO1QiSgqaWs6eFPF0pUOGpfHT/kf0DMpLv7VXJ+HX0saXar7NCFZQIFKmDJEEJMOL
QHyQ7ecWlxhcbi3dmQlfyv82MxOJHJRQUSd39V8olid0cEIjnLj3NS7g5zUEK2crP+9F1aGacfTH
uHuUuWd6h05fS+Bl1Krw/WNN5uDjaDEs5kv9h78EkhqFvD1Dot+JD6msXzQSugOL8nLcHJJZdcjm
ENy+i0blO21qofitD7LIfX5LDY1g6FbLVDlv/7sb2tQ1Wzp1Uro0sL4znZsbNDCiEAs/so/AW4xS
2glPRE4jr7Mq8aVQmc4OgQ/rqRKIZHGHVUiaUFa8mrUY0lwGopIWZ8ufTPlD+9tcNikF8NhyarPc
T4f6u2gRZA8fuur4kaIZqf+O5FRSqWbjuaD1uTu6rLcEIw87uo+snDzCgxzsOIWcjDH8Jg/a7LK7
zHMe85emRYoQ+mp0lzQlnIocLbqvRvrrBXAYy6rPLMyYxam/QXUcWEuZnTrZBAfJ5Dyz+aktyrTk
C4qDg8IxWUdoIetNHEtyKS8gxBxKM5BmVURPT1Uu1caySroKWTpaB6V2AHdw4bfTIYO1NNr8w2iN
GVuOuaVwSMNvkBQcMa01DuyeUhuwW4lQToNO7cTrQ9nRQ4RH2kkDBwWYxyZw0QDbpfVeXudumDEr
mVJlquygkLok4BfNB9NWtdWLFl9xvDbLkVO0jomdZ3sVD06qt43aG/6BTnGZDJDxx/p+ZRefJT+D
FTnG3NkDR+7gjoqAGnKGATZiMUV/Jhl9QPm1PD4quPaMxGdNtYPiNRYvdZ/XHaIVuD6uf05gb/ou
igDYbGnt3UUujI4su982ayHbtah2NQdpnqeQZ29MvVPHflH5ut6fG61lULR+XRm8RB8W6lhiI8gA
I9FsjJu1kXgOkltSxyPynM7Iek4WpDUG+/wgWHnNO2yOeEnv2Am9d6SvhZ/Ymv8qk38FbfAaF7ZU
j4pPGSH5GAD8w9CEGBkFhWpzOdSMMo6niY684/LKx/+befOHC8I9DmGHWpJ0jxt9sLPJucJpHswm
gozx5H7adhmjjU0lx2/3S4bmvY25FYUeryHW7+r8tNoe3zgai2Nuk+1AfO9G1ov3TqJBrZIWnQwn
nUS/klmfLq5elVWtb/7Y5PyJ5A/8UnOef+fQ75dkE6j5MfuC4w+ubUB6+w8yFlpKST1RSsYTuys5
BLWSFNX94BeCfhIL++Rsopi2j6K4tXdqmWWUvC2IZ6IvQqLDLnCOj/nNKDspcRkykqi/dA9lF0ZM
0jkDMN5d8RURFIJsdNND3t58ryEJI6STNqhPuBaAFOqGxJZ+rafJTXRtAyxvsCWoSuXrn9CGSHVv
BF63/4ZG4xR1J0aYGDsvIoFJSUO0G/y/DNzwJ622bh2tiQSs3AdYMXhS/p0TLPQFodKK7LVX2rxp
cL8LrbDCVPTuuLTDIlhBcaPMz4fPuiCc4d+vwb9rdQ4sGJqic2ohrg3OT2wJ+73IetOLsM+85S1+
+xfActMHSf02pYzUKrwLJTOBE74jI8L2fBeEzz5zvcGCHEQIsxZypGDiUjmNcSwafhcgOzZa9m7q
kdU2wuuyrzC9BaafS0XLSIyxE6O/+yS9af+K2XVLrr+HfytYTRTsg7dkm6UuzmuT61BbH9OxEi7D
Sn1H2toJ8A8jzO6uz61SOGl/Aq24/ItLmEqDEE0X0WH7Zl3qWlZ5MBep95TOwwzGTNuZvMeUYvNh
HW/Y4R89c3PmozuG7v9zZvhsM2x+h1HgN2cDAShmrE0gYpv3baBrMd4VMKXC8jjEeZ/FvYcQ0dtU
SNUnM93+ZXobbo+WPBwwm1PY6oQBc1qysghqIMk7EqkJhjrxeCzLNaiy6aGAeuDUA9nu3hKp8DOO
qEypk1VOCsGMCJ6vq2kP/nPJASfdd2eqbU29cz3TiEu8h47ynUd22AM7EfdQZzkBXu3/5TpPB2N4
8Uc6/C0c2VfpKWWRmttWy1rtkiV3/WIjOtbCUJJKR3kQ4kRFVJxgL5oykt3E+v9DB/ZOSB1NUfEG
C3oMPpjpdA2FZ3RsLBKpdMVIEHV8VChXEYiXuOCWugwIykbMqJUbaxRFWJ6Lvx4vePu8RDMRk+fw
mNYX+1C2JoQENBPM+61OQxbJuEoNB9CKXFryDZe8g1fMqPQ+lIo184pQ8xIwLt+d4LzPAHB0QzG+
iWSTM6jYzbWB7BIGAW+kOWAuiC/PiMmFIsR5TAiiI8qFxtyIcW8U2Yn7ytl9qSJhUmHuX64bw5OO
Y7a6D33SfsKlzx6DmMyQ81MPlmCqsdAfr12NrDktu60nb1zms/X75jdGud32goV7TYmJ7Wxul5/v
8b8cgh38CGpRCtAYFOwt1XfiYeRlJ0NzDktOS7DKe2F/B1PFHHJj+ELAlO0+nimSHwMl2lQVH3ya
whIKJmLqSr4j+U3BuiDCaM+mDiWEL/FceDElCe9SNnmWfXI883xkq7zidBQwm2r0Y7+l7JJXSNWJ
YPasYt2JYpEiIufTmUgjuEL7Lg1fzZ3Wa2ccfh6uFlOomPLtq74IPuVQ24VZwV8f/pfhNpKGjm+l
IhQKT9JrGfdQz8fB8uxLxCH9CceOC+nhgjIsdv/H0THAe/EEMtOxtsfaVVVy5y9dklC+iBfD6nr6
9GBikw5DjaoYW9WaN4OAVKLtJD5cBHQzBwlKy8r3AnLM8TeMN/wd7/AvNEMZZD6ZPDpqaBKKan19
UZWTvN9eioipyMBN8BsJT7pK1+4nZOyXeUcWrMBmZ/2pOVJf5JslzeKlvwSdVnrHDBGSbXcQ/UAQ
CseAag/Hkw8Tj3arUQuPH0OL6W/BlMQQzlzkgCKkhLE2G+1lN0PnkygoDZHgXKFz8qZMHCg3rzqa
5WnbVT/GQrXchQodopUkX319h+KYGS9epieBYP9ag0aeygEcA/Yb38A34SYXVVMON74ZND6E8TQu
h5a0ORKos7soVS2bRZZVnBaseM2+lrBdi9dpMWaBGyfa+wmTtH14jMwes9o0o64o/Lx3yLEinPnI
oYekUU1nc4Zj4vx/QcKmZSZBCAAkggcc84DcqA1qI5fA0xLD0XJz94P635Vb1SQdqjY+xggicJ5m
Fr7eRVYAGqCRHZd/psxsdVloB0LkgG/nX7knmPJYxsR8xLlvLroMjtg5XbP1uUVc4pxyNO1WZbgW
1WPaSsBuxzHmW37dHJnwO/P89lhPLYzDSpfBuyEQPgK2yI3dFXChXV7is5gbDooXANUzxIhVdqoX
jYuMcZrV4h/59QOCjlF/OoQx+pO8gd567YkkgcOjd7TjEw246J8D3ICLpOHyzlJP13wCtoP6LfTK
yRehefCttpq+7N01nMsUhKV8kIa2jkVPy11fHfIq9nv3jwIygh4QzVQ1a1+INjPAN1FmaO3Juv3a
5oKz1UepkEledre8Ll9DVEu9dObrGB88fAGEJT2B2OnQ54PmL31/i5PGze7FrXyI7R4brcRTlojH
H4totWKii4DuvJoKyA2nu6hk71ZrGs7pRnVenmwUOIe42Nh8bDpr9AoUuCuFtodKJuC/in+btnMm
2N/Y5N9+hw2tHDPfmKZOJ8uIoNMWOoH/7OGshgyorHH5BQ4sZj9yFUsrgGtRphhsrvno3vy2a1vp
y5wDizEqiNina+eiOwpvLiuJ44gXB5iBMoVovvY907GlTeYrFFjVASdiPZT836dNDnpiHPFVIN+S
vOK51u1j6Wojycgjgj6BKMJShdmOY/Pnzwz+vU2xIcmGVvk5j4o/9Wg92aHSJ2XLZccA99cwhyRM
P2aCFVgjTQ5aHmRs+q26Irb8Y5sCA5UxF/2rR1SdSC8pRo6fOQSmzkX1OR0Ha/iyYolQAeeA/V5Q
M8ZEWH9RT1D9XS+pp+h9grZDmpCXVd2RgmJ4Ke9L0H8et8OXfywmH/bzkV814Zseq+LTyOhHVeaQ
APOH945UfQhpa6hoBn6MdqgdTEH4eCt9gqudrXQrKrTuvRNNzGoOlybEwbUfgpb3Px6reUKhhM9T
1Dy/4DJbDTy44eZ+/AmCJbKvLU2Cgg1CcTLjcVFBrHi3sbUAIn7y0XV/J2A7tAq7GD9Wl6OhDtNX
R9EU1pcSuMJIe7BtJ6ze4Lk02eQyPLA0vG1qmkw0R7FgHrDyIJe6VMmfXWf8EuKETDqiqAeqXo/j
09DFXntzkiAi3oqhgKquBuq8Nge/YpfNW5PaGHXnwnDLWeF3APGkdC52Ui8pIJ+YKKy3CuzF2LOX
QUMCvucRac7UK7Hnbu82bSKDHc8MMrFbu2/M2G4KlK4qCqkeFAFl5UMvSW3PZT/STOkuAGY/uIUL
9fzBJ6pPGAvay7/L1fS4HA7badO+Og15WEhNawnphfhZn1YAqsi3dvwJ+c+ndE4G7Ysz0bn6wA/e
ABNow4aciESF7Or7CbX41fdyomFhSQP1XSYA3UYOep/PClmLoqUhjfnOZ2VeRYfzL28oLsWjIakL
bs5dY18/6cUHyOKoswbMt1K0Bp46IeG0hY2AG5NgO+bQwJSabHkswGsVpp6+nE7OgEeg1dsqSEQn
Ly5+GuI6MKhXZjmtHxDzOECbz/zuEJXqvSkeKUwuyK1+6S+vFMSSQOobHJzyQS6/iG0Ykc155M4/
/W6KT1RhPvxt/YH7SxgJriBAx+5PagUYkiSuu1MGbcGKc3i2ht8KqBMetsC+rhrV1ZiykknK009K
Zp9BArl4U51xt1P0q8blvjN0/3/xkMzAaTO2+U4ECFkU/Vg/+YQBRE594U8zpyoGXVa5KOK08q/T
Y3seu628aJTpF5BtllQEy7np4MfGaDDT8e9NlyQfmJec0b8q0vni+cLLrKnGmkBKtXWGn8HBwCbi
lSs8p0cO/DJbmjhtCG1SpK+wvQnWSuTWMItbEcaDry3kLFvYVCO+r2EdrNX8NzYOMTUmLOvvYpBO
rt4BXTNoWs1P2vuQ91sN5Uct9ySGhnKPfHfAI6GHM5Xk4JsGZC82CBPKYT7MovGA8r0BqsLBFK+p
V9NKZrRVqJoSVb3n29UgnM2JEaiJYoHWFaL8j5VCNd3B7xlV6x5C+cl3sTktk50qlMtcylTeGxo4
Fnd0unj4bHGGJUsvGo3gy2OQ4LlQXAh2nyLVOW7YOX9G9ie7MBrR8duD516MWg6U9FsZQ9iN1uGT
msaboIzllrsxMFnbzeiEvMKnzoPbtntyp8ZqC6vO0cVLiZz9GrtQDGZIuyNH3IcOPsQXk7xpJx0l
1N5wpjxTBkVf4gF/p0n4G5D2YFNfQvdnTC8cujjl00+52ikG6FOh+KvJHffZQIgp1/Vn7M3Inybm
8gvpMfi4ikn+YFQ/G+qf7lWxguuTky6YjTm+ZpbR7S0bClD4eUun8k1zm458rnomDxKCwld8aGDQ
ieGiHQy3opN7YvUDPrtDYuc31cfwKLnAVEGKCUZmo9Kml2AuDyVcjTSsnVD252NpXax1WMiKH6pD
GGoXMsMmxX+PIEhAYpczlZxXpEBcP0sZj8pN9ujCCVpKDHtTz9sLlIJqbwNqA+h1ckvRwl/IwcyP
pSvP8fWgU7Nz5DzvqzpJER//XMUJP2jbcSzv9I6BoV0Ki3oUFIRdaiDL7I/4asGwTY0X7bGvWB+I
clvi2VC4B3q54eON4AgQL8uDGUc0N/hiO2fiukCJjtqBTf2MKhHdQqVHCHGNhZhXzNQMdb5O51x5
nps1pp/KgB/zpUu8LzJZ7B/Slf2tpkulIPjER5k6RHwH3uopIntE/NbsmG7BPtxmC2xEKu8Deoyu
vh+Zn1CnN3QwLpp70YWY7gCzA3jPfXI40TZmSCIjPbWI4FSaS5VVn25WF52VYNWrzjhc7QYTPG/8
cnJwzEfQ0WpszSljGMuB2tLXI/ex/q0Pbo/AeZIpCh8/lo+zCR0Id4XOQtU3mg4JUqruHc44i/jP
tW1m9nw9MHqkVnezn+KamkJcisi36fRbF7dbIEy16dkNNPIo3XfMvpDfGID13DDTKQl4X8zFuav2
zkCJMqZhjg1V72CMsQHzcEK1fcyv909srUVsxPjy0HDzd9/sPscBTrXlLcez35tU6JimGysu81s1
Ho5uET4/omNRNLuN6pL4avLbLA5bNUXZom0sFqk41YTUwaGSNEZXiU04eQjEqil2kQVG9KxvF55M
11vHCxLfPHcWLWjKLYvvlFNqGs2AsQAgg+7c9BvJYBPhTZ7Qa9i3MpXwvwj0YiKTNu0UHmS3unUk
fTw1sNtix7uYZJxarMqTC5a+a9s4ky9tM6L/W6hh2XW+UpljloCAGIY/nvvW76KCG6r5LG6dvX5p
QCiCuz2m3ofBfVXdKdcBR7zH2dVLRkfB/0ztDzmQJUZUXjLDtMvbVd70BHBpSN30nhg3uX6qMMuB
ehAtEmBPP4QZH7Ol0C5cwR+Evtb0lwXJMUrYHX7fhc4sihi39ElGr/kS28aFfbGFp4AbwIjIq/DZ
L9BAR19fzS7GKub3UYtir274XTO0FH1j28PbIdkjenC7XJEcohoST+GmiyAOX6oJPXuyEIWk4C4k
kbZ1LdsgnSjYBQvRiA6OnfR2yz3a8Mn9Ir+l9KaQEU2ZAlraDnPywDtl0zy2vLb9qund3aL+UsZ+
cDGOtyKwqjgU68V+acNMqHF4eCIVGlLhJYiLIniBu3ad8S34KfyES1mHH9ed+xZw7Pjh6SF4LC+Y
TRJGW+eZPSYd9PBrXBtb+e2PTT8yd0ME4DH89CKvmJf99yBXvBnmeNT7VioNsM5x4bKYIDMcVDhd
SBi7NVklrwpPouyBvslLj/VpgWsmM/6FtiUV71fZ9I0IEIBC3BxXRmFplpM6UT9KY2uu4YP+jDJl
F09N3r34q3I50WQPwsh+DsYJWJgrav8Tio5SzzY47aIjMtTemZsNmTHoX1R1Rv6FXsbFPCiyO/+S
usxykzFdYZu7HQZaVl2BVqO6P2Pa2BU/YNZQAkhR+jGsrZWMIuADlXxGx8W3U4bDaNuiDDRtnlht
rj4l4IcpqMBAcLAi4sWC//OU53Rh8+m6ycZQelJ7S6AOxpBiaSZahoWaYMvvdc2WrmUuEzcgIDYx
C6qAaDtc9rWyj0d1Mi0DffOcZaxbm5SiFRSsokd50uO8QV1p0rji97pcd1MmfacCW6K5NIuzEd1U
LTONfMMn1jUeqhkavpIpQNGXup3N/QBJQ1BREizsY54qovpKaWUcu5JHWLXxttLxJjZKI7LBe2iP
NsY1/oYSB9C1swWj8CHIwAKfD+iVQ7Y69Yj8bpJu+9UHNiSMq5YiY0NRMy5VxVKKFZEZcaFaBG+p
j8T/Lu88ZHpDUjIVv77yYENBzm+PPDO5Qs4ATCwdeLWgfDJXVohL3nmjo4vqPadbAnr0+M0m7Osq
Ndc5qnTJ03xT3I7sC2WL1IoG9j42I756b9LR/QssnscS19bdQ4hIq++7lrduHUj+JCMgu1OKv50Q
rt9jJ3WiYh8y0Ewj9r1FuZ5phh0RYaOXvpY2eh3XVBHtKHEOViXvMEby6fJWd3k0RM1AQUOyx9la
uYe8flpDqixvTwFqhvLByo57kcDP8KFJOVSW9FshtFDDSwHT/eeQqWJUn12d28YPw8F0k8sN+D3X
TNyAp8tv3UX/Y3MROBJ/EJZv4ec3Hv79ABHQvYZVZErgorCsQcTvMrbn4FnjvVLeWkvchd4PG2kc
cYMtYPO1y3s1HhnGxkuY+KOyUJTPcVt92YQHbwU5kKbC8RhgKe7NEFPtnuSen/YlEey6STW7N55u
o+u+58a7b5H13byp+DmXmU/G2Q0/+nwH8X6sQhBL6OzbEDFkW27xLlqbvCzHCchYQ2TwbAxBgz5A
w7xCQ8irhD5MNm8TWcaq0fUvONG+P0wQXrnmeTvtkDbDDxRVab6SbJ5TGtc28tr1T3WaUO7tsOf0
YblEXshxIecoIxnKfrRl7GtkPpYXHFNy0WXQ3CMTfl5A42rdqWc5nQC+u1uQiLh2d8zBLatd6bOR
x+fMVRS/X8YGFJWd4XlbhA0/YnYHm+F3eytypflQ0vKYDxg5gYN9xwE7H+Cp1W5BacsfvJAwOCSP
VGmcQJfFK1SaSTIcIM/Jed3zMJGsIfPgkEf3DdFhQQMmOd7d4gEGvSEGca28ufm+/nCFT2xCJ0go
m9Zuk9c8hc6JZuDVmf9vUv5xa4ayCx2FS/J+pqtquwoa4ureXEycBzQxt4oHqN3nZbhk3CHGY5Ha
K+BdrfmRMorBJIdieWuz7qmyxHRRW4WBwT5Qms8KcRiF7DCiOtcdlgqifY+5pzn/XsuX87hPjdxY
J2kRAinp6JeiIOZTiTqVsfkjVXiUC2fPX9EMOaN6Zj4fH/wkxlWmG2jwdVx/QkOQaIxsq6DZ4WEO
j8+JiqjC/+BdmV1LzpQVuLR47pP5marvP02T29cZtlau6YRiVvGFuLzwaY84q8Q3rloJrlPEo3Op
NJ0ksAT+Gr6XCB+FdUE/kOEI7oJsmpjwhgDSo/9t2RQ5flBeFy2YzqOlyz0CmqRlJThWg8AcLJHm
CP6IK2TpnO8LrY94k0GNrFCu3SxMzWsRuTY4hx8kwcw5LCLJVFAPedbntbbhVdWvlq2Ww8rKHiSJ
MqyBQAsZ/Uf9dXkyEKsbB7SSxut8mzm27hTDEJrn2+fVuaOwbt75d0D/YKWNfIYSeIFvDj6k6CIO
VvEc6aN8qlf2xEHz1uHlszkrL2Yx8MzfU5j2Vp31IlazXMR7jTKvGdktYxTpNnioa9nTxV/3mTk2
mjJIHK7DdfaNU1k6bVmKmgeuIsdq4UtBHjzoKXyudp5PWKIXD68gruSuQ2ruQXLl6HPqPSHlKbv0
/NX8zOL5CFkkdEogOhyEswWGYvef66kzI16xBNMU/tyQ5D+E86giCNHFT4t+uJJBH+VPgvHAg5Ad
l9RiimnscpsfcuY9Wtp8QJxAGs1YjfGNDAVbA+fjH0rYtNlDYICR6YfBxly9vskfMnwRE2As6UhJ
UEbop/zZYTPFhQjhVkl2RSbuaAZZRGGydrlEbqbIL58bktZLaazQD0BmFhVCJV0j3Fljqm+UERBg
eNRggisebR9p3saULwAn6vDUxXzFsJsccOir0WMfOOjMJWtjc2mqAtvfj9+euVMT6h3TRY1Dte9s
FtQrwQgWAByAfIK7Ptt6OiyAaiWnffgiF3SSC+ZaYIvLYTF9cW2YbTzVwmNTC+e2PtOibwru7MQE
gHFZVmJa3d0VUPMjZ5XtxhnlkxT2C/oIoIai2bZT4NjEpAb2JUdljIy8S+Kf9ayav4SP6e8ausmB
ZZ6wP0ADY5hmZHGRXO672zVWrY9sF6nrN9uEajBQOAbNbYajYXRVMOqNVCbxDdogJrlLlqwm0YRc
ddJiy8dXKrpBQm+Qyos2lwG+XlRWPjO6szstA/Gu8pTkqp+bsjD7bEExOGD9jTElv/zIY+ArxV6o
ndy9NbOBAHAB6sAOpGwvyXNzyawVEkkV7R86eSKZLMyzVSYdp/RxxO38RGFKUab7NuczcB8lT7Eg
VuVyb7UKAQh9qgApR1moCqfTZO5wnXMUEAmC/OZmUdBHf0WzZZwxd3hur2sB8FdbrJsct4ol2caC
GApJPRGAgtd+wEUy97vpyXCYREUST2g/TpYvCJeEsdY2MZvslCfsvVe7Phb8HjIGFQ22WWBEmUDs
KEytX1eECdJUyjjdxTU7Q2bUoQyphrAdpKjXqu5HtNL5WDY1/UzkmSslpjf9XgsdLoJXQU/WxVr8
0IfhQxA9xr0Zxqa2bQLrLZSqBkjFUug5nDawhVFrWL7ulcruWGhdmr+CAbStLPQuhtv+nrRpKyCy
iRquDjYnaO09D/3DLC2dXoKmWRN8ilbcR2usMiIpCSZOT5UjeH9tP7pokO68Z/fUJYtb7M4P1Z0S
fP3S9nugDPBYNoJFYTbAj+r4FlZv2z+Cq8M7BYXu7uyeYAUEDoOGstXYOrOUEr35V/umQZerDFs7
pE0FJuVkiLDAhL5PgDAt6jtfrLvAHfom2l4eDetQCpPQophqgU1iKndFicdurGK5gvxb67YDy700
25g+AX9jJIq371MrP0AERv0okxdy0iVNZvJqVk/gxjt7U9bHHWzHaLFAQY5s/Fmnsm+DNzHzExtp
WFbUvjKO6QwgcX9D/KJmo/cc+fe4HvQeVxWcK16wcKNwNN85oS43jN2VNLUnN/6YoB06UHpMnc7H
FKAXecAp7lH0Frn4wa3Mj37azgbkGyFFVbW6Tgs7O+V01ItzYCgsUZQyCoKexxNnqTR2/VkgdYMC
nzxxq8doqxaW8VzE6A6XzpZ87B/9PU4PtU8/tj0Zthbm3mCQXwnRq8qW4BSn4RNSYSxji0WjOsLA
rF9fwkv6CBIQXL+hOPcrIKEiQoQanEfn3qSW1p8bSgg1pFH2XFFMq4nlR4TKspmM/TYs8/wDsnQf
c+1nMLuvYI/qBqzeQ02eQs/yv1xlzUmmRYzLE0XlX0T15uy3D9jWhG9l0zvJgRQGned7NvQsshpF
+MefVNeCsgNXbg2lrjXKWjEs4W3ycNYvDuWRkP26rwBUF9lCS0yfCyjM0bzSxEWlF7cbFmtvhf61
9GTtSW0seDlZhbqPUBHpuyU9elC4LgHsqrDUxtMjHxxgybB9rl50a8tQ8vBTGJ6NH04w2KZbPU1i
+gqFMGuHKuCJEwvU7HzxxAJeaDcXvIgxUwloKdw1U+WTnVP2z9/aYCIT+TrSdaEd6cGEx3rNk0yh
GAIuBQvl+8GGFTKVxdHgG+TsK6bdnOyxJ22+L9vPBZsAGu3W75eKoeMi0AIwhel/LeVMotqHcWCq
0ovKlJHGqeUmOtI0AJkuO3pT/ROl8FDnAhaAjk2P3QPLEJE2LBaYxFiDdwl1xdmkXp1qQPWFhdZ2
ecPA8H4blnbi3p1uXb6veWRbQLPQs6nNRsNr/hqIrSD5G3ffXUoj7xSOS2X+NffvKIZD/Swx01vs
haimIVTn1xDA0VuKvI56iF1xjtYvprXU0cpIXnY63Vk0byqHcoYMoPimjMeCQR6xHHOjCFUvZPut
pdnDBUH1Z6aK5j1OH7hfTSAQvvUie6J70n4yv7GStk+oGuh7hXqK0KkcqGvveHn9BEfkNmHgHdL7
iV/U+UyUw/2QNUyZkB+R/iisAsvcPHskfopB5WxBjabUdD9xE38dO75N+zNPH1+d0neOh7IJQgdS
viAL1mCWy+xF3mw8f3g9UgMn5FSsH5CN/7IripuL277mgCFIb22BxGJBZkaXX1u4NBa1fM5hmVqV
Rj45ihEIJRwXa322KCnujdmbAIM09LGemXjXIBvoeHqlu7UeX9gRBHOOXtlvOZ6tH0jc2Njx6y+D
CIm1lKHoV3qFvS4daw1FIt4na1gi25+VESMmzlxjneJtTQNiVQ0a8b7Tqys1p8G1sytORvGCFRas
iye4X1x9Bh4q1l1wWMiA08oVu2uXgggp0OsicV2X6Dj8/yYEJExPug55CxujVHNZh5vZmjDM99KW
j9KHlFpyAgcAmWh6isPpPY9QgosEPULr7/SvF3qRF1Cwe4uQiTVWPXqLoOb6DLP/OR9fXX7Ml/D8
eFgj8eJahDCrrOvqilSpyB58y2A62HjVuttyBdDFmZapBWs0FWorF9v+S9lYq+uGPWhj52EoColu
zXZXuPMjjv+oQ7y/udkh9R7jCp8GpvZ9WiSYf80zsnvAiEe27q7nAKvJasROLu59kvFGPxI8KFCd
onaJEUYHXzIByYKIO5n1Hf1IiMR5linAHZJzp+iGH4pcfpej61toIpXs6/TftQGSamRgPeXCqEDC
OE5VoK8WMQcyLnHK07NtttnM9L7Q5zqNKoetKqOwj0v2aktAZ99hP9I9lUaY0OrMeS8GOqQc5dmf
O835d3JTLPZgj8GjYawqArh/Y+qiZ7sLJTM4XxsH6Y1JoM6Z2E6IxDp4k6gCl0rAumNXs0RGFPVA
6xYt6jUsBvpu4e8FzlNGWEE5Z6fQoNAICT3o5TkmF6H5UAD+pEe26xCIwppOiZQzY1qsrn0AuMqb
iYr0PT5v6RTmmVTPyWd3xVTTld4NFWQ4/+EHDLLaUglEsIuUMdfxF9JLd3dlYukaIAlVvDSk0jGX
n0UG8VuRqAzYdOBTCoTy+EHvgK4yja39fKxOniYyYNJNALilqQVGRSD623T2yEVTZNOTVxWnsxso
CZTn4L5fTFYHKYOt03L72ZvLCtQl/C6TJAev7mNtx1yXrmCitxa7nyFQZrlVYtVZX2QEeG8mO+gH
NFbHz5OjcyleeS6IQhwrDYIECx/oxMCZFJHEo5GAtMcwVDnzoix7YgkJtmuQnYXBWQdrFS94zWqH
vwVC9Jy0udnpmPNIFZNJzkQDchAlWoR/L51RPxwXkXQO9h6Gie0yvRy0wT2NV9X1zSdMtXKQvyEL
ZHzf7CRMxCMnK49RTUgpXEjWjPD3v0+SSODcFFs+sewap+E/MxHmx5Z58RnizTeXVgiAOT5gp8no
KChtovlL9F3ERW62imLxSATw+qSgjHRPXpKnrazxvqGoCVQWqq9F+1VceQ65TsvAbQ+SelfzJ7ql
pzdzWBfdpWphR93TjCy0LSGZals0vQEhfhZ1EzvGTNCxhrcLPYd/NOHPIZM2wTmRMpd1lGnyUckD
wFIkBu/kq55zBQbvX4RP9OCvmjZKQn0GcEuspxxQNHPrXpXf2wO3ETx6WenzZUM9vlvUA1fZA9Ey
5UhhlGTdjkprNQJze0d1uHUXH9zxnWNLBYuvCvAFgyML/5tW6CLo7JisQpI3oK3afcXNhgK8Ea4j
UZZuET5UR4mRkmyeOnAkAG98MjU2c5Wy4wt82HbkwCXeIgyYcc7BI3GOHNPORJqtzwiG7AMTLEeK
1xLe+mP9V90c7MvsleDA3RjL+jNf2jggwcCWTpQR7OrIfnP8cfLWVcOQGoW2kmsIAu4hSsS42YeR
tggYZa0yGBujqD49AuyZgcwbBsD50h2jzwQDbsiONIxlGrEBdC0AXzAkvfS7Qzp+n4cAzHj6FGKl
oN1ap9kHXEjD8Hk7zmTN/RIqeeNFn+GL0tKAdounjWpuxGaUyvZsunZfilicISkrHo/AuoL3Pnek
2vTnODMR+BU/CZUEcSvmvhsrGpWieULAlTobjERs5wdAf8sXJd3d3bMwUS2EvYHa+3PZBnUUBsan
kO+uTd//vAQDhQUKKHMZcYDszHRkTJx163q0UeSFCI5IA4dyykP6zjexN53UCJwhSzvJoSlnoIf/
XUbHJYO557mEicE5b42TSGYKYbWEEKkbeG5nR4KaGw0AJVH02n0vELAI2ezazdOGsG9IuRXCB6qk
EFrhIvhSGfg9J8zA45JenleHWi19Zq23CHzn+qjVtU2kN5v8Gky3ZASzK59eRgvnZdPNl4Ihr6HO
0AFgXJxjZzvVKYMs8DzK6f9hx2UqoNnErQjeHV1maCOnrhIw4Wv1IpidCwsVVB0JJQbi8ODL+SC1
gnqJyYpDOnmmodN97USKZJPH/nasTHbf3+KWzl0aRj9KfGFQqkd+LfGQpIRdyJkLPiI6eoPOyg1F
9Nkt51sGtsoWC6K2dnXJrNzR8nVSlvpAYO+zo5bsFnOWo8jUkQ38XQpY1Ux+h2FNfivjED59+ztc
jg+/dze+pOc7grRHWCUsamPuavQUf/lbsoVo+KBQnhe7gYl0ksLkuLpmxRmT1zCtN2QI3dxYtaw7
J0N76lZFQ1+uXZbYstfXCJLEQEJRbQluIo7adoS2ZCs2IEKV3tw1XwP0EuwE5I6MhHsVKi3c1fHE
WeJuT8uKAvoLJqwkAaNPhk7Fds3JPa0UNnEYNWRLGM4m1bvHbia2jCjGULGpH7R0Glg1VjKBOZTb
Ze+/N5sifEgfHoTyZ54XQ2MyecaEh69gXKKlc8bferzEDxgslGw6JegHrefxipuWwZRdHlAtOJDz
MQ+EjKagtYAf+9j7HR5I95jMpUbglY4rpG4FsggTpEA0hbJ1NthFejfhU2h00APfhB5I5sAhyUAl
hphvtaC69v45XM9emIQJUHOptn/fu1Hlun7rmKobqBqJ+qo7zmJI6rOPJuLLtJvlQcVvLvHcVg4N
HgrvcnBCj0fgs7KyRbBz9podHyFRk7cOLyZB0pJCx3hEAIPW6xdNXz+OhHNlh8IWb/gHgmtRxyfg
3zqdb/ButoKb1ylNjEMDtDpTeQFPVMMxMaFViW3wCu9DoiAjrqo4Z1+mCu6YefIpXNFQPBff3LU5
Hmygzh4Kw7UVLGp/jDy5L5DAWAJAtBL5wAdBQJOVFbz4YptpN353hzb1oW04kGUKYq5ZWVVOjEYc
cI08xnotSVi4w2cCtu9kodxwj2URifBdu7zRFXa71rEeGIS2oIsX47daR6CnO6x3Cdt4L2Q2nIpZ
MSHCLAu4bTczppohyHoNC2YOJ6Kx0BYs11qLT/UFArSGIAVxmaP5J4P3EXZZII1qqVP+dorMwBdw
ZgAIMiHE7ZfJW0Sx9UEQvB8SVMnO8B0SaQh8vk+zZdRfp/JmKurLcgagKNkxLlyz7dYtn3M813pM
cgP7uTJQrKGd2zyK1x+5rwVSKasaVjZN+S7tFCj94KpxtyKxOCkvmQLBPPKCyAZIyW/+xzkDJdwW
itrq3GNBY7Rj6XQmP1doNBXA1CMqxTHm/AIqpUsbIU9eHHBIy5M/viExSs8W/5qK1wDZs6IdirWE
6XZpGGp0Q5CSkstjZtTCoeQDNp7sOHUmF76JOCpnfIU4eO/5p77ZI28i9/E8ou3ZGTu7PSL5gtSj
Z/zknccdu2z6LsGqQTkZlUiWCs8r6f7T2rtWpGFGKYYI4YHiJMn4v9bami2RW25eekAcrSLngshX
xKAjroQJyofATsV8dsg1x6Wf6/U+sG8FFLYkJUGoqH3u49ZD2c2sT1JQTSgDdBX6R9Qqg9aNIpXH
ZBJlDufGsLUOFxBMSfhrWNywVrgJsGPH+hXSojmdDYy9G0lP8emeUPTBWbq02eDSjver56GWXxSg
RFq5OiCwegvUkw+rMJbnO4jcHThZBdpwo1MVenj+B90NMM5XZoCxmzSZhyD64qx7OcGWS+6xJ39i
WXMN0jBaC3IwM0mpeag/8gX5Af0GjoaPrGWP72JhbHQNFpT7SNoSLz5iL0qQq3uOu6GGsmsAFRnu
52ThBmDTFHs9IwwZe2NvM3tNOyPmX2P9UsTPn3K8T8nlNH9sPZWtBp03EcaYtXbPxwaOKkaNu62/
OnpgKupwAnmql1X8upzid8SyPkMC8ybCrVDgpC1MireAwERnIUwLR/yTjqr2Jxt9oy2XP/zq1Jw0
tNkPQNMhRqy1lnsTdwquacqxh+mVYLZNcGjXySMg2aFlY7AQ20WGMjLG7y44D+j0RmAy2Y3PEb89
u0Y10rLCsYXXcQBn80L9jESzJxTeTbnwDRuYhellvr47IgVK7AGXb6YZuFL5w11zXeuZliMLa9PA
VPIIg+eOPJU+Im95KOLSJYSWfNdtQQ+tbBJMwlTqAnrWobI/u4cY7MwZzye/mUdasqCm8qzJXhzd
QN0Pe/XHfe26yn8oRlM/5n8lpIM9AidO3VqnXMlDohFd9BwwKozVZdroERk7jSiMlt7ThkYGXIVy
uUwCM/u6SOJQWwMUqkhkUOsRFruQGuT10va1tVEJOEit7x0xJjrMM9ZU4mGeyUfyXb87VbuRvaxo
Y0gNFRbnGcu8REJuv8223AsIwopscg4wI5vBYzBwfPATfsmssAzFhlidkCb6NCYnsUfpECpB0FIB
iFB4EvnIItnerrTQwZ9sZRZlITEHk56qZ/2OTh6Yvb4cXx+cKGWOVd+iR7BhgL7wf6+RtoBSkYaT
BVXUj5YNGgwuhy96hZCWWv40rslh42Oedx5pdpVhH8VQheNDIQ09h2YD5ytxwA/Ak9SmNERTeoop
hCDrdwiO8x5to6XQzAN3Q8wOgC/J5ECmpwCHRhXZcODGE3UTApyj56qsU2krtmgGhY+v+sUwmtbe
NeFIpZexIakES+e/jxi96mZr6zh6NZXvGHsvFxGhLAP7joVDL0sLHcb7BtWhZDvdRwzujQDUqsFL
p7gyzEDCww+mfNQxGyLHgjEHhCwDpcstEm3rBVwsQuzzmDunvnOVjjYx+ezC8gDdPzDiptQ6PEvO
ulaz5apcvVLB/7C/UteWr1A5kFYnnNZ6i58Z5nR8/P1J05dTAkmnr7LXGyr5AUrqKWlyMfE/bdCf
J6dHdxmpzIhO7Np6FCBE5OLo13yBN1soLYO59juWagRMLBLCTCRU+9M7/p7I5lgHAhYoS2Qpfok+
gpuTKuHK5o5AbxG+bpfdbgh5mwfWiidawKi7DYc0N7iKkAtM+/Hxoc2VGSyr95EQAO1N0CxKps3O
SHSd5hPeOEzIKPlNL+W2CqDFSBtohalWBs3twhrXRGAB87oDv4fek5VK7NDLMWhqjXisfwXI1MOS
wN2WVFyPBKt6vC2HxRcTQbo7htK1gKnTVEdAKb4E2p+PYfFQpeljUHhNYPjrr2gfu50TFz4+3G4M
vpjFBpaS0G0zCTsNh+9dybxHtKtkLKvgB4a+OJJaxQWMpIZfa65apiPT0C9IVaIE4KP8jPjCJ7NI
u5TaJvFgEff19kSI+7BVtIgEqtFaFkF7qduS9MWUBr+yObroNtsEdtBF2u5MyE/2MNR787xHbMoB
r52a37dmbHyHKuudnEwy0jqM1pTecjmK6cS3gqQNBroUJDCMoj1lnFi0geZrawPesyOQzf1F6cpB
e3cr0/5b3gPJTVdmc1LLUzBhnVG7mYkdq4Fv9y/R9P8QkaejRiPcrajMIqHH0i0t+0vH5geFHZVh
BHpaAiAbaC7p57OrlvFRXAsANgAJkEgQW/FI1hbhFvuPqx+zpA33AP/G6vcP5U8HBQfH6TRcO1GR
9JR6ZNcF+waMujB9QB1yvrpRSdACXvZ/rL87pgr/yItPW5dDYsac4f6HSxx/B6J5C1mGB099ailS
UhYwygqnGM60Pa20gIizsg4GRElSnD2B0RoDD/f04FUTOyaUsdvRmRC9m8JgYPy+btrLh27Hv6Mp
X69af1M6RJFthlhge4VVQNrjMH7UP1xbOEMwnzbJtC45xsAmbnweEI4U6yD4wNmgPuXuCS/J8gcS
UpKYrcFcjd0rkToestZWULg55+nQlVNOe4pjYb2d2/N0U9r07X/p68AjgqFrFXTXQnR/BkjXQdAg
bgI6oq3H7b1XpF1Lrab8Cx+nUt2Ify+4f4AzlR4j42DFbJ10tVoZMpZNCMcUlmHJjMsGDP42fSxZ
JnqnMlVUPmOZuofSDk3tHCLbI87JqsNnLPdN+kOZiX50Dzceh69gJRrmfX73z8TPGfGf/PPMd5yV
jpXgBkbkpV/K6/HNd0b+Q5XeJlMxNX4aKscFKeCtMIvmGBkiA1/nVPGEQq76MxLrFqF89uef8am/
ZLFN4n6+93nMzz5S5sv/Xw8K0Z2jq6626iilxPKWqFLT7ASpolFsh+RUQ6uCs4uXexE/cRnXdLel
K299ZaJrRvFbQAnSNvyxNLe4C3pPjI00L0HmFIs35mhstp5Yqs6QhvlNQJ6J3lbyH6MYmEGK2d7s
3FP4/5KB6RQ2zw4BCnUGwAkfmjzYyUussu9x379bbOHk+RvIwHjloJp3XLwQSZQZIMF0/clyReuO
6YboToWr+C1eruI53YkqVRHfv71AjXzxrCYHJo1J3Fs1lheMJYWG+kNg5Wd459fg81kfLrstQild
v+7nRPFIWuWlLUcoU3gWPg5uHZJkta7I63kGYOxdm8+3f8xOGE4n/xv3KSYt27Z+IWgbpkfjdKct
s/3WsEa1mg/4aRXwnBNtCmfaWUYmK/1pgW6RilJ2l2bK2Go7UF0KRu6eHQy1okg3JzbKTQK1my+N
kPOjMTxQDFxAXM0vxM+Vwd2W2h2YWGX87OgQwbh7HdnqfHDZyIjoXtwspjqjaDlgRxXYyWc25Kqr
4gYeQV7B1HjoqWFPN1ZmUhjdBsY6ojUi99ZH46G9M1uggbODrDPI+qJfp+1u1V+lZyuU7M3FXlIY
agxmMdlUlfm3hW21b0kzhYnqGftpKqhKyLPG0t2UCWlgQk3ekVwdAhCXBs/H9cVneeuB9SRC9vTE
0irzxrzFAzWhlmYMUrW7vh/hNodbl0nx05woW4SSV8iMAEhEiMQbX5Dv2QwmC8Vvzk+qhSRDM8XV
Px4E4m726TLcSQGK3+QhgPPpjj2Q04Mc7H5RpTlxcUt5HUTk+pupsjCMwaaG4qOh0ZldSMoTYwAf
loRY7gulWSzu3JFPfOR6Q0BcPTkEAsKtxm28nnmUmhzcOX7RE+m/GyH714KciYwvA6s+TfDOA8Tg
Z1ScQZQ6bd/7XSKXYmxqhu10F9qkXcZCu7WnEWAdNrnRxwFf71ft7OX4BU308A0Q5k0uwvO8ommT
JwDNmlQvVPvliXalaPskpagKqtuudbeHQ1dejSop/lDcYuzoeL8ewYD1ao0N033GsQrZw6AESLhm
65ul8ITSJvUvF4Dkft0iIzOJSRB0dZJLluwtkA17X2btvpS3ypUmBrvbKHfMIyzD7qIUkloiJm6C
lGfZvq40Bsec2wRVMb/O1aIY9fKzlmNI6CnmdaCmcfILVlQrtYiAuSsgTjJyEGNZiZr4+DOVNlA7
xhbxx7zUXWWOhs6HFxL7frgoNfNyk45Pxj4fERUDEtNKfan5BAw7Z1+pPUWlOoDiXwKRCrfD7F4g
ElnvcveiRGDxfDgpWktMbIkAbAYlJ1hQYpbTY90IUhGnRJCGRiE71Vo1rDwlfusW2IgWMtLFVSQM
acgCtRsIMIPManZZtTqhP+ME8JRhk2PYa+8CsnL1yQ2xuNNUrmd6OWxa8rL5gi2/2Trm88h2GX/E
WNhr+r4hcjowm6OG/KVUsBNoqY/WvFCK1G0g74RyiR+RM5B5XUz5u46bh07iDIFX80XPmxMpJMEj
y0QX4udHqlXcp2kt5F7XvZsVj7vFE3XCTDPaRej+wBJIcPcwMb/OAhdnlRByc/dtCexRqGrhfRdv
TjuDANHmKIBJxX6J3I8gf+GWEu+cMtcrnLbUb13fSj1EE3zo1R4GDGlgu8Fr3DlRj71iaYzqzGOx
4mz3583fG4pK0gh5xbBteDn08o1gWa/ODBDsNPqig++Y8VvZ4/3sHYmdsE+j38+200TSFJkbzKmG
3lzYHNQu/TY46yFXn39TZMbUip5ebqMNwSgmXqB+AHB8C3Kg+mXqwN9IwlNcYzXqzJkwBn5wPuQG
SMKnK9hzwRnrU2YrBCqPFKMkMJhLJrc3bcetiof5wgaZIDUrrFoRlDOxry2k9X0Ik2Z57dMNZ76u
6+o23KVwOcm56/yTj9cGLuXQJON6kJbgSy0P8PCGwFZx3gvGfoK3K3KlyXt+gS6ccFP2LUiJxlIS
g2uYxRIH1YuU3EIaquUtsY5RI5Km9ZDXzjgXo05fOGwNBVJkRMVJ9BX5LZkZhoiCKMK3Z2rpDnIC
7VCekUdi3sJX/7BUlZKNzfT+D767y6noe/a6xZ9j+neT1MenIov3KXupTV8sRtH5IckljvRDYpwn
D0WCrWzwqUDYdxyUi0qwEKwpXIOQSwXftkobU0luz8tEJPeFgtj0fKJo6rnFYWCiYp5aoIyL9mVE
uLDmh1wv5HahAWSbUhqsk+dY5kOQNZ6X57mL2KGLhCDKZMUsLODXqg91/ETX65KyQ2RpHlKCnmml
JgP5WyStpvss9M/yZV1zPcwjGmgd5cPmzwwL4nXQZQEuk13E6vi13bvCAySD+Frwt0FVoHiNdUVG
as6Mx8rah04WHlE2ta3/Kwh9OdnJIZMx6B8coU+Ffww1r42yGYYVPaSY9ZENkVmAIngw7VNKy8wo
mFF6wO/43KqClILi6PINELe89BNYzW2gYP1GhmCwslNk9xpoO5bDu+fbutVt/iktmj8EEznn+dO0
1rJt5+0jtoc58FKVk+ep1XR+I1cg4FB5yCXmke0zXmHGwTAxdH6Y9vBXc6C8I3zAwzsOsP+ydDX/
tKOpc2HUq5iRUVEyDZZW7YSU4a5bF6Cc+Ss0aZzxZ9AETK2oF1fHvIHpELp2bLfvmg7ZfXgvc3xz
/eWKvG/iqI+qxN7x9JlyhPIUGRzaDKAjAQstZa9inRdr/6vA3sDFO5U9WXHm8z1Yy/D6/p4TE8YG
XfrRMclMvkeTpXWuEH89VopQAUoQSPlDmSlJ2bbu8ZEzB8zuDW9bVK/sIpOzGhaHo9WL6yq9CiJk
JNwOM9dCrrDCrDhMfCwJI77ZEg/dtgDgF9SoK2IoOk2X4DAADHRQ9Eehfn16/VdhFR+7aSa/P7zM
2R01S0r/cIrRswQDx4TPRSEsPztFKAybkGmYi2tj59qKjyfytM4Us4tD2TgWhbEZoggsTDhuTsL/
sNshqqSSxjobTnk5lBGtnDarjrggzOYHEwNyQk/E+EUC7C/dgMcT3+OSnJ+YqYm+c0WDkheE5pT6
us7D3EcfILRBVVgxecO7baJx1JdZQT8EJnC137Vz6eYYomEv9+xGE8rq5M2pSk4p1kcAGrPuxdaS
pT6WJzrYgCC8uxrDvTRS0/TGzdwjdmueaLxT8nirMA9FrAANdVNbrbT+9BkCdAGoKKlpl0U7txmh
xziDeo8O62gSbB5NUJN5cUPapvXIlV7oYdKWJkn8WkrPYdJc+sXuaoRscL/k82TKiyzXpIb5myfR
Ei8Ve1aoZ2C9rnNa5BPFBSYEUGjtIUUS0xRhn1qMYBqxlKX1QeqRXQiCZ4Qn8l8PET/p7iCbdCJf
sSokvARLipTqeSPyHIGDiBFUbsC3LXJQjZ08HEJp1Dh1c/VqfpxnKBtLPJKMNAwd+FmvoCArKPfu
AjVeYxbNb4J5CKMcPL+xGXYYq2ary2BIHNtmJtcRcLu3G8dicotWONJ/dDhDckV0Doep2wj3o79R
UZmC6YOBSJwRjxx5cLe+SNAMvobQYUDcJwao9yyGwoGF8BOaLV9Ki1XL3YH4iwpQODPhrLebFLUi
fzsD7FimzuN5LYx9RW+ES69MdceM8CJ8s8Ywg7QffY3iro74+9ZG9PUBorc/Nu9oUMz1m+xOqs1N
BiAMN8GySJiDkiHIxpL87isDmp05jWQaKj/dr+AhcDRM0IZ59EZJAydHDQA7Nxw6LQUtxqnetdhl
gJZXxuO5pdOicenLPRpGwgTt6HSTd30Ii2fW1GtX8gxMgRzwDL3skEUBPaktmxyUZ9uNZZq9mQLv
DY04t44oR4RfFGFeLPkdQww9nYKOM7OUmgdhgenwIfirevYRCDmQGq1vQ2PoFh5bLe5x8Q5mNKZj
d1YnKHxpBeJtZOjb0gMl1pisX9xWKWr34RIrDmoB2l3JTFh/78C2bgx/2mWHD6iaQTC3UwgVR+Rj
kK5BCYmMeAiUdv4ii7BnYN/iT5Dxka9XaNGCMZslIBIc7D2BK1wC8i3/f9gtE29uxtZTMFM8vVZJ
+moEUcOIIGb+qct2p8usHPN1T7vcvj6iMRa3pyEYuW7tYMYj5tiVhB0xdOQvXDuhGe7GDw6izq52
WQVeLCzSCkhVpu2l/GgpR+FvnRTIUVIxfFB9I/Bv0hJ9v9fnB+kr0bBDai8TMXXTmbVJsTZFPE9I
mC5iSZYatQ4wqjDFDmVr5wyAFjp8r4jK2Y8gPeTrXICl2DddXLD+Y6CG2fjEZQYE2Nrmc+BAOh7q
11SpRoP/omCWp8PsJoNcyi0qXuJgznuDwMHabKeSaEo7AyJXnUIKJ4Mtg7VCMy3ATXy+U/JU/Nds
imRwSV194YRxNYef/d4QzpbfNIFk1vewKMN8BE4RfBhgM7glgv/P1UwrHvBsYv7oIkWjbOd7Juqb
bG8Zmv8/j2quPSUKxBjgzTjvq5+/vk+FHTmJR5aHKWQpNy2T9pDu1LpWAAKFUDjZvP32tstZMNnB
ikpEdu5TC3Vyc0k5aKcBztSWADkr1X6H1hlimWPQbKWgjA9dMxWLWNsB2UguOmTUrAN6RKS0MBMZ
4nUGZ+WyW+TmZY1DOfFZlWXhQp5W1c6xfcwaAl6t3XrBckGfSB6ha3tfsJD7cBkoQE0W7WEPor48
02hp4roSNXGsSzlT8yAHCK1gx9Syww1Vzwgisbfwo5MGGcq3wLfWovP1llILTbKbqQm8doiAJ0+F
TsaF1sF3+16f0n9SCFQGPPktM/kdeoo4s7qendk/0df7CejBVRQdyunM2927c/QT1QlW3nU9weEi
10LiB2SybpQZLgAVYhObRHlXsW9ydwvs099IFdAZtWTci/TJptikk5FKIMamoZuuXtqttlXD9RlD
D+/rdGIYst0ry0F/fS6JjiRlNqGTXghDJlVg5vvBweekUn38YaWnbTn9YcW7081eKnVK0idizWAb
BJ98QKXaP1ozTBepyoopTfgaRVbPC44llLooDQR7QwBHg4dkzr2KmpBkRAn1e/v8Fhh6eoGuBUpk
q22eGg0vUywaow/EKqxMbbkeJzSMc1Ag+2dXkNq9mWUXFzxo9+77VXohfp/OXb7laRLJMy4p6l4G
88mcV6YyxGNQhPG93bf7J+OjUZbhaqHZoiKHEXWSqSL6Tl7oi94mBMj3W6wTEuoMnFSBeAX6uz70
zh74OJqQa2lk8ncq6tej7lV9CmUpJVK9jnvSmgDOdtnzl4o8nTCITrNl7frsZIprbr0ez0/c7+Lp
lNhJyL+sIk2Ojjm9zawIEWBDzUjvoW0c773aawUZ1IvAYknVXrvQ1kmDMHrI/EzaBOfeReJy4GGE
1dmeQvVj6eIi08OgVHMZz5FvLfCn+IwQqryyy3KX6JZ2IABA6g6EUI6BnZYTPjSuRcmddpfFIjg5
iAZiZYBhsJO9nvZyGFjg0FlFBEF8Z5VTKVSGBgQmlTU/MYBcpTwVzajW8hs3L/6ggoXnay7xxT9w
xu8VS4kUCd+xFLo0XxK+ixvtb6Nhk+eKss8l+dSopt81pP1rWrOd762vYVaXADZDbzNsRrqFthS0
l7zVQ2jxTJavL48tjM3h60zoksdmbpmjHILItTFNcVj/tO6jxN0z0nWSCr579X4JykM6T2Bq92D4
IR6EsBGRqv0KPCiT9sXrydBw5G4u4N7/n8LL+W+GwUVZSeT9pJaGwLTT9F+9x9NxydHR2au+E9xn
Zykqy78cG3bheMzUjAHKP/YQ7+0xZPBLzqewfk6iEM5wvu50XMLml+DJwt0zXVdxrdCozfxhEgax
l5X9OAYcvMooKVsvdaBmvfxwEjepjlGsjraV8/AraN+y2iO5HwzZJa9oBvnM9Ic0lyicMXyYb1wC
X7ie3OmuqNyE8J5ym7hYdJxQ2V002J5mdbZCXx76acNNiYiWRIqAE45GQUkXCf3OeJoCp1kSJ65G
HCZ8fiQ6FMeIuiBXLkMb1fPvW218Apjqyj869VsCpeUodtjxT48FqmIQRLdXclWtuwl4PdpB4+QA
j7df8eGXvWfOqZ52iX9oPVIuh8Tb/tBm+tDItP0kgNGG/G4LmANv96GXe1OTtaRfQsONkiVycGJ1
jt0DjMoDdd2Nm+La2kP4gWHeNy1YjfldXwSepxFB1EDFbFB+W+FX0jt0VYTccNV8XQ0RUiHOIfOR
75ErDqerdnO8ntsvg6iZWNA501w1Ih1KV69dr8bD9K/Z2sSOX1MHIDL4gKojcPoeMfTJ+I5pjtdQ
0UztyN7lWPnHycRQ9PXqwgRO1bem6VP//vSqf9O44De7Vsp+i1vniNwtgNi7c92h1pe+Rj1/NjYx
680ATCzaSTgsCXQKW+kmJ7c8aWAtVhYysR2n5Rhe/TcppNV0iyfTZTNyJ1IsCfpFK185mR+xRVhp
RPm3HAEjLt6/ffQiQzfGGCev1xiT9pvj42FgKIKcmEhDAGcxoO70G3mLS0+NfweQfSDogDXyWWBE
nijSsABH8h4CemHVCVSmfdNNbeNskZEValgwZlinnHOI6sXvCS9255k5Qjlyd+fk0mhC7D8+5r5J
K0qjuWb3s1x81D/GCkexL132ejh6NmbhIRkhFvtYKceSrXreYFGhw7QUy+dbNNQwsO4FSEsKxybM
aI01POB0d3B6btZ+ehrPzxr+9qXAQdAhMZ40XTxiFIrovEUCPWy39mh4HyOUJw7bDe7YsnZ8Ol+3
QpI1z8KClP/9IqG8zIO7+De8qhlBBBrFIPVzs4HiHar5GqatXx2RqSonrSy8i0+XMYNWy16UFcr2
FiqXXJ4ozWDugsH9kwijoGK7XT23zLWkDS554vwa2X3wyWBcAuS/RHqI99nLIj4Q+ShQg1LFlUzU
tzsyyll3/mNuSTooHo2ifYiqEuupmoGiLhnILXrPXKsuz9FFiRp5Sr8tzRZCAzF9tbBLZZkb6nxV
5LEOEUk5c9vKpITptV41XTZycSWEzQpo6I8TboAU4bn+Fpn1WSYb3awrJa8/JWETbi+EBL7DZauG
YuhLwQf1D9GKsQz63nbXBLJbjQum28Om/WS7VNZ24IPi6ZapvOzTHr7GuauwXiEs0ljHIiiLofbE
YuHo9DXuKmuAwAFEk54rUDbTgqG3FseKELe5c9C7dtS0zos1ivuRlhGu4KftoLsfPmBcL1Qz4gsx
oHALfbIVJ7xSgZkpuP05aOK80sfCFLYAx8hhvu06EtljLn44S3qr7+XHhMzXKNQPESjBLKkeSzfD
kwKJnmE+zH6S4BIt2s2jZm/4QrzGFUltNMZSqw5xJ3GkvhAGHPgwM5tLm8eGwPhQeD95F2m/KEyE
ZsPP5ATM3YQzQ577C9VNwukMGncMA502MxavuDoCmmYimDql/hc7eYeVr/fwlNBU2LyfJK57qvb+
DtBMSRRyiZicDJXgjb2tCoxGZAj+S+IwGf6s/zoj87+BStpFGPIbKLEar2Pagdy7RHH8m5c8o+Vc
k3GZwRjTVQVLrY6lbd9F/UabV8IF3bdukAD2YJD7H9bXtyTZUxJU6F5BZ8rmRvEHgYNoIc8nVAcA
4xoA/P7ZVK1q0u9cIF5vhc1HoKe5Nne0NwLuLYxGK9fVAXdaI7jvpkWRkRXOYBrmXKOcujqmNL2v
7s7OrsAgmPv10q05jwmfBzPoQ2rdlUK+KW3DtwDv+Cz7Wz73vd7fYZkxi1qa3IS4bjE34XEFhwPb
t/Wbi6XcUj7NlOEDTEANTlFkZ+enJ4gXpWPsvesCWW+rCyHxcjGVid0LSUrS1Qyw7v2lkE17hceV
CYrHNabofGu0brSYB+9ZWE7iTE83+Py2jYC9GumLeLojF9WozIe5v14r/5dMGwyPATHXGtkoUjK9
zddVlQw7Evcl2ScZcA22uz3toe0o+MCL+Y1egxPhAyfjeXFWhUxLpOehG/aoMa9RWs7R7DzZv168
ZuS6mOp4ACn0KicbfPGzArnxTH9tNx+HFtU+ofZublwkQg9CQAV6NhcsItmxf5D2YWJibhr3ttHx
cCi7gSSIBXE8kq1avSPW32AEH6H8Hqps3umWunVXSNDqhVJC3+/QVKIVTyiklIwqh+cKfM2anC52
5p3ySPstS7fnytWRiZ3q7PIyw2L2vJYBLvLzjrzJnHDulj+gyrQNuuFP0J8XEr9JR/CXJVt9/qFw
zfzXByEUykPBRLm3SUznzD5rm/H5cFRc02pOHej6XmdG+LJEy3fdxOfcJ4ZwUD5bqZB9gJvjV2ox
yECC3nfKDK+SPmwpig2/39h1+6C2qtlOTRjU8PSa+CkTktmG2NPPnI1BZsOlz5BCW+zedjoYPQti
i6l5ew7Ozdcsu9+KVFt/E50UR8bSZRk/U9FnNs5/iSN4BDJPO4+i4aWm4qRGq2+PfKl52r+/ULZJ
4hMPDqZH6crtx7qad4yQ3MgEPPUbylPCiUGS1RTq6vK3TV/FhFaWMPHJ0SKBadKBisbDWrC/X9WC
11yyP7Ux/QwgxIVn9IfPabY3qOXCnRJT+Q293T9F5bU4YPkj+1WmOjqVj/3nBgjdPJhgQ+jUUp9h
Hh1nBQRiMOltUYS/eUGIvqjr8dRG7o/Ugp8d/gaZkSOXMbkmfXo/PNqkEZdlhSylkukzkv8ntJ6p
ON77tsCdcg5p+pHIRTH4SavKr+NKd/dBtcTPthZYxfF8qUwMzNa9h9Y67CbVXWGTg3n3hkfwZgJw
xYBLwYWDJHpdx3QiWnZGFg3NHzPuCYRWyHBD5G6W0yergv5Z3m10Bd/2OJOlbopd/WOaYyKuZ4wH
sV+BZOsBUBJc2khjaa80P+X1aERPXVZlw8v3kj80J2c7Y7cf6rBWiFDGVA6ZKMkz/+/EH7Sd7UnV
54TRhWloT2YA/cBaRg4OmpbJ0vpOk9d3FMuNOPli2wwo7ELGPPIuEr91D+Hb9o7frcsxWGXPCtvm
OtEiK7QNfu4oGemCa6z445oh07XTbMJrwWWFLFUFoiTRzNgiz+0XJZQ2rpb4+iIOZ4qDnGX9LNm8
jm5m1zYYJZGJkYjrtPaEnbVfs4kKsEOEeRs6U2uzd3pdoWDL7hOeclhGesRcSQAOjKYE0LQ0vj21
mbjK0Qz9OcUS7jAUScODvml0aEmW/Q4h35eqUFbrL0O53mRXHNeoeIkwt4FxIz8ML6fGvXi2Ec9q
s5LlG0NKl+SOnkyyzlUx+iAN7Vv7SjU/lu+CBkSE67AKvvBswIdEs/gbeQvPmHzkYPqnZU3eYp3d
sMQBUJcZu5p15zpBeNh6Eh8RWTcMMFtj90g+36QaiN1f+wkf38QcpRj6VKUpHAEAvOq8/Inkf+yM
4a5R3r/xa8i5gjq2hmRHknKQUUS0fGxbqrvtG9PVctMYYOxTayW5Ou4CqNv5v1vqtwmPTLQB775v
tkOCLGhrjOiMXjUDfU3evczs9u0xuuzOrIkmoe9DqOiTrDn94Fi22MUgiQ89IXGHfWAieW8kFMfs
1Wm75NlS0ezqESjyULFxsCljCZo6ZTcF2JI700FphqGraoaNRNAKLCIUPJQwZ/yPRQncbjDTfLMu
UoOLISZLkFSM8Y/ouq3mSm3xpAJ9Mg2BfKvJ7GQwfDhwo9JDV2nB4I0qxTPmKSjUhPEh+I5OtN4v
xFArlKIjOixbZILSQLOP9lJcWjnnXmN6TAMgvImFlG3tV5st3G+8thUIWeKsycq5TTRpKSxU+ll2
/ptEGJ5sslw3e5RyU10FlURkkY7TSkVFDjIuruqULKaksqDD8M/NvQyCOAAGcNalJF6VwdYI3uq5
hLypIBcnCwWfTWcIXpo7Cnhm+c9/1vydSlKi+avtJmN80mt8G9EDe/ijqbqtGbhabWXW7npX/IQ7
KJwAyaA4qF5MOxQ5icXeRfojfwVQ8jpqyIYLVRg515SXSh6oK+u9gjMg12NWO+ezL5xBMHmRZXMT
TTffNTLMZoAZjWTOXVvP0Um/QSW6g4driDG4E8f2/ZFvXbAb2/ocA1CqlpVk5v3n/hu52e6Cxace
DjTkZUIeJut1d7Gzg5qDwafMhX8rKPX2+vpbwM/5jqEtvgVU2WtqRZ2pc6vWLu0Sd24l1yLAtyBg
FfO7uQGd+VPh1DUUBIXAq8+TMGu1mK82xxBEQVWra0onLkYigLJMxFuS4ZI9Es4hOGVx4nuxIy32
vTTDjNZnmBPwej2sDOMTgHgzGR/264X77yG80x7ED9Vpa0spwJYbUZco3WmS8ok9Bq8N/Syn7PLa
wbgongH4e6EZEGeSkmt8hesNdcgvr5XZOlXAbBksaNb2rK4/Yuy7L+lzPOnIk95Y17TQDon+f2y1
JSfThZJC2Nf3Yury61n7lqAIQurE6z7D8aYE/V2c9kqQ+4r0zcIeFlTpzazpdYkvoDpL3aG5M65h
zgqnbv1oO1GH5PXvhSVW1gfZN0ZpnmMO6aN/iARubX/SuQNcZrRZ02yR32Fqi3t0GzpzPrTJ5NdR
15Z7aPVQGN71I83TpoU6qDTcAguAj/3DLNQpF7ZwPkaCr3N/LgNIgrbZEh550rI67z1H97NM0Xmu
qHUX5fV0/ZfhBY+gzvOR/M8CC57IovUyfrRflsyo1/BfAwHI4D3dZvptfYCNXoP7dZD736pDdoFU
h6VkswR8628VX9MvkIt2VWe5q4hBhq2A7O5NrwLHp283Zn+MatfC/O1DJDxyq+X2qJ8qhAtUtX34
1FzIlELYZz0o1MGKiqN8w1boK5pBhwvIOQea2ayEY4yX/SGqEltwhSK9Cex78pe2kRMNchhH8AXq
2Ux1Hz6+hza7iK0O99tiaDEeSlPDUmAjdO2Lu06FoVK97cL9K5N/5LgsGGPGJgf40tAriaOo76JS
NfNjaDqfc+x5248r/AN5b905x4VD1/VLrfYq6pw1modrWdJpZBs/K9G/6Dco5za0UwtV8ggcxIU0
5S9rR0INSr34WqfLFvLDDIYemEdAHEcaPk7CK/kaBlKxbdLBMR8sWf5eT6VWtGuJWnIGsct0fN+0
qWoKRsvX3PR5cQrs6W+qyWfWWWnqkdDk99NbGnhyBTAvQBaLdKspw+dq6TtB/oYNoc9DGbWnywb5
HPe2HAbjBOHnZBW+Ef16guWtw/MoJZ6jD0QR6VqfCNNqEwQDotAx0TKwpcuBk3DBAZhcYnmKagEq
ZZ7VE2AoBYpQjbxJ/dwxfYkVt2t6RzavjME6+gsl6luO70yujVMpVU/ylfccW/h1zPJEvClEPD94
9dAssrfS5vIkAZ+OIEbdHt1rowfei7Bq+Cqt+J3wSJWzYxVetXzP65NHsA1nfEe5te8figcR1SiI
1aqZs5ULvWcczeyP6G8msvyDyMc8P+NYWbI06/tzfI5J0SsYTl8D/CAnsdX6skm696whz3JQQE/R
866xsJUKhlUQeouH5YKd/bjty3WfLG0BSvrw9x59HsX0suelypp3zr2fV/7o4lDoLv1/q1klZRfZ
lvTBSVOoFsAdmwl14FEBFszmYYWswAJ84HR1iijGpxFok4gcbnT10pblgt8O9DUF3sG3fZNV3BME
YGjI3vlM9mWWvYGNed9Yta5t8ioWYgy5iJtNpH17AsoBI1jGM5/015elF6Xk4v26r/K8QK/gUhQI
C4sm5+0AtgZy7aMPK3EyBrxRwMpa7MJV1Q5rTKd+0ec3Pang2PM2FYS/vj0JhRb2WAdOPwnYeB+I
yk8ZdJKY6+DvIXzUEVf64/mrRmsZU03nAOL/hLUscvy/Ufcb5ATxIccNmb3o7Exxsuxs5ZSAFGvJ
85uMbB5wdWf7K3HFyuO76u7UcmSLEeSvNoU1FlY8oMwEGc3YhXMcGNpsK9XjWW7AbiZ6mIVoslak
Ydo4OK5UfuhsPFlK0FKuaDp9OPIuXWXWsDDLGZ3n0OdmGD90M4SbJxkQ6C6touKMqL/NUVxxiGdg
hADA62V80L3JY9z/JXx4WBUGtPtRTvjO32nWIa1oHYktHyu+8BYv4GUaq0Hlo3f8af4idjvqhHOA
B1zO559icvT7Lj8B8tfkkF/aE90DoSHA07mEzoHkxFS3oAGlZ3mTFA0eSQR8dj1l2AWRDv5N9Ch5
u2gFvwn8z0KeIhSuFSDdI5rWb2G/6dIsQPUCCX1iqwBptDkaBLRae7QnK5WkXntcPiUVyaEp3zRL
eZWZaS9KvbITImCrRAi1b+gEKTLFnqUNzh4PiV2jVBG1jC8sc6A7xSWcjS7TehV6IBSdw2ve6usU
p5U90qWfqBKLyIaU1M+LOmn/vmHSfX+ts+Ym+Rmr6sg6soSrwWA08cgo7RyAQZ6HnGs+k/DFizO2
rYjxiHqUoXYQ1q0tELLrB2RTJTDx3vVn6LoGOSy8s8CQwd7+xppTZZdgiWYfdKUNKdzlYPrVa+wT
vHZyYxbea3OG7XF2Lajj+yG7aNgILAMWSey39aUvwijdmLPmW8e8e9acbfAdcCbi3O1QMwbS8rG1
hAJaHn8ByJnvmoBhEkX49A0AwPEnI3Vq8eW6rY/dezkQL8PEyVK5A4ARoYRk2OsGuOco1F9oVXCz
e/JkVjmW0TP+gdtvMeT6VL9TQR7yWV+tbkhYHmpZ1ILQb/N8a/GMZJtvprd5vGKGF+Ns5e45Etjs
p+HNlcmlq6kF8pJBgtQt1dq5exdbTbDYE/lkwgKx07BXWI+4aDmJwHJPNi7RnhTrPsxzPzYQotXf
BnNIBhSihYEsM5Z/XHzmQJo=
`pragma protect end_protected

// 
