`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16704)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPak/iHwVkUKXxdtqF6qlW2P9HJ89gT4zeosXKnzybBKQieqC/gfd2o/5DsPHAPbzev/0PcRz
xqOSTFx2cCO85netIcsPSeo1R5gyOfXUtUbsDtx9beEZ77ElHZlwEjrh1uzA8qqXv4qYnFWm3COL
ylg0gXiXGrlci7dIzObZ0xi3Hh0g54y29Gbg0/YDGwZpu0NMMlDWj92ACY/sabb+WxgVWuSMiTts
n0Jj469aPeE7n85MUVcFGnHpH1lC83f7c+yLXGHVmpNP/LBRyncGWuwzEEAVEK7fmnG/YO8pexP2
OTu0j4S37HZ12AQK6eAg8XEf+QzZkH+fW2pmcgAEnCsP76H0mFuYLN+AMFNB77PuRhJnUI61uAND
b+vL66kfesQknvp+xDJX1/PrJkMnUgqrEvOKh3EGbR7j9XMA3RC5PItgl7YIcEVcR5UxI4qFNXEj
RTJ8Ro0Wk9frjJj1IpMCi+pcHwtzLy5B9idmKFbCxAjDqPm2KyYXeCBK3LfyWs6S7c9iP3R1yndr
owv0zgKZ72IRDrS3y4i3JQrcjCgQAiWIBArGibNOKBTjENjNcgH5ce1f6T/xnCILnqwIEn7iaIv+
sLwH1+XFkZqRHRF/LPE0pW/KY1GDblGoZa6QyaLksKtsprakVBfrSYq9RuTEYnKaxUxy7xfIxKji
IZ4Cwt6kOt3gsAnknx3SpFeB3IRtA/qcpYgJXN1nB+UgYxDYa3yUIUCN6rA+dEqdJj0MHs1laNyw
ILl89ReLnG/H8WvBCV1M1ezW66Q3MpX9IdCp0Fk1rB7D109q+eIqctn+JA7KSBKYMw2fy5pH4izi
NUvltEqgrPDsW9FHU/1IxVB4VvfBYF94sVvhq1MO82ko3CWcRqfzUqMEN9LoV0JS7VYOLdofNFhs
rbtu/hMAEkbVXwUuxHYs8bmAYU20UG7CupzEx5ng/qw5IQsElAlGPj8oIuEAMSIwe2eylTmPkrLD
9sOrHT6jnumTCv0SUhrfYnxx9+QwImKLCBsq1lbW4YMHmWfTRlajpcOuZTOxAkC8ouV8+1+YOBjB
+B7A1rFRNpD2FXoisJMmnffAJ2PXoh49AgGLvE/41HGapMM5U33hgdzE8MMoUEBQQWE7hZouBoHq
+QMbwSpmsWZI0KVobil0vXMaCVj6TAhEfqR8XOUCHhj0sn0kuXX+t37UfAz5AHKd1/dq4aHw8oYC
t3w+YiE9iWAvI/cPLYAwZkbGzvKoSAQfPMlYXVOYvWLmgxRNwswIH4eiPvYShafjf2w35rYKMn8y
MpJeksw2gU9vEyioY4Kjbcgz8KLRjvmhCU4M30cQVXa/hrON7a3kRwagQXCbelCx5MeUOIPPxjXW
Fd7BI+++y5oTBNz8/gxhAr6EU0ngCzqEspgg0mos/zokq9DIqrvnMFqRopZ3TPpyz6mjt7hlseso
+l0k8zGRAeDGeZr+U86lBuBWxHLaHYWG65Pxs7SDZaxtUWSrzLBNdQFTI2Rayjr4IG+0HVQn1g3a
oxZyrZsisdFGyVW4++UJ1xYGlpLs8n95WAq1GxEBrpGSXIud6Bbt15/9Z+VxHb9LzQ3dUlJbr4e4
Dl8pAraLqxY15Kzsnhljnd5k5fVAhO4qUcdQ15zQPumInWF+xWMvX1ZdtB9Ej6Mawo23+f2Zf5pV
TFAXZRctnmrV1cCzjR2ImYBPFzhXDYKIXcchAlAlb6yuGBefnAtBDvDZzk/7M62i1zNVmOe4uSnr
3FQMQhzsgbcAbdvJZZAS1NLZQoOJIzKG8dbnB9FE1bpazFublKSLYCB2yYB4J7OaX5sQ+kqOyX9W
mwt/LgI+fkgV6alPjt92lc6CMF8p4iwkCLLqlC67joo59CvY+P4JXx6r2CmvZyYhXgctHLm59ZAc
xVIBagCiQUqs/x7SSiBOALd1VnRUCOs5l7tx3pscFJyQCVFWTgwUSLX65tf0alwqTCVFjixGwWlp
Azn/+yLI9MjfYV5mMo1lE2fdbDkvfUUATpXM1MiVAIHUL2ykN3gvZo8Fjdt144BPfKvFCL5RBgy9
ysP9f6EetZqyNjIxLAc9rsslG4XMnjiWot0zP2QkyhNlcHHzUC3jS/WfUWGx8HotU1Sh2lgtcaEk
enXuXDVjqARRGFKb6BHXXWvwzO55JyywKWSj5gEuInM9OKXIHkQcQGpp3e3pbQ6/vRj2pWhrxnge
t1NWaM4sVu4+RV/NgbvxXW7wbp5qys4y6rRwd9JxDTa8Kk4Be85VsuwKLObTQDHfwcP0JS2pSHy7
3qyiicSh5Ddc87PIAPFzRu5XDhMDbzYjGJvoBI/lmPAjimac9eA8rusQEaQS1xhOM/qKMHNupLdC
JY4nzINZNs+P8dKCMCoC1Yk+JLSPt2U8kErSqSgmNg+7VOASK/br8koISGlILA7F6pnIaS24kd1m
ck9Xky4D938QoeaioOEEtRde2nh7gOWg9zarJnz2ihsbogyE4zH9QCOE7JhEZ6Qoq+jPmBM+5HG3
gupoIID4DgK0IpmXoy++TZSL9LtqPjkxkVAuZEmrhf5+ZQhoQaFLRPSXhOZiYoLyCA8y+NqWfJFS
Jh75R9F36dPQ5GslMYSOWk6Qz17AAwJaRHPspU2e11KQbjzT2VOXxva/La8n5GRO1ZWn9VJaISJM
P2we8L+BZHoBLYAXXkmGPYafzxWSk7wYuwHMSFGWQ4rCop7EHup5cjXHl87DM3X5maOlm1nN/e2Q
HDsIZjClzfwdTpTjgZ7KwP6vQIZa0GxqJKObWoXcPAAmfXTCPrKCiHYXG/yH2+eN1LBRdFvGVX2U
87eY24cLwTDnxp6WAgPfZpsqPDRORFurEr0TS62lU8FnLFCey4BBhFAph5gp9zL3OrRM+vtQfvtC
/xkH6T9CsFpX+OKljoBdaWmEjtHqkOPT0FFo3C8i7OaCfGpVCAF1BGhNcRy6/0GVOxxQoYBawT+U
ILz/oFEDzyo9hJPJiCVVhm3Z1d9u9ximzBT395ighQEjn5PmRPfIz2nMVYfV1rr2QXM87RvekMA+
h0/1U3heSSBqHHPxV6PKpnUMSTa96QtxYqxvjdN2ioZAEGONVib97DASCDPwSsQB2SmYBbJb0PjO
WMxyDMjEO2fjMLW9Q4FOGtOdNnmYYIVdjvRT9mOUqIftxVyaTC1vYiw30fqJfbkxQE3YEKBKj9KC
OAX6LCTykgcpNI55dNbVLZViMTNacZnV8VFb9AwYEl+OjM8Q9L2nkmIl+REYJ1asZ4mQYZir/hpu
xaKCNUUW0bxZ4S0BGybiVdmxXKGxn0fm7X3u5cWAc4q8p5vXuwazWdO4yRO2jlfFmoA4TQ3DdVWn
Y3Uf5bODCUK1zxfYyKR5pzqiesjIYfaiu5qEm7VEOTzuaLOXqx8wRivp5D34Ileez/+0OkatEWFD
qTtnlBniIB9W/U/rYB0EcCgieUJahBsFfVbuVzclrS56CQyWt1jWXYCBsVOX8Z9gvQs9M9G7A6L3
yOAY4CEmXgso/+w35dfeLQS7p+J6BNWU8zitClibWckAubiNafIKNT3fsds9xD+dEozEPilIUqG5
iLAXID0CVrhlenqfKfJr95n55xGUMYmdBfz5DgO74Z/3SuHagdC2DEbkV/4ro0ko/he7MyNpApyN
SmbcZIRhdA2uxDtLe9fIzZIIEL8eeiTbFdNO5IfPsEPKhKCKmHGeS/KVfSmThGLlNtewjvhpr5Ak
wrdnJui8+IuI21xjNAsbphOUd5WUTRSAPSwmammaUz8ep+bbVcAX4ZZ9Lr8s/CbG0sXQJNUXapKj
GiZYF8ty2Qd/pt6dRlKmZL0wQ+NNy7gduDNyh2cK8KWG0HEjxe+TkmGUvFUkh/My/nVI/o5p6Qkl
a2rbw7UyBlVrTOA/9wAd7XhqRuSuxvQPTvsDfU3s64S4Uj6iQrJfg8VOTdcY6QOoR8hNpj/vGjCq
2N60PtoMbS4v7dyMccXfkmcmWPZXdvydjNAcmZ0BAXdV257e7ToM7kNAHQf6gCelGUa/y4ZNLpPn
ui1olmnDpUGHvaLkzeYmVI0WDrDbNxroBsP4Gx2sCfPKzbYML4yM7FIIVh0/9WL5/Y51XyUa9y8G
QdeYB9e97w7ek7L8O4RJ2uFXn5418+WbTMHX5s/OiZY4L0jhgn1o4s4Uo5p07/H69xEOLFysnURi
lHxQmN5mccaMab39CXdkTQGKRT5FWc9l23QRGKB8x11XVen+xEwecRuzkO8lyJdXdKkAzJ/vtUVa
ZX1LwJXCLN0qtprIHWpUvsObbzhN2vlUsaNV13LwGokH1uWMs3hEJPIVC9zSpPf651xUKknYWQtq
ADs/OqWOXU8okmDh2bpjtADBiyJ/v0h14BHHahYJEebUvZrrLSHvA4uslAa3dEtxiLU6mpD7BSFR
4UDHzTI/uQZfMN/UUGW0ijVs2xC43YitLcCSWJOloMOd1BqRhHZwueFKpc7yzCLy/GkEsLN/P0lE
gsIq9XaRiAWpgqR85D4VBTzmwKR7ULwR3Z/lj82Ts3zGT7IbMf247DeeVJVjNqEEFZj5g8LI/jvJ
IY8R9kcrLupcqH4IBVchT1TVGBu04iJEFCvf34k6F81jqChgiDwC92hxoAxIpL1j0T0ZYYA8eC+n
XhgnuTlVU7xP+7td4zmIKgKxhFACAtv1eL8hZUeL+quaaP8Q1esko0RRXhJkXqU4CJKWJ7ZF30PS
+ZpqgppjrytH6p2LAtK7Z0+BYP29TJ/IJjlfSFiCdnDmfU0F1YjfI5n99jPJcGjYItari8GuL/hb
HQ+JA4DroSsQgn5V+NI32oF9NDAIsnSU7PjsdNT6xLTshk/kEnUgAP2zVZOBGrmV65XsPaKKatPj
OFvKp2+W+s1/+ispGHiAJWWnqLN4Mftl4+4CgWCqJmfAJzBkC7vxt7T4GPC3h3zqE+5jcBv4U56L
QIHCXLwutIJL+llKIRElowqZAZD0hdczeOBLWPdOxEkuQioq9fRS77j2AS87009QMC4L65LVtMUp
etsVUWV9zX8mncSOpOYDss+s805NYVdxRH0ZOrl5e9klcCuUBYsd8iJ2fqQXEimee9z3MBhUUo51
f+hZoItbuODl9dA2WzGn0EUpm0MvjrSe7gBXqkMqD8035NRi8hKQW+sYUQhvTucL7BuatqqzHAoy
Vd7KfWjGGCn7pJRA0VOgVWD6sYwzTlxgLLPZa66bsV804n4rnpJlnHCelzlCEhaFXOTIwM3t47Fd
gLLFurxoHqccLjvZQ0NuSXkc22LyS/AdMH6IkuyWQm4HQ1lXkq3hrD9iCXGmbwTl10pNCl5ee6q2
KflKTPquVnJqbiRaCtdYC8jOmPLBQaOIpsZLQmIRLHSykYj6ekPU5Haujl72B/idHhvdQ2fYg2pn
6WlZ++QRrImuTWl+uVvfH+QA1GxizJ5C2guB2bNUAluASQV0L2RuhSRT8p2fPGtzSEzUp9hyMSg5
QZWWGsgGjYnI0vjLNjbGM9P97dG+gh4VIYPP09FIgrXG5k5PGZZ6GO8Oypy321QevodDGTnaQdHr
btcLUqnV3jb4ngDiMqwUkN+Oj2kfTV3HI6ZpKZJcbutFtoB0Tg2qXVIW4eXSLwx4BscR5Rk257nW
Qu0TnNhzLsPOoUBaHDVa12gBcxSfBhdtECOZZzzBFt02LDdKtw0PytjoM8eTGDaoBajL3tMEgzW5
sYGO3SYs25ojzf2chti08qbS9sGPbVBHofWv5O9haQONRtzkjSbxvMPkdlzJ7XrVhAIgmd47ZlVo
xssodTbcyrcZjdNEuArtxdf8QbsN1Dt18cO02g2c5DlK8tR8Tu1V5+x+eFaLSQkTg5Rdtt85z8vW
ITLR6+c/NJ1jDgLZ32J9W1nEsEbxu9WrtUbmO7K2tQzb+OPoiQJHu6wnw89+zRLw/cj0qS7EsJw7
ftR/M1Lk5AgLefQp5e8G7fYr6XUSTa/ShkxMYUDdSTvDkPtrBmIpk0xQ6OzflD/Op9l/QINHxdVU
we5mCt+v1CP8drEo9onBZwNzWTuVh+3G4lajX8YGYjadzPWJoU5uDYeCiI3JevWQHEUhLiu58ah/
jedkAMr0Mnxra1Tn++Xbvja/rdmXPf6RbjO19lJr+Jo6Ush2YPNZhmKgC88zN4usOwUaq2R7tfM8
fGRSiD64YJ1NJSsv+/WI5dHh4PnouLMEG3jfywyEK/sBxRulOfMCq7+FEZQTT271I0JPjW5JffVU
vVoLhZbyp2w+Zyz1eODVl50JFJqI1auH+URRkswhQbMDm6c1I7/Uiw6gmKmdDSwdM7kSTBxledFr
bq1PbFnBENTX6/g4b+mlai2gBAT5TfrapmIlqnZJlEtY59Wwsfb1D7kEQDrdjQ/e3x73dE7XrSRx
xzkz8hUlL+7DBawlQ69vlOhSmhb4CaDGUva0IrpoLi+wL8tpN2FRfN6ApaGYIEGkmgRxc3Jx1RoO
OLJqDey0Ak+45lq1xpqQwXo/rqKfe86nIF3FfD09lNch5OqGKi2EWgzFUK1uj5mcCgZRA1tYbjVR
Eosixa8OwsCHM9BZQmz73GAjfl24jYjnM/QU84YAG330BAkDfWMlFnR3RMqV/0BWuJGyOrpv/X4A
+5IUY93bkj3zi42CBwAzm+b0dNcEr7HfGFDinvJylk1mvnFViz8TksPYeXCdQUSzpBYj1tYEPju6
gDkA895rl453ZKONXaB8C0JSd5UI6i0xXufAgKN2q8Rx0AqftIESrlomP+IMqNhQkRxjauw90+Qn
VPqCMeQPtmu0iXrXL6Ptm0jPLRGfbBHV365sSamzK0R/9kQgv41fPN1oSHMfenG7wQFxXD+j9Guy
/dEuBu29hkafb06HTQhUPTNO6mMtPFlVYv9M4+3gU6pCw8ItpGytgBh9PKpu14vhfJ8sLup9d9M5
AILvuqHY7CSk6ToZ0UZhPHU9AbXniKPXIwKg/vpHlT4nsJ6Eg8gO1QxFl/oRJ6DUrcka1UgKEIGn
+Xp8wg6PwtQRfU/6WmGsItZxCzASmjx7UoS/46yCfmjcbk29pbb/vnB0RCnVHtPmucj7bZEIYDcd
jTKYRfyD5iLWC5nuUah3toUVijvtN212xl7fjlzwEs/AV7ZVpfGo6drW0J0L9q2FHBYYY7kTTctu
z5hLUPwWsl2PBgvGLPE33wlQ/lBrMvQzRWOcNhqWZEV8ytzv8t78eCrZD7W0wU/3dFPV+IGI4/0I
C+Thn7JBtbGlBlKARnPd3L4A0h7wLh21Fw0GikW5TosswilK/cKAEWtJueILXJRDHA0vbcnCM/5Q
Qg8FPHkjbexHpsa/2DaOPj4ryzcOwMhqVrh46BovX4UrA+pWa1tBJ2RgDOGJsZaSF83KOuKXV7+x
J62alcn8WxrQ/mctTqFyKl+1slPP1iMaz5DCse5ezxVWTasgQPaDoinHCP3Olnfwosvj1etkAPIp
7tsPfkgGfuzcHEREWAGFIa7sb3nkUAT10nCeEWfgSpRv3og1ZGrYIju/c/GUJn006vK/R3MMTHiT
IEF5OnWPjEfVh3thMs7Vd5RAuc5vM2qW0Wn/I99vbPAPFyEOpWeZ5jzpN2v7Tj4Tlp+CfROy6QIr
e5G4dHYb/1WO+vps6dfSVXX+qYVPcZmFqMVFoUsKp/5yA43eEUzkz07wxuCjJ3KLNxi3AeJ/WpvO
EBFdQo589ANpW+kRXEjLgGRHEtf0Q7HRtAXrJIP+0R0AKkwfPkJeeVvA4GtDLr3DEGPY8wI2ed/q
y2/+OCLVfSR15xZlWFp4PXcVi8OS3X8OgzN9tJYF92OG3ldjPhufFZagWgVeFfv7bZXm45ADtzIQ
4mAtk9QOmcgYSzwv2mbSl+bQEVKP3ix1k74Xe767kId3lEErp9/NAsVAgTI5u+m4uYKHLiLVLa3n
4KGhjv6aWw73HHAriiabAXqNdR4t5VAMsDkqQ1CAxlzw5APWh7GS3uYUBGycCm5GqLqUMH6ryG39
E/m3E+SfTB5+F+YArdA3gAfdg8z+r9ITJIXItxMguiwCqmVJPzzR5rTp/E+DEEkATcv1msjc+iVQ
akjbcidW+xZBsFqucl31SaJTYiKSOioFBqvpkdn2ZZJM9LqOFqoaccAFKvDsX2RfXQV/ZLu02dhO
mMOZ2h/w96UVUs9QamxWrnK4aNr7NDvve8aKV211WRBdxsL+qfhYKr7bKMLTAODHuZQeczO/bkG6
gycpPTXOkPwfPHVmhDWf3A+dyewqnQ+XUBQfkcHZHgN2O+rMnlfFGvpiMzfPr8k+nMWtCsfM4i7q
K/ReqcW5l0OemeqpWhzIn6qqg8ApKcGi529LXW30UpRhvDxXChq/R6ZrwZT1oRs8rs/bs6XvX4Fo
Yea4dz+OYso+AiHyTgAVz3kuON1gyVirVy3QSjmmoyze3GPgjSmptShw72LwvbfqrfKN8TSRLMiQ
Xi0qW2xrDCO1MFQjN15bySqD6hNXX2FHQz/qpYn7n+rKWVVkSoKDKtoLzonNd690Zai2qEQKE8bk
F85/UYf//Gz5PvlzV5LmdmhAKemwFCNv5NQjo26eeo+osHG53uzjneqQpqB+/tmoKMfIFnHCXIUS
+6mb9L/US+I73/i5LBJnaHUPNOWdW48R5gMGEHyhmYfjRoDMRHUQYykHTPqlCFFuqzskQXTa7MZF
IOK6N2QRBO54GDXBXb2rI4eyU9HH2q8V8ZpH0j8WLz1KhheNYOZNWkpqQN9PumlJbId5MQ+HW8TK
m3HAuE+v84d+0jgkK25qmX22E7t7I6eSS+OLw8a8Y/B96f9WDl5IJ3IOwTRi5WdsdP5KY1083pJk
3TPImIBdwaP4MOF4PdXFt/V4dOoIgMRaDCiF8qh+ynvp77agShBtVe3HmHcBbKPTbBaKmzAqIKfy
EX34kvMlBESoTrqksNCAuFiX3Qi1q25zuMjOA1oMut2tHg32iyeHT9RmNCw8MmtuBMMHrCb7ZH7+
BnnOyfs26FOe71f/6f4cP0q9zDLEbWZh76sb5mIGkBR72TifFX+q+CuSgvoidhdC4eSkSOFdEmU0
zJuMghrv0jRMA7zha87Eo3wmHZ29RqGd4OEfGh6VKEXgcdecO2dPLfCEYZgLIq+Hc/jPkdzee3l9
mEeLcOflBcQUHgY2DPmi+xM8KYZ5aP5p1IWeKYjc84y2fc6sEBmr2tbSOXEmEMXbRQzLz4ojX/us
ci1wEh1xeYilca/hBkzDfwvtq/PQ/woLxhNUEaEgRjOKnBENK9zeCa5MZ76Zb2JTuh12Bn9GcyDw
62jocDZfDnN7k3/zkJsZwf/dLG4gL7KeQA8Q3JJcGGgFnnTgzadgjYw/F/PN6S1KJFxQC2by8wqz
zAiG2UFauaaMnh2d7cj/kiSwaj+BHCqKCpsVkiUVQmc76sDNJzEWIJI7YudNgmA3SEveKG+fdS6Y
S6l9rhJ3bMeM4nk0/pRBiEjPIc2NT8tZwUPlrvmFexzXWuziOXhPdbSAOsJ/uRp+Jt6R9FrYM8h8
z35TXizTLqibuqkrH+iDM8n9rrub+F9TaARMZgxBa3kuhsU29A8mBGuY/4647Rix+RTta0ssDRP2
vF8tJf3B79pDWfjOzG8jB7dvMd4WAg1vg3BWKfOs+kRSsdwMSA1EZEAp8gk+jOCh+xtzLL3MAYBI
DWYiXEOZTTY/oKnbvIS86Q5uxPotfWnQRxXn9JEl46eB1LHVU1FhWQFPLmpVZ+gFAm6ej4EcMpOB
5trEbEyOm5vwmOhDhcJV/XL7ud/+TczEBnMbI5BbZL3W7InSV0zL5C1X1vg0acPcJKY2Q0FkHd5d
wc8xZL8LrOYRe/GeNXg/37+MtvqkAzB5IESP2WrRb6oGqir2BBK4UE/0q+jsc/2WKPcnM7R8Yj0V
cRnh8gfBxYGMm64FJgL89B0wXFSa/eHaRlDaXQQl3Wjhih3AC0aDs08lUDZxpqCjjPx8/NPEvuzu
S+ViWCkK+CyGVCA7y8bmMIO0QdROx2hNa8K6eNDmzZfvVl/qtAdHlVT/89YsQ+tu3IdN5lrdME1o
Pg92GOcR3y9TAb4Jl/XMWlXhZyDQ+LSM1VLb/9kAvGQj2RoXTTgoiU49TGVYVtIYn5NkOpEXqzgT
LXLpBPSRUnfwtra1V1mlHuynPA7/VaOVBS4wotbKK/3oLzbUXwl+uXa+4b/k9EWwNSaEdfgMviSV
RZwLsn9Ani1qEn6Gyd0bjstYNLGtQ2Xv8ytop/Ffapnn0O28fiauDjfY0fqgzVovHwhPri88jBrU
3KX/5tIQfD/npQ0WVRJNDAZGcuOQTh0b2BW2/kfXTbck21mWTzECJvJdxLA6SZObEpPSoS6jqyzR
I/NwyzQ4zqDnkvijX8Gzab3X3cs4kdXjmSXioptXOFrT28pDr49YBrDIVvGsl87i5EagGDIiv3EM
8CbZlMf26LAD3PC19fZuFA8qH3etIYoR8zD1MGzQVf8MVQZtNf1157RMispR3nJQX6ErB/+EklVF
j0SjAT9BszgSAV5CTrM88wnuR5uXMmJQYEAga9m3486lqRpy7eyqjQxwQ06o7703GbsnExeJQxS/
22hDW9bAUtJXIipymVbm6UrjzXOyHZ8DJYsT3bCZY5HhRYLWcxHYWSJy7O9EzbBUSa8vhtHNWM5h
Iy/kp2psza+JZ1ZvGf8i8zrDtfqlvSAVsz8fPE8xobYeY4od3CbaNHfQpz3wAaSxMuNqmQU6t+I8
pVyJx76XK/E8S5gOv25FftWWysYxzi6idLAJxkHxGxbAe0PKXGjJv/TB5u1KT8b3XCHxsr0nFAt1
yTBJELBJJmy3SFk3mehvdjjtnikmmDGmsZ3G1v+fF8mRQ2dgcIBiNRYjXsF+F9u76MI0gNRlFT+G
v+VoA/oon7UX0PM/cE5g3o17/mnK9jgBx1BFXE8t/EutILxyE/E61S4/A3kWq2h/6EnW6IL0wLqW
ZkJyZNJfWoZ2GYk4fSab6yzxkc4RCVKkj2l9WGeqqV0o28M+R5kTia95KE01YK1s9Lyj6Up9aaFv
uW7RjbW3hcXwbcfw/C//hSY10qSLwmsSA1o89hlRNZcyOj7HV1/Fl4QKvQngHR6OqYkqBCfJ9/IH
XtdJv9375nHvAYe1+BPMKPW7GS+jVVNRR8edUm7yy2TE540bTWZjyKpnIpU7jai08rfYSPb0qQnC
HF3wbrIPCLh1x7Z1hiufLZsvFNPOpicTCakZtLbctWEvzj/YeZApMp5Czz8yTcLdXZa4OIPjwar7
wjhjhtzHAATt/gTZ96om9scWwk7EkMWlpps0Mxl6exs3jJQvIDM04Y4OpeTAH6SdSuytZ/OqfIv1
gkkg/Rd9fiaVoAnOPc+yW3aAeoRcWLoheCWU0L/TfL3UYW1Thwo2zdmOxSIeIh35lMF2Rg8V3/uY
VTm2z7On1UG1lYhJCjjb1ymN6ETxom1eIFgODLiwzyBY4hZY7TV78FK+kWLYUwoH9gAftt/TJF0v
ispuTgWD+y37m6hW5H8SxHz1rw6kjQY9lIw+gj3gbXQwkCbzJL2hQlRKj1LmBF7EQWy2u2PZEYQo
iExvjVztvcog9sb6xb+uuXj0qnQPY97ver6OiAcyIpF0MbSFIQMPHRRkiLq6oAsYo2J6ThZKFy2O
+2pJsDZu/YOwED0eu1AM9H6S7mr/idSmLwE3l/leFMqT8MqaYVGzKRKt8rR2WiHTWru5siWon0y3
Hh0DBfeAyND+TIwEziX0YdjzXtk2B2Q8QA0qjlQDmX8ylLh0MvXmj5hIRO6fm2n9Te5t6Nk+7vFD
oT3YIbtu8+V8o8u9j7HF5ZL2F5oaKTWq9L6e5p+/VcvRQ64q9AfJA3/w8bNiqMTKvIEh8EgUhkZT
0l5NZ5ZhxUZPB7UT/TUJFrV6FNz19wxtQ5ZKbPvYmsM0PHx/1rDm8jBat0lUxUeU+fju0LmZN2ir
r4dN2qeTii7Jps2hWaSVThvxM5TU4H9eWCC8YYWt9CU50TB7dm+ax3wz81lTtLCmEA9UzHLiCK5J
vytG2vJ2C6lxMZDUXCSoFLj1ixHqceP+3omaF19uXFLopU1TT+5hKElj7DC1tHfT9gqlhSarcNoB
vythnUTn7etBKY5CR0WeUKf5GwWf63wt0LQjXzpA8wRL5a5NW6e4NhAdA2bofTeSFgurztkdubT3
9VAnSJbFsr2nSZqbuHdLd8R4EQxrXKH4/ZVxGwWUKQIvvKEWlj5PulAx1W7978SxEF2v+jXQWvDp
PGxJVhRBMoMMDPC4Qr0rzy99xWwIJeFa8pC6WzXHHQj4gcEZG8LghU05IDk5xZQ6VJzrFcJuh+nD
g6z/8UT5l96YN+cG8J3M7geX8KSuC7wToYelCr10CENscrc5AFCVeIOsLwS9TdSeJZRYviIP+HUK
LJhvY+8Wbg5TfO2Ay17XjqZ2u75oaD6y2S1CRbTREcNezcINkKx1uSfQtOiy2M0a0+/7tSweFXTW
V9ILcgpkRRy2vGao+yPybmwbQkCABw2dVefuJkKIHifH4CKtZIR3rjezxD78hf+JYUpjpzbglTnu
M5xq47bQTOB8t7gLfVyl28JHc9va+dkMCRiPbR+YymvPaL7BupQPQ1YT8oHJpA+pl7SnThHtD92O
C7wqOrAfAjwB7/10hq7TRrEWuuU7TWL8xP14yJLlt1KwU/I6E1flCw4RsBTgU9VqoRxKmh1iTVR5
89jlCevWr3xQLUX35l6y/KC0voBtNIVOTEX1B3TPtFO9l94CRzaH8ZX3o6C346LK5xxv3mY/+eg5
6Oyk6HlWLcjBq9aygkqDTt54SdFOrVg+12/c1ww9hAmQNhjrTU/dyucQFIsZfHIxXlfsmo2eeYmw
M7nEC6c1MiB7LcStwN80jwQcWUB+AEeLyjwG3VHEkQpFGF6thdYlfKSO3jKgOyHH+Cp/nfMY9otY
LhQPUw0y75lOIw6c+ThbMGNVfzEK9c+wmHY1g5Zo2jkeGNGbabxwdlg6cWQpZl8GKgi5Dj12m2qS
tsU7wICnhdiKIFLSoHSdqZzYSx/Y5221d7wZEHJlaVb4gW0aSK5G5zXmlKEdhUNmJNcMY1fRT20A
oSmXGPUOTZ4jVI/JzRg9J9de6QuhH41An0d6lvxLBuHmKYdpYzOMGsZiN8DQgYip+xwqcAU7dh6w
Woh0uKNnwoEN3h/icdG4y5aj/DDLLSK3Un6cMUFbByIvoDyP4S+WUX72T5o/zuClyCopvF1KzbkH
D0i9Ok3RE0BUqKU3MYe9bYyUl0aijYDsH63F+S/5PJXOR27bpNxJVK4bQ1xxc5ljKQLJTC/svAHn
QpWUxkGZPY30EosZ25FsPWcOYRbWFTHeuXUhbx6aeF0A7Fm+1J4vbBBXDUZLpBIRUVFATkwEt9cq
D5WnwRqjDWWaWKK4lV7Egj9yINiLJ4R+aoA/1TmaUFgfgI4jjs5f6x+sJeuFGE7pCD1RtHXpq5DE
0aWnNMLyI1p2MEqQFEqtezFbe5BMEuIL1dQBbuDIJOE6elia5LGBRsrh+l8lbi9LLGFnqzjjCBaD
ro5GArweUViaAqoISosV2PhRNly+/5NFMCDvaCSkP6Js+4a2Y97q2vQ9js5EkaHQXkMfTQoALp79
mP20Q4hTN3aTWCxTaKZkHZQViy6uXOnmc5+zGi7TzBxZm0B+LZFmBRIZirwZDkh2hBUSen3fweOs
oCCPKPktNBIB+Q5WCPHH3fVYBgj1uHqIAVNdO5mAe0II9KLW4P7BBrD/dqAX3Qj2Uxxfg31AOjz6
1MYk4URdTSBxpgMtdvthoSPzSr55C+qtQyFZqGEUCSuwPW4XLNBjB1vVu/GBsg3i4yfXfiAME+ul
D4DbJldlT8eA9QjrsKLONwyWQ1qRpepLi0Z0yrmG84ARwykCUPLByavpOQ6Wk/M2mUI2ZbKPfF9Q
g59BxN8MsxN5dSUoC0gkDmGlt5GEI6YltMJJ9b+Ft/gK3xWmuua7KLO0vcfUZvp8dQcMhkBmO1ve
Lj1D7Sn3/FJsMB/G2Pk282npVsTtdXYJYjSf+/jzkC9T86YRQsq2Q9EAUIZlAjNoizjV01eBSp2u
A2axJLqWhMhP3771HJ5mIkAZlD7T3OhhkLCpJmITcDngof/dPBopjJUnBKgZx/beuyuH8b8KW3Z0
Q8qD91mwsqdHwtL+uocKjjnOD6fWaK6I0lfwSYoL4XP5++TiHo9VxGmwTl/3xghflN0zXGX+VK4T
VayICgqFCuL0CS2Xfe/HTORybygTjTtcsI5WsL4HRbN7trpHY4dok1Lot8Yndj3lDpysvCXcKdQr
671Iu/LlKmNvOBIgp6VEImUt6FSFhA/HJ4g4mGhQtTP7ILFXTqxRBW4LBteIPX9C6Cev59YRmFiz
/ZmoWxxG3emBmqqf2ZNKzF1wE6xm0XaKrZ6lZEBuRvyJaDpHik5OnNauODJvyTE4ECV5QBck0rFO
6qzwjeqRbdPL/wEiOppcxppj/aKQ4q+hccMbguIx3/5kGeZ/vdCGTk5M8NEsAUsoggKHd9yEUdJP
M2fqdGUZ6UcD2SSlAZhbV1Zw7oJT/jzgcb3MqvxW3rUXxygAhYnvt7yT7QiGyYctuBZnRx8qSqDa
ardoMmMhZwda6F39gFUjnbpJVyOUi6MCx1pwSlo+m9TaT8h+p4ptMVJjJL4D1lMnOe/HvM9wQ8ag
A3vzk4k7Mg1InrNU77C7bE0QSRuuKNrIQZmQJ7NimP1/Oi6ZK2ZMtGgjI3eJ9iuLvCDjkZ+vcKLF
/yI2rX0iwt0aGn2fHTihLVPtWl+LEe7H6GKVjf3RGaxTbsrFHwB5kIL20to2CxvXT1QNptpgZwTy
417TZYFGJiBvs00tFU4kvYZOUliW9zpjVrehLJEdfE7B3h8aObum4TCaaBlty/bzF/Tww8/59rFs
OddiabNNZAsYmscivBGgqNbLL0UGRQcd08Q84Rm2q8f49lqVy3xitqgPo1RuZdwalIMa3Q/ixvt6
ocWIM2WkKmT1OrRVXRICivvsnmTETjZZMgx/sF+LIwTQgAPuWcNVbwv4eR+I6O7RmeLxE/2JwtaH
WbAbr29df+Hy+5zf0W4XYyndYDBl7d0G7iawQ50nUEFncbAR25QI4R+q5ph7KFH0l/PCDixujxxt
zOHjoFeZalFfsKu/Hn525B+p7Flkt21mU5eOIXArFwKYSQ4/50aqfl0oswitJKt5KcVZHd8+qWZq
aQ19T4W/9wMbiI7ktiYoMNEu1OsJqGRO2sn3kTdSkvMhYOBirQruI8Vz6Rsz4ISuwfMjMjw7XNNT
EybKBDttf3JqtG/2kzEfrtcejgGl3IRz2S+BkeQbVNt8akHvSct6zuUmuhJ5/JCQkPIl8TyvRXRa
Y5O8PM/t4oXs0MaKX9Ar6ZM5k7/3TVEGXWPKduVg8cMKlW3oishY1ZAd59HSTHS1PxiQWP+gXySo
5N5exZxG6wZ1Eswemlonju1ZvLSEhZTvNkPG5YvDznSk/cwqw66U4httckCrf1s96tmG3p2KWNPM
5KwgBwfHvtw0jbnBiy+b+4tCdmx6yPqGssmObm823JLXTOBnBzbazl07w18ux4VbWvr8TsRddWdo
pBptouukj8tJRZ6jIt1ffB2MZRNajAEBAhL1kInBE84Num/vEw9zwP/E7HkXmq8gloY9FSqHIwuM
Lh+C+Tzh4p1sn/L3JOwa7On6ZpWcfanicC3Im2hTBKBuIlAomUuuOcSy6a7abOqhBzLRO+p1DCJM
AMc3ntKiMKjf/j6vo+rhFqq7N6dkiJXN0yK6rtYqDHqinHTvjCz8wQM4veNev0VaqOQX4e//tYs1
sPNl2v2qRHVFoCi8M+z+gorGXuUNSpn+s+JxbYa5MInPsO/lu4jjhL2PLBZbLveU0836KZChUVpN
6NEk/zYd0I8bmYFaV2ZwSE3oopWoUQAqvnZkb+YUu6LexNQR7yUdAdktil6TsJRsMHCHQJow+2oN
O3MU4OtkgjodXD5A7RU9Cm91Ch5lK11tu8oWS2PQrlZAorT3RkH+kRcIlxe1MRHrVY+tlE7+M99C
Vj4Uo5Olh09DGI9Tmk1ORVwCPE60n/+w/IRma4gHhEz4669/RAmn2updh3ydAQ3RRYPlDi7mMzaQ
CWgofAtBXdxX+Jyu6LIKMnQ/LxQrqtsIzeR02faZeNw7HNRilz5Fqwe332h0hO8mSu3KZM8yjfq1
D+ZOJSuu9SHzA6SpSlOCMvT6zVI5yemhgb9sCXCee6u4x0VrUXX3Mgc3mzeeAysNIeA1YEs9Z6fk
AjPfbrAx8DZlylSYAr1pXgA8m0RUWWCV/53D7fBpCl7Gvf2HVsHMUK+RessKluVnKKZ6T3981Eyq
JHcNbbjZN1wdtRwUxIlI0hbYp86Bp2Qs+0hOndjSrjP8N0HPQEQsOfaS4XdjrdLXTCdbgD+kkOed
4hdN3AAV7tnF0m/m/62i17VJXwXdGNxOeZmho0wZOQFn+j5mvt6RFSQtEQrdRwCj4X8Xig/+2S65
ALsZpi1JhKUqaZpRrRNW7YOIF/bNmECdDzktXX7lN2dOpGbr5uJNN8hi5oWWCkt1/izg+huEdsTu
+eOyltOC+GXFmZ6w/ml80ZizRswrwhYSOVIPg1X/Kd8f5ZDXRiaCjxUbzSaT67vYKyqGJbRGL6UC
abaySPlCm/M0d+QXjAu36zIZAxX/FimtuNOJXf2WBenpYDGy+mf+aYrLTkKnxKEQdtGYVonLuqq1
XfyrojFTmDoeuCPJthrSUniQdzLljCWJPfF90nlS67hm1zFWa59A8lWkkFHDCtx7Z9CBytMSFsuZ
e6vfHLIsjW7e7g/+OomoQShH0I55U5OM4jZUF05YGzrY8Alk6GJQmgRMV1ibZxPX4jan3HGGX44u
aKPMbduQNl8EuP/mtIc/I5uWoIy3B+dW/BQmqLioBLCnp/nD30t+rzF0HUk/7VWwjqTs0JPoFzUy
SMUQG4STjaXn53blHObAlQ2sjUNFSRZ3FNRVcNbPHrXDzAxdDNLo87fUi/xkejtvczDd0O2AsoQB
pXnHDwM8X0oMqZVjVPs/7/foJKJr6laoDl9qMbm2Rhpmi/TNezNyhQL6kTyoIqemWNQzqlDs5VRY
J9jivyC/qIAbj24wzKQ97fH/bb96CB8VRE9RM2rZAzVDGir/dMTOMopw2UYkImJVW9rRUMsKgzFD
DTUbd8gzzhlT02QV2exLauywJLbgjj7+NMDHs2qNVlf410XqdeSttuBxyAtpU84KX0k8Zag7jltH
l0Eb5md0DhcoC+KGKIs1pBFrAKAHPRYt1nWgZMhhD2/Cr9dKVd6Jkl0+aAMcsA+Vy+M7TX3Yz4Gj
MLewH1wVMV8lCP8s8HYNDNX6vtxRX+MpgoJjg9PO4ZWFE9bgL/qAt2SsT1H8jJgt9ZeYYk2rIooa
vmUTw9805pG/hTHHZlCDG4NpH6wYMOKWujsMg+t6CyP5oqNYGGvbpL5cGIHoTanvAoC+UxPACB/i
iOcvPtFLJgduQnAQuV4cJeHBhT3YfLGkjcvp3sLDdDDhaZGRbbzRki4J53xLuM8c0U8O7G/Emsqo
gW1kwngD2EIe6MppSeH8opTtcdgoMi1zldZt/cQ3yt0Db/6rSFAVaKhAYL68+Mdwd7eoCFCrO+Qv
tJ8qQRql3g6yqjU/4ywMU7iF+yHJC9oDvbsWkfIwdYrT7iYKejXtapbZuLpNmQ7Am88ghxaQC80V
+eGLr3g2qW2xnj/enuzFTJmWhVCqR+OSRLAgDvHfJRywh7Xn4f7jcvS71dsQCcCsUSfmGLPVLyqo
LtX1x9UtKJ7Qttof4T4WOrA4zpRnatuqI9qnd+6eRQZmjC64Pgpagy+ddfpeenoX0uaLLRtxE/t7
PyHcT5o8XMm/t1ESy9yakx4EegnojyGhYBm0JDWX0w0abpqNdWXAPGQrKkDVhW9VNiSn0bDwgs5v
BlRwFHrutCE+ul8yxLHzINytdThsMY57vJtLVDBrgX4FxxjPtGUJqz3WOnTspZ3jkWIX9yENwtSk
SGc89m2m4535TKwblZ8cRhwLjlaRjg7wFKyCBYkSPGgnLviOcvfzMXIJBYzXoZtbIbtJCvXsU1ru
6vUx0biBSC+NBxBVJZjND5bAMd+hQDBVnROoS6mvovS5SVOHOXt+D3Y0bxusw1FBfKbZPYDL1Gqn
1tiCgBszQDJa+Hw0WxGrxx3aa8Me7A0csr9/jFW0pc51cED7SY0Uk6g/Eu40n94hParg9AqoMGmT
tv27z4Y6/LIb14nzYT8/Zmh7ln63Uz6eJybvn1l1XsX104pI9T9lbjWzsaZG6YCxkSrF0TEZ5UNl
HJzjuF6SE/BGKFsFg5jbaHSAPRlBfrQNl+7l+uFqx+DJScefbSLqq73IMjgs47H2SVAED0qT5NwC
vS+L5MxrBw3MdRQ+VtiM69V2ug7wChqwGTX2pkaaXEw8rvXXTt6+OmlNRGgKn/pt5YSAAhWAcRHa
EOSsioHSOPEC7X2Fa1iEd4ETiRR+9V6NuSnYC1ZFqpWSF+2ANxMGvyHNDx+IN3K+2WtV4Aqt7hXk
VhB/PnOIsQbFWL5IlizHN6oyqLdsIWimgaUCg6NiUeN6K+NrVlBvddoGb5r4LZhI10ilKDPvvGn9
XjnoKDKmGVrz8ritZK2II27Gn3V7DywnWUSLg6/6uQbi9eysqouaJWQyHOGtRPawm78pAm2fd4F9
7VNA+bIG3X0bNbu778U4QIddz/zyMfKkJpxWzquFcc7v1Cmj7495vGmeek/Qnw0sZlgQugxHusAV
YfZzai2M2Fb1qEORbaaf2yF4Gqqms9WLbW0Pod8/sq7kSFQmjijf4xc9zaLStdMTdf5lGdSR1cm4
88j3M62LuwXdhrVDIG3G9vDPlAadNgFzWMzmeZMu7Nf335SxhExTe0aKBkt+eJ6uBtmkZjd6x3qm
0pPQ3OcnfhWRhHqGw4/EqiTjiQBdEOcDpmXvPNMoqVCe/feJCUJ/g+XynMlIyThklu4JIXBMYxNK
uwydEsJ59iZvQoORhgBEw3Yp7AbGmDB/ylYTunWRxGctsWZgMrUlZL3t0XQaT6c75goFfbCN6NT1
Y1Xdd4nJb2r2Vxfy+xa2I8WgXozDx3CQPRghGuZ2GnoJS4fiDtQwJVu3Hte7qu8KZrqy72LZfrn8
HkUy75mOLa2FGpD/QiGyKqZ7TnmQbubFxSqr5h9GoeVeXP5CPIrBXJWVoRMmUXkSojL4Rh4IWp38
xy6TKo152iwq2VvAjwAOaNcgHhBQdGzY/S6Aw3Y9G7wuwt9Sr8hcG0dmnx+cp8i6idYyBT5IMoV/
CpcuDL3Cd3P+fyFcWOP8matoSG5oLP8o5PcPN1DSDLEkyIi9zMQaHkuPWP44iVjjXOD6/3ZM3kvh
ipIN0nBntzAGc+FSnnQ6uqGHEeGUbYqTc3n0EQ+ViQbQaOgKAvJZ+KYyt2vdMezbzUQGx9zasz0p
au4Fr/X3L+0FypYxe1Fwq9AaL6yWrvqfSJ/Bu9P9oUwY2Ns2qt+GEKEWkx4YsTwfCxnFnqv7w14B
XxL00uQqvhxntzfJPPgpFNjx8LGSwBzDbcb7h58SobHLtN99OW90m7uowWUSa4iB6Ldm/mPXP4d8
gDv+qwnoaLQ5dexqDBvV187ja31KaHNqTXvz/djyC+TUuRF/bWJMd9v19ubQV70jOuty4jq5JQZ7
QbdVmltu35xN/cXe4NB69ETPgZGlxJd4w7CokQlq1+wRfubjl3QBQ52seHjGjKcw7HKupAGm+tUB
1nk2w0/CefCJyn/y34EkoCYjC4fV8K56nPtN+VKKGzUKs5SZ4NBDpCwOw5B4eht2tIul8+eInDtG
B7VAH3qWnrO19soNvt4KIYyZNSWi3pxCQa3WhW5fewZVIgNc9wMNm44nCz1Yl5t7OADbfD8En+ay
0j5SvWBoG9caJ1eKigww7R3tS3EYVcbLVViEbbMNKtG5TXQeHi3As8HSiw16P1SdPYUiDdKFxVX7
9+Klx/E5EL41Ta8ZaUpR1/XnStThHkTKQQwbbqg7l43Fbe1H/3HM09NIgaCngbqMqL4Y5tAWrzjd
aiGIGBVe1twqO621itA4s9b0ALVsKvvsY8XAafufEh/y0PV1TgGNDItrrLC6i+CnIZHKTXhuAU4c
R1dXejzvA4JKtPz0eA5MAyOS7WxZU5qgh10KX1nNhuglusOFgwzMIqI1x2fdEcNgdtv7GkNkvgMl
JtqvtvXE/zdQ8hNXBQEM4cfwh3yVKdje6HjnLAbkAnleem6GURLWC/zmAUmuJ8cgvaKtE7Uc0oGQ
kYgTA8IyNxn13cBLc71Tayt5FjyXLjZ76hpWnMruWnoEBz5qpJhDd3iZPEr3uzj0A0Bad0NkhmL3
RorS0WarFCi0n+47cVASSN8Uk1qECTk4fI+L/VVj3OhEFs8i9s/YL7BXSQGZ6htmjJEc/VxADSSc
qYHWkR/2uhAlEhT0nWVwqdXh8cfWidIKjf5P4+zW5RPt5j1AWAv2HYXIzrjtY5AaqgGPUo3kkvz3
1+neKqFaUs7MQGv6Z0xi0DqWEP8p8XpB+Cfg5cKcrI2CTHeCVLK3MB2Dzz8B7KnXGDaIqW8yvsZi
JESbDC6Q5ObA0sY6eROy9sze9EpDcSQEYrsjoXXGCAq9qRwa8BqEwRn5b5TwRZM6qoOy4ZPtP9gP
5bqtUe0ze0EmNvgsYtE8+0Sg4JIR4UYGyGxYk2BVH9kUuWURbHMh806QdvURH6Iyn7WV3BMDgOMS
qdUIcmkpyQLuk1qNHNxUIZ8dRT36LTt7xYu/3MDGx45riCge2Rla6B+4QsMJ70yRTXqmQCgZQygS
iSRN3MFOgCmpAJMEc6yrxpgXLs5mn9de4mHmAEO53zzA46Xi98vCtDUsN+nid50qIABmbaTFiTpo
dZThBnQKyaAu7lL/x1VTDvoaEa4nG3qm5ZzOOIT5iy2li+kzfI2bK0sLtuNUNYM47Cy9IpXjFJY3
t4lFw6glzItz1s0TYc7GnVmuR+5omqdjyHeR+E3LTeoqYAlLU5YuSmIU1URFOSy3tqLx6s1lWaMj
65cmnRaLqexjC1k8SqmZY+/vGzHpDc+jSyoc7QddcSMXoJcNpdA5GRaZCaBkaKVoMof/CKlfzVJe
w6Lynl/b1ZMsu5ZOOiQTjmVc1OT72futYETfCXrzNfjBLWfETZok9m0sguPISvT7V64OnCgzacUF
NjUAeQGT4BH5uQ7s7/hU6EF643UxdxlvSKKaKpMXqOBSsxZgMIMpEYKU5U0eCxxJUNgPyZEn69F3
/OuinfaMXEoaVixSQEVHjYUAHTXmcWuRoyFjpYz+U3dbHNQeIak85x57bQNjOLwazEL/YdC+oY+Y
MjK1e7lve0PIHHi/ekylp71WB4fR1HtPcwTzdcGbCPxQgbTN4YdwzCvsguiQHwnJ0DzFX6daDS7+
lgNyo4rtd0TOA0zX//JHo01213Lwsh+7OXB7gCMYH1Opwm1JigK5eWEcDzJA6YaJlzb/DSXnqDzt
wFoX6PFt94JaRKkQAm/2lSD+I1OWMbnh+lIEK45tXfOQqgxXCopgwbgyjLt0OnZUOUKIAw2h9myJ
SRNCGPHys4Fvi6vjNcP71lv4oMTfkQh3GyUOexiWxquIQBbRT0PLqBDQy5187C8g80AqcaAZBtwS
qsEedCaRwV0rOcycRvco++ru4tJvOZJPOrZZhgJIqZTMfS1v730swqNqm4ikVsnDlDCEQam5l+yb
avrsLG7ij/hksoIVFWLuDGWCHaFMmXL+UWtIR5t4yluN/ucyCUrTgiTvUWGbp/KWMJAyThCwy48i
dA2GdXLL1HHgdJkAIlFMlFxN/fi36qdc9seEj/zLMWg1Gc6DPH3Z9ttQp6b0C+/dMY7yMkg7LCgP
FY1PZxdIcahKos0qzAVlOgiEmXq2xXu03hooRy4086sFEhHVpKq5bp1NQvLpnmoVqp2uaxKvUMzk
tVDKp34CYJGZbxJP353baknpzp5ovOAcqWPaG4Q+IVmgdvZWbfi6wbZ3yXwMp9kv8mo69YQen5Xv
rFmx
`pragma protect end_protected
