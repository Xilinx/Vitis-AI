/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1082544)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2jKg85EiopJdNptgajIwKj8qQENVrSSQ5SzUCKN8+AP81qH3dBxNzuAH
u/9dy+7afGEGY14uWZW9FX00jKdmB8GRM8swqsnpiMiLlEqhgVCHrl4yZH6o1PHuQ9L3rViYd2dM
pzkj2GuBAPEjoKzDGMadHqJnXNEk5VSYwTQQSuHUDB44Gv6InkH3O5XOq+hVUKuP1evVuPpPLLwY
wj/8sqLv1Pecn/PzUey52uxNANvyU9NCZCEFXy/lg5OSYZ1iY1AjXM5ynGFAxlFEh15wVDwH2cXn
Xs0yVCGYnMvjKzS+J7QIc4ntHDSNteNxp9T8z2eRLkBpK1I1XaryPL66fO28pAgrS59mH2xrB3dv
5isvqIJBZHNuJE3vxV4apj086ErPke5NPMzsA2052lgjRq0sM5x10UeCzsz12vSaTDUNt/NuWo94
MDeX6Y2sOsVWDTclDkkVAGFK3m7zSJWIm+gY89pkiaEfTTdmTKY9OfIW5hlbZxDzObqj1K0Bs3NX
fTNAZcUh6SuKlGPas8nx+ThY4Lvyr9oCNjmj8+j5RSrNum3QHPrsWNRN2YURZk4FyjbobMbiGGR/
BiQTrnO+QK1Wb4EswbqMDhI/o7RutWLmFvxKwsGGxDCAXJUs7U9Iv6Owi31ycJ/FW0nyzv40zBfq
DS/Vp3cTEqbrHSeWXMdzEKGoL4r7gjf/f2qixVfcGCV7nHBni2e79LngVamtCzJegx10tqN2o02Y
4hNykNGUcZNmsM0+08gnJrSb7wDhtyxWhLJTwehHzZgleD9HPhA9kLAwGRojftbRbCFAeJjJYPT0
owC5BWB2lRi6WWvTYQBJrU3L/BzSQEhgWggx6ZhPrd+lqn69/naTy7XAnqU0RYYGJKQMSF9UCYsL
Ux+A/IUGC/QrNVmjdVK3FmdPep2/OQMW41J9+kMM22ncHME78560bnbdZFltqYBrnwGQv9U1q6cW
qDAkawT64fcs5GVV1swzJZAs91W0DCNjpiCSix7p5wxwh6gGUhU3o1p7FOGqYtjB29LQwCVmr4OM
ByGsdNj1XTekiB6Q78ELDBJ9OBirT7E+AnRZ2iMK2iUZ73zhBGwRAYHT0KKTTKdk/m6dVcek1Ckw
UnQzyDO/u5lkM6czN+lGTGOyYE5Pk6FxDYWhMfDkaj59U+RO/XERHDcD4MtBSMduwiTjIukQwnaR
mzpZCR7Q1VXLP/VoJ0okDICGFdXIRB9CAGlxm+LbmUiWpsJdQl10b8L72HoRNmy7r1VT/sGWv5kY
raH9tMRmI+iz2qNLpzOlcL9icUxYl9AUDoqtB9tFfx3zjEJYuTyyf9VykJ7wbs7ITmaSEnYlRo7Q
T0Z61XSO1/uENzZn3F7O60MIwe9Br+GMv9gfxL893zH33KRBWVJWuqtN6TLXsCespUFZ9y/7PK14
PTT5Lds755kUahsXSvf7EXAWijCx3O5swNyTExt3mukAUF+9JVxPSwzCJIEb9Pq2lILaE8gnory4
g00NGJLD/nbF89FTtycIN/fKWSIKhQh9uose49M8BIj7GkqDIVmrsq835FNkugC1Rtt3+k9OeWvE
7GeXoWP/zhTNL6LberR0m11Bca2y/pt/yqleIommz/Xp+VLlwdN3KShziDadqosN2WrJ45MHkJps
Q1ISeKL63WNm1klZ5mqCGcw4q8AuhehgbXqtSx1EgpnmzAHBR+gOlEpLDNc7wXzntVTi3dsoMxjT
ierD01ttmwxNe6Rhi1FTvGU0QTJaoDi3o372hOXb6CS57XFHA0cksCvE16bgpgklKx1oMdigeAGm
zSh320bpKkXTJfFyBznl9z49RqF1krTJ2xlrwTD+5D57UW1yA7wKI8MJqK0oFnMrF4/vrpYUW4O4
YUqQD1ckU9eJL5aqHKogceOowb8C5p/koTsbtjhDUCxLZ7yQjwn6vdUoxy65kCLUZNQbGOeK4mEj
cHj8pSidwKeQnygPB9VaivL85t1cJw1PCw9KYv+k7LjZ+uFuT6rAhvFUUrwjUud7ZuRjVuUN87KO
hINRLetv1hOqdvzXjMgMEbo9QcgfSk3Y/IE/MPJ4TF59I9TH4HvaqUZ8KD/ivmZd2vJDrJoQVeIA
3wlgYf9hS7suHi/6eTCQJufl4RY2H9oZz/eqRJ3GFlkNHqgwH7F3w9ucVFVaYvlky5V0yO2ogygp
iMXoz1Do/tkhk3LXMQbGHAFEGmzzX8J0x/YYJ1WfRv1HlqLWJN4hYnTkM1V5ysP1HJiGxUmCBi2Q
7vQvelX5utMkwQ2bD0z1L++Skutvd3oo9Sk7BB3zMWayz98q4t2PX8SyFOx0W7AjvXT84nfzqFS9
lXF0o7iQSTU8ICq+LwGQsWSeNEZlfsjk++YQTY0GQ3QS9BdFmrcg1A0RwLpP7K9WqKeFOaSV2RQ1
S+GnJun3OiKxYTPnV3/TrQ9X5IzFUEtwmM5BA6ESmMfmD1Qn+x0Kdoeca9sDgkD3XnzYvYleWk9e
K7bCBE5X6Qtj645MKcGB/07hPnj7sXm4Zxkf4Gp6maDY8uVMXsBAJSkmdUo0+ZCQAahLQm5Hh30r
vuZwLtHjkQB+unGjwUt+5AIQLK130kQ9H7vfzDM4PqoG+PU1cMws2e/FEnzHrwnLtU8HTAOPFrYg
D1fzn9XipRA09yOujtrM9QjX18jX80usnkj659wBzlmqe1tPPKs0yrrQJgvf0qAzb4cLkt0Lk7k6
y2RKG3t40eyC5G8V5iX8W4R5G2l0WrOZCsIbp+E6FYmLYacm3YjabKcUmbHhuR+IQhisToNrhmFU
85gjHTBpi3jZ80Q8rw8Eg1084sxCIaYFm0F6lPX+t/3EGfaliM0ATiqULqmjK0yv5NbxDyO7So87
+F82L6J9IQzeyK0bvftjzeiCPQJaQwlot8jRxTU0LoCc3edG/M+LUC3iFlkqDvcWWOMufOgmQoXM
qpPamSMVpbM/0NKbbgj9uyF4QAA73YcSHaRHyLxNtIBnIAJ4U1dHTxRJRGIlxLZ3NR5qCZwV4yAp
UoQLPKCe/c4IPbz/hJg4QEILZb4PFioUTmAUIwUu1pwQcFfWORhq79Tj62Ahm1ZpapcxNDeCO6xn
vsdnMqc5EK5t0g5I5jPqUgFENv+YU0a1/jRVrlb7cu53NS47X3v+GuZFJjs9IMxdKiezFRGcv1jK
7aevS4D3ZfuWOkabztaI7M66cKplcoJC4dmndJCpbWklPXS7gtjU7WvFdOdsaLkHf16SA3HSttNZ
8AjFXVSwjt0bp/EmnvqXM1ylki5jsUNs2UwQBTVk+JnjzrjiYZDvapDe78yE5sRlMV/Gf4Cdr7pi
+DzETnJgND7562tdIJqPBy1vdbGtReosz+WpwIalw3NAXmJ3baCED+MvG/M4O3AGnVgTz449W28P
Y0slxP44P70YcyAXq8umggYvnUg53UAbcGVBzqVjADJiFh+DCMWnt9zaHRaa35/na0BSYHfeCj3Y
Rb09+Qye1No60y4t8ef0RTwEgDPchhc9J6YsbCcPKxu2yruBxehL8q+v6vyV8Xr41Ukh+/DSNQ8D
LOxhA1J1b7ghrOvWW10Ze2XCIAFBOGVJoXR1bo7QLStPBuj8vP/uUINTnDcmGTaEVuk/xfMneHel
eIJvl1XV+ZRR04SEohWp7u/360+6vwNmylgtPIbaGFKJwAs6beAQJ1grLsmSxiDp8OVKUtJ9Yb1y
XtIdSuy28C1feHLk86Cz7FIhV2g8UkZnJbHbTsE3SNn1iI8z8eUo1Gjj8XbCFZrlOpfujvuqEuWG
gAnikEHulcDsfe2D2Fj3KtF45JUCb/75MxXfVDYMOqoTh5jZCScT+C+7KfQAtZJy9OTqKgATgUvp
17YzGE+Y8NTlLPJnlr1kDlPYVwtphf//WM9LWyHERwtRQyqnkhJP7+scye2Z5VM5ISFY9RbrUEiC
+1J/ctRLWWNAtntfmRqpg140S+NdxhDUDh2RNJ4k00/+DFZoih30jpKi/31gAQMLbA69KmDhrqJi
HOe4790qFpzLI7Ynaoko6Oenu5Z55YSN0jb3y88HNvqBZV7D5MUVZsjvZH9hli3ra55oh+IbvctX
DGbuhkPOaVJTIhEUp8o5loav/yI9T8hODyAs+TSfYmwQuP6yxyRLrZOxBriGd098am83KtKupWCU
eY1iOmAQhTUdo8vvBt7kzlAJBJCfaktVejUTKvRCMX9HnbgOA50I52jNFYohBP8vaSukX9/2Od/u
aDZAe7+uJ5TTUua5+vBSL0uMpk/YF+338WvluPCwxv2RoWlcRvdNJrjDCotuxiy4ni0AQGSbrol0
XS8rCaDW9C+5VLRPF4FEWyXwWevG6r9MvFF3O182Q8QvVtT67mA2+Pvu2uJexP/4njaj23pJxPSw
OCtJYSwuULgd8TDODTSd62X2mozyi34q/wMZ7M+5/28F/swqg35qU0vUKlv+0H7hLd3CHpAz8Eqm
ulSurjS/fgVrFNmDKUp0Uw15noFKoxG1m+ZohikPTkkWOkcDciPpdW0zarQKEiijWGIanTjC1Kdm
MsZGTADJ6kaAhsNOdtvZKRv90759ZrcU4ME6qLNz2s1zGRWqDsPCxiA3UDncEmGB485KII13dyUU
sRW4G2Yq3ZB3L8McSK70+hpsxD3zgbty4VuJpLoJuh7ksFLVGg9BKf77/ouCh+Q14S5XpG7tg9rJ
CriGsriMrnb64bpMo3azsKutCHb869tlml/D2UuxLDhfDuIzwUHTneei74v/bruCgt1IGgLfTyNo
7bx9SX9vPxJi2vhA60EljefnWCVFolfh31TenzlSKgV0Cu4DI3F2L9UF6tWQoA4AdQX2EjD+njYP
llh08nTKmwsXsV5Q/ji8XbpoH9QyggPu7YkFFL2HxMInPSjcgpJLInLcv6QPvPOQUoJnpb+JQdvV
lcAVaO+hU+oWgAzPFWUy9S0a9SszsweRSKGXh/li2aDIOaPlN1a5yl6JI323NRkC809wYkPnkfef
gnzkDPm4grP5wKyCnEKl490Bv9z6vhQVSLG2sEvuDT5ScpP9elB/ANu3Heo2mBXVGrV4J23fHWbP
pjZXTE6sh05Ian2ycqYu/EjVXtGRRem/ts7QekdSwHeG2YXJsQkmf6ZYtJgsmZbZbwWQLHdn/Qcu
Hm/hBaY+k1VseV8CB6DJAzF8LmEFVFr6SYLXoAiku9VMO7Fb9KS68NRT1HizyGXhr6Yr5I+8hmWS
w+a8EZXg8w8Ra9S0hxABXyUJa6zhmcjtFWT7xQkpIoeExNXssnXEtqNDQPLum1f2v/eoI/DQINPb
cz05r4zFBtdR1L3bC0ZnC9Gr9QCudGHgXlKC2lHyAZzVFCaEF7vCQhgxe1UnIzpWT+MmD5mKImlR
xdjSvMqmaXxDFPN/P7uuTmMSG4Ff7LJNmCGak6PW+25ZQHymNUCqIQ2oh37xc1pE4wLkNWu52CHG
wFrh8KAWSALr4MUNAprlH/E1qPbcXvu2WmSwnlHVXDCPnMDFq7+aqTcMIiDcKMaHpApLj+DVK/kd
EkmFk9zf1DYkKvebgpGHqBsDGDffbUh+BDiIXo5DoQ4FDkKpt0Uk3ckVMmYo8edfRtuIhLeEUGsO
UrrucuG51bZtZRYb8otSp2MncBubOgED6MEu8G/GxUumSEp/VNOG+QMZIYTiQLb7C1fV60vXpOvx
G4pfwk7miaSridyUcdTz87R0xQ3RchKuDYKgnXi4IQ4PrHStQoLosQC+v+fCACX2LXdJNjVwne7d
smLfUlgPKdYH/eU4OaJdibihEyx31DTryjXZAVV9vZ6TbrGsp9isrrCVD/nKnG4amvAICqR5jLDx
nax5aEIg7Uu6cvVxMd7vO5RXy5rdmNXEVVf2zQT+7U1fAkgWsMPnVkW4lwDDK4S4G1GNpsbzr2ab
dx9mrbqciXagqojZ2S74oLDMVzWWU4yWaVTHXv6jv7j00N0/EbtvhbHVHObu1JCss9MDh3MKdlTd
XsIf8EUS+dp5mmYcA6+VWjR4L2zP5Nb41PPvXFRgb/rYv7uqqItOMqk2KY7DNOL8+gLr+3BpO5TL
9/3BZS/uadFK5EwqSC/q5/q7vqhZpEF5TJzDPCAOZdY7Jp6JxulCL5MHJ7TFGTfLLkq4PntLgSGn
5KtNnrQbndHT/lMeJeCbe8kmt+C9G2JgvSTqjm4jjlx8r8S8r4I76TIeyj3tRBOP6dwm8UisOMt0
hMIZ9cHOz482BEMX8Tcuuw5LAnlko8SFeZPbgU71JQxGPqNnRL32qaPC89XkbR4qzjW13zA95nIT
crIvaGqlCykBweuy5o9JBeVuV1FW7d/k9v9zmxZ2vm6LiKw1enOB+8zSadx1lYy/zQutoF4IlCjA
AlMLgddN21Llu0wTO9+E2zmOssq2TshHxmQhyrHgstRkRtGjTWr4I7834QjkSrJtCEg3iaA6VlP4
c9zatRyGlqdfcAo8AGH4ycUCirmzqsdxKNNRXbVPQiEZbYg8O0EmJIHSU4Bd1qmnKJRMAtkQ+hyG
7tRq1kGF+LgqWsGvtvgOt5zrXVqqR9vzJ5/RiD9aOErNWdm+dULjGFtBA3KpjON3na6aqO31x4v2
48tjIph8oNAWTMYnPbivLbBu7DdxTF8/ktzUkpbAwogPERy62zySMutmoxu2ZkrLLfJZCHmASCdW
4nID4mPtkFwWJvoTDqfAvUYIO/izKKLhfSERMgKqa2+mebh0hoZGsBIEGvB59GX67KR4bk/x22WU
EpHWrCaONHyGra//NCNxaHEsIpdDxX/uYRBgOtARGVO1qWdzSRO16Z9EphSZXYyXsHOG+8MRS2Ob
0BDI4GWIs59iV87PPjPnoB7nJJ3oJCnRNmXITp0xHZ0RfbqgTH5M2UWaAME1uRnhSB/alR7kMW01
AqCnmo6zAKaSsm1cLyhuOrlGmtznuyv3k4NeBpurcai0/MqK9DYMyxIaBijHsUlFNW0EXmAbY/Xo
KzSziq0mheOUZwK/Taeaxj0a1TiuWrVAhvZh1VQYZdJfTZkomQ/R+mY7HhAHDUgjTTV5618FAj9K
VqNFYKYMTVAb37hYzRi8Te7sCaW8ZhpS/VUQ8tL1THb/+DVJJDeo84vaWQ7dS9AQ8DyYeJ2tiiIk
Y927Tq3hmEYrBKRGy6O2S3e4Uz/WSXeKYjEdP+AeqZay5aOy7/6S/QIiG6z2qf4Ek7loGl8oty5T
ZYuw0leqCm5tggl5QB6iNlOlqXj8U+0C5yvSk+1BmBfHR0B1NW2cSfjrlEz9uOZKtXCJLwuNYohs
NGPzz+JFrbKnk87gppvy/T1VT29QGQ9O2lQiGvA4C62zVWP2HJXsW5SUYTsl5r1vQVAX4EyFn1W4
vY+Ykw3M+G3j4fgQ1mQhJI2WyfY/FvBOI2LEPEO4fuKjYCwivHZVE/FBSxlwtOpmLLQ+n/+E+ybJ
Rnwj7s5lOhtybV7EWhg1BjqKvInxIpZSC5eFBoRedTqAsrS/d37hAocSabZFi1JTRmJZvD/wuNB6
ZEE3cbkZ4iQlsYj5Xp+nUZJ4p7onV5uCT5WXN6hzmjfSBPd4PWQeHrXA66QDxKAhHlIbIUv9NBhR
FZyHM7GVNY5U05dHv96FsuOa3AMrZTswv3OEIOEXm6GaOcmQ2dr387fk8toZv1+7ZuYsEzFatJp8
ScmrxGPyP6XE/qnKnplrXPWtBW/fbQ8iAQanF1drnJ6ghs2qRe3XSoj9/VFJh3LUA/CgcPfZLbCv
Vbj4nOGDRPO+A70TJefXoFnrTc4epQNGheM+8q8WBQ6y7mRFjzxzl0NaErbndVYBCnQSL32+1Jvr
3H3qlIfYOHr7lMg327J52ujSOy8k0X6fsHXM6rNTa8499hP5mArb0RZwCR8Hl9b7iCgvYLjX6iYd
se6KOpu4WLLJWM63lyPcJWLKFBUWzvJjseAjan3D7Hbb64QJngIh+ftxupcu7zeIzxi5di71ZUdB
Hi+SlLfj2KR+0ZweimuQU7mzurtQA+p7lN3PaVR3+GcfZPqSpCMjKF8Tx0Xj3+C19IGpeOcNEXnG
icjdPks6mNT0QG+EBBd6+Ezd8e23eYDyJVpB2Q/RiH6dHQ5AOSMY3zQLvEpp3ARVUC9RfjK+U9YM
twlggAOW+F8JSKmzMHdORmSsL8vUNX/VNJa4wG9S5X4FH7WCiGHP/kHeouCvg4U6+hdQfnVVzI9B
JMrjq1+7CNggl4R71tW8MFk6n4h5UhG2bNZFHy1do2jOPiqHIrMxF8F4JpPhniNIlg8B3wY4pEOd
Zpd70uagUFwewlBXWsgibYP1D6HuANi6VOeUKTFchr410DFDPk0n6SOUWtUL+HmmQkSco4Hz4G4R
l1ABVJ+pxbfvnpudwvqZo4lWAmSBMKKD5geRNi4EGk+nwKeaNP5flXpRPXqH+S9eMr4RURGNktuJ
o4g5A3s5cVdvhh5GL5BybPNlBDyPIZzhcpVYZ1FzFcROul8hgkdwqxJ9YKFKdCf0Us5YyWmscRwt
1I9y9Og46wmxffU5VbnSy61O63mnWG9ZLmIWBak3AbBtET7HYsDLTohc5UgIwuo/TXK9xfXCjhj4
AkRjkzNgQm/HXs9d+0OE+WdfHejCsBM9X9kMCJEG7mMbSWGRPSFZm+X/ghrW3wS/b7z0Sp+HuMH/
FJ+4XRv6cHXuql3SXlMv9+keMmb8oAS5cHkLKVAohP5hF5qjFxyqehjIu4skcmajtr6iZSWo4m0x
7MURgyXmWGWyFYfyiBlwyGn2yC8Re+QG1Tc7SK72jGTRxjIrTGt5sVGGrP46oZP8qt38nJYkYMD4
oodejJdBqjr2dawnMVKcVGH8EgDSXh0ibvUPLcxcICQXMv9YtupI7EbZM0Ic3oIJnzf8lixm3X3f
ZSORs/c420CwNK3KSxwlJS7W7jYxDX3JlmhLZoQKoGd5dRkdrkIK2EK24LXqPu11vzfrkwki+SY1
33/87MVINAtYkMoNaNqBcKJfxtA5zdbqkxUbnnaR8BvhgfXr1HQ5BakkXxFp2n0B/C4Y7HE34oCG
NskLrvNCaOMfQX+ykILezR/JiaqFD7GhCOhAA2en/D/AGPQ9TTGwJBdBEtT2U7jb2+S4Nju9LJU2
F0o3h2tDcJWywV+dpZuzQYOj9MpRZCZXY0XHKeFUPJGGXYY0HisEWlWSGLcRbsKUsM2hsytyokDO
0atmoQh+rCzrLG2StEdaeRzagsJkwzOE0RfSsxrLiSlrkc5EUPkS/k9q1nSvays9N8eBhbf1iA7x
IcaQBLukj7ReBD/RHa3R0wIeJ85bN9mS+q1Jigs4PD0K3mddEMo1dJYvIhEHFF3XmQHBUaPBRUJq
fp/uzw/JICAuHwCdqQb7cWjIgxBHxyKgHvHwAIzPpHspcBHHN7O/mZMgRq1z5rUquybwQ7N4FQ6Y
igAnHtZbVbTxvPGU37DB16Y4DmUCvPbo0EAIuqLD2SIGSqDU0c6tU7LnFdlNOoxSIKViqxsb99za
RBhR30lEt5+cdAZU3mOemodvnmLLoEguaV/DRqT+lMhbuMQfKDS7zkpjW2Soposq3zoH6KOAA6oz
AnFPNZvZM5MNZ1VDyJlKyETkol5X9RzLpBIlRNul0oNc4jBqvRkQajD/pu/DOikMPLSgX4XlNVXP
bVQXGWrMcxuT+ey67pvsSZpRvx+jTee/G9IBzKYMMNvrw8HDvlI/0TGOdKf/oZfThx8NcQLIf2II
veG9mAFW1oHWrVPnDpGLqnqMKwaACmQ6W6kq2wyuzB4/mdd8litMjT+FzUvNVEDJhRLW3E8/jFob
cmSBaz++h4NUynwp9uY93Kk/8w4XcgkjTTPQL50MYKHS6JswvL/AZdMgP9mNOTfUNdURElqYDWBB
Np5Du3u5IxPYTC9jjWp/AWb9wJL6RKEaSUgaXa1vB4uXr2jK3xh8JswUG2Y7TdcsrathFsNF3XF9
qKdcetI+wMN4WFc/dUFdYEOfdKzWHvSYVKn1Fb5y8CBL/NRehJwaJOzQZCUnJg0nkN4IqWqnYRFw
kHTYGz5ABCoMwiVeuonZQpDlG0hQU6mhuZo72MikYYZTDyASm6vro7NykYltlYX1oMSHh4nwE+eI
nyun0wjE1eRZbGMYNNbzhlPCAmDhhq4k7fJazf3wRELbykSwrz3XHdcrn4+xM0U+sGMQOCMCLvH+
jntESd0qOxpBukniGFILVtbLU+qzYwpMME01pcV079WQxt19bl4awP5VazA165eWNwz1+l04yvWN
3fa+5kLIV5vSWgCLdl/SvNqhUZDgExaTNzh0/OgShp23/PuvUKXo2zgDI83CGwUiD+PDKcY4ggZ7
qz78OCPRJdTVKlGG48abMCR1wqcxl21cdGpgS70JU7d8Riq/zzaloIdKdT67mYCgVF4IT9IE/xQC
+ZiW4IgNAnlGBzMr6sxFsF/jcVeE2oilP7uc0SWrjxpNviMFxGRPHxrRN3MXE41u6kk+5I8YRq2l
WSZqnvpEkg2hXqQnUkLVi9SyQmOHVmDGxJmzsTso3KgIW5cV0mDrWPkoYutBcblAAwvYehHUo3QW
OF7AFskPVA/Nsb0IYV0APXkXG9yKyc4g/5sLoq1AY7z81bmmsQFodsVmH3XUiezeUBdtgBmq20//
Nb6TMvvLAJseNdf8DjIlGaHTKO0xW0k7YfCU6UZQkkBSxwim2P/rcg3ThO1DqmMZf7mVTDsXzwCg
q/02Zk3QYi8DCVP9qLNqxJ/IBaJy9wIy53e35RL80Y3tTznOHAZmFt66LgMDtV5g0SPM1Py0LiBp
PkooTJhQjrqrvp8rYPkD8rlwI55kUCiztoEsUhC7ecJb3l1TC6EVOnFHZSK79kP3FndLEi99AIfM
wE81L3mTztvakNXsAGWzVbGp/CGKRjt+DWKSrCEMOvuJqKnmhRBPPnV6ZXgh3FJQydmw9DAUK7qs
HTI/8LSkg8E1j1Ggo0bugsYETqWih2XdSYccuxnV9s1mnTleDPrVDJ0hKZZQ+7H0v853MVeJVEiT
52iLGnxRT5/XHqbwufykjZl/2VE2lyChWSkO7aamavRqrpa7Orxh8OafAtN0Ghtkvg3lYDOxFDX5
e96veKRfsYrObOhgKspaJan3lxhNyHA8bGFuIYqR/XbUFWkn94ma3PXAirDpUQWnrlFe5ZW7ac3U
CSgi+wOPbQC9V85McclGx7mkNmiomlaYprbBly/dc8piGQhX0cOeUgGoH/DPlCMYE5aab8NxgZyh
DwI4yI4+xjyRMXuIEf2h6hayWPmiMVrJsTgZ3HU1VhqSWOK8Ccc9iOA79lClIa8/VjHQQ7P8lZEU
5Nli/j8NAefrq36QGZn9wnscJSRsfsg+3OU40tzVohzJRl9INFAWpCxcdbRwQSRrZnqspFiqHZTh
EzceQJQMKuwIVqI7HD4+MT+7MkNHqelWvP1VICtRvW35Un91RywyrVcUljNg4TLaZUmUQMavun6E
/z/MqhIZLaEz0WlNsmc64ywV6YzFDUeMyrDxD69gYtWn3bBTuh9lpRzzdMidG8kyYiUtKm/owC6e
FlSFPxfHiUhOb5H6jgYJ79madHoR9cBX4mQ/LG3Png6wdffN3aGTjIPMfZ/NUBfWDIJRAYn73ugr
NnlPgXaiblrENTWBqnTyYpUVr69oP+yx4dW98J8Aiab9Ia2Q67nQlJ+MDS2da1gDYLQeDS2xDnqd
6563ZD+8ENnn8TzenShzFIvsdm/bEOuaySVgmOFjUqCtwIxazrj4PGl92BiHO7cewA9ffxwq3QGU
B+olSe6/PicyyCJMlHttso91XIW+430ZIVa/puE/8eBkoXsqNVQz4c9JHOtn3Hf3BliXtSkuJdAZ
TdscChKt5IIx7EDCCPdycyXYbAnv4R65q4qQsndfxaXlvCadMNNBDb1ARBuOk29vv6v11gFAW1Yy
CcpAeaDVJ+eqhcP8eAUdYyEPoc0R0qw2BI2APUXtwjyvvackW1zKLtBwBTmM4rc7o7rgN/jbHDnG
R8/Dv8Z06XWC2+Gws+J2TZMwZR6Rw7eBYEqC1EpOhrxNMdHRlaEIeu9An5wi0Ow4eFDP0OfU95zP
nNQAYJ9B5uA9PnxOAnG445hjp5Y8iuPMCIJ2HEFtNIK19z3+FMx4zHWmVAVtKBAlZEClTqKJYSi4
nVZQbMvCwkIDhRVITBQxSn/elde5QOJH/ATcyRnfsFoUUJ50XvnD+XHitBIfFPyz/OkjGTSS6NWo
Y8Jjg+t9FEbEdDsv+vRGKBw9ZOl5gZVzBEd0EvcEOYt0tazTJSKHpe46MEHxtuOEH0F3fzjDqqU0
YnKiplHryQvi4+O6sJp471GSo2T64aFO9oxMml1D+Ipe+NIecX+hkY0Gf/QHS8ocgCZY3wGJPNa4
IwomGSnGa2dVQ279R4VuRgMXVgA3b76clCOW7CSqR3srApnBdBR01JbEeBHPhgQb6YVM2KyMq3/c
fwwX3tRMqk3aa79Sy2vIpGYUvPJDZ54c30zsoO363wemrcwPMuCfBaehq3AzXa2+4h+heNS5vZK5
FJ2wGiKLEiLpy5DDfOaHeUojJFQYM0ciqIXKpRvSccOY0YwoZcN1q2SN9cCdwC54mXSOD9p8ypO8
pojwGj6z3P4oFWuZZkTMUiQkSFr5hV+UXxNh5BHB2z5IcymRP5LnsYaJ4VPwvtFJJJb7zMEpwRfw
9dDybaX6Cu5mwBPHKmOHR0juEatFzp05cumv7hVM9xuzxTbb4FxMBbDn2oMZrT94SEBczo7TzO8l
YLU9msPXwqYHAWzjZjnEdeU2ms0u9mdEf+q0lDmzN2Y7HMrlAf8KUKEdJKgleLeGlQHqpGIRdJMa
VfvchmdUQ9aX2b+JjSaWvZa1UxtJXz9DIbCKNzlomOL7xRSh+c9yrvgZM3gUj+wGwPkW0JutT26S
R9QLxTW+/ep1WyAj8eaooz/G1uNOaJtNwCrgKwfQvA70eFZMr0JGbXT0om/HAoRlyPgIz6hDMk/6
krtnplloKeZcZ3Cw86qhkUqpG+FZPg5w2nD9lURMmUhMbWrapijTQz3S9IgtH4dhHD6DXANWjpyB
/J9y5IR75nsNC9T/1Rjhn5J3Ev58WaP7gcxfY+uS7kfJ/l3Ies+1fkHx4T6CCqSdtY6lxD4doTLz
0yev8w8dvniTsUtb1J/3B/KLRP59qwAzmS6M/qr0tAjjJtQuTrD+7NhQO1X7T0218Y5XrqzRg5ip
j1NVbNnBxf7UMqFbEN4YPAIdZBIkKM1drZ1Yk6HmuId/tB7JiEWTCCYXe791MBy2GfAdyA43rTLr
VCcFq8kEllgLczSO/3jL621oUKHkf0bBILdzg2NYFN8o80rIqF4oda0330Tx1TA4AEsXqPuSBJNS
UctQN0DHeA7FqwE1JsYQFGHGKKSnXgqNkVvVmTozOE9AusEU0cUUobHgjVDorfqq8FjFPOG/3Ii6
qPLyHqDQe7oFVxZNwO4D2g1p5hRA+zyCOF+0bd0Ndj8qAYxTRI2cvRB8Tw3lhDKAOpyqd6dE+Npt
rNsnlVZ+pqJJZlg8dZAQ0HN51zYQaVY9Azdp47njt0MAiWLCY5zo35xtOqfGvSbKt5kn3wjRNG9C
aot+IPv4+TTNCcYhvH3DLb0fNg8o0TcWZiEtuTvomSxDjKdl58gM0RGcA99yKla3rHnKEN/AmOBp
Vu4ot5N5pWFuLtbeyyMCBaIbYrsPsHUYH4rK/7prFCTCxMZS8B+mcunye9dE1d2jnc6pE05lfIjG
gt4X38tDA97+7CWxK3GB54LPH8OCqJKB1ZPFYl4+QT++3xvZpVQzBwDObZLp4c/TNB8NgpqsVMoc
LKsiDca/yvVA69znZNJuYSuensldqKnGeEVMbP6fShQ5GxgNADvxaKTgZU3XM09wEQoenzogc6Zc
m3Hb7WLOfXD7EZcVdc2VDzv41qnIokiFSv45KBxVrlQc6jg/R1/EliYmZspWsvNds3DY2qmc8e2D
/rjavpFoJa4z4afSvSST+dyInVArr5mmamM8iKi+tMonYTbIXqwYZcOCJrZMRJq/XJ8Nx9Zmo1Yw
sn46OiOK6bxn3x5f/mntbXwZ56rCGijtUs1JfV+7fQqvvICJSXEk4fFV/trUFpAaAntloxaL8ife
QgUY1lUeHW7ThV4DjMM8niy5olIaCrvlQsC7RsKKI4wv1WnxDONRkzrRWQqOCyTFetYVbFLYG/qv
O+TjGHRiQRkAmjVvu3KfgI6JQomKY8KnJFVJgs7UDyuHAw150/64xp/j9DAsiOj0bcC+Syjn+Fnn
yCNYg5pLBfOl/GJqUrUTCDU0d/M70+GrMIXHxP1spfhsWJemWLWuKbVcBSr86dMvWwBraMNC1P4E
khqfT3Wut2/hHiEUMIE14jr4o+TaYrWCbVIx9hBNRGCJiRqrzrQ+vOeQXB2TQDfNniquViQ5xKIt
RoEhsTzT1gnEFOU3iP3+2d/JpVkrdRqLO0NgAWWUJmTSLABjFZthIYLf0onL7wQ6Mb/mP+6A+JX4
hKMXmjvvRJn1Jt5zU9vynZbbJmG6yeTPoZZv0yV5r/A5xrVaiQXT9OfBeuiH7tb05KZgzJg6W1dG
I4kDeEMb/Jap0kIV3zuFI+vISsEZ42qt0I8QK+Q7k31WPdOkd0z48ZUopCyPsyshJ2o2v5MQPP2d
NLvavsaoYzgnFkLLDyC+lCTwXVaQjpoGu44fi9FikN4TKFbYe2SeAC/THU6QQqL5nBe6/Ep1aXZi
H6mOYvcL8k4XQDocu6Ajw6RPOy0hvQa3crb6trbFhddVqtuvNGh2QLOE1MkAwWtGlq5OY3uDWsV7
uNMJPHYM0bTw/h04Isa9HWLq759Sfh92/wG0dngBPjGYP0+QQOAvVmNSIA/q5u9BUaUIlNl9xJwj
HWMNEz49U8lZz7xHaofOmuh649UiSHl8ehNgxQ5Xec7QTc2a6yWtLe4tPNzubavXjsrW3zOzxfCC
erd3xmERDL3l/gfcIPpxS0/Ho3zfQMpAuMz80HLlPeP1RbED6NkZFNi3N5zTrs/0VCD+7h5/Rsd3
Du23+y68+AbmNlckK1QoYRvAqhb2cIJp1xbBXkuw7aurMZLBpPricLT0BvGl6TrSxqg5I7jx+onO
knvY/jVGd9D11qny2Wnrlv5mmzzvAWyDzT4r7ugkiQxQOZyuG6R2vBilBKcHdHezigcGNRsXL+Tt
LKmi0Wo5oVEbgcRpj2oYoCHS5K0x/8qhCf9E6p1ksaUn9UaEjtJZUJquWj0LQ7JNaWkps2Fr76xc
IiUUDYGqhy7/pPJEZFAcog12b/yfKqa4613BNRDnmofZxdcmECNE8yvEzOoudS1zIup47MLpXNlF
Q2L/rSca/axhLxYWyMZZaX1uHninheJBWnkacbVk9XoWdBxnniX29TGO07A3AS9wkR9V0VkDUBaB
Xh73ZUv1SiarQDjI3v28mPpKtq6EKFheWZKX8EMCVK7cSa9CtRSpnTEGleQP4TOjvAR4xPUnVbJz
NN6obN2eszRmRieorXN9iGYoG5OWI945XSK6wXth6xTSl3UneUfnEcxGIlgT8Y3O3vRt2+nn/yQ+
FIkgvyBVMNpw2OrazOvjc/g2BjxP6gRnSOZsK4AL6aP9Q1w1lTmMRci3CzzQRVorz5F6Cblah470
l1jtiZ0FgpB9ghLAe0l/ifSvGZRnfWgYm3gTCLADkwjuynbmprDB6yzT9LWXnsG9U3uvdGrQSlwN
uYfITccOx0DUlpT4RTdBI6z6csh6Gl5AiWWKTD+IvNuUxWPsEYHoYtCBzNIJN2kmdk8itqIHnPpp
QfA3XnUUaB+OUFJwU+choepHXTJpmUTZTWbuWdToHR0JFmF5ZRsxZBiYMTl+2RGmf3t0GlJyOylK
EQUNRhkiY3aJvBYqzJRIWebzmxiW4c5+yT1iI49YS8kO4LpdSMRngFJXifEv1Zm3hMx5/1uxFfvA
Y0FqCbvjxeizEe2spbbvfClJ/YHgAK/k2lmzOQ0N/IYpg6ojwEdxUNmmPTXyLJVhmFtyUadSttlW
LjOYkO41coHpByVoEHoAL539ACcUflQlwZf/nh8l1JaBeRoIcilg1b2ZYmij93QVC6AqMp23oa4e
AYPCUeZZopWCEH77nCzKLGCKr774tE1WpLgRCANeMprdLhSgIjwKZVK7Syx+90fQFmv1r5vtJYZr
bRZBjTapy0YIx0oi4JHAsgMtEgziOG3ZUo1mINpiz/EQdlitRgULqoH/HV0+B2KPlfAx5wfv5Fz8
WrDECczQPxKSXNj8tTteVuBpjf9N1weDclnF/FalcO//QEg++wdFOZzjTA9TXliTeRPjc6z1cndk
5f17CySYn/Fxh++2wDwG9+ZaYrfG7Nu9fhzgoXgbNHPQxjTMGWi7flmrbm+MDEpjuUO9IBZm6lFN
PrcrK9aHvw3MQHH6H2KcgrLQJOkP51ZVBmvD5r/CUZJuBsFQ7KEFw4sK01iADco5qoXrITe/g35B
lRYRB8dUICp6F/Kx4FXbkQJ9D7ThejIuTsWMho96uqxpyO3zqOWljWvmNn3+5JcKA/VNJAbj6qJO
QsWYFPQctTklrfNxifp2rMU21eCyWWKXfcKq0ZLFfR7E4nCjLUTBY4dMH9UJsLLHxwYmN3P71ZCX
O5Dp4QVSkHQ4WLDlhO7PPYQWcAxFaH7N2KUhqHIQ2qpRjUBQXRzf8H7zHav1tHdQFhUmdThYUuEY
nkYyCWRvUpon7nBIvzU/Z+AGrKmZIQRjaytiE27mCjYgqIIQxePRW1x3BgLbSRrIYd34bJcNon6e
XWVzvP7IZCumDAoypUOwxO9IzDIarOxEFItrgOM1EeVInZcl75BoZZwYjpZYsUy33m6ojcMLqEsd
kZxwNAVb/4apEE7evb05fk58rigUN6kgbaIb9QZ10QCe+V/UsRktpUdZhzDdBc1NAuS1Y/ddtN/S
Rp83Y2EsmU4MqV4BV8NU7fOWL2fWpeckTgnVzCRSIUoFeDDqAHycBYanVgWbYd3e4MNOJw+jAKr/
4z5lbuOGUMKgEfUTfqYCek43TBwharvrmgkGgpV6WBnqLq6iN8E+KDkyD+NBRuH85db1jklI7H3Z
C/+Ip+XQTPFGr7vl7Dkhu19i9EbDsOFG30vh8LyvGpP9SZSOUp9A97k1ExoGeLhFqfmZhndojrlh
X3mdI/rC8m1DXqVD/R6bJdT9sLQ78JHlH2kR7MKcpt0X7U/YluQi8LiHJW0J2KPhJjY1wQS1kdBP
bzZ+at51bHtrNk0T9ztD+mL423UBrUdtrzjet0yMaxZyOSHhFRCNwUq1tvGJEck+tyLT6noZJwB5
Q0d8mgmC7L+1vBC1QRKE1J7/xI90Ey/TbkoK1VcqDoV1tv/WQd0UaXXZoqQold6drMkHDpPN2OQx
xvdIidsrKutRenUOGIHjXWBxqW4paj6nQpWGBnqQiSqC8w25Mds2pdsyJCavHUgdOTEwv4yzkzQs
T2DQqKpLL0k8Zmp0UvWyrO0MxM5C7FDpHM3/19rF0L1K0ZWOlcE4x5u7TY6iAMN8GAdOetiyIMf9
WIsa8XOBzN6o7o26M7gaGlUgx/UNwZ3D4+pJKNoFwUilfks7vmI8Q2vaP3IEN/Fca+akeAfoBruL
LCp4qL3XrhddbGlTUh7AaDzr2pRI8wesutZiMKAP2175NL+3Ay//eLrzOcYX6APpdOywEoT2HVTr
afyEAXJGqUyt71GwJSAYOxYiM6rqb+qRPxJtlAakukmFyySX7FkQe/F6sYoGZjL4BrDTWDCWbT2j
c3Yc84oo+sssM8orDPxizbixmkosyzPLZ0ZVTbCPUZZSN9ERzaSc1GS83lz122/Bl8S5/4CMAdcv
7+1gbpKCfvj6YQnCamqbn6oKyetHC8pBPrGwSqOPkLf0csQOVs9qIncFNrB/4cKa6siRwVe9OfFm
soizNugR1bIjL7BQlcMNKyRahQOXqmaGqPV7oj6lrADaEsdl2cgCXnd1GCRVm0hOM31p/depGPXu
xOfoCquctSWjsvdeumghmUUBBPWZffdScHcRIlL7FnsbCiLwg9g9yh+DJtj+DQ4XIxB/HZY/ma2E
e/flx4qIIP7oLDJsyI/+uTFEF/mW2iU8HtxXvjVKw8ufAjDfnrQKVxk0wb6tjQ+kqBWu/WXQlk37
LSlA6+lrbI56rQGhpuXR8S1zCT+t+RBBYmPQ7xm8PcZ1vGZ/DpTP715LJV1s3WgjTl6lqnby/KOG
0YITokNkEZ0dyCjnfljSSgmchIaPXFqOc2AQEI5+7RZFtkPmwhMFxaryllmLl/ndM1rzAMimFVdv
wjGVFMW3C8Via7EOW0MRdRXsWGslwAQlMnlh3eCKPYWcaiIgfFGLfd1DaarUHPvQ/vmLIcsJSg2n
7UL6QSO7+ot2siAJ04AFmsMKJVkeaeCvtjwYyxSATFnpt1EroWW7pgQVPI0N0ZRy6gBKVx7yyQB4
205cIC8QN9N3tK/nvQgjAvzRmCrgwdVAWH9IG203FUsag7ZG+xq3lfaVeRWX1Y/qZp1HXJkSlvQc
Ic7A6hHRaneT54jfQn9tiQfj6v7hIhIz22+C/p5MpcQ1KTmykrFEQiPBSY1C14k7H3dQYlQvIqzq
Jjidt4l/QLLPDKchNLJgVhX0Dh6VVI0GWz2xaSov7K8KRKGpFGxcFJ8RH1kjzXUTd7LL4XNpKB4A
5o7bzci+2lPlDvoHklXQldkQEYVkKS3gOZKkVJkzVhn0KjmgPeQVRDK/lRc8nkKHAPYIC8A7qfC4
6u69q9hs8zC9tuFh+dRNpN51JpJg8s7eVbf4lCrn8TlUYFew6BEPQJxHKF/pswCIabY9OJhH+hVN
eZOHx9artvT/W5hvQhX0Um/YntMEWfmSvUBK59KepTrHyVJs4XoX900rKKbsgRcolOU1cMkuUX+Q
+qgDKy/SzgowjUoHyRZ0n3Q+BdFF1qhQ4MhsNvbUCaYNIpSS5zlewxX9xeFN78NHpjmPg3Os3szE
uStltZzCCVz9dXm4cCQe8Ko9zc/Ryd97yMSHddEVnkaqGJpjwbVPSK5B0Nq8l0wQC/867NhQeJuJ
tzFmCFQrNTLBJuUrEt5VD4axtFacrsMAXhM2aRLeqKvjdBNGa9bwTUVQgqffANsmYwF6U5ooJjpA
GzSWRvM2+EXbaxUnKp7qnjjfIK1c6Fhnf78Q0tWDVO/Z4kA3AWZzwpzyWL3/aDhRD5omap0C4sMk
/XOqbLgCH4qjtOw0mptmtmJRPZIHtth1kcL/RbFkT0Y2zAD2fMiWJoOAcJTo9NAzpqTFkqTirytG
RM4d/KyM7OCkWGOP/CGwgzyhstLBhcrOBKtihu08xGTLckijZLQJ3pTeSGTGiiezQ7Z66tDc4IR7
aSoC4lz1wmTOUPxRjwVmoVj1pVYUs7f7rL3H+k4XVMp8DHUumOJkAu1e5D8tuo2/bvuLq8NfsoK6
nrLd2dAKTfPsrL3LQLJ2Lpv6QEvSYOEG/CUVdGxnGeZVGMWB0i0RKG27/Erb5YOnSRWA7HIsQAGn
O5q2J4GtFe5CIbKrGIAQp1NebOp+pr9FpIS+/h5S2OC2CcMgh7uW4+PDDUAgA8phpiaM9YNniS3i
bETcdGtZFO74btVWYpb9AADM/Jfs9Es23+jmyrPUGByMcDb4EA+d+UehoCNFqAf1EUt2Ai3Rvw+m
IcMuh/1T2U3XhlgRxnaXu8bMFdzYdjD0yv2pnxDIaU3L5W3G74eaK9Q5t8bjtBX4k2yIh3KAACu7
pq1HgBnso/ZRxzzeQVutqYJpnp8STCf+SjTCjTjVq1S1Nw6WreSBB3f/Y0xfkzSRspadO8jEcJ+B
VSSjHq1JH/jeSvsUvVmPn3CgGNVuZoFLZk5jfsFFisweGJQ/SmFcLhbShrQkNWskJYI7C2dR7tFw
eMRZE9yXpMSe9pESv7OJQysS9zZhXZECwoXnNW4omho9cKPvR3DUaUPG4aXynJ1FDqzKjjlXOSiy
41htw73dT2bTHxSV7r0QWm0mW5/ncN32ojyH0kjzqXJDV1pJvSvbnVSlzQpbcn69UrqV4e8BfYHF
yGqWyhFh9yZQQ3b0DjMDx8EFe5uMDZlLExhdD5LQzeozJQlTkKxzjDmOLF3op99rdvYamD+Ehq0h
JROlwp/Tl5/SE434J326/eJeTpHqFaGyS5EmcLEuFR0sIcDUgrPy261t+GaAm7gEYkIZ7NBvI74p
ViEoie8GWbiTKtH+IPatBog6WUeefdmOnxyncddeKRfODmrB642yIpkBDVtiqM0JnPdLS3aW+2Cw
xXrSxW9/GWY9igN8nnaC0C+qLYiSh4i1lW82bMRu3ID4hfCw7c3Z6LCWsS71BO+4i4MAGBXTBTtq
n8m5/hZvHlkg2896JnJkfQOcw11koregYSRoXftyVGtNoWlWmy93vGE0FLyqqkez408O+4PEOaAV
RT9BEGPEq4XHtEyGOpKul92QnTQ/2wJzpREfkV05xWorA9N6fEtiaDsyX4y7eetMXKq46MQBQnqd
J8NNWWTsNHrCwKyxr9Y/tppxfWqggVxU5dKMv6Ax9kIIE56Q1NxWHOSwk17r6H/SLg1Tn2XpNslP
wB8r+zR2+I821iczHzYcX5AvTdI5iH8sNMOnxG8AjcK3RP8aFnuhmR7TGpAMw/kqq0X2MEgCOn1w
fIp3wTpOJeXHESU31JrFKgphk8OmlpSAJk+b2vz3EoXaLHelwJ4PR4EjT9fBAve3Wxk+PcWfMiRh
NqQ4V/xfvdhzu5x3NooljVwCMd+vKI9BXrnCokOTBSelk/nN0njMOJr7EzduQXLgdIZNufdOhkFr
JzAPw+LtMIv1nlhmnZkjNoNNjyKQ9TlY7uKewkd/w3ZMz9uaVYJN7+1jh8frFmRPE8Ijk24kkz9R
8Fxv0Ri2+7QZDBP30rj+TQfdIGBZfFUhP6eA1/VlKRUuGO2I2BGNAogjwBNcUyvP17jLMbof3+YQ
+cPkLqtEo5fIy0+BhC5CXsfz3w8cxM+InftyVX6Aq56qLrbQJ+AB6SZWv9h7Sh+kk5xBxr+GHket
hSngPAY56+iyqtMf3i1zJdAhqx4M0LvhWYr4/CUvJNUTNytVZyoXIKKLSimses2kATLn45iaPrG8
0vn/BeNOWoHlA9DCJ83/zrCAkb0R/e8hiGXi6jQQZPsO+9/n0SnpsjtAvfyFry6qSkdLpS5WG+PR
ZQLU0mtQPzDpyZlNRKVQIYNy0sLJJMhyTTez4T4qKe0w8RDwIFjxnxRTaemFIkyBAijMyf4d51FZ
FlB/PYJxAaIPSki2VSnWHp5kRtgoFgYpCi/7VBb5c4OeIotQjNTDtfBwacmIs+Ulc/ix+jgmLzOc
akRguVWvD6qOCv82b+O78OVQdKVMp2eDBIzNTqPxnztiMNdWlnr46Uhagaf/+iTCbXjH63snWRLf
kIFktiM0PHlCwEFRnWnyVPdf940XoDS/p/mdokv7Hx9IIR7AOtt0LBvBHhFdnPnwd2LNJ+g1a6CT
0vhq3lid0ixSy2uipdHTJ54Hh9J8/xQuXIpk6IOO9idOkOB/ajIxxQBvNEXB0QUvqnwlnOyeZprF
nKasJtHy+CO+t1FTGveB2SqShzr+e4j3Qv9mDMxZWDnAhcuIigLkRJYV90gbgcqjDFjBkjUnUZOJ
QYd4lrp8HKEmHh3WjVnLG6zFd5o6PgQqtpcPaKcfcGXWyBuskhRJD9XrmoNL5bWRVZUruD0kqpFf
NfKlg02R3iSnyox7fjCrh9dNLJ0OPkI9foUUvDTiNXVq23orSt2NPEvnvFC+yzwbG+f9U7e0b3b4
/lNFuMPU4Fi7YK5EEkLo9BX9mvYUJH0XJbPJhFM4t0zh537EvB8LVFe4bFsqrvnDiuGv7VkTnjwM
wiUhAMzYPsfvPudYTl9La2eVeamfd+EOHkFxA49DH4SyJfTyWDk+bjjmq/lEGuX6dMMOe8ST4peD
3lpSa6I4BLPot2hzMr8Z3YpvgDp/VFlLh76PuiKBjrjFdk0KYT5XDAJMS4dX0jP6tIU9YLLFlie0
lD4GFrlmYutNLMGYpbem11CqwhyQsl+RA3UdyirSg5qNCnBgFrxY/a3Ihf0JR8Am1paNAzM36+IS
B7qxxCpTbhQjCVXdWNAJEWiMn0tE4oNbWdRTAJ7dufhR682yu3TMA3kJpInv3OAfcz/mxwqWfnlS
LNvrMzaSKe4UYV/ODjCE84/OiXTHpKRyGGolmlSm7wVk4wXcRRSJ3vOnaGIegzKn+gE6lSS1b46L
sEwgIzR2VfYE9sAhcqs07HAdI0xNZvAnsVQZkB7Ss0htmPMhP+5wUhSF2on7/lzMRJ6piUNz3dT7
iuGPdJJiV3ABrpGEr6OPjRWBjnPEKLobjQUpOz2tYzspsmCIk0y8km7xxkS/ALMsGPJovtuJxR9a
i0YRlpdkbPEs+qy07RwejANXTUiwckA+AS5963v9KmuCPc9/TP04aVNfbqgm1sCDH54itCMPMGMq
6omsGtNooabne1yvU47F6Zr3QlUhoEZFZNWRl3N2RczCNWmbbTt/+roYz0TogL2ZAqdmJ8CqQ8ot
UTO/BsLvRnf5VSNXvDTQ09xgevhruKRa+vucGH3R5iQ6fJggqSlLVsXSS8WBQbZYLi7hWxYIbzxt
yEznQ6nC7rUherljgNZ5oyb8CV27/wERqoj9kE/39ZQNEEJ8+5oGrLBu/m7J2t+E5AnT75k5Thke
WPW7ATBwbQs7w8tlU2AMn+XkbNlB9a8JoWTvv4s+zm4O9ed+Opkyqxy1Xw25VYj5z99IIJCkdDdV
ocQG4yqIRfhmfhoOQ5QP4MhShkxZq/DPQ4CzYDfT/Rqv/LlnLUrfj0hWch8mjDIzXBqHlgZcMfc9
fN4whdlmTePEfjxIvmIKrebW75T2w314fQqebYdOfhltxGg4DVeNY2Wka7gR7wJkBd7H4W4lu5Lu
H9DUbeRVkwO+sVBAmRBOV8V6Qqk/Ts6J0pyct7oq57BGC+IiYX1hsLZhcF4vrAsAzdwfMkkOF/8n
SR/dFWsGH44A5dwRpnqWIaISYk6EE/AWxK6Y20Q1KJ3JslsX5xWzFLU72PkZ1G3exKcqGJ9Euo0b
hawl6yLI7D2AwTaoS085ovbOpgydKS8EXOE1C6FgdUUOVNtzG6lQXOBT5L/9g0wQ8YShpuG4+RDt
Vu9JNP2Ox8du4vj9bKNAV7KA5NsxGRtLsboKDfaNmK7+UGCpXqBshuiIsamfze6i01+/be8PncMe
ZVF6xy6P6vc688QpS91v1gFpS1QzagFypzdyCHbL/bwc4MdzDR3MZYJvJcVcxHFlSJYdPjXwG/bc
6fv+4tfW6m4AIzZITPVnz/wGVC4VE5qzcnd3k+79PYutMrr+mLqzoJD0fbDKxcyqtaKMFh7+rVsg
x6JUqNdyelLfr2elL/ss3jVBarAhIPRoaSjA8Mju8eCZY7JxtIjOs92gs51Q+yFekMWSYki1EQzg
PqUPYm9fwQxOzMqM32Pb4asr30MgMYZPP8R1T2S29oVcQ/r3r4nJqVMS5XAWxFy8l0bLMX6qZOFt
Ht4I0Lumlqb4N/Lhh2FZrpGuKIPLZOE/RSUbIxIVygNXZsy6a7xBdEUd3BCF/Nw2dFVxtoYlnet6
7nrQlKMKga9dHElt2znOJcs11ddJDPjJcqemacmomz3JFR2CKeWFX/BZsfhmDh3qWI3iZNu49ci5
cTvcGd/NhumV5+H3kSzR+H0IjWxzgaa0q25DTJYvUzBaeGYQ/yt9Bso72lN8OiGn/oySRE/U33vG
FXjT0hD4gSl9LEQ/SYGQvtYzEquEcavm1aGCKb9rDMj+WVBO9TvchW+1pha9v2lHMn3btFc42cef
JymsUtbtqD5OUDKdthUAZbEQQsE2RhMFvbj6TgQq0wjfvwp4avS1ywCa2pxUQZM20XlRMsw3fLQi
J5lhmr9nJKax8MDdaunueyiuUympgSluQscQYP21IpbVyk0Atl6pyOoQl8TzbNB5ncKYfZ3PGlFM
kNF+Car+4iGTOPoWGuH7dBFL7n7x6X0K6oYpvzXGaLea5V892GrAFsggMu/abY850gEAbYUFxRlf
DjScLrujbCP6exOcFZMiO/ZTopxux8pbdudQpsXlKm1yopyOpwk0mvq9JT6M4YlcXXsYPY2Jo/Ms
WEEN9p5ZmWKvpABiiwGcqYlOMID4CkxK1JntphxZww7XPMjEq2Haq2C7o5T+3ojrkK+gRc/KLRms
7Ld8PXYPR+fKKFWEpK0EoT+YR1KfGpW2jIbprWgv88Twvyrt8QNkpcGIS2FK9tHi5rcsjm9Q0igM
FL4pxh5mNfQcNgqRT33zbt4sYCyv5u3WGGbggMVH1sa1lSNa1Utarr82TOI9ed/BrVOhWeD0j3LU
zazBJUy9EAGlgnJRkUmS+Hb9mGX9T/VaXlQRSfXXW6MThCVfSRRopAMLeYuUjQKJPBIsa8lA0VR1
l4RcZ+z6N5MM3g0HBNXW1T/XgYoX2pEYFMv/uZdbsJik4s9mD60xMFlDKEMmHWtUktCuZWw5VVHj
sXrWcJwFICnsrpbp00L6irYfaahginug2MSkIU8H79qz7QBLnR4vNd0M020MujBFsNvhTS759OoR
ZsU1ss+ZjUEh9nCmZHZ7FnaE/sqfWN5RSWxeX/qi9G1Ki1XE9s75k3Zf7wRUhCgZcrWqZrDPTFq0
k79TRrx1H/1k1+Qveee9A49sZdJCmqg3pnQZ2hg8I1DUoiFA1TiEtMJRULJxYJTAzSKNOeWH3HOY
/xG1Oucg+KBPAXMOBP6a6TuuQeLYHhPnIEknbIXSKGCbTuM6XpI6kwTiqwnqLiWyekLJ2+Y2GIwV
iDZzdP4xGya4mtNS7OTa5fQU8glxnNksKPqtVCPOrigau9DiGEZ+nRarhJ/NlMGp//rMR/nPwBJ1
Nk3pxqhzMYXW4vTzNw5a8nLXz55bLGDMz5L9yu0j/zrNHQAQK12mOgMmgw5Yi3kCQP2nvyxdhdgA
c52bmd/PXsLERubLaoNHVQAkNHvcz7dfmVWlDRyUJDXypwI3iNh1CV2j0alPeOAEJqpksKv1VEYm
POTfczZP0/6xeS2qV6IjUmwdrspOCd3YZW4j1E3hRcTH0vi1hmLUnmZePXUoTbnrS/ZDLejfhalS
Fq+j5IfT33ammjL1823xeJRsBLvAZ3LO4qqnrmvrvI1qulsAr5iJO8vbQXMlUX1ez4TPtMGkb6r8
0iq3x+q1h1Ikes7doAZefAblwyQFScWTUD/nuAj7X/3Bw+MbmGR48cPiB7SA6COjgx0YomoLm+GS
aZAdxvgINRlu+/hseXujP6+PYj8ax2IrGLOw4MTigHpKM8JNeIYEeVOpxetGqvZ5FfEjYMXXNtY+
YF8WdmtsohCSkU/CUAxetHaRUgiwiSrTY1/N1yD71OCAxU109cMF749+fZGbcK9m4VofVmj+FHPQ
phqtGaF5jWB+FkFR3Huv0nn1S7jzl204pBJA/xZf4cvwmVHm/mQwQLoJAzIrZ8jnm/1PVFKnnHA4
ImtYRml9rD2tl+sK47fBrF3zaQqJAeJAjoGwMm1WFXnOPSE0AbvJ0uRzXFWvdRwkOfuETU5NgfYq
Sf2ev4w65KTm7mrPtVROfOdYwblb2ipaTirDqGhuo90nO/QPZt1+A6BrybszLxLPATA+ZRN3WjZ/
U/VMWYFapLcOe/I8xUqxW1tN/w/2hGuTyIM22tgqaAZ+53XgTi+QIvGwqr2X9DCJQQkUJMd6gcWk
XRuQWqK3Qln4TrjWbod4/n3APpybetQfE+rxY++pdNQMlfgV08XHXokpfGCJzkAgpVmYaBQ06xQ8
bWIGCpPKSJfkf4jotu19iNeOIhbpSFeVL1zvzUFFb7ssEhlyoJDqzlFUaWIZdyzFO3gNv0XNAp7u
TmnCHZLh4fkacIMtyUwjyuYi/xa1LMcuOJhKkn6qsX137lKyc3RJBP6imJnGpzwNFZIc5hOz/TG4
OTspaAPpa5Yq3zKA/HnnS8T2uoWvTQjxQnWKF4ERXPkivC50C4jYMgovEOuNX4nGzJYr7bknWWxE
C0LBCR01bKQJZIn/8ydW98+knt18VmiHAuBE8sPkuTQqivpvhRlaG2aXgHnF6LvKkCl87QSPQavm
RmsYXzYuGkYSYY/7pDFD6wSOUs0K2ncPcjGgOvJZ7ZDVHMEhKmdT4SIvkTVK1QbxyPXAh25KfcyX
Y00Mg9bKjHAWKoMjRiyD52YyRWJ7WHis9409AA9gPuHKVB4RAKc2hlr0i35VBRpy9uloZWaMvWQc
9S3da6g1p/6xwMcN6j0rfzousB7dALPGbgP2HLxLaS5X9lnVHINVKe84oYsd0d5XqMizxeAOct4n
JXs2pIZYG/rAIrO/u3Gq07Hy6ozVrfnZlXmZ8TfahZtMadIYOl9YWk53lYo5LWLkwmh3onl2cH6F
Hi5UhahuVaF7vs/+ACTU3c4XKaQMk9d+IXmmRd+p5R9UhB8Vl0Rl2xM3inBWiRY85ondxgMbg9Dq
gDBF5UDRKoV0s2o6AjHav6HEQEoegZP+w9mp/tX4swXh1XTWVN6mjYUaVOqbIBNB9qTOihLpiMR0
i+GEazidxmG3Ig/GMicLFVWq34B00xYrcIXFfRDVqmba0gMXFl2IfEx7T/sHwd1zK/uYIawB0OKR
S4PdDL4dkD4Cv1sSz5OVOvAb5l/xdoKOj5BpxGqyc1qUeXMj96TTW5zf1kuDKgzYzho6+/3dzGeE
/h/zSxSZ2o5szki8/2zkxNRQKk8XE4r1c8FkePO+KYHdc3yBc0GzrbmrcEqa1IxX74k/GFGYDEr3
cffLvrY4L7n/4zzPTicr5iVMI9I2tQzFLIutlxV2H15qb1JycSwt3dgiKoaGyZz2c8kwiS4bmuRu
2ngoyXDvwEZA20l6dV8YR5hj8YeM4HPELA91sDx4uUSPeQymAmROwVErfX9Sjm4j4BF/DlzI7Z61
lkkctcZVLe3+yid4H4GAt+vzSTkGXHqzP2KZQfBndEB2l8XFIAzyC2gXLGUNFuVr8rff8PzfaIi3
4GdcootDWsmVBuZ9v0G2UkscafW5kjx0lnEzmDgueefTVypjoq8iUxbLbYU/BZQP69/sjux8+3YP
kelJtLbTJ2J8NVcW99ht+pGe4zBTNO6xcJysUHENfTNrXJ2+yUtLQc2daabzWd7S5bXdCikZ0pBj
gyRD0WD1DkeSlu07wg+G+D+UYG4ESIcZVwQlDvUvRiQQK/lM0sca9hGOEIX9SwUZ/5nxqD8tMm+6
On8gGSMHwDjwUei/Fql6HmDDtzBknK061CxyXMQtDLoT5RDMgrDNZzenJXSE87+VdSYzxFzj/cQV
SLJJ36F4SupNUwAaZnd+5+mWnzNCXTx7xhDo6/WJrU6iDtNJ5RKQydhmWiT26e6JeTcH7oXjxCL7
6ThfX1ZZ7UdBGUpKr54dZV8Sve2cddC9+hGZL+pZxL35LrZ1q0fFPNMFso1QqHRdXWPvO19pVzbI
LAm2l0Q/vg0XhzJ4pBRASwE2ED2Uf8kOas/AW5hG/IhP9VK4jFusbcpqqrhLrZGfpYCWM8a01tz0
Zu/MjyQf/+/74zLKOZrWNDiLF/6Ilri3EBzWOiDpMM0QfbYorNfKVJoqteF6DuWom9Avi76sMJTN
s+ZgEFo7ADx5A56ggmRwONhELkhaoV027VX6lgZE2uZpFY6G92fKM7NrX3/PxiGJFnfsWXXph0n7
tOac7ndz7lmfHsZ0Ck+DSEbjtUO89YZE8W2y0b7aihYkpFKFduUjHJnrS8aLETDom9HO+Y2RJIwc
4i5MT8cV5O+yHJuSnDgb3/KLGmO9Sn4DBM96zZkqwBeJpxejDbChlpAR7Hy9LEPmPylJFpwuhFlH
9s5IvyFJHZqM8O8ngDbhRXn7I/xKzppFOkm5esIa6Eh+mlCnm5Y4+LCqMRZG6062TUM9KJIbOqbu
G4M+dVPfzPb3p3ZxSgW4Tdbvtoj2t07ZcOXGdnjMOsg9xVHQJrF3w9pYfol10RuyIHoiLWS1gHDX
mmPkzuJerB3PXda0H1jF/nSbhB/puN2/flPu1TpCDt65DBP4VHennF+XgpP6eLbPtNozApdt5qls
an3q9G3ZuG1a+rqfhT7P8PrurHjja9BypYRvoTTppuYs3DB+nlv+kzWgCPHrRmzB+Lkj4h1WkWVI
NGBkgl5iuS4SHWshf0cHBw3UHw5SVuSGKKeNNJUpDDk0goKw3q2aoPpGZ4I+ylFXo+c0jt43pE/F
8VcH+yq0toV3bBHAZVZfTEebQ5NOIOzgLIbmHTIx1loI9ky2q7I0Ji3vumRpBYRQNUoCLexmUfSG
slJkGvICo5gvqL8ecn/xv8VzP3UMcIQE4Dcql2wME55fZ5JxPFYPZEiu0PwBtwZpAp2AwKHT8ro9
8iozpr+KW0YQlicmFBxH2SFiiTaNt5X+1NvfeifGp9lRX0P1MEUppC+Bk7GL6cTHhJW967Mq9TZ5
LiE90zerBTea2oz/3pd8waYWNKPlXJv1m8KKOv+X+c+y5hUT6QdVS6+BP2CpWHIk0yqUc5pjgEco
3zvGaIDRO/H4/E2qzbAPcMaOltriKtIw389heNNit3xQRRCNLNJAhKUO63eZ4ttt3NiDrqP7HGzj
2JT3Vsde1ZbdpQ8i391iTYryn8FRnRSyj8xO1Dnnsj4GnTnrCtKF4Nyfe+m2xrgHFHJT/UBAhhPV
EeZPwLNKMZYel3q3genB36F1V4/XV89O4B2r3BGItttE6unvPQ/e1eY2lJpracLckjpi0H/F0T9b
fP4qTUhO30eO3z6Cn6CidmoT5YncPb6Tz9GEcnAHiCCmHMRmG7R9ClHEXuKqsBLuhV6UWs4vs/ra
KMcKauz78iT9X4Hp/97USjXaYkZL3S84fg1EKBnq6NUMZsX327p+AI+WUc/kg8dtnpqh3f56W0vh
UXwkqIA0f7bk/Q/VwaSmuACAZZXrdh1tzQXoYmMhopMVOQJ6V9Kst0Y8NTDkRRFuPd+u/VrFCYcJ
y+TGs/Tbc6cZn9AZPBQRLj4rPdX7ntzwH3iAn05+7jioS1lkZSVl5iHj2k9qIjpLYqdC/i7zl/O9
mhu5Z9c/90O66o1PLxqwHau3NvGeUKnJ7f3tBhfi9a13En0jtorx4yWCa35J75l2moc3I/MB90hQ
VrhmDxfDlDu/5f2/N3HrwJp/gtu79Zjj0Dvozx5RMV7sm+7ZBrPXnPtT+3+o9uR06qf6SL+g8nMw
7Nv8C/Ks6EeQgRSD61ee0T0j0mUqj1Gh58+n4GJQ8o7O8duOif4ZqgSzCfgIGSw+fBrzhOvGOUk6
Y7qDqaSmAhXgFMIngg7TJW6FDkNcVxxQOggoQFXbRVx+DBVEdT1BtIN5HlZ9GGgq1bC7jLrQbjiM
IXSe0KB67leXGGsPqFzgB8PDDPYB0bRrksf1Mb5HUl5Ew4CaHmDqod84u8rEdYtn8nZ0bf8DDuIM
xW4NW02m2nRpUUOt2Y1YLo2bvrcrYPMu9kKK3VFIBhpBmCaGrADa6EI/ToXVog7GK21S2kl8vYhw
LhhNAL2BUFcDm+6Ov+XFJjH8a6kBziMCCbSpUapSG5F+GHofKwRy6g+7rSrpyPMIF2iDCGMuZ9rV
9mIu1r9qchVCTZxpyYlqZn3O4wILiDFbiH39Ki8JETWVNJGAR5LNbVSKGLOx69qc5djL9G7tlkY7
sF3Qq4OyS7MrPhO2UVag4gRsuRD1BAFMUyMSCsyZQZmfAOBPpt4rTwR2ywpQOs4VgNcvNtC0b1tD
Iw3ZskngvDRN0tFQNcLeMTJrxv9TqEqkIumLzTTc4PvGsDcgfuoDw1Rav3odd8BmeL7VcjgPic+Y
fG4DjBr8T0RlOgquUQwFwuZ5dJfS88m50vVHbFaNAs5bfGCmGL6MccPGOsl2wSm4JOkgcd1F+iAU
8dmV69mFtIxPj4um5LruHofU//u2fsmeaxjiyKH6NxqKelsyOohe6H2wA8OmRFFuATHizJ3qouCG
1s2ZukQsr695yrZQ8+g9/zP9RwvLyzgyrPS4Mr7e1gMOlfOOjbpeWyXxiBA2Rw0hyA+2l8S3YU12
uJSO0IJRcwsrVu2o1sITu/DoKUSRMis9+K+qGlFx6sBuww2o5IHMhCERM8eo2pDDswNovoqIhXxh
kXLbfCPxkX6H0q4ZQLixRiX6rV1xdURtzB4KBrCO+/UcXADx+yzqjHCqIITaL0LdLftHi67xIfg7
fQ19aUo/jukl1kAzjPAHdrE6O72CoBOTfsFnxUQx1WIxjzTbQwANV+CFO/1qve2rPx1qFaOoV19u
h67mpg9cyoemDWyaYeD/Kdmghu4ciDnpnJI8wydfIj2+/3Q9IcX+Zsj8WkUdPV8pxbwBYiHnOPwO
qJoD7xDXYdkyp10/D0WHBimVtZRymcA9oiCMr+8aOP8hjfleR2+BzvYV4/GUoroYH99Fkb5sowjQ
3kuEI5cLAOW25ObJyTrUDhl/NyR3riifiPfg/EK0JbkI2D3JOe9NPDm51EJKjp7pa5ktqWSZCTrb
Eri5FtzEw6r0D4cfLEqOx72UxwoIZaHsgBk+XOij09huQzyQbjKlFfPKnFYWa/1CVwB6AsBYlBV6
ThG0t0f7W9G8ozBpsN6BgM/NagVy/owcXq1PHiZ4oKuzufVvboyl8KT2CzckiZGbYXyCv26ejAtn
r+ftR5ErqmrI5dlr1Lrr2IL+QPB4fA0Z2c0d9DAScAl0CJbgZ7iBvRifhtOFlP6b3VsUNs7FZOKu
r5iy/lc2+/hy6EDfhdip62U3rAM+FA4WGwh685c99rDoVvvxalAJcCnviUaRQyUrBmvZmJ/0m0dr
bwzgIV1dDAxm6pnlRdFZFVAVQOVJdLRxZAovi8+wmthewlI+iVlhkJgdAcHwA23e9d8HL1AfqcZc
2JoIsDEwlQVAS/JhOj0QmqFb0kYY+N4YeVCOGy8cR/k5YrRaZ9d3QC4EfRbKVP9IpP8/b4aqC1yB
uqYH4BfM9ovI81b1lzV848vPoiHN8ncixMtRL7n1XFXOFMkVCC6CN5bMYIsAgXH9n/jpftq6F0wu
sDYIkzGuPcLydBbI3j5ZOim5gW8K/sY+iEBhMOAqIK3JYLwbl5pJZCX3qL95p2AIaj6eVOHIQUGu
qz/3kRGf5ZVOIsKz6o9dxIhcaps0uhMb8RiKz5Q3CEjbqLNTf2WsTysomyCO6UVJNiI8zQXcQXo6
BG2mmAVzyGPNCJR/H2XO0qivoy0RN4Pk8WgHTbP5U7JRFclt5tJzCDn7pp4Ms2cFdrJh2y9R9Mbr
FR20F9ALRe5y00gUNd2o/J/MM3S9VDnHIrrBbP0EDsdMepGpn+P/2SxdTn6rXp54X3FaSlhX/FGv
qYjZTa/uDWrODubQcvyTfv/YKeGWV1H1f8LVkMgQhlJTtk7IEgysjE102Tg5iFTCg3XOZRFc24OD
j8HDI3yb7lYDwf0E3Jt3wncSN+vUQDddfyIIg5KiSNPapwWeTvnPfDFy71sBuxS12g8iwCYgV5dh
aowxeCdrktEs3etslvLi1tPDYwj49mHKR4MRtBIbPNeaSHu7O48eJJBfKo2m49OQx3wa+hXa9SlG
kBezjo5aqumNOjwsq4lr8722jH3+/peg2hUNB6ByRZZVXPBJaHWlwehi0vi+jw5vZfmmF2Rc04IA
6KM5Pv698Nfk/pwlhelF2g8ykt1GmV4NbUJn2K8E7ne78Kb/iIXt8QJsUsFhdLgXVtfpoey04SOb
kOL6NErz+WXiWxi1QaUekAi4/bxV1P286XDFoEzPakWKIjviUq3MXkRELpIhBnzA6S3Dt9WcI1Zq
pENAqW09uskDZBOxyrbklCTfXpMjMDJIfGJESJhdFDguli4tOloiAaP9wnhhUqIwSw0AXJaVTmRK
53yupfHdwiiLOUpvQSpB1y6sGXEaRYbrS9TnIb+3cX1N56OWq33qop4+FbOgqqslfF3zWlYFrIEn
bu/NFwlZ+C8POW608AiZinJ1gYlVzcDLpNFnYeqS0fOnxdvpRYSXvAoq0EiiSuar/bmvMQnRjFTn
yMtChjkdcqyF9Nj2MumYAK8ZNapEInumHrodCys6e34C7ithYutsvfiXu79nmkrPwZ3KvIRWu8aX
+S4C7xXa2etSd/6QpdRdgRymrhRBjwKec3WG8yuCcKshODu/3rv+DccVIN9g0sZJBglhEHySprv4
MC1ynLhasZZlaSQlvpWZSdL3v//r90qZ+08NHBRonUv1nzg2zmes3iIpGmcIVC0L9iSiNlYE7Cky
GTvak3pY7ugw6By9PBFoVPpNHaz7pDMp06oIIBK2mf9B79hsXY6sWiOFZ3KAIMjpdLmiSRmu+wc6
Y+bOjGPPCkkrFQQ4t4gzWFt05PynuKvua8L9WUwFO+cfG4tutr6VHEyeE7O3CGf+T8pq2C7HoOKJ
Y+/NyKn0EetNOSdd0ieGR0DADzgoYsVGL9OFmi5ATnQFDLkjdyd+LSGXN6ShUl9vvfBV3bSgEBCW
2KUUig0NZRCkrgYCWhWwNCRNwpC2ScR8hkJu5dd2yiG7vskMgav7OROBuaIHgoTSt2Ai/C7BpwkX
jnm3GjzdLHqOhJMm6ls5FWWxAd5kvQ+KcbJIeLD+EkLsvhWiPlqOYq+HaKNRI+8aWVbAtgO1fJIr
wc8TK7HFZ/nqe+qOEU4mfcf5pjfx6NF2BINwmZOPA/kgZAL/HCbMV60gkcmCmJnMfGA6K4GEg4u2
/ld8fRVIC+kXaFhFn8PDLMTU8lrgM8/Yv8WyYIBm2dCLzQ6hoNkuS9ns9htLqcfjaHgeVsooAcHB
OcT4d9Jz7XVddCtXn+3EYpjbk5/YFAHjYLjD4XMIe6evMM6rhkJKJrnR3qFCgMdFMza3goQSkWl/
87ezMHh9E7QETJsYkg68EzMI9y0yzImgrpyajE7LwjOiwGhp1mUyNkf1Tm4e71e/SJKxpnBcdwme
qYBzyKZJxLz87TPEVH/2jFOc2TMfNIgHwbewUsyoHLLAQo+hfcUFijrm7ZLFP/gBfQ6dhZf7+raH
umVpdYRev7pQjFgmHUZ9qufEfwmE9fqpr6Q6mLWWZOUS3PLrJ5V0rixodh7Liz1MNFR+i3IMUbnl
L87tdrlNI9uhN4mWylu4DFY3W7Zqr2LhawVKm8TLMdTPLFBzg2ZqBFDDCmkivzs/1iiVMnyWqC9u
xjbNHpv/ZJWhU2rbIS8IKv+eZAx+jKDjHHoqS8NY4ut+nAtrrdjQ3vYhdDMQOn4NU8CbSPqRrLQP
MYGdd+YtjCozGZtOyl4cjgLKs+rS99fMHJL485/dEtzmJL/0v1Ui4l44vWrTJzVYAaGB0/Pn+03H
/htTAW/lNuXHykbFunLfxmn3TN0jpQQExrRulLQtYcbNPMgSrRGx6YDAbdfYjeyv1swEGVJMekfX
Hj0ETOQqh+hKOVroto0kgDNFqAADDBCfRIKzUssKT5r/IX17mmGfzTGsh7dF96fg6UJgl9/1HK0k
IvqW8mY+0gSjRtLVRmIDrPnyrWerfpAUeZ5a2yJ1ufbF82cpRpDNr3Rr7BCESREaa0P9msQNdM3s
wF5R1h7CHaFoyRiBQUdGFDUJ/tvYo/uVCotn26RSvj5s8zGO6/sbF7ibSqKYp8vdZSird1fZz8rd
Fn/mCmIS6bzB7ZYPGjE3Gxp+Dfkd7DPD6unXnOCpdE2lcXGQUsb/rWJroAmiXufIf7fl36OVIo9u
Ay3dyKve0OVj4x2NPi8sBMNuXzv0pminD70Wt0LemUDr65a/Iy+cr5Et2S0fuc4F9cCdFCJaYD2P
qB16875/VZXxAH+9/Ft5yRy10X56Osf6fNdxkpp/loTmUnwnPVW5KIGdIL6rB494cF9zbg2TX1Pr
Uw33xeW3Qa6TMgnKPcmqsUrZuQc3zvVmQXq7zY2BhdGMygxpX8yMLwMAqaTUKk3DlN9FK78CpmL8
UCiLCnAboIFXvygiIm73T3aIjtu27WgI6F0IfQdRcysyL9+5mT/VICSDy6+40Hw/LR+x/S46Wb3m
ss271KdtMj+k013uT+tz2GAXee6AvLdlLO6c6v7dfmXiwaU4Yn9CmHnWCEIt43HvgPlBtv3yChNR
T1uw385yYucWYiYM/FJgWW+Lr2dwCimij15PbzwJDEI8LdKvsB8zBovhl25RI2Ktyw4LtNEq4N8i
/hYNgBvED81pqepOGklfaXdQu+1GWCJPtHh5WpsXQCi/EMemu3Mtr4bLKzX6keOkvmnxcs/8XmdU
/DnZZ2viruodrw4a9dYcZ3I+Fvz41Q2No681vZEMCf8AgrT7PV7QuCW7TnwDfsOZwqZ479dvxa4L
WalR1E0mSc48hVk19JtKppJS0c+fA1jUNgqAz2OQmfBqHg76MPKpr2imUuPy6S6pUxWexshgGEly
DDyYWdlbBtca6pGZEw2Cc3epKXRgyTfwpfvCKmsTH5Cuf8iBXotaZGudrwq2HTdCULO75RWLExZZ
xAt51pTEvZFcr6rgOv9Vt8LELrrZLboUQK5ao4Z2n/mmtW0uVitWiN3xlsBMCQ98sZv5iqeboDoH
j2QwQX9QFIntLoV7OJSoa83Xo7uqO9w58BDVuNavMgRU2mgq+4Ir4y4V6cKbq79lBxeXRm3MmmCk
5IRzIfqvMlItf4j+5NsHVjNzhKHH/Hi0tt+EHPsZrzQyDWsCnq9nR4H/TY2lvWfEfCmdr00swScx
Es6uHEjB0MjA2618huOJ2utl1MhCtQ2gp62h3rOiVKGSN3jOemjnTPeUlh5qdJwzMKluv/0P6xHQ
OkaigZYjtOwNBaCbGKxrxMfWqMKMoOP8HZz9iDjenGTfWcduCgK40obUrlSDUZq1MmRV502edonx
exDOicV8ZiOSofBiFj28wTqyLLQa3xPG017xNkm1kC+wgfTyI5gUFg4BB+KsPGe1lAQuuSxeOaW9
HUDFurbqKGswkEO7n6pS1PU/UW+KijvyTL4ahcgRkUa563DBkEZOzpJeyxa4C1LoRIBO36K7yGIU
753THsstz4PzTJ70tc6Lm6WV7lOE0pKTa7gZvKGSK3K2ciod5t9GerCEtrMl2lExhJeaQxWJUKpT
cbjA8Mn2m+U5pePoZOPns9hXfp0wpKEyDggIG/o7i9+HHywvCtEKbhg/GLjyjHWuprJDMeCX+wQi
97AL5ieHGWvefsUlDYF0ujUCEK7tawV24Xh54xSHiBi9SLn2GFyysn0EF9Ujg4sDUmAbwstWvPy6
LOe81dzE7hEAJP+DLjpddyY2fP/GKvUWZPSh2nslhksFZzNwfxz8htB5VgfHerbPTR30k4JAzTOg
Q0iJl1/ycyJRxO9efosKrwdJzgKwB4kHj7DUuj5kFQFLxjTnr8mdYSFGc5q94Lp4meqiW59Y1HTM
HlsNlji3RjsfGONfdxO1H/v769all5TqssKUev10M+iYGnuLQOw4u0c0/glrKkYV22yq0wB2f3c3
Qh96puU3mum+xacQiXtzNqvHo/EfHAoH3bcMoIStlgox62ZZHepHthdqQBchDAxw9p6iZ5CXAP4V
5A7IJHMBR/Dmn//QjG2WwIYcabX6ZqZZhRw9BacXDBDuLT+B5lKDmZ3hOOPAWM7KglB+qlXocuiT
0AoFazstYtL8ZwitwPq8FUFbVcKyJDZAoKN2zhnaBa/nLzFf4j2JEqG0u6rctw/3+7KH6Xxg6U2W
Vdy17LMYundIpsz4NFWCFbXRhIUNqEvCnExXWOqRjocuIJJQTFbf1MhFnlil2f31jO8u4NK8IvDD
Ohcc4VcCY1Imb5Qf+Sv5YRIuj9rO4CsvIE4G0TogguzEjeCHmYZ9mePrira5yteS+JItaKY5l8Jj
3EGqnXb7XwjOL7mx5v0GEe0vlz3isAwY4/ZBhRrdelr2mkdmNtAelvrdaEAm8RWL+Ps0dUL0aVAY
Yia09jLNE9poJ6rLl1Tbhtusw/V3nkUwfGVTT7VQqID8m4hGXYwsrdzKtc269NNlKzs5W2TBAX9t
HOcBNSReAiY9/okxvIbYqDdNl+TE8JOGBxeRul7Cln2lVIV7ip+e6jzhQGxaYYypcgHTICly/8Vg
l2J20IOPirQaVjyL3jkJ7LNpB5MUXvNwRRpKf3We0qcNcn8jyweyKr+oFTvgLlAQRnKZC3x3PLS/
rmIUPpkxc+wpdBWfydgW5hiAKOcKL9T/tw7+fyySzRqoCyWtQyufcCqeS4L0eFoyFrDN9SivixXn
lA+7C73tPtOKlr7nbzLolaOI6YQxYTDO2aJOofEEHki1G3bu1ULJuuoUXYtlmhoNSJEVe1Skgbou
kDp2AzDOUmnF8uaLihXHmClW74vmWNhCed+DNnGZr8kPyah/Xkd0Ak4BKn5Qt/yd9r9wGBtVAUSf
rPHNPsjOwjGPn8nVLdTWuBF47dFrL6nsMwWPkbJUmnmHA4Z4uZep0XB9Vs3AV7PRa9Em55pikP8V
1WPFkVyP9rEC0DZ52NmSnE//N5mz1tiza/5tJYmwJvoZHB0GTUJgoMxTyyMsTQa9Gfeyqa5QljuZ
V/D3OnC9ohlziQHLHX9Dt+jOo0Zd+qQOh0rn+VOzBItxKByLRZ8h6llB1p4tMxZuKNX5SVKyVUT+
XLc4W1SxRFxHX676Gtv2EKTveKJ0uLarztYlpjvAy8MbOT2yFzLmKe3vzVka8pFvOTaC0AYRMRFS
zzGEOBnHwE7/X9tqeM48LT9WWnJ0/1DvYiIP2xvL+6XHVvBELqxUwhIoIEfG210bVmQUHs6OWy6Y
CmvUCWmUZNeJWfgjEoVhiyIgwYi7J/oJHdRdPV0azDT6/cj4dAiXzbMLfh+4ZnZbchTfyoJzVNxT
MNg/2izCpVJBeoTpdH6847wLjI6xD52d9LRtoCeDZNemES4O7YWOlpAM1ZmvTurkIY29U8MN/HG2
53LqtXAARGR1KsvHNulY/2Fw3Dva//ydtRaruRNRik0M1jYplMhHE60T5aE5EAd2zcQo+tYbAdhC
J6/V4bkAWX2tmqufTTjt2lFCDhbHq7e7SeGpGgHXaiFgtsg4jksGwr8XVBfY4Doay4V1DZu7DNdK
2XtieDSmZDCVv6ESCK+krlnuEvyaYjL2N4g3JADRXOkvf2lrycqpCjWd8SZdZXHsY4mFPYG3DxwZ
AYKsUo7N2WDb/vZrzCKBSQbk8+4doTT9wvkazxFTdHLHIl8dLn/243mb+ASRQBzzw0e10pH8ELHn
Q9nZK+ATQUgDL5NxzB1AkevQ8IevGiQjIriQWynGSCsX6NjQKKsSsD+/ZdGGF/xnsoa6tXaj/DUC
qDBpub0Fm4e893nzTAb8wiK63J9XbnM7iHsxIgLk4FuGhMExsVUlqrip03iCnbLPB9bH5kjPZghr
o3buypnrptVRPRIJzYZfyLOYjOIX3FMsJy8hTgDYee59z5JoBo1L3Y+QdNkDqRqR04l48x6siWxM
ROq6s0r/QDe64nY8AjqN3a7uSlE7UkVbokVj3TkO+nDbC67tBFd6JLMnSQ6M7kuwjY6FoSRFiKxC
8r/Ph0bzZrJh+PLj95Wj9jJNCMFm2VGYnI4aM2K3iKUECvr93NCXJn0pA8ekPFg0XyPcK8WwgNaL
gue04Dz2XNwiU9r4CDWJg5uIzaB2TC8WzX9rGyySdMhylV4NndjFBbFapUnRiDnoa32E49B7h84f
5QglyRUe3mh97W6/bfCRsg1pvu7DkigbLeL4hBd9qaDcjsQbRH2+HkNJIgY+YjYakA1WEWpxZ3sH
rW4y897BQnRxKDyEoFvaAEWd0Wx0QXwyYcJyr+OBYO3gMs5mpXRjWnX4a7rhwAO04gP8TyhCZft2
c4UYjcOO1MFNEmFwXkfWGIbu9hQun6dccWzo1HzccKSuxVp+uqOTRW8T90ZMhm4lOaySjq4iLQn1
pvLOUdePEzqWhPQPtRBA1pjpHIfSz2r3h2dJcZUj4ULMOtAPHRB7C3QHGkhHG5DQvYl66BYNGFuA
Y6I+Lbcm5MCbIUSgOD4sQ184F1LQ8L+ANZzQQDq/BImbjyX4s+cS++i/+NTEG7o14feUpv6DIZQg
8EN8FgBk8QZgTQzk4Qvf9uRTdAUUzWQvtl6tXbTDSxWD5aUeXlV3sK6RduJA7Mf0XRlWAtiJXeb0
SCORjWccc+gX2NOnLwXFZpru6TucXY8j9a76ck9dujWYi6xmcr4GF8oX4kTaO+0f6cyuWaUkNREV
cwkvnvwzBkiuEIpP5sLSZDDFdDRVqkdmLSyKZlvueo5pM3D0lVZgxg6hhLvFC3A5mvopKfjGsLZ+
GrZEOequDFubYojOYIDRhEJsSoUwjk45R7Q/jSXorQ+c9xjOc9DKaJrbzeh1yi7ll8E5pjIFResx
q1YC+N0yZArBNBOMkYLhXtMkNmBrKflJ5WrYBuqSY8cJ3jUNy9F0hq2US84ClOTjN8ZrCyHpU3Ch
fDvSAQxNWoE0n340W6PFmP4+bWgRpNxMiusRyOq//Qa1vxxL34uTYzFTRJM2K7HgCkm0e4hCDVuA
7jKEfg3MJpRNHB0aadazRaDut3ek4Qg8r2Zt6gyaw2sBjoERM7xUjlXKNzqXCipWmuHhQRQXG0pv
OmTiQwPdME7v8W+LBeWo5eTA33ZapipcOaq27AXv6ZoZA3+YUZkDa7rzvzZo0Ipdocg5ukeizlFu
Nv1I3avdTjs0IwuBCCzK+lfzwP+DuL2uK6v7Z2SHGxJCfebhl3zGkV3AL2509LeOdTws/ideI6dG
2Y3Z3/yUDMaq4NiRudkpXswPe35Ex/2IiSsPDfc2bHi9lvrX+KEeyfSnztgJxend/WyXeI07Wmnl
lRHO8/asACcWFOmDmQIjaVzsv1Mt9SeiXeU1BQDDgBkhc0x8rfON9Atog3wEymsllqKu/xsSLMPf
exnziOzwRSj/aZH/bfvl53og3Qq6lgAvLoySQNrMC7W/Ue161zF4o8RsQhivWnQAiUq9N7EjCpFn
T3ggUPB3QWNfhYuhHdOiXuSJRlcLAOV4vcP5P+9rfqG8+9yUHLw7SMmbeRgoQsXjCM5sseAWBhsO
h5xJ/wzGRNcXSBwe/i21eioNaTTBuCztfLlsI3Yv+xmFIdFwn33VDmrZfsfiewz3z0BCN3oe6EV9
IlVZTjY3m6Ag4nKd1jj9I6hW9l78lI0X9oCQ0O093dwueYWMFM9GZzLNKmaOGO6uNcBR6YS04Otu
et0T9/Lx5AOvmTMEXXtnZeLfqNe44TT53i+5TigKoI2DIMyKoX+ZailFZ2b1TZ7sYEpJnR3mxWuW
DwBuu6jw7eP+dRU+idhkpzAUIyPK+RbJaBevxRb/h0KqiGWHQBMm0QacAcrcZOy4CoOrIPeaP7gO
EDzYSZUIQLogaU6tR/2BWWtVhZ9vopgd0+Cs+yr5bArc8+vW8VM8DB4429fRz4m4ycKGRgEk0C3x
DcEbbD0x73x2HKbuFO2XvMmkiGPGLuVZPb5U8X1rY4DVNS/a/PNfCXa5oygDwCc8eq/fWTkJMKQf
VSTDCkLGmij7zZ2Iodrgb2DwbQQb7jcPp+w81lr73jiLVwdTkIkm8cGVwUqaRBJnhMP6UIN/L0Q2
oFQ6AhsQtoCf4Tq+BqJP+YmSiJt1Q9jiDfZIeOuHIKoOvRzdUDu4HlBoLn0ebb9ipK+gasCoxI8G
7x9bYe3LdJ0BKOlykdndATXkEQpdyk2zX7AFNW8WG0zfcfYwCS57QELzmUKYiTq91oztC4LWRw8g
3DkzIDx25QrVWTYvj20A9x3Z3VFlsFPwHCM3j9Az7tDJ2MEegOfwiFAbKF+S0LjLqqilbhdDJonA
vB5dweRc9PGIGAe2QtsfbiW/nqG/wJRgfhxS/oQgLprSoGC+pFxSn/9CKm4Jy8ayNZBdvI96PSTB
woMxZv9UsuakQkJmnh8hThw0wvToYdikHrWSfSoGTDo0NaPVfpolbcmfjzLyxOhhSVVdR0kwqi9u
kzpG1g5j55ks2MMgIbcpEpXe6JzLsic/edSiMR2Pn97WVu9A4kV37n7TLe9MfxufHJcKa0Qb3NRD
JfX4lvNfsVgiTlrF8P8xS4TgwxAkJ7Hm2zUOp2EieqeZYMghPvrNNcANEPSH3pEkicGlkvmwlhYF
VqkQDzN+A9fdAA6/rS5J76LoxIPF4e78mG5TC3BDRvpjhWoHyWqHw0Sbk4Lgje14CupzmBx1K017
BIOFlQz4i3X52SXqS+eR99BvZuJOdUYr4QMIpKsTiUySN6I8BTTTN7dHXcehh1wh+BEVIQWCY7KO
QsfKyzFDcv5FQKltQtlJqiW1yDOE2CHneTYJrmEiq3Y0eHOxdUuldbnuAi/4fZB2Uu+G3DPDRehz
7KmgU4dco3fEeW/KgLLFhzDjzMrDB+ORP/w0v+GZeHbErGuk0O2EUZenlv7Az+QLRi2A+JnZsdsA
fecYTZzJN5kkbiDUr/anLXZdeSYsxyJHOhRDnP+t+GAQXYiX5JHN0vYe5N00CeVvoVw5Mk+ztdUV
YGBCAZM30ytvfKJNmJKhWOWcxl8MbODiLEyZa3drIMEjf7nJ6iXcO+jE9YLaHtPwq7dHluOIMsk0
JlQAO5i+IsAiJovk5St2J5sK+dx0qnyTQVXG5u0WadlRkIG55mwYzNnBHmTC68R8igsgsCsQZB/W
WSxMn7AZDgrFYA7Q1S2ZS/d3oJSMnxNfPD8PR1okaRTGJXYz4KqXSk30dd7n6gsV4HLdmcizXiEW
2Wv555RXEbazyGigAp7pyszibo3Nadi7uItOyVO7NSrOi/U26ylAu+OL9NUMw87Ap1oMEChJFJ/J
glKhDKc1RFOuzqviv5yP8LQQ+LycIEizVmKccNA59HlFFA7ouD3Ge5k5dHbpsJPUtiuUVEjDktgj
h8/Gp/X8Vn0k0bFmhrSXD0zzBAOoP25k4hEcHjC8+GnfPwy0wdI/LyXQaIHshsXEoqIPYqDgKs2p
8AOsCXa8JfWu8VSCTGqvsRLxZVG/yoTOCFHNWs7B4sP7mKpbw0Ps8bWTNXkXkuWyjbNtz3jLVNcx
ZPInoynpVqceIajon+9Wd4m4epQWjljhAA23p5oc6Y75Va6UUkWzrbEr+SEKpjfUFCkis2SKOGWK
RZEOzciRtetqs6Js+L29vxZ5NkwlDEzi/ElhORlypTetB6ZoQUgGXVFKOkfTFf2j0i6u7Mk9jk9H
FGc1AP8k3q1unX7n7RsBKUEkYcIcvoxHVqwPncSDjl/Rd8V3fc1wU7X/n/h59GUFT9eCiJdkG9w7
/OBCtwA2XIgXjdMKFL1QQ1pI6D1op0gM1PpAzr9RH037Tz2sT/djs+amt6pvmqTjCnLb7OSBAruy
X17KHP9zQhhGs7ogOLlwAED8k0yuV/fS3KuiEInuAq3/hTBFJN54aGpW8cBFBNApsKT+n3njoxOm
vfQTsbZUgJEC5hpEEWC6Hxw2yab4uBwmWnQgOEBqsgX4rwRpMVoLHJHL/XttMJRvZMKWpzzfQ9IZ
yBTNUDs0UwVgn9IGl3020XChv94kf2mbVJ7d+ACM1c4Qg3xKZ8mTCUtAwrxXwbEwH//AXVT94jrm
GRgkr3xAYvWLwQM9vUkJuR9Fr0UphAYLVW00se41gQh8sIbDO4AIHuQz2PEibgxE7S1sc65mlzQ8
cFbeyZz2AvC1jEmhs0eT0iRnGes20O51yDn0GQGBj2C5tvaYB7taeGZFM5f8TpXILaKty0vMACJs
SPTvMUPT4A2kUpK9mPANRmJss9G7vN38hEEiaojNQON1l0I21Rygpnl1PZMhXtY0YkA2AOYh8y+e
ru++LWSiD5P+FZGfRBC44zyAvXyQ/q0C1tiDYOTh/Ton0N5At7uQbsISkcRy+X3RYga/6Ygec/nT
IPzrhUQalN0ue9knwLUb69mrFteP6n/INdYjJV7LiKbGdjDgrcF1SBPyH1nlG69baj2jQKonmAv6
Xz4od2PsW1GuigNE9D7mkrgUBzTVwOw5NR9kRvR3pxFgHF+o7mnFrxEx8cyQF/pWUksBah0HiV4i
DcsGkULEH2RWEsN8lYNwOmN0ObCVFKe9CW71aoy6mMify3cxbOzETGLZpHD6E34Z2UQeGepjlNpm
OdJ//5NxYohkGJLtRFHYvGifkL8GTeuxSWM6z2IW2X5NWg+Bs3V+CC1zjMFo9kGnaUgXBYBgHqg2
aQCYJ75tPeN7EK3wprga4byRuKVYM3czqtFK9wmSUIXAMkoo5XAhceJMPp3THtUOusmUpUDlBPRe
7bzBA6IRmxH3/lDIv/TYRZj3+2BzlQ8vvLpPTcTeNZ6pk9Ap7yj5W5CP9ZLJFWMUlBSiFm/paV4k
TO5OOnXnaZ+cb7m8cn2TH2PjVAj8IAJTmz8ZU+Kmf3T6ZYS8WCqfZavWtjK06iK1rAU5OnZGY0Sg
Kdchbshaxhf99yslyJYwhpC4iRj32am0DSGKTHFJr8Pvpykbd4HZh5UVev5dbLwPoWiti2iVlGVf
HjJp4J0Op6jIJQKs4m1bcdQBn2pYFqhrpeqMO1NIG6NIUtR23tPbZFXj8W9spu18MBDyAP6ybp9h
NqG8ayL1FGHqudZ74iXPZGVXaNz4uHy0E2S8/LuN8KVMzt0pIlh23xeu19lcpYGdb6WeaQxOAUl+
pQM/537iNHpCWdUWe6uM3zlBdFuREVRvvgbC+uOIdjJXL4OOAT06n1horY/sEW0Rgmf/gKUviiyT
4eu3eYq1HrFgMUDiMsewDU/lKZsDYCvShARhTlyIVBays2syoI9ou64jzn42h70pS972F6T/et6x
FrvWejEF4ReVk7A9Rw91OY80cMMj1/F583r5oYKpunh1HUSxOlbhR7oXroUOj3dZkfX9y1Y7p/0+
6oCmFdSZgn29/Y5dKsG8CKlUV8hGNkUQ/vEFRFNiHS27+AvlkHVfFsNrtC+q665//pU+JBtGkobB
hmfHkBoOgASzlgQIhV3Ef3AD3caBPyo3ChfrINXeUKCrrsgAhFpKVO9Irernn1meRJO315vChN+i
MJcK2FV6JVTz49DofZCg+WbWl0HUWaIqKwnBFFtyJMQszlmYU1cqvUNX4JOMQpZSVJmioRkCVaQ7
JQ9+klqmQKYdxHmzBcxRB6DqhsSGS48FtfH3Wy9GnHqHhIbZzPDi2ueh1OGezXiyesolEi2f1Nbp
tyOKvdQQMDjPsH0+YVggV4sieyM4vXLicfGT0A937kIRPsUilw9Ik8DEmztuPo6rwgBvpCiE/JdU
XQ2IIzN52tM7+N20p51PvGTOlLfnFOzahzxrjhdgRXyPXsJOpmKM+LCTFfRIEaeEqpFx24QpC5Mt
7EzA2u362iYQ8qUR+pwfpieqWOU0pJF1cFZJOKh/lFQJFqDLsEfwFrZTpX8qSDwmuEqQq1kfJms7
Hydg8Z/3dkx5kuhYjvBU6q3gyk6ZiWqSx068nwyOn983YReaH7L4rrt98jYgiIPoQsK7su4v4IPz
JmCTHdrBzL8e03/gdmDyd6xdWJ7lntOayCYLO4kNWZJ7rlYRcPwbt5U7UApJAeoift1cMq0Zpxwf
JoUTvrJjMEe4ccumKKFXNp5duA7sUqlef6cJtz4PXUYKL/EofIWbOPJZewR/k3kKPoJEB93KKfMK
Bj0Tf5/7SF/GqoXhywUIl4YpEWTwB/3CfdatE1XKNWgyqWtgInPBYq/BhsPxqqlOIpee75hWUNej
27WlkKJdAE+SZItsFaO6eDmJL+/sJ/RVCupfVCnSgt7Tw6AQcjto6fCcGgsseubT+YbZT1weS4lR
4wLRYMgzMn7RqxL6sxq2C1Sg0icoHUdn3QojnvW3rstctxmjQi8v2aBEAjulHwCoM7P93gGivNWo
1oMosJs3xw3wH4jwoMUDaPusTu3pW0C19cgDmlLEDo7sBMXjKuYtUkQf2J2PH1NeiotyXLw2eAC0
W9L5YMVLpAUY2nDXnrgKkx5axg+rLF7J7z1RaApu+lULK0YuKgmHUF2VBpPWggQy7uw6z7YBJb2t
G53WzyxJyZv8xQyS+DHAK0pa5/sJKFNd3E34DCpBQAItF0cQ0VP43rzKawkBtihcEZ8UF6CERKLz
PWjbef9KLKtrmMXCU18j2Z/dWYAhpCFu6xgtLZnTjTs07bSDgSE+rqDDCSH8fsb3lt4VabPojBlg
V7qN3PZAwkjpzk5jq8/CebKlhx1Aq2tMwz+J1mH2GSI+Xz6JO+w661FXMm8epKQ1hw5z8J28Wlzy
zCdS8re6ptXiwsVsjTI4LhUjHlHCLtCFBLWotsrbaYFdgRQglrPl/NDBZHejSdjejTUFVUBhpaGZ
jUGCcbwvBblxocR9Q/l4NLN8YtLoJUxJb2BRSvE5nPfw83IfCxSay9I6EqMqMt6mAVof3zhEWWjC
TcqzW7vrpgNd390577MILQQJO2veFAxoWAVxy127a3uDUL9nmkq3RwSQEewjCE1EPG6oLJ/fyjj7
QBJDVigjNjR1pxBCtmMJdLRyhiq3RiWQ6iXpUUkeN0hNcdrpHW2+9c7U9hdegNf9mMZ1ypR2RZdI
kKRu2fYIIh8saKCMAJ25tpaJGL+NR4zsDZloXANlHHxmUhFyUpp/ndS1ppHMAzMqdsu/HJXLjWpX
Kq5WkNZpEPPdXWTOI4mzkkKj/B29SG6yoM+VGmsdFeTAs5NGepBAhgP0EOSu3XNeLCI0ecJA+GJj
QQ+SmGE8GhVy85FUZMT1awQxAaRbokkL+1rnuDKWHsU/Xx+7J/NZv5zCxwEePtFZtDM781bCuW93
ertYbVSdUgLGoS68+UkxBxYsF/G0VrFzRN3Uucb2mDa9VmRuHFcS26AsO8hn222xsBc0n0VOG9zv
ic3K/ZPLQSzwKLSpK3Q9KIwuFiCgApoJb9VyE6MD07BbOR25DObyuLhUlHK204SRSWC2YPhV5ePA
XQaltgU7fxsgCBykQxYOP5Q6bDXRSG759n8+4fERKtDvn2QROSjB9x5ZIUhjZncppsL2jsbIHXzG
cGIlFWk8KmljCxlQOi5ABJl8mc9SglQ/SBVp8+6UGtlgn2co4B44xEsK2UFu5cT21EKK+Xv8aZPJ
tQ0dYkMiMhM+sa1W8i1erdhirvDywE4xv3uGTKrN4HAEBTm6dND4VF5W+IuRDb+fcuriPZMK+5Fr
yNookgXG4MI6MT4e6OmhAsMspnNNKUiZakoKC9B6GWUbm+/ItzE7MYZnjkmFB1NyZ2xo5nZZ94JL
PQqfnFNFOppjce8GFPe5FWu8J6XxOWAZ2f8XY9g9Mw6ffQgj8VwcMxLUZqCiWZ6CJwbfm73YzW2+
b+wGqsGqIQGCY9lzXtIm9AaYGDkZibqs1XUPek7xIZQRJ0YY+j9J7Dzzw9YqE9IATRztSw2RcS6B
MaPi9bEgGN1bTaApko0qBpaWsR07qmrm5YavqGEZZTIxfQ50ssBO39QAQ45HXvCYXXxbzOM67NB7
QO2LKFoO7vaK9u1GRuYbitK0f3Tce7v+TYt4DBQa6OBO88TdIaSzOSKuVBfnYnfpsiTBPiL6JuX+
K0zaDUW4DZxr/iK6FojiQzMIPuUXZYLGpmGxmFQFYmjPYMAT9PzTxLPuZJt4/rr3F6XBF46FdEBC
pn112ZL5eYL95rH8naLhtfx3wfFEGXxWQr1EdSqh5XKtJRZDz0qKXf50EMOVjRPcfo3JidZCN0UT
dd+HT/enppg8AsuP/q/iWDJp2Om6+X2O/FsBQwtE9oHGnJl6/ZGLTGBHFBGTyJg2bydzR0me3k/f
LMpmZ8TApBCUvkccoqjvAE3AkKx5LgzWZ3JD2LhMp5EGoUdtKqrTSpuzHyQxn3dul1TmGik4dmu/
dghLFCKdlE8r3ALQHzPN90vpQUkt9FUe0izjKw22vvnlQZyFWQG+NvdXXNpB9kRg4u+rjsObD6l7
DPqTw6sz+zp26/QF/WloIoayYppVi65s8vCiCdvzY8yETWOvzmJqhq6uSMzmvDhK1R2Y3W5ZUPah
2fkJhyVW7SqDiZ7NYwU6HlWVQiLplkYfxt5Min5xZ2I+qv23yj79xK6ktkBtCMNQKjv+DEW7PZ3C
ZBdnsK3dN4lnR/ZqMZUxVr0zZqvVGdtXKGxF/TqQsU+bThj/meaQDjt91vrK/cH/krgiOek8wkta
6nziwOdqzMHHDEkRsCJJufbvlP4SFUIlAf65jWEHehwUyGnGoOB7ehdCzgrP6cpm9CeP9ZSt+BOC
CuQbkWqDJhsOAIktiQ8ZSRX/IercsqlDOby7mdz3A449V017XmH8CcCJqESMdZVVcByJpA518SnJ
BmlsBiHzktvt+sJaZusugVB/EWDX/KXsb+3CMIpKQrUvIJuvg+WJF3a7pjqvSRscnRz3imHh13Sq
Z+1asuM9LWQoiW8i2P4+Z1GUMBgvbL3e6Aw0wsZBuMGslzqctTdN9dQYaX2KBpk4sPoP2b4VHEQx
kSWEgQIjdnVKG2kvRt3Ud5B8MInqogVOXOB9I4Wus4aG26Nu6ibp/oSL2INhH8w6XcPXAcvgMzE4
3hRn2dWum6wPv61tZxLA1XZKz1xCJVt5YsshYyb4/l5erm2BPwj1ONfmfs1YuMejyuRKY0kY7wv8
pShqSWMkIpHnrD4q2mGq1M7pcCamgP/YLRm+A1w+gvKGYmHkEE0SRhlNQSntaOaxOKZ7f/UvEcxF
ace8v99EkYdzA+PXaFUCusrrNuA7Ufg2GkyWf3An825HGMG5BF7PVSktcuCnYD4weyiHzdGeFyeG
HStDfUlEikt+oBrVAExMHSTtm6mfueYqOOTU9REScA3MerUKW9IvDy1HbUcmulQ2d6nV8YzJNZyE
5hp3sFY8yfQRJu4WiSoidlEx4B0/4ROJKaUEXFkN37iGlqxbm2UzPe717ktiyOE3pC4VCDiATkYL
+X5Hi2tTRDhLp9JkX6YPcUddPXwW03DpzNAYXVmQxpxE3ovIEMwWatRnZ4KNJVwAlyv4jY6C/8Vh
Ku31JqFKKe567+U4NRASEs59mfnzXVW8fdXypk8n/YhqXz3sKKmaFXPvo3kQ+OuC9Yn3gRY1v+Hw
fh8dzgGv3091URkih2Zr1J8XVItGM0AwW+1u1wZGg64azFay0KJ+cQDOC+vQqNJNaX1gGM6+b9yd
7Dtl1oM4JxVMS5HvzjsEXWRE3ZXCvY9PQR2p+WpmLDnpXrJicpPY4cTCm7AGWhXfEIwD8o2ADMu9
CN8DyGxBhgXqqOdnpSyQymVCMAAN1rza34a7qwMnyi8jG6PiIxMu+tBUFROWlawH7+EK9F5Kp8y/
7wAsIJy65d4j5wRvExHQlfbYDnAkY9dKKF/vOyJ9v1JmrCanWxnKG/0aGMfydcsus8ofgmwg+5tY
CLGMw3vaneFhY1QgsoeCzE4cYHLXWgl3OOnDCL0GZOQuVU1MqPSO11V0PNN3SfRLMMXHkNy0cCJ1
HeVOXN6EHJwK/WdvR6YlMIfX1RHq/dw0qSqRPNXLCUGCt1MDk7H/6vYQdGqX24UHh6dCyVQZtdBj
yvJlEZZJ+6mD/NOoF2xMad6Mgw1u7YjN6y+dkfeOm8eEKTRiCTcW256JKtAbcoERFOfxYPul07RU
+qGAn/GoNdh7m3y3FHmYnpydwKnyUYCCqNxHUTYTYSpqlQ91QXiGNp+LwSUhPV/laJXS33ShHi2E
zI0rvEYJfA+elQQD8fHNBb/tp+2vo8ubdgzVfkzuZsx1LG3QRTHqtr+u02xe2HB/2xqWjcEPXngE
ycxdIhcadD4jlPKUqbscYX8o3ma7VqAGbzPpKgvFQZwqDZ3Sb0LSKZcMbu48c3aN0hLMTgz7JfZB
MC+iLyETsVcg6Gr9JS5vdrtmkU4nVILrbbAFmQ5EZXebRrAR/YENwZAthXlS82C/CzBCWqIG2aHM
f5RfPTdo2UtCi38rUvtnLVL5d0fFN9P/yHmwzXXd74N7bnkacTPI885T0mwgfTBXdd/vxuviPJFa
SoTa/S0Q1ewXoaCfHkCxdmsdOW7gai8iZQIUZacNoCmXkbOs43YIInIoQeuj3gR6CvE2TK8yt8CZ
uDRncN/OfrK5/Zid3xk1E63Rda/BL74M1LTdUcTvuC9oHgwHC45LbTG880zHVCQcDlaY2l2PNslX
3NZv91N7oowd8lcPeP40PWCCqM6Cn81ttWFaFdbQaJuFvGe61XM8bW8YHnmoD62mJseXGOVoFyd/
nx12uWyDlUkZJOzlm5q3T2CPjAJYa3gLmmPURRbqEFEyiVlEWsw949DqsJqh6hS6fBcIa+Py1bkD
gN3CvjwpLWYKMPa9Ko1M8TWELbEHsh1El7r7zluyhx1Wv4IDtaqi2yk0WgLNirYkuLXfEY8ANlsS
t8eqkrTVUYHN+Wp2ztJonXJKmrkQFALBEtleAjDLaRgw2BosQUL8wT708x6pyW3yqdIwWW3y5rmu
IODLIqk8pxpaViCVMovRd+mGawFhaPdkTVdUUQ0HD0WzSyMtPI+IDSpmG+WfTymGL1YksE8oxzsT
c//K6MHQiEYv29I6xsxC+xnVcJEh5sX+9OmVLYWaG0bhtaF8m3HCaNIGscVhn4qE12NIwxMWhIWw
Epdwk3TjG7iRoc+97gdnT1lCm77o2r+h/HTqVovD4dMYOkACrw3uNMWkZP49JLovMkI95eSY+aNh
cmOMqXRgREUzPvSDS/qLDGgtC9ZNTa8+Nuqj9okRtnTcuar2qa27PVGQVnwNHtsi1C/ATdA0tFsV
uFdYCci+GLAGJtAB83zUZTXHvniqY+kQaLkYE6O0vxnGt2Oydc9/iHFnoEr9Ej1Cy3E+/KJMWIDw
i+ddSLK4xKFGyQKfv8GLrbT0usRy4vShFQZFP9G0X/0ZWKSo4Qr+E2XBHSMnTZ5IeNyeItNjFF/s
AJYDpa7ikY3avcHsB7DrJJmFtLyDiRadyzbKTSwDTe6tVCj/ug4qjIlwUDXrXEwD7jBAxl55HnIr
fUtNS/yx/MGIqDCnv1fmAvvu+XgSKlI9po01pxyMu4bdrrmSbWOoBza/NuN88nifFeZN6ffuRiLa
k+3aEBU7dm1GR6A3ZU00KZuw4f6D4f8IixXdQqQmAlIuTTDn9+UYvLHzyGMw2rqNs+2/by217qLD
P6v00i7b39UCEx91tYV7aVzerTnLyAOJOo2yg3pqRY2DonNK2IqOlgZg+DZPQYnjB9QMw38kWe4u
mnvMDg9kQRA1fVdSbXRonA8ytYAHkdFfn9Tvvq2dcBMavic/f41Jjgvknj45Khyelih0rgGphbxJ
Ug+PabKe1U8Wj0RcScWhvo9VwvP4/KAUF9TIx88+u5zVACQ7urDYBavI1P0xKd0N6vfS/k9AvRbn
wrkZRCUDXoUDim3Qt9A1VEYDHVdcZHdVPcn31BfmsjVJD+bSC7ZcqfcJAZoKLLdjrIDOb4qxPIOy
eV2+hFdVlbVO9DogBxkLfZDAfTp2TjYZz9TL/Dps9iAq9GYmxOyKhgheXb8nnUaL5Y1Pk+R4oXJN
+gHpOr7fai/d+gl91ly28NHj0ZBfAbSJi553hpghLHyB6LK0xm313YL57Mh65XED6vEkKKF45O0w
xlcRuxvn3FVh1LjV0C3OEhAnCJIqoPNgEeFSMc85rkR5Omh1tqMhl+1EH0zlkF7DRO4UG79ZGYZ/
U7P+xb7RvcyT2hf2C7UYJyEl2aRxIiQiZyuer+MRXK07Vs3NwE//jlfUVXzLBTYwNrTtGS29MqzX
xsRzMLS/R/KHolWDEXuTJzTDYSS1wuK0sDXcF/KE10rHp7z+lfNMy30cNRCTWLh/60bQSyI/PXAU
C24m0PDUq10+7HwgXJYnaad0es6Sce55gItleWsL3w+l24zCiADL8/SWoRmV0JRGIUW0IrIa6DZm
ULB/lPDdTPxIvG/ALQl65crG+u4knrtNaNbKH3CIWDoUbd0b4v3zoaxXTiS0snciyqp5V1miHE7i
Wrm6MMNwbBVVqCQ5QmRMPJH6fPRbfTSNzOHVWhSEbDhqVySCio7EG5YNdZ3TgnD9arGwl6xgAnv6
YJWDirW0RfUyEKpFKHuq5FL/FqbvtI8RyuULAvQRXTot7IP4DBymuyjomVeymvBqjWS+QNwe5IYv
WVk5C1GB+J718yqn607FQ//zlqMm01rLG8fijEZnE5XfY+cS9S/Yb4Rf4jhkbW9MANp596TYCcJI
y4X9/ju4nVLFW+tLa+De7YGppQ4lh8rQ9MRpZ9USVHF++HYC72Q7HkNVYU0zT6cvRrfya63hHcLc
4YHkx5zOCr+7Sia8KTqor0X5uvRfLTpFEFiWxUrhuU2+2QEAW95JmD6Yt0KBFHWJPh9GRTuRlIYA
dfzL7TXYRDjn0bwsxMjuCIW8gSBPVllkQi8Xbo1rJ5jzR4EQDzE+QwRKSvlIQeywzNUpmtyRvnz+
02YPYLZfiuVWW8MT1dAS6YB89br8svRsHFP3ISpJrTI7IvUBs4gkeJHucfHwPJvk8vtmqqmtHC49
tWKNm/cuBHOVs4PyO1ySijyCmkFLMTRf62gOecFWNfd55I/Kbb9FIO67mHTkoUNIBtKJTst1uwqz
EPm7w8PpXT7Ihn4RLXBOziCjwE1HuV980A6OJ8bN+BhQtil5CvOIelhwTDkDvCH/O+ZfrjPzMtlI
8XceQoqHUXtcT/9PykKIsl/zq2pUHJdGAWgEbpXaUloEYzMC+3qEtHPQBM7KNL5OT0wGg17pnUe7
o8k6VhsIsRAaFG0KxdU3U9pSaQqQFQBbmlcu3rLuv8kJbIcI+hdRUjEUUh51dB4lXxjv1S9jAUJz
ugauHac2Xn+Wax0BRVlyylEsIbgAdvJMc+rd+0vMJ9VRlmfwysGOPArgj1J3K7h3+8lRDCjhEidq
Fdz9fnxgRRM148DIaz9rze7XU+JEKMyGF0+t20vfWAEn0cujvEL8AWoCsAbHagXl0aqi21mTG0cT
5Ozf6EYyXP/fYSDzBroxg8wHmdgoaJKBnPQqcIAcdKaVVjnBILDYmqCClCTa8dOQnOnxX16usLp3
xAKpNw0+pbqH6HhHSRuehJz+VQImRGa/pamy5MWSYP6Je4hUSp1q++QfRGhzWJ/sS5Xl+2grwqSW
qf8b4XR5p+7P/Ko+VSyaWW+WAQMADpbZfbxRvXcfqj9c/KGikpGoJufIlXIHwrDJwLWUa2qH+pr7
m5ZzNeCII/Bkxj3WtEfptcJUNMaoOMosq+So6iGX4FuYhtNn3YLMf6QU9Sz64MGR892fEai+OUII
BuZlnYglyte9yxiNM6HX0XSDLUJGdlyo9oT6dyVmeEEqtRUaQscGJyRI+6vC2iGpFDxSNCPpdMY7
AiuKCcSs22CPQghKUna8LhGPAoO1wGdHLi4fPT4xcoqZTMYxxh7519H5Uc+Bh/j7tRX8KB0ppR2H
IjAAMtAOMg0JraJgVLElPMabrHfg2JcJdEsmw1mHlZw7qRzyPMo1sdF0l+IxTMnSpnetR/PIOLJP
k17yOBw5jleJg0sPk98oYtrdz2L++JJ+FSwyPhFVANrvO6/HNtxN7XAQgYANBLmSj0z9XwU5dhyr
TqOrwj4VHcx/oWPzFf3coQiiLQQK+ZLQNdGazLs1v4hD1TBrk0Kzpq33oCMTJogOdaHJ5mtpsHz6
0eZI7Hry13gwHwP5FgAcgNPspXSpT8Kk1c10NeEIPkZpZqjnNENoHn7x3v4P0KqZwyvWQ/IgmZCY
6xALGUemKMTj/qNVj3HHw32/FGW4AqD6bbia/PiN1T+ifYRzd470W5REU7k1eWJ3TWk9yro62lnu
IybHvN18hw1HxjV6e/mbqAaxtvEiyj5w/8mAx6iFS+fCBr88oVz1boHNL3fARGhW1t4jgETls+/M
0kp70YkJlFKpFX5x/O/Od88ktB3lE0OotCDAbhYcOQT+rBmyiDKs3zvbb6RB2bXHj90p9Lv8WNMi
lKGoVP34M2h9NWTGP1W9QXi6LryT5lBxKQu/un2TEZy8D4xgQbaCvd7eGPu0vXaU/x9vJr18cH7t
SEY9XpwB5TIPzzzbLs1me/fuYNEyBl7VgbqviuhoI5xTZo8YNLON02BT0+Eh0Yz3ubLM7xztj3VP
T13Y0BCJsc0L6OLNjnU2BMnHbcalWcNDgqii5ZWwTcK3Q17VH1BEbqfYFjx+pRnfgPBYzpt35vb1
dDsx0ICxWF6BYc7WtzQji7RPtqOM+EzT7zDJEIxHnZAD/VIQ9T99coMksEABPBm0pl+K23Zm6MBT
wDoYuFgaO+a0b/suNctqyk9GAUhCkcri4qMqqBJi9ys3excYFwUizSEX8hEOjuc52eFPEolabqQr
KfVWdyKaSG/f59xaBKyfhuhBi0Spt4ogzopKOiASBVUHoerocHO8ZYB4bBClNjAskXUeIpAKouwO
pMpZ/u0gurAZHgCKuSnnHbrF/SrsdZ+LdX13IhpipGbG5giqCtRv42SoaJ6KsJq8B9McVVZ7Hgcj
/wmV2FTUilpqTegIt3UMLAs3w4CHlzHxZoFCklLWEkiOOW7BuxoSX9ZV+XojYtCtZ6EI6iw77/P4
2gnh07OfO0cX6e3I/cyXQDZOxMFVKVrWKKq14VD9H1QRJQK3wJv3vCmR/hA4cSfZss5W7+qMuwj4
2qJ1GiCquHZVUjlO+8ukGekLJAJllwKojvN+5CufR70oWpuxXsOU9Df9QPnRV2OKKmg6s62CF7AR
ZYwZ3s39IhFyhPpbm4XfDBfWqUOOPcfFoeDldpjWlYj+u6AGgiQYVRAs3L9EIwGv2iRKgBNDr0ar
1EACwXhdWk4fwfJkSQUYJQ8R47xGhX+Xn8NYD8ZA0hKz4B7cVYYK7g6OsUb3iDIgG4VSgvi6N6gS
jYJwLRnYXZYmvfKxTw0cm/Yqf5y8O3Rl413TEn1GnAdGxIfbzjY0q7uV5GqsqyTqtBnqzl2e8gvJ
KD9n0vxgqkNt/DiDTM46BKW/llD3/IhNP09W5Ng/ltUzzq1Djlkfv4MMnX+GX9jW3GJQkh+KeEWn
CyAF+0TqY/SEn/qABFvtqXO7NTGVELEmD6MMKS3OZfRDLBTVpG1/0KwnUmbHXdlokcIR82CkN/8e
dSLr2U7rdhKJ6oivr27ScQxGE+eT4TfMkqAFGyuMXExkqQf59YSNXbPUQlZvtfhM86+eRlQUK4o2
Z+/fji5tQ2fkdE1byFJ34hQyrVz7lz/dKzqyKP5pGVj6tGKqjj0IoCSno7ePetDk8ncLtz2dQR8F
Hif9ANLpurf7PQlTYDt9TOrH8IoAVwXkjVDXwywrF2QYW+tQfhXYd5vy7tl5A/S5M7iwPWYwyR7r
ReUl/d8PTC2K+76zp/w+BYjCfX0U0yDK5E9iG6nuk98Tee3SLBb2DwE7rwLEfJhDAVWjVQws6dT9
QsMvvWxC3mf7xSdremYKIQQUOx6qpV4IX+oeo+raDqNlSh7UGB5RQ5X5m8GnmAsEu5Xpy9NxgZTG
6MwS32YGXN2XhJhGh5FLiu32hQNBOX92uiJuPrBY/E5q7jDaRgsDJAS6kvfsx1fGU+RZEyI6sM1x
WO8e/w2RMZq+1skRb9kB/8lS4EyHcw6pju9np+u04U5FJTmP/WVOGZRqpulGLGJDFnhD8XyHuHo+
ZyqVzebEeFFngzgGGXfMm0Vhx6ekFefrBrWToncDAxWNZSEwzCwYBbsSfKxBNc/tq25H8euRkdZF
DiqQCX4JQYOYDCQOfdvjYVk0DFWy0bw6BRhf8NyFxVyKbl0EkXLe8eLDZvhidtcwHlPACPRH4a4K
PDoidp7WC59Iuh8ao+8+YEDvMXTf4svJS+2P4GXfEMPTcAta6ovK0RX7hIukX2RGrR3mFYPg08Pd
XrpoQioYgubV3vcT9wzKJhhaTwK1kBdxRgf03vNuCbG+UCThdJmVsaEAX+YAKNZuqfcYfZ0wrp1b
2FqXh4Z2pYdXe0o06hOa4ofDsv/U1oAdr78PRIOTM29q3KGgKxgxpbmpHeqHv28oD3gu4gvXF9Oe
393ZRYlGqp+LLu8kyvQgcxTooA+aciGOZzikzEJ+HquMRuLqy3GYosLbncxHNGGH2JeGxbn1fPJw
vofa8dE9oAL+hGbk6XMUT6efC9a/KqyQ3iogPHyBOAnYE0j6aGlrVmKbZ7CEhRSgxZwteVdtOAHT
JL1xM2uZvVzolyzqOrnRPqlWFvarerrtEbfIspzXaAYXMSJhde2d55j3lTCE6k5n8JD9rkKMDdAI
Bb2KrFVWDKuDYy7Ap+FiuVJHdce4ifrCjllYUISopyL+I1tlUu2RrFxpUZ/PMIRlWrvpYkSVneG7
oXirp14ohpg3LmKAJC8M4Ive/dem8w1L5DlAP2KPsWgxiq5SdZp4P4rQIuWbG2ANSaHvt2A5QXTa
i1L4iVTXlUksWEizmzRzDnEANylAPF8re0kygKqoJDqUK0SUlKBOywvKBW2NO68K/ZvO5HM0drWn
EEwrJthGWf1BEhEH6TANauCvTLLaKywbR0eWJqPjIYmKc7ikD1HOIdL5v9rEuIVEGOd4nIMvu5uP
dqQd9Vy01ejzaNY8W8O59IuCx1IG1EIY3zXIG6LwCLplCV4JrJYATDkivJ9CYnqrtjMLxSBDJ0T7
8vgNJaLVP4KqqbYIDxU1hVodfqwezEiVTB8LgT9yhLDo7P+4NKfGPPukjf8AltXXdGKiuTWFmCdT
fehHN8hP5w6slxuT//TAp8Lh5awTC6hltPseX4RZ9az6NkYEpaGKOPAUXFGNltYS2ADmzfBW/XA5
Y0AdkLqs6QFPaSVRxROWGeWGxSm5p7PZO2he3N53gWrrZ7dGLmV4yMW4sbxYgDWPL6r2lj8j6UwM
73Yvumlri2GyYY0sSufFHJK6slFA10AtppZn7JXqpzwkZNzsemBLjCTrvbAK6UrRJv7483V1X1v3
9C/n1QD4JjUVECnY/tlDWFtGgAihO3+wD6lehV/QwjtU0hKr46i8KDtqDqwPTDDb/Z6gODsaYeRy
ue41g9wnbXuhXDVEICF/vqIM0ClW7mJLxuzrNHTRt0JM3jc8BPs/u4b9+Z6O6ayBNAemK6eVQOVb
11TGAk5F5AjymYyVtxE5lzYGoJPAAECB4OAoJ75hjQkovJqeHMdHV83CS0EewZSIJK+EeiiSsvIR
SHTrRFa2/pxYJY+3YJdFNjNmA0bChdFNpDHwlq+Fw0OhJzCQtCNfZuRNMpAA+Le1MFw3bpjZ8Ev3
Q9iDvOTxIk8ZDVUihWuYsAm5dnkVevDj9UJq6Muz6W0oPQNYVCZN5CCXZ70fKV46yscuVnhbi4Si
3fsr9iM1Phh9IXfviEyY2L+SZMktKepst0JQ+AfEiRDIDNT7dnZSpsRFDFsFBmkn7tJNxxY320Vf
/fcunkIqvQ6ZAdoIQJ+KU3h09au7Y07fxmbXqtBmRBWMoSbdwloEl9swM9pYFxpk7/jCCTP3779U
Jnb9d1t0StLS18np6SGzlxtSxcVlLWl09KM1QxV1voN3WnGjQh/2Up9N283qQTMu8uToY4z61DFe
8QbJgjeN/dmqAQUqPKV11H060aSB2aIkkfZMpBa3zmQWVR8AqO0gzdvXJZZiUxcCqPunOELaLR/m
dDRZTrXPeiu8Ldih0GNs9nePg6OM/Yz9O70KIxO1oURssNK6x7SAeCXMpHQTsZw3t94dujVloYq9
x1HkqB3VxRQK5PnuQiZkrzFpbyehzz/olClRCasqlYWKW6EQevgaps1yBPBUFd+t/6GZ1Nya473P
HyW1xYshYbiGyw8r4VqL2A+saIjeEyLGF2J+JhWEfA+KmcusstCM9XRNrgvaZBgfZML/frwcHoqm
PROdney940WNLmOI0x4oyLAmAItoo272FaVkSf2Zoy4hhQVuaUY8oQjB0iKoFkkB5IAXQNGLyQ8R
OfOaWu8EvXTSAF2LptgV/Aaqy3PsF1Ky4QjCc6NL+WvvVC69NyTCrPD9huEoNjts/Kf0WmO19wud
SmjZ08HfXJZl4viqyO/TBBKV8qpGIqGm9h5inGLph3lCtLSzL9voW+gI3uVCMDzuGh6woBK30esy
F9+oy21K+ncotIHJyFAEOV9HcZusMmy9qCSJ3m+6d1OmoPa3/3Uf1f+FbzABwfMc3vA0F6SzRrwg
sJGPoaM73OrjY3NpelfeMfHXzNV4sSOl5fOciHxeZhIvfUb6NvlsMae0hHXk6vDbuKCqlKcxhisB
BqfEkukX9X7rdr2hP+RZiK1yJVz8s5cBUxhyeKBuacKkQBdOtctSoGbnoyNI/bdGkUHYkF1uNn+2
oi75lxw98FAhwrAN4UuJsXh6gZ0Hc4Na8amwjxzB3fhIYgvaH9Gv2wShIjgGG7AUrWpgEpgW0/X/
qbS1b0cls75RG98sQ/m44HFgoL4DQz2sbx0gkaJnYSgNAUHNrKlrwhcFMiFvVJsGslUCtDrZ6DWk
nIxpiyaOfjn+fv6NqMhX4OgLxyF6GLazZTty0xXAlQd0mYswaoeJitJsFStd1+F6hlWzjMmAgD5T
4Uph0PAkturB5kLAvfAbfeQVGbwhIdOXhLq0DUT9eQQBeCPwMXFoUeOAfWJ3Gs58IW2UKUYPqoRT
3Pnsv8LfsDAsXAAmsyGCNY/3m7e4dylWgtIj+HcIRd+PzM2/qunGYSKOAh7k8SbZIq7c9LM3olZb
Pfpg5lS0QDRpp/zmLuC8WO+n0gTR371u6ebvAS0CpqCZXzpZI1y/YtDiVBJjD+pGNCddGfqTHgcb
HBE60rkyICB1yChJlKfMTgOBGERItpOaMHHjNzIt6YKBb+EW4TZDaIVVnO3uTzMsk6kfCKyNJzzH
4dLCuIeXnuoy6ltaw7vrYAlryBcMYBNBvmGOMCWn7tQ7xxfjuP+KdImEp0gOvz+2NIsAxXsCYyd4
6XiR+eU7eYHovRhED4b/1/s4BAypO0s4Xop2rKPHuhHRSHk58p/s0bSWNZaSoUt5T30LYXG8YgkT
rEG4y1hbEZFdAGeW3pliBKdoe2YrVip9+YR/P3ucAbbiNGCClsUgk84bJfMyZYsXQOzCq/E+JBkm
7CVk5fawWrxfxP0g02YGw3Xnt+1Ld9pwZbc+HiE1Ptc3PHRFS6GCiIrmZKdcFFNCnqvgAqZTeUFF
FbZwP6csnlCQwWSlWxcuZBmCzJ0wWpUpnHCSWyQJEZ9IPO7vq9kCJOSokSHOLZTANrlrO/TzY1eM
OFd2C/c66DkpnGSjxNlJI7ol6ESd2/17yfGoV93lw1DrZiE5lrmDL6pOI9YgkiLXD4Nrjr55s2Ac
tTseb/Qt3TtDutI1sUF6YJDim0w+nUzhx3lz9gQBRDZBGSMIrTvokXVyEFxsg0yfkFaPYLlnz2wf
v4jNaZgikB8yB1H129PQFFaZMhTjCQIpuh4kgSf97LWl37k+fOjLJjx0QdaNKt+PGoxnk+fcEkIF
3eO4JfReWVXD/KP9UCRVtyp/lIqAOj/uLcMU2JvqaqfGNBBrwKUSRWFnLfrxKHkj2Msn5DBYsQF4
nOW+oFjsV/zUs9J8WbvpxQnM7jRlzdrQKkup9m9Ob4FUfVU9WVlBvQoDrR0mmW7PKF6lg0Faa1yx
GOfo4ZrGrBemJ/z6yqhL6zaklbFik8XFHosjG/mgojiG8HEvMwLVJewcPec+q0/d3ucArvdx0ZBO
8Lg7cMXWF00Q4BfVnqJIrzF6Te8HSMPRrIB5kq5rga99g38tRAcK3sH2d6LYHIN7xH0JGT3zLyyf
3YxrWzYND/rC4lMMDsIsM6ZPZ2YEYIXFPdaO8NGUxfiocDMMjaagCcrvV+eTyIY2cBm2dVNGduHC
TbuV1kAbrc05PjoQl2n/Jk2b0mD2Y37Vbr+BmFoImnUXuK6WEkPj4nPnAp4dJnUek5uRlnLuVXW5
wf0q2rfy0Lg4C+vyMUiAhtz5/0ZI2dLl58UO4uINleGUuImYgXWSOF51ye5mWS3TZi49q6s8qp/+
Vj6fxELj4SHK7IO2uEWlIzgYK+7+ByiX0D2XVSFlTtzUSP0IjVusNLdn0rE4cvbFhRFDMTwZz8ni
acI/N/XvHTIe4AuCgpRikTmLflKOJw9uxG0TnU3pO4WxlWDFe1lQT/08zkCz+Av+X2HW1ePhW4Ts
W1i+dBUYu7aZdnd+Eqj82+VM+PAEz6BpXSaf8Krp8psUhJtNyXVFZ7/hJKJJV6dlbk+AYCaF0chM
rKnfHsTkpGaYm+NhQlSnfWyXgDbZuDuUn01L+Lec1NMqrQXEb/Rd6kLqr4bmAp/pz7uE56MOhDLn
ImkVeQEjhMeQXDrADXGqnGMZWaEujVK8d3VaqLxdbhRDeLLb92JUgZ0tmw0tWGkWdG5YSI/Z2uMO
EQ+qFM+b70B/gx9cDkCWk5Rk6sAscgW/11yBybeN8pz2cFAwpTqFkGWcolVHBdJTavXn+zKB/kfM
4YaguamMrGdDQKK/Zu3V2/5ySYyYesQLe/+y9wJkHKQhWxcSVJMz95pG5/6AsKpKLCak/YitmIq0
K2k0T/YVER6/AfmzNuKE79apGkNMpPjDmUol1d3i0KcsuHDXd8vscQSES8NrVL3b2DMHT/eV5mkR
0OQRhoquvDspf8+W2sifgmXBAdVpV4fRshUcwqLVvZmGm7mVeuHFGLmc4gL3k4+vXP5BUDtiiZef
GzVPNfgNx0K5KOvhhQW3fVVUVA9E1sLpEeVrUk+kW0FAD0Nf8raJKqcaaB75Z1HCTPDMBBkl7NzT
nClKsEFQci4Qsfci6g9abgS68GBHtOSsc02olueFw7wWC106YHDQXClH8z9I0/MoI/u7dGpnicqS
bDeHpI3coIi/3RGeFWrQJSLIk2pLtb6vQF6qQz9AmRnjf/vEscimM1pId6ftC0Xn28rrfV5xJIA7
1YGYupNRK7ChCWZrtx0B/Y+W3Ezov4qAOGuEFFTunV5tyj4eOeoRqeQ1S0QCIgZSGAGSGhIofPv7
D2R17huS1NHkwxD2Jbm0cLxEDxy5CRJq3s30xTQrXRgXiRfw8YvqKCzDNKV9XXl5Fe2g6hAawXl3
EcUIpksoLL07qbpypLPXUU4uSYNxv7pEAiLT7RIWnzq7FFM4c27aovvfzgRTtbNm3oeveg7ddMuj
UhR/iyasKKEdBdtN6ymfITlH/JsRFSqdBp8gt13kofZHCdBi6NHVmTMpFYADctnb1PS5LlAvwr4j
CdxwUA2K7iL9hATUMkVEA7Nr2um38U3Tcc0OgSBWzdo51zOrcdwaVSFgohDYZtC8Q/pr0m+ux9C3
hU/sF654oahFqdf8dIiZve2VuT2Er7kBMJkb3zJKFpT9vLq9mN1mp67Vp/P9R7TV7raIJ+o/i49z
DRiXIznIF3aHys9Q9kFDj/81Rcp/+jLgOgX13lIgf+jSUNfYLOpGnD4JF/W1u1jLBT90KMeeFXAq
FLhCmWGXHnJcDTthfVCPggpdnLyf30J77u8uThbaUK7j+XjIzeUVjTAxnm2MwiktyUMlkBXurRzt
2p+RxI0A7iuDFt3pZOohhOlLB9iAedMw7DMs2irxvclPpYDu6Ay50RCTRI+Jyolzc1yUj8HwAfzi
0p5pp9pdgnGLKQaY1YdRuVob1a82To0JsC7pmR0UvLJEaCvP0fKQpFU3cWe2K75/OxhfhgrNdZxs
G1czULEFk5+2YM+v5pmdtKNFhQqrpcDbAqjq/VRThZNLLzv6HemyS5g6N/IqyM4ICLRmcWSOxEWw
pWMDQidWEBSuwxZtH7zXg8WCyaTQ7P26RzRTz8I7RMBW/AchbYt1CiTnTsSVNrT8aUlwd8COYoZT
qhmcYVTN2VGxw5d4992dzRsQ2u3FYJizOVli+Kj6OCUUgZzwOJxrtOoY3FwUS8CmH/DRE60iiSn4
fz5VxDx2cznHldeCVwfbgtSgPDrUBwDneJBmgnuaaxbdfABEwMbc+Xja7EilXg5qfYlsjxqrg6VX
AMqiyxkefO96B5QJo7YtvpNOUx7GAXS0f3i7Ba93aMwpiJqGuTEPj3AwyolO1Lg3eHcHBTVCq1MB
Vq8MfsDa2DCigk9qKQ/nRwtBr/LrWCRXzKnotR+6TVCVEJLJsBSyYk1U1yIsGlQpkUKRHnnTdWOt
s6Q/BjfMxvXf1HbvWXGAWdIdUU/m/rJvW3MDVomMJri6LX4+uHnDc5kchG/G6IQdtRzZoyInbDW0
CFnYqS/Q5j9+IrqSLe+N3Gm8NXClx74as49A3DKc4+oqLUSZBhiYIRCK+Xee1Oh1O3+8z6A1nfvT
ZUe0fpbxoI+0LOBMOkW487RPlAPyCsjHnDSFnXnuXEt3N/qN2x4Tepkxbw5/EWb6AI65WQVFX0ui
2fFpgwkG58LgPezKdTR2qqlipIsl9xzNOofYcBdHrr0bNiy30MV24BYcGOg5pEpNUo8kRiUKKW0f
9xuVWyfXo5/qrHhRNie4PX+/WOp/lQkcDqg6hIwWUWjrQ6ZG2K3pYdmAcg58APUlLO7LKrEtJCIK
BKqnS5VbZoz74CVb8EoOyAlTsX/hipvZNjA5gBAbgfCdZyX0FOVpqVDdz/CJym2nuAtDEFfmcK3L
SqcZxQEWP/wgG3UwIO8rwKVAJDHbgyrmOO2ivmxQpW/QSy+m/UQD/U0nhzPdpo+CJ7uBV1Vn9L88
1KU2nmu2l4pg9E575sucFosF5mBd+qDsCQ7CRYl6s/npCsOqh5CReNvM5jMtlF1Oodfgo4ExyaHn
7/b9rMPlffGjzi4IA0ygnOFUyffpnEtFCkSXBayLSx3d9fLXw5DQKQQc+sSt9eLbpZ2Fzc0jC0Ji
ZdHTTpLeUy/Vo+iwX7MkQOae+xQZkqUTboqOtr3EpklTQ4MqMNqKZYCnSwjaV0F4W9kfDQSjcIRo
accbdtlWEMcbRaeL1E0qLQ8JbrE78U6m0BjiZN7rRni9wbH+Qki8yJ0kkQ2Bs4nLauID/lLioTrj
IUY1FW4lSGjovj8nAjaYa+bGq1HdXNNbBUyrKUiTW111Nq9oEsFM92HLZgNAYa8wmDMMa4sS9FAA
990Dj08dLCxU4gAIwX8TSciFdKpwUTC4emSlJP8BCk2iFJPgsMSwFr3DGKfynCJWoSiUzWw2ohJ7
sZePpYstSg82ugYPaTKKegyw+mOSwS7REjUjQqdUxjuZJcNngAF4bA1kSo4EynBLQFlRXu9zsaiJ
rmjyOonbK2LbOnfDs+eUUoviHQRY/mTYgwf2Jm9DDXaiyrY7Tg0Ui7ZSV8Ks8j5fOsVlZ2iYY9YA
oTbMmebaINZXNqAKf3OfH4+3UFfCyLQ5m5qNe1H6TlXKWofg2SnHU73buGBNuRL3BO1P32TH4Td4
qL5cM2EEfTxDWz9HLw+2PSiFstbFJOVgro0YDoqSZ/50H7WQRMSSjFNIqGLbGbWlk7/3zCiy20nW
QQfXMAgShgYczdzysNgWstrSGKjsbJM9dP2tKytx46KLrsQ+VKFa0/NabPfTx/GzK7UZD2RAkKwo
+syRwj4t+XQFcwkYIuucT0vuv4cX8GHgFUYxdxMH5cyOp1rl/wKOcqP0uI3K0fv8TiMKe12QDY7/
BsdhZXDnvUpcXUpILFTb4o+C83pMDK9QI1zJRp7EZ7MsyFvrN1VwQRtSdIS/ud34UafKXhP+hsxO
hsd+TGM2bsFYSZ7t9Onu4Mw0l57/+tfpXE6YH1YJ0/Zi3eRsKop/B0T0xYGUUYD7RvaMXCYrMoMZ
7kJhHD6kZHix/10QfHlJ+mAI1e8F+7tERWv45iYPYWlICh0AlSq/F2d8F7qjQS5ED+ZJIwiRrMFW
Csm7jEvxi2hoUKQoD9LUrVOzItIGSFldz+Td1WwaKkvlap8ueq6s5gIEklnvW4DBJMwOD3hmiNf1
nZU5kugybddEUFHP/N1J/ArFKgxJsIsfNPwxmQaCUNU9KpwZ5sXUoEZRSTQ+aui42oBOwlL9YL1W
BEAvEuPCxEgw2iUH7CQ1zC1xiQb0pGNJVxQGB7V9qbhak1JjFpHtqNVCurSSkF0UsBTNUG0KD8bY
L+blbjz4shwr5hJ1XyCwJD5Pl7us3qP1zOuvjNZpSrIto0IhmMtq3X06SmQY6w/04re/baOllBAK
PV/YM4ZjUNHjq2yOYEli9aMEmcxeRnk1j9Fg1aSq/0ppIyIwws9YMiJmAzYXp/rhckp8f7oCpkq8
LspddCPjxs4gZ5wdAYT7B971haS5BOVTC7aeEgilhb6blx658ZM1bK2DgAx8rP32TggOZHooGgba
HNqRibx3ieNE6WMwms5jDCjQe+l3o4lOPGJHy/TSXw6gW1BxT0sqY+TnORJJLnuyJmD0+0RZ5XnS
qAcE+9PdOwzYVHfcPc1vKEqBeHGVxQYzUJOgu3AfslSZRZvZUy8w672GoUEfT3uFzCy0TKSBJjaj
fU/eGaN8Gl5duGrADNA13DSFTUQP5sT/IrPBFowjr5vyZh8de211i2g30n2uQ/8NI4x4hIGb1Iii
VXReEaGao9HJPPRlpeW9mFDonZKf89FUPawV/UyKx/C4dhbtHwmK9oceGhFNwC2IEHhUaVCjwDeA
Hw08XOHWdZuBUZMeB1gAIAENoG4QA3sQ2gLpkgpvaQ8u5zPR9OkTvzHGHMUbpTKN8YOZcMuZedo8
HcHA5Mglpx1DcTnBXY1Smw2HH5oeRJvzHNtgjd7KvQf1N2XZYWjqJ4UTO0w0pUtVW27Gw+TA35HX
Hz3N5xW44VMd+cWpqKYu1Fq8wf5ENgReaiC1kmmLyDI+THiH0PfojCl9yuixWyViHEtIhGJZaMY9
Wh+tVynp2pJExfbv0ca+23fd7Qgk9wyu1RZEwMsfbaH4EFAbympQ7ev6A7ZeQBVdFENVCHUdwgQT
AT8rMrS7CX48OPEXM6Rrezk80B/mtYZjqBZKCCxi+y6YiEFiqQz0+0ua8jPeFbUxOspi9oEWuJhb
AxUUsFtOEYxKo0tmonu2acDl1JprSLtS84pgpVGSgpruiMzeedK6hb7hV5ubs/9LQrVNCH5deDf1
ytjOVtfI97lu3iFASgGGJwwsURmAqTPKnuZ44YEB7vIC1bZ2PrvNzX9pJ6cLPd/xn59O4rg4ElIu
NJcsurqOZhLNYgWneF3vGtAUl9FpQ2XyN9oNjUGcqbjTvPB5Xpy8h3iBAsDVCdu5fBGPYczBjVgS
Jv9lw9K5VrWONxxPHqp5jBolSIhm3KOMX91eXwaQZHIFy6JMocN55r2tw59gdBSe+PnaFXN1X6qo
6NnNL9f5NVlwWS+tiL1GivCVuyc9T5FCRZNyvqhozaIWlqFBYr+NFcnpdYJoMOQ3g0p7U4SFJC1P
16I0iE0Qrlz78u7OLjz23aThWfLCYLwtod5nCqdKLY+a+v6lKVpsQWQgIMkPpQWdxmYGtOiIv3VE
YIDRUJxak/8D9WVs+HFsTtMjBu6apAhWhxhvanynm9aW4TvU7i26cA7WSp/vGruc55uuZtSPchec
Ke7c6w8bUr9HqLduaTyioog5nWqhcwogTcQ7UPg7v97j/hG7DnsCRtoyn5g+1CY8MI653CgQ8gd+
4LPdyllcOkZpI+BqgrPzq3oHNZeNSSN0bzDcCxwV2VLwGvjHVktzU8Q/yfXLCsOJplpBsmpfS6ma
61V7BrjPqBb8+mqCr5YbwK8dJjRRqDiuWtyLVO8jrTLOqfE1rrW8RthJJtjzlFMi1BQqFs4ANtpt
m2YJQC+B+BiCLxyiV6Z9r0RiIYrkucC2/fg4Y8ut1wqX+2hkVPX6MZGcr2b5NE9BHIRpOeG1P+Tq
8BBffzpgQE4RX1VdQWVQfVeHEmChnG8f9XBzHkg2VyNXpnjkHU3nDEEMxqJBMDKKoMXxVT3jT1gs
9N1t3HXRqCNPmwNExZOdTLcg414M/fchcgHNactS80qjX6z/1g5jcQd9FVt9p5EomqJIBOOjnTeI
D73XpKpwkq9Le2xvgishCb1z8KTY2HPLIlJ98QntBkL1F6XtkTJgQLpEAIqlXqgKcocGMGubZJQj
WssOMqbMlQPwC4/rholjS9QOYYlG1WfQAzyKIP4XcbmbI2SsLdWJ31a6ZdhgATZrjMhIOrf5Qahr
eaCrg71fGzirU4OLzeXu+pevmNk4aN6vj81F7QVPFoMq3Iz6v9rQmokv0Mjb7Kr6pnbU7F3d3bgK
ndTFLi6o5qH68UrwGzKhiSvVO20hwX5fNEKglZsnLHwCy0ugCPsFZC8bHzBlOtmUnfoABmuG2NZb
qCtUTKglNuTVvsRvIKNf/DYinpmjCPpDUhrc05iolyMZdloW/YiqLbi8go5oZQh6Ilof2eKVHJaY
6H/lns1rC4mxkjTER28pJseBI/BdRs53RK3jtIZ1R77ZwfrcP1JuDyIHWBREK7OvLFhODr2I2mtx
Lm1E12oikmcCyWxppI5vz1x1Cuv0YRI6L/cF0Z5vSFTcAxl8aK5FXiik/angkjXWfvYSQPuB2GUL
vwmozSJgwMCOUqBQaYzNEHQltvA1DJ0PxquBaQQ311oepRJSUoXZAZ/q6IHqZ65hDwNt9VfLvAj8
YfHMeBj8y91uqC6LGbwxeKPd1P+YNbQJPZULU22qyWO+pYZjFFCpl9UPwUoG6843o/Mli3yvcANM
/YhrFesfWgR5FPrxCWlaP9w0kPUHh/PoeAQx5L0r5HLOtNO4qa7IDEiyyLpGbXgRrj+KvmT57H3M
cL2NDPgMw57xsg25dN/nI3Q4RpB6ltkk0jCTf+qq4J+7LYBgW1C0WPSc+CuczGsI0BSXwUTVG+nk
HspsKJ0iVAj9luNVdBOZ2ABp2Wy7pJj5CYrOhfVzg+cPuP0+1Ee+ZJw905582adaYpV5iIIeb5nj
+/TVxz8aqC45pzeE2wNom4x5+6rACJ+sdBQ/2U7hUhvnW1vMoIfHjWun3vF3JWr1iJwgkBbheke4
V/cX0Pz0oUn/aklxMmsWqc8aWgSYqoxhjkgADYxHVLiZOGoFgGGGoEn/4TigCTl+sHL2oaH+MIJI
AK+MWjtBkLWwZHuJpxHGT8YQTSbKyaTWOK7ttttCt8y82LT3WFFUI6z2oSyqGG4jD1Zsp9iCEMma
0EJim3WNls1t9EDT6ZQFpPPRgnjj4xCVDOv0/gCIpFgzqTV8ZMfAJ3LwejmUQt7oLyvm52sSchBG
uH0c9lKXyNktVVe86gC9utRdl3k0RufcWaSQzrIkeA8NwhosFA/hA2B8Go6zmAk5C/A318xfxms9
Pt3OsrQAAlqg2fCJlXbGqkYpdPj6Fr/YfQnxbubmZ0Notmt9wBe1ulmSsmks2ZlumdiaMByToWRH
HvbXAhlR05Jm7P/zzQfgQTeQ3A3WmPUVYaDk/3xnjiUX+F49gA+drz/C9rXMoXsLkfktYoLBB8Yq
koiR8CgUPE9qGMbSKvKN9aISRNnqChZmDTkkH8HBYgcs3iPEcjOi+d49Vjxt5FCkT540UjKBI2H8
M/OT4WeOKk+hTMelscXSe5KYMm9GvDqmqTVclwMg7klIxlLrlQsQ24Oq2lVpz/6yA3g3k664yRpc
4BxZkxMbQjoKZV4lDuAQozwGv++zIq6m84ct74cvmEc/yY1800dIZ4LdSLb3ZIrjVBxcas7A+RSV
uzmb1wPxoh33JfFLU+jAW236QnozQUOODjzkQtKNKzesSv/ti0sKdy5aMFc4yLjtHYa/MZR97VFR
zqp5FaQ+3jhVLNVfItMwY/bBl1hm8lXCgf0QRZSOzMoftk8bQeSF/I5RGLhuxyxMEfBY5cvYiseN
tW/a2Nb5CegM3u8tJWxqlwA+oZnyRLbuYv962G6XmI46iBdPV2BpSN6nFh8QXT9SqYV/k2QDRuOq
CHrAXvyy+9/XnPo4E6NQ/gWFZH27kTnD6Z+6gPzKPsmwm4Eo6hOPZkikUpli3z2QBzvGh/CAZGWB
0V7yVvaXxbRVZj6hn/95G02Rt8IZMRkv3pMFV1vmU/I4OqUewq93fWxIUAehobiabeZhBvB+tI8m
uM05knLakF/KvOyMx/fo/VOC4A72ugOGMQZ7i7NnIO1+zz4xA3mk3grUDxbk77RPTjw24VtWy7hL
XkH68FEgWZcubCUkA978ZbH2qk/vTzD8sArUJh8VqvG8nxCO3EJNydxveOT7i0vqEA6yrwtF6SHj
T3A321aLKuvbxaFkWe0gbQXFpId5gm4zIdwsjW14fqgacFWKIjneCHCoT40ilFlybXHRgYTHcAMn
B0XxWOhJrlG+hqmhuek9mbF6yrchKD1cj6+CJjSvqxsEtKEn2mBnjjBgHWsOgS84OCvo4+3/syVw
aUIkFq9xRUx/fhetnLwYnNi0/G3BmsoEk+utbEsEEO5Cj5TovWnXYTKos281H3KHy6WODdyipMKV
LcARgr5p9Lzxe/64BZ6FRGkDQcYQOBsApQ1cG6lKTSFerGZctZqLEad9lNj4oujbEZ4IaQNFfZo+
L4kwcKWt/Oda2Mb4aeFP/LjrqpFlmjiYwHlc+xAyTdRue81AkgvpZXF5weYBu5C49Ua3Mv1/cxNV
r+0hSt8QKhM1qWZn4pS5ghNC1+jhyFkI7oKkrBtKBu+kJ+Y/yNveFADj4uKdDEfRagooWLZOdgsZ
IrK4E/ioAWRNwBt7p3UxMUhtMlxtPW6+S45BPJ0qe8J3hD50w32BpZ6do69Fwi55uS+1gZpwumd3
qMcw341n4bPGcQRmGHy4bV3W4eLv6w1cl2EBnCVnBy7grycsQrgc4pa55ZTexvsMcOL5O2MXKRf/
KmEPjHKM+rpYcw/kIL0nXlHKnEuy+SckitGuSxd1lb4CjlZ1nPUIhoFSI/bpNpU+pGed3sB3mN+B
nCuqLSHItlZmQEsPTI8wEhu5RtTLeZJHK1gfqVi4S1gnb0LqWfhmplOYD/eML732tMU9io/IFad1
VX87+aancvphRZSI1CV2+ujNByJJAqypZWyr00aMqdvdw5NeBFEV9YDBRLnZlpY8LNMpo8384tmb
iU9qjekiW4o/G4/WMIHXA7q15Bx/Q0m/5K8inkHQSnrHTnRr8/+ADWo9Nl5GuDeyCP+lfMaadDhX
pOJHTtAIwL4RUTBMbrVAyWHhgdax+2wde17C5yVQZO66bB7r4dWozKD0IFkSfwMApcSp/OpeNqPO
QX3Jd63yhniHJyxyj7lvZTBezlNXpqgP4QuuWBzOwn/3xzTi9zp5fhepS8xrHpd9Pkl7XOiVWLE1
/Lo3pdxI0mWrjfc/lnQrhBDMZFqDEIIT3VLJVkgY+A5jWCPaPH1DSCdWiNH3dsiDVLgj2uH/5fVf
TzLmAgoImVJIe7KWrL5mZi4CTOZbz2urzFXXilXu9NYheSzxRkclSFgTVgyn5Z8UFDNhBtcmpgou
ON4JYCh3Rf/usdu8cPEThrKBUnTzBBAtVeOgjy6DYPmyyaNs0D200i1TvTZyOMg0bFA1GgXxLjXd
rGSGuf2TaN4uCfN6NDDi2Dclg9fcA9dBkKeZW1cQya+m1w9+Y7tx73uFYoTLWkqeZSsVHYUI5Qf5
qfExHIVEY0i86I1LyF7QzK8TPXtSnyGi6am8nThJJEMUXLJmtplQwa2PTRxW7hOQkoNN6Ap5u5/G
GO27ufCEYKzGYJN7oi2aaOYxJe/Fq1ecjvUx9Qqny0jUJ8yfHUhHfODjNlPx+Y684j8q3emHj4rO
n+3Uxu7tdIwsSKZHU1UbbcNWGQwpnZ5pMgJWmAsKOnnCWKdWQ8CJrpEsftNQcVvULl8wL0D5nx7U
p/6utW4AzAKkt60R9WhO9aGtW6acV9tIxWlQhzNHPcp4MFPoLJpEwIBvIqng9PeUEStKXheIpOte
dCQFmdNgS1BQsRTDSJxpqFGNhvWuHiT35i3WRxyD2ZjeJlM3eXGtGFGRSZ4ak45Pn8wII0WJ3+/K
vu08Ft9tjHFV9jzREjQZxCx5K8EHTvoQ3tQx58qWLtFH1muXxLzVUKeanuVCwVPORFAyGQGFlRoR
2fT9vnxQc4BF67JHMRmc9SO03TeJ1etwl23Y5GnI3KgX/rqwzsyWjFuWNFDH9dV0SZ9UhodAEdV9
WVJpdG6unxJlxbyPH/F7ldDe4sjAtf5NW+yst86m6ZongbutvBgewK+0BOmiz2x0PPSid/UiYUZr
PqjljXQe91ggWH2g3xTx1mpR/LH+opuXPvIlrX1W580EVsEWzfqpIP8MgFRi9yNmzh6HCFHb47gN
ywqXmjC1NlntWnFMW8qsddAADfuZ2PKxkaQWf2N6xjpfwEB5MgeEO906B35l//a/QFOz2RkYPXcT
hpGeOqsNpWkC1JA+XR/yyU0po59rqYBysfHjs1s6AJDgSiieNt7N7PX9Cri08iEkop60hjBVaexH
pmvYaVg39zpyd4Tm7c7Iy3fWdxmeupr9uko6knEwY1bm0XP4iMsYZb9gASQyPHap+RcQ4PvXW/cu
iPcd54GY7q9SZEzx4FWFslVOcpZKG9w8s+aDaortvl0gqlzz3Vaq7pfnQ5emzOHc+ZOfTxF8d1AX
QTSYjxRKYqN2PEZ2CmNVAyhTVK9o1rC8y4GUwSSQnN8pb087cZLuY30wIa6Ad9V++HLsgpFzR2KM
5zbo6cCGa+XpQfpnpH5MhNkgOfCuAF1odPtWM8s6O2s5CxOyeQPKtk64HK+0JidkZ6sqXh0zOfyd
EZTosCkWcFKRknlggq6dackRWq2BEKsJ72n2z7Vo8lPks2r2Q7GrqUoFX5VNKVBZLv/hmRw6igyN
XcM0uQdo2zIly94ptKaW40UhfP46x4LmLe7TI8US/TNXCI9kN4u2tVPK8tCBSQmLjeunOMynotLv
WzH5sFW8ADLjNUQdxlG7ba8LjDqByZntOMRJZylHp39Nc1fwvzzA8q8nG+sxBoi/GpdX4/nxMXjm
AIMqrjtNOhyqjwNpsBiBtVI0q6/A0vG0ESmeulQTZ+bf+CtXIngpvqXt/QBRYdlZFdaeloypvgoM
6ntFuVuNcz6C9qHnv3TmB3VXmjELdBKRx4OzFU9LQAX8LOUEEVfduRbAOOcoBw69zaVmYXEU6zsG
esoN5ZvGvZs1dT+ovgEm+ZLsZIf6SZ2DXwlUUJuEL8XkzPjGaZValxjUpgGZCB0de2UtJYTrDmze
ngSsGXwrAIr3SFU5reVsXgg90MmJaLKgb0ozzNBliXEQz8J/T4DIqo7YUtU1q3tPJ+D7CFbehrvf
DSRvZN5HnW/xNd7r/5J8ZZjsbV52BDVv14tk9uF0OiS36QFTi2a4ZW8+bgV/gB7W5F7a+VTEsAt8
oUq2XSQORn/Ts82BDnubhrPkiy3mpXWY56AajyNxexWJxPWUDx2jDNJ1guRLDreJLKsmHITHxZRy
aZHjOgBmN/PzassWyhFhQLTccfAtyT9r7aiocvQmUzbS2f3UZgi8m34Mw42CYwCDOC1gl1vMpZHs
o6y5Jhm8qqA86Ps9pH1qTK7UGVqX8uwrETXHarBdNxeWCXE36nH1lYaaVGvaV8biQV+8k7xYNsiI
uTD1VaAd0WvqC8msqKXpt3V7OKWXyJfjG2Kp9cPIG/GvdaL0uv5ntx2GXsrck225Sw+help5taem
1PTFJlm2zM1WYDp8bplB25pzHp0fWkWn/Ik9wi2Ttjp+gm7ryHTobSYLSUPBWsn+0/r3t3tIF0e5
lfjSMZuf8VBQA/Ep1EYnVQKV9tWQgbSeOfHLv8XwYVesn3khkdlWol4bf2awAbl07qnnK6hNulMb
vYJxlX+uOHvJh6w6F6K1mC8rgnxV3QWYaZmLOIWasLWdiUL5X4b2vU5FLzYZqG3ll/ByCGIUFIpe
8ZVZDbLNn7LSQ0/1F1YKKXwPB7zOHR3eKubzxxgX9R0B6+9vbrNmwFOxgSNHyOtYjL/8vhESlyul
cjN6kZerbrD/SLtpqRQ0jVcIN5J/5yE2VZlwZBVKcalmIoRvdZJzeR+aYIEEZgWoHAvLyaYApmnC
+p4E8BZPjuaIOV4sF3iYPgE8sfruCMA7+gGT69xNa6AJV44pITTJYxZK6I+MXZpCY+4LDUqJ2wYT
vrceN6KAI3mvH/y755kOPKRqiFLGFWJccQSnI2hJmdRpEsgt5G4KEEFJxu6UfR5vlu64Az4QWIVI
uiEpMrWDDFhNC7/ezsRzPjk2Hy2L9OcdnKkbFrS3U29PsQxTYPyJ6J+AyQ6x6NHhNEQVMmwkJIPK
8tzp7qpdrktlLmUASidyWIFmzYGv+iyQnjZvo7qdngdbF+jU+k3P5vgkKBZW2CqN06SQXwMcFdJT
FG2Nu8swEmUzG+u2inejNB+poASwBcEOPofx/1S/L4962soEuJLW+VW2kUUy+8tW+PC6/DyQPjL5
yLHytHfaNeHIr+CsqAtpBgP+pD1bLeFqbYZZi0HNFsxGXg5T6noE7E4VDLkvNe9YBXq6Di6KqdTo
dXgKkIECpjrSFqwkmSMLqea7879gjttGxijkPJfbFuTisnKh8ahJ+OLLHdu/xuYEHJbjDphX+Yij
OdchqvglhIHQuwUSj1M39Ctm+3YZcsXlWVf1i/EZzSemaVDiykJPMRrXbU6/uGRl0ih0F3gQVuYL
mhduaNdRhxtYjJ+ZeDPpl0Gr2/dgi5TEh7M1aO0t96dyQviuMly+fOzkmxc4Vp82pwGUm8c5itEN
pemsTm11MAtdpr0J9Kr+P3jTaUcKSaTe0JYXOJTyFjWHES3GSvaZJOnjBzYZ3xTHyyHINTYmHVBH
dGyHFx82QFUghs6ug+sO3dBYKORjkD3Y+NcN53u/3cbQYXDGxE6Vi5f86XDDJD6NkYOpWCjtTVRv
AifUsx+J9q4Y127l7OwG+kmuXcLX9cJFn+d9xUcsCW6ufGDEi1WIpc4yLL21owRt2Z20Ri4dQ3sA
+9Du3oyhXtNTb3MfNxauQylegG4IwgE6rtDWFMRp0NlXCV2EpiIu1tJbktnHC1nNc0PUc0GQ4ANy
qjW0AL/ktt5/K5g2LMSGKnPmkYzP4Usv7nNd2pPLYKEX8vU/z7UO/ujjdn75bLIepqKNmDCY1c72
m7wuIdnb6J7fKndHe/EJacGJVlgyjqNG9OWIvnWzdQQNU6oQ6/U3ov3eaeqHsYURnH/FIenAgQ7i
sZeZWIxhyA1Ec4EGXUzJYBqqf2/2YMBv2j4mRpeU5R4DPTBQkbB9fCPWt+/EhIAJ57CSIBN2ZYAN
s/olrd4O4FMUqXqqEC5W2yrPFzzlLzzahrOhCHr8NfBYdbYb2CUysmwf0E1lzvWgDFowXGfuu01P
rMMmEvdRp6c+7kDazEhAqNnNSKOJQNF8+Vb3KbwhXSy+Wwb3x5fOKUrc4yu0GF4FLF7JxHtOoTtr
Dj+QdRG/GS59Yr+w3OubXEJiiVPs8+8XQqvHA0+bKfrQ2+i8xFMD6NZu58Hidr6NHRKsbf6zqBc/
OjiPRbifW32u48dUYSYwpKnfjOXq+652JUXd4yesa4krsj+krq52Ir56cNL2hmK8Lit6NAPFD7bv
rMi2yCtKAK4EHfo9F8atbccJJuCRaqRX/PbwHaFHjpbTlogl428DVkySuoHI/+dhd4bxkVwuAKDg
twOkvmqnMqcqLXoxAfBOB9XgXxHYeHhsRleQ1O2i+qi5yh+Mo1avHX4ShruDCE8zailWn/jRbhfE
sz1bfiViRf7NyW123WTsUaEaWqs2roJpq/Ib7VDcNPb/My+BjAHBZ+TM2prxPydyKNVADkbxecf3
ztNTYTl7E/8cTp9cnwrLp7BZDpmLk3f2/uX3JqvutEnwwlw/RhCfSpRUWbIetbUJmRGEuHArF9mX
SBi8l6k/wmgDNKg6AM1sdIw0hOc8xoXajouc9V22xG34wzsD65gKWhu7R2AfrwAlOYCWNuw6HUdn
Pv/vaREICPF5LNog+0bt9cAxtBBf5rRZ3KpxIey9FJLpGMY+4aamFZmdCV4qlFGkCkYsSuRVTJ/R
3o4BRK36V8Fqao+rnybOzeE969u1bSNCIfvEWd+29yS/Mrtn/90rYYh5eL6xlz2waLpUxFZs7zjh
yPeuRo6q9HwvRiEPdHloqU+QjjSZOi3tanhOjRracYlp4SGKA7WzQB9+iD1EdnuLTLK86vVK5ylY
/wXlLctxvW0E1Let+t1NyxJDTi7aEtwW8GGLGB3INHrNglwJXNNUtkKLTOxmz2Y6j3HhwnMI4C59
weUx63ExFPoHVDgreoQTeNHvarYcmuv+0KIj+gNua//lp4wEB7lCyzUIlubIWv7FXYx5+xh5R5c5
5jlKmdwAv5jvR7396hVO/7NcNfTHCvI3tFORNdGLcC2xhy6lGBVj7+90EWb8ccIlVSziAtL+e/GN
0PvzLenOBi5+7mK2HtR/akKKAf9kX7XbOrysJDSDgHe5GLR00hAJD12Ufh5IwWdP/fnIv8z6hnji
l2CXdaAt1KFjOhUvulLRup7v3M2xAUitmpca54jCAak+IqTnlnWPYHL2OcVxXkl7ftz/MJ/OKaxo
FwmBN3gpvSJJRjz8jk9cxoulkZ8cmfn4fnQNX61DfxlzvMV3Q9lCOb+gFfR4IRBLDEHPgBeNiKfG
/GzBlYz707yYVbL0ICTCzWVtUIWyqMh72s3fLA02YaYmtchiHX8w2l8Ibp7y4CMybBC5y3tGgDO5
NK20V9AiUu85SQwnG1Kim5G8iBccLmPy94FM009GGWop8yNa0jiJ1yYqcdhbcvvSkgpVdZTsJZd8
WvgX1jyzQvp55CtyTeQBKesD3b0RXgh8sqPV5zB5+srdTYyZowXwtLhws74vdvjiOTXp9dQJiVIm
dQgXEu2P4QtLdk5m04kYWtao7Gv+uOCHKHVCsHrtBnBHXqFAXVNcp1Ea8a+sDhmCDOHVexxxFXDt
oAUDQEPqdoM/JsLs0KVE+jQ78IzrE3UzbVMzMPKjbzNZcD/RcPt1VJHAPjn+j1AOItaj49YAlA61
Cq9/oC+g3xiZOf3xxojwJiyLyBOOnq+a/BWMuQ08wlULY5snGEOLQAoflsdJfp07Baw7xA2Pofnq
pt0XNjlvx9QIQBka5T6cwDmOs+GjUIlUIwE6/vIghzZ/TsrJSXz0sXaLSOCU4EI+k4vUdr1+BWFu
0HSqKklvb3t6u7VPqE6fs8BxVyVgsR0XTiZlgsZ02g3c+y6PKbe2rMAoBxERkMkK7CXczi/agYst
0lEf7z7rwcQ5wDBP7Cqu78E38bjPl1ajJVSDWu/nKDvLX5UA7UwHkamFUWrrF+5vR1PhrvCGKZXG
uxFocRGwCRqZw+DAhSFrgk5Pn8KPHA6wTPOfQrwOC9g3alnXNswqvcOwWj6mpF/M5n5FzLhplkeB
fawcI2lDui/6eOT2VOGiJ0wwPIUlDdDujZ6n4uSpWKkd5owYRR+SWJ/TQA87014sFWzHaapVue6t
MEyOyykcdsicbo6C+kxdAeX1PK+gn6TAKahdswWm5NX0vnnJth334fdAo58H7lIU7vWWYiHwAhys
ijGtfwK0aAg09gMqfbRyLdGGfKgGdYQdB25xgCbRlsZ+nSj6uDoZHT1AjfkNjroB7ABeabncsLCk
t1stq5CSsUKnGDEVVNYRDLwVQlADtahQvd+N/07dLG7Axr+4icEIej/amCBDHE3/l5rwpICDZrgA
peIzb+Cvx5U1uyaZW/sTtMR+uZuUspKebfqSP9P5EpxoZLuNK9KpZb0YcXV/hZXL7G4otIsBsQcB
cr172uBQD67JOozH/ud6MBrN/mFG9mIpYg+S62RvzMgMzLKzZwMb4BzBeyMs12hMz9Lal83T2Mm4
W0iSNLxH+7c8fWwRi3PrBdB+eq3EcleLr6qFsON580ruTj/3CCcAYRlvU3Ci6EC2CHkfMrNYcITp
hu3YmLA2EnmHV9voOxCXw/9RQZ1hOOQ8ocjJ27ju2I1tRiY4nZdM11S0KgQddYBtPw51DQCmiaYb
0Xx6TCJzOcqVnBBtdIzcsz6iJNzmKy430k/tkMbIPCh2PWkxwjwdIPbP5XnGVbSBGthmJKwgBxp+
fXaNP3AjhYwc41phV58gJh6B+sjZ+uI5Rwe+2kcJIyBNAtHeYvtIXeLLdRoAoEfpVeRZnB3FKTTY
Jqkoypln17yXSQ1gZYSOisheIGXK26CgoWDaz0Nx67+MKAfJgG+4J84zuE6l2/im4UJYSCGFje11
REwC7Zkr9jnFanXlM19KolREseOUd2OgcCTRKdmcOKZ6C7zpMsW+pf1R1HOYH8AVCn/y6vfIDr4a
Df8aTjazyOsE3IzxEVsxWiU4YfmQJOePOdC11AlrO/JnEKFw0xzjv4uBVexdq5LUEpK76WJwpW+e
xrSSG3Ell5ln3sHgUHjP1BjtpD4MXp2rc9bepv2k5bDnYvZBFo9q+pmTOTwT2kDwRaNPk3MT9WF0
piTsv5MXDcnskrDvORGmKzR277x6b/d+Cxln4qR3phyY/GZ3vhP/KYtRM8nd9OYR4Of8quuxUXum
DRo0xTXyVbVC27WkEZ8pWyvttE/bq76alkEla85ktk+XvsX46YN5BmR8AMw3RfGHoAreMbZHLaJ/
7dGP4HccJH4w9nUhmOoixvqHA1UtbfG3VikXmE1nQvfkxAm463yR3mAfhFUirmJHumQcvqd2HzEM
zTTyZOFBsQzZm4xvdK1Zfkoq06TzTCGosCf6Ayl4Y1iedRS0wUjb0RA3JYDHgH7GLNX3XX4Qs0QQ
Tzy7fT0A5esDaOMqjd7NaySwsEy8fjSQ40tHmvD9PS9ZG2r50vg+kM3YCoqX4bgXQs3hTBob5skT
7c+EP4GYDjNw2ua2ZLNJgEIgjyMEV8rkgCqriY4Y6bKHD/p6Jc7DOQ0umXLBNF+hD50YHQLo7ZyW
hwr3tuPnK9CIcZ5ggvshtGwBx9qPj9WkEHDa13Nbu92DQQP0DPf8aVmgIw2Ek9p8zriQkCVWk0rL
HC20CJiqLoqXPsUsQdcAW0ivKLWzyHb+264/cc5NosQka7zgskjtxnfnbjbuRXemp33YJv9JIxhh
aLXekKK9Up6FExRCcZhiYlXCs8wH7fXBgVokvwFSmdoNLiqiu4lqvdQN/qSJc+hNudC8sFHfJZY2
qtk06mO+Sc6BREssIJQOdlLy2AefhroS9ToPGaGzGKncfxx70QQM6JzDBdPoRCFYVHj42HmjuU7+
IeLp+q1+VHBPi3N0otKmyao9NOEWFqLHVBSop4JRCr+lH0PCPdXeEODGsCeDq87OAorriDdk9nRp
z6nGlaIdq81ZuWpqK7IGJDUpgOwtup2g6LtiHc1Xd7vlAHtQnb6x/O1EuAWESrpqRivsyGmrlnPI
eTNId8M1+bH9txqi63ZWmoAco/BhWV8JqfsTvmCIhKTWFOhh6d+NfQ3xrZRVeBLln4/wDujh9War
zm1toxxXOabf2ciRDvMdM424pWpHazv01fn0zzmP32T0GBWSB/20NVaKgFhYSkIIgxctPqnn8RAX
U3NqL8Hp+I1y5bmGJZj2eefnClk+Sx7BLKGSK40NP4JQH2elzUAFNN/J9fl0i26rq8Ckkh6tnyOc
MhOMDhXc4pJYsDR4JHDXWaZOfWo+z10LI/jwh4cl+ZyUUFObEXL7lu3BBR5OcB1G7jZ+n2Jzuy/E
FkEHvw36+XiglSFssI+JPkFB8sbXXWxyPBXNflP18r3mXAsENjHvqExxj8gsJXH/+QEHh2BJs0UJ
KI6R6EtYsUoPJ6gdmKWGQQ/1ytB2bAzquvIcEmR/1tI8zct/rrv1JSsKP9xyXuXIeRlJ3rykITYu
49PhG/DLiKsBbyu5VjjMkQueWhFpc3vroPZF9l9E0iMfWdkuvYIMNAYzNhs1cX43YtU2cl01Tkq5
N3ZXGRMcbmaQgkuT29ga5rY9jTN0+VAMrpINmmoko5drJ0iF9R/Mt2GgFc8/G7qPeQg5p1sgM81N
10iEGCYVOOOtc9XFRb9t57p9fHsmWXzxFdCcN4HBSs9w2YIaUQrGval5Oc2xpPT2WTFirWST8yNP
CoUPXzMUEFEW7xvc8JXoVvkS1yJ3nb4/7jaxOlpN8nIDXHNh3J/kMWWYNQtz3gVEAVETkvK2VL9T
Guz5NTzJ39tYVy3xHPXEFAPX273PwNj+cfC9zcwPg1+WUn0wEq3wAPCd8Mph5XtrdZwf6tDNcWtY
pT31xZyBzKSaMB4+gCaiPvaM8tA7DgeMnfM5zUS9K16GWezWRxZOK+bRjCsidVXZUKWynq8SC5bh
rJDpl7uDefVr/bHj8EEM7vQqiSGmu8QxE0xVasGhpRIX7ZSWmegswu3z4zLYYF7zABsQG3SI2vMG
Za/Wug0nCxlVfcScAwJRXccutKpJc/SmCI/TlrdAq6sFWA2zilPJinIT1fytbSJY7ll7jdYStUSs
7PO1ICyPidLsq9tf7fCMrgGX+lNIX5ivimL6TE1rbt+mGrNyJ9tczd8+LH80Km0gRrbXiI2JC2We
hKP8Ea0m1cvMxxV5CRrEqJCICICDGo6NGoDzBgzNnb8ZHW1tsOH9iZAZNq6sXELnZ425UOQ3BIaU
gIV643VeJcyncOENnOMizfC92W7yfEEMmU1+p13G0Zv0plVifIHkBjIKg7w5GlpCgLqVbzvysHMe
Znn2BZMj9+ZJJujtnCkgVMelNJTjtiPR0zJypKc5OJpkakcbqYvSiNAyB2I+sQctbxDqlbzXEMa5
TjZEgLo6Jb6426dMCcAuhFFcvnv/uRPD9hOD9G42AITkokioQWdP3fDcMxNqgyEazOh1fWQ0vv0t
32LVk11DOIYYBk/qdE+dO+G39LGifT3EGsg6SPJ73E0fT/Ickf8OQDRTfvllELvpvHKpVgoHXxzu
ZfmVFYud7gJoueNnNCunwqwrZnIYJ1wf43nA4mIjKUtuA09PcXu6fNgylkMo44vU5U+g7e0XLcsf
X9WaU5paF6iGeKObLDPtrf2nqqTkb+ai6mMDshWdEaOC6Xy1rSEPV9O8K6KgKWzC1izJVfPdjfwz
q/WRzhiTUiKivMPD/uGT3jxMuo025zacWAsMr273jTYXlyuj+bXb+i2ZkWATeDey7Rd+IEvoZ/kd
JvlbsRgQDk5FEm/O43fTox5kGTYlftigRvZKgs9wmf8H5MqRlxwRtfY6AyrvcqT2YdEKKIlpcL5X
bGvPbNwBOgqCAgO5jocxN0dt3zXZff9QY34PosmgIDZq6G5/y/xFQSBiJSE7/7AJbgyg7TUyNzxo
m8VWBxlkvx9ostb7PzJSzO0EBK029jx2xybQc6ev+m2R48qdtM0+mEdOsP1S+7weEQtiKKmcWHVC
b9sgUFYtGnbO99qmRWwLGc5fpyCgzrOI1BAIGAJJ6F5Ea52I+KnIrP2cdC2XNSQBLyWgedrFAUUK
USWhVwiocIiGGyBUnDSd2Q9IpZV0sIhmA/6l4TxgGc1JAAsWI/8pM+CXLX7TlfCQHr2y1qgVEWsA
o0zG+jPKnZgv0HX+MwOKVChlLnC+KGQ4RMnoW9SyblCFsIgBJjQ4LepeKMwqTG1PKwgcG/ZWfuj1
9746yt8viEUr9rdXveDzSGbsDLpjK4kcu+xZU/3U7RcG6xGiraom7IsAbz98zbyQEgJSdjcp5LrN
zUI83wVA+Lu+35pDn+BJbfvqzCtNTv/IPlLBfbtI11p0wlY1JNAqgTEWlPfQ8kAmz1uUiPfOqIHk
9UjCKPvT7sziUUWxhjlFG79NmM8za/Z6wADo1+uxu68AmUqoDey31atR4c4RQOFGrjdI9tjnpgtu
LGhYgXY7DAcFk3UxtKF4EKWkMvKhtMQnKQm/tvTOH2RYoTx2QtqaU+x1UxHT56rtKpvKzyinYDjI
Zv4OY4omH6LIAiDXOoxXnBGtdvM7DG1VHkaBW2R6UFe3yAO3ZG+OicPjwRB7UGWgQGznSG4KvULz
4XuoPsR+Bc35wQRTmBowvFx8kW/LpOB0rZlKNNhHIHc6V/hT0H+BDsQTsAHRh5BEkzpwPhf7tz1+
ClMwoLdCUjnoUljhTtGlrHaLNrgPL1kFPOnWjT3pyY7Ezq4XROhrsx5DZ8donUjiPMopWOMXR4D4
lKB1qg1DTBqfS26PyDraBhfLkRkUmafHs5NRg0YJGIszN6PNq0iv2+PIln9I493toycA69CPjCvQ
dlfx/rpqKYbBoMgMNU07g6JTxGCBtfyzRvEGRI3FPTqISiqvhRtwmK8+gwLurKYyuoQ+ELXDbbHT
CHuFXxRfPPaCxv8ZJ7PSEwpo7j6DWLNNAHkOAJkx8XF8MzXbta1COu/YoYXSTNQYidRxz0OeMxFp
m5krL39L6h3pUQQUUoH4EYWmQXiSHKNumdnHaNqVOk3H5u5w5Nkaw/6os+9ckKMgMacqQcuhN67T
qXmFUs+P3C2rXLZOwS/C+Qp8AvCefhyVo7LvcRtyBS9jorBI4jRxEgE9OBZQ49whoQn81l6xwjBF
zF0t7SyuNm3Z1/p3j25o2+IorQQqUH3CxtFh5sBA0NLOFloE/qW1doHFYhR6sZD7x+GxODMeM7iR
OW0CH/T8S418E+riBzVGg1dHciuclo2dFX5bzBHRnFkGAWucIpaK9ue6zLRmMjW9iR2fLko2xBxM
fTqbsdKcMKRteE/SqXPHGIHotLF3HgfsGkAU/vqGSUtrI6eWj9gACR3ljwPZDr1th696nU5e3UUx
W5OFwj3xQYKWulGSEu0NLnJ4A5uLY07F+tTyIxaRRCn2yNGYvGD44kOxa5E9Q+Un4vPMYSalrqvZ
XqIp9uPUlpmc57j2VUpdQ+a/GJdCCc3fFxWyNEqzvPh4YNuK+tqBHZsgbVK/5FhNWFk47BbvF4yn
+VIk0MLxkoi8wDywtdJkjY+nRmKdlKw/iuwU1q7cMPdDeFEZEtua6J3Zh19mw24Pk6DLQR0l0WRx
H9mJB8p5gH7h1B/s5K8aB8ET5TNJH9VzJ466Tc98cQ4+b83qZAMuIyWGeFtKckytP907cum0MfQB
CIAkGCg5qh+wij74F+9GdbNyP7zMzeQ9AqDQYkAdMPHdlUNbBqw88jCSsigpmGQKugVT2c5xJVUz
GmQzhsockSWpMlQABd34t2rripAYPGSBZmSNlopatUQ3e36aTO787epVRneVFkSkVbHu3SLGxNXx
LeLJ1gvC82os1T6zed2ghVRTiP0ZIE5X/FCeK74opKWYEmNvt2KW4R70E69pp69mrc1PnNwcpP7i
raKhYCI+zieGxfme/zWa0cF89+R181RmDP9awWRH6DdFOjJtf+0np7lH4sxprItyvsAR0UWPno0s
t5z/jOou1G+ygXrnq/Q+Nl0BLwcWi6/2uWF13qGqpMqZ1w1rP+KugS1bOJNL+vkDS4LzwE0L2Ukp
dGn0681KhsAlXwJgcsD7qWh/BLBkE9C4KBG4qOlsdRS5VDR7QAxyg/j9VFY2M83kwo/b7S4OWEI6
MK/4Kq4FxT75vtcZcaHIR+cVrkkeIWyG4d77nSt2f3b8xVJdUIDqemTZBSlH0YaKSzIYdkGbQ9XK
Ff/Kmx1QEmbBI3xipL5n/MRWXWw95rKNNXVjNTcMUL8Zj9ftM5GSLqBeY7ITAbU6muwyhIiX9G2M
3p7uw4Rh5Xi76muxX1wfjiVJp1oRLpmotM/yVAdL4nOwoH1SA5GtHSiyx0Madxt0t2VV+SRlxnFb
g8sBQEnpNYQt1CMD3LBAfYNR+fttRBZWs19YA6rBG+cUA6wYu+TmgqlMjvhwdSRUZ140ZHZL3y4l
bYaBEcDVe25W4QKj5WMHfbSyk4Ia5HIb5gSBMsL/pelBoHPkF2nppEw4gaFCIA28rQh4rp8TJxgm
0i22RlVEWB+HNYyk2RE6iiQ5IPpVPytoZis55ShZiSr3Jh1pZOJ8eANGCAvyxmhkXkM4Qhvgk1O6
qsKBn4BMCPvwT6E6Lv3Ufz+fmkyP7ticSNykFoBtO9gVAQu+DIYWN+kXALnZ1Ns708ZWF6XaFjA5
yU5uppaObN9gRqg/gRn9hZ0ecxzKkvS/lrkc8pZiNFvFV3JaR0LmJHMy1RgHdUQqRt+l3oH9L01m
rIneP/myVrJ/xhcCxAfIvaOknJeEBi+dQ2JP+AIYxj4Az+DlpqdB1TLeYIm1GKi/59sjNJX2rvOg
+rQYOZLTje80cdhUC6peAhfCKp7ej61X8ReJ+iKwyftf+dYyFsEN6rBlO3FnfknRoq2v8mzO7q0i
NsguQFShtHKfPT653eCwoOcJCxfQqNTjx2iNpJSffW9wYMOc0yesESBNf7idiqmf0Tf/2llCwkOa
GZzEgd01Z9tXyeHd3Cp5QMYPCnYWT1dF6aP8sKzf3T464+2YKGur9jsvF6YokVwlKDsc7bGZM0La
axTpdpr1OrM9PWHLBjC1G7wFaUpaylJssSqeOyO38+nShnCebYLjajaAp/h2b/YR7XiOiDLw1kKY
RCW5yghyfJ2LUAFlpNfchMJvhYdNCX9OYZ428lclhKMp1uMojxSXuxDtAopkINhz40w743zQIu8q
xh5gvzhyskb7NQPzdZ5S1wCPwTS5BjfN+lT82xIK98Xg8Z8CI2DQBqXrU8WLpG6QoaPpWqboWzU2
cHfqHEzvYiuOrbz4O25/t9kb7dg+N+PiLHq1IIhq1m8WyYgVg5PIeyjvgzxXPbTHOD0I1Ncur8AM
jI9YEMYqfsDwoL/wHI0B7Bmqs/KtzZL3PUIvCJdD9zjHtAdSBoH/oBjD9Gx6gxORNh3nMDtWxdsO
3REL5wGEjUHzbxfAY/MSgNeOBB97F/eKAS5svAyLBiVsjpHdJRhGSwaJ01PS7lWtKdVO9ZLw2c1/
h29pN/vaqwFjq9iDs5gyUX6AGa2U3EzXIPPj1p34KWtBcxvu9BYDYiueL23/a3pdM8mdITWJjcSd
yAPwo5qXw00EvpgCbS9DMfbPG/+Z93TF2WJnsZzVV3Ug8ArIvptzJPD8U2ydgMkC6krM1L/fytS+
Ia5+6uNwwenekv7ysnYVl/+WCeqio4RPzzeI86izIUKFUtoTNvDOlW6gA2zM/IUqrWzK/9XJs4Mc
AV5qaLTAi3U5oUqh9JfDXCTxyDMwdljWoawNqNGQBfPG/ImntTwB5ZdXAbP6n+lFPj4qOfhpUufv
OaeVe7PAEmi61SWT1huiZQh1KlgVAkBgqBmGB4ybLC+ixbXKUeQNjdbvhq+A+i2OeSgkikLjbOnu
JxqwzqXasY7Hmeav74RnIiRdUtbohyTwPQW0Hx2iIAcH46kzkKBAIi1rQftsrICnX/BLIYtH56QB
0bner9bc5j+iYY+XxD6VElikRTzm8JbNqG8+8+Z9OAA4C/aASTrRtSK34cMtVOB9W3WY1MEy7l2C
tSlKkcG9DFuz0DY+LFixR4SGN+iBbFqV0dND7cF4hXGJQr03ifzFWG5kry3KX7CEZZjer1CBbfbO
EmYgG3zPQO2Tr0Q8czGSoHD9z+jO+LU5iYHgjaH0p6mVVJDLygRqpqgXNMi6XVuK1kHPRG68b7/N
5rgRISi1MKbihdKkDHEMGeD3I3fQh83IZsEgSy3ZH/AWekLWFZiz8e7HT6heiBI/RrMXcinB2F/w
SEj6W3R4Hm4v14t3dgxC/bYllvro5CJBZUTK9QQySY1ay7IPC81b9BDkqFIRIR7cfpW28gi3fkPA
vb7RUz2mliRzCHMU7HxXZ06EQtuimLBuwMrlXFJtAQgX76Msq4BiQpGGVbsJ3Ooq6SiYzeEfYWzO
X+ntkqgW7gNCp4xOtW4+DRVNueLFG9w9pHgDz9DKSkXR8KQcYlPbHS1kgcl5sYPVDGEHznDRxhQ1
5F2gOWM/xpK9YQyHp4QsusQBiRO0oUfJzIxRZzsjWFn+wCvvqdL24VAomNj5nZpVcrUz/loMZ4eO
Wo1Slj1GOCQQCv0nvqoCBHAU0s3rFMjFJ/LJMeUhrMXHDZDIlhKugdglFgTutoIQtCw3PXxpQwTl
dnzF/LUrwX85SNS3Ym3xnwl9V6Oion2YK52qOsPPsOxdJhxiKrTJi6SoBK2JnhnSrHeCK3OG6BXT
68HdtkMpBxX8mZdrgr7Yrv5bRQCGmq7Nixa/wtXlvSWY36je4VKp9JHHuYeHBid9kvCMGxsyvBOz
+Mkxhe6KDXnnMbSQVIN+E1Rft+UNc1zV9UXWWvkcrM13T8riWrEc5rTYbiOUMwt+z21OQlf+jTO6
cjPzJMUUsP/OsayMQZmnRBjJI16iRNxFRG4hs0lbzmdFr35j7+58Em8pdvtX/a8TASu5/849jHdT
fG7VhCcXhgeta0YlqCaxwmA3wDQz01Dpz+2gtAbQ1Y5qrrAszwNsbdUlrvr8SexFAeywrV2Rip+4
tWekPihFtUF/PjUOF6HkXEtuee72h+K+vuG7H3nzj8H0TPlnXEzuIfHPbzLAzOsUYPN2L2mVWT5u
42ecGebqalXpVmc/U2hEtSTyKeq0JCxo7G3DNKE1ZfLarvPwnriTLi+Nh792qOBfgmrXkegZZTf1
XuFGTK+0N5yY3BHT0+vZTNrQS2pUL4Z9zL051lGRaXOKUda9D60Q9lwjPiFkQMfGSpwnJ93T/WlV
Ik50E5qZfLRA10RCqB1x8KzpDFJM88FuaFMhnmdZ9BnSxyJL2T3h+/+hrIWbMofcyhfN5tIMf5XI
LcU8XHzr18RaPcNC9Y0QS1yU6aO/uACjKHzOlNgjKBUws5HqK33XYLcrVrU+y21AMyygQjD0lxmJ
Wql1LBFIQ/wykDCGbpg14MmyMYq9kBALBVvX1RGnmlFq1mRnnPHHlVW+971INJWBNdBzphDoJjcw
4nEzRqxkaLCWlCVPBBG5pY2M+HTsJCb/nb72IQoISuyk2FrOM+XlwiqOqO58ZOFVM/RA57fWOgLb
Fz4XC+eegXCJ6j1IvG3ueKnzN4QloXQxxlvD3pyrm91+1OA1D5o6VER7GYp9GT/HdOPtJm05Ci1a
jA+Q1wm6HT47K+jz+98SevvgSx9zv9J25QFylwFD8d7M+rptzqHI/4awF/FOESl8yW3vwOfMVcAU
bLDwutSK0E7s482RSM3jY1RIRGdD5fWg20b/+XxA8tbklCiLAPGLN+5ivtvlxxpN+a+k5FiZXIsK
QB0VghonIxUuhcxBzLDmzeeesSexAPnummGnaMcKm1IW80wTSF287fxrTy+xu9Xqt+BZFYtBvdgm
ecgQ1e8KEG5Xf2+TGJJoYZVPRgKI1qedEuYzbs4iED8V76a6bzYTrdFYthDx70QSWQcHc2QpB48G
gsbX2RaFH+Rxyl4cHC/Xnm6uWf2+UlQOAk2xFbsxBmV3Y+Pj0z6FTbx9FSbUVrRMxI5hFvBu7LMD
yKXIFgnPfwbOQtCJv8mXEQJXGfZD0ONegO/X6VoHSAnlhIjInsRIW4p/vLwa+YZraDpg/OdvIcSO
Rmu//m+ajkgtaO9qr2xvClgK7+5vJf5SqQgPIWwyat2v/V95113b1c8HZ8uHu+0BDVgzzZ1FBu/4
JYLNMw7evUCCD8VmXKfLw9/vR//J+ysxNuiaWmaPVuwOqRcu4eOaE1rAezhRwM2yUrlm0qJns64+
C7Fi4QV3/UGdSAQgUIJpqirHcIAe6/jE4QBFJQyRch7+a7IMuMh80mN5s6wEIHHDpYfdIraq+5cu
PLqSjfo7wjd2KJdr/C7hK4pmmizugI3uvSmvkTn1+1QpdSKOIQ99OIsqdRIkbF3S/8oMcMPg0Y4P
RKVFGDwmBRHxe2woXDlhP8SNhrjcI/fAM3BMhF6bXLaERLRWN9sqAyA1z9FGvY5RHsYQ48x/yboH
6AvlNoxJ5dbfuYcw8lbOChtqELB6einc95Gw/otl5NpZOtNU8ynicXjwb8l0tHryfTOaWf7gQtP+
pz3klLeF+bibeIfFcRWXEhHzbY439pwKDzJHBS9HwRB6LBBk9gmb/nK3SRYMN4jxonF8bnnReRGo
1sGLZvZpYvkDl3o9xn/nILrGNMmP4Vs9gufjzM4GVgUFznLtQifEYkPFcNIpOTADeT8eChiqpSKB
eyg9Z1Gu9enjpmZu9Svu7MIHk15cGTo6cG8DASwBc9DmQhA2P/+r0NNBdJArFBHChpZaUTJ3mPXr
cyR80yzNiqnq/RYWsUfjmsS+yjznXZj9uwNpXEjrgHJFoEaldQ09ibUMuxkxbkcmXQ2QqbstPt1c
SzTWxSquzrLZKoqqjBTq2t7LETiqib/VcHIxAAprSSQMTZAZbiNbLzPnmAdDhB49kru8Qxa4I/+H
x85PdnksUT+USHA5IxKVmuiJBpQIZOYzkh2eWHm5V6YYpx/GZf8e9AjjRELciW2pnp/0BBUZVY2/
ugBeOx4VlrRbCZ/V1wXYBeh+64oc6hN1h6SrR+SKdWo8sdbEbf+kU4M5PzWaZc22M2sGmlepVjjY
y5XsacFP/qLKb95YKhaWb5fVyuKy+do/p3j7EyPmu/WMVs8KDi6E+aNrYQhqTibh9zPVWqyeHHLM
cxw8J1Y5+XtsUmTHSA1jVKD8EU2wIRSrLcaaOaet4sAl5rIlleSr/mj55/QuG3Fm/c6i60i4YWLq
AM9IXhJXUZCfJ441E18O8A2LAdklDSWsUe4MXH4004erM/OZ4ED/Q+pajCOXyS3wZioNQvs0z/FX
Y3codQ6f95r7FUUNUZsIbTlKHiccBXqjaEenZiqQBJWhGv8GcuK/U14+1G9JH9t3rVsDwizjFbc2
x+0Bp7M4Ia2vILvxp7jfJAk6MQ4Rcgf33/xCn/gL+qVTRFdLv0Cs+CnEQy9uJRXlbFnEHfAac7yw
zrZ7FCqQL8nJOGv37P2P6bfnQfMBVQ1wH2ZU/Elinv0OhQugLG1muQp77imle+uMslCSDmlt3Fx1
15hHiCizwqxC6TIHQ4U5vILduqWUWM/vYN+2loRD9foypcYX5uurKn7YcWMEigtH2sGpD+dzoXFQ
No2aqXqVaBjNVh68RMITO6kTeWYXUaKdpS69JO3Fhlui5ilwARUHmrBNRdPND+zrR8g+7cZs78mi
WvUT7zWhyE1HRTlGiAiQgPKWRJyq6Rm6o8ZnQd+HrMXfetqkC7zL6RYftxJDtWhiMZJiXYEnFh2G
C3z8jBzaTcB85kwKmz+becBhFzr5pR1Wlwi3zhHzhR4iCf4lm/Pjvg0+Z47jns0IT9STBOSidPhI
fLF+MYKe8rk9jz/0ORZgYFgEObnognbRNcupkiQDbcPj5FraYWTod8dR0rVEMQGlRMsMmVIVukCi
qXBJZ+O0TAkC8UUsiaWBqXpcJbvmFznUt0Em7hlRTjUHOmGqcIPFJdcRoQ+P7UHbUCWHj7RTTfg5
Lp/N6LSjXLF5zS2G/kRogUmohIjPpfldibajaQVaQxs5c+X484rmohNKOC7l25pP3BHFXjlNsHUV
bJRMZX3Ti7clYLsDdW3yhi+gKXTRbQY4LeQEuNu4yIW128j28D8+cgSUWPD7aYcWSxwtJQxWO7gV
k8NG65XEhJv0W8Ioi8939xcBqoKGpHREDYdUm6KzDPJVHUeMed70sChrvHD0RuncF0rgAZVs4qYm
gcQhg/Jo1ut3HDHhi1TS4qP7cuclU7Kp0DbW/WPMlRnN2/ou4cnYnGR3oHwQOQKqXLjTlhIjomJk
LdUI4NrWFpvPYHrjedS7D5D49OMfIUNyg5HPo7V6mzI1vcps5/da158/d+oFfIIgzh7IyKNxEFPu
pms/mEXW2YFytsqDlijuhVCkDlLgAhhgqFly5MwqhGTyvir0P13jOEgn+cmBkwHit1n6eBNxQbTY
5C/JvbjckYHEFY67hnaojcBnEbrINWqZFa135dWx3EVpbsc3w/5AILQhvB5+jny8DxWHwBw+StBJ
rwfbQm+AbgzbjVi20VvsxIh2ScTBiPcdPRm+01BimWKyrLAz03wPhqg5WdSdiH+oF3s7S84eOBq9
g3ucAefo6vTiqrl8oXQZL6ij/yFE6uj7Aus6VuVMwHPm1Uv8sIvtSS8nUrPTkFglSUQ+he/ijXFo
TT2GXS8m3av3JhzjPt0dQVH7eOUZvcvM3QYN7tA/cXAgAGG+R3GXlwD74LLeF/BKP/XjmEVZOlNF
dQxAgE7L899Zjhw4o6KxdS/Zd1+mwUKvCIY2JYOu1wjbq1Vp2KHUr4Uhaqi1shvaeUMMWnch1m4u
lYqvSMOUPWFLCJzUwDWwMNae0vxeojTu1w1RBLGl4RScOy/EGrdxMCPqxe9LaMIhAVKm6WmN8jhK
d7GE8W7FZqbOi1rzGOEMA+iAPS05Ap0apX8zXMBl70dk9TR1AGw/qSu/5PhA7HQ6qLZcBmHCPbaf
Tn8kv9qGzvElBWV1MZBLZhoYGoD+3tdgLlT4kyOzJSQYXCf9kREpEbwEQ15JgV5W2zNJtouDy4We
0WQQ0Ldkz2VA46UFpjC7150i6SFjsBelKUcCYM1cc02Ad5DMz1jW0aSXeLlJqa0q8NT03ei6NT0B
Ec1L8xasTZ0qPPM5Na//G2zMDJolENoIhP3gE1A57FU8P0utLdlXKs9ZzFj+YUqf1PRs8czxNtGn
G9xrSscO10OEBpg8CgPxhk67tVKts+0w4FtkcR2fDYRnq7qqs7p2hF/a1yXhjVPdpdI5ey0jxCbr
BzfLZY11iPMA4CBtBp4iF2GTDTLIQ1hagP1S6W36tXLZKrLKwsuO/HpCWSHM9szPWX1JR3897I8g
UywzMttU4RKainPtUH4Fff2n3+n+9S5U+SNEwm33LhriBSWvZ0MNrJwYfXGJckpOX40m73kY5Ni1
ZLLyqY/IXLm3UBWw6msQiV/QIPBP3SuImj6fpA4+uPxKfWtfca/f8RG1faFb2Ia9pt9aaaThIhOA
WvKXfTC0B6ZqJhsolzR6CXN8sVnvchUgTUHkZ+ovknfhFfLwiIOGDvOp4XUuBqsP8rhuPEn2IB8V
UDnokENaKmWDgPrvAGcxKBvXL9OKxEiUeRO+xNkRRig7RLYs655C0yLpla5DARBcA4iYBiriXcqS
HLeKE0oLq6iwFxQxB4JPs8Nnd1DPnfcCtcM88zaJBZLtvW2qAMyZ0P7+WO81bGcpmUqQ65Hi1gfN
Qsb9nX/kYQfxNqYy7IEzAHM3h6JTb4hU+VXC6E1CqUnzXKVHr1om3w0ZoDb/CFBOqbkXbow9EHV3
pKtp7DpjxLCZ4jjP8uSsGZbFnorjK35FChy7kyCS0Ozjd88Uwn3Ye6heItTQnGxSA/DKrT4nx6EW
HDmlqgGwDCekeiM7CYV/p22tLjUIQFKiJ8EIh2JHd+HKa9zIbCzlV4S2pWkc9o3HVCkElILmEpF4
7fCWESO5XOVsKXQviO9vBm02u4l2bO5uIDd1x0q6ina//pZlvqzYZUcShNhrvDemhjzWSdj0h6OL
envhYUjCN6B0XvYne1Sutw9T+VxjVhbPoQJfA0Q0TciYnhOyL9PvNtOaZo3FmgUm7Cx/AP29IKgF
0tUsldMXOSV/5l9bJ6B7IiiURwyZrnwAXWonC2iwKUcGo/6HQ1Ape77hEdXgfMduvNQLfjmBrRec
rs2pxmdFxOtN01S5WI0waS9D69i3Mlsu8jJeIZIJWKmpjtRhlasN1wcoJwX/iwBxMGr2TOuMH/Ih
ydJ4pfg7IsBv3UwcsgrU4UMs1/6ibQXFnSiD0K6YEAm41lo40oZledaX3yNJZwxzASWvkoHDque4
eiXBniXG6yKLRL3zsc8n6i64HlHrbulyQMIra4qJPtaJcG/PIgdEete0ZgxuVdCcB7gLR80SL8zk
LNci7sLnDsl+boQO1fdy/bPAdodUjhpd9naW95gx1tSjDI6MdaS2UN4zpAEXdfUzCQJAm4ukdZMv
QnePKh0NUClwNBlBCpdllQdne+K9OMD5/VKrFKFnWnraikTSu1QqfJNuCGv1J6EzmS2C/YuQBaPJ
axxjyatS4UgwaWJJMHicZZ1gY/t5rRq2sadm5aoPWkTs1pPPCRA+DLWt7JXg4GLQvjamDkNugWeP
MEWsHYGx8aWp0wkZeLSEO3NlF8SLpj17CrjmMmgexikQ40ZxGHmM6V78lhRRwv8o9S9UnoNeTVdB
ay4pQGXhxvkfllIvJfnGeFCq3QNeHXsooSn3lI88qfjU4iZGu6pgSAR6hhgT3XhepMYBLClGSQBR
1d9XGO8fiUm/93+jXH2TcI1rtTgb5KnPuYlAkD/TVIvUOum3bQyFZ/YI04RhO/Asnr83JgpAVsKa
yRVNqarbapF2RbPBqVBotoqQ53vbAF+PSVecIpi58r7Pw7Si0Vq6lSooxDmI6GGS61zRvFCteeco
ak3D2I+6TY8TUndRb/Klja+38NgbwHRHGMg8GSI03Ry9uGbw2st4XeDeOEMvCkDR4MWEwTzkb71y
M57jk9R07VMf235br6szbBGq4SKbz36PbtfAZ3Ak/kbhtIK57ZEou5YJPQA8TdwiiqTHNE24BcMm
AMPKE0XKHGTDQ4+/3GzCPDAL1gyowk8V+gaXKVGwenB3ZmK5XtbN8gJqe25h371pWyFqNWlP3Dzv
byV9yz7C4eypxtX6XtuxTRwO3qn1ddjzmEuoj4r1XnHI0OkvuCLv3qS0SbF5UieST8UmdR0GJjkz
kElFV0agNtYMovr0TqiNVV9WzNvn4Ecnwo6R8/rafu+SH2J2VCQpprYUmdosn8Ty6Ht2uLC/V4/L
C/4z9G+yXufKP+orLVj/jW4SKP7hGTcMWEMruxz5SbZms9T8bCYUO10B0lP0wS+aXI6BaIKIOv9B
H54jhPB77CBsl12QKmSaVOLFQXZRm3ly57aK5t/q7BYUvaGVh4q7MXeifIVFHik8k4W/ns29+OSU
9KhmLhnCV6hUOxzln0ZFwczLWtJgjD494qXco13CmYnyj0f8pW077+8I2pmeN54oH00e7PAhWc5H
OQkxOgKf2hytd4WvF0740aOyhuigHUJpcicWsA3lvOmMU4Pgi/hkklGQvKGtMftGE3/feThUOEHS
zuaYoq2+Zf/Vcb1JvaDzA4Fx2enelJ0pV//MChCAQbXzxG2bp9y40p5dunz84O/0Y11ll70hDNZu
BJI+EkDTu4ns6QShqocNVloEvTF6uKhGl9+I+NnNCN+R0BmA/MpMbP+7qsGo3NZkOKuMnd5AZw0L
ZLm8gENo+/jlazO1tpQvY5BjZJAAkhZdIfH0IRt4VC+Es7mJjOnUUtqs+JJRKlaJRUZmgBldg53S
RLmaoR5d7Ri2vtv+vvJJKtQV+X/itCRDQ7dN2Kvml9ftGi2phZ9qAa6/cPfzvVz6d+f2alNzRL6W
Z4JII3fLrwTafgnfCRYtZKobebcGRGdYZiVcvMHJiblC6MfS/s8RmzkpoyJTWV0i+LPAwCOQK4zE
0yU2bjJ5YIsHspP6DBJKQzJ/9lPanwRw+rufje2wC7FBlJOTcVOc0SiLynNSPtCT0fLUAJPtZdGG
ANxRRzGnGug6pGpN6QJgmUeM5kB2o9SAlvI5YOSalH6zsrp6+/4L0ARawsFY/ZhZZKCaPPJNaLM1
pGLtEkaNWxhhmM0rCGX9eTkj7LCdHTNKcD6TcJrJaVs1+qNMozWVzawhIIsqjnvT2Xv6ssd54s5H
z/yqyeMNJQGSgU/9t3jzxpCSaBVDMN79lC883xsIgra2A6JHfU97dZ7RqvgxKj6YCMv7dvsFTmBO
ESU9OF4UbGBC1g1z44HGh/bck9W8MM1vpbydbKQWVkG02wfZuuX99BQAmntOEYeg4Pg3XXRv+fj2
7Q1G/LNpCm5Lm15REjmPAM7QXhBJnwEehxC7qcK5yahBkd8/RaoureYriIu4HIdxkoemxmPf4xPZ
LgcUUFWyfI7MolSTuRmuWutgHk8etFnR6Gb8GbCsuKNz20iucbXAXLILiA7vgv8P++tBvtbuFfWA
0SXpp9bymP97gE2mI8j7RLNReQZQ+un5M8Y+UQ8/QOUkreKRyfSecDnPpgm0AxTN1VTvRFw71i5T
oyDVaKV+qbBB/8fe5vXPFu5LCYAJTQd8WEvcEyHHT3VVEXX6deEhvl63aOZwgn4rm1jNXQWUoKwD
2HXeEG2Spag4iWyItYHPjVBFvC2WNGVUSznF+2m5z/Si3NHbcUr+a+EOeZZIZ44G8CBT4zbbCPfs
IkoJw4EzMRsUUy4oqwcbHD7Sd+8lwgpsSULvAGmHSt86vfNqIfCaeoN+sPTmfwHpK0uv6fZf25LB
FurM6zE93iIGBagPWRfhFOEL8d7zQsWrAMTs8porphzeZuqsP/j/rWAn3tzi67BK6dh9DoIrc9WB
JeFLtwqL3Vn4/GBN8xDS8tQ92/T4yEyK8jmm+jIqgyFpGtEH+ioAx1cbU4djZ7OQAb3HOeCm1h7J
785p84seC1P7TD20Tj8SjpqHax4TZZTQ/6ue+X1a1wK+WNrab6o0ofh+AwHx6Csij+PUH0EpEyyr
WCxGOl6RGOPJWCshfQBj7ukFQLRKYC9WI+KT+UfDMCgsdxQfqElKnL8RteNpptoC+k1rABUm87R5
cKWNPxjpCk+XoLEhnd600YFj18qdUeQNLeMOF78rgr1VKTclN3upz4/YHQ3CEtsrT230lohOfC7q
hCmkROZgfYHAVqq/3GLqxqvj4hj/CYkx6RehaTVa3gqq+fbtzhvkL7nh+AKHLQAJQ3IGPlDEg1W/
YASYJ068Kakjr0I6DgwBcYecIOXh2IiF3B8D0CX0n8SFMTVcHt+4PHplm7hFml2pKnhORC2DUWuk
4f9eVio/IeTFmudEcQIGp5JXI1uapnSc77ty2VQOwaKS1rEvpqlqXWe7zLLuD5Q7MTc+ChLMi4z/
waJ2JkRHw4kPoB/O9Rx9udHEOHD5QF5UXOFBZ4MSeW/HVdHEWcRU8ym8Ouxunc3Rvt3HT+gLtSqO
oY0C2l0RLAXtesmul8lqNjkjAfs7xWpRUGd2iHwfZs4P6Jszha4rHvROuhGCSIdQLPJF052UlOSR
gvL7ERMH6fblwJZgSSQRJtFbIqlGkwxHT8qU/OcKw8SpWZ9Tpjj2oc6ao1qTSSBVnpNS522iw9a9
geCpKuEJUCom0XFblVYOCBuAtNx432vuKLHWHVhbte3ZXTv58jA72yjKeuETOqRBVmQVX/MiJu76
cFhH25lYuED51omHFZuLdjY/HzLxjye/tpx4wGDrlwd87uTs6fhPLu2FpUfsmvNF/uGZfejkDVO+
sSgAYeaVfHGObPtgcskyYbZFed3XyFyt/9Cr/AcxMbV2c7s6jXEjfOElSzjZ/3z+f0MnsIO8Avky
TN823T231LuYu3SgWxiMIB+arUWqjlu38MTIaUuPsXfrmhPadthtwhusPHapp39j0/uVsNhiHWAS
E3zH8OaX9txIfidW/4Bj1IO+rbvZIXtneuHDlgnUAJ54FgXO92cIXnMBwYUiNFJzgaX7ummKQEuv
ouIN190T1xpJZPL/aL9+aipThpqaEwmY8+PIy/4GoCCrMI5ytMlaY7nGXH1gzmMVQYKp33ddsZVz
vAC8uRsRBabncZjsDBjbO5RoxCvp5aq8j0HYbSI4/jmmvec603b5s0GgIXOQvpb9a+WQcwTup4BL
gulYeBSsAN/u6rHlD7qXs9EAQM6HE1iAyaijmOrnh9Wj0DDnMDnjRKW61KEDnb2at50fsfJ3j2/F
SlNprg4q06AnlfeseGK22cP7bHZLGG7YS937t/GoK6G/kkFMJY7EMe9/KkQVBOWAl1pxQsW74l6z
4+FvhMtApUusNaD3VeEaNhjdx3B4fB8g/ZauX5JphggPx6msNc4t9yHcb9Lvwt/lIZGRuJXpdxzS
SfjCdfkWo+wT1BaAgz00HDa0F9jNci3xtrepYnWS1D9dTZXiD+13v2FHZ9jNxG/ZIg/VJq9ZnPpl
bFdGgi1oVUcnDkxqxDDgsq63mp4GfU8YH1rPIEW7tiKjmJa8aFA00Xmd2I54sWBhSQIp7sM22nzN
cXqZGRz2j3VqB+gB8iqq47xXv+TnU/THPp9mhJNJ9SQAuCAvqt+FAsfJd6YYAAB+tmcoCaePpRTn
SmP2hGX6hh+TMf3hW2wMmzlMnaHQXrCeyub24mIgqAOWfS4NJSa81LG85cr8NVchLYW4VX/N5Nfy
RCFloAeAAT1G/OZYbEfQc7OFG9tD/5zKGM5YxtUIjtCpuIo7Ud+hY2KAdnSmagzKTrTwvimJ66v4
71t3FXo0knlhOmNqC3s/KToK3ZO21nuvoiS9o4KWKg+RZXm9DalnlKCFK+odqiwq6akl3rrLgv1H
Ywx5Qr6P/EhgS8oShMcSzZ+XrbyjFISQBpX27gddY0/h0Pe9IGpN4ko8pPj19Jo9oalwZ9ChrUiU
pqlXTLhsTLSPXp4gCVmGRp4ONuaprBaLItYZvkT578VRKWGWslvqya28N8HHmGp/LMlBGRyODSAZ
cejKM+gLO8PFqeK+gpCbEhn4URzFBusmXXiVR76mlOskfGHZoukU3lZgQosAAQGS2yAeztJi8iSD
8JC0P0CyjhVCNdQBh2FlNAe2vchet+4CIISWfD7gs7Nkc74o3nLJuflMGzhmy3+O2FKmzJ+TtiNG
gJS7+Ts1D3mlMuB25UrkBM4DTcjDJHQsXaE0I18rXxo3DNoJQn6MN4H1HdCyd/b7/ieR020xrQyY
9VBZ1nwLok86d1fb43fzGBYdrLam9rAbXDHk5dyQ39k3dVUfzOLUhhteehBnD3GyaDXARjy4xdb9
NJNnNttCl+AaHdMD8q+aTI0BPHDUoN/FgLQj8ZF010uk1kjvgmZbNm6h8DzM/dk9UvJ8O+SAkmLV
XSDr1e8eIGrOyw28dyO8s/L8bMnzdEVVJEn7yJU34daPE2SDkHKc0CuiUhYB5dkB8M4KGE6wouM/
UP0PXTY8OOF5VBt261VJVyQ2USD38ea9yJozQtM9sh2HEkx5U6i4UxAHKni406kr+JGKI3lAcarh
JjhIe+j6Y16iYINirIeIr5g4cxrg2vNwNAjbURGlrcISuyYYEtD/mis5F9rU0XPIJfF7W0GA15Nz
f4fi2Ggp4r7C7bsRVAFJCQSrx8EAGsPRh2P8Vly1HxxBgfoV9/IyoGnqsx4OyGY+nyiHMNAeGcoQ
vEwRZKDJ0mBO4Xn4owq7ne/GaWZUdnfJ/CqPL59hF1ue3tRQgV5Ft0u0RLnqjOFcgZycYtC6ZTH+
pvl2CHyyzZp4L1++s25p9X6UZKgR4bcZoRU5Q1jVzGnKcHZV1jPNdIitCH0TbtMr+hPcEeWHUEpC
uMP+Ig6CN/JKSxqgKDLkp/x6NRK3pyiWI/vh1bnpxmZW8aqnV5P48v1jkrwKm/iVplJ86+56I4rR
2sZ1ICOMbc15uCqOUda4mhMHhF9hc7BPZ9wp5lUAt4oP3c5ceXAOVoxXSDeOlyukcznbu0+Bt21P
Bc1olCWCkqegbI0MhHYKY6u42Git3TSAkDMqECXZf5XpLU4W7KpGDmMgTyf30ohCYWgKhTiZLwUE
TEigDwSk+nV/0jeiE3xsloqRFSWkLO2kb3O2YKnWtKFOZBisYKnrg1lw1g0MsAJ2ofXMHSrqWzJq
s8Ytv1MjI5a8W8a90nB6QRT0j8P6sdQPRsPxUK4k7m2O3suUFxIZXkR5Cs2o2/ObOpmCkPjGvSnG
j7lTJ4SsMBW//3PtPdBwPp+CIxBGVJkJEKTZUx7C0M4b1SxTuVfW9lgPUnOtl7NXnYT3VAaU8uBh
jlb+hdFFyIjy/UG6EXGtYXrXuC0pYzHYVRx+2Ll+C4C/YyFVi6z5iU4mc/IFdjQ2rkS1/Qi7fjdK
fgr19cYss6pEy1m2R8Je90HMKbrUtEUGK/cBa1zuBYZjQRqoW3MTZ/puQ4v2SwJ1F7S9zwhnRgAM
rnTsx1cqX4w33RoFyJwnB9sdUg/EF3ONIG/7UgFW40iPunmBw62e7ixGAsHmA5lGkq+f7cHC+j93
kfzxRBley4lb3rL0c+iP1qjTv3bH4R1uKeVTKgnpRdtl/KNe5UF1cV3/g8Esi/ErSEWVm2JfBRM7
pk168YsMLWImrlcHujqBJ9aT2osuJtkVbX3NL+RcOYg3r/6DIegG3KzBKWBx5ZlY9C4GKacspo3V
9pMG6mX2Kx5mSZOubaXTbkng00M5S3dj0ckwSnfC9DK+45KOUso5xMTOHOCxQBE2EE/OGQtvBu8O
AV5Zga/qeJIY8oAJm2zmBai0DC1CBNc45VrfwtKX5nNvNxsj8cWdRmxLuctJt7mnMPxrHjxwMgq2
aC6lCuiRNaAQwkSiSNVVrt0zIWi8pWbwWN2yZZ2+0BNiPS/Z1FJEbTcZFBPl4hpG0oeN0hY5CfQ0
E9pL1NyO/2ualyPpwqqOCDDPjkSwL2eDLsPaIv1Cxm5xbsCLLyHKce+PoscCgp/qAWAq9/WAx0Vh
bvx+xXZdMvc+P7SZNQ5278Rmm9ZoleWNp7l1dVPbiK14pJTb7bQ1r31P+/ggg6C5cvOC+pR6yKpb
sqw0ITUXBYozd1uQ0FNkLYy/9E4dYwh/sEf7i9rT6ry++1nCdX4EaWwVIBTTgE9V8utJh3uKWntz
OHPecNI4XVvO23+Lp2EnO80L0/ngCM0PVsSFlmWe8v12Qd2gSFOmZ1HAYl6wJp8fPetA+fUe0rHa
oyYCz7ckHYS6YU8kYJOsBDKywYT5A1WcPDUZANkA2ryoS8jP4x1jxgR7wGGANSiQpt7V79x6yGFi
SzgeFSolVaZ9ngz+LKMchq/1TPL9Ul8L2/cPba67qw9sDoZQFS22cxRhfPbNxNcpVZ6iRFpGmGZW
wzTkgMyfWZ80MkikemJaO3ti7R5WtX8Rr/szCgrD58lm3Dwc8jGh03GG8zx1YugulPisrLvv3v8K
iQaugBpsGmAOD4lvdpEvcr6C0TIopXSlrICDb/qI4MD6D5iQesug6rGuF4po/FuzEjhFhak5rKs7
4aXF4d6qrcivOYpC0XvrRT9EmaLs/PvscsxB1KF/TzhP9SIf+KudiOOgn02YsKE+9RW0Lg8k2tBY
Qk79YnwMd4iEU6HopG0lcfw629CVuHb9Y7E1PY51EZkQjMM0F/xlxGWK2Kno6VUUlNkPFUCMEXpU
THBf4T62KlUiIM/LKrzHBTCMbHOvgpnS45sxgp3TezrKic8ceuowKN96CAbSSdfz0jJbLfiyRQSM
lLeM3YA1/LU3i/v7z3Gqf0J7MLOLGlpBF3Usc0mSxDIgzBm5m+DxljbJr7YKhg5pZpHG3KBfzues
f2Q/dS50f6pWI2KLHMtL5JmPZRVnEcv3ZdderrGXjccm0feGZ0OcZj2p2nx8iFuLnhut6Uds3DlK
X8TVqEJ3sbJpKUVu9kWSUBSuZ0mtzralBtO/msQoV0LCc2bdXyi/1oZ1pjW1gB0o2AaE2SByQciG
SLRiyef5Lmkm8yK6MUfsZRNZHrVdeHVH6vdRpgUitGV1q1GS99wUKXZnIPOBMmhCPacNp5vQvKx/
cx5KGJAZkv0jJIX7ciWA+s9jiXosxS7yvvwI46WnXKXcfnJnUhQEcBT/e4q+YTUCxf1BrnZlHgDz
YFk5bFuG1LyggQmXVD8kuBiXOlpERWGsfc3R/TZcSmN1ZFiJIfpClf0L/E+gqHmPC5wcr3AIi1ZG
1wAMCfZfxyyR9FmONNzpYkuh0Bqaot9HHiU3275V12sMXzw33P376/VR9gXdenTVKPIcYDneiNeF
cEaKCj9adTePnFKxg1Pnt5eoD9q/BoVW1uhEPEwbPmZylCvKw/49IiwG/B5bqOXrLFlyk2Fqagvf
Zdfaj0idFiirZm8rQxRPe/TW5r0Bt26K2Vd+gbuiym1W915uwhlWMR1aECCE4bARinUtdhAcdWxw
gzKujyTL4KjmhFVzRtLSRgPxMYCmFQX2iUg8ZrZfLxJX1C70GM7tGb2vFjM68bFyg1HB6XyN3DQD
FySMhPSFNq874YFC3EDz9KKy0rXUm+c+xlQTkaThtx81t711i15FUPrBqcOM4B8JP3INJzWqm9ON
rT9oO2FTMZNOq9YydxRLrqlB8xAB2S4bZLbGCk6Re5aeLWxRZtPaO25ZWJKKQ6zD1p31eEwv5mki
8NVB/LjhetVxLrrzIGpC9nUM0lZ3d7UzvmY4RE8aLCcrGPNdBVxg00kLxfKQZCTjbVxBC27fpc3r
PLAkQ4OdH46JPep6YTwMVRbyIcYb8nLkkI5bbDupXZzB5NYQwKFtr2hg6148UwvhiG2tAdHNAm5i
YBINYoExEQBadgGcJLqSeRkMGIQYfvE54hqhfApLpV3FPyiEHhfTKoj57JkuhkgsUfVzSMaucDPK
STC6jnhLI6Aw8SEvM0Pg6o1UFqCNX0UZxlrVTE73Uoh7cTTLrLo4vo1sR8OsfKuoxMlAyqh3Eb2K
cZ8ajs9wvUe8a1EaS/aLCOoo5cG6sSB9e5saypduXvdluB3Y2g3F3j+GSl99ul/hoxLuYrrqV9ZP
5aj5G57pXx6J26978cK35XlYLixWU8FZ6zf1V3VEokf/dMInyxRLRk/V/b0qMYFft+Jmp4VgU/Rh
L3iB/BZ1T8mcoSgFyUe5/D+j4u7ZKFb+dwADr0Nxqe/RasPm5wAwxEkuD8TgXsHo7dYl3HtuGoOM
mLIfUWex3PfvBZQxaQabjKILV+W5lyrJZ630s1O6CiPYuKRPEVWg+TVrTt9UrvCKM9rkrWtxOung
drVi5+qxeeddLlzwtL495dmrRsXnXSHJXkos14+5fEJmcivPQtw8CYpba0VzdHV8lFlQQv/exQfv
L4zmjvhjJMjVifBx/A950NM9sGOspZ3dEeYTnyxcWC4rON0K6WXqDzLMtNP8Mxx251NhjB6awYAF
56MXXl1R/YBGGkCAa6g1mKOmr3092dijFTqLF7Y0H8wNoueU3HILIkf3X7uaZZNyZmW1VV5pZDA+
nowO7rleWKQD3bFs9uJw5b1wCxBpDtx71eoAEqBIymGpu6lzKrHmojc0GcpQoATPbOG9zbo8iIXR
oR/jFlXhE8P2kxM0h8KuPrs8DGMcnacJ7Wd0wkXHXv/uuOFGZBIoisQ8gyXjERY/p12jqXpbLOBk
OFGFNz42kxD3XRyL9NZgXOtFp7MMwdk9b22T+b9L5iHBj5Ue/WsAoG56R2t/xK6BdqajZ9Au0Xgo
CDpK2n/MH4TvXpoTHWE86gyx/i95gPMCOiUOb34tnFIDmXQdvv+e8Xzg2UT7CzGxp5ZpLx9sOiX7
Ojfk6XmUat/bPXDs38dXDhaIj7w6MdB2JRG2d4Gakxuq3/L2qS2ZQ5KIhN6MwNv93LI3MRMgh4/A
ZmVcTT3N+TbU9ZQMdA5z4+0pQvp9jWbsfM/B5hRTWDxxhvHOTMjjKu3UtwE5xjtVzCWrAc/fgYWp
jxS2f7Rkbw6/dLsoE7/Y6f0ao/6x8kJLnhYLoqO2Zj+V174Ngh4Z9eGkox+V+OJtdpLFNFgGsfvb
LxD+Zd/x/JK/u6rRsYm//pg4PmYPnaqtyI4y5SA41Q5GnLLs+xrFiRK/3ps5tx4tu3wfryBwWsps
qE1uuTcORkV0Pea+c1fdjeoO5vZ+xjoEwK5j7oh3CcJ3AiBmYpHuDrnfCZfBwVytkEZZ9MVMSFez
OIKevWYkh29ZoZUJ/Ty3IjtcXjS6AmIgzOtlhu2TGMmjL+Ih5Y8CIpmt7rBX4RJ1eSAjGAyzcJpr
lJ+iUNvJuKJ+IT8XSYlC00hdqQNt4y4ducQ/rIDOddJqbFTcynSbXCFPBXfNsc24DPIIA43VpBaw
PbzEpRvl8gaAm8azu2V6V46lYwYXo+eu+nHAKh8Vy3xZIWBudzoIhICPvs+b82xpbIHFMTrXORx7
0C6KGPvb3b2cQbAp3JtTRWxJTsawz1DNJyPZNaAhqee6ILawIrB9MyRgvZ2Tg8X4P4B3cWP1wQcF
Qhe+vVEZblE6tQb/ImpPHVPFDUtx6DH+XwoBLrMLQCrOgahLnHC2YuUdVFwDNv6RvwI4bn0WPQgL
9KAfIoqJbO6Efj7K8expvynDO5FVcs8d3WAznaeVzEtyXThemrGWvGf5fqtB98t+LXmqh012uit6
5EJQL4RQDdvc5+7X9knExrJMrXPZPAd6N17dYM+7E1Jczq2JpOKEQK9166BUo8dP4NCV1W0yhnWn
kEssBKC3pVvRgm20K4x2Biqiu3SfXgGXFpv04A3wKyB/mlweJD92E08WmYoJ5LKl0PVTYn95c2Ze
az8Kb0Kk8SLsHNq4qoY5hMLLRv0DSbHcQCkEsWkaONk0sY7egc50FpZkP26Yu58foaUNoNG19GGc
CvVt29KqYzvQUEN1WRcl5KvgDgWx+zRVwn79RsLTK1S3wFbSbdCFmn3oOc5R/7+i0xYfj5vPgeSS
cyBpzknL+QqQLdPVavlUxhqMDC8i1JHRXSLtJQ89sWljnSmx+BZzYDIRytA4yy4gcTrZvqmP1cqe
hl2x0RIOJmJqqGPZvZHx5EyH2H/X3TSIuaQT2r8QFQ1CkSd5KL2TqxUq2F3PyQUWbBu3xzO03TkY
5rfGxUKTDOMEUBjkaJ8ow08X0DiMWRtJwE9lRvIZ4+laeRa62YmRLFjxad//74f2CScQ7tIHAoZT
25QFajPE07SoGuRTcDvDqoK4ymxyGBjPf0SqqzIZXTsYx1f2JEgZxm36Tq57rWt6kVEqHFa9G38C
paXsw99DiNZTQCNhcIxlhqc1ei5Hmk1OZ6wX2Ihp3xpZRpRveNLARveE062wlMOO3MSMqtjii8Ei
WGKGh0nj2qpRquyYMqYz7TFdLYHNyu7/5jXR7dfI/P7VbEYGcA9fgJ9+GwRV9iX7TERATw5nAl6+
Yu7P5/9fo+mNW7lrquZ6zNKCqPzUkIxYMdAtbKH+pWwPA8eJpoAJP9ac48xb1/rJlfIggDiyb9Iv
tRpxVm0pSsPU980rQsnShyyhusrqt3BbUdnQNCPm84caMoV6ULAnoJzFizz02n/EUZg0qg2cKp6G
7G9hphwKQCecBOU6t9+I9K0YLGr10obFIF86I5LqkWQ8D0mlc2ce56nWlqjU/ItBNYnhMfCq7J5t
i2/vzL6GWSQey06YUDA3pSthUPJnNLDz9RESa/qTKmKlBrI6IT/2nuDn0Jsx8bdjmZfwaOaDbkoO
tiPYWeb2qZs4cf/MNu7D7QrZtzBN1miUkGul9XWU16mSuqxyzvSGgwer6EeW3U7mmFY0lXqtq0JH
G7Vi6NRfbZzg8WeN+xd1pJ+nCXINS3pslPzVWs3ia6gb9U2aMijNhqF8/MUwOhyhn0fErPT3PjPF
abfNRKy1N7Iy+MPvr/WMGjSr2NxaLPGuk2S4/tGxn3gdA1z5HX3cF/g03gjouMKq9BXw3Z3lU7Gf
F3WlHo8QNKg7LaUeSAHggQktq/wu7MieScbu8mv4vrz1qYCcDyfTR8YI4W5/J06vEg7/IUrRQ4qr
jUX7piQRIJaTdLlaf4LM7j3nj9v6RHtwLN1G7VuJR22BF6f/puGgCHEEfMaBfAn+idk3IaHLEPXj
YLzwaAwRFsxjPd2+6IX4HnsaeyUWeTvKLFSQ+o0JTaflDCu9oudSTg/YMGIO06t37SdPjq2naHDj
DRu2ahFNLP17wrGhBHQhSHy3lvMXP0pMTKLR8f6s7FtuO0ed6oRrjZfvgPu1UIf9UA+RNqs51WSx
TGJ2e6QoousN47l0x1+kKarVzDdY5O9TNTgqe34LC+jQ8kiX/yyU/dLvV9JqAJNfaZR+06NNE3La
J9NJNlDRh5PQj7qIo9lvhpOdXFfWk7ZEtxiIWtlDdgdQh9fBxL0yJas7DyNHNkZCDuTaCk05paRB
7B8dPYPLvIHYIKlZRuAlrDX5wtfXEM3dj89eyrZ2mg2OC6GAC6GUqpuMbFlgQBvxfg0Vnp8Gdh11
0ZK7VXhLG9UiG1jYx4nGeAfHIt/zssPe2d/BAE3UX9zmsh5SRDmYXxCS/ehg5w+aUEUVEL9GN7MF
AbNE1A72IxseQKEwix4P46ZBxvj7iWcDI3gbQYDtr/eRr6GYwgS4wtB9F8pIg/Cu1KOzLMTj8Hry
WWooQcCkX1ahDa8jRw9eFdXY90EBxuiTKwWxOV0mstnm7TYrEjksqX4ZGSXKumMFGqPtsZGwXXon
p3PJseefeEiS5f7R9etrNHv8Phr2CipWrzZk3He1Dqg98cpbaugKxRyAUNyvUMhEB8gevNfN69v0
TOJGkGvgfEKwEBbGbGpxIQx2j/LZlY6T/XjYVR1oQQlbLT1rbcSe2D7JGxrm1/haiiypRV+rI9kU
AElNTglCowsxX6QW7UYvJqlPw4h+HmeU/voZ2FnK/dEFIn28ZUmJCzeX8NrzxYK4CIMN4OdTFDD+
NEiRmoWu25zQpxCzgM39cSE3wjoxYk+sovT6VWTFTtxvYobT8d5iL/3AzhGhKCd5+9byQyKG6Yu5
8NO8Wu5/GqaXdBNXNEohwdvs+q10G9lbCo97CZ5QOccQ7rDXPQZJTgmAHb+QjQf8U0l5Fs6nGspS
EH/oRVpcnYWfjctJJKvVpcpik0m8bORIJFWnQUyOFYCAjsb1XUXZUoK2T0yeEl9usAn9H/cV3lxh
PZdntElU1QZG2w9Fqo7WTAAelgzuwpLrtlXzsd/m0bhoCOl0L4W9BtFZJobHH5joXJ/U5RbxXVLn
WnMXt/N6t3DkMO1+OXh9NxrYAgp2htWO6sgxBOpCYoBbidEDZw26VgmTFuHHMW1lMX2sxsAuTBmY
dUkogKd63gSscrPlxfKFyhqnjU/+BT7cV7DfrSyMdoY+2O0/C1qE6FqANf7DUxWxdFze1Jzvook9
+EMhf4DPajs9fyJ1WLifujcU26ymZMeBZp4QRXln8dS0gu1dz4UID49guOaTxOmqGfgfjxH9BUKc
e8M8YHRrBdgoQubXLKRH8GvqkTgl2x7yjW3ru3NeR9gy4myifvaaBe0YtWy9RpsJieebmwGOtGAC
p6tV2dZUkVTG4wdIJT7gwlypRo0AT+JJhrnILB6CA3YsbOx9AhzoncLTVeXvxKJoUz+Y/i9wqMyb
JL7DCRkAMiXeG9FXW+CIDXABeXSOOk32WL1pST1AJLClU+mJlNBAFBqSGbJSGv1z/QIhUXzCEITc
uTDvF8gr7yaANseErl35FgU2SGvk8IrgIWOzS5MNGDSMef//HAHmmCEt45mCjl+OgsmM1QFuJ766
dP4j3MOIbWxwSIbvt6T8+KJrVBiKmcpDwM80rfr47UBr92LPqwNSSAspg0b5YE1SP1BFeLkJXwuH
eF3dWxm5LKmP5kgqO0I6RNx+csaxF7jXn2+OExCrWKJ0FxC/dNgZTCprk3hjf1auIAvm57lupA0U
WfDHaAWLdSc2h0UxNP1bbCt/a/ELx7yuzFJrZHY7YQ6qBNm9i/ISUMlkVd9WR/WnOp4BkoJ/N16w
HF7Rn5yuzyO8jXZNB/4qjrEEiDPwfsjJwkWKX5NF2TNFNSCUr5+wtWdk6DXY53OTHBLp32v+QylG
ghEIAgPZFPpgL206VrCVS7QN02Hrs9TvpdUSUuI0i2aMVOEwNfsLaFHnhw59+Ra5wR0UAHtIMdFJ
wkXZAvKFGLmAcjlWaH+gZ+Rdrbe46dqI2NhJ4nO2wOp/hhnHbWDc5jHf5QTylLoU46vCOY8SbdmV
VeROe75ljubndNYgwXo2lYUzdMOA5BTWJ2vJA07PXo6YrtxLCtM0GIb/KHYv+27vEe7ys6SnBXF3
nkXXxhWEYgncHT1xvqnUJLpjbqbt8l43xU3TosxDLJR1LddNl3EGP7mkf7GI/6zE9pNe9e13tEfa
r3sflKC8fXjZ9s+xyaAMnnBz2Lg/fyU/ESNki9vadJ/d0RZMgVPzMt1Kxg6Bi7CBIvmv2Rj2lGmY
AilXbgraVCEv39zWa4Bw9q8/6pvvI/5r+vUFQbziu5FJv1qI0WlATYuQrc+jrPXFu7k1MygapXxA
FynJ4AiY2mCBcp9vOp2qZBa8JxVyi4Gf4G9zq1bZ99Wezolne/RPNKThwq2seYmtYJtq7hHMVMiy
ZhrD/+H5ev97i1hfxcHuk+cSc3Tem8wBa4MPOcJKHKkZSzokItYRjKjuqHUvT+u2YrcrekX97FH3
J6duKCLBnxd5k+BnJgbePyUMXCl3BeZnGeRlOwOOiykTw2X8qpOUAkDi5ZLrY5EBAZ+H+Z8znZDD
KrEVBFX93UkqWUfVvRx+JxuOPqppsbLlYXewSJ/XPa1zx+ed/KDGK6x4G4KJ2LY7EhQtpMgJkKzH
nxpiHIeTO0/z8lrVEeCIi21IF4sJIhNC0UNopugigpAjNUCMqSbjNwk/wazayuq31XRHd8X4H5M+
CR/BcBiyFTctZZjD1YYVDTqXRqBW0conYC89fANebJWi7qaf9DZx4dr525EG4ZpqyDxeudxWxj1J
hhlP5qol5Aos3R5CYz+Diilz5hLRHKgDqXEzj/4vb38I4MytUSLokibBuXUUCAJm9LTT//+aQWty
dwXjs/Eocu/1P9Tc4SQiXjSYk8+9/i7cLotzyBEkyFCRuBFAIh9Rixhqn7oUzWt6xaj9do2QCwwK
kdQuc3erQRUO7rdrRQv8r4hMVAMp6vsHAD3XJ9ounIHE6OqzZnFCtnxr7iEBfjYZREetTfXmvFzz
igwfVjuJjv/dC3nwzTMSTXlYyb5LyA5PA3BE/uOhHLCANqVCkvLNBS+l/v/cnrAfapS+Oiy6s3SM
vHgYzFUTP9O9igO9efh24Impwr5hYAZPWLvw44XwBbKBKJ6OwjaqbZJufevzAY23FHnOFsmEn38W
5kyAf2ECpN9br1qZcKXM2Iudbnyd0zB+8mfpvgRJoEvISQczH3g3nCEq1UloFujbo15QXJK82y3/
Ac/5SRfpvCjdpn6hAt8Xx3QGtDkv5oyAwT/czvL9Uk4f3/n/3y0gEIrJUDbFURZz4fjLPpyfdeHy
uoOQaC4elpHEe4ECMzvV4ECUhTckKoP7RJB2aKN4a0Apbl1sqGQX7qIXTuIWCk+HsAAFFl0mEMwj
e5YqH71JxKuiBJkDC19ObGbQFm21iJg+kb0VukzJbDp7jutwRKowKswAm9Z2M7E3R3YWpxZWDmKN
1irFu28SUz6JhfZfl/vpArnyPlsad0H25CAd7TPcDRMNZT8fIXGhDwGjy81eRkoIhIpoq7h38+lg
uvfwcNH5YOLeDC86+0Lqbk8+LIMBPq1gwCobFatwdxwARPZ6ZJ7qGjM99s5T1qDb6JM5HzimUC4L
UN7om63vIvuXSeraCz7hBsqHrlsKvHt9N/9giucJU7jeBuHnOYOanF1VDViVi7RnZPu4tuSuYNqN
ws8o5JVDiB1ZbYjPm4tpy/CE0unMse8ZLKsKmvpT7qalsJ1wa+zc0xw2vunNfJxgGUcWLrXD7YhI
Nu+Z+4a0RAa0RIo3+aRGSzVGKgH1kdqlogsScJZgT/IAc6yA/pO/q7umP8g6aAv9DN1L3JuVLRkh
hjj11WSJMxLjc/waiM+dR6gbHyN42OerxCCKT8DaTDFfiaLMkRTGQh4aBDca1GPZo8/DFvDX1Pp0
V4FlrFPVYJVd68Hi0GGTHrWVtgXV0QMSo/je7j7yBnUXaJhCK1+0eWR+5syl6i5IExgZXVabs8GJ
PhsKf8FYNkR5joniNb6xQaw3HOi4aEXlkRVmlRmA1ItfA4xrdt14+qADBV0ZKa2f/69CIXx/UoAN
fUQ6XQ0B7o41PO5xZJawjQQiKXPBhFy/ziaceA+RWe91xyZJS8mbVJINSbwlo3kU1CiyBn+UiQPq
EADPezkM8MTlboNxawB0ulkAf3tnYgsUAmUQOJGMUFKXjEKEIQIRNhu7n4j1JPJsWtX2bkaXmo3j
8WZGT/pnnuT5oWQaG7oG7Xu5SIbCuJw2tYYCdokVqeU0EPChkDkD9naOSfT1U/3MGEAMtkLHKQYy
K8WnpZSTC7eMmBzeTFglKQXdLZZ4J7L/WUjEjvOpwqFLwt2GcJrFA93WbYZw8ce5uMb44tLfWuAp
DpmRYuNlhTwcp7pQV9//YJPj/geI6MVBDdec2onLFQNvdSrYJhdh3Xns+kx7v926gOiD8V4OzXIS
nXZk/H18D0v+jA2ggA94VOwUlJtZRWKY9/N0VvNURL1PgwI0Dabtop3Y1sekIZC8jJyq4r4ujIcF
GrMfUq3NzDr33rY718qT6GUsUlpkLOLsR1Dfaef6U3gRbPXvPiEIt/7J+s1ZezTnv/fZXDeisNTj
nXdNzwRFt6L0+rGYghtbO4/2p/JA/vL4usQvhg816dXhkWBh1ZSsNtzNBluGgsFwYIb5uxKcEsJR
K3GaJUgOwWMvQSr2WKniPuhOshVzaIAbj4m5CwodrL9kmSYPEMVLZM1YI6khIMcu34qrUhIHt4xZ
HknqhautPwDyAuAbJ+8++xZR5/xDkZYxcRkMLAxuOZXhDnKjUhq6NHAd0AE9Cm3U7f0uBXoFp6/7
wx/SBBzIxDxFxaEUqCbHT3cPZFi4FRxDStN+/TZTOtK1mUxVPU7O9n2es/bYzezW38Hkra0BbKs/
WXjBd6h1lWIPc9bbyVjGWV+YR4SuOg9YWMvrO6EoCXU8/XHXLZt4s+tJDpnHXFVEWTGIW5PGmmXq
jzCohxCHqd6Xo1veeGyusuFB955sxfnx167XyDdIM+FEPNO3oIEMXE0pn/tWP2GpTaMssD1DsLlX
DUpxEs3iIiqI2C2VaqAqFTJuMR4scI8xc0NCN1oCI5I0SXGgbWHKs+3Lk0BJXcz9gwC+7902Doyl
sXq1Ur4vJ0noOG+O5VpRctxZf07703oNZYMkkWC2FcotHSlRa6fZoJzat6awdHCT8qBmBcCzls9s
ZX5SuQARZBrVwugmUA2f3+qHHkgnakl62UI22KJr4yGwulutfG2Q9g6GBLZZNqeC9pnCbSS4EHqa
OPOlfBLgPkAppFPz9OheQn+pXrtxymCmQeLODfl7HUvee86AS9nWNSzpGxpZEj44JVeONtlvQYHj
mcJ7qm3HG27Bu5s3wdsP9SKhw043kgTt3pRfkH5SOZFb1yGERIdTJz5mm1R93xBbEoA9nhS16xG/
P/WKorZEdTJ22JALTGdiuTx+T3cLSVY/oGxBmuQkcWlkkp3SkezrK3I2R4aIXEctkJfBJnZ2J6OL
uIG9KK8vy6XJzwYicE7+BaSDhXRF90+n/2bwyni+nVwAw2vcCOHkkWGNXCXHKvo2uFmTYPfUS9K0
7mYRWAjbvp1mq60OTyZx2wkIX6ndiq2Aw2w8TKCS4oFDd+IZs52kFUomG6ZWQ5/VmZ3KdzyiVEO9
88pzlutrmayxsYYs2cF/8I5Qc65KFrpKe8TE3fMazcOymH7mJUgcsxGipK0taNdcFOdU/iKgIJ4i
/moC76BEUjCyQYXdzN7V6QoHKnYkOpu2e5sOEeL0qiGwK+SDUp8SvsaJMdg7q58AvOrl8k9t+qqH
mG09QMGzZQwdbTFjZdPPZ5IrvCbhn2Vnr1fCUnFwtcDVjygoCurUK0hFrbhNbzf5Va+ADmRUhvG4
F5GLYQOSVHxaumrZs/I2GU9pa4GzsfDyKQETLDpyC1qAQeOvEJH4Q7KnVchzm0miRzlHItAOXD7T
FHNGE30GKWoyamxTx0EViPR74iWZEt15jqYmNM2yKLNE1jS4uaiC1+em8CbtpavNQ3F9KDd0WG6G
XL8pRLeqtSqmJTO+ifU3AX8K6wD+x9qUfd2G6nyWtJHQ8TKnC2uMhBjdfY2GS/7rJW9LNVwY7pbl
MrCPHqRiiJsfO8GxSVoVfKCzlIMbmBnqeZkncDDwR+aBAODmMtKwtwvIVYn4el9PcFicBeQvmPaG
buaKyrR8akt8jjupG8m5IFh4FFxDrD8XgfE2CAQAjBioC4L/BtJaLoKH9brbrULsQqZ5BJAI1NtT
8sevi6DRpa8c/uOnvLRXbJAn5zxj6QPx+M97TOwsalaZ+ckdyEPGTYEcvLjqHXJJlqr7KS16mUCp
ixsqEGRUX6B0KbROWg5IkwGYfNFgoZeJ8LNVoEH3ZhRAxJDjx69kaxkyMxLcxMkbdl5o7e9uVV9s
cM1JXswolRZ9AGCa8m60dhZTTTtzBxyugWLIjKAQgdcN+Lx4JLYy1Tg2LEZUgUY86UN3p+9Lzaxo
oaI89EormT93b5fQjYVJou6y1spPBvMr6g+0mhZmmNpiEzrgRKdvOHLWPHnolISE//knXfQN12ux
6RCOwWlNcdIL/A56jX348Gwsc2jcpVmm29xI8p9Q/7wQ0MGEdLUrAy5rAZXCQTxsHyj8fOM3o9Nv
82evsWzwJ8iU36E5tEqz2zgD+hadUrxspysTihzpay+wlt7bWQJYztL8b748KqzgviNM2vfxTOIV
ZmiUBda17wtOoOXFEas+F7cuC91vL/e6H2c31UE2ZUH8YxzQhGBRqlCvQle673TveYa7FKst4a4f
mF/Q+4t4qRuBncPWRtHELlDJ9gEEYYFMkP5VC83t0G7vSd5P3gq8nABr7mI69bd+/m62W8fkSbOQ
q4wjak9x8VmZlx+9xBob6E4q8B5adIHGeyibMHnAiUXMU414jX5ppUrBBnGqCZ07+sYabBwuo5v/
id4TibLwTdXDkWMlkJlWE0m6SaG9soJ4PeGTmW8cS8krbOVacuzcJm7rfaHjOTibI7paFX/wfyJ+
6tMd06B+cFfHyLjl2BEjj9YnlCoM3kfuw6R8QOpQ+whKP+MFw14AlUGbgUIsKYzHu73CR9755vsF
G99nogIbYaopnAplSHhu+pcjkdZCH/9cDnD2Xj53Gtl3+BgsX7TLt9w+TdpgGHws/eJ9uDWX2Sun
pEZ/Pd0dORGrf8elG+SQJoo8QDx1OzhjlGHT/E1Kx/RdDIodeknMHPI3G28QJACL4mcuxrXkb/q/
bEsMCjwk5jQSvcOmT6opwebftrCLmRYPwXyPYFWjTeEV7GuNygyRsS2ToSdftt+y4xEBQzc8X2b2
oydSfLfyAYa5omA9z388BCaL/5t+EkcQZITlFSMCxtv68O6BPlkGD8oUZYrANF/Da9Keemnw81OK
vxfpLc5MG6/mFC2eQV0MGPlXZrBaR9WUDBlSUUis63k/M8h509EQlKgrw0LH0FovmjXYC3X/kI6k
PG8AWymbFDr31phjISYMuzJIDsvN2wZJ2oP7sdEehqXrdRCHPEQqBWb4Rl9k82OffplN59Ub486X
YDKisRxJpczOTFc+4fkhOk5AuBHYgwcf5DjJkYdtcXRv4Tf5L9bLR5LbENBGypnRexx1jg+wYX6S
7yunKz2S4q5SOCA7UtlsTqiurlcyxBMmx/3K1o4bj0dx977KN/bjx9+e4gcys2nIczlKPBOVq1eq
pI1nsBiLo3IgHhy1woVc/u+eswspkgMbMwKbtLjC/aiTd+tL9OJZSvILoio5U2IuWqxN3CN17tpK
jsGhcrjy/ummJtkpAJ7iblUxGwPAUoqQkx0uAi4k4HqMWkEtuC4HW5ehDK25fMp+8Y+xTkF8vHz3
GErhPpMo8zRLuasrULsqrioaSsYO4wWMlfW2YQMDBwA/rv7SrJWGiG2dE8P5g8pWNp7vB29VfQT3
/F1Mnbd1A8aWY1D//OgT++qmSqt2cKAnLTvR0hNEMrOaCZCdNkZJD1qGH/1+K6fSFoxYMBBrmnd8
Sa7RTqdmtpbk7F1SXoBtEEYI4JS0HyccAGWbpsfyGJwDLH5wXy7P+LQDV2oNJ715KKO1G/0mM8Yl
HLXUkbUQYtOJ1GJkpy4JUfHEUAaCHk6/dkRKX04wwHcYYnuvYPEdgWr90jMyzvj5MfYvrEFmoq+x
3o2McJEK71wEu9eVTijkeOohfEfWD3WZ3h/e10nkVD0IAL+ppVLq7MwzrjvR/4hJspqqA+ecu9zO
RYeDoXaf8Ggx9kASrvkINdRKlWlSw3JKKT9n/DcFqqWQTw/93cZaL3dPuNyvgs/DYh23tb7m2Own
9N3hxOTs/Uxn9lGtOjXpKNCwUId5TT3HWDarOz9neYDIzAXLuHRr9bmB5el9xbz9M002aMl1SU17
79INpk0uwj83r6oixjxuzPtqXXB2+ZkrNOWIwPSOadNCVlCIiK4mbi9TQM1JtpIKwTz0FVUraj5a
9j3n5hWhNLPyw0HTcXpQ3KFKa2Im9RpCbJQc9Ex0D/pGSLYw9Ld0yXGlIjGYodTdT8JHT1RsTtb9
06xSLjMVVq6rc7th9sea2JEOPWvA3DRaVIBjyYpIwR0vMRmMTRBW1chcio9PNOlLkWERhl/67RL7
hDAx0yJav+3I+1c/gkemlVxvuvJ7BJLMxPZWxjlzDSSwk8DE1UsqAjJlWG9mxNzxHYG2jVVwjriK
ZKhn3LwUCsNrTc/RcBWmMpR0BbS94n7EvbfFtRSZFD2xthAJWFy3xwHP2an14FNQAHfHLyet9C5s
IabFLc21DFIADoJu4tf8CL0TKS/A4QTyvtuj3EJukkOwfDGrM1JZZYyVPCRhmyQjuiuFIMF7aXAh
XCc/diYc+W7KQYhzEVx5avZbRBJmCoSRY3F+REiXuHfrSs0z7IqubsLtKnDgwdlibdzmcoT64fLq
QDzdj+qYsCjg/pg81BP4xDL3BahBXLQEoCWD3BiAcFW0CLlAD86oFaxjVSGkjqLLohpv2AbzKASq
E4OoM8eiSQGDuXa1JPPf0D2MQ6VekyLRUbv20ip4SPsyHoXxyHrP6yilVN8t5rxXtLM+U6ZImVDm
SSJ0ocruOrCD5VF02VFJ6eotQB6XF1q4K4zUJ8XC2g7V3ob+neUnG7m9CfVt6Gssv4bqB5L+3FjM
rBOQQsTevJgEpK7WRB3EuzewWSR69sIR0XE9jJE1JubwdoHjKHcRxfomOPdtxtxR7ZFAnVkBl4J5
KqEfnj0GzklFOdl7ROrQhk04mSFQRmG2e9M5mi+u+uMD/P5zJY1geQxmzwCrGzcF+Zbt0aSdUNAO
4OoRoLSK/TMEiE4Z6Dc6uYeJI0xY940OxfUdQIJSHSrp9T2ZFx4aK/8kROLrxaa+lk4HoE6PJnjc
D0beaL1tMrybyDK3/UtJgFoxXx/vO6OtIlhL+KB+0foGJZq6nvmGxaaUNYEJk7DZFgi4E0yCUKYo
dbt1tJmlobidMhMUz/p7vmBxPvmo8ctYN0Li/SFWafvh1wJMmo81+pxmodDIRJrPOxWTsDb8j5Re
sIPaBt/StZ69M2BwW4PRUj73SK9YJT81QB7ru5clzAopQ1xoiOYhYw0BHlxv1TaSEBtsDTjWXiVD
/cUqOE194Z2wvtsCgWrwYkS7WBOob7lHJuUOiALAx4cECN7WDzbsd0RqYdcln6+wWP+8rFgSiCL4
NvboMdaSwGtl1Tu7bbI4xuuFKGtdk5jHU+QuZSo2v08p+URMuSqUlZT39F2wJmSpOnV442TQJNaa
9fPxfSWdWvjgjiRvWbmxdsNHP6uMQRXLTd9ceO+yFxxtQ3kK4ysvZlKvWnHhy7I50oBEqO/FM3wL
f+C2Y5yylhfgvOmkClwdU35HfbrMW+HO/fynneSUGoGBeQu7rJqlfxJian2ZYv6WIs0uac/VRsSe
lqMTftPDP8aMZHGSEtxvY1jIw/vTKgdubgKOfPXSIYiUMOvhmIY99GMeTbWGbQo4cQNfj8sJq8hW
NrLkCDzeA3TAUmcZuFhVK7fcEVibmBuFji4f9GUESISD+DKfRW1dxJWysfes1DtQyARtGRga4Um9
wRmeaB2UlOiaz1Jfp/ra1eEWK4+P/OhGqVOKb0iQeuiR07UHywpAo7UzU2HtR4pRZZAbG3gbxp+w
YLLaDsmBgF4x/09ZfjBonrU95IWRapepqVV1T/GYUKpay3bi/YEkd1TUwXINiGydVF5uDdTux6Mw
93hQjpyGBgb7Ac1BAxoSW+9XP48opqlk6iONNYQJp7Pmf1O00rk+MI1+lS9jcVn2b2iq+Npo56e4
jDO9qDyFtqAyGnfKGRlpOOxDqMG1IXmK6+azg7U8E05zR+Nv4s1p3/XiHy4+G1M7N9sqsNpAGz6G
BU/wg+lPqygpE/ZJY7VMXvBDDqdcENU+hf2mrAqSRJkhDsnp/r3C5I64lI78tWeSJG47OiVAq8Vc
fo9mwBoKzphhFIy0ydamG2KmMEPtE6r5XZg2QVzQRUHl8Je+4mIN7m/Fks2WKnGM50ooixXWiA2s
wfjK57qVGLLLZmU+PZm9sT+K9y3Jk8siV+E1VzYEDbt77ZoGwF1iZLyCFzpTf99fLJWi/W4m7K5v
EOcp/vzhqem3KdcNzjPh+jBkt48B1sCM6RfE/P/cREgWIoPgbeGXrshn60Icg9/G+FAFu38k4nc+
aLTckCzJDcZ2oueC7EltYrBbobEOEMISQaroAUirrKvRCpgrnpUus3JXY/hT3tDgqiSOZbkV/l1i
e2qp3pq7f5561cxIyAzlGbPM94hLqgpkKHk9c+wKeDg18rcywxjvguJoUSGoC9u9i1e5aQ450TtF
7sNQevfNqEs3uGfLpiBtW1Xi4c7VkcbElPXtg8PDJ8vu28nDax741FjKa8TpY1Iw2aBwgJNkSO4o
naw9MogUK3Tzk+Y7ZUZAhiff7hmvgOTcSNyKwOtBxRFeHQFUcW45uxbKGVXTXJM72gKLTblgSByp
3zSnqDY0Fli/P+ZEddP/hBMUh53iP0dx1V1dUyDKjjPG7ETpD0dul6Ek/7EbjM9YjjqkZsyT0MqC
XMFO5NtV9JGBAKTiNXybhsh1Atzus/m6VK9Yq8mNUz2Qw2YKMAH5tXeQqedVLdwwkgLv4s9xa61T
LqnCHL/ERhSRMzulBihfwFLhJiixA0gs34oHsoL+wSFY3UIoDgEuQGdXG7dZS8FzKs2ipLZ5laJY
Kae1PShDttYrmPHaSvh5IXseNcH4eeJg1t/fb3+exU4J+jcUvOdEOGHrwxdqlHLY61Adc2TjF7cM
nqfx2h7VvoTvbFmLDyiQsKtq94rTOmunFZCN3Rul24jfW+a+7a8ZDwIhVdl3a2VTK0igd2WEwt7P
Wb+VzhOhWVinQZTyqIyuD+NLMIjIzg2eFakR6eUPQNhp3dX0rfhBhH6FhAoxcxDjVJE+tL0qweaE
GvmS/OXDYGQnk0kHc/mrqIyUSXgabzFTPvUdNH9Jt4H/B+4GgYK89xkDQKkNy/10E343HrcQHNWD
h+Vb3FXjGQNkilo0qmdAmgOQVERxz9E9NgrfZjzh35qZ4IJPv0cX0kE4F+X0uGwHNg1KPrC7VLzo
ChNkiQoie3ITtnJoH1Z6kDTqMftEKesEbHrSxOfklWQVJ6pM06gwh/Z+lRt3o1SpcSL1vo17OCCH
I3OO7NcBJNhxB38SxIPFenGhTxEa8DWpJ/Izm6d4hqPmFX0rM9fY97F4dvH7gON3TAjquN0/5wZu
XatonOscGo2FbaqYTv4PjBhgcSRvX1kqDVPQejecANtsK6M7VnS8TIUIJM5ujgrUK77nggKWa1aM
yjhdsPNrpZ4eBW6O1M0On+xDQ48I4f3yCI71ZkWbASXJ5EhlrgtQsJ4SdHZhtgOAJJs+CW1AmAa5
aezbG80W8B+zkNP+12iJeR7F9kWwYm/HVNQ9GvT4r/n4NrHzT/ZWolzR85PGqGkFTv80yoH6OLxH
0afaEjYRqQDTYSyPpyT2scw7i9BM+u0F7Gd6kKauL9fAbTyUbg6YhmzRX8XyWvHHpmVLDs74w+WF
hNK/FjfUfSv4cdt7VIIh8jieTtIZ/n79/AVijgr0C1ExerV3mD7dgo3AAApmj6Lg0hXeJprlnOD+
TbmSb74eBGOK5r4XDlCi59+NK+MfL9DqRNvhru6292kvqgAPCK/AonqEDECax3k30+do1ndP/beE
pfAUkxAomnOlFGpSZKLwjb+d2EHk6lzgnejy/r+7IfrYRmVfaTAKYsYiqPvTlP6kjxI5aroH1AcA
+QOOOGPRmQA4n8KtUiD6+Ladr9Juk5zK/yAZzAhdVTaC/Oi7jtqGD4imwMnJOqyLt+VgIUGeOLWA
5eDugerbhKlWTZLwmhOnQyTn0bWIBE8S3ct/3CmoHE7ARSPcwLOAA8yqXLKMS5WBjdH+sP3md7SJ
Pooh37wsVXZjnvzVYRnRCrOJAWk2Otxu8o+R0+IzUILVJ6dlZWt70TIkYPCtz83v67vUqKrl9Dx0
atzbtViljQtMjmX3Lc5qh7DiA0OpSovg1rZQmV17WJ2IvblmWDKnnbI++vqbgyCg8d1CQKsDp7rD
yWlVsoH1Mcau3GeDfn4Nt7R9hStqWhlxaJQ0Y6S8xzPhEf/58aoe9ip2RrG1hSCmU0eqQeaQLhlw
dUZWknyOi8YWm33NoJOCNpsez2lw6xSn377epa85aVaFERnZ1/bETl0waLAH6CZr1PLFJcTCUS6x
wo0skSPNGiWek4yBFLnp1zDGKMWKM8mXm5ahYAWVrkS1fLoNDSPwtCsfC/68B4zWobJuNtpL0A6U
wvg57bve7o+KlShItg/YB+I7S688TxYo9NMbO8bUKCWUSj/6i5KzoffoBgnCg9CIco1w77QEi6O8
e9fMLKXPTSxd5GWFmdDW82ucSw9Xlx3GgoWIfX+fEu93chbEl75ETjN+72H6pnC2So/3bep7WA0G
YHZ+uKfyf8wP0WL/uvG0Jo9zH+wJc+5WCxjlgAPffPy6XbqZoppFwV81g5NZLD8tHUoGVBsBEXbt
c4BlGJkGhhJLgroy7gskKJyN/HGGumK4USddAvfwU2823hCHb0SkaX6ibpP89UVCFu1Vc62SMf3A
BYx/avFMcVIbQtgBPlQyWCNxCCO6jmWcX4mmyGQZOdIokgSqEeS3DN8tKwM/tgeWZCZtRYIS8ivD
1PONCrY3AVHEsLgsA1KfOCvu4RAvfX9vwHkxh2Pw2L5twLLDtkE+NQ/9CI7k+yhPjwMha/yKb131
9pyUgLAyi8jGdieWo4ZtIlb6sWDJTksoDjghxOeqaUaUOOQu3QODJoGOGB+6d9MvsgBRuWSQaVu+
9WRHnmFNNE/uDKXRk5Uh3Zg4aHLxWiMkBtpng2yAYfXEOso8ijauw1LFbptWUMl6Zn5OZMN4KBcW
maOPzqCWQzW2keOtGaGlqfbHjAEzFeShQPLJ7D99QjzBQVARvCXycVCSNmGJLvb5rp+fjznnmfWe
s9KBkkb1OVBAzRSYs4YSm5fgMamtutVMldUeTNDvGHeZtdHzO1H8ggnjzbPKWF5QXMNnxtvb0pSP
5iurqvjFtWFQUM3SNK52zeIEvDFFTjxqjfjIshqIQCVv7cfw4oeYbMIzO93VLFYMeeTHzXdUfOWg
CVRbM+TR2GliWExT5Fex2eSVebE4tz9zN+yPW0Fbi4qh74cstbtRCLF3NuACRM2SwgFRK7farCva
13Sv94cJf3wes88QPscUG8FhHU8+mqBYxJLkwB9eIgpWpF0jzncRq6x9TGzxK25fZ42Z/av88ztw
LeYNsLLB7DnoFK/e0qX3DWMClQnOGBTea2h/kj0mBVQHSITem2qFneJrMyBEDraTCbIg+0IiTqcO
3n5NjsDPP70Qsk+t1mfNQMu6iesA3djwsJ6FQOZ0A0eiW+6iXhuIfjqNlqYIm+L1FRhfzvblg2TS
tY+Ne8Xo+n2neVV+tQfOhIosCV5JbBeh6Vdven9pFpjAuTabvYzUYyMery1RGJwfNyVMGUp/cvF1
pzkkH/zUkWwG6D2qolBymUIL44FJ84/BFLvEbdrt/GbtZrAIMKKokkmQSyph3PfhYpWrqI5rXxf8
kpNPF59SAZFlMUDAa6sWPBoUUNUhX3sCS9p877NPM8DzEG0w509Xj5eGsp1ZQxTEnckYC5M1J1rE
mulYP4YsHT0n9ZohYX8abPDqsFs0TaqQSaDoHrS/Fii0uHc94wWV85d7RCqp12X3zoyCqYVGe/EI
A9oaLD55R1biHGtkVkaYPVicr1kIrnrhd7l1pOkrrUGK8dT3udEZj/vFlEUu+zqHWXlwXro9V6gF
1Yrzi3srIeRI0hheyofXt3JkMtQJxN1TsYmtxcR3x4nv6YCqOPk9y99oi7EFEG6wGu8lf65DkLdF
xhi99SnFJ13JtVxdiB9AmoCg8akz+Gc0NjH6EBB1omaRBD4zteu0wvHKLUA5vc5BUbPlF8KdDc68
p9xB1M8ZWbnxdLE3zT4hAFAwIzeo/G/kpjWVHkZGXBsCh0t7X3EFlBGHyDY3RnDXETAuAeHJpuM/
hdGygItD1ArVGazkfM2SD7Xbg3zHwwTNR6ukNn4zBd+vepAaqLIZC99t2ubFLFmqyZgZQZeDqIOv
J89kp1af6Hs9DMGZOQm4UQ1OIgFTJTbua2n4wMkVsTbE6ibovCIDg5JwKzvif8u6jNouqRzTsg1v
kVUBu9e2a5leCAEXY+/oadDYJxoL9kKBS3VjQusmg7jra4smwdCVtYNvBokAHKtBUF3L4S4o6T3d
02kNf6LOgS2zeZiH+59L5XZsWCqKN5ECuXPihFFb5zSoNk2PnuHtrB21ZKMMfVsn3174FMmeyLUW
m87iI46VEyEZYLomC7GuycGkwMb5no+hUhoRSpvoejL4pgAzVSlV8lUHkq6HDknKw9p850Y/H2Ta
PzrOfhhwuVy76nGLWZEEgY/3rAABzosWX8fK6zYOHVXaoVa4NEZKrnFi+pnNBM1gF1lWXVZuSkKy
MDwJsUmHMKpdmfMYy+uXZB4sBYs1gdMYbMp8HdX8ZvIugXpIPmav9vxZlB6D/FQUctZOa3qXn27M
/xGzZSw7fqAxodITf77uAVzJcfT4JSkd6R6yongQ+2uqoT6ZqKArFHd2J4Rjzm/9tlW+U0JwP6yK
v1jz2+/zsXiBFjte9CpgUtRUb2O6RRvxkFqAbn1dlBVqbTBlG3GGKDGNWqOKW4ckGKEIKQpRf6r2
fgkvhIKcPfKF8MSCN2qJ8eVquShIOLDTjl5qKepoqD1agcy3wjCIrbX5FND0G4vu/Yl7TVEQ/YZ8
bZg6E30OIfRJn5UCS2AM7AoQe1aMweB9yXghN4ILx/RvE+ZRCBiRKPR5V4ybn5ktq9Tw/H8un6wC
u9frkcJEj/hc7Ll/8+0GO4lNYWYuRNf94ONlt2K9iySs9mJl3q75+6Y/NF0MYsnUjAf9lIKuB4Ir
0uz7SaODmnBlWf0YMHcoerdZrAx4C1YRlnL5NwvUuhlviAM8zwjJQgq0lXK2BRDUGMkVGW6OzcWf
Gb/iaAWWfT9ksPuHrjn9UARPi7PulposY2kkZ+DKmZuEIIomgbP3/iNtKtUOkdJp1zsO4UViLiQ6
HtYbil8myWwe7CMVxRrnsigw1sZiqOrpzGhNesp+fpSjPyy0coTBwt7o3fJ+Rju/h7FiaVJ647GL
l/5a14HPO9iFRxaPRf1IlItIbNqDHo/0aLit7FaIEIkqaXZkY61jVcy6EQaiTRimAKqYpcsTW95d
7zf7CEMWZ7KkvEgxid6dbuXDsmzKbnZh3UwFNTDEbsE3TDrd/mdnpyBs+EYI3k9XmfBs2ToNYIT7
ZqCFTSjGwNCKU0RrpdV98RP7UEeAUTtdIqcLiHk+4ykiQYVM2olP95weyletGT7/685VEEFuSEQ2
UjxBR1XG9/xUzWArD4N1jD8JMDfdZCsnT1kCYkCdGPJdVL5hRIX0txQ0qe6Ooq5ICDg+51Rg6iJF
oXqvKzBSUoO1orRNcXodTTLzDCoH0wlEOZTdRYjdNef941axFDob+1QFBE3dJXCG/NzZE2OvTi0i
kdC8hKDQswRbmiSRzvFt+Ths+gXouXaJwoAMuAGpvXk5jG4pABaX8D7VY0RZCXW2fYjwNW7exncz
VqnweQVJP5YNDtE7UJv34kzBQVHWcQlGT6oqF6YRw9JGDsJbNxzMhTjmGRJODEdJ8wnD0LyW0j3d
CRNOPUz1zloQSOIqUpKZrhgpM7vnEY67Qi4yP2+E52/ebzqUM7oTRtRx4ANtZtMaYrDUeD17I+La
ipaxeu736iQEqCZZgTXQAzCp6ZWDLNILZlxu0ZbdjiGm+EPs2rVs4Zgh/a0thGn/cKK1Q2xmqiZ/
5++8NVqLbMeIau8njsn+RwNhUxvj92qbKCMRwhq0St8JoSzWzOn4Z/PaC7DY+OQ53G7H/rBVolw3
ulpjyBs93aHU37yv/suKkqq8+1GyswDwRwNCuOltW9Q3pwQFuGNWocOkaBnBM0/JsKceh48vGL33
1dLn+wWalTKyMLcRz9gzlAZiwfkk7D97ZNMmy9OSeD0A7YkNsUV8aJ+54G55NQqGXVrMfJphh+pi
IujCnr9oyW+hkiEQ4qvDlmWKhPReCHWyKbj+fElBfRS8OuO13jB4PitLWB9wuhF3CcY0O2VTgPAE
vw7P0NLdhuvgE5YT1UIfNQP03xw25eeKw1FC9YNWAA6KS0rudkZ9EumtaSCi7hlSlCLSenh5acM6
6yBLQd/1KLirUG5IX6PAp8BcnvvtyPRVBNbctlW/YwkNa8MHMEIA0n5wTZmx7nTy9jbM4tjSxPPS
/1QLDyYNEAycRnGBnLjh3Mg7CaDmNoAN9T/wTi788Y/xHpEdcmtDMrTdgaqx0tr2bFmfM+ml2uCv
ylwgWVTrMwL/FswMS+JB8FW93DN8Nb/c8qg09mntUSPs7mCIUKjU90QhfcNI/C79DE3C9SNWdNqa
YjOqftwi8TjSPsJJIXfyxRfEgD4qRaR70HrwdzGqpLIgPWlwgRuIFh4as+o0K+oSA/aGhhPivRAf
5/UGTp9HkRXkKXb2TQGlmjEykY03as3ndIvtDycuSiClF7hac5KDEBN2USnWFMPOgmOgqbiXnXjm
Yyinb58dAjUJmjksNjYNlCkIHwgS43ZGS1PpN65z2qfPO5jZAeJZFfS5hhuzOIB23XEl9I+DiNXv
psr4v+OXhGFL41mC2VGU2sC7wlFHVRg0yWHFS2efbzSAizDBHCJ+YVs8SZ8wNaOmv1L90582MGuf
4pr6XX/SHEPUlGFaIOE07gvfWP9x2MJ05dCxBrhUgae8OXQOmZFpVjIX5JtUHfZyU/LcN36QLT4J
t5eLljWq04leSzX05Tu+IJ1uA3M15KNxixtO0CyJG5EPjyRPXfGpnQG2JdVANJxMNB8uZn/JxUtv
yqd80xU2hz+tv7zR7oCFsuFV9etfi/Xn55pV1Sr5ghndTj61XIPzS0m0hbU4jbkL5p+f3Z8VvdNA
WA54/9MCaQIMByAKr6A4Yg2E67L7DPfLedpadVOI6C6q7g9Vp+tIQ6CwX+GL9BrXsYLg3b2KNMqf
t54PEVDrUYc+zMlK2QoV4TO2kPU0tRsCzWNXU6NNrYmbmeE0oEPJ7jPk1tPcHjpJOmBzPKY2wlB/
CCZtNaHvpH1mqnOPoJs1Ndr3xhLmi3u8js8aWj5p+nB2sMTv3Sfm7DEcbV69TGU7r+kJSjrVDoNm
KaiYMlVmOc4MDzAzs3uE/5D2VS/eXXsFXKymsNHVV9578Aj6jfgQj5ISjrfqEZtQ+UT8hiYf1lvs
YrSqUqlnsf78f5pWycTRlOiZzBjgxprVHuyEfC5j/MYGKRo0/8jmbxhqiw50xNM7K1ZFxabyqf3r
kmdeuL7zBLAkjbsat1xmGZDSfYP0VOXOJlCVXbH/BOuKgzJGGUFv/s9vPNsZz8dkwCR2DykUEtlR
oesSo4AzfkJccSm4iVNSgSt1ur0f0kEmKm9UXEKBuz+bFpnuUdchlk0XFcsQP5mQ11Kg0krfWR28
WbLtA81RBmbXRce9fUueDucm18cuuJ7R3TCNUAItbWrBGhmGq+PLu/Emf0Qif/8NlR4rF5o4Fkqn
YcJiYo8i/7CJgT8NHSaeqG4W5R+bxMtd/0HrApQH5rrRpck2aLX8OSwImSbTkz5rhSZb5wDCegkR
5gUErMqtUEz2Vnw5VkuyHLJmmO4obwVr5ONMsgBf/k2eLTbZWYTfkTrLGymsndDFm94NPgJxDCUk
RFDuHGU+WdTCj4clanu9Q7Z+AgIfX0iz6d14dBPMLUWGjWjeKSAyiON0aMeq2Fy49dXtkZGtYbaQ
sYoczm5AnCcJ5gniPSukTQr6MmcE0Wi38gMOk+zhaktvcbhsqsp9L6qosV9Prqogg/4HRSk6+gMx
aDv74x5ODvnemXZsNNoF2cwHds4zNb2jXL7rzNXWPvBFh5yQmOygbmmvvVQNzIj/fC1919tZWL/0
v2vOQfAkC4zZL/Qmy5MOT2fOXzXtv+jXne2QwmsZZp5xegT+uxsWTWnQSlrGHEAOXdfqnDHtIrxs
TP2DU5+7NTDNU/pp+gA6q2ADRaOmYgDXMu47/5DUBQtDbEAJd/BReq9XffaL6kZAoFg4IjBEyF4b
wNvHAjDFzaKwzuAUV0tnuB2lmZFFwwkj6NxkZZCMrCzqCD5gR0MuvI7CU/IINkKP298BFyULNcEG
dI1nKRgKsPOPJti+CLCqwDnu0gp1y+hC1UPKwUrR+4GgIFJCOEbZkRXUVyJR7icpZeikw5aOsbPX
rbWR/s4THIXdVe3G5equ9r1ra95zCXQU94911YT9FcdcloazgiJmgAGbWiY86KE/Qt5UkQuAARY+
MqvUHvbvmb2CpZvROtnnwts1ZynE9YKuaF9rCK+vot9JLUFdzZ7cIAj8V9AEIjTr1ASDf8NCgyrz
2NFQ3K2Zp1/K6klHtLukWB/qUWKpovK0Dh9LAVBN0VIuuYJ6VE6CbP1ZwHdcUsY/4KLJo2FnVmdt
1AT1Ug598MwIpOyrm+YxBaTtEeS5OfsPLygTUTYCEygzWAksskeY0RxSoBW49pryyGRG5Jyg4CmI
GMwZe2ZE6KvJzVdmNsu5SydXOqfU6Bys9T6gyKm1LgE9YqV88izpYWoP44LcFLvj0w2fGvmUMlTL
SKWutLcQ8UywTGnD3z2xWSYjuTCEKRMNEPlpS00GFWCo0Z7y3uzwVTvBqekclFfZXlsNAHKDbZGX
l1ZvrT7UPFgp6YIMxeRvHt8AvYfCFtEwMwPNsqIHPfsmPmi1Xub8O47wIc3AaLpMsibJBo1O9ROY
gvCtgxPPw+8QwUJQKqfFExqhCsPDQAC+CaaAOKIF8wi3hAFqI0zDg1cMJL7w8VevlDuk7YuQB+5a
qf8CLWX9l8Eyup8jY2bY4ZvDZ8yvdZAsi84R5T9B5HrSM8hQS+6XfjfZ5pXk20Duc/0nmgXye84B
fPc4978PT+peHlgEwWLL0Nlu+5mxW90aiK6yc4vEVPTv5V0c8bH1ntSekJcmHYM3FNu7/3hxP1PR
/CsFEvoEqNfS4YGqQe0os7WcdgumMLLcsrw0LTJIIehfjuKp6NTmpaizno9XvxyrAzEoN8LvlZPJ
f0Iscw9Cnf+NtQNKIzBJdA5VPypOyE+shEnGUHE25j8dv8DYraXYGxNOfWZ9pbWQxD050FnlMtXl
TY8Q4WveBhKYfEcJ/nwJt6wVMHzTkouLOOUESOY2OuyLJ8sC8ymZza9yOQCk+HDD7dw/UkWZIArq
KWbTxpkTSpj74pTKgpNZcm0gBOYQaXRlgWz3SUmrKqj/T+3nV5vNJZw/JmpYba6hSTrh7TGJYO50
cVlZqHQVqXCUcRZpi7xoBdWXQV5ci9UVxOG1jrAIZdc52X35nHDgv1m8wroPe5R4G919H7LKfw4U
I1ZLiWA0oOHTpxUe49ihUt0kVIcwBPzRl+cmRKA5A7AcfDLlsxCP84T1UsvCchgMcdVvPGQWPkWP
cc8Pvuu6D46lEBL8MeaII+j+WzLi+aqcKEXywdzsVpT8MhkwE4cuwl8X24rl8bwTZjWza0Iwrfit
GVOF46mtpLOoGzEQzrijWVJMYpGsllCTg1zoiuyQNv5EzJd2NBV9fHsFG9fclB12K7COBt0fQZhd
DU+VC+wGDpJ0sAPDItcf2bc1fu90iazgSlgl4E85V+bz3/UqLgDn/CihQJA1TfmqKrakxAthR236
qtvekAhlPdZpHblhuCm23788/G8LBDmCVRsW1PUMffMq6rPOshKmB2qEjMBwHe4BpybIAT4ESn4V
m0GL2qT4hQfWFSgheXy7tWMsqqujnPlOQOsN4EHuQeeRSrGBpNeBozafSYwHO//+/o9s090Niu0q
kvWBmV2NvsDEC5HxdZ/xhNgLCi6XUien/9rPuvoQb6O//jI3jsKpp2D833HjkT/Bg43kEF6cCGos
k3KAAH4W8DHNr3pjvVIYBbEU2gAeSpq24q4DsqypPE6gui0OXAAV5F3gLOrQ+tjoak3FkB0Kj/lP
6H7NtQ+WfTZSV+xHsZMaVAdOI9XdRuQkp07aY30Cm12dvRCV/CFYLT678BnksIVONk4YuWGGtErh
n/q6LYpbDZ+YTOmFTvoMeqHHkIFokrHWUF/qyVVbOphLm897J0aOSCUbbUREUISLtQXtmiSIck9I
fuND4XaWcdyhOW3XHPZ9NcofTbiaAlGc0Z052b03oLQPp5Gb29c/paDJ9+768ft5xR0MarHSVnu2
c8XKSaRrFiHonhIaFcPrqw4FPb/DUjiOe75+8A+k1Nya4bPMHIben5RYl5/j61na1BZ45Y1krc6t
MInKLjmRlKQvhIFHm3eq2221aqskWLxo7sPCNojJsI6JAu5IceRMH8h5EA8y0vVUA6p0opCi4Wgq
NVwaaEocUxYECkM0w5fawA7u0hshesOS5Bfb3x4jzvjjQ76o9JspZ7s5oo2FkmVpa9WTjkEoUXvL
+EPNB2D0fTy9e9DshvFk5c1hLa+LetnBe5lXu1Ipe5Fk+0wT3rRU7oqP0s9tH+uocYw+wyXPgecJ
yo2cKXn5vmLgqm/U/iwo0wRS4RzF4h+DoBbpTkXmZAnkdLNurtvwWXMuwdJmmgCjZyij4jnoH4yu
LgZmH/VYgwP+A2Dp0hRgqmD66xhAGRy3PSYUnooPPvqPmmPliCewBwC0qyPuPHnamkD0pdtiAzFp
Eivpm1M+v1RWaQDYlIhwzQBUromv5OgRaNzyxMsAN2HIpBnID0LwKL8awcf5z6YCi5YdSRZLa/ec
M2Y0zGr+bvrZOtWIAocarlWFpGIeSnIuzwmedNzaLG7VfMpsze87xCjhyI/CAqGs1XP3ru0BMyHo
RyW/kSCrYFbgxT/m5Hh4A2bqF5KqQxUA7E/Lw7ZJTuK4xZykytaFalTwj+/eT8p3S5Lc3TWMAzlU
e5OBiHUYs19hMtoEHquW1WuoR5mbmBr993Jb+xhAXmt1zb/a9uBvsv4u/GtYEB3FsUZNl4IqEfNT
YGzaV3+e6Vc3/61yCknnV0c0qMerX3PkYUryJU5D4xn/uqyGin9qvAZqJQ/5WAc0VzyhQrNwVBoz
bFjnJAQ3mhK/14fKsnhFEO61Nc7ikLJUlushF6ZiX7Xx7jztuzu+xzZ0h/fwMvNHSqHg0xeJVUYI
LHarH/LvIhos/9KdCUfiXZht3q1VfOnNIeK/UQU4HZpBEheu8u1dmqdOG3zFzHuQ4jW5AK6gz24O
yESCceL1x+kLKsqNXExyjTIksy7RpKMvneJfcRjHOv4MOmzqp4qpRg88pIS3kybj3Ls8Jn6uloR7
nOKmqI0u1lOBNxd+zd6CWlbxWWfKtgEvae49bApJp7WdCKhh3eHoKbOvBGq27UaOr6jkxbNhqrDm
bNII4VCwI55GoAk4U+SpT9XpeiPIc9LxOL/GDY6vV0UMmfk0dzJLXK0yMndNxIa/ieFlBeBZD8uB
mRKPceA5xFi/v5p9repu9qRxElyei3ZKLdwKEM3qtcBG+IRViNdi0PtxXO5Y4O7e1L2Giaq28bwu
9fxEavflY/UmR/RpgdXBqcqSdIb1d1R8uKZiD+QpJ2/30pgEfKu+yzLmZg3VlgVc81g9NVCPx56o
UKYkng1kdxJ4Jw5M4pl9EZpWTb5XCKFziwjEQpWgJCXuPyH8l6OgwP0puNiclNYzHyN7F44nus9D
FBkFUZ4P8AbQDXdP8gKSZakhGv/XP6RSXPiBtjRK+FFSaDsEY3FQFuCDYD+xqmjlBYp8Czsk/8t3
H2wn9bYpvo6nq32tn/odZ1rrGfHXRWOwKRCqQvnBMKNk45Q2yF5UodbWAYOcd5MuVTi/BbQy3A2h
CGCALtc5EZQI7hwZjRcGVIlNn7DHa719a2yYioDiw/x4NZ3jSdPUDZBz+0LraAfNwpjBiK03L/2K
D/XUszq7eOQLyH5yyPEKAqY/wzQfNqSuBOAcLp9LwTJ7WDkF7zTevmZHtxCFG8izxiVb2FP6ML4g
6ioO/2Zt4TQJa6ibXXSJIf5v1iG8Z3EF4Ajt9aw7p9sCS0/1044igiTPSQy6u60f3/PlEcXDSlMG
rvuaqDw/+7HBQYfin/o9GYMGkf7iq0H91dSE017zMcalsa09KF2pRN9J9C6zi2nHRe9ok+AHOMYd
aUVDYrrZXWlqJuvXCrcJTgMrNz4gKeSOrt3K33ZpaAM+TZHwymG6zzCSNxU24LfLSak3p4KyXKdq
4GvgcE3K+w1Zr9beP2TpidCdTFJsFMP3usWORTJ+brlktLDwO5xcFjLZxd7B2TmWgi77znRAIe1q
XnWD1KovkkGTgTuCCOXBRekLXCSCYJqQrcIhGzyMjnsy7PRwX2QdCeKzFqA+YH02LPFDq41tyLGc
3+wOWglRMUrp8XrZvSrOZ0bbfjkseWScIpJq0HwT3O2nlXtsgU7xiXafwiMrI6s/PZgMcAvYaMnZ
epaVDqv0+ddB90uBvMshZdCELaaLrytt9AQBI/JWpg9x53fYw4efHB8A8Cn0dVzR0YQMCCAULTLi
jVhOkr72yA/2DdN6dd3shbjKOq8t/M3gQNgvZXwsLQRp4qD+7+trUhReVzWhetGcEet20ETDybbD
3vd87MuEtRwqsOiXfNKCTFDUX2CgcLNZJfwnMH1qsvaKTa7EdOlGODLxIe4eeVvVkiTAIIMQZV+d
feE4rk+zAwLAnQ6YnLw3V+XDbF+hDzIkcIUIFK0r3jQ8XyV72obmv/OD70xTDTEv0z2K8cLbOEE5
IYI7FmqrIXeeFRk5JBtfFwbRLehecAlZhbiweB5waYgdXW0gsNfwjE5obJk3ElGbP6XQlPOv7T7w
qkZcpkYD76+44411+VJjxS0mOg/e1K84QF+NZhrSkT7X6TceJhU3aeopbNH58WpsSVmasCn91YHk
s2sC8vahVtLahRnzFDyhvRXvLSmO7qgMxQPS7NI7BkhTOnJhLB405ebN7iXs0nIwuwE84uX/PQXr
LCv4aR5EwRSqej+Z4gOehu7AafwNKX8bkJJL507wr2i0Ook/G9MR0S4FeLqDjNRJqWxOaRn9HLpp
XD5xFuuWLiPeAnQaUWFm2zGT3USntLMvEyAUhlnuqB8b23E5GwdO8zI/u6i6PzwoXvJAz3fo4sDe
06u3JpnTMJEKlb7Oo6DMOQcqVtYkrdbCCkY8PnFV2cF0IIzUtLqWbfQRHRFKMSxSeHV7xo2qlVV6
E8QAfLuagSbIURILj0XTsn1M0jeUksZ73AoYdOCpfOBCMV/l0p+krjf21HV4bjBskiHg8ONClQPv
nbUscqOWAZ333luoTCtwHpgD9CIbRqzE0QHXKg9puGFeFqVKiMh5yZhqd/ZjFvGDoyO3T9tEj6zE
By4AsbBPqvgkKw9hKPyf98p5dQdb6RA8DDv7s7HEgK9oXxyvk6qgy3GtqvT60B6fI0iARTVEwx96
pr8u7XmH2137L9dcHv8eWjqJ1UCxX7pc0l5i5RYFcLvWsVM0kqMYWG1Ozxy3r+96jkU1OdC2r7O+
NJ3mXWKIC0t6SeY7zBzZ1QKi74vmEALqADwYtJBy4CLQ4cfVZIbjQLmSQ/6S5hc/uUC3NTADTeqJ
bLeMfhdddBxxREnF6bV+91hPD8udoJw6zmGLt5GuKJ/Y0nNiw3w+txu+P3JqpqdCcUAoqBTYnf7M
SXmMtMUfHCH0LmJQY2YDg/67goPfaDMiLsqAHABPLEAHE79w9sHQUrRcDl9E8pJp5LffU9oI63KK
JKS4/K6uX9W0wR67BZ8smZU/nWVq8o97PiRC+X1FOZaJtJ9NvarFUTd635sqshRknJCTa+3jjVCZ
oidsbCoX9dT7AZgIrFKhsOSjhm7AvbXTZmK26HRhyDP8edDarHafcKaoTxGPz/aMMYgjYWeyZc8t
e/tRIfyh9zX0i0txioBReNqIQfHTRIFvMcmxLC5Jjz1KRYBDYSfNfAUuCnI8eHhONd89JuPl2RhL
3OcNMrJo4plk8OFyierwj3LQxwrnhJDjOfr7OKOWx6WatNTlU3CUJwhNPO3niaa+p/w1tMX4FykO
GwPSOE96kky8ZzG0By3yhdztfV058g0NCO40Ka+11ZEwSUHjf3kILSFze18oHINjQ2bP+1d5El75
p0LzExRezvDEuD7YTnFaNc+aBuH7TPaygdIqWmWlw/ixOzQjmKP5vl3K/bYw9UNmXpjuSvzkwv+M
elAY/PVwtdyajx25bThxkLiPsQyMol5OEK+khdlG66A1cWvOznV6oNU80hZYI4K0ija5T40Qchvj
SH/MlZqCzXsZhQXdGqahOKVXwDF+12PAIp/Fsf4B/ZOLXSQfflLGVuVIitUk5jV6u5Z8tzs4VCIA
Af/CR+FXka+KASS17WwWGDztkyunzPbFKKbsaw8s+2pB2M2WmqVdggfY34diBbZqaHT5ug7DqfF6
KfMgKMHJ1flHvEpXwiOT29T6VwtzFBMiaAtTYZ7DejHDdr2mMU2qnR77NqCc5N0FVZLyZmQrAbm/
Kkbeflvxebrwl71/Tac56UPvUr118Zf6qGY2ghHh6Os1yIm7yjV/Hb3spvwc8NSYaoGWY+LkUHwq
g2Srm/ujBu/EhJWa927PxCjFeFN+SYmxoZ1ZDNapqHc/vbECchoC/YXUlFpESWLPFylPYQmfregV
H5G7KgzykTuHZVey01deA0P5HXUmAe5x6o9D95jLlSNaSEVsX3yFrfWgkgFjiH4w9O57rh2pS6+P
EzmX39cVaAhJMd0EzvP9kT8evTTuZG1vIeIZiC8fEbo9nOIrEoRuqKeQMb4K08qTGuBux61nXPKW
ckxwthq6A/75ctbe5J3cGOhrtHT/wiQpcfcW9bmwJcNGdmQ6SJa+S4aAWguKpw16GzG0R+vbevHh
1zrp4AbzbMboso6T/s0AQF0hQqgn8+MLvoFZRI5ZG4Dwrr6rkVP0iSxt7K1+JsCCppJ9Gft9aT2F
yoPWyf0TFRn7gZF5DhUsj30HC2BiaDv7d1zm83fbuPx7+uhje56yXTAgmLXU/t1giWM1YYROdqVb
0EGITWv0s0TzrUJ7CLCoxYLYhFjW+uNXhxxswFcJfzCpKXt6kF3nOLEr3/4RaYzb+krIii7fAy8h
UqRtMWa5ALY00wDq6+k1fTcijkTzdjTTdr4BaCvkWB91l4FXSIk3JJirDz13ytDy6qoexLwo9CaK
/j9kuQyWyvbOakOlQqjLpbMEmRU+Oy5pXKILPHebG7Hri580rHdVspDAajZRr6NsHpU4JCNNjnTT
89lu8eiuOz2/yrw7IBFg/JEONH8e68Dd0oJhBufemJUAMe1sx1Ugw2Zx4WTcYBq3DeGLPF74gARh
ks6iNtO5lGKz2gQ/sYSWbJZpCy+nKkbar3ehjCYo5s0h7fd2Q/E5neizapYY2b1/zh44sUhKeQsc
6chokxIgvQh+AQq/jzP/nzosDmZwZDw5Nwbo1JIyTkCIxEhcrAI9sHRtCtNB3mJxGo9OC7V1uplg
v62FNlCrlZhgHsOybcD7Xmn02XyIQIaNWJe33/XBfLYtOBNwctKaY4ZnB+NmC/E2+jmLPM3woo4U
i8Z/Ruy/pTv7BjEyuETTplLlfDQ50XK5OeYh+X8PtJADN0X1BXoHf/nd0eXqTmrYaU9LQcJ4plQh
z/ah+CR8zH8NrhTJhkEm8NQynn3ChNn289BHQuIwNFNmnzyZU/TKG/MwU7DxBP/JFWZJwUzDq62J
iSKJfOyOetRQkD5My44NZAwugtcYXCNQAERM4Uzhcvlv1eRwLlNk2lP7osaJ6dBZ79Gp5kHEknQ3
UmkBA6J6aLzLYB+/BxaQduu8j8ua2DiEiA3A7yc8xFcv74LBe6NWeDUCLiXz3p9qFkMwcluj+uTf
ufEnTgnoE6pqu0xOL1NjW4uTHnMcZUcA7gEZwszPcC/rDvXq3Duyoc8PqNu+YD73p7/nmC8xOqmG
xRbJzX0pVGgaxKAk9GNxi9Gh8Zpdf1HK5pNdQ3zn+4bVSnodfc/4y86dVDpuH8buCBfjb7MaynUz
tZDzx7YZZg01N66EYlFgj+Unb4FUvsk+aLKQYolLH0BFxHTVlaRmwthHzxvWtQnzhQno5hN5GSQo
7oiAuDAY0XBFqNtaEcH4Fhhgym6CSHwrAfvc0GK2GD3KjG5VtKZXFRrJDW9+kpN5S0/vOw/KM+0A
xzM98zjNVq3pIrYEEacyIv44/8eRM1NQc00wPZTsUR4jkzQfnj0o1K7XWfzXNzj38dgZqYvZYMrJ
CxcuUnrL2gE7hFBwWDgRycI0oFyPC7oCEXUEKrfLs206JEedRLO2EeD27q1Um61sbEx8Cb1TJJNx
qcL5SMiUIK7MIVv3jAVQPDxZ/NNyEpL3gm1eY89WL43HU9zLZhxueewos0e23bFd+0g8Gey3fPc2
nO6K7h8r7VWUM6RCQ06AjJ1R9wn6qV+hrkiVDSFg67pFdt36PtE+Qe54xhIGds+mS5cg/Ny9PWT4
JbS0Z+DyKrhMYnoN0YIhC3BMwJkjNeUR34tDQa6ijdK0pOuXwwo5DbmbbW42m5dT46he4rk0IKyo
3gJTeP+YGY1BT7N/GiXYV/zZpwKr6fQqcHEkrGBVTiraJj47cuYiQ8fbLtwSMp2V+LqLt8pQ7ukt
2ZJE2uDC7A7X+Xu7OL8f0FL1yUf1Dzw+RMTJJPHihtQv6s0/BIXRnhqugP2ZTVdSZ0ZNhcHNArEv
C7iMpfC7ERar7HSgMUE4f81IUeZ3Po7BHcEaGwvW7TKWxnxW6O/7DrSUc7wsONkVjjpvaLY5VLHn
9LEoN8dvKbjMtsttN2pV9iB8+1UNkbOFbKXm3vecq9a8WiIjh13cBoOvGxYtugQWsfBFTxoWPzUP
KP2UJCfTD7huKKy4Fx1iAuElqYFrNawJ1wYv5vnik4bcNkBMlAbqIN9WRcytW5lglN70JTULI8AD
h43gmu/PLN7ZpyTvDJSAZrZdDT3wqVKT7rzqfnbzxPB/4KzkpKnsKD6N8CLG14YZXyXQdg9/d6nH
+vM+h51nPwjzOZcQ9K0iNrTatvnieNBIFmF/QPt7GvlmSkhyj+XJ1aBfYULKLbNMcHRLOabLpY6g
6Selj8FAdT2GJPdwo6Uu6Pe6PpRl/eTtab/TdS80txBX/QhS3/jQaylpH6wiEA/PTU1MjYlCnW1p
2YeCAOW8xC7LHgUciIQgz3WiF0Es5aViA4sc7eryb2xfbAlty2sECEvuvJXCmyOguvQFi/VqH94l
1IGdvdPVXkvzBoWF7d4llXmkXK9O8y/Ffhe+EggRYldUfzXUs6bmBAEJAQe0BPJpcjyXsouo0SRJ
O+dO2nBCKU5ifMiiXchUpWK9Xpo0NaBxCrkGcxyib9RO2jk5U/gy4a671V6sBRtEww305mJp6BEo
UrMxdpITSPtvx49zj3ATVX/Oyvb2EHKkaHqlqBYo4ewCbmxfD4IcTlD6V4a4UW3JGq7kv5v7KawG
sBk7xx1GLES/4+PqAmc2VC+drN4r5HQrt4lE81m+z4ZUjpR4OnWL923iIWZjGFehbUejfXg19XuW
apU9x5MR5hhTM/v5qJcZ+ums9RaTJNzRyCCTC7xPIMeU3jLypgArepNkntFAK6InYbpZBUmZpmPr
Gn/qmDZmgd34tL8qSKhw2xAjHmOafO1dQWRtkLk0CQFelTIQ/YeBnOxhBlkEKwdyQ72az5UJA9vq
jgtnygu7PqKLgPOACtdBVUbFpR5H08OHc2WKK78YuTcOMTwLtz01yErBQiF7WgANEmH3qaytA3YN
C2OC2GygyKHUcIfCA4o4vOK69M288uAK5xwZE8woqBv02DeEuBZhAxY9Fhw6+TsT6WLfjJEAhSaA
sb7S5JQ7YmYZyPX0nAlwMJLAL+Da3ptABDIRIL0FK6MhIS4VFzXbAy9rn65y5DMsvLhSjwTCDTQ/
NPTmwvoSwH1Jxn8V5yWwms3h4Zh+LBExDgSLva0OlPJaul/k+4xMlHSriaa2rUCDjQRCeUb3Q6Hw
r4PEUrK3Z+2tysoFOEWVp96s4xxRu9uVtgqThvK0N0GiBOCqBM1w7AAqLVYEwrnFmZJVkwRW5IPX
AMorAajhfWtk5u4vl19QuOkRGKtL6+RW6rL/fColqIzua9PA1W1D9pbI/QYWtfkwnMtoh+c4XGoM
QKfhRXV0cdCYBg2vuAw8NZYjZXfG2HBBaSaEhCfdB+zBy4vJNf7t2L5hpdnSDyU1Oh1Ui0UbhIf2
d+0IFG18Tj4yJTckjWl6ayupJfVrOkLfVzLkB5ikEsb/aIF0to4wIg+D2u7akNF/b5B+uba+Nl3v
yvDswN15LhWzKc2tQ9/2HpoP92DdVQlhwnmD5b02PYH7iRkBKL52EpuSoyAzaVotjBQ8sF3WWQWN
5xBHJCL5o6/NBVJHyHBqlH1A7DR/SNCDZUuPa+jhkKUfGUtlSZIsy4+vWJ5TOruLv8iE+Da+qcqS
LFuJXi05EOzGIKUS7ZeLiDOquLD/V717i8gznIV6cK9TurqoHhqmRO1OzfbmKEGENv0ap4P6RACH
5GjwpOhlM2fcdFjQkNwaBXOtOISr6zHWpZbQmAv1EB2zhjU9QKHIB8IR4aNOLQVIY4ZhA27Y/XzD
9/vaBXYtRRT2ab+2k+QpmAjy6TTur3msohAK3aTNxUwbBGXx4Y+ikMyGClHbEEoPNFpXPM8BEvHo
fQb42inaGzi1w+YXdDAlkZf5AIMfkwTRIQRV6ktCG0t1apsskiKDrMgpoPG3xSFrzQIJONJix2CJ
4Ye4gWzmrhahvW1+o9C+ZoRzv1N95IJFR4UTBHCC8Rc1F+RixzIUmPxu4x5wurbGkfyFzwys7vsU
S43nAS0EzwnoNrB76oEvONNfpJYYKHUaa4IZ9t08OOAXFULcHa9WJ6qHBK94W3baPeLVt3zMhfWA
HRQ5ov89b9l/KWHPnVD3pf3kE2QwILqVnk1CQx38yMkbXMuG66ZQrowmNJj3T0i/eArCXXmZPqLS
6MObByFqXCZpZ6gtYHVjp2AuMDtcpS7WAp9SaZ8OB43ZLjWuMJnYTSWWOPKR78DFbkERzxV0HKBp
z2/ld9u/0LVFZKh713enSMzNCS3LW6rQtqDp+AVnU6hBqFbZIIZC3Vb2F5HAmLvfb0Nim+kWi/ln
3SOFUiFAHOs0n5z5QmZhEFea+O3//2l4CCUIpBoFAUks9XustJ+yyxU0AQbP725CL8+8U4/K57zK
ElMbshW+vMVTBoimjlQr/TucTacgULVS2ORz9lUyG8sXnxpSUrnXCGBvuzx5mFSlOPdP/ybZ0Rys
jZrp1+FB/PgmRW7J+1D4/il2KyINYTWxmhWlC8kl5dhAdZu8dx5DNYnIOyLWgv50K8iq5xES7DAw
WgF7iQhfCMaZ3znngkYXcaIwSrTWtq0kMqS9r4yRZ89JGpExGsP7b4ARr2LBTcyJTlkxkSLxZ3SU
kkZ9DP7JgsH23NULOp3ybtBsKhWWdiYDeHnt3iqM29PIyQlpYgMTqHtITZ+MgWaMhOwsQWowilS1
SBq6As7oRhDNVhhX+GQVjpO1LZHBdTT+Bc98BEAUJGPAauAGF1zr6Hmuz2f55yWt0q/Ovj3coive
Ask3QoEFe4EVRhipLrBJBVb18W9+8gEUkmcDQh/4ILe/qyeOM8Jem1MmyoNgtre/HFfh1q5UiLba
BjGFk7Vhoraq78l7mOulx7g7EzyDmAW3z5EN0WU671ydrapozC5EcUwbppSLI/0WRet/wXL4xrJ0
uYZg+wTDCG00ENJ5ShO3p61+9Yd68PPp9hyrlc47HJ/SMFu5SD8dIWWfR5dACIslKldD1gYV0i0Y
6Y9IKvlrYZcaIHXb+LfBTgKH9o5Cd6ZVeIVwdMX8s7Y/6QR65RfAOKpwmBBf1qdJB/064j2erNok
bCPWz/ZEq0zYPmm4MRnwgvQpFCVf36vnU+BJRo63yzOcZ/qmVI7KcoFA0KO5p0bD9iNbNHQ3qsai
4UfCk3Mzg2iBDtVhJ/RBA3EXk+40bTiaAcBh/Uw3cTGPPkSI+572Zj1f/khAO/BwnXF9x9wE+WK3
jx81b7baWofiQBu7D1zsMjGmLoqOIkZ8RKRaky2n7wODBgung2RRS5R1GqAkwengn9ZhlOIbc/n/
hpQN0YSdiDXnmxw90ARJB6Jl5qF9lcgT8nyQI2dg4t+0as5k36k/+c4F7YPzU8/vgDiiOWewjtbO
2HD3ePpkL5x+eoDSCSkqkEBaMQ/wO+R8I2tTMflh5sE61JjLeOGD0OYi6Wi/OnQT2zkF9aWbvVlm
Sx5ssaFHgsDOR3vhXzZ7wgJYJJ+lGaSB4ZL5y7mousIvET2r0jpVXZy9GdgfBByCEiXMxHLZP96E
KZb5uMi035fET+Hizq2X5ZA8oMWb1jA6Ga4M38NzFOqzBOsx326SvI4wrVuh9pOOig2cqx3erdh2
ONdnuWJBBDokIw6r0VTogPLomj6r0QG4al7CBQu5j0V4jQlDU2RV+VnXOwXc4l44LuHQX1h41nY+
/1WjNZANm/kVIaUWe9o9yLY+q6mTqVOB/5lNdUzNLCrT3RYbyWqwWMu94BJZzZQeJk+1gFhHu9X3
jj3Z4SYVh/JeVbE5ewVFwuWe3ch/Ej4Lo4xiJCGS7Pz091BsP7mNyFkR8KLHSnt87TzYPg4NV08s
ODGsitY83s78hBMjpz2M04hYjQuxw1fGBOQVnpekdOtNBq/1p4mpI2rX96g/GfKprfNoGjIiqNvo
t7ZFEK1g7guecTG4javnl1Hg2KJuIIlDBoxqKKD6GgdGpqq6YzCYHrsMXyAseF4wRvwFTusnU9bo
xsYxKOX060zuT2rlPcenEj8rnj5JVF6sjvHkpXukBq2BMn1ZKTFuy3PHDW/DbX8nx+JjmzRMEwEC
4EVzCliJqy8fxMvF3LlX5tQNzZ0LKdHpOHVEKStISEeQ7YUkpXR6ZKcZwKNIfYEfoCgngsRYWast
CZ0mEzluXvn8ghYgM4b9WnShkRPKlmMVJ6msZZmOhGZ8l6RG07azz9qYMe+9icA1LNHbfM4hriLA
/IEOAus0fgDAZl5U6/34Nx2jL5ICSdsXAtkLyHNjdgmk9M8d//rAiAdIooDE9kYar5zgeMaNYmME
l8WvGycjGNXc2fs/ox0cZmBluPd7A/OCHdKFRsxpgJDri8IthqiN/60K7NnQ6HgJrqsv74JzJLim
kW1XYB2Ta9CCRBGjvv66C2jsbA3Gt86MSgvxn9iErb+VgzCe2ofbsjRkpt8VjjTyfe3sFp+ny5FR
UUH5bE0oAiJ2mU2wo3nKMiyxZtUnWapVDruV5cUNvdG4TF3Va2VV4Qhyze+eNhatMh9duD4f3dR1
W3oI8VW2yxPkS5oLcdhNa6K6rUhBTFA7qpzdxrj09oSAv52OP7zeSisOpSeRCDnUzaGV007tKOlg
zFASJBanIv0qv1oSif33CJYuOdQLiIcwveT+uu+uss7oUvouuEzfLOfoB6Hy02aTYZ7tCkIDcbjG
EWP51ffnMGkf3Fv/n1OHGDBIvtsWSqVnR5IaTqcQ0ghGrgkg3avj58HfyNrlYX2gURMdLkGEDe7f
X/XPEXoIbYh4mDgdSHwUYx6US0vc7lfElCLrNwEfvVzsX1m6IgTAD8hdiskJm7Nxc3+gXXczdwwC
akDbCzZR/LnOaGtigRl+MoIf6g8xalcu5nVV9Ybuvkwy1etBsJNNPlFY3+bNUUzBaf8NTW+OxygQ
ZrS4gJbQocfLCABYr9AcbBMEqB/hK3azrY0Wo4mKkee+hzefT5l5fAFJlKbsWwzcy1Y9i+VWDENR
R0FRR0jtHFBhz9k/cNxg/ff+pcGpYUG9na7HQCZFzZyv4cDHnV6Q2buwli35QyCxP9aI0OSG+kWA
YX6rL6Xl24TgYW0rzPIFws9oyk3in95xIu8SRtwWzEQrEUGcv3UBBFHXfUCBHZIVhm2JgF0C0Z/1
+zp1fFsw1LeHDiAxMYc+ybchdUd/VX0Hv3FacpNgEBb1DpULWhni8c06wQDvIX3XBNGZMFxcXDkA
hptbxwzMfBtmTaNam24ZdDTLAsaA0VqpZRBS2VM7olQcyZFazNMgph6TdKJBjhpywsN8DmnSY0Sj
F0ofFfk5uFgyQOK3EKdlX/Emj5h3u/syz0s6LkXQTTxrquW7gfI1n88XfAoBtOP8qq3o3PimAsAH
Z8y3yW0HkYFebrgW0j7PmzLE0l13cPF8sI4S5SO2gQXN3lQ0kOU8D6WG74vLoTt11ENcZ/d3RKlT
efOB6PhnxrW6n4lGi0Kc8gRVrKap5mCdwAp0IyqSsHSxHQMadOmswWRJY7OpFtXx+AYdtEWPiev9
Qoo1TPbE7M3sjDUd7QJe2qSdW0u305amsPh0BGI0rzMgM8WK8dupceFSNOXbt0t50xsyLVHf8tYy
fNVrlBx9o1RigdsQ0frJ+WMMP1t6E9XCtf7SnqZayJ01aspn6xKJHDzWEk0geydmhX9aoZjs1Yr9
cQmGkSoW0+eLGbj+iQI1G71+0GBRP55kuuL39zcRaqdizEgu3V4WdArjjRpd1fe4AEmi6Q8MwaIX
nJQ3omFKyJk0S9odIDmZTi9Tjr1PHYgc73CnAF4mDz5Y9Kin/2VWuug3rj5qjjHJba2qnEymclc+
1UgYrCEJ698bWTbtc12RI3ABEE9nOnXooUA3bvuw8CKvlQKbdkkfqA1NMnB5Lw3ZZun1GYV53ff6
a+DFCJb8kGirADYt3DNf1PdueXteJrCLfo0FAbBSGdYOfaw9qKSURBoI6zbucOkA6Ax6t+hhhvqM
4Bn8/gvABFOz2W+gDywO18nLvZm3WyQiv+W7Fq32VTEAKPt1k2gCUPYET/pQxyYa0vqrCMS6bnTv
Jb15fC0wi0aKMGNJMWyqnYmjcMT8JEyenZyTrsOibzVDCAZdus9uCH7R2axmUs9F/BPbanbjvnsb
0Xyt9mpb/QA5GeeUx2Q1xMYBj8XeZyg/P1GTHyCyWge+mxymhbr98xviTVvQz7TkwSZLZ3QgQ3st
i5fOvAQRVW7k0qwaFfSEPQJaEbC1eyoUJUKSYGDlqFzhW1uOBQ5NvvgsnIh+hh8bh5z9HdSOf8+V
/8X/6Kin8sx6gmOUdkkPfiReAHJK5NByeR+u+zt91qHFZvFTaoH9YNiTRPtloCBJWCjHyfEy7pE+
lJKhWpB0VsYaLCrGT7Et6tMMv5Zlh3NjiEcAKEVuNiIKHzryLKfy+yUhmj7Jo8Qx2hRWYQvWl3nQ
MwnkpngbiBV104b+btXk7wdzpKEQICFQ0keLyQJDi65AIzSWP2/KQVX3ADfvWIDD9ug/z9j324sD
Wgrra+TxwqdGijRLKn2wFvz/SH+Fr60s4Uo8sDFY8yN25P21qL90efExYBZjwJ/u401wHempKf/I
1H/7kqguEA+pIz2Ul4sDxH9C824/yBDOUadObRYIYQBhRaDEB2vofcY3K8YCAODTIIKjI8dbL+qS
FmE8EQKruqhgp/kw27KhZ3gDBhZSnctxJPJMe92ACnhlhmW/dBqDKEanj5n8Fn0lF9xkJEMP9Ljb
tCFWyAolKHdZi/LNUQhoNFypUewax9M5grfkksk+f2bINSYuDPFc/f4AbeE9T7p/wbvL2WAcwaOs
MrQWburwx3wSF1aHHUFSb6BqBTrJfRCgq5/j5aEiP3T4RpfJfF1Xr+yJY8bEjO5zcex8Tg2sRxG1
8cYyHqCDYPKIfMHZWRdY83uisyWYXw0CJ3IiwMyIysvGtQHTZAt1vYDGFLq8HXt55Ax4MPCT7GyY
GSe5aB/wjg/Y+P89yPSHrtCvVk8ak+WoOYSUBgz1Wql6Xf5bDivoMfYwLGMMbaHAveofxj6YjhDV
vLci4oHCcMhhjdeAD38f0hLoQ+jgYtwbWruPKifT0l2Gj11dzYopUHbDDmsnEUDk3nXuBGKLRAS6
jUUnUxAgSh27dKwiWvsTVHp4S8TY5S75TWTntBUaw4c29F/BrSlOJ38cF+9zDKpSN1s1/K9FXBYu
knADUiY/Gk8d/0bi+WOFZ6Uwuoq5HXhjYjXSl8H9ym/KEVfPJpI+rKR4naOoaTTUPmIXG3/0E4Hd
TEeNi3xwvOBn7SDUy55jVrGaYyql/+L/6l5kmQwqKpv+NVVa4hkU4vCzW6aQ2QjJ3c7Hl1tCDfac
nC0u8KXuzAQL0nm6u4z2Go2Di6npqnC2H+JM8JHzdwYF8N8dHU6Yz6xNCzV24U8wWUP/KWJmQO8P
FS7JNMsTnfeOQBiuH5Sp+TICSJrj4SL6epNkW0NPojiGn4/tWgJU3qZgHtmB57at58bQ6irnNPaU
UrBQS0KZ8G+uQ5Hplk0kMF4HBuIHCJtU1h6joFWk/GXBxYOq1HbAUdvoeKjXsHQcRbkZ3Tc3oJ1q
z5bLbKekQPWKgudXU1gSckHVHIvdmRmWYQz0oXwMrWTYucdhrfMY0YRXuvIr8LRWYYmVRU7rLC1N
W+t6tNqb4zzB1jLUg9SP154Tm1wvINiwxDr8dfiDU9PCrGn57uy7p4W3zQKbsqfjKrwX0ldUmjNY
lMfYr3ie7DWtGVGMY26o08KI/K+Pn5mlpXs9aRZh2BwSNQbovpxlebXilEh/lNdM+fQNZkDXzFZ8
wqNBQOV0j3aUFYDuwn/fKJUFpdmTwvl3LkqxQqY634CntZxAU0j0ti3HR4T+8KpByXmbGzK3yTmK
qpe8Arbx9ykox0cKLwfBZ5gog7nZ1q8oUaPn1KKd1wFLOczO5DsuciSf8ZAYhu63iovykPbjoHQy
NzC/BFIj0rpJuaQz8EyLb2JvIqUWuoqaYsovnP+PISW9w5SAmjfxbDkDfMc77IK03tSiBOgP1MD3
j1GpJ8DdzfF4trx/ibRAF1S0K/NF3iV7g+n6qSnkbV4q++XSXqtJH5FJZ3Keft/MvSG06zcpX5+m
2elICtMwL2mpqPcjEFEItEWjzmZlH9otqXCkZ2frgIIiAIid0JlhXKsEA8Wyk+sWF/qVbVPvunqa
2pQgbR3cYRefQcSHP84XQVVkIWXWSVZtpwCceOoQrJSHzmjGxzAOeYed+fINJiP7dbSAAHynpXkd
UP0E/dKDV53IooP34oFWjLpzpjkAgYXwbN0C/lZ2SipxQdWneXw79+604dn1DIJPjQogumY4JYx+
aM1V7O+3ckERLHcVh+/FFFwY9kj+rtmqOrdNtDaUDYZHMTknQoAwJkE4vKcvzh1ZO9DGdO+CQTAg
yoVu81gdxL/0MH/jcdiph5JRK3yf6nrDZM0sCWqr7smPTu2Oehi4BqhQL3jY5e+HJObHfTrWW55b
ivq4nX+3Hf+/qrYvXWenBRxBR/2k3g59U2sP3xoJzeg+cJpJZs+QffA13QtGOoyPNtGCntzkmZ5p
p88Em8cn+0B5i9Y9QcYogpQomzP0jyfBymcRkf7T8HLZLAZgGBf/kzAGJHuyQTVl0x77MevZ07gQ
1PMBbpSmGDthNwU1oOQiP0ynOoirDTO3722o8x+3yND1MSDpT5JTbCZrjgZxwABiKw8r5E0i8rKU
RuuVtPsqbVulnWeD/lRdireOMsZB63eqw6Or0/CrbBMbbqNjZOH2TJFSm3boNVDUEZGUc+kpTvEi
7SeM/FMcgFY+ovUNlfX8ebRjS2Olyo7B6P+EBtIGnykl5rMrOKYDT6Qe8QPXu8+cj/9XxRWJqhNl
JCVdstN2ZhJcQn5kNBCrpV2iEBy/YTczgHy2YTOMPim5A67A9CtFK9Vh4M6nSjC9znjyBByI3UXv
eh1o0gMl7lxsJgwEgqlRkei2jiH2rxjSpKCB1T5Yetgx2aqW4B51xVXm9TUnPuzGBa8MHsVBNv8M
2ccwljrF9jHfXn9fFfRduZsOJSdGjWJ3QoKSQ7v8DMdUKxRhHKp5G7GTZsxjhtYCJZfpaf4dhL0b
YOZ7fK6xTVzpx2oFl4GODjUM2TvPaUr/wCryps44FPRI3gzAPmeR1OMK2a/5G6EvpnPOjSHvDc9p
ALqxXfSOi/fXn9sGIhMWAUXYgE/2QvHPeIrBoEG5pwW5/0umzh6cvAYyChxZXMdI+JlgMJI3q9dx
4HtLQ+1Ar9vu01y54LA46lXUIPN6dbtEuRh0BRQ65GhAfkRLXxDp7vj56qbxLz4eXwGD54pwI0hN
2Io+MaWxannhLTb1WTo2R/Jvpf+jNZW4Elv2XwGxklXM2dc+8xV+rjhlPLlJ74O1IkZz+vAmq1eu
sHF6SS0zxH9UZEmx5hUq3bATe3lUW0ReW5KzPLu89IJYZy6mOD7gccCl/i/9uKMmSkCw7srs128r
UL4qG+6M8SR35Ecjo89VRTsZcP1E84DA6LyMzl1LZBOTkeKT+OSRWgNQ6LU4ys6lukoQBeYD9qP+
Fj1J4Ri+GuH2UqWIZy3F43sa4OeiuBCZ02IQz+4cKU8NpHg/6ZpQSuKIgM+aIW/REFo1ZWJjq9QL
Zx3nBe7GD1Vq2kliNl2qe43kVYrQg0PhgmU0G2CUxMZbkv39ffK7V2iFmCzbldbLgAHbcVaPyQAE
iXC2lwDG6Ehtx5OHWg8LRLkgt7ETopFvUlsxaxzTXRHpKRC5fqnZXMd5Udk6UC1Lhyh0bAD+3ehi
3ztfxHmvjiNtV8Pb7G8K9XatdDkd0CK4r5OYbHmvA31tm4HmQhl8Cwr9cq8KYhTIPHMiwmsjnRax
qcyZsEPPVhevzm46KStSw5Uugn9Gn9yVEJeFvK5u2BwpqJZ5KvFDgyrT1Oj1jnIdFoLWtmOXlH1N
sSFhSEUNumHKOILrbvQhTMNvwBIdbxwbRo1sITjT3lV88be8cQshum4POJFiDMezzVIkmMholE41
jsYfX2+8NIDSvZoXZJmK0GiR7xLdAhJfP0gdbjoRPZzZxx2C0sP5RHReiSlSzN3IMJMphZOg7ghm
zidZpK8Lk+cqzAwrKwMhOJDvHuh0O6CqKG2TetrQQWEtMjqi9QPlL0yGD6WWILcBVHGsjqJ1rZr3
DG97+cd1pH4ZhYUtOMYELY8YfwgmblzQ3Y4JBq6Hyhdm5YicbXScTjX5khRm8kr5RwoJZzpAyVZw
rW+wFf2PrrOlAd3YYWnYqo9pwlAfxEjU61/z4zItr/JaYi/VBT11y1VtyVb+9NOuU9WUPo++MXoB
yY9uQEyf6rMZ9hmH+SyFC0XwB+fB5I4nmRNXreFQ/q4CX28y16ZNg5DmqiOEjfa/HZPqBUzeJQSE
Bmw2vJY7aTcRMWD35mwy+k0JuzMTQacFE9bsYCVeuPgfmKfudwq3EkJWODlFPozSDweWZ+jXjE8P
v1sZU88C7DHLwHWnEypf9QpLMt5G0KfxA9JiCg2Jwm0Agh7SpOmir9yA/+jeTyFETfPqklqlyYcS
9Cu3n1xu5oYAZNzrwm79fCCzLy+9efXLQAtsqtbWE0/7qw1gpYMfcCAVlPtzY79rpIHVY4lvXPQ6
TqAG71EPDUrFNexborBnraTl/VCJ+kyQMCzFD/kX3v0Znj77YBz1dd+/JxwYxUE8qtPKrH/m/ACx
LZwf72t8Iwkhu0aP8Diy6WWjXwmbZPk5dtrJECZXzKZdOmhPcfeBMW1EyttQGLv5zARr5Pr5u4/T
DJxli1CUIqa3jyjrgbJzNq7VG6SW47uYgGY6reTIdU7OU9ilLVXhiLSUJz39ANtAxps0C3F8d+/b
06naNQ/WhK6e3+6aMffHnXNJlAEIlOH9SR5sNU6bwaF78RMHmSmWmZJdNDUbqmB9dc1GqkEgvgOQ
4IoUvA+Tn8oZCYl7SL7IR8Xvi+izh4HOKLCLXOYdbp119RzMi/udAkdxR2eR8qOy9+6NqgVltDPC
NoOXKKIkYxaztPY93/e4OUWpeLa5S8I9gN4/AcA2jf07yMYn/u+qZRgLMruQHwUVuPvwiC37bL0J
3CbDzyZcxfieut5Q8QK7/my17LlIoTxxf0s94KoUeKL452lBD2pdUR0U5WIxip2U4ziOUzMVyGHy
g5NFPlQLxS7dUwhvNxVcf8PFD3X9F7eMy1m18ccgr4bXa/bVZhfqAEEcEJge/WtZ9nOl+r0o+gAU
jQosye5C8J8H7JllsuPa84/tgcvuqCGSE1cxqzr0affQ4glyXcdg2Wef2emNFNJeyNsOUueUyOqV
tOEUcY47bcQCK1w2+UJDuwaQqI9GELpe0A3XkbFWMYWSKnziHhq45of0xA+QVNnJUyOestwvWNGB
vO5Lg33L+qllXiCT3J7IdOXHV63D8wV+o8KYWbhgipzXlNGLVobWjFT2Lb6HyToufO7HWCQyIoAB
7BgWdxAPHt7WVJenE2XYryVZKs9p4yzMV0tnOxVNQsoNLfCdAlWpuVv8pYaFPn4k+LrW0wZfVNsA
FsAYDnFbxlj9he4qKl2TiQX9ZgW3IVGGLrpdvyOPBbsMNQGKbTkXvBpUp0I1e32i9fnxudXDLh0O
PkStZZ6QWA2PUAa+dGlVhcLc/uzJKPV+o+25W3+MsfvUHmSkEcc2YgDOK8WpPcTXXTpJM/Bme9He
w8Vx8ilWXhpiglutFeJko5MqNxFulxazbwn8fsfHrR+WaWP+iEeOiZczOoeRSETsXl3PKPe3cyjP
y2IPs4PDnBgEyaWOADa99aLIZIYd3gFMruVyYcVfDvvI9uk8gsbHhF73mpAo5jAJBvOiU4L6z6C+
FhgFlbgiDbCz8S8TsCO0GIQgDeXBtAra6KIT6piiEo4cTe2CWbZkuUJeF9FTfEYEtUYK+h4MD3GI
TAlg3EJ7O40+M4dvU7Ww1gP6JJBbaaKkuXnsThPstyR2aq0B3K6o4a/YStQOkVbLGIuvMKTCcYpK
9ib5KJDjGi9zdZ5B5IcaxYwdTETDoTXras0MQL7wasOdvaabLlNUJhLchY8++I7IZxWly1qwp4Yr
7wt056tQGGXk2q9sD9gl5ZA1aSdW0KxK0yid2bq5niNzlBxw795dNmPi/1n0eBkj8DC70YMRzBYp
gH/f4BEHTS8ACFA0H5QZOOFc8fpoYZdnsrwLXWuzgb5ADEdcycnXDnK2K4h16KpTsUFum6/odYAr
ETtNU0DyidnJeEDgXlB0zZ49SDe64y7ZHmUC1uwiVDpZ+krAi0EP2MGFGgR2JbB+lbbE99+HiKxB
zbsmr5AftRg7ZKsud+banSytNPZ+4DLdxholVtNB2F3KLdQ3xDmYE+fZbFHQThjdlWkL4jlOc7sC
a+q5znp3ZIkuEdVSvb/YxOhqN/Y4KcT+fWRABVdY6gAg+6icIC44mv+hNczj0VWyeAqfew+2tz7S
H3gDx3z9MXbZvzB50noRctMkbKyKrwFs4f7Ec18FrSy7jRNlmU9F8rlueDTu4skm3idZ6YqRXAvr
UY0EuwgPNLSvOfneXB0sOeapu7YTdP4Q48aS5IZqZVaj/WrSWCR7d654Yn5GxnZxuhsKHuhbjqmE
Jp9IC61h0Sd7xuLkMJWFfJ2W2KrGeSeDI+nX3U61QcwWLzEqaV1x4xnrwY9UGBBXEzKTd0KY4BDD
JVkQr4Hp78Vy6AnsAdMG9131bDawCMTZIO6smEdFO8XsftvbicMCXJD6A4+UTquAZbXBxCXR1zcT
UWglZCxdV4OuhDoqaFyqoH4UX5GYeHdIoa3DSPdoTDheF25yERhZNFiX5c0q7vJ0tkPIS5/0sJNJ
pUKt5UzapLrBMWnSSpx4qfEoFuKeD3FXutpH3EDV5M85v4LuIEl2HVZJOZSmgVRJwU811fmFzouX
givfLS411HnsuOu+kYuu+f490UN2n16CsGAxZ1m1KG/SwTUsZo/V1Ih+OUwJtg1iuT01oTGpjSv/
PV+O1hcbK8rmoZye5Xlzje11Z+LUghImlFXo51nFFTys0xTe4xv6L9POzfpOxNH500rvoWxRDitN
d/GUxvw56j8FuhV4MQILoicH0SU/rmb4+smhhHX91wJq/8ZijJQbxzhX3cbpz5dA4zgFJDTtg7Ac
JtOqXnz6e53WCrSdoSIJjEZPmLuVq0S0SiWZSW8HaEJEjgSKXKKEzmir4uIlrSIyP3WD82KX+gKv
bAM/QV8Z8k3pgChwQLSm2CK0kp4mYRcVgd2vZcHV6J6A/G5fjJ6g9xn8ixT/MmBz12iFLCydYfdL
TJynejNc5DICJu87b/fDYsuERb4SU/VETDnM87se8S6jDJb7U/irj9fki6ZRZWZnov4h40e6v9Ml
mACFJW+KfBGb0syi75XPsaKc4iYceZykKGj1Gmh6HJsMBt/x8y/r5M5AV5SetGAsKAkstjob9plu
hXm9y+3BtKzU7jbuIreHhh9/4WZM1DIXQk/uh9q+GaTkJ1Do1HBmW811a/+kO9SJ9mNjncuiwHVq
gMh1Gf8v6D5bK6Q+wifDZaOaKjW8U+35rk1CelTyLE2EaBsev176xUgHsEfdfCKb6A/E9NCaqBjh
FTEbj3S60Rkdc5ANlqzTgQlxd3MWNl4FxAFHCTVkFdBWo/CtEmjow6yzleHSXjPkZdkJGrjlfuCR
MU427FOAPjAzoerqciDvKxvNDAkOZutrjzvsbo+xqZmqIw26svOYLDj0fp8pvYfvkzs2TrAmyK9g
3i8cFImV33QU4fHsLwyTyPbn7DegrCiCbuKHP8quF1Z9ucPpFbXA6GdFAdRcC2fRkTgLN2bkpKk3
6JVABBD3YWiMOBAtGQ3mbvZYpRalU9s5GVqnRKm7YFQfLBCZZWa9XvozWixKOOXHXVHFiMp2mXXy
FMtuM4krYUI16YFRgvroco0cKROb5fzvVB9Bt6OZcxwxNxC1SXBFcXdNER0TWYO+us+PK7fLjHwL
qeCGk/UIZdObD0Bowgf4axFrvNV+Zju0Meo79HjnLLR6e+/Xp6YybO9+n+Bcp4xHqshzc38ZgPXj
5MfXd+VyhcyKCKRaWSR9X0RuqxEoX+SQPSa3cy6cRgcmc7k/hZgbqaxPOJyNT9fVY1rFKkKPT+ge
+/1ka3SiM4TArjj0VHjnWm4opepkhTOMped+AYnqW3JkwRTSIabcuEEin3DGioFzU5m1G5aAjG+Q
fz7N4f0Rb7TnPfX837aJ4V/KM5qo6fccr+Bb78CS7spWBCNpPpSVlyUrzrjrcZXnqbVxKq6hIKM8
mUg63dwWjoBiQ9rHLdkhL3cZq0efyJ13YmKeWtU3lO7HxCLZyuwK747JRvVB9PSD9/VlsmzE4Hoz
L2yU492EU48pXF20zlkmRT/n8PPUDDueW0QfsWkhurYsnl4GpMjC2957LdzccFXqvUAE1eBsJ352
qJslGWcrEhTUsfiU7zgN+V28pzQziBuKPs5Sjxm8mFD2g9iZiqJXF86TNlqLdmg0tWglwXqKbxtR
i00uS2BT4rZkKQmd9/2xB5qCYWKtT58rS59+P/tHDnpMlFnYSsyYNPim7PC2nqgHTDwoFEcn6/4p
bhmsxVOygithrUq3Obk33bSyKuXOKmfCPs03b9RQ2TXI1X+d7x4XjmHyybomrb0ac2wuWcy7oEsQ
fs1VqF0VwEYxYesA4lTtBFnyQckt7KJnZjJ1lJjn/adtNi4WLKwnD2hEZPUuos7kEcZLBXGlXot6
g7MjmAZrafAt91/tOCMUJqUV6epFHuLfjCZMk/tHfye1g8TR9Tz5HpfMWeCgUu+zYCQlZaiexA92
FuA+2+s1VhoOPHehBGVQKOUGu9SqktLJGi17a+K2550/Yfs2p84Zk+sJHrx/WBpa8AfKpt/bZe1x
szgl3RmUeAWZB561RmDnMkMW/Y2xeb+1/QH9d531+py3IEojZrsrsnOkMJaQQMMi7H2+B3+v9fWO
Gore6jZwYxnMFrUqhIM8LQYAAKqETJVXuOWo1cBJoIHN1qVO2flfpMmh8R9dYCSGFmzQNyLPXv2N
8c675aMlDDWSL5eVVFK0VeJpHYNgm3OqFioNS6NSRRSXpxz5KZvsIRM62WM9DkwqDRaJxyzvmr/N
VAyUcN3FzbsFUfNwFv3GVIXDo4Q/MpEdh6js3VJ88n3HN0tqAa234NPJld5zCwQ6XzKK5pr6vB3w
mssCtc8rmVVP1Z9GNqn5+rwr1916yL/2gAviYxt4HWcq1ihlMB321qpqXwS4rr6FWw1VzWYpUKN6
WD0cF0kLSteiPMEVvWIRjoWBNziL0/MJSKCD0knea+6gY9MHSxIkZ75imS+SIU2Fs9HqKpkyfatW
x4QL2ENcb560YV6v9yuTGHeOww5CIv9xrNl8LDijUe+9fQfhbQhCrZ/chYma0FXu3V6Nt6RpQix9
Ge7sMvTw7d7URWRg1TFU39cphJNW454RvyYCCjHRpv7i61e2yiej8XFrG3p49dtWnuNCG3nKkGOh
VXm7Uad/Z8txV9295T2gxzUrFlYIYuB8Xh8Tvd5sM15e5sRVuzmPnH3rYP0wZtxSRjulwZYYGJYa
8uIZtj5Ah1JrJNdKa24BMcp8KyAAMysmyYh/cmVVmzrRI/7Q3MNx46OmHYM23KiWtOdJ13FILnSS
0j4umpufvG+ufuwDIm8ejv5Z21M0rqFqrHZSzqUxSOaVplX5EHWRznDxdAezYzFQIVaSSsmHb26w
tOgISPYrp2omLEH+K8H16QmzlvTxn1JO5HJYLnqlox//YxjMCZhs5+XDxfIdJHTE1v1iRhyx0S7t
4bL1r8iMFttZlX9p0yN/3rzX9Ch1sVhkvnFc+OK01LmMuT1C1OXnZiOhip+8fVaMz5WHSO0em7og
xJHCL9G81F7WLXTSNXdfx59Q6pdm9f3qMnmdCqbJG39q9XvfbfhqolC3dUI5NwsITT+L09QNAutW
7RpKuEOhWDv2Ol87R4Add2IixYQM5m6S/VMwKUtWvydwqnPKUmYGXprF7h3ejN5fiwJreMsW00ly
Zi7khVsUMASBjnwAUp5ySQmTeYbW0CjR21etA85Ou13y3PGy92njjO3k4/yMdWmGCTBHLN1nthqn
+tVFffAuUyrnOfc9dNkvS2cis/CQBoi8JtP27UA2KNYTvbK1aeh/Giw9hX8loBsfnT8r75eD2YvC
NlWt8Qb8hJrbIeUmmtBvJfJfa1B1neHjD/TMy0cupPsguiQMKbaOQdYjLjX3/ZBn/xW6X0p/gK0/
qYtFT3tsIPFc8RXXN1E0ruCbOrRSTTp8f+e/px3yY03T/SmxvnSwVP44dg9vtDL//bXHW0UWwRHu
HgWlDCUu4gCRSyJsXu0fjiYnuYDHE2+l+hWRDBHCnmlVKE2VXjt9qgYN6wM8zNF4o2BptYpgsUWG
Rcsome5unvqdB8VoEO43FQzrPSK4ZpYmTyaDkKIxjshOzow2YW8GYc2ryrD70QRVvSQsms2k7JA6
0y61SgEx92N/rbMiWLTfRb8JMLCbSVARyCxyRnypGUqpL7vYmllo64vV0XDEAxxY1IO3B8o8nfXv
5L0bZLR5UIa7mWID+wN6XaoJVO10oVJHQR4orpnLJAu77IFeN36+mIBGHcxpRXo2oZvIqE7E36Tz
SIzJXUB8fDFG6NzasmaocfW6oPfLOLKlOzViMnyBfBZpZDNtmXyLP7KDNdYnvlrG2P2BsXA4y+UX
UYmWv+LZZugSkksTkUij3WGoyr4so9zYzo2c8jEkjIP3JXD63KfjglWkw38eRZYRtlKnpz65N7fO
JjT0XK6e3av2gtVto9KRJi2V2Zjit5rgJhApejcbIhAj0Egbmt3utrQ8B9mJifTwf77L39hOX5Jm
hshXjvoWNtrdRt8M6gp7CWNycorsSkc5dD1uzAdvO+F7Ui0mL5aq5ELq3DZo5SoXwbWPiq3FLeVa
jqJIKhzKk0+4pNyBW/kBz15UNjBauHaDexvt5E8CapoDubE0AMXyRePsds3nFREziPpYF63TQ8Vt
DV+d9Y0LImlg6hMIysyuAoBGy/RzN9UhkYu2dmibY0bOkigvPjZsMkxMi9jEPkc0con2H+sQIG3G
3MTfPYinDuVQEFTxu2abttLvq6kVitrN6tnVlZj/9vSwUDoRAfNPBAodvHrWIwcde5mjNapQ2tmW
UD+duMDBrUM7Tz25JPJgaM3zbHQLyKBcCEiNZ6D5KCR32nVHlHkOEEm3014A2OkbUdip2GQd5rUY
KG57dZwVJ+KeZ//W/uW491VhyYYDoCy1xQbPwnishjB1L/xg+IJG7W5CXOhHoGqDtBvo1ZFVhMvq
ugWMsEklKh0qwncohK9FlfQ+gp6otG+UZRYooPNtZg//UbxYB75AkC9DDMVcomhDDmER2ax1iV+V
SRlrGdjO328olE8Ljzfzy8BHoAdX3dIf1lE0AfXBbofzaqXF4A2tyLK8tJHUh4nqkDWTB1rLjS6L
6J772Qn23Sa7cgt6/SmSr6J12SMB379rYFuZuF/66OC5Lcx5PrviFgdj/uxDuV7hDX9YybAmsdKl
OXjEfwWdbiQhFjw050BxakfIAm3c2PhUkqWbaSU+fYSQ3yj1PLXjibHOyRY6piCRhch5jBycD0ml
61KpKfsqjynPMBsNTJ5uLFcOINuVIeyoxNqrOYN8LOgZyRZ9lXXy21qh/xJPEDFH7Byc82YyTN5W
9b1MOtzApvXL4P6MkgN76zZXd1y7UZcUeUnH1N70ixMyjsxQn1MV1YViX8maiKC7xHfExdhCoHt0
Vy3LTp1/2ql/hEEijfeslK65Y/vIK5oCifk1wSv9ZhknET251JHsfK1Xyn+1S/Y4adbpmTq2B//V
Apa+f1WUfCd0zqb6uPIGmlB3xDi4meOVG3l/VCzH0lkIrrjjQrrA8LE16OTX2kQO6oikGDVfZSsA
4kyldzbCmkBBEoTOBXmeZVBF2YGYrqad8ew/0PR4278Azrq3HBYLuMHUg3J6rjZ6xF0BLeKukPNh
7zjm05j/BWH8F/tLnBDUEn8snAeel14T3JCq26DdabUpWBsJdk8cXPrOkxpuE8isnIYKZt/xeyxA
Y1VNQCS6xPMMAcZPbI4raj6j6vb7G/4gFiSNBuxb2lHd0sxdTN3sLXuUbPclGqn4A4/gUfO2EhBp
HnTsWkl159jop7Ld3aMQs0I/B9L0b6LTNv7RlsPAz7vjSWw1/lyz9Hzge94P+/PLigsniz/TPSUQ
WxBb8V+Q5EoEm/b6aumfvf5+u51R2UwjiOAlwlgPmSgRvICGJcP6DxA8h9c3ki/QxRAt6A5gxmDd
CHi/3utCvy1PmxW44OVrANqv8+BKvmv6+tguwmnKbjsarn+7CPhKKMb5luashsgVWGqGdr5m+kci
0DgUEFqIX5EFsdMSVQqzgfjl8mzSDn881vYtT0dcR/CGcv9T2o/uGYOWCRrbhsldnn5edPtC480i
K1CUtMnqpPVn0+8YxSyrSpMOJmyyG4FDZnrt/qeCEuhpbRTLVOJPe81pKXlXPW8I4CBCWIbQXABY
SWVR5nBJOFq7LhO+6+08uCJpx3YrU+oie0LSHkJfycr2Ctni++OVIAWQshdwFFz7Lmodev6OPYBE
RHazSfIW4pq+jSUx+9UVo+gYC4W8azjVClsC2L2X/W6Iaw/md9Hf4BEQhXpdJu4h1je8jQjfg6ri
l98NLQdbFd/CvR8RZRTvre2gX9H6apIyTjglNqTs+LCFasSITBYkR90uIKtAH6AYKHPt3yhdR2ry
dPhsJQVw/VqsmAM09swOjhp7J3Qh9rkvq7DcoNJKMqh/2Pvb9rBThHSnjhI+ExRcXKzb/PlL9Zy4
BbaJZ0pjvl2RNuEE9s9bGn3qPx0UaxCNDLNBxqNMQxrIFXkCxeLCdVcJZ8sA8DXzYJzb3efXSedW
9EIYSBqWS1hnQGY+XfuZX69StgymprcbeV472Vn+xtUMWaaJ2nIIgLAkYZjQiiF5B+YhWQpCBwUk
EBM64qCfpEDd6mPso4fcSycK2UmCCbodkbouLfgEY/GopXQXorxK4tpPZVQUy2bVr27dDr/8+xwi
AzHllIhk57WUMVeYTUlFnQSX+s/1kwmg4dFQdsfpKu1ngP7R15JuJtixGh6zq5hwOQZ33zAIgeY3
vxGslyeUZqteQjUKVvDpi+3C9H0owBkiVqTql1UyPmgjio6yxQgZaVztGP/diQiTpgVe84ef+LO1
ulsCihl/EEaUfOq9/lAUtyAch++8Bqiy8S6fOtvR9rPBc/7eRhF4xWuXIhhmEVqu/eC1YI4vDjqA
EgKk4hZX3cDIeuy8njFTS2kqluE8EH6QBoWRZHWonIT5swpL5Ny5mjI9jiIRTwM/thayzlwRP48G
1Hyj+0xP82kAKtL3pFIOwArO36w3h5eMHCntIyjpHOAssuOMCvZ+kO6YR8uJshJT/3prRSMpW1DP
gybE+eldkBdhi0obHaI5dDW7UB/lzpzWGFFKztTvzIJsIWmIDoKKipeRTGyYc9lgSLpv86GTDTcv
ok96ZFBjRtSwcKEBlD2sglFxnV+JvEv9aXt1+zpYFq8gNsBw5WVvOVMD+3QRFtfJ+cKz9IHgffkE
BThGusAGAS2Ge372AHfUTARdyTAYbXhJgg+SqT2oEOcPx3mryjzLVjm/mhgYncRQGnhSYQJq6u9F
EAKygJcvnjjK7H/eROuJverkCM24v7VKOc2Db5Ef4goRbvLN817h4jK5ZscKi/wXg5D5Ix90qwAk
00kSvkaiU+7eKPj5eVWWm4pIf0bwUyv8z7zZK1wm9EXTiekQCtQoSvCQeSuPbaVQbvnyqwRLbxGM
X7BrjJxXKBHmXtwo6nBiGj4TYUWS87fRXUEcqhT/bk+ymr0pQeJxko2WNjReIFud6lKVeeWsBxVS
rI2V4cIeXrP2Ufc6jp/Knt4/A2Eg/8NmtFLxXKeA5VZWaedcy5AwFqiXaWrYupR0EARYHxw2R3Yx
F43T7kqBrXosFVYaDmW9uAS7KMYJB7/W1E/wRWiionbCQ3kLMvcxgCL8xoJuJChiJw6xgiVWqPCE
Wzy31PApYEBecYhssduX7Udz/BcUbVjPAznLcQypemgt5W5yN161lxrlKuKrDuu6oQF8fiB0dC7t
LwBfvkVzYvnVR4UcPebbzWPHYE6d95pzQyv3nR+VvpLWtPfbhrFtRCr7Fp2hIOi54Glrl1ryR2zk
f8FC/9l2VPe6ZKgTEAl2O+kYuzyIRRnjZDRz/YZMZVa6MOLYAthgYNUmEcjUs5kE50pdfjLVUFHl
ZWWzzpNZREwHenr7dk0ywJhTexyz9YKz9Ee3SSroFfCz7h9QqABfea7hmrKqQPOjNor5Vvlzmf+f
P1vmQMtI0RXuPaHWRzTf4cPghqcFLLHWscqK5P2TGmuw+itGgU05WXhFKSwwSXchRPPKQ8Y89U1W
YiARNgyEMCHpjWjeOJ8+OV3NGPBMC40p37udSbHgluZvMS5YpBFGGahoP1p+7qnwrl0Vuctkexfz
KefGDUFpw0SEuzN6Rvi45MmO5lQgYhWBeuvZg3lFqszB/4CmQr9eAJA0rCBej6ogqoGjoKUFAVxo
kFbuv4EoITobtm1vsVWtSCw4eSSxIzEGB8uaDiT9iobYetCPqidmnUj7IeMuNLc56EpxSM00TNmo
YQV7nDya9YDA4nyVsH/viUagKJ6yUIzYkEvUuaFgJY/LNn/qAI4t2R3XPgH2yMoZbVusJX0dEdAV
gpyQtnpmoUExenSxw3Bx58UdUJqnjMXPhNQXaNk+EJ/WPsdRG5Lfyj0e1WqqP+0QvCWXLJxAELA4
pUxWNZLVgMWNyOYtd05ZETSd7RrX1TYUz83JQuJit6OummxSpT8sPScLcPbREtPsl2D8VV8UKthU
LT1une6u0i0lgh3cXtGzNAFceju/jV1pLoCOvdoaoBljoHxBTtRtmP/KEv8gupn88KVK5lsIaid3
xkG+pNw7VXGD5z5A5O4WF3+mG1l2hj0Ups/Njwf9lrWGH7obzPsJNLwGk5niTi/ZLm2J8G+jhHzT
ewTaYkUvejOSbEXsEfJXPz9bSd/dmH5+oAV/aY9hsSjjsBpMDu0/1jorJIOlTlk8F7bRHstF9Iu3
ttzPDeVil6TbuC7YrMQmUVr7487yNde+c/+O0pGDEHmLWdzC+xYvgGSPLaXWOSSKappUlfNBy1bp
9bHLyBmkchVVRYJrcxzgbUKJyGz+p57R7OHExFvgZ+b1E15LN5sbidKtHoqkuW4nqTiVgs0a4y/u
QU25IHP2G9A9tGIdEPUIZmm0yeR8puJN2U7HsjhopTfyrA5Ogl2ISS3k5lt/jfN7cBndUi61RAKe
uZZTYL2etWMf5taym6R45xz3qAbLUTK1+gKkH/Jly5RPCt2/yCFy54xQ8TaZYjC+EqzT9uWyyFjt
SzBQuMsqufZHC6hlGvGj52ENUHRPUcR2O/o3mTk7Gok7XrTUwCs47I6HZc4/gY3u+Vuv+5+93/AV
9T6zIuQNuAb/qdyU6yimu0lRlmqvdKN+lZEjb8kAc+7xFy6QxddjLboMITLev1y7gaBef0Ky4nGk
gyrjJH+PW1J882tHfWX1fAgfcMxGyD9YExteqaDjcMAtlTnxZSwhWRviETmTyKd8U5BOVs5r+j+g
gKmEk5sToSgK9da82VTG+HeVqdDHNlDqrJhsHKEQQHY3kME19r2dPiOod/S3WZAvdB2jHKVNDQQk
ZSHI+B10j3AY0xP1uYwLlvuNnjWoO2DIbxt9Wc5VmFsJVj1QLvEx1qUtP3avGUxKKzys2aLONG0k
GbtXnbMHGlyIQrDqWAMU/UFrak3VMTG3F6rYt1JvNVTA8jTIEiISbGYFUicGBDLpi5BUeBMVwrQ0
9GrUEXL4UJr6z4c9G+la0aOOylxovO6G3bg/2R8QKFEkT7IqnEBqEmLJEDmKbQ4hFf+8BMpD5+Jb
1UVizmln/P5wczBgkcwDNrSxvXj/RNc8Lqga6ebIBSoBZ9Ab669rD9edFdH7XUDc/VvJEfh744i6
pQiVPX6pdCrV9X7fQncSqZSdrudia+EQBGp8a6VLkw2RDMa9YtpmMgMZHBQ9bwdOYQpNuTw13oOm
CYnO1vYH96C3bZwMxRyijAZACtcqhjecmKwoWcyVKnvAjsKx6BM2yTUaYt7drS9JLSEGS9NI4UyB
/FvfvdzIkMowgwtafAoF8CZ8a4xz4HfiYFHdqG4ZISkJSvcPH2kOd1MPskNSYDdtaSRiC6ILAuq6
pzKXm+JZTvBOW3jGqtySmWCoMj5G/U5tbThkCqYJg/yX0HjM6VZVz4N0xDSUm+jQ6xPu0VMCdAtO
YOkRSGg4HbebutBWZ3Wg1fVLu94xgBfmQzDHdkYnyX8gZo9ZJweNyngKziNMKKJEwg9FjsN0FIep
9Dafw7zJfezhSOlUwhClxWVEBv9ohfTt24R47qYe3xEejeIs+vKdsQIZLQt1gQ6+8Md3VV+6Gsk4
r4fhlMJcEZeo4WOS4KuRvzOhktrq9v+0LSstduBN72DZny2vtk2eULfn9u0CEOB6VIGGtjIOSFyg
9vz8UYyCX3s3PBykEUoHNNbeppJHAqu6okXYOvx9iRpFaloCJhjLkzxrvnAvwnrORnwM3W8FE2uV
FUFZMWpYGSs12UfCamQ6BS4pCW55HgZR5K0KAjppv7xsK+elMRS3S9+r/3Vqjb/aFoIe8zILWjtm
uL8avq4GCdQYgiHh3kMYQsFIZvhOpkNi/yHpK165kdlMA5HzPiP5S7539w7hTuNA9YaXcNRWYZrB
3sqz/wqJ2fCLeL6NXr0HxYeKfVHROTO55Uo8Cg4cq4E6XKMHhZ4MW8Hdh7QjM5hvhgBfRXvYyGrF
HiqtS4/nuNt4h8MffICkgaUxIAiim79uReVMoZExbTOerrqqFqzG87vIFxXiWZAoSJGA4xUPhTO5
0ZGVBxaerwc+rijlbzJGUvQLs17LczuEoRlFi50ITr93GQGdUejze9DaDCYbeMw2Cgwi0Bym2Ey0
o8Lhf0hl/doU1aRFh5ZIcCwtEeIlSWKy6c3KCu6YIeHLCnKukC3K+LBxpaAn/y7CE0ZIrzL6zOGX
MCicjrG6wt0EI5mqKnVuhf84D4xA+He3J11VICn/U/P7wdhZJtmAyj6viVGigPFsu1azVpyk3pUT
dhjFyeVcPW43W2T6qz5lEFVjre8SoHFOEBtE7CBP+LlGnqhy/W+0a2xmdGlEJ2L2yUs94QVpnFVP
h8SdyhGjuctNjjRHZ4EIamwsXbXeN9X633HFOtoe+L4Evk2EGpd3eAWug1ObzhTCA3rjcGiqMeBh
D6cN2N1iqgKV3IZlIye655yS5QB0GyOWVVZbydwOadOSf/c0fMC/Lul3yL33epjFO8GsyKnbpBTG
JvOWmsA3CHlmoTLCXHqS0t6sxszRYCsnm5jNsGppSwPiD84Q9Kn5cKsbML1R+sMT4XJ9+xKvhECc
J7AYAeakB4Oezhlc2bpFzZUuqwMwbLWUyY3E6ddrANJ8pFjzJ3KQ1B9K1bL+4Od194aKj0lqJntr
SX8U/2edruyHfpmLrKf8s7TDTFZwG2l35FzRblVpAurIgnsQQRdVKoBSHhU1BSaYBvQsoBLVXkmA
8TciKqbd0zkvgLi+7Uq46pSBJWYdgTK4a8XBJjPU0xl0pX6rrfi3drUDoEnuXMCLgdbxNYUPcfng
ur/lKu8btjW6DzXcdxO1KmaDX1i6lX1G/CZSmslZ+QiueyxXJzZ6zg0kEJHgNmGAp688Npz6Ad/Z
hshr/xzeZKpdIY9brZd1lcxKdxlfK/3S85vqZFYpDEFY/JEV71PITJGmuGAgqsiyVlRCbohlWhDI
gFaDRwDQ9fFYHUzyJXulpAZgEJLqXTU3YBtfKqINjRsOp19aJ6nH+RWhNfOdKW5tZzzCQ1GQrp9H
bqrBxVhqNUVPqW2j5BGxaKCYcLVenUotf8+wX2VqqfWCtym4JMvka5Fl1XwSLHA0HChyihkUbv9L
xgHMvuDJF1ef10XWY7J9Zycvc1dN6UO4aXAQCbG+66v/BFcysDaJQInXXjVXrW3sEng8HaNwimA4
PWJLFyeq9EIii+5Jf3YFVCulR7aTVJRTSLHI8Osbt51uVo2p7ylfd4Vyds4JH4M+ckT2q+pGHnyG
tmJEHiCELEEIriUbpzkDx5SHse6nqAlHw2xOOfmpwwd1gSwPzj25dHczFzDrSHRrW7YwADnMVJMJ
EAw4Q3W8PWHPnMr9Wo4m/dwEl4/pV9vGpIn80OhLLviuYRIqHDzvhq6VMarHOrgjVEIOBriWdLkl
+812wcKJRha7jIA4zc7KLr8sVFFQ1lwqGq4NiOySjZRhRAw5HoE70SVT3PMOzuFlymqYgXrR0Ibf
eqRJctHuA/geyFf0VXlo7q005AHb8E0schlafecgVo+2bwmZH8jKmXC+7HGNDvQWQPMbkRAx+WA6
iKq5/nOkio7TpRKm65lkujQ8RAwPJGL1VrGVoLY3Gs18+8g9g639nHKubUnNnFBsSuHNEDtpr027
qAfwh917BzWSrmud/OJe9AmXVxTCzDcuj5wVtiPapHq16qWJpn9ad9pnKlKeb0fTmzj4Hz0UxUIu
DzHgfbxYab5SUcakxt1E/TsYtwG1h1o+HquBwxYq18VvHAZwdp7bW+93lrmlHVwO0GF6+YL/+/Ge
tlA1Yymv6Spau1dkSUpo93QbRFAJJ0mlZ3SmhrEo448eF4fC+nv9JU5ZrSiwpyYerID41mf7OoRR
2to8XrSqF8eNkp08/JUdu7RuL6bJH3MKeew+/3u21ZtWibNn6M2bKRCFTKs4AyZvI15XcRM+1I9I
YHIp8k1WUugFjIll+wFbaOCa2gyIm9xixSpqZv+L7S3zDGH5S3RY7qw6hkD93HKmPX+CrIdm6Wmp
U8/TJYA3Vrf0PJRawb16s+IdChedjIESk7DlMwGdEgsXI8e8MsvSBOqWvJlFphMbn5reekRK/K3F
3s8yIjoQMVFl6Sy/YYivRtBPrhwGtwlsjYyWz1Y+QI92dLF4Q4ntWi5A1rpzTcCQrHSIsCwMVcLX
xd1ybJCfX6QYhXeSS3uersa850bYFmRgxMLagC+NJd6Ns18TQauDCbG6+ykvuBz63rlbBwWplx07
qXXIwqTGgoTvge+Z+ocyJ8pUm7NzcaUqehrSTV+afIB2OZFSusc2hxC0XTzgNA7RfGwkCT0Is8bq
94CQXgUYxWCHYWfi+Osdawm9Nk9hejaSUlQBV8+qGRSFCxRm/5P6VUP2jPAbI9DJbeVzBCDvIOo1
uR0RE+dqiBbrOi2s1ULGlmZYj37388RdgaDj8wo0b6kRhnZOia9O1IOVY3k4MezS2VPe6dRFt5Zu
kqlfiIb922TSNh/AWnXX8fYlDH39MZoZy0plwVS25eQ+RMMGCxpJAxrnBh0UKpgoEXTjRYch9Fd5
n/gqPMdwQru5u0uhSES7aD9Oa0Q5elB1zCtw6Urvc8CktYdWO+nyD7wjfLtVRfcqUQxNnGs4TEJk
bgC84rNqPnRLC4+PtY9VSSsCtvmeeKhdttdRqnG8kp2DVqeDouR0sB0VrmyTyY6DO+H8K3pzuXIE
uLocDNGuL5E4t6ejHP49aWR21WFtgeQ0y/XcVRXbuM5MYnqotXwGdbncTE2M4WBAb2XJg1FJYfe5
yLFls64f3BsDlYoRmo6Ml7BfEy95atjpuJFEHCE12mL/5Akr225rNVeqtOnm2lA/qVKo7IGtj9u8
g5/U9tzYvVeT5R8xq8unBrDWSF3Ei1AlAi7U4GAMN5fvOK0I83Zt2wbuYotHDYNQ+zHWaJYMEeht
ipGCLD4DaohCeMeYAg53Sh4M+IX8kUetAVPItAIUDQNYHhy+KXe2uhU6F/OpCvvx+NlXQNobU/xB
bu+RCeGS+n74BzEv+dGQNkTz1cCyDKOFkEFMNO9XhhAOVuj0eaEshk2LHIIrFXiJyqymsFXKHmvN
XJ3rbjl4X8p+/Wbj9qdQ11NBhHrad+/ujBn1R74KnIusVnjb0ZcKrLNVsB56u+FDV2ke1wNA+SiS
X9T/GEWvCbHCE2xlSaIAdiAYQhRR27kokRBXsKut4YAsXP433XfxggVknfL1f6RRvEaKAX/6E7Qy
K8TKXuwTVvq5eUryHEty67N+aCTCxlGv3cAee7hnbmds/s0mhLIJ1AqJLuUYIcpsGzFNqCb8Vywq
O/fTzJ0HlSnjwN7qHC9cxGtGEd6qRTP7NJzPpAWEQ9DAeq1lW5HCrIxp+YTx87wt6Ldw2PPli8za
tUkmlfANFnY62x7sNDXWPhAYqMlSqqDolK0fyrYtGafGCMpKFUqMDjDy1SAGYN1ilOrBP4/lTi18
1dlURTmfoa7kX3+bPakWt5S2WDUzLZH+XG0K7vKwMAM0URV7ICxdy1wioy39s17HodVRIeI6VsZn
KQxkYWlFnOwq0YPup0UHlb0uSEOxF0XC96PW5XHbSLXtRU5mBMh7e5E6B9E8imAEviZrczFZBWK7
bKWtPsDOSGrI30NfKML9wRovMMM2vO2DinxBWhsh6xcSBcRKsE4kUbgP3hloItqRVWwjQOyJHjGn
asutOsSMapqXuGzfOSVFp+JD4Ep8aigRFStMZJdNTl515FS8yAX3Bg9ENfDYwWbWcNnZBO61mSFs
R8EZv+4SsNzhLnfEMI71JJvIhplEb3Kugxpg3Hy6m9ab+PUfwG9GGG27HubCQEpT2taTjQS7JRY0
T3EzVpuHb2IG/0YvW0aVvkgh693LcmLaAgAy4+cPvvECqZPR8QKWHZvXzF+h9T7TTo2vhHK85DUB
u5ObuYIQBPguewub28fBzsqmQrN/vg3BvU8ovyD9oH6HHSWHY1gsowjPz6rEILlW5MH3dzi8/LeZ
pzH/Bv8Sg2gnDqOWbHtP2bI/pUMacqm8DPsYwOLWXdJl8Gf1cOCzFsKMMKnDW0Yio66UGsMbgCfN
QWRS45BcDZ8son1YdV4bc+O3OYLsLxuxqs4WwvaDvPZi0+4Kn4dFAt+b1JJtbWAAZ6DsOjXLOaIP
ofgE5QNt14W6kE/+dgcUXYdkp5Ic5ZYH1fs/Tha5yd6frXhgNOo+u/WXV2ipsjnvICGnedfZDswV
UyHuFLwC6xV7LkDh+UvBnA54noaxAofPmgl9qW6P4BePvajOHJyDDvQxJAqVTpk9Nc5CrEubqF/O
7laf7eDZuJGXygH41Hp2sHvMnCJoyPeed9QaabtHANqM9ZzF6J+nkTJZDVImYTSKHxOaWdh46Gpe
7M0Y43BugWiC7yRESm1F+h9xC1C0646XHnhC3rxKWeg6Lxd557lUNQPCEos80nsFct9ehtXpXIWF
9mNwP6exeyBgvFsspRYGGISVdlC0PWxWUCozQXHNnRS77uvFdtPGSd0dBl0pWBzfWzZTAm8oop7R
b843UF5FI8LeEZgUBFMaUAojvUMklPWCg32ei48xmU8HdMjn07hV0E919MvyOrxENI1PyPhbq4fK
lbs4m777u9wl+Riz4Z+IVptNMHEYhYin5qlQHNO/euAxhGX075X4x04tmA4CoBgJQdHJG7SInvHS
QPlhXuTScIttTHOcgfTrIArvzN4fPk7ck170A0fLBp89ad1p1MqKSHD1VR2wMUw07MY5JuXIbVJ8
URvYkbp2sW0tBm4z74GzjfmP80TQ0hKOsGSBXiS3TaFyULMeq0FGH7Fw7OmFVu4AZ45z9kMkX1dr
13ESVsfRAWC0mEDHMicPXOYP0nWGeQWzMOiVkX9JCSwdQYppxvsra+SRYBC8422gEsV1VD5PPjxO
wowO1oYOYQMq1SBpdYPc1PHJkb7YzEgEa1vSWI2LZI0Na/Z1gdZAcxr2RTcz1TYd+44AYYJ5upk3
jKpHtghXt2PV987JEoHce/OS8PXjnkwxEQHS3+ebGytvcodKDmTAknIYoDdHXZBAqHQVFRU/cWwj
zKBUzbi+ymtt+Cr5Bu+/FvOrdupJbmc7VtvfvijkGgT0sUtiGsF+j9h+YfmTs+iWHnyuDvA1agCq
n8+aB2EvqDH8dXeiES/Z64+H+3m09Boe27WBKngHXHnRldIssaDhj3SAkkmt2jyEA1tjwCYsk7Z6
2uAZOqDesD/4gzh0e1CYb6IDdJOVI5my/Y6UleE0vN5Oydpfkm0e95PFRGmsqCm0c1twLii8odef
MUIxME6AQcE+uL4H0a8WzjEdznvvBf94MThqAAFntEtXF9gQRlyYXuI1Kmgtw8fQudXlxkhZ983w
C77e/k/jzO8prDHA5oY6iYVb/xyRjTG+IL9G7h0SwlqO6GzAB+aAYxohp/A49vld17N0DuK+1QPU
cCcLxuRgHXQajwQ1SCzXvRwix7FuUDYFP/RpOydIyahJBz2AJN773yoWQ8PI/CcyAtuAml4RH2QO
14Moj7NHMUtHLYEivoiewGqq2QnJNTJVM7DKciAH+bLXpUocyH5gfyFLw64///ie+61pJB7rtpvf
bpB5+KU79tJvmfGfsaNBme1g4LPzkVdLOK1kvbSzkyP+e8nlg9+khkSwFP90UNC57PRYM82c2Ghq
v33KD5jrXt3zphj++JPe/CCF9QVWg2PUmE7jSiPicfaywIjK0w2dMyA4eu5PG8KvunhEg9ve5Et4
BXtBqh5GAIcVqlMPfUeChlf7JGwGjK1DZTWPoQszSsw9302CeN7FIhOM4LkS+fKJsyQPuX4seri9
PCDpcBdwIbkdFYbYUBA1KGTFpY2MmiDl2U2hH08iujf+UCrNu9bh1ZhON4HVjNgLJ0/O9Hqyk3HJ
tE7hNYUrZPZJWjKyKUhv539JXxeT+ij6mHoXW+GtNzuSi62vr9GvstzqHzR+gF5TSJY0jtL/UGXo
fXmuia3G39i1K9pRfh6kGZe/Ix6ckeUV7sMLy64++Sfkuz2msN5XaiCXEsxZaT/8pMur9E3GoBQj
Gn5czCbG6fOTBezbbGBm8yKdNN/keiJMQTzH/yXFrx2yGMmmtKxjHi6iVC4psk5V13jI+l14XpJS
PYzQ1hF0Gjzs+aNzstHzVniMbEquBSX6HQKoa98TX12BnZIqwren6LNgxW9shth02AIWs+BRph2Q
HjJKZWPAUZ0pOxp/Dp/63/onwLeL0gAK1Ttcw+s5xlWfgbkWy6Y4yIGQSaiU9l+K+oNtL9/NP5zY
ysGUkE7h2ev+xiDlRrxjO5QUyjaAOCRGZwS/0znqdMgEXImBfgMsmgsZQyCYIUtWNkFjLw8Xc8s2
xDp4HwCK9OFApZlOQe44beVtvpsdxA3MPObxxlj4p1rXyCEmDPEPe0rj+d+0nDeTfzPD52IlvPEU
yi6mpbRuczDz/UjqW3Ua6gw0VGB73tiXBf3l79OUeCGVvy/27bwpJFZnvuwnIGKyRnDS3/VUTfJf
KXjFRa82yjldy2NRtmBYNJSKuYSsbKNtU8RfLMmmsPfYX4DblZX2M7l3zxCEe3SLtAx/UzuSPtcU
OlKwtpFtRpLr3M62m+QzG6wu2Pclq/Q1+KOnm8YlDHOPWLaiXTKlEptadDOjYoDtR2vqdzbswM18
2j2tpM0be3EeqAPohBLFbEt/E3XtsNtdc+QWgc1EfWHzV47ZHbLKVZJosIjSJLxmCnKGRGSEAwPS
Got2ld9764xMXnJksjTTnXvXnFx4Bi3kUP//hR511H9eqB2UUrCogitubw7wY9KroWDqb6plAUNY
mPlTzsIgEI89y5LvuZzrKjLUz2cYizhkbTl1P3oGMZ1/fmNET/2JdF4rCDA1SXogVdWgZ3SncF2G
yQoUqPH7w3/o0Jj/AhJLxLpPweqkKDbTNkU+V2Q33j7YDPYw+Jays6AAFvRWDEUH/cMIJri7mOYL
fs9iAAZynu+64av2tRhHrnkVnVC0RifALGRCuXxyQzbwd+Yr+LW9YpM+Kgpr/cbZucAHi8uEv/hp
kSyyKyQsT4MMU5soeETEHRQiWKddvhHNidxHGR7dNRGNX7wbcRnFcer6AzRXSO1MXLNDeDA4en58
tv7Ts+wEsc1PPeSZNFTuch6rlac8rdrM1toAFgogsI6bmVwgKGrpA990HQxdoO9Y6HYZuiltpbrq
mOqJKZouCR7aikHl2uN9UckRJ1ahhfyB9AQbzEVm0FdnoIwfpJDq7IGF/8njbGSrn2rtiyy6jp56
QP+sfPcxBHHz4Awz9+31Q+lbnrb3KJXiVF3Old8Dquuj9xD0BxEkhBRe0//19cr2ALWye1krnkN+
uc/vNUKbhJHbxJyzg7aJdegJGwXYJi6VHK1Y4X03R79r4tQIfwoBGtNifwgowxK7GjZoskiZAoS+
dcXRlmpP1Ln710sZLc7T9FLgh+zS44Zq32rn4yGik8zhjKva1ISFA4P64bfaACbkksGvNg4jx/2U
tHV/cX2cRTroNd5jZX+iaPiyMozqtO9LPoG5jTGt2DeFizCHVkYvQ731BYocTXQto8kuECz8qCPW
htVvp2TdIto/wZl9Ns31X5X1kKuAbBLFBLPGGA38cTlwNtGivvTs3LdWdsgAk07kuqjzcuuSgN7l
dRVrE9zcks72o/B7tvMDYkCc9CBPBiFafu/T1XXR5Bm9k4wePmsGDDK4QkC4nuj7voCYXNZCSXBu
2LWSGBcx2SNh4vPdqTRPnxBCgLChZZAua/kZ8rM7kum+ami5AB7nLQV8107QCvuq82tdY96M8DMH
dEgWe3jb742pPhTRReWRDky4QfazMSSWz5ZeWxk2f8eKt7NCSWU2NFHocb4ZsV0+Czf7z/rVhtq/
Vk09GLx9IIHPoVqDVQGlvAGArtFeFz3ilc0xTISMXj3+OGeh+yF42IZuiGoSatE8sJix2bKpmu/g
oHsbqslJdrWKHb3jx9prTpK6gDdo7ODtbqcHe+q44/y+wc5+CuEpv1mQhr/9KpnorLimez9cACRb
at9v3cyKyIRA/7ckhJRF+ipnqQK1iSk9/j7r5wsShXcsUB0lSPbutIXjinUviQv/Z8/tWpIJ6105
fH1gxnNuLNPW6rjt9V5AWCdU796oAkvqUoj47or8DKc1q0/21d42JQS+TbgC1eYEmv7quWC9nqms
VZod5cAV9Xxw61RCf3H5Jbik61QHpxbKfKNLTFcj1XZ0t/I0dH/J4uhTkHCvgmjofQQEHkyb7NPW
4E3s9ZdQWDNf1pTl43WVX33pwrfieMGPDTGoNzu6P9+sPbU0MF2qR9Fd7/G67iS82hiiVihMEk/o
ipPoag8GtTD1RS0tAz/dnESWXboSB3nBrmMtxviReEvXX+qcv4NWXiHM4PJFJ+jAXL9hgUxchzzK
Bvdb8mvnuXynFgOKQXdvhDwfBXEe5nPZNE1b7SNHWt13JGDHQseh/9/NZh9Ek0mlPJ9nIOI9JjlY
WAECGr50rKUOLU7SrKt8cVUXfkDrbP3oz4EEM83LqLdpNAthkVKFrzmOhE4rZb9Y4IVKb8ai6DYY
RkiPJ+GHwNu3rzg/jEWVXrVPp+de9DHR8efgbOw/Er/7J2PmZZnsiK0Ih5CwXGFoWXjWuNTKVM+g
87AWPtSOhXzIxCXj5gLsKbjv+DBFQjPB91lzGg02goJhuGnZHQ1v2VcDDM9pMEOUEa9olt2jY2L/
rOU+2D9AdsC0BeBzZtZnBYC+CSOubUet3jEwD8jl+0Q6+s5FPonp5RzRauvBt+uw4sAUctCcOkC1
tdUodcvB/CK4Sk3wlswPwkFOG0waj1REqLJm0D6wFrsHKPAhJ6zVEBlzXDT4QQY3T5KTrEsx1xd7
QsCmbR1qRoz9+ox94qlMOU4Is1CiFoE1nnswEjz9PlVw3R7BjKWkkRSDNxC3ZKfNrpVMu1YHxTEY
HxbcMiN4+2o29BlvzQmKyjr4hcBw6OIYyUB8kl/hR+3vNkqwvBvOzvbK1ozGrW2QNuOSujJ9WI7h
Ayi4iOHXtbwt8UnTK0ki1XE9XfifAUo5lcRYfpcrsOSlcgkkOwLN0nn6tor7etoS9ngwH+FFj5pY
jOrfTWGDIhXHB9Rq6G1+fBqxcZ71q3jyWzwg6LVAaK0Hw0dI63HMijMtazeqwbJaeRDsB06D8E2r
tyaKaeyjvGTYaVW9e3LdbLCYvRMzGPgk8Wba5msFz/bpsS/2Q1AeQVYycQ/LCxPgYcCkgj8ns61G
sB11UTJ1gpC9HGpdkk2Bmik09sd8z/v3ZJRvavj1OvuYcqLhArntHP4iVCBu4XntM6NrTYXXLh9e
1ahi+m6N6CQ22zvMXGEceH125zs8gS8ZlklwtmXxTybsQA52O6QBx55jWBPM1JF+dsndWWUnnF3o
L0fJFNfT94lD8UIljCB0XP8RHw+kNA8MGPbdqbqH9bsIVaTgQFOfuMIWjujUWSs6JMiuSeDPZz3/
dk8qlDZxim6+mBGJBuR9gM8OVtiUL6GnGYf/ZJUffxSryCdm/H/8wqYEOc50orKB0utFXGsRfb6P
Ck5yC+mOBCeglnLGXeQXJ4ZAI22rskS7NohHqaoxXQsMfszbsBnWee73y3Ni31l2+23WZAFhnwi+
bEBxXj6snKQwDigOwany0o47sH5BkXaogtZVwtWG7BsDH5+6VCJiuc2k6vnRYljolTB9SX0Lf4Ui
i+UGVbX54MF9uzqQjwOnVIr4lZ59vz6LtDC19wfviEU1z4qVwP/sBkjc+tUZ9R/T2AWvxtuVPH1R
aiOcj67NAUHvWN/TqYYXG61No71Cdf3d6Kw7hi8BPxq2FLsK+fbPQPmNRMOsj++yYEArflbu/ei/
6fdyizhHOa353oRjvWSRYXG6LP1LJz3hZ25EoIt/hbnHPgvhwgXpG0u0AdLCuyQDQgHsbmAWZGjQ
WLJO1Xud1S++aMU7TpqE5JwSST1zzZBpbiyQXfuJMbTTQewDHAyjX9pJn2zlFqa1lRZvFCIliy3J
0ezaCGp9btBWaWNyKyuh2CPlD1VqkXVCnl6Td3XdZhXj7nOWrM6PFTjb2T+BlhuowQsks5ZExY5j
boXP2D7Hq7VQDuf19BqnUPlU3uFXJobCq6aA+ccq8/kHMEEUVJUj/cPLl5tCDrYuIJARsm+7o2NL
LZXHofdHFP3vugYoN3elIv7sbF9QlBH2PeuCHmbU+kCtds9qe1gkWJLEvKUggvxuJ4i8kGl+S3kq
OMXJpWP0UnFxCKs4rn+ZBlvT1IzYAX68K0eV0uBegj/wLFmKi48rGwNiT/5u8icMfdnTUiHzrbbR
eRScFE/EVykUhGFjZkoITVehO9f0ZF90gkNi9/Yg44DaOSdNlyLncmsWLDBjlL6gXe9t2/77EBbv
nMspCIRoSY+WKy9B3X5LtnDbUWqg/5zyhFs/L4c9XemUsu8VG11+FnFpHqxCBwg6w81vZWrRaaMQ
SxmSHUX4fDiglXK741wGHL0+Qq36vfJpWcI54aJ6548CZ77C8qg0kuQys4UCl7Cg+PyS07wOYQ5F
nV+/5kiXmZCSv3lwkp+Un1QJ5RcOHhs9/IX07Qb/Nu2cw8mKOFPHkdyWYuoREyanHXDTBtHP6G+T
/395m/EKlnpSAd2SAIF+DhIph98jcTKmNjs06k3GRJ/dFB/3s/iQSwPGCmHRhYtx0oZlVkGyBHVo
4l0xl5lY3PRk2io5JYHypixsvLdhrs3QU+Dc43ylGCrmHOtfGCZo5zdA9GrPNWr5GfN7vpYKT0pA
lxX4D0scruuw0qKR5jdivQr6yJVkTDR0jzcxDZRP00YrU6y9XsehqiEfW5jdoCBmCdGRLrzTpCXR
ZQoNIztIt1mqKsxtSfm7q6LM6TCowJ5cjC1lBnM+wvICtrCMR9WwfL7D+1JUldfoLy+O4PAzBk1k
AnOFUhQxnmHKPW5oSJTacrxE5al/mDg3u5gj2dZgT4EHTt+moqMsorCf1+nIZ7eeLaTJi4aO8wEs
cDizy9lz5I8xU17045KwxrIzkCOR3foRQ6Zi7roD2z75GUf3H2MqkbSuz21y1+qlXi1CHYfVwFeu
L1Pr1ufisONY3qVnSzo51uwsUJOQLA0azo8cCL5MCncBw/su8fdQXbJtq5s13HHFHq229/bAYTXJ
x7/R1FYh8nEKPQWDbd/e4UxtH3fsET4UUsnwqhOima0DbQNIElz/sK5uPkCSopLIEdko8fgYEbjG
zAfjDFU37h2QC/4K3Kvr5CXoK7wFpy8C87TpBgI2ZM13BvdUgtzS7Xr8HPFaR4dalcO0d4JHDJrW
1iXXNWE0PsaRDUNowGmLLPVGuWXvxUDElXBt+Kq746gWI9Pm+r5DchmrEWQDneVhSO1eZl3xp+eb
wbYS9+T26JXVopQb/p61r2JYFjm6n+zTFhRJIgT6T5TxnZUlYXRGLemZpMXePy89fuORjX6yieqb
56hx7m27sSkRXUGMNRnDuYw09d1XA7zhjl/ymV6i5c+2XmHU70qYQPcV9f3JLHfAPB01sZnLBskK
t1Xfy9hO4kjpgSjdr6XWSNV4uydNHnNABY9iCk5cxJTnJpT01SoieAJoZ7q/e3CoSllGLV7Zg73T
o72+aefJf62VFvVjn2K/buKJl4mEiwiOzH6McBmro0p4A6cmaA19eNfTzshJoOGt/Ex5KVUHyHXq
HcwkA8VABUXN5/bCqL3bmm06RenNevC5OK0BT9H43jacQf+XyEu4Fgn2Zt3JB8N7w70bF7u6seCp
s6bIU2/KIqWR9zLOdED7mTcPuU7gsaG0v6tTUcLiM3iZdy5IhYC2u0+JU4dGwHrzsKviMNzgQWFr
/GSG/LJZzvgZ9YC/SokqLwoFtzvtJokCMx8cWcrVCtFk3xzAFC1wK5u2fqnUrvLILmIYaQvyjfsm
4drF4e3oJwCn9gMfYBI9y9KyqezRVd8vEyniJgkCM7DiwUq4kI3InGAS5yBDkQO/aslLq05Pw4zp
7+CGWNsQqMkJ3zK/Vmb5ocFymedR1RjpJFdTcFicBwlO0puSLOI2EuAHfcatzAJcgr+ni1ww26zH
Z6TAmyG5LRPR+HyCrnQ7d6GN/wVr9XPn2SHqMFwPHBE45px7fBZ2wdfVyTRDydWTCXNZ9ZAnbF/s
ZTvidumJ8Z7NrSxmBtXSIdRth2BG9orhB0mYWwYyEi9jqraZyblnj1B8c80/pWNc3KdO09QLAai6
KbqjGlHKl5S8u0NPO5t5dX5/TtKfxrofXrAcvMJEjE0JsksnouWYcr7AtrQqy9iJw9BmsSPJiRf5
w6/UssXdEy0YHfASbl3YJc5ePyBfT5yKH65ido0ytTpvdhNevbMLHbHoalUwGSKhkIwIjMEf7pWe
vJQxXDWoOgdzOWBvJ6eOfYb7njXp0xkk8S/XU6zIxqDdl4Kp6lpd+uvV4SMl2/GoQd1Q/w8A7JHM
2DkQch1Qgo4kEVLtJky2s2t0aiMdO3GI/y+cCevMUet0avH/9RKU21Wu1s83XWaYgdfKrcM2sb02
HHs5IPgpsnwtS/W5V4x7qWQNa3rIlO8rGDF9PAPjtmYEoT+o/zSLO2NMJPmU2Vk/lPpxk43mP7JI
tM99/bL2+7wzM0Zmeg6R2LIeB85bwxAMrkl8zf0HfqQjiqyH9FeXP3g9Shh+h1+WgId8K+fiFmFq
wgCnIuTvoUtqz1nh6z/qR/a+UbWcHhIDBVPqzAmpUHIOLEBvVDbBmLOnZbcuvyoYp0zBKnFL3nCA
xUWUB1Q+a+tMjFvNf7JQQnMxOded09RsFYuA3B1si5jl34sFsZnDRu0Y+219qMdp6rVX6pvgVfzL
JQYIChe3PijDOt71csotvIt9GUJsm/jyOkejNSREVEQgpDwKyE/gs173t2hUDW4FUVFMe+ZkgQyF
2uVAnjwHbsZcp0Pw2Kz94JaKYFNq1B8E1kDSx28FtZet8QSZ5+zS7MLyQclL9bUdr5w+X8PGpSTL
3PoJJio3cTVQ18F1Tq9wo9+JyZbsOjWYzP81A5IJTphZrkWc+gLb7d2dBGIxoTY5rbDyxIEmDFQY
oHtL10UArWx39sygqXKtkk4B1JLAU+9NXyDn3rQY+wBsyECufJy49Hj4Sr2SE4WHef8RnlCaoqQy
A6raaLi2AUPv5TafYRQm8T7MKr/fdoyqKA8nc3H1X89Q3ztcQnBBXzeXiXZaG518rnWj6X6EEIBo
mPcuwEG3ktdl/UJJ/O0qxY8aEoCSR3F3PBJtZUqc1bODoLMumm9mzoV3D66mFsOa3C8Z9Ho8kG+a
J4jWQFRgOxMlQwi7bmS+68EL/eKdcKAK2C/5jjVO5zKBhRV8JdcGONcz/pLzLd0pNHAkwEyHwO2W
g0emxqPP1MtTgkZx5DwkPxDMJiEPYpN3DQa1syuRztzjBQMS1U+TwGl2tAfTGfmbMPKAcfBLh8pI
1TIdBH/uRCczmRWmt9tf2e6C8RKQOZplLqKoNywglQVnrgofjWd7pjKK9FJcHiNJFXCCgeNZuvjT
26L5bnwyx5w/7PXSif408JyUAoxOROMoaBJNRlUc+cuz4VKRaDmJS0fE+J3rYbQ1vcND+A06kL8I
/X07AD12bXt5S031tVw00zsnkRBkKS4jE75oGJ1vrK3qyDbz6GmLAM/NPKKCk+aJpDphH/GdaCuB
8BklnQa9EJ48WDSp5CFBkxUceHmJ2MDh5cCMmfE26mgHPFwe00rM7lOocV/20BVBxTR2su424WO9
TqASp83g79BQiwhE5uksUCEFktz012HYJj3c6NcHzFTpsnOdJJaI6SK4LlfIS05nPjdYXJeXLdPt
iKchDkmTVqTLs8S3l4aC2XH0Bfwp473wy1tUpcCPLyk7jS1FdSlcQdXYSA8qXsXnwMxVEjle/rDc
flGeGRWdfoCzQQX8MmXTe6pOZhi3C22s5opHQ7QhfXBQhJSW3JNSPVIsElB029ssD7Fl1IYGEkpg
u4Y9qVftblBmUvbeanfDEMi4CtHXvPhHH3HS9FW+4a3JG0yu/0kixuQXFRJMWifRcbPQ31aDER1t
RAhaRVNiUVkQOiu7Vjs+9UtC+VFqcs2z47DyJ9TF33WL2b5G0EZhgNiIoOXME0Y+TDrm7zbGtqcK
ACUvSzBbMHSmOgTfaIUHYzqw+WwBlRyVSC+AHM7QQLaGBeBtaCgKMaS7ndJA9uvQHls1pwAyh0QS
YG4JONhbz2yQ9YokhQMh0hU6Jn2uwKWuDTfhGZaDDHcrOVHsh81oyFiTa/PA99L2pCszqO4xusYd
or9vaKTJ4UR4nc7d+ZBSfu/QadZPZeJFpxzmtwfVfU8tXo8O6tb18+guJ5FLr8eMJTBlvzFAwLpG
NnDfp5J1D3lLs+tvGa+H5bCo6f3khVIvilr7jt2fl2vKPfpMTgW/gsqxxyjSsJbJHIhHU0oVxwjb
/9Mo91CI6FoD6YKdZGFcrBwe41ocLwjkQJf9UEs6MhTrSFeY74yGfVXRHMLdEPZ1G+/JjDEfeZvR
jBnhjCqKLwjGqvCfmfyDGT7JfGn/PxmNpILM12DLJzLLvabFay7dNZIWbYLaEqQp0wjoTLmoW4P1
n3cTr5sd5+tH66BrOJlNlk38r6gdCkHwS18YpgM+kIHyXN717EJW+Xj+gzOKaLxRmHStDjyvaWZw
tsXNxeU7O/+KQUoqas7pw1eOxdxAa92SL+afJvDiWfl0YailCH7THTxDTDO4OeMUL7yAOTZSPWJI
6UVRIQ9zfxqtybDr6NOA3J2KMQaR/dori+wKOrANr6c0dAJYYTLGPRDHtxqWOAm3SVi+TxH/El+p
98PwEpKdNFG5Rv754mD7BT4EEHuU50F4oaRpR64ExLNLZzJ8F3cYqg9ExE7DyNPD3ZJbSNGkjaMv
a1TiA7v+KjloioEGAN60/hKkOlVAfI6o1zCAb5ZP+xxle1CnqNZcxbVvmrzX8zkTV+7womu5vs/k
fb64nYP1SNQ0QOhld8/kKg9ZoiFXm8rjlhXp14SZHYpyyXA7lF7Z4HfD5yr6yauRCxLShSJDuXL8
ByNxqC1uEJn8ntqiMrGjpBDwHt6NVaEPKjd0YiCSOaL9juxPrilh4v4b/JslypEHphJN84NSo0xC
JET0llVIsTzHPsCupDvdFddxw71sYOLWj5MhrfHpLHX/6LR4/R8RFZ4FMxZnGRq7s1wrTRd0rJ4q
NWA23e7/FZnlOMKmjGqxFqNV6wzRdSryzpZvgX6fGuNn4TBkbdrWiQhFAgTmqaL07Y+rAi37znTx
zw9EP8P8GuOvpqhge3h1yRNbTQPGA+nFGrx39VW13McJJHS+6fOPZGGGfKSlJ9mm8pIXsT/qEBK9
TlFxjyQmv0kT4zjg/q3c225btm8NvuVN9YjZxKu4W9svFNJGtSozxws2iSlUJ/DZZ3NUiCqVQ9tK
t3hAvQYI56ozNm5Fo1bTiNAIVpoTEQdk+P17z+EBe946griqcdggqaKEDQj1StIsPox9J5Zm1lPF
FOCqUVuXns70ZmfRE+FMHJ0FOMAUcdP+U2SGGpcZsxyokIyVb6ZHWhpqAj0Hl/sWyZVd76oRJl8p
A4fR79y171qBpxjETjAzjl0jIz7IHju0+xIj/CtMVdktEJV56yw6OwljyRtCQBkwqzSnnI/+pF1t
RQDRsAg59ji/+S/w3DGn7GiCJ2z+Rpyj7z6QO0X8YL2WZ1N4T5QMUU6IjDmUrHsFZxIWfAhHUy1+
SvDWJDnyr57eW1wdEcPbiFKc0zm4TfaMAZz6o40qsTnGiEHbWsS+fmqqR8JSQutOcrcFxcJyn4pJ
1LiK0JbZ4xWk0ijDTP4c8HtlRjqx9g1tkbTcM8Rszio0i/1ADBe6qdFKeebeD8aGj1A2uP7scb7R
eEOYlpsKT9N+3GsyhSQK/XPDITG+H4eLapJI6aFP/O3pFyi/hc9C8EVG2ac2UC7YEtocbhhTFgsP
I6b4XH1Q/TRNM/NKrbRars6JLD+aYRVvGazC3P1nYj1Diy9r4W2KXR0NMxdRJYO+LH3skgWQ9AaG
zu67T1GIoJXt/EEDFfWe4ocLrJPzr5K7btJyYeX208PQquqKoAdjqzCcnoflU2te0+GDOzbTQeXx
3rXybEIIcyc1G/S53UsXNdewnRM2f7ZS8/CxVsdItcSv/x4SZ4aab+rHhUCHuZWKvuEsIX+GsxoP
83xHjlU4axEXM6xZH6yzdY5fGgnq4J7PI1GaQGoLVIcdvoAryTMOt5RwfriA4FkdJLURl7fd6ctd
SHz27vxXBo+n3bwgyDFDXCkM0RFJf622igwcoVZOcIPf595LbEq9sV/7YWJq+WOhpo2OGba9Tgo/
TgIBwjf0vVIKIK/6AjYsvxgShsLiWO9bWNrRdBz6zIOl+Lnrc462+8VjugajPfdroVIttC9gAx4F
XVpTJc1UnetWaUrDPX3OvFpUd5pK0pnoOsV9yclJdvu9snkDwIiVQmxYBOZBt6TK1WeMGdkzNmfK
fGDo/F10vXCVqmWPJs/LQ5C5QyW5gC9+W6DYomRr1saYOMOAcWsjm6WxKHAYgoCw0shAH1cT+nIw
Q6ff0+qk3z45diHjafQ0pEt2CBanXJtrBIdS7KKkJdRZnYHUnCuHwuF+pFoUg9p5r2Kjp2CNMGxx
NrKSJTXWfBcKdDrRct00a00DOkyEGGJ0Nhwjw0ZSoNK8T7/QJnXDIK5a2zrExC4PLSYl0R0Om3e4
wpoSTHFFvhohkstJlu2dZaIUKaoa+smmEA8olLfGF5tiXVRyOqi0IgzUmWQzYPGU5u0PtXoRSzcG
Mw4iZkUjD/UoXscy+D1LtFnBo67mRMwUrgUAjoRDQGOB4K+F9HKy/B9rS3FpZJsVMdgt+pOLqeOo
tMkZQFQtam30HO7WkEgz8eOD9OyBdZqlSL2+TL0mVEtQbzbbtqXybIrTjFsrfKa7O/JFgWLLgyMr
DyrAP7FPpiCFiODCtPaIBq4NNDr+QwIIKERvR4mhjN46DFNrfQaoIuXc7/HbWQE7/kpXzwctfs9V
3J3GzlA8HpFwLl9Bc1iuMmgp/kQXyfXyaVlwjJzlQv12ROld40b5/z39Annmmhp/hhK0Fix3tStI
cSkFrZybWlOrwUK0wz5lg8yOTrJaTqQcRuX5v1gv1C4nePDe2Pk/OHhks2b+0b8Oe7HvqB2SuGVM
2V7DONYYzzQhXQf4ljIFxx2RKUTiBcAe2UVHsY/WfqbW1lUJhtz+wG6ugFrXbltOEGfwyLKoWrHt
oOhanj3YqosOLrcCPgFg2OT0WszqSreTmpfUJ8BnSBpEx4Sb6b2pFBY5dbCkmQ+2SjC12n/J6RNL
67zP4wRo/qvMmHV9CNvvXS0XSvGFytshUFpax+IEaKJ7xyOHWKtJbhjUAm18uWRW330IwFdm0f3J
pSLp8yweaErKTBT8KlcavYKpuBdvpcZhIjep2tPYN8DyycoelugbG9DMMsixtVII14xc2cPLE9Vr
2EXNPXxu+eLIy2kpwf4KaPyiZ5X2dYxyZT2gXaF6clT8OyvCFUAJxHhUGq/tE3YINzFQFJv1/cAZ
lqkksF7LEzXgG49DXhYuIB+FQZ+2E7H5jb6iHEnEEx8TowVJxintwqc+6L3D4aFTZ6UG2oIy/nB9
8MsBhyf4+v1sFVZeeT+k20XFGM3Wx6ArV91+9GTUO9qaGSVZcJbIweDI2Yk3p+2mbFE2WPVxduTq
bNlAiC3jiybGChdCIDdAwTuHXkbt8/whfb6nNRKw1Vs6e61w3/d08x1CtfyY66G0TokOhMiDUM/n
OJx7lDPIBKg+VkUZOuDBmydAUCWKo6ZGPyWrjaAokoagNqIszNhJyzH/712HY9uBZOB4kEtmytCd
YNwErH3nsoQQ4MNzByCZ1vPhM7+/xvc32EkUFtxuP1GDBPUtqe4orDNLZjAyUW6QvOFZfDQjz6vN
+NxxQV8VDJv69kipD6vGcarDUrfWuowo555h+YUc56P3WOL+lDuzfUaEHVtyLdmBACdBFc5rm95n
1XO3LV8MSQefq0EMTJrdQWmD15HugBLhBiDk7GCdlNB72NDig1nx47ghtm0VE2dhvLdKlFasehWq
EyPDR4gvO8p3VMayFSL8jns9WD1N1kbmd/VJtS5sdaqD+uVI4C2/uMEEqNcI7rasGsQ4Ml5qpOoq
WymdQo2QOBxgVZD04A/Hxn/bhDS4CkZOCWgrLHD/Y3H8mwa46ED/hMM74mRhjUX3Aw+WiLL+d3n2
yJPpWis2u88PI8UgGYInsn0hhqqqqPCI+jslSyjDDNHlDnfAISKAQ0ybnBXR5HxECUZBcWiP6Pvx
keGTPjKgnbKZae/phk7gq3Dnxto4Sc8t6TDK8MbX4qnCj0daTD+YXdvEMErOL4d9sNSp/S2qnxNQ
+D/blDe6ieOFrCjA4MH4gSjkn2abffWmxq82MGEojNWcNR12fiPNgb04IJ8vIrS8gGp6FlUp5b2/
3zI0aYCS7cFnUqOorbFkiJ2DiqJeK5FxOChlO8PJ6MjRygDymkiNPwndcBU/vU/ukAT6pyRWMXgY
7y2eBmRCaNLBBevvHsphMGklFK3SAfk5Vncpostf3g1r6ZOthF4+q7DW40HxgOUMicbKL2RjP676
g+AlqT1e/Dr9H0XKLINZVx6CQlDDHA01rY0ToajvFg10y1End5iw5xysnuOx9t/U8jFpZS8qNkhL
VF3b2mTBIpY56ThzMGgNFnCDIFoCR1x/JlJ01A8LzsrE+lo5lMv8KSP/PC35SGILzux/ZuDvWsaP
OZW6lwLvOZJLsRi+zXEmox/84V0PX8Tdsix/zwMZTTBpFKY9kiLt52MuP/wRsmlyag6dbRr8wjJF
Zk+jmr/Zo8Ftnqd0pjg3xVp6pHkLS4PXQTOyv5nRJU8Y8gvr187o4LQ4vmsBu62tRZxxnhXhQdYK
TOxVvh2nsr3ZAs41p0/rhZjvVrR/fOSPuQ2aJMpetjRb/uSdITaGqBT6tztUmwLaffE6bXnFzmZe
qUCsbfRLi7HZR8gXG57W0OStgiCjyGeeo17KqagODH32zLkkxhCsFhWUpbLp7hQM9XqQB4Pd3W+N
H9g+s5QELwiovvGXqtaqSUd/CFCHEN3F2zaRFlZBbedjtAcBuwZuqQMgKrpRU92ar2UKFHu+flTJ
s80OhucBHDOk6ye2lSpM62L4Hh0fyTrU00uyNuuiX6qlgMSJ9Gsb6c4xK+i2cbr9HOYTRdhUXXtt
RmLNYispt6IbzxKHEaptqAFKFzJxakTDiavMHxT8B7wkJMX5uxol+kSNH/aijUzcowlb2SX8hBLi
u1UQzCW6PEln0t1MzaXLDjwXHYTwuKkuC5BkrcFPsbF9yFWx7N3gzww4fl+r6eWOPkk1HJst48vb
JaUKjj46nj84y1N7tyAs2MNL/OmL4XJszu16HJV/vdGIJWfPAnCM0V0jBQ86wQ7v7qEM8CsLO8BF
QRpcEPkwps9cUIvrPWFUikbUWokszVGTDp/GtMjDEyGG3ql58byj6fWfLg89WI8zQx8rrha8Wyr5
eS2N1r/I4bmdWyy985M9jeJ9cfG+BCI8/9hSAIfCbf9dSEDpQVdb8KE8UMuXI7lse3nWP9knFL6n
4qJaS2RKlio9VNAZ882YaW8TPqI802bc2qqaEEK/EpwHTr0/0GayIyLbg1RENhSTwE8pXmt18QZp
RcVKKmnq7eMaT43SA6CUrjWaFbZu1gGo/4dVIVPG4N2ahfxALmxEjOFIExygtcdei85+bH2aqqSw
fHw96bV6u3dyw8mkAPILTtjvgWhVeLWqaVu3ufkghPz8kffTyZtYK8KfQIgLciYk1XbLIbXWHjYd
mYwwO7I0eEi1GcYJDKx00X0alHvH90Vpnla11oqGhnDA/M0vhkOa2b/BgmjeMVrOEOJoxXaKBfSL
/k4fY87H6PaBewFElfntkNgJyDbBBB2n4oV7gFrsR2yxPVtmgT28yVNQ9cBYF81umhDLAP9yVfq4
NaIuhCy9R/aU1OaK4nqf6eVClkYVCaGh2cZmhdukFv1WKhIT38/0iVWZRH0Pv5cqvSGcKNm6lfc1
/ThihdI88mQPwt3LzmlsN4yGKL/i6hI5aV8osqA0wm7D4PCfnGv1VcPBECRY/MumzDvHuIWIT4cW
Ob7hitDIK7AVBfXSlc0QneWGvIIP9jRIr6CjiyfCt+v6CcKEZ3Dw4Tt0aSzmUR8KC+FJBjyZoqAP
g6LaRr3wIVhjYkCRbzGUOS5+YrYrXHg6Ds84feIMIlQUy1qqfwTdaHHBm/gwSpQguanOgUg0aBKB
8hQQLEwjQwYCFXIihVOngnoTW5tOI/8EsiXQYd2uJZCe52bM6bK1QYAUG2lO5qsgnKpFcvVYaR1j
yu32Dj4bKrQOCR2PDvW70zCt6At1E5OZKwpdQ+k9+wZrJKQfj+e2NLbq0SLgHIgsMrDbONuJMATs
BGezX6yH0hAgU0eyzDR8BF9GfPaC9fmz+XL4XROKO9sLpjWPJyxJS2g9H8SeRLjVVP7sdTNDwCZv
erulfnl/YhCYWcy+rPTZLZxsmM045GevMKJz42NyNF9tYNrpBQyDYWCLgt2L0Mv65F6agZc6F27e
MiqdHaO+Cid6UiDEENWyIq1YTW/a0ZuKTCLQ5Skdcjiv+huBs/qBrYbTes+8F1UNC3X5wq0vfgsZ
vlEvuqPlMPs6+yz4YtXs0TpJ5wM5RwdNmfye45a7bnHPnHIILdcWiBNm3uklKO+N6P7xVW0N3ZB9
s7W9nNFA/aVk6+Wf8Xh4IDbeQNYA5RA9eTuo3KOyDFLuCQ8Dduz33vE6sHBt+cZtvQTqNvY5D4xw
yXdyfF4WNHKVnn5JmAgxHBGv0LlX1hIlnBUjNxWxpHQ6ustz4RIh3tQMLV5MIOOJYUsOOspepWk9
Jfsd31AoXXUpZDlSdwCV6DZnLI1vG86LPae16f13z5xX0ffob+5C5CGgkNHSU6oQWPJS13loGU0g
cbnjFZCIllpa4sFs6lECD8RDlNzudb/9WZ86++YL6EhAVIfmZldoliv5WyVi5eUhlUmwa5k+kv4O
bMBq4kHqmNUm1gPVx4aIPfSzuMYrBBqcmVJCjGtqciR73hRZlF/71cOE6wU00YCBeCSR8DvfVsGR
bZDOBy8LM7tAMsA8pqng9j7upua7UforJIymSyr+VFCRZQZECQYRpSGMT59dBCUxgtSjmXK5JM2V
88ZRBEpBi6Fj3RAz2Pw+/6ReLABbT9g1E9NMA4orDfDHDw8tNeUA/vRj4QKyta+qMz2Mq3JW8yWk
dgdsqbtyJgQpCf+1+rrdQX07KI13Vxkp52+zH+9Ll9MoVHjTHpYfcwRWyKrqEyL/QN0w7oEse4ve
QugIbvYBjbARX2OgCmvGzkI3ZxQZc3VzulfMOI0T7CeHsA+xWCw3WSfcXwQWJnBWZam4q575YNhd
KtoJVWKUUHPGqDl5rIyIV/FxVm8f/RJLFsSF+gwVkfmMFsMD1ZJ6K3LOgdZp+Ykss29nHF4PEzL0
ZvTSWM+3mmS4SHR+W82B6JNaoPZVRwS69hy0jr6R3Ob0p1ya73KwOS+xakdzfz1iVUqg7ys8htgs
Bdf99ifmTwkzAlmkL4rhEQZ8807zXpHuPoWgkfG32UU5cPhsoCldB8FgOayjD/P0rNrhP7irmzIN
NibWAUEiCHgu1GvRr1ccVNrOilw1SXlg9jCc+M40QStGaHVMzwoyeF0uS8C6RBy7F5M6PapDxv92
v7Y4imO6HJMCTLE7+w0Ixa4Y6GYMs+MSodlyg5VoxEtgsCFNpNykepgo6PVjsqfAhJuofDZL4eIp
7Gglv4J9iDN9DrtOjFeBp6f5gYVeWapSajJRAet8gyD/zPR29f7qw56xhY40Z1dCbOG1LZu5Axen
wraA5VUJfY7+OJKyt0JIN1sNS7E/ai+lqMTNuLH7c3NzmLrXYV8SmJFhfZRSO4lWvBci3W+i9iCw
S33MU0eP89GhhYU9Cmw7PSxaJwVektBKOZev1nys3VlZjrSvwr2kW8gHGcUAvwfRv521uazejzh/
pqDRrFVctFu43DnNfsGO+j9Hq2VAEjxFHrh26JST+SWESUzmT4I4DmzawO+RJzhiigfAtb8tcqCU
PyQzOMm9KDJ6D5/tH/BKuPyyTeH7k6DjDoksuP3jms5dW9ebp7Wr7ECIytHn1VCeZJp1sGxMelAX
1BgFh+l47TXYn2MGUM3puHE7LjWA3u80bQQz7VsVu0SCmv+rTkT65foAg0aldhP4nH2vA7EOuflz
cQuq3yAHBLYkBC9y2njp8f7ptbbaImflFMA7ceW5HR8UD/eWkjrRB43QI5bE7iw112LQG+ZmxaTC
1Yr9WbS9yE8nczjB1ey1rvMQrSbZyPYVXJ40/91fB1dB9D7YvVanXonI4j5PuNQVHHMxrwNPHQWD
SyhoO+C1cRECIBEnuBFttW+w5MDVp1WlxVTlfX8YEilRxDeMmXD3CcWgJtzYRB1KnV+iAPbe1uX4
K5tL1hklTUR++unFM2RRlCiMId9AuIkK7fYGxZwzzgAu5p1U83bLWytaZcoGIXeIrrmpDT2cAl36
3mSPLTlLbE42rJHo+9jF3qErcEU9c4cvGH3tOxJc5/k+v91TnKu2Iv9qWlb5/Wak0bQaMYzKixFV
wKbBxXWe6pXjMHVmwPsvBaq7vJKCQtmzP94jXY5RTqUQdvn3fnUWvoCRMQYN1eKBXXymsNJVPKZK
P7oIhQyAw3MYyK7AbNrzJ2UXI1uE0JEEQkPZLtWwlo/S0D/ExNx88e1HBw8AJdpW3KHwpkw0+Z+e
jJiQZXe3aaYV8/yPdaLfq6usshaXSo9mImt0hxTn3xn6fJCbPuuUu9D8X6TKYO78FQLqButxJHJH
Im1Gj9jZw/V1a8s9gOYzQq/5uWyc0Nm4qCA+vhRMwn1+TVV8yD8U2KQ9SLbQN8QgATOlSzNox7Nr
wjKoDyjwUT2Xnbz57YW5mQmNfLImS0T8wa1pT8xVSAdOAllb26bn2DuPggYhscFLtAIoGsRmhjtY
pZPG10OSF8mvOKmSA03PNfdgmGj6+DoWJ/d1MBL3NjyZ3n+hIP1NcIGIhDUSgTCCtU3LzKAMZtdT
PrxZ+1sqbtv24cXdUj7tWhepgafocTdaeacCbC9REyLsKT//rR4bcgfNgV6Hs+Howp5YtBQZGYhM
JQOX/bnNTKXwyF9BpIu5Be28/4NFV0qdozQ3MDyTLQJwlGQLzyeCE6oSVWHJcM5niFlTCmQETV2b
99llwiGvIN8NNd2psliMQqju2z/1V/7C+AluOnqhNjIsNo3KEgRaHb/Q7b0NZz/jvDLDDLUmsTeV
v68QKyRfOSdqoqqJUlsJUWopi+RaT3rzRuFPYH+M5Dl2SJr68pp6OLvuJOgBx+Aym8PDJJMEfjnD
eepSLahXP4BCEommATkCy9C3NUBvoqoiGDlQNWthrZuoWPutq9M8R3LsxaAU7Ug3RSbY0be8s/xV
E42ikmTZ1IAPZz6wh8pST3TRHHi7Doituzb29A94Xqsg2OvIQCTGoH4VhSXq88rYMoWd6Lm6eUEc
2gwnVwvPWKaCc+0yAAdN5cbppC8tbhGleAf3fFB65hw+xrvUU7zJE/F1ENfjFLp+IP0yNMVVxaiT
8VLqVUrdGEJcI4irSJ77kevJokhbk/v/Fc2EI+8/NFwXUFJLcQtZvGDQ3FoT9YQIchsmJejuoYjh
AWmFDpS+wSfJedF9hzWkzgA7utKLzZPMUVw4d6Cwk5M8q99DgNdQr6dEKHRKhD3L7hHKKSPikNYK
xc89xA6yBAjou+ZBq9oHxQJTdxNXuT7TnRU4x7ri26BoFZIEjKGs9fsN78EjmVABjA5oBVhLBWBF
C7t9WrSABnmqNxkRhb4/8hJ1eqyW5oT59OAKb+5alYRvYwH+jY6lQWKj4c5JBVQEBO07iEml4B86
cyU2MS88tLzQX9iBWxd+YPyk8rsA8GBNy3xRnHxN2aMbeD+pETatK8pRzjo7L/TXGiG5D0L4d6WL
XZve8uSsfgxlroY89NQRTREcRf9hVCF1y2glaGwtrIgWADowxCm2U6uHKqvuF/P79rVw75rgySOK
yQ7YOmo2Xh47ukw/6qW5fXxYmihv1Vd1nNmPSvzJQL30JvKTRY+IXPSM/ZUEZaI+cd8Z43bsPlvO
yrshn7jNHQ1sUJodHrwsONMDuyeRmBhi6Pmj4R0shKByJEfQIhW46Jd+S/7+t1Dvm7tZ4BH+ibZC
lvufjbwbRIhppPWz7x7vYzMYBokpOMa8v098aoJpoN6L7Eeu1/k2kWhkrD/AkyDCUmaQUiocIqL2
gTPoQKL8HZfXIBRMNkWYGkTikTLLoHYk1XX4jeSe8rTozpnzt0yIjzSUXkjv0ee6EOBLmxIjh/+2
HwNCeiVL4VqNEvPUNO0oaD86ntJs5kiow/le/QEPpBchkRViXQhY3seGmg1BLGtb/SsMmEVGWvRW
nAgwV/BXvYEXAACC/vogDj8xOxkmWZCNQtC/xIPZVxT/CC6q3eMYZfYdB3bD8snzCfRbIakqQFbB
uNg/ZU0lgYqA43tFzX1wZn3/Kyoty+LTBylhS6pMtdfGQJNhNxLF3f1MKwyAUHd9AmRK5FBILeRu
AyISLs4zoyp0rg+aqP5NFtGqGSps/4aZZga+HhzdEB0oJYIbqNglZtwMET/+oiFpwZEGYQDiQ7E/
+J+jcIBmvTYe0ziJfHtoWPDirqXZZXgKF4ywdDX6OmCNTtpQoU1A7QLyz7d6WdXp7RPCTtaciPdP
KzAXwJI074zuuI2PwkUT19ujqrehZaIF+211SZzM23Gn/iq/J7osgXpx7wMGYMJ73Bsgqg2DZ5eo
PW/rjDaKrD22HyPJtZApwzm47H2oSIsw5XZnAPkBs4A0Xz03gc32AQ/FkEmN7Jhwe26YG4EZC+vG
X0LlX/glWl4aECrTA4aNW2lyKX/uJJRB/VAfdbVzkzjCtHhTOkHMFNsg6X+/WSdLG4hIoRWtMn9A
l/jMbZvMbtjYqwraKJFIEUxaUkBMKrH5gPd3ZxTkO1ga+D5+UGRMhQuPDeWMBPe1rUVZOGxt1yuc
3eXYI6SRaYqHIFs6rYd4lQpPuuHDRfhljpvHRsb4NCcII6b6c7mUBoDpFR9hQkg773rDHteioOoY
e9KlHd6K9KV16Lltg5M+0aM7gmV+6MJHOohNHzAHBE3YRI3+6obLgSakS0GUaFYaeySMkxHbhxAX
jWIKtC0LxX2NkqsIfV+eeQOw8+56Ple8GlNwLjSEM0v50/Ip1S8J8P3nDzceIvAFlSrV+qQDS0mW
NNk5Eop8BAsKN0MBjJVMpteFYF/jfSQvUwiUomV5XfQrfkLVtCmnVlupTIHQ3d5LzoDeHZ595Un9
LRIz2qyhyLVbptEAxV3WHWvrRfvwDlYSES8S+pKWSd0yzFA0okV8GyvvAdJ9IwPTAlHaGOHuOKaK
WIoKMX0ep8A/JhnbXeG4irnp7uhBuNhiC7IVxictSp9TJrmXBZHawECv8Dk35heLe+vjGw/eBUC8
4KWVcZsgV1Pwj+xmDQ/gt//YX2V+OIDGmu2QiZnfFrTqbatwThDIzMKrJtMX4TvwVnf7t24Nyyei
Me305u3P2IWV39sPlJcVuKbSE7SWV+8kCqeMGlEvb+W0P4uXo0w6N9rRio9rYW332ROjYV6klVHl
Rk4QDT7mVFsr22WdvqPT9eaD2eBl2hr/DNXQRl2ERncZKz8ja0FwdDRnSBZwyujwENUXLgB8rRen
rNIu5YmZJZmLtPMRYUkOUfKJryRXqh5U+gCv9K24ZlgZWry7CU7bGEFXceUjVIUj1OpI8SC2+uCd
p7Ti6UylY3Z8QSPN9bICBTazmq//g2jq6jMtAkWhQ/YBtDXzUtv3TXHVmrRQP5CmrDi57TCsXEFD
N3iB4HIx9QgGb5sF1gCY8pCK3Tpz1QaVxE31VtjvSKKM5pYKW1I866is+5WDRxP0G0Q6FxsKlta2
xZlBt8x4JjFHrtzp/NZeczLXMD8iGHe8rsiUK4G7G2k1z0eMb41QLEOOK+2T1Zc8BP8b6jHtCSb2
R/EF5Nxkwx55/TgruO+MSv7ld9rgRx7/RdUSSGgwzFgWFrAPsg9uXtFNJ1NTBPTNAGBszY9mGkFi
/KLbJJaVGkDBgvtB4RVTbv2ozNTi8fqbXpvlaC/EqDCVEJX4sWMMUIrCnY3hLwIlj9tiwQ9kDdQZ
g1NQW0MCsq1h1Ob4khVi+v3ERODcVx7q8Km2fNaWINUM58Lyg7m4df0yTuDK2paeCd/GVnUoj4pz
nz88ZB4pgJuAnAE9Y0QQ1YcvoeBfSjUnQxEjIGipqef2M0/0tWHc3LX4DKdvLoDGtBzjNsKY1Shg
fkMrIhMqfay4pWsifj9UM1Z/KGWlEvdJb1rAGgi+dNPkgc7rWStS6ArGFSjxiVYSPrV8ifcrIy9D
G77sDamgd4nmpmIpq7Oi0gBnmR2b1s8/IYPavoMZoWQIkY4dYfTj5gJoNnwYW2eR/woHd8MGy1D4
GqNOWXGpIR3tc/DrLYvmAPkogzCQBNRyFykZ8E4tUKkW6TLKeOBlwJhxcc/IFiJca4SRJMn9PKIe
IYW7DzD4y72A5sX2I7YqRoHVVDapb1QOKcD/cDPlTD35CMIqBo0NF8qlcLpAFWfQVVgmY8iIzQ7P
Uk8Zf/1P4u2R9toKhxuizOYUX3WoIzH9/Hsz7y5H+kg6vdTVlm3Fr5j0TnX0+mND+byn1/NzD67W
BKDGDn1XmcNwDUoZIjYl9LC32FWnpGRV7DxINW9+brlW36RLQYGq2/Yz9wg/TWSu54C9CTWvS1eR
1JJohSrVEt84F7TWZz0xqel3axl7wt1nczQ+1A7ipsBxcI2T2rUwwlS//FLJ+CJFCr4T4wA4VAqy
DL0xv/4JGQje8auTjksUYCrBjUtDHO1SrJiI7IHQd3HTXQGU/OAvYRvQ+hrbBW9o7s/LKfUDk+LW
AucKW2ZIZpQ/1seDGPTD9lczZUjcGNq5Ujio03QPIwkqC4bFptIPxSSKBfjJetcCHEnpSIIQHusg
tbRCru/2bOz7wMayX9QAVCNT+hea4qTq7mpQPYbX9yk+/y1lf7mHpqXnGdQHZJpQMtsbShtMj2+T
Dw4sEu1JQJcijNwqJ0qHijNxicDFiAO0Gg9Wc2hV4we632AO0SQpjzWT7xLPVhhFO/oNQtPINjV6
Ub4yAF/dRFa4uUEd5QD0U+NGw4unsEujokXZKBHsbX+0RIbrnZi8JSxTzuUHY6qv0lGxly8G5CH+
8d/XLTY1ExwRwVXFZStGAyUqvHO6rmCFLkoRk8qpuZ1s7Z9ctgrLW6wPJw9BXCX3wNDpRIhd9pSb
VgoicN5E5SHTti1h6HXhi7eVgOJTy+C4b4Kdv/s368Yl4mAYE1tT76uEU3DTnUgizHZxcVC4MhDc
e6zQQ/1UtrK4W/dfqhcpN2cCHS9jSgGBi+QLH5AdHl2uClS7KGEfruxXjIuHujvJF4YAtqh4UsKM
HUkNbmCneVsxhR70Ak7ZLyVZghORYm47i6vhH1ne6rdsHWruFhN+OJrs+BxWEAnXMRvHOOU/KkaB
F/s0+QK72rnkkuYn5nmfZkyo1ByjlgkbXuPHXi5EOkj/b2a5grA+66ucjf+kQlFDMpfzVqrnpNz1
BH+zJ/LmGqyTnf8FgI9PSuElxFgdR98SuNvDwg9BpFVHY8CgA9AcyAU3TlQRqfE1KXIQuSP1nzSM
2304rVXflKQ/IfoTPheJ9KTPnydCNYQcZJl78vXIqENYFyDdJrU3+X9CNVp+SSsnHnQUXLAJBGYo
srGGdQN6+cuTwsYJZqtCxfjxlckB49AFhp6esKwLw80BngI6NWaG4DYcBbKxnW2uQJjKZvJwLNZP
WvwledF70BiuSphSHmsK5JFeZw1S2pgsiH5UU8VHVAhYjdfXvpHRg3Xz2r830fobut6ICGrZZy3L
GIYXDovEUTJ6RmhionnOQQiebbt46z7mli9HJwC/xIN/RY7SULI5+z49Fj9DQoX7mWPk5lcJU+QQ
35aOAxMFff/hzNKe0HPGYQUNMldBNrJpyTWNdCIhS19nakvLUsbfgS7o1OtyeuKcbi66wj+PxFWt
tJd+r9QkSP+mWyKES/pmTGUEQpeqoOD6a2mEd8TPt2c3cpJwkXY//EOfHQ4No1343WHWAH72btX8
Kz+H/SrPgy+w2/892+/OgVkKunvMRidVVLLxiiSNJjv1iwPAK2SZssEStqxrz3Ah0HrS/Ya5Fs8Z
09YCv0wJvmizFspYl+mNxRwNTCCbTCfVgvMCUiQZ8PScdVqWw3fzSvRX78HJNoYUdx0MAKSNh5VX
LNOJymQ+oYciSbUi1mnff7HA5YHHq+Ipx1MlYA19VpjYB7/qA/qzPtBi9B5rv1hW+wzi1+AXs22c
8i5ikPI1tcEh6lnvQZjttJKaK1vZvHEYACVBvJHsvU6U5dGd+40rZfc5BLnh+lMTul5SSaCT/GXA
SQFYAGUG44nqRAJfmbigByR0O2mFrZUtwPAKtvk+NHNNfxfNF9EH4/Md5H04cbyyvavvapd66uK6
5p1EJBLWE9p/BbcWNERUoccufb5kd6/Mt9wMhYQIdrNIklS3RjEDYBCYWmcO/InzQPiEdlyojl6Z
8dyFP/6d2kzZcF5r8gCjdOD4G++WI3M/AmQt2RzoKSAzcht3RMuu/xhN8grx2Srf6DLkuJ1iITSQ
X2VisW52+RnVP6l6KjIW81XO5brGWAyM3Dj1PKOWNmxTENdjCQM1k3gOFB3SqndhvNO3HT5TYQvN
NTNMUqyWzSnDsIcZK8FUwk4YwgXHQYrq24KBLUj2EGjkOG7WlPcnltcpzv+tIPSOfmoKnoj9MLS1
JNDmqMUYpvJ3nlZknggrgXBJ/hfHmavzhtE2k4/JlMBqyOb7YCEPEm+Xdw84yI+X0wpcBDnmhOYh
w4jiuqDQSFfcHc9nfN6L9EofsRur9kLKCHZQBI+3524YE14kxMHg7Penwj6MbHSZFQHXFyvX1j6U
9xyZmoG8xnsMNY0kn1tq1SCHmqGCpWItngbQf4De/5khe4oCogNFvQwg3vmWCSUxYoeNe8geisJz
rQWywjRJkp8qnd3FW2+Z8LhIed+xftXyzGqY1JbghClTqYoA/torn35kzewOrgHobsTgiIpyc8lp
t/9Ij9cEA7e2JgRl3CquIQ5MxpMU7KATaKSHycdWRtnjkBJ9dSAER2uSKuCDR+FynxAfV2VJpwSs
oVHtWLPyXD6BR3bDyaWDANR6EoVRvPC0HYg1UsTxMed4wCmo8B/uEW0MPJKhPAWUES2Q9FbW231k
dDpyF+Eo/mAsOj+GK49ZB0VXAVdDTotxnLNvYvRxsqY1iZ7S17L+xaxXKH1KJTn37e2xbxhL2FHG
UXaxkjzLsof/na6MZi6BcKJLSqO0+MVXvEzCakLSUjk9pH4CRkDlNi8FDgb9ICt5YTn8CFesoPFC
Hy1jYp45uNaIXAA1GSB2c5K5tZYtCNWf4e3LAERZ6HuWvUhmTSoADjj3Uw1TKDf6TctrzxHIvSl5
V3cufta2GsGBkMVLQEyU3BNevpfEAXS22+LLVxaKfxxdofPw00g6wHh1nnaxXEPPZ+KFxyBkhJWK
fsSt04b++/dNTbRordMhM94H59h6EvcZionSqFHms/OsGyeyx/MNlRlTEJltIj320MYPduIXlMR4
aayHoYb7TlRLHr+/Tp1WQfDS1f076IxVSped9dKl2wVwSN3JgrxPUjYe2v7fsazS/zIgtAaTpDmO
6mrJHIiq1rP64BBsmsviI2D7J0FDkum4Hb/X3cGSz/jBeJgms+0VK5U/P7shohjxk/I/jtOh875u
ktfyxjzyQKVs/r00tth45q/ntGIXdrFgEC6ZHpDLN+TXn6qcSYiCwtsX/nfxP+1Pwmh4b6wGyOT5
o1DZiZjwEzLrw1V/QEEwi0AMneQ6vRIsVZonQe4j2yVZDpEBcyQ9nqGCsUEVxftfFV0jEhbPjtTr
flsCkut88t82GCtW/SffDVKG+HsZTSbtah72IMCCfBGWRoR1tKGqqieKIrzyHzIzxt56Fs3Z09SO
97KCYmObDPBmEhxf0PVkX1pwv0Z4rFW6mmGs+Rol4hSn5o3bbOwPqYbyw0+B5b6S9585VcpEc4uW
y0nmF+iYrbPqSctV/uT84lNk+jtmnhYe832r3jDc3YHEpU0ngvKn2CM1IokydBSN82uYXJBn53RJ
RYEm2/HFJEVPNEJlqyc/w3Ty8MMsXgld51TUMnfuBTS54LbUAKmFX99iGBU8D2L3/xSH3XQKvwwo
C8Ia1ysesBNROWdTCo6PBStQS+yOAXNIj8qV4ToTohi5qk5FISR8eu9gW4ZEjuS4CZeBheJEjR3U
XRXsulCz/bf6c27Bx7iku0CcnH6tQ0uSJ4yxe8DDFt1HIFJgjmVbCloA1VhHzC8Vb/zxnGyzZP0o
SpUSh8d/w0E3cU1CX/V7ydgga9oM6K3t9nfk2HPEqO/5H/NtCwaPD1kkm4OOEkAiOmgGeOKBZCfr
kN/FiNDEFVAYAg+KzSDj10A3NA23SYTjoyQZ4OdRUalVXteMlIq9KIyMo47Hy6POWCPYmMkTZyWI
skTsBXq7PZOnm8KSU5NfDri4QyU2odGvlQZokRogBYRYaJUm4v/k57AlDCJQgLyoV/yvZRZh6qsM
TMSIzIJLdZgTOf2VcbGBdPpFo7m2gw5Qc28Lgfzf1o1nx1HsvoU7DMrhv6MeO+wGkxFr2bmqhagw
HBEnCB6V8xFoYqawIqZWG5JVKQggUeWcMymWbkCUYOdnhd6UG7ME/6gLYhPXWdCR9b+25aAccZE6
Gdl44MhdD9NXmiFAYn6loKvDd0UboRiJi6sFo6vNSuhbvxjl1XP8a9yAr/aMjIve3mZR0RepGYmc
6CYUiRlKy2vjGXKsD9pPpOKkp1fsLmXgox9B+U31xseikUrjKAZzTBQSXP1aIGAMGU5E1INSO8eY
1dmpIJqAPvLdmvml+KzD44HrPtYGcRDG37hitmUYgq7TmF9IxFej9EnQK29ROyN2yk/LknA7CafM
3BXuL4uVx3phrtGq3uo8srYslKhDycrw5qLvbX2mjJui6gOAUNQJC1PuNFdCHRXYbag9r7kTFeVp
cu7/s7anC9MrVmb0+d3Xf5pfhWyLC0lBum3fwAWbBlIhASSGAIs8w7gHCxqttJ5cQq5kai5gjEZ3
z810P0MMWKfJYSZVsbo63ju6Vg0pJO7BIEQzlr9EQE4LjaQoKIhLnLAjKQB/ZqHrFxMtrWlXSqGa
PgYJdNt7ekmFaJNLiOnu7LeckfpHdvEeuIbOlwoJTopgUsSOlZtKv1uYQrmwjb1jAO4+omc+BssS
BffE15a2WQR90ldnjV6gsMXHsZVlATY0rQlbcNPB8ADD4OyHL2/4fcihRgLI/XNwB9a7dDdvaLq3
XJH8rtYliobrWn712rmB/qejxWaIm0ZkbMNR5qX12peP/t6zyNhYHZouhw8LgWaW7Bae2LCTNOtp
d0gb9dWNkAucSs6ks0Rheisp3HYLaTCPCy5AxlgcIKXR1wh/+84woE1SlJtLMJqW2fIFPXomKpAT
jsYa/p+LG2HhZLXNUYnpmubINsYY4VS10il2qOmUvN3gOBV4DuS5+Pv7t864px6T/8CaxRzP75Rj
5FUBtrEeoXnRw7LhsHvQmPOP9thNR6AIto4g4O5RL/lVXwMwXxefuKatXlBDuDzFXHUvvXEAH168
0JW0u6/QzHc+NwpXwu0F0ikQMlIkdUmVcOtG9m1btGcJ43CvDaWznhPgMRo7UjZKLRFc4ikFH2si
AC1J8jOp2gtskX5mBfpa6nA08pZXqlPVBYQUxgYmXhNYDeWMqm99NmX1EgNv/NVdbR7XTdbZHV3Q
ooQJMJPikrzh52EWVhba5OUg4RdnmMR9NyEz1LUm1/XMIWsv7zZi/74SfXz5cpsmfXeRqSc7K0gN
6IamaF1LJq5hLGhxxrDwn5gOMDyzmHPHQ51NddHQrCnnadGS2gjzG8i9xkCnmvCBsfX2UgdMxxwm
a7nV69+B88UgAHSA/BdBDjhqWvM0+EBSzFDpGLtyIgyNGIW0F5WwFCavXQFsqjPqToDpAT/q7QqF
SxmrVanlC1mhRHt8YCSY1eKRZyLY3x0EZio87NQNe/gAGFtYcYMFCNF/X7EdGUYVTMCaNKySZEKR
wag4QhkEnVQZvqPlsqzJsDojqlctQdaHTz637lzTMHHF2bERAgiJPwumx/ntx13EHl6AwTDt+wZE
0OoPjPabCT8n5GhgWIal+wKMU46JxD5C1sIYtM8AoUlHifwRWqYnc6z/Yd3wh2f81Vk+8Hx5IPI3
2z8aPm28MRR/3dTRFsfYbL0ylZaaqSC1OGnT1mWySjP8+4V4+6IjkXjqO0qFnHocZj2YrAz0X+vy
nXUgCV3XzbPGo59UDylOjlc9DvL+pLff5Ytd978pxLEM1lA6cDaB/lxOTF/+FxoNoUToFok6ysuO
IpCLHG9e1nH480hNLkIxkKtwCUeDAlSQe3bzdZ5PLrggBqPQqaZbNIv+NSkA5Ql5V0SkgwQSbzey
hO2gc4ZJGh89IpqXuuDJMqPazcjlDbw2lyeA5sXFC0ZWWxdMc3zXqhlfnJtWtYT6tuSI0fIkFp7T
gecHdjaZZtAIcA4rENE2Hu/WcVZ9j6ZYGke0u1DtJ5CFudx04TpjVGHwP9B0/v1RS8uaTj63YP3c
lE3NRBEtqzLAEbj0P/8otTq0+TABzx/rhQCPZGeg0ALJejQau2Qr6qsKbASgogHPjZNobS5qm1rF
YPtJWqxpJQ2mOPGdazkby4TF9ktWBviCifjWLxD0qCXBvPOHHShpqfnXCGv1YcnZRfz4swQhL9ZU
f/S+Ds4FUzc8kFQPHviAn5dvV0uedb98hyGKQe5jg0T/G/vLs2RX7mtYNGmqCsQ08kAe6QR7qMEv
1yEXRnTmEIC5X3fJbj+0U+rYOjm4wFtsxA9oJJFHSCr5dQq+4BzslWpeFcWKpfI2X56FRj0xiQsg
M3r2pfPOSMt8Z0CTs2BBOzkgTOQe8zjencCdrzBa15pGqFZ3eomE87REMhsK9DNwTEB8h2cgx2yF
ImoOZqdDQHgfX+1UNl9LGl+/gm+wb1yUy6m1+c9UkZijtJYqu1cohKZwLUdSvi506fFlTkv5RSQW
hKHuexUTsdlVYPWeX1Y87yXjO8Vc3yK/M5vejKEvvX4YWuunVlluVrP93eymqR7mex6D+fYZVn2A
KUyagwNZtEiTmM3BsNAZFUhUuTtfVAmgbeXeDS7nNiKMRiVAMyrP2rRDt7dHT6IrHUnDdSbtVsIW
c9+ARIYCMp87J9/Knmebp08DMcokXUHSJKb8MAmOYU7Aj1Qypi9gMDhYTz2o70kEkj3vnLPrsbtn
jXwawBW7d8E6lVqHC9mnmBtwlkFoOl2NajILiUww1JG/eguL8afClV4XOSwAk0M5XOeOeUB0d6O3
T0J7pJowpX4NaYEJ14TgeOBlYuHElABsdm1bRztBDmHtbmIleoCWypJgNh9SZCri4Crx9Hc5WnPd
TtclTZ54ykFbA+3NweiFxipJ45DtzDp+Q3iDSMfV+xO4jTjT8kHJQLnFy45VCyUyC/7kTodOh+JD
mSP681HGH15ZuEyq7DGaUZ3GcZZFHui83mBJtwUGxnPxisZbqqMBKvezfYLgMa05WU7XyBzpjhF8
j98/RfTN3h0NV8Yigcvb9gxe+kKx18gQrnIbVpjKev5QQ8MAP/6Gh3mZJ+g5aLnzQ1cNzAm5bsfs
cHSsCnWSJ/rSqx1blLidvAXX2LB0nGobGyHHIio5QGYEyt6Mkwyfnu6D/FSw7zsElr5hacuNTxoM
1OzLF1zunljEz3mCPFFHdXIJTQa11Zb8DrEHeGp4hCUr9MiTeAaju0yQoeBS2W4lNiS0zCO9GdG8
DyFgLDe3tUNPApeuWtz27cUlCUgW8pzJHdM8AW1ffav/xLBdds5oQ9olBmFp+8MMa1V3I5n+DxXB
0iOrClI6ZMqjWQLotQVsx+vnjB/hRH0zE5qt8YW0M0ROpFSIkjkXbbVZLukyfNBiotOlvBEeLFi3
nIX8LDcyftq9O8mnL0Pzuz6BDCR1GTDdt85BdINcLaf/KGIAOgIYbwsSuifCwDd70yq1grvSL5cO
C/7jOCYmEO1AYFOgB1kr20lvPWRA1MFFxFmxNxj6+bFfwj/sGzL3lpCwGtlJoiciNPR5rSWhgCPZ
6OEaKD7O9YYBZ6xm67oJ5un3rlQFwBrq++O+PMSxvfJ/mn2VmyGh+IrlFjAEXsPyN2iaq/5z39Iv
o48bOVsH5pmwRNkc/NGgDlZv/xIpQG5pW+lnVn6pTHpk2dm0gpwNkrh59gvUVPB38Ilx3nnXy6nL
/AFI9BW+TDT4ccTVz45eDN5so/IslMLCg4hI7SD6DsdL2wUWdrQMvTdEpwJgZ7+XnRIO7heVRIf1
p2/pG7mU1mPDR1WztCrfPj9780UzkcZh2tj+VQvCf/cql0QQ8eC4kcqXv1+wTPlJw0R0rwIJaQii
7P7DhNrh8AgPApq0c30BtLUDpL0sS2qrOOLIHbobaBCz+XR69AkVaM/V4O2R+7CTUr1D7aVgmo3v
a4Y2ENEw2BhnNQFK+wANbGORaf6IiVLXqoG7XMTHj43ChaFHd25o17iMrQMLDAwRui1enR3+pcDy
iOH1u4CrIm1vPErlzP1bSwTYli6jjzm30IvZKZLW+TPQpK0H1EIu63StN+wZquz8BSajdS+93I6R
E+jpzUUI5TLFOXtSk8ZXTln3sMbMAKSFZz/m54rCPCLcvwXAqxPQ05Q4UwKwl+b4HCdkSIT1SZoS
9PUgR3EU7gmf/mNtr9GDPeLnqlBzI9qtABq4BZj3gYGg3fS6HxTqyw/k+NWAA1CLqie/Or94P5Jv
O/UvLAcenTKXj7wTfV6WNks4xQikyIKLyIpp6KL1WnVc6b5S9+l6FMvwKZ9LQaZy0TICun1kEIF1
+QtKB60N5GOkQuJCtBpsgo3TgGJcq4YXpNkHvrUMmzMD6G143XMu5XBqL1M5hW17RN7NW9CAka+g
enSpVOxNblAoIKxOuJ+by6mClOWLUL4M50ECaE2PLaL6NrKLUPurw856OrgJvQ260dGMRADmAJHD
12e6480mRnoLKbBRH9Rn9yhfQuV3ucJX1fYSlHdDlwGgBDcobBF16AuvKnetgdain5biKS0X5i1W
RjAvbhKhvSpvaNl4T2jWhcYJj9r1lU2SV/GPQhItT3ly0R5qfzk497fN5ykNSifUfriW0GxqDxdL
fbyNbmvNZJ4FuMqbF9WsYqVvXvQPjMEULftdsMZFrIkbxzU5SI5EPFH5PS4iT+O+6PyAkvyk4YAc
vcQUuIedEsN/rvjPlotDy3+ImSO+O457daqyVkInfmkral/HmojqsMCAczUqtodDihNUwY4CDl/m
dFvbBbZkQNgkEfTFWPlph2sSsH0KITdyr04wB7kNCrzaqdd/tnGw0iX7+4gWFysuvHQ02wrUxPYV
S3+bVy45rdQs9D53lGGiRQGALNJrxa0eTMW+QB2VVGzsDCtU6M9M/KzBtE9NzQXb9I3af5+2igPE
UYWDZ2+2vEmpoeahlY2UaSCnxXFfoUT5SjaAylkCnlg70CResQxCxBLVDcU5gwiEwX8v2EXJDrg4
9ZLgtJIYGiwZfLM8Xf78u8JtjezBGXtF9YLjx/XpXSKlq3CDDlx11qGYoBwJ1T1yPD8jw6XXnNZr
K5jbNn+SZ69YdDNLlF2R+t7N6QsodBZXCXgbhPOQNIY96PAm0MRvQnx59u6xLxKQ5VSRYxR5E196
y87u53ir+vV2y3hdQmj0byTn6srf5gdB93jaDcd7O7TwF4H8hRKdtFXMKdhy1qlwOZPyRTa1zMoE
uHtM4sML14r6NW+0ktddW24JWxyYDnrbJGSGYzhvoD56upUpDqQYeWludid2xl7eLCUzYh1fLMF/
yVQGQvR+VwPHMCnzY7ZlZ/MjjAd55a7tFDkSZN8JIibFT62yckqsjZM5wafoYEUDnM9x/iKEEXnV
OqcaD0eX7xIvNgmR6UXxZJo2nDjPoOjCNK6/3WwH5AiH9vGAiovKQ67NddhT3GFFO575t4sYx1rO
/noqMs3hMzReO9iWwS/Bldc2Ao606bCvcHyVBl4LgJCjl5FK17I62pTzf3PIlqKhgK7mkiUs27uM
MxJc7pvmT4lrRbYlgV9SBI+JfgXmifRnxptYy0wDhZPqSZO+RnxA76ExR06ekUWJtMiue6PV/SzM
icQh9Pdw300CxjS2Q6xVG25I0+FXSHs0kt1ggIHbUPe32sj0RxrGFZzFWPRPHUkuXCjNPzsi7h4h
tVV7aievFqo4vmt7rQZiHBrLDv9xwUMBiCISEAAiJXjJ9Pzcnp6gF63Zk0xdgcMxdNk35KSizPDQ
3fDSrAnlGMz5UtrsO7bX1DGqGlAWDBQTVq1w0kcC9xyze5GfIrXVEG6G+bF+oKLtPX9qBuj/RSfO
AW34uRO5+T5uitGFuIbcNa6/r6JH8YOg4FjfYMBXAramd3kNA71K4Jm1vewFORGlG5utr9DJBauy
iQQORl2m7gv/zSExQXZa4H1KxPPyC3+FD5iHAT9SGv3ppkQD5V2OQI75YfmqYybngxpHD1OdJlSc
x843YUhzytn5z/er3DQ0rtQx9hljKZAqimM6fcGu6XgAw4pSJkgD+3nmmx04p5IKt7Jr1Cu7Ckp+
8JJMmrc4P4/QPqfxCNiNffdDMNv7Lb9MHUkb1iDZgL+BaXuGevr0slRNZx6uympz+NiexIyL69ll
W37BR29lBZC/3+uL9UrUBhoERqBcNqyUnhCHgUejh4mpo8+hOSYFn1VUpOBeLodGukmmI8CPm2/h
l4a9oMXQweB76KXyYjPRozT+NgcIHxVVnasF+kNpylVwe+cRY5x7Jmhn/wkHMnCuz3cCfuPZM7MQ
3qsxHH+Nf9lXm++tE6IolUF2AunbW6RE13u9tAlTUKVT5kwnA78hjIbMbDyDO5cUCqPRE0o8uRe9
T73CU/uR2D0gxyFObQeJjHL3niGu3rheGs+S4COlLxzxrGKk526fD7PkyjoZceehInVxxeacBmEI
zQeycEjq/9TBzjSGICM3Gh8UeiO5YZykDeLrSzc5+ewpPspanigL2ldki2yJ+iH4b5rG+mDY4Vxw
5La7rNlh2fnS1xZn6tN0Hkc851E5SY7GDvQ7lg+rMEY0ZZ/ILh1W96kYYFFBaktXqs4KeAQJQ5zv
9D6CQeQgJI2WDWcljr4oxoW7QXjXfG3qaKnDXBb92fV+/WGRcQkT76Tfaudf5Pt5ad8tHoQLAG0O
4fDspAdU8u2Ye2SImvIZJMmjWbtT0AB+cUa4dnScI8RUctbJfkLTKExgh9xECrhOgTxIrn4IC54j
6sL58eCZw5bsuxmrIQZMhiAUYVGwkm2SZoxfiDVaw9OTwb6qej/6vdaKD0MGL2kJ71ppzVhf6FgM
Y37E9YhP8rLzSOOjOopomhtgsPFCpvh38V/FNb/x24+TxyjbEU+tKA+qZikmRVcgLzpqXFTh9nGQ
Ltic7Zhaj+YPKrTTARCmeNohbgkstw8kSCpDCIGhnXTfrbYuMgOCt/Iid2+p0hgaARXgeod42sDR
lyI7LSdluii4yRshhGcDe3qpNo29ZWQ5zwI7/NZv7eSldu4qn21kRjk1YERE2XlcmsBbhKLoa3E4
A0pmmcPlvWVadi2/gkjcNI2fpnK0pvT9qbaPMEe2wgekDgtb6nooeAOuK5sIx15X1MxIkq90Lp5E
1hH+agIRnlaHoMLdtjO2j83GxkScBJY6ojT3SbjQQ89UsAeJVXnWBYEzPPU6E3TrcASZpGCQN7Ow
9ISsN3CR0ooaL1HMjFSEvuIs536EFL87lj0KD6rk+Pc0B0Jc6LFpZK6eUPFyOod3pk+QnOphMAXw
l0R2Iiqa4qUsuXF/KL5ma0CUGN6AXsPUVaGdrSQn2+tWLpF8T/xHhZ+EpAZ5E/WVotAAhQCtAwbH
mGDfd8Ks8PMiAeV4jTx2qV7wX5rGv4yqsD1GhLYsqczCXQaIC/8KM8IP84M5nlQEc0hwiYoYBwV1
AUfBzQ7/mtb3enBuas4bepu9bCUr5DKOeZBcyapZC/sNul3xOPzt3W1TiKjKZqv3FcMQTH8Zbr3G
sSV0PL78zCoT43sN2wohD9DG5kR9J1pdglmgfsBgY+q09FWbxggEnMBxl1H0wKJh9bzfJbDoGR0H
D9XS3DgmetO8byk5LlSxuJxy1cH3AiC+229SA3lMmwC1cajBRQn94+TexNbQSCK4QRcY8RCg3M79
5Hu/yyQWJI7qsw36d10RCyVUd2HWGGw0Ch2z9todniy2v9oi3K4TbvJvfl0RgDLOz6yhUEFRKmx9
kmESdpX0znoai5eDJ8i7jaa9SJZDXKSVJpgOanOX//+eSK786MJkL6GDDiU2NB/QWSzjJsvxu13n
W6BFzqgd7kqVTMoukSx4AnEdWTcQWGcbeVHeL2gsrwb+PlgaMJNeOg9Rh26eFP5wUg0dK6jcsXMw
xKd7ZjoxJrn0cCaR5LdercwVByPFyMBg6fsmgWzr0gBx4NwzVlE2Wwg4YOiih+SJsMLUQ06x3UrL
9LF1IWDPYJp+zB2GdOplgt77/8qpbtLhfBQ4IACg/JdpW5Bs9+hSwdjIjjbkk+7ZVpcihgJWeBjC
dBkukNYhlVuzWRFq/34v6A6Hg+ws25W7+Avn/yXbbAjXzNwOwL9RBdCqCOebbcpsChp/UkC7rPeX
7aVXDFaytB9xss48bOWe/gGyJr1vn5gXh3lMC83+Of8yNRLDa4kJsLxoAMQBZsWHbFbDMPPUYa0E
mzgI7rKvNgreH9SJ2ZmbFRF+smB7FvCidYLNUuDxIAxhpGQcMa56fev6BofZhpgJYh0PQSnx7Acx
9JfPzkSs75ZQWsIfG00A4/EFR6oS1Fo9C4fhuolbj80VgI49HnHf7qIOivmbcUE2MATPeVEVT5Uw
PSttu/mkP/n7Mn0KjnfY/jojU+M9dQREOnxj45h/y40Rlk6L0yPlMx1ConI95SPQkzVzotDWoLYT
uW7LL8kYYnPLMpsbzWXgaO0ChiPuvY3aVYiTFBv16jghbPqegRQf7oIQ0LHfjaNAbEx7GpEW+Auy
Rf+mMGtRjkZxsQMQMp2hpWmGpqI310QYs1RRtHkOr+Jq/J6sdTzWwCV92k3PTAaEP/W7IPrVGjFB
Hh7HIgAYmDJn7WUhwSRpXPemXleoPm9ReQvhDzVsiGyXbmVUuJtEKqSboyi9atG6O8SIiAY1wwxf
SlZk6SU8rWBzqZm02HcoOWIBVsFohlU9awsYKvsdepY4Io5Vc15tikmU4EgET/8J5S1zysffV5kB
ku+NOxudnkNPFpMpM9EtN8ct/2hO6gwGT7Z3eIlna1pPalCX6MMXYo7Rb94iHANAfRT2Id7T4yHg
zRnu2mMr+SeiComGsbM+Adm4hOk5D+BvDgLwgZLEOLl/iNg1w9DbsPM++W5WsLwFLimAoCvUwBWN
Ag1QtTx30JG1n7Nt9a53bLhaVCkO2OkFP+i1MEHmjpQ8O1JxgdN3rcXU5DbhC4h2150xiBEW2OMA
7L5fzcX5b8fJEk6G9S/9FV9Upul+0iMCSqZMeBBqaL/4W9n9Jfu75hnqaLqWIJ9truu8rnjLu2+i
T/GVKmkxW9ruaJBQ4KqnJIj+Auh9uWJh2ORS6BkZv4gFsAs0tA0G+FL83BLAmjoq2YFmLVEW9FD1
EkjdY+m64UTp5ztTcvTSYwxqKvP/CqqwWR0ir2vdj+HjghkuwkaWBeOJ+N6WUiOBpwzwh20xKuts
IPWvAYs9z+YGxq3hAz7siIZyiTVsHo3MO1UEEZPXqFx2NVjW27KNpDAUs9y2sJHXqQSwe49Ofe2/
z5DaV9zbO1PsT/bAdu+u59Im76+yGxcxwmMhOzptn9b2J2b1X/k/tvgSIKDtIfVT59qtKGYtbwRn
Mh3nm6nCIE0aBKSCaMZSCYkFXs64/G7AR6WGaJ16N2eUySX7oryx/t1Tsh1IOpnoEr+Ch+qiV4oL
WS4jtkvO+Rngqg3moL8t5PqexedYvuvdLtVVi0J5g2eGgNMr/tWdvlesYGU27wnEEf5lVAS99CiM
CVhYZcji0R5+nWb2bozuIg5ht65l3ZkhqWDZiQAaSl8xnGRE5kDJ7LTNn6wtaiCCFX2TYqv1AabG
IXdFcigOyCGeT/VzKSRD8R5/W2LamBn0h1uYOo4yklqPh4pwQ7LFQUT/6VtiA+32i4QyIjgrHNQz
IVB5w2365SfhQlX+bVd38qMLk0USgvsf+ftGYg8QCcAyE6qxrozCo1fAKpF0wyXkrsZrTWcKo4aS
A1Bb31xvQVSEFnNUn80HBpkigiHii1WJ7bCqv7yPJ5/niBWV3/X02uhO+nD/5o8e/etD1ZbJL03b
4gz6Rb2p9U9rL2VNSLtB9+FAcB31gg0cphR69QNSN/v/69UKfGCVaxE4WOrVqTH7E/n8YPUsl0gM
pxfp200d3oZ+yps9QE7vVVpHCkj0SVKFUMoaRodKEEVVzsVq8ojdE+yfEzG0DB3NmlBEPp8Rj4bM
OfceCSG3gmK5PFNJPFZdecOIf3MMaREZC6JPzvrN9+kQJ2626IRzj7Gt03KN2iksLEjfmcFaxPaJ
dP3j4yP8htwN1Wz05rbFgakK7dFbbGIT3T6dmk2TTB5+Gs3m5lLaDRAv8ypS3gwCJBa2e+CDDj1m
2Gk8oUdbxEbeomlAAWh8BWYt7RGqKepd9hzthBbLzkktfA08APlx/W6X0oR7y5NvQ8EoFBG8u8zd
rQVBq+2itO6ioV8pDgAi9rcaLjEXPMnpQ3HUjM98YkQJqU1XDUDLpKFFf5caFr7qyr5zS47MBxj0
AjUg2N5m0MKNSZt9EVCFV7NGP7xlSD6m0XxuexUszz2Ek3U8jroKHR6UnLiLh5hNTdqLbd7kNoq8
8LJ4Ewi1XM7HroJ7NSUR9CDatZRpkAOStrtAt9QCXz6vG2VVN1Zo7+Hi6seRs0WECvJaUuV1iVVz
9LGZYzQgPyHnXPQOJKUnAN4o9d0J67Jy1wepRsSEQ1qjGahbhvnYzjM4uJSFPGkBfVrRLwNhFcAF
HSYZlFEXAJad4YV+RrDfVCsjf6PtcsO4NO7fp0pqKo1k4TeNQZW4GKxxd0ttZ8jCJQ313E2m3AKK
upE0gWb8X8fkkuVakCReeHjU6qmfodzLYxfdgGuLFmz0rle7jzHK4QkpcZSMF4jiIsEhZrBkdxNc
rhR78jX/z2Qb8CS8IuqDyeNxj4u3M/OADHpgzMx5ZigIJHxjjLU6EbKF9lfIFFpqB6XxpWpI97T2
eqAwjdi9Yr6LALW/HXL7TGx7Gf9mHtM1W/NZUxQaAUxPdL3gobW/W29p80xl3z2V/3wkbnVNwmTc
VDfPqqj8LO4MRVfGWuD5oQUgacdV4oUl06pgAqy8qwcryTuTKb2JVTSxF7uyJk7SBu9J+km1E9mJ
mTRZTFmvAGu3A8ws+Nbi1j7Ka7lsEDmWqQa7dgU1gVJMpZzJG1W+XTmUKG3HrETDJ19GKoVgMACF
nIE3hlCiHfVGIioLgkZIASbKCzE/1jHdXvq0aOpCZ0X+T9EXM8B5w/A+5cOtzie1D/XjrdmhgjyF
lN4QB+OrzLeso/IETtJFVR0ECaX5vQW3yJu2VXYM8sR/5gAS5UcqEjfiEI3heMz6Wxt3XrPsgL3b
OXtlniYqib/Xbr0xes3H4JqpENHYK4Jsj3zRg2yDHK3r5Zx0TkMr18CwBIu16nj4018qs8i9TWQF
nk9TFe/F+tgTr3tjrB15YACfhq9TD8K42lLAr8F3wdvg9Wln1gOqnpZEBBVP+mCLbIEiumZfnSUi
Q1ze4dkcUtr3af+IbHDcpufHFljfnbD/4/yzOSWH7tcEhx2wyW/sLhnL84aWfEJsLj11oIpMyA4U
79OK2JNDqPSVNi99oVz1z6g6PBsZOuqshYnAI4z/Y7gtVh4CJhyGDm8ABt59uV+VScPbuGmMGNdZ
ugPiRUOIGURYUMT6xc1jotIz3nnsPDQrCAAxvLoxKuXo7vUhbKvBldbZr4bGxKFePup98Tf/ju+v
A08Kzwoba3Png4FnlMInPpcNM0NjQe1VTouqPRmYCoJfOLB5Ky4S0SSb4xtm0k6bX42QHKzn2XJh
3C53cRqINEP3lQ5Qj5Nvqt3rmxGHTS5U1p7XpiSmWN64eHDNYJQSTBsQQz2/t7hPHvpkvFSwAgRr
JIKwrn6xhWP+/8kK70TrSaRoyrFjp1YBd6/1Dp1BJYOHkD+f32DRTxy/d2dRjYoBt2IdQs0ZXFh0
1ZypU7w2hiu0L2XJjpQX6KFjQwcP9TDpsQ15lbJ1kZDWHEwyrAA64wS6keX6ma/jAvlvt4EKKDSf
8QLz9Uo1UGGGlkPATKNgyJ0Lz8JNKgrFDmy2Pll8bYDyBoWwJ41WG16LVxq4NZUW8CWe53ySIbln
3HAjlGbx0fT4lPWkUnRKWLkuom/APbKN4RnXR05oj52pOeUSdbY7yE+sSzc/3+Ih0CdymwyD7tnE
tu3lMHJbiHx/NJcE6JXRuDJvOd3IIuBKxS0TnhtS2PI0dS5P0SA+q3RiBCRFFolqUuU1QSTsherA
QWtjTa52k0Xp5fs2cdib+lII8yWFVEzgwv6JQkfagNCfhTbHmJp1BM6LBpZT7Qn/0KzPK+svb7ST
8C8vlQ8pBLkM2l0hHAdO9mL9VUs9myQ4BfrtM2PS6UI7Zr49uP/fzayxnfyuwz7CdGGmYdS5Sc+2
kYd+nC1bXj+L5ke3jzhKdcNMH25Bsu2pGRZk8bhFAsK6n3PBXs5lKyciaO/Th3UXXJCIFVsQc1FC
g9rtmC0zn+JAikbAKYSexoj0sdy48o9QiKbyIeqO58l2zo3ro1MV4o9F0Xr2+pTmxsGuCqUDdtp0
M+N3O9Gx9+WqeNZm1axTRwn+gvwrkBzx6iAKoeyvMNjbXa3yikUFdXbFmGu0X/OSW4atRz3W/etn
BP2qZNwAP30isl1bE1inLmiFcyh58EMg9mgtmGm9zoe6X9WFLXPwxs7hb5figQC63PNvqqAvHca9
FdTeLAPGpGNK3U3aoLDCvQXj+tOf2H9rntQhwMIFLAC7EpD2qjj1qvNu6iy5QWOqyaD0b/SeURN3
vaa9h4WqeuYt4lQgAk/X+fV9M8M2CBb8i9E5Vb1YzDOMRPfjrSwNGWFOr5787GdYbLPnJcxDIW5z
isDbwdOiHssL9O/u8lFwkmxKWeEdcEJzgGkTnacZ/0B/DXkobz9QddT8j4JyRpWKS8Ugfz0HEzEC
3Z14qmhYp2oGnWQIEa3XnorTsuHfLzzNFtTSKQT/HO+0YtqUs4bHTcBHMFbOosS/UJBeWyLU/Tl7
gMKwIGcu12zMSkBATMX9krf/gtwcsv60k/amX8xFwdB33LH8BQEBAxgMR+dExUfQ7rc2libnR4Gk
1TwsCY+Q9TJQj3ZluF1xhQnxXWuRUkT9Kk1kiACcmNc+qH3uzcIT2lO0z8dHBk/PxWZn91xxUnAT
Og+hrblgNZOpj9EWiHh6pgTop7rNPijJicIgyQk4fISyL58Wa2102ohxvcXqYNQ7GdFhFyvxvKRR
pRWCX3pxZM1Wy+5PFvLLWqGtIGtUgNW7B3Y/ly69qNGbmq452jIMk9YfZXP1xa/i0an9ZwpSz0hF
AbyktWT8UkxBfjOtAU8PHZXV3HnEeobdFNDeAEY+atnOsT1UDLTnZ/L0HgJ6tMhEuiXS0Zq1B0tF
kCLCWegrPKhLLo0p33+KbqEqcCx/V5lfhGLOB/ll71gBoRCqsKHKmQl/VvaLSCQ5PxCm5Ne+cglU
MnD8Ks0J3tPaBXAHpSMPg9/rKzt43SIdVPAqWMeP3vhCfltux8wEG56eHhyOeFyT8szfV/ZAOpBS
P7g+INuNzjhNxSrLk/2FLvzC/DV99jR358Q0ZnP8t97PXn79250bi92gfMPkfiql93JujAicxKhh
LhFTitvuDX1hbpWeqSimOiKsF+qsPJ2IsCkDVFdR6jxhuMS/Pbm/KyPCgN0BBnFL1Etr5SjCQE0Y
rECUNTUF8cJFsnc9sf9/Kw+iJlrMhMWjlrfQQ9TbyPhxaxgZJAKyDxBc0TPRJh2ke4WlNbiSN3Vk
9l/rMpE6ugQAWqaww69XE+++WKWsH6ew0Am5W4U2/LVXZ9z/6p2sVEZvWKEtXFCUkiqDMtFBw0xA
tJreTICQmVz4czBMwAFanhecQlVfU/J2ZH8tEtNecZzeheascaB7RlfH9a8gEqnQkm0fIcB8XKdx
qin0+aWtFQfVA+W7+Z9jyOKPWw2BVpUPqflsNTls2w2GcbLUjcTR9hhnw/W+kViJL1AHgEYj69Y7
nMgqqjtbEcuvWf4ReMCVcCdGVhkfcNXpdqOfF/XoB4n6PwdeMqWWO+YYIei8P6eCD0DfFGlSrlNZ
eFVRZm94jEq0gezD1+QycjMa9MkhXs0j0/rv6g/oM3RAsGIPWTvKly1qSNsfCyAeQrn9a/e0dMw5
bRg6XKQCqBR3cnbT5oC0Y6gBsePfLfeNfkZg4dA/mjmVbRR26YzNcK+K+LSq1M49yVjHs4CWsZpw
KZkM6Sdt/rEm+Xorfa3wlN8bDxO5DsWLbUAbuNnBLKqKVDqeBiVuN5AckcLQcyBLrsOhxkNudxAE
CD0LQ8LOVSp2FgIRZMhQeyYmcrOJSdT18VwlYDtrqMDMwTTVP5DVKcWY+onwTdUHss0zxgutkrFd
//JLU3mYodR7E/nd/G5knbW/3k34oYvq+1iFwpf68O30ogQDrq2KhtCghzOWFB3KgEghjcKbSdTE
Ph8JNqiT4G/6/H3H0wWe6BnyyoCi7w0SFHfVlH9ArCBA2fiS5gZ8cQJm1FZgGkbMs2H93H5c+SQC
emUHaWrCFwzsRs+Ho0nTzX15dCsMXh6cOe6bSgnTs8uEIUc9biIozc/ImsGfcOG6G9zRGfPtaMto
Xc1SDT10lYk6neK76IWT09Bahfx25ZV6isVcoFdTjtk1Kb8U2YAsCbYf3E26GPggiXe2LWNplv0A
OCAaqFOqCfljP6LFXyyEk+LAmfCuwx/C5kPfbUGC5GvMwyDYKFq2iwdtlRW6tMBS8cNRmIaSxVqr
JYKxTtOSWpqMFIEnV9xgtrYsXrd3bK5A1F4rMorj9WpxWmaK/3VL/WR6ybuEp2ZGpJpAZ03Sz8tc
pd7gpH5kdA5QX0EAbdFD2Z4bUuzFgTjzN8VuVmFJBgXyGYei2QF7vtPVRl12yCcTtzltrzlasq6X
C5K/LQdzl3mpFU70sV58ybPDDIGwt23pGBgdg5oWxEXqHDBHiqHkrKPqwVXDEt4+M0sdCZsqJ4i3
ElyXU2yu0afR4x6MMan4+gQIvoucCOrP5AYb6Ix2RcE+1n0V6PkqmLdbK8UX40vdhqiFEy+S9xNh
SsgoiDJh+4oIfODWrogDTaVa2sQ6ZkC2JtyWVgMTZHkDk1Etmq3tguJNnY111KQUbTxaZUyBI7JB
AWwzRUAwKQZIiKVi/ZJ2skVZbUjIaZPmlReKTVOvZGPrY5qExgrLPIvPMQ/jBdYih6bjhXCEGov5
Ryfiase4QPzqJpJI8cLfz0q4nQnhp0R7ffe/2RasgfdlsbP1VqGCGsE4jchJH/olH/LeV/iG4hSb
IaTNf5OAlq0UNffeX0onJR5XcPlr9m8e1+Kl7tBlMzSToQzDFIVOw7W8ZkvNbp5w4Zy8jmFbCKk0
oO/DO0cMmeZ2EEsEmC+8j6d0FWRNE2fnKZt0JfmAWs4jmtTJHpx1dBEdmbkArhwHEg4tyoPxWtGs
GG/pPS0yjQ7mluPZnrc2hYA8xA5JeXcmDcl1y8oZEPWtKZLmxq4+MiCiHxFjI1b/FJfI1WxKYGtE
IZ0eO3rbgGUKnvbTY+0PF6RHbFxPjezNIkQcuGN5JouVMnqr4SLVGTrS2IgthjZ/oUCDGe+MIaeI
ufWAx+pEYFyDXOp3tbYbSsn83DnJd2GoY1csxotYw0Hfpy+mk+WUWGFIrbwdNX4YP8DW24T4fhc3
M6RSniUNUXa0DJfgy02Sq1WiYJPMu1Xp0Cg/m1aUahNu20U21wGUupZ2W8NU2eNcJAOiz6DibnrA
f8L6ZR4KjwN6A0Jck+713KT12QNf3H9/2UgMaZVMv6y8E4Og3BRy6kv9Qf2ztp7Haz1c9O5u2z3T
muXL2bVoXLdYqqNVx057XfBJ3fi2FK8UU+uJnlsFBMApPwgoS0AwW+vFgLgBZpAmyDEXSXsPZ/UA
lWwElIoISitsB0oPt8aiFyDwFRuqPVA6/SbKC35SHuEyLJ1AXNHvCRsHjvxnrpj0wGDH2fD1Rf6S
uSgqUgMjHTR0bJ7hpRgYOVxzGk2sWuYzbuhsa/lkTqlLty1SA0GXCVec40Ban4M7sUNT62e2Zlwx
7dm+M1DXs7D3BTADVBXuhLwKN9L3a/NvU5/PSGay5B6cogG1Nm5ud8w5qNDZDDpAVElWCIn5woAq
/L2ThJD/CkLolUaAjnn9I/J8o21742nKMxPwp9f7yqKx4LfrIfYZaKxSL1AiDsfWVARpjTdga5Z+
4Xafea/cMZQWYMHufPZGJyINUVMwv99T68CWaBgiD5iQzZSaNxIrfcLo8tFPD2NzhEjwSjfegMz6
bF+4ZU+ZTX9huPKWRiaUePs4amH2hJN0uwpqoPKFlxNlF4JCCP7+rfd4NKXxcdHAwXoy9oxfl+AJ
FPwQ7pgZwVdsIsLj8MF5OAJT29B1e4SKS+kmgPeclmtTzv2htH94ufntHLAEvvPHMTiXCsFzPqS8
tOGR3ShMFFBVmgbChNCXaqBkkdGI8ppWpQj3rak06OwAyqXnBkv9Ipl3TiX1oZCivhicGlm6I+IP
14oSByvC4lEO0R5XEUoCm3hYu/8AfwMVFg3XBwkD7eVz9ahttvnnzeZUuozGJHMGPME7IJoELx9J
spffxxMsN5sUNuCSIVzaUi9tD1R3Ll4dXKylkEctDxZO1M2NQFram4rBWpZuqeMy+q48+frquRUW
DYtK7w1g/031za/Pl2UCZqbtWCx3e95OP3LNITDtnUmJndfye8YBi5A5Ffu/VIGUu0WreXpVbR0M
mKcf5jQHJEGcvgCwuG5+c9cFU8DyjKlept8OrnkCIo99Jv042E/x045VxHfm1iBRUdZupJI1n8ej
1V05UZgLH3YM1qiXiVD77uZwxAaxkMWO9HjZpVestLz5BagPeFCnImmbq4RbuKpz4oKuSXoU5UeK
vEyE37X9CbuOt0QS14bRggC2qtG6VGYSIwzTj5+FFpOKcCLyey9QpOoeOKszGl6zTQ/RRWS8lC74
dTSBgN1jz/v+lK4IcU+27ruHQsUPAYgrw2me+tqOdq5ZWNw2O+UZXGoojLf/b4rwY6egT+Fb4dba
eVtnQxdvW7jSwmYdYxgfgUb0WECqvbliTj5YbwbF9pJCq31RZ7KSBaPpHXQnt9jMf3x46bAZbu7X
jYdFr2SEE+oM+coIwiHxrtlWAXuwUZbZnQnnmTm3iEJJaQDzJVY/55Zy72LIoDplS73l5oY4CpGv
ecKFBKoLW9tBmT1QhaFUbNFsTKHbw540CVbFCwhqsFwZ5wroRvc3LbQh/mWkOR67FLTU0UDfVExX
W5VBiCns1ejpLQ1qR8AT64y/Q6arZ4s8X7Z5cMEBa+x2p9p+tEu6xTNdUk/duvq37rOYQRm70vwP
CZUxJ0taw2AX4THGfQ4mo9PKVOpYQJoxYD0ZO6pZBmZkiTuEwD8kT14YCf8rnFhDIB1+VfBk4+yz
hhwUWhXDFYL08fLQ7tG+Q+XM56Vdi44ZmKtMBFGcLlq4hNeLRbuORb9oUXFSLE9iJM6DnFaxG7y1
zFgymzoHVv3njXoyeaBmInRD+X/RSlGlloABC69u+Mre8ugGReJ/UiB59T0Q7Y1i2yNmsZpXpBHB
GWooDo6l5TKmQMbk5keylbUhyYJyLbaLIIhc/pfwg56npQQbQQmXNAqW2vIqmmxjNhhY1er6kz2t
p+Y51MvRyJjrxnuZaD+qbfdS3ZTgN9R/WGVsz9Thn35vQWWk4TClzmm8eMbeMU6wFw6PY06XetvC
GAqAmOnDceYgjylCMsPTqIyGRUVIWh5/pFcJ31WxtdW86VTI0ayCnt5NbeJHxvxYbMpicBa4Rubs
HgylUZHq8i8EoD1u3VZN9o/xB/RtGPg3BVjYXByql+NOFpJUJ+1Cc8vWHg7etPlYj6/iin6vUK0b
lA7UQkTlMtAhUOFbdITSwmnsKHNNKXDIs3C91KUV5Ehr20LlFDtfpRwc5FH1ven03IXXZVDKslZ9
ILCcfohFkElKnwklLcTJzep+6CMpNAavGQpQQSRJBV81xbtPNCA9h2pSIlh9KoHm4clhrvLfY9Jr
i/fivvmAVvX+d9KKLCJZGUphwuezs+TRaqEQbAwykLYrs4PK0vS+hf8Mvt1hgBb/7xfQvyrs+jRF
mkSqWQYeTWrNTavZ5DfZg/L2GMFyJYb6HRlqHndk7eYprSrOb+vJWKRIENSgcbHDVWgJpRHcGdTZ
myCkTsGmpBusEWPQRalJopjPfhoqvCB2wSBsk0R6Pr8+QiWCJqaurcr7RayniIiGeLOQkp0gAsGe
2ZVcGO02VayvMJFtstNulqshAlFFQjJZBSiHhBo3Ws3bal8YsyC3DzGclJ/ixx5knFK29is6LXN+
SmDeZYWJSwQjz+g45Sl02Kojv2MVU4tg4CNOyLAoa+WH21FqqeLcAx3WmSwOuW/o+GsLBJOgRSHA
PiYzF1I9KWUl9FAshiMsFLAqCGTYIECUlSURYtVR/RRlbPCv5rXKHt3Vjyv9AwNQjyVy7CQNIpMe
ZV9nLeZ2fYonlTS/7buGUlWHiwnMz2E83zz5hF9NuQNELdk54e9S7LngQjgRjiccMITGDvphRG+j
GYeQGAcPCCppWCqLxXllgOYRBIk6i4ZZjCLgYubvyvXPNu0VtMyGh9t1qXPbeV2tfa/px5JuWTSx
YGAai0ecjzdeg4oMum+VTiqNNKDVehUlwolxQZu8bmQg7877/ThnIF0VXBIpdwAQVfRXUsF3FcFk
dTqKLimfd4xcdK/kBF/n7XWDqZjmH8B8kDE8TcP2tN+MZPhnpLh+/bpL2jO3/2HM5LOqWzkuvq0O
enJe2siJknd0lVlW6QDO19w9/thS3XMoubO4j75hLvpB2CM7WaQXSdAKKrlwC2wQ9lVfOc2NrzUh
h9fiypRzRAhjOJn5A5m1MKfwLMgFDx7krhDYoxfEbMrdC2mhqURPGJgJ95D9PYMJ7NsODCDl1tkC
8rtt5qkrlBv67NG3avkdRtU4O95opMRndmGAck1Q5r80JVwE8sgEI7KDjwVyDjwi8vIo9Agb73Ph
wfVovNnL+MZxPQOwpB0ofCj1zHKH0ombVmpe3lfmwOIGIgzpTZYsWUCNya+WVwGAsTZCOfS/57Qi
7jhR1ZFw6cVxjvSiyMTw3VfuVw16ORzI58z6SklDOwWX6oCPwnNcf/sLyRU4MP+6OUQxCpX8BK9V
yil/QSQdYcQpz/DSkWdGOBLJDQdmKxECIzx7JmlrjU8yjsuf3p+GV/Df953ji65JcqLAAxGR3xh8
XwsMi1/I56GJjPgXwkIDC8yy4G4MBBkgEZlBIEaUqF8jXumMVlXnPZOPg3SBExBGsxcm5Fi9Q6pu
mHXewvi0IxXeHqrnGt/wcGCOqna0FE7tYfwbIh/oexT460mA7eR5EkjSFIQQscY17okd+CAM01yE
cgOr9iSxyU23sUADnUYYJVY480ndenPwAxw8VavHfT4jGTPz37buppyO2kGd640GrrtR6OGIg5pl
E6kAD9IpXbWBGgEvVpQTEogqOJaYI24dYOm2lZiBbOA6byELMrOIBs05Ki82OzP49dfsxf+xVwCE
kMa+v1/TfunwwsZWUqjcRXsIOtsK90a3XHGavZ7ny1P5sHBMDu8YWmf5PefkFcj9N6vVD72gO6u5
vIbLuze5XjZ4Be33civoWh2DcHaJZL/HyU7fxdNpLVvEROzoQT5faQAod22O+qK0kNFjEiyX6kZO
1ru9RL+Lob1gCnc8at8XA9figOfuOpwbrCVGOLcxResGPtZCURfbtoy6W0PEM8SGpi0GtrIfaNVI
ZQ2UXg9NF4c6vvJXCme3AlQEn+q+nMS1Zm1te7sCdLZajTXCounzHo7ZUr1X+Wq6DtBIOmWcIr90
+CDclXELQCEDF3VzwTGbo9MHAjEJslxJdOg4Dc7go84f9P9PHogqan5I+RsIN5PdcYRjtTB/oS/s
PguGuEaOaLr1NLvrI7+MjR5i1w/f8Sdp/8ESPKOnoZ8FRAY6htEPd3b3KjXLopYOPDq8t/K2LcKs
F/rsvqUA8oDsytL9/c06LrVuHcNvNBGb6UvkyGK5Y7usBzDYroZxk29RF5oHoPsfGR+FxHR6KMJk
KhDsrcFqHMesB2ahndFNhrMEcRaU8NcZwIo3CbV+6npEdBSb4KXJkPADQnePR7FC+JStt/7z5Xzm
6uvebQQXs/TDKMxPT7MxUm7ktycXXQ24fWIz0jNuMbXgjDQXcDufL2HGb7o0z8ixwwzrJljEWEtL
0YSlHQSix2HpAuo6J3Lu/ouoblbYw8NRdFnOrJt7HwOXV5vxc1OhhB/xxqY1HxzHA+IXWHV5bUtR
s7RtE/VbQ/4py8OuGdNuy7IiBrXVTOVbaXe4ziUHvHeWszdrHokY+K3v55kBaTf5JM4xk1YFf2X6
oy47JsadO11xfFv0+yS/CXXiKOMUcOuv3KSE4hLJYWjzK5tjXlDO9EaENuWBpfnwPcICLJtUZdaH
TVt0nyLTv28EKC4lxoRwdRFfh2/W01Cz1zY6bZgcm5BuEv2tU5645f//WQPOptxJtMyOC+7bG4s+
v+WEES+NFOUqUdnOCLyxfQTv9QqGFqb2xNza3N8js9I21CMI64LVGVAbYuNM1pJ2pi0cmds33qVM
WYXRxdYyesbEZrJo+fZEgmtfIkx+kDzuauDQ5N2r+llT8BAJjr9juqBfxxWZMSa6Q2YRwpW54EIT
QDw7tjtKQvHxWu6gL9zXxre2MvBv2t9kLeG1kno4Yxg5wQoCDln6lCRLmuGZTz68W8jir3npf/Kb
dCtmyDapBumam/ZhIeb85+gsVv0e5M2cFQs1YeJ7ULY8qPE4+W1ReZOK/okJ+hjhcEDcxczkINa/
MDu6IQ0xd5KlMohp62jeCpodizvOJZwK0Sk1mjyG7kgiE2DC4SIlWjuGsc/KE5fx6o+zNosq/qfO
WWDUEHMLsIUapdnuFsMQDX5nmNe0TSzJZkj7DlT3ub9+hHXP5TSIQSyBrJV4MNcMGNJf4pQ6sYxz
ASX9ZVtbpajNYxPGqgNxGbg9C5IlbhocUnR5Upb3VfK/LVRglReuLmrhNrp/SrSujhwrLxZx5YqX
XnAKkk8nmLONU0jkhksGh2s3yZIDzDac9M2L7J79FbWGQmOtP72/OGJ938x1aMeor3ux+nbiSR91
LBZFTv3eOB85QhHgjVGSezGrJmcKD4gTFqEz7q+XxFMMF0rBPShl4/9v5iA5zwciqZ6PaFAfLnoX
sYA46o3Fl4QBY2oYz0N7ubkXfl5tYwCL5ufnIVtfCVxdJTLUPb2mr0rEjR+kQBndqhFVRdyjwhD0
9xVNcjUWxEiSwdave/YXkX21P82pK7hyMj0NdlkeaoZULA7MEjlsV2XMDTYShIB4s76tLh/HUUD3
57qJ1zbv0Yp99Y5LVsKv7uG3NZpRgOgCuSEBbfrlQigqXPe6qQshQWFzcjDbY1gnXKJQGITmUB5W
gKhvLvixFyCwMMYJBY84Z1hdOgaga6mXZHFlgH1IZwETo4H+RcbFbrPZJWJwvzqcRM7vwW006ZeG
zNEoD4F0aMsfu8c0iru3CU4WiSUcxSy5mjzHIWlz69E11EUTQcxEeDBC1IojSqG+TZhGzFqmyZJS
FKL8I7wQUtvDPUF/jG5Xr/foQUR0+SQROK0VCUaNrQQlhncc39FJ/v+gaV24IpEDPrCz2KJzzUkg
Y6lsizI2YjZHQtpUq3QaRSUZE8AAf6ekfBViduhhkOg+yK2bq/UbAbLvQ8+o2oRFZIJf3DB9Sr7D
RtTqUoOV/Y5CaXUR0xWaoKJFj7TA3IvqY0O+VtXQbtlTDR1EOEKNW+ChThdrbSelJd5f/DvCEORM
iVHUr1kvDeAzlnImuF3r2cNGVPiyLnroU482uL+rY++YLmS0x6cj6NMwHjWa7LPr54iD09QwyFTn
DyKoxsUuXVJT26IQ5TTG1G/P8l61KUY3nwDIshqe9GQgxkCu6GJ5mVbqSN+0EE7/z8cMSb24ZHZA
b8vfnepNjHV4SpkrVrt22XJF1PuqP52KsedwttpUd8CcE1WD/GmytwQ6Qu08xaOWHVs1cKHZcA8D
XHmbhFSu2OQzcAAiayIPEr+zx7hUhkDA5CJnjceQhckX104kg4wMup9BRtP8YqD9eN/Jhl3TvTqN
gZ09NOQY/n+SSDWx/PNgOT0POspN0d8VWsFPzCPuP+BdSyzZBHhzPdgxqsNoGsUi3+NbodG8/4D/
q+Q9gHiORLexpke+CUhLsE2bcj6d4cyMkLO0eNwNRy1BuD2YyAJXvVOHzUpbjeGcT1j9Kobodkg4
30ZG418PSwUTy3GRWF9vet3drQsjONFrGoLdisonxlSpqV2pgNv7VnW7cbOej6EwcMOJNvTR5SUv
U4wsLvb840DVRyA4zkyNrzhIaIXIUtm3gHAw0hvyuOa9dHHQRvnVkMgfsnLwYOYUNHDRPCWWFPdu
47TpW0fnZCu8ob1IoF9V1fAFb1y/fJTrIBVUWXcEUHCfVZnnwnSWbHbBqinK+UMcSWY4LWuxnKGV
GkS/ofw4NEzFhxC0yKVI0adEEzd2PfiqsyoBQt4XNTbdn83UVkajwwPIMI/AYQw2gl+ie6NGgjOt
IcYfMsl8yWk1epc/YkzKu/73m/YNm0P/14H44OKERLT+VE/Lq0PttrHrZUSvZn25BCqgYUetyp1w
7mBdhclqzQ0z4fXrSW3CiTAuUCka7VCmmpELDoSC5KyWHi5efzayOMBlv3eFfRdwnSb4QjRVf3Gc
PQmfJbTNERNChukESseE3TVUoPZAWSwIXQQ/Pqx4pFtT4fABI/2Jm3KcPxWlXtxipzHLnb4i3fwB
CkwtkPvpJb+v/KDuO/BL8NQejwZcgybqyubeFexYjAVyOCGD0nB2SsldigGRKm0nXKPc17PKVa+H
oRWognnFOKp/VDR9pFyv9tGXzAbTW8ev6AxOGl/cw1QiaBwSG7d+66T2uNlq7Q6PhKwtmLsDE7T0
VXsyeEFoiYRdBPv1bkmZJsg6SYOs+VDF0+PABr2t7ENg+lPWurBBewDm6QAq0W4y5PqdWi6pdm6F
+a89e0mxG36g76ri4nkErEx3Jf5gzqWTL/PW3fCVSCsxYaSla1YcW6KQcuujgxkCw0eRIBmxCoL2
vYFB5q2/od6ZaLA6JkPldar+geRK/yZBwu7p/+X0Kaj3emEVleyzUWTqw+p1RguIk583jDxgNs+w
4aa5VrtZ4dAy1uDot+jJjxbMfsN1qBMsJfLAaPj9x59kpiZjzWmDsrgCz9m/CmUjFJnQovHdBPMn
03vAtPfAj474DRY/JAkCJnynXagSdWZNjObKTh5BVRhWOyJBl7Oo+u0vcvQZJX7JExnxiL+S9aae
OAnpw65NORARUaJiI9enOILyN/LLGHgj89PHHdw6XjatbGhMcXoX0iSOjSfyR01S2+YASCSopCE9
PaFdyJPZT8HArn59ZJm8+Yurfl8l9jKJ6XOX19ESYGNvLFvAaK/lhJ4t3DL3sCRbmDCUBFJwbk3f
JKcV0tlWsB8xn5VAGHguFp8IW6as790ENoZIJNtLKg9DrGeSzX2vXiR2/C0eVbhThxPMK/ujNhKA
eixKYB0KiFP9D0dH1kHoKIINcfK0Fiqbe1ALvZrxI3XdW4poecm1ZvMim9pGLm6qL34HsdrSeFxP
sCJ3wTkKcmyuJ9OipojDvbTm333tZ4VdZ1xXLauQUoUadtBVmMfSRRbNGmM0BqHqtlqDEQgXLITr
UyQOYIWtnaZr1cmBHU1hUelQFiZ7dqHs4besIQFzFvz1FqPx5iVN+6tZZIgQPWoEVh/LSYEDRjF4
4s18VEUUaLPEd9YpdQ1rASYogmBCbM+3NwiTFfkMU0ka/NgB8zkweqDH3OsG1yHcHnmdgcR91oLD
K2TxlwG+qdQSeweqtHRhrTYs1MYt/CoEZa+aRaQ7ndbIv38nTHGkRPGS8w/ektkQGXyC9ihkKqvI
Q0RCAFjrJAtxmLD+V8JBsw12KZqm0PDw2gDAgImRG3GjeAsuX6QIi4dCFvbz0y3UHpbLLJr3etFM
+8j2eeTvYdSSC4Iv098FlKs61+vIy136nsmGMCB50KCx0/5n+XpNArdyV2Hb+B10xsou40xqHLr+
WNV75DS2sE7rz/36MXVpjGHpsdFVGhhoeJfuQ68oLwXak6UC4eoD/UgRcx0XoI97vDLcj5n1bEos
ZWkELIk1poq5lOVP9+h8oZ5DAOrgz2KvKGy8NDm2wqI7WabffOeY84DmHDtsoAI6v8pSiRs4v9n/
uW57a8/Qucs8Swm98r8cYaoG0mULFA5XMUhRrYFuHkgt/wlOrqHi0Lf1m+EKIdh1l04Ce22K+lNO
kLfG0K4w/L82N/FFaynQlDHxsRDpamZVd2ZN34OeQOOZycHTXuIXEsDk17jTqpA9xm8fAs33rZTT
jM6IYoEo2vgDwTPNeMWXLtBVFDxwwrzj74s84x4Xq+ZlqKX6aSns/KToJpTNXi2p1dnHfsw6a3Zv
3a2qTF6Q+0xlmkPaOQHiRqPqpbsor4qybARta6D7qOKtNbiD1247YkYmeHMdyClwttEwMsUxhreH
5+/t+WI6ur/JVDSLKQ15MxfRDBVsLxoq+lSqive4be3jJqLHfSrcaEB5TFvagheXiBmEp1O9bC0A
UW8MNoERDhNbauRVtXRKO7OeHENtU8waz1X6Zy1NLNKfCfrb0eWqzLa2I81sR3vHZ8nEYJA8HziD
jSQdbio2/yKEiIF+ou3T7VPL0Cm6micg92R5In6n/SW/aPRXGfciz7V02Qp9Cc1+EoDeBGpIkSvZ
5Pd8mRbM/aszkooJ/a40MXqbgEiV/qXBbeGm7dU85TTNSpIlSWlQSViPSzujtXGmuei2rb/OcS7M
txB5ydjPa6xYldgr4Kq0yG10SNtD7Rnad4CCx6sNteZvcTCj9z3rGxnj5TDZQBTieUtT9+Fsv/dB
mQqqYUa7jOBx1BOmhOGwLb4on1syvrT0Jpn99fJV4Q5fM1Vm2jm/j1gi5GLuzVRUZRu3hYWnXGWU
Sqqe2onuN9NxzRV/49OascQuyQh8YyVsNSVmu/KJ1fUQbWvHtLuWUHygjB8hEOhw6lqS5ITyE7wp
pKwqlXfjd40gWzHUGEV3PlKOZrtXbRiy8vDZ1aBCiNNB3zGMVoMCPFJY3wmr5I5//G225XJrU+Lx
p4G54EqLjw1CDugBOpeE8Lb3buIeIwWeQAazN3EGo8evuQHbNljxFAozXDY4QT8I4ZkW9CE2hchk
fD+y/SwR9cDiiVxtVDEwLQl/09a5YOiEAmz3pzI8crGcKaWaxk9c0vOzBfwV+wavrAAN8uO0ndUU
ERXDkkm+PzHE/OjuODt5U9jWeqS0whIK6byPOWMIsq5+JSDby1l6r0gI0YB9Zg7n5lG92xlYA2eK
HZnFZX3iElNpcQBCAVf3XiLeUQcxNQvcdsMH1w8lPPcQOkWAJM6wnAG18Z77P64YjKg9HdE2HFb2
SFU78kV9JUcabY8iHnMw0tuqaB61eUQeHtCOLimIdURwTZ4wWV6k4U+bIgaCK3xPsIk0seDBpekD
qOqkHFGAByN0lXlWFmHu3EaMHatcwi1ToydnJ29K9JvZ+syzXXTPagY5B4rmH9+U2bOByP7578wm
RV9LgeOw2/kY2vYteYUCauQgNx9fNpQzeUjro2AT+pTYf5h8tatPf4BARpfWBYdzUVu+yrj16nvE
yXvRsK++q/LJ2AtWKhmaGG9ltg96UCIJ1H50Bs+yw8Cq1ouHoXgALOM6MNa/2B/2/eX4teTPnAu1
iYBWHEW67o3gEM1upcK64jkTN4532V36OM5MqQKyS4cRRU2T8Qb/J9q+FRuQaIarZir1LQGuesN7
OcxbycecR/LGl9WXUqQ3ixeWD/xNZMBBeuXEFGf7GpsFUvpWsLwjJZOqna1oIiAcUiN0nD79UXL9
HVGGWaMfucgb/+yCt6/k9U7qd0D26P7pXFnJ1qC9/Z+PF7HnKLCgKoWDNawhlcod4gcj+U/ncDad
yFIahMMv2nejut9HftAQEsNWHvnmA8i33Z8TxCkd0dg8T8wV63ddGUg8dX1cfQwrFATHk7aNhJnN
ksl4B733s+oxDM31h53vMjCLqs2kkDzsw0HEd6xR3YJmfK2a7tk10OJp7BgHdcpwssnFRNuJCk6d
q20xThzu69cfCNFXMGdd3xWM8YVQ0p2FKVgy8JTUJWmqudvBX94zS60aUJxUh356XjmQkYaKPyCR
SSIyz7TId/nlA/u0v3eeJNZMuJOvzW6nuLaemIMJAKbQY0JY968pEvrlvOvpEt5we06YwQenKspm
G0otE3UrFfAiNf5oVqqI7N8mVWR7sgZMyN5JYnK1hosBPpjy06pQpnTmx2kN7vBO2eSEhPJZik+P
iLgsTFOnGPymhRz+JTJziNx9kKt6LD+sitP8y4Hb+bJF2SfLOqZrYuSnWkKDX2khgNDwchNnY58Z
YKfv/CS/MUWkakbcar4UzM7u/Vf+XNPDAUoPgCqr1IkmYXG4CK7kwksIGT3I5zsRQnLP5MB8OENI
rZtV0DK7xj0G0RlARgpQeExjBxLhappwXdKB1IeUPqJYevmcMiBjLrs/N0dsQXbgaAZj/0uQQ//L
N50vbyqLoe3cawmVnA20q7ZcTUXJVqi01+Gj+ZiGY5wbIs7BXqVAYs7pkPjuKK3yq2sg75DJPrdM
x7E39J/68K2kKZC02g9hMBQoh8srth+uz0QBvuKGjMYy99VpmscWTTcE5QPSdLEVjWwjZVDIJnsu
HPtJ48hXUxjWTHHCBBb93taPxN9VX9zz1ryyxNpsjcDt1IcNUN5mooIJQlzVCUitYYKIb/OttJK3
7ZCvjmJFjx2Bo9R32ZK2SxOdS9sw3HADvSPkALsVhPNnfXQ1Q9TywkpqLhugRVdxPhfUSa1R4l3i
cNIlAEIe2tMVuhGEnCyK0oBxdiTtjlELHVjM6Yd89uXcQGiwzolMd6O3zNKOd1wBjPK4TpeC6cjx
+RVEFM0jRMhrEeuJf742RiJmtKTL77WcDeiUUnAB3Nwo4mLtstcXYVKwVwwhyrDaPRNRJOKqGTY1
ikCGVocUmi+8KdTErY68XL1bD2UoDVfkX4ja/uEMnEVteX3Oq6Dy7XsXsYUVtXIAARQK1GhM++28
THgQM6zhDg25UFHYF7Pcm5x/nMOtcI9b6EsSkWB2oM62X4xAh+tyRTZvsGzs9f9r7KEfEcIMpos9
cJATBo714SPTO/5AvgQzU1JTaToLvk1BvAQIMxw3Rg5slfZrmcyELMN2IprJeJR0fNMJTw16kQXG
axkI02OqCGo6DTZDkwmefYmyrXzrrHcl3By7hPjrv1Lard945A2sxmqiQdaLs+ddf52SpbtLqdht
mLGhgRgPq6JmplOa88iKR+4KNAuohtGLH9tvUSZDm2jVawS6ltrnPQz+ahKZRmRiIWY9LPeXon4H
RzqoUva4S0Io6aOgOnZUcF8rdfQNYG9FMWIZ5bgwlVydYz52CW5OFeNDHyz1lh+rGe8B7dbSE5H5
Uo6smWeYBpZsNHVGOcDkNMR0aHz63yB2lPqXbal1JBt3VdwO/C0/WtS+h8VNB4HB78oXNNiwJSu9
U4K6rlXQAgiTrjrttCth1Dx5+NPq2yc/I7JYtfV9kYn0cGpmpRqELCoswGXNsZsdZ2EiuNf/o2eh
va5lkHAhXDv/Xv1oqLDP75BYJp/JAd90iTlBr37MavODCUkA2/7Gd+OiXW9ShdaQgmmvK9OANJG4
bD2nLdsrXBZtF3X55QOq5quIUZxgwSGdgdowSk8r5/wbq5SejI6D/gnzJ0aJe/pvL8W3KF5/akL8
BD9Cn/Pcxdg4X+il9LncX9tvTaBQJsIjsmoCDtOh8r/4OGDMQ5Ib7StExPaZB1mN80+JdlS/waxe
wBdLU+TUDyLr6hU5acxwPnfnVWrE9krZh/x+iiqlIRoA6gAourE35LhvV86T+VyfINKbo7wFeaAH
F6xRqGKH3hgurmM+LBOE7GOdgyENWtxixFvvyBXk/e1YJOct5cNMFZOfHQZe+VNQ7l8SVW2fa8ix
DE+spTj+5TKvrAjwXobw6hQvVn6RuZEYWavrhr2v7fgSrrKj0yEIBJNQ+SyKHmNvOkX046GSDudb
ynDJJin//6JrvzVFtd3CgdEYoBC86jY5KNaTbzSFsCNYaL2c9NAiUnYV7a3Z8LN/h98ep/cJHt1W
Shd85nj98zVHutaHE5ENeQ/zONgGydOEQIySjMyrS1Jz2jE/gy3yHsN4wywloK3QYv+F+JpAmF3k
d7A2l5VHQsYRhGlukVCzP+YWRQfXmqmmV17ZpY9Pe7J/A6Z2UWa2usrVJb2L3O9TFzTOhXoiLTxr
yF06iCzB7Lqt3cUS0DHmzwE0UmEVFC8o7ibyuzLtwqqqedKq/GRpzHymGLi0l8AAKiuGu4Sp2soQ
zC/PShYbe78kIg9YXl6fV2seq3vqbxZRRIzwmRnUjKIx6OHYqc+jIDJcT/yk3L9Yz/lpbDmOp13c
LMlKlabj2KSNzFgNXrjHlAfIiW+sTtORd7N4At79CzECq1JGTqcpTJGo7gz5H/Rg0bSsbGRv++YV
YoDqTMhqTAAnuy+cW40pap6D7teH6l8wLiTvsN0hUGodSXijgJDNBpdFTR2HODIYCtPQsceaf1qY
m6eKToQ7ZJ4GXbhuZdaoem70MMNh2krjPYfhF4wftPaW9/40Klg/gvZOq5NTVhtaC3qoxzaZs9Iy
tcOPP1EDAkZZ2h42IrtoCg1tzsRsy+DVmtmlzF0s/QPIcnOEEaH7JeQta/TABhzahGnamIuO8E9e
1h7wgJk8MsZgqMQXjIrvo7P5Ogz+9M23Bf7cr6D5wLyJ6Ud1/9+KugZSPX+v8vJu+ghVHeogple2
ngekI2fBZv/7seMkewdUWiSnIjhXg6r20XyTh0un2AF2Ydmh8L0piCRCE5Q5LTm2tl2Zsydnfyw+
B7vCB0JOpBgF6BudOvxeQMmXbAh+GCLV9+3swrZtl9BCrgkxiFUahfpO17doq271aIWVX0z6U2Jp
9Hu12Pf/AUIVYsmiVp/RztLddu14nqm/j2+TxYjWIsJIL7VsEUXgejdtNmrNgeUfQJuLonZO4D7t
XPa+EmVih6elEAfrOkrOn3ETn2fuOt2ZB9L07dq/mhhkD+Nq4zVnSFUUk3FRl27sKLux+YKZq7yl
P8SVawwo0oI71mMxoszPT8cB2zyenrFp8GsbeZ7XopQ23WQ5NrDmdaC/kCu9RfVcYf0bydSgqvXr
+tbdPUAm8f3nquNd1Cqin1XIUbmjS/DMR2otMyeQehM/PwzRTVVXqmyENod9SuxKujdZxNehNike
4iflVkWUA35xscVWTAkjVPEF1xW7f2++7wAchqVNBJz9e+nyu/scfxGDl9JuX0f2WGO9FEEeuoXi
ul5X04O889hRmHb1ucHm2wDt0yNZxaP5qZOqlCxkEODloWhFLQ4LkDXKOkyILDynn0RDGLOhniuF
4KNCa8eaN9EbF4gjGzC352eZlfFtnkeyhP/S8G5WT0iRxpg8HDz4QgJ21FpLJhaTtHQJ3my/WgIz
PtGGAN/Et4+UdhPd651cARvmv3QZw3hy4CNAlPouAhMUTmpacYDfplEhe9/6BhAc/Z20DFcMwdGY
WAVvvBlGzGNmsQQO2sfAzmlI8qF5kTRx6rJBQk1KX3ozP5Wa4yCCzU5CB8LURBtrC/h7fgJ6JZp5
K0rvzSzY4ALyK26Eg64mVfSFrKs8kpiN6ChlX/LPx8l040yScvEq4qPtYxrxlmsqPsobe9wBbY/M
Kf9GQnNcZhodEi39wXLpHWPvSBY1gdJCK1Fvjpd8bWdMmctyJNs4t4GYrM0BEjOtsQ4oy13Zodei
l2e/L4vxXK2K9E/8Rc0h+ulbIdBeCbytyaIXvq9kuRMZTAQiheopr6i3uJgXKami6hynRP8d5lxt
uqagmo1jRjjpAXCyNOJK/UTdWZFCiEhEwEYCVyffD4XHREsKwKlBczMgRyylMdprlnt34nyaFTBZ
yNrsAIYFDrRsR0lM/n4H2XK7x7HCwioaNL0nSM7kUI18upt0KySlPTdHVGF9HtMoCDkk7KIdMd1+
eKlWCUqUUJI74NHQN+iNVqcnxIOQjo+4NVMZXMIKS6h8q4ZH949OGVWuItGlvkyQzofD8a2nsfFa
59l9KpPWGTIdiF5cunRKLj02YtdHd3TNCTYSzyvNX9NUxCrDkA2AeEKV4VuC2J1EYLMAMrfLghm1
M/zFYtmFxufYLAmNU/qKpvnNP7+8vzZoCDIzb/ZH+NDl1kJoKGAAozLPtmls86SM5n0vPK58jRKI
Rni6+nlIRYOLWWFOcbWLpJfA2nayMqDj9OC9RdgIMLrs2P96C9kPpzRaoYbGCkhTr0jt+NhlJYd9
wQ4S4m63uk73VsDWmjKa6Yd5M4FqlxeksJT6ehIGjNb0iVbActJxbFJj50Zg5TPRigHQCiFsQhRS
Q7dzF6t1yVhVm2BOFH2U+7gpTIDzAjeT6xKdsqa5wUY2JNQjdjcSZlC9eWLRxl6LMtJ0ps6YaSR2
HQeoldPlup82FPBVtqej4+tMPeg6xHOGwPTDALizLbiuxWA413fiQv0SVlGGr9Sc+OyZLM8K4C90
dwq5w2n55oeXSeHbPUdyP49ETFsB2Dpq1imQ81YEpeZNFvwqONMCTTToHgImSyiVwRy6U53jspcb
OAXzWELVxTnOxn28upu5iDO560e6TCipxRT5jmYDZnlRNiFgNbF/aeR/DV+zURMij+65RsO47D58
oXHyjePVG31a+rPNCfG+k7HklLJY1oHyxOvK6sUhUEsCy2QMzuOTv73jjkser8J1TutaFtgzyCVb
1sQkAh7yFNAjU2CLLUhiA1uWVrQR2SNCNZDwuQtLch65I/h2Nvl3qeyAXN3QgNQpJn7XAQmVtAAP
bNRqTwFff8D0k6gQP32V9myG2NdzPBz30SArIn8k7/a+Xrpa62rDzWCiJSSYosxmhWPLHvTuglak
w/cgcuQgzz66OBa0obet+wq8mIjmC7TZaT0C3prnNMxZgCWU7BOZcvlE6soJfu6LTjrOwlBcau0W
40tIiEzOj2PNoQ2FZZ2UHjqjXfK9EeAMF8/69yXgFw6UWOKP0Pxx+iYYp98LvFASdpFOVskCdS6k
wpwdBOfu0QaBaYlIaiqvZEUCubmZD2fot3y73oesiupt1kJmK+UaA+kgtv5aHa8MxIyoYhjX7Pn1
RavNbHV4ZKDg0AfmWHYP/2baxqQ3hG9cAxAVemuY00Gk+/5NtJddzRt8+iM40pJre608c094T/Dd
7MKqZ93OTnFqta6vfzVLxbia+eQBAwToVmmWW4SXHRbH6SKcdnJBO0l37GukUHNbFHxK3HnkBJp3
K/l0a0JQHtzu1G5+5RUdT7ZWOs5EuFUUEtwUSZ9+vrgsI8DUh57Ag0cNAdnlI5oWvHOKX9VwOx+O
EiGBTrVi677cqdDQKQnByYpSUdF29l6glex21BTvpHJ7qYJSPPbm+UtRRgCbmpNZ3Yct1pbPRyCC
xgoVWMXbjWGL+BRE40W8Ln4H4UpI3qwqSjtHpXY+oQHuqMDynCLiukGiDdVV2+lidi51G/vAJ3cA
WVLqOKVJHcS166FR4F1JGC5Kf1zeXCpiwp5FyoIAYJoXZpsh5A4m605P8UoicDhafLqLdx0EQ7Bb
DaOHqE9AGBtkCcTKD2lBgstfblrDQUQAN9KjBpcq6BJ8jDoj92DaP6/UQpsyBIMj+LEhr3uQRiTH
RUc6ieV81ZdHYw1HLXwJzETbwDSOlxwnJcbz6M4Rfp+Zm2JlxZWBlr6zUqMVH2pQ8EzZQ6EPqGeP
JgWD1oZp/uBMpHzDjw1YFX3g7n8tbbce+kzgkvVLyqM9GvjEZWbF/QOu2jQJbry41qekY8jgSem6
pPrIp/Ye5EgTHqjgFu1wUgWyrulxrrvZk4eqZ9w56Py8VQAGYmyqTyuUnav8uog4W0OJaXGhucMA
evFondaxt88tdxEm0Fkfv89zuVoJsf+XLsSAewWRLprlxxHX03F0bte6hfbqcp/5IoLTp8oiZ5mm
LjCX3HooHeiecszw7S9v4gsnJH0nmsA1HGc1/jJ0ejC01boAO4bbfOLxoTK/rlg0jo7YJEzhV0dk
8XCjb2tJX4RUFhLBXgoDrpFmTmkhFUq82yEnBV9GLakpDBjlEXAuj7Sd4h9w81hVgLgNTGWsfSop
PakGwZryZ4TPRuRnsyPuVHoDDeOhrChilR8E2447S0gmgRBVH2JPVGHArFFYeArd6XvS7VDZy08F
bbXBAz2tekHakmSmDcqDlBNPKgVt7/faDFjonUJvOG8I9P3hWuKbOUgpmxLzEfcBBYxQPEKP6FQU
8B33/f1Gta6s9Gxr3JW/4ecsjFYOkuyBwicveYV9A48A0eI5twxJwWu4h4OOMQ94qOCNx1GDnlWu
HBJL79u3WSSQfFUchJ0haxtYJl7eKO0DYBCXWoUBqrKKoOYsGaxSq85QdK0wcSnrZghr/udN036x
ruy9iHNr+5CuFD4R+WQoBluAr90hZnPb4a6Z+jqG27itxYopNb7S8Wa0Ocj9qtg3FsX9RUCRJQ3L
rh7KKy882OxwLpEdq77KyxDKRIc4XqjTk8wtWGCqO9pllqproE7jpHT4jkbWy5oSzbPuvMTR2YBi
ChAEQplFiDYUE3evuWvefwf5D3BZbG9UDXQw3JJSJKeSUahrnFImxRBB0YOSL1SL1Bwmwb+HJ8bN
LSrkd13z22aQIBZKlWBw7BPpQhmCGrjtAlAir5VaUnYv59a7USpc3pkJLsk8x5AcoU8yjneh2Xc9
H5j/1aCex+agBfdIrtItWjHLXnTaPeUUfbHYn+pC7O71xvZUhF8HCncKvj9Sf1nksXsC0JP/PIXa
DiVm8ICgFtfXVU+odo5KUNLUci1ZHu4V+uadEUBOSPDdvtkO3uwNEO3+U/75G5ffcmI22Wr8dP+3
567WykY1ew+0cHNb1G+IzFBGEXd9MbSmo0I//gprjgNu43aRM5bAkSIgu0+srdD3x/A8J/vLG4X4
E/bGopx9gTteQa22cy8g7/QnqUR8p33sBEsww7ML6aFj0vh3x4TeXenOgT1JRGSdeyCDpCtzJ08B
2grWQcuhz+skL9AEPQttBQrYdRWS/6/XusRwZereo6hqVp2IHMQrN74JL4oNwDApO6+eWeZyaHei
o1P1NQH90kGUash/k8wgTOqcqkm05f9fz9qT9NG0yuEJXhJxcN9WIpcqmrAcZATUwkmmq0aBCdfk
aW0onEKdQSmVmAmdCpGCQzYxgWUkA51FRWakl0NuD5G8LtcS7JJJ+VW2cGuBc7UY8e6VllEjQgI5
pe6S0kCIVHYUDvmxiUptcZGF9FPm/797b0VwsYtMTFjm+cndPU/uOQDnsIz3mRU8QGb9w6wrgY2t
B8/h7eax5VJVNf4bR4FLnzohoklEDSKlp7JU3NU4RC5tU4HQFKL32zefMM4Bd71RkdpNsmVgrTXF
hfGHIhvME27VtjsxYz0aRQkfq/GBuo/fAdHk+0FAyEZtWRkrhYq3rxGRZ9q2pCDU9tBiboF22JfN
TQudDjK7saSClgDbyFO0bU0m5HYx7hxbxS7WA2BZl47qg4frS1TkXB1zCD5gUQEf/sQKMNmpb4OE
zjOMGWq0ceRFOgsuWgaZC/gGWjyVg7ZbFZIAziLSRMXHVoLZwOma4b/PvW0WH9bSs4P7W4S0BWKA
0w09+6D54FUqGYyaGS+p697OR33x2kw7WhH7oj9PCciHLG8qEUp1uNrWIqNZVn/QDV7ssdWKAXfJ
2mq2YNPOTfz8w59PnfwE9pmFldzYYkYVpJhXfQcLilQ9fT3w17ib1PgzouW6VCNYXjyBLAHDRBTk
Ea6ZRcadtuEoII8rFLo17TycBbUYXcm6MdvNPOwPBExRpJTYXPULDH8dBmiVAerYN2UwNIdqqwxh
qVTXP3j8JWh8aC7hqlmKv+JKg9JHxWT818Mt1sfO7udQVXzxdN9z0ZgGGwCZlaOtdlX2gXX0vHPh
1/f9srRaUtNP89vJSUrEUUxl8rrRhsJPTdpj8hyTJGVqROw2rxmoKPH8/3+m3Nz0QSl9ltotsjGP
p1lL7fEnjNgB/WQ0hPWdJmSACuBX78pC/KC6s0r16URr29ePUOSf/iyiX68N/3FH8M+G1L5fZMDf
y8m1NAIdbLmge4PobCbBc5wxCwknTnJzmaibZPTOTRzEsbEHeHXN4xYToXCII7KgC9hKSXpDb9VZ
3rY8MWgZF27KEX5CMiJC5zMbYCW8fIrVWHPz9vIdD5hgZkNaH8rnGrYrebOoJhHnTV+uI7W2Vh0a
UhW1nvgD+9Y8DKGOfJeYn4siA8W7LgioZK55xdGzhUB68f2ftwrEu3NMokUu6cu0pLCP44S71Zst
5aLvKHAALgECr3xwujwEwe+SmjduPUz5tnlr7r6wsh25hWQJHETHvGy481yqN5QqfNZI+ghpYd4Q
FV3MLcfiph6stH6ADh8BwpRWqKwDzKV46xoEt9SrBCP7OlYnln1Og+xxm7+PteQJzYCQDWPOpX5F
ixMIvSuo9u5Bn2Z8/pRZBo2MRue3r/tRT/Q6XIzVGnbeCR1rH57NsizcVWPABY4i1JsfiZ2ZwGk+
aiyA9/cKIOdR48proptfXSzYUDmuZ5qI/UoRJeg+o/9cZW07Ft120hWOQyykxQxPoPcdVW+QR+zV
P24RruiFi4QZO0KSqmw+rczgEKlZ75INTh2kzJeZX2B0mL2fcxWGVORe92Vh4tUDD7j4Ap8S7L89
inJfSdfxJ06KnNCt+ab7YsCSvpB0Nbd0uxE57Mza2MVwmD9NzU6HEmw+x9iZempu1S0S5/HsKLwr
sgVhZqMDp3M2BDl25HSIGEm4iVLxw85FqhL468D8oAaw4MOOuOJnHh8E0WZNjq+tmppWm7n0YG31
R/RyMWapeWFvDOeUxO3L2Q5QVsucRHNRbWITV3drKEAwsSeDXh+lWgmgYtFMBQ6xeWB1PPt7iJV+
L3QlpktR9Fhrc085aIee1sz86NPnDka3+7a4vRXYxQyrjSfH6BYhcuJuLI6+okGDQ6CXxAv6wHUj
3DBWUY7TuB5fCfBboToiU3vM+vl7R9BOzdEsWzEWPZJxIKV/qdja8xNJtCslOsPJDaEq0rCFPePn
Y554kmlfPpNf1XexH5kILvgvEyxv6LiuB6/kEsDCtEIr588WqPvVOA1/ch5RmRyWP16kABAdC9bv
JoZjcm5m60gLVh5ns2zqlL9ir1mgBesCItD5LpJ7r1K6+I+gJjJOlHOcb94CyJsI4OYxPQugA3ky
7XKr3JELCdWK0JztJ0afKQSLjq2Y8H/AiLYQ0jFM0VqNPjc7cUx3tvxOYAerT2wviSJNcr1CVh2u
n5N6WYtBYB7pJOh8OjDH5agZMNAyUIcYLKi6J9jSAjcOhqduVW1EB0sz5IHWe7/0zLqrBGifB4CB
kPytetqbMWayj/5fZ/Uu8hQxRRUdXvrR7vrZdt5SM9n3PztKQe0I14RM7gkJJZQaQmj7H12floOo
aXluGHZye0qpzTU1gwNl8FYi4Chh702oRMmxh0QOcTtwlm689pwcMpE+x2RQpXves6jBApbLfdjc
uCdJHMpJGBh+AHoBK9nxwQrPpKCNJYeVx019B4vOI6+GL9+WEP8Lpte/SJc6cdpq8/HPfEKmdyOi
24lIPt5Hc5Mx+leqkurnT+uScjmuGQQsAA8AGpkwQLNn9wGtf2jwvjZGn2HyuDL7W5SV1Km4FPIl
EHMq7fYeZKVIGHxaEf17O68jBVuaublVd3OW9fZFQMyf06SbY/fZQCDY/D/Vj6E2ShnFwoRZAgM4
VWdO+XKSo0apKwwF6ivZaNnQpeK0wOjs0Ax0cHou0Lv6bOmf7YSOQCrx5atiLJtl6P6F0FNL4n9/
ZwPfhqmM1WKBYxklH0+8oR3HZRZf89qCNwSHIm1LH3yvgf88OASTfaiftOaqcCGFHd375OY39MFH
MToMKJQCcJ+nnYTQ1DwQcR+PKcpV4ZRjPjiIhxHbQjbT9ugw9SXVawNeNnj3hbINMou5zOG712ke
D6Fgs7n/nAYj8qbSi3Ic0PmVFK0ZD6r29Df5jPT1udTAoqGYmy1iFPauiIn4lMnvzTt2O9wDUScL
uzB9wJZudrzUv7htwsRpAhJrmJcglUq7LSeHJEyW7/G5Uj9vYS9DfGlGOCXcyI2GlfGzBLwT0fBz
bLhZnahtRbY2A09Mk9wiC+p9rtT+majryYOyuq3l/bb7y5SkfGafsrk+nuWxpS3knF90tZNq5z4M
CX3rLZbJog+scCk2DU7RB8iFZkv6MAkGmSXjEbmovoGxInkfTZ8IlgwApYp1tzq1us+crP0/7vqH
VLTzF8H3OaVmvyR0ohhyQT+52eidH/gC0fUjiz9jsNt0Abrp+vt1isbSqzc0YacsCGwKqmobGVAC
FREBt0AURwuJin+JX45qvdOV9Or3erpXy63CcUtDy28cRZAGEpdA5R+BqUstUhmeabGpc6U2do81
XNiO8wuQIYHj7oTrR3NVcQAk4B5Z5Z2oHlGOhTUNH/CUJXruYM4aIK4g4UsgPwWCFV0/1C8ym52d
BA3KzhoErRzUh8NPk4kHHrpuuyFJdfJ6G9Pjz/syAEIoecAjvKhAbjJthXrEt8MqlM7BiVnvWFFQ
92HkpfClbznOVFOB9XI2QQoj9gX+bk8Ri1z8rOopkmyQqiXgcZas++YnjOp58ANUkpG5fxK43ly3
zFGzLSk9CT2lnOVec1wLSPZwHO4MZJw+OLBfr12CmXXVJrzH0xJElKGj/aXX5ikGvTEqgn83opi9
6n9SOHArzmgjgSpu9MTb8ePRmim4w1s2oQHMXABTakSmRia5+3stshGhEwW/ZQvOPFNOGrUvfckI
iVMIs66S6AGH8DR8k2ltdAlgyBfuqORs932xO88OD5oZG4C7OtggNJFKAbMyDzFhpsbaoUN8/N8I
EH1ro93dtEeCoFo+q9zkz7BpFOCjNui1hGWi4Owp6nogM3LfcZK88rZgzsOygHkyOKVnfwOQyCoA
rIHD4u+df8vRiuoRDDczV0T44jPdWAmBBT6B6ivi15sL4afHTwMTk3YCOAIZs8qxMJr5pZY0LUlE
MwIns0VVYd+8XYd5nfcJwhWxqGD6XAuofZ4GKmoWeZtpzwUzRqjCtNID+WVHAwS3GlpFzCUaFV68
wtvbgF2FXrwvwgo54TPCjdfX2jymnZt7vV4VAIlTqoGKyRBrF10Krv7QEu5dMWlHV8UNLZmtpW3X
5vDI2KhVfoYGjWp4YvKJqnlP3IgQKcbMmtTNowsEbx2PYEML6SkkWjciezRjNpgTP/CQDiC9vGj1
zclycx1CWz2dOVr8jv/u7tbyUTLKd3QhyzdDMqnX2oYLJq4ls3s/TsoLqMVDz00ckcDVRxU/QaR8
RvPO8ttFV1ZWnTptE7ZpH8unw3IOVVoHV5yKB9hRbqDpCDLQ4ccnMfDnI6bKTpxReUz4M0RY1yGG
ovYAdbWE57uOfjfGY6VDJ7ve0Oct6fFdHOlNnH7MI5Eb4GfJw/v8JwgN+/bEuud9RsJdWoX+cz4G
RI584hBuDpyU6LsomWWCGUuDITf1/vOWC2vdDLdwa0O37Tf3UwcU9NhwAgH4eWZ7+v289gUL2Has
899+8pNEA7v39+BKRRMMSCjGY09ndFF+Fqmfpn1IFXtoo3hEt4pExDUu+kM9fcjVcHEdBJOnCfQ+
lkGtyGUhtpZtPrqcmapQDW4E2ro4iceXnFs+/xtS6hbrWI93WQsVRVZCgTYFd7xOoNZTvMgYHD4y
zu8w3gkzeb7VrQ14YSifFjIhouFRaZ8NFJ9jPyhvuYLMZegK1FGhdoy4zLZvIpVtmaKWsEn8t+HY
KvIiDn6u/UiZ3iahXnQvOyAxDa16KZxCh24bxwGL/51mPqNIk5ukaldIef2X/Acm0uqSHpORoR0y
xx5DvdfcKFheUhy5X5xkGeMWDm2Jse9WR1h0MDu8BjNRyDhsgcrHAI2s2p3XRYHLQpp8pd7Edt8x
Zh4t9pQGQbDTLAlpEpyIfPIuKhvA3ZOooGOOyzatr1G81K+icqHFaLMIytOGS/PXawv139r/Hx8P
hHNm6S4arCAHBUxR976xAMdcnRu6ZV+Z0zm/wQItt5QTwUcoJ4b4slLFQSFVVRIXS3XtR+ERKNwo
sJ4eO0pZaoXd9eNHgCPvZgW0q/hQWQJuNaBS0fgDqEAEJit6GeY4HV/HdvTdodPy/teCVbySKkgR
UOU5qDF0YBN3fgUHzVN1ujHbpt7z21JuOF2yXxSa/buk+vmPlE8+azGspf6EGTdK925S/OxM0VnC
Wtxmzv84qAyoiPZSbNZoxyNlzQzZjImTHlQJgYURG9FOmqmXBYPkTIYAcgOFa/LSyU49I8dPUi9T
UkcTW4KWrxbxSGO8a89gPwu9bsJPAIHrHUdGU624/zuxRxoqNEZx2j8ER9ka4MxO5B9QG0Xr6Fbf
EaD8gAaLC1YFV1ZEiXLL+jAH3EH49Az+ClEzUQXyGib2llNiu5FBnNLEgeh/kYjX56KMwiWsiT3o
pDYgyP4m4GJnHsoyGdXBBAogte6OTI3MSWH9Ee19/a+G6zKmAnlaB8aGLXOpGNaIzrGLUpAwAzk7
wUt1/gieFdMALxvrl2fR6z8SKqhX7fa3AqtYm6ErRT7ccppuoDe1wBjR7UmQlZCxIl2zVjzoT0mA
6DScPU7lNESYB5Kg1SasjxNmNuGp4oV33/OhJYQcJ4v2jjKeLjWYXKKRTNbOq8fvphn9cSqA74nR
7Q2GQKyPlLXOnv0QlOFhdevaq/zk8/H21dGQHWUpZ0dxlmWsNS/utcDV5z0QYAToMr5zFHqAPBCa
Jc6MEtdv3z7K6xtItZQ0eu5V8EcIOf4lG6X8jUpZpqUk9LWAvCkAQKEbn9tEo6vmFhVmNHSb7FMC
MbMmZzDN/BFv/XUVvT06Dvcm2d8lkfd+lMGBDeBYXCPf38zzvY5JQKw0xG+0HKTpEbLGykjNIDtl
hEvN9cODoFfx1jOfFTqYzw4To0Bp2eJFmQm2PtvJR34+fWOPtP2Ywjf2GXemXRMOUmQXhZbr7R7c
u1EvDsePd8bBZ6ymMk+qNgzsSoL0ZmH3TeDoeoVjHhlEDGl1CgeruuFwV0QkwWgqtBpoKETrld6T
fGUKkiQ1urmjaFTEa1YifytJ8MOaeUFNXXBVyuIvnsfrMBTSQbUui2Jkit4ciN49O86VF4JOK6wI
VFOUds3fGQR1thrBTOeShVOzV2I574T87s7/7eg37rxzXQp9v1Y/rjeZQ+UoMDNbXC7OZIorhcfs
DALucxOs7ywF7KYV1iqmi/SJA75SYKrSGKfKEgUi/NZR1xVC4ZTOrTGTayhJSj2IxqWHRGjv7i2J
788Vurh2GagGhObw7S1OqBRR9ugC4G7t20clAdmh1+//V3j7PA+Ojjiiji9K/AE5c3C8LbdbUDWt
phIu0spwv/gtuadjKFscKqUJJDzCdfc4uM2euc6/20h5fchCQTHFGfxLGQSWNlg2cbLZhP4lbOBv
6izD/N2BVXE1lw0mgThpzvdqMQwEc803+bRfAWq/UJjEgp5xpphMinIXipx00+f3EPDKeTlfxiD7
myCNwT0De1mb3NhrYUaUbfTyILPZYNZbMWe1BvQVXO1On2VeaPFVNWuvFbNTa1M/BrG9imJVF81X
debKW8YGhhR67zF/IVJt3JHa6Auef/HJY8o5yvlFSuFcZYVkEeQg8dwRLNxPcf8Ggh6CcWAFM9/r
I+F4lxY+UJQZ54Pc9tdC7LaBgaeIKqXvX0y4HJks5M3XmcOqKAAQX6qjrpIA7tBVnRtErw3IYm4B
DpTBPtP87iqqsSyazNrScjcdCu16F30qu7iEWmX46cbo1yBEUQiElYVnVkTpijfeBaHC3Q05PUTR
4BqMn12ZLAqj6E4v6T9YFnAQStVCgdG4iFLGCMGpHDNFt9WsfSb9874ra7rC3zxjHiiVXINOLfkp
r/It2S4Fn5BQ3+72uSUmgc9ME0QhUSLFcmfjAXiiFf8v+Ga8XpEqoRjNflY2yA8b6qCxg6q/S9dY
f8HcDyCa3SLcU/1B9CfsQayQ3lQbe+fW3NwOzafaHU8lKEBKRhXlyJIH75hjGe/eEOehKW5lm36V
mDXKG5UVeKR0kVHwaMwm9gMBE9AlMvcejyiXlmNO9agNol/tnl1Vd6abFBSeJBoh5FUDJ7n5wABl
kWfqeSgbfaWYdMxxmE9pKmqoOh3GVZJ8/2yMhZ9r+OSOyIZ8UcNJZkcrL6x+zrmYw3P8tEdFCae4
9CD125tTGreOKNxX5QojGaN9ok8p9PUSOOR6nq1LJK0zdi1KZH/C0/DlDj1cS/s+bZOkfxC7+Jko
aNJnCQU/vsAb+A9avkK7Tjv91DdV0wVrj8cB3R31C4fft0Bh1w0yYDmuvdGmr73Tmt5dPK4jiRdM
ngod1LngUlWYZ7VQPM1v0PqHCxbqktb3dOM4LC03VTJX8aRPuRJ2elEIgiepOOJGPAplX5P4Y3yU
vpeZsFNDkMgW77XcuAEC0JiP7w/e3sXZq7e22BQr6QV1SjvwwsUKNmVtzfST4ibwJ4Gd6ue15zcy
P1Wv3wNZs+0NHHzZGcQcujV7ZhFJ3Vs0xa4il/vpJSDnHJXlJzQF86eqKlrqkmjqIikm9oh8PFj7
EZXTFSdMk+W4neZbOG+kf8WS0gKCa1+vKOprBzpUMiVqlT7TaFj8Fkx5F0XDDm9vsQDcxLIlI+gg
AAZWm8gQ9KGtk//pkyPTrSJXnqmi6yvNrWHiQi9ApnXvKMQ9BOnEnrn6y1ActV7asB3E//B+Fv8O
Sq4/zYM8XVq9I3S3ZnNX2kpWlNA1whZ4HG5YP9lxYKtXmCQNdS/qYWXbiwzbyr436uu9uLXAvNLO
1P2gLhIpNBx8kMO7cm2idLDYBMGaQZIcRDHg8d5UA+aC8MhcJDtfzrENr9sdY4LmBZ4EMmRQlSAh
4hdnOgrXeHIRayrQFgDW+Su0ypSCfzpdz3OmBvUUk17p92qI/WQqHcxqkq8GDfr+1ZV5H0VWtCcD
9DhioYqZ5l2z6njF+L0f7PbYeJ8Hz+qvBknnDtZm4GMxtwT4l37vwfq97RfZ722d5KqJff5yZgyU
PZY5V1iIhdCuTN2vOlEmI6TuN9g0bBCvfvbTWoH359yHujsXGpGgZ6fCblzKJ5sTTOR18oe6R2Ya
0Fmg0lkLeXfgWh6WdhZxu2XFR2sy99cwEvEXw8hYa4s+vLV6YiIu8O3W4ycJHdXVQiLG36wRmkoG
YtjjquC8aGzg8U/K1o7MWRVtivJ57vTOumBZ5HBDUNYsbibuQC/ZGKc3s3tIiFshj3tqngtEhvk4
fIZLaGGKHDexFlSuI19rd9Awul8v6QEgYTj4Jk0QBniU6mq2dAKI1FTfU5RWyDDa+r9E8AxvgpF3
2bLdvQiXb0gTmMZ/Tg4dd0wmrsEaHBXSnrAYx4N3JalpbFlomPmCBIsKdzhh5TvvW7mgZvbvoUi2
d9CT1gI226UOqw/rVm19U2t6FH7WweRP/MoUS/ALMPPu+D/Tt8fw5UNsDM900r3DQ0WM/Q5eg+04
58ZNBB66/fjkskoEDwgfnaiZKPeTsxiSUoLQFhCf6aCG/UapGK3ldsQ93oRFaMQIztDqy53A9kM1
wZh/6Milw/1tVyhw0+rDWDFXUXbpavrnW5ozN3HyILuUdRWNckTLkKvZFXZMkloDd+IDx3OOtPBm
zCBOFuwVsjJGaBUghiOmB1cgVVzAvmS/T+iAjLpqKntgA5oHMtq3Of2yLwC2E9kaziK5yI7Z6vnO
Te0rtlYfQQUYuSmb6DpNa496Lmta+RYPG770RbBaK8xZITmkGlZV1FzuhFjhx5MfRji4j/OPdXqe
tQKXd444RD7as3qt8MFX2Awj98Z1m1wG1VRjuTlpbM46B2CS5SHFSuO95eJF4UfnrOqSPcyZGrZ4
xKnkCtzF+zSjlRW97nHQqrGt0wDHKBG0XxTCjpPgZWwTMHNUUnO7ThEQVDlVK4lqvPwbJPXqtoGs
R8DAZ+yoAlb1jwOyiKQX1Vzf5/iaoPJMQ/BZNOu33RElRmAsbcal7OAdoIam/KDxgsQCnjFXtuwG
0oGJ/R/ioZCClYywkET15VmTl4uUWoVUIhCa7LvDKfx38Qhnt/DSJT4kkRtzAXe97iG8Yh1yom/Q
hkSdK7Cmn5khM3RXfRykiIt4I+tfpet9OgsYdpvuBYYJeO/IoxGH50vPaRDimwIVEuNmErJaeLkA
Wcruhbr7Y5ut+Q+38oD8YOtAvPC+NZQf2y6mmWbydtlJ8JF/PhzMKp11irW3Dlid+FAixwObUG+p
ggIsgpd+OqXDpUgH/uO2pKn7RNPPTi0FH2j9ID2cmzn23ymc0ZTyzNZPirXSNdMimEYDqNFt+OHa
0oNMFwV/t0mPDiimp2HMWHohBN+ymsDhufpf3UkkDJiMlKjgX8Mvcf+TzCnnCShUqoThfFWLTm3s
yFUVKtkmAIB5I+JjRRHH2KhjXnEscBhwkiZXnPHMZJR0asHODvfT+GJC6bd7cgYvclxODZxeqcGi
qa2Ol7OmOVGaStwJ2rBPvY5yKKwBmryUtKT0LYw5mbZK3SZaO8+m9xDHiTVqt2vpfQb9U22fhRI6
L08pxemOHC/PATug+tsYisMoSodY2x15Y6SZVj9ik7/d3gr1AmHg2uCgYBljMRa+DZ4yivzaln5f
YTEWd0O9FeF9/WqVp3wlnbIPe+vLQko7sdVjyzCD36AM6fcZXdCDV7h3i5mBLjOKbzNVqHvx19/B
Em72EsSv4G4qMMWrQI1NEi+4MZzi75bJF1AQ6rgLVwvcXzyfKAfjsfks2EdCq31gj1AwUgY8fnXV
bNl02RVk1liuf6n1UNlIacw/amO7h1J+uO6eGxIBgPAQiBn+XvqtgGywG+XOkQRYRR+Wy+jBiBuK
9trIq0btvwDCXGqYLUV/Fdn4l1xCjlwcGtZNtPt9EPt8j54rIBpbJKtWVJmHl72A2LKO7d6fdd2r
i1msuWJVFJXA358RgKkYiS8bct7T+eo700Q/qXjzigoYXKfr4OdnGg6a7IB6EnfZsSCXM1/+bIjp
auXnNOM9nFgZQ2pcZ4tERC6x9t65cFM2EKruovSoYn7u0EsAabfo2WrOhnAyoIlxB6zFn6BKBqS9
r31XZcW0XD0I/6H+fQyCchq/24S1FBlndfMlj2hTUecZpkNR/+2LGjxrQNy2TaOHyFvCeuIrRBgI
eduESQQLCLdHJX2PHlKIqli3AqthRqRbBvrpkmnAiGovBWJ2w/rqX31F+LO35ygre7nnYhUlfguE
+BekKQjsWGtU5djFeII3nn/+JuMk8fEnspQmEQLJ0pSTebN1vKSS/io/5Ap0ZJzCItPi5jrbI7sB
vyF5aONtnZ/M0Dz9BHrOaR5lQ5aOX4S/IB0kd+1sywrMwRiU6SU1CDJu2wDYJExepnWowE7BJTFg
3c523XRm+mmiKcM9bQ/zridLC+Lq/YQGYM/s00iJm97rPjcnpseFqrs7yM+3KqLe+nJ779lS3Q4+
SocmdxQGZsa0NzrKBGaKYxxMjzd5X/atQj8kOnrSLrYtbNHT0JThVuBtrG0So/ttfZXc3lSsQlXG
Ylbuao045XaMhr6plof1P6aOIYgDcjaAjSQvR6YT9FcVaMAmpxdKsursL3YVQCOAcqpyJ+e5hPWx
zNc+K8aiWNDkiC7wqgH8AUbtdZKK6QQkuUDI5MjtM7vvs53rkLYrUKgULgx5/XdRCpgoSR0XA0UJ
RSSobMbkG1TKZ67SYxsJx/eIKMgrnoL8wvSdQGMbF89TUgjdZRUEG9L1qjUV5ASUFk0j4wYZPG8k
REG7TwDWXNTewOeiNafCMWWG6MOT/sv+EIsovgVn3R2PN4wrLtInvorQj2mPufdiRCzhi8x8iZTe
frn/COff2evkledA7ImE1Ft6RnpJy1W1wsi8/njLtBzgSR9wB+V8R1TZW2G7FU8TtX0bcShwRwbF
pgXWTtx7NHYShSd5D5K+Vzu+/Ze/jBHJpGbOxywMpvr9Rqooxj5+YFm0+HNf3kR9nzQaPvdq5odh
5JcjP7YEuSpiISLzRqQYsJxlEczS4QhiklgSr3I+tJZVRoXVd4jFGQQbzmXr/d8BaMQp5563WuPk
o+FAt+sOM7xHV1O/BAC/ij1LtNU1z7Xzwns2zDFK5gA2W61kwFP6K5SFfIPoT3r1Q8F9mrLJh9fu
wC3EtGQ4oVbirD8qS/g+EwVkiUOvgM0Fr1x0NyT0yikCnnfttLwnVz5n/zhI3SMqIbQyJgSx/zqM
YGmprXFUJ/qn5eXG39xMAMYZCb8CGAmgOdC0RAFjutMhl6fyUQ1ZY8ZvxX5HRAByJWo5EM8KBEhe
5wAZZWTE2LTp/RBfjwt91nSH08hXg7skQLzrtbEOsKtHVfMQ6NQ/FJyvMdwvJLRBTb8upFlgYdzn
Mx9sEyLHndfbaEHA3EqGHwrj+lLO0btOQYsx/UxQHPLg5Cv0qBoulTqQdOTJ2wH4gmTFoeulj3Wu
mPKxPO3QnPcWtW5WB6tj3wWM3FE7caIfWxpKFh1onTAt1lO1FYyPpO3JbzliuVGGhXOgfqppRunr
tZMkddFxRVtulVeeF+G/aeJw9CTjAsK3xKI7mn6/3fR3iJKOLmQAwkRJaOo1BVKpRugyLEhvSDgM
EHKlftYfunyisNbM7MTI/QBiMDdBMWHNMLZhl0a5rjAzn1tjxYGsCgQr4WH7Ib4gxunoaNJLmttL
qXIJ+9ebTUR5Lm3wgYtL1ZWosu/BIKmN8NbroU257H8ZVtDuTBPozo/O2HJXBgHwBbS9VyAcZfu4
MVHiq4KqTK2AhFEowdaiBTLA1L+E7w/I8sIIKaX7D9cfKcJ2MckezsUw8LHTvxrhZO0OV3Mca+GG
SritO2pFzxEaOAOKmdsFJK4kyt0q1ugQTmxxzDCsToyWawwpWWbKARXskEb7Ote5tRvmH/AxE6eH
0HedS3X6N1TqqXMA+qgv+eDweedTZBHsJTzrCcPmmQ/ZMgBqJ+uq1H8RwR65ej48Y5TLlbB2o3q1
dH4ou1LL4v30FVStwQSD8lHyg+GET0PvYXjHUwrxmkcU+nuKkdN39cGXpz20b2GsYGacYH74QreG
yPnpAI5LgBUTKunh3XxdgPJXDDKvKoQ2pEuVw1ynXGqToglizSD6Sx1GEKZ8IoWuKVi4eAyre7iL
EetENuoTdaZ1BixPU2k7VX60N3VwDiJz3tL4n+z9Vbr+ORBrdMy/pxEyJYsPqu4C465+xJ3caf9k
h1Kq8z4vwNdoCiS3pfcTTul9NW+bCEp9+2IvhB2C9sqxTRsxOdLpwybFs+4ihyqwDZdJkYEwUJgx
pTAQJJDpl/j3yuFWgftB8OAgQh5IaRSAFQhbLqeaZWpDMe4cBbO099hoSYKlZrXZOA58dunoOEqe
t88mtSguOf+TbvHLr4ZzGUTXVxfSXUxRyz5L+rZbjDwm6GO4/L4T/uHbaqPJLT7w/+lXDOebkUVO
o8qlUfqILwCaHhx6d+Jj3Gn0HV09XkdC9PTQuagTlH8ew9EcktWkPQ1wzh428X1nFnrVcMqAmROb
iSYE2GQ0jlhr0YfMdPU2KsvaNZp60Zyjeq/PoV0AzTRu2Q85tS8Hv5KpEQOQTr51CfJLrzA7FI1F
/VH7Pv7oKLjHE1/uXzPnn3wyvLA+W6mUlE/rRL7SWvCZrB9oJ9Ez+i9Eq2yngl0y6fN10W35iM2o
tQiOMN09SaDcHCKLUsKEa87AgwEvCORc2MkjMhMhvrgd9iRvVrzacogqjviVdY2G4nbNHxyx9v2+
C3EZMmiM8Le8CkQrTruqL74/1Bi8F6fU6AHj2k4FgQ1MJtH9X7E751P18PKddWj0OS7EGtBTZHS/
aCVGqDeympuMbA2a0nWS+2qZ6wQREdBfk76A+jEC1y5t+PaTB7t1OS/zyUGPHKGEHGC7qkGaeA9Q
NwHk9ILFZz6dPbSvJPy1iYnN6FB81iu24wCu3xL0rsF3Lv6b0Wv2zzM7qz3oL/7BoPiG4Qn5Moe6
prQomcy7GYVuDAgcWbyfOucT0Qb7LN3OSF9kyHYg/JAt6fTtUgj2GZA28RS8Cp4DzTjaXJMwqz4E
SofdYNBRH+0oQ9DCgIfalaaVydMVCwpYBX60TlA9lJwNYrn/810uLvo07p8c71qtx0Me0M0xtT7+
MIQDQPSzbRs/qz4lwg9tqiYhb9IkDEoPaVDXwMSGT7fz42A5EgnHIuD8GhvWoN2/Tvxqo34N0A7A
PefNNJ0H7WlO5fnyK6EktCh+9oC0fbfxnbwjrHBdHSVajsTYaje2hR2X+Y5yEoT+f7+rJ+ocAVHI
RKbjy2RcSixBrB3r1DEaXAlkgmdYR1WSUxH8nKneBsd/NTfxUjwH3nc5e39ekWKVYvMyWZuX5hnU
ply6pnraD9YUL4dCn6TpmWMOTtrA01MWs7+aclggdpK5kGNQGconaGPViaV6xxK0d+9HceSc7BcO
X5d1d/VbyPDjzI858uwHV3TPUdzy+F7yBFbIiY8XdNGemjnOwuZ3cyDNtbdJYZpSA1rVxMEUxG+X
Oy6UltOx7mjVK+1qXPW0t7c7Sl5/1KjShjn/Af6Zrsac1wa5ly7j+vHqIgAcnJCT3B4sYoUliEih
VEI4Q92SuOtCcKP86ESZeq2mQRfrCmntebC0qBVHmyPclwtXuin68FO224ETCChr8kq2W4bsUhjT
L6jmoW7zbasjIPnQBzuEL9oK4d9DxkFoDFjE80zis6z6w1yVMXZbRZJVxtXtDZxFIjE0pY8V4ZnF
LKkUfLrUPXnwSOFEeSge5BnH5A1iKP+QTLgn663HD05UTwl3SzGaAyIettIWZDQ3raum2pc07Egx
xXizcJX6bjCKIqm6xzNP+QUONiuaM80i9KDgqTJ4qd3uIlHcbCv8a+ZHa1xFhvZZSpqkJFc9lt2s
Wx2H02whpulhjJ+pKQECHbtWvsMl6z4NUCkEACVYKOmAug2HGJgc6mlITXkhXPUePCMIx4APySW1
zm9I0ksieiX1T+LgA0Neaud466BI2nmRUo8OeNh1kaR2L5EUBYiENXp6bRKgNVeDCJ/5G8hjOV9l
wQtpLmoYjrYTTG7W8/HSETe4Ew9zSgZCs0+s6qNkWckvD/HbsqHmX06yaUn76s0O5CbvKYsS80ZF
ElEp3+RuYLsn/V3twaFBIORQF3WST4cDUuhGdYvTRLAs8Dg++SCW9HFjFQYO70hdLnai2Q9kxhpN
5jZV5isY0IRtqOdxSI61SPTrJaUtjbMl7C7kZeVXzfYkTjNgPFvh02mtiWo553Y+H2su9+tiPW3u
tVFdL2GoRBlMfU9FsNb+6NwVXClUMCAe/BNjvjxliKj+4iEvb5xp2ia9cUaB4GaWwy8sklZtakmE
kuBtboka8zGaQlqCaUxFAoLfFcEblAQSCOrs5QN2rzi+QeTTP9KBMsRRolsYq+f2OsUpJLPNya6f
7AHmPuhbVlxT7d4KKz3z3er07X3RzC6lNxy/Sb7wo/WGLgOqZ9r5csjZwDbT8FfsR0LU/UBM2XPY
YAHHNki5vTtD8OYpLOfPysR867/MexMrhqFpXurhxfArotGHbPiiAyH8YlaJZ/jMqStirPs891sp
4J6DWxLhH7SXa8zVbdRN6ZgRq+CzkNwl35Z3vNKxBeg5k1PYUM9HVcA9hGrhQYJym75fMsQrZbcg
qU74WXxuCV8LWuGIINNWkHBVHtDk6HtZDppAPzZ42vSIkUWetmwkekAVfFFmNLZeLU5Wc5CRVmQR
CVRxdv7Ce4h2crpkvJV7cSVjHKqhMEuWAoUZjFLsA+VEm+jsWp2V9t1UYMu/HOMRU21WMy90FH3H
XvTeYOGbZimhxKEm51YQUYuGTj/d2EBg3yo6auxJl1fxy+5yFqEY3A2/9nu9WJqfEVT+Pe1R61GZ
IN11zf0jN2pLW95fT8x8r3VY1c7ufnTp0ugs/74uJTwU43l2S/Dn50XOO7ZfGZBhMHiY8GCsblge
MxJw+lJomhIlVHq07WWN1dsyg3B76V3oj3Y8bIVdjEteyBr3YB2PHyZZ1WI6thTp6K+eE3Fwx9Zk
9Eh3rpFM5+Qk7XjI33A0TWxnDTCmVxNCOBqv8KuJt2wvK9JLS28QJHxJsZ5Q0FbY3tBih+urRgR6
ToMc8LLICz4tP+Dzr1oHa0/Ly7dwN0gr88dp9uSdNQ6NzXOXArmHm2XUjBhr0/1X8JXHYtv8BvPr
O88VF6FfaenRBjGvPa4isl1YK++tUnh1oCk7xpdddB5rHotIbkglWQHK579ejQHuiZUNl2mOhebG
+NIaeP2EPn0DsdyLV66OPtYdvfewut7K001Mqodr2u0A+GSceBeqLMNypN4kgV9S8yY7xrL9A1k/
Kai6QxhhkCmSM033MjZ572+p6XbdFQRKeGTS+1UnbRM8JVZdlndoLDrbQ3dN5Suw1A2dBDJujzKN
FaaMQg/0m0ZX0C1m5dhnaOo77u6FF6CEYhDwjVBDdPMBPrk1zWooT17yGK0iE75OU5sSiEznVAHK
pjkNCtrpzZMz8Tll/BgUUj4yDkqI/V9Y9mb8EeS9oYGZYWnpzbwWvQXosVrP7bt2YAU8bms9RWUY
QVBFiauTtSdG+QNWEFX6U+OneHyS4m/TIltd2N6gT92afJsHv+2emWyKNJ56kvv1Oart+Eokmgbq
uyV0Ddf2bjmmj22id/MtOc/MCHyiEpmyS74XnMORzwFh23Xf6OyBh1jgKCqCsUyw9ol83or0ZjHP
1HKonkteJcndXdUFfBniNyK6Gq560WiUiKKM9fq7ZNAXrwT6tJmzXD3x0HbOFyighrMIY60IquQu
US0Pco3QJJZpC7Y1wtWp18sPTJYdz8nJ2K8L2lNXYcv9m0ZiEBWfxCWmpuaQ6l5fyJ3mJoX96yWL
IE/y1Th2XYsmV60ru3b1pGf+l+0BBAGXNvUbLx6hzCf8XCsVr22WGR2RtYHlBBvBy4sPSFYAaFxf
aBFhdDLVvHFt5VCj478SJNyLzzLmmJf9rYu/OFMW9m5BtH0HR05K7ZUGj534zu5KYo6cjrCuozDM
VsvYeNze9aeP6L5sE6HysOkeMhXX0L8dwJ2TOI9t86nyqo/MjnnMZDmEiUVbDx6Y8l81Mn2T/VLm
SOE/805ecw/Xn1v4rWdeuCg8h2a6IGESR/rwrpZ93EzT5U+/rSJn4lFJpN6cbZ+WH2VMb5A7cm/c
1UL8Cb1Il1U0nKmEuWI9BWECW0bpYxIdID9BIIgmPR3H2vCc8aMw7UigDPm/hn6nAyBsh0orNBIi
JaX2/2HjafAQ2upKwj2lcyq+uDBWDE983kqzuEoufy2lXd4PYLKjB2I+pjkl70y3S54tzi0lc6ui
Xt3FiRb1cb4nzA4SXLqmFm9OhC/5Tc8t9NYAqXGMOKyUcR0KhfwDreEqaDVAbJcwdFm/nVakPfXi
I6Npxd6gqc6ko+/+dcMcJ5uCnio9SjYFOzIqAoQX8wXQJR1qNRefOJ3iikFSTafmi4X+4Zf84Hhw
qjCB9lsuvGuP/sZmWZ/BDLAX1HTHwJr82Kp55yIhlq/z3rLWwN7qcPvZcUlqwVM3X3udA/etzdsw
uAMbilFcXpDcluoEZm3YqssV0m7Os1SEHDuasqMjeqa8cchx0zLwYfJJPEqruA5Uw1LQjeoCYrhE
Muu5LxggNzPxTKfRmOBWAntg7Rv7N2XdVAbSrCiBb+tPGQvqq0L3NZYoIWI0g3y6Zjr2cpgr4q/A
NpM2LmaCBk62tedQeC0W2N3h5Q1q3B8ZAlai4tmn4VjxShdyaznbvb2+TQr7txGOH5vkfVFg3k/B
O3YSoQhWKDqN58WT82ULu+/Gd6ICUelEOOHeO21p5dk3qdGc4K/ObrjAHBNGbdKJNhaAvhcvMkyz
/0ejfx27YGKAP+MBmf0vdoukBz2hr++1eXF7THHYVZu/k31b2eCaSWGFDH/z9i+C1JQcIWrXIkvr
0qJupiYDZV7G1Ek3SUqwijp5jfxZu0Vg5PpKy0EYgbEUUReXsTvl0lLIzHuKYbqYVjnHUgVbEfeg
XkrvqFJhfUz7UJWR8kaSr/8nydGUFV6WesRC8gcIZGftBiJmofWyPjkKlbY5jLkRvIW+SOilFLdx
rPEHQxavyNh6oSplPbBVbVMwy3i7OSEu8zl13KaGmCsrxg1haPfoUJtp18EfH5EMfz7+K1S078Iy
l/8EsI+MtoLGUNouYom98erhxdrG58D3VB4uQSJR5opS6qqJxgccmokNExgtqzsl/eHfmurt+gcr
C7MhNF+rkQ+o+7fjOjGEVFDezWr14LrauLbmp72WONBcwMtmelcKDoFDMi/cV46jhIpGZ0jrIak4
XqsnfBeR//JgO3JVud2hK3iCcEukahZCk/W83lwianqgkobep9/jiT+V36dnJUjbRFUs7Zr+urOL
qr+u6x0yYi63XwdNuQJAglmKo17Mbf+7wYMpc+6g7yer+4D3gwQqDSr15xH5sCVrRp8RXzbrq3Db
QR2cEHoCd5exsVxhw1XrHHEryeWC7/2O9rikzQLGgmMjIQQc9hC2qbBh6nMtqWBaTfyQtdFyXn0a
ewXsbDYVX/8kr4BhiJGre4RLS9gj/xuCqF8HylIMItO/RAHm/zE0HSGHsgV/QXEEpnLRUJrAoM1a
JCsBqbeh+qOMYr+uVLfFNI4Ql4tuRKpm+96oc41jqVI5xAn51H1pDVXcE5CrQvnzrbGYgSZfJXCN
EUFoEIa2Zir9Vzzy4+R4Bi+lpN21YGNnaLP6ZXU5vQF7JP910zEVCkh9n7Pz1qEZDLUKrCAjFqJC
YPhPuj+3m5Z6lH/p12iQw6P795sf7in0/lhzaQcoel/8fODxRlkY23w0v5hXMf6VDyELUolIBzrl
ftJAawBB1gETUcAD0UrVMf2yKmiAa8rJIthnhS9BPHccImPXwUh+XtigywII+1aVz4ruWhKEYkxy
M1AgGi21u8o8SlYcDfy4/4oxPQkfDzkN4NvaXCWSV+fiUnSJLAarQ4tSBNwF+qO0OP5paeCY4+/x
gpG7SZnjyOqpnLqeRjvGOHSqcxCaBcirv9j2CkDIS5RzWUfHmo//AC7y2Zix6SFAfWME4EBEak6L
ehPnqI1ZaUD7ZwUHiW3rZzuuk8kNCWJeNiS8sVev5JNVoDlKlbTl09+g56C+QZQWVzIZfA86yXQj
rGS1rEbQ/hhb4KW3k2hNFLSEnRWKJb5dknrG4dVliJglVJ2xd1IlerRIuHgbqoqY77TsSYxQCSMT
timss0rdZTYBcNKnKfuV/4B6JfKGvEq6VNcQpoc0Po43qx6OQhzHqhTPRs4ECAwzmtHkmxKZzDoB
rBn0G+Wo7A0zLhDGUOTM/z9tTjJFrrDLOhfTiyDEL3m8R4ZgUKjmrYENjbzgsaxmf1HrP3Ir8P4o
3M07Mi9zhpdwsHmrs4OH56xCkyN9mDIT61i+9aBW9w962bSrgbq5tyMAoSRiyy819V0J3AcXTv0D
Im8Zl1Mm9GTLSvArPpTPwgoxfmfA0e4rJL8IafoS4EZS/pWnhYU/FlhN6nnVlyOf80/xUPFpOEnl
mfMDV+bs9JVo5lezcJ3KER+2GbfgEEGBMFbKPkjLPBmEcOthTqpyl90P2SipGnSfxuR7CnMNl9tB
Z6Jhn+Ldgvsp3zQkF5qWWjC4tFtEsYQ6WuOugWIAh8o6rZjlrO9iXcxA+A0tOH5kfOLrsEWsRtPj
v7ItQf1IZeyUS581AEWrV5+2jkM1HLjDk9ARLUB+82xkfItd6TQGzw5rgjYS2tbqAPliSeucwFn7
9uc9ZAtc/MMcHoixq2KeJt/YEOFtdNjO1nfqMqc7KGO/AMhRbN4g4whRH/3XRPD7pGsphrcNEKvA
qgz+VZxoztULb0BsS/2AzUGoH5pCtbyfkC7I8+BoBsuMcfvZMSsWYOuHilWzCl6HS76wNexKkEJo
B8pNwpLVzRpyeqznrb5PUpzPBCNjaMsI4przcftuTvisqst1rfzX55WM55pufzueMTVswq0sX6nz
ppeLZFiNScUeg1wOKZJSvFsAXwny8TSivwPm/wGPSoSIrRMqdvvkfMOQDVk5qCk5fzYTqdizYc7n
ikrHH2cTQhdrJy4kmNmhUf892Vr6bPdtvLU8SdrEB6KBsU4uZygAFMr+EPrgGxYz0ks6KKQ5SMwG
XRSTmlJpuYuL4boTH5nUOVNWpHpaWDlSApmTbOw/73K89mPKI15ImRoCQf/zj4o0bjjVsnBaoqQ2
vcujoUyAvFCrMMlpmkWcjBmC/GUMmky/2UFu3YtNJDAtoD2wigycMVHg1kaw3yX8eqs19kC+H9KJ
SfhbFIdnlhnxT3NPEq5sESnigcoRS9KmXYwGUTK6RAVjGEdte2nNK2i/WsXKfY9BrLtMC9m/ukWP
auxP2zAA+/FWkOQGQM+gFpw1MT/TuVZ9db/wTOYRmuvlEg5ZEJLBTNiamwWW29lj9Ps1LNOtiAwW
UDtKnkBJdkq4AmazgbWzP5gcgtDzFrTS6dzHd+o0qDc4G2VcnNLMofFO5bKDWm6Mt1m9ls7ZqZCY
Xqfwpzoeyo3KuSq2ppszNdGyWO74+5U2k8fzcqCmbyPpbRZoeuuDjInqjJMusMruHTKCw/bVwUG5
cGaAxw0AhhJx5QJNww2e8wtgjPeswtwQs0KwRS9m8YSSAY11XIqR3CZkASZktputWzQRFDeWZ6cM
0wtsIESE1F43r7KMrWwLt6rtP8yb/jjCBJP60hgXLbnPOd47uj4CbGwvl6GzpQ+DjFRDj3GsTU+d
emYiJE4Czy16dDFYbTPJwFWhirfxefC85DzayfWL97U6D2pSk6MSlNkdZxhOtwd0jLvUP5pqeUap
e+wo0AiwT8U9sOqZsVo15zjYncxkDm9G6Xv3WuDFyNoAGnSmOsN4hPUwJZnDZ2nzthMUPjqF2jRu
ZhvUgeT+rxiaZxaIwLvFkg92X/oUL6w1DmUtrsBAoPiGtvCcHjG7OjldsskbC6uPCAMtpp6SgDwV
ec6FZ5S1s1wSQv86oBksHjLwXlUrb5A3kFwntGNOLyLTp+++H5dVo2JZXnEu42sbb+hEWgYELC6O
W6D2+U4ozurj8BN6cqnGuueQcYkc+ZL+VFto/M7jUxfUqfjkGJMKbYlaEFRebMH2nZKxiMd1pROl
IbSJVEZams96gMLOv74cc7FsRBHd1Qi+XjYKkVGn4Z7jhPqouo2Upyn6oCYkqiUTn93lMeIdviiw
L6GUs+YgobB5l+uHXPImsIk3SjE0TA14E/DbSuY/uigu5t+mERvfNlnUChKZZq6Q1WbMVSRf8qKx
W4O3wjTZKwfX/L3nOOo14ZJBb+b8SzSWZfT56pP9afgzSc4VeMjEuHwhH8PHFcOqEIbAPBj50zmr
eNoZ8YMMmoKzg2ZC2/WPAsm1SPutImVjK0cyh4i6OWIWhfhA/VzGa101AGQSjOv3lT9u/HUgAAT7
+FI9iVGhCWDhFihK/NMUC7NhO+ikRiBVRd2nwBi08yyeZFHFkz8h+LVXmd3IgTzlvYs2i14Mq7pP
7uW0Lni2g2ybYnhEz0Iz5yNdxeJU5U1vnHqD4SdG6OpM5OIoCaAgTff4+VtVGqRB2+VPM8hhKVir
HnltxX2FvbhrbWAUdrBYgr+WZMTWmpXmKH9hmhITbIxM/KFmw9yNkzNYL5Il32krvIS2ey5mXQs3
3Ezn6lAPB8BPjovUgYSqtnB1BlXgaqyKSqK2ClIHXwh71T5PtjWnAqIg30EREKqJ73y1dGEkb/7c
PfkXgAhcUY3ucP8i+bErdkiuFq7TigUxwA2MlzFgTvmyxC+ntMriDtQfZq8FtJ1YpiuxP1HmAZ8q
kLX1KHAyfium791eGwUfKzCW/Yid/gAg0qFzVpCqTXjpJZn8Res2T9q4Y7htaN0hNJxaFUFFLwdJ
ntHGpsaosYeTYStSCBvxSfDWUoPqzu4RyQK8nGTeAPXAMoS5J5k3UXsD0BUnQZ/BKxxG1motE17J
2iwRbOkJsRJqoamdVKvF/h8wC+PUqZ61mgNBLtsIbijwBlol91VvnEQyIjW8hqpS8DT6buhssJo7
XW0dP5I2pIOuAeyfEINPJaVDMtoKJjGws7hLzLTihrOxL1gpCzMvFNyGIP95IlylppmBhh92yG1n
WePARxMourWyjAVW3/+UQIsaGXjPgSVJbmJNxNx7BRzg2wd86yyfjyH9Flx6W+A44dziLGhUumqZ
XFuaERFFWZQA6SuAXhH9BCNdGbW3VS+Vn3oBGPJPUdoQiWsyplyuuVQi5PK8cf7f6kmGVoV2B1+u
iwmegCDdg0S3kv63SdpZylGtbuCNDSoQwW0JJa4Ku5tyTWDWTU2ArGNAPaT/A496c6jGN/p50a0W
Nk5RNCMEqUiFBNW448Ejh0No8HWapJbeYZjvy6qX5MPv9ngl8JVm+WV9uDb+4xI5yYB6jyFd4UzH
0nBNOnh8nEkJVLJFFcONB4XZy+7aqy0NFX+JmIy0jMXHDDa62egQ0F2AgSQreReoY45a5841+ZoW
FHV2rPIwOJmMOQgLzi4aDFXpCTiPU9zMEiQYNsB4n68xJDoTKJe+aS08CyJ9HWIw1BcBUF185Ykf
2WDwcROw9+wbtJct0nZm2s7DxBgkq9vaFNIhQp2xjsYQBJLRda3X1obBPoitTiixTndAqfDF8hvE
QLTXfbVadzEovQDFUYG+BtEsoxnRVbrhpTf2C7eFbUuaaQiTB71YRC2Arl6dCQBJjb6Uj3M4Xn7e
sBRuuYW0dctBXXwReRbdvw2v0roLgaW/6K7MpGILhfj/z6nkvOv+v3JCN+YZjo/xqoXQ41H9QOMR
YzYH2hsrYtMrZ6Idxh0zlRqFTcMAp1INgDmKIEJKF8kn5/uwQAa8mfmUUkCDHywaHJwkb/ACnsKV
RTVDKuV52UHDP3VvdSasu3NgOOGCUMPgd//grX60YhjxyHNHMqpAx/559cSxro9ZVVKotFpo7Tgd
Wq5n/7fV/9t5/7U2J0qSv6rCZ30ebnRsitPxywUhCRj1hesNAcpRs6Hf1l4FWN4GwadTyX5bNn5k
ClSF1d9MJO6b6TKS/loDZUnN1J7s10FwJmZ3yzcaSXFD+PxJiVzYDOXsIuWImslY8FvuD5M/Ya/K
pfsX7mX10fRXQ5LwbAlvDK/DLshHExkLiEeejqlNHqj2uoSSf6+9U7UQ1BXCt4ET2K2Sg/MOs5TO
HL1AkBY+EJjawKhBEN19w8gX9NbjS3Pi/QIYrIFuBDTCzCthgdi9StZjIskot4LhQ3G3lBmT0r2B
01iI+WDPjZ3mG9P5GUOzpU80dqbSA5TAu+vpaaI3M7vVHmUbrB0ZkT0IwFh2zGj+/2iaIVaFV2i1
yEMco0e/N/8dHx4HwJTS/h0RzTKqZbhprjM3vNT6F0bTm/yXgknu3VuB+8NvBDTKgVEDDAduYHKs
0Dc1PZ9NdCEKDdLJj2L4F5gLAeO7fL9LizkuNQ1iG93zd0Gpsg70/fK3y7srjJl309nDz6i5XoHP
IZIe8nyuhFn5cqY5T7snp6SDL6xrDU+DX+/w5xBJXT9at84xXP/4qRjgvuw3NTGiP97LE7/q6Pto
TrdI61UFdRmEtu0FU5ekF1c7N3eDTdQacqnrlmZvzG7z5zXd0pGydf9jxUwGKOng5LCO6RhXOeyd
bBvj8Wt3DJWnDmGNutjKq0zKQsrq0L+dNcSAG7JQHRN18LzNUbvnt3W3XOVHptcmCReRm8bCezJN
bDhKpyIWaSoBQdExWWds1Zz6OSlahXbL2Aly2Zw9w5hmp2Dzt+L9Jb5uI+jiYSQRS04TXq4/DdNH
7idhTZelKHhsBDbdiwIkcKmDP+UEDrtHBroyzzYAJ3sDpRPDEBS+fQF4JXiEy4ESkzV7tiQNLVLM
sW5eoNhROl0xW7CTDdGskbnoajAyM6aW0qjmmu0K/C9oCXMm/zUA+FcGigyV7zo1mKDcIXCqP9Gg
sjKWo5IrCoYNdyfcqsKClSEgxqlQXPejA9wkaT+rUbcUqrBCLMcGPU4ONB/XtMbi0R99QlKt8Uba
AmReF8K0AGPO6wIOHvYu5oCqBLEXLSs7pDaZKQTBTtFSbllAJ/e6fdyroVpkBjodkpw+mn/pBUZS
qaXbwG5aL5JUrBxmV0u61reCLvepnMScRCoeh9R3sJChzErqtlCJMfgWQ4mPfGXCszntikC3MfkG
UgGWXEBb0o1JskMaRrhfqdomR+YfDd2f8LdNcH7CkPuDssl0ISnfXV9WlbOADM1n/PSljE54e9g0
dKJ1RsYiRa1g2vZhe6UqzXXuHDTFoxCwIfZwGHEqMvJa3lhVuw5n7bo24yXltnNPiKakGE5CuTDZ
ZruWJqHH4ollRMSrrrN+tz+mUsTuSdBhxMEc+1GJNUb3f8oyDrp0rrAVjJLTnIhqEJu7OxeW4Vux
BeOOmW1On4To+iY7Vj9lLfTOlYJVLnkbYsyx4+vlkBSRaMWsWT2taCR0bml40p9IZ2AEBPItJwpv
quQ5id/id/jQMfGikGRQp8qM8+lkAwkEZy0fHk0/QNZr/trfnEExIf4AaopKvlcymB3MXulG4T6O
DOF3Ie51lZp7OEpOXMHUd3uJc5pTv9PG8OOxImMCVVicM3nHyu0Och5indMUkIGnUVTLNE7vJZiA
i9cWLzZJw+axFDpzStTePmnLqkCFmWirhZ0WEHnZ0OA5JL01RG0bFtpZ3iYr1nWx9STy5sAq65TN
TOE9BKgNrbOEGuhPJAkUJwmfJOFCUwVRPCOqKb+cf+6bTSr+kmip7Kz+ep3M0sZpUBLZg2NdQdt1
wAYVfzLXYan9tWKMaFG5c1MspLMot1qyZddc/JOf49XIRQi1yCC8c0EqbaUSsnaNLqyub2RS4GoG
JT66QVD3z0jA61RMhf6DXJXSOKhNYtb5tYsrUkLR0DY0wrYuSbyh0n9a1MmIxUOxBtBUOmdUvRu8
E2Eqao3+mLVjm40qeVHd8ameDxYaVa/ZX1f7PX8uLUkbnaBSPem5Cpsy3RQPFL8Mb4uvUIyDIj09
CVEr1ZmT1qrewBTXKx5UPzPjzEAJ1HCL4IREW/TsrA1L5zfLHoeGKslz9qlFry0cERa2f9xIsZXd
dz+ANWZ1p0ViPaS/FRHF905LOBxop8o3f6HdkynX4zJYcJHCiIhnyzdQb4LPAgdrFgRlrEiiHoiT
0jHazh+QSnjMrdvWOZQLCBSQWX/Pjhlfgzqqm5pIGP3tk1Yhl7VayGhpgP/umMJ+n7RJtx4vvn8U
RZoGG42GcogNRG+BzGMx4IGiB/AiIByG4BEC90yjaUPmGFxedYcJ3KDCZ9cuowfDeEVY8klXR/X5
ohzyxwzVAZCj26a9n6MfKHhc/bbkPDi9U6+HtyMeck7hUv8ZX5CSO9xRPXh59qODWbGZ+J0vcoiW
3qi28pTRUN1i9RQEJWousvTZwEJaVdSZf86Bks6KwMZEjV9CWShaDUAk5euMB30c/X1E240slxvd
GcKpb6AnNIZhBlSU3F8slUbRo12TLwovsduKImRhOb0EX/I/cf1ZnstVRywY34GYZemG5dZNKjRa
w/9Xk1V3/JWwlKuHVqRXHvdIBOi6ikCO4GSy4uouLmESpM0l6RUujr4cI1kYlprwDmW3dcym2aGv
Tq2xhgZ6C6XBAzZtZWUQ1vcH1L+5Ygz1hrEVYs21ip5u1YfAuKauctrG6BiAZyz9RCiHE7Lahq0s
b0hsE3S25kozgtvh982aVFiL+gfbTtGTb/kM+rTToBR3leGnR7bLMlBnyh3lvChhOcZonwSJCuXW
jj+1Fr+/1gIjifrFnD1EzJ8/C8h12BhG+LnNCmalM3TS59LpKZYVspBvsWJu9pScpaFNncGBywam
/PS7gYmQYGB8hWoNXRbCL0Ea6VyyE6Xvs1UO0ilycJp7Go0EazFlAIGIDzL6eF8J+6CkHNrAl3Ei
x8Kf9IrpBTsSSNsr56RQL7ndu1eiuKqYezWXpTWrVBRd6I73zGGGFuNq0TLoWfGR6dS4AJcZvkqR
8dUh6zsAvsLoe+aJF0Jl+xqFDgcR8M1tcpqmTdIIcfmuhHmXcG1VH9GK7fXLVLKLBbiNVF2Wjb+g
BH8Qf4vnDdZPJc5ahNqzv6EitIi1nQ7vRTwFJaRpoXBKa+rqfKFIRLiuwTDnxnFuopQu+swrxhR5
WyLVzMZAWwZtBz0BqhzV5wXHqR3aKv8Iysc9Nc0czrvREIixVBnHeWA0MGt9C9czBCspkXfSJH49
5iU0Xpy0jIw0ayO4O0lguQgXrfyxIWjPGFS1p1oqO9Zxifu8/t08ZsdpxJOgD4KmL5Ub/XQXYXMS
Cr43gqqp/WhjRiMFhDfMIxX0IL5LXAnHuMeokd2WIoxuXPVsR+eP5ZG/h3KMadeYXFFVsPFrOXza
oexvW/BDC66rTPpT3C9fZFQCL7L9kt0/vXc5ZAwbEtgTTf4bggo7wv9NUVXNODhn1c08hj6g5Efx
/mniSvTE6UVogATGx+LsDWU7B4oLyw0sp3jX8+abXBkkq5YyYtBTwJmRYRROzftakpCEoNfKZYvY
ahktfYH+mUROV59mCUGOrMAR0sIoKiCJ+bASXeywFe47zgi2T46rK3AiPd6Ul9m1ppiRrx3wpukO
XpIZTsxVn5Hf0Pzaqdj7PgJm0hYXWr+x6aXPJfwRZ5U4l8TddVXcaPKcD2r6fdjjRzUPEsV3KdHB
vv2EUvkUHhVPMIf88yDL6PuXDm0aJlTowfnVZcIBFkxhDhRG3WBPSZH5Cvzu2Y/PmkTgFrecvS9I
9PP4CWF2PowDk5vr7Madt6L8dW77vci0CyqB+tIczKIFTsx1eVmhuUg/ODZOnAlb/ugq/pw3jn18
MDPT8pfAj3A7D/JbKP7d5I41qBFkdCr/XUjZ2w9s3DCqA/EyXuTcSRItIOv2KJE/FgUXzmNcF3HW
cEMzKdbl1QBXmVtgTy591f4RLTIE/OoxXdGYQ5EvpvCnENRdy1Y71YLLLBPaesy3vHYVqDqw4IbA
2XwDEEl5TCvM7uFuqAkzwY+aTrKuovCeFD8KmVT4LMlE4/nf1NQ76P22kZb8dh20EiAaOsRY6N02
MNRe6351n1qM7eJ/pqsRS1xaVnvQMN28C+kaMmjt3eCl/6ZEHxRMjq6yGC5182xXHQIG4OKfIThN
KxFRW5gN1SBC0+52csAOUeFgknqV4/ZTM1WZOL+iVdlzNicuY//9MbNc9H6eUEX42A0cxTNyf/Nc
RRqG3x8xn+DtKYLgS2Rz8LYCHEe+ZG8fgqxkscMNsjvLejL8yMLe5qPwRsB1MF5FuXM9yIAiZkHo
3rC5GiuvNZqKHw5eIkeLrONVNBm+O9HoX2cZ+pOH7cZ+AoiN+apWppqgcvvnnANUgIBZvZFr8D/K
Sq1kZvxjS/Zr8nSjM4IdoND8drCBjUg0YT9yHIhDlJu6g18qIbcaaUWVcCHo8i1nNqJ3B3IJ/ysJ
v5ycW25NOAVANhANZjfMQfZBfqPHdLwSkRFpjIreACEoNVzV3yXtnM4J/98KcZW2lSUlilB89zRE
DsQeFUnvK+lvN9WP6HC+rcwMt5FkpnBbQe0rVbdXcuyF7VW6L63MTvI/6sDunnwWQkdSf0czrNCP
Jhc3nElajzYAn+1PlYgUx6hUE/LMHHtnze2xurkhwQAFUuUJyaPNXbxioQ4RQAYN+qguylOkNzE1
mUClsxsn5cddJulilzmVL0fClf/idrk06C1pIueo5NfZYnKxkzh2kOKRiF1EWhmIhzIkhcIwyNVJ
WN1uTO7sSmwpSk2kwfI1Drmitwk3OWAyNrwWQAvI62nf43HWGqiMJx4GF4DF/DqgJGroIM3uK52t
3xLTnwfaXyMeo1qf4W336OiKBF0GwSbbNCLbU87rQUQBkbmL4QjW3qrnfUCUV0SyflCH4CbpK3Ic
f3meqGLlqUmBDtLHiDWDEA57Z7LfEAw0Sj0UWHeZYzLsWPspVxnAWG6CWZehFJVlW6NFk83YIpfU
uOGLakTblC/9AOl90mHB3D2f+0L5/uwcyJWufmxytkXklyW/k7DL/fTo3cj4dEGaaVAUnbL2A1G9
fsdHTej7q1Wo28R5dHI6YlHf4TFOG8jx2i7hAEAyG4f7L58iq+SBPb3A8bxdjvr1VJCGqf1uCXCZ
nvs06mx89SsgpBSbQDAwSXy778pZ1i5rSHNee2jNwXpJU3rPtN33z1QoxFWGyV7jZcUegB3VLmEf
lr3eAK3TZb9Mz7oh08HprTr3w6r0P/zPvKhN7xvwQhCjC7DU2ECXFKGeJZgbNqTm89oO10c/ZBsi
hETv8F2G4KZsYnKi6+X9QuJ73/gxGqF2li4F/9itLmgDBoSjS0PsTMVlFTdMV1b9LlntptApYO7G
KSKWAbKtBrSH06Kwj+zIdWmLc2dmrATyjjFE48M2HwCqnisawprjtqC2G8e379K/vTRz5WC6MTTc
EHF+7KA+Y/9sLt/xVPEnI5A8tAMhrUVQsj3aY45u58Jqc39vJeBnGdbur+SKflT9ZrZM1sguahbj
5MRPuWsCPtLkIZJFiUFCXlXv8k1Y2z/oByWs4QuQb1kO1EgWyMcxXzP/1mt5lCNizzN/TNrYAqKZ
mI68nCE4WwnX0vjH9ZBPCbzsW+TtK4t67Ip9RD6TRVlosD+DE4+sh3XCiwJQJOCi6o9E842SduKC
ZoNVj04UGdY50o1yZ7clUSpKtYIqoxQOIwbcCPmr0SPbW76s+mnttv0mUpiBs2zpFKWSG3WMhyAd
fajMreaAjb4TXCRJlTy+UMYp7rHJzCZaDuo3/F9rLSmipJgR2/xIjYrQsK5XHnoi0/tHeLlslhfG
xryGz0cJiJkC1FIGk4hCiFpK5pMNHISH8zkv369UH2Lw/NsV9kxKNbE7pFBF9zL9Jb1m/FSg+7pG
KMF90FZTsfEFIWx4r43l+z6WcOdd6kgw1mvDoubcrEbFMeenDXSJXYuRiimQfFiTWWUUTf205v+o
rLVu/GjoTxLQwmWqgaNPZjrfGRdYEM4jTo6O9g50kSRKB3EqyTt0P20+Mx9Q8sAQt4ZtpKLtJrXy
gUMrk4br7DOGKSXdKk4c/QyTPk/okafGk6+SAZJt1Lxd34CEavabqBO4DYwzu9s3n3npBAaMSArl
yDv3ci8rp5NGF2TIJeTYY4EfZmR2kf2Yij5RUxwlYQ6PvS/7Eqbwj0S4aB3Wu2PRL4vFBDQ5VTOT
n3BH/41cngND9EKIKo1hRKQ7eiH8jTgnH5cCFV8amGUlbdeNem5EMiKj5AoV1Tn+PmPZvCAheZok
UnbC2nlAUVVonEQW5yif5GbDacObXwOLhKMIqIXdEQfPSfTzIbmj5NUjsJk2jp+1oa3zEfNzPED3
zzAXjEw+X1961AcBNM2z/Pwc87Qnlu64J86aQjXcIegVH4tUFvTM6aTeEWndXqaSflVeooJ0XZLK
ukHLGI3dMi10GoDZ8Fgx7DVd+6t04VwuQ4NKgvozKfgNFpMnEDNs5RWNfmPb+ynENt9ttFukg6nn
BJoY6y1W6iz3/8w5m2Orz9Lrs+YixFd9QMWFFF6tJAkmWduUH+IFTQGovW+YgeMxpbNLCFwaeZlj
BPqQ1mDsA6vexMFS9ClpCA5F/koQZPERbCrmMgLrxaGmbLTSJYRqP5OJE5/dRZSTVLoL7lTKIQdR
EjEVwOq/dYO+kyhI9BZ4kzAT/8dYPCrHusfff/H6F2vn8p6WKAY/QH1SGro4HPFXyaXBad7QXL8w
GvTGoXykn1S+cy0vHNa1eQfTGZdIWoGFDzuRTIDfGfMYx7H2pOjTBmpY/XVtN8Ci9z2W/DAAHevF
oCEXU8SqO0Y9dpWoOZ+Zh3gmiL7pbUjbDURMdGhw8Lokyft4MQRW8soiQtoSxVAtqyqZe5xcfcB9
gqwv9HPasMY/isewsFSHG5sz0XEBu09JAgniKTOKy/S1Skox2qEIMllGU7of/DHovRgexBx4UP24
3sPpmY+HodcDk0A+w35c3k6W8Tz8C7qHIWTV3wUsKVNzutcBDf2KuoQKCVp71Pq4C5cOV/kCZYv6
WdnZ0EEP6jrHUu/o3VrBLPvSHCvVcGcuvro+AfEOi/g/6UGDv4liTKw3Hf0wTwJqzAuZV6NlSAeM
nWbxcK/Z+nQlbfmv9iDHv3UN0bUjqdK83uULHyqhR2UPIb2+xZVqByHF3bDCJ5tz30/eA3mv7B0w
5C5HUsEhOg1QCY4kElFgl6/lS07wYH+13Xg/CVV0L6OyMdsrrDnb8AqdGeWcGP5SZhdBAsmYS65r
fXmJFcVNPQN7HS346ninTf8MUfxTEpbji3w1DjkQ7L8JJufk8XuoD5++dYgV9l3KYYWHXYxi6Elg
akXOVykwIZl2MhNv3LztW/yZD0gZ9rZ8c8YDlUt1sZiRIhlG3rvbyJE1TSDwMNGrn4fmf20CPeI0
XYm6mCGkyR4nhocjxh/p6qYKdnSvG/puvBTMe6bv12DJSU97xhfqxr9lUQFzUYfUd9DRbkE2M3vb
hDxw65+z3mcyjmEKVkG4jj458N8SKoEiC6Htb76Wgm7KrSWf0xanUUWXqRDF7DG9H/66b7PLsi6q
kDVFRIFMLjfxLlm2IkbIcWbyArtAkIVzwKhHgGKRegMNSyKModuH7FHUXE8duOXLEEenZVhdLcMb
sYIFbsI5eDKctnOn8yIS9ilCPmWdk8bgRcKVfAJ8lqx2p4kogrGUssao4vWH0ivJpWLfaAqQuhpD
uNJfiDjf1xuMjlQOjEQq/fHsfuxuLzvb2h0N1gANsG46TzW126zw5g4+xvrOR8eohvGUZIXOkmU2
OTQ30zTSODLbv458SkNiibFcs9O17xuznFd91L9nSb6xEFbe9yTW6BVBPHBIbB0qe8l4yf4nphWb
5RAKJ7jH+c8aI7NM0KtG3X9lTvSABijxvX32lKDQokASil5WVr1GFiUJ3eMLSN453nhaTPuJ+pSZ
lEh7QDAnQZS0ftBPhbpFYynC/vH/WUEcEbLq+NixW0UbzaHuRnn2ls+j4SZUohyv5BWsdsVqn8td
rFMFhAXhJYFv3Ay//zLtk0kUqhF330WDNE8wmwyhVAkCV7NgHykT9GNKWMdflznM0CNOJGoKfbXS
v6e8Zql0HYuGAJgmy7wahmy8yYbpOrX2E5Kf3AiJ9LOjZ58D0c3AKa5Ou/aifm/HrxpaH8+GtHEf
3PICjehpnSDaFHXQLdbQJ9x/5KtOtVxtbjUsT+RacRHHxOc8Gt90wfCG0omDFNPW6NSymUf6d8vU
LScQqZLsgMBptNgUJJT6tjmDRvmBaF7fNazsXXvptVr7b/SjttqdbSPOGvpYDvab2ZUTD9ruTxmm
IFMb/18xc/LfKMBNa+curtSOvKD4EJ2N6akfRACwV4fAXEmMO8W6ZqwLSn4b8aLpPLuxJ2HtCq3E
Yl7LBmnDBOxe+V3MzPikUPv26L8einMRdwloKp1gbvRlTud8kP0qdjBaVm6MeeoK/9CJ05P3E/TW
w6RIKwkvZGsxih1+3Kc10PoBUWAdoZNjC6lyaumjTZq6Bk8iMlHPxZQWWMbY2WI8R7YtbPX1gNBR
cJzERV8pMnNxJOD4tsjgnQbQ4nZt6rE7NxNk7OSl3qLx9yu4ZU9EB5e8L/wOvBmhZKgqSjaBXSOW
xylWU+Te4ET06zusWWZqj2X6fjOzC38mEGlXkv3hTzC0xXwhL4CWv7rcP8TvTRPOCjJaI2Kuuo8p
iu/cnHC3IA7VICNctzjwJ3PPUOPskgfiekPbZEGMbWKHxHkh2JoPIpbnEFTggAF9El9UclQjSBkX
JR/rghDqXS7AElE80wMr1s3AtRW0BXNfN3b6b8sIy1vkaP5rOgktmYXuULyzcODUGEx2dslDA8P3
LfcNU39tJdVyIHmlX7FmgjzRyAARXrsypYnTsn1R451L+mlbfQ5z3/g3JGRRjHnwJWQVPfHRwrJJ
uP/mtlicsk5YEhPLbienFptJjUfYz8f91GDU55JeFB3VTfj0bTTBESE4pN24p0LcXUdR2iK7iIwN
Z11zMoLO2IfREQBoNYfEegYCQ3pDwHBrqge2yPUycpm7uaB+3WKbi30FAxaspBsZvW1/3m8inc9x
UchpiFKbD49d3pQXnRvg+mr9UuLFJ6+fpSUdFKU/F09RZqeEHwB58NAc9G58waxKbHfHhFE5QVeJ
EMVwE4cxhtlQ5Kgfd2RSWkFLEZHD3VQORq83dXhLnHCfXvav1J698Ar0IBAn1VMJo1dSxmSj1n7U
fTBIIpskIfOl041+npdztjykoR1zTeVRP5ruE2PdhGysecX+MmZNlZZYo8VJDGxx7P2wQFpL5a8Q
1R8YYbbmqmoUWr0F8KbOfeALHpjq1Chr/uTyBGB5C/wtIqzIYpqDY6FXb/Hi3cpiXlDPmuOlXS/m
/dBnrjGlhsr98AFmYF07CTDQKSmx3LL8nWqdnIWht9cJmMjXxYsk4cw10/aJTaSnECHverW7mnoB
gv4dMPG3ynhmpoiPMXSwdlcTvdjtQ0jFm2zjYsc5lCV6gbC08B7eX/RDXzKA68a//C+s2QJW29t8
MYAPz5iu2C3vHqU/m/DCrvRXBJJSajpYXM06VZ59X5O3AuFWBDXJ1WkwYPDHVfUlQO0SsRTpTqDD
PQIs3j301q5l4yKkBL9nOPP8pmHGABqlQxhrsOHGd3pn9mLtviG1UgCs5U0FsGODLWASM5wpZS+8
NnUAoLoRjIxQvX0YZOGTnKIwF7CVemTJED2vuwNE37oUyjQiCPfPD92HSQ75CZawx5VsMvqzSKvl
sy+F6c3vPn1D5duMOx4RUA3gxOqSJ6p9oHQZACbswUQBLLsf/2HENv/ukz4aI4XdX/5lISF0QYBI
mTqJfEKKncSrSn+OlRcmNb2kHwdaj+HbX389IZmlv8eecvXWZgHBaXO5Y8LV39Hc1E9OgoYwzeHP
xDx8L2WxV4e4mdb7KjbjK5vpm3MIwfLt/IDxA3V00j47qUIsZKuIRMkusthskIMKhCVx4Wd9hYbO
ATcMfe+70/SI8BiY/hVer5zBzxLWpKh4sriM3Vrhei+kthxxqRo2cW5nbXOsANYiZTFo3ZJIrvMA
MF7OSvjWbtLqfETvbEC7ZLj0AjvEzhmuzRoJIcbRtsiCkGV2aUxguFuYh+JgTUSLAJsvXSPh/2s7
U3N+YzIxNIhqOXIjZhA3/G/keLygodV353AdWrl4CWaMHraXsxyzDOFVpmop6st7ePu/SQx9OgWm
kov3JG8bb+NaizT697cyUC0GsqV1J4rlee8kexuCnvoXeUTzFfPRWFvUW85HzZr3DtS7nNmaZXna
xDuibU6/m+Or26rpfR5zE9GuEC9AlAyfbmEYQzlIG96ZfKEEHPUzESf2PWtkGCGd5PMINbH42iYJ
BupISAGgDOKjIzkXo9E1RCpRdQeg3xcRNh8FlLZu47oCss+YZ7ZpuvXk+nwnj083SizhYcQJbjbp
Qy4TF+IpAzLW2cS+gyiGq2Xf+HnmohplgX3lyaHCzgJWNRB5+ZKXFlfurlCws1lUyUPe7arX86JR
+L6Vm1cTBVcehXYXuuj9x6hnBSsTG9Mtgl82bbgT1csZuTaRdRBYnAT2ybBOgpwoi16pPu6n3EmX
1Wz2/tdhctXu9ln6sESzn3m4CZQZHqSbD1BJ09WfZQ4qmqfe0PPrCfYBMdBR517irVlAVeOWJNP/
yJ1dhRtA/9qCPhFc+L4/VPRZBDd3YIgwky7nJXqSNcR8U/gSnGqgCAH1a//1hm7ME3auI6c0BPzw
i9lXZj31DVQFhYj2X5iX7J6UpdTeJu8Mxw489vHMt0+VYyEhoZ2DOYuK2u/zK6cGdB5P9xvO3y5i
4KKgLS55w6N7BqaKNkpoFX7NqpVAubV8fsRb06z+LAUB+r9Gy7KBZGhJSLKbor3aBCi/yCnLX4lk
WUW+iQtKgpF2Wdr/HLx2cCBSCgGRL2xUmMFNafmLo/sNbWgrkGL09AwbdySKKsGKYojoeEi+t8Px
I9kUSHQJCUEneJWWTraUYIwOxLyLen5vm3VMJDJmFqR6ormFnfgXs0/30hLnnvmRJLUX7M3YypPx
boFZYsLR4k7fsXnB6Q5Sfq2F3f+1DORxBnnyBvcjZ0fpQgyuKXJpcwds3QRvRd+/b+JbnwS7vHgY
PqVwHx0hFzokasAtJX0QVYyvGK6DpKRfXUhkyYqb27C4NMUzYN8US2Ryj7YPbsBwK+bGIDzvFg0s
FTG9EOd8eTM4b0Ui4yEE3xS3/nRbBsoCdBF4szEZhF3QWZE5g0bviXGoTU1egc2FqVvwScIqrczQ
hiQGHTAR5lRKqqTdBqwMRFM4HMEo4y5U2jv9V8LlzdeACDZVoTuvcmU8wIbBGBZZTxDezsmA/z+j
IFcAuAtENcU838m0HHbQtCXIqLH6TJ+M8HiXvpj2iVIwuFY18LylkoKpU4BKeAm0O0C/M09EzVsq
4mB75rCgFWCF2wRz3PtcDV3RXuI5qMWDSFP7QYUIQeHBQgUPw7Sw5r6NSv/kxxM1FKh0BSI53C9Q
HQvLGejRlOUX8KcDWckqI44N/6XhbET0Fy75yd4RWuPNaU4wdbY6Amm/l4i9xEh4hXrN/S0E6pHQ
KHrwQaMNlZj/OVETe5/qccya4PJho8hivBAq771U7pjl9qc0BUUR5JssMkymKmka2HtI/vSh5aNm
FHNTRUF/sFsPVfRLz5OlzqcpbVjKxkA57bIMKi7ljn2Acb3sZsrD6vGaYmU9d4fNNvcP8fcRACl/
299pt1zEWpxG1lAtxFxNxZrt2UFmsHOTXTbUGbrxytqlBHNs9gC8ve3ToMKphBAWRLBX3OJt1oat
6BqIz+YIYoaRjVT4LLb+pF3rl9ENFKryUkJKgSPUlLH1c8u0CYS36zsTtvkesv47b1BeFg8FDAQ5
w7FoN79SQIkJbCj9X7j/zNzXifycESMphns9w+BLgkq9UbG8cLgyAA+QPYu08YjpGCP5gj20kbCm
2c3QxsD3ImwjF/LXnw5GwY8ghog6iDcCATsT3qeDQ+ZiE506j9uvksOFTkpElgy5mTTGPhTKdiau
C9Jg2OVV2HSI5UuLbNGwEnnnbkwk8HWc1PkjMT6lpdIMgqLBQ9DTg4tkU1Gp5U9CMFiNRMg0WXbW
v8DC74dwjKwLLXE+Akg7565qM9BczCnzObM0w5oBDlh6NNjRUmTC6wUM7UtqXv0ZvE4nLSvH2/+8
/R0KQB8GBLBMOoUPdnxoQ/QmfP1he77wiz5h/M0F4FM1S/SMolefo3xaYR/FPlFb0O8twZn1Nn8D
j3B/K0wRsiKW6DQ/op+K6IBGLoB6H8MvYcCY6EZLv2eSNyr/tpzAmuUHfrK+3hHXP+MwnWh3DL+z
U0KN5KEvMQOpX22nLE9DZIrdSHQ9FR/TusNDymoizAoa1ym2wrQ4PgcUr6DvTYW5elXB8gonV3V4
qJdVlU1rITrIW6E3JYnO+d4niU5w/Oiw95XW397DVWhkwpCp0c3z8gJYg4kGBaHUTemrQstnhDmW
lAyWdorid+WhiGBH0ytlUtMNXSMn7QHTzZ4JIfr4MGbgBHSGM7F919YtM3EZkomvlEjQoKfO+s+Z
SESINQr0w3lz6nJdE10+cUmBjo11dj73eQPjUNgTPup3NGlTLY/Tcvl4lIXDi2H6Kbf/TFd2IYly
O+VqiF940PdFmULpdlUrsbpu2SDrAwqTIptXjrzm8LBmgAaAYPk+fxfQSMxfkULZ6XS1ntx+YIgm
MHqMH3N77h9A0HSTD2Uqw4L8aC0IHJB8ep3RvogpBFyV9xyQ1CYJQVdsssYv9jyCOa0Hn4es4u7q
WVslMdPI7fM97dbjVu0DNtIav9RmT8H6z+t3B+t8wAT4tAzhacBBTXYqRgpIdV9CuBJTZys05WpW
K3LJ+78izbmeZ8tEnqN4VFbPlpkgp3+HqorJhY10zyiMcJga645uNQRQx86hzJvdj5JZbNBdlB3P
YXFltFpsu0eBWZJkpFXzl4D/6wceNOEQyvXVN4Ko9g+ehNJvSwTq8/gaXMgqP9jGJ52mVS5/efHi
DTA2bzQeScW4usYIif6NhNqpJsDkL/MmqytEC/MXokE/im7Mtt9zCT8YA0JTUE5lKu1vmHDRA9ZV
9KnzVCPI0so5ve4V6eGrgTlkcEemiuSlngBJOmwq+ThoZ5v7VofuzpsijiyLe5l96NjNyOcRjl1P
ugW85pN5HRUsTy1QniHYJQ4J3+To++xfUWJbT/bqhSgEY8lHJd5CEtxExovFqFDBaE3HqKpv0XX5
qG4Ws0XKCulSSeuJbgkjxzMWnjll+r+kQxZZKLq8CtqPtb0+a/qHI3wWpy3fiBagPtfsqOLVfzNU
7ln2+GPWaAtpjwh7MBfICEPmKChm4YCio82mhgt8fh26xOXxpiiM/kocuP1r7nzKkIUl2yuUXRWG
g3fcO49HT52aP6Axj817jCm0t9DMBWl4tUl3CffZ4lfBdh6VzoiLAfF5Lm0p7yfmgm84wRNLBeoC
u8HEAUpe5+oU5RMlStz1tsbPRq3eVC/wCNgw1dNyMBXM/jnJWk1AO1r6YxNbAuaK7lxH3+AJoTkw
F0H33pm+XBvCUe03d2x290qXNGsY2RD1fVwR6i2o0f3pbBBpcs7Ztq2A9Y92gMLIEGjXFBnLEiak
1wzVo/Vcvy4vD1Wow6dJVIHgJTbVKCeH8hknnOZFucHNeczzmhsiLEbU3zDMGQx2JncbEynU/2ZH
pL4GBgcF6FZQql/LXT3QwM2Dw2UBDAw4FR9aajZX+7E29qSQBtI64/o87fyBIxgwikJ6HnoUOQbW
68md7040xgw2uC/H4Yc/Lll6o8V17nXIP8ZASu5I7m4BuDKLJoPtEs8QYWwtEkHsegRO5/Mn3og4
o6pPUXQWvmoaGI4lMxgbr8o+i0fwNhgTj6yKNNF6VXk1PBJXpkPz3ST/i6wM4pHXfgNEJXvWbsXm
ulwycvjn5CSj+b213wKpAVq6Dcvge1vp33GyshZQuc0AnzaORhhx3js/NNOuyLL15ELFlNYxCD3s
dp1Kc0QKM/xhtc00uKQPp/EJA0R9BcoJ6tKo6Jtbx2o9c8JYUui7yGi1UkJEvkuVki7W7b21Nel/
/nHAu9zO/rzevnodPRtvoQ8RwilEObCwl9G7quOCFJ1E8KvZCe6MFb80f/Lpvz7SRz4UoTVmOzoh
KxLJEsQirln14jOC1Oh8KJVJB+dAXK/vN8BrG3LmjW1HpiiSpZb7rmACfDrSe79/IZg4BKSHQVWG
yZbHQH9ttnruWOAVtzO/voCk3fyurezVIlyPnQ97ypJjEetj3zt6oEFZQ1u/68mcJrFVxZQlsY6d
4xA8GWdSKm2O6BJRZRA+zAX88Kg5vgDar9h02hcvO9h8MlvTEe0RckRlS4eRlhClmtUb9eAYTZrf
C54IoX6HN3A4pPIoW4clNdnbqnIfiUIlDHTHZYsc5es9wzkdPa7Y6hqWK2pC2B+YpS1m43w9qwQu
QOvnU5E0NlFBRhcBBEyIM+f8aH0dMXdjUzyZQKtxuCD9/wNg4ge3MbVkjHCG6+eppQNgHoRdnaNx
ZzqL5dahMPPOwp7WEjcJtv54iHRmqWMdLBYE7SrgOGGL8KfXTy7MzBTh6YTIyKcTzMUMGc7nJqop
1b1etqWJ/CP4LrSTCXtcEy3J7TZiiOSGkJ2KklbB2M4r64MGvyfwSWe4eG8hVCKWouN/Ch8mlxB2
AXJFh35eKwGxK5wZNOg1prNQPe/I6MnWCvIyC6nnBIAT1DuIIv3qKWXKjrFDkj+i//Dmjfd+WdV1
ReSqaVHZObX2t1ubaex6VvFh4iNNDYoiGkdLxqS1bhclO5BJsXQnC71HbOwcyso1NFFX6TjAeHRq
PqlPiDTjqSK9GlTA6wD0UDfeDl91ovnB+7Xz15tUahDhKAF3p5BmYge94CFCx4gpLLj7JtD1r6z9
fqijdsiKZIGBb5xSbk7osYOBNipcFfCUvigHMS9Pw47o2z+rgkge+R6YwwSbFPqEKVhQHrb5nAxo
Qjz4PyzUkEUpaayC6M2GYJR+OFWpXJH+OdzX0qcH7okTMVLH3yAw99mtj17ELKQsJdQrkPUOoc81
KPuQDD/XinMeKMYX0tNGa0mzKdBt/penwTcayi2Bzk6PJ/Oof8Q+F9s+Sp6C0UG2U2l78/7A8Waq
tC8M+fsQnmdsDnDacyQh9YIyGCzq0G6V5jWHhLBxme6SuTtyRdDnOomZZWTSKVBuKqCB+Hy8cb2R
ZoMPaiF/sAU8oTEbBGWYbnxEepMVeGc0kqv/gvghjgnsaOLJCdVfF0ra8PH0T1eC+G3Qi1mX+G9m
ap7mf4H4etFpZcJ77eYrO8DGjtzjZrsrqBkmWcIg63FqKtfpYa1KkMQ7v7NmXVoPyShAyIhvo7PM
wVa8929SNgwAhZHPN/I+FlOt7XtZ5V6tkDRdh00hi8LI1AmIkYTDRbngv2qYspYXAVBQp9TXBU+0
/Q2gcfHRAAHpMBhW13iYJdbP06TuFM0+KYr/Hl8QKdspmZ0iKzGbA3BWTvcaxT4r+aWzqHh375fp
2TdFI5y18w3dfWiv1kWE7Xlgk3QOWyZ8aanSIxR9o6vbb5eEsgQyxPXOKoV2ljURstnGLCu6GiTW
oFu6JuifZKQvMXx891sMQyghbKIIWoFUz3Js419nlfVL9RfaNfisGL4MrCk8E3SSNb3QAbQDvz/W
OdWE6geIZHkPk4aJgLLpigKutAL6qbMOhNgPuyGT9k4+TZzban4hYBqEEpGiSaE9ot3N/hpb2r3s
hQI3RU7zO92TksDk3RPvyurZKuFYBVYYCQ2sxGMNrOiZ44iRRck/d60RQiaOyxxQ24crfvfCkkdm
4ozeytsg9jjyx3kWE6EF8x0SNg4vdcBpBlmCFmsLfpa4HhpHT1NHodRqKmk4hGAQO5YgDrbOgNo6
w7my9I+92+8SyJFEihDfkfDoljVjQeQ9SxU3U0l5N2RnceIOmsXANdrHXoam7xZUP/YjTAKCOxyB
U896QhIpqZC0InAteXtKj31YS8R+oRNYhgtwvnAcLg/EQ79pDuwYx72wjjdaXKHy684BDTPNXim4
MQP/LsAz4fgqQ4nRYwbOWw8WR6H5c1R0b4n04VPPQb5BT/goql5ERDcmV6x17PKtLxn5Xk+eN3S1
mDLwkAjH/UsI4ZVo8pzr06ffzVJnvL6ExKEHdUwiUb6ByjtOnB4iUD/MRtKmdOB5eqCxMxKvjZ4H
PlCGtQ0dpElLJ9CBdaunlmOcdlKMmQptXNzUEtE01pZaqMxDNIok9sf4hsF3i+OMGTxmfH+tjFhU
3/UhV6UvVctxlJfrBtY9N21C/IMEDBdZ3r4bSZYGHuEpIS8FEl3p+Fh/AezkmcuBISRqP8GqgOl2
LcErqZ+rAhEG58U09jJ8lKzR/Swi/+AlMKDwUscijxQm+p0Y/iO/GHQLHwnrArS4Di9kGhGxet4Y
jmJ8UNAFCuOUhrX+hiV6+/LLmKH82c9mMVYsVE2vUAmdUvFdCIrAB2PEqqhQ8sAlsPxQK65QTJKh
5+eX0eGjdvPYwXKQGe8h3NrrCWURL3Lsy10tCxBPwOCDAEp9vxzRDa/VJalVBcbIWuWm2NuPJpn2
8UG4T8vnDJChIbmsyrR4wBGZDGE+IqlBPxEIAezKbJKQaXHFbXCrzS2jPoRmUoYVT0a5L/4c12rU
oaOxxUZrr1Gei8bjbbvHaMb9cyxklSrWDBXsfUAZxeBjdTIX4X54Z1hhYxgGcUWt7kwuGni6/Lw7
w3FTU6skg2RPcgsI2bbNh/n54zlwf54cjaFpc9MPn1dgS1wmF3m74hsOhB4um6dRkzRmSSOkScND
p3cDXMsW4LX6HKg6WB8dvep9aF+lgaX0BS10ZzuKOaKb3hDHT2csQFAZqbvrdupjf1AznbqC9sJ0
U3oEFkR6FW96Ln+vtlI5xRj2mosELkmmi3pbMJvF0dKVd2IQuLnZ+fvOgOMhFdAaHlmCwUEvy8dX
rex4LnP61Xk/xScqRAEm52LO/ZmS776tXO/jZlmnD4fHzKuavxtfW5ZI8sctwTh4Iv6diCnqRU8l
V6hsuGF88BQ1lPZ1gcQZOJvVQ97s8KeTHhL+C/5MPvTV9tXIgDOoeCOCAy3go4MyLE4qwpoR9H/G
LIlxklMI+kLDo82/JKtaW9wQNFosr7vHdHccVtpgTju16MNlpdXOp0vREA6LX3IMDM3iZfFdj6K5
DX3UNF1C1JWoRkpC0X8MJdoT22hfLmpJD8ruPThk4iTMXM4zCIQ2Zszd6uKQlJr2TZzgtRNQ3spt
67EC06vfNTmLvocAhRHM8Zvt2/9riTOV9zP5K/LhuZffiAoAfB7ayTkeUfFP0tFd55yhjOdtZYDs
GfPx+W1SUNfBOxCbJU6V7XLsCuolu0D66XHrDs+9ab4KdnUyQE5GH9uc1ZkiK0hxQvnrs68MGzOB
Vn9/shUkLykQieGtyayiSKcFic3ia/QLaWLZffGHuvTQJ1YI9fZt3LE3XzfbMIXE3LnJRqzF6Cb7
Zy08xu6DV7E7KweqQp8JjlYRunWmlkK3Bz638TTUjj4cm55eoYwKOzEuvOFgbaO8p0RfN6ks0Kl2
Ikdcm2RzgzdpBGJ7KxO18PLAy95BiWVEg3UqtNoHIFWvtRD23sp3oKoNCki5oZv900EVaooJi7cI
tIkYgIJs4sHcZLuoxheai0EUGeme20bfD2gSldPc/m36/o1a52/5EqD7NMBfc4gPnTCXsYqmzZ0k
29zVkwvqsQvrDj5Cdu6XuM9IbYQua20Swo1NW61Xu3zVChBsKsAaVzelhpQCkuuKxC4rXMmXUEmU
wDkeZy9BScsQg8N2FdWVOhk0fP7JFcZoGA5hGDRULlftwImDHRul2ngOc169VDTL7HlbZiPXmXPr
hlzE+E6rT+ZEXp9k7gcq7ya2lvBm9oAOhh13AO6aA8gPxhq5Hs4EZUCSo8IGTxoLasHSTznuXs2X
Q0ty5eEqNcRmZ9Dop4WMWUBibc0/QcvEwYNkaj4t7rEc+ZufSNv5J3u9kLGw+pjz03wtseA6ToIB
alsGE5bF2FKlZr7GDTTzFb3Yzl904XR7RhO/DIPNTAvaBnTtGOIyBuzMufaDrA3gmGbFiKYGp9YH
wrPST/U3wNXneDfofz/KNpGMdaCBVyRZVPZNdqF0NzySfhjKiUJbJZ7hLGXNF6FiyTb5vnYH6430
vUaFEMXKVBwel6azMFHhXPK53G1N9DDcDlwScXZPTj1R45TohAjkk3eSnVALkHfoXHw7jJVeoAP4
XRypnvm29BR1HeloU7xoxIOKG8W6sV9yRoTmXegCIJ/1IWXG92vsYB/A+0YQIxvd4yk/VfjmFg69
0tZyYMe+MbBosoeP9tmYTChz5e6iZP2cdMz0D3uoH5GJ0GN47eNW73ynL5egY882Axx0Kb9DgWN5
xPXK/iMmnSOYPeS5OK0BxSlZ2m4Xxv2FglEUX8EEIMVGW7ZmncTVwE/cqSlBfkIIC63x2BgXWRGl
i4K5MU5AI4Z2lsuRs4m+i7BW/16tRIr3EbKQYFbf6ahK8bK+41s/y1yhmGJgK3pVIvBkMGYev8pF
Pmpan9fZR6TUEpQJfV8+Ht9zQ1Ugkas0W5A7qx5Z/PMfa9nsVtoJOcYAZL3+Avff4qUzjnInaUIJ
5feaf/ZvGKAfSqOvJYGGrLxc058pWpZE9a7xTg1A4r3zEY6z5TDYVt0w9f7DLcZEYlXA7Fr/8+WD
qy+g/NyzkosC/kQJ/2ukLRT1po81VWLYH4oyxa4SjE1YcNRf4WU4iBIEP2ZwnfiPOV1k1uT6Px0D
vmtn43HuSPbx6/apXTL3DepPd2Dw9s992lj4P2wVw5xs6jeo+CPAiXxAilbUxB5C/Mrq6LXV0Znc
mED0A6VWmdUth0Yl6zffDTB7hWNQhYUGDwD6Nrm8nL5/Da/dwLqoKYqWp2S7tAbVtdNWq9UJXe8T
3JqBEWvNjLO+EPW114riu/DoIvz32qL+vQY4L4IsCKKGagBBT7IzvmSwSHoRW4V61J2HrLYen2bE
pEWNjIG2paFRSlVOuMRVGNJHUSqGzbIQ4BM8qHxm8jr6/+oPeB+daNfOUUwrM5Z7JBkoVjSxSAnD
kswACdS3PX/9J+0zkxE6BLxPY49zqkxc4imU4uyKK65PX2rnfkMmNsF5GxKaLLgpEHtUqBjsa7b+
Jz+jYdlGDDSulz0O6SQVCb5wI8ksQ2VMMX3Opd9MYQI0Ju0caYJxsVGGPBHbOUP36EkrV+TLpTmZ
x06zLCat37kwWXtxuU+JZZZhAsiFzIj9ZYJRbcvaMgmwRoDa0j984jtd/pSkN/aYWBE3S0Av/821
y8Yp5jllznqlcgcjv204V1FjyD1C7GTD5lalv5rk5l35F9cQH8ypSUmIsParsTk+LIJ5B5hi7kmP
lQhT0EWfdXykkVpHNIDzghwLHR8n6SlA42oy8XTO2Hx19qy0U7sRWNeZiA9EeYLonC4tW2apLXkS
nDrd+J543tsPeXBSIYo8HYTo/BqRbtUjWIOGrulLK38EYVFcsAOA9hT4MqM8++TnXQIU3rRyASq0
04hfAw2Cjpxu4sElACA1uzcFoWbNdRjwCvMwxEsMMSsm+HZfL4phR/Txw8Xt3M/Mimwwbfrtf2X3
ultB+iyT5PgYXeiO5se4XXxN/riM0XieZpfLt2DVtalLEzH4SG3t0y26/65jO66eymKvxu6j1pGk
VZ2j8tJoYSDxmYOi+D/uIEvhTbaJei1B+6EJnDx3mvu2mg0srifor4cd4RP6eIIkYLfMUX0HN+El
ALHZBnja4Z87zVoubEX0nrDJHVAXDdZ5Q3Y21sdiYAQLLwj+LqG2A2iSPl+Vuly3G2d0LfZMYsAC
y01qJZbX6W4XvsnmkjWm7nfUySETDRR8zmFXsb9cMTvReEZQXlhNwVNrrYy6fHGwJV2cpOfffkwn
baM1ueO6wfSWOYKRkCkpimTuwc8d1KL8oL7dB4Zpf5ld1fmv7fOokX5Axs1pVOg4jEUMTSUm6Beg
7M135QCpl2AzV+m2dtZ2XfMbt9Q6p5+cBJGlj8/BVro77QPahT85gihOolPYG8VcCe8SxoFDg3NK
iwG++gYrYazUyj7MKkyMb0V94UUCFILcnVJ5Sv5fo/Lnvi2H/NRiHUedI/auV0e2fycy2JcV9Y4A
t35vbx5bKQVrul7SyTZlv6ijhaP3zWiOy8FOxytOKW3AG07iWmqRxRkDKnJTl5YVLJ+L2Pi8kO/s
Pxh5OhcCOBgAc6YBvUsE27gykMbFDD5r9Sr0DBUJlIw22vaVZMndiy4biNfl/hn9+Pe6pWDqO7u5
v/PxMJm0zZGjmgWPXo+HVdf8PKR4nnxVk/03DvSXTuFYhYK81lUg1s3sfWBuOVRSrlXe4RMZKs2B
yHVgv/y9D2i+1gpFWQ6CodpigaGb3IxIUjfkyEIrh6TdS21RsHodD3Iihe8bJCIicUIPa6DKp9zE
8m2YVzvDvN3gNuF8VyUbhjENnleW7NP9mtLabc6EZIKx0BVxCVaF6LpKXD6dNxg5yy21RWjGEZ7G
r5qkFnDk2pKhevUco0a+j8hiprTcTSdw4o1TD6Et4nSXStGAlP+RkOgZs97h7hkwauu6LXsk8Xwl
IQpW4LnUrw/FiLVdnTeYpCorrHohDXxZAWl202kofObNJweLQOa6zElgsk7KrTbhxnQ3fQpGRh35
YplS45/n4M1MTQYYRGYMBUdR4mkO9sL9PDj4IUe6jeJbvNVbr35yNQaEEx+4LX51b2nulEMYSHQ6
XgDZ13dWZulSh2OAbFJybnqSIYt/3FAXaWZp2LRR0mB9Nu2LDU+0LvAZdY7zDTowOUJDDia3RAi3
8YSIjGWGn4vWR7cpW3gRFYOxHBbpi3BLjEmPReJOCspKC8EE0tRcvOxJFHYhxjZfs4oRzw3YDrVJ
HqSszE0OSTdhI15ayISC4iuuNFTafrInM4Gqg1yBr4JfdPG9d8yVvcgNITPU7iRHMbwm8ro3Y7I/
joh+aQ8Jd9pDv7YTNm0btA9ciwN3ZNMzyLZj3CYwd8NcXXuY/NWL+RXDAC780SSXgyuh0ZdRnNKJ
1+llW+uMJ0dz2IP480qqWTI+yLSKgNfXt1UbP5DzrAVrk+k33odq5YAmes6K+q3bwj3JTW3HpcR1
64NH70WHp8hKD32vpdXuqyeMoPkAQ7C9+rC2TBkLtWkKHLiujSB5QdXRP2J+1+A8ctq+1WYvYfpT
Kbnh1KliOVzkBhW9WRZ/Ol4dIZHO76aS1DCMv1h4i0e9eoPhyJxUL1Rps987DBa6aEz67Hogk+2r
vppaSUfLWVQVZbvnz70rfp6pud2ijxte6BIhaIi/y0VP3DAxzKqIz75EsKHMpIzm+UjFFc74dCis
x4F9T5AV0NOXJff2VtmZt6HrHPGA1bu5YGZcByKtApN6QM1cYCZyDwDXOZOU+tJariMticIB9C3C
dV5D4wDOpKNEBPtIa7nOcsnnrMHYHTwAQ7wI4G8ng9V8POO8OatjQpZyp4HNegEbIza9i2zcnKsS
HiKa/Jitku7vj9BK2fByNvMNxFVlKnhT0JhB12T82Rd+j+hxI+iXjyjm/On/Q5roT+fw+Bcn7aln
TL9naYA20v1kyzdAJzwmZQ2T0I+gCmogPT9E/4kXu9t9/NfUrG2UTFNZrvmWYCG4wDsdGg9t+1El
WXM2bsUTLF+pRkL8uH3RjnYvPJ+Nq6ahKVGIz97hFvwdNSwpdguF/T5LLpHRKTt3mEoB2y/tgTYG
6tc/c8rHHBB1+li/GfjS1JHLzV1HIT3eUSCW4H2zekrlPb19uJ6ttUPmMimlys7mRkic2WnfiVlj
9jGPdI9jm5iPkbTd0gaxyqyGWbnhol7iPlQq161uGZyfEql0xGrOngv+r+CsEDHn5Br96ZAh3lQ0
UjdrYqPVKHpIMzCnk/BYh+q4Jtx1ji2zC2P8BvV1JGVylFYLYpaC8oIH4C6kC0/RhmjB5QjpkcUv
GjL8fs+zSafLCkNV9J+UQRFJ+nx98hFIpx8G2str7kGg9beDJUrdrSGOJWiaAmgfzWmrBv66dl7E
AzTxmoyoEubcvTQrrY9vhohz7QKSP361cZkZzORZ9aGOWv1ljR4BeHDMLXZcM1PBAhHbULzxGWxf
fCV6ZXeQ8IJ4MdUtTvec5rZDNoM+iH1J0FB0kIaW/St127uCplIDQ2OPmf6uJTbYXsXRwDRBwGAK
ju9530jPKM2ACiGZ4rvEgsHDKOZ0Sgv58bnPB7f6llwGPhA9W8hT1iCnthErrZPJmfyoHeXH59gp
qU3NFBquSqQ50I+KUMr8WOZoQaK79uwC41pojXncW4m7sAn1impV9+sqy7/NaBajgoujuRQ6zzR2
l+ebwRqJqL78FL2y5EsziSzq9Gm3GYaOQrs8wWbTSOarXP1J6+wOW7Oqw2ykSC7YayIbcaTR6Uza
dY9dyWyWBjvuktUIpv8sAPnYDtPstOdSziisRhLkHPZBYx/ee2y//RHDtH1BRInfbbtyQjTtlLUt
dLhcAt9xr5bI3417aIQzEjEXTDX+tbRebpmTsL/HgPR2NJvLjJqCEm6FAkuZba1Jc0PaqIKQOqFv
QHPFgyVRheX6BhzLB599r2zWOmtaOTY2ZwIdfeX8DK1J1X4+6Q1pyfxtlbx9wpj55fl8g+ouLDls
WOiCS9zVVLz2L4jsVKUwWu+Hz0tYpBv06YqjB2zViLw6Gh8VuzPWr8TSQkEd9Xtbq5Nafst2Jg6c
BWIWHwCkFyiwZ7p+9B0p5adxjDtg5q/N7tNUtJImHXHLduXZt+3JWJON3xuNQZFNtfegKjTRXDnm
RiIkWnYIWh03knjNFDJlB+Im3avupRqR2u4i148IOemlxTKbyfA/1qstSriOU9KL+slErLp2rjRe
cSrwomvJpzdSGbqqKiJ6OdBrymAvXeaUC1HA8Y/3gK+kL78TbngiCDRuzGdMGHAMVsiPQLKh6m+n
LnaqYF/j7XbMIAs8svl0SQ/LISGSYBXq4qA2LtVvbo5oxHQaP3np1Jdw/t5nYxLo6PszwZxjh/G7
AfRomz5us59aaHUGPWw7Tisfw4xongG/LhgXHtYWLV1l1ZdqRLoyOfVzgaHmuy2uWMalkPyuL6Bm
AIFu0X26AY2UVFgNBCsW3BMJgSlzVdDCf3MDcRVCSldkdN4H0TciltI3IY1/EzET9R6FHXopmSAX
vA1cZZY0KIjhIpI3qm2Hlt/4d/KCeP2ZAq9uZmRzfvC0eqzYOszNP43quAnJiJJH7dNno39ks/AG
k347f3fkoAOVhHuOE+yD/UbrJNUuTp4HBr3Ikilv64BuKhcg9rWVx3sYPXA4imoGthR+fn6Xchvd
1yaThLR9NR1B0S6SOCQtz124iIptoahouPKmor3pTG53B/QQMuqlMbn1bXhCWKLguHzgCFlsaJV/
gRn4SrNIU6sLWUpuNiS3jzQrn7TL6R6b/uUkBuSkQ3jq9yiL+SZ/bIApOgKIw9We0cVZrH31chSA
QWCAkpPhpeLkFp1wIZOeKqT1ki9Y65hkf9KAPPtpc8jp+3HUrKRPf5C4XRgkXnsdPTsCgyEhBy1e
0AiJeRONGCM8IKvFRo3KqlLa1WxSe63ihUBNHV6ciTZ+6Z2NTLURcFsu5EZwftMKuprOTrd19UZY
5ZkG+JBJJ9YgcEDcfTwVIprZjJJXbvC+011LqTpi1SC5r2VZruU99h+n0JJ8/obEwenFiBIp/Rxo
lK7CQePH1Pa0FlXV+5khhj246eljQsASiyVBnCsQTuH3eP169PyzJnTmu9BXwhwv/XnH05yIFCF2
D2BNrtzHL2LMG7V/ie0X1EbGvKEiMt7FOqjI9R+GtLWAMYmo3krYyH+VrIMQzLrYJEa1sUpvqCPL
M2mk0vfy2B9ZDRAEhUnkR2zEWX/syCKtRthczqb80A6QHn7HxzUl01AQJne6yRh/Qr+hIQEkythQ
Go83EKRiQvtKwoxo0Lge62iLGS6g/g9dpPrNiBiAQRBwBwd1/X1R0JvuCY//l5FAHoDtAqn/ura/
p4qz2tJD/DWGHfdY9WA2ZMCDssRXiydDJASZF+pNrQWbKhSoNDefYHWlAet9Kmy2Yo3prYlT/Rxe
NJHTTudUAzgBTEIHTkDS9vyte6Ecuuxi32KikLKQcHJ10nEYlfI4o/0cXwYaoVkVK6/6fu58QIoA
wXstjfzu+n52Vuw1Guv4Yfu1IAnUQl1+mLPEB+dQr69JlcC7Yd/oAMKG2uByt8pC66iUhAdzvf28
5UMQrjNbJJh7slr/YhVpxLprBwoae/A+2xGhBdVElaxLZVnxN+vyRQv8E/Md2L+UCsr6qrOqQlBA
L21f7jVuCfsnOw3hzF9dX4PYt5OnfF3ZethDAqjDIeglhBdWYVcRzoqvpJcOCFcUxw46do4GM2Z0
CZ7slj5o60/5h/AmE+Gsv1450LHQAMG2u6b+bsyWOcCZrJEiMQ5pcP+oKisVA9Fqg+q/IGISIWb4
GSgGeaBL/rTs/RqQnbejdlLstI+JdBFRXaQBkaSwUHHa838lB1rFZ795e8DivbCpnuUjMtD2iRiI
NaplX+w6F5XBfzJSUAP06DPBvqml1wq7/4C8ujv3l2ntrQIfBloqDbN2cMlaT8OM67MR0MmgvG+H
k1JX4pfWlTzl7ROS6B83R4j3UqDAxec3bSZvlnSso0PWd4+OtVk/nxVaNEM5SwCPD2RYjCJRsH9s
aCYn11kYORUAYCybTqSDtRcQZWkcJABWFHubBsXGEVioedfFMSt3+OfgB2bH8W6jYDZ972TrhxJD
4W23/WIKgrN08+yYV2qq52TMKR5NkI0a8mu6f8edyXroyShJwgbzmV4USOF9QaLkYizkWQSWDvLX
vAyK+o0lOufKElf8jcY44nucv/peTzePYpP41wZZ8joW7fW5YIqy5+APzAEuoptl7Yt0MxplYOXu
zUV4cncHZH2FiHpAgdKuKcTCnw8RJx/HNsEsEaLDWlf4EQMbIohVnkbdjgDaBZxzxM5CmW4VOFlU
nyzdGfjdfPrifjNvmN60NqAmYYlQ8SiCtoaBUixvC+Bt/NOW1Oo99YdzEiiREWuQFLojGVyeZg+z
4qzrcWN6P8Cx6Kpk+q9aUOrEn1GGycdno+/qsqPBrbmEuUDmXb+TyRI9xAxrj1hyTqvNHxaLvLuc
ulBFPhqHexzACiOXq3qrat7zFob3MhXoIAY7wlpGKjcpHlx0EsvYWNffy4jGw0ZnOoU834vVzdri
XcBDEPZiKXB4MH5k4OySjjPjeam7KhhAhSGIof/JmNkgvTOu2uYos6+q33a2LljIsm2S+lc9xmNz
HFxqD2+UIOw98H7lPwrU3JDTPDMjPu/a0knKJ+0ryJM5K1wm/6RYGN4veCyGDLUTlDuBO9WXTn19
ZSmlbtwwoGLZgPAi+Wr681KKZnRdx8CMsBBhGAd82jo6B68MJxb2AfjVi1prWLUvlP6/LqiFw4pe
Rf1Zez8yyi1lkKi5w2fo3PbFfx7TSRTI41qDpBOL6KO/ENLYsX3ehs6MRF2K7arIkXYDnu2ed5pX
QHioYGzyDGgCaM3BT6LvGf3Cdau6z37BZeK3Sj1FMyJ7F8H038NDaIdEUPZHQaaQR2EoUdIUyV60
v5L/278WplqYiZjhcSqFUKe2mG1YOA0+UrJn62fgIyvnl0nyIXwuyLc+YSXOCKTxBnLUUUJNnw58
zr3mladn0nZHp84bvveyoYNjOPAZ9lsPLh7P9aj0COd4WmMq6npKVpP3okaGbybpMLeTE1s/uux6
J3UvRaysAZ8N6kkoaHoWcLFsP8AaXWA4Y6D0B3RQMULlBi4jveH6DmRj3m4/5N1RDSwjSmDbo8hE
rdpC4DxuT6foQvv1tSeWaYlPM2PN333MLEBA1C4xtb0k/kH9NXlSO0iu4sOwkWJFyz7cspcFrOWr
UDP/1r9C9TGVRZA3S6UNkRxdZ4rWYiSJsCLvzW4N5R1+41rpKPVYiv7tAxGoG6P7ExwXkz5ZA1xh
f2cV1uapiM3g17PQni+gq9fWfXp0maVxj6lZy2tfCC58GhzCvVItI2yU03c8AfUHuhMyn5gu20uo
q03deiEcUvZI1kgOdpH3AIwa7tw5wvTDxQz8mQb5dwj2opRWGsWa4U0Iu4kAn7RTqmIKIgT53fMS
y/F78vmvaQMt24yTWndOvWyclYIQ3ufj6q1MwjqMqRxoVm+eLcZzjtSGl0qxJqgG7J7qju24rZPi
Zf+JAbrWYNRjCnRT0WbYVsByVZ0qxcfQf7fv7ChB5gQLigU7gjStmPrSVXx9pjhdN1cZ3l2mj0BP
4DNNrY0gBFog4eZOsQAXqVyYoJUw5bxXyFiiuXk4iEiGQwyfvr1Y+9dMZ9g93R6IM63sBARoCpg2
gbJte/34W8I+COZh2wW59LFe6b6zcq664HbHfweOruzFFHL0OILpgHlUJn7h7x71YiiA3tcQbMHI
h2e2pkyVmGlzMLqxLzYEgiw2Rw3blU9j5Emvy8PHCbXJet9+kqB/mH3iFHeEUP5iCioud3hKIjKE
iu5eFgmhSL3mcHlKmilsBRjso8MmSNv0hCd30BwTlSqqRLi7cIjeFO8u6aLSsa3IHI9NlXd/F9z6
qCV9Dcqah9W54DyOABLrG2GBVJhRx4CL/14teDgxz4cEWowtFqcjbqV4NIPZatqabHNw45hmSaLy
zEjiUoNBp4kHVNYvqi5cYHzON08/jgRZ2k4SdCKNcF30lOHz7M/f2jv3+zOBqnb5TwhLtH78t5Pe
fKj/XgV84T4KTWBUUzw4Xg5QiC9SyA+4R8hgDM+DfLyia1kNk+BofLg+yt5zTzp2EXCtqlH1eo8l
He6tXYEbU8xKdTwLCJQJz8ns4rDrbz4hCF2LBv/hHFKQsDHuy00eUd8LOhmVzyWobr8pBXp1qtlk
j+ePy2OkrD/kg7r5cA2Bz+smMmoEEREz3GvegL0iY5HuG0knhKSjSy1yv4FYLkGOUXnDpdMrwpLD
p1bKbXrEocEOra0QTzXXXDzIxImZLUUgOLqVJtkxcfmHQONmfHBjkWK+jral37WBb/6KmWPgdgpc
2bmJWSEPn0owqcT3Y7T4xkf/bHBzXcSXhyErfDGPr8VE/FbBOxo+0oC4kmDnHHeOwW668d0kgWrr
NaiwvfrdfGfGmPIBPRKbGn069sy+jzB9mM6iDWUKOu2wcnuPdUFV1ber0UveHGB9yJIMTS8zfe3y
bV6uy6JB7VGIURaCCZoYTR4hukTLwuLTc/kv+vUaisTzP7Hj8ncrIy8G0eew51uWRBsoM/dbuF64
B250KfTRSUSRy70iKrF0N/24AGYsC26jhEya+OZfMHfSiAh5nWHym4g3+iT6jcZ6JfvkU3oovFXg
KIXFStReXJqiYr6+bv5rhj6mXhzbbsXNpILZDMrE/+Hs9/qlnA+mcrXDF82QIHbTHH/4E0PjAWGi
9AUwDuNWN5TzxlMfz//RQrgVVC935gfz9bPa9tSb7aXmmc+Vdi4UBt5v4fmZn/kSZLkN+h9L35bz
ProIEkrlsNbohFWUn5j7H1g1i7cWgoL+xABn7sv8ckmkcJvf/zKKtlhhZuYf9kRIXCBEQCOD+okX
9W/BXb4lnFiWdTbA+2PaAcvM6/XJZl2KgJzlKwydaFxs739ci6yPWDYF6b8PPKHAuPLyJBp+iCz0
J22i6PzuwoLc6G11jzRlSp88HymhMwydOAxIMyiqIAq8sr+I8Zmpy9u4s/mm5smcYqAPmRCw81TI
kNpLva8Jh1aS1DctYGQ6F9nIOvLP1PcstKZsJJOQsr30k0RkVLlC6R2AI056NF3COEBIjiDAtKEy
eGC5oL8YFo9JLjjwNdX1TB/6UJ/a2Pf4rKFcXKe95EP6ntU/pqZAh5MQmyFrDg/gSOGwAoV68PXG
ozvSr6Cpy+HhVTeJeeyzrxNu/ErWsjI6tdtG5b+e95c2LPWPbKmvdBFApfbg91HJujHkST8Y1OyL
ORNtDeexNrKyYSWSbtN3lfZJ1ym5/qp8qpzCVrilIUKg2LvaekkRd1kjm/4bYXpqnfU9yYj6AeYY
NnxDBEj6IS+ujoj70O0N1Sg4rOzPwJJQ5z240IVI845MLdoBjQUb8owUfwkYwyguN7mjgAljsbl8
lqbnoHqbB0gk4IiVhF72fOeHCjvkaJ9AM27Nl7qzkOY5QLhVyl/bSknGhByERapIQTwQv7ecDydd
tmW4r1vHxU4pQI8gqxD2qVVgzR0UiEfulxEnvGXOmhv/HGHunAHgAXIBqGtBFZMNUUAm2ilRP8cx
qSCZJ7EHzA4ljvWGnYzRGkrVueIkkxwGbz7jwVxf2g4PiwkQaGrUruCvrLyvbXd5vrmHxTrIIACa
q+3xmMQjeZ7AlFkd7ZtnQTMcPwBCcaya33dAmwDU88KqRA+Y+ndtKGrsmjfy8+/UKP3iMh65jlv/
HflxTR7AqvR43nxZyg2ju0YpQXmE1HBxe2cpHKgKGdtIGeYLqJJXPN9IxNI+Rm+eHB/gjJrGsJAV
7x7doU611g84n/5kriGk0mbdC6Fjw5l7sMcp8I931ZkeC0Ml6AnoO1/v0Lv0N5CcrWQcFijgREgX
P3c+VEA/8JGfK5ix1YndfuL9uxxR0yQ7e/s9m3kpIVaRVpgkE7D14gcpV5jqG/bDPv9ihQaA8bjw
R6x8KPNW/302bgDGsMIdCjicMnAFQAZSuoB3ysaFfe6bStqB0YvUyWXgjke4vpnbTJLMViH4y/wu
Mu9f4t4iGfBN+ddj3qG0hGd/EgwACxhlWS37bcwcptMQeHVDWerFN73Nd4PBHvdS6t1A3VRhF2V7
9EHTwmR38MlWtlxlE7y39VWORVgY184t5e3om66mUXDJ/Ev9zXXQ4BcmYKOSSri6F8MrDQXDAwgZ
DjkoxgZcBEEuRaeMaFuC3EndMYrQu6UUQCE+dNFT35EEeWF1MMDNce9hot5Mj93f/zj04K4ukiRC
I5LeYEEc2dmioaMGaNZxAT9xb348/wTb+8GpS7aCKGzdxloGZLjxanH+DH3ORNZDaIvS001Kf5RP
GUgmvHYfn9ygEXDVYef4BafheKMq/FfIU/33KzDunKA9WZYYHZOk6c6Z7liu3giXN/mqUD6KfSPu
0oAV7ceVPXhDryCKC3P94kR3t4DiLL76wJPyVwqHmyQHfbp+fDfaxBo/3DFqjkmz2FPbMGHlAwZD
xqB7V+PJdeeUsNPRVdQgNgYfGHZlPSDcp67hDSYDSX8niKjg5TfD0pCd2QgnzY+CjWT7yG3Fe8i7
oAXeEGeZhg8Wp1DmM6jR3BIHo4ogQWXN7sXxUTBRKvqgpETjqfXRSCiQXYjr7oPBC/Ev2A0N1oDz
csTx45m42D7iqIN4o9j95M1hfb42ro6Eb2vOsglOFS/NmmmVB2CElOfmfRxClQTT1PyX1qTvyDEO
M1SYRb9VfVa2UcsObrarUop3kLvPhOwl+4g0hi2JGISnUpgg+rtIQry9yHjBLftYpH2HbRk0X2N6
flpZHW4J6HSryMjAoBJAyesH3nr8TWdaDj41NO2JZEE3+rklnGgWncHwAPvLaG1F+bWd9V8Ui0g/
v3pJIvWeFENOe/OogbqE0im3i9zuB7yfMfa+fuBl+pB7vBNhYxfpQ6iUqG3AjiqE57b2UzyPi7mG
DxGP9cd0Mw5NPAJXZoWBiW12ulUTweW2KDRRKbRGd8xaO1jVyL3ofQJTU9A7EENgbwRN6nfIeljP
LmL7GEcu82OcKVOmD5EXr//hUHtB2QrmlKDc37fabgHRXN1zF3cSe7byFgwVKEWOhpfCe0aEdKDj
rXGSp77Zw5QmfZ4Tq6I8ItuqVL93opISgQLKRhOKX/MhA1QVFggj9aF9gtnr1PW9M5zIAlVpGiEN
UJR1ygc6A+yDhkfjZIw8QReSX58E3AwGiO2O68tx2Hn6aUm9znSpCWi2Ywza1pwAPUuwTZMsBx3B
d1pTvxRJsrVLfugGtmoxVs0Q9wOMnArKzyxl6v6lrPoVsVcxJK9Qrxb+Vn7J3URczT4g0mjIMTqN
6VK9nVlC0fbwsMt51/giRD9k2a99HMSKnUZd4o4nWLkwpMofb8qoKgzj6nsK9wCxN2m9kXmOstHb
L71jUFHJsibS71Cjh9pbTJLQRj5Cyw8HJvMmi6K98akipUmZn6ys2w6FL7fW50OUagLojB2Udzih
YrwC5YPVQJwAdlntaH8Is5beEAbjMUrkeCXcnqs4bQXxNQm3pJ0TYuETOFGA9OquiOLZ4Hv044uD
SkRWZ/IG3OmFqKCyK265K6nf1pxyWnccquuc9GGUtaFj1B5X7fcQehpvZ5l5gPE+aiMEXe0LkoLs
Smm16x7rBRz3B/CyOkrLGz8ByjrWUJuxcB9N+GFRUtGeo6idNWMz3VvQxTYfF3nQsG4HHjSoKUq/
8NwZ3gGgxMKMNPe272/1S3oncQuOJ0G4jI17wXXdsCNtx6FoKWrrzMAOeKMHEFUKcFOzh5Ikzq9M
gYxmZedHUZkihHNXhEKdc8PVSs+c6okjLEZgKjUs+1Q3Jg33Sgek0lqSo56GbItH2nbsIk0O8/s4
DzlXVR+wG+lDPmUQkEgTdN0/Had35DtpEglE2zMj5tamWyTXB8hYdKiN/e/I4jbYH49qKv8k59CJ
OhcJ3Z2bK1YmMRYi57GqmQJj5n1+0WUEsyyOJPDckeEPU9/HsU88k7/xglyMSwyJs4q4IujLrd6q
tTwhWZm7HVjlSEaYzHF1A5I9YQzMKD2r7GODyHQrb+EM9AnaW9sMx4XrYy7JO0+3EYFGe7HaCvNF
NVjcpKdxTd3ZlCGFdYP4kAnjsbythO0aCuP+49fazN/Wt5L6LpTxfq8E+ixN5ByUQCp1MfGQiPtS
sge3VFx5cUaqEFKTAHOKCKCCm/+H7IL5CRGaVFkc0CjlcnnEQvdhNuQVByI/45MVZ1CsiKeFQXJt
eJXmLvTUJ02kzEDg7cVfdDQ+PN9ookhs/xcgQkpPjyG2U+/XQluobxBAokXxkI++wj+QG3BxX85z
5IARaWFD9I0N+/T68GuWIfr0coNHh9h5PNW54h6P94M27fxiEhCTFbppN1eEK4SMjlgYGQ4ZVeGI
hqAsynf1Syctrdk5hJOuNo6fWtuKh56ZoJucsE3w7mNop/pR+aC3mUcIMHn6aROykRZ5JXyFhd3W
mrCFuOuNSGEUUSrExytUCs5xs+6p5GigqU7p8Qg7JvOQEHBOVKkbSiI5BrNODp0VPOdj4aZOuuLk
YQsvsNCsavNIbYozPEbibmKcCn/I6rWUA6sNWnK51h20JSdyrd0eE2jm1Mf/TWBiojD4ux/i5BU3
ijWRzIVQnnazO7s8MIGUAiz54iFVr+CsV3G5cSE/ahblLPVak1ueSX0NMWzqI4Egjlf6/b9aG9Xz
3t9kL/HoR9Wdeet5GwySR0QURzSX4ubMQ112OHv1DCB7x3+XFbmiXLLRl1VNk3WFo3pyeQ9xwKDy
ALT+kEcPapGFz3YfJ8dgS/fOzuHSMnbwpvwo/UCenJETiqctrX0FnxTFv2LhG0NHyYiNkQdEuNor
sJuPI6XhNRAXSniT39uf2pUIqdMHM+K1LFenDYMma10GXJeokFj0vm3ZHfMD8R40lk34Rcj375Ni
zSiaTl6a0w7mlVb4IAMCP+suoShX67HPyegck0dWY7/CHodyje20CvFnyErHM6p92es+aSj0Vztl
WtxEsHdEhUphRIofsXgC93QAVXD21u3YCJXQnnx7O7hcGSn2s9fEuAOmnbLxdEiIF7mIRlskKnHH
b1jam91o/qSmJ/BFgbKEQiEj+i6vkzdovrcXHgRCJzSPapghgWpTV76UY2Uy0OtAtcqWPwU5jner
77k4vgsQcADGL30ucT5nfWqAseaKoR8h7x3TzHd57mg+neaY9PsdCIQLzu1+322BmIHgSEB/QUBE
+Em1onlN2fcXiEqgrpJ1x2Cpsf4KeO2u49iKG+vhvRpjuX4bUUTkz4vqLirnRHONl9jVIR2twZK/
BQoPAQdO5YavYhu+UNKKMGIosw5nqNAeLjDYyWmxgnp1GRGEV2frHaIMzXiQa02Jym0nU4LPwT9O
n/J5JHqVI3I5yPNnZ5WrcCWAzsTw5XtPVwsz5gaGyuhlEyyKm3CsDlB2y71c2OEDSYIoXYcTrb9V
FqvGNl/iKXVVniH85agEQt1GkHrltNBwwcdiizrr+sd0MXoXNyrLxw8/vewkjzUxzwd9RmHEalBl
LLdGgCEZaAgml9AEt8dSbcly6imPb3STbmGQLtk6U9AJFwjbdehalHCvvr/MPtDVZpDD0Bo11/27
WDcziWoL4ltxNWnRIgaQwHZBAgfwja78bqL+Lz4011mauowjZy21NRJCH+J3m8AV3ziyCpwS2FiI
V7PdiHErhV8GnF+wNdgwnG9mQaxJj22gED21aB4Iq182krHr5jJIHHZAiM9jDxcRv5fTP/gjujBf
UD94XONYLc3GDj1d0CrmmJUd/dgaCgeNTO15n+Ef1egaNYlSlGvNsv1TuLCj2CfFN96xn7A2g4Yy
yFlYbQ0nkoP8qf2OIxruUm78eN03mB/gx4TTUduvlAqwjDydjRgO44zK0X/sBvUU0Kxij4DBZDe9
1AREbsUNjnVopOKXG9GjYt0MkDJ8lvH7N3PDSqZjjmyy6Ah5IRMDCOFS34cflpwCWxP1YiZVEWFN
w+8ElgrKDetr3oKSqu1t6Sh7va0L7uCfqd4oi2lw3Iu0SVrfnOAwqTt1JmjrHCayFX6+5Mvb601a
e9Rv0hVsP1FqlvJvNe6DvQ81snZAqA6j1Q3TcA5M1B5JUS46SS3jCw5WtgodFX7/QqHHilBadu6l
iQRBkr3VTYlxdGgKnUrHuLdxTmo62orKicFXZXIHQnXvDlF/Ij4X/qVdIHJC+QwT7xl0jPdsq0qh
X9+AGWWE/3eGcu7RzAolfHXLRtm7V8ziOwFBUtFj9Lh89u/9SchzH+fuhbAKdNFVkvxnhvkNkYy4
b8B4knAAQ+H3C9W6gHANYAGdRPGgJh+BgWE8qphbMZ/niBq9ulEW4dBw+f0UVE9nMJDvs6pvtRsQ
ZDpLVXjnxvVYHf7Fqzewo2b5dLfCjXPkEQdk86t5BQBv3SLbt8us4BRyqJTW1PGPK3LwTNXCB0MN
KucY6jLRVPg4q9VeqpURi09Fx1QMhKwOPOJR5cqP9RWhURf7zDyVLweFmIm86R6lwR73y4BgnBXD
xpygLaDskZqUDEV2jgMZd2QhoS9Ze7U/ALdZu0ftMSOrX4fK5LVD1eg9hNcCVdEGyaRAXFAOwOWg
cST1djSPwGSIJj90AvuyNBRLeWWnJsUT5ymq1nuzDtUL7jtAdb1yNUSTUaVCIsSRoQ9tHdWTRrEE
beiBcDdcYybjHpVBa3aPWUTRh6xI8DQfFkt0iuOkUVXc6IzSKR9OFTTsxWqdmtJ94XnHVbeGx4M2
vrOnoyTgOra8Bv6OKDe2L31n/QPy454Po9el+fNyp4Pr5ycckjKZP6lTgH+eDPKg+AnL/dJwPIzR
K5l0g+RZDWa3nD1C0HSTXTiEgL7Pr3C90eVdTkCE7XiOo3NGQYPuZN1zzNRwBOUDWch5WAzFCzcp
RulBCnJcoYazKkHzfUEnzVzIzcTkhCL2POTWvMyHlmxX7dr/BIOfBvN04tIkz0MiNDr9nKioUTwE
js5ZUKeelEaFaU+xIZ/dkMrSk1HNS2AzScITm89CiplsycxSciOr5B8OAM6C1uuK+nuLMfOtSPPN
K1WYnRqLSz204JuQCjp3xZQN/K6sPCRjv38ChHHkB9irK1FxkGWBme1YVa3c1MlYMSAiksx2Ruln
xRhfvk/sxpvFNepD7CyKoc+g7h9sPIzuDLuKeHb4fvt7tqJZubJGSw9VKxGvvimn7awsE8YgiO3Y
47ECbDsax3j4iOlkBZlpc6QoUauRMQ5JMqMn0q4lH5KmNpDItNckcpcRrZPIHc6/yN/7Fj3VzuqJ
doM2VRdbJfeNmefKpwApUAZ7OvXPvs5f5stQJkKQHhovLXgvn7e1+1nDapAk6r95ThQU+j69qrKJ
x1SdMEMp4m4BpmYkXxuABZY095L76sD0jj/R+pWrVustf+numNjCZz5Ua5o/cOAxYnC3QDXcDfwd
NbXsb6fBRPx/8qwyBTscLwSsueZmAN92ty2HO+AMD87FprhG4DgI1HbKqAl4XrqRLwvceHm/bI98
XNYBx+hvTp71px1H3gRfHc33lbcFnj+Ze5x/Z0IPsc5M9StZkL/NeCurqvWoIo/zY3nnhVbDbpjt
5gyjuXX3cczo+iQml254inNd+Rt+xetr0qNRjFrfIuWo9YAob3AUpbub8eKLhYi00Jkuzg1PlqEN
1HPQVPOWSLA3oq6jrEZ2O1aH7kJ4uzKDnWRGyRbPgOrYbR6vtI1SKTvPnpKk31nw/GOMXIILq9ED
OACWOGK4XSXuyhgKjzG+pThgECJxcL/bVxqF9NK0qOF0/717a3zfc4tMlMp1qrmNTzVysHg3xP5H
ko+tJAX68AGh8z97YaU19TmbVHFN8yuEM1HxpyNvl1LKlV6SD1use+ilCIXV8q8/71+9wH0Hw6bJ
Yv9skxluhs52+oNBdWjuHWZcF8yLIfj5QL4gcaF+AqjS6h65/OskBKlyACTR21ZhTclOwCsWN2yf
rXpx4WZuCg2D2Kl7HNGuGEUGlDUUwbQbrwPKdPHSlLpLUyZh9wEtIKJVb918FIVL65Lb/L+wyOVd
IhlZICWq/trFkB47GAuVTl8xNzxSiOVdKVN9/Pidu4qdjKq1CWERRQJ65fg5ssx2TuycgO8nAMb/
6zl1KeXENxAEo1EEkIt8qUKjiZuP9A+hF1ylyD4VAEIxrE35XwFxbS6VlHnOulT0Lhxyzq/n8Hq8
fLWiZVgP1c7P42q1B3v2aJbKdmE6MXVpfz4XaHLB+l9xd7N/IrVFd5/GG5lPbP0/R3FYJGBesp/a
vC5QBzdszxVBo5ma8StXcky5H1I1x9YI/nmPuDXx67nuHvWwg3JzZ+uF9zFLddgUr6/dkn0GP9B0
g1/I3qlweYerekEYp4TXGRODACznpp7BiGx9wqb5mKFP09xCKlmdF6p5JtGkfRZbV2LBik2k30mi
Tk6LUFXwxNnyaIFN+hPYgXHQX4lhGuaIKodC12kT4FgRJvKLjBs887aHywUfoJ8VVitS9gwVRxg7
HugEwSHnHY6wADiRxWjr/2mErD4Uw4EpmnXbFzhFl7XLKhCSPiESQZCBcLX7L90v7YavFOk9KqOQ
5R17TDIRJ0/5woFiMYXM67aM4KWoDz7ZWj66IJ6fUma/c9n2X5hVJnShGxVSiaVaLyCsrQPVKzW8
UKfTH1mil1tale7tWb/3T9Z6Z0iNdPSLubqshySxpTdTetx3A0FTOPwk/o16ulG85oeGKMiOFajs
lD0gUB0w57AI979lKn+ntqe4WvfdnbZcco4yzGzythQpTM7WtZSU5P0Q1cW7nCAqWnyYFMa7VumK
dcGC/szr9faBJjgA/j9379wn3ZZ2MLWRKJJW6yVk5wt7wzgyoXh941k2+2ajOrN1eqZ8xP+KZyxE
H4DYgw7xByPwH61j4NtxvJbtFkB8A/XVO5LHpfHLqZ1UyaKNVuH/AKoFkUhse5yaPBRvv8v2PrLb
r2F+BH5b9Z5sIw5iQd4CaMkTgXO1iH2+B5G34RqdDkoj58s5j8TFCAomuzKTKMJ3qB1inJ+lgkbg
mSYRoGWWC69RhnPM2AhIeMIz9oMMAR9I896uDq3a2i6cRtA+yweWDfLsSFUgxqD/6/wJ43ke/tOm
oQHVT4gbLvv5oXf8vJJOV9j94vEQhLlSappTMIiisMCINBx5Vl/6j6T6QkbnME0RD+9W2Gl9jquA
6ldv4HyfvsgJ3FiEadIdDuIKaOij+/tG0imO5iIVWzAH7mDY+34PD28COqNYtpqr1Gt8HaStMzJD
UYW0D9a6aHMwgG0veP38HXSv+Dau4GBBpPC3sGesi90n8o/c+gKcgHFpbxO0l7AqclKCjJSLiRWN
UKGQyiodZi4nGLtViyRy3CZc62zGcK4RlLv45GIpuOHTxS+JcnztRDfVD27yGdazkMOfvIoJJXL5
R7VWsK5cwZtYxanBoT7ftCyXZq6H6Q0limcxOKC/e8Q5EUz/7HMlDlMJleT23vo6caQij+dRL/vS
QlgLoIisdNo4lo+Nsl2bHQzW8OqbYr4dqFJjDaHKwFubmI/pWn5Rh7UlCOug3K7HQ4cuInwzN2zc
IPzcacKtaruCGOxcZIOMtXIWoS0oGm1iYkMVpAWGeFBIBqTuoVwy1+cpP/Jax2mzwaMp8nZbrXw9
ECHmI3+fHBn0Noa/OWM4jHvin0On0fPdxi7c+WC9LJAGumPbY4+0i9brOI3ZnLbRHdtel4XUjasx
oCUr1ZzJqltIdIWMrqHU5pZwTIqDc3inOpHw1b6otE7xv1wxEnlxqs8pJUsp3JzXbwibYkoux1Qn
AJcHVOkTAlhJ6c61/lVE/LxEa0lxMdL7aSPuPYnEDs0yYQh6O+ejjwl5zLUIl9c3oLWe+CJnXWIQ
UR3F3Dyi0S6//0USA/tuDZrlKOSOIK6dg7tAlDOYtKyt8DVBO5zjMswmL4qetxcW6eytsJZ+8oaE
uqFCtrsfEC/3BjIbhZzFsbGbNLqzP8jvc1Wb3jXp8+QBbb4hb2IvuDAlsVJN/pX/FHR+8HXZYWNQ
bLn//ktLl8kaIJpa+C4Z+NOMpmxFq9+F8pWI+vqQGAmRY3JA+Ttj2Oo22BmLUcRpslNN5sh5xAWr
DXFGEEJqNf+Q8aWrFO30j4+LpvNRtJUnWkVSEhMWPTTrJq48b5ML4tpDuaqzLqqhYzELgPbKKjkR
hnkguLKqUchLOyHdJAFekjFFu8+gxg5fLHXSlhPDVyg+SxvNHhZ8NKqmMFZxDTAzwoetIFAmEATJ
AhTuUhsz0NM12kvQ8SsyoxI2OcTQT76kGI73m1xq0iLqFMIPWo9XFWCe7R2OhKp7y/36SM21lrF9
5ZmKkHiiFNlFlA94INwbXIixstov3nzkM8Q9LtbdSnpyIX2aa7nnjWNbd+OaFoggjq+x07qrMYei
nR57rW+ULkXnoS8pxm+QzSGIQi3AAFq5oybQvQboQayMxzQIyp2gYX1ASh8i1NS+o8fKYFHFiCUB
rdoGLD0gaqxf5N6omlLgsPguE9BoHitRpuJgaeZXNVux5rTmp0OZ4m7YSApcmDqpWIe5P6PqisN3
ndY2ETOMlWybpi4H4tHnLUK4KgS+plJIEySlyTRpfdITWZizurpJa8eGJe+HvIkCKjppzrr4KgZM
9v2qkU8EuGee5Fp0YgibNuXJz6CZJ5uvWKzMiZBNJrDEN+KFFzFf1ouDBxDaamGXgonacHGL3rwF
qMrbildpvNYFnLM0gQqC39ASM1sDGU7CBnGOfmyAFS0KwdxsTtkbllAfBNysGMq9Q5lKi57VL9ud
YC+7lW+out/7PfV6w/eObiWeTS6cyrCPJHFJNSYZYmT9jF9OxXFkzNuTa+QzxZ+Gu8ECIuWGb9DU
gXxsTSP+ehKUxSkVakPXSAgGvpb6dbGi8TmwvFgRjsMI/btB97lxcLKxzAPFG5H0dAafVJpN7HYY
rISWQe1cXVw6ABAANu/TQNczQuwUrK99W15IWMPi/dXmqb3wjqwsVKGmuj/UFy+6NIAwlR76q/OR
1KsKTmsQ1mMms5IhFTPX5TtwSZgVGXCk8M4XdtmdUdXWFkjDPlPwrJNY9AypcEWBfeDKbrVEiE9A
+S+AmRByCGd9jKqNI4kGD96Yd6iBrDTMimJTG1gI+SAi8VVOTRMoBI3JQLjzXt98FUMYaCoRHP1/
iUB1CltKGD/sJwylKtnOGoxYxsV7mPD7/saxvBK/NJB/ugRBZZqz14AkmyOPvqshbaR0UvR6XKzP
UZKKa+Z3SfOFCcWiSsAQ8U7O2DuGjcGJu6cpKComVqRaOmOgHfHRBTbhrS8iWbFbr8Tnx57MVvh9
yHKL2BvDjc3C5OSm2K/m/9WHj/s5DQWn19t29gIQ0lpPfaHkO5uhqWI1y6SsBGtx/yD/GHaFKzHF
JLT3K2wUQ7Ba1Uny/WFRwbhskVCtMNv3j7dwIQPwZ7ky8eLw99Vc7h6FiZY1jGMhu6rVt5ZJ7She
HEGoE6Vl0upiHtbZ4NKiGsdQhxemwQvq5TmOcA70pv8Usp1gJsCB8uVKOLhTIYi6A7afNuqbn1oH
xoQz6vTaM5wvzAFpHwut3HaX98rfNt3adlhIXA+HDCorGypN92K0PJuXEIn0Tf6+frT9ah0uotbn
zB7T6XvD7crXtLRkiCo1s0eFI9gWXI6Q4mXbP+ja6lKdoAd9bgIBfBlrCXVa3XTIWZHvFAIPLfeg
N2ykNcCv4lmXupCjNVYyj8huXH7eE8o3o5PQpx4erWRj5mbdVHcyYgT9Tc46XHr793BPoOTOST2I
7NtbP6zTurJcst8b3Ug7R2pUaox9vIzRQQFvs5WN/B+o55Z7me4Nh4iN3eyhNye9DWHn/9F99ovQ
68bgtLkpehTathBqI5RPuiAKUnA1gDqB2eKizXd6IGo2QrBNKhIrvRXHP+T0a58rSo+qjZwlHNQF
7VcUIV/krvC7seyGY7PjsFsW0id3iup7aAZPkqx2Bhuiz9AumvsEFxJyix9QyflVRi6nDWhC1Bhi
g1frgM8vR/H1Gm4wO4e/HyUDClhUI2fLpdKBrSKx7w1BPSTetiMI+RF8+4R/RquK4DX5NF8gYtxs
RlPO4pEbq4cFRVKcve3jmz9UOfkZebYQ2TzOUiW3lOoIEnTBJq1dpUjGjHFtb1I7PrVH82MkiHW3
AfW6J+9e6fU9TAmCpqFI2wF7Bdw2ezji9eYHsZvm49KrMs9R8Ppwdp9k174EbBtAs0FYS+6jDZha
++/x1EkNe1A88f9jMXpxca6k07pbU7FWlMm0yF3XdhTtoo47JMwx1kQBW1eS/Kxhl/6I/1URQVmJ
IwCNR6ESbUzZ0RWAJlitmXgzLSLfNtZ5mN/6qwH4eU1c+irg8xAHfF/gQ/6ca4GKt1OfNlJsDzhu
Y2DMYL7a512qZ3nQmKb+RpZK/Gf2nHUf5bSM4xeziYrPq/axtwjm/b1lt954NIHavYlkjKSZswCh
YynI7MUNpRZn064XVjCw/3IUz97gb3/z04i9VPGxWeTtCMpNlAPBVh3gTl6KzJyRZmTBzB4fv/qv
hEOLGgiwDP0mEf/hEH54tBEGUU6SfCmuf2Njs0rgzoc7rKpb9EVw5ExybEevnHc8mxHIEo8b2aXR
FdhUcicfM4sCxSjOWJmBRVu/NhLWqsXB1Gj9VaLvrpXBjdH0+AmJt92vQp6yl9PTQ8VJ2Mna7sXR
F6oOLWTy1yrZ/WdzGwS2NQ/M+OJ5fS6Q3BRgj7hw7qVeQeHZnjrfO+THYxol5wIau0Yy9595MlqV
08FLZIybmFx6RdnW5KOkiHiQK4e7WCwvEaebE5ks6kjHG6Vr6QfnaL6q96+wWKHUVXr6pgrzHswS
JyJ31EdvzkN2Qj2tZb4YHFYVk4In5wq5eWYFWtJZ8DxDAcQ6727DZisI1+WzkcUNmEmBXd+GwJlS
I5qtyiHLmaZNegSnoVwmJkTcHGVOqmcca/LA2ziHorEuyx6fI8P+Dv5F7saiYPyodFlwB7Anpx3g
zI986ynOJllf+qhkSE3hs37RpI4DBCDxikPJgAcJXtHL5tPf+l3U7Vditw+gyZ0+CI8tvyrJQFbH
TxrR8rkjj5EKfAgZPE3P3i6h83DQJYy5nhX2JrWeAiEJuMpzrlgcIPM74CRlS17iMfnVzVfo57bB
5Ccj4evuCCviDNEr8UhEheVYK/rLr7E8WajWMrYa4ZRHy19vF9UTUHLI2CFi/ISONtN7sS2GG+BE
iQu45GIkLrS93ILXaPvFNNsIB9Sz/dFar54sWY5d1EnB8wudUOqJkvKS8/9XJ4jXWniUp0Th44x8
Heb3Ns5rBRfcWjyBJeMda6KfGqG0drTR2WFx2kIZuuv7wMHLiCY6zpaCYtQhgdPef5BuhQsrRFo1
UsP3Uj+3pizuVaj2lyAT8PY07an8wn503x2q+AaMKsrLHWL4Ce9YIGiIw94h1pdMxFzi7uTCWenR
EAcz3O+0oZNyCs0V4MvjWdvCHbiy4oEUslx70pl88brkDrvlC2V7UdQmfIDaR7GBn0R88oXrg0qS
mnkR/lXHCIBpAbZhI5qDoTEVyAos11MqNaYjblK33kfWNC5rZFt+LlVKU1AieLP9HvjHdr5JPnQn
J59oHAyNEI4vlKi78wykbNWkLh5FD2JhwuyUVnD/kt/NjsPp7QlIgGClhGMP9ffgjAek0KUMn1u/
8Yef7q8ovqu9MHphAic/J6VkX77Knh0keUZlwOMgFMySUvPELizHdUn1ZyPvFsVCDaxuxlKNzooI
wNcmnMlIVeW77AWeNZetoZFCO5jFzBMazqpVtJB0cBgMLrb4JGJKi2lyqShl4YadbTTm0SuPV6cn
VDUaRrGRwX5w7e33YjbtQkCKt9+IXe0JnkT/AmSIb03FzQlfxTf420o7Bu3YAbl3DP0ge73tmBDF
muFihx2hKGcQdr18kcAqf9ujeLC7+GUiahtfu8DJIHV51TZokC+3q6QVEmQa7O1n+pKoHLsy08mI
0MWXOI4NAy8BkTR+QBWsIAg9eT/xiC0p3l/tMp/mKMyIEniSD5rAaqu+92D97wEvl+2ULkWN/PjS
fyNFh67QLuCug4DR4boNwy5nAA4yEeMH4wPH+xjq0SHU7gWFevphDzdZOPTENBqmSxaI5B+U7Gza
j0Pwlevd7G6eyZjJh9P9iQ4hdlgFHn2STODbyIpz7GiLY9rJl5F/n6pgwSgeLsqmWnlH2x7XCRVS
Qr3vJHjrbYIXCbZzbM4llYBFPlR2JyZMgfFbNejZsus6Y9HaTRGyjNKrYqXAb6rgJdDWxdX7Oy8H
Ou0Oc6Uy87V7LKrK4iMIvdEd439pJaHMkiNSJbxYtI8wvCMHlasz7ANxGCTT3cj+qZBk7M9l5lXp
KAAglTBYBq0TX7X4f1jRWbw6TaMJStEjNbvNG3VYuZ46QCPO0v3GQa8NNxwIGbMtK/RO8D12w1X7
Gx3UDiUr3YcdmanH6mJgc1sYJUgb4DYOGzYvFIaUDqB+GU+r2b6jW/Icy02gtWTTtKLLJvg1IVbv
WrAf6zNblGjAURRygs0Wa6hDijAYh3aJEdUVSjB4HROCeG1Zbl4Cakiy56OjIMB4Au2uGt/s9tA4
Op1YGAjoHZGOpvyA5ztgF3gooJSYoX5m7bZznGxrrg/UIBKAEuJFS7/0PSKgp4mVdVe/igoQcj4i
WkSyxAvgE6WqyEtjEnIDnD0+D3bwVdIg+44A5CVI2B/Qxr6vU+lp+1nbhe+jmZRx45x2pJMrZXZv
BukYYmwlfwdDcf/6OdSLFOTpd9HYSHUFWAIBWaJ2tHR+CsV1d1qJleX5U4/ilzIZHKFRLyeAymv6
LVUX5EpWBEm5effjjMt8wRJqSnjy3IcYeHvYudwu0jfH5JzYQ9gHvwjkMkcATnpoGx+784EZFYz/
oODClqvAvFoXXieLQolMYERwuV/LVGnS5gvToswkABRU+ZkooyLUNWMP5rwM0nY+9RlRHRsYHbUg
VDr1qO6A+SnndaNTdwNVCaCSD2DZHlFeaUHQa31XnMDERNlBE98omsqU5BG4+WuAOXyLSLu414FJ
eeldla4QkkhfY3W6p0yypvqwPteMkOOmHf3gFBexx9eUrU883NHZKX2FLjvCvMaCOTV8lXhY3Njo
W89xcxyCkE80ciwPrKcqJoAxvb4u+7LPdCnsfA0ourglsLz9tPUYo7/MIkTHAKlvmZhCOGzP1Ovf
eYxOsYb+mEBKQJLO2N66Q0mUFTMOVXLia1UKd/VoQbNHayKeAuBS+8Njh884GmgJ96rj5ioWPwhU
Inl/LJNUK+J5EWWtDqZ2UwoLtwbhklbZZ7KJk1xRiHNbINkzPQDbYICrMV+ov9oI0ksB51dfz5ET
dVLugWuJy/BJVsFxhw9wXKlr5BOjGAJ4m5iZTQt6sVVHo/gSQjlb+h4cnu1d6XIFHIcMCKVsE4+K
ZPIzoUYl0hCRCMmE7aQiHDKN8Mcunp7B7h5Ub55L9LGS1/cCSkl1kNoooytOi0hHgAbjt6Xyruvg
/jSvhD/kSfMhadEBuUhlC/DDqahAAumukTQXzZEehAsgwIx2uxFvHuTWsjVnqv3JnAXYTQXXTtJx
tLrVulYHDdk/cqMV3dbWX/w1znH8etD+aplXfnyu0zNC/RezJk3bzNJLPIDT/GWY9DiYjPHhinVs
gUQTLDCcEBwJBk+CwbM/Rv/QZp3yC6C6MOozL8wb9LGILo465nwE0KNJFsGBOSST+sPJZ6rmVEf6
HgSZtnRDUpy7pRGvxkB4st5502tcTrewjWWS8uOZp+HCskax4M5JD5/WAeIbLSX5ml7izDDOPLRN
vFjicC+W3TU9s7YjtKE+vqm2DHY4QJtMp0996JbBETL2gGxbda0rDpqrgUcDDnFJjn/hd53z8866
Ex9CoYJ3Q64uBeE7JdBkzPE3/ZFHl2nlTV4fHzyN8F3KsMuAVaxO2RL8mLn0yxIM6RD4NYd+zOlJ
Ros6DlOde2ifF4wdSMjz8bxJeoKaE4Y3uk3iTAojlDWrE7O6kpLgwSRkIu/8tizMMD7wFAG4XPB2
yTrhAJdnLhggjRQE3vdDf85OOBvrh0Qc1StfrxVJ8NjlDG8gue0JD5y3TcOltiP8JC+Ph7KAVCAb
sPh9tC3Ddn3fC5LpVM3XO36lwMUApwmxxnSywiqDJegHWZen3tqhbJfWZ8mal/AmAo2GbJzZhbLr
GKgOcUmShDRCqSggm6s7i8xzhBSj32ufhUNoi0UrhAeNM89nLdQho5yEQvO0PnrowOU4r/Q2Z0LB
w5lN54ikDmSEv2w8iELjg5n6UlDn0LC9RZ0o8M0kLqDbq9x6Wtm00zPZSQGm+T/F70FzUGHFyeee
+K5dwIZgTjAufF5jLvZeRNnoCJrjUv+AxsjDp9JgOlx4rcofA+pKq0TY3Ne1jCdxC6K9vKfrCrE7
vbTwO87GEYlVZ4CicBnA2meXnEG/fUJutvzCMQiBBFghDt+hLtJ4+hMBykEWRaM6aUL4H+L+D402
xZvQant3MJZvrvZ0yaS5lIkEg4YTstXPHd6hCgQhSnETQ+m/rVBc4Pt5ECA3rS49S1xJOAQ1bEd9
Jn2wPsaHdgdR+F2Z5g3LKJt3EVysEfmTO2Z1pBXSHCFY6dN+l1W0lkT1o/zp093fM6Cd1ypA/c7J
GIVEyAHsmH9K/faHutYxLXzAniwxfZTJ7V90hx9xIZc2EncXH4zcT6yVCxXEqyjW4fah6HeFle6u
2z5cVgp11d6iaCElpHuZw0ZvG691W7VJipLoE+9MPjB/l67VHXqi+WkPR4eNzRhA4IpfmYOK4DmX
G1w3RWRfoZqiAY8LnS1pUpw+Vh8/H1ZB3/ShU/mE60Bp846AgVcCZW2Vh/l79delnacD8NnYAkzU
V7e3bkXmx1/M5O1WNantiekpeRaqcRil1T8lQwgy522rUl0w2awIsWqiGNkala4z8LM9Xzhoq71F
Bv84eYJyC55ABe/DON2ZgymTqaE7NARR5aX204W3RufZm8vJ/WCCZzkueydJYtOWk/D49DY1LXWE
rfNSc0cfpdtNHLUcbVOhHPRoxtqjTnMx4nznerb90Gj10zmUzBbrgcIJF5rya1jOmy45JNynsILF
1wHeXhcRovkmSgPtyN2DVqrX5YkdNZ/SNCRs79028eNxGFueXkpLuIUHzBrGLrhnaPgwnZWYvxYB
RNWXSAN9bfQnQNPYPI7jI7GyQWpldtbpR/watb5hvapbMbMdUpPVfqCBlPeupfIfdpakJQfLAALC
JwyizP+1wsTYOycDLWidw7YKXLI1ay6kMJGXqZKR11h4keDIRSHIpPusAsaiuktV+oPq+pw2aNbi
jbT5Ll0QkP0VDjCpaFAyAsOELcgJb7vn1ZAVRk0cu+U26LNIBkYIHXriHuxiAHNJ32wttCNnhWMv
uIr+x6GMZb6fjovo1S2Mjc1fqK2dYbjay4Co/WqsnpOOKJNgtcpsZlbgHyVT9F6h9cE4vitwecQt
ms/8ESfoC1KVERpm4bdZfi+p7BR8wpRyMEQX5pzm3ODBh+sLRTOi92F2NirNSko2i/xg2fXIErsA
+a4EVe0SNW9hntnq2CrECmSKRnSiEPFanix8sP11hwE0+oymgZOkacu3lYxeQ9u0iUIxgIAwRlmD
UvAMQboRSKCFF+IlTWHjPZCeRcNV5opgyMy5QORXaqpR8GVDF/5xtadQaK9axP1uNSTzi6bBUEmA
AO1pKlvpXO2C/eokbRjswXpLVNPaMq4RKo2lRIF5281NsY759JuKOrGbt0beD9oqzBI6fPa/Mb6W
b7WxWcKIrrLeeTBD3OhpIWYmjbJudCg3MK8Kgimg6ufhdlmh7kq8DMpA9ZjdneZ8N+eh5mLzclt9
Tc0HSHIqt/PSGUQTw/OyyPd3qDTPVdx/FLmzSflt0du3Qn/L9yYBXhOrl66h8f4aWcbEDgepfVD8
oPR96MSoTkpnGdyNgMNEV64nHRMapJfXm6Tac3Nm63pNHvqIKpFL/M+8Lj5TmJMebNRi6FRrwCv3
613FqO/C6MQm9Oa6RPIKnkCRAtD6eBpDNK2T5zPtcutASwq5g/5sCSPZLQnCE6WbLVgCa4mwcgxN
HVcGLAd25e9VkLhHhZPVZpJrakdloS8IVaSNAzj9U4fWeLA7Z5CdllbdeL92EUtSFD5IDwLseRsq
80UaftuK3bGJl9a1FSseoxKmZUxJiKDMKm0trjOC7uOIYAKcxuIxnqw8AgX1Sp32FU2Ne6jcSRdr
DwHKiQCireFreZimQETDwYTy32Ght9oxXsTa6loALPZUIqIC7eeCvvfQNykfy+dW5CJmm2+qK7Rx
PoZjdjYQWeySKdT+pV3su7pHMEIq1n07Hp+4iwvRJ0LffuQdR+v2AVu3Xh9kLqjsf1Ps9iMCwEET
F9Ef+0CGXEn96Jaic20dOdKDXI6Zvwl97rrgyBJ3KnLXs2eQ4GflC9hJuMREag2UeElo5amENBoT
QueP5fyBgOF6eeQCNOUKHzbrE4PLPPU2Ts+fWeud3cEGGfra0G+S7ifq6d2A8CCmlosK0BZ72n3D
ikY4f0xfmULDUZoGSO8ScqlvfRSkzChCCiDjRDiHJNywqaqH1dX5NRvVArCu0kbsGUkvIvwYV/me
6sDFn479WAA+stmsCQhm2MA7LbBRcFyaXy06D2gmowHHGLGYwOF0WRlShrdR7AhWItGZW6gzZKss
uJW9snr52EXLuufK3RHus0tAIt/QyVpon6iP2nK3t37qikx8/Qs5+AIV9BxJ3Toc47XwYjXwQZV6
rLdcrXZIFonOzkmJP1brzXQQmOvx4lDC+pMExWzYFF4xv9dwZglbyC6GOq/dzll/1b6ArUmVY0iQ
VD1lfFl7Ascz2E6ay0zZ4dXjJJlwBOH5nWgMMvTOJiZ2pWZ7WS34ASgMHQ+BuBoQ/5O9D5l13XpC
g/uMW91jaiJ9rFgvbSd7thko4pKa1EW9p2LhmUN1dE2cNjMJR0QT9/OH3lrNOB01NJ8M+gi9NZcP
6UENLIkYqs+GMkHcEfolQEEOgWQYumFpV4RBWlivUQbB0h5K4AL3Bn0gtA/2o2+K+onvelfcIo5k
4UeikjiCxx3Nh0ZqM8FDcKrv4xBNiQcCud6eoMtSuINc+QNyR4CUTRXvWhao5Qx8FXMrJOrXq7J+
IiXu8GxI5pu+IP6s2aOXIlN2LkU5YWxe2OfOrOJcftIMfhsviws4aKHC1fZJh9mIu5QqKtALVeED
lr8YEZq5kaaBkcx7yX8UT1ylNMspLTUwa41RQD79IYQpZ9ia7CZmXnyIi3bLyQqPvKGE+1GlHIEx
oX1MUYG8HoIoDD4juoF87QULi7OIMsHtw7W44ewBbWW9TmqKqyv9xwb4+DEw7TIt/cDcFCzktGyP
K3GF4R64sK75WWxFgkOhFJdcLEB0KHGPAS64M7vsKDO4CLSyMpgC4H1F5wrKFsfScfNHkUkswbrP
nM5jLzM3PsFhUM6SE0TRS9BvFe4J9MLrQsAe1vltxQdu/kwGvo4lnrvDIOCHEmxEWY3aqkhX6fqa
AlBO5ZcffjOV6342cxbUUZHyXHYZuUYpvui/rWjOYFnPacOPW1wP0cIQXcaA/gYkPQbhbI+Fl1zK
7S/wvkFRO6UUy+BrUsFT5iXdOwtuTRgtt7moulltClWi2fSX9exXtZTuFTFAVX7E81fZd5/0CgJa
bYE38Y0I1KRRsI2IRVeakgSbDtZBtsR4UxkUPRBpoQ6QbhskGwStufdLyllr6xqK2QKaOUxQ8rFX
ip9VJYjT0+GDfkX1C2Iu0uxwScGZE4P261mwJqGzudDhyuYKFB0/c0FfsdWeHohgeH+yaU1zVOO4
FJcqH6nDdWOpsFxlkXOycM8tA3BWOFrbFtCGHneZJSBN6RqU/ZVuR503VZzKHdDQRvORLCLg+7EL
FvhoNpAP1LMsqSCGpmxGMELrQSO6oUhcqum9KEu/shDRhA7B5RrPT4s7T9M5fAlOkirp7F0vVPa6
m93CzFSPLuvoOk8wVLp0J/t2K1YVgDwoCuRzS1OwLPwjWNOXQp7rKT+ejPeunMzg2+0uxVv0wlKu
n79hKoG9eauaKM3wOXZrWAFF7rdrC9jJLtAVNMAIOvEUz9eE7BFrkMF2QfA/xOTcuwXUaJO37lkK
/I4nQQfjr6ezgKdEEaA0LgyxXxhTTF0C3SCEF7yyikrILEVFEDgMYmyKomXSHmL2Vx7OHxs58m8/
DM+BVbVO/JEeAusI3nC8lk+/bVtajn+xxBcv64sVGyTW4+iaTwqZBYKk+yHJ+FMCFS3VCqzYEadS
DaDvOspm0XeT+/XJyNfc1HJH9xOlc4MrqzhARyVK5h/WDaTF4Ls0Y88MoUkbPnQvMhvy8RtzsNHu
J/nf61Sp741XwNQmmz4j6y+/IsIxoA3azukMB/tQflCak+SZ9QeY/hRp5cmCUsDEkb361bQiTWox
pOBOw+nCz8e5ERanwb5ATEr02DyKUf4ZBdk7K3WEILtSN98/8nn74bHKoUDQOvBcr4/WcLzSAnaG
aPA+9Q6BKOhEDFDcMI49aYuMzWoYxdVkHY0oGctDSinz2qAd7sOv7SHG4eDLz4YvhDyqkOjU7MsH
K4rbtqzQF51CAOX2dxSzHkcin9eoLsc9Y6b2lz+6uoTdbuzTEpeOwOZqxWyQlgzsNj1+UuM3KCer
261/GtooxUwK9MyzTEys84uhgvzXsELL+9iwIJm7UjkNkfgbcxHA7GbYOebiPhv01yD+TPIXr7qu
dMJ7L8UDwuWcS607wq5n4XtS/AJU1yObde5dbfxubuo0SCpZkAkGF3089fdzKEqTWaSePnW7opbv
0jpYzceK12YGDCDDzvCc3IarT5IWN7T2A3Bm8GA+Jnjhlt1xQ606na3dXrDtr1F4DP6q0S10REiR
T+0t+pf53sN+v038neKqIdA28O3v0s1jhZ0xINXlpM6kWdb6jrR7i+epQtNGfbSC7z1moZhzF2NW
P85a2i8w3GllIG3ECPnumAEgJHLXklwcslolxo0DtNsQUL71otDuVZPt3vCjG0v0kfk4k0g84r3x
vAhhVhJ/XIK04zyBFY5TpXKqxyk5uwPc/bYDBNzJDk0pSE+pYqmt28eTDhv7TLYwSiZ0bRRaluiC
C9n2gDtij3tCFRRIKi+8hl6GNrbMgp5NS7sGXA6AUCpwg+w2RecJT/Qu4Zkpzy666lcolLoZgkia
RaBMJfzXYZU0hGIpX/yhTnkke5ta88JuUKCZu3r3kVd+eaZJdkrpG/pfY1es+ljyjvB9uHkeUjj1
yBWflByeFaSFZjzCWa3j+jgyyJYCtIl3u5x7to2p9YuQ53nfzmEB0hu6hxfMufkdVx98XZeS/XIZ
379gdvTFuhbBQ0/Q/i9x94A56g1st8OmF7kBEVdZcuje2+X+KDao5QrQbO2vsmdxbmSsEwfvaY4W
gxhHbnH59hnt6Mj0JL7TsirjnyV1UU+KMGaJleOSNj8OS2lvpLz/xVRHa0zpIdw1BhbyW8kxOlBb
eIyCRVQQmd28G93BfsmFoUDGcrOTAF3wQo5w6gR2GFyWz8i+nSIAgppa8cUMk/DSJRIY7pGbujBN
D/mIdtBK7w0LI01+VmPN3PfXK20wlJKluyYB4U3I9dE6Uqc4kaEZeM4VOU49U3/JfkPHDAOfhWFz
Y9jplx1hFrAv6r2osWuB1g+cJ1OuXjD7lPp7hncx8grWRTy2kyyMcWB81yedib32ogV69mxO3s24
8Q+/HaYcpsPf/5Phq5xbvu98l+g7hVtdDnApA1ivhSSNUiIrbfcHqd8Shm4oXfL+/iTsNukbGKCa
O4BB7rSYKRKSy7pn+g/QWwc1B/I6HxHXotW1aLr7+qLnFkCxUniwG8ZZi3Fzo20feZ539wwp4eTA
cncm+eeyapoN34G/mhTWxV8NgRzHozCG1Qh174QbENGyb6AfKat74IOtTg+g5pZGTho7I4Q6PYyM
wcLt94T76Z3PdxkjcprGeKH6SuRoOVcDtGN9Sn2Kq9qWCQXRI/s94IvEaHN1g3yQsEFpRpd6TbQy
sIFWnsnFZk4KW8R4qomm6o2K6CeQ3u6Ylk3t1LMuE43mbg0HQRXETfaD/HSAe1jJDnFpIRCLsLXM
jXpOf6bkcz5Oz8GeNK7wAVTP3sWxdQCSQJOQX6rNRI4XTox+9SvkAFc2zMKJPWvDpM/HybMEIU6w
Wzx/Rx4rIaKrdd79MnMdv9c06Gd27/DdrkvI6xUw0lyIKET/ydELOe4qEimCDZ1urOLf//Pqunk4
DDsTgFaf2PDUyt9r4hoh5PpeKs/MwxiZJ+/G3e5XHOdIjGY58qaqr71HG4CbdlgEcJu5hZ4SiG1k
stiawRFTgCucyu2aeL/8scJdSsUuWDaYej/fEmNyXKRD4zDOHHh8rq6eeVlZj4dZQMEe+IeSY3ox
Lh+wb1WSliL6vKJJbSsFAONzSvX1REqUuqtri7l2okeqv6pYIxDDtMGJhrq7/0noqLZL2aHH7pxw
VkBWT+tUM1cQyHIjuLE/ctJc90tK9CHbKm3sTLy3BP98YQpxaN6+ftraYSdTzxm28kZTAdFgbnIx
Ar87CuAnifJvcnlJhooEa1+7iW1tgEZz+f8OszWIpK8pVC8nXn9ppPOVmDtmc24UTXi5EELz7Dvj
qucsIGJ8uA2V3vhzaazNwtjQH45gF7qy/X5i317FyWGv0K+va5Nv8dSJiZmwBp80LqvjMkDahoyA
ht47fanaztLmQzqgk+uplFTWG1y218yqRcR8UkOTqg7nZ6e1Ai+35gHjRnMobcGY1CyVgPpMueB3
lXch6NuvW3toklnf+3gk3I4rCphH4fxZNZq43d5U4mjO80Hs9JLclvdETIJUwaSG+15trnUh2vwJ
ErDt0z0mcPJlu9SQz2KLvGp8rx6Z1S/HiIi3EHVOsDBjHGSdY+S2yqwtJ6WRpdIBGnASCas5zaqv
w4Ke36a/Mn+n/1qCI0H1n4Ll2zzd9Uvw9TbwxPgBSpvYkw531NNq8O+TPhxj1Ec2d+X/UXExAjRK
L7VA/hBhj8ooS14r7az/E0hrcH+KvEqgbZNs+aMSfzhuyh6aJBDY+khYupnII9aYLQg2kMeRNbcw
hsvWh9CqBBbpMsMr/gVVnRsCA4zMeysDc39BbIaRJ4NULP4I3aex4SZPEuwLgIUIoRiD+Xdw/9mu
7CDwleh3hJsmBvUDUdfddKqFfL+5CPr0EZGNY0EM9XDeKxSd+l3O1MV+jX3Niqc2eiB9DFEmzEfF
CrBbtlgnSgsm9ZY4WI/23JQ13yV1azRshlVXZvK5/AtGRLiOtgWakWow9trUyrEE7rt2RJb5cCz6
2Cz6DrG2Jz23/ih+HKx1SCBCOnzBaHbYjjV65lBoYNtQun+woRS0Tz967V6aNJoK8RU04VS8Fysv
p8C41c+v3Pzp7DA56hRFAQT7lpOiAj+neqETU1rUg1LXMD0ZEOcKa1pSNeprXE1TjlMS78dhhXOi
pdtXOjiI/VIdrNgO79iO/Oi9q2GiipS9dsJj6CZqInnySjTEzo8Rd7Sp8oa7Ps1RzP9xVXC1DjMw
IITJqHVZQnIUEShb/waHscirJZvpD9FLPDeW47+KmqsXtdPkx2ElW6cuoUODlYIKqNIXQkXiQsY1
tfMLM3WAvcolQ0wiVgRYwQJsvsHNnNn2ZHOZDrWNU+yrGPQ5GTygpv2Qgs9GhUoQ//t4HFytlex3
jRI/Szamq7/qCrnnMCrczZERHuY9MXTUj4uVH/eteK5IimfK0Tqy/9LXp8cbVls/abjlI/ekOZdK
WYs9JI6W4SNfwP7p7TP+ckVZsnwtpm3oppbvmSao/YQRAJMgxWvjovDGRl0InAraWeQ4sAdXcNEk
git37hWCSqsssrV8BXiOAjLEyjKAgewJF07c59mc48fbl7m7v61Lfu2BFk3brdoeLqPgy27cXpUp
RWfVgKYvcuCV+2HxOHeKLs+DZyfzSrpyn6c9xJNk1AHOwNwatUl0a8VYLUdV2LrVpLCobtSn8qbX
3V0OgzvMy/qBuSyMmgyV+0Fo7U1z2NpNnSig3eE8JshBmVdgyMxFUib0Tg2gvHYar/Ln3LtF609Y
Vwwj7MmofThmt9qByX3JotAJP+G8YpVxFGIMo6P/eaHjC1uzX2+Nlj032gILy0osCUf3/yGjGeRV
p7tswZ/CQhM4f17RILIJ2DTyv9rzvMMgq5Cmytii8r9f3EeVgX+A4FP0TrE5kQ5AuFlj/8wFgA4I
5Hr9elR5OFcKy73GQs5Bsc5C1oBNvWmQAt4B82PhHJjLub1JOAJQxKwNrXtJJdDzGpKTF+xFaLo+
h82uMmyO6RQjvDfscai4UhxJjdN+4RCvKEXc4Fh1+BqwXjmj3rR60wdIf1RkZL2bKPG8VnQcxWOS
J+DR5lG55q7UxUJRnrRd+glcFS1PHeI13KIbZMsW3PH+aKD7sLM/NwqZBLMY1tvLwH9CcpeCUGC6
aK3xWF4YGkTRLrNN3vJc1S2MI7c34C8XMjGmXGTEMG/2H9kCcjqhD7DWqyjJBpaC53nWADROls6a
vDjQv2MOze+fHB00ZsQeUBKed4x1RWMu1bCwkX2bHmioUIjSlh+YYh+aPCNMzd+HHlzrS/z0mQuN
Ac+Fz0rRz0QNXzP/cgeR/I7sxuDmYkN9hmaN3XGNIQLyIlOKVvWVsi8D7y6f6tEzEb48B6G0ipUY
fRiHwBrT2G/FHJF7QtkMDvkE2IrOitaSUEoK+MG6tTLZXHU7JFPX86NB27/+bv7biBEVPteeECmM
SiA6dPHAzTtdAqtZf+rrqQ2+DiaXkydWkQtAxYw0Z2OeyfW+tCjG/Nymdybq64GQvCeV+Fj0kmch
nJxaB4TmRBmqm0k6ESeYD7TZjlsOPbbLgrZJqX5ZuWPQYZtn06mwZ3FWp2BkxIBMTcMNl2swZMQ1
bpEal41N35rpwdSWskFDOWsAHE8p6L/5w8Y2KrF/quOgsfGveLuBaC56u+0QSOQqHYzenbN4PmHw
rJLTsmyihsWovwnbQCCYR+qhdh1l5M6Mw9xN084kasOXHB8PJsCUfnd+9NwRWyiM11WhBs5em+bW
WTy69gLioEYWyBPsXhCE7PcvFXY08GXI15hipWA/BlHl1eU1mFIAOZcYxG3GCprYF6P7RLmrDONE
yoej44vwGWoocsnJgFpZtYpw6v+g3bjGM3R7i1YUd+ClvLhxXh+Z+0fNgNmlJHFGizK8kQVvQ3jL
0NJxTOh4C3YiDGwl4FxBcL4BdFwcgL8Ru4NMXa89DFQx8sVehs9YMCJ71AEan7rK3dLdlVd9YdUt
hQsi2987FFaba2bTj8EwpK2za3WGP1I9oI/FTLxOmLWX0RE9E2SzvH90JsBSPnIPvuwJ+XVhrnxE
amKpQ5msib9WAV8IxYsb2p0rTKJ4lflrmUy6GTGj5yPfGMKJJkFW+FmNQsugVeYUDOhh7wXqe305
hm5wMYo1oznKNvFntbJ5CiGP118YZk6MPPB+hJevTaARtqK5X7Wa4R+Wqulo0iRZj87wpSVvK6UZ
krnLNuKtXOv0zzkucljwJKV0mlsZ/l6EssbwPvhY1CsCKFibsJszA78EPePHIkneWn88ni2jSJxI
0/uVABnNQbIJlW/Ka9hizczW9pHEKt0n6HvPIvk1MlMrT1O5nODoT7ZOo9A5UlYBPr+DOxLRvL6p
ypg94C8nmDRpb8SjQd1j98FL509GmPp0QooD8/1gWAwzkvNbHV7na2LXqPEyqPlYxYIFuAWGgb4k
zVxow8bHaOyY8lLCQe+7hv4XnDPkPmuBThnXbvxtj+sLQLr3ycSKVB8BYX9232b3c3IgXtxP9I+i
SjOJ9CY81+4e5qrzloLamisShMGBqILqyL+GGqO4c5kWeMfgqNx6unhTHbSGaTK/VzJXa9huF7yS
Ztp5sA34eoxDz5KTUfHTE/hZX+tIUqedmSJlBr/e3Qwiomf7a9qv8KByFyjTC0zRC7wwg/dJ+pr2
c8QV7R/jaXK5tAn6WfOGlVPYod8/QsF1BCX7dWywWLzmrpkwk/JQ+qkWllag9H685Us6HjbMqE8u
T7eyL8XFDiHKph2NbPhTnXipUo4VvMb/ds7NMQtmux5OAgzVeOHxDvXWOUK/64vKqNUDTc9qs6Gk
/PQ4LgMXi6JQYV2037yWTnURntBNWVgNIit3k+T+uBOgjUwI0lzQ2EOhqFLJ4W97W1FqgcChedSu
kys9/yixjBT4vwiiat7F/UywYWfVHcJavcjDvC/1qIkbCcDano2RnPaYaQKF4lxf5wPDZY33nWSe
zV9pQGh2fmXIIGMc6stRitcLr702hJbmFLN7G5rpA/uNquh16AYO92nsb8k1bXNxu0PbuM5zUxqR
a0h204R1SBC4lta6onC3IIScG+5dsroGggNaKojBr52Wl0KsTC3QvAgWeVjH5sjoqa99HCSJtBYk
xay95Kzud0sdcGjc8/15PWotZy8GpQJb1lc1DjTaJD76pQgd+SZFfMf9GQxxCKoNAm4mbNRnBhTR
CU9kx/BUDcu3ZGEkDRiS98wbH7aiB+P9Gw9VGV4ZSu+o0RhoW2Fb2yZj4cJRCk8G1MGLPfSbg4td
coPpeUP/h7wi901qusApNJ+6KBcB8wIu+7Nh5kt9Ur7s7TmNRnZaWiDU9KHNdfzwfN3OYuoBQwne
2hZt/IwX/zIJL2aM2w/GluaFiL9en4fi8Un6zfk7aFvjpfatd6CagT51rmqnK2HxEIIkBPbm7sEA
nxfvgchbR6enFHfgd2PwSIgJm2gyEvZjsru6l3LfAmMnxzT4n4+4XQluAVouPVM1yXJJ+tB8lSfI
R+iDkT70GED1lvl4mFPmB4UlYlQPM3TiWFgmyHL9+tRcepxOERHymkeR8g3TKa0cBUve8jlKyMNL
4Z3opZbsGkJIEknRqpjy9g0YUGa1OWhfobQRQhPPQ4jRxxbCb+d6h5OWxc++Rx1c3YQKaQMDDI8a
MfeZuIgUSzmODHe2XT1RhEb6DjNeurlmW/NfQP1/J9NOaJYlms78lliqM1tAh+8l6KT0UPLIi04K
BVQ2K2BcVEY2niCeVnszN3vf8j9jpHWgjVLFhpyTf5pMS89FX7lI6VJWo0RGfJ+yudk5vYX/Diqs
PD0NUkOm6BIhdvBqQ6DIqt6rOBita5hHNUseDDmq8qGJzOFs0mUkNmEEnR9bHRQV8n5Qe2A5W3Xm
6nPh5+IOj8Peix+YM+mdSc3FjEszyK0kBTWKDPMMlDNF5uprY6UfhOH3+Mwx2ZsIcr46zGGc5d8T
+KuN05K3nR1nfZFchiA3Keyw/OgACe62+zJd0un9lvlLqHqZJyFuUu7peJ6gxytg1XNnzcUmT38i
KULzJIj1hOcTo4ZZjOOskM50jI08MuMC17uyiQXkhr/JGXFsaQh1rGjpVlCgOituZawXOqfWgpRp
esX9zBPcS0cXvPaBi9mSbg6qGYVAEwyBZcXfk7tP5qz6W4+ebIjlgbTtjs84hy9y0+wt6WrgkK+/
5AB0JD5ABuCK1Z6vHL3jZdDdFzMidR5JfLHoUfxraPlqmjFNPdwGJLHh+SrVYx1eWYf8Mpi8BX2C
NfcR/h7nrYa1hmP3xlVqOcNmlsHYzOmu80cAu02jpEzPpIpCyAuAWz+EafmxsvcZYr75ow9bF6xc
rIombwBc1mLNludqOhCM0txPygmJw4ynRU+eiqvixuAHBW8Wc6STKhzXxKBaUcz6LpBFSELQLDWn
Qoq+A4E5zcVD7xBC6FX3/76GB/S52r0mvn5NA5Tukr2MvU4deCAtrpLk7UnYs0GmQsrKHuDN5cc6
Eey8iIzguujfzfhrSjEvOZyVR75l2+AWP1W48RtEEyj4Bf6U71N6zZmfypdyLi0xbve0nTQQzodg
PAl+XIF8nIbiMcCiglBZKuhJwr9Fe9PZk6NZvE2gxig8KNpCJTKMvLy+qCsnZQebFYQ923k8cMQ5
/FfD8Y7u9SWkHdwHMCvPN+ltAWBho5ro+JzpyIxKYax3nZ8ZDzvlOWYA8WvBb164Vm5lz+jy/vjf
ALU6toKK8y+TapmAdBGv58qzLU1OGGLH64CtqDjaB2m72fArQEpu+cYcbDSi8bZMjcKpR0a09rzh
q2V48X5QfhZLPdf50egz3wn7FF6dxPvdyTJd6HAxHKrAvsxCTsSXN7yWQ9rKT3QmMBWaudo9Fev/
GDeBV8MOUqNgV9sbJaURBolyJiJyCNwWS7aer9dwpatBpPX3B/Cz9Jrv5VGYB7T8elnNrxLhLTx1
yD6eUPRo+ixgj6MnFQ3H43rxvkXeHfqaM/7OmPccqCjMDp8w5/9pQtcVh/rW770xhT0sMcLvC3H/
6zTDMNzv4lSdaqpx2WHZFUfCtfnS4LZWwxnjo3PaoJ9cLgjRdND2L33eoUGubJ9Tk3GroySQZV55
O3WBvZlzcTw8g8quRkYlzopXQDTdZ1x++BppmwF5Fb90eN5ua/PGIN3jcuYfUzNo38NutXe+u7w7
ciIVmgxb4yz0Yv8VjY12+JoeBSTYQmDKwfSsmebB0oZ30wsAIQBPPUqEmzAFk5dp+fuA4fwE7qJM
zl70htT02EvwDBHhKkr/7Jg9+2BXbjGx7fnlnoh4e/NLyGCV2VM++RxjjdjaCZGZHYQH7ei9kxpO
f5Y+IdkvfZpMP7wOQWEP5q+S+eJ6XMOdwzK1/a6ELPt3zrB2ebXWAIWmr1XkS882waoEWVLNqtmd
BcUP3JzxgIQ7Xk2RPw+Epz4Ryg+8Z3uh4vxDsa1giqpBjXDIB7B5pXTaydw0+vjR5VxYQK7B0d4a
M4Isp1dAK9UcjhzVgxdw0C83Qf/ZnbybHc8DFCvsQs9q1LUzhfVzCHOokjiX6iN5O32QWPEdGHc+
UrZ+3tfnESRopC+QpH/e4GY/QEjMx7ERKTDW49OZRf0G4XApA8vYk8ZC/c+J9kgYS3EIuX7vXrNK
sBbwAKjXIhTQL/6oXtmtu0tzHS0r5sdMh0dOUbfISicZ2yi201Xgfm5NZo8IsxE2wLX30Zg7kyuH
BY/YUf7YiKkgvhyeSD9MZtpcedIQjWIef0qpGw8k4ETBGSRON3YplJTmsecWpLENmffDrQMj2RZp
5hLOsynLR5mhWLM4tarKAOGh+dZefh2c6slvy5qQ3EYgocue+1p3OjuK2POdonWQp6hGjmiyE/zh
NV2Jw4BXrsQxQpdizxLIQ7yOxIqAHR7DWl8p8Bk2zfZe8P4mAU33vRio5GyCakKNUdK3TiRvAQT6
+BVwTESBuWB/p0dezZCCZY907Y3aPlMmv8+u5vLn6RKkE1j+Zo9zMyxRn9rR960GrHzmZCELBX8F
OYQuI9yWoG0GL4FoU0TVRI7DuAQtLWRsgWKB0UWqeesL840D9kVsdijGY+mO6N3pyy7oX7eXTA+Z
T6kVnrBfkS4m7QIFDk9/O2Mu+jYs0LuSpxKpH570twMJEtxwpMKc9p91cq6DEUN7zyPSPpZeE/p8
LSVB943rvdB2XSk3+JJSQysI/TtA4veJINyvIPCB7L5KpYJo1GkzC7qAipOHU3n7A33tiiRtEcWo
tAyArYgTlwiU67MaYqeiqbTzfnLR2BYMhMbdubuEdtFZP8JPstVPdx/NUCFmXnWhxlI6BrxZ+sVC
XSaehzDwE1LCzsqJBPKKJmOvdjuE2nFtXsxkrFJarJv9+SUpZWbBOJVO/ytTaoa6D1/g337lsxN1
jVapijpOVCL9AWAqX0nba457iEX9fQjFRggAqh4oC6f2T2CyGdDF22/kJO7lRUb71BnvXRKEeoiu
WXjhFw09qIhNnlIYGuu0hj/9NunpUi+N8L8+dsZ1cQrK3DZZ/pTIyui4SrfKArze1TJK2Xf2ny7I
vdZzTP5sJv6x4+BNbBE3Juf/S7Ic6M488SEEdy/mtiuNunh1dZtdhYRyXJOn0/tfKNHkxKAmVIsp
cdTzNECkPJGSH1/mh1mEPvml2u6VRwSWHVKDvtvXAq4zDmf5KhLfHpjjr/FUrRDn2aErTqbcKmYk
w9F8tOV8VTnWAHpNYc+g3CHPg867q29Gu6D5DgP+nkPzCGhhmmheCHVuIWAkoeHkVl2iMrZJauxg
Hi/Qy1HptbKiBkQnTDBgpMH7I/cRQiO0VV5FjjwelhamdykqpsQhUpRs19VgjN+15Ntw7xIFp6P+
d0RIcjV4gA6VYKIqSKZS+hJ146K2DJ+jNMExexOd+pbWelNA6QJnE+RNjI2SrSAPiVPgYXWIEVuI
pnREFRYwE2i+NUcYv5SLFJABD4tr7E8i5RXeKntSpREFlnNuJEHXdqJ6FCrMJFJ64Pf6ncqHErnk
NKnmFqTrt0iRmeO1349blMfsCHBZA+hq8Bb4woDCSNsB/mLoknIpfYQrL7AV4F79tlbBNSkee4I/
rS8jEM2ziCuBoqsUFt1mGcWDJ9v1Gns3cbD6Tx920ByUl8DdE+uhvHuZlNfOnviRuRKxbwWd/cld
eSt5GSgO+hiq8DJSo7XyLdNJSCAj7eLYtDqAw9u1YzLF3iDAZ+zTqSILNr2UpGc4Nu+ON3YUOzUt
mZu55uB45YGLxt0KXqGSVjRA/smKkTQEmtlyAFocvvL5LMhZYW1HSIN86mDgV5njb4fgD5LJcD7w
4ObAEOsZ/ZzADWiot1aMIuq+AMtutMc6gr31mbIi3Oijl5ERMPD8ts7+wB++vJKkTOyk9fi/jwr2
kAXqKa9pMZVT/8bYyhhg2bEU5kaJGVmcAMAt0pRB2YLNgRCfShz+Y8fo5qCAzVGmh7cwnQc+u+BZ
lCNoq8ab4cP7lC/Pr704amxztkwce4HtdyOrTFeBFYfLgV+FJmMau2ERIRw0yGYjUfuezomhnyaM
JKrpaz4AF1U0kx0GwJBtzFKcXzPuTrO3EuO7ZCUrsbjYScHS3Gnr4dz80yCpKHfWl4ZLIi8yRj4/
7K+KIoLYsmMvwcauIUsMh1+0PTlji5fhdVcJ1swgwgz0kjYb5PsQGEal2YR7v4VdaYPTj7mEbcAy
A5wkZzvMlh3Jfv8FhQ3vlYuNeoBR3+z2VbCoI700uvk/B5egfrVlDeEE3mOyNG2FSNglFwDAF5Sp
yPKAXvxwvakRmtGN86bRbr+QsDVOneoJkC9x1mNQLXvCvqIe/w+EIrH9i9BOeJ0hudRT8kNYaAIv
sZpG0KVIFBrStCd00bOBBc+Kc9fTZWO55UoBfmQZBaSe2+uMlFuzH664nOGgiTkfKJxzN4xTIAqc
WLwbV3rhG0oN+/8X9vGtkEOxGrGOu9f+t1oNIl7D7L9NAhMroJNsP0fqRyd6s6kzjJIyiwZBOlSW
ZrvUNBxdFfC0PEc8HUnJwMHCHVsNucju2WI/SIsjUWnd5ZSbWPZn8tA+Rr3Z3BELZ7BylGjcU3Lb
P3STDZIe6zju93vnmLAc7tGbbNpYgZQlNf8U23PiI2XKhW46KagSx8GzLuYDmh+H1tYP6Ch1CCW/
yG53SknNRPpGMiPI6gX4pi+gf+CpIyvkSg5+iqGj/TMQo1+qHhSprkbGEPuISUyC4CbUFgG/t7Lz
VdRDXbizGRZlKCBDt+xCjcFh4y3PasOXAcmNOrgfwiwtQU1frSRhAQmET4mSmL2Yp6ELFbesKnzx
qlOF07PO0F6uCzUXFQZWaXtY9fbBPyjAAMkM/Lope03DoI8v/6XG+ZPBzNOAaiZtBvkXqaokxe4u
mKmeyvVWyCqhq6jj3v0EkRUWNvA1V5WsxZ7glgNwIuKK9YI4w4e/oG70g0RplzGOfTyO8dinKFMb
XIARP5+oQEiGnBP0GZwHUHxB3armPI7BcZs9jOFMCNfILWZiM5FgzZYNaHRqJguXLxYC6KvmJVMo
Dhf5TfE2CQ8Hmopp7szCVzgcybYCP4oaDVW7ER+m3iEleKx/t106O3EwEqyx4L4z51RAT1dAbM1n
luu8TLV5iJgOmXHqCAyek6HhndCMzHpn98KDompD3ks5F2hDwWN7AxedmwH6BI0kVQ//DVkN0Pe0
UxINQ2Au5ooBQp9vXLfZXw5PTD183vJwjZyOq8rv6K/cAW8yB4rcSID8by2/gO+9ILPOiYyeNXiZ
BzMBXIUVKEM871ijL52CUtgiyPyV9PYnBnmhtQCa4S/LU0U45/Qs46sNCC+/nDIamRQEdrAmx3Si
SGrjhS4LH750f20ekrmGauK8qs8eLh4v9fTaKKj5ClbpVLm5nnrA1FGa0tMkDhze8ITzNP4Oplfy
/ELqqOht8tsJWPie0VIzBheVVIcjenAPontn4QF1jLTlt4w9SIcJZAiKPBCK+vTmPIlwgW9DED2q
Gm95w5hkxC/HGkCUXxwtuGJ7V94URoJ5Af4pYZgNY+6+w1h0UNOUbfsc/L7yfs1LMaOiFistT1uu
K1YwKrWDALDVcDParV5pUycxtICQY0MDIPDfy0sNQ9EhBL/y09j8HImbtlP3uTY4TGJhpVHnRsng
zIJPn3DsDYfQkgEQ10AdkUns2yPs3r0QG5bg07otb2qCrZYZHWBKLWTEpx0UJ+u4DGKSrnnNpoX/
nYZ2y3uF/0HzW+3WYl241ehWAJ8+lbEpzv2kD0xRBdra66kMzqQBoAro2DS/2vgBrY4j0P1fjPpU
0GZoDJkGg2s2omgp3WwDkwUy0d5rNjbEiaLJZoNY69THzs2Jqhmsra4c1fA0gFYEFDXoY0Usn8Bt
lwib1EkE8tpaEH73i/2wcmdhOLfrYlKazPzg/AYGyxndMWWoKRYLIFLuwvwoz6w38oKV/Hop7glr
vl21dwDrZS25IaQdbxaoO6A3yDglfoEedieyTdeVyJsCWppmiF0GzJd7h98Z6/0HYBqBAIx8PInX
L0/32Xc9cFBSwhWmu3UrONzGU7zxy6nkhTXJwyrPNOzrJIFyoigc6Je/zek68c9lwPtGxjx14QT9
Y1HwjEZXPd6dFaZK8V1GUfe/v8+0VCt6Bx/ydDgz6646ahmRxFAsk8itkZs1qhWL61AmZZeracqA
2kR6gdYNvA1OH/dkHuwsb7uYD5b0ESGQISWXsTv8Ri9PwSvlSaH4XmJNTVWkQkoZiQm3A7M5jTE4
M0q9KUevDGxQLr/ssUeXBj6h8wKP8zkEMJQhPGzNfElgGuwpgq2O4zcDA6mfZQJ6ntnuedfsai4s
4GamFfIACVyXJ6JRv2uJwYAHIwIQWX4wx7oMwZevh5cWoMdCs7xcWXimXKzKukEFBhHsgqodOqr3
9UnHUggKyeZUtYA15a6tLB5pPBYV8z7Z3FafZeddKlDtMh5SQrGD41tJRuY5BerwIJ9QFcraEi2g
ckvjWFAqhLsw/52q18lni/iVQ1wCGaVumIa9k+d9GOTlLHHsYwZd+HB/iGGaEmwcIj+y+cpIOAZg
eyV+arPUMU5inAjlKCoECgFMjhK84WkRegmDeEFHE0kkhAkVZRJysCtqLIgAMDDVXJXjYicnLfFP
EToE2PC1d9Y5yOCsnPhVoCAyFwv+CTxH8l7KWwDRPfSQPiLgxSFJ6JtzNzrZg7DDC1kX5avPJxpH
jU0EF0Gu1Xm7w3yDxUKIXBHDP2VUO+biJKh9typ98kpUtzjhgLEZv3xy96anauuGY/morhT4CWeE
Fkvo3oPq3yNgRzcYSoaOKJlJTwCukJlHDGbWDe36s9KO+Gz2W/+AN+lZhMD1JmwJtf4+2YSyrwDC
w70w8HWyAvc8UrTG/A6rN3V0hWXlRuNUmhieCuVyfwdcN69ErqFrZ+GbdGuM3hHEE6T0igqX6yCv
h2zjwLoTjTtxXFGqUw9aEWpgns+bpxhuCMBHTz6KYImm2l+ymar07vtdxd0tNMOWTLOhTsBP7Kil
ChAXray+nh5HP1uiW4oS6fz5j5HljKo6UsG8hCd1RBLCRKIcoJ8Gl28ipeSTcATs/zymFgGzDmtZ
MxyzYFKAi6qwEwmyWRT6ykWgB+CbuB/BgOzZKYfVEMR/c3wec8YgCmk5OfY0NrSQuUx1KudQ5Avg
Xtv1rW56AsJLIYLm0SPdHwV0gs3YiAVw73UzGzN1D2Bl/yJQeu4iHE5dGMxpRqoxZpNBOfessxNU
cxlNFD9kz2MLIUvApWkDt//gCmFMeq/lDh+USg03U49ixb/fce0oMnbXz+a5syZMjMs95iYDYHKW
TeIZp2Zu1MCE+PJUKfNQmfh/uM4MSH6kMCw53ofcXzz/Xu6VHTbf0qIWRQafjaCTg9aBdx3W6Zs7
mIMzyRrsW9o5fvdKyjKiKlvEAo9CUf0VMhYxvNYtLXREytfgwTK7Sx/1yGWjtqQDw+HK1l6A1SsC
3yi6nT2QvQ3MpPxv8Mz5IhppL1YK3f6hB9F/RaT7WXd7SaAZIUzIpEF4tkkpRNo/pqEFFC/NzUeQ
3JNhQirsdgIgt4ZDnem/pYs6G3zJww9+xUQ5insyl+XejTFj89JHZqhRBA8U+QCRKiqh0u7SWObI
HE0t9KCsl88kdC2JX8FM0k/XlcX+8Bw1enh5tB4VoXOIrFQdtQF4ApyFeKUK3a3BLukqNIOqtOqi
IRMEPPq3wv5kowxpAXi7zELgcQwn0tvEvY+Pxhy+RL2n0nPzqBHlN5Lr7E6Btf4iZ5klRKVFU5tj
5aldVTbUqTFC7y0tj/pa2StwzbTKC2n7q/cfL2lnOniltyd5mBqzNKk0IOLsSfUwihg/halvjInZ
vJLAetwl36ezgtF870hee/QLa0MEvDukXTfXOt7KYsHxFkDknrqlPPIb4fD61hRvt660bDzaGV/w
OUajs7k1hdmgc/6ipItnM+dHAAYOyqvKHRoKpAs/0HeUt05GB5pBN5dXwi9sfJ6MHmqEVJdo+FLG
DZvaSzP2G7yfn/Yy0S3zVb6srw1E4tjL5cBYR6WRScL6FdvpY3P6IJQQqEhHGUc/cZwVV0PqTWP8
qwAIklUopBAXRBzidSYcoq88D9nfPXetn0/DJJH4gEWhzUvJBdAr+eWacsjSVI4e7DX3ZUtRgQl/
O/VwH3qmj/9vAXONJeKjcJI0bmhTC9bhMKd7hRXtmJSm0tdPEg+UlUQQdBn1e1JfA7vtSRlGsF4n
+LP1C9c+OyhGBNRHL1wBt1n/EA+aU4cvoIZvHjc1C/GZpyWxvMZdBAzijdj1WU5UCIHRUN5KV8n0
u0KA1Ozf3syl44xQs0QydUlsuyrTLFzZAVHhtpsdbV0LXwm9F1udwCAey1CjCBHvICfb26ygIW/F
so/oHbT7RTaY49lvP66ZCLSg86dR5gSc0xfSL4o4x13AyaxCJrGEELg2tqk6qwLncWjVA8ulMDz1
Jz6cQ+lB5MdlCy69XZyR6I+nA155CwmPgBOOHkiFwc7AO4i58ce5u3qx04OM5juCNvDJlqHu/ju7
psUfalgdMim1gQZCAKa81Jvg2OspozgMmnL4Ha1AAFReRM/qTGO/IP9Nn4R4ieiSeiLPRnihSYzT
k7T5/CBLewQd+afjLwDbXbh6QynLDB7hI0PBhaHsziM2OvZSlF+BDrEBlsNH1IBojfC5mq3oyjEH
xffAVLPPw+RmwlzIXgUJg+fW5OFvMUQEwRWyRSmAnbe8NF3mZYlrpL47CBtAjllSktPcgnp3jXoc
T+o5ZzK5j9t0iqVz6m5geSVYZ/MEqGTYrE46a9lOacM/D/4qSWLX5/GVCWClYUMA/qsCeI4Iuh/d
G+Z+e+kyDSMzgg87y3CW2cAbullTMkPu8EB0wBZS8XzOJTHOyyXEN8wKCtLhNeGKZuT2qqq3ZoKQ
lv48k2LDid1YHJEkfs1bJ2UGwrkhYgTt7xc8X7rZV68mGCa4fZd04RVN94KVKqFdEXxeqfeFM6OZ
179RsyOhIg4PNMZlGPyPYGgNv4vkEZKv03TINm603c3IvJTdbCFA97iBSQ2oUsKDCdaCl2xw3Vbh
wNIq9meivLNubzb7D/JCKVx/+HgxsN5xALv67KeLHYvl23SLbo2JSjocMi9WVViMOUbB8lboD8mH
be2DGhwO+NOI6ozkhv9i6X5SAQTOGjvkEXZVQpR4ZO++z+bgwSJqfzvGWaHN0HN1Cp7EuCa3scF5
I2H3YnshQ1G6Jl4j6LVegqpvOKls40UAeKXeHDt+LMV8r08MCW+xrmS8d6RjCDnlbUWeJLgMASKM
EkRoEHsihWbjXAWl1mBGcWr9lg8lSNM73hvT5fTzaKjOSwqtISlXvftsRK4dEoATAYhuqMhR8hRz
H1Jzho2/WHkWfjXVLxijX1KG1UVo3iP7VxazXkJvFJq5G5CK3625XcOE1js+YItBu0JDTUPRrpch
jf1JUhI/eUt+t43CoYe52Kjca+hd5Ln5NCMjSJ6XOPuZRxg3dJUxEp9dovfdzAVxkEjON83wOI+g
z/3yvUaeuJSxY8WiLJ5J7va/akCYSTmg71sXx5F/vwURFqd6WOf6ZAy/jEiiYVLotjo78FYDP9qZ
2PZxqwBfdIyqVUOpDx5gPqYNKFEsGSWFZq/sslgiEuh4DnRkqYjryquwsWR/3XyeIF73OP4nbnuq
IEC83bXJVdpnaVFu/E6SUXcq3romjAQOe0o668G4pXenDzqDfQTUbJflyLNujykB4UtmcKwDLSGR
O3yki4d0kYcK1zaCGrGhEOcqxDtGFeG89XH9KCXtdvsMvIzvo8p/hrijxE4tHYt9fAHFIvzz3ii4
MWj2vwMdVrPkzbb4jeInbXrWQrLZ5nbs5td0r3I1jQmYv5NmtDf3e9jdVvkh1vRY9vp5sEobyTgs
scRy8JNtZtG/1h6uXaWOCdJad2yeX52wZRlKm/Wf8Vv9S1E9khHoPwa8ZZcJzamNOwzFtVQ38ERc
jt/rPW/DnOD6C9np6/iEgjO7KOKifuOGMOFnN5O5YfO0SzViKSCtEzP5vgokWV4Ssa1M29s3bTtu
d5pQqjTB7idVDjJIRfHcCpy1O/fdhjiWf6fzWVE+6rcm4pq8M7ovXci4vxeX60OYSCWmo5RlAgEN
wVbSCaP6bC2sXEhyP3F8McGScAwt4hg3hLTBbY3W0O5KqasMzP008jd3vH7TT2Z8nfy2UZpOP93T
GKoBokFMbLjSTcghmxE4ceqtYkDJgJWrRVMi4pBYmB3BIOSze8H+xjh0to6cALLAj14Q8zngxa/m
yOPExWfAzOVuiPgBthk594bsr/hFm2yIrtbKaFcrux4tQIRjB5KfajdIIxo8Z+oUORRFTmrcSwrm
IrypAPjQGzqZGHclTk09B+92J6QEdQ1MIQUb+rbL0yXtrLkD3eAZ1DuuZkwT5Pd7bh4Vc0yvQ6cE
zywyNAB5qcmcZ9xU98yQYyDW64dla0KNcChHDfCe/wfEo/ZIEK50VFdN/wA2oZU6DO+tUeyntY+e
kONmVmeB08UyfnvGPPUrB9xB2TeuoQivHcXY34gg7B4jLJ/FRz1BmR/7Mdj4JZJUxrzXdgTuohuN
YJA2FGfEx9D1ZjSp8TFUrKZhqIAUBPdN/yoQ8+8osvhhw/nPFOgOx9JtwAFzNRXirp0tqXET6y8n
ECw5dz4gjNR3sicb1WZQl9sn/h7N//xgiAw3vzaNCZazbB93nZDCxdVpScNRdUZZ9MQW+c5tgz7a
jSvLyv6QENwu+rWcQM8prFDu7kdBfdJtZi7ozQVbCtLZbTDXRjY70SpeLc5/ZBfs5hJFEVmBbwJD
S0CmfZ7LUt6lxQf2G2VsbGV7kQBg571pvuhVYfDVjFdFycvNN3KjkT+OnFHidG1cAnylw5AO3OCs
n3q43BcovQmKbp+oSacmEqXrxyIz5JjcMzEwZrYcrpe/7eQjt0PRA+EitVtyRJ9kiyKg4jNsk5Ta
FcFU4Ge7C2N8i08QEN6fiWii9St68KVrfWvc3f8b1j8xsjox0SvjXxLLDThDcLYkGbt/3Up1b+y/
coU3u+/K7H/8w1Gvc3H3hKy4pWZKLBIAGUd6dwyFm1fThKNNgYPbxp6sFrIUqbP1NXnVwQdrb3+r
JZQecpI+7r34MiFcgivXckbW7y4kPpc0pXwzCds9e0PIiGU/2s8gaDJUouw3KslybnAd/UlYfRIm
2pqBwHp2PxZyD7NNrR634eGr71/C2QEmffzW6NuSeTOleoFqF5qK3yiGIMFPUYcvc4Fd/xR1EQTK
y9GnDvo8BvKK9opMP66cmdTykgRYQ64YQZxP7NY9n11ELbZ9yOpPtISHv/pRjWYFYNmrqhU+AMI+
LyQbGDiUugMCxxj20pyICYD4EQYfGLHExGyd71vs+DOL7tTGXp+1NVpFHBLiYxOoBXnxrx2EIIZp
Cihxx11PS1MCM9hkJI5E/9s0sMgIFnZ3IERkonZHqqg/uC9ttHFHDa9v79r8lXSjqrMSFJPh8ye1
92HyS9f5NHLQvfmeCGbQcn+yVxwyW7gaE1y/ZfvgvJCaRO8r+dHA6qHrb14PslYVh8njUhTr3cFY
pAlQuKCPZEFn3dOX6/tY0x/TmkbLZ5uPXSl8EIdYadRCToNvTcDVcQPYjf/sWmfX08KVc5oOMaHJ
Nvnt59z6hogHzNUe2ku7V+o5TBpgVgz85WAMad3xbs6LcFVvC/K6oA5W7yfnzhDKw22H0MK9Qp4J
T+2uWnzMzTSTNB4iQgRet+9GL38HvcChvGnjEZt4Ya9LnH7ZdeiL5h0d3cmMT5XteWROdIHqlwVI
NKml1lUZMbUIAbgd/j4kxyq3M+pXf2n+LfVWldnYisV6NwmVqlkQ83BdcWfdexUfg92blAJqveMB
Q2ERfgFnqVtEhJQ2faHf/uv8WQbYICRxUmCJ9bAUamjrJMJLuuqTKdCbtO8jJ9jygZasOnHpL7yT
0CmhrOculaqHgS+HdGxBOjrr9IByKI9pjpr/47N/mwAgjD4F2DoZ9nALUhmsuD2HUUyNXg/f+CEV
0HajVPFwP1oclz7RvDDeIdT10taPw3FWdY7lkCn2WWTQnrGLqmdqzLdz4mSZ9njz5Ds6v29tkPFz
81ss2NhJqjeXhl2kWHqZZbGUYYLHZwsq8nPPUCOb9zbS2jeXY1/uRWEiCZlow0YYho5Vz5To4puX
BBdYaZLaz0aoIYXLMoqmiORDx7+aNdJk94R63KC/Dl/JnVJvX7qHXK8o/+0UiemuZtUUDNcbbi4Q
7vU9bgM5Yq/ech5WtR1fwNEjb314Y/Mx7aPzjPDcEiIE7YIl3Qlzj6k43/RY8s87581nCoCbM2cx
Xp8scmp2Rbq4XFcVPMMT3kqAtLM9h9Tpgi/S4DmuAEp8BPisBLr0I7aGMYrAg9wSCdtvwsrHo4Ln
dR7ERRVQorCcaqM+tKqngq6dq7r1RaksTsbs7mtcqPSdoMWPlblmqoEFlxAYZBSa4xhg46mhOy4u
g1VnkWjmWth5vPIr4AXO3KmSZsbPTzYwcb+6/BU9SEgkmErmpto/EGSt40sy791p9K+am7oUWmUu
TVmFJZBHZCCDM4mMnJX8K30C9E7HWIC8O+8+PQdCjJNHe7OUT/bvO9qrd9Wa5ldBYEAmg/HsBzJw
yQDitx5nf7MnK3Vc0Gko3yTQNpMANj3SaF42RRsnVFMAs8PCjuI7Rc4SFDhJumD8wS+6YAsWriIS
OmEMUnfyKUUH9GJF2kEIKMGH9bnyvkhyVt/roJW8CNUtCi/S5WiI7eVikCZfauMg+CHvERiJQg7/
i2Ru0dGqaE4irYX3ey/hUM8oYtffpVWjbFlU3fvHeMO5RofJoahaYb0VMuNO6OPXCAs9/ItcdHX5
aMls3DAdU48VHoWedYgdmKMQzuPxJeLXfpKwP1QPcnUMNcrEMZ0qIWolTHy//81dOooHs+7anpTS
oX9q/h8ZzE+weq8CUnmjPVM7xFXal0WzrqUqH1Pd/4GmhpajSiKjKpO0iS9szML/0GJVqz/nkK2F
O/a7Rs6u003ENofv33a1vdXzwzGrrwURULonMu7EteVrye2RmSYbPy/e53lmAIMCiJg5Npc1r/qm
Zl9sdKjmHhGi8s0+kjRdtZ+0aEWaCQLS5WzhZzigiRJrwLGLNZkcVPsMYrWkByqQ0VxFB8xiYfyE
iHBhnlScmyBzQlP4CgGdv8u6xH3GCTPv4eCjEvhjDfts9jIGSl+EUKax6XZ0cpuz5o8Bmkulpl9u
InyV15s6V47vkk3ZB+wSjwDPOD+RDcldjQDGjHLPjC3JZaTg4998PfNQ/wN//PN4ESEQ9sK1+TUm
fJR5DmPIqbZv3LVK4Tr9EkjkQpCdgy18ER9oad6vTgaYqTaeiMsl4Q7q+QmjrIZNKELbzd4gvf+8
ZXKsazYlYMYSoY/M7qwAO36/mBDI0cIIJ6EcJvhajSv2+iwyFmGhN0XFFPNgovxFSVfKsvfDYVIZ
tOl0dGUxG5vucl32fhdwEI7xKtPHSZZTW+PgLDMYszTjxEzPWqcek8pIyOQ4buZvsvgIdfzbNu8V
Udn9GAws+ZnbtJW/pm/pF+u4qGfsQO7iwJPNANj0NAULYpVaOdxKIsUHubWvRHVI0MmER58DGm5v
xFZQZZCnWaMyeg51evHaNsE68C0yz+F4J2xmcJoKiJW3z17pgW/VX1p+RJ3RVBFamuF7xTrXQr5R
r52L+RFz8mcd1PlpYY8vOhsAhG1dxhafpgvT3D4oGkWHmaGKLIh3M/TKp7vIcCMAWgyinRAynPui
IcBcvDmIdnIDq9y+ldM6Rm93jyWeGBt70tx1GDkLe+P3LdpNrKLthjqtQFyOC/HgnM7ZyRpiXUWS
fLibHQaGoTVrXsRDrzbv9dxiVqbefccr6Zf9qOMswFzjpE5OUMqK1MYtNzahXU5mQ1FQF3ekAdIa
hvSoaV/DD/DqfmfSfaDiwFILurKXDLwKAzSNxEu6VFb2kxelWKs715NJq+hAmzZS6V0/7JZtFzl0
24b/P0XOA+2ENBDqTfXmTRfJPBHIg3RFvRn92R0e9or0+OI3IIfaOszt7PqOrua+8AGPTkkWbvyX
UkoRdtzsZm/acq2FqyAn08QqHNhTudBBnKN/bFrgcggT7lAGEyqKvb+t2peEOcXTj1uWX+xB75Gd
dxwO/m/fJZqbTtWyiVpbosa/s22zl6J5bIaIK1+kfVPUPZhw6A8nh8N2CwhfTkokmtKS3hNocZmd
ew/mW9YXaxg3zC3su+YDssOW9UY6/YlhZvH6P15qE3/0kfrhho21YkCfPwAF9YMZtSJ8vrrlrcC4
zgjqDxHexOuNYAg0+Cv9lqkRSD4GOVeqccKf0BDxLjaer2UAFmLcSn/ekn/oW27TGoTM/E+1DXJ/
iv1Xs4fOAmxelPqPkwAPSSauPkgXxynd/l008FbjBkQyRgO7OF9/L3NzNjmQMEQCF7Nvaz4aDg0u
Hb65g5jmt8pvaw1CkBu6qiiaG2HdX/ci8suGvZm4NJrO8IbhznYqeMmcpTneD06tS8mWpXDQIJvK
c9qGUOfxBcaosbc5y7uMB7tkS0aJC3WgG3RBI4CT3b4qds3Dw+WgfeeTw8ceYEuRumR50loL2K7J
uIYxNq1tOBgnXBTw/VbFtYsLZzDc4ru61etDriyV0mR9obOgpeaQz+oru1yF9vSBE6ACloJnbFk/
cY4knr7qUNzDCvL8pjSY5eLAedzseRqaEEcl/bz0tbYx3lRnFo8lnRO5UI/HXsB43owqOo0a88Jr
KdvEAV3oTn/GZrqDH2nrxvitWlsXY7efTANnaNmMZzDED96IUxJG/HNsl8TzBmVN0WChFdKwE4Pu
JRHGhW3jtNna+5GixX/Y+LDq1oTltBcLMK8/rogPpVPcXmSQ2RTtuDrlAGLfOqTlSas1yF8dazEy
wjYRoKwdYwvuI47hj8EqwS+XPncOg49f2SH9ymbjzVnTfpxlka6eqh7KLulsXatUnR4AVrjilZII
Wfz0jA9ETokU/+F6jL5a2sXNL/FsJ2Onf10lMXAgA/Lg07+SEJOQDHFC2S6G6ERob+tsUqKzWl2i
kPP2s1MsZX2if5abiv1S6Ah0DTuJF9KWU4Zo6tMueg2JIz5UOtBHLo983+lq2qwPCSEz6klW9aEB
Fc8ka6KNr8igPvw4vnFvyDeIB3yHSi/tROy++a7Ybq25rFaL0JoZ/yq3eGVCWVlzzDqX6KfG3EKV
zs4mcz7tXR4hIa/1NCs1aihsbqecXBMlRlH31Q14cVu4cJYIYisQJwoaSdxYo9CwQEwmsX+GQQAB
FrGiVhbio3JECykPfDL/Udm316Ga11pD4BeIP8gjeQEO1qYJ6RI4OMlDJ5SKtMVb748JKRO3zzps
GLIrF1Z+Vpw1cgQUW8DAgxTuwnmTMJIQyANXV2HErIxgMNSoeBYr/62lfUl3s51GnHvnhY8f19eb
0sYy9/pbkp6qPD+9PiHF7FN6+2OrurHfM1bse4X56K2ynson5FtdGwXCpN5ENhjThE5CsIegYR51
zRfZvNiOap09lv1l7pZfnIIoon5VGyYwQdmG/BbO5Lih5dMktszsWNHL/kneKY28GW7b/zOzXV1R
eRzXTZUYSX0u/uwkhDSFn56mdqlbRSCf5+8IA3bXu1FNcTAFNLZWhpjONUPgZCPr0gxYuhAyIVYt
XXiXIivbOiO5WJQ0VqexNhbVVaDxLbsYixLlLzzGGZJsF7LSvGn+ZxBR4Z2YQ3FkLu142VBGZMCI
vqoygtNBqVJ9HkIv/+LEpieUn7giOIG0+XCi/mPxGob3z04UAYkK3DOzEANyAI+4FSRGTHIbgXf7
FE+6/ljwkTXn6Gir2x2PVX9VEpraBXGdVW5zd8+z9IYiOcc+vy/2LwzcPyNuaZm6Y21gplShKs2p
tSCW9VYXPrWsfXGCyZhjkZVBBfrSzlmUMf6k7D3HOgjFi/Gh/VwoGNcK/MEGo/k3YJIA0FiMLl2R
YHPcV1Yiy3f2joiw2UAi6hoxsKWUl8ffl2+fDxSgpXCVLfJ5uw3kQ3vMlRf2o697T3yYKPB6jT6d
bRCR6jcN/fpZ1LIFRb+efp9bQ3CLboa8j8+XOgkl7Bxx73x8nI0/BawT4DjQ/TdXPXDioFeOUQRS
XuX7ACaOQl8WNXisCLHMeLEzbdEnVfRSbSMLGlEPsFQcv/fc+r+TI9oNm248LRykf9EhLK17YcCn
VK00F2W+dCkYBWkVYaO4g6E6Io0QNxbTd4Y5XPzQQWbDa0Z/4JHZ9Jc23u+QmaCs0XEiEMU8pJmK
DIMGcMk3ffnxWhWz+Om99BXQCDmkN9IKOB2z/zXkhmkJBQtiJ7i0lwagunGzRko/VTNmSLMs4h7o
57Ynk6qiSbmf7/NeIXdjqXl1Nx5dQJpJFqSsFvyB29IA06at8sIz7SA8KSHaRzSLFXELX+raGb6x
ydmIk3PVj1xiKfBTPdrIeZPuFrcsM2HVFGRaObmnLFgRsPzsArX7nbVcy2efYJu5TwXvXKKPNG+T
8Z4MJRQmMqH+Dp2ed4kmgbDqJX5SrvmS/Y1fQiPobkOxctfigIRy/z0RYU1xjfDvC6Ly+vM+gHVT
Ydm+R5CQiNuPrc8xnroPLhVbObi7LGE9uf/wjTM1J9PZOQ1W288Q4NOLDxa2A182pPT5hJ4gjtJ+
ALDLTiWk0IY37tpVw2I0ZlUIU2tmZ8FKd5Yp/Si7PVgqg9cHmJbThpCeTMenYGfz7DKSs/VWa+Qj
XV2xzJW2fKcrgVi9Ag4h5DDd1kTfFZXpNuQhb/i3A9fyRxMU24g9SlK/d5Un5zRJPmaPT2+tFQDv
sleDTu6l9okWukUxHZwb3Rhj/LiqcqBDiI1dIj7hFicswr02mYeopOBzWNXapLnQM0U8hy7AmjHr
rskDf7A19PjqJbGdVDL0G/Hi/4PY3FzAFsVjqecvilQd3HUu+hhHK4x/V5AIOcKOiUr98CnzSn73
zDsaCU2Zb+/yO0aRJR+6wIAaqH/weBSTdV23iuwQ/u509y1WPzk8xT7HWATQpO6YwJdYcdwkBBDh
aHfQA+qePquK2c0zEsKJVkkFU7AqA88jl7RWX0pklLpnLWr6MpLb5+xed+kMSDj446noPWxTHt7U
k8+CbXy6pHDS6RRyQgDAy7k4naOUKfpikTHyCfPM7ZM0cFFMqrYFwzk5tAbcbyPQQDtl8SPLkUYo
nm2ras8WhFd0VHWaOFlifqXhnyP59yw/SfqKUUlpM33/Hus9NhC2zrl8A3m/a/GTlW/4y0WP6Rh5
YjQHBtMIQaN0nOReXnclGKQxJVRebt1p27/2GiUImMuHa8I9MJ1gLgwqvQOnPX6TJpv6wvpeGhme
K7vctWmFIEknCv0XkLt+DHrGXVeIFImJ5kc3uCdyKJlnX9FSVA+ba4tYP5njbqMs11XzAOVnwJSw
crjwvGNnynDtemrRMGNT1DqTA9Nkbv2lWM5PKR1Nui/yPepc2bhCgVkYR4bG3EHwqKOK3iu4qETi
CX2t5XgBIZW5XOcXRoV42x+4w9NmFp2V0WmNzyBV2cBj1GF3u1/uztCpEqy49WdBHzP0By//pp0h
Ku+UByHbSAU8z4XziRtf3OHEROBIzNSxNBe8jdibkxTuZedykZuQOh8Dmd6ek7kVscAVKcBHKN2X
QVOuRF8GWcU48hFrS/2lC/4bK/P704QS92cc7wCpowOqLmvcEouWCd4yTsvaE6zQwWMRTR9JOIlm
2B2iObTg1Y+SeLeQCO69R+1BrhC0wZDqjylr1z3sivzsOJvVR337pClxI9FYZhwOFXHz3jo91Snj
ybCO46SZRpgkpCmVzRpbNhui3H5MvKV24uRxzWSABc2kY4gQ8kq/WnDcNRy6X51xnNWsj4dBMFOs
WHaec9Mvl4xH4Q1dpZJONUAhGeDhMGFVFPH4tSlkICrsWAz/OPiJoJ11xPm5gMfFTq+nELJVQ0i5
jiKiI3hWxn0EX8Ki2l0eCSf44SZSa/bPc2rAuFfF5EqX2wztGSxmafyc9tf0lUVs+Mgb3lQlD627
a2JprhxQR7zSHEudHkvyPcowQjRcDaJZRUA72KKfpy8E+AKlvxJcYa6zLdtC9y165R20kG3V/Wd/
9zxb3YZtcvkb4eg6FpY8UFmjojoimwIR8En6rU9g4ox3x5K1m7s6b+9cGP5Ty1/+1Q87ybOnx8v5
t6lZpDd4sRcSvtQfa9pvxBNWL8+W9NvPSHVxCacHr8VjAjsrie3cUF46JjhnVfuMKvOsfj8M/YLK
TiySZcbLhevJrV7MYYtHs6Gact+AvrBlozoNB0w/swbC6F9lKDhBIGUECYzTBP+qTHf9OgPi0wmH
QTkF2hXwtL9lz4IBr1HLW3lFpaMJYgg5ERp/yt7dXmPUmZWeMKLHXPmYoHNb/FGrZZ0PH8BxZoBX
KFOsFbajEfEZMLpAafbXtYC8cIAuPVuyimrzs7P1ixgy4NdOv8qB+HxUiGwWfQTUmTcqhJAT/fXZ
cp+uYkF2jr91eO2Nlm0J8hu0yBcDt1rhx708wfqxcPOpsCd9VTlOKJRoQBCHrGX2djBxBQ9bUct/
QoJ3c6in9Ct7RqYj5sr7sgpfXQSiuydOjZnCHh2bsanY7rFaDP9UK7CryThxCUWr+8MiOIK49vhw
PxWo+qbaRMLUUZlZ0nX3kjuKdHvWtZ6FlHGX1uLKbVLyKgRVdAsXeUcIclPZpAnv6NcD1Yz42qoE
byiqt0H0Sk2ZhNnLORRr1xzkkoxWq+CtXsf0GrON4XZng6y+ay+tL/H5zYfFKUqdcDqsrgXqlM6g
umy+0ZVK/swssu4n3JjlbznKDIZudXlyaaCyjN0GMVWyGChNKmfZfk70W5iybPQpyD62qrPenroZ
yhz797exif9VUiAiBMzFht6dToWr/t6IM8O9p2BxJonaAwDnVwIFXKpp7/2lo+XEMLTQz5E69KBG
/E257+IwPJ+0jTuVxXMV1hgJDFGirIHsc8/k9vSSzWYzEfwJGj+iGT/7QqkGSSyCEziA34ZJ27Pn
q8v8sfJKDK6MmY95qjQUCn3voi0MlnMIdgxXJo0rIsfTg6YmNk+KADAMS/nizmP9Rt068gWAIiQ6
T6BkhoaSUqmgJxaasUXA5nXu3S6QDMXwMAVV9Gsk6JjwOMuE4xO/M4n3Lc8z0fQTnYfQ6p2S+OjG
kTJTaN34CZou/f156FhpWZ5nSkK8NOPoR9ILO97F8Kmcq212i7nyiSfsuo6XFxj3PTgTL2F5QLjX
6fe80ZsdRrAESjNsIVJB6D6zoBqtJcYX/X79Kpczgyfdu7XAL/bkjdUBkQEVhJB+638LtWQY6RmE
thiDjEp4rPDRFUQHQxAjxoRRsjBVamVouIf94tWOeNoGbWQ8KZnqRS2/H9BYySZooPUJ7XdlN26o
1oV8wbBJgijPUxPvxJi74L5uqTT/QL8txwEDbwTk0+1IkeNRArnH/krEhRAOUgSu27X8IOnERqBl
x8KUUEUNzdvBR++Hv+UlTiGQ2Y6s2q/DCxYFozrMU3FtXdZGkFtHu2pfbdH1sc9s03GoIpKy4i6l
eLijNrtO2/smJGAXfqJsToMl06gM1c1hKqKGxJESHhSvslE3ixv734UE/qB6LmVDkvZWz+TOs841
wzA9QokAbkOLQSJaK1t9rqosxjxt16L2URdK82Wlmqu7mlxSADRsaLUUsl3PqKmbqtr68GLGY85Z
iIvGsuVIr0f0jcB2QncbBzSW1W46gFJicXuEsoq8dPSSRRzPXaUPUI7B3yeLCNgByIquvC0YpYuE
QUtId2+gYP3z7ljWRJj+fTBfkd+pidqMTvGQfRr2IswpUSOViiwERT/THrAmdHKabMngG1t08v8m
0vs2W0/6F/p6qPOruRMXA9nqaU52Ks/T38tLwPvq5Vvl2V/a59pDuMruTmBqnSFVWpvn76PCjcK6
+QGT7fDKl8X2lFJ31yRUbjX+ugvSfdKRqjZFerbRpyCzgXOf/o6sGQ8D3gCtY2iJskYwvvhPpcmg
EjVN+IeNMYM7n6v5vbZQ6kIHUoTmKGlsyNc46K7S/tOHCOV7nXphJyF1FpFZZrFoGkscQpP1hbpd
uYS9HilSPAQkNV76K/6x7HDp3zJDnQfVLALZMwTF/oluCSCnjvqNWGO3uX6OebYyBFNgZlIfWksy
a/6+ZEj+KF/76a19o0BMloyCBA/T81Ciztugn2/W5jyXB1EmqDTxyI1XtbkwJKILUhEiQtYPe02b
ygZDHQNwBU3ZJmjPw0H76B0/Pghn3DwZrQHtg6LbnbpeC7UCWCWj3xWVffkhKa4Hhn8UklfRWN82
DXcprs79DUiDO/s5MZBkbTfhgHnAdTSaadBUOLZ69zkJ70zkNCK7HcxxrDWjD+EADN3GhKFkVNj+
hM3DTP+ePZ3zNQG5EN/kpgHluSHrf1NHpw0Fi8x5jacv5AyX4V7HhtSjvIo7Y80Wf9d9KcfrrDJd
+bzZYWF5jfUjEkDZ9uv/DmS/pVmqdC1sB5VEeQIpoqJA7GudvTO3uo6//zZOasmrzZLQBBR13WI5
pH+731EPvLl7HBLnxDBwnvL6FRrG9f3K5SUTC6L7dtSbidli2VJAsNKP0e+6APHRcMkker0+ZMet
qFcIlHSGcKo3aMd8YW01leW209whn/tjF6IEz1aJxfEsL4H4bec6QbH6Qe5RhecN9L95lC5I567i
lofub7Gaoztmqy4NDhU5Hd1Wf4uGX0sReXjC7lMqYp+QCP4X9qf3ACTV1LVCmnfqq7tA9kHeFPmb
/T6FqfVAblQkLB1E9tOAcz1TCD86r/81EhtJzPnI7oLtcMrDqb6dOTmJLnxB2+UDgKvx5x/83a8s
h1BjU/uLrU0GxNZfMQxVN3XhpgTsJnzEjXESpyqqjjLSsCWV87n6drf9EC9vH6tYeGHmgOJWiDfS
AuibxRFq48viUGqcPrIn71wXL6qOACjKKxZVvJIU/USQBKeiG5cwDR/sluXBOr9NxB3KpAxkv6V6
ZyDKsUgLwRqmr176ne557KNP+pfasZAZcTsKc26Lfq3FHK+QeGoUXaGc6JyXMPDNdroG2TnRdoL1
Dr3Oh7hK7Y8zeZdpVskplKto9rFLp6+yw7/uqVYkd/hC0Zmn2MVFrC5PUxCWHjsJW4iMOx6wW2MC
9Tg55xC/rxjUzyPelsdLg+P3G7FSbb50DOgWg36O1lXU5yxddyau13PsTZTd/MSsNWFyCPSSgTyi
TlV8S12GXsrpt02OI9r/xHquSKFYn8d/keovc4fRZ73pMgQQweY61eCZFVBi0QmJHHpifhp9E7E4
7BS9sQYQLTa3x54RUJxKcOK5boxkXrDpZIU5tR0heVkC95xaQLJ7TxrUi5eyPNeBytG7jpwbWq8g
kY1Qjh09NF8Vf0Poui1xr9ZhzKbMy4GwReFIt13v3+xhh91k9CGchgOV8WpjNo6pk8nNxRJ6BGc2
mp/QVHRg4Lksvu8C42b4k+ymhyRCjVmD3LG20kfi2GiV397UM4Q7jGnvpgLXNWbfl00WdozOks+k
I35xxUgv1D+ejQ7maz2DXE6MUAzg9AfOsjS3EwJ1goKF1Wc/z34N7hW4rN6jxIDD8k3ExSo6FJMD
jRPNLI/KU7u9r297lUCQ0e4ESJ8oMRpuJbHZO7BThVuipAfIIP9pGgUXzyFoSuMzYzbvnilzJC2h
xaLh3jf6KC9WodiUb+a2YR3wjyiCVeeB9sUUN8XVBY3VIsrqdUj/yFzldbngoe7gpns2VCrkTUHi
tK3DhGjK8wuMWRO+EsMpkNFXH1qMzcYw3aaToCjJ7a/7br0Dz0i2kzaFD71o+tX4AiGsUn6UEE+m
YmBs0mF+kawFudMsgMXeHfZflRmpehEO/j+77+dInvxjL/HF9py5Zkm3C/2+dWyIj6wy+aHF/oFh
/Z7UgJjhkyZyE8l4MDd7t18vXrmCvzXzCoQHq4kxfVAHUGFvNQufGgOFE9h6ODzklEu6MR9lhPze
ZU9PXiK0oejO7LCgzHedWaCXLMV2ACQ7r8Wk5FZEY3xB/SmygxrWoLl4gh1Rw77LENtora6kgG66
Y6EmUvgYXtHAaXeAkKNqJepXvVqiwYGB+MKeCo4Wo3sp+PZeGvSBJHyWi27fvMI7OFelaXyj88V8
k8N9SN1aRyVztKTTUwBnIJE2tyU+vIl4Z7P3NQdtCBEYagWid8P+xgm1atvHCQy13kBVi24Ui2S5
L2dn+8ts0zHbP/KQiZxsTBoJORgqz4jB2FV63jmpgfABqzTLjAIr+lovYQM24rvVNB+5/lzauNYv
+4bMCtlhuD3RlXWM0WgIzF1sjENpFVQFBTs+F+OzGPz1DZqvra95paDQb33CLPp80JAPnB0c7cf5
FnAGGBFhEX99N7dKBwyuAuAyrBWkj2YwRoF8MhLSzqej2HIX9v45MEoQmlHB3iSFbRD1Q5JX5qJB
MWey7VyOKE2EPvjaQpbf2P3SED/rt7h8DmoUMHKFdMb8wVbnzPIptNzyFp3jPXz2NVRwr+ro3tAC
6pduWcIueYC7djXwvWtKKlVWxhG8x5pKNEkS2FH1jXFs46Yi929bQjiL6FL+obriPV0LAljGHJKN
t+H+ZhtJZpk+AurSf5svoeT0fK23YF76sm61hb43CQkvywoc15w7EfHj2tsFuE4kkn1JobfVh2A3
26qdNXfyjo/AFbfUktOjc2FjDqu4XbvameX+y310D5FouFdECnO7sFZ7tVP5u3DzrMW8OexL0Bol
Vez6pcdokBtKQStkL8KtIwzoa2lZqKEXxv3CF+PA0oVAgAhPcp6xXTpPLRnpEWuIFbG7kO4IGgJB
WAqX263dWbNdcpbQVsF3CuunQvNhXgJ5XrhfzZ7xXL28wjP+lp8/lEWfGm+GZYk9yf/lAyHutFq+
ysL89SrYw1JwhsXen5+44HaG6ELfBLyThnYdWoOlPEmLY2sCAySKj/DpbYiANVxre5trk5jndmyT
XqF4rm2DDvLE5w4HgNgRDIvPJxUFtfXjs8t/tmUBQqmbWb8kUSVbWWuLsnFiI668n/V9NDOa9ATN
hjBrKJw844e2Vgp6FvXHBqcaxVLfks/s0Y/BGEpk6pSt6nhfpU6XfYkkPNYASykc12qqLtzs9Fm1
u1ENa721f616ZH34OiAQtGo2+TjwwLutl+1Zay5J9cqhWUiIBOEiGW+4R9FEox1IFdjZMnyRHxeL
CYTsU+GRwzYW8ueOmeK9vsL0DDls+fw+f+vinjduAjivOczBT7LIOGZX1QdyDROCG6eJa4QZj9KP
tqsFYaco6yNWqtOkNgiM+xiBewM1Pf07hieHqX2w4pfzruumN4zR20oew94wfzLWs7vyoLapTvZ3
1sPQEnialxXbmthYtR130St0lQC9ImAcOg+XZMjfDY1mFMO8yUgY3lYj6xXilusfJUQSLH07RcRH
zevc3UJTWfBvJ9Gl++0QY8DfULOs38QNcwB9/NhzbrSKayP3bo5vsK56MVOV+Qh/Ep9rCRsK6PGC
kKlt7B+FONI2/GXDMScZuFRpkQqO7Z4POaEXoaLoHqx//++xVKmMFMKrE9mgADuxqgrDJZhx9T+/
4mFFRsIdoUKMde4V72eoUvJDmjsaBNfvfHGYpGoacmWQzp6s9+lvhArQSry8eGy2uvBU3bboqcyw
Sy7cZGKSiiyxNWZffQVGgQlliyzhU5CMgErR7clV6uxBfOTQKUWvspcYCUrJzMsHuWXAflmxckDx
N5nPufzdNTbu5S7wAAsV2MmkwyW0XXvMmxhku5mMH5KQG0hEq0GZWHr4bQw9w2V0ItsUCLuhwzC9
8PcrOcT9GmEzLY6Jy+/QNFBHSQF7YJK6MDqBetYQlUNqnE8xChbWUvsYv6mW9SCfj34XOwd8Kj/r
Zp+4gRq/ASstkNjnqepNEnTuYA3vTPwVQqYAYu/kE80i+CvtBbq8AR2E2AQyF0IEJOG0ahRbvKea
1jIQO9Pblzvz5KO0dPT8caVOpXqOeolMUnRfZi78GT4WYFtB7aLgZEs2FUFaLpT0s95xS+g+364m
WOeLGdCdIb8pjFExPN2jP/3VtpD1mni/tVuxqlA3oFF1ndvH7qymBPzlB/tebDACySzzIrNj8WRh
DimQRzfCWdrpCoiRVghWDO5+yohN3Dh4K9zaLXMZMkkrMFvXphK2tYhmyN1wdLiGXId2BWGMaKfo
rwiVotA4vp/nA1pe+jv/BF6pyPeQ9R1/98qOHQh/kU9yQy5IyNz5zxQ9gwSFXBl6Drm+SghVAuBD
aBNUaAMgn9i8IOAHVACYge2Yiwo0iaku+H+yyuFFmlzP2jzbL9V96lF8Z95l4gbIaIkxaYv6ayFF
JECTGN0xOGXDnnLP4NfTLtU4ZhckZeA6ZIJfkwl0Xa7WOzDnqAokiOsaMwtvYw4dBS/jvTEjH0cp
MKT8R2Of/1nkZNZ+PA/WemNsmBFaXk++NC48YcWNZK+ciQioraiLc/8m2uR99G0ppnwvp6tJolaq
msokPhNkgqpuKJO/IGqwir4nARP9So4ydW7o7Etc/0WqwmnTWE7qcsfoSwFb2OQNHXdt8tCQzj2L
akqd6phZezhfA8CruqMGffNV7sklV5a5WdBtVnnKpX07xTN8ilXlzdF2wTlJqV0tZPn5zXAEKSIZ
WUyTvRECOdKZGlMRhE6osdjxLj9cOk6LLKLk4HIGwICKossxKLZmFCayCXaM5iKYAk/DqscLugaR
GJp65iHdpG0he24IDRGyGxr9YnsUDhhb1/1pET2GFyD5FgGNkKrgAQiV6gjhb3ZBCHcUplilc5/+
QlUOSRqwOVlvzqcJWaQ8oFf5ebg/iiTwaCI2FlsBGO3JYIgm0O9Slrv/Tcl5wJ8d0bXommfM984q
NVULARyjBKFDcZaFyzC63tZWSiZjtF0IXTX/9EKh4L6xUSl1uBN655tUz78QCu5KSfXn+YjT4+Rz
pO7dv035lLr/i5XW+TL3NEReYK+/FznX51hr4fLp4knmFI2zLAjp0Ttu3XMGaJRpnyy/lTLcr7GW
GN+DELLxgeEZbnar4Mws7bPBBjLtmBv84ad7yFSoe9GMPMtcZvoxlSVRuT07qkZpi5oSVmKHmKPA
veGB4eUJ6H77FYTJT4jxyTgrFpHatNTALZ8lxaLltSgKdMjaS0Pf/K85MgRpAAhRYbgTYgCucvHp
4OQJO0L50VkrLdH1Mlr6VYPtLHuA8qAobfx6iZQ/a4Lkt5xgzABEqODAkvKSmNJDeYk/Y2/eoAkm
USNr/ROJGqejrH0iHMm6k2IhzOkIsgt4wY8afv0+7MAaldbR5HVy3ipTKNkG+Kt/3BEtIMbXXDLS
najOfCKpJdflvWxFHUNhmRAJxr0gcFWE/r/dj/CLvJBPKNP/Hgp+lL9vqO8esM2GmcQa79Rh2BtT
olzLPu6B8h5MzrXcLEQx4a7ritGVRVj4IiWnALBVSxhbMCo3e/+cL1HugOfE9FR/GB9WYZJtlEav
drgIqWkq8v8R7t4qgzAtx327EFgVh2OYtvbFFaan5YFvqyiOgJEp211miBeoZqzPWjx6g2kWr1Ss
7sMariYQtk4d/+c6dzuxFgzygh+YAQVt8sXMGxl2QKOT69ypvhbvrTqByD24flwinxsR192CYUDv
5KvNESvkRtZ3tjL4vxFTGEQYpAAp1P/9v3ieWUNdXTL0YvV/wU53QaaUrDPVaYXoP3J6wo2U1r2N
2QviQ3MiEgz1G8fErNpT6Zyoy6KC1chVFrnc7c1jmngNRU442da5htBM3pegKkCknD3CXMODiWsQ
uEbXFzJkXIP5s553wbtKkLEekBQXENB8vF7oEUWFKpjRbI3SVb4LBGA3nuCDf1JSaiEZLfRVZRi/
QeDbzed4BU5++3OjUraSDtJIrCiGl7UPlPo4TqqMxh+l033cge8ljEBkY4AEy6p+sCw9IOo2GLty
+pVNL9CaG/3A3jGLndAOpEdDSCSoCneC27X5PjKDm7ErCmWEAyQdE9GZNonOYNy1kfjD6R5RJcD2
cJO3hoZ5nz4Ds+8MF4y+cnDe7IqZKM01VAZDKDl8Ee7ijkXixDfYrt12yWmZle2sFmY9kziplx4I
9W5ggmKKCn33w1CVtDSzZYxZ1Q6dGQSGUN/MWdUHtIe7iJmGdeZAktDExE6ZVnPXPWprRXYfQdLc
0R329qooqotJYDp8/+q5G/JL8bVSQuvC8XBTqcllS2zHvbjgsuJKuZ8VsokaM5ynaF0bsAMpnb2c
PcaOBFeDy4jI37QByx0w4UdE5vFSaVRgYAV5sdHdwt8OiTodZLczL4cTmxa4YI84F3r4z5042YIo
VZ4tx/2QlvI1t4gUDGM5Vei8AeRDNNPm6rhuY5eKsjz4Q7OpOv0LvxIUtb6SiN2GpfVjLda34nVk
uV1luP7346NHkdLwLesPBpJrYXCJfH3vQj/b/9W5kkEDiUgnhsMIBrBOfFPJ8ag3v64mKhyEwrVa
Ixv8pFQMn+CCKDVD5OYSQtChfailosLfytMue6vDiNepNQKFwfVKE/NRMx7DTx+WPp4pNwVTzwYz
bfZ+eo8C6mMimH7AE8Ux3rkh8YjXGtfSxZwX/Yd2y30RqEkNQkcCihjMExOBWKAJ79vIOMmeYfOT
rBD0GM/xlyZYdkp2X3KitAyxXd6f4XeShGrdmYQd7FHx0t2i1gPK/HzR7sd1JEEoTPakxDcz/9US
sYgLFLY2+5UCHkxgjaWqildAJ29l6ipOU+jBinSpiM/Em4GljM8ohn7Fnb6DFaJewpxh4UVVMqvr
9frtn33nFe+EzavoDwMmk5dxM4PmD/127HQ2qrUkGnNMSrs/DJqRMECcGqUxFcA/k6cHOZCTrboE
3bJwJlW1Vy9JsRtMqJO6e82ibAOILIE6CVTifXL33cueqmE0cHduNa8R5I1XwPM186ohaIv2QoMA
25qw1gRv4nNhfF0BeKWmAuIAAd0NmcvQ5emq2x4xN7V5IcQ7WUmSY2pMbRJyamZaSXaFNkoJEMq5
1/c692fWVDGC5QnFdPfCVwEZ9DxN3TaeGP9mQVPedsYDsxc6W8IkMGGChjvvpZnYGgDIlV1a8iof
NjpwOR8HCltqUsB3p/TtUizUxXM8GRhhAE1Aw0qpOgPwAOlW9Aubbaem4iw6yiD0fhbkNtXl1AwT
zn9XI4DDkDodXrE5fi2/BDLuDJkE5tzWrm9FbMeMzDBYx1GlbzdOwIQEPto1hspjSqDjwRlWlxLJ
EENDZPqM+e1kbCD1Qq1TbXlXukV/o07i5l7TXbhl/4I3Dx6Ptv79zRgUTlgWzr9a6pB6qVzy5JhZ
hWZCJ2AqziURA8m3snfJ1VGwNUewh+cCuzptebsSR5GDR4d3ru074d0EODn+0EB1IVUlgGRtaNaB
a7SqstI1Qm6nqCGyyUhGH7Bj0pLEhNBwzZ1rertMtA1vUF9ulxijKEm8xCz+gRQdrdF9psJntMvv
IhvAossw9JUMSxmMUcfR1r9NKOQxgDR1tgaC476ZsXWvDy1AYBhTVVWJU+dSzAya3bFvQDK1NFm/
ZNqbmBjjJPg3aa82oKso3LTII32cKuq4MpIYp3iaybxE9EDitHn6D4+3ChB3LJfFqEysrnRrvQDx
GPOL1tf4xtFO1Enp9Ak/5HPPHBgH88UyjEQ31n8AuToe9A3U0kIC3Jt/beRElDPbvPG0rFrYUxfZ
/1WOWimM/8YcdP+XEslB7S7SF7o+J4xuPWjeB2eCBQZch9qMt1ia5Dy0l9nIR5g0ki0+IlXijyRC
/4iUouT2Lpe2k+t/2ymnbKLcAJyumjlZ++CU4F/Sp1LDXX+cN8OObXGlew/af84O3+XZsNotTeMd
BL63Shzk0awXDvzCpj08tiZpBfJIEP+V6lrLtBdfZ+9cd/UGyHz9zOtUgbJq4PMvOU2RRUYIpDCn
D2efENV/xcApq5WOo9rgZUeE4ERyEoHQtZmecJA0bwIrrmoMHIDp7M2LcfT4wV0co6yP5tn4hMrj
9jd26ZBZMcgMcMiR+8rzPCQOfWNE7aZM8t7kM+z/lkCPcOP9BwEGlPOf2ExaY9Qws2X3B46DVFIf
ZFkAg4dR0ViTUXkjSl50skHuiwiGJEGp0Ms0h4peF4fBwncF6uuY9K2kb0v5jWyUxALxIDA7otE5
yo//Q/NzIUEKB9K1ppXrTD+JMzzZH5eCVN+rvfDlTKisvy8qI8GX9xFI42aMKmCfCOxlHe38jTv3
3i5uOg5dPsF55xzJNDVLQuf6Be8GfpVzjmPMJSSBAFZTnZDX9yCJB9JMP4AETdx0PdDJrjaw38lX
KuwME6yjdIvqVeJSMkdZcjzU0xhHPI+t2U6a2EjgaWoBKSX/kma/YFlm5MnZfqwENSR3wWmVmK6H
ANgM5bjmdZdD+QIPDy8CbClH4TCLVUn+/LNsN1GnQCxJJgMNkVSWb74py0x9c6BFNAGtg6dZlFxz
jJq7l19gFyY90vnY+M+eLWSVTG9xk0K7y0lz06nQaiDL29OrSwChRK0fL2/JG/it3dXmKVHRV52A
D+jUaBP1IwVaGzscpxTLiXWruD8BpPb2YpbzWcux6urX6K7Tq/KPL7c3/U42wkFF/Knen3QrOFlt
D1ae9kW8j24Rs/M/pXl2qRQFtbBDCOXQ0MsC3Cuh9qc9G+srCdNVgbiOfZYLYSv8tIKzY8nSnn5q
Tzc6wO43bo9SFBeCJTxOue3zEambpU927y6hLgvWyZ5MbvG9vGD4MVAaX3G19KlfG5bUT+TDPm3N
9FJb2XpDP9ZiFMW/J5JBT4HioF9DIpFTbPf1FCYlxrIrqEFGmICMF6Byc9o5vrnSYFUvRJPEHFuI
6HIU3rv0gavH2wztlpsPBb7Mtq2wrdHSaisDeOyBkPvqLry/Ztm65ggcvstdK4QCGj8K0JyqrbMy
V16Rxmh4IJTe3zWgyzhNKA0JdXrlvnWPGEVqDi89x2NVVkVlr16jjQOAbHQ2+MjT8RkrpNpsEtLQ
aJpvW2iaG9RlRAtGvhsHNoFgcyW3FIBx+9UuMB1OTAvrgt2+uDLJvUV16MEvKVmIR3KNIOOLBqTM
EURS6B0e0BLLDt5M4ILpSL3VQ1Mjxya24Zrl4g8a8mb7r7nPi+sZZeASEkTLwuXlCHdiqfGncvw1
SgHq4aQQWAYNf+vwgniYsk8rapLMo1DQXrXAaUOF9oxDNvGlGSDeH6fr0o48ggrm7A93/CPga4T2
BMjH8EsoJFfYlbYSa7UCeNSOk9PE3tcVyWVplAtFgHTBaEWFSlY/uS4uLK3ul+qK01T1fJyFWkFu
fqfwX8Bqr8iOfJyMbWaXsyx6BsvUGJcdbZxn+e0D3CbHdGJTbohH3845S4RhG4cQg/LiyueMjTY7
I285ovIW2e9lKS2N3EeYEb3klWvJC/nPMfb6v5OPdr8RfKdKeDKYUv9DAQIbCI79jIiTvXBi4bDs
MQB7Qjjm75FXdRgW7N8mWtQOKn6sbdFYTYI0w8nPQb69FJ300ZXkQoZ/H7xAbenRjQc/57RsWX8X
mhtJQdKC5B5pxOgkbM7dTI/Zwb4I9tpdrjDiymgEExchd4Sl73ZNpdevql0ES+ng7uqJ9COyN8a7
MYnF4aeak+P93iMabwFGfPnUOYxRwfhV9m1Hmx5mFIyOSD89WHOhY34yD3V5LRJMdqIdhNsa3UnT
UrlUZ/qMzWnvl96R6lb4kbWyg/Yy6utyzYBD6iXHSZ8WwFwPmffg6s7Rn6XVNpMoDookc1Ly97sC
hymD6gFIs0bbQxvoJR6BSfAkHnKq5Ez4grgLVb1UhKHY4NZH44Y9B70hmXB9i9a04SKJPph7WxSZ
q5VN/B9YlU7aAjBLM+cYWOn33KD9U8qO5M2iZIswpsHp2Dtf/5QjeVC1y/btwPQCACAEFavdJ7FE
TEmy9wIZP1HHfAzwklTWrlCFDl+e8nVQMj7bHeyDVIBchtUICUlUE+25Pj0t4rv70C4kPVkk7k3p
8rh+xBhY7oTni5Pc7SNHeDi5S8ErUIKw32Arp+DqX4ZPHTxWsBIvAs0t7yigDBeALQHiGgP4PtBm
W9nDKaG0LdJ6UnTv9nFmYOGtUOi4Tbx8mI5ZOz9xl9duze6BZn6UDPSur6A30I1AX/FXV3knIax0
eJE0qxc+fKNAaAVN1aSNGDq3LV5dqKBZANI6Vlism7QLaySTTuwMagrRELatjziIzIy36fJcAhu/
ae559LRrStAhSOb82wcB3NifBnb7tbHZMYwoHs4YDoAVYNzYPkiyvK0RyDcxMmbXcRGIsGJmreJ7
CvQurHbMr2L/IlYsnFUQdj6O5g3oGBFw8JHF0lj2AiAO0Cw5ciU6peTur2IK9C1XuKl7spHahHwU
hOAvRTQN2j8krDRmUoWxYNDxdYEGramW8cTYyi7R4Rm1aOOBC0YE146+jacxXjApHwpNGRnmdwRb
B7xEtcEMaRHgTPQcEN52hC3nfv0LNsqyLrZ20Wmt1WL9+Q7V9MNieeF9hHx4yWfmYDZBzsOaYItE
QFFSekl3w7jWEqH6gaE2vPQFbz1l6fxOvniZKze/TkBxTC9//Jswi2psVV4I0MvBPQIsl2YtpEBt
K/3T+yCHEhBwgNq+p2CKsZwPmYkegVQsHJVIOsp85WFNJz4DdI7O5e2k3XY3VSrDIiUuB330yTgJ
whwtu1AbkZK8Gu6Fdg4HLVBdHRa3eB2L+y4iNyH8MDq1aFgRq2DQU5R5Xy6gsnzBvBpDZM5D3/xV
R98IQQtSyRzYnR2uG8NWmKMBaQScUKAkSVe7HwDwl3VXBgRM9VyDLqft69tiYVaX72rSpn/lBghh
lESZ+f1og3+HI6Zv6WYPIUGTKUUXhrlKl+EZrX/8Ae09s753zBtXI3ibxpD0TEHvA1nCJUNGFUqY
I3NxxiUzyqAQalcVmHFklw2sDwZifmWytyP25XkRNlVArA/TexGTA9OmFPYgS4txmJ0UuVutDmh6
gCGaOREGyxmtjmlvP1BFNrkgZ6u4LNr6ZbY78h2h8VHrgEGp7GKeXt2OThWzf56pKHBUnTzeNdFu
Kz2XoC6iZXh/JZxqfW29puGB4sCSLDZv9c1Idn5u+FXMtqknZsmfWjCyGo6SEHRHfyEhkNFlIegG
lD6TZI0P7UCjWOlNr30fPEvDCoTW/kTDX+ASNjuj2MIXh4pWhOfjmLPYwnST+a0pfAWaDlVJbkE3
Bu6pSo8PGoch54Ce1cHX+0dZfAE0uKJ4FpJhPniwaHi+3NbQAjBrCzY+gOxLRMCjZIXXGsvKMvKo
5biqDKjQNVGUlMxLsV+k4vquuWYIy/789FKEHcG5v5F3KjUD/RHN3kJhUsqRi3eNYPOAegP3b01Y
ODdH1npySfZwz65978ckbrhfYpCj/GtvE3rCNOrh6mE6sY86FUyBk4znAwRHu/Oan7GM0T7GV3xu
BAzBKhSaNatOlgc8Koq27NE8NM/hm9u6UIOcWZkJCU/4daXZPDKXBEqPiWSWBo3udgIo/X+mCpDQ
7/ts2uXkF2Q4NnLbR4u5bfH4EaTx6QSfAssooi3Yj29UhO+I6CR+KTtUTGbsOWJAHaRcji2gk6bF
05Z4NC4eRPZArTBfUQXAMeYwuQM/MGsVinkbGRCsLM4H37c/VpASyWL7RGDkQGhLUJG3j7xqcnsZ
1w9YonyonbS7LploEFW4vxJO3nmI4IYLKRHjwoSqCDRJDoiJveUCyLzWp1IQxSqhUOVAy36hirfX
QE7N8h9vL2gDK1AsKFZAO/pSymxdPJpTTbLX+gY+wEOI82KVGJz7CTmHiNXnOhDIQGicm+SBheup
HaTk7+zCxqCXdGweJuoFcAD0zNK215JP4yJt7uYwMIJb/CMmO5RqCPjyfeV5kOfXbNDdiyxzHCXr
o4c1Dj25iY3ARx9JoRgi0KPVU7HPi0A1wQ5Dlw9bwAfxvTX8EJ6yFOPHlaQ5XS816az054xpmSTA
EP5lBT1sh1iSXXypLADGX4AyRsn+17QRpo4sbfL0rJ+I/RFVEp2wSQT5saImyl526/nd7QXGE4aL
ZGIOC9qpfWBUUAbOwE0Z3E4+i/W5V8px9KhSZNOwF5iY4BvUVPkU3BZYVqKGufYsMJ4bgF5JuEdu
9147XeFtGyLxn8vYDc7euYTsSNcKw+gOYzs1JezpWukXTH+5oqZVVXWKAbwoIRg3RgRnTJ2McWOZ
pSbkpCKAEik/H/snzm4zPQ/xIuWBkEMGqZ9/WYU6yPTOf0jle2ZOKOeJt/O6xZOj2sa1ODmrT9uL
9EwQt5/pUS6ciJaIcMNH24/9y9+wCkKPX2wwJJPmHaJa0v36kgjDGMC9S/JMuZy00e+emIDbeqDV
6b0u8wVMcsZefuindxCDlZES0m1VtQ8+OrIpt/E3BqnReXLf+GMpATXqXAszV2i/qFL5kDWmYIsg
zS9s8sQdSOOP/4P4rhZUfjBzn/1/UzI+iFIAq84wVgL4Qlo5IMPxMIiZvi0aS678xkteD1BftHPR
8JP7LgKCX7wQPTEif8zFUSzwTtzR4hnYj7vuxSQV0utejpknuicQZKrB9D6IIVqzsmZsjbmAmSAB
t/a7jwOMFexyNAhVdx5Q5pLh+J3ySI/H26+SamG8gN0Qz2HsQ2VW4O94UhTJJjLYqNVoXicMPBl8
uYfcRV2McyDwjh9m2Gm5p9U/ATa7ZJbPQboWRljYYo8mAh5sl/hBvrzQByCalDmfj87DmqqeB4m3
SChKgZ4s57NXbRtmn+kfLinyU7ZUV2jfKuTS/c8O+xBn4XRFHue51QqSZ1ZxwEaFluRUhLgfBcuk
Aoa4DJfndolHgVRiHGlzJ4jBBacrkOSC3yq4Ba76ySad+yrTuvYEEVWT29/nAtEaRYUcEFBD3Xxv
MNAOOEJ+yX3/ZT62VmVLVUPZVL6epXtxButx0ygqmLQTctaAzRnWwxuOnOxi9O3dkjlM5aQJDzQi
bDoTp6aU8mYV+w1sf57saLYZblrUhBLh3/2jzdOTOaeyevFpGx6Nspn9ZfzYxvCznzB/tzr2dh7K
cbLeZ7+0hRt57dHeToHPae2ymjqKSN1c8rOWZBUEzaJACRbnUmfpIn82PKnWC2h8wJpdzW1X/fCZ
04trtktJtx5L3ZvnDf/SMv65w5Io6eV7y+pWg4N/F9aUy3LQn7fPUYBQaBubuiR21Y18uv4pq7/B
tTriyvtwULszftH2+yBV99yCQ15tCm5QrMs7GalWHLxK6yw1SeVbWKRjhy53h9zg50tiKJUmtGPm
qrVmMXpaLQYbSvMncR0qVdJwzLefsMqlgTRcFPdExLLvp99GduydVym+n5rXNAl9R8exYGOp6xRW
Xn89HNZ5q8N6pfrmerrxsnx+kNZ6QBVvSeyB7aeh9Sb4+Be5EIe8JKDaZ+fIwDzphferG/9zqANd
OH2OWh++v/x0Vr6d3pqX3JLq1JbRhWIlgqDKIEAJBADmaKbqUPWQ+Ww4Wy8Pq59BS493E1RGtc1Q
48toeFx8ZPX8xsl7O/9KYm6FUF5NxUswgnuPr/uC0xrCCizHgrSHsQfAASil/kxGsLCTZDtAA12A
Tqox6Flr7TsQ3uliiZa8ifp3+xuTKkggE2ck6k5xKTLd7tQ2mfA9ACMTmhn8nsh36n9tPtRPl+P4
TBrLu+/GLK7uY8FSAThtzemPBQbpN5g8WrELaitwkLd7Olh7zb+5RTSwI9DgQTZynzfF8PJ8ZFey
M5bJLmGDoEUqaQWInjy3ibEV/zSNb2FPbH6rHzUdB47ZB44pvk8K6B3dnP9BD4+96XxKGC9tK6mV
jd8ncCI6S/VuHFmmkOYzfyDR52GsPsYoxi0aUiwPwuT/Jn0ygnRhDfAn58lHuRyYhrzzb3cRJQvH
ETwtoOc/TWxq0JO8oQKxfD/3oOzSfxPzayczOSSzmHBysSNSXcTsm4y/7e7rquWPB3R7Mst/OFmv
DaxgPBe9Os5n3Ynq+n6z1pScqDwfKQv4HmDZdCmP6orcUbP2pUANRCkoOYffEvNqPc/YJtCu6S/R
sM88NZa05keb9GrUfDvl1AcOOoEVnCJ5eN5Xz1Xihiu7I657VbUiU/nsvt9Im3uOGWaVFO3nxwsa
hy2Wi4+ITW2JYpgPZO6aE+Spm2j6M8RT2Oq2fE4Dy4LqTFgdV4Q+T6eJORPBaH16f6snmQ4yBqa6
mgj66DoO5Mk9c1aDwYi3KStz88SiWlERKgVoNAOGNaN5Hat0OsrMhtk3UWIiwH6SnG/3Rq8u5QwL
8k6JKRmR2f/zZK1NQ/ZN5BVeTFj/iN/CY3TuIbQgQj9f6+kIoF5OzEQVVdA0sKgoTek6su2kGAUX
Se5vXUqOCcj5pyqZZtqG6RGpHJnoPrXxqY7KkazjxVdHojMZ3aJSdwnuMjIrdgFm9tLz+CsaIvpF
gvdnu7VdtjfJxlET5vujzF7n26A2XHIyVrxTBpZmUQ6c3UvUnns4kiQUXRJd2BbCeRzBQ0YsZSEb
Nv9VrrB7grATfw2ryp+zJguq0cH3NOk1mpj2UOcbA8LTw4Gyx2SRJEjnhMNbTMfokMJCyKUYovO+
H9Tw7m+MtlEUyF0seeewYjVfAcuEmyHgeYSPY622NxQ6qnPvnk2F4pFglnQM/L/mmyx3TGhhdSD/
/+xqT1sqRhQ0gshI4El+QQZabVXxE5H/4VRzOJhtBblacd57mzq6XhP3pAhtpm4vf+X5md2MRZcX
b9osxe6mkO9SMyQTEVm+MJZsF942nXtYPPzah1YTNj/avbFTJVqHM/ejc95orNThvRn+jIiTtBik
F+/3PDiogy2C5/91Gza0IhSnyI+xC6DqWcoM+vITYgn1tlmxALbglPExyANQddeC/E5uQl9R9aM+
I69R0w6IA8sthbzpDQj7+nhcEcomcA9t0ptcJDHS4BB7mDp3r56LjnnxjP0/wAl3fOpB4EwTp15K
BI5++cikZ2RAKojCJtLAOdlw1PYMXmsUvohqHGfGDZL5FBz6sptfX8JRImaekp5VLYGy7Lm8VVIJ
WkptSzQB3rLgQmuYPIwCNQ1X8+8SV0wyeHPbITE9E7/gRun4gbtM++oPKvIg0TEsH7gALuCVXe3M
a4u+ubgmjHs+bDXMyC5FVrFFqq10ROBCIJ0rV1+1+huxdlIkjJKPh4eT7y8SsQbRHZ5h5V/L1mne
A2bn48PcIsW+Wk8W39FGR7p2zKyV0lrjrj9FcQW0XfHPItnfcZ0dsz/zur1rmO5anTDwYFcn7QIm
V7tFvzaDPwx8Iqeea3P7vYUlZsNyeoda90OrBGHncoLyftA7c6KbvD3CYjcqkXzqigCHLZzoAljz
xG7r6fer7sDGG5x0U0i3NlOhyZIWEKkyTnJmYDJ47b3sQwlZpmyCjbJmYWx1jm4UQDGAZl0syiJu
f8E+Jvsg2phyAKRTGeuTv1UAbVZWCorB0Jqy3Htj+a31sSMAQoPEwXFi2vs74ErcjdlRZe6l0MMV
GOoGBFo1L+IZkuUprv5O3vX0kh8SPxr0PW5JdCK/DISgJVkFNheRtWu4/FpnuvDV+950cDJgEL/k
kViA2N2PCfsJa0l1xFZl1ViatNtYqfokpuLEHUANBfBuSYwZ4WumMxF35Ikv8sB4XmPp5Lj+dcM3
/+vaR4RihArFjFI6R26/fu2dM6U+KdydTDPxXAFdJJ9JAmz+PxW0YkuEng3lBDAWRnO09DLuehCX
5P1yrHd/fesiA5YQpaTlUCk5elQ5O9K8yEVatOd3xi3hGOlPRqX5D2oB4UVGAGO197DsWvjBgoxX
080n2q7a2/IkowFxT7N41alqf39vQ7NdyPNK6xUQZT7CDT2z4LmQ0oZfwRFeQblYgkY/k5awF+jo
fz7waVF3/yvH12LkoCRzU7/3ELMoR/8FonteDsExMzZEU16MijIykpPbT0NFh01JGQE76R5wNtKK
LD5q91c+Y9rX/dEZTSHQtd2LgoNvTmJoftAzUPsbNCzJigjVYEcIrfthOgnG5PeWV08qSTQfKOTj
y7BaAMc2tf8RBqfnz386JZKmO0QKC5t8aSC80R+lcDAnjEB/4WWjEYv7XDhUsyKwL73Yz4O47GsV
D0ifMda7AzP+EjBBDHfJHmiAlvibOIKc+F5XMAiallczNwp0/24PaAmO7A39kX5iUf/8N8UtSMh2
YelrtyG8SrNbmvz+TrfyFoNwfJ5qNFaTH4B73vg7+ewa7JepsQS7/0Njff7lSwGS7r30gLGv5E3v
+rEYpFY4FjTyxHZKwRazK4E3QpSCE4DK0xRUTYzb3WiWKKnyLlznx7CzvSdqkOKzh/UIK3g+ycJV
TOybAMuqKPuncaODu827UdVPlzgjlnL5x968VA4ZhsMZnZ/2ci1n6WEXGRd8QhUN5ngePIKEp/Qt
q0whgUzh4JgcfwqRDa/oNhFsCv3j5F8bcQo0IE8XRIOQ8GFxA3e/+Dfyw7OJSOfhsLHq33qo9SOM
JQtOPw47T12+c2yNBYHayDX5xR/7OmwdPOYf5cpZ73tGhmyMcbnpabmZVEkmODenqzg2+UXhLZ8V
6Lzy3HimC1ApFBgmOeI+78YemxJkwf2K3GRQddr/5MPAn620lycJVPuQdBxESBzzHMvD5DO2zXaC
lTRwukd1af1a/ChiGxiBTqWx1OA97GDzJmSVbeHoBeKFiFSkToMbZIJYHiSiYzj8oX06iJLcOx5k
moS5//EQ9zAKLjAMW7/ZX5eEEIB8jDr7j9+hLH7N4K6yl86odBGGq/ISTQ9jz9evQUxiVSWcSOvf
zMdSg6nzK3RPkeeOqXb/a8/ujQ5xdwiFRcA6TRo11eYuvFuxGNovi5HS8oANSUWbGQwc3GPvsT/+
mTG4PNLlpTiRtAcOl0inzTL5LLZVt85NVusFNnrTNaeOZgUm6RK6OCgVDvcbuMyty3os7rMk19uc
pJhzPR/1F6vU/JxQZgF2uoBVRx/tpn7Fp+nSoC/WYBIkPDbAAXHNMiBVon+Cw7pMVZxmHfjAee3S
hfVR/3wt3e6ZFo4gDiOHdvtnmvZjcjsDz3uGo6wIUXV6mRRoYwuOPUH6pUMkIZQFylpJJjpXWX32
Khlh0i5SuGONGEBkpnsMnBTn7si84xC4sPr6Fw48xbB6/cbNOi6ZhVU1FF4JtHljImp9rUUYc4MB
Wq/r+shJNbI2LtcSdvoXbz1nWP1vfxYeVlQDeGU34wKORFYoL4Oi4p7OfYPlX16+sst89D2MbhTy
mKTbOFCF1HXg/qcdXWx4py5LIIk5GP87TUtDXyDav6wdJId93C7HsI2wDGqij/JeS4xbNbSk1Yl3
m4j8+0LdqZvzzhd0jgIJwv3rpUqXO978tJ58D0h7Kryayt3FOJO8kdl5vsVfD3KTs6BW3mL52YtQ
dXJ3/zlIiKg0PBRKRHwckNGJRJiBPVBmfDwQ9r+kk2nRGJVhaYbpOwnxbY0EyGnJCRhweXmnUn9d
FByoscqrplHDnnxaGEgrcr9miqhYdKn1mdXmcWJAs9padUyos54hm1KG8j9RyzOuziqyCFkiFte2
HHvhzt2XKS95QzzjaCyD3kJdsxOiOrhG9IgEPvI/YfsbCAUy6x11bviCi7QpwCi7q5FdZFdocY5J
gdQDPKSB1E8Mn1+OKjmscdaXmHGdWj6EZiIBcIPGOdw789s/H3O2n6/wQr+tKIhjHK0DOAFDQUaJ
o7ylUxHHPIB1j+DgSnj4+/Emt9OrKRlP/5uD5KNjd3cnmbp/MlzFPWFJ30M2BX9lHu/MmgHZcvFl
5gtrexLZSGbMxzgFTaNyx1Kg0IiVLWtTHeK0/s/oRRuMyjiykA8GE9diFCWOamt61gWngscjxhhj
+xU5z8zm7aSGhBWQj9qTq6u/xPrGfrV2RPs8Au+qOkT8usTMv2oGDOlcfLtY+JmXu7P7oZFGAi7E
FC2CubdwZ74qKBzmZaLRbIyPk1amKJC1imXVcdUtWstLdkkrsopSOueizQtgBVNZfnbiXkhgeA8m
2kt2ezfNwcpwjjW4mVFCMm2JaDW6Gs4XeWWWdpxEHO0IoeptJB9yb47hS1Fo3eOVq2SaGkfc6gb4
sjKRffkn9Agf42Ik912vEzBNFiwY07Bsgc6ejEl0GFvPX5VVrCDyXzSFLwRa2+23iWJ8FbOcoOHH
U12iYawBFkU2KpPQ0uatLa9spWMYLIKw2weH/JY6VDjwlhgR+ka+7At0hzjxP6WAEoYBBIFbDhMu
SQhLEkW26KRK5G8H8uMjmJK4onpf9rafqlLYLW71rdTRIZQG295LVsQ0uZ3USxa+mjZbFbdXK7fk
0Ok8jjB9D0vGiOEEYnbinH57K2DyQEaKDZIAz3oYYAM5cZe2t6upIXHinQBaYe9wsqzLe1yMD5rU
sdjMIzFkUjXFhcEfS4XvNI9G+NIjgbHcFCUt+ZULv3psuoC/kWHuNcS8Tdwh45vb953mhAA3Y3ri
mdn39xrH8PNT6f7TIUNjfmplohs3b97b9IbnYqMAjAtj0LpwK9lXsoT8hvpabtK7JUtlaO6Avi/a
hZsfcrCb2eXPbqO5WDAda9B6gjurvHFnFlIO7KeyoSiV7YZOcVgOrU03owbpoGuD89OnE2xg93Iw
ztICxy1kvZndHs9Q4Git4gRdCIxtcH4X1TSrqg5zXvXY8CtQrzlpDiJp3/7N/AeSx6A6i4qkvTLD
H6JpmC/wKgOzBHwqe7v8svlTi/wSmE07zmehP12mbEPyfWiWwJsVzqamq6pAH0IlkRTgewoCkLVg
mXaiQJzlx4X/RhbdcJdP0r+TgkybIqO/NgyWF0W0GsnUTh8+E7k0d2t7FmrJYfbt/urPhE6zvj2O
xct1kpGiSVf4CH19smbqal8uoEEdP6/AOsE7bUllMLbhq0p/RcmfRJervHG4cUr5KTLyLCTSFKIX
Y5imWF/ulMzoQjaYDaKyNn5VXabPMwc/3+qdlQwSe9IQMi6Kcez8avoryPETqGOEO89DI+WxucnY
pd1Fb3fozyGM+UMzeFoA7BOuO4RWvlDnd/+gRyi+iYiTmg28ntUOjbvg2c2CQf2fXwaue6iPXO7C
uWvjJ/f1ESr4FCsO8gSdlhiIlUGK+pEOeuX+VPKz6mAZzBWSXLHi485CNEpzHH9B31WoCSWjml0Q
Wn7VdQA5jag7zpnIlgg7CKx6VwXs0I7+TjmSgIYwt5KlNamDMx7LT4ISKt+7BoiJ/v577g/8C/Yw
H8qCGvzdsCLkm+VvtcFzvvNhsP7c4JWzY1IedzPMBfRdmUS0ABP6bKjqPZ6eTg4wZIgQ/dvmhWUO
1/H1WnPrn7pjufdtgb7r+0RXmfo2bogX2CTifbRbKX3wA4V1jYq5XPiZPTf/e5DabvdpjL1gQd33
iDVPYKBgowy7PyjyTuWagv45yb5SlEofhmXkumG1kI7x3q+f4i8rieIq0XVZ1rcYvCp9e3sBBLSD
mda/kPwJjzeqTkgB9uKs6PYIfFJHs1YpSDPoJIwMACQZj8pHeWfiWoScAwtiXVZPwlIQs5/4C5Vv
Q+9IrZFAcjy0XN5G8zhviBUuWEiaDv3jPDhFuf3m/UuFYDae18rHuHdSgWNVx3x9NiBAMr7s7Gcg
wWiMgZy8SOZ+NtwsaX60ir3NQkALRiEgNbukVxNEpgPnUr73wNPT7qx33llsLtvfpM0F1BlMsC87
Xcru30bn/syeHwABxndC+xPDjTxGTH/6V2L8+xFf6Fxrn22omXdmqZWIVn6XwMODipizKJNEmqoi
K5/g+08zpMfW/3DHRgYaN7npK0NcnU5btArM5gCT54cDNhZGU/Vczvh3VGw96bThn0wck56qn9Wl
92Yu9v3kJ4nGWh14hTHcWpVYEuDch48AGJGr3uJdyrQ7QYaeZxhhnDuWw1IlaEjeI8X4Y2sKR9XM
vaaMI8TvCL8f4dkuM0gbSyDnf4rnXMx6qvk3i03++MaJD6BS95NeZREYreGOpnmo/V2CI/3hCslc
TfXOxXKrgJli2R8IZYn8t58RGDRZi71ItwLBJ2FBY0oAiDR0UovI3uB3kG6T1xVdJB7Sayk2mayz
aXynHqsRxxiBFbBPK6x3VDYFMFvbfY1nQuzZq28hhGwOsRZDLM3RR9gsCcLnCcG8XgqV/81jkfZi
as0/uKLfoAei9CpV6ErD7hS3OxjvMVTT3k1HEpO9ALpn3+PSRdVRJ9yiB//Wo4OSk6myNqQ9Sbyc
nawUyqvM0AqkWsCdc1QTUwq6IsqWWFY7j/lfzhT1QDATPeKZC7aWDiCOy+0n5qIYOodomn9luMEU
oiqHhscNKZ240yzrzIWfsllTYbCDC5QG1gWlKA/3UAZyRgy8ZaguqOiDaoqzq3Rd+ZKgQBaKECyM
34j2ZhcU+51QcO90JgzeJSMTP/p47rKOm9uBTvYyWCaRGFesOpyaCAK8FT3TP7xHPHwW9CxyzjtD
hYpnriMq6srJcMxOmzsI7XgWUfpF6QjC5HLeYv11dN2MhKEC4S7TUs0Pc1DmfUBPYCejEZl1lGgA
4/A/F59BAF9Y1Zvr2+7hBcCDOGy4SCYKiYQpnigYUrjeoXfKoH3xWORzNPp91lleZZGWl44SY81f
J7mS8TN5cc97uXo8rrEA3bZyol6VBGZv1eopCdMPpTAo2X4JujaMi+Mz7BEjNdyPzOGkN1nF77eZ
gt8rzYLZ1kVJb7Ng+WnVFm08BOP1AhA+d088fUaZxQ/9GannEzY9KQM9WCHbnhTIZ8Ih2AJoRCwE
UxMYrT5SuOsqD+lsL+oT8c+GSRjoxOMTm6KEB1KmLYUCORuZdYO3V29qBDJvOXroGP+oMemlbbbB
wk1DYNWnb14rZBl66ehqrZHxiNWzARc1hWoHZ/yaWkRbEHUghVueq+OhhA/6GQyzC2OBcqqJ1zJ+
W/Pdm7zVEXKzzJxKLi3PrTXDhM/y7Xp4YHShu5m4VphqFJ8jxEHnLiMtboaMZQ/WfQYzdY1fb5tq
z5a2Tj8N/HjE3PgCi2ICEr6IDGKbyiv5gqq1SKBnXItdXL6ByX+fLJ1bpO19qdC5rmV1frXnefzR
rnoTkxPORlz+0eYAL/qW0V9VtmXTkDax9ZaC+wLqM5lJkMOV2m7p3lzq2HOlD9YopkhUEg0h+C7L
sbICtOIbgqpVY8q3LGo38H2xr98KkzBTxxWbXKs60up2Z/VQKdUDDOmTuO+2mZ67AkUfSKSY9LwM
OxxVdAD3CmCH5l13wvLBx35FjsYeHEweOanjTOWOnit+SeHwuBcrgFjR8WUHyTtyWDIbcEj6t8WV
MrRTsDYfzDIdIAmA8iXvw5i6wNM5r7v2ZmhQ2U2EEBwGHLuTvbG+tzb0k61Bqd/MuqroqVJSOYGU
FZPDe+0WrjamoCUaEMJzoHqvBvojIkxRhKQf7cDiYUW/SEgbhEoEoueh5NNBuMt+BXsEsvcuW3Bn
9miMQRHKQ6oMA+oqHbVJrPveyAoz/2Eyh3RAS3wlXyUb5Y0E+gaAp9PSmfEVbBRugTIrcLFso/My
6ceg05LUvCwRItnR1ZhFQxIYT/FjP8ECCvilDRHUShiEDVCG8L1bvQym7zgIdCFZ9OTCnmEYChr4
d8JQSCNcHIwo7swvxenXcEY/Po5KWwjnI7j/1C02amGDpcB76K1QFTpC5lTATOQuOUIIjfs15WKn
5mvdck76nzLdp8ZfqJyrSwGGSyNngT5038kY8GvpNMJBnmZGjNe+OhOZ1/GQcWSmXG1XrVAJJTNy
7GFoa6j28f5WX99UoNV1rchHGmg5yWz6NBpjpyftq2vSXmQ8mC8t9Vv4I2WsOpetQH6VP0v+nSmg
7ynOPmeebMe8zeNMim0mDjoyy8sm4KI3THF/6couf14A+2fx4jJJr3KX00EsKXPxJzPU7pCRXdXF
n1oFm/cfjNGZgY8prb0I5khUaJc7WQIm/Ic6Bwv2cLOmRTeoLE1el5blrDKqiedW0NEqNT1tvMGy
YtByPefNY6DeiGWT7Ul1rPFi7vB0wLC9VGfOJr56Y1PFmTS+3Qi50RUo4Nd8dzeq0yAhdCeR564j
2/uasf5kODa1ApIoJRoj4zq9PYuzb30BlzN71TsHIzE0Cnr8dsscbVetHNaOrLhL/YT/WxZgWEZW
eA6uTdWZonF9WBkqES0qAE2YOQObL82msUXyXs7M8/olxJ+spqdT7DD8mSCuv0GjL5ptPA2RGUJh
qgS3fJZleFK9kWSaeIOtqO2egY+XRPqMYUsZkKlBCatmVVAWWJce/mW3t8qwKMMlULCFq/bLS1ls
b8jhbpdn8NiaNYhAcqZulRI0JZl+2l02sPjSOqbLwbglIhezpSz5QOdinjDKYL5hw2JS+oSS6IAb
iHVoSu9wlMl4CvCWZodvOx6MfzK0MvKQf3XR3zP+kfg3xq8iJuDLiLXjhtNtxcXm8kUa/xybpqZw
Mi/rOGqUVJUqNOfAAAk4Gr7862I1qMXD3AfL7P8ABlVqDmAcZTDYYq5PEaPeelNMaMTlMyxLFK2h
DySV8zdDbJ978d5otx0tRGtpCNS45NynvZhmYNMCrCVOY2OouBsskTPwLFtaJJg1S+cCy98Xy4iC
ncHRS3jns32HqjzzmLDszfXzvgG4fGXochdrMQZylrKmjtO2MMcZ8eA3uD2d+AsC7t2vQ/lSbhzM
nS6SQPcgHy3XkXiwLkYrIoycsS1GSRwx0rT7URSNYBQcypelQ/7FAkOpmwm99lJvJGJWPakxupkR
zwxVlYXM74aRXjV9qiLtNivtfZYAYol9sop8Z9GOXoz8Iy32X7CjaSTqpx5ZEN1fAn5imZCmk+/N
bqQ8MRLqNcNC134nq6vMYFm+8hFH2Yz74ixmPH/stiOw+nHK0rgKGbMojRcJ3nqbUapToNLjao+N
NcX+lzkc87r2A0kKxxioAXvk8Mb1EuCzbruCjHxWjV8bvLAqgC+s7tjtcUPIan7BIhhKej2JsMhm
Pvo83bptgl7rgpdJ3ywre/Q+EaUzRXtJMcLJ6BHNwAGWJuRwS9aN+DcsYH8nl+Jv0k6XVhXu+pog
mUiGjinT1a90Pv/0hwf4m6MbcRy6d30+YO7NlLoVQkGqKlwWwoT8WMm8VzKiN5ZKgxW28nn8rgd7
YtWcHvf8qZRm2vKZiRRTFC6MLK79WVjeiZ/H9k8I3wq8M19WtWfToRCB7rpVc4N2GJKgjHbI3wJK
8G21TJwyaJEaw0KLvYOGaltlFxBsBHwjLUApVVGk1aXHhKE1Jq0AITLlR7aaLDhq5TP1jfdxvhWi
x4zgw+Tmb1TsQNc0nBtT/pqiFV2XfSEFArloLlp1cNw8i1XQTJSNNYNfoXKqgh1nf+iwA4ibUkXf
NRGwJ1eve6IWKnqA1vzm5Oaq/fxZj4znZkYBPbcEYY/eoLdNnqC/D/+I8m/uQp2J2M1Yaqh9b4B4
GKElBhCAraRPeqsXEXUPvehk6+wKKN40Tn823JhIeTEyLANZWZXPDOjpcZ8IFzBSAjvGbEDbWnCC
YRNNY82UalCzKVibHr7OQgNs3U2xbxlaEsunxAVNS3kueDQDnomZqzOVEYyjsch4E63E/wuF/1+3
o1rr0gmM2cyewdMLUOoLZVDYvlUlsmipUBxv1ONsYIn4Mc59IYeLF0NQM974nsywptZLm5Byor5v
IVxlfozPOZDz+NAjceSbb/jBOPaXqVO04Y7ANYwlrDnUvnrYeeNro4WD3qfAZNhxLFreUI8SND3J
qpOw5GNLwPbXREeve5Bt6nnDfzdpOaC1Wjk18/o/53SCMeAeCgPC+BUQmBR+hQE2CJuqVzEEPxYB
Iw78d3tWDr3KCmxUymehGGuPky5b6bKBXQ059NzxLX7/Pi9Ra0iY61RiZ36Z09xpDCOQMfV1JqqR
8JigUv8Z9Us0lvUZG0AGzskfYvQiRhhsLy0SACX24acdrOJsT38aViTYdY9A7rWWuscv021rpmTV
sXjcXvWuc36TIt05Fvc1hK0ffVOk3VsFM5D64kqJq6xlEb25kwnf/2qNQCOZKSzx7A92IC3RDIZs
ao3hzZEsrOywRVufqgBlL3gdeSpgr7cqU+26qB8LU5wPulAxl2G/I+69gZUQBIqGZ6EEtiZooYiS
VynrBdXqpGbvk7dnG1Hz30b7nQrr1aGLxlJ3Sh8KsnuLwx3xJSrWd9obBNZiiY2+8pOCgyOZCnza
QPKxZKxUUxp4yToAGe2iNeTaFkV8axDvcyZiZNMFwcvuO3ufqtDcpfedfXH+RtitemErWfv0VDyU
Ugat0fL+oR8fMQuVghvn5tTYEreClRRdHU20stNjcwodAVJn/gotLEnVPqtIDzpVa9u+QefZ4rB7
knmzKGuXqNOU6UxD7/39/GOeaDPtcrsUK0HE6LJuFZOdeoIH8j+e7MdKB/P9VNodI14c7OGV8y/F
ia+StO5RnWNYTp9zUngSfbxUMvUgKrfC8bzitMu1lSfWUgRULpLElckIZz1+KognYuvPb6RPBFBj
WMDG+bxXt46QYaVkt2HqvzVjV4O8NRbcD3CxjhGSBQ+khHMN2VM7n8IoIySXLqJh6zoZGWeq5g8p
2F5ofXgYCQKkh70bJaAUNi5aGM4mMQNANCAi0Fmn+v7qoYNBNErrQAMbHwHs8mNfkPgmRd/8gvq+
KPg+Z0H8EqnuWorhXjU+wOOFAUOvNfKntUUz7L3f/xc8QNPltgdW9UaPCeXmQIMvW3SWLXtub9ZR
cO2iVslMIyeOMquuMYy5K/8p+okMESmYcEhiecj4LGhmdZRTGg2zIzzDJCylRsbScCVxOQs1+1G5
RrJIi1a4Gv+WDibMUw3N3pz9/Mqa4mFZnmzYfzEHwFi3YLj3+sacQBMRyx/+nCZaLmvJRg9Ck3B7
sO59KzYWi6wM66gcY+9A/gID+xf2R7eGr9vH7jrpdadRGBV2UgjeIW7IkmhUORbr9LIVINNLzHkA
TFEkaCJJOR91eG0xr4aR+Qb/YoPWOY+/KxO42LnFbIGmJHoLf7tAnYCUGvRZGNHHqeqokXZF6ylG
Fo+G2V3lJL4uxZA6LixurFfCyweLElpkWV/60sFkX3LLzgDOqwhe5DODa1aWEMyDYezSObmp25gS
JSHoGqtWWMNX2YxQcouvSppLNcmqU8ULB1j5WS4/23jEeND6iRfhWhh3by1z1W1yUf8N8RWJ0Sqs
d+aAv13MD5sRbrSWX7Aj2GpwKZ9HvVE9FuzoJ/NqjHo+axapRF46OrKjXb3kubct7F4v78diO1Bv
wXh01T4JAz6PJh1fjaIPnI1Dz6oGSMjXIYbW9b+b2guq6wrk7153rvSY4dXO06jkGPEcatMplw5C
uOw9rffYTfcxy/9NVFr5wByY5l1nM2A/PWf3fxi1WHD9wTZtDVYGdS0BslcghsX3xOEJH+xImtk0
z0+L2KYVtO3+EqiUK9PYaBXPLb2cRid4W0NliOKD75ocvtsFpT6A72ndKwv80HkmLQi/EN9ll5Sa
w9NlutRoPSkYk+OyVwiXPsZd78uv9m/aBB5Nde2/oCQGlfUBgTUzTtEQLctf9/nH0gVWqvZCrjbb
/GS/4AXOV7r1vjmVYInP3wLGzcgaQPzwUa6y1dn6fhiakTfFg24MMkwDr3ox5sseNqHsbUF/qnsB
bvRTVJFxoGidFtR+3kYxXNJyUEad++rdt6zU2R0khB/h3XGOsgTO7LLvcEZdvqlYen7ujue4nsjY
4lfdvBp3HHDP+aM6Kg8n9mJI7Wex1O6UxZhTfZI2XQTpgtB4YZbOf+qOQhX+TQW3bqXBrFIkzPCj
xfmhZWnq7DEQ8mY6CS0WRPPJkyDGDJaasoLDDzX5DpcK19ETl0l2GDjJowRZQpAJgubPOtrTbfb4
oeRkThDBtSMpVJcER+Xh0zr5yTGcVZFAKFVOU6qndX0BKnSxM+crAJmD7h6Ck5E+brOP9TiLm4dx
oqehhEIU9HgpsKOjBjD0VnU+2YB302dFlyfMBdAX86NrjzhZNht1a8v7z8FEPtaaQiiQnWV2rw0h
1j7M6XYcr1KTvylWO++AYyPhUcB74gs9rJ8/v9ZT5sn7lMXS/HOMZrDaKcywQjwM7stKp7kM4vPb
rYsxirqp4obOrnRYSrwPE+lrpEefoIWw8IZGW1dnWTXkHzrkRMSD2CYchsNYlwnR1HWrQZfv8u5Y
vejufibSI22XdwhN5cuLwerlH8GdEjo6mhzxNUdKIgpP90X86azXGWpY0EMUFQVoC176LGiPQXhe
/WmAUK2s5FZZ+z4Ykek01VSgZfdaL6gF7ldynOAZkhxZ7UYvxb8/lFlrXSuXd9t4YGsA0ashTffH
HI6jfqKrc9DiJAOQYclAFF5MPxNfSnxFNqxHwqarh/RF6ju65I/9fs16NaedMl96GeGTxREBBb7l
BW2cF7APLxZj5XRj33szdwfJV2C4aU6UHTqQ6hmkVEBmxdtbllm98bs9H0j/1UVrfM0i3qIFqyy3
Rc/zywqLNAjPAeLYUWs+rDcvub1gD2/IgDO5+O9naX09qX/kGzfV8hK+m0G82OvNOBqxsrJsOZS+
TYFidIjS06/lu8pWcTW9gq4KeAnfpuWCVioMgVMni6RGESc1uIPZQVm8KmFvfC7pwMEghJeRPRPj
vPdJbXBqRdhr93LxQb5ToUpVkxU2Xu/wDWQY0oEGpaVcTwLdLO7diaMwt3usBD2W3/ywvI/fJ59B
4o6NC39Kbk4Tn/yUDNqh4LIvQ86W9p6T6Hvp5gkWK1R1Ql5ESahY9mjWhvdm5D08AGo3kYp7l/2f
ZdTLxAIlgt6Y8p67VrZcFho77zYGC9H5+hpJ034SpSPEjJ/fLeTF0sSpqOTBMC2cr/csA5HY/eg7
S1Yv8pocdWpNh6xaWAPEByZWt1/LBUOpiuAx15tISzxIBQkeBcl+QMcsYtmNViCRGlXJLmjMHcVM
jzcoDUZQlaxcpVtNnAtOlv5DpbMDYH+3oomUsuphtu7hm1uts2yFZXleoctMgRdp0mSd01JQUNW1
NtoEK18/PJGdBhUlVMsYXKbUNkltlJ0QVCO1ahaCTKDKfN9LFD7NB3zVtBs/Ke7crlvHSdQMv36e
oaNVSRSBaHZG7M7JoE4AXmqG0rZbcKNOGLHr+zIbWwbq6XEqlOf2ubiY/oAvr/XSuNYyT5dgAnka
iMvX3sggMCcW+bWEa9sEY/62QdJgQOnOg7k3JS0q+Ha3TeYpn5rvwx2/e5F5slF3YzLjIM//pHgi
OpioQK3BHyhdqZzJv6Ov4ay2ph+I9VLwU6rhyicIXjN1TxlnML8++tab+hDZ6IGnIFCEpYVHRt/Q
RMm5xq8TNe6CykoU3gQ9BB4ycEZyWYAqVZ008SzVlqPUvrb9UTdbNhQhp4UflLDv5NkTQRkK19wj
qOfQ05djaJpVyZKleNe9IiAJLKrK4mcY7f/RCWqPYc/uj32Y9wLkh0+rzseHZONez+lkZbgRzmI5
agZoOjEqrVOtSQqlE73ovnHwvqu0F67c/msI1ErYG12h6rNMdE/3h/tpFul7AuVxI2dS872ho7Aq
WU45/Gd5xcS/gf7hSUQWf2gvHXpw3ceuok54a/kLrPqH+Upp88phESklOOhJs0BmIpnJ9CkRHOqz
KLiY58WxD1vPK3Fz2jCWfZlyJy2+wKvk4rlLPN0VXdJ+Ew1L+JoF6guJr7rBbBNlVIg3yn3Bl5ar
TZbfFujGR03KpRscPAmRuqszXn0rcuqN/7C7CENzjGZXyl0oHLJPk7l6Dlxmuw3NrHXy/hr4gbZR
qlFqXnR5v/w3KUtkt3MsXV3Lp6M9LPuFgz4mHGcQBRZy2I5LHm+s4U2wheSO2tjiGyTofY4rEcot
vGCSEepq6P21ZOMtg9K7UTHD6Sx6/yt1Ctar8wywPb2vge7e/dnkdiYywQKXWyqfYeQcOkBmq3lf
yQ8PkUwol1n1V6rrnw2FXfU92z+ZoTBOweAhVim2M6FM8BAbjwJZxppAGFJ1h0ZemG1iGGkmGncL
9yVfEpyEx83t/vrb5oZKCR9Fvt8NvA5KvPwvJCStuwMMEpoj3zixi10JCQapSILStfpBYnLcZvkz
c2oNz7Tbtvasb5f5mPJ/P5t8KHc2cTGOg9B0wvM/BLNNiCzAeHTNtqBdEEdCDhfSQ9/FY+KnC06s
1Os+Sfl2E5VHzfe0uQ+ueFBwQOVMDHJaOGdaXHMHCRO+4yVWu2FyM9m/HfZsmWec632wGSWxGh9J
M2QegfUR4MTR7fgneya/2+0dGniRguKNFq4SJbrd7sEeP5pcymxf9RnK0roVEF+6flLY7lpUX5ys
F9OayOIoEDmK6qAwsVJpr+TXLJBVmkEuzbXoFm6Qtpe2F2vbaMGMoMfh/Rcz0Df8Fp4YUlwjZ654
+sVkHaeING57c9rAf9VJK42sOSfE6FktXi5s0TW7lm6GuQwLfLmcipXHWxbJM8Y0JcWg0FSRh2Jv
P0biG+aMuy/mfijSOvpkiHmRB8KQvf7tqNhu6o00SCkww9SIjwjoo3RSR4iWoZaVG8+KRIXD0wJt
vO3fjQ5WXPN07wBm+zKR1AsWHyhhvMb8sqwqa6MigcBGWe/HC2QeQ6vT75x6oXF8rkpe7JGUQFe2
VhNZqKq/V/LGSFMvuWUyS28PG3ijX4pKBKUdDOgO+lKTwQdpupPLUc8X0IAwkBf1X19J15ROY9n4
iX29LTmaejqcVWxhSu+Ng5Gd6bffXnJtLIpA2wt3qTy4qAvfoW3CrfKC2qAHJTV3488+wLtt5JOe
qY9IRJ3Bdkgmu+ZhYwyfiuTsOHl2jdUPclxVrlmLnMPZ12OPbagm4PdmgPVF1zyhkVvAdRelxAzj
7upFG0DFXHR1xro+b6yaKXzC8G2jRsNR8FpcaxOzbKRwMPJnZWCsfFpXuRODW1ifFlovjvQe+Zc6
latok9Umowu8fsxT1a2ZhGhbQvN7Y4dLQgwYX3feQrJUDYmDGVRPrFdGVTJ08yLTnDBFK1NQXB5I
J58pLj6JyPKJCuFgmAyZovaBq1cjVOG6c+Uv2Fzuj35Q1mt6dSzHmbIY8N6+xBLX73VCD+9Y2Mzh
vD2QPUBsCRO3qgsG2bjyREfip5XUyRq2TuWABNNa9P1vjvXH1ZCleEIMs7OxNhwYR5KtpgRCtwq1
0KF4jPepCEWpk0B8DzpIBVe/t43FWSgh4LOYl+Vd2zaSoUTHtrXgDWoZUtnWwMCpXqj8v5eQLXEz
kJpbYQOMd/aP5oAy47gQae5C3jOBCw2/Vhwbh12RmSn58RhfcoZzAikfm8UZsDe+IeA3SHzAbIOp
IVGAmpVy4pfaBf+kjXWIIrC1FoHToc9r8vOzJ32PdJrTB6ex+aUcBE5E4qay4Uws31YqyMXmwbEu
+60F0raWpUG9h+Ypzl5aXleTXYpOInwxU/8Uh2Kc/1wzUyCjD72PWSvIEN+vgCJU9EWhN1yYHmX2
TAhFd2xv2h6Gv3GqPVjrwxvCuEQddSm90iH8wp6JSxYNT07CGHwWHTVWIW1aiNrObTOZjvC+yzes
pA97BwT3UjJOGMSfVD0doJCr6uNawV9uozE2mhtJXm6enNWB931RKqBM8rRNu4aociKVe2ILT8da
OWjcE4xFvrX8g0ZNwOygqgL0qOb5ctWvnTgd7Gnl7dLHXbylJMu4hViApsCdYdri0uNudmIZmbt+
Zg1LjOdfucr4E+ENd+JZ5kmPK1sA9Uej5CWRYwNvwrLKuwnJ1sYTvZoNIxVO0a736VxM0wi5MIzg
U/sIBr4ToHWyAv3N2k9H/Bvhqiuf53FJeSnrwgf5yKt4EyWWOztar1DqAdurDmBCvWd/aGqoyew0
gwTl8AvHVIaIujRPFOcfP/VaY87SYQxdj2iy+etnTSD9n7QGGbonWFuY6dUwY6r0CAqXB3GlNntL
9P82rqkcwQ5l0eNukYWt5IVvS5GxAUO9xBCUtvsXSXHR22wEUQTR9j8aO55ujL4GxM8rFg769dda
LPdshF6jFUiQhhAStdJ3myrDwjzS46RFRIhKdIPzmoyl01GkS9JvymNZAdEG8943VUPBFCZEyfox
uq0C/knAW4MZAE7SR/SwH8f2eotkx/kYGrQCrE5LLxJ6L689TJzzKh1D0Jd9I1xqMmkqdPs3i6AC
DXy4BMEQCz0uEBr/zL4icfB+kKDkoESn5l/TkJ69NEIobWPs3QUYwOM5xrCkRYh52C0q3BGsGBX3
llpscsbtCjF2d5H7b6d5IMfXVF3vBzPeOwwUfSaVi3nwntnyQdidmHy/gKP/sigNWrSykh1lmf9B
ieDceZjZkoJGnP6C4h4PLcIkH7tmZ1MiH10JUxWSa00EnI1VgA6FRULDtoUJtuV+5CP+/n5xCugQ
+p9J4jc/Yy8tHyLujvvUL1ibj9zFGsW9GFhzRVEHkT7GsaodM084sueSuAPF2aK6Rtgt8L1zMUpB
22QJ9kr2pbq2M9TwLKZMVlUjZP6GsGNi5hxWrijIzY4pPFr+Ru94wcwMMRBLifZVjG8QeyxcI2n5
gQi2hHlMO0mVHJ1zPqSJLPscLAXi6R43lPs2UKf7FiPUFgNkyd4+RYa47zXZIlxFKiajoPrwrHNd
8SBKrP2cwk5IosFfCqFafISEh1MPXT3VMs39BlGBQ3wr35b+IY2mEvW2vhWFVgZ/6sgohfrAXYqA
iCgjAAMIZpZ6JSdQDq15+JknT3CNqciOzQzAyEAXvmK4sUxw1l+01c6IyA1VOIJ7tHDcYHpHDg/3
NtI0CSZuGd6dmypcShzjZXnX6rNA/pImEOXeyoOj+tKc6cmiIA5VBpmzo7FG2px57rJGjy/1YcH7
C/V/M42X11PBkT6pg8BJ4Sg08WS4ncj4lVbjBxTHufJfJwOOiLrKlXr7JcAU/JYctwsrbfxyV0I4
yT13I+8oGN2JOLhMK4eNTwh094uAsnFI4uvIZzBTpLENy1vvObIQGIwYTT2PESbZO4dD9oGH/nkE
98KuTRfQhsUpCNkkVJuFirl5pZFiD2g8pUolBIWlMXIqIlXPU7NPMfeoSmeLtRYF6rkSiL+rA+d1
GSvuyoQfIYUIxmuFBHIhs+4wdHptBPefQHcuegFMPVPFuTpidaufuY9IqB8UxQMv0+3h7qLHI+F7
U4LoCuD43KaPSMzwDUcjL8ABvk2ZcVx18evoj4Va+/OOvow624wWgMhBghsgNHDZK066QVWM/BGs
YVrBT/1LWmyqS0161XHBZaYDJ0eFL5s+DpgXyjTcj4v2dkHZy+/S1a1/5xqrHj7tbbApfiu1LS/L
oREWt9DpwiJN/ZXeLLbM3vEHVAgFF0SddZmljkkIUpO5aCihmfyJ9mSaAerj2d+GDiNxBXG/140S
qPeqxb1YQz8x4Zc/YrdOGD9t0RAcDnHKzz36HzKk1L8/+bQi+9V1DLRxR87PbtHU7PMJZ2rrdIPR
AD1H7peFAMONwvzlaYq39A6gLViqPnZ5EJALFl5JJsR3fNetUfSrbgRhpCuC8GzKfPQfMsro0KRF
JQHJrhCu7x0b6fHv0fwxopbZyWfqjxLeoKSseWk+Dp624lIHw9D9ney27LDn+nwnbwZ3CMQcrf51
/EOkMkeR/cOzIea6/Uam9mG+azjEBTVb8JgozV7vzf8CwEE2DLaxfKwwuN3FJiK0CS4tfiK8fJp6
kk7eHYLEy05JTRw3z0bwahODVGvD0BHr+5sOsZwhoGgisOzyLpplhKsz6ITXqeUUtc8qFSKTTwIf
BLA2CJKEtQUMFTAarOm/paIe2uMSY1qo2Z2Dc3kM6VTy0s/c2RsUn+dJvSwgBP7Zu/iu0Yrq5i52
jQbhPu+LD+b+CUcRONumb0Rw/qGzYObG5gNMIYogJPfljDCPu2v0BHwQONlKqtSExMP1s5aQvczW
Oz0WQn47gS9daOPv/M1+51U1NEvW2zNm78UUBi3mDz+lZ8toQh0w5P1ECHGOkDJffAgACGyYa71b
09Vu9LocWsjmOZHJxyDyjx166QQNM4RaC8z764HCK9DJeWbIdh3rgMmeTGhQA9z4iyhq+ip8VuEB
w4RNQouT/au4dT0/Rx1q1XOpZgGxHbKhjdLEJHTVHod4SuPz/YYlx+P3FOTSPuJpDdGlg0leajNR
fCEW8lVeRzYwoZ5xflZFvwzBzegbbeI011NKoinsMg0ljmsAunz5xRa43KxuKn7JE9eZ91yFa5f9
QZ6OLMNPnf0JMAhrsIguvTLeLlIczk5LCN3cH9ikcU892GxGmYrKFeR7go8FDBAMFQW7zyEL2ecm
jbxLmvkMOlPrqHjNb3O0h5KiksmHSTZ8/JOhyuyPr87MD2UlUcCNmx872mcnCthNR3/xqls35Ah1
3nPWnCS3a1QgnLnPzoS4s9KqdUDQvaJn4xw3kjJHbrUSev5M2ruV9cYOmZrUIZJ3TdCWitH218U7
xBlPmLpQOeBalJqC93JzZ4FgTz63t+YW2UXnyXDS4yxfSGaLfRIWpi/wrJwCF8oxcsgZOapw0bxK
S4Y/kFK7YftM1UGc0x3mN2fLJEfa8JmELkcyQDXsfeZK4YWDfJsgb2Mh7WNBfxOdq+jk3oK0Y7Kn
HbZcAYDBgG9dgLqwNz35pyTNJpDs8eIpzEKMKbjTu73mZYS6C6D0EJhGk+f3XXp5ZHzYt8LqzYJl
YFwTGcjTJiSYm9xzxnuthXDrpFDIfPgRmaceKzVt6olAzKiW068slD+CgP4xvfv9y4bIegeSWdQ6
oFA6/hHmIHBae+IV5DvyV1Anfon4QBxylJpVqrhFMCuhFe6GyO6tepPLcjVUqRUcUQ5iIru/lVEk
uenVoqa+Uq6/b202VUYkyealnjXA1pEnpxJxt4JVY3w93zWYuAfbShVFH8V6rd7hHI+mL4q6rimZ
Lq2ZlohL+V9fgn0NYeXVxdSmmQqwC4Ay2+eb8roqsy++QSwIuNX+SVPagDEHP+vfdts2n1fW3TYh
EmRS3qnlCLyWRMknpp2F8k5vMU0XryTyK9+RFJzIXlp0rSMPayUwFq8dn84/xwApqThZrLwpdUiw
Fd7exKWQqBNkGpAmn4ME0lwN9YXhMATDcY37/GJSBoz+ebFFCcBkt6r0JIov6lGAbMx9J/vvGY7A
oqe12CCy3PMyyxuxzA2Cf/OG0moUAnl4scYa96vSzIuvLYd1c+24OGvZoUGgfEttB2p+QSiwJDvx
TFowg2g1i/dDts4hEIl+nLlzd2usoZxzjHY0Z7/IBv45kbK+PmDGDpeeRgIM1KmVJtPocdAADIYU
SmGFUr99mdQok1U7gagrgAtyMSFHQMSMvNM5wGLuFoaLSBtUuzoH9VUGJi7c6dYaRBrOmvHKenml
jOG1tk4T8RCOCT6WAHCiqyTXvdCEoEP9wJNFIZPRZcU5VEpzugMVf/xHIndbPz7BGnQNbhGk+j54
1q4tORxg5ZjDOjntzYkSzcwz2d27XHKxEXmJCBM2J9o3wc8BH74fd8RafcfGngLsyIbw+eS7pXNJ
Y88CEfOFpwrNO2NU+sNWE8LE9ekNXwIrnR0HFYBKfkdAs/s4c2c+gGOAzBpdbVPEEP8iq/O9MmfJ
mJ/FcN9m8xjY4nhIqEIxe3o9EqFde7YvfYGgPIF3WZG41oi4U+zkL6C0Gbs05zlA2oyeHbrHMhxF
L78OP8aiWJ9lKHaSsPCPZqH9ZunpGS504S5R4U9t8zxgT+H1uywqaBabKf62xzPd4cKIaKjfsB9k
HtsN1jcWyhsYHI1EgykuIQDHURkRHimaE9IoTmGf4lw4VjTEZ0kMb0y4KFUOCPvvwJ7MBf+59Cx9
K8u45QyBZkVCM2BtzGIdXzlfO1eIE16uTNtz/bvepp+58lTpu6bDwRiNT3QpnQ3ef+cW5e9V12F4
r00SbJ+FmH/lkEtxpH5HxkFeu4MANvgaBdtpA8mKacvBJ8p/5PNiStveZlzX+4HQscmOrKK38LU+
k3Ivod6TsoLe2miiTPMGkHEHtTCL1NLID0tHwFkUxRWiwvWbScS6HVWJYL8GbHHHgykD3LUp9qPE
a22SmJMmR/w2g9r+H5o6omR4mOrGCa/75d0qVzdoRoxwBzFmjQWYy6yBHpB36Ft1/WDtM6kOmV+X
3y67MKQHmdRkPiOhF8bqiFny60JNi13D5nfy5D76sIJzCxTtbwHhy2816Iqogibr9xhCBUwjlpOW
snqrcbZbmfP3G2pcZgGx/xcAan/oJpCc+hrfhuZ7scJ5yDrsQdN/EYYS9A423DS3hITACBjL5ykU
+q+UXcitnKCjHypBMgPb90jDi5gqa0yyDEscTpeP0FOx69akAbdTBGgKh9TVFpwAhL34zHfdDDPf
ohTDIrp405OsxecTFCfkGOuz7r3qm9FlvWJI6zQ7wxssqzUJfxg5B5sFMwPwQaGbbdEwF+E9m5VY
pXJLTqSpO0lNBpMWuo43gm7bO1O9N5b0FwWmMax3WzbhbWqVTmZ8uBGAr/ISOb/NH1HcvmsJm8N3
mTRhrWxzqrwtdnnJlUhtgXEFulGeaC5iSIq90qLcyprJ0jDb6nDEMpViZXNKwYwiK2/ECt15MW3p
EfcTAkTL5+GTn6Vwcbgjue3qSJdI+yLAvuwWYSErysXpQn3R/nkPdNzbrWFclIEEEGK9UFLwIFHK
gX3n9XfDRQlwMirmZzhMPXrKUOMsZOVGDZSI9Njto3gkuClIcvx11qvY5ceVqQCeOLM1IeF5RLuP
O+7oxFRLGuL65GxJjxWHvxq2e6Dr+6BR3x7HY6TohCFK7SDiEyuGVfL5QIv+yIrnIftpVpcAzG5A
E1mmv2fxg+QsUNOqy6frfjWSm7EnGW5QCM4YSA5UYLAnkKvOmNaQ7JQHfXJwh6o5bL52XgIh819U
m6cTOrabWiUnOWDC2L7R+o0XOE/MOPOW7YkoZHsMb+UHZaUEpxCJ/qekTpUu/b57CFdb6EsQ19J9
4+lUb1+8gfkp7DeCidfDHrHMvN/tl0q0fhc7tSXjxMSvCApDKvct9UZMLSPEY7sQf9rODAeZ+LIr
kMr82szBuOanKYJrg+ntlZsxQs3pwM9qkdYagDYMcKb1w+3FIuPYYJ015xVtBnZ6g7NxVQO7OXl1
3vMoRXhwk6cXTJ+DaLKjZijsB5TbCSYYMWQTtim+o806vq9A2lfG/sKlE0av5k1WKpevUBDBM1R1
i0N5yJ8Xt91Tfv57RTzbdGNlgiHLM/WCa8+w8uIQhV5sjXvc+YmbB2Oc6ufXI0GbxCioiGa5J2DA
XeVxTLhZ41pQsBUn+s5WvBfBtChpOFa1ZqGEMEIFQdTuGzAYP1tW1J7Sbail6HCpvIXq8Aj8RLl/
7S0Up9kkR/kJblt4+OHdT3Q4c7oZzKYiv0SrmsCL9zhqzpjGClX7YuOrpmt7prtzskuXHjoJMixB
iGeqGHM9CNhueEP0JudgyGkQ9rTfXbTGrCUnxt+m4xX6Tu1BZzf/gVDCvnvisBrN1Xjxl0Z2vsYF
5rdcXABQZDDA1o/HG5xLx1EXdSsJq1Vs28TCv5gH0v4sj7XjKqDrUqtu5R0u7IUQLziWIegveZ9R
mIIN1sYZj5IoqfA1KtGluYgwinOBDUud8TDK7CowBVwFKOcd1gtR/aUwQkvA9FrLLuQbuTKt5Pps
UsECyYR04goT0mBlG5SX6qC8Z5HBhPxErtrMiKaB3tFxLZfj6qyqjq9M1103sWz2a8KiFj1EnhFH
lZvIJYhIevJdNBHKjFwxPZWej7SGpzV7hry7rK9vMQPE6Mr0e7AQlXTyF8AxxHk2WLKH1BXferSO
RPtXeZpbbeDQ1GkFB8TENBfRbtS8dOqWHS35GNUD2naKwqCLmM8aOmQG61+QZpyC4a+DU3EcxGG1
vrk703GsFuXS7TDeNEZBG32Z1TaBc3GQnuuRIWlWOJXgOdhK0EmVETOsd0ARSqSRERAhkAJnAJEr
CJQA031R4su7mQuJRTjZPnGARCWL3OGWQtvNkU3brl0pBO8wmis6kGEnWLqrX9jGkvp5wd/614GH
QHw0+gK+68pnNlQe4xIr1gVictdZfoy7+Phk66jxtQcsTsxNxT3VFd3HBLWZZCL6Nf/yfuEZ+TnT
ftD3rghAHma3lzox1BNk2DA3ljDsPEVPh3Liwpxb89YmOOOVyb1iw2opsK1pWcnBhC14WijGs+Jf
8Oh3/UkUxSWWzNtDNf9snnUl/P53I2croVrd+wytGj++nzQ6VVhEh8gxBk7cSmxmXPSV/EA2mE0c
hDmxMtJmiaYN9Tw0otVl01dDOxkBLbi9+fr8t4BmmtC0sQCRTu/RLqYNwlDD1ihbpUbsNfqmTXNU
D3B2Ednn5Kh8hcK+l9AqDCaA/8AIaEMlt+wb4XZ64eWpZf5KzdmXTzPCqdklIWq3NriALnQPsesI
KcJIGAO988KvvEOtzrasNopYjSGaODXzmdCcbjkeATG41WQWdnminK12H0yYudy2nOxF9Os7lFPC
7RCEJZ+qW14w+Rc+P2l2uz1aABByzu4vBQL6XB9Q6A3JIkvIcz9wMbtq4FqvIClD0iDG+sKX0XhI
bXoxhIaQujWUuZT0pxMsWqERiWwyvcOcfGtrc+mDMwlvNjKPfRgPdhx1LdDh2WLlJp1pDocd2038
pvdAKK6chdJ12OhDDvOjXr0pQO3GFGCMbaAbf6MCVMzUQqg4xT5XyG0y5elnO7eAt83QVKFwv24f
zbt51drXyzI6BGu3D1ekTs8fNa4Uxr9ntTIkLz+WWCtjlmDNqLW37cSH7k/DWm3lyF6uDFo/d5Pm
i/GkCMBAg7fhg+6IDEmPj9vOVdt8C7wzc17hD0G2EwBpEWeGGGhlSyUUEpk4n1oiWYZqyLBB4inm
X1omvmEkmpAA0p1zcXqRkhu9oMmFiU9WOcQo5Sh4HUNcJyI3m5uvg3sj7mivONsfoAYKUrdXPRAt
3SSpXHOomkmvEiZZo+oOwRSU6NIurEyAV7p7nQcdkKT32aVsh8GFdLaqdXE6huKbnoIU7UHn9UVv
2XWWExO3/JyAfTw1tmHP6+RiQD6QsZsNOVmdNesT06Q0weMkj2+F8DsIv4Cle+Q20tWDuphjGX+x
nyPxSycObQS+yD5cSxpZyjnasI4UnhwbHwQtFRM1ciGA/0uFrwvEz1eyEwqaIng2qlDdw5R98NBs
DLNLrsJ9sTVKsys1XqeLA+PknlhIGmmtbPJECedZty4bQQo2PcImjbgsOWECM4se/fWy7LCWY0gP
g29sBkVhN8uB3nyKhyaZXlxLmylaF1yW4HNL+r4uSR5RuwVh68ckhpTiILquFuC6IeR/RzpbUTPM
MHUbHzr68CQ+TWsQt5Q7nTFCljLd2W1Mc7mj6O1hTPSl0AzFM2EYVjGjw42Hu2ysK0Db+RskJVoQ
9hwuQqum6MwvegpZV6MQZfOmHbW/HXr9HLfLa1Ah3peAjgJLXMHjKK2EVaH+A9tdHJAA68jzd8Qw
N4M36A0cU9adrPZKXxxHtGqFv/hVZMWATQe25xazF46SyRtp9f7D5KQF5PYdLyMrslV4ReGwz9VF
dLBkBFPNI90twVzEF8V0NGhAY+cPnHAsdTUEu2HKbBFMFSNKBEv4EYbhUxkFvZUv6CaipyzUFLWZ
8gz99Ai+4zsFUJN7uoVysqXpy4GxBeTbhC5BJe/PWTxPRhmZIJupa25qPnlwAqxtP2Xz9HHElhox
DWZAgbosxTTzXfA9GVWcMv2JsZH5QRdwDnPdsRMjWJu/NpQKFkiHbZihb4MlBKxDP/fuv22K+F3e
5DGbPtKJFIfqPdE/w16f8r70D8OjBvGtXgrBxoWq0Q2VWfnxFwZaMqVQe4tDtVw3S/5v/IHwUpK7
XSj77Kl+SKDc20mB5SrsHdRPo425+/GCpGwEDDRc7uyEqp8bQ3Z+ryK9VaWg/KwNq8P7Gu5oOakx
WOj5mk2a/sSrXlCmb4dqfrRfFHigK5d89q7XY00LMtiOK8EsoiLQpbhH4PjtTSsF6T0tFRREQxg9
D54DbaMqjVKFmg6B7/M/T6jJ8eY5NPUmbN2KVeh1oqczrRtitKA5/HmizfFfSLlDKtymDiNVVM/Q
NKLw0/r9ilrTw4tdIs6E5+sA3wysQk/GbyVhrXwm4iw2RYiOoRz6yc2fEDk1FpURfKzFF7QH7Blg
+1350Ngbed9AmByw3/RwXDy59xMTrLUyS/+cRI6N1SKZ4YHAPHYtoX/NIOMD4FlugMjyCTAtIUuG
Wx+OBgD7WGICn/iEr3R4yYa98cnlmJSuSB3c5YJEyY+fyM5TfbZ3V5Xq97bWbmtP/dSRxT0NpyLN
2HXxJIkeM36pOd471Tizs94Fls3SOzxf/NwEp/8d2ZHHvyZ9hLcAb5smwpUY59mdZ/TzYoXzWwvz
Q5VLbg9EygXpfVPJjl/Expfw8WVmiYM7b7MqtqdyFamYvi6xt+tGidMfp5nn3ML+/BMmRkDI8xW+
MuZW6KUWUzEZz5r5O2oQ4J/yiXV1WZrMt89+dp983fhVZ6Vyaqrk7fgWP1VxG+dlfywJGo8WQDW0
kAqBFyOKwbZpq6SiKtQgr3PLzZg/KavCvjgpzvkmoRjDprFkt0YJ1l74zHAObD0aBoHnlgOKzfh7
9bYQ9To/wyz7aboUIj4W1inukBBeCZOjMCvH8NcQA5P3tUwvl0DejORLB0gpHG43mRHaBO3MQtQv
qAvzlhghEiF/mBwOpzCrOmsLJCkzWiAU/FJDkyvt6JFbXlAwwxmxqQLG1ul9oW1QO8vt6fOPhIxn
YGkVkAANJFEOSAh/mcNvNu/tWy1VosMkO5oug/pltTS5EHUVYFNUzOxyikMYF/cnFqmZ54IJNF9y
ab1qoM/YlirDlNeO6AIFwa2D2Wx0fh3jJmIsIKBGatdTS6o0Hy4CFe59M2rP2kWTTTkeamd5B4kB
WWRQ5bU938ipiLG8FgyKWTeVmYyWU1LUn5jSlWrw0mky7otnt+jd75IQiTe9XPf9R6ok1UYdqxhK
6wF/UAaIQuemG2YnLMsCHDzo86UHlc4HPPs6Nfx4j2bk1F2U+uoUdtivIhUj6C0Jyalm7YiC1qVa
8JC/LY7/ZF8CgLTQWLbLgCFQ2FCsh1qLJM+kLMX5zya6oEfsiCh5xEgYm49EOzyfi4O73hyFFV56
U8fkhuVYNeOnBpEqpAagU1YxQzm6vQfky6q5UoSeC85jt6Dan4afBeLmLGFBv1kAcPQj0w9LRhQ1
dLpaJbH2zwDQPhVXW3vcvkLx2Omz1ZBPz9LkncJ9ZkkrgVPb/iq67j3IQasqpyIl0eovx1NzPDWG
961vVrQKCxUZEW2gmIFxUfPF78oXtVzKCsAr3jKQ4H6ru111nO2TMwtSXBa9mYo8EJae3y0ORJzl
koukNqVaIu1wOGU9XfFJacAgZGFROxoLJTttTBJFopu7Pj+6pJaNzMMrO3LMjleYJUxc2uu4cqyI
aIfS1jRWaA+vCGqZ6wscLP7PxHf+zNqHZFCp/QW9YdgwpvSpdMKLu2zE3AD9Fnn3N9ah70J0El4N
D4FV27BABOFWOLIWZOiqW04FojJR0YM1IItrk/aEvZASnSYgbkB9z+oncBJJ2k89JMDKIuIT9XBU
XBmuxnCXUz9pvQEQGL7frHA2Ut+7iPoT2TCtvkuh0eU4QHsU4h+L44Vpet7TKSpkrt3Uoj4aMA4d
16TdeQ7NLOSm8Qw8FszKq2zemQRRqPCFkxV1CZAfkxiNujaXRp3ZODiVR5UOZOEEfSQ5mK9HxEso
ve/I4YRGaW8ZIu3yfHKvuCTjvXgS+CAPh2eFXf+hNMC5kIu+pO8j9eOM/b4jt9lPQd4rvb9qblsj
MXluHh8yz+MC+J4gaklSDqD5xd4SgTp56Ug4FbkWFLFQq2YNavpRXQNDrtRub77MIa//BDgoXavO
GUIRO/zcK2wKIlMOqQw3wU4QQgK3/wmCTvTkd88zKHj9y0epagMaKj6hrtsl65IqXppKtvct1RVS
5e/4B7U6IGxe/IIzj3i89yEowo2g9V94fhvTUbTX2dn4rDyd1BA61ZkkjiEhDDGlpylRqC93phWt
3Cra4zk7A/RbkSp4x3G+XfikPd1abGhEjOTz6ghpQpzKVcTn+uOdVMxstQ8Dh/xlTNKJl2x67SII
QbVJzYZ2hLLb1aULk8ksk5F7fhxBMFy8I29zSgrwuNeR2strbf8dODDzYNrtzBUb/bkTUlGbNVB2
fMwyyz7UWvfp9S/HxtLvnAU/Du0FA/vXMUXHLVzk296c0nO+Cg+2s3JOudvuYm4hrhnSbk0mrrl/
ixfzxSSoXbxYC9HReBpYB9wAI45K7A4ta6pag9Z0JOyUyaNm7zsaoz1VnNQmEi1KicSSIjyQ6Niq
WrkiTbZFZqNknh8RWUL1aI/dP+mmUSvE7+OozV/Nn/qUC22Q1CAqX0myzlE0EHtp7EYhzV6mX9q7
qOp/0J2y5LgJlbxoDFdDzjIhAKT5/7kKE5IO5Ev0YzV548pWJO9YZGrNQ34IDDSZk9uNgt3D2d1u
TqFp8QUi+7oxwGmLTd0tHghPYLbB6x4kfBWnODExSGPw2evnBuz2ZCFaIa3MAiIqSNuR6yqhvXSj
GmdMR2Eup2+Bn72bb3oy0r/TFKg5MnbmJ97nHma/mDTeoegZ7wXdvw2Nv/65u9gayt8fs/49ojcL
lciSy+FqbsQ9hPayvLyn9DtjbAdIeFiFzpe6IfpwuiOfOyOFHQuabYWvQeDFfadNEPTCaCLBgm0s
bdi8w1q82UvuRT+fSb2jh6upkhEI57B6bxeu/kqO7R8O1CZnbE5VaneoEsFigvQ4oxe/6WNnTbMa
fvGqJqkyhV4rvSgU3y7DrVJg/zrd3sV+yhVoslkb5ZXRmk9i4RZb7PIOIIuwnqtATUWpBiYp3hOR
Trk/UngWvnnD7Y6XSjy0a8qbV+PaMU1mTC2Kys3e+Kvs7aw71kE1P7U7oKuBh1v9qOVGZXMieDCt
8OmV4MTgCBiQDPIq4R3YjJxtXOpKuDQ4MjAd5pEZDDihXbBul5IhDRUQdAuaX9RcbVW3dtdRs9JL
U0AUbjYL+wOwarkLF9MN5SBmeaGxqqRGgePnWY1I3XjEJPMYq/glQgSgMBzoJuQ5G/5UrZBZb+vV
ef25cWzFpS0sKRhgj9zvP27G5MNuCg3gd108xce3zN0yoEQY9kXX8nes/xIEsyMLZ0qImp5kiqyK
08rAQ/2DRcZGDjudj9aGLvYE1EIa+csDPzAwq4RN4m8ovyc46vkWIT255edyIyM9mfOBeV5NbG3T
L2TsO2yroupkUHqHMx1AUXA7xy9dr1augUTdKMJ+yFIxmtcCpXLgPtBQepXkLbSrbZKp1g2C4oWt
Jc+gIU8tBnfSTnbPbQOdprTGo+wF4RT8dwN1ExAIXoEdwigrm5UPEoMeG4MPxOtd4a2iLF6nabXZ
AfmPTuqBYNbUMvduwKTH2AHpp/SXTaW88O1wZcz54M6+qEBTcW3yk1NZP/6UzqYWBNJ5kS+gR8Tx
H8zgtwql0Xte5ZJH+JVr+q3fXBG1AbBTVIyzyWNa9AD7UF/vknEtWHlQF7RhjoId+2xOMT3+jwu1
TgEOGgiym2TfIzmWJgvdpa+QlT6JNMe7dgCeCqRupq6NgyAfpYikVbJLpuxIA3LytumRA7uvgmo/
hPM1WU13clrrgkcZjq6zDojS9AllPA6PNhy4AxKn+G9p6RNeKSQJmF+itwUUo1RogInrAvdALzsP
Vj7vrZYexjf/k7U7ufM0/5oP9ouoWnn4xDzx3ZXpFXbQwZIC0KH268p++aMdjrBUa53ot8UWiXZo
IYz2pdjWT2Bg94uWCtzONyUZibS5sU0ZHAOld38J6fy3Qo7NXfOb+4B3r0CzvTmjzE9EwhMrb7g3
e/UT1IK2b/mEUwpeAr/za7sYvjEeA1amjyJwZvB/MptF+QTtahJR5HjZxXtoGbvVEFcEGkDb/tBH
uUJjdPP4dmppxsrwdKrO1PwnjwY8gfSUpYoIz7BsA7sSfj2oWGhxgUfCRstPH2gUx7UXsgsbInTl
N4m2rV2DyevbLdyswmqu4gvJZxAV/LX8uTAdQPPgn2GVszKg10PMpWAOqrNDcKqFG7P2kt7h3X0f
Q9s1eBrDiwwMMqPG49krnupg3/7+7TfkEwoC4jxpak6BAegPtBptsYjxcFp5VZkQkknwkpZA0Akb
4aIL/eAZrBJeJ75AdS1KHU1RbZvX/kVHDSEebMrLA5BXFzbWXAF/stVkBrFgusvj6In4aCghdgzy
deC1oiX9f3NzusZK8giJYJ/gILuPOhXzR86MoWTo2z3oy6iuPYd0joJIViQ6ALqYeLcQ1TMjT6BT
lTlctV3HoiD9jQhOhaMlCfrufthY6ts+UU/wnDI6IPm1BPVJV99RF0697YFjvhFEa1i4DpMcP6g5
swenze9uFQT0mRh+wP6to/m3vqOeT5xf9QC3I9APUnCBUMoYEaJE/OV9Snu0z4/dTGr0gvFQR3zQ
7eVJm1Fu14Q4FBAgdE/mC/CtgHg3l3u8Lb5s9FiMjSeajFfHeO8iL9IV+NU9wlrIRaN3n+cnvVAk
eCsIiP+aM7G7iB3Nl9M5TiNuMckgUVrLdmYrhb7fsedF80iWsxxDsMzOgp6GsxPWrKZPHVixV6Se
Ha7JJlL2VjY75+macLZnMNFW1KOWTza7uxWbkbuMZ/PJ602eUkNHWFgCPGOMVFfQdHcBiYxG2mxD
QifPz9MGSrILxQJSWy3jvm+hpdJxnMhBnOhQLUX9+GZGVjSteFpXSf1v4hrsx4X3pN/ov+sHxKaB
zZbAtLS96tHSXMohADGqLWBqGUDxfIjZKAnEK2lwRia2W5WCespzpC7uePmEV1+QDK7yzO6fO8Gd
6RkZvsEqKiHL8JwtGRSnYLhcd7lrXOKs9oA7pIQPLbadw85s4vmYBNri5SAEtFYGO/7C5h+z6vax
PQrAZeSQ6Z7VPOmTgu5/tXw4vp7iQUuCDOEZvSdnou4jbAhfHfBxU4+j8OWqsZYL1EOzGqhpkUda
15l7g9vQiAOwUn+8xdFkrcGX6fmhg6cHeos8/kh0q0G6tDJHtBWjFLI2M6iRTD7LV9c2eL6uFEGJ
lC8je3K2NnGE2em2VqwYx3ymP+sZMGtqB+lavK2D6OtUU4KegPVxYhnoxZ7tUZ5dvQl8FH2Chl8P
J+xmabn9sLbTmuk3AmING9+ckXuNH4eQOECeCCmGdTilVaJ7EjnhqQfZD3iLiAdAZm273/KFud74
Hppax8NlT+TJl1zOcscaxKCw7Z0yKe540HdZKmUoTm6TodAa5nYpccjDptKMxP3weW5q0J+rou/C
aFGJPx/jqSSTceGWtxK2mVffNIwsST67Y/PeljbxntaahGID5wGj+pn5gUshX+E1e+8x+yIKaT51
AqMVoj7KG66JmET/OS4mZnrGrdJjxviNprWqKVMDRsQcJG2xrd6pwgK5vT+D1SWQdOTduAVZi1sh
EUK0zYKIx5nd1UoaGp/RLwp6CkTHtiR3vnYzSjmc8x5CiJt2ku9rttN3vDobgd3UZTrHz0qy201y
nJK/TrTauzyHWkihl17rmu8Ob//SFrKS1htD9KSiUYVg/9bfEe/TC7zxvAndGixN1aE7VE8R5oyT
f3Gk/VSbZeGIg1Wet7sg3eZ0t9S3Gl+0+FiVc5Fhqrzm7J+JE7WUaNGMaz3YmcLetrLVm7hPJbV9
UN1VkCzrKLaO0Yik9r0rE9tXlJKh9rVB4ArWydxRpcZLqQMCt13IeC6IvVFJtIJNkbZcsDghyNR+
585z8Cv0MRNAYpbESjWM1/PXGRHrMFwUfCxCBQrRnBTZZT3iUGm2lQAgH0Ef/n6/DIj+V1NohwkP
vv5zhPBDPsYeR7gUrstKn5gimqHS7UYpNoX8leo2ekchQI2EdeK8OFI5ykKK5PVcdURlJgTnUz11
vufoHQN2zO4hritBaXSBrOOEx/A2ult1joKLzOmSq558Mq49xnAS4t2xbSNWMgnp6ulvgJK/2+X4
Mikv3u16lexFYeBJbIJ5B09m5RtxP/YADbq1xzmcczg86CvDDVr5pZ5lMvUea2UrAtOXcHm4vjuv
mEkOtHTjWyEqai3RNNodIZjZBFQ6VFrIk2MgXmcwR71GAX6bGZveVvRTwhlMYfabPKOErmMZiGAD
qKYXciAZa9uniCMX1uHWd/H7FDQWsrmmHJlSUkU/HtgCaA8/+kb3WyADX8H1EtH1JRLdC/X06wEK
SypRr602qlPyHvjVZxXLqwEnrxILPfdxvD2bRLqb79PPVFftguf0DRdloSnY6gz8HVhvFg3hflVD
eoyNyxgHyJoXaQG92n7jFEPd97oIvQy99bmLiSgjQN+fNkJSty5IxRHpdcWKc127x+C69HS9D5QV
eROVBUb5EUF0VlUo3imnAxgE8QFmAxiZIbr3cn9cl6J95xkz33BcadOKZhwyUIxNoXVCglJAT8sS
XDD0hhQmbXSrqVF/lFsDFAdHWVJEQTR9Bu75UmMBkL+ThIDDhdavZhuYBHlS/NPs5NsiWVvk0LGw
0Hs2ybjVKB8UlRGgpuJ+pPqQa4IlOgQYfgKlHZ+9Ipdlt4vzXcCpnXDwo8sydwk4Jko3koFAAOJl
XlDqtCIKvw+9rEuaD/MR/BpuGwSs9zD1Nu6GENEqIHu4/5G4G8j2FSY9+Ks3KZUzk9ha2c0RHhnx
0x6OzKyyBBdOiAa3QxxVcx9btOhmqSQztfJu814inbQKY+C2CFJPK0lBcHQWTQIiu65kh61R5GBY
ETZqZS9O/iqQSjPaxLqcs+mQpF/k4UlznWfHXKyUlT/jHGyrzdaQ4vQKs3cCKwj1v5/8985+tyNS
RowAyiAlmWRnJ44uW2+oCOWl1kGthPd5m+vQGcpSNqyZV8Wj4nxSYKxpvbW6PfpBxAjZlzazA4QA
BZwntxhUqeoI9ck3197zIITtBU4NqqaX1leX8qOQ2tWc4l3zFO+66AS22q3POpKC0apJtiis5wUV
Lu2pizP77R+f9n3dk64/ulaqeQd+xJLnf/yIHn5ikBKKR2Go+PkZz8lUB0U8DzT2KyuSAzjLDFD5
NeHZHR4rUWJw5SQHb7HpvpDWlLR/JXcS2FsKMt6jXLX2gDo7TxOr6h/98wxh8FEV4e2uDowTnn/i
/26eDc7wy8/tVUiAyCd/2cH76bsb8OH+GCV/hcDRQGwvs4/f4pFPZTCYF5rGsYIR4UzcpNU0Guxb
kS2e89zJQIi7hzXi2r8LVFARkAcb/b8Xg4/G+nqYGdL9eVDlB6YcUsUTrOIubWq4fQFPD3sECfzX
JEuIZkNn2Nzm4LJAWXdPYFSEmCGJe86kvM6HdRrCeKvGeaszoO+URXXU/QmiHTdNUEaBjSnk7Zqt
4bOEh03T4AFOsWLfGAlWDuyUB1JJ0mQ3kjI+xH4Ge40HiR/+oVnZPtBoq75syD7iM+dhNMq9M7LV
X9FGc52wBqfUvSIC5gei9htyk6D6Azmn5U6JCXVzWeJKxg/k4CljgzLwJt53I2lV4a5NtKK2QdNH
9S++OrNbScqyUqxjMG9uUsUlUSdRUUjvYwh7suH82MSrmJ7RgHGFbphnpuD0WPD0pppqVrGUefBK
7BMVVqJ7V/uLCigMftkQ0NsJH83X/zl9L+VX9TVHeKJmDBTs+63XACGJHk4KaSRbxHS1ONEu0ulK
2aZpmNb7QMvQYAyj29hOcxmqQfOHDT1ILIcT05aS8lb8mTXFsrBKFKoi6MtYs0PdcHUuMZL0cMjl
w+NbfCecm2bgCYnn/IcE1kP1hjhEbr0dy/QjlKxc2A6kec7CxBWtJLkTiYIcdIDzF8Wdo6LKwFqp
TAA6V/L7OlsG6H7WiFWsD5GdJWPabC+3Rt1PoH9wyl63Uw/YJPnUm9g9AzDUygmUa0LTRlRgfXEc
Jf0J0VEcHmIKlP3/gN8w5XuSR1TpgLWktxiW3V7t7T8r6I5LaT/7Ji86wJVn5BROymoS0/885C/P
14h1ZVCQub8evPEa2yTnA0qC7yQSf0O7hbMER46eRi1xmhZfmWtAAcQqsoiGirUd59CPYqUvveNL
pKPBh+1lQ61ka3bS0AJoXQUsysNWA1AWcEFyz0svhmyh56PvcLdHU6QUPm7ZpptXZSooPmEQBfF3
/PWIU0UxcB4NmaaPvDCmDRLzyep5ZzgTAmVDqezRDwUzOHvDpq+0jXinuHlKzWSa+pRobCLfKth/
0Cco1rXKqLlMKZK1FMmeOA0q+lHQ29XjB169nSeYle9n6itVRe8+ZpKwVtuTaPZYyqTCsH6F022j
P9HGlQCNm1vM68n+v2Y+qHlZVEX2SxqfMqSI32f/0ab2ShW5A/8QCDBovHYpckTXkzkhweX3Ccwj
GS/Z2ZsFKyVX4H4Rm6NZZ8oaOVMXTFDQakwuRJhQGOYklwNY6TFsFAKJNaG+G09jdT5mLE3Pj8PT
cnPbPvU9lkE8/P5s8m8MH7vcREeBEnMNpXLYcOxtG8wxJr/KOdZey+/9QW+430LHMIazhupDU8zF
BPpjZVwVoJSZG28KTgpS8olo7Ts+rfenoDKYSwq0kz9QV6rHwTJCvGYwD4O6CHhtVSLlKetKwm5w
+ioMmrGHE4Lj5HiTjqfaH0erEENW4vJGaqqa0WrEDnvcIOit3YJvvbpq9lk7VJadOJG4n8zxWmgP
iniONXYjIrgEFkTerFWDrOvPmnh07cY/DBbr+PQLmH7TeojCxOqFG8ImHdNhJ5ivnp9XIYFeYwvR
GDqVbmN5cEXe229IBDHt/eesWrgJ2xDiEqlTpCIuPfmqsi4xoXY8qdvxirIEF9YTJb6236LU47GE
Fjh1+TvLBIG6dalUQilNSfkMJMxNypmpJy/wigxE83k7UHNTS19MqJi3F/OvHEtjt89JvIi0hPXK
2SKYfgBhtGKtYv9W2HpB9n0mFAf/M7T0JxI6liK0Zcu5zWONWBUIpf82c/5yqx0xrz4pLoaFICx4
gRRCetjotGBt03XmAM0lrNRyepm+dnuFBnwyI7vG6HHJ4L32ZlUVNLAMtUwhjdiJjX78rGVG1o3l
TDEDEABn+5vG4oEIghDyHuktphrEoaxNkh8TWITOU2F50b+F3iZYJ8RAKL+2XYv7MFFxybaBvTGN
8Rx8azp+j4p3XOTIbzw2Eml/KQx1z96oXmMh0Zdx2HQYEjNI2JomCbVpp9Rxfi4jjUaluRhvbuXU
jG7d3CXLycSRmWdzUGdVCp7UKOV3jUP818uTDfkHgFynxGgn311roPApIEGq4xkMZqqSBiPLPJrE
uLtWASvK0SONheIQzgTG6yhSj//vw2qe0shsCm7VB0HQZ2q7e+asbTfoZt2R6RSLOu/DcP7OBK0v
tZwztCovrtehmtSYS/loBsCSrV/nHk5kX7QrwSl81W5lzEwy71YFd4mDVqb1BXaWgkydQxjH9gus
40v3Gl3LQEeBLTlzzCODiOHaszxpZvmPCYXnWTxXuw9TQcq8TAIYK4KhpkW9o9TgrJLYZ9hik6VS
dGV9rHSQ0NR293r1DF9caTPr5bQMzNIw4aSbFUUdcmKY5c4a6jDftc+RCYCXUWR8SZw4h5b6kHHA
mwE/Lk6ERZBis/cOTomatfsGtDMMvAuen/fF2NUmnXD4QPev+pgrCkTmtlv8HnIdtkgydSSfOkQT
NADJC8fcSn87LbAJ/2vmP0hA6KjxRLK6Pp8VraBliJVKg4vdM+W43Vhhq5rPM3NYIyS+JfH5zPMi
b8YD4slyJGvzTRM497HCSoL3gZbc6RrKasL7iNxyfTcRk2IUOktfS78Mt6QdQCzivQ6lA+rPBZdA
2Lu9IpNE2eD/vsgQ83+kJdrDXvIulFdwEtoCir0ArA9hp1KFKw8re37DwjJA1PYmRt/YBZCqaSDU
h8ACThCP0pCZIj7dN6cxAeoiNxFFOC7bUE2S4E3p3CNwV4r7NpI+GWesbpfkK9caDvyRGea+Toxg
nfuurjxLEBriLN+zkA5tx+VTempQY5MXST5Dy88cimS8NUg1Ni/72wMb+d6JAM3vQP7BoPAwy4r4
WdleUF8WdUxYbmou4I3ydYVycTF3cpnaqtIpmFJZhHmBKEQ9fAHUvJNlZa3AVlqo7Rep14Y+n/w7
Gcs/B1FVA8K1qZHej9BknS+JeqB7f9+i7oL6nYcO+gCfaYPncwyXU2NWA32wzCG9r5A8ODTtD5yL
7uIBlLoUAqb+XKxJJkpWAGBSQYC6Ldhmm5PzH5u2Hth/HkxdlMjhGLhLADp9awhIs8FGxZiAvbrq
luBsjjeI6X/MeIs6ANk9AI5Ge2Bn9udfIiH46y2zgJ3goMhlMaJk8xkaTUDnv86zo37k3wiJdp+a
9aa0yC1Zgb8beLF4rJ9EaP7QZAl2JEMbHT3oaXJK+aD82ZdiPApu9/Sye798ruyHrug/aegXyitF
9PuGV/rIGep2j5NDT9zrH3BwptEgaAK1wDrOXPySoYP0VgSuQyGc2wOhsPkziR6Pjfno5RZtv5b/
SAvYKcK4Xwz8V9aVKawALFypyolR+MrJiB1nUzj3TjyCD8QGD0//z6y/rJw40ANdGiQaJgFaSN/v
2fN7g0vQUwsAxfhha1fGbe4SZ0CRLayTXI3Uc9TjJ23i6BIdSsR2EvLv41IiNdgR+om1FAXOpLHp
EXaFyPFlwvQoQi/FXTsYATFJMoKvtxIZB19dOz4MYLfRw5HMOLXCSSSshM7Zf8NYgTRYsIVvjdPz
c8F8O4dadED/6CWohEn2TzkTiyIcfeohr17pC1GlLvB+AV8P4Ri2PHA4LVUdvzXeJ4GWnzEGFgzq
6TqOOu9Gt5zR7nOKHzWOozxSJiLHrF2Ejh1/mlaVqZ40M8X+Nv18L3f5ETUJGZqDUuSPp8NNXKNV
JYWFwmKA+k6lah6wo8BH5loDyx7cuJkK55fomN4NuMKpjQKftThbPP/muZJ06hvw/1Z1y2CmO98H
flVtBEAnFU+55t+h4HJixYngxdC8P228qyAUti37qSRA3zfFXzHCSlKtL3FCg2VaNGj8YZPFp1KA
HLGUjm9miG7t7FVwQ4Iox7I8qrIiuG810KT3mpvU4A4pyitIajbNSxTliOyY487XRGsQxR/+5qSg
Anu5qbvj3rMPtzUOPy+V5Kuc3dbapy+Kl5IdPXrTOr4nD0wUw3JgVaSmh9lHgJZviAn8GUZYzOoc
jdRXNbnQvHyOW0Zn+KtEu6bmD1qRaYOJlqZN8EkN3wiAyHohrY/WsuA7gUThiImgVJnk95VRO4uv
F9byYDGcRFEIBlPiDkPNLqEH/C9AOttbZgFIIIEGzDkD3k4DxsmWLQUXIcm00OgdJvAZDUzUxbDQ
JSogp/AUF7zBF5ZWy1AQKDUR2lbvsJbNQhWqVWOoJ4XGxHsi+B31g7Ku6C8HwQZLkvlUdr/HQ2fe
G+s/pC9wvKcnGZ8AY8/q9gcJtqykVKZ7KFbjL+ZV7TjLfy4iRFJ3FwX8mQhEAo/JLxdsUB6jdSjU
npfVZczlYlbOSAyCHzd2TyoTM82+EKMZlm8cbAm5k/gVNyDL9QAwPaqDfCtnKcesdomLdGbS/FXw
R/oyk2RIacoxN49Uoed5LCH+ZAAkFvyOz5lfGhm+zQ/sA1wYOf6FiqtGOUVmiIJ7UULzxV/SPllx
utKo1u9TRmxo/wWbjDQxT3mhxsc7KbOARuyhhHxLIRU4pG6YTNA+rvhKD+zay+WfvzcW0Kx9ZdGN
GbwX5gSd2f4bfDmsWRn1oFHSYTU1GBfbXoyNhfwjry7697r30N7T3h8ex4bHENoAdDgI3JqNihH1
TDyPhe+fsIj2iZqpQGRZKeM+7NqizpsiYsc/oRMGYvD4+qVLACidJBRvsxz9sezJbVRqOd/EgArq
7rBnYgsOPkEQ1DxIOOuwbKrMFhcuzvrVD0mCCvbrRVADGtuy4B+pY0MRSjy4z9X5evGWILxVgsVD
PTp76K/jZ6BwA8WLNs9QI/uHuvweKYNbUdQfUA8kYAPsL1rnJGxiU2YLcdg8YpBERUB4cYjberTR
m48/j94PEsa10Gaf8cgFMBjo+q15NNbnDL7n0gNSzTp6Qt4HeG1zIfkBVvZtsL5c6NUdpJ4gjHU6
Rwsi/SmZJyEnO0pLjTxEWUSk+zJSJoj7WFtKXmkGjqtWw/kgvX4pmxdWtdmf6OPPbObmCXIzdugG
xUxBb5KfmkAMAlHdJNxVNJXJA6QTR+lh0EEroeKEnc8yCW8gEdMN1ExHAK5uP1NO4anTp3a/annA
ihLpwszsorolJ6BlIC/nKV7ZVL5sXYtJoR2FbaWkvmk0X2QjtRuwLTzd9X4tOsNAaND7e88vGHiK
cyJXOwYFeaQIZCK/9TgLAkiakEA1Zk2YMI0BtXOympOc4IwpHvJO65/4w8GT39HV1rqKXMR7Lta4
7aujEAaKh8G/LVn1GZfs1Yc6xgt6w9rqql5J/AmcS2kvLswWYGDvTHj9g6pkyk224O87HxZ+vL7H
r5dd/cXmEyoGGmOzB5YhfOs0zrq6yGZsa654yvWCseh8HmjU+DepABpqW/kfyxoBreY/SifDj2EK
DCeUR+Np06rVH0O6SndO5sodoD1jYS4OHF+YbWM0sj+wmqYwm5alIXUpsyI4GXctj/D3zXTNBpyY
tH4LUoXS2oVEBnXMMBh/fhCCSylits6L8qIU2+zTWRoD0FNI73SEqwWvfxVTK/Du9CA2kVjTNY3V
MCL1orW7GIM6+pXHCJAKxYuvj0+Ng/WdtAMLf6ueADcujO6AliDVxoz5deXxqKTVgha5zNj8EzrZ
NlbCI8gcsbgdJfqhAYaBK5zQ3RALswA0gM1t25PPuqxurmXUrSvvcZ3qnT2px+aDc1tMdn6Q/cuU
yMdCcW/GBFoGmUBZAMTpFCfrqZe1GTeKh5jTJsa0Eny4vY5iNGEcPstSskrhQsHUBjyCsqQ7/r8v
eErzjNCqqruP6GpLrEyEd7ibfbefALmx2Y8/Bb5v3Gn6xNjUJMupeYxBUGiMOLALdyB4ZqeBf2C/
Zm0O69i7qoDE7xQa+5zOW9gu7jTLsFJggwUCoLfreKlKJ6vM9kVnlm7S58U3/VZcCk27AlJyfUsB
G8DC/KuLj/F8+TfnKrCgSzgsG2lRysN9OTj7gJYm/ruGXTCYyxMWLlB4gupCLLKqWmPxKSr1TByS
xivXdagTjgZuHZcxd2Ut9HnzTkLHhW9UNM65qAWiegOBnzpiu+UXeL3S2+49F8NG0tMeLtuyMGgg
8j5xIItKXMw1k34g50kToduNMsDyG+dvcX8k6miU63SqTC+5ri5APxdYiMXiSzR9pqlTVCUtlLTp
ApvIXVBUhNyJavBaL5YKmHq+d7C9Dhi7NZlQNxE2HIZ8wJzttAbNO087QMgeM2moA3Hrou+Uuagp
Ouuoc5zgU6a4cGChJ/WXx7Lcq9ePvE8NkQkbUlfvr0+XW7qomVbMfTrWWDqBSSebAwCTok8YiOq0
NStdwrqZp4cJxIyJhRyCf7kDCMwZEWsn6DIRNl6S2lzQ0qXn9phktDEGqXVG9b4p1FDahEfFYpIg
igN4p9DnSd1HHdsPNuQFSabTkoAsnkgrLFMAb1w5DweEmpVYd1Ydsdr+GDxrxICKh0SsH2iDTaQi
uaZmJrOdsK6uKsaOSDp1syEaTZIIQrbBw+NpcLxNAqHE8vCOLadU5/jBLVvamRU7umxHKBN4W9Kw
oyADck4+9kYXvWH7l3dwupVaMRjToTVj+6Ti78WE4OUi+bnd+6Jf/BVX+ZXh8sJnj+l1P446fpSe
lNnAlNK2PKrSXRds5AWvModjwdFjrBVp7tnpS0CO3eQYa733yYmMYhG0+hLRERrIDg5l1GxUBPrX
yOYGRtwz8pvRHlSrYd+xaPoHmDmMowAeqiM/2llWEOLPDv8m1TxOQgnnsrSKClrwaWJCgthfjil1
/1cZEOH6iyWapEefFzDTCq51CqUOYScmdnc5Wr/eLXtSMPDaJsB4OGwGc3TgOiyl8P4y1xdxeezF
l9TRWsVNI2xh8pnTj/FmfP5fXKosUlhsK3vp1VjMjTWv7hhHo9fP7arsnSGYa0mt4o75hda4Ze4W
iRuHXgYnbrKQmYldVNFcSW0WPHSVqSsfkjahfE2k1NgEqzlNM+GZk1QKhnevYOXd1oi9o2c1nahd
i+BNhGC5z0sp3xUwwJsDgBLV9apIWudshVVzvZ11kkjj4nDiih5xj8wH9J4T5kPn3Ls/JYCAt4K/
q4w4RS9TGDv9e5fDmjfXYhrnjvptHfBbflpMwjQVwkexmGFPr0U5DX7Z6/Jlg21J0Gey8WHIGzMR
MoygO8Tmt9pNSimHX6Bz6kXMIwiYegg0Vsl3Monp7e7arVQZmGRbQSOvMji/zgCM4vQxeIXm3OfT
7MVr+izEcGCBsmAX8ZFxxTSPNMx5e96vymbyx0SzhcnGMiGNbwrrXf0sMhdZ0Oron3iJmjXJ7npI
j7dxPolGMr7ScUljxqJeiu5z8gs5x+V9wh5zS9vgdokf0Rvq+x5Yw6wr7ffnvF+E2H5wgB9784Jb
jgXPeM3xb+wTC/w/HfhjZl0+wpzMyg4EHXfnjn2UAlUc4k3/BIOIz82UpPOqxyHzRqzxsJ98Nqty
XBxQlfMBnzPzJSRokW1wt9aXJe7Zo+3rmlMdyw7Tzjjd4NsMWEMRg//L93W0eACQGM30JmHh/g3w
g3DtSD2w1IFsjPWHfuinLGEneBdl7jjqV13Mzgi5/GH/jxhcgseHFJN+hHLp7aDYIQ6g+Zc3+JfD
u2U9alrLWxW0E6JKQt8clfeGZUT2No2S2XWRt6MoJJby4dcitUL9bJeHFvx2txQJve0zhyDLVCap
OWupBxp7dHmCtcc+oJDIE6mUEhcLRzV9Zp9esT09Em28GjjJKHIDpXagVADAI4iXimzhaZTjht6N
QQ0p6ftZTWErG+AhyJxlzaFMCNb8W2MARWYA1Lxs8+zfXueISHImRAsh1sPHrag3zqvVj/9bmcSi
t9pgIWy2Yvgi7yEtJkYLxCBAEIXiJmuqWBqfmN04lLhD95IhmLdvrijaR0/Do8A+/6zQoGrgnnS6
z5/7AdHCNEIFE3sDyQhrcZNrZCg94y08jmU1vo+J/vdbnYWPBnOcm8ZF6d4bsZ73whxyz4oquJSw
hb0PRL1eiCY47xJ6dNIbq6qzI4zmaNblYOm/RzczqRMWz8QjzdvE1kuVB8gifYPT4Pvm3pBnAorw
oA3jID/AU9RxJaIyGPc7xgL2uGCvRkxYewiuTfhsfdKPIfJeYG73cDtMrj/022FetCzE7q0lDLaf
1UNBmBXXSgwrn6bC8anLqdIAMdeQ78Hg2InpPLV20HJ/LLc7B1QWh6sykuq7ATdfa15miIEZgrd7
K/ThNMGeE9Gx9Zvi9vaunGYNYKa75RLAdnuTxEpLsH8P4oTOXNhyfZcYxojygeviT5UfwowOcVqs
B/OVriiGVlra7pPESFtt/TEz8/sXJXG6Xyys+Zdzq2Jl0z1la1gjTjrJLYVGsyIz8MO0/mKy5q0Y
5GkPzTmmwGkkoHFufrB26FyBSZCzDP+je+8x4Tv94WapSZ7FiRE4bQy3azCywV3i4nNCTx6j8W0r
Ddw8jv0npybHDCwRkASf4RBWiIXbkwZR6BsjbN9aKBD3fLuSV/dLGteCIS/UxJh0+a8SSgx02Aq2
PmR6ELh165orVb++zvBoBrjkGutjXh78SqYIww3xdYjiUcgmp0E46NdLImKpB7a10D8/8snpZiT3
hCUa9gzTDI+zGA/iMnlnX7NlmKxUbTdPjukLxOMdiknnW59fq1Iwf4Xx/lhPYZBMfE8Er6+jfrN/
/GGi6COo9AAgcoc7lDV5us7T2v1BnvnUyJvqYgzAeuDFGhQFqbSU5qOj1D+i/MohfRNPd4wwjY7H
VEH4YwYjD3LfuAFFkPFcr8oKAxxCl8axoeUzWL8Zn3ltHxKFUICQEQjicZcAfnNtNELXqlEUsCp7
rXHp0fnrBlPHPAagVkHT5FohfhNaPSQtuB4E+H8EKq1iUJlZy1SBgKV+2EHInpss1BOHfIHOcXAB
MNyhgcj59Y9Hy7b49T21xYwndn2slcgoTBMJnBGtoxZBSIbcsZfxoLRydM0o8fGYx2k5VwVFLzim
O6IL9HlKmabYvUQXH3XEV7RD2J9ou/aMFcTn1scMpT7yxiKS38N7x5toQk1FB+fU0OA+d4ikH/AF
+sboXbK2jLya8prAQIzMxsW+uvrXoDuaPr2kEmQVB0zTY+YoP+5xG13pxQCrUFzOj6aqxh9JT96C
ihJ+xlRFGmpZNH74Ze5OlRPtbO2j4mK/9aOxPMrnAr3F9SzLqRJrrcS4ngRGMjfNu+0PwmiCTUUm
LgVPmIpDfjUEP/UlDf9jS9Dqn8xmpzHglQ+fl53nn+bZgZmpVW/naEuVb+LqIq/CzmDH5FZB5ksG
SAJSQcpUXFtmE4y6hX4UljMCscswejOKEvhtyqwBwcT+4ax5HQqbGpjzGSpRlu2HAyhlzaUcX5Qi
zUbCr+BLhunmxk4PUsQCI6qeROsx4DbR8jaMiLO9MH+wT+v/DL4/CSPWZZ4xDKGWP0HqaWFSW8gi
d+dv5jpOlZdt4mpa/qEgEfWc5nKgVoBMjjV2QNxevLLMkrSZKOMr0c0z6YmIB997DQ1/9ejwD28q
LkPUfOQla2s3XInxaRD+dpfu54pIhbF1gmLPzBn8zx1RXFWF3VIjiI+C4tH1oIZu6l+kqJ4nQfT8
g/hyeuX1xn1xz3hDnx9wC1vrJv0YbUfNUuULB7qiIq51J3c1GiOlEIwn3OOh1n5iB1qpYd6mVwKw
mSKkOoe+GqsYQtcbgEyTvEfGuZMSSzfdUtACcsWmf8sjig9CJX7w4vM6JaGHKmk37B83/Se31hG5
T7kisvyyCEXgvMsdR+VQlGOB51Tcnc21PhOLEgIV+2ce4uMjpUIY4rP99Yjp/3r9psyl2AowlV7Z
p1da/lJinvBiOG8Hixye0IsGvi347BOepyNiopONmkxRn1AmDKiT5Hojg77JQxwO5XE90Gf8myxQ
fc4+LjFXKIiGi5v0XSAD/6n3ZhLsFbsf73gAVIIametxMZSIMUm3qxihF9Edx4rFlrBrFai9BJwY
NGX5DVKU5PczCzKNbSZX0wvhSvKqvVv9B5JSPs2Yd6hMJAbKsDpzkciq03OCEJfe9rJgsI7CHM9h
5SbmtCvk11x1W32QLq7MYzYVcQh9/RuiWAlyqan0h1lBcydE6V3zJnAf4OL2G2n18KZW+nVTw3gp
CmreEED2kDaHhkRz4kiUfhPmmjVNfeMJTQ2JXQpKkFbilMm9pActRH4na37K9GC4vxQ9hOz/8jPM
y1DDNP+LL8q/mRL0UiW59cmmbYlBdV34tOVgC0rafwFf4Z1KABJIhfvmQaWLwExuIexL5nPik3ts
1JwPXvqHJEymN29H/SsQVuyCAUKNzocGevuQV0K+kzyjT643ZOJ+Mj2YibehuvOydoC2DYB6DKac
tIeW5v5uviUAaZsFEVooTIyzX0J1Yus5KZ3evAnXloclB4bVcwbDnzCmNVs9HNtyT+shFbcSYcAS
wbjpgXpPgZZMJ5xDsMaga4ztrVILz4E0FcEHtxgaGAMx4QIDyE6Pq7/57ImEgn3i286IWVpMpjvS
YvJg5I2TV37DY6zF+Oxd42ORhAaXodM7UAbJOIqs7BWUjKSuZjTgBpDRmIJrnznPvNTS575DSf3W
jvqRLZAxMvnrk7c6PhrOYz39gzKVE4gXC8n51ro39+ljDdIsVxvzcss+CEKWAOZBrTrmMQyFKeib
gIB3M1ivcomLPHBIYHYflYbStA4FrcRa2GCBRzvWNKqeq4K3rvt74R+rmYLuuQWZ6bR7CHIiurbu
+QcC5bbb3mDSNdVKJdtkV1xFuIH6FQO3Y/2+pP4z5BEDxYZCU5yKf7aX3wtYCnCFiP/Tto4s8wWu
8hTxP2biMnYIzt6zR7fkpBqOlCdJCjgjNBeM/SrFY5F0y6DHVLO6064pIYy4XeKkRdYCO6EbVGbB
2R6GmmNn+mlpYRugRfkLBvKVoT/CgXOlIZ9750OR4OHbWpWYFniynduvtsDP9nXlDexnqluZzWYj
7iK3Al6x71mIZjv6Hl+s+XaPdWgh1CPg8pLZBEm6pwGihDNuV19257XQoq+dwDH0GuGr4fkB0S67
4X8nN7R4v/4vJwSBNBNGKvmQkp2btRKmor0HGe8gnWrLOjACQvCL7n+uRU+Hjp284lqXMPSDW/n4
67N0GIG65ReC66vm6U7B9V0x9JZqpAkpAnVX8BEzS+SB1b2Zf8dCQ1wkmz2UbgBxe2pt9XYZhnd2
D0LhV28D329Iz4RMrUm/vJXo4sCvbJL8RzjIKu1N3TVkekVcfLFYwNJp0NTvlfgIDpK08krTCwjr
0R9kkV+zFfKVFeYUHonuQ71sc8BY7wxn3DoZXerhCQJJiDedI5w+fTeFQsYP8sAPRdJkXFrwmPtV
InB87XS87hBAheAaX4hbqRUpCHU217p4DAZLmA38XG/UGsIIPYOukMaupXQIftaSZXGsQy8L0/XQ
Eyxi6IrSIsgGqOc2yWFky8SvvlYgWj8FLXdev8Vx5B3SzNCIGdAqk6nfL9WGoc+gK65ZbiFWc9sm
M0LemgSeKoOVoPocMGOuvFLVhJGWFZ4VW5D+9Bm0mLI3iuh3x+oXlXtC/I4Ywj2k26Gwl0C6GGlG
ZrTJeBZanW8Wj9ikLLetG67BbS0rEBBK2qI48g5z6BqaukMLy3Naa+VoJeKd3AZRK2IZlicAA6hq
/Ui6/R75pEtLAuFJ/rVZ4AMp4wdYHJcXyGu46LW0Jzt0zuCOMp2RIkX73HlQFR+rGBkzjIE4VGEj
iDVmJyov5PlI0b9A5QENU7PYMdLHHUyipwFEfPSXB4JZOALTse5/C4zlCuXhGUhC7ld1cV2nTPlc
sbQBqWAFMMdK/l4DM2Wvdc1XhR2rQSpObITIvTrcN9DcZ2wUcNCahj8v0ny392f1pUnHh3Jfc8MK
4KcYkc5t+vSPdt9m69pdLaGdsNYjP4H7KpBW8A9vfBkEYDrGHkQDkSEUGivwSR0AwHhEZp1XCbXo
MQPeAVRHLpvqlNZOq1oLSQ94FgvCHx9y02Psoh1vhj3FUE/YDG/CjcDEI+J8lFZQKVVW8Yri1dc2
az/AjW3Rf5chI/bOwIMPxhKwFcjFiYOYH93t5mi66PfaBKkWM8Yv0osh6H+MuuRfaexUY+7cVVo3
UnJ/fTpGKeI2xmS7r0ftFs4A6NZpnEfCNlK+8uNUNAJheRl41n0Bh80b1TkUCF2we4ogpJ8GkLGi
JPm5b/eTBjv9l6BUtPV9PH/st58sVej3zo/mjoW24ZFkxYP9L0M+22X5aT4LCwhWzavgtF07gBbV
8FTIZoco5BXvIczSvog/+iLyzAqbI3alEJSOD5bKIzy0pYdXz6lIaa9XMLhckctMfPliNLBCsOe0
s9xNJeFHGdodtHlHwSqQS4llkaJFYWmPAZMB66wu8H5461XCcwpbavsVJU2eSwSOK92T+JXhTS2R
rKFjd82gMk30YrwyPdoc9ICwr0J9cW7pSKyrAllnN6tCXc307twl9VguLPkiXLSxIass9YPdYHAw
xvXUFBooVBh2Z/glOeB39fbhfJCBTDnyMm9TuyK0daCEWgq5aumyueShc7zTXPWMyez3rhqsuevF
xqSYalxDIeY2TtiFDNqZ9wVLmC8ta7UGsMCZl94KSEKGydezdrOv5uTFo4Q4NFAl6HOM0G3PjtzH
/1M9gKz2+Kon/tFpJGZCeqMdvsvORtCWC+mTicO9UnmLhdbdlSHm0TnPhEvKP7nQyKAGv7ImIDjp
7/K/leA936pWD7PNfrhjWNf4rTcrvvfvXWjpTwxMLp0kHuJtKRrPk6tmdJjd6XdClHm3QDrytPAw
bGdRFKa2/7oAl2GRT13eZr6ptmF1rmtZWl2fvII19c4W6fUmQgFfOUatyYx9x50yQUShFf2VgfN4
natRcW4np5vPaltgQMtaUXEVzi8ZquyRfjyBO9CJN2UeTSmCZv1efn/gA+G8TFg75o6liC2EzZr8
GLue42Clh7302mQoJxXDBbCtiGcQzqqHlTc45UrxYIXsKiPkcRWzKdAwRJ/ThNhXLkUBcD0yYSUj
TgpUdU0TJ7UAekk5tgaV4I4oBJfi5GFv4mi1qTXC5/bdziFuMpz5rBI6OnDpX12o5lhow29sYWCr
aUq5V5Lm9qh6baVLfcjyPti7DgjlH+WoNjgJwA3/bq5fdWNaaTnu7eaXjy4bGq+l3PtOTQsF2ETq
hLHeRx7xxCWIWwirta8G1KWUSy3tVwo7pARPuwh0/codOU5zrjsDXNLzqzqiHkYSvafaWUFgXZCh
4dQY7XdDmtP33rduoIA0QGA/TR/hBnKKy4QAOn697mmZ6aBJWm4hAg+BKgIcfTo4lMY8JsjLK3sO
ie01HjgffLFGVGbZZ0ZIo+KwuKv5SqujpRZZAmzl3Yz6/Bi2PlaalAg3pQmfujbb0p0piF+7n2FC
Sze9D9GCnfiWHFQT3eHVUiCTm2H2E7Bb2dwWxXsXKDMii6AU9Zp1+XgBdpVNCJ4WarR8R4jNDmSB
0ManXB7RUNwtewYRQY73IPcJhC3/GPAezf/AR18014sYe/n8l0vybA3lH7/FlYzuuv0kuWWV3ENY
ezLmkUm/gebYGxwgsSTP8n3hR7Y2gJtYdJHB7cEC8/MCTm+sD58ND+tJlH1M5IJJ6h7v5zFolEzX
SQ9JQKNan0o3DAZo3GgTUdPHpKVe0Zs6xeew/AYzn0iOUYcQWZ4QXZO/FCYqmcjKXsQlQpF7d2e4
uOU1yxupUN4N06xDGgevrYgCe0czQ5/lcniKYi9s1jUNGW04OLkYQuMUwi1DKdwpf2D9H2v3HxNf
pimtv8Gfu+PXq4aa+YtiU4AzQ9zwr1cn89Z5yLlYo1UthOrIq2gPn+ae12OIF/Nv26USG2dep/R6
h7GLRzvxG4BykzKlS+A9l6gr/D64AE9myMzwmey1lREIzsNJ5wqk6RQBr7pSFec4SyI6zI4qfDLo
nhTVw6sK89frQdNSrFPBnmSCG0acgEEpLJSD/s4+Kf7YrIrkPm53T616hmnW8mOlsAQSMPZAugSL
qHGsvAJVneNXu5MKrt//8MD8ZpR+8RD7VI04XlZJ+rwX8EbZWWOLVWkV+YcPf077nBLV707ug5rV
knfvOsRdycI2aHJaioxYwnrudR2xCV0+n4/0yK+F0zbrz+8cUKZtiofcaOfdxZ7g6BEPpxemcJKR
KGRBaMgEFDY+N6hoU+7MV/vhPK92ysN850KfgcMtrPd8aHXcGZqb/KQTJFjcuxPMO8fPv4uhrorM
wRtztq+RrJIy8PLjp5DGv7pQTNyHwqvFUC3P0/Nuw1nlJcmzD5AL0A7CPj7qAHGrexx5n2GXa3GS
iaFpSuSdEEpRGeBgC5vUgx/cCWJBFdH6IkH4IOnubcfMZCQ6263U/oXC+2ViKLsV7kqGK1rt9QTj
F81ZhUIl0mqarmUAfiktgvMaE49ioqHa5dcuB8ukkVDMYGMkrowkNP2cwmdyjan3sGITCtv9daf+
DcJ0ql/IDwFXXFQgUxMpQHR2Ff36HRVmgpW/eT54Yx2Pqpe1sRhXnDUle471eE22DzgJN9P4Ja6r
UwYaQbuTY7YSDxrCxhGbWxq9QUlawBvaKJM6CqG3oa0kS2CRkDbYhDntoWzw0mC8Syr1r/903hqA
LMETeh0XpBthKQ7EO73xytakrK+VZqYQnMkYXnw9PLO1UK85M1q4Xu/57U7iT9w0Nrn56Zf4YTwY
TQb5VDGKp2JN8z48KQX7LQiDxI42/6Xiw0HI/bqx10hC3IMULqJdD55ooaeEeTgsktm90K8LdgyN
1gU3ZOenQB8VGTkjLW6OO4mCS4+O59KQJPOsm6xI9ANNgTuCshRGjXYukGuvBcXpL7s59lQPDH+7
bz2HgRNq6kI9f1P7rNtGsiXUoeWCuVcPDQ2EgTNWtQ7qgmwphvrbD9Oh8jyCHIJTZFJusEZ/lab4
KSDBR7K1DgftbK1a0QJQg09paqVfZ15j/FUpWHcnQ4Bjo4v+bWFA6Mm3bALSO3kSMWqT5xwloX4A
rbLU81hKF6v5XuH9dXxY4gqD895pELv0dTZ+DV/MUkrbEcE3nKF5gtK4/i6A2eaFk/3q7uEVA0vu
kaGrx0vI4cPObDWsPxKJernzBE+3LbowGs7JTGwdPTw4uS3y85zYv9XJb6t+0D7VAqJcdgYujmwp
CUVyOFOFbJHqgSDdumlI9vDEoHpFze8yIpGEpumBOv4lrzrzoRg988UqwFSNymTdFcHb7IshK0X7
L8KIzf42lj+qGCgvDhsq9Oug5L+4nQZdfx8RgLE96rDMtoTgTyKETBklcW1q9Qhd6GNlYmJzCNot
BmqSEi/HRCm3ZXf3Jenw2NPZwv7SfrpqEVsT2OcmlhklMxtbV7m4FRjBNVRUovC0/LvfcxIgVhaK
X5Sd5wALVap/WbhyULgf9U83YdX3B7VQGMZmoj8E5sDCOJnD+1R7RO2iQ5byUI3WbnWQ1IAvNCQr
sdklN07vdcEOFmB6Eest7wtjpFp9zimetAMCra815cr6ckzVfNTQfvhull48rfDpgV+9fJEbtR/J
AMhscl8w4Vcc1swTcJYes4mh1RzNeFfgiVuhx9OK3ajCbYOybqVtnST01Q9OLL1jDyCfQwjehjYz
X75jaToicJU6vAzJk5AJnSGkaEaB3GFbf8evCrkj5w5/6Bw0XzqcwABgOXaHr7hc3aPD43Ziyv26
P1yZ5qtrGuczBHA5yq9oTJt1JAR3Vd63ENQKLTEQPm4SIwg4Pycw4E8LK2bRrZLXpTjXSaEpaPQT
mpXsha9tU4ug/nGtjMViTAIJZFDAJVV/j0d90Y6FkrE6V8MSG9XkGg65z6GqixlWImstnFOOwDmx
0DZGJyjbqvlDleSd1RHwCmB93sYLqIscSAelY5UEc8G5LHUoqc45vtKP51QSzpQuWvN+qdbOu21I
CGp+Eo08GWczusvJbl58PdQ7ffsGWgdoEzQcQ5WSuwkpKsOCGl1f1Y3wTmASjCAlgu5b33ZudSlp
jWLuO0NA6JQJ/wq4kseh/tKKvgw35p9JI7FdW0FA74sR6ShUHi0IfZWzZ4OaiSSmLxDMs5ewHD7L
oVbsWU6Z/qFAUoXsuMUOVlcFA0myxr3e6R+/wpH4Td4TsgffA/2k8CmAMuAuaf/9Vw5zFiSMipIB
DgHSLlDqankRyzgT3ZXm4nW9uZv4yFhEiLBAAvXgEo9cbMjkdkTEH9cfNXofp+6pnzTb8PSQtvQg
uIBSoXo5N1rcAQT9GODrN8+3sFL8e8T/5EeOm8bLE8i37+9J5TIelAwxJfz1EhZRE0zZxo/duWHK
S9EgbsyOq6judYSRdl75J5locYVpBj6xYYaT6+vq+WaBHVi0PIfx+VBp8xGFrZ0GeCW9rj7OurEz
DpRvSIpI6fws5J7l2+5lUAdopvTqighDCTluyAJpugb7g04exeUPCjzew7GLnW+MrnJsEUCs7VcZ
MMt0LbL4Hj2JPqmyN4IVlJCNbrqHR2S6jLhWj+VQAAGeNouoikmJkkrT57TojIQxA2UsbTmFUjOH
bN18gE6G0gVUp8vO3oHZBVbmli863CuNJwoCFGzQWOzjvOl4bsf1WPGV7hjdtRsAxVkgfF3L+ryn
z6+fymEdumf5Pg7E2O8gWdFyBEeDseQuL306Elm1XNr6pa8H8C68MxpLc5ZlCW43uXdONuO+gNOu
Y/763S0UOefg4H1/NR6pb5Fa5SvsxVpYRiKCopeQafKDWRHxbisUIQNAAo/Garlh9OgG/lgj8lpe
a8TgUch1c/ziSwPfBZKwxxiYbwLfDskZMj8sXHZoH+D4sHfHwcoG7jcmis0xTAhi+NnvyFhaBNce
d9tLaoecgYyzmOC2XnWY4Yh22SmSsZ7PCn+URUAfcIsBG0hf0Xkcq630KhKM5KcDut1/BjxfDcmj
yxUsqrj4SnH32IvWdEKWAkDGoI07P96ZoKLs/aWlKBB1FFa/OPnUDzkkLXUu9KM79uJwPj8SkOf7
v6zAfPLyjTy33vIW83lO7N4iF5XeOX7RsFmLecbQdJC74Yc9j0k2FdjDviC95O6fQ2G61zb6J61N
ihjx9Y5OP0oq+vwz8eWJDhmi6yMaFVgwxgXlS7KO2gHzjrIn5sB7dBrnKgQLghN2imRCgSsEkOri
qSo/AtIHc7KrCXqKVaIzV9TjjLmD+q6x1bTFH1av4EkxltCvTSbdzH97ojkJjhuJC+j5OnydNOJy
KkiI6yMVcowTlPoMtakHq2QIx9hKG5C6nhP7aj8xQnjn+ybT9STFkYzvqpcCEZEkpF9M4gnk3Y6B
GshTSK8d19sIsm/sgGdrxzAH5w0E3iCfgACxVPWtkk7MSVfmRYNHg+a72owIZ2ipSXsMdavjxu1t
M1hwJgfLLZnLWEVR1qRT8DkrkzYQ5pXJRfceHaueH9+PqBGtOGGov7Hlk0hUevF57CpdKzDR/Ryp
uvNq9AS/qbmo2cRL1Z/WUdqAym1LKadVM4+GL8wlZJ2MUy79hYcNQKFhFwxUHroitNY9bA9MGFQw
KSOeXQJIlM+4X7oH66/psQygXsM98PNbdP5R0DxlcqD0Ry/qGZ65ke9+j/F+uQChmk/iYe3zcoEm
sB8rN6OGmnTEhc+JjW3YG8x7+v+Jn9L3dShqdJEPP4JEWhd2F6/nsVXFyylqwVo8XNkHuSpNs1w4
z2YHQdAjv66yJYpBSYmLfsmSerpxP2zlZkOztvqWxxuVIZFCqru495VBeuHcBtD4rEZkT77OoAwA
PB0u4D64MbHrJNICToL93D854xPfAO3Tb2yG890RcxTTs6crfD2VpodAc8SkW0MaYbrTmAeNz0tM
guHmIC8wjjvkqU1o22CwL6OjJocttGgCIhG8F82DQ6OaOwN7yx5AhkYNlrYbBfQLGW0cqGC9BdlM
fKPd4SPZKemao9gbUfye35CiewCeen/P5u7XujqYlaTMFeF0cNRhgSHg5UNtcNYwKdSulp/11xTN
8zp5e8BcyYV+VwIMmJDHwlbpGvVeuMafG8M5FXl76I8QOuJ/oOGeqnP1ZCYL49kbN9D7Wy+cGBdN
AGx0IBRLfbaVoZszfP8ymS2WQr2niJFMuvZ79O0jCWwXYbOnK4hXHShY/zivfZNvgtyZ2pGIt5h8
O7dj/bvcGtqjZC/s53UP1/n5loXUK1xuHbl1j3kBccl2nLL92S/2H8NJJ6tfytWapu8O71oULwnk
Sm9ke2iorry8iMu8Nho9PHkv8Na/z+yc1+FspK97/VbxKTdZi0DgPKU7LTTtpxxFLrce/yvRHEr0
PQK6lTTiykmRPqx3epYczKNTQWnxkU7qwOfp+BUgi1g4TJ4lFFyXQikg8z1JT5qh0SZpT5AEkQsm
Bzs/A1TFYAzW/0GusprRBrC2+1RxZAQDY/XndzfzSNcetwCLjrtJbZCDNimyLgnf/E58IDivUJ9X
uzYHNW++X6N50XFF6neWB42HX5cVj+27VwJyEVnDst7Z4bTEcPVEPjRJzYxhNTZDAb2cbKywnIOx
oWa7uRKEzGko4zNxsWi3JQNmbkGswIZ1NBbycWb1YJX9UOV3HyequPO6tL668T694EuhHTVa6b0W
CaMwL/f0roa97zyTYghet2Y0ha8/reXcq0txU/M/5R+5/NkuGVoaYQBi96Asn+2eo+Oyzm3wb1nJ
tptSgKZNtR409iZ2BQhpg0BlQZu9edBs9fZggDHRpYQKTnLUBA+aTL2zmwVXatYpw6ZCdJkg8lZy
5oEzNlJj/kM25NADRc+YWpcwApsZerJk3W6tkNmxHsUe+vmKBClJTDz9eRlrl6CbQyK9Epu8Jxoh
mEVGBr9c64AIqPNrW6QFeLLFU7iPxHSTNvlujzgpeNl7g/nLM+dLUGjaPiUd5GMt8vLmigH3VdfS
Wq8fOkix4IAfUBYS4dk1sPx1MGIOWl957ojMNDI39YuzcaC2yDUtA2VViYVOQipC0y7Gb95w0LBC
TiKY6gFIMLRhpIcjrqlBEARnlq8pWelJnFhSzGxqAgJtFHrc2FYBbQSQLe7B8N6Ub5kuk//v/WhK
UWtfngYX8jXjuUSGSX06R58xI71oowFbUh8ucfFjAXm58EMAtACJCayK1w8qSrTbqHq72KMf1DYb
OqQ0Q5jZy+HoKJ9VtEs2W6A25BaiOpy1mSEw8t5giJ0laa6fn53J4YAfaX+EKBZc0zWTisakOhrk
NKnco/bhe2NtJervsExpXAtCBPMaJcl+HEF8I6+fpqzziBkZ86FxFpVrkzwWOe2hHQUpYC33IMLk
r1uahxjPSA7WMiUXIM9Tgoyo0ybnV9vkDRFumEm+S+10jLclXaT9+o8q3RasLhsPCloP0FVQOgpC
FEzysjShq2jxTFai+GogXnE66xUYfFlsyUWRS3SsWnSHSYDX96IwTKHkY1NfPsDG3R6ApUeTkm9G
QcEIdwpw1UOaf3CayJSNjb37M0XZSMH09vrdV3kgn1A42I+X/bP60UXBaWzTlEgHRzG1spcBFmTH
ZtCeW6cJQ1pSJdVLtoKMMxcpsYydxlgYFWpQLrm3gX74uXqSgPzap15CUnG5OxdCgQgJ3Jj9bQ6M
CB15dRqZ5RcTiUhWHeqQeABdmihoCjTmshLtGW66lBYtxqx4GHkJ/zURuF+2EvgFcLdK0HVWcglf
OHh7BCqXZAKW6Pzp4/NCCRwxBp/A1kmFw1S1HVU2YsRHzXX/xaviP2ZL7VvOeNdOTP0gIGcQalRe
t4a41UNgzivTy96wkB1COsRaLDMTzi4kRRg0AJMZ6eJLJ2rRFh/yh4gJqlYQXEFKlvs83DWL3kJ9
PqEpPv/3tb1FU+1xCsp9YO5e52g13iBILb1gh52nAdarJyUXKgnRpr3WIezZXsPyRLOsgdHYczkK
JdocwiRjZ0BupMG9SYl4hQ2n6+/8sKfaSWuElfrwxlgfkXQf9sRK1FpINLM8V6WXksU78el40k/i
aS1w5saSoQToLbM5YSQ6wKt6MMBerGd5mGfpeDYFSchZJ335vhnd+D8WAzLx8GjuM+uCjOg+ce4N
KmnJNxESMCwq7OnUzUGvy6UoVBYW1Nk05rBNqCUAZyR2wisS1+sNH4VeWx+eLQs8Vg38Zm/KdfxG
6+4zUHf3iZwXK1xs8CSx5iZTrjSGQ6jg3kbGJ3DnefFAnPbIrMIsOWC3wFVghJmomPMQEsmFvJ8s
1KqianuH4F9/KEZ+c4sMa3/mK4gVK6ni31DL1Yz8+NyoRsW72xXHcbKfBRcFMD9yV29XfJMDznLY
xGrEd3aX0wzeAHyICoUO60OGIyBCXycgq2NsXmjWxG+uP4RtA58CF0AMFb4lL3z4OD1wP273XxvJ
7F3huwL+Qu6JbbREW6OUfKIqrsj4cY0H0nO48kEtmlXTMjTAtO20rRJaB4N2ZSu9mJ+HbfkI7njk
JeEJqZ9Rt7hHX5yYDdw/VilcNDMI6eIJRrAo/52dklzxI/6lGUicCuG/ThHviOUqXptWcGkT/H1g
Z6+opi82FV1nG1uDrU3sWuWL+7kl+qdY5lRo5RUBKqpoZJyE5kUmrekgaHy6/wI25MIqwRLO5NjG
sTF5O7EfDkLQQewd233ygFJcd0xDalQU9BRlbyW3ih6pXoBmyYj2Ka5xP+rBZ+kJgBp6b2wRWIHB
TsNGwiNHPJ5xLcB+fyvVCI9AYfjDr8SemQU4jrNzMRDPKySdDJSBz5h3xD0ksHmeJpsZqRo8f4Se
W82LzN2Ckcyj7SN5hbqLxGaiTORM8NhULLE9LXb6YbxYCNztaKjcveHQM7NvshuxftjwW28syE/7
BKuQZmR+0RnkhJKf6ZiH4bTvMtT53V2dM8nK3Zblb6A8fD+1XFXbwrwwHX6lKWeJvQ6H6LaZ7qDR
XPPtId5g6qr1tbg/PAMqXpYKImQPkYJay+3n8PQ6dTsv7plvCBQkKEIp64FsNZZEtMzvFAJSvXyn
yXxpL1z4OjK/KaN+LYV8Rg5CsDaHf2LcBaJKTLF1eS87hKWj7jGQ5Eu3r+JbpBZHlkKYpBXW7sVc
mXMmv8Q2oqrOp3kzx3rHQO3DVmmboDOanu1jbUkimZgFwc/UKLFoAr/nikbUHUYt4fjLDsaEZPxc
61P5meJfgnHx6Cbvk1PV4vg0W+lOpQ3AnhfizUE11ZcQBnP2195Z1sYzJc48gDgmkiu6WwhCaEKz
bZnNCR2LuPTkC0uUG5mnZkwMR9qvDWziM4IcE1n5jjEWsNbpzjlIjdEmI4g21z1f2Wyz9pZC7tfI
Jth9zrArJ+6iO9WfXXiaEF7Tj+Ixi+IoL3cDcKry2pjAjH5H9qCNHRGYLB1yefCKowDGXDSiNX+2
55/TQIiJFK4D+GxzBNwuLGBhriBxlF6+pbKnlL70k/6eHyTvUc4c/0a6avDfLwrHrSV75kvmwYmc
GcywSuXN3W78ZDXK3LopMKnkxb2a0OI/YKMpbGzIOQ70txa/+TVIQC0wqGMfzvjVjhxjhRqF3AMA
tIdH/P0lOalEfXn4r8ru+YkJ2m2mpIJwmdWVtdk382OFo1Td8oHEbLHgShBVmolfrEP+ChnajbLp
40zIBFGjYJdXcuKaX34eW0P5IGrNn07g1DuIccKmLU2XBGnDcs1XPr0kL2oI687p3jiQz5jr4+Uu
+Wz7C4SBhvENHFXYK6x4Iy1BDrk1G9jWEY2euhJ/aU/hjmrGh21mFY0V/pDS6Y5eUjlPC21eLcQW
hiDcOG7T9E6ekD6nDvTiZPS5Kd3BgSAhTtG7t/MoWbo6FtMnYB41ls5ERCtXjviLKhmGlOjCvVo5
/WBGq5MKwyfpsq2UcXQyGDE6gEgj+iYHAZ5uj0Fvc51t1NIaAOu1vzCMX3TZVTGc3aBnsqkBP7MJ
/IpZTtm5uU+XWNY9XMePf0H2iO0FjPGPHSt8UKYaWvLl4fOLETMs4rZy609ZslTB3Bi6+0ffzJAf
WSMaxh2ha/jAEt+gY4IVQM7cCepjG/xMhuyKjnarJN3FlGK2w6G5Kn4ePF7x8TcaHKQIarlsnndG
KRwp6yzfpxf6Og/wvXa/J1leaRvwlcW8vKx/DHUGNdUKs0nMujfBfv/r3Wr3fJ+i+QpX2PCC084B
Twypa3yjbY+FzgQksGer9VW2CdmkEJENnb7714Zp5KwDvDQqKW/PLqkUXsI8ciisb81qtQqfrWP4
QD749xuajQBi7qT5A4ybFaAa8PmKMqPR2Cf0aniex4lrl0MBfqz5CwKM4nxp6PvYE6mcVdvlvhP0
xjiUrcypneTWWio+blyYt2ZRVdvctK9omjsD/l3UQhtd3qQazJBRpkizzMwuql70KKtlrbXo0J+U
gH9iAYD8M0FtrMpDBTqvfa+sr9CegX38SXJ+pvdz+h7g9Hwzy088Wf5CQrDumJ69CBfSrUaTmsbi
j2zQijAiLpyQyHTUZa0/dffJjTv6F6bTE0PoZuEJub0y4ic7hKakzC4C/ey3hJ/bi3OG3WDuz9fi
XSJi5GVJUdIZA6t2aCxQASY2vwNM3YrEyJygGrthZUTOyD12RiwGVWtNsFPJd0nae5jv/d5e53zk
Dc6EMF6KVNFY8x1D+hPGqfuHWX08PbdP5U9Ex37/ifCe4J8G/hmxAbi/QPnzj4TI0Hfs5jCUD8mh
eabZs+Uo58AkElmbiZ4NPLTJ/iKGB96354xZHondk7XIBcN2fKlLE2FQCBDw+QzzWMQM1a7ADUbf
kaLk0s3CiYGDdpScSHAv+pPB3xAhmrN7dztSNehQInFYjL58Gnp+wkvnzxnmOK4ZZkgccbBaAaE8
cb6GqWfUe2NrZP9geZuOiaAVc+HWnlceOTrH09PGDov2KzSSZCqZbDqKAfkxndYAYEgOEzapweH6
MGhb6swdXmaZgHdduyIueVUECtOOzY52dqFj9mQZFUCObFkVNi+YTi5sMWfxluIQK7DpzFTnS5dR
GMQK3VRhHlwfaMcs+qh7W29RPyOpIbxwmgw/NP6Vf/P8jVwLeTOkVNJFd4OXMb6X8kvEdmI2CYSz
+KULplxfmTqSXgPy71yUuL5Dx55z04TmkV4C93kZXtvd269HmRMgv9byTVdnzYA+Rt8/0EkEM6Zy
wSstrgjR2jYtPzhzzdkwfPL+xBjbyrqUl17Cn4Qix+i0UZJTF4t8UXP6DHb3DK7Z0smiCaaSgt/q
gJl0XiV+WTgfb1kYizWRDstEhr+sn4ru2TWwOFDubUHxZZo+uPB4YywLiPeDim3tzCgaXCpvqZyq
9Kq0gfQ/ymPQ2K73wrR5tq8mzKskkD5pNPLJgLATMNHxn6uZutAWJ67sxo522qiwSXKa096png+w
EKKllB39l/33FSaKPo46rRyl33Wgc22rDjl3Fq/4ClReYSyuMfqLQIqRx8YBSpFn9kSDCZCF6K8q
/ytJqF873L+RxO+EC3ghRfwNfHoKiEMpY4jOtBsaidOLQ+xrmS+GELr6V8Au32+cJr3JtBqFgbqX
tpKj+iM27du8r7ogNlyFr8xnO0Aza88n59th4RaPG1d+oyUIvRODhSkFIFXoOroQnWV1CFEKi0Lw
QN7hFuhgVLVjdiWvWSaGZYP1lPXJB0DYtQtFBh/bR2LJY+qef5Cf+OazbK/gNbqJOYgYZ7+hp2gv
FsGJJX0wy/RjSwHl3ZSlV0f6/WxJVjTzr6WeTEwPKqRp2cT7JdjkVZMCglQ9p0VBVxlnJeEPxcjl
bFUgSUfKS2Pf36E0iGUm2LeFYJJl5pseZrFVMgbKiqNvP43idl5w7TuyBdfm/uGnzXdcTG3+sBx/
QAV9HPUZ9g98QfG9OGD8r2+56Y3GpA0af18nUe8i8i4BH6RCSOOVMG1w9+kFZJwf/EdnE/LbeLPr
lV9ngp+iFhWreneH4Yasuvb+E9uTYYHC1kwRSYmJAWXe2BQRlO0P6KEvxR2IPng594SIx+nJpD9L
imKiy6/5X79YIaQmKamXsa3ZkHKf5JX0RRUJrueCcmhy0hrsew3IvyYvfzxU2KFoEJgiYrS3S3Cn
5BfUAAz+wYjuFOJ48onSiTzaZXxRvyufULKXOV3H0TAOBbLpFBEIpUrvuk6A7DcDs2Gf/on2QIsc
LVKfJqvp62Pv/tTYrGGWOKQ/Rljg7vgzWZVdbuH7+18tEjV4w12AkqmooE0hUcx4ZUj28Iftdpyp
G+CVgCzW50MGlS1o/MVS8kK7gcG22XU0aRg5IbC0DxWwNKd4lUeArVlm5WFQljJF7G0fvgZuWjp0
kx119mwJyhxvmL9UngNZtWF6o8tGxd342mSV9z+0vdMn9H+D9TjRJnP+9LDHj/qcUktgOLJKcamv
k4A9oCBrsdlJsTXFz1zepjjKm+aFfFdGUxIEFH1o5mG1CNAgPizW2bsD2zHIe8ND1kXRU5l/05r0
VbCHPXEfwn68uyw4o4n7jhB+ovuP1U8n0BnIA6hDSoLh6Bf3YDhfqk15vQglOPfPz2+xCUWH/GgA
DrafICclXGxzvEsXCAJIS8s9rj9k1xJoqDnjYWUpCWLlStNwKmbfSNpQZCVEnkSEnVWDNDhwwoh8
j6klX3JxaZ/nbdf9GP6dK42YlFc+gklDn1N/He/w4Rj1gYyMgQxkrnXTGDX0GArxdOuhuc6szK1f
EVfWj93iBbLWxNZVVCKhAL70vf2iQsBBi9NhRVmC0zmnddWKrXR1bsOT4/IN+Wd5GNvzLeVN2row
+v+YpVkitAIMIx054tqpUg0l8pTD8bfBelD5jtMTMLqL3VRYM26Y1/DJrvGJ9kZXIJryAff6lr8X
ARBaFH3PC10PftWVk7SprC1yoOz9b0LHVFMnPkSaouH9fOKOvUt2scXT3WxjWuJvjL9qhEEBViIx
VFxHoilpKmWXBCf+Pe6nkPp7zOe2pwAP4NNGI6WUOaqz5oJ7DLHeedZN9MNeHuZv/I+HDp3ZD+ip
X7G/HwrzbLCyAspsT3524siK8Qdsw9Z8+Vf490Mzxn9Tm8EEJTLqzG1yN6y9fvYePzonXlXzi2+A
ctyYsJjIDf1Fkj8jMhhd2sWbtujHC9Zv8dL5izIsaoMftVKFIIKdruyIRO0/QowVrGMCdXDp9vpo
UceDj8u2w3riNt5q/GE9UjZx1+RUr2NrxJ5KPd8rtHtcPdISZ5Pg1+dZvzqR5KomQpDUbY6EVmiO
wa1VS8k0ZEsFTqJsA8+35SM6z3P1faDVY2wy9RwX1+IeyPqkUAFK5GPF7vB38CwWZBUBtw6thiNz
bMQc1Xz62d0RMBv7Vfxk3bfGX9/OQ9J04IX3acpR8SB3li161K9qbbUBSAwzNIuK0oOLL2cFPxrZ
FMS/AfnO8yDSCRGdCell8YYu/lOR6aTq+zQveWg+uvpQ8ZZmAc1ZN03JFDia2QFM0D2YshS2U8cX
agi5jTvv6XWZnaed1stIYq4rM9tXdIET8xfuZsR7y0vX4gZIH1ojvYE2k8DAqe9W2F8BtOzAHD85
a64Ppi6o+/C+YHrhG2FAOE6UcX0jy+ff1kFM5/ijRHyjDtL5kMbQvwiYNQm/homoT61sbPU9ra+G
FsRG7UtA5b7OtrZCnlFWO5LYvqr6PAD0J8IXGElIM+aoQ3uXmfKg3K/+OgSHxrlAcrxWPymGLZE6
tcZB98JxxuzfrPqrqD5ioTlcfX/qqNeA2o3CD009V0XV62rDUDx8rlG56uxy+4MLX/3d/ZlKANYX
Cp+Ex9YFvoKXnLMImBsjhXRxULr/EnIAZp6NM88owRDVu8EHQHW3HajOndtjdL/mDGUDmWtzvoTe
zgQCd8oZ3klv0wCSduBZW/8UUVLvrs3ioLIrcflLHofhVN3qdjdLAKulndgwdz1j/S95O3pImIfg
pGJE8Z5XtVUSqW++ePxrFhih/h+pLLT0Xq8V/aNsZQAvqPQB9EfX2e/W1FfACp2u+fgVYD4aRoTz
5gmkmMAalGivIZpZ5qXt5EYtEaBL0Z+Z1kKbL4EpdUB+8FQO821d4irAHiTW4gXEDRUiPNFtmVV0
46eIJF5+6cbg70wFv/qxgvtvO5WlCAbtp3U0Ph84+wF+v1iB5urnvnDwRyNewqIt5lPJj8/+2QyO
Qmk9DUx1Ao7xi+qUz7wSWvMlRGW1yM77kiPWcXu9O9E9SfeIugcUgntJZ+jwHJK9+okQVZcp/hmw
s0xRQiQSjfZNK07KYIYo0IganKSMkhVzwV/gkT54Hh6PMmjtub2SwYSY8tU49m6+XAsuDyHz9kAK
+6MgSWJbOrM8ADeaXYDqbOyixGLb6UDgL4Wrr4ZkCT+0Yk1+tPczr63gca7bmz8zfhN/TOg5qGaG
7p+NcCUAaPnarBtP17MSPIf8sRWZZChz23fRSggFu+Pg95cQvGoSKenhcWWUdvUERHORfBVsnLFc
Uxhs4zRcpXrMmI29+d1Mq+8loLJo/U5HoPAxn+OP+QljBL+wCD8Z9cBo3mcqKZTM2pAWCSlZvuNz
bRqLX0giUnyuDu2lXBRB+5e/su/L4YFYoOm3fMv1cTP4wDjARZfh0lT4YjYagl4cUiscC4/Aaamd
VS2vn76/SfpYTMTpvCuUd8Z1LA+FfNnQYuvqnsqaKqXj1Gm9/+gHvw5/ronn+bdSvBrzTSdqR6dC
/6JDsHhnw8Mm+g/ulkPLyRw5LfijQljogEgbX9D0NG8cUqErKiX1rHuY0RJn9i0IB9VavyEWl8gA
zZBrddFzgTErqQX0bkHWtFlb4gDCCucbmlKq1V4gjVOX38/0ORtWmKOtKH5wAnBCkNFXDRB1TUG9
Gx6Ff1vTrn0IQGBTuGCkJknfAsAEUt6owyPB2fSNr9/SGT+RzqlDZNgWuc8dtZxz8N9zBf3T88Bi
oieS1a+1sMgQkofq/Taml8U6u20md9JliDjrMpHawHQAIZgmFvJk3tCJrNtczn+5dNJKkOQdFHq9
YU/gDKWEgD/TBgOV1yXMLGOxlhTJnmKNKXvoQ0vnj+OIxMdfA5pp6V5QXPkAnHlLBg4I0iW4dTbt
Qcjto+jxNenvNr5mtLokw1OIqxuYQs3WrskqijhcXsLz+DZwGFXSj1pKOdJBz7Yk7yfguvquQyAn
EPqUargkXFxr+8I9CuzZFQzqBaCS/0xjBV57djmYm1kmzwII57jxyc8aipMypGeLDnykTNYyhy41
uNZooPShYzku8fbs5BoQDG28ki/QOY2IQkde8xoDtRCtp6j4U6P/hBdznOqQDMl0K0rACkif49/j
MyiU04a7dUHNNVDcRaSGYbLYBLFQ9p3ipPqBLl4lw4W539/kQ7T066SoNjdScy80uqHfu/AZzbA5
hqDvry/6RYfpoeSDO+XG9x+ZMST+MVY9Bhek9QY0Vem+41KF0mchamxzuI9rqlQeUJgpbxCocM5Q
agbQ9Ixk6mVXZi5Fz/cj8KK6txiHdVhHp/+JABabv6WFfs/REEZp2FJNtXNP2wavt5Ryiou+NFiU
bLZ+hMqywCEEXolRjyr7JtIBm3urGyCw+62kIvvuzseQhV+6xcIW1vKrqX+tC39SGDq8JNBsXdIb
WcC/ZoULM4wHZsT36utUGeoZva6vZDd/S3zgQmowuB/XKh2RXgnlCIAUabh34wJxM59LYKg1f2I2
zqiYVwBK16FNx5miK4LDrA5AkBav3YCwRo2Y/h/T8VJJk2vmbMnLOiicohmmCSiDWKRE00WN/5nl
f1koDLnders00wETf3UHLovQNgM/5FKNRF/dRUXfi3/ZNLNx6uvzhSnqfqGxdKmhC5fNdydQ+Mv9
TNFm78rTB5gY6FEFaAPGM7LEaqoLezNA7ilf5py/GHWMunHTYziED6pIEBES3OCWFShFj08NkQjS
VBQOuN0+xADyRhNRiLOOD2WIPvPcB4jDno2ifL+TWcZM9uymhOMphvK9DPsKz9TIgltpdw5mWMbA
lpITQfcl4sJruUFrWc++F6YMAKm6O9Wl9hb5V+35uHT+jBCS4y52RkkUhYhQxchkC81dVPoxLelb
e2Ok9xVNTEC6q1mLuep254GNUcWIz5AfyQw6N7/uyG0fbOvezOcNU4sP6WigxPBU8wtDRvHx8IEH
ECVSiP0Wk0IwYHjS5Ca3qbmb3QkDmgoPazUu1PuxLjRE6rXVrpY2Wr4rM8wM6R8J2bczcgDSewH9
NT7uXkAZy8GDk1qGSClZh5++KT8sGLGZlshr09/fkhZPJgGf0QVcuIOhGvP1WQJbEewrmKbzEW8C
MLJ1sSD1I6w6tcnU9fwpoWz6q1EUz91IZfMdm+tm308e7cc20ls6iqhAjE9PVrp5S1VxR4xWcDjk
EN0dXDfTw3Yp4kgN+3KOhxJ1TpLDONTMrELeSeucHSSewAg4ORKGTu6AoARXevPMJW8SSuRml3fG
Ol0zJuXYUOKoUCEz9p+KWgi4NDQknwr0Y8+0INuLucnSO1kuxxtauQbdtIK3d27mifA0i9YYm0wl
I11eE7VTQUPqKcj10ighVWZijY7BlqWi6cKZ7ioH9U8olEnf6A1ojBLat3a8HBrCBEWNPbRFphLx
rg/Mqz3tCQpWbc6r/Wrg20pGIk7YgcRStq+GpYLfgbvohCt8wrMN16/4GWfTsxXzuBn8D0WaicHz
+M13d8H+CHJZvRrsOKdMkLVpuVbzwlDs2qm0cDJMiMelhepf/ukVJSo7Lauz9lLoQzZmELg+HVmU
l5LUHV5lYa+w5VkM7qLu6SlRKP/w/Syq/TXoizyWLwvl88ecn59zCnZKsGaqDj3e0TnX56g3qbfD
aYFwAa7DLcDwe8K0KVqTPoBxJKWJ1IfRM4rTVua991OvrmVwhEr9t4mSY47jUeTgd0iM0Wa8unGj
Mr5SoW/bj9wOKK+4VVss5JlgMusA15jrrcvxFUEr02PvJOgL37VGXPX8hgqrLSEo7yDTp4Q5SaFB
xNQyY8hhMVSGape4IC/1Gmc6WOCvEYb1hO1XD5QE3SaxpAPARZs+9TzMo12bE5fmyWgTBjJ2yrus
hKNAe7u593q90X1bats21gPRSskQundFvSvzpB0B7eJVbbbN4kc2kB+pnYU+agRtVda2rgbZmZEF
losnCo5SobQFkNH+YxuqeEN1OLVlxoqx7sDAICZbjsvHQowcER4sPq7Di7XNmX2t6OMBhu7UXtpY
ho9q5qw2LPMG261xIqW7py9SFem2yTBenJOCHQfJ3k8DPKTH+o62EhsanVTYDqUa3N/pqc4Fhp57
JO7o7XTrG+v+txnOXFjspGXnQQnWGPv0eVbgxCEAJT7UBDkGqOP4FylhtBAwIP1m4YIy8AAPQ9Ys
Ozl4+jbGUbByrRxs5ohiqZ9w9FfEJTS4667vsP1D8UShFCMjlKhOJkTg+xe3r1m2I7WYYguVhpM/
YdSrP4G593KUzq8G9hsW7zkckRLVwFk3A+JbvI9EbTyus/8lVs0mMxiusQZYvfAflHADUfneJ5cp
Insohujiq/rK8TqSvBbdrUpGgi+AqYoFPRkKnZnmlfZUpW4gK8qh0cFTYalyOdNY2FJ0cK7gcAae
/T0oF5gsKe6mqZofjt5vLPA275saYIz4+71gHy8sxO5jZ4PCNbxpob4qGjZprWiap0yEtkLB9KxW
aYN9JtqxfEsUVM1TRUPRAgD3R/l7x6nmAkwc8Nf/gPqBD9W6h2lNEvMfHoRGCLf8eIIDvZY/7yBt
wySydvKq63RUl/t4YrhTOipaWiBeHQdNoYz+DTnwEJJGIlYElf/5iBaS05faQvR6OftglflpWJer
9bgk/tJXI0ZZ3szq+U37mIayHmvjnRCs4T25Qbm5I91++UUoY0ITGbdTu2/R9CAid7EE+9D24lE5
Cbuu3RsZmMvmiKA5iKPzT3LeCVT8kodA6f55lqS1aa7Y/yhPXn1tO2zIDbiOQYiTMz/MGMOXJRLo
eaiCKjR3hXnXPuEsxNeZuGdcTSL7ZaWZG7CXfLfqzs+1/PUP+QkQfnoX7+6LQKB0w9uLUFu1OeqJ
/HT+UqXZRlwZk63w3bkwQfCkU7TaBFlCLKjN7FHV/yD/utqCsou4Mn+5MLLRBAnKVPz+7Sz+jtUn
e3lIo3bjgqIX8TDfb6nO6atOMizvccQxUba/LW3LXv90zJxE5TH2AUOimwmyIP1JSuA95UBeUYgq
XWnI39lgKZeqLZX3DC/NeNZfbTXcjlrqLAX19eGD04FKO1M5vLT02UowT2aeprSAceZfhukRRlvS
UQRfW4idg6NhbTUioEYqXhsdGEbXrKM2pttbzq5hjTqdQXIN7VlUxkSbNCLySajiXK1vnE00Ypyd
eR6stjgUWPmBOF7I2QErc+TIFlSpaghTI4QAqJiEfw0VLpxEkBT7jTOjaZOjcReYcnRIWQB/CjPN
RaJ1YTSb1H6f9HXNztonCrpNeuFg2LAfmg7LQV3p6CUVIN9KqEALHsYlUUTuqKUEMTWRQ7LrBMgD
mBDDgBA+/Cc+4eZwXrGZPKSnmdG7NXqjntNpXLhP9ZWmpCm1ZTmHH1YDkD6V2sjlS7GRtaPy1UCq
8L/s5sJ3YG+DMgsCLZ4cRZ0zbwKNekf0Vp+WAOX3A9OretB1BWkR7jRnXFHtvPWciGb8MqlQB9GG
osOdqERcoYwxFmSF9VwS5NvWjL4uUfhS/59r/0Bkb0ZqJFCib94+msDO/6PRgtqkL1cy2+pcHQnF
8IXcnkyuwVJgTgVxNBHyDWq13sOVRcfAm1CtcagWZfrLAQ/F2KbbOsrFbs6UgIcymcBRIe5sCWzf
Yy/RfqvrTp/3F/GiHYN6DcZjnR/Ou2QIqcyGBiN5SRgbSio7sR2t2InHUZl8fwrCXryU9SdyzRq7
aieGvozATC/BNS6KhG7M2WlNGWjwsBbDXZfFRiTaUWMPCdhxMS31W29CoPazIhQIj5UGAeRI182Q
GILLboFUELIWlufqzVDoFuPZ7k2IVh8Bs9FEaQilsn1NpQgxjLdGoH6jh5RsmaQLtcf+IljrELY3
xkFfoPwBX810Cd2pRcjOYJ6ovy1yQW+tOePCIFQm4q4XeBryN+fd1OerTRcIdMZRkql9/rzbdy3y
buWVaghHrtKXq8hAFw67hMNCsiesuXFtyFjBS+X+A3dFZLAjqCS3YX2ghi3GO4mZyOX5H8IlA7Zh
vRV3Ri85TT1gG6j/xOD4Ny2rRNxLQmGujU2fzLTzuhJfPjDThzfivmYwM+WJThv0gCzv95ZvYRBc
TmjJ3srQ3wMEflFDHv+67cavbarjdgcLRE+0qanh72OLH9VG/Oo7dPZ6HM/XXIy3RLrxivai9E2S
zPQ8Gz6vZavs5dy4139zjiBfaDQT0x2d5Aj4rMS9n0q8YUU/W9QxYczK894I3FdTvovsQuWZ8iy3
n690sxffTQpj8mVK4raKDUkx49/V/H3OY7o6H5vDK/7vcoX1bq/G8RwSl2hjmViOsTLwEuIFGn4v
Hh4EaydD8Nrg85gm16MlIpdrhwXVrUKsAt9gt60bYLG1tu4C/lrU2sJLTkJts0dWPTVoTIjnFrJ4
W4T8UP2zfVJinQhz55wtB3UJpZJ4Ore726jF/4Dgxcee3AVuFJItdPHU78HQMqfriNOqtQOlXEh9
5BUk8g7hyP1xmIXaOxiG7FXIAzyjqHH8DdWByHNj0xayZ3THWv4xSjNzx0LItM6k7cdBPubWhVlM
s8Lz33zW+slsOrUfORp6VQER760cbqd+7fvi3Kp47d285cSJtTJrl/82MomB7/xcZGLQgcy+L8iN
44pRaehP3sWwDKcZQiWC5FBiHbzY1FmaxCbOqBKMNqYu2EWXaeqGpryxrxYIBWJgghJogdbL753C
Gool3mlPlrQEGVyW5gxjvkNFz1qSFm8s5Nxt9ax0x3BW/tlKwyci31IwnYzGPzZdWJY6Jnb96KGt
GCIitEr/He7iQaFPCS9EsEmyEYgTdkpGvDoIM+DTgSbm6GmtKW1jN6WXQ99aRGIQqgnLy6FxTqaB
Oe5y9KsYOaycneymdRQmxwDBO2wHZe3cVoMzKKIKYPt+uWoq9a9Q8S/wVa12+gI7csTSmbiAa1Q3
QEEqve79xOnVefov0ePCGwYKiVln7QQohWQ0qd/IduZZwZCj9sdKMq3PXtNIeSPrLcFa615VIw5u
/5PMBMw8X1ObvCC1ksnfP8y8NTxDKTHsN2h0jk0KbWU8laEh4GUuiTjyqEgZ6Q7MWScuvRRKaN/U
LPzfVjkTA1T7dYb6AeS6vpYfBasedv+FimdkDpFqJIjwXgGXEmsgwb4F1owWZKxPL9gG0+v6TJEx
Xd8dc2orbZaQ7ICUUMsM17EEh+8L7VSFMt3qPk7uESsUG0N5apeowgAH+ZlMm7NvfKjCKsGfJV3W
4JWXyv2uEpiEn8toJhMkA5jgC6eqoEiBQSPhXKocPw4Q6qz0qx4F10/AztLZvCUjGkqqcEnGUbnZ
u76tgw4ipEQOO2JTSTfUZQ9AQTLLkepQI9mPGhO6lIAK/wPXG0tOuM8ZWegS+v/mC8rr4kaS+KRH
T0+FomE9FM+jUVbdnd151hk9vEGRpXLMOQb8a/Xa196wy0rY/wsZrPBfTCBEGScE+QbhhxZSH0s9
RmB28XU/n6aEPPUFfKl/3ecWIHh9iSc44CVHAzQ9sO13Zr4jqzmHFPeHXiihnZB7ESThzmyHF/d1
PWrqvUvpZAXvdktfQyebdkPW6QVqePIgZ8NC+SyMsLLAVifv8XDDI3XL+lQRPQwOWy56bJOfskZ4
hLJX/jRDYBb18eKAMDuYhCA4ioo/49uBQH14xfYbArX5P12yS1kmfV4EUrdXN0Nc50e2+mODqXZI
jri65A2R9hFgLxXuV3TYNqR5aUNWEl65X1MNz9mFTgLS/D4ovaLUxoq/CWnXEux/pbM30TBGZFK0
SYTMY13eKNxrTjoPeO09iyhdwJph0VUjVGl0gBphAoD0d6SCqTVEYC2CA+544MKI04iwglLlngwj
jX8E8T3aRKm/HFZ4lgwc4Dbshpl3SiLHzrlIP18/GZlnN9iuBzu5F320gQLI9v91Cb14SBuXdFX8
W8p+mA+BC8kXFSge2ZD2+YqCRRvvWq0I46xRP5ltmgQ7bhrMs+/uh4i2zlpjSNNEq5KgWa+zY2mE
XZ2T0bDvyYnKTfdWKG8gX79RFfxeEzBUwo32qADjccyxRe+IW31AEXZvP82L7gK3pLj2Da2e+JIC
bN8y0KHYoc+nXKM9gxNexOGtR4uS8CetFF0Aekh2uJhwXg9x4WamceB7bKz8BfNJL5poHjzYsZFc
wkpHT9Q0GcJVkaPehE1gP9JoJLk67g6HEzkg7tLAyPmNwSpqny8iCSGdbmfCGH/EpO2Kx/xA+69L
1OsG8ozfbok/3mzgnZNKVD70j+nd02uN6Jyrgmk+UKWdU8lihJoGcKzTAdDbZgEij4Vy4+cDCBBC
s4PubIUsPCHE9N9YJoNk3vZFKft5CAZIkDjqNUCdW7zkmt+5sGDbKO4+vDawwJDWfWGdGeeekvsT
fm8SLqjuuzBs5y/MZfapQkAP+RUSOAyihDGtzuhneLj3O5tzhsA54Maha9V8UxtxqSkElk3HF+G5
kXJDAy4bcOJ5FTghiJlwdQrMIuZhokNZcAY0MzbOv9ssMDgE4PnWG2EHdSrg72Rkz0CuEyi30Fjp
7wPDXDdcp7g8+jwnAXHUWDrQtQVAwh5/CR1DCKrTkSK+BklNhOleFD3ij4Nu7jOacN2IAJ8FFjna
tVMY8h0KhpASxqTWgIqBqh1RwYgPG7NeoMSlOEKAJmDXZRRBzPeij7Q4nlMDqPum2wJWwMzNRyVi
ea+fpMLKzuo644z4dKkRsI+JB5N5806FlrqUlht4HtCprVIO/jN+TmGaVdI1MkVeeFba7mG0fYlO
rlH7sLNDXVlS/KhNcsJOxK888bpyPZUMjM1afEJVQh/C37t1VZ7ssRk3aWEbB5wD9NO8LP6HQW9p
5Zy7pU7Jt3Y9t8H7bcXMjO6/kgeNLmd6dRyZ5UHtMVjDKwbYGIC+ZL1806ZHxNGK1U/1cZtObPYd
BZNZ3Ys2tgqLTGXbnrYNrsALFrnhIsVfOyk4fPPaf9wg28WMBhfqX7/1THiGy1zGPXE/GdGBKi2d
pZqD8yQICsNXj+I3y+X5ZygqF172XfY5S76OpOsuXCA3B7xVu7GLV3hK+7H5GpZznvhyHgUtxmK/
89EtPr5m5MJ16Z5YTs4763lio7dI7hT3JEhGe2iAQfNrSCbUdl+TmuRZBHsZ3g2ut09TbZc5WZcO
jUernTiTObFIqzDAu7H5LfqUpnWzc467PPv316l4w99ZOFTF9UL87jWiuItIqLDNTjUwX2u/sJxv
LksqIGxc8K9J+Dc5cDf5OZS64Pznc64Q5KAZ8pBAF+1vWebfovjf56sqhGAoQlTWX/GeKahALVfV
kwga6kbQC51UmRSD+XC0Skwfm2K/KqoCHcku8GoGUkXj3qUQi7hYftIHXV/dXC2r4oYnEGDqOB+0
JWetBSGBz/7K/mFhZgiKV7cPNxfh8jY2hNu4eDGoeZJ5n1LHgQIqpM4I7vxskGGnUOTs28rNGUMb
fpvwulJp4GtAaw+0lgIwwq2kVVtBQ3inHzLs5/UWRKjpM5p8ZslxpmDdc93YV9mJm8mMTHmUYaDS
Kj8xAoUnxwwHcapUK9Emrm0eIz1t00KKDs6FRDs7EONHC4zdPg/FmgkQJhgyQzhtAz2GSM6V/BLn
bvTgrIWXqY/98SDkqjN572mI2u+gOHqrI9s5IGOuwza9eCCXHwtOwPL19Yk0SGAOrDSpv9ECrw41
UxhUwhGJU/SeeZaKxEtHHw3wRnq5IlrVsJcoTNekZtUD5LCsVEfaVohZenJoiO+NObze69hC6gTa
pd+fMwN70AfV5JWXO1AqaMXKvbdaqF/VZzJ0e/G9VhbOEfLFdzsf8ttJb6xkL5R+4lKI0K72cWob
LoyYyrPTsfuajx0uLE8gT7Ca9plUJFdfXtOY+DJKVeew9HcvHrCz/w3NZlu8oOuczJ0F4+odSFI1
NBpdvrVtGY8EmSyPu6Dbm+v5gKG4+W2RwTrjJVbwa3xaMPuZPP/0wyaUrtPZtkq+n4FMTmooqp6B
nF3BKtLnayNM90kbVPaMqAe7h49ViLbnYJKmOy8zq2Nw/MOAvOtAn0dO/lcWc6+CKVEx9K5xjlNL
/iwVCdQugoZ1WzffVvpfxxlQgm5JuSvMUyb8HCZ/uijPfd23GEJNM8+1JftvZBauHvFwudGaGBwa
7Kfjurn2M0SOE9JLuIJIvsfaNF+nTFy7SRjc/uCCFcIdcSNaSV9L2tjlv4LebyC15twYpxnWP3T+
DV8k+XQMgSlvIQCQTzjxM6KCce2HIRVGzc6XH8KcMS04VYU48I8Im//pq9H10z9lfOLi0MabeFSV
ZSAbdjNalhj0E1q8B+vdItmur4xJZ3kA0YzDguWjYARTcpUt9/up5+u/myy1JJBsScv/BHNcs5ZY
/l0KO2lcr6hu4cqi9Ok+koCAxWy7g/rR/gHOk58+1anv86uYeMYIiv708UnNKqTsep16jPzymUK3
EJely9traCbZqb3cobXuhnppoFwJ8sJsACRT5Bj8Q/toTXIBGFTDAmP9VcpIOfZrcIh7FoHpmQGo
ZvcpLlIlh6kJLsqR0TQfvuEwY2isdFVa0bE0cQ6jb4DgQfmnNvtbVwATmhC8J0hm+CpY7UM0Ubqc
urO3ZcgNiclAavvJQzS8umSQXoQk1dctjVCnO4XEpCgRmhEJb48Jge7gweHoxs5uQREbNfH2M0zz
qurNZHHdoP5SphRTxguD8d9zfqX6s5tj4iAfLjJnr3LKQRBHnHB0jGNLfMdCjf7Aqvph6VM/4oma
oa02i/jBfDh6JDq/vM8RvHJzqk3fvUhUt8BQHRZcfYQD1DWHG++TE7K7rS1gFwIpENiLzQ4twved
91MBck8NXz4QlSh0Dq2181fDF536bAseUXzqzV26pVc0GLAi95LjV5x9SKzvklx6ftrrofFdT0UI
fxnSaKjcYfOjYBETY/1n+RWsGVQMgpTwck7DOUdjNp8dO69feoZjj/lbNX0aQghF3wIqaMhF59Xx
atGIVhBT3/NLTeErFZOYqvXeRmcmOkPdVIpkXdEMn7ldrm1AApq9T6PlQmjcgBL5q/hoyVvEmlbK
WF299kO+hyOMhYwUgSlJ2ZEg79Q/KBbddgC8ALVOWuAVLCuIAdZtJ/pPZcJK/H+vkjnjfz+GoVPH
9W4x1kPhFu8q+zDLVCOdPWEWnbd+mOdWsqmp8/KvbQekzxOLm97yTqsgElNh2oY3AvXmvt1noUQV
Tca/ciZu3U1FvHIxrpiMaI87nNqoqi9Z9veUnnXf2T7eKbgIGHBTtEw46FmLizw1wpBPxkHecBms
7N9fNFTMxRDSBnYFHM8Nx0Ltp++Jkn2/1Iq+0t/afNsf0thBqTgyyRao1kRhLJAfxyoFpHV6h6fS
7GiDfAZPt3MTTVGlKBDO5nYX4K2pYFxWuEVihA7AK4gM3854Tjwru1iJrJU5hmgNY+bmZ2elGvQ8
CLcB+bvxX4UwBo0ISg6iG9aM18hOdELAeb38zpC8NtoZMs39HGnKVR1v9iHdbEowHujQKD1kiCEG
OhwvQ4/ZI03aF/FlMX8M0mzl0uc7AvyVEajm7VzhXaU9VkknxFwRYLaV5DMpM5LBcL96L5qPj13k
K4HGDrEM/lS704vbQaO5gX4xAGqPThMc/EqPDvWl54PlYN/lWctgBU4KMbP3j05OUW68Ca3XIoM1
Sg/PMNI6/cKMIIyPTpjSik3AQ6/7aLAxfolhZHAGM4BCTRNbVLDDSqJ1Y/F4AWsUQLi+ekjfo6bc
IuKedLOjCDiwQgOcbwiEQJuaM7FC37XYTyKyPRqoYVJT9fPIYXcq6UeQY3q5ntLwDBniHiYfnSsS
/+yN7/lq7Zr8GdFEz6ZAbaQZ9XaM5txo7SdlwPm6uKOTWU9REXt2kOB1lEcU25xs2SH8b0QXNYhN
WIvwCWwJIYady91tkn8pVR2nNXyj5699FUuM6+19jUG2cKF2YjX6V10QxAWtbNiKVjvWMTbZdYrP
UpNK18Ih6TJXKP5ywML9pVaK6CWkJyaeXtOUarBk4zsWPjUC341dOrSZJJL071z8reKUjv3yrNey
SBQqFtmSVVHpBqkK/FE3wFNG4cfLymf8IcjTQMeV3SURPXN700JxJRYpErQbb/Udvq6TkontLs8i
TEzlJJ4grutc6VlnHLJ2PPMD4X3nhxYy3IXIK/FDLrUYkfOEavf4SdEM5DmdEFvlEgTHtwW5N3P0
bNolthVf1U5VTFftlRd49NJesenZHYoXZ4X8unyvMhOnb4Sw7gAlmeJbJXEqXhrVq1g1qUFw2LSG
+cRqEC6T9rGkjWz6p/RdBeIhjg71DIl8sPO9nY2eHvbT//t1sO6Hn7SY1xgXgFhBF0MdxXgErAP1
8bZNDnezMxXcPE9sq4YHpHbqbJlFV2LPflSf+2+Gsx+aFTRFHICmmj0miCF18+RVY7or6Ey1z7eU
b2MklaavyrdQdlOAYBqtqL84PeKIHUup7A8jvAMzwcpPkk1u9tb9gzAuEaGV602p/itBU5EH4Ooj
TO5mAxdE7QsMeacMbc4UQyH2dGIIaldstYBobe35DgiNgY7z5xf8v0HH3v/k0XgLda/AByCQUgvP
uZg/h6kyzbMqxyJKiT4ZNvjAvTvT5oMrHaGv6gfS0McNc0ZH/x+shrRcMPANAwPqMDXNT/W7QVUx
DZQ2zq+N0VgBL3FXwe/nS+C5/EIn1/ej/oo+TcE+ZPeJ0ubseTF6c5HXa8YkDoJ8xKAjDxNIR8Sz
kG+qvpkQKtG7BR7NlU+JOG0PYvHhCpKvo9Kg2uVC/Vym3kw8TguctODxvl1hX7kWP+iXGUj8Tc8O
M58aXhZFFi5CN2uGaAZu0DQOBtPi7ZC+qxqpxWW2508Q+F6gLbRM2QlihNT/NdNrFte9h+rddDpc
iCOIgjGYgpwv9YQ38RX2mkyi8mN8s4sihUrKYxrlbWWWFDPc4OR8+FmxWoJK8L1LuHL/AgZBJcth
9lrXkz5NFlqXhYIEk3A6ObwAzK/C7+xJBkm8Eij3bZigjUqwgzthleBcJuxZ1yLNqnxiPsWh7Lh/
A7xwm+4FGMI4J7DIGMYxaDoENySNWq63ekPi1+7GcxVm9TQECen3ICuDcCDFH8htqqBqoHeKWKJf
Wlfcf1d8CpV4qynzMKid39qU+cZFVzA3Zu1991sp5Ciq9X3qNf/1LSO+4nXg2iEJwuhaFurxBSX3
4h88dI3ogJl+I6PCcI40VN1WycrUbmZ4W6Z/cWBZ/8U4mms9SocvibsHwGP+bhiEE5VeDifFEa6S
RgiUSPKLwsA1S5ZOgQ9ripKMPP0r9pstgrRte0o4sudR0RHSGz1o2NsOtUwAsBsTm24NkNKOQW3n
ZytRw0MQDFuFgrjXfsQophJX81vO7w7D3gYZMd4MtiRP4Ho8EdMt4beRUtFd97kqz/+/cjO58V0E
sYYTGlVSl4pv2xhHF9Jyw+4D/zpZ01c1MBuGipyd9cxRnR6gaJ9L9nC9q9+61TRTz0wftidDyUvY
jWPVf5kLiewCR7Z/r+yAwbDZc4nkdxUeChgL1r43BqlY6jC1ZqtdtOM8xPqy+i0FxN7DfhhEO45X
gZzZBJ4Gwn719PxRym82K//m/G/WFdqNrWJud9sOuxNinME4aXGV6hN3DlxDeYK1JDjxmJrmwlP6
WxaqCB/BZg+r3gGlLp2kuH15bZz+FHsvrbiGvcEQ6ggDgZtEmNMaYKSbS+Dxvf04xZ9jngkD5D33
bnZkYiH7wK0Iaqg6MPxV0/sEZoOtXXhwjOL6HhCg+1HbUiliGSvVv1x5L7iyJljUfKTHc2qTk/wb
oqgNNi5c+77g8V0lX9Braw+ulUR9iH4Qnpob4sXoVqv5YcikIvixAYKMZVLu9hCWR8iu3ijtXOgU
ZblarBAO0neJvd+9JvS1XOVFSeLrJacVl8rBFaEWjKra8LdcgUTxzNcECrvvtD0nh1/fAM7cH1Iz
ihyaNmeDjb2L8SXDJAXXznHwkYN+g2SBtHyJQLtREmWmBwyOg0zgAYIbIM2Z7IpyzhIafha5b6Bu
f62bCbxoQcKGOTb+FFRLIG2GXeJQmUfUpuTDaOZc8/vOP4FIY741lkHOBNF5/5pXdl82oNoTxVcs
vLCStTMIXguYwNtcJdpkS+l0+PNhmhfM8LimB/OlvIhH3WB3thazcLcXPH0gEfWkOAk+NvugqyxQ
WEudBm6zROz1YqvJ+4VFWSIW7jau9UjId1NTkj3XTFBZy+lcwxsnxI9KUHupW0HQNHYW1t2UKy5S
uiH+4ilwdI69Wz5+G/PNaKIMJz5KUBa+VX7Fr7zyXC8HJGoLQVVkAhy5LzrB0XoCOqGyKW4wGRiq
+aM5IjedjyUY85FRBCq+plX6yPu6HF1B8/Tkng5wjdJlEyy/iZDWUymOyKHFsW2Dd7Vg7N0wRw0F
FYvsDk4UtbDC+snw4zDWG8hlItXh+REGSsaZ/NDo4vHLsbhy+FYxl56/+V7fzlsPZ8U6hbteV+Ce
ps+vVE/Auy5D98dAAfnlWFJXDz6Gf6P0wNiQiOu05vmmKvx+kWAWOv6njvDzCAQZZssivI0LPOY4
67XXfUvZPlfUYf5xKofpHO5iaBWpuJcXv6YaAv9uxfKY6tF57u1wDu/UXjhi8fSgsQrmBvCJ5O+Z
qmpdyIeTGOb/Y55BExxJHpCIXhS0jcUMFQP/MuQePFrMACExBL9tuW79HiHbEJzhYcDqr+Qg5VwJ
ILeZkUMXWkujcdVznGw+PR/NxP9Vs72rXBYN3craR9mCNTTdgOxou2+uY+O7MDKAp/XP4GLcZ/RN
kviTCCwTOQLwDyiSK68kgG7FSToZ0a95rHOBn8o+zVcRZQdVrzJiBMqopxtw/FIpafpvRD0SkZAs
GLbs/zxUu8gguaH5n173zZlwTxk+UXtBCOcFxUi4gHBLZYqb3EdTc2hXj67HAI1ErLDYCniIJBbO
6FBMXnYtHWc7GRdsURTpbOLScjvjwpGOYY8S5LVctVGQQpc4rX/yVqX9jvlEOxJ/FmclNSgavm5R
0ZqB1E80VC2XV4sRIryLWcXyXqAEm6qwAiQpR+uAJ1S8y4cS4ryg7qeM95Xp/W3Cft/15ZWC9Lzz
fPRFNoIH+PL/MkEcy1sGrapiGtL97dr37K+mIwxIKBte/5L9ODQTU7awq1cVsiJL6HfdUd19XkM6
ge78DA7+VWMCOdTbQgElamzBzB8EmeNARPIJc9KhKDTeghzixb/0GEbvJPwErpkpfHtSwyF4iFco
C3xaKQ8lwBqgRJ3dsgiNjRIqhSWSLFGH+jX1pZjkhfu1TTOuq8VGq73jdsJou/U+SxyHQ7H4aUrP
jf/1P5G1/sbpPfsekINz0ykMCE1bsqYiCJHgviLLU2CisgXbnE3YYmpDzDPUVB0cThu1XjVzTCzG
hpbL8icP/Fqkx2a/Zc3oA8rL3tngbPvS7/N4KApNo5OGsbxybUOiEfB338fnoa9BG5lW4V+MJ67Z
Zc6uldqfxbDQOZWGgFn6NV6Byl3NVRFHxA9nd8rEA13lQB9vD84FSOT6XwOiKOvlIhm4bnuZm9tV
KIOD/6gC4yICI8qnPOvzJcBuGzeN1r0iXY4klHlwMrTnEf6+5tTWU6PVMEcWHIUx3QWQyuGXqLQX
SCFj4yysqiflKa66B5qmyvci1kU/rqrPoAa0+8IXdxh4+Wnc1PqLa7M7QoSWx/8fbiaAZoY+cp9N
bOaEvhsCksSCxKKyTqrJ3D3IwZZzoL+hUCOAlxuwrjvBUHxEXkvtJZBCq2RyKq/3KbWDwg2lzJhz
PWQy0hpXab5suYErmNHa8ITkr4EmRioo7XQWO7zzke99sbT/wg1vkxTMThqKNItcXZ2piw1d7rfD
chsU+xoudo7yCfNbpcpT8/oPBFpsUwtRdTJCHT+bFJpUG60Knz/8QsR0rw0MPkr4hAEWd6Iuwa2d
CG2+1pfKKlpSZazVB5p2nvM9T646Sl20adSgdj8q7nd1sSMVJiN35C9xpi5derrfsoJ4IQ1BmJoy
KNRzdjj48zfXt1IKpki53c5uDh1Z+9xJOPr9DwGjlU4JckkIjqWiyL/bgC6RVYZALP3OmvBrS4VU
TbfaGkr3U9ysYyJwe2Vk2uGMQNI7fDiQzZvuhBOqlOau3qBtOEAcSi7hQFMeloKW+mO2gsOfEiah
v53gY5RrZ/+KNGEM0f5trA6XjOD3lbAVjM+jM7NvduZ+JQef2V0q5tMbrOsX+QWbh1ITWQ8hSwsS
P6jajlgv4MKRH7Q2yh30G0i8PM+gjUElqmbxTHgkXv9AYnmqUybTxfDv8zsy7G/2Ni6im16knr+x
iJjw7U8AjjfE5d+nSnPeGGwKl8aZRlcf0kMjq6GkRcG6Hu1G0QwXZHXpRbvy3xxVarouSoXcK3re
68GAVU/8x4JS21yIOrz0Hb9POu8aBAMi4yO0xshL6XfpPb5XjJiz4MyWf86BM78mzQTL3FFHifVp
LGoZ957uFHUCTfmNsNDLJ6Dr1p7GddDoJS0SJHT0sjyi29EA9naOGC0OpBLdvxR8H58xYRPs/Smx
MaMoe8VqDu/scli50ycDDfO4nUVyC6htkkdd1HaIrRDJUSDqboiDTudGC0OwoGYYMoX9uA+1KHiD
suEJg10ZdLOdxsTB8FxMXpch6oWUa4hOIH4UI5XIM55YpdBJbAvsAfEa+ie4AP2iZ+KIZJWbYgCJ
uUsGd2936N5Qb9kCMYaT+Ldwh49rv+RTpd7CH2HLywYij00OYUBJzHL97QZb/Pg3z7EikklEB8ap
iy4s2+V8iZ4UnrjbXRRXeCl6Ab+jzTXb7iwEROvmu9spaooB/YPpGMFIsoIhay/73Gx6CLj8xKI6
KErnNWyRhDXZoxdwX2Jed2h2YEc6Rn2g4YIzMEoTiu974vP8y5JYrTkOGxPD3b50tALc5VLa4hb6
QWXrSKm2Tw45mXGf5lx0bv785auhtaS+H7LZ33STgSYfKyrZTx1HkVgv8yWhkF77WR+oWWiswEHs
skkI0b/4qcMmO8P+YuYlYMxrm2xZuWNIQxf4DyVTZw3x09fYRJY/3oH8pG/qNMLysaV56LY3fp9m
I+Ejkskt7V/sstU1AUveLNAJ2sCRhMTUfTOEBSMWDTE1Y0necLX6pVPbYG9+4yl3/QtG5VSP00Ob
TE7+fClXKKPt5xEuVUxhNRmEgkbMLETvH0IpPJkA8XpgeUAZ4JutfVeaBEBCLP6SPCI0gpKQ6bGE
EaTSg2P0Mgxz6glteNaswcfHm7Wv8eYGv8d7uVH6CjkrH4nhvK0iwAjmLrm0lvgwUhCUUyG253F3
xOSJphdUv5foQUZkpeeA+T+ZeeQ3W0kH4ejJRKcL4kdvq6SKckUrFnkYeU5s7l1QU/kM8CGYnuK2
rJKG0FdZH3gzmM+sv/MqczXq0LqqOqWhT2cV6sTezYXznt9w5J/49QV22XiRHEXnAoGi8sIHnAmc
wk9WvJWG00ydgaq8EjOgk2e59/kGEe8PrmS+j0lQSj1B2GPO0a/Idadq5lhIWfLpkQlR/AdVAM66
dmgggbGp1BcCKq8qbPbZ/UX2n3jGBGhxAPbSAy1hE3ZuDI79kigtfJurwOs/lomWTNZWevlQjp/B
HHX5t2+Xrq2U+f+J+4ZniFYJpxq4WPOVHzocKfSlA2kSNL8qgTJP6VdA1AgG8YHgsn0Xz0Pxts2G
Gt3vCBlmA/qWqQpxeHaOQZpyHMUAHDh1glCBhxqNn7RoizbgVJgHNXKGI2FIpbJpAnBhspINNAdw
Ey/HZYWO0pDfyjiERlBgI1al5l+JIhd/pKc7Z887xyJQVBZnroiBVGxdBqivZxMBoyeSH1LM9uPC
aJK9y3zbjDTPnXgxWepWSekHWLWTU7B5pqoRg8IFS4UXbK/CFh1dXxTXP8S32ouDuZABCHRy2Ql6
ZT0Bu3saDQLa3tJBCuVfaL0PwlJiheYmjThhZ65dk1fRG6ta56FVM74ABYAFwM8as2yl250AA9lA
plT9IrZjfQlXDBmKSz3VaRijRHCfdd2/iKb7mvYB4IfwHrEH9mvKjADfPX9JRCExhkS+oabE7OwW
zdpXEu9slSOtnwbWeTm0piv+6hacemSH8kAn7JLP2rTIoJkMkHoydqyIVQ5Mbh6052PVtJqd0LnR
c3P2RY5Flzq83ru/bEpqw2ahhy8aZ9wt6A8a1FyArgymgrSy7QuJunvHKIP11mCSyFLb8GCJAFRH
rZacq6jCaWBJVB00ZgXNGfEG0w96zZmjiTk6wYLLcwq18mwTX2ArXOhrHxGMMvWXF2O+u1oYfypI
d7yDQUkdc2wc3TorIhFSKgc68HzNg9z91Kng1AYlmhJFY0TawWId/VcIygeqcF1HcswSTun5kjmI
gx9vmAeoD77/5PoZ2YfUXuZBfiI7Hj7jsAcJDLODt4Aao7N913Cqcm1uMPpqxcVmJGD0zDhfwU2S
9KKY8nm0ZLeFf3iDbsSXCz/3ooUbI6jrtTe5g31R01Dfzx3LEpgs3g/kFzWgSpy9wRw/LWhQ0Lt/
0MbdnHybAIp3b3FgtbKbQMIMKQT2DvtaOhidkZZ4BvZLlub7N4RQCF+sRU0YUn+Dik+FphpdchxB
r1phNvNgQ402Eu29I2a8z4LRSCFyqqAE6JkAP9LoxVsrqbEWEBquSol6GpgpWz+D4eSY63pUO0JZ
AtQmlQUgXLDIyONSw/mKWUE/CDjAkNBE9tqnVWCLKcxAae+Zk0Gz7Qy7Jcfn8Oqwfzqq4YramD/w
kViKpqvBKiWi5wlsiqhHH696yMKThYZFVW2EVQM/oEPa1SQVWZDmsCpv/RdRCfi1Qo/817LekAsK
KcWcSNnarpXBnInbBLx4lYDYsCm/t4LBq777NxV2Nk9XOHpc39pqF+PwDpDxGnwr6Vq26nN8MNUq
RyBJUeZC2kwQ7s8VliQdRCeIFcC9vRWecFjtcrni61nR1O1721mIkIfksG0ortUj8rtz1j/+BA66
XGwdCbS/lEqoaXopfWy8dxjVkbGSdQb7A83x01/PDXtxcKhlEbS/h92pmaw3SHnyc7ARUBydG3Y6
WgCUozbcur286QpscNlGz6P5aufcCpDHPVCHgWmFz35r+FV5yvYWJOkIck/3qQNDF4TEhj7LJt8Z
ssSm9TAluJCOw36psIFcgioIOTWT3sxChsdVivpSj9dIjOL0Kkib/HrdqX0Dc/XMhGvZEgiHw/M7
6V9a4xyLBuR/qOBkb17AW/QtUkPjnbykMex4BSmkiawhylIlYss4hdmrsUkkH+qWxg2pQPajy84Y
hMZ/mmuxQgz7BWjNznoFn06DIuqEcd6/F2GSOh/Y20iQyMdyGFr/ETS2wQCFS4YwnFCI511uUFtV
6S+2bNoR6UOawOu6Phy/Vdl0KyFj1MTrBGF/rXVLhBOf+rl0O6Jov2NITYHGc9MbGl0xMiphnJPu
AFkZ2i4lTHHMcsjUC9J+RZ1PQEM4pLTZglfcZpceF+hVUnKk+wKnIqHteR1V4xQphdsriqV38Qvj
bEVs21UIm6KWezNm+S40Osn4QlO6lshxRcH7v4y1+tcZKXwUN82d6e6+1dDEZqXstVCME5IBjwaa
ToabBPS/lz0ESdzq1VqwXyvD6SEzdgl7bKVTOYgp4DVIpVaKe+9s6kRFPTzcWqy2jt4LWxS0MQmv
TX6WPTIEkJa59IeCBLqhJ5FyRqgSdEe7OTU1teWBiLsbo70y9lr8omuOZ8nq/08jAhOgiCJlU9uU
jfa86OnKpfAoDjOQaYsqKdm8TXhy+3Ac8WqrYza8G6qhF8bMzeCoKwlKjUpVA3SHs3qEMcEj8P7g
M9KIM+ea9zg0E3uksLqhMOqXdRN3Q+AfiyIxyvRlQcFIcetrEe5DCi2pFSolkelslmemK9tnqDu0
rnfl512PTqUW4cAsa/WEIIub/O/Znr/p/m1NY1+I7tqA7zbxGi1qOaKLYmCpzCtMNKuMN8A4+Qn7
tEJTB1mqLXu/ekgGO9oUKapGj0/qiF2yCntaIJKmkqaco8W5agfCTODehCF0Ks7DF6iYZ6u2GlxB
RRgDN9EzhlGDC2t7ytzZhsuWIDVQIb0hgbDUi/Q6sCx2p2n2nVCiYBDIb6VY4HvqfXlYm7XmijDp
mg62Sb/kJvsLKuJW695RRDouVxdn6D6wDEThcfVK8vhdbl5Gr2fGgzA5XX7B3Fk+tRWttuQO8tRe
Wi8tk7nYsLy7PVjEqEeb8FGBGr0dLvPh1cyibASh3LwyQf8n+f36ZaZcIWUJeSLwvxQa+0rM8oUQ
FISHzFt1XLHX2gOQeKOG0i8p5Rlg14oFrw506RMwO4MkovmCTka1zLXooPjKe9tZgTSK994RKR/5
TDWAcL1f4zm+rbPYuYmT+QUPZQuv2CdGJ4apEnMRJC4bld+V6kEGXW2QQ/7ANOWWKrValvj9ld8L
jd8U393YM4o4YbO7lJZOkkPnnFmUKpt65Rcmp+22NTMptJdF6mWBDrfjopCTDBLD+19guwxG4nRG
xU2yJA5a5HquOAqe0wtwJl0y4DAwTAYmJD+gUHIzLGZVBYSIXxB9U4QqtP6NNneszbOKXdUPTQrY
oXb0PxNHue4BDu1Fbf72RlFmlKeuQpn7lgqIFoIvvpNelcs8Kjm5uRBX/edrRQscrT8J6Yn1gqaZ
CTRWwKQue8TmaukwXQjIPuGBqukoXyaKaXkp7symmO8yWbJeaJxNNWXdIXwT02yru9Bxi3zlpR9i
SQRU3a2KHp79axcH6+QvRc1+DjGUhOpuLYqRbskGPfyHbfCCSQstPtfTNOGB/J6FdEwn3j+Q3Bik
dYTT2wYS1j7BP5bsEhGnQNXm10K5XS6fQ6J4Vvb/SdKmVEUdYJpQ6R+j0VDBAQV/bTbSbj+tflWY
JGvq+yVmSnuUbGDte3Z9DfIESOUQGWvI+EfLqXTa4BMby0vXZf9Q5U+jqw2Tsye1K0cNeWh5CJdM
D9W8dU1D9P0KuCggHnOF99XkL5wUsPt+ezhdcEyXdBFSSyiFqd075J9/R3dTUm41DAi5M2Kmrq45
DexjfTJKP6UD28X026wLj8/Wjs65uOryDUPm0SRhI6R1lhxpO4utvcTu96LwGs2Cu+IM0K+lM1BT
Pq12+BdJqVsc6kG3cYJyKkm1yBsDABfDVZayKCzufkb+iSVE0vxKfrJtWkvZBOc9bvx5k383qcRv
RNgc4TSr3bfdHCKfNoDERJ9NBMjTj9pXQmJ9CK8DBmy/urf68UvaezYzcPinznh2Db9ZLSj9tG6V
0tlojJ85q1xKJ92Y0mT88e2cMXwM+l+R/jW3u+VlxMOBZdY7duXd8xuS5MxMeCk6dy53e+zj8qrY
9k3T8i/7eQ+LLUq6Z1aqOaz2p/ct/q9SEfMOMw5D3uKTqtKcjrjk7ssi9TfqpYgYl9XA9W5WlLUs
cd0kvsqbnIphkpZV1g8IaUuX1xp3LCEP4Rt141GsuNgJ0ZPWY4DITbHjpXriepm8PvgW5RHzOKfH
GDmAHzfbUlgAkCJDPfR8V4rQU4H7Gciswli3nwi8ixfatdYrQOFXiYXRfPf8h/5GuX81GjS8P/uI
uLO0Jkfr605MH1ZO/e6IQZoIGHrR0F7IHuMxiowHoJX3dS19g+1owRWCTT0WxznyZPx2eVrwsGNs
mcrUKx6emj3ekyVBgZLhVIjS32AFLwZhbwXUfftyZB8V6KaKzsGNR+KZRUVnzp4nByeBT82Mm2J+
F1OrXccKeZVVnhQmVhI9hL+p0VWonVbCwnkmAhJ9/oqlknoCV4ubZKXlAThPiX3tIDB7I4kv3ngP
YWfXkVzvYEel+h6hxOup+Tq3+UazsAu+WNPpKM5rq2mVTQ8cfYAN3QCjonK0MBBhykuzJA3KmCSU
hX0kRIbz6p2UGwj/X9yk/21KgbhjmvvGDqw14ZiUeGKEExtjWJZYsnP/7Ppj1mBqqCJ92DRIMu6u
yKGmXaHpchYs1G2joWccFlt4whIqLqFV8RCOWqPmtbQSV0xWSqnhfLAtlEc7+hBJbnREi8g2cI5F
VvOhbf5Pn/lSQFP+68//pM11VArmkHjUDwANxuu2bmY1s0dgBdJlKN/xJXt+ZQJaAzzW+ipuGqU8
VdeBDATpbHrOtYJdWp5oBERIziOL6/cExe2TBds7b/9pjOk1AtSs/epljeTSxJqHjwAtEPwcF9nD
IUT+FU6m2jmGxqSoKsKZhe0MAHnFfDXG3l9vmu9bpkxly8Gi1qw7IMRh8BPdaFrZ3xw0oUVVCFpD
oYi6Vp0eS10jVZNpl2TmmxB2V+TeE4J8nw3OZT8v1eYlIiTDxZlcc2pIgxO9vOCgbkJHJavll4aF
kRbwEvC504x4tCVl5pjrr/r9bVB3pDsnVIeRIkkOtRwApPvw+qngiLT2YXuSFgl/4l1nU+i7D8qI
r9cbjptzlfYleRCtcWsecrq7XO6htNkqdA4qvkkqVU5AjNQMIZftCn5nKBYN44FSYBE15XCQDcB7
pVt7eDulZ2/HaqyQL8bNcGO7JAokcmif+YnX8ID1VtDDux/B/HtwabndZMcekRCW2BGWejKLKbWd
/nucClnE0Ku2rzKdZHUesWAG/YpE9HMpjba51elU/Uaj/r+X715C4xLzLEjotD2DeWFrVogMAaYD
P0sp99kFwdSESioioiLBirDdymaGLjy9yPqmlwp0zYpesvWChH8rkztzYQ/gQhuJxTFgZuE9Izmr
KlM73y1q1OghCSE3YfSRXWJeKPi0cdk6AHJwcfd//YM/iDPNmGDS8PJomg4qCpdkOB+FjsbgHkaA
UDZpbwZwAa1fpJfF3dx3RPhbBcyOKzwrjD6tKbtxLAbG2sAFpTUwmNA4VQ36G617dCKodhOXCjCE
g2VTXMFvYhoT+pMT4xD06tCcxBdSA6rQODqnVareLAByfoub0zZeWF7aGzBd1gGHQVAKTEmuinRD
uY3EJIIlwPTKjH0V5sEVS9OXal7RyC774UGSSkb1rr767e2hoWWGdVkph2q2wKSU8lGypLHCtDEj
BBJPW3aaSSLM95BB7YEULHoLVvzLhNbLTvObZIxF25ryeSrhPgS7hlZbhxRY2+iEZCEVsg8SDZsE
Nd7Xlzc5rKrMUY4Xhvz9hlSXF00VG+LMYqRmcwWIcFmAwqHkkCuSbo7tAxwjFYuks8Q5zR0A/7ud
saCTN6/EZHDJDLaC7TVSobduBUtE5l+NpfVckApPgU1q9h8bwunS5325b9YCSK9XPWL3YB8Zf2ur
g4PvJJJsWlXvfNPx8f+V5vMvWtytN9wn6QoPs3WXzBHPqLSyo5HjxyfUfT8dEKa4Zy9MfCrIBmPa
5F/LzFR0Qh5H4nJNT+BRMeR9dSSE36uRptZNHGSYxCYnIQpc/bN5+q7h8GNzZ+QnONRF7ln4POAI
I2xY6WYfEeZrrrEvDDtH/syHUJmK2HLtPUGTSXLJI/S1AC+dpQ8TGd+jHmKBfZjeEBtxKd0xbWPD
yabqYScK0FqQgE5m7VKwdtWQ3/5QyXRf6pWqnS8Qrm8jFTrucNWlTjqLObwQ7TEBDv+EHFN3esWz
PBLQcXW5w9ZuJ0P1ouDNxmicBXhf3e/SpJPnK6/CiY2rMutyZUcFKMzCXXSmXViBu3eFKPVXlKHb
4TxWNAnf0BngcfjDcI76XdPbMF2tFqwxcOBgYZgVSwgB7ON7DHrdBxpW5vk0AyyT3kHlLY8h1M3k
SmObcEbpPiIg6BoZ8vLoxhErYo/pbBvSKlDAdGFheipYSKvd36TS2b+ipy4HbQDLZLsIVhFogu7J
G7lStbLsuq82eL1pAMgsEpySV1s3mYwojsOmWYwSGlUarb3ottOE3WKLdfmd47YyB7Oig/UwDoI3
hmu7ku8xTwiMX6v07zZbcPqs5GxSHxE9Ch16i6yhWDpPze3DR0VelqrJhSO3CfsFpaf64a6K4hIx
hnq3pjsGiwtFUfswQBnxyWa0d7gKs7GMb4b4JJH+TIK8uaJmC+fSL5qJfc9eHzGntxXYstfrtOX3
XZrQjbCD3eK62CCFD8AR+eBAQ3ff/bhTcRfuoKH7yrcmaqYLC1wVhj/7Rk5dEX7nweh8Tdh/dLCV
inQ/xs6vdxAwQaGH7noTwk0xp4rR1oO5IZx+D2FC1hJlnb0RW1ZjhIOTe2moU0Qpu+8g3jRg7Aqx
hH9M4Iph/fMwgoag9WeF0K2zFiA7CJKiCFC1K+D6iYM/mrZEDcqCqKLp50Qti9IobOKjzqykJ38k
+H+AA+3HKq1d16bLWwzis1NpKNL3I5IYDxOwu9i4stlgaxkLMi2zC7o8gVy+oOaiAIicnmHDugWI
ZYC2RMA6dBoqSdx2MU5u3LsGeAUytMsp4i5h/rCOzXkuyk6yPAkpJ/qHvqE51d/aCLT6iFZQ8zat
5PRHlk9hiPsWqCt+pM67JGYka/u6JEQEpDzq29Td5RFpAd4yL3mSm/cLIuA/QsP3SLstNnPLpY9K
GC9joFI2DS0gmrMf2vXid6Z7cPd9pRn+JYFWfwnV4LMfLmcIV++CgECZ0ltUFF0i7qEuFwsS5LbY
hFwcbugh1FK4mlqbO2KroDt1cZOOFnJZ559kIPPfp/Jttr1uBZ7ej9WeLTarI40zYIbMmkIOcaVu
5ZIrXzswJGIdGetHyzvXhM8umuHojy4yQ8kDskWasWLtmq0LUQAKiFLG1n5vwF5aAjPuDNWVzZEK
PPFwb65Su8zZj00DeoTERQX+/Asw0gtKWfUzU0B2JO8NX7et44B89v5Lu1/ArAaKh1qaMxSUJjRo
vcM4jIoZLuenmHEQeo11Hpe99T123WjrI44MZDJNlgdkJ5JxDTADb5Ez7deH+1tMSTxZcd275QtC
QUv1V9pKM2lz5RB61a+JYwZyw4vsHtLPidf73F6AENSK2o24Wj9nXPWF/pwHEKDf45ZSGmzClIYe
NG/YfywIQDG30G0m+YtH4QBAzkoHVQqz5UgAxVPpgDP+KcJD83fhdn2gOLvkcqYRvSfCfFSz4gdZ
Sbx3eWw+wKRAbe9n3gyOBnZt3U25hvv0US5DWEBgNSQbFsMFzjNVVuzHUpm4lUhv5bwLhWaUEo+k
iNtGg9PJhjAcG4s6oT1mDuvVKIUhgUyMe1s56xm2/WdK0RtOBibx/akTshrNE/Zd0e5ab7ubbY+/
c/Z8HruHerlvKF6fglGlXxkbqyT0kF4HTs/jF0V9YE7Vh0T19fcnoQhCVbkZPxPhOmJy4/OOreNu
jyphUleWJaA3bdtDB7alHJSjRfvvt5YWAWztqvdxEEdunc9KLJ5FhSMpGhBYrWm75VcS1V0b0SMB
PFf3dpxafClbs3zbnw0uSewyy5KJtR/LQiUf8SQ/BL58XNGxjn2yLNwBqXnNI2XRf6jtHSPwTXqU
7rodF/SOig+51zbSwX6TKoRXnugqHIoGDYkbeDH7NNsfuHoao400xgIVPcWHIKj5T2w2nOjN2yAI
9lPXgMz3pwYczMReYwBtuUwusAnrQ9HLmtzbB0CT41DlaYvm3Wi2Xgn5DdGLhSxLWd0LLF4d72fL
a3bSwhdbn83Go9SIAjvjAxYKndObHAZNS7enbF5Ow8pHk2lhwM2rmQAy89SevCOqnNf3Cj0EalNH
Xl7BVKDpcS8FkzpwvKJmKYBhk3+0ab7BNily0880f++WH5cfLHDwg0A5Mawd/CFpPoKn1Lw2ENuM
eLTJ79nU0o3QZ9L4HTiXVgtq18stC11HIELJPzRbYbJVgVat1VBSGOxUb2/MRBufOB1mLPXGkedt
//u5EQDtZ7Bo4FLOazg47ucgXSNDNS2R+MQ8avjCocd2OCLF2cZhpEVh7MjUk2xuD098XwIsv4ub
OmNTp83kzgSxPhk3QEhrIml1yos2YUPhOUDDHAVzBGwng1EdTYCNPIwGmH1cc+8vgNnMsbGNCMdX
ETOsNJ+3bqHEvh2QBTH//BHq10KC8JYBAkefXfe+jKSDBsIPJicHWYBztEP9AjZIS+MIgsUCGJmG
VagRjvZdG/o2C4+TX5wCvV1j620L1ci6S7vJxmiB94w8/mJswNkhRbkZgCXQMLD8fjA/asZrwpvA
RvlNvs+TOe9RbfRXDFNez+DWmDugDDOI2+702Jx9AamSSFBeyeq0UcYDpUBKhCERbLmS9t1Bar/4
valL6LkDrqHPfdEyeBJEsjr/B4ENXDDkbq9YK0U7cAerxhbWyCTfLycNXfKqgplHRvQrA7q2KCkC
tpKe8OGsHJCgw86JQNyFIsOf7iZVs9YpRygZ49+e2ZwqCVUdUSD22YbfKxG1fpkn++NZ4MPOELNM
NTkbF2xBIOYjF4PhqNWDFuZLKonUnM0ZA7BLefrofpwU14k0ADJ3xdtQVbGQ/Wh/u6Q0OPjxRfnL
EFuaoJnbm418J5yXRrkK1G5DV+orUEi/4oz35tx5o18DGkuaohDs/5CTwdVnYiMUH/BKGgji5jdF
sRQhuwMbmlQFktNtBzYga5h5qCiCbPFeWXLuhoZc/LqnDO8X1EallTOStaMsjoyXPSZRpT3iomO4
Xu1ie4f2wxR7AucarbsGc2lsLFm0Wk83XMgGxLWv3DDhywW2fgn4caQlwURBn2oX0Tg3O0yrWL0g
INEI4qtkqRZh2mJMZt4rxdttqaBJwYLNbcFX+DREivy5vUkAO17QAXZWkQD9wW1+rOKY4lPtACoi
QYSzvFQRrI0H4UT1rEGZFGj7SjqjcP1LIu9dXn8wMW80P1rn9YIGivGwzm+mGNIRpGzr/bQGtzq7
IKOzMPc3dspLcqwoWXuuYffvEWi0b8okE5WWzM9T9h4CFiL3HCO4ErUcH3DbJuNgavHfTiXxZBSj
efSZGXhFcZL7Gx99JSFvFor1wO0OohJkh445UKrA2wDFrlG6Eadk80mIZRJth4kQLHhMVp/wcuSn
yPD9Xl554907aoqEdwQCQXt39NaxecW0qFOMYMyYJR2nZ99/cNKBnxJlywZPcWXezdAItfA7rhjD
ZM/3omZDffQKHIG0ggbmPRmXG9OY9+7vBSbtZbpOhqXO/y0svvF1+hjqe+wXUEbToYTRH4SemzBv
Z8035OLT3e5Gm+b93jkCXe9MmD7HBJsv4/XpXv4em3KMbRA14rqFAXsXVnQAOfLgwmlQmHjfE236
LMMV+cHqE/Xv/rJr1mb8WN9FuZF//AKvvhKuils454PZoqh/68dsiswToT+XyezSfF7/g8Pj5W/g
ebGNyL6f9eHhXhOlZM7OVQE8Rk6PR7DL5YTTXjPQcUO2H9WP8d319JVPIUODTWatmjQX/qjZJJPH
mD4yuAvzOiJqKr9r5iYURWHmhWbtmU4mqNFBBFYI4iJoE5j3S/uFJmYRKDNEd8jI/Z4M9or34KRn
5/WMyL8tRFQlmsV6Mw3FQkfQS4nP5qZiKsk3ScW9POIHx16fnb7xZFfypavNOw1Np7jdXpC5lGh9
yCXO9m+yYvLmEdHqORD04/o7mrpPS5R/6CWROkDFZja7jlytOhfZ78pBzq2czMlFwXviAReB3l+j
5hiDlP3nCiOygni2YukTD7GON6EQKqNSEvCQH1SeK3UQZX/MjXPZ7JzW/BrxxdHqLmJr+roc5NjZ
0dZfmpWQC4mXBHbsybe1mVzWIyY0wHfi2SAAchFCZj3PkH5xLzQiE98Py4IgPa3Y0Z32R7bxV/ke
3R5I5/K67BMCPhiFkYEYouXyxHdthv02b+JK0AUqPdtBvP3a8N+OHWdBcHX1oYV3GbmITrVZmMqo
z/g1hxoa+Gytp+735tnXjQUzIthhnkQcgCWQnwwRn+uvyIoj8c/HLALWrABlhvgbW6LqCI2iNx8R
oSWzLOc1S/vLCVFh/gg47qBz9vtVhgfYDtd8e4F2dcuZkd+l6fY5wLi1uLckHEdP2PVP4+Jveaj2
IIDFsnrx5uB2rBvsLdpMNOk0aQy6YMVk16cHuQC4ROW3BfNCzDfu9BxxRfZz7BREAXa/8o5vwDxu
F5TzSRqgwqRn3jSMukLKbjm8wk4UsYy4wXzmsl3qLY9Z+Gl8uHOH+HHb/4bouGgpQxIe9O2DM9Ht
8+0HXOkPuxpk8EpWoni4RpcgxKKem64N4j54J1lmu29IXaLQFSvxHkMG8kn1NaE4xi80/2zZWToA
TCI393Pk3a9Ks+mKb8D58VPfOgpi2HN7y/7eyxj4ATdMALqWoBhfTciU5xWApz9zIGUq61en8jeW
angF7HHpvAGLIBbgNjq7VGuvOQHKGym7Ufl0vero3hCPUwbwztFUlYe4P8Fm07p4+07dzo0XJzYr
+HCsiyzsyzRNtFQsy8nUJHFK0PLSqacamAl9Xm1TubGiH0PgiHy1r1dHoAPeEXo5Na3leYzFaoac
94UF6QLtIXPWzuRwE2C5+ClsZ7SssKjvPH5KUD4gGTYmxuuBcYQiqL+m7RW3YYSOfluButCNHdvM
ST+tq50lh741uCOMoe7GqSsyoTz6TLwmfa2pBzLi17donXfaYsLRct5VvUFBVrLcYThAjje20KII
D8ivOeH/Lb8hALjJ1miAu9F7/kcTnOpGXKdOQCa1XZcJjWbhU558zyXf5W5hbJ8SYxsLmHqDMijk
/MPUj/XuQUYr9M/CHXTanUoeJhDLzsIWez45DZgau39AXVDy4I7ryv6BldsubT4bmbdaZu4UtEKE
KKGNwxx4vfWeNlOjvI1jKVSfBOJujdD4xeS8p1UFV3tzkNZG6JxvgPPQR/7QgNy6/eYhLjMX4NNr
5h8OeHcUtcuzoIVdg1Dj+aMYYXTRt4qL0eGJknZT9VHHQslUX1055Oja5HYr6Dx5vcWPuDlnCA7e
4/OZOwjh7dQQioG3lVwWCWjf0Jmow1nUzz/Y9jdY8Gt+nUl8dqDdU6RfllmK4FX6pv/KAI207EVT
dxnqNQOy4/qZr7/OEJVQNVJkbRH58q1IBF02GFrvK2U2/lLlgC8z1+HlcGyzfFQHpgcSqkhANXv5
YlOmbTwqxinDZQ/ZQguzzkZ7OyjRjhrP89VcE8ryWBiQ60bLyKKeA1x5GOHdvsMo4tIJMPBESnsr
9n3JW4Vpw91BtvqCm4HVjyF8cXufAEUaxSZbTaNL1KUd4wUedm/GsF/TY29Nw84lB65dyhqzbITa
s5c5IrOz26yyPYidCwkVa60MaEiL4v1R0z8b/7kDiOohUGtYLHsHm1T7PrYMP4vWE1DNtXlbhB3h
q9GYz6dtquqhv/S/csyAqHOm9wshvRK9YF+wPeBUW9ubv/HeNcyZ7FqgDU455UNN61J+qIN01hHt
HbOfTJufW3Q+XQDeSjOjK7fcApoAhbcP9xEdhHZ4zGu/7A3TdmCjE4HG5frJ7KrFtLAfiyBSDDzS
L73Jm1htzQhDuuotUQGog3BXWqiONCuEEcxOXsi0T222MDk4U4LGBdDOpRjzyHa5/PGcnU5iD3MQ
ZkgiDrBqCLVn0J0hNUwc0nIiPPIXdT3jDcJ+yv2vGIVhd9N2XiGLqYlcOCLUsMC/PDs0h134Xw5/
vhinkO1JM7fMwZ6VvadQKaGCkIDSC3qC6rK8+32E3l4dfMzAKYSRqyxW1+vbM0ldq4oDMbNFunRa
sm0d4VFpVyhS2pa9foTMR2FtdsH5J73Okknx6dpzn+e8hMVsbbsL1LKZcUooVKFL1HqKuTUqd6wm
KHdPLNJ7Wl8z1JwQS+IJVYjfAXYfE5/vlsR4yHVGIqctm3AxSzLtw0+QNuSnrXE4nCSIKTViFjzv
H1PEdr3vrlFLitpFOfQ1reN2ciC66SwbIPplhE78MutodTE5W7SDCV78WY+BqGRSrcIEN4nGEwnC
3lqu9M83RTvYNc5o8NvkxebXCcYRrV6zoEIgFvH+eF8LTELVZyWMYpM5N1oDDMmS4pBiT0Sy16KR
ZxRzlRK3DeMyTh0tS9ORNNIcjgQoTKq3CCe6jfTow2ilc0OYpMBmRL1YkrEk/7W9tPj5XNjaKY7G
Z5ZZOf6BMvcGoFapirM8ZPbm37OhLQXsLSQrOwBWQTEW4jm30Xzte19ms3BGekrYEywqZjJWrfpc
iP8P8aAMc7uEtNz76xs8APbEJVj9ZbkdSegmkA4uHTIExtg2mQT45lNp+IoaomG9xCzgfu314tNx
cMaPTD8GxyhCdtm7cpMCTOhsMbncLgnf9n8BIeI9w8RKYarYYQUQdbajk4HFtL1OeW8goNONPktz
HSP6Kc84zwleIpikfT15D1HyTfTe2IElyQNevB7qFoD9UCK2CQSlaEGVgTNjt89ssnjjPmZB3uPH
diqhnJOfS5VU8ntt61e8ufNCyyha+U9BPF6OKAd69QnBb3OxBil20NSM3eKsNMhrO6q09L185nTq
g/XujrOWOCmEoJrqpub+v6N6DnbA1SUr8vbaFSkwk2c/C183z2qaK3/FwmZpeggAEMaq6Y743NFM
UYrT7X8Y2ljWVw5OqOPWObSuQzRfFKg3qLh1MDPkp0RIx3EO7JJwwGqBRBB0kr7yXp4Z2BjxTpNa
Df8ViSlLJWaGfn+M/mFt5McVG3tCy8RCW8eMpJa0e8T/yOfX5ZEPx1XdJfuYpNL4mnaw60cT87T/
UmG/cnUemwaQe9OhpKC79AyAhEz+CsjPHzXAANyFwoUSr8u0GdvNlzM6QNtbFrSrUw1DBJzhBahS
6yqlzfxOzgemHFvGkOqnfSDxHiI+Sc9t86ePu4s7LDcYhy9fNmpk/RfAcLo/aNTIl3nG63cL+ZrR
XdTGS/nZes5UYqDOOVmVVdQ7veSlfLZ7GccO02/3PUUEQtLLrY0YuXUUtzqQbgZ17tFyim0QNYnS
Gf5whLhced8Y32uRUjCwcAv5qS1329DVZj8+JgSjZUb7TcICsSEFgYycXcfS0NdWdQJnakHJxKF1
NpJtw5Q6VWSjJ7/ZsROEFXFEw1VN+tDjrcFH8bcCPcsic/rjYn2BuyydEnrj+DP9w0fQ4Zs0IihJ
eq3EadRSeLSTkZ4whisZYS8HiKCQCIo0f745517uChwg+hf8ksS0bH/a3FxRjLxMEcXkBPTrEVMM
Y2iKepz4SbuaBoXN0iAaqRaisxZWofmaNkQRbEyvJG6DQgZ+9xod5B+G9fwlvYjzTWtnGKff3q2t
xpEMzRRDw+u/ThEbimiGQzgPsRKJyMaweOLPhXW6NSXYd2Ptd3im2CQ0WjDAZGoYh/i89rEkW+JM
sMx6nOHx/ybuvMf9dnAPn7k8HmNhnpRTGd5rOhseNg5z6Y8DCJiNCMJl4B4jrep+9ms9Jk+BI3Su
aU+ZBShg1qhd9FdeRIP7fzv5IPFxN6aoeccq+HSX2B6xFGcy29qPl8wF3BEYbcCmQTNg1OEtzhFo
2nuou2if3jlZNTxdoCYBlZ2UD8NMObzsgMCX+shcedWOTgdFsdR0nPiy4RAVA1iPyDnQh9E+aYk6
kSVf2crLHVKuwBw+IGlOJ5fr7tM1Bw5TOYbhXVlr5aSwUTw861VxhgIkY4YGpPvSj/KG1H3zS4R8
Dl6TA3mWA8NYjJKQ7dreCkf/1ZmoIFNK2+td0ETA1RXyw+tCPkDB+0RRgphTP7hs2T/ljTH/6vU2
yREtPGgr87Ysaj9OZqObxSqZ6rrtsGwXSRXW+f/nhYjC//g8qhLqS7UgpUwmk+GjLxayDMrQ6rd+
hVivmun2+CSHYfLvXfMZZfSbicH/vWf8KPQADSP4L4YtdABIV6Pcdaj6ySNFFhz+fOfs52/DJeiH
NmCgH/SsHfkQxzs1elCMq0UCtyR2YPqygkdLGe3dq7JT1WgtPU51CPFihkJtwa5nL1sehlSTBkXT
KWfU95He3JmvYTuDZR2mAKKkAHWP2R++L8D/5i7s6PZecQ/2qYKCY4Bg0y6bFquERNfN63jv5DAx
gX5SaG8x86RM4MwFgpxEIilSu7FfU+E8ntcJJFZnb5oz4MobPCXaC5PhYLJigeVQCxnRQkPR8rym
87S4bpOkfdPzobGW7fHfXl9624qgWBGyuDKEvkBzn+kjk6XuldBex0DaXkyaMasDX+RsY6FgdSGN
rQDbHrQFJ6I1eoFpH0C73k/yPL6AmgGdfmh7S9GBhesLHcapNBNzw7u4UhotUILQmmmP4uJGGxz2
tgJUnYOb0Gma6mqncMi4w8oL4+qK9DDouEIYo0Pjs46ca+MeduW/fp2iEW8KL8SzndfvRumrO+Mn
i2o4EucGZNZ3mIc+3xtbxV8sK7JuNkW4sX4mOfMv/qEoMngX2yHFdF2f382/RPNzve6d5Vi9osQm
XgD1qfL6j4lBo/CZRSE3xTo0V3Nc107x6oD36+uNwIJr8tkWgyHMC5gbKrcCqBYUdqtUXtVrfLDU
HFeTrUylgqKZpKVbZ6ezFg/SU/owLpPYOa2QEiMdCy8KhndoUTOIcjUenh7+5JSVmx4MZQE3qdtx
hcjv6lEtYpnUCUB650ZRWFFoGu6HcrZp2O+eKT/7TQFtpM23Xm0d3nYdpdzyFQKew3M/Le8Nazuq
bo0vUOoP4P6h8RDK2vp38XzOS0YhxMNekEWd6XQ5uTSG79UQUjzDjoeen8RLX0/I2K1lz3+Tgstl
S4njoUHCXA+VUFa/B1aEyCHwr6d850sS+Jkk6pXEKbFpr7m8OgntwgCHkH/3ZXd92u6N/O6RVNfJ
bJR2CYpbyu8AFgeYZX52o4bA2I97hM39wFhXaL3aKKRmsx37mSjduNLauXC9lveesXQxhkRds8lC
Ece5js9obV4fjrkT2s/xJshqGEZTgOgsHUvbsG/Z40MgbD3xLMsJWY4LSPElGef1rXIYRwF2Fm0G
ZH+0NOaoayUfTPkRksRbHILc+FjQ6D/qyJQ2i7kSqdL/IenwR7RWLmonfihhhUCAzV8xWa1XxHkv
9t4wqk1IWg5CkUForv4FHiqtk/jFpg4GRROMf6+DCeeX5wPfuNjwe9Sd1ZmYaVHZDc2fNzNDVxXz
K5YnjUjMoGwx1XdVKTQmOoPRo9y+Q16miF1eUs0XGqeQTmwZJkJnT1ltdXVmrJqXlzU8v+vr6YaR
BfUkDaYIrvzrEVVBURcuIMswblqDjvu3Wuoh4tF4plFWsFbfuOOK+yDCdUjCm/IYodu8rjdK9Wy1
3Knl1WHCW9J8CN+UscInyEE/DL8YiLxFX5XiNWgB0rRy2hMzTVXON7oAtzFKwV7w4tOgYEus/lEE
IyG6FexrnPc96eLQ+c/vpbuFIO6PfmgSGNjH2xPHJxQ0ji1gyGbiqrETAINsewQDjcOKJfxH/UtP
yvgD5UQNcKI8jVhw9mUHGVTUuc5Ac1YcBKwGfIRtL/2M20Ix7fWEPu1Q2PO5Fa/nxfnjRfm8/tbf
C0AkLeLJzvreodvcHPBZmBiW9NAlx+CxxCduJLHUDckT+pzlM9kyoK5GZDcCsBNfUNoMQh0mLnzL
NASTrQagPxrL3dHXV42JoT18QQq5QHCLqqdF+MOnS4QpwmYak0OxMc/WBsLHNe/11W2jVAT4gJXB
s5/XvDaBmrzXpf5/+19pfBXvK70iT9JP4mh6qiEbhv7F6I0q3H0MIlZpz4HtQqwH5lWSle9WEyXV
nTxjEwuKWae5p7Q8nXpkaq1+7S0eiQui6VWRzPJjSSEfGEiEeMBaeudVJKtivIVBq7Aj6d3DwKnT
PDau2vzrFkUv8+xwIaHALI9oo/n1ph8qKi4jPdvYBrH2eC+Oy+mbZBjQ3R3s8URTRFncW6HH3IXT
M2YN8pAuY30GWazEVqACsXXU7rQNVIWVb8WV8VThlUbH63EY2HHDfkLzWmqIne9nym6teFW+89WK
yxQE8Ig+xNbeCU7HBJG/WdOaKwZK7So3hExcfawR0ZkhYFKGdmY+VDOI5q9kBpvpTHqlJeuKRova
BFu/mIkMdW2nNHJVOyMTjeiYkkNHLigYvzTa88uakdegrWKmh2eSxiE1/b/M/eWMatoWhJ8V8CTO
Ce523auQWeEOtFJ2sA1b/Ay1ANo3U/cnBBgj2gf2h4Syuxf4coxT2IODKqiRZYLk+iaQuyIYD/7m
NnKTq2MJw1o47UoMGerVriV5fLpOrX+I11EBeZHfuvFesy2P9j5iP6silTco7DpFiFNjfWpCjTgQ
BmcpabCuwvlZ6YYTgAGJsciKHMhBVMJNq1ct+EfF+vCU5wTcSWmHSkOzq0yBYFc4sjgplIGgwY5E
822q/R226bUnDiUNAiFLZH5ibNdJBufsD1lR6zuVjaNmjp8GQUjhmonaep0HX+lDtMSZZ6QIRHxc
m3tAjBwaJ1LYh/MrCaer53SrnVjwdEw+nFz2/W77OvcvxsSHLUCsfULOpb2GVjx0mKgG1gcvD2gw
Fdl4qv3PZsb7n8iSrHguVGrHCVNEUtExGjxd+9poduXppmjAjT+ehOjUNsiF8M/SbuLYrwJtRVuw
DdvBgcWaW8lnCEW3sQ3iqiTf/6MCB2W+TZqQve9q9vIFJpPS+5qZNSBYC80aKrw2aJqEx36VL/Hy
VTl0GfjegUoTydJLg/etZnW/1BQXUl+zBn8Dtj1DkO22U7a8QvtT6LHOdcitaad+dE0N8XWFK1YG
gYxreIYzKlHgAh7t/YdkdAvgv1eE2hVcklaZ/+Eo8qTHyzWw3pvV5/6uH4L2iwb9bHGp6CDpkoUE
5BZF5Z5y0MALt1QEEKI5MSQ0cO2PJ8GFYm7wBmKHnxGH4B6z7FMsnBJFupCaHRDMZDHi6kiqWUwr
irtza8N0UebvSyScEgqBFxFzIANq9kPS5oMaUYXavAU0FnjJTjoPApN28B1j5gAorzFXKdsBpMmU
zPf19i8rcRPg++plr9i+IpTfsQr1b4FF+2ug/3XZ6cEjKapYMMOkoSsfMnuixOV16A/wpUCMnM2d
tFoibdhoRL6p2HgwxI4nUUmlA1sL3ncehg0+50wKc+BOuDzaBJDhPze9hmNoV4uBdt/1nrkZ0RNH
EolEFQHUmgI5NKLJ/SVBEogIfwl3Dcg4MLE+24o/Nx/q8g4zZdvk8TbjB/dDtV/3yZV+NX/vikoM
d9lQZU9P0IUUO0Muv8k9klw+rsgSCSvBmdO+wbxBGZx3ca7vFHPFXohKmFe0swZhKGw8dFL3LCxa
vGT83L8wNgaysA81KH0/31R9NnuPnLo01nodTOofnr9yoBq9JI2rbFMo1JjQpyUS/jbB3385FOEe
efRxUT69p6Mb0a81s9kMW7Y7Q7oPiAuGrY4DD3gynKM/h3DdnUYJPp6CYOCbgcB4F+IZ27XU4B5I
q8bKXn+Ney6sdiZfCMA79SPZO5jUVlXSXjC+CMRpuCY65dK+TB74bdXXUK/CF32/Tx3jpHcnZL+A
lNQP6G+BU9gEVoGDhPmhyqUhxwflSTIWwmR/hDy/I9c6URrPoqsUlj/gyRTuK3IEUZkNNdn1x1fV
evQQX6EOLR0xNaSiMh9JwRpIMi45aTbAMnjvHzg3MysVKwAlbupLjzVm5IufHWoGvcwVAJpjD9zP
pIf8H9C4CSyeu8tslGY6mFQzvPN7/BSqKNSOFifykeh+BY0t4quRWa2sJW5Onrvd25aIrTXqjZ8S
UElmXIJo0gh0rUS80E3+6Znj5U2erAA/YLkmmqsJzjtak8w6j1EQahRHMhcBCV7hI1j79jWhRP90
CLAOmzDiBxK/C6m1oO6ko1tStpa7ma0yN8jr2rDuL5nDTlrbcWVxaZd59ZefwybmQfjFBI+g0oN5
Wt39auSgpPM7apOdyEogs/9XwPbuYdSIuo8qp6YwbxIDWXCxmxAntE72LKjqsmzYVWi6YPNH4rYb
c847XELDxWCz5A0oFycneFoZvj1o19KvRRE/lDphaHRG2xNDH4fYKsAWOyK26mKL3uUkayesbR8w
Gj8mCayg4VSHj2KKXnjhnIo4rEj4VX5VKZs3YwphEWpk2WxDgibstGe04EphkmuLfuNxswu9p4K1
d7mXfdlV03By9T7Clm8dy92lYTiJtkH18KHBU7oGx/G/34Fs7NjeHzMjBR3bl7gUjNKfzuHKTBYB
AR27FK6mCDFH74leiR77gnDQqwDLKVVsUp4zGtsRVCyPjfg3L7iwjhj8BLK3p5WZhgN4t/r8DRAS
uacMklNCmf34ynKYXFfKhsLAltDLGU789XNUSRI6ZI1uDi+X+zkIu2c5lvY2nKfUpHddTn2BCD5C
g8cPJvKnz/d9vtc6DzQVRvPYu9AUKzjp768szuF+ZAb3Tx2Vk4mL29etSWeH4nOAwnR2ma9jiGSY
LuNiiYVjHzTmzBQWQVVCZWeELkq3VJDDWhXU55YZTUrlEFLPm+iA5d1vcLF2CUeMS+cJ/Ri1CfSY
2mpFyaSjaDF31J1R0MNn8/7mEP2M7Dj9QNblpTMF8ONQFVw7mcXzdKIaajvgyyNJk0Fx6LMpN3I2
Ip1mUlxkaWisdu4YDFbk1dbquEyk28JqCNzFDckVKdV7+JeQD/6ofS3SNsiN8E8JpjsmrWKgQQ49
iF2qc8a3pAdNkOVGioBDeqmAj83ohBVca35zIfqwXntH2ReA6HVLS0ciPaWHtA+UpPn9soiclEfn
cd/1eiUmMyqhIWyCaCv3XemQTHMrood3Ni4HABZhqnmm017Rs8BeVl3kqfAF1e1U8HRMWAdxrui2
FujX0O8JlWJKIwtHd/lVMoH9drnhGJuKvjlUWCta9E+vKlvzG+TCckV4W1uobV1u8EP3yuOcJASN
PCt4Zx9x5dFoiZ3onTc9cyGwml8gbgb80qLZu3AWg2ZTPQWZyqOtSitvDN2LPYPeavrQlsgfSpkw
5CTK03twxo7nxJlyjiMXbmgX5F0w3yDXGh/YsQmwXYJa5yJxUFz6xe3PhinXmiUbyjms538Smd6e
ET+RoJk6m5ZwCjw8CHOkGC1msIdBulgngj+olWK6mMQnCHL2Oieu1OiWBxLqRYoQaBVp8+JJ5dEi
iIkXlKlV4JsCYi/sagUpEm4H/OEavaLNHsJT8UdXvSlXgaGy52r/ngMZhEVEKzfSzIICWz/E+hQd
q8WQAcrYlRGn3hMosvyJ79ghd7d+tVShmfWDS14C4uYil653W5DsgCsZ+klOkkEZ7U44BX1kDfYv
reulajJKZ6PSzFdFyQihC3by23NpVKWnKHtXUc4aJHiMQaGCAEmr38DTHrPWIyBOOaoa58HFnq8g
XxiToIVMzKVx3OiNCyFeH9zBhuBblP+JN/0TQUKPQI0rd/9GhJ3Hlf/5vwwFdAGJTtitGgW0TS38
kUJDjhu7UD4nC+ehto3pAUgr5cuRh7q1QfxPjOmT1/wh3U8zWBHrhPiX7jpLcWSC6iL5muL38FQI
KP16pB5GKxpKkhtloaSJ+3zI187yPE8rj+4Bomb3bx8LcO74RJbklmpfmWf5vyOrqlP+51oTDI1e
cwwiJtxnpnOUfTTv3RnLrA2Z+gny8txIRMnAz2rpPfY2Qx9t8WAx4w7qz0Dpg/itXEa3ZUOk8ED5
VEFAX+eRV16eQhUlzxIAaoS18HEYWNbslnz2MUlp78CQXKmY8bxDzo+yfDWkRCp52y9NRfbdf4Jz
yOw4bd3TMaFz6RwkRfyYw1VaTFhVDxLYP5OQ+8LbwDzt0p/pjT/QyoL9ys/EYDMYjZP8i7HJbFpI
L3IwNYSo8Vzzzq3uL1GuN6QVh+VduzE1a6mXXNMhObTkpsN9EfDb2ldsKAQqyt38DJ4hN+/JoPTk
B0D0BMtM+JvvBJslwMquExYxvtqTqBh0o0JBJI8ii1qAPcftx93hNS/0csT573UJywBAdSiAmszY
KBVSSHZng4vrsEqKV6O4edr1hQkPaVUPkeE4WIxWGMZBSKsiE9HaSl7HyTBmkwSeF4IbyM0vUoUO
OFv3wsf8JyZgjCgpO7A+FRoSyFh0qzj6PdVxdHMUAcjQKZdVCd59lXpD+wI/VANstSZxtllCKYGn
+HSxrGPB/nzpNNhFZYeQPEHONsRqGahyciNvBtXpJpdKtf7CZQxzvN0ICzH+sn0eRzTvIYYMAt0y
TeS5/b33Xqxx0k0BvfhEAHS9WF+XWpBxrTgmgFCIN6cLiUG/bU8W7hGlegTgxLQAwToVD4hCsaRs
jHNspmUPTucv4oHR6aGZI6saykVIfSfoca34ecN8OngARngTbDSutTaTEZhoNAHGh10X0tIp0pA+
KekyYsjF68qEd0ubn6e29KjbVoHdsdGL7XyIKqFEKyfuUjcTLzV93fmRg2JZDrM1eCKGbUMP4dFB
rIX5AQrjbrrm9L4m8eZvPjRS2vzvoB7t1kd0cld/PbjJxhsWdhbZMKlehvYk4DZAKuJO4CZs7Qkw
d6F0ixykeGJBeIZ0a+ZPrQoW9gL/k0+UJixo/usR/hpvpl5oiBE2SoYuOa5CaEyK+nRldB5io3Dt
rKTcdX10B4aEPvUVhuYPWLtEHFVestlYJSLA/mPl/aVa7vVO4VEpFDr83gAqmdfb0c99Qdt6Yggx
Z+xL9rcFqfZn5kly3aPm1U4dSs94PVRIE4D1ucY8zFM3yDANQj8SFruGV38+xzRYGBo9TKLXUw9u
CNPguZojSn14LnfCfxV5EYnrZoiQ+e1AxSxoIKQbpWWitJOL9R8kXTLwgTw3rulhsD99hFIH/SqF
qDwlQcviKJBI7zoVcRipURPsYJCr9pSQ4JYCTl/LJNh03jWCbaK6TDlphb0CfmjKWvnDKs39GrZL
DjAMLePMLdc43xzVqVz7gPAaU/5pJl0M1+24WZARoN2jDEFAqLjtZ3f6g6GafsQ1agrrErh2gG9i
FlaMNGKBSEA5XgyCGJpL6O//e+Fyf0md06ui7cUor2TMAQkLeocU+HLKpGy4ApQyEZiS4GaHhuCc
UKiXn9afUYJTQwQwA8bIix5u4kVq2tC8A5XRDO4maLgwRBzSrSXoUOp2K8BK9pgppsASaCjckwvv
V6AoqUEMZH/ghUC1Eh1j8nBKQa5pSVrEf3HjvbVqiYCj+3gUDemmhze+CmbuUGY84X+vwdYg33bW
sryThy37Z1zuuos1yGIp6WUWhSRx1qI8xOaZY+fT3UrwLOKzCDMJ5BPn6iwrKDz57iqSIfbwA/4B
/pcgqVJtV2QBYzqpAOaDXQV2mepQci7ELRL4rrSv/9V5AYDbZaWhOb1SIWkn9LqwXsdxWzAswJv8
172DEieRdTKV3z4yoYmkZ2ZYSzxaoIsLGONN8LjrL4uNXw5GD4kSr0jFS7KjxlH1HzPqE9gE+3fq
icur24xXyJuftwPBXSQwVddsHQ4n5Uy4iXXD7ov/eUgiAnDSK86IFdvrfJE/WCayeHt6cLVI1IaS
X8nrKEHEwYQWucFwjyAh+4/jAhfxhnsxcwq64awViqoUHDdqrzXs4U4x87hnDGoIQJVxvMhbdtqd
dyWRJkVvuXA+69uSGu3GT/VAtUs2O4GuIHub7BV4yvk7qOubWJHl6c8zJqOdTNe4R0ecIw0wJArv
PF0i2dsNDjcuouL340b+3f5URGAiUkvOhm8ZT4MvegrIj5Sx3mrkeQZ79MPbM6ojYi7n3WGH3EEg
AwlCUWppphJqsdBzcmREZNk0wCnHR9dkB1wnTV7PpJkrO2jNgISX/HpXqPQNatg+RLiDEODa8mcH
tmlEntAqm+M0kDFPzGYwuayW0dQ/DQJpmLrEcVmir10BuLgWWRh5PU9aVvGGXazQ6LE43azqc50o
iuk6f7XZozyvmqEGKvbDvwOznJmfucoE0/PY/NgwsvpZ6ajO3kRgC1eEA5J/z99tWg9q7pdaRxZn
okzBKD+OrKujyzpXwoeD3ubw+wJTT0P9vLqPakMqwEw9Ae1vNOCmmblKRrFW5jmzVA3z8CBYO7Vx
i0astF3Xf7PLhLTeoWTGPKtbfdUYtKrbSfZNYIAwyJqTj+lDlf5rwazx8XgEXPz0JD2XGRK3TGnn
8ralUUUWy/MywjQ06pWUwAFIGagBFXFzB4J7kwb1ilBRkZpjhlrbwLy6CJbELJ4GmdVDrDkT+Fjx
RnJDhGeb+/sauaRPgkYG2NKW/FYous1OjmyKr2K1Zw66JMmsS/woQ+ztZUzc/TZyQ5ph4Pf8DSx7
jBfsYw6KQDlI47hZNDKQ+7zF4EVnHnyIdZbz32wIEBzAm+0y41sFjKPuMw5Qn9GdIARdp3V4mrs8
n4aDmCeavFkBbW0tjI16bGvNNDeunGKFMx4tfsfjso1oDqWmVomi+M47VnEhw39kiuf0jrm3lrV8
+HOwdxtBttFbB/0nhyAb/k/1/SQRKXfnoM+QMO22fwuOai/ELKnad4TUP5RFNXgVgw18ilA9mPej
FUAn/syLz00oOKwF1UNqd0xSB5UnMJihHEcEzeJQfpb7rNplV76QdmiS48LIsHaHrVStRfQ0qNIW
cp2PGpogAnQ+GFQ6oLcEEGkGyGyiUG2JLgn4dUuxL04h1sHYEPDHbVNRK2qCH9bNyQz65955FxVB
MYRaIHa4AqWfHBnQdw96TPffRfAsCkNpEjadkH7FIJa6ybfM1zinLtdtA1Kuie3yJpJ7Dx/hkbeI
9iNX+u5ZeHR4e7tKlmqTr7MtHpVnDlQSYH3Da7j1FXfoG4w6DseRnE24BhzlMiHdZdUgtf9sjx9p
06kENgl+AkXiVk0Gv3mMfkvWpRthUOwCKImvDgDe1H1FYd0KmzoyZi4RUqkMBojLWqtuO/3pZzZt
dpZkINsoqZYVF+5UzE0Ip91H03BjiWIc2BWO96/3hR/yvZdvOqkaY4sJVuQme+Bz2MHJHYUgxm2i
3AqgYAww8I6J799drhFolnUPpsI/KYmAgSYIItm0lHljPtEsyndMEzM9NU50iuU63KGVIjIOTKqU
/zCzhvrh9WNl0qG8cKtWhgZwRieGUujLJ6/zx1lZ+/mJW2Zppli/pQN50GLoxdcY3gSCUqJAaw59
HfSbTUSeDJ58V3hG6RjmOcsdtXHHyHXSPOsCQCVMopXws9Y3gYrAS5J+qW5jW1gEsP+OEWfnb5gp
iGKCHTyRXnpbiQJ5SZIQNFcySALeDgnQsP9kfQVcbgZA1lr0eeLJh8nKlPZ2vltPciJOjCZrWOCZ
WxrW++jAoZr71YNKVOm8xJy7Ga+0Eru6zsJVONFLHVwgFJIrIo7Z93hA+w5aradLvio+CCqP6URy
qVYAfcUkgzgOwNtrPxMTHCDVakV6DAixXpQkI+32xlWAFzFiq/XcUXIRYtYB18yE9aLFAtqGC4w5
BeGLV40ljfzllayTLpXMKHRd4vIDzn8R1ydEVm4pEyO8e6MOgYiy9+SRxuIleOUezoJh34I4mvbi
uaq8sgPphyoZ3Y0gqnqxdUWw1b00Cta3pSntuzc/Gi+pDv7eaIQtpwWRBr34rTld3VAiPcivfb+O
SlS14t4+SFdrjLAxxJoVFIROpM0wH07KMDvlk308FGp6upA1AX5oyMImBcpLZaEhT+K+NQH4Y/Su
XNuAuwHYCplwJZuzkNGgIfvs/+0kcXiYHj7b/AQCU7Lc6/ZKT4nSORc5dG/BSIAELRDdLdHh5KU+
GPoJb8STlptTVJklBOI2KxSKYItaLNZO7+2PULq6OzcXUqh25XlLq5fiesgpJYNTfhmQWNlimaq8
JgQeXRK1ln7VVm10bQ6akfX05xCWD3RtyqyXDQWVLfCVHdxauYUVqPIXYY+QVfLhqsDoy3g9/qq4
VPXIL2drTkX4iw8tV8jMzPmRKYvC5ZOd95YR8BsIEYg5TKVxeTM6AJGRIILAJr6VabAPNgCW2zBi
ECJA8VqhuGS8S/EW7qnGkcrwfjQoag/xCLOKPrJWFDAZ2gy6sUrLuop+INWAKxyxuK4iTqLBPCSU
i7TdlW/rImzgw+EsJWdXIKyrlP04aiHTy83F8Zn47sTfxUGiqdUVkVbNqbi0u/qTgPOTqtXmvsUn
HmXBvSj36pUhJYcV9H/gvyfxOtlbtOrJamMnhObbVT8zzFudvpoRnOe6FTm1mgSZs3kJobixPxGl
h4xcO2VcT8T2TdM9MeR+bbLoNjMz8cFt9WKQQri9UclpkoxAsl+IebpAe43Yv+O2vKVviSSn5H+H
4J3aPsgWcsuGXaXdjsOdL5J5VIaDKR852Tf8pF+NaDDmquH01PP5wJxSoLIR+3Bx0Ky8yLSHpguD
/LuTGgLNdNDUmDc28a/YQsbw6wbi3Wy9m30n+luG1cC9bgX0ki3XH/mIOoeAa/mAhplsWs/TDSwJ
IdVMhrHm4NZJAhdjmHw2uCvo4+Z9O6vlA7dhF8eiZmyqTIiH/hh/Xb27puGJDTzFRrW5O5Yd91P1
YZsNMsVQL9C4WwSLPsm9J5Es8CByYfxAvyIwL6LzgPq/QOA2u4YXoc43wXMEHHIFq5/LQ+0LJvnO
V9gF+i8TDecatju3suR4I6KjaHoidn9EeSL9zlbJusGgFHTgKfxfYgMf3JP+H/1/oIWQNs/IB2MI
xDRZXSKNyGr1oLZ0V+K76WHXSzkXOsWjNHqUdUQavLouHpHQl8VU9nZ18ASQCkEq/D8XJwDe221J
6LGbEuQYkPYDx4OFZJdo0gd1J/jmyAabO8w97tyFlcKPOi0ld6Y1OvJdTQnLQUrbfjbWvdK0qk4M
7ybfoiub5GOHOPQJgv7h/Yzhw2zhivOarxY4+lPbuaXL2Bvt4w0J74fift7EEk/y4W1z7Y86BCeL
oqrmjMTbM4b9oiEWyBG7FcilRFTcWiPmaKaLCrCDVicm2FsYuo0kL8V/PHlfIRqTYocNQCFp2zND
1GwkKCDZvyJsY54fdIJ7zrzVToWpNkqwz6D+4grgI3VNXoChH4N/piKXZecaSqZ5ipjlrNf6pexW
SpqPHzlv+LNev526HU1ghCydNSJtwQtzxJdjoOE2xJyTpIcCDnch6cDCyHMafcOediJ3ozmLnWej
jBkoUFu3O0o9qPmS3Pnm4jvP00xuVmcJstWH+gGeKV/SQdpJVY8vYcMyn433gsuy0eR9YS+efcjn
FSK5r7U5bHeMUC5KFKQ5ZAFT29dyLWnn5ZhWau5cRD8m/cl3VMP1lHdaQId1oxIUXdTRmnz8tFZ1
oqqogaA+IPYjGQQHRW7FDA1Zn46k9hwLRZHB68du1Bep4PYvbKf+Z3M2FXCFaWgNvpCiTL3c3dkQ
LmpxtoYCdl1swEup1XmfEqGCd0AEo0WsnU4i7BiyyBK/uMRDAEzsO3tj1gLQWerJDuO6mA3tF283
AiPlR0dxPUfa9V0+U6LwOBmeLLg59qa5o/L3Hk7AVzVpD1C3gFEjgDoD3a28GeT14+xTPz2C2tyc
kbNS2eZ5Pcbh0Aab20YUQIuKPWFv7rLo88hPze5quZyUm07DqhPzm+nDDpHb/7TgK7kagqToFdWB
3QzX6UwrK68K817hbNOc5VRuRYEJUH73lxkHXqLcKgRtTKZcO3X72XCgl8gDRZYTZl8TpZ4cvpw0
cMCdJDw8joWyu1jAdzaXIQgZ1DpgPvaTqcyPAcuzN4Naa2jbXdMmGKxd0dlO9F/qWbChWPiLfwB6
RORPw/OXjQWLwzY/oXqaISqdPxgDj0uErfXNUwUxsnyNebYdHoCV7/QQUA3Vge94es+Xhgn1zfxr
vJKDSWfC5fIed2ZZqtJgFEl8zbHfEVPrq2GEQaIcd7Ewi+m7qWEfXAVeo30ayOeGd7LWTQxJvyt+
NnK1n3s1l3IvcDaYhjs2A5P0Na0IAMrqdIpIoGNRRTLAPstQExn0oOBNP8Nwq864Cx7/rA/ky1DW
/E5eVWVwooi03mqXQRbsPG9/nf95BbFJ4XMqFA+9k5+2uJKfySsGspzHuDG2Q0558EpzgVMuQ6po
BIneDOxbjfB7m9w58W3AW/gLB+THLTC9Dw0zaRoy9z1bZFL1KD5zDkDy8Q38Tm6lKzcH3h+k1mCQ
UkIGZ/A/dCQ0LrO39jxgQQbbgKl7qiUE+Lxr/FsI8fzddfCgUgpkq6yyGgLl+i3sbodzELjZ6yqs
kR3ajOqHmkpQMm5NpOm54wdf1etRWpQ0Ci3wR4A3bMa2hHQ6bMCGrMD4nVkQvpgosBRLHd6r5izV
m2V0iT8WgdW1nQMqZ2SR1FjNeCMQ/ee+ZEt+uw6WyJ1o9ZqzMZW4WyuPH/XCkAe/dJiQuJWgAytb
SUC/YWFJUX4JnFUSd1bBdtrvx3xmu/1bq/O1DS26Ao2wLAEdqGycSFORqvctHwqj64K3SIl/kl+l
U8hf1OmAFIB7ZFohH83jyr9zZAORyYEyZ1EFFeVXPUL5UYLiWMdjMlWVe/C9JhRSJtG8k5pWqWqs
jQAVtxAKfwpyxh8UmEguJglsva0VXo1DdQiT3sQva6T5MRHgPvdDqXi59RFC/iuuauBjR1mAQJq4
wxCf2bBdq9S1wa3Ff71pb5spUbJfvs+KbsYa6ex5L1xO6BIyUvLbuF3LlAC9NbLT0hJQR8lB0wKD
c9NrWNjf57uAEorxPC9ibzWjEehu67mEXN3OqxZkfOz2oas1Cv6Kx9h6tU2dltOiUGW+Ekp+HDlG
ArtWEkQ2D2q7h0VUyp3a7hALZP92sbyNwT80IjLfNhvNVWcxBENR1bwOKgmIzk8qm9rWSjon9OtE
VMTCYKHvMez26G+pqJGwKM6Ioib2y0qI8bquw/bBs5mGvpG2wdWYjNAw4q10VBVSPCHVnwzBACmS
a9eb+9K7sPIMJGxqLdSKovcjiNci/8WlN0t5THRO0eBznwAPpoeHSp5HIpqG66Jby0UziDyn5xOW
tEprkIx0u1A7kgnNX8M5EAKDH5zoyC28bi3IkUzwz644J5/J+B5OhH8X3AkKKDRTo9W4MxvxfHD/
OTM60FUguy8/rZkLULtf3gAl+myLLO9CZHh36FvhTADPZL95VWbZ1h6TNmScFW4yeF7p/ekVfPa0
fiYIOGppJlBNHLEpofAZH7FNVaE6VkHU/qW+NcoQk12i1XgbyXj7/5pRxiA15qg+InLPADvc3fe9
9n1Yq+5ck+TSDCoPlh4mnnhzBwOMEJuoHLc0WhI6MCWqIpIRImCw+6rxGguBShdG20GHYWgDd4oX
YP4KXag3GpQE6xRUIQNf0zVGj0sJZbTRXjSg7c/uDNFHNKYqqPryzijKRMXxMY7ip1X2Q6SM4pOe
pMqsUcvPB9qc8MMSDlFV95GrHvN1Fu/cMEwrg0+tVyTHJqkm2rXZpNLrRw14vs16uNLIAzbb6mxF
szCexdpKrsteUCEyyuzv7HwzBZXL7B4yNvfDMSY7fTovQvaHWJm2PDcFIdwSqnjOhddJ/JVTaprY
IleAyLrDMgoTjeWQaYhdpmJsVWcZAJI/9Ob0j1v2o0KVTNw2ekr+Qf/OcHA9CJvE/etcRTMvHzDb
No8fRA+De0sP8Q8rLgBKTE0xD1K+CSD1U9h1raHY3VnhFdBX7pW3OmqJrlgC9ZaC+K6651aK3s/+
y03doGiaqY0jW9lyyNdEyzK9DJ8wK5/gX3nNoNrXluzwtwjfcpzq2vTiV4u7Q4XtWqaDG75mG75g
2nz48wMcs9r8Jiyq+Pgjk4nbiNP8nCt/iiiImudIzekvSGA9FW0JKDrB4Trx5MwbZ+9xGjZtLJc9
muQ3l+N5ZJ0rksuvGCncYwbNjv7f3c7CCYTMJORbI8cYw5x/U7ubT03ba+fM0x4xOKpKweqBDgvn
+KaxZNxaxA8sMDyEW9PRns216Z9BylxBECyDqMp/ecVd1t/6ynATK5IyT9uCYJRA4xmmFr/YCHqi
o8S55RYCWeRnitE6S114kE2I1P+ffSDWW18C3A5Xfs2eepURO9/N3guiCmp7lLuBSK2iQQjSq5HJ
Zz13ZLCYYWxA2G4rBoxDYKi/vaLAsXZpsvFchdHGK7mWwjgRQeZBdRpkmKIJyJqcRel9tIggDdWq
nCO4juf2gyW8fFNChu8kJQqWeDWoW9YNnQrapuRF+1MXYmN1teWthnzQ1oQY9gjkz4SQ/enuAXeA
UX5JyVW7ei8y3hWllNtoQ0ZGCob6SDy5kKkKAPUbGy8L5QG7tzGZgrfllTV+mIlvs/EuQ/0jscwN
p6TYurXi8eA+CnfjiEYfbynFm2005TQfINkFN5GT7jQ+pGfXcA7amyoGKXHOs+IVeafA3ld6KlA+
WEMAaS0U31SwSlF2SFHzC739NP/A4iHrfotbnSBzBg5OmxqxKSqH+1gQ492M+Ay+AGjxzhAgRCHN
qvF4q+6egrQJCYNP1gNoV4VaBX+YexToZjSTv9OzVJ3QOtcAxMQKOKYrgQ18ZNxR0ZpSFAwxjfl5
Luyi5qkUmvDzjvLQnvHYWPKqliZksdGpHmNg3uDcbPT9BKaxIV67A9L0ka1DSP3EGUuRTRrLZJQo
ZKPOjiRnlYSf/0/YLJ0U4lP6wYenkPycPrBBSMsDf7zKE9tYrqRzfFPprA2n56TZ61CEZ6pzBeR5
IMqPA++4aIgIrDivE7vgslfAx3L+J9Cbjwrdh0+hdZIQ2PLSyKZATeta2yYPvEz+en9gVgaRoCxz
UEQif5dSvs7tEza+8SAFuYqxlskxRCDcnkew1CgMZOlcN6fdn1NkCE6pu+s2cftB019U+AX069gg
iAfr8f6Y34lRl9nVFmkX+EOPLlaDffytYb5Ey3pb2Zw2ApZeXSjTl7vVzxEU4ec7eeKjFPfWSqMb
/7Y1bCSUX0m37gSwMK+BntC/2NUnGL4CrCU2bnBq13E/JiCq/O2TPwl6CpH7Mf+e4i8VYwfaHu1s
dtk4snXCYLc4QAjkQGhpYLHWnz5F153E1iupNa7sEEpaAYbOa8WF5PqdAxqt4qLRjqcvC1sjgdIZ
rIfgmz2ml/sKq4ilY6Ztq+A6NLUN0+GwtD1JlG5v4V/xCK4Av26oxv2qqsqrjt3pOMbUvSGCOuEK
DSFPBx69nK0a9iaIzCT1fCia5Ti+clXuzjQHd+kLn1zCVU1jHtE+0Adm9V4QnIW6yGt8YRI8dOVd
WZiZrmNGVQBvHHl038LhPOwThS190btHBwzns2DEp95+J80Y0Lpi44z5EW7Qac+U/auwTgToezGb
El6AFFH3BWHE/BUdEEs4BPHPNPlyFyasISKUxQ3wNJ3PMR/+wdly5REYJaBF4QKVJBHVV4M+mISa
YZvrEc8Zq4WgbpeKd/4uCNV2sjIMEDPbYT8t9HQ40D0jeG2OFlbLdrTAn4fYKdkwh8BUmiANzSbS
v6+tFwqkCzTmu2usY+QkAgcT99P4NIMTpOOWr3n2wwF6cjdIqs+4vM/8ftKJYXjFdSI4IRZ4q79V
9YirqjqrLI2SssGibwXA97EaVrdNeGiGnKZMhPKh7ERqOm5ZGB1/dEM517JtAHSNrT+yebCeFtAE
VGGsXSZJRlR/4CYP9zGQbU21b4VoKrbVWZJ4RstMuzxc8HBdrrTAEYg+xg7ccLXD3uym6ywxhjlB
UugbA6TSkDEK0CJpmXPkEzt7/tcdMoni2ueb7tt1ATnQzvYWY7QUIDdFk5NuuTBr9OeVuQ3g6ImF
OSxGpP+9OUdBMChUPSDh++KWUvBxU+DNS9CNb/9yfOdv4pE6xcXq9ZUqOo3hoFEd4Z+PVJFLRT4B
i/Ft1hXlbatnbhKeOobvk/5FfsDc6Ml/IsCMftABFYogZghdMBoLtGwyEj4sb/sFSEwZ7ufNTwe4
6TS+3+TC/2eSJZ378KyGhxEK9D2gKWBOxhhxi0w/YxjrgR3QlhmipW1q7PC6+exS2PTVCdZ3T6b4
KgMj10eTrmlYFEA0hnF2VyfZWF+yh7LwqG5a2xcVn9uESLXnX9WKNk+BJxNtlhlZ4n7so0egLyqD
IR9FCSjY5MXmaAKTC8mv6JZrq5wGUcD0dflXYyydjMnzIJU93XOg9Pb7KfV7IBS8uYAEcjBqle/w
M2W31wGYFI+5pt8dEFL2sQIGYf1m5SMhQheJFingfZZ8Uk71Q2MlC8QfyW0EWdTnahqfPpNBtVI+
xWJ3E9RUM6XB5N18yzHvDtRh4W3NsGM1LWQa0HiIld4tk/TNuKJsdiVOCb6MyX3qRc5Og32L4Uki
O+YYz9kfShg1EfWp30CWRI2COeJjkMUEQr22aXBicvnRSpWZgXXOdcEWzsIWUzFEKqPykEcec5CC
XKzQ1UXSKAQmpD3kdEhNMU/E/hc9uxtYNPRnugLJ1Xkx/i2N6tESAztQdCfxPslG/5M5kIyARCFC
3aOSJTHklgHkLXmSIvYwQZg9zgDC8e+rN6Seym5jNVBXakWkkIGiXWFtLRVlLO5+OvJ+ITzMl5Bn
3JgP8ZIWl+MYcbzWDD2VJzpP3Brq0JcikNsJtVimIYm4zXjZElyOtGPgbgJC85CkZv8pTcxscEy/
LhV4w+Yxb67OhHgwlYY0gXDsdaQho5OFPQuCMY8HOjAs0oF2ls9XF9SdQ/+HvAjkTbqOV8VNW/HQ
HqPKvHzQTzrJYLyw5MdY+Zt+w5vcklO2Drxng7A2r3r2oJh2jR/6gcWBo+HZO/c/HHfAUt4RkR9P
FqXUii4+TSMKJ7dDNNHLCWGsYnV6ySVBwRm4mlK+p1tVhKJNc2o6URz6iZFQHo0yL1Cf0TbxoZN6
sMK0XXhWDZniH9tGGjS8kmykmdZPo96dJfpFZ+OgZjhlKdTmZu4tWH83aCazK0A8dic/dIWWMWQj
H+BwftPPgQOeGY4zw45vPWcW5R2iRwnn1mFZFj/6fyuMsEHWjsI9kbuIE/E5jkV39R9ze0U5itrX
KguXc2zuh2TWkRTNJQl+D5Nhw2nJmxE7u9hoj1ILNJZxfBo76cDQukb19a8GTmHqn9kCNDhtwitx
rjr/f/h/qftvyLGloGHyerWfghii4BeHt/YRKICL4DSt/5a02UGa/07jMPeDJN0O41O1SDzCttlS
j66J/hGU+I6/kzMP4nRhVbMz5K+Zng/sxFTxZ7eXTxNfkAWh5rxtpszJqF0x/cUoLuJGT8TaUZP0
wpQ1HusIirJTgfnMH53TiRmx2N1VzaJfFj7zwPu0sYhps9mRP3vIChPEIcaxmtBA4KdtkZ6kZj6c
aRcXG53zNyWoJEu5KEI9d8fUCGdGDax4SoTyfoe5iTut+D6kDYvN+Qz8MlqXcjRh8DTgaB6g+hEv
5cLycUfQB7dYMk5b9D56xiMG0vFdqZkQIKwmoYaFP5Ags6IIiP9gV9VhJMTNKTvvU2RUc+H7oyT+
CRJeURWLvE9rCMjKYlUOiBC5OIUdiSaK4CZaJlbp3Mhb9OaJf0E2BxZotZClUhYe8odLY+jY+DCO
hqdVsj7QoJtw1AVD2l0eYWGWRghf1TV2Tu6USDDO5Jo7vwgbhZBHY+A75YiNf4HxsxxrJbn/KgYv
2ndWogPaRj/zapTIyfJZV/29t648EPxC3XPylsa4ZMtpVr+9Lo9tv35mIoSMIafFh2Tg9A+URMS8
fbHRrxOflW44R5tnScroyDampCZptUQE54YlHcZS2U6PRDnnryqvXp+GSUKQRJbs6+WHJjKs89n5
y+fy18S24dOhBgVqCcnOKe6VNKHAcsL4T49xXI2sA9nNrdHAVhw+xzEorAd4xk5uGwjeBGwBEMQG
F6kWqZOV1asI2zEGYcHMleqFKJe8CQPw/MVOJypL3306tochqKDSvrBFjsqv4MQ4IkiD+JojodQA
IFnFpagWj9nyWSlrTnKvzaYurcOiuXNeAXxuvBHoinJ2O22gdALTJXIh/ZqzecSpImAqDsPYE75y
tadpRLd1s5m2qh09zgGsiydppKlbjqSaKG/UFNzcv6utk4XnfbXhKxnmZLCwMR3OXqljns0GQFM+
lTJXveCmx0MPGlqzu8kVHcV6woDudIUwnkQWiJL5SQMONX8zczQKWbCShswn9xKIiPB7J5CMnHwK
wf6Aso4U8lv2yq+O1aPbVE2aSHXyR725agcnu/JiBAoxvdwx/YycbYipHpX0WFb6dgeYgz4JZZfI
y6ZSTdZ2nZgY/qTaagO+JcfJZJl0H2W5Dq5eYrn524tgBCJkqsXL61OOhKiwulSyFFcKEx5/BAMs
V9A9jK8m5hEQlcI7l2c6ani8/Yyxk1bBkvtwdMzCK1jsokugjvKzvX2KaTUwacr3t7jSKpuBgfZU
aPvEGcXs2X5/RlhIMNLd5tZSVeBSlW7KJX8pNiMr0cOlLuglNkFBgJTdoQiegjanb4cJ93K+GMi0
4bAjMUDM18grP/Ke8pxQ5KxcLxV1gZUctK0+nh6I0YfxDqxIuQPa3yyWUz2sPaG2NgyiWf1uQtBs
hswJeA1e/gOHEete+SkrTy27y4MAThLgUNZFgmSdGASXyXjpua8r1YLoOGSXl4XuxRAIwKb+lyFI
VyX4ejyrME75Lp781f3fh4nw+E2QddVWJP/X5hFnfUjKeJc7nWzr+Wscxqyg/UPW71SX7STgv6v+
38nQgvMtC2m6PlipO1TB9KBACECu5fMLJkVhMTQUIVbLPl/ryDEkhtSmOrsS+msTOJ+Zp9HgrSn0
QoXbv0XV+9vtVnSrNR0UIPUoJDZLZTOvjmMeY3VZrtkk+YtmMJawvSeC2qzfP4S9F3v3NviJMkbK
qLcPgItqBdYrFH/3Hh+pVIi2gRL0Cj5ElQRRqRgLYRcxw3fAKV4sYE7PCwiZjE6XtSs3bS/TEW2R
ijq8pra9YjL438SCNe7qZ3nWp52SIFKi/TjyVm1MhjtLaEbQBK/lokv812h7FSGQyIHgrHCxASzQ
gaf3eOCiRWi0YsehGNhJu4nRtbpALtQBqcjmp1SQNfb3YUkF/HqmAHpV9u4W43hndIAljRTsn/lc
w8FurlnOW5hUDkFDG9brnHCLZH2i4us7gZnV4d8alP9Wvt+NVAR5goTaqe9hL5RLt3ZzAKlK5MN6
c8liQAvv1UAASsmyVKQfP3/CuseiV+wWYAh0noCO07eOe7Qc+2n5srI3w+2u8jOxHc9YDIJSNAyr
E7bLa5kYYJQA56eEXaTPhuDT55U8267F3zDRbUGnVSP6wa+gTsV0lAZ3b2DFtrxrytcLT59YmYeV
P6Ozj41ppBe2ojWrROJHgYqNMOWY85YA8dZoe3vB8yszYfsX7zZIwn2SV/CQgQpAvVc7pLahSzkF
CT84XRQjpAWEiWFUOxCxerrdYNNlNjCSkIAHqi1WgFJUc7mXqk3yhOZATxheSz35BKnW0vUQNeWI
M/lhdhiVb1sWQ8aL7JkpeWsXaY5U4HZCsGkBQYvd5JHb8KGEJ3PoxiF+UUd+OrrWI58guDq+S5/g
MfdvEglsGcknJVmbbUBnWwll1GHBrpEaxm8s9++L+6nWbPhrbjYiM2nTx48Fx2ruOeRPTxoCVlYB
9FwOH6q3QklIBNZJzay0Z6usv1NNiLnEkwL6ic6pi8+kq/CfYMZ2i0eA38bEEWd1q6Kwbxa3L/Eq
evOy9YRebD5eBoRM7Z28/HXrtNFRHjYX6sx24nrnwxbMH9PN404FpU6rLOcsjIC7DWYtP4UDMus4
ID3RW+nyPqm2MrPpuuOwjeu1dipgL0o6AOB6u0kyff0FwhhwgKjBaTsV1XIT9FW8jKGPYK1j6Pjt
6tdLdbBKRjPho1++VTBJaFAW1OCuimRx0RKbgg+jfLBeTTQOoe+1tF9Q7K9qEBe8Xz0JwJTkGF0K
prop3g58RKMxcPi6l8hLCYv08jXmBLb7gFjxMHqN2KuF5fQ35WLWkod6CUcKkBEQntSNHwZhNNzq
f3jGsOPIYJlETBZwfO5V1g5wrHCF4kY5h5Dx5FnUgikVqhCbD5Ce9JF8Y1sWRYqSJG+t1VkturL0
aK1f49/fFgvAc4xXXptzgMh0JSlwua5fIXgRT1DzKfp7fNlA4GMNtAK5jNVnKoqN+WZErOXamXMz
smv9EUIPo697WCWjUyW7nvQmRf6+gIqg/rQsZFYACVq9Om+K04TKie+dZiIFZPavLoxgBPvQl5oC
cLpdneLrnpkniT10SkwtxXQ/H/R3iSypzkaCmjlny2po5VdU46ug4aikjJY8IGtgASFOqOKsRQVt
NydsV0do+KAANjOFLgeeGJouA34w4UevucMKaPZPX50UUtOq5Jq+J1ytn7gLaeSeEm/sUX/4V/Ov
Pb6nXKeumxJX07O3SgslX5O6ylQQX+05AONLfhOQXCR2Gj+c3SNJuOT+M+ujnJP1jX1J0yDJXV/C
1x8Min5OyR7uAefVYitXYoVIoZdF9B4RyMMPB7/DT+RHYogMcqHhyZZqF5eZEwtKvSxiJHkygzpj
cMJxBJuMkxrXWSyb7wR6FfPwU2gJ+ytLQnnw90RxlGJ7D6I+azXSezgM11DPZJ7TeRNkqIGUKD+I
yI7DzJY0XiuvKfN3uqceN4I9zPwZpnKPvIFlZ/PGKsa7RLqOe2+VMgoBr9WihS3noPBGUOpLkm7I
7IqiYqID8H7t+Q+4qessizrknhGIK8dK6m2kAGhXm85K37oRul0ZaHfbSTVw/znVoWeGzSpJ5W25
fv+F1VqxfLCTB4GLXiBxXUiLbQwlWgoblkNYa6PI7B6sl9+nySJJSvU6+ZnKiFV1vG/0Dj0z++Mt
1hO3W8AVm/bXk/+VeF4DL3D/eyRr/adEQpj34qLfze4PGIiELMooovOHl1/7YeyHlf6EfNtWtebC
7wytgugDz60b7q6Z5+OVfFyUYn5nvd7f9ZABEfJRE93PkCOSXgzf37DKL+2c2Qx7m18jELqq+sp+
WkVnNidFpS9KPjS6Sz3P5RQeEOuIczfHZgSWOgKBEuCTgCg8xD0Fu95G5LDJ2uS95sKD9EP5tNHp
52bi7MUpO/2WYHxacPcunDxhwIvhtQoTlMAoBj2L4j+MZrbgCDLFRT3dMuVwVaDSRQAtYvKZG3lO
EjP1hvcqdiXmpyU/st8yTGuG7xMhihURkwoVadtTOMrH8IB2NdF32/mps42C8ereYwtxF8SW+75P
S4s1WQfzmFOdubdb2kxYDukFDqVzCsebrRzfq9BTB4xEOVRV2RrLrBfd/QfWdBGnRCmFI4Mm0yIj
lrQOfy8i/L39AoLU9XZ3rsij5TKOYhkr+eX77JEG6cTDASbghs2W4lQTv0z1H5vHNDInz29Dg+OM
qNamiUeY54JmmDLYv9NPJEyOzcn70Itta9JlKo9CKVjeBzBmWk18epQ8HIdCL8VichMFzBASR5qL
HdbJ5qjDwYuTCHQzkO7fTwSChlZQa3A5ZdAEU5AIBObReQipHiklPQq/eB0ClXcAlweKkmmxgRA5
MHuv9EY1afQ5ApWT1vvp8j+L9hGrnx3wA3Rvb6C0fV73WXM1rzwHL5sV0qnaa6iiBnjwou50jLQk
XxJmmDLDpnEiBmJ5RUUH7UXMWuyeMDsSA6iTLrV52cQ2ADth7zla6gQaAkVsXMc0WpBxZTmgwC2W
E0dG3vv0UTPPY34e2qqVVNIHlfepbmyO5c/rCacj5QtnXzT0JgvT/aprjgMuRhz/KXWul9vAcxVN
xXQzKXUsbD828McioIMV5EvIx0MoD/EDydlB+uuhcW77hDB+J8VGHhBJze9+hGd4OI/fiG3RLEOu
b8uTuDlKy85tzlXN1LN6FYqKears5cxJ1bWh2NKezPPDjzcnY7VAcgMR9pSAITVWk6yuZn74yYCM
/qJ2G3m3yg1nsbW8HZ47Bh8599KFVgpifokQQHutp3iwv/cq4uw2rI/YQlWAC8WRQyQNH8/lDnrR
gQmJmZFLNhCvyH4Db67VuZBUy5igrGg+lXDRX38wzswCXSZ26GtzeuyR4H7gz23L4Ymisl7TmX1Q
DbOEedqx91gZGmYVCpcBLxT/hWjeWwIRgtBL7P+EfsJdyGhHeS2QF+JrFsEhTCJ1UZN4GycaUwFB
i/jtijoCPappUrHGegwM3AjuEMsUZA2veGQ+zeFD88aS1w0WW6Hdc5BYd8+TadB4EjJibLQfIlFB
Gw3Hf6+fafH5UEeQP34gN0wNP2ce/eCjf2SIDcQ1+HzHlhpAle4SD9lWEGpstw890isd5l0JCVEh
S5JvizQyUa9JPVgpWpqvNn/8vtxpHPzkQxASX9PvLU9MsppD/vUYkl9catzGXpfmIE3LndiFnSTT
bDrysm/5hZneWmbyc3RIawJH2c96KgVdMEqs627XzNkelTW0dg7SrU6MRTYfDZe+wU8CLRlmmTvc
PgROEJFJmhWS5k3yF9A9hPqFDuHuZ96jPStzvzfyXy5oJ5YZWuf02HO43mFUnpHl9It7RVS7cIFB
9Qmmw3sNAT1qpSwliEFQzD4XJYt+f5eHTGDpvgssODPvzyOCDqaUCs1APtMdvH5QwluklT29TMpW
HW71083uPJ40YmAetyBXqFW6v93UAjDN7r/avF46b+KhRI97+2pDbuKguMJFtH4PWsoS2lmQEDmq
hemv0/5QrQYX2XaimZhKnXj7AFf8E6bSw/i9YR/a43ecb17LxwjUoiract2n+RhwjINMK/BF0xq9
8AhJA5bjBIQPaseyFUvCSwwpD/BASwfjNrEJm8HCRCNn8AUf3Z6zGiq0tamRW2PWJEBD4KOQqF2d
RFUBuQhRvHj4Ysou6uH1UDXdDPcmIKT/tTkrQhqWLIMzDHtEUCxNQbBcBncpNO9WexLShKSYmd1v
WB2oeNuXvkHGSA7GYYF6QkR+PCU7d8hxxR3/ixS4J0ZEx+AzhU1oPmtu0Ym7wcgo9tfUdQvDRMDG
1+/8NDTM5ZhbP6YYeIn0b7kQkkraY/1xlC5Fi2V8PB8vZKcaDWVSb0H+/yKlC0yw4LYqDKf+3MCK
OYyZgImQEfR1sinU2XNTZ2XkfHZKnAU5HbiTIBtm6SF1+zOPb2Ilw0JAlqxYm1vdNURRdIe4rms3
SIEQRuoiSJUN3dqHRZlhW6mXcVRWD3Zth4nS23EDgFgDdYcaATOki3mlo79UvKBa+/tuPc48067/
HfvKf7tR9P3q/ejXWOMrUCVk4N2L96/muohVuGIvXplAX7Snd7QQ+8QMknfjHeIVV772+JFBnkhn
rKh5qpJiSce8csI/kTFGPAiIyyQgvu/+P1MVFcjSbkDFO1TnNWKKj1J03fHpQX7bsJp+v/E4dx21
9keSqfNesHZYzjpPgGo2hkFykPlY0gZ7kMYCyALjCUUzGimwjEojAjowIbCqGGEcd9o0eRKYTpZY
HTxIXOPdKcfP/m5rO0X/SLq3cqNEozyHKVHL5JmDnJcNJbHsb4b/pHunlgSIDObpME4bRTfJbNC5
a7rp5OybwZ2JCtshmEA/zMHStRXKhBk3XkY/kmJvY31KYAxYv3SWiBe3onphWr3yg4KYeNPWHHxX
yybcmoSo5Bl+iN5Od07kT2HjjHBRNmw1SwZaxc5sIpJOhTYGs7vTtvquouH3GZUfFED5VgsVYSFQ
cMLl4M1yDAAZc/KQNJmBTveE47bBWHcWXOWPcQCtGKamXnWtvdK2EuIuWj2eAKv/ULWxXjaCaRlV
I4ko7ivWfhu/qNHIbjpqPryUdxVyNuVQS3VUbpZ3TxuaiTYEaA7jUMHItEX0vX3apwFg8eJ9nqf4
DwfJMhbta0qx8+G3n6pmwyhguzYcttdIpTI4jIWoi+ZC8qdJXiG4lXrPayqUf0BaYB8fkJFmk7Vm
9tb3OWJiGUnki/rQeh9Cd7w2aAE0J/Z73ZF/eoQk6ThL1uHXD49kOtSk5qfM572PVWltm36O8xiB
QbrNs9LY0RHvXBMi/u2RRcI4USN0VOXt0VVysLhxca9aCKmNrQhtLmFTpKoF+yFwvB4/ZHwZKuvd
cAioCxDG0lvqJBASz+riasv1ifOK5qLRqQl5tSgonq2nUOkjL7qZMUc++TJJUwBo+LRhHgcr2xVY
StDbwFE9op/dwmv31dF58WZJOgxfIDg9fGmAaw74jKACGXwcn4kgNMPjyYzG5e0x2M/rGqqQPvNi
dY4jZimFIcMQbE2KlHfT4cIvoIVziqR1SqamHkaFYNTOEOawUVWOpwKSl6HU2WS4QTyOplDyMb3E
JwLbtabypnhcUN1VpTxx/opkt55Ts8rDyQ39+gCGZsnWHK8EMW+6lTb0bVoTHKbwHedqQnbMBSFN
mTaM+HBhkBxzxvDWu+2ZfyuCqC1Pz6+KFFhVc/kBWzlDWoLAA5oktFRzNzZ3/+dpYLPcqmSzIbJv
ZGcORRaTpqvUZ2VwpVekoyTH3bhtntPGMm702kFlu5446OV8WUxuKPzLUZGrem0uW7zO+oEbx4ES
wAKh51iZtjxc0hpUyXNjWcSiuXteEc8s5LO704g9XD4rdfJr150oFHvAbM8aPhY7FJ9QWBWqXpZl
Y/Q+WN5lEg+cdQvAccYVqREloIfgDFgIPw1bzigJjMJ0WCRSCLZIFQN1l3Xiu3wwbeIWWg6XZeQA
tzmrEq+hwCSl5htHLQ0JZEUGb3cv9VfikkXZqqoyuPHZcCJ7AE1JDazhLSfOBTJrmq7Xj5Abyu/6
J/xswkjEaePMq7Pfq2FiMvOeEIWqAwYC+/jkmxUsApX0Tpwx5RgyrIpiBrKseYwOozwgfPTX00S+
wEVXBdo5tbZtliyw8+Rr11yQH38/3blFRArivU/cBWtRwy6Ju2D+Ml/thrE4s317xk/ShGgfOps2
0Os3uFC+8eOw4i3xKSDfVnGgrKRPAC9j0fjHELQWSCyrUWua858p41yQ+3Ug+zQG3FQr/OK1hR0L
4P1Z42u58UgO5+z7Yz3HEfa4gq4ZH5el8yrklLpyAIgVdT/NkPpgbnXK5iCu3VaSB4+hRSQLW2UG
UwBNE4mo8tma7YslxT7jR6OllOhynJVpeBjKVLT697S/iHFfDo0vv33dw3XpjZziQzNhLLQV8czz
nMLUswQ68piQAZvSonuZvUOfKWncOFy/T6GWUYVT6WDdLQe1L2OshOHwUkaZ0oL9aThl9c5e5Ha1
nwaqM0nFNeMPvJ6ou0OUP49SgkrMsmG3PcgzEqe9Efp2YwTLPfvN8HqfHS/nXdTdBCQQzVP9Y9Hu
chuX46blmqzr7myL3/BZcRtk2tU4qnSWooTMaifxAOXHYKTYRp31YffGTzA6f8O0l746HXUQMCei
YdcUi6Nq1Q7YRwLHR8AKDuPU0a1x3mLhgApcPoN7EDXBp4qtTQMGVwEENfz54+S2bQY+W5yfxIjZ
cFFzu8QtACh+AK8C34R4PI5uD2Pj34JyuN9jyBnermNxhjegMjijKJdPWS8fwHjDer+QiAAbhNbH
7x49XSmUA1BMv6dO+89mQWcJG9Vy5dV6PQOtcuFQs0JGnYakIsOlI/3ZRiisRQn7K7xHHTC1avZy
ti0JsBDLaRwrVWqemIkLf+6T2VaOuz3uieE8vonDIO6OeUD+w0OPMCwRDySxIxR5EV125J9/Ddkv
sPxOubou9tQZgFjSrIEvhBHoDPZfKaCRxf0NAPgscyK/kywGNYX7gfyqSqCAwZF6wODAr0qu6rxs
0533AYRqC5+OTPOHaH8HbpS9ZM0ivUoUPnw+6zEPKm1p3UqW29N+ipIGled9+EEJ1bovaeLWpE7d
eZ30hkrh1kEA40oYEtAelIv73U9FbAVc52q8AiwHice6Umc4G1W/PT8i4THTQDH0/3W6bQNYpozv
jef0pLmsnVxrfptUwpST7CSONnatmoFHAzl1no38GnaaUUKfpGrBrTDdQ8ChGn0p0KZbY7+O4tUv
dDJZs7PKPmfvq9JHdUesAsGXNtWaxexALoVTAaaPQamBfCKxHXANRotWISC0CJ9S6MHoKU78eb6v
BxHDzV6CLmXSD/PQ4s/rwE5sUi5HFBB7Yghbr0/3DFu3rUg2yjWnkf3/gLHcau06AteGAglquWJK
u8XBu5P00vnfc7im4TDRAw/IyQxd4YrdtLhdv6vgSOF6MY4Be206yKNEid5PKewu382PaJC7wF8p
Dvf65Wb1tz8FmiAju7EdoWvQYbIFp6tPj1XEgwecytURYvBNoIqRSF+yn+QJF/UqUFIKOPj4WMWW
zVjwzgNWYBwhM2Pmx0+PMCfZHFHPLl160QqIYHxEaryRv7Tzduj5wA8Z6zOTwzYu3TBjBsYwh7ys
Y3lcm/xImRYUAdh4UwR8Xumw++gFrnsIK+Au6TKNpuTf5Hq8BKTuYU80p9ZQYr6mCyuTuxWKzsai
IBbTO9Otp30yUCvZmM6y6opW/ioEGhrjHPEVU2xq8zgMKjeoK6auw2zKcErWeCSfUqhJoQdqFxgV
LZLU6gqVEeDJS7G6YrX8Iylt/2JOwsKdSU9mNoz28iy8S7nMzVs/4XUiWuOIf3EL7cRQjTrA1zj0
rIRMYCb5ezjS9ePY1Z4WLGYWYoi/ZOvNICmLYQCsKW8g5WtnhFepyN0vd29mX5gJfx8Qr28wqmFE
OSWbwW84p5qTQlsN02MTq+8PTVgE2P0nHRkTOcuLfVo33FtI8yPhlf12VWH7YE8ER9rlF5WrRCas
6cufYvAybZeDAI3JUfjjnWJTauziNQLlp30UzcKuVdgOUoH/nOo8f5NpfD/4XD7Jodra99I8c9tx
JsaBJGHLrbNq7juEXqTkOIk0OlvDf/42UZYpmC4GyRt1iN/qh8EmJPKLotQ/F2FwVjJP077q3BP8
gLfp5KIDt85lVIi0/jnnXxX5raTwm3x/VjvQjQJdzkw1128E0O+wSYRYYWTbLrJ207OSkLT2QhVB
d03iF/ATuIjVIKh0sr9658Fst61wuIz+b0XvmW22SDbqCLsRJIvrY+OuYWIiAZFQkgIbuOkuRsPZ
qg5ggtkDPMOvQPIhUN0sjJ6tyRBU1ooFa5HOV3G9KQOjLcTzt3Y7edtQ1kEnv9qbGnh6fnYYWXoh
JF2tFVWJdahto0S2pMeUQcTUqxhMenHwbES6cfN2lAWMWcrRx5ued1WXeCBCGqKQuD2x72wpQYCZ
gKY8RMycZDGNyWscOP/zJPERdPbLqok0rz0mKXKbTWtm9rIZ0PNpUNexgwQgfg/qSACEH3bzxyuz
rrVZnqRADIiDbKnf30ePqe2+EmnK8u5igbLMOHiF/YeFZqSaaPzt02hMPAn8BHPu6Gpg3L1lRAYn
2tzb1xxfeScadczeL5Er4j1xLhwoJ0PUVot+lqfC7/myhIeNAtLRq6HI83sS9N16VoOktlzUoAZp
6kAqOfavBwh0wjPh6NAaskN0f5BMwIsUfBgvB5naRp362b2+A5uk4idWQuNsBIj0AlVu5iysPOzw
w29zK3YLun9A2DcORkPVi1sI9+5xFNyVpyHgc1ifRHm6+hFKqJ91tHMYbNNUupefJmZf7reB+Hi3
Clt3xvXGgoysRJGMATluyqWs07wZRY5XC8P6SfMaOohSZq8Tkx3ZHuBIyxgWnmpBYdXWAIT6kuB0
OxJ2ME0BSQaZzDAgmMoDx53NgdprfHrROtB0ACgT8bvbHNQgPtrPNaGFMx2tC4RHd2JkT/z4p/KQ
aLJqYnX4UAj1vWq9e5zbziiUVZH+Lt0bukuN7sBWxiPUbM1E39gzGkV85k11SjAOLmZdkx96IErp
amk4HIIjOt5Z9T+GV2qvwVkriYu3oXqkcDMuD9uXnWXg4S7lKg/SPd5rTbSDtDMYtCUMxp2xRrvk
j/DlcgvZ2Vh+oo0fCo9zDk3dhfDuTgMgdItVaP0SDC1ZPczdgGhdO07G1Fg8w2C+Zq+/DoAiNjBb
nFOdIS/G+QpGSA8wlLilfykaNsQ0QzO/0yXo+qmsiqKP9I0dTa9G54IqbgzKJNUa39MO3T8QUxc9
edQD0GXwY/aYV/wIOcyp/nGvOG+MBQOvlAbsN7He49OPnbRVVlRyNaFtt4+FDOMMqazCp4JPZiqN
22CcQWo6PoYyVtbSlkG4giOiMujcvz81KOxRFFDBJdLen1bcc7gqyp9nw3gCEf+V7HkcpY/BnPrp
Z9iYOaqRWIPfFY3IFNjNZ1Ua7cQ/xp1ycDjuMkyjjWFW4Iv7H1cwXxlJotEBrtF4KerGDpzjdI1G
+Faea+0tkKK4YpKyRcbjpY7TcGIuNIo+9jUQA8R2flQx1DjjiUIY+6upzmiFcLrsbTnT8AmP3spg
W7/+DuRAtsYCEtt2iKVGoTPnjDgILpYvFelnOEz4WWKH9uXVI9L+E7/2Mea69E8KIkhJRr4UMN5c
xHSDHtNz712A/oNAAL8PzWu57NaSYq+PK/JtIshnKQOzNmmu1d10Sw9zKsMerJdrSmMgHZs0stU+
a9hL5gqzMAwByVgv+CfBa0GEKlLDwetGQTOhy5w2o82wW1Bxgqo138qojvrSboGsm5StMl0uzKn9
Kl8cNCD9boVbQ5vKsPAOAqA/2eBBPtCEQGVvotug1W3++4rtR1emcfbX2Wv/gqnEiLqbsiqpepBr
b6PNpkQgOfllZ+9diyDz3/gwt+x9xzcZ6a0NFePtE+cSlIYJOgflZ4gIK813humTDn6UrU1s16pz
vUwp+dJSRnaefaV517O5J2ESx1LZ83HXh+LkYd8Cc7jLdTXFTB+UfQW7Kk22o8hzE5pJuxzWILE1
yUVQjmsn2ijBNFqx5LgX7W+xx6Xw6yymvKUWWV5P0+tfTJ4iKT+arUKZFw/BxrWcH+vfTjReO+a1
GkcWk05NWRagQeat8mfKosa4dCkZMEomtwxhN0Ayg+hcQjYKibNHDBSpuXhRwc7DH/xur8DcaZxh
FEvi3ADKLbuaZeumlqcGKYFNQFcxyoDif409T/+8wGjve1ph987fXbNkdc08HhVy1GNJ0LRJWH2z
LeLX4IM0ZgsY2sPrpnKiT4OdiXmEiAsKxcrsclxdUVQScFOQOocTqv9cO/LkNOiVUdE1N+5bH2SR
eMN8ZcsDAIXbc6PmKmeG2/DD163G/Wx85MqrYM0WF7OYueVuU3hTf10tGzrN31tXmHIaAvJMdLFv
aDIwhck11CoDV89htz1L5tWIjzzfnRy8e1cb0z0dDDArUxle0iJeXvUfv2pcxMyq7McWwGKEhJRk
Py6ZZthKJHS7p9wXLL47D77mEf6+gFnIbdZ2A5af6YVFX0o1A+h7Q7uL03bHlT75IqaWgurG1BlU
QNQGj3gP4hqtqTt1Bi3576Kyo0J+O6oyxFkYWxWZBg9baD+ERwNWViNWEQoPhe5f7ZvVXGed0t18
6nwSzLRl/Xa8y81yTxPC4KS0R/DmvX0PLfSAsPdEgMD2P9ZIUN8tTo7Q/EA4+YYmPzIqC/B0P9rR
fKYm7US6Wun62mSrJwY9vRCtrmq4wDkFx5w4gFo5IO77K8JiIJaejQT/Med7LF18qzvyvwhxHljd
XkMhhbPcWi1tFAV+aulc1YmWTMxhywEUvCLnH0nMASzGT1tTmDZMm9bYlD4Opkm/Lrkb+vwGeoT5
eVu3+BtTm5VBgCALQUAG+Y/+yZcjFl+8PicQQfLIi+MWk0jeo7d8C7d3wtcOtZ6pGkNsCBmRI2tv
T9JffddzshO9em8gSTQzd5y+vipKx+wtgv0DS0S8Ww8JEe1sDbNHi/zY1EjfqpFkT4bSWiWVE6y6
p9MF+x3bULdTUTh+hSIU8qNf00h0/uOC2URQjHdZbuYfPZTnCN7s7GmNfKjl6qJYS82LVDydMPNo
eq1ya3/8dfvHaDJxNsrWoH0YSKIzyxFmZhQ+KOLlFZvaFFCcnxFmFpfaFku7/25+ynS80H4NM7Eo
tpAPe2GCcofi2l0VlPYIxSVLA4FqdbFcGgA78x+nKyu0hFWGYFbbCDJdpvyt+u1mvTBAOyjRtSmo
mjbIIld7ZQ6wefOYuDc8YqfgCm2ICoyUOrxlwTTt2/mEkMkhzyRs5W7dv7rbuMqHgCTETmWSsml6
Q71jt9pNK4U8N41hHispWRxJOIuanKbSrrCL5WKDtVUwlPuOhxpgiUg/lTT70OXtMFFML6R4G122
Vimje+vQJB/NYC0q96sCoors93vEz5h3bikCWeL8TBHH2Kjvfcz0PKchROgweaCInHS4Ior84n6L
y4Thsb1mdChMYaYjw7/IFJ+tJK0pgUym/eJMSBtiqiiz4aU33M1rkD1piQDSIibfumwRS5EpD4Pl
/PALXD23rUPxEpM3maTVa63QePLLCXjY+GX9nycuHy5KID8VvudR0rJRXmMyayfRfrI1H+6ca9lx
37AVKcQlgCN1ZIBSIeyj8Kak/1+eWpgTxReQH+rZ1NxcHd2F5XzQqLllNazPgfKXd834d4u6IpcM
sKEC0Zc9k32OiN1JT9ZRnJxrFs1jN9s/ixgVuuwvOB+nT3yg4uTpLIk0WtNNFvmOml0OZXdIz0OP
lrRCV6tksmL5ObFuQR+QqK4RqqNcsIwa3owDrESbKxGakyPk34eOl6OuAg4gAjI3ePdczbvnFTJ/
3OBaIRdzKiltMWqz55JoBWMyb8+iuRKfbRA2g2iWbg+sZrnF2FrYyroAbAdjDO8pA46fK9dlWcWX
S7BhhtT/9N8ATtnP1A/1VAw8w8r0c8LzK2llYzd8ufPV/qgW/jhZRm3ROVrSoO+lilgB/6w2e4UW
84J+Z4dTrZkWPH3w2nlRPoCofIz/fMdIOb1FlAMBRAkTayNVwqJ+5XEMm5O2Jvz8vAKTQb6l2QKO
RyN9RZSxPilhz03RGNEFEO+F7tyA1zvxwvxCDmhXLavJtpN3+OEhwUsy28d3GZpK4eCtl8GVsQvF
Pcc8u2UY4HNGBYRhtHhKXQ43tqC6F/GPkNcrELZE4qq+44hQg8f3P4trTmjlNpCkQuFt+C/yv/Ul
MzDBKtw4w8BlVlGNBfJ2N0CaqA1v2mRocvS9joVNTLJl0wkLlEBXBJTPYKR1Auv10q/kHBbtnC9l
/h/zwXXWBgkqALO84E9jfq1ScWOsksGawkScmq6Y5VSqwnnGFihviGvVRlua+QBiZPYgZ3uoSxPI
kaQTPRPNXfpc9yRgYL7I/7GDb3oqrUxdqW0x70PCTNLv8w6xz398HJ/6+fNGcyI41F91WF2TiHlJ
BUR2NmZvUOIt/+Ky/4YT7S2KBg0kGelNSjAciN/A1Wm/CkjEi3l5JSXJTHGCFrNwjr/v4O3VWdXO
jcfMQ2eBt8NXROTsi1eBjdGlHSXT5o4jYBARJqLVioT8AMNNAEVbHI397l0Swct7ATgSOcJtDs/p
SGkcTviWJTtZc+6mube7vkw68ZuzakiavqctnsS1nDRYZuTUa+pU5hxyeuStG9iTXl9roIbLu65u
jlHsWqWJkfSpJhQkZ+AaQree9SQiwn/sTAepsWrxsal1N1EAMUIU1VlMltIRbh2VoNIEXrW8WrAv
mm+w3ZeUq2I4BZGwykYtgfDMRjRxjSI/JroAMU02wcMBgg5wMq5950PF0X6CWN11m9pip72ibKxM
iEku8z52N7r3wMHDDZE8bI2mEUppMaxOwyeC6JBSsXmhFvQtq2uAssuScfmRgz/wzGLGi3zTOUrK
CXgebIGgdXrXqXcNY/P3KgTmyxzeBkJwI4Z/g/DfOAKUu4IHPwaLnW1PEqaj5is4/8TYPI6GaAyb
9nypCcrICLwQ8QpbGU1auwi112rFdg5mmWNnkPUbbDOtyFilsK8lvhnQW7Bx+kf9c+egYf3loeg3
rweVo/dUW/gOoyvabqT8GCB9eh7sPUy9JXSlosOQcufnisB2ZOCwON8GxthdnVolu3gTPYSoI2nO
UpIgNLBKN0ijn8GHj+/tUypAH/mlMTH525UfKfZkSAlpoOh1B1wFfTrFXCTgq2mY8ofCjq29e3mO
khd0B/17TS02KQOtgUS6/WV2/tBtTxJKxIYayolxUV5uVBAV91gqrVCuydrqafqdKd+MX/ri+znq
wRf1W2XXFKumiJHXDE1ZiXQx7KGNvcJVMjd+E5o9DpWj+5ryFMtT6FgathM83RjZrwNVQYHtEmOj
HW/ElbAKGTPEqCQRB6vWUL7V2dG8iH/3Ena1p9FlyqiA1gu0GMV3Rh7JVRRpnKzaKVlJmyjtX439
GkjE4uEZPjOZzz8PBB6He9BSX37rlBtJi8+v/ohctlVCVjyr3oQSKXbZiYaJ9yB8lmDhBhSvNga4
JG1mf+NE0cIFGWPh8T4MY06cYFBGc6o12qzqrplToBwh12/oGEEyCzfufNcRRMcIV93ApXMnKycs
qpHCHD8s7e9SGXL6VNcqgDjUuImL9SqL8LK2ZmP2x9BwhgoF1+DhPQK4whoEOdHIzcfK6h1NUFYL
ZOHjHZVPi96TLbeARvJkurcxVdvOqBKuThbpmsY+M82mQmhuN2Kp5Cj/YGXuN4Ms/JuNfq1XT/lV
TyZhgDhp85c/FHoPzsnWXRFwNU3/oXP2lPmupkxZQY350qjk2OR+qESRoDMDT945QVem90XaVqP5
7cm7C8mcy87HGLPn6DZ2y7ZCG9DN0+7sP8bEngw3c1l6ARPxHqQaGAiXdF3n2yZ2pTeVGEhfbcPw
HaBg/cxh8S24OjoZjnuNQFtfKgCfrliwgC5hN+fZ6WnPnEgKSgZZ//+qV7HivgoPtO6Nd4XfR1Wp
eyKrOa8Lg6wU0h3D0LpaztNmu6QoaRz+6SbLL9tYf3oyQHs9K6BlzeHNrNpYawGtpjBQnh071dyu
qiDXZPg0mju9VSHNk1Ypth7w6aeU0V3/p4D/+XujWnoAOSpvz1zC0OXdtVsYQ3+VN1KeN9u/OtWg
YCf3nKAgPsBEQp6IOpU70au7z6X93kn0XUh55HzuJbvRrlECqEK8gvmhtCdgX7eM68NTdKZs3VT6
yMj7hhrq+Xenw0gCOxw704kvmf/WspUC1PAK4VCo2ZpUgBG1F4wX7W9+0zGhO31B4HEgHW8BDq/w
ZV5uQBEpNfbHiXP5699FapyWk0B5k9NUHkgsLUmawF+EquEp4NO3TviVABXtgL4oDjIz6DQGvbVw
8JaX82RUZsncJ7il6Wgq8sKOKEgwEOCvpNiQgl8ebAADCgmDd9G0RLp9f50W4cQETngeHNQy1tsu
eRUxDUBSh0yF9BXH+XbBVyvhrkF8E7/Db535ys7g5+wHCGKMldU9VBFP4FrsROe85G70BPdf0mZX
DnjqhrIWle/AJBjdvjr7PmH8JCo7DcLWiegfwKfPt091pPyE4EdXff1PHEmFzbnzV/3Cw2CDxuBV
NUAjGokl/1SQlcqHA77K0bKnzgvisoaBwjXLq3bgOQNXdMeQdkYbg+EQGm7lvVcnw9VIWK4dUywt
lBj85ZB64ry4nbiWXr0vQa9/flUtO1Xcwygwy0A3lYVTZz4chPnxxsjMkmbPYwS1SOVkrHs8jx1P
MRgWGaN0TdDnwTjOMmoIhvOv6vDJOPCAcTKT1L+redrQu1Qw5klLr+kb1WoPOtEWPOb8TIaGTtvq
GcVtc4Serzb9swNAxzD1wKvOjQrUVUkAH/qap57Z8Cfa1EhCdQBSQKg/nxU8hNmfVVqOx7Aq1OQW
aZPB3bo2tuAn/tMEB3Bylj2j5AoNey4h+dEc5VgD1h4zRiQ53PKTbdeOWAhS49fkPA4NARToGJCa
IiwGjwuLNkWJaWFgoNugnB6/FfMSsWNAZaESJaR1wKx8yxVkFZnkgQ54ZIp6X5PUsIIQi3g5DYbE
F7IKD0L4HlKnDQH79gIarXI/HHLykvl4o3YfWb5/bGPIEeQTePxj5Dyx623pRRM4xjIrl5WNGCa7
SOmAukDVyVvk6Vyoo2IOGp6xq5ldOMecvjw5PXUMFlG9SKFJJaWPmLAS+/odI6Oe+j2JfLOiSMkc
oSKFzfFZnU9ms6oqCckTH336/3bL3L7RXhMWu/59y0GKXsbTRaTMrSat46zI0JKN5d1ePbMmGK3d
xsSgLVVJRb5KKFwL/PVESjF/RJ0EGxEGcQaQdLnGQU8nkNT1bzBPFkpQ4gPIPgp2fYE87XTHvsJq
oVB9PJ48C58cqlp+gqjDMfWIQv2FxvS+HkbN4ekJ0sFpi3vLGuxYYq7LMbTGzznYBvyQWZmnEobE
JyaGi41mtjdk0hOYY6ff/evI0m05VCHk7dZWJMT2Tz91oUJcsIgDFZfbcB1wEP8rxGtuPFZ6kfcs
IzbrQExelzQ5kH8auLl6aHNwNA5d+j8B7SI5e3RWXIIFBAuIOetXTnC7IchT29/CxIh/IIhc+VzX
J3qScGuWDktyZOqM2IUzozsSMSPhSjmIQubiJw9SNRCTJvzu6UEF268KsKLqBeJ4UKi039vjK6wE
wHKwlrBWfmiJRO1HDDdtQB/OnINYQMKJLMUmJj212zMl7Qmet5mzYcI7BsVK1B9M96mb6MxTxH3u
UPqcbmPK7CJqjqy5w082iqxzOIEzUQOZHpqaFQxiSiaMsOD9QZF+3EIpOwWchAskbcGKHj1wtMFc
eznvnDdTtQJo54sPEytSETvASOcPKUjhORe3OHpFxwi3lis2HyuUFRJos7yOdqhzeghVwVul9CYI
QUJSq/qKVGsXfvpJkyHSxtSd6Di+isQCQrrkm0t75+X2OgqkZ8qbFGRlZh4q3NOJb+C7QIK6FRz/
NZY1JUS8rXsff4IXKGBGnuCd2n9r3hNQCiaGT423AAbPZnj6LysvYoyCYje+vaYNFOrhrzHUTCkg
MjaDmGpWuNXH6szOhYXFCVtO4GCnc05q6lLxvWTKb5bKfFY60kIUWjkjLCqzWQ1yMomZCxZpScQz
mrRYNf9kq9+QdTLw6BfpJxt4V6V5zZNEanIYYVvG0vLR5cyi1SAZXUckn3hhQ5KiiBwW1+Y0XjnM
bLiaUhcveWzb+Cr6POS6oBdodqYqUvhCY5z+GVRPGrj6YcrIty1AzsCkFgY6ZEsvij1JlhnUI/Iu
RkmYumYte8kin1LNjPZnEwMKGEBGpw3hY1EF/WuDhe6HEsC29uLGcbgvEzvZWwFFmuYQg3DYqYmA
TESn0LUU3ejjymGscPMrNJ9qeNOaqTnD1jk8h1zFGdrZbpaRqztHeQTmmgsl/eCcvnLlZq9JLXul
qbAarP2ZPlcSOP8PYyjEzTzpdrO3HcNnWVQj3fqw8HzjJzZYn2PiyD8kx4hIijlUj3EhMZlluJYp
lCgGGXuEslc1dTlg975PVFqTb//yi6fiKLdaw7MUUeC4JQH1BOWT4gek4+fCgs2KGe6svUR7Gwmf
qPNNxSGkbfFdjFEnCzCjpK1Wl3/DEBgLTsPQcw93y/YOM+jjWetilNL0wXF32D5O4xUR/8kcdoCd
sExunCn2JR2GwxOV4/1+b9PgpEcfoP7JW2kv8GHnmf0dRB9JkG+iRYSnxyaDzVTh22bBpxNqUfWA
Yxeu/OAIvdTaLWVzeRHT2VbVHFC2khoFRRBoFtEDdcOv4UbwAd5BmdYQW8DyIUnGyrHmoH2xXQL4
KgEf+SEtwyoIBaH1GSCWgAJUNBwTxWqrU/8aL5viYK3mpf1qt91tZYLFzOoX27a7mj+waeSbJUjI
OGy2wvv4baEx3MP3ANuAfvmXZf10bBUuCClsrnTRDYueqkdrNY0CK4jDTmRlD2z/jNulk6LvDxhe
ijDCbhYiqNVzYuqB/wd0JSttGU+4dpiQMD9TubZPSnj2ZNRIHTXH8dAZ4SBh5ukvXoT9oiIfttmJ
Edh4JARw6qLm4ETTpbW0EJYA5D8hQo999AWjy4DMb1959PMww+eU6r1QYYrx47fZq9UBy522TmR6
TEVqKFdVMz1+PNeNZryOQ6h1xB+5D2nIiww+7LkzQiM0O99hgSe/1Gia2KPWde3Ro7TOLYk2JNkz
A7tNCEROmD/ywJFJjmfJhXpo7F7HWglwu/dlSuG9jVb56aMbGSRdabYMeSRrjC/sR3EPKJU/HKXg
vVXJ4nlnmQ5MHUx+X0etO7G99EMVH6rnAhUnAFesrfLQYoSyICfi5aT55dPPc4pnbhG/NzYhi+mW
nFORW9oWH9KsFs3C1AL2fpVqIf8oMf9OK73Jt5GAA4V0BHIPtl1CBe15b1t0vhM4Zwtxu4qjHwqI
H5gdumnR+yj5VYacJxAzet9IUtNDAJwgelv5lLkOfhTMwej6b0gKQSxytO1Qz3dnS1PQtjweQwT0
o80QixFlgv09qtAhi8OXgOXzMdBhsgacRn0zpcrTON4fDkhqYEpyLOqjcezABJ9nVZErzg0RzvxW
ImwJF+y1xYycONCDIdl8BPGjGsJheVz5We97BohBt8+aVAysvuwndiaGRjKUDN0YiNXTVIPkSCKR
Z9D/yYQWc/bb9OnaH4prE6GRb3U3hESQtOOXl3PgttdwzMrvtN365sR4rBQJn4AZ1aqyHJozOgdj
ZDk08cvMz7t3wKO0nQRSYE7Js/f+p8H2uTFVgAn96WfIuabY6IwKD476TzhP+EQLxCtl7pKezQnI
c99y3oHEpRj2dyH6yxxYIoVQWkNDcw0KjP5LrcGYUi27DMCWNt6me7wc2SKBt6yNI7ESPvdhMs7L
96Pe0P25vgKaqn5qLxrUIRJGWL+lHMWVYIsDsfGnqxZBVgHMg1wp05uGJTg7OgvymSDaxhLn9tcz
h51l/mcW3Yx/XOPzXJyTRdD5Thnf2TNhSAFdCmZe7ycjxM6+mcRhTLN4+hFyJLSWZnqRzOT/mvKG
FT4lDqE+wu/zr45gZEik2HuK+5TqOK+9ys1D690P77OGTRfCx+Ay8/mt1gqCuCc2ZJxeLUtklVTn
B5Y0UBRLLCUDrFKAeJLvIB0rU8aBYd1KOcxzBF36otyrmW2JuHsneKT3gaYU53XeZ5WpXjVfSdFP
fq+TjfyR864Z5VC/HY3OAlWEms98skpDwHyof2UaFbGKBy7Nhx3LdxYQfZ9AFpooffDa1X934WAN
+WrWhsuls8/NJomg8WaDgeiA5hMnlcuIRF1YsDT5J90wDB2cKDemWY/Y8ay7CW032/v+XOqvwxBW
2A0HFV3TZX4dQA5NabB/UcyI3F+gpeXdLaUCZy+y/bJ/xVu6Yyz+tFY+XwGxRrvUQZTWhI/4+8ot
XytX6GsIyjK4wEmcCpH8Rm+gh821FFIP+sSAMUby7qoY+9ETUhvvclHsIzYVvO6ulELzq7oChfmw
P6cM50rxvRW3+cPcznNAqLjnPta8SZFKS9VOlN3g3OsUBYR9fYgRIfFA6QE1BOlKXqYS8gwZ+qVM
TY2HIFo+SiHjPfSrnSL5kC4jJ+gs7mnYvYRTUEFNvl2oSWGSWOkI2pFAncL8mh2GmEH0PDbBJpcn
Bn05xn0TEYkmXvuAIqmb8GQJZVaY2xg0chXXZcfKRE5TS4/Mk3YQVDimu8btzKzxlXreDt3/nK+O
sfp/ZRHWjhecJgYZH1AwJPb71zaAFEnNpYqbXbsqxgNF7zjXBBPkDvBQMTPreHnsIHq1B6smHpd5
GZThzAQztrQc06AHtVTAn4YXgPRNz4dL9tWXqOXCREfbrqdJ6pXhMl7/mDDYFBOHe4NMGcHFWgMD
rBgZPtgHG52FHIktkc4ZZ72rhccApYLf2ZPqMrX2zIregbhRRLpUMLMAchqAy6mU4+aCRnktFy8v
BtSGkoDRGTmlgR1uu53qnLU95bCsKG7BUe8JNwjS8/17uy51aYXL3Kf/X0+JzKmPfHW3AX/BiWfE
slB3gE1W0Ohq/kabb0MZDeWBBaW38NN5UywfhB4E4jcifjcmI+XDR9ZQI7rUZ1n35pcx13o90wVQ
0QA8bZ61nmINrR2eUKWoYNwKiltPsduq3laD43UoGGdgINWrUBoAtvUIOXNtAxDNSa5p9UKg/cNN
RWtdKGPYQTP3nYuIMvTUobwV0793f7VbuDxiIDpSxF98Diz5W11O4M0w/pnjrDZFJNo9jRevtu5a
PnCuixENMbjD1dt9lm9278TUyHnmiVg2O5+yyMRK0yn4RmDD3/LGNmlZsvXhWHjuU77CmqOqqiFs
Qu3jnpCCD/wNzDUsKLRiAJKPrdrK1XrWmGgVV13Rw9qzlDjZ//pLXPrOjRbRguwAgQvSgVz0UuE5
P54wApG5jz6A08F771QTQyt812lsNrtUZkaPEvqAhNQmobFC/0lCnro+8qnd/IJUi2NNL1L9e2CZ
ogxZHpTxpqPaWW3cQqMoV1Qn3Yrz7ech9Rj90241gN9I3IuwXwol9oNBe5JlFFxXdNXQ8mOZYoEC
ABSCceiK3xn4mkxOgdJMjTd5/iJPHlln0TflD93W0VVbdlp6L3oCpNUvdeyYRU1CWJ7WjAc01Drz
zA1SPeJJFs1t/+crvCKTNC2uwywcW4vRNOtxEPDrfub660w60QOlNPFMInMS2oiNMF66bw9LwhmQ
ZZLmQ9Z0vqMeXnkM4LYwFME//HbR9lJXmmMb1kc8DJRSLn3gPF7yvCz+FUwwNvd1aCAbQCKaD01d
l+L6j+dGjplTQ/sL7JowD6m8YQbjvw5hd1seKTkiYnFJkvt0jiGywR+drjsAmN6uxPImUi5sNDbt
bmfO6/bJ158jL6ZE/eDqAdw27PQCx9T1W56OtrrNOK/UT2XN89mOuLpwnuPQX4hQP8A1gmajURcD
HF23jrMibUurz1M26wPcP9fNrihFo1Wu7t+jjcsiGcnu3pHdyWXWiHCYa2FnbCNHQZ/F2QqCVzdI
tB6yda2v+g9GqWtCxIkb6Ekx9sxRBlDejNoXReGVVWYebmqZ8ff4pE+OLmcmOCmIeSJDk7a7Svk/
MvnJZfcTlIBzJJh2FKBRjLVG5teVm2zZoWYPGCCRAAyZxHbkUmrAi+P3Q2LtwJtCrCe43Zx70e7n
fFGMmNllggAgsV2DnbBOzbJfpAt24T1t9EOh7PlS6D0I6goTSMVVRz0UTkkRKT8rM6Sga/zN8Alf
NqeXhLPiAJWRvXPzHLlSTNyrZXsgAsj/JWKDYFWMApYs7Kj37gPQ/vi3J5ORLkhKjLxZgQkhyeIs
vkIIUn8NQQnf2kMzXXYu3ssSC/xKidzfyFEvodF6NN7R+nPkkEw7WBWf5nIaj3GBmv8McWI68PH7
6Lh6QKyxZgHPzXbbVZzh2aRL9awgQYkReUpCGGwvbp9H3y/v55nztD7b+YGM1icwqtKeLw7z31Up
b7Ke/WNKlSuhy2wgsmdpytbrU4OIS7wokHObq/ygTB+rZzsPp2oPYHT0RYDJYK4240/vmeCe/Lui
Qt4j1FRoMZfc/3S4WUG1IJ81p0XTx4wxqoozrsmRgIUE/9bQrlPQvFfRjxn1gSgPN/RUB0xLVUDK
ZXLVXAc0Tsc4XbzHaC34Z7smeMhU6xBr+5iZrGhutrs4lbS25G74LVmVB/e/BSk/p8kq9ZvtpciS
Us2k2QcsgxguFgr6csLfXgw/aNJUV9e03K16GJRUMYJzCKbi2+emvkaFoJCbROhMXxlFwNVXwZk0
KUWQBmHyXgv1WGZOi9NuRf+bajbYPNMQYijRFBrFFgcaC7TnfW8+UqFrjJl1CYQogJPJFJ0G5k2N
1R7R5cB9FyFs/2BWG4eSszJIhtwndaL2C3PhSI6KKMWXeFPVVjSt7s+7LNUfv4GNLXZrcEBD6zYX
46130hKScZBVad+AzK5Oof15lC5u8DaGhUQDkZc7HsO7rWjVN9xNDXgelU5DBjP7pNIQDw7QJ3eg
VqTQUJjpFotVs6EPNuWeWKiODiOKYUkXonr6DgQ42ccwxueeUw1nQXZoxFOZubHccLyv1f1MVVA/
ivwKEmL2r76MwLU9y5oeUsix7X1S7XtCxzobYyFXgiAXRLWhzsXxm0AaTH4Ywp35t1piq2D4QTLz
a/ySmlVA5S0ZzSGS6tCZJ+S6J5bbKujEkZmr7hUkvy3j1JHrOYH1EnPxBMenPqcL6YVNQCWujAR5
2l7T3cRwaTkXf3igK/AFdQaZfk+hse63wA5QO8Adyl7Om/9/WELr3BBtKN6w9rw1MspbmrDDp5s4
yVMM8uLX5HYmOEVSPlvOyZ1MDdPSdO4sJaFNArpwRKm8vzWKiHQg37hRb09O8/qa1r30dmZMvoas
cncP2JJtnqA+EttqStgYrlV8Bf243ESXi1M4AbcLPbfKJIjV3dcFtfMfgXNcFN5wBRyoAgeWe6V/
zi41jtD9VmAypVsQzDCwnFCIbTylgl+AfaYy08ibg7A1SDtj6t6YjZgjptwl4GzT2dz4wqJKomuO
f8AAhLbCcQEqH1Xg+/ZJlbUwOWNTVza9iAX7mpLCMcLRxXxSPbKu/uQuuQWloGZkk1mmMRL3eORd
fXIlp6S7Zk5vQpQFkK+a26qm5jdXvMlK7QR8HeKRn3W7B0/iqpYtVjFhb4FLKGRhJr9uBT/iJVUp
FdIduDao4UYr/gjL2+10F0BkmBgMkoxcYVHpUP3bIzZOlDSpXGKBpd+I8P3oSB0JloqALB0Y+a0V
+TC0YEDqJn/qz6Jw86pXg1arRsl8LR4Ir20j/Sb6dfwVFm6dn3FyamwyxUpyDNO9iYBYlP1hURGB
Mjro5yff7Fr0uOKjEgUjSqiNeBIrGfqa6EiCAORddsNFqvk/IEu4ijl8SRYgs7Gzo/qxG5WIuq6X
kREb3n+8FwLtW+ovi3ZD9Cu2cXH6Om+hQGZw5ZxEEk5TBppy+m//kKP9dxyHkwHEJjJlL36PjvMz
Jk3jAu7xloFPSCo7N9KR1t2b/5OfY0W36AqhXiyLNz/32t7CMdRTmj9fAJVHpppHKQVva38fcVqh
s4vDKOAoxXVK1kzfBe8ccUG4z8jnMVr1nd/Qsf/C6lfC8OSo50HUOyo7BrQXN+5Y4pDbHw7ayDAa
+pBI6By0hzvYvdPNJQZxXcBvdEOUuCpw8qnecflmO9T/BI/XPPasr02KtOgHE4OKDKy3UQ0lJs7k
pAHXEfhLKP8ExhxMdb8MITK7K0y9KdWVQAl4ocaO6YpTNBlwl2cFzoDigwyMpHVnXB27dpmquNMl
T/He+XPk5P9zGqJNEuBb6/5LsOZt1fAdUica1BFrywLvUO7L/cnvFbLZOThMUgHI/25CZ5HfOW88
yaSwrc/F0bPzrrQtFUPky06pDp48to43+lTchGY6UZYplz8WVjDoVz/ncJKZmu0vDMwo0+skNpFz
cOCZzE5LtkwZyXG6o/jQ/0UO/1iM2EXN5MgC96RcchSl6yF92RUDhFFlUyDH5n0pdfVDudnbIKmV
aRQSzV2AbjF8ti0DYKuPsAUaASho7GVIfjX0BKg5uqnNT1aA9gzWDgZqLy1A04vPKtgDA51ozcmb
fU6wvHqNT2lCDtPdSMYxndYrchiJk75DZpL7xsxbFzv8+UZ5MOVUmgal4rLsmVrJ1pLRIvCXRcpV
5rtsEAfj3RigvYhkDjKgtDFA+0KUdPPMWM7Sh6AbletuSlh0U3LiJhnyRXzsbrOD835jfIqGrueA
1is0yCqOJzR7ISR/JJeS7plQ1rfx4NZHehQrnAFyCUfRH4fwmnh4Qd18kRODFddmtdqfB4S6lcOo
PziLdTVJ3xN6k5YMPfI/SBFU0lL2Yrmdyayn4Z9LZ8eVQfcCcaaI4fx6pkO24VamEPCB10dpdIhp
G2r1YhlovuJKDLoTcWkBm1X2lueQYL46XL5OJ/b2QVY8mv9phn0Ng/3geAQa/bEyfNMvbBmgWibM
d6OWzv+1F6Zo7IQDXaVnJQMManu6UwBH9rjUMXpIG3EVAunVQRjjibYKeH3uX+3RNrqaOCZPqyiY
JihUI12HOFw0WSzAxSWNVp2NeW2XYVD1pWKbfN7hGafj8by1DV9DaigwVvfDFSQNm4EJkZ3xGixk
wbmWnGf47MX7vBE5VFD7atHBJtLczCQDTYv/6q+AW1yk/0zKI/s907cT8dKAHt5JukWHyUzX6oDb
javE7I4cDCTE/mf5knFP6S99DrIH9trL3gdIZiDuEn3+BwZYlb0rKheM+hD5Vy/aYXVZ8AEoTk8H
bQqEklYtLk9wkd3a54d9PXwYJ3lKNlETHJKNlsMUXWAPbNPWPZiEDPvMW+1BAl4L2UXblAl5mlpN
DSAoic6g7+qwxmyUKHYYgEpqqKbnCeYMIgfjSTlyfHEVROwXY4UmK89eEp0eKDMiEa2W9yyX2rnw
KrIofAmtBvLADMeZFqhHDOFhe2bZ5018qwdt4/DpPQwNbeeN8uuApEFHXxwx11VL3fioUsVvlnCw
stvcqAZWeFZRgSD9vdD5DRw3T9objGUgQVUeYyq77p3BI3ntQdTgg8hcEl423BcLG9g31n4lvoLQ
UphQ5Y1hwiXsoiRLVXa+DzdUQ/Jep93erHSGcxYbUcm4INCR2rcVw90QVxt3ROMLG8yaAjeK8T05
cJsPoCfpIwzXIq5s50KQg/WBaG8AomqfO4khcOQ7VY5gf+lgxnxsNrLysu1Fjmjeog+A/qh/Y+sM
oumFRdvipcFtDgaB4+DF2xkuEpIY3mA8mHMat7JCiUN/baevOBfmUk08g/HZJPO41dwr1mIglzEn
aMzD1upd1Cz0nmi9sx39n2k1oahKuJGycf1s3FhRYTvCJDgvKpUk4zN16GAtIKCqGRf2GiRjq1fR
v/XxS6vig3hjgnUHnInyQUt0LSRNf7UTelLGMvRV4r0jytazSTT0anNP0EA2tIa4ZEmxGNf1sBvc
1xQjFmRlMyEZIiMpt/3q0zfZ2XZ4jG8r5lFX1cOko8e65wFTKiuKncLt5POapil4QOjGUrZdwGqA
tgR9OatWVBZJ6xl00Q2zoJ+bIZh3jdB3NuhWmmSfe1FVzMyd+Ue76S/qOeLRpDwfExMfq2zx1Sqe
D0O3tmkE0zEFc7qpqIqiJbJ/rFqIVfh9YAQWpuZDXlojJVpYi+gcMaRDueQnLiWiIAksXLuHmgiH
cDmujnb7hHGHduBFo+hDaU0Ue5bgN3ieuIEuFuJI3zeTH02bc9FtZYEtJFhPCswoZqRlcQsPz091
XzGv2AFbBPoHj0FwzV1Z+XkHHDGskiYRre9wsfII8tDfpo237+cw1ZcZO8I2ZZK/GwjFGy0PMwr0
q7aWrnsErkV2YK93tNuhp2GDLVV3wURfGGT9lAyAqvbn3mrD7O55XOnmmeW+NqRqO32ZdAOu2oWo
+T5ByptygyAywaQDRjkOuYNiKi0IaxIfu5aUnRcvlsddxE10YfSKqlSTl1qHgmrqWpmUnH3/WOQU
g/H9M+X9wuhn7xlDLukFauZBUS/iikcElWZZ9MAENsgMhwLtSyX/LrElnu0kf7B5Gkk1juuRLsiq
wOfL9bgMr/Z7G+VKleVlZBgB2b0TPiuzADpVzMdD2gLZa1gY5ANfSFLW+up2JtjXrSNwrETmw+3L
5i+44nHxUM2GSr27GeMKLnIWzKrD1Vu0TNN/e05NvfKX15UcmzdSxnzbGCiGgQcxZIpAOd19IcZl
y+YT7zY43opr5vi6pWTgj8d1UBqYqRj1E3kr7Mm6981+gPdxfEeF5g+OrvZGdrgkOp7Ipbd9miMJ
g6XjXzOUgJsCbbSXHqrZCl+7GRaNqWWXp+61WcA2gm3P0Ka8i8ROYUWfNiHQvAg7T/3KoI6fGB7i
AocDeaj0lTtHokEDjYahpdKtSL46n1fRC+BQ06kxFep9e0vewoSkzV66s45Dn5T6+UeOcwgP+VIw
HjGkOgjDZczwHv41EsKh3Lh0WGHmldcxMB/iAQqX1S4937zTPNgNsM0ITpHUT+B8WXTjYJOJ4P9N
TxmIIM975abj1tGg1B1Cts/W3IGyqiWngq7HfH3lzvDsZOFRIaAHdp0GqhCi7PyJk2L2DPUJ8aev
o+xxjBCu63ZxUuOJ6j9ttqU7/OfdsxafSdZLMFfR/YT7+CxsUzS/lngL685l9m9TH5jUx5aSqJBA
eocWKdqOjUNcgKyvGJGnD2sIfUTa7abs789CK/S6AViA24FulgZwNCPyzogVJqMyeBWofE8vYrvX
kMkUHN4rFn1I1I1TfObdJQ7Lqbqu/m3ReUjROPJW8+VMt31RW15Ooy6wlL1ejeDDc8PVvjVI9xBR
zr+7DI4P7HscO6k6wwaqazhpB7Ih8JPiNBvLkaLF9CnPwLX5VYitrujvhpFT5Ec7sdmaNNiZm1dp
52RRpu1Cg2Gy7NN6lb+cNv9a6TmYvuwriVRWqn9sDpnC63Oe362tR7m6I3t0egfScIWXCxwMawcM
uyJWnk1iYWoiZDOIqDevMMSZOKj+XCRyaF9HVqkBKhZMB9y7Ixc1kk4zAVqFx/DW+fpHNGuFPeEy
Gc342vWlgBLZynWiDF2+lP/lE1OABV1M2cLGYt8hyR1T4pZ4lTQ6anUldPlI4w5IWKnsC480iqt+
JBz1PWVyixYbW5nOp3A0pCmp0YBeffC2GLrZjkjIhLDth8eht2ogQAAJnhnB6e2IZjCpx4A93CJp
SjUQv1lmIeUvJEEzCAc52+PohJ+9w/TK4nG6UWnpnM3FvH7tCIjy0+TR2z08hlSbDSxOFjpqZolz
1Yc4TsuPx8Hg5aCGWB3Mho1HkJvvzZ2UzFOWVbt98l6SsgcSWLAF6Hcs1MqcHJnkEnqjSQvyN0EN
ryhUVQQr8fUtAwQCfIoBhfmwbZuajIDb5JP2w+4MRgFEEM3eukXF4VM5kWrRAi+9E9jFfqupGO3V
oyXqjkXYSjPC33YZhHigf5nTa7ycRe+kc88J3WGBXs95zj6fBLOw3VwhszcgUDqumz6ecGmGvdh1
nY2Agope8RLKxHCSs3vncfHRrBwWKzraq6j/1211o6B93yBZFv+mNHrUj3ewZ25fWEmUtCqQHRKo
M24l12cbz1/Zfc2GD1UkfJiK6sr1v8j7tAOO/tIIlf40XPdajs97l8K08um0RQk9IA8NLBsR5ik5
Sl9w0IOMXxQN420719qt4RrL8je7vEsWFEYEIKUvHUplJun963MrRrFUt1+OhLj/oL9JLnFnq4Ck
3XO5F1wl3m1DE0+/35CFZH+FxsbAV/YPxlK447IvpuMaX2x+OSsUCwQO9May3Ev9zcnxhqlyJr8B
S3tpXEZ+vAXGA0aXxhS9GvHajT+wUFuUztUkEflIj2CrMFg0La+WpahEPzrAQZagnVd2cYu2j128
IKAMvp/U0d9RrrA1xFe3KJLaHzZ5IMB1nDsOL+PV1VVNPzVTQYXCl2suWz3vDV/UfV6z262GlG5Y
nlaIuzjWI9pDotPJKOHTUCsLxQ+HaJl6XfG6mUXjdYathV1qcEx60C1izX2uC1MJKV7TE7vpuIn5
o0MKzKDe4HyW09QbKGju9B9cSZ6Eq9iMHm3x/RRDX1aXQJ5S2KVhhcnP5o2rT7E5e+Q8lhMggy1V
ZqQqMf7ITai5+MfSU9ssvCg0eJ9tMHnU1+LNyMxQyBzaOselIne+D/FAmXYkXtJz470xeC+FCQG2
q3IhVv4lzaYmBj/jWzfZkCBIfZiCcSTrDcNn46HL+Hw13Xm7lHiQZSVbUnWOSZjdBbvYosa5e5cG
L4QJM+GShHt/vQZOs30xYXoK43nMe6FMuG4ldtql07p5MrTlpCgs4WIMjLeaFcoAEmLTBGUP0v09
LzpgVAR7dNGHUezyKpm08NLq8KzU58AO5STt39p9drGAHBrIU3CU36BI4r90XQ7WR86cRuK86sHO
S/sxBCuTxvtIsz2D6Mt3t/w/eO1hujpbc8QDb/M15my3Layt0O9I8tn0jb6OMiA0MXcgJhOKf4T8
NqqIcca3LkTyMNsmRno2uLcY6lk1FPY+LmSvvoIEeg760n2FltXzL1i+fwYgjLygNziMh+p45c6J
pWvWfZOr+52sPX+tabGBhUvA8eTrk6zXTs0d4BnpuqpM8f9tqhX1ICnVI/eYcC/G2/ftH5tMsLOD
fKlrhpRrvRcIMGPC7yy0oIBqtU4f0asDM8GONQPLRyYUxe/dKdRTRApy/qqUNHIPnBaapggvd87d
RH8x9NKWXC79Jtbkhjk42TwtWcLc8iKkvREING6XlJs4jmDbJSdG1M99SB+4rScB+SiRtVIfJixw
k0asOkF4AynMjkLX9dWGzICPFI80dhyCB1ropi7rZ103dfywL3OM4RKdbcIdIdJ62qUgyTekdXfV
FNGG5FCRofkjLcuhcvhq8IGIg8TmVVD1AxcYyhRqL4c5bwsx/cl3PSxiV1shqpATQD1YBaCleDVc
rmahoHAajHfATUZ8mFVCvLTg4YQq20qFMxBLMPv4GUjsszg85bx5Jf1oAoq9iPaHDOUvf6CJahjR
6TVt6rD13Oq2KfgAiGsf0ONnTLoZ4qhxMvSjsd6NSDysX63O4nnnPVpcKLHYvfQtVhEDwVVBTe4Z
MftOCa09w5XkaIBx3SAUwEYuKBi9QF8H3bCoum7lQVYmjuuCF9Y7LZ0K1/RzyXS06hWtWeMtPJbl
qFif1SNS8COXuSgRmgAutev2vg+0CEDVm2amdqJipl3tjhZl0fmYSgyP1wy6L0oYoo57u9byoH2b
4COFxyP6rG6fOPCxIfs0Cd2VtL//IWsOSitFZeLBJoYeGR0Uw7jpy+5F2v0AnE5u0ox+9Em/L99h
wmr59rHUllUur/l/DdOYxT1E8qApejWBA/T15X88N4yn+Loc8PIzTiJ9mah3V4MqN1enE79sTYQP
EgEOORU5DVLEphlHS3GTaYLbkLZEeWeuj5V+5d/hqsKAvD4hmqYCtKc5St3QXti8+CY/UjnDjITm
T3tMvxuj9IR60kLbgovZFLqmj/BLkRjh6q+KMSExk/M32RDeWFgckNM99rG8mit44mvi1TuENjJp
V7VkiQ/QvGK1RaxGDwThs7o0mLGnUq8Gwe6EGf1AJ/9spzcoEe5xszpjL0KcFcBTKFBYE5FScKEV
gsJ7GRLqwSTPyn0atQakLbhZZXZ8kiiESZTijn9c/k9oqYpvsgd7qkaEaoPY8Iv12o9cY/7siLAW
kN1jrpAKbrFw8vW5CSDtzUmo3C8ACkMW6571VpEGde7EvVLUZQwT41TnU9k9VoHD8Xpl67a83/FU
bL6La/mIylldqenWWryOAJuzu8y3iWz0KKUaXxex7CzUAeMfr2+WQR+2VFiGytoJ8DYfX5VcKEpu
+p5eUk7kyPbHZjahkUdBNqIY9QMiEQOCe0KI5wgy1rtPRn52GF8b6WzfQ5lKCLOzLuiltNGSs5vf
VDO4Bg23Bw1DwMBI5KLTQ1iwJ10SmPiTnkDisv3oHeIOARbKnTgBKP/wEARKK4x6IqPaSsc25JvI
K+1NAvQKW+3h+b2Fn2DvvX9Oxt4dLI2mWMJIgl2f630IKvQl03Q1spefo03EJYPwlKz1emvs68w8
zfitk5ctVmM+bF53vjuIxo0lCp1fNeBL/Zi12lU3ysHbct1hkNMfSeuXAPjRYet+l50aNcyZ7Rv1
IN28qebUmMOlDJqDcBx/JfDKLNRO/PyNugi6c3ShWGMs+oqEiLNLO5dveGAswLOkaXcbLoxqkezK
Id992/RCdPkS71UpiZjuiY6Z+hBN0CACdDSJbMie9FbBpGeLgIPnby8u7hbvjbFjWrMsEWZrfxsO
SQ6nDrVmFAlDcMmmIBKOMUyOWcXX+wR5wW/Dsa1JSgsmWCo5tiVTJ42E5L2FLqeCdds0eBAzKWKv
rDAgw3D4ll0j70P7wwefEvQrg7CK0LVPusU+3dtuemdgqNEWDii7jRv9J3vNE2WrxFfVweG0yVhi
wrC6dGrDG0mVG9CGoPxdphH8YnP0ZpvHDZfYbeWbDailD/lY+AhDJDWpHN9vqw+YExytgi9iYf0p
MpVouHnfXWsjzP6+hueZszrizyilqUAW1EcArI/FryKsSHXUSitunWEBl0rt6Z2+JUv601j7Js5F
H9TszZUNCAWI5+XfAswqah1mrk9jhKwC86kijBb9EO7Z9c91DlMoXwUiDFdVm+uPqg+fphGNtjWg
dcbY+DWrKLDvmhtxOEERcYvZpYRifdu5Ygl26lzojJfq3MTWd36Tdvn/ux8fq0mF8UXKF+TbcwuU
qvf7aew5f02xkvP3iUp5e56dnieN3uwnNMbeNbvRQ/bhQwokvthKpDQx/UXsSGInXHztukZWDe2P
fkv4n4vvDLnPEji6+G/1irHJGaDDO7kRJpX0ou9tXkYAz9OWe9TScCcty2wCGRs6jAp/UatiX5qN
uPPcs8csr8m12xmM9plVmCmsYEKrvmZTW2G0hEXqyZJEKr/pn1GwDv8s107Ehd0MppFXR7Gk7+LX
y9Gbi/PvfAJA1yoJ5QiclwkJDTi7rIggbA+6RTtX4A11Bx3d/v3cggNHnxUEYc73p6AgKq8fgBUX
iXgkMZ2YrJ9Y9tXhRIjocWz0uatWGQWrsgKwWj7cfoEgDcTeyUiwVgjCz1CRz67TyAypeih5Fw1A
p2WTUmwWVjwrnBpBW5PgVJyQHdY8YeVusYwhiuDrrD9QSWCrmkHHzrNt4M+zQSFOyAuqIJBeiVi7
+HDaWj/BrfHZhibWOd+M2dEDagP2Gd8yHyrijdPhi6Mm+KJJzEGvYJEQnqbbsBuan/ePx4BkGqjh
Zi+7/Dlyvg6OZZo1tU0szV5t/Tcz+xt9kE7Ob9J/EY3mRfWT8zKSudcObSK5dq1oTbISM61WRqxA
o4vzCMN2C87QilFbd/o5QLepLKAhrVlUp4bY5IJ/mRw/txQxTbcPFO5JrFSj6OJzdv3q4QwgCZYh
KxW5lnzhGyO+XYkz/P3BBI7hrW8teV6PegU+fQ0Sfiyejz62T/d1JbP46kjB8h9CA6UNSjhQSy0i
/3CQjUQaebJVs3mTvCkCAf5qbaNdLAeGv+shVHyMfLZzyN6U2git6QSpbCJSODSLhgooajylfwHs
gArw0yAT3LvbOsEStYBq/WynAmADuGXPVnM/yuUILvyYeyDmqGN5YuYNVK+xbgC7ABTcj5327pbM
04QgT7IPl9FEIBfndKCeNW/xq73tMplzLwuEw+I8XHKBi2kZIFiuPzqr5zXV/jt4yLj4mHquNiw/
BoQfyDGLNy0g+AglDPgoov1TrQvP9dXV/cSACFTnKQi2wb4zglfc4QXsKCfTL7nWpkUjG33AG3P5
eG8P3YjpRNsY0BO6yn2BxAnGckB+fkqjbr+McaOLR+dhfNtP0eBd9IoAYANCSTYrCMCaNebY4EGP
9BmZlqjibulHgrfvdBFHN1zRKuL7Z4eSGkpYB752LVyzCNd24s92Y02fZCJ/mBYcdtenysAKhdcP
2I/5ki2riqCAKaPASqQGOSzomezqSd3JjF3V0P8PuIC64DiiRcvNLZRwYmDnSu+uIWHMpH8bO2TT
bZjVyiTLvzRGIT1IZgJL4ksmM6JxMY4Fb7q6fiJDDgZbY1iTjyFfHDqwgfA0gcxgXXyLcwd2JahS
OSS7o0aeTS6LQESBz08w89BiVlcmCkQs5ryBcvVpea49Oxa2n8GHEKDehj/kX8T44W6i2xrCwwR5
bkJAmPCubHWlLERYIVOFY4A5DLT++ITLothKscd3gQwWh+4jOLXMnErjytqMnNaBX7QMI6SmvctL
GpyNQpHK0jlnThRyjeQuxYHzqoCr+QS9I2nybAvSWpnO/RnfLNHx/BlQ39dPY8/Y2QRMew5/CF4S
vXD4cvK3WnsxkZOyspBKRPW/bCe/8wgfQwed/FGUIUqPmRp9EQBnN3lwP68+1/ZF1DH645QVNADt
fsrW2z5/TZz48hDdcMMHD86zDifD5+D/37joCXwAHmMFyhJ+kJmJRO2GQQ8pHeNEPovULep5Qqxy
qZ7k+1N+c8ubA0SR02RpPPmtkqDkdOdCur93ZTs4icFhjf3PaBo/D7bU4G1BTX5EoJqpeaNeCHh4
r5vq5iinIWoTHXOeyH05VaGYwc2BUpgI798SyGaMygzBfa+xq22eJ3sHz4jlR3+VaX56U+NgfjM0
KZPoPC9rXyRfYRi4RnxsWPaSfFpXwNjUQZPoOuL18E6Vl17wniNS4DJ5tqqwk6vaInfAsqoCltPz
Xyc+T+zMZDIunElnnfF5dVuQFfR1e7ytNU8xqskAglqPOaUbnKvYHSpvjDPCfhbmqWVntfobkgXG
McofkQeNCBHU29P0JlwCvY6CH5WGG/d7jP82/SqYcdx8LIbeBsKBOetPx10kNCYeu6mfrECw+0Mj
Pb+BJ7aWCqG7BtPtoSPKzCSCMcVhQIaeD5dJXEfrBzGrgnezXaTbH8iVyrFtGO8oRzkxtRt78ldK
y7JGxP1ahxIQB2UxGoI9ESi6qtym5wToddBL8V9+mCmYGblephPXF2GN25x2RlGlMh79iKZiP5tQ
5v33R3VvV4TZ/H7lIENhIP2dMOUGhiwN0JqUE0dKMZsscVwHURpBpMcIl6vPrRFjc3pckWLwWGOz
o9QzIA/dnbFoBSfUm/TTVaHRTmlXCeWlL35OSBpnbDlsEnfcwAZfYE4SyNDyIul/srZacRbuE40D
Xe7FnIgtq+NCCak5ugKsoGSfuZYIOcfkMo7VwgCIVIc9Kky1Jd4+PwZB0ZjHqu7494+XyaSpjJLO
d2quvskx2CgRioN/Povcar+3d3rSE+62cvodMXoAJIYq0ssEbHRuOMoxoewJLudLZWAEI0I9g5VM
Ra73PcKBr9ctmgRlGe15RaZ53uGhCL2tSDkXmEyJmRpEcg3+oDgTiA9c40NTBD2CDKn/nZ4s79LD
4DNnNgsYRghGjEwS1iOjtwqKTJtLt9LtrJZPCBtZerry1vQdk/cakmJELEVCSpZ8JAzcB6s/kuwu
pUZe6+Wxmxs6QVaBjbgvNcKP5Rot4vRLUZKEeCWDNMa0dtDl7zdMeDSJVry+bYCw6LCcXcnRlHIO
otTvirrQTpTRWlmmrOABiTRb2fjfIuO+Xq5aQeXj1ziV5gomtBNGrxhpXfesvY0XIkMaP4e4R9wb
KMsuJLlG3iDguHPSK+hIH6ZgQpCXITlMpXBLncFUEeOdRvNyzsGk2+otE3PwZdpKG1VYpE8f+zha
k6RGxLmbzVGYDfOJxzs5NSxLRRUUTVlJbVRa4fm5DNJNyc9O0v9q2V9LQ+IWIQBPPl1bdjnJ0/ty
Hmieayhz/PS3cmdDqyjQIIqMf3i7GqtJlRywh+qcMyQsmGQlOFHZ1DFYl8GHv5LqQL7NfH37ukxK
evfvSHHg+qxSIFRX1w1lz/uu+99rdAsxEIuaRP03Ni5RPc9IqT/5pu1xFj8C0+AyFcgtDUi3E8Em
vO4rXsoxBs307H0D+PmW8JGs8femD0HODR1tDwZFF7gFt9eSSiFMaclfm6qMQ+zY5/m5j741MbWa
zQpAVC6y8dwJwfzNmVFVvdrkHIlWtPMepYDmkbdDTuWRT++gLt2M506c3krCw+OYksd0stq/FC9t
rKdFKsl8rKkyITYmCFk6TxkJ6qIXC6EljXRwXBzNEE/tSicyTFLnmAntwjd1pRPk5Fd1V5ON422W
PWV7dKEvwP45nRRSzB8iwg1nWqNOrzAvDc1DeQAibBxBTejeM0UCIx2aJG1ULSKPPV7m7hWQ3KGf
sjBljw/GML7h83e95JNORCv4gMB39IVBOn/zxYSjdnNGNFM8OF/c7bfkPeL5MetpuDwXtv6J/x3+
OOsOuaRjSSVvQTDTT9CKYamCfSqJ4cvoZ5IpvrkNfUGRmbjH3dIPaU9VoHqT5MwDxMC4eBvs/4CT
vjI/qxzMl4ArZj7XUlcW25Z4IpSrmK+lF6JTBYbWqr409jBqd2fMk92ZToifOnVGB9PWdKLjQcIO
ju7Sz4lat/hvR8S97H47nlMcMEqgI2fgUiikKjSE3EwhclbVnKO4gtOQm9z99bsQQavVPi+qD9BT
vs4yP6+jEKnHtoS/mhTCcouW5INvESEZCC14SOJsh/223b7V4jIPdwoxqvR7PMulcfaI7bkqyfoo
tLFY9wJvBhzES59XNHqY4wufjvUMRbFJh30ypF6IIfNQpvcGYgLbbPad8xCIhzjV821x6WqDuA2E
jeKejn2wP+e8dHkx59wfvMk9TheIr63vwQGX+7zQn12sDNo9iIPnDA1VBsxn7nl4e5HuMRDChdf4
e+OHvTlBUa4pJ5HanbA+3h5eV3nnXNxXelTbr/oyaM0zpQ2E6Fh2/Nd9Fq98HjB6kjgfx76cSsmH
eEWZ79/bipGghhkMe77bHMhakDnukD98GgNPctO6kasWl/pKraUX0inQBcn1ZjYuSyeAYfqsakXS
+4KtSkWFei4E1JheOnMrRxYflbWQthZEJU01Bjd8BjqItg1zrI0yCMfgrUopi0PtBuJLQaHnEaEB
r1+0W5nXi3wumA0z3hQI6M/pI25Jl5/VwzPDWcmXttFNf/Ffwzogk2LiaCOXDLRsTKiChxtV6YYE
MCIiGoGVHZYGy18iCJ2+xnwbgRMtDdCsul6IV/BEGK8C1zHeXKAeTQlwuXNMQMeXgwvDyuTtZYR5
PbjWakapKFUKyrNlCafiNryszkkKHxWH71sAt7g2VrKoUuQrITbsN8Djv0QHeVuuYOVUxUykmqZN
FPyfCT+MNIqar1oUfNH3p11My97WIiotASAkfyZLEgJqZx0lAtF5gngmBSd0U0u4UxAcaWqryC73
qKwutCJJnKzHx+WE6iXYq/tm5iLZNBEs+XlyG5bDLkLxqHIPLcjOPZK4t1UpaKUrTenQpi9ekJn+
hkNV1hNxT4zsAKuBwXyCB/UGHbsw2YEu2g7b4YURbP++fQniBOjt6k7N/dX6TG9e2tMCeollq072
bjRTfS55rF0aXv1zdxasqoaqKhnmiEqdHafQpwyZ39Pjgu6FoDir3r4fp9BH0OvN0F54vQOfKZ02
QMUBgq5rBWjDIhDY/U0OSwD4KDJIg4WB+AjhgbspGj5vVWK4is4B5yHROfPyLoL6/FpUsB1KKS22
W3/LYtTqDnMfOFPuPT9M5MALuFlyrcGER72xVVNjGdnLZqaUxEnS5cifjvt18dS7esOKlGUUUhjV
y6yjb0nvJxPrNz0qa0jeGuqnjk+d7FJnyY+cFvqygkkRi8rwCBPRN/LheO5E3Txjc2eM98jgziyH
T6EafrZ6Ja2/ahVlriRx57VLerYFRsM0Wc/u9jhLklYEAsM4oM5ghnHyqP3F5eIeSvvsRhbiGfyh
fndVjPZqIaVqFrUxZYWShk7wMTATrrzB5jKhQ+uy2pbX0JPRd0U9Qwhjc/oJIkcB55pE2Xro3+FD
2mU6SOUppcyOv06etjinbDzf0pd9an4q42ivEmBVBJz/HcdQVQM08if9IylBetsdloLyqWeGzmUg
ailcxyV36QxjdCRbxZjPYkEtX0r0/VUTjVhw7HqsO2rV01moRGbkQCHAJau4gFFROcW3h4xKdd/O
9iRUYR6cvhzcrIrbGPeoEZgO8WLufwBCx/+oNhunoDTW0QELoaUGsQyIwLrGg3qrDx3yBK1rd69p
haFbcxl007x7SzSxxkypMwM5uXFNcAqba/2F33TRuvQU2eSDs0OXQXcFMnT6H0oQHB4Lu6ZOP4D1
IUdCe6LmE1B5qqYyIPXriw36TtFXb0NF9zoQkn9YfShJgkNjiv2V2dCEUgWs+LxNrvhqvqky6PIU
I3vrUiaudXkObeWqFNTAmDJCmN15sqLA73Xi3pcdRLhnBx5UAMdJfUUzJ992zadF/NogKIs1va82
mQcqD3UjtkDbyplopjG82wnl4lavcw0m+TZRT9ra7MkOc1brrbdpAMEex0vZbiNWCKjZzYymrzj+
68EuNMYR93Og1OnoGFub8UG44W50WS2JNWw92WE0arMKTQUMD4UG13r5eRTxb2SrWHDcIcqm+jVJ
HgXdNgZDYiTW/cPWpNbWz1U5i7iAiBuJBkT66kTLPhOldwEovooUeE286B7cKW/Cu8Di9VQNzOvl
1P36cb66BseaIL9qy7ue+j9OOjvhD2C8atPMcTk3YH7EfAKhMlMbTTZRS4q7aR10LnI3nAx5SoLE
UKzNFo5KMWYAJ20bPPIZyDby6zAMDGl5W/22vXr7nqoS/4KHzbd9ErlwKjAdd7daS4BY1CxLzvSr
xIsWk4E2/be7mP6b45LULXjdJBS4dcZmb8CsI1CXoy8auUbjG28YzcAto1Bqf5+6guGhMwT53e3k
FgjaG4vAyXPqm1V6WL8uTKlcSLVtRKVaGeXTJ6La4VTLH9GXAbOZwAAXxO4jqQcT1ccdwCJOYV08
raMcbq6+mtFlUh52N4mAEE5XACokwO4ALzUX5uRVxLd/aRwIi4Zn9jgWEny8vK6RAglQL7GzT6Pv
RLcuSHNN4yO/xmbmxg7UxtawYgJNuY6B+5K9fpFYcYGVj/y67ww5rICLAsY5mWQWZ5PAqDgVRTpE
apVApq3w2UVL9xBF16Y1GBKb7lLgW/pGUhoVljxz3xlqP+R5j6+19xI7JvJwNzWzw6nsPhgJ08CB
1QvZeW/wJEy4n145Zz/LF/WyPpDaBH8gpZeALfr/JTPbMxXeCwjwe3WUzJPnsBB6nTGbbrbRTc/6
IJW3R6swo1mqcTrRbTgw4PEmDil+nQRS2ZbftIfyi2qjOhuZxhrWnZxsLTQbnpfIyDAPvZZbgvsF
3RQg8P+wnKsXJKJY0l/ZqFKjurdfhxgVoC4MgPyUj5IdNOvpoZBuFEKfOE7YQiqohok+NL/Uo/oc
JG3hNDMi2tP9ye24r7fu6JIeletMSrfIGyO9WpDCkOjRi64ZQgt/+ElAhNKEJPpG3PYFjmoqHxG6
/wU13KoT64cnNKm7/j+xaPjQt+gSmpUghgLCDWhOMU4BsHqrWBbTeMPvKl3hm2zaeNMGv6+EwzSD
e5JEEkYK2Ee4re5gK+qIroxAgq1jbjz/RrLsKCBaaPJqhSzp0eEEfcMxvkrAASfi5LsiTHcZs7k4
AJ7Vr7kgW7toJ5kCrPi4JV0FXd7PalaT8heHU5ta0O2pAusneFgWWTOD1w7nQai+yya9RGA8HNDP
3umBCz202mDpd1xfWDlZTn0aYuLCzAL+lj3MGqajKgiGrdMcL+7TCU0c8e6u/1jAtuUt2n37Mz0U
VHuiyOlyYaGbdfWiGUKBnzwY6VG//SQGkqVSUj6BG8epYUtvbevyZOvHmfhYul/FXAPB2+1KsAZz
lRqC380gYs7SkVvIYBmYf2n47r5gXZZlcSXq2qGxNzwJGlYW5e41zCPMgDlDTGYbczFR/ofm4Bet
onQtj51jb92QkwIN+wpmFlQFk09DGdO664xlTwbwky3XslicypAArlN8Huwa0JmOqP+rhXaaw10s
Hxn9+WmyROw+pF6b8e0xwPEMh6lgjwCIlF4ElGfPYzs1OY1kseVVM5PXWux2bqWvuSMIhm0kXD17
ychPUjq7Iak8sS5+g+y+pHnGmIZYDJVkJbk1hP8+vY57kXCzuVmHm3mT9phigUlObaNHBvGNPAsw
sU5p+nDLTVosJj0GwgpqVVtCAYyx2EZE2y8+ueND+cjX4/luZQfzssKrTrbyGx7Br6+uirQ2Ehhe
aK3C6IxUaLR8yGNBuRNitGe/gyhtqDqDi/IuXXvL7ZxLyPBegVMNfVhWEEOCAc7454jpLeDT6gb7
H52OfTQx2vkIBnVaQ3xtCY81/P2rQlGp5Ui+o1mFxjhe38Rr/PoLUsVwveb0uK6eIVARnirvzezx
3K/BIK6U75KP7cObwTpFen0bbdz6JCZIEBhyx5oL1JoGh5MiPaOIuI6IKPvCGeyYcQGKZrfwTP7T
yYeQWUIPGvxAECRih0zKUZi78B7CwxGZyUlxNxbP/D6KBxsaR9HOzIs8Lv9UKf4rCsYFkJlxRDOl
7NQlRfqxBMoKBjo3BD+Xyigy1wpABIeG7lx+SDZxMgYpgP57PS3y+JU4SEhtQBSMzG08BqirMjpc
Ge5Q18kBMFv7vKJD3QoYYu5CtbaPKxxaSvz1/+0/3wpbeqt51Pch+2Ye3dxVgCCZmy1lReehZSfO
fXR95imEBGX5HNhYMKUEEwNa0qOLPbMjJ5HFOYOZ78VFXvj6QohqMSexhoG1QfwjgP/w70NoshR8
g8RZdV8dpmjUUDmR3q5oLqs04KHDHxWls5bqBTiL6Caob2+2Xhyx2dOg1VGhHg6X5JsbXXqyKLDk
zDpEzAnzRWIjnmA+agLa0qLxLaKh7XkpzzA/rnvx7v03LKQnUGpRHVXRpRB8xhZs6sSkSOqxF+g8
RucMeOWy8jck7tDKJdL7rzp6VEGFK69g332b+PUef+JQHjHlgkhggWKpGMZsTMqYDn7r8WdLE/1m
JQvDgbwrJIzz7X/W7nR745lI0f1QyqYuaqRmb//ragRuNQxPEkYw6+Xzjsmy+Gt3RkMoqywEKMx7
HKuiVz0A+3IZwTgE8JlLnfR6DYtp2BhRJjy+alnezFPrZsGp1DWgnxkX82OrRgRjBnj5cyNaMh1i
hk0cVzh2f7GEkZ9SfbE6ZkE8b8PyEjc4OO1NnzCV5+rwCbRoQAdsc29GUjDdDVXTrxDNTgi/DtkN
sU6vNnmJi4J8/4GzCdG/eELiDXzBUcGUH+Nmp4HNm3C1jTfI7WF5vqyTwPwaFu91eXmrIlCWTlSj
ISg1reefRpyAKFm4dF2yKGwtZYluaqI6ZrAldCXZVBfhElPv7lexNQTcGVUweRHOxQ45u4/Ly6Lu
0DgB66iRtpM6m0UWtO8CJGPrzwM1A3Sr1cgdphkzmeM5kWsxXZ18Gq0H7t/O88DHe09riiGxDu9D
TjS6QYebEgXlWRhyVgXL4oMOfRdeb+161WiAP2Hut8dAQwlSqAlExKLZ8xB5VdknDzMPZMMSNjsl
lpFC9hRKDot13D8WU9IvfXL/f8X8uNnpeNfLgIpuJc53Wr5LfarNiAABG1IWvEtv9u7/dDSbJPeS
JXaLq1kb086zHgyyUhGwA4j91GGDteMnAd981f+Z/e8YCdljcyFqWrwUkX+Iui1mIatBQ5HsrF0w
3C9EM6ImOC6ErpuMOPCW6t5BUNwLrNyo05TYIyXVm4PqYTWt1X4zsUFfF61FCHpoiL6lH6X22XHN
sXfufPlQdFaxyV7ASxZKyvoQqLLrNSECKZTwpA++lVdhbJD8VCwQYNAVV2UiDq2wBPbX4CE9ivRb
odeIRCpCjzE3jWWeuFxywXVRvXKbsLfUwTMLf29L8yEN5WbJUyqlg60RsazmBMj2lLq7iHZSWrxg
HsukinyALJBZonDh1EnCdPTLVZaI/aj0iya6PeF+zk0ADm/iNwy+ZxCCasdCuV/mE1nltsQgORiI
iz/ECmxGS6kxCi4j0JN+p3KeyG2Y2YTKEZDIgcVs/h7hozsfclSGimjFFrMAcYUOeCRRJlIMHiaS
svSIyTkF2kEgk/RIjDm12CvRgmuYjgSBEfHKhNwwAHu1k7m3FVdHyCzjsqJt2cCYbhIt9MFH2Yf7
EgVoeXQtTYPaul94VF517/Y2L1oUsL91NPEiHFjFSYlHqIMUvU3LcAusGxSQX9xNoXPMMBkJjhWh
HnTpzFunWfj/6i4wB57AuLsCq+Pgqla3ZjqV4ermZ+2AA8A1awoQaONGHeoLJZXlnt45a4FI9NkZ
gnjeELmdkgaMaF64W2QyoE7cYYZnXgRyqAjP2Xchel3dJWPXIsBobG9fVaRTQe28YDVbNsau+KbK
xneXBY6cT3D669D2k9UBaiumPVzHc3lYDGGOwUl8Ls/m2NZvd6E1OCJJRkfnEwGhE8a8hcTSFAv1
td3ezoF/6bD5UnT+5RyKIsYFFyjbKGK3wqFYnkFFuC7a/WtJtsUzb7Sp7aez0k64IaGAguBPnvlo
BK7wG+qQ2IZyjdRj4MLJ7ER2zIm4BrqkrXwM9emOR6zVlTDpIfMtDU5rgfpUQiVI0ydQrYHCIXQQ
+lhGKlIAWPCxtYMsUr6usNTFPEsXwGSNIWxisBItSLBBLoDX3hMQr1yEmQo8KtcoNNnAExsjpwp1
opFYzIRUkrUEeGW11ahm8osph75YiN20xobAchtPKpSQOjSpi2TL4OEnWZw9/dl9y7uBz6NDbqSF
M1Im/bKO9vEdI8vqiZlIXFJ+ERqyTcSdiUZ5dPqjCRLG4wKffjFOhEGFZRTfy343ckZ/Gb8f5Qq5
yqgXKNByueonSH+LwKaWsMS8bbF1h97gRx5Karr0XIX2u56yGcTYOQClLVWzOVpyEnRh9pXmQZzC
inv7vVpWrzNXfdcjjSk7ydVQM8YqPbG2t9wawQ16qGTbktVVfhTFwbGae8Vzapezo8CIBUJDGBK1
FxeyXIjsfTsN1g3Vil7U2TjKvp5XdkGJ04ojZ6n4uCuPdlAJp9Ceigk4hiS4RJhqc0NdO03gvru2
M8ccGrNT6kqydA72riO+pxI9kO/Qv6GiIpTGkg2do+gzkEmh7axEYLPhc/p9jJP/VEl4uHSCAwu3
9R01noKi2EBuZe5A4kNrOhBQv5P0g5/nbaqYJ0t4G84eUANy2WkUnjXCA0y6YFITNSX+INi2B1X7
wbaTG4W6ezLMw/CnOwkw5sOjh6433iBfQF5dyeCj2amkLob9wMbz0k33fJg1LnpRpsC5nnGBwXQV
RVYS/NIPKjH0PEHY/IJOGRHGjb2U/5ZbfY+C0yiFAm8TjkNn3cEWKlOvpStK6l7XnltwHugW16hB
OB2urMqhVRjlglxcx80y0ABCFuHTjQp7c6ySpG+8J0JJ+roYg15d8gRno4lOHwO9hm7PMpey8mXG
3hAI6TVVowbeR8o8cSS/8DWVcuYn7xALUGuwG/JGI5doCas48V1U/yrPS16GTYRO+aHjyMvMkp9C
sRUlRTQk1g3PccFQjTGwYTOeIcJaTx10ZsTqsAZqc0XqKAbCzVpHisofoYWx7XkUxfuTip+wa6gm
8/k1MT9DPLLNMLQv1y3u5pETMdxuHB95OJ7OEZKo7EytCnYkKfHPKEdLOxMSVq3LW6RMFFisfxPH
YCLLr5p7zHeapVBFxc9G5IWwgqycepTEvaQ2R3RG9hj+uKQFlrOJwbekwePRJTPVWOZewW38mXHY
oMbp8x50zH4udb/x2/jJqCQ88Kdq1cD0YNuhvU9vHfS113uvGi98+DVdwvoJdFpywkolhql5+ZZ2
Ub4gHv2aYW2akt0z06WTqT6LvjVu/zjBha0BdW+Nqf9NL1eR7onczyJ7mnQY2rNUpvMvPpsXEPjn
rNyfQ1GeGpZqp+F9JCvQQZLp4m9p+6Zef9ZOR9T5H+eVVbcEGxN+dHiTJhwXUXByD5J9YbgJdNgQ
VO8lHiVxwCP9er427KGScg0MAdQyQiVHRcdYC+T1CyoOzSCWITCaD6zkO8RwBJmcxl9NaT6hzo+7
MOuk6EoG3TEa+/wzjil/bc05Tx+ADuMd2YF+oa5MkaZImH7gMqPmikpVi4QHg2qteuSIdeirTyR3
se07CdSjpDQ6H+xequbfKFPiPRaW25xe7QtybfwkdkfYDsomwYD2ObgqkMxdJENIt3hOwZhNrbTB
Twa6rPQBFbNbS6afXgB5l/ZTY0W7RFdUikUbuAMMIfu8I33/wOxiiWJH5VAWYrZq/Q4oWv56pRqU
4D6hEFegmtz95C4ISahxkMMnSzH5EGVZUBpW6cTZciafEU3tL5phfTaBqkuhci4B2XbUdAYVwt3B
UkWfZ381GvQqhrDHXlzAzhxQ3SQPoSvsRywzSL6F3EaTEvcDGuGxB763A8SdJ9PJfvb/hun4k8CX
bODlvKk0znfP2zKqu6ZMyzgfyvr2m5vyjyxFj5DnuB3utQKafvoETXkH7xeNDlfgQl74Fhu/xnUZ
lsYGKRV78zt6ZOWsgp7Lr417j5yB8npxwN2WmhsT4/KcH/n70vKjkmfqAQmyZn+OC+V0RUhbo6+x
dqItnP40Naw3VlzgKm8H0iNGHOZwlPxK4eT0o6UM+TawbHh8YE6C66fie5Sj8fgGrvew6gHwHYSq
603lmvGe+5ITJ5on6WQgNIDAN1qmqP9uqWohukZdFze7XJOf19AJdzUNExGkyTDpyGC8efWaYETo
YaEPYAfyp/Gf3K+EZeEgvsiu5sV0YaFmfYqqbmOdY4SHjGJW3U6nXL4S5U2kPMo8huUHFDz/V99n
wS/MSL2+ierUxYwoLQzlX+4LVXMx0bTS2j8vnU4XN9sd8cDzp46tGZTgABVJlr6R+KKWTQjl1XKY
3g21PpfbSlYRNMjWIdOagSFq+W4feXxseYTQXV29bahetvF3yj1LRsUjwM5JUdP6cSh2K8UFTQJ/
VdXbsY8anpZBkRZOwh7uYa1zGBV5v/VHwUkCq6zGJV/nphryJYDpH6n8e9Q/5tojKq8ThsrMIavl
XILnEI/oKKIfpmZ/TGea+q6f8yMveGSpvD4GYtSN88cE6z2qGfyguGPlK9cpu3mCyNEP6EGOE1zn
DkKE8BGS86q0qY+Cy/r9mMl49UIPoaFIhl/t9GBH2rPAlChofAkKynT+Gy6Z2Cm7vD7pm9Di+Sw2
xYAIpVCr6PQUJ+ypeo40xNwzwAMRvQEgsuQZS7l1Vwoc0mWUAsVi6PhQ8K5kOYHrwp/DHxHZ3N4Z
t9LSpcv4W/cndAREIU8aFVLB57Ttf8eKbJ4mdGMncYUR3CmNwRkqA2Fi778+8ltgnZWXgoy1XmXe
SYsDr+IJRjfnEh3VNeg3t/uxyF70yC7XsJVwm8F2Z1XJzWbJd4YXpgHRk6JZJrxtUi9+igIAPnLn
TBsAnRZ0zZQd4XdGfGXW2MPNJwjxmDy04N1jWHmKMDfMghpzbAD3Y7TLiWBlDrPfjO/hG5bPyOde
aorws3tbYL4ObgNlZR6dtrQZPzQ6peUW406H6gukwj7BG6yvxO4Rjy2YBPiPPqZxxhbp8N61Ighp
HOJtaRHFFlrH79qYEqSwu5ayfYB1eQ6A70N00VWpBZlPhkdWpFvXOjUNfyKt6rZX3qplFdH2Qtg1
wFC1Gf1nTcgRTtBRB8sYkIkgtaPvW96NLK0NQcwF00mXE4FSjJFa4a5WbXo+hwYe1iDLforKGMTM
VYce1t+NzwxtO1ufAVJQyHBmX9oSxemS2A9/S90SIO6UWJw2W5pL+CYAq3Ugk7DPqQn+56w0tYtg
rdm1KtTlG4nbVU+FE1R2USblHqCrZ7vRql6oUD4RP0rCtF/OgZjaP+Ovo6EnUvb+C19y8DQddllJ
FJtCkl4XDtWiqurTDrvY3XYzIbqboovpBQVBDbysDdP3EOXOStKJWW60MhrU4FDQ3bBI6qZzip0h
c+bIBkAUWha4E1n5zwk6oo4OR56qLEvn0aku7lX/avpUKXaylxf3q40LC6Hmsj17kbPMVeYDR/TR
wa/nagxiT6BAlUvP/IjYmVRfhFTI9jcHKeJ9Mm/MI7XVBDS0rJrrleWdmxkDURTVlZbFKpi7wNS4
RaqonGOhNC1cEjqMBxLA67zSJ/36O6Qz/4fqMFoCHf+f8YJGGZuuo/wDHIbfSPqarDWGpiY21vbk
ql+tCehx9T+5kArM7MKbRL6gWy8ZG6NkaiJ757FJVx0QpAwseJmlhKKt/9bkBPMXyr7pSwpuYSkH
XUWWPKrTneaFkJburNEVeg0AGb6KHobbTSgFRmg3B8QTXheQouzpXscj5lWR0GToNYqqeyiUbKfN
9Ek5XN09dk9xPg6NdeIjXr7h5oc5TpqJhc/Z2FJQhwMxxbSo9f2pk8MPQW4DEPkXHarkAOEXl31W
OxgJAqHxbMLtNCGpcCtKV+kvfSU0oLeT19D9fmA3gyXnNzxOKWvGvPh/ztQnp9cYvSjHTe4hdFNz
Tf3W2Q3nRzRJ81l9aIVkraEVx8g3XVZiKZf3IzC9M48uePZ53pkbDB30/iPK1E9maeMZK1S9rArV
3zz3QdRIDzuk3YVWs79AWsP18XGmq6eedYn3PFypIOwPeEqqJZjv/uk1h4+ODweinyRrUgHTfCVW
7EsZN/hdfLxPnwIKtVrTzzCO9YPppl/x/wRuDjdCIHMFAE3UpJVor1LGYx4Ogp05JUGIavwtKwV4
TsL+kNaSnx2en+IqH6qPorqQ33KO9ZEtbWW8Mlo5AHvZ/zd99h/OCIfdIEnlakfltI+k0HgjhosS
JC0IYyQYfM9Dc0GsjdJKJ86B70TLbbGDHDwtzOpLVGyE2+b6kWNjdIrv0ddD+tYsiLk3rTTOvbo9
lm66j2E6ftiGwJmT8Bu7Txc+oYcfdSW+QlJtIt/Lw6qcOmtVTbRZAHpR9J1AhL72bRMlNN0qUj+O
Sz5OTKTIugYlLW05Dx2VezvGQfhce6MhqANWtMTuCFbilSA7FBHJY1iPRe/MIyh5whmkcF2DoAp1
i3/AOfB0CdII0bhYeV2VVQ2LFAIcddgPDnefRhYZ4qd+7+faHg/0tBQvm49j4cfHyy95D+dEqUBm
Gsx0WoybYp0yFGU3TWhi2GOEs6SDOO4nVA5HR3WXx2PrHHg6Stxt7W9/M6ePsCoS9safNK950+Rs
JxqCm4Q8JajCPcjcdkNNPZlDFBLwjlR8ypfsDFcpoF1ez0bGivYQEgiRp6Y0Q8iRvsOFEbB72IwT
CGrdBsdUwx6SUA2FhkZ9oMSCDh9hUwgbsw6qH5QEbLX/CpdwWudioB7I8Vgx9IVWyTkGRmAgx76m
duuWJn6yeZ57/NkEBQyoTjrP0FCItcn7wyNHHA3aZkXVyngYHLll1+Hy48SsD4IP4sOfsbPKGpcV
9LWTHBR0pn+v+EfA/QoYqvvVsC9eUuv/h2TCvSg6n+XRBWE6k8k/XV/yexLbFgAWobPAnsdxgKKK
Dz8/CG9Yp/pATqauNaFlQOWakvggMNqJ/laCzJE7P/XU/z+4wzQlX99Svvay384DH8V2W72sM7yx
L0bVCop+KmjJ/hzwq534rAGp21b1w1KQLnJYfosuqi4jHoJEtBbhp/mSghpgYAtO5bIpsv0Sns+s
QdwFoRvlq3/BL46hdInp2nka8/HgfurDhhAzJmJKNoBQ0CGPW8i1uwJnQIjgXRPvjgH4E/BlR9dL
9c1FVFosVxAUj+kcEoUeJUBwUBB6Qye3wM1FrFu28O0K10j1u7o4NF3JMF0SK6mZOjQtViI1UxlH
71YFJcyNY4ccCT+dJNALpgztT4Dtnk/xQ5WVjtUTIB1vnnxDena5NDUM0upVtHoT85MtTUu9Mip7
YDyzcw5DqfGCzohPfciFgcnlIBJyqmkkkjrdGSRUcemkit8kJOdjVx5XJITZdFPpsm5a3GAc6nt5
ER/SB/FXZAU2rOzdhOl/YlctJKyiuE8S9/T1OoUDJWTDYkHEJ6kLVulu6TnOHjdIzl/781a3u+Qv
N9rTVNeldmQdlvvHdwwxVH3Xl7OjsB4ed1GUv0Lnt2NRjX6Sct7g1OGV/GFIQpAvtfWBKLD/N4t9
f5AoKJ74KFdViYTlsPpzCbK0QhkhazfYBV4xilagDIYmLlecur8aJ6HFOhD6wG2Y0zzYvrz92hK3
2TFzUfUm0D+xdVIMo41B/5SqKJ9qIh7WQv8J9lOqbDVt5zab3UQiEoS+/eCKoEmGic3euoelVXZ6
C9WVxIN3mluRDsAENANAMp4Gs4UwZzPrVHIYgJzbOu2SIO3xilUtgZxgkMEw+kKtN5uNfFexEOSx
8tyLp8rdU8Rvaaj2sIq9HSy0WNmMvD6fSzTYAisU7YqCcAlX8gHIoWhFHhmHE7lTpJlP/tkKYQWz
Q9Y8++YqC8uHPmW/qu9RgRC1TtDL3r66R+U8zuWJnScWVt9A+SA2ujaGUKrdZj24+0yE4HJ+Dgk6
KcwSY8KPHGbHVdxqjE3yTTRoDm5WYlzPRtPkcgxOuh8WeYuwYa1f9JwTkDniXdZarkNrmBkHRIdl
jV+6R7mJOpSo+sBtNE6RWO8rKc1hDxbPLbAQ3rSoxCjxuvvUd+Y0aP1Y3mNpfuQizi0ocRyCelVR
p4uqBJxzDrOnhfeP0CfXQ9/jETYBs9guj4sOjNj3VFaAutXKB/nMGeHtSuXG8/aMTF0cSJBGVoG/
rWuNptu9j6TRR1dKWxDVtsdT3s2as/Kunw8WfnjAx6hBWQedG9Ve9x5d4cjTJIgLQA+wP3Vs1L/6
rwmBy0lF5XmGUlZTQadIdR/5UF3DWPocCGJXh6I/ScCyq7sNKMS2MXlqJbIPw5XOg5es8AlIRSXX
B77bkzyvmM+4Fika20fuYtRBkdMgjyrZsV3bUFYmsolEpEpbL0wGR/+e0iQ8T/JqW7Dim/lEyYNU
tikO5Ey4zRAGN9m8b1c2VDFcU+AczSMkISpxa3r7AXwjq83da2GbO7ROTrtfzL9D0tTQT3YPX4ey
N4HQcg4vLUAr4n7iWFsmkbaaGqF44jIiiGBxTmmJ6rqhG+kn6o+jgHA8HRxf/Rkq6K3kbM66eRKW
riwPK0qEibUUwj1AkwkKf4Whj67Qy+5nfJB2aSwXn4c9AiGVy99D/Rw2f/KErQLy8kMlsvu+RvyS
dDx0GCqV74fA+XZRMQC83hcBBCftcV52rlvC7f+RjwhmJmxq4x+AjTbV/vBp05rIGW9w0SULcqTv
WBbr+bAqP7mIZOVqO0RXCShvVAFwmuv1JMBDPzAU6PCg+NMCRsCzY+9y17Q1F1c3TNONc9cH9GnO
wbPYL3n2qo+2BVF81PsLHLUaISJkxz6WUUY9RRvdwLhwEUO+DRny8oS/6aSGghAzoQMJSG6uejIm
ETCZ/982RcWNWa/pBp8W+sAUklYg7k0aYiNRkEGE24ptVVl21D1ZDIlr4ineMOvuNyltOIO8gS4B
4R9eS8H5uSrJ+u7vYPuIXwtoiT0l0aEuoFlRqhHWrzBpER+NmfYZOFFCVL3B0i4WhBhX0Id1YEna
Re8lif4uAN3FGhQlNWXR6L7ljrV1HtmYg5j7suGWAodOJNzIMGEb23f4bPkBoPy30QdTQ2QFr5qo
BeGIpp3c3Ll7sbEhBl+pqnRZMWk9D0Mgk9hM9pMQJrrGQEFnpsi660Msifacf1pQFYiFuMgyfaN1
f5h90oQ5IS3iMW3hCYU4T3CU/bxc3++9keFlL6lrbM3tKZNWEqbdHJpWf2IP+ml7kUaP2ks137Ge
TZSAPuqB9h3ofHksSIsslZI3LR1IVajIyv2qH2DJpyE7cP45yd+OkkEqWuc3xCyTkk6WL72VXzzN
TccMAP+iuSXUx30jtiAXy/BwxiAHYNxbnwhpwWYm5Clq0aOdHvJBnEksbA81x29SIMLwAd4uZ8fy
sMglHpKh743k45Mygwq+iWeTln5GiTEyEy0rH41tXKQUJe4Hqj9Dcuqudvwkj5o/cYUDhpeFujJz
ekIrJEePmg4JLJd134huc8VnzfdqzVxKnICpmYN407P09dliOH+5Xd+KBufASYnGMKcxOKtWh/lg
82J9wvRy+8Xb/E53tjTSPrVqatoOa0DhD0B1SF+/J9VCwkAP5L0/aKsi0nxZJJSPVoxEsmPq1neD
QIIa4XNNDKGWS/G8HLUo4yfWjhqXGgHnXkQfxlD675H/QqR8f8HQ6bbCSxXED4uFYGD0LUHfL/RI
Gqb+r3RVI5topyaFJAPIdNk4LyULCPIOqWZ7V+tzBDWhJo4P07kXMMx07bVkWHJ8QNRiH66h9cny
RbI43rcNOsLVFx9MRTFUOrXsMRDf89usKd0t8ZJ6WF30Jb4Wj5HrlE7MNNzTLG/7iZ4XkH+0SKfB
+Ej9UsYYeB4FRGDfZ+04Xp5DgaamhmkjGZDJEg5nxd4Zu4Hc5q3EQTisFYFrCBv95WR+V5WX44ve
8rkCYq0KtyHOdZhlFuxybuqRbNG1RZkZzoFTrK0yYDK1oAabSJwGVorINF9j/gOOODtsvatr/Z/h
7+Kw7MvmwD/OxqkYghozitCOPabBBc/38MRZa51PiGVUGH7HSbIi3v3a2eLILyjCKOCyE2Sz7I8s
AFviWUx9QU1dKl6jZXap77uJw/3qHPtATdvbJd51C4jGmKrSscxXn7k/hdnyHVebHHTrdF3COi86
1vgf5KARVevaE7y4bIkhWJY7oPQkdBUIPXMD4U/+KFWXjhrrMPiB/1+DnOE05LvvZu8bxsDoyUKO
OpFq6Nfos1bMLy+tMIMXHYn8hC6DZgSfAuaT6zFG8k6Sye0+c2fVHYSiHhByrm0++ysX/d30QRwj
SUbL6P08eG+Q1eUNF0hW7jwElhSpDvi3RzVyqI5vnz9R+SNqbdMenCevraARBFTCLiHftro7tylw
ooiE/CCoPgD94ckqBZ3nef5D4ksUPyQLiTkUQORcHBFZZDqN7nxGBpccGPmgiGaecexzbvNpuOMA
tJd83XLH3hvsRwzNY/1+3P/obuH//rKGGUsGWeAJbXsy+4+MGNdWVH9AgDCCDzCbPqXSyAtEKmsx
Xz2j2Onx+2D3FQE7ptmjlxA8TJY9q4s1P5EdiZpslcWYy/neAQCdrXw9CM34TkbyQwgqAGKeA7V8
YRSch8IidO2kCgfRUCa4E1Yjg+KnCBp6qWe0nBJ9TnjQZcy5I1u9LjbnLyQ0I4TlDuquyhzbZ3uX
xKeg1ypuxrF6ZjL/pMWAax5OjQ594dhtp29jftakOrO2FLbOn5JKV1x2Ic4dAXBngzXsaBtxOSWK
nHE4GTEon6bIH/RYP9zT78tpkekNg3bzmnl8GXKvpxMw7ayzL7hil5/tB8lw9kEs3oXrCryn6F2u
UHTBoWxMLYMIiR6CposkUQkLuvc9qbCLeRCVQB37vKzy7wNLHEfCRyoNTuD2YxhEQi8Dba2UN0bW
4AQXeNzE1Ajiu1IxTxcaI1fNWembMWQub8REzggszOOvLKFpWbfRkAbzvQ6NaAeD3SYVGrUaec4V
deNVUTW9+fTVQvxa6sl5vp7KaNjykY8LCEH2VleER66tkRrtTEC1tIaYLRwz1xLMo9pMhHqEG+Zg
LU2u7IFsTtcGfCvyI2Gac1FMhWI/BgOlqdUM5I3Mwfi/qefoE5zVT25P8ortOcOZ68FUWtCC7LGJ
eDNBtSaHZI+LXN0BosWLT9zxJul5+8Oda333d686GR3sx6499/LzVCECOtQFFR5Gm7odQjd7DLrz
ET3lHuhpK/x4Y2TNOd2aGtAMydG33p3TgsuiS/QYsEcJypI2wrcBo6izm1kZDDixC+dDDogt4c+k
EbZ2bfAgKsOEUQTmfzskVMUFXNTh7qPvVmQ/rKhJh/oAhep2koVMVoiqsxrjUoE26CbicdjuR86B
uRcnhFWO6Y1Rtk5ow5YcnOgnSS+E+nMr3j1+MhFrIvfIgyU5udMwNWZTxnrWS2X4xTojfbBOaJYA
itDex4DB1Ds3Sw4rK4TRXr3BweXJFLQqyAVqay4NRZFDrP6bpLr0mcbFuX06/m5upuCahAan1s5N
1T01n7aZ3HrV12iCLuyDppuKS9Q8hxRbFxEAQqSjSi5gILOZHCyU1UvCp3rx35I6mTeUbCgpJdqT
Ydg3yuuP44bs2UrJoVt4/Y5yQBo2v3UoCAF8VYIUcxxguKqyMOWDi+Zie4gvsMHDcgTgs/zDjwe7
YNUt7ShVWZ9b6U/pwcWzo3T9sSUcsYXIDXDGh40EcziOPb8Mwax4AhTxvTGw0WVT+4XeWbT+Kea/
ewvehlJPREk9sGynpnpOxSjsB5dG8SE3uhXyY1EwGQj+iXERIV/oPVskdMNHNbDqzsxtZ9hTAMis
RnPcrkdtZjKK2di9pCrpx8OyOSk5oiHDSi11K9Slpb6Ih2EtuMcqgSt2l8fnXCa4KkzHQhABgrDE
Bk+I2ZhX4Ah+DwtRYXRJ4cPks1QeWeSSV2BBThxJVNw/aDFV5XwwvsIiS4MTgh2EsRzF/xGsYXN6
fPPXSfnVC6rrDr228qMtg+C1YLi8PCa/N01xDr1ZhUNFXID9bL4mh/BxZYpeFB085J493dpY4iCJ
qCHqA6CVrQsRQOZRl3ffnVBRmfrNzn4YgRmUQVCxWJgv2a4SRAbijzr78CGAXMiZYMtiMoOejNbY
ig0T2UUbiSMtebaGGEQnShqpcrHNq0lPf4t/+O3C9QB8ULoOnSvBNG+SbJ0rjCU5vrfCuBhq55nB
3ykytHtZIUCO9ZSa/TjN+bAQ5b8zgSnEaq3m5XtfD1HMqQpMh1zK1FvPXM4ca20afbN++7BJMuxr
/DsgD+YOSp3n5ubDhqmmg442pg11YxO+YVxLY75ffRNbaebMPGH3tgoAibsad+N6RktQkUeaBL4j
pEsokG/1623vJvyGV4x1Ef7HUwMNijLmzcVWkz2HIvQlab6gPTVm05lmm1bvpKrrqHZ2ooffP+Mk
FsNjMVGbiHllaNZQjPEtqB2sLNKwSUlpThFes4jSTNeOOmFehVfobV0tdoH/ILMx5xtaqrUwY7hD
icQwT5QNFnaEiHEP7Vpp1Taa+z+YTxB9PKSVsVq2Wd33SNCgcHSnJrAs4FbHWwxmHdo5gpM4ZYRX
Px6vQn8z4sj9liDs2E7/jVdkvIVgSkWj+usqZmlwDX9Ofs41CGqMy1s2szB+IqjPFQKTwVQNrLF9
UOTZgv2n+zSVoX+szCrUAxQ2L04CuMgalbvY1iE55ABjfKyKImzwkjLzTiJDaICWHm93vwbbj84C
fOXQcWxcSJCmSnwE3LeLxSWs41bVt035ZWuqsV49fMxDRUTRg/E8amvpC8ovx/nbOHLyrV8yB4eL
8DsG87KkOUkWxjxem7NoFRoMy8i8qVgjBllPORUTnv91xQCqg3MK8BrwMoHXFOkTmRBaTNCYM7l+
AHx3FT98qphQ7VYNLHdhGWGYnSgpE1zaP5YpbZ/0BXy92bNqBYKZ643XQc6SuOREN534POke4tl2
vmSDmfmdusMZpGCO3lKnDQMwxf9ymWh3Ia5F2o6zdiaY11USjTaVyNUTufueY4He++tsXbiPmCVY
Kw01vlBRSweivzz7P4b0DncZQEyzgUewjPpNI10ANL/4WlnWBUlPyk7ibqZNWyARVwBhaogYMyRa
BJxd8Y22KNrUQMqHaEj5dSvW7QgKGqEM6+w58EYd9lg6kvRadlcivp/NrxE0uGwAa7YaUDltZDfi
IXkWCNByJhJWgH5B2KvQMxzwFcePlWzTBSDELpYNaMm/QujUiQfzpM46Narp0DTAClBFWxMh0hip
Km7UxJccWmsAz6gJnXKgf+EWaOCGSoi75IQ5wml1Fc1XLgnGXYo96w4I2poFJBsTDOHQ0oW1QCKJ
9rb3y6+kRBufdTlHnGCwy9PcTSTptbQqD/15Od6YL18XkKZSetxQL/l7e9ThN8mZye+Td/LPIfqt
axPSNvAUlJU7uCRiWWtHb5kYhvZzou0JHOcDTrRnjFxe0I3gqohvFL9k2PSp8Cp7Jht7OK3iq6Pd
jJuNw2IBzJOzPbx5qXevvurcrmiw3xe82vFOhV3fMiuaSxtKBN2cA2+p8Er20FTXkmUbBwCWHhIN
LojmW8jf31hfTq/idRM3pJ6B4H8I4+WdK1/sFECuMpJgUq7mF39PKDYy6aci+FOzouVk+pdNQjdO
Amoqb/bzYQkVN+0UUApnhstP7CATbPRcY0g69tTRrBUCAAiWChKHD20Zbg0NS0feOUtNb3rMZaq9
YRYrSpxkaf4GVvS6QC0rmPUbjcMOtS0V6LZR1/BTPbvWx8P0iWetpw1+aPZ9oqi7xUEIHoe6f442
OuHkXcFvktCnFSPgDh6MZQonZBRbdp3o07xpuNldozk+8qCnJL6IlWdfVX6d6QRhv5YBw5ht1+Eo
fQyKsN2Aha4r/r5MPG5EdfIWZqr3V7hABuwkf1HqTbNU2/LFhYX0h/o+hg0+gvuuCEgk+JXrp0RU
rqLRRkHXI/eqnkiunVFbjq9ZRNOqrg+fbO6P8gHBj3Pjo4rQVMFcPcitaT4b7JQ2SeWKsHFbEhWp
r7uEh/iyHQqEy34FP5YHu8TUK5zC+NuDjtYdO812Qx8N0kW/izbacC9l8DnZYNoUyTP7x0tEGz5U
dzcznlIxlfcpxvalvNvyu8rifmwOL0uH6gTtptCaMcRjYooDFu5QDQ0a+ToH85gFHVuLaIpfxF1d
0tan7uXLSaiIWQpmuJE4t7yOClOZ7STYm8RfKYVfXicFjAsqanlu6uGmr0mXf3e6dml/h+YHQJGS
KEoinXVfxKSJhTekFWv55sGQHZR0+gVZE5Hrp/CnxVO3YZvqTBHVcON2GlAhbWA5vETjYdsgRxiN
9xnfXPy0Ek5MuqZwbvElRvDbmyGTxpaIAwtLBZGDVHhUB5UNbCj+jH/76+pLFt1j1nNU5KXGJi8D
+8bGn/Qr+NduSzvbZSTfPCp7LjalYbfmlMgj7Rj7YTqlDr0gOrNY7qHf3TyiIlcLJakaJIkiGbop
rwxGpVh8hx3YuSBYo1hapT9lNmab2+SQNxcfc/3V+G/38AAVAo94irYweMobNID30syEwyqiN3s+
VFjtHu2+DT+TatnPTRk+LfZ2n/DYsgZ19JWzGGE4WhrGNoIs3ZGawWVpeUkbLhqH3lPVNVsWZ8nb
0IUMq8Ne4pxL63J1JqHCFpbG3KsdknU8vfZcY5T3MQD3Pzf2e93a/CjssXYfst7o0Syuaud7o+9h
B9wtzIIz9eQikleMNPsFuaps7plJ1wlCDhOZFSCsF/h0vV/yo2tfgMPoGB81VkGXkFBBV5CRHCXL
MkDr1kn7Sxd8mDGH/M3yfHoO4RzeoARtDxRy2/cCxOvXG16M6ztZs9KdfmniIyiAGvQ9B3MzSfs8
WMCnuf54x/EXwHFJcE4L4IpPjQg+3KXjVCa6r+EybBwPlo6x8HD+Zpotg2I0WgGEL0aK/lFtAzab
oGd1UvgI1h5daNqSyBwuN57LUxTIVJZaeXtbhfzmcbtR5Vq5QB/oEQLpEdkxin7y8m1C+48iiYc5
ZOa2PTo9/4O59CShw3hiHA6XHA4X0+LoIc5yL1LLVbJ0Dxm8JE/FvG+2OsLS2PAdh/ygexVDgDU4
OqdmW2nulenGW1/fKXrDpa4ujj7RiLcm+bPHnUr23KH/tborJrr3+C+80YfoPEqX/b7OJf+4MZcv
QhmOyn/2pZiFpaPtm57gii/kYFqC8TbUZVbqfEKuUj+sv32Jjl9BZ7sq3m6NvfJL16VY7YFo9T5q
z0z0tcGdoKwFMQznDHs8Uak5xA4Gx1+rMn31++z2HxwWDoRNru9NsKarhH4JaCnR21VPMtW/WTwX
oV9PEUIGhXR2ZM6JJIwcoF4SC02ddqAQhjB5IjxB+rK+0OJnuMf6zSibRpyrr5dfKzMeQhYHRE3B
S+CxKe39T/jbzc+Jx80AoBZw85etmmF9vHaKygR+6ag0NAIfzCoeUCtL7bg5u4vPVWoegKbTF7QN
/kjVG/CeneL7afihZ5jzf4QnLPhZKWSoqi4nNCZw3XHyhaYuDi21w2NdctT0Q2leUDkj8A0u4AEJ
ax9UF1Du+c1v9cQqhNZHrKLNhU7jI9Pz9qXgd+xOG9UJ2Ocjv7VhLiLgMpOYj6pOUrfAOZd6orqe
YD8TZtNb5J+SIu42P60QbR1bXZ06otgglhYXWIH5kN82e90FILkTf9dOunLQs1LFXAMrlezYwepq
H5zjt6uX6It7FEV8Wlz+jVYXPxSkvG8+QamCdCzne9yFg3ZZFXD9G9Jq8wf8eAILbVW9W4MsdAm6
BbnMXYmnGWVGQEGBwkAilcWYbt6M4q9dmgwW5ihKRFOoNgBO1kXNp8e4jqcjRjVVtyvg4TWPID0A
ygYZVBNAGHEE5NLEt85FdYtV/iyRvRBYRq8/q/jEDz6o75AAkhr1rLJIpxhPvhEr60O4UjXGgVlt
bcN09g7Sk5NelEW4FI1xYft0JgsUn8HBQRoD890JAXrVis+jmEenir6xK1td0KJiK10skE+SD2eq
V0kY88k5qOEwIyqe6z6KbYXl8wxkHpqyTrjPQ680iTJh5RfPRVK9O4Ryl76ohKAwESb4Jx5+pheq
BGU7nsePCaWQhH8OdbG8ugOBohBtNlXwZPK2i00whjRIy9e4cmNkWUaN5iiK6QGCDlVZ0dKEw4sA
1RYu7wm0GtFidORutQvDjYcE2IJA/rvQsXPqYuaixg9a8L2QGSXL0KMuPdat0xvPTrtZLxFjbEvg
c9WhJMcUWhi2pXqDejNadf4C5EuObpKMCal4EGmYD9L/721jaBWbwnhiZ4NwT7Nxni0mMWgRpZ2T
ggY0bZazlZJ3NHqntEQQahzdZtWjYdEv8ZADN9GYY8e375cxwAx3Egm+be8hAlB+U0UmL6ym4iFe
eS2wDwwBHhiWjCAlKtq7e/7yVtOv/mixG97zH8gpvvr3kNMkLSdTwdinMj2ZjJlwmNq/mYOLDAAx
2YeUqDD3cNjXtQXVNI1+JWYFlCmH77qZuAnoNhhwsSjRjNhV0rYseRC+5cCQQF+2Zllp7cu6VExN
N2p/4s8hHu314ZhvN+epZfhlw6LS/kCW+evk0Pv6ERkWPHpTXry9/jy+I3o5/sVL8wevD548xm1X
Te8Szjxi6pjB1wdUfHJQIH/w8Blxh4rUQZ7zLJYPBIQ1DfjJj+atj5eEluSw5PihMwcsgYYpEuDp
Ty1++7FWZRD2jD0YPAjDr/folpymPN7GYFCv6EHghZy5mwYrKrKy+/g+OrzKSMYTaWGV09qWVtyP
igtgsrOGDrsX+p8qhCWcStI7fiwGVdVGizgkfzs0dVZrBFetkD2magHfP8zSaDBthvLr80XYETed
Hdjx9cVk9nCcTcJWgzwbTm5d505aBBd2ERerDGc7ge1z6HnZ1Lf61CUtIV9KhnjUTLW2tyJ0JjnV
cUxR+oq6J9VTyI+075v5tMZkkhrPrH7pdlNWPJZuRGU6Y62mW3s9k8JH10YyRAe+m39lE4w6T2uf
mnTJplNu41QWYV4v6ExSRdnMyROggvzVGrsb9YO3e/SugTtU2vu7TSljyn38SUPPptIKllRyWX7z
PxZoHVD1xCZQ7QCnND+aM3SvmvTnzwNu5oJGJLlwLU8c8786Jldos2vUfXnCEP8SbO7yiiQ5O5us
P9VmqYhp94NoxIvptzAWnkTJmhgmH5/T077TcZ1lSniOXidWGzZ8AgVusvquw1JciAA9NnBXvX/4
NhvHqwz80b7q+QOhp0evoKfsLEUdvjioAa5tD6Q2maGoNJIdbapnpJ288qqt7yqWOfBgwytEwX91
wjIfY931GiVxReyrVZD626HMFAHhXWIAW5LtzbMf5+LbHVmQXPy6F+efMEGPF28Pkhr3apWKPSHg
pUrF/WIimhR5tZHyzP5IPLD0SSIiM+018zNWElY3bNbbmRiuxrXH2YwTc7Kl71DmpnzCayKD1nV1
dn9a7hhM/LF1sGOe8rSsYj974hEJGSRsiezNjMvk1PKBPkXmqpmw3qNMttodJvAarW+XcMz8MZZ0
wdjFh/Uo9/83+iMaW0z9HUqwTR9H2AuAvqoZwPsrsEgFAjLhY+35yM6TvqFBDDRaZFaMEtFlLz2w
ZVxYHAia/tIH3yitCTdm87xtLQuiMM0FjU+NEQGVgAmRmwJWu+2f0wbTFjP2q+GVx3QWQIKE1am+
Iy3whsD6Z+TjEhbVxqcz4yt8E4RJ/C1BxYPqdnvcrqatgdczpraUprvvSNEaL9Kp6FYUMzZPImTO
ifLYiDi9btMpqvMT3zsw56atIpDdIbtFhgfJ4ptLcI83M1GFHLiRso9IcAXJ9x7olxpkHsxKGQU/
CcCy1I1PSP4EQjl7+YEsk9Rg3q4T8OTWpWyP4RC9fA5ww2eCHgbKes2d1H18l/u9S4Nc7qD9jcVP
wF/iFCSZb9cvdISoLO40AznlDEXcVopX8G3wBemw3VLBwvO9AferWJJSu6Jfl4WJLYVNX3ZaflKy
7e5WuP6zhWSyy9jiZv26h0v6mWQVFHNfavgU9WqQZqapMUCIJwomoHXWtxXxL71uXc/IMFmeUxvL
YgAUjDVP4Sq+TvKSXTol6oH80s0Rb/FVzZ5Knu1QJZBrvXNZR1+FEeRYsyGXia+FQ6zRWBROw2N8
zAC3N5o1GvssQF6z32bCMbxXYaw3VjO+kc9H4deryrQaJ0WAnwqOphVWD4h5FvjjQEvmyh7D1e/6
0Q76e+BZjF6dxo4XfO1RfxsoT/KOYjbTpE7Gv5D8ESd8cojoJevNOQYftZcaYI1g9cW8HpuWMd1h
9SQxo3zwiVYVQhRcLzUDV4IdG90P27k6rNigtlCsPLM//SwDg13dfq2XGB5NHbJE3tElgLHccGPc
BjmZCdcEUVCgz5wZMZrN7fsxVvwz+I02+KnS2m49Yyy9DpX8kg/XZmh+OcGWchtnf10TBufxcTnO
B0inB+Yv1SkzhhmhDQaDzLZgHpPlp3rnmZ27rj3SKetPKYk/qFHqI1EP4kGNbUUeLmplV/8XEUbw
rJjZYmknVmm+pt/Rgg6gx+9SvSKd3AwOY6/wLosVBOoa4R8HAPRGgS5N15OsL15v5kZvnV/TYJuq
n8bIpPWiQKOZ0Fg9sujg4dOYrnZvqo4/UiL8GjFwBbQhPkMjOrVtbDGA03Ep4fWDfBqjQ54pMY55
zdIoF2DQQlw5khyW3OnOJF8Yg4wyCLTayXYSBsqSuWXofpauqxOqZBm/BS7NwrlTCnd1gS4wcAMB
KQEaBBGXCupU9wpRUrYhNZDgqMPLHXWp6xxlnCaO19tsX5yLzDxt3S2NVswSTrDsMwYRwVUATPGq
24tttWKySFqRkIzGl9Adp4NUjlogswpQyOVYVnyC+iGW2zwLNCgYNQltT4hVc/c2H/anEVuk8ODA
tguAXhh6pJmRSB++sSwyQFDmT2itOxcIMzFA66tbSQFwJXb2ajnD7ALpMB9wVDEnzk50PMrWQSGJ
nnPAaHBJj9LF5K5scNNgY4lb/9GktBt9c+CPE2ii9wanWMt5+U1RZHDG5lhNaf54uRcwyamNC5ej
dcaxIHI6Y97NksuYCZw20sPDald70lyEij4xZd0lOYNL0wEGoDFk6gtybZxXOlP2qv6OP+M0eg/W
jlKQO0v40+srABpphmHp8sGKroL6i/R8n8Vol/et66sb+DgMDke+omApOlJCnID6BQi82zhCP346
ElyZrjSa8uX73Afp6Ar6GLXvzWiMHbTu130/ZMVLomtyfUrhkM0CbgN4h+BCPhU7wsJhpwzhWafp
Lm/puZBmHhxD/choqF0b4z3B0dZ2qP/nbs6eNdaFPA9/VO09AQjC44sN/gAfNhl8VNyjAUMfUF/N
IHO1fHVwTqAfBobQ8PNH/Jq2ORn4xMa9yorUzime5/WZUEwMeq8wyoYwCIfOF58xPmivB6GSnlFk
18SXdBfSJGL6cWKdhuFSMoFB2IupBPoyCCoMWEGdHXTf9/OYVhqIE1eHxNC+fWer+ETtJq+5VNYY
/1XqUhGRDikThhNwquJSPltq/zNwDmWmnJx7lnEd1CotlSLPMhmQvEOHz7Dz80RQIBXTwJjhJ8QH
zfisJACiMjDYRlgc1Fm7MYM56UuHm9cEn98abzOAOyQN/cWebqoahsqEelMG42qNjh0Nk0skgbfb
SkYtxpGqBUIxqpg3+n7Uej7AEaC0pQsVE+UDAtm7szbMdVO+ZJNib5QNklsR2F63JXNgDXwuqE4t
a854OTJ9bWEWoAxkEInubJDYtsyE0UYiz47YNJF7QIx6Lch+n39YmKGeoEbqN4YyGz92QOiDSDP5
0l00ETN7+R+oW6Qe7rT+JBkNIzAPH6d8uFgHgw6rHKk5kMvLPbDsABsD8bXaYqbIJH8CA7Cm8Lss
Ui26J+KbHCuOnv4P9mThyx3850cdPTUzbSy8OFmIJxWK5AqCsUU1XSZ/Fkra4+Cxx8Rkiurr0fhB
PWoG6S3fl5fVNkdd+HLYB3ekPdanLlQYzu+pVGH8Q11vf74u99zrjn9HA1Z0TMdWRNR+kvrgDmrT
SR+67WcRvRqSmoTN1nqNzbAvi4Fd+bEPSiOxsKSgZ89rwO3QxIiBD/et4ylYUdss114dd4xPmP4l
19jZv0J+9nIRAFdvzaIXUE/PYjdu9N3FqxdbLN8A+8AJ0bGJfxO+7VdFTTN9mkcFP2TZEmpj3L+e
jAiAtW5a5n7GwsRVHBEuzVKuUt2p87pzp6js0kAD/t4J1TSdFqWkmSr5e6QNGZVuAsJU2+7Xpidz
/L3tzEZTdUKdrYy6vA8lHnOL8Wko9HT+P0IXiHO+Ca/FBo4bgJzjiCgnrGhNzxBmUSnNF/Fu1PkZ
vDjWl1tIbBWzMGgERu/Aui1rib5I9cs2ZyzOaxD5d4fVu3vVN/kD3SE2nP+6sa8wHLwoMtg7bL2D
yMQXHK8iKUbF233JJD5Lyl/sqdQSvSezk/P9ps9zW8j5UKdMSIb0S8feOnYvUYfGmo8lK6+FtbMt
s9M1+ceIZ2lgoJ6ZcfB3iqIhfBD5SX7Jnr5rsGrxswjUnLVgoKEOH4OLxd4hFPNVkkw5ZFk1m0Qy
/TGeNGHL4FbUF8W8sqBGaYIfyKH5CN4/9jbpfx8H1KdqHI068j5lweg39mqEK8DH/OcqaQbJ4DUY
ut23OwhxxLB4IEfKia/VQaRrPdfhFP2/25R1nUnhwvzqkN6ob64tOi5dKasNuGjs1/Y6K0sIQzeC
xJMCve7dTOIt1yqUKNPJlpvH+FqFIJGiIZuMovDML9Rz5KQFtFp61RgLJVWJgXM1v505wOIRaFI8
LmSi38fyzxBQRnZCAsv/A2xTmEbd0ueA6Xpa5S5xYTqzo4I97AjF4vvy5+wfBlS3PvQMvwVfGnvm
y+S24C6etktaEVB4BQNe1ry92iC3r8cVppqIBH6UHxbRdHGP2/fnmONsri31Spx6dKcPKnaqgJEA
VQ3gIgMASQru2ZofC6fG7M2paITVFblD/Ojejy3mYselxJMQLWqwkC2fOhkPLGtj6Tv1tAqnTPVT
pvvzyih970d6Aw82DJl9av+gwip6lyA1oTQPDg0rs1OM1wQtx6qIoqiNu71TBonMkcfTnWmwXQ5A
8XnBD20e+QZTFy3vy7gxWKmF2iA0h3HNrKKOi31c0f0Y/ADoeM+0sR/u0ceeyWnRd3PyyZMMLLvG
i5mbsh9rmPsub54MEAr9KPtPeSoDcZ4n5roLuTGX9Uy/hz/Ycm86e/I8MTrDlqtfy5l5P0nxiCIK
9+7NfGtk4pTVRukvV2+XXNu3vv+pKuwbJ+eoIr8Apy1v1zTfyZL4HMyqUkSzNQzXDS+p0kfYHIs1
os0OSEQfptYL3XWeAzxdwB5kqnG+i+AuUMU2dzrFnBs5dA0iJc5hIVYWN6BPPUQCXHgMolwkGjEo
FKgkZW+8XRu2G3ADQZzEJMSvaqA6l2zdWQbBwsCPC6eegBAt1ewL0nNJ5y1AzDKRgsVEM3FLYbki
Ovggdgqb2iq8q1wkE7DEDj32ChLGMht/8je0kQitun8UQubKR3W2Gon1sYcIH283fvYLLMwT0FPR
5xWGbPeQY3PW4wT86KalRfw6k34QylOVNGG/eKRYVA/Zyyk7VteZtkxXW+9INkJAS/320DJmBe4i
GEFL06tjUY7jC69Kzne5Zp6TsExmkoMJzRoOAMdfPbsBnJzNB+9mGFwA8+Px/vBoS4LMexMayG9x
w92RLgJgvB3jNNgce8XPk6IwuevzJ3szvj2JSSltNxCNRnVtPPWb/c92SkNK+2/AgwZIfa4Hvcx+
ozL0rw+wDpkIBiaB5QRISDxwy1aHEWqWyYfY5zcWZVx84BLwFk34FgwYwvqWUPKHbAdT9OqLLSJj
F0H6fiRCpAG033fx2okz0ylyPaFN+iLu9o8BoqDSlyTwAG/udiSTFJPYLrct5yAKZP+vRXj5GEhM
lGSUdvfx8T4tRxbm8tL/kPNKW8zJF+fWENxRPONVyRIK2Lw6ahZaEam8wBj4FPACWTLwBh5Ti084
+qmqsNDaHQJXlt35IC4NKsQE5M805xiPMFt0dhPTrielMoR7Tsy2JZmeizre8P/0XqsXxRIgijYh
0bwUa/GiKWcotKMjdLM3tTOk5M9rNsNWUq+vtSv/dFIpq3PZMBwvWbFvB9KFmA6gireA2Z9l0ga3
+fg2JCS34kg/F2YEEE3k9x8ZgWzJM4Zwcn1jmOj1mmO+k9lHl3aIP/N6EIuZLxq7PEcUUq0oI6zs
qy7kd/szHybinObOiyeG2so2MlbO9FM972fmgsPre8KyxmmMcjgh7vty0W0kwC5evkDc73tByhA+
/07TjiE4yfcWdGL6Nl3wQPAcXsG1WbTCrGyIQw2q58RdKdMkltCANWHyIjQ2pUlPyC8QcN9UdLPb
byHbIKi3GnUT2GgkZLfpfPO3qKMgXA1uDicAo9REsg5c3SON9zS9YbXmGBkM1AyvegfJZpctFT0R
zouvOpzNpiPmlCVRopYIBZh2cePGPatkOK1VEQ2qYg/qp8svt2ZCEOd5w8V1OrBawCihHCXeml64
xbwm03EhlOKYgxkQ3c7UD5l6d47Ky+SpiqvixiP1WNBGT8HmkVsk9+Z4tN6YEfuCqJ4IrpEFPztG
0rxREne8f79pOm3iXFZ7F9phUUJfo2cpbmXwdE5dhwPYjy9T9MYfoV8moa5akBzMmEUcVU//fIka
twtajR24eUJ4WZrcPGm8xvAwYyotgvwpNN3YFmOUCYaHEe8fwUvV3r9ywY7s5La2wdAXZtXXdYtS
SFVfdo9CnaSRui7+koeM2woTvm4TrZOpZ53JSymwvpOTZTzzg4M9XcXKi60PI8QK9D5Fa/LKlTCA
zMd+hyTn6eXKjhfcMWYCnG9nPkcIZp+6SsTMAPSCN6ujGb3rGy1dZzMy8o9tHDbTqxSdiC7ZJwX8
sDfIhxSDHwtugrZy6vCkDv+LEPq/A9/hvnqFSx6yJ6TKKSHCB2NHjAb+MZqQVrOd7kWOOm7SP8T3
E99Ffa9H6eKps4nv/r/Y/G8gT3JTjpwun/n8zt+MRhqSlscmwMtzF7MSyzA4QwuLP5tQeg8N0wfK
jz/VzDTWIGMRe4vp4NMdDr6jamRomgMSfuub2odSV3CAIPobGI9FIHxbQtW+5ZaaBFIZaw1rIuBU
5vRulOOA4bmRoBOx1/N3a94UAuiCgfbkuKLiGa+JQKUiDHSEUgGKbkUk+cJNC+JuJ6ASF4rFSQGY
zAHmOav5Wkuq/xBzyUYNWGyp7JCdiTUsAL/XA9hnos8oEwTgRm8SC4/0aKIg6wMM9naPAGqblaKg
1pfQMWS93DMIZWVZaJe80KliSUcVnePdtu3LB43WLfk/j2ZiZ8Yabq92s28svGXBlnmOZXV3YdsJ
SC1Se89mKNAGoBHVnfJameWzLWSlyGuhGBYsUQq0ca3OHL/OryiWheJlb3vkLsXr0PxRHGO7Uzv/
XARZbe5x2/KDXgSUuCNGlybbAYQR1VjAU6AhWa8sD/U8/9cbcR60C+kToFMSbXVwUgypOXyzvvmj
v4wHc332E6qOTBIY0iHXcFcKjOYAZY3bSfoQLcs2si94eU3dQffOk7Hze4HU3vKOm19JaMN6IuDu
3xLXH+t8BdwONAAkWvNPBVdnhPV8hgYfPF4uEcVCzK7eq7UQ9uU02pEHyWUko6esPq9SJTllP/FH
HKGh0FdSxqwRthVEkvJbpSKenLUKXLSPRjBkD9tJ8j/RMDIWotjRGuOpzBULyclGGGTermNcYZUX
tAOVEsvbBwZQfMx4hBqjyEl/+vK43DQu3wlOThe7f3w1Qx6woj1PcA9MURERGOms5dXlA56EYVXg
oZ9Lcses9GM+kcgDcccWFyrtV9V/4D4C5Al/m5nMUqqdx6DzTubrlU+D05djeBSu2ApGTf9zjg4G
Q5Dka0JYOfPsrpuWBlEip4pNOJyOa8xS3Usw7E19brLZBf9DadNPahdKmDibHvSCCYEVVtn2t8We
mIGylEfgyVJqPKzMJ9cnlphUa+znuxiKNBdAtj1b1AlOFk9YC/rwMnpd30QS7q+oQqPUpK0VF7aG
dHKf54DgLsLSCVZw8GOgMJz/aRxQFaR5Wbqzirn7aBgI2FfESEhfQ8f/qXkVFk/kEabK4cw9ocKL
W9gBwxIbZDs10MNYsEesjD1GV9JyRHn/kZRFZPsp4Z0fMSlfw9hG3DhJdMIRXUZO89i1pmTExlwG
ZgtjzrgrrmUT5lLO1zAb2sDASKfZR/EKoF3f7dYzEGzoWR1ePnsZix6zUHz/Gfc/BYUq8argjmVO
lRHmyoPi6qJYvD419pnKJ0TQ13aID+zCszJx7ebLX559Lht5KYQSI+re9bv6V3sv93Y0BcGPvJcX
gk2H+RYmeNsS13OweVQ/xSxaWDXY+hnBpAkEEedZkaf7rhIBqvs/fyIX3FRbIDPySJtlUEXSOFj/
thjCAAKyGKsokf89Je/ykvA3PpQsgKOSqRfwxEKE7LgDsDcr32Wr341o6V+2mKBEemkRcQk07K4b
6cbBLZ4hcpa0JMI6Pgj0pAlL223R7oslIiLuX9dU9eY7GBpZAzMr9BCBuLC9E/PEwRBkgH+RE64Z
aiwocGUQlLvDhugx8rBG1PFYGMox1Tc8vWe/2mUo4f4JBdfCZvgu6OHPwoAJ7re8s7Vrjauejgv+
DnB7hjWCD9ZrI8QOJdFFne/KC97AcsyMvGDHWwQGObIvCm4mXzStk19Q1qLLESdu36Y7cZsiC2Ex
/vnfruEB9I+LtNYsCbZUf4baEJLQlUG+ZRNDF135JRNhge3QNFMAjvJhQCBE0jRiaH1VLG2A8I7z
U3IrcXYF3oR8rLbs/awkTm2uT62gO5aHNr5snu1DZ1pxQzTfL48dwVTe7ZAbpl2R/by8mdyiYOEM
DIWIYSoiiOgBXQCcpksD4f7qSbOVkqvy43DqfCt+mhZmLJY4MJq2asW5i8SG8njGoV14BvretUnS
1m3PwZIjY4pzIIOn/EMP/O4KU2UU+IBx10hFMb3Pm6oZbJqyFVuVxSthpGW526UOVNll7s9x1lGV
d2r0hCxJH0NWDFHDOIYKZekKzCCSCXYFV/v0jC1qQcJRePSVsjSMtXoRmO5ABToLpKqbrpGXNY2D
uepn5TqPb8z+vyIbKWPYFHTRVlTpzY5HnQRjD61nVYo4jzXuHjp7SfgQKC69LebOkqhDa4SF0HM+
wsuXn0O9q+HvPFQPI8t1B/13G5ZSeB8XtmLUD1V5RDjDzDJmd8FS5VOUBzm11ps15OG1bQmLnK7Q
PV3jfimK/5+C3TdIn23ZrxsjO52uRs5z9SheJY4iURre8H8oYLnMeTi59Scg2SGFZgADtXZUUEOZ
zRXLGt7kuElCS0W4Magz1sWPVyCPGf5421iSidmZWv/R//PF+cXF3PikBNLjgOWXiRZiFUHzYWhm
pxBWFzWMx1bor3UC8EdtriYJ8u8T4rtZRTVrugZ6OxXCoTFM+VEWVGcx+H7MxhBsYSHmEVyHmX1M
y8bfRafIe7UIlB7CbzcRWJLRkOucOzoBYWp2xqyCQiDlV5rtdAcqcKd1kc2zNEyaXX/Nx7kE6ha2
JYch79F/yB0bVJ8sn86wJeXZfVyrD66iVxl424yZYYQgZ58StfhHg3XNEY0n8m0g2a5qmdPyRzrE
jUZtxF5iS9XUAtR/xULNh6/2h9ICIJhN+u4o7eFvLwG/QgjfYz/eCrzUCQuimVslmQwVwZWeIOzH
5jXfuRQLGRPzJGanBbCrNpkI6bflsMTNXeOwStQVy6Iv85vnNIfbDtvru9FpvrjOmAviQ0mBYwLT
otjEmz74ujGr2xC4LkzGIeg7hhAxczWJnbWA2zTthDF3fGr16E8cdKyp4+2pCpH8GsTRtrXx7yev
c5YLnNlyH03T1RoRZqD4FYNbY05bopPuheJIk8n66YfW7+LGtQ63qjx8K/QeJ/xSliZ9Kn35LQb4
IcUJcKU/fpl+uciu/1aZ51tDDrUG3bxCrFprseGcONx7vIj6hV3p3gY9NuDaacBwsJaIJ/fa+l/K
DFj0hciZJQ/RYHkFH2pPNYi9dy7T+w+6ETsg8P0WwpC25tcKC62PjCe5o4Qxf2N02y7bKKWkPfn/
V9LXyjFeCmmxan4pA1tnzbFTAkUoHQQ7CFOQVse3PKFiiJPOKk6nNY2P3AvsFysnyK9kplskfQ8T
/ocAeLX/vGj03pOSN4jAvj8bE32zK0tq2FG/ecE7EySGJzNDafGfL1EJxJD1edgBw2h9ykiuLhYg
x9iYMfttDgNwxdJzgERxDHVB0Uk26O6MSYR/FYT52/fETkJB8uHb+VS//+mGYfZjNOaLBJxcrnED
HgF0RdyJSk8OlQ4bkIuTbsKBQbgUT5cartGN5AIhgvwcUS8sV/vMo7ePtJOxezPd4KrB+/g2e2kn
l6VsTrrZhvA27L4bMCiP4xoPPUQP+ECSHz+/HC5HMv0JFusiyTebrK6AnCltbenfLrkyJy3pYQfm
y5sUNaVrRzLrMmCNFJiWJQyO9i/BnMmVXlChKWdcDaP0nXSt3WE2mjswhIgxU+H3VwVOf2pEy5d1
FHJgNsx9XfLYnMDE6o31NKs2WkWCgMXNzOQO2YtnU/qHx4bawT/bSEo1vuWUqm9lqw54u/ESim+q
I5wTbG6b2XWr6yc4X3d/NJfOzukF0eY6STBgOYsPw2gmc6N/AKIfzcMqERhZyNPvoKidwISwF8sV
903URzTDr9Yaru9p11nLByJgIQGhnUDcGdMFJyR0Y99Je038CZ7YuOanOxJVLctz9JOhWgGCZNHA
Eqs92L6mZ9NGKnHhfRfVP1RYn+tP8idgdkkPuTj/JxVhiX/hLi93Z5t/cyApUicR31ZfuSfWQ79X
90ATnxJoljbAsL07R1nw2rSVpvEbrTKgOcMGg6R7j3P/boybKgmtL4HpXbN73Awn7E8HAl26E4MV
r7kogSTKzouQue+3cddDeJR4ZYAW8k86myPBrFHqfNOTwxbask5rPGh56jDZcplBmx6sbQCL70wX
eqYu6rqlY+D3caNYpk3Omfgt+iSCcuKJzkNSE1dfrjAHiLo29xU/j4ALJQIXi61o6JOBQ57hijsD
817hQrQ3QpGfBPsrBWxLDJHMmsWlqmCTnkxNyXu6/EIc5rspYv78EeARMAqcKade9ovrTdRD/+7e
+yKEN36HblgQWKR9Fq8LjXs/M9OEju0beznhCk7v3lJQj1urENtLCCUJQu6q76xtzIjNyrOLIF1A
1kQNTDwrkwwL3T3Ao4aIslwtwvbi5/QhnuC2Ig32oaMO79TtzyUSqu4FOXcuY+hJ2U0+Pgm3rn4v
RYI6y/mFHtW2wi2RnNBlq4j6NFAkRdga8GqcBGkLfrUSaUbtB0qtLT2MU6W9mFgw95Z1KpJvjrPG
U2QOTpUwNJp25hH6O21yIDsBWKZHSQA6OKVGd7aQhpnVlO+TNs4dHJ+vJi1p2zGaaIWrEZS0dwNf
ZOOKDOXQQh9ljip9Mmu4A0HH2DF4I6aVyaTxfzWRvLHVlOCb6VgebIhmwqcQSmnqs03DuGYavEUy
8VY09xiFktRyM9/wcDrqmB4M4Nlq9MxF7ryNN+p0jA3PSV2Cwex1UwavGo4mlqhLweAo/6aPFUcv
KIVsZdP3KI6IucJ6vowbEXJdf0jdOTVUhjPsyV3wqYdL4EKAj7x+QoujhemLce40OYkG6D8zgFWq
LZTzP7ZQd0nPWmp9zG3rOkv1j+hknAnlYyuCglxFM8dqhfXqRJ5fdKB3tX02hclFRtZ3vp3IaLm+
OmgIIzOTkWh4zrZ6UdnlMiw4Kbh5OJZmsRBqQ9cle0KadZTju88E0kRVZ7teKZMc6anhWVpFccPo
l3191R7OObVYdVWaTZ9clqPcN0obS4vrxcyZR3RYu/79qKIlx3y2VkEAEB6Mb+5V6+wiyadKjpoq
86HYDjpIhmGozcXEf5zMjf2Yw1vNCIRMyKkQpuoU9DegjiNRRJy/DZxbi2Wz5ST9qkDe/lHMHJOh
iO5h/cwW/TzF1guyYtLiPtTT7nicXsnSMenDF6dKxo2UhvdGoN0D+YHkvRRuAHHJXA0MBP+W9MFv
xsLiklRV786wc69l92Xgz9JrABhOQxtJRCCouu0SKIE1PymRQHUUKlT1bQmh9MYnw86QomXeLee4
yjLMsWqXCnpXxEW0JrqwB5PD7xmARWK/1+ehiM2K9TBjUpULOrkahcnwNXl7//PUFdMNL0pofkzt
gD4T6RDYK+OnGltnvUlk9zY8zDeZPFp+OSjKzfjdeCBUEZyJtsjSQ/gnErMj0TudK3ek9BA7JOUI
HJ/3Jr/HYx0KRJ+ciUmLxwBsMYO4Z5BgFcwyT5V23D0iXpxbYlHT6RhWNXr81DP/Ue1r0VJpxRWd
fns4qai7c/ohtPk8gtTjPpyzbe21yd3IZ+/3eGPoMZBCgpyN8hchfFhDihpMDZ9o2FBaluinhSoQ
4BqsOSYDW97jLQGJuf3bHsSrlZR6yz88QK61MeiP4scKuUGXt1dK4ivh0JkfDfYgMPOqkatpgKeu
0WoqM1lNCqbZyJPW6I4rdG5jB5WdXUy9eSbGoYJJOmMLr0FLOhnVt8+fqMkGd66Y1aPJx4PKczSI
yLAe6BCFtkkqKht+11NvMmy94XaRYYBz9wubqDfl9ADZ/JY/lPqUdw5nkMgC2L9DNXV7/9g3U0JK
VXbteZhbM0A4S7wX9QQNawzUidIxTtlNq7mAJe3Uk655soE5GHSMa9E8smB9ydDio8/EBrwNGUD+
fW6TOmI0prgjlqFC5Qu3VcZvOl09J0Uxcxts20x1o3DLq4stXcLU2BpWGZhjzVeCyVEEbQLrpOi3
V3XVBKeDy2AdOBCIIc7q0rqBiXJXV+zIc7x6mPryyygna92VI8raJ561wdgKV42jS/AgIp2ZZXO+
sNvbhp3r1ihTjJFI2LKgICVu511rt2uxG4Dz6nTgOBMdTr66qCh+QahIqhJY/+5R/WK7e3csQd74
iwHBnSo0dGHgwzAh7I5DtY3I+epbGBb6jjkPnvhybh/0R6KES4JHfVhlo3iui2QbvmIHSIfcbSlo
K4xnNhARD3VGp3GDcGJ+t5b6iuzmrFVlZ39IwOmX6Z6CezLeq4xCtpF+RULyGQDfHjGKZgGna+qw
fOof+lSPMRQ7Qwdt1sOeQf6NRgwXHr6lVKzhQOC6cSkhrdMuhhU3+shHHVvxYXoSFEzgSyEUcb8P
Jg9kZPZdUxPYdDYkFKQgodS0L1vT6pbYTmH/Yl+GG6kxsmSb/1B+MuwWttTbyZUa/Z+TP11UawIY
wDTMKsf889fAMwZctqjNnAtF91ZPrtCVJLqsIBcW7L3Baf31H5uGV18lLNnpywN4afQpqXngXldb
YypYnmwAJdAqL74LDxXF/XxiGhWd4zNrqlGzfvnp3xPnGj0Jl78HaMmpX/UYEz9TSDTq4pQL8blo
JSFdX+jHUD5qElqJcdy057tUzqH0c9blmZKk0HH3i6SMGPMulWyoXJ200dpVBwXYwomYMRwC4HY5
VRDqnkQPwx6XoIWz832Lxy1Wik/yjoXMCDcLyqlV2wB001x0UsZUMiFmV+BDXLDTFPD7w9uWT6Mk
ONSCQ/JiwHQzyuAFP6m+T4/Gbk9YlS4eIzSR5FrtLmYTvd184dFWfQvyFL8wnmfzOF0lWtGGAccJ
aBd1xnBNTtZHYw6oCpVYE2as8QFliGmLDNCbjGYsSS/X0hv7k5J1Yx4+pZV7n170svHqszkBNGZB
WK2/D9UIU5fQk7gjkSP9ZSdTyp5oqLQEjoE5v4ctEA5AO1HorRzK5zVdnqjr4KPhMFVqStX6+8KJ
YF3GVVdE5zOvwsWYz42qNlGNzWfk6LpWCJUVvgsUcIgqIZIRO/oeD5rq7w/0/BDw/IVwddv1A4tW
ZfUPhhVUpqJ3+WkwuW9fjnmRehX9Sx7Y4ddpjQgLmDkTKk/TrTJZ429IUjcq+JB/iFJY2SZS1XIQ
ENeoU/cmW8+FJkgnjq36YOw/K20x5djdNqXxdimpmqjfKhr1WcOtjmT7LXS5fwaH+AnYtxc1GLa0
2uPQsYVVns6katFNpLLdbha8+l6lOjd0pEpaOBsnJQnGCAA0dvJKhvKnj1Is8mP8m76mwwVwwjuI
ccMlnsTSZleOzO8RD5g6mCOe15iS0gsd0I7kfPVanHW1LUpNRcjCAwG93xPBphIIhXDtEXkBPbjq
ZO6wxTs2EwN9KtgnCz2GU3NxSzkj8WEmF6g2kzd71VUYkdbFbKYdBmU2+UFzhg1GtK1crWWi+zt4
WIuaHN9PVPoTB1s7CTHO95s0vpqkKflik7DqD6UgLgx9EcTiqvQCVdEzdNFhcCbrASBRqFmFDNqD
9J6rjqmgCZcTMrJLS6kKSohH3cMU6K3I4s5dJVJOaMmxxWEDLjYUZgCGyJfN2Q1BosG5WNLnsuM2
957rl4HbZCQ0Pq4w2ZiyG1xKbbAFoaH0Bfro1bi1vvNxlOF6fit/VGZaV0trzA4sTt5W60UBCTVN
pFP7kmN67UL12raNbiHwBT6BKFN8bXEKYqAOse/LSPF2dY8uqqW4EC2mytr3Gi1Uis0K4rzgUHV3
MWieIHeCy5vXvFQ3zYxoG7jTVUO4dzHgpwU35QXVE0Og1qqsN77HSZ5UVWoeOFKfwKV8j5aHHiPZ
+6cXWLHY1RZhboAIKXbQuC8+EeQgCa1uCx0YaG1KWvRoKRnDAbVcjijC6YB758LupCmzGAbOH3BJ
jSopO9qlCKnAZyNZXR2M1k+u5H4giJElAntdWk3ee9OIBtSukndqimznIR+/nD+ZjPK6nQgeMbaP
Cukti76ThtvSH/Vj+gJdSvHyW+eKCDnorBJPwKHhuSaGLSSloFgrZ+/VSTYlCaC/GE68YiUn0u+l
quxuNIoo4h/2PrmcOzogr6d/m/UlTty5CkkiRRhIGKg/jC+XWDIvNJufWmV6IkCTTYPWh9XiXi8M
Y1TX/uNpCUDktvNeDwX0fkdlY2t4sKSfrtghl6TYpfIYh+xOT/17XT0K/w5loHeMm92zGrsjm3NJ
xH0TUw8EwwDS00xHRhjIvv2Hwm4MbqNGcE3+rOgS1mMYS/jvMIGYzqHVaWa28j5GQMaqqhbNAeGJ
wEj0C9nywex6BmJaU22gBHjiNIh23Hz4csGziRN4e6qnGVkZzUMHoq0GQHpPRR5W5n6laRw5iF7A
nrcHYKh0Cv5zUtXQtwZi7bZbnxIULHkAYbfCR78dz/q83oA7aq/Nci35iDyBuUs0yYZ5dpm3e8GK
21s33oZz03z0QQthSXvDrTKMLnlhKv0UOm78vn9k/R8SQpwEAUCE5ltVjtzaI2WN2v7d+x9sLD1D
U1neWo321FKOfZN/SLsZTi191zvJ6cM5uMTBMJFQZkuSGNvWkJ0sjsRqYreM2Fp9OhJJQUl8KFzE
oMyRzEyUgD6nqlEMyeu92dPjwUJcSTnykyJcZS0vVXpSgEI0Kt/Wve6q95RWGoi9SxLvthMONUQU
JdAVu08ZGn85Rkc3ibP2DgYO82X3ncaK0HMJo75XJUMUGzBgZOAxXBhRo4QtmnUKqnYvN4jOAWOi
4+3g3IOPVBewYHcMP79ckzlhNaw/vlTBzpqGmRCTKqnws/Li2zf473I/dgxyWsy6zF3p7asemLCj
jj5ALIptUgCUyhS8tshHDQpTSLn61ggK5O/DEsxdGr73tonYpnvbyxxmRjXzQthzqGLl+or9MOml
qomgteMK8XIEeVxwQKMIlysOJo+CQAPAAhf1KCb8Hz+WlLEAMtpf7I15Alcx22HNHrIi9RZZ2z3J
TAy1YG/HYySf2cCUixxn/eYcBqtnSaHtPnsahZk7qTuGh045KO49oXHCD61uIyDKTivU+OE3GhgB
A7yKH4iA4PcCYB1/E1rK7WUdMaa4pSK42eLKszXWHb4FEe+DKStl7JhEb181IaCi0X3mzMXiNpgh
+q/oeSqJAAoC6Rq6ATgDEVaP3AfIXu0W/EwVHCiJGYKAxjBecW6ghdwNURmNoceOu2kT1g4IitUd
g/uXRSnr5guRcq+5O+ECSO8i9isyIiMbrAs3oY90jbi7uDGSht4fFmLaCWmj79roSUjmK5B6XVIk
lpj6e3EkRHUNXWQ8R1PnjkQyCWmirtErQc2JjEaOF11UdrAy5PDn9SG0SXJMXUmt5PbP9kVOPtrI
nCxT5mXjN+KmLjvNRY5thlY5B1e3DVYnR5i7u6h7WQYwzjvBZuN4Eo/xAWDImyIsEcGySlr+Fzq9
NOrt4QkNLGiwdo8vpBi/Hxeo2sbRt3pN/PoT+ZaQ+bo6jC0haxbl0H2bq+6eJf7AUOiksqBxAZ3B
qsyA/73dKPVAlS+EFISzpEyLmeOwklwpKcbgiLhCkgVhgFhh2EyYLY5UUCo6BZW5u0ku0oGpcM54
HRCT83jGC+WDRObZEPHlXpgHaa52BIEbGEF+S10liqjegheXDIS9wuOV7VIDWHYS04/Br3VEsHFg
CIAozQBCBKAPIjhH8jd7pce/3+U3HhrkNSYOlruAxuTYg9tooRZY1GaHu/dfXJGepe9KfxntBbcN
IWSiiiHjihdKvxHEGkvsEeyx5+hn/a74lXkw+PKhmrkmNCig1b+i7hlwFGd4qqx3nQuPvwvkAGmb
fyWsz7YAijNRzBWij7Ja523/DdU55QJAE/peiqz2wuaNYrfz1CKtED0hDqTtySpARqWAqmum++3c
L6RBlLxs80UMVTNIJavC5Pz4V7/bzYcBMOrFHfjDYrqlTAEA7/zui4QUhF3MsD9GFkjf/x42MAnd
BwqKAB4PyaXthOMZXUGXOkkJWVgiO0Oyjk1dHyIeF6O30Hvtwc/Xmo29rw6edxAvE0ghce1Ahfr+
prILVgdMfHVaMWWXg3UToPEgS0ly/eRPPRn54K9MTyUvo2Gg4vS6iQyb90NjJ2vZvpE/xmBuSqy8
xA3X+GXNRqKyCGqCfFUMu3wVy77kOjJEeChTHyqJ+ljGEBSK+G7InPXB81Chh3IkKehAEkJYYgIc
04+sr7VQ1Zzv3uRnV3S24Q80g5H4TpeH2k9QhLZOB1HckYNI0csSGRGpQ7CN9FvJY9Y8i5zIm0SY
MktZ2OQgrBM+2rduS4Ajo/uoqYkU+qJn1Ty8C6aCzE37qY/z+KTc7AKrmiDa374BZ6TRQJS3HB0Q
5HXs1LJA11oZHRq5SCmdpZnKXic6oXnj8DEYws6uaY0kNA0zreY3fTdaIK37JvHPQzKUWKn+kHMG
gIBX5YdQiXRTb0bAT6FPYlWT6W63o48A0tHBolxL/ktkIJVdQALULzAymRbHdzdk+DQ/+hYxsrmj
3RWL2VgZjREuqRlDZkFQ4TTP/qF+SJkZW94kWQloNtenlNijaJ604lMZrc99O3lDPRC1gLgqJm2X
U4IUywZTPnv65FT4B4Mb02YMZ4cyL6//ngVg3G5v4EQbwNwxUYI3tR/Ww/Y6bQBzR/hAdo7bw1Uy
xdjqSRvq6MhIa3VzGH8O2/Wppt1XIu/Crw3ekayx6DHHVqykDmpPDVbJ/wkkVBuEyf3PBqhpEZe7
aMKT1MvLZMcH1t4Sn0Tv4Oqjjt+oXOsT6FlwlLj+AO5oN633xvvqSe1SKFt8xNPVj+Xf91w21Msy
HqsQn98TZWzo0wPx+KWe31awkS1Ncf5KBGlqk1YUeOQCh/DBuw317IGjj2b8eIEkBhdtFrZhUipe
mL9I/FklzMJ6f2xuXqb+Yb5IO00I9Cu/a1+LXkrWIll//obHtg27kErKQT4Vr6vK4XW6+2gCnC5L
pKgGFtSi5iHpxmLC1fC7ZPdAVi9urmue+wt4DGyoROWzup5N3g+8QexAXSR9JCJSLA8FXQmg5RQ9
DLTLwhe854+Y7jichP1VOaCwBr0tlgwCXmGIbN+FLpuRE3gtDWIZv+Un/AQdb0psgYeibD7YQ0oZ
FaFwI1ZEma/trv7QUoZUzpwNsJbC7hF7xx90IOJIW1MCE9JY28I0dEvM4f7jwcvFjbVvp7RrvXu7
VzJT8Qdn2DhKUFQOscQwpr0iRE8R5/yg025IfkJ03pnQVzRPAFN56A+9iRt+X6ShT4XbTADkC3j7
VC9NPWa4IFhWxDzy4jV4+3ZPKJ+2STKlVnedJ0ET6rLwiAf9j1iEaFspr2OOcjJO8VUV3yAQ67Wb
cZKBe+3bKtpJe8rQd1t4iG/qMlnRVIcHRxWPs9d+LzUC55dXLISlHL8jitMaUPZfSIg69SCR9xy0
DQ1Ptntrgze/E1ID7oJk9dmgDkl8++wzKUhrexlBlNQevHTXmnZQwPaxshrZw2E96Y/sNCwgQH2R
IUo6STQZ7kSnaOqtDfvmHGaxePUERKff1tbm5Vb4E9g9BjJBl3qC2mdPLYZ9I3aOCFe35Ad9wGtJ
TAU3v2QAaTvBfv20gGMOmlksCg2GDfrW0ahn3Hty6luS+OwchvAlNSgPxNJ5zAQNcxburJ2TsYfF
DvgkC7DK07upIGx+gaqzRhkc2ooGV3/bt36kOL1JgGSZM2B6A4qTh6xKzQ9Rc2bmxXQB1MiV82cH
yzZQ+PeEHA530ze+qG3wkzuVSi8Q9C1HX32mZD8+CrxBRDTyi56QM2CxevwPUrkDl9E3NOghY0h5
AziNV8gr3nmOVCaP2+3X19cXFjPaBi4oKEKt5OCuEofmS0Sf1PxJrBSwe6nbS/HrCTMJzIu4oQLi
4pSgoBJ6Dlgdw4lZY8vzeoYhdUS/kPaolGht4brevQDqbqV41ruCFGTesJ/nxlOS6ggajQmOUYV/
B22OLKih2l5d1HbLZ/v4fSu+8rH+I/8yDItjFir5xGIiaDCmwzB6503pXvSBAD+b4oxxAnoRwE6R
QOGd4p14UX61VyRfnc9qP6LydBTaTGkhMk519/YlwN2vPZyclqbYr+jal1Lpm6MNzHVh4PNNPZCB
L6tXuNz2JpCcOedtxSzPzasfj2isET7aiFtNxd+sT37OwXuPAXzI8a06UVrBgb+m7zDw/wFKWzhN
l1U3YziC81i+YRZOkihfls99SiCYjvyjXnv5D3bjbPm58LA3gF1XD+8hQ9P74WwgUaHowyd7DaDG
powHD54mVGelMUcUgeUd0+x2CU1h+nxiB8EXnGEAI9VPvol5zB9KJRdOrM/Yju1KPFAv/w/Jz3M7
PVQ9AaMGosYVXbXS5fgnjYR4xjRtIgoFpPYAJuWYUuuS/4I7MBDWimRgnVmTZN4pkDoG5Z5LE1V8
gbXJk7FnMrwfH4fCvloWDvCIo3y1xxViRc7althWiP+sVajZWHHJeTlqhIiZlTWPaOU5FZBqekjG
1Ltg/Cnuy2xKSd0DmjfMWCp1C310qHC07are/jSUL0qh/3AbRfKP66uRf+gJAl/PgzsrLH9SqHAV
0P2z3hDjS8fS0NRuq0cLLnW5TQHleoXZTR+WwXq5/z1ZM/Jk8BJKu/q7rpBSNGisBM3sjcUuPqd2
WHbcci2mDfnN+Vds3MbO1jEPWIeL5ppWUeOoAulmKAG4eDKJoitw9nKnHLyoCe2453Pu6EJdpEFy
id+2XsHjssaPILOVW+0pza6zAWE9aGkcFWw222RUj7iTjfXw3zzGl/kDx2FZW5ED11chLKvoosDM
txOkclMrfiYgKH5Jiv2V0gURfaCWPiHLZtOJf5W6fTVOwuXTxSuHFwpZ95cUJ8/gDLj+1VQeLu67
m5PgvqSa+4VRNqm3pSGgoNhvVy61nNpheyb10QhCykgA1kxAL1u6WRdx9B7NSZyEd4nGRDeadZXd
kuv0dTYw3o0R9aUu3shcy+aAJI/qzPUjQBt6C1NU4ApblM/Fqt28CeFqS5oUh6MT/C+fUEC8X1cd
gzrcUqPKnD6dCEUz/5FuLh90d1M7mymAiBaAK0lZAhqgOVeCmv95MpWMu/3mokPJ4CdyWpVjkl+f
824dkQd2/Fsz2tVEtxjNTqwxlO7YMkeqruIR1r+Y/+AIfW8RbDV//JAHovGSrjn67yOf/BWoRZak
7Or2c+qWcgnMdqpGPnrnqZqBPbfwvvdbazolfwA7fSGHTwSIe3nCLlHnmf9ZQ5u9gkmgX2EgC+H8
8qiovxH4WE6jve6PD348LCYxCt8vqlhOh3xbZtzHD+dpjBU8y5cNi8FQNgQ/KueYHBVpDBW8rawv
MATLlrtAaSWYWR9D3jamSUJsGGGUbJJHuGiX229gTzlrP3Ncog7GNHC/tHYloETTlO/LkqLFOH8O
dwnAIVjUYA8uaIhOxEYeF3QmHiOFtwqKKM/aXeuUz1hZKIFgTDr/Xk5/CfADYHTzYXqdf1w/qYtx
ST4UIM6Uo6TGRRLhu7mx4GrndBAGlyVWHRtgrnjYZ5emBdF62OEqDYzeOOLSOEfXzL20ywxKgqZb
t1jVgz/Rn17W1C3GgUQraJ4Xu7+AVlYBINWIUPq1jedebaJwBPGgkccNbs22iADCo/dPtSwYuBhK
zEL0pFvyg3zLIzWVwOGfRjnhm74mvzhqQWgQYCnM41usVajStjlrg1N5QLDLcbKzG2Ge7HmcXVMV
tSiQYCcHMVeZWsqv6DPHDbS1UeH2u+MiyP3Jng4XaOOQcygRTA0zV/AXglU1i489LEOur/9kUB61
ieD1xHGDB0/JFW35AUKbWoF6fj6FivV9Iy9eADSen6PAcizxPAikXFPxkx8gO4o9w0LMkGZByAEK
tFveK5ix+Km5oB2jFHOyZVBAu/zJjT4+SRXsdSxU/kQKPEMh8eWhCvogxYaaCXwF9SAYIVB+gY9s
LFYKQBw/gfQPwiQzaUeZvvh9otbitXqq2IVmCMqrJf2JOkP3l9D7yQtSdXXM2o24BFMfu8Chn8pi
X9++o9eQUiEy2UEHij+m99qGfZO1d0Ht2nK9xUaGqzk1GyY3VRj9EuPMAxH7saymhMqiMF1c0d28
HRn7nX+rY6PuGYAEBbnEA2v8HAcWN+kudLIthmwlVJTAPIjst0lfYm02fKWfEeXyB9V9SOdwVE79
YSUTllknxjNuLkh42RkBm2rS1kpQfBhXDKv31bJWWKG7Bv4Cw5k3rQI3tDbluJR3Kuwbew1COwu6
lVsKcqaG321y3N8VhqWgobFfrlyRltnj+5TvoH7xt4tdl1FFI+veqrJ/b19IXqGKZykyT32CCnOf
naxeMy8m/pSHbcIHkWKmTDiVw2WhCDE5aAiGe1usHMtv0h1NLx2GR1grZmxYxVV4idsL3CNEBqty
CCYRg0gNQ007C4TyynXkjtjoLTVF9ObF92j5IaH4aTv/UgA1w0DvJP4PV80Gm3eDLiYE8sij61xo
heiR+dhtntRasxP+6+jEV+11t75aEpJ3A4IsEZsj2fc5q6B/K86zob29dK0Pib67LZuKkUGunD58
p7oEf9Q+u5/gDsZaxW2jdhDyPdLbx9UMd01n7wDIcNZAZdOjXXopn3b/xBSdxkwLqEG891AN6QbV
6/6e7ZISQyjwdGkdL6mIB40zyKNJ/6LPAiGOrOL0K83YJgouUfrIdW0Tu/6AScHds99yZpZJxphV
PHahozNAJudIbxzPDScRopZTL6VAkDcm4iLgoCd+pP2hBFjOXj5Fqfot3O3iSyFyldu3zTeHRxKG
ambCzuUfpuQTYtVQaM0jnAPnwMz8wOkjT28O8JBaZ/lD9pyUjd9JgsBnCZhYVjtSeFxpieZ8zQnp
i0Pnb33FcGfCFKNAmPkCV0+FhtoePzGYuAHjFpWGdujuL+++Kyc5eHJmGFMga7yiruzSAaFic9rn
M5ygS+bf6rmUDFcPbRXI3uGVRkUgCIzwXfNnLUU+r30TcN4jDOQk3i7ihGZeNQPoOkEHXDRWMTrf
4ECBPZiGsVa9lTV9sN3898PmEHP5VFu2eBM5ILdkH0StJiV8s+TnjthI0NrTCVloJdcX1zLp78A8
0mCGJc85hc6utHG8WZmzBLqrttQsT6tW8kSRuYZxLeygv9Ew/oEOMKKBk+l7BesypJwdNaJeuJej
jnRwzXYXYbDXpTPpLpSK7ohQRn5zeIWaEuAqDbnZkgbxZRh98HC2BUqmQLPLWYgw+yYgJ9IBlx15
Yyc87kRN90Juh2LtpZFGld0Rc24VP56woM64MdUcDXre0a03FnEzIvqtfAyeYMYNVx3w6P3QIM9C
ATWP4m1Rah3G8s2ciPpTFI+xxn+WTois8+T90enOGCH11Vv+IXyyHe8a1UBl0Hpd8ychTBVoo+K2
pWkQhsQOCHsOdKLOlYa+IpxhX36SbUlOVvHO+naK2LROXpAZrXtYMUkDwl1oK5RyFWcnSN3VRD25
dI0+4DN8r5UD3UOo0yA+c8zmfbMrxzeU6+52eSJtYGd6x0K6qakYG6zQETFx1AUvw/j5cgyD5ZbL
qZZVkWI+1PZn81+dwNDo2uIaIETx8aYfearKvva7fKsOB/6QBj78PBa1DE6INPSoEE2Uqbckvges
MyoweCBFJOlR3Dr1/FLnxLM6XrCJ7uaHq9P9JGwP+dqV3jF27O70c8lFRw4s7/vIs9u7K31fo5vG
0YuaO3Kq9bQPErJpWhdXHe9EiHRwMbwVgBX9TgmwmzFUJDKJmhqanSffbrRBr6+ErlcNhNGYRGQy
YVSGmRO/6WJwaUqNtQg59VsLbNbJ6qz3LpPL+hsynKUsj0AxZROdE47vlMO5CWdAqTqo1uDICOQk
kf6T40TcsVh9SaMrgMJ7p+IBGs8x8amwv2vOq9aUrmGdUr1pcwWKwlZLcvxavm/hJsroQ7CA3ZQD
6/uRS55z+Lw+8TfNn4r2aVQB4rK5HH4YmpxOGP9qKshOEGcPgpZj7ItWjrMuB5shno5LVNiZ8uUf
6b+RzbYdr1LPCDLE/fysbsPC4XB8A8x0HlyWV1iHPaElB+439viipthciLabEbFSuWtx362WXPjF
xlaZE4Ov/dSUOC6X99r9YvPB/SNGKqQDhBzln+sy/lZYBtoH8qi/sc6jECnTSqgdcmVAWa1LYcVV
qPahe7QqIBq7cSCVp2nLvwy69M/04pLT2Y/A7E2qU3+Hh1jjb2q7rLLUIx0IoWWbxW6aqGLP3shC
9CTyAdofCHVUwuMuyqZ1jYq7zunFyJCreV7CAmjCjT9r2wtCyMp0v5jZZnTwrteGcwbKn12uCD2F
dvcNwDbTko8eN2XBw7Lm3G7IAUQzyywP6eCWktWZ7IzcSiDq0R67VByMZA/feOvjr4hlnOc0Yowq
T5HgmkHM84ZS1CEi6Z1YLid7G6B/aI8GwhC0XiZUskEDfE6f/HcaBxNigmDoLTQSUau0w/FmW9qx
Ohgn2A5eAR+D86zaQrVe2qaDCWwtFeF39aW/kulJwnxpdib4Ztxm6BUXVsGXG8+w6NeprDnp7yqW
TkhRWQxn4S2LVjrCV4FcEtRXYMRcyn8iWsCOUVajrBNy5isDKAEhOo8WUGYUBgYA38H4TOZdh8Ge
YPRqeN5Lz9EIeeExvE366zL0rTlSSS8Iw+uKnnNGv9LHS3IsEYxPf9nSYxKPdRhuSHOB6WcZOFnV
7ujvRxMSdA0tN0XXLOpCCU7ufio0O3508mDI5QThutEJIFGDzEYKzAabmUE/QajZ8fhVp0AlJgxK
j9//teZsjyfqnJaE+tR7Smd4K3xvaynqqNEo2vVAupI41NpAETv02M8gxZlaeqrwTKUZQO8p+4cA
XI5lc92y8wnbC2/DpFIt1rwteZtZrtEFsx6s+38OAXoBXoJw2de4XN66p5R8cBONGs7Fe40TuQOW
0VA0waIkq2yOUIBMZyuMNsW2BMZy65JBls1je8wsUspIOcbe4IAMExCnXlULpo4DHqr5V5IUNFqb
ZxigUWplZs//0T1IP51fgsi3eH6yzEt2+HZDpzVOXiM5H0CMxMLYmRbwgr7D5SfknJhfwqa0J2Tn
4r293db3zaNrRCkBdaC+LDzL5BIaV6/jx4RcEIKXZ5R2MR9wo+KQ1YdqD45NucRQujY4KPkCAmSH
oEzsdM/CqrIlkzIRlTTAgItCp46cT7CFhNISeyTmG1nPoMKwKodlVvMfhDylv5WDo3l8sbNbczEs
by/s69MIfQWz0v7+Jh6ERxEup743dmzwOeN2QUNmTpLVQ4WkNZ6S9sHQx8bnWYGy0UfvGS64nLyl
NGQsKThp/EG1QB96gJZnldyAmwIFX/vKatVLav8Q+s7/3GW2PPM2NVN25GetXN4WoJZGMXWCryLj
2A9hGQ+1jcI4yu++ATzWEnJlCUupkABFpjLkfYU/hCW33NMsTl0CW7l3V3KV6772WIPtcOq7TVkq
37sikRD4ew9H6dQFjAwKu7kQbBhYPZPYvAva7nBPcSvjIlRFF0zQYz6DzhOL19Z32vKb/w+KRNx4
mruiayhv4zQzdJZqCDPAEb77pIbIeh3+F+VLYcYRe/Y8PSCNG70vN+K85Kgq1N/PgGqIFuIX7kRF
PCpbaz57Bneeapveb/tgcEek2JXaFe/vefhicTkU5JG4xItV6ME5nlmqch/RgdTmtdsM7+MxAt4a
lQIP1ZQlxqEvhS0LbNH7KQnRvC3/ZsSvBB4DT36d1570en0QaEHqWDYPFPVNzUHs1bw+VrglcIff
PqUYRc4zhwScbnaLPUSZAztqV3coqyhSfDtn7YUPhifFJ00vqCz6axIjlZRQhbLdLrnrEvXXHnVj
a/zMhkCQWZJMt0ogPU9dY9WJJ0S79FhAoXeN7kcedMVhaBnv4KsGdgN9Ah3RUkMZvVsSwNK5o8pT
0S7E3I6B2+yBI4rwAET/kckZfRz4ZLs6RHL0ixHzNkpD9LcmsR/mWe6aQUz/UQEpifISU+r25551
u4Pg6NDn+bbg70Rz4PJ3vzWcZvlhn33WcKAjDJVffAyIbFz7oDxI8YCQdjVJ2bRY5ggp40/as3mS
7BuRaZCRwsypvzzoIROIX1Zfm/8GS1RvozpUhoR+r6GThtB8d6o+UwLd2p0OkW36pPNdE5YiiMOg
te/E4YL8aRUxeMbVhHKkxTdK0BlJFiJRydiB1mikYiJrE3N0k70FBltlvW8Kz3ltItPZ9ejAua+2
Pfgl4J5VU4OccsPqdWbug1aW9LbBrH/3qDdpOA7iPBMCz/1Q//EkS6NyfmcGj6VR9JEdFBCLflOq
qWCAeml81/wCKUIAbaXQ96NMRVAQAArH8mL7WG1BjT8FfmupqnXLpgyh7dmGY5/USUqNAKJTJqkX
FV6jBhTJ81DmvqNHInuoalY2CGBQYwNLUwJ02kcEZh+ra8973SQsqYWGi3hXkw365fpwNTFPSL+G
P1gKCe+eeH2DSv4xmHrTdjjN6fJAjE8b6Qqle1uJtsZWOqqM6KWIlg8DteSqO/GNTKK9gozuJ5oI
f49D+wMTCAKBGEnvoLodz1+rlioUTqaSxTrMHy4HZYXrI94wiHwv5IYowv5PexVkYBbw6fe5Yr+4
oAKG1VZdBU8PIFB85fk1mJy3Z6i9dXDi+2mKHbT0E1XHIw2Qrc/mf4/ZtfueUBbV3x3dxpAIE52S
toh0HUP1DO2hozqGOwOqcWjG2jL4GjqpgJcAsi7/MOKJ6cxN6/04kSHEnSNl5JUvfPRbqbIRDfGb
cYIlVHKtf2Ew3xsNne+6k2YVwZ+4A96wmOAfx0w6B86DxKbOOe95dJfvWGmAm0t4hBwQQA+7uI0K
OdfM/yjw6ZrjAlh/NHYOlbktd5Pkgvj+NS1G2PtlEkTBvGFOQOc2iPk+JVatUOnzQW1KrEj7NBxS
Zw0phVzp4U4Vaq0/1/OMTyI3Cq3iTWosSRsF2XZviiayp/xRFMjqj39OGj84em2FnZ1sgsbJKEYm
/kMg3COOhw3kaIjC0C8w+trbmofWBernXBnG1UnAD/Qszg9sM4cLoe31NP/UpgyEaPkvx1HXQUC+
qvIKFyN4rIuX822Op72vHLKCKxR1m4yutpmL/8zgdWZbCp9b8q6vsLavChGHztSG9q1BGSj1922c
g8ckdv32nk7spI1ru201w12NvMijQG1n2QwZLKyl/Xy8rHTpzuhZ0kd//iSZgU8dTnrVkkCFRXT5
WD/vglZhGuzUIhuYmgKlQm0q9WIy9OwpTbA2X3mCWQ3RPUSmVDl23U4uCAfV63i3auYY53Bob+6y
kIj8hJunu372iCrsX29nzPnw0CfdjZ8HbB2nQ9c6yyT1hAKFDct0xyLlEBTY6Dsn9XugDeCvTktK
SGbWygf0rxtAoGyYAXV1HGivjbKPF8bap9G+TLiU5qpF4bId7G1mWZC6/nR65MJXo7rHGRlejXxW
jDdRkt6drtCvkszThptEn5dD9un5FS1h++w+90JqdWMzPGAytqaRImdvDPClOkN2PHrxL/M8yA6f
EMsuPNvVLPxt3D4PVxNqj+oaMF+mTNABNq2EMRqBRTD3szA7J4r9LI2GH7qvOcEu44FLFYJCFWoy
TapbkUI9tAitHGhisAp7StiZS6Spcm5LylOr3Mz5x0k2x/i8yowwpu1qdSGkYYtIMUjmjQhVGTpc
z0chwGKxl+eLGIBxvHEXOjQxo31zjAMU8jkNV+rK0HRVlKs85Swqg7fiM587BgkTgodfKfY4w6lE
lrboPWIHiSxjDUAt9bT/4jF//XlficZrAosyY539B5CV5vAWv0T2TLSDu6qumX7pk6tfFrgnp7jW
cbwaHfOF2BIgCe2vmKBMG2gsC0O2nCvLhQbPZUG5XESZGLly084TVTdNV6Y+cjgC2TpG1ZXL22m4
HlqCffhb4tLQ+wuj/jXTOF9wfeVVfUsG7eu5ZclEU2V08FYbRJA+3uxJ5TfDX5cyND9JX7jQy/gw
VdzZQCUPYJo9uQkFZBHZCIrBeGMzvSKRrLbixoKzf84Ti5MvzqeSKixoZDcMBs3n+E0KUJIDEcji
5Hw+DWcfY2ltwX+ysNGlEOuhtOsqLcRcYmLbVbCsjqlC8ZRXGN6iU4bKzjlx4d8l9nuPCoTPqhT5
rT8gT40LhiVjXTpodZtHVIfSCF8kV04Ny7rY65g6b+9++SuhkdRy19FxM2HcaBlKJ9q3tU/j9OIE
rItv+88JZSJEx3jgbPj3l2zAoScubki41zvTXudVBSoE4uXNE9zTFUU43MwpG1AtRvfaZqT/VwrS
xqac0uwa48RISAFzzCrEmkzRVdRUVHtXCCu9lzoMGhoyc5d+kHtsmj/aUdXAkelEAAs58XyL1YD4
uW45mU+i4/qNqbbNOp8QdUsNBx2I0ECuzKrJ3WD2BkLVaGHgKmmBQCLqVAkM1K8ulnQphYvZdCv1
4c+InI1Z4UyzE4uwP5jhyneWPVKrytWLk2GtrBmxvjIYXwW2ML1Pn5MoBCTrkFsAJOvIs19YfpkG
8F7/LK5mIo9uwVny9CW5Uohs4bPldMprNBJKLfkCe/J+W8BOXQ1GUF9tagnUXNjdG4xIq0yERodR
N0vikQ6y8zu4vxjDsFyhZ3IEQrQyhnH73at91dvnNv/V4dI7TK4GIeUHy74TV6PLofebjXa7ik3/
wJIZN910PCYVKZUXV24ON+mWlz1I7PPwNCKMPbpiWqmg5oX3aIzCZaKaK5YnrgaQG/acErtZSkNA
HPZYNu6L9OasM9a8jZ+J/mXPnWkVu2KD0U5mBgHPAZvmHQno8QabuKg0EuUyxSjil8layYdievOi
KfkuputiEAkc4MpM3ur6s0cS4S77yvrLcpowrFzyD9bb63kQeP9VH15eyaP+dyuHVOvsTshXQi2E
BV5kQ8rOhRnwY5U4EH1BuVWlgiTIiO3NlzkPfB+mMMx3URdbc7ejQ5ojH0U0PZzulaN1GElzio/n
HMzOvmEeOfYpwsm8kw32eMFPF/u0bhJSjY8P5O4kJAYBUMtA0Ko+xmQdIHeEldwIKwqi5VIqtEN4
QhRD92PwSwRY36BD+fsLo525nvjox4J5413rh65B3rTv1gg/I8oypo9n/4avV3kgj1jm8SRcAB++
96yeb4NWDJ6bil0vbSnYVo9Y8sm5ErCNgUmK4POouiK7rY7pAU/I45UEWTZ7iB5k9lY1mfVBw51j
TNxo2O9iusd7FZZnbRZdDt3YG6U8wbxyzkV0DTlH2RHX4Q3G+bH6dABQsOu8UCYmLT9RB6tNuyzZ
eTIvFYlI5PxYZ3jxzn5aT4PiYzbHqPDZ6+qEAf6v342DsWaJbq1Pxe+UQoaH9JcZutEzNkzKuAB9
tjNypTGg6E40cn7hynqrBlT/UNccSv3cIm33F43OzTy/2Nwuy64ArlJfmqMziqADX4tEo9+qpQp6
3PArwIWVMRMBhiEE60B5s44WyS+II7SWBTmvCNorojy4UL6zbUc1X6bgMWy6KYuGLHa0HbrA1NQ7
YRVE+f1QzdLETt7s0x6tyULZ+C8DwKTNINHHAPWCzHnJiRqwjuVKkV69vkEnxM+d7cWTYHaFk8Dg
SO434/T7MJNJHTwyWpWlVchL+Qef5Djmc0K+gyaupsBqJ37BSNrei2CdnYTK6BZznbuGXwnkFSvB
HAHsjtByKy68YHB0/Xo/WK1jyzgj+jM2mkD9cExmcxBrmiv9ztFeMmyh0YvqDKNI0NyL5lJ6r5ug
vpEsqgC3kaSuYYJjX8Fqf+OH1VWhCs4Tdd1n9ooj85dsx1aViT2QusD5uFVvjX8vc3g68FiLOyoQ
Auw14H9OR9euh48lqnMkcz9Tf9AEBGgr3wSw+/e48GckJ5TNFk3XHs7A3sG8vCD/YGPZtfJyzm56
aWi8WFsXpbeQm2rgzEvg0ITXL+Y9S8KQADuQ8zrotiwLD/3UWehlk+luWtO1bGNP7O3+DTqcexpW
wlZx0kyjIEGnVvpWxamyo9OdQP11IQEl5Fg92qrvqLG6Jc0mUyQj//k7hC6JhymUmVywNbWW827S
GiUd6VO2yxdA65t8ndmhGj7WODRvNvV+yKJJ6VkG8ZmysgU3I/jyseH4JPx7wQO232TzodrNT/5z
ekeOc2Bgpc1WXp8SWcuyJuvf2VWzkAejyTZ9YF69UpOXJ/gHMILLHq+I2hV8ETCn8Qtr88TwKwPt
3AhDHPCLRAjRctWulcUtpnE5ZL4gT1GgcVKQxgE2cjlun+VN7YMavO+8b9AiQRv13dfoasIcmEVK
YT8nn0GyL5x6sWa2D9yagJXkvS3/D2ELROjl6clxBgRjYnV03xv6pnNdp4FZI38DTSVne+xAMxSf
wQXdY9/QN2gOLtie87EbV2tKEkCMZs4QT79IZonyMI36KOpgQsUxg4NdAvv1dk07fpYmDztE7qVX
F4xfzYuWgWLl96oypKJ/5sYFJH7zDsXem8/5GYESHi5xOF7KL76VbKlK7H0Bnavzr1N1kBu3zW8f
OGICxbrTLzYkcPRm3oHxBY7lJUKpxVQB9PkOCzfx8HlJf4bXJ+aBBCfC3AWGtU1kpYW2FCwiYkvV
qZUxdb6EBiWWiFKVOmLBdRel5xNILPNgdB4tEt+J59ri0Ub4f0GjOx8dqHpLMC5vh6avDevmMCOo
6zVrvlgUzX+KugY0lBdYEkFs6DaNtxu8WTcSGrCtROH5nJsOlZCeGEP2mYHt7CMvovqAjarkaTuO
3Vb0R+mcn+3jKJshVRUyaEKgrZzAeMov8pwAEv4BNuHSj30M0yQkC7foQk6ZSGdCelTBXKD+H+7H
Zc0zO8gY7Ps0UXeEpEF70bhp+YlH8LU9t/YMNGFocoPUjztwp7PaP90Gxk66tkS/9JWlhZM1Qf9u
ww+amzqRMsZPyACa67AToEmD5aA49LeeRRnDj6l3aLU/Q3UOnDEHpBORoAX9jYaFUl/XOVMcGMxk
uGB/NZS3sProyDY8o6iseHyYNHWQR/KkgKeWc17mw9qV3DKP5606QEFBrLkh2Oh7Cm+YC3ftKfGK
nrlJDvfaAsg4TY0DtTLMUJK1URXjj42o96hO5NwBHz3gRAAqBlgEUOo9R/mO7z5u36Vzvv/9RA3+
KSCbhKoAc3Rue/YmuNg9blbYnDRyHB2u2KHVnZHX+n2vtCrzSTJLWg85YOyeS6TdnwHs54UXg2AC
zqoN7ms562XgnZMMdl9eoYv1La06nDVIGQjD6gvMZgaIN71NvFZ1uYPiP06IR4d2YMINNTuU2Xzv
u1pwAboxqxsXt/X1xsXKOXajYZZY2m23XptxbkZerd78JDGfi76kIoQqt/MG8m6bGU0uTLhaRPfL
jyJrGn7+5aZKrihBPsDEzwVneWVCU/jKns4uACeX5EzZyiiHbaNbpA5kbSmfWNF+Von3yA5yLfu3
FUpaSN5nR63yXW0ccjgL+zNf0Zod2ZMiQVpNxWq+GXjV9q0n46D8wQW3GVbDFfaPo+jTpie8K9wT
Xhbo15ZmzTZrHdU6fbAJUyWmQ/89Xzuk7ipkNwXIHmy3fSzzPSp+of+fB39HvDPqoV9gR2KjgEFT
KgFeFBGtgOLsbXM4DJn5JdE5uz3vE3xPALHiv9SbhaKC+hdDUj2WVYLA1fP/67APwEMsHj0SLwlk
9Z6WM1PZ6b74VKbw+5Marmist8Bn+PeFuBCbOH+iXRJ/Oouw+nKZGRi6ZS2J3UVIhyATOsPn6S5g
nh+hwPlZcTc44d+yX99/aiGQTzfwlfnO904tyA12+o45VwkZ+m42/GYGhMSMgzSrjzEedk37T8SY
0qXF8YBQK7yYlvqWUbZE+21lwmTjOp1sTl9xEQFT1zxvR8YO5EUWAQ8Fc8erwN3DBMHVp0gcOAST
2VO9Tz+7wHcJhs8ifPjFu5oVp2gGLrBqa/sHgAad3HYKZeNHbhNJN1IkWEYoDezDsOyEXq0VvHBO
sOhrwwVQP9pPBF8z0j1x/TgDa3HXdxj01FZKVdZGmrIqsSelxxrUVRriFF8OoC23CtSa93d37PEu
hjF5oadQvWSiFZjklG1JvJ9ZoobDqyku9vOYoYPSodgl/4ekCi2MzM8acTaS0ySbU+r7we0nMUVn
Q28u0WKxECOPEAN/Er0BvlmZMJcr5qyxcJ9QuRJ35YP+3n0E9bS1q85ibDXJ/IOUACZM+nGsymy/
IM6OJYsIXjGvHPBnz/79TpWkIEJzoJWnEdfrujkDJExnCnhkcjY/vOfYdXRqfuj1mMqoHcb8QYnD
caFabrgzbhZ0vgQxGqePyKKRdmA+WGc4LdwDf+ydNg4s1GvkGU/rW9HfHtiXOTRqyqzv68ez0+AU
x9FSvMkE3zaXxLhC1nJgAjdJQElYPbOBokwSxAC9qvR2vqGwXPDjEBNXoHlVMoumhOFhPairiii+
vCpA5TdrbaymWaVnAW3wAQjxsQZ2ni7BNmR3w2OF5tKqyO2vzqyFPrSByCvk476idCq9dlTuUTKO
BmVX66s+qnsaX8ZQHvkhNU4KfcOkZdC4CbLcLpciLBPOkQoVJxHQ6JMw9EUaj/vbOEQOx1U0zBhi
7yO28amF7/yIZx9WmzK3mEeKUxtL/3rQa68KtX3u8aYLytlVCZGw1yw/Fq5C3VRvp0ba4vbT7XvS
fcTQJzAIT0/YGdJDSqOAnKa64PEY/J6wx0QewwzmVtU8nNeFYd5VuTDQDiz91wG4CqXwkbk9CeSF
Qx76F7aVEqazQOXvJPyHOpnpMuJanLCB8uGCeFf7n/0an+b51lzpgX7pWMgSv2/Km18vxFlPbgLT
sNOsGf+FRcsMCAHcffSkOdscqaiRDOQoH3WNLIwbvzJ/kMhq1PzO9SZVNKcnNA+l03I69N/FDKrS
nOE7NaRbXQlJ6uLORMt7fEHWUAF/vSt4ZunDUs4ZCuzajuprHhA5mFtIgcZsS8Ctpsts/CPZwEbm
0O9ds9dyRc/KSm9GGnTEhATbsMa+VrlIIMUyZa1rcWzSuhCsFIy/0xVsqIb7uMRR8vu7lr6W1dDe
Fo11nYTyvTJkiGTdir11J3EYXm+OgDl0kAb/C6Xa/DPgOj6RddY1Hj9eTFiv7KAJU1uetAT6rcT/
UzutZGn2ba/yLn2gj2JMJ+Q6hPsMFqUtHPs/QC13P61Csc+0lz2PFnXA62UsgTPe0gGvQaB8oW2n
TjHeOhm2c/6lGyMPWG9rtTMJIG6pj2CuoShF2PjLLKhgxPzXhg0eewaoH6/lSPmyzKtK+Ih8+ez2
hiIJqPx2uRRxR7s4ETbToT5YTMlc+PSpZgWu1PVOOMi13AtjJ/IqVlIHzDiKQngPjmYf7YnnpcVc
b84cqUIUDR7UUI9g4ptfQy4r1mpFlhEmQiuudpwj6M+wQdkQc1Rhk6O0dgkhTWFVoHMwec3QWnbY
AY/4ETleEqD8UglSgYV0QE1zRpOfRC4yaMIAlmdPni08wrixo93KgbuFnfahzGQ5qnSRxKLAjnao
CBV2EW0Ss0meGwisjS9ku5XICNEmQGRxkFLT5dCj8XCIDFwy0nFnqdb9Ckiqa59mDiBlEurhnNRU
4hXGJQ8odFPaaxJMKPOftOnnbNJLjyzDv1BZ4wvCDltgB581VZU84EvbryyjJl0wMBVmAVi9uQT3
eOOYdfxoserffCBcGRIOqWyaKTZ0E7w+4j8p7Kr/75aeKUXm0hc0mHBDqHnBR/auHscr6UWeH1sq
ji8TRtPx0MH4r81pK7ij9plcRpDRN7nKNGwUADGDCxl+NH0EQ5qyEDSU+Eyi+lrgloIWwy1Rs2xD
6wWybDQ1J1Tj+egIeFA6pvmC8ucyRbtqeHx3NFkxj99YSVG4k1W/SuH+RpDnRgLa/R+lbMPA6aPb
ZmR9aAqhE8k0l8EfdfMLBXuksHE9rEhz+4Q1N9Sjw9vgnYrpKvEq2Tad5MZWcCsvabN9adHrbJg/
Ito/VP6G2jU18GRfGcYRjmG/NAi1UxV4n4RAbeZBcjIYA56PYRdq+GJul+u0OHAK71FdXLX22OC5
RgTtaLkvaC0lkLeeyeu7pi775Hg3EAghlRSFR1iU4dz+IT9XDYnYiGIkO0/pJzE6uaCbOUBg9kpy
G78mt3IJ9hPr6E4oI1yqe4ci7FHdPS6bvKwixpOMRLZ6W6hADogCd4SPeC/1M0jQZS9rk2U+2TfM
TX66oIiQq9n4Vzy+Ahwt0k4rplo8BukQsAIrTG/guQBhyM9dKSd3KlJFylaVr2n4+C9npygzLfpn
l2AIQADrBBZ9N5RgUmDL0kqYsyuX0SZAow16Nn5mHt//2+rVIroV1UjBG/WXjzN6laT4QoPiZnEX
PJ1Kr43lGz5ZdXxuC6lRAILHp/aFGoT0kCSFZK2kYyBTSBAGNXhJhzbinWmCGrlLn/msrzDsSAxq
8RuD5+ug9eMMcjal5Vy++S3lx4sa789yEewNLjPxo/WO3zP/Dt+hfux0KQzfDV+15+MRCv5LG2zm
1aDzHiHlmNgSLZo+n9cmtsNd2DlE7/y+DN1J40+/Uaz9ElmAAlqVJ4PbMkT8bpYZSlGS4dqAukid
bEnC2aanIKkzHYclRIIcCwqXkPv84NwSqB+ETb90FTP03SJ7NMQJfgbu8tVcut9AC1yTfmsNmJZt
6uKRjIk1BPxJIV8FNKrR0ehl0fKQJS5BCvzHe3yQe+5uFJ97FgcwbmPGtzfoqIOrPyTEKPT4iTmF
clMYx5v3lY1Zk6oL5fx/oVeRHvfSDypfH2bE8FAGI+e5I6c8Z/GNYwri+ihoyn2GC2kaRwoNrOXs
ETBF5+RwYrukhP1CqD+7v6rfpfrtQq+iGjSsUCTLEoGc5WZ0THq5n/uB3fYm2ZAh6P4ZNJIxpd1D
AULs5IHEE5A+PO8Max5gv1J6EYJIGxj7d/qk8pAQphfcLEM1pCkp7P61ugiOaP2SnP6FeKEJHbYl
vdYX9SHqOKv6+CAw+okdT9/8DykfCrpfp+6wE704eGqgV7XxjeHfksaj3hytyChju5B42mHOMcBQ
6QMGvD/dmoPSkaKlXhsir87YO9I00z6KcXlZHSGhjQu0LGlnyoPvDRIUAF1k7vXFsuZVRf/Z2LTH
1RevClRboTuobQQ6TTnT50LFUwd10COwKgqdLdZO3gsZgcP+4ZBBuBm16oZaPgocP6xb7Ijqqd6t
kw6Mql+dVYPcY6elFEWXtff5qByOAhYzsuxwGzNywhnx8yKs7Pu1GkjHeJaL9ixkjpv7Cq8vTEwV
4h2sis4qazdoAnK9YoXKL31gNcsrq6dJw0ADBnYoJzd3Y9tGPI/gqhE9pxuRErymFr8C3dcUsVJ7
cJfl+4f/XdGbt3qxD6tPdBZNELcOxpiKz6nz1LEl9DSC8DlrEUS2KskAOT5quVXckv+qExFRdl4A
vP8z/mGLA92WbkJ418uzI3pcFF2kxMXYF03SNOegma5hYkWNgm6Cg73ZKv+n9CY8PHQXh/HAefIa
r3ICDy+U1+RAuSSdsJOYI/UPFltPNAsPyP++91n7NiiyoQKaNf+0OJaENI27qD2lPo4aRj1gKCYu
KCZjhmqr6gdfTokMVUoEPVc6d+PngwSaXXiVRneqk/tGW7DzqPLd7+I2GBjLtycvUYXLhUhPYBTG
qE2+oQj+hvreYmdMyOQElJ+odW5nEc8ybUmtdaPk4A9YnZG058YrrHUt0gmY2ZzqGALRtiSAngsC
JhoIRaZ5EyAyCVp9Q+ySW7riMNohOWjn2iIK8nbuqlaUqxhimG6ZQc/A2wUCZILPT/ue4lAeJtDe
HTGHzFhW2Jxj8JFuW/2ani6lboJfQmGgD1pXnIvHMnF78gUzxDvWKDsqyv3J07eGtgPE545eFjc/
qHkxEbW93VDZipf01CDiUoOpu/RDWCjF41ZlEx8QzgFHgjAxAcegocG/pYHDEWzgBRaMwn2igbFQ
qZiYo8SVM0l3YlF3kfAAqgO4I6W2C49BXxZgDTw/viwJzoApm3pjnHUOLY8LG4kA8zAEgZEXXwzx
Sw2O+uNPGCP3PZQkZ1jSlvK82yuHLwoZ5iY4RzyBTMgAhGqG8jr/uN4UCyNyOL/AXUvm/+0N+vE5
1xeXl/rM7OMXUlN9stEmUndmftFQwtdM3VkzrA9j8Lh8Jww7j/PRoLsiWw+1so8w7TJ8BOMEx/8X
lAb/g9YG6BOUTQpj/Ok4pot9OBPzNjMkPCUeWaIhBOVSkr+/pFK5JLR61ykryOS7hoC/mNY6pYvI
UwfA59ZJmXRVF5VpMAwXonltpM3QrQdQyM6tbIASUVGKGZ+gyhCupiYNAHa6NunPnYzy64v6V4zi
QqtoJ6bRmLXOj0Z0guSBQFmHJuPMNWhNRqLLCRcQbz/Yf8ee5T3BMY0cjIqenpTWrnlPHc90AMh1
Quva4Q0JbkE4RZJVeVBmHKpH5AFE4kKolfuuewnte8g+3QI7Bru9tkaVdSaLu32+2NQDd3YU0z6E
gXsJFoBSFhFnM872cLe+UE0RGLlJFV17jHY/RpN+6Sks6wX+s0VDtnnZuTOFz8fsiZz7C9FkH/Ce
4WuAATAFETxxcFsYSsCRC5luUrAJ28cPbvRtL6CbhsGXsPc2AzGJSJqQW5ezcJr92N/Dd5hOXZog
d51vNZXl0rfjd3gQsa68JtVkz3yKoDRi/q17R9EHVTEH7yx4v1vu4ggd+EgQpAMOF+MO+s1yvGiy
r2E8Xi/xEMvvuxG14QLXizTgE73FU2gqmNPx9fQFWG82lVGPy/sfyw+qeVWGoi+caWcQePK1gK+1
F21sWf2yjfBp3dmzu5v1sn2uNKcvDSJnBjkNuxQrkABfm9PEjsRj+bU0op6hc7zlT/4OtSiRahMX
7zdAxZPzVHNZp2N8b7UcYkst3L2QmfMYkRrH0EUAatiOMxxgNOqWHtJ3ad4X4d24cMg8G+OeMuyz
A3lYLGOA0au9m1v1rkGkSwI+CPeCvOac632b8fa22yFykYogpSoEfY0UuhBEqyo2pL/eSqxW7AGE
8PGci8kqSudiBwddtWY/X3iJPK2ShLoQM3H9sQ28zHHK9t0kmUaDQepsdb4ABJx7aTo1LWneFbB4
LEd1lEnHqSNjiCxYKpmbrzwXU8FZiWmmMtFWGw6bMdwMkdM/AG6q0OP/NTQ0iRcNDdZT7tMSqvRf
6t6nt/s8eaB3pbdfX3hxQ6myWzJ9TMNrcMVYeGwgS2i83ZSH+hsKcchV0Nw9Wfm+4DOhHH18rt7H
Tus/bGbsVUfYiQXTuuQKFheEpnPka0yCAoqi1SKszShxH15+Ccm9ykx12yA8ZlqB3ER2YQN+ucZe
FdvVXkpacjYWV4/tHivq+eS/WWb7ZPpqaQiJYc1zb358Jv4ktjl0aM6Cm5d5zsj2g3H7HYHGsVFf
2kjgGS4zqpRldQ71pq0l4qmnkJk1Czf8YuyyYZU41ucQqwWrL1KPNdy2yutCkVgfdf36CMwOjEia
5KMaGNKUub0eiCrwCz3CKapiEbea490Ow4+foxBykybMZeNIjNOC0xc3/cNAdnPd2TztORBSI5Nm
tGe2x9t+/3s/GJUv/eD1j8IoSXbjvY4+1B9vTDJy5mjk75TmS4idi64KIgV2P+DV4MOl1Zs5XqbH
r4BNNChc4pUFP5th5R+aWfyue1AVgqy2gvdv2rqHkBfIQLpkuxmA/GuDDnDsVw5CYmOqhGTr9fFN
CBw3tFFBapCQMXQbh6hGtw3rz2OhaDUEuOYTn0rtJylrD3w4iF82MjHl2mCpaCEwQZSMKghZDPeK
vinyi6NlCrgC6L6rNTYO1fdwZwhYdHr7PNsQRHxvm+iiBGjdxo0QfGllkMC/oNN4yOZbVrLUGsd4
bd6+J1BXxNVr+QQYkKhrJ1Mas98Q5laR3sjCzIIAFfKoMyIc7YgJL5M+HRXmZei66786hz8xLo8i
BsdGsO8wvvKpMz2m8O9U5ktwFMNIb75baD2t44ecke0DInPnGWzkOIzr6fl++OXMr666sb7o7HG2
SGfshxlrFmKQjCIo58ScEae0WKG1m4URIYQ+2RxIhIXsZrRm1f5GBw1Y07vFN7v8UHdBwFn3VcVx
rahxE9FY2DTEP+cyPUPWMhWO/FhogiAqfQmCIsaTC7N9OeP5rQ1cFfptJU0tk58FcJumGWDW73S5
yiVGg8Ls0x06Bne1swelAEpq10Ojz5XbG2oEhcq/montftHb54LSzNseuB3iSyA3WsvUqctgjqwB
4ljeRbVvGPZ6EYGOKgG/uycHNDZ2XzE+hKl8Eai2YAJjw6EyuK9YDmmy+wT744MgxmzT462fS33m
b8baLpB+ugpkEaYgMZkx7aDYwYntddbAQBdbtZQHbgVbOIHF/tXl5z3C70uDPrhbGEiiNRJS+pk9
zXv7GJxiHRIB2OkR5UE+hu6RHjPX2JDZ2KBRxfWQB35BFbBAVhzU3/KgDxCLaDz9d04z6DW1iDsk
MwYPJwmppNc11bw7X2+kDDZT8UPH/Lkd6TERQN0hWQgY6gMmrnctmful61U6u8vcELJfs0xViHMp
ekoLe02Qsw0wyhWOdLkjz5xZ9KJ+PF2XvBRLnBW3SXU2cm8b9ylc1iw+3mkmFNEeAhlIIgmHlvJg
NoLpzrtxR+EJSyBdHIXueH9HgwDZBXEtUW2jux2NPmvnOtgF9J8C9VadYcwxlyfL7QTOpyYMjo/6
RJH7Q7aTkZ/uxkkoyzNFQm2miVHMB3IgOkbQLfzvZh1PZs8HDH4j5mhKjdH9+I9/ULMbsykV4aby
7wjKqQfIRPs0NEfHcCm0L9f50yvMDzdMy1wU/WU4g2MFPOChAdBVBn9vbDH1OBnY/yy5SCjienEf
M90Serg6y4KnKp7FuSXARMBVFLc03ELejyK4IOsqYgYOJ3RdTvl4dLVed60wghIATb49HEQ4cgRu
aiLTztsztkHI/a+1PfDBfITnjxmSRoSt+uVvicrpUY0EVzhujg5V2jdnga28xldVCZMicSxTBcxk
JPpzs2MauH5hgfZ7z1B1NAl2BGNSBKSVqVten2SczJY1jC2UoI6C/QCq7mlXM35kQvhNrsBA9KBS
ImN1oUJ0enKad8H2Suazp5vb80c86nxwZK1X+eh1CMZ++wMjUI7IbTwsFPOUprVP+z8l1tBOY4D7
a3KKrqN6GjiE+36Lc5PK1qIGeefIhNeYrn0pfG/GB5IPMjnUH1dAA+Bxp9ql5DYT59eO7iQ8kd8S
qI0PB0vlRsseZKjEAQTQsylYAqt1h6pq6mWgZf4imZY0fFv+HgDyqoNl5DCC9ND0ZCGo/HU3lp+H
Ci3uDN54w9VFqKIuXHyaQ1sztoq4lvF97Nb9jZNwtXRU8xntdzW27Hoz2QFzrpV17FJuBpFa608V
1v0tSyBoBIlXiTadMN8pnYImF+w/2RzRqUohB9MPgEcQB0AWVpAFjAEEBaKmS1QMG0PnHOQ1HcjR
76hhHxyeM45UKmf/U94W/JEMGwwfR+bUVA3oAa+FSqMwJD8yc54I6IhzhxWfD73lJJV1ckFXFf/A
lhEY4Kxa0xq8jShsF0wR5MPIGQsApM2xkrilHV0Bog7lOokCRyCiHPqKewhaXHRMf8aALGxF/y+H
MtLg30qXP/IOpdY9mPeNAkI9v9L32i4WOqwcIqIS3mNX5KpURgGcVU83cb97qtsu+MwO2hN3nNHr
3r9DXRXSObi86l2ozOL8itFidX/3jWvtmEAZQqt802IdpYUbV32NdPYJObl39tdQSuppiT89R9CV
Htk3/3UwPlW5ias0KkcCG+F7KxN167rZIUvGHZuoCil7EHS8/0GNSdF3Yax7+DE7NPKU2U3Ty7Zu
6W2uCQrIKH330sEJNp9oRHorVGC6tcs+BCFJ7Tw/2Bk8uQDmwEkFAIst0iwU3ONM1DPh89EBDnV2
CtUuUtpL0RKQKPJBtmKAO/VTNqBxxNjngYmiMUiMxSAVYmMVo4VOy1O7oQCiRU9OS0AJnfAxW+Ix
cSCmV0HvoSn3XCA2Zn5q2kAaQn+IQ+uvFpYjyP389KCvkYDJ7wYC7B6NDtgERxx5nDLws7RA39XJ
D9EkA7OaA4A8K1LzckAi33tbewYsgy8kpGE/uYGwH7PMfLmY07/gMAdSC/DUL3PBzdZrMlTF9ich
3Erof3moygVrwAs7SQdDB2xcNixe4TZldjGD2ClGkmAqjFRFZTh0KtL+y1awVuOv5ego72rIGr1F
7cnrziKm6lGG17EAtAuQs2I/gAQIAsjf/VVTdxEXXmXBcoM5Ocg3x341S1FS5V9QLQP6ecsVSQ+Y
Bz3+rxx21p8F4uf3o0mJqJI/OJ9Zng29Mi4UldJGZA1umxDCKFaBZDMSSjCxOYJdOOzE4rWlzsc6
KIQFIgc8B1xpdhzqKxKRPYAWa8wOqYmqXpIF/aElYa5ggWhxTmFGLyzq+b/TjY7PsVD0pUzo1IF2
whENJkHrJlp2Il/OwSKGdaDG22nyDnkm9GvRixP82O3zL+V/eFkRisdrGiuNp6v5tt5YqGgzEs1n
KE6pDGZ9xN5qC+6FfpdXG5yGuYRgFY0gmgjaZ/rPWCsQtsaouqhihXhKxNHFGUF8FFKomV0BhwS6
Xh15tGsFNnwIKkrsWPgOG18o68M7eACNaGyi8xZmK6sYn1+EdcaZtKLKq6FJXgsiFwVIPSzAzeMM
G5e2lcE8HuUACyADog7uln5uxdBEG2YMtQzuDI6xiQAmqjMf/ITIIbzyC6iSVG4g50tFaOuPIsmn
fS7j7GNVz6GBnfMZdKHH/bxVONzI4/QSja3hgISSEFW8N9Iz03Ffl5/Gm4fvxp3pYziO0ezJM2nj
lS5r0Gg7tLBey99KFwQIy6lNec8ndEfF3q3uFru4YAhsjmSTmiJQO3KMjVAZxYwXNxP3Kgomc0iu
STYSYYleRu2ovaU3ij94DjOlGNZSlafvvACPOgfIj+/TM6oCuKY+Wd8J+kVK2ZTA+wyCe2puFnI2
yINu0R7rXwlVVYOTteZAiEQnXzAVF5YiuyGNPOzP/mIj4HhKybFRLKV8u4Bt0QgOaCzgeoE8FzKn
U6BvIxk+i6IJY04z/nhYUzthr14MwdCiMacIGMO7ZBAN4JzerLmI3kMQLqrEixmy2adeYIehOn5Y
Owo6vEcggGysRqN37xBBaoQDNA6P1K/9DcUfR13heNiCEF3Gbwt1IM3gBl8Ak1rmTSNXh3S0cH0z
XWzqdtmSLQYeDQUtHxMP2vyl2i+9gdPKMjaFxWV8WDcW49HYoF9TGFreaKL0NYu4PynXzafbDG6g
IliToC38+loxPsEIFsAJmjoOx7Trsb72LD3IOHuMnWWKVngqpM2JyZ35dl0e9ODwbTeguQfeaQgM
eV0SoJMiZL1ZzSImWGy0oQzrB6pb1MxQ757kW4+eJmG/tbrCkshaEahws7a9qoCNcXQJ0TwvTtV+
gFqa019Pj98nKygGPu9LvPREZVQ0UX1pPfiqT77B/3fLG0rF+o61esoVPCkQs3n5ZVHT2MkHgzvh
UI0iLFmB+4YfBxAzttqmI+CZ4jJpGooYU+tjD8RyY5vDwq1RvDZhOddcAxfT2sDgqXPD92zyaby+
f5Pmxd0g/EkcLDTxs9pBb9BvoGvVPKuhdt7uBAy/X6E5EWOY7JUnxRyffZF07RNcDDP8isJx+99S
Z+z68AdIl8JcFjwk3IKrIJyoVCpcQnIndF96UG7x/WOS3hlcAZ/p4QmfaE+rN5gXL1eDpeXAWIiz
IQZJftBcE5Uty7RQoKCG18kY1tvkafrmN8uafjTXrnKA9S7YTBt89PI/EadLi2wls4Xie6hvBZyZ
8whR742RB5IJatmwAObTUCyZiVnPI4AgYYMlVV5GXcN/INp/3bmURJIovnNIZO5dJgDjt9DNsQft
/XR6jJQlsl71S2y5rsEox77cUaVqxN8qUD4mGpcDmYWm9bnEPnJ2vXqclp+DTfyTRugSr6plTu0l
ypJHeHbp728zxiEKCcn1wXI3LqC0CDxE9u1MvY+M4u+lOTwf4XsKpal1B4HQSR8Pw0RugjO/QsaX
ofqF1kyOZtsU8yvimXQq24EXdDgZI9JQXEp/qlbQ/LUu0DXxogykMzLVgvTLrpgT018Dtcp5THqa
AypVWg1NRzrpTQCzzg7WCk2B/2SMbb2M+JEQXvFDA8m1L/ZbZ4z/O8Ib8V3NGPNLOE9Pw8NXjRei
LHV24yzVxkOu70oycLoeZUT6C4A4EO0/JRCgFfpsWwug44iEcRAqS18+FIgrK5N0vIDiM/URznfX
SvhHh6gZCE+vuzG0c4ynbyxTrimH4KPHiSRvszhBWx2xRSpWJakCK79ybNrpJJANd0WK8jsb+Ubo
MXdvu6Gzh/XWp/mM89AIvc4NHlHD4kQ00nH6oyvC5GdelaIzn5HgLkurDpox36ZbDc7ZVR2OQ2B5
ZXEm3bt3XG3IgTdgabLNyUUoZRwqlHrgFh9bH55gH83EohMnGzyrUACY8/TJ98nMIR2NJI/fXh9B
VKV+RQXABwC38eGyjDcdRdxiyApLxf/s1lGehzF+pcsTeiQBqhQ2/xNvevcTGiZ2oWNNwLcz75hM
AOXt7SAO2Tgi4mIL3mUB8bZLtbrCiM1DvU3+E/cVoAs9tlOTPzXNj6bv89fz51FY9EyTI5QNbR0m
TJdEEALJFiLOC6D5TUZ5AarfVyCEzQhcsXfzqISWGoJZhb1538X1DQD0Jxfj8DnkjtVB49v7OGFi
3ZgPv3abX2e6LqUUivk2s0dgk8Y8nnUBK3UqBvQQQTczwWT47w57csvOgYBo3m8sBs6uIHYDx7Cc
HV1OS3iyF2FsoId8F/PiWCtD0kr33P5qmKXRKiF2oReOUShapaSvmjwwuMybhFCn7q9V9duvO1G7
ar/iosSucjcgPyw8WABKsOY9Ukrv7sGAXEOe0xzCg/kvFVxifFF9QNj+SWdVyPr8F/s2Q9OtRjhS
BlOYqqObGRYAYBM0nXAi8ig0LOHNjjIezHVsd/PABELoBbGQhHLktu5mfx6MVrWMI7y9HzDCPpoj
NhGeG/DSLu4rr1iAJRINohZn7VdjZQbjIEkCZTduBF2kGi+m6XMHIAP19AazH3a2az8c7SAqY6Ik
yGho+LqZ00M420mW/9CIRCLAyOJuBwmKw6vBhkKbtlKpe5t5kTEk41n5nzDdHJdt9zvhnUC93B0/
tI/Bp813ZQ6MWW07Z9p0xEcHJRTAVE0m7/32Vxtw4z6yA41k6gMQxom5oc5qng56g9SYPhTtuKge
j9ZbmVoUiOBYaEHpPuDud1i5Y3DONyprdZGdb2KoEu3qnCNPeQaiC9aLE6sYhxYspsZA9DFNrhlK
DTTZiJ3xDL6NA4oZNKGe3Cyakqq1xEnSlU0gRHEnNbRafUe/1B2CguEVQlXRKH52IeG2Oj58EKjy
0PQlnnhO7lJFjSpLkbGFyonPmWK5OOPswrNg34tzTmgRFF+7kZzG+tP0V09wCNYACUjsJSctAnof
zpmO7KkKz31bgWgV5grVdL1O5rqF83UAiFKOCXYsLa+/KXgUKHHiy+kQwiIBMhyVUGdO3m+6sQVI
OXb7ve0ZywbCBW9vE1HCZqddZC+Wn6VG03K9VijwBltiOGpdWFgXKSFh8PFKSiCXEtlH1Pe0OhGH
FwjLxoB7wnvsI+1nCiNZg+zdgw4b9RB9qdnO3sGmMs/MYSDjnmOcf9bf5AVRUvZWxIa1D7ZS9D2a
s4hHCv2yZPGsmSgcJWuLweY+UdXaLLfOdk/AOr/s7343i6JjjEcw2jnyckT+RkDTMFkSZbGuCtH4
SBPHgPYAS3XR50x3cxnKppl2zMKvZyrPGVsdkBWSUIIp8NBgq0pNpHhDazcXuNt4eHDxqvAqKw82
cFxP7ZMsyk+5EERY/oRMPgRAgwSgJFil9xR51gKwK20Ii3FnsXM0CC9cYsH23Cglj++AbROfLQdx
gCEc73XlalR2jqcxqseKTQsGSptUFuIMjl2yfJxncJ5/7dWJKIycW01GAsfIMb9HU/xkv1PyjFiJ
f6Ptc74fgTXXAHlnoQ59JBqt0wUDlLVycAuNBMyduXnXQX6sfJ92oOcNDr5ZbHlSzDJhrLgMVsix
C8PkNgFOaTv7p72uoOCK8oL9P7qDONAT2qgB2R5iexd6DDT8uAhIj9l0TLD90A9KtvqfQxiuNN6l
NfaWyb/K+C945jIaiX1p4QmN5DIqeZiDuKY6Y60av7342YHIec6wqxd7uPH+FbzTV8rkZzYiVTya
vTVw5ZbnBN98hJ8zCgXMgzPWMr3UVdtIHuRhXGbwN78MLGRj34Eu0c0WPXfQ9Uv55Lh5qALcv/+6
NRfJ9ztiHzEqX0Z57TZEI7P9O39ja5J5lxmTnOgT+LZoFP1FGuRrsiUn7xfdVal60I3Z3LecXood
yJB2y/ezEOPZmNgs4VTbD7uQxdfr6pyY7KH07+gixSowDOTNjJVpbZJOToeA9SUjGktqYDkwFJpt
5oJJh+HWlqkQRsW2kPTLRVThJKHvF2Lj+wWY1P4HpXgvExiOJs0YchAe/Diy8lzEinqoALVgVx1Z
i5pqkib8NKLhYG+2EkxGBuPTmiCp2rPqC63flkUuhzUsBGGr2pRadbJWUniy8D+Umza8MWQ0POOI
PnDo2ggzaBx1CwNwdyoBmn35m3Fa4YFfpZYuA/JviI3IenMDHgKgRPjZMq5QDSjjB7hIIM476sb0
3P9c/W2VTIO1F37rlHNW4KNA67RIJ300VTvMDQbQKEVJPvLRg9oo6E3EiYlxGzxhfsLuE/2M4EXM
8fMl2V2LbjIZZR6n58k61iMoUBa74bQnBHAuphHcEQQ/fKZ5/apWXMZ3Xsw1RCP0vxTbvDX+MCOw
1f3dvwpWVXmosOzQTtbUCtQ338ryyGwy7jbD1SlUAxcEMbEP54EBZV/8rHlbsZQ2bLyFuUo3R1pY
MA8R/jFm2ryLwwcLWyZxsVzcociivE9Uv6SsA1c+ko74rcd92uSHdZ177WzD3ehEb6FKk8auD79v
6Y6FM4gMp9/dy5mnZsKZFUnwjCAv0uvZDOHoUsVMgjo3oI/4CIDsMugEDvBoY03UsRZnHXQJEC9B
fQ33/VNE2tF6iktLEehOOpa7Sied8IS4XAL8leKYH7p6Vrp5WH8E1H3FdNmbNRV8CTQ9w8aevg/N
4+HAeLbc0zs/nB4DeQY+lf3yWWIv5921cSRcbJpkExzW3VWO+Rm9EEl0BSNRYBd8vec6aEJ606M0
GNmvUyDa7o8atz+X7M4jTQTb55zmqhJmBF4lsK6hM5vcalWZ0ONTziy/Sy5EFq7yECeLuml5c0qA
beddtBUS0IBZMQamHSsHqmfmuvimGtEzHvFFAdRM814om+xaoMLRCiPSI+QDw+Sw464DfDB06666
n7ZsXgVxij9Sz+ehuo6lI03/ajKFMB/YK0emUE3uMgJTFRzeXagQegoLTreFzhVusO1cNMM46NO9
fwnB2fYwoKZ3EndyfhRMtbEm2dRsSl4B1Kro0cVsNLyGhmFEqu8nCLHAFwXWbc3gDEgCcPc/VjKp
av6ZlKyyjt+1XNj3EptIER371tkUiUlhq9bfMRRCA1dG+ajWLahWO9S3qkvbyKs8NhQzFfm2uKeY
fVVtp7KJmEIc/fxQ7Jfrf4wNQLXSS0u85X5khzitJtBq9EQ5As9rkoHvJaqGQVYn6hLkI4+MNfOj
0IREyfOVtJvUQj0coQVlMWHlFFWfzJzq0vMW8tV9bPMBXT+BXBkIwpQiEIGO0lKGC67P4Nqm3WJR
FRbcnUD5amLajTAzE5/H6gmyKIsYT+yPHsW5rFN2vqPm4lIG4SwLqvw58I/xo5qpVDnOo/vdiQFN
5Gwq4llMwSUpehweLzjB/oQR+RePXBEt/yy8oSc3G0yXCNgJKoo5Wj5V5NrkSvJvExaZBicdot6P
Xi07KvPhkiuYvPH6OdXKZZnHqn3YIMiTkWXGLWEHL8bonYdq1NFcxff0P5AAarcizIU/lCw0mmSx
W3AguKd1/QT9/gWoU5xm9X2fw5Z9Ji8v9lipVzKQYM+drTjatsd5IDgZG08R0OYDJsTBw6+fMfvC
8dX9Rq9rtqdVkXqxNr8uQEQNiKc0FRJWH2F/1811/tlfRsxK2+w6+roV39Hzwu/ieU8LvJsc1sUl
Ppmb7aPoagxQXbB0wPUEY2V4X2neYCyWTSOnyWpG3JjLgv5da/10V9wDbh1dN2ZN87JMiVILxNd4
Zi+8l9OfFVLDS1zs9WK2YWKwo3xCwGAZnIu7j0Mxw6Qz+Po90lSQrgwoC57mTPR7Eu3Tgm0Qaxx9
cOwlwTqBh6MRWm50BS2onkQfZ1985U471LYv2xVqsTMQgkTYHWQvwADrYKpkkfIluE9YtC0CAJW5
z7EpgZBFXzzo2AKk5YUzj20PdHDSyFUqOUUG8IKpazOX0AX6af7VsZiaC8MP46thSaIS/cqibbVY
Czz6j/a4GiaCCWmP05SCuTI7vFDhM59SITUrmgK5jBr+qhtjIqOrm5+iWhON+PBk+Z4Nms3DoVBu
bOupdWNbxa1dD5li7W0MRWQFYGxTA1yLTZdRF6H2aeYNtSZzkfbTOe+M5HiKeQD/3xmHCbNvjXBH
2xMJ9scHcxOnOV/S1yRI7w3pVOUbnHJcVOKH8Trd/kByz9SJXr0RXDltbz9i/hCC3zO0c53q+KYl
hqw+Fdh7G2M3cksR3dJqmuhADsaXv1ZecRoZLGVtQw2BCkvtyxXC+0yw9vAp69Wbgn5hQbaRiHYs
Zxka6v4kaaHh6bpVLeMgS/LhfKmId/UgYciWuxl3dI4K/h6w5eGxb5qA8XvLX87/pfF8UdJMyevh
aSBcLkYlsYOi5E9yW3OVaoJTvqDJfN3lKVja4dBsTPJGufcb+107p49Z2+nIHwrald+KH2IxIEqG
J5g6iIYIsj6str8jvzMrvREFnwn2GIKGgaS5iMVnQLBDnbNtAC41Oe6pHsnYsNBKJp1auS5oSrxs
poeRCDXYs/gRfvUH16EGtl8B2GP0weVxsHvlDdpExyYcVOUeg/RC05sbyZKebuzBYaBI08EJxNaD
cu5/cg+BjMGv3jyN69uwtQ/pIBiFeGFGmL8jhApVfrifgN7wyxnyaCaLQbEkl0v7q8+qdKmlY2mT
FXF/TRosXVHQ3bts4UQkUZx95AakAhgjJynj/gJaHIAXITgHp6Mi0NiQSAsDguN6lIuJfLbaE4y9
z8Mc2KuhTzUm+v2eKz6m/ZCEscS1k8F8C4Ocrg+vKMMSptRu0D4XXG9ts8l9/93tyX4afJStkkIz
e8UWiZspBPTmJFtU++lsh8QC2YmmDNx5jcnmv0qY77UTrqIPiov0essktcmmktcB7H6zkMsS46At
i2iiux6bCSPGn2p6Mm4H8CEgEO9W5UvM+JvxN2tp1bEfleEJofkTmTkzJzRW99htf9C0KbuTvQeR
FSnuZ0toYlAWhnlHFTw9JZ4c8QNQGNPTO51bt7aXAcsKHM0kzgdarT9BL4wfNd1cplH9w8Un/n8i
jnxk1pjHORQsjHAwA+yE4gwBziD+K96bSpXauK6vRTk2gzWq61ZJzqZD0n1awrhcgV0UCM8mvD0H
MhO/JzHNbWhxDvd9+zcfdZaioJmSYMsAKJlzM63GrTqgcZT4Scv++C9gxVgTj1WnUA9b6tldIrwN
RtZnjUKhWM/VMwvprFdWrBoDffkgxCg5NCnEhdN21uMaWrAnVSrpZN0qk8NpqCJ/rnT3XVk8WZVz
k1/JUe7uztFIv5IAPSgnhHloSjZzanEm80L3qjffxJ5yBplbZxHZyGOn5rlaAonln1wNQxL6hS0O
0eox6jzJMdVg+Pnk8gKi3x3+NhoeKfRdcR0AeVmAA+AxDDQ+trrr1N/60QoFz70C/6iOMTZyekLd
y5riOTf53t3jFlLbUxX/iMPzVDqokI+4fgp4r6Q5LepWgpj0RdrLx6M/wVNLNjufNjSiOGiU/2kP
qx7Jx5rDUzyH5+fEcSA8PaxwTzWGKBSqD1h1OL0URJzpGPOkAIOBxBOTWR+I751j354p9UW+e+Yf
yOttt+0i4e7S43r5LzA8JU7RKI8+vkvWmwpZ/j9F27HIuElCzdEg/6nNTsIdoJGGu7seTOFnC0c7
rywj1Q1JOMc8WXqSTuqsNet82HxlMDppeGhxB51w8CQFg0Zo9i3kYcYthg+wMEl4D1AuMnRyNm3Q
voX5F2DBsK8M5qRseP5xEZxtxtTB2XU+B4opd+s6SZQdOWNyl8i9no/b4vFMQ1He2O8zWnSLoFY1
HzJcmL2WiPXlMU8eJmPApiOduWSWdp/0M0xLo9unFKNoaE0/jMNDmzIDCGkvkwbdFNtX1EVaIli/
Y7/wi0gMjCsf4kej3VBFnGvQ4wJHqrJY+IbgqWYUojhMFzEw5iHd8cJ4fqc8Cnm1IHdbq02q6f4T
AKdQhtLf7KrXJHcmkXGiUsOgnWB3+XpAB2Mmq+RQaYMgM8t4BIsc1bv1jjnMnAnKg6TS2e7syeyX
fiyUvsmCBarRg7ApeRoNSl7xlO2Ksjoh0Q75A4uIifmYFvLvSGOB3i8nWXXHbTc2D4YE6+xmFknq
eFx5nbUNLcluGxkXDRrDgYqgAowIT+D4/edSTWvGXNR6JlpM05VoO3W2u0EIGwSXDSRz3hc23fTj
RGiQOolWdsQQJdjRcLnLoU8A9oTBAgC6ALsMOU7qO9jUC39vL08FXteQzZfKEABUl2XIhdwnWk6O
qGKbR+RAyRWzvBT10NqWV5a6p2OBFKUBY0XCt01EcZgWuW2nmvbVIPd2X+cnihSH7d20gwZmkIFe
v3BMD5vf4hc9SSLfaJMJ3kcyXno0Bqzgfoz9HjHniJtL/4veD0T3nJK39/N2oPI3+q9QFZyPWZEX
Q7BKM6wL0WToiHdOXj+rtfpbDDho6IgUNKCKfx66XHt+e9nyfZEnZHOEjQlEQjfS1TUfI0XCN514
LkZYD9aU800uaqwtuv84MDM7h3ZR9iyPhyokcEVKhzfwn3vM+EckzwxZ+0HS0fXFeT4vedlSOhlo
c8PUwZdm4IjW2sDN8Vdh1/+WkIDB7HCZpSfnymy7XMMDVSPIWXNpkc46IUeWAAty80cYJgMeTLWw
wh7El7BPFC2t4ahBIV6wXOZyMAIbrPR8bCulLeGMn2QRm0494PEfjHBwT2BKczY9lal434uWvIxj
XjfK/jjMSkCmA5taknntYkCu+CNtNLd0JbpEOdLTEFCtr0FtNy3EvMS7pOKwn3e7rQ9C5HLng/M+
YRxuOjnGiF5x/upGD6tnwTlNOxQ04tqJJKzTezl3G/4H8XOrklICZC8fkaC9kesE/fUs1YhP87Or
7PbCf4xC/BxQAd/7RhlCrxkCRQ/6SkH+9JDlKh7opup+0PCcfz3SDLaw7ga9k3CDGfMDAXSg4hYm
QItfgdRcei5TepvPfw2XRtd8TMoq8FChzqZd5Dsub0tfk5FgaSyFXIXKlC40QckRi621u1pRiPxK
LT1ncO48OKdBMaJJG/WWEgZfoNYyJqDTpTrz6VMvo1JehSc1IgN4OMDiWPe3YAvf1hQcf57oYkh5
MSmiSBKnKRA8pdQJ3GLVQZVCoDHJT2h2i5zs7guLEYO39aaT3309qRZKQw/fwReDRaDjtXmzwHn6
eEcN0dPClPUAk4A0ok34pPsBMFbNfL+uS9z4fWFy1e+Jp6i/7gGHRrWl8XtrddLkMwak5lciXD5Q
tC5KJHEiysiMyjeL5HzP+vq7HXITTLu2zS+QSnsh1b3BOnpju+L55tE8vv8+F6bfI80p1h67XFOc
RU4KaXbhIbJxcmhPrcqJZN8Q8IOIUaJEUgm0bq5WYibeEK5EJ77K4Tzlk/FcfJ1MRoNvSfDI2u5C
hmgMrJuZiGgSRIlx7NaMqU1cINFl8SmqjStymYEnlAU2LFEOmRZrUCIJ/ZSvYhGIl/9nVmgKmVfE
keZEOIg+t67HF1BZyLKfIdz/9bPGm/jjg8loal/ezfV1RZJ7WTZoJ2+REu6ujjoNTzX7v46AiytX
quOYdpP2Ak4LcwxAYtzG4AlqcOW0gur6YsNhAhLxg9HbwsvoJh3ErBzJOgewaPv9KpZHkE2eSjiO
iJbLVaxVxq4UVdKACIVSthwCoNZJECdKaVDbZ3bJPLZrOZA+Lx3skuG7cfnH0C1hRKWN6tBGxBme
4a8OFeddnshj6Zw+1vIpvC92soPNqWpwdaI11T7LFgNv1K88Yu8Aha3ihDp1S9cfqNnlp7Lq0mR8
/4UGQYH0Winl5rYaGm4RV/F7tpNpWdPXkO88uzYjnMeScQpz1RdbdCnsEA+7fkHshYOKvW4TvyrL
e8E7SwxRAFZx8TxREa3rKd2/2lhcA3i+QxrXFIxM4nh85eFvFBt72uYMeKGzUedeRNcQBILiA66c
WUUKolVQ+NflEB99W76FYJxAom0dmxZ29v/SHVtF+Ww2AnZhtT4hlCPBwpklH5DrGhl/tkSvlisf
MpSJeAK1lC0R7SjYmz/QyVXQn/uJwJOfS4Id8vYFRAi5Lp40tFhnQ5HnwizNSUgtryxfP0mxJcw6
Wf+eOy5sThpilSoUhUG8Vo6l+0LG5Jp4pS5vDxzUI6iALKZOIm+3S92sCa5efEmxYR7s18+E1BQc
2jzzzQrk1LjUZK+Ai9ErKWlvPb4cGO5S6Z98OwdWVWU+zWAQhbckqxzey68Arh0+zkczZOwLFHM8
RvBwnOlT9pjNQZovGcsPOtBZw8jqwLmflaSNaxcreyZmv6pIfczk7TxmWmbm69uiQvzJq7CP990Y
igWLFY4DbzZ7agb0S4ckp5H9Q5c7JLZAj09J5q1YOu1gBg96y0Z1i4ZquobvcYZ6Oqjbbv/CeANw
pvr091omuAgZRmyPmiFWyF4j9LsYpdCAcXXSaGcFytru50+I9z33pvHU6Ijg4dmAj5VI7E3eyuqU
QmjCh5kH6QI/u8yAMRTLKsLDT1Hb6ReWP2Uc6ybmiMfpqOn/cn5OKVW044jBVndESbeGj7n2Nzss
51sREVUTw0yoOhmzq1Rm/OrBGWvUr1ss7ThGe1ZFiNXBezurTnz8dvYUiZ8bmLB3Y0p0XPrSuAQ+
ei0n3OPY9TrGi1VVaV01dv/B00pdDXbuUUAfRaRP4/TwVNEp1XvnT3Xl3/V11GKH8SkDRc0Rxu2z
WAd6Px9kT1HduLaN7gXbqebu/X+eHA6WzY1P84I6xWH2nvpbBeUGyE+Q13gbfJiovkOyjK6CHjzr
mt0mav5pGD3JPZRppQ9N0VMvGQeE24n8uB8pxYEjmp5r0Dd2Eg7MvXN6fkQBvUjJsxtps+IER+zZ
9pqIVVYonY50Hc+1WBi2fRnhUQi9oWJ40bMmCEgaAqGHW7wezx4He+ppJqmwbbCV5FPj6vgzr0hU
WsKzZo2xxTvQ3bKA4O8dyATom3G1+S29xxjMot6SFo2lKqMowAT523pz2j6vu06CQP1r3PmgWpQz
gFmjem+XLa0I0ZvIPGRof6a3sa6C+1QlCRfAiG73KLukzDC/qnaCznC2PRbLFyhLsA6BzRcwMD6b
JmznaNkxPBVcCwBbI7jIK4dsiGNrB1e5Jr+veCQXZxM+Qv9j112USmjeLiO53D40r4XqQfs+Q82F
vUY8C0bpOYVoL5MTXIZ3NgY3tDe6zI4IAEaLr68pmfPV47SQnMxeFvxb0AV2EeSw+MjVojTJ7MCE
FaD5y/es6CxOUinbhVpjWgcvtQbk7aLsmaPhEh78UpB7s7OJ0Z8qx1RKIfKckHgYN51llpF2I8NH
4Unq0r9DyvlMKHklLEXL/RbBPD3H5B6Hv7iWr4NHwOgjhxFYugfhFEDIg4l2L17e7WVIbRFZkXO3
gO9NIjkrmnu+qwqAXaTmWVDbzpHySkhkzfdDOjWTuApE7AtyiZWmA+x3DNEfc6fVAIvP1YqJoDqK
sUCEgG2lA7b55QZQTIZd9sWpwh+yUnaw4ZQlOLB3dLsJzBIkL2MnQY/MUlXe1R6De5HIQ6mSRtgL
l+jbp4I/Ard0U15/nM4IPBXcnArrvihnb1UsjrNsVNn1WoC9qbmZKCEUE3OdHikZTDpxJnZ1C4UL
yjc/Qj3L09X07Fx5p8INhPPnDNIAyAJ9Z/ZeOxJ02cZqBxigwC+YwOQRejU2v9rl4kireuOFUxa1
1ExvcaoZf6GqUqzOW8mobiIg2T3VE/2c41ne/SBC5b/81RdNPJysZMiQhABWTxwHK3w91ngJWHN9
ay54B6HSRhlTAtTXt0CLnJ3rW5w64XkJW6yl9liRuF2xFYu4BY1P6kIsg3Od4cpfV9i94Z4FJlTX
Lz8SJdxuJ6txE6p80I/J6sH4wRCPT4EI7uK8oW4UEP4j0a7ZVNWLOPDLuXhYsIIYAyeiQJTGmhTO
y0lEiKsX7jxO02HyM7+Veqsuw/um+j2as88XhUvknpAYH3MOl2fKubGzCmY78XuR+lsYmQSJ/sF/
rSYEgjWKiJQhfUjRSSpud/j72+SMDLtuveb/ATyYOe72u5zqrjNLkNWGr9Fz5I5F/pfIt+TQunOI
SNC85jYYzKgFsLP6UFxZJnMbUybQWHo17P7YYda18Zq6o1sN25J9H4Sxb+OfvHbVHTIrm0HSnweU
8237APNgVPG1nMerR5UT8YVHj0TSzjDsbW+h5KFFdqZ+GsT7nkLjRX/W869cwarMHuhkxRM7CkCG
gVWJ8zkRgHHlooNgiSsNOWN2GS3n6jl+uHEGTfZr7bT9yCgrmYarJZuurqfXmrFvSP/nEIBEY5VI
aS8VeGxSH/0QDJASupEmKGRsfmAQD/dmsV15xzK6//qxJOBIAO1zINHay7a5/HbP2gewLCL1gJKt
mkfaPU/wN0uLXuKLij2bqe1affNdtIzgcHCi3FVth8AMFmxf4MR7LmicizTQ5RTYPkJPiAx8JpSK
9yITQe+tB5dKriAcflJNwkJ7r/auLE+gfWbDyKWNLwDma4ZOM8n82pGKsfE8WmxuGRR3gWmCNUQ1
yVRDwneHxFAMvUyrkZ43wNT1tT3Gdbf38G//NnFAmSJ1XmWJXPDgWNBdtqPfxLghO0nwp9pEQaiD
haururOaOFWitwhaoJxh73LgYGTbFimnxsRkeMH2oiuYjSsfDvYS90HhEMroO/XnYXzSL5YK3w0Y
RqpmvOw43tZ/Ao9wlH8R9TcwSEnhO/v8sHAAoBxJFjjOPPYJVKnSGzgI03/Ruq7+rQSkrWvALTw3
Bo4nkH9QDSSIav6GBDIY1RDUfVN+DC2mX2QEIom8c+HK7IKR2uBA2IOPUQgjGTef74hgYdFA+HLr
qGNJYJXHIToj1yOp+4qNdMDVbMhUbqj7NnsNzaeyLoPgjzSnGMRrshtc07A3oRqS5A0kcFe1o/3w
V2IdLc0Gi6UM6b+EVN978oDGOuhLpm+RHpB6dTWyxmniUvwk4wxqtuOIzkXM9DQYoubdjw8A3kS6
53loE7qMsSaizW4sXrAAARuFRvChYBbATvZaVq8JOb9d3tT+yzJG3KjWRu8THIMdi7bmRJiK8ApI
NJJC0ZUtbNv+y8N3+Kq9x8lFcqPWwVPQCHzLOD+JlnVhFM6dQShKhiEsrI80ojW5pc4V5u6GQ1TG
xXcyNPUcsCn1wIZAACrLl0YfPp2Pzfg5OcXLsoJzD4JsZVVmnxJy4cTyjRsU5lwD6K5ulHbb6ntc
RRW+bFSutFlPDM0Vik7vXBNmxpBdbSrzgqiVqb8DkjF1uflMMkmVrE+1aH0rf8gDOqRIhmiBgsj0
kdtmLR9xRKYupgEaRCQ4BvacK7y0l4YVFLxYlN5vej580uQ17WJbSMfQuqICsS2ImHS25524fiGe
gSAwj18otdtjXDW79pFh0kzNbBqUUEX9PKiNRZpcCCGD/VlQ48D7y/gEWg5Uuk4zdOOlwV8gafVT
v4HjBw97UdkICEoigY45ThvCbD3lp4zp2lvF4WDnmbAo6wIRNotQW45ClplPnw1nYGHgoHlEzgOx
o6Q4ObX3e5PvT6vw5Mi+JL29riHT198FkOlX8aFoEo2BndvbslXyzr7KBoMw5zIv+D6zzScI3TeK
Q1/dRqpVnwEOq7Uj6+2Af3QhcLMBkwF2b+RSSc3Xbgbl7S5c/HlJFWbGoRwRBu0AGxRoTRhvyMGP
sFGr12WY/0Hx97bjEzn20CM6ybDethKCItrzzHDDmEa6rTmoeBNfLgpwhwRfhgX7WJ/udOpa5IIn
gn6C21AwR7telicSFWv66wx6NqzChygKpp6lgC3xes8fs1vS/iQeF0ZHXOF9MFAF9p8ovOKf0Hpa
0QN3sKoK+WW9kauvaQLTU6Dd1vR7UbqxX/E2wuWQ5XvUKnSF+pQGafOGljZ9ZTIBgUvMuDWpCG+F
NZ6/UAVh19wm2a5CGGlBmW/UDGOIWRPu4vg5s+OJbifSccw5Q+ohZeDEhbt6FMe5Fo+TCkWKDcvC
tC61UFLO/w5mR6BURhJdtmpNnuO1XQ6DXkGRTBQXVZ21nloObTkKDJ9d1drlfMvVTX6znS00OXSj
9PNsu52WlTr2cten5hqzH9Dk9roQXMDrfEizxwkwmZaBhwmwisWnIYqvIBtxhfydwqZk/YLYgvLU
LxqNb68zy69et2ALuGUMfQln7g2Kp6bO88SNjCeT3cYQOXt3ZwF8us8FKQZMJJcprQG0RvUjwb2I
fFQ8+JNuIpCqGfYk9ce2CJWSqbE7Vy0HyQ3o0AVTlxrBsixcqPZdJ70+xv6fIJJuNqZqFPeQE54i
E5cQoctY33tVXpVDthuJuLPWct5SLxKunlAX8wBxRqtlO4az1hqGdE1jkfrBmb0LRSg3uhJnvFon
y2ZCGLkc2EGDatLPvafsz0eqV9drzYJeItDaS44kAhkwM9vlpJkhc0tab304KDHRZaUBlwRWSY/U
2eSPYrUEG1E+c7+SQxaeU5vBapN0CbIilhIr5KDOaB5na11Dq7doPQq65mvWsFOtBW3FWJiNcdDG
DL/h4hV0EGmhiqRSgo8Bmq/U4GfbNIMzPvmqGJqhP0A12H4XJAwH4hu4MlQhUC4eAMFwue1IS6pG
CZhb31q7KkWLRfxsbNrsJjdhhE5Osc7kwXxPB2l2yU1uy9n9JaZgiyZuh/khACKn/9aGp3QHeqe8
+bT3Xqak+kGwjMje4TYD/n2UywyM43CFRvRyywdjIMiEOaNFKZM0m8qiCaq1/fHLW7JX2QQrLM5A
2Mw+xhkVZdLgyPHqD11dXOMHpI8xz5Sl2KCBwkQ7r4enea0mKZGS322JDYg3aGO5Sf56uv62TPbU
AXqhtTPR4cO90ryN8y8Ejkp/70ePlPfJV4mJ3V07JaJ0xh09XhBBszj609LpvETJKEgXRe9ktTeY
v+B3C7dLdRxb4ZTcFdQmIG9WthOPV2AyUFpzd/20IvUiJbkmr8Tvisq0uqYwL9gEIzd7FVcBwdHd
HePWSOIAkx2rwFbQ0127NV04jPjtdvAYX6PYRXKBbl05ywLrtXDEUV4GxGWL5bvzvknnvRH+3ag5
5wPa3+h2Rf9NjRSRTDahWqAwIDafW/v9isbX427d1zQVp4/vmqs1PqHun9MTab/3nwwFnAMgjtCa
2JKciXkF1zZTZMPcJQwLWPAUnbltw7Qfd4VyzmI4aKV3aFM/+kjWfKMVs71JDdSjyY7ZktY/BIOn
Z3ajSLKt/s9KQxr5mN2s4o9ZAeFRaiu9dt8hXnVtTwc+/+5yYA7+07CZG2L3RbYuJWhA5iyVieZb
A+tQqnKsO8Xje4tijceL7s3ZSd601LRivPs/Qwdnufx9H4XTe0rac0B6TtvNgpZpx6N6c+mzvIew
7ZGxL7iQSNBKNJ7W+lEDwDbWllKCAvjpjLLiKt5qYOI6ZEMUNQNyKMlzVx9LLgkl+SQV50/XEXhx
698Wy+j3WMedkMPLlUsnN2lZYiHYIA4jBjQF+4+DZBIIM5gPtthbTScwzC63wZj2s82MIssRz4qF
UHCzpyL33pZ+pGr5MLluPJd1t1SjfKIfiib7kpBHPz6nAfOELoYavx0tmRzkkS0pkjebwVU0jnYr
ZVWnIPFw6bpjiUEezbAbLVwbQn81WXAbW6Sqp9IfE3vsXxTuara4igcECAM23fVcUljitLEMfYdy
WfaSFe/UJwJgya8PIFhWoBAFekAXRpJg2R6V6m91cJX0gIBfdOdWUDMejUHGFCHAtVS7yfv7xs2G
QvwCKMUyvdVwlSWnorXBcj1JnMHmhBo5GR8ypOTRDYrcera02xy+7f26DtuNE1ygbSSbBom9hX4x
KMbUmuD1MNv+xJkxeNZM+j4xb54qupsoXfBwJXefb+n2eEViB8fPQQnCdyQPLm9rtpOrrPAvV4WP
rQ7fm9ghR/x+ZzLiNDt9NfA2idW7aLj8UgRmhLrnI1Q/GEMzeymGLis0l5oi3MTbCmEiCakHa+g1
sma/G8Ofa7x6ubUbtuMELioWYwzcdOxXuJUCcz6uNQ2853z/FA6hoqrGLrtHq7Tlx3eDrHQTqcIm
XtmV+67lJPPcQWYN3IuH2vn9NwOheBaXemnqk7RFsfZTz2cvqDOOiMZW+wp2FYbOFf88NWUL7Ztp
jWgUt10iIjTuzMW4mGcCIuNMgFPGrhpUPeK4e89QjP+GejQfQqLdYzLlvPcl2sZEC68z/MpbG0zM
7xj2QXGc0QYi+Fq6F3+EuB+FgxwQx3ZPgH87tSEwLX9D7ReNnnh+q5Dz5F1lf2Tc52KSY5ASWB83
nJbnt3+T4ZjbGk8QbEV9w3CPolLUoSrEQyb7/jzd7ZVlGv5KWG+E8jtWz1UieyhA/hEzhVL1a0a/
zJdX1P6TBYXAG4xHw4Ga0KNh269/u2Zuopj/zqIkBZABz4c93f6zPe8f7NadmHF4EKia/Zo58ohr
mQr/RiSS94EvNu0b4U5r08M7UmGsAvQG5rklHJ678TnTXHCNqVXyNPm+IkAiyYN1YHvZWQc6gKqI
Js01WQZ4WaNlulF/V3bsKtEgkWG8qgsTYJ+J9f1lXvlMSNtnBXUr2hGpOEZPHDyRip4eblvuW81F
0kWOyL3oEsH3/Ra+PI5s+erc1MxIIxYAlOJob+y1jS57w1JEMXS9JgnlOU9fClVJ1O4frL5gxaKy
pnkyRx7cf9AnX2wDK1san1LxQFCdfva7u6OIbNHlAZUqjl4B5sNCf5278Y8MvMS/2zjKn+cSs9Sy
WBIegfQ0DkLQVgvypMC1BqL4xhghFNLHVDFT+sqBKVykofgYyt2FjFIezzLiLA311cfhrw8JSO9p
uCVyousUpKd86WrowwNIJ81weUuGTc+BFR//TRO+WCLqpBhkIllK/yUzJpQVe9UuH98GX/rGMKU9
BkYkgDNR/ZSFGNPYiG8bppaJRxyt2QFuI29QvYCs3VeREjcPKK5aAtoF9nanCe/rHvXXYbvs5iFp
GqGVgzBr4RQ2D7/vyCQAU63cux684+Ur8GRJ1bJcPGOgmPnkj5KWRKYXvPKSAJV0/DFSU+0YbizB
+MfZQGWgEYXn1qCWQloxn7nODgE9C+g5cNfAw+ivoIKzFQDS46U7WU7DXIQq9Vmpv9E4qDqfHuwD
GJIcSU8ycdFnH91zYXPlVjyXVQc6NR5Tll1pbEC5MwQ7TWeV2qn3oaQ8zhEtq7FbLKQV7xxFIL/X
SxWdydduvT9oB631LXRuJqw6tIS0c9kXxb5HahX8Fqi8w6/FexbuusamAIYP5l1zz9SFcpQZwdhQ
SyBvATec+shfUj80Mjk95Bwpjw7QaTDvOtJ9qLxnwxC4bCUtjyBV8VkFtdE2ty5namGIzau1Z0h/
5GoVQ0ObgWJb6PW2Uvxz30DHkd9me10Ps3uZRetc4CYVf7nixwq2f3YohOzm3I0j48tFn9fHNaos
FDD12vk5hvhZQIhzQOkMQ0SQNQqJ/5Kjioh3xpHgOzxBvP78GoTY9gtEf1Nxp+RWW6lun3WthkY4
7Eo5tLkojEY/OGjrbbu6GPJQCdGyd3I6ZePOh4+8Gj8+pHrn93Qd/cZL0Q0PyDZLjgXF0dLm8y64
uAMWRlOPl3/asI+MNy+OB2CVgSx8kI7RC+v84G2/Hq6IlLJ2Bx/HQKzBAAwVzALWYVtFFm+GeFRG
QHU0lObiytAJjHnE9VRi34GgLd3OlArWgCoDolsnK0F+Iyk21dFDtmEu8Qnm2aMrhlvu46SIH8bZ
0FMOa1xL6AeBSYjkMQ8vyMfHO595BnAitsJd1OdRkIGvxJQLSGr7SLbHyr+UFSNYs500eN5vttys
237OevqjlxtvTb/5MPYvnx55opNCEA65DCupyfGyx2UDYAahwEbFsI1YOZo1Bdf65pDHgdXEoiJJ
UAqk40mbI7mvlypOUN9kasjtBNU1ZTum6GHKSU/NCxoBgkg5/V2siBURr5omj0SwI5uZEfqvj0UV
OGmVbRv3nksff50wLzR+BTKag5FWLXSYhLC3yhxaUeVaSq+VHupIyMEWbdKchn4c9xkZt2ke/W1P
jmOobLkJs+wW6mDGTvfG0tMiyGYSzmtUhmbqbY/abdwt8fGzibu4Pli/07/EtJbg1qedYSOd5dg8
cr2OJaRokUD3815Ck9wg3GfjcjvqkSLmeC0etRvFUcUYi9DVhlgl6/lLxVqJKW2w4JN/ByfYLtmh
NY3Oqy2lGbhb7oO23WE4ntLa1zJ+8lM2ydcKGFbZexSjvQcVc1x2nooA50BaSDBP+8+af/bD817b
BTH4E6Rlw9Bad1eYqDrJkHlt1efxv/HDSt36MlpEOQu31KUVQ63oUDVYADdchJz874JWtsTq/py6
gT4s0a/G2Ic2yZIWsNFnrUGbcdnfGjankU1H8Lo0IPjgYzBXLe5k7by9uAVFtdZ+ura+XenYsdwY
MCt4ojp0y+b5+4zRsJIVZnwACcLiJ6AFzn7Z8804wjS4krgrPxysAnHTAB548AnRSHIHAp1pRSuE
GFY0cyf+vZkfN559QsSitvMhk4Kt8x50eDjoafcaGM389lyZ9idVnGXnAdd81jleLnEat96i+rnq
ZaaC0o5uEB4jAp5p7T1O5L75HX3Rzt7P6USdJCS3YXPcryi1CiwFueB+IcCOmcdyTqL7Ku89V4AG
EAMlueximW1ldWluGXKlCP8Im/ZS+Hw5yqN3cDAiDOeqtsPgnA8yvEkXdTGp6yAonEOlnSkooqqP
ksjnAWt37NXh7ZcyKvKR2Lnn0OtLvA/IBrdJLwzkNngEyWG1tzMP/3JmcHbLD6WQme44RmThJEhJ
cstfHIT5+hFnnDq6Rl+dxzl8pNeHl/+ZwhizV7guFb8o0pjk9CPC6iV1yMSxtP8bT/3rgBYSXwAN
odjowlftpCLtzb0k18Iu8HMzaVgqQpZROs6xpcyrbbzs152jXDVz5JGxBqXTd3vSog6iEuPZ1450
qJkjTKlMqsLUSX3WV4GNsgrvZ93FkG1if9CPwBCv9iVmMs9Bto1AlQNVN6M8tSiLhl6boaCBeJH1
YRohM3Fl8xjCZk+QuxfVNxdrEP/T/hPpuIHOW3dgHBLI4AJEoTdY0h5sWK+3sU1uI/VmqmdDjXWy
06EqZ9C8l4ehTLyo7uCYWpg652y1c/PBxpA8KFMSuAAXo8H7EYtsKQtYppS8AkzBdVaGf1Zx2H3S
Amcc37J0YabFGrd2+khusu364XO5X5WJNO+p6ko5HpqTJwAwAFCeckO65nb8mMKHjQUCl479nf3g
qJl96o3/P8+0oD2MI17GJmTf9YRsdN0a7452vjqoNTcs7rgG3pRqMGrMQlVqoLEiUGe292XnGPoV
fgY29cgg4CSIIefnAjbrTb77Kce2zFuE7I1BmYfQTbJyACoEjJiVl2GeAm7Qn2/iGsGVZg/1jfX/
Ay6XbQI9sPFO/bHRY9MOzvoKP0EuhyCioho8KX4C0r551KuiKVq16T0N+aXnYI92BPGb+DRWM/aW
SAQLwW4rLJDkCmh/rneHhZh0odX35KkHPuo2hEaCI6u3GNCdz6RHr+QbqKkKDQthCVi3WNXW8yzr
uZxu/wojpoK37Psszjq78wBb6I9vz3xHruPMwdGlOia0Lt4BhkvJPTlj9BIkTZb3rnaAyrofrScp
PZ7Ra0rU26YxsTVMWSQ2hd+IFL/qGBT16NBQlrquLHtJ1DLJSFxNQWIRsYeRkRCh2JGo3qtsLwOS
eMWmFH7q7XackbnnwNeE2/AQsl1Hwod5aDWFPaSj3wpNi7vYLpAknCAw6bVBgWgYwf3oTnGWl1JX
dYtGVL/IJWIx3z1d/yQ+nwdeJulhQ4mp2p22t8BKVDTBKKOGYSeANfNWm/veGZwhvRbsBMphe4bD
/hy0yr3W8hSBNG5S4R+3N80gfG9klys6ixECLnbyNxtFcrBhHiiwBpZnhGyoooJLj773z7jCrrJ6
XTdHLx8/4mNbpAdeRqP9S3hB5dHJH9Y+pw5ln79BSPNKV+iqz35cmjl9+Uo55V6dH45FH+XcLDnd
aFFpDxVwatlrlkTad8Ymg/po+EdoV5B63pZ0W9HbT0mBzQyTI9K6XKsJn7nxeKhPQq99vtIf7FlN
MI9PP3brFN3ftB7oh/VqKK67HfnJtkVIrZ4UeiQHOWIjix9b+CK1WuVB+d4rjINkQpKIg0Mp/4Je
3fSLsDQwDjbfFsWn70r8nqSwQBvJqE/MTR31VYdNmjCSBkYT43zZFeJ0cn4MeOdYyyk9lGjV840Q
Zaft1J815wmg97+1PEMTquNAds0sr+zRQOymmm6wzY3xuoScoyF/kZeqSuqdH7ewkvCg0qKJIFyG
o09DFOGqUs8nmtHP/lDvp1LoY81IhsOwYGK3u70ZFU1oYDlC99QFyqTfbg+x16IAEigPHE5Cl5Pd
7RuwUW430u8QNB/T8i9N6u8WOw6I0I/+6LDehDfi/acGMe8WTyF8Fh2if+b5H4R7Ozqpmwqdqa8/
hPvkh0+aMrGbis2m/BJO8n0VSjPcaoRHc3A24uhmjJe33jMJrsqTPiFlpTn/lzZ/q+4Xj4X8sxYN
wQbTtLWRa0W2shOVzs/EhJFrGeeHroK83gJJrDn1pSacCbDxv7oBI8bX5s0xCRSJywY14o+YvNzs
323WnCgHjkn8SRnVM68F2rtY9Mfe2oNNrDZnmtR5ub8XwZcjLHkqku4POOSQfMzk7yF9IOzYeBID
nXkaOZTQYSjfxAHnHpXPDaDmF23Zs0WV1QD8qzhTZyMPsiMtBGRVzZloo9ZYd7h6vlkd/IqGRHNq
wzrPMAlF4A9aysbTxVq6rfiHI6rzghSKdisWea/8T7YIf4/4zYsMO40GKbuebYm7k5Qp/02zaE3W
iV3EHZTVUitRR7VxP5SBg4NxLEXGQhswdJaElw7S7x37m0bYQufP+BCinOFecdlmA7MBKWDTdDaM
Wrd5kJZwTVk0buL1yDF5MkQ7sDGWV6EmkeFTzXWBzMNYe6ZcJU+yBTGmLXTgaefUifzPHUvP7o/U
IqHg4UaqWce76+S7gDi+kA4p3G5fxETkivVnWSKrtj3FhrfLVs6tU1VhabOwz3NClEb51Emg+PoX
qQ3JXVkh2V574cfMq9beBIrzgX3bEByBpo8jvGDOICZ+cwohq/HEeLVRTjxBxeRGuitXBWN1kbc1
UZxbhUlURxAuQabPPD1aYGTGYGiyy1CYFHSSGp4IHlW7RrKDWqTjS4nEBnDo3431swxeLBeIUsvE
98e5h2y5mVSmzfCaP77t4a4LeG8QbGsbHyRDsvr1Wepc8N2WvjMGDOCLT4hkYL5MgvzSO+zFrP+D
qXgL+CEZYDHT3kYVDRLe7v8FlGK5vzX9A9+E7nEOB/RC5qNed8CDQiqzS02WOmzr0Yp9tUZOVfC+
LktptNACXccynCeb8ktubwHh9l+rqKPZs5ins06JnepP2RduuoVMtmkSnvZUhdU+mz2cPDnmogA5
cwqP7/ktFJdlwsdnK2tn70+m+YoeNfn0LLiknG7mK7ijA//Vpcv+MwlfzcV8xNyrLHVVurYjxWqJ
Z5LRqUD899lEhijP6NMVCUWVdRZxhRzfMBptT39mu5yXMVa9SvcdvVdFyV5+rapakHSi7ITBpc5s
fsMT6o13tuSAkU3ylAxmxWGJ1MRrhbY+UYlYiiIGjy6hFnrVBv9lq9Xi3v4ofw0xxKVqJwyFy8D0
EqtlktACjpv721shhxuvk29e0D3hJad0a+X9VFqfIplvl2ce9iwinW3xV/OLGnJfSRt92wdBVfwO
JFZMWJ2z4lNf7VNGQQi91MhvpdqJvOsNENiovdCiRocUhD3Vb+ssvtpGdfLD3c9Yq9ZCFmFa/cR0
mqO8t/pDYYr/MMdT6lKgetuyXDSOdJDca/TiNFtxtXjHKApaOIbeGL8MmEylZLWRxmSvipyA++cD
pCfNZ+pPancs9bONbOzLxl0FJno2TOA8UphWK+iE3AElOHl/lzD8JQ6IKXC+s+OCc6B+U5d4IlTQ
mnGSW2UAF6BgPAU/fze4vGDBJiMrBhz7fGDfjcM5GFAeXaNqFhCafI2y1P7UVVAhoRLytRdcG12u
hEiJhkqAHeJkF5jCu0NrdCUMBYprRgX+WN4sDlAFtWvN6ZnyJsDWy3RuSo8dYLPdlLsfAs4JshQk
Lua2qdzQJeolrQXl6SQRrN4ToirV2JTZkmoHMXv7cC65Ub5KeNuAMkiVzc2zWSU0WGfHT+6TjOaE
ASx7ofZay52FWpfFfqZ2xfP7Mcuhva4VKS5UMTggrsPyzhCIJmw+UgQsN87u4AJUiIbb9igijHJb
Ev9myyk5PHeMhBysE+b6xyWS6WQBxqufdqXztMX5mKsaFonORvWNswZYjFEE8C9xBv4SOGU27uF+
+9NxP4G4k7NER6Yg/7MdgQryMIXmHJb9Ni8ljoVPodXmVU0sefCOAoDciWT9YswYYlqX+pkwGYI5
yiwRDNT682A53+dU9pm9q0Oe5g3mB2TbkXsYewFAf9jkRmvvLgLO9ii0zFutbntJu3CKcMmzA2qd
rSuFeVyg+5GYN3Mnb8d3kmcxph6dS+ZHjoW05OthQWS0gYfC6fZzciewsQsMJx7HPh06fXim3Swb
3bfzGuMF1b2+A7BvqKGVjHd0vYnKEB0ZXYoDoZ4Y1uazR2NiiIU0hQt9ndZVWMDQ6NANjFTR9HeJ
qsCzWvgTNpDMdjYvZJLgO5Td9dv3QbyddErENF5HGrA1O1viha7p0kq5HJRv1EdpyBypiLjgZJFN
W2fHcpuO8NT+wZi3upH6KYXysnPqfVjunJ25gzlk3xKKxSNIlmWfB76R/g8n6bRCGGu5K/UeRLrh
XcBPIqavBNammu3dVTmbdNmYWDvEFnsSvc2gsbFPsXdzLq78G0vpMysfzSxwJd/QEVO9DTQ75naH
Mxw1jwqjq3JDDhQEsf48of6m7v1bky6UXARiOJIcx/IvyVDR3v8T0MDDGdpzZVUix3AOQ8G/TJ3k
WziIh+ROWk9JpFlsau+h3NwkhIa/FW8nCBc6tU3DP+Yl6hck0UrbTUsIGE+UgIPQ8tWiuqVtQRHX
5MjW0e6kJoXTMGzHVUkMR9IhCRhl77BQV3oYilPAOY6ewJaigzRNeQ+hudienpJ4v6ux6YFJytDq
w7Yjb7+yyg+5A2lRsT/+R4C2CFm1Y27I2BqHewZH2UBVC0spjCIiGq8sULHQIR5py3l5Ciama1eI
L9A8sYJzNb0PJonsKXE3KoudF3Zilc6UNBgoCTzhiLhrcBQy0mTXVG1AuPOPFugSpH1X2RuAvxcF
nhbNKAD+Gzu55A5eeeu60NH+NsMRL8Azow6lk3UaKfmvqkI22DTVpGOq+zl9gLHXGOFO7Hkg4iHE
adqYiZoFhZF1BAPGKsoMSjwNaEGefLGqa3/6TOgr2KqVPT0r7WsLSXMD9eMa8eY8VnnUrUOl3ocy
PlBiTCcnyvI/2JbQ4RxYHenecC5/m4Rzd6Kqaosdb6eUNne+WY1n0fV4fBGXGTfJfBSr4pAAJKri
rVtwELcL/wtMxd+pjwBimr38j0WDcNPj0SrvEAEH1DFq3MNFgLVbcGgwQL7lp8BCKSE+cK8Jsl9T
5X7WlPTDp3aY/UOEGh4fL2WhCO8p91s5G9VzV1XJAzHxCO7ROvSk4D31eCHMeJ4ipY5iODF/GYNS
ioyFtuvg6L75B0qxeVs+dchzMNxwS6cwujq2m/lX6RODeuhavrU3lLYfOzuWQ/14Hj7coVZi6w7f
xIMmd9O5m1+AFd2jg49GdO02l1RKkkI/wxCd+IX1mXZgHikPUmgwk+IDZJ1BHOCOrbzAeeAoiEoN
AeoRLle00bb9tzrNf21aWdyJdFLBJF/fUEpqbY+4Ej+cKEK1i1qSYxrvGQ2ADCW9CFMd/DPg4W/R
L54dqRCjKCUrPShHfDhztzk4GOkMfcD92bvqKfii3s0Gv7h3/w2qUdZb6+28agdLfUpNiqLttiDM
/lkAbV05XgeFVyRVzUDf8jOay6d5JXK3p8JzwtTX8bHYFAStWDN+SB/OqAH2HLnm3RK5Bc+jSGOt
8t1n9I2GTDbwfFQeE6e+QgehmXSGFLrc7vQG8L2Jr3B7vjQklyDGb3pMucBwtLybYiTd72U78lJN
hSeOQXpZnxJggew7M5Pi4gcT9hM+zk0a+GqBZ8gzXg8Vxwtn3BkFYs0973BMYMn81+XI7IFOjuCB
rPcen0FQbUD8oEybko2dZFh1zc+BtRvQ3OuytMDi83JrXYMofZjYKa6CmBb6hITxCv0OfFosALJu
CoyNN7TvO+eSnte0Wlofy7YVKogSGmtfi4XgYoWOESZNvq0SbLD7O2kNwAXJj4XWbk7tm0Ltp+Ei
t++LwQ1OLtF3bj5OICFwbAz7kOeo/cyoTEPQtFiVOwJuDqagcd9XPh1ohmxEjb1KB3d1PDFvNUOM
btIwfXCrRE3mFAOnN8X3WLISxfG+YOqkdCztTRpXs/4gA9jC9cWjZZQsgWzg6fzWkNTbnQoXIKBR
IR0NuYpBxiApVX6KuqTTnoyCthYziFDG+5JaNtPsTXmik9xTTChL+0ra0L2n4u6mf1eee4E2I6bS
lvHaZal2l8fyyfumBBVg/equ9lLklhfGm9Z+YaE3mByaDgZ72s5OgWeZRvvdgr41NMPNxn7cRP0O
b+BLIk6V8iswRpgYqZA3f6Z6ViOL1k81Fk2EU0oq/SYL9o/tchLT/MDREPacdlbStSW3vwLSOjJu
4Ivv1Pul+hZEn68lv/KMdSJO5db3ax8ZTtXUkASeYtd4LbnV9RX+iecZB2HZcLpgBDDOgZLRh1WU
i4xFfzt1SLtIp4UcQmSLLIjaOfRWwK8czr95f+TtiVxRBpzYorcKvNjIeo8ktv6Z5lmXFpJyXsru
4SJFAktd3FWjvDfZlmiEB22bfzy9Gls+YIEMokYC/AOd8h4BT7mLchRkK17+HekLvOn9SJv2p6UN
dTn8sid8x3QF/fVCXcd1sfleOxT+P7pvC/ROyxAOEa/vAkIhwxscFtG9SoWxz9BAIOeMEKbKV/VR
U06fowljN/VPwOJccyI2hjY7bxOvYo/Y59uLRuGt5VO553iG0h+fs4vwc76vYR2tl0EoTCg/0z/T
lOTKwZg0stGAJga9RWmvphsQjVlseQs8mgNDSS2niKfuxTa28NUHTa7DwUfNFDFmS8J1N3EFEg/3
cBFpaLvXXUsmtwKDERuK0XUGJ/4T8sOkL/aCzxTRUUt8jzqjetWqXWEIBPvFg4DBZjQtwKJ50g9F
uB6xVml7hoMrxC9T2C+yPI2c1e6DyGCrUEKd/mf/y0SnapCVjFUg+M8/g2zq2xDLf5ycjo0et0mL
2bO0pQof3J5qMq9sGZT+hZ44s/ECqxl1vviJ+8vsDW4KrQTMVgG1PhGWT8z26vBCHZdtaPoWlS8t
OHi4rimz97L7LemANR62EFzrTOju9YCCLAo4WvYXut7+tFfInHv0csc1MpgUFIiEViRbajCca0fo
0gDiOMuLdyQAnbtks2S0yLngcSLYNsLxA7PxXBKtGcZhCbi/E1bnq1MBaYsSM6ZP3PjlP3SU9alG
BE0K+wc5Y0kdpAU11I+DvIczFxOdNsEMRim1zv4nGaeNjE7o9wkihNBeEmxIVzIqc0dl1YEcSphW
HPRDdTHbyIeadrX4b3nX61SSmvM3OQDNlfT2ImENpiwxWm5gL7koyqUPus2M/1BCF+noCm4CWeK9
Gxu9glR0RX7EhFXT9jJoZpfJSjsvNjcicFSoTj23Ti2F7ZDSKG/C6H+d2Fq5vdx9RnFT7Ms4ixt2
n/X4nkY8Lz4ZpAR08W110VrATK/FSvr6OxEd2Ug/aji0KXMVCZLLj8KqsTSOg0Vp7KYA9+faeNe7
xn0MSzEv8EzfKVTwdHhw06q4A45bHGPrIU6fU0K67auPALeWYV+CRNMrQLq1vCQQgNvU9UswOCMq
aIiEy7nHxCpPQ9oj8ArjUEv45D0/8/uEikjtkvAF9x1y5y34/0AY0odB3xvMg5WJ0FNraTP2Mz2U
pckzKvgEqw6hLGDYTeFBeofnZ+liYYtdXtQrZCZI5KJ7JR7xCaSUuh9651z35QOEE6fhS9i1yoln
7EYfl+zolQ0Rr8qVB/HGA8yfGzDUM48RgzwcYyMs/EgvMARDpjDryaMKq3ZBW329VxTApRNOCENc
yAfywU+GYveTPk6b+H+W1Nk7whwIeWoCdIrargW3FNbDkJaUiEwIEy6OC2CrjCvfpSQZLjIqmYMx
d/4aMXzVZDQC39WX9mdt+pKuJKEZcgLvcBS/E9N54oZroxOkuykXEW6anqCpO9eUCDbt76wg8wtG
NhQsyLs/4RPiRl4YoU7hPtEbzk8vYLZEbfv5wfA2jCEWKePJjMr9JHKxwv6bu4S6oCMlFiYZvIS3
4HVyRN2SEGGWkYg/5XDO3lfmUSvriTvr8Gv6ZJuvDC7PqwTyjRjHUgtMlmRBS1u2mFMCK8iSYwyt
zK5+5hvfJ0MmG6xKGdPk36aZOTPFcDSeDdyTVpoUgNBfbbV1DGXQ5zDLQxrH4iOMsm12pXio7iPZ
YyRqYEJIna9Uvg79EDUatqodvj4xUBS8dS8hlW9NsGRwLdI5H5VhKpEqkWBjUnTXFJ0LQy4oC+9k
aEAH4wBUNKcdWtmp0BMA+MBazQLrs+L8lLJ/vso9UxYiauvje2Z3pvX5KGRF7HezUwyB7mnp70e5
gaRo6JLeB/aPoZ20RifvVBPIc2O5yETzLcGQ6sPp51JKHPNuC/5tRCR8KfewU+LN2JsT9eKYhNfK
mNrVixQrpf8sdCQm31UoAl33NIXygRXIuEDmqUezAYt6ShGGJ2H2Eqth3HMFhralNhi1AHXNpiDK
eKrh/Q4hOVpvbwCJLwMiiMiQobIr481sxDHc1zFu4ZwzvQlAkoc20UEoxujR7Dm8RxuFBuFZwyTq
yv7ozBPA/A4HPMbD7g5abSw9QFT3BRpBki+TfBAqbEyGSWiX+ASGXtCicwpnDUF00K2DYV3M5jtC
ICO1Mzkudwfn+PDhrxRSVSmLYsM3SEavWGzao/xp9FpPb+PHFJ//k1Iw3rVxU+2vN88oY7nsiNXa
BKOVCCuy90jvQag48IP1N74T9EfiPrdOFaxWL5gHhOs4yMnUa+cWslk/8QuHgdxDB2mkBbZONTNC
QO0Auu8RpzzdoQ/oIvKcthWW1MhPszygwGNmn2b1DCULOWneZY3Dr5Fs9ECXIrcZTKlI4Vo6R63A
yx/1GhVUhrXv391m91DOq5YmqzHmlWGxZQvSb0HmtQJxj0sLyrplK79C/FHTY54VRUhYTF+b2b1B
e6qW/LYY8Ylk+ghT3D5swxNqSoy30sAMme6yFi/lQ7IAeyAzk0v5AEdRSjNlH4zFNwAqbtYAdWEa
1ETqhbk5GQIlGpnfCRpbl85KWo3cvnLAuGeNs3BjqsS/azrGAX2jqIJR2iFBVXQOA3apDvr8Benx
SHbWMKBDjpuE91NVSVq5QNwlVWZ9c1yAcM+R2tKA89A8CekRjH35SWTag5Z3J+v3XjaSAbuRAOYy
DYu/6VkhoRBPWWU6n0kqJNRpLSjCs+qFD8GGduU4VsoD8JJLpmhDuHCkYNlStRA1mqU9hNlw1kOf
2h8tkX5lMmszpK0OW9Uzxf/Dp1Yu+eKrUXj/nqeFAtt4vtiew8NYolHPBLym0dkjo4JSYcFj0LOy
FhEUPc/1gIBvtwIeRrJ0YwioW46kvqgTx4Ka458U6Wlf2ERfRrKheHLzgqk2d0/YNn3dwr2jNUfk
02W5gfN97AeGW01NQiaxBIa/t2n0ArpMQFgIq0/p4NtM3vtXqFOUujBYXRim0pzce+HMOiOGvqHi
HBxLj5WzdqBQBHINR2tQVV5f/XoTiweqGs68e+JpVgRYbRAB8IpJ138ArOL0tMDoxPjF6mSkuLHd
2Do0E8EG7hAECfZtnqk2tEywVOAVTGjUkdjH41Qoq4fpmKp4LkMuAOUM7nMExLkHmErk5rkdZYZl
9k3VUyjVpf8a4MxdNvaUaKTlVvpJ/Dk20HMT5SaP8F39j4MjVsF77H7qYs6SknkMSfLwFNNyIwEV
8TPOxsfhyPu4QAcC23FCDTGgYoYOfsPY+QUFNwHttKwLZKdXIxYhSZgPnaYwtBoSHO+NR5YhtY+2
lydsPseY7BJODYKkcL4ecV59Hzk/BU3S5DvRvjlYoRmFAdmd3uguF8vZxxcxXqiP28TsvS5ZlUOV
AgsJk/3giRO8nyU8bwubasrvIc+kA/r3A5CKcPe+olnqjazdYcLYYVTC27t91aQaenhg7Nvq/M/t
8DPJTs/3x/uxn62n+isFb6h8WC+7SJqaKRlDTkDWxcFcgkWT3kRIl/NSkGt968w41Mh21f6l6Qmi
HexY2safcRTCh7BhOh87D6kVTdw8P4uIFHyswXbGIaWY/gbORXqvFpIbFy8VhT81th9UW/GyPPo6
+cuATfLd27/Nl4QndHFlqO1mL48qLnLpcfbHTS3KLPoshsh4pxRtb38ByLJr1DSm/d2fEWqV6EQz
JiP/0v9Ad9bhPqiIrddDZsxVXyXhN6alnMmBaXOfIVwS3LXc4ebehJ2w06hcEYDIRoKcUA1WZoco
IDjEYzpfOjGkZRZnkcmHIW4CfJvYlAHJ2L6nNECKTn+DKaNzcoOgBupoh0PyWrQ2rfSRYvkd15am
rySzXYA9Pe3N6Glurcv2bom92fs0qEz2aijGWQCiq6zzLuUsyQlxzR9uUZ8Uym7NLIw4B3CqzLuh
IH0bkuVwjLbR7Tcg4zL/pRocfj6rk8p5QqxPLp8cFV/0EQSxSFuKnKQBLLNRGBLQptTFxwr6ezSj
WHwRzAQsGdGZDAVAJ7xr7xchM9FkpzWWDtnx32vIOZJAF8/y0GKHQVdUCaYLNN51oCKlABsIzd0a
0rnsaUco/D1ZpP5lEj8h3kI2vV72aHGkWDUAcn7fYBh42UDW3aJE9+Bxt7lJ+JuQiItQnj9Yscwp
IG24AM0Q1XKFhGF5Zk/rTZ5FpwvYqPTLgqcLgNokeWYWQ+I53Ct3R5dIAc68slrsRjfofbl2RoXF
RqSU8seaSYUo5C9XlpmVz/IKsbcdi6nd9ejRczUxH1YR6lc7vfADnE9dGZ2E6M5xcDQ+F7g0H0kx
s3qBO7N92yPiI+cNfoVY2FNyGGpyGYQVBS2L2tsLcix65Hi0jStDT9ZyZ30LJnHplYZPEVSO/0vF
b925Xj9KGEfsaictubGPGrtUqZPriCn59uLzVgCsSTjyUO39xU62IHfuIXcpZO5sVPxwqxSlCby3
yq8w7SIMuxc1/0BEbRn1ufS2bMqVnito52uW/M33a0PK9F39dsMTkaHtbisqaMxRr+7vNn3UGO9O
ETXy6hollp5S18sZgQlNE5dnLXU2tfND6mCVuSfRsbhvd2jNCuZkkirR7oWgnfmSgzF9ExkSPRiK
r27+FQB2Z32Glrltd/Jw8IPSNkrqewekyEyp0TVTCh8hXLNsW5n/OxsYqX9YmSGStpQAR2yquljw
5sh8hgItPdi88G5yE17Y+SRoLWg5vSfFB/jZYAS0OoL9hZNUIwvdvce8al9GsSe30g4BudVn9t52
J9OalnddAideKoB07B4kGaKrR+7bAue5/sI5veR/Bj56JTOkYbSK4qKIY4oUsjyrlgh1PluZXnRp
2H9SC2eR8RQQwolfKFNsbA7rX5PaAR04lxs/laCZLUUaNRw/4GlE7mfmn5bkn3EMNl6U0esyj5SG
u+IyP/YAUXJOv9NUb12vSBD4jyQ47DU0ABMWb3OfvNyysm9Aj/BXCL8++8SsAIFBB9CYvOUCAlC9
D7SweGTWeHAj4rp7Rmj4LL+YqYdRHWjq04TMY8Fn9jZl8ItMc7PcVgIhpd03SLb/sZJGNRecxMQr
k8XuFOaVlZrimrSoIjVZsc6wi8dxEp00gKZi1RTl4yQHgB0pWXAAUMqA6dc/XbhLhsSPwRMJs9YI
0WRuB1OJ0wX0Fjf/AaM2t+eLPr9r7nIndJkVol8LGS26AZAcETCpxc+7KMNcCD+EatbiXfrXMtsW
2fKUDwQRlqtzMjrY6Nva7yuaT2AKcmxT6jG/eDaojWrlGfsONkSsj046nD7NVmOyNKh2YQ6I5DBf
x6Uib9h/UISoA+wBmtX/oOjrYAsxZO9LiWyEBGuwEpB76+Bkco9txs6fpwiG/hjUTmo7PufM71Oc
4Ym7QGi1zMLPgFVuE4rz5/S+/dMR4e57XB4RK1d8elIoUjJv8ShYzqELgpSYuYGoO+Y+4JjufEtQ
IAaz4XccgO8Gl87qpJn1ybseW6gtNxw3pxP5mEG4SKQA28YqsLfEivXFxhxC+DBEOASjJJ+f5qTO
AxKVDbx24bA8kJ4CK59r4hySNQP1jJazm43ObjJXPb53dZWMK8RisZYYYNISM9PBwLazeB+XHYLd
b0n8QRPCSm9tHTwLqZLrMLUlx2/yG/8toJYlZg7B+GEmT2SfzDiuWL4t6pdKnvqTp2I+KCDTuKca
KXyS3aN0+5g0ERXjG6EWXg8OzW603Pkzh2OJQQHXm9T+rrTsXKciUqSF5aCkbloB4BBmbX159xmm
oFMQ/YiOW69Jy/hQpHpEbNKfwKqBXT4tN1cV7o2gWEDoYa0O+XF4Fw8Phvc/n/8JwqaH1XpJGXzp
E+BaO2wh88ckn9aaygBZrqaJjt2DZ+1Rg5PWko9MYKlinh+2xb4W2CameFdo2kAVdurQwl2dDSiP
sX+3Y7HMRrgWGu0lceur1vSeGvFnFhrn00LhPFXLWbjX+GT/lzKCe/DY8/DepuU4nH5lzaw1Di6+
GTPmB3iaV56sE2lBBeC8V8F95Hb46EUpD3mYVJC+uh7dMGrcsT+w+OY7bjzXlEL8NExoV2vwvhTG
MAH4t9FMSwXxnoc5fNTQ4CxIyv/g7r7GMwfoS3JmNHfm8jKBm+3it+7mbMJm8zlqxe9C9nP1wlfG
GyhxiTLbx5q+IcQMrobhXfS3QyBpmuzDjhfKczFL+BDTq83FdtKgP3mtOUCODp4ykyGywEf3CVfE
+r4s/Jsky1wb57xYMO6EybzdLbfqnMZnGCvehN5v5jwreSWrHYMhy5DLTmU5iBSM6XcilwQlZwiu
Eo3McW7l9udSM2eO382ud8NyomvMne5V/U57s1ZWqg9i0TeuY5WCHWYUvCnc4liuEC1JcbcVynQ0
BOvUHqnsUDxRN7ykbZpTlL5XrWcs5x3zHdaOz72e8ngnnm9UexzZXm400dNrrb+nxY9aUDrzeI6t
aeCSSIXhHl2ntFxrOsap6/+EJHcknqLh3SWR/5kPJTsWixQpIOTsHDMFP44Li80xMfe2CoqFwnK6
Kx6fz/nRFpBfNvcqOrdnRQK+BlRtLJIe7EUVdBpVU1EjWhuioKfaJVaycWazTf57FjDdMQraU4ZJ
kBcPZQeBZxPw8rBcYZYHA1SSZC8nP2EgrPymDZjFS4intmPa3RZ2TcRuAdX6B7UjZ07xjwmWbzRl
NQGvC/7P/Jlu0E3R9b7trPM1zSBEpCvhaOovl75tNzFTAFo+f5NQXNlJEYWh0qWEdAoL9H/Rj3PT
FUQQnnfyU47PBUNaZvrgRG3h3EWPLV9rZf194ikagx+nB7YdoibQfDehjhg4uhUofdmN7tHV+JJJ
C6VOW/Pk52C85h63bG1iBb2NvRrrbzEsJzZ2Ox4t9DQRvvcCWasIRS2vTSOqU/89EKoJe9UwTRvd
Wmlac2G/qKBEiD4ySvtRUF/D96rDbCbJVwiKxsffD+b1Tipque79jTA5kYY5I9+ADfRbTongRRIN
hFhuU+mypixnkmrpujU0Y85ZQFiehC5fdIYJUe5yhdFJfeOwbA4JYiKenw4xcgTNP9frHiCtWLjM
b7uDtm0YjvsxMH6lP+ZfHrl5b6Ey9K7bRsYAFI6kv7Ehxd8eml7jfMbZoDqKfBhH1tiITr1nTmFd
Ve5Jo3IanlE0dEroPd/YGJJDZjnaxW1amcsmScxVSuib+AJpnPltfqsl35FdaCBrrqFmwt+wMjMi
x90rhj6ltOzFerd+tIeORLgHfWndp78jtG84IqeGtgbQRbyy/fu663Ytjq2PtlQi/jhG3E7zulxq
yVNPsG+kFgE4nZ1W2QXhRLaTpFFwG2PuB2HacS2HYOuWRS7wFh2RMrLhuELoyMtC6CDBLYBA+xvW
NcejHw7sMImLMZFdtzsQ2e+AS1bDayi6n+s2Qhamvx7AR+YPjKUvX1AERYe8JJFdLxMS0hYqQKu+
RuFjVHE0Dqs1Co9nNbr1NOo8zRRj50V+9M/dUkjwjvQ4jCKcKOCiFNRaYc3i+5ubk2EgWTUXfYnL
euDvsD8O1NOrjyDNPEmzY+EUGaDSu/Z15EHxm6cmqQxrxX3XqZeorjN+u5eEwrb5hrzg6JKPGJ+r
dhicc6Nw8F5WZHVyrI84c8bbWAtOGQduHjQRcSw5f9QGJ/JagApP3mBJuEZ0GWZPKCdcb9fRobxr
7OnJ3qnTUdutBoB6YpuDFBTSge+4XTA8YS2fRDyX7hLd8o3R2dUkGxmyJqhC0n89FoNmhKxMW7hO
p5xuBZzYi/at/FJeTuZ07sWExtZxUA9J5tkfpSvvZXe6NuPXkiPMQjzDcxiJLz1qZow+yIebvk8e
qkjnt8MGOVQ+0s5fYV/oLapVsIgmItzTKMr0Whbu8gxKBNExENo2gz4j6Q2LncRKQRAfsU0JCKth
3uRyDUF+Pammr+oqfLGFvkWK4tMoSy0sJ8/Le05QdYlBeru0s6/rEUluI5R/vyITiEE5UzcK4pu0
Y3XEhBgi5HifFQ3JkGgESth7sbhU9TBbHQRJIpTK4rl6HWxl8k/7p9g4U4o/D+edZ/QuzYLZGwur
D40gpZrPEMFwlJtx9t1KJRIlaiHUtCmfjJazlBOJ84J3qn5zgP8FjdEIthd1QLIIWOJWS7ua+DBQ
1onjpX+Y717+TNbB8opGVmYSgkefG/nEveHxJO3xyuvAm+ENDDVYXzCSj03tPxEWOnuxnz1NEfvK
FS18CPByN53DjBlFhNMsCDV16BdV/EHWF+ArGIkIckOvgeWWe74PEF3AdKaJleU1IdxseS+GXvRd
P8VXQ1DUvhiAu6R02OkE4Q29oBhc8CNj5Sj31TwVHZM/K2s4+ikACbkgs3W1t9TWHtUnvlIySSdI
+ylSBvTPaZXl/pZ7xD+M1jm852GbLdTJZL0ePp62X0wKnlh1+lcoiz7flbOm2u98BUWQJ9SaoARf
AhnCY8EjNMUtqk5+cjl8e83pmIycva/YciVTnAw0ftKCOqdL7jKxNlnbOU4S7Fv+6w+R8OAl8Wjp
daIy8jJL83ySDIUU2UMVfDSIhJpFSAXqh8Ku1ERVWG9aRU1e/y0Or7d+C/6yaaPht61bHnFVkK9K
T+Uy0bpY/fhjCQk7+dy8+YVQbUbN7y5vPYW/hTfL2MAXaVmNUnCnXsqe9uMfiWbdzTW6P+pzIEfi
0uixAWIV80D5aVLBZRmD6CZXj935PtpK9iP9IFmKNfXWZFSsCDmC9aaZzvGOMtZeC/qbO7XWy0dX
5Z6tebBq892KGSsJO6igXF+yDEj5BjxftutTBTcw6Z11Kp5bIqSe+Z7RMmVZwzZZCrYrYVSsjQ2k
9jWiXDDqjO6nvDQDuc9SaRdFYhNTZpKJPX9gibPe49gUe5T5pb9HKek4v+22lmG6dsccFdIuiF6t
ekw1FAixwd9d6ihzqcDE5GtW4OSWqsg6uD9u8rLkPlFsXhq2Mo4n5GqmX9ZMEDM3xKuCYPksr8A7
kxF9AXcaSntz+mjaSa5KiwrmtiVqpUXi9hncH1vzCs2gdro1odNIupSN81AlezE8puGNh+iQ2NRT
YmIB10RSaBQG8gWcCE2VDuDvlmV2CXa3MeIvkNoQPFpKAiNOcdJR/8vDa8LCj5TIYbtOo3nobYRY
w/3jODySl2BgfQZjnATfM3xZp77H7sTOfLjM+ql5Q09BpI4WHka8Ymx+UrWuSIstgm+LkU7jR3HL
95O0cruNjnypKVoja8lnGcKc8ZfhJ+nHxKLNXgxOLA0FV2yayVNJmYLIQJCyhOxeooMn7V06SmPa
T0VABPr5rP6RQXymlgbXmeTSch6oV3etZkrSY/trETqNDjR5aJC1G9oIuN6QCxt+MiOUXZ1nZSVu
PR9TwWF8QwXIv2L93fFb6BJFe1XkA6BkAUH8kl+PWMZuExm9ySrm6ZN2EpLZzgbkh3logs4zvq3b
kyMYLk4Gl//xPXVJSwD/ybmQEOtnv4XvMwQaboDhPaTYmxUYnyn3ckEeNuRlLEiq80qDWa8gYlOI
AGY0Yta13WU5QYkVkde+BeUYSANE1tu5onxbTiIJo4XLo78FQNPjMaQmylWkDbCsvcMijse5jYxO
yUXNtgYK++SkgWcU9DElewJJyDv123TU9ixTDfUC3blqomINPsJ5gQxSfHQVr5usw4cojZ5K7NrD
sjGp2ptRTLyUkSpJRPxLoElGUox02sCUZM+WfF2Z2HSbadx7iboXwmET4/sVYYFf/9wVhs90A+ls
QxKD13wcicvDvEjNRQuh2ijqM8/B/pvhXLuUn5CayhgbX3xElXYJmkfSHDFTVT+b6/eHRBTF0rKy
Ojf5JVUfDZzGdMPZnWIbbVnyhRzcirBs8+l76VeDrHKa2g5FEsFudtUL+YJ4kAfgaTFvN/S0WeKr
vkMMHY9dFdfj8gixAtox93oOnnSQvk0YeHi6t34XtU+whhOoMxvwN7Qp8TKrhQLLtJ7HY+uno/y4
w+wDUY1jNA/8dgtGxsD4NJaHuw/RNqptGkoUQEeB0NgGhsbjDeSYLDsyWRaLsPMM0aa0hgJyQ1rv
Mn6x7KX0Vn8kFhNxmRLfXRZP/bip8V8/cHykd92KnXSFGNBHXsZ1oXhkiLL0OCWaQQnPuGzd3kUu
fzANq1XOo9hjYKfg+4aUQBgsXJlekpOJ/NVsHN4SSqEXYRYzAUt+RSDaX5dosBL8FjrhuunlNGsN
vVAf2DENw4AxxixHX2cgJn61BY3Euwg+0Ke4IoIqUZ4pT1PjHKp6hAbvcoUBdJ0mYPl5fzJsxTPG
qQjBK34zlCbrMbp9Tvt0PlSIEHp4gCIogfmLIrv50HC/22XvPkPXiq1dcma/7nbN8H/+jL0WV3mN
6dZJkg7nmCQo6NdhnwSXlIMPyrvll1xKskMBpE8CIvgHS87WwUv9LxRpaclaNnTyCtUyz80WgsKc
d02og+BdoSCpv6yj8VTSd3JMuWp+KxBn5CuRMt3nR8cPznyolc5ZkSxpB60RYFpLf4sSi3i0jvrX
LGPBWkvvk+iVprkp92FwK0zNcRJ8w324HpP5T+klCQTJUTuey0+/h7s+arJ9ZxejkbcWPcHy4F06
o3q5/mkWk/QN7mEj4H3k55mLoj/+zgRCjHMDAw5lcoepHQljGLFQKK3lZpSFy9DCor0dneozOv8P
qC+a3Vo4DFcFL0vFdsGDOOET3IrcccUqzuaNFGR11mMGAmbKQb7U1kpYtUyc1/+LB4m314KrmMdg
p8I29Fho/TNZo4r0EtxabRIjiTSWhbnEOcyBV+MgSmyS1ue5g9W/N/5qA5KVDwz49vh+Ph/DRTWt
CrW2CN32WqoPXv3YOq6/ppgILTq5dxDIkW6yO/8PJF/43M5bNOu5kj5LFcYr/TX+cJwjzxRYkMJs
igZ5RJgmFAJ3rRuvih0QYTgyRyG2UaK9TsGy4aL+PYunY971GlNoGlXDxMxwXCfet5mrYaXtKwp6
c0WTbvX/dmqQ/n9f1KdkQl0Di9f3liDfJ94kgr79jdsW9Epvz1L1AjpH1F/jM+q1Mj30WFsVaQAv
isWxUPGbmsNhohpkN919KvM4bexgFEUhJsTqle2KV4AZ/E95+ZIldRywA8N8gmGUJXlKSqvugOUs
sU36PjDEPZaKWRIfumw5T0LxgTVeA7Wm6zowtdXNMoIA1104nTbmHnMWaIhRmvB7uGA1TWegL+wp
HD1ADys2ZkAJ6KetO3ISfCPKguuCE13v+9dXx2jBvFptm8Cf9rivKpBgJljou+LpRH5Zo/5EOcRJ
gkOtn0kr43ZiShmrgNDKUyh0NcmruBULEwNxEH4So+ofQxOoYI5KQGJ9XroqYvZGRF48Q+iNyV8W
MCh6ZdtT5oHBQx5RgGr9HI0BWAxD1680FLCd59yV3UJSxEYiMkZoGZUq5IJRnnHhhBJIlGUIan2f
y1u0YMTS5PjYGTYBTmnkurH7UK9gKtD/z4DIVGDIr/ikfO1vrEXXbmZnmga7Gq7pIDDZf2gChp9E
WZK08MdZJfBaHBhSUiqXZXsrofig1jQyi/syCUSO5eA6WkBcqSZaBeSNndWhZzu5V41FMHacGtEA
0NcDmUbKgPvfDtWNwmdP2sT1UfixAPk3B6KtyHbM0pAh7UUO6YwEaW5CKteRcQSli3cw4+8fX8MP
moBqilbB5czvasX7GVSB0U4MsVQ9PXX+kXmS29/2Fiy/WPbrYR6rS6SWQ6X9E6xLP73gII0J/5s6
L4vI/hZDJhd+bokAdGX43NkfxiYVHsGrLdZTOmZJYGL4ZPbvAF/RwPcCfGn8mDJIxQquzv/EuSPZ
ipR8/3PbuacjUt0U1ZEjjsuXFU4KAyh2FlRqbMacbZCOiUMAWx0wyO4HFMMCBiTbiSOtf+MCEGl5
cEARvNlNmcJiJTWXZFJ28//w8WnJpzhI/ChiSYPGjxpI2FGgE51YPhtHrWu9kfMjN2N4AsFzCdNm
l53jtMxiyJloXSt/BRJPqxqZ5ifIoDzfzKjd3ZtioVkZQ0pMZ2XiNNiApWbIuhHF5H1aTxIJ+VW7
1bWhl7gwpJJOnnQcci/VIyivFVrGI30qIVarPpvDV62T2W3C54y5PVKSK+/cTSGB8zcQ3p+zAfPk
qfFjapa6Qj2l4+Wk0uiXBqPi5rYA5V/XF4W1BmfPlP4GdLQuU1gSahuJyrLFc66AlgfRB7vNrYMM
A9aAFnVdZXarZM6dp3cQ1DaGL6ODQx9q0YFm2jYGxTurNV+Dcj8AeazUJCyBbOlGFH9LbY0PTcfd
IabbmLrQAB6p1Cc17/CITHNzLHG94iSrtFa6dW09TWKJVCEkjKcqI8tsYSXqrrEaWd2WIvWm55eJ
6VdqVa/VImUZ2bfWXSK0FWiCqWNcBbzMd7irckILmIjBGZhJSPayduX1AUuNEVveEIG/hWXZGvYB
tiSINEVuuas3u+Jp3/t1pWaV98yTP7ymkoBczwOAp4VWC5tx8CN42w3qai17UcqqDGcwhGBA7nI6
b1o+dVqPNHdn8H5smHQKZwZkZb8qJu2ZL9ku+3zl0ZrbYXA92U6LzlwShLAodqkR4R4baizBWtY/
7q1RkYVWfZ9uADYBFT+xFEMC7bHza7a9FTMp+GudUwjkLtJRSkaT7TNChkYB3w95BW7xSPNuulI7
NX6tXj08tXnaBDAqUAFrmBg0YEhUz7uACnQk2idlbkEmrO1iXd/IsbVy4okyNBOBIwte3voBj7Kb
7aTuyVOCNht7ztMIVogo5Vbdg/i9xMnUKDnY+Kp7BEdchVb9qPlfc/EZth87f3oGg9rf1jghiPXO
ouu5+eEeGZlG20L9pSb8CHzBMt5Rya/9GUF9rfKCMjcKS36nE5+LS7szr1ya/sxNaRWsJLpsn7KJ
LZTTq+azd3ZiqpM911vGPRS/qUgAtqhZOVhk4YNHr988UzC71Bd5+NntYlzRDYDGSK67nCZqxFMq
sYl8uK0Flg2D49N9NdTEZ509i/Fj2IGvDaImAUHGSgw05Vyj6V5n6IQsV0dnVTjMhc+qYNgQBN6a
f7ijHWIe6O7F5c2mUt3znavwDvTyK9D1SfkYLYiqmJbWGD2AcmM5mPUeiXgsJJksmTsX58armrJn
6J9W7dTybBNsdi+wqRpXnsyNkdyzDfF00VIBNoQXpQ8n9jQRPz/xb4gplCYhNVacp2NQyPxp9/v0
gb8hYBbjva1OEH1+29FvIX311lNmkqVARgLm97SICeEf8QL4/AcE6i3eoZeNbPufJTMIWlLj1ljA
BXSP5wpFtBcPt6k8vdTeq+B3gTo1z3wYkvzrgMkR5PlQJhlklw7IQgwG5RT8vNStSVqMmPRiMDdl
72nDimOj2IuySHCOa+FN8LVVCYvAPEtceWds2AhcM+bpPfH+qJn7t3Sxi+vFn2GqATu26Bd9A+kk
7WChbV2GjtuKMrgV2i7R/+rvBVgEsSv7tMCaHTt2gNkNYhjkvrnA0/aUp8YmW7H+5xzPbYdL4qq2
+l/JOBealIlM4he9vD/FK3sPF4WjbuQGhfKJSV5UqNhzDYtDEZ+vKwcP8l1OSSjetgjviZ6ExBvt
h1uzROaNT8dbgb+jKlWmS+vogy1Mh1uTh8jRTjn89fKeJZwW3dkC1aP8BIF0D7BESC3V/yi8IwPp
bUa5vYiYrhwmpUo06xRQsvpp8Bz3itqDxQRsJxAyugnxyhwe2bSW5GWH5MV6/M/4upyIr2SioVTb
PUCfDJgNKbYzW8lCAO0cM51h6L+ZTt/Ji4BbvoKLNsBIMRQk7j8rKNeMoGqmlqiqhNf4Zf7OAaNd
LIo2sT+ykOOWq2j7CHriyz8PvzXMHePAckeMhHaqBEf6W7bRq0Br4QjTobnSWFw0ZVguSjLLPs1K
EUbajjUHrhwqDv1sSYUfGLeSj0KelUl2VDrnWGqS9hc+Isp25VLK8hWyntkzEe1WlfmYl5TCcYTb
/a7+cug3A9oN8ryeNfY7oKhSamV51MUNk5SumK1CjCYoUOtv3B0gbFGakJBWC6r6N2DQc5AWFJcs
NHuOCqeWllUM6nBz9DCMlbs0lUI0ARrsAthZ0ZSGL7GFr+ErblwN5InT9n8ROPCRuTJPrk5+w2TW
aMTtbWb4z+GP9wMe3H5P8lncyQJh5gcvIVJTgW4tA41QyHTRjY5Oryy1Xw3WV2s/Oq7zcYx588wF
XWv7hAqRQT8ImhaE9N/KfxW9zjzJHxRG8wqeQv7xvJcnsYKfUAaEbcCNe8rhl8/MO3KvjCLh5nhP
+ZqobubL/66f2Kd0iraXC0cpVQpgFjGxd3ZqzSAYUkMjPCiUPChQ6kAI5R02IROO6SkYT5zEC4hF
0+JWSpsEMLyfCfb3TN+KVFBONSsk/mBKSaCAgOfeaAfbiSeG23ELqOgSlz4YwReMJbjBSjXXAfcX
jvhBcxdv7FtbMW1lCAn1x707tI1KHch5qFUtA+BNMV8jzO1bhIW6oEQmnnDhzl+eqD7TSkBwoqrI
VafcDedPOrFxQrz7fHZ5TaEeI7YfM0LM1OxP6gKgHTFjIQP3SKgAAPw+YTdlmQOx8IB+DsNYB2VV
q94C46mF/9LM/SoqqdUBIKUwojfoeI94HYDPb8vMyEb+awH716SPCGiXOnSWQejcIUBifjnWqAUX
j7ZtV2g5BchlZ67pqgoinwSgYOPKM+QWfrAQFjSQRJMP0jqUizVRQ/Oy2IDwH7oQB1bkTAPQrvU+
5GeZ8D5dtl7CjqAak5jT+w3HAS71qczCuKoCnpW6pr0PJFlxE55pI49SrFf/RobHKH2FDzQFNQcQ
/FQnawyeVMCVAh89KvgUnlxc07a3wz43YHnjqp8avkG7H9TbZ4GNdAvI64wPtMGq1VYvYlsSC+9S
ZovRcYRj4/KYKSPpMnBsTzBEmwIpMjlJPBmzjxMxLfh85XPesuUia/lx0/5DztZHDXGt1uU3hWhx
mI3XcagapKusY37iRGz51BVYdRho4t46joXfFxlwrSeiUDoWbvBks3AuhpTDP5nP2y6ITGepad42
aqQuduq9QQCONaGm/oHhbmCl5cPmne7v91KeXpypYscpPSAN6Ce3ORkY2kE6Mpnf1fZH41YUpJuy
xK6MeotUh1rBY8rWc8Tgf5FozuF4i54DzM4ZjtlknGASEp7fneSihvTEfmqcRC3hIX4IK5vP9Raq
YNXOT+1OwKdrHOHt7p1Pglc36UoSdo4hY/h8O5nHufntXGVim56b2Ann634EAZwUiO8LOMk2CGSC
bsa44xeGb9Z9vjlcCl1ko7BaXJGvzFGmxnnGYhm3svFdQPOAm4L/XuASh5Ug2gz9VQtusGslXytH
Tpm7cl+GtaCNbzDOZiH9VmzizGGwQKNKiPjKX9R/lPoE+qWbV2E2n+j5+lQlIZxXECKb8TamspkT
V8bui5aTmWEL1SX2OVtPDmSpbKpeqBL8oePWB3u+fqanA8q0ZL0tPFzPoICFkzvfIK9d7u82DKJ6
Fx6MjjtoMivJbwbJvbj8ElevA+NppbOAUTT424CCGku1w5os+gIAM9QqyDiDMjHP5C18m3oJMIYw
noaI/Xsdy5tTicuPTZ2t0voAr8i11w7S0NPYZAPmB0TU/HqnF8WSnjtbRO5c+1T/bRailQJFL2R4
uKR5J7g8U80euJFyx+3MMczT9jyJqsVhAZJ6vQihDLYjqcGcnWMnnWpUj1TNKH3BIu5UR425QJmz
f4fiRnZqe/j0sd4IJCyQRSo6txHtXb4sALrGuKoCcJDCItMEKVIqujC7i5dd24uftkyK/G+KCJ3Y
FzWFoGNayZY7pbLVX43cMeFI/G0BBe5lxNMZatMxgktJgdDtx9c+H0mvQpK9lkqxVdoHcKjWm8qk
Ni+2Z8GBCn4E8XId3oel8s2Rnd4ZRrbVd7214WPNbMrC+6pRVvvXWpL78dRupav06DoLJCRXj8gs
kn58Az57rJsFDpkwRehuSF5J3C6Kz0/EuDk2+L6vnagGD1+VxSIzoGmKDeDjjIWmNko0Tf6a11u9
TWJGnk2yxjwjOvXjIG8CpgrVbsL8eeSrskNY74r944qqN2MA0Nbb/JUHbX242tx2ldbexmAvMxJs
r+e5eSKV7V4BzGvg5l/eqV1/iHNuuMUFMzw7WwPC8/3Zsp3ewunO6ALr8/0PdIHPGkxDLty6t1a9
dqhw3gzqoiHQg3uLlLSjJjE5ktB49J1crUnydUAn3/ioFuN7jx7RXq2rpVmW9sIZMe/beXxxAQRr
Gpuv1E0XQygmWMmLpIjE4znXSVedpjFTdg15hbW+6AyMaXuqvZKfridPGx8E6mhthqizQKeJJLlW
lMQ+dZmHrDdLFxMEm2BRYzIKUKWlU1GvgDkpR/JV7nHy0ZVnsV1i0jDDr5W9sLfMf1yU1pG2peqS
K9vRVjebgWK8/qW8+rQLNg1tv6U5dxamO45QYttBzHhCTxMvFC0iQanDBeuTpHw0XxEgfxiymn8R
JvAsEz7yXyBSXyWKeFh7DhyO2UjRH2chXRL9ExcW6IVZvUB3MRdhLccRm++Z/QI67uotY/CYtqoa
6Q0D3ZZadiYioU8jz37EZrMicY2YMug91/p5fhDdL6xM21DqFp9OCYjhdz+kJSkmts4QcbYh7gyv
FEKijMsI4eQ31tsGyOtcgJld0jj/N45o4qvRmayu8q6XRylX+3PRou8w4+lhlpN4bV6SrjQzi6DU
T1MmWuauUY6VTZ6J715d/bt/9DPDeTVduMvNoAVfn8vO/JMxbBRoL47CRPc2Z/LViPiIsPH+fyVQ
khAvyxng6plRhMzbg+WajvxZdgHadDcaQl2J/SPdcJhrJd0TUKKolJ0saXtpOJcKfrTulTxE0t/T
nF+hFW2A44dP7hiJezhXfOT0BYB3mwrmHSFY3XpSf4qmj57DyJiAGjyyR/0wGbtBqhp+5k5qj6DY
OKQcdFvOB0prurbe3I5k8BHOFMlSQg9Qnpkddz2hS9FOQgNCuMck/SdtoyHmDhnhmyK8Sn3ylSHt
WyIxXFw3s4OxwKTFMm300illPivciySeE8n+y9KYEYsOea7cBFT9lShUecfNd4q9RCdlTlo9OahG
4Z0KWyixSzEeNqCVrM0Ydv8YPbtmZsOMgUp/Rh/bA27dVlv571VLhi2Rb4EIy3Yn+FcXnUb0BlhG
tQgLbMn4fmdGgFcgy9RMJvc5Oa6xS9F1JhkHjbaSK4jG2/8ORPLLhMlBFrtjw9f0wloy1VomtPfr
wHmJdBxjSOTUoHmnZ2tV7N4LiFzEwu55O/wfI2eASPtYR7zaejagEr3nKu8ZVi/P/fTrULSeRDis
WJsMdCse4C7hTqclL0sh5d5SWaJ7us686v0ojnCERd6aSVqQAsQvNJCc8ONVqmP0nVXy2Nev9UZU
eW0QRbOT4dbsfSYizv8J2UUfNoM32KqVKeNSN8nM9KfomsgqTc7oMhz9qLKIQw7umb9QVysJn+ml
Bqh3LG69PscnkQ+WQ7h2gAHB7MArmqkNzC1EaceybrHCLCGsMGR5NSh/vDtGvDTVtQAU5qDdFD1h
1lCx28l1WwZKVSarmlZwbPNhfmLnHhCIw22pCbJKXpwIhmdmRTbae9o14LVyCtBiVbXgA4Lp6/ec
eCwLXKL7Ip7DaXul36S6NX2P6b61BUzqfD/2/XLPrc6BJ6oSV7S1UZGTcmdtXd8arEJ5y7vcnWsp
H8H2HaapxnRje/QYx5buxOeRqmsUi9u5br7XP+1ltqldv3cFPDBsxAtChxtkcMBi1OPO2OT8GjBj
8d7+vUwj0D/zB/1boMSiXlwDOrR+xxPlXXFsDCzuoOx83/kXkYIRnpQSCnDO1hXD9f5syDL9BXVB
A+hYkLdIWyZneZjUvDFrccTjqx+RlBTCc0lOM3SElWaR7y0jXQqR14Ht9BSgn2n5T9Knx/1MVQaP
dNquBegxK2oDhJrtwbDGR/Wzs+dfwZ5gfzFPx9IKhPyGMjxRMEMfM6/2nlmyscz88nshq0j2Cy4w
TTBs4gcoDHmzR7C3tIml2ntRJbz1LcXABJQ5X/gdQE3q+zh95SHoV0j3PJ3Q8jNMa/w4BUsNw8sn
y7N2i61xnOQthEMLtg0YmhK2usZuZrS9JhbDa5ePUkyjY82087qnb3+LRtz4ezeCA1Y0XJROrnY2
i/rMuNVyCZCQGXDyYUZzJDfh87InZhcRs7w1rUSye4k7A28y/6D0bHcJQNeNaCxtifqnT+mADCOv
CaEbR5IrCJRss+FN/U4q1bdMOAYuNjB9oF4Z8ukgXjbun9qEkS5hlXwMHgshlGrcmRw0hu5EKs24
6AKExHpdj02J5jyExNKgqslObYCSqu1G01TTkmh9GRItqzEu0Bmau7iXO9JPvLhdTxIi+7k4DBOh
FwRndqd+7gq2uMX96QzoaaKwpoy2uUGF6wPOEcqlRQmZWZFAodm3ECv4fSsR+aJauKHdgaiEeLWL
HixxWM1xM9JWpWlgiljvEg0aFvnZcqMrWpvttmC7RjaS1sYdzAe1qoRUr12QZPfh5MuQw8w/niH/
Zt50HuS2QiMHbmG+xKdnxfd/tB4koAyWWgxiE1dNqOPj59hh7A+l5RrNaNa7sb87t3Q7m548rFcI
B+4ihdWNMUvtdBuGNt3uqVRBlU6F5hE1Wg1szhdYdrnGvPOMEdbtsIKjbSKeq5KefCMytaic+KKg
HTVJQ9uxA7o4ylGZjo4lfJNzeB777TqLx0Gj+4YNr1naAqfL7p150vCKVaKlExsJ+6ApP5HUQSgo
P7czV3YedFNTCdsDf27Aru9YDME27JRgEvtsfYPzLSQbjnW1i/BIvHNeMhVKx61uehT50mywyMfU
s0nt1Gv0MAUwI09byxzVe4a87jA9092Qsk+/9ZnbqFT2+CsYtEtPHcGeBSuunylH/QP161p1KUSy
eiidNul93cViUAM8K0TAeHJCSxWV02R4crH1Vu58G6HMKbh6lT419r9WYchiXrEJF8UK54FcnjVD
YzOqnLhwHTNUITNtxHL8KsNYUXwiCx/WfAA3rTTcvJsrKtIoHYI8hoHibaD7FHmuuJSNFcvd5HuK
w1rN0aLB1my20+DZwRTblVvrbsRj539CzWOARIVxFItCJr67+4nib19e3QXqHznVlsk9CpeVM5oi
eQn+aWJR/0ak60KQRlc9ZHaaaGLtv9clcESymrlKUxlAircGWY9zD7nW6DbRVWibOk5AHNYN385Q
cJlbrrWyfrW47fIlDwZev3+TfmVCxu/NeTDfkFpGeh5BgJ87EZT3LqZFMmbTnfd3odTzW9tl2pNH
A7MnBQBHbGtN+r/h/otDw+fBmzcorsbqjoZxW7wEy/LunPGsBinMlYH3QENZ8X3+OwDhxijEOvch
nUFyOJtxzK9y+uFLY5P61dIsITAUvY0d4bxJU+dXaSHKDscC0Yia6bN3anE3Rim/UNwWArAoRIQI
JSDSe6ZZvznQDbNUzSN5z69+cPSL2L84dPVS2fpW7aY/OTAeck4P/ZTU3jv/GZjr+qbMo7cRxbRp
87yWwhle2EC/FkgZrhU5kEd48x9UkLQcx5h2PHCaPhB0IlUZP3iU68G0mji6omFoOcb8T1vX36gJ
Snpd80WP/ydzvmMxbp8Ce8M+4RTZpMNi8yBhllBzQvKa5jnM1v8mMAmS2tySJbBKHFxxjv645vD7
hvw28PDzLu3lgth1y312Ut4r0zb9IVOHeD7ZpjXs1xlmGRCtiJ7IV4LRagMSVqMsvaQvFRPB7+2E
zQHcHImLDM+wpfE2csBOZMbYBzOUYuIj7a1NOhFizECHKs0+Rd0im0Y+ho5dcIEENI12XdPNrc3N
OBkE6IPewMBf7VOYb3y5uUzdx+0Sn2HX1h9bIGeWT7H+RvPfXwjEdGE7KTtEyN71zd2gDg8YU4j0
iO1H8t40+3utqlzzRjFMkRO97F4SukHeb+NpNscNGdE9PsYFamlP+MrBUXMofeMR2p+wV8gNRPPy
X5thEij51pkdYMKj8FlNviSzxyhcC6VDBDdB3erhCaDTAHtlatal4M56Aaud6+Rvzc2UeK/uCF8I
5pW4qzTXzgZNbil9hkWKJ6TpvLLVrnyZPZlAETyKvhGX5MiM35lA+cW6NfMyobiJ0TLWQ4rpmUkA
vDfT/wcDrLflMgzGFwZ0pS/Sz9W4fs2PcNs94nsFk6ey0ktvtBCieEZqqJdQgrbCzXPHk/EMshVd
TSNQ016iljsZpffRpiZFOJDdtAOFL4AwC31PP02mqMIHshIDIGsw+P5rZ2gisbG7TdhvtebSdzp0
f2ro7qSTiWZJFfcqZbA0tQZ5oILqKIjyTQH7hBhiZz4GAobhkP63RBiCTGeoC0UWXkqDmNJPT0c9
Pq7Xm+OETMg3vHMZgfzeCO7OnE1/A0JFFttKDM9P1fHRnHXv1YYhpWYTSQVwk81UwauiZuJl6kf5
E6ZtrNpe2RivGMBINK1OuX4fkW6jG5FJiGHW9ZsuTKb33UvukF1fHIx8WHvYk6KtrwOqbQ6JMd5+
kDsCbJh0xYbUFvM2d5DeMNjExh2U6hQ3KAYrDZJ2/HgIQMD2wt7L+TWucCOrz0kV94Vut03NRryv
nDEGR7sE+DYH5vRYty30K367s+JkvE8UpVypiusJ8qAFD1gfRcYY0bde8rnoVIoMOgyhdB0TnnlM
4YgValam6yrFCahAH+7w5eS3Zm8E9BTJtYhL/fa2i04Dfsj8O8kHfNMzXF0Wm72cJ5mn2P3tbJB3
vQOFXVveyA+ap/axBKNCz9Vg7/GzNOuymRO+8OFQYR+jxjz4/aUCDC8i7R9q756T2WkFhKAEPt7+
kvTXQkGQpvxHL6wLFVcu/6lopmx7XDqA4qZRc/OsYAgwbghGrbPOngLgTPiDpBP6LsO64IIBKkPE
A+KXCIDlX6692zVfu5miHi5bv4kRg2E/9IODeVhc0oUu0vfspBEDZYMxkPkWfvw+zAqYO1zr2euc
XfhYyxcDIPDPMNMUwZsHwI59m/3bDlzymxRRizR0eENrT0l6N1gjIcQB4l+liGWwqSbUfNnKRXuP
5Hp6DkKFxbfw2M0DSFPyi9L6xaDq+TmPQcgj2FQ7c5Iz0fYu2b4DbZKjSsQyfOxem9pl3WtYMLNl
bN9UEqr4Q+fv1y3ev6IfiaUqYzgzcTSMzZqEpJyFov5om47KccwhUj+k53ITKgxLNfXlbFdQbiKt
FEB/AHwLel+s4C/Xv+2iem6r9GNFfU+pv0Aw7gx3mzEIbEJbs9X/lCgIWbDOj0NYHNXV7vHCkHaN
XK3pmXwzs0wltajJqMkl+npqOQmhiJIoVa6NfQo05Z2quGRbuuG50N5eL5W0AZiUe8KeB+jQy7wA
6vPkJlQR+EIoIR6P5QDTbrMRlH6LolVOfmyCgQtLiOULSq5dDK+Z5WAqtplHfQzNgDo/7ueEbu1j
s5w7tRtwOD0k6SOuOcrd0TntQ2B/KQBexi48UasDRk8yOYpLuaHi64AfCmjSkXLVgmJ6zjOa9Ad/
RcwtTIRxL66QZVksOdVgTbv7piOpw0Gvh37Br5aJzcCwgq6bApb9CDUk8pkea5+wTIVDmuR7mR7E
weMtBddF9Z8pVXJtG0007dcBRfXeAC0QcfFhw4BvFdYued6e188adwsSz5lwywksmzw7OPPrPNWv
/IQgBtDWM51WZ93ZB7WHHJnWiGXcPeW3WUgL0N2tzUM7JQgP/r8vIB4v3aH7fBnbCRkgauHVulC8
eQEgirjbdE9YPAVfnbLxsIW+YXCmh1oADGSOJn6OWmGd6N3J84OCoZhOBPIQCP6jaDoSuU1p/9C1
1We4yAGf7+FtnVH/Da7BDlOFMJJGrkPfF7cObhMrHPu9oSkRzy0zByJ46RSL8wKv3FmahorpYprw
Y8hxG+zm1OX5wRDgQkJQHOJsHg6nLzvHmQ4PGCb2XkLmYm4A3hF+8hS5AaXX0r9x3xr1QcnWPeLv
osi9zHJPrhQuKm5oQO3lmFgYZ+fY2/UfB+rKbqlOSI2JYdtF8R5sQk7JJQUFWmImIMdfcoYFlTeu
ek/woC2CHymfh9yknR7nZg8+zRrrnNMuOtJkfQ2NXsQlB9fLh0SvJisxey5YkM3oFBGt4799Lzg8
AYn4HLmYR0C1WGx86RsrJ8upjrmZCseGZBdozInjAsMUrYCy8vHxyy87Kr1kQjZSjr9/YARBmojc
OMQ2VEpgMKE/Tk8cyU44BsA7UdROxn2Q6k2142Nvh/RCrl8HpACd/lI5LXkb1oVgcpPkbkBau1Cx
/nsoHYek6MLxOu6DuxDQ+RBWgD/HqPD2oNnIhmYA7ypaqJNQVH+JoMKq4ilV8gOMhsN4FTvOwJxF
T6xxo5+f2ij/aQGWhBA2cDN4qY55SivLxqp+wP8A4KXDbws08t6eIMmzaUU+kqRuYJwolnpNxoCK
UbhYYGpSfMqXR6j+eQxPEj2indnC7oPRBAV+ZhFkvhYMG04ySwRtIN/Hygl2XCSh1RukgKdP0Xah
ykSk+CmbxO2p0c3tILaxCoOm5jvHxtue5TlQRp5t4UhC1A5UxNoDREBNwvH/Lyc0VTkJ3sXjc5rD
99aQ1KAhCXe3teSn9RnnuzaPuJLLMLS7NPcqFV1JqPrt76iltaSCDv+G+n+kpb01L3Fv8t+fxApF
KWtF0ntMU7f4M7fQuofl46DVFct6m6AGH10DL4b23v8LYVXyK+guX1tICEC1gbO2SwopYqIc5tHG
oJvsrVKxIc9RLci0GtjjtHwApk/eZiJSmulOUlUzrSbSth5CBvX3URchiswBGi1pln3fjwhLLa8d
KfcyZiqgN2ncFzfAx3R4chQuzixbk7MAlMiRC0cmrEaatGzmE0Lt9dMv46phgNQa9PgrBTa12mNb
h8OnkSuo1Uus8soB9J9BCwniqK9+a9g6L7RqTQ8A6C3jYUbth4lFZXz3rdzVgy6X9+h5H8/R1mFd
RHFR0yysFUCHcQ+oaBJ4qpHpnMZrHHD+haCybOQ8filjB7Mlx3/YaFkVvfA/Px3F8hyVB0WIQHfC
KjbAF033rOGDO19etbB6ECUYDlod0zxIDNvekpf+qF80bqfqsae3a53aD7HhHysQ+klUrd/rQcaG
hdhTEvOdsVkItMNp8WsCUDixNPXJRFeY18OV3/rXPqDR1EuftfCrGF5APv6MGNRR/FStd1uv5Mzc
abbNA42nQvy6jAn6LZEpbfgPf4l9NoSabpLU5haiOAYtgz4JT5GUkg/VAeYCPIRKpeOKg5ulN+N5
WuC1ocN1fcXfJWZGDlA3Rxbrfsjp3NtcCsXX8I2N/OowTPZ3FD9mGiA60/kPfE1/qh9gaK8SFG5t
Sc2G+5r/spn8me6taXmYx/d/dRbNVZFDl/5KIDSWEH+3ThnlPm5OKy5Z3ocHQLrmGgVUYm8LigB6
qii0aijKUQ1+46rANYfaYF4rFQ7EL1W9JYLSvQM+yX5sW8h7LG0yMPQXmb7co9EldIl1PDuYvfYS
H14lw4bJuOgPBVqYqAlmsVsvIwpam0nC6GUYkxSCcgYVl39qCYWjp6MAfSL4xQOV/JNs5X9llzJn
xlFKAtB+lSDdMvrACQV9YtwGubYsQ6tE0OCwLOme/ImhLAePRqXnB+7gwYrWekfsSK0WQleBhaDP
k+5i35nTHIHbxB5k7LobhUZ0m79e/r4QPgEtn7QAaYhnUywq7kTa/QTjkKDih5cQXTUpe8RNIUzs
kvBU/zQfV3Bqj9TPNM/mi2LF6fQQNCJaklOeyQybuvOqf+dmQ95hpesvFASEnuEhPiM/TScR9T7N
qyfykaTExzhXd4bg1aoDcf4W3kRuLs5g8t+99uN5V4A2bRDXohLqpwv7fKyVS2HggUnqgsdCm7Ti
pT4RMuDhi9pIfOq0rR8+iK2JI70iTOJ33Zo+qlQw0fFGSn72ikW6fc+yRP2gnNqMN1mt4jLA26W+
Q2itpo2zDiGqR4pdu06oh//xWnyJNwtFV0t0DoV0oCwYK5yre2HdkRiExZnp0GiO/9pe0kVQb6/Z
cNZJ4dOR4/tfV6tA4u76VEKhuzavIvPo1GToQHUnO/KO5kEHQ7n0Q5sogWW+qky7/UPlToYT7QF5
SiUzYSCP/L0sSb/OdLVOYWP7CHpZbGGciwT3BdYtvgrM7HUwykC7X6kLRvtewuVeyZT6Oa5h1s65
eb53TmzrjgrA9PnGh2LeNATu1cdOVKh1ruBdETgcfB78pP5ojk5JlnTxrlCVetXUjvvzPybrrneK
mNePH6Mferd1fuqTAOhLwA8nI/SJmQ5oqwLTiF10XBHSIm8yoJBVfzfbrYUrPF69dAetc3LYO4sp
3z3qUxkxk4DJhVSy85CrbITt2aT19SXIcDh9JkmZlQ5K6SuQxEojPdkM2jutkdnRJj8aJ6Zc7Fb2
/mraMjmcIgq8U3Xthrh7XZZSpeaG1acNZ3ylBaiCLXlSwhS2M24ftePpMTedbpJrZALzL57HjNZD
95KUpUfddds3l1ry6kgGPwmPiX1aW9EMw1esnzmoIyYWeNFhThi54kk+HfgnHPc8BYCS1HGkBA3j
6qXNdrrls8eXfaktj7wkRvEoNJX9mzukJgGH838XDp3EaLyt+yXk9HrRReoaQ3AhorclQWnaeH1m
BAi/BOmYFCHiXhieV7eyxnaCMBQtZ9BQT+r65qMefGl5VfdRYQIk8581txIGLtcjRv9Db9p+L+y1
6v60yHtSV/TxGfXS4G11J93RKPMESCiELNc2jpTff/k4xBSCsRgk/t7du69RxK4VXlNZqM6fhhgP
m/sqNs1ho3INdCfK3R8FMwr9m+n88rJJ3p4zXdfdMGgpV/Jn0z7lWOpJusjYHkcTZAKcpTHYqw9H
zvcXS6BlICpwdAuyt436zy1EyjPnbDtc33vwZR0zrQ6C5dxdLemsbeKXS71aaERcoe5QxJKdjNmG
nGCbByQ8oJGxCnenqrmoPOOkqmwRf4F2b8Z42UU36COQVBxsR2eyWra7wu1FmJp7b3Vch/0EnHCU
P0/svfMGYTttyRIy9fDF2fuhUaOV/UgVg/9l7Sge1H7e7pq45qGUQ5Vrx7oI3zDxhjjN7Gvgao6y
Ozy8L5AoBg1v5mdE+aXPOynZPnwM4aBiri7h+gv1orKO+zDKt/R2lZAWAOHdDwxEjVc7EiCCW3Y4
zvKtgVigP6epR+OzvjCe1E2wMJQi0C6w9vMQeUxBegHT/dGiGIxIYB7aVI6mXh8R+blTEtKr7Pi3
2vZYDGpgWtjnBWhOqbfIsHXGhNJVm3zZ1e4bJFPO+qCodI/OKKcQrozoePlauLRDk5BhwAqERY3e
NjEL/bMqgtQ9aTxlKPk3IzM+mxNuX5STw362n0ClFB4Noto0pEY7nDRLawTeIu1ocijuPtAAua7i
xkGIn2D1sM8aNxmanZHadgJGcRHMSR4ekdhP3iRgbEuDYWNhsF06U5gkxDzeSNww1Blmdr0fC7t4
zLdhnuT+ufikRWkiNMLJI4fKK+4ll/RxZ0NVMjaUoINK4LMVMTrVtI3UbOaitXri/FGaoTPGMXjY
nB9R0jODqN8mUc/G8UeJsEZxtughTjyXXleuOw5WVmx45FcnBYBiasyK5qnj7EOSfvcJ+yEeQEYq
bX6yNukAzLmosZbvzEwy7dFpIwr3ECDAiAslogMJcFE4nK9ZG3Ib5sbiZSoFwxvGllCBqAR3eIjm
dyhvnvtnFI0BVxvAhbYD8IhmmMYnuOCjRDUPl1fL3ljUHKdhSI8Ju/RU5syPKlVMBvT2DrWV0BFx
fUMLcX6OmWS4QeMdwNJbCfTyXY4qJrtKGs7WpIfA0yIqLDSbQ2cfdVs9YzAuvIRVbHox1awlriwN
BEOiAhGa/OUJ18uYPrgolkEdoepWHz+2HlY5dDzamQKtMYYD/mNcTCV3MAiNWhypj2N4H1e65COz
oueIDVaZwDv+eVSQkz8O46V8nN3eCiGNjQauqyHhsfXAWaeY7mJDcfYhq+zOryJTTSe2EyyNiQYR
/4hqEltoWvFMXBDMee4QUWslJ2vJ+2xcyZZ4TKQmokauD2e73Iqfyt66V0wxP6t/jxY15DtpYyLH
Nu1c4Nvl9Vbp7RUTu2WtFMiVd0BmQVPju/GoE7JZPNxMrXZQ463s4eMTSjYcu/aCsC53QQLWuZnn
MELUjCEo07at3EKOgGN0BbnsCxkT4BIbINDVKzUL81w7EappZOcfHdP2CyzycsH9FVOoaToVbRTu
a5hi+8s3bOG8GN46ksqGHLAwRceg/g+WNxaStgctwPeaK9A8fG7bEYdmKbckjJUn+WCYh4MvXe3o
CMnf9n19kGxZCW3fQgbKZciNzi9/FGpWZstUtzyl2x7PJ6ZcN1bxvo82SiKPbrcLVbiuFBCe8jbr
Prok3CAnUhsMMhwfaiTKMZtx8GojQHhPdtkbhlBd8QFuiGsHFGFwgQ/uqE7tsFopwBzOAlcI9Ac8
EXeSohicdDSREvJ+bKVODs6mZC+xy2eiHJL9TAsKgslLTa/RDWVB6Bo3KeFonU18VfLioV9BF/Kf
wnWioOpr0BzyHTx02PUqe1dAbIM7bg6kryu+T+usCZXg4PWI5+ON0xtpPqvQxYa4gMtOA9W10MMJ
vKsr6mQkl/2O49WHZE8m00qjYEvb1HshScnktWQV+Ze3ot+eGIR5IxyqgF1aSwbs8ZsUfxydV4YL
GQSqzrbVwGMSdLALgVo8IPx4E4EGomv0c6Y1kPpyo/skQ2yPjlVn17QHmOBFy9jHw+mE5F9qgI3U
Qxhr42D9TXUE+h7A0yIB/U2Hg/W1GnjhYVCdbK9YbgLmkgtoSHINZkTPs9SHyktTixmiZxAj0hGa
eQCBVGJdyyL13mb21yOPsiJovtQsYLcyriaTQDlmIUwu4ZNBnY3zrnc/69qzJOBo0y9xB+f2o8KE
B7rhIPYcYFSE57Byd6XUcTSm9m2rJHipRcgwZYwwS3VpwQLpjQ1FUSQqAz5WvDrnM0VINP5/zdac
Tfnwfmji5rAu2MRgvb0/p+Q5skXecS+etE88NJtoZgHOUcwd+xOsRkWlMztsXRwmmdLoK27qEAcU
RBRdwjSTP+xxp5qDxYqswK+C9TMUMD9Aj8e7sCf0x0m19YRcEBzo7Fnzfuo6OCluCcZHwTs15WGe
fKo0Vaqz3gYUMstxuV/4FYmwz8gqXirjFn3CF7RMjaiFWM7RS58u50Cok6hyWzFgxLQ4ibbtKIt6
PGoDp2B7RhxyuS2+AysT84XnaDofCwfEUjYB9K7FcbOjkgUNoWjFA06+p9TU+SCQYN6Ur+I79gKP
7tcICyuMLGqbMXvwDKD1cqoABTQfltYRS/k8vYWdb5iHfja4tKpcL7NlrC1eoONApDtzq/IEWk3b
N3G7R3A/GzPFt+9y0xrVlvhItroivKKHq/XWuIMbql76/3ZWnEVI942j7YvCBOcnDicQMOXl+4J9
V6Mv1mgAgLHlqPSCLV29G5sThwpbtZjeFENJTRkmJEjSk/HbtMoJhm6dB4I9DoCmxLJnfXZ7NOTk
W62iIZxYAqwbUG0YyrxfL+AL6dVQEtNs3v31czrOwaRgR6f3MofZM5jY1mqgO6ExnD+kimUcX+V9
eVPlJAnwaKcrQIUaHxVbv1DErgqIi0OSak11TvhBY3YP7Em9HLBPoOygCbsjq/eU9P1ChcaYnoXC
+OqPUgV4C1GA84MtdxLNEDiNS+aoXh6uaIiVUdW6v/ryF6buD/iqO4O8CyaWtFwxvOR5NGy+zH5n
4Y7B3ZedhuKO+fJkUtHYaPQxjb2jBUuA317ZPa8rUaWRSGOM85PaH45pFa1WHmXVhPwR5lsaiqCO
uT23RXtmwT4hNUVI6r1nNzvksQ0BvfrXEZlJj0IbIaf3iJkbzXqV1zm6SUqiIhd4CSbl6zhj2zb1
IxAmtNpc293I4zv/euWpwi+ew9HUvOH+pIBzYtNigVOb5jZAHTM+K11UQQn063CdcIZRTLqtIc4y
gGcK7x/G7orV9y3ksFknXcreT4iyxH5sdNBB3CEbFlMLjFcqr6BZY265iMR/RFvwAHJYUj0DeN2r
C8BoObtwTd4x3SmFzXuMJ9xdFFcyJydqstNHFj9HF6jDPXJOpyAIcshW1yn3784EHexVPS0WmOlW
I2y0mD1CIH6o4ZpS2cu8yj8caKqAUpWYOn05Kd01uaGrz5LsUOMjXs2Lxp5Lq61YbhE+/dwXGKxQ
KPPNtZZjnt6/7fRZGYhAp5K0QIOLpzuwYJCkd9J3YJFGuOLd+0n2wzq+hAZUqWObviSCo1sFXVq0
4NJLq8Tme9GVP81PTAQmRdMlfXJ6onmJoJzl1qmi4dzTXEBmDO+EHucSVNlSWro8hzzrz9XTKSKq
ACG183Hzm0NtglDx6EfYiZZdN2wwQ1rxp/8CAoQuQSDYZZU3IeB8l9wPVNZ9IALEMhxHO2tHQaju
yvhdRzwxUp4as4VQWFFvc+bdcjwF24cO63wee6cLRuZCFNf95x/fLfadq6DlyBsf3cS+svIde0OH
beDLkkB7xgu4WP1HHNmOqm5Z9XsKbQGa8vcsDVuhgUeTjNrsNiFmARxSZCsrFvBtyyGS+RDg7Zon
YsJ4TqN7fBqfQbppajvJLxgNP6mpXgC6Qeb3wQq7lmdH/ggkHWNvwF8cXqCj4sM5RyCY5JX7j9XU
JfOcdkmqb3LBd4uQLD+Lo9CifyQmidrTF0UEp5oo44LVGF62Co24vsgTqwBEp9YHHG9aVyV3PTbA
9sd+uEDFrfH8Zmobw6uRPw3NY2cexBbnflV3ATdntaKVbM+O8mU9jN52ykDj7qKvI9gW3lVB7Ey5
8Otk4avNJdA9s9TXL8kVr10mtakryHJEBQrEMeEvWWQl3Q6xRVkZ58JIFzUZNce8f2ZRCQlyKgXD
x13N1PLu9HYvcCvx6PevpTiuqLwEYKvPXkrWND/mu+EJl43ZsuNckVILZaHSK/ArkCVjfzsEaRV4
ZiNwQVd0KlXN17NtP/S+JafCzjPcoE712K6Rhq83tZ2BNaSh6YFQoVjUolag3fPZGs8clJksmeGv
fn27q2zO42nnzzBb52yd3exhc/Ba/nFoBhhYmR+vjgQKbM4oK3/yGtHka2sU2iXKLv1gz5GahI4R
chE9JfGGX5PKAMg8/gBBdLKOzyAPzcfiJZVRZBpnhsjzNhHANfRvuao3Qs60FBAr4lOlZkjAfCQg
mi355ZuSUAca1m9XCoXtBE22XPgLCzAem5Vtp/W/X5uI6bxWZJSqw4+DgKi+C3XLxIcPAFzlmiyj
DysvK4NPX0AHmJxokl7asKkoDK1pLVcaTlGXHMLSZjvbDbMQjSya9DW6BUSrXj+aNbNx12YDRdgg
a+qESpIcb6y31UiFttmgb+JTctmQRlKvTy1QJ6xpclrNulkCmo668F98tSeHVbpTKDQbydN/BFDm
RWHam+3DCwKCacjEkeADWXtdfAb6ybtfmJRiCCfSKveTZl0JyizUW0YLIKIjK+PT3bz0U8Q2pelU
X6tIk2TqmZHje/yeNtFAbqDlClgTwz5A0z8WVsNtKTmvt1wnAxt8ZW6p7WUU6jbkhw0rLX9C4C07
JP1VTCx3+/uFKatMgNgcD0ao8+igcbpS1j2mKrSrki5U6YQX2SFgazFKo7iPfRvGSX3MQsFwHr7p
+xmDz3ifc5NHoPcWhMVZjvKniASGP7cfqeou5FRssRDmY3g6kZDtGjJAd+7wY7pTD7ELQGvVip4Q
S+EbhvnoSirnNU6enmzDZnNfTsh6e/yFDs4/7uxn9722q4mggTuXnXX3hrmHyoCrvkD27HlSFXNf
v268O/WLk0pPLlvK7hBIqOIzCMOCjFdSVSjpvLBeFnRwr1fmfqVTGWFSvTV0nIp2rGjd57PLQZQu
ETIOylnWolFYuN0jbr3r84bTFak/j9aqHBIYUe+ZBp3II31/A/ajeVyTf8M7GphJBHAXlFYwVzdX
MTHjAKR7UiJ7AxBEGJnlSMc+sipUG0/AwaCvuYvLE9s44t6rMfc4gQ9nYq4x30mYu/+50LEwUwVi
K2qq8uu/OmrmYUhxhY52q+daNR55U6bUMNXEoahLxwOAV+ZBo3PSmhEsubi97/gjQit69ZD78Loc
cWou3awPmLDwHmOdLmAMl4zeUPNyb5rFHUf5lShp1xRVsWjUpXxpSW3dhov+ff2FDepj1QtonzkT
XZp+XsIaqe77T0ZAw9v2q+W1/LBOBoAYzZ2b6a5GluRsRn65zUC5CwjT5sp2zGWKJDLtdaxw8ZqU
NJWMFmormBwuIGDkqcmGPYoUIrFJT0rvxBjPxRhQAHv/Mgam3iXBNKm8u/CdySNPFiYaVXtw6Avb
f4fEUDCK0mJzMMJxEKgSXonI+ds96au8/dn725ZEJ+0jPhtvRSQVROtTYaq1z2Exw42rjEuqjxyS
lIE5L3OODRyVPiygLj+U7VLLbvuhs92DB8kf6771Z2+Kx0y7kGkxu7FE6TxU3wkCF1bVhp4pc8+9
2fPQaJWocZV2PlmqiDQL4BqrAytSBobvSfxjsbHgKPP2Xo7rdu4d8rHtxfLeclGIw/xvL8eSVk4b
MkrU+ipf/a3I3sxs/QZeWjjvUfSztD2l3SsPnQ/mysDEchN9V2zxOPv4ArBN5hx1pKBHt/1YQqPa
1ehnVMPC5a+PkkCErTlNWYvX4cnAAgeAy6tFV48sOSD9n/9aPe+dIPWmBAXT6Nu2x+5vfBFvssfn
AAq0YVuwHcDwTLPQ3Nqoqi+H5Y3aCOob363xxP5K/9yQeESCtwbc637EXDBwrq7jgTZ/IPhu6B+i
Mquq37aDRZeR8MPcffuGvON6xadrshHMxOKjs3Z5TeGITO43pqosPzo8mmZ71vDTl+RtTq4drkCn
DiwSMVrMgP4SRNp/M+c1l+otwrx+2lUi7zkf8gMXfXqR5/phw86oDKS/+suQ47Zznw8p4KTsIzx2
pWjmzKJzOdl0UWpFssNjeCoHLnEHfv+nanEHTKX03uhp4Z0MAq3Z5k/zcNa/KUsKKbs54PhKvOvM
1JyKG3NNKxbwRs3cIdb/vGCkaXhSXHm+WPktf0/0vBnJUIe+9WvR3OworiWK9V2oXNRHT7vnGDro
67wuQRqwIzPy6TJU/R7k0kNfvUmpjLQh6z9XPQ8SHQQNt592z3Gl1N0czVxEkg6ZbJJltQcKpYnE
0qjjatyC4z2oGusUDFRYkMa/lWif/3kAK1I9eHCfI3qj1F38FznttSZopS4ksTbom46h83ckF0wz
ARusTwaDsMgVoCxPqi7sYjKmkceewU9jdQ8LuzWQVKOw63VqLOqQELgDyAhtXD5t/r80TZlsOnwB
3lODSizG7UrqOgTNtQOCf6y4mggPV4HV3+GXDdJtWleP9KIbOvMXOkTUiETQNoGUyVc6rUyWky4b
d9vRgsrwpTmwZ7bcrBMBW9+qxvkTJ+EuZPPM0dDHczvF2J7D7JYBxx+7ycJeBElGhsZrdpJsdxJ7
7H6mukdAFeHx7YuQyq+vqtS6dRFAfVM/RDWFQPSrIzoHJVb6t9mYrQhQ0TXTxCEougbDXQ1/FZis
e9MYD/CzSIc0k10/8OqVfKCW6iDosOUZz0FZrPZPxUA+yhhsVWZlI04Wgh6Y3h/bnFb1w6jEduXp
VWK9IjykrU9V563Hm8AfxX0OT0YqtryOgNOQm9OSMYoTAu8LcT7p0S0R3ZmsGJKAKK1SxvkHJJsO
dnEMeM2zId2HjfgC1PjiT6A7UFvYfQc1kx7O9O20IVIJeLwCUkiy8H4HFCGeRv94crzSVwG7mA2f
gfd3+Qs9Z3cOfeinDLFvIW+oZZwLznnG43Dx0iEitug88/AXKg3daZzGqMZKRR9Q0xLltSU9M1sw
bztmeUIy4wYSWUqtdB8ia7xbHLtceKsGho6dg8QRFmEdImSdHbs16Ygq9XRcahaYEq2O7nABQ6IB
XXnjXLKDmRDTgPVc19fJzpswIW+1tJ0dIYsSQFiEmMQEMMnuOfW+DuNWoml4s8WvwaRZe+AfFtsM
d3xmGBOHbe+tq3RtSoLJfKrrPvttQeesNSO70dzZdv9aQgJAAEvdqyertRxmVTXlij7WX6hhdcQi
4lXSjOmeghGBeBelZpODuKHMJ7z3T6nu1VtqOo+QO/qfUM/p07yZmFtw/oZMuO33jlz1i5Y3AbFz
LcUhkRgw7cyZ+h+N1CgjDkv2U35odo6powLUBoLkO0QI5ZnUaxNi4pIgH606HRlaSuG9Bt3pfIdj
+3NDg0NqmRpdMlyBD0LQ8GVDgIc44GcCe2Dwg/bieyuAy2ZAgPT4hmWuXfmagc+c4uZv0AS6085Y
sbGswwn1e6JfamimlmRy2O6lsr0VTJ8HKEi3crsnsB09OiHM/bDaWZ+mTTOQ9BSjzWjyWpd5Y+c9
P2MvHa4g2gp1buElaiqoQv0y5ry+CD68MnGRG5KuBFF1xclN5KLXr5SUT9r9PIPcNhklhrMBORPe
uQZ6zMify7dJvPO0vyHtxLP49pCc7atOynk5xEytrekv85msQP/nJ2OgReaC8P/UKCuSutmYnTp4
AmHFuPfX7iDxd5ogzCgRVtLdXWnJlHMVsVKyYNVPExfDqsBsXDz66Nk0NdHOtTKc+3Z9tnyOts5Y
w4y3ruNIYN5HzuNHVQtUo1bE32igIU5ae3AMxnbCB5uFp5Qopr/WopKPgnIgEoBgZH4NV5kny+My
9gnQQtHrTnH9osVSGsP+xYlW52d6PoHmT0pGIdvgPVioZ89Kc5cEj5OvaDLez50u6sDntE5JwXWi
jSPmeEDuKg9UVGerjmbvuDbRO5ECqsZj96pE1DoB3VDXhfFge+5v1x/aIICs9zQyD5OraFjnS69+
/JNQczRPZypff106rv4hHlvZ5uwExVg+Jus0Jiv2EA8iyniMdE6p7BsrNT+s4Jfror66JDLQgaft
HB0IDzJAvJ0LpOyBctAph9Gsx9aap3ViB8WuEjc/jprXcnqHCUNYtwV2WTVol5ugyzEDCrPyEBlv
S6Q5/YwqmB5rm5NcUkp+c0+QFR5xk/yziaLKeftRDY4G/BUvinB+AxhpPW0knKZ2By1QZc1oFh62
fxCGu9/1idA2im3Oo8puZrLb0PppVZ3DvD2n5q8Yh653FBg2JhYNZvdvne+J+EkUZ3H0xivUpq0Z
UL+UjY0KgRqilcRYwWxHEhPtx8+APKifo6cM0+khA5fEpRDdTZNyVIYeMjo7PmkMfg1Q9ANgmtmZ
rG2HQj05rk537HB9FAtt+74GBOxHJ+/cq2wHrCQmpGtUxx9qdfQZcfU1Q9Slcij4HipxNOZc+/4r
o42jStffjBuDCiW+bA5pfKaXbJmA6o0ClCqGRWfEQ2XXELf9g3TBKx3zcUJguGriIrlDjtCfmX7l
dzE+42qPfRWXlaCrI6RDOm06Voz7GEyIHq8vWKV4PoUDrM65p4jhNr3HdU061XSh7Du6H/3I9V2+
ska3n5/jdjVaYp7KPpmbkvsIpcQK3u+CIOplXRC/0io8iEHtI+tM/6lMQ0Rfd3MYe14Y8rA5/mjm
JaWPKPBR4KazarjoWkfKf8PU17zyfZn6ogrXKMNQLk5D8fDKlf9Gmnv9bDBEJQZHGE+wMrMvkfBT
NBJmqbYsCuR3MbnunzNG8blOLMT2PSYskjU8ZC4bJS8I0Gl3MHpl/RWJ1wIsicup5vVLbQfSF5Vk
bC9SiaUjA2hzqbrGFyC27uGoWlTpPAVp5xPanlPF1AnO/W+K6x3N1MHM+PcEVx+LkoUPutOLeuAu
CXYUnB2P6S1Litvy8K0xd+hn2FdE2EemBUUX7uGdFDLqpCnO9WgsEOw+Y+dkSan+5uJdMSVBWFvm
aK24AnTwZUOAjNqB133vsOMGoGNVZIuOJqK0js/EcwfXgz5OQJgqnqR3DkA2omVyVLDDhAFAGXN2
VrkrWvuBQY3Djviuve7AV+e/fxwvtjkgkq44bpW6pzOAaYBd8TylIIzWYuDKqPVQyOHn7cT4txsw
hxJIGj0oo2yOjvYpGgS6CPqSBZIRar5ITlrMKRoKvf/I8wyONTEMDysEB8kSGeEigOSz5h0GyqfT
UF58Db6OJVYRiYrGLZ/r2mKhj3C9qGqgGuUWyWuomUi6jZZ95dLuHRF2UL8S+xSfe3S0W9Q2VwJO
lh8q3Yyw/EGmU+cIS1iZzw+VnOarQ2B9HTr8JFXkcqpYrcBZBAniwskMm0tlGMmiOtp9L9gC323A
bOIS0aEJr+I3fnBuDF/Db776uBtbHUseRItWRhnOe574vuB9EfNPVl7BwQvxYU8nSIfZztfgs6Ue
KZ1+5nrlFSnhytQdaLE+kSgxp4u63er4ih8JBIVnvhvbU/ect3zwoaI2EmkkqlGfiENsbsaYQOmE
5SRtfWzHYTv0ipLxCY8X6CZtO05DW3P3GI8j1NlEUKLefONPSkJUC4grA8eJJh//mI9hijwX2AGM
BqdN0cjsdM4YMWnhKKGCtzfiXkYGrZXynd9FEZluo2H9qZiuduYdQkp1+FpYxfuXvEaL71m+WdwR
XVSNDYmIluQ1e25cA9UqoHaUlV05vJhGU0fCGkAXBPBsMig1SSz5ukRNRxdYspbTTKoT92CZU483
w+mGOu8L+iaLPMJZ94/u9YFT7UhWPthqcGcEXXvcLstcEIjuT6WpLeqQJU/hprjoDcPLXhMFo1UX
QbgivCMJi6noPzATKjBwwdMV/igUT0FTQGj7+Vq+9AVLLjTYJxnVK0lLMg7PHhKAy59ZPob54asu
zTOyABzVISzlTObnRi8Z0WXBBUgvMRfz+FvxE4LG2+Y71Z6Vi9M8WfyQ4o+X8CMydzzsURJ9vEDH
BY55QqewXCTlK3wvAmiwx8qt5bmOiSxw5obNBtNAja8lEjuAEMTQQyRj3ZGDPYIORupX2+NwF8Mo
D21Q2cif94JidkQAL0D7CYvZmUL+tqh5tdLDfMSXF+VprF++1ObzvXU9qMRkUpcbv9NXqKaZVsIC
QZ8wEygZKmtn2pc69SHQnEFZ9i0FcY9IV52idVSysSreS8YYMK3s4CzyRLCvSfEZyAFvCURKPlhz
Ntw774gVIPEgMM6k3y487GXBwAI14yqolJwtWnzp8tSYdnVszk1dUpwXEPleP3/ouEjXcJsPEhrX
mjegCjJRRIlUoEYsfvwGDD9ceSJjUopSQanWVhhvTAeGtyFkjng0qoqJ/gI0kF5SYa+XrV6KAr83
orem9DfNU4XL1wf6gtOd2CU+4wKGIGs2nONuS73RHn/KlZMqdj5OCvULpAl2f2xU6JjLKT96xecR
3JjThC1Hoy0C10s+R3DgNFMLSHdF8DDL6XCXfvp1ula5wELn+/CnEp3l7sFgp5N8UxY4ME2w4BRb
vy2F70BtJTSQVQOBuIdUb+ZKsRHbsIzNo/3OgzMEwHitCMwv1O0MjvtjOIPVST7d3HsIvqx9Cn9z
UlsJ9CuPWn4rn/vDBPhXowo0r9RnLUGl/FVdviZsgAfHb9YIHKhVf7/6NLeUEHFvAGrJZuxvJHo1
DAG2QbOalmddJz5kEPrIoETrdwNzPWlmtsiBXOOJ+g9Jp5RFZ3ujGRKKsbpvECdjCmghcD9+e4AJ
fwbfQwTzC5kjPLz/8RSFQai6qh/aiwpQpkD2Ogi+vCRoJhPJu0w++SpkhwdY2dTWpgHyIVuFU7j2
2QPzf3hH7SxU34/lGfpzdVBX2+KtfzRaG0S98CFbsndMoipRPOa384ouGKkE2tfRwrboHQ1GPqMr
FfG271EJuSB8YZTDDwjFZftMAdVlpDo+E7w9Q6nqbYQ4KthCKN4wsVbT4zOqwzxfdZy8VfL+rG6Y
GhDDmfWDjEaFEBpyHT7Xhb7usXph1jGxdOB/NUQTAjHzXGToCQXT644E9xv3kXF1hOGs+N+wnT2g
KWtRAeDFcEAt5eZDj1Dhpx6dIvS1Cmy6wSeFB1NkMvK7cKYZVLALVOCye62d5JXZRy617dqYO5NN
5FK+1SA0pXI60sGdnlUHkgJRZ26VWNSN1z89Q7PcBKe/jrtqt7Kw73MDDovAc/NI/CZm9Ye0lSdx
4sKe+yfuqFD9OuxEsrktY7/2eXl9TJz7T0nuKV7t76022EHJvabMUwKodMsPX5GuXqDM3NZ2KnTy
sFx9RgbSWerMF0A6RKe9vLwHqsP4dG9Ci+rVp6inn+5419cjTXZt6q3QnUFm4cBIDN8FHTB2UrQ2
zMEYiBVRRWg6EMoudURz9QjjHU4njydBbDVWiWHziAMjPC/LP5vtjaKYyCoAEw9B3//aiOEsFBmr
2GJWjetvitiGrRwwGrYcLTl2wkv6sS0cLLaa1NWok65rHDgk+oh+kwyH3KcjCDXXmOrivdxsXDAM
RHa2J/IlQBC1+vj80Ln4Xg3YVLUhm/uFPHlY/bB5AjIycdK7kBDM+r8tlpsu0Revob8yLl2sFQsH
d2yC2V0VsUw1Zl9d2JM0ez2GQDoXqH/dpYgtRrPxFeIdlVz70pX4onA6Z6WaWRRt/sNo3bT2tz5s
nV8/jRgaNyPsfHRpo4xquhrf5sAj65CIg/bbcEugIK4C+aOwxkXi4tPm/EhJAn12lGQl3t+18J2Q
H9pXxqyxv0jZYR7qDTVP9fqZxr7wCz+qzH08jVzAuspFB1+mZlCpGoIGed1wYelXqIvXxOGkM64d
SqkqRUNNYYMPlte+3I9hLHdGf2DmBaEkiIrOdJBYHByQMhAU/XLZIgI6+cNSWlLKpPp4a9eWrsM3
0mw24sE1WF1BbTQZIgpicJfnrzPCiRCUg93bTYcDanJwS8sol+sY1eiG3gdeXZA0yZvu5C3B7SYy
AKeyyKGZFic+IGHPO0e8brWWwiAw0sfTvsFXwjFru2U6wXgbIHFWrbfLM5dlDx9PlBpozSRC4Q85
Rr9MIGfwBWuStfWUoM1KQnn4Mhxz1rsNoTUTNHuH9F6EMh7MfhkWv7xgdPEiTMRSCIAAB7KohNKI
eJcmN61JOuxtClP9HCVIAFjz4gMpeInbxv/rR9RniWtC9ymRs7bcPkH+Bx5vAdLXaEsZGYTDok/q
uuHcJ/pv+DPz2NSXg8AusScRySNMAnvtzXBSXGtaQ4kCYDCpnTqVIjGvIX5JUuyTK16XEpigmk46
CaI9U5cPZz+9Bhm7a4eponn8X0GFM49j1DndIRoeqaSjo5yXj+242VoySszol5RyM5/J00z1Ij8T
6HQR/XpsqbXJqIId8jM9nRQMpCgGX6KKb5jc0CuPQg/1uZ/WqLmNRq/OsyTimNtqf63h/L4ennFA
yCZ8KfWdC4VBhnfiWLMgZaDUT220VPpwEc9EA1SPcUDfRzimKjlog0+ED33ntIpZw7WshCHnGebL
aO4tz9S9GzIQOk3+/RjwGCqQm1/MZ3koZhYYfKrESE3DSL1LeAN8ex/phMr9H7ZVGeXijZgKLEH7
977uWCjbL5qKl2zw2WGr0mbETlbKD/VRpAuF495dooTsVAnZ+IaDYa7qTBU8Gr295dOqhZ+17mpm
Cw2bLtB9KDp6o5pgEpuwpQphjyhCH1iLgHhRHUHunQHkoth+45BMNRavZUve55vqFaX7kBtKF3/f
ZE6TFRV/7Ms6b06nb8m+9lw/7Kzqo3nmHaCtkQNQnCKjSL6sv0KDDw9OUcuyQnLx+5J2sgSH9VlE
eqU/iQaBHNrQD06lfQIA2r0NwnWo4UP/J4fehy79yUdBzggSGl1v+PcsogTV+odqmiivOAzJasFw
b8q7LkWyuCNwveN3vvVxch2ibta7ETXqQij2jgr2wStfKA18+D8VYa1Ln3BofuhQ65PN4OkeJ8k0
HHbxP+7zUkw5FiTs08yb9QvtGgwyUZzrFRBpRlDq1n4d6KRD/wijiMJaR4Afo7SXc6VSYxmeoyEk
584Yes+UlWvLXsd3V9nkFZmPvcO3qOUSuD68lZws98UNH8bGcJaIcPepRngUWAN7KVI/PTZfo/Mu
oRtode0Yoiq/qbFK0YOQlOAkiyhGbGq1p+oz7eu6+JQ0cI34w6OKXTIsMabsZr3MYdxDWBrNR7C2
8U5LzAglyEWuGrIrcsldHd/1A7FMow6DKQUAzIe8X0JZ92eKnsxBYcNu1GA1n+gbozEWKexEGjzp
Ro5zWOeR1stf3EhKtrBIHaTfjUQXaTh2AEFkdKAMiDw0cxV+QP4MbgwfuVdP7F6Ind0kEtuGUU59
9G0hjyCIpMTw2yGbGfFuGV6usN/dLVnKIbYcRgoK7qH7NmrzOlzPQdfh9wKmZUwqvfd8awYu9h6w
8p7kPJxX8D3lZdy6/RkaJ6l7H27UDw9D4+6eKCk03sCJSB5OhoPdOXYBynS/EVZfuEw0joBGNoWu
30DD4r57C5BDHhNIyjEhs24lgg9QTAsIzS7qfEvbFosKHGs5sIR6HUj/vujH7BYlNHfn0DihrZ0q
/mlNs10heO9b3K4Yj2BmkuGsX933aizMXv/9gUvcFFo1pu6by1ppJbWNNg/aGudwBTCeRmOOPnPU
9wBalPBcskvUzcV8zGQXSgJZ2C6c2uy6UcWxLfV6pdZ6zoGLwxeAL2VBVXtdJU5hKaSKloJvVB+u
Y2+wy51r0AdohGYOlFevjflvZorEOw1EgffMJSNeuRIBPKzfPOTeBppuxn6MVYAcq4QssZq8iUdf
LJ5iQvo6LxANOs4lJKA9HuMg9IryYPTMc+wyODWJNItD6ETlsUKS+V6y6zwZAh/G5LVHyQ9qTijS
NJ09XuKqcl/Qirh0E4XgbpJovnV+WWYKdaXqKN1udg/gYyu6aB80LS8yNcBV55wZJsMuwVs3nh8B
5keDqdaRA1L51U1HDwVKXMP+ob2VL6Jaj6pLuYlVNXZZxVFzIQiVI9ftX1cjPAwGimVCE2j3yoRf
iTex667DO5P87DA4UweqFsR+A7K5RwD07bCpz1Wg88ygY1EBL0WndgqaA7KZV6Nte0G7royNJ9J8
CL7Bwtg5MJ7uz3uL+TdD42lZzNEqCyMnrHrjLx0YvXIjKgy3Li8BLduCiN/3+pvWdHibGhcZovEY
ElegItMrprECzl/S19nadPmgHYuerYwVl+VZ8ZcKFellH5cr/RnQiJF1RdMGp+m8WGEGv/S4XZ0x
trVaIwQDQ5OguAaslQ1YwUW3L+oVNudZP7J365lSyho9bGLcb5HmbJWMO142kAvXHvSD1Jpkyvr2
L2B4JfgIZMQtYVtQbnh5VX1byV1oif0qwXvGW0U50pqNTzcUSu2Oz1b4DpJZqTXpeaX1sgbJ0ZCp
UxoZmxtKcfZuxuiYYc/GYzObYtyKH7e+mB0gi0BnfZBkZu9bIUZnx9lOicfyyl0kb7PugsmLrM/u
LVcUCXwAULdUg4SChFNSE//5hRT26+az39cSwseQrJvnYkMftc7IsqO34vUajMkmyKXOECW2ovMx
ISgi7vivy+781I9cYVixu4A/trTi0VgNq+gyCqyeoMIQCK61Iq7upo/9ahFSory5laCXTBUwcHg7
5Jl11kbWJ/qe292NDlpOd15HJHST6OXU+XETebKt4GE+Mv1Ly2qFTS/sWmgdCO7X+tXCApXFUw9I
yMUQz675nxNbKat27Cdjx2jV8oPlU/eNkztoh+on+KO2oH3b2ahmbMsjkwbUL3cKd/RPb+hHGpEC
GJtaOLl1gwgyklLaBPD0DzXb12H1c91oakRMhVkjXTgUDfsKEo4kxMzY/3NqNWDZoLcvZxHHIGb1
kFTb36tsphF/fuMNZY32F3+VUrhbbPy1CJzpA+AqesuxWrMHNdglA5grAuQuyo7D9+O+rwq76x4I
tBTgdlbW4NWYa+6m7oXR14HlIfE+hMhJk5FZzEi9i7dI6RfImVDutB6hzhngQph8ZLl6lGEZVT5Y
4sMm7FG1MVEM2XO/7rUwIlrDaPuiqknzh+ocUhMeee9rJMUB7Zo5/v13yUbX+30MoyAV6ZykrJ9M
dIgLEakdhc+53IcdCmQLFhaxZPuZgtuigimzyyaC3nrT1ja6I/H76vmcXJ2S4+qJ64pcST+aItiT
yMzu0CKjXAmZlW5KyV1CIMP12nZJkhvQCTdOjFbRQ3KZYD/rtyP1KHgqs0lsmCL5nuCpTPNVVFgp
SFgCJ6LO+p0ZY6Hs7EjfzHVZpwo1mi7Y/cLaIr1VETg5oEoJxulcjq2meJ1D37DryKOKGLAIxH9i
0pfhyCe8jcIRDkVKQ2KxojKF/vfEjJXRWNpVOIW7+oi3nMqXSc3ADkEOK0X/pK/POka0fCIMFGMd
uNZa7zCrFQMGW4EPrTuqWo5dMAaR7CwtaqA71ShWGYhoDedksUqQFFQpSvL193IFl6qbMEFRrFxn
ixqBxGnvL5u1D4TWApuCwijQSJi3SNP7KzLQtRmYIt/q65Dn1Y5qlTItLvMgT5Jabf4UtwkcYRBF
//Qbapz6ycSHFy0DM3WREQaOy664Pb5a0Kd3u6BiPDLT1SKrKpI58kBRrAgBZ4LpfHUzjIxGqKLg
zI3kRBXc4VO3KYqAiYj8UlP5TBFVZfLfAp9cIr5xJtbhNNezg+mFEx3SRg9Tew1i3//wIOiF7915
uJoXIAFu9m7GeCf12TtyesAJyt9ODLywIvAhrsRNi3VzCusdm7uNEojS3wEAvG2bDXRZKmatXUKD
jLhQfyfMkIXZdmZ6BOuSHJSAEdKQLQYa1jLY+c08LIJJXi1YcX8wfnXIdPkZmslwwbUtMKbeSsK+
qZttK/YeInqi4rq9RKlHrmigyf8p9IRLfZOvjQE/HfHG4LQSmAfaNUgxhvz/lc1E0MRO6BqBUAqp
sFRDl6o5FaIt5rk1UTgpYie8fDa9/GX4TyGFZWLEaJ1QmYBT/yN29Xx7+FxH6L58MyTQ3SFeXzjo
7VGpokxpGG4gCw5rI78TFE0G/X/l6ISwALeFRv/HLCnlhb81oTaERvfAyYebs1q6vAtURPlvzPqb
RlB44Q9JsV5ZYmNQd6EJWLDjc8DNejIsVx5Yv3vDUiSNNyagicjgXKuv2mPmxA6sUYNbb3NR1J+7
lgRD2hzx7a32DGL7oKAEqee6+LbPKD5lsaEo42ZQhzpglDJMW65YCFdM7zYk65Tqo1yvF2QHJnLd
pT2imttXLUvd6/DSV3esNLxJj3RZ0zLMPmGGANOOoB6UEhPzL41xTABLaDoM6D3N5g5CWngkOIfh
htUm7GMFftX9wB0ElQpSWwW73EQpQqrFbPT3xGLhvnru0NuUeztl+7vg3wXo/Prl6IdJw4zZ6PwF
qB71tkLseEJlZWQLVogtLNHvgdgXbyA3jGMdSVV36pHYWbR2oHuYAOPXB3jmX0mE79LGOilOzeW9
UJx9BgyZkXVbNuTs2gFVnq25sbwPBZFvXz/r/Fwy+Lc2ldzwUe4JLOJB1hBAEgsu+gzX5J66qZ4e
DzuZdvSYqbcGthMuIXyg95N/JzA+vm+ZuSIm7c447Q4H4tg53prElZ/HlboA7poiDEFVCu0f4pyI
CKa/ZliV6Y21PV72DmIlpJNRygoCsR9b+QhO0wtp7QoU/XgjLMwGl6N9fiilPs/+hNULIrv2rb8T
9I5W0OgGhPOSVhJVTASMuGg59ehSfDKHghAb6F0gTZ5MMZQy3qsBzWy3rleji7hb6k3f1p3fKNDz
hYmdPeGYJ+hGAEW2m1gvS1icdYRZdEdYOig2e3Kr0j2+H9xpyEbsB/qxzAKA/r1Q7hTmaFY5V5xU
8A3faIhnXtSqYOKw3bWXdsE7NC85ZgMwkduOnf/UM81Mfk/vTAuvn/kpzsuGsSqpF59p6mD7JTvX
9NlO5uxuoJJNTSR19Hxwd+DKA+e60hgNh6XndZFG0ye/20N9jcySw31j6x0UoocaO9vB1wAne3xO
VwvHBwBww8SygFW27BtGSSXaETY61cgLREfoNT6EaYfWAD2wYa7UnVd0nHjMCJh+80bfx5BeNn7F
+bB74xj3cQ7w4cj1cvOtRF/Y7cL+V+Dx2wAx6gvORSYmai0DHt0t8dGe6INqUtB7sEiBESDz98Z7
k80fJjSbGvYqk/Hm+hitqCmIHx156Y4WBG71tm8ILELZjIqHc3+168CzrYsB/JIOEDJcMmpeBo0k
oXOzDB3QBZlNPVR1IK49JvnxPY/HnxvgK6K6RDVS/62lMnw53Xk1/QNSp2tV5cwzQS+vyLvgacc0
jJ9Cn5ar0IPaX+cOExM+k0ZamGIIa/Q7GFYxPbFlxhZlOIwUodY7zvKX1itvr4Ni69XI2SU/Hja+
oqv7gJ8xxs0Tot2hUvCQ3MkaDlWSgxyMnxiDqzHtCxV9AmTrxM9Ek6VdICx/gdc7pCfX50IhH55P
RNDX29vdwM3QMIjsNrfRG6tPe460Hv/DDDyL1B+tJhK5KjB7GN2fIHtQC6uA0kt8p6BZ+hQhx+Js
O0G8WZ4cYz2luHKwgoScLtfIzdxOrDvc7+k84rZHSfvA0vQwCI7eCuleddq1Qd4PUxxAMVTviqrC
6L1eW+ZtUfUETdcTIKRPsmbryLm+vjH7S/wmBt1yzPAH4aTdnoGrpV4OWEHSNtd+FnKtBf5tgmKs
77uNCv1NshfoCEtKQS4/jsbGWJVQvi5Aw+14dWJAowUhvCaiSAQVSV5vlMY8Kaxjg5zHJbDUGLnG
gy7XLKHtnEx4GPC9gzkSdyBujRwdztzCqqvaqaH4nuIyWQEGyYzRQrH+HalPkGL3gYO3hMWLfV9u
e7naFwPPInWReSc2tsoiiI7szsUSx7NRsMwo9Mx48f3QKZ39nCDTRe0HS1zyMaDv7ouc0AAg2Tw6
iEx2kcbkHwmkfn0n+fgwn/AWAUL0TApvpSJ9759GPjyNeTnH8ae+zkXwAracSIzBcPWBqKvAxLQT
DFDTf8AAMd+n6U6iT1Bgfboielsjr4iCMXrhJGu98J17lw7DU6LAGL/z0p/Yx6NPL8HohHFD4IC/
VVATvA2vxPNmTYft0K/Qiw1SjbGfsw05m56E/Gzh8bFdaEn2UaOZchUiSvdsIjEb9EEOEXhCY2tC
r/dbxscGDGuaZrSLNjOOsjPZr1ZHrU/2RyKO3JbBeh3knD3TWmhUwRsPlo8AYz4FSxEtprpjLH4K
PXCh/hyBI3ldagYyBUs3JXEck8ibifPm1sCKXAvZCj7zjqLvVdSCHsWpeOZ7iwHWsJlYLYD92iuK
EWAwnRjbhRqSvAyRnUcD2OEAmaz2jpUyuGPHagirmlzyvfUoqN1mv+XcjiMfxar2SxorUfB4Dd1v
+QHcTT7V66UGF5AxT/OmvrQum5PaynufDQKTYLOSvJJRWp6ghKdqUdwLQR36eQqc0nulrLjukRTv
wn3qq2OfQmrr/jj0wWrK4xxNpu87cfZ2uU+IplsiEaq9ILfYAUslabrQp1+tBj2J/vkThpKgwtml
rIYBOHL1p2Jcy2KSCOcYx9idBFAZGU59KIU9DMF0isTOQGMGsvQ+77s+VlXnMi7Cuf27J+90D/F1
zR25viocinbEiPkXHyhnAWprmLc2xkHIfEp90TUjvLKUJpNnjlCFutQaDD8A/I/MXNNAEVZ1dEW4
o77vWcJFD+8LojGFRHJEuDwZ4fJC8lLT0SQ0uDw8QH08/FDdSHBphbHoTDq8YY5H+uceQcYJEoeP
UFtjFu1jvQJoGuoSItRvfEdTIMP76YrWwc0HgfEsDoWH9DTvTCiKNvoNplNEIRp0ElthDD6VtptA
hFact40A8Q9daFTnvRw/4DvidMXPN+mBt6kRBdV0DH+wQv15wBXAEz43ZxV45eITMl0pnVtpkpjl
Bh2IRyG3sfeNvfh2FzGDZ9phVRkeyHZMloAbPAXGc9PrjsvRm8KGAS+OnloocYozgAo46H+SP+gC
8OscRh1YiYXjJZA0jfyxCG0wil8wnCXpxM7lxLqidzVeFOlJl90vJmfPQr0ld2a2mAGHLn3yFMvE
kuuEbbWWWPEroDl2yUinyJj3lYgzLLq2S5MCXjdG/dN4MBFxYsHSs7lfodNqh4X6UrVbfyRqN+iS
SVMFsi0LU7NrcMb3vnemXmTHd9HDJSjacTwvpqpvm9kL037KZt3ULojUdzl01FaXEWL/2N8NvXVa
lFm2h+pwKOSBYNHR8m3gIzpYp+8K6tQ0JM4sMJ7+Oc9kADG4fC2Ih0jgpolhyNBdHeoJqa/1uUeH
bFY8dLz9RUfVHXBGsvVtXuqAI0d9/ZN9GiF4kXzU7do7TfKPSTCV0fRtuUXa2yXnlL3x/S+ZI3lg
oYFmgB6+SwQ0T3ke1RKUPJUSqQKOeAdoC0PjS6v/lCN938QH3Lf4ul999CxcZ8m5xrnYNmCqTw8D
YxIlwdYmFLSD35WhzVmvxSZqIWS+urqrzbOHbsazSi1z/Z1FLGogpybUp5K0YHzMKUeIyBfIsxsK
6tuYqf2xPJxX3IOh12LI/H4ohuScyNlVbsxLAFhiTuXtedIn0b2R7UIpQ8q1JhP4hu9tR1r1x3+n
Fbwexg5a0I0NmCMURDU9vP4BmiKQ2ohz8CVze6h3cqaypR8QoHGEGyxcOunVh9nX2J4zcnuxGRMB
aUvoNor77gkH8bFKjdY/hYV5LU58URMFwYrettkxxpLVZz0m+dhD/4Q/vw/QwY+0liluBEPDpG05
TpatzfdYHOluuJBoWFh4w576uOJXPNh4/AZ62Ev2XyyZRJuZ27Wu1csT/q1kEGQuH250/foUr/KO
xvptpaLwBmFpmUi0mPEdDVyHN2PclQXlPjoMIu13FKfmvPkN30HegTJcDXYrLvJUlPM60SBb0mGe
nbHsyTMF2FZ7L3hgKbANvJzDLHxBPcL+P9hMJkF4q0gU6Hb43R9099ZV0DW4bnSENjbhIIT1SaYu
F45mkDK3/AU0mHT6gxcin0CHPYyEUXWdS32a5vlzlkGamcR5SoX9KyQbhgXTs/s1ABK0Samwk3J1
Sd3C65lAqkMMEgn0wZNvExgzvGVaC6HEd5PuwUGPFIWeTmRME1RwTgRuZFhlaUwmJF/Y4UeMc2cZ
tCZpCiVckibu8TdItQrW7LcJ7WoLcyqoG6gLqJ+rOsKXwEONOaLbEhuItMJeGEwqMaCHJooH2dnM
xc0ulNqf+drzbCSyzZfqyBGvNLjpUJNXSgyASOYBzxb+J/txh2kh+Rg4vdpv8OydphqFEDjxTNP0
qd2eA4t1JoqRrI2YD+umVt48VVQKbTK1eaKjqiH9D+2et2bywkse5e2DkmOS3T83BpSxtx6QFLxo
CLgmVQOVE8+socc8D3H8OEjjMaRVcax66enAhO2f0UdQPsF1/LHKZge+ci09kcwDKyFxqPASCb2c
k4BUaZsHxoiLCoPeIZW1Q4owiV7feBscVJYlfK0+ykrzBCgsIWt/3MquIVsa1FT6Gc/gCoK4kHHa
CsSV5H1zt7qZJrceH9LpyPWWvppOyO2dgrnTyIZIcadVcuBKyZXUNlc1VKZkSali6oWcgmXoGA1C
hhRx7G0yxz66Mnfrb8nMz62Ay94wVMlLuWyyElDHmKTcXptWGV+waGo1ivS8n43RuDnHERRyieuf
815rpK1F76OaZKxj69BAGYp/JAbHmp5UH8hEEyQmFwS1RTgaZD/nWwzybi7xQ+C5yWTdJ6bbNsP6
xjHUHdk8VA4p5L83nJ8TqMvj9hEVvNn0ateorboTBBM68lH+4Rs6hug/ZeZG/DNfL/d4M6c3cwBE
VvUvte8BE7BxiQ1MF/NNoHPOLnyo9jqAA/qL5O2RXweZgFM1XyIMOu1L1pm1nKIeoqHrb5894vyN
iEl6TuK7RVb9F8owaXTgQOIlUvk9t46xRIK9ijM+RP1u3KrrEYCTGFtM++HLHlaEfteMk6T1BcUW
8WDgFDAmpVpCggmFsjDaVviwqCLvqkZTvlRLZwf7IfKMQqAeWoCkeI0WtZkNUEQ/qbQQYbqToggW
a6743NIlJw50pUIYKgf6B8k+40GKnT/8Ghb8DfXClbyIgZdosm8uwPOtLKjxK7NvOAvCGD5bqwF5
QdEXdUKfe3b9643iXkBmOJ2a3bsvcWbPpFqtpq5YELGuT08L+cqF6V2jOH3BN/tvV57Rh+ElTJQH
pmpisHWXt0lx9/IP3YrYKPp+7Zfd9Y2xSXHnbw+K9OnyyPh8raSzAH+jyoiAsg5pzLuY0Wq8+mqp
HV5TUdMJ2ypBchVqC0nYuKOV32sykYLHZBFdBBAeuoTkZRKkuWPbj4OAc8zLZx7M59STYx/lijkI
MF8DFxFfb0RNoGnISI/83rUjwtNXv9cjGOGCuOnlsZSzMOXGGuhuCXiNKDRlacDYfFIUJEow1/Zo
I3NlL1tj6NMHSwL+XCZHyBwfgWosuv6jMfdpwrpiaOaCLeg16gGc69IcMOpZSx6FxfenaWjjjg9l
qSyHi0aGJgc0RM3vgQo6mMpGALHvpJHaCqwFiDjuTQyNVMp0ZXyNwHKrkaG7i6r/w5rLRSCpmInz
qc/PIzHWuIxpIL3bMlBdT19XSnVX0SwrOx7ybi2UO49UpdX4OwNPNzBFux4QYQXoBE/4t/3RSPCU
Z/tNtlgLH9qpu8n4vdmaXdDLof6K4/PWpCQTwWkwr3BfOEk+UVGwdOCTLo6c0RpM5CW4n4YCozKX
aCZ6svf9vl7fqDVGcVeEf2qCsqobq8z9uEYVmJGZYwOCiflT0nQ9rONYPpKc57ap15gptAtZDiAR
g0s//w3tndIZRRlVYnuf+YCIvMO5uCpkQwGusy1YmiBhIUVBLPYVRkx07siu38qOKM91jJbFsG5a
nH6evvG1m0tVBvSgllcpKiNI1VNMcW+dC14B2kQOHv95jlbfpQt2tFCNtfTYYRj3/DjtZU2tuGF5
tWk8pw7TME4UTXk2Z2OB3jk/AUHWiI6lJVJKVFEc9AzktJJt4Lp548m0t9p6VX687Y0WLXCQoSx8
cAWvF17v/ceM4y1VXEMvGPZC4kTo5nY1MZxmIOQkDDlb8xDDwIfgTqk4CLWRySCNrrKz4LT+o/pZ
oykldICcCIFD4I0wkT+WGEScA70O6uCdixraxtNBtmsvNExZjdVrHpza1bCOkoqliM0BQBxdNnf5
ceV+IHMf2Toui9f+Eu1Lg/WXcZ+ayKeZFQw6SEeILwYGswnwxiSKhla3edNypsOUW2nPr6BW+n26
wuIDVkJEPT1N0lymH6YGRgAk0Wq8JOuxb+NxcmtdaBk0CKh6QmapInCqlmb1tADPiIjqgkXkKUAN
gMQa5/au9uZtMxQw8d/P9HZN0FKsqYElhqOYq4MWoEmYJiNzViBnV1MC2cP9OOrpoHOVlYbOskfI
QKmctxPUmwROaF6WGmxHIvukq2uakpq3+cKkV0emoJ0tMQJ/9NlwAB1Q7hL7gd/QCKEY0O2MeevT
ojzfeUdfQ1QEY8RyyMlrFkCk108KooV8FbPvNHANtG5gU4lUpR6zpzdZhGXNjlJD1nQzqmJiLM3E
utxdsQAn4UdaPXkqGIO6L1B0TThXFPLOyjENfGQ/qpdFBmrKPpF9SvovXhl7YiGi552UWYMv3hXF
ETgivwR+ayukvJdkKqN0K4xAP7+Q5oEORN4AdqTgk6wyumDhSkRKE6PXlhC8JDsOD59jvfv3qR5v
YC8+0+uNLzqfv0HnBJt+7KoqFO4x7mmSetIOtqhsh8hbDkx1DjOKrrBnjXi9vbwBwxPzPNAVJecK
yrZW65TPIBWHpDUzz30P7EL5DO5uv+3xtQxR1tefuLdtQQJJw5Jaq/KDiFblO/yueMV1tUUGpimw
IOprrOUpkV/542YaJopOIV6INxFrr6h063QB+AlhtMuhQ90dbo1fr5ZbY/ILoX+HmUJO+EvyQNaR
TtUmowphec46CMglRFzhXUl89Ynu8a0Vos/nP9xeDYUT12WS7UaLFSD5thFG80NgyCmFgGenc665
y3JHHzcfQ/38VqaXyoXVWLhi9V2tpia6zzxh2gRWHHkc26lzxFLfRfdb4Tbf3X0rSNHpPm9WGxW1
y5/OLAGf3bFdrqu99Euu2+pRHB/E7zri625tCqp7n8KEPClk0dUT1uLVY4X8M8MyW6Ut/vHRFqCX
JAIKaRD96rTUDX0dRx3I9K4QNkj59M1Cc6rP/6mOMrx8C3LX0La5yWUveXSajEn+nrXPOuJfz7HR
JsstDDOnhmDQpE4XJuAGZKwDXDPFqhO+cZ1R8H6Q37g4X6NlwjD0lSbX1mKE+6VTZOx3lkIDIdXp
8Ju7xA+26nrkQ0U2LQvGFWlAUEk2f8VhxCsk50qZBNibQFXi1+ksGzMjbBWrM3EUdwYRtDAPPGqa
QZvj5+LHOTSWCiMbLO+dnmw9QAakIorIxWxUALq/B6VyRIHDonGN976s6JMaEGn0B+ia+HDRArW/
ysnD1iq530TYD74BFIwgchgsyH7uO0Lnu+J8GT8gnXA+5++NS9NNBM+MGU/Q6LaIgOaDN0jWm6V8
SUF+Um4BVUegWuqld2An4opzBA8GfmYrgeEdqA2FdiaOTAgcxCmdNcNDmg7X3Ic9yA46vnR2KVoa
i45Qvxsb978rlzRtG/G6IH1/NNFVOja+JsT6QQRm6+njpJCZOM/WCjYdOYqy3+zarOFMszqIyn9B
WAH6B+I3bs4Sg8z2BDH8JN+mk0T000MP/i2cmyT2i9C3IVVR4VPuMtPzSb3WNh8miANUSZTiQ0Gu
EB3hrQxSDLbkmWQrKFaKNoJu5qKU1+Ka4whwiIw/gsiBn9kcEbV/Z63x623MtHjUgVnUjDpY2li+
dqqei3n0/lizmqEP96s2xB7uK2KYJoJ8+2cFU0wP089Np6ct4Po1XCM/9wUsqsKu5S4FAI2CDzCs
ZbVQq9iD1Of65cf8yx3/+9FT5Q9O2HSbNsQXYIlx4LcWBZscSv6VQm5M7VaW73ZFK+K9P1umXqrR
crcoVeAWGIp+gpBa9wwr+WmE/NeSOBVBVlYdQv94Tz76JbVZ2XVzYuEMtyMu7cbgS04wFDxE6l+O
WD7sZyrwpydrsC1l/cnFHlknLrClmuSwEk429Z9v+sfp+OjnsWUkemNJSEDgNV1mnM2FD39t1uBu
hLSiLUpMNoZ3yj+zxSt4gGG+lXpzcQQxvCAsJ2roRtFEq2LrU6KInjUdxp/DyfA/gpMPjhkCBIsP
D5qNBizm+i/ToK1C9J/QlwcaMzyEcQb1OEiBXByNjeqRbMHHYaCQitbCrdzy42xgRmVzDKYAWBUf
CApJ3sNaHFBY8rCQs0gQ8w5rpcrSBVJTkjStNrz4gZS7fj47jxannH0yWfCoz+fXIlzkZ1T1++jg
AEuEW7PkZq7neLSKcerFrr/u6USLmc1HXkraq1xBOXMsiFSUGMr3rv76rMWPkK9qQKDsVnvMkHAX
nD4G0uQZhUwh9H2ovr4LZpq0ZB7HevhPCMs27/wkxhNQgnekrm0F6rQW4kmD0pHrAn6e/ZcWsOAc
Vk2MQUklPVMDerGgl80/vzInJ2v40qsNneTPbQSlWaHnmMLFINe5Xwysg/V892lRnYz0SLxwTqrt
OvE4ytGOCjVi0+ElLbNvPXot8jc4DgQa3+FBPOZFWZ1XPUe6TWI3cLyrbcJcJac7Jmbaq3EJQQyQ
buEmT/HJNi/g2JAGWgGw+bI3yE1oVFjub0Xutomo8cuH8UoI2nm+sTNXXyMsZG/y28EgUJftohMi
BQLfKiXYxmA35OT5YUZv+DD+66yvu+jrBPul7r+DDCsMgZSGx8PO2/M1i+LIW6o0gT8gpOc2bkJz
9zawiV3M5iGtT6SquX441zIqRbgkZ/M+kglUssOMC6EBCpibhF8m1RPBRC0bpMsFH+KbyT8xdIhe
68nUnOYX8llyYRdE3pu3AUwWZEEyWRAJHOrgVT0TKHD4itsbVH9R2pMxk5DXFSGDerIocvs70rZ0
jahvkGhOyuwHnBPTk7VV5ow20SB8rOhOQTmFs0Sd70qtqSk1PT0KAUSfW7UuXxh4+006UHIP/PgB
zjN7y+2Wolli6rn3OiRmedoyCc7MJ6Y5aHmZ+7qxntnO5XA1QvSUGtCP10o11FibAM7m68kL8T7W
VciTLBV6PKWR5a2lHsEP7Ygu61GANK+kdRCyZEilVlSfv4wOlrGi9vCqW/6ToKUFwMPN010n+JRd
xvj20uHMsZ2kGv0QPrK7iQvMvdmU0KWADV4iYTk/ojJ6N5k9l5XL2EaXJwog+6Jg4EFBNfqCzD5A
mArbBf1QZCEJVL+XBA6S+uRePCuCb59LSH5K6iss1WkpocEJhw76BqIbzH/A4ZGcwokS54gDGg0R
6oqevsWdqTi1MYcyXIWfiab634AfLlhqK+SKDa50Hyig8FguCSwNTbaZ6K0dIalBPto0BTYVybpm
Ed1N/HUxJrlx+JuYUwWlvlca6f/JUmqb271xhplo5+8BfVBPd0XwhnT0DZ592tR0Pfke0WoZNm40
kl9qhLcMD1NW0AHQtukT86D5juCRxKpnfBhuWkp2+5dGGjLH5zhV5gqXgDKH0XcZwllBEMg2E4HY
gVNEiBRCXGvFDd3GLhAGUU4UR7MghcyBfVJwgOh7AcPlarcHNK0Szn3l3B6ddPwWkAAPySlQ+Dj4
573rfZ3/L9WiUsQDBw8lz/Q8KKoHafAlhLw7A+w/Ez1a/iDIMpPwtHOM1lOT1zfvaVwePHEOFVTM
OJVIfH4T8z2mF5VT8fuXj68wgmMhQkkRXSPF252oKWZJmh3sJOo+4sNTjp9KbAC/B9qQ9GGFoRul
Fk7NTVBZBqc/t/7mAeznlOghShmney99R9PAL9UOd1QaHu0tix/+/zNfxcnU0Zr7cH2cM7r5GuA3
f6o3L4PmXu9eHqU0+evMoNiu7EyaAX5S74KGC986BmSFFdjgXR2ZGEzOj3IY1daVfToQ4IRIuyBk
4cT6pp332b08S+N9R+MCrX8QcYnc7EXOdwv8CbJFNicLLRRBmRElg+nDK4kNrHDZV86BGollGZeG
e2Q7a810SIwFLYMqfGIoI0rM69TGpimqdUMm7IhjqI2XwEqxKL309+0eYRxjDadDqjzGgBvqHI4m
dkr6vwMuP8ZAifRCTQQmxDzW9Q6luY+H8IAZekvfm2LkJxR1X9dBdxLWSLJKqmqPA2pxDj6PIkIJ
kBIkaFRHqECTYUXFO+9OZ7su6gQQzrI1LvyHfj0ZF5hNGdJuIy+D7NUeQNBdyNQZbOlP4ggG/3zF
4gr5kbVLE233+zHpMf3qAYX5deRD6VO4fqzBFxMUVnyjVJXJ25rroqEmb4Qyvl+ZX4fqTqKQGueL
DpNWHg6ni6aExjKtGvR/d3N/k2iXNxZOpGD3nEWY6OZ1gEC1vN56s9TvlFnnS8e08XyZsRRfr20g
vxEHFZz8rd/D+VEcJefQzckVioAWUMMBCIMXtMVP+Aira7myX2p5LxlEIo7mFyFn+WfLX+KhFGxv
z+emx5UEf8kHq0kqwQoUvwC7TSmPdhq2rsFYk2CDSrvH4yqkfoIygaRYT0j80eF1gKqXk+Hqr2Yi
/HZKEjikEcXfcQkqKPOXg0Lhdq+NA/eNHgPZ4zWm0wPrX40jr/oiaxCEJ+Yt42hXH8F2kBt/e300
88FwOquiTeyxzX9slPNbY3FylG8wZwxK6btEU3Lm+XCGCgpK72jESrYQXWQHX7CsrlXAmY9i+PQZ
t/70gAIaoYzbI3TKrapxFlXqGm0eqlxxZhhWYX4M2LDI403VC3uV936McIEuKOgk6Y9G2q/IMXic
j9w002AhPBuRRro5qhO+kTX3SDO49PCPYw9ObpASO1iRI4CfsL71rpqmdtOEvbVdJuGZ7u6qTrjV
k5sx/wlQHLlWj4m0b/yVWAjBgvE3CoPr5C9G+eV/Za2Hq87pg9GA+0w0QF0XCzKAhpcCZmPe2zYt
oEbqhNFwah4OQc5Pv28bqMn/ETj/+/k89iHvpCWdsTkGzvvuslP22R6tvD1MoWi1POH7RaUKq8eo
vqGUO/CppARm01u/7UiW+lM6PR4D0vJ2d+guwHxj66tFbW+dpXwsQEWXlIL+bvQIA00f0Pc3sRSj
+lP5XRtiqHbwv76IgVcbMdheQ7SAzkjg0u8lNuo8ep2bF+/LEN4Qn+1utmJkJCoPCuxYXwyoqiBN
zhVuUqzx7Ey6QEoFxu8VyzYdA173/p6F7LaoWCuB2zDvZ2GNbmq3NHYMEn5zErnvEqXan5D00WdE
cMm3btd57kvsNuyJv3V72spmpdnTj7FKXGP+iNmnesL8By+8HX/lq2YLrpdyawnP4Q2T+9Gts060
FjhgIyoEj1B3hqkg5CqGx3YdMH3h8Fk4+WBJEMRSMoihWCy+O9obHs1uS9ntt23tjS+1HPvGktH2
1442kLzfDGc0oYC9nMr58HwSo1JjsP4B8pm5jtmvEJxHeaMLHXtAw7GWCKX+l1UmeYObls2fTPUe
pAMaLEH3AhZ6VROi4mkC8xJERwony181jT8sRc0MkJmw3fI6jyoGVAhOeDLhGL/113NG9S6D0GvE
9bLSdpYbX/SVGPdRLcNboGk6PIAucARt78FYzn4Tqqy2uOfJeQuESAEvgL3FtKxstJ1Pb/f1ScFw
jsHvqzVyV8YmqwdZMaCK7etCZ+Ce17EtC8JbDx2649qLnzbCk2Pgz+nvFCp2pTS9yZ2fhVDW9Te+
WQbjoIq3ujADJtZU6Dic0XrfckbcUzCI1/Gjo0u82j/IXUF6fGp03Rpc+/klFa4Q5jyTcP3oywuu
iVsr5ceauOCRfWPrINyH7xfKDaM1q16+UvfP1/0/ZNGRiNXBsGAT8WJipBPhKGqfIkdl/EBx5mWJ
Jb5ZejHyRpjvDYoJEn1oNRM89obKT06y4OYUjLk2yDmqVVSPYmsHf+aC8Xj6eouyPT21BBUeLgkh
jlyYAceLahni/WOiJ4XVaagVzZxQJAm353ySZHVu4UffF/SznXsvJAvMzyBib+UsMU602duka11g
rowhpJq80klg4vQ+w4BaWmuIuG5jNkyuClvdfeITmr1S4/vNsqmcmm+gAqTLb4pKaRI+ETu3vrcy
WYBA5s9qraGVSbBbsOn8z6gQzYNCcXWTkXw39LFOSw1Bd6uQsFZLSe95WdwooEPEB+HL58DPainc
H+fVKTZTMesOit9i+rGyjekF6wssfxjfo2zdMfU85thQ8/6kfNDvExLZ1QgjuGuZGKoVjSlTJOEp
vzoMUcaClJ/7tAskxwsq/N3T62/+uX3dQrOVSTeuQBqlV4UiOBlAVusW821gRNqBiXuED8mdLc3U
v1NGU9MlR+95uuHT3osi5iteG2aCvW2AQalyHLdmYcp/N9ogJ84MQG4x4KjLOpVwxJwOjT50pChs
D/YffnjBt3auYB4YfV+Pc0+a5B/pcCdkGXBr+CUlnhQjbjPODsj9bxgqCxOP5S6VyB7Tmdmx+lFu
gu8BhoajbnrtTOmgSbmzgciZ4luxRdBkApccr4zZGA6obHnSdgoFuGdJJwEC4OmM6aw7Y+AsMxYY
kuTqoIeMbPBxgM2953ks+JnXmfRH49nRg+qGggiT4tzBvybIq9v5elJHYjcSX+f0P9rGj9379sJY
AdnEEgC3Zg2nJdXYVO2s+AW7r/SFxI5SsBbo1ketV0GS5HteCEO6JZpHPty6LMsyA9XF/8IaOL6+
8WAbUkTx5LW6IZx9Jgl/siCfZLLhlGmdE48ex+IA/OIbIjsFW7Oo/YupErsVS/VD6Nm4m1+4m+CS
0PcHWugsfWFANNih6wsNraDzRMpL3ta318Kn5+j/HV/WMW7sWC1QN4NYLViyJZv3kNtmSim8N8qK
EtGjDAXoQI5DdlgTc8bHpe0RNLY/fRyNGh12SqFQ3uacrXjFwcTzurLv8BArhD03QeAtex6G2+5w
xNFynOKaT/IVSj916K3EiTMq31EqQR244Gioh9yHr8cycbeGBjvqEi2ZS3pxTu44bwWEUERgLODS
I18XstBq5F8Cex4iQPDv5XCKLbjKTG26R13LHCV5IJWl5TqoY6ZEOTTKqMcGEAvjfO43r46KCBAv
rjIM+zQUTfk9aa6dZYC9axQG9cF21Oc+S8LJl7KBGjvJ5n/p7P31zP4QhdaoG6R5GQCCbyiiszoj
3csboT68Xx3n7f+UMBjxPjTz4J6HaYeuLPma1M0OY0iB8qUDd7vVruHwOBwjVqYP+Iiyy+lgT484
06pu0pUGttVokQeSKmhTlUrFMx7kfqecr5vmUlVRn3uGm6KB8ZWtnrLNn07YGm67jk3WEQYIjtP+
vWducuSFNflqNIEyR6o/2Gj4Qs3Jz83yupXWuZaRS+4xnIZNhOtQ0FXQ0DdzippWHU8XF2uAUigH
piYmEvSW823b8SyVCOcPPAvOBR7xjiJ6MXreVfVJxE8WHZOWES0tYslqkWQo06WdlrmVdmBOZ3Vy
38WeQXorw2xbYDBaWCpjX7biI+goNBV/e0yoapEt6rHbJ0Zmcr46WdUQgHbY8Xgf2WeDdxd8Ng41
A1hpQDjNzEe0ko6ctWZ6ePa3MDr1YGY+3mQ+TtAQ2u4EW/+1CoQ4+1Fc49YZaPx/2DzRdYR7+M4l
REAQeYpVE+XJyEppdTRQynr0lWkSeUe6XYJhzX/RlgCE1e2ulsOqNabKD4ybPZ4Rwvti8P/pzFJk
2qoBiJUuKYfj7VRd4tJvNqf2n+CGsgI0LPdQ0QUC2GV3FrZHkGSOy3yzaJt/sakqyDduEyhr2gu4
puAAWtm7ZVHhwDAJao5Z50a9Nq4nukOv5fSNNz4mu2AB0khh3N3uslDbGVO5PGhWWmDEBXiHFn4g
vn/n47k4ZzLdkW4NB5LE2IfROiGiInI4WxiTHYy0KjYC/u3b6xsGNWWCYzxwlIAw6jPHkY1eZgw9
CFHBM94HsAVKc6cbiEi+jWmSbEVqaEHiYunBcD7+yLf4Flr5pTxFh968xSigCAGcYH1pZ0oLbbzU
g+bfpRBr7nMsBciehpRWcFYwwTq52N10fLeOtJgiQMIY/KluMSVKUfr6OB12RM5ICPolpQj4+vdO
I8i9pSsd7Wn/E1QkcouYzFG/pVgzWiMSqkIiF5wRnd0G1Bz27gdc6lGSeFMhzNGJFsx2JqPFqDfu
R6QPYf8ewm7Ksc63JkdBBTNcoO27rILhNI4ULH8xjJ/udMc+9rW7rXtp+/sqEeTHXAMdGY82bTBO
mRCk8wzVuLKfwZXuAEFyJZsykqgIsu90GJcqh/lMTpF3TGVAkVUvIh15qiXMPKCHi0NGiWcg9Fnl
M1FsnWLMOeOatzMH2AS3hHPVPUi0H4DK5jeBAnqBPVyKn/pHjaDgv0I/dziTkfMambnIsae2YKl4
kq4pjrmKR9552bHzPrnWcz1QsFUQp2z0cdER+lZ5qwhRaJD25dWcLT7V73HpB0CXVQEVme+6IBks
a74uZ1UKgpR1UVEXnPGmGPFWOP1H6bdgFRMDF3fmbrHx0EFRoQdgo1FAC+gVyXiwu6FnpadBvVby
6x2HghmuKsfclr5SU5cI83AwZdkAH9vvmqKcUX7uRpVZWwWvki+DqCtKt6PPhNa6gH4VJPYcyzFl
z3/7H7y1JZnyMSdVXB5KnD/lQ5Ojj9sbNfidBah6B6wQi1kpekGfV9mGv78En070Vv1fjSQKNaG7
w4doqsFmkZGkRNDAsBGwGg2LIbqnUChUFvZffpUvKe+TLek8Vd1yxsizz9O6iamHEw2H4qB+vNRi
JLQFE1rcVr7L+mngxDBqYhzw07aYUDZBJnETla2QST3+Nikqn6HRJ1gvhClILpaHr90YNNb8/CFs
Hx8O2zHrAPx/3yQfmnXumDzUdE9rzZGkcyhpZS7rEiUXTJCmnooroYqYGphDxRJ0O/BtiRX/mufX
KJguZ4/vQJ+96MEmV66NOI/PhfObK5bUWUMmHwVV0Hg2JejAH9G7py8thm0Li4yUUgEd9YpF7lfC
nL4PSiLgG8uo+62RUsYF9yA88XeIcEtacIB6oEP9WWHMUVcjxmA7ZNlqC5l48nDP5riCrJhTFZso
V74eCCea69CR/2biz4tPsAkEDQd9hGh8rATMTqpJXwS3LZyZmT40yYqfuuPUaUGFD7UnkWggZhnc
5wi8YfXP4Av9271ewMjJ1XK1hOji1troIMpvsH75rF+wCYbmB9E7+Y2RKRcad3Fbk4vT17C+31su
X/ppb1dw74QcMagOSMSVUEle3kV2h2W2P7FujRKGeYP7N+hKFfJM4kfM2FIzfWh9UZ6g8GkimNjy
ZGKrHGeOTkeHiGvOSycsYjvkPmu8caMuPDuV3CJK6IbAZIudi88B7LuRybhu/RTEk8nFKTqcluib
EN0oWC3amEmVIGvWiOZ+93ZbiEZcyM2gw0qSLCU8klNs6ff4qCgeT2DhmG8Wo9gdBnI7mtsP1A28
8wvDMgxlTHLhzKd/oYDVDXbTiy5S/wDKr9J7ptwTEujgGX3gtuW+lOTXlyxFao0St/YR12YV6lZ9
g5l6Pkd3jnbL9Eu9/W7eOgXSulE96+fRICGwkCWn73hNBJx416qXfGUX0DPwB4n8MXr2mB8YnfU0
BnpQGkg41ZY+qPAX/irPmo9UVMPHve2Esw2TjTCDw8ZQZYu2fyTCi4LTw4NMh9R6Fq5kBfY0pBXk
00b0s3LrTv28ZOZ5ZzUEN2srz7SMybEYXAl6qyYj93b1g14Ds+pFBjP5GYUboFTILZR05ym6lEtp
9+Y6fZWRzCUaYiwPPlZEDrSGs1mO+v/UcDed0+TElZHW15YKbV5V/g6WizoyTttsL/BRnYkpEmzB
+LtKFIweZE7NM3BGWFY/RNnWsyqVSuH1209M5KZOHB2dGok+dINuUYnrBNisMIpz7yi5g7ODnlv7
p0BK4qWQ5Aw+P0ZHCBAaiBY47eqj17mXQRkrk4EO1FUV6qKkP3ZYumvwidRgIKixOHapI1jf0RPu
UJsNPw0qjQRbSkDdGdeeoMssE7Xbs3hVksfbq7GP6n4+lzz9/89JS/11Vo8oiPoBgp7lRnokddDO
HMEhLwF+NZvmxyrQbas6y5S0AVVlyZX0UxsbV53TBhfrUk21vSI5UNWnlCOSn1Iy8t3kDqohCnwO
0c3S7YidSu8Ecr2+zxX8WrFXDzGRADyMAtbIWZd+qND6sw0d+1pKJcCHmC9r8ysYLHXhbmJgtUmy
qoX4uQ6rq0Hi8TVGLGhQiSlLStpqd4CAj/AjKtt97hFmQeWGsmTVzXhkz3VWKo/jOfbkx4gn2bT1
Uctap1tIXtkkJzj02HVCzOHwSwgfBNIluWDCJalec91y6TnD6OuAAe0zhfDHhK2cAAWW4DRkBfuO
6wk9BkTRmQjCtK8niZdZUdRmR57kaRYfj48aRcBKATnHZQbpq9yV7AxLt0hgPUleIlmDvmhfDcZI
QN5ri1fv/jqQIofmSd1jNu4uzv0SWujvjZ7Z4rrpx1tjzMk8Oofkxy4xSGQwe63LveUaeA75K5MT
h+WMvc+gIe+0iu1imj8rOThZ+9Tbsk3j3IWuoCNNVXJ16I1cZnqKezGiXEjMsohqYC6tsfs5jVmK
0Ou336nzWDBhCRfnWVoDg7kfgfnGlAbtA0WxaHmdxstIOVKZaqbYDPrWsDkAcaJ1G4n9b749sDoC
/BLFh1rUBzvvUWTPxQzVpw68X0hanMG5X6Xe7mhZV8U/jZQznvAfqioLUeSEH5d5HBFPgiUZ2AHt
N5EMhE3SVHb46WF4pmBvY0b2jwvpFMmUyrrM50ZpNAb3Ok9VfEBBeEEzudC7MM01DvXmzB0abopM
aqtbDRkrkO1kpf2H9tVI/g+FCUHEZjfW7c5rJPtDCHf44bGU4/2F5xKh+cXC3fRQddNXzj9bob6N
YKwTj7pTrWWHu2bdiEgKFo7iefm4jkMo9CBJVWfabl2zVSqtZ3BRQVgtWwJLv065MLHA5smHXUsY
VA5AR36gCCpcf7cH/sZtkxMh5h9QTNy5HzzL1gqGcXcZMZJJmdmxy9nZU3bK7WrppULXGYkiRZIg
eslWAaEB9xJpmdeIaiIfgzQbN4glh3PnU8kbULoQQzex1EG9YO2un3DG4/Tm/SmtlqWg2teaLeCe
b2TNxt2E+jTIq3iUu6C+o9bxSIXPUAvREME8nW+GxupudbRylWvc/CzR0cCotgcY06QO0KwEuTAd
WaCGxayowxm/gDQ8wa4J0KJCnzswwKOOdiwdOy33EXyEB5OJn9BZH4SN2gVK7Y1jugrcKgIG8+EZ
Ih/lTySglCI/CkuhYQbW6CyHudDMQBI1+Hsa/l7sEvXq/atJThmo4i832mu4HKDd7lq+SsVyYcY6
jcO9Ijg1xWP85tL5QihsBbJESKNxFPwA/fNf+UwzMojBrs40RPBCym3lkPV39sbtZJTsfGJTAaCo
FkY0aOIbacNYkRJClLCoyW1EGB/ImjYDjxgRkSYCfg3q/2H4kturvsgL10exMFsU/whqCqG1Eq/w
69jrJbz6/Nfm96uH+H/kxDHfQvSbw+BGACwTZayyX30QowsHp5sOQTlsNr/lIZo6VesMC6iyBFiH
6cjyP8Pxg82Uni8f2SoEtVE5cZKxbV6P2o70rcBkzlEMhqE3sVERmlAPf2JpImMuEERz4sWSNMAj
SDdHF34gcOaAi0jRmV2azXbl/kFF4cxVM3wyb5FMy5d1DuSeNdBVprMB6BVqmMvHcxIgf/M9XcN+
hqjkebxroXVdDr8+Xw8uVVBJ78wJZL68+U0S0nwn+FSEr9XsXL8nncf/1NicwS78zDqtNqzwKFWS
q+Gi65IZjl7wcVC9T4lbPsmSPx0rzWZw9HRqB9wxcbutYniuOIPXvR+RR2ZLiRcG4+d6mnssIdLW
usYM+xrbCPSlOQVNDQsBGyHZyIztxMwOUzhJKkkpPsyMcFUli1eGg+36hzPTYSM4fDUFVqWgSJ+t
OdQpKTc8KFX3CMqcN64ngk8Df2HC7+7DeaVDHksL89Mv1TQ4Pv9EqweAZXSiE3+JVzD/E4w2oLS1
FYo/x5vdLW+hvOPSfL4M+fFkNRQePca8y4LHcJsBY2RSLamGt7HgyCllVYaSGZmwXmU2Y3sVnwS4
yM/5PfTHAIjZGYDB0aNW2E/AuehlLnA2uUGm5iiirqZWb4OOlIj6i2mTMwOIWV//FVQ8UVPDl6v4
cAWIkcKv4W3zSsbF4UkFCbpRpPzE14l9zKJ2dG4kmHDbLvS8bGXQQ7gQgJSroZomMR2/X3mTHdXg
6vpB3dAMqm2otp6jTCLTvGNM9F9YC4NNY0A1uRcVB5OuGhY6qfY0RCbdwxh9QtNw6+x+ckVgtLr1
2kHd2fPAh2tWN+tUzo7S4sd71R5ww+v81PNuU0uVgzg8F8e8GdsY+osLTQc949yWjDmLBGNi7ZBp
+uVOdvZyaxCsLS8c0E2jp3WupAKlZ8lu4Hq6M5NPuf7kzixLdFh7XWUs6YidIGNhF922Ew5xHBxd
Q2up28D2tBIf46+sLqF3mQA0JOFGBnngLYuApSHHeVWjE84d/IeM8gijyasv3jMoP6Maojv+i7TX
PBlZHYYDroZg553gmqe5apu0y3qI1vGpsykvAryuNsY9DvZxt47TZW2qFbu9gEdoTVcxrLYQoy4E
xjr+K23zP4kl8UH+ChZSASPnzLCFlkcQAwjLTr3uh62vCvYnHMsgAhSrUV1sXlpbeMiVO8kMtg7e
HJ/QP39z5Z0f4u9Rx65P678uFqSMm4zHrjWJp8Yv/KIMJYXtC3HYXd2FbhWxQjNNHLCfzCR22i+p
qkgvmoN70gn4U6wi9sONgrDe9K2dZ3oetBET0ZXCxLFpHApALAIQsxbzzxtuL3qt9XXDCUfDHbGf
+LsJQsCtGm6Jl4LOCKXjWVCNpTNlEP9AnQlinsMV8JQIrmzrshS+Y+x+rL0NieeOGAlmdSiRqner
bGdyg9f97lkMFTg5z7dVyFD6FErxvv/cWD79jpqeRvDUl83qpzVR4VDSlDwUUPGUbDlta+tYQmuc
cN0NBP5Jl4a59OzLndCt+zYtXUgcl5Zw8wC39mOzJlyQ89f5akfphEkCkAipJQ750XlmA4uV1ExL
51xqYmXaASPGJdSMMSq70ToKiUfwlkLUgk/ZTdFYcS3RCBnLYOCb+n2U4BkTN86Ll8JKGkHgY4NB
DZs5OPGDeCcPgQu9Tr44YcdYzNvEZDabVdC5fwf22X4tJJjsv82WBnW110asOkv/9Hm1HWkA3BBj
PtFzV2xjSzPnEqy2YaKGsJUTtezmyP0mHaPcPLN7CzgLQWjKpcS3ZBMzDajRGOppVVd7Ae3um89i
qFvMWxuiVWTMD+v01jk8lkO8+ECGPnP3ARvbS/VvvsdRopMBLM/0cwbZ0oxmDcq37WBtIIaxvQe0
jluy00OWuoEZebWzwrVWZ+/VEB97cANSDh0iCEU1LD24A/HGiCru4cg3fplbOaCcFfg2Tji9BNNv
NABO/y5p2nnGbgZ4RbBKHKcalWnTNCr/1h2TkTIjCIf9gFhlijrWZ2hgkXUOZLs6zCVbZfqXEWQk
SxqNGnThozy2TKeqnGsjdOgtGmS0GLjLitpaT3R3Pb47dwSRZFQnBud5BR8TK3cC3dyOLohjwSn7
jsBPF4q1XSFCfrxQu988LnxiLdlCMlyHIIrT+WYjsceetNyRUKQN6rwl9EEE18KGYj3Issu/cvtu
8qiKn+yyNvPlI6gx97YuDu5Em5I4Ps0mRmysggxfkM/ZSJXjOtT7KSYP7rB8QoVUXpR8IYY3s0S/
3V5+5hkd8BtUEYGIt2GFHNNbDYOmkuvgtl3vi7qpoLEs6WquDM5RDkGS5ukGl2OeBtxiWlOb5ppO
LcvwVQ+Tz6D1wh7jvlaFgryj5R75I63x1nZUNz6RHmjGK9Wq7AFGXJK4GbaGN9k7YSLrGhW3lO16
tlyKUizBfj8Zyf91CWQvekrfZaBu7aRRz/4AYP4ZiqFD5xQJ7cHtD60JlahpfyEhSNG7PIYduVCG
WT9s70aEryu07OBSQTnCC7aDsVLXHaKjHly6oawL6wyHAZQ1DEbUasKDUgKn1+iq9ZDRCp4t1H1R
NSPtc34Cy4Q28TJjnJP80JCxW25pRCP/vU4uTp7ah6NfjItfSBW0LPXarUMxGcOnL1xZO8ByJIHZ
8vHo+B91BORl1+mZKG43D0RsFR9LO+xLcj22plT0tX1JcTsecvzGnOp29itMnRU2B3x8U8MA86tT
MuF0Y3XY38s5ZLy2xY1CTF/0gND1zYDVsclGYkYH31FoHGsVSXzsthxPhFKOijc3gCXMlJ7TSxPS
2EiiwtTvM05VfWgxgxleVVTYwwqIPtk8X94h8TlzKxrqiIUAtvaP2vCH2BmGmgOQxdyu15FfQbhd
rKNgAilwEjMUb4KF7xI9gyZmywa/dh4uAAEnDyZHa9rIp19Dp36aupv44qhQcoJHzM1hGnDC7Is0
s/9SEWEUayj8l6r0vJzR9Z/yn2SMAoD2YwINtWvM2j0qwp9jrGmGR1I+Rg1GVvvErAacztrU4R5P
zhMX5cL2JEAbvfqQGo07/K8C2BBs1bj9J/pdpPexu2cZ+G6UAaWZD/I+RW39OsvfWs3Q7n6fE3ii
hD+bYW98zmlukhsh0/EFKGwZ1rVz8sTABNkNdUFyGpIMrGcD1lLu7tBlKRDlxSK9C2MQtxOJ/ETy
QKCFpWkkadOv0k1bm8bskj7mPiu0WHLNMraRH4kTB0+yGfzRT/SvID8bbzhjDYRkUCkSIQoHpa3t
9C0/YuVbn9mXNgdDvHXi7OzMAD953hMS1NgjR+m2/z86oARmXjhAxOClgmKRAX2jj1PpvWS9spb3
6bcMlep0hICc89SLwD7e7kn9TjTwY0ZGcMLO+lh/10anMYpyqu5wnEvPmmOmPid5z3I+5G5FRw/Z
CeR/RyQfa/RsIVBPxaoJCtFMKAl5TyGwVz00PywsVCqGzibU5fqpIS+5nfNo2hEH6y0pCNc3GCwE
cVTVp+wAn3AQkIyUYLNifSYqgk3urs36RidPh3re2CdvTB+xVLVpvU6WuxQW6x3j2Ke+DBiV7jMp
n55FLcGqHG8Qe24jUOmuazOwLeTUMOb1YMb5ZPbo5DCBQQ/qoPoh71BJRsMgw2EqYjpjR/25kmJm
zVujaY5O7s1s9XKACeLCuhQIHc6kS9V4+eIgJ5jdPPew89uYc0xGoMyGeVJ7CYntsg30B2YHy8Ln
pUx0rkQHxi3vvLoME84n3FHduvDYYF1NIy6QLMCXiZB3TwQV5o5z4wKnyQnMI20R5fqUJYDjJCi3
gdlD+lp2Z6XUrSJIkwTwpybGAut33ILE93LZu3ajnXuqahV7a3Qaa24RsxC1hRvVTPmFaG2yGzgm
24eWV2TNX8tT3YYKIirIxYkSTBlMIGLjA3Eis3n38hS7F+we8UI3qUMDN7Fqx+anw2noPscbYeJl
Bdvt6brkpgHEhDrJoejudIrR7NnQ2Mb6+fDaDjIEySMyKAA8M76PUPAp6y1vcwF4AJZtvdqTBugv
iAmLwYD4gw8q+SJOqd7rGsdMQD1Ko1NNb9HL03Cgd7EiuCny3sU5G8xRnS2ulq1ldZdG/xL3bIGH
oFBNH0yyBLGmArzsXJbrnxnbOREE2IA60u+346zo3pZE/o6y4ho5nDzFO5QAoi+noQEgh96H/gbw
gNMS/NFlLCAmu2th8KCMFFN7ChgC2elzJfzEP/Bykg4L1THP2QSZ+tzKV5c0jlKQuz4oBXb7tTuJ
rEFTYW6Qs85119ZyOsl0PXqrj6Lsk2svIRdUz0tFWVPBEfbk67J1HFreFtCCU4/FIJgeTJsSp4XC
/TNBLExR30OjYBcoeccFHilBFg+NJCj+XDIjcntlFKANRTlXSnHL7D0xU+kpLRyQ5WoynChGrlsz
08yEoF3oCh660YcjWHBwFabL0ZPDvW4yg6Nie5wuF1IZspnRW9CBvd7N/DcAoOA79qnqka4Kb3dq
WuDbM8nu5Wa3gt1j958gtrHzwgFtLwUqE22nPuMfW+Y1kH0sda/F5tTfDwdcuV3U8do31LIuZd4o
MLx5KYa2vVwmPVZKIMRlUTCA98+SRGlnA1+wn8NnIp5MVuO/ajWezh++SKEVVdT4x4sTquNmjGD8
OcHfiQk8afMkjJlgZdyVsW5iVGgzOcq2RNGoUFOq7pOsR0rw10s/pl0as1ZPUHkmTKODbOkGSUSk
IFDhBmlPhK1RzsskJnFVzU1OXru+5V9SGGQjdx/ERotHTHhnTN0JFWDbNGLjjTvEz5iorzQ9OHHd
XEBsI+wcugR4TCKGcDYyCVjHY+V+zu1sFd9szGvWl/YWj+jRZ2dp5M5UR779WQfnQpJoXfejdiFH
y9/AaSAtwiYrBtmTjd1I11fcRClJC0c73vu8inNf5RgP16Jb0BhAY6bCYh4Lmmgv4H9X29+zZZgh
9v/mocOLJrO2cwI4dJHavHKhjaT9S6g/tkhDj3k0vdmKj/B3Y4Hsc+5gcJOCLqoi3SfDB/XlkQav
2+BtBkaTHzr9b/NwY2QL5koEqLNnkH/XTb2o2q2WYS4vesZmt07DxWY6/EWSFTetFem+xlZ/Jf2g
AlJ4ZYsVcAWsT0WUa/CkZ1VrlplYi1dMTog69ncxsDUass+JGR2xVuREcUOHcMUL7zqt3z1p6SRa
VOgYsh1Y6p0mEnQrCseHnLm66NUfS2mSiRCp5WvJOosmBqiyD3GCqKlfKi97PA9YBJrl378CcDCk
tuPalhRVv+KCLf+GMr3pl5/IlchTSsEKUmCQtxl4ESgKxlvrHFppZXaLovMBL3YgvGHSk2Wq+NNH
VWn4fo0ylJZrkaOuKNsg+DYfHG8BkUIy2LdPKWvQLIUq4r2HIsPSWk0CZBsV475b2yyIeoyjgkXL
wmVER60KUTWR+tCinJUwekS13NUtyZjNQ0MEwCUwKWuMue4cfRvJyfA9dyp4O+fvQtY0MC0AfwMb
6hG6qlVhzr+TKKxXAG0JdJy6YOBMfsJ3Zs5ZqhO5N+PYox/M2UbV47coNIOHlgJ5dTGxJ24i/p5n
ZFeirMMY+CNuV5uGGib6evEObEnQLKlXuzfr6Sqost7HAy+TC8oHeUWBy8eIyr4RxuSOc/9KRkiG
Wp3QX3sAD16ZoPDhDsVqd1u9TD8FwpnKzf86eVMzb/846Im5ghA6eNqWQSpun6VsgTzbfvzGga5Q
KGkYilFBf2NscKg4TNEcTqnrjUg3WIl7fgx5r9XJcwaRTg+YbFVvJAx/7ylhDh87wgE6EaJq6ryp
ABTirnK1RLqzQoGuk2/nNmTxHttrbmm1lAaQPnPROLyCTDq4VU5oMdiytSr8OK5VfG7FIdGtHe4N
8Je/Nn07l4XrzlKkVPUen3UCTBSzZZ8GpjPC/4Ml3YNFPcaEhaeCBts0E4MWq5/t9OI6pobZFF85
k5O+Yh68+rLwLmH0fGK32+ZOmoqsKS1G4f+xgBWuhVSH4OAJD5WdSKV8rsXGjLUxFV2tLH5l8m8T
4HKHej82DUl89buXGq0WXFRfmt961/7GKSV7Yk6o8ZSfZGNqCKNNjBVAZq/QO+H5qbOGkzuMJitL
NRVSyfXsZamKHsAQxKet4IK/j6eWbQmyFTEzDjyhfylJDYaFBnR+Io37a+kJxAPhlh1BlEgIocZo
o1kBqiuVSnI6GFp38UlpjnTie2H9pWjh/3pT20KRBUolAtZIStpr+D8Em3764Mct+/mf8eGiITfm
I7hesNsMrxhyf3wYL5AErEb31vjrGcTqZVyWeOSqaLcnOb5tK7dzlnZTLZGpLaKpx6hgMC3ad5cc
AA5NrF0YUgBVHxC+ibhyvKXKMQKdh7xgtHbdGP7pIz6J+DqwVTR0xzUOeKwD1HOqvyanQag84K/1
wJdRDUmeIqlFK8iaK4I4XaArQhC38KnlpIeGxnLiwZsCl5YdeK9rRnbpUF0mXJ52Ubd5s5+jAz7+
b7nxCh5LmxIPmsJTQfTeAYZxyXuhEG9brV/lvOrLZF9G37cF1CumTtpwFAl7Cu6JNUYqU1yYv5Kf
g/JaOflAbwvtGbEdzILGEY7xRxaWkqNgLPYKGYZ0jPNMYAMIXYNl93wLbUW6/liaxmbLke7zNdIK
zhCxsjW5Rjy9grDNlh2d0Gm+NPnf4bWQIg6NVuKetP82xqCcn8q/SlTmEGZ0z0c11vGhSVbmu4jA
YMcOMUdY7kf+hkCLFFYC5kyyiaPwXNBt3ZHdd+jpVPkTtIFD+bnjKy542+TMrhCFSquvfhyKHw+1
TjSx83pAabOndli/crlu1x39OMjodl9RDfhm9FIDxnlW18dPqgkB1hTNxCyqyvYHtvOL/PS5rfFe
qPoqwRtpdsFRWSx5zodpEEdEZDamZq0VWCsQvI/BFFwBkk/k7+oivM2I5El1xTntboq2CeQP/uxk
IMjvbzCA2feQ9FFa5Zrx0tlBw92EEnBxdY9zhdtHpYw4wPfq/zZ+756VcvOlHAqcylTjPBXEkKDG
I+dl+jppDxCy6Z/kIiN69ODvdCE6Q2HBD/zeIUx0SSJNd1B3tANGtmsXRu5AGBR+iIIqTUPslhq9
53C5D4u1LEprcH3zpXRxdNiQ2Kq7h0jpnqhRxuYZ9Dg/rlCbvPXAxV3Z+1QUVLy2BI59h1AGlBHt
ZO3goHvNrAe1Dq4uL22IYaTYwBdr5V4IEejiNnFTobpzZLgeeetNquNAmtg9Sw82P8rzt5vnv5Pb
6n9Aa3//16fR2GZOI92hg3RYhiLTUeMDukAGCXMPVRPtkZ1ED3DLma06mtGvYeJ77g4cVwWY7rEj
pv9hlyad5PbZXM7lGln82J4Dx4BdcJZGWOEVyRdONiCYbxodYNNnbtI1CUWCCr+OgKCv8QmtWBXG
rMnheV9xW7bWeR9ScK9bObwuJbZyB0GycHEgyOdjMHafjUmnrytlIF/Uqs16KuxvbSaSax7woBUH
IwODpS1nR1XJ05CQz4fk2NrzSSKX/iPwlFNcDeBlPxa2KlZndULs9a3Uhnxrkf7/UDU5dEdwdHNa
75/WX1/YahdGUNucTPD87TFiVMA88p1S964teFmdnXSxNKw8PrBxShBVFBK27TZlwfPYVYA3bG4H
0XydcUD6Mmzw3gBBXDslPwrgDPCkaNpZqtAU40xgXeeGfxhLAf9lSs66OUYcHo9TjkOIRS0F5a6X
IanAdPAY4G+lJR+wOzqiYZfLFrYtVVfUPa83qwOgHcIoR+p/eDjpD/MBbOAWD56jwnLrYVC6PsD3
2sYUaEFTA3G2gm2geJ01jNozEZpE61XzChPy0+bDU4TjwVjDsA1BqTr+vNyaHQ7/6crT+OK4Qdgr
HfXG1u1x5ZucbSr/TgvImVt68saOI5DWENcX8G9OPAqzjKJaYEjnS4lrnVCjZxt9/Rarm0TChg9A
Hqr17HHrwmFcGdfUHA+uAfLCdtWaZSyeeyo8XF/gwlLygywyM2V2lhNZRU6Cck70VA+buFoTOSR8
iGsDuBlummf3qO6rh94HPyF4D6m1+TWdzIBqHjQKdBCg7fqoXL56zbT8yOoQJQd/VqximFqtqJhb
3tJG+oEyplTS+d0h/HE7KQ9DQdD4jlRfldXVqM9h6SyOGp0l4czsrPcAkXmLdxpK87XwB1ehu0sB
gsbsu+gOyUNLN76wSXZ5iTT9n48lfGPrrmqBjw6KVXVpma4TqOwFDSOQYe4y5CowjXuHG4gLwwde
rKe1ROI7kfvidkDDwVgGVUzWXIYpoD6wO1oq2UuVDTbKXR+/FgDLv/n3K9DDCgkQUDfN4sKocf5u
vqIiS/S/oyJfu+JTuus1lzlPQE+MArTVve0gjIbF3MASicWnBiYHASBTtAMFrDMAa27oxGYQTu0S
S23dEan1CoTS9IIFRDd+BvELmHOZM3i5+ChBpRn1RvAanhfk6wwWj4M/XzC5u4YNz2L+0DViFDvh
yCVuUeW4b0QPdMk8pnFmM7zNgegfOtPDbNWilkPDQ104OVQOZEDJkRoLoby70HBawdyxVZiPx2WA
YJgBTku3oYFxuEKXPBGaUtVB9tE6KCBxwk/3Wd+gaARlBLfht3KQ64psA71MpHJdlW8IoZEJKnK5
uNDNqDpIduXUF8dK6xHutByCxX+MOWOTcfchUaIf1NkV3QhrKZvRlTtkuZpq/2OSjmUI034nyIJ1
wUexEbnss1AmvSyzD0lAj592uYr3Fv6N3ay2Lc9WKYOZP/qgnjVr/Kx3It4NHpgnom9mtAakwDVj
DY4TEU0+eaotHYc8ToEnxu9GGc8UVGSwrwjAwBYRZraHtqGcsXzUysfHVKJGDa2UblkAHRoX5HyH
ot/TFqZ0l8JClFszhpAQBrX3ja0JJqhN9XmQAtjgUPgkp1mvc+mXp7z35Io4is6bC2Tf3SF9/RVB
0YeyKnEX7EUvcbsTxAD1I2itTJvEOeqsUHw2RMNGs1sa1lW4G2D/jpOpEAv3Qtd/VWRo9xbkMfEC
JXore9Ox14aeMv60xvG1Z9+CBjOUAc2wd4vW3IqjEYWFG0JFjLlahIQEd/exDRgp+n3hiKZ5azwU
btLQFjygqGAOX3ZmA7j9OixQn8K10iJrQ5H6WJONgsl3wi2mL6fIAsHDL9cSLBUePcobJ4zaTvcr
9QQ0cKccaVXm8Xw8smcwleuoQAhUD+HJ69ikgHVCPkrzpMNJfs6wK7utigNqp+fUZHGJ5UBxwJ0l
b4fBxDGLf7WFiivsTF2fhu78a9e6+1kMV6glU26B/+cZN9qyGbegGTNINBAAmMMOU/NXBVpEHauL
yMMCBXSUsUetFTw/wVugOtVgjm0s7nMaUNa0a8vavcP7s2lsyQOw+iK63WNjCN8VDWz3YTxzA5v6
TglGV31lGkd4lUjhH4Dkq65SMbWUUF/ptDtwcXp96SY06DnLooKUJE38XzjeeiJOqUhf27NO02PY
UaT+BZN+28vaHDomWGXtnHjKZSj0wJP4ElpolMPNBlmiWU+tFhA+fUYpGAsTvsOXfgVBuhPftyY2
Bgo2b5t2A/DW6mO3P4cwmydkalO3AkjxiSgWbMCqmobE+fuZMFXeVWwZEBUkbAbrXPxAQ5rJQ2j2
rumqU3YqzkB2FS2AUl2/mGZnX1LqC853jN94q6y40xupho6Cmmg5s5KiygHvmqMwGhoaRFJpqWmY
BBwMPEASz9LR9Jb8OQ+e1ArVIjMFoPOI52iY7H6FcOozEbGn+7dTBCzSa6d9EctNG3/kemebSSoM
peobE2xmF5t7kKGIM+R+//zj7rEJAWO90yO03X6rpeJCnkWd2DglfKIAhScNlT8wrHskGMyh0DzY
X78wxk2vkmYn7Rr57xx9VSlgAKPfEQBvwN6tgXo/qPoA8b/20xh7W7VvTrbIP74BwvodCwsvyPXw
wTFaUeKAQP4DeujnyruUSL2nE9LzfdCIEnn/YySpPFuTFMsBUtDERNuGngBcMN0kSTKjwiMJ2W62
rixJXqA49OONO6tx8cUGVfNJAb5esLPZzSZNCLEAwZAiy+XBv2uc4S77xJoJB37QEhm1JVsrC1Yn
15jhp1GOuGWDbBtLQ0f2mmDYXKe3UCG8rni0ewzJ7k22EMguuIS9N3hxzLujiDrIDqtlBmIu1+9z
KXJch5J7GvLVVao65t3Vx6xNV+Wi1ENQCMsOeljmU/ElWjfW3zCTD6o3nqXNMxA7oLMNBwtXkg6N
XiALnBZ1rIKAIGuWoo1QPtldsAqys+X22IEkpto7EvGK6o6IzjFRELW3GBNFmmpUtfe7wXxUEFZ1
05/nGnX8owoDNJQEsIhoAcaXGWTBZXBokkvBaHsYXVWjjj41RxFadpYssUVckkSfZ84y3IkLv3Cn
nNnJ/J1fTssWJJBXXqQVA0xkCdVuRvtD6i90yJ8+hKsWRvLk7fYxc/3IDx44ttr2nCyNzyg4gReS
ooI4qVX5q++SaT9jWfL4pXnTVvMgJ/Z4GSkTPZ7cOjg+VSl9OG3BYxbUrXcmwf5nP58hnfxPj5Ej
+3wUz9yDG07Sab6OD/wE4W/P7nkJS94bN47m7tyg5pSKG7Dzz94w+fagYGeTarmpuenVotihuHE4
v7Xf2YZ7XjY5EVxUkCnkCvWmkSVm1uxKVBe65z+OJlG+SVPwW7BHBnVy3nVPO7IcIz00CmBnmZI7
lDq95qnfL+3pnnNXXqLTwscFG0EMfNUN7+g/ApCM/1jmJsluaLXVjmi9z3aW34NFfiAJpDLj22Pk
Y1HPpyrFoY0x62NAT0V4+O0amSmlkNLK6nyDdLN8EkNmiV0RS8bq/jpj0a0zTkY2FZ5XpTgVR5fs
tDi+VDcz5G50S2t3flEbklD6eefwtlGGqIqdbW0TvAmX3ud5JQ031SP+x7yd8K/D33pAfAp7RYI9
RQOeYot6LN63Hb8ENuY0XPPwrC+7ti5DdqkS6RiJcqjwkiUfHx1BEcVAHqExmbcZvP0U06Cd/RVS
WgkN62nAeS31aBBIW59sUy2K1pZVHGUaJC25YIFXm4PY4P5W3XsGQmVudB99fCMDNh896NyAkA2n
VSMihvUc4Ie8+ihZojPrNRNvj85vGxJk5xP7KGLPyyOonM7ESvmPJzns0fpgRfAsmj4mDCdtP/3J
wZPlq6u+3kKH9AXSSyz7XutzJW2P8y6y4Bf/G6FAxdRmcQtIfPJd5k51QVuS62ZMVZeyXD0Ya9Yb
oZNbSc43p5IL1ESBzQRMVqVc2FIbPmpMfFYNN8ikOH2/q4DXY66n7NsP4N8g0fa0ttIoueXA6pEO
fjaj85SjKyip++WZ9smfaiedTTsALk1pL6sEhnn2SVoihaiLkMqYB6g6F5h2fiPQCPFvKp87GKoG
1DpARaj8ok9HahKYKTMmsKypqiPsGpIzEx7FFw/Lzff4gStTuatQwXXAZ7YZtFdNOXSmVE1fDf2Z
owBPNeiQRoe1uMZqJLzWKrxrfpc2uwt2TTJGtk0eYHSfRaMeZrb9lPrmsiutScE0oECUEjYQ9Ggp
9XpTXc68THcbvse15tP2nZn0Ujfkty7pfqRaB/2CryeKfugldu0KLcuUTi0HdIJGJ7ToKehEr7Qa
VFKOFqBDmaUaqK+Pfrw24Ci/UOadj5A/FEdCMBAQMIeQAr2Ou2fsPcKKBBds66qWNTxeuZUG+E0G
9Jlg3Bm1XLln2Y5kr3u6d/fgZeSeiZwrbiGm+XaeBkxO3olZSOlrGfqMszt5Dfx/6mpqKf0M+D9X
9h9n2LD6Hso4alNohSTIyaktoSRxT5iKpEA3SDssXv0DQzvzJ1/qnptPtrl0K8vIPQUi4CxxC9r6
P9lV1g2EXCBGGRsBJXyggwyITIPD9JF4W677R7jwj3B4fPKblZt4be2a3+fL7d/bOT/YsH7KJu5X
7yXzrmq8TxTFv+uZSzH+nxngfVwk3zyUzgSYsjuy/3xEtIH8vE86qZ0wtR6NBJuJMbrqF/MTdWYP
Dv4PlQRAVojx8ERl9dgMWsPQiwBkwUjgmtdTPixXJCUqVce7LWKpdxUGIfe+2Xteo/PpZNav3YMD
A7HzYr0ydKJpO+BESbZdNmcA3wj79IWNoFFf2qPx7B373C36Sbz6/LqUnKa3Uu7ntBh35Fz5yz/l
8N9x89siIbabZxG55hLmXN9oeoCsp599oXWsptO0I5IcWg51cRvspL9sDrRx7Qk8CzAqZ/a8VHAk
LL3UE5VID6UjhAFT18/gshHwNelwupwm2XZZLNGWjqioZQejMREhR5Tr0uA3wmTh/SC/6lj37MIv
VlN4cDTiLSg8mgoVWOXBd/ZP/P9WT02+ud1A1m1QV++Jmhi2aYQExwcTmgxpcp8QxO237ri/b7CR
NY6BZcx46gVdqsOB8KIR2MEkSKc0kQJnWFhUyvoUSYSEOVxcgTwSYQLOe9WB7rNMMuCqeqEGQ+/X
ripAROC8oYOyGDHwuDqknKA5c9R6j9seFWmEibfLpMBIYDA1qG+BvzO/0qp6iowCRZwdF6M1eJUG
AIQZq8HFbUI5LjMhRmAIu9nLCPlXQDRhuV5+om+YuXEdKP+KC/ypLGZQZ0stlnl2/0sH0dqRS6qr
0KSnr6zFmJS4z64Cskjyct3soXC/Rdq+8ejaMMMsKo/pyQGSCCqA0gH+OIone5a5TjM/d3RgXL2l
2uL8bvJboQwDNPC7zRwvIC/mXUchMpCzZRuIveXkSxdH5/nFG8McIyLIEq7HKSNbXrZch65UChxm
1anmYHY0dF972zyO6F4Ch2yR18RlNZujqRsjn+oYUMFJk23tVledJP9Gjz0ioz89ACB6SlJSo/ps
XmFuJZhFh+Tuj+4oOC8TenoWOvI04xUsXns/fmPe9CLlLIcC+cuJOqU/acUih3o0uKIhuRmMyN7t
T0uBNdfiLUEA9xwTHqHNnUMLFUzNf6OgtpCi+gdisdNvnxdxSzePBFpaPmF78ukmtMOo4MAcYDjE
vZo0slpirqtfxM4Vq8/n8yCAIlj/qsgWIEsnzTGBcVDdx1ACrxkGdCMBEm5kXXqU93JIRPWX6Pa2
b+G6WxyNnTCdsP4ZWgfmhzzEtHB+D16YF3gahjIzrPU9B/NrjUKg/lwaoNIpicNG2DrEpq8ISr54
9xnKpWG6pGD5qR+YvyoweVIchuF5IJulPjJk8V5Grv95c5GSLhn0Sj6+zQQnqYNtqG2rwu5ihJqH
yOAhN9mi/btQh52vupMW2+nxEiRfKP/e8zpXQN08BFR5BcpD72Qg2xWJxlPXtnWi0MjNm0my9VuL
p43H6WtBF6G6EDStcEnNhpdILf9H9Xy/n3LNNddSl1XWinYYHaoDmqJnH+3mpNiluThPWPLfuIfq
akrzeLY/rh2eKdafi9997fUvdQNlQoY33/7lVnLSwXrPUmI7xS5P752WlV2Ym/Ze59QK4J2ieLka
DUcV8c6fxDcPGcZaTV9L1OO0GjJ1o2t1IJod5XfViBAJODM4PfEzonekJW+k/QsJkukvBSJbjfxx
Cl1SQiDHT17aEpyi2sgxftmDd6Y8u1eKVioly/npvLJchbVovtOonhT0OxH3CLcAd/wBYUERpqhI
O8IhOF26owvmfCvlE82cgs+YDCZR/3fczKOVGcG3UUsFFIAkt0I5/expWCyQnPHMJpn1wxilVlGp
9WJDlOqFN28dzE1NLzDl0UZqnmbDbTxqRQbjoCB36iWkKCmPayRnghEw3eiXcbhTgPMwGlyJy5wm
cNWRolmuxlm0wX3DnyPV7q18IAY83ZmJXhHvwn9ePRQT+ikOtj0nzJC+cNvGxarkOn51qkwkrANg
IvWihQBEgYtl3PM0shyZn6cAlYwwFOvAUeddSo/LAkUA22ggAfAeT7WeoR3ZAARkw6W1P5lMsfcs
Gc58BLoy79rlRx7wRtWdEHGTIfJ2ZMy+8aYKdzoz3hY8W2rWdyrmLyC43yvlIM0Oxq7uCK/K4Jmn
pwM2Qjuu606YadRNkz0e25y2i5LRgNF2+A4m6Vw/cSgikZinno3oVc7Bfvbkbc+j+FusBHYGcG5f
KlcbuSBDgEkkm5IkZF+t9znmKggrbe794tAqVIAuYH0wSIT5+GLTiVa/8377A5AJBeAl0ynJ9Jor
AEiaOUZ1ZQOJ1uNHNhiqpm3tozHJ7C6wYwkixzh2IyYxMdASFbMhRItqDZQ3KcPkBNQK4jIImxEL
GyLoQ8NpLLq1l7GrZC/e7nxckexIKpEK8EJjlufMeUkCWvNXtTzkoNEjt/29pQAYURZrUmhTyiNn
J4C4TbeJ8IjBNo6dPMwv/vve2fSqanQt6FsXsZCkrO5FiaSpCevneBK/YsMD50Ly+KqT2P/D9j8B
hbKUZTr2URdtPHcGbYDDqsck/5Kwo4S8VqNSoarsobNZPqm3U4q3z6Xxb/WLY5+/qRTm4clxnsNd
24S2PWHxrOa3yIaivmKWbRsKJf/2Dektr5vkL4qkfi3JLITh/pJul7jXHpibjns9p4Sc5BGtQ7Pw
guqfOI//fjEszZCR7x/SvFQIM7eKoy6P0mdhq9e9XjNdtTAVG7p0elQZC+Cw0kdaLxqiifbG0et8
MmhmY9/l+2r2LqDa/P7IJMVE2o8JRyFwPDEthEM18NDknUNsYQ/gZgDcfpodKJsANH0kCoDXYRbD
JxIJJvjGb5AfZ4pVvdX/oyZJTpCxl+KRQ5MouAHWgGWeQX4ZR7P9QRwEXhE7fxfl9biWj5TgMFwW
8AT99/XkPDavc2OzWpkmkc46KYLFOy7TC2a+5YAofOiusvNqfuobNfgbceKsaiP/cW1jBILQKJ7X
pSg5miCRNIk+wgsvTEDbb9FMxHvX2nF09ZLOgkHRsdvBR7UtsygJmH8017QvP30CBVGsLEsGMxPv
1l/11TEObVhhuPv0w5/OYnpURZxV7EEyOlfA1/9CPY0f3Aczo8YtodPs8SAORIh3vTy5KdCjjVyJ
lAk71Qjqqzw75z9DlbtNLE0eSgy8aa8gze4bmDI92oN/Vr1/KA6Z4O+5+b/rndPWMk2pHXO1Ti2O
fSRyGUv8tB1CKFJFhpERjLpT+E7MTzKc8QnfiFUvpJxxMIhFahKuhBTLBKZmKZL/UqjcwmxsK6JS
nozFNmux3Ok1hzZ8zl2ugzPc4wT6iREAls6tBgtvv607/tDNU7s3Kw8QajlfeVhBXbNap4AN1FZh
8ycroexRll4NA/n9OsNQF6gWMDAspMk0jixY0p+5mgCmhMkthRuPX27qP7coWnztuktxUjSjw2n4
EGxo+bLSGu5aU89cHjiOMFB8i4+v8zBHS4XTS0qRNiVQb0CDUlwmSAlxkiJ+hCrZe0ag/J1NxgYA
+Pip8ya6MDCKDv/nmuNsUT09KjOCg4T/r9L4RzfkoHx1EWBroqUE2BI3pDzUtp4fwxdxNjqtMJZL
VtehZy4qONcjBAg0NiyINtv82nMYiFWjf+RcfY7F4yXlFsoSDuf4eGAMqJ7lVw6pIu/lcTpIrr0Q
vbnZDz4759GIwvfVJ+7HCSHEWfkcdVTHPhTNMnxp5giZ4TL3MPVfj7hW4HtOuhjw7aLjsT+gMoLp
Rvg3g8KhqFIc5xf3xDfD3uPBCx/CJYS7fLZR+MQdHQwJS92QSzQBGxdBN+yDpokbavr/4Pv0mRo+
/Q7B9CYpNPMIaTwTsfNKn1QMqg5R/JzPctQRyDfHJMSI8QpUmwdi3yGGtu8mDGVWM+IiFKk2oaBQ
40xckblNoBpk+nXLfGfYgwpb7q/NbrE7BEVAPXyV5P0h/hvY6I9RqhtbKiFBIoZO7FwRmmSblnJH
jHZsUPkHqb1l5si4eGFh1LILIa6dYgbdxDWQ3R1zkCYVfVhrHt/A7o6xSyX8nzzoGy3u3mriTYmk
/eJ33KTUJhWkUKFulcc/FWz1xOcG3HJJkCsz65tmCyZI+n8IaAyn34aXQJRCilgSjmlAkLiivkT4
O4VzwEHHdGUpbhcbr/bSVyoTtSYuf/c2jK0glgOKVSVnEju53bpMfAzejCSay0/asYIgd5Hh9lMi
TlRUxxmuNAz4ZKIlDPk2G0gvfWSn+LvIZ/L4u8GJiHBmX3zN/2QKevUThTbBtgM9kew3yQyMRDZx
aAOwvryXELWpZsvB4OxarRwLK1ZjRjpzzsD2J1C+dpkQ9QubQn24OqnahYofW+ULBxAv6FEBDUGQ
xzVecMJ2DIlXCntmqFKw2ucA8cpGa3CHXUpmvsS1z5KQQuI4LpcpFzrw3gMu+T/XuZ6tGOg9/eAz
lJD6ZFWIvlxjFnGxe71uv9XbYYRRL+Q1EJBL2qWTNpdUUKyv9UoIuIG/F3ITO2VG0PkYn9iKFXW9
7sdCMcOExJt6SqaCnrt6+BqDzReJan64qg+cvrej6z6fxrJ2pU1+MA/sT7/4sIwksYI6fzpdPod0
vw5qxkIQLTa0dlbF/0mj2Y+Rr+v4dYDchMMLU/njVh5teDlx+uNu9q0ElL2Mjp7Z7QtH0L8Q7ChI
dAWye4Ax9EENxjbtEHxr6ysw3noLX71/NSzN+22gn3CLMJwh+FK42NiTB8/sCu+zc2G9BNma1HLt
yT3e2BTC6k0cI7PbkdrZcY/885Mj64M8gP+WwSXFlYf27IN+P+7y6OKzwo+s1OR0v//bIwORK6ha
Je+KouWSiUo5FD85JmRt9gh/FYBl99dDHTicw8+XTCTuiK/MzAzjKjliSzX+nnBbfhUOM9vDDrOO
1l87fHXx2zwMzT1HxyLd8E93JPaN5RwEPj+TkLeci83DEDMhgzrcerPMLt8/CQ6XRVJavDALY5G6
QCsb3wLJhhFdWedPQcDWijUKDEl7zEcbBdDVlq5ygwF1RAO3A8nM/iQ3DXyaHc4EqZMdiAmgDtkE
kPAOFRjOb8gIyL8EAh5FA3FaG66FilDoGr/kPWJXjZC4ifJkves+MYWKxMoI+LmhLQKn9lnNJR8Y
nMW5d0dNed00xG5JeuypZ3lNISKohqBMCVPzMHRbVWT0SIIjsY+rVNz9YUitw1CGNddz+1YQ6zzP
PFieqXAkplQVNIv4Dxjlv4nUxOzM/q1EJ02wUYfSqMOo8ueRf6raAf7E43Dx2AIHf+iK68hLtZfN
RThIR+Xt4qAW7TcZ3hk1rYo4BzBmmPgF+PcysiW10rljx1y5U7ZwuUZ3YbkLjldVVmD71dep7p6W
nUmg4gjwXwmjxXLtJiT5uJod13LU1lz0R72sDXb9rWhIZF0i4AJywUrBFtQyXZcTkiFkB9bmkr7y
Bsr8n9CEUddLQlf5DkLk/CvKjPUC94TRC0hBVpIZL0Xgn1PkdEonsfHDLwPM1nrHxQiPXYNkISj4
Ybd6/BAW64XuHB4kf/bN4+HJ6ZK2iSlkDXC2iCMCBufgZmxAIvAhzMZRIxXY4v2uh9Tu+hWBJBQy
OrsGSAAVbA2pVyc+TbCy//SGjPNIL1+D1wfNrmcAdZ7o19lBDdccWl5LqCg6YDOAJ/eQSZOaIcsZ
nhGvBjYhVKN3q8lA2+28JMf0WPIk9NzcjPXlRR2/uKwCvwXRLmBunwVIBU0IQRIl8Wv916o/jsvz
jNDeeo4WbggcFGElnOATDgnE3eG+a85Qzu86NZLq3UqZfqyY3cESInOYS3CySB89dXTiYCDw/8cb
jRcVX/G2TTW1lXfp3zi9zhxm/FGg5b4y2Hxp+fBZbSfnDWO+3lZKW/XYxjlthRYkGq0HYyRpkn2i
5x+VW9Zy0qrn7MlzTNRwyVoxtMRw5Pn1oGjpVIRUVG82eYey51PxLVrm/RTX+ot4bOhV54x1QVN9
FzVJVk0b4TMZiI5jG7xuzu2SBOP6o0MkLnLpMQouFBS3V9VET96c6zsZXqKDCQ9TmNOmfyDtx2VU
u23JwSlleOmn717RkooBerjW6IPyLvmJWZjZQ73pEJLbjwYNteWnWFfvGvR/bLTStDjQagkAbvAL
P1PSDVNvWFs5bOrfrGwK1D5TVQSbLc4BGUptBaD2V58/74OQjAIBJpkDjjdhjIxjR8wvJeswmSkx
wkXUOh9pR4OKGYgwJqnZiqKXHbIk1N9WSEQpvjyJ7oCf6PpUEODdztOJNmuOeHudNkUJrwIW2PCK
GrdvhHDipypQB/u2Dod1dtx6EnjOM7y6gjjXeumk2Iltw+v+CCirO5XPb1T1gkC3MP9fRhJMCFtF
OcODUbXBaKmX0UCVfWOXjm4l6VdhhMJi1ghq+DTpalw0hVsAme++EeJb5agxhKbz5uKYkJ7+9ua+
cg0dg0OSZMVTrT80imEn2fOi16oFQuVdwyJSASYD0yQwrhmeNaMwM/vvcadbLeYpY6CY8VkEpSrS
wpqaqtn7JQobvMxWwprnGUbX6uaXF8gMuNGhgYoks+eTJcSCGZMLGKOUh4Hae/844keFAiNr5KC5
Sq1D1NyoOlUsRsKofsx+URSl2mrSdiiGylvmgMBcCrqf8QrR7Zk8u190yUN4zgmoxjpFWfPNhT4+
hCkV2I0sk8InzL7un3S//0rXgMkLV/muyliqPrJIXDUex92328YVtvHXhO0TVfpLu7uphVXedGkv
c2OURAHw6Bi1zdXte5cXb85VQ3k5Rtxa5P4Uz1CjtCZS34j0dGu2vVUs6C6Tak9nPsOxH8cGyxE5
SGCiKEbZ5JB6udjhfgFmXeREOQSJObGBQH4bK6vfX0rho49qwjYmxKo/3jv89ERIHeun/St6k7P8
Bk/2TpxsMinSHRxguOcnJJj/TWaCRGcFuh5bygX+dp0BkLmRGcIN7ZBNj8OOX48DSA8KbG3Jh+w+
6ewCzSS9wUzv6owYjfUkoxHxuI3XhosYxBKYvt4pePx3+DemY4Raud8RBpkEHsthvGbt7GOnFfpC
9cqi3IPrlv4AUFiJihQRRXPC7hs2tY8wvxnFwTTJgyMDo+YtbXPhi+V7AQ/TLWWBHlwni4o0b5Hx
091UJF9e580TsihqiIUdus+4OvBKPa4ijG4l0wqRxPCLgiCgnlg3VRPbyhR8p4c6VLyarKcIeEde
tS+y5JmqXn5wOEuXk3opQhiUzf22lAWCzEMyy/6gc1Q6p7zO8+ZjILNyBk6l4+IonrK+4J5bkNF6
ZolMce2dQ1IKv9zKnk5D8rMqeVrSyKngY5iXRroP/7qc/e7e9Oo6xHMSbMNt2//AbwC0DHIDKj7x
qI1MgN3hkk1m3dYIQPi0ALnjuLDvRS5iBSI8MpIn7Euhhp5OpKvFmskTHuQI21NKXLQTLVJEiap1
pNJfjJaOxFrZobsqld31Zw/e9TEaUZ7Xn08aT38dqlxcgOlR/qlsxZy+CKPzN2lhrj3xvrlcUUR4
HYgVEUWSUqWxmDJDnSadPurYzOFWXcRl9gonaqbAWhFj1lCWAV4nOGp+s70a0+TtRnRsDpgyPfhI
woumEveS9c5Z9P7LjMkeXzsIKCUVqgkO1R7YURDwWGJHSM05/s82Iwp5oN9F7HYZDrKDLqiSR7g3
jNAXRROFBE6r4i0HvnObkuKr3d58HaIpOmoIJiPb3UzULqosWJDziDtQ5Lcc6x4y5VR6Wz6rZy6r
BDzUoRHzlE0DTlLAjjjV2WhQH6EKFtjleCXqMl0o9XHfl7ge+5Jm67tsbS1Nm25QPJ8a/gPVsEfL
0/Unfca3UcJomZes2AUbn4tddVgbcIB6pT/tdFdPwB/EcJho8tpfVb1DtRgP8epBNfl4LxR84N6O
ISKkU5EIgFIgRj7eBiCXCJFhOxX8Ar0Q12/3Lq582qN42zYBEklLbDxOsK+UePtPLmDirxXCx34v
US/dO3A7TlpEeyHi85/CeNmXsiqIvTPbRyxInLLn41FIX0WVtU865Ue4O5LSmqgZQheiFRP42cW6
OsFkzahNzWKPCetNrzh82JnrC/Eb1PSRK1AadJk5K9zt7n9TTUgPJ0ddJiVtM1vBcrd4HCPj4CT+
nQLYkusGpsUnBIDfuw7ULidvZWCEk7m8dUjDhoqv8RXXF3CFeiRb9vZsI8BEla91gh0Ht2HQftqB
Xvd1e7BbeznShgWacJQlpJvLf5tOcDcHnt4Y48OFZ+kPYgEOMJm4k+p08Z4l3efmnSbPs4UFaf0z
7TKiU0xDul03HV+oCcKLzRLbehLZvu/iz+6IhEYcbjpooBemA7liaq6ct/8atrZBlvu8hwQdbYwP
15wCzJslHmGQkNQ2vyC5TyfTxd2ZSZxW6uoJjhKnfZ9udwc+qLivLKQEnJmE6FhtDOaIQxYkNMIn
2tdD4gAcdgsPtaiRrrubwwBnYrzs8gYZVmBy/+PXsgeB0B9FeXZ6CeiwukW50IEnUrT7d64jRZdy
TK9JCxBvxk4/Ka0GXEaO8VVdHmXgP5sx80NiStNSdtbdFUU0aA0Euxh0p6usF1v+D/5ma0qX6oVI
vvsmlesd3c5s52JtrNLyQwg4q+9zfJz2U4OR29sEb12IugrfjT1lctd2YUUNvyS3Y0IbzYknuHOQ
7b3DAiwz7wbXCijEUQtltbCGMeTdU6cItOLPSCPypTmTsfbOs7ocimpR04yJVnvhjDcKmg+vdGsq
N+i7Aq1/FKM7KHhZiy/E5Ui+NfNgBHQZp3+0LxEYHRVtndZLqmbsexAmZ4+Xl0aGzaA0sFLCUNOq
0E2k5sQKYaYj79MPPoEvBqk8Xdv3pMzuQHF5AWBN+W4UNLAxKVBVyJxfR754Vwk7KbgHiyigvmx4
vP3fq9tm6rzgTAxzAWGWFzrGlrDjXmnjvuQFLw1xvK6FzwzTsN1EVdegxpsn63bfLKN58U8wg05c
d03Iu1xtt8lGHMkQYCMfx3nI4voGoWPxbY2HLWw/4RamilQNtpcJT6faOa7z797JqCzGJ1zvXypv
OkfonA2SK5G1zWL149L+WyG2OWXAOS29BGAS63unjg+f6awW5IrRucNYeCRCoHo15lB/btEKw7qc
BxvxPeqTvfD87wyFOILDbG37m1mjjcVz55Sd/pWBeK3Yyt0FLEPimmuBCqym7mjbVn5jbTajswHL
ZOHlGQwStVd3StyGI1pq1Pda0ByD4Obv4/AvKz7CMei0v+H9VaAfwEuZbd8841kv8sHSpBu0e70o
hAYwtuBSyDwAZnR8jMO+DZDzljSks6W3e1kj5/Mm0YWQ1YKkAsCQ1CCC2orYge8vXFwD4Oqe410u
b5ytODA79wXXHq8rXMtuoie0wIiVliXJt7X7/DU2YYydWZ8NvD/Z6/DuHkQdC3y2QDMgIAbD4vjh
/WctBJPviOSSxIejWNp5jHH9mQYj5L0RW8N86dV0k29IK5ydNylOigHIuIJ7sfKRh4aRHTfm7wAl
UyUE8AReoHz0LfPQn2Pb05bRkuOiPl/eiUOoG2l3wfAuzGV3/rOjejzqC5AOYveqorWSWIRqxdwQ
anFFws8KIedb51LVcya7jP7bUsTDkkqe4PA2rgKyNt2ZWgSeXH/q6hVznHfzaUs4tTZQrwsHF9x5
y7b3PEQhSrSCHUcDp5Czq88J3ddkuERQ0Lmv8r88eJnq4AIYZiQTNYqvwAqusmAXTTgdhYpWTzVF
1pt5WXAjQb9DzFZRoTkcoTDADmVVUBvUu3UduevqT5VNjYcBz8bJAoi+pNX8TsnEzGLdc3dq07jJ
415uBxr225CkW1qlOvxDfgtuQgrdt2urZXwLiRoZsMEmIh5+5nPC+5gpOzH0yjvDM1Gg0xUX9oMj
abvoCwYeJUc0CLbk0bybt4+FLftertggvmejfOvxAW6iK1ZFqr2WNTfH94LCiVA/VfryESrl++kJ
8Sv8InznYCp7WBuGJ5ue0FwpW/ey5O4ZvcxA2bBGFig0ebNsL6lhNzN71/B28+hNezTgKkQeKLIM
4/OF8VFH39Q99V5GK0bxSpSdm/6WpGlN318EdOeQCqBIGZvHCSDS4+HOAkweQ+etsSv9N+riMo6d
i4stQLP5yK3hGTcsBl9XT6GyTECuiOkxBn3D71nL3cakt5TqT5J2rPCKK7ZbP23fhCD6Pq4/drGX
wmIQGTDIG2+xBfovX7ziBSOLcOsQIUfkZmx5493BkGTR/Db6blEc9JG5s83YPvspmj9k95kbfNGy
zs4nUXxypmH8w7ydnmYaueqQPUsCBT+EWpTv4PcuFgwJBEhqv165LqcRuGC06GdrT6nhp5mDzoAt
Fdkf5Y7fvFuUpWHIsVSDnQoBjLL0Id98GKzcccgIAJDXIBDuglsK7/TMF18HTOKzc0hiupWrGKZY
cV6Oy2FvLXsTL1sOEtzVXSdQfGDTc9lvOkYUt92qytq1g4izu4fnVx4IENc0v9u+u/RRdBh2k9iN
2hnGE2zkQder9sPNBVYxtheJVnjC7jjcGa103ugAXk6gvJRH5DwTdEL6RfOneCeSLYWYHsDV6dzw
2ohE9iURCnVzayWUYZH67JgW9x0DWkSpSt0ofRA78FvILvqRLksJ3iMjz2lx4xJa/V8He9ql9WFO
pB0UhJXLZdk+MtBZku6ZStHtu5c6T5QGVRYaX8hWVriG0txZV1u9zrpCP/SoULuGaX7F+QW/pExk
QYgiSe5dcG8cp13CI3vEiaF6oF9BfIdOtxoPPaFsJKltab6fixW8+psKLWBjO/StQFYYLcNzboEo
ZoG1Gpnz63U1y/Cz9EBZg4gAUQNxBfpocQLqWpIf8kLt8FjPK+/C3TE1x52fQawAY/Fp4XYlEhqu
1ydPhp74BosI3Hv/7pe4OKTZGFZTFo52UXZuG93d4lh2SbSF5ZlLZYO4kndqm87qWqmhT+mTxDT7
pENiwyhws8D0VqsY3iZmQecWvXDFCpdLvKk0L/hw22S3Mq6HuQ8g0Loi944WUak3sO6ekZls6XjY
fs239o5VLs9taVgcPsW5wxnjaLxlJlBSZl14nVs79EMkdYfGa+EeoG1QXkj9Tyi4Ze+y5vBp0ze3
o2YcFhw7+U/bh3uVBv9EKczD8CLTmklmQX3mMr9naT+4FNcHgYdTpBlwH54ylcJKJE3FrdZN1uYf
vBhmD3eqlRCxt8O1OJj8JTf0Rr5EA6MtpDgtaw4PdB8vlBm6qDXLiraFKM5cox+IO5u0WaVc9f4u
t+2DRlnOPXLIYBcBMU+5hypOIe4W4ZLwkSbVXqb8DTaUbiDhGaKxHKQu2nW3b0khIbwaqeWTgBhs
+cGGmhrx4ECm+aJzd4RWHtDjVA9vh93P5cXCnUc5bA8LPoq/exwmaZAp+qwEofg4u5c/3eVuynB1
ZgzsiZxXgLBZz+IKnqThkjN9jTRdK1WymhVExxL9/h62mXToAZIajYBMY3dJ5ODEczntp9AHsisL
WcP6Rh7ZvIpNvhXLgEi0bWeHHAr2+/0fo7Cfefohm6GZ06qGw9H+SK6dUVBt3+lCKDeF31RWR2Jv
t0jf8eLCAYUoT3Vw9o4SKCZBQjCe/St1CRIpX9eNPf3SLA/A92YxsaY/DG+9azRGTVRB7OnxzS82
ls0xP3/UyuIdGHIbhzjE14HFdCq9a1XApn9D5STk+YQ3qkDq7he3k0Z8VRaHAYjGkRx67zykq/PZ
n1b/TeClWt7s6DjobiuQ9xwKKLwRw2MnyMwjNLpEJhZFl7icxBT46UsvQvqJlPi6x0E8krgHBwA7
qKvBAg4mPXXB6fQimjJc1dyUJ4zzCyXdypaEvpIsNLonylaVFB2LmQo2iUdz6zMz8iYLx8L6xyJj
5IWs4VY1eWYcBDwsk7akGAXvPIAZEAOXBZPm/6KwEJWiemjF8COTIwZEs9LdN97Oozdmznp2iirA
iV2UpcCED/DW3HFc0olJWkbbP/QxtP+k3LV3AWeXn+1tjaY5zT9W6XtZgpOcUYKhTyMGcmNxi+gF
u1j8pDwRU72XT2sC0NZY81yIRcf8vBO8nqAi8rG554nHnlSz5HivPBiYLErVN1L4xIjSaGurVj2O
Kw1bT+U2ruM4yrWMyjZkerr9dPWn/BklAMbY8wZ4jrYCEuQgcoGvH7Glim+LIurNmnp6KopYPsmR
7NX8AF6yqux4xhRsGIzYnADj9g1iu5LogReoFOng8MBD+omgnKHTvj8YYqJOI7NH8cOyOsgjRnfT
4Rk6ykKk9x1LyxTMIWxF67gZ1EYuB7zt2k8j3AyLMna7OBaO561RryPn9YmpAIU4rDF6fScpQyUx
q61FWWLUgsiDH6Qa/xGAg4H60j7jqklcPHVqpDipIR1VCalTcrXQZaQVHhUp/uPQKX6ePrmohnUx
JdevNk3hmttyzoftNQP2jAjVbin2r0KrwenC7oaNkxlMRG92MXh83W4YcY9ejiMDSdxqx48jYcan
l+CZtRD7dySRyPJn7qxoHhLVwxg19CTp7M4+mXvZG17/XudWpeOMQRGJvpifplrL0XZWO5WBRTYE
9mP9UQx07rkrCdfFYrASSkW3/fRxwzcshZEf+QZYQ7LNC7YY+fszpIw/lWL5vafphmfs9EjECKUq
aSfkk9A2FvkgJFMWaKsSOILawQPy9F2XBGTPorY1iFYP/gIIxMtWAcmXjZWH2875BgqeQ1S5hoZn
6KtrIe3hEe6v9R+lgTjpKTeye8pQTRSU/nPXTzGWHhp3a1ht0Halux/j6YLwcAAjEXu8JYbwyN++
vXIAhrg8+T1gzzRVWECCVpuHKLWHBuyDHGJcj25hcHImd52d/O2UUocGJedrnNULfw7HxLWP0VFk
eJFhOtvaGuM9hmILq7AdfaXi3nEP3K8fFp5K7CKsF71BFr+uMA77ICGnpb9vxD7teUXNwpXptN67
nDEZK8/R5co1a6BSmYp4HE0fq9DPSXplELr4pF8JfGmMdHQGsCH2NRuud8NRYil41x7/nv3Nc4ww
yc1aNAG1Auf8wEGMc+YOg3cyf9pUbG8vbma+3Pgk9GMSc50xR+NzTtBIkJ6Df3IucMpawiAgWgI8
cQduuIHQeymUCNRoyA06WMan+FXkT0zDD8GjhPb/E/QYXw5wbLUOsLQyF5TnfaYy0047ZqEMgp51
AzYFOfs1sSk11Afz8b/t6xSNoU2pSYolxsYjJydqxfn8ZXVaK0O2OR01uF4tyZ48d1hg4F3PXvV5
ZE7CoDuS58rxf9obL8VBhLKQBdBcFZ3elgEM0WXC4uZPoJfh1aQlDsOAQMzjlVzhlqtY0ZBXXhhG
V2IgKJ+rUzZ8dl/fFy/njgi0Z5XqkTROnU3l8NuSN6o0n4vtueA+Okh4fDJlNv/v9I0ANSi/DIR8
dttP6urkMy9T7kQNJsh5kE9IA4oM9nc9GtBhj1a9fs7B6HzjrcRoImV54kEpvZO1yLPf36E6CWAT
7cXdhfjhdXs6ahMVnuw5bbJAdoIg3fCNYtnuZX2uXstYGvku4iA3mZ3f9HXeKowxVN6ARoAtAyCN
vTjPElAb1zYjyoxVYGKjNutJCDaXDEX2zqeitclqhLtWXnYOyEoWR/lCPyE7qzRdjJX/K+sYEY1E
rh+ynmvouEegtSQ99eihPR72N9U/KdMXWbk70vTL1BmSWpQHkTdoljnE+PnIBUg03X1TcQaQ5VMB
JNCaeQrkhBzO+1Idy132urWdd7keSSJ6+EnMVxC6iQwOgQwRN2efLQe42YU/m29vjEjyVUXy1siM
2KqmgjqN0dN41Qci+KlFFH6EwhVe6CkJG0ylHYxsAAAEwrbm6a6HoWrLQcUDeg5I2Rdjd2INtTlr
Pu4zmdrsdOflZNEBl1woEwL2idQM4J6SaeBSzwPZjHgtMneeWXmVqG3bPnesCKxilgIY5d+yxdU9
B+Dg21mNHuJifWE/2y7g0dPk7PhnT0RBvp5dVI2PyFBpIzsGNQyyBLbk2tX0ZQgVk4+YqMJeVjT8
l7E/tZb2fY4psTo3bW2bybI3RDNtqdfIv3QI6KVfHWK8UZE5mE357y7VC2Gz7KNUnxOFWOc/zYKt
TkkV4iigpdrQ733LjHRoS6CMQGbjl7SbancT6eeqLN/zD3BLgUbCli3RTJQv6Q4DW1kfzY+/hAHv
XDwMWHjYCPH2bpAwjOK6aHEXcz/jVblsrfgCsZlUcDrLdd2nQgFPak9s0jqQkqUqykJS+ID1LYve
zssFY9lBk5JGWn4tf7+pcVwMCrdp6OKpafQ1YXUW1XX45xwODmqG6eLGGSNy7RVBrBUXgisgyR92
aMWdiwom2hj3jU4PNeqblY0jRYaOycKMyd0ePIR9GMohfhyKAt5r+8jN8pUG8cD6r33MKOx9tgV+
HljJ6hWfxlr1Hj9tQwvydAivMjfSdAMJNWr3zfUQzGC9pYq4aprUR94sX3fcPYRTmxDq/fo6GSfY
9S1z0ZzqF5BEXJUfuJaKj8IOrNpUflfW8SYaOXdKVi/Z8oS35NcOAU1Pkn7c5n6mqvG1zJbKl1V5
jat1+JGksqBr8t3lfk/2FDe0u9fjnbAPDvjifF/Fb/pysTIt+FeT3cF55udcBLR6Im9uAeJb62qe
0tWdUiqHcM0b6kOuy6Jbu2SGPaa8M3eW2WhMmbWj08GTSNHyuyRtpFh5xyhTpHR3OUEAUKpf6uAL
XE7u0SNBiQB5dXfLcqm7P8H8+jn0oWbDskZJvaSex196IMbl6RwBQ/we7zPgWoYzB8WYRkeoAZJs
UyxkIyisrNp7l8b8M2oyxPjXT6PoG1CGGHVvOPkzfi3dAKvjxIVyxibN8IhidXfFt0oBkcH8FLqh
s1L3wxb1yqHa16ZDWVwOPsjeI2HNIf9tvTOs5mGx2Wkysi+TvKcBc+SpzZ7H8WOflSwWdzJUR1PB
cax+63dH2TPiC8IN63TFTQXGp+v1yUthMz8N7pLaSc2ItW1oKzuuOLOJxWZQntaNxzYa50bmkRDV
xVIcP/i1gCSa4kEJAQQQIbrxQy8UPw4c+4Zzf4dT+YfuM1L4nZDUOJutIoOjRN1ndgyGeQMF0Rer
xovsBe64xBzSYZGLTcMh4gPQe9/osXT9vCpDOVxh04RoSr6zVN8iPvxAG/s9dw377g8jzFow4HYb
PHvsz6YsSgY00UTMK6zYpF0I4llOJzSsoQkyXoFhPtqlVywoA9OMbeD3zFyPU43ZuE6A50rcE20d
vkOuOlFBwi4scGQHTDV4OKIQhDtOBoC6fUSPNBkDLktD5YsbjFet+7MbGG3/1zWvpWnpXYEh+7om
vSPmtN/BGYWzgaBeOVk+vhcWM6bp6sEnoLvRssDU3HwPT36Jf4aKJaVVoTjomQUWN3s/OSdjEpMo
c1iTv0MkZBa7sYLiJNNfHdND2bYRlQufp6caoJQgSmr7rYye13rqDNc6eSnaosrw6rEW3j6Sx/zN
+QG5NQwqaFYOE1iqNToKeGrFKW5YLUO6gg48UDDBBeRiQbuVKGUOBRg3ApbM5P2VxFdr/oqR2FUb
w/yK5u+zeAREkA4afrIqcIRC0V59sPxxHPw1kS5urb96ZMBNNSeFCPVEeBDTuxG1VhgQoPQbEouh
UsQXgex02fu2D9SE1kLb0l+2r3/1kNgwN1TQfR+7Dx6+ECZjDqe8hKr2x1Met0VkcTsGELyoh4/8
GMofuI16v5SZDHyBy82vnjgV4v5mmCyKAyhNPg5psxqTux40irhA6HscB9EkNqhzDUvEyPfRLf7O
RtuxveI6tds6G8/xva50QKQaPNpI3FcIuz6U/K5E1FKKA/Izmsor8QQ34DKuDzdawVT3a4g6Ukbe
3+heIJWmjOJ78HvGqeZHW6oN6Hr18ZrvS4YMAW9NnU8LuGkwGNK+AiT2QUZDaoWIsmVk1lvLfw7a
2ac4VeICnHrcrqXClXYAwiHs1OFdJuNpqrF2yiF5971NhPozaRJdxF7PO4CFTeku2fNOALMleyNu
O5cOuVQu+4pw1FJB249pAyXp+rE0HcneNByTyN6IxPrPFTc+j46RVXGpFLreUQXbUXvM9rhv4Hkk
7ulE0j8dODnm50u2OqUSJRkQFb+GVLdMahdj1M3oVY215sblZel/NMBtT6/XT2B2ontz4X+2lyUy
4D7QHc9faPWVq53UGG1kp6NrrD52yhpKtKCeqDlyJ0ED49xRXlfCfuTvlleerVUH9QnOC2oa3FhR
acEwC321NKx3YnnTryN0LxLINWx03d0i8G0rkIe26y1HnegZ0AI0i7ocZ4JfzXw/btoLLpierME5
Xuw77NIUNNSuxiJbwzArrv7dDkJtHJPnhaLm195EqiYCjGr/GZ1VnrqXgWhmm6HixTNPXu0iM0JI
Sk5bme6eWEE2A4UhaPJ7WZ/IMApPFLHhEc0/NfhYDzXLUuBD1c5CbzAlWc3/g/CNPTI+bundZ9Mt
6Cs+HWN6kQm/63evG8xRPqptu6YdPeunBlMs8oHaOq1BHo+V9EBWxNaVvn6gkmpFBax0exoBfuip
mSQLOOM4kv670HlD+5WArU9w1JGVrnXmsIEuqG+PYAurCPOh3aDjhhDxGRCgqnMYdXMvAh33/ux0
OusrqLYbMXn2FXki6PIL99yboIPLWyXow7pUc8E5SbgBeUwzmT41WKlFXBynf/FG5dBLP0EqEKkF
9gSRMYcHBtQ2gHwxfMb1Lnm+6Qovl7jD5k3FerAZ0QKbX9GfnHfOaYz3Bhz7/ItXFqc9pXDTyXln
3bL/kf+nQY05D/YrTp4G6mnCAAAOpVK9v4mOV036mDc+hAJ0p0A7w7WyERNcRzhY+/meanVeOUuI
S2CuxiSsTE4iCrF2KAoqk/smleU5QCkx0l7tu2z5Zrf8EGXtP1g3uayujXcnOiv9nq7pUtip8fPF
Yxj3RGe/Q74yg9wDU19haN/cyQwADMZ+bp+1oCGBQ3Le9vSNyaNa7fD9VynK9OZ7V8kNw+WuktT5
Tbdfelx3M9Tv+TGI0C+8qnSDS7qPUNhavWZyRrUDhJa2bXQkfj7p8Jh1sAe+dowtGerSXlErTYbg
/qTnyL5so+EHzieneFFWyq8G4TxboFiYrnV/I+y9L+jQnxD5K9/i0ZgArF+AG5C1wnWOmvMbr/qk
tMXux/+6MD2h6KLruHaILsdUAOVaxWTw612GjdfraaVqlaVrrW2pQuPhOmcXfu2FJwEcxzOor7qU
Tk+bMgDeZH+lMLDGvWbp8vKOtfTEWzUX3kIdb/Qdihyluw/3WfikGlUDbUCGFvNocs92bAL1uQ11
KgDV2dCaSxNKpj1pduJoolfRKCIPtv6gIqDiBUclTs9GXsUYRijImcqppUvMY3B9fM5pvQ0yjFid
SWbXZUXPYl+uFMmGE9Qi5YTGdMXSEPNft484sfaAp3wvzZjje350QpzHPFZQ4j625j/tL5Go/Kf6
U/BrOx9i0vrSywgWEPXBhMnNa+1iCnNusb76FvFyiEOv3YG12RbYUWDaCSuBwylsTdM+7W9Sc7RB
j4Z6bV3oRpCMBwrtz1bBt4rXAFhPObcSjHBXZ275P3SXuYNYQbjqhsuXGsiA2O5ESLy6Oi+wKn9I
Bt9dIyz/3EvsbZ6ba1PB6mNnJiaKn+PybXfIkjVWvs61oSo/qu3Xnro5ANOuZsOcGc7cC8NJfrZa
FgvocM594YtpUIAm2UqKpIrxOInh5jfqXjP/MZjw+6jhGJyp7hc7m7t7A8Eb8IrKsGGDYiroAmON
mUs6pw+BEXqQcoM6bbisM/sOYQR8HD59fXqevUO+PL3GArYhEG707PpLhxau99e3JzjnFIVqO3nf
YTPwH8GHeVDySm4mRt9E8GZ9is/CvWsUvFwa6jv6x2YNWvKJdI6Q4BoX+7oWNju2Jls2GMqWdVod
/J9nr0R0PSS7sIWZB+zwoE3bLr+vLdcPIKjU07u5qm7SViJq2Aa9MPiPqExt5NW4kybmAgZIoRtt
b61pDosUpWGq5VfhZjt4Z0jowbtzKphaULmbtmqYO9mnRYOAUAQFSfI7rAtyTiIqFrl15EgfkdoT
d2XaYbLY5rKPa84g1WkpkGTQUOCC8ZUp09bCqIEMxgb4jf6wgb0O4ov/JJtID1lJWQdOWHQANgPK
nX+ZqxKqarvwnG2w0Fi2G74SciDwfQrGi9VGQcMc3bElhNyJ8h78Eulj+sowjriOvGuugKVJwWol
eLUqEvvJsV6WOTUE2HyO0VA+TpySIWFMpMpgqjpoIXNbrBocMqNACaKPXiJNYFbs8i/AwHr25mYr
tz2+vL9oO8oB1u49GrPYqZRc1faGoqcPfR6WPr3qrieTnNKWr5GCpdHqVPWj0gU8tdv5Q5diGcPL
Y5R7IenvcYDJCKOdbBfY9wt0woQFfY6RqP0EeMEg/vmYDRHTGKjR7Y0PFY4JtHfhNT3fAJqFtp1+
8I/BZ4V3+7poGZuJCZQuQEm8QTvKZCpUzuP5yGhYyeaqis4WsGXdciCmdaSbdwkfp9Dtd24oQFrk
X26BCPH8Qq/Z9AWmGbq+35MrKkolic1H67rCVnA5gEqNDIbdJhauWBPfraiHrHzxE1nrk/wGnkX3
ozGvNt1pJDR7yqRIIUzdd5HumOrRPNsprvcy+kgNN+vPEsDVcWmlTWPykUDiX2GOrY8YXp6tnbRl
w/pqjVtI5iFUqQSMSX3oDIw/IHnPrrN1K/KGp/jWY1YcYFo827dJKKGx+3PaMBJU+BnKLCKiRyOd
dwCPpYjMSlYHtU60cdHBGM92PhfFJM9rweHmWAmOYWi/kW3Zzs3gpwA8898cIb9uNSQboEb8lJ2X
qh4Hko6Oz9S+fc0S+6R5dl9AcGAOaNXazuVmSTZPUb4r80dfpweQUoSHyQPHEc+6LK1xMWcSo8pu
U1dwBpGNFizy1/tS4/ePYE/0wJVEEyuKRLgcPce7YYDEYXsmOu+1ZZBd/m9OjFV0wdkmZpa7xb9O
v8QcGE4/rao80yj89ayvG+aPc+43uT3CAKW3p8UyddhC1I8x8AoyLtMoTAFALtdjsRI9IesnEMjv
QPHvO+tkT6VxK+JoFmZmpm8bNniYVYB0g4AEdXKXjnVf54K4FK/wUUR8hZb7qzOJlE5cu3+6gW3F
vaa1msuB0VlLvb5OxSOxEZeAWuNVjMYeZhkgZtDHaGA9iIJCA4CX3wY7h63ithsGJVxW9NAnc3e4
1YzJM7AvOlha9T1AoflW/MCfWAb4EAswxNGo1NP96BR+A2rl3zE61iG47Ww+aQnl765KNWq676Vd
cxgdBnNGZr/yc+3toU6hrjGV8q80Q039xufGc6RwTz7bNftXc+XmyhzqcixA0UlC7yZmupTCFuXh
BJmTChSm4NdyvXHRF7tRCWfRHvJVBFpVEInawbbETcPleVBSthgPtpVhuLi3QHSblRfOuBZTzdAw
Fd0dxdBJXnjWnxfjQG/uj2lvciro486LZHgCsuEdEIhtnC18k3J/upI2HsMzO1gcpfjuT/QwV7D7
qHG28hdQ8atYRupRG/53qwXPXnobG3C7Dws6FOUVfvffkN+L6zk4CRIIBz5Ldey99v+v+LmTRcZ1
3iSyVO6QTr2f6EWZlgSpbXr4S7k4SN7gco9Hxi7L9kbbQ3wEXZU3OPF9rWFQhMKIch9FEDsn5Cau
GfnjlBESadeIz3EHRMtYr1Rmbs4iF+dg6NAyj7QIiSCCtvc6d9EO0fZwiVFKCE5BHmhWomAFt+Ge
hKg/0uvSAeoy6oKNUs5faW3mkQCp4UZ/brvLEdDOpnc6Qldw2Ewwwiqf4jDUxs4CsSzLWxHlA+mi
YjOYzAfHsGprSb1GyV46S7HlLUHJn08FkWEwkUcioA3XttIz8Fdv0WSxelcZLxvijio92ait71gO
Kxk7ftRNVaPONRcxWPBF+nBHalxRlzSWSPU4qTZLvv94/GOnQIgZOSRQbMh68X8aKuU7xlB9QY8Q
yxONr9uZRHTVrdVPOvYZtVCYtVDzRoelTS9UO5UfrlrszzEY4/RaVjdUN6J95XD6JRFWrpi9Nbup
y0ZLJ1+SvTfIkuPURmi9QFhsADxOt6KAVOK1tYq0x3LqLs3nwDIwTMvwOiCiqUjPZb5AVNfvg8Bb
RQFS0C7LrAndgLkuT9yVmxBWsueVdrpZdCbIMZlLxiKJ+XHFg0kzq0UTbzDcYJ6ZNtF7e/M+hIqe
FRMcaRHT0NOTlC5WOLqajCo3lC4ConwxxjYdKpTIsKxWvCBKaJKndJHiJdafxq3GKAWjaR+o7JqA
QpgY5BNMVbpUfjUUxLshUkxLAW8MoVW6pe8+0NgavncGpfOrr0zt0a5pbK9w+iC/BG5lqg9XzDKn
n68BAGABNDS4OHluQTN1D+kmhDUvUw19anE0Q1g5vJa7vznFYPXE9HiH0mIT9oLbCmnlGyw67lAv
SfeeXKxx3SfVWVN1IGKvekc2jGjl8crnT3bgGYj29v0+T0JNwxMJGNpGX+XWFCWsokXOpxbfqcpy
OCqUYlZJ9ERWs9BVQ9FfYPNTJZ3Ey6C7S8vEWfXtPI8psoqHLj8WUcRBugWQuPALWX/zda2DpT+7
PHiZ7iada5iJEP5LDnYf+qqDb+2WJKoEoS1bpS1irqoBNqTOXaMWISEh02GZsrKSIn32lbmV/3jc
pjyTGAavUfiddUEp+bsTelkB+1PHl9EV6bXiG78w6rV/rCEqNs0Vy+xSHMYWWWRpDLufYgUcEILa
7Deb74/k6Hezds0v05MdP9yxI+s9oQu+dzyEJL2vgE/YAJEKB6KQWCKlpZVrqQd+XWNrTPGuh0Tb
27UP5f1zgAGiJyb1ASqGtoI5LvpYD7sgKZDsgRBCwVQgwHxHTIE3xv646MYxNiQKgrkX6n/RqCsg
PJ8hTlyonx8r5R1FzMKBFR/MTBQi0lljmUddO93RYdDVoraIwtGcJ7bxZxZnwQI4j/GbMPv9R3DI
y2l2owgiZs64LF6QbUDHADYKtuOv3GSRw5Wm+wjdiG5uNT1LLCYXWkDmma7OY47L+2SlAnyt3TqC
nHM5VUUtxXrP4fr3ZWkbgXEWctU+vrVNu3ZmEUVHFo+3tZe+BV23yLja+C5EIQqy+kmVRZ6KMnGi
SczJSiDyMHu7gMKkf7dR6HAeEuIu33A7581MsnRgMWLUa2okq4wTHSqyLDcgzqCGrQXjftLKF0TG
TpF6Bc5KPnnMi8NrGQ0BsM6EgC3pBtz+z4UWSayuIJRnjv88+25cyMbEnlIPw7IIJr3t3qwTH8PZ
KxFaXbziW8v9L7og9YB2coKXitHBniESqwoNkpa3aX3a7fDqgCeqVZIAcylD8+CCkFg2dm4pSecG
1n+el6Zz2K4kAX9Kl9t3hx31fh/VIurLRXCzoYtqvcmiHERawERlUrj0zxS9jtUkhBMz07PvWrAf
Y75kaVTvYVbAy5hoxA9j0Co49VzNYv7Cj2dNGjrKFeChtcnvCTmp8tuPghg4ObeQLbp+k5p1R0aK
ve9q+MwVkAxt5WhQj6VsxDRSK0yxI3RWopuI4Lk5v9iLt1c5z83u9ysx9rAk0UqX6caG/GE4Cf3c
yYekKjplZRrRFSenGb1kTv/gAvbgOhssMRTwiXX1YSjvHtoEdq3U6zcWJNvfreHkbwsYrtdXEylH
yY81FEnx3Th60SbSH9W2WFb5G26KHJ0fbVPId97ZkPEL0dcseJ39P5uPUHShzUBt4s85j9INYxQU
YnmPkaEl3q5eDeAQjBp8/o8QVGyg/GFUp6Hq/c8L76zbKpOBsC2wFCahnnMUxb5kAksNxQsteYsG
1HSVILI87hgsnMhR7sjoAPMGl1GuGMbPAGRGaZOfSEyHzQmwnpglBvNVLMKD64xES3tRw6zyeFva
J0nazTIXjte0ZH0qfUT7f0mD8GDVjcKlqVA9W3if4hiLTHB/zw9REuKnRnAyRTfFULFnvfPKBsY7
wv/rQxx45KRfWLQe153NHmFhC5b3BReQbJ5HQk7q7ewcH5HZYd6G3AXzFvZoHBfXZXLhNBg94LyR
icB/hX8EpCe5pz4N0g+g3U8PeiGSaLnWuiZylzXNUafY5DiuQnbDPNlngeJZsVrFWi/BXXSbXOFL
CkmhcSUwyKerCJfjtjLb9RrSE0+nQNe6m/Ax/VTGTB7d7EsfRXiaTbYabcdn08RaQO3mFQ/TJyvw
cHI/ixTnJQvdqU5IN38QEPVwAxt87CP8qKLfHwExSg5y5Skcd4mkvoNYJwiDU3DUCMipvw1V17og
uigcx5+58T5D+/Ng+hD1niiLghIZc2Qfg+K3zIuqmORQ9rebNyQHCYjl1EeAaFrSC3VXkaGVrgyx
PmtLcfv5xxJi2AW7BHbf6EFzQOuTLT5LR1tm5wwco3TNTU5ojwdSmYDCeocdlc6oJovcoU1KyxCs
z0wu6qOJ3O0Nqe/etEFT9ylrQjhEDvQ5UvCdSnEXEZcri47sxO3fs+cN23QGgZLo0viPmdEJFOE9
1G05iDAgJkFSPjjJvrJQbO+zukawppJ1Sn9cHvW1ZMttfJMrshT8U1DpATbkE6IPriWDSmQqjz1L
3Y1+xRZz6BY/LlLvGLsfqBmd5fn7TAhoZWaYh9F33L/IUCeV4WTIYTqKm8F+5fsGBEzHJGJYz/Vr
jPjK/QbpQMg6Lss1qgF1wqHAZFyFCY3DTLq2HGgPN6kWsL23+V5Wl25aoKu+S07WYzpphPu3PLBq
fQqBlFjHaaJJJqrUuv32/SNiLj859SCcQgQKAqTzd7TALfRuvSGadK6CPw7KWa7O/aT+6inujcZ/
TWqx26QwQGHe8fsqHA27JuaNlhLbrD0G17udDZoM43SnOJSu2+pFX2L9SaECuBdwHsMaryO+po7e
qYfh9D6gNbLwp3IzheDlaCcq9ZaHDbax+gZuuOifkdhxnTSASaVNy5HMIWri4kF5I0zprk4M9h4R
b5Z3PcuwCySa8of7Iks1USdMZtEVP9lIrfic3U9qAEjZL0ZJGeQ5FpfCQcyCqJ2J+clgvbwAsFNO
RAjL/S8n5gJbK8z+UhYeQ0O5g9tsaMDVlNANMXGTVL2o3cWeA+xZrduQsGg8x1n3k4X41OzEOmBj
4mDPgZG17TGH04HNDMXQ3HpilyY1HLxRe6mUq9gMQtADPXz5hSZjfSBGY/AxhS8VGMKsESSFOuAS
AOs7E0FMqF8BhKJ5L9zF/y1cdL1Q66a2tqLA6bULCaE6+ONbUpkGwaCU0z3mh2uV9BPb5jfBmWI7
lNwVPVEkNyDxd3SyINf+SUsao5etsFySyIbBdrMIgyxQokcEgLEOJYN7WlBvv1s6aoT/Bc0fCPnh
1bgsQlUMC0TQkAJa46gTNwVf1rNrCqKbsJPwv98iJ4VLvs2U/4tI338X9hR7KhUeshPZg4GUO5D0
xChsLDMKybYtpXPZIeszFpPM8VQcxOJkFPiHb0HLJo+q113eDi67u/bG2P4wVbPd7TLJBERqhiaC
uy5WKignsbaT9l48XOBy0hDVtmNbE3+1/8ltiC6uGGTLm4HMIsv0gVVT8O6dwjh7UZUKjeDF5xqA
Te8rrJ2umltnNFoHI0xEsspt6Mn3cduBZwRNPN9y8odxJCDcogzZRyx+1G04poc/cB3OeIj0SfND
xxB8mRkrW/2vOMIyhVrB3u+tfSFS6eo0+mKSMdyohLvVKtZdWCpqqM7UqHX7Tq4eb/DFoMhQ15kq
he/KxMAY7wrhCpKaApIuNRS21/qNuIlVYxDWBBUAhFUo42T1NVKRsUcSpZiK82se98jUh1FZTDz6
jQ0S8kkjpAN048kRbEIYVgnASzfic4Q5MEtuwpeaN1br24WBtikjhK4ZD6T+mfLb5lht1JNEd/7R
DgE0Ad5T2iernlsPMFLIp2njvCtzfDn7aLrCo8d09V+dJE1N6Qa9R9rOvTDkj1qMwTO/lFl2rOAx
Gsnl4O7X/LRhaeOVVre0BA2AJ/ywn1FX2/fDQ4vHzSWzv6sO6VDxkrUKupnw8c9R0UDFyzj405q4
IqeIeBTxXEtPkETcnYObsOvKNdgmeGm6bLzE7GafRRZg6EOblM/4z4zv4Gds2m26OqIilT+E36Nu
qaW19KwFAFBAr2ds7wA8ifz3GkdB/P3z1zuU4bBHWHXIbvnHNLnAOIV7F5QMjuqHz48zLr61WsWn
IcPeu6p+vHt4ajscQvO8l1SWS0/lsMJxzBsKkvCA6nso+0G71sdQsUM/TjqZ6ffwwe78yQ8YCnP+
5Lqc9qPsaMSSe53QZe5q8VS+eaaLXNmNXjGqd72vojVLk6ra5UZT90oAYwyRvWEFAFWqx/dIGjxt
qdxUVIx85v2TxS8DithJ4LrfYiw8v/uvp9dD3HNCd1YcdeXJ8qhJat/LVUENRu3eTSBMSKqGpu5B
B5h3Oq5LYYuSZFLkhnv9wclxgl1OjuRN4BI4RZ/YczaAtsy/lhsaj3rvAOUG/tuEKKqJu+XmXuzl
MU5oJOepED0zE9/bfupEGPYSDPkQcMet2ixSJtqcP17dMwiKeKT0pMemKCD1Ak3QBe1ht3PoKcZ4
rnDXv2siOTh5IBCI1NBOijL0XB9u2yOERBEDvRjYgTYUTFU8EEPdaNedpufMPRwglBuUtXqUln6H
l1pmnNxNO9wcYXZ1TGFop7+ezzDBAFheOz7/IXtHp1hforNX+mDg7UxqB4iKBL71QIx5QjhVYyeX
Ek86Z8UFFlIBMVEIDCqn4VFOGBzpMY2wMRMsRGiBO7vINqy6Y6DaQl+ktq9BQ1bpiBDxQADcrY44
6dq3bgrcPa0bqmorF6KnExdqXNG0D5UOvwXq8PwTDl6pcemuCGO087qaM9t0gMWq1NqIc3gS1ZTS
Q9FHwVG7dz5GQlewwMYl1rQSuPaHxpgTalUhHRLTFIXoSycZsqRMKDM57SvN3y/PfAftd8tEJ8IC
AZotxsWdb5Kjt3YsFqI4yuBBb2dy041+RGr+HTFUUUDXXw4XyKtotmnG4RRnGB3G++F1A88uxqg8
C2VYEeFyX2vwu8gKqQuQY5k0Q5CWd74wDeEBdZp4bPZl7hQE/Su3cWoN/O/sNg4eSYDiAbF5V6HZ
siI6Ao4c8AEJChmVzwURy1E98C+ybLxR+E6KO4jG6re0IFlwVVAYPMlb7BQSyoCYd9ivr+YAkorb
Ik3jvzQ6ouRu3r3nVYtvIJHcqpTRsWhOB0kpivIlYfuL2MCjr5t+cLa+g2PWiOpP14CBR1GXOPXp
Dk5Y7rzJo/6s0o1k1w5TGiMx3T86hP7HS20BTBTree715SmEdXXoN3GwVVnfwqmlcKGxvkCVsw41
6NhEGfFfkxjM9I5dapTVIIGtrdrqMSkCN2d4qiE1NyiN7TZHr1rEGiK9tpZmbEBYmT78XOeOV8Rf
tdUSc5xe0Hhum4UR0+foAjVSgvX69eNecq/5wSBsntm3i8xnuW7RjC1sI8MhFdPUO/0oXWkW9YKo
zM55xTHLrOTFcEIl+C+X3m0imtqlK263d/eEOjMrgCYjdKG0/qd7iYwMas+RGclBajY71rCGKUFE
JVyYS7tqVVxSMwoRq1e8SeNocXW6ExULLwP3ZK3ma+QMN8fjv0sPAkJ66c+tHSUl74TgPxC0atvQ
tsMP6x7d9I0sHX7UV86R6s+BO1Aau6GnHu49K1T4ams6acaDYb1YuEpAJ/M58NvqjHkPh+lxP39h
sYhSUNv00QeAoVsFsb270O3KDImCH6bRaCTHCnIFyEMSV1B9EeOSOfuOLMnAK3sWESHnWOOjJwZ8
aaSaqucokdod9l6VcHAvIgKK2gvRgW07cjjmQUg62FNpTC5pxzZ5VOVVXQ0AsLlXNGKJkEJpocdu
DCfhj9joVad+nKnVC0aJiz0Vsx2rrXBHRc8VFU6pvH00KYnoITAv0d7w5XBKWh/ofu+cIHlkuDiQ
7DqFPoy7nllSOcX52cgUL+CBtBFoOxEOLwyUkblY7QdnlTkbcUKpZpkklNnHYGFSX2AZIvqN7HWi
JVxd6SU/huaG+xjPpO/MRJHqbXRAAf8cYKPS2iHb6MvoRWd5S/ruVYTFz2ymL96HwbNjbzhW2uRN
kpb3+W2WSkVsAZ/uXtXpJolYcP1OnT5IOMSgl2oHGmaQdOE3uKRhuHRl2BCMv7AJqd/HJL4+f5/z
oS8shfsSCXdIDh47QiRlc3Pn1jQHPHRv5MXDs3Ek/69WN5XRJAlfpIlLqYY5+c5evdJMiiZo7IxI
lBMWAzTanSHrXMiwikNhQWV/a1kUiMbes5w2Be+fYNd9GYHA2PUDoMMXApe/BKWtWkWUbBH43X6m
BhRrx+ynlSIsPK0OCW3kbCkiZK7MS+RdOaNWZ/bxSIODnVc52xecn6U6JucElf8g3Tv5AWXb7ZTU
ZHtUUiqMpQQS8g+KqxiUjz2zJL8U7jYzs9/qDpwedbZG3FLk3Ux4Zscf/AXDgA1zOMfiwrBMFwck
JBOLxPaTttBK9Le5hNcGMNRFFXKFNG6kHyp/1TxHVHIH8XkPeqpQm9wp9ANtYnQAwhzkpMTs+1yW
EDeV2Sx1ojJOgqiPicEUWh5iZZ7jQoCyHhbtmOOc3KvTA2i77shVc20HZ2cgCp6ubEufZKgPejx4
WsjzEBf7SyCnkquHvbJi3a+hEWYgCNWEMRS1Y1OItJ2rK3e2KJwoeDuXzEoblrWTP5v2F3eoKd6H
A3KnAy+OYq7z+ORz0ItlwqdfG4JVVAM6xc+s1N5G+KrCdF2oycNsBAQlZW/38wUZb7rpqhnxgYOe
1SOigua2IYG2UyIMFOCABdj7PHvby3Yk1Vp3bMtmIVRJgc5AeCHTAgWvXX0KcqWjmJFhTbINfOEr
uR+Bfgv4touFACYZ9+oAvpM1aybrFX/lBVVZDF5+swEZPtnthnjWsV0Vv8aWMXAlP9KbQg4nLmtX
QihmqYjpWl2CUvVapslyjKWllxMfV1b24yTtwpA4QFu0SvoNXXL8JLMH6+XzGQrpHPzR0Cvoc4Eo
VbC8HAt/7+U5jf1xEpjtAv8KuIqE9G5gnXkB1FZI64+r+/HBZat1Gn22ZcM1l/Vvvr63cBzRhGVQ
NfciBY2GXMf34/JGc5Rg5NUggee+ElPMcQWkcIbGKEli3+K8sPHtZvMtDRdIxeNKFM3wj9KSZJmW
iRREoSc99YKbS2vz18B7B2jefEMVaUqNFSTj2JA1YlGQVx/Ph/rhuinkYX6qANAIxRLY8Byx4J9E
fB7aWo6mlAiYzNAnXcEOSWKQseatxhQhwc9Y/LNtRci+ys35gZLCHUbsDBVuC3JFmhJK6WY6o5ka
AFm+J8yIznt6GkepPq5ebGDrap6vC2eJOXXjvAqhdA+Yo/4kzmi2wO7tpi1uu1illS0w0H3p++GK
iO2kG61GBKyx3CRs6E8H4nX++zAxWGNI6duNDD09CYw/v7fzLNPuFvobzlI24z+oVCXrBcMIv7/k
vbR4lMGbwui9rlxk9Y1RnayrEA8TXUAgL+zMsawekJfCvK2F5koqDePs0T0be82qFKolVAyfONwF
ox0RwrXkwbjsPOcsKqyOy/ayfx+ul/5XLrtyHqOy1/xG+t/92VJYk+4kajbGrlAeCI+GZNusj/sY
O1JUHVLgJ6IwY6t7b+rosgjdnRlbYiaq3rme1r3dvnFlG9OKrFz1KiSAD4N/1zZx6tVVe1+Y2mP4
4jkSBBBQ3mR/kw9KnqftvGwObc7MXDOYGjZX/eqtOhpcYQb7COXW2S8t1qJk1Q2OrafxvxCdya8F
0KgMCoRN5jVb93qXWL9SURzvESgYlHh6ZAWQLmNdqvkV2INGHNa0Q/8GJOqmLw2Y0WILhBQE7gII
Oj1zIxUZSeLdumaoG4yCLlsTAJutGOyHIImQSmu+1AitlxVVVOOdLglWnN9c5uEzEv8QAsdeYA+1
hcwvpEQKX4v5cD0CevMbYx6TwauCHQvw6hf4Ok/8CFR0cC/4bGerltAg0HdLkS9PjrY1MkCudsAu
+RroY7jFoOACGmuls1awDpin75RE6KLktc2P0+T2KD/3PYa4ByAfVDYtY8uWWuyv1LqQkr41e+8D
96vkEyB8t5aeaEO1FSkutRBaG9NdzAN6EGmcZI4r5tnCe7g5ftXMXlBCfw37dhF78lS4rK/dNv0k
d6/p2qMTsR8MPJnx1/J7+oGpNuUetgOguesxA3AfuyDVfTr04oFC9BfChURcEbcsdYOkjG142cZa
a46hl9ASkOF1DywkYroae67thwY2mOlvND+WtHwBBuCRbZRKra/2ISuLYrbLm6Ztv5BL9NyGCRFM
8oM8xt9JCuZfKsYbfrZMdk8ZNmm0+yV8nBrroygIx/1UbFAP3O/gEZOqt+Jyg8PkG4bYgPROPW5E
G0BosdgeTnQFhjY3s0EGi6+VMokFPFgVmdjSlnb1871K+FsWHD7PUwdo8cM714q4DWfJdSCwfF5b
lIuLATRTyUhBB2wFGsk+QQ5Q3QmFVNd+iyNvkmnnM1EgubS7B32IuBSHjBjw3xY1ViqVPWtNifqY
wEJyDx6Qo10hAMCPWU5MK+20vqDU2agnIGn0+R6HiDYMclbCl3JWqul6jXCFcWmu/rUGnEAxmkXT
Q7issg59doWkxJpcWT0kPS/eLpcfXLXXYjXQ2CHnFkgie7C4+mcrMaMV8PupAW1U4nVxWkHXmkLP
FW5Iduu4exbsSF8DLbWN6NOg3YnMoIAjTbLl6kfnwINJEH9gFNnjqP8DlE63W+bwPxJZsQD6LprX
IBpcyT6SaODtF90cZKNf9U/US6qH6S3IaTmGvWTomiKHHPVS+dO6VqwZ1CV6KOalwMeOFO24xfBq
E8gQOesaNtUKrI9SIe/0hpI/dSHbp/zdciR39iJ+kP8xKipI9rPvL7Us+7Zx5GLgUxyQ8V6Xz9aN
bOVZ2xyIumZsyZJ16eCEpmkO6c/tKxjilGkDmx816BmmobY4s27vi/HMJh9peg6hlvMBjSKpLrtf
dPFDcXpoxFOauAA7x/EiD+gVKggmmuPW+PVEStZ2gx2Eo2Teh1GB8rWv/YzabWssA1WKVNYtQRvV
xc3iXXMm27ikAqcH1FYEX5xbXnNN+Pht5E0R7P9ZuSUAhp9AE0yxwgrWOQKpPqXAhtTG6onX222d
dgQf/NV2kCpyd3SiEb6aSjM6d6cT/ztWqgzXjum493a1gjG2osk8SwocuUBaWIEmT2q9g2qGRMqE
EYiXSmbBWTGpofwGXjFoXeOwmv53gMN3lZ8cEIp2UiBcigsYcYMoYZWpJleOMVB4bHDQR6SJo8eP
0vbeCJRC5ODRtRYc/fK1zizag37kKfFwbuRYdRiT4gYqCnflUEYOkQ7YhsFrX5jhSMSh4dMDUfdM
6QJ5/vfgl7raK7zZVQJouura9lWXjnJpw/g/Y0Cs9KhnhHGYlo5qMBnliNfwCfCIt/UtjE6LWGCb
70H+ArKcyVVXdHIFzLh6IhbQCxo/q3IqM3Y3vghKm9Y08SwPNeuBgxn9y/tXnTEj9Vr4c8QTISvJ
8f/YNzQX0wrdyR4xeXaV9xk2oxY5VBefeN3g1ceOKhDojR6HMIg00FMqSaxLg8gsxmZEHUbx0J+P
EKPRcdSg3jCj16u26sAxyE7pIo01s19vPE+XbQqGF6lHXeB/qk4c14qXOuDv0XM5275JCKEe2E3Z
+Z9E35t7u6GaCCZuNV+lIKUJwFK3PHxYnifd/15ehV2eA2PfibaGO8NTp3g/CBK2yrQPi3vzkwdJ
XucVhslwYStiaQ/ME9W7jmhhwJTKfeOeubVAesqkuFvqDQnsSkbUW9G9FHcCyof7yq8R6WW7DC9x
CdRMzY5hFJUwVBoKl1s9KkVT9jOh/P+RPu3TwRtYbzcZfML8No0DZZMRWLaRWlhHnqW+/S5WPRHf
Y0B+N6wU3UTl1nMwRZcomzUeCDbpqUrHAGRmvkpFMiHgU52ikYsN6Vo43FfVSUy5f1N13XBtYztt
36C7c40xpaKY1zDfHgwAZ49U8Qft+G3AdJefMCFhzr72SVxgXglzvaSepGUNgpiFFA/6PMQqASk5
8kwG4QozWXy+zxrdPfSwh2HB6Asm2x4id097eCgbQJses2MRj3VBkTqB7I2FBFs8/2wLgNB5xqYE
hRJhWg0NZEh4nQ618yNdsE5mYUJ7xNa62Z6SkBNADg6pb9KD9ru2nwGIPss4WpPkgcy9aPsR5oqC
ii53gXIA0gJ9Cd2g06/Km4ZW4YpOVA5WVuwPberczjJS9WgBGfLtYC4sWQpj3gSpDy71u4QsYGCR
0dvvyXbWfSH0Z1+8AznGrufofulg3W7ywLxJykO7zXuM2GCouF4rvAz5TBRyLFsmj+2lMlerpYPl
3jV2i+zgQeF1yJl8CkuFPXSKoqjct1eUWLt0k9GCyHwcuzSZ9D31YXb6ZBCsw8IR0tz0GEOTRqVl
cirIVGPnvgEWcuIp9GZRw/sarlpV6TjkXr5EOZ65xb5L/jGW+u+1CM8lRMM5ADCwUPREPCEROzkH
AbNlwwez6fOcdJKFuPgo8Don7I+OkJ1kEyOke8VPMxeDX1Q89BOzu06yn7YmUkgt8pEUV5wWCzz7
ZK78NvuV+FgRKuq39/PzURDJYRhHVTyQKTFe+1Hwjcyrl4kNTVy3Kl+JpTJYyauW7VA65FcgQpgC
UjIInOo48lmv7fIWVfm9b74jioWf2BahJqHh68/mwtwkg7IHZ7L4iMRdDxArFeRUEN6OAvGxlWn8
QmgjyNcS2/Oz+oF/p9cDAKLW/MXMTnguBGbuGCgxLulq1zw1VkemYXDXiN5oIIcBDRhI1FKyE7iZ
LC4r2eKzjsQ7iz6o6cQY8dUxTo5ZqpLzrTnykzWRoy0qLTel3q1D+XEbso4nhhdXLAkvXRRW3trp
btBQs6Fc87gBH0/bi/5x19bvo7K8rVLVZ5nn9RT0T29Q3ysuxC6co9GXLeBiOM5JdwNAnjjI8PCT
HmMxHRc4ihNzMYBweYOK8sVWnmp6XuudttTgoEYZmSUF7AQVZwW/8vs/Ngd9Npuzx7wQisYDaybl
WxTVTawMQsPT6eGeqJNmOD4oI1IEJg0ghbZfu+cfHPHVzwGA8/71MyHogf+pRU9bN2z/vpIx9jRn
VGna1pD9s6dJdgrLHn5v1gUwgNBZ4GKrJlhO0r4qnFw3dU5xyeBBjvGH7cQRBYJT687RbIdyhF3l
yWr+VoN9jdA4rvge6F/YzC4qSUACyY7QxkW1uazckyIcKi6/hKhQbQydyLYE95+JTFSRqBPOLiYs
YtHTyP7MM0ajLw64VDqlNMhJBiYNK3rJ+2eYU0ge/Wojgc9pCVA5+SWOaEqSBWbgHCRWFRANRMoQ
u9uhPfzFgrIVYBd94V3tw3hmNy4PrmFc4msfHNK1q8c0yJnACz1dxPO46nZIqHpJ250m8O9twzBz
xK+nOimDMmja0Sk67VG+I0UEgmkMiveZZklDH9dINV9oQtWq7NMbiSCMIEI5HDnwZL8hdmnSTf4D
pDerx247hcsvrioo5Fy5hPnXnlvqVrpTbAWyU6FCbrj7BkZMNHgkd7EocYywOXWDYLLgD7S0DIwu
1O+yr6RgfuYOkgng280u0wi9bse/cHYZv7J66Kf2G4UEGlwF60SPCepbWBpQofa43xJi1DY6gtJZ
+sXQSpHJTrL7auiAqsjdrl52qmPs9T+iZ08XEc2J+TEyJV9W92cNE7QdN0NCWE+za7WD/Ol2v5oF
wvygbSrt3YUIomOEx022YvQ959N2YAAqs1jXYRl1yj4uGOmvp0pXR8igy0ySlxfU4jjTWG3We9K8
14cfvKw+vwZ3xAAlcKQ5QWMaNyaPnVaAnHQG4JLl9iHtE6Flg8SbCLlvIvYxYGSTc6clE4qPrhpl
evYA63hCqXq6c255N4hijYSBNafpxM1R/cc6Cl/W5/M5dNiGMyr586155ZbkQdWLI5mAOiZybr/f
RiC2XBbs9V+a6ZYhY9Rsm/pzdC9fpiBYvZ3KC595Jwb+wEU+A/BB5SAZ8DKlWvzq+RIRkyZ0cNdh
Z+81s9o5mbSrPWVSXWLChyF8YJ9orFkaXIJseEpd2b7WOvgKb2w+NiBalsjCGW2VzQlt3H6K6LX8
iW7r1nEwWnuTyQJQOj0LBEJXdAHdKPEEObMnlMD0ELPIY+9PqEMWl+dLFBmXDLB/xWm2WSOYhFZ3
RQUgSrV6b991TCGMuKY8tu7cK18vnP4mrYrzpEpPpB/qaDBp37qneZrC9O5VgAdm9UfC++AzaNGW
4D3S+cpCN25an9eD5TRwBEhINMXkNpQop5cHM4Hj1/8YkjQYx6jup1HltsexILDdKWtYT2YqC0FH
+W0UDb9u+1TJItv/OMxWU9MZNqfgpXzwPVRxL6tkp2hHwmH6c2L1gR2cVuHWwUznsKxaQOOlbN8S
gGFaQ3JJBv027Xgcc9ef22iRAHteuufuyvIkLR+oEbXQ4nWCIDELnprV+/7qpYtH/BiPVEnByOhA
m1qMRd3pBiDWu5RsKuqtLwPDe16GlBwLHyhAY37BkjR9n9ZI0AGz9E2y3HlkOgzrfEM402e2X/OK
75mRuZX5dAFckXiEnRVPHqhskr6A8sGB8issuSbg58Ls77gazc9vtTH4dpapJcauCo3Pf0Eo1ERl
Rr5qaBdsCEf4nzvjIxJfZDk8wQiKQMY13VitBDjSQ+TmkgLqowJPnTmcnfLytm6Lh9ZIOc4WUb5X
njrWP4l8lBYl/mVE83Os4A07BjoDrr9hCsCP8p9HBRGJVjifRAzgQwhRZcG0tq6hRAJhTY5vM1KE
kpa5n6q/bBH8VLTjkm7d+j83FUDflhrE3MVhc6gRH7InPGtMZTaJrvACKejhGBvPMFCQ2cIthz9I
1nEPpvGxMk6/JcCbwtSKOFQ7bMqrWtZxt02XIig2MRuaTfop3LX7EF6ToDyt433cPlU7IMmRf/Cq
hX5w1uWArnSr+1F0q0asOi4jbORF0++RFg2leh1UqCSPVwtISBRIu/beoM/hE5pefFjTu323VDd4
GuEw47NkaseQPhUxhGzryjtWv1eBwoDdFd2LDzLE62wI1swha4q46niQaq3kxEJdP5MRAfTg/NHW
oFG3RRsXUekZzYkRwRWuO4Pkma0b4vyCAx7FMxJHUbyik9ZX1MtWgoTDv0cTr7mkvKQqk4ftWSaM
C9nCS1rXQZw3zg3gGSGPsYItyJqNjM539IZDyefX49nzKUPErPhPId0kiXfYZhripJgaAZVfI6xg
49vMvEM6o0aGQbKV/FAIj3ibc8ktXWuCECnuFMQr9OT21zIchQvkoL91Bpol5pxk1jeMpEoJM5zd
kzY3ZJFrGuCePMfqb84QQ30NzZOJspfa8sEstnD35FykyJ9za5rqfQCxTQCy2Z8MEsxrMbC/FXz+
PO5wAJXZXO0PUeVbV/bjrgQq3TZXWfVaKxhJKKOrSHxzfH0HJDxptOkdxNWglwdrY6kwSoG1kKwd
ZwwIoVHIfRM6pYMQ31tztunm3PpNTRueG7kyiZxJhr9dXHlfobqOg+cdxoEurmJ/o6vHFg+me255
dwRqRhaYezIJzcI+mc6Nlt7OdNa4/TdK3xno25hi8E8FShGPGE8UHfchXtJOjesocQCjK81q0E5t
WRJA25fGrA7Afe04/tDFMGBVu8dczdSJQEkdUVGE1k5pgXoY9ahwtaEya+zJ7J911bE6+iwHxf3B
r4lLPwcklkKy4Db3CefRr2OZZRI7t/46tm1Ky99h9sy/Qiwgki8ie1TyXqZkSL2Mmis3OVWHD03V
Ar2vZ4q++L6KSX9GmlorjKM4glAruNPEs0MqBV+DEO/isIcxqYj21zmG1XaJC0TlGUbyNpUDoCFZ
J8wBpdJ825sWcG3Azh4yZTdwY6iQIMVj0fRhUH3Q7o23BvMeXSklA7nEd3scmReXmx6Yff6pAA4k
BUjfkNeJD3vIqSanllnU+88VnHVUr9+Wn45QwxQz0YYCgU+KCVyiIb0S28u0AvVNl34O9+Ui4mNj
usNHkWPWG1B6x3sMWn38PmgE32xHXceP7Md1lCoQt6DBJtV0Yiu0KT5aI0pJJXFr1krwYLPuL/6E
Xv4ujg1UgZnvF5quKT0rdjAX6/1oNGeJKU62JglBzS+UJ9o+oL+KpopwqQ1bakaiZJcU2KP2DcAP
denXDUjfTv/dbOW2Dz+6qVGjXhIEZMleWRTFirCfs2fDclCKD/A5o7YqfXk2EA777w0RoPdI95IY
mDmsZlNLo43ZTcJw5pHmcZUS7jmyPUxOaboVNf/4Z0hk6d1hKjC/66IZA4oBbC5OX9jvGg0Jko+2
Vv79Goj2lE3g0tCJQmr5AUEifU0zE04LdmFbvD8D2TV39pZLvPSGMW5q1Z1HACdrMEhP10R4zCGS
S381SOXpGoSYtOcuwd5FPjQK2BqGEybhXqW6ALqU3yNt5gFmrP/QEYqQlE8wKLXWGwzDgwEfUwJC
9cFyWjwatK5nv5iKk0OVrc/1gR6FenytVs9M9b2Ovl735D8vpYVF4gZwaB0tRR4e1fnv5yuu02D2
KpxpCyPuvrFL2BBe2egUL21vhlK6/WyEGzZrOTguZASzJva93L91N1DwB+Nn/q5iKihczjBuwofR
SGW/SpjM7Lj6xUHxE7vFpo2eexVBr+KUjCDYUrET3s5BvFY0oZQQvE8FrXclQjPjdSDrAiMeYkdK
wlS+pC52UzeTbcqHzld7OW/4ipjbSQnknBwuHCXwcNA1h5ZTaXDNhB1agEViG8TSCZvZdP/ohP7o
bXZQdhEPviJDLe44++7tSgvHlU7XxgHyhZO4Lk5XtzKnrVPJE0k8nHUcloKKPL4VRExSfM56cytY
P7J+dfDu3XEBsOy+RI2vK9AGOh63QSo3kBKTZuy6PeWp4pu2P2SgadRlAgDOdbL4FX2o5NRquVeN
Rd4SiCOJqRUNkF4RkN0ED4gJY6N4ZNGBAS4B/AWZpTlvgkvVUfScCAP5FgdoxO762Qv0iA5coIxL
Q7gIvVrAPU4rN9jnfF6JU3nYpROxB4J8Soe4Aa6UrM5FisKlb+O7w/aclG/iXIVGW9jhYsWpQUJq
AHmCkzy1HdcYVfcMquxIDKyBGMF+1+hsCRpMoh01/NojWBgqImdTVPFL28W14DGjozlEvfyJbr2J
yfM2QIVjUxmQzIGFYTN0Vp1d0tZA1E0xqEf6aq4dPJlUfEO4meDZv1snDWIEYcosE4XzDh+PsspV
qkCvIYHyxYhK79BCYbRwz3p6HuywDL1qGF2xaDN9IbG52wjmZmoV2nP2fI3A0PazGcf+XhzUqWIv
XilknxoRcR4J/xrqAzDxU50y4ytUz0zS/oIPFqN399mRu/0324BvSz4C978/jHvcg2tm1D4ExcXl
wGNxXILJUnGRfDDw+761lIZrm35sTg8xu5mVMHCryIDWWf79jEvb3w1PYF/vADy/M7U3wWaoOEBg
9njEj6C7Spw8lCBdmbiJIoPE2oWKmsWZn/VHds60q4fIs/Nysa3a45IDXr3e5CbGo9kpOtqZb3w1
DIvGfIIa9bzmz2RCQtosIIGHR1inn9JMhiDNxNtaKMAGvh9jGXW9cp5jBIP33l+kDy8lTW3RBfmb
mxKvsKaGthNPBoTV2HDWR0VEwMjodtuE37Tu2HvtaivVGybBa0Wr+tj8onEToyGEA1Fb/Jjl3PAk
2wuviJlbdBvg9RjG+yh5UOtd9d1sYfV7RJ7k7lR1/MuMhCRUnC6icDe8l9jQBfZzFRI6+J2RFjW1
kmf4KczWOj1iVfVafLBevRKmtfGA6rAgh+OuNTebHpKB/z9jps8u2wBS6W3Pzl/lLf9cY+uahsGe
EHEh/9aRdy0Kuh1BJZBBRnuliDsb5bgaOMECSj2TDmg+bTCttzWVZL4o6q3Pf+cJCHt0cFSY8Wug
t7w5TQKWYbojeALlcy+yUeYXWKIfn4bqkiCSsJclDwGDzwi6x43SMk64zAhiibe4q4IPDZZJYMw3
NxqzQSJrY4CsV2rtWUnbEo+ihPaFgQM/s90URm9YTDKJVyavmCTn9/h2mmVSyGDjIJwvzp4V6BVF
wqtkE1z74+cv+PkrthlrBEqlkdNGO2/U+LWpbsGP9MOb/Vkucftayz9uElOHTzmkOmjICaRMQsfL
NSu+t36vxHlj+GU3WX2CbFUoz2vyWdVLPTgcJo7brsOGOn+FbPbUzqAvEETQ2grksttrVIXeTmMX
ocZ+bt3gzo+Q3cfzBZ6kiAk2+nTKH8Zl/juBFASVDLblL8GwoWyOWxH+ifM6sSfaWfGEuBJTDop6
jS2+zmXtfu843qytmf94VnnCD++0NpBj6xVbTsKECG8e12tri23aaPZNifytRlPppHHz0PawFmpN
8wvWai7W6VPbP5Hx6o5d2pcmNaYtmlB+90nz4UGnsa+DIeQ4cbiISpTFrtt1Z3uZxCiRqVamEVkg
FY9T+046NGsZmXfoMu59IaosjQHXTg8vwNM4cG7rmZGf7nXHhr2raOAFTMZHJ2kfwWNpmj2X8EjI
fsHIuu7BIq44oRrRt7DI6HWozsuZOFaJYm4LQ8Ng1lt0NMI7wY3wRjTrwNqp6PVJ/m/8txBSM6RO
F6QUrt8+aRxAP4ecbPaeWaYPVKWdbBHBhx5eOZjPH4phXbZyxbW1wrvPdDjqwwhr4RX1H7T3b46N
B3wkjdp7gdAGnikIn4B4mA0JRiN80a0enSTI5CFWYXjrLDPfzDNjJ+Xw+CVFiuZpquSAFJE7qVrV
DdDdnRwD/Htd+s2vnoemwW96P69qk5vrCBDDHjTPy6vB7waq6iaRTEfSPaL7GZQyYBA9V7HPUuC/
eOFPaAPiZTSkqy8co18hLT23H2MDFgBxNsyPzTaA4cvfpf9YVZyz+OG7Ep92Uk1dgV6K/uP8gObW
axu4Bavki+sBnYMm39drdMJdtf2y/FsxJcs6w+jXLnt+tDcL9anefps5eYK/OUuGYXaotijoT4dQ
DLquVzjoChiZGKFp7sZDoJ4D6219ntec42hpv716Wwyu8nLHC4LcmLxm//ZQO0m+r0ZgFiacJ4J0
wax57Y/FijRB0u0jTPz7PVghnOtS43kiZ5xuHZ1NP0ZOiCw7zyiYBT4gzKm2v7poxY41FQ8/sbQN
5gXPK39cGYGCfbQgVi5H0y4MieTf3d/k5FvU7O/F/Gi6AbfabslrPkWnJT7dAxA4pAliLmvL5QE3
3qw6lQ/FouAQB/O+jSAIbJf4IvjMbC8/NunDVpzao63hmHPFIvT2C9aVisepbPOOOQR2dvnSEILL
eXPT235uGlgE4FBi++ru0mHbI8NYA2HW5EtRzFPVMyBN1O/l2T+EbGb0ccARrxy3EjueBcAggw9g
k2pA6w8drsy0HfGQrnE1di0NeR6uyPBcTedt/8IAtZsKawu1nmPf+U9Ro3Fot+btjQEARaplj0Ls
oYWc4/ZpkF2eOmkv+oPsXRLfqTFJb4YMU/LsGz/6DI1hUA4z/6+e4x9Mm/y5RFItAIyF2frktwu/
dPhV/GusXkW8lGkeXB94sEsluQQYtOOfD0iiFQQzzhXIS98mQk0ziRAZEioA2oZmnu/WbaEZA+Yi
nbjDMXZS+EmDxWjGmgbR5eXxwAajOm1Wwk9YeXUia+9OR0QopKLhMf9v3XvZUiSGFDhaFCb7+TDl
SWsKu/aupf8GUxyrHP3VspP1wNhdFAzV59rzUDdPf4ypRYQf8Mejp0ded7XbEAiVYDC9R0ibib3f
zqQ97MUVfvoH5YonNpvO1UcSiaXtlKN3iuqTSrG98oAi6JH8059Ciqo1rWQqOkgR6d6EKDMC3uOu
dfajV/z4dt7hFEe1qZt0xdjqRZTE6xqddqT2NKfhfhV09pd0TdBYHok5mqFMBFvJAiP9JGh2KHJI
MhjcLlP2q2lm+MHmUd+aDAnWvMY6EPWkKZS6QAQ8w8yGpbLVy0td2RjKrWwPAOke6w9V4RkJ7PSK
cVblNT+Mb77F1UUl6BAz8U/jTq1l5eBNGrwRIQp8QWrvYkpLEFfGrk9AKgpasVf3JYN1MXnlSbFA
ptDE4kexWP4hZipEiPaYi5sOutyjqdkcl3VlkKxQsezFXkaRQoCHry1jVhn/eD54zwKKrdxafh9W
hBB7QYy3nEhqX1risyqAUrNdKcM8HPyJ2p5Y7w9URH+WJDps0r2ESVGJxWEhTMUuHh8njVujrXtO
UaDrVmulZQsfx2tajycSTzoEvrOEq1mLxqvPZwXc2DQwNgkQAh8X9StQrHIqG06sbSiGEchRFWt/
zwzjFyuwAyZqDyOctnCfUvzuMkCm/KIfoHS9x0gfslgg9WVprVVrLAwkDD/osNiS6dsCGCBZhjQf
42McYf1CQZysEf8akQISKRewlaPY6FjEeIbriUz/bTkx1RIBCatT5UOrFFoWaO9Uov1X2j7vJ2+C
SDyI2YtNWE11B7uoGoyXD5lrC7sRaTJevcd3t9KXhWu9MKqPG0gRDEhON3w2ppH5nwYjxnqXG7m6
9BPOXQ73bjKbYHLCcZBFUnKp1JUpYSnN8kgx/fzJOQILiuar8tlMq3Xs/Yt2zRkl6A5lqdHjcgZP
K065kolAWFvA2GiEBVWx4P8QqSsWa5D5lLCtb0muSzzV0v26t8aMdPOWV8a71848q7cZ/8MPXqiR
CLW9KLsCfkPbMTZtQI71KPnVNcvZ/ngmDVepUyB+GjmGSHCGX3eL0YIo0an1JrYk/bB7C8IsSmEf
7GoKGxLWxaA9lTvY2zc4yDNU36sukiyN6P2TD9yL10ZVNFRRssjYBSh4ppin/NqO5qn0qw5OwG+g
QtJSVmzQsVuYXkk/Xq3XDqLidRy3awAzsES/AqbLZu9XVAUC1MpHDP3vs7Xf9AnSqsODtIxGAzvU
Gk2+HXC+EjNxZsUabdrYTKUKea5tpdbJhdYJ7exd9YyIYBnX3x/A51LGQ7s9dbZjlLrx6ZIzafpo
qt2MAcw0GmCtpLw3dm9FwKtBskJtoqLrmD0L0QWi2Frn58bl1zWIoiRYvxc441WoN6HIR+PIcZn7
VQmbOLf+8j+anIMPVEcbtysASY3O2mVW1aZwxZ/XhDJVzwNOuOc7ZBBi7je4KLSyURVnfWt7GI5u
RHeuoobflbUxDNK4V/8NubtDL/Q28R0K/PKGhWqZgsUL5dICllKxguCNaD17G2eAaXXEnb6cjKe+
PqlkuQQq5zq/jRPyWf9KtKRx8AZEXkIBkeB4iOZieMYzrxpkrxNxOW3+KwKZhbcidTmkB4GVIqMb
z3ISoZPyhMgowB6bemH9/Bd44YS5DmqOgBpDRo+5yQ/dtduzTGOge/3CHjNo04g2UM8KGCUQLYqU
h1GW35rRzOmFhJNOzC0ubxLgMXudpzLFHVOTvBIFRufNJPWRPj0xKhW3698DHMw1/lyZCuWu5m3g
qiaSFiAJEZBZ8s9FalFImRaCoYiF1GQY8fujEif6sFjep/ne/p4MfuehAu+Je+PLAkxSGliL8v2V
RwqOCna7T0LqMh+2E0ydryL8QMBfbD8ePRbgt3158VaiBtgYXRnl8HqudZqwZ6JlvRweTmQbGS6U
ZjthEn1maggW2S4dkO5vSbyjKLNp8fdxuP10JrYKk08HJf0vXwNjh0rOFjaK9A5OEWmwmuXY7XZN
1fvsWGhlw3Cnb+eEgHix0J4i0hnoTHQk83NiFzQ+n3eg5rZsOL2vBh+urHntCDnOFNNYsItrTJGC
94wufBk82jHtKswI4zzTKK++TV/R2OstQLq+/09BFmNEtajPfOyVEhx9cbD3OrWnVqWx32YcoBez
1tq1K0FOmpK00oHQ6FuGM7Dg5XJf5nrM/ekNQdJ6iViCsCOr/a+M9ohtvOMIAiBNP8Ju6KxB6SaL
5MoZzwpzrto+8ehTwBSjpWlgAnnPujLggE8CNEDKketqlqrQ3HFtlNUDD0hAkSfSihezQVreisEV
YL3s1MpZ+zbVZ61NRgmGF3cbIcjszn764VUX4J5NI3FMRWSVk6u0KFkp16MYVT95QxTPSioENnP+
KeOQ6z7YEBbuWLEwWB81eX6SVRFztSqvpKaFEEficL3HUhvtsa2LKIdmYVSm0qMv5BjnzlUWvkd2
LKwNzIaEW7KON+cE0//w2qlWuUzO5M+6+tJs5FLdftMiU6r2ciLjGM98ElCaaNRKEW7+gULct2hv
xyNtAdurNSCCqCRRT/pQR4RiaHguMQr/DwMJg4H8fV1vpJZk29UruYiTDZxC8jhpZdWTSrFqZMtD
CZ0pzUiQCqJdMNSErHRJVijBIYiPt2JXU+AuR0Ui8Cu5Nu2Y6TYsNaV206ignM4xl5FWnDGrxl8b
fQ+lVtMdNoejFanMTvvascautSAConOj2aNWDdRcEEkpZCvd5UMuI32YIjQUWvnPHi1qonFx4sWE
2mY1hQ+HfV+5k7TxA7ebDodeyuRTUdHUnmFT4Hs5ibt1a2RWaqqMrvseb2e0pRLQ4c97+0rL2FEB
xwU/uxk1uxtHDlUXWzSjfh4NDmh6LYM8olDPpDoHcVfndk0oZPX3BSBNco01EmxUpwUDPZeURCA+
hfkRxSvjf/x56yOTJT+cQJl2j0p5MRdrQ37yRkezxEGJ0ch2AlsWeUauvuP1NXls9cH2iPWE4PYe
abDH5Evir8NRLDwX1iAJ80oA0g1f2RIXeU/FyGyvCFC84A9XUbAS02g0FjnQkxX/AqFlbgtvr7uG
tR1DFnu8jXgPlDI6qPncUhS0NEHhQwn8LRFw1b1JzU/EmdVazqNcMMmcaVmvOkK5FRvwU7ngFzTz
+MTyd+NcdqbThQOHHp3EB24By90U2uGWyCVPmW/c8AF3zPkrmCzcrfiVJ9B/E7oZ4JY0WiZXTHYj
INTkye1+rdI8InqVvKZPgurXccpG274fVZNDzZIuDrFo2ly88ok5Nh/+x2nAFd469V/IhH8/392Y
1eyzRiqnMezgPTh+Zs413KiIBvNks1kfjg6Y0mqMWaPRkm7DzJQibihxYHLcDPoxIELCtCQrDQKR
IAKtHO+bY3ffDXec6FDLgE9vw4KQtmQvJ0MWDsDH5PWbaPCeloVFDcpFCPNWeBWfbTEp+VSfScfC
JWw+skV952zZmYHXcrAmg7b/GN52UKGpvTBiTYWGTOYIUHHZH1+tVQzHFs0KBN3AXJndnD2l0ypW
JKFMPESV55C2j8fmy9G44+3CAew5TcV6jFSEUgRP4a5g3AkMalYcKUKQ2yjTtAcZw9qHNeMmue1j
AkDsHOQ6ssmK8A9R4PzqXTg8wUxJkw7QMnpTYEXPEmgbuMpS8epKzbsb0LcHsMi7Vup9SM0K3mXp
c2tW6INCP8dEc+FdRQ4YOk0qJVnQybwBUtlnj+lz3n2Bup80YlWON0iQBBZOH/pBiPQ51d7pen/I
tXzfW5ndkRHWYmq62tAe2982OUL+KmzPbQN07U4ed/jEDqMuJayRrHVyOncAv/kRERN4CMzcHWlj
ZCgzDte1DN6DyIxNZtc8Bt8yuxrcl2bU42PIQ77UpO8VjEx7OQKZXDIbdTtHNatAuKzc10SOiu9g
U79HsQLef8HUFqYZNZwc1T3tMDLTFn9wrB54qYJKdWADxRXzr0IXZCsaTUqXspvJDpHrXe7/SngW
k225CTq8eQS9+oj4C/e/4qW2gEwG5fHSvuyQulw8206cRW7zoZcIOuVrl6ylAHQigKcayHk+Ji37
jfNl4/u0P3fvFTrtm7WLOnADRYHRSYoY6X3k/WdeZyYUpfZA6SCyufVCIZnZruGUtFsrBl8bKn6V
6NNI4g29fYdq1FwPtH3i2AqgXzOXDCUNH5+peSCMbXlwxPWfrUUPOqUZG1QhC7jfYhel1AsBnQrg
KIqWU7RhyXwp4wROiv/wdrjbLPGKPEavBU5QO/fhpN1e5DwWgysm0NNmOVfTQKopkkJPk3wEyg5I
HMyMs7pk0p5Do0Cs3AXp83EAFj3ULc50vDyLqfgrNje5vsK6knD7Frx44SF2IkHygP9MDPqe9Oop
/X880MOcJRaK7Rog2npYeTkSbGkEw82IirWCk+pH7qJ5GZDDxw7z3gb0pe2txlgZwC9c60LVRu3J
IVaMM2k8ZZ3XNU0+lpA/R1jtuY41cyi3Dpmx1y1G46roR1zl1uugPwUemSLcNHYKvze+TC8JaLHH
sYDOOvTGw0/AjtO9uA1rT1tSe/6TpE+wB7+GJc6nZ4sXGXaPX5Ry/E/4siJ9XYyRGwKs6Tb6he3K
7WYuVqlYpqFLxJr3JRJx1ywIjDe7h2GAUDUxwN4zl6WHkjsKml+iNRublE0JQx78UmenoWXVmWbt
tPI5O2nZKbvyCt+TjsjbTEodL4eUJLWAQSLcJeNz7OGhBhK+Sayc7dXbKls3+eAbVC4FRcD6CvQ2
l5dCyN1pCbjXhOaj4wYVJ0oiclaZGw2LTn15LCU/Ma4HIL8EQEZ8b7yW2V/ZQUc1hsScS/GQF+6e
Ra5LTsbOvycJ1yAGWci4g/FKgz9jKtD7gJYNrC8b3d8ME1JNZXMb61odCUW/nnB6egtvaATwkX68
2gXXzrHujriKxv9gPIdB+xNxh+nKlkH1OAYn2YUp1HR5IhsuLsSCiEAqcGewCL1zfYTOUMIhLBqC
Ma1qfnnWpJhObwYEK5UXrscqw5jCPxcwVRV49qQM6Pjc3JNGaPN6w4Rr1Ec9qycAZFmAgUXj8bH0
JKzTsx66lE/tUL2bbd1+ULqfZO/Wcdu6d4HSsBKlL1NFD78uHJDypPWOuOf8vJG1Rz7qrpLoAQAO
HHLWmW4dm7U9TTWgERIHpYmPLasDQSBJHPr1tDPIRoIE4LANvd+fftWAcD83N/D8m+4RLGJgYV78
fmi8DHy+FJJm6qfDqaYODsWM/WYDEPxhxi8AM/XEF9QQrq7SyJXKYpHaHY+t4z/NV0Wh/B+dNpaI
9dMQk5FwGPLVHQuclQXml24p6lwg1LYW2qcCYkyBVNmtAidAiKQwBz73fq2M3UdDN7Y3yjNWdaMY
WT7tXW8Uv7QqbEYKlm+lvQngmTjCjR/8hrlEdE0fZqzIfYb1gmiEdMMnhJYBJwFZ+RWOqs++P2Df
u/AsGuhNAkw9BoZ6/tU4htVp6leNnKDz6ORw3pB5B8HGP1aJPa6J1ClqdsuknOgmRi8HsK16rTrz
RFWyh9WfT4YmsLUr3EN5fbiknlX3EYOPbhIvK0CIXPyeBIy2c5+Phe1XFuCXuzc/D2XAU23HRzAT
3JKGxjxcDdUyTTAsGi25jjuQKKExbrHgRnAm01TvTK1U3uTEQ1hWTyiqp7CWY2GFyTozsBfg1XH4
wKFGPnSGE0ebKXAaLRPJSyIQ9c02sENSwBFaymIi5Szp4oIqfomCjViU9TxK8FraoAAdjfCwgB2+
OMZ+CM1g9xv7IiEMNqtARBW6osCJvrAViHcdac3UxdEeQsH0047dGdFxEj5NItCWR4TTMS+LCZSr
kY87nlPS2O6THniW2y/AFb2YYNArTUtz3KALZj4ZpdJAWciLNK2rZzI2xzODSTottOsqLKXg5HCt
S4pjrr2VWEgQAcBITaoFFpZ7DA4dWDG8tF3hMdhRpxFsyA8Vv5w8Mag0II05RLGrERU8jd2Lra84
5LXsdojqhCbJ0nr/u7WuhRL++f6h3GLeMPyzrhUhauk2aUdx+gi+nffvuZtrXfZA4N9CgYq0jVU0
ioeJjoADQ/BuIpvS5zmFy85rlxtoDipHYXypNzzqv/mwV7wA5UxJ8QKNWrK9eB02NqSe9frHtB8Y
nWmp8WpRsa2ecHazmANqXGKs17Pz6XzRKFluCbFnKfBmWyexgvFGuF0QC+yraLxd1zwl8ABPOJyB
q8lF+GNFyveu3pkd1WYFu+5jLu2fe5oV7NhkuVa4q5Eib1dtnRU2SK2nIuEjot7h/jA18/P38NfO
AEZ1Jl4pVcD6d1rnvaAe77pEALPXvZBOM2CX7WVMcuY+gO1JP7+tRZNtY82hDlSwtQEaFkEZSskP
FO84euC/l2uOfJff7onieG6V9Ifvfg1ievkCA3aAdpzl/042V2lNS6bkBDtHBs9Q0ze5m/TSloQ9
5XQ01rSc4vrbJTeAPjPMbFwGYeAom8F2/pHTH3gGRYyf/r4u0cTWds3ZXgJPmeVq62mGSvMPlAl8
fMMrdYgUEQAwcknwgLT0qGZCAE553hqyGkMxuX7+R3x0X3ZCZMxVaO7hTiswuYLF7e7ayQEl9Bp9
9WLeLf08l0hWMjEbPtJhoM4ZEwyj1VbD6716VGXUpERjkyGBR0Bca+bafVHADbcKkcZS/eoY56/H
mcZhBDhEJTbZI+60eMPkeXkV8KNeXXGpDEoSLKMl4n4EHmQvlPip9HGGuxwUF6CO9UMgwrc9/ivm
kqPiXYOqLf59EkD2xB+ehcRsHbtXnS7z9QGOt8iamWqZUuiiahuvtGEVIRuGqUKnVpwE4RsVYPVI
pR55Jc1z74vYpgZnmwsj+tZXdOjIFjZjnTCNZDDx/ockK4aIazT9eKJPOKqKZOkjwCHUlBYqdU3B
KH9ouB32vvcvfPu7gYwg2KvGxo5xJbSC04aRfwq13WMwVhwrRWccFofbRICE9PWE6HNHPxZkYKUx
N4zd2t9d8hYm3i0fpz3Vs6EaY5nW1rU00UanZ4rJYwGY4xgTVSQfXDziQCrqsuL1MpU2c6lX5Cla
487RodlupyZC3TOKvNYFKSnHnIM9YvU63tunZTUagYBokkC6i8+FzZRD66ICWhEilSaGK/v3SngL
Ys4K9uX3Wj41Fp0wLXfPvEG53B5TbMWlPML+HpJfmuy9gvran2lrANJoI77hwaZrptDriHgkqnOg
mqDvnBG/t6SnMVypO0PQYsJ2TcQVyaPrnMc9tEXi8SIFjpwMxGpR3ke8YVuqkG2V6wmcSsnVjkKE
jR1u215HtcDrAvv4ejH1yoDSgLTgQizjB6jLXZ9jPu0lMtMwJeOCEZxhts1nVFgfrw8GskUbrZDx
ZOUlQuMxa0l6WVuq225WkQ8C2RESjkbefx298IFoMlgh52HUNlu5csdj6bfJYwnLUqyNkVTENYHt
MGbFnGk0Fi6mMrYioFZ+2VfeyXq3A+6JSYxG8VTKoCCI3bCq05/VXvYeGZORg0nHgGqBcR/rgFyY
dDQpLm9i3f7WRzJOe5FOzoyP3LZWff5shcIn9IKQsv8mMCXr/VEyqi40TH4ZCmX2aqMh4DMZNBxE
1k3WfEKmWDK1QXVIqcIzfJqnV5FaWa39gzx5mjvXRMrxoXFpX/+0oA6uuBDbsmw2/TzVXXSXw1Gp
Qs7unIrZyMJu3T0RZaNOuHJHZwNG3mA/JrUEw/u/yzT1e0Y/8wD3uUbxpllt5d8UaiUbmqhLiEhi
X4njkBTVqBVBYBc33FE9H/TxuAXkb97tbyZdRPk4qR1+QQWaVCIOmLNHKtZMxyhYU0FdGcNxVQjw
ySzOscO30vETZZAsgBjVJm7iZwhLBu6BtALb9F3yocwRJvfv84gBq43w1keWR/W33i2VTPEaffD8
AjdAssYN+f9fYMVq8Htcolf3NZM7KSYHcVsOF6+vKDUzQQ+JeTRXwXjpUuIUKEUYMWVRuKIKFOE6
M6Vueh/xHO4Lb3ExwKyMqpvjg8wjTPokDvyjEcNDOKtNgiR83cJJW1UW1/4SUeIdELeC+WDqJ95L
DCclhy2SbAvaR6HJS1UDVB1yw3xVNVEnFTnJ6ZC3uXDTRSDwSnnw3SrcYWs6UQcZiKmxB/SUtBZ3
qcIOfZcsRYSRFiMvT/L4K3Gg41pHcY5+9YiSwcCs6BNDc8kZLFPWBGl+roIdciOxJjDgWtiSUWrr
/0t0kea3KhHGOx8TEqJ4GO7TM97I8NCm6viICJt+Ssw53xaRhG/krmwxmKUP4rzDMl3z0rol7rem
s8Nv7n5eKjkwXUpA1/tx3unDvRKBsYsDDsu68DrnGhS+Ip199m2g/Xmi+T7GZ0pYIoocwF+64Muw
CqavYudF/1OCkQSNvRKeK3d7jyx6H+3QaQbcAx4K+8XHJerZYWxagiyoDDluemqMNy4QKomDJKp9
vFMdBhBjf0aPQ3YGWG7SlOUPvj3V0RZ3Gp14G1aDUbvrfx1bG6PwCV2DX8AsemTKka1uDqNC6uUk
rkE9IgWhBUUQn0+4imcGnOPQPlGWCCGn9O7Ne7aEO3cfZnLNrPsroPNRoTtoTWtB60gT5JBPZsej
kwduEwM3t/Cvw0Rt/9FFhibSqlIynycnczVS55ED4mxcud4Lc8IjUO/ZxtUH+Z9eU8Y3UvGmNxt3
bYX4pl7+Nyzj2ijzCBDgEcBlb4NG88xNpPaFSgCJEXO7LJUIOUGzeND9kiDX6vI19nPP7uAbAcOt
ez7LKEFQN8LzCClvCZcX8vRX9PRtTUxGjgrI1o7RU4KVQMWGaflckkMoZZBaESgkVJO6MS78zKU2
9d0r44/r7pjJZz7hNRINdfTCQPKCe20xFBCnInzyA7D+E6SgtnaXNYjXkOydfnzEaPEXGseInfYT
daAbWE0TXaTcNeRaR9mUGz1llaJtuJIPbR4yPb4w2yU1UNAiLQqr+1KZab4Q/+n7MPl86JRt0exV
xFR4L60JUOMAyW64wnA3gjtdMSZ1ayjdIrtAmBoBlFD0BptGDbIAp/CKzCecExjxW4gxkepCr9aM
/+7tV48SAfaT7IcTj7XxRGoEaWDPc+75mRW4GTbdS5Ej2hBoQY2xF4g1Dm5RShQy7Hqs2ytW/HX/
WMcKM7o5O1kQ75hz7FzDu7jX+c3QCtuv9JBsfgdIVrw5v58g7OOCbkXnYC/RLb2b/b8o0hMqwlo3
27RVuqT25hipXeQQT8jS1azwrBUMI3Q/rcgalfmqiUNR4rST47e4jT2G+ofItRpAGiGB1R1T2ofv
iBi63WgDT+q96MS3syRgvKrGg5j//5nPEFh0bycxALt7EJhyGOdqDRNuH2crLBmr4v/HhSL3ZV6q
uHsq6P/p2idXlGMB7otgn8E8bRqi7Gx5lKRdpse17yCZjaf2ryuqjCtfl/kwp+aSgImwl1aI+zG3
cOaqcKEo9U1hMUxRE76hBHCdaQ+dvynAUp+fhCUA05xfu4qrtbY1qscZmkoH9/xddTOgjhy1TO91
lvj19IacFgFLTYkpm1zsIMEPDhhBfs4C3O6HqWvyEKeDmNQxr7JfqZfJ0woIsoZHsS4zIzgWliE3
bvf3z6NxzBvtuT2bkhwNGshCB3QiwEIWkn/DmoiI4ZHKRZAaOr9EUoPX6L3LsB1UO3AHizP82T3g
dJn3HKX370Hc6FY/4VotOvTZ/RKLLIZ2Ysxz44R6J/yG5neLrNpZ4VVU0NpWfWwUrR5gKHxqjZ6Y
8AY9wOl8k6V6B8lngNGfOswz2yEBVZOmhCMZUlxLCgBZ2aHZE3y/3SxXh2e5Hwtpy+A4sU0VE3pB
GNbaw/N0cdLHvqiVfKsHVnsqVx0iD/lFidzgqwJ6neU3CoWRkvZ51MbbxTRIcjze4vdjEWwgso9E
IbBbC12bAq25Ex2n2vIUxJP/Fdsi5JisOIlVADcU11Sup41XnhFgDRpN00mRnHzZSjmRStW8irce
x1H9xrN+RV+HVrvdi/hZrjwHdNkbQ/Yjpta4a6a297mNS2fGFyjhrypMLz5pPlZFxHnI4FOW0dUl
ymGI2dKYoh9+f0zeK8RWvkNo2RNkmU/SM7SGD6mawQHqyfIcZQlyOqtViWGInLf0SVbkwFqC9KXV
T5BtAPxW+rFaMGdTseHvWBQ/dWnTWVETqgknWdoovxFoQ1ChKS30aTfL060IxRhPMUrAAr4TnII7
LqtHn7sm+Zb/jk1KusEUr+oxHh33+m7MfR40REgdl+QT8sE0SJMbx2Zt/hZTNfogZuX5077F85ke
mOCp7qTgsVSMz6yMnOECa+O2EwT73VA5DPtPzIVte/hrWFOmQvP+KoLjNg6UMV60DDj9lvMv/P37
6DAu8xiVEHulDEkAaNcWRwmLcIxp5iOrkzv8Xh11/nNZd+ieP/o7Lg1m04SZWC6TroU7UnIPfl2n
4OskOxhlqslaPmJudVk1yxh7O6mieYvwvbm2gER5eWMhOVptGPR/G7aO/feQmATuPQM4gIiCuHah
pFtoTNXIN2y/P0BS+ljdv0jTriv5LVtYb5PPBsASyK6jgH5UC69zufBmzqpJCwvhhA0z9o8nxGnl
K4Y+4bldBvWPj7H8/BawuV/DmtuLCb5SladZVwygycCkDy0XBBkFqwncv0Yei8tfWAOgfA/5ALam
wuWAaYA2Ybwxkb9X7bXY9ZZhMZ+bKZLty+xvJowO6syvp4ZIQIIJp8CaOS2BC2+vmhKA2btup6Vm
ubGU1hx1/YLGFL5rk9wF4LeB+Fy28JtAuiZWnGLtDuZnLQnWYKBSFFMwFBhWAqQkW8jeSuHyC8Ex
E1pIFwALUNTfbdaON3qccJuHZL/rtceAK7NFCTcdsAazZjwylP6aLWFbmFib6K5VloSHRMY6vsf6
ID3A7VujugJxvEsmV2p3QHA27Y2rTNkNNV1lR7/S+3BjMLwwLSPF3ObhLcCaQSReuGvTAFWngXI/
GNAO7uxmr1WeuuwzJO3znAIivqFzZhlcW6rJ5qkvfeZDU9V6u6w9YppT7e9TVDhRR8+jL6kyPTm8
h8VzrHAa9YbeNOPeKB0p2ynzrlVznjy1rWremnTl9iQsjs5iHYyolYwc+IOt9fU5Tr/anA1FDUhY
i+c2Om32Ed+hk6ZvXw1RExqHNZ0HG0vHChqHZhCDwqYpQcXhVmol0ShM4Leigy63ElzU5FDXtN0h
zT1iaT62OgNbGJSQar9lkCR62MhZqY/LIMtdQ1YLXs0kcGsT9sUYVpdKSdfcRxgVQflfOCT5PZ6y
UOQf2XBwfFKSStXLSCMyXe17HM28NV1trxe+/fgGUhrdL+/LnUwLKPo1xqYCaq2AQRwO3ukPza6d
9kqJxxDxanG2fQMfIZ5dIqT2dxlfyQc95+TC72qajIFchvKmxpJ8gBb5jCxFUDgqAouR/TaWegqo
1c3bkUadAnmz5QMXbZsaVljdieqPSHbnxMMuqRnl5j3Ca/viJuYgIHoPxGXQdl+dDhnAtdOaAWtn
4W+xOEhTJl12OkqrcShJw0fBrssQQrLh9sHhUwMA5x7svzHMm4o6/lV5bPhWl7UmhnnOm5WcOFgl
8ODnIKoH8o/X/zPAifXs/oKbYA7rLmhfkkcrQKiBUXsjWUa8t5ZOY6ZhuPwN+DE1VKgMZcVdy5fC
iyjxv1K4PlQxJ1Ob3Y7nLz+Q8kFjGHMOsxkwrFJu8+BCSlj1Yg7SuH3mwmY0bsjKB9vm9kGJ4rQl
/YriApYMigDykuliZtNd90fKJgnTo9PY+yr2NHxlSPmthDA3PGQUBlXZJUkWyYIXkdG4BFycwrCc
IB312fl/l8RWzg2xmdMbHo5ZxDReQbbnDoM5ERwtnwds3nEZjIOg9vk/NF2CFtsSbXkIALGxrm6Z
QIqJH2e/mgpZVdFslhUSgxbxWyg92e9CNMi9JSM+zQZd5UEWSS94c6AvaX6JOoGeatNHzj+BJ64X
AOCcbzN76x5D0LQnqTrpB6rvPvupfnSZlmJOPLP5qJUBmrk7VYpSCOBDZevIvgTS6gOQx0FoZ3mZ
PV6RXqpusoTNq+LJUlG450vKB+TCjR1wFysmEsMRUCx+Lubc7b4fZshvWPyCXh+AVZ6oZ/uV/hMo
KKrg9ZD8hFdiVFquPclomiR/z+jkCcIZp0TDDc0Zt2Wz89zpSEwXoDJEuoRXaznyv/cIP4di8uTq
tAJAAAzjpmBM2JumF1IbAeFGDqk0xlIOl1JkTCUv1QznJ1JyhE4vk77chBcoycFo3jA/mXgZLUTU
7wQ1mtgqNLJFExPv90h8V57bDEgzavGESaD6Dh3SERVIz0cK09XHNg5MAGadbcftNmBciy/NX65n
+19/QSL/tQpm8CVevb0otW98zPp9eELl4j6RPkc5yAmMI5JwQYgpd/PRbzl9XXG1aJci8VZLyDTb
VKRIQkzCPl+pL5zobkBNNT42w0AN/GpqcKU+pSdZ4gbkCDZPl4rgtNFmLijRymACLeOTcSscdJQc
RFsTJ9Wgyl2+pNHDxeen1L6tYtyRcyYlYjFpCVdwF8Un5jn8d/ZIsDTaCkaaYAyOrdBG6jij5Nl8
BcUItjr8yJli+eZowPxSuY2WMj8SD8Bc5dfaaXut8ISj3u4LRM5I9jXBpdxn6u2r7nuUHDz18wUo
rHKMWq69RkI5WYEam5moDGtsED0Ny/FoJbSkgAJ3jfEwvEUbSckycNrCo0l5LxjVSBM9x5oTNiRg
G5rpL071ZXGTIQGEW8hSROat1y6k/oV5t1GBw9FhlIcFYMR3D5JcQ68eXB6INPOSTaw0/aCtNGA8
btaRJJoIYlMfGfm0y6rRjJOub1PhX7JwdkZO3NTGBtQJhrbV8O5HwJ1UFP1+eI9cumX6Bf7WrRcX
m2xnfaYzeDZKiu9QidMOJsBKJfq9fuenY5AkjvqkMIUMAGYS5lH3yyIImk0prkBM3PEYs5vPZ1Fl
lDMf6fEM9UAKoekKo/IyrFFNaUQNa5bd/Px53ofowaFy0psQyZPAikQbXIg+FHbc2ym6nFOksCBW
SMmFixTemuiS7sfqRldTV8iaiVbOCtVTPJbrEzTb38jWAHZPLoTgexMokySzA6TB/dgarI3axYVB
siHloe1pvr7QMhX2bTc7VFAvSw7/O6AV4q2hcHf+Mf/EvEhfGjCiesIIsUiHs5W20bOLAEN50fV8
RgeVomsEikbKrkT6eHSqq1tVN99DuWwnKsGGGgxPVZvgWBZDBnMHthmhFoDXvfyn9B/thSEGcWeX
XMmsBQGtxvkIP/BPinwCCgA+M8Ycvubzl8ua4RjEgZrkHWvM3OgHSFQT2vfGLH4qe/4NsBS5Fe5z
fynfHq39/B77UAULdGIFEBwCTsVfHRVn4EXkgRgFn8ae2xD5C7Z9GEGb3LhPM5NvKMKx+qffgxlG
HE6FYYsdeLS9nH82GLSnei8wFX/3iW4b8iHrjiYaI1xydL+llFPquOcmvqiFqYuyJMB/Lv6jDYhf
eD/DsmOaqG0S77xtzmp39LLgLhA+fDY+E9jmMgvQUGmZjK+28tPHFVERt5PW3qVOpXMiqWcgfm+V
FVYtiKW1qBsjjgj7OfaU5eRNBsCqc4JipQiGCnkrYe7ooglx09tsanhZ739DMlR954rnvZvUyunL
bjdJIbaroGXW9tpTYnLjs2NN/JKulRB1+KWDQUq65G04Z+VnmSmnn0E3wwfSckql36fy/r/l76DK
GSf5lPK+Aqmy0d4EDw+2KXgyQTvd1v8fXOElo/ojpXSedESaEBsfWeNShfekMUN6tpYHpaCPJ9G2
9T6MavoEd4s0NMazOmlgMT+kttQBuUncQkJFI4v3h5/ZhqkibIuMICJEfeMHNxND+9kthLXZNNvs
AOM093K+7PkvXVFTQ33IrmLRFJ0NDrAIS/RykghjjxXsNMLScn5VcEUg+G1GHmcqvtivYLgBEyWp
w7r2gxehM0B/V/gdp0t6HtauiW513Rm4siGVv28P29nO6tRnscGkGfFrEXfkb6N0I0QxuCbBxSUT
ZEV26PocKYA6Z2Rc5dvm8x8Bp3UccZeOsNL2wPHJnc+QmWcopzXdVxT12voOPXjoGSf38xbxSZ0b
pBl/fJ0XPC8o8RKRzBkd2qoYaFsqbkbSrQ5OZFHGH08ETXBdjdSU6evIUE/rgWxLggDCTHfsVlW8
K58hAk+dMneGEB5p2jm2WL8k+drmK0VlEQ8+JEHTm6aT28rZVgzCWRYzjvsy8k0cHK4EvXPlmKps
wO7qcdYLn2opEq66NBTS2PuIQngMmyIiMogNuvJLB5MRCk6NSymfWDF4akyyL4AomnxXrcVyT1Iu
0TMYGlKF73R/hGh+Lm/52nk5sPD1mZyrQu6ruCVMxrkACPkyGrcgYgEY1UdfnV/4+7/BvBw3ynIp
BwcqwCG9gtqoj0mLLyGh+vf0vFi1756Fo1f9rc0v1NmXlKvuFBLhT5WeMqtACkzDj2jm3WRLk7Ym
6GvdYDthlL98Vrm/X3bgC83yY4ycgrNRHKg9X8Gu2zhX+mUWr0PUcP0FOKFlFnX0vQ9iFhbSRdH5
XORGEuq3OkFxgDxDWdLwnbF+JTsoRHOvFOYDDW+zaKl7UwnYD6pLxRbG8lhQg6G68LZ6qGOyu6U2
SoDnob10pSegkXrxq/cYOZ8quMJG5gjyyxbE2eYR5YNFHUWSIPcl1lHD8MiFEdNQlWWdNt0D/NU7
fxWmvUUDwvE/eYSXTfeZZByQLuBlhTuHvWnRMItmusm7EO+YKbuidtvbJk1m/Qf1UrVkSx+3JM+T
4e/AaoZ1nc1aZ8QN9LZKCh+hmXqyurLm54HswmB71eLT2KJyMGCwffQiOyCR8RKF0J5FB/73dvl3
bYXjSjePj8gQiMPggKoWwQThY8P99uTsy0TGajqAxNsDPl7351vhK6YrVg+LuotFoiQVfws5RBX9
LY2ySez7tvEEAN9z/sxA4HSWZlBLMSAtMFnhFWHzKp7NQflpOKd/1kf3F4auORDUjs2aBMqNAvox
/w9oJilH6GX+vLLQ+WeXNuka4QFENyx1CV2gKmKjLNyIV7cXbbjPQGHdX2Oi46Ifsf8PsZeYrtmL
3Kbpm+HJzHuUtebDD7PdgT0yporLoRDyfjrkgfEI6KUUYgzMt2pWVa4IkdRfCOt+xu0r8zWAWREb
x+RvednhozXodeNdCJ7CYMVY0c9duT8QHDCZJJYXGQAivwpBwF0PzegXryNZpLLGDUvSc7uUI+xQ
BJ+XZZd7mAVinS638otSbVkqXmMcqLkE8KExqsZbftfWDW9tP5Y0uaOH84160yK7bo1iTECDgyFT
elfYwzh4D2YvXUET/EAj058uirsgNsc6dSZgWRwMwVw791sYl8gRcMgDhAWSxp9fwdwwq+bM4mYz
bBpnNPLTNnxH5LWuqOdnYpMvzzLm8NTk5DyxseX9VJAyKKCefcPOhN+DuNlxtyx9nOWAzVA+MrMo
zJ/+felMznxCXXlrFbpeszwycFCFp0ySPsNpVMIqP0ViqWcHaIQBYXV4ebjmQ5/6O+wcAKeNryhv
cleEp7+Ovna/U/3trLGgh+29l23AVoOc2eOqeHS0C6f7rVA42mXCDwOnswF82pvHkSBI7l87iLlb
m+REt1Lt9jpJJkh9l/tT1lCI5RrXbex1u7OT6EgAN+IMcC6wlnjWMMOeElvKZ6tvyK/F85MRdPEr
8Wcy9xGl60A5pAIp2775m0uOSlqUbCXP/XTKvkPk2qIB3+Wl4Kor+ToQW1m2H1+1f56TkO1pEz/m
amRgLb29QJfDQqsHV5i2XWowWaMIMGE7ZbY7UFETo/7Sd/IAXiuyKZ9Lf1Il6PO51AN7s4hgrLL/
5/IQfxnsx+Qvd8gh+gIaTyjfuQKY5JIV9sLW+sTjc8WesSk3Y3Do21Fo6NwkSsIDbEXzhfC64pvT
cQslC7y41aXFvj63ziqmFbv3HfPQhWlcer1NfVaRk0mPhDDmlfXIZXLB3X3lAmHQ+4TKF9/nyCgs
frjFhWyjnkSLcpbYOKuosqIUSV3jh2zmWmSzGlkw4xN8Bk8FNWvRj6mzj0NxXQdgx5spXRjZSTRy
NBAV8IOcqUEqlVojSpiUtjC0xNpRkvRIrhS4F1OAXErwqzXNzu5Gjb1SP1N8k2B8ww5oN9tJu+yu
852HSkzSvcBbWfEVGyEc9mN4G3aTqYdaGxZ4BkF47ni1w69XE68ADoJkUEPYo7CBdNBowcyi0x7o
dM8KNE0uABJI6ujRNOSC80GxDhXxlcNR0mtxRThNVPncQUTPHPnqaSKw7fTlJorDA/lWHfbIjD3k
g1mCCBfSMCdp6H7iZWwmz+K8pjcP5dDbBFDKlohnwUsOesPIO8i0I3wMtG4U+bQSn5XZrH0zIvTo
LMJECdX/LLk3SMMV7H/Jdga7T+FHnyI9A3+k0WB0fc5aca9mVZoHmEIHv2qfysQpgwB7h3DQ0MjX
q/8l+5iWH2cgEzND0fySlvMcwkyeFOESqEEPy3Jw6Rs4SO7RyeqFum+PSvqk1WbJYfwcGQgYF6lr
eSJ0t7Ftumgd9VTFU9c5ZGE6F00Ksvw7iZyqon0CKUQ/e8/QszAcAoTZ8sEUQIsREw0Gq/qJVp5B
OMWkPxn4QbpfecNE4WwEU8Y+ucS8IRNovltym5izcE/PkjJ1QxziZniBP3yQ9fStRrvCGI9iHdY0
UIfaML35Lf+Fs0e/ZaEn8UPnP5GTRPDSlYP/UAa8Dhb6+ub8zA4S+1rzo7LhJLuBeO7hYYcaRU4J
U+j6SS8xFujxRJ6jd156YIHBstsofNIWOQ7MmEdyWFkTEx/VvXsA0sXc/XS9woUqSdNSLLJ5smb0
R/k8nDqEfLEKVuXrJs8J4vYmsyiSdsR/5n9RWNBg3SMIPS79hgt5B3qEpiLhmMSGhao4Gau1lh+A
v0MmD5R74bH2wc1Z1sG2Yu/dIEDBWo7YkZ2Rhqfaq0uQKqcXAbLojy46yxwQt+/8oGQdIbwoBfpH
LbKrTUKV3BpLreIO0y7K82pjqrWZ6uvl90lDiQA5vQ7gQXufwsV9RRFVpA1YGvWr5Bj5OGVqRxGV
KckGt+B5wUkQM6S7yaRmicAhvoahYlQ0dhNLcymsjSYj5SSH3AC80VsIYfxzoEmeRYB4fKAWVZux
lQimy2ExXff1HD9Kxcv3g1Dl/jlzYFWayzzK/APGNc8OkG5N729HDq8f8yOOrrc5rF/pIcvbjcvX
hCOnzCRFl3c2XZFK9CzTjGI49GZTz15V1q6LbIy8ge5Y2injFKgcreuRhXS2+bdLAO3PLlYckXCH
mrDaQX/DCWl6X9xY7cx9S1h83kwXTuQaupIlWhy+i0/TeEaj5ldLnTYSIEYC91ZheGtgsUHc8JNh
QkYrxO4UsDIR8Bw1V9GQMdTBXYu2LyrVXjYvccXlRZLyW0oCRhOYpdsq6eoEOI5nzzFKwvcJMVRN
2lbgszA93vgcq2TDCW7frXRnHegSAxbgnMzRUhwC2gBgZxTbe3MXKgo0RK8B4qs+jY6T4plUCEiN
m7kj7rqk5Iba76OX7u3a0C+wf8o/aPGxYCh2lBZ+4DC11uQMRAtup6GJSwoMPIBazTivJJ+QpYNU
ecPDLpfPFPtYDrF/Xs154z54GY2H8Tqi6By67fIEXxAOkEcpVIAU1BXonjynq0eMS2bAvnpzKiZS
hwNUEhY4Nr4ppWTmNZRu4uFCgj4DI+dNWbkRnOHWbv2hdjvNW5cDa+3S1HdwbZrjBQfwy7TSSdvP
QoZZDFqKXl0EllK71m2eHrHS/97oDBm7ygwhCddCCoIH81AZPvgk6DCmebC1Yy9pqLm2Geb+4mEr
JdXypYQIGA/oJuytlJCBeDo6Nb5qFGRvabEnWj50cGfXFcONFLHOXChi/42WBHRuSi3txpOIPJ27
QaMH23g3kXnYBJNh7xwC5+xUoVaX87EHTqmGfBKmSmEF45TyZkrpOBmXOxmyncUUkysDLQbkmJA1
1ueUVH+Njb/fhxldAWzYJ2IlQR0KfKygEYHIzuxtXK7UCpu3/QCRNOCr5eqD6VKRlIEw76ktJ76q
3RR04Vg/g9xzuqg+8CwXeYohUXUOyurIB++cQSJAdj1lyYWCxZ8+U8WcRi3lTzKh058+6BXXgP6U
K8nG6kGdK2jk4p/o+guR7XUGT31hmkgaMKIzWXsQqEs4WjtDU2wywJQb0bg8XqlrmX7Zvn1YaOXc
CJnSEmm3kxurjMFSzGxOlCc470X1oXFKaqWOEfImQPve2RUOMnhE00tIXE6MKgOBMhApizKQl8fc
RLjOUlIm5SDQm6YFScsMDtlwnJIVkd8GunazKcEaVVUCqOa1s7g+CfV4gRh6WFrUzM9OtO83wu+B
ifPh4QLJ1q60yHgBMBaZbLaf7vVtmPwGwJOMvCu/1q4E+s9XaVRbBLZ+gWzUdbhy+KoQFOpsbYOX
QeGYAlL2dO51u2C+pSGMu7GKOLtrhSKDyUNGr/LEroAglNjSg9KJE6MndDOIUxrW5DzjdVnmub6o
FEuEKyhLsuy+IFPO5S3BwOqDjmnREjdYw/cYCjYjOQ1oCeU3W/46ELPWOiiLK03wcVo1hU4danAI
u2IFH6d7CeXTKyvAm9JLNzmYVCNl9BP3XQ0tRDR7ZUrFq8ffTstk2DAi9zGnTmIOR3DJLqQxJDo7
dUaJam1BWR98wjPYRyGwGhfPic+qWrk2Pd1P/Z8YJYXvH8AZdvKbWLF2eJdQkTSGg3v98Ogs4qHz
q1y3G/6XAQ/6PuEFHyX11zv1EcvIHRPuCtIypHBUj1RE2DfQyQbkCi9bzOWlkfBpxPMt3wMulBMQ
T+BI/1qJGbEZ/jU3M4Swnf6XYzBQCNzTjb+VWRfDcgRL3hvg5Kw+ltWnBiCiFb0J6RkFZ9/ATJAC
AiU1cikIARpc7d/jN12jYwHthhbXGCppXJIRW7p6J2rF6GAlXtr27fygiocx6Gb9T+r5G/P9EbiX
fN1CiczfhiGeUVKkwDLMQo0y1mW9/uA4BQjS1nJmCdjWRua1nidpx1R8pyaZuhNzyFAVRjC97AgY
35IveLHbuPrqs/NYmBs5wyD45X+URtA1S1XKpo0yb8oE+gCDMjX3W3ot7hlxqtmN3zNsd5pCPqxG
NFAUv3mws//n44Hu0Ik1OYS35Z5lwI27wsUhKn88eg8mH/eXorK/4HYml4r6fCGDJWeERtsDkfCw
bKVIa+86UVudIWtxOLYklanQrKjh7nolJRqhSV3bokMCoDTQRCTXYdpUIXvds85XmywThjrk0928
9u6n0joN18bZWeW5+5kJ7kd5Un0jWIoueor6QfJn1b5/l2ZH3kgqSbPct1v2SC8njoeRTdYNdWLi
DxZWpHlgs7yq7E57RykFMPxFKjuwWUmsoswEWbZ9TBJtVe7+9gAggNML22CEim53Ww+3/k5q3E2f
yC9AZpCua/C9RytBx/woVLpvdbWdesG6jAmCt8S0wJtq+CqZmcJ1TacNawRodcfFOh8g/wnNVYeN
KgFJFl+0vNu0ob66ftyiNcYL7V0+1sD9kwaO6ji7GgMeDa/JkG2Q9DiviqzrdHQuf7LPyrUPHz58
MqIIKs4mdVyKZkTADdlT+MeCHLMprJu/YVhgzr641iWx02/UcmacnNXV43lSj2mHCIjArjdACNQJ
eTya+D1wH/lVLBmYq2QNrjFiRfOGG/qB4X5KDkYrcjpsZi7OdTkt9AY7KNN7NVVv5A0zQLMUI/XQ
rwaCbqMA/lvnAsUpzWlmC24ZO2fvXxefUHcRL5+jdmgEi1QsVLXo/NVMSuPw85curXgVRH0u3qvF
cwNRxGrGD5iIv1VwmEtNAIKYp/IeCpo6NMX8zHYhMo16Kzka87ep8uolR41yluF2gGGGVGHQVS97
wiFHkaDWWf6Ul/aQ0gZC1u/63EA1d0dAQhCqnbbgc52zbDMOtTh9pGdMgRaymbmlm48KuOw70oyy
xIKyJCM6ScoVG82WkhmhGzUMIe3gBHz9nTOHYW8cWjK/S+YlgDfymm3j2P4Z3Y7iQUa1a4pjc7zS
O0chI/yjz74qpI4GyW5Bsvo3gDSk7GSoiPk1zh+iiZ5lmDjNArIBjZuLS8jPzk5GBz6mPUUchDtE
+5r3wupYDOWdmiylMyimcUZ0fAXqk1hLklFwbUHVG4aNv64OqTiph9xTlm+IHeOxSzIhJHpfKh9T
e8g33ApY9gAqhxryjLhjh0p042Y7yc6V2aa22LR3sMbhJk4e4wXz5XBzZ53yzNQS5VTM4j2kzmUC
RUEDRIC0azwtU6Y+2xmhMh0dgUQVqNpCZC/Dk9oi01GnjQfpDIcvPazb8sAcFW2rhE1LnWsU26bA
dd6jfT/1lruc/GmOzveRDqgPl+oE8mIN6f1VFTfvDGcFZ2vMPQrjD6u1oRUfWIaLL45dSkHpmNle
7iraTZ5bbhY9OKiFMnyoKPBZLWH2GDtK76y6QHOJdOPIAFMmoKn0BhDeHOl2YRvacjCVAAzfcw9s
qGyVL4Nl2bNZ0ykurzpu2t+d5N/uimYJ0+nglqDrroFfICoj0XfT+qhejMPS4VoOvhTFg223+HQK
XDt0mnrsQyfiexCVuhGKSdkR6z6lAKW/LNmY5QLVK/AZWg/wgQV2NUH0inMAqwZd0SLjMUTOo2me
UpR1yx7f0D+A1mlqrzEkndWqz4iP/wso83bq6jetZleKIVDOYjPw76jKLXy0lgJxkjzkuvEmBpE1
/Aq+aMP+GCikFhurP6Ap02TQp3/opKMVbqFv1vKCWH+egkc9vbA0xqzhRsG7huIq4WAPCjy7Cp4Q
DO0PQuwJEZHbJJz9valy5m95rjvkJAS4nmoJfDo/SQl3hnSWWQzD+/I1eT2ajWgYphvlgen9ku24
v0iGgRJ/PGHg/kUFY/OeaVn8tdwOk85BFV4OUFAaHEQaxVtP0UfKeuCLKQrCR1vOkfI4pXFEo7c4
61dD7Kkw8SQd0ycloDeIk5tbDwHkPhsX7ZM2m+rYtJF3xNi7CH0feOrBcYiBos62YJMHdBoP4jKR
HJw9r6rGT6GkEgeENqm7h0RN0AS22tbX22nCvOjrEj0wWZN+U6Ju429yd1b8+6tMBJhZUEDIFMb8
J4+kEqyIBu6vWF5mftg9NtB0C/qXoGr4kq+/8Q5QcHOBV9iKNIod32GwN1/r/tAQY5saorUF3G6K
YegNoW5JuO3ugG5xn1wP9y6t57vnysTnzKoNQa7vI9fio0nXZwS7ng4E2YsQIZq5i9bsyv0o4EKt
UWeVNv+4tG42Vuer3k6ltiASZajSFKyQZf9KrIoixBrmZpn/Ie+MhzfyHl5sJskWPJzn0GVGHAd3
0QaU4GdTzxfzN9Zp3Mw0ReNTK8Ib+kkcpWyOU3xQ/SsbvPjZFV3trU2+3mYej+6pMNH50glX8emU
CFbb1kcC0zwtezX8PKx/949JFQuSmxscMDTRl2XUw2xHAmFcA+sJPYSoMXA/BDwSRduo3kY31wIy
qFgCBy5QhuMjbtZJMM43HiWwWZqMBRniVWDm5Ff9dW8X3fTq/WfnMg7nzwSxMbe9EgGqTd87jxSh
dVbfM/X0wEy64FXc3JNz/eamvTuI/bYhUvhrWRfdg/zCM+4tJvnHBmXWhbhp/CqYJZV+N/zwqfpJ
XJahSzOvO4Ea2atqNDQjIWHB3IEcC23dL5eTp7TBso0QhRmwqI/XqlPg/Kl0w1Lkzwz8Vm96dBn0
ETWBiDcGJlZp2j467bVxGYgLiIoUc5G/KV++ivjq0+peRizVpFo1ruRQas/CZAp+Ynb3D/hlO80Q
VOzIYLdpawQfIoQ19zf/mLujdN+Hv3PdeLGugHDVQstJo5tG1WWFkK1dBBZipinujR/i2Q4IQSvl
TmX2cmEb4gH+BGSQXt/EyUjYQAUq+u0tgflLWCY8hejNdnF5etpEingL7FcWm8X/iHFgjlVv1hEC
fR7v1yGrQYJCESuE6v8xCMrATfiVOt1eloxA8pxikngvD+gNw1zgti2XeC6rjHE7kZm+NlH3IGu9
fbAs7mp9E3d7mBP49rMJnx7yyMTTVdlINfqusOIGSt8FEcWwT1fOfsR5O2DOwM+efFhcoF53/EKz
7Fqzm/GbZgDe1QCH8ZsRf2G/RLoPZINQU/uRthQOOyFOBhJJlvkPTvcWhqkDA+smUYmr+yOldZsm
TubvwHl/A+U+Vn2AMVBwPugdI+I4dOgA0cjArccDwWIhPgnuLHH0Pu7BCSYab0kZ/8ilHcQ3qyfj
UUB3joF5yCWdky2Apl60annP62SbtqZSAIpN3iNECTHhLZpTGCIIk6MkOEgf9qq08ffVOyhbjuST
nT/UCvZ+alLtFW28HZNDs20+qcyr1PzkiClESsgfyvNNfxDIFlIgS+so6DZslkGQARYkyKZvX+hX
pYi/iYIsesRUXk4T8n2TZA3Uia2EyvEtAlC25L+919CTltS09f3z1ImudxIAlVk5c/gL1ntyf7f+
EsghgAEPxNOHSgSw0lKniGvyiwrfejp2/EKdl4+Sioi2+TEPJRBz382bFPnEhzd6qSRcldvHeQJT
rhmNxEiPd3nCDZJqjXZfhoMRkTfV6ZF/PSxgY58cLLaQpeDzbYDx7WaujtgWJTdbPRMKbWNkq1+k
dH3ZFemcAEqJiMk29YLkncvBrTv/Zw3zWKpDwB7/zvkG2qLeMp882OzbL5Nh8S1i5ZL/0Wz+7nwh
5fjUYK9rPE5rSETZ9VPrwp5oHEIkTaeOh6x6XFRBnhvRU5HUQAERymmQrC0ZYy2R4B8WPoyyRcx/
HvygxXpYKY9LaEfd5r+igprPnVLvtDYLKsDeS3uRMU7jNvM/0Z0XzgR+Xik5DYBhG3Uz/QxuU4h4
HbtbWDpPT7lNOB7CBFDEsAa1j8Aw8sgr8rC8UPB3nJ+DIgie7fFSviPmt7G2hZw3mPU4rM+4zapp
Gj10hqncdgrZXh8LVW8walbDJObf2F6puAPmX3nB3iXbS6bphCuvrn9w4JekBJzBZ9grsUO+F4Nc
AjDxHRA86kH1Re3ZlgmYUKly/g/+BMskdqxb1hYafwd5DwKbnRdTGTBwzjkmJv+yM5OdXjMY7pmM
FnPWA33LMHhYMIgfkn2fG1jescip5nM23K8Ig2e4hrVSu34fOG7uL7hLmDmYawFu/mG06fc5lGSP
Z8RaJpR9uzhj54HvHCOcT/zbmwwwkQtIvMAKsKq5UtabNbcB+QOdw7jfx8J8yXEy1fEq35ihymua
QExiVrrCcReRzB11kVuJZ2EnMEGzea304wItv0PNeolS4yc+m8276GJUNvZiFGpb01EcmAU9zvbe
WdjhVeiPypvJlf40QqZZ9uWAijMnmQmoLjPrFWCG+aE1vXZY++27WfGH9VPw+uvlSRNoUvR6gvtS
3O/p79jy38+4FcEdrPtutbYw3ldo1926b5qCZ1WHsS7CSezPZG69NNIdtcVKsKSq+NRGlZZWkUoQ
jlQSDfkEcdi0fcxh2xEdBExTf9hR7JhiIggVbIvGF0V+YhlQEvoVpBXXf+H1FGtmcm/ReWoQR3hs
pSB2SztB8G1pmkEZNIrI7nhXYScfkZXPtvejaMT1eB1mrCBTvvZGuli2qph1y/4nakiupzwjxR4E
WNvmstp0C8h+2QqEN2kBnJyl27QrxbYIwEltEzb87g7/COSPvM2rIjacxrCxcFfR+ACY4os14lsc
pwQ1XEYccb/274mcdMAd1gJypS4KDU/PRN3im5Z+o1W9JP6VfwOyXifGoWMV/3dG9Y6wzJmeRK69
X6T/w81xt3HW/iztE7CTFWwTV3nNA2yTLfG+EuxoO2ci7gWBm1XmZsNso96B9lfnofpMdZ8RZIKb
6QVA44F4USGJ6gy+6oPIB09QvRDRep2KRlNShnANrfJ8WrGFqn6r/I1sVgV5tBYJM2HeJQYGsUZv
lM8V5Jfc6vLPQoSeB9hOeS9veVi2r+HlL4jvTwhtGo8H8+wRB/r6yeJox9dve6I2ncT0SZabFtr6
OnbDeS/7f35y8pdbo/pF/hi1geNZPDVi4BTq0xZ2sQo4nbubjvzniI2woYVkr6lxzJDJEx6NYu9I
qqD30mrRsldzdI0ElxCWtWKHtCpsVrFm+SD7kDUEMn72Yw1YzsK5C7027f6KickfsWJoGaKwjBrS
B7eqJUuVEo8a4lwoeCYXDPAJAvW6dONHe+eYfcL/tlVYTl2XPPKAEJsiSbbCk+dM3OqSNe74DE3i
p412Jpg8KJwQ0i3RLIg7k44vRO4T63YCoS9a5CUhtFOx25RaEAQmfL87dMCe2OsW7Jef1oQ9th1S
CaRIH2KLDEUrZaJmBDlcKMnoky50DYYgCRoAfPQ2/583W02ITAEhsZ5spkfc1fxl1H46bdJgU0NN
ZFx1B8eQiT8PQmw3vdlJjxPne+KqaZc8vmMIFA+pENeDMJpZPIGB//rdh9STE78/eL+Gp9PT5+bE
pRXAYGz4ORSGAMrST2uSpZrALQLgSldDGQKWklHAUxQLAqzzTSMObzLPBNW9ft25PnRyMgWINcj1
Dvtgb0pcOCJwbVebO0iZFApNTWoFu5sTeXylqwKQOU7LOXe3wpQIleABsP4Ow6o2C8CNDWRfYflS
AFEeAEA3mSwdxtHH4REfXoydzDs/gV8H15WwOA9uv0PWiOlVFqooOl24w3rvjnQzG93sxaJem4mn
vB/kv8Q2QnlKKSbRaGvSFbsZWUgB6IDVnyXltQj5oWMdEIo5Cqlxd+NK9zuFpCwe6fBMGr6agI6p
Z4WuQtksG0zyrrz+9DaZGsvisakVxcnKlrEDA6fpfWB/D4eKu++CcAx69FMRrx1LSHfkFvYwGA/8
J+hFEWHj+aMSDKINY3LUgkodg7FLoYLZs2/zW6iD9hXIs7KXqPZmtwFvmK7jSiddYyGLzqeRs76y
s/7mVqgC6lHIfYtmq2CfsIXBk2BDRzKtSNmeEYfUbpLIBeovQ6vwo1ZsKrySYtUt4Gz/dph3pRWr
3gx6R5tp9PhV5FifTp1XReI1ZmI9nrIR6zd6J/69YRKkK41cqhxr9YmstScmPSNskEhi4njkDwFZ
SMICcQ8uQc9Y+QwoqXLSfXH7nWonEkfno2vTeKcy73zYv8NgZLgatqeQVAuIWf3aIg2TVx7HHtyW
1Q34YnK0HXiFn7Pvy8+AapTwzFrfaMu6hskn1bxjMeddhVcZxCerFUEvBfZp49DrlVVKgOI+vS7A
CqO3M+mnixs6Eb4swN8UE8X2XemAPEQ7LEBuK7ZomWKn5o8k+0pr2TQ3EjTcn7hNUjQ8Lum2Yc9o
kdQlqvK/j9AiQwEvj0ZQDFB0x46HzWVHq4l3tybOCIoEVHAwy9b4aCavlPJtCyImd3ufZjZU/E+b
P1k7UoHP9RtNgvwqiwL5Ok99GXUosLzE0ir9y6ZLnLWZFqUTuGdswIk77U+RTbik9In6wTiTVZ82
9JQ6/VGqEvHB5uVSlKQoOXwk/4kTqOFnWRTa9ZaPci/P4/7MfajasZMXONaqpbiiRlhGZPe4Uf4y
e3o0FOpukuv2Aq29nHRPqbkKLoby/Lk2yq8vysoHuad3E4HUTDZ2F71jYt2vJjRw5aO+1Z3vnzSZ
BwjZzTF2kSnIcIFKMSNiZLiefk/QyB5u/+nBRjGsAJxAqsPfPk5aTxiNnAZLzNiWURFpeuXvfjjv
eN1m51TngrsKL2R0Axo9SI9I38AAKBYHtG0i7uRq5H3732oG1Ht53WzXopRqi2f27141sOM2+T5/
P6YEdz0alzsGV6bvq8lteowy2ooIXV7htTVvQCiJN9VplrPCSvUWyKw1kSC7aaxDhcxEQ+2gG5CP
LUViX1X2+YW48Dxw5xZiR6xa0xXxtKXVAEeHXsexODQ7Q0P6/ZRdKyeZqdqE9jOOXuSSyMmhYZfu
6lHe3XMATyC35NPs8GpSfvRQ/tkS5CfOpkzHgqGlq7DCjqZChnQkw5WbTPNOJrqHy5dauLqIhHlm
1iGS6YWz0zvIQCnsqCXEZtOpJZW6F8GiH5VrmYh+++jCkNK87Yxl6Y0hxOv/8z9aOxEhZyt2EiFX
BvupUreqN4Z/I2as+q+/ZXqd9m9a4+NUqDg1Titrq1Hgt70WEkl7kY0NeL7Dx467wAD/+Lbk3Zks
baqydTCFNX2Wq0BgeIJPSJaR3LBYvBrFIrSTp5TVIxAylCnvoRVo55fPEKFwRBHRjeZ//um2gWYH
CGpdbfiOmyhxamTARUiViCIEJzrdHBFooznXEo6IzZ8rMLHTggXKpwi1sySMCS/bFOYWH5FmBapy
YC+YnKoyGf8FyFVw422FlcRs020x8gM3cjF8hwmqS7Gv2fGxMMzXSds9zTvqnAsZuN5Ogf81gCbP
y0IN82aq2otsQRikunwJ2NGjrUeJcf0o6gVOzhtRj4OtzwAo/vAVOtPxdydWdhJiZ6Vze9eryaCk
rVBeJ3Hjhk5aQyEbBZay8nW+QEuXzDtq+peBGHyCyGwXJ6ANh01Sii6sy6Zj1sFFhRB74rE9hTrv
7HRrWVfIvje8ApjuXyjTc1Y1pGyfvQcfxZnlIEGbIGuMy7cZ63BMAjI4x7qRdF7UPEOUyfqTakU8
FMkLN2a6pUP9FVyzGbfRICUtVZ63migBIpFn2BnCiO4fzHIadNhK/ftsEGtF5GSmjbCffmB6sPok
4gs4mIcXAhAIcPdD5X2H4GLotPnTW+8kMKKy1CQ3baJajCWG8e/twQQAGoZJ1nLSoFVKf1Gowtrq
k9RVpcvUbVb4hKqZEDqlHAHgSs/v3jAjOn33cMVGzhVAqK7geUtDpCY2ikcefCq7mMNYVXhMubSl
suJY5iS9cjKJ8WzEMQmUJ8S0rnSuIn7+UdOkBENba3gTg5hdd4xvMJJZCdMGXsOevJDawTeUsNMp
MiYDyHlrTuwk9WFyMS7I0LoruM9jhaIkxzCallQoIec7G7zduLid2SLXftqzfjam153uR2Jo558f
tu7Rg6VbZsBQLNcnwbKPIzeoxokzDvQOmyCGNA/5AWMVRkHhOlrIEX75RyBpiz1cG0NIXicj2dma
WW1hoo7xq/tBTf0wUoufwk6q/nOIYSTaC35nNKrc4iTSxx5Ly7COHuBXKPAbGbfl8Hd555IE7kzp
rIuS2p/ukgmj/01IhFnHE8e7nO2yCXSsSvOhLulUibE79FsO3nnSVuDHghtemHMGyyMNcWf4d5ls
op7qQOuXmSmEzmf9ZlCygkl7ySMZf3F1nvwmDTzmuyPaTHa/2pQ2dG9c4g8lJNiHBp4lERlfUjxz
vSpY9vnJQ46Yn6rVa07yO1jv+D01BRDSQxDtj8hd5ViYf4VCh21OWSEzaplQHOlDjicrEPGFLiHw
Ffa83UJQnD37BuFCWzms+sI4cH7zn8MlTDBqmf1qIYzDvag+O02uvNpSYNjcMU/YPsaX4vsx/jbz
niaPTRtCxXLN/kkndb6abj8Lh/OkUfbdODP9GSzqYm5UN0oZlMIYt45P4vDOATf3Rliibx2Kh938
JpqL4eX901cJHXjLQBdfWh7n8uu4Fhkxdqbzb66EAqOxNiF4+mU6PLS0M6xKfSj91Kf1oZEwiG9X
cJ0h+f8FMw9jMnZNvRW68b7e4E3eN5+4YCuO1hJUK0n22H60GOjus4JvbnQYpQ02iBaWseFPDQym
lbEZX+8EIW98bv4Mt7v3/7TmXIV71MP/R2oAGO5D+KN1LGKQNRkPd49F7G0T4Y0rVms2FMfIFwV9
LAVlSYjOEULvo6WkKqZbG0s9Xy1hWa5tqEFMAf0xor+Nm+1wNXD7BfYukklkrCsY5Tvr94OLFM19
KOOMOtLjxgLzu0gJznP3SP5WBej5ReApMBlCQitFNtj5k11AHt/KuuGJbVN4By32oZrHx7EoAken
TWSaLjqmoZq8OeqlhLLbe67IqOLStqU4MZNglCM6tOBbnV0YievvomeXFxAWptgouJd9Kewz4uDV
vqWPGCvwzev8xejDB00nUSOFINrajofZWME1Y2C1gKaDWuLlm0mssvKB1tpYydWwmXkIDqIfJz81
/o4Jx4h75UPz9OkERlE2cLF+IRxhjKhc4mjTfdZN5T4VBSObvF96Ah4G3Zg3tqP9oBpqwc07qTOx
ZBa/ucYB1TwL4odxkyXQmJ3ek6BmS53BF5FZ6mBIwQq3C8zSn8hGtRz1s0PM4sruMmdz1W0kVVCp
g2b8Amdun2uA8euxDqwkCfrCDoDQ4vfZhdw4litKvAze4Fq6Y/d+PEitMfZ3P4DZAT3OqFjhoAJR
RpVNNQ+egZ+gLUXekO0ECKuzxUhRzYgskoFrr3IItKa+cdAoh6Z+z3gN+zCalkb6QYhafulwl8QC
n+MXZLY8Y2NP6bEDFVSTGXr0wOWCCPMzBjfQTlfPvi8jCT39qmvS/0aXbVdurlg+le4pzFZ3HmRm
zvScSVnai8kalQla+xEPLRbVTNVJeNlW8pEFYxi9Z7sidz2ZKzNu5LSrT0znM+f6ewWlXwMPKkDB
YWZS3iDEgr75F+0ZB5Dq3k/bfHfRCL1dm6b8biUoXVL3dgIiC/AbeIZWoFDFTZU3hV2ZkzHZKIi9
QOIgfwyuW2SBh5iEJvjsUeqrgaCj2+XJJH2pIM/HdUKUFg8HbAdIErhT4PtF4cEB9pO9Qb4SC2rw
A1YuFM2y0YVcbFrOySNuL5GLqLkHZuZ7V7xKAEY71Oe/tKdKrj3/8HEAzZbtd86IwEaLZReHiyf8
EZnh0Z8cKYzB4IiXnPLoBVj8jON7p/8VynkSTWaKiSII6YzRdjx69v3B1UdxvAxsi0364lV60mfa
s8NB6fKK4LuLh0mNkjkU9W9taVQIx6fIFSJobgpDutTy6/IiCWTIgpvdWZcYpeSfGB5E3FMD3nLM
WXXOZRT1g70ORYGUd6YmiZomz6913CGIaEkwtW16We7gQKHGfKSf41WGQE21uNaVqjH2e8K0KKFH
eiaBOUDMea7y281F1eYu4cFTTW3JfCoC5QerXHhDML0I/7TLspIKbDDOQ2dUX1SU62I63ye5pn+Q
AZVqTebDCWHpBQNnL6idJrNs64sqV8Rq5q7PpFq0DlHyo8mS2siZPZHYbEEZ5OI2DBWWRhvluGA+
QZEnctv9MHnv6h2RafFI2JhSlhYFCUDkhseoK+HbLI83E/iX63HV2NtlF9azfefqAbbJl+Kkz+mP
enAFs+tIYd9czEO5VeDlBZmuQUF0ME+RsuBn38IkGWpKWd/IcsOluuvsYe5Uhoy4KRG8lFvNXvAD
aG30C9xr4TGnj6MJWNg0Wa/mfdBAN6MmjxhhLlALc8qpMOqPQ+EBOOUZ6govKVrrFtpZ4sB4FOMu
YXvV4lHfAYgiavVROD1kn7+0+QsmzQCY6PB51Whj/vMDH//64u4MVgfi3zyCIvmZTVdRkTYCIs7K
NlH7R7SGvhvBGz4HsrNIv3QVveLEo5vNRsXoLr2C87MFW5kvk6fEcp/ySj2aGx1FFvih9ePfF9/r
reVDrIw0QgMCb6hoghqvMDSVG0+Z1kfz6BV58prasRONFit5b+E+/DCjpOzWMZICkZcHyGcsN/8s
Z1s2ORBn8bVL1Uy7xx+uwKF7GN3g6IyGdL01M7v0W1KbmvVJPfWJW2NdGWHDGNpvN6lcC8OXG3ZB
ce4NxHZtGq82kYOIi4LmYxuvvTiGESTEMe2nYK6vwnVWe2mU2w8dz+VJ3Ioyq+D/by5wfkJ4kmpy
hz9U13QrvJ3Pq2QfNtcPBzu1D0nT9jP4NEKkUCb0LuWc0aqvPuBlY3qHbUCDFLNgTptXe1DlUosX
qQVgFB7GPzFUckeQOOBPUBTGI0W3LQ++eYJrU9U6hXZatAjIQeLYchf0FJngNXjD2Sh4ClhgmDH8
mX2+VWI+/ZWRsLUGJzuAP7BPixb8yt6TqtMxhLcOsW4vc+PyrAHyogAZ5OyiEG/qOG1VfiZCSW0z
7NHwPD0CGNrx9cb+NBvytOC9RfMfhfOxyVd+ln8/jvF1PKl7Scz9HI+6gEiJmbBQsfNFE0BFPaaD
JdS9OQVZp2Cb+Tr+m5XuzYGlsSbdAqxrc0jhId273/sRkdm/FbanSm8p2kl3NtdUree/GhazmTbn
hy5JPBCmwuRl0c0vy+Q8zES0hZ5sw6Fn4LScopiZpBlWF3DhCwgFeuEYCEOUcOG63PzKtqlGDVrA
vLFcJ4xa4DgCASRyBcN9aAde7MuwZMKhOXOBPFEuht0VJ4plguhv/6T+K/Rr2Idw/WVQvKlZ4X7W
A39eolQ/x8PzyfgJn+/HcHt6GWKy38p5mEouemxYavx6WRtuT5PgwoEi7CzdhN9NlIrg9AHKRE8d
QxdYYHBK8AROrozVahg4bn+toct6HZ4p4KQZ/hELcVxRPXrqNxp+0a5ys4q037Ug7ziP2+W6u5qK
duSNTgfcIvQ3yC6scefVtQBye1/Gqc2vQjo50KyAxnivJJmoAn3WTyzEZ7heQYV+qK9kKTk7DjA2
udywPmqfnU4T6KxK41xwFF0G+/T7q7Z9xluSnmyVV1ehQUiFPrDD3gQuvvskYF+Kwyhl01UiArEK
CmXK1RS6YFD2FHMqYvobrYxXDIFu8vnV5c3s3XXKlq12I1j2SN0pcpcNRmlF4NcrMZ0hMdqm8042
kobc/ruIarFWhEl8IG5gIJKqipE73Q4caQ1IMyi5vH7J2397DO2WSZouU/EcBTZjlOS5DL9iKaEC
888+A6iF4PKI0BUUCJfDB0WP+gxYBHcNoPtXIGSorJy+9/jma99M2e5o0olrIwea2lnQ7DBuI4lq
TF1dglZd84yIQGJdp2pVT+f1yJq+nAhV2itOuX2oZdrktVAr4uiOT20tRRZk+cWFPFRlkCGkEl12
40PQjgKfYNdBWLcoC5QT5Dcwepcug5I6XmVDUdaAaKMTDLlB3mFzBzQ7fHDKwe7vGhj84YLal66P
MloXLdyLKEiVw/GS6YNzVM+wIGjGJ3kJpIsmEqiHjnA4pmy6Be1EcoC+VDloZLFYhzYd0tSmSBvw
teFj9OKSHWzZL2AP4IpeormvXKa/OnuvYYaGGXjhATy7iF5wRUgXxtuX3ZbYCDpn1pRraA4PFw38
FpM3KFAz+QKuMxZCU3i3T1qZOzBXQvH2pdd2aCxqVrzlAbrcTvGq1nC5ttcIuean6dtGEf0T1XeL
k5g3q0+ESrOSsqkslbKzt0ItiL9ZgSwc0wTX/QVdumFJAq6nIn7FctvcqcH1d2lfxTT3cv5QDUmT
/huR7iKfpRL89mvZTrH1x2Rw0ls75KejlxtJ1HK08M8HMJRkxbkoFPQHUrxwXIBrCcfhseY7LZ/6
6YEc26AeTFnNoAWl+kMmmVqv+3mBl6xrs+LyLU1sMKMqc795xBgs2IJj9LHHfKRhWQFtesEGXAiN
16CxA0PwiTpV1WjPEEax4BLoU695eGd2G8sw2NQ2GUu4LlYlMbhsJ7nC2xIgGJ+2LfigdSQpW2af
fdrOKEsQGabKExY69sBeOLOo6s3mRBfYtzTcfYQXOgNzxbdYVAI2KJpDwhi9sx0QF5+LmHbzsRvB
ULadoFvEZyfsmlmZZ2GMAjz+EGgOonumus+sLSOklH72YWs1iUtnMSIz4s03kSgEpFZtWVgX8/up
VLI9USgKqHGCvETX2cV+xP9bIyS2xLEXhJMQjk8HYKFlCpNrXbbsim5ZRnoaaCNufcvEClqPaBHG
xbUH83lq/42duZgxNfy4i04+Cgs9MQWKXdOy7N9rSAaTk9r3Xaxm3PvNZPOjYVx2DC/It75p6sLZ
c8ptQeeTsG+sFSzlap4jv9av3iJDWCVqmfG13fM9H84eND1jRj6tqwekTuiVjnqhLHbAxX6GYEUB
QRPAJU3zWStSIBX+yz8EjheI1ImYGrSPbhe4jlqyocAbuJ/gAcKcqwK++aJgs5oNZjEUZ2OFvu2c
skvrx8s3rXOANQH6y8rzQ9fTn9imn0nAdL94Jks4G1KRiJs+vk71IgTYQj9V3O4ASezISfuzDtcq
vSk8KdwHjXwzC5gSUQtCCsQLCX/ZCw88f9d8VulAjwaulG9e80RiN0oypJhw74rXSQZMpxiGDQGQ
BDq2zZeMHJPKwIZNTCem5pa89gXEq+3VXDT3zKXzm2HR0KZ1jVp7nnoe+v8Xrkv+r0RaRo7/Z9Md
In/cc4JaU3FfdNdDbuUFpS4nSMSRVfu1jIqNo1p0CRiwmoyNUJ9+UbFXqDJphAEqYSu/Lar/tVZ8
eQ1gQ+aASddlTywGA4NYA/0EAJ31Qf9n/tiCz8PreWFHQirCtd04u38jog34+GG/nhRHiZLvzheX
bYvNmvwIXPL29Z1jILhLnxVh8b75UTKxoQbpU5RukCuhexJlPmPSu+t+EiGP/onomiPzIAwfu3q7
gSXssivhRaj+6XCbHk9tODxkHwsGtIkv3GsC68nTsxGqXIHEQfuWs/d/OZ/J6D4C2EIKr3VO8voy
ODmN6bDJtqX4zgMti0HpjEE8bknTBYRjRUBGcIHneoW1Ug3grryoqwnhSj2d/WW2lmBZAfdj5CGu
lXq6oe+Ax+BmHF8RdRZDiOCKHK6+DgktLBNGNxOW3CbgeV1fRzubnIw+Dv9W77sbhbwPscpWeKkl
fowq0DBwpQHmwN7GCy+3kQmqmuRt0b/FUHQqcLMPS21fNbc6DlYBwhh2Jv01a0xodE4FlZi5AXuZ
yHbvfrV/X6wHdjsqKRWw0gtTWJZyASz0IJIuRx3Qa+aV/j4Rl/xo2nwsZYSQ++/wkN2oO+SK93ua
sVdlt03pW2pW9Tz7rbiP8aJdZAK0NFxuEXJJUcsI7ZDZrBPlHf66KlerZ0ycQseVhI1FXK0u8XQX
VygCgxqcxnwq6+i2xajBh7G0MsxHg5MK/65QqDTOT4GagRzqnTJf6KOJ8ahjVWjsSnC9Yw9TVQ+/
LfuEO8W+t2Nx3UHnIjtbV3OLSCMzpxzIMGk5yofrJRp5u+6bulgpdTWbA80QFLiNW/g5x3V0Xh+0
zwZA54OhStNvU380kfMUw+sqF5fPzenSpYuQI9u8D8irD8RpArQXXwHym3EuGzGzkika9dLYZexj
nTjyR20KsYU7ctm2niBLV5g6+CTEP8g3ZLdpNIfyiKHp2qP9XzD4P8WXNS1zQp9ciUcSZG3pf965
cnrPboI423+RsazumVlgMrkbhm7d0wHWYj7CvuwFW2UIpU7x20K3N1HFHp7uJ6BytO90nvEYxZf2
1AkMCFURcIi3NwgE8FbHxTIi2A0XzvuEiGK3/B8wrlShNVrgXIOdzwH1Y6ph64uamMGycI5X9fXA
1KjR6zK2cclTAOye7CemCaRpkags5QU9QNcqIjEWrZnZIBpiRjUBI5490i6MSA23OD9HLed9RJ/U
63HE6EYr6tUQ3HUAzX5xKW8Ph/IaZlmfVHQTXmVzaPLnhunWIyHzluOTKNAXMAuyAcK2kvZJ0KcH
OzY8lBzDO3p1jK0feeJ4swt2DXD6Bg65RaXoqfbOmcWSIjG8e3DL4tEIzJyXeSJY9sYpJEYmzBfK
SxsZEK+FZ+8cy6tc7M1CgvNL+8RdWCr4X0pkQW32M8kEWDC9Kvc7ANMMXGPFaVURTJPv+Z/Ryilk
emLj8P0FQo30zqSm5NRnCZr5+oNGvSYf+KicrrIobhiP6Znhvu+NmcmHLs857ivUaGi1c0qAkjU6
V7adWv8DjoyHetvCpwPFTAKTqjur68FpH8SQZqXDQD6oAIfcACQXIgdm7ST6FNCjn4Cqfqre9XMl
+WlKbtegIahZqtPK9j7dlph8R/Hm2x/dLXhUKLYw0gxm6xdV22w8VU8ob/mbe+xx078HoaoNwz4S
HZYTpk9xbzQJsE5Z4uMJk53l81/koZekH3uOL37Ya7cVH9fs2PPZinVAwlU9qbIGJEk+/pZkZezr
bbgYxdAZAoP7KjsxrtKhtpRR5tl/1SUjCZa8QGGcqm2eskwxKMRcbMPh0h2FTijc5nFHhE84A9k2
i5dGpeMyqcCGBp+WmGowQ1v+HVPQnPBP+b1LO387Mugz3ZjzdehCMREB8Tn6k67s2twX/BYUO7wL
mygUn6FI/xgdd/LX1qDXS+mWLGY0OtQe6E+gh0E6awViMKjXyv00bjS2CIE9q5xomqJ5TE+C+eiW
b5aiY+BEl8vzyuKkgbMZqioxgYxuYfhohZK4uNozpg2U2QnVbJtlDkz/DedfRPO6vjZpuDbHxjT5
hvHrfSo5uG0/kOWhUpLQuy52PYNVLO+5kmQXlKCmzMEBLFPsrqjMd7rJTYf2bY8Ox6iWzm98BDld
VFjpU+OtFEEjA0B0VW9FYh59P80Sf3QCSiNqqrrJhn7NB7irg/sE+MO8MyGvKr01pGa2FpnywxFb
hWEvX5c4Tgc9iyqjR7RI4cLTsKpsyEZXBUs9Qc0Gi4YByC30fmgW6MiUt6nY774W++SbjszsHfxq
Iwb6mvWw35p4g7U0g3H2rc/mF8tzgms6ds2HexEVbauXBP6f29wdUbkEuaMYHFJ08qh9hTWTp0pd
mlwicNocUMD31iEPGsMulEHlr+HT01UVZMBK4aYvm8aoMuBeiQ0wPMAwVWxKKmClIpvaHRitCQmN
Al5eLiwh3O+fnE9O70fXiKvaXPMYtxkG5aw6IXirGqn5s9kLSLuXg1azB8rXMn1ANCGYydSsjMJW
CEy4spLXet4dZN1+4W3NrUu/VNx6g9MMAtQ7op6w9aAck5MmtevZofNdQaH/1V/FMnStDPsqUxS/
Z8UA1c6r4u5nQ3rxLTJVlKmHBMTJYMzPBZsqk8uOtyy4GZyvD3IIpqjE9j7b5RB2u7pOkzt4D7+I
FAuKjp0u/BRHNzeUfF0IR5O6yoFX/7zbMIGzaMDN63+weT1gaLuFQ8+PSqW+8e1fLmupkFVDfCOB
XRiumrbBK2asfVOqGzbfjzwf6/PKv8NvAjIgArQT69hxSjzA3diSg8vRxnPWdgoM4d5ld2E1fnLS
MgGZq/jDx61OZ4v+vt+oqrSrsHYDcikUzeQIVkp88QeI3umUT4kUr7hpvKAyfH8bpSxjD95Cocg3
eIvBNmioLAZq5Ikc20zvDHl04qjB2iW6sjEMwp7pvMqMlC42N6W1iPY4tIJ9MfUxE+uois6k+/wW
5ePceUrpTJgkWlafJv5BrPqYTtw7xRo6rzUEM0kn7UpPmTAWoqd+ssC/PR9USnHiH268nzQUb53c
uDig32AfsHLN6zV1tsleVGptDGP5iWfA5Nzk3+v6AdP1bqFHplPqas/pUM8rDlkbq5yKB1VHb+4c
T5HipNF2pQpjdZv1jGv2pdQTocOXJfeBFBq2wCc+abJXHxlwDHVJCPtzgwgqHpiQH/xEQsqgIvq/
jvUR6embJ1S3o5MIM+eciZA6rAwTanvZOM2myTIfwNWP1Z9pFXMdox9RIB8wqkQslwXJ6y8eI/fi
70KSIzB0DseQxpifICBR3FwC7H+ZU3FvCSsBqcmxxyE5CDL1zbn3N5FCPXYYIrBo+Rgo4vMAVEAO
w506UhX5G4OrCsFC9IE3B9sA3RtQmZ1hDPlOR6GT/veHLrukRpnbo9bpwh4KFysWfGfkpdY7h1Oi
xzW0ImslDkLnGyfeyJzg7b7UmabNFeYpV3q3se3EIoivbIizFcC62/c8RHk6FH4Zvq9Uh1x8y/AL
Qpw4+cGyXVd4xlB1YBzjQ8NUYu5tEUTxHWk2H8MW0D+LlJ+7g1S6y6xsQU/C2X+OEV3QFQjs4tQY
yEhqABWt5rBJ0MJ8Rk9DKzAJOKqHpCzPFk37S+jUmBxXMtx5uae68Io4zh7OmRbNx2nnpc1NjC3b
WEiJiaQeeO499ec0Cxnvv4Vju3ULNnGnTg/bPyG7DF46vfNVbD9w3xLJsWEE+N/74hkDDPP4eriU
KLsn6Gp1Z/mxOxsO6gjudlfkJQX1hSErr7U6jGxgoCr3rxp1m6dEi7Obki6N72YHqtPuEi+/xqpV
bY4SQ6zQic+2YUVbFfEXHaGaLb8cUWbqhMz6++qN4hu8LVnUCUUym8gd/5tz27mNvBn02kPhS2ui
WehH1JFV0Le6ntt3OwlrFdeEmczxWu8jKbvQmNJe0MKQBACUXqWZJ4sLMuY0TNU324GJLh8NsWm8
HMI1+hBONiI0KJ9wrzX17fD/Bjw7fVHwMCnUuyCz1UM59Ny6SFtsMTz9n0dj7fErVVUMFJItl4Cr
M1ME6oh0CQrwut4bZNO0oRELFkXG4cPuKuEUdSwSdEW1OKmqcqjoRc4Usl/4E9cQitPXDUUE6DPq
vsR2NQ9/ENJaY+wVRSb6M0w46qiLWj9Y43F3HCQkWnrMZHwnuAJinzWylkbUf14/6UXSot9huIRF
l8MW76nbwDF2fpliB6NP9DFuWQGj0hed996SWAFeIYjqN8EfRuLpYn9p0obldsT5obZecVzN+ML0
egJ4OBbQxoVDC2oT+zTsEG3H4nLh/0njOmUWk74SU4OPAjZVaLtjM7dz3pp698gfYAJ39UZxtVFL
dfIlhJDXGhLrTMQHNsb/0VMxLiZBSuhvYkZrUZ/r8qaj0vw/C6ZgFcbZ06W55SR4L6iRYpvGuDF+
0FyPdxQlPPNz+/ETBdoB+cakBrT6p0hrr+/EroPSFf1lgM2ca7XWYaZ6FRDn/12EdMQT9ozuny2d
4xqPT7NysMufueJderaF09DBBfQkP4weKVmItefuNvXYyCZTGjp8uL98KMXSUCqM9boAu8eyjf51
RZ5ZA2utzXk01c7+1gKmEHjnEvPVISkzKNhaunrQkqUawUHyaaKvdK5bqokgzwj8YJvW69DMJSWz
3d16jS0cuzbg3YydhySEPOuQqJf619czoxh4pIS4qPN+JwYuuWBt6xZZCPkqVygUupeIL3FMad8Y
36ekqoSqswOD7//4H4Eye/2Zxcrc2kyb9SjAdMVFWx6ND5eMQ0gsxH8r25UBrTViDo1cwXdzDMQv
x/ZCngq4EbsiCiq7SqL8pfrE3OoH9sCoIAHEQYsyEirtmUCHijjZKgbMDagBuaJ0RXBb8OvxriYz
FEJhDjzjj8hbI5JxDDX9Gco49gtkhMwvd8N8gQQxcXCjKCM1wVXgqWFopJ9uyWZJWk1DxBRTAuJb
hHADIa+Wog019F5L6PZe5bOO9P9/IfOW+4v+EtOHIgiFP32IHf64aJkYDemTPdpjtpOHWuH4UkIk
6N97FL6jy+rCcI+y1EFmV7RrHWnkVZKxnae68OGaYBnFcSD+MW2mx2ClVrBiyjnLx7UVpX9tIo1l
wCoc6lOP1zbpzljwC7HikcKVL8OmZeE4EabEJbaDuCCtxObYy3xAI1oEiFCrMoOCMZeIMufh5UWi
YD51Bws9Cep21528DEhSm1i7LhPa7jT2ZP0ySEtwPxIC+StLb1dGoDUJkRNfytOkfXVffUnPIHPl
YVFcxZ50Fa1V0/bFwhau0rKudPApIMrCUvyUsEmAaHHcqfkRzbpdEmSh1oKKQCrXSMyTV6NzXWYC
3LNZI/2XNWP7DXOeLxnpxslzw2wdfUC7xvEjW13hKQUQRHA9Esa6A69mqeeI5zkeLdilJ+ejoIG6
8fse38xqbRlRqwJ6YM4ls5IcK9ipo3KDhk3ETrEjXosuZsiT+ev+k54NsPIB7zpLAgmyHNAL9hug
CTPNcKMqLjGb9ML0fJwo1DgHv2yqUQrDYCB1QUEae2v1z78AlQ8yOiCBXn5HelX6h5J4dopkZjfV
qeiJWxDFuEC3lFtlelM2YXg0i1N7K9ecHhB/CNXuhU2uDbfwhUBXejqh0q3eogOS1+qRGRXrs/KK
FpRcPMorx/Ts44TsHWfXEHiG3i/bN1AsvcRK6kcxrXqo8XrBk3uC/wj6eKxRnGTtc1Bo/54BCWVM
2f3wvmJTUlawfY/fXOzs/JEoztEJ46VreEbYMUprolD9tdEUhxlTMm9CPq4GqN4mQQHw+uFr4lJ+
z28UxcU+OFyiKnR9bsjFngLh9oNDOd7fOX7OoLerP1Z7zuDVrHAJiRnrSg3+dVkJfI1TUMVVPh5U
kKVVwFKajd/Q4Vd70tchlbyMcL4vINM81Z3A45og2S2KlEkuFOMsm6I4VEWCZKzp1+iLl/71aPh8
9VGXuNTOhkYUQNaWhfB7w7xRR/48kd9LIYWyZYXjrHbVH03jXngY3yguO2wYHOtESLIIeUQa0/u1
zfguy2Q8z3nCt3OsquK+YtTu+tZyARUwWfame37/0sVgKB+hvOSwHMhaFFdAy07uDxi3i6B0oyx/
I1jUlRgyE7zMzuMQ2rJ9Gtf9OKY7bhF40in8Pma+R/VCykSetfZ4cxp06nsA32KXzu0RMIDNeDna
+zm/ecXx0Rbd7A7uKDy4rHwaXodokM6B2bls0bw7RIxcw6SqPA4mc97yVmV13oVUOkEAm78p/jSG
KcHuA5lkMRgysh2zluY9KjrJGRMTc2B+PnMXDD+TxXzljtIAE8v4lTmQ9LH3KulGj5yi7uQLqXyD
XV9SPrkQN6tGeTqukmw12L72T7YOT+/zp5gCYI3pLqaAs/ubPD43j6A1RbV0wgbi1PyUoGPXS85g
3yM/xWtaxPk8mknA9Igua2F/FmapCOwkgFDFKaEwjvlK6muiVwTkL/QQ+9apfqTQ/4c6g/t42kPK
4OnOinpq5W4h2IGHpSeqgnNk5K5G/SlcHlqV41HJOUgKQ4xIc30oxOYPW21CiYgC1T4Z9r6ldHQ8
3SrpP/pIchFIckKM3rKj+dZMZ+tdg7eYhEBs7u86F5XPyEZ19yEPXR4QpCGFfOPavtMF+SecfzyN
EzCK2eQBMdhJHuf5IIK2G4+8rC35NbC5cg9dU9uYHjXauqcqk6WdMpdFNAFCdqewpnJ8WmgrCgZ2
TZafLu4zloGuUQrAEzUvW1zmtGWJrfFj8J4UpwFHiWZy903eQcWu+aaCspw30C7XTf77f+GROa4s
WPepVLCULSzxbbcWyjdELhM0psauDoQoTN8qiGa4soGfANSGJVSRwyTSCjZW+f/GbWucH8H+Qw1x
nt8ZkEZ/NjhMKhbhBnX7rSn0hXUXpg+KgN/i96saEnc34GPRKdFXv5QId9PeqJg3rBzGVzrlrwAI
gPH/TRIePJx4ebiIPGK36MivXgXufHM+gSv1b0cM4Y3CtjrNnjgE06w4qaaqh4DrSjyubIKVjC+P
ptlji3FpSstxk0PMGOxmgisLjhviCnMPiZE1N3KIcJEY3F54hUAnDFyGbLmTCn7HkSaKcFI81ycz
uoWAR8sUOFwmSaM0JQuWT7XX9S9b2PorKdA3NSA//lJHQ3nMYLaUerWPBDtZ3TV1f1r6/jvF6Wz5
YzW74MepaCV6lqFmTMi3+mgBqoBFyLHbm+/yiAiXpDGP8mMSw1tZVKBmP8aHBtZ+xQqc9EkuHIU9
pYraFiOz1vgGr02As9JRnk7nQj0tqjngZXBj5bPhE8+yD1ZshQWZmDsBDj4r86fKQPNoNoX2Qkks
JJOko5NNru2qjIPfWJ+uBqbyjHBb13U2N+kh2hFgbQmA97wujj4byfhnBCbOI5Fk4CyHpJORGjGZ
tkyG0zO/j0lJLQdWKfIMkpXDjDvaQXBhhXqxFX/hm1ffZRskStV434+GL3ySQipZZGI7I7y0n46v
8ltTirw8jIsqcK6/jOxt3wlX05/EQ7MeSDcQhU4s3C5cXrbkemmbdgDsbs9IFAX7DAeul/afxeRX
kRlW63d5zO6CURqfb2ZYmwjCXsxbj5hofl4SJ5lZNE92V68kZccsESW6t4QE2HmH9Q5dtOmCuQv5
rd2E6OaN5XTAG4rqdjqNLQJnfebIDaQYPH5L7PpnrVoCUaq2YhHlt1t9vPz0BtL+QzFj9i+s0mjD
/B0+Q3BoQgkD3+Q/iYRznqNiwDuJmNUMOegsxFtXW1+mu82nfZeBV1zwuLcn59T9Y1Q+tnK7swMo
d/6QY4dNtzC6n1hAKMUgGBUEHjcpXpWxDKwifULNvzGHOvHYo9QEF8ac56c37oirjt0kYc3Ia3nQ
avga6uh2v/hSsOPjbskI5767ztYIwM9hi5JR7d+b92kPEf5xOBzuH+ZXlhY+YSuLHJBY+9D9PyNc
Wl/aX8twB3C5iXlP5Q/TJ0RPj3WdrnTVoSEqLkHkHL8bnABSABaK7bijkhkLEeAAUSKzgqKCDqgS
cijfMK4xj42K1I6+SJWKwNYubZfwEoSfr8ZFrdasmZ+GGe/u7GXvHPu8cG6zn6dvvBJmJ5DKOJM8
Err0KbQc1tYpyc8O5BX3AeoAcviFbC03hPwFnOsQAfKRVzIjwwTopgjTxx0GrnrnDTMuF5ALyEaz
qhyDQYYcAqDzzDMTmbpztjpUNffgRCHj3pUd9NzqWuH4ZEbdDAS/e7g7Xcp3dFVGtYj0ohu+P/5n
G+0dXzvzAOM8+2i7tU0siOOkyxyrMNfBCZbELNPbiG3zsPNCJ+bRlEHG8EJ0rcAF4I9txLpt6DmN
UlBe8JuxgX5QK5DHRssF/MRO2oeHAoVOce0+FkjkXDtzvtQzw+QwUc6X3aNGNbzu5Ael1hX+Rnai
h3gSwj9+RoT8ut91CeZGPyuxlLkOBJahGLGI6JCdb5MtW5HsW1uyX+KPwLEx1e6uaX8/TFFzd7q9
UgIZXVdNByQZBR0hyuOtmE3FjmHhEt9JJZ57YgzNX77wxg8THtYkaGovPIa59M6jK7Hojvb9KEPD
2EwsO/IZduYVACw8s5Ug/NH7anQZxR01EFn7MXPfCIYFkcETwqdHPjDcaSd3JGZ5DREwJnxD7xVV
m1QsmQlAZ5k6f9walOEARZgZhQqyZ2dTUueiSr+bgYZsyjpPVuPNSmd0FYJUjHksfNRXY9l+9gIa
yfQdo9OHOqDyZq+njBF1Zovwlbs4e4Vccz0DjAHkLM2NxuYqDrIiA463MSvwrzuyziJ3baWWwJii
wFZdn+ALHRrlL1UUFJZIaSCGfwdUNgmKxmcr3B96idP1Ob9mk5PQkvFSob7OKByGGoGPMXuxTNdB
m6inzAhdvp/wCW2vke+f7alOMTaun6nmTWcNSNJRvKGUGJSTLNzUNXeOhmjjlbWSpD+xf6QTJ195
K4hBVX2EzGamskvR49pKzwccFTE10GHU7JEBEu2upG3jUDjtJZGqeTvNHWJh3lRzYZQZ+TgnNBI4
n8objHICXRTlh12LlFEzx9l6IXOF60IHlkEj2KxaRV5ptAYDlBCu4Y1m8yOCpFuYmTAOsFOMqGyQ
/bxRJD3rP+rTDQ+h8IHfNxwVXxbCW6ABFfUPw7UiKX1UyMpLRjwxZ3MrEdBDwx9aFPRSG1/CxZZD
ki4+f7x9d/grddPBvhWdhI3yJFLetWShFAjm0ADjoORnLTV/mCN4XMvVkpgGEoZBpr1fzdkvA92R
Yzwe3x5cMJ0WPfdYu4MNlDnhcl+pLh9L37QF01u0AvFDInKGpU6oUeBBNGq6+MPDEQbm4Gg8HN5t
ylm34Zc4aL1lBF0cejbYwEsXi1WTRianSD3QFSmA+1BYHpDRPyUYGa8R4eDZsHhdVu3upYXX0t1k
Gg0xXospQdx4D9VasNb7yqVJ3kRb95H2mAbUOo3kswLBZoOv3U+al9Gab7ek2gPR/ZGXPxFW+NXJ
ga1ULvcbByAMfsUUeemgNvcltASrlkdPLWzeCbbofpQTWxwZC/hxVsjjR+7R3HP0GT9lRXUZC2rU
zd/gWMUXe6Q3gS+O0JBZQIZgQDoRGod8ayaPMpQEUUQkek3AGdcbGp0y7ACJvR2sczCLgBuQoUFg
e18cMIsER9lukh+vBqbRqbqfXQALSksUt86CiCzpj51rgG93nSgq8+A+ooIOHperuJf+J2boB3tE
QO02pJ0Q4MNA/T8hIQngwi2a8cQ1HYCEU3eg8K45yHbqlCjYc0P3nXQDB/WKci5g86J/CkwRuHAQ
z/XtZsASuXHEwmBUYIWZzXqLtFvhoOfVkELs6wveB43deZ4wJOfacwPqJOrsCoS1FUAYaSWbH90E
AIUKGFW3oMeONytp29aixdIMOHYurJp5WBDWD4aLTzd6SKmRney1WQVrXbC1CvmGaOjlwYw+oSDI
GdaNYoFBdc1OnWn3H2XcF4pT5EDXA9C4yGLGwMa65BnwY/xYy7feTjG3Toz3/Js6f8JznujdOVut
B4PokCoQb0/S1dVseRJmP/ZwsIAg5eK9VsWXc24mDjaPXBDhX3OLsGZsALbH8FJ6wWGhIRLTrIoE
xLplbEU9XtvliHF5x1dLnqQqk2rWMcL7n6jjoPr1U4LxI9D5xIcVeADhSrWJfmu9A7x/j5YuKA/l
ljhUEYFpGj2xK1etH+q39AT3PAUXU1LdAeMDIdyyue069yRiAPlAAYMTrzur3gzCA0GhKbZe6sqM
h74QI75z1KYOVHFqVcFdxBtLVwJDvX8MELrCs19C5o01nIMGKgUCAkUnCkao9meNXhBAl+7jDD0/
0BNB0BuhwU7qHdpogip2Zo5nobRKbGfMjx9jvjqbHBqVxZInnG7XVO7lGWGROk7aMzjkmqK/WqWv
I2gRND5kQIIwlgnhinoWmN77HGw6/fRUxF/K+vG+K/PBLeQsYGkbd0x+nZMvrsZq19SMi28kvw5e
RecTBREnS+49yhOVPOHcz/5g5iIKikx6xPhG4ylS7w7VYyQBqTCq2qgaNDMta1LqzH4Yjweiv4xz
uB1L3uqivBOXMMeFOsJ6H65W+tFOSwWTwZhkaWpKnUXegZNRRrXpxMGpoL8vwKKFrZDjKMFPIkw+
DAd9diEwkszAEof4jaK0jSPwt533UXwfdGkceEMn3pzjDBQa3ecNQF5ahExCMorYUflFKtMx83Td
1jg7XUJqySQ7XVVnICf9f+2d5AoIVwlX4WLFpkWst80QN2wfI+ijOZoHOJVsGZDtxd3m0iwhofca
K4jv27mMxqLP15fLH9U7Sb58294+jEpdj02NWUUzuUWiwb0D3//6TRXYBxxYWhyaiJkmsgSBEujz
0m4bgU0UwT8Seqs9UHkTvk6bqJX2xqJd7lN6To+8OIkPh2cAanrxLCeaE+wtaNgyVtv8JpXHAkZ1
sjVbNBjnvyrwpSAJJxOtO5g0gvBMfa3tQButkmAjgUsBJvhPw/9mUXTyhfRxZUDlltUFRMLIn9iy
3YP9XIw3ifwgi0haYzpwXRo7Rxz8ThJpayZqOjkqZJAHK9nosnxSntiODfzr59VfJF5TcaemB4lf
zy7B2D+B7wjnK5dUHHF+lIAT2te4ULmnSzHS1+wXRt9YHXZxUAjtIpEYm8OoKQpt1xJskvjWuYFp
AZCvoGWF4iXXQdb+M7haRcu7JbYFggGLc5dvKcEg4AcQwZBMTj72NIt4aONo9jQeSkyehfPF/xQF
KrGhCFlZzXWd+zKjF+cK8GY0sJSA0VCcqjv/wv0RuQyGl+oNSQNIQtPGwkjE8gKF15s605z7NU+F
d0JUaVN4d3RfvrF615sP9gRCkNEIT56XdvJUWM4V9FPWjGKQCEEvgUyd/mWh4/fF0uEyJ27KMIyW
C2AsQlcSYVWIoWl8zaama4x0GKURPtaK2fkTArE+f1W6oWCcP+mnR9tmLy5TyhiQuNZwFV18qwj8
72AtR6ujRpCvo6MirSr+jQbkDrAVArBEXrgaWm6OX3xSyrZ874lw14XX48OTvzDfasuLMf291U5J
WAsLaMr/UR9jUw+eDLnmXcvfkJGR9wfpCMufuKFMmKfYtvH98YTZWnITbimVofVrdErPyOCG6fqL
3nwCQlBIJpPtmo3jym1qUzF6H+i5Bk5IeJGakPCBoBN1W4qFJhbj2YFr4QHVSu1pSLKVgmRLq6de
A7CRQzdr98Ko6wFqOgCZfGnJirW0HB62zzRQpNNji61nW1PZhB+u/VEEKc+0OSbZBNp61xUac0BD
xqvarfVYkLkG5oopoKFHItRHkeiQwobb7HPo0c5uxft16GrilYYREGBx9qapiMJo8GlVi6FSQxTr
ci9CgxY56XQO0I7Ecuv6ObffYwg88uVA/t8EPvnDmTTex77S28/5RjoxMkWoXcY2DPWz9qDX+XvZ
zL6F60iAwo1ZX1LJjMajnPo9ttw7RCWYio/vCLaN+Cb6B1WMQWdUo1kQsydsq27sz0yY7iqBtNdX
0ouKQCDgbMwJ5eXo6RowAgJ0l93xjRk1sblrTK7eJEOh1fhgvl6sCg4opXM/VLoQVtdRP8j/Qh2Z
JlXP6s3Tvt/8vS5fwPiX0jJaZX7xvzNblp9YfQfLIe5Iqg8KihHdyt4MSMwmGKDuLj99XTZquEk+
4ff/InAkvt6++/v1DIGkbWa7t9r2gEQFGGhv0Cgl9dcy3uroHZ8vFOTGOUldqB8vdonxouV4Msui
94HLdCuhRQ7Lq6HUy3sWUu35OqH7B6a24tzzndJIa7YIo2QxpqcPAnGw4mZwpqzZbiGJ9FLsPRqr
/dBaleuhfsMzsJx7EJFII/qdhD+YHwFasLyqc9j9DM5EH58ZEFiDA2LWy1BNp/GienRKQXgAz43f
/QO3RuvEhjjSeqwuDb6576WLb5Q4cfRd5ezJFkjz3xtjA8kjUMDLz7jaWbHqA4ecgiL8REeb5Q7u
HlngPO8zmIaNGjYYsdWcdBCB92uvjltLSJvaOcLt25wt67dIm3TCDcOTuU0ERKhnEqWeP89kQhYo
+PogDxA9sJhEqGuUOneXYg9e6vqz4NfNAnRwdhYEFBKeTTBcSgwNR2r7n/oljWAC5Io7xJ7nNCmN
UM0Xm5utdEypEFan2BeLBkLt+LqqhxLhtx/gEnMx5HLDbTQL6JdehTayjVSU6Jzyv0PTXY3BxkR1
mF9HYsl9mEKRqzWfz5veLe3Nx+DBcztypexKyYVWYixaeupbnjXsJnjXMtcdYdEOB5KONGok3ltM
GPWloVwT05kMr/zlV7RTiYjruHpXjBp2AEV1NQZUh5T27GH2Af7JoAKNkprOadmkqWwqlu4/mIq4
xenOeDXdrH0pn7/TuvKyg9vFMYUdPAM6MffEiJ5YEoStgr1L/lyOM/gh+K/b9lgRxkVkyPXlEBpF
i8dUHpLqSPXkb9npTe3cQ7jwF1lWyIwR0Pd8fRJxctfWFueXjDFVdAgjOfeoQgYzuW2hO1XdN3TU
doOSPF3s3MGtK73YQzRiiKF/Nm2i2p50Bq4Wcq9ZeC/P8v9jX8tTDbph/HIEBu4XZKnQLL1Rspj6
BCasX/x6XLrMpUKVvyE7/Id32yKucIYwjIAjOp+oR/Mb6Vh6BLMHeK0U2/0Rj7ObiBqlNf11k868
TNQUy/lrorr5LBoIrkJGAx0M3HfembvobkMswLcG+rYS1Ni8YJJFBEbTSXdmA1CCu3LaO2e7RAOM
wFhn6780ypOkqxru4Shn+krhzxXYk5bVho5ZZ0eymeZxNBp6HB/qvHHdM1hIOr1KK80GuXcjXf9J
tdju/Ddcsus5fr8l3cSnd1NPxohloOODGHYvO+GLMcYQBLEO6Oa59OLFasioixrdUbqFsHJpubdI
v7JYAl+gDsvHoRONCFzREuw0fdZZDF1VeC3K7rV+NfwDr7sQpS3E8dYtYzrz+oXKi/9LfdN6eQ1K
COBsQ6dzSJqqGf0WkDcLxRz5KqXXWGYlx5NWraGLmmjsyT8uNoFFRlQok3m3sstquxxCcZCM0ll8
GBp3sEShCdv8qPa/x32kai1v+5wWBoDoyQDZLrm2CZY9zgQQjc31cWUjTF6OcVvYIziDQk/rwzV9
0qQ4SIYpaSF+JIRKYRd7DR162mXTcrFUhwUJXawNuuO6hyzWl6vfKjK79oYkJN5LzHYOvYn5n8NF
EnwDmClYq21/of3hXDioP+UMfbmUD9ye70i/9oYQzQ8tEadtMF4ckrbhLYvDvMnP3/tFEEqNu41Q
fEJeeVonN6leLU43qk5Aqe3H+0nIYpamKuDx/5h/qC/ppu4pIH7PDrxSPb2isEgu/ErydDqroNev
/VGGNSH2W7l7TTeyha4nMgv6S37/zwO0nOPFESSLju1mhYae8ZnHyt/9d1HQ7BJWqrFLkhXsDRLd
Agr7pGqbGTiinGVN1bybUbNCQyDEXGQcTsAygNaI+m2jmfeRcb8DGMBowN5HdxF7lQg13BeJ3R/e
Us+76PIaIoS+/oViDxa5aGqbbVv0Ax1JHblOPn6NFwbAG5ISATGKezTLeSKRTvl0F7JROV2WmDJx
xvyKTk+rNp+2cR5wTETec9qhJB+IadgK1NyqrUnjmLO9en8QCFipLptgVikeZzJA59KQfa/6cynI
S9grKlGXLq4qLeTvcKINUSN0gZxcfKxhs8SMIxcPB8vGdIHfNKQx6ZzEssMlM39ADssR5b3tVWnL
aq6aykUGfQOcf/YLL3sGfvHej/V+2RAmiV5GFj1V/u1Rsn6mJv+bC2KvGnaaezD+2OmpeOgOJfHt
0GCXynd1R7IeRegS4LHloSpAVTgu/l62e42OXMh7TCbyvsgSIDUr5I7Ow4bAeZW4TMeMgl+QnIIa
+CSZdZzC2jQjHTe3DdnsEq0RL/OlYf9P45nqIn+AH5EuMgQKfQlGE3J7I/Rf/rBjM9bJCckTeG9O
8evw55Uti0IgSYaK/3EMBuOklHMP8U4kQERx0WsbwUbgrZi2wRvzwfYlDAPW2k3s1LUNR0kKnvQ1
frJNxwDyejVFJUbR9hJY1S1DrNKHzqVPAwEWXxmqVTiOP3m7XY5SAkhA3GuU70iM1FrGZoVvpdaU
npfno3OqVpt+HwHuGlnlQm8bcJPB2GNpPJS2agX+6zbpqs/O2RZ0m9LKvnvdYySDXhJeJ/eudC9+
49OQZbVbCOEj5VRqAd60sKrmQC1sadm/TzC93DOmlIvAV16d4v1My1ZUF11V0K+kZfDGvZxRMlkR
QaiD294HJ7ijfWhiVgkrZZQIUrKZQ2PJxPgDRBX4uPoKMyBJW/E9h/NsJ/3ns7PJNamfsdatFIYZ
Iy6DjCg62nl3SiKWKRQNp2LBm2t2tEOXWDFe+h69Sv/DqCHX88e1zJz6tmmrVpuSmk1PPoHvhHty
9Lt2XLG0rzr1FF1rcELm5RDRw78BmQEJ3je/rG8lnw2ce/kbBAIdDHf+TXNe/hpq1zQ5vDnazXvb
rsglU66SH/FqI4AkihGFo+vdzbPdVDrnEHe6hYLUQ/A6yVT37h9vTlad//VyPWeSL1fqf9ZkePnN
Z/1dSDF31bbXah7ni984Vx0Cp8ye1qyNVc5rTNopj32pWTTy8IdHjSYrr/dMwQt62EUXaDADcnA7
dsgpRkUR5v11D7IHlSFDDF+o9xhzsIVRTm1g2sfjvA1IixCmDC9V4MZ7m1lv7Ii0KSIOwlH4QbT5
6OpsLIhRfeBMprihS1Nmpst0UCJUsYGr2pYD5Rd59vMQtZAkT1A3PVr6w09WgPlyLUnKXsXOvzAm
ShA390S3GV/XsCLMnAbhAi5F5wBaL7na2eZSRer8unJ/F6DKIYUHWTkBQ91aUrqKrqmfmQTNyEll
35hd/lsM5ko9jXbuDUlXAzlrDN8+vcquCvmkjdOAM4SIFSImGfh0exvKAhs9OFMA3Bbk2euZuLe4
ejcWDA7qIuT/dG67J14NI9xnYSnBLuqLVuwh7Ct1+TmtcaZHYh+6ETYGcxp+8Dk4MlYmDxihr3zt
ssQhzHqY63tfnN9aJ0eX33rCA5QvShREr0S5q1OE7x3qmhqHRcNdLEWtiDV38Rh/z4YKWbHRgTQD
bfYnIp+osTbvbaU5Ud0+Ymkmapvfx3O+T4w2ZTzL3ZcvOfmmkeEiYIKkzneV2cTTwedulhrhJsrT
J4TxGTT1vtwgMZZMgFkRPlJwMSvIw5fcy30iR8OaGFyZ+1mhKOJRwY/bNPX9IzgTRA2KVuW7t+ZR
Uin8hdR3p69gkgOX988B7cARCEDPKg6bd4XlseZfM0+89C2mrBMhb/VbsTOVbo0SSDKmX+3FCzWM
fHwu2lzSshy83PUb6QxxG3bY2AlsWWf6210L/yFSLHiKA/GG6xwveuPc0lszwYbuw3gF0P8j4Zvi
bUKbgWcwsmIKSecPryEbKPOzKFNOGM9YKCuq+LKp82UdC0zZGcmV4ndCfQwFGh0jDdXmgHelGpzR
MSoh4KjJ48juX6evIVM7GKq2Iwa/p6ny0beL1odzqQFZtL2v51xrDbV3dRNuCO28IBNn+Pvz7i+F
7pp7J1Z6qoGO06deCvWo/bdGSfwILSuXJiD4JkVOn/U1+8N77ItqmfMQGmoZqVKPK2rnQKquKrqc
d68jEwXtZmsxQwMIiAjERMgCGquXKN4CfdzaLdt56nU/wpsZp3TjCV23BQXZYfK7WgIuEsk2KjIw
pXxNt/6ygwf4tDAm3+duRtKtdJYqqzdRbpSjhuZiT70nvSyPtrpSPlZaPPPFmatEVx0k3YIkPdcV
qjEKi1vWfTm7jRZhlOgdF//hVyPEIU4lHpNO62bq5FFIhAA/XZfuP0YDXGZQbcdwImA4TLf0XVzs
y5R1Bzqf6y50hhWxLhnfuY8nBoG4r7JdoGZspIrXFJjTRK90BpwjwCZWp6mT0KE7Wbue2im7vu56
ptBiZhS9W9rIOQJrPstgRbnk11JwK3jtCzlemw0BEzZEti62lf4Y64ClYKBY1r2ecXXzKFtRAL+E
wuj4u6Q1lVPQWIz2NjMzc0vRgGzjOI1+Ji2fJ/nG6j4c8OFTbvMKY3ThVVXyuCm92VcZYlZdOgmm
61lnIBLHYI18S4kTVIkRqgCtgGD7YPU6NI/B4WxKGyFZItVQJifE2pkhSdlD2Fk2/4nFcPZf0Wr1
leFSCmYNSXVa2fDlL2yNbDifhTHHhYfsy2uddsjTwAA69XjiKz8UBKxuQw+x2eH5HtkI7Yc7FLXH
8J8ij4iDDCAE5+ppcmQ6BJls1KIZHkb+9PFLFVpaNfm/W2eYcehTxvyuj1nSgH4qx2iYQQX0TUNV
GyOOE96AsXwgLXiGYz1egsdi/quoHSYlWSAA8+biOfchBsBuOIN98ZXaDP2HRDYHeaHLZa2jV9Q4
4xxwrum6HRhnqbRND6M0CnuDqhzqUWV6KOzNmyrZ6Z6JLncaZ8urXaS3+slPKkV7xggaejMl+MWT
Kg75xzKWiAD/vRUs83LmZCpTmjgQRah/iupugu9S8j/hnEVSJBM33S+5CngBUaB0HimQHBMF0sih
rlUty7VZL4+3oaDnKzpcMLxg99UuvLAww3UVxzNEYpENokOYWLR/4pEduTq5MqyyK3tNvmIR8Q3H
5jT5TtQwpH5IFapGwonOVpezpSMz+O4/89xlzVzhQBsa9NwCFSpEr9VIjNPbMK3503EIKlXsWCLh
RZc+G6NT8JMBZmjrQSXj42udJgeNUGNsT/AAYeFGCL2Q27yEv3+uXUUQ5Hcc+7cQZioZLiUYM9ld
HAuQEok2Gf1D5lSPeJcvX27h0mW1QLiTRADC5RcbopQK1u2pxQAk8xJTTQJBh/s1Ayq+gZoQLhyb
w3V1MtMDwU48Nk356jRLx12aghx3m9r7oXOtru5nEicg0x1p8abDeuPjm8j1SpoaXp2T7Z8xn9Yd
hkadSSm/EByNDvMecP7wCU4fhF+DjDs0doWyAQjkkncNbUs6d1oJHKAZA+9aNy40k/8XhNGBerxt
A04k+LF3TPYhfm/9Z9HfNOofGIyCDg7EbJdOePWCKc8CJPj6GShDmwS9AjEI3oaWaEsIzAOEmvUu
LsDcJ1AAW1SjJL7vqSeqsiDuuTG97z08uNLKujYJ2DK1RhtZP7JxQQhzrzNeSjw9USGWFDfFPplv
35TgEWBpfX6J2wfq4OvR3ifi+V4DZEmIpxA8iZ20xhWH7axM14rKEIDQechJOPdj2RxtAJOSkKd7
of/29kdDPUcoKke7GuCCrVjh8SCgACbNkvLj5E0sORzkl5JkP8Dimm0Ri2W07VqmmWAOXH4N4m6J
Z9kOqySaLj13Si3o20GEtwgLkNO7GWidBUQFFRekvxWXY8ZX3M/WGzaW2E2oarOdqBziaHMful6O
p/AZtSGLV53bwpx/l1umMYhjd+qHSMXSp4u4obTAdTSJqdvkLIEc4ncN2QSwCJoWcI+tFOxXX3Wk
YxPk8dPMxCmrODDOjfvmSttyA3ZfIsLAejZmov8dzfUqSi2JM6Vw8L3XZh9rCoLuH3e9IAwARoNr
RDM9WeeFylmPXezqgACFYp97rKe19Vs0czrogVrhQrahxL3xhlQaebDhFXLFQcIanf3HoMdt/Umt
GWQ5tdFAbvF/gU30h3hURG92OXz4w6MM2c0Q7ahJOiPVmkk0DFKmX4Qy9kLPEfqH9bxZtwiwBQNm
r8R8cpuOgXfjxhUpW9HB1Ogg6CeFujiAWWihiPtyAoMNUC1EOjh2Y7mhNYo96chFsBOg7jFGK7e5
clURCTq7qMLm8gh9YGHpDcmarEWbX7x4ioo6eUdETUxggj60TqQ1mUZ8XorN2K9WDSlRkMcPU0GQ
IgzZAgcJsL3ahILhChjk9Pkfc28WsF1R98x3Slp/YmaZVE0lTbAq2LmGHpitBBwxRrK7N0naR6Fe
R5IvAMFPLZPBcYBt9nW1s8dkaQapn2DXkoDUPAIKUIXX0U8qZ45zfHJ/6SKZc14zBUF+Ab2z39ra
I7DymlNofstni+vjKMwKhYVTq8U8h4cG0g9mqiOtYz9giKozdVM426m4h/aXoYEkrAjsEJ0b7Hp/
MLzsAk0T2yJfUZ7X1E16xKvnWNx0pXHVzV5byv+62F3wRIfNf3Z2Kat7sfNf5cwzjbl11XyFvaWL
HW7v28d3nk+hN/L/yiy9DI2u0vbW6DgEOjerjoovaIxcJCz1dos2+W9Y2hqqWj9qSp3WlW2jqG+O
qdL63evd6+75iYIbOrCIvhD+fuux2IaZMDYB/WRvINiNopHDKO6piHjbSiNkLSpF6YK/6ge3Askv
dkIgx5m4f8bMvkewWH5wo7hRKx0fpPLpZEcJNi5yXfA///Y1E6bP5qtYuCsZHd+I1KJaCNvAHXsm
Qj3GKsQ2sI3sn8hZ4na9NPMmhOVGqLVSaOMyOiHYfm0tNfeWYQpVrUXiZIV2QY+Y38LDj35WWlHN
j+1trNFB4KRuLyqH9qyvC2R18zYdRMq6N1kvFGSc1tIUumdgNoLZLUEcgKTGV9cZ7YfTDRsDfhQT
ZlbquJzNkoyGcC+mVYyHcSFngKcOvuY58kn/Ldg+WhDoS67p95Z6OgoNK6JkHs2PGtv0LoMiq0V6
PsauGySnKRwTsc0S6MyZ0/09MxU5yUTZqN/RXJsH49fTQsss8u1tiARm133HzRWhAGVzNg/cwZkH
B2LmWOacwdxgT6BLGdiegEXJZScL5xrvEV1hklFBxEUpJdZVNApmGwcXf/CMjY3vEAUCi5CxWaWb
uFvG5DQW72Cg2S7TAFKxzzlijSIJG+44LD8PfBf9HYVF8/9G77y9G0Tkdx1HFflJneCuWUYQe7KU
fa1ClirE4JZjdWDLwzgtw+xdq/XJRsIV027+RDhJmoJf/Lu4IyONVaIKLtYcjMQIv7vRHHSW1mCn
7olNzI+BVRbaFyAzy69V7JQvh6dybFzbFFm97FUjWA/W7r+iER+/psLS2BFo32b0Kwjp33z5rhvK
CkeLq7T+1N6hM/9ePyoQbF8WqzKobHt1DLIavHITvYMsmofJSRIAxMWcrb9oXmA467EHjf33jPyL
vNNmpFbDdZDjmwuwEJfT3zxCkqqVN2snC7c6c2qUX82Qngdp8BnRFh8c2GWRZ/wuUVEEigD2wq/j
DamxWGWm3shohf4d1M9VxW/6jNMSbxQ2WgeoYtS0w2zmiZ4K8/Gu3KsTlPsmdo28aVtyOzmIb51C
VKPn8HxPjn4RODIl9BHMPAjKtqrDSR/y0Mhpk0dbbRnMbE5rry9fY6ZepRMrH6g7YJpdbHUFv5y2
uHxKvZjwiNhq2BUODExe/EWs4B7ZADS1azrQg8bGxHh7rU37cJ3Yt5ciSLdmqpJQsGtfDM4z6LAt
Q+eAInmOWyRbVEDZDi6ail2sVGY/sF4oqazkBDwf2IAVOJY5mUgAO4597E68LtFjwkOC5WcBUsJs
tdiqeZpd+0FP4v8hQ8Qr8TuHsOwd8rQTquuyh/dgB2/XHRHpp20jAwSEnvU4JvqrQ9ZyZPvKe3mI
3PXzE9b+I/DwrbHJRkABIkh6s951QNh0GE6V2v1DA4OED3uKE0u502UyevfujcfvOVYvh3UkRR6h
uSJFj7zKkOJoWJRLpHv4Vt85GXUxduONB+OnkiFE/9+/z3IV/MnnCcJH8PVEHT6mC/wj1aHudc+U
7rvFGKg/G/gfQRSVnn21zVvLWJLJ6fe9lvx9q98CxexM5NuJZCyNqhuurQ3GrzahtBUyzmj7lY4z
GNblRZSLjhF7v83h7WEP31owNgyYbXQs0FyINC7F/nKT80XvQDcfVUZyhvzdVyxqx2/8RxAhPcDY
vDtlAp3gA6Guf73yWsfaVkD46YSdFqNshK9JfMOTic9s0ZEmzfu+JuGxAhF4z7yGflLyY4K8wzEy
Vazcv1Nw23i+hf/8DHySaTmw7e3us7xqchZaXgYYIGdiYnQ+/wl07y1vsC6fMjQzVRVtGmSm5FyM
qe/RCz2Sx48ZYaWUvN+uy6GFxDZE2sltmWI1aT4Avm4JYhxl4NPiWRXQy/3+RKGCS0c3UxYTILpb
zpyz3dqbBfheC0Ooo3fB8Xn8mNiFGj+FGe0BgUD0tIG/pfO1g9to1bPQKtA4SEtDA51kfmYg+u15
JIlTZspK8iMLFbloRyngtY7txqxgtvv7z8pbTm2VUpaJggExcMR6NSUn/G7hQUhX2XdtHgqZ7znk
15+QlozRQDEWgNDJUZGSH7H7lEzGGV+4o/XXHWwkm3e2Et5jMtY5BunDe+azxLjsuUUdeTIqE0RJ
iktFNSJKaQthlmWNBMcIf1BdFcEj0+0K8zZg8AdYMEww+pENSeo8Pw9sEjgXcfIF7kjn10eBpjTx
AzRkefQpccwc5XaqVljvtuwu+laomnnI/qjUO+FQhh4QidAcqX1LpkiFM5s6Pf+5xMKDF8Si4JTm
qppOhrOHfVyh8XFURWQwgh8TOlSyogmpJJgLLJK29ZVjEeFj2ob/yHStiZdv9MS8DJI8GiMV+AvW
0bMkBpsAd7SM0ahAD7D4YjHmS8C57jM0QgHHtoHsqvCta7v50g0TJE0VIGGz3A+YoPyCLC39Dvc4
8ZnfNKTQsvCc0hKG/JeN7C1hZyBeztnhuh41E/w7AeoHKjiZqOaa/acU0BQIoPfOm8FnOusZ/Vos
xo5gzFLlmPuRIE39jVzImHLyL2eKGZVjSC4bAKEec8AxO7iZezH+UV7zSriUVJQD3deSuJro2Jn0
yI0eQfurSXi5+66MCM/O6GMaxqOCPAT0czJqNZRbwD4MWJA4ddJdBMK1LTvj+x4AXbQOgCEkoGnh
d6J1ti6TnrTvGtlP4KbJe5/uaA9dzn3GkOcRFpC1dWE4FEIQDlGgm3kos/nL83NY3h7WgQbE8hOJ
zkyMgQjNP2/N08ih480+bYUALxwlzNBNvqhBK5lDdb/yNLQmbxtl2CXTNtYHT0XjH6Z4Jk6M6lD8
4V5S1XEbc/L1Y2b5NynplzjnFlNQzI/z8lvsPEzVRMe8qSu4hrzubzmx2eQtXG12Xi9Fhcjs6cG5
E7QOmnrAqLY8LaCqURxofNHv9rQqWP8srdXvJxHcXkq0ZpRedhYfjMlv/f3zwQ+bSmYcuSJ/RlQM
6+R1jomrvjqB57FdRYPAVEKcsavQGm7yJjXtqvGaycjp5fPZplDSHNXpoBRUmg6SrpBJ0MZIWfTN
ZYuPJxYXJK29F8D/wFtveegu/cqNTZbpErEW6w2+7fL6DERz1+QK2aO5L+Xe9N143dMKWjAnz68D
gax5zJCX1Or2+Ykme/MS8YQAv+IYTrDhwGs0fCTGb388haKcp5CB1m1kLFvr9PfE7CLJF9ohbznE
5vL27o+97cbmGmGaepnaP5Ll5Ed9ZOCfeGp8C4K8hGXqWuttpAt3ijI6Z0ncXEIMEG6roRqR7rgO
ThGYe/qmwTa4IFDTCG6Qg9j58zEcCzZ5sl2KHc+QpsqF8U9VLmSlxVo4b52m5v7+aP4jb6SbQ3yl
o1zxSW3jwwZS7NrIXfTX4kR2zFIkIAxMNWGv4c+bJHDjI8ficFFobLx8JjA0bF8XbmXs7v4EeaSu
oIAkFF6n8DAn6FQ49U9vrvEHQNchqsszWFNSu+qZBNTKxNTYIeG/StU5K5WP3KRbhhQ0L2a4FFzk
vmuWzR2dxPOlax2wJCK1zWPwMDTGHlfs+hJhdlnLw1tvE+SeKPWvsJpVw7cx1IU1pBaVSULJwVp+
SLASPLcQzIg159ygr1g1OlBfCoIU9Y+T4+xFA6VFWcDRR9tLwKNBTYYCzcFE8qykB9C1QdEzDrrY
r7kT9GRQXsh4FU8tuIA7bpA8o2ii57wYqaYg+Xlv+KAnMjmzweteqKgZqeogdLkA2/PCovZw9qBT
xk9QAndzNFcM9CDrNScQwS+M6LeSCGQeraQRNf8z29R/Me9/ZP90WUTKl7PrwYzFH0mJ2qJGyB/k
ggbkdoAXE2fbNGLC2BdBi4rMc4mdhlV4OK5L6bHP/MGAj+Y1PGLSqgswVUqkEADpIdqvl72xUIlN
buSDwIvqnph76hcX586BakrYSkU+Ia0leoxE/NkviCxC2zMfpfAZT8w7ge/as2d9o5yiKD1GVtAj
5aCy9NNC5SZ638zCMR/euEojrriWMRcIYXstzv/C09fzAT6a5E4r9nbMqonoWeu5ZfIF7NJLBzDu
8Wj8bSZjTzJavw5tAjBZukfK2Ba9nLucZpqECdFf5NL4tkcAWCwKlXqcKu1AyfNAQ5m8IPTUmQLN
8WLHK57OqzpSDls/aG/LtgGFy+w5km6QuoNjp7UZj8dd9BhIwUmU1NSyPehphHv876TFqYt85tI2
OoMPsSzJGsh0sX3GSpJP9w1kticzKnWItfCjtzR0q6np6nZmP6+HZ7Mjg3xc+OcJ7H23BOTPO7aF
+CVx2cHMoHwvF3/Q4Rwiwvn4vdEL+nLP6EPw49zqVRr6jxW2dIHZxJirylXp48uMqCKRMnjLjy6S
NACvUzwWl7KeWRG/QMHbTvd6eC9ufiB9T4lk/URZZx+Z1QnjtFk5NBH4k4ME6WjZRPHuImxinZuQ
khjnzIothnoIHxtXi+9HteJqtk73yuiBZeuNeHA56VjSjTXCGrO/K8eWf00rdYxIsfEYNTzjiev+
M732mKYbtmBktNlPDlZr7ndeboT6jNRjseuINEuzUgBf7pw7jgj/sNiW5GxRjWWvwgzr7HX2HKIc
LxuXmUtoUJIFvL7EFeoDpNb8oAwUjLpxn1H5qT1pSvF9+qUW2SC7ixHRqcZ4rvKGzjyLFm0/o7DH
D9CJE3KykYq8/sTzjrlCI32KL4jln+JfCVtW0wrN1mLys6UN3p8+MHbhLhFl0pUGn2QCv6ostsoJ
1ZpysAiK2PCx8rtRIUdbNeniRaX4jd42GEMtdf8ilW6/4yLVYWMULMOQirC8au91Hp4JTGzWr2V8
FVs4dPr5Kovp8f06hfPI4nwzQvlBT1FXSwHpaOvN5FXU9B8CABiqVlKemttf/lKTpHwZCDxZFiPt
VriJ2oyy/QMi7Aw8UM18J1ELOCHgZYIYV6p2VuQ/+gijGRoxIupQJdKQ3rTZcb53YfJFGimrElgM
MmfrPB6xuWmYNyhGzXfuRE6v4s2zxpQyC7W2qLcloMU6S/NFbAo9KEFiTiyuJwvdBo+jcZfT+u6J
IXgQ/FhRR8NK+u/NECqGsjDEoYRHyk4uRWNjI+Hwl5hPYKQIPzv6Hq337J2uvHsAMYI3X/DfNrgW
9EsNc7S34w3qbJ8RZe/Fr5EL7PfOTvH1PIjCPrE6XGrnebCZ+Y7C0CRV7zC6HlNib8caMcnNEp+u
rQZnStTebNc2CUj0+g3HoZrqOub8gUmPcC9CEWQbS2W/EqxwHjePl39FFkaF1ry9/NL3R3up2Afd
hMRIgaIjc5CSTJQmtsODnfqLnh2GNZaubvN+fHoTHoMYp1oabDF7bd4MeNNuBuw+CRK8i/VcilII
DuL1SYHeDXoCTk8sG31IplU7pyjho3iXrRrXKyu9ac4mBtcgsjJTiC5qFTwIAqWmUblc7cBKmujF
tILQUGX8DSd+LQVLgs6o4TVZg5Q1iW+qHzdA2C1ImyKoYVt9CnPsrK2Qcu1IQaMwl22iDSpg95pm
cPwsZVm7B9UoJtssQjLd6K66KNzTIrx79k6fib6wKXwfPZgUzDEQpD1XznUmfgPFaDGA7FbVUokp
+ELi6jhQ5nRQ4qHzyqcPClQyw2bdmG6YdsWO1KeVdYwiRRgZ1U8ws24nXl78ciR87LRqvUrRmnxO
YHg6aKbSayPVxL04JAJ7G8lIVEyJMeB/XjPQAfFJZcPqqXoWUCy5vYRROdlc8os3P/4QIdNgIXJU
+x7GbTk8iY10c59dPW2rdlTGzmjGKeW4GTwO56VgSyHFt7/k5kLVsaBThORjbRCh6InzWshFMpN7
beABq9P6NYK+zNz2aynQbMrfu/f6+3ytiTZNqKYyQfgj0h1AmAEEj6i3xYzE4lZrmykZrMETpITC
frpR/A1Ej/SscLp2mwnoDjHC9vPC2X55xp4Pk3ki0+JDML408/RqhDz+yYVPg/SNkkaL8yzcuNjA
6Um5XIJTW6gTXUi8ONIIvSJPIayWhYmkRnZTyHF8dp99UJH1DCD9IrBpp8s9PuYGQHgr1dGTwszG
aQp9OPNcEX+yysdBATRBlNTXHIwrIziBw6RSNE2hFk2JfQ0SegDMYDdVQQgPcdZLAi0aM2K/Osi2
AU6MeUzleDQLKvfOHsUcYKAMAClPulsMGm4KcW4v8sXJ2Msj8k57BW6ilFhdyo2SbRPnsi1T8pO8
6pq1b7NHOsC4aBmflNEMoZhpu473ubuS748pSUlYYvCXo3ir4aLac97luw3DQNtPlkok3HBJq1BQ
5a2Lb6G2y/Lx59/oEyK/GmxlCWdZ0wnuBbRIP0m+8aQd2cFQ0K/SNuNSSu17E/0J8LQZuiBMUCBT
5rBP1WbW8DEEeKhZY9egYqv2Go5x53M0TTYuPE0RdMV6jUABMAdG38Uwgtl2WC7a6jy4QjKr3jjZ
fUnQbFwAYlIG6UqVxuzO/lx6QTJVkubyzE3VOZT6awDBmDyRen5lyjU8tbovTViw/md+cKYo3NLf
RrwuK0ZbleIsSjG9OKu/JGRl39yLO//889Z5BvIj6Gld6z3PCJyJqwN62Qg4UjO0M/qQCkLk2eFL
XLABArbR0sJ3KZvV7fzUkRgg4h5mvSIHT1ofgajAsjsjsdNJql3vwh7J3VpryHOzXJVXqSpB7Kn7
YCVxNnXe1bQZvY+H09KlCgLqQrzw6B9Oq0QBF3F22Y0zFr6ZYyIuxY1mX9wnxeFxC+iuN/xZrlu6
lkCw30YZeyIWoaSNaYSKFbf4Z+PHjgUgF6lkLTHoo8YaaZ4KJNQVINcZFpgmL2gRPKrZIN8x8CIw
Z34nWjBDHgCqUiFPp4RUorRVIZuLGPTsgCt33hc5tu+26UsB/mIfM8S+pIDEpzg2WfyCH9VZimjj
42+5aJ7y7VlcTdwfmlOaYhUbb/REYmaJiFK9Y5dsR7y/TN5tJgE9/VpCEi75IuJzPAQseAnDGAlG
GUzOFhD7JRQJiAbHqy1Msx5+rw0sMcuKJX9KkHgZb15c6YLJHpb9jjcOaXHT2b99jHoe4ACHBUXi
qkE6xLU6mHrhQoZpde6zgOn0PS89IqXXYePGYFpddNf+7E1Q7jda8sEbxK8aOaxcUf+fPSrLtnHy
B/vW1sDp1HgeXRT8HUZF2VnhlSPSO8siHbC+Gl+8aLjUXy5+MmBXIiGIeuYSGmmqs3xPRbKygRNV
y+MgF6Ds2P6g1IJixZ09R3Jg6IBE+OnUaRkZ8XhkYw/WS3lruItWyLI4h1ToRRSBOs4lDVl2hz/8
oWACyb02VHe10uIY7vO28HTTYx6YTU9PhLfPYdTlEhuo9uCy8msRr5vC8mi3aKzFZA4GTqD+a0He
E2topXQElZr9+OwpitpTlg3P+xc5SWLqqeSL7UdyfqjkokJ7tyd+ylj2NRKraJKIt1VLY4uYiUiD
fqiUmvoNg3cUKg/rJF7ajQADirRGz58dHpitwOnLheoRrSdL4Pwc2vjaBqNBoNjfxa2HBudJowhZ
L1BcRJFMhc6xE7NkpjSoH4Ew5xFdlbTon1QKqth+hdSXYmUWXoXq0/Tafn7cIq/IjZS8IQru1716
rQUZRfcqfOGXm+WImvQr4B5dMXhGYDrNpT/3AEU5DRJe9QGSskz904qHaeC7zXeu6cP0t+hx5Kdg
BkP4/wwrHTUU62CaYKXka9m706VAKP2zUMfgIbN4RqVRs6+JlJdLjeEjEt96mItomQdNiS22Lz8z
/lRingUxELl49XsDEZbv++PZz2P1bmR4zTUloKef8/31MUuNqghEQprfxmi1L9YeppmkqSp7POi9
CNyB9HPSrb73F+wbXffT8Z+Wo/OUzVw9pF3Q+GzMayAnH1w3xUOHde+3tWHLK3WBz3RiFc+FhkNN
/HLR+v9qIEg/V0Yv9k+VH3INEMHZWtA79q+jT0jmhTAdozvDcbKRFxPRbsgVnuf0FAoC9w7YTPvv
ToPpprjRQsFOebJFNuUi8OJ3/D8MJu9otxtEBaeiAPgJAZ6UpB7VNT4+6FcJltI6tpv6kmqzqQ2q
R/OSWb2C0+d+azemEhLAilL9BuJouD8IQYpLlTHGcxjWNSjxjnF12Si31Rue1NcD/fayCIz8aaY9
vPPiW4j84ydus2MTEUrydtXsHD3P1rSkwUMzVNS02tGkb675WL33pOFOAh14Oif1os696XRsT7G2
4Lg4l/3BWz4M8pDm4Rjmvktiz2r63ayna2Xz79GizLvqp8/cOlE53Vy4dvXYWSm9yOpo9cxRWd6+
UIN+XFj+geLuAPn5CjIs+TQ5fs9FhetyWsvdAmOg5I8aL8w8D7a2z0Q3rHc9ZF2M/aEAh26a1ohS
eeHqKOuBSc/2GTleEcQdKwkGwy77SiWL9kyLXEoXpnRy5ALe7CUqrcHolkaR2pU00G5QW55x2nzj
HZ+uCBvGEjYukyLdpg4MBtAzRoYBt882pHZvQUaviAaLeFEkfiwXqF8IcHGAdRhQisoQuQq8FA0p
UXCMOxP8dDbQIkBvvWHY3By3ebgNIM5zjCd2FO+/mrwQX7zezpbcOEbi8Bz10MqxIC2354bay3Gn
o8PjDYBi947Rv/oH1+OUV/7M6SB+uP03EKCLgj1Tj3k1EH3Qc8kJZF44+oOd6MMmRP+RDiUpnxw7
uLnWQRpCgs4rCcaXto9JlmoIxwCUyosKTApSqOhyyjxOthgmdLN1FrWKuJRs6yspmw3DUPjaRCl6
rs3DAIawAikSRhX7EM3dVI/fM27kz/74FHtzNHJPVjMbquY/8AVV58ZvWQd+ygHIe/f/lo21cv7C
L0bRQP1fPmZ5JpJsBoi9rDen9pYpq/F1NviFUBGu0vSSlId5vKnBmW9whfhVdOhefBih4/7eNp+j
ProSWRDLoUNBNRvmL4Zmax0IHfaOfnSglRqpsU6JwDJk6Mv3FozNIZB9HskFAN09WYijuCPQfPqj
GUjMFV2bEql9op0lqXcpdoiL4Ld008Z5OmlczWaIVtyxvq5i7fmHYXgMsvlPnHcSRpOyskppfo1h
Sq4L3NkAs0dvX0XVMZSKehMvyKq2OZHYpzitcsjy1J78gt50gh1KSYKjw/A/PuP5lgnpSkUMnQu9
coHa2C8E9OgNFLv4I8xDWauMDnR9/jmqzntcGnH8mlq9fHWMuOQk4Z0GYCp2CusiT7Lz+hxkPGvO
j3VqXu3ufhylwj0X2H812DX9zpltbKnEbqqcPhj28NGLgOS0STSUm8d9lWBhJWdWn1SSi5BtwYeg
ZfPU9dYeHpz2JPMr8aoPYsO9nxXE1uek/0AyWktn8HetB/+5wDpZkcSmGC+vUrMv2Km/RrD84hXk
lC9TYhGa0mE3Lnmi1dfJ9rGo0mOSRtHwp8xCtCWxul4ZVi2+JzT/QW/Lnmj+I6mOItcOB/gM+spe
RjFGw76gJRW91zb8EkTRizDvasG0GsoCcQEpXbPJ1cbiLOutP9qwgt6xPB4N3ypQixpvBOaek4Ek
tKmjZp7xbK+b2/OfpKoXTLLAaVG1l468MAsrzIDLNIFGDYSlJ5nAq3AND/mdON+DvrzZ4UgHvz7z
YrT9yGsticrEdCormcbrQS8pcyxCi6BEn2bns4zdNoQCliVM3ikxceJDs5Ckkm7dC6uMkMKThcPm
pmS7kPCHsaar4YRr3zHNYGdTmLKlOO4shu2SZJ//Q0JiBTYOswIsqckDfWzogkN5R0CteuaISlBH
0jQScroQBTPSxb9ffSH6AS2QbpTmg0m8U3vhBXSlHzkUB7bydZdw/s3xhfvSY+sjG0WzG1Cn8pqk
3PIGCG+tIYm9Ro7INQGdNFHUEBRbaKu9+mPW6KRcgylPczj8H10CvmgI/p5f8DlC7oetsUzRfDmh
TmVgl1bkKNa4jPfEs3V1rMRVu9LfCAMtL+VSjSHMoCmUp55YxjwQ3vT4dUS6befEUowFaLkZRMRJ
eFNKwtzOzQmNr6v8aPjFNJ80D7axNizL+GAgG2+2eRWJTGrjKlIz00ewO5cw3EqZMDlb1oKA7SvN
CQ5mA1DTsdVE3QnZ1icNmfKzFAd4sGLX7+bH/7/i5UOmgKo87rC2fma2qvhVdQUxlVrd2H/bYr7R
fyeORL6c1jfxTSJbEVAGQ78jz/xxBOMi8zBtrKvZu7iTMv3gVYaPG35UdX5Gx77gvW2kL/8h6LWX
xYTDje8LpsRzRQKOVgZxfyDqXJYzf2kklEbkd64JMy96aUlz+kKWUBCeg0UHy0+cEV7XUIV0woLB
CiJZsyUp/3A2vDirBg6uGUrgAcOl2MJq3pom+S67S6y642w7hBoj7jWkYxRwxteUXlhR+4fG0F7/
gVYE6q+6PvPQUTABQxilBov94/pVPGYY9YiXrY3Ew7FluvCfLOaFoitOxKEstO+mkHONJxapYd4t
TKlvnlOmi3qCSpAThzCNyVnMoOMNQo011SLwE4/kyJJzluOBlGAQ5j3qfd/LekkTaXf8UnKM1odm
S04yB8KnVej56i9dIVySq5BEwdWr6dOnukrHF3ZSmsWr/VSho05/li2cZnaWMMZCX8WMyI78P38s
DbbzA3IbgZNG4jJRo7XuTw8fGKBXuwYfKbPCb2mS1bXWhXUkN+imACePPCqDUa8BSvGcmqjpcQ7B
IrHvwiFINY7CBwEpbZCFPPJtQQnd0D5a+i+tptOvzQDtXuC+6Jb3gAe7Lv4AG7dlrADmLN5IIA4L
08TT5KpG3XkdbRQIAWgHtW18OF81bqxZYiA6hbF2hZ/d3KB1lzkytRgooywFI58kW75MnucESuiF
EhRO1T+3KhWiHstzS0nf1Ho/GIga0PN8Z+pqudeR75ceYgch9puUtCojEzioKW51fCZmdgdPBaKe
WhYoR+NEmsST7e3BZZgaxL3L1z4qesZK2mjGaSRCrx3nXWtZuE2/rsQnXv/rCQ+mGk44lnwERCe3
tavpvZHHJWjLitAh+14UEfHk34rj2enEAmJN3OvChGkIuHVvw4uUVq4ba7JRYloe9e/SgPkgN3OH
X0MnRswf5CEPevXCj6gnAAngzTdTvxhWvknwT2P23iQTAtbWhEVJNZT0JZCP9noHGO+boSA8jEWz
PV92epGFXvWTEa6vBWfgkJ6p7HBcpNH2DRnaACtwOfBcn03DySVDETKyiqwrePptghOua/UAhns1
vmXSLy6O7aZO8ACfHXbbzHItlRa5KCc+l616wpdl7zKf2H826ueCg3xgzCUXy3hz84QjM2z8kJNJ
/qOtM5isL/k699Rgv9ZuVjq4MQKYWurc4IWoHpyFOgMZZ9WkdZhijcht++hPeK1OW9Nv0EJWjY+s
N9b4ZBjusq43NUw/Uw+uhmqCfsrxB13hAqCybClENG32TvR2TBVHRSX6s5sDLDYREHZGKNdtV5ox
UcXPqrdhlxbBB3bRMi8CnlHiYbirRWW+lmLwoMQonGXZp6gy8SP58jd7BAp1Vp/vGbCIQ416OuIU
dcj3o6CIOzgCHEgyo8UWixpmYMGYPoeP4GMIrh1t9rUgDBLwru9p59099nd8Vi52iV38+FEVyFzI
sk/3a9ldLeoIw7Sw6LzxPq0vVRAe2kdettuRjlvbrmE6PhR7AuUZAX0UsCDoqceD1vNjdkuodTpU
eg+92MDUfvBm3tiExEgmrWIPzDoMyNXi/L9whYT1Rv5MFx2sRwC3kedbaTHUYp0bs7Pic6GYA5g/
cxefdXUn2ALZu2Yry5BKbNsRh0SHY7gNNf0688+9vZbNQbrpnfsGlUug76f8vt0g9qgWrlAnYsw4
aC440Kl6eB6QnWfV0ywDnCC7+jtd7g0wIQ5FMHUa5f4hg1L8je5y91Y63BU+R38mt7hSDKCOu1pt
uH+HWYDvgy4vZvErwGL8bx6wnskQuNvWWhlehkd4wzAKSCLf5080jPAM0hnXxDHsKrUddp+1FcZi
bH82iXqnhW99scEfekKyvkoCSzR5hVj+lRZADIRxan8WeUGXbnOgqdxVR2IO8QXisQeAhTNOEP0U
Z5A60ic/2CfubM/9VAPT7Hi4wGUXicseeM19nSm7okRRMCEcWtesHHUOHJB13mZ1V9GR9pkkULzT
RUOTzxFb8DyDLqgQeFZ++YzrqMn14IvP6gzmkruX5YggVh5T5qALMHrGnDG3txaoQnJjMpTz/JfX
cwCymWk4b9BGbG+tQGz29eseiKME5XHkNsQ+JrQFeGnuuSydJUG6u8HjlwKNPBQvu11L/LuZ2SaP
X8hcxu6a+AUXmaNYRNVSbbEC+BtqDc6Mb6Wj0ihwV11CAVC2Yp7hN+XTqxW/GImNgPfZ/cOjU9EB
EpDHcrVQzbfICpDyPlGF6+/QsIzwSQwxLPjcFjgi7OvXuAJ7y1MSTqUyWGt0UX/qH3g9XH316gaH
lcWDBj3rQHHsf4TP+pnCn92rCb/kC4E08di9lG99knQRn4OS21ORr4CJojPnGXNVxhs1N679xQvb
8bkcV54OCb/m3b8rg85cOvRI13jRL6Bc7f4xXvuYWHWES/olZEHulzLjANwCal+qhOAO0Mvnr9TX
EdFK1Y/MlA5lYOD/OD+f1PZZs4A8Vbs1hwhca0xtEWDq6zVLOse4o3Ev1zSggE36N6J+PjoJGJ1n
B+6fDecE35dPbypD42N93qrGAP1BvgbjAQ4avf0c01k+AHZ26YiRDyEG+HnSaP6XWxoPLNKv8v69
9SYlHxdlz/QSucCsLy650Xp2WWfzi6Mx+PdSlgtBmQcksnj3Ql24gtGdLXq5LyZTIux0zaEQKmoH
N65Fyet0fNR3C18dyGshUbhLHgnsyXi1ym8vYxXUaN+HJJJBd3BXQ6snPezuuN4KszDjhDYp1odJ
NIU1Yr7FZ57jk6dRI3YuiOiDutobgtHGtVQseta4mNWoTt/jEmli8NzwiDsalRdP0f8HBRtKvYnK
4fa+ZJy0TlbvUnSpc2crcmWtzvOMgz8eto/8tcx7Xf2lAbMOkrGRQZDIaEBKMI2x6iCk0Nvne3qk
P45a7o+6ITp3AyVDxIYkrNvILEoHz6wja9wUfuIUelNOpuaUn+FK5CzhgYUv3MI+PycCkW/5/ded
hRO46wF7PU8/BdeFrq6T9EH6GQCtHLRJsjx43++YkFCnEqOZdXUcW7y0nNtKOu9X2B/Uq3anlntm
y/hINFDI0Y13ie1cfuTYjd28GUqI0MeHw3To8JM3fVT8q5kg3kiKZsTgKyvTapE1Uc6DS5bRUray
Drxs22lMnDyb3u3oZzSMWvj+qlE5cCyMQ7B3NzH52u44WxyWOXiAVTRwcVZ3pVwhbo1wNJK/emtB
pmyceM0ORO+rLf80kIS75l60n6rv3MMzrYIjnh/aIDmmvEbJ5zd4GuPBHB1rpBXsdW5mROxghAoX
wzRwCzVopd6OSBGjysNW+lxz9xFxlkM0yBWivF1A/+fB04okdOLJJGHFFPAvXTfmPwp/DMQQjzti
e6AihYpziMwjLu33e+Ah/6RoZmxVF8AE2LjVH0bRfyT34Lz132oWN+Dm2TL08ZfhSUtASKLw70V6
2+BmtBqKr2FubSezTGzi+Z1XXO3a+g17iFtwc40SC2ZBrao4L0sESI7b1mtROsgFF8GdUFuHlMGg
8HdFfgylgKWjvdDuUChO7bMJk8WWpFDub4DaBHJgcA6AXlkSzk/9wTKsxPp7W+JphuXwPB1+6SzT
Xy08v1+PSPxz8ajFP/NnOb30ioH7/ZlFGoq025y6ZkJMpecWE4tP0t/HOtztMmp5eMtUjbj1dWRb
YN3KMKx6jU3XVj2zv9al4ZFqQ8iW6aeZHr/fIqz6e3HibLDcaaYiKEl1fMUZNo7n8FUy/0GCwdBP
ues27m0aOGsIaMEfJcGIbdZm7GwWst6dUbQ8CxDaUuGqFPfG3bKSunaKuANUDprnmytrmhBpwBEu
+48z1yElP8RRpvaJ0EOLw8wjAr0oGV23a3Phu01RGZSB6wjHy4+cUyGrW548zRgj2CIYDSbKq5eZ
3PE5IivScNnGMfwjnc5dPA2rjxFU9npEis2JSxozyLmzCNeOGMjX87+JE7FVycYXCT19SmDTgE6C
LZe6G+fiRqkK5MVhOphu2VRN40+hqTEQKt6SQa/8uBSkf50zl8HM5MGWRPQYsO2I0V232Yi/RFYG
ZLNRVMgRQibncvHYPw396I2qQKOtTwM4q/XJIBctF/Ty+fWn3wkJgQ7kcRnFl3GufWcdYPM9QTxm
R205UBCNQsPEMCzoc5MqI0+8n069Fe7QUzRBpTBK773hFEZbgndfiSzAasFO8kza+KSicrvZAVSU
qJY1ekzU6r4HcqOhzFeafZVY64Z1KS1ejLeUk6eyEAsHQzbEcs7nNInP/AcsoTr12vfp0Pc5wma6
6cebNvh1af07cRgYHEkRnA8kPGkzgWAe0tQiOxWxCNjmPzLFMjkmCwehgVfSGbFQ3KMhO2KW3WJm
LveGoYhSbYZVEnKLuqsU/jngpqxz6Ch3ncASYBbRQj3AcoLEkVgP/l0YhvnHhjh0QfOQ4f/PqUWE
jptLr9fUJEavfHooHyKZex/7TsApS3uQeCnCgyVSeZf+1KJnUpvgEnYib6jA4CcKYjvYYUtv5ixU
KNqa20ZIumb7SjWFznN9JQKY5q6sSweopP+NRIppAMJ0xBdfew8cBqsLM2XM+KFhwBiKtqAr9MxE
iZqhlnF/cHjJiqHcvhhNw7pout/nqEOzInbj27h5dEi2r1gAJ90rjjsXuKECMu3P1gIvWIV6bLRC
idEgc5xT55QIsjRLvJonSjhYpUTrphREhStpVw7vrZVRu3ZuaJdymspGlJiH5236aL4SNl+juLzI
J3ZMKJu+s9CwJZrC/DzPzxSFR8U2Fzfy5tufcLfygpV5A9t6DkPPqrjW28hV3IjJhx8fggEqTqAm
FSgIeWASuMPblWCXfWlW8LzG8Lw5rF+uJm7emUh20CdQmU86Az4GyVVRBpw8eJF13XKw5DbmOKoM
LZWBw7mYGblcJSCgAyaH29hk37Od+UTbjOquELECE3BCwZPvCHtiuQUPie7KxrtZd7hApn82zM86
+BIaGEvIeiqAoCNhvcvTptFHhtmhmevZNN/byOQyYxMelbK1vqwMSG0YCIDZjDjG34MgGbngG4AH
p70rUq26jPD0w3iFgtsOiUTR9mzQtQYQNAxTg9bUuxIy4f2eiHpIL2/G8jWiywd4d9+mpLymABpM
LJ5TPCGXp0a94XyjvvjKSv/6vBfTja7Z+mG1qf4p5PZegW8OHHPbewoVG5CK+4fMJpSg7RTlfwgq
bJlA9DakFiYcDUchIhMwiNBCTm1J2PvcBLaVcxiNJjK8R9M8HJ77JKpG8OYPHpXboqViSeEGVphd
k95P7N9ctXVDRtgR0iDwcq8r+VY1bUoC4slHVbEkpKQ3gs55Gi4IKs8bjLoJmOg5tEr4UwJ9VCjx
q68QMHy2mIW6j3/UWY9D1WpGjOjyAG3MwKr04w8B58k7Vhr9AeRWn4om2p3oFvDA6VtSje+/L23u
efnZ8fQApqLtHfokZ1tVLuwDvumwtbvrVXaNmRMRi8fh3LBlzxIHrfTNne9NZFQJ6ej8jxXTT3Tn
VYRUtPNBE6ydgOgTm/PEtVzg3MF9ykyyykfV/YeUKRv2owFzWPn802hBCpCJKkJ50W7D3fGITQ51
g73Us8zTw457/f9FpuvW+XLO9VMtkQQzBtZW0ny+h4qb2wVifRsFVeOg+7Qy7NQMw8ChD6C3ZlM4
0aMjoVh2dCPLC+5tcdCW9nbPp03cO8Ek7oYCkNw6O0Tv0ZAqtktcBJ2be7L3INZx8ariuHKgSg5c
A8YFSpXfkUG8Dms3iV6q6Gx52Q36DvIs+AQkJNlXaTqZa/+f0GUozYVO6flF3FxOXXTEwLO8aJoG
lvhmDewkjRVvxCukd/Zk+xRZ96WasLDHPtJLZcAGqxzdPIRIxSE8S7IjGP1mn72Ltmo3B2V0q8T+
iCEBTgXj+PSot6DetzS0AAoWjukK6o5zgS73YWktoMyPBg/ymPMcWpszVOdyRUj6qaucHnVq2mAv
VeCvhGhV/6Hk0OJK1B55kQbYbP22EDeagx0YWkWpefFRsGsg7oYIZSuZtA43MneZZJl2DCbVOxkf
3nWLZzAjwb+/deZPDJN5DcvjNU4IFTuvSF4KXnUQ0V10KOSFQTFjOJxkFMhIkMILRzTcJG21jKmn
e1WX0EvDreg8mn67A4nszr2BRBrLxcPq/6ymoYICqT0PB+uTwhEzwTYe/rERQ/SZ6dPiJX1Sg1si
5Lev9h6dGdgIjwgUGCL7zyWBep5zjS4GtLmnqMgI1XoWyo8fNoA9vfalvOfFlIUkka3Zxn3/Lhpc
l5PAPTdLNNq+eOhF21EEkYcN08GV4XihRLlSugznMFTOsVt+uUOjZwEHCqTB46py2LjnCQKugJwp
cRQblo7EM8ePoOhhtls/7wqOYg07QI03xyuaQEOwblEJyk5pFQhkXpqxd5KQjj0C1TV/2xSHr6Ca
yKeagyuqdzPY0wLpvw3MLNJE6GM0ntoO3avoLZ5Z4P8q1f+amnFEhawWTJlLbqeamb0yxvD9H2dK
Pr/FnVzcr7Npq5W6kv+shEkD87XGhrobY9v/yA8qNwpAf0RW9x3/rs23inCpbbHQVPkMLjovB64w
J2zj/eNXo5akDpmuuuW1b6Hsv/s5wkKPs7SofvZhsmLk1dKVrV4P0Uv03LGplZoXTSBKmCMVdq17
l1zj/KhOjspbci0XsREKsPZU6dg3j1fETc5mvq5M82g7VQ91D4uih3uEiBd58CKejymVpthjCcTf
J3XMZpr/A7z+sEgFreJGN1NJX7PRCT85gvkTlt5fu55k25OKc+hPK0HZWxCggGiVjc6kEnB/H7WX
Nz6YthbwcTmOf/BIpud0Wrjg6xtJlgtm+BEb1g3oaCTW3miNB+SaflavuATltR75UO2EdSmo8rEl
F6VKvrOaaO2pBb50g3pfrP0RlynnnKDn3c1ACSMvL/OHMszPVbZCY8P2Mj7hmX+O2U2LU2zVezgA
YFIS5LKS3hOnpai9+sIfdwEi/ISe01j5AOcKN/8yxaw//OURCG6Pi3q3/7wugx+QXFrhdM8EfYJj
e5Gdne3vnnypgxSGjIjK1z/nmI+ZZ47xyJI2K2iEbi6Vl620zjwAdw76dgXw8ktzNAIavie0b3kR
1aR4xcHQrbSJPMUfFI5zDlDAb3OFQwQfkevmH1VM+KNI5Cf2CJh49EiYTEW8f0iOuDSDiLPYQDOd
eVllypJoGQo54+dAn20k63VYhQzy7PqorHsusE3Ovp1mjvZJds90yuSCMOzumrN3dfliBP2otCmr
NxryoaU9yCrt1a8fClZWvjQwx2RFrj+ndo95hK3dOIZGxOjHc6Z54fu1YrJ7H6O+IsG9pnbBkCvk
9KRmx3rmUXXxmbDznwzZOE6o1xZjnxiHotPOFJfntshG2kBvppYI7xxCV3atWSCZQO0dI4ZOcI7p
ajCHhzwb0ip0u7YvzqdftUngwvmXdINxnayXolEbmwIVFeXA2XiS7DEYRy88sVtNVYmenp8/xf+i
QOju7wQ2AKlszRNwKMoeSD+MFSvAhQweF3iKltXzoix8gt6GFWwmBqRvVvZ8OpLOB4tWdFhdSVlj
wvannacDu7jOXntIps0i1uY7FuK1mBhXoe11Pz3bEsRIQWGMI4xFTWq5qaY/egmoZ6IRXMGzr/ne
jk5/ktcCWGPnUkzMaie9wBEuKMNYNbh+ki3PFrzx3Pnbs2SOPvyop6qjH/3I0cWra07brucVVbGm
x37bLXjyNJeRpcVVQDagioO2Nk9TzpGNGDk1TOPXo7MKzr+45GGhlubgQnIeUZgjqHm+ZVbgKopO
UPRd+XNhzEKnJXVooU3hTl7+yLptIWOh5g5lYb749ELZDuGNVdl+E5QNMm0kGGUnqQHPaBuj9Seg
kXxyssf6dP4ZgLiX8beKiGX2crOxZgQzZL2TDOj6hwfqcw2mVU3hepT+kJ1q3zp/H+buRnT4ud7O
sThsHbb2dtNy6/OsWZ9rg7W+Lk6pwPS2U+nNX3IYItYdS2dNzPI/Z5aMDr2DSdos3ptQimOBSnwo
fl7/2QEwRCNFHvcexYrXthWy3IKJxdHzvDbTFUUVxKtSmP6kEPphQgkE3RLRbB4DwuCczXxoh7uE
bt1L6McI2jzBW/OQmveVgWaBtN7+BiaC5wNtjK6jJw9/XaMXH6J8uTZCTSYDM2L9mTDxtS2sN884
vN/Ajvp68znbFORYsseKMa8Kd2i+F98ACAJRzrrV/ObcM+5xrHwkecEgzFQH+hnhbyBOzthAnUdQ
kn2dmeJ6Ppfe+9t8C0M9wtL/CxTOcKSkFVuCoUUivTEvUeqIEAJPg1dnVKa7F7PbDyndZkcP5cmp
Y8HWACHKKw4ljUPqLr6YkAACtgRBHTo+HoJiA76pF+WBfKT3Y8UeeuzenVmMlDOZg+TCTgZukpGd
W+emx4CLfPLjL4R0YxuQSoULDVusqjtgedQNW7PftsUzD/JQdIWToBwtrshkcsYXGHw9aKGoVdwa
2q6+vtizWIGGLPbTr7qRX7+Mcm++pVwrn1/HMbiIJYCF0hWQ4dfOA/076iFK+l6PhVtl7iOQs/Dx
x4t0vhNAKMo6rFZUSQIv6fWHPOKX+GifGie2+BvDxZ44z9Zbg5feN4wdwaGoR9CV7JjbB3Dl7GOc
stUk3JIUEeD2e6TRJviPUcEkSn4YLE2ycre2z+WlTYrT2ABV7U39RpZnDJOiBEq1PTNwRbAGRUvl
rozF207jfAp13OYiM7+hPMB8H/xh9z4nvPTov6d0Azj7X+8nlXAlak40yzJ5+XMQjpq8STnns6fL
eaVAgzpz9luAxBXWY4ziLIq3XXvozu7jAlK2Z7LQTvwDMhZRMLOSfwwfB57oyjzUd/zXRiTINOPE
k6x6oBfAisxjiBJkoC7GPxu5zdcvUscW65UcwGoIA/Vln3Ma+4eW7goSN8BXHC8Yxc3lfMS1DQjf
dNZ6gqSczuydY1LmsgAOwR1aZyqqn1kdu1eV3KFRANGEdzr63M3aMflE3l0F6f3WEEgp8TuQYG5k
w+EPltrjAAmPSNuw5tNUcrDG39X//EfrcapEHZtvTKDCCijihxr0TE4h27PmuWKuNUaPXvg9nxB7
+nVd+Pm+DviQYOBd9Wn8tM4au4BX6SgLjnK2J55Jj1h4x7WF3EYsMzJ8dfAjHh7va7aD/zI86fQS
J/KsgL1bRJRNxttEvCrDAGqDXUd++O/ECMm2spMryDqjDUgyENkac6pbypV5uug5Mj/mKCxm7Wwo
EEIyWyQGxafP7JW1YHN28wBVMwZVhk7itLFxyqyY5XobxncgCq1l0j07HLsQ3+GWhu0u50h7XDnw
8qtpaDFknD9BeZaVsCewKdkpGv0fUP/9qACwLJH3JAIBMDH8zH3MDl/LKPywb4EZABviT+a3ijUU
aDWMZFdzSyTnEkZqulxnJLSoP2wEncuan2gEnm0sb5d836NdHY+c2qDfHPY1HOjr8JqwdvT0JJBZ
AbJ8VHEN27/8khTTMehCqPO/vh4fPTw/bm1fDtR20M22WK1bDNFhPxdtkJGAI33SG8z3sx0NBczs
hCgta26gSdGfmFCYRTGCBRIIvY8l86wr0TnD2h18Bgf5cz0F17UFlLrnS9JWX+uiDFz3yiPrQ+yp
aQ8iWwUUM6jtB1dJy1K0AYXGDCHaaGy4n+62DoBtcm0A6HCa0sDOnNCwzqOsnUeysK0sTFE+VYM6
wW7ASFm93391ai6H8KC1CWEOk067rxAO9YGdayEQTyYdmEpp+YSLRfm7KWPgmlGfrj8Qc67squHv
YfsgXcgvGzEdBnLTS83xgXhaEapxqcfoUWzGm0lKZoXzhy/hjyVLCGZdyshFZDO9JDyZWR+4AO9A
JgDA/rNs+2FLKNlAdgMGGtLmc0TumiutR9cZaE8nWSpFDXYoOFQg+9Uu0bP8ppY9jJbOSjujLzwf
F00nIyb8OWEFyNGL06KNQoiRldUFYfn1a6R4KpSK7bZD00y3eArbsffQLLwi1YjkCqnwV+5uGiqw
CBItEa5qOWcJbt65y7bCjREJHsVDJeSiP/VNx2Bbo/ZTUH5/kYfaXFJV136adSGeaPDB9NXMEeR7
jYUgt31xU42ElWbNPKvRU7sM1yC+h4cwvEWQho2K0htikqWXeVyh+Vq/e2XIgNdC89VUOdpbUQOD
pUGkx913CLk8++LcwAF+s6Gq9PWMdR5ChqUxBRcZoABhkHKlNNLEk17nU9d4irGMbAOlel66f/Bz
SuVGam0bBEC0GCWIOOt+UmciT99z1UFjgRZpEgMk9R+vzRpn++ALRBdyEJh6LKMyHMYX30nJmvQz
bfSy1KfCsNAYkYod5u2EijwvxFpODPnc3/tOJUpw2nuZ8mMQzdELuTCWaSQzdnnqTXEH7SfFd2P7
JvgFNGPZcSKeDhpTA7KaZxvqNlYd96Xp1vxKlH8r6Ad2hbTIhfLqPn2AEvEypTOJELqEZly+onkd
RcfJPPdFRD2fVlauJaSlq0b+F53RsFLCddyAAHjDx7K5bTalljpkIQjV/AqeUBJ7+hhg9fbau0ik
DkwNk3PwSJCEEMf0QVzxfwX0GC5WRy4PuCrTFwmVumormBmE+SeFPGq43gK3eJm7rQ9V3hnihZYj
fQMIUooPBggBqW6VwRFZXT8MyQH/El7FmdCbQflDen7uJnnLsTmhb8JphPD6GscOv0EgYCxBeAYM
sizHacFfdgOfyXEFxoWtzOSqcn9mcEsBcxtvFMnWEOykEYtvpqTYDas20+FqTf8qfpv1CAutd4il
Lj3ASMkixK2b6lemPL5UTgN7A43vaBLFEqZm8qzLhC9F3hYCzF3fWLPfovRoqHvKW5SIqUdhBtND
fbDmebqqotiZR+43EayVOobBkoM795dCY5sTOPEf0ONGjnOzrAkoA1Z5Zi0oM6RYvoVDdJGN+z81
kvtFh0EqHDIrQWDNf/SkPYALY1PkUPzotpPnQPM9JEBqW4cT+630AgMm/DrWtEI1lmiiotafOGt3
eEu1Kt7MGePy+tmRLe4Ubk1QouuhlcA72LZ6RavqtqaCaXhQKqVIO8XQwxEv0QUpB9PqH4RFK/Qp
qin8AgI8/ugpp8f3HTPvg71EXbAwmOZpfS/3DP+WTv+RxOgM4MPCAaQM8Zpg0o9aZBtlzN9ZToKa
ef5rLLvKxi/Lzltr4MejFezSdL0Q2sCwvO0Kvg9A427WtmJHtD0F2n4FuBLUSYDTG4Cpxnh2OhZL
dZ3x79KpbzdQNwchPcfxTOsnw/AekpWnZ2LOyX8J4EbuDG8fn0IL4Z3nr9/dSSc6jxCHktc0WCG6
54+hD00swajvPjQqEN/iZFJ8nYWgSD9qyLCFykA3qb+/qN2pttfwlXW4wpCDrD5EuAez4ZAUhLOw
9mmN9BVGCceK2K/Y2cQ5L7XqGbMC93IWWlePrdwbkNv9f+4vpGfXxKRwE2BntHXPJT1kvB59+/i7
rxI+mcdWyrx1UzOnqAdGV1NNN2Isagm6DY5UHEIEYHD7i+hlTaIYf4WOmG/VI2OvLQPPWOqLw2mA
19D0vXJnIeAZNZyz4xrtPVAV+/TSr9Zkq9O9+DenYdDxqCII0mbCUahmzn1zTCZ0JhX9UzAMnxLL
smmdhGUseOQbOKszhV4cjw6pDazk0cYYSzdfKWMf2xROcos6zEaV+bsIBbHJSKIxrAp2NWoesRQp
hADsLV/yCf22tARKOgmYXfOY11OxpA+0qlfLXufXwAxfzyZA2y/ai/ATsUrZM2AjZjsyvaqDJBSI
VsWG4AfGdE8qUnIjr4ph/WquD8zGFXxwTESxjUyKLXm8xzhnkIMTSmFxEPxN4R5AidzVulmqX487
LKqpQUWpdTJCnMJPZC9TG3lmZIklChDXZR4JGPaz9N7DnUrNwB0jFEbGtj0SVL/1BuT/IjbdHDVf
Oe9BxVH3/m5VwXEm9P2gWUsxO2qH2dSYFtzKZChF53QqiQJ1z7GlDh33icX0D5qH5jQ+LiCtED/r
4uaoykFT8qETEUKSJlvxyX4e088zOM7ZosZZKevIyZi+b5aXjNQYZr2hsjhfz3Orx2rQ4IaKAJgs
/Um9/VoOcCQN+B1EAw0QHzyzNG8mI6R4Ay9H42XFpZQO5ygZONQkEM7a/mAE8QS8wcDu8CI8JEPI
Kl7ZgB4jGOuzrNzmTOSV+XrrDP7p/7M9x5aa7q11xn4s93d3K86TRrAZfnuH+M+3PFqnHezU5Qni
tNcETNBdC7Tqg78T3srLdT+kx4WYcwHiIiA4ttbjHa7Z9o9H/P1GIGl/A5cHTyQgKJ6+cbMzatTX
CeWgLh+xQfE7ClpaEhgpsvu2a3GqOE5vI/oymrGPJ8EgcHoP6NWgcaUWq+85EOX4vu/rd/lbVNSY
CL/49lQXidEHopeMD88xBddsOmgu+5tSVwUF33h6wUXeONxwNJS/6kIbcXRVixr3JXfiLBWcl/gb
BS3+7Nlk76yr+SGLUgoBbYY8uMpbJaNoW0SNHZBdivOiSX+NWdGnHrVa2UkL6N/Ikj2FVufLFwDI
/S024LNpVyVEaqrykh46pnrZwI95/rqkkdggDauO9NvjAKnOzHdUDfawClvIJ6ttchd4xlzIDFZy
LyVXSkMOWc3NYfpmlHByNJtWjvViXKbcuUvOS1/CtAIffAIXKCCteA8JXrgTJXD1VtCQ/kp0YWdj
IFWijPNkwDTSm29vfDQxSF8hkrgKJvxsBi1yssmPzi2fb1bVUZyyi9LkL/Hf1eyjSzhhrNvJz8/W
+Lk+tFJnasDWV3KUsh459BaheinMyM1Kzy1hyqksZIBQzrF38AwGs5pRCpHmWqvhRsuRW1eRUhq6
xCaPC9BTG0ypJO3cwk9/ZeWmYKrxv/g37HGUriPNeAbRUGkwmKjRL6T6MtVUKa+LHIJ3xZyTnyeA
IqUJcCqgkMePwukAvdzQC1zJDk1Ohk+KWDyhUKamR4vbZy5OkWPbMTZTHUuKMAfArW/Ecc7gSWgb
EV2JltTr5PgPlEb01EeGxtnIPlA0yIBYITzMbdZNWzUHS2RZsfYCu1eX89FLK9deyuLTp32D5gSk
Ztlsx4c4MHW89U6OgLfviVw2fsMAVK04IMhHP3632Q9eG2IcT3lfzVHW4tFLnbSwduGnC0vz9bfL
JxdOHc743FVy8WCTKtTvAASblsdK6GEOyz17k7E6UrTxew5Xc3/29DdEw8+iBuvcWvdNdX/wV8Ru
tP05w+cPW+7/si7ZvRLlXSnUGaUK9r9lohqr8lulDyOefUP4dDKaKBsndW4Jj6Uhweex3//r0WIX
Cx69t2A/xcr9SwFBkTMYxL9+iBvITVD0RkpuCAvBtYvcEkb51zC1OB7dJFjlGwfH7R4AAWDlueG/
ZDA7lBM1jea0v9Tumd6/7ve6XScMU9t1dZ1542C+LRWbDdIaXlfCPjdz/bsAq+y30FsylWzRmLmv
uK7TYNwg2BkZpYI96fajXTYLf1e9uIWphPB/CuXY1arm9Urql2EMSXHsrxEDXUPYTPCss8XYsbMx
aEis0Vk6c5rnhjoNmE7fjedNAEK016RgT1U94y9W6ZnH81kqYP4ovROflXsOtNYv9iBO/po0DyHC
od21R6QOmWz4FVNjKDN+Iag7VY8RNGMmHbtJ/u9dRHmGMhx+c1ifv9A3c5QCNKcCFxXjekFYYjna
/nnDZbz5EKXc5thM2h1V8wdI4S3oK4lzwWMdNLQpjBI1wHRzmxHridH+nYr04IxD6gEGH8hJ1Wel
vQdct+GyA6n29h/Cd4vT3Yma9HqPYK8abyhZnJHUMvilRxggMGF9Wr6j5LXbs2aehzsZNw2NWppK
2b7orK/tAbnj0EBUA2itzLDGz71QXrjXJl9hNceyM6k9JxEFfQ0kETaUX8CptfDV8hXiAWEPJO4i
FQng0eeTbNR80J6OEz/9Jm7PpirEzj8TbtyHaCXJPPtFD8SBltSp+3QJByUkjgwl1tH8ZoX+Gu4m
0Cw4EDZ5lbXHAZNeCdnUSwmzVlR/wKJVV3m3/OOoqRMm0ADpEEgiTkIrzxoTTkq2cFg96KTXOENt
+GLZXLxy7bUz7Qalts3BKVv6GK0lobokhCj5ArYd8072wkLY/xt5YOOcZ2YMuThY3uB48DoDIC6j
n59uo2dbFQki4drY03lnZPiIRyUmjhUkjpMX1UWV/sS7YC0ZH+0ohkczb+r0EX4JFpRxBMgkgHQe
ErNIBYmdLu25/rvSeayldVqV6ZetravmdXo+DsGkFLlbh93W870gfg9Dpd97b0nMTgMjjyubikCf
H3NYvROodt236PqLFlolvYhQH3VmeTNir8y9F3G9/1jmtsqSXc3rjjPmNKaqktDDiqEN5WVZ2409
AIwTQazPQAbT4BbJtsQ89hhSZ64z4wBRD3V37o2lod3YO3Pa6GOzbhczbhhXM9Q7OlVJo8Ok18wW
pP/ycs9jxRRxCxMbKfJqfCwMPFnVgXLEMaIAOvtZDv8C5GJYMyUaxuaUiUadRaNfILnNlwEQ68WJ
eMaX109Vppwj2reCn1WVHWYxc7j7ZqjrIDGPHXHQWQ3GTbucn76gNit/jx9cWTltuubOPYnsv1m5
Fh3wpz7NFeO8fo5DVbkzZ3s120Ho8AsPV2zLTWStUDrOj1mukMxIrW0jUt8YQr3NRNhv3mvrfegQ
iMrV0Kedgf5pSAZV7QlJRGuRPJTwntNDuG+9Vt7j60eyYJUc6hdMbaXL7UbH6FxvsXtYrVejY/kW
z2ebXfOLLqxqGvJ0CSr2U9Wsfg/ZcjOrZNIG7bGWHf9xfzB7JmPkEDCtyOS2V5XvO8B59il+fadF
UVmMvVAyYdgBkndsrlj64Rt4Pfq2zH7ZaR0dYaJ65xdW0Zpciofnjby8IQewm6fTd2HDGr0LF/Ls
CwGGWIYW8XIwOYErhM/ERN8aRClJrOCR14LMkNMgW22FCUph3jtO+gotXfHHLMxFFJDviS5fMI3U
RNuYzBsYt/ct9w/ChUW7xAikYeQCDlT9H/3o0vif924xT/u3djRBJ93PL0L8fVsSMvH9atiVNA9r
DOZ7niIKqljHf+RRgJfCyNoY1TH79vDwsIzOFr0JdekcaUyl/f1Veli4iCWVzfH0l/rzFefp4HAr
T5bonkOEmsb4WT8bA7KLFrhK5pbj3+QNLha5V6LXkRwnxnZXTYC/8UeJyrng5TS/xyiZYNE3I4dQ
IGq1MAg0DmfEUDr6uBWCsgvXB8nKdW1pvMUEczOUmmkcaTB1KBFJ2Q+NWe+6NLNrnk4+XRfhTs6H
FqMBPSlo/AxZBWpG15Z+Xe0doghz4Clhf0cNMNNCwaasTRoGFDhbnDu9MMV/5IkZ2VwJ/sbYWXJg
VKaxlQOJSRxSQGVABxUokhQRJVJ+40+5zk0twlIjfe/jShv6UKSGrNIemQJKQhJGM8DNrXYTnZOu
e+7cE4mX7eW2AY/YNWNqqzbd83DLDnONcbpv287n+hKy7JoOJaF6I0s448pGtubzcJf5ZQ+SAx1+
+BNJ+ctqNq8omqekuVwk+MI7nicV9dxQbrCvgTHvlsB97b74qBfTh+aHhSDN1l7eBYgjKeYhYRCY
8hgk75SkllFL0UGt+Jrl/hg52lEIDUna42BaT0pnh4P1Zs8whIdcFOhAerSxJLKMfzySknwOP6+C
axUd0hkkHhR1bXN8sPfgReutwUzcyi/QWjlmYrGU6VyNSnx2BcQXVi2Y6PUHoo+jw5b/JudrPa4r
mok4mTVhoYZFFaRyUhQCMgT+sozoTU53q7ehbxbssrr9qpIZmxZ9zALmmtLYQzif6at6/xCvM03k
KG3BUkxSIV126LHk2qyeN4kh/FqgR0JcDzw2Qa7aeUGVfWiZ3fWAkG1xjfqNUV/ftFMIfi19YsMR
WSklPvwJlqqEXNxXddmflQE+q8rVCjuym/Gd7NsUV4XTh/K+h1sUe1kknd+Jxk/q3lRzMCZG/f3Y
TY6Ofj0Me9ylSnB/6xF6VAWj8bKBjmogdO4Yn25/B6a9IOJkoMjDB2CWdHDPcoh96Mfemjj1JaXn
L3AhjogFQvnvw7IAbsek9rBQPPsPRmECa+KluZGyBQ3pcQOBGH+IJIIQodKML9ELRAbnZ5BRBYFi
a6aIMJA7EwWY95wwly0xFRbLw3eSPMZfrqFBIjHeAI/aQ9uaPzRTk2s08+PDbV5MqEr1yqLqLlUw
1L7JtNOw4CJiwrevAX7nPr+7LI4EYc7keT5L9g4v572Ex512rJkVQmigK38le8XbWZIQuh3cFvb3
jMRHUo4JAMdSJy1/xp2fwmsOfqYMNnQCHtvsVUzrTHt/loyROltGjJ3eSZjhJdORR41z9cKWO/wb
46DPzVJDWeBOr97gMXl76vgt4mnus1qLTQULJui7g55ToS4R2Lh7saxp9rXZZ0XfJt1/er+/skLE
ZOKJuxAASriUqtfchfrb64pKv6vmg5KnIkXrrGyehiEpJFZoU9sOcL3Viw0FuIgIEHdofWGHMItm
pls1B9g5DWZVISN493NQxi4FswOx5Fv9SLChAgpwk6aj+W+/+HN6O63QEDa/xQXJBA+ptzta+fmN
nlW0g7O49rqgW71LGNScpEEOmLbmKjDxgZRq6WoC15c6neL+aBNZf4RwBIOhiywGdb2fX1PFlln2
FXPuLAWC3wx92Dk8/e6DXumaOoVQg0r2SeW6fInXtYla9glgOXlI9zr8LcB03fqMg9/HjMrtbtge
62HnukGqzisY4s4FEug0/zg2VyM2GiqF9dEpre7++FjYupHW3f0KjSA1yYj2ucZAtkdcfXd6HJjg
MfxdVnm5QJORX/Jl+Cc7Gvb3VTPaPsAEb19a0RPOhzsmYKZ8xnVMp9tE3ieCKUnBWPHpBADBrD/o
3l1c/nTwT1sGmPoRGILKVj08w/fxeFnfUCyl1z7kHcf7eWUCOVoAh709ZsNvNVUpP1pgPHWqa618
mUsdysLG7WTzZG81G5GGK2qtmryI6nUYyyqOXR9qW7N6GvA24df5nbBJlcA0DX6O84P3qNs4MF2D
fv67+QOoFzgbgoTpUbZ076j6dcPEoVPVKiL3fWzenBEu6gnWdxAeuiTN+c+//lJUb/UuJSORFwbI
MMIbxl+YDNVY8guDGAsuq5JwpQWragRVgUkEXik8PiXVqCdbBNX24wIsQZJ5gMn2ySoCMiOUVoOV
frDrm/u+2kqRd4ROsWI1Ry37Hg2iu9f0EQGnecdYzXYggKcLylJtKGUrJRsVjxaqUnkfCT0O9R9T
lTeS5BGjeTwn0QPrlFXFont1CWug9zdqWyu04H9ICB8gw0/mh48waNli8RpEagB5L8Feq2qaC91R
xaIMURdCZufLVmCPVIsnl+gtghxaxMxTP30wS/O67+k/FoN6nGq/oIbNCI5dWFZGuAY3mwyGee5Y
nvn6NTq18DJex2KCGeeTWZGLEHrEy1K87UiFnHiPWLyjGLkwxSYbtkCH/aFIspllMnrF+xEAsaRW
9jGYMezGkwLccvyCsVN48r65z0tTqbXTum+GBxiXP8V7i/7+5HnAJV0kgICEkLOFNtanK0Rt5cSV
972b7dBfNtdsFWJaGTMesY/jMBZVZW9FYyVoom8OWYzzZILskKIjUse2sGvALHIZukXX9irQoj/r
zbNxvEICG47WdJnh/ftxjh4senwyru3mGLUZmC0culEqTmnEAp+7lY/dLvdLAlwZhhAiXjOWjvQC
acS5FLjInB3WTF1FRK18tGdQ7qDFG4qe+/I4GV6Z1iw3OIydFSBBgXl0XPMvkuiuH5IP4OR5s5/s
QGhDU9yge65Ci7sZo82+D2hBodmtvdt7hsEFjs7sFwUDoOvOQKvKh7oiESCazVH3SZDl4peoT9Z3
GedgvRHFeXbbK3SF0YDc9cCwwSnSLAG0JVjE8KaohZGrJy49MgpXQXfB0EmZaY9MLR4hQOupwtSK
I9nSx6SMlEpupB+OWekWltDx1cZYa/vkVzXdHgyNSIMtYDDmOskEp0/ipK9wX90DVo7bnGk4y3LL
i206Z5sH0ykvGXIxkowshrdALNQtWCYwSDf1siCD70g2LYDZo40oCV83A94jJPd+XPv1y1INzOIG
zzEDQk6PybpSDqN4aFy11KF1YtxmjxKqUPzvOGj/ynqUbcaOVhXHsBCLvmJBtQzf9CuDkf9darQN
TffGMOqDS71fZqv5I21g8dTZxnTFPaSYZAa0otgJVryQj2EwFnN1Nt4fvi4FzuTVN1KX6442niJZ
UXvwD0K27dntfGNE6uUGdwFUBmTYf2DzqKxURQNcZcmpUBLyDWSJytWaTgMPRVl9u2bRmdQ65tub
rsV04ryxoa3koBzuaIQVfpHUHqgSTnz6oypTvOjz94wegS26H5VPV7ICLuyD4D2W42O1l+7sarmR
iJC0YWRxiv5B0xPkp/KvTfl5Z55x5+PERuTXAhQHtl7HWe4yhYd8eiKddS4zIPUUSq6otAFjmhE1
Tlg1jNlTkOLYb4GweCpUaMBpL99uO4ZvbtaclE1dZXXodmg+llkMqy9fKdnTd/0rBemA8OjGJqKE
MdscKMJnhqFmI9Hu5vdWV/+PXkE2kdS/NV/ozzBA862EDJm+9CdrgSECLA/ZE/H4sLeRjHbtVGxF
ZvHacGAlO5jGFLORnun0C94GQN/WHaQ3nzTzHKoCjnkqr0rnOLr3+N5jM+CsEa4E0j9PkOZ/62Zs
/Y0FZ/lwv9cXAvl4/i0gnd9NFjyX3rReXbpVX0lrxnEgx6H1BblP26ZRnuTDmGRxBQ6mncuSUdiA
2jCaQPCF39pBEX+uP0TmbTAHe1vKVRkigo++eOSmZdGxNeaPu/B9AthELCCdhx4DcEm02rj7YT16
oKGZXX/RAeZ05/n9cOgUpFD6neu5Emc+ZW87POKE4P78zAZlZCx+p6qOn4qUb3u7f1oA5Etaqmb1
8ySE7N3JAvnjIsp5MVp61D7//yBsxb3KjJTHVpqDB926wP8l2zfGnHM164pOZU1YM+2B6x8UZFVW
11LuZdElHyvrt23IdMoI9uRV6LxotXJbbrrkptsE53JG0sxr4si657ORxhcWe2mGqaXqmDQji1cR
leTdPrTpsVs4pfT+hytY/C43M39swLxE67wY7AKCnRBzIUgqB/3+BPclr4MY4e22zUJFAmagUXtS
luKFFrKI7kDqL6eUiTE09t5FldkkvhINFd3rzuIOBku5vgnAalAZaJGSdFSdf3nqd0gcH8hmnIYX
p0ThbCKoIG0Urh+hp1f0j5BzYfeDwXyf3IsW0cD0rlCuWu2fpZ8C5pEnMkXnQLIbMOeW62yuzsx7
P59rb1xNFMFhODMAiznublW381sxTBD7pxAOQpHxjXrN/GKIkeXq5XiU540moT8EUEwOgUuGBz7Q
cDPLJZKpTmr9ItxrjNFacEDUi6GN9vFE7DWcbnL09DZjJTFAwfYqeo0nzouVCAcrqbKf4JdJsifP
B4WPphWSBEr1dt2O/nHCP3r+3csiki3kqI54eoGjuqQl7XVf4uCOk+qIDOPE+0/5xKsTLfA8KdAk
UK4YqjlOr5x73cekRzJfUuw8OsiF7U1947dlJit6xDsPufJvucwgQI83Tw/oShsYT+UBR57TqaqO
J1kB8U2wWCx7U+IQrZ2e5zC6Oel7OTESihY4LXIKvhtu8WYl07L11DVLnUO/2NM9RoPDzomE3WFl
CQLjiy3ikpfrq3nDeKGajnpQUYUoGe1k0Gxm7ya+Im5XEFQlhcq2I1QnCs9NjRqbKpSaM9hl7HGr
FRL+UJiovp13YFpCIweNClC7ybvf3zQMpUnvHC9qv42JVIMqocRCIWlJnuwyPzjn71pIWSfYjX+f
3kAOxn7cs5SQh91w0qN5gBqedvPHKMFKY/Yo3YlElFGQaVGoCRikrTy0FQMMJHnlJ76OygfxVW3b
GV1jQkZhraof11qysmmVqVkaum6K/E/hMQXQ/Q9cz6Id51bkCp96JhfDPmC0RahUkXWrgZQDG4Wn
zaJy2EfvxoKmgOZSbwajp+3RE8qsZoHcmZzi+s+ZZ8fgiN1hCZq0VE2MScDslcCF2K/kLf81biIY
TVdu8hKLo1xzEwASvbZO/Gg27geP2ySzlDdifGVe7n8i2HNFZA6XoGvB2TV7AmlHqCu8zZSka5YT
g4BR86TUDrhkGrdPSXgkS1Rq/AN8wN0g647vlPq7CywelL/UGU2YAVtRYVijH7e30AAXRA0+rqEZ
hRyJc4SxpG9pO4AHM6JAEvO9V8XrHPdyFgFE9LFUUTOf5tP6rdOHLBJ9FeGkWs2d63Ka6U5a1QoY
rd5MQlZ/BVU78DuGhsZysRV4V73mTszrYIt8wiOC8FuHTRmvDWURd0d7h0xjD1WeoaygHeUSkEbW
fOE70HuR3M6izza+p5Ecsm274Cyvk/6F6IGVwSdCeThyq7EjTVtQnWnlOysPfoOR4MwQCgskjxQP
bMyNpZ3GtXR1wVvfFctqsz4x+Fm9mxGmlZTUA1fY+uq3DpTfOKHvBbCbzmdvLRsgFyeoPpEPEk0c
9c9VaA2riMFfD4y+pvU91CkpNcrXtvpYe+SMBMVBHafMbj3l9TK1pfSmd5f2nkpILL5T/1ax+u9m
Ke/g6wwYcM6twUMxJMPAch9lsc3U+OHU6p+tliGcn7jcBEqZda09ewQcNsUwVpFhfpRSU3Dz/adV
+3V7xmUjjK97U2m9SwO1NMt+3PrnVRMJO4EFHfsAXmtO01RIJ9YmarjdGb6Mpag5SPElVWn+sB1D
9uR4bJB7+JzdxkklTjgk4wBTyStKX8otlE5S6JHs3TVjaSyYUqK6c4tNsQtQBKd63ZtAycGJ3cvr
MC/z+cpOrenzLFsuw9yBYMo2E6cc5GzrzHxabupyabsWU4icL4p5LCHPT85koTgKuKjhxnWj+VbV
XhrSZbDXTmP9523rqSd+RdJnZXoQUQDVjuHSuK2tV5GEP2fL/42c8dog3bi6tbZkgt69Y2CW+YSK
d2W2PTVitIpxjKJfnCu91EFt6M0ZBM0MjcAo4FdIik8xXL/Oe8VroMLihD4gT9ZGyZEXjdCN+L7G
mq2qT5CvmyNFXYCuPRNkk3yMnj9xz+E6qfTS3nisyvZsQZCIcivXS5tSndHTm65Hkhs6f7vJHC9+
NvtfFawYsZ2dMeLxZv4azP9esvSV5OxhuCoyVjnXLaVsLEPzM/qc0o8Fd5hfdV1WskR1akBdLFPV
gxPsc1HAyV7SJIZu4i4z53JHlgNLAeqvTarxZAoHI2Ro6q+irBQSrYRJLuN+q4Tb0Zt+V9X4xOdc
GL4siLk/L+5mLFWPENGt7fpz70f++C2ZB82p513jKvpySJAAEnh15CEJG88UoHKvtxWjPLwt9nfc
7WyUmMNByLqHAOpKGwxtghlq2cVAhp5vJoiinVCQwtow/AQSraOllJEQZnZNf2CnLBIA6NVlNXHM
LXPRZRLj0n96QixYJMjeDXzDwfyES3c/wJQZsYtwSf3df6Z8VgfhSJZQcJMn2hDOyQcbJdKf9SIZ
JMM5h+BkLoDDtw8X8WnwigYuQM7bhdUoCscwJIql/5gqggfi1pndmL8FhhLP2KekxDmrxMgGBOnw
pvB/ws+Jt6HltM8dHbXARQW31ciwk9eDRhZQAQuAGtit5zmW3CRifd7F12480F/jKdn/Kx9Ikz7T
kUT/BwzklMH0RTXrSDWOi0Eqta0V0eYtBVxYPnvctHx9ssC/xiiesZnbVyfhy/cTwr4YIoCvuCCz
dibO7Zy9dV9euzLYKAMDGT7MAEvChJyYTedv8zorexTqrmf6ZkPZUS9E/5gF4gsn+e16hxs+GQn6
J6QoIDRbf1hh3Ww6z4AxZcPISAY6T1WU9fC8LIJmmLUheCRW2RojmsYikT1luG06v/su+6qGWCt7
VrSjI4cQxoBmKsPVUP14WXf3XojUKwsLu3W8UHOt0tyUcwDi0MFNhX9evGnRLnZaAKKeBNS51hXv
M2FAIpfonpLGWxOLKGY4OpuEwdWwzmEtGlxZK0uo62SAHC+L0v8sGxzhOFbu/yG8pDoa0dH5yKrB
Bgws82NQeg8w5yBV+8wLgPS03nIKMIXSCQWJ4lubbyKK031x8eqmzKhLudqKE8B8Pd7oZagtRclS
Eb3vDxsXNDRP8U1gmUr9t4qmRufzC+sdBXUoboIr+fClOIXQzmYR2RDhU5LymDDiS2t3DpGo0foB
fa3VnR5cKKKgDaj8Zd8GVRYcNUd4oBKj5FHoaJRYDzNseqLheIwoUldkdlWKwb/3SNc9+E0dzCz6
9jYWctpf47aV0NF7SxmlOHv+8wrhZyww6LJp8rAFBkTC+abtPD1K4BsTQAXA43TVis35wmUYRH5a
TrRq4VnRjuLqGPqL4Op+BmlBgNLh1Gzxk6ZuGwHggbO3HEripS/FpKGIPHe5eRQFYoDOx0b3lBJ/
EKcbpe6X+G/U1MLDvQUDQhpsbyLGApqZ+AX2NdtvcDO6nkhIQkCO76XEcrX5efLUzmVYvj5A2Ymf
IGh2FeJ+w7aSKY3bW9j6jYYSSOqiXApH9/xF18Ath+YJstw2xc2I7g0l6q5wIIFvhNQwj/kuAxFK
B0NryERqCTDXR3mj0WhpKWDgw9fRwM2RYFI1IcV7+UcBrWa5wriFfA9yIvwxZLCsmrSXd0tZl3Tl
QCezPKXtngaBNsNn3nl+3NoCqlNo18lV7xvw7c6uZS/eBpg3r0rAGdg/UqHzZnS90vQv9qoMK8hh
1NPc00tDCMvoCIF0GR7pr6RIA4W3h0/sTuC0HrFp6V6kB+Zr8koHHN8UZVCPcVZAD9ld+5hfR3Su
zVF2lMbZxnY579oxThOekmN17+7frV26yRNJsQe6pq77H6Re3S7DEbPsPPWxhBRdwmus6YTXoW4y
AI72uvingKYw0wLsXqYAx+CUZ4TwBNMRTqbRqJOIaK6puEJtRT8rSK7QnDaVm6jCGkIbYKvbybuX
r+m5CkWL1ZT2wPQsyrGr9YCba3tAqeupxcV/jWeSD97W0+yqvlkjUmyc51bJcQylaQUyfTUc4xnf
YKr9wQrNDXIK+xOh8F03kmwng95qxhAGuqy4uddLbVoSh0ZSGgINQIe4mNt0iEjbvRZQMCnOsFPP
A2u4aIq14qM1IBmgAtjKFqywaFP6XSaUG50UPk8vPZtlnZaT2t68HDwYMO6HU3C2a41aZhhfTm01
O2SuryySnLyfgN3NqGMy1Bx1FNCkv48qj3+8iuE903OGBi7iPVzyeI3ZcPCgAHo+cw101OVC5Fts
3AyavB0QWbZCnF0OlvAvII0enyBduKEhdduku5Mif14OvM4HN5Jx1Ra0+QBLiricgc4SjGbwpFbc
kLv66L/YpJGyZubdxu3uZe3iq7qUZ6PR4NmBLiYitNg/yLMuz99BTz1TCsI3vF2Y3JO1Uu+Kb7x/
bgt2n4tbPiBqGMKG3qYWBaZE+sj487ztenPqem7x9Gz31WHEqhkBB85tYs2M7s7U6OkIeIycPf2d
Ih+ttV1GsHAPc9kS7yqNHzUmylXKyzmIelPeHGprBUN3P1xHHHw/hJrBoPzTs8nH7GPlZzIsg7u8
lrXwWbHfjrEJ3MUisQNPCDqYh9z4hly+JCnJVsF00jU5jDSncl9PH7XWa+z0Aelhix6EfBrGUBS7
rrof7xMkl1eu8sgWj01xU+OVYFU52xIMzpMPhjJvmgd3Mff6jePW06+fbg/WknPo/tZiEVmwhuW3
kGT9s78lCEevDrfePC1mrNrV8WUP7PE3Eve2frzvOJ8MA0HHLJzW8yAxOAkgph3Z4s+2g36KNMSh
OkJfQ/swykWeZdTytdfpSmlr7p7inxa6XMHYTStUbZ2CySPOfqj24hg7ouE2KufZvxfKExID/jOW
e8kp/IRYFWthJQx+RDG0XFhFtv+zPah9K3aqqTMCJ5uTqNfL+XKHurabkJAmJsAJX/C/JfaZ++4i
MGodnjxpdlm5wBDvZfimUXUUxWb0oOt79dD4gfpI3YvjYJQxxDc9yHLQWu2KWL2En78QuL2M6oTD
4nI70E7SucU4GKJmjFZaVdRy8lFcHlcLZoF1XuHIeLNUQpZVcU8/RpKWUikXCP/mPeQlrmpTIK6r
fuA7pUTrw5btdV4VaxmMOj2pNIwzVaIU2YOWAP5bzREu9SDGzLrImsNvsICw1tIE+f8ddbYwyb9c
9bCTJhLEe7zjJFz9j778XZwshEbILl7Mqq0Iuxul+2Myz06TZmeoI2YT0k+OxqJ/sAyP2CIVZ7n9
vVExLtUSMHnMdM8ZF8zS8SB15W2vfQE4D2cspKXSlCts2cR8o8TzzcvmvrvPI93YWSS9CyzNWRxl
P6CW1fXlzsz9vBuJJYRIAQ7Soy/BTpAEIEP3ZD3VrsC2Jxidy2ibPHEWPgArzc8d7DrP5U2JUGbn
L/wR2K7/ZgmVwdIU/2iD4uxMUhtu1v3EigS6EMnNoXS73PdZGeaNqk1pZ0n5UMjdUGr8KNk4Ms2F
ZRNyoHt+FHf7pOQ+eE56sIuALaKggPSZI2xS19VHCL3FTmYwQierxZGTlLtsMVwQkVywIPVlGfNB
4ewEv9m3wysUxcKOBJMEse5nheakmRhaeHeT1tQmtRb6cvwGeSVW4ZJ4yQf/9/eN/+uEoNuNxNim
Pam5lEoVxIy7Z23Rpo5NJQjBoJZw04iZFFLOUcwIpBjTI48nsvvzzcnPHRs80C2Y89dMhcOR3m8/
cvafs4TdWW8xtJzkdI/3mcT4llPWAOhOu9CEY6JHV8XnMihlCJeVg57OSB1nk26L+KslhZVM9ztG
2fhw0GfLciA9IHNbMmVRGZpQ6RvHPp0wlH2fZ2OHamTFYUvGmQmWhlNVaBS7BVvDUQQjpGjoXM+o
QVMFkWMIk1BIg8atMVPyQ7TCBbfU5n/unm3pdQAzhedo8YbLykOaMeS4ADQXrT3E5ONSly2hXXvM
qL5p3ZN7sAh1Mx9lAnwjEkz3cQKrTxHNqqV/3deOpvCcJM09sM3y19ag2EmfDsoz3QssO71uVhUC
HUWS/d6zHdCN/eu79tpplCKJ0F4BM0Cwl+C7Ssp6+Hr6RtBKsldFnpiZDwvJX/xAr7N5PAYVC9yt
0rYXZPG6zx/eiNktWPXOrMts6C7dx6K/ti1/zUjHc5tfVkNT1cAE9nh8MqBTzrzJm8ohNl8FkwwJ
4lG7BsslUCs/l6Xkt4USKU1HKpe+xi/4S3CBja8xsKXoo4s3IGLE+Bvejpq4dG2J7OyMldVvlgRq
h4TSZ9zKUAJxFGFX9Y3intbU6aG8ZGduz3Q7pMWoDoOwoL7f7Etxyd7IBvWyk79K6F0ixBHjdpBj
41VTTDobe3iY+lsz7aO8x03alhqyINDBge8F2XxE7/2Oj1/EkOgRpxWHdlCe55Nkxb3m55yjaRAi
A5IhLy4CuS2A1ERHMHq/r8Un0LoCxOmtywJxHC+kogTiktK97akD8pOs1zjPRH9gJrcIJv+TUudF
qoWlm4MeWFU2caoqwUxNctJE+pH6Fbjjiv9okqhlHFss8vV8FoR7ni6UqdVCRq/NERPfPgJVJ20B
JsntomEax1ZZpX02dLz/yfzwQELuQYc7NiMBDwbce8rJP6F03Oz3fW3mwUmj+gG1daDJU3prv/bI
GfrwtwHrTF08jhz3CN6imx0sk4X+72of3klhf/zXj+d4II8CupCCcAbz9KGwIYTrUjftIU7M6JtP
9JuWFETJ7tnamUA9mEMxzoqw+Ebggvae3awsUba0EDZ1McvgwOWZD0Ca6inhVxztG4uwHsBDxOXw
c+RLepsw/URSj3RNodicVaay8FrxziWeI1RAQwHVj5MmzOaUuct8bhcDrNIvAkSlL73fpgxBm6jB
JtIOhZ8xZXkzbp8feiM1ZQuGawXek74jjl5PozOFcZXyGOIUCFjOWyY+DiLe/bNXFoFP7Oia/G5C
I6T3rse+UMH5yrL4xASCuMvOVwgs7RT/MC37nQAWYiKOFNyDKam/1Tj1gwPExJo1fHz+dX/H65w7
q7NuH3PMiUOKs4x37DgERYc+s/An0ZY6IFCB4LMuBHGzTdi95Sq4st7LSo3Zp+98QYhqkhuSFc4l
Sx2+zPH0CQo8wC6QOKho245RgjeN8LYEMcYcdb9Yxn2fH6KyEHBr3nkoSr4fgyQKUOegS2fHePhp
QnakDEGomsel/vUdwxOv2pBy1ZPB10L2V7NBTBTjh4cKTjTSK2s31XOqa+idqJ/cF11Df78KGyFa
op7W8JQxSMicZe8/CW2tsBzLD6B761MBw+q7tfJwXxkyxUYrEwC92GkHwKYgGF+mDt3Un0TZRSeC
gWQQ9k5GgaJ4tAim5AQNAQEVZwIoNldx6hqgyj5T2owc70TMHqRLR5qA/l8Xawf4OzUbyqOQf2Fv
Yi5ZtmHbcqDs63tfbhVmzWdSyigQ2Utld5sKoHksR/fpj9yrVIG98ldVHql2Xq23YWQk/TZttqaY
4KGf6pi/QZfhSyPGJxFqmLD0UJnXs+pnKA66r8vgUYe1IYq195wjn7lXpbZZYtBCrp9zkTBEclsh
7+TQknhs40Z+msVeYdZCOpU/1FKB/h2495CBvBDvXw/YqUdQtldqNJp+LVBBVnNnrE1wHc3flVGy
5lV8Hrj/926yr7nuZI1+LOp2sIGJF6is7EpFCp1Noe1wgn4GU/Sp9RsqIA/ebf4ya98nS0M1Pwc1
EvuawRff06MrYcmhtRRpey/35CGlfGXpGb5rEK3L179RsYo5uNuQIKAhMyE7+BG4soyCduUklCQG
kIKcuNnwt/D5ewWu39b5UzZrB6lzxuF8BAIlq9agF3NK6fb+Ulip0ZhPgNSqPosclowKXMhjn6TY
/LlQ5Ygug6S4yNhxcJrogyoohuHgYaeyH9gjGbB0QMQcArSp1BAf30gb+1tcwnoRcY3Sg7FSiXpR
ohtsmv2mm1g+p+1GW+XR9yCEuEJLFF02/4SU3TBT2i20JimpFAVTyAchjW3I4Sy0nt/2vzoK74Fk
grvQTA6FcHK4/vXxtg9gQYD0TYnVTfxKjDbpU+vpVp1hJxW/3noE0z2ruiGFiTxAsxJEcxGxYtFM
wbkGLO+NLzo18WTAP9AgrC7lkqW4QghCLRCuf4QBXd5JFv+VyqG+1LNuzXV+wqCc9ymu3toKHRPI
M08MYljNoUrKzhpeutEqAhUSxMb7Zni9LhkjgOAt72AV6YZOc6DsewJrvzz1x9J3/ezCjHuGuHqc
3Rt4JucBpvXYFoxbHZnt1aSMafUy1vLNNAO5zRHS4+AOpQ6TbVec/n+bFnY77oiqFEaDb5hqMTm5
suhOTjJTlsVm6XSFcJ+XFWkK0tJtLy8ViBACnXG4QdY4KyJ56UvcgajTF+Ikcc5Mg6X2+tawDQxR
gGKFnTa+GNi5Q5AD2vCteppREY31+JPKQN0dKNdpy3l23/s3VnKhih5S82bG7U+t48sfL5iN34WM
oIkxZzrnuLxnsCv66jMAaBEpf9lXzt1LLFlgsANmlZh+tD1rr6o3SsdRSoiwRTgdLD5kzUuarO1R
ubeesigFV0qrQAh6p1PhjYV4buW12E5ocoWKKhojDQ0TmwOYjbBDQ9IpiwgvHW+O0NGO2qyvOHUi
5fyWPbdQWwo7qScWhCS+In1+yT4rLPqU/0WN7d6oheYPnXGEpO/wTH6AkpGyClaE2Fsyyz8zjXf0
vR2qWdZEfcz5Jjn2zXlbbR536kL/EfBQnYMW6yjnuH/HiXpqp0Vh+jc1f18FbLnhff7U2t56K786
mnfhapezfafntA4KVVK4P1Iy/ih4h1eS/Q49BIhfiuB52iU/RWDPFRA+nifWtmd8JPEce021ICsH
PR+wImQX3jKU6BW9Ku4eCGPU9iURoFsdTZdD5DnbJW5KCWunpCcQYmCfJmhSpjY/ITVwXGGIJZAM
4+biBFoWIpvOUB2t+SnWhn9h+zntmAkJA+SxZ2cC8AWZvrMhyI1S/QOxnftjzVppfdb5uMZ9O9Ym
5w79vQ8NfE+suIqIUhFmGrARGgmqNTo7nUHZebxELC+OKlDYjyfAKqIhFWWJhK+KZNu0K5soKSLB
aUagm0UzPc/TR+YG4EbCYjRWvA6EzBg5zbQmt6uzH/w5yldVi+TUDmRR2WzUrVWcSwAMjCtpgrah
uub5r9JaFjz5sSu0LRazBHU7Xz5b+7m+ff6WsKRM4ODq/GP33PvVIQcurl/4Ub+M+ud/uOB1MyUv
oUA79+jlX1d1FIs40Tct1DS6DZyyS1gbi82HQF6nPyHuICIB3h82Ol8p/hSyOA9VjoeNOkCtz1Zw
mMr8juSE6YAZTqfHoRtjtst+M0UJZGA2kgqQ9DS0MDO0KncHHjOr5VtBOKNcOivkVYFwFb+f7Ntg
gBZeFQjvHG4qPZbYAnV/EJ/LpkD62Q7TqWN1DJaQ34OjhByxHeNChQ1vFcSJsRTk32mDJ968zFZF
gZQzdrY97Eonlu/F5VIgG8uE7mYGRAte44MakThr9VAkGIyYPxdsg2f7XG4yN5qgxT48KFeRBhEH
orXH3hO7s8Vkb6SvxzLK8kJLOJYGPrebaSHDjEVXJC6LB8ePQ6a8W2Btfck+ifNpudJ+UlZfmZEB
f+I6GPguxa5GKUmN/C7pP08rPaTCNrtUjm26JFYmverXgVabl+ICywc4jusgaCjffhN5xBszNujp
woAJ+qhq/d0zSbIbQ/wiJ5TB+fOLXJbcv9ZNdhG2Yacq7NZxRylIlIWTP6d7x7fwV7BIBdz87nJ/
ivlGvuqlEz8k4qsoLBM2x+0KluOMH9VDrpiWGx5h1noBsehpWAzHOAqBTFuTXRmNra4OKskV12I9
YNULqCDinnXje+P87rf0P/7k4g7ul+hvxShzYWq+H1LRElKAp/q3KrteyHfGzHTGn0XBf8RUGwi6
hiLd0aWrlct+xIUSk+Ir0pN/FwvnlXjZSGRytNpZ2nNjJ2JKaKt2WIcSkTKI6lQLuKYJUr5nCxkB
oEzJ3s391uGDc6xBCBo0v6CzYnzq47BMPmmBLefK2q+xLucLyMxd4AJC0EBp6gxCEv/MLk7GifxF
vSea+Ovhbbf0zzKvydoHhb2pRiLxznPkW8AE5fK9xe2+qQwswGHZ+1L1glpHtzE4eWr+Z/aZWPBC
jj1fTGbOMsZVeQBfKzg417fDII+l9VP4DCeYcgq7f/sJ1iBLJae7gX1jlKc6kN/jdXThCbOcfWDb
kI00C+mbcMPatKDtQ4O2kl0bwpeYjcKYQZnVoZXE8qAeFCYqeAIW1FR84IbocMBqqexpOQBN7xUx
5L6nMnAQL/r+35q1c/w7xUxd5+GozXsdNnYG7Xcpj2zPFK4QGvZiAF6GOAYiINa3Z5jk6XalqeLI
3o35jaXCq41OG6+vrs+Ph1Kh+xA/08ZUuCegBY4U8gsAfFkwYtni0pYUnucogSWeV7CEHb5sszkc
rGSO4LPkCqjPrP4IbI2tO3nSUZwrW/v9WzuNNU+SxVDBuxj5PkhvLYAH8oceDdTPRy3EkwpiyPB0
DPDhjyCw/2rQKZIkkSQg/r///i0dU3vJZAw0x74b01eFnFqvhG4ApWlRzZNLIxOuqZCnJtA6dm/B
i2znrRU6oZn9f2mIQBel4mMb5SAu1+KzXMCBcfsbnjU/ZHR7gIABao611HjeeeVkK2TFWOoqtKm7
JMfCFs8j6I1smCW8EVKz6eiFjxm4Fy/VjNEpR3T3zNpIWefC+ZwUkkMDQLW36ezOaAW3wBmZCaoO
5KRIuFBqrH3pGTRqbAL2hyADASw5OnSiPGxuX5wl18SnQa9nYQVrY1stAAX5CaAJFIzmR3pnJcMh
yIF3ijvxcjYhbEm+hositlXRI0C/IHA0/Z+g/jOBd8eKKLeIQlg2qiBwh1GuVARs2TF43hHGKkgy
rxyGZ1FhSFsfZsGUlh5NzgNwq58zAjwtddDkKbbT7fdGHNgopXxywiCM9i3MbXYZAe3g2MVMQ7GU
2J+erg2x/dQfo960SmDqDqvr0hgaIM7ZsxX882g+6Pw7gV7psFT/PnCoQI2ATvzGJaZHTUBClKHG
HfGSeKkXGVX/cNPdaPvJJCyImwgXguuYlGDtJ37KSv/aUaxzH5tCneMPyvZxMgsvhn08q8Cg3FSv
xmgtqHYoLRA1NgmmBTsasM6nPI9nvZ+nHuJ7dsOd0ZCdPV2ro+yDMZdyczY37GU9NWRGvPPCWGNP
YxLWBRc+66rEBCP1rR+RWgpwApRFcu93ueW6JxbpJwGwHV97oWIvWm3mBo0I6MGVTZ2oiyJEgcWI
p6zow+Xk02vj5PqaVt5rBT5CFJg+3p3xAx//vmE8uVA4PistiPlBwGQCbd5xr6VxLZeebS1m2Z2l
M2dezDaLIZK2IAJf5uDcMSDzFwhgrxcvr6EvK7f3HMr17+cfn5XkGGO5BMtSHBcQRyOE2BtLa9wO
v/+63wSa1OvFbJZhA7GxzKFVE9lU0RTIHGKLVIsPAs/9vUQeI+VwI7/UIZAykTfcxSJrp0suS6fD
NvOjFCB+Wv0EzHMrGxQk4bzKqB3pjLnvh9pajzLKC4ohnMx2sSm0LC2UghVyerK4HqP1No+/fo+h
O2IxkB0wX6vPGOj9vt/w5GYwS/oLdUpsrq3eGiZ0O7R4cNqvk0wGY40QBwb/02ptSQa146WX9PhP
54a3TJObeN7TKZkgfwUKQ5/SLVddNIo5g7oJpNQnNkvKufmC4usmS4Ln/v5NfDWOdoJ23c1pA0zg
twqdBy+CDLbsAFNyQpCcosYsvhAfZ18nNo/aZ/8Z8Mlgtd6PtlzTOkwdS3llnGZXNT1wsLhM/jRj
JjGAY3Zc0VjhZ1uesye5vbwSsgdOVlBfnqWR1hEqm2CmZ+a57WJLbqKo2n+dfPj6CoCkLLX4CXGT
K3dhlz66QePKugkZ4sXPvs35eWYF8BQeNix9fT/uKOYbv4mqneCfEubwe+HtAKJ9pyo8PWlhAep8
t3bWTQqLYVKuEFr3IxkeqFrqsmhpTPKByiUItw41d1TA/ZkR3uoH3iDAqW77macsK9RWLTDtBzOg
UOm/cmlTlRUsMwovoMngPy6imG8D08xrlds9p55PecQY/nEtnO/x0s727w1D7g6v27DC951u7qfA
9HLIg+wQzHzBBOOI4+9kehZjpRPiiuK7WqoPW77OxNOBj2gKZ9x60UAyagYTvW6Pw0QtC3+ocMR5
zRJvELf89nCfn2rnI4ZVOZ0R/rw2E9bE7XWgu/1xXD/ml3vbqDatLkK5uQ6X5bEb7MAYHfOp9Mod
qgBpj5LDrzScXMu3umWaSW1p9EPsoWnAdxkFqQpdXNwe7g80zS42G2dqh/ODJfmH5rJJFUoNcDLi
b2TsNMBE0d+32ajWUW3MI0sdV4XiAbKtbuoonorkjLiD2gB/pFM5xJHMXPEUh5oPjiJx7bE90FQW
cG0tWUbdy7m2qtslGv8NQ72nNpZF6B7mRj0gqRsvezxkkEg2A35wS6BX8CdkW4ojn0Y5FulhXnxJ
pVz4dRvKtVEkgyIrQNClhGAlyp7uMXk5kii+0pH3pqBWrnWkpzYdWUkAiq0wZtvwnPhtV4/SFuC4
/FvSSu52tBHDESd2EUuqu3sP5I5mRfMiRtVjHqKZN4b87WLnJ/tooyxXpCn5G3GQbY58LXJe2wwK
7m4SZtmAtFjOLh0MTLoGC4y6w5ShSHrbw+a4vUSQCFfkOwoII2oDt8hGvbopYgakuamASx22v+yz
+v1Bwr33GIFMNMl+lG4iCW9q/rQQK7P5yS3Aupk22n7I80AhZVhKeAWdMfkeb3zHBWwudMfXwapL
kCUFjXqQ7nlvx/52lnajGUyWaKyCrooDYM2tw1ZFLpBzSnfAAyqo4BXqs6A5/Joy8WuRxb4Eb3ZC
u/TSpskX2BUKHpe2lxKmOjojrkXeoY5QbGhujkjo1YpVW2Lnbd5de1cUBaERazW8DYwMbPzT5VCS
4kD56J9c1lCqRFaTGAvr9JwqNR9O7NYtIxh/AZZeq2gK4o0FBBjfY+45IcckvTuRNwWJX4EiXDoX
59WoZiZl7oYDLsVl4KRb8FwRk5mPVBS/RwRC8qR1ehovHJXio8xWWqNo5JxytY/fvZa3ndPP45hF
8t8SSu96SyN/M9Zw/VaIqUuCNP2weyykYS/kWS3ZT7kLrv5HWN5mzmLvs4t/5fHGRaN5Y50MBLzK
I0C4ndM5HEMZqdSfZMa/aDBX+W8XcoYojm1eUEL+QNPGSTK713yjH5sdcLbDtnG7khxY5gmKZPd+
FBf7XGMTGctP+2xjcV25fTINWKMKi7bLymZGJWmqoHjDpS8zsRMKXm32wLI5ZHKM6kbbaP/RI83l
0wNfWbd9p5ECGz4Jgud+Uy8ykjADL+R8Czxx4AJ7hFVMGmtLe4enSFbFsrGTC4W5n1F1Tc2/8k5M
4Azp102z+TmZjq21qpxlomaKZnX6D8ok0cX5NtgiDBzvrpxw0bkKdVtlHy1eiZsbZIDCZnGftxsw
IWUuTNNWN2asifHXbvvajreaDWiJewv3fhRwHfrA0un8z76g7jvvj+wRnQQQYJnz3+eCE/3YPO/h
+tvz9OgCYC1uv8HzlmCrKXmfJ95waQB2KfaOenbdVdAz8SXIDkh87MjDIF/g/RD+qmF9BKamrsbA
2fq9hzTsKUVJs0tOdyUFqvLHmoZlzyh0awzrrd6syHMt8vzI7G+zRoR4CKqPH4S21dlU1OqbPa2Z
uekSS900MyUwf0LHTQrD4s+HoZcpXdUk6/zuWx4JM6hoKgbjkNu3XAngQqUac6y0Bi8eaH+vZFz/
58qSSv1kYhZ+aOzqmY3Qan9lNRvnaQJnrCrogsNzEU0hCfGT/+kUpH9GKhZrVcQ/lTLHnto36kuy
QxdzRTGhznBnbAnzdv1HfB6L9+xGa002S591xEOChXUijFnVXuu6pcT1GdJX4jHX6JbhEcNrAVUs
cYvrf+CgbAVlTmA0BVXqrIICkprpLKWaZdekl2PX9BAe6AdMFteoC/KvmRYMpwmIYe2hM0C8vHrW
yZbjpVlqReBalWXTYVYeaD20/IwAp4QSyY1gn6A9vNDkadFNy9SgBNmEZuMtMcIZXY2E7qoBoVUB
HXLCGCWKgT+4SLOfJ06yKLFUYeO2EkOdtkelG9xXiBqZDY+pp+M4UUR085arDqNYuYFFX8lxPzf/
o/6qkOgTR90I3TEh5daU84aT/4j/ogJmFf00jQh3hTh/vQP/mPyH6L5RFLgJHHCDOi7eb1EOnxZa
IiGZvndweZR/g2spuqvlUsG0rT/9HgUfZsJzbBSzy+3/qXMZSrJ/kvwis39QLqJoUCzieGIt3Ckg
6IuN6Fs3uEdTGDOE5YyuDIuhpGi7pWvaDAeoRw2P5Nb00N0bVx6ZGA1FNtMRIAXzP0Ak2mIbCP+r
BAcrFkH1PLqrPFWpKttOJniT+7VyBeGyDkkR18kFA0GqXxsJAfad8aZ8xQVULb+h7f6diJbTV0PJ
FGmNXmTLY5WYBifWbtZoWE7NyOHOuEJGbzcPMUHr3Qz7MjUeFApdznS64zcwcXnebLwSbAimYUth
Pcyw6Qj4cgC5MabsKPRz0q7yamUUPLd5OhXKJGU/gPSD4x1FvVJNxynQ/oXCziraikR87WpD+zbP
8Gr/gLNbVsag3EtzFACEMGpzqsoGEOj9ScBvnq02iJiWlf3VVfXibi1dAz1UZR0VWWd3uC+Qgt4/
8/MFh/68+mdfiLGk7go4wBDhWL4Q91LM0Aqf0ih4tC/YRtoKVCZYpbTxA0+3+o2hop04TrdsatBh
x5yZlGO7alAFlZFPiWX3PlV0CYShx9yvV+PF5rmN6kfgIlWDTBNQ3cOAIoRo05J73lFQAE4mbk1n
Ez5vn64qKE7eeAUM6GCybnwbS8x+t3ga3F+H4Vj04baGmuHyAO7Oq0RQNp4hIIFgACq7FQ2B1S3z
mi20znIbmkJi3taS/5972uZ5Ydc8vEJIWUOLuMJSaa8t1Jgfcvu1SZzRwWxFqyGnuIFzDp/fzY1o
5xVyuuFzEHXYnU/PuvZefEdVIOneugxkY+gouRVFKdFhduvTlHc9tvY69R9NiRAAkDNkoB8U5ggY
RifMpTc/jMJZIDv6wYR5lQv666dITbH6qYEbySJJq2rAEqkjhLy8ti0w1UVgGRXWXYMLOYS70Ibp
I8bqFOfuGh/VayAsaLxI2dFN6YlPLGPdrN3RwD7lCTNH/YBJ7quny8GLwOynI4xVcFHKTZuKipsG
5/qGyVwjq5qNzMbtL11JNo+MHy4zjKO+vl/lfk169iwzWmVSbdCS8V0sSEZYh2cNKME6kAvb/qN3
A/St7d988dX4xBU64aFoorHWszGQosVd91+zSnoCIHxZpeuEMnLx6qcIjryqAVNEy21Gv0NKHKdW
ce2IzmcfUmuPVdeQBqw5pFP1Bc8LQ2dU36AK+a3WM7L/V4cn9otGUxbCz8IHHiL94YDIoaUvkmJv
yyQherWYpE5gGlsASYAjYArlNUJitVxfDgrB+M1wTV3I745vd/0OwOfiUV8R0je9wwq0WsIMzMm0
/lqVTUU9uD2N2la87sJgEDBCFfpHcCsuNI3RjqnYGhimlU3JQOIlftGyqjXmM5KnyB6yByQmnreB
w4ZbYgfckBR5ozc7u2qYbwWSt6wNsYxxvBKV4uqW/SRRIK5m3e8Tk6gtDN13sd/FglqrE35QmmQk
ANNA1xj1FQcCpiFLlHAV+y4yXAjMvu6aqHHwEV6UqU3XttJ8vOickkVxG4cJoqFbMuj8Jbg0NcqR
qvuBPTgZmUNryuut2++MImyRZGPXPTwhBIHo3YB+HzonAJ85czJNPm99+C5LC2K28LlKy6jTVxC7
3dG7Fj/2IcLZYRFxk6er8hfq8Jmx6kv2M7F3LuN06WzwFjNi6fg4LwjTSEc+42LkP3XwkeR90rDZ
xyaHhVZCAtGLLK68vR3AkpzdFHtlpEZJIKNiTf0NVFQtezmv0+6EarQrYcS9lk7hiFnWvHPZi3/X
vP8dkY8Yr3dc2PULxYm6mlBcwxscaJj7o9tSImr33sZHruAsMQE/k2OzKvkgY0oEWYQ6z0qrE7lL
/QJmppD2pV7PcxwBNyEyCycRFBosJXzmb/reG5SKMStsGdEYM4K8nRqYI7ZYiSWjKhyISh5S1kqx
8tv+6bDNZah1NWh7wb0fIRCyRA28RMCmuFXdziiVvFzYK2YjWXTnm59tkY3ZJwVe++a8BuaxL9KT
k9bvWc3FRl5uzEjemmWzfD5BQsvBoHymaEqFcp031NawaYL6CCJfWYVNT+IdLTpllqBQYTlhTpWT
FFYKDg6eXSMQGAF19/ZjRkWKyuVj/pYeGZDS/EhSM2gRIeq08Q5taRqKaQMP/S+CO4QigFK1NX9W
CsqG3I2RujSxtNJAoujncgwBMQ9Q0wl87Rscjcc5Z5cqPs+sJQukGZs9gscYgdFnwywJPCNTB/lR
Yq0C/JIV4VYfTtELrHaNa7dcuWHOcgTfSCoKt+1+UHiPTzNr/K3JPt9AqhIjEoqLlJWZV01DuLmd
Fy1WLP435Q6DK8B0q+FIhn7nY8xFu61grdto0MOJkajiytqzvdUPtbREK7lHjDcd0rynNdWKUvJI
ipbk9Bok7bejFiznFle5lWctwJ4/0ScnllGkJP6DhvdqcxEgqK6EYDlmF9YZggUfjyrR6vCdq4DY
+p4myZrwYtcgi3iwKe0wUWKOjuaKm303SEnrEMA/O1cYUL9JeBGJyjPeUde1+7wsQaeEd7s1m0HN
XLFZ0LzoZvlGKGC3uY+EB74vHlHfUaBdIENvgosu/Re6G/AbqE1DdvUfwgxejvFYRe6VaTJ/Qhq0
B/vZqCtRFfxQRsv6A+wIW+Sv++Z8aLl0ezYmfmKdB6fkMsynPD41+nh74NBAB9VoMP9STXsNNgyr
LWPwANy8F0YEeLGXRNB6Lbsvanq2ZyjDJ2zwVM3eoliIHea1pVfnsxgpPQAboU4TbywVAexTBE2B
Cjdkdr0PuSW+RE9k8kHkc6SogbbzzQkmiVn7gQFI+1qmaX1g72JTWlH2q4+T9ZFdgBrF30yIgZfK
2hgq7o5ClP8jh7VkGlzHcLH5pAfZdni8oxcpe9nXHmFUssiKzXGAN1W44yB1rrPYq9oZaxCEYA2w
NMDC8DkftVC7IO8XK1DJVA7JRaW1srJqQxFadO30NsTF4P870UVKxyJRF62KXewPDKh+spY5a7Ru
/CVMyDTp8JriGIHpghpgb0vcZuLnOTOYRGtJ7xzw8Aef14cB7/9JxJgUAIx+Q59NzzqsFzTRdjL9
FNGLSDi6wUaXemHGkF5hpgTwPmEl3p8HHcgG2/nIEQniDd03PaKqLAQKxYhgUnsjIiIrrNE1P9/8
APAHxH2a1CT9N9xaABWHtwBn8ZP2ELsOgYm2D6OV0CR1Hi86y0W0jSeLoMErN1/1R/CAB4gaNJhi
ZOSMRxUszVkd/NYW4CA8uLoiF+WXl590MOFzfvJ/zVYp5RLNrE8GlffCehHoNODVto2qabaIHqCG
yKeXwpViJTsVRQwqCP0fpY9S9JdnAoynhlfpfPBWbv9B3ZkfqmkE2mHItr6tlq9P75QZFufr2w61
UEyQDdoZWWVl5ZCfT/Pv30c4yAZeQiW0ZAuZ5r/7V8gTFko70MOIZaaDDuFeWkrbGTP63EAhaEoF
ZxKeY3+CLzwk0g2pWzhh0bMw8o9Y7UhsSqEzne/ndqi9ETHvsBE5dj7zjGhhvhuuAmOsEBJVJs7T
zgT84V1PZSGE/gFgaiA5QWzW8O9tM386b5GhoEIs99BJew7Y/UqkXL9+EHtr7R8Wf/rvwa5GX2vl
2bbbl6NCxlmQd2WctLvbM1VT4n3xIhTSrjkjw6cN8XvW5T01dbYpOmdhi7K6cZm/YrBYMkx7xReN
71zq5GTj9MxLH3QtFf5ilnSuKQ4nz4j/T/La39PAp1roaZREA72oLhBCT895fAfwoEk0mvAq8Jgx
ydFyKgo3bPd809rPGq0P/ccKNM+Cm67ynCN1vXmEoHYrTibaDvt2RzeLO5UAoDWMp9VSHKTqv7uz
0rYjPOulLy5LrrG9DfjJ20bq012oa3kYIzn9AI3zGlXhiC91jvljmgXFtqEJlU1DOa7KEhRXQULG
CRUQUjDEq3RsN95APjgDVaJNfEHQm15ukgZaqREEoAwxM7BcZpnLkMPAOC5u60pJvKfZ1JT8wS1G
P7UCSEwXYS2x3/aY9HYmFXnHE7rzfoDf4j9jjY5Kvm/ssipG0mGL4QlU4nSN9qwEmxJLIZWANcHY
/XUkzBF7xiZwxWERYgO8U039zPQOagxXMz+uXKhFrQQGa5H2nAmweA9nD/YehQqLdJAu5FOMvpbY
aElj4pWdbsZYZuNYiIshkSI5GMbC0/njdcLiMDq7fm7WQ1AiqMLhWjx+BBxI3cdA84iLESWtK15S
WkUCHiJdu4f/ff/IKcOaqlUojkDSIytvTWvA7cQIgVTT79owBizIZvE5OZU+Val+DzE92uXGAjPK
xnTPoB2PiKaz+AkmycIbrotEVre2yGrO5dmN8icxsfKJEmwSs9bv925Q3nlXd55IpByRJHDZTxeC
4IpHxVthYsn3G9BTt9JGKhzRZq8SohmB+XH4IcBtpAk1hKVA+xtqA/Tb+C/osApChnRMSLVyvK5B
ahM5gha33vfIJOyCs+G6PEM/M4f0SLCEWJV+JJ0EC+Wt6URr58MD4pyhNKAqygqaIoYMeintdRNT
XLWHq3hAnAg9UjQ2FvJQJ610IdrQ9sJHQGZA00gdHaSRQY5zyGTyIylTRg8Ytsmta2Ewk+kfWcfb
PU22k4dGNGQM425Ze4etPE+xQNA+TOBVJIBSedY61hB1002KZaAwPQ0uPpYs5HxkW+2AaKrvVYzk
EjYE0EhiCi5FOMQDgy0aQHq3jRmXIrQmxp8wDa50+naW88+pCAt+/L9vBbZBKKwsQYnIk5CgPH+t
W0ZIjgfnCA4F2MoXJlZgKF6Dbk8VEGKN/Kmhgw4SSE0qO/DG0lm7dtWEXrV4TdwyE5GDDHxkoTjG
VgJ/cSJLf0++j+tBRnqwdhxMpg+aJhm+E+1/h+OfhIEPqIaPFMK8S1TPnw4NJi14JUn/VTQLVoUF
hkO8AEffShFMsoF20GuvbchPYhaFOqxu9TtZOYrGtjb7QE0l8W5GWM3IuFQdemj5O3MDEv9mg9Ob
aiRIo/A3CRx/v2CAmPDXI8BoR1pB9u7vGPwcAi+dteEeBGocsWuvn+NYXwFs5BmlnDRXoYug7k8C
rk0Mw/m8BQLhELLxj9c2kWEswU6yGJQzez57iN88YjDjP6gjeWCCkbh3tTVzUz2l2rDLxHts0gAh
E6bztUyAxKBow5EIv9Q/dHBhz9Ovr4YNMN3bMT/FxVPaImSzkcdxf78qBsJcEg4a8EX2qQRzt8nL
6u1Scq808YKrg+WQIfoQJvCeexvTmY9mPsZxpsvthXoh37LhynHmnI91w0I8DFcAn4jtC6SFc4QD
yYxwF7UpLKtIUEE9NWvTINXdaqs3Q4u1Cqj1mertZyh/830n91lhwEkJzmLRE7TQMFngM/37hIT7
EnifSyADMILyAO5Z2riK5w8vtZNaXYDTMXfKcgkTlE3TQQczauNO6XdILVRIDdmj8ZzYiFgfWt17
faG1civ9guDyr4ouJ5o1BmDqEbyj82jGEL5lU0DzlJrZUD+9p3AH8JQFU457q+OhHM9I8IZKD/Zr
5FzKluneRglEwVDoa5tOeABQLp7lp3zrBj5+2mnIxLPfZaVgQqcY2truHcmVToazqALI2M4K6/LZ
sxb22roisda4Pd3AvZTiOjRit5kv7bHYhzcmaH9+kSq640ahuXjd+WafzlMTOkpNinwmtqo86LMz
w+AgfPCKtlQTbb3NUZVKbbv9YaBrC0vPPI4iXUmfaltf2oW9hYoeBa7hZ7ld/w3/B2SEdyZkHzE9
poxLo0NcykCMSYNqMCJ+D2VuuxGIAS7UHps512MucNn9V8lTKQXE3pF9m8XVidIzMt6pX3krv3lN
/i7vxsTq9sXdtdmMIhPQ/9BlE1KJ5btk6VBPSicWARty9rl+oqC6UT+GkKazMijSD2b+KebR/+S7
/3UU8/nmV5L+2wgaubIUVMn+JrXq9z6VmhTWOpnBcGDKWMURZGwcp0HKoZ3Q5THEfW5FskoJu3lU
w0ZbL0sGzaJJ7KyM+vws3LAIr2zZuFAaHttn9dnyf6uvhxwUIdgfr6YXARzgAKHNvbkYH2XkCJC5
cysbi/rAcTcl24exDFVcaTJToeSHFN5NKZu/ICFf/TNtj0+No94mGxhV6TygdNn2aYgY2Nwo9gE9
xfofCz58z4YWm8Btx/SFvv/Cjj1U47Di/JBaCAMT5w4369thnKM8VChBtz061ggVf7HYOBM7HUpc
7CVp6i3++Fo0z+suYgjMHp4lC1OOSqRQia8/+VJ901Q65ys1FkTQizYbarLa4hKhsw7gd/AdwKL9
e0zuEoJr/fEdOtHxRzvKfnL0lfJx+gFQ8UR4Yv+tLR8wtFnKlR13whKk6zRpkFXPsKUof/XyyHmM
dv6PLlKTpUsB0F0Yhkjk3rqxdxUJo0hFLtQiVF39tb3wyODWI7s9ubDAgBOIHsO0qEwYYeih6iY/
wO1eRORNCocXdrr49jTqgeecIDZF+N9WBp6PNjR6CwKMWXCMEcyKLX4Y62L2iHQF80HARuJeXCvJ
sZeqsKaJyPgmCdaLl1Kmd0RLPW+H71r5FZrHKsA4mi1fkMDoeuwhtUU6K5TpqU08JidCZ8LY75tT
EY4lgkbV8EgO1z08nHxyt+T459olnm2l/jxymkNbBmh0E4dM9iS93gAHcWwOe7KSemteURNv5bv3
dt8YyJpwrsuJ+wsVdUbbCs0AWonJAaJ94ww6CDluMBwfQC1xmnMhqUci03vAIaU1y1Tt05WdXZFd
I5XZadlF5p/H1hjwT+3TYBH6WUEzzmHCPCJEowGjEX6LMIRYY1PhLdAcFO1Vk0cRHZCjPGXOiGTe
PMQa6+S/jbvmDIgofUu5UbYOJYjD9Xgtk0oQabKciaQuRRPjzUgQOCv7UWyTxhKNwrY7RD9oFnKQ
tkeJ04QasEMqM75US7v21W0fpZEKOvCNUV8BNyIm7/pfrArkhGgBrnqECkTfpL0BXwjo5Rp+Hit3
+ltG83oWqHMMYGFtwteYS7c8gx2XyJxKzWF+P0FirxnsQarnG/atQQn9d+iMEmasKkcq8mVD3TcY
97mkbdSE35izAKV1vuGl/WoBfAL97FGQEI105191ahnK+Xo6667oG2qhs7Hx1/gYAY89i49p8xaJ
ucKopusYY1o2QUtijq2xmzKw8QkP5vNV68zipB2w0xZdRIN/fWLrbFcl0R/efm65I8GOyjmCdLfN
i/j7pxZPa/gSHnO/olmJ4j82hnnZg3rbHBe+lhayrXaS8fvnrUEydLJrowGGmZXvBk8QR5matgvW
kqytnLv7Thz1y9o8bmSCaBzARFV7zTQTRUcjT6SraQIfc7WnnPt3+g7/71KoH+aoDQt1BN7Hppw4
3mVgEu6MjxBsKkz8CQ9acqLCKDj5RQvultikpFJ6jCP/154TgKjSHzCYURfCyb2hxt7YJEFxoeta
SXceF4rXFBnXs2fT7rCBqtejhCqBJ+TolBDYxRVtB5ZADnzu0imRuSatUTJCVdwvBV7LYsPq8Si8
Ylc5xPNpDMaNKP9BxikZYnnE8O+sTB9ympY8XEwyoMKOSx5zmIXlq35NK8NthDlEIBEaheqxpfjb
PnwI5VyX8aS/rfwx38K7b3UbcPk0yMjvpZLlH+hlqGyKiI0bkBS80shoIumhcDaPNAhsPYlhhftf
Qn9MbUd8uD7kDLgTim84R4QL7FXOZPknw6b48DSrs+F4LYDbd9wROOl4eVrCDTDWmwjQrRCpGEts
dMWylY+ajcUvo8xZpUV9zmL6fgQ/lT7COEzCyv5cKR29cMxSUiKlMLXEKGu7VWjvp3sxd1QObsfx
qL2LLBcnfJ+XOm7ZFAaA0m1/5e1ZyK9ZPfReKMoLhi7PfQ02aVei5YVa8f/PTZcoV6fGKNjCif60
9ND5ulYKGc1HMG7EI4ehnfILTJfs16oPi6ZimlWXjTYyKkRm3dhSwIqiWtUru9HizvVTNi0Tac4u
nxsygUyDfJ97ULBhisMKgKepEHiDOWrGSl5GKebhJ46DPG2/hT/a00M9D34WpB+SRyNKjROO/j/z
oZ4FTx90GJD5aW3DLwlEejVuyqXuTjCKyt7clbUHUktClF5hQLyJJP2r71V8pRvO6j1i4OtBfwdt
KsQjhLfa4QId6lnN9w7OOu38U9rgW1Cbvec7JWu8/Nbu8q6J5ub7WGcOsOXkxYIQMny+xrzIiLP+
OX1wXUgL5rdstsWpZCCL+ZFjob+WLYjGY4YbJCLvn8qy7VTZK8qY1wnvNp0jdVCdsrSPSTnmTdIL
gzHRnSHMou1X4ILZdFz7JKXiHrGfEVFIRDVYfum1jFvBCVNF4xzXB9MKc34Mb4vbC6tZP/zRyDyX
TpxqYMgAb8lQA48UoPglcRsAhM8n6v04NxL2daanOAToMPOnz6V9vnij0WDejm/OXbX4dygi2Wi/
PT/8juFwQ+zj3YT7PO2YBwYaiM39LE4fzi8y1dRwB1YqkH/wakq3gioj7foCMOvSSzLreg6V/cCC
ZiluFuwvzkNfHxwYa+pMj8GTJ23LG9XTJdx8A5gLky2v5VssjfSG1o6AZwMooOVFpOp3iJH3sGQ3
o5suK51YNXlIqrAGNnPoiDvd91NYZ+hnuAWDt6D/zHoQiB8B+fxc1NpN5Z4hx3xpIZblI18gFSrH
kiHglvtUCyhb9azjCIc816/IkGnLYsZ7fjHSkGHWMR8dy8wIlj1+8enhTfwbGFQkph2lmaNqbVq1
hBCof5iOUD+bECcHeAp+Fb0DZto7fElDCV/xRodbHZ7oon12i+EWSrLpE345y6ML+byAB4BKZJPx
/6cgueVm05HSJZaEPjf5gm7vwYL0mOfFFteQMVlkOwedHtWl31VkLbKyPpGvcjVqws8uaPe/zP56
XVZanGMoRiIxM/kM7+zYNApj0kI2Gdz5kcRm5zY3ykvpP7KqRKKzHZPqUr8wXwnWipqsAKQpuCY0
iCloK+3OAoFV35UEiuYKZzH8Pte/+VldOVKij3IqvOxPt5QCcolQApoT6auBaX/AQ72xFXCPDU+d
p8TUt6S7+mmTh9Ag8OmHooFt/Y1KwXC3E8Q5hnE4pCCZvcjZAMjv9k8d1h4+ZmBfT7UKCM6ZF2MO
gLC6P7zrSGcKE2FCkbf5WcBETLPA0x19l0hipckXmAVdSJzlB5+PGNUekTE8uuul4GfvV2MEWwCh
UtRF9Ejq5n/ZzfwKqSJyaVolVBdJvqlJLC5DcjvjbXfUkBDrIjmQTASxH3Yqu4PBPy+NIn+ISg2p
q3NnVZ/Iy/4CAum1upm50rG2BWRB/cRTI5RdQTwtK5LUpmlXvtMMn6aZLhjXV5440JRayTV6OlRP
08wYwrEimwxESjK+sr1fV6Wfil5gTfpow21RkVxj+DxdjrO6++FUc7s6lva8+oegKrT7sXCRWbsg
AaatBY51AEZLcwmNZQto0UGeCPJLAYRSXcezbhYXSp8LgvqlLLkDXdctb1bze88g3fmy3JYkaham
uz2nmXFGi2oc0fbZMbs7qhbVj+azJFts+9vMGiEzA+XJ/OQZT9zeKvXpvwTQAOS30mau6qQMMxiG
kBNcqPc1R4hKX2FCpege3ykEvM/qAB6U9ZwHz0VUf4ZzTiG3xDPKHU1yB0aqbL+amJqodO0Wdi6j
yJyL/HHMq0/Dy09/p5jUlmT1hME1fAcRwSkSqvNnwfEmqSM6GdjKQPq2zqcWDxxDbXo5KgqCblai
GK59bAuoGAvJyofwUu4+CVYJQfHiWRwn0HcEzjcabTbugKTIBlgfIjiq4+9NnKdOKLmN/H7a0mtZ
23ycyw8u3HdygHU/3isAdNAswJeMiIUnrC6E2RhnsATbR1ZlXOouTTeZLO1Q2J67K49gQCqL9N1K
O4wrkxyhsxOZ5zOnLTLRkHDrceIQPYHXw2+0DxCSGUUz/XcCJmT/eJuUs0NIeFwK44CHNVtYrAwK
MCSbTlVZymDIbmCccwp4bPgMMpuVJ4pmYYabNKCCHxzOu5byS7IXrUL2d+p96+zgQFNFXRCndusM
00XoqVzNSHlFmJ6A93H0jZ92Zvy4Ph99rCDrzs2zABqRzanQqjLqVkyuHsd+L0blXEvNclyD12Qm
p8WHoYTVkYZgtjhct+gjS41Agzck+9Qe1HXPzImaeH/i1c+K7M/IiyWwMPPp2oGw4r5o9aqKoa10
ae5AWkS8FUS0zb87fl4mGigCSK+vUgtmwKv85H3l70yeLHAQ0MJbighsWLIWNZRkVdfKoEBHxSK4
WH88A3sPzDdhxPBe50gFL76u4vnt5v8cudNM8aeXbZvK+xMp5O4WXrVUVz3xS+aoUhAy5M65wFf8
2k68AXzIDhbvbtWXjTKRoXTpJ6P81NAeMMV3nj1wxHKuVpf4sT0vHe81F5XModPX5oGYj3cVU/Hf
1wRKvpvyPBVrNNxxsF2XWZ3d03RfuTw6NWcnSyxfl5v2diW+GQTeI3iB8j/AwX/Ti+lHx/CC8k60
FcRGsQ8Ve8AmDc0cwTPj5ZQcD1ncZR4awKGC4pqzsDYLi0vnKcz11HeCW4cXeacjMUm8hepfIiaH
33QI4lCs3V62Nadjn6f3wrHqXPBzXqwwOHq3eqmtWbIGGFaemQHikTTsiGG2CLi7B10sUYrIC60S
zkNFDKbbV5rVz16+sd0Opy8nthsS4jGBpgB7dn98VVBntvomhUbXCvBcodsnqYFPIjaM5dK/MtcY
G+jLSYByhLmkcJxEUGpZYjOXWJu2b12UEaR9zMfxF7p4UmV+gp7F0GzpKzNKi+hNg+J/cXjy2ziE
fMvlMzMgwViamxiAV9FtoDcK/IaVQjPnIdHI4DPzOL4CCI0oq1h7QGoB/n2NgHlrEwdQi5ybJLrv
P/L2B0cLO1DUTXOpOEDIy0Gy4rpuK/El4y4jCKQ01hXd8cxVp0CYxuhmylKrPduwJ2YlPWbb2jCm
3WaqinH3OLsqdQotZtjo/Hmnrr8JkE9H0soKonQfU3rns18Bko08kSjIPmfXnctxtNa24wK3s+/D
d+l0Q0M0ddJ24od90Jp336lg8iYoK3cTr+KgRsjE4QoE6U/J4Fx3tv31AcARvAFT3+us/NZfOyn+
8pOej57WT3Bli7flN6buNpXHP1fjSWFsC+tGRP0o7drl+Zh8YXbRkBr4IxQTbOd06vI7cWJvRKD7
Fa8eWfeNCdtawaAROomBH8Lrie0t5WhFt28zeoKodhUBte7NLiY7urh7EvMaeU32LRZ8nnIAOOtD
NRTpKAbJIqDX9ub/LFwkxSiv6kds3HVVnQ7sV7Xj42NO6ftnfMJl4mSLGEG48FCFcn5XGPZSWtwm
qOfAjCgyWqtaTL2OXQlpzBDj98s0v6b61Mk2xTjj8i0r/6jXmaM9xxpGRZTBDhpsIZo2+P6HKgyf
tdZjG0qliYxrPxvE4J1kizMflIbW5V8TR+EIOOMbL9HbXNsQm/DzJiQVhPKnRDL/3JrqW6RDT3OW
K/acS3H85+TuxOWIozbonzzd3sGuzhe45BAOtnPUUPax0Wh05KjDbOaNkfuDehw+rQhDeH045NFx
2oNHz9Lw6cZdnqDjpE1JWOzvR/olTwtrlqHJjDm49ry6Ob8t0C4MagXh85cvUZkhMhsizY6OZtfq
hBsBapyTTAkdvhi6VDtCkaWwf57mFRl8Fru9AmMw8qB+Ub6+KB2NJw3Z5ELNPXqZVglRsacfiiHZ
gSTWpf32pHgPpCcyJD9LInYvynLXOomi/YFPG6JdDM1iNH30qhFbhfeSIW5D8aFwcU/aLyzzZl1Y
IQAGQJHwBMBDsnRikqvlMzHBDWCWN/dfJAcVUDIkqQBSxxbWx5OPVyi1GszhOUTSKn56pgf1+n70
BmlH0PupYVtCnP9rMe/zq6NpoLPKX6SwTp8+5KZu+oMLqGcw2N5ERcndIscQt2hWjFKXq9EZiUiu
82C/bPVSI8j5Ho7a8iRo00eThsFlknW1UoeZIgUwVVSTQAWi94yKJARkrgHrKR1agVbRgp+R0c18
9ogTt6IMApmSGaAemPpZiWmo0QQekktJBKau2WnRbtnjfBf1oEX4Wa3xNfTKgfuyXgxUFQVDuQ8W
/HNE2kX1AN4HVXWfpWTHAF1JsEOM96Fn/cBjxn0lLqLjuaaiZA6uGeXgZic7TqFd+xoYLIv5wtGm
nSI9UZD1lz5Z39Q1vgcWsEIYk1cmXkwLHIfpDKlk5mxoZK2cSObW3aLBgLgsLExltmavlQKeyHTt
/fpYQghUTOLdimGJGix3bzKXefnlzDfnzy2A7Qzj0QWtNn7ePK9G3WZ+7Pc/gDN8uL0I07pt45cf
Iaz5m0FwFsJ3dO/wCzuZVDlgoWNRpOK+25RoBZ0LdQK3D5u+cEEO1N0WID9WtX3bYPxF51sDNXwe
NDNp6fzcRaLX8d2JPvlv5f4mC/jZfKCzQgGGhovBmWcgPcA9g2uJCutH4aDWIZNFgRVsAmV3kUlG
p8MdF3bVQUdBXzlDl9BhelbgYlAT9jXrCpRIvLf+3roM3AebQPAcB4cckVY9YjiDZ7eC2+B2vaNV
29suoFWkPs1KSJXteI+d/bqHsU1MrczZd207em273kYO69lVDESLKiPA3HM2+WFxTnZIzy00273n
TwuWzOLSHdfnoCtf75kd2nhsjjtV3b1E7m9rIwtYyEzGqzUxn2aASIb0FdwrYG0q1CQwh0XIztgi
Cl+Wl66m5wu9SVxBJkW+txblms6YWFCUkK+xyI1AZSKyH/TqapgrSURGyBwyinUqpavXklIUVSMh
Q5TP4VP1BcU3VWmwDovHb4h3I1XuSiGhgD16bULtUJb5hksTFpqPIGyU4lqtVtlGlypByyKtIrGh
pTfh84rTBeP+Z0Q+HOrqSjxnIYIpQHdEMUPPH50WUZU2KpMXplP3b8xDOSeoA3MPvL9dDRY8eHvh
eY7PMANh4BzvFIMrIfK2OArCPqnJTzaeqgtLtn8gePcUYIKIb/jTk5YaT0ccDamaFH54Oh5zqR2t
o1/7HCTntjzizFsZFg0Mr/EhJMEPd5eUjhrcwcCDeoU5S0Oh4OKgM/NN1FIAo8bqnsKuc0p9aOSi
bfIlp3LMFtjg+FYk29mYc4PO2LHVr1d+kY45MMunwFZuG+qgqM9wznNdPygjK8xn82e6PNxFSIP9
nNh9yKZwoElQlG9De+x5AQHb0QkxCXK8n0GVyISKrU2HKzZnqubGK2TcC2eJXHUiNQF5yZs0cKgW
AAr8Bi8Q4pHL3nz8Gei82tFmSj+bPuMV4ha8X8msa/qkBTdAI0LeDzVx5F6PNkj860NLDZwp0m4X
/8BSLimzdTpX4sCUPy9ps+kROkinWOCo1f0LnLyYhO+6Or2hehtUDO3tUSxwvRDVkCuemsZYX6Ck
f3cJ0pVtv0/2VJBUqDKibVIZ3jpmhp41S3OLPOpN9UsJhIXGfn2hAXFpOzxObi6E7gc2mrd8dpAu
OMhHddvvuRrJfcVvby3h0sn/5lFtFLALJBkB8zU0Ndo0A3ahgoKPU7BgWm3kJXO9cSEIe3ctmdLP
yPiFCxnIPHe5tq3HyE9UInGNmmJhUoCiPtKc3J1OLHnu6KEOOrLylmeT9UHhYVZXmE3Q83ynPfp5
NU0S/EyhrHLxcc/brKS8jswmm8NLRdcJqCUEt8NDIASED7EsMuKhVLohVcDgrPwa6FsyDIb50t+N
R/18tYsAckGx0NfHd2IwYLH1U9wBQCl8hBb4mOWq0QNXy4gPy2PbvzEpv/rrZJpbJIqj+DM124rk
dFO2mUqDjaerLZFLKyi8d7Tg/RBodSmyVH12nSELEKMHunEPmh0WggajKdZBNnrGrkBIIb76Inc3
nsXIx/awHF8P52f7f35eUf87nEVxHlHaTdsAnYuvjLfG/96gHBDGDnB5WE9hn1GoT2/Ui/W8Ejcz
3H0OHccxjOp7ZL6WdNv4f0nQ6NXjHCRJZmOo4DfDWjnYR/8ASzQTdc4JedPLsn9di8LyMx7W+t0G
chwZA2HvXlaZEwxp58nH0dPlJLqRFBfB6/fVdCkzxGggFZRzFaom0esedmWgc4BcQwyVQl25ZZMd
qkzzsOh1gyLIUq3VoyhpByZBvchzefcBfcdd9MbRSbL4DxrI4ffA6d9FIQKuKejFn26BEAleKxxD
K9kAW0y4/iXUmkllFNxK4Wygrd8Zm6ShH11IV1WjQMn76NVuKwn2JAPLBZjQ7iIaLsJAasfZgNHQ
sTo8Vnq43/Gxb5mirYYSuknjG6A6XEm6fP7H3oXeoRo5cwSqp0C4/tjj8IPp9btnWAaKh+2WHVZU
EtiX0mip3iSRM+oW41MG6Ac2f4QML4CyKFyn1Fsyp0c3Do5j+y7SKf771ZdyUQtaJ9pCUDxDP8EE
iHBUCtR2P63BldzArIqpS3AGhV121PxuWtDkTN3ReguY54i0j0Xtlpf/wX0+SoU8MQKDrto9iGGp
nizHQhk6VIEwCM0yaVms9vDYKTNqWF6MkT4QUIqRqde+ahSGbt3VmXeb8MTezGhSTybqAbx/WfNz
Ffpw0Ne9DyV4BnlYHNKACCT6yYFQqnv6fv7AEylTzcvidChhwLF/dDt5gfpvBPpV3zt4s3n7RkPa
VU4Qf+1pSKplNG3RspK6rvquJeYmXX+YzSuJrAwCbjAxZ/XDeOi4wnmLm4S9UjDdSNWwXQB6fBRF
x78vLw4NfgdrBuwGmnn5t7XAkUx0zVDF3FZX8P03oc0Hn3nZQLJHrAOvhWwJIcbT6Vs3CiGEul7d
oGEazGOwUbk566qgFoRL4cv+ZG2PxYbDANmalFlqHTG0hE5fcVbYrs+2NjU2BZICy7u/PSmZK0ta
7NzTridQy87qmcWwOQREiKL0IS7+4LSnURzO71OhFws+ediOB9ylSn6Pxxul8PpWc/tspAO1PaFF
fwdNE3tmXcehImRorZuVznKkH49b74XN+JfKuyurstmo1lOI5/OuZJ4oKjb/pd1yd1in0LTifTVO
OrJHaE7oSHBCFT4QhEBzDA4kItfI9fwT8r7QCCpNEZq3JUaeHWt+fWAkClkjkkUCCeS2pdR1CYRw
y28GBKVI/voqDBrTw68yfLVV7FYI9lB1I/ma1I09DocOIr+dRg7ouZZ5Gnlhy/kXap2xoe3Sbl6t
jpyRBDwPAz09cca+/OaNaNnlNjnR/t6mktAj4Oz3GZ5A4riiSjrC5h7GoXpaVNl4m0qpbhwCEkOw
x8ukC0Eter7s+xZNOIKnbzs0mA05GiGXCJ7vnsx+cABrS+6CsQKeLnTuvWsAgxcXf3sQbIOCSS2E
Ba6rPmi4qtSu52rLOfLDwJSjsrXxh7lA9yBumPnwq7vwoahEVNVA7bL7KWQYvvVECOeqNIkfF3tS
rKBFny9v0G68RziQhpugqXjfB+vD54sMqpCo6xQo/Rd+a0xCYLGpBEEs0uzmsQwzfLOPYCVuX4K8
EsomFbJ8npP7TUNB2W1CCRoNxJw/SWD1nLf7RCbP3olDs6HgNb7avS1KVGR8uFPuVSvuuyvJ/gAI
pLosApF1dn8EHjiRZzUP5IY22Fzws1LHcTtv4FkkjELCAYyGHI6R3k6gPnZVMGkCupVSjkx2YVoa
gl/H33UrirZn/g8R8hlfVcYyRyqFXB1rxHSaK53lkTPklYyYRVZPhij083JsvRYC5yBwlyMV/afK
jSvJlX8NZDThpaEUu9fO+B71Y1Reawps009tB0BK2Nm+zlYgMNDz3x3WsyQJciBKSoV6iF1NtY8F
eyDD/RV8VFhDz2CD4O+p8Sbwr07DHfzT7I/XM3pgkCgcwANS9aZlBrUfuy3/M80ldvaDFlEcJ/Qt
sA8EkbKY7cyvRhLTbk3p4CdkP9SItoeeQQiyt2HlU7IXcAfQUSYamlfJVc5t8WGu8kY94so1+762
5+AK0+vjwVjhDVkQbQqhcGRTMP1Y7wrfhDUjHGLCufpf0kdcdQLkq+O5WXvh2jqQL9uociuU+kNm
xayCIoS7L2QcMhqsPlwB1uRxwXfzZT0Dz2rANGQTEqmq2nmA/EAGoz6i5SmV0Z3VyZhEl1WTjhy0
04SZ14IcJ7pUFlGOHYJi/5gJTfA3g5WorYrw17vUNMrUYlCctiKukHMJJcSS41XpxOK13lv7XNHx
xPKmKzi5DAPbOgFXa9xVt/bCaKST1AgnvzEvMnKjUPLAiUeWggW2RiDhEQTPhOEG9ME22ZNhsx5l
PlFQa1I7LGSN6DTbGHATdLEh3ICht2X8RWdEaxCOSe2wuvv2a9rDRh8H5NyO0sERnYwebVoWteJe
wEGxTujsRN0UiuyY+lgG9IyPaE34We4vT6Am8kFMcxkZeCIHwWAn1mlXj25420SGivGUiLQpBSTq
I0PaoOOSsMxa+5nd+XkCtgoxsCTXpQQ9h6Urp1S+BMFVRcXlLMSTp6vZ5Eg+QcIRhTxl1P/DwJpu
VQ9FCDd1zR9EQB2si/kaGp9khlg3JHnJ1UKNNY+7cUaUCWBSX5dl3Lh+gMra/c7VBmOwzl9PkKVr
SrIq+Ml8WfGaGOtQjHpwszG+8HYeKCxvewa04dgb1e6zRi5u2xu4TEC3iM15u0kHvHGqMkDom7SZ
282ePOgbJdpwjxw8OGP0v/UU4vO56z40r307pzSNeXhOaroWT8G4FBs7tY0I03L4dT1Kv3WPGIwv
rboYTXpJH4oE+CsVoRrigXPatO2yb3SiMBSrIbyGB76mui+XXaZ4q8i7dqg3NmhBP2aYIuE7kB+v
A3vG0yrV20fZfIRMIP94M5/hEt3gS6nbNw0CG3Zk8kMFu0NsIKnD2HRM3mgXo3CD52vflGLwgDds
Vcvi5gpLWbvuPjTlsBLKozgWSidiPnjHS+Szwsz/K3Oq7Voeb0zCNdUd3ypT3OAY7AKF2vMEhPX8
FhPypR2jrfU+G/T5iFQ9xzFg2TLiu8th/jWhBYbEzOEUfeJh6fPsCXQyzYBOehdnLcYfkloQiuor
4PH68X7JAaAFu1ze7tAyrrc2WmLO7hq0zqzjHkbc4go/AQ1ua1PWz3YUwnViDqtVMgHzWxvlsHK9
gqwaWSbOxAnJrfdMXn8y9wSCo5PRKnYv7BImfrGMqWMH516sdbogzU/gRrbjdaiga51JibAZj/5E
AulqVZZX5L/+Q5WtFLXwe5VJriRHB1cq7jTOy2l72P9bFePXJpwMEq2kmgIXPKc5Qz/sHmoDzS1i
/ACd1d7bzcEfIYSOkdUQgFDDyUOIsaRuFWLWTly+FACzJAlkEKx5HOGidYN9vqipCbp7n73liLJN
QxwooNedI8J9mlhdTfw4hd+nP1afY+E40w4rFxg8YDhOuIyxkyXOQ1Fd00Y3FMwQwIcMu0HZPrgb
CadVMKGwkSTwejLPys8CKu4rcVfrl0jyRIFxjl8CM0gU7ShL0XgtsVbOwdijxU1a+Q4Oul1M42qJ
2mwmvV7SYDgQIdKLpEOxwUAIX7zH9ChiYIKYZE1hGJcIpbAmUcQpaGJ/tbjFZIXI2JwB/FnLFWGx
HLvizhd4wRudlUFedkBGFAzVQgG8WbgCFf1aeOjeJ7hlXvmNfJWgO53BP/LK1bMRnbjaIQc8LbvA
YlIzT9B5JXd3lr1VfhVhfUXB1WMPEAgCaK21vvPloHn9tkYc/7fkZRUV2Mz5GY/XwosLFVuW4Bpn
sS+mrHw6d6Ak5lcmUT5xxTDOyIUTMs9X61zRLWrcT608GwpQzrTRpZMXudFZxtY88V4jVKcYjv4x
GVk6RiFsPEVlfngn/wtHJl+jhUdQp62S26lyARGDJmwh7aCcivaxz5/+2LewrjpSrHtoh44YApWN
c3MAg3P/5SmeVwb82AF61WxJLJtKwW1TZ/Qj/X6/Yzd2/rPCu47w0fuhAkZY+lcHeA4MSx281pmj
IcJgyviDfB5pBGgWTNJPj0027U61Wv9s9TWO/25n9Sv6kSzwaWTTaAhfHR3jMKyxTUQ//pmfFAQt
G8moGwLM0kxR8D65cPtecQVTgPrt9SrFQzofRcoF+u0KRf75F0fum1QjZLwtpOlHW13ULLfuQI2V
ig2gfQ6w3Lmu0BQQRMMfbuA8RU71UKmU9fxJxzR1EiVh/Z5dJVIpzKP6ymCcTnm4ozl81xTfIeus
D4qmV310mGMkGYB5z8iUGaqCQOeS/KIRtKLlc0xjfY91GdpKlQG3awGn2Y3qax1IQf5kB4la93EC
7S2PCUtOlLad5xtoxM5uwXEizQaqdjcLOD3GhzrbRUSqVvS8Z4Ps2Zdc2geyKNPks3IgEvjtq8SI
rXi0z+FJ7LDmItdbMHxq5u9aptkC5zaJK7C8yxwfPrNjv3oyVmyBNFlMtG+uau7e0hWBbd7enCtM
xEeNPcsFzn9yvkpFCRszK0i3JZ8JBT/Hn748i/DOYZr9dTZPd3N8uyeueQCQkCJJoLsPxjX5IIyR
ngA5LfxfpeCP+Fr5i5KA8T2RRzYcD16YqToB6/obAoV1iwFxNJ8oS9y7uGSk4PTG9jFipFSJVuOl
W3AXOYAdIiA8eIag/jakDiu2M9KGWhhbN8BoO93SjvXwx0cxtW1q4sbwCBRp6GxQgjzO7+pQbY2v
+zj8lCRZQT/5SKD/AcxyBRzCYKO6Dast1hCSiSE+Ak+dx/wiSd86xtFw2jEbD/byztK9ywa3Yge8
NeWluJKIzJLU203kZKwKL0roONV0Opc+2IZRipz0OtrLv20/9BsCGvp0aHZjrFjmxtp903IJV8Ok
MhXn7bJ9rzpgqkUmm/4JjmeomnZLG0tvVWBAu4YXnWGKLqcwXdz5iGNUWosqqouao+f+fHjI06oq
iJGd9yUDCqBXnM+6WYqxvEm7eMi5XTMX5B4dWA75w3QEN3/EHQE75HvCQawMFkaMPEKdIpYeWL5x
Mlew2K48ggSE4KZg/fOQnzF1cvEdUJ2DyW/DPoeo3IETFFrZVhqD/xe/BPu/xTn+V2JFnUEG+208
NMafr2eP95LUDzVwZBWJ8AAjJmN/Qj1xca3gz7/cWHRAXXmL368xWeQ5ZiQvTKTFpVIs+O7J9U0s
zR16vpHA3gq8fIVmebx7ap49N2Yv4fYCSU71Zz+vc9XSFGX4sJEDstg0dodcZvNEkvybogWNJbDE
FH4OETlwDxuAavWY2JTMqVWfcbzBZvuVTdfnUb8eX/OFnDuQjcc1aO6rLFbIB0Efbpi9vIlecTL5
xc71+bNceDaJTrgOiXmvUUK+VkowIc0tkWV7n3AjVt6NnIFYAR42shbG9WQ6KYL1uS8tWa1as4uC
ehS77jwS63LonUs5aM5hLK8XZj4b1XUZwY2jMKupA+yx7OG0JnSHGASjChZ8sICW1wo3IEOGprl3
OcheZ9PyyenAPVsNUfFbqo0GTHk0RQwqHFpV/HwxmrtV7a9zxCmLUyYnSPmiwGQGTmC3Ewdp2rLb
4THXhC1ic7d2vVb1y0wsNfncuPwndInzNc0whDWY+BsXIxYKNdp+EiMfaEvzOJfiNTwlnL25aUOa
kUcjd3DV3WeZm0ihS6qNQ/tp1hJydKzW1dUZQ9kHPPJMpou8N/KSl0XzgdfVLXgi3DZnlbDQhVUD
ZyZHumsy5g1l/1zR5InxDsCI1u2nY0Ah0MN9Wd7+fxuIbCI801N8Nn5r+f4sQeSmJ1W2ppOQyqVi
6plzTcvH56zeJyNryeJKemgGqB9V/OLW8E/PM9S1+4vBn1ab0cVe1ofo6RZciuufjcqz9sO8zGcI
bVfPZ60GNA1eVPa1cKyWsLuwBIZLWz9JR5TNiTy3gr9rG54w9GpIWuRQwReFfZwiRpTitrLMoM9d
tMK3nHYDQVuFL4Tb3pHU8FqGtU6f+X6NFnSr07R2RsQlTTvTvFRTehlS1LNs9jrR4GRADsQj+zdt
jAFrRyVeiJp8/zetRhh1WPoFd4pH11eFDB477OF+JrAAqUlIkk0lRB+xpURqNDi64J597Q+WBx3q
a6aNkOnFc7W6ofWZrpNdAeppfupFLC23gA4Ock8ncijP83+bouIBLt7+G7YDE7YhqcKVh7y+IHL2
uougl8B97WTsYk33dv3F4RHRuCasweh98QM0B659mDhwL4ER8WXxLL8RVR/dPUGWutJU6vW1/fbj
dTtgOa6QGwgBaxZbuZgq6tU7JrRGShZlsTm9TxyO7auU+Maeu7uavFH/Y0r0DXSwp10jOevxH176
91t8fa+BQV875KRkxIQSnYzsZ0p2OD11E5WrX9LqWXUO4iTEmLSDCUvNKgRh3zniO9HMiMw/97uc
3/f4eazFd7T6BVNuxJ+0s7xghKv3hYVAP8S+Jg9kp5ns7/eOPTC8oVhLWCY5pN+7K283UhMm+2FF
ic8kE6zHSHOEtCs5TTSyQv2/GsvZvwAyl9zcRa7tedZnvQBJgC6aOkz64woH/3WQK56Tn9zaplEO
pxL2o+ophAB+zgRcsiIQtfGmY3BVse1ZIZTa1mGYzlL1WEEhbWiVtRCIgGWjbkWzxR5uhpJ3hglU
IyaaOYx3qcFpG0neXzymUFrn35IBxX28xHUhlf+4voZHZG4SeV/iQJtCj0JrlGybXhixSJ+91REc
K9DNvZUGouGKqsxE41WEXpBgBzdXwXq1SgPdgmtCgcZjds4qjzJzN+yBHxaQqX+Gd9TmeNksad6S
KOHYORc7Wlaf5nIKwyLgpMWq2klgLKvI4oNyFJuWNiqQzoOTl6wLRiGra5LaaW6z+pthUl1V0oqp
GDp5yFUkhQpWf3+7cJ+Jm8bjxQa8YjuA2i/+rTY6OAJhdGvCsY1nUPHo+OMXz6JB8FRW7hHXST1Q
LnVwkFBOaqly8jbBPp4VkK7vnj1qIbeTGJXSbD2BLdtLabT+OHrlh1AxCpqDXoyTcpXoJ6xvK69E
KCHEEdQAIck+hkErzDUzNvanfoqJ6YSucx6htm9U4zq+bg9AdpZ/TyamP7mVNcHuGz5010rWd3xr
zXg8mTDny9DcojzHpAwvhGK89HQ6ehXE6vv3iLxcWUngOp/K05wbZsQC3qthJPar1hJOpYsYotNm
0G2QWYnHPI3glGXYo3ikLQisb8Uo7L4Rf8sY4jz9Qx//n1lcoyvc4mBAPzOrxTAiHgf1EJ8v+Q7/
Ysi0osg3RQSCaYOGCeKoLqqu1uNdOnLZ+ybFWMbW7fhHvj2qH6IoGqQoizo13v560EGLbvbZ9lhm
0JQmpmA6e1hSi0eJnxJsZ4g1re0dSwcJ7uEdNW8EE2bgcD1hED0wM35FEGcjd4SS4wNzLmXK2IyJ
4GLYVkBNvE4e7WQA2zZHOy58IBVy7Ay0gwzoRuFssZB1QLP+9ooLFL1e93Po7Zm2J+wTmcE/KirW
ryhbkuZtTFpTJwwdcUAc8t4sp1kbbu51/LwLNeWO18tq+V49+YmEcn1sk0chUa8sb/WSuqP3xQLg
rrroC/gANmq/lB6xKgK4vSkbE5eLqY7XbxBLgch6bL40G+6BfpeQken7y+l96vRq/JtpF/14397z
e1qQUXGThzL/9nGrh+a2lXFALsNVOWkJhIOgmKapt9t5+tpLX2lKbjgFCs19sjuIp55Y4hD42i+1
jXQIIaErVuOh8jQ4RgLEiCz2H3vpJgyKfeD3wb3UFfGZNBEtDmVyazD7rlE/hw8N5pQEMN1vv4m2
VJrMpAwyLIDBVABJTWVz2Dhl7UlwPzz1RmQd9YDzCjFR0RkDXzV/3Z//Ha0nNi/uDyP7YnS9s127
eE2tem3Jom56HMot4J/Qpi9r2UlWWgkp0xOOiMvsaud5vSDN21c0StX2ec6XmW0DZMeJY89pvMNV
FDGeMpAroNKKYodkhM/1iT1KFqdTrd5dfPiAtvQkLfjs3lEpipcdPKhicRcJfiqh0vQQ8L45Wvi0
XYsKVGENIUC1rVVco2qt9LsTJOviTzScHXhyy4KhR+tv1ggv8HoKP0xZ3A/+RJv1TiVZk4zgFdBW
7GyLAJuoMI6xc5bsKQisJsMO0hq58V+PIyr7uC5UaG4MgGumoeCFY8fkt8rvSO6fDcwEXizMyvvH
wKgfdN663pceEokV43st3mukxTrWDuVkNBpQV9Zrc1wJbSyu6e6fHnkZi5nK9eoi0vedIEejAQfO
90B8AYcYHdZqIXb6JwGbZfJs5Tvf8PRFEm8dA7dJpZCnufDp1kpHKIrwSNvTjA9m0dC8YbKPwOgF
3zml0OuGcGJ9KPUYLLxAkFoOkcT2I5aTFqChnFVwRnYqWxuQaNpvSCfEbTqw+9vJaYKHimOtrS/y
i0M3jxIK0W9MIk1iWn9brJUsSfnAIMc5IEfSWBociTG6YZ4erhDvJCfdiGIY6X2vOO3eHD/zjxYg
6dA9GbIqCanNurNc0zommcVIyJFf8mKa+yKeogNQFQhsU0TEswV8pLMQX9ah8oKiec/BOaffZFCf
1BawNzZ9DIbLWpQr9bEpXeSDgCNKp8nTq4QJA/RvGc4YcBLc52yJYpw82ga1WokigR5l9nfoUNgI
K20cjLsdMtxZW8r2Ls/+aajBq+5htMHgcSW22xzYK43Vj54tOaPl7KI34Z13rYJAJV6t0ovbsAgA
BEUHQtJmqBPqpbOicMKgjiZAiGOXfUYqaw2jHVrPmcM7P6qo8uPq8Kd9iO/20vhySA7MGGHxOCYN
k66l/HoO5KSucoCU9k5QpLLdi9rAqazBC7THZOI439RzlgdRE/O/2L7zGAOROKZyG7Id3G7ynoU3
RIeBVq45nUSvB5lS8GNtmxojiiLULuXM8sD2sQ0Gu++HIJhWjAG4OW6HhDx5XT6lF3LQJhaVmMCt
Q7Th6n22VvVfe88yk3h/I8DRo4Evi2eAfwP6Mt0eHVkQ0rWILQ3GZ6S2tM+/XLw+xkQwBj44p3mT
RW57VtGo8cDwrcXcdDJzHgUtQF5YOM61+McZyE2UNKsX71jcBA7Nf4f1lv4ltZxo6Qt0VGkXDrPU
YdA7iJvYfIGMcNypo+Z7xKBMXwnvq7C85/v9zuD+vfKWSuhpFT9nhwJgJUWASxgiIqyOazA+dirp
T1K5ko9DfLeIRr6/tEmttWYuIJDjPsc9ddk7IlM8DtYINPgcdfR/3WL3YrHEJiQkzi5xQj6IaUw1
YNn4vrFY5beAR/XdTIPWw/mibLmqHuOx+ACHTCHG9evx4ninQD/u6VMt64fhqzpatWuW2x8SrOTR
vyemkSxnq8HneDrWzl4uCulpCPOJoVi8RvqjM7wHQ+ZC2nzkA+uxPF5bscT/+K64f352QzeyWW6Z
iGg+YgG5J5klYz2aRVOJClnGt1G5IdUOVRxGVXuf5X6RQlWprXgiBIlN1VLs807YJgyZltImHrxK
MZq+yIoNaPVqHU7YoksnqvODnFu0T5iMujC8biVxuoNW4YM7VOCjvwI5GeuY1oUq/YGpVauudRwH
HtZE4AW/hYmG5hxj1ZSPDWFMps2YWkr/0V/qo5tGk4GKM7rOWt3o82sclu4Qel3z7uEPh0aJ/tw6
frtwZ5CQCgNdVxL/Gk8amPZ8bLWuDiqUqaxDpjBMQqObm/ZDKf0wq8U5L4/+kFk/gK50LPKOzRHU
eSaX0I6Yal45oey6elFFcnMe20Dn23nI/wUqD53/BPzp1AmNw2i4OXmszEDCvcyWhVqgj3aVFTxy
OkBblxiZEzmTViRFPPfFP5RmbSLaXZ59ht4ZFyYhYponj/NiibGySIC9txFQTe/H2J7pIq16HGlh
yHvTcr4Smm6x6If4hCsKGat3UmG6JN+bPoQenJlq+8tMb7bcJnpFzAaNth/QfyD/eTjnzu0omfqn
DsVBzI1OUl6pnPPw+EhFA/5dJBYE6v/7PXrBsf3NzN0bsyzAhHDYhHZs5kxp3Qz+YdlDWztkL57H
4eOX1bhiJFXYtXrqRgrrKPZ5+UQqtTEkb5leqgSH75A7GAjTOaGowvLcy+ClKPn6xxfc5wXFOpUB
neQgN9rGclCbGKCgWZ1VATQWTnp/RTfE1sPKKGAjqe8/g8KOTII4J+XgI8Yj5fZAa2oFWSWQzONC
pyUa9zPYqA+eE0v2jkrGfOtW7X2u2N1SZCDyhdQYtoJSLiRzOirmtq5155fbNDiP7dgkLEntr7fM
457+oZxUVOy0ysQImUd7qGan+aO6bT8CcHFuKmntxWgebXkgpNyyv+S7YeZ+snOiQy2dVKuAmUHA
8Ztm7iYUyxMTSzee+i+rBPg3M7bUtvFNeZJKy/kVAp7LfatmLDHilMG1g/E4y7d9rsGrhFRcdGBe
jYosWk9BfqPNrcl204Go4Ky1UWLMyX3r8LZWoI6Y/pQx++VEEPirXIbeHO3STy4QAO3ZRHRS4fZm
QFMCYNVsXtL2rm5Cq/o07ACbReWo5dVN7L4dnlvLScWkAMByU67G1JIHok+BzdyHxaiT+9x8XDtM
31WPBLY9djE7kdu/Sgv87JhPa/S5bphzzOSIWIiiMo21ceIp6a1EawUEsNsOuEhxUqVMa+EuLaFJ
it3/Iq2XQ2913UxG69UXVH5Mekh5R/cdIVBI+exXEy4F/jLjbwbh1VFJHJgxYpPfiwBALed6L3iQ
RTL61NjODjneSQ6f4p9QN4hz+mrfOmD+OyvBjlmYT5w27mQR+0LFpx/FKet8aZt6GyzoI39Oih2X
ZkR1om1CqX9tm7zTGEKWjAf0Hp5unVXTX63JoIQvri3LpXbJlrs8jmLo67pfxuPF7pWJp4TW5DgW
/B3AqDsUKSGo4RoqMuOeU21uCFFMdtkYGwCRTaoWVEVmLoaoqkak+doXyzi/CC2YBqgLsYky8dH3
jN0ncis6g8Q07pet5zSkqRwYiP1W5/m9BxyFV0YHxPZUuvUk8Et+Y0aZpyDev9YmzTt00p8PaABw
SnmreR3sWEZYjBMkHyjiEM21Fj+GbbifPytf7twYa1x+ySR2yhS2L6dP0VmhWaE1lF8pziTingRA
w47qqAPkMRGvv42Qqya4/dD3Wkvjc7PVtlINVqd3wmBHFirHzSIDkY7pJQNVAoBw6xftidilCS9X
frNwU+AQ/zzph71D6YLFsh7+CNl1lCY2Y01Z1JjkACWL6H2UOerQRS3zQJwvpZe/gKC8RQvWKF6g
JzpT6GxVvp+vyrdxwqdqKlwrZAcMPLlk56Ygiial5ncVnWiVxt6LLH9KGesmukMn271fqfdDeB6k
pblBt6IMREWtAKA2plO86/GsH7pcje9RMce+jnousCL2hTRjD0O593lhTfC8sWdjYUfJ+ubGuStE
wCz6AiTWyIackxnK3Hy5wMgusyrdw1bJ3e6VNQOxLzAXCvB8yQEUKFxIac+1gmYMniJo0Mxy8ynq
PWKKWmjVllYZOPyxRKNffTMFVcD8F2ORrpeTYZUnwtSZO9m3ZRZl5RPJ1CTFClKkxe0Owj0NkmFi
MPY7If3YC9uLujaGNKQsTdzGX+lH9zJD6tvWHs+gs+hrvkVxwUMSUjQVkoQEjFQUNC024H9OmmA/
JvijBG7dbXkDNbqqwKgWJP2U1nvY7qlEBJ7Cf+AQiZSTZeBAHyH/tBTNf4S01PL3RxjFtFChf9u1
DShh9k4+zEP9z/IZ8fopyCVvcvxUl5WhI/LPVtm9FrhZocCV2oM/ZAv/S27J2EB4ejdQwMDukasl
37xJkM8/Bnrscga+TsVA6pXPj8WaMbGVFS5N9NabimjGJwiOy8hxXWGt2L/oYgzC+D7fkp5/qmZA
OP0HKY/aFKNqm3bVqVatALkVIFzhVIGeNvgHxZqG1FTrl3aF5FA9nASp9iwIP86Ik3j08LMGx7yY
mbUZh5m0wvDinVhNvJ4HqZNsGHuIRrZDNFom8jTrVQzGP4cvciQ8UWOB2qBuZ7uOMUTSLrjgnVC/
VGjSdYbYu9Gq6pkECspzYH4On2/wC/FfVzRZzvWPLb9h+AQDlxYev0blM1o8FX8/257aTItl/6vl
HFPx6v4NKbqIeU7n8q1ZW78DsPbAaY+jHObm+IFIejALSPJukcNHEMOjjO0hJzDibKj7N88crbeP
KQXlwbC2jMIIwQrTM3Y1CssiZF7wFKmYEVo/WtVLjukVl5GOe/CMdR5dFRy1VUPH5gM6dt0ev0Lg
VpCOT04ggxn/JKOfI7GSV74894OkXS6bLpQnBSpjmEWDSp++bzlj7I7sI8zCblLpgRIW6KR2+Z47
OZvWbUwW92WNGyFEtd1fubKtRF8WytjOym8rhtFX7d3oIVVn5OL+Gzd/Ark+opQD9ymuJSDKevUO
3b1dMo6gtbnOwlZ7if8Q3QiaO8l6i2Kw3zsTcK4i+WW62p6LpqB4GkwcZSAMLb5d9UFd3hriXpoz
I681r78rhH8oBoMxoI7nrWr9p6YdSckmgu00kxsuPoGjccKYs+Wbnd38c3MPxZlVBhRcdYIgls89
+MbJiIqPcMPd36IMrVBFkG3kUyJQ3deMGuvRglRLKS250UOkl4r7jdHIocaRIGFw6eXlpOdfsGFv
zWM5ne/Gwuv9m78od99Jg4aK7wpf3SsynKrLdHgxyPUXr2dNdPgykuMTirJrga4wxbyZQmgy7MME
6D4Knomf3zeOPg38UKyOx0B24tco75WqnsxIalCr3E8jEzWkMwalen6BdEDnOoWxCq9mLvGOw7/O
yr0tJFsp1WbC7jTcb/uiYMRZP7WDgjGM8w97r9E3LwtNokE4sVm1QEmLAUzBNSY0CHtjhvf/corh
KFH7wtLev2S/dcW1x6N+sVoCSu2AZS9ny9CTutVdGR3fRvsyWuJb9xEKYyju5I1JsP1uaISIwxD5
OcXNTXwdkUYmMVF9i4M7ou158M+hadMX+eAU2of2uRYviN45Dt/AuurPUHlMmXAGKZFhra2joR0m
KS/E+R7j3kt7YFshxWkTIw8dRTF2j+e2z6Y5vnCxm1EONvISg275cO1xYempv268+zURWh8wMgs8
0yinxQkfuCgG3w+Vda40c9G1Ze6knA+FEqwDRGza8kQRL7y47OgG8tXtt3wfygxrWybl3eIaTPqg
0A1ZZYJO03uIKXtr8lqv/Y1HzJhw93wrjOLNHbCtx5zIQrYsv3zDOb060zbgaPdz0+LdEXT0NTDY
JNctFntGNPEZLE4stMRbiNlhRVCXa9an8/QdqI8ylTM8huogcNmPc9T/N96+LX9pm/6pkanRKog0
WX0meXv/7jhtXwEfjchTey8tUnQ/orLEmt54SgD7L8e3kWJVcCdecMEDpWXJNaMD5/5V9wOy3QDb
1tz44gbnXNiFNa+9XA8Jmgvx7NKnBm88pFAI6NFLkiM8GehohsR6pZAzKhBGjJ2O2sw4hBfalZZo
mplVIMisy4Iv7OVpkBtH1HuKwTrCkqIeBGxA3zHbt19qP+1vE96ooVTeZCj7buOywO3r2HPCqyER
/yoEyincaVPLg0jtf+uRhOBQlyBDt6dc1CrHolOZtUPnVrPyVkGfG51aigfMz/8eyPVwhOSNaGaf
9Kbhz6jfF84SBSCJyWYvAO9sMI5RQ7r/zMwqOnrjrLQrJNThrs+qYlZSCJdoP+hD6/3tZfobzUNa
8tJ8NLSLcgi0mGHTY6tZfveYHmfeM787jOyvIq8Jp3w9fXGa817SgJH2B+DS1LfDzTIe9Z5FuUP5
d2wlN7IRj95iDisoBbwSn0TaxY7X8Ikgm0QiyTvuip7QiEqx9muyeNy5f8xFXuXRGf36lu7Rrnsw
YmZWX96mg08+koP1/W/fuSYmRf0dGKkQ8NextyOLkizpIAOtkldmqSGDNTsqb1UgkveQyfjg0Lf9
9NqoBqxFWyfcDMJeT9o6nTKmqA0FPSz9UBkl+Wr7gbVk5n6e6TwTsAWZUs12NWJkm8OBaax/ie2Z
AvknPJ7QWcDezfY4Gmyep79GRyhr7zsEd4wiQI20ndTxV6B0suiXmGfE/fcdxbyWdMN57RpDAW1n
2tzu2GYToBtIfwsk1LJKCHsAVk1hF7IrhRVqZvNpnubuUBtqR8c6Lv0SBND0aFC6o+F1WLCjGxhD
aV7hziE+InE+cAU/Pm+F1446dbuahzAq4q1iFpLjc7LyfPlLm8nIscHLWEIemx1XDrhfVDEdrTbY
/WIgQGo13QT1Bzvkw63griOIRdJDyq6F9dCnUyjM6yzQDGkNnPi6Ha5f0E/l66muHubk+gI5S8IJ
r8lK1yX+epYT+gO2CPAoEs+XEmlFQgOEVZbJDz5V4tHj7LSuWwhCMbFpQZsxddxWd/3bCHCvMWfp
fyvXq8V30hBfkU5mYp0GHx70L5TdzsOqHpJ+G0rrXRf2bv5cUDdQrVSjQMHsy16xZ9RijOUwotqv
DrMCu00es7oiwTYV73VNhvixCfF+9IKKjZt6zo8x9zIjGD05xUlYjAWJ3xlb2jQUtqfdcDm13hzR
zia+atc2RvZVgfwFkG4W4bfAa+dIbFRE2meIsYExRVsuty0EVpcCSKVZOhCr9Pt4oPb2nZJrjHu5
wqKACiCwzoofbepuDhvh0/SPkwHX6sC2VhR2CfpNEp6TjvAZ73W40OEGEl2FynhCWM4eNvt4dwd3
c706rEVoVbW4BgCTxL9boIoMh0GrVY7d5vRd6C1HqXPqFf/c6z2wTv8k51UGbUA5bD4JCGd5q0pq
29uQyMUZ/ZmFBlJEZm/e6SSLCg1aox9lac1opMw5jNMCnNkBOjZ8/TzvB4AT4uPI0+K+V4J/feoj
mPXWljTyITh4F8rUx/w3qEMTGIQqvR6HzV3v62Z9WkiU81fagKpnejonjP+RmxNC37s6N2cp9QcQ
hOwsF3WMt6VK2ETfXr1nnp9EGyTv9wqaDugRaLhAXKE+uN0LSCibc35A669vVyBSvSf4NjGeHGVg
vKDTzHDrkp7PwCAWJ1pxW7/v9X77hPWcpXE2IPO3HvBHK17pCQThIU9X4sG0Rwpy1qzgWwRbOiAf
RHA+WCRtxJ2vjrqY9NvA26PfCtrGBmPI7Ny+pK0GTKyttqJA+Bux6DcXAg4Q0npB0NvBGP8GY0It
3YGGejdN8zpqMPGZlfGZaNtM9nQd3OXC2pxstvSXKiQkpMlOMPfjIJGX9gM+7j3DL0SBg7mVLX9i
X+APVIMaMBWri4xWMpiCllMQ1DO+aw8a6h1W85LORjFc+UcAwKocXJ05J/JiCkowj3LJ5irHOLss
EJSMBSP+7PHK2lo00/GMcmCRXp/8yvMfH2P6cbEdVmuULqpHnlpOM6NK6u+H98pYX1k3XghHCzq1
uBef8a9s8T1vD8mhlYZ0NUYPMbl4ygPikR/GBDcdpJZoz0o4YfIn1VFJ1bzXXvp0WSsFM1RtL7Yg
o0rrI/GMZ92tJBzQlV1yHQqR5nZv53gx0Gp+IcINOV9R73o83a4dTLqY9XlHVHCJjKLy0ELzTJIU
lCm6StnLe+Pz8KXQjzhstIL8ZC6fBqTShbl2zvq9tS3KJ7xzjZ3pgy+nltCNCKXbyT8BzDn/KG1C
3GhVtMyyBC5G5J2LtP/aoDlrQcPE8hTB8FGOO/U+cssk1WgrnLJmL4s9oVckc+/iw0hu3OJWZjpX
jpiyKln3EUwwEB3Mi4idgiqomSsD8DbN3K9bfYt6Iodym3WJKPe33w8N0Lpxxe4TdWjiDylcbMKr
3Iey5wO+j2TGrgLvKrsXlYcZzqt1ifwnu9U64EspKYVYMQfGwc7gOlXhJXV+LRxL5/FC9LOVbAf6
yXWIg8nih2Ikho6zeChSh5aKwYWFqOIdHa/9xjYTitjfXhOYvlDlEVBP7YyySl82dWNEXE593pwX
eAKCKXEH1/K3YljIs8fSCJxLbjaT63+NbvDZ0OVmELYG5QUdR6r5Q7V6a+TQHLZUEmKXed4MpI2R
12m1TNZEsFYXZt+TUVf0Ob4IZmpS5UPBw5MdEf011TYYLuKjGUUT8SpVkkwCtKfo77fnyUuosCCy
/0Lm5kJ0xgUwOo44IS8cI+sar92CMJrQo467NN1XRhuENuFBazBteI7EGOlJnm3IbEaHMBj9nFJh
dltCeYzJ2QySB1gCC0SHShoriG7jfPXn9nMV1sTK7XzlEI4HG9oBwO6wIoxT1NonydLojTuGT5T/
oYvMlUlycfODQmtEU8HBFSXEgX7lrVico+59/pFroGKaEc0KG3EhXx5k69i1UN3vUmniaNPuWFMf
Duu78z5EvqUTkq4qKewYVF0Hx0kH8jpKpqljJw4RFOMuWbtP4gghaJX2WvmJx8YbDZglhzINQE38
U8Iaay9Ep+UfmFgk+d6jxgLF74yJoQJRHJfwStOht+RIL2uIrdf7w6F7ayCik7HPJ/s+w78oXMW6
xLtE8E8mJ1vpwb+ysgrEFuz1lSVXxzv+ic0eL46n+1IFG0Zy0ht7IKH64Mp8XdYVRgSDLrCsPcl3
PFtIuJ8/yZyn21cYpCi1rkmFUkNQEgkU4LecpKEOsRqLzlqKnVjjdvqIKBvURudYmQ7Bz3yq03tn
BUStnWx1tluXoOJCEM6t2Rla7HLdYQyFswgqbonOuc9lp5+AsCLeAPBIoA/LjmZtPPxJY2ROg1rO
eQ300NxbpGX0kiiyGCKwbMMRG7Hpqv1vrP4dILUfhqGRPpF9BO0n5JejUM92HPsDi/IW8X/Cm74Y
6/5D7k23qofM/nqqj/4p9rBY4vHi8E+L10YCpC28t9J5IpFsYPRRidd9xgIHO0BL89sA+C0w7Tm3
Gdtimoah9/eucMUDBe5bRXRB3qU2X0TvHJnrGntyDyWFrnooNrVCFPpF/l7kLHlTAOy7qoXdSQDe
5Bmav7ymzrLjn0NStI4tth22nSu+0HAa0NGWPBTPBATiZ4/ECHb3Sn9vbxp/wiB60HH0+ip0VF7m
R9nODdwpXzlyArtl6FNpb3E0l8W+90megtaoUXnRhmswMk5r/9Uhkw2VDqcc8Cb8XAsiLEOvACnH
FuxsL2uRd4UtUgkWw7jgTge6vkHVurt+wll1TFrp0kqer9piLortnd1XVM3NtuTbG58SXyf8xs9M
Yg0RUBPMntZAsDHtaNTIWoLPoEllEax06cFIlGpAoujiSsAAlJ08rUhbtS8ELBtYCDx9xSi6pyPd
bj69zVej250b1D0rOr2Gse+ZwsFLR/YyWxIvTMP7L0LpZQk1qLv0sK/hIGwMk1kzVw2O1GHYMD9f
m7GX8SxRGJm/cPo3OQtahRQo4Ja98i4U3QH9q1okdjY5hFfzrdPqI5s4Y0jhERQl6CktNM865PGe
AWZG2o8yylwBxlyzhxOtIym5oSzu38s5YTqhUGE+o1Hof55Q1nsouI8dikTpTPclZSfMnEdSf4M4
0M90J+nynhHjVp1L0CyFM5GGRdMKawj7NSuPNTEECRDd8CXx5DJrPZh2mlkSnVK0Cr1TnyKA3t3v
d3o9+I0QbCswS8jZ86EfjHNE3nYHFGvJx16pDTb8C+XhDkEYBXmb6lrKdVy/Xg3/ycXpWVt65ZYi
8Q9OdwVyFdGUvcfOrfYzkhf53/8PmpwyiP8mZdZOCLseAUkbuKoBdAVN4HmcotOoW/y/6PXhYMr2
15NZ1JYkdaqaxlJ0OKdD+qNgBZDwpstZWfEqzu65TuwW3B7kNY+j2fTuS8mdNlyb0jqV4VspmBRL
hZp0mu+NmRQXoCO0rBhWRBpTWBIGWgpF5pSrSAZszjZ6Z8xV4tzRYADfQp3PfyjUEFmfQNeQjtKX
6v7SF+SxD6C+ElRuWj8iIFptY/k8lxKUWWw94IcazbxLyUwf82tNVZmn+95Z/gkaEd58aZg0n8pM
NsRNtg/j3jcr4jdI9JxrWCBQXPV9fvvfaEo8Xqhib649b6vn3TUCGDFnezA4U9e2kCKw8I+jDcQe
HoYEnViWHUOQCROnQp0JCwD7iJw+Z4xHO8o29JRviZ3hFRv0A/52CvAq1Es9yt+4aGwU0HjN5nmx
QSrd8gUYLps/HP4OPYAOcw5eA2A45ZCeeMGc4qMFyhT0N8dRMy10bswykEQcW8hCAs3wj0B16Ylb
o8kPZ2hY46b2L1s2OCBFkDV6ZWSidVxvF9Ux4ASOcBMxKh8nJ0lkL374K/n3miu4mSQKqVWkR+KL
UjdYLuX6YOhrdW/lw5FZPGD+KKCvbKxWZfjH6NFVPBEZiVCW4G+Gdf7CaT75zJxiF92KAqfh271G
5HCfx25tF4uXqAhL0KOagcX1ACJclyCZv7ovvn7HLGFi8x7usOysFU6GXBGIg3ZFT3TBna/pL/kA
rwKfQk/F0BZUvs1smYocbbvmBJUPRZAOOclIp47/fVKZ9e/cHqdXW0vvLiRHTH3r7dQjz7U/gB6x
GNpiKnQuxMTp0QhjJ6Hx/wV3WZNEad5LvPSEG3La4pOt9S03D3aIDiDHtMBxnwWfmbdAFmAbDGXa
T/kMAqnKYjN3rv3xBNIagcLwfcai0cUpfeWAtv5zGgKTd9jiJ201WFbkxzVMjFw4iKVMYv0Q5LlI
yqBofRsZaKh2dNYd8uQdY6biaDnBeCcfepqTFLRzt5we8q98iRT5LuTyUI/SNP6U/VLvCfZ28MKv
+ppdFAnA3y/ipS+7VH36HQU3KoNxNiTiRaWI6KPPv3DoPf/hCQC7F98z45KfsFUCq0vfFpR7XG27
dlj4496hA2+PXVjZEWI9fYKLEN+2fPhS3FsK+KVXV7JXuWjwwesHbHEW7YaVyQDwrXxQMepBaIGs
6OI5+TjDZQb2WsH+XSyF8MuExAcvh/g+Gls5UIfziqOpM20xOY5nW5G4Te32ZhaP5+jQ6NqwpM4k
YyiWsbuP5QF2dvgGErUix2yXGYbPZ9XTQlFK+0zzkdsDJneCjy77i65Jo/fvF926G+D2qpgg581Z
44KqmugA9XqzuI7cX+vvmTLDp9/JjHPJ6oX6BvVDAyK8To3a1Ea64LOqUGNJvIcN4cEarGKzLPu2
q6QRUkkrVbkOJIOfZEFky4HXXsftViJz4KqdlIGDNRAZObACdWu6vlwnJA7JOCzphncna5CL/Vo1
/HUxrFDXqUZjTW1fwAzeIaMlmk9ULzpoufOi9lMWhTuIUshr21wJDrHbNKIDyt0uwoJ2oiGv3xM/
oBrkL2+n6mF3AQzhs+K2haOFQcP0El6hGm+aKiLpVjQgOrxo1H2KrOt/OYLcP70spAytWygui3Yl
u87TftDu9Br8bP6O7ZD4FZ3eDuqM7BdLe5lUsNaTo6ZYf8QdUmaKDDbBtoa6+0OFdVmHlQoV8Lfb
aUL7cIdc8ddPtnZsF6ccuhMhpqWNtXUnKUSvCeGKHrpD8NQbIWlfbL+CIN0nvcs47RFb/7lOaKXI
KbVrXhPLC1RUlm2ZmC2ThttHYGpbwRMFC/barP2zQ2SaRpF+yimbaZZaI2o7XlQncFjhyatAf8H8
2ZfAb0s7zfU7lOY8jaEPtFKKow86bfV7Bc6RveLCXoDuidzkZ5SpAE4vGkq/baY1CS267UGP8FXP
/82jpAHcSzPzL0QmbRkQcLh5BxmAV1PXv5cyNEsizq69nMyJFIe1BqPw4eU7HliaT54tcHru2jmF
UJTV0j6O2p6Y51sFLkVWMkLT3GMnajUAR8vTivlWKl5C5yTa0yzBX4ynXaiJhXktdXOmAEVNXFG6
rT7KI+gidfRyx62v2JoTB7ErOEggVNJqVSPSQ8lPGtYGkcEevGsqtRd17ec2EZ6TeI2KkDqchzc8
3FZwE6mCre19f2/Rf5iv1fEZzo4s4yPKycH1oBo66mSEaghaXcMZT9H4awqLt9xczD906Lkpv333
d1BZZkAzQ9nIpz3hz1nNvo/heeAxe5HwsBwr2J98A1gFF8/hFdy2LUTrFlbotuDZdLgWt+aisfmv
aW4YicZPXPsVYNq4GJNFKjbNKyNVZgvlkODkdhbRBQbXKZ90AfW/IRPCBduSxnERgdKeHi6J0Nja
+SOWIa4lGTqz82WoM4YHysU+6qzm84z2TNB0Rgeq2X0CDCV/jpvoPFBa2p2tntHxoxWt3JtmVXpe
4Boexce9MSz1o3pXdURUUeeMZKBw+6Iss5xtjKZzou/u+P2XynFCYbqxN+is5inV2+XRf+xqLos8
923OxI/DKAG65uatYhMFR3h9aufAKD+o9z+WeCS6WO8l8GsAhWpb9TB6Y0bZYTutHxAz0i9YSf1Q
Nx/ZQ77lj4cQgEyMnpQBKjU+jGRs31mqbs/gzqT/s3hd/bf2XNq2CgimU0/CH+Q0Fbjkyb3Viz1R
Cg8sJjAv4Rly7W84ZutJintiPk0XdzjF8yGjr8KxGci6bBawPzCMYdQUsaBixhpEh0/WKvq2N9VA
MiUNq9TL/LoshbxAqdLPnnTio9/rE3S0QB4n26YZGSkYW3xNe5qpBjYtPDO1wZfx2ZFOAZyYrcgf
g2+5tHvI6ezs77REKZ7k8MKXLjNqTlSwOhDl9B/VniebRk6rmy54tBXaK43G2wxWE+O1Dv/XLr/5
dVzviOawoY4GDWWhPOIn079eTty8ibyndZdrelhNZhRp+t5Cayg7XkDUdIDNUWiocNdxWMiHeEVA
dHIUvTGK3vfs66yNC+mw0+szPQ+mv3Ivaf+xWJkS1gpX1wX0oQtJoHokhTvcol6ZxlubF1fwaSPb
mtQ/CfoMRTTosNEzGzKK5yMiDlwNA4nlWbrRN9dbmyEbZHMPmsd5NbRq3DP2gLI8l+V3XDpTcDlg
Mb4kJKcKeFN/h2ggHnmS0AjMFqJR4hAN7QErLoXRgurXVbOySoGzVAALLzbLB+N7HpE0kJazUmyw
V5w4saLNX3fnZzp724P4RRSfkmzprBGPEJR14mh5HVHzUFROt9BqKGpf/kQIbG+ANZJEnSMsOGWv
9O1fVBpix/1L3rrQiBv0T+2CZCSmuCfaTmEKewDxNMl1U11SfGYhni50PNp9oqQT7p1uWwHfQ+x5
7Ewa4DiCWoezVkPsaYGMYEDTFTIkM9t8VBIo1sEUaKFJBovL9Mbd+FTm8FaY3U88EL7reSgjqKbv
XWeQ42Jv1vI5G9zrSoL4JEgqkeziBRWtEBCodNlX3Symf5B/JVi5r76i2jgNboOR+oMWYqPs2nyI
LW6errFi0pqnyB5DOpoCD8fg0APf8QacZZrTwutMASxCvvKpirEVABwMdz8K7cpvuAz//vUg9qyq
lHW69kjNhM/tL5XSbPLg/2M/BUyIvfIqDRh0EYuTnNygZPLG70bbFhPjhPmFDrZLrad/UC59Td+b
EQWpKXdxZmnoY3c+D33ZSok+VqixG1rQz4j3tooXnZaBmwZo1Cqgt/DWgEaLC3LDU641DYAleUyf
ms6tEsq+pBL5t5nR0J3IFBbBcMWBVi0HLV4BUnbeLaTWpR7F0IfUgt5JT6rs9egQNzjzLRDon6AK
hGvT100Zt+QWjTykOroKcUN3psUlNlxf+/je2YQWOQcSzdr+nhcoj546n3mX60jtn5WnuamsK0ab
IF9XdunWEMipoIhbIq/vShFkeKi8VVAE5HiSDI4kMxayqak6fctbEkwqFN19x+DyRDqWf0fE2bje
M9amVlGQ2hWLWJLAH745eVXS06HxSJzZ841supt8RPi55kABBysDCb1plG8lfUj/FBxXLYjda/wv
MwQEMXUKWMtbuhX9EYX+DN1BRnLx4oTOCfmABiwL31hFI3KacQ65ezGfSMTNG21dCZBR/aYCdIZA
jOIr6tea8vJ6PBLJZeOuBI071K3PyH44z/pLCS3DjpBfdEyzilVBZHLiX7KAjt3UquxBkN9U4KUG
zx3445Wc5tZ/By0Rc942sYsiNWe/4HTL4+IbtppX05uTFSAapRVOCFaKoo/gEWzvVGYZsBm0ZWN8
jZdcmA+eUzUZ52Vu0MjPB5FWm/OQ2OQA1zECsWUcLLGTLTj8iUkhj82HuhhyH+L7YMztX93Env62
ACOJ1ARLa1/K5UqBDwAfBC4ozyHOFEqjdRO3CoiUHo0FhCHNvwb6Sq3/G04YHfNMsBF7iXHUpw+z
OUfLTM8EqBZjswtlWSA++ewESxWRj0xmhDt1HjA+q0BI40wCGvvN7bpO168R3SI5FUL/jrKGu1QD
0lRr33NBjzoxrE2kFaWpc91seHk4rN0blnP+qjj7mo5R3JScF5I4LUex+JFAP9BstGUC4yRL8cSh
E6eLgCRakJxBYKJx1GUkyPqt45pr9e5EPJC3QdDv66wLjBsaapWNfYHJHPUlUH1pfauivf16VUXf
hPqBEtXB4ly9KkwTRhG+9iMru9WoioTV/eDDV/zqjVV4JcIVN07uleU04A6hCTM2J3LHtQVRdEdG
5d/6jRwOb0/KjwUlH1wKHDnZ5dsqYe5Slq78jOwfvwMPiPBGZdBfHaddPKg08xIbahYwR94dvZyp
qmcNO/nWcVnQWnPo05GyrMmyA8TSG2i82EuI651hk2cH1zvArONJNrsaEjQwO2WT77PjGIhJ4p0y
2n0xFIkZaQ/q5ZjSbF2R4F0hDW15A6UfsatWFAxmpm6nrNJrTpJ5IKdRMvJS+hjF8SX3LDHWZ/NJ
mmm+re1Jz0+T3xek+UwVtqe6dci8XaTzRi0+KdpCFKRf2+VLCKiDs/dOz7VfjH10tk4OcAoOl+KG
jjRQ2YEezY/3NP+lZk8ZltQxiWPErbi71RQ0XkYnUeVVLmYhN6IeVTWWeignNOp/jYvO9CK1Hmbk
fbj3R7rFijJIDoVnf3S2bobM3CR0hXkMCdwFrWHhPPr0T8yK+zOpMp69X98VGx+AAX3EXgh7zf6Y
oJlgFczTfL1AdlhZc5fJLx9kideb7IIBbl3xFLobzCovR7mEWfJ5rB+x6LVzb8+Z8WtmOJC552ey
7pYv/xWtVtzRplMXJ3SLT9OJr+jvrQ9NsnsOTYBUiutg18YUDhPaGArrmvfxMVBYKHcESfAUl9EJ
h5+QUFt5/O3PzvxseQlzAW0KGprAAlLxB94OB1haKZxM3nDtj4p23HzDcBQ6mxdSXUZK/9hjXdPi
eh5DBeXLB5FAi+LGb2WkMc1LxTgoSImCen8pF9IvuDLU0dR9iZWklKzE74o0mgS4oFwcn/QbQz9f
RiTJVFcu8chXmeVtVz9vpkqG7aNdJtm7/H5Ac2RoSMxkYdnxoAfPI54nvVRDYblVT3M8yS/JMsPT
azK0IiWqfRIyFDZUv/z91wK9cjvGGhX8yY7K/SscaH9/P9rAwTYRXrqmah5mwBZ+lul31MdIt0xx
9AO+Hng1daCVlzSIeLZeC5iqAEGHPl0L49VlETOz1sxkVIi70xvvDbthpdnrXgtM3MRGTCGAttZd
RaW8DQnHRAIDq27y/9TAu3SExAU5Qrsv8UtHCbmYMFB/QYFoYerV8RT9gP6cB0SpD/nyNAbmilmE
6Nov+Z8ujIS1YgYDXYLUMuVKM9TEEJ5mVpOqKjwoV+4/xUgaN1QC+emTxfq3UH5oLEOXufli6kd9
Pxv7Jh1TpNk0lR+VkJC6uGBZKjZuyn/dJ06BCscH2+h22p/asgF5azqi+D+O/ZC2L7dWaiI8IyXe
z3k1RxRgOeZBVMbE6iaTLSbWOjseA9LH5LwpMxEGWViF3hm8OIF6m8+n2WAbZOfNb/MJ0hqlu1zw
olls/mrCWXyhfudE2Z2deDhStO2eKHs4UrHynadcI+CmS9oRQsKJwC5CXnfts+xVbvagM6rCI9Lz
EDUCmoQ4JWqExRYyeiM7dM+Ats5cR9UkcsRm//OmuKuOV3PkfABgiy2tJdoToBdqSISFvnHZQv6/
X0kPjevPB2hK1nysJnG0XnadUYjY7/tirV9gztAFUPNYvVVOYXY1lx2ryrXEV8HJ+B9Jl6eKUJM5
zTCDGEoMHuXyQhlVP8ivFnfoPy86Nexbbwe6yOOLyJ6FiES83RfBJg8EZGHPfLJUfvOtLISlFTBs
PpPrwHJ4p5dXJEjkEAgePhL2tGsWRbJoxVJ9E31ywlamrSHB3zP76g25wjKGYP3C3lZDz+ZQROf/
F85+qd/mQIZ/NW/niYnrfE+qDl2HuK0Kv7+54ReMsqllnekrK3VMHHN3e6wZmnD2bxOEHTNpP6Kr
+EAB8LaSWXydXeGODYdxxmYYrQBE/0gcP8FOLu3WIPgwQpCE8lZW/84K/9bU+Yss2QeetNsQrnho
kQ0L1EXiqjkHt7IxN0XCdQ2hXojjKwCpskaz/LJnUHGooZRd1M4LehIeAIQ/RZlc8WSTqFohf6VT
bBKzo5wvB8J8gtZLIZIzDy1I7WvN30k7fH4SRWRFgwRpmDrZLIOUbJWwNBrI3PE4a8J8/zE2gHaB
gqwSofySKI3n4ebkovQK3pWsU18ZqN5S/fQA8sgRXbdMs7YjE/SdrEkNAzLo7lzfVtpSi4gSbkA7
A2mlwAzQgiZvTqRAYONCYkEoibY//QZ9n5GZ38zEkV7x49XrND2tza7zFecvH32tIu8FnnsiHOdG
DVqA8uid9ckSzg2FbusIU/TG5nPk7myONuyGWlnuZ8DN/HO+Xiu5t7EJOywCbbmbJvF+pyiAW8CN
RidcZQgViuKSpYF5E1MDb6w9CDU0MXG7tdoOsXRCLbYMfdEZdv+ABzvgZJwpK6FSc8DG/WwIVqee
QkWiNawvem+UIkGqOLcLOgG42MSDYHTvCw285oGKCusKOkaIk7h48VR4/TP33abUJgefgAn98EiH
K0ZeBFUd6QclNgx4AE47jxisSVTr226u/2ugYlFr+Z/d4SoBrdXHy61GIgcupwUPYwnRhuUq2eNl
argn9okcv0f2u78FAuOflY0zmuLk33Qa5Qlin+zcS0+BGCjqRKiLQEC2mIkL1iQvnP28AdtoL1kl
ZDqJVAuk/DNEbsBsKCXQKs4ACW/gaL94uafRnFD2FQTp5NgvNax9viP1Xq9JyFdgG2sbRMCyiMzV
H7cd6n749Bz92bMO/9DQOH2ZJcgyAn39rx2ralk3gjkyPzwY4SufFRO2N8/vXR4+YNHMkOE8ICsr
LEz5IGLu68XQnAxCB3iIQe2ZOyWc09QsQdsKn03tM8h9Ji1IhNAIG7WgMkFPB3++cblPAjY69JRb
KoLzARsgjycctwl3y7Kj9iwPXCsstNdUVEYLfaLtIs9YuRDkIQYNO4xgdVgZWvSpmSqn4cPcMMOy
BJatelv8iYpObNk/ry7+Qg08v6KcPeq5tCtubjO4EYnBwvf3/pg2WTdz2n/mrvuzloPda/TekEz1
+jm9r36PUqI55uTsudJZuYCmGf5aRGudNOwsER2UT29GO9A7o2n80e5j9p4FV4wLVvKWR9eUwxBZ
RVAC6DFiqTOFTSZ1A7BsGTsLVwkRkMskyurUpUrfVdqomWmG5ap5/8ZtrvxOIwhfXu0nmJ0f4JNL
5oWtJn/aOUyJLybxp8aeB1+EmGuPDkmfA9msd/FqA525KlWBgD04AZ3+VZQ59xP8+VsVAlfcztGq
RPuH7tHfKh3eRHpR6D4YFAszp0L7IUXZ4s8fQ9bb7YF8tenK/d0I2U9VNR3JXM/T7aTL7Rf9fr/J
3uVCtQ1dbuNcgkcO0GVID5nHRYaJVQjBZlrWDRvHYkj2BB33ni+KzjmB4bQBzzqM5gSz80m9lG2Q
UHeS9Ridd28302AMbDSnmU9rrl6feXmNNoej/IQkaZ1P/M8qiDghToGop1p4ygn4oDuNf5w7V1JV
7L7sxUMaZ05aJvFV1pLOzNZy7cdW493EGCCl+x0bLd0rKWK86kQAOOw9fijRZjQqb/2A5KjZ7Xzh
PDKTEumIq9Dn+0+iURR9DxaE65pad/LJ/RmLjvVegyUiwKtRmSo2gVivhEJarnpDZeK7HnU4637V
kbJ/5Xg9Rb221XdT0f0gTu5oqP17+6evByKfSmFrtg3Tb4M22S27vvHilFYVasioQxZxHg/HjZ9G
/ztRQ42V6OHkBuP4wEDnJJ8RDrAHzOnH8gYcUrD93JbUD0xnugluLhYPTPx7ZKe6Z89DhzERvcY0
6OX2nK+UDrAX3t/WaDelyL2jsD91qmffc6gqwFYYR7csri/R/Y/VaeEndly6qOYO+I4UiopAMLhY
pNh/L4Rg+btoVL9Bo9Y0iOe2B7ResC6cZpxxs1grm4ffF5GQ9BMVQUGi/WBVGFOMr6ODvP/Inm03
nqB5j9p2lhI3XFrUyrGehkyxlUXSR7JKArdDYzz70pm3KvccaiDmlpuWHliz+TcnoyFVU87QTJCV
LDHU/NDFbjnGzelx9HVnksH3h+u5a0u5h0Vb2mpCRrkO4BtcG/FXZqsv5vvcEKryMamI6vucfxol
ol1DE2LMiMZNmrPCi4ibmWTYgekeyMdSDxwtcarez0rY3WU9+T5qGQdwy9cjN4ZvwHCSAVuJGVBz
SXNgftb2mi2on6sVwG2NhTuU26KKmWk5pccX2VszsCDoyG8lWJuTzfzc5nOsm7OlIRpPOGCPRJj2
rR52MwH6npeA5zDRcfeo92xZtDuhhzw4XdQB+VLZnw/tktrR6b/1wT3NgLT3SZdpHw3iDmlkBywM
72d7W5fTz6CTjJkFrXJK6jIHxHe/c0roDN1kNiDpwEePJZWCx794Dh37cFPR5Cwf0fJp8QgA13zU
mLBUpUOrBgcsF/SW5h76qu1gF7wl4qNDKNA6KkhJAXC0VHAVOj7a7NTqc2hgpm8Vgz7r6zqzFRpj
+8Qki5pMkXsjUFy85dgsR6vHe7NXtov+jazsEVCzXTVZ9Gnwl8c8iU9oAV+pjW8kyKP6Sift0T/u
p2aO9+Hi6kUxHW9sCeollwQKm0rGJa/VBFafb3+b+xlozZzaC4s3mXZ2SiA2M4x5oXCmJN93tjw+
nFc03bGg1tHXch4QQ68KuHz8kP8A60t738Dbfv/GkN/dWcSmVfA64KsRcOFt7jVmvEDLXwe5Vg0X
4RV/SxZgUWaFVD6joR5mvvq5aA7ayfxDfaCzx174yXijXpaJMlp+FojaWW4+lS47AN61SVQIcHw8
fnMeFiysGnFbiOsxAIAtt2SWtu+z9nES2sfjNL8kpYDQifo8ZX7Kqdz2WiXFD+7M3KWqrXbDC7Ko
iPNft5ec3TRtu5oL1timw0yNcsOGl1NRhYqOzw8uMvSv2qDAEZlBnqNm7CiUNXGrIBY4ZMqdPan0
K3lNXBPUUFd1k+HPG9/bT+wP+wLDOvFSRvxjyX8hU3QXCCs3JBZ/DRCXK1BhIm4Exe7Uz0YwFErm
Pf4rSrz5dcozLrfx8+cyfPC5JcMNUAAS1kv/hpPU1H2+gkiZh9ev+Qe4FUXNr4wqJCmn+aO82G6u
FoiP+akrZnXBaPFYzn1+y0UEDvXTnKiQNfq4BnceXIgxYHk/onuYsuQCJhvwzJnEaNpKsjcMF4go
sHxvHfuy2JxdZkHe9b3sgFc15Pt7wKLG9vXVd8fVbkOHxLDZWJowwNuxS7ue+cYGPcfbzzKfeaay
zTok4aAcIIKTKBan0um+BRpldi1AP/8bANwbRz9kyQxCibbKTMJIhF1j03ov0h7sYl7911FFh+HI
i1UbLW1PqATGN0PjI38ak9ObN8spZKPXEoGT+n3SFxbtSEVSurfyPcdVGD1p1yrPhQpeIUksdMsa
KFy0uMbmxwW0KePmc4GZ2zGyLEFSRmaOxMKyZbJxjz2sHd4PiSe2I+BZy2V/tUyxTwnjpAPSkK3w
HtrL1puefGOhR61d8Sc3sf6GSTLlZW4nbaUkz9nj51X5KdyDVf8+4PL6yqkdwDRH+54mOx6hcESB
1p4iFMnQTWSAi/QuKkYlSvBZN/LBCGzjKYqvbU5wxCb4Ud9TLtGbBhVsWKpgAPRipt+QqhyyWX5h
XhnyHtai2fer60uyr8JzQbKrzwACttUyq8hBFzK5RnLyIQ8OlJuop4TfAQpkEN0e4g8MXry6WXMP
psP50np3F8/aKMDPPc5av+Jl41yopKEroYc6xBxeiSNAqX1AzhCOf8PVAFoJO0FEdxCPa7ZphSn1
rzUm2MdmphSCBAT3fQ/rnoER/RuqNkrEb07HCvzDmIikyWBrtO7Gnpow8JH/bxDPjXSsY988E9+c
49aph9DcZwa/Cp6912xFErKfgs2pDrQ2Q1sP13ABpAcF7LyhJ3JvquaDR5V9SZTx2CEoHpJ+5/kY
wDjC/iYQJc/bMzulCFzDJ7cOxdY6lskhxy+hxNO5p7KtngxZRdVUdPiY3YMF26+JSjiiVQugosPW
8jI96VoOXqyPzq8+VfyxWECjSYv7YhsL8IesNUP4xysCg0jvgs9AVVXa7zbMSx90hWxx5SLCuvo1
z5UhfGX0dOHcPpy+k95W47/CHfW3YiEY/QFIUFFhd3ranv0LbNEBTg6nBsjVsdjF2go8NVXJyfo9
767vbUhTTO9/JZxZo0aSVfbCnAXikqUIHlcBZHnaE24ahmXlHrVVNGJwhNsCKKBdRoIkp5pACTFR
WW8bjVLqDOtrj+i2+HxQQDmhdavNvrXuhf95NiaIb/gg9vwBa8Z94lMsI1jJWuDwErXFF3cXC0hE
2mQhwt57wRH3LjshznkFLCBIZ2B0vFDOW15OSvNRBRsLGgOeuDuEv/7GnFYlu/8Yp4R66SwzcBVX
PUBtOjRlhPAGVE6SoSJMlm6xtqI+bi7QsTbUlb1pJE0F/h94e2MLdbW4l7b+NgWhgU9JglnWalWd
Han5fs8KTBf8wXrMHW3mbt3u6n9eoGky4yVuiuhLXXpHp2BI/pBS9TXlOfmFXuCtsAYfn8nK4dor
O7bVRdH9fTjDF3QbMcv2cHRPmYQ/YW5GBkked6J807ny9tKRwLp3yBJcmGHw1Xrl0qLCSCrhsMcn
RNO7FRCxr0vUVENwpdXISgLjbcT+dunAVD37AzFl0vPC6wkx6gmr+6BCtadR5qHi48vXwGPiQY88
fCM4VLINjjl3x9/oiPZhWhhSC2SFNLlism+8O6O+VYoo4t93X2WU4W+lBlEmsYes8a7Iv5QWiVf9
vIKQjLTSLqAD736zVj//WJsPeIFsIeJFlSl9RTZIg/to6frT4moYYKr6/V9NAWcRqa9+7YjX5BqE
N9oX3UkvRLaIWaO0Q7jQr8ySqz6tWb6iKwpAQZIhpNbodZmpOXRwhyEEyUWFKb0GqeXEcZWcO6wx
AxgeNXzg8+TKQp4YJmucx8A1ESJX7DXnAbssbpKHDnfwZ37NWqzsr2v6PJKMHz2DfqmIFNwgjkfC
UgSNAK0D2mU8kZ0EWda6CpTQnaJCZ27scw4cdZYQs3wNAONiCIe7499D3Ruqfh5/ytUy43rHvC/k
qIj3825nQzf6sJI1XmvVhYHMA2WQkvs94gUlhsmGB8a0P4bFTIrPSRqND2iZ55CbW39C6OnCKPgd
Lykj+QGyxsrmaxQkuWvARLIN1zdGu6k2EB+wIJV9TqGQ7pd18ulcawcKpygjTYWZmoVWEDzb7Uul
x40/oJOcYyPhqtNjJIWF4AKhjPkvfYWmSVZGVcJdhrF2Qnk7RaywxJ3h+vlqeQUC2mLHjOUbHdiW
P1eL3HxKgoD85ynAk7pqk3kJpTqh0qg0pNq2KPKYeBt4AieIq0M0+hyt8kX+ABidtgE4dotOLffx
mZGPtq9SSJaq+qUTjW/jhAjohntXe608NAH5fTQsEZlU6fDY70zaS0V7XamFrUJQyPO6f4OKukGS
TFDdli1bR+fNjj6BFVB+XksEMKRjH7EukMC01M3MwkJ+1DrAnlyS29YLo/AwsTcn7PhXIKe4ASlH
toDpEQjBOF0Iw/I5EnQ9We0iTT3tJ+0C3ZinF0t8U/emnkuVUoFaQo8hcc4mnDtuxLVHInD2xi01
Qy6GU5WvAGqWkVSKri3pG7HSKxwNKOjbTCOCJC6x6QCQ4NHQob3MAgYm5gtrIAJyZF5Z/6EhI3d+
R8xi3IaaW762yNPr9ATcu7TH6K+6pLxfvjt9Z5Zin2KBQB8dq7/T4coGPeyh+MXXibOEqNjSCQLd
rfPSIhvbad0ieNE9xkKsyGdU0ZtFRfMiNA5zbRgd/lzHmUKhYI8zldHjFHvBDIdPwDGmm8xyedtZ
vsM2Se9Q2IxyzyG8JAfMTFBMHlvngtqqIrRckb+UEGjjrBmc4uuhRb47GOh+lnfKTfySqZB/XwA+
8nxC8bYFnbd/gBfuYEYHfW9SpiOxheYATuWP6xDwsjNBokeQiESPQRrBkIGOMzJX9Gb9EKn3YlOp
hcxVW8USRw/Kkii94bTvLVzY9GGPYkgDZbl0KLPX4Oj1xQnUDlHqxeLgzakzECNX9sbyGkJ21h4Y
2Hipuk0uvjb/PBTdc+S3i6sw0FIpWlW6uykjgweEz0B3baylqT/TdZFmLFZ2pxTQ59R4c+/07wcq
nVL2xc7RenP3cGp/YKikR6FKwgC06MzaXFXcXEMN4Ij88uw/IMdonrlT02tIbN/vYHyiGbrTUN7Y
m3KMF5+x+5OR4LT2kJe2mApLqBWk+LhV7VNegnnqSIFpSKP4oWd21gKgxUXwQP+7vPBVOTeO7WQo
uF/AmnCeKq0ZSURKbzx3CXCUBdBUO2yDMMCzGCpkoI+uBJRWEu2xMIEV0ymf9wGIhygl5lFargiU
nZ5vlYDb8JWXdIvbxFQvn1FCZ9K0ImhwCvwxWZmkvVzr61G5Hy8FlQ+5v1E/iK/JobmTT1NAe4sN
r5sVXIrMsfZgO90p6S0+mc+7+yeI5HG3eVtcJ52yyl0U0I/mZOhBSxjClJ+x75rFYhrBHxWdmm5c
r3wjd/8CC3Z88v4gJ2PAFXtkm+uGSnr7jIxDq+cy6bF+jFgfkH8KuVaqzA/PfmxmFY3oNjcuoLeV
KvjwU5fED4kePzApQoi/yRt3X3ZUuoSMKmQPHYb1fAFk2bnHPp2uyGyhiB2juY1A/4kvmFxsuJa/
iXYxUTI2v0Fw46UflRQXi8fyLADBsislt71rLHozsFuKkF/H2L9MFMaPjJwoX2UsbC4ptxmMFjep
wdGzhHsb/IX8hvBgA+1yaj3qJMKYpTtfQGZ/+wUrf5yYWE3hQfi2JeM/RsDIeZu2Ux+WnYbSEAvr
5dnZqK4XTdE7EjrtS3RYMVAv1qzKblokEm+uiW7+cboHYwY3KdQ4/r1ao/90MeQTH4biLDAbwU8d
IisyAEH4tDv1AqbSiilZUzsGMgECrz2NHDFs2n4P3RmaI+EHWtQ8NUDNdM2VngssxMlCsGjE2ueH
NBNUbh2pkVWEBP2rt8QaEXmWgTJYPn88ESYos0rNz1wJmxAMgRLToyvXMZLw0qA2c/FCDkmeQSE3
c5RFD07t0Ei81x/zzq2rPSb7ISiEgghtbSpO+Kb1IZ9zIeul5MFq7F8O6YLCavlHDhO6pO2td8j9
CqvCCyay0fHoBs58Q4mEkXN3ruCM/5/mXUXXeoJZtX/iZf5+DNCgLGLiLwiUIhcJzmCApSlXmXkp
B1+jcERiJg/SpJ8Pzbfy9LOUKeoAA2mcN2dYf8kV1+/bxjf3ek6EBaNEAAg5DqVgV8OeE78GSyDU
EKupJTcGa2uVsOklfn3/Ggyt/XxmXdF3A0wA9UqMC9VJ49FrzeU9/CBAWyibaJqIlOvRC5DCpOKN
ljK4JJCNelY7536XpDuHBVNmFzQgeyt2YDW3+DcvyOHZHNZU3i+hx/unHH1Sdmz3RioaBg3v/Kbb
6FsuJTOMITXfIDtTG8/3gdz/tWlBKIO+D3/fa2pjzDCPg5lSqVekho6atycPPftT/tgH5jjuYXnT
3ZprZUXDKH7TTAlUCJxgaxkqI8mwL1Vi8AMhrpM3gA2NlzutM4+/zvPmtmpXr9lbeAm2IrZsePJV
MY5z6wqe5vBwf1MCwk2+uZxGRLodr7kOrRirDRpcZdq959etrp2RXE0tRy0R5uxU2XO6lf9t79Er
vj5wggnxYUN5lKT3XPjslThMt4QS3wBKAV4lFoFG69wGtii39rZzyLTNs9qKLpiypA8/e233dJNm
P1d7dxPLHyCntF1TmXkRxo3IAy992Dc0vNGtcDkdLNdt6xSp+sGVSgOYy9L/57aK2zc9NageVmD2
fLjQr2A1PnN44PYXE+qIX7h+oCpHQ+leDsvvkiKiylhW4ns58iTxGJpRdz2Si+qJE8iUr0+O39m+
iglB8PrxckbCw11rPHCGSAfSl2DJPTJR7WYxWSrT3bTAiuPdf+kRtsk+IW4skCJyDRufFDIKhlWT
kWM7yQy2OvVeZDxWIlesjKjsJPYZ87aK5A9TMXZm+o8bEcmd6mPF+e3NUNP/FTsgQrYx8hCwtrW/
vKDsbS+hzFP0FghG6YlgFBuocZubzMNBeV4EyCUXI+FfU5thFj4GeFCOrcDDT2pYMTfOmbuqrCsY
l2JDDTDaOV9aFFJgLLjHZPBNK7elTw/xCFrUeyzzCXouRMC/gykn9yVguFLvrn8trm4nvtbvACJm
ZWWS6VIfzrfDG8cFOKxJXa4WvNDuA2f2FkTogiraaFWbbQ470NivqawwF8XLHYQTDhI1tZmJaA2K
wjxYIzLrRv3WaU5iBmhvUDyzb3ixhfrm/6gMucG4tyIjPvVKU0tiqbOtPaAFIAt3U4swz8nxEjT0
PHT86qDdYexQR5Af/FxyOM1dL6W9BZ+0u2Ob1MeLXgYa/jUHuUoYfPLpLVMQUEdUEbo0xHBk5YUn
b8AxoHtCJLdRFaVf2j8riMTdndOGuDQfznMQ58OS+dWiEhYpyCciCkw1K1ugQHlOAaICdnwRFoKR
B6dLPX9GhKmXFz8o5PGkLfhu5nPvYFXeWBmeUlANHtLJ1pTN5zyjWlsfsEAfrmY51P9+t2BrNJK0
yVYjGvvdcE1h/9w1vcSIuaop/613lMwhDXyYrWk24jyIvxgwVFz7rw3nSazcgaWiQJoChL6/YYQS
gW6yKofA48TqaA9eJfuoq/X4C1s4td0b+KbRQt7HhfoQIXpfgQxgosqprKqY+u6A/pyfR+/e4zAm
8jpbSwrfpwt0mxpihyI47nM1+3g1/V7HPigPw9ggWvmqBhbgGnYx3NiUKDgjXipdxh/OAhWwl/hq
eY9vlrojfz8TtroU4PIWl4KhygN0ZyFFUw3TZ/nmoqNhExc5sEKfiJ7Z59mkPKRVDek4ffc1H5Jk
LChr7J14ZL/3/C3J07mqlAVZRflmfn/jb6XfSrZiDc4ggLgAckMJVDY4VwfLUcyrAeRJ2jw48rL7
WAsVlXFmPU/gk/2t5PNgY7nU0nJXaxWsF2D5qIrYY/famaHY1jZi2Q0BgMWCVerPnxHDwb/MlzM/
vic3fJ8MmyQx33nVJ2tbJRuaO112+0QFN+fVqkeiqYHEhjKStdFnTPhHssFjGBt/FkfNlLphrLWV
lms0tWMFQuUOEM9kEoVk3a1lqq/SK6birag7bSDzSmsZlGfjvgFrqmIjcEXeNMp5fLjsF9sBJKo0
tiQY1xRTKv5qtiRBK3t1GWfqH/0zbf41pDwVz9T1FwS6EI8FZPMxjbPvvvp5SYxCp9TTDj8hAIIq
gLpSZ57xNsKTM/z4kTh28kQznmCzoWD7+ZZody2o5pRPJ8aUHp7Mk0iInEdR2BBlVA1DnLf2LllU
PCx0GdSFuMdUv3Gd7Jq0QG+JlIriErpR/mL6vEe4sgl3ZmwQv64z03degbqHEJuBsIuptroAhNxL
719WlOPRvpgdDZ4yGUdCL+CBzJbHTlJwnSzA94iz7wpJuf+1XUWFKFOTy2+gsrbB6SMNyb2zvUbP
ptU4Rt2rmkZcQHcOcG5Py1aw6a7sN7pMzlSKQ10r40UFZEWHl/kWAMWr3+cnRu0wYbdB/0IImJpe
ArSJ1drD0qizBFUNSZdmnqHxoMkvZKg0M35HBFOfRlwV0YuTIB2TfZcxNZuRSVelnWUGR4a10ARr
v/zT5SH4eEihWRe72x3+jMXx3Knvwi9ZCtKNRBFJ5GR26G+ibm6st9dlRPunz/Io2HXFxZeqTu45
J/pNOFKBI7NcSOQDuSVKkmy7Gi94pVpcQTo45E9CcuUC09Azm9ukk5XTAHZEIjlCMF5lV/Wo7B1h
6i3uo9HRU8A2zc31wgab3sTOgKHFn3AdUEdGT46bErODo9kmnyWK9mgEoFC78BCfsrATFXB5Gr+4
lwtjE9M0LD4LPRzFEuU4QPt42/KgdnJVn6KqUmV+pnCwX8TWzHw1p2l6wi3qhEeukJjZlOfFpQrw
K81f+V+jIFyVrejv4w5XN7MTNr2kBZSNZeZTIEbTxLl4M9j78RL4CsM6e0Jw+pT7HkteI9z2Vi6f
AmDf12Rq84RIsdytyUECXev4oOTbiFnj5ka3hJ59YiEh51CsAUpkWxcxmslLwkTeNLmi6rkmVZnV
PMvtvoltSeU5NcTtEvDQBguYssWpksnklePVWkEmp/S3t7THc5mFXcnsvodHGIS5iLezgRkAtSCv
6D7ev3rtvqAzoT6PmNFL8xtwsAlwB9fOTO+iigxdy9yO4yu85ozSalVsdMjkJSKTPbtAXWcn5V5I
lBCZPsk0TA/Rbqgiipyu7GePnoPZoHZzcUA528xREg5ScRxxXEdU2NwSgz3TB3LnJfhi37FTHSgP
G9gGx8Fl2WqGIfz9/x/Jau9gr7noxrGjjWW1yDb7akq59da++RrQ0vRozgwp96gn0EJsQmYNbXLq
HMNfSicESi1nDW/2V4C/hYxCHivKOEpW/DnjBGoQv5FbmqWhUr2eIwE3EN8XbVW2HWDjqQvVgsuS
DXNrrmg2xt++HsyF+vXFIaydO4hE/UnfMzvNpOOKys9aq7b/B00BJk4AbHP9jX7iF9bCVe83OgHp
Vz5zTEEJMNCAd+8tNlVYKxZo9MwOpq6/Hl1O/AmibaYs5Td8o5Vd3ldLVvBjQpmMRpYzCkam2mZ9
UTqpBuD3oZyxAOOZsKMppWGlY9hR6zty4mTlnHxGBdtfpwmif6YdKiFlKBGb3VW18j0za6jf7KFV
FLbojHBP45XHV95/qR9OPk0jdR95J6EMozQ50RAJgR28fk8yL95WkEbNXFphUMgFKqokD+lBISp1
9xwOrX33ipEAjXJzWXkqV1aQy5EJPRfm9Nqth0eyfY9UleeskQErXdu7UBjbwD3p8NR2VF5VwJD6
wO5RivkskdJnH8kVOqbBcE8uFmhQxBXEDm/FOI1wuwOsZrdLODbZPHKOeIyxloaOVM2dGl5scnHg
9lKysijZYYNAcDiJnptmpnl/GzCiniRbE8wYgVnTcsh9jpHU0MwtrAE456tEMIPJdBio/nICQuFK
6musxRA8mlhkxIDc7aNTqcNP2Fr1Z8qmlHCxeiZ4OXgA9OxpRArua0XuikQDExGLd6TKr5fZv2Wi
Q8aZgwRU7vuwescJCiKSxRr364Pw8YXAEAiHOM7OyeMWzddFYY50GLOcFO+wVDsUF4Hd7d90VSby
WrheFNtzDR5gWUilrwiHlZLC5dO1PXFBXx6wB7xbd6MbjgBm4Cg+NiMtqa9z5cnTZmAiq6kSoyRp
DaPtSQJGqAg8zUlK64Qvucjh6fWPUZcN8iHI105dL+y7v2SncG/lrKPN46PDPNOBXf7GObyc/1zn
bv742O52VT/Za1kCmxTDOm2/2GpoxCGBH+wZ8G+CF+CsBVpBNHAOMUH8SHXbcYX+QcJ25SCqVnrI
Ah3uGTdIj52ipuDcyc7p9Jbcfpo3cGR1HxfMxN1Rkv7Y17YzNfqjFfTWQF8th9WmVgqCy5ywylf4
nluVF+ZDTU5cannVffcS5krprgFiQreVjLTvHuqvUefdr9HaX8DD8X4w7p3I5tVA7dBZCX30qc/O
CsJ+8P3zVlhLMsDETH821lFxnR32EJV5ukqV1aPqyrlmVm0egL5wcRevGzE4WPNtgrPbf54haWIt
40AVDFNDXiJTZL7aVEX2DyxZJQ3LxZQWNlAFfRF9TCLABct06ISqGr1R2PB51GAdJVXiRcNUAV4F
3wLaQ8Qa02XKRbwQt/K8kE/tl4inz/xTZpUFntlETz6n1pIQsJFlT+JuzEZD2VOyq9lyHQt4kmWO
iRM0iNGIpGnon5l7bnfT0gBSgy9FygmJUkfRDlyU7r7qzUeIESLzNl91Gy7EspiAy7DgP3h6RsU8
+hUw+C5s/rgXzBOYKdcStvMWrwukb6NrWEh0vBdEBvMwTzt2/9ajnjEN/dyNkPNeyHkfIoFp9xNR
+WE0K8ZjzKnGV3eiVlvN5Yy3norzS8mDGvBqF7bmOu48rasC3aeHW7SqHbA+2l0YRIzzt9VBnJhV
okEBrXOt/mQcTcJqFxUctRvIvB/8+KNRIKDLXWjm39Gu4mBzP/qAQ8HF1qMaW1uj0Pmr1GhyrSCS
UKO0z2NrOCg/+ZuuA04FHVb2Xf9a37zqIJVe/OEQ6aqLTrL6qAsMuKSFZS4UDQVpDb3ZwXmcIhgJ
6z2hrs4qUqc3No3ViO885uujAH7pGQZjAtLTU8SuJ3/2DoMURgv/RF+27mEgi136Yixz/+TxCaPE
/VaFGhkCe9feqkYCaOintjagDCINqAHB7GGbQAFRIYa3njOzi7pgaIHPbj/+QAq8NkjQHvktBJZ/
JgQxKbnjPr6Yu53DdyE+3Pi3q+aQgErXcCoGsV3pOiKae2iaGq4YLCXESm9jMaDFSAaA9P0uyiW3
KTEEbhswbPDBGSvehxabbLDCVL8ayUcJHOMaba7rNtfRUt+6SfPhsExJKzzh1kFtGNpuaLRWnsY+
4MBSeGa3ARqmIAgU9VpOCmQ52MQ+QYRWctKE0pE5QDP+RpwvwgJhFdtb5h1oIj0NJaYF4DiHVc7U
NH8wXW3R/qzh5UdjYsfW00vxQdesUpzNMJCp4AMTJqfAh76G+VPnjOT0LA2kF/7ZH2cM1gA+BhcR
kK9Cx1ne/wH0CFl0NQO3ekginainrxL6YyAl/Hmajb/AwazYdTekT1KV+VE9f9aYoEq2X6MUSLmZ
Dz9hwjQv9BKbiDLB9Nw7wklo++3DpYSNDRc+rLV6ZokCKYsFleqIIapWJT8sgk0hOLuv+BrzDTa1
5tofKx6H+AQ062v2V/Vq4bWJkGIdiqRVuEVU2Zo1kNBeE7Tt6e5D2DawnYjSAbghkDN15nMzlC/X
Jjwau4WPkix0rH8Fs/y7mEgzxzESw0dH071maY2oijGdE1/9uE0HZaqi6r+JmixQBFOkAJkdonMp
dEFL6hbFVJfxYzdrldIpdxumdn655suQC4YfRPX7XSVgdvwCYycjL8RLPFNdqu3ZFI/GYwHw+h9r
VKpQT/iPzizNHRN/86hn8Vc9sDUFoDAWq38RefXRjnZwGdWepk0grQJ3jA8QFudJXM3rqya/KuMn
vBGrT6AtBw352jQ0OHABJWoxcFtjeMv7ttdCZYIi/WXK9nu+KTW7qRQ86JBZ7LzyKJOjZSeySUUh
dDYnGBBUQhLGjsnnzVlqeR3hEWKrB+m1bIv0lXuS572YF6+XOi0eElcwNKpTFK4UqO9c9WnDjplL
T/9ZSFZ0pw+RoJ+uTNddmq8B7bNMdg80P8DErO0IuRwtYqr8Vky7O2wDGnX52w/nV31ucSrHc0qK
uA/i/uFykGywysTbqf9LsSymTUwF+6nU4cStlb0Wufd7xwDi1nlhJiLJ1pLwAadTxLy6JBAaCjzv
xOXWjzCCUnqnMYSYQFuv3OyRfqIFNDAwShN9D01XLeI5J6VHraargJoeFQR3HSgExwZbeoLewRtC
GEZ3Tds5/oct2Mc2YW1tLYXv10gL6/t1+euMTqxEZ4nU/MnAXrBuwp9IC9gwK8qgcsLGYwlHqQlF
GtuARirS4ZTiA0gLIF+Iq0G22+YvTCVEt6qr26CJf/zLLTVlLUTcufBXovF92tDc8YtW9uEl0CFs
/hUzBCkp0bdP2azYnOklbFZHO+0FWYh1dJQ0B3J42HJsElhpdd3faMlJTyFyHb63/9yUggjxa14X
WDWFJ8h0zByzodeXho18ZmOvxjNeKEiEW+nf1GzOBLLbJ9QMrjN5Yb7wqGr7JuKEbezsKbB3NvUP
rHHdPzydPMINSBlwKy6XzVLYxD8b3ojjni0gwYiv8/sJynjDQxqLIe71WE2DVCEBV5zepXXV2MYu
NE1H4bfdDxdI2wLO83oPUMMHtNQMnA2Z+Dc+yaaN+aLcN89ZW2Uo2tEPH+0rFKjIpTbSL4FendLv
JVQbeKNWtjSVc+FMqGK0FJI2lGXABVZCuWaNp6ZpfP+yCHPk3MGyFA2qZK4KwzdEeyp7/3ipHj3P
u/qAQ33X61QZLj+tRU1oIxZ5kJ7BDGNgBB2FrtK1I6qH3JkhsojyxmSGfC7btSOVZ9vJAI9RMGb5
jif7zF1t8VViYQaZw5GWv+qHXTN9pi1mI+cIGyZwdFtCPESg5rDuXeDsSri9ELaRduPucr3rctqv
3Ns33A9/OI+FS/UINE+I4da1a+L3LimKtFxdb14GtVTjJun2j26SzzDaQcU9a8w/pBU54dLCS1ly
bCde0OiSHLVA2zKVoBM1yzad/PF4hqueUjO1PoiTy0VFfX1YG0e3LVpFio+kK6MymrodYL7rssFg
d+8Ev1LbfjdN50hl/3mV4hMnmO7tomzKqW2GSPAoIRjmb9Q3a/7QXWAHWghuEZ6Sfdj+0UCv6kIC
kddF13ioYxeuXR1k8pQmGIDwGRA/C6y0ILoe5XrgGnS5C9m15r2LBco+/peqDUWH581IrOzCOdjH
ty165dwGhHqqKD6NDa22HERoM/uc0KjDbWMRWLUCgM4AoqQf/CJgR2guMFHLy1e2tRfZ00hgOTVc
0ZDXEo63uEKDy4nC+G22MO8HhlDHM1yUrhIh73rGueVzYowIsPdy/TAjvykkv0su4lS4J+p9AZGy
L67wenBTVn24qxG/2nk9kwV2tox1fVxgs+A2DJV2QcMvqfBzWDvyJQaopUCx4h47VRNKA4MM5tW4
Q0YeqTCsgV3jdkjukf63/Qxef3qqb954QJN/R0CGE1koYXAKy6LQ47uGm3r6+1r63hz1W4Xm0fa2
qYRkUWLk7S9xF1y/kHEzBA5eD8c/voffAhXhO13HW8DD/wr6OZColC8xGdQmouFHd+AgAMVok1SY
BxIjogx7fC0Nxk67bHUwnIRecfkPABUj1c7iTPWu1bODxxxdubKcMvRysnBUM8aKNhRG7YmFzRIu
8cWW9kCmj+EQaGG2/vOthkJ5EHJ83GoyxOMI2NG0HNCuLlQRy1KWmOJYnOJaiBhQSHumaaqVF/eu
DxHbbNhEjs1I1V/bnRMCThmCT/xTV4dkPhoAMBMabD/5q9lpTwZgeYQ4KTGtFzRBPqMlAUGje1OW
nl3qqIXjeCULnfi7YrPI++oY4UQIHK3BhN/VC6IAf71lnpRmOvLhxEasH96o/IZwIAPecIPnernS
/nR15exDEg4Ec3iqCooCS54sZfj7HDxcMZhodwZF3lxJ3Q2mcs9IwfV3SJkxAdoGtFUv7ou216Vd
FXt5MezHrDSLaOJLoAvrP/ojivdak2RAsRt9hT0GUk/LGnIYPRL9rSjJMDO/5pvJ004AUszqmnZb
3uWnGphIL5dpFATIQr9ar5HeRZD8v0U9mIW9V012q7/5zRa5XuoZftMIXWA7/4sH+f2tIE0KHg/r
QxqTlnTmdmyTKB5/j5n6xKRUoz9ZilCqwFglpXySgsLKZeTrUtsiaPQS7/feFUJFl64SobL6ByQ2
It3XOWa68trLofESHUdZ3AYkGbZJznA2k57eiJaufjP6fZ/iX9tRggBEdp9i9u1y83km9XHFSXUB
iG9JIx+1/bE8lU4Y9sPqvIND3purE/zKjHz06Vrv6EyEmLRLcrPBhEH2uvKzsk91CmQ6KeMIDUQv
HkrPCJnb8jwDcXA4hnzmp4V+GmCLvRyD+DBEZPCWaWHQ2i/gNWRobs4PkA/PlqrBUibD+2Ensrjx
1bYZm3xu1YT2HN8UZmzQbRbx63Rh2PYoB3nWelfpA+Sa4LOqOuqqReUfdtQbSkpMMs1eo7tRBtQ/
HTIxfivydvo8nPabcLbpW7nHvazcSifkaFBmBvsON2VZYToDz0NX6dnhNdikoNKaQ+ORMl4MyviF
GjdReH1QwQoKoKW/p3iOS5lStQiKDM9oU0004tHJdzcsaOsA7jZvcvyae66hu27OLUbgLeswVHDj
ls0HHN/GsJkdrKs9Z4xW7vodSlMNnN1Ddva2X055I0h42xCcNPvr66sc9tyZaqbZtumarx4e/pvj
7bOPV2I6XSp+iKeGEu9r/Wzj9Nz19iPVfSRRUoUSyI47dTePy5NfloNJ/EaNXmZtZkr/1SzUEQQn
UUUDnyV7Kiaqz7VvFPKg9efx0FlMWf45V+ntL158KtaOYvbpDJpG73pU3wO8hebrh2T9EJDqhSBb
QhL3OYgnHMdGOhLLiy++kNeiFgiJFVrayfSKfRww6nR2yRHOKrrXx3VsaD3zOxx/xo2DlF5ksJ1g
k8+8Xyi+QFscalHOeK2U+YF5XrtzbR/BLaxZRO47jATjaWralQA6np6bxv1FiWIekLirfgd6S40E
j2spDAvF6+H5uVd+kzj3s+WFbCmnJ4jzMENam3jfXuJTcwCIAD92w5z1ZrBMeOGfYcXQtI9STbK+
jDCQiIkPQRcDt0WPuIOLGCQQD2Fok07+I1X3Jfs2UedDVUSXl0hnc+7Bzjq3oOooTjNHiEf7KhKO
u8pA2N+bdoaKa+tqjzUN2lQTzMCmRiO6qo8gtxWuJhOjM539gYOc/Ne0F+hT2DIsG2Ed1g7U+p/L
iP4kas8bMxriVqitcOsPiwcYCnHnrio5K+j5wXF13jR8NJKYsRjTk+jZngG3NxU3C7UWzJVCnx9t
Se5Myy9J86Pd6x90mP7rDW/XpgVHJ6/v2L1tE3INfKee3w0XO4NvtZ91SvDdyFyldyli2hi83Dvm
VReMEpw4QFed5jloY4RVadz4molNmRMaFdEBpP/5HUtfPMSLvXnihEOsiv0QRORNy7YyZbvchabn
Ee+t8ryT4vjaSRnEKGqtzyrco1CA5fz4gWn2fVtChKy03m3QFD4Rrr4s8ZfbIv1sP3Rvr0CkJPBD
x3B9hQG/qmZJqPT4q0YAG24kSYaVz1rTXsO0pZZ6DE/2x3i/cLeLP0z3p3xGDB0c2rbIbFA7EVcb
fm0hU2+/eLjGrTYjxDfPorVGQiN8mRyY8C0GLvnez0vh9Kpr++Zcl9g0bAbOfiNpHmLGJ3pRXdDr
nPGwMt/rrsyKUm/BqmNNBJiAj2qSlv0/Sv0ic46vyWY4/la+nhsj9QVOz42JInRzqHnNaNpbg1yF
MLE82pMTBAmrHwOrxJvn1YXBIzk6lRDK75AnBitJvETdkBtTGUK/QXQ2IvsVPyrxv5IaSJgZjrzb
im/s7r4kwLNv2xN5GFoxonCqsy4wNk2qxz+adaaxJABTQksZpBVGTTlqfVVdj5jdDJp0EyZN+cGQ
r87HKDVXcWRIAKqQFpwgM40e7eC1jgEmAngrknRnxvqyfJfOSbc7X83qLJ6AK7wXK5cCyePPHccb
PENSotvib7Yfzp0Iwtz9ohet4P3056qtzbVegr5GPw2ed+bEFqc7hP3PWnuW9lbxZg+NFJ4KHBoV
9+5TFmWvcO7Vt+f6NJ/y9IiTIL6Fpyz89y25q9FIf9QV5gMT27eLqSyAmbOvaHVGs8tKlz895BN5
LAvjFPEOvPcifCz8iRAMDLOJhcaz8mf64sU13vK9gi0ag6DATupR9yARegXftbbMFwBUecbgV6o6
VdIg0N8XxFd0b3kSWzLxcykhcQjWVNF0CkPZqMUYt8QJF11pmtabeJg1Tp3gIo4z67XAAuoRij91
JXwQCTEoljicnrMSl/hJLYOAVQbIAzKoXGxOSG+IyC4v5nWxVxhq5vCoseRiIUTmmW27Q2zDsZlJ
kSNJSG5bpCtIVEt48fQ2Ff3nUa5BjxWWJBzv8emaT6jH93+dAPRyqsyfgHWNd/TJaJ7E5IxaaoFw
h2+7ceV3mYX5x9uyTNSjG7uU2E0o5hI2Vd3WNz3BZDRjDC2VJumxoGcxkKISlHBBwoa7L4N9uouJ
Wi+9q+vPdJ6o0aXwS/gGxju/oR8mw6aBLJw5vXum6wZWArYiJ++zM2Iq/6isVSeu8ywpuMOytymp
rvxujeCjuS28022joAsoRcuY8zh6cba+ijZc/0Jjw8qd52JVe3lFJ5bdOdu4pSMto+EzXdO5ngat
MDbghxl/IEyFzXJGa9jKm5FmTAbtHu4NxJ/boHFE+kjfLI/XcixONI2/CAXHNzXmcQK5g5Rqt/t2
BQUyXLqWKb9egTEZ8GKHKWtZCsI8UASnTNiVyzV7WWYJasq6Sr1SudKpNuswIOz4D+zVryyeOakg
DpcNREw+qy4+ip8O4W12+BkL1BbdcTjuBFigPAk0BLcCa90sVHkbDEqxTSVuH1K7cEVaCQ4S80d1
G6+2QTUHGahjzXdG6uyDI+PWCaTqeTaRNIVTds2Sb0Wn55WkTFhL4As/W1KRu83S7QMC7FsL/fBD
xJSesNKKfIiR9rfee7XiuJnwxF1fob8yqgV3S9Zk2PoJdogfyL3Ru3kgPHUu8J+ypqJS4YJe03qq
kU07Q5tTovlt9VrD34luLsuaBjeJBkUvcO1lBXy0gaGIFhGr1XdnvXWjNJq2nJqdyBrh8X6bnV8q
rsl7xOCMnxxY76kjenFgpe8RUALX7IUzkaZNXSsxz2/h5yiVM2EJuygHS7Lcwiq8KMH/bpExqLB7
oaGgMmPwC+6Iv8s30InGba95nJQE5YXa6VGBisKaVH/pwb6mpV5akt5sMT6YGnLKINp8vF1gjdqU
Vg/XwjVjdXXImioX3qwI1xQFBZ2hzxxHtnx2DAxcSz6S0ba8PuSlfCDVyrrZN2B3C73yYRZ3A3Do
lbhwbrnRo2Pmyko2k7baQwLv9HTxg+aNaoq6lYRWyfCxe6sZ3QBJqLhai/f8TOoaM6OvSFqKzLo/
DV9nHGrsCugo05iFHiaVBJ9PV3PJTZ1mrzaZy3HWb/SkJhWoUunBacAvh411RKCkkNH6p+4I92E1
o07j+p5H+2Jr2HBmWvrV6U6zySHwKw56V/TvpTf6Y4Ri9U9x4KUzeQVaGFY/i55SCitxktybTzKC
NaQ0eRhnb0OYcrbn3obhYNhXjeBjHJ3wv+5iRz9yUG58+fAVRl+kB0Xt2HYpSuachZO1u6ag1gq/
TsjCbML2oyBxhv2yKvzAjpZzGXmIuN1GweqOkcuZ5H+/C3LvaTxf9h4TTNhz5BN4AgTZzPWKW58h
Jaeq+9PtqArTJE55hjsGSL8fs5YK3RRkKsjKomJb0TiGXCgJji08PQmxV5DOO+czCOLFIk7Kr8UF
SX+FqBRObd92+VmTMz4zoOIpqyjQrWxshJ56sbQA2qPBoILRXtC1+TaVR2pl4OSTW/i5IKOM4v5X
+xEd0hP4JXSqVU00kq4QjdjmXwJCqB6uh+OyQMhUp9HcaMGCfv6YoCfwnXBxxpaTX3w/fsQvXluP
GTZZbIezDW4O6wDcFsohrzhkvWl1ZkIw3WAL1R9Op9FMtjHGvD8V4wmoLGf1NAkNT3d3/yu72xZX
/RZzUQ18iqN/d9lLzzjiZUWTMbA/JJBU2rwiU1US1gakd92QftrtZvO7eNwzORoevcrMW4n+4AEJ
p60eA1yuQq8TjepWPhANusVN7KzV5SzQezplLG5QJyOqSAc3vPZ85yxhcwaUpK2g3xofDimd9sK8
g6wDfiMUI1cWwwSuefgeJHzGhh9gs9JT9Zqqh6zSzDKRck3snu7Segu1o/DpWZGTwQdnhQneMX7M
Bf7dOkpiKe0NbIWcEknc9QVO2N4E7nSc341XlvE5GRwu+swlMOL4A4O53KtKyWyl8YGFX3PF1eBP
ECSvESvVfG2X8SPX7TaKK27YXEay0KebWOLtMy7nCFdsrWK6ubWysQ2V12vKyKaTNJsrKtsQ+W+a
f7oVqPFXO2hhabTQrZbicK8w/yDO9y/FyKAEI4OrQEPP/b4U18oqjO9A/XjfFipXU1gyuLrbToKH
JK+kL+4ZOan8cphxXiACApjOrCaICI/geeSV4uOve1jMJimBJcNQc4FUrscu4adY8uqF8m+G656H
LWDy8wGECZpXrbrd8KZYt2b+RHv5jQe4ri9p2B0IwlTLOxVNQwYZFVbTacbLzFhclHQaz09v4iPS
qOfdqCVrv6oErDNx0MJb0vbBAPJOvzIepg2prQKIkOYmDb2gpfHZUndMi+YFUnWgCHWpEaeQ7zno
o14dF00CUQoK/bEOW2Jczf34YLkPdVWiqAr2wIYZN5mlreqQ/Nm5Cw2CNehBO/x3su5fH70oiOmi
B07sOfMbZk6Nq0uJeALLTjtLLTGqhDnazT7zCDDRpQj9P150aGnpy8xokOJKRzPlktkRrU8NmqnG
shIz8a3TXDJnpGHctPftL7+VVxD750snx3LbZzLCQcL22WeXRgsKsSsx9K/q3BDYmD9Tw9AuujbA
qUKnh3ndT75841lSRB3GnowvAZTeg/KtCoVjzRwhBDAkgXAbEKc4+o+iitiEZkk9jwryIhFgDGZ3
JKdAIrS9bStaWyUS9CBybhJlM8w8xEc1pIkSWonf3S3clI6XbTsT9fUTxUclqaHnY4Rpw83DWvbs
d/xARBCA8pvvG7OOXP893o4++Ndlnwl7Ow6RlsfDt4IcbL5d/W/m2j2LnSw+bXUI1jAZy091GN00
e/g3RXn+ynKoThXRqbJ6fO7YObaywfJy2RMLCpcnzsreYW007a/UqGLbhdfhytxBYBe8OgaIofUj
uFDkzDX0/WP6AwgQPwVxo6Xj2ajwhqOg/9Le07Txj81rMV05yFcGBjGoznpZMmc/Lt8LWZJjgrAc
N/JRmf0cG2VM3h0ECCPCkhhoVSEUbA4WEE/1HguickOyrY5glkh6SpCOamd4AZ8pXt1llxeP0jf0
BPn8c39dMbTmososVYSL5Pofdp9ev8v45OzXRfRWx2cORHcV5dhqLY5yUViywTPiLloHgKLRoloY
4j9Whna8b2K+EZb7EPRk+jtdrCKvG8tCwVlGrmkABKf48wYv+GpK41DOSIBBXXglcUyS6k9BjJsI
KGudd9X1yZlPlhveGuSiV+Nl44DjZwJ5UZLx/9sH/8fE3KgbCxhJ+1rxQjjpm9LOo8DunE6lT2du
GCUmm2R6rw9LreEDdwMvbsupjoeC3vPZVDWzs8PpaO68aIaFYfwWk25iUGO4e0xkfQfY0PFZ88v3
He5izsP9HVNJAIz7BU3DZdBbnC57RIZGeDA9pdl2Lo5tEfar2W7wwQQkdTfBz/cdnvaH69+8s1eX
vgnXcs8iuD1/FocqRdmgOqiDPE6FhJ2RoegSr/6E+AfNLgEukkT13h50Rn6eA6+Yroad3nrHnPp5
CePJtCBf5zdUbpc/gBv3V09eGxLNsOgFhJT92ajErgVEchcGRxF9PmansTMIu4ELoftVuRdTN6mq
ZZ5MQrPsLW4w21DBHO8fc8Ymw6y37goOOjY8L/3oW7WS568K6E11xlh7TIHWoUoMezdG0sFdnDDE
yHdv3b3MaKIPF3jFroepywMkKFBjrgrWpgNGBOqAy5oUpvKINj+o2EfOX4Ccw2BHi6iDZD1CQFlZ
yC0hmdr9tCiKCyxSbJ3m5RzBgZWgIr603fjFrrLu8TSlh3phv6jd5n+4Gbyz+wX+8xkaFZGomYWD
0W6sqSzDDFkMXPiu0iPZ5C1yWXcKCinlOBE+RuYN3Y3c5GQ2TwxAImhkTfAu74wOzp2V2Ge+LUZ/
GdZZPv6inalPReZndi5LosAoY4PafiKsNPX+IYYgfpYULunMKf6beXp8S3jIYdWNccV6LofZZJNI
3pwZ9SAHe47Vhm2IL+/9jt1AdgYBYb7R/B5seTxxnsYbAxOT6YM3mEN2KQ4uAU+kspsPJ1RgLyGc
QNiayQJb3JpjfDJ3FKRgWVlfyszISgtUTw9MbnB6klsrUSupqP9ESS9s5T4+FKimMLJVJ5Hc/x2D
0b2sszicUTcea+8O/LfsJdGism7iylNy9AVZOXtPap5DCfMTzEadeM4fvkb2V4DDpO2bBO65RCEQ
sT+eEu4Ur/cd0T/plMI88UOAW1n9m5EBRnMNNtCFCZPRo5M5UTpEOGOrogGi1/ZNsaPcRa+PVNWP
GeDKpodZ1tGjQ0Ix7PB7BDJ/lXktDVDEoJHN94GAwP8HYFWGyy6gkTQmtb30Z4PW5kxCSHhVaP+u
K+G+qiUs8iQ0SJ25W+4NxFzftv8OWeP1A65CXrhf1sx/PmU2yLCBh0YfelxkGpsvnj5vQymaEiy0
kc2q86ZH7qS/kohiop1wUhwh0Au36xjPqrunBCchoBUKEM3GrQviOZp0Y2Z3n99btkpIX5GCouBX
frlhnmeJP21oDQhiB34VCZ1UoMvawo6B2td79uQxMEMjG5gIEKsLMwItU5CNahhQfglrLS+pJGVL
5WU17sIZSQkPLjFuapsBBcVhPm3YxVqzj2WbowtdDty6FDoXts6vqJw+JfcXvJjlpw8mEdt4ssx3
+ldrAz27CIwvntLbr5WOC2PhAiXXtXIJbERBAtbAYdWv/4IHDaR7cdFomWpTXDumrylXSbc5FmU0
YjGV1f2nB/8g1LcMSB3qFPOjI7tOoaccU8ebYqbtfZX4CD9NaOBG0xdYuZWk7xCzaVfgt4ZC+KJ4
K0L7tQzJsk0eFnphioSMelXnz/viUAdveIKqMfZCWMTq8oOxGA8f4O6CZPebEKSSARgUk3UlHIJr
DBWcbqdMeFTSXJNPz0XMXTE/WOR1AYIQ7iqd5Ktfz76qumiqh7ge68yX0Zby3dalaggzZFExlsb8
trRGyDiDt5ZXqq2x8JVjtQDjEETKdRYd1almWNVIVAsbyFPndSLzhzbXFm4tyC3zBMCd9+eUb1AS
OAeWUQvYC4MnaL2LpVpYghVfxMTCvD03xs8JP9hXROYqc/uT6fOzwPqOqgKVlFSUuGmpy1jQolki
1rXsxUv1oBALgqYIuR5wQtCqHPziq3mWG7ZAkcbg/jg1XFB9H1E9fKrKABB7sjlDguWTTHoMDi6v
9oehaHIq9WJa6qeHNDHPo08HlYCyyhYjskXYlFhnS+/e7xxfFnrlEFIUk4JbZnyjeWGV7esIQvgy
Aq8Y6ZeNoLg1iABhZ6n+Knk0o5LVaFtLnCJHaaQruBmK9fxOQi/606XPUjlkai8N6eup35kRw+MX
wiLG3XRmwtVimVRSaYdX/8FJUDJvF8i34XyMl02kreJT38l6RnouecRL95L7R2SA/Awvnwq7l24A
q6wDwiKLNbm5MoaPt4LqkyWe7Sa6i3u61RF0ySuklm6n9GUE0dyp9fsi6RN3K0s7TxA4lpaJGB1j
vgi/o+Ma5iMwB1v19GQPpD6R801IJNuXEouTeSk8Gwx5GjzjuZA/fowlNNiLH74WOv62sIR9lNSO
m+2adeloZR4vs7LkK+aGmXJT6poNiT9Ou3MH2XRu549GYENJq1kKbRObMCvoLEAOFKNIlPy4vYrw
nSRKrFS8xDJV+0XstFp0otoG34n+GEtoAKBlMdHIsRED8Ca4y7R1xIPenZSR+qWV7ssNouqP8u0Z
H/0IX52k+IXkgJuV/U0hQQBr9wdJY5uM5ofJ96qr17X8/C4lRtywMTXmAB0ZHb4Hf83qDL2wmPcw
hbwZubdOH1gQHlN/2z1E6IeIEw5HnCr9slQAZzlehf97qTLlnFn1OrnShc0TO4c0WjSQflNPlgl9
W+DxhjUNDGXChKbKKBdRnEUcV93lCGZ/jpQGUNHNA/33iXEmBUekJQqM702Cvgdj1Ir+7KKzkKdk
idDRd5szEMr02KZPHtJiJ56CV3Gg9x0YGffGXepNFfLlth42Op2XzokLz8R9kSmXQ9AO5cjKDa+h
O3XW7IyCQqbos2nPcrtXTZ1bkY5DJZRf5gRHVDnyCSSIvAPBcfjA9Gjzg9ouXQwWpzyEKOGRK+LR
gxh0kl9s2b0DoRTDkP+A7RaenyYyE2wyJREDSJW23niyB7zSD0Q5MS8VQEfMbPP4CKG2hNgbDF6H
Pp6UB6dT1TuPNf7IA8MgMOhpZUS28OOLJDEtzu+ZKO+AQOHIc4YC0AVYsPquwNgd48lXOE/Vn0Fn
+DCYHQou627NAlsArCy01qsuA6i8yPkwC3fBTRzKp7yARqQSkYwL5v72N3SEvK5/QwavLTjl2Cyb
C81sNEmgvTWKzlVnH3/mdIP1ZwuqbU5TIQRi8a4sCCCyLD7WIIfd+aCJOlhXyKr4LwA7FbmFv61B
FiwMQpngKl2FW+aVGdago386wJX8N8drCvcO6nwPadKyqw09FZck5J2u60+n5rD7umcKlLDJoau3
rA/xouMvaOI26Vzi98EQt/HU5NaObzj2s9Q3ul3F8geHBWme1LKtgP8d+hKV1ks3BlsrRet4/pKs
xBzxk0WBYpQerKsLhJYE82hFR2EWGMabjg4tUvw6nqyGRT7AzWq/BKHKjh37LXax+hYWtZ7cP/n3
yTMIKESl8+yxdT3ZzSpaNYW40OiqGUFAWil7qRf92+XECWM5pnp3gt+kSEYeQZnWEBV95cOAKP8i
LSlBdd/Iich/zjPueL3dp0RVkm7ZAxxIwGBFbi1Q3bX4kv2mwqFDecUYXPKLrdPlFNbV8FW09q5U
nIRSGbo09VIPsBWlM1S3I7kBGAg1x8B+KRG82X3lUpTocOgOihLb+ek1cwbmH0KwDvXdPBCfNQco
9fPZfzxG1UZPrKSjMFEa3+zs92zYUavI0JMOHXFXV4z/YHwqjGnMQFcrrKLjerYLDl11carP00k8
BerIR1vR/3EwNNx0Fsyn7n4+K7JNy+Rk/TscavriSu0D9BRcytAlAx3Nv/39rpC9Nqi0FodNlXhL
DuBOXx9V2nTfieqOt3bSJGTCgkIOdBVZTVQ3y1JHU8jsT13ORr4gasdlM5enZ+GP0bVWBujWgrs7
cqcg2uCKOUZUHRuAdEO3FFOkiZFkXGDbKBJg7yMuFlus13pftv8C69p7wIUmL6tDJkxBKfiKeL+t
N+aEtLt6NMCo+t/P/YQ8U5HX2Tv88eFuhBtlhNo5LKQOLp7ADfBeDJcvijHcnD2g14AT2Jm4xWh8
pUOkSh+yoHBa9wMjxh3xXdnWQx4DOV5FyX+gcSLdFIye/A4VlpNbcSybKtiNiZWswmTG0HT/+QwK
8JjQDk00nsOzWcmGfxYkkqzXVqX6rBR4WXiEp+5Dd5itrP8HPq5ZsljwOZdFvMuw6lwcF6i0Sv+1
QdVe3zkQ8DTDq/g+SbCRkP6ar+Vk16uQ7Bjci76UyPkjc3kUnftymWUlezwtMxQipG6JUIR2Np4q
kqWS9pHvOnVQE94szqjz7yMR8NTr4eb2+/Jul+BHboyXFr+lq30JFOzXpUvQS4/pO7Ji3tQg6oma
2eL/8Ue5z14uTPAskVN+tX9dEIJ0kwOeJkcE57Tg7NA/o6zYf/OrjMQEP1c7REVDv62fohJg//qe
SqFhuYJNZ9hCMLQ29eznWcTGpBGY/TdYnxEV/0SS6RkByHjFrKGfSZVcRjsuyiHKXGVB6lEy4x8J
mYSYatzlWOU/qafhVcGokj+4ieZpsBJVP75l/6Wi0RgG1Gx8Y3D1jf84AeGclQ1L3yCy6EGmEOzV
9Tz0450ks/cQsYKeyo0eT6l3qARNTl+hkPC0f2rlXGJcFImvbVAtmxe72IOLJfoeWqnxVTltGXD1
rF1cdp32WeO6vs3NhBN0XZOD1BlJEf95Cwic03+OW1i0stYAhUKkaJ4AfU85w5FGgGhutHc/RU/F
RMxr1vxYEyU/GGVku/MTdT6wHpYBsWP5+N6Ylw1xIOyV0xXsfSzTr7yzDy0/q+ClX4UjQ6tIEldc
Ik14CPPM0aedlWpDZxauNCDBSG440axMbqc2D5wI3GSoqy3UytNxxcdCtvYl34hr72ipGvzKVA8p
xPxWs/YHkLvRwYQGGnrZRe5+BI4AoeBLXbfmxs1/3JV7/cdnyADTBM4dg0YISxsTsitZJpNO21PC
AWj5YPeBX1j6xBL0pICx4s2QXdZTszGxYng1QNVlPh170gmYYktnOVl+SI5uvV3bIWQ8a40LsjvP
H6StVvRA+FQc3S5p0yk3ADtmRfwqXc/YEmupSLuYIbZ483jTHelE4emxzqRZKUPNBpLdMHxqnV1l
uFyMwxXic1YCsjMKRlWAuiWHwLyKH9KFYkSI6L2mzb4P/pBbx0o2C3k4OATjfK+MI8/gt+m5HMWJ
7LYukzmX+3K5jsKIWN4YZi4Ny/iL40YAnf0P3l8Gr0OUv1UkDgBGwLuPGQ596VeYN/z1iW1346zl
gYGTIh4JN5cVH1IJSahPEULLZx1SlBpcHvjGKV7f7eFh3xJS4Dp8avhQTe6DR+Bf8lONaWEDbgbD
7aMsT+QHAzxXHltMY0ujTno9U1cCmu+Ww7wngZ+dYIDXNuMa7lHWwu1NEXS5ZQee/4eWIMLHDuzd
85PJ4gpYVVreP5YYoG98y4/Zj9w8rAkOGLUjCptcVoetD00AYBQaCzYGIIhcByGDZVHQLdtoDCh3
Z30tgAeRbUBczJ3DQpYBJp6oho9DzM2WVwjqg7e0lJu5rjTlpbbfYFHrCv/Ve0EG6XzPIgorNnz3
QG/EVHqvFcBfmOtHTWODtq9ZD1YDtK38uVvag5QRUmOULdpmRnai4ncgdYMYNqZ6D8sLYvBQwMr0
YfUBM8v1sgMCuXU1JAJqBW+bfw4r6vpTyzAZ44+wNeYxY+hFjAVLRglAunajzaT/2cXVagpH7PaD
3xcqGlUZ/3KTiUzz/HfdCbNgPWA4ce8GR7j2+Na8U/IVAmHywCppoMImO8keGtAbYySCuAlGTPk6
3dxQJD3OTwN1DTtoKeBiaPC77ejMYIXX8rHRwhRUMjbgoessbnA4kXX/W+CAYeeNrrBXTA5mSj3S
+qpRuBrS9T/lhB27nOeC1j3HOCC6erE7UWQSu513/Ph8ZD59YEoMeduIIfuOI2FQzfMOQF17b3H4
qJnsVyARvA8jN+HaIZc9k4a9qkRg0IfU1TN/cJphN+9keBPIWQxklcLyhF16k5Lfre/RbKf2CV6l
3DOn9GZ+Hi7xBLC5P7aFmCdxU5nlxU8HY+nq6Nz2775noLHdus6ngC9w+Bi73efJD4Vg82k/n60L
rDkjsJOIVDVGv7zECLREckeJdVAaELyLfn81KUk60IL3NloKBZ/eyhhO11BquF62r6fqIhwOzFL3
T6rg4Vr2o1dVWx0xa/sL7Rno++TbHcl3RHsxD8gAxypxwAgVzvTBufo/0tYX+QF7o5eT5C6iZoZR
KQW3jJlvX97KMG0A5iKkEy/Q2PagQn8Q3ENXOTbidxN0KANb+LniTdGReIc3L5Q1fhzQU7+EpUiA
Anw0gFhqWfsLybOgj5QrrAxnQ/8nTHrxHmT3HxeWH9nxcDV+BFZPIJhhfCoCCyUvQJbVbutwl7vN
RjXU2pVBxPrUGwcfPhCriodXadxW26TCIgwDAelZX2sELxiDHKEvGdr4s5h4fQOW0bQ5mWEGjBKb
dd0sC/nzAlEq75q0GLGZMsXtRGDTiBMMwhK/R4ftypx6eA2QEO/Y+XAEb3YBjQX2tBt4gcgsAo85
jJb4OkZX/LEinVcddyVslVmqrLEUkgHwyj34SJlSSYCeRFqvjN5L2kWNbVuOl5DLginuEZ5k3DRT
D0R+BvcP2AkVd8S+ixrodQVMA9KZw4/hSLuQoQ/IZuGf3uKQbj9bIE84mysxXKpwqjbPYG0xpdQA
XxOj/yvpgCkaRr8k49nbdiX755N/WSiwrtRaZHf7A/slpn3MXEShefGI/cOGCOrkGmge/3dz8qPV
C1/OKH9vhrBE4VDi8UPbWrbieXCn8uZjZ4QntUsEZAs1e6hIPlnmRrp0Ydc+YgmVaG1+cvlBJ2LT
1WHuOCQXuxoUsWpRDWb7UVT16dOJp0BnGwALtUccwvAlg0NZNAxZUR/oEDvSyvDjWqtPNi2JYAr4
61Njj7vtsn3IkY3cGQQW2Sw3RgSMoN4NRy/npqgzWpxfCKBTg8GIoLsjmCJaknVnt0Vv1aRrL+Z1
CJ4ia8qiYRxqCTDpMUslPTlakqOQNk/kdmSGdestlAPokbGuZ6tbidEnUdhxtTBXCfunJCySpGlA
76LKzKBTaWnmGr4jmswBNtzDE4CfYaWwoJSNJ7QlNtkTaccZ3lSpzUY4HXRmjsOdgzNLeBV0LQdq
nuvov5zKElnbgVHmBPMy3XlFR3Vgmq42C3mV+UeSUUrdji96nE3dY4ZVCBDWII9LmCNeRUmTulRD
cIBftdI4JBgNj/cuhtik9T7bvXZ6Zqd63+TtKF297H7LZl75PTqNThJZtc2l8LMaXnTvfcXcq+lB
QG8Z1r6gLr0b8K8vtv0JyaOW9JSboEBevZ97Kbm5sC6Iw8/RgELB5qFPUCaTcgo+QqyJBHwiXlm2
h7jCXv+5DIrseRlJ1NRoQ5k+D83TaOGzJ3ljOgKc9k7FBJ8aiN8z9FIYLBteaQYSPNbQgJDKFRYv
FCCgTKXTCvb3f86TjOg8JKM4Nu3eq9WtHq5bc1yP0ml1xXmejraka2oeUo3sQfg9U3PL6d+VPByU
3lWgRhJo0zH7Sxu8lE5ZXFbOJfBPeTq+yK9ELSyUtxAC9BwhHmBwdXdq+nfZElvhXQ2aRVsot0+j
yu3gwzxu7T/6triHOYuvpfNLGXllhokbvFuO2PVu/VGwYRHkgtXL8rclFaNTpNewdT7dhMIbzPr3
hLYedRWfM5G3NnXwxvTTtU7CbzCufZhtT6ZBq4VQVgiRbHvklw85bxBbwZ0/DeGmXjFdr6jRSHNg
oni0rLGUHyjIUYSSBOKYioGbXCvFa32IuKs1PSAKaQbG+eklQenbpynd2EUhnYjV+AZvpM8NvBOn
kbEMVeKG6BShKH3E44lUyBpuwI6NLN9nhTlUi//p2AqRDY/o/07XLIvpTJ0XWMvOrB61KOrpfa0H
PVPVYv54fOp7JlF/W6ZTJ7fLFHWvThpeaP15oLnP1/obfd8u4IHQ8CJN+gaeKqa5l57T+8wDkLGQ
ZtyzJXQ8b0fnCnuuSz/6re2jbR9X2Q9jtwchCb8wIVyoX4NWXOwgljhQE/ECHSLHGWyVlQBoqOeH
5m43Mhbnt6AQUQPFjwrqhsmOnv2NiH1Z7DGZ/Lwp5FQAel1BnyWtTO8PfxGNQmOUNSLyVDNO4qDi
7M14PBgflL0MLW/Hd/rLGa/JoYSgOFCT59MeksOeVEAzDnINgRhwtUGe9au1GiDcfRmyc0WZnZ6j
Al81/un+Lixqhx+bvJxF6p3VgkDDD/wn+zljXAJiSEEuU25VBht9RkOrouenJhe6+viAEv5H9Vtw
XfvWvuWl8x1sUO9gKCqnsjlkux57CfQKb4xvUv4yQG1SZwIh5SA2LBFcuobEuelA1X9/wDn09hEz
ben7JhftMyot5uhK1ngslqpmmBamGEpDusSi7lgDec9ymH1wx7DwdXuxl6JPkPRZwoHhdG6kWKY/
7PrCeHbeNIC7wgg00WoDOmeA4+dLoREILE7z2gT/ENiX3rT5VVRHAxBeZjzihbiJ7onQXGfz/ZH0
O1U/Y1ntf2TH4waY4X2hEgoQn0ZXv+YgkC/tOegtKQIstifMBWYzhhqPf4G6SL10BHGImQ3Ir+VT
qmlppt6dmk7caVxhpilA80BMYcp/k9HVord7wLtff8Lrty8+U+sLN5z0QXnD6Jga+ombHEyW7rXs
1cdd+gcaSjvHAXS7/rhdJgbJZUOT3Kp3xqDzk40epBX97r/9d9ALaULCS4jzjzy9H75xBGK6SqPU
FAf2qYv9YZIuBQQgx9Kj0BoPMRfhf73lze9NJurCarH9WdwoPkqpluGCpPzztWd4ge//MEui6cLD
M4a5zx0FM7b83onIGsRys5XNNijbDJ6W0V/jqKiOnfI0Rq1UPjy5wQ/0ABkzXcuYI8qW7SmCp6kY
LBpV32JTHyoiTng+pTd4oLetgZM6jlgCzI+xxW5j0Loz0GpkINuyDcl81C6tnNdFcsi5mD19fDND
OBoRBBqQwJ9AAfUOjtS29m1+LvDDPc1RJC1rblKwZg4vkmSvEWVsa6s2OgWEKFGCTCyo5Cuotmj6
qsHskRJfh/dIb0ITfRj69y2GJAWtREHwKOjoZEJcGk8OLTNKoS2pd03AmU51TnRUJNh0SxcxByHm
Q5HWuGqt45QdfmvazKIzxg751KtpDRFpxcY8jABYqgTQcllnD0GWiTNt1OFG207o+lkORrspVtjA
PeoxfujwpNNNe+cVf6LLql+2cCRef2yMQMIQKWT/S7o8pJmMlAggA6/NSiy5+o4s6qT10O4cbrvN
kxX2vowuSZ5pCQBj6YH60TXAVLTMDAUDhKpZQ38mgQLEzrpFWSDxvjmJ96n1VDby4FXb+R/GmwcZ
1DWUySX/E2jm8vS8qzVMy23TLLwsZoHJQe32a7dEZ4+yRBv+PWfGQhlLY0KW5nlh84KRyhhLN0ce
ZzxpjFuKwz+wTbbrrVaaLb0HOjInp0Qr7yIamQYEZA84giYXOW8KS1tbcByfUIokYsltgHac6sjy
rfQ+0YESc6V4e9pLZoqFQHgLWtDw/DNtQTktI2m8VdnTM9nFYwMahPngFvrC2fHCMgmWaQNjky35
Egc6556u70KLVZPfSSKfv4cDAEkLa2yUsB2bKSieyvS7YhbJrFLfYGlVU+U4g0i23TTC4c6pzy5+
6dZnBE+pGpDAR/a7reY+mzdSNNnhsNxXsxyoaxqHDY3YaPBdrcRPgkWmL1weCxt/P0QqL3053rnN
BhwFTsmPikT1Fjb/RBEaYs92EE5oZg5X6RkTNoTYmidH9665mXm0cFta8R+zOW8dBTshzyvAKPiz
H5X+5xbTC5DnwfAkGK+vxk4qNyZazv3wS9GzzYIW9MsKjcCuP9u1d8/pqMnKAJqlJsLfGLvQ/ti3
dLunQeIPmy3+CTk02n/ShZr7C6toTdRLfJ+xod0UtYnhSyJCTjp7vyMVjef8tT+vlGZVRllRW14z
UCaqYykHnRNcXTMv1ZgAZ/ROTlJ4szAlTay/unOyjQSIm4PZEGm4ongN0k29hr1UiAnm26NoO6g0
Nn91IVkozh0OHTWOBAcBORClW0Fc85cuufVceu74TWW/Q8xwWgc26p6vGa/tb9syJt/6wRORbkAX
lL3pD+9Sp5K0cyEBV3IPx/ytPNcPymSAjswu99Uh9wYXgsDaR2DWgo5lgUzw6zUIwWG27JPsVKkv
O4BIERM1I/yjQbSs7raYRgQEpl+sIDIkim+UHzMin9HAM2He8OQ1EXodm58uK9UtAJrPzNHT01Vn
/IxG+uGhHpI+Zs+J2diZ/EVcW3KH/i9sA7f14vg5WxCkUvey9Jf/iAmw01+4ieL1OSuMpQJzNx4o
riGoZx6W9xtjO3U5UYEd0Rc162lHiHUboi3mRq+dNJSM8M+mild3Fc6IkiTB9SZCF6AWE/vrU27u
PMYEbcyX9CiIhl10JChC/AHASdKGvVC4Y88V1D+F8aIz70aOMbBYyCiQt+P7GhaV1HZxctEtBNWl
2BdOZVZ5cevZgUeB3Q/AUijnw8SrGOEwIa8P7k7ZiI6jGlnmDLKqkprnKk3+JsLiLgk2Mbr5wVsq
NHnWkRXg7FMIXau3o4I+6v1gadKWcztP8kAcEsDVf4HeS5Z6pSDadkx56+tprJYcbMo+HU7Pj6Lg
tpZc4QZN9XSw8Ctnpnb9XBkSvAC+AEUfudPb2QgpkTDiylaaahcZXUDbsSAWkel9Cy1iS0UDblfn
FyUD6G98/VU/ZGkmFA39Vz4z9V0hpR6Ca5rfJ4KqAZqmYwQCnGNidwmFECgL05MBAZPh9MRFuF69
8R3iiQ9vJhqATA2yJQbEBHUwVhstXZE/brQZK6GbOwlec8eFGmjqdJkJ0mX8UMsNrIvOh1XHC5IW
T8dNu6PXTfjpuQhcBDAcU+VnQOr9eWw1tvCUAuDs/AnWkXpamhJ+srE8vNcp0LMqvER1/+J63DdR
+U1JqyN3QBEXa8DpWgqIT67hxExiKXHXbC8VsJTwpTVSAh3Srjw4pwT0yklCPEL4JQU53k5kNV+V
9mzrKCzkGghpNJNUK1gdhVI3cJgWea4IdtvvS7ibydEhLK8p8KGtm5sv1tO2eBHnkd9XT4CRp5Ki
UpaynkWOPrNcOXmYETWYX3EH4s41U8J6Vw7CdYMduSQP5qnLFA/DDkCxQnJKIbyfz7nZ1ug2hNMc
ERFrSXxDiGYs/aE9IZvaunQKmhkdk+EUWG+/zFZTyz+8YudeOMKTagyZvRu10Z0o6ML28jX34nVB
w4KwCv9mZpvSnLZ0hyV7vGWfpNMLR4glUmfKbVwpGHbiK+TEZBHtTK2vEow7TcoI/N+k1jx4jMvv
OTrSW/C7leTOSVXwv9Al2kmbyguWQQvFZu/SsoFkXzS8U2S5+SSWijEUSqx2GhC8VGEYPLrhcmVL
LCGdcdWQ4q7DOe/U+D6hChQNiYxeBIWK3EkmhhdsVgYtDrtPWAnbP5OIke86mCGDvyiNarr0QQxm
cZPDKQzgBwm0uhESollojd3Hwe8PH1W4+pp8pYbp4nkNWegZO7vykEIGbAGtbqqR0nCHI3EK1bgA
y0lbNXsfQ0FYOxgvh98YjSkR7Qv9QmmWSxzxgSYptBfrdT17Jk1U7lZLsRdU8HRG0uumWhjbfbit
vIjBARY2EVpQPjbAWP3EA5zTvwFgUo+jwHqlQmnc3loV3pPWMqeAgyM+2WAuCFoupTJmNL+U/Rj+
gc+NXUzjbV/T0/FI4Vm092/EKc26nvHO5T7p1ui5idiXrR2EHezB3h6OhlvvFKGT+yCucrlyWd5C
3Fu1/7Hn0AK/TqX3cjvA4pWt9f8JGB9XhjCUA44sVkMm3E82oCwEpNH3VnkNICRjMqoarY6aK0rr
ewb6vbzwybKlUwUivnrsFVGwkySEta9YTDL2G0WbDfGZwNwgkg/vOyCb5N3nRtIUXms+rw9N5FZp
Vh3g3gChrYQua+Y8yWwuCRIQMII26Q/0HJDz6nXziPlz0rY6sxbwAbtpvI1wXicNAD8XGfGij+P/
mclJAVnkpYtqI+lnfmRlwal/TI3h+OEP4iaqNrhfalSoJosuYgMV/EfzMmBBsmIkp8+6syeBTqSu
HmiJSihAK7g1lZv4qsEOq8hDvXzXbpf+2mN7egZRIO0vCLhndwuCGZiMksrTdrup2eoNip1PHHh8
9t9/3Q6VLQwMpDOUXzId8/qf5MhIVaUV4ryS9Wa9tS/+HmnOcAcMXYvJI3pmXhd2CIJrfQ2jHm9A
XEHXwsiG33dlKnovR9M1YRMOLFde1yZCMbeB0jV7Bs8OmlyPuqrPz+sOUMOaAYjc+My5pJ1ZT5Q6
LoebPDfCurBGlQ6n56qR+SEOWzceEb3GsWybnOzBmBYwy62TAMMpD3xQBD1EMep74JupsoVeroW5
sZjSMx4YPv1uMXcEgcRAwdj66jaPwoTCz+wHpo+abE4wanVR3Rum/reQGHc8Ze3Sc5+nj8t1jUwL
QuoiNUb3B4mOXfwexkKJP23IOBVG0iDuxsM1TetYs9L+BwAiPAXZ7inNiGlrAu1jwmblaMA+USt6
2ZsTBkJmG/3duHDE4ibI0tia6yJlEgxpf0hfQkN+L1kK7XlpcxpeX+KjGMP/E8C4cRNHgUX7E8AW
yrewKVdiNXsQxZK/3yJBfiwuWasaFNwV0Fx81Ol1+gqtHxVHJTi5OfTej60cD+NJdIbRQX6NH9D+
PKjeczCMExDifBhO1eQ7kvWWW3XoN9W4Rdb3yyzpbO3EfTKy4xf3eTs5tBGgbZHL5OYgvfehLi3n
IusRerJCMcTkQ2cAPIix4AeDWZ0R+BPAvulE4c8goxwW10OsEA+ZxhSz0hY+wyi3ySOMEY2Mb+nT
MjLIrKCUCOmIFPA3Vf7PCWSfvqlpYmUyHHkY9e/BZCliOr2iuxg/5/U2dMIWkCUetqbBhiEw0ZkA
Qy/XcvHzbWEwhghSTzC/y7qQ+4WS5ZUaQCMQwkL56Io42uXTOh/Ll4Mf52yMUx67sN/mgPEesxdV
SwY5XL+nCRqOd+GQEAECUsGS0z09E4P1UDNsZvybn0F/2stkYMYa+mtunn7a7lG58nAZXHL6OPBm
W+CM7F55pw4RJaGDkRtK2HgJqkxOIC1zOxneG6ilflANZ910acjByeF6vSlZ8ZWfTe5ZDgnmkuqi
iuuMWdB+BlmaIV8Om8PW+XueHMV/tPdj7PchlQ2EJnuyI82OR4onx8njYKGQEQkN311Xs2K471Gh
4QmctxWOmyhjjsoEILfuUJFDhMQvbZkKd7xf/7PUmIhFez55GJFJIMFzPomtOcXJ3a/7oM/MWUcc
DG/wCJ2S9m0ss1dKq5hN1pni/w1PNbdjdbu8O9pXB3d4PiRKUrh5favtCm5m3LTuKDc2fd77YPbh
eqsVWrsHKtwKAOJj8WHTbCoBRtKvkPttVow2IRmKXvvX2HhHmvTurV7CJaIUteZK4ZC6HTywPw6z
biDO55ssLHg3VXlJbiPaf3SOu0v6sHp8AxW5T8H6q8wJaG2elOJlRoKBi2BweWFrGhrySJFL3OTH
foPizjgSHkX6Mb15fygvTNpZb8dUSI5KCzE6xipXwBKOUSC0vc0s1uWiV5VtzqSwx9R4ONQ93+iN
KyQrzL52/TTUo9JRJ+F6DsjE81tDNA+McWI7y1BG30voJctuOJzwArJjqDMwPPVR+31d2X/729eF
ZDMqWon53BSv4SSaKFkNFFAO0k460mHgM2r4u9fuN5X7CgOh7ByqKJphhaHS4C+yzDkecMGZpQp3
U3LCVt4sprXQRufs6VES0ZW1uGR8ZRCHSNh5stHcTbQcctzWNOP1HqYJqfmKiIlRQZgMWycVZ98+
Gl/cmVmx2oG3VrGxnxuIga/gNuQys/kKC0Y279GDoovjA77mgXRQHz7iBhlV293fIDz6VRJrR3eS
ftgXWfZ9EIxCXJalocYusllRwaM4RoFjsN2aEWvYC5AOw2CuRIi7cZkaSdL77ggbn5dwYBBu8GpB
hqPsq3SjJj/BPlBB76ZlEmWA8UgwE49y1Am0/6pqboY9c9aHf6ZiXMRclJpGpHqVFSe0I/lPsryP
caXYXMVBQ93McbmgrplHsyBtRZVJxk8Plad9In3eThhjeL1xCLrIf2hRZjikVIpK6IyBdUs1JE4x
P35wzeaL+3oT0DhG859r6BsoF1fLP1dF3q1dOub6suImi7plkiWO2nQl+dwQhh7nOZAIFTx894MZ
dFLZ47uu6q69zLoYvghj0I7sqBx9PNXax3J4qTF2oSYICjy5XZqCLyeknyY7KeKDt/ypWxRA5Dju
vqxbnqkBzNaNN42cZvBD3NLzZnExwoAfx+jpTcpNu7xKhcXxzQ5STfFcdsEfoKOzOnoCnEYWPgy3
Sp91eYmGmmjyOpFEU0cHlZf9z2Ut7/QhgaQQtWaOq4LceJPmvd3E8JmqMnQNV1wwA8wfIvv7exFL
2V8+ktoeokS2EWdn2grmiMjKPMWoRcqm40FY3PUAXPJIcT16yrwzDmF9FmOt/ZBv40Z86iOESxWQ
0cSCqdrLi6L/0XpfcOd/0DUu3sThRiTnOjzdEFLfE5JWk3O+1DMLAVUhmKgErAFlveJQtkMRPkps
tM9uzeZnExOacuHmlTm/IGDFr73qF47dRQYok09ozKOIqzQdrkb9wuzK1q+kljRf3gtbNpRcWbN2
9+ZeFhkacJCQtfXpTr1lVJz4ewTfmV8rxWGiSLEEO3bwLMC9NrO50REknDI0R8nxTn/0GPJVWAR/
yOrK9L6rNJbY5oYA6SJYHwAhC5UgA3Nudv5jSz3z3/OYqLi3w4deGMOvqAuQHgshCiWmOlSlNtaB
7M4y8zfRF+fbulEpnM+bcsUuxx/gjuxfV30gT+parG/yCCs1LdjIiws3VH/PSl0jTzyOl9kkgwWY
4bu4YN/pqak+WdHGm+WiA1GCtQdnKofuIBBIeTVNon6jlfPezEIgZqOSDIdBtpM7kTbrs5OvOICK
qDJT+sQwJsQco+1weSRQHbSn1g9rNklqrkvjiLvyHc9VwmDpRhJdpn2Tv3/Y5fy5wQcyilhNmPxC
RekrKf3YbOFXatbCI5/pgPZpi2nCHjY6TF9a9OVQrfSPx/9prwHcAa9CVWTW+sdH2eYbcGc5TeoE
DNBeOKiObe38WRuRUU3Iu4XoR15VBIArZZ4SwnIPoKB0LkLU3n+oJyc3k8wUht+EN2/KMVgN3HJa
QPrCEyth/7YkmImiPcsG/LGbUkkDbwUlSCjCGXahjlE3wXR7zZ7ovXuuPF2LczdXgqztCdlQB37w
gZ0FBd2ksYYTUPHpU1EgQ/5w7HyhF4UoEh1/OaKhhVQ233ICLBnbY8z4kvHu1ufzZdXv5m7ZURIU
Qs7r5QvyTsXqI4U4osP7zx3oHeuKFuMImqTZDQovXJ+3FqjnST2+b8l4khqx6b22cGjMhCQZnoQy
/Y8uUNA5aHlD+MFVlxvYhmNPof4lBJKStTG4C3P/pe2QAePCpMTGZV8CQ8DKAP8M1IaV6uG28LQq
GPbEndREO223bgaFTVB2Yje1hwb7O5ZiHnPPeBoKG8nAsGgHpvq5naaEUUOummmOAfvhPOmcTBnb
VXo8xov0qvAuATXb5GVcES2sKOaroDXQvFflvloaQuTjwCWL14pIuFpUdNzR0aAe72SF7P9JtPk9
Wk7HdEHiwxDP+VMEz8lqJAQ2Az/zRDBtxgilvKFdMVeCQ5yqbMcmp0ILcL8jmso3TQRUXktabrPq
8pXto6KCstkeWAl8ARhTcZTvH2jpvxMd2QyAgQAi8wAv3l/GVfvudqmupyE5CCraCdn6UKeqQvv/
SX9PALHqOjpPdfSTq+7jeeIT2Zlxj543c2uhoG3UJXXE2WfniTCoYug5R8OLUhIDPsOLVzgieR0m
yq2NgsBpXKfUpM5OVj6AIsJguMM41XcECkrPxQYcf7PEGSmi5rI+3K8KlOMloYB0SXFlO2xWlehv
Goh+UKIDPkvf/Sy8jgi8PF1jFP50hF3G/VNaRaaFkdof68HTKFyTPrQ3htIP5EtqqTKRpdsPOi5B
Gu7XwOC0x/5vdf/ljc0MH/pnto9OuBOkkhNFlHhMtlJVLfsvTBUtTPkYbHxhOqwBksYLuIqLbCEZ
7rihZP613siNqeG3vee3+qr9lS0m9/wthtYVjqk0BpNxPqCPXTVtACIQ6HOVDx/0nFNQavjG3jMa
Xe1WuX8pS3KxgkaAkm3NbzS69QXbGvvEqV7QJbpS0wMF756L7dcdt1mkGKjzXHvuiFddheWJYZFT
qw4/ct7iOfVUeJGSjcEfE37W6Uc2lP0/u1ty3CoeSqj8d1uZc8klMsAyHG42RA6BepBHxsNHstVw
Uoc4TzLNtrV4Lgh18J7PcPDXaHz3h1yzsWf3rFfIaP8qGccEUkoSYPgtv9xEShPsN5Lfs1UNLXZU
4b/SprpN8PL0Ebgmd3VP7JhXyHret7Gd3146akvM1KSSAZB7ZV323eMusUH+wM7iAVumv7USqojv
cCD+LEjF4LL151A78oB69RI0VTvuVNS2YUJfRrR56aArIbjiEVMp4kjFXDXvNyWH+fVDnkQaWDKF
KuOsyOrwsMGllfgc647ztTubzPhAh7pzeiribCXt8i2NezWR+WaKgLMtULlvhArC92kTTSkWqVSv
g/bo9OjbmZEURbXzt1Eca0Osl6ssBCj0YMpxcI+tngwpzHVA44z1hfQ2mXjiaYqHzvtyhB397/wt
cUtFW/rCC9wiDiLO5C2XBI+L0dJjPWUzamSVz171AGTLDshO26d2wUd9DAJM9wlAzZzIv+e6SmTv
9FXWhipNM47XxIXU45ix2OyKtzGNcR9p6yiorQAl7O/9bVECPfmQ9HTN7Dh0XbCqebG76ZmBUZDk
Sg27Le/2jvOcr3vnCB0pGlKVH1DCco0GoHt5hGdPCoANiNSQVvwXFUutJ6pRbw+pW20iD/wfv3cS
HZr+qO29JxHsiro8F3unASVlk8utAgGWdG5NmMnVCzsH6qZW/+lUPPxaeezvNzP9Yzykp3Do87YR
rTeW18iGbrkhrqXdvF0NDm9EPwvHF63+ETbBFlgrRkEkn4eH9sPm+qXb+O1MNtY/0/6sn+eBhJRo
H++bnOQwxRkS/DLL9qioIMjKlMGDWaDzIN0Vmf7XJrjFGwgYjx4+8vb+MVBGBgocfC7wGfG+THS0
o8WIGab75Y/+4ormTckX34xRfcoOta0MtqckUgHdi42xLjbKbIG5YQhAPpHpBk6dA1+RFUYtJPZN
O7CTZ+MrT546Ngqze2rLClbYGc1qurNzuM1CQsDACcHkzKcYncemHaFkYJiFuOEQsI51ZPDUKBv4
O0xJtPWT4bLAbl96SZrAof2Sno5r6mazNV5eKM8q9dAm99AFagw3iOnt2+3eTcWs5RFDlBHsF/vL
DzH1TzUSB2276IPwR5O+yxvIxPioDXP2xKC+FVDt72RFL4IwbN+rCcv9yQX+y7c7sHGSX4STQ+eN
Ke1mK1P1GtODdhdkYIstGEkH1GsrcWwD+2JN++VB4C0q2BJMYbbFfigl4wOyQg5A5S6XUud/crIW
V7CTaYiL8yhuzVfggBFoaWHpU5jDxh4Ysy/YSLutADrpWf6kfdnRwXc1cdJdD8Qye1tolt0MYuzx
lBNUb49yL0XvprmQnK82+C43omrgwEIb741nykYB0K29U8FhvO99deqn8Yx9ZI+QpGM6SPEYA8Jk
hEKqof2JJ4+XMgsEmfmY0R4Zfb9XBUkGCXV6LV32daJ8vHzBWvdT21vAPbIiqcra6872ybY1VI2E
2zuoHDOrEIeQGznLYtsbi9w02w1s95E7q1AFVt1WeloQUXZ/37R2mP6a4s06HxnMN4R4ptn1QtsE
dHEbJ/omZgrv6unxpJvpE3T1RWPpwY5TfO7fExGawvxXY5enL49uxf599ZUIVu1PxWuYiWyk3IEI
OhEcmr+98qMVQioEhSVVg1VkHb4UFSw/oVPNxFhOsIigVTnN8uKdWHUelXkEn7edhVY0CPwgo4ay
1EWURjSGiTXirw9oRRfShideiZNbrRTe/XSKH6CTdH7P0NHHcf9bFtcTDR+kGhMt7QyxWQQTHdZr
DelE2Y62/x4rz0v8oMmmPuoM1Jmh0mCK213I7vNonRgdTB6lmJ6ebEVplAjd3Uzf05rn60/NZeos
9SrrgdYHNXlQdYLgz3oembaJUBeiZ/et+VF+lgj4ky5/1c7NFf20i0EMJ3Dmg7nsxC3UWQTGiqn5
ErXwR7E/6DH0b2vSSFmvV9yGavj3RuoZhe85VCz7GETEbb7yTpHtyLOHj3KWngj3Ooo1FbalODxS
kYsiGuV0GswoYbVJbmsn7w4auJDxnDIkBzQqfyLthR82nbetkGHvQKIorGEcJ+y9UliIYa6c5tDn
xrjeL8UgCoZ9FklozMDpcw/Csoywhenn273JHr3rOdhg4ccohHmp/pHgEPWlK5b17iNb7IyrmI4a
hAS2cY2pMHqwdR19aq52NgagUctsVnakQ4101kEQC1u/bNEQK2SJ0/cB1TJW2HofUss+IDG8JWUS
+ZMyzUiMvalvSQHrVB+mq9yYHUitjq/lCSJRzaGki94dmYNEvn9fd7eribZyEhy+8ClD5vcx1bBy
gDILMunmGNofavP7cquVc7JjtyYdyK6qePeU9k7dngk4aCnYwxHtffecR8PLQEEKdeQW6By/PuBw
3vcceJapsBhvMfYCUVgpl88B/AT7ZVojX5o/TAGcJXrNT537j1RIkwnN/zkmBdYFzomgo1A1sdc8
JG+S1X/Wn2UiN8JKGpVxc9oBm0gSW4vcGZZdWF/+tKMNcPYW2jksKrqfCXBDDlSbIq7LaLNt4mfB
0WPVrbTxRP3pwpeLCgUvszxxxYh4aS3jH+djWBMVNmiP5N3LT9dl8Ibbc/wSl+DjdgLpBq458ffW
RlFeR8FpCoUyxXoNmR9iX39bI/kkcNEnmVmzelx2bN45wgphy8aTFVv59OpURHupQPGgicxxDPqR
TNCk98KGKOd7F8vajVGwdgm4H/LUKcgmWwmGOmnUlI518NVjy/cnciaFZONEWAdVrjwbRybHh5LB
qYmn0pu0wzI9L5HqrN7Ucvavfl01ozbxwLD7jvkUtpCzuJyi5ZQqO4c6pGPdmeWGMWTnV53AlL+q
doBJJAsI1Ij6FQ2nNQ3JQvVrKymGHTkU2U09ilFBLeHp8zzyOx5pkymAckaf8ur0YHNhAvbLW4Cf
SjQ4gQaOMho/+bhehAX5BdpCa9AXy8ES9OZbamPSHSIuFyHN4BlMm21InN5W1H9K0FiueDhJq9fV
qy9OQlOd8Xuyg6Z1KR50YVhd6hHzOn0IdRdcPL4KUFuxNQEerlkvPeSZBhGuWeR0o1NuncdOG3CI
sNk0vAojFg6b3NgAsBt0xskxt2lhSmKpdg332ml+lRHT3FSL1Rk7UsLeHexM7ptXnvQUMIQPaA/Y
1IxxsE3Pt08Kb3PMgSBjWyqyC+58iZWM61Lxpo025rM+Q732PUO2dN8vKqmbCeA1yEBneahDrEk5
Szw6XWpBABiCa5Y9pAsJvWX5+HAWWDZ2NGF0AQKQloAtki2D65aZ82nimYUQO7E+VJBvxKdPt4Wk
y7LJgUjQYDv8ovtw24mz6N/U/gXHzOgwLWqxVt+/CzqewHSsq+EK+pxaHlMDajF88Rk4VN6bAAj+
MgUJVE/1kVqZcQ0MX/YqEgqdla5RRWErpa5BbyOrqLOZsL9srcNvgC92HxFvopDb+DtTacEY8o6i
XpH6/H8sl38I7267Haa/92QA4e02eHeQBGgyPyRxTuMrO63wEYTOmMVIvler/LFgHmIDBfRcdCXE
Ho2CIcg/D1A2PQZ55rnZr5ItH/0e1fUbmkKofZlLK1hsoS6Fb3ib3I7TcNDoQeadMZkfMx1ieko+
EUlGGoh2zVNsdMotmjzYxuhThudodelZ2C50uGDSdd3T0NaOYS/C7/qRbqC9C4gfFBE9B/+0sXQM
sSXYOX+aPzDtoAyc3ddwuoIeezDh8MRNcGwHDEdA572tOd7ys2qUB/7UjBLswvSv4iZl+OUlFoFS
p6EaSs64LMXAANkCned9AhLoiWamf675Njhc1eS68Jf5JOa5wGDdR77f7KPQvZ6wrHS02H7Sj/13
WnruYJ0n54oykGxtWy1hagbCKFDsSblSgFo6bxT9AUkFMOTaz/37WBIawMUnEO1LV1+C1JvzJvE0
KkNYlORWe2Bh8uoHU2j6zDAtpx2KhsoKr8w+T4aaWxaE47KZq498J47EYhrzlMxR3Q7mVtGw1TKd
uLEwef8bIXn0o+iU0hy36A0V1p9jLwKVpCW1hmi7FoK8iOqR5xsqDTK2gTxjcM3YCOXcyuENoN8u
ZhzwN8ynY/JEPafHR1fzowbn9wsB/tVtfue2HDdB7x2MUn6B9OoLzl451drVjNA8D0gplyJ8brg8
9rZeuuH9buqj91RKyyGytMTzPWAp0kjt0IAOJrb/t9/hiLTlXNvi/weMMlMqldN8XF7Olmj75rRE
wAj5mWTChmIIlcg7wRIC/k59NsK5lpVh85La3ZzTGnRFxYckkWMhPY8qNwY1VEGhBTUHzIgpnwux
nAT0i1CVEDq16DV2OU1cRQrvVxZ7F5TUf+84GF67WO439wjnXsEn+xUxLy2mddwvcdwpp6qT7Ok1
DTaiOHxVYIs64pHU6QYxhYcq/Lo1jItXYwvOc4dtwMdbJ0P8ruBUne0eidwKeXfcha77Mw+LF5B8
W2bAbh01OPRSRx0ehlRD6Ib5yiicB7m/egBScJsb+7km7syGN7bh1MBaJOnvbd1AQFdeVHkYsqjr
TsEquaNEUCgVrbUA3p1nbjgoLEry65Vbr3Cetpcj9bc1lW4peVfmyD9qOdRLhkzbgsR0ATK8MVNN
jf28zj70yLvWeJUYJKGou9f/XXnMGQgFCwncYGKmyvDW/r0ingQiz6OE4YZ3yQXRXX6TYvryiTfD
RZ7WvC/pV+YQvobCuOjSg20Qat3SlIdoiVKOwEMEYqunzXQJAvrHnIK7j5/wuJJv+ourEGFT2Z9Y
LYLvq9fqPVcANFKRknTrVSLnp6TmegO66o5AnuM0SiFOhE7tR0oodgSpeXkhUTgLVmhzGvT60aKA
Px+RAUcnKcAOdhnVYXqBesIdiftMdI+icoF9Aroga876phXL4Y59iIKfsNN/vRGLFF25e/IFw8Hs
hLoNk2p+I5T+zFSrlRD7+oDQpmqDq1z8XCAxzY7MIIlw7wpOBjpaXXTrBZuCl8LFk727zEUobjOg
ro0vpSNNMaGyzfJ0Xg+vTVE3VUh5uYTkS6nBhkFFpGEOcous08uLeDMHCZAXdSAbDDANI/FRmGEO
7Ei4RHhwqzAQYSbgL8kERp3BHWsqE2A/etWxmivkAduDM13MQVAQzEpOTG5KvQOMKWCTyYAZKG6l
iOLWi65Ye4rmVdVm+GAY6W6q+CU5G08RisGEjYL8WS8XAOyX//U32q73nJYRyFy5JWmYp6XkT8U0
nfU8nN8LPCK+RRRsVzTcBTm7d0Hj8GzDrymlONR6ej1NY2FBhNsHDZvMsKdzAjiOBqL/tCIhi2kE
xuYcqNUbnVZSzH9tcIVZOZR8mJD8hKNlGdoQVCUk4mKnvzNRdqdRwNXTDbLA+0gDgJ9WVvPrrnfR
mX4r7gSVwZ7e6k+bk8vFlzkIds3N4nXuDYrYxzKVC8443pe2R2DLe1ed9Z6hUb9h7bbn8J6Pq2R/
YUjzMfGDQ081K2ZFIzXNacbc6vX11ka1066qqCRl2cj9bxnJcxmoVLpWO7l2UUVYCRJEc28aBKfR
H+ab48Cj6n12vKJ1uon1jr0NCDszVUBXrrHuhqo1aKiIuK86acYelXwk1xZII438tzIjzRvmfcma
HbCNqerwE6EBVVGMCgdoimkr3G4dqJHkj85nBtwzAGcU8FIftlpLELVDVS6lxqs+TiMdDa6rPKOJ
dSYm2iHpyIO08YYlS/zAOEIKLCT3mL4h/XXT/DsxdXVAO1mWyYux/kHztUOmXkVBvON+WTXVoOq0
/JGIx/Qy9XdIa8QyPuMOlYf+ftLPCnKN2oiA37RrJG6Mhrxl7oHKX4wXnn+R7Z0OwcsAYUWolWex
fkn6MI68OklZ+7mlLrRrBfnPxgzS0JgbbPPZkMPUCFRCdoxwCYxpWwDFge2pKtpY0gD9sCT2pYgp
bY0RI8cHTHBu05KUU1l9PzL16pinoURqiMqn8/0aWAjaVeIEM7/XgdWSujjPWSdadXs1bvL++/yu
Wuz9E7iQrxraSGnMuCgIgNd8MAx81r8keccdP4M2/xMuNNcWP0AuEiYpa1nqbPTuDu5sa+fI2zej
MT4Du2QShWTWD9eqG/FiXENygAE0+UhBDLaIENr2s/3OrAktlfpLdOC1EtqH5dYtoRm+Vi9o21Uc
9OD7hOj9x7WiftfocVhrkp/GbgYomIuOwmZUJa6zSmz9Y52fD6sOF57UNFrikfqm4a3WyGnv7bG7
2QtjOhsR8LTQI3EuFcOzKk7clyeLp9bXOlbHazruTPu1VgjAEuevCjgPXi4S+SJ2lHaR+gPoZ8eg
yVP0aM5+xq9m2u7STXHNgImg1wM8Q5c2xup5C4l/rPamkTndYHJy0JCKI5k6qopQWwra4+9iak1i
O52zc9y9pvoSikRhY0OU6Jo9n8XcbifohqZffAZ28C+3xj2ZSrHXiwDSYWn5N30Yc+n5k1N1xAZ2
YPgbGpeQL/JjoiZ8d3kNGQXLq4f5fhAgGQ28YweLSs/s9qsYk+R6mrKJ+XlpYPnr2mJpNadxYchc
rQoAiRFQa7H5X1k1VoNcRlPjt0C1EfWfQddFYTWgMQ9HN7VC2lD/F2T0qXSqob5QKt2dAjqVeygf
rKMgbBNINsQ1dK/pfbdnb1/8ocyowdC7FjJXDn/OJGLVITHbM5pTBauBUAsJU58zj+Y+t4R26zY4
62orcXED/a0x91ZDZlhAzK7lyJgP9tdeFjzO9f6kJQM3w0lpmExaT8N5AaVe4Jgg5d+VxZs5yfk6
A7pBnl95aIfb4scghO0V3r3k+tjFKhJGFAFUtbuvyWJGzaPh9itM6i4mM7PjwfoUAvihY+WLNGDK
knjY19yrqefJW6/TIGCSB8FjuSkgVExdR8+nCwObB7rWpcaIKrVn7xqyo4dntoXknG/vwNZTDs42
GFN2LUcEuLOwJFVj+DZwjkR1Q7/PYPDm2dogya3phSj4kugXL0UGSc6la2zOKjnOm3aabNNQ4faR
mQruAFrdcqTA1Mdx1RHF6Xt21ForJk2jcsk5RQD/qacDJaMABHvI6yLuDiucUY+vrtw0FbCROuQg
vZj9LsHR5Tgv3ZGpySBV3Fpt/DWDXIKb0J5q0vf5Hcvh31+7clN4mSQvSklhzfcvACaYfV8Yw24g
3zizHfWsyDsySTl5zEbL/V2uVbmj9U99w4soeiiXp0Ki5dxggeB2tf/mORz+U/ec4WExE4dq4OpM
NTjX7C6rY8O0Tr4CNv7ffR+n92F57iB7S+LriKbfC8sZzKmJ1wzoyNiAAHGTKVWqj/MXSCj+HL7A
0iKT6pMt+Cccl4hwasAFZgy4KtvTElJP0gkU4/Ugw9OWmUDUkHRwzEEgmmyO+97l0kpldUTOaruS
u24EiylR3D5jMlkX57OFRmst/d8SaxFUKYq7a3bh9V0R3gFx33Or2GJOYJl5oFVcSY6YxXHDquzo
MsYrlcyBEqf83PcN2St5+RmXG+TiahXvzEppHsVtisDVZZmkZAAxH/Vi4M27lE1xH14hVOpbCLP7
tTYMBqbUt0QvQNgarrFOWN/Z2OKyecki8C6Pj4I4g4A4F8IJKwcuNyLYdGLubT8yilz7Hm3mNBtr
DpPjmpxSxToXsMcE6E38BRU7qschVgxS7Zsnzf7Nza0EWZ8q72NO3ciJG/fSlAOSA4/pDYQKUiS4
q/h1dFK3JQpRAWHgly7NQQnRQT1fPnAPcKcWrmXfKehN5iW8YwxMMrD8bwQogsxQaUoW3t2IW3o4
PdkoLHzIjW1+AutKJmRDg45drifRsH9BFN/Q0F5gF5PrczYRvV6DTyFDAvARw42uBHs7eLa+nPfA
ghB+CPPuHle6VxPoyw39CYg6DuPgKyWK+KIUR9JBu5deUSwKQpJxx1wpY7mKT5/G8gPUlP5WWbhI
Q8N7gMEzJQW/kchn5vpyd+zRMOBRSYjpGgARKo1XhN9OL4kYIpGj+v0ham1HqxcxEAOmRhtsUm2F
hNFdw6Cz5/q892kEFXNHzAEfUQoIqpvomiUPhqqPSiAfMyedoBiVYkeA3Zxz7sBr2HVbWwv9cO3Q
IzjxhmpGQlqjTQ/BKWua6LBC2ohdZM0yixn2YfUNTg362QP7KgHg/v73peZl5mEzoWTnX+xvMJCD
JILmPkNEM4APXeX+ujH7y/Gqu6wCksPD5KjZFPfyNlaJVaLJxdDSfdonaH7U1jDKnW1iGm3QeCfK
NMaapToK7FoP07/xekkRhym/dUbQtg0o+Z336GPElPkBAA0yqM+oED383OidzIg4U6txDvY/KUWM
zstrMA8PaInSgtwoF4bRSX8YP52dsg+sOVa4aQc+bwSuZYMEO2XLPMOHJM3yTMsDASgR6bkXElS3
6SMxi9VVW+7MmJmOs1Y3khQy4lPcAFYB8Lhwhak255CnC0cH0W59wQC77gymCq8SgX5Ymk2Ofgdp
56+NBceAueTNSwvWP0QhuCoYKZpxLrBU5WbeCNQSBtfn9Ys0QwNTIzSYe8P8j9YXXCd4NSWL7xAa
NZ+fZ1vXrl+exMvOgzZfHLrKec77dACf77DyKFX1c1O6KF5tJWSeXBouvCskFVrltNvyKYhsYsHl
iCHbWDx9qqCH/c+56O8vPR0HYmI6lx/1QzXZtUWU7yi4f4dgnYeLNuNLVBHyaUtu//bx1Az4zM2I
/FmhI0urpI5aXs6ydbMMqvWx5nkSJ5vi7uq4ptUojVnyuybtuzMy0u496hbbyqSOanB4moIcyhbD
i2/tm+WTHvz4t1TqIVDfV4EGGXxOtlf6O9VXgdW5//DszzbU0ynouC4+qqzzikyEeMaXDGumOy4k
tAtRHRKN7J/gw3UHNEk/ls1/CGjwSh+M19eQeaGLaaXEmLtwuCtLraImLYG83LpMPeqAb+KVWHSX
EGceOFVtSwRrrsdocmwExrsuWVLHjDhZueh4SJIfBeQh7RgvefuqZdPPcnpFcdlKRww+11iRt1MT
MmwUbm6gIZgXXxd0pB2WgXaFlI4OTD7tc2OF2/OasMucpulHeURyNL694WCwF+HVqNyAmKaBymsM
Mg2JTkZNGkvRlWEvs3T0kiaZzewA+7+kS2tFVOlc3T7u23nZxkBvBFW0R6d5uR5vcpHw5yNCQ+Dq
mALaTb9xnWw99VaDwNVpukyTkeJLnWmMp1KXGBwT+SmttVl0IY32Iqcuk3hyUYkSe8hB978Z3VbZ
zVghf6pujEu95dDG1yapXp6yrLmlltgby5u/qfLxSth4K2rNw1pakmK6Olm3rgAJYoYcBnjDlgcZ
NLoOynzG3kpThM4vzk2/KSZiBPyEGc/vZ6v9bvEyqFYfXKNH64bYfKJX2uMttJEo7RiXTYP43IAS
aDZLy/vuKc+w7jhPPYOorQWK+nmyhM6ULzVdQG88UM92SkS0X4xDLI5TbQOTBNELvSjDogLuIxyb
NJYcpR4oaXyoQaS7IL6qRAuBe8hU/zaZ9MbhrRfetj/PmkHiSQW1YNi7r02fcC5LYGfRIp0aqdsS
4NFFVSGcfasDyOYA3YoNiVSqZHK6ajgPpMugf/d7Ga9xZ1w7M6qjSbQEt8rKHhFgAHwJ3TkwrdE2
35PkcXJSV/d8+9OA4LM2LYBNIcRi3fHIOX+nxdRm9fmHpS8Br2/tYnA3TL8jjYAKPndc7xkmDCFk
T7yvOQ+WTUdyWoqHXFQ1C0HCVlE+5H+EJw087HQ7LcDP1oHQIgfyLdVy0GWssLtoP9zWHsfX89Iu
H2xJiJg+az+5hNclDBThvBk1mwgqlHrTK6CvBsT4stghYrcBUTFAVONu7oUdnB3Vk7vr1BPgD7OC
WFkEbQtsUO8DqsH+y1gnglOsGgr3atVg61dMNnFd5dgqYiInXGxg2A02ntk+MlQp9g9neR2Ne89K
WrqAPnIy+PzrUzclTE61yijvtOT8G7Ym+Sj0Qv9tr/gJ1VEr0ZblGtJ3UJaPCxBz9A2Fy2DdnDjp
CAURDNGaQkUSObLkdnVnptz8Xp3rgDVh7foNcm/J0r/1U6hDLZMlglxIIJa3uLL0Vvt0TJjfG9yf
IAKbgOhTvEe5rDiaUiV2DFkr9K55wjkhXL3baKR1Vb006dYatX/GxWJszrb6+ywkXuk1JlquxuYb
vegjlZ4r5+02whd8HAftUOD5GTS4oyzkVlqvNTqB0DCXG1aRprPOHicbcCGU/b/4YSmw3zs0o/Ty
GjK8GHDVRhcAD+3LTPG/SBgH0ivTwYN69eC4qpoojX0zOfEjn3dpS6hiIgH5TlKookDtQgSX0wKy
GIVfcrGc8kRqapwW9SwZiNX0CwvNXyvcvzwKKAD46656lovmgFOqp2Cb3hJz0Z13tfOeWcOBDcO2
vrmuUz8GkkCqfyP0dbQOWhCw0fJ6YRZJwen/q0VX/eBY7bLZHdCQsyw/Wz8dKiATNe28Ilj1eiHI
RYl8rCCCEM1bR+EwtBDOSc7rInDMWJKA5GthYBjJzwoAp39OQlz39jhJ+VhRDoxA9p6nNjdmADUA
lmu1rG2P0BSdfiyIPaz3NOQkQ73EpA5bTRPM+34l2O2lcAkLeEMSppxUiDzxIUqBWlpGz59HnIB6
VoipTgO9vAM+0Hwm5updusf4K98srqrq/TQmOeCRifaYgxSnLj095ZIEo11rEeSq0nJ2Z1GgWx/A
65IrPahJUtVX69173OfH4MKpQDzViNx4LGNfVcyjqlgoRrpKh74R54bVRCLTeEqnwP6m5xwAbOEY
OLRCzj+Z5d08UdSWwDL27PunB6tC5tKj615yeSm4b7VZUMbRa+/SSX7M9JEeWGO8sYUk/WslcLP8
xSH9AgBWba/NjoLjoRtntFircpYNgVJrcYdOF5tEBYwqslWBJn1cHKgwFq5Q6LAtRnnhVyI4H431
yTuE0Ydqgj1bTCEAcLD5lsjCIsJEMDtsZTqghFWL7CrMZ0qE5R+8OUBqmuaxHULurxgJtjyfdZBx
KgkX5jNiYMG1t5DCt0JQcVjW/LIqnfvfrgE6f1I5flhDfRii+vQEdOMgmgzTpqwzM1fXD2bjkwl9
Twr/ajzbveKI7YIqOgbai9Ag07Mb5+2cuY2XX/ga4iVZeW5SJB2A6nLyb+lnvHD241o+i8VbJZZf
dkRY2zA5HVwqOe2qGMYLRZ+Vv6aC9MB79ck4jwRj1L8L6T9zrotoCQODRm8I/5RnxkBAiFNzhrvx
WXRFHx19/FNw6CtFQTBT3JNMoQ88j1GRb7KcQrtNpsZsszwGIUDI8MBX7jc42j194BkztYY5TxT2
S+oqju9Lv4rI0JCONPWBnSw192ikKwyyWUfJ6H/yhrb3yX3uXyKBkj1EAloBcouZ9vAfdZo4U2Fh
KYHFgdN5gQTTAaUS8DXbFfpYSKfBtMEDa+L88sH49+64LSGQr8uOldsJz2XmX1gQbMdJ9lzN6L+4
1XKp5SIWHgz6MTZEWoxFEEY9lHVfY8pCeYdLXWNiyqSjqrK0miiazsp5DEaHdPrrwJlfcRvSm/jc
VyM7hv0foCVFerNSjXloAll1v7EJeXsM/R8626POa55TaqDJ5CbyvZS+us/xbB63+1nNr8O3l5yT
ldy9ikXwIRRJvCoIX7V+EC5PR/ED3MAYv8h/NYClyijZIRwaWqSkK8djWhlHpGEt1OwP94KnCCKt
GllKFHaTuErBpiVYs114DH+zscDHADA3ZAFoV5qPg1fG5MeKdRHsrUSfnnYlCi+o35V+/S9hf1NB
NPWUlhouc8gMzYPOorc7m3mWxmz9JJMgd4JlkaHVBklHYcAa4rdw1gKQCGZ4j8yLGOndbp5zXJaH
6w75qKPDNN9jHai3C/fPfiTkwy4u9G5NDNklWI8AyhY67makx1tPHoFBss5cejxvYnLjKgRl4B1R
RwQlukH+BqPJQLmCK+RQuErqGOoouh++cPHgwXK1+KP+nKBtj7454rHJBhhC0L80EtsQH6Iq3ja+
8xdKEVUekyeSnIDy5U1PuwCbEmr84ulrg/moc28szzrIKNO/TPuovJbc0dycWHiY8PlmtlUXe8q3
gnx3bfjU2/EiTC9MBgMkIj6dr/gbgGLrnC5tuGQlHbIE31rxy5yh/SonrbJ6Sx5+12zSgPXUp4QC
9GGBc3kqalpooPa8rltEU4+bsCQGR/RFexG8GkqIbbzFWS80gtztq9HdckCUgHPPWvrM2gQNgWkE
H1aisGZbCdXAIm20+H73OXZlOE2as/syHu9VNKu/j2RegtbE37mfOE5fiUqbSiTCaHE9atEi+dJt
r5o5DdTGGV6OPpNtsIO794Bcz8LcJsABWLWezFL065XEzDbqullPx/c0E2tsACLxvBdXyqIMfK5Z
VUaNzx4osPM7rFbbaFoQHmlRhEUpxM58bNZG3H1/h87ueuu26aEUL5yaCEMZE0qBd5g003af5Bcz
Yce4vtKiCTQCzyIKzwCk6nqjcqUnxih2mie2D5Lsui2fSMHlUiu8tRosS0MI2YP/WMe4HKwjLisO
DBLRZxaxOdr1rwFgNlLf2qZ2zOfTYUVEzlfI6laRq3GA2O/N/INwcXnTgxHQD5OPdxe78ejbVxij
EUFoBl3+rSH2eEsDRLfcAJlgcT4Xrz42w7i/BGMqBCqHwP5NkxkPFQCtS4qNJb6qE161ZDMFe46b
RTfM1e168n16N3wtjQAliCnL8le7axcxK04GSgrq4C3FiuC/lasFk+XN7+G/iWVCzoaU/Ra3e9oH
VvDlqSW6OgC37xmZ0gdpV1TU7b/ZEY2lvvAuTtaXKNQEUgT77LG2CqhBuT9vDsYIR8W0X6/2wQKi
KLvPZ9F0lwe0g7XE36WAG1ZOsy0lJ2ujWxBbuGdvhvpb3XAFYB98oD2vfxyBcTw+CFWxzFyn8esB
V2T+onKbI+YI8ElpFe/yjxYw4SyfGarne+gZuDOlPeW2ntnbDi23oJ6i5EuFit1HPEXNgZTTfjou
tcZEKpk1JPA7RXIFWm1CwXpjwODqBCUvZPsBeYb9QyV/hRvilwiV6/5n4g9O35atOnEd2bqjjuhz
qt680qaLfLmT3ZcSN7QXED/MysICI8XZbQJYxhng3ajAklT2TmTMPPto/QCE02F75zUbjMXGtycs
JCi8J3Nu3G9R3SO6QLNrIBrr5bUoYQq2jHU6azZ7OE/suyq6sJqlKvJTpPSTo9BAT4P+mi602dMV
5v+mSw6GDIGci/MwWpgeg/rY8DOyzvvDSX2nCGzbdXB1okRX2+mfQLmGOU8A06LsiuyzsWNzJWe/
b3YfEr3r0iy0OgKfmANIyf/JMUF8djuTAJoG1DM66LYMp+TscmwvgWs2B8FTGJQ0C4MONj7gabJq
UBcUK+xmH8nCH20NgODR42AO7ziZ6g1z7jXU4K7dfcV5ZeZBC1sQlYwE9OpTIz8DRSonvwxj+t9e
GwzJq8VTsp2PbZDr4bwmUQaLNr+GVTfIA5s8MbnnxS9Tn8MTPUqC9Yj3EBbbUbYbF6zTtyJgD5Tr
NXz66gju7jYVWVcMeQOOzQ4q/MO10qLFjAtZV3eeaWEVwELd9GKVM1wN3nR7uhMw/7FWp0v2b50/
/HFm5eMG8r+Mt18D8pDx4jBPrlw2EEmXemN0XsRCcqgZSTE4UZ8SYhRkpyTzXWvamLs/05u4N+R2
Px+Y+rg1JLEkYs2YyYbRMb7QonbCZJ3mJtFloYEshFCadSorBmv8sIXZics6KCujHZ3tv9fnsNMe
0aye+pcSEBf3JSYDSDo9XXJnGE4E2yZjxoqM+j6b0HK2a4OwegFZobyNdhtxA2AGKqsCO25J1jeS
CHqBkT+nVaRSu97aWg+oKTGexPv4KyAMiJnuBbYG/Iy+BQKiRArIoFScF1XO61B55ky2yvPgkgI6
STxhuuE3HuQFUjubrm0zGI/CIn514tRd+WHo5+LcB4EEvFF4zFxwSl4X0In7cBsdmmGzpL1q5luB
mVmENZbDOb7wKEdWXPYz2gwCd8/F9tnrxeL0CIUTGPLlJXMGHvGDhtRIPylCPjd0TEF/sSI5TWl7
kLEo2nvNoygUnxMJIs/MpTtJepbxX076Oq0qqGVjWzMcSUJP92OoxkXzyhT2vf8AZkU5aBVTS/VE
V4ANn0CLJ9JvjlLm8cLgHcxtgys/JqwK603lb5olvwEZADcQU/C/NKEWDv1W2xPudu15Ds4fS8tu
5ayZYAnqs3oI8Lydvihlt71HiAT4SBaGyV3Yay45xlMdi5anxUz8R+nEwCtN2cUCAkjiTiAYfS4V
czm39U6dPVFve+mM231b+ufqpEddRICXG9UtIwYiyh2fPY1UmLNpRpeF4nkzLdy21pPfuQES1JUQ
hOpTU0GV6fP2pM6szxpHmcEvn8a/nsZ0K6B9NCxLemfbFR2NQ6s8+UgNDZ0u5ELzC2FMZl4mqeZj
Cu4x7GQEF0kL1J+ueSBzhrD5X8gd6dUCUyn7Wpu4/ek1o/7FOCHAMg8xR3rxkcay8+KrDRzdHbTi
sLwKJz/KaNIUo0dRceKQ4BKPQTjclyBJqhEqiZluXjHItZua4tbp8zghC6cC/tBWJ7BdJ2+oLrbV
ZAA3Va55iYvcXBfeLbK1mHATWvEaN8Kcw5/oUbXAtrnrMDEf/AaTX+MoAx82zntguX/iyWgFO5S2
bXOp/v/QGIvt1RofVv/9AvLgfAHMXpowwZb0493i0JuRazOnfLrakJn7D0cy3wbulNX/4ieqScbh
fzwYLR9nTVWIwlgLFZ5Qvssrfo+lN4GBTFkUHMdb2E8nZVZnxF/vFG/GuF1jewE492RXyJoD8PI7
KJnbTwXgChbu8uelDqi6kuppe+5vgZcVR2i80VpKfKmKmJh5r2/j8BXxatf+Lm4lTttbmG1QIYbL
PhcbFP8edlAfCXjYnL7VcBGI5Tn2ePfxgL7L6sHS6skOEb75t+Y0SVmV7xwoXelBccEg8mcjxkzN
dw2l/vx/t2IibfreZQJko9JZwlEZNP5wcyfci/xWQWoqvg9/ofKbQovfnYDESn4TOafHnXlZfMz0
Tj970lh0FqPAqixHVAtDqZShXKYzAa7hlm0H7sq0v+QB0gHA4hcWJ8gMCpASqW/3CK0FKrI/vUPG
2abhj+8V1FZX4V8rkQrfreh5d+HdPLaogp6ycQJ+6Oo8TTMNl/CmH+8jc8E42SNOO2pN1/7q4bru
M4AFkOLE8lDhIzh24cMxNrgfimdi+8ltZxO5K7qvsyAKAxrd636v+KP8FcL/A84/r/K6JG84Bm/j
kBR+W2exSpqqxJANdNXsVQ0x2kK8+zNTY0hCLdfvtn/cUgygGVjqa/orVL1V5aBOteeRfUE9aJJ0
AgFU7V9dtnrj+R5gEGByZjhIpLzMNOT1/sqQmsgvEplvOSrVjaGXyIjQpau7WTd4HF3x5fcGwNKJ
CIJZjCj08xwUKrniO0lO6iz48f6v4Y1AEnAsVy9TgFx906Rxiw8lLaClc5MU0cT285hznA92DywO
AlIeOCNblytDP+tWB6FGQ7VmzMQ77XxBGNNREN30VibAjsdm8CJl7g4Z/o5sb19BJSq6FONNpAC+
lVX3H2E+3MS+ixXP5v8ru0kxcsrpA0RHA6fJLKOIIFooQEte4mpjntndy+OFbmj42sJqnxYW5dfe
bKFIzjyq+BUWLwpmXCcgxPBz33G2BtOInzwo4BRsuCdE4e9VFzTQOslez+ZMRfmb/2RHV0aTSWgT
ylhIQu6WkDDf7HsYKIy3XIBCaG9Sj7wOjghSZHF3s201g4WxhgsfA4N5LQM9a/s/v6EQPXIAefmi
CGzBe9jjJe39mueZqN6HQ38IzE10HHm9J5D/BU+n8HJ9iYtK5dHAn6IbwYbWcyS7p1GaD5NSObrq
zq7MTjgdDd/GfL20aRdZeF1TgcPWZwEVzk9ST76MrFDVf115x0PhFtmwSfH6ECproYYqzSilav3Y
Bz8N0+w67vmlg9S+Xkz+7QD61uqYLEIzzVlXunTFs0oqi2C/dJcb0mJ+mfVZjsDvZ6+z72Muwyxo
Qp9oq/Tu3uUxs89JN69LXFML2N1V2LD4o6klFNn7AT3iMTZHnex0IOgXlV+2XFBLn9rsg6Ksgk+C
xTabMMsLGOe1w2VdAcuM6+8pOagcNTdM4+xkI1+y5Ah6yBCWQ36pXepfoZJFLE7XBNRXU2i4PPvJ
kV3qNdiEsyx9pL/WMx4C3m28RYO39T63ACwJHq6jhRua1umcV4DAaXNRaxq11cpJXsfsQkki/MNv
+MxuvgwoSURQLdc2X0ssplmUVFOHfL4xkeaeFHOoQ7wPVJxq+0+Pm4Il/ThbX9dZ4FDvTT5fwNIA
QmhRpjybhtQsZEqc3c1GzyuPgL+eBvIoY8fEWcvPi2pl7ibTEa04qOHzQuIDp1Fsqd8tJkvWQvdi
S+7B6iSm9MtBKjE0toZkwf4sdutf85tCmAbjHJjCx1l7vxbKQj4IizMey9ZeUE91PIdqNY7Jtazt
508J9E64WSJL4FJ6Q/VlN5MOZWrknh79LY5pv7V7kY1/dsOH6hfkhJrjhs+yLmPKRCVxIr2Foilt
GDKDC3Y5xDvs5Hpf6ATqJudqhv0OmueFzS9ARHRjKtliO30WJFhLYMy078FmksbAtrF3SY14401k
iOVBekRAdOTwELlQNbCITGZJQ4JBbgvIfs8UMnECu2+13nIXsx3qmQONz68hjsJS9v29kH7PaCqS
0YOI8Rb4YCyTibslG+/ACzYfZXyQ/NZNLv9r2BTrgFFUK/ge7tuF5ZJiE5+v+LdQo6hVMxBprUdH
cO4JGs3jzdjlPec/8GZD+bvNKCF6/W4CrfaJSdAQ+uvSWCO61uvCqscuPg7zIIXeq1tNz1i2PAQJ
nfJ/nwvdcYzRR3aH3CSzas0h45u8RmbcNFyXx/5+OdwGi477eu8mFOZXmAGBTlxgz36/oumO4Xv1
y0B6s/ykJM0t93umAz6/aBACsVCF+dgI49ozSKoPYDtSMK9CZtwnrpW80rjGpaJeufO795EcV6fr
CEUX1zS4FIgtOy2kbECBjYEOqEeH3KrI8RR6u1r0MxFuiTGov3sOtD0bWGyRLWtC34LrOlzVNwSK
W2AOFqiliylsgvTo0EW/U1z4442SoswZRNDFfA6k3MKWmH08IAuX4ugO3YfqFequiQFF7jncP2Z/
C5RWie4xpjFOGBu/r7qGxdV59CA79AoOGEBX1uQZH8QnFsuzDICNemqJ5p6h1oWadS4gLhou6WJC
GMRW2zmSkt2q93EGc8iBdQx1BgWgMf95c/T+6W5iAQjq5oDPj5z6o6z5GLY5LKeppLOaZwAw6FZ1
2UtbuB2EuV1wfEX+IUh46k5EnskX4kfALkmJUxiXcpzjpnH7iSc23357SsHY2rc57fVeLE/YYoTj
PGXJ1r3hZJtyAqz8b2ELmzZrRhXMNx0CDTzz7s+3u2KAB86jM9oQzI/GdNEg3eoc65KChT5oNV3g
dUfh8WHettxOZ28+pAsi1fCWSIgVT4x2EyM8jbCpL+ZW7MIwqRyhsg8+9JnvTt98dN4vvGhGGJGg
ekNANIXrskoRxOgqfaokfkFFBIKZJWsiCAV61VkjVoxiCSCZzfiSgoqOCIclGvMQmLIf3Iw0pWoq
Veyfpida3sy4/p6yGf+srmU3/6IRqXcYLzxUk3Bb3SPwdSlcYzj+RUL+NaGO1bmWSmJ9ovByaKfb
YNll5pa4YZAN//EKCQdHcMQQj1Yg3FqgF64KQfeTHmGTGsbDvMYGpTVFwj5UKhW1wx109Yrea2uG
Dhr0JG6tgZ51utIJgAN6HwIJoXcogW2i8Ro0AT62rh74kPN6xuFCj9K1Ew2OoEMcEYOQ92Uzxe+Q
LZz+hsGPWmD83qX5v/HG6HwgbiW+9fAwfFFqZcwXPmHgz8Jytu74MmaNkTFSb0sjRgsru+tM59J5
Uodos5s5EgqwDabjHZ1gdvzbj3q6mlSra27MtCDmuUUhTjqlyZp65RmEytPIvTsPt1Wt0zbCr3xz
Tuc/Zq/F5NUHPEG+cHwa+ejLGfDZlPEH8oGoFoyipkcfVFWPN0FTEAI3tLKirnCWbQQYAxiiBpLX
efQi55dWS5IEiuDXzDtIcMCIGnGIIn5SvoxY2gZts5j7SIC1MfHJgz8KuFdVOSO61CYcjYpEd6Ek
HqSuHH6VwiV5mlgiT3/wAyEIzpg7yZsqUWymz4OOXxw1EokCnYFWJLxhWptP0J45pxPC/2X7ImXJ
X/6iLYNrv0jgGM9hfO/mi3/qAXbylA2ZMuqfodDTJysEjejSiBz1ytT0neWkHzvm3e1rEYqeP8la
eq3QXLLbzyw7Y3DHHnx47YJUtM+mid7ZGH/YIvOodBcGekiZIccmJyGEuPlpCGNNwyIW3jC89vUa
Krk18zA7322elPVtOerG25PgCFOnAhNgMQX7fIJXzObB3vXXptCKt2BCOzWkWaddsipD9Co5ZgdV
S56nBVzP9f/zICVHXhn23FhaeoBv3zS+ng0fdkIyV1S+CSfY6UglmHWqctT03m6OJaI6LF0Qz3uh
O/1gti/Sb3wtfTPrgt5vxj3Pv1AyuLdH23Tf7BDOM9h+VI+UHbtTNRbIX9mMFuY807AaIWPG7Z8x
89ZH/sbwRPQAcRD5Jns0o+VG+OzXHVpRAV9a02L4u0x5kywu9KsU8dtqYniCLLW4WYsGGj8kLxCX
+4XUuKPp9EQaPCIfkDyhrRC0qo1eM1FG/8EnaXmuxhA8Xc2xUCtE9pBVeKofvbHDQlngVdDegK3R
OYZpuPyVgdMI1a4UQCJtKz1uvmFqdVQi0lbi8RhRn8x2s7rzGhHG2C94ntrOKJFD3PiCCVCbk8jk
ogrARnvNMW+hXcR+AXi7/CoHUonorLplr1G0CVDLQLCTGz5zOnhfqfydR6KBkjSsqmYbVxtp9HQz
sDh/eBznXcyctPPCbrK8zI1YlWHVtlc/1rBOVwcApf1N2WP2gjDjtkq2Sja5gXngp+TX7qJ0q0bn
gt/Cn9NK1EatvxZew9YMAjH3i39TiptGzinqOmz5pvqqH6rhZxe5DEzgPdqUJFHK8KhR//sXKJ8M
xj7uHmqpXWXRz4TQ3+uyqbrWnaZSrQKHIgd+9FAGT/oaoPzGf0rAFotTW+VfsvmzNOrg/WARd8AN
otAkyngy7AL/6BkYj3JFfry3b97w8UIHE5YdZT1MwYnHyYX1+oTRZpLCdySReVWbpJQsrmOrzhkN
OxUE6NZPOYTwIrRxI5TZ77zFotcqI4h7LWpcYzHbsMDAppYW8V0V1CA18axSIGC+waMHtWXP2tSN
3bhrZRx6f+iOegOdnaHz9ntObrrjc/qavzfYP9dhKyBeXxBu8YjSddt8nKXZNZMikNRFUT89dewu
3VfbkvdpbvyFwmbC4DRyOuupyvO66DCVQuPuKtadwyfNTbs8+X1Kfy6cx8qoyVLN1g6STD/2zph7
3UIN8aKUCXAVK3CA6tVHP/V4vu91+IwBlQqKi5EVdwQoCWQURwZSyf+pFMH00GjYjQI+NGINj/fC
Z1SSjT8zfPm1SIGqZC2YvzZAijLa2RWnosBkFaiTXerN5Xx+WU7TiG0kTbjdqkrdBsGj/IzqCBk8
jvwEW7G1IMtic/6qvPtuB1VaeB4lq+ZDfK0dcOwDbB/bWqZ7rfoas3Vu5LU0mOyDljxmycFMwWEc
6f9ACLagdRfb5UTkll58NjZdaFHxo6MAPuKxUSDFwIpNq/iYg8WH/9+ZtOqtZg/lUDfidl9RBLFq
11E4WwwQ92ifD7MoQ0sfcNNILBYCpQWwVXLNftp04sKG56CDZo6lZVBnlpNSgmMgajEYhOVE3wSH
Wrv3fAuFCFjKVAErnwtNMtBeWmccht7/VFs6llg/8UtQpni8dL0lbMt9ZGZWKXsgV3brZnPKjaWk
cAlGzBwFrgC4PeOwtLYd4oCOuetRtTTTKS3DasMIqIylTZb17E5Srpvnbudiu6EJHwX6Y+DLLXuS
0uSJN2XgzBxfT9jHkBz6g+BFabbfOImGjUHBVdLSSoe/OMCn1cwt2y5o9wfybPnYTqdFgdtiw4Vn
n+Z6R0GJM05mUrmZCqcc5lS3DMr5PitaGybkNpD5RX04YdxoJwHmze6j5M4CxMhCu3szn8KKYjdZ
ELTMaMWJcPcGuG0GYT7ETC4QtOiIiXA+uVVzm7nd7PMYuo+fgC+/GZd1KM7rgNTX6K9cPVlV+JAH
eJqgIOiZOy1ehYaaAFgnDAPL6jXRefSGZCo4UhJZMLZMxocd57yHQeenIje17U7x8tOHg1fuydc5
sUq1gk0m8ta1tz5/TNBC9SxewFSZyHSEkU0AcukZ4aKsdADybl/95nuADUO3kLOm7cx800B1yQt4
cQ2sHDVLCMwazG71TpGhoNUnD/Si6PuqUTOAdI4hh7TesgRI8zld9KTywx3ceLWLDQYew3GQ5ESU
A9+z7pijBNkiovpOGDL+V1VnWzvZ3/5Um8A2Kco9MyqdpIzkI2Ot1IjW/EHFAwW+wQ6b9XHy5fKj
YJyxmyr8w9jCMiW+4nY2Mrh6fOU2baJ8OqNXAB4ZuUGcLOYouW/1MamkGuAWCEqsMqHib5gcanYY
lbL2yCUsRGNms2y/ZeEzjYuSx9If8BLKP08d8U6ye61yzXYEzq0QQnWb21vbkFNT32bgjjf3KWoP
l1EJHpRRPZFFdWT8FYOe7ymULBLe9dgxfWLsUbueMOGlEKvhZo7soOJie+yx8w9OuWxa+TDKKk8V
/xt4FQ/wbQDyjDgQt1j7H9SuOjjlHuj75CGUF9/eW/ye3SOhRkKPH5Lvo/cgVqoNpiTO4NpGTJQM
63AFy/bg3+1PHSPkEoAGkXW2Zc7x6ZdGGUNlUl5JbvQSvv3+0bgO3z2GjuDfYxOTGnzOSMJHb9+3
qIQH4lJ6i4JGDmNewKDT6arHdLT9P6V6njw5NXQFFuMRKPNKI+mI6lk9fLL+KZw1b7BSEYVu/0MN
kHKnJ5KsU1G55ATsHioPovmGJi8ERPm4Q4Lh0kybxLeD0gSl/Om9P6b6dgSg8FKNL49hmevVQgxQ
4Q6hjqJhjBZo6EusDtrq3gYzR7Ec5gbKLSUVlRfib9FL5YI0TKtwAeqPD9AH9WTWE21vuZE8tWX7
LH/Wx8iXRrbIZcMN+h2sjDvjfk7kL2GFTQ26wY5EtwC5G1X8Kftd5Bti6moeSTCMS5iBM+lJNAmY
vNzlapWwXCPDCxe5klJa16vmdadQI0AupxAsQVNI/DZjiQKcQWJuujhBeKbLoZBYLy39WtIS1BH+
WA0zRX1LsXKB0Pmdga8JDA0Ru4X/2kXbtzM5bugURtqedeAU4R3dwZxMqWUenJN2gN7guxsX8s2i
wLrfp5K8nJBU6LS5rQ5Pm1r54JlcLgkVL/o7qj+5srdMzsH0MGjROMFoQLGyGhQzpwXGLnrOEaAt
NwcehpYNexlkqMWjp+Gcbtxw9jDDEm/bMMWW9HVP9ytNrT/ekb109emJ4VYOCXGcPyg2VSdW2QBg
9B7k7cNOULE3nsU23VOP81sHmqMEm84VdDh8cCMNdcGYUszxjsXeZ3HXd4uG7LUtpgfrffMoAxFz
Lootsvw4xpdyghz80+sdR1LuKZUD9We3JQGBu3Eo1gRgEbsNihTPm3Vzv83stjkcvESmQtJYIz1F
XY5h9w9GOdEhsWh1OerokIGtdCausKJUaNYKMe51E2J9kVKRAs+b+k0tsawun2ScnuULbAqUSozu
aRDpHO8gzBD6enGhgquev2r80exjjYDve8mqVJQWA/0FnjoEUoDA/hyBFo9xvkEEkUSO4RZpmzkX
XqNDRaAlYlo8Z64iU7BMZFxz9xhZx62HI0bvEvTl1C+FRZS8Iee8cldjkY9TPqC61A4DK97XO3xl
ZIHdJh9MCof953QLNar/I3jMAehTYS3IiKeOVvIsidYJVxlT7rmiBgmoqz4GhHaO22MeHZiT8Kah
u7Z8lSYHCNLencBnmtFPwlyXegIN2QjKZ/ye05HhYS3Szsx1JlJfh0lAU1siIKhEVOR/qTCqrstH
Mu/woNJnYcwcpcx8MG4B+pmM44e92PBcHX4UoLVfFdqxzlMxcrjmh33XDgSMKBEHy7pKfqv5EW6Y
ucI+oyrQdAIG9fg41RY1WvG4oCT/PPMOJ9S38taLdwHix9xqItyWKn/vUSL2YVrkungS7g257cTA
yYJHa6WTuNyVrHW6Zl1dzb8vA5FKAyoeikkSz9PieLhyU/ihhGGKfrB2FhVXjmR4Ly22JXo7dUII
Ytp4qs6H5SaSMoVJghtQyUC+ztUHE5IeY179rPwVtnWtKYLjzB7sJK2OBI2RJ9DuLKIpHxPHBvTN
e+w4TTvkSdYhAqZqFhV0va9h+ydH19JA8pUnc1HuuIhkYaulz+3d4baFTU2bPs0uH1znsRC8GU8f
3CZhzdNvkPMZKWMWv2fbZlJVnkWMGzne2PGHInZ7YvhRaQjG8T7LCtVWNYmTjkLJkUxYeVSUgIl7
jmZOm+0a8VYSifhWYV+YsgXUt9qbxiiX7SdzhtXh0gOXBdvlqK/MTrVhQ7M70cNY+NeN0rOX2IJf
ZhgCEvcwQUUZmnOX1DZkiHwU57PjMT9YZJkVKA+eruiVzj/CqQazYuNV2M8VKP4134exo+hQ5FVw
vIiooWvlcaY8vZdgWHUcO8xD2n4Fl/VK1tTLUZDrNtfjib0RfYq0feRmoN/xkrZLK0fchgEHMvwi
UICGNDGcp72iQRgg8x6oLyvjZa+EOwr1RComzoQt1JltA1vF7eZDoOK9j1YaSwhslbIeHUj9FNWS
BEjALjhZp+us9qzhYf+VOixDuTusFJM5vk8PIfXQxBpga6uFS+iEh/TV9PbXJxprz4JbJLO8Xgwk
oJXXsVEDyNUQqRZ5SY4ZSuufR//mMp1iZDIApgESa/bG6+DNgQlttvKieK8vTdX3YIjPEtgZgFmV
M1UK/HcpoftdLdSnZ2gpF7m2VzSyUfcNHMaPG/H7rzCC04WGiF7oFnbI5DPGdnC/gRkSpJ3vmUFE
WYp4yWOl+zwGPR0v8XMOo3CoY6zDBxcfocXVMAZzEleBfWZzvjhCDVD0pBWZEXaRqhXN3kDSGJEs
k4a8AFv1/lnWBtOudSXN4IH60Za9Yumvac7P3pch4v/DTf+thxZ3jcuG/LXGiqBu/0l5qUinIKGu
dVDsKjVzJaG++Odpt5e9fi9y0u29NlvzDU+iPuGhcH4TnazT7UiPLQTHV9EWfx+6paNDkKhoaLgw
PJHX79iIxkYlIDdvALBU7Zlsmyy++5TSU6Fbaic0JD2Mv7lxFUA0Y0dIrVd7wG0Mk1KKerhrhokj
b1vGvNdWN6lF81YkRTQR/gZub5hHApgBPDIUnUYM30ZCwc6muWp0ZsHLj0v/umNvD2zjHgI22J0U
QlQNG/lRBl+SjBXZ/jDnx40Cgz6O+2bzmqWbOOb6ZweCx52j3CI2+QD2LhrWWfR2XmoQoB82xyeJ
uJu6x2KyxKNyl4tN4Q2FfNAV7ScsqkgHhhf8VSxql4RoObnbdkFb3LuJOSQXqVzkKNnTagZrhvN7
oiDi2PtaeR7HtgaUC8iOzrm1GpatgtMTOubi4O8foty8M7AMoZ1QfiYqe7Ej9bopLG8rVLidJH/f
cdHxp60ER25dB/UqCWCYjYANYMYemkTRrE5Jqv5lFRMKc7RQgf9vEO+a3nXfXp6nP1IdFAGDoluB
8bjSRtjTb/s7imPEFNEifrkZN1q+PZPXopI7aE75ElftljHyn+/ywE9npMRx3sh/SRxTIU2OAogT
8p27hDNsCb+wWyJCSpAo64eog1+wzQqpSW0R6Kmn5vYtSyUccHEl0NgYK+2Ee1WZC1ay4okCjdJx
p8rj+lNq7nuBrPAKejCKOibe1ZtZluPpyy8rdxAe33NewOGKRkZuDWTL34jcXp9h08yiKKp25ZXa
1JFa422fDcfQiAvdavzjqvrCL7K5AtFVdabaTYa5aT01TnkHUFlg5edBjwXdwoIFOLmneN8BqwDz
3dcxH3T5zdWPIDed6hU+y6QsjKFcZ1ALZMGHbec4B3/eKPfa9FY+4UgCcigL+Zb/hm9RVIDaI9t8
2x3E+e+Cf0eGNFMJxV4EWGTrEmvHjhk8wBblbW3mC7Q86aFpIBbhMP927vnwQSZrkN15FpBYAE6Q
Uvh/iswn8jSmyNFG9u8UnDZXm2WGyW1cuDiUoo2iOsRcyR3x+/ET7u8rWZe4wzyA/yr1sHT/I5Pv
ExfPJN6HT8Pp+YtMeALL8Qrqji7wRlHEc+hzamNQj6lzSNvXkPkfCPvq3oQwIWg1oTN5PttjNarq
Lw3Q6CUjK54YvxhC6j5LJVaXm7TD6FGX4s+umbvKAcmV6YuuHPw5vZEAwE1uZbBNRhWRb9Cuv2eP
NTDRvoaTkojBhz48fcboEAjwZ01h9LTbDU9lp8F30yabo+mYg38VVHK90gq0sD3h1scg7iAKH3wD
Qf4VIOCWB6wquaZbsXOTzxch0WqNiaisWXkVejwaMp06dpsE2AiNxHCU75GhHByjzd46TQZy7+zK
rN3peLUrh+kPprDlXek9MH/CW5HKSjjcEyki31vUPKotr5XE2rlSp76EtoG6kdMcjyMa7zlwuR+3
Mry9ROPUmpxdaAUkG6LysTsgL75IxLVd4qIGGHYlXJ/jx5Y6GelfwDsoNBjd4dCn+d0lKVZ/L6Oe
id39DCnufvqkYun3JoZbXUpoCgGPM2itWsWKIsNIJY6YAfBgssCmQ7/hB54NlayNEbeHlB4xGZqM
pibqLFQe3jbOjwayZwCmhsYO2He9Vwm+G0JV3Km6N9oq3q3iqBxO97fC6oFAbt+qfjDFei5XrQMR
lvpTCju/YMkg7MXOeOHgEKVTAzQ0GL4eObntevklVRMX5zFhg3te2Um3DN4s6i7weDk6PH9iptyB
LBqfFd8lmmR2hdAP4kwIx2Fp8oYA6oHpz0eVOId4xmAWuBn6a9NCrVzT+qnImxJiJoeWqcp8R7Jo
UMozF6H8C/2mrS4lTmZ5qvRKU7oJzgj2APD+CDaNynQ/pge1JuGPn7eNJUIZpj2FhOK+tt6jtVe7
hR73RqLr4N1sOY6v3FnFyD6pdjulXd5znO6Gb6C7pWKiaACq9F/xcHClJTPGHl693f/EtcEfrLTh
90tPMVC9cWGYTTxqgtxuCC3/NDywOM9Aepnsol6Jv8itP8U6kv6I0u3t1AOXgF4lkRsIL0szG6fQ
uJbMU+cmENUCyRjAo7YywhWLzK5rF1PFC9ridA2yMwbDwDKTbTFYG+QP89ZCldxumGe0udM/KObY
xW4VRSTXpa6FZ0KvR6Y79Osi1BxLPfS6MNUiayiHXhLtmhgIRpnwVDMr1jgAPQqM8XGO9jnew5et
S1UvwCILS4Q9vXGbQAIH5yi+TMfEzRzgmyp+AWa7fkv29XpDUQTE1Xr1z7LS8H9bqmGbHXQiYmaP
aUqn4BuQPwGH/JtcISNfqP7kgXjnweZI4KrSoDJE8UYAboGLPzrE3pRACnC6LSgUu37gxYhxLtvl
OqbrHzDJDNi/j+gi/Lx7kj8A3g0eJzmEswQ9Ygr/zs2IXx/eANW2qkWFssjj9rRC3D62Gwvh475O
JVgCGdBbtXbCnzhmbuu6LXaCPgR+dkyBfed81w8j5JzDvGEPN0tbDYY7P8d/DN4PPVrtKLn/uTUm
vPbwc8dOFtIBAfetPNMrygex/WSFKxic3XgmMgPSsIU4j/On19kG0XrKVy0ur52IES9BnrDLtlNQ
xrSzhfetXoV6lOn0nwRUxUnBAQjoV5qpJ8E9eEVbGUqpeJSyUgkKXwrwvhyRZ2x4T7ApimMTfRlr
BE7omTm7DJHDthOq7OIIg8cGOK/jEM35l5Nc1+isMM7DaaGYxJJ1d83ZDnw8Yfbm74uM9qVEHG3W
sKY96t41EyuVNcb5Pb3cHxDrNRXeMn86o8DZCiaKa6CC7Nk+JaiQPF0Fyl/vFd8s6WruUo9CvFOx
zTBnqKc2+DaT/32a8ydTz+NafePD9lkStAzW+sFYeM2BaFX0gj1OBYwLJG1OayFHeDJBxHJpkxLc
r+Wvx/wOkrTBtotCj1OLH2DTsVN4uCcMnq+5qPsqkwQpR7798sDY/DmuhWDZUzJbPKXy6jIOCcjs
Y6WSwdWbPbBL/hyE16kGHd89x55Z1mH9642HcAV3FuiOqV+TELMXblWwMBEUqu3QCTsszrfgqtbo
AtPRJwAUoBuVLVrkAfvEsP7WMoGbDEV9RlaRDABo29AbtiCeH1ZleVl7MPFuF2RVYKF0kIcSu2IO
3fGQv908CtSSnLMV3hVumE7Bm6Iu9ExHtLnIucxSYUSxSjyLilHh6VwrtQEx0fz1bH+zIPZS9vA/
TLV4sZsb+BMGOCHr0T2bgXH6cKxldOGrjy1sWTOHrhFcvQAz+jQSDtcWR1QSnpJrVjJYMmk6qL9b
YlNEIP/eCB2xGq3jwUGlSOAM3kI1oQPyPhHZHruUbd9IWA43MUbGNhNSD9XP6JQU9D1GGAdptevL
ImPaanVrl1av6x3GYbUC42KIy8ND174E860ppXavJV7O+r91zp9aEQ2tJ3Fy+Wb7t/fkequfshH8
AlVLtX1KnjkclIiD2K0SDRON5SAEACa6sgH/rMhscJ9M/H/wtDzdbG8SEfAZG0oks3n21+AlcAn9
tSYdzM9XU1ncjGCqZ0+o27N9EHpgZ91GtEeNEvNR6Qz1cUWHY5Pc/cnyppsY/0znUNGBHDO2tgM1
TQnXqcX9UZ/mRZsD8H0B1D2ul0rxtIFeRBPclv1tEyrWWbNa8lYGKRiDR9Axr/j8EVIW9CVJD8Vo
bhJ5YRQ/utnOTRnqX/0HQgxoCa5ChDNo6zJxZQuVJoBmPEl4l8TdFfa35ytiI4Ld8x2+5q985CUU
eG85I7IeQm8nMEkq3HLMwE+UrG/hbBVUVQv20YlpPgqY0Om9n/9HIV65CAdIzeIjk0AhW9ZlGR5b
2pEQOXV+yNz3+3W8ZtubfqfQTnpKQk0ceCJ7SbQOOAxk4mfTElPn92iLiQARuYkqF8c8W7gE2KsH
GLpnzSQ0guqMv2YEujkObcHS57YRzg8XhuBegAbuUIVMc6KA7XkOaiEMizOxal+cZDwhCxbfdRQD
M9kyYyjUuy2jID74KKjQ/6/ocjN0vwL4sTdVQdjzkFFS5jpU2GuvfhJgH+Oi/StrVpwzQdLWQcBj
gRR0+fwA9LGkaG4dAZGKmePGOUs4bLfSlcQRV431Li2fRSKHT5F1oCDHtjO+y8/StwsZoRrcLqi1
Zt3kiMxudtLHO8Kz/iW38tjgj3gp7UrDoO6c8zlZJFWUxg87KqTAoSxTL3y5JDlyOMFcaNknzHQw
sUIkS1D/S8rv5x30m3KvjbkWG6W3xBYm5srNtQOAhjAM6h3JKIG7t9i93MS27qSYvABWnkHpJtaw
t5/o6XrJkGKT6P+hwIYvP9BO2+NENzUIgOtaZfRKPESF4U0C3ndlBIFSpJpZsuNMYB3CL+0xHY5I
b+TfoYy1TLDDj0P8/JKgRHaDkRocdbtaJbDirZCPS0SHvRP6Dosck2Q0m7n+tQtKcwJ9CJeUOcNJ
dJ8clxwu5LToM3d2LAM+8NytuamrRPsVHV+NAxOOeV9LpVrODwcbdGoPXzRCoa8bvwFViVwSPu5b
ZcLgarvPpTSMnStfrR/FkXQ/MWv0TzgEfxMv+delpaj+Uu+TxLorkisYoVsw234v9VmYRiL9hO9B
utYBV0L85BL0m+BTLCcXVZFkehk3+ZK7nPf4/K8/GGx79Klz3Wnptr6CJIZe6rFsxcd72VzUcF07
YRmgLbtDHVs25wSrjIZ+XuJpMixbz/NrR5jP4b5KnVv8aQXq1BxDrTe2VIus8URidCMhkEEzOp9m
q1uHi0aPsvdJMvC+vez13rwnkJJ5IZKS90DAEvGO7klDMNIQjufIabd55eEVtZMdiA4GnyvLc/lH
dR73U6smqzp4YbWAdlcMvb1DUNWoTJiGnAiCYfvGWbq8BEbiUKjjyFPWJscI0CPv+t8BzB/bZeAB
IvPwHOV12fdUa8STY+nG5SWCTaQ5pC68aulTCGdml/PLEUbEcuZeR4Yy4POdoOXNMQuhPcOdN2TD
4CyZI24kmG4YBV12V9ZpSQ+HZqMQMZvM9Yo3IozpTPz4txJH+m+2EVrJYj/RqzE1PuqogHm7wPNK
5+UfxmlnnUwgKe/Tn/LftdFKyXYxlwbF9+OL1mHeJNm6HsrofrVYbzmG7/0OL0LJFCI88SPByO41
+duj2NZP5Dp/6+j65AdEdiqFOHCQosvjeKFrKUEjGaXuL4X2RfAdq8ro11yEjMPeIrZMhMWlhwd/
AZ1Gc0w60YIOCLRdLUnaXJbdHWZvfmn1cDzb+tBaT1vnPteJqF9PFDQ7fDmojouAz/E3EBEF8DaN
ey+9+P3BGGsjfJX7RimX+mNTJEJ/aqNpUXYc1lxW6LccX+pfvk8aBa9tLW2UOEGaAEvJ19Jy2kWZ
Bp56XCV97psmZjc1uHI0tyKbBUQ6vvrsb1ke5DHZ3XE1CljLy2N82Nqx/vdYCv5RYiIJETIIlNBA
WtLADAAg/wU6XabjGW4byCWSFC+QAlVyNjL2V0P1fEF07ZOdN/0+y1ntDuCz2nRfnKCnvy8I7DQS
Vha8AIG+4K3NuQhE2Vp8MOE9QA+vMAUQ+j8WVwVre2jMe0xF2NgIT58kv/9OTHicAWGCqhidJJXI
Jy7SB1WXQS/+Wysk0dB1Gz1j0naX7Zm2Zou5rYVxbSLtvM75yNXmGMI0cQtsWskb/fjt8poflO7l
02agw5QvFna9TcCRFDVqzPAbxSML3gJPQBy8/12QyjVOK+SskajhE1K2hSbvinTOLnRA57TJZYYJ
sDKj92JTxsHSnTeqQJA5Ao3GMwrYARxFzkGmp0vL7Z/xxdJA8j6uM1U66IXVew3ZapOR6qyp3gBw
G4C5iLcSHUrTfqrPag+88MZcfO7r9J3NBwM19hhi9qQtK013rAhCUuf6sBAZg+d6VdstibU6zD24
MWwDrXd9IJoAnuzFnJ2OcWlFQc4R3yGbGoL2Vrk3xJqB3C6tqv2dbXIqjsJdYXe0SW3Ks1knyP7H
9Q+zzEs6NwA4LO4s5WIfEmYgGjv9qeBELj3s4UczF3U9Dan74hLF+J5UXQKLF2G04slCsU4sZSv5
viydJ3GhbtPzVJaNZAT7Q10vfWHkAR/L07LLBgTWJdiEu9LF765P5d3HSq7Y0mk+Ymheyz12+MDW
56Txq0eZ4/DzPZK2XMASweiKZQVQ4DmhJVtkirI4rp4VeVHc3noU6+w1qMJnlU56Cpha19nxt03Q
wsB6d91/DcJG7hmwo7VUixKm/gWJ2izMBUadoizOATuwSwb3zjgUWWZ9Aa0FBU806qXZEC4uLMX4
AMpsP8KDCC1106obt3R+2mZx5IW/vExvmSOvRSeAwVFtyQtKJKRTxCX6IFLpvdEfrQJhHv0jdsD0
GsqwL23J7hzwPr4CCBLPj+uvjElBlzIA6eAqM+8uBjoaAthIXw40MZgW+asbyQBEAIPswIJcXDYN
Rqz+NOLeuafqWlzre6KSsICLoSSSDwHPuz8NLnr6Upe0sYHh0TMGS8joycNCLIbS8q3R+vyCOmwQ
8VZRkoTxJ7oNd7ddfaD/k12GAKH+fG3JMpgwYGEtrKN3o1vxoU7VD9HaoZCaeblBZfaN2h4keZ2L
7L3m6XtqQ0igosdZ5xzxI6q+P4F9kAol21w9Eyre5Oyyxb/XfCFWzmpuUdWxbhVa5BT+FRzZQm7H
PyOlKISrTTWmJ9l7d6lBqkygUQoB9xPz39/hebiH7ZYdH4etCGUeMLRvAG+W19gq3Vv7CJuogWvv
9DRjytWmS8YmGlH05cT2np26i/TIDMIf2ouuKL483mbHaW4NLsnHcv60FCNg8tBdzlj5CbGUH8gp
ha6YWDlpgiczFwVT8RLgxDRw5OJlhVMn/ArIk2xmDcvotb3RuV8iGlBxPqzcWmT+JM1vO4xKB+D5
RCJzcV/OQ2ahmNHvJfa7YyDT9IQUmMsE6NCdFrpaiI1e42wjcvhLlRCqNkjRojnxXprtZG4c5KPo
BtNCOwYV+1EfREDQ+/X4Hlcmg/zlmhVr9H3mC3VLjhbYM0bzp0SG1F7VXcbWGFrVhDkWfA82O+ds
/pKRcp4VhNbWgzM6kzHCcdB1LM/wcoRt0UTnc7St0DMErzRCX177ne0Ug1Mcd/CwgpFKwK/OmB02
RpueVvsBnZEq3dFOU18fJ2XZI3WDkL/crPqc6/cLrQtfeBQ+x4PZQy4NqcpIk5H6oKvoUAzIoCKH
CWwdp+/JLeCchzQ6DYvsqoS3bVzididrbcwHOCfUIzdgeHdgXOYbtavo52nLwSN2cvV2/U5XxRIl
8eMTTQGn5P0pEPa5prd+vaVJ+W4VBhV8vcOAmRwTVII8a9g31CM/N5qOHgPvPs6NuyqOgMNLk3Xp
Pm5TbBVPckrWUTFH+eOGKE7RI7ZQ8wVqUGobSdi18d/4dKcQk9hxgcS23eVDdsQnFR3UyX0uEvnk
gVfT6VKMeeC7aCF7XZnngbFGc60D5MyzPKgKKwK8YPniq77+6hAcl0wrweKfWjQyyJ2TyEoir6wC
+lWxM2JF3rvXN4Six4ZnDv1PJsDv4mBtkuSriwkpCTugxwecGGZP6qirGtyC7FisleIs5cX7fKlW
op0BD8z/D9OtZauv9qC6YRwP29jfcTwhHmPokcw0+I6QVVA8s4tNnJ7M7Tv19M6rp+l7iNAhUckR
kfApXyIGI9NNCQg/j69buuJnj/D1N2kdQ3iabrOaX1oR7VzyL8l/Ho4Z+yKG2XjRMVaSV7KCvLjK
u0dFxTR0TsphG4pE+/9x/8dEp/q+poU4ZtZVz6ldHQTd7j4n1bvgTGH7wGoB4dIvqykC1yIZp9Tp
sX37UcIHd941utBZ+Lzwb+NC8otkPmXWZZI6hMl0Ts54iG3mMDVRJmVHcD/NuRiwALcQQC2UvDZg
iwzrK6Dxc29EwMUHQWVNp1I3FZq6mNE7z+g+CWKymwGDj8ujLqVLyOdA7XzDWfgo13bKCD1R0XKp
+JkXlG1qctntKy9AHlhbMnUpxhhL2khk1vmeRINGV1GuCMFo/HRyKPV/pWqO9iOAWYGPFTqSBbwY
9g4navKaoisY7Q89lbfkKfMPljczdzXNvsWgI5Naw4c+2vsaf9fdEzBYeImy1Wr+LSOnAHnyJeVi
JXj1ZjFhLZ8URMHRKmq2z7DqNYEzIi+fx9yF2pF8kbBgYguddp1hqKQ4kJ28z0HpziEl7VnFNaPO
mRkcXCab5kwknRn9GwTaxTkX+JTEpXd2gddWLxRs7oGGgB3klVVbTbX/CWUviliR9gwpDUDE5X44
GK2tAUnjK7sFNy6zyIXFguC1J21yWi8cQ8MvHyeqgygEpynG2caAshc3A/VjbB8W5hNqxrnOtReZ
zgbAi9/ELMHn4W2EEVDxapncWdsGXKFRyGukp8sWqzSKroBqzgQ/ZZUbiTJaYAud7CfLoGaaA38K
pNMsWjnGfeMTtSTowG4ZfY3jP1IEQQzSHpIShhWZHM8sC5IYgplfSjA+V7LzXJ84AYRujIeDSoft
UMWVMDsljaPEKS85GdIvUryoYBHFcn1WufCzv/+9C1RtRdiGErrE0Im3dIbpBZ/eCYGAYovov+wM
Bs04WPS63FOAyxZJFTfWDpG0hUlAII3jzWuOg/A6gMymkAycOGg+hvczJuk91kTPPtM0NXBYa3cq
tse/8OC/K0vZI4CtwhhGEicippWrFjJf3ho0NfzjdZo8MgsE7ng8NZy8y363vfJMDr6+Tb8RZU0g
j8pnDGdM2hYkOffl9csvK/QCiSxV88DOjRwHziY+qouLoJla/H1nKNWORZAiQUeb0krTdoJCX3SB
mHl51w5/gdn5rBjfLIzJeBStZ2vmYjInwjEP8V2+eP+RPDXZPGKLLVRK2PBrKDHolq0rhaPJyeEj
1TK+YhQgMq4eONiAK4YlO01rmngmYgfIaKc1a43ZTyMtROoGAfWlpmC82Jnw/XllIBVbyV9UNzyI
eALU88pR7vKSjO0Jpp2EqCjExCMkfzO95GmPbSPwT5Ib4Gr6LdZiAHo+412Ku/J+9oIONRhieEaF
5D7Cz6eWHVQHUPUT+YocJZM3ztESa9JQHEadPDrjqq83Hy6+mowtGJXO0zbbna/qvYkttyn7XTpY
bxePOCAGnayT7VQl45BBQF5x88k6cJtcVPHctuaowewxekS3JqZBBNzM3wTAEVptIdyAC8GoKAV5
lmnqu5sN/e//sYJ2cCw5lX4W/f1m4gBu1q+VDoK3hNFIcxuVKpT++Ok/03CGUck0CCItRxUyvmFX
+06DXa1ohoH2bpX0ijmlQbOq7Xm4vM5L22vDydp03zqWJsRyENqCBRZfAZI4mkEi3L8wdQUq3U9H
/5+zcgh4ZQ9jtH2WYqZIGwDvLVE2i1GpjS++PvtQkc56/dvuWKOwtXX7cSF4y3M2s26M1enpMuSZ
dWAGDm9OuDR6t3DzFI+iOTbMWZxavN1dayaccwGABt87UI6RHvnq7776wstqpfML6YtuKMhemuWh
b2Mo8Ms1xXcywckOUhL9hYxg+MxFlJcKUVUanX/2qDT61nkI+Tc8HTO4yCCqjHnyhYE2FX887YVQ
zpm49G3cHMKLUdXjQmCW5gYe4AF84C8xcXKnHIzZBqtlqux7yapBTcwXyqyFPvz0wMo9QeyPsUw8
r5tmhqXfcucg6/6lB6eO3yuAgqsR1iA7FIdAS1xLVjDTgb4tZCGN3KRiqX3KJ4bk7amwwm3yE0aI
l593DsuPiSa3P9rbV7loHvwwScjBZ/+iImUUXgsIfbvkNRiNhtDX34HZCvTKeh34UpPq0QclIGYs
qC7r9br1XponefN4XwJUJN+gIfjl8zU8g/9d5RiiclnueTHnv+OuO4yMBwuCLEN1Mb18qo1wswFL
pz4QRwjZQh6gHDmsWDUY5FFZulrk0xzzJLmd9VjAJ4TCmqveeS6vpmg31LvQyGK+onYQd3wS6zxu
3+fhjPXys2AP6Psczkw8YM2X1+6s+6OVMzeG/fZLI42mxHIXKpkmhtrI5tG8chVgBzo8H+V9ETwi
vZSoLfM7VZq4d8cS3GeAoXmvTbhS7VaUHW/xt7iTSrxVUI3QZpEp3XUm0TZLv4bXVxfSe5hYlxHG
EKPSNyG2rPSRsyqVWKNBLqpL26zQIvpZO1E1b50UZ+SdyfXNUnu23gBZkT+QZPcIBYha4/ZVK6VX
f7RACkjCHULhphX4kPkqJqTasyopdyDppc/Xe0dbAc8lHc4BNErV7RXsRrcN9sdnXUXUONxOuGy+
p3Fjk3zSOay40DheJ957BM5fCwKEh4pd/uD6QQIVCmnCR8gNuKbReL/IlnLnZfuU8uaFiVgrdtPq
taBeK/ljqY63jf2GA/k+EaBhxojoxm4jt5Lf3fv4vjkEX2VmW3yNrltG9qY27GkOiD0CQoYHG1JV
SeN1JVGhjwrMmRHtxDiuR3uuOYG57mSrBirkZ7eUVqBgK6sWxp84AG/stKd9kg9Gc+DF4Xo00p5e
xKWncE4Z+Vjfsh60p1NONCsS1OMy9N6fKNkjl+C+a3ksfxJi18NDMAmEuOEgC9Sooev1HkqrmZUD
kPZy+MsoPBEuO8k1V6G5XqQCvddOcxQiHi7TL7bzMgZGaw7/OKGBo0uPJtbsgefAwkXC10Rahl2l
6Pw4TdE+xVTz7Cg59gOvFp6esW8z9Ci5+gvKxbhhqi6PWDqsjzNSaUpqJg2Yur/nyC9TTG9Jr0Ex
M2zS2BeZ/Nm3dS50IRYSIZXFoC3vPsRGG/H5HPkdDaZnnLtUDqa1WuItI0+qWO3W9AqNHwCT1XOA
ufTNBmhErEzo5RDN91lO2ucLZmeF8orIJqcw59Cm0tOHhbZZ8j3fU3efUO8Th6geVKwyUyV4UTy/
OWjVlrnxHplomDGhyZJL/CJ4M473AZWGyzPnjvsptAj9oD8Ke8a7vvf8pbJBAVsaOaV5iBjLpHWD
GbO58mPM+sVk821DuEM+ybeofnP63TwKah8JkBzLWgXkrk0+8S3w2/GjRPABQZ25yIxAhtpPaU0e
oD31ftSAdLf5GN2mPbBoXZ1xfGBMXmCIVsWXMPmvmocpES7h9IpkHrj53QSiYXBdUT5COKE7tpAf
+hksiMfQp26vk9mgpR0ZqKq+DH+/jKfLHhSWcU/K3zvSuLZKE867ekBsiYthPvFHlhdkSOv0YXGQ
WgVqikqBT0lZPlnxE764/GQICSIh8r9VDOLObX1qkM7mefEhT0ioPn0DginL0cjvaYa7325L3lxt
861rdJtt9na/N9Z6Qn7hYll/y0un+MC5S4tMoeCtNkrhI7GFSvq0czPNB63pmE+anMvQlsdUA54u
dh7wthGHTDyw0uhmVyWh8JsVeMbira+hDGpJBa63q+NA9G/RRP5oLlHduJLTox5/ewJVt6fRj1RR
ZY0/EAWtTF2bDX6j1aLPDVFuqsaO49vvL0OAIngc0dJ1/hRLRo2ZHrwws5oxXK0T8zpl8TyuEzad
a4UxqEIbPw9YVysf63czd7YYv9ECmQn9uT6C6e50iXnu8EeLCm8OHc/0YMgY4lk0OXgR2+pbRAuw
aTkd2ncBaQqmPZC4lh/44h32omyCHtWgb4BUrI4dI1MDXKrzljqQOe5igSN35GzArxWwTgWrJekY
zgR/cclb2Vh2jlln3bVE8WnKI5MbSdDAOiZRf7fAQoZ/eb9cDtc08lmvPWBCQTsl95E/veSrpxIM
9XsQzi0JUqc+VOMJ1NsTBQrvk5n2GQ2gTt9YYFPdY2PMnCUEYj1mHRC2++b9OS0k8s6mYnM92yeb
dtXQ1biq/xgU3JKQufSjnnLfCMhyiQgR6Iic+Apy/RJbFcYb/7r/o+ONyWttHLsB/nT76XlL7oIq
u7g0lru8csMGD8zJJUl4vIV9Z4WW+vJjkY1tzvsLuP7j2nqbTb4bSR3jwvH9bqn9hBAlMPh3bXfG
JN3W/AXApMjUwKHyXkrW30sww1zH3kJp5NfB29kbHvy7ld0I8j7aNfk/4UYZLM3MagjcOwniqMps
Pr4flEzLtO7rPQH4iHCDuH59t22o1p+vUqNfOPFbi4kfhvqQX4JCP3UkT6Ib6H9YypW3LGLewyrX
TrKSl1XVZNzROILiQwhJKIvpfChFIGf7DiZQPdu37lC7eRoPNNwIQRHy9FcwPF+haf0hO5fM3Bfw
3HYcRuqVT65Qc8HYWCrekOz/MVCjzWJvmf5kpjY3tc3SxOWg0Qr2Of+aS4ubc4jtEiXMImNe783l
LqnDk5+6r15c//QHOyDfvL33QIzoe4UJWLPcu5xPfnkVTWWD3sWaMZM549K3hAHG/mSu2attqIcP
CTwl7m9ZWZmEjwScdhTYvja75rBK0fi7bDRW3IWTy0EjyGj5P8ak6d2tvmQox8EGyrnoNNY2l7RK
owO9pIvSSf9gye4V7G1HraNs6y11xNcu5+o1kLdFdf12Mqjn8+jFQkN9sYulOcQ/j8f4OGCuKDE4
XHe32COBG07tdC7SG03Sy6ILB8m1k+KlGlZMO0KTxSraVhlBIBF8WWjvcy1gWXvihyiMMxKTRVqT
Vtt1dSUgaGHnH+cgElLYmwBRDPLfXqTRYKUhxNbDxd6lyNPu+u546hVAwTrj/Ni95yuLGKwnknFd
qg0tQ7guzqkyenxbPWGm3OHcswqXSpPmf85uavMGIAcqyEtXTj0AG61x/Of4V7/RZx0ZqzftJpcI
NYBFhIJirYK95MnSJqjgZ1AAgD7x9O6CoOiyo/vRYyet1uOfx5bae7KNVVezNAw5bxIC0bZhX7H1
47/lsJOe1xycU+jcRVww3McfcnFYFxfRtDwNdnDNol14kLvFIG3l9g72DBXzbfUK4rFO7h65XfcS
n/uMQAWajIR/4JHrXJ9S3C8DcFfUS8tbup6JBpWFOSV5TJxz/9PLFMOLnKsQzDHbxDFv8rYZy3UT
rYvcXkXkGfO6eqP/DXgAEl/Q+E5yhQMq09Ph6fOjK8oyJJU8nM0M6CftoOoffFgwchCXpXlzACzB
hU7dl1XVEYle6cthXvdaRjlTkYmfPmnKxk49b2KOM8/Hd4DbkaGVnaZ54K0T0NR//gJRYiOO3mSL
q3jOSh2+x1fZ8jzyuIpkF/Q1yv/i03iUHr84rZ68TnEkiPKlFM1JLEGBZQ2jrRWY3xqY6y4hQeWj
WOnOrq70U5nVHUr/g8CO7BEhtCASFShqfRdBN1PpIaxfekceE5GbHhz481y+UpzMSQpZmJbcIVTf
AO7bYhiPBbHr7xLq5W2PigYiUBXM0incOh0tV+OviAne76GVGYvKaNLO7xdU4MVUCDJHNCOyWdD3
P1VwpiHo0o+6X/zvOEw44MuMlUdCt6vNpPH00bsfc9xqFTX04V3d8i6a24c6ZyKmft9FUkPoIKtr
Kb0my+jONMDX+7szKo8HZPA9p1144p4PW/dw1hPOv1anyz5Qr0QsazB0KI6PNznBPBdFldK/9gJM
vq4dZTmnmNUklxiEapNORYJhzHyy9EZp5S98oDpgtImnOHgdchzWqat5VU09cjFZD9R5Lyg5rwmN
XPqmcovsQsXvtz9CQGEREWGY8ExchHAJlj2Ud4esZwezhVLWS/GOoS451YA3m+93ujw6EBk3W+kL
Zg+Gu8jQmLpSR3KnHe7WudRyBDX88aq406eE3LB4DcNxFulxkhxi+NjkX+7h+v7pmjh7d2rTZRdC
YxZceQmfCck4kSIbyFj+qzFDxTO3mYwhMo+Lo5ily+0QDTTiNkZnLHPsqRGq28SeHg/ZoopaPHdN
oZ67KY3rDJJcJymAiTI0pTRBpshAaqAPBrjzRHPwA3WPB+3go/WMmO7LBGqiHx0eERyQns/dfbWT
cN6ZMFHDG+x4ZCQM+gbJzc+OuW3jWTIXCRuXBn12rJizPlnbPpnNlCRBlQ65UIBUQju/ul6YjAmt
60pHlaCim6K/6CsjSRYmaIJU4Fm6+ybVUaJwFpKoDdSWYoicUSoHkZDokHSjMs0ubqEc/11IIWAN
LRjpiPT3RUA1Vd5e7+TpVUO4kpmBB+CMR2ShOkUa8Um1Nqupq7sTPBcMgX5oBOpzRG2dDOXlQ+7i
mNWeyLO7Wo5nnGOeFktwoq5VTqLcNvRMchFafGTq9S2Wws5XNb+3E32HtaWkZS7u+/hSmsYWnBv3
bV7eQSR6RMbFvYqtlrBhntFkRnY9r+dOdWdmNZSPbcGREDSbVNclp/2l3f573ILChm+uFgQ4XG3k
sF1VRhr/4sgz2JI7MFkdyVc99uvXJ6hac2k3MFcgY6m4ceLI/hB4e1YH02JrWFGCAIA9empCP0bP
tQNtdlODh5CghtL4XvW+1UZE6457zl/3+GRNxwpk4/c4MLY7Lxn2nOXTXy8rmcFOufjzNF3BRUFG
Wi3QaDa7UuARckbyBdkT1wv5fLnWjIXpLV5LAzJbAQWCsel+BpvUquVfY4otiObJaYPc7xM4b42T
i5LIAblKXDatziBSGjNHkntqmr1nDcbCmKWioP0djXHrifi0YhHK0MA8vfI7iENEhOea9NV6skdh
ieexRi3BnBkS3DQVm9HjnqABS36n8AV45GtdIlT1arTAPeOOyuo3lkmqM4WaDHC23y5hhETbmgI4
3chCyYC7R/1YOzd/5mCVgzmmqc1CLlAmB1YIfaE4df3vzyOjZJTscjD/afl5CWLmV8flQlkLTHXI
ew5A8IjDx+iGKHBgvZZDebYnZUE4/+AjvaiXP0GeMsD3fvJmam9NSCW5x/WPT7sh4KHPghdzTUJV
DQFR0Z5ykHNJXOe8x8MeFw/InNob2ALnU7WuBEfZsQ116X/DDdfa0V9P5Oe1hPW1a5rJCI4rqgCh
M/ZRnPr4PG1eOyaEM84h3HEHUg9Oe9Xr1K4teKnbNjpF2QxR1kwO+S6zyHqTBorbbSLSDWy9XUu3
7rv1rdG+GYnuYsPSrC2hkXL6Y+TRgI8D8Rq2MHIOpoEmFNg6lSxY83Ow1RER7LF7z5npWT4lIq77
0GM+Wf+YLj4BYs5fEOFKG9h436dE2rjcJFwyBiP9rojqeyj88QrqXndlc8l6odQu01dyeiAPBE+d
6mprkkuR3+3KMU4o8yY6yEO6s42OEOcNBEGQ5TSQKD2wyE0oCHJ4Pm1VMs+3o2hQAxyKt1P1IX4C
Yl60Rv+1gSgycD4LzKNY1268RjJq6h5x1m1HLfDisOs6SZSLySaMWygotWbtOASwU3Gx4TqhRGB+
o4oRfbePU+APBmGgXmdxLKNcIWuyZuYDD7Ui+RorjCrOQZO1niyMNertrIVYcdWO8BGNDu8wpThY
EVesRVkpyeL0J5Fuqb4asl39uC7tcHanWanVJ4IqY32MTv2nRs1HuX69T7rgEPba4gLW9l5oeXnj
4DT/tZvBkYdfMQLY0ft8CiPLj9ubopPuhybNURLTG0inFJN9JP7K5YNTZtK1HR18gEn6TDu3TK+9
BSvc4gv6vs2BXstukHELxFKmFQE5anXhRmVZeZPoXaYoAY2c027MkC6ebO2QW6o3UDCa6Viki3lh
k+0EyxUAfYYn2nmLVIUzhOPinbhdM83LTtSiCiNn6OsWDtleMn1hUqUsAxYZ7j7nZPPdG8HJyfzo
5m1sQ/GMzLCOCkaHlJ7mHzIG8fGdMbeTHcJqSSmSOeaoDIVw4VQIjHVT2QMg9qOimpAlJW57hnTk
tDiQkQajsv4IxF9tWlfG6506AZMji83x7MamO8BEAwXcNK/CHX4zBjpq8QeqWmvnvyJZC30Lfbfl
2FhbIdJ5wC5XG0GEXm/2l4S7TfN9sdBfl3wXa5npemD2JjqABrlCBWZc5htJWqeuoaeZlt8MMVxX
YpGgr1BNaK3uMKxDF7ovcIP77yZEaKVa0TafZd+AaGQ7jPdza+5ErCksPOKayBSSacqWBjFXcisk
HSYSlp84akO1ZGlc1cH5/KXCvtaJ2eU9jCcTrfd43P3oiGT7FtL9A2vk+IAlQHTTpsWEw4ujPJnF
m9aNTgHn1rqSYjop8RUSomaP8EcLcnwWIr+3J5UnbS3h76VRUKC4dqxV0CvtJp2Y77S3zCxzWITK
QZ4i2niWieReuBjqbircDLUHTgFGrXQo8fxdCsJ0IhcFcziGR36CkJD9z9qNifoidEwQYebTPTCc
13iNIDKRepGBzkHOENFzrTW/i8sPHEfbzwTsk0fL5P8rTEFMDTs2Nk4R3RuTbzImJnPVlFfUekLw
KmRLEAzPzallQyt+3PmDG9q/kBwlay13d23mocL0JiqxZfjb1O8bNzGuus6bUfxvDqLfk6/EIyyb
JFEcegf+YSPUzGYimXZWogcFz7T1jpBtQlc80U/YOTS55+1vIdx0jVejTdgs2cjfHrTTzb5YK8ez
NRyCZxdtiJ9Z3r46ly2b5ccAX9GKwkKyBkM3WwNY9n0IemrpJsLkETUhdxWZTxFPd9BjEQVrGwD7
7QYid0p+Gk9yr1tpjQjO9oNhEdz0/QbTF9MFN4P3KBD5it/mJ/1J/+9ebxfGdUGbf03GV3LOYBg6
wVcFPKtfoGA3hQ7Ise3emYngWQH4EvwOc5Bzu6KlrmW51aJSonPrhLHISYS4OqU3rdFa3xsiI58D
K0T6twO8DE6MlIAXtmq7ns/jcG3HXdCDjrCW7eeaK8aUhFUVI7z/VtC4XNX1BK8UM/Qb2lC4eMf1
qJv6FAiNzEBHnWfzR5F4RZxLqpXX+KnNdXdXQtG5fGqaI1aWxtbiH01A5X1t4I28gzj2+sbaRLqH
Bj40h0aa0d2dQYKwQZW1sGEPl2C70cft51gkBPhCpE3vwXMV0Vrc6qHCOLi92HHFoF20jY6K+B0d
Z2YtHVVbwdPXIX4Yd3G8GA4X3cf/I36LGwCLDqnHv60xq+YP3j4/zqTrb2d6cmr8WsNXG4gFBDPs
jNUEbxdbcYZnGtMqoSCk+0hcO8qFa+g5eWBbm0+jQ2TihlcKnIaVue7hpY95jS3LCRntqgne5+Gp
0+6dmh83edrt5qeIpk8d3+YCAxuXdWy+ixx25WPwVG5boYWKqyMO0Fb7DEjz72pSHjOeRbgizhkJ
ZV278QPV1fUuYyD6Y3fssl5BnzkIsix70Ug6rYC91ojODRuEm7thXtYIkTpPMfpy8GGC/oHF8U/1
rllxHxk+pgWGLfdjkMqcQHjjLedlx81KIaisni+ZqnDldHzPXVgqEvdxRdp6ARUOn3+f4y+1GKEn
3aZ+pe8TG3bHcylX/V9t3Czwjr2vVbqSoXm9D4kqfA1AH4+hut6cbHpeTunNiwhZW41bIGUH2758
fMU/LLCPh/ZfNHW/FvrAy+gz/LurJjmhug8lx+cpDIBG8PpUGKrnwuXelawJMI8psyVErDKxteOW
okFZ0mfwh/zkDHk/jczOrv+jlqX5sOFnWI2h2YHxzvjcx8MGV240qjjVj73f6+7tQgAr7RBP/1nt
t+h8H67A7SNOE6nbcgL5fqgG1DHuDMFxu8WTb5eEDPxxlVP17Au6knkB6ptqp32q/+OST2z1uOeF
tnOCnudmTAGJfSBZ898DJcdaEAZgvtTNrECGyCmqWxc37OKgn5dRfrAuCZVX4TEUfchuz/ihjzxn
ExuZTngYB4miyknVw0k9XE4lssvG81tOUdlgOnvGTOIjXX1RkhAyJrPUsgDmVztL8EOP9rudRIut
oSTIOHe0aMalRD+dNsdZCdtoDKSrSJCavFdRPUCUMdO+BTz8hsjz+WxgUsx0zRrCOeev1IvTWBJ3
8lwwSBJG41h9jewE0aFFivbQLBXmZi7JkzhlJAXCwZvAKKD6XehTLwAxqRTKUAGSGST4FBin4Pa/
gnC9DkxEfKeQ/xW1nVL1iDfZtXydU1iNNH3K2LUcoe09lAH8wNwyOYD9jDbL9Ue1q5cLCZAgnFq2
HIZUfhAtynVDT4Ai1+DmbKmFYYqzjjiCmrbzL9npFcJZKExN8D4FHegzldyQThLQystCaBR2YLkI
7k1WZR0MnouiUZC8O5Mcj27/KV1bnM1tMbK7ZpMUoJjWw/WzmDizHyxD0ChMC+FzLzRjGfVQkSjR
hzyEhMhSsviJ3+r0YJDJs8vzjE/DKvdTF9l9zr7x+jWgA9qtMj1w1VjZDwEHcTcINw9g+FkJXLsI
6iXAdA6XidyEnkuOeCjqDh6RUeZMJm5aAflsCgVfeZm/DfIsnIsU+y8l8zMLXg4lAHEPdOTJLdgq
MIXTmALyLOZ+Tk5NjfErEZC+V4COoY8JC9jh+fpgZuZWKF8lvWx0Mq4fAXybW3LSeHIlv6+dmpD/
VYhSlK4+XMEg/6CbyX1cK5DgUtlnVKtuXn0L+To0R8QyKNQnmNIkKKAm8Q8scyg4lKuORLRdWdw8
nagdv1s2/WUk6Y5CSKDcmRs8BqtiZp9eCzt5FJ9R1XeNIaV6dYF9fWBOD3AN0yZPdk31hg6TnBtL
k7TOfSY/GYTJtpXL2ZJW2oDrio7/pnsZSPnpPizJHxo7SwWqUJPQKXYIzK98MjOM9hSk9IQwsigi
BosIgcL1+I4wJqHyzlfmsIjjU5SXLIJTSOo6J0095hLeqGDJHdPgRCcLJY2Oh30v7DQMnp8nciyh
KPcN9cS54v7LWLPLTGMexInJOWEOclS+0pBX7WHnwuk53an0mhWYNr1f33T8OpdJVoski+afQo6z
ZYgSOjZull9uwLD68P5oBEKqxrfNo9vy4Zw4Qmiq/S3OYWqktB5mfxi6n9GdCevAUyxD/DIDTT3h
WKTf6mMYr12IilPWaHkC5aPFPeHFoH1aLsjINsAGmbnwtXl3zVuuah7htHoKxE2HNa0qxfZzjgD6
UBNpYQO3rLaCEElAP0nrRmMJYzn/RW1SBb48sJPsdF/89Z5HkarnqOj6sR3SAx9bN1i28RsESIAt
IttRCS5BMk9LUJuO1zgk+//1e6IdrKNiHaTNu73I7nZ1pJ0ZfytaMpEUUaUQfAh3GW3EDg6atbjx
e394kFJaOQe27JwWR66PASDXz6hpezxHwCkemC59mVLXNECx3bphbUrQt5EUxoUFzsZXwU6twMQ5
PpiRlY0TzpORVB4sUXDks3YEgAzB62xcL5wYUCeOq7XhEBscIaKuhfNmanW9ewXEi3WdYUc/kHmR
mvh+6ow3CLE9alz5NHadjdqN8nBPaOWPWwVKJyuUe2DdDXOObyXFW0Gz8q4+ozxrm7ELpjEPuR5G
X4UHxG4M30gOxs9RYF9mYcceyoIfSrOpbWxfNXR6W60uAlJT1GYufKt8pQVUs0Wx35+xOYgztbGY
NoJ5szSkkLM5HlUlSlIHigqF5zDsN5GGMLK9SdPGtaQDMtDpTei9L0B44eHkF5J/ad/GFRJdMsV1
FgntY9GK/DKCi9BOFqguQvyPIccSNBBgSLB+2pahtX3Id/RCmPeI0dnMr3YbDTVclkv0CqfOTI0W
/lV/pju6ImaisMgoydlYt5UMsW0/lWyBfruyYNhyeaN6SfX2sK4Z73QCDmk7pGh4wUQ8xduchN6T
Q1VR3+8bI7JO8WbYqHEnELz+zagbenNRMNorkzmoYD8xeG1Mqk/vFfD5OjhhIa8ZfP8s8cS4zIfd
IQgKNwrj6s4qqXm9P2cB+k9ca9ZKIBI+E2g9pMQD0tJN2LuuJlY4OmmnecuwqCaouk4SSA7OBxfn
YJNLXjEy25GhIml2Nh4Aclg6G2GGXbjLfj3AQR0IdBxcRnbz8j5uYoxHpLFuSf06Ql8YWMx/hCUz
n2roRTBefduCKLxdLEg9hmoE6lUQu4rnYyHTi53qPo/btAmpHZfe2g+acLZ3ztgcxPzHX3Ow3hRV
DT9qdpjZxyik/LDjNz9BTCDB0oizojCygJiopRN8xwsITSccCsv1uhxctfK4uAg0N3YFBZlZGhBo
d47Z522q7FGAfVzuM+1U6j4hgpHzF0ZsJiUcLMF+auyVer0M2FW7ghWUxuJHUDTJEkDr4jS/yh48
Z2/V61HsBxX2dTSOA9ol+BejvZ5pSIn00Mx6OO60SWqFXIyL3wbbe/llRpzZggkUY3qtsL7vEzhp
HCL8LiENYLHhGMQilfsudl1Iz8ZWRD1tydhHQD+Ufb448JBQnMRTZBAeRcQzKzi165MwEUnnoio+
UfLkuPlzWJXhgzp2/7akUqz7Ljf/6RkwmOmo7Q9NISAWmGYOasyD9us3m5XnlXnm5twRaZcwQE2o
jVk0r7RMgJ7ck4gJRNbgZEj76O53Xm5DQHiO2qbJoY/u07QwmvWZfTk6dG1f1PmaYrTFZb+7XdQK
WG1r1POkIHRGAR+0w8YBhcWSCIwyKJGw274nnK2PwRIRx0V0SlDqRpc03khb8cvcCle9WLUenX8w
a/R0ke6vjsGlDK6mJ59r/E8PeCUW9P0ObIsrP8ufb6xpNZUePfL6qsPqFvpj5wo4xk9g1M8zF4xm
GeZym15+u2IF3iUJl+GxAZobDhoedXOs+jEH9qezsXkhxzfCWEVAts7TWvNnGD9Fksn87Uz53LiN
v+im6v+XVM5YX/FRjI+3Q2Wv83fvXWA5U2qKGSHuNgncmVqUo39/6liTpivD83vojGf7uc8HyNlx
/ytu/U2IgbWcdscyVzR9y5oK3Nd2JGYqS350nhkT91bbQhRDTKTlMEW+37PddYUssQsvz66Hnnuo
zcGEksRqwEJmvgFSIteyW0FywNURXoBvoswP4rOPLGlzUs4vuQjdh/tlUqRpXBGmx42yMygWLNHi
terNZonsBfGBBp/VPUu8104YuB3PHz1CNItetT3NyMhY99uivRfEgUta2mpal3Vu0zeGJ0oalDlH
BFBySPF0z1EZSNX0uxZueTN5SnlKGzHksZvNui8zFGbXAUZJph/qMb0qfdtpOds/UNQDMv4NKMHS
yxaOkzQODx2vEvyZjm7vKCWVczUO1ZF0DSVlqRAI1CrtcV7HwufK5oDZXY6hj196M59cZrG7ue6h
4TsJPtWvRweZOsyqHj0q0cvFuxBJCcfCxhnRYmdSGv7ijIf/yo6UZ8iIKJGLWkT19oAK34yKCc8o
7WFL2pd+BLnP/8c9vglwhYdGKgLQJaL/YoTqgSC9JCG+xQNB2+ogiiKOCY/E3ujFLpesm3t5j0s7
T67PB7+zf8rZLMReZh0HBenkxTBSAYWj9qukRdeTHAKhXtKKrAp0aapBnH/TOQuwzLXR038s1MFd
3AixdOTUOV1zHwmSdAwoNP2i9IcBkF5ZpLoP5IhQYNi0WAOAKH0m4UxMwC24CArAXalZ/Rm+3Qv2
HNcN5Jdw5M9eV+A/EYqwQKHkf+9yE2NsZmk3w4tdEiuexe3kI8YaKl9CYWV0t/eOlu307wwOqDRj
xLDOFoIxCqK/zbybUCLJRcna4Xlx8i2U8y++o5KONT7zs8sT9jxruo+H/IH8P/4Egc2Q0lg7AP8M
pdwHXfVVV1ZoWk/06iTe0rMz7KyfHAurLjRiI55C41hAgyfovh/Xd0NprIp1aDnffO0qL7A8Vi7y
HQK489t/WVvtlrvkg78808Bufrfm0yL+ZmSztFsQvM9pJ9OwAubRbLr4p2LBSJAlDSo8wvJPnRLS
XgkCOK1R/GKDYQMdkk6r0dFDnH5MhG/kSJJ8Eq7912SdnRU6MiY60PLiBuRwo5YG4YG4CCIYb845
MR0+D6b0q/CfnR9JdxJfavSQ1sXDHTo3xIcunDZ4esWcqgiGx+RAI8mPbsiiI1mw+dYR/ONzUN83
RNsEuytue1A2MmXT3CHzRV39BzNAaxo6NvKk86KZ775hmzSWYX9OKL0/cF7oCkMYCuw5keZ7LDO6
X0GXGQKYQ+WjIBREdx3WwxF9frbCvmdjeUOoMH7J+AUzi/afU2PuU/CPgFzWDwTC8XyJBHpCkx1k
yaK6DnewBskBbyRsWkaAT85d4xrF4fvkw01s0ktpM7ftrVb5IimLupwfpWJNcgSwt2MHei0zjGMp
hOLNUwBRcbi44wrsfbbbwGHgenQ7XjTCfr9FbIctOs1z/L5z7zyfFZN8/7Kwsv1UHavXn0+Y6wEr
P+oENM2YK8TOCfxgpasCoYGWWPtpFPsG9UtY+tRsOWeE8W86j50UaxY/ULUlarwY1pLdvZ/gXgJw
nLgV4rSRyTDAabReUGEb17F4hfQrX4HdJQg0Ww9XSQY5YHrc66jOgo2MX8YuIGMS/YZJp5p8mTWc
Lp5NDY5oXEhXgqPKBLm41cmOTmO99R23diggjKjR9Hbgdeyw8zlHghc65Gvj6Xz8a5RilqNwVfxV
E0HeSzT4ECVJDu2g77j2IuMggEH3ow/LBz2QEAR7x+wyDl3my8OlnB190DldW1p8VXMa3bukGJpX
6z/P4rbpyxKBcKvoCWg/yQiWLPo9OFZGuiuVjc6zyrcrTISFTT2xc4FG2YEAjQwHwpV1hXAk1xsN
F25BHuU9hducGx/K9ae7F6xESxdKDlq55LgN+ShjdHN3mf8JgyRK0J60wl88lGn14wB1OSrFAWTm
uwPDBgOatMg3lKwbIvHOCGDnVhEqpTL0tbvtKiz4ffIMz9X+RrftDdv9qer89Pda8fNkNBW4E+in
DgND68zLXTTAYAFnXzGn4jqKr8cYFUnH9cxerEuX3cyU2WmalVbK6lPEUTvMxAnSeGkKf9mP0f+u
tS7q+o8PzkyJPDxrFhqVn7sRLX2EKu2SXuKWiKoOCVpl8AxXXVYHZVS5mJJ8FUIP5fHwVH7bwQ4g
h4EgvSSbFvB0hlTHB8E0Lbwsox+KBQS6uTwHP0NWCbF+llKzoCaeYbBw6521sqB/Km+wrwNByGJU
ZZa5Tj321LCVFsTO8H5Qw5urzdTcTN9QUnFQez7BJyttNkMYK+t/2dOUHSw+qQJis11DkaLjl0Kl
w3/o0fkQZrLO9smoKWBuGiik+E6dQVTwIXaJnn5ZX6ne/j1mP16RdVuP638rN8iNZ6LIJ8xKWlAR
BGOHeCyYkg9yT6ycbGxy/Mn1juVI9Gzo79zpvZQCDfXaKl8UKHYaF2E/3p68K8JmPJgmLp95Q7MR
hybbT7UKkSUaWlkWG4bA+x46+w9pwk5bKQ0tfROmlMhLRvFgoRh6wrOPjare8CpOlhna/wqOlI/q
UJzMtAvMm5IGpfZUiGTX/OdqsUSkVfT8vbDbhNWVPt4T9rBTFhp46B354gObKeLIyCgK8HbFaopm
t6BnWo54xer89H1O5UAA+LGA0lwQ4V5lrpEfQ5WmVVryJ8U6wRt5ME+QJgZBrBQOCe3FUFMsNfTq
I3PO8FUrfgf2ucYs04vaPqwE8P7EUI5ktTM+L2eJhm4gXXi/yAE2/v7EsK5xBY/EO42Q3cYTD2d7
c6Y/ceok3WYl2Mr5jVA9AT99R2DkaKfXZ4IV7SmaTAduzHcgse+q/iKkWL8EYV2tUFM2AXv/UWKG
0UxcwUR70aLCEte8xa4h8jvUHL2YrNsmV6XTKfJQ2OEMhQCKLH9cOlx9lT6uS569nxbaBXudScTP
x8elO7kZ0Ovn37WKY7kdQJVYxWfn+D4dfvo9zwrlZgDTVVj906Es44MxeTQ/bwbdPVfLNCmLGtgE
xZWXKFrtpg4cmLntklyvya3SbPqgESY/0m/8w6kFsum0KtEEbxQfWBpV8m/sd+D/ZK+2qkW7rMP1
T4O8oAZuJOMRnrJ0QkOajbMHnvpJjtW+CpC4LaouO+xH+QeiGVY3lkJvSdBvfFgRXcqGSc9LWjAE
gGfYb6AlrYdahNfU1GqkhLDSt0UDoTlhwfLwiwVMQsYT/7SCufAEWzby7mttgDj0Adcq81clxMWl
Yu07Wht4jucygm81b7/LDOI3D+m9EcuLCfj11GDgwqU7vx/UQy53RWXcAs5Yt4b/LtKrcSzSFHXf
JFUMbmsECJc1uv9HthbJww+shb90pyYhh+bZy2fY0H0vkVNN9LWerFjm+gh0HCPS5eopJJa0SB/j
hieTyF7qdZ9KQHSYqjmOTHtGvFG8qP0VtFeQNHWk2G/ZZdRTUZGdK+ruQCE0kpyoyZdXQXAfFsde
lJoN1ZfH45SeXl1vkrUEyl+axju8PfHaTASQQUu/qenOgAa6saUcz1E0cIJ5LG910OZLLu7OMyMi
qdFRqH+GFCHC9jm1ti3xYWGScx9FjKx9nDw8noL83uyTsAqUN5ijv++5rQIv7BeVH+RYuhkxqTbB
rcw/nC46x2KrNj4m7eLmsA+TwqSRPuFZ1Ww6votX9DDsIBCZt8xuS6NucBX2CKS0fDzXLHapo1Z/
C4td8SnHNVbkyqQEMsOp+nXSAsg7XECUYqxqnVa9DLe4Dj9Rgd503rO8nEpiEesksY/cqFvLMIK4
DR+eGfPSmjI6Bnbtv9ZhnqMkBZ6HGWr2504jqifwuE2OWTZK1mlB4hxeO8vhyb2T28NUB8jcGMXL
LO7QuGZTsgeAR6rfoPIdQ1jkbRIml1rVn5/wNgDSwXXZqwU/ziCycFxGazshM1VxRVVk95t78k02
7jijgGzPyZ6Y1TvIcqwwo8OPgpyJ6BPPWA1cfAP161klczyGopcL39ZMqZY0tLn21vOwWCFphrha
PJU/6eDozEddhl6XgH5giDSEexZw9gOrxKNKivpFNfqhNsc1oPLz/tnGrN5Gl4UGRaEu6xejGtRT
i10BlMXdS55o7aFkOat2heD+Us7dom6MZKQkVghdD/T6Bt+BCtrnBSDe2mfh+yobY5jY8EsaBpTL
FOMbuuJm37JAvBY+TtMrwO0JZUQdDY9Q/7IFWYUwLtx9WeDjKcQGUcxsUy8JfGs9y4K4vOkNWVmM
I0tWR0snRxzDyYsxzBB6kzYGjO6J3pjIurxX89KBvtYRyXSKGQX7s5uEYm3iaIiGZw6oxE9tMbt8
oZBY9uPEptBc7uqRdZk6fKM0UfgHkdzCHQIgWMvVKyqsMD5pCsWatAJFHph0mQazydE5qvSxhEKn
raNS6LCgiDsNuDnDwYtc/wnVcau+5mIRunyyBlt5UhJh8QxG0o/5LSByvB9Vll1Yt8Ar7diorDZr
nNylZ2yg7+5K8BHgA6dSa7eDk0a8hsknGpMCYteaC4AOJ/5+qNRsNRGIuTkipsF/NVCgaMnzGxye
cIMq5T/YySvFdcyOeTwCahFuXp5aWhM4RnGW7UbeOz2rQq4BtT/nmaJT0765v2UCfTLq+kJtotY4
Axz4EKTaajqzE/g1IOAHM+84SWkel7UizvPcjoS5bd6B8OLTK62B6LcCpTenpkawZo8drVSdTm19
D6H2LzdqN67rz12NK3B9/zFYZ23SQD80mVNshIQd44pnULUI7rF32WnEm70Gh/A7rF1WfAkpJrVB
rAOKSsq+L/XyMXCWZ7NQzG+yw0iWW36EsSJhwPULB8uEMNC/of6Kk7YMdt1sT28B1+RRH4qorJ2Z
Myp4iEa54TgdgfEZ6DpFjq7l0yzGSNxIUeeMP1bvf3Q2sXQtLHKL3NQdRVoTFD7FUJgOk3+xxMZ7
AeI2JM9//5ox/c+uPLob+gABXPStV3NMVDZn9U4lk+gtlJi1HCw4FY+GaKO2Z1Nkv+xEM8Ojk+R6
T5xnPvgPjEPtjOC6O11f448TFGcQBqn/RmyGolUaxUZroMVrpq+dU4XPiWyRXmGJwSND7iTJVI+8
Rq7WLraF1K8R0/hGyxzFuQ7vEVT/CCS/k0blTrbbCEcFTSEcNYAF/i0od8SYZwnThWYFsbgTlylV
82sMcxYEOnHdWmpvjFJSo2sqsUpn5y45Cj4YgPo7TVvPBVSFiu0lgboH/YDd20StEdxH2TfYPeqL
czxyDXUs7YbYPggxcAbatig0ftCa53fsEg/xCMTNH23UrCPCP//YSee52X/u6rbCgFBDGYFauNYY
AVOLcztNfFsbvIIStKEUIHHeLRZPfQbwkcDHsEfTUs8VALPQFMJKIjCbhzTxff74hcM4JlvEQ/d3
7cbj3HAACSo8Q59nhrI0YDxX2SNWlEqiQMtlQ6h7bR7kgRBI7pxKXAUpCukJf8Vc/1v2x0fLEv2H
wz8X3Su/T7vL9XgLluhCg8qc1HRlQXW0qQneoq8hReDPzxVeALPL+lbSrXUqrOlV7IxWXKIy4lVM
eyx9WrzR8jm3EASvUGPW5DenP0LVOWpp5c+TN2dZXjJlQiNOOIRWmZpBfV1psZ2/msBDWZ1NBgbX
YA4xDBRp7gUr96gWAqAdMzXaraQ27LxW1fV9Fh28NbYQirj5+TriUTMuBIK9l9O9boBUv7GgfAW2
y32jg93D2Nyv3l+P+ywXBR0sXdQlLjjicjo4unPugKTZ1UnTWYaFBj+rmHSiZnFCrAJSFpQyMZXg
i4XJ/m93xaev/lUNAC8hit3OR+ozmjU7ymyUa02+y8o3A4SSBhIq4jaFk7dhGxWuomFslh/0IeNa
mmF+XvEcEAZDiQuudw3O9ibc1iSuv0ybEGvHefBuhl2qFT7VLs1ZDqlcpzerQZKCXuM7qcL5f4wl
WywT4slR0F27zrzJJYCRfsyBCE2FRR/Q8+VvJFmwMVJ9cV6qd5pHEYULkmntefWMrettlSaL8RCv
O4vRgF/upHDMMM6U4p9vU82VrpGsWKx7zUnzx6qnXgLkn2BbqhHADPT6AkjlzPXoubfBMM25WP3C
dMDtmLDKmeXidoXiZpvszyuy+9SxwU6FhiDGGUpNUR9yNdtDlfK2B0fSo0QPc2s4vz6jkzp7dvKr
lkRSVidwgfY6z3rbQgWQX9ZcAO/ZgvSulBfaYNbd129vXg8ZkD6c3JzzMCg1HLaFj8tRztIAMGaJ
zpK+rDPUz2LITcMBIDjvCVUTfMSrn0ZTpDPaUeoxH1Xztns4Ub5Hu++WJpjHliyxaZAGX86bX9Q5
uBFIfbqUX/c/qKCbA4D+JbY7WpnO9BYNxCRK57Bttpe3mtk7s10WLYV/SGZmp7ur8WM5mkxMru8P
6Kssi5wssgs7X+QhdnJOYC1BPlUSJ2joAIn6uT4zhHVeijDkZ7gTbWVWg9wCHSAzjM+5sq7w3T74
r01pvcLcvSytlqWFHa8BKCe+3OVAgNPPeWlZGq5FN00dZlQi7dhy7MzAC4SIruOjAO7LrB2xC8+k
GrWZxOtdv6oDFu97Xkb21g2/Pz60Er4J3Y8ilnzw6Nt+Bhv3gl7v7dxmirXXGOZomerHlfbzi9rJ
2TYUY3qrrzBbN8VbaiM/kkIYdkj9359zw/NtLEKUUqVFGLiROvbcrDmiD7mAnNYg/sRHJ9eKbtj5
uzPphKcDs7u7IXPzaPTxEabZCl7jxv1daFLtkjiswckY7jkmQlQWlkMLEN/j2KXUtdJUUBc8WThD
PToFZLh0HJ9vNHzE97/JSvmqZfcWV6L6uXbUiszX0yBP1qRA3eSnoQItVgNNXz8W5M5oPWQUNe47
IWj07brI5xW59vdZZe1YK9QvEWMFDSZUtwrEswGl8QG8t4wYjyyNHIIAmplfzCLCO/KzvWRybXHA
GHOAEPuVFbUENL3xdkgnKOYTRbvpP6bIK8PDelNI7zfFh1bBYcm8J42qz11T0Vcrr47UMVnKVKX7
VwQxh/ykfa3/JxFCCW9z83VKvtFSgXa+tTGMCV/glg12bj+4NwRHIeGJBn60vWRF25gzFzB/Eatm
2Kq6FQsBa8vY6rMznNwsnpVDxvNE/vhcMyoCwzu+JKmSchPRMGdFnQqS/nV49xeOWCv+5h633ijb
YEUdpCsewqRsQAlHOnBDleklkVB0vm2xINgJZ0moA1K12Ai4GpIkWzOQBXxsLqC8MoP1meYt9Myy
wFzeuB/ZuE9wJ8oPFMp9gtVNDeXAuBj4kyXwb/6iRnG6XbGjZCSyzdbBV/t7M2u09g2Uhn173Hul
rY8LQNUfVOVE3Gi8uEaai5mwFf9OmLDd8iLaXcNn6k180VgNTUfhJOyoDR5sX+XCW9H6mW5K23mO
uNVSq6FtG9O4S522yXe1Omk8P6CpQEA2RBl+jrsIjtkh4YlkQ0AlvIiLMW1Hui5Vz0kHDYZvrspS
pxyuUAJVO4Y/x2M+qfuoXWF3B9pmHLHDB1qsJA0YNwofopzn4yUvYDVpITfa+JtROyMAmWYDkdiK
jkxekWLIayprsBISKn9gozP/5x0KNCRQXkwuC3cHI+JKQ5zpq4IrL+qR4FQBCLx88f8jz6DtWR/Y
e91L+rG1rb+lNYaVNMi2mtuKdzp7/XaEuyEJGwxfkTFCBb0i5A2lsxV8PlA+8zyhy/u6TfIYanf6
IFbb4xJqjlWKV4hEPPexIz0VzvdI1ZNiljfwr1TaqA3dcGcp4jWNkFH51BmkAOp+6LUXm0KhdQxN
/Q8PTzE/qvcp5UtrX3E96Rs3if6hQTvpue3ERn5OwhxNgvOX9bduG1HkH6JApGWvEg+Wu8yAsh8R
0RGIGrr52bqLWQqthKSiC2agEoAxQ4mtCAp5Gs7iZ5gAgis5wUqtAk7TP6AIZQ1AbO2xMk8ltHkG
d/j/PBIhWEDMa8BjOmhsT6rEEExYYl/1+mdlVl8XttS5qXutFun9tMzq3ynkpzVl6JrG3QHdtTEg
Y7b8f4nBVrcGIeNSavSEa1dJ/TDjW9vTL3F80qMsWlzAYR9ZtRUfhEcz3j4O+5Zg2yHnVP6lQERg
YdbNlnIHF+KqcCdcI2s2LF3xj+vY0uXWMHD4OrUO/EKxa7vy8981EJcRFx9bATKAO2alDOn7fRHN
7dnFCMI+LKeVMD6Qo2VN4UT1joAey0qGylKNvt05h+KPMa0vg9Ed6o8z+Mzf04DQnbT52dIQ4rdi
c+05/EpC1v+tj6x5gkZgr1PtqEK+FWBcqHDfAYyIQ736K32s+3g79w/dAJB1L3gGwuXgc/7bbbQC
/WOjHIebszxzldO8y0vyNaxy84Anw3lYK9FBtnWYlHSWf7dCMBW88AXxVJK0cCjg/0Y413fbRTu1
GXJmL9bn3VsUa83AGB5ev8fEAdGgOJrLSG94QEfWX5jqO+kymgdfHL7NfTscRLCcteX6LmXt2i0r
FRAZavIsx3r1qmG0R465+0n6AHeKMo2KvPe7EKyehReGdoRX1Fd8tNMvVteIV/WT5u4Tkg5ZFK0X
sfvMSFQqVtvZRkdAlwLuW7Is0pFKbaVBiOVYJi0WXj0hyyDE+mhIFRjB1P5cUs4tHemDb5dpiS85
VxfFT6v9F5znQI8UQmdyPy26MbAcRjuqn+OxP2BrOpfNltktgf0rLZ51WBpt9JZnVqm7cKylOlgI
XU/YyubuLKdyV21eASIERQGx/rbmmAEdom29todm+2p4hPxQKDxdDzrtbU2LDYstPcA7HXA8v1do
ACavG63rClrwFoYmgVelRIkGgT2H0JGbuBYb0hPj66GXeOoe12K+1dEUpYgic7cjF1VzTgDCIl38
xx6rj8v9u7tXXw6qRcU65T4AT91ZFgOtcl0XsGpukrOifKMIOl5MAWFlccxCgrW6ts0pieGsfugF
zilAGQ5Ujghg/8EF+HpgaGI0lgMGxXm27CkAXbQKrq9ey3fg4i/nrwpaCS2DpnNne89zD9CBsEnt
UIuSla9Hb8qy1BdmWesYUs/hLHnyarW1++QzGgjYkmEt9FK67QcQ4p3x/xpjmF1aLtXX/Y6iqacm
EjKrfXK5ZxFcCXb/A9KK10K3uY5mcf7wSIHBaEi2S3NxxMyOcXviJuJtsGuEXutQxyv00os9t6+g
YqRKJig3KlQcIk0vHLLyPiT4BzSlM52/WGQW7KYWWaCKFdfbOhOF1lRQvotg8cSpLQYr9iErWtHx
2Bs620ight8vhxQstW3W2MZfCarshN+TEg7eKaa24Ber536xxCt+be+0CPqJNi2X9BGr4GdcGc5q
Z7jQLGhEoMGMODWuMG/b6ueEf9oo324XnrXvJXm455wuM/QBBuFR45KUEd84Kdtivc3gBsWSgO4Z
FMELjgquEQ7iWfCWxV78JwDAQDfn0X6/ri0JXgaGL7VYZVtEgPXXN6d94wr8/WrzdryJ5Y2ILSw/
5AT2C2moNSM8YHp3LbSWEL/9pIvPbCx04XkJxEIrPB1GEw1WyjOH7QhNDfpb+WgYwU9pMVvhR60Z
bnnjQ2aKxzraZlrCXjnnzUe2/DcI5ny4XGx+Sy/vt4yPWiEojenDen2HfZ0JPaDMR5AHqmQu2VJr
3omvjhzrLa46+zegHuXI3Q/Nz0b/G0DpF3jzDsKBgmq314W0ckfEwKh/bl/7eMOL4GNPk129gfqo
S7amabP83yX4zO6bAGmWeXtIxAC7DCASyD1Es+h55rbKPHOtitYW3qrudFwvEVxjVP7QNBr+tJ9K
jW+MuGxkKY7owpb09MuhIzAoyeFrjoXGlzjsjs096sEasWpJ9udzyC72XOplhR5p5daM6AdwY7i6
R3I7P7/NmiOZWgUQKDsi8Ln2+N/QQ6TWTLTzg2yzPBtXzYUOdAug4IsebEL6zuMx5xvqVdpHnbeK
WJykJcwbGtp5UFqWLvlFVlEA5bltBeVBypij7Shox+epvfulbs9s3Oc+ICby2ly66vcU440Hmbm2
Ds4baTbi5C/VSL+a3JpJixct7uuBVlsAaJBw4mLRl/5Sv944h3Xlbd0WqutzAbEWLrLhbm/BiEjk
OXtupaC2HFQpuTMdo69em/UqH5bSkW5aiVRx0RBaTRTJP5Sl5nwO4isBqJGA4k6wmn1UPA1nMXAt
vXikqm6gVQMTnu9OpG8rtHmlJQJdtNOn3EFLZkZj9U7jP7YeK4S52OLBXu3l51U8qHOA9r2nLRx2
LzkeJBbdECTc/fETsO9nQHl+2lWxWMrAf2vSC7GcBzPkYo+sHYoWubOCnbaBCqYQ9IQyIs0FyZWO
HzYuRR/+xqqp0vZsgMNHIKhZjfbhDdjUePbrMe8yVMobl9I7oT3c/D51+wDmQkWi4xZjN8N3PGLp
4Ao05BkiKoywCHz+lsRmmC77hxMsDgoV3BnDRKffUcUgdUUfGysgP/iGqM0gjpov5l3gNoW6kzwX
gezhNSNwu+HXk31HQcg8rscgjAQ+/RZcqTdYkuaxRYFt+JQjmCoKhbCH5X1O/8s7TyQDo41zy4zY
u8BBr+mAuMYLSZkYMYNHm1ZUw7FR752+s7EpcG0l/ngnuYMvO7rk45NUP2PZ9ogpulYVZvZK2N/4
yG/lEoYkf8dyl8XdtJOmR58bAkfgrubfmpdKXE8Zkkb3xjyH68XMOwxM0n6bGrUEXsm+RirlD+Do
r707RijQ4gpDMPeP5V87yeR1rh0elIYyxfN9tKXP4EuQ2VtpCdTBfQYw5IzkwROQRkj9IVR0Ffgd
pIl1XD7nlExHwOGR204UwyQe1CgAunpzVq93XdUEySkqBx7fpV0lCJYE0QAIFXTqprb/kHLriVmp
CXnWfvrPdbSRagChYXXSJJ1TEhvhFjPHJn6v7bOje7SgS1/nX6oWvszKLMP9aqlhzQJaQshnq4iC
oAQkg3DvPuBzvwOEYDbnWxfVAFkOkIPemKL+z0emfAgjtWxyQbTkOyRxNvmSdHR+KJ0dITx46HMO
aA11ECDNX2N9qs5GAeu6rJvIXO+HiWs9NowkZlrivDC8DjC5YpmiD1/nkFKF54rRN59eDV5yAQ99
EEpQFQaIXC7wO5XyqiWMovcuUXuNCor6QJi2n9t5qSrNiQkJBITKaANin3/95Gh9L1deece7q4R7
/b4jHLEzETR6iVggE8rNjiN6BkNgs3ubykF6F39rq1Upeadd5eSVcrNpKG8qKJ2DXya9g42EWF4Q
/gzD4cBTPVEaw8Up9JmQfxOqAKyIQYi7UMiGzj5qQ/ATPySryQh8rVkssT5XzeK+TJ4NN4L3vKm2
Swda7Lkt7t83diS3tOfo6iSiVRLP3H8h/wmlXuMCPZv000tpkoiVpWmmEe09Vn+R2M3dB+P/fCCc
3Syta9pyLyU3uAK0wwrZHzrPOKXeeDbpubXkHNX3JnGfQxPcH/QdU407GVSVuwM4wO4dk/W4Hdsm
MW65MQH8kcDIoKh3rICIvY8IS8BM+58mPPaz9dAhvJ5udm6X0QdufzczYO6jzdXHCTFxU2GEg+m6
/TSuRm65zcnFXQl+qrcDc1OvonOJXzSjcgDC9jf4wsg56SfShnM4Oc3q/cAXebkzDPZkgKS9kWZo
QfISR3s1jll7jq0ordPJc7g7GvozDtW9LLOtW7/b8ZMUAGYr5tsYQqNsEJ8inWYWDCWYNgZ7MbBr
GYPNkahLJqAoyQHkcr8RA+9P2//mHufmCaSB493mtcj0Z+iiy7+To6saP80D7ebsPb+gj3EKTcD4
n1/QQeRlkQ+0QtXvMjKorj6zjw6a9j19gYVJ3/T9DaslZZmyjuUe+96g6fS/DfHKqG0BXu+Pebza
VGEw9evRZtfKZRqWpP/e18SOzN/nylC19Mz1kHFRPkhy8729jYV/Tb5qq0IuhXqrDQ1Yo6LSK+pn
If//2JPlfC0x6B1kpmEOMSZ0LEXna9EDVFN1gV82FshCTTGX/Eptv/4gVQghg7SuSvhT8bqioRre
ID2bq8qZ5O7pvJv9UHzEdH2gkjuvISrWY3mciL4w5PvOnKateSDnKr/199c4en+isMWeVNQyW/+Q
FD798gC1z4pbp2RjSSM+Hl+Tr6iEviEHEwUHCTrvmc+cC//2GgZVlGEZ08oE/cIFCOvzpjNNZ7/l
AgOrz1lIMAUhTsFQaHSF51P4XG4oehFcAf2Wwp01odtMG6UB4yO3KBa693ofRseV5FMCxBmJTggh
t0vGIVtt/Wl4ShpSs3k/Q5+XIuIIeu676q44UnNdq9R7088tfvDQwBUdRD/rUNzv80Uood24NJIJ
HyBuk5zqNAaE7H+HlURBUfjL3la+YFFIiwDlCRWm+s5igjDV0qWPpP88l2k2QaEnu0YiA0rJgHwf
hWbtBC9lP3mgL9EC+o4AkVBonjOWVa0esbR6V0zOmKwoAsx6JHy8MkKV182T+QUaTNEvUN0Afryw
fFgiVTmeYAza4XcQtIX8Ek2FhEOA5Hg51wziwyF6wy+kY8BggL8UXIgNf0fiApYtfwpcSjSriqFE
+43Xnlu1IEwlZqzyVkt/B0U1fqQ7cgl6WnV89l1TznT3TBEpJj8mBSEEQc4Fc/r8iDzvQ6RVMbM6
zm2aLyI979pOUwa67B/kPub1ksWPYE/kNUdIJpQqJIPhti0rQXhdsFHUAp/5q1f4MnpEqTw0MkD8
U89U+rh9xcyP3uLk1J17O4Oqu5woEuKec7iylFwDck/5RqIYiAOxd4+AuBtIUYZy6N7DNjGbgQi+
KcHpAYIcS9u1H5zkbYolB4lJ7//5fctP5z8+t046w6y+yq5Cs68XC3SRad96w3tExYFvJcQ3AaPc
rt8E3wyaw0PX07XDyguIescHCM1f0QX0v4ilYlsJC/4y0goq1JHFmSJb6u2i2koAHMSje2b0Xekf
V8fE9ErmhY7PE+MM/7RqdlaQX0+BidUSmL0d9SI2ZH51Ofg3DnOYgiVMVrqG3ePfqJKFtNANtm3s
F0cvy2ah1uzn2QgwinPFLWtb1BuHgdO5xPCSPLHqKZIULlwo26VJD//iRTjb4C4L4KH9bZOxpFDX
31Zs1uhVLRWcw64i018aq43yorpfn9LJkXe0P8fDEo+WDQL+/xPVV770IRfTXM2knPLZ/QBZ7A3s
BsTZwGKbaFAAY8zxYgGvGS8JuaWCrqIRB4bcqud/zn555nf4aVZNb+hqR8dxYIIzfAgeSbq415C6
vj6TfdnH3icFNAacaswKwD6OEelyLwM4s66FhYEIO29pinmD1GVIOpnvFW635wCoCzUoxwcZzWLQ
3yuIfTArnmNudZp87JQQRuXq/J7SHTOD6vYFFMYJwOdT8qqXqvgRNDNRTqdLM79eUJ34bnQHo6l0
rID6dFz76sorMmg9ujfqYGpPL8MAnmfhReCN/ZYPe0Kps8xB1hloJzj+zajXd4zCTlz5QltHqzLU
BsbnchjVV8db28WGtpZa3pPZiM/yTzSTsfLSvwTOzHg6SsTq2iFhgBXunkxPM6eSeYYJJvenhjQ3
gCn2t5g+VUWQhRJ7kkt2B8PsHo22jwr038nA1ZaKL62Src3mvLXvRx9VYV5HJ5q1pfoVy3mmWgFk
DazYbC+/g81p9ah2Y/WE3t1ULN3QKaWC69AQwNGcbGNkzNDeGHLj9alW1460sZFl0uA3owgiBTJW
NzENqo/MGQgbk21D6uf7Np5IqF9MG0T1nT1b5o+2M8/LYUTN1QKk8dlBWRQu+WKlXbUt3EWxvZ+e
sMGOtm++hysjcglezz4EPWJbIOxZSOK81Wzv1XwC/VB8aUgfGR3ZnzS3dQ5TZQj7tdcHfydewnwv
8U9UtGY3gfjjLZsnZ+OpPr6/hHPbtrWMz1diLJX6O+Am1P2LvaQJPcfTRDJ742lQ+K7jmjq7+0Lo
iaNvJkBbvdVXvTOFicaRR+h9YWnEziGUZyyMSHaSI+4kAQWWmL8kN63bsp2bP7IRV+0Ccrpd2AUs
JGrg4mImMCJNcZKPqi87xlkrn6ywLOlXO4/uuIh/V3hgQ2O7R4E8AfrzjNDEG+3R34iFWUXpJyDi
LxMV5My/h4lsx1qfzjhBzBxeTD8MOiTKpcBCYKlEIy7+Wip00pmwUuw5Ob1NF+fR9vF+hrUlvshr
fgXlu0FZuDlYBOWVuISGtWAPnlfQ60zLc9cF9tIdcY+i+bKAqHu9pWSrICmmWEs9vBhWYzIR+Yx8
f2/QOTE60tJOLh0TLDDKKeZBRTf3tMZ9mfuL+bmscnYcTdFHAFtwoF13kicssk7WSykfkUlrKq75
mzqwKQJiSqH3xGUYTHI4jO8zWwniO22OXYfc6+tao+n6LZQzGdSNQfFXkYJmS/qOdimjkVNMLxip
ptAr2OSpNOIiQB44BuDCLx6Okyh21aGLB1naUQuugtI3ZaQNBsISSG+cQom9sOvsrYkrdT3rrI8r
Rv4SC2T1lWElDyCXjAZeHuYeTvApsJLgIbmkrBg7CmPiHR7+rkuUlhO/7arIHZ6vm45xRlk1YPYh
vgA7ltC9VMUPPjwdwEKMbZHFwT98o3FGqrUQeyWxVf21UeMv913cdYPhE1PdemvMVb01D9UeTSI2
2mLXiNYTtbBg6O1TqsNYIeXOxfrBzKMa6LuvxMAmGUvBmAQaXPLhegtrN74odyCsRBZGVSJKmyHc
Jlg2YWcTVjaKIAwGaMfVKjVAzjWkBUrME+LZNIydJ6wF9gP/2vRVGHJ5msNXcuTdGj++y9dhLX4g
hCrgMhzpip6fVxfvQ1KIXGm92OfeFOFMatfgP80WCudAE0PixJJLOmz07Ti3JTfR3ndC22eSFGiT
bxm36HwF6N0upbZq+4v+hpBs1hcAT9iclfb+7q6FDZPdwWUy7YvbHnOWnEQoCopaX/hziU2kcoW2
atFskgAZbbwUQ46SGpxyyzgfcQInAIu6UMaQvK7HKRHMj2Lie0fXZW6uZNe93S7/jlefEPUmCMum
ptTDgcspRDGc2LJbt4b6Mr+XWFgDffBQqlDhSHJ8P56xtA7RaSN1Pqo5DvJhOtc4UKivJL2fLIxa
YAnOWvVoGlVUKwFT380CiC11UaFY/D+wwbRKPzWjhkM6VJpZKiaUhuZocHBzIIwShdxRAfNjhr4R
EPxzIqncNeK1YfJ6KNA71DTOnhs3RVtgUAGzN94dwaDLcsXy1ygFESX7LCe31jCCBVjnJE20d49g
1w/nUnOnQtJuj/tXpSvGPPGwKdKiROnu+L5VbbXR/XF+DP8HQ6V0pTG5F+YvVwZa7b9PrAytxRbl
J/tDEOBGCugF1thEUODFcf7D9ra3jwuEjEaKtsiZ80EbBeO6HacPeT7kryk9zas1jQOclHARgIkK
0RKo0WDvl2iU4zTFqJ8BTHGvNeQkk4J4HV6VN5Mk/yyHAmuF4wU1qBuaHxFlAuEiXC8ptiThMb9O
nWXmnbbtWNb2q/YiHHFt68EDZauj1Ph7mo7ACPgK9wDtIJGSElOILJtdUVbSQdAi2YSFHAhj/mJC
icg7QiAge+tzPWFqIhVusuBDXBGx+63JcAuSqW+wifO8l2tyuXp53Vtq/1Exo0blNBPnAoQ51m9R
ECvVT2WAJFrdMGfI4pjgJrzpawIyC/BM+hSui5fpXbo5xjOi0/ua2wL02UhTWWHtTbbl30/xAR8S
6Uwn1FZSiIjm6Sn1/tXsy0CLrmd7DYUy1QRXpI8D8H75EgVBDYh0wCejbJuPiwbz0dPbSzOPCM29
EfyrftMZLZOUQEs0B6aRyPdy2k+7je2xkhtd0OLrqLXGH35APyDoGE2UAZ5m8QY8DTyHhaKQRscS
lotCLq5y/d4uLhj2f9u2RpQJdedhoKSwz67z7yawb953YuBqiUAB0dTkO0tdKwPKD9dydWqhPqCX
SKwMyTkgHTOB5aQ7Hn3tiQrnc/z36C7CrGB8D1YPYQrBU382YiWe1hT5HLxgD2hPVliZ8DiVEDbo
0psVh3t60yxwqWhKOElwk4cfY9gMC07XC+UYOJOkh0L6cPEeu37MpbjUj35RMQLUgq5IafeaPdrv
XvFurVFAMNTG2yuVpvkVAiYbAcjk3P+SE521ScZlzbOFMtERPPCL8HFhObo0YPFu4rbjyZkh4hE4
rv56pFMtlRRJsVO8sHGCf48bF0er+cwmqtg605jxfpdfpsdpxAt0qZGkJ8b0XenRmbP1ze3/GZ49
jY1cCogaDWGTMM4l8PIbaCJH8s1hSWLYfzwnzwwM1mKR6x7NpaYFVTuBZVp4VuZm20puNVOvWxst
MKnzC4B33lg1UUPbZKyBFtFNHuqFFjkdxbDmaPVC3VCk/DIgQXfcPNYstxw6a0lz+wF1OTJX0K05
LEv4bseWyeQz7Y7gTWdtQ57JZJErshyKYVZQL/MCmx0R+aFVHrV6LMUso8aydkZ0tnaBDJTfvjXd
fYwlRt+wHaMnPWOOQiRROfWhzlefHvRdBcyUzazyUKiKlElqioOPJlcmuC7aVL3RJ94TeEjBHZCe
zRX7mSYA9VnMv2JHi+/p8i0QStYOan+C/AUcND48bxkz43+pkCL8lViWyR8Vq2snet4dADpSHv/m
l+Kovl/oD94LCxUAwr/IYgU/g2I/TXV3Zp8JAFUse0cZ/fyDHl/XmSZq9lNvsG2qeJPoZ1iresD1
snxOPGPeNfxhsOmhWWRpU778j1WfeOBjjloFM/zucBBzjVjQIJzq5LsKVKHDuCiaHM5PpLl0zX3L
rddBdkwo27Dj2S+o2spWFogJ+eDHeQm+RwE7kfKX2Imw185b+Gtvz0ZWULpOc8Gz073qIcRApwik
NFV1j49WhmcBu9aXINTWnWYXTqktzZ9J4mY1ElwC7wO3eqq5U8Cfli/3aFmKlUbxu2G7YTAcV+JV
8XIpLGoZRdBv2KgyH2Pw5+xYk4GAlPN2X8K2hBkBAqfHAHJrY18JZjcY7fUlNrTb8ZPihgPPo5lw
vAsacPiWSrCSyJMRixjcnUoLYp7NsWE1teO36xDEwiIscRIK2VxGi42RgXj0nziQn3mhDCD3sv2X
3TxWyg5g5xT7FqRovVQaFnzPWzbm46stXLXitDWlgxNzLBAHdsdyvd44/5z443LrdLl5GTDiIILT
PKjX/ZBwRL3B6/EwxUtYuOiu4+f+u8GTtfyG/Hhm+HwMLYLF2o0ngRt5nrdpWAy+B5sP3TkK4wmt
zZGwrjiT4LsaKzUr4AqFhfdd1ZcwHHOWFbj99SyAFlvI+TAhHFwLW1Y4b1qGP8emZyxLC0y6Xar1
0yjrzWIfqtjKi0jr+HdSxiLbFVoLfZqZEqdykHObvoavQlPNNPPUAvXaJNFQbCJykFZphH1BdfRG
5gPzbmXhlY/Vj+p81c83qCRCTvcHY5ARedoKlx1/xPpdmkcH+Z8wey+DUaLmppm5lPrJj+hJReJr
9Ss5AaacWkyOTZ9ekJHyBoFbBJwzxmaaZxtLSKMlK9xhiCAJn1ELQaHIuuo8C5lAaXmLA5o6MAAz
utZdAe3SBCA+7TN6EPT3wVwAg9LcjkScU4ce/6sniJndxEoruOV1eLkj6Vh4VkBGemggOmdg0Ewg
jCnuVnNNQ7SHzKr9B3OSYhKFkyVdoR6OAwSzZ1LMh07m0PeLTmEalebNzrMyVYcAnX4ZGSnNm7Jm
84C7mDJ4oJr6DwWNU83oOy7etEBUQaIU4uueu2K2ePp07Fil8IbogQFuFpJato5oRlsAN5mamIUs
quubHdqiBSipddtFpyTN8vnmKAKyiemtHw+L7gSLCoHs38ovG85ZHREBhqFafFycppTMMhHZX4rp
ZGxC62lMR6+2av2EzG5nsVv60eaXNw2ug36UAZYzOBi4RqImwRc+bE/HM9ecJATS5IwVzKC54iIl
CkuEskIswll73OACdVXHseIRFapS/eKc12J+bKrMUxEHypvgNEtSGb+/DVJAVUcdquvtBDPDnT3G
rph5q2qaqjyzlh5W2saPE5pQ2iDqi54AuAAf+UpRt0jxiDUU/y2c1J2Sy3iet7ZqVO0uk+GfQBH1
wPq02SnQN9pbBQ+66MONslmK5b/cpRWcKcm0FiaC2Jm+ZF33eELSI+QL8SFJQFcwjIXIBN59E8VA
3XFo8t4DBfGWgQQAanxvZtEkzC0+4LURqp/Xe6HfRyqdrBI/wLLBMNmQ02Z8MQSPTi+xiJgSFQ3E
pLUW7xFkXUAGBH5pnAkK8OwuvbxVqdI0q+6PQFpRYZFV+KEV6iOlinmybjc0yKJ/1m+hxpdprqQC
EUba6HRmBrU/NHWKUGGO1k7kSxuRaoob6BjRjTauheRuA3TYsnWnbFK7Sw45vHieMaTHbYQXYPBB
P+/j3JjRGjfQ9KWTcmLtIPSYa0qpmLiL6P/latTMnTs52ZtjDL+Y4OBfp/rGJcxwm4fiKBVFb4Kh
cgYdKUdMy2Cx3s9VRruqgcyQmLA5Hn01o5xdvi6m2OdQwRv+WVzPev9LLnpW2Cf5qNwLQSlEqi7Z
sBx5tZtn4zOZadUxH/YdRMJn/s0qJIRBJ1zYkU/mWK5mfkfy6PG0ID7WOHy6Hqdeb27ZDTgejac9
BbRPX5VuV4aKrGkOWgBYMSbAp9vYmBUO77T+8WwY16dPnx4HaJb5CHnEoWBOgltJPymS2ha+UNWE
oJsYLxO5ad4XZtWW87mcW4nxHynIumd5+ij75QWkvaAu4TUoQLoXgdfa/6v3ttIZrOUeMl0byakO
+eOBmGy5iGbG7qfzwf1DhIHT3y2N64gr6O4Lr8Qh/GrlgVI01WEtFjCoy9Ko1R6YJ64NfKuIZbDV
pKQulW6Z3CIl+gBpI0yKfZXkowfSRNM/nnJTkRMcA6i34ZznJwV35rxd0hm4e0rkh9fUpOpi1Mv2
MQgZJAjwo98u2wTLkQxoJ7qcpskYpg+IFSN8SuBc1Pn1b3vRNzGm7CELXti39j1rtg+Agccr7dGb
ziy2uCvcIfZD/Gt6weq0jd83a4rYb3sQWCM67mDfkCZwkqjYq1H1VQi6H5hglWTACCs0igzT+iuH
IQF+UGFSd+2pjS7RIQ/ixTLonfqZQLgC6a82BIXnCMD13+ubu2eEqKZlWosUqdUoadYjkGuVKnIi
DtmyamxvLtl5lmLsZYx9Bb9X14brHbR0byhaVY8lPYsjfeV8zmUlrXLh8uo838xuaQA7NmcMCwS6
Lamu5xnUgAQjr2LnjflxtWmL7rOHTfzLnOpWHAgmqJooJoI3R1uO1L61z37X3ZaZ1/bbSy6BNBPT
zpL3Pbr+ka+xPTJZZnTX6Ybdu3aKNFtiTvI+Xst3rCVUqvXsZLV2ZloCTW94GO8GgNMib/CUNP3w
BF27NIfr1Ilqq+jzPNZ8hIK4ovbz2GQGS+5CIJ7Wj1kVTq49Age33ItXUcPReg+iLiybLoUJvxFA
YkI3IimUIYPd9RsKnVdYIiyiT6GaJoICu+9yrrZpHsA6Er4cmu/b0AH9kM4LTVdxdyM8y9qMkXrW
eUHJxXX3+hXd5HLekFiXQNmt0wQ45WNiRK5m70knbB994l7OmwciAMgJfwf01zyjzorrBIO4uUFM
qdcMzWUygrVclatIQrzszrIRDlV8PUqDn587GHK5tG97i5NzUbCjac4DK5eWpOgbMSprgEaL8v/j
N61ySq6znmQ0oM1gel2mZfl+7Bxyh/2Pk5+vNZceybV1mqrdBH16QU74Fwco1njFTNxXws1QZu6K
ZDQMXylTB9ydhHLetvibYEWHjzq9utkptuTrXPBwfe08svBa3OP2xyhMtz1IfPrOlfW/gmfTLgI1
DAcse4BckWccDzPVlRKQaNgq6y8hBt/T73QvC3fep6UooeskiREfLJW8MZvZY0CC6IXXaqCKxPEW
HDAQgVXL3ilVs5AIuwjLaPe52DjyiAsOrk5wPGLlf24U54oXLYDvNhrs68LIKx3AnBJUw1CyyJfi
Y2fnXGz5xTG4ThsRQ1sQT5vNJvEMXncUfNqMBcjMTkPNk2xNNDIFof7o58KfzQXMx3Dvm9Pyr52q
xkRFciCI9G9cm64fSmx/dsaimAOzuF2rdDUGOByW9Rl8EaxSlJQQSQmo+HnH/8GEdmU4LjewfK9k
1k6fdBVfrFQPCk/nFoyVZL+03TGwhlai7Rv6ry11Mi9hm1xUjHWL36ofN4ZET/ZGQQhdeaP5TfIj
c/6gqEYZntQif2hgf2my0XQHjTEciW4tRBBpV+tzuYg80mre6d6skkbd4dUMsMOL19k7WdJse8kS
zMu6looQZo0ERg7+FyCNdVa0hipx3UpiXNNBaaVxhM81Le2Er2dg/8YSMtPX2U5XvwAsalyoZ27a
ZPv1Dr9c4x4pzZrKP4ld/vXyfy+muti3PrjT+Kxk4WsDio0WAoPkiNJ/6Lri70sNO9hmvSQQy0/T
bl89jJjR/vMKO9J/Kvw7S+ehrxhaQ5l4EThxVGjJdnet8WZgseNqEPuRuG0zDeIrdQAReGR2tppd
v/GkeTP98nJlPdGoND7gipSJW52dprUtebnlWdcaayautlFtLnjmYqcEnLC7BMYQX1C/SDJTeY26
OIJHuYP84fWgQ6jivKod+nlOO/rZ0tHCYF/gSx7ex/xJcEOQp42+503iwe7iAs+4ukpRX4O938DL
Z/sMWdrgbJWOqfgKtcCYBDw3xeCi6pxFwXi7o1iMpGkyvVRWw85jbIoJM5QxkdttzGT+/dhcnHOO
Qt71I4fS0lcx2T1VqxbKblj2i0tK1H1OR4rRzCIsbnPAxZ5vzVh/Q9Md1bFdiXtPUJsLOS/TBtVy
N6sgzSXyt8M0ngPMDK4tWL1agazGQs32n2os9v9SXx+W8N3f9urkbIzGu/QWVW24qg/NkexC/xmd
5TSXA/gupsfiev02D8RJcpHgGV2q22no5+GNJWah4/Lnx403mqqqATGJv4ZhXJXcBSOuekrGDUyZ
Yrc9G2BGDq8ZO2HJoDKvCNLmpI0qR7x4GX3aDZxdmr0HTxnEjIQScw/QCmIyJSjEC3Jc0gbIzUGu
na4Cdv2mTGb0vzJYcB5CbG6I+NASnLmEAhCtWiKXmQeswam2fVmNiL8LnrFQ1Wnwnhdc3IhRizvQ
CHoyiU8vpsJyrQP+eVyIC6O/1ljf3EUVhZs2CSca0crV6qouhGoobX5rH0MjKneigLLVOFeABPOA
5nJhAbxaET2VSKHzPugK1jzqVhzuSSZNAIejxuel+lpqecNn1VDLxc9ZmUXFhPHGFCk335bXwqRq
ryYuUA244kgzCSDFU/88zfaHdpeRWvOuYQs8Om6WrESr6x05GE+N+Y+SiZTI3QLY6ZKPwXjg7cdo
XTMOjJvWpOEtvG0DwfmGubdNfTgGkIJDYlcI+0SYauQS2mpsOZtysj0YQ/wenx1oeusIL6k3/dSs
g/gzjRUGFyvPNzxR/E5uZPOfsMVTUm/TZTzXHK4PX503GdnlBCTuWXnT1fuJyia5DY/QNp9FG9II
OJAY4+WGlCpD08/73ZBt4N5W9ys8zVxz5CJiDrD2HkpIrmrRTYCSjgAfjE7EvlCDYkg/aF4IR2Ez
lQu/eJ1fZkKzCFODDyp3eJt3Q/NiNQPnqkG6QAIIBuIZ7QafDG9tBw8hru/ui4x1OaFtHQZwpd06
kU/oVNLJVVW5OjWugw28g0ImPA7aBvlCS98Gw3uF6YBR/SMiB6LUlDyQEq9XpxettKpy2WQ6ZdOf
z9GbpB4Rn2sh8v5TkWyHK9mbzrKTDcQ2TDSV5TMrKuUTMxO81tA8KfhHtcA2t2yTJv1HSm+Cccee
aiyHg2QU47oamuHRv3njaF9QSc2fG4zBHYaHWaXZADOX862iO0rc/xktkt2aGyKdoQWODW6kBBwh
dQghnHAEDQ28RUmn3b0VJzUvUg5LdV9Ec8se/3Ffk+3YQIuTGpgijWnAHYR1V+2rpsOiZDMPMFrH
Mu5ortRkbYSip5nKFglknbUUT/XaOya2qWe4ip/2hV9GoOItDUTD9CwFHPERYA7OvUJUnSc6uTx1
FkO7PpSfukalVpds98ysV0R6TutKvZSlLGQh7uULybOSLukdrnWjfivgvm/6vXd5tzVcyG7ADgHl
am8VvXeXgQU7Yoh2k59wDgyU6j2fJ/Srxv+wke06CFoGPLedKgRYD39MoOLnlqD/zBN1Ud34qu/v
FHzTaLkm2Lk82W6FKBL3QRYy5v8yrO8l1eAzhElWxZaW0UdaCAkxMH5B1IMr5TnYzigG4bsUzVkE
PH3Zb5YiICzp70J5IjfsxIsfdO/KYSNL6vNBxEir4cT44xUU2//uf+G2bkC1ANhi0WGU3/wWEMDf
bBGDdTRnLL5jMRn3s0d/boqBKvI0u8pHYhPuhpaIiUmYafoMHsy1UqO+iTfk+vtJnps1k9jyCxP+
6IffpQxQWrNTbHDSOfoM0N/UZ0gWX7wyNT9K2u2uw1vdMhlW2ehUhLNSxMGEjDOgm6C2F6mLAfZC
KAjXDxhQfzugcw6FPEVps1vlVa9rqs9/N1qmEZk99UXLOtedbEWy4GqkK6e6lTj7QOsHvW9eymdP
63viFpHH/3y2d54jzfmaHA0OXCHKW6snxtazJ6ru6A3SraCQDDj9U5RrsxQYuI/pqxA5CkqGY4dz
7xR2a6jRJNbrtbW1Gi5idkAw9rhcOVw9IOu1QnTU5J2ulHw6v1/KhZ9+VZvN9je4yuWrjdbJ3opM
1v4omp+Y8aH65fA2l4KRiV9siM7gUy0sPUqLTgcRQNxKpUJs5iEbILBa/TOF1bTXv0qnhz/RWp/p
cwyxnzvbpmwkh42ehgbiksEfXGJ2J/tphmrRaioKh9WCQne4NrZ2jsdwbEmigiyQ18vglM6oXHcq
afY8KcBDKFrs5acXaltZLW8bHd1gfmwTs+sMWBglXufo/xTEjycZ6fseaBQ1qwQI2+1K0ldUmczY
wGOp+TD1FlwhNdMQgxxYTuR5vS11I2ytpCCDyO0X6rvK4UjNq5N1zbADukLuih8SfkvQuhaTGXtn
+tf9ARTolrevkgb2dh/c8PIpJlEucN1gz36zNYxuhJ5V2msmhN7rfqOiVyPxt4xJrGKZBdUNYvyA
M73V00qWEAMZ+W8fADUpl+FMC9cCHtyzZuKXZnj/Jo3fa1Q2m2sRz0EaW1dpBZ9XcutqH1W1BbzC
iBjrIYpT/4rvQHObPRz1IThNq3XDoNKG5V2NfEyHpqRuNsm07taPAuArYK2vV2M9iytCro+5BN7V
n3eJia+G04KpH8j5sy5OuU0GazQrVssj+0v3b/XQMid1bBwtk/+R7bSZZcvAq39mjk2WwvNmJ7wB
VMhWHP+Rtu9u69edl4dGkyau3Gbqa7z8RPchrGn7ctOUI+OWAv66IfkY1Cs+CvimPoPE8ZHB5zxs
saIEFHXR4zHcEU2V2A5Gt92fzYmO2pUVIbNCkNusRTBBbo3kOZeh/pHl0O5VMxh0DpSAXE9WTXaw
RlK6ktHzi7N3ntw1mkyXdQBSdeN1EcL8+xewaQCD1iAMBzbyuAsG9nZ7kNd/uCDQXHTAp33IMxZz
qUDR9RgQV7n8hsUu1a/3zLS9cjoynYsMVtcSzal+CE5fJe2Q9KWri4qes5hcjRcSUbIpx244HG3D
fYygUwOTCCSsYwA/zz+sIPGI/Pd4ikheiMuW9ivfWCj08dr+ivoT2Q9XS8hHnuGYMYpK1W8hUPAE
D6jA9jDpZ4aByMdz45OrwV5dT8JaXj2yyYwBsXtoqSlXLK9dfG3G8qESEIEnhnw/JJrfYDfQ6C5n
3sOgIS000sOxS7+22rgwPxIB7APz5ZSF28U5HA/vNAEcqvfHOOQrafQCUsoAHFv7GAzfXFFyWrGM
VIa8LfnznTCoG2EKtgzy7Kz5N6rVGDPx7Gglt+GcNmiZUoQG4UIBdE749+w3VwGrJRcJRNfNceUE
vS2j8R9WeoeYQi07twOAf9zshaRcmF/tq/m/bI4jAivKHlXSgsAyHffaJHL1RwVlYB68M51ciQCn
CqpvDw3/UTYhDkIPLrkg3u4bnupJ714wl2HllgVkcJy+n5//i6Aw/iRYXyjyDiJYtlpPvSL9UbMI
frNS60aJsfLxbM3PtmGmnD5Dtsw4lRpfNwul1SFd0x7IaNxctebXped05gFNQArsfAOEJg/MJAGu
1atth7cApE4tSKIaML7Ie6WpniKDsKBGBjRVoN+llrOTel5eQF+S2yfRU2EBuIn4pBxpMPBEWDDq
MTPIrkYrrpIVapyepOoNIlWoJqZF6gyPpA16yvM9v04xMr5przx8qTy2a3TD6TTtCoixKgCQ1NE+
cX9DAMk0wOeV2lihf8x8nFsyjjGKXURCztfnD6xP2ExoJPdO2KzvNSBS81aPOJFb25gIlTbYFkY6
19RTlLTDvQM70PYkXkEAJMPDYRp0H4p8sAvc61GYU4aDQ8tcPw6iHD8BZu+YNwVXddU1d5RK/pUx
IwhaOlgG9+db0hCFvn7+SiaSzfuDR8Fq4v6/VSO7H7aDUiVqMGgv8r9YmNXeydEq6QnL+wwsOBvI
S/YpCWRp1rCUggbKgEa99h0C7R3QD4BQJ0yxM3NZSdHIuKvqL0IF+3sAaabk/mH2Yolyyy+IQNkk
iv68TRAiRaxUPYmIIIhKzXxx+mL+AQBO7rXXghBOBsk2SVWkklPLU9HPBbOShtif6UaQywtrCke7
yYv4X3Dr+csR4wao32M0Ow2qjMmDPEX3PwV2zpLwm3Y5Tg8GGb7CA45W/LbRxyHR/JMQ/XION6hS
lXv5qRm6FA4oc7GcEDD2CzjYviW1pl9XNj0ocWnJQMIiEFT/d+He00Rkorp+zGWAFmAR7Xvsc77f
04Mi0l9ewk7LI2mwPB49sU6jiyVqbfu5q0amjNlAW0arT3qlWn33CNHEt4pzu2lD83k3KCT+Pduk
tiTe565Sp+ktjSWEabPtOurOkkwA2bPbb/ng1tck6mT8NmP7ceef1kEBH82Igq1NXFGGsxqs8Eim
Hgn/2h/59G7qJKRPeAOL7/thkog4s6xmktm658gaQ5lHfmSy3hUGZqojGEv2wyq1uRbYYcouQ4af
L3Kr4QQ6Z0xCBTyLlBrNONv5as30oD4QOsFMULOde+e5of2j0trGO2mfqODjbaS5A84Wvhken5qb
OgC7jx2Qdwg/HVZPE4i4EyH/VP7yWDD9L5IO8h/uJy9pNzsG7StOkl2h/IAWaooZGGMRyvQZ98Rg
09jjcX8gF6ZJsTjZ04l/RhXk/vq/yfmLv/+FeUCjNwSiURkUQtM7zWERsDoqCF2GoIRH7TYqQU7z
ojAqWjBgMXlqHT/e7LKcuFkAq/oDUQyMoUGM0d4Eo0LxY8Ny5Xb5cpOt9C0nu9WuB1OY4gFEPkt+
cBLSHvJXf3tfyi9vKyg/oKS3VqBFph+72F7ppR1LyDDCfwlbEvdUrzSYeph8YwdMYHDzXLQQ/daU
vEzXJ90Jj3GohCpY71RHtkddoOkVE99RMP4bQl0+3yMIt7g8fN9UIDq0GWKehIzcPhyXN/7zxwFk
mOmx3yDfwS4DLGOZYbq6tywCwGwxrWG9mlirM2yzT8kdsvGlmt5IKr28LpHa1tl7OrZ53mdDStJz
f/MJr5OvkS06K5ELmMfmEziP/ySjTLjvHr9ynfDfiV9eog9q/+SCZryBPIZOomJ+3ONDcnNUXaYJ
jSAs+9DUvoh9s2JGgf3E13Yp77BEhpqXpS8i4lKD2aDOrYN6MPBuWN67zgp6UDORBPNMcBIMTxLh
my9qDHCFX7J7Nh+y1NVufijkO7YR4MO3PMrErC8VZN830B/XogT8xppf8qb+3zoF+DIfAkjyH4+B
tkTBCcP4oWXr5Zgtl2RiugOzrjioBUhHk2I4VGjwpIcvAnGQ7gf7hY4Tx6kGIA+0EY3TQWu4Es00
Tin0/agAkNZVdVmRmsM6VNXEAHvyZdakIW4PucX9bIu9RjIfFEJhjk9kJiBE7BNxusm17XGG1xNu
2P5lAEhrZKFtTy2xsieMJPdly6GSLSLhlkGSBegp8CO+CCv4T+dtsIEwfMpESAEY6TTnMBbMHHCw
Ph0INyb/8TgYD2SdefYebVNfzACTtgGaG32Tzd53fFlZfr5zeGV98eN9MFXTg88V/NlBbgqVlcRM
jOnSb0/mCzraBvdyhKu/T6NODW5TquP/DAc7/IInxiMaq925HRrNsYZCg0J4EgoqyX8FDKNmDz9x
aVNjM4gbzjZuEpz2lKUXmakvVdOUdpEBaistnSu+TpoESh5JXSErbILDTTNi6HRz+CI/LuCjkkOO
NnpnKrXJKuUTC0FcwcS5aEIqChjazA+d4WK7Aokwy25AdldQUl+vTpm3bvrSh6eaPq6WjT/ALtGO
QOWrUazPrSuq2M2gzdZetKyo1GqmLdvkk/ni9g4X8yJX2UkS4uc0kMfhCer9QtTjm02o/PHC+uLo
YLREiggQGoUuNPXsF8hBrumXf2XkxFMf3rqS+Sk4uSL93yJvBrjoIjluDv7CWrc77PfdwrO4263Q
FOP9Rooz9Os/MV2N+87XlYOhsWN6NUUSSJE210tQ5h0IPyxSjfGo+4OfsmsUllK1eEqabFK8vqu0
ARxtgNebHoIoVWwZObJGjDANcz9sDC9/Fdx5ta/99yptEvQG0ZxQR23+Aw45HhDS3QfR6bQ+UHQv
Jq3IGjJXtfgt4hfTE+ekKyRNXDyhdd+0bOQiisx/H1DCOHuUfynq6PMP95GLqb5cfvZ2yUzhrgQ1
LuBP3xQfMhE41I6OCouGvG0GVubNXvAd8sc31mHMWCjrNKHjKi0yzaSxfFCO5bvuy06JmlJ/WQHg
1jHAP1bEusMTNmRvzlrWPV/jeL9ARvO+lip3p/w7peFnls+z8a/1tZ/IM+SF9gFydZKb6QUIciXv
Vcz86oZMQSePEuRhc/Olhb1AP3cBNmvXfXBFFPRrc4eeRYz5vZVse/XbZsR80LWV6HeZ5Z6X0qmT
Jq2TgBIErblYCIuxFnjgoX1aWkreOJcbRHq9mjzdXb4he30LcgLZ/t1eNxIBqLWceA7vjYSc4quk
uP8RRFF9Zpkg4UQTs8XDd6nPfFzDbttHNY960YUOuD4PRu7AX4JPQdPDF7edJD1uQYCGPxuv5LxK
QAhOGVuqarIBmKbwzYCizs6VxtPQjYlxjmQ1VVv6veZ1eCTg0PWADpsyTnh51rGsXqBAqDxVxVlt
YI3/D66fmg4rSVUig6Sh5TadGznfY17RG8Frh+P0VFDsAY0VnqOJyho5psillxhMtXBc4cP1HnCx
AHNcAr5DY+LfIfpQ8IbNzN2K3Q7az0jE+T3S0m/InmYeYGvu7wZWCEITQPHm3pvynDX0OUgHKY2Q
3RHum/RCzLLyUpbiJutjnDIinVDoIgCm5qBzlQkrw3n4QGUdvHYAXSOiC+ieiF1pNYBuywNw+fT4
xG0IJZnivONDFALLuTlZSoCZnAeqznSMephbwJXYSi16Zr/1lOnVxLMk/Q8sFjaDLBLtWwccyv84
9vfRv0VZ7K/D2VwyARguEy0Efea41ArxC+5wc+gE8oNyKIno5UlJRrTAtx7dTc6ByoHtGpywfU2P
1IOmJNpJoHmO2j0p8baQEW/+LTcIjy6+CplUuM6JTrdbC3lEb43EOY9YO9Z/t+uzmdBeX3FyVW7c
iUxeZF2/CM8t32zG/NgjMk9GsXysxqd259LDp1tuE9o1kfEE4dqodun5sYOaWPpoVyNebwZIx3d6
gOTF67EX6gIhA++iod8Fpg89aYNvmSvwNvIbVb7UYF5LGEaCpUIU7OIk7ZzzRkTiBefTz38AWba5
2Vw/sInLWQI0FxrBFCPSBIpylfl74tmS9RkGB/cIUSu2jjYCVCxcQgcx7eXHisOhCLZEgiUxTfG7
I5GPJtNp7DtPOB3ePZmKdoTRgdMZ740kQLzVWN3P0MO9eFup8FEw4lFWC4vo6dp4Z0eZrOyF422N
nikMyPy3di1WczoN41vsokCh/6G1aIlzmYgZODtgF6Eo3gwhJzJb6An9/x/KYgpgPQ3kkPPf/Vc2
SSkgutvZDnvLj3BZ254LkIoYhtyZHUnN3P4yDAqRtXRhSnxw6irL08GDjNhAhuInYxPoMqVwdLTr
NhEBlOfDuZNyHLOglISw7WKFQiNA0v1NU9eLfxUGO6ZfMPBu3P0oZ9/osn6IrzB2Qb/++PNoW/xT
2VbF8i1CFDMBFsw6FUmeEcuMh8xNJ2V39DUyn9CLLMhCYUnVCGreEuoMZD4kjr4WSq2EkIEh5HfE
99lHkmcm/F5PyIKCXvQfs/2A+SZyP/o5IffQGVXGRzM++cyujK/Pd/CmxbevYPFZQIqy5vi7zpms
MqsVsZqeQPIaygSelu6PpfGaXdxmLXP4cqmSqhER/ek/Q9ci4xLzaUhfkKsfwOGVCm3K+gxoukhu
NF7jdaGngufjTnIpTUilXKUMTGPxXKAuJ9+7Dk4RRzxlv9n8haxWY9DYFeSfOOicyhs+ginJxHuO
E4X8rRwo/BmAjBUMc0B9bZ7ZXcjwcJsIeDARAjjg1TDsHDxpw/NZXOCLWYRy/OlCHIo3n2N5zaEW
GxWl+8uR+4gbcFh9vHXYFaofQ/ZjCRylbyIqaIEzTbW3fRTAkabdq1W1+WW/d+nPuonryiVSNPWv
YQrvXada4RU1cP3iYxxkWdM87w9D+HAzJRTeqnM/DJIsuN6EGSbuaimBmSUAE/sa6OhmCDZ4hyEK
3ythEXtNsfcn/foubPOPudmLhS9hwPhidc7ruvHpEpwAbvOJiUVLeIVPFA+kLaYbbId7ozyJ3mR3
bdCh0AbXKd7WJayGz0El9qM6rhL3m8ALWT8vmgKBk/r5iXaAx7amlKYMDfGGdoaRr22RiVKIVGGr
gzf2saRjcd3erfobab+ObmfB1MCxZPAkKCdoj1SUX+6IGQtI72H7tAJIEmykdyvmAG9Z/aRzKTVa
rID83nDKdPsN0Trs4oLjNkZSCBCsD7IbmY+lHWJnFSoY1RP6rdRhBv+8h1JiGb3RQaw45zDV5AFh
H3DDm841QddssWNzUL7kI6wBKsMF+sR+WKyxqTaC1FIa4zjtYqCZwdEw1FsvZR3zOPDzhFZv9EnU
P8OI0Fr65tj9pped6iYGA+u9bVEMUZ94N75XMFacIWHL0Rt82//pzAvRPCGu4rRAeS+9Rd9/6YPB
IwKIge9qO9Zlqq7qyhNgYQpj/40l7Wr5Jxe2BP0q0LVByOBqw3pbIRRGXyQVJbTdzcH+qOMfgtSj
bqK/mSh6gGvHN1skCfWnp8T/qRBre+mT0oXCA36ghd6MyA0qpBTcTmYhoscVGqlU469YKxdjXuG5
LbvFF8PUvuh6eSW82ssEFFXXOVqarNwmDvTWRYa/W0I4QRILBDiLESPPoL2AHASI+BVG29K7wq/7
sqmVEzGlTrbduSBSGotrKkgQbW8serNcW1T9/pWHWTNfdf0e3QVC+zcGkUgRokyafwifXmpvU/dG
l/epV/n/FezPqM+9r7ZhVkz1WAfAUTTdzL/uCVdUQZzTSuPSnsF3TiUNEWYiqyaM0NQhrvfibZhG
QbY6tkJdjJYbadpWfCMGNODO5omtqPUg6y5H7g+R0l1RrrjcrpHXVlQeaAdvk/3EPt6z3gLlgLQa
q8rOWYQXclw+MiCM8NjZpymZWA60w82Ugx+7ElZNnjBKqsLFKPzEEVvDHOQ6lr9Rbkfc+2GwZP5G
VVD5HP3+aAvNEvr+/zNKVuGvXE0C5LV6C/EfmW8IipN/UAX7wT7F8dHDALAd9vbr8/GB883/ils4
HoVpnam9oqqzetFAI352NDcpUM0JB35YsGFsOJQz4p+J8rB4RPaCHhoPElLM/I0EpERw0ZCz/kn7
l0Tpn5Kdd4aZbdQTp40JJqhrfqtd73A5iAENu0XEJihwbYuUnlk4j1llHWLeoqxnrVNi6IugDeQZ
sWefyp3DXCdTbLc0CqqXFHaGYO3yzF5tCkYsRVDKpohfSRZQjl3uxKBaAxKJUgI9EG+7/4rAeYsp
tN/cL5W1UhbEgmEUXlPVLx6e4M1MutIQjndoy7RhDa2QxvXsvQn2gVs8VReaDbNdPMjAS1EvSqHM
Sy8u50RHJc+8U7kyfZmrAbEGnBu8oGwsXudlvhqEkKESE2in9Wt0AyKF9P5TDaxFqFjzJZK8vQz0
y4LUE4EwZaWl2NdVIIBjL+DacrL6vh1fk+4HAys84KGyqZ0k35crJG3gXXzaflNXnyPdUtPAKPlP
evFFSxw++oAKrpfAYhcoZvWa/tMZToah09cYtxkcH3yh/F5zCIAktI/JvhyAuPQl52c2ESZL+32c
YKhxfJ6SPKLr7IsgVneDCyFP0bxmY/tdvLGGmrqRAUsA5COoe2W+CV99FobdEr+7AGXqQaAAWBWW
6d/pzladYDUF8YTFu/4YGXTnw3Am7af8SGrP3fXsl+OIXODUJEK/BlQXkWftQw1l41KNfxGw1Ts0
kAEa7BCmGgtpiQV945fhG6Pdtma3GM1iTGZTOIdDWcck++UFfeu3eV+EqsKYvlhruup6SstYVj4A
AfkJUz+GiaWKXKGcgVaGx/M3tqgBDuZoOHNzcUS8lm3ifs9CYTSPAS96EBDDk5TW2JW9YEuIxcn4
HrINKXsVhaDp/Vad6aBAf0NkuCIOWwGjr5dS2i0jiRZi3OHbWgaOlJlHpb1SDrtVCI73PB9B+CkH
oAdd1AoYZvoNQWshqCYrE2T0Qy4vweRX9PHdwSvS1sFftDGoKhohv3NFkvyFovylfGfqh/fK1cig
Spr68ocvy40Zo6xmrKszxp+e8+4zHvFBbyH7BBH8/2Q3zMCpvqjJZjzcGDxRCb5CZSuXemcDws+b
evQ71iXERam0O1YSFYalOjYnYf5j4y5SoC8Edrjlv8tgVhLAaVAbN2mfaCNDVGgGX0gYHEmSI93y
vxtS3BPaJEI0TNdYWWkIkQuAezbLi/Q2osSc3ets3UhPP4yONHnUEzAXePc+rozFu7SLljGCUG3M
r02fYYRVk9HoQC1WtFli+HW7qYiEfNu674gYXTUhYlChO/NHZ2mf8KBhjiQG+krE7uTMt5bDgHgg
TCg7DsaOejvUy9yBfX8UU1X7Q1aDiG/DgKZFAyJuwucfgc7mArIMldjTa/xPRccm4uaF82zM4+v7
ClGh6mtWTFe1oTidoPw/g6QbvtZkMFaCol2KsUP1p41FHZ1NnyOOIbcArAAKEozea2/m65xaQxU4
bfNgiExQ/uC//nVZZyVVYzwM3PAPry71zsgquqs93frLu7AJlDDRaycDsoubqvpf8fcRmIHMmWkC
y003IUiE9FGTOLi507UDR+nbIgZecDUjJhh88BEdmuPxFRtZdb68RhhnadmGmIfPnLK+fp69Psz9
eTI66X0ygVdHs1Fk4JpFQf66M7LRfcqeSlDtYOkJ72TdSDw4X0rIPHqww8YI3h8m0xul8FXxu+Yy
NZp+UwKJZZRM4vCnzsIJBQGJKEg53+yQNqsqosbB9P5FQkyNAccjP2GSLZvLL2Kb9Z/zl/Z8W4zF
Qu1H2YdWEkwo/D7ui4sKy9aCzbN1WX4ItJMlQyrv9VryRa2bMgB03d1FD7mZVw9rGheK4hVe9xeg
2dwEsVi3e4PP8Pjm2tAbKudFy8qLxJpv9g+eFZblXtLo2gsPG9OntNmxbH7Wpe40ZV0skuDLRvZz
0v5Xj5b2KEEKEMkCWtJMgJkKdas62+gY1Ru+/QznHr1YJHopomuHivoy7Dzw0krqj5MKK1arhC1C
ve9yJQ5ShVbNduR9ibpthDrCorKssDcAXXIz4Il/1F4gC/iRC3OvfwdJ3PPOhgv6uv9+URpW7t1g
slkIfrUos6GDe36RTF+Xr02OdQ+pZD25RCnX5kF4gNbkrKxtge9fyOSXnk0PHyxX/1YGTIzo8+wa
OjAmuz/8qTlvP1OyqQEcBhZMrMDcuxgqrH9DoVTDGxyi5RBFzzEgeq1+xE5d2P48xh+t+JiYwe28
MJ8M2CAFdJoRuZ59kIf2C+vJodrtgYq1ZXz9SCUsXK7D5aJ6+llhBmQsABEHR8AR7ZjUGQjVHGEb
tn6rFw+ilOo8mzxpV9Up2ZMCvq2ufpK+oUZOLwBgEJ7GsF/YPMwXxvds7ZsosIIStB2R+LvVYzfr
afa1OyCoPXCF4mMyVF0GiUaWYbSPw0w6iNOKVEMBEPlcTGkLTUQ/Yhxm9uyFYp7wV1Rw4NhNtFax
/iVvDP1ScewVE8Rx2iCL6nA9YonF7obav6Mmy76sB7YDdIv2RMN+S2ARNul/4I36B5fBZmiu5/af
5UVnB5N/3D2Zq3rysdtA4Sv6G3uXA3ItPG9gXHi6mZFRz5DFIeYqAE5Xu+Onsu+APLdqVKiM1dwh
Yt7h3MCYJ0V44UAgA1NqoVfinojaL/Rg+3HxOtbqt8qeiZymOAJxRWAs6SYVhZhahpx6mxppJPbM
0cQicQko0k8LceOSBwmYddhorIqI1xzMuyrxQE1adiZw25OU4jqtehVe99iXhDXCmxCu5O+q4pvK
GwykESOa98Q1i+e2Scde3Pw7J5ewVekQG1RBKGUQlS5D4kw/CwQAi+L2p3azqq5Abh8aJS6is2Rh
VS7+9n0aFhHWwN8r3MybDutozJl/cUs9IqceRwSoHwRehcNLweKfsytnWrkO4Jre2Tpaio5Ha5bx
kB6779HPcOsUjKgA2jILpBTChmjbfzv6DdYl5uSV9oVvE6b18+L9X3OLLlKDnnBrRfHAXpmtQjgu
qagrhqh0xKuLHN/6pWF37v1hiZcq+rGcsN0qPpgcDPxbYYYtrV6gJY5CZCaDBJRCedxib2/NS9W0
pE3x9VU2yyPNqI210jE7B58VMGbClI3cnUXUu24S4ZWCx9DxU4ubukYlpZlNq95613Am8705p6le
Vh8TWZyI9MupJf28MhlwpIKktWsbiBwwoaSUjtCVWohHmqZdo9V9D/FFjGAJGOqEzCNKSuu+FOF0
Hu6uQCAffZKgCMX7Gw3474ZU4EyEHa8tifUFsCC7tkgUw3sxJoIL1POFdKPUN5nI/WFV6rpVmxo1
4guHNPn457LBZFoQlDXuKUfAydLcmnv2XSHydl/SdYMtyUSJ4bW6AbTAfJC2Axghgs5G84YbNoL5
B8X5ygQd5jPk22jub0NUwiCjIO/s2+6yyUZGSBD6DhSL4sl/jmpyXbmVbleBe5l01u+4T0e4KPOY
7bqby76Q6GzQ5u3d4WcUhcyDZqgptaOi86lKHz/c2Hkjb58cvfHB5561xEwgqzp7HkgmyzglyGnk
GPuiZLtR5Lqz4grL/YeIkd9eGri+o4YFq8ZUbL/HCpvtajO5MJ79HCsyzyb1du91pt4f0c3/npBd
ySFO4D5sGBOuyyA+epQ9y5x04eYKbxZkxxlZsaVoQZ2Dyc1MUDudwDztYk+PYzDJR6t0VR/oLOdn
u056ERc+kjXfQjVXUqU4m18t9JUHNBCGbtDIInCs0+MzgGTyQSF4BgkxXsLvWSMA55D7dHkJVgz9
LN9I5LVxYhiF+0QG3Rb8jzYuF5qCBJvxp6F/gxnX1IaCcnnMuSiZnvg6CHupIGcE9YIMnZJtZG7w
o2Q3ND5v0bb1xsjhHgi+yh06n6y5XOXbhPaZvnJNIzxmxV5P4JCOda+9vN7UQhX8+uiimpytaGwB
t5orO3AOxSWsqMAU+TentfMELt3YbZlsVzbF3qvSrJoUqA9hbmDTEh4FcvLzCxo9Qm9VZtn8aZeN
Xjbq5bBqn6uvKwW3u8weai7zbsidTkrDuHs2p4j+CPoK4z0mCfjDmwSO2IowU9WnEb8kPytuvuC/
l5r6J+jTjg+cnhxcDaAjWxTqek0XNJWsnnEoqFowzejIiiiQYRsfg1+81CPJ1uDFb5Gbmp2QR357
0adn9ZF2IsIzXmXpKXv997WI3F0o2gxZSQErfDIzlztdVEcwPZyis//yUl+xvz9i41yb0+E5SldX
E0h9XeYow50DyoldAryMkv/YOME+iZ67kX3BjpXemxfrrnN/AM2v5HUQCnzufDlxbDJYIECqoG3Y
0n2XfF4/hwW9GjRh+VkJXnGj6ZvHkICTRH5qgnc7kXjI36Ic0VGN2ckRCUs8eaudlGgvA0yq0ExP
Lf24oBm2uYdaXilo5JGUOHjDHHJCQveLRg5wEu/GWSVN2kIohfZCeoppT0RxQNIQJRAhotrCgSXP
7aVx8LcLoufIH5kme5LFU4KFKwdJh2lWCs20lHwHIQXGjR/WL8tsFchj4+jAXFOTQzxoTHeEDd+H
sVlmgrv/tK4KV0WHz68OLcCKDMUpfz710TFT5g52G9UNf2uOaCEUEAtS+/LajmzvxER5wD9g5YLa
UHyxT3bY/m+/Z8+Dwfn3G4CX9fN5XRXtGX+Qq3xYoF+auvyJ2O2zw651kIwvZ9xmE2sJH6YKXxaL
z7gObBBIjqyAxmhzVOlQgeRB8HC8t6RYXh4rEq1BNDP9r7I9Yk/CBiqJa7Eoi+4VFinCBbqJEL76
Or9pZVuIOHOgv884a6w05UrEEF9ivXh2QlRImOgjcQZqekfgb3+CRYEHszdD/EP9cg/bWXX+Yo6/
ySpoiPHN7hOF7saUwZDuK0ApdvfFvbAE+tnGCVFRHvVyHsFYe8p1s4yUC0frCHfntmwq84qOWszI
X9zggZ4vKmZ+Qs0+XCAHvArF85uX1poE+wagrRm8YNj/cDPDV/53DKYD9PwLEH4mt8+PGpJiFvvG
i50VnouwgPyolj8A3WIYvXDcc2vqkaSyWpDqVk2bFUV9MkX7ol5Q+tNcHsVeFWqZVmqYRFgAoQOn
zeXTBoEI3zwLRAbED1fFejoTYfMu60A/QNHbh2wXbtlbTkBOC0Buth0LFhf5Z6xfFHzh8TGcL9sN
MtrMebJCPIMwNULhK2Bx9fgjGY6vOcKf1QQt+0VVycLdyLwqhavtvP7P8u06iMd0pJ4HG2N7Ketm
YATNbbHDSMRWGer6hdXboBMh7m62fomVDBVrHNWtasmmc1+vMNEXr3RJ37+6U0AbMIc/ErecspYi
5mwFd5bDZ3RHE6uZ7t1HZzZQKfqseECY/5iDA7plcOGGQfN/l89DOuvK5GYVLUylzch55J28E4n8
ncAJ75wKMGmQrFTAK83gnvOFkcOmvIVmdxDEDxy7mfUgRH778s8+6zcZIHkaoPZ8B2f3JHjnpYJi
oTK2wHnrfinYHZt38cGw2iSu5aPlVzJYzfPtIOJ49NZ8Unhrq2ME1lZvQfJnmXrr6N5r95IuejFQ
C4eAJebfiZdsUOrysmYBCc2sJSct85ftWxQmUsvPwXsm2F061KxfE0js8lgbqHtvJP6koWmQmoyL
B+L1fqNrusV6/HLwlWbJBHmXDP7+shRGRAVerhYmRfShdWQel3GfFY7mPG7P0j+eWT70aKYIdhM6
b2WdrSEDxz70CdLghUZSC/mffcEBKNw+MUObri1y1tf0zCF9Y07j7IKSwiqSUIwGwL0IGYqdt88Y
4OueeRJ19JNoYdQnqRjHipXVhhZyT7sdGduODdzoEuo35gYHfXvzbmlnO4Qh0YVtcaRgtmvWEHse
FpLKigKnqRxPABnSY2X1xvByCnZhv1EI8kJfk6iclnNJNTjhvUUdTqxtpdvLFWhVIFtveuADqzQs
TykECFT6brEqMn2Yk4u0rgJL0J+FN+lRHnnVO/DgZXmvP2x2HpJm9kokB5IBdCEXbeGocBarRAs3
/WG0aOjo8RKBsbfOH6N1kt0VnB3qMC3vK3uwJQDdoY4IEtfwp7wFOcFHGucF7slK2TLFJIdU9eQl
769slom1aM5/Inv+v0G5wFfgWVdgjIFPxvBQJW07CSxt+K8r4GRz9JRBDHiiGEcNwX3LRt+mV39/
Dqwr8eRSDiyMRB1k5VKZhTMjZ+yAHP8zownBTDkd2Mm3KxEAipje9lwerqKOOQyQNSkyd0xllZpb
UX5NEWVftO56BMhfQ3tr/rfPSYyf3wfNio7M8a+E7qLpPOV+F3RRNGXG2lgi3UjG7/Dzcsly9H4l
T6cT6iRXYo+jxim9EI/UNNNG2AZNEttL3aTlW5le3xBGuV2v1Ax0dJDdGdLdxxTN1EqFtzMyvtVp
k61u8KYMa7/nFCyDGQ8UVrAbBXRBe5d01ZtIRVJ/XHPcMHyTeWzpM6K2rUAd7Zxtmbgh49FXTIc0
UnmG4j9DFN6pB4/+osPHYWObpiolBn2LPcDzOfScqAYhBFXHCsqG7exhqNYQ6GQSsVtviK9MO+eh
7Dck1pgZsCComHXL8SWPpAS3bI9qLoypG7DGEstofwXyR1B4ZEJXQuboblvdvp4XL/V0F8hN6Lli
I4Mk13xmyxA/F1sRZ0l4639OoDGmHKOO0T5n6XmJ59zyjnRMbcXcLxzWrZmroF+n/+iG29Bi9GRE
35NkhhYCnd57SBJ+e5AXW64H+tngtHesjZAC74iCxDkZtrQG8M5z4CssnYef/PDpdsDMPQ9rnDE/
stRTd5Nm5kfFxWv7DdEHMLsB/Sl78KXZWkDYV9uWesyqJo1Jogl3KD/ogE0Zrvc2fq9FPNwpsHHs
AkG09IEJopL7acdBxXk2z7G024/QSgpHYAdnlPSeqqKajXHQrXY0yRMCsyhIY8gI1YLwjCgKiNs7
CqNMORqvf+QFCxDtQogQ4FllVJMwimzfmy4+EacptcKY54VDxAS1W1qMTHVIW1TiTj3o9JA8AbyM
IzJbqeXyCiYYbFCATypzqfWuYI1c0b3n0LWqC2U8kBSp6/jfqYL78zD69D8p6x1NKcnP26p/hdPc
jbVjeHUIOllStrSpmissO1KVL1G4wmhejxoa+95glm3stc4mmY0LhpCyQLtv2bdGA3pNsSv7Xk7Q
VRcvokd4OltcCv0NT3yEQO7Rv9B0eBmZ/QWQ7fmAqbipz8BfY4TmvUzvWAcX7JHAKFpeKd2Hn8Qj
EAFWd8yzMihvNf/lcbWUE07xGMSnDqHjPJg5c+XC2f2kd3sn6wt2hRGtFuMvPK1aeagEDUOoMfWC
MQgpgvoHkLQASQTS3/Jg1ncAPAfa3NOf4yYBMWTevrUb5DBclb23K/hDJ5D9m2UrH9yjGZiSHHxJ
UeUU8a4dcz6TKVpKyqqrh2zhGZ7Ev0V/hzNP26A+Et+5pk1ZWfdWn4KiGMEDbf5drwQxGO7mXfwq
YITYRPkgFZlctlg/bGaz2NkhS/7GNqUnLXCOyBxnSQJB4Lz9L8Q2yYxkqk+H2HQH3v829Bzmtnlq
+q2doyteqQFBJoPaWItaT2iIbwXizwBoO41mJCOS2PbwaXN7vV0ITHGx9ORo7QLRQScCOqREdCVC
ay/IDUN0S43XTnXps/4D+YG7Fle2UG36i4RgA4e1ZYDA8SPOzjyJlwkqgVRLq3k2PoCokbjPFM99
eS0E6gMkEO95gg1LiWrwC4ziq7A9FDwiMTYqd6yzg0idT5TDwFcLnB6QPAMXfBx+fON9wGRWaFLq
BO9jpl+LFblaas5As2VjC+FbMGPEcaRT5VVf8FEzOE2LrGEmwvzNKhyTrITrdCHfgkRcZLNn1We3
wrP+tzrFIN9xdrbUioDAbesx/gjTCjVuMU1NPwwj91BsoteY3s1jVxQHzORwXGfA21SZOWKUiYW1
b3txmC2NHrNYNMYPKsD0F0F0lZuOb8Vw7GHkCsyTTe8CxPYUEqpN2N2nvmZ2gdLAmgbxXxv032wt
MmDLOPj5QcCPtN0dn4ohS82OMh67kmf9Y0KMgmsqlb00ekmOTrRrXa3oLF7jaayB7JEV7Jljm7b2
LvG9YfL9lE5V143LsriClcUhOhdG3vEuCqo7FmzNQKAoG72Ax3hjV+FEzPqePbK+LMgZZC1zvIn+
69XmhAd9duDbP6XtylPkifBO8Jbd2UB2BRGolwvhHYeTJkmeTcj8sZ5om6kPvN2DOTSwrrgnxVx6
YiiQHCXslxn7nHRupiDqvQeLWuFmqXAPJLVgkE40E15gbMlNatFaSYfX8+Rv655FNK/ZLMqw8CMg
yckotZNy4TpSRvTbVWI9YDvcO7bTlNuQ4mTaC5GatI/iNSlAfiM10g6eTu/3yyM4RyN0zDR3UAj6
FvjrCnO7/b7fuFqeJUpO+FwZTffpmdLl2AQLw4A+qc5ImI6x/OKudPB/Zwq7RDX2BTa/34travKE
OTnYG04wkzwxwL4XG0YNzcemMm5+x0uKI8S6vbqRLtean+fdxmYi1f0Gg3zlzLDoWU8NF7Nk/ika
KxRMX5AsG4X4ac0U7ldyOK4KAAx3tMGMpO6s7ofHORtWhEaenyMk1EwK6sw2flNk3G2e7k6JZf4T
P80rxTrOsmmdfisTEL9tNHVbYRhNyliyg/ipKGKy3BfA8dDvWOuKz+UvSan6Px5qSoXqzVb7HC/A
8kThkw8vm7yvEO5X4tWSCHDnU5kLj5xYrVYLLnwFi+1HAp9YtMnawyY17V8cTPzkoZTNMn7U40t3
EtphJJXLEH7z3IH95wDBgxHEBGb1MPJiwtR4Xez1ABPFzhi6n+n7vDxp7tHsUcT9Wam/EZ681EmH
9D8rW/PcRszFID9atukixocpP/WYVIHoyYoY6qkqx73yU4jCl8OZzMVwA2t/QYHmgKFb3rTUeimW
tnCkt0TvMg80hcTL3evAsJZfk9nQ1rYhMytRVMeSb22jxy4RX7dCeJ6n9gkZeND7S0sNJTxqGO+t
zhPuM5TCFeBxO3soS1EfOylNhRzv3QTO6HyWG+P4zRrn6WxO7Z2tBgSPbAoskes/6yM399fkM5QP
nCDB66/I6YQqxt2MY4lf63Fgyss945J3Ihv0VF8YOBhitEI7MRiIpq8dPuvcPA6lREm2Vc6xkzNT
43BYcwhGqugn4V3NEGUtEs0XyvkvOwhM46W/nKAJ6f2HUqgGbGIppOg8CU0hnupLMY89KFyI2GSL
UtN1Z4VOuw1q3sZv2hhdPbTVSZ2obnsoNhcjsZpYf2A0cFbQ4liTy3x41qVFpiAAXG1jYHA9TjBB
7lPG1o6cWg/BVJQvFCUN+u+Z8+q9MB9upJLq+d2r3rhAOzCagE7X03hmpUL9tKwUBLrOuvSP24Jv
fEbnEwqu9jtWtLZ71nPiKVICOP44YRVBcTlRnzk6VB5eC2IkYGWH077VgEm5gwnZHprFoJbuIHta
qLdHr275I38okG5VLIP/ovLhNSvvv2VXiY1ik4h5y04t14QVpQ4rGDVRzyxL+WrWCqhBzMrhTaBQ
01VeRWDWpgyKOQ2POxetFSQH6s1zN5SiP2wIjDYsmTpT4SyTOY56NOOedfo1h/RG05ME8xBVQ95L
vby5ZyTQzOKzWu2/XSJ7bPTQ6FfiQ/Re+y4bWYvYpXV+m61vHUEi2kdK4+GLssl76aP5mTjMOWb9
1Lgk0BncEJ+1eZ82+CuVOt2oj+YtT8QcJ1HY7HrptVdfoWeV2qH1BXA3U2z5Pn7ZKbvxH/IBknXL
PPgPtJCQiFHlMb2F3jehPE3GjoLK8D77uupj5JsfSMf7ZPY8FsUbdKd7B0YFG0OD+b8wcJnuyC5I
Rg6hH4pNmgK4GkPnnpuQ0YuJZ3LYdoYIeMMm0DRYNAaVZlKjfLbmmieH+08M6Qj/9rkbQj9A2C/3
NowVDOKwjUTuYVENvn+uM8L5d4YUGE1EKkWivXbpMlxfo2SBl4DF730saIQjCivz9L1r3Vi4YhDa
4b9ZG8jFybPyP9woM6J+BnMNgpASsWKsWNkirwURD4q/kZ7JUdcXBfYzMB1WrdjBW1BU3WoSa1H/
ky1yQcUvSvK434nmQmHCrp+Lkss+nuZJ/6cvJ3ILGd/1SRBr6ycbfVnuMau3JTAG1NryO4Ykkd9l
DHrG2yt7Z2j0oJDaxVy2FJoR6xcbxYmypCBExOdvkNLwmxysgpD8R97VfkOGEOtpY0lPUoQq94bu
dV/jKqsetl3BXXkP+ft7ZeIw9JhTxPKkpnn6UBMAYHo1MB4bLUlNh0AvEvZG4eiOat8sJJexI0qa
/Tzo3d3Her0yoKSGrfDI1MmCqnqgIwjLM8AqLdi7zBWMytyPcx/JBa2oEHZE/ptdth3eQ5kYQwCc
KZIOxODb+oWEXJq/Mpnvsj/VRTgw7+N/qvltJOkZfW086esXyewc42aS/niYVL345yGmzzBjpMGV
fEGk6lLxEAodu6FVhUa2F/wAhlvYvvw37Ux6750malC07N5dNts83mlOe5iGBgyw5jM0PVSft6qn
m3DCXHTL3esIWy1VFxaXcUAfqrujcZfV+D61Sq8AiBD9yf20UltV+JplZ+68yN6ecd3dRclaUjvA
/hhuKZCsIeQlKc0q1lNSuEhiyRQzQh9qemqR7Is8cS3A3Ymk8EEpKngcsSe1E1J6wrydp7W2xAl4
3G4bBStdfMgFaOSwpqWM4DM1Ufs1ht37RA8LxaRBkTK5nocBSukILvvh05cZblKJTXj57JVTyw2a
/+Dh83lF2TucNFBWpdxT4JPBHp2MMaVfcV54/ZwHasDe7p/qFBQrRWbqA80MI2otiNAn+iCbxhhh
Ko4InN6w5WjAAfiqO3+4oosw0pWhti2bQgG3dfxmlIBAUk78zhfO3Vk2hS+fWzpqNiI5j0TqDQxf
1C2HrqlczLvWs/I8YCFTO/FL901FQWWaSs3FSYGGE5IvqYmDQUuLNaRg3NW6gL0Zxy6i/9zAXrDC
7F/AjG5og61+rEnM++wN9tlYeN46+xfEQl+rKDe0anL4SjmzOdiALBRMRhb26dq8kegoipGQeba3
9Xb8Y6ZPfY8uXKTmaQkBH9puZkXdQ85OLhctaK+7zhS2ohyiqFSYu6nT5Kzi3gjmA5Ri1ZzB6dkO
wk/26Z0ysD1xr40mUD5UfT3KbGvCJ6f9mT8PcwZD8Gt1PonQwaE25LR3sc60NXSlSvEwvIeI6ECE
LlfsbRo4kHczuc76nfFL+n6Lw5HKt2aIBTVASfRHIFlybhNZPiBNx6zpZC9KwsUdBJlbcieVHzvG
gLlFJoNgr/3W5OWYSU+CngzzX3aFi5y0KYcTp39WZEuQS2JvW0X8lURoa40ADXjNnsT9xXYLB7n1
rIhZUarT1h5/4+bg72rfAFBlS7BQgk+LpyUTG6nzpskImjBBK58DaEEl07Xk/nFYdE5kdbIeK/A/
8yX0KfFjm1YyFZ9vbfighstuoqwG87PI5bVeU189y5iK9GUFTwtweyE9fNu+xjFjETC/Q3EYEbmq
w932BryGSRBHEvNVqyEQngu5kSRAtHs82D8kF5+vuvTYE8TSNDMkLDI1aK4Tjwm+cnq3ZX6RX8pu
7S4TyyrrTTowFyDps91xZ6AE0zUf76FmwXxeduW7CFJ3GblkklUAnOZtJIHe3uwyYLZMQ7KfO4sL
eiltT6lp8rKIXXmXFlz82F6cfeglSJW4TpGBjQlEZpjRYHfoWx6n5oohdhJU0ylXEDMshKLTlOQt
SZJ8jkbJ43a1dLYTaqIxhcfxh0Gxp13p0UqpKVTezp3vyE0CXkfSD+jCnxubVoozbjBBqTJXXQbW
t+McyNGwi3U5tntDRVU0AU24udUphUxbTqzTYHD01l5p0YNUOOXNg6fI78zfI65bAP8xvuNu7kXR
gjkkT4zzGv3bAn1Oh4R/y2kwIkp3i1GaDwy7dgA1Yc12cmz8UStLFC+MV/BiFVtpyssRDE6kJBEn
NPjjrdA8UAtypGmGFzIRjjr/EhQZIqu50t/NeCL7HyeusWczAEGpl1e1uajC1O88Ov7XT5UbAc1i
Wv0iQ14zZOwEPH4AVmwXYqBd6COdwJhS8nZEyOv3yC0ktnHPNBQKUfvQm4hsbCck865wFarJaEH9
jJl+1un9uVFYLniyHJCM93LJVuaHvnAWFGgZqRgMBMSe29CpGUfngfV/KgSV6GAQGqOMRzXLOYdA
gLEZ0thV/PFrlRI5Kt+KkpIHNOiTas7Dif0wUvukkOkUtYUhq4We6w7dLj+d79DS1QrYSRK4bj4C
aVGfLDfFNU0PFNlJnMxx8nkcfS5mzhz3Zl6EF+MYwghVSJxfP/op5NwmAgqYa8ePcMaiRSq01xPa
F4cpNyBVNWCbTHSW6sh5UUjEMwwVPQ1H996R73ahwbhXdjE4ltXG6MmRU56T23giT7kLoa4FW0j5
TlUcUZOnQ7CNxLYhMVjAaV7paTVU0M2ftnQyxhK5MIzeGp47CzbeGUh8ivua6mI4iLgvUGq5ESJk
i5jAVotorU+IR/ML8jy55N9UUe98ds+EIzlO7QDNZeyJmmwFMpaQTivX8Nl4xn2yENYeOeE7K+8R
+RTjzOwKHiC14XykKCyfsbs9ghmIKXCnl3R++LmGJ5I0s4IAgQFW2Wiq9qf9UCDBFT6NjWzrJyhN
d97nEkgfGi2sXRHgyu57nO3cRg+jsE56Essd2+T5lUFw9hatZfxa28UozVscO3APoNDtaFm6ldBR
nn68cxnn/BxbK0uN8LmrQuVt3n1V43u0Ek5ri+VRClNewE0gGaB60A9HyeiWtnKXa8Vai07wOhiJ
JWSvl80JcrV7QJbfl43QUqbZZcbcXMRreReQY4tctO12Sjy0SNzqVZ4vQu460ybWTMCiy9f85N13
35uZltNJdJ6Mn6xlnzQ5PF54kzPZzJ+DbDmssTO82DT3awFB4y0xOv/Si9o/kgCys+DBGmRSbxpp
MkVKCRvL6S6vb1VpMWdTEebgvhfTj9Fzf5UQbiLv7vsYrWnPkKGwklsqJ7aL8Gn/oIAyGkRQDrhQ
4lymF4/fk3QPPStQS2WSTq9gDVb5EoXl+5X/eOc6epwkeO/hJtAC4mlDrxgz/S3aS2LU73QEnko5
b578b8T6r7OmrPpws/Vz088SsKqa0PtTezxdsoAdtWbPg056qEjtgQGNymBmFY6We6HVacBdwbjT
3qo2LQxbPawORVDZiGRBU4yq4AU9rgxfWMsRvxyMav9eKZ2h3qbfI6+CSBbUhUpbMiuuaD0B1ALj
DA4LEP1Q6QpIZniLHL5oq1mAOVXxzOVhJZHdtTlmn3h2bY5DSSc/yGfv+AIjBcrVNITzCnsb7WpO
ntaWLAQZtVO4XisEv5XTKQvEa5LqbUlK1SdiEX3/XWLx3swptvLITx56d7rjApmefMhTXHEzLWgu
YJeNEEMf7ldNCHdwj8YpKgOjMRnMhtFWoCc8FHPvavhdBg1QqzuFb+vi3PxKSZF7pjTY7ta5PKrh
KmpXYGrxi44zX3iSC7XBEIqgbzsU91/MEPPNmlvYSfHnJJRGMVxZRqWhM19nAvpK8tgm9HnTyhMO
yEyDRcXyS8ka9sX8KE1sXQOvlJRWRamJmBKO/4PiqM26VYHRcsGz/lKs++rrDjBybjzPoOob783Y
tVc/Et0K8GcrztGa6LI5z8VxrtiwUS8j6atUgAX2iHOyRIaL7L7Z6cwQTeegWcU2w7Ry6C+6PgE+
/8FEzsr5QyT8AoPJZmR+wRrVleTBk+Jo5KhzeYbxQQl52THZB2iS0lXV1zZ/UvEgUvYIeIYsxHAl
SUGW4l3ITO4gUsn0QSL9iCmWEnBAS6KXv03o8X4bob9AzGOZPHRgbsxGSlhCrBGsh0Cmx/Xy6Y+z
xeKLvuAGDr5Y8KtPQkOMA+5eBDzI6W3QaQ30WNM6j6HnG4DhT4cpcLIryG4skHg/a4ELLqF3Ooz4
RM6gCFB1EZqSk/QiLIBNknVpTxb7ioqSsNjiNKUOLx8sZJep613RLr3JKvd3jNMNZa7Xp7XxUiVl
g2H3bvqBAd/YtdMGyNRCgJOs3C2rmIdnvS47ptzIXEFkINK2Njp/dW5Ptw4ujBnL8Eb2xWFJbTJ7
BCtztzYpWVm4pFtO0mktxjyojKVlXcmIt9x5DgeAFdA3kR6JuitAT5MiIzozqN4oKriL5k6hhZx/
hLI8QJqyFyfFTriF0LJsZ4+doTa76AgpVXniHxx2ag3z6slgp/Xbnqoy8ohVAFdzvo8bDPxDuD0T
P4hc9B2m+Yxj3EK9h+NWeE6rQf8JQ75koOT9YUPl50BADWjBFOkrefL34CdA2eCm5uum5cEcuNT+
nJFKNAukbPNIsTV1yxLnsS5QokLei2AMP+ikSHXrs3EsAcBbO4R84WURRU7yFwU7Jfx052oujI8s
j7pOWUtIJ6BrhOr4rUzUrHlGoBzOrkMU/JCAhi3QMWJV+jhWynXUjNoq34eWZd/495F1zW9fYspi
PSH/PUQS/r0P5/EPgOogqcL7bSYI2x1TmA4K6iLHpsqX2lpvj0hgSmHnYU9jyHnfG6IXKLPe7IyQ
QugSEYDEwDsU4kXuCSC8hSoMg+dA81SoSwHNgyc85nfHfqsSPgAeOy4lDQM4xO5JCzaLFCICb//Q
qfMiKoPhdQuNkwlCROmg2tB0MPJhi33FGBqBnjRD7R7/uXrhXOnZ9xZvNSfhw1BGE1DlINZik13t
5LSmJoUPSESxmQ0+CAV+kdnDlZvFaTr88W4+j/7D83eFKT1su9hmvx841lQsuE0qGT6z4TUcYgIP
WN5QZ/il3Aaz3TZ/V8bls8UbJAxgvjXWJFXvOjwouJtkdzATOJS+UF02mGGEN94jFUbe6BodTxjb
Tg2LdNA0Hx4zFK83ppmPZIk7WTlMPBhk3i8sPGKD6e8dWRyIeB30yKdmBwJ5iVogjoFo5n89VyEM
KPqFoot3tstNLawbPiSyD+mNY6zwWiSGsGVdmLkvWL7e2GHZFE8p8JEVaDL8Ndi9gYKkJYFV2KHB
Cei9VeBSh1NO8NfEgrJo8XWXl+TfBivWWMrLrZdfqdjIuKRlZdkVAuvhcmAcGUD7S9IJiAjO7uKs
u0GoWss0+BIEkwD+sB4OCgNL7pp21iUMrrZsq9MPwrn8SpYnv0U+6x3pX326YbFnW+2glH4KAA3i
3BMVMgh1/u48t2DEAzqSNn1lFu+hM8R65qhEcnxke1iYRX99K/Ok0Enzw+hfgg082U+8u2qCWU58
8keWKKMaBUPxyr6EnO7B6BXV3lgWNOd8UahiFFZsvA15zatzCVQsHQ0DEOwlf1tDoc2ZCJU8RfC2
zxtraMPeWJvWty0Q5HXD0rYeVDSBxaIlQ6VrAWoEQOTuByrkKV+T4F8QuKUHbNpc1xW8TqqNdbpB
VuNrmLYw6elJLBmNa2wF7B5l4ODYCKnzPGIbRnUdQovrt4kSGmbrHuhVjfCFTNHQw2jhJvEZyH0W
kFS+VB8TXEm4OQ1aXd8BDQhDKqooPhswU4fg9v9Ze4x9nBwcayCTXt2sKZ2hwHG2nLy1QbfT+wJW
Rbbjw+6vpXC6c7tDXCL1P8hFLbub8Zq07RoYwVTFF2RvsoI3OYjrLAwVLVX2zO/I5fxUup5TDKdL
Nd2yUwnFxiXP7woDz5VU6kAfxqrBjO/lwhcKQsvpwQNYOVSVRr2cEnNnCk64GatsATNFWyjTQwCD
ZuYHMXRXqQGe2nRq4B5VQPx9rNcJ9nM75pSsHGZP4sjksUuy3N7IJtZWfcCjf0ztjBEShc0NAtOD
attiAozdkmXcQVbzgrxp4NyBovs6mIlY7bvlt097bOHJ/75TIeBi+cGcibTyuZlQ6sFl1HeTl2Nt
nA7gUd4uq9MggV9a6ep8Dk7OtrjCNLya66c6KZ9KseAogSt31CoI53x0/jUe0qxNWE7O671xw5fO
OCGJ9q5RCEGZSeBlRWZL/msez63BOfRMrbVI+sthjTFIKpmbcL2wefaS3GsIaNKvsWCBx/CJdxUz
VWB+qs3X/uJ4ECFwGZ3uD+FlHL7XlIiF7bqdC8GquzEcS4l3X3WJvzyMVamqtadXjQjHmSIlUpwq
oXGAL9RaIOA8Lc3UERGugqyAa5pCOxVWKQY+4RTLBs9uli/XCCaY4iYR8wSwsYL1zMW/gJYOAIgZ
GfaEnYcrGPT1NbDohhAW790bu0PTQUNgVAjCH59ai8K0Yt2U9gVj908eUzyntwx9iQbLNbwtYH4Y
aZUrFW40su7edsRwgTgOBrQZWm2q5wxiV80vaGERvEfVaHEsPQbq86w100wDW+skFSfUNCLhhxi4
YFR27jhnU39fys1xn1kK/iuZCx0NTOIn8rCS/0q4qk21MrNBxE3zJNZT1yv8UYTIAzolWJ+6hS1A
2pbtzUYwgk3e/7Io8aULKCXNx4CQzWTPpRZPPiqNacaxpR+UqrL3B7GCvY0pFpBeoglpKN4CoCZ1
a7aybA3iPxXjd5eim6inaJTHhHC+ysZzifwjugIQTtbrbz27VYt6BkfpWauToKFSoI32eBTrO8SC
DnzSK0dkoSJlE2BXSADi3WNxyxaKdXCSA0qchMTsuRpQJJ3K18orwLzCrK0AXGs4BkKAsMJZMsnq
LFVjtbkdNY/IsMiqcxzjOIEmn/Yy7DLPDlWAyhgvEZVGmnRxI5cs8yYe7ZH6rPosURUFHua9Xvnd
FvzeSRMheEBuN2ibiUCUPpYqtfTKwfqtQIaOtUMgqwMECx/Km/hm0a8AljnLdJ0rMNKdeC+qHUm/
i6NKbdhKL5v0CBrjMKUUDqQYzCiL9LyxNzfrWvz3tbXmZdqWz7YjbloJn+xOmaC55NovPcmwCek2
P9Nk2Bnhrb3uNIo7iz5ALC6YEdGbAazGLhSYO8LSdHZl4mHKpE6e8UH/sZvBssqqC37HY5GaqAtO
4TpZKLnvAmUE566iUI4pyI32dnWByPD+ox0M3pfxnEUHbxlo+Fv6eyplR7GUhGKNUqGeeEbyLgMi
//bPnx77W1o3Ur/j6fFO0Jg62n9DiFeTveHFzB9+9myhqs4j/vBgbZDOnAoBoeWtemOJanJnMVJH
rQdrNsz7ddrhI8jxKdSvpr35ll02qODaHDFt9Rx92kt6xbQ2iZNO5MeMT66R687JmC+ycIARs0aT
5jMMF5kSCV0HM4KRn+1YQMODJdsPvT5PH+I9PCkTflRufGAKPeifYUMTtPZGc0N5MyM8+IqK5iKE
s2g1Rk6TB6ChNmgRqHo2U5E69AHM6DL2rsBV/dxlaU8nJ+LRhud959KbcukeHOzoFtoC5sGLZPp5
9Wnyd7RoDfQyPN0YQtdfRYZpkMrVMvLef5nLhrIkMc2+QS17klfgwkJxbCRN1ocoUDZw/7hZbHZh
A7A3Q6Et2jv2Ac/oT/UUojFY6KVIlYTx70F4/hEMHkitTstH6CdBdOZEkBANZQaxLMI0DtoIh8Vs
l+xNWWwy8iBWZdLAkK1GOditC3AoOrmzEG4uBnIMHoKqAPswx2JoHh/NbBSqWy3H/NFdUSchT9LX
cBvk/g6ieAIdX6GN24OL9Y1cr4tFCbZIFnsds50NUPINOHal4nRgoSTtjJlwo7QjIkGc8pGqbRKr
xMfmbHheLm7J25dA5ciddUQ6/yXgMxeb2ZFB1GncmB+hlGtZVypMvDemLggZI15rNkXacm2pMPxk
46+5p/IexeVWKSKr03+li9VhHQp/vU+GY+v5dm2PkNA4gWmHHR+enNOdMj/BYRgxwcCWjDwvtwm/
XGiCsQlLtaB5eDGQdgX4I8i3Lx5FdBk5O7PzkMLf77O0xXGenxzcBZG1WMeum1oza6qkDR0zlShK
9izCLkDyygI85PUuw4I8FyDRioPFE+b6Wj9XoPcDawjJPmhC9FoJNVbapZZKsCz7+D7LDSWM/sBV
NjXis04LHP+a6yX5JopGFL29W/OVpkHuw0nQr2WJ383UGZwaoDL0L95BDgTp+KR/HhGFvSSSotOW
oCH20qxD1s9rDUs52d1bJr7Votv4zom5GtyhI45NNP7bdKS1ee4k4jM9Up+ygjFJEsCasmXeJ5+l
zyHQ5xZsWNZCKuB8dHOG2IbfY2PnvUkTv9ghQG3Xmx1IFE5LXuVoCj5gZzB8/VAHUOtf81dPuyUp
EdBYlwCM48NbBuWrtakBkZkXnvQQwqfxIJ+BoKA/W3bbiNxKc7YuEWXcE3/0olm20g9cGv2RgFkz
c9d4PZYxfg4/Z3GQP42gywrk2qDfsn8fFSDvGClYhystRw8rrK2lmDDe6c1hS4A7MNFz/ZIY8izr
pQcCnxVEIVkhjzoc9J+bZBkmYTdBZ32DjehlSbXtD57Zzg56/Faq2u59JPiWzWPPZ5pxAvw8bXhK
HwwxtfJHdRemNox2qmadmWOMkZys3qSYdOWPEksTfXLbvU8Mh7BUzV1xDSPhbXPFxHQcMfltI1dY
Gbc7qsCDCHgPPJN3K0MTEdduaOPEZDXE1TRBb10V6/ToEziG4t1aMBOSBMFNAlp3xNw5N9OGrpei
bQEIwmgDrSUCmdto8FpjjmytXRK2GzwQEEReryvVILBN54LtGzYdcmyNl9Z8naeDe8zS6nYZ+H4E
YT6RsvXNoAnBVT2xitnh+Io/Ehkid7xx4Rb9XPpspsEf3eNTvvMwKkIOCzQCM4HJ/Icc89/7LxnT
hPpe5GoGVPQLD5JT0KMnROUiqAnVCcEgn9ygXFwsESPjYVx7l5JLoz86TcAAetZeWqp471+Xq7Qs
+6qlGMwHpaz4ROrek/ReNmzZ0se6C2hMqSs7p+0+Q5Ol+X9wEljuJ7zXA4DQbADRniNWHKfx5Dv/
Qud7sIXqaF7q39kTXiNoaTpB42p8nerQGG5p+xlu38gEgDv/25CutIZNrvd0a/Fc8ygYaCSHzJk4
8uClYsxwYCa3ZdD48rJtaDcja9ITpDGm9G4//SQbFKT5oRBTO1YhzQB6cICyv+8DBkeHs5v7jsX1
oV4csuDAVYWCXFV7L1i86FWZ+kT7DgqyAeHF826QHsoYSuK5dCXIqqUqu7W8btnHhvaGwTLgEwbr
G4Dn9glYu7XmXdUK5g3EGMDexQRjtUm21I8WuxKOjVD/EEYYAJtKtWVOOQ02a3A52jF35KlMSA5n
9oJiWuck8o4Z/6Na2YonJ4D1o8dTC/DSEYOR6jqpohCXlodWC8evJ9/uoxcN6Z/1fLo35D8I2DGk
IbbQGM0RFo1Ytq0MlyI5PmT0onzba7gaYAMOIOqXHZcxqd3JunVMrbILI5ApBv5aPykzXZe7LgKd
UFMCrnH6cyq+Ugw7mNQxh4YMptlsYFM9P50MF0FPd4/69PewRWWsPsQATBR9VfOqiX2n8Zsyy8Np
95F9qNBNSZoXFrSL681iAvwU57krzCXZx9azLTkkB5csnUzFNPetsZ1mRG1ICSxmoDIQ9CjJPbhn
KU/j1Kiyg8JC0MrSvR7zst2VZ11a0GAQPjLB2biTagQxZ7/AzNm6Uf+lfpvhwQtTCuAion0FxzNC
InUWYnUWDf5N9kRnk2duZHQzscLxogsSszzn3XW+jsm2RNQ+6C9FiQq2DE2gNFIpvtz0sr/92A2H
g0rkA67OlNGpLNgqIV4TRqooipZanGucmhaGhoiK4WTJLjj5NUGpWfylPvncmxLcXZXZaHu+2/u2
vVcyy8qqR7cW/dmHiDnnBy9RfNrzrE5UF8v8hjEjuXF39At+10r88/nyIDHbl8dhkEx2+3vli3UX
pj89mgdT4iOXT+hXtyeR3KpPk3GzFKmydbl9OmWFdkHLzCzkfWyN9d+Ym1/Yyox2DR2sCGY7K/jw
LU8jA2tuhjCXzV9mfLgoNCV+IG9JdzXnJh1++q4WmcDX/FOGpe1zO0E4mXZz1Xt59HmrDjK7Eppg
pnNtwHLu0swrN1nlNOFvp2IWMOLlTk4sT2dc3zpmBQ3x4MG461jXgAUgbaGdmxZ+S/UhBi+pk0EB
KkIvRP5PLOMrMA3EgL1Npbx6n6JdBwqaKujTChtNW+YXkekfyWu2WzQk1hDV21rNo57EI75nZVPi
6C9NNhCNk/LU8dyK3ULvWjcIhiuYkrKEwgQMkPC7s6MOoGYG/HmaWeMEzGgy0cwExEZM7571pFKL
+cf2e/dJKw6OoNr6+jw2Z6jflqlTqsYT8pTXdC4/JMol+81Qp9+I7tLVa2Rd4G8cw5VEwO4p9nKx
Qym5/2Mhb6FgiCVqyqnahcwk2kMjW9Jy/Et0vZlbMGhCaZb/oH6KtYrh4XzRpXoP/soPSgKe5EJZ
CjvOyPQHXBJlRsWqxsihOLQh61BEd0ta5lvcmmUdR78Ud4wfLLQsmXyBlRYuU7+MiSdL6riUE5kv
o2sCwwVnX3KQE/lLxVVgAHgmvVbLuFTADVrxB6yLEKU1LfToieNU1SNedsEaedifQpZbh3w/0q99
0zIeMQjmJWi80MxPIyirSL88vISF+t3AaKi2Kc9wC4G9vI91v/13qP1BphBhD2AcJERwZPkSzkr/
lLuY/q3Eg/7bo0ragSvJtIzr0L9sAqIwu2ZLDffgIWt1uQHgAx5EZCVuh3oBEOkEkEnHY4VNOtmu
DfzjlxeZrhba7kR/5sSgjfclsI2ZJVWVXmrmD3pN4rjdtxVfZbyksYVEq5seztThfO91GXPtVw+B
UVEwsaGcNblpFTXtb2p/2UCecDPdniRx/y3CDCxnlzVOVPW2+oKoMfbiFylSj6f53aaVnnXDdyj7
/NvH7nJ8BKoCcVxa+HdkSVjpwffWVg2nRfmzSGYXnf/B+HvOEHbSgje5iuRdkN7OrF+u8u8nMObX
6xVEX465pcUQUTUVUu6y4gcp4xhHA1BGd5eaMPYpdNsURFchHBRvl9ElBnjEzJUsx34lvxIRHk8M
8isfs3I639/qIGYAQuVzqHW+Ywkxa+Ta5wUo9AEoc1XdQYPINv7EQGUgpOYDbddKVIFmrvxzK06y
RLkheVZzsfjbJQU7t3stOWnLciSmqBm8ITUALWUtP7tqtGKR4M2rlcnaM7Wc/aK7IhTmo5Mh7vtV
lgDrOHwPL0FHUpzlTjDUL8t6sQyalYhzYPiLB0VapNe7aU9hkXl7e2pKTeqGD2kAZzlojKdNVD2O
QOAXRRjyH5jwu/6Ju4ts8NBdZpdak2cp+BzshtH6sJyd3gg5y4HGwD+LaIT5Dhz249H8s6Co/Ghy
FlW0xGxyyWV3lstPGmQvlihzEOCwil1He9fz+yFeVqkj9HabpW4XJoV7C0ms57FgcjZX5uWSKEuX
Uw5qbXmBS3kwsANB7Sb2SjPdrNvqBVTw2MljYj3qFNa9cORWmk1iPGPOl/QNDlvE+C5vDS22gvn0
C4gdVmh3QMu+rvxnTPME0+2+ATjLvYzMOm000piUi4a/meEGwls42R8bWKiPJ4C47xJZchYCi6fV
DVaeBuGzs40jJM2Dv8/Y7AP5VA2uaa8QLu/TuGQPby8zFJo95NsdX+7Ap2fd8kF55lwJqhrkXsRO
tEc1EXpFCZ3BJvQU/21AHILlCqpFw4wAjuHNDUWt1ckdWdZYYrV92r1e+hcqPwSUBq5uLU9JW07R
pvoCckh6QFC6WIl87zywRweEUDTQgr3RkTbAA1u14lM3NCoIOyuF3N8PCcHcaflBWLmWaDEn2MYU
Jparhzsge5NyiiOZBDWto5K0s3Fo8gYELSnIkpV5Qc6fWxD3oBlJu9mmfgi8CdvqYcCV+AnJqJY/
qV/yMRYAiYg+OipYdJOqwbI/W+Kf2NVaJhGXA5iHRoqSoOGZHWG1HBG1tExWFIMADqr1sOYNDf69
Peal/CCWMEpFbtFwnTIkkwWCtWpzxAooRkUOqfH2kz0MiCucpPDri0uPxwYJz4YuwDMg01So80rr
MVS5QeThfHqPeLu3pHGGA17Z+f/6yPGbfvM71oFIXy258N7IponSlI715cio+JI+he2Yuuo5mxii
anEcWs7J0VlFBVpzawNWu4/nFFXEDH6Z2e8N4wXHeyIvA4xKEHcAkCruGJo3r+9pf9RBkHQ3nVqi
Ktr+S8OEA7MC4EujEISMt0NC+8n0ywq5Om6QTlJzpSW/cyC9w4xSgMhE5X9FYWFKRkLvTAdJ9SAt
qgTrTkqocY7bzDSZRa8gD9gwK88fK4zYqxdhQVea6Nhlchb6AR724ArLn9bQgaW5Xzi44GCOIba2
XYrfc4+93/v4CWj7mzW5Ejy3fFckxrejZvAP9f3kOB0H6klrWNVjd5xcLzbglLbC3hcaFZOobiWf
2NdgyQB5YHmE72xc908WJpmMTN7hVMFY+/f7CZk/4FgjgcBVjtsdoA2cY0DodPe+myiZ+Nr8suXZ
lV37Zz8M1EVrif64rXEhvL59K4iZpClqhRxEFEKV2Dr5vxKosmKvFC4Boc8kZKt9sGmWEr+y3Sci
NLKsmpCoS7Gs506E9/WWvFiYTOyJkqLtXdyoU9hPKZxjBZw/SJy6PPDMSYXz5BQoHSZ+1q2GqemC
8bwomWxCG5F5gcXuxUsLLXrQh3Dy1vsOeQHyt9D8FNXho04B44eR9T25rCDSTx6WYOdY5mgP6QAg
YM6TXcV5U8G4b3gcwldAsOC9O3vCx3K5xNW9DA6cqABg6CLQE7wucdN/ecPTwU8O160iWg1WUKQ5
FLnnfHVnP+OR68oCD3pKYN7fdULBmm3igaxkijBHdCgs/VaeSX1vG4cAFa+Antqz+OqdvyU0ti59
zipoxP1viMmLFZV7SkbytaksBFos+d5um3t17JycbDHIz5HB0iKQQPSjsbmzAxSTj/XEPiVs+ugz
Ez6QdzfNfUu4UwwUqBrvxzi25p+qjL/jHVUwNkb/Y4t7hDzsataHWSnYCfOAlmwN3JGitrbswJ2u
2mwTk38MxmCjMi1dEP8faZHb1se5mOryh72qr5soZscCpW4f5e/XITo0St+jLZEcSBCi/MNHC1GH
vqPgeld5cCm5/mB9b6rnN5pxNTPC0EpsbAT8OK9voxDdl63uUbYk3nEArrsjonXeyAq+u0VlE31r
4k48ikuGFpRjyFc2s7jE1SrJHu93ZXfHUtBVRcFeyF6SmPgHR4Y4+12kDdKttMrioj88qbUrcZqe
P2dx97gE1STVl7u/XIGt/zuDgu+CPsIH3WZifk5YnSdCjWv+aNZBCxHvyiVHRaL6h1k5domir7Mk
9dvcP/qP7auf5PvV4hbKTkSngJg7l7nmDDFchtjuxq4HqPPpYbkRCUhoa7f68RNB04clXfua0KjU
GlkVLpcZvmupZ31hKZpPQ8vn5lKj+UEXu2Q3BHNxjrza2nH8z8WaunNQOAYCkQWf2HuAG1FmU06B
CHSMZc6Jy6KzQnOxXejuOEqOkg+uG5JRS0mqGwFAlQNeotCOmw8+eCyu7hL17GgLrGzXALGIx9bm
AURInRanGq7uoFqys4oXxmPBQ6uyKRBHxpxd3PmfI3a8TUu2ChvrMvShX4L7+WSZkFZmx7CUZkV4
SwLP5eSyKdDmTA28qM+7Sjp3GgHFYsvGYPyZzB4d/gf+llhMZ+EDvMNbtItF5pjCoE97k3Q/Ws+Q
zDkOlpPb3c0N9U66MF1ftz2jFpyL2Sou1XFH1aFILx2NMSKXxCLV+YU6Kva2Yxm4ABpYZ6/+bpLD
JOB+AM83hQd90Mc0aHRmAEBVHvzCVs9dUYLboixKSsMojDMVL1i+5GGKBQ1C1ewq6yYfZAMsUA/I
UqX/fZ9trS0bex6tE/n+itc+Q2ZNWBkUdA1gXR/iHFS4oH7e1y2Nx5wvQN5CF/5cgLX5H+nBieAz
WNc443Mg81HLA5UaRjXdg/jfkZrVYFHC00PS1/sEW7UXp02ufjqYlWBftphfKGqGuyehG0uznXeo
jnfI+iw54yV3wOQOgqo0+/JYzcdWThfZl3+J04Pxn+oAaTTl1UnKWGt8MIEc8gmqXT+BDySuXHz8
iPvuLJqer9ry6D767d8q79oigf41cdcOGmelb0r+eQOtOrmuv3fKtGfxe+pvQhOINnLxf+kCk9uZ
E4LuNz4GcW4MmUmDnFLCorwjnlNy+NGmA4z8/TbOBWLkeNY7WndzjknW3DOSI8rlmFwqb9LvHyxh
Pkks8lyNfmPzsg0rerZHq1yq7qBk+d1WB3EuUnov773lq6N8lwoPguUbPUuWX3MzISKuQ8zDFOrs
bCaMENjhUxetl9seqXuC8rSbcVbCRXsNxFErer0gEavplxfReXvf7odyOF+Hz3BrMUNaDEnQWAO/
7oQdg5VM+LY6mKfo2n5Y9tOKhlEEibSeTpxEKFzAyOE38P6JM1CYE89v2ovFmqZq79mfKmLnM2II
t7cxXCqSKxthPS8NEfSNhUfmmwmh4wR6DJ5JeoYpmwwP7E87s4bzLgzf+TDBqKC/WKJF636C/1kX
SnGeAJ26wPQxp/RiXiWkPMiCrn8WPi5s9KeqJbybVJXjZt6Ly/82fng1uk5bUhw92t524ahnFtbG
FLung1sUWnBdTD2LeqTtYQN/MMkAI7AX5+aVgnP9aL57cNxSX1ve+6t57VYeHAuCeyj5EMF31JNF
x4GU2YVl+5rLQhfcWteLRCSO2KNEbYLxAHTBhTujV0HBtV9PB76gGUKHhXgiXYLlpMRzmo1/3CZC
lh5CCPM04mFOkaj//Jj/4702ZzAZyHRLh+p4oVph03+5eYKCaHXicKk0JXIUyeIbsj0AKSa/q0Bi
otA9wyjz6R3FGCmomG292SQYa4hHCmydaXfTrde9snzjA/A3lYp21Fo68/i1BjDspd/7Fe1dJXVv
QTQA2lRyYCo7lUr1M+1tDa46t3nMB77kvlTapH+lQDpeJiaRUYUOyl6bbSq4c07kapLXtrLIcLRZ
Ddr4ZPtIFOTyPIs+Pbm+NLtpVzza3oD7IPYqAxdQnXa0grNhJ9wexZ8oE7O2tkDKtzeaZaNC1O9+
goiH1AZG0RU3VyuhQLjaAfwAjKKFBsFEBoW3jYTn0pjL6QWH/LlGXY1Fgc2WZSVbwlIs7+sTAC8a
3Pk0kA0zy+ec92lnQiwpMUrXexFoqRZVfZ1XLDmYJ/40NwzcxRfn5EfFNmth8Zb7U03kcyrxWBQc
EwTLWJIjIu0BydW5rA6+qFDghF+G8hv9HdcFyyzNBhOuEmkWfyFuhmw6rB53Z3U/xKKvAsz7cyRW
ugjqwWW8+CLB2oV6XdUK9m6ltxi+0aXgZVA0sBC7yGjNvZsYu19DALwOkSzPImfZ2nhv3HAPggLu
webpvtSaKBQniagQqnGlyX4MVikOC991k+XG7zc/mAYYp75afhDl/qBMW57hgNLSvh76JG/2RjNN
oNq/eHLf3ZjwXP0NrbevbKKiKZX0Ui0kdUstCtrcwkJ9BNypKcl1dRRSWZXaP/cPWqAryV/Hc8bh
k7Ay8NhRlF3V5WGZl5g30z2xacTJ/E7Bl6NFA/EocR/UXvzIwcsi+itJyvqLsW3urHoeLArYrErQ
x9mz2FmUBx4OM8AyZKdMuBLHA001qztGp6Qqb81+nYwnzO7mGykuM4JL2JRu2w6cPNDDKpXxtaHx
icsTp7LqRU7tfwsjEdCj3G/8Klk4tIu2zN/tkJ6vYHw5C4xYTmfcLOku7p8MzhQzkqjMCTHS62Zi
srwZa1B4kD7VxonpE0eX3LnAv2M/xU0497QIeMIrvwzd6Z4EfGvO7nrl3vAj28thj0GJGrauTNVA
G1eXNAtc+ssONYitGdU6r+lJ3i2E7+WM/wLLnUr/WfQzRZzbHErRzk5suX7aOo/DdRlJXOCzHLa6
vgJWAL9j/+pqCsakAhEbP2arHqZr/yIqec1JzmMGvu3qjOaqgQFh7t08K8WBrZLR8B9Jx8QZNW8U
IzmW2VD0y8S9wXaYVQVTh0v4AAYsbKCKvBzKLp4r4XC7yMPcwLteB2orFMssXTpQd19xG3087aUN
GI6vuBNwJGk8hdW/EDdU/Pu/Jzt+mBAGlRBn8g+9jWkNbDFbep5+o8r7M+tJx3MBu+xWWKSpJqnS
3uCdaaIC795NY0yo3wOXmoDKeMWD3lOwB5fzWjGYTFvJt5g9CbcxCbmEjvHXax+/enZy8qJTm2RW
DbqUOzto2DU2xQlIYLgeF99bfrY3VfWZ0ULb6XIKhYOy5BG/5Bq3V9oCUdwIZiYgUko0CzkBxtSF
/cmoW62AvuZufdkYjuOfpuGh8/SuY7fAlN4HCkl8IfzpFakJ+wun7QXKMliuLSGlgsoGZ1YI4dfN
wldO6+jjZe7sGiYBH+28w3glsL91ws8oOKMmIayBf/VRGKq+8BTVAN7fNX2PGzxJlaT1U6R+jfFW
J0anqRo9UkyxUL9YVQ8haAI+RqVUFuPIf7JovuR5pJGa4+yL+UlQkpL1mwGq2r2r3EtsO9iu157R
th7GO37xR69yNTDNOVXv3UEoRABGccrTizfZHjQJJO6GytXMYm+HfJZKG6OmopNCduacXIh2PmyT
aoss1l1/EXh/6kni2SNeBwABboTcluzXYS1ImM+tkH/0d9tDzK8wqgEoQjtbZfJzp1Cp/54OcdEw
iIEzwgb2gf5OfrnRq0NpX9l75eKZ2Rb9L8HdSx+SBHYPi1rhulKZ2bUJfxe9gJE68RlODzLMaFyC
LUjxGPhWRRzTfcCnXcC3CrIyqLf128+9M1bTxjMPz9u4PiRivtKNpOUhFSMT1JpeORHxjWrCUp8T
Z5EMbg3mygCl6nfsJjUEurn3dQY2WnENidtv4aRU4PvSBdWSdtWNLaQAAe80RC0jP+nbs5BSVGQJ
O1qPwhrjOGIfutr5jNRgsPn5xhAMY8RqPyV3Fdk0h3Rr9n7hRSoSs7h+DfGf0BzIQmmmqsnAQ1ZG
73z8B6FvQxCY58qub/k4EjFYSU3R+UUPcjRx0AGTCt/J3L755F+/x0xZOtd0O0awinpx0cQSZfsE
U8FZ8bNPQvhUOLG59PsLMze1t1Rht/NcEM+upPPal4/pB3yekDR/0rNSfSEZl9AgOctkjRBjWjLk
v2bPJ9rcuVHAF+FV7XHcXqgcAhrFLKiBxmQtXGlgEYqOscedATAxJgvBNCVdjFZhsMxmi8bgE2QC
5mRJwvMrowKNHz0tgKCO5+Q4DeHJE+MtnODLnQMOdFvsrQMG2YfCzpwKBL7Cuu9g1VMZiMWRvaZO
t/en0bKYFynGI0qC9UyvXehCXffw1j8EYFDxG7o3erShIFXV69Cw8g7yQ4+cKWzToiJ4q//ZUPSH
ltKpN5V/eKTMnTofWLhqIMV4uVCQui39BlsHpPGbM9yGmGb39Az5UjjQAmEpUzt7im/QzCAF6StN
+i94CJpIfsxftJ9SY8BUUW1kgNFgxCeY8+Bv8D4CquF1Tp73AQXr2TCHoC5Wv4j+YGBW/bOqye7p
ldf5BqolKL6btNtsPNh7HASBCVVKsmUCiKgW7nwlrWhT2ZS5vKtP36WAfUmyOGxEM4eO6d59BfrT
GpCh16WeLf3zJCT0sWwud57yqKK01Reqqerp9x90VFpHg6dWf6iVJfHZR2b7kBMJWLcQreUuqJTk
5aEMnH5u0yRbKDzpAgSb0CI72Yle2LiE5FdB2cVWf8clISN7J0E+WQIByyCzOP+ZpMY8L0s8MGDm
Toq04upltC8mq8ZeR0zVC8wyLRNRWvFo3On3T+JtrBc1fPz8NBNqie8ErCoNK0cFou9sYO40o5mU
yY+k89uo/X7vdFdrL4GUgbY/9GIAXmwbmvgbBabBZ+LLdG9ASjugdUYjW+B7uASUkbaSGF27UXNh
k6sM12tqJeAqlKmpK20vwNxJvtcuXsrSbbmfy/ZqIrc3K8V0o5ZgQJAhJj4B5BeiutAg01+2NrdK
L5mM0+bDzGSQQ5lmvfc+uqyYkqXoeTal3DELCHpxToMy1tJ3L4PBNhjvB/XLGBpDW+GbTiTzWj0b
lGpYmOfE/6mZ1raZqcaQ1ROucDn7SmQgRxxmRx615UXb4UvulxFd7QDvlOIIYnE8JOXdRCMbyP9s
bfCLVN9Dcl1kszhn0cmbWtTkh9P9UaB/TQ4kbJlsV2S5NYiWjKbZ+6t/k80lt/6F773ue0P4JyNx
T4jigwV/VHWOLQvz0o2bDONJHQB8/9EMgzUoPRrESHh67TqnZWVVZN6DDfKllx68Zuu/AV/q7tC1
noVcna1Qoyg9LX/Ix7f7tAYtpuBg7iM6OJoDWj6i3MhDDNB39Ke/a+VqWjLD47E3MwFRDvlsX3hA
uEZnSe5NQGyjo8H3O+pVfrDcHRCYkPik0RClmV/mOr9t+5mrKW5PSa73CVWkn4h4vhGsYj6aiisE
y8sufkk5q6dzNwGJxPghCWBwvDNH0bmMOUWKMUy2dEhKE/kSLO0Esqq8FrtPd46MTZ+ocJfnyG0r
FUGsBHCKwjI+uh22+ip5nS84fe0g7rHkC3O1vRqRm2ttAhISksB8toifi8AR+oGMwNXsF4/v8q/q
IU13vXeJBiQx6h9uEXRM0RKdENa7WL0/bUILgp3FpkHBcfMvGe05rpl4dvpySdPQBV4OqeZbp/w8
0LMhgoK7zAxwRByz8Ef8iz3GB4LnuDjZDp1MYnjaVhquLwIxYPrSw3F6a0VmIa9Mz+8n+DsyS2MD
e6JueoiX5yQhx1hqQH1pbwX1ysMpHHKmLVkzRc632F5/Wp8ISckz+IEiArEyezBhZih8dbVQT59K
5tQbGlUikF/NvIfZkzkgOEs8zlyVFo5HkY5/l3D+tNdIed9duCDRJY/ASIIfxHccZolVLezjykjk
A0XjkK/wM96orRPK8YzuiVD+cZxELct/y8CeSouw3mOhCV3bBuaKe5rRTCIKKPpAQHkRNuAiKnis
k1ZORGqh3sKjSWt3VxHhif19EUqKZIBI1OIjlS0BahakM/nt1605vgJnsR3AIHwM3pO0ur3Ly2Me
OZ3+LPaJ1PIEVsVmXj9OdN0DlmEeEKmYIfPu6dmbUVBaq2b+RwAEWl9ueV6/aYqnb+dmu6QY32Hf
GGb0SqygjtnJXHZqdg7eH6eW8QgOxRezLNfPnpoT7G/mBPC+76UK79DILQeaw50tc1mRvjcotgcL
sCD8k69fnRyxLf4pwaErnF3eN3nugkwKXAeT3CBEoRQRASoOUUfu0NGTDRQ+vXkwclOprWUoeWMD
VkPrEoV74+nwUqaNRFI2YArf6zizzdu7W1KR11N0MQxZ+HWTLpOqwZyKCz87qapJuRB6gfzgPfwg
cNUn9myWGx2bRv7c1Ddc8IGCncXtHl6FpCOSKq9tvqjmd26ZEyYXyS//gSBRSbn4BQ7sPszMzz4c
bRehNKRhObxqEm7rXQDQkQs4Jv6N41yQbie7fVYpcYxTpu2FXMJ9IRpCFbcI8ulXIQj75Nt1qZvl
JwBR4FJv0AQZwi1B7Ox3OmlUiq3jLrJcCB4IR434fwHBXCCrr3pSf/PG1YVKKROxl4XX7m/7lxHk
QjcQu700XyiEZ2k7qGNXnOHNZHBwhZ3CfK6z2XpNihnWFoDuJKUVofqO3FEom6zVXiJmmJe2XziK
o4uW9cODnIdBKeg5SN1155t2b+s0IaZjWqPeciNVDSzFDHeGEivTOR58wfKVSohQ8KwRvl1FA+pv
M8AdQnqkCu2UJats8uF8cg6GwTezYRhj01hlCWlJju+oB/Jz5l7jQkUoGrKs5fJ57HFvWQjp2X2e
8vPs5mF8HU1ESWChMUkMiF6xKGvzWrOBeY1e6ONr5lnMFod0Ha2QbPCNUlU+ETSgiNHX9MsGMmgp
6ieIbLEVG8evy8GhMVb+nr4ijiQE8sRgAI7iUakxaCsLGOUMXT/BauuYQAvVNZZPD+vE5wIsFIsn
5iQRgUOvSTjrw5CoeqJGcUfQtJrZAUvXoMyprxic8mVS5HkN8GsLoInddf6o5eyAAF72D0ImL77m
VOZXiuyDYgfuwqTD3oS7o7WT8wD5R4hvy5rVLhNpabfDWzAqbuRFMN37Ecygkub1gkecQrX1XuaH
pcQlkJKKDh7mfuQ+27g07qTLkgaxsakeSak/DU4HXOnGjjUz8vFeuoYmDXFANmPhHZhb1wxFWeCH
CNdqAhNoh6MpFCaLgExUuFYuGYwxSQ1MUydqtkq8dBZQJCZ99MPjCrF5uV7+aDYTvNV1sZAIOIYz
MvBKJENwT0RSt5zKYH9N1OMnGE3yFfIdLKNo4UVyBtZxP8lp8Efgv2LRsDABAAU3VkS3N+hb94Ll
pok6ARPrmzNRf8MhY+VmYVuRaWGWWJxOBJhXZlqsJcNffOe0zINGM1uVt6WZ1u5l4EOeYL8N1Fk0
32JjCVHfyByjaiNBUp+uNYZYXLWgcDkVWZsT83CuEF0KZmE2VoOE6F1nMIyaC5UefhwAnu78PT5+
ODWZ1Qnsh4lNmmqZNpyoFnSsrY5JwvqD6Stvg1mjvLyWhkVWegn6nMtI4kF1B0lFJfqdY12cFcnE
grUlJIuDACH96dWYMyCmMWwRdKAxwlkgKrbJf8gjllZM4HiVQUuAM4djtG4gPOqxA/SXCtasKB3O
bYUtMNgaVP7CLHQ22qzo9COFSqq0rwoDSX+haTGBiPpIbmSJXu6TzrU470i2YoTGWSCJ79KarDFO
WHOzBwS2PykblW9SpdGJyqk/pyc4Ei3tcMOmf1P2yPPiZeWBh68tlR9pGpZROGK1o7C4f+ZHMccj
tG43mVWtqOPMhS6KL1WHc/6wO6VYmxWlLuftGdVQzbArlgobz3ooOj1/yIthfMvTR4Nnhz6AFa4T
Gf+iYM9F2j/CxSwIoziVg7xcyL+BdkFChIYkjjM15S/PGBZI4QrP7VW0RO6JLwkUg43bu4r7gZsb
skAWhrdw8qiXN/Ud7ElQWB81raeBRY2IfcQ8AlEWhkyBOSuyb21/ShxI5bW/+oz3tnsScmVdjlS5
s72ZjEtbmHlEOAYbmlCoW8tx1gf8lC184B4qxUjHveuT4x7yjeRj3e05vTG96kksHMeJHBxnL9Zg
U3xFb2ADnBxkwQqlqpLltdeQQTkXuqU3v6m08G4QagWLDtmAHcDeWLxA2UyIU00mU955x70u0MDv
v5EYGBzRGr9q3JlarLYTssPJw681psXndBiTKU8zKO+o6+pP0lOu0s0984O7ZqpHEX6EBTGnnlgx
B4T11kg5mObfTTTUXOVw3P2nss7dsVNDEYT+H/BP13n14JmQLXtvBxqZmwPQlZYBBiMfTGFNARxP
612QqkQlZGIHyShkQdf2imvXWIBM638mLHpEsJXG2uz5CF4m/ZYAYjC9ZtOjQUWxPIX7xZ9CXoVg
VHd9K7NdqxZQWR7QQeVDixIMBvdY5Tz2xmsnsBl3fGQ/cK3P1+mYazt7sSsWpXF8W0HyGd0GK0QY
enNHA8YBiSuSt7pFgmv2iu0ujpYwUT/UyoM/CgXFP44tp/4QRt69utHI+KiVhz5IhD3uvjlvevss
ElYOY4xtquT8TQ6raLaQNCyP+ij9iygIxJTDjVQ44Jf4YFX8WlGp7dGXDi0Az8Vxr1AGxzaCQiRK
Pb5j+QOIzUL4szcPfyG4BeB36Pwti9mreVqzbcMge6alGTyo60GFZ3xJzEABuPKlxegVRvQBZjg/
/jlkkgc8mk14b77eOJysu3Oag6QS9iDerpj2p7O/05vfi0+NEfdD8cqk5lFh69+k+ayWve/Do9Ur
sMXXCYFOB1MTURSHMSBzBfaynBc8Moo7hydliXs1SzlzKk1fIhLUscjRTtjdkiArzrqwxoDTICw1
LQSv/l/aa9koOG30vUdyCfMQFdtwJ7ztIjHAfuPx1Kp7RZNJW9t4SyBVvDlHdukKzDjNLppqPJjg
IA+j6Z6YwA/9RQ4wJPKHdXk3VU25K/79F5PhrU4Qbv+cRgtX5H60TCSuKzuUw9oIupEy7bgRDM8F
+t0FPiNwdJkuKTDYmm5jEkdIc4Cghj4hYMMaRMCHmVDazs/o6swUigc0wxs/Cq6g2jj1FIRHvwiG
ivoCC4V37ni3QQze6R8RPJOzPh3XRqUWG0PacsIhHYrD2QmAq8NnMXd5SG8o9CkL0DUxKZjBCpU6
hqS9z+DZC24MwgncET/OBJqaHd0lm2GY5sOAQ2rXt6u2FZHRUlHrpg1GaKQOt1+9Ax96Nvcfbl3E
qg8O6hkrGkGA+Jr6kf8+6SjFcTtXfr1pVR8bR/D8+wZQ7/RGLb5jcoMTL+q76kiawAI7AKoe7mnN
RsnoFmlMgnH7FIOSheITCimIfBBdYYqSVGI5KPFTp1nWsmEzvLc+elrjKRND0GFpOPue1hL/6pqH
sU9tNXQ6aAPl6hDsflaQOg7XIywJOUWB2oeOi9EoBIPOjRDEx152SESAAyp9s5tf65ss+rVvQZKN
pjwtBDSLzezFS6RJREtgDY1pj2dCB8uWyPpJj1tsRl1CX0SryyhlS7tMFBdIXHfbwyDzk9sEYckl
fkKU8Hg4Wn3Q/d753Bwl0j8qMkybQJeyC0gmiRRcbKEiSKywWvggWoklPrh96aLbgkZx0qq+OJHN
0QRh5z4n7AGgcP3mjUXmgxEtM3yxojYxtiNBxVatFrb3jTEHdvERFL8u6Ms3dSCJALi02ALjHIsA
0g1/UOL116gJng/zci3sqjnKLabl0sgseJssOsJo6R2bK8HEMR32rHZeCiEx+/1fg1a5rFN9Zu/D
T0+u97rws4XKNB7bbPXCLLgT+trMrnB8J6xZ82BcT0vBRCwbwtMFW6kDkj1OUaZur4twclOF6enh
xdRgW1fd7oHSG19Mn487xI+d/+0EYsFGT+5o6vlVFWq22zK+89kAM7J7gSrnkhlSiBzWXX195NRu
UUy4WCuo7H6AgDX34eLc8Dm77Feu0yebstvec+NsAAMMn/p0YL78kCk7H0d2fJpBTA5R4o14/Mem
aaeR+H8OllxDsC3qR/w1lCvUT7Kjd3iqNVhHC5v3R3oPFcK8EcETVVoYqMJdGdKMncxguvwB0uLT
1HMQgwhP6FO3IoZ8v+1dX0U9JSEwBSLgdSVxGPfFD2ksq4H8S8U7UXspmmzgOVNKi6Yys9Tnhh8H
Gcp2iNNirnE563xrldXUHO4OONzBLs2obdjSGHMoqJkkDdIALwIOP0FiFkLbdAvKnu73yK8gcGaG
nOJAb4iTIJbeFEQm3cL5AKaOFmFsFKV1WObfJvxIW8ZEgGscVWecs7of5KGBJJKXjbppOoR5pc7N
JOhUWtFFbe67K8PqrmClStVYyG37+3pNJd49CixzhMCJnWqQBXfU0NlZ3wPDPzOemFpHmjDMtLpT
+VL+cCy/t7kavmdYFVbs6G2ph5SP1k8/NtfzlupU0ZsLrDFHX60UL122u2R9xoTuytkLdYz2KycJ
M/WlGHAdSXDrPW7t3E3BImimGzv5RGjIcJlfwyh0LnnGI6lXFrO6wokH2TxSd9fGQZKEe6iALVg1
J4pr2v2td90v35xpS0t8Tfao4Bl9obwe1SArah6DnPX4J3vFpmDn/t3AYFW84dnbRyeCM//gLvjJ
N6CIL2ZNHjrowezzbfz5oo6Df1jaYtBQQONpiQuR3RItyuVqoma7yk4dLJJY6p4M7q6oYW9MuoGw
fSV1b+qww8/9SYWxXym7piVAwJRbzlt5o7BmTGuSNmOkWrJLPvp5qt42qcA2jzCFhlfmokM9XmBn
OQwHZjpgQ0rX0t2zO3olVam5nQpBniN90DS2ghUiTXxGcHI24Gc1zNDtJ791NpwYT0cxf2NYmfG7
6q47u03Idmg/jaAU3ntVmI/yyja8npDU06PtqYtP0l2UYemTDdeVDvIelz5yaye5ZmhbV41wcO1o
IJa/CvqkP+G9f6CSuUSQ3Y0M8yn2JV+JeCr4WwI+e5CJooKa7fxOCGY7At7x1Kh4kIpse3Z6Xxql
GfmrQPYTn4fBQF8RrvkGhaIrov32SRefv/VVTTSAqRyYFy4m9iRZvF3o7iPlP8c0lxe0MBX4e9EH
AGhF8iZ6eE+pQ8hUzut7y15i+5+OV/V3bjg/IBstrpTopoS9Vmn9iby9d3lN6RyQ8qazGv5c/qHX
N9HztnrrJyD0P2tMsJjS9LW8kX7D2SnT8gDYFmj9yq/C5eOsCTlgqtGX176INzXnoLtw0ZnX0omp
DO1G5T+ZqYT4PR/XZap0w0Py+qNO4KIA/3twcV5WMgkCh9yRhb+CSTPIMtqRMKgETrFQ1ymLpPVb
WJZBl2n4ZU3yD1qxXPVqVfy2t7j6zmTWYu5Y5EyQzKI3tBEALohEAGzitT+0IVQjkmE3zHsKPWLc
jVAdBW9p+Ge/sciI29yl39ABPxi4MGBMqaF5pzhP9SfMoqGJvVKM1b9cHiweomfkJtA/o/DU9HCN
Vg7qMkvdZW99wzCqFhg2c5YU/Cb/tah3T4nvFY/HLOchFun86QmNjbHOJuM8sXA+quGKsp3Pcpp0
QN6aWPBuBQNv/b3wbcxWoBefOgWGf0tSYsUG+oxVojjlrCH53lM3U/N50h1Jnf+z/y/leRm8nYP0
MzyI7f7A5gajYDlKmC1uSYGwHoPtl8G+X24UAhBhfe1dyyoK+tEWqSSeXbcFsVGeZmT2kScryDpu
czwPK/S5ZvZ5zp19b1CHJekEWrdzDtC0jft8auGzTpsgQ5Bp5MSQjUIFlFoehjnI4Qcfzx70BXfF
JrKNxOWAVeeZnHa/qJ8MxMrPOpZdGS5ot4jHPa7L1fpCKeaUxFaaqZvaI+LLqZOfRnh9fkdHVaBI
BjYSU3CJ/1wrsH8WmGQK9t0x+x6vI4CrgG1Tkb9ja1o2LOkXxMoG1z/8Y8FPGuzaoEH7I9rsJWv0
YYf9zEtAIJ+0iDkR8dTEyYUZzVy3Nl6Mq6eMUfEEBprS1vG45TETVHiqb5vi6GlyGKqb+rWehv8P
8JD4XIRNSwbAg/4+FHMD2NUcFgUwr6xBZt1p7AwWmk1E5oKVGTpp9MlaqLrb6W/7PYAyv2uJE1zm
TFOJMpaED9bGD3P9esOLRSar5C5Avr7MS+rfhDJvdTnMALU/Uhjg+LFIkMLcsBAg0rlISxqUNaHW
1dquMi8fdy/T1z2XEe/9H2kkGPinTMnc+93tVQSjv+fmwALgKFX2+nQNUg3pLTAQSWalzjL1zz56
79FhNTnoMOgk9lkTIzE3dacwzXSSHjzjMv1xHb12x4mNu10NVLvH+1uBol8Pr+k4EmfUWopkX1hy
rhcAb1ZS2j2t+deRrnMSn84x3k76tT+AXkZmhyDcCaxe8PKLLN4cVvvnV3RH65JUPMAOWFpntYlO
vTz5DvXSja2A8XsFsBW7QhYddTdWtj/7yq2g2dPfx9WBfLtXxq95kTsCvemaW0wlFqtq0vx+V4o+
o5F+jl5UAME/+fdysEK4DY1/UnceD1vOmSemBvi+lB0Cg48bo+RMrgDQaj42jzs5Zf95fPs8S946
JI0+NZ/iip0P4zHTf/EsgI8COHhtKH9PvqbHEI+qAroH/Iy9hwob4D7RrWy49A+zImiEG+7+9bHB
+G7A6ra6N//7hobf09fGwDyvXO98Rd6cmRqm+M8z43j5t6u9dcO4Fc/Wl3svsKxZOl6NW8G3nQ3h
CvYp9UUUXxakMLKEl3buJNAniHm42y8jnXkazJo/wpRywfAUcZWKzXObdJTmXc3ZdvpPffkJdrlC
YY0D331z52+Yx01npYvXNqOyWbgWh80vRsSnEh9ZNjwaEtu5DG7kwOKquGog8ggQ+uvGLiAcpEnA
ik43D0w9aFKSkJSRjPsknM8vAjUKM4yL9ks8mKclHCcvu5Eg8HwLup9o+Iu/vUGZ68PRSFHPTZbq
5VA5wb2ek1nQe8NvDdcs2V8D4lL3/nghshWeiqHBXJ2pkTQqxLuvjfUjXq105EgOiT+xXqeyHQbf
sns4amqGF1C8Yj+Um7KMur0pH40n48p2eYnpmIFRFfv0m2WFZ3KpsPoiynL0xT6widYkYoGRTZih
3dOs9HhRV4y3US83gTeduDoiRKA8VpAd97GFS6+Co98nVO7CJ1bZ2RpxOSBgOxHfgPIR4tuAfEsY
wHug70gZwZc2cPHnrByVhxmvPROV4ZRmoKkE9mcWavZ3kvRa2ytAJXSpYbw0113/M/gUcRgrrX6j
c3KlPNkVVgsNpNb4cAfhaspnrugSbMaOdgnhE5UB8zNBi0jDvA+5/yCL9kDseVXTyPJBsC7z8+Xp
kQEtsXc2jPf2J9J5gcplsPE+vRyRvbycfMkl5rpOAOzKxPrLZ4Q4U+fvUJ1y/iCiyNRL1forcwFE
Vs5/PkwRkJJLvBU8Q7KQjV4dmKO5Lzym36Ej7kWq+JirsPF89Q84r7qyxdFb6wCQjSrEJFnGcgZe
81usbN2fPuS1TgOMJK3XXVXWhBg1zObgC9a3Stu31Ec1pz+6RnkNL4k58fFhaX8et3uw84mcaz2b
5JFx1uvGLIrNEy5I6YBvLpJOTZgkHNBtP00vOsg5DZWbyn0jS2OB68TKHSPMz1cezZoPAhJepEJJ
3LfDkJIrY33hHmIZ4Vn5JMrYZeaFeRXCoJfk9B/8KaUmyvp6xy+qjKASfi2fRx3An8Cc0hGb9Io4
d3Tj0FQmRWyEugx0dHpJSBXtBQc8WT0QRKqBbEETttlc05CyH2u8GSf7oabzqJRI+B6nLNhYf2wp
NuWizqR+cSC4QBumYxhNnfdtRW/9Jk++5/96VL1zdJoRYFH2F0dGlDQXUKDX6fYs5yXebxO3HbUn
tBT6KFhVstXHkY60vU5Bn8ouj0FOAa7/YHes3UeOOz+x2IH4c8niiPGN6btlslRxIzrv1IICr7Vn
yt7FBAUz4FAcQHtC+sfvxIU7dc8asW6gGItkYSSi8fP7fi45oJA/nriFLT5+xc2gRCTuez9y0/N4
CfXrn2SVe3r7aF+RTxNAo7d/YF+Rdofet/WSr201m30xcGRMXx4aPeCpQETLB8uI1K8z0+SplKRY
qPRfNFOSfdVDbi3oLZthDT9s2Ji3Y47XsgdPBiu4z6Z+a80yMipkTGEhv01RJMDKNF9MmEcwXJ9g
E0ucCfDI4kOfcvplCgrMRwUwIDvRm0tJJXq+wWtqAiSLMgoQf6msH3bjxGWN+W4lYC3xGoj9Miah
xuk4ZhIfp8CalwMoaswHhSomoZDj9bBZkJTPxZz/XP+AEEXrf7Xi7HLTH8NitwXMMj/RkqzdX4GT
ECYuVl2AV/Sulq91M3H5lapTnh/KaxvOm0hCw9OPxLXmEnHXypkLMAzAVCEPqX69VuH9rwwwz88w
K7vmDqz7muCWcnULjEWenG6ryBJ79VDdE2HIMHyGHAjwtTVZa4MCSQGWE2AZivvfB8OOmvN5YrXC
wRBEgRRgVhnFOYtiMq5QV2lH0/tGcUsxKQX5BcTBexFurgfEjqlbRCKuR6iaAkT3qnjFcoBje/GV
hg4edApvxsKI2gz9QiMeggmqVUISBOKwr5JLg75qD4mkQRS6oHUn2ml3F8vW1+nl5g20vdMDi0T6
fA/KA+w5bAon7WL73kGPlT1AxfBhvBSv84OluRSm4qKb1D+l84ea+3SHC7fBHbtpiBoCha6XxwaD
gdXVg5JWCsYsB/6Zf5PZSqGtWVn3Q2qPKxwjsElFWTlpYp4r1oJeZ4L2KxIu8EPhF6iFNAPRnF1o
tQa+nd75EiRtkaWTygPZcphO+5Xx1QfqQ7C9XcF/M2KWy4Shkty4NMnyQP3UDjW56nFtyNHB/Uv3
GcCM5UGVbeK4Mb8hJpX/AxIyLMGIBwFcLxUB1u1LqE6mT6wQvmiSk0cnzerzUJdau48Mq03iI2EF
QeyBz+6GATf8gQdNn//xyhplVRKxOWrZKt1alaD0n+R3Shrzo52tuWLwfWzGx8LAP4VZz1OSaOYm
LlyoYlAuJB5gfR2rKcZvYvfYsylqE4Qd4ugXjr3fU+yXw0GFG5V44UPGsaeNmodlYvheSJtUGKW0
eMajs+HZqz33kSIrbX1WyTTkQMfzqbfTMOl9sLU/U0RfZiqU2e738kykqb7UqKeRyuRVA3GpvGrF
DrkQ9ehBiJcOH7mTnPy2GnXIvNcq6VuXSoU9u7wF9wfyBwa4T/uIxIszgVBovYvHkPTtHbE431dT
VXGypauaJdw4cXOPUAdivtFWjxiuzICqGMe/jcP/9I3nEYDFOvVmqFg72hHHVzJn2G2/2+aGcVc5
qRKHfT/T3OYFrCiZfJ+mdCIVZ+uDuCsEPhtw+vmgrX8oOHt9/9F37c9lyUmMI8MT4qs7YB0zu4Wa
pR76qai7Ia3HdUGfw7VpUz/w2PJVSccN10vZyw5Gkbpe+//gZer03z5SH7B+RpYCmM8o1rz7jXug
3BvP5N8ZC1TLXikzSIv/ookUdYc85HlU6U1XLfqAQnUHRqqolPxpn2/5KZxOmq9dnudD15Sx6Ssq
E/6z59Eqh0ual7YJnUL1vzFOGdwSe1epP+fxA3MH+c1jH1xprS+rGgfIHxePQIsC7OxjcRMVwv1y
mCIpxQL7/g7gZl/43bNpxj4KSfpFzRWG7KwucICPER8YdAxcWgDHO3b7Ts4X9iaiunadPmo1DWrS
4JbHFB+YjM8WwG3qZGpWAn92YqZCN1mSvfPrIA9CY/M1yiser2eV3xLW+D0o+rye1QFAK94JKeBb
NR3ShFgoISRTPVuUFkWVZ+Eb/gTs9W6pjJ/Gh312ysmRgkdcaARnaGYJaB1esi2v+UYNm4s6X4g+
VNZhVUyVBzVairGzxGnfCkkkxatH3gnIYDan20Wmr9BXGjsk3oMcCvqrPsVT4Qf1EiqeQS9PCsWQ
Kk/zmN78L3yu/TJnTH6vPMTVZeJ4ocesNHaikRkQ5cBH1AIkwZTLDceKCPjfiS7VgoQ/c0ZbmHJ0
Yl+80cDzk2KOcYLYYYdKNNY4OG48mnWCn+RTOJyr/11219YUDCi9vgqawahAVvxRdsiCglCPioGf
xxSIrTYembR1fTOnylASR4LshCQ87RLmDH1reT+1E1J8QRW1yZpIj1iyhzxx3vRey2uwYCR6czUI
UIucbdxjrn/S4bes0AEdtMvyZy6TNq42fgXw98+byskTEd4ekspqEhoXomyZ+gGo1gIzMNJP4kWq
0pA4876lGz6e03Q90nIMQe8bjgKOKe24kC6cYzxt9PzlMY3szFo3jy7gr3Hz2tbEEbzRsjfpxLtn
Nn1zzjc3Jze+mpqbpC5sTNMxNRfITLmOpoGQ9HG8mmqiJg8W+50bn0TgKSy/wssHNWxrVRsOY6Sw
AacK0JQ4fEKWPtmYY+FzM8dQJqCwM5amEh3dM0gn4qf3XVCzP90AaG3pHpeR4L5zOsIqFLlJMhtl
OYdUt5cQhtMghhOEk5b5r+GmZ/qi5uUN9hyNY1oCXajROKNh9W0/U42I3iov+dVULuAHd/BSRSaW
LoLVwCdh2xrK3fDN7Y4XErAnhjIaIUH4uq9GSKOrdv1nn3no4FBNDmQgWawnRQ5u3hFgG21p9UYT
1KYxCL1CZVldmhTtWiQQ+1rKll57A+6WXLULEcjhKLtZDawPkCAAo4DmSaTkIFhzSZaSai/cJ0oq
wosCmJtUfDEOuOMhnEuBwQrd+rgeC2itj4Nyb2pkWePlKhFjy4J44StFlrUXJmt0Qp8ne1oEdNkX
4gfRRty3TmqeyL+bnBUz6MD9wcVRAA4dgDa94Hf7AJ97pnH1clutr08oXw593ilizdKPQpTWVt73
U6yPDgTa6fU8lkdqnXHRtpgpSoyzyV8bgvtMBZ4iNwX8g3CTj+ZhjvQXIEZCR6KOkUBjemNOpaYd
TInqR2ZxOKb3WyED5KP+TWv4cpksTVowZPCcKqiywHT5bXt+yiIbm6Pmqz/LA4b8clicw+0d7ep0
f1uHisFIcwJK+X+5ycJt2L33R8A4OXMT2S+ch/tel1HuRPvwrsoJQPywuH1Ivdi6RHv4Q3XbzqBr
pkpVXy0eETtUqyhvUqCqHZhTxtVgNeXI0aCnlozmLS9T0HC/NeQ8WbblXXe0L81Y9HPS1JoM+F8l
AJ3PvkBGiFIBdNU4ISsaXXeocY3HrmK5AjWavniyh9wcjKr+yg61QjvHA4PsrZbSh6vR6LrrHanq
rH0J9m9PzpQTh6mRXxTlrjkk0Ab+CjFFm8NFBldbrCY7dnQ+YuoG1gHSfVdzkib4wReMF/lRNv8e
yGe3nTd/dRKmwGp4UtKPUecsYxo6f0L8FrAEDcou5cUvCQqLmVTf/ewCjoikC+LfDjVca7wbfsVn
biT8n6r51abqjPMPBHsyOW3UCQoo0LD+uzPsVh7b5KrMtqboKJxCj150350CzkLjlea1h7bmsRcf
oNcerbMWANy16DaVbri4EvgOvFYSOh0B0457/YrwNYzcljhL2Lgs9cBtz8xCscOr8FPgZhGk14dh
74f9sqOki2uCl9iaNhDI3UxvcSlRyqLJ4uGVH6qPhbKuWB/qXG3/aVXcyAT28MSfR+p73An+u6YR
6R3wrhg8KykCxsZDNBzfPs71i2QDscbZW+mNXtTgGT8aLf0Q46Z4zunl5baFxHiiKYXRMoh/I9GI
3UI413bILXB/TJ3plIztl3HdxhH4mLooNkvR/AF9G8eAcoS82OolzGRFO6YzrhHTZRlVFqRLxnQA
8uFfFxUzbGPNCaTEydOIV+Pu95Y4HkIHMvo7RxdZN6HPL9LNNV8pV4k/FLHWsg6MC3QKYMIfRk5S
bX5vQIFTXk7ZY6Cct5PYu+9omLmkKn/79tpfNTI5pbZIKedaTzgiTr1ImSy66ZRKvs0txj0qa3ZR
D11laUJVfSRc0meGnZI46WNBYdm+eAV5N94jnN5Uo9OtnmkTaOfYosAEiqSxqDMd32vFt0k/1oRV
TAkwz5jVgEuO3y0RYQc45VofQToAgCjpI7FRB6TYFX9P7DOw1CWjpwzIgjePRcuvSPuITUSUEsxc
GfoszWQ2Kxb8n5LcMioAfVnzOtSD6mm7mwWb3myfAQLG2vGD5diIE/2Tnoem0tmJWbHDVavtG0y8
EXPA6Oj5ZlTpKXqcbHYxR4CCrvSHCbG2+lIe0g9LM9Twv7uYqaSOeIii/d/Fy3P5VKMDTeOntZ0O
S3h71P6Qqgh9AcMRJPsmzgHxZXtki76lu9dQhB9e5s0j6v/haIl28gtkzTJqXEhOQhzLI2zMBlrI
CkVEJGt8T9RIpb+9Qkr0KpkyZoxtiqhVYNyhppMbxMBChHj5IJp5QyHktLvpvdPdkhY8w8+4rTRY
dPLWj+r1WBMpj+B9XQkin7+3PA38vCVII/cBL02E0BVp5kcqxKnzV2GLdIZalw0bekLmUrJ4qk0v
LF7oh7eTJorhJZF1PzVoVq2kCc59SjA4B4QKxrobtkKT5luPkYkUcIjO6g+CjTr8rcvcfB0wHLGu
bstDEiw3KMU5ZqELYCMhALb/byXFJ8Fnf0eg1aGwg9qulIytBVzTvednbB6E2tXfhWD+KT3R7Eb/
+sTszP4v+KpiBY8cXBrQ/VgN6nC8wupmJcMHubDC03JiWy4tZDNABsWpn1Y64vPkZWn04esMOz+4
yyTSw15dLjE60NtOKRbXYovChZli8i5qXCIeq+fxNyXP3OhvdCbVF2FPLq7n74ssNF5ltWJmBxgJ
mrAuM/4JCnqNd4e2ZHG6fFYJBQiqYuFf3jNpLZEcVy0/p9yzwLrBb0pQPhfR3fi7H3H4de5a2Rio
V0oNoGabm8+bzh9BugXWRw9wvwwuTxZ3TF9uzPyYfBtDrLGx4pwTABHdjS9gs/akCczJ7hxmkQEj
kqpas64jzvINagy5DPcvRWO1NB1sPvoO+kwBuot3WJGO2eQgaWKfyse7EBZFxUXJ/BTDnCYTj2AU
H+I0qdWUCe0mW1Sbb+/69zp9WgpjKzp8oBbKmRQYgFQkWf9i9o0VRzbroh76qGaEUYCnnvJe+1Xq
LdVi6peBEzBBtotEz+pRyf2TkhbRqMTRqPD8XeaaXUYB8LbNjH4aUjxlB1wlCLOIwQFP/MMwAY/R
WIcPDRD1YQDO12LJF8td8TUPuj064THfmkYWENeiK14kqLnq2aF8gm8fjFoIggtyHKRn7XJDhbEA
2hVs4w90+3u+Yak547ySJ9BJ2cdgam4+40ax7k0rVaE2oaoJn9OIG5Pn7YwfF/6d7CFjh6DWLU3l
Tg6ZZuGGFVDnsQ8zlCVZ/wq9Zyg1n/GLVODtxsDrTYg/JIs9e6clBcO8SkJ1u2n2Q1+Mrj5Jmfcf
Ai5K+j2NexmosI+C2Y4/kpMQIZ3HSEBWMASW/tHJn6qrHRY42zRLi7tXV/APa/ADzNhUODo1Detl
Z9lJ7Cga19ZdfxeZjE4O8SiBinIhnD/7v8bhWkP0xu6km3enRJCQGxtneGgm3INJK+CSc1jCd0dU
2niOzbf2uhM4PTJUitCyoZCfUL5k3cdKdLkewG7zYELL2gfLycvwFVEbxHMfmxMQu/vQbhP5kCSw
L22C+foJyjq3Fp4+442FKKZzgpgczmRsV4+8igpSqQmT+s6lUkAayJou+PgOPN+5Y69eWgKJ6abE
ZnvH9jKnLMrZKQpEgA055F5bMvF2RAO6QD446UT8/83NngmYL13c9pozsSPh4nZH3hVDckt482fj
Mr3UWTTvl/YJe7oaqIvGJFwe1sRkNid4Znyf9x+2PFL9XUnm4hmCUCF31L7Xf+u2umjSnk2alCfB
q3RL6fZSMbRjjZENVTrCGWTm6Ax+R9Iyf+XnxQ1dwaBrcJ75dg5zM0fEqDoinBAUtO6ZaRMe5Z5G
e/OLQBBkq4pWnJjqo0vUYf+Mlav23PLXmjrNlRM4aUU+Xx+6jRgBLCk2YtuRxixETggrOhqYP1BS
UBJOgCPMccC/hC3IoqrIi4xQdxzrAdnauocvYHOr8A1Zio2Vc1/AEbL72X3YXb4LpAAddYTy6RQ+
JkLR7biGjVyIX7YYIq7lmk5wEFT40/K5i1t9/Cc6qoqt6jXHbn6qSH2/0zCD+UDLjyD2E+7PHUfV
52SRmrZBkXHHqQDVXLt+afm9PlEuRZgY+g1wFfbKoCnvhBonJ+RSMmrm/201RXr/4PQ7c3Q2dste
t2c5XVKQGeU8BFsQ2MRhatZDUUL956Ob/F4QVt1GBJhqS1Xo3iEGlG4YefI0XYyG45eRprFCfY9s
wY6NlkeqgkemSehVP2xUzfpGcculhjKrMsGwgBt3MqNtGciLmkz6jH+XNJm7XEA80oSUgdoSvTw+
7Wtu08X5J3KzoFfULa6hoJ/ptCegunqPW7Tq7IvDucA/Y6MukzSX1y8JEdbVUxSjZRCx0xMBB30A
lE/3F0wkM//swF2riKhPz6cd41FvILIQZyrNcKqKVmhEv4eZoiy2uR9VS5MEdbIMv0+JPS7+VngW
iRbgIAk+yPpEXgRO7s7XaRHmfh9YUm+xFbwy14VPDkFRbwIa8WpxyTbkMlJlLMf6dlmpuHvQu0pL
2vC7JCfHWCPFYRJl2iy7UvNlPGCStxaxTJgzw3E9cXaofANBWq6oVgN0zyjawd4Exi0T0LDEaIkt
h8yQEIBE82VNTz7gLPm656fzTG8pk4BpShZI845H13znUBGp6+2OGm+mE8U0CyT6Gsokxct4DpjK
jrvRjf9Gjeg+Y+jLOppup6lYGUsAUUkUd9oPyYlpyF5GcaFrleZ6jQOE8WS1Ubp/CH9JZzcJFp4J
uhuVpzpnmUAzL9tdeZ0XH5M8FOf6PjUdzhHbnk5oszR0ZgS/ActHKL3ZXFkzUCMPUREOthPCMJx4
tGMl0tNtlkBcriGxAnpuJwVipNRPq9Dp7Cu9RaQa+CnaLKy09shwytrim9WT35p3hgjmiWGvymSH
8SCSA2DYN6+tw9h7AWtP5KQripqT43QDEzGZsXpRcFIqo6GnFoEtujk/gGmIxWk2cI6IpmToBTEY
7BsFEYHFGAL1FRAh/0ASuuw6POEtGudihh4Jhm1bt72rkTCezpenSyMpUixlo7+5hzUmF9yO2ZmB
b3VE+S4Qs/HrI7rEYRgqKIXeuJ06gwDHu0jF0DDIzmhuHpDkfxLxziQKPtMnXSuXSPp6D3nzzxKX
hLG0q1TaAW/lhEB3xoz6GvrMABElNrbF0eUsma3e7VqvpREogixvRDV6onGhxTPN13dyvYGCIRm7
QWEZGmM2nAbK/kyRjLl9LeVFfPEWM4Sdga0sc6Rw5YwVXOaH0e3DPvjie/DP4mf3ZPxWhD5CetCJ
kyD/irBCBFAHHFBlpDc4ooBwQ+6a2bL6TLTK7hHkfyEWoRVfO5qUaa813vjd6SB1SE0CHA0YPsB8
H7mK9esLWxBHEY3aH/DINncKHs2SAvjAcFS2RP6WA+dZ21IpnVDJOeBXdXT0AEuCQrDg+1VMrNy4
zxc2k2cDBUObzh7irskvtl2Hh7uNY36c7HWLq4DgVBTqUlBy4cPBvbStiBWNIVSoynDmdZH0HIhA
h0h5zwUCP+Ps9fdN8UjRywSkRqF3PO5g7gwBHWNnJB7qQdee8skzNitwJFt4VC6zT+UvbzAJjtlA
T3SH17z/+hIIv+wImk7as0ogJ+Epifz+MgUy9kPni9a1+C7BNLi8SF4ukBIiYnwRNNfNxv/psznX
DaLagVIRszmcov314H7lHau0FYSGxW51d+0pqK2Xoc21xl5FlRRd3M+jrFAbxL+h44a8cFDGBhBd
QqAMKnUA4eN2fgR6sNYvBDV7jc1wn/nWgFyksrna3Oruq68J1ufjrCAV+LkGCYY8qmHX1UZIXPMo
Vx++JSLp49oebtI+vTMrPnjIe4II4iy2hXpkXA26cfWR0QPh+gJxrWqlpvIXbNbZZVZxicq4DeR1
/FhdxwWeLmDXc8JxG9oJGbQH6e38luwgEpLbISoPl/sP4llYTzAVZO55SrS2dDXgqccmmezvIh5L
u/OhQGmpVanb7TuFQH9lbuU7pSyywx2ZtJyY7Vy9aLzfCLGZG3HXwzfaRDnwqMV/vW2lB/3C2HEq
E3cNms0xn1B5i3IYesvNDvBTsSnGU0+mn1G6xYOvoquQkJtX8xDBLwOb6cZTz9SX/+Yhu1p6PKeX
ZsvrYB4AKG0Y+WvkIp2TyRWvcGU5DrA5abvOEdi/360RI+p8Fgk+XUt+WRPvhrjncNnDsGFBRv/d
fxqiuAg2LHLNRbjI/TZgcksIpKaWTzJZdvNhwIWvw/Drf37YyfWAKKMzXpaGuGzaF0SI7hMd5yE3
Whi1R4oI1ACT19TrCt/xZeSyca85FeaU/axCPaExi70u0QtqNx5Ihb/VNK60CFho5pP5uApN7TlB
bYuJv1DjFwkN+C7AWxFrcTp2JD2kIH4488nbE+MiheDhnQzbnpXSDOULIH+nJ80r3XwBKWgQc1Hv
Iefqlt3CcK/A3oNlhkV86dcy27gFu9d419x3o/6Cm0n8mp994nnBgAirELyoCh25FrlnCFkBqmOM
H0ceWBNYH+6BsMsbj5+flrKaugmwLEoiFUjCb91/AJBB0t6VLv6s6S2q2nx/eMH3voQXcPON3Ih+
qq7pyk6yKzqCoRw5L4tmIm1Q5oDJQkFQDV4tvt9X1syBe9bzSwlLXErHczc+IUMpF92yFwcMa1pW
LI9iEBAOmRprDMvkXyNJbcJdMi0y2WURSC2gco+jKybVBTAXy9lcaZZzITFqxKaCtZK5+le0eg4v
CAve8Q5vhWQunxLeE7MiTDiXZyYZfEK6DyJfWZrVeovNw95ZvxWDXsYsG+v2VL4WPohlCpqc2lLp
7aczyb19OfRue71T/KErmGIwwfAITdujbMQ7Ribu97ExR9gT2csvdI1Zp4B3ypW/m0gnsbb0wesM
Jtm44JdryIqRDnzWFwh5kLNUx8RiTlBWf6WTm6LVYCMcwyGtxCY6fk62ZdISrPocIwT6/8K1QH7l
tohjdqASjPwP6Kt/ik6jbmTCx4BgEic2TIj8gl5qyRZPhippDLkUDi7aHVrvWL5ISoA/ZHr8c0Pb
pycLlRY8XiFXjskKr3MoiEgIP5Up1nlmm2Qic9xgtveyQoPft9GOTD//P1HDFPa2fsSE4CXOgF/J
iq8Dqh25jqZEC6OzYmCfKPjdBWZC//t0+fddFF63ujzB1kYsMmrIpxMpStNzO0TGt3NpJOvE46m0
5lH5Y/8jG4A4GAqVk5SgDUSMtyfCCaLrcZopmu0N0fHNncWmkXyArid/9kHVyH93SfZA2Tz/feKF
afVB4XyF99OCSH60yHWPGoU8NcCOoUY2kvWeGapApOogb5wuqYUf0vlkZzH7DjDW3gc/wOiDeKbz
UkXArra4+V/rFelbTn7xXtM5kpq59Zsfr/fLg2TolUgs6CdPIGCosCoFwj01CWE1lBC+lG9Zv3ue
DPqLOqqGgpxfjbYSN4Rscbb/JTapwPaCQpxJ/fRWSiDL6XfJsGhzrm9kPMCPmSkLmLIbDW/aM/FG
mxTrlvc7sY7Fe4wnrDFznE2H5uTbJlzNchTemYK3ulYFpPvFscn7z+CIJ4SCzHZGV7M7Ig7/HxoD
0gjeUeY9LzR6ykL7ZX3roF1e0dASzDrApns/SNTTjigZPeT5xbsrrBNuH1kIft8AwUe7zl/BOg+o
qRYJbH3p8hO/HOze6SMeRo0GFvs2Xw4oy73CMmh6cvwG8iz/9WVT9k19fdwuzv4wmgq67ZkhV2/e
sOvc3M5/h3P+prwchiHkdhcue8uSm7tjNctYVZ6aTbUcFrMQSks1OgIil+8yi7PHPT6ZSxeNz0PM
cgvW6+aSKhnpFUTvprKgdAbVTQIMCRorH1FEPL5cvWSY94F/LxyVbBDnP7+85154UXHXv9AgC1P7
flX6qYwHJtmfbOhfnNceEHQWaKXxJmFGC31Z0wzcfuhJUtsJVtriwCs9n0HjAGDek1aCEzYUfG5n
lqw7XkZqF/eXKscxYPh1QDK/1VIstHKGPiQAUk+IcLlllzG0K3C4CEUW8J8ABLzgokZK4DtW1yV6
Rbqiyi3o5UPKZKru4kO8ifyaFJP3Yt22PDUfRatQPDEuQcJ4elLJaY0ZPJBs+fbN4OB8Ipos8JAz
MD8fXPpqdpvXtKLG0ajUGQMPWq1l1oL+WbonjDVISjU/hVExKBdryIoz2wDdiG2Z9/pk9li2eXwZ
rF8Lfxep0rWyFno56oM9J3OeksrQM4eHhSgeX//VNcP6PBpXQiDKWS92iF0mUZkiUxhZ0nVnC+u9
3egStOqyT6Z+r28KMkns3BGO1mX6P/n89zrnJpQr+VZGLjWFKZsJdRZ+zARhqCMPkgPjUnFDmf9P
L6JCiW6s5JyAAwdph2iixxgNab0fQ595SNW7JBRhen8917+pqHxG1hmySa+ug5o/Ke7yUF2VsoYH
UG3ko9+KzaQBcs0Or/OP/bH2drl1E/wjm6z/G7Kyberu3T1qi414MJqmEFhYj51GAnHIOjYUJ3B+
+mZ+Ll7mibNgUXZAydrjjgFI9V99RViAgdb4wtkQ9NgbQJfUKYY0SMYam3i8rvAhi55xDSa/Zha8
6/6tBrH+dXIWs9cP+10pPgH3kYb6jwU4F7Qqu4kK62ia9EGhYLFf9OG4gtS1W6sR7Je+gXinYFEY
0XO6zYINgYNxxI+5zFzygHxDaI4yU/jdG3rP7qV5q5C58mI+sRpzhm3wQG0KydPxdqP1FBvsbTWs
wO300yaGZqXo6wT6qnMg9MoHak1mE+bJja52ia+x8hkDPeeC3TdXVmCVo1a/o5BWvvvPCyFrl1l0
z1uggSh0eQihPdEWIdpQN/wQ66uUTDwVf1vihO7e5O7gclu7vHjkPwlnyhZgxnPo/mIYcUTdfXxb
QHAbvA1GLtGkt13tkQaT4ZMArDH1svOo8SrJLcZX39tn/u5j68f2E3k7UUD0LvrvxexBPQKN4b9v
VZzwI4ZyXv3Zhba+wsWZ1iCJvPLQU69ad7xjTFC90bV31xZPM4uEXkEAWGg5/3tFvm564Y/OkgvD
3mp7sFv7ze48FYd0cZaAj2iLRTJhPgpjHRtbO5s/T2STWa2acSFpHjDfnCyH0/va0F/Zg9wUJtvN
U3zMhKNrmp3O4X4BWcYuVopnGDcbMK+dVTfTRky4rJ7+FcV9NRHdQLZjaAI3CB4V2SENVeTim6n7
HqAQf2faq49Rhi0szBxEv5F1fCDVkLb1J7ImnpWoFYMqSfB6uj1H3CU6ZeCToGF9RV9IHddCgjRZ
mEm+pdn7Mqd305Lbzu+gYelwwtVltjjtez71aJzb76SMqOSI4A36m0lBGOQbEF59ENkApZFB78UA
dTnhIBEDHP489svKy3VjpoKYRTpo0imn3wDLPIXtdr3yjUE3Icsr0qnam5xC64HoIV+U/TnhiI4D
iwOhksvjLDShjpaOBBqzYmJafh0PFkMRt6DpmXv6hujFet9gqVEC5pYVR2Y8y6MRh8kI1WhhJzOB
WyhY5nQYy23MH8kPwt5BPoRb4cWlcV+QEreg8JdJGYNiixBLxbwb8WiFk92td5gLXxbeEMilRLvJ
zVLbSoWT5Fj96FPog2iyeVrKqVlKVO18Fk5+pwYqT7rf9TwDOvXBvKbUpi0tx0W2uOV3EmWU/BUe
93y+qjj8t/jKmXMtDJ04++JLgLt/RHXkHeucxDtVI6fpfhgIC4vJwISmVvxsLgtjNEeN/7xaW+69
FbeL4ggwkk2xGHZpMdcBOBVsXytbc2i0N46orWe0X2iSxHUmBS50jiY/tEtTer7YDOlUw4aZIlI1
kNJaE3nIsG/seMB8T8wcZ/ikgnFZ8/O9yXmlBVlTbQ1/fJ7ZPg6jIQ4bgbpP2aGKAggCbaedDByv
g2MPflbw6GNMr18wLphhA7WMOR5loNFc31QBxsj98jvcRwUKzYaGW8QGdh1UNnTR4YSJSL59EtmU
6aSAxT8uBrOHbp47Wv77N+vYt86GQHL9KW4hOfYjU58G4VSEHT1SXQ1q1CBsrsLTvnqqYtI1HR+S
PQwjZul4CbQ0n7H8C37HiO6PNudN/8TVsf3Keka+R2JsqKj3KgwsRNwzzy/7jXfEAja31ZXEMPB5
HJuDi1qxB3DjxubbrDcWV9TUbBJ5I28r1/Kt2RuSLYFZoDCt+9SZtwNeLHMlVc6iy+mWNEinSfjK
JZuT/lDVMR+VoDvwRdFpUmOQraUCIh0FCTaMjgKns3AQH88DxuuLE4u7Cuj2i7ikxihcvI4n+Gla
XmLv4eTrvKuPdQlXehyDrwqHeiPxZ/xFrZ8mFV/8ctnrX4rJgbWiieaankWxR2m0rO5+76/ErT4B
dmYXjF14jR3aMy4YvVZrrUwszSdufkxiyf2TtphbQ8XOBmjTqSrZeyBhSQ859mrBf4oKm2e3mZNT
Qv97gCs0RKBOYdJy5H0wmerRfjYR2B4uRbNRkgG7Vsfdc94ONbLv59hZNkpiypt5nHBx8tX+eVdi
GN7wzLkVTpo1DcOzTX/2kDl2c+EvU14jhG9vw7LJ0568FU2Bf2AHl05WkRSRWocDvqCcORHnRBiy
MT6edaYoJNeSc7TPcNuCOid/O9F/z0VV7cXmGYjmvPozmesvjlWwKuEyrmarRNycHX+dlrUISpmt
CYHKB5H+RzzbjIqwZQUmpVQsGz/j6mD57yzcbSzB3pMpj7Ee5IrAEzET9Y/DfYJ4IBzdSNMCyUzi
cwsq4m4EX13FsxqJXf8GEmsupLILWolp8wNnVSTkuN5iPX1ENSJfXxTJgl2soPIsOoFYkZKh1obq
Lp6NCl4aE/mU52X4OT2m9UaIvfbxGlRbFej8vUF+Pd6EQGghoWUnIpDTsaGqil3hoLIzbK3iF8vp
xT5HBMwV/+TzBTrNRDYeGRxVfR7vONdash7iHq+tDav+ezbdKbqiICrLKBhxUAM2tfzeOYTSYDWe
AID6XK/6gk8hm/qgmVfnAjK2MLnH0A8nafASe5pbUkFaICYRCdeFRqpcYgTUB0q/dlBdhcDSqq3s
ela4z3JiG06IZEC6t9KDUvrdA36gr59ERhlD5a5f9ucfGRAPeZExSWQPTYEoleFbKqni0M0ppVJV
CguE1We6N6AbkgbKCBavF1/ksCR/4sQ0TmQlBW6NdmZLY1qGbN7xLLmt7l/fVssOveJjlkEAG7lu
OKt4CX/upXfbvQP2roCgJx4bA5cIeQrioRaLNdUHY2wYmIxItUm/AtG9TzCj+/xdgd/aiWJihI1t
BQnGxtF7cnIIh0a79QNLVB7dFuxUZNssTB4qDENOwAxC0/JKQcpVYrNdpXgdRbvkENoQJtotCobc
ycVc7nYMERlnuKXToPoGWxfQJnAYT3fbNcYIrnVHun6BjfCzRzxB/ckAAbwQ5HBwVS52zOPgM9Hu
TcpWmKyzjVBiorZU1FnTENnMh+Q7d7wYfKd7Z+LEbWKxo9B8jDUp2jaB0IDBgVo18ca9NYIu1Zhc
uKQg7c2M+tpjDlm8BgD8d9vSmdBK7RcXN7G/AKH8GqRk5FGdqECV0uTOL+T1pOe5CByLEMzdredw
7+SJknQq0/aHCeFQ5SCPVoz2VTJnWbHZyLkLLDdnquNKRewzN38K95hlvtTowLMol7dgahQ6avyA
esP9CLKul+f9/pwwy/oQxLjdun4+0baKZ83X2Y5oy7QSvs7RVeEWLQgiEduiaT4JdWnXG5KFOI2b
RAhye2m6SKStR8plcWpTW6/VAtxnMC4jWbNBUcsMrGdX2NKLbwNe/7aQwCJLUUryHCZKEDTclC9S
VdGUHOvlglPfpS3rDdEnbz7T5CI2E8gQIJk9pGPnXTbMHVjkFaEtHbaHXB/hyeXypHi2kU+oPdyE
ldIKNaMRDi0tS4kDelgUpMawIEE7DSuk+GbpIy5ZOZSAvlrIXwY3x0nIPVzR8eeehfvDjNaCIeqG
zyhZNdIho4ArrJW3cmCB/a8oXxHfZILWg7K3rx9MCoKiqRLQr+Ji7a0ki5geIVFwPbuCAtxM6sQ1
QhMVsf1G6RC3GXWfzZ3b8XL6R+raTj0lTACA0THcr0pDuoPq0Y7LPc6cTzHvO87PWyf2toaqLg61
gSxaa1ysBwmnW0LeFRfmTBsNocw5Wn922rwwyrsKYLwqWm1gbKu/Dwz7IuOU1ME8CmESgCoVaPYC
RisGPihryWGLGbytSk6UmPu5kNmLnLff42BRrUuueNr0BQuXjqIHwLFm0iQ7FKMTpgRe14z3zjJq
63aXu1N5MbpN1PNc8vzQr216cRI9oZJJcBo8BLsUfNmi/zqzVx0noFVN3CrLsi7NkuPJbtSfiZdn
mxhg5CB7qT7UOZFjbLaEIp3vCzvOCRy7ACi/keShCKgIJPREnn5rFsY8NHa2TAvERNxCIykX57us
v4HsqeO9UiGzGCIk4Oac6Gw2DYSa5yyFaEC120NSFWjZSfb2oXaxKxrUQpvIpuEE3MAFRTO+n88t
AG6UWdn4yjz4gp8ev8IsKHrufCZ71JTUygpwPvjiZ2bYOxU7Vj0JBglYRcvbWju1u1b6ToVLHA6A
Xmqs8dGkjME1OxI0eWGw6GJIoDeHvxGkcoUQrAgA3w4nhSYVB3dxOvCaWm27lqGqkQzdlZ4NZsbL
wmTpmxcQNwXSf6cimV3WHWv5bEupw+78gICcbOnH6AuHBbomR1ZszkDGfmtAQMpmxGDs3dkYoKHb
f//FrCVqopnTHpH1Eci5MNh+sQPvNTVcBhnQ0fmQ+VAOGtKC8AjdX0E6IITlWzszlB9NvIXO5qkG
100C/J2gfZMabgU3VTc+IYshFpMT57Th9R9wW91G7hjC5stO4qSu7DOML6CnAP6Xiw49dv37UNlH
74JoOJ1l0iPyrw+d83ZQkzoHYdtgLVvAp7a6PMigAVR7l5pEq9ZfUwCoBUtB4mUAdyThzsAbEyeA
2kh39CJovDC6hXTgr7WGKgTtS5KwNjpiWAePgQTm5K9P1x1I2xKVURhXgafpvmQoLOPiE61K3ZMH
QGSzULZKjD4yqGA72BayLj2eFlmElAZOiNrYHhlHTnrc6QynEq6wucMhL7MrEeqcMoMA8wFI1gaN
AQYiqBp8TrkrElGuMqToHUvJIZimdldTvBgexU4/kZjUQay1Pwys921eA1ibROqpPzpHJe4J6uvO
tmmKHbSBkEOxDNcHh0T3PmklQK4jQnmWOKLCPGgRaEs+R104V8exDZ/aeFSWl7QF2dkYgIiUxtOD
CNqA34zgKv++Od1iOUPI8vhU9Rw9gnrZLHX8GxZHUmg2I7mjvJc+OVko/3FOUznnlB33j6yooeyg
vfMHROAkFnkzQHmUzQ3vIsXXWuT9NuwbUTWRQo9xqOZSVoXgjVGQ8/WolgZbnvdBpNOiz1OgDdMj
am+t0q+7hl25g7D7zV9TTurAuWAM26p0bo5gCLRu/KKPsHZ4BvFNkYc6QcBzeQutHhR8WDnHaCl5
yGs1xz0FYYSiQCOKM6+c7Rp4eBSl0ifQHzE1+WNAK2dLmEnjRO2B//NTIU3l6Tjgbv7uJnLmEfqg
kBLFiZhG89xSOSaOXNLqaasGAsz1Qba0nQwxOUJE3KMQA9KdpNY56LrVL0RZ4oCRrA5UrVTBXCCC
LQYvk46UJ2EPLic2H6SHMqbu4DJqo3fW7lZ40bPf6SAW606h+OmBmd7rGQDK/HQgYdVuiVTa2QFf
P8k3A7PCF0PFXhXzonY8lzww21E+JWxzzKvc+2LlZ17nBR2iSJYxaE/RYCzi8UlkYUaKchyy+qmS
DpCZ5KIaSosri2qY3y+rhrYn2YXnnmpzss8mWYUJOqzG/8u6bFA3kajVR8PqxrVxlujt9AHqqogV
q7UQT0Ccu3Ts+wE5l/prqBgZCJ031O6hKkC+A0bHFA6Ua3FifXu7Z5vxbZSBjre8w1+6Uu34Cd9H
UoXRuk3yosIHvo6vkoZeh9kTzhwSLsUDXhsheB9WKqrkLiRzismzZhZL4BGrZl1QsjwtzdeTgNS8
hFrk2Tt1pF/5TxEuUGgJNXY9FHHxmvmL71Qzg2weHu8emX8pQ5W5+u0u3ZDchKwmR+KqKqp1uFtZ
QdRQHhKvBlFmNGX3nECZfv9XbYNWYWunsZtKSylJDL1gVjSXBu+Nwv6WUKBkn33D7JzEpiw6DidL
W7+MD6aKum+FklJ6+lOqyh/GrNGYn9ECTp5agwfaKVO2u7F1N+f29W462oVfqWYYJPw7DXhb34xw
E1nEvwsJBiYwJf+zGlCS8qtpzRB0gQsOu+xkth6AoEFSuzZEA60kqBIhuf17TRnSd6mDjrPBj164
VgDpfPUHXJ4lIYfItQJxcKFFzyXhKbcZlUIRaLdT4WvDPHlE10xmuJppIh7/79aud0f4RGv33tE1
WsazXMuacCsKOOxaABonGn5v+L0a/7vpvQsTuXuLnuN3NBRwsikTmZfsr9PmzDB0wUJa/S5rL0mE
D/CVgk4gHBXrv84wemn/0i3dJm0UsZy9w1l4oTUVqIZ3bkog9iWbOCkteLgN9H3KWABLkyRaBGo8
rItiJ4YA1ZPhyRznXPRVOQDO9vb4U+K4uXiE6rDslX69d1m9JPb9AqGg+mxGjZqXtguE8h26VrLx
2kKpyLto5XAoXUhQtElXa6KIqpp0v9HWR2ups8OsCogEmJOTHp86zoZHn5cpsuB6GeLPCQAXlM74
sQCzH7mtOAhvahD3Xt53mJPsvxI6vYRiwoeW1OheKMlc7CBotjmBV61S781NAoNxRHMgMOSIWt2B
IYAddgW5OaYKYoZWItupyeUqId0gaeRTW1EPBa2xg2nUV+zG2Kzg87gn7gVCoc9QgsjIL3El/3uy
TihpInrC8XCCpEYmOI2vhB2mgVunv4/3He0pYTMwB5dX1JqyAai7i6bwg8dquQc8U6Q0bznitxqD
hfGNtw8zKy6Z6yhCk+TPyzUSSddlFsVfczOyP0g7f38yXXXl6jhPtAP3vm16Y3cQTz3m7soGSNZb
CIzreCt2Is8UZw0Z8tqExCv+uHCpbQV9QcsmISoy/87CMnlway32EtnY9AwTKmk3mJtcAN56GfzX
O9W25HGRrJHIhMcAzo/AoZ97kJujhawZ8orh9YGyeMWoRFJdjQwDDZLNRe+RvfM3AZQH3wru+m/r
SgnmYSKh2jADH2GkiQtCP1dBHU4mbCbLytpn1OdBjrJi22DbwA39+Ixd0/Jf1Gx+K4tmHxuHEtC1
UIbljyuzBzMGQ/7BKlJbI1t64b6ogYKN4ssNoeogsOTBus6KQE3FKzG4O7RcLtSLqxy++cWUBf/0
yFeDsMP62LwmOm5qLjC5vl8NRJVzO4SozNNwNZN3qs7sLZSifX+9EwgzaUw1A92HMGSa7sQPZXJU
TKZSRfNLOxub45n8yUPtuLBjhSGsjuh/5gDlfo+rgWQ2Wa/UWIhI1oq65JR4dWH6Vh6r18viz8Z1
GMXNRBrn2Fv4HLaPgxzcrPV5cqxLKzw/vU2rFAwOwoZu/2q14hsrp6SzuEg9Xoj25Y3pHNMsUJ+M
+kqDiSm6bShP+7L8v0Y15SXc95aDQc4tZHKn/7XiIMlNeTo7A9IG0Et7M+LEhYxRcWfWCI3+MH74
YhnZ4N8uparP3WSNMW1I/8SO3T6Dy+vfodqaEmu6PftCfCSmOUq+l+hCKkVzcl6NABjQbBGEm5ob
7rFB6ejyGTJsA0diGwdhD9HOKEiNterLQ61aHKL2r+rMMuBZMgIRKgB2yglR4n7dtOeFBZ+epiaf
yVAzKhM1GwqkZcEsRpx9/RfdaTKzcbvaJJuEd5DCu5ujhFQsPEZAA70r4tCeFXxMho2XeNJQEm+f
0x2G0hkeOoNBXidCzBPxxO2p55CZvghB+9auD+Vqr4WF+Y6TrTVZEdawJG9NoWrKEOH0R64MljVj
iIH72Ny/VgStQb2ktRO4dNYrEfAZkJYRvLPcfw+3l/07ibDd0zL8anORNEf0QVdwoXbf+fCDNwWT
ydOt8bljvh4VPZG4gzv44R2Dw5ZNanTfRNYhRtAebmF2kAXgN6Sq1UIrzbYU4N8zMa0bxeK2PDaC
L/lQMXeXu7rD7zVBOUU4wG15DVWbr6zwf2v7UlsAn/4ZXRHEFK7sGmuy99j5//AdE7/EKMwhkskk
SgOBncu8GfhtZs9v7PNDTALkZpgROdt4fD5C5BBJ9zhRCjeqTyQx9CcYOzKu9NTCpr3sz3PTel3K
55WdUm5gmPNxGLWip+H8mO1WUsZoQzMGliWD9wV+Mo0KMlInx39dg0YV0pIDeSnZhRK3QQthp1qM
z3/1wiAp3fDjUjL34e/R15UtAmWQiZkV0ChEfBzmGRrYcIA4OGCBqIdTWqZjBo1HrBglu8Uptgrn
afERjtNkS8vsYyhwTYhceQNUWOVNQrz8oZ8+HMehO9bxfZgNLTdRRLaUSqFhM4zDO6ViEO0maGg7
zp9lVOJyJKyh+TS36Bqc2poZ/CJ35knKcMdyIfv2ZiU0lTQVWZKBXycPUv1bpUt173UWTc4abkwl
vybZMk+Xd51gh8FZxx5l1cPz4LtwHadxzW1ZY/e1QpwrjDmh40I1Blb+VWZ2FpswC5H8OdWXKWcN
/1mIJivpOh6/ujJCH38MfOHckBIuoW1KJyc4NVbCGE8RFScq/wB86GaKoIrcx8YyMvJiZ+iz6QtY
0wtmUp2XTgvGd74Ky44V0wnAo9POsqBFmKXsU2S5buL781XR1JYWK9fyItbYIVODjTZv77zE8sWN
wEOU5nJaN4Xx/vqKMbXsHGMfPbOgGrAKDrtKtQXxTBM3RezjRrwMC7L+JzfXIxy01rRQo7tt5e4v
9X9PjluCxQHRWiFuUevO11WpuKH80j5LVGXZHX0lj3+i5De0tkIFH9nvaw+I4CaKFomy+RmQ0I0d
rfi+suZAKNkquc/Nxm2DyFGrZaRolQp2+k2sR0p4XSlNUztbHRwDCR7QCh+QpaLCVQhgQUWcPBnU
0cwKASruuCmIiR4/D3r1uslNltQ5rNtojaMKIiT2RByX6knzyVUpNli63k+742ERi7vW2CgJG8eo
oBULNxNDwMTodb9wmLW3BGFXF9i/LiCY5/1xC4g3o8iwig13jGHmIWMjPp8MnvyoXMWR+l7WyXni
LqB3WYqE/xtW4TvDpufApuOIAfFJOCpxHx0p9325jf38hX4ovPp8ZJeA+zYJ+S1lWoK2T1+orZfl
wJNVrjomIf8HwOxb2OOGy+nHwA6HjNcJDDJL6GuCfKaIqoui92Ub/Lg0KJhmxvKQX/bZsVpqCAnd
xWzgRURVN2i1Rrp+XJfBb/18rmEOeXG3SsUmAOh1JeZ8A6+6dWaa519BQhoUw/BcpaouKg/qHTod
F/WQlVKUywmvANJz4WoH60o4PctKQSigZRUjHtbyR43vvuakxofVwsQrzmQ+Tl5rHr4AO0tFvaTb
mRLmWx6na+cP3Oe8kYeFrR6uDV7TmoQSuS5SbhMt8D9GNYIpciWAKR1o9tImWmIZKSERQm1hZb+n
pC/lAIqv9LKegcWSe8DVSTDk5iVtCSb26L0Aetlj9eVakggfVvIlG18ITdLk3tRAXMRz+q4no0Wz
2+kB9oTPy1p/2PbYoXdJqM9ZbSlH0S3n2pUkHSOEMsQYFrQAtARN7/HNmN+jy9pFRuAA/u2G0ep+
v6/deGyQpIGDLFtxU+PgHYepgZj0vG2UxQjdpbzfF3jDjb36ZAfsqp5z56QcOo3whaUWralxGoYn
CeFXi5pAEtPXPkNOeBAD3J4R1F27BbbCS7bNStJWmsHu1mPNsmhSKq5FnnuOl2sBstbb0T/e/WRt
x0pXcNiaWJuoasds8iCi0fV0V078IfmGQmY5ai9MID93E3T7+uG+wIkAof5xVl4n+0AzITqjqmjM
Da2GVEprET8R95hl2Je4TILswrvKS7gH39uDxQk1erdkfRWj2QB0/6rPcrH0oPzzIP7RnoqCRyIf
TKUQHjINUqTAEYIGncacZoQCN8d2Zo4Dy1CjkwqJL4To0m95BOp9JXxNF6L07Sah+LaUnIdJ7StY
55YUuyiD1XNQdGKnuB+3ZaipAEMPDyUIIOnc/s1kJR/p/jMwzrusdIXI2nQp2nJo5bMA3r6+T88e
hZPOR+078sKO7RPWKc0yUOOKs9N2hwEhkTvFx0AKafIzMtQFUNiPyiKhV2T98n4OsJJHbCCW6XIJ
keXgUHD0V/rKgyJaTX8D2tfbhWZemfiCxqBtbY/orsaisqOG3C6P6D+A3G1nkuiRg9GPcGZxVfda
uv+mqF3jo7Ro1Z/f1pbByZ4BP2WDS/HpXONH1MV/sAnClgLqeYCpjAWqsUGFTdU4XfOTZCPF4+Pz
JzU/h7hre6NQOwyXDS5WBTpHj9DoTSqfatsu11w4MERZKNwjzjmD88Clx5HjuZSYvUszB8I2LFl0
BJ6ai+yQrtU66AU4NwqTPD7YeRTmk1tVqVKn0YiYp+lkxrKdiIK1pj657Yx288v4haQUILZ0pkFh
9W6Gr1hlSynEmvkKM74Hhc+lWsWjKOLMhFN0jyNWh4HEwST/2FH+cg3/OpYVFP1Yk+Lh8ySEvm/L
kD+sGG0EgjNgNKALoM7wI6ZwRtPFYAe4E6BWzGVXaMr5UmV0d6oVDfCm+ibMYSrWitbnmICYQQMw
CtpOPeYpEJNXbQzJHv6m6J0xJsXcUzlR66njQqj8YodulxUdKYnNUfUTfOjDoZ08wu1hdib6ZFzF
jNJBWop4hnn4FnqP/rgFkeQUpMIeEbU/0C+yK3XJviCAi14Plo+rb61kIQGYEz7ARZ1w6gLyoKsA
LU+voyHS0TLhP5EJ1DwxGye85QAvU4FM8EOd87LXImPy8NqQFuDBJGFvtJ+NPUgn8yA+w46f5PRb
dg57ruqKNpsBBg54hnSN67xHe+Oc4IyZZzRXgVkQRhg/W2FoOqk2aupzgbSTDbyuKKeTVpfHDLKg
MtUAk+xyu2+HVaZhQeyMbYyQ1vO2DpLZVT5Z8yt6DMpKOZuarV4QmVGpl6QvBWU2Jviwqv1vLBHu
ow+RRlpe9ZCG0/tLmRpkVpbcZPIBzLZIXDOp93f2mlfmLwNRQdXNNRBuCYKJAXZLXBXC0UyjFxpx
csfpJmHmtLhumGWq7VV8NdVgfemOoIjN3SMU8ioRT220yzjsiyCF1y3eebLXMdzkt5qLvysI+fex
+VYQ82EXVz4EL+aZ4rQo0d3qSciGGAJZdDccUPCEgDNf7hOFSraibmk8v0a2GiVIq3ZtGB7w5Xo1
+UEn2clIGuc4os0Hi7DQhYfwCLm991hS8ran1v6rXYeQfv6qUXpWdfVMB67Wj1WRZaZIN5JgGL3D
VAfOU7npn1Rac7FzaoFJR+/YKHgEsTCdRc+fjxWf70sRfJ7xiD5ojSdfk6TdkqMA9h0bOgPXmAbG
9LisjM1jvw5LfTfmujlryprHatGO4GEGsM3Ac1f/WFGPAWpFEWIGOb9bo4YtKIbaCTDSzWEFwgRV
VpjckfwqGORC2XtPVtL8RQzQAxRFnBF7Ib+NibQers/PLu5j9CXbg+eyqH0xx7a1HW0kUlufeoDf
bHIdrV9sEMHRpfN8hQkQZoJra1rlIKnG8lxmaC3bHdBZkq1wP4S/4h+nzBrueAiHeNXipk+3Xa5j
elpz226QdlFNtZKcloaQb4o1rODHAks9t7v0TNNq3QO1cmNr8CXGn/ADeUcVaSycGSkTJbLxBtjH
vrLRgGliIbR9AQp5BGiOPxWvfkO1hgiBqQuxp22F6p7U3vIV/zsn7K91Ig7ysUZeZ3Y7nUMJLLcn
Rza5rj8re17gRJaPSW7bwAlq2e5FkQ8G3wmaNF8jlUyORjPFGZxwQxRQVpX/inPjwO7LeOpP8wdx
WMuU/wiMo590VWu6kaz75Rhar6Mchh//1diZXeR4b9sXHdluZ5rWFxX8Ld8qgE6ORULU8Igolhsw
GP/CcDPo7wtBrkgh9xrfwQF8e27XJrhHxAliJy7RVGxSM1bC+68RR7iwhe03RaJC6m9CtSQGXMjg
FN6oSRxsz0beg6D/B3p3K5Ze4opQsZpVHa0Dp3Jqe7lTakTU86VZRUXcox6aInae1/9oMp1hpGHK
vtH2p72+Iv/5ncE/eyL61UszQCEWyAYo2EePkXV8oXC9f0tv+io0hvasNs8tarOTZCATpZBoeYp6
6ctyjOHeTQWAEzPkw2l4QetBS5njPyMTfjQPRqm0ae2FYHvFcib39gYPc+wWmiimr0mtIuIjk/zp
C0MTYvnALa7sWIiwBMybsRQftlYQ2lJWWMiJ7jfq2ipqu3n5W9VYB/XPNmDv5vY80MzgkMlfSOKb
265pUwMboLM51AoZviMZ6wTbALAd7XFL2wfOAP5zzJ6eqFnZeUcvRWtLEn3RWfbky7/yODvRTkpR
siLaEAKGTM/Wn+s1vN/iiUeioE6Qt2O3xVA3xIxNLWOZOUc2lN4ThfMkKxYBefpgePvryBQxN0cx
cjEPgEtnUX6TOa2okKajnGNWqO0w8jYuAhn3t4/QEMHYBOmLnDgMa0sFo6yXckSHQqWGA1v6rSwq
aVEc2kt8qE1S3/fnfUyk4FFMcB21VLNEPkRMPMW3eNMTn0zdRHASmT4Dye2/Cdy20TNp3jkbn3ih
Ch8gsJRdslYdZ4kgNDzqB7bzAM9hHM1prlAOFNNDO7QCM71hS1KPDPKj3r7nPgajLD2zyeKn5PL1
mGrZvdCt0j6BXMF9Se9C6kb/E3dOQWSyP4L484CIeeUsv3jgjLNLORjK5BK5FOna/Fv3jVFtRx0J
aoGcWV/XP+gvfvplnn8/gOatVAnuCeil4haXGRJxysVIvO25K4dsfy7z6QcsfBeOTrPJH3RnwaeP
UNG2mZM4anh41hoKkM9SOwjIU3q3ZCVxMUJTm5CDpIJNv//P2k/Or65hJJN4cAOX6wBtu+H94T/R
9dU2QA9/OL3vlZUSx6Lij3gSkwrYoUJMPC4RsxZ64bX4OpO0xaPLSczHLM4n0no4Ivxb0JGigb/2
CJnu5eUo68WnMcRPe+g5wgZ9TZuNj/9ck4jlKl7pCIdkE4H4arnL59zOwUla4c2Sdl/x3cYUp6b9
JhelC7dWEifa+hmD0vxPV0KEBnu70l7hXKUs7P0N/gQf9PEE6le6Y8YVYwlTNs8cKBdavLMfMesq
NQgEunjYPsc0k2EP3vMT5ZdUYlyIMlkAvtabcMhQ6Bk/yYsB9v9M9Sd1gSiMssMTWaxsGi3jiOZ8
Gsu2zCih5hZY0Cz71tSvhwgm3l/pEFa16tyJYux998W3aP79L0Nz4vTHRUO3lsxwyjO1l4ERm3hD
WHV7gzDQk+QPW4+8lJ2L+BnIYl8bf74sbwdEZW0rlwLKjRX6ywpWDsdJdBYbdOREmXjLd4ZgQc6s
whGUTvSBt/DUrKR05UCQgpaxM1lg0ELJOFaY+YpAx+zNMJCHp/hU51vew7nkzPEsSMKnEOog7Nx+
8UAVZFgBASJqqCBFlbSbZUtuM06Al8dHIHilF8jbapPbb6njKGWEIvNe+UR4IPlbemYgTXid+TOr
1KC9lnab7FLIPPoVjOd5xdxaeiK5kMlYFXWcdjZK3NGUHTa8s64p0H5dQHHZGfZTzJX3vwx1iJjm
JIaClpPICWMVbZ1RBCiRzurLoVk4FkXPROi6Bc4Uq6IOseyrRQu7Eqp9HFbIR3ObHxqytXd2+TIA
0d3bLa7/uR0V1ifgcHvrpuqKxRo+X5AsmZuN6LhiYOKmrAZDz0gQVjwszDoTZJguyPyv8h4W4z4L
WLckQPzSXjgEYX5ezE/pujA7IQH0w8HZJqSWLDjLMb3mpNlawjaDrJE4ozdIEa8MmmRG6ohaXysy
wJAcJZf5L9jqhoM9V369En4YnLvaX9XNUCPxnWs72CSHHgm1np1FEcP9slQQMuCrafKUSPjIKtWJ
DOlW6xgnm5HjiPbIy4i2guko5aiQL2TA3Uvy+Dr5J5e/lB+ww6Uao6L2t09KZusZ2RPAw5lkBcJ8
gXT7Zij0O03FzeLwqCgP7eZ7w5uoeUQOTlQ13FsBKCPB7MZ8tvIJfYRNmILSNqmz7nzvQurCvcer
EUmAN3NmyFTOOh6rTwjHvsFkV5W2XxF1seiGZA794DFU5BzW3NfHI6O5nKq62FtSntT5PLVvFZid
oU8vC9B97B0rjCZHsyV6IfK7nMRQPQ6XySXt7/bED2lZxQj/Jfq3vt53+ddqUyAx6ksWIaOFsCrT
DQOZmunr+LxjIDCYtKM+/Urq2E6XL11SA3/sWsfwN4QKACfRPzuBSk188nB+sl4F9JzxbrllG+Pr
zTofFEYt0D+WiehS0EAA1KeTd02gjH1NBtQZiRad2lh96kii4FMd9aIP+PE2D1vjwO64cOcFW52Q
xTtlotsB80nnXivWs3Rcb2y5aHnlNTFe/U840eqCFqFjPqVfz/pDj6TNSZJEdJaoUxWb9OgvA2LW
fuXMVHoyK3kWxLVmmL+UYeujfnNLIhbNtoUYwZyfj7XHp2y7/1pPkTRul4wczY1REga8BgKr2M/s
mBSTCggl+OBiRzGd8o23I2TMlbWnjilNAn3L/WCwBUaj3rtnAHlkVoQ/P6L6+pq583AnAcCUZNbs
1zt9B/BFBZeUXuKP6hDC/8SeW8RHBK50ZIHPUYefGpRydjobT58caPZA6/iViBEkECLyFV9bt0G5
EFX96evMtB9zvSOE+ryaI2mRnBpznJPkApDLSL04SXBbpRFL8CMcjP3Q/Y/hEwH/FzuYh9Eyx2Kd
yc2VlnQbTOjjwr6SJe87rIPeuwlYqpKXS852lqNRczPj+jpY1FOnyoob3/yE9rU8Iz529cdzHrj/
tQvytetdf8S0ViHm/zn58FqM+VfK3S4f6URiacUs81ECc28NwsTNFd6+MfN4Nx+G9VCW7zPuMK5q
pGHZEPNbKIUAuxRD7q5tPhxjE1PHV72JEhCr1X43G4emKiUzrpv8k152rxkfWQlMiBAfZ//K2F5I
i2/FxoJr5CsNcj+7DuPxfrw87iH8zONYqv0fLFOErQGfu/Nmla3H8k/e0dO47gPPXOWNH1bVAJI3
r/bxkr+JZf08NBdta4TGYk1dlBh/3SuuKtjXskoVtcEDcUax+TNe+t/FHc/EqgygkubBkNSdes5q
6iCCv4mRwj7VGcLT1S3HeYALO8KeEw0EDsq+wWxAnCwG4RMhXHg2NgHsvW+MILhKIP1L/JQbRkaO
yCh6tWan+20brlMmAuF0aImr5F92kI3k2GH2rJ2g8EfVH0ZoDssdsdFbTVSakXWN1zTiJFmyKcGw
STmKQ9sjCtCsYjRS9AQ2xOfT/26bSSigF6nr58N0jm4YPz2lawHzcmhrL7Z5BH1nAHEZO2Ltwg4W
Y56pF0O1JxIHFVilg+Mcb83hUFKGasClmw2SolCsZbzCZ288nIC6PiEWv7e0VW6ZvfNgLsiWq1yx
p5020rgEYjSDHoO6aUjDUH6mTuPNkf1gkUWd+Rzi5/TFb/60kQ2ev2XwPUfSwbKZyc5lGwupO5+a
5Ugop/1JWliE2ML0wCYSar+5epI7mmOawI2Gndf0b51xVaZm3qXRJGE5/s0Px+LRlAcXoDBK4YKQ
soX72WpZPjydQOkxmEUmIGf3nnF4sEbKTB6tWDESIPzOCuH8Ld22Kd7HpUNF3Khc/j9+hIAGKfz0
eVGZkynNJ5qs9B28nIr8MbBUA/mXaPuecA7zOA46WvXCMnzfj7v3Gc03sVaWHjeYAEQpsALisLAC
mbRK+tzXw7d16Qvexy72QmvjK553lybk+mWBMDEV3kTX4pp5nUljJ/FyBbO1wQXP7LeZLhovqrx/
jshGgTjb1uR1Sv17iK3T5iglQCCNDdv5XFRKVOLv83ouDsujMlp8gi+wCdmb7sHCWPtRHqtLT4el
0gxNpxgt1jImU0EabpqckSQkwfX+60kikngCaa2Wbqjram8X3z+SkSoOUsjOlVYd/+n6cdc769zF
cJssLJBcwj1Vj8PuOD5U8+VVLuVN7viuCq9e52ciGhzVS7SaPhOzEYizPn5Neli3PgpytD/qUbq+
wPE6nHnOND7u4p5rMmTGh7hXd3Znq0/gOltJuFhemOSmT27LTkPJqFx3MfP4okIvI6n+COY9eGn3
8cM41BypqBzfLpxpSxNggnTCCeGGAmMgWZtXpi/fJ1SA8PjAhbRQJPX6s5tdB4xbzv7VBZGyq3Jz
hq8PvG3Agf5m06C69ZYIESqjOeW6D7EpVgqi0HwPdhzsPKBmIPtaSNqWxbnpfCQton4Fc1aueF/M
SiCXZBpesiHmXK2p7Iy1VHq1Nc4PBVOKY1k+6MRruNsfDTazAxq6erT0tjx7hmitosqVU14OtBOe
fj0moRPBdhq20txHPnTvc9tUNcTCbn52alnkfm4RAHQP1hMNhBl1LX/tsAm7kaxJII6n1MeZzE9S
nPtIgkO1DDiR1DTkzLkK07PvJrbtQ8Y6wmko+08eihs0peqxOzSy6Xx7Ds6GvyrFRKe6ZSKY9W19
EDKbt3lvV8CKWdV/RbzMoW5relFFIT4eUiUjwRE7xGqu67Nf1HuNlkLCNk5PjO5cxXpO4tN1zDpZ
N9RKPHzmo/YoI9R4GHpEJ6pouczOu5AICXx+FYN/hD2zLvOf/Xa8Yj4XbnAaPbh4bIjLquFFtp61
+FCbXihSKiOBvjQAxy42DhVcit50+C5LgIW0Pm/G90XhzJdnNLXztFOV/lHth2Ynd53SvXobGQhF
riVMlhet0mfg81tRi5ht4uILT8z6BLwfolUAhtnejOsiPjjHmj83yD++E0mgXpz3QhBX/j/+qdhu
Zv1qqpYN+TyOgY7JmselJhmoBnKf47kRoAKBuFTg4FzeIapIKVLI29ULTKlsiAvNhzbQKybYs/vV
pro/B1iOLIv1/oxqL9AX41Gy9331E9stjO8YbAuAA22h7b32bNyPr6460rvjk9/QY1obl4TMdAfO
1rSkUx5OO1xOZ/zQZhxInfrHIUJHIMe7J40AprdeSPADCxy56e+KpPJzlEqmx+PXyKJQeavnmFvk
pNMddodhJfF8fQQFpaBm7bYhmgI0NgC49ya8WBR8ncEBrTc6W4VguKg9GAPLxsivhwfavTdcQFXG
8XMxmw45VknrhVUnAhUmW1Izg3AZQWkBczDEYtcAfN3cAgVpKsm/uuxvvZ/WgkLFYCVLYxlT9g1j
rKWYS77kzwPaxwQ3gUBwqXVtSNgnvEKKLt7xirDfVSyOvOKZpcRB4yReCKKeVOapFKJf12RrOGEp
9mBKlvHLBvVY8LlAC5RinY9jjFnMFfqT4pl6+sr2a6YUtafC6qZ/OjJvsQcN6QoT/cs0wrGyZE3f
A7wnbnvMYJRQFt47h3miE16TKZkaHFtzzK5Md+DjcPn7Az2klXOeB7P9QiewmcL2CcUW2Y8vCdWt
xCtn/WzHLzypsL/Kxzt4Ubs45PtjM1W7XrcTupeT4Ta4x0YpJyqy3U6hR1gK0f8qghoq6YRbyP93
WUQlhnx1F02eDhMytD/7WQewWPC7ToHp+KKbic5BgupGN7z4gCsMFJzZg3PF9HgWCQlZwWTTD3s5
W9DLChnx39ZpRfRILcuRoyIXZZnUXCRpALFxGImzUfIJhNCC5qfHb83gNiy2EEewgKrPq54zMJM1
CMgDRCMclgvmQKqvR6E06t1CKEmBd3lBFLb4qA5fZaEQdKntXu1fdts0JA64we52R/BsLeY0YMXH
hTWZNCj7BPc6170D0HouTS+uY4MmdNV/TLmdsjTTOemj0BMwY8tjSyKEgqOk8CNDNoHKVAH44/ex
DHxn1Z62EnD6pzIVGWLD8C7HO0y96B+x6ks3P8mO7+KFNXgUZVX9BXWPFkXTQoqH+eLt2bsSXb5s
oJmNPGPCen+TQ6G0jZbvzMUW7lYQgvUG3JTwmE9KaWhTPX9RR7RlLHchGo2R14vxj8Rwrj+NY7CB
eRsudH369l3hVkSbM54jM3+47huIy4fchjeGnVUpGfrlZdqDGiBgcjgmg/6sT0CJaTy7kOjcO6eA
YMkJS+dbXHRALWrO6KslWv4PBsgUIwo2AYkZqh6mz510/CJehl6sh7SaxK1B3yQIfyQCjcuOIF1A
cFJ34Wz1mA+Hi0a8zRltmNW7ZfMXxw6JgvtUi4ItuKRbrrjDl0rlx13ln9WNySNwuJFhgL2c7jKY
35OXAOR5e6+kofoD0uf9aAtuqCwgiXcZ759pDG4Uw8Jh5k0DYv3iLWRPg5/9+B441+iN8ouZa2aQ
avHlvziYvzmdOqKD6fre2EGHXHNfySEABMqzWkDAazXOQ+fOE9VPrQqujZDOI7SR9UIpgey7obev
SqoG8Sc69Jt6ysCat1hebg6YdIlAxlIm1VZlwBm9+fT3l+TWHuYuebI+c9RNvKx9qO3xaekPBELB
JhAABwplMLqxdvaDTe51lzZ9wVzmY9p4B6sZDhokbCc4+3RVablnrEjjY6e0XCRGgzu2Y+CzTYxD
/itcn+Ue1GXkTq7HRLc++OC8jL+ZEI+//sUQym+oA8DYEtEIspk0OhSEJdzxly4g/0ILyAf0yYvn
QD4JV+pBfTcJHeKvFdtS0hSPWoUKQP2ZJOvz364btH90vm4nVOiaVyd2ijA7sK7jkAsLTpU3rzXG
ZGHCAeqiGEgDvt51uR1/SKpTmV3ixW/xQTvWer18Vpuk9nWoa/lPDskkLFbqCblNxpHvL59JYFWS
nWvC3QE+s/6aruQCXK9Uy66AyfvbPB7pxGnWZOgR60iA9iowbAWhmCRc1ZSUpK88v7Hb74LbGvUO
gyL0t8MkQQ9SjP58Xn9c2Gnos8gyn/0HW5cOmWED3wk8yEKAH/D1x+Iv5bPwQCTVH3J9WfejvFRN
TnVCLNKaeygT/UBzKZwC9qtN0ByMnEuE3xpWlZ6GkQXkvjsdnTUC8VqAhxKByyRIo3C/0mAod06X
cWxfl6NDFL2a7L41Af9225JC9tzZLzfgB5T1d8QrjajWrVQ+j4ANhXDv4CzG/M8pPu4nMX3evyC9
LoNoI1kTrCuUiT84QugRewyUJkCTixByuZNSe1GdNMHHVbpExOSBKt7bvNfGQwZbCIV0ah10uw/N
6QxmrtYescXq4qKepeLeabLjWaPRBVpC8BRx6Pwl0LKeSVABw2yTSd+TeCEDGgq9skABS8XVEfDs
i6VbeD+iPWCdNtiLQaMg9tYY0HL/EkYnTevPAZOU9GMHHHu++1SWlmFlc3C5ZqxeLYtO/HN8Pxmv
Cbclizcn1vArJKQbSUZZylK4HI8ejnFucGa9RP0qPYacwV1UjtA1c/jxtQJV1j/XeYh3x5sWE0qL
O10tDPewt449VfWgUCprTzc9Hv4aZ0BRNbQO02z3FlCa0KwF6ooQvq2V59eUc5n0jgXk9IvL4iWO
QtZ8/UzwSGwPzIj5MwV0CDiHcpZ3D/ZamrJ+WeXAenEq/sB405a8MKuJRy1bHMrGvXz0BqbKPhHJ
MgHepmmOGvAbf+CJweyHUP9TawcyLJ1hzcbpwsXNlOjM8Mq8uCngh9M6e/ip0SQGcDATAHk5Tyby
+CJc9ZDUVVZO2jB8dRgktgU7ikz0HvwNZT1hGmVvc2syy6kCjivkjxr9U0LL3WpJsK5xWjH9jC0x
HuwVPTB5qezXRxGGE60a1vdF1zKutcms2oLvnRjZt/ZByjpHFDsBQq15iMubM2jeC4dDkBrfnsok
Lzf2xFyQe0SkbxzZTsR4VMlS7KAZfrDWHkztv6d0LJ/xqgZqSC1NHcxIY4ZbLR0o2hXChX9khxo8
Y3mLhiFlOdxeeOyFkMy13DQOeFhmc5koOc+TXDFzASEgmmh7O+1+0fhvK/BRPYBCJ9mMeNqfVD4+
f4RhshxxfBVPDhxcDg3J+TViJQKKPJH2Ck8MAx9L4nH2QZgCMIn1282Gh4192K6mWGLxPKnpursZ
J7qNcTzy5jp9rPuYthdKlC1aolE4ew8pv/d4x9o8qA4kkhxtCqXTVHYpK/WWP1Dh3/CKM/7JeUJR
tC9SUSAfQ8eX8CVaMsvAgzqH2ledbVB0oAeXc6TO27V+q4sNhP0/qzhtx+0VVW3RH3Xbeydh+7Rg
o+GbEWSWbijfNgBX0neQlGXzCsyAnX93AKs8t/+BbgWN+qOzrY5TVrJK9aMSmwlmUaEe0sO/26Ka
G4DUmg8ua0mH0utAcfG18D+yzI1lDNU3iBvB1PxzGBm7oT1vkRvvnKA5SuEY/774aaIi2AuUi848
39EDDAsI0bg5RZG0dH5QK28KiQljrdU0ZeWv1h8knyoL1uWCPQD7xnYWq78XmuC8E7FyvnRXujqK
8P5M+mP+7p4Qrfy5lksX7kBwz6LGUgTBnGPmNCk4sMwGnjU7Bvpz8ON9gjQevwV8DKhk4jsQYz/a
nKNzMCC9RAdZv4O0jLGDK7WrLlvaZC1sPOyB4GU1Pfp6pzSVrID9OhBvdkVD+JGXiF98zQq/6Nm6
lznxnQsmNurzuq6HfBxYmAxRQddJwrXhVjGeTOLIwxysZ1iFK6rsoqglQ7in1Sg4RtU/KHAVd1vS
8MkBPZUIWC8pxP/brI3xdnE5VYln9i2ZRgersf4VwmM/e/FuCZ24gbm1vWl0umLkiN17EG0xH3/c
NCA/1jPJ+Qc6VJ7hTz85G+dju3a04aMPJrDRdmd9lRU4eIY9fupC18/UOrGem6XcQxdYvQb5oiVz
3ANT+Zo4Y6VxxozX+an0eDhy/EvFbHoAtiUOf+PHvweynpL0/fumZZi2c2c79UweNJaxiLE8wZBE
ctSXHg8pZYVPGd8K5n3RfhTnDPoXAZK1f3kqGlDY7x6VChRHXObfJRubnRCwYh2sOUbwzQaBrYJl
xw73x/w33227X/BbOphsI5Zon2g7rTdOFSZg0dqhI7o5fBO30hbrJnIB/cnMGkly56fxuRrQZB+U
F3simL/UT4xe10YvK3HrgDzLy2QKIgTX61zhcDCX6514UVTkAPQn/aRFYGxyKcqniMXxzBkfgGRy
fKvJekFAvJKGbXtOupvFjYOOM1yQBnB+3qCzZXWb85ahGwPw4R8H6OXr+pRCkzefGTdQ5kK78t5J
tqN7/4RbsHxNGrFMuijE/wO06Jrh1gyOZ+dBsZkB5uBP2HapGltzfCdzf7Q/rqmnou3YPykTpCzZ
pPYr4htVhbivO9vYBLryhWGpzZVOAWdT5OKOUGLeG9VLQszUtkYshEejDwggeCeBeQiaOR30QHc7
R/Foq7cwim3gU77B0NnBzsI41caS82bvqvOpuxD5SiFM9q+DyRphSQgnZZKJMbgqnIhRRC58/ZlV
Is4R62pFTU2FFjnG5cSfDdBdq43j4phEQoDMKX1BhnC7viTSYnLVI/u+ZuVVUsXH0WQACI7K805o
esu71Zn+XbUK8Yy8Eh/D0tps4wNk4S9YS85bxInm3ezn3N8FW6VZELtKud0ncXOiS/01mxSjNjgv
sW/2y2jMpoF1ESMyDR0VRgA6jmlLPgWwjC9/i0zX0FRW+k3Kf9tPHRLGQWOAILmwhP4QT1ROgqFK
MdqG5yG51Z0MI2SJqtfl1MRdUIrXr4HicK01hOplwbf9/KnUo+gBHRJWmsUDdVfEIEEIEfgCJzO7
jaGvwb42tFH4n6DH5F81ZbSt/dRtVPy7HCF9o55pd0XuYBa1mQ+3/Xk0ttfevcaW7CJJhIe6iK6d
lZKR/q13CXlLLCrvOy+3w8qygrd7xXQTh6qtkaaWziySg0wbcD8FgauXHS1sgdvf6/URzzS178Qu
StTEJO2886nMQfpnn1fX/xvYgLrNa/m/beZBtsBuO9BKBP9gXMRNAF02Zs/7VdstgDyklWclt6Ze
jK2PsUXZqpeTiIKC6r3D063weX+avmU2W1G2vGvfSsqGpLGm9CnIQZfDXA/MfPePf08bNR/jUxjR
1VhstL4RXYZSTF5uZrlEq03JZ8wFGJayYrPdLVUY+GoJZGSRmVGazizHXCEuZCf+AzMJuqPl8LLK
ApYcj8axSlguPrrPXZtT6ZJqaoqlAXw77CchupIEQyDhccQy6MjovSFCbtZZfKnbZRgUtI7Hm+84
uRbGCRT4ni8rUuPPMEM4fOR8pfVjHyIJmoZFzciZSbp8CLOfgNmw8DC+cvhUUR1CRfacB+gqO4sH
KHw+UNodL9GSkIdY+Ty1y0vIVQI4/B5o99ASIAEMKcrKJVkmeHgXnvc0xs8YdVOgJrvHqNZq/fTE
7VUe6unfYPiSv6/+86cArU3kD2ykLmxyv/kxHQ0LpSp6s0uceeAIsTvwsCH7+T/uGwMmFvEyCZvV
UftP0/Zi4DVpqB0a9Sz/Rqm87Q0L25PwoEszD793qrqhhCARtP3AmzUAjbRCdctV3/jZP4D/DQUO
Q57HpPiw9eW2neUV5AcvTh2SMvRcLrGKVCnfMhAMuXfo7as3JeIqDm4NTaNoXHn4x+U8OFN0v/h1
J+gH9FuPZ7nP9zoIueHr0qPeeit2Ao1JWq2R5AGITjlAcKv8wB60ceDL4wpjpcFZQ6uMpLLIK+SD
UBWMcl9WF68U2/XMW/6pF/ShWFLQyUkP9BCM0FuIpJEnafNcPjh4q0Sp3TcVSlLq85o4DWYLlyCm
l87RWy0sV9wTv0Ya9gISIXrBc2OEN/XchdYKXa7qzd3g0pYNuplU5AJ/kotTZ4JqiXfpVyFQzB/S
CS1pCAmHpScp3v4OtFUs9Emr+YEoAwQSzdPZimiOVr5IVEFgYPycJ4ZDJYFToXqknA9+uWzTL1bd
HnPH4VESaI+N2Vrq0OA+E8fe9LLSGNQvRH3N5TXLK66gl97Q/JrKujOd1+eFUQHPXO6fgV087CnS
EUtBdmqZPlaTG9ZkX5U8aLQMl4yE9gcrDA56FYP8kJsn0Kn1U7ve/54WBRFQvlw2ZAdH2NBp4Ni4
JFbKGpntE0TDAO9kW60wk3t7Fo6YVhJTR9IwMlRpJybrwl0TKJlPiq8am8qOvLohGAC9UMEfSHDg
42GZbZnzUK9lLEYJN7zBb08cs2Mw4fxE6fzFbC0B0B0MwHy2dSSweeOpqCh0U+tCQSeb2Iz7+tcO
qGH3uCAEHIG2oBwlfzmk6h1663ZYADG38mHFH7NIlPWKfwjHIuh8AXV9bIlnYA1CWE/9ObVDYZCO
0QiugPDiCcN3TIh9z/ZVVt/zFcabAHs6IaUOA/bYqjmLLVYvaKPD1ndoa5hVFq1t9ix+NzHaj6Z+
Mp2edOZ4Evo6U7DAMCvPorSGi8cESa9esDUVPazzOmStPhoqjN7RZzTT078kHaLI0x887zbtSAGG
HA+EeNChh0NLBJKBKO1GyoHocpus06FqqVmths49X0d2+2GIsZxJcGcEz7O9rNv+p4UuH0zyjQ4X
9mtmfVSluPlgdiI71DpBbh4EfQObjvl9HpYxYGwWXJUD7CWelD2STSRRWPgxz1cATh8xK6anDcuK
3xzYMrWdRrhz7HKv/P4o8a/VbG/tpnSgO2zOhfEfc84NtfyDG99o+9TBPELdr9aJD3l2dxVDvGnn
uYwZbjMHdFsXLSn3/52rdbe5bf4dLVIehtWACNWFNwXwmgIPag7vnWrCSZ8DaY/Rp5NyXkxgXLDI
zV/NH55QDzTi46j//rFg7mi3bWEo9+8U/RFN6h8q/DnKj4b/LnDMqVM62FwBH48Ilnc9lTfEaTGJ
9mIAVneoGjJFFPur6vyO0qt8ObYHhmEMZ8NY7O9wRKy+XJxlVpE2Fl98fiDTe25yBtfJ4xAZ8vbD
EhvcItun4GOwyMz+23uUGm75E2DbeaCiwh9GE8pFnHFIRtFrL4EHRPngRAZ5ve6xP33ejH0GvpK8
aV89TnEC878klB8vP29A46G21GF3HN3TSvhRfBYO7JBoQfwelyRgr+LN27r3iYeQvHKj/BQf6IKJ
jV4tMsYOXUJ4lNV4XG/MJhsaAgSBDdQ3fyppF4BDp2qjjmNAIIEdQFFK2lmvX2ge3/DbWbNz2lvf
W/Fk/qPju2pIqWyQZEq0/JKs3ws0UtIiLAsdKdY6OxlcAITKsIOcerZd3QnyFiwUs+lYbnSw44od
ICuD/54gewC4W9uzqOey1t022WLjp4RVvJMo7g6C2vjKxzL1H+wrj46usdMBjg7BCzcz5+9inCM5
0VSRYqwNEl9nQla6yAoIzkj8QB+6NZRnZ1qu9pSpz6cAtZKszAkfUKq64pxDjjIMmTtAv2hXb96S
fJrDx1QbPHM3kpfLrR3RFLfevoIezX4CMlM2rKwoi5oqLszVWK2+Jz5Gzm7uWeyf/EqosOaKtZKu
m2L1fASRX7viM50eb7376d1LOx9BR3g+LxSAirajEusgA5/Kiww2649fG1sdyMQGN0MHa7IYRyf8
P/8eHAVnrQ+wAXx9kOnZrhx7ihmjDkK1JsZDLG+1EB6X8zOflxjxmWWt5XaUxnOc+cNVITk+VHyi
qTjnh3vAjt3o/uBi0xsYFRt/QtsEGxJ+wuSEKwyAuJkJ/8YkrENvcSkk6gMJyega46H2b/PopzX7
kHj8JLT4It40NjYeQTBWKWEOkJ9marqnQk8uUiU2XCu+VdTxJPuRKFFmrLmvTqtW1ijiAGvVfjDq
+vjGenmm2+bgQDBQLCAFfn40cMbcmlvRWbZbxl8f4A2UjODevTmgl+0phJvNDduDYX+yTtcgBrZG
soPKa2wTLku7Xq5j2CjkL+ULy1DbwBsxBR01QmQu5yRrByeKkT0ed+vl/8QjI5Hm3KmxrKVSZahN
3WiSlLb92pySgiJTKzl0jDet40jH4y+ex8SNTdUi/P6WhOpW4nXFuM1gnsyczRNtNd0xh5K9buMj
4Tdu9xxGW5N6843j+87svLquzqiSY7Pv/aFVNcQrhAqPu9pCoSDF+TNAQ/pmgcUc/lfE3Xvr3PD8
nFz3uxvZv/VaCe0Wkn3AOfy8HTWLnyVbXc9MQQ6hA4sF/Z/0iKlwum+sjdbuumhqyhFropqehCkd
/UKZaBQL08dorqjY7iGoIzffrknonnEHGV2Y77rQ+W4PjnlBcBZg5cU7zO/yzyvZHViPFhSz13VE
D8ArBWavoUEhwUSNlLSSxC6csE9QpaemNhQaMGY8cpKqKNRJpJFnXH4rTohcUNaSHJTRY/bDoi2m
gvPju296p6jkAaRHeFZi1EMqTzYuV8kI+2fKBhWEqmQTags5llQxg8gWr0jc6xa81MdVLxbeMfpx
b9dpP1Uit30zdgncF8BYnrLOkb7LyXh6yJb6WuVjWJmZJCAxwkMjXk5l/26+Bs1TUuCEpkA8ms38
i92VB6HhO73WevmY6EHZdv2owOGJxZB/Ui/0q9H7QkGiSQtgbQPlrqFJ8U4doh82ujIrsOr3Q4ue
CqPqAmYgJX72tMk3g4tUAVZXM84EPZskHsUGJiP+I5wgxmCZbOiUJDBwd36z8ccJtlbPm1ZbJOfd
qhK2B4URxyLIULb7+v6AgAQ+ryOnWCT3BEhthCztF7ZKoN/Cz0326BcaLEDrt32ur18dxZAl6I/K
p/cLxF6/17UExnU7Lsa5e0VgyBxefXRceZUioKUEWnXptH6BuMTW4EpNblo/5kHOOgx+SaJRTmWQ
oE0nMuyfxrzGJO8HEiVEfiJlGwPNNmkcjGx1LG9M4IxLmj66LsFv9onEH1u4UWTSldtlq4z4Zeb7
PVV/yysfQW3zSGwDlxgwlpexXR0XygPKOxR6CPmlo3XXEa0I7zTxmsYnUce6QF25eQXODMzbV2tH
2ltzDa4c74F3jzb5CipzIYNnihLcwWuWqu5T2rhDgdzdFPoJdROf30lgPmenCTOsBLD6bmF8XlS8
mjShFRs81pwUvhZEHmgqzfpmeesNqdCVes5eV+qneTOLN9rcE0D7G+PotNV6dYh5+8OIUfCwI5yR
c6bFnAG6ZKn2BF1aRSdiELMZrlofGRS0YMMc6raYzXjHwol8G0Twp9fHbvh0SKddQPGN99YO5Ue1
efH1qbQwywDgBicIh90cgwkkuOhKWH5jA8Q2Rda48v8upeLefca4ywwEu6VET6TCTXcPeEIHL+rV
3/MTUPLUvwHymaUFM2LxdbIQD0VT5JHo1EG9ZTozgh00xxVNGvZFEdmeIpp5I13uJQDlcsl3XQqm
Zd0lAHIgWAlo8ndkzKwgaoAkgjho55UncT/HR1XnAlMvdNVuy85y8TiMZpInqIw5I0qF4IwtntSM
HsX6vnGW+N2jkNe0582TamgaiIz2J1yhTR5ed7Y3IK+6PVuBeGqJUCdEuLTUQlQP27H74uBkngMx
ZNgMEfktZ6ZQZISov5M7EDg09BNCtuCGgrRbedb7XjR4Y9n+hMB+xFFvOTtBu07M1g8eUrjHShxl
0BEYzNEAMXlI/MKtMrNjLCAYkHx6qUXdvYJ1Ss2lcv4GBLLVEO+6DJxWXmsQCyCNmCmy2mAbjqOQ
wVrR4s+plXSJV1JtTKXqHByLvpaczc6O+HmHudT+BsPZAV5MJQ3AU+gpe+FIXIAwXUUvxLbgTcCg
qaFrPypQJPzyqALaoYKIm55iVp4TAd4G5ABaBQF2TP2xin7n5zUv62XsCu6y9cOvi+QI+zLA1UHD
G6PEdOF+PGPLWKevbxReaTXpuXIK7IiPdMKDMBpvyroFRmN9oNaqlkutow1W+RZaXDabauB3qrRJ
r+mA4/hjfPfEpPx7d+uU8hCrdJZmnh5awqKMoRmjMLyZ+lZaTCl48dZ790jEx4IoGroi47q3hJ74
YnH/q7UEx4f0X7KRosTpeAdDFvy4vk47V4lrVVDZka9zV0r6QyAMMTXHw6NIEbTQaqpesv/VLD4r
+nXJ1zqYqHIrjV69+Xf+NoBfIcreu86b1mepDPYnQ7OYbGf+6C5fqjw0GIvN7I/1G4eRDyFHBLts
GHT3lJQ6fAHFaSt9MAzZLSWW/pxYOVxWOcFEcZB3BMFO0DDXpUioeAtelvcjs3S8LEj+4B28Gpm1
7SPi0T9bD6goNt+CK6SEdU2xbKYBnsu4ZsrxNyQYBoN4Y5/oyMG1Qo69NfZVJzj6NMsilyXewBTz
WZuCnhdkBHxDjfE2l6VKjZ4m8zVIYaMnd7TnJU9rn+UupzVCm/6ZsYeBskAFsLwEwWHMbZs+pnr7
jKcW4OwhclE2ScAhS3Pegjq5s0GzyTtEnEPPtlYhVqAUbaF/nIR39wtGGmqP5QcOzGD2hUBk3oMd
GVSqglKFKvMHSGFC5nxy/33YOasUEo4ksW3xTDBgytlJc159WxqJ2dX61IW8DaooPhbcd97Upd+e
UMiPfh6/28k+b2168Pfm7t4wYtGxfqNOA8zx+fdpHVawYefdHZldQXg4/DlHbQ3VwUg4ky7wsCNB
AVv9PSJ+OuCEoRczYY/pLFgb0TX+s/pWwpP/hmDR6DNWhGCfhHy1NfEdeXrNkpTJOLTpuW5X/f31
NzIhdMdTvxfqrNyWOSChH2KVM5bChjXIFf313xfspSySe6r974ZHGUyIVvcMoCcjm/x9jk+/SVTe
8OY6SHE48nBwl80hIlj2mKDV4mUnXT35nEqXVpzib02bqum5SlHfjSbxCQjPzYKXfzBPkt1gTwAv
iX2EQubkuCTeBrD7EWGJ9gLkaieLZxxedzZXLN/sZg+xnVNw+Vn4iOjXRbsoQqhI1spYkcZ5ScrB
gF8UJpzVD5HIoqwch2nro/xjH/7/ryaXGQ4oeNgchgCFlagio8vzGXUHBLgJAdeU3dKAv8AymTOQ
IA7VOiXvlNq6Oca3dB7+Y5lHwBUbd1Qsan26U2pTJv1fCmv42OvojVpdF4S4zR+uUTImWgI64G9S
zIwDhNbPZLo0JvEBjDvT79C0XnzNH4FkOxlJwhiWNPKpNnmQv8r9g3dK0EGUbthvtsAhR2K7pSF9
uoja0HUCzXf7hLIKZfahF5YvpSLzxXvB2gDrWUSUJcAPN83hXOHZn50mPqNAIhItzZRxJybviCqN
E49GqsO2TJXVC0jbL8B6BZf9k8Soj1enlMNvj7KPphce56SE6pY+mQrT0OEw9zjzPjmAGdGILbXH
WyClgLwXuDx+59KZ7sey38fGKZeVhGgzIC/gh6ypPCC1Va9nowKf6zjGclP7ab9F1Xqs7Wdn7MIg
Ki5C5cxDuIoVuxYyX3NrsVKr7HgGhw1c7Xt8uyo1XFSPQfbKW2mI9qxv0bEKh1g10Ma5mKg0vZAA
oPLsB/lBUBWCRSGMoCRLh1wfv7W/4enB6926K1xwLkQvk4yIT5JtCxIByniELB8I5LEtCGEltZkb
+jHnSAU/OXd3LupbQawaDWg2P/6lygzfjB7bGpF86oZLnEnDOdvTr9IKvuU+Nl4EUlr1BhIcGqcF
pORVrWfVDfxyhZtvBeZ6MPMl+6pa7KgJIXsce3KnC/GrdZ+cRFRPqOWIDel4Lgi8vgjox3Ec6N3N
tz4MtMIwBctJECO16a8AB7C3nCbOCbWIbQOeispUOMdThZnk2MS6eXmczl/mCQNZr6cDHT5jpjYA
wpWcRDAJXKWVArTx2ZOCCym1eOEcR+aTajFk0nJqlOpfviuN/5VBTKpriUl/8rJMLUbelVPB/BSk
lFTJiQdIuFlx7cTlysrbdcMbucxGYwFXuQ3LYCUGf3skovV9iauqwpSEIQDRjvaELkIujU7Wy9qv
Nne+YMrf84PeR9pO8P3qi60v33jBJeyLXZy23iD3BeZHCUZ/SOC+zdv76KpzC3bbv0os7OA1mKJo
gF/s7JW0dGxqnbsQ0jGLCOXNwqDAISfGKsuU6TCXEOrXQUFyNJ07lGOBoUyZnwDmExyde3GcVVdI
VSPzCY+dFSkkSDoF+DUa9uh9F5wDjsp32EZcpqORQwWUYJkOl8KD5tzEq1NrWm7w7xiEWFxvzQHg
FbSaclgSIBuc24fpNWyeM+46jiO/3yUwH1NDvsJAlF7yjShP6v5x/6R/FurAVRErmw2D24dQmfoo
dWSaQRQd/T9xk6C5vvfnMvXiijScNyYamxizLxbSe5reSpYLlcp790pjHmF3mS3UH4n3X098T8Le
Z9AW/9C+F7jLboSiaurdPsPxG4TVbIesGudZnDUVR8uQUk2leLl0kI4oK8hoKqyiyKKI5MCaV9P7
CWkWo3xoDAmENLxhMyuJBQ2TQdNNdi/MbX43Q2ToPetzDrTVNaeIlAq5L+Xnbpi6OBccJLK/ypTT
ajcewqi4kG0ed4NdxaPBmtTftzB1klza52TjNkBakla3eE2X5mVCwauFFVavcygJjaUKvk0oHaOE
acOU0FTTTLKZS57yP4dEr5yB9/xUXeIgGucOd3vD3UejMmDPZuTPw1Jj+JBmaQwSMt/ap5DAoG9D
ZGROmLTnPgjcQGV2BbxScpFNdJIDOnCVbM3D/KlCm5n/aW07OFcqI9p36O9+2oXl6w3HAJtkOHHl
HbaWMsTbocze2+9vns/jWcIIreNdqT14x0JkCN/bpyYFlIs/1EwMNLctfNA/Z/7uwg0/CM+NLmsd
2D5yYbyKfGlJGpQhVN4ES9SqyorUNXIxOepIPNbGKVZzQhSFOYtoBLXNBaRUTl3eEzgVD5LfSx+L
LXfCKukUkEDJrK1jzWrEXvzdOPhtQUBgdChDh33rLzjrhnCxbl7suKYJNGifeG4OJbheOeLxw1OS
ErJCA0FwPjph/vkHHUfN9h9hySPaoACCEbDj+To3w+WJ0lFzwGjvpo6orx4yD/F2mzVrn2z3FXNk
8spejOB2rrDEzg2tmlQzvLZjMVXMxYcnw5cXQHHIwSx4TLl36vLXSmPm+8X8fX47R/SLnHsVHUOH
5vuDnhVQIEn7TmT2N+gmcoXDx9mpjqMQq9cqNS9CL14GPZXF04zQhljkdBYjvuW8t53Nq9uySFk7
sln8RyKNf8bkBrQ7s3t+TBviNDXOqeCMewuhgaJYEW//2WgHLoGSG+DH3zxNMm3O75pBTOz7BfuP
lOS32K0RbkMP+DXhbUAW++nHoy8NWi8xPBJ7drOAo0iCewW3hWJjCz+tiT52+WBhd1nfrAy2iKFN
Xhe7kfAFNjFTHqPaF8UuEmFtwn+UTRjco4eN6R8qPnQzrLrg9rs7Ioh9muJbRVcICsoNw3GjX1ar
bp6nrcNh+iIoU7RCe5YU23JuW+FRhkZcNvhmAxl2Uprbd/2j0NzYaiQZUibrHR+EuoQsuqWFle4X
8YUsInjlIN8kG3+7zda9V6t3kQXRGmAyzY9oqlHNap905eFv9EXMlf4EiNBANSguOXVtj0Wd1sMx
983g+K6rwOxW28n89bpVC/lrJSL/bOJKwYN5wWrXI1Fh1tE1vZertdGx+z8irM9Nf2ysz22xswZ1
cVgJcOvNCdDfSfOLBuCTB421n5Kcog2e7IffKUTg9q7jFW2OMJ5Y2hSQOeiKC6Owt47LLm1qeA3e
vdc271rHny7xWic+PAIJBbhODOv4WgG9xGrwEWUVSwctyZvFSgh/ng07Decx0pq3YF7RsmqqJmX/
pQbXVOhWNg0mAtM72AWKReQuavemiQLajHRyps4I5p3eCjP1+9HAz1YboY3VhV6CSDiGx8iuzy9r
1wsLcZAiBeDjq5Z002gC0XR9QX7Yd1pN0PYVjdpeb+kuklK3N16BIpHweVlxRmhbq4kCWOx43v2G
hO4sLs/9CrCPG0Dm3sK8ytUq3FAItGEF1T0Cx1FdOw0irf6GVGPuY5sLfzNplbsM14CXmRXH1nxx
13GSUCr+X6NpGHkQBgWshsxzvGr7+k/HjUpac8ClW2vMRTeNyggFne4igCr+abKuYJ0Ac1sx6HOM
6of5yl80qBN/h7dswlN4mtQ12QZo3wrxzJ9bSKXqk8F55mSRXcZjtzjGuXsPEb5mEzIUG9X2jp1q
X/FT1/GXIZJmGTlu754iBm9Y2bVt8SxxgVCzg0D1c1G8C+YR+ZhdUsKbZvxG0Gv00CekR/RYOywZ
wMS0R8raz6YGxl9cxHH5vJ41X97i+8qrCYxsfiuIpshujW6DGNl4nqusfXIOC18n0uM9s0jJue5F
RJzQduDtUQ78RLkY0rQdQAnGAtxOos216urEP+L4wdU3U+uNRllnlxkD3SiL80jvVMJT6uNym0ar
weKt9yg+hwwMvA2cP+PAsc0A96mmlA1c/6JnbGJZRBy/lF9tTJaHhsiRZxqP4mM5y4IXFrJqkLJr
bTXkb+wElrJbNlEHjUL5LAzd3KgQTmJkuHer3qYg4E9gyu6ykReCzT668RDn22StjblTXom2104a
eR430F1wOapSTl1yJBjMSVNoI9lnYHRSDZ0TxeIkM9zac/AOdItCE+4KyN3ifOvDUTrumc4oKGI7
Zlnhk2Q7R1qN6nEH1CASEsFdALm8hbv2w3ESfu4UIO7paVvsXv4tHTfLLsBhT4MkDxkeLirfvfdc
isRCb9xQQbwSInOBMsSrwUpX4zaOoYzors7lpDEW89glrcMOJniGBLj/S11/kohlbqg/RX2umDvY
zajRYsY+05rY1K67y8lhYriGJ1Fmy5t4QdsNF7HkkjPjnoACjHuCDSxbUfpCkFt/bRcxYwQx+IY4
7LsDgcJ7cBL0SMHYvM0DJKbrDi+CXl9yu7a9PxOdhARD+gZmuk9GHRIEk93NoNLc5DBsgavd/gr6
gbuwUne9p0VbKqYIqZWLdHMf20y65WEcPKBGfJoq1uDC5JZjNBOBdr55cbXbY00HDTexBDQrCnwm
u2W0+3/NvkpM5BssyF6mpVFSic2UyFodeVXrNO3rReMzrjF8MLfO73tdE8VP2g0Pom7Zf8+Xpni7
R7/EH0NdvePipPRPQQc4vbJmakxif8C2onGxT9uAiJuh1xWsBEhc/DfwYvnc4qEJ4/cAlXPV3wkN
bQh3d7ecAgez+q7xZkUdqgbhD5sIWoNaX0DhptB2P8F10g7W+m9y1lC1WWzqR53Zj2EeE/ZIuAGJ
azdBBzPBd3Ny9uNcYJCMY4AxaLYONEz6a5wvjIcsyroEldYGiytRbgqB+q2+C6cXKLthngpQtMOP
POB4K7zatstryLxay6GyBA55PAxy0RVLcxcf4v40rS5yEFOf81PVu+fQhp7cTV8gyUenWpiExyTN
x7GfHtPHTMNXHc8sh8ndNs8EK5/s8dkUmiC2m1KHfMNJgEwfFvn274vQLxwoIWpKPecXeL9kmFVX
c8453FrogGuuXdL1hmM5zzBp3caRSNwzAN020sK9seo2DtX+ZAfRjUQ7MzEl/MMbeLUIW6bNURBK
nZdCzn4vJJLgCy+jnKz+assYaeBG0+3oqSTJf6k/LpcvHSFWPTf3m6QNThGklYL2VfDc8xYqz5gf
KIeqTmRfpLI9Q6bvN1nfv6QKajSeV8QRxcOLhxfLO6L6nPiFnE5ChH/Tn5gkQ2MkNwgrp8in61sq
M3BksTLS+5WgISFm3+KchJD/mtexI/xiD7BwNO7Jo4Syz990E7VxzOfX5do7t32W0cErdmznsZYF
hITGhXDv0V7yPDQ0LrQ4eXq5sa7lW1GPRxEx7Ku1MEGKP/T5Fmo2JHXQ3Hxr9RAe3v5JjJYDFJQM
3TslVCEmd5kSwrkORDyRchA79fuU3jsxQcJqxf2VfX2nOzz8vb5uIIBejr6v4kryJHeFSHBERpuh
D86MBjxPAt46I80jZ0XVx0yftIMzDUwQtdHe11XJBAyyVaySIc7WdybkUJAhd7VZjPCYbEEwwGs3
wb4ffaYL1qOV5jsv5g9OmfS0ICVvlF+rN1ypEbuVMg2pJf2LVhbbHBFeBNojYwKZGsXIPwVfDI14
r4tN3us5qTd4dPrac6dyHAGNLHSmi4sYf4FoPCakCMSfYPanF+YccLJhz2ecDZDASlSwU2x5mhmk
kjSSkW15b1dOhPFbTXx+3wxcuI/thU0fBWbshU6sv/7NEyzJ6rJZam4vFx1rwaWWx2h+u5sNa7eV
W1kD7jdKHihADL8VZHF9txKZQ2ibB06JtS38SdK5o0DCHq8zHwysMs9XFj22jSDVQVQdT/1x0g3j
Ny9zAIAcVMg1R+i359lvKrfDe85rwBLuAAXEcxs8ZPrhV+eGOVEl+37T8BqUmgI73HsHxziIdZuB
qUeTB3cz0652hgiT/hUG9WLN4FVPQe78pChhWkVwyBqqgI7RXmZQgQDN37b6nyWSCjj212CWqCo6
9av/krMLvCPOlMzyN0Q+IdTWXFtHmQo9nstn2642458PHmXy51FG2INwQywEeAE2RnqSeIT8wwRk
dBwG0TztCt1psjK4H/EbFj0g0fzKRy4YLzW4CR9A1XvhxpqrhiUtlPNpxzAtrrWq/bp9qFAHYgx2
gyx7Pk0K7grFTASV0+yvBAOL9+EE4XnFYF9NWBxJdRyuT8aV+gbzGIQZJVQnXGB3iOCcsUOXccV+
+ja+nDsQP7RJAb6pG4Ejurssw9eSlsj9kB1+OoiRcbZnhfsujrI1Ssx8h30ZrZbKAx/e57VNkmO1
bq11CupEokzsfrF8lO7OOtpCp+7yt9mdeYgmLoSwiE95ZLeYf8vSmZXVhqa4FHpHj47Ww86amYmc
54cdLrbo/NvmdvUnMygyx42JgMq9OJaeObOi6r6ETQf+owyAIRDCEMC5RrUKRl+WeoWIK95ptBqN
HPu1yOYa6aKzgrm5BJHw8qTm8cNnd/+V5QfoFIAYc0ycfkrb61oTTtwC6YoPD/gMqfTINetqJ2IJ
GwLtfqceJC1fp1+xOL9NZ1b3QqRhBPpibSyQ5WgAhEWiIb5SwTSy5tgcMZuC5Q4lHOvow96bU6NQ
mLzyoiw4cJBrIZ6m5We0qlmC4dbp36nqJ8FHRNmd7elQeYhASd0znH/f5aeeJIW3fp2y1cSV7keu
YWsdZfxByZAOCZRFwoQ6nA8dWrT15uA1dvW3/UJ3R2mzSmLFIV28Fia4ZNkE9mSbJAsRrM5vr2Gq
P2f6FOd9IigqBWGh56laMzNU4cE/vWozXQiEgCfmLpEiwnm07K6Rxt+b7P67DlB6Jm1p06UXvtBL
fzhREXA8LoE1XX0ivt9+yyBNMsr76D9SHhi0ipvL4836sFqE91RGLVpkOcGycQ/3Y7nuINuwP4ho
d2Ptd2/GP1VCwDf69+Dm3rZ5jpyVD4r9ZFo51MAKhIlk1n6RAzTcGlTs0ut9kyTMPa6IvdFQ4LDD
xwIUFm8TIW+EmjcRlLTSrkMRkGEiTQwcHhsrjJOsdmnQ4BzgJKOUfudZPAiDVa5zyIDBe+skCZlf
BDxIhiqh51TyEHpHrxgP1UVkUvWy+vXvzWY8ouD2i2BxiXV+wt/Sie5x/39vFOCssepg57a3TDbk
NFDRoK5nqFMdKh38qNanexxnEkmZT37+uq5P7/j9lKeDEgRGaKlDlYzL2vQDpgWW7BM8KHt4QbkK
OfIMi5oI29wuJOnQXRwDVWL8B+qbIGrNlzLXoxCpN8DByXZfb9QoOKFKXQtWYRBoCNb94GhP+qa+
aH96XAXh3rN92DrLXI5fEpJSFrmTFlGPIt/w57FuGRFwwbJGywlP6cBHMMbwR6I95P2uUAhIw7Eh
tHnI3SEyodTr65815z8Q0FfQpdjgvwW5tKPxE5KRbZXjv2huUQGw/y2iSoNRGnfkBo4//dCpfxtX
liIFhP9uAY3GXnonlUFrejpFmNgpenSEmWpdm7SWNKsEaE+5vblMVUIm6nqd9eYSqTMA2TF6Gb2Y
CE8BQolDgAtmZ4w5BjrnLV4KLNJerTq6x2V2JBjZj++sIwX59t3thKN0ekgtcBRD3NbeADJSZrRA
IAqGtEk55YWHkI5VbaKMk+jUCiK5NVeri9UbSqnzIvE+K7PqRrgVjxcYBrUbZx68AyJzoSC3cJNm
sJJ9uPhUYPPb9yKxlY7Nz8BpCVVTC2BK04youfUrL2NPI9IpE0JNPr7KmLjyCWM1QmpzL9KXuULq
oE3+T0XEsWbMyfNp/isHkEZpgghE8riNJ4Woi9avoBcR+xLO3pR15UaTaJOGohh9V5/5HfTfT7ZY
AJQTu/loKiAOjVVYkFfnhAuD9WC9XDVwWf4VSdV6i3q523nxpTaf5As+zAWhYLGSMfdycY6T4R3k
fyd8v2qrIOkyCLNXWWoucOMCtTyH36Mw3F/wl6ScHVHN+6jy27aZcQAHud1AclIhojr2U6R3IbSn
5lOPsIdaOWNYyFGbj8jI4L6SygnS1xaIPpRPD7mznUqOwJVOxP5IRLQYAu/Lra/R2RfgsWvizcwL
gBwyIJAUoDM3rp4vOliahcQTMqb/S2VbeMNxw/0WV/6VFe70iNwKoA1kWfNhDJJ5oD86MGzTeyqQ
R/RNVMOS5Ge3H0ESe5ZnM8GojfIM6xQTqenbL25qRVEjHZPspj173RDTV5VU+lvuElEBYCWi/5iR
qEUYjcn4vfT1kywlBvdH3LDWYTuJsu5NknUJVTdLEzXhC3jjJMdQVzNm5sHPy307D1XUCEKwRVqh
pMjga4CYvzCQfrgjofXm9Ho5Y5EybkXe7tmWb6PkMZXsIB7KuWbfYsHe46pE4ta6hntFpobvCc/z
G1Nkg24Fzlqniry2HqdP8V6iRt0jg/GTn0mSjjpf3iI9k9Bw81hKwWNW7SgsKH9eYZ/Zd/P2O8H9
5xdXDNXtQ90jtCU/yLy5U3YDNeL3yLROheIot8XWqKIc1FcjNFFc+Ty8ac771ZpWlhVUc+k6+Ko2
RPt2di/OtyFTGN4C1qAQalUr45MKqgAxUlD3vUw8FWoDKm4hIkKe3Rq2xLV5PjEnuU/jvRksI872
TdlXVIU2YvefzaEcGOoCwO7ToUAbWqXyTJbuWVfg6ZcTH1m2jNQGsaqGcLSZGEl6wO7rb7+wkc5a
ofOZycqnHEM6yu0ZVQunkUl8PtEV9V11wGCIsWIaS2TVAvZTVI3OJqnOhkw6iqa/SvHRfMfYZlOK
SPOj1UFsy1OnpStfpcHh2iUXySnSp5qFgmHkjIsgtneYEb2KeFDyUiiMIw94yokh8erSOAZxTf9b
JEBWLCQjk6Ul/bVbxaK7lJWc6Dzjw8Nj3F1SGnDV9A5BTL0mAzGOWVp5nrR9N3UZLDhHc57RfxXx
y3ZKKdyakJeT9kttgAdbFUMEbGWIkodu05gx+NWxvfEnHCyISYVsuxqoUZxib7PoHBOAmVZ4ftLc
wRPwkb8WlaHJaIi4RrP9GIQMRQKUeXHbAMNYFdG2KoJRFE4yTrFfwcmsCD/D3eKFOeWYjQEHs41I
ywzxt8+bCkMLUeMv+t7vXHzEIy/t/dhUsCw7f8S5eNc9JdsGDDv+65CglNYipZrc4ZeMG0ToamRo
oLqrbm4P5LUb+N3zH5nx7XbnGWkoX7er3+t3fZdYFtr7EhklZnD6OCtLN513ugmbIB19K45ElOqJ
0pUGi/29huJPpSpr/HOXGeDDJdw9FF9wA2eyCbxZ91drEJiFbHICN3lhZGI4eughLLedcBkP7brS
gLkBDBeMfgsP7NcxP7puKajdGALgWqA+bbZ/GpipG1jMSci0o2F0PAF+/jUDJnOjwx+ts3oL2azY
3U1S4QACvvgGsqzJJXoOvb/xkvcDmCQCbMUGzv3iZKdH0iBsGRz5QLiBoIv2T7iyLGOO/evJvzAI
ZL8ClierBHbZgt/HOpbjv077O/aD9pIwvdbQKsHmLP62IlMRvqrmXP5RxyJt+HR8/00G2mQZgPrr
VufwbFdoQlZbm1Fkwel7qYVv2wMAWjLiIwt/nfKDs9bOYQQIIwW/Uf+Tu6zJDKSNCIFAT0G79kFK
Wr1H8mgmzHno0uRlfe3CBvJs6AXkVI3OG9mbybRbX5K7qCWV3SWyTxMVk2lC8cx4Jibz+n393sCy
643+MNSojMmJVEygSBQmoM8LS5A3aAzLLtS1w0IVd6cg0q6OrOFDqbjBm7CkOtFGFfKImEwzzNmC
e3nAVqdm5dGdZ+x6/65En9XAN9HIiD6alVrt1VPeyGaCKvY+c9yDkxLaEdHLY43XwglR3DL6e11y
6giIzV44i8OVToKOoZ1jjVxxtls/Whqn8BEuTM+HJ8G2nXBT0Tu4G+q1/7/gEFUbV9DYDRL/UvFS
RdXcVPIoxdmgkeNMVYe1f+aLqiYfLo6+QXJ0DimLq5bkvYCtKJLQQYX8u2fQB6mZZcEJzWBoWHc5
kVEYtZoDcrBIYwDYnu4DgcYWJZlcadG03i+RJ0OTLIDD320yawU3iaCAqziXWA4hFZ0clr3Iszyt
12L9L+e/snq7MV4+D2sMYgVgusqtXTxl5L5ISnZdDQr/lbsz2YBQGjM/EzbCiYtL+K9/z+xyVQ6Y
W/JjOsMvvI6PqSKS6iULxmMV6zpiCFQSj+Ri6eT+jG+vBDvdZaBPZmH7Z3eQjwEzKHMpevAutKMj
QRPrh71KvrHnBOOcuIUFilDyonv5FV7aSkC91Zbn82EmABBags2UwBliQXMFKeu90mH8XEeBE5Cz
Hkchf5/rnZxpr6xftOgozbJUpXwydLTncz7uxe+OQC1NOe/BkiEz47WAsIMiWlQzjAAIZgWkLaua
ZMkq8deq1sLu93izYxAkrupH9t7SAtmakETdNnYnLo4yunfwWEkM9vLeQpUGmULbV1ZRuFqJgWql
RuzXjJOdnLvSYDJ+Dy6+qiu1Wc8PRQyANcYwnNbu4LnFwNK3w8CndRLdMpI7PjjSxEmujroHuqEU
SfSc2REM3TO0p2Dn7M/GBwGpfNSi3VTq06bZKJprIz5IG3aPlhOcC/8zZL7yIwJpD7f0xdSQkNhU
GPPP5b5AK9uHOq8gvWE5X5HxrxnKballlCHUHMzSVD9Rrk4JdFe0Ezx6BZWKgin+hpP7ej/LjiMx
PM4tFKWhJqH9AQtpx52rggKAYRCnZbd35gIiTezBOGknsmW4WDWQXIqOL0x6BfH/2S5hPDV4U03O
9ZliEh0Y0fctXR3UhxnFQMP4K7OEdh2TucQh3XkMkMldGsRatds0u7wj+2cfP6TLyD67pLWTPrgb
UfWPFbOkZhKcoVFv1BUuQMSCOeOPtX2ErCfUqmv195QFrA6J1opTfpC/owMJsjw0oUpcvyXt8t6s
W6vIvHNorSh3019iR3g0coDhsRe1udITM4eJEAgcyx/epbY2bjrGmnh9kVynSu5/BIVyQk5CWW1c
Qb5hgAJ2N9E2Nj3P80E9zqhl/Zd7pzMIeY4VlFjBa4lwqU/K7xbFxfnlhRJofaTqBeCNsBMrjk1u
CpGpBZ2094Va92HSE2GjTUsP8fLfVJtbUws8w6Sy/a8Jxn8MzgEXj1mYNMW0yrX8ntAJsxx8E2zR
QRPEROMFzwT2j67iqvnfwOQooEld4WKbf9D2iC+Oayqbt5VhObncU629SiklJ1kJep1BWB+brUcl
49vuXsuIo+uVsBUQr4v2FN2EKTTv00rh6mgkNV5Dhp7SvgoLSsFeq3k9e72iwKlRgHQqjr6oElCH
wz/lkSj2yFcRFjmdjQzZn0l1im0GkM+L4YmAKZaJfSEd4HQi+avYy4xgJjtvqo4nPngPoPJS13/b
1gOll1CK0RYRfd9y4Y4BQlp3avedeLDLo0wLUNd1qn42sX+606/Fyi1BNGnMcxuUarzGZrcecAmn
dblwCfzrlmoWqmfEyH5CXNjoYUmFY2AZKqSoSPS3+nz4kPRkvH2IE8zxqCUqLD0iOk4NSXC9wiKv
1KOum1fBgfIC9u+L0jIVXXl+I5RlTePCGogaz0un6Mek5/AYIOtvsc1HEhk+VmXZE/zu9S+hXo+s
NrQSoMAtXHaf58cTuboSKOb+7mMoCGfwWCLobJsc1BLtsuKpDJ7M1g6caS4nmoKzHeZI7jOX2Ypj
NgHaw8HIIYXFTLfcv4n9HK2Kab3ag4LTz58HUt4RyaKhgGBG0+6+KGHHKnUc0yZjs5sKaL+mU3B0
O8jYPqj0SlNROYYZmdNvoe06L2IW1o84RfHXj+oVlA071N5O6VoTvmZNG3zZBZfdn4NSZiaZra0R
oj6nvtLLwjjtuFn6ptaRj0UXZQPOvSZerwnMpVpdJ3rVEyAUSawp87sWOF1uoqrA0BD9+cN6Vmvn
iiqi7Fq2F0oHiRqtzSCLUciwj2kl+ovFqslINRoHDMzKgNxgkyQO4JK1C5oSfWWotMzfdeASCYYN
dBJHY3vABf/LkdER8il2xlQkgDV7lzKA+rmTcrI3oCq+21pIEEmq0AGGw1g4IathWbm9JsVKqUNi
pQBXj9Vwzfkj/ACl1PATKSL4j5PRcIeX3W5kE8NoZy6fNwIdIq34jE0U0HKwtUjVe8NhGENCRI7T
DRNxvixI0I0Q9kQHgYlWNm6Er2tpvhGePJb7A+9O3SWcBiTXuyLF78+44gHRRzm4C5gn7Soz3Pkk
VulujLLuDwpVw9/dsW0ec714j8e0tb0wUbmeYODqVZR/oLlvx6jaYJBGkeNNPM0YYwLtO/qWq3eN
ASv83ZU1Yxqw4sIBAhNpxUtSDjHpPN1npRtUqmy3FQ/0R0+ygEBcKaxSsKEPsvV3LlVmBGaWAUJ4
0JafBwUnfOrsI7bIU16M9pako5bprgpGi1Dqujvdyck3XZ9eOWX/m4LDRyW9ma68uF8f7TVV9E70
1PcNrcbvjHzoRNDqgvMby95yWAr3d2A0lUGYLaQgJ8JSAtr1NESk5iv8AnJsi8Jh+jFDvoDvIRTK
u13vYDy4QtYPC/hX4yxGY9v9eXZqkQzpIeA+0z4vglmRjYo6HZQeDTAyT1PZwrDfo6n1/LgQLKvt
9fQWRfyq/qaaau6NvD1s065Z40Z8P4f8GimFOXENHKlwHEqIw9rME3BtmZEtY6zow28fEyRXKMAz
FvvXVTFUogxBaBjdlYrYtBX6zE+k/tKNjlmCnziRjFr+/oT1HuYLGQI/nXC6AoaCFMFQAWTzzgQ4
XTA3UJqUCKbBy6rhMGK0+xza0LD661cujD31FQGt4tFze5T4hgjV7dldERi9cbrysPzkcMefRRRC
VwDYsEo7ngq/9zbZx5F+EGmaoRDNd4RYcJc491/tXi2ILJ5rBtzOki2urzFqyFH/oIMc1AelMaPF
DwmZnDUTAOsp3rJ1hjAqPQdmso2TyOP1hwQAFGqpV7JZcvdsK0+NhY9dbUZiA0Q8FaBfk8IsK6dX
PhKYoANOVTFNbP8JmXBBmnjgoLOaEAMXAsWMj9oUKHM0PhO/OKi0jnxGQHPBJPRK8UaxOmJvu233
W/rFfyVHBAiGrvjWkwcN/LjVNGZzwtK0MsgS/NgI+rcLNMVYYvCdxnzqP8cmdFnsDWcAx0dZbtvX
Eueqa9oluKzcM4MOUVOmv97POjuWKHfw9FO757onjxX767gGueiN0hE/MlN+bXcZKJtAevhQO2MQ
prmTzDhZt95Ui61N/Ryw+Iz7P1VgWVIJepTnyAJ/EDwdHYGyitLottdcg2RLSRxHc+p1vQ/lIlVk
bc4D6rQ6EX5pj70XHhgl1tXXGrxEarkGcqclma6FUZsQmFRjQRDrGDW5Ubiwf21XSu6dJC+v7LGO
6jXkeyFrF9WwABCbf66Fe6iqMkecVq6wRKTVkvV8wKTf4auBIfFucTi+kVR1KrrEo03TjdMvNpoZ
T4s45krOMG0xj6Bex82M20a4QP4kuxb+VO3IcR8/q1vzMNMiUIN+0Nixv4lBYq3g7I4NX6RqNfWF
adjTg8XeIHXiY5t+6iyqb3QN6u+kxiDRwB9BCct9WcOO3ksHozrmz0hj8zu8l73X+4HDpAX88Jvj
jFVhP/oJDbNXyKOv54vMOp7n3+UBtHZ5kO1TzntOsrLkKHXnMRvwYbjNyL9fprKEDvUPjXSqTRgs
l35fHtN4GIZrsoGkWs9uaABxt/rP3POvTNyGRyuXpCnvCa14PUUGy6GtppPyrnFOeddyQxQfHkrF
XPNiqdpvNhgszrv9EpAmcdDds73HEOH4JP6cBinFFDO18zoXdpA7JogIMCNQIhCsjdkZ8NMAwgiW
jonPvo/uUNbPWyfdMpGPo9FJAHNB+jngxhPdxrR5v9errw0qDcc2C4FjZfuxRyYDqMnOCpJY6kzt
eh8yYo+Brs+8sL+Nrny/R/fCxpq0RyeljVfIJbC7tf77oph2i9akpHiKKbu6Y4G2xW9M9r1ivRKG
09XGgzCStLCLBrgOJNvOIH0WPHC+YR+JfaaCXPcRw71kpRENI97D8kiGS9keGSjUl5qeCjHhH89U
sHRw27zUz+QLtoDEJf+0hatfn5Gzo6dJl7fLD2Vu6ACQrPTkS9ER8YLDydGNffc9jUCi8ykh3jHl
99V/NmQ0P8HqXxX7y44vroPZnZhcBjo7kdYFMai25IrT8TpEG6ZrxoZh06KFOusLtJ9L13qGAYNC
A5Gw5YtI82ESRlhifljvIy4GCKnCs2YP3UzVQQCLIIkwetMVXxvrIikU468W6czR1Sujt+C9PYYT
qqUTWRd6z77sc7zoLT6t/BojcCky8sG6Zuyq2q2t0uuWrLfVAfPR4xNWJZbDYWGPKOWfawkf2Wrk
1NKpdvY3GnLB7F7FYEQnJxl+tWlPUSSe4uta/ezy70KxVunqhzNyCORfbNZnvhqSHLu914iAGMgU
OPJFrhm6Fo67IRfQjK8+ji/YsIyN7t2DgzbMqJAAEUY+Ky33XXwNaTgFxHe4ZSjWhf6hWbG14GT4
pAnMn9kGgzNrq11CYsRqso5+0UMS6qEbqCFuSo2wnnf+gIjLHcJyR4tdMqHt0AOiJioQK9ELeh7l
gJV0ZLqDWEV4F3OlVZyyeKWtTpAHwHyyV1hvWvSXTrUTCrpSC0EufinKgRVn/P8PaKhnue8qKinJ
Apj5BSjuxwaJQJBjRBvBfebOiRLHEppqC+SoUua0SLxdSkpUvMt7a0yb52e05epX91EY4RlvrBCa
2azlkTFz1O4CUSSzItiGM/bK7dI9/jFltgQ8U+A9fAD8l3hwbaFC399yvjVADZQBMzrxNKBd8gtg
E/8phhRyA0jc1g2q04oZZBp8BnXVGE6DTxvaURY6nYXwqZWaYh8/tVseip7I9tV5XModGpiQ1u8S
swgW9prtRTKcOYBkV95Wi3qHNuQ/CCw5axFsQ2hRQYbhXOvsJLRkLwWOZULShaI2cYgSjzJ8r3fi
HsFK3OvCj97kMy9Cr4222i9eysLspO+/rO9vYtCTZzV8uIoPL2BkPRb6YV0EG+b9vubs8capqTuP
h5efP1XLrVVRMoHXAyU1dtpz8QtbbTXqHNJmU7R8GJXgd4YoTD7M8qXkcLPFaMsCSLxA2YUs2gFk
6JL4i9S6V3QSml38lsefyfhPmgGKUkHBOYZr68Tzk35ZPoRokelCODbTScDdkdV1ugd+kRdFyU1c
tY2JldXpzq6JFmx1wW1YOW/QNFxf4pBeHOhrfQRE/WcV6H/dY6ioDxNs3zMG121k6tmpYbzO6lL5
G5l7MLdR8MGM992ybjqDX+K2COk9woq5zwY/0yCE6+aG3QIslKzSM8Rm92z9C0+8PBdbXr/3U4N+
qU+VzM5+ArosRAAXzYR0wIhTCWx1Smjk63yrNvOhlRRG/7RcG8/ti2dds9KdeRik/iLN/A74JM05
zsyAQUiDAPlV1LVJTEnRhBPdRlyRMHaBkAFyCLNSx6eNM3WesaNlymlVQQYZcnqeZjN7ZveER/vK
euLHjBmBNp2oEgE6prBsCW/zmHNhB97OzEGVkseu4Bs3qc8MfWQXz8supaiDJ3wq+uUHsGkr3dkn
ysyUs1Vf4g6GS5xbYe78NAWxC0uzwHrMACyXyijRvpANmk1zbyK9CU736CyZlkGxZ2hsaF+GbY85
FRj9m31uow0oLbXyHpmEKLPraEukEfAAt7wKW7X2+82Sx5v6xLpLTUqSrZh9WTBaZqUveglRWnOE
At7uMHLtjdfQLpACQN1DixKUhFsCr7HMkn8kMLA5FVS6oUgzMMLvxrc15agLQHx7pIU0pKlWPmso
HDzdNtnd/lXNYI+7ZKcJEzThOTsBrDMz1mKVTN3nDSfx8Z9B8UEgLwLV79sE7phbjTfYZTR787R/
ufCAaPqw6EO6pd8nLXb4bGBRVHijhBWubeRT/0x+y1WIkWkIS2NkxbTg+9PhIfzibq7qXbFEwKdb
LIi/ebvxr/q1xj2t1cZ1Qan7PIFSaW17Ds3O2UDmP+as1uONTLEMKoqLzgTd5pR52gmbGa4/JRoO
EXCY0R0VhHAGF3zIx7Sn1/QI13yQ4kldkzt7W83/p3ZRkjgOCt/jjM0suZUVs/BzIgEc0pMxLG9t
YRB3HCfjzNmyFfY7/aWrPWdSrK4AEeSs2Xki9YtlIVlMy1OtNDtXjil9NYUnth4a4Hh+h3YxPzRh
h7Nyf7uWk9roJM9i1mzHJom+IM/TRVh6oeIaORDHD4dzSYWf/GYwE5ef9kBmgse3v9SsTzB/eQJy
FBeUunjILq3HovigwFhboF4+FlxbJjZNAOqDCrFpw6x9nVn3Yz1eOuHc7mwkoNgVd9T1I/1c/XFu
uvL6i4nUBffGlNBQqFVa5KMDVWhjxid3MeQbxhSiqRjybI0LOb4sAvlPnrPV4L8CTfio/Rdyb6Sq
NwpWS/UaTyWbpek0DIcoOubWnetmx5b74tOiwb6yJ5/n8GgQVFqAIHYSm6XJib39Kk9gsgGv0QK3
o4dy6sklU4oshIItNH8evEOUbBQ+zBy/vH19WdRHoFuML9rA6ZgL2gyfdr6gDygf6Cb6rl2Y8LAs
h6931V18cXMqe6wPu6HAtyt02WQgH0ON8jmHh/7uHqsU4BN90rwRuyrjkkI+scuZ11wMHgvlctzp
lLH7LvTKg8G4AXNs2bP1qHGWjl/jDzP2jhkMVF9X+KZIgK1IPCyTHHEmJYmcFXiiksFOz1PX4Uyf
lpBosQHvztqTNKHT5rjm4kyRuWUF6m1rDnCynpQj17kkzyBZqMhRcKzWCk4h6qbisAnSYum4q54f
M7CHBgBrgD8AFFYlmVKRxPv9dpvoT8gHhfcByYHBxAfjCP5tpF4Qg0ZfAdz+99s8jYnS+55DRHl3
ePqUZK50obaTEGJrrfobBjFEopP7q9twJTssq/F/PSqLAGPICbx/h4N7LN3vCW3yWCsExaI4nSwD
NeM8zhpK65I4aUxgJ6ULHdbqL4pbmypCp+AfqSE7VuMgADmao5pkHOZRqNH/UvuuqpPHoi3WySzC
rFWlBdJ31+dXifzkQ86BYstaepzcjaMH0Pdrij1e99E8b/sR6WIZM9RoxUMSJZBO3oDZ5tb6BgyN
Pd4yVkl17qvrdHrWaX4PrTpPCyJwk4y0NOKvbMo8hjJg1SjJrEBZcyWkA6ph7iILbmyQS+27d7uc
EODrczsH4JUXXy3TwGHBy9kxDGivSFalXbe+MDcklZih22DyJ36TTtNzmQmnjT1RHaYGd3Lodxqt
Tf6eNIswzYgO8XM4yRjAZFGfMjK7Z2LZgCnMasV+7aENgXfXLeH0PYycx6MEHDpW8OcMqjYqtlem
4Qb9HxLBqJ0+jvaIXDOxZ6CRrOQ1cySDAi+su9vbeoC/UHIh/fw499qalv+ryeJ00jJss6ZNhMqS
Pj2gt0pjmXf09aM9sI1uyxWAVdG0D+SRejEPsx2Y52uExzRgpwTfxl1+NMO4nVSW8i2OSZUX7GQ3
PKPzKfk1uA0wmHtrBJCe+LE6XEa/itZK76OIpECWoNooG6Ofsh7Ed6v6qOMwb6yjXKRuz2NgLTfG
tuPe770tbVr5LApAkTYHrXc5iAxvrSfX7IjdDJWIbnqhMqr4aI6+ZWYxFV3N+6s5BeglW0cmZZvM
lPLGupkATyDLQ/bJw3218bJpPpS+x0MC5A7EiNaLcaFu2Y+AHfiDnz6p9MJvFizMYzWPf4hoCDxh
+IQsV4L4yhqcLhnytEU/+NOsA0lZ2tZzqHpLExuion6QO9M5CVD9hiP6+zwZ/mCSKC9Bk0A7pfnb
pJa5SQ+DHg9Yl+agrYTYDsbutlNxjgxifv8wzNF49SGB9lV4GEAkSX7jNrSN9rxI2t9C9mXtrgZL
LsC+QbI4coSdV4Kit1JJuSoNuI3QVs1nLdPgVH3a1/xvNsfsuTHyqo+nRDYjR5D2XR18ez82CYaQ
VmTyHiiaJxdV+lnKV9zLd/pa8Zu9Oy/9l4n84k/HwVPVznQw7IbE3JpMaDeLTQpMvAtX3ZGH8UWo
hVPSmSQzT7Weji2zMZxhyJeP/tPBrt4WnnTkoE2aRVzWKItYf17Axl8RpHFZY91nOV/PML35CRmQ
/97Hv3RmNsJR5d9AGVC6TLzPaP4GCDOFbEVFJ26c4MREn0CgPKDUc6rls5hGPrY39eEXVnn6F3wm
X5ZNRZAsA4U+WxUSVQdH7qWGU1Qvfm9SGNdYIIQ5Xqp9ugj80XHkXm16gWbpstM5MkWT5ufFRhJT
YEkUObQxm8EXucv/s65KVvrG/Jo6nkLT2HWOpUzZI6hax18/waGQnAP0fjjmK+cy0iedxyatcvF+
BGlMbZ1Tz2YNWYKZDbqLP80eZGeNPwKo2ycnL9JJSCpmhlx5nW4ID6IMmRzzrmOwCbYg0PyvTMGn
qrOpE+KnDYA01G6VxsTnnJ+A7zaoIOb5vTwwi9LbuljOi2K1RbOWNcP8Q40hZXkh0QEgtF/wBlYO
/AJZkZ/Rw6N4LWNYRusvQ7gfCRtPGuUnaiWUOid9sc0axD4917NVMBMkC3C0Y6njSsB7++ahBw3D
0qeTH1AzJJnzinvvu9h3RI0Yry+HNlXR+gkHPcsPvGFUAMRsunnFp9No5nmtGGh6jHCBHzOD8DmQ
z5mGtR8ZuCESW0KO4LQyh9Wy5UC/11JFpl3T3da2DS+DUNyE7cwvcPGSim3Rz4AialpS2jUmTmBF
snUQM745kuNQ2uzUIbcjxvq2ih9kvNH1Q1CDAxc4OQGMBajMgudDyH9cKypz2S053ErG8Kq8D11z
t1e0ufNVcHVoALdhcuz64txW/fpB08aLtYrYwYG+QEOraul9yCjQXCRBVRWPW2BdAWQoRERQ4gn+
EPCmR028Wj6gKKrvMnLGId+Z1Tgvw91NIvRo+5fgpEmi6hw47m8kNBgYeoxteCb4EtBCWBB37OIU
15uQpa2NA2V/4OSAHFwU2N1zYlN9TG3lDYk10K4FFmbHhrpfVfnX5GdxXhcoFsifIptD+CA2CnML
7FtC8R3Va2rIaWl72wHL58EVOBiE3d0C+iGshjIndliwmQ/y3BjMAca8rckxnKoqZpwu/1mhiBcq
Dui8vTBEo2UnQ9URWigv6ssmGnd2QnY9IXsWjkvMXPAfGQNBPBMPpxZMwdEUc/aemwcx8m70RqIZ
zzvQewTYbC2W0hAKKVPCk5JNG1+Bx42uaA60NOVHHG2d892SDfkV0KOuCzWjcSfV9g8t56Od6t9s
tN0ncOlqgKJzHYVE04NTnqWvPzgiRF3WLKuMmh7cps5+/KZJqxY3L+kPJg+Q4GGMZ1EIlj8FWX1r
IxTkrfXUYDM/cD6eDq0kdB2cmAiU77Z5JqHSlVpaSTF07BG9oH3t/Hdu1Md4ELwvIDMSHXMR4A+n
H0bRt16PDz5kVHjXX4IqioxxOuxaR0WoDy6l7lq6zs5FqiavQkSw+okISGGTkU/qG8Mj3I9J1/f4
dTP2Zy/qra3D7R/wd5jqvNxL/FyUfgPRdoKCjkLRJwVXnBK6PPMJ6CtJ76LnyijKg9FUFHF+dynz
gNLqiXfoITPrPJxS5pGsUb25NrD9LILB/8THB0XxI2bcLFJQllQft6R0hNRszcChhHDluyu8jqUh
630R5Z0nilO/6PyWXRR712HbS50gGsn2oS/lmvWLD/ue3DMvAWlW14AR27heCKwMQYRnRw4yLpQQ
4RB3iKXRWwrrXy2lMVn4CmMg0NvhzmUpB+fAQEYDykq+eVAXixzCrpDTeJluQE9qs5HuIJCEumWq
360wkYSKfFexo7RA9fAOpLf9MLdI01bwv4YSJOwPX9a8hBP7CzhpnyRDbfTt4siQM1WLvVLDm01E
m/Mgxc97qjsN4H73d14R3IPyrtTBulErLKxkI2HitbUEFprF/Ax9oSqd3jrp8wpqPSWF2iw2z3xv
SFch1QtQd62rOfXpd64TGFvVEKyScbSV5QNE6o/5Q+bm3peOO/bRR8sOg25wKq8nIuEywTTubE1F
VifTXnCthEvu+sUYp7RUsO4GooOqm6997icfwCeVky8TjzMHmpczo7Gxn2IB7+jrm+Mg8qGsflyg
FW53IqH4DoEr/OVhAK75ZEdK0KCIPSowYEkXNvuKGnPlZPnT3CvbpdRMBCYy+YeJXfi5G1rS1f4t
X7GoP7o+zSDqKwX8IZEdu3yx/VTSbdZCUceNGDkkLhfJCK3ZPBcgj89Dx/4qo5K0RD8NYcRULp2W
BiCNDlhfLZRuplmKMgusIdCAsg5erPrHNvChkXGUzUmRlNLrj1aWrU26bQtUDX26JKW1DBJHBVO8
NA432b99nHY+UMxR1chtd6nNekZbZF92coZH17SI2el4wuh7QgcJcGMoBrp98l1Q2LOkptfaDnwy
zZx5kXPGukX41XwwK/7Ck7U/j6nMbk0ZnvZMlFAvSrn2M5Or3e7Wv3v47pbiQQTLb1vpNlw/hXsf
th7AOGQidqcPbr2++xevRwGUxkZRN1rnBLwUBtioKc0fDtxrDZstTEGNx31CXS/CLLPQP/EeaPgu
HfFHiWEgZ0pntoFgJLpl7IlswLm8yg9Wy8D3suc8pLMABSPSxXYBAwPHi/uhhqPdVSY0Z5YiCJ6B
/lUeCNPnLRcRLJcAXu5xXFVDvBJ5OlJDNNqKxd2OK6MNZAdW9sOPrTasFqIuPB2MXtwTaMzCq6Gq
RLyZh7+Efgzbi0H9llXOSYDGzN2x/zDzeCsu5HELxGTygd64f/wjE55ndWGe8by4ntbo4ikPjk9U
uUZXtDSKu9LvQkWXVEkvPbdoRtK9FBqzaHKLLMNTzG48lQyqDl5gIVZ6ZcqyLUgWyk/pzgAX8jj5
wSqFQVVu912ksUAJ65ePUMfcRX/kcycCKySJbdGvPs+gS5PAOwAHb7d32mnFa0qbyF5lrQDo8Sp5
7VT/+ZX1Z8RoRAn1HvNTuKaKUKOY0oSRuxQWqE/+porQd9jObDtBe4F9gF/6yeQegF5Wb0ZKJlbV
7S7bBPd/vehxNYDd4nIKl/zNSleJf3O1KzS8QJT9xjBho1zrI7vKK2hPz5qJkXrOUnP5/0Y0oldu
iKfO5O4LDS6PwzfygSmI6T2oop96a2NBy2dlZtUBImQX4cPeb5zwYQf2ROlUT/UKOnJ6kruFPZ3j
kDA/FEIdyKJWCnv1eEwTQf5oXEsoy1+HyC5VXiuvX9UMGpKudAb4YaA2E1J59KBfQOHEmfD4LGtY
iRoWWbleqsWCKscmBvfPvYP/pqE/F4Sjg7EOy1tK/81QU2N8KdmHDx1nrPzpsol1DhUhbWSUGiOD
J8p7Agr127t9teS3Sefu0G1L8AX4i92kUXjl7TJOXtKwdLPT0ytJqcxMdIOJy/YGje6QfyQbtxHw
0nz9bRdZ5E5vNqGB07Nfiu5H3nHnmp0lAJEmdZw5WfADGc8yZ1pDcJUrdtLuNlCd+9ACa787UZkQ
rdUgZ5JYPzYmyVhqERss0Oq3LwdlhlXXUEPECJlonbVotuArXPCqWXuJUAErZWNUrL4apd4jT4Oq
zJ6E8hxgm9IPe5Ptf31T0QO7jXXrA8R9epmLQP17sp45t6OoP/kl8npDXuNzWBkKQ1J6v4524Q2N
1hxvicK2CSquqlCiSWyhl2DUuuR3OmKOyJvyiv9sBVDipqbaX4V+jXs3yX0G6qpu955cexRSO5Cq
lNBbMXDnpriLRtXk2CHQIhIt5L5OdHah29GkhQnoU8xpw+cLHwNpif/IhbWauf9+Fuo0/N14HBsA
Trvx1s1cLHDhWEiHngYVuX1w+ibn9R5lWrMqQ0Gzgq7agJ+NWfZm0mK/9moEmqINGQKDO3X14xKV
L2Ns9LuMtIRWw74LtbxZJlInozszgOTpgzdBKIHG8yNZhW/MpGyEfJbk++St4JqTQUfU0ApLfBcE
enSlsAC+idyuJ1A2sDdXmg2rm3tscAh9g3N4dPoFzjo/JnVnO/f6bz3jCPJbtKn0ptKsDHOnkSQJ
xuRwZR98E8lZGiEqmjGsreZwp/aHtwFyOrcmwy8kSKVLGUpTcH/4mGWimzv8/z7g8gH6CJx+iEpL
efW4Z9UlZ/BzJoILziwYtqbw3gCMK5YxoZb+99Y7ld74XQT3EiDp/Xthfb20HN6Xcj15/hM+P2t+
wUcLcMXCyKgOON/sg9pndPte26hGErL5h9LaqkMvq306+sxd0R3QBW0JK7eXtlc6mVOYA99XMe1+
CmZfEq2HV15hIlEQU99oaHe5mKi6pI4Jjd1JteTC+/+aGJ5m2WPgzEoKLT8l4GyziX1nHe/BeAqe
++LgSWxPxOHMiXdf+a0D0gLMTmarU9HNIXf4aYLjEzk0ucL7TG1IEo3Z3R2+8gC7LvQ62YbuQQws
1R2e5w8Poa1O3zlPpIP70U8gagnM7Th2UXK36Uj6G0qh/QFTTyDOOSmE/2ofyOc8mNnttNUademw
0zrqoG3o/yhbsOxZEykrKXSzagheQ54MTovOUCC8DHNFwmaypiHJtr5Pm1hohihbHGgUSMc+tskG
F4GULf9J87pTx1Ck5FfDV9YHuN0RpHtYxyflmwzOpTgDHx8/P7QYjtd9kcnRn6njNVGSmADP4llS
fbDHhFG5Xq6QgoMLlS8sihqQQ6Shp+IR05/OKzuu7ha063GYFfR3QvjXDOiSwPzwS/Nfvcvo7upE
YKE/B003RCCGDFh+G495O1rs0anOxMVugBjf9s/zwEo819rWoYm8BQMagOz4b9wmzHfx68X03NB+
revow/m58AE7cApVSts1uvoPVcAwnUU0N+JE22zVyC5xN2C2LKwW5L5fSz+aoSUXvP8X1077f0xS
O9yR6i1Ic7OqNIfgaLiCxavYW1R+bHFdPyIFel2csIaRqT3hJZ4kIhWRQpOSQeQ6TNmDHdz/4Jf6
9Zdfug7WWyTEavwoHkkksDtKyfVpe6DWWjvbduij2wc1AVnOg7yfj2OjQz4cvhWXbV7YNy5e5VEm
XmpLlnE3ceXFJbyq+/PrLAuLF0QC0R4Ih8+goni0xNZUG2tLLG8nfh+7K88R/ICoSiOzxOPkbkY3
v5vTnpnxM2r0NYclgCGW+iYw1G/EnkFFkSQx81aKO/qi5Y73Bo1atTV1l4fQ682rCVGn/d3WazgI
ROcsxgAEl3wEYD9iqz6OjHsxV0f5Q1sBJE5WodUyF0lMODxY0/4qZyNG93nvI5pufTZYrKddJx24
gdk1KZ59+KunNf0UgRnCIPyUTb2sPa7YtPOTW5jvMibNLJ5sCl9JAIii05Ys+bmtRw27mrRPHj5Z
/5qgliBFgoQk8F5nVzxxBtyf5V2Gb/19C1VlJn8liJYKc2qpGXSWqdgzkiDz0/iagR/RGzldLUBk
6N92zPqggtytz5kX1CAoZAPRx4/QkWuVzfp2GBCbdp3CBrWnv/dGWmr65vXmTmQYc0r9vNem4Xo0
hf0HI1909VjOsi8lIdHthZCmdE056vTLf95ge/UIr8vr+yAnb9jlv83WqPL5w47i8abyeMd1fiht
QI2r6pncinW3Sl/ibwKHKrQ0wBU7+uDLVVaIfdgHtH1q+9Lj6rUvt54Z4ciu64TUuYzR1tKuxKOV
4wvNKaBIFa7Q5SQGa8VP58t/Z7xWjN6909Dwl+/6REr7AZlljomTWsSDdbaN4K2GB4V5s/oBmWQ0
/DIg8DT8uByDhB8EkAIcRc89vOD2ecfOevj8vZNd27z/Dx91acNwWora7hr7XSYxmYdC9Cw7V9XQ
Ksutqz4XJqD7BlRJe7VrZcmvGdQ/5o47p9ewiAlF02EtD5XgDbEJZ3cO+SQcaUGiBKcnCXSKdw2I
pq3AjWbzC2latVspGuvMNvzG9QWoNXwRfzkl+KIVsFEPqj4sU3Hb1ACHWOjhemkckYZHu470U+Lu
Gg/WvKNGg/FgKkMWPS83EC42Wy2ufgxdQmSjQZDv3mTL19zkUWZEwm+H9NH95Sh3UwbB3rk+4euM
SWfaO5sJ8lfTcDZD7jooIlABm7xkKR8q+yOOrph6TdOtoTFa6vk7uAFvL2sfPSighG2gh7QGPRT6
cXS5UUJtZIjqzcOSYgRWzzM6q57XI1z80gIO9onVAdm/RmHUCkCkTe9zYQ6keYZ85PktDSRRsTKK
tx5+b3ZMPBvjM8XQEZJFKuysRUKGnqE/r+LrdNDj8VsO5OXw+lM1KgG9eBqPKTNs1LfMWSJR/H72
2GCTfb6IlxUqut5w3ugUZ1lJoGTqL8Dq2CyF0g7HiqrzecbD3LlkEq3UdakbvZjVVlg3yEukGo+u
ZO8plUoo5/erHe1WBMIU4GNbRBOebt4oSc1R0gwJPJoxvCBFK9mRABUdffHK8LKoQFXNW2cZ1YjI
TiYvbeCk+vzPLZ5XyBvhRpCf7zr3o6zMUhiOXctxKSipne204a9w9qlKECGW8Lvk8mwP3BseF6Vx
Ph7zMsQMSpaxxCz6WYroBUBYcXjoMMr3oN0EIhpLDVggTc2trl+rDXaK/fU+TA0AXhRsdxBrT+Ex
uVyfpB3knmvV8UUd6L0PrUwEPhkE5g4ECY2PkZT7ig9wfiSews9BKD7crqM8CjICy89sHWefO0uq
BhbRhSOfnxZsGLR00b1cllsU07oqjAyFB2E4obnd5mjJKA+iTIxlFnz9vzIToGVjVcWyXV8DFom0
pIPMiETRGx9ZxPXZP5oo/kO1gfGqG+A/1cuuq3jMe/SWjHNf3E07/m7wBs6FMnGkETEy9hMgEyuy
b/41MDTsEzVdN6PtkDHYzOUukO6kTeUUcJGJ/0qLZoMQlxzCsgazWPMqVxb4fkxd5uWZ7gkNVc5J
g93v//Y0KUqmY45m1eh0e3nvkCEEXRv2OU7T8ldPq6QzDoLyaHy/GrMai/Q0b0IrD1VJXyfez3Ie
7GrQ8ITADX+zXO+QWATEQrKfkDcKaK2L33vDjvE0j0rhgmKPVEZQJU6LsHZko4uRwdqr2zBzGMGu
sntFUvJf6FogWDgeDNzws9FKmeOurc/WgJebTGEvqvj727fFxcq/jyBW4nVq+V7RpGN2G3A/S1jN
BH9GCeJwmV20SfEtfF1tVUEBqidXKjwMmYjNPfCipOpbt4nU0dNTqCQ1m7VTp2AYZoEnP/Gaitzs
M5VW7hyLEIaEGxcqS4NVro4bogJxhuRko23BlVTkCOcGm5s/JwfkqmRuQe3mbP9cfuGOBkDSTncN
e4VoKaLSwKyNp8QOq18VeOYgJxzns/0AcPOs3X2+Bf7EwowXwYzsrud5XQiprvG1gfb5naESGmwI
TBExbD3kG6cmWGuGCVrSfFDMiWxNbINDyro6v4DfXL89Gz1urZO1WX3f+P85+DMuT+DOD8uj5rpQ
2dpmxHoU2mWqLLwCI15KBBaOfPMmXQz/cXP3wEAsVMmwsKgKCA/13CGYqWgEuKvmyE3RFUY1cTIe
Kzy6fdAlZQYTvRDSuKCdfJj/EMsakZ9Kmk2sOQMbmzhq/27asZvnJYc8c0hlsT47czn1uazx2gGv
VUU64ss/ZrsiG8WTjggFNvNINNXXgaxH8ZfNG6wFnHjMzM9Jp9YzA0wdrX4Lx7vI+wyJu4p8QGyX
503bF7QVwCRxyqVCFfm7KcFsK0+Tfh1AwcLKKK9S6DIKAcx7Co+tqgb7Y4SUvcneKT03CKGmsjMc
ye9DMc46OIKWZ/woje6zPYPuRNYE0nUVxSMhO6qaDB77ZL7UHTzP/AcC9eeIw9ciSt4PFeQism/b
pf8QKgdxYBpsPvp/08QZ9QAh/fcYUnezTfk/8/0lMQ756G061LNJjH1aOQNcVISSpaB1eTzdldlz
2bamuSUeNPBfMEMUkLvZssi4fRewHjpuomn6rP3j7ISQsXl47/uq86kSJxRaZCLWsKNWJ1QlPaYh
N6Pxq3tHrDSvu0It49z8AEt889yzzMBl08lrOwpQ7s/PFxhMCzaqsVbFl8EvFpaY6Ffga8VGeKTD
RpK5Sd9T0MGVoCSl4dE1frFvZ1brLA6jiorzLhUX9V+usEuAmTED/Yhj/4zkmugEBDh8x5mXH6nI
C0pGvtwSjtfRfvK+Qt/MGdgdZIqCP/k84ItXG26Lc21F46uMSpHFWUs9+k46LIgCEJceCw1cQBKw
iTZcLPInXQBDehcbTEj/EXfG+3/FOBwqC6DPUbUSJVdbuB9w6mneuzKR47ZpuX7nHH2xxIjJr1Nb
6rNq8+vmoAkZnqvotX59K2gcPtCrIEuFjbnkWkF4PvwTlRkbPtUbN+PqX4qQrfWg1Ir7GSilZyr+
vNI5Uv/vVfl0MCRG+j6UZ1QPebZ5iCVJptrlEneS33yq4bS9VgT6sVa22rfyaAY7zsc1/hhJoYhM
IFui9XXfO1TrXpgVJTrYkcHR/3WGFOwalp+Gxv7qYGl5Mfg5NXQ+jErdNmVZj//3Ksllrl4EzTkk
5ARk/3luvctQjKdhlIVdFCTkBIjCQRubTGjhZCb3PxnzeanEBQzrIf63oEK68tb9p9AxLfyU2pGB
6brsfQf0I5i0STHa3e5CeNilakT80UL1VTCxPZypaR9KmRO4FQ7PrbYyoIpns5r6epSyA8gLjBuk
cctjS/kA/P8R5FBGsZTBLLkMZ7nU37TNe1ywgWh3ge74LjX1hsCRgxf0FmsISD1xEehC+YxxfT7C
ZKUITDaIVBls5rD1qBpQSc6+vI4vVnbsdG1RCTtg59iEdHc1L+9pd1wJn+3BYim5AgzcMR2w45aV
v+dVbGp6RiD1f0Tthw7N2d3yny9wO6mZBwhqt6Vi4nv6On8WNfaU9vd0hZaSGueF1zyGE/5oXE3L
IUhhyExhUrOulyOk7GQZQlPm+xbpDcCohiK5vHJEU39ibS9qK1HNlYG53vml0BDDsuUoP6psQqgH
gQhVzfL3t6QXfUa3xhKZ1b1Up7rb4x5UWOmsFQu4UdU14krkfhwvvCnVMh5seWuXXBllm08g3nn8
vJ/ITK+fy5sBeNpI+PuEcD0Fhw2BrZUzEh8/y8e1Xx62sLMF8hPfX17mnogzDSUgh3vUufJxg+D4
GxTmimvVvHDPaoFcZhOmEd2amFk8cbUf7ZFe18tb2IjxArxdGYr+mzSIHdouYCj9hWDLyo3+odQi
plVYrA4u+uUoQdUmM4DchSvrS4J8IWXTQbKqGPtasWQD7xXTbETAYHPE09uliV2n2UxqVd76/TVS
T/PHrW4DxQFhnkeHhMYHgASWoKTOCvtQrN9xHA/U4U4shJ3T9Uqw70sxJT2IcEW/GuRmbMcIcwnA
1dhc0AoX9Jiem5hJegtp+8tfylwjU8ICO8CXgrvuiQLjObN5JW36wxPbhL6caxwJUQa2SLRRUR28
lrCa+0CNV1IeWqfwhbGskvJmL+qi0fL2o59dwTEw8PfHc1CLmFFqHwDkasKIZu/M49PNt/kHRXXL
/qXUA6OjtQDfdpiIG22gnxaxZVYSe/mXx2Zljb+tKxUxTzmabekOTcgdFz90TJGEIKlTeZPNN+LD
YHkkAdDvoKRnJuVqlCVWVUi+7+bYGcNwG0yeCfWt0mYUX+w+xF5uwm8IdXA1GDEAqOSvJ/6F3gL6
DnZiOicM0O6BXcXuUN866K+hn0eL0RZ1pA33CnQi6h+VLmuA7Vc7RxdTDwIoRixmHI6qnWRCrEdS
ZodSzW7nO3DSzV0xOksBXw21qgfTvoUp1lNi6Qbw1agnyKJQlcikSgEOM4jkPNNoHfyaDRFnulTi
fsm8/FcwaVvUpsnUDiIIzZDY9NtMnHulQx4R9M4vasEBLcxVchwqstPuhFDjpumwwjT8Q6zZVQcR
gfTK+Dsp84jNgUbOGgOjcjIi/YtZNORjoR55fEBhN09m65iWgpB1OYVQlGgOaOrdTDZcbgN0ThoT
UBTLoyJgaPsPqZY6vfS53c7ePKEL6uM/fr1NX6U9m0OdBKb1U7caOeePXL+pQbFftqc1aWPDmn+b
NKzduUdjuJOquf1Qx/tyFgasrNYNsHBV/zMsfqOjMRFv+X+KjiBax2y8nVHpCvVL5STat/wRpAG1
hg4qGPfEr2mBRcmmLh2k2kGkZ2/1LkO23vb4giMbCyiQub6VATgv0DrXkZTYJc1MkbudFcnPTARo
c/gfVPmfKCqKxCQyBC9C6/4VZf6aQ2ejWTZzjak2WjJfF5+WLNk0q+9NawW6Mf3e4PMxp7U0ajNA
10fujzXbXjyHSXi5PSyGDzBza8l5eU6UWj6oy2F42+q37esN6rL8DgLiOLNCnYeI+Bxp7L50K5ao
Qa9bdUTS3XICb0m7oTz/T+HICkS27Bj8F26HnpczX45gfpI2cS1LmhqAJxap/xS2BeOKMTLEv1Kx
o+34MMH8JLhF19UmHfqpmlIkYFBwyrDqcWp74V7xdrXcYnGx7XssWQqrHbp1ZqbjVhS8aI0Z7KOA
tsxsaQPZaFxb9W8fz4mheRmh/BeXeyc5tu+ibAaaUYuK4166nH/srHp4gIXclTO+p4HHScaD586G
+1uAXancLvZ1T/as7rHrr9BfOTbcXrMj+/u4rR00Kn8uyczva3e8F+T7XKEUcV0zR+n48qxNDHOC
4OAUedhenzA33NXKX+J6BrvzDpvMOuN2rxhNwr7mXjN5nxefBjlh+/hhAtLj8Tf2xl2QLSgLfvTt
cw0JtSYr7QA2yzv2Q6HisvD813ZVZre3o7wAd2V0bCsBDWzxgJ7bOOTEcEZK/n71H1W8sAc2pLQE
p7RTeI+g09jPrdtIlE4GtKcXt/Bt1m33+3UahZ39sTzZqzdGBQbWxy5ZqUdY0U35KRW1ELYK1nGZ
HXEsi1vvKC1X/v6E7UN9mjvVsUrTwLiFWLmoE5YeTYFgFS0pWBg2ZFPr11Ar0/OrsGcJr/mxKhOD
j8+U5mzA4URPoFn0jYQGDdh/C8jjH4IqDKmzg8zSxp3Thh5OFivKO097AF0rX2OA+TLeRWlyheRc
SwzLou7NaWcwSGeNvfkkcAU+UBW698VBLlc+s/bnJwEUVJWkriG5BLaBiyxCZeEu75qEwoOMgvrU
gBveaX7hOGrRPD8ARnI5cXKtoD1ygnT5UCB+UKmYkX22sOIPjHzh4yJ90K2BN21SCcsFgNleoxYP
5l/uCWg8oSpg+QDX78ZeWTkyFjMxT29QfN+0dbik/pwJlmJS4Vl4Ja3FA2hRHel6Ff760fWNSyxG
ZaJl6z0kaEE493LkmrSVan9sTELThuvVi0wwmIr9zjbckbHUMgvf8B8Rvt0bqWkq27TiXr1bgN1o
Iwc9YXuVTF32dU3O3v1pXtUh5KXlh85IDk9YMB09xrKNnUDyDxd8/QWrkmrmNZ/7Iw4UpNDXb9+X
c3YUPCmXdWL25dGi+lwgztWyL4XPYumbs/rNWPPlwWAJQNzKzc/D6jTiKdv/Za1IHD+iIVBRGmB6
RZY1LaNMsoUUw8WPxH1zhC5hpVXW0kF0uHQFoHVHD70KrqRFwnjbhBRlGft4Kp63pJ5vSSmfF+wc
F/l9P/3BpR5uOfpagKsx8QuddqKbMai3YSPHyesTTHk99zJyJZMUsUZ9jdPOHN/Dlx6t9qTFNKtZ
y1SdnK2l/6YiUBwBxVunuc0RanF6pg8kPa1vbC+IWpBJZxR+zzuRYwTN/1XmPS5NJ3vIqmW7s2i+
gGwG6092AKVnrad82ZTm9tJO13LbPZO7MpEsfXGC1uRHJO1hH9EeZRiRJlFn6ZFYBDGuFDlDxKUT
Gh6a3Hx+KAURkPXOHW1ePjLPovJxH37ZAKB6iI1eHGpKe8FwDqwJctkzHjhJbYrPoTxekZjJy/PZ
WeXonA+nNj+aJasYhKWh8TpMJR/tAftZW+4JBeOX0Qno41Tt6OAGNc+SyiyiV2Im4PU6PmkC5Elw
MuGE9WNXYFUF53ge2rCCDyUsdloOmOUUB6feArQpn7ai7Iv8gZh7vzRDyJ3oNucMv8VckjRn7P44
yv3yMRQ/x7FwDCKvoZ+8ayjsz89pd4YIrHcC9rQRDO/xu4N0jZHXYwChoPkkMN9cgpN3dfNDBjXq
Jq/75pWehjSpV8I75nE3JwUZ4ki/gVhulNKgNyb+EqLOI0A1UWl6mIdkX8uwVBBzKUSkMtBHCYhl
CzYxk1kyD8JBhDHRlBzMMpyxHqxe6xhIOrnGhR/lUKTWxeTC7Gx7AGaJAZViiNZ4I/+cP9/CFVE3
V3FN/tQXRwPnER7t3wZV02K49mGS3J5f+7Bo465gMSibUmTRCUnuzrghtZO7aOkcW0bgM/ZpwDzl
AHFVuxiFqGqj7gWkcB1NDMs5MLxz0WoioZYlYu+5pVzwUStrCLp8YRHkrl8LfBYI3iCHKHO8gaPR
2Ia7AG7Cff05wGAm/wuY+TMJsbZdmqy//qbQK2MhOXfuGSUeOUHtO7Md0YaiYaU1ZB4shUyTQ7YH
fzwjhtQ/cHhy5/k3KhThE1ncHqbPmRsUZ877OpATzV09DF2f1pVC9e68Iu8tGhO+nILQVQ+zoKCl
zkBQuzkQSF0JksnMR2EALmnrH97BKk8bmsUvp7fZJeGhNkgtux3KjXx9OqQu7XksjhHEh3O3lL+W
nx3vFvvmb9242M4cvJ3RsMGzuCAoc2knITfl6pXFar2uCjQqxEj1pfICvFn8X6S8K7LD4/4/c9mh
xRtFbx+oVDPBwlBBojn1d09M8mouO9FRm6AOW1rUqD5BzOryRh7FTqvz6lPzvghVhtPQmgifPdEp
2Ey06IxQnWVHicJpWok5Fu9o5vAWLP2GLEw8kQC7tECveiGY2Pc10/8+wAckzI52NDoRs8QBQi8L
jmzCxGdLNJTRplusI2FoJML6ht30AWIaelxkSjxlC04vd+1tmqYNNkbWLteZdnxqHxNHWihis5Nl
BaA2Pmy9+vxyJFRRJhl08WBdXiIa/zY22GNJ4TcpFfWHfv5cxhNSws+zg2XDW3loZzvV7f98u31K
+vv4W5yw/5CDvYJkglCkGfltvkzefRL1Jtu1sEBrzdo3iEE6+p8vuz69R32yC/WFt1TYVf9H5olX
EuhtwLTaNRwuKIJdkw8RySixC+J9skue/Vtf1R8HzEvmPSrvg6OFbKb1iSI1x9HiFZBZE+tgpwub
Hijtx7lqrEnjctHE1ufZACaBM0igMc5kzTGfzd9wpqB3UTTYg/2fR60eWyRJ0bJSd3xRGnny5jhI
J5KSMt+3ppcVbbR5ZCR7PX8rkbi/m/RxTdVUv878RigFFflNxjOpqQWp4y6PMq10oIGjxPgSjJlY
21A3vF7DDgYG6a6chMIsXMUxSwxz76XjG/AEuvrjU6AVoFdOGK8wVUx/xLnzjmpqdVLUjo/CTaun
RW02EVzWChN+w3Oav9Y0Me9BG1Nr7xXEGJuNfw3uhK98HOpU7eG1Za5lmourEP5olyycXkzCzks6
LzIjf26LdJKQUanG7fqP3UWpSkJ57nl+tafNVXmFTv8h+mz2bJRz8zz0l6vO6Uc4Dz8b8yqlSJdx
JPEJGl68Ls0mi9nlZNS2VfqGjtxHuauQWVsaaUjjlmoktnI6ZTfDLZlLUGpe4g7CawjjH90QBlIc
kuexULzX0EZjMw10dF+7IsxVA3u+dqqaJ6o4xpWhyo0b+35scnoC699b4dU5GwhmoBsohNxbALzF
pVyw+clg+kQnQh3DfaosqfPPkElIrJPKHZjwKoxdzF4Kdp0GMhzl91XGyEzFmAtQ/G3lEyUa8YhR
9qD9057riyCfIiOt/VZTumUD+g2IfzSonFyBupBmwWDhJKCExyJL2il7niygzsijW9ffm/kcC11v
Nx5eWDACTWojBBIVZdi+Xit5J7z+PW4FPr/2jbaUV1BIJzxdLUgBmpLkAPEWboiUQyh+P6vNZnLW
YxZg+fPPM4BsCZBVYE7zfxVSJtpycK1FVtmVFeThTzmMEN8rCuBtwM0HK+Vr3//Bcwi6ztTa28BL
cOqCuYySuvtTJc48iNwKeQHmL2SBGKHzzKeMJepNESZPErja8SJZz0Bu4o3fX7ecVm30W6THAXmw
IUMvnLr3lpSj32KKzWfiLsLUM1UF4FUHZ+w92Sr/dOhCRubl+Rueg+lxd9Pu8rLmVjc444cCaK47
HLsVnMyGj1FZFppygsuHBDyRJR95vWHPyY73Rq1DyOqScSJeN4gnH8Ke3EJJzxyn40a0/dfv+JlE
akpmP/g8vTuOkyxOrSjCeKtnJ26OPVgBX5zQ0fC7IOkqmRDmR3dSCrJsw1kjRB4UDaqc5olz0A7p
YMOO5xfQuPn4deA5ExOKIg8GOGQbMVRRFpe/rCeF5RVY0VE5zL0A5J1u1IOqK/672UevF7mt44Gh
otM+pbejpf1UwYQObwR4tASaLGHpcggOzT7ZlSafHUpw/Pep9bQKreNExnILbYndyURHGykS02c+
Ivhctc4yjxcNe1/SK4aeTXp9i5nZja+O3RER4+ClZGfCAXJf/fmcthpYhkZ8YyTaqhyhuGKzxQnl
46T2qYzjouT5gS8rthb/hYjcWmOWaCxpcBcAavDFleome8BiHwuuj7PyFn5K+b+dnUJ6InHDmlOw
u7HZyjMJrk9j11g+FQafhhuGYPVBLYCzVXJiGojOv9FHr1DaF+SWddm4hjhIrZtJE9BAcPbj/mt6
oVja+o+mgW96ft6uAbnPWnujpfgBt8N0KZ5nKJL4xLNycHzgnFQIE7kNC/fSH3PTB4JcMgzz2uTM
OOK1437+C4SaRnDm5Pj1mQ/QwJZ5YC2G1PfxKtMSlvkk5g16VxvGAqKSawHDi0d2vb9YeVrJg144
Kk0RwWQ2XoObrFEbZ7MrTYM+eIAk3N/+b9gV/BqRiuQxx3hTDFAXZM9pDw4OZlPbHAjEWFEpApQI
eElA+Y11nrL1dk0YkNkHnKs9XK3AtaUe/oWVdMFBaYRjJqz35VKJq44X5uwrROisI+Xui53rxp1c
BOyM4LZDdYk1WzYnr3Bv9//YUnXrL5ZB1EGsdBEGH09XMKFdJiGNvSd4tIDBYjTQTgsX6oOhk8Aq
CER7TYCAn2WXc84VFKykMA6c37Rud53/jVc/h9BjIudZvyh45MF03ejFozswmUFye5ClCFci8PM8
pXCnEStJLGiOUsUDjt7CImVPkA4If/uD77OkGqKVcAc8voAzWhYnzvjEAeZrZU/BN3Nn4DMxTST+
Fn2LfT6aN2F90zPUVt2BzAzUNeEiUkFGHRoVdsTjDpFvIeZxFgggmZ/CGjyM08L7SFBXrR4mvSG/
YYMfmtgCedRWcVkNBycJW2LhiCGUwuZ0bbTCoDUo/GIqD/v1Bu13OJamNPCbDPn+3H5qpm8E6kwf
JIrgEJeItEKHaqzZ0zZAXEbAjCJLL9Oep7YK/SqD9v8cUIz33WqZBrcD7lcr/e76Lo6xSi3m0CKY
fD7VGsiV1D7r0yvodGTD7sLVi3M44sxXt4D5dSfHeu8gZgPkk7WF5zQxuXEwuClY07ZoyPXKCGle
CA3gulM5NaEOFYubt1BVdrR+2WQgUazCtG4P9NG3FdGnqfdpyR2rgenl3rY6GYBteLxtpyydkvsQ
Ebj/1CH7I2ayfQ7+PRtDhmpYz+xCUu8bU74OUkFzR9uoh1JSXVCjEwmiMwryrMPOiADv+MYDvODe
fl1+3yhqMEZQNeAI0hzlePyjX7/1cZLoR3tca3zdf+5EEfVgxPnGjwyMJhOontvnBbJjeoc3Eq90
s83h7YNFV4jJ3LTiODOP50jHemPVgaLQ9YdkuiIJraWI08Lx4/84gbOgAY2hVY0PTMvxvrGRTjHb
XFU2VyiZZ2fMqlI3/9sAtlCYP7tuvmEAVNVnbUAxb192EFB0VQahGgxICL0yMSfnrHJGLCeDRhvb
+8t+0Ey3YZWRnzSj3hk2ijZq3tQvue1Mt6XWZc4UfVmhmXxwpWCknEZwfkdjkzgs4ym0qs9KxTLh
pT/zulCiK9wKH0kaa2UBGILdiLZPMolb5UMAZV/nELnb35mG9FVlaTxsn5B9PVFtQeSvuAhhyBKt
o2P21pdM6qHt6x6OQe/u3K2IoKJFkMOXJxWd9KIrCelilmNQ4IC0TStHxQGuNGwwiceGSUVS6Vqp
vs+XIzu1mGhSsVNhDaYW12xcISruhHgWW9X2k5mdG80Mh+k2TVOrN116TSVxnh352MSnjZkNBj+q
Ts/9vpXRXZznsgFVuAEH7CZHTzceDOxLwWn9bBYQwD53Fod82Y6g0/HgPURS0zVEtAQ/oafJj5Sy
tvoRTb6FsjPh8T/XgAbhDuUJbGVICruQa1bqXGm3VOoa6dCkSUDNshhcEt36JoParnNdyIxWHzfQ
pqGCAFpeujlD/UGahQ7w71BnV/donTBad8aYt9GDZZTp7EXz3Hhj+30f0p5w8NHL1b1FZKHCMO/R
wCXDzYQtr3O5MykGSZDU10W38tKJ/Sg47kE043Bl1sdoMBFAogiRbbj3G7ZhJ5F4tPdEXnRqcze5
zNsAZpG9Ee8Xax60CG/2nWgRhanF7PK8GV8Tt26uqbe5lHSVogDY1toOskN72CvrxWHW2LApwaWl
nQZwGWAOxQQa/VZGmsO6NqPkf0T7gxQrMr0Tqgx4u+4IZIygngK0vIyr2PGoIgoiMmd7ZdELEbLA
rdv/VVyQ5lwe8Bc8m0BxWN7HI863Ck0hBn9BF49+Ue2m/06HcfEOPEkoTdRuYJWdT5ZDpU665mLc
cDp2QRaWrYXWJeoNwz+jPs2HYnRHxaa5oXrd8hm3beMXS8FR2CeelH7WFkvjrtEZspRtG0Ham7BI
lcnGci/NTPYRdkmCwIRSq7dVZQBSlxaMICnj/l7rtQWUqBXZyU9/ZneWV/cpJQo/MuwNOCS1roUu
5g0LdsU9CE485QSI6D249+qJbBLb4ds9LhpVngpVis63UpXaTsXk2DtwHQcY7hOIFcqkl/DlUWNP
AgEbrSCAT8/QbGNPepRgMMiV1JpAIhBqqxk4uCMyLInYAfVUGNMO/CK4P2wfLy4nqjQhtpLwPhi4
RgPijiB4zo1sodhh1d84rivfMYTPGHTUy6UofJNUa05Hl1S7Xsw0GA+01M/pg+eVqjIL1yPHehhP
vX0AgVd4BsNixbrXJjNic1+nDQcTjum8lAtU8IQ4//ON3SeG/QmbL37vXwlNvI0PBVeTWcLes/24
BFQgP7lnYpZ+1sb0LmvZJf/2sVQJA+mgX9lVy2MEGqEvlAp+22lqeVm4PrC3gpaUHhP/IhpRl1kE
TpBua9Tpdp5twB9fyVGvGS/3FjDQw4EiwzA17XWxzSSq2dkeaT3lRyi2ztjK5VNg5KZBRy38OFHl
+l8vOn8udpkB5IM5plbMf1OxMsm5r0Hd4xPsHjYaG5X+/E1yeaVgu98LjR8IYiBb0gsLdohG2Hh3
VAoNe9FVVcbXXcpk7+FWzHxqQwMGsnnH1m8R53JsO8btWtQVhk9eENjOeYirHiG3WhewbTp/1EaQ
3d+nPgRo+t8CQeIb2bLmN8sGqR2WbZlkVcBss3UFsJd7NBCYA6DCgu9LLtLg9bmcmDHl8ncVNHul
K/smtbxMJE0uj7L5pKtq/Stu3XObQsaUeGcjP3bx3mwsGYFGhk8/8VnA8JIvKz5oX0GNEOiv3J+i
uMXzeGXMAV/CDDJQ0QflNoOrl6iWayXEkB/w3yurIKmda053SCUJnOL3SVv0v00XKY842VEdB0RI
lGrQOarsKg4oC2/JX0OIdnMW2yT9H4poc0sfjspZoVUoaLTZH5zHPhWRhxX7JRDwlBTGBw71oCPr
AeNDXg6Gy2Dn8EzjgcW9E3eS6GHDeSXcmLk6hKktfMNDOUZLbcBzJf4dP8otNa9dkIBmwOTEZw/s
wCG9PSNBDRhSrr9pU0VpQOiNFNoKi6tm/4UuokNDKXgB/Qdavo1OJqw3+BBLaNb3kr6hqJEqGzw0
ro3W3k9d0IR+50/+qanUDJVQpDnKlmBlJQss7zgmvYTP+0uy1ZnFNHBuxi1iSlGsvfgThUVmLwwe
ivY4wO6yQcfegmB7lPpyxHmpGWdTLJVOgXPErdGfNNDehfJY1ClMY5v7lML8+sB14xnxv93gSSuX
3A7pDXvSVZd5q5AxL+Kxp6i0/J+Y0IYp/c488oH9arOCbVZ2tMTVdzzy4pUn0KvuEqkO7IqPBjqY
J1P5kt1S3LR6qLjLJGN/snVNj/lsnzMJnncfpTvXj+uPUHIkwJc/bhz4Z6FPUBzwEf5gr/7cZsUa
PrehEtvx5jC//ggTP3vRYA9/1F7uP4b6llEzhXFHKnw2dnve2ap6TGM5Ee1PGMkHPaa8XyS/L19C
2OMjKS5x08t7lF1uiJbDzrcnMV1P6AvBwGpF8CjQby4xGYX5RwL4IXsz24L4+ECHj09yzVpiRP9G
G/pfOIdQKxYvQhBbSJfSlbHAtMVhdwnXP2o/NvH9JsFmrD7qCCGzN/rsaTY9xcljbeNIvmHZ8awR
TjxaqqfbNX0pIjqbENXTxJLxVCTijoHDo3oFP/Pcx83ZXctv7p8KDYVvIXCpN7FkxNWPtI3Hmk/u
ITk7KMiduvB6G/3KHtTNFgrbpyCkMVso9VZ32KRxbmpdYj5wzd7t4WuKEMsk1Ks5QALEgXoorhRl
5Q7cYo7LWCwS0Pm5HOalxzLUorxN2Sgyb8eTzzofaz2gT52hmIAtm/08WQGUNMIfY5/N7DiBkT29
lFc+V9ThWKMeP4CFNfMCcQc8rWPpwKPmJF0o91hnk4maDCld2joJGXBJSRCTkhnzqXf1dMW8+Jqk
45AASlYDn3VibZPjmJ2INKu2qcVbRe73h06JWyjE6dkW4JROB3+WcUDDAEeg9rD87WN7eA5anVqB
ZQTfPsF4rkCTLdW/iQlRKMkOqkKDxH1LoWchROdmuipWKlZCwPo0YL0MvrrLj93jvh0dkOX+cvop
bTXJSZlkgfGQ7/nurjlh2YjNOEKMaIOxZhsOYJK6UGce0nIwSU3VbtEreFwZLeUOpelPEgBBpkiQ
nohYwceLLW4xKjKl4a2+mRPdc3aDJ+w6Zta1DYrn2A+2obas47y0cvpntOr8+FnN3Npb8FhtL6cE
Lbq8NtOCyqqtiB42EiO2TMMASshxSmVfrhvR5X4WB6+GVOEM0J6k0tI9iIrB1PIJsvibbYHpXYme
RxinTlgZWiL1X3IJZhIfZGYY+fkUw/OnMlO3zspMBduL9/g/CE9eF2DSF4HF3GhTwQxxQmK2/gon
jbug1yUXkEPPwhLLgHQRdr3YVHmH3rJUzDzY2bnsl8tAlPwmxaoh/WS5/RapYk3YfA89+HaSyukO
CRkL6xfhvXphjFcC3BG6tsfBxSznXbrNa2svKogr5Cl07+Rt3hW55zIHbgNOmk5BQIV18U7Yy+O7
5W4NDfabX724BPC9FJodzsnh+cugEePwPWF8z5l23pcjF7ElBgZdXSupYmktrae5UIYkaT/GwHio
YeOTRBlY5UAXGjdTqPVp4P6uJsTev9G/GjXcvUi6SQOFU2JrZf5Ev69TbZ6TRpbM4OJmfa4WhRK3
WG62pjlwXLO4ZtydDGdq0OqTWIvk2jjmQQOuJOszIo3Jgngs++TKGV4DttXng711IcL+d9v6yWa9
95rKbZXVjnur9xHIbCv5wrxekaxDa/ELFoNzlbZwkElxtdULhYRfLf6edaYj81kh+UJx1oFnllgn
IQbfUFHGQxfSRSW46GR+usp1kAqtsYOkgvBsrCcy1EbstUzVywYG71171Uv9hbTAD6RTJrk64AU/
YBr0Pu+5R3iIjH9zm0+Yss2Mf/+TG6b/6++hJBd4MAnZxuG9R2HYZ3x0yorgKPBIQv/gBC+n8KQQ
T2gs2avkOZvcMlaOcODZ4hFMWffxagpD9JndMpPglOETJX5Cq5es+ry/Vrzy2tGfSnlJCMfW3Ggz
NsL9+bybReDfkYLopaDhYl9gZXLZUfahhqunJWfLWnFfQTivUD2Hb585U5bPZrmFffRbmgWQRsvA
OqhbZY6nHzEAtubg7UHKNe+5pEM7cbdRRYM4aY7ZIpT/JUB9sTpbrMZIAuSJhT/gg2mtT3O7PIiO
YcS2YynhQC4Df3zhP8285jcYWcG78kAazhujGdEb5waDL4jbue9LeVagBWy5t6zb9VVtoAns9MHj
hXwhNKc8griHx1W2VbqCNMTHYgYL6O9nsWxTtE6S0EXIKXa3homMhk7qXfqdmb1uesZYvnRRTfwe
phseecdvBX4FZc3OQcmiUzL7pCPmZTFaiE+49tqAVLcUsesvSc3fLa8eRfp9PUwaKcuK35CmN6la
R7bt0+sjPaUOh0lGOjiBZVrxnKamUeUGaBAeEvkLAgITXgphjxiHU6h+fKs93DlxisHnwQz+JWsk
eyJgAh/qRMb8ye2MaR1HtoO2y1OBfPsUsG+lana/JKcNB7iflIFKjjeDUHjlDm13lYGoFtnrLQTO
4JjedHS2+an0ikUy7myz6W+uMzAEzTxQ1yGxHrGK1HdshBoUAr/AuM8bQp6NsbLuV/byH4wDcAUO
kgXeTKH0vJ24JW/mjErfkfnbks0oXYHn78kyQT9yRtObitpQHClJBZoj3VfcQYaPcbXIQeM9AX8v
uLs7BIQeXvhErN4O06KYtDkzPkPpKzzcuvyzaUWFYCWJcP46YO+nrLlXm3HXnvliM/Vjs3RLFobe
RvQiaJULO/T3U3x1RgvseRSieNztUprd+GB2MV+tfz85UEA9EM0v/Qtzvjv7ob67ZGP5cp7MbSgS
CywjVzYZ4U0UPAEoO1QL/CUvFw4xGppXyDlU5ut4al7a63+VwQpv59roaC4YUGclFh9nCS16Dnbf
M8jyEG1mXmyrsSETXfJAJSiNRqaemiLlKVMnqR3uKx/doUNYGd65LWI/hhqzMkRngDu+n4YaPfqG
7kj/ulYLjHazzc2f0M2dbzLiVkvI1N0MYF0lb0Fj1hqbVRTu+WRoH9qPCW6kJvdqENCe/1tdD2P1
FGJfai29O9QMf7Urxn7CXILs2tWUpQgtQniQAyDe87ZKvTWQ4RYQ2wLKsurg3PveTfeQ9hLsdnOx
+gPxBjcO58L/n8PbM2NU3248gMNaOE0hmhvQIdxGRmJDI+KZV/stZ/W7H9Y/wHHHfpdiYQ27oc+D
jtsV0FtKEVhwGAntzeIxM+BW07rXoBUtn15Wp+RgsaOCxKcgkhhQ58GyvB4p3WXtDwc78KEwVJdW
8F12ejLNcHfBQwHXX5jtOhxcKyBcavW0AziQcY/5ma3VSirGdQN36v9oyVdcwDkkXQv+alXpiNDt
d2WGtFw0ZM30+156IgzdHZ+fhqftyaBZxZffhtwh9moBNkUeJ2DgGyjfe/uWKT1U+P4aJkkOt7wH
22ObUu60QCWe/e9Sk1TuQhPG2RzEZjfX9YUJDvNHRH2UAjmY8hwRdv0GYJGsxuFNp6R2vajHGno5
BkD8CrNEtBevdXDODXuEycRUaa+g58SKU3vutvtEGtvJWa9cTl1snsrH3QlYu3o6FeGah8hwh1zX
DqFoxeLAt08hAk2dXEqINCdO8evOJglbhUCX3wA2iqi1aClFT8PfwhF9TADWb18hkh/trjg2yd8t
e/MHVGbmJG/9dt/3uU/UhJ0DC9LIzijXM7R2uPgF8LHq45ozp0nYfuCPNsFzTjsE4aPqw9kWPba0
fxwgvNN4tph+nTgGK4ha4nvbnZ7j6TGYS2ISba+y2S3WsBsDfwGb86ZnNxGdoOSPEBQCVRL/REef
aMzRvRhy0C2INLiaAy94szqNHUO/K8CyY0aVhZWfFVVwAUT/X393+7DGih6cjH0SvKpHeQYmblBG
t0tvzmBM1ujA5d0hhAxMe7udXw4sAYh9lE3uZYQHhx3/ldV0NPmzMiHbn35ywQ2A7eR6/Dtgjd6f
hUimRGwtOEdax10SLzkSXW3tvsuM6BuWr93OL/8LTWZpiyuVUrxn4K7nmBDxTh9XZXd1z7PCfYtC
7IN+yFc9u2jlhGaV/iJkgN8/zsUluHXZ/NDqWB+qh3xHwfpeZAQI6CdlMQzzm7kyIrp40eDGDJUA
Lp5VGdHSEfOVDjhUfjGodlNl7i0qeSJvDESIDWVhovR+TqzkeSDy6mIU9YGR1va0dAyOFJc3dIb4
pVhSsuOIv4AwrrBtcGJzlV1uBcMZha3wAm5eqJAzyrvHcp7H0Dzmzbb0ew2e9aYzB4DdXnaX97Tl
RAtEsMJgJkA+x1w0X0SPTdN439UJtnjkKjNEqLepmxP8Qv+RFpiJDz44ALh13Uxp8Q1L3VwOPQhz
wG42EKydkuUldsMJOyIWqPFZNJVVqibXDT2l5m8l2dXsNHAyGpDEQSRWo1miEWOlTxoAvOBaEu78
oHqvUFCvbb6t8Oops+kIkyvWtFUS/CrhSR9I9GBaeeiZiICB0KFw7biXHwA+btWchJreQ34iHNAM
9F8Aagh/d4jbSD5qYQxQDeauSZZ4fhmMzkIphezptZPufwQw7kZAssnt2joQG5PSvEQyW+UJGgn/
B8qiit+gWtsPpfFcMnI0aiPChIZ1VTBMDLSeRaa55+8fwkN7nH3RzHdZZOXzAOgihX+ZZ+p5l6LO
ThicemnVjG9MGX1qqkbmJ4bajIRTHIH2Ihu4+2IlqKCp5v3+DSPQCo2PRb1wJ3Z1nJEldudfCT+p
ZiCc/gzDYL7FGb9IhGEAq4TxHHga242fF1IanmkO16mCA3wufgAu+/4LecFFKLETmUr/LYmYmZ4n
48DV0y5Qx/dPQU66UPROdVP1vyC160936/dCkbeUi7jniq64QFXfbfh1l0NbQngdLdF9Ebgzsaqf
s4FA+q/ttm0+s1oJwEQryiEyAIBQiZu8vXtpYB+bOjrHS8T0ANhE9Hc8lrv/4JD0pqotk6veG4ai
L0fJoFVNfhgEW+ACiW/ev07lFWbPFMKK6iF4QYOaYpP5dhBIFmyDb+6MIECooVGkb3FS6LrUUmVq
bfaW11aEpVkMlxcKuY6WonbbgyMVGKym+m44yTXNtXygWMuiJvEs4RzUnnFsDf+y3WwNuGDpXqSq
Kc4a2fHgI4kQAhP1Q6S3Y5UBqhqZgpc1WANGWftQ8+8ZTTfQWG10NKb0bAUy7qx387qKTtfanbEK
k2pAYnAgdSm8t+A3ausGjKwCtdtwrfM8dhM+XTAElA9gMSePSvSpTf54p6quInw13XuE8Sf/xECj
xkPMrMPv2aYl64DWCgdUoyyPKOsBn+ce+i3SFoa094hkCAEtosYwy/Ih7IJ6GkeyUw5Y83xhS4g9
uNsk21YFUMupn6UeooXQyLOhs9VCWcuS7QxPFgcC6RpcbqmjbPPh7TimH0Ix/Y/iRgJe6DUtRqwo
6tqGmcLPlNy8+CIxspANwxj1sMFRdkhmjvF4A8OIJYuft5ZLGhKg3YXsvDIOtTd6U5Q+yWCC4uGM
JNIwRUpYKuNnmmghGay6wlI/QHC6BSH+x7u2Ckibo9pFPW5omKTXGvIJh8wZCKxMiPKHUWVa4fPt
tPerVQP/4P1HNvH236bgPEKOclVbJJFhTe0yLm7HMHi+2hMWNI8tjh4fLqCpKfwUMQHMHXyZBTNg
cZV788Qk6V/a4Abp50TEHS6HkWSuD35AIapqBvOguut4YlSFoLUZASxg38ekyjykQHTf3d1kWJW9
uNamC/SrHMhjl83weowcSFVevkosiBRYAJ6WhOFjJbtCDNNVnyYupZg4QWBcaYvAG89EecmchoYY
Ho2cRYnpyLiksLK5gJHCnXijwQdOqQTK3xRzHK4hTFrvpQjjQLP0HPR9Znx6/QldoEll+VrDxBNu
cFzFn4QINw9B+xq4X4Ji2tVs/HKh7dVMajsZQAiEVDItPDEoLqwpJdhJ94/zkGCctlqX9k07nyqs
2rcAr2QWJm2kv9r2Z2kyCvDFsWqpeJ35Lpfb5MZex/e2UqnQq2FqEurijwrYCql3OXg7E/zDIfYD
UdD4ZgseLyKLWkPgQchk6/++ytJhjnwjA+rYJp3qPicp/POH7OHxrQ1hrDql7+OnpIt2BD9kACxr
nK/SwVFYAcCBOxpGkIwJf4e60AZHCqYZuenD5PGveaUkw66WgmY1eJRL15WQvtgAB2nxqq7pfkN/
MhgPWS0yR8Y1ocKOurkONj9W1QbckddhNDQU+GJqfghLPOBKgmKnpKt6/QMGvrzYLJc4EZC4jlzI
uMaEvwzAgq+DlY/45dRtw1JoT2atNvQTNHTYpT3/N5m5Y+o10OQPdMG6YHh1td9Ys5PlGNJOjPNK
pGUGrAvNZNn0Hk84K5ZyTDXKZvwM0i6XCzYg+rJQzKkA/spn84nnib6LJjuU4mratu0zIhAU3gjU
zXCCJ6CerJk6LuG1z/7PhDhY670F/MxnixpkyMt60B4cJALEsuVsWJD7BDts5ZYBTarBb2x2iL3N
q7XlzlXY6pGEzwnyZ2J9FnrBV+n90cSTxjBDQowHoTH3Rl+poSTSLnZ6ulPJp3U/R0t7a3eI1m2g
ZFmNGAErVUFfjs+JorTGN9jhuJQZtnV3hjdcim7NhvoDVDb9jw4CBSmhMIup5efLgdoILfBllGHJ
TmyHsf4kflErp8yJqlK+U6guQJfry5xg5f0543ug6RgjJcLm6cM/eOMug+Z6h7mFVzAVoefEwI4j
nZZeV/yqRF0O8K70WY7cYm9xCW8OPTt+1oAthRIrsheajk5fwY3XX272pTryAk5CQgOW6hgKF+dc
WOLaXFHn/MZI+T8ymC0jofRgsz9jRzqJtEnVYRcGKei0Whw5CUPHFndhYRJOCHscxBO9hRM/1p4m
qWoiDgQ4f05r7S3QsCx247Qy3DCafWD6sFCmTfyQBY1SRFzApDh851nuXpTIMoi3yeojEG2mb1By
M+hh97/z+0E+Ios4oaEVnAmxJONR2eC58IdQPDw/IbNaEyouCAohAuxe4phC1YC8h8KtXvqMOR8f
tddJ5Sp1hd7xSk5k2lt7DZyTl2Rt5CBI8piiNYVX6dwrfrcQqQwBpGE9zHjw63EZTZIqnHXihzZ4
oahgvgXXHqWXY5U3pL7vy0ZQJ1JPjLCUgKHC9YPKGThpxAbU6Z5NxmxZ14Kmdb+SaexWb6rc7fJ0
3RynGYPZhHKJHOUWVIMad72+zZbbA+3lkreviMAE+CYIEJHuQVnSamCi0moRNW7m9RNKD1gmJZcn
k6bK3O/wonu43wATe42x49pQPUKllXy04P4y3VdFlzoDNP2D6i2a8CXexCDGj8/yqmbV5h6w0UzF
I5yec1HEffnAHiEgvQ+B+XVf/utkYtwfukgOh9A0VgGUbhNK3WOBnflnB5Cw2VS3Nyg63FStbtHM
G3CHByapwHb93Cs3Na/BveDyDGCguND9Zsk1Iyzp5gBDMZRIOevtJGiP3sxZPAEc4Rr8+ah/MYiQ
+BDSlaUhpZ5/PYZ1ReGHWgZ+AmWiTxR6ANaeKwvUME9K8iyHZ7LC0GacYEBY32qKyezskjpcWS/q
dbqkOYpb84PxDzEkD7sdsUYV1hG3BzIawckEOjTmngrey+HP3ogDfayLRUdL4pSs4p4j05tLufmd
N0bZ3jEbXDQqqPnOGyj5IPYIwER4yxSC9VERP10BKXSHh5W2Lvnt9ET92jFU5vigmLHT59RoWEn1
49rlLlwhkMIFfqHGHc5V/SUL3ntAm2pUD9NmYq0lcYm9ltBgPnsfBvVoCFYSYuXRKGLm5C/clRAy
fod+uhBQi9nF4NobFoz5vvisq8rIb1jOshBgDI7DKug2vv/qGFdKNNyUDBQBIUquTQz5bRr1vQSm
vahSUWKa9Ys0CAuKuDScEuwRcPuK5FzdRg0p4RmZtlYYJcyx4gYjQy9YD8cxUGVBlow/l1nG+EZh
ay2/3VQ6bxFl+nXm4mNjvjKPWNFekl3fb3fmmSTGVkpJGNil4dj2GVvfBaVUwJQgFt2KCH3AcMqd
1PLyaOxgQCNxzWuyBDNznpgz4mhZIVYyjFdJvXmpZVWeYwDc5eTyOXAUcT/wrvtgdHbr2xiFNtcu
IjDMYAE7Tk5YzwBOoEEG11FXCQ0D7DCQJrVuLQMMmHIPxl/viQKYRhzCO2qiVYo5QmQoW90N3czh
oKg5x4/Tx/nHVU87SzCTWHUh8sMr3qHNfVIG2u0xxkTZCsn74WFeHBdwP85YwFHJ35+s5oFVMQcj
xiHhGOJ3ljzh5LRzt2MjTZKfQfqI7ZHY3jl3sxlUGDHo3nX8v4OIUyZuCtuYCgRWZ1g+joh0r3UP
S6LmcIKvWSvFMnuotcQJGxBta2A567ijaPLwxxWbYzPRisz9b1Xn0z59WUZ1mqAwJex4RNA/RJJN
YoOxZwd313uDn0k1IVUcxykYhIQfyxSRl5nPWQQ4JVIN4bPvLL+lhv7FWiukSeJTlJ8w9oofCYrc
00/p1rQh0l/7CeqSK/sAC/IuNJlFsx4+5v5M2+nGoeu3n9clMPURaL0Pt/CK5gXO77icLYr2O2e9
a2AfF33Z/aWyDBOSZuk/Iicd7xUYdS9BrpO5vGLNekSUV+jryUydI0jA1HPE9l5pP3RwbNbniS7j
PQAe1R/F0Y32U7+Vq2oz1n8innWr35uDUwmSkoB8jKBfdqho+S9z0fJDir02T95pTUt6d1Z+19Hh
WWg5UYUOy6iHMaV1aggaTqg5CrcsAJyQx0c4gamKUeq+Hj5gG1HARPkBocS0G3/ksEOwCfeadF91
G0asAs/WpYPqbN04+xkOtGjehwl7q//aTGflMPukS20pw39sokDdGzlHonP6yxSt3gS0KdIoh3eB
Pb1FozHEck//Au3v+Du9vh9UQx66724LASwkmzTLfySp+WyfOl4i3uH5w+JNjZDD7+Z7Vb7j+DmV
Sqgy1hL36clW14nX5vg3mb00s9cI3E+FUKcJJ52L1JUQ/pkAmmEE7ISvzhykYvtFCuHLlt7aa+cE
sgksYzRmqcqiLaTwfpKopD6Vz8j7b17T7z8lCJsGiZ8Vdyisztq43a7h1wPtJC92TyOvX6fuC0sC
gxn+csU2UTT5eKd+Csm1h6mVoVcCO9iIbt0DzWqyUo7ktRwUQdixOKYTllI4a9Eyp8Cgohf4708a
BX4IRTfeg8vA4vF6WQFw2HYJ7SYohd4vf2brkwhxos0ZEqawzdfcpav4vcL/hsGabAvCjfwUqoTV
axE/Doc3qnVQBSSdwQBxtMDxdADVLTQb0AeKGcCgvZOmyfqHqDBW/v+lURH4+lrzhN+sSbBRBQvt
1Yz76J1lLUp0dNMUoUr0YvW3BK31ouAxmBXN9QS5WCJ2aF658WXe39ntql8/Y5ucE86x/zgW0wsn
dbv9X1CrOGO89PpIjoUTDeE1hIAuBQpnxPcS+WF/FJkIOQP8bsPSKQUugg2Y4ur+nUYA2Zm2K6TQ
U1IaZLjIkgfltEwrtb2LpG4V/0kuU6m5t14PJBJnzFcvafxWeK2XZ0d7CDIgMFsxfeDe051eEV44
7RS8q0aob+Ocn21O2rDQjJRa7WKU4gvRyoCt4LjcWnfuFJE31V2jurTB8by4SWEEv3GGeC6OelsS
Q6AZOnw7d/MzxxZffalqK8c+vhIvA0nh7Ju08X7llFARwQyR21p1G9HqIsWApXpr748Hy4cCiJmv
K0v99m9JOf/R7iiEyV9e1UisjHqsG/LwMynDx2upftl66v4KnLZXp8k5FhALC6S5S8BhPG7XsYff
sVusGfy5MMpn3Xyb2ugHo1eCU6DdBM1OVLBet5oEpM8VnUUh1ciBwQcLgZ93gRzYn1dFkglAESZJ
foDibFbNWBgbU5Q8Vl4IuglHV6mgwQRIsWTU7pi5Tcw2jifFNB7j6gQjEmGYaLawkhwhrMyqcwUm
IQ04t3zlK0TdToM/6JNF7IGjG/IWyc8NircGhvKkJ1xlgpzpZw7Iu4oPkubaTXw/KNmZTPKqnQg3
gkvAgD0/70PS4sp2yH0ba7K4xdr23aveEcJlY6gwuRFPS1WvH/3eea9lXgguVBq9zhSthB19F1qp
lC0nsQHw8W9byWu6qTpGledabv5NrXBiZdTaNHCF73VCmPt/stUv4u3i4Cq4Ln3VC4S1vEnenRSu
yw0VB7d5O0CFwlJ7K+UcsBeNoUug6aN1salVy21XdCV9a8A/q2UvxTzXvpFhAZzsk/vBtcNWxIDt
ub/yX0r8OLgqpSKhQm2HH/uMdjM3bC5GKZkMIPvlokHFToK7TAKjHg3trMkFM8eV3Sznt9rJzt+S
nGMiyZG8eRwDIN1Tm0NgudZdH9oNOGt0/UrZJNCJ0S0z3B/GtcRy30hVWIkfDuVbGpfoZTsJip8Q
OPQMaRnycLC18psneOZir0bMFF+MLrRTeOHMEGsAI1A8LDJAxPo280u1ZwhQkNz4sbGZuVthlWV8
P1Do3w/7/Gm2UNlaOqM729gaNgU3E67LN/0AzJ1G08A0rsXDPS0kmRDNICERf7nn0p9sVUCX4QaC
ZVOWRlKhIgE3MwbJkSE+BKnSvjH9bhzVLro6SwNJvnaue7tbIGiFCI/j+tSI0vVqpb5hwRrV/UHy
20fCG+cKgz7bt97CmTjIQtpsEloo1xn6g4s2dmXLzfhzjGbMGxcj/oRbJ3cNx3JmzeMiOu8yCb6X
Lt7pA6XW379x+/VUDSiu85iCXCK0GODSYeB1HWSCBosdc6+rgyabQ6fUpEkNv0XpjYDDwhDDWVOb
mguRCZ/KRvjslvIKhEa/xzQsFfaC/QK7ct5pasquZkmgu47hUfgoFSJRqg4fEjxQh6dN3LPnVdS9
dqEUIjSJCA1DKU8wi+iK106IKl98K2vx/ZBdhtpFsGGIOLbsiEJVZdTD3XoHCAaLUo3kaMg5SF+y
DNNCjWzKaDne5u9fPygNVDBrr/32yoShnsGVWiQz4OKQm4gB5DY0vv6iQcOb/V54gea2v4BKgoy0
aEkB+uQ2MNRCGIOn1mYM1Box8x0NdlS0FDuKyx3lMmIzwJUM64k9oI0usOR+UoaUBk4zEo0Wu1UR
5nz3GJ+Y+LLHd+1XN60NxEvkUMX8HAASk+EHTUd1u7TUY+bRZ4zvaHPPj2Dvi6Mo9t2O3YNb8iBz
OMOUOx3JJLslA84v0OQwXwWhETgnQB32s9cz+SoLU69BEB5rmSa7a5RTwtAvqne0CEQ22qb04H2z
esVR/F7smlBKDlLn3X4jR3E5MQwVHBQ+Sz6O4y6ba/gT8LJ4aoWxtZ366QE4Yrjs26lij1lHIrvi
+V0IdN5g9d/PWkyhqAEbTncLWe4U1TlhzbHj15uuo/Xyv6/cluCyk/7aLwmwI7xe+gk1tWY9qwxh
J4qGvZBvdsc+sBVAqsv6oyA581g0lbW2DQu4lBDvEIX0SATo60Cpk0fg+5JQwTDJXLH0jXH2pvJu
ttqqygJSGCee9aQYH71f5IWpuIE1fV1hvxrd8LOsBtvq5AsKOw4KWuXuPe8Uw0xxrD0u/kEstTqH
QFs/guyzu4mfd+MIsxiCy6+FFntwBRWslbOMOo5ynewc74sJLxyJhGZerrsX8I0NouEYpFSKVH5R
K482oB/A6cowGL92D6hQ1xYjp1HjutR811G5K6Wh9euvwy1qdLbRayXZqboMUB1v1yvo6P8WSmWs
kT78WhTDXM6oYcnBMxxavYrQ3fQfOu1XbJYq0WdwfuWIxyua8qsSyZ7A5yAfguVEJ2ds3l8QykRj
YzLO7xi/GUuJIcM17kckVkoPwuv5Oj4jFp5Dj6ygF3vsvQdWPWlqbdulXR5PzpXKLpBl4M+wOGSz
4LVLBra8+tl5MAmi37j14XRzZgWQrphN3g0M3M4CmgneBnPmHinOR2g0cnnGpLqRVGW10QUDOHvd
0KQWl8vbjHbolbdYQ+3HKqHxovWmEQo1OEhPjRl9Z8TmDdCFOx18snXqGXSY6EQ0O0m3CsZvEE3M
WZ7RGcIyVVhm+Vs3pMrwIXc/YIOqfoApDLvCu9GtrQNDXsOVDzyRBOv5KmHbb3MDj4a+a9jUmbaM
RpEgwNsX6yHqpACkSodsby+o9RzEDsw04BbsCOrK4AXYEl+VCdlImfAwXFGsfbf8lfa/ZZiNGbF2
+fZ+HejvLXYKu4lZpeqnH9dZAVvLvi+U4XSULq7cF7jdYdc0LVV6uuV6cPHeg47eWPXNwOtBg2Wr
m8hgsD6KrNmSXFMntDax0YPIMHMyl0iInJ+GX3gt6o/KNxl6R9O1cJduE633Rl737LZjP9MxMShe
wj8Vd/zJKMKcG3g4dmUU+mVNWVMH+IFwEQd/0gmjylTGs3IvFFdn+jlRvuxn0m0HotNT9a3Z9Voh
ihbkgp9soFGTvEyxZGz68mow0rcgCz0fQI3vke9MrJBGZcNJJ549Vqs1F/Nz1EL4hEBLYFQACweA
KxP23N7lZVJ3ghA6YdaRqgNly5bIVhmIZbg38x34tWzm4r6lxsNm+rqXFW8dIsMPH/Oq/fhTYvnU
VZa4VNc6mE+tUhIuWAiQvDTo7J1GSoKF7zNsU+6X917YUP+KYMvuQHi+G306RsUBQDWCJf6YMerd
z7TFWU5b0e4CH8DDx2E8fAZzrPG7UWtkNRcBITUIEH+crkySILohFHqyHsv0FWo29HkW1r6ejWHQ
LomV5zASq/Z+l5eeSa/RYYFEHA/3EhTaTYTkDVfXGVoKx7+61hUHSw63pb44DbwaONT6Ce5EVpFi
Y58Fh9yzCv+oF/acrm+Fq9+d2xfOUYyDCSJVumfSz0dexOzOI5UACW9xCUHYw3+G6kqmjBM+pg5d
2zy1Cu/qMuJxX3KjKDzvGwMd4v3h7eLI6JHG21sBaXpGSnE0S/XhVRQursCcW/v0wcijZuCBKkjO
uq90KnyKEGGHgeQd6PUmS0AUR0kVk7/g4nJtX0VTTaPEd2/BIF06vOCNCNJSm6VXkOvomr8sW1/u
Eg9kN01BYip5DUmDVSd7M2G8iTJAdnffS7rrI3chVRD/bHqW8CTNHUIksgCzSIxhGeJAOds/CwZj
v6FXHWGYz7Kfob4L9CN5EKOCf3quDET28aC7cWmMXdomfRSk13btYPZR4F7rmUXenkb65QRXrTaJ
R3FNKmcID8VT0jT8Kfv7Lgo2EC67gUv6cq95Rtr1hHlpJnvnakn95C9iN8d7lUk8A9FmMFo0k8mC
n3KBT3Z8Gfbd0efW6M7vUwLrsXXRAxS1FcLXc8dSs+l3aKXnHBrQLTQ2vC48a0m5P387f63i4LDD
E4B31WNjih5TjLQj+xs5/fZuBgxDysx8zq0WWLxHs19MSOTb6fyyWm4oANPBuIzUO999XrdxwaVQ
NY3+Fjp4K8uZvZCLEEs1PtmmwGxl0xEsHhaAbS09kIUmsvHKfwA2yetPMSTegTmUWIJGRUAlU4+9
BEq6CH5tKAaTBQGeBIpSBGmDpf0c1Ubf5HvM40Zsv3n9i7wnWQjFRmGWKtb8ou4DfavmcxXIdYo5
q9+iOyb7tblw/A73/qGa5ONM7X9tqTOkowzlt6KLnG1PXgS4E5Z74vE8P1y2TlYl24GsSrpXsgne
TrEIDiEL8Wq1e6kj64Yk5Bdz2ArnyTNdBjA9s+36h2sfJL3Xz89liGNboxHNpjrdZmKpn3BQCuxs
j1IVCasSi3HCRzDbWzqWkWZNwkVVizogd2W+N3HHDKtsD9LoFMRqPL4b4Q2Kyr++WokZ8pG+y1lY
4ZBIF75rqDvSxiPnoaQgn87aJpg2t5bN8G792evQRSR/YsaCHBRFbHbBpVS7lMM/RiaCl1A2Hkvb
8Bz6rCevk/VfJcX9Qu042hto7LHT0fj0Qnnib4cgq+ZvGtl9rCw6FjLxAjs4NoiHEnG7Bi+m+BQs
IK6zSSk/BgC/RlQoVzyU7o+BlQw8hAgAeSifSQgiZAKClaGxAAcwlNvtMKeO9k3JJm9KwnBlyJMp
pOyl5NTydgmOCQC4kLPYaTOPxJO1RSHt9Vxg/bo+/VMU3lbM2dg4zp/BMo3LutY+Dq1Bo7U1AA+D
3fd+oUIdAKX3C7YcK1U6GjKcSnWxo4Gh/dMTwfNYJ16Pub1J7NvB+ks51+EHsOPVqODMcoCLidzp
l9/4J9EKIGn3BNTke4F32R8mK8jVhb/nP73KoaQp40B/ADqVPYUQoSA9xnbsLH8utEAta5dqXUXL
QuRSl1OC0PpofAMQjoaXpFeJaz0eIXNWcb9pffj45OxX5VhfwHE2ba0UGpCO7s684f8ugQ5yRuFY
MRhuoUwijke37AimkjajSKLKhV6wdjs510g2+d9lZVqUlnMPxawTk4NPpyLmi6AWBe6qDHLaQpgQ
4gVzlb0/c5k1W4MSlMHWucOFQS1AcOmzJiRtU84Z/zwDM3Qj2jhv8Ly3LWH3FlmxsgvDXvZMFx59
6mrMwzSDx9mNoxwSUbg+hzqZef/hrta8/EjFO8nacI/1iH8UKkR3jq1uWqcdKdwxRZgYWxGI7vH+
P5iZ+lBRk9KykVH/Sk2d2gnFUdJrV9ybDqpvd4th7/YmuoNDFbtwofCkyBrQFrEGC0+PRWcYh+kv
etwXS/fKcwxpAbpsvly7oQf82jJYjdOHAnvRLsQY5Nxa+TD6GqDDRba78unpSbAM86+YifV9g+n6
P1c9nvZddjFU2rAwkKSOMws4CS+BaY4n9ZyN81lkVLCPwjU3JTJt4cmP2WOg5VAImXD/6HUXFVxp
po40ubATGQfv5EZS9APoMdt9S3urFFhLrh/HI6he8/7U9eyCLRgwvlxLPgT80uj2w1GQAnqmXo0Q
Y05ARCqMQ21tLMULlrwctu5Z9Up1J/kg1KN9hPgyOmlEHyc3crWWHqjf6AdiX9Th08rX4REl/Yr9
FdgzJ/hTUrNXS345lDL8t2O/JcfjkmOQT1KFnVwXkcoN2P9Lm2BToT2kfgCKkNcK/u0Bpqxh7opK
lJ78wtogA4WOhdoiWSoD9203UEKuLFgMTCcczcHfax4qkyoqi1shee5l+p/hPTBttjdgAvZ1T5Nn
A5OzC6XP+QgXSAws4AH2FTXq/WqDBoM++BfPn/q3KxgSy9vYIbzaSsSy72DZoTiw+mZf+FVptMHA
IspW/PCviH/ZkTdYeSAUHSUwbncBoAj0iuTm6m+tucceRwsSjPtQw3nOwYhTXQFxRBt0gPvHGvxs
oA9FsrLTEtoc2cbkgwTJLwkUT0dFgstszoEd0877+IDqiORUI6MVU9TtaTh6C4lB0T/sd96fTijr
rYJq2zPl5GYNbBgmcM+BpAINUPaGClyk3HO5KasmfBoVh0XZK/LYYiSKaacMl2QJUBi4IAeQ7P7U
sZjVidamxZPBBpMYdgo796txpL2riPYsFqv4egRdtcOirjyQ3DfQqMluN6a/kPwq+UYBwbgJmkQs
Qg9Ilu2qUd87h30kd6o8CIZRKZ3JTA3fhEAKHeLz8PI8/LBMS2stqgpMr785VdMuASn7WlLSbrM8
to+vm/ESu4QrsPBGc6P2NuPi+6F7UW9QW2ii5qLmH4PCm5WrBi8lsQsha71Hhhq/W/m6OYpOb4nm
nIpSNS5wXja0DLcaEFQMwG2azUEsxdERSSGf3NYl/3AT/3pxufPyVbBgDMi1UHlQA6Qjmg+b+6Fv
wzgCPlMsd83X/QOcMiqUIzPvcXKN96ptYTdzKo90/iYs5va0ShuZK/HKoH+EP6FAjiQPw6IpfdjI
P9ZiuOu1mc3VgESYD/iXCfYwsvvfxaVv2+Y1uW6EPl8d85hCCahn9mwHbJQ6vgswB0Swttd0RBH0
cPIc1miBKMtvwSDuJiNFPJUFHaPXaS0Lnshd2eBZoYUuvNl9L/w8ZQyVGv13T+moxSTSjLmmh4oV
O0vjiH+7+urLtdDo/IfH6ldjI2HsjOA6MMygiZPtZONpaL1KVzggJMAa9w2YuUX5xti3kA7xj9Vw
QPLAgf027U8OqhJ2raDpFJZpRRQDtxcmmvsrtcmD/75FP0XPv+F9ZaHdJRz224hozVFaSKXeBFXq
7DrHscdxyF7Fye5A022G7aAENcgzY9xqFo00VqC5z16UM/YoH1d9aMAasEjHDbo67mJp+eiut8gC
tXsqQD1e7lu4oKIH7GEJraic047D8AuQzhxF1lgX+h5jXwPGpEQ798JDN9iipCiZgzfCJ234jx+6
2hXNZnXEmpw2UaSHVX9P5mhrCs+pQzKzqS2rEOPOO6XJC82bb6TOq9PienKbRVcW+Bm1sNYqtDYg
8nMsYtwe6Pv2U3IH0/KsrhSLa3C1cRZfSrqXFRgY3uv/O/4DlgnvXtusXLUMiVni9RZ8OdSS/774
DuD8YIGnN6nXlhZjUcRIcX78OpCISlzsXE/+9Eg3S9dcEx+itbQj+iLf6b8fPS5LUvRlEPM0L6tP
fB7bN8KEes9xUfXTJ1gR6E96zBVla46ZPoSmsMmcw793AIuKOJdWsvzjPmtHHO0pJgpWBLS7kIi3
gabXPLu0IYMyjFK23cIud4dMIQljFiZuQQQlDhTaM4VWgNiuJliP7xe/ORRpvXNsMUeCe/a2ev63
7tEOmQiL/Ra12qsQnkU5YKhVATojy0Np3pcI4bskRB0QRXLgG9FR/4uHac+SuJVVC+6Wou6q2omu
bMCq5XP2NFSXHPLGkorUaF7CEUz88G8x9FT6cJzMW1bPNN6pVW+1ZhcHCa9ufWK0kEiy8d4U2f2H
0iThGckopKQ/w/1fprKMZnG4Nqjwy839A/jEua+3lC/3YhVmb58DrC0AX8ErurOLtQk+GmlrcjzG
eNljMGWx7q9EqlDx7l9BgLsm7/qrue4LZfuVRCwiMBrXSVekFjBRrXE7Nj6QS/2yhi4Epht0fv+Y
/RlkE+K5ndjNcTAdketaooQMnc8aJKAeKWA1PibOWlN5NvGvk3hpriQmNthxFBIhwPOGlus+Nfz9
J81TZ2aenIh6cg4NkBVTU+gP5pKkpiIw9ygE7uJgh+ouaKR2gO2K7n1RluEp/Os+maxMFDVk6Eti
AODXO0aGVd1QS8o+9cWBWEHnSFzLxdXnhpvDNzBa9pMPxOijIwbd1S1XMkGfAJywrpntqOTGZOAc
9mv6Wggt74dqRkflzypXOWPGKWYDqSINqqEMpVa3whaJ5rTSAW1DhF3KaB5GqvIiad+jHhIrwhXE
9SAZY325wlMAvVTRDyMs71YMzuFrvFH3dsqbVsEzGvOYqstuBOuJJEv3DCCYmqFQX32lsYXo0xlQ
YpxSsfeWF20c2QdIQ1ZchBwbnDdEc0KxY6TcdhLC0fEz0X1IviUzPplPWdZyIAeyDJpcAg2Gs9Ah
6LvdUXqsuZvGReyQ7gNrZNzQzeshFkfDcV7aBw2Vpa4M0R2/8eoTqvL8sI67TVXOmtIJnhie0mrh
USePftpll290X8gUKz3jDQnp7zCc6LtWmkDpAM1RogHoy3zKN8GEIIbzGdOMmgP3TISecpozrOHL
eZuU/CbuLPEwvqu3Wvfb3/V1UjCpTuuvnlxDqlf9oTtRSvDbkds8thCOONx9oxyJeyAuXlCRyx4X
3sw2Jh5k/VrYWjY3Y+SalXov/+z3SmHvkPyPGJK8zq6J5RyxetZi+EBeivbUd77Mogh8/lA7x1Bg
McWGUA+DLzmuncdrk8qVS0hDcCFOKxr+yUBl6tFOWBKpk+O7DxzbcwVTv3Q/AqF80QofNWMPN0Jt
PZ/Nc7btXJqhkwSyi+in2ZzL/FAZCqS2LeXITudrJstZnIAd85j3CU4b6pBomG1VI2RtLuay52Ca
vb+KhloFqEj7rz7sJgshTnZaMMGiUKmWtiI2JhLgGHPpAqORgbyXHkDCjT003i9GMiODbwuwK9kx
40M0rYfRiXYHvRBx18Nzg1LX/cRMYEuOQA727vtnMdYGI0k2NM4/TteVeFfboNTuIqfseVFGYVjt
lxECvBFTXJ9tJOR61G4SjqnfmiBHvB2ilZ45Vga81sl9uEQ2zoSZ7mHnkxfVtADeMD52qEJEM8kz
pQ8/+im3sH9vwKg+UqxHaZpiMo3jLLuMdNFvPvSMlvLokMTseUMUsBHlfoJBk0Yk7128JeGx6spz
nu/IsjPDdbNFxz/lKwaAOjVEZViflssX3RSKuGS46mA6YbVjnoQL90jncyUgQtSNVf/DOvpWedVG
D76W32snJgsVX/cuJy4MkBHhLGtkMV3JOq2urcb78PdRO2FEpIbLKOGPYCj/HobXz9Z3JGnhLT+4
U8yCuNMNAYDxb07xSqtEKE15V0h6lKiubvr+OrpHyiH6eK/jrLSo6hUb/+rqGdyy8WRTGwscbbv8
DnWCzFPcy5i+QUbcC/cwBIgCnqYOTbCbcqDX0iX4397ctpySQu+AeJXWEN1o5C8OrgyxTRM+qozS
3s6W0mCjCxk4nCB3nfvD6/IVFbhdQjoSLo8+XbDxLQuan7pe4RMeK1iTgM/h7HmH09x+/r5878No
+L8RB1eelzB0zSfk3FneivnFxCtnutfOZm2itGOPj+EROZl4FilRDTNYE4AZDcxmIQ/Izx/2+pnu
+iDvOSihtDIHzVVP40sJ/ercfSHLux/fdlTIM+xStJtdx9nnJlqWW4Hr7lw5/trCvDk6UhE8nNLz
kaRVMWVjWxgED+1YEGr/Cbd5UhJQfi5ZajZQbYftqMNHEOW444GXzBPD/FMQamTK1j8EIOr/DTFf
hepSAvExVAf6OguT8IGDh4RmhH+2fdhWped0pQ3bwiO7Z+sOIXJcLGeam4tC9kKOK2oPy0eLtyVT
AM+sALq8FraNJVn2TDtzjO+H9+fI7+BPdBTBrsf34gAO9Fjja7PcY2kKEnvQNOP1o1Ms4USV5Pm5
oYu6EJKyOCR9w1348LmLxeQVD0kMx5mOp+3hojQOA5gYJzI3aqbjQjuuBCzvrLhF3UfId0j3FKF9
THah9o1kbPUf0LCVfRuyVFc3LZcraReo1GJy09+llYI7+xAUyWRS6fuPl8inadf50eanJ1iY1RUu
12eUBPXqdkkSd8/QjZc7YODRMqQmRgQ18MHuR/9CI8vxzfJW0RtwvK/DgdosEr+ml8FFGgAWKOMJ
5c7gA6odJ88LT6oxNSdOC51Yz4sMYSJF1u/j2TmJ82nfkOuSlZ+GICPXhIFcvLB+ce1ihJCR+noF
f8LaOj1ymzUorn4qKHVyx5CdhWc31IrCMIRD1Qlx/OSCY935GKl91XavUSsZc4VmcGR3+rkmniFF
quDtG0v+/oZXasjd5aMdt6MaLCPlWd7okYhyyA5HGnJl+qvTLjPgBHYCxnzfYCbAy2Dq3HT/lz9j
1JR+yIs22+0I64dYUA+N1T3x4E0TbtVxSLk8D8Q/+EcG1n/deUzIbrLmOF6CPrTAXakrkahRjiJc
bY3j1qSUNpeStpcQMhm0ar9XaQag+k/xD8/kQhof/05h30jG4XBbhRGBNftxqpokKpbRYN1Mc5mg
zkFOxGcYqktlZhtas4WgnKeM9u8USVC9tRA5gNs/lgdUW87b31Z+oKtfOMNCjJlAFNl8aizeN36v
PRO/0rdoMBmuRqtxV9ruOBIlKmcrFm8l7WnPJrRKwdRHkih+xe1r9k0vZ5M7qFLJhvb4j979D1IJ
TXUUctY01bWVk5PK2sX16Qk04DmkMN74FBBRAoHbJOEA3SCuXoLSJi3IzFm502561A2gNxz0TFuk
ySyltc+uo359JNvgeOkVwFxDNjAhv3+Ko5xTXDQ32coe9+ZVIeySH8LgQUMwYePUOt2ZvzcPwl4s
J2kTAmyTEBz71C1pIeXF9+5HY76GiU+nykc6rgCC6LW3Q56Q4HBnvu1xmKM0cKQwcK+YTr7jb/d/
5cxFfYH3ELxuJHP62YufGPKwfY9GPr8xM4i40lD6EctlgeXrk9G6JT5AozLrLev6KRK8t7YST5Lk
G3rLSpSYjoi348AaDViuoiKBY8g+xwOfVx1klCEfg89EiYHF9VL00kmR8pXIPDrdTjJTBYGZNMxj
Fjh/U/UcMxVbJGFI29Cynjj9NmEpWUQUF98Q+1E/QSPC6MlB8Z5Ab7chUcbqTpZ8w1T4ys2mTN/1
K9ROeycK+rSFzu6Ul0Zs1LVt1GL2ETs47LZSVs2nhSXsYYzAtiCFM9JUPftkttDnXRZ0i5IjqMWM
G6OCwNKTu5ScMCqbB9IIgZCexy/raBTbyR0sRuHmyRTJmHCXg8Nl2j6EF/hQKJnV57gM5ocUenVe
8md6hakxWDcEAPxrVmHCE2KBgSLSrd91YbIJjhmnpZ9iSjJDtjBHqXe95NpY7MqhxEyquQKAgZiN
2n9umENLdhAypOTTUflKxaqbfvJVfvzFkWuiDmx7EPHQ8MuGpZe1adv/LPGgWds6a0ylvNcfswK8
Oj+OWBd1WX7Rw1E3dVww7E5FKA7zo5/C/tzrdE2utJyUG0XM1HsYyu8BkWUG5j9ROEtMzVV6KMgg
LOL7o/ELoJgJ4BibVWhfICXUIkbH7zkhWglYqhMJlyJgnMWPqdBXp83fwIymYMx0M2FINt5iDVbG
wpE584mDXPZ3wqJziz0B+87n076mO4ANgUV2cdMP6pyLF3N3+PiZ7mB05FuVzFW3JY++YnTySYFx
OIILbYdwREmbFRbj4qPHiJNodEBDXTya1vj5u0Y1FlpTZpmZ+vGpv3VerlPzGASNVf8fZtczVz09
fKWj8Qjr/cHxstM7UpWKvZr1f7yODHMPBmoTwOTdJc0zfQTFvGipOMmiO1Fb7BK1NLrfORzNgZCI
NaVM8r3x+ocUsuSNd80En2apd5Q0NvDFdqsVP79oYdHL2GsYEcrVf+N/pqioe5XJiulErM6pnWyg
xtW3UqrDOydOBbHGHM314tQcYPPWaAOW7PRxcjUbwoGvs4ME6wRDEK99ccprGIw5wv8k6gD3NfVy
XptullcRCETdi/UoKHm3P7/zgL/rUc/hVC28EH9Xiqxtb5j2zYXv+D17rAXQRAZbPlvlUDIQR6Y+
vYcRoOpJVODk0z3qFNORrv5WwLcCnfHuk9+LS4NLzGIao7mTg7gIwoYOcrKbp4FkcYcs+hU4y+En
zgi9ZcrRbLoKRzFX+HEkN32MCI9SOiRaA5bRZJosYBfa4u6M6iJoXumfXEae63sTBozhTXGUz+oA
kI4hoUyAef9PUSouD6jvwCCZDIWuevn4Nax5e6k88Uk7HY5sFBj0a2oTxxduN0vFj5zXtANNgFux
pi/oAVZ7zmPBajZNZWR91T3tNblTQ3GNAxTPKiR9QfRFFVs90C1pSP+B0hjYnYQWETZV7Apjfe8Y
1AK/tlnBcUx46+ZrjS6x/g7FhH6GRziKd4ExyjHntCra6OFl5YFeXrvVB9BJBN0cHtR44l/rh2v8
sRCGYS8V1nzS520wD3KBPqoDAqQwZeHN23Azqk6QfGB3y1PpO+eWpIlDezD90BjXtoVKWSOf1Plz
X7XQMnmfAZTeb77WQ0Tk9/MFf6wr78kZzq+B7BPGy6IG9rgFymB6Yhtxshd15np3/6VBsDeg0DGt
kya9PZa71rWZCAHAqZSLFKdMfBNX7v3/zaqhUXHFMVO9rhQuVm9IScNHUmQCDdihbk/MXbtMIsZx
g/mJTfIBsoty2b1v8l0OqLYVxFNGzUYGEip+GoJs8EJkeu4Amr71LI5fsBIFrWzTyVeRRrFfopyj
IaEK6BI8PB+kc8Y7F49D1ueSumrH516czsr8lh/9uLMDggzIr4TZUO+nVstiOOBEgItS+1miHplG
JxDFphN2VYbDU4H24H5bnZrcrk8olobfcMDYEVyNQx1lqerHZhwovohHjFwckbx1oZGU9UAQbbyt
aIHj/iajl8ev4J078kBTl3DWC+5eh1Cx+/j7izryKeMhzIDVrskMGNy+Sxaewr3IxJLSlQ1zI3IR
SbxEvnBNhEhBX6ZazMOpJ2uSxdcSVtP7lGac7+h/hAFAMH+dYaeZNYQpXCddKNi2ZsnFHNqHWB/Z
rBQekSGtCxrhEkvFtpDsIHehJqL6lDhOzVzMDA1h+2iZxh//B8Y1YEh3zIuF9Ihz9ro8fZqEleYB
7EGY69C4Y82T+PtU9lfemKWaIqxXHwaMwlcdNom6pKxYLmLvZN3MC7TILC2FjaJBdjUsXBg30Obu
qn2DCg7vTE52xy+B/0yMByCC3xfBu49PhjraFDqZw0OmyihG14X5F6hLxu2tSbyj2IC0nyisOou6
FHWprpEyaqbSfF+9FNQFLKYQSknUchr1bJ8oys3RdCAGpA/92CNoH62+DYMHZgxACHPzhVmN8qKh
LteSNKuEvidyusovHizuYwEPUBSDjR2h74FD+Cb/P6FpL0XtZFaNYHUqICK0VkGazoQxuDzQfS2l
CqPxuaDikVYPBB2OLaxaK5hzPax+m0hazsEfG32rYdhn0n+sWwksNr7rR7JvEyAFarlUtpTYsOHa
i7Yfq6HjsP/NnxrpubpGsKeCRuoVfVShBmTi1K9iJNAlfKESWvBHpl/cKxBsBSL7xT3YvVDGrfCS
Mherl6lFJoUgR+FIlLIBYARJYLK+8+Ti1ByRl32nQwUUpmOfSUfeiGOt6V5xDi/NBHGPc1vYi30v
a7HfgVa64WDgyt7caKnfZEWOQueNeIPiz7VkZy99n16t8QccmQZf3hTg1KFp/WAylpZEyyPC0WS5
bqcLSQVUK0eamibSN++Vj6eNfSnKj6GRw0I7uo4YKXxOA3H1sVT7IURLuDWOq5OVMaw9Ygkf/IDq
YkFBe4+AlcBUYRLkZCvoezWuan+WGSMhoaiJHonxFd7KcJhvDDxG4IxlVBCzO33zWKZA0KPmB4I7
y4K4/JmvyGCP5VjA8on+Ss3hpNnzTBibvnTKlXac/oTORTwJxp5M2h5Q0le44109aoGWeGn5xNPn
Qjli/RKIsCIdcNqCR8yfIu/vdttkkfpVFEOE9NEPAd2qtYhPSXPaxFw1Ebr9t3nhhvyTbM5ltXVO
hn40RzlSmOYBSVZTOzpaahSFvvm+fmmELOzkptrF53/LkUQoxbYYdZTMkGMQ+mXw5DvMKNfKDiu8
ar48zHeadhTGj+lCkYvsRYyM7qUryzT/LHlEQuK4PKxwpG/2ahTAVj+bgaQJCahSqSEuzTu76CX4
ltk4k7YmLmwIefBvEZBHggY+8KOxzI+u3rmt1oQ9+aon6WuRlVfsPRTDzIuw9zxt4nYBSxMqPifH
U9Yb8tGTxSke0LwEcwhDIrj9SICaAAoqFTp9UoZpAO73SnnAjNQ5MPFPe7pnZBtbczrw902Z/Frh
szn8FnJ0ejFPAGvFlm8pz1fkBhYweFixfIga8hWmI5bxuMX9TGt2wNV6N6Sc1gM0CopEA+rH0OEo
thgd8ZBCUyhQno6D8/bXOt2MJ8pNb1OMQVTob+4lbJPCKpPR3hPaBMsYB593NYcKR0Lc/kgPSrqj
/TmonJ8lqrdD+Q88cbAtqQN5NI4r/BOZCsBtqU9d/NTgD6Jx6RCPQGqfADQma8il/QlgCPD05E9I
mmK8QyEhi1j5VRK+gcFFID0+5FsgD2PvsIwP7RmwexEsCmCmDeFqyYJ6GJOqxDKF+dwSXpm8Etup
oksJKWN00u2UdY2f9yjXqE2s2bFUisc88gsiG4FWfRFVSay/mWQXKg3eIlPBkv4DWDA2CKqHO9g3
n8T0DXaYmumztIWsfQjVh8GqNj3LKqSpdlUzZ+ksNu35aiYxettZYVMY1HUVSu9+0rz2JqvyyeCn
ObEk4l4g0DN1cmhjMV7eBC2YQSKSPrJ+jsvHo+IX4rUOwJSnG/3zwycop6inIc1hTgNnY7UbiGpl
KCGV3cp9cZUva0NjGM4vzxpF37GVZrgdB4f/+QfCOQGGTMcWL1i0dJl8eNRxclXsDjl1rRT4G6Fu
mx/l37YIzMkt63jazAnNIKi1MO/q1ML8niD8xyJPgrt7VJxO0H4Zynfogxyq2JDkdOYnFku9yshS
yPUo1ifcyS6J0f441s73x04iC1Sl0huU8eaA4v5OUyI5XufDdElPVQSgl/I8JbxvM/YINcUCocVb
YjftrvTTPPHisKWCtxN2sszmU5JeApJ8hDPx8WWBMa7aeWjEEc62wF3HJSFh+rs0IXR7bWY76GSV
irgLa56meFMIeWaC4mOl9c7CBzzHU28lNJjl0zkp3hTsKO6n2HbbS1IDX//3Lbvq/dbybjU7mx4a
YUoEoqAjXtlNHr/WVRVuES/HuMR6nVAr0tAk+dtEkI1cOudn0VMIuewD7h4q6gacQ9IfTPWt8Ejh
mB+1W0ukB2R+wJxI0G8fl98BBqDr45xoeI9kw+SWAVvkL7/U5LkY2kBc+OAXiObvpcliIw4ptaW4
KlLQSmVbAAq9Q3uFSalwvWhXUXrqVmwOX2ew5P+vmbxLYN9KSb9ptHSC3g8koUS0uFU4A/33CRjB
lKdlmAjj3vAhqKziV8+N5wIfaTmVngr1upUK2BxvzhlXQiKDJNZsCpGyGhA+ceS2qNkPR8v5MPhs
hwhZOIm1ibM+e+oIs3uZGTLH2+XdDWR1w4oQ2wqr4ZRC3FVOTd+uS7NEMPl3TnYOPf1jYzZuWMWa
U2jQ75ubKCj4FhEaiCm3LdrLe1bcBsGHv/uNKG5907E294MpDJlGhZR1v0UmnIhr6a7wmG3OlFDM
dJWoevdi5XxIQrO7PplM5qoFJVLV09SSPr6mO1wH9zCFBHWSkQTro0nycVP5ZgMwh/VosGKF6wpx
BKeNi7oqJVmoFlqhao5nDsdjz6IRGE2Fa8dxr0oEIJcLIpMrYraFFnUn/4iZHsGwNK5IfemJWHCz
l++AblnvxDRLaQd4tZmHIewNYmI4EuddIhQGVOaFb+BBh5GmKKNNsbvr+qQI2JPRuMypQqssrpD0
I20L4QMPWEr4kg9JFzrU5/uekPnx8qmenLKnrFxByknMPVJnIZXRjDpUyT92V48rJcHvQb6eUkQd
FIkAKoguLulZzWibj9vOCjCwhx4UiS/plPAe7daSwmWfeDv/mwd8vGhiquSjYfvSw0fOmXPOwmax
m7RY2499S4m6aa+hq3XvNiLzQtH2NRAlVkqoTLkqnn0YMpIRZILB5GNQMpQLzal7Wl2yKfzz3Kyo
677PY4afg39OUGBXTCZiRbKC9wmJmbLuFb6X+OnVg/7HhHoupwUG2IHR5r2znmcle6BY6TLjd5KW
R7YA5t1Rt7WRY5WiKPicf6rw3lVO3K6iksb7ANOt9QmVj9ZDeIHZHVtmGNA0jqM0WclE7Z1IZguR
nhh0P08Wx8alh7Ihpt98+U8+vfhpZMLDeG7ihCt3RbUBVX6Qj0PMcCm9/iiIMsTOgHPDOF160ykM
IBJqLXV1x+emlke7h3zV5iJipfv4gXFxhXTgA70j3AgAa6QKCk3hg7uLhQGkREuy0sv0etWLBgjv
Sf5kySbQtJx2EmFk/PXU5/XBYbb/cYwBvb3eHwtaNmE+FzIHZYYuPP9DenkEOPUtBA4jSv1e43hN
7bKAWEMseppBsGI78VC8pBuI2rtZU7jo0S/lNADjPORPUUEa5n5wVirvYUe/l6kQCKxVpL7mvNpS
vJ4XAWykZMiLZtbaCEOemPoObFCrsPve7Tvl3s0cny0XteP2jk2KTHwUB9UnSAsNh7d/VDdG7u0z
wiNTU5l2KKSQJEw4037OYbxZeHXHVTGDrHAZTUkD3bkRFLlsI/9Hxw/wPxMtvOxDz0fVxUu8kNBB
sNG+QO8aSBihznzamjGzl3HzJlTmsDrvxll/ikZJvrHW0sp8LlhRarrs5ZPz0UtV+3tzmkWoBthq
3lrpTBZMToYcmI61PziSGmQMvn7PtujC7migEETfdyQ1e8CqMvvTsEFBscilkTK7Xh6/M0gSheGx
MWE9V7Cd2haA07bjC2MQe5QxbkheYw9L4aQNNBg9JTgKXbfuAqN2clw82zfMOOqesBcsLEMm1l05
OGi1f5CIm3nYcxj04NjmYtHHKI02bV51xsOSb1HhOvg7nyJKmz3PqY7nAEf0gqwGaY/x4LI9YwS0
rCtktuA4OZZF2v0SQ8GQe0Wpvuo6CMZhJ//Imz8FfCJS//pcWNbEpEOUZ2JwCJkc0EqtI7ic8YQg
9aca4fnaMg2ODX3XNNI9MlUz/7qzj7ZPyCDcSwvesdFCKB7p2Ee5ehFtbTX6DhYqjWOBkvFWqeSo
1/adeXhCqwTEH88JEQntSUplH9sGLPtzZJjfbHGU1gOFrfbBVrLAvd6uc5NvURKwkmHB8eS05sqy
ER6emQjUW1hj0ubim6ebnBK5lkElXn+5hb/SYmDEmIU+H2SFR11iKMmCbktWYDN0DBh0+80SbNND
SdAVN2QgCnwEDiWE8uJ3Z4Zj2/w/X/C1SBKMWn8J9+nb7dGhqvleBWOLff2VQwLno2WUZzQ+pzPj
DA5WUhEYs0e+4G07jld8AxXq0qn58F3bOfOqxCvuhinbRsQmBnqMl/l3DVjMZ+jJuMtYv6jwFTQe
tgu0CGrfAfXY2tZF9jo35oasYMYz078Y6oPc47rzUwg/F8DDZoyboo/6qMWhb8A5p1GaTDcxcJ6z
Pb6ClBKK2O2jJq0ZVvBTXV+E4dEVJ4KXidIHe5glnIi/hlXLd3TTy8dN3KRQQiILE+FBSFYXPbok
IOcgY+ZlQtTuW/P06Q5PT4p4ZBXifeu//EqJv7cPFALC8BL9iDnuqLsE9YSeVcJqjKMUxIqMkQIL
iC+Wb4R4AReE6N7ViNm1yYvRl9HSvtgqlMiemq7Z+VAs1eXR78ljskG0ymesQfsjcxdlBjejaIyA
z42hNw2EDlgZY8MlbEYSAbSfJCKYdpkXL0PjT0l4vJFg7gLTJH+Rkl6/Jl1oM2U9GIIpcPqguVU4
taBXEY4zl0uB6IUOa4bhSEgADqSprp66CNNv1XKgK+tMnm2UDSJiMNE8UgUUedDry+KLs3wvym6V
ECMYyVAISe7fuN/KS/nGC9KspUaahOdM7oUPgc4qwGePLBnQeZgEbuwLZu6Kf7jB+xYSZE2Z1pnP
384u9SCc2hab8oFFaf9NiGNtP6NG7cyXt7yVbyt4FLwTovm0OYZISP9RqlinVQPS+aSDB86wkuMn
VMb2vrGKCzrRvgmNvcE9Ps9UFrR+7tO3HIy+Yp87X/6SmWtgiH6rj6SzWTHAei0Q47SUTYoUmCEw
FiTYEUkuSgJbA1AU8SMYjkRekuZ8N+vtrXBqIqomMl49VoYSTrOgdvjMpb67oeSvgcGhdZRdlvTz
BxaAWBlvGSHUHgMDg/5l4eGnMj/JG8IIlp3ClYJAZ3cvVwU7XZOGoxFvvDNAW0pVYqBRXkHBA8u8
liBC5rOqCNpfHt547CCju5zms5r8VnxSWFw6+2AbHm2iQa7MG1mYyRPPzXH9CFtI1YPTbL0b9PGK
agBGeTxFWFwdmnA+YJel0T8cPEw6JTuPZArOv1KVQ2MWHfznFQexKowfR1Abt6SkhhxjPn6iflEC
pjL3/P2Lij3O487xjfM1t4Hn+UZeCxcpMVSVytxdii9WLQjhs41hwsYPdi33ZiZtcTgmvlMvJgyr
2gP470i896PEDY/aBhcvTnnSQrxo9Q53T44N2mrcy1NF7/5bnAB3IXI2nQQULaFUhkwmYjJNABxA
jQBueKVeF2sxJkny0IITQ//pTv+cccaBXwmmOS0VpdboX7wpuat7xy5P+AsRmtkd9ZxNNBEdyJbV
7s0MOd7LssBno9Cc44paA7EdAU5ar175IvYtHnppmteAGmn95tpp3VDk56ZIVQ0GYwW/3LLiOQ43
5Ijsp3mMP/4ZyQ3cfZ4+x/XMq4b/Kw2yWQLMsumdzlbRFq/ZanZDiCg5K2ffkPMbnt3trhnYLd+o
leiBPbAkLOkYrknDUYHtxIHxYaEYW4aIoarl4tyztQQZwuCMOtHYo1+gw/gZ1FmwjpnuW4xXgdep
x3DCbEkXm+1r8hqgEkc/zc2RI4e7tS0sZLB5GMoSehqsJbq1FoPd+BskjW2nm2m98Lq2hwutxKyq
+DoWK7R6FwCq8YKOW/QomARm2ACnwmfwZ2hxo396GX2qSEQT0naiW+HrRTvUD+633ZsLN2AKtRGk
e+rbt5bQ4MJ//3jdSjzBjylA0xuCC1cH8nbAg8R9eIwoHQ0ZQRQFDNH5+ym1gcPQnGxX9TOROUQf
MpxLLA8OkkeRi/1dlqAIAvtREhl8aleptYAhqxmURfW1PwxLhjDyelUcf54IyPI3SR8lC9Xpo+mc
76vS63edOpB8MAZhOy6abb7JPsBnXst55qIcN4bshl5lG3MwzVyaVwvgc9vVw6ZAzSHnp0Ue+W3j
S+Xvy/MKnIWtdEHXFbRHatzPS5deRULzzBGElaoBIqwe2VUlGF0V1nBIX0jkEFgCT+aVXCzYCp/0
mU1udpC4PzKMo4FtqoxkExRYqJcIOqfIQ72qh6S6twDTILAKykAaWTkOM1VEVlPGJdlGsYi/IZ7L
vgJCsR+Sqbk1LVr+u3itCoVMe5DUkvTXgvQboPtVZp0xsVREHvbFhqJKdlJc271lOo+ihnICRnp1
HMF+2x8iddX7zcyMYhr/UNG2AX/Jnj1tMlOhDSoSL5eGolreC1yg7lDC9ipwhbf7IYOJhhxcihn0
95e2Kj1G9Mmi5+L8JSlDS5hcAkOxmon3uPnMRpMU7WEE4J7vxibDZfTpWFamiZJPbT0I+Sd/q5ET
lhpGq4UFmOF0SifRa1FswV4ceYZsVHBkAI4sby9yHdhgOZcHFQYakcoamkH+gBKxWu6XO4sT2ph9
VCYsY0v7OFwVASF/B6IJ7dxM86Bc96lk8juWq2D9s30IcnO4aLcp4XhVlEKBYk7NhnE3hzZsFmJX
J2yfTEve336gWLhG1LK7uvyJQBVMJE9TcBjmI28wpWb1l9UYW/Ld4LyGOq6WCWcWUKB32u+ugPK9
oMXGVpbJ2BOK8p8ki0dzDqGU8SlVtZcnymwrSN/bsBpHIcUuyd4dzVKZdgaHQH7F+9wdyXzmf+AW
1bB8OtaR7nzN6Vit/gq8Fx2G/4uuXj1+NUoFRW23fjlbGVVqwZ7Xr2wZccNh6X0WM1PkczpubVhi
RZcoV/7VpUusRAWfZ5OdR/cePiOQu4P3hj+RCOknHjGGPwD2ypNzrB/GGjhTKtYEQhFpUHSz2tW7
GAxEpSz+YIi5bhqrFGHnY2E+Nx/JvRshVxfznr2X39D2HTt6riGLugschWB1SCSw+/Yt9/eHAlPg
vlVaa7SKhUD/61DgN9oo5UHuNazXZ6B0o2RmSgji/tC3Zzh/TmdSUAOtTb6xVU8ExjDNtCJ9lkaY
SjggioW8Vk+UysDFpqU1qDNsCegsOEjHHUPy2QfZtTNDpEzC4Z1FxexzX++zdP+Pe9HpNkXUe9Sw
IpULyZKMVkALWFci7lneWTzFrOwCGWwkyNv5QYUj4RPAvQnYYaIQKmJ61qw5X24O8sT4ruGDh9Yv
0jhtljaiMeEKQ5UYYVUYPu4lW5YnX3imnWmi3Js1RUOyDBLYo6V3l30fcX80+wAzuK9V3vC0py5w
EIg8nsE8iLEDfcD2SuznZh85rmXSm39xghUD5GOehYvnC6pxa3m6zAbGM4Z9f/ihrPfBuslOMPpr
stO8RfWZFc/whn9K9tX7dVv01FSy4Trx2GCrRkAUF6HRfGZDHvhwkUfreCIrensnkQj4GnFB7Q/J
LE1yhamjR/+raQVpR9a9d7ZUO49nUQN0Jz+cUXJta5SLuuXLYH2dkZHilKYExlzNbq15ndA48+o6
WvjddByipWnCBtkhw+wGLYL02rwk727kpJVgnOtckMatRQEL3WHwHXSKh7XabmR+mqBqR7Rz7y8g
haRxxas38UyUyrnjggdRbqLKow0jr+CJiZZJTUcHIzV7U1Rx3Xohf8d8a+U7PUJEs5HG7jIpn8O2
IjCFlugnLzaKRu0v9ZEGLoQCAB0+GWiibVBF951depc8RXlmZUU3w/vJnCOCHof+YrILiIxEDA5c
YGWz/SmgmFVevsakZy+3DfsjLQpPx2OZD5Di7UE4dC5eGA8xKvhhidHiBKrq3eDFsvI1NZrcBHCs
LW0QH/zaE2xOHFdKvPpVCPBBjMMeSg0nzPtuw1t47W8rYTqSLSd8DRrW0mUl4xQNFfUj2GVnYkfD
Uo3JJB1AihsvcglT1caTbJZgMXIR4BRel+eiK6VJbgiTTCSkhVR4HPT2Dn3h5+btVAntlryNSDj2
0Lj/xGpS1UuQBsiyy+uNaG0/zjbYSdLXuIEBx2sdMFh4JX/InEUSpnK+fAkSdSVXBbRywyuUy04n
fMjgVwHnMBt3xuM0DbJMrF199FbZpEaXXMbOZfOCFxowg2Io09ubD6gXj2zvkrBVtg0OIMaBU7hl
fB8dM+CZaiv3poSqFhfNBois3aU6w8gLZc2sC8HqP62EV1ry2vJEl8KUx2bussSN4dQkmoDwMEi+
5mhyjABRXRQzFX6aLapdgytSq/890g2R0LBvMJAcYe7hM7UUHrw1qOyQ+CEdcyBTCW7PdSUMgCwI
J87S8B3fbzEDCObWvc/1ZT5K8DqKVXqI1DpXJLWFFkuxFSgN5UKF2nhjqxvKZ2bWIuIn7+SRmxQH
y5c0oMKzStKBCF6LqVJ01KQN34gwB/N2lsMaEUU/NqOexckPF9/992IddwjM2pTfwDR8Axe7maNl
Dx2WwBDzAfBOwNtkv9M5eGj9HNga26TCvLQ3kM9aQjQ8++hw3Dsqa2njAA+Z/h4+pgDwEs6Q5XEt
0gw+zKE5J4NedlQv8pmMmvg6+cVpmw4CbqPZboHoZtVQhA5tnE/5o560VCpqOrG97JMR9NJf0GwV
67y7zFUPWqE75WHbcY91b/wh2ERm7dghUdBPNMbZ5ykv3cg56wQlZfOUAnp5DummLhX+vkiDycEn
/LPgzo/TQhNiTqo/n+vjftlI812UscbnLuQg3YuBRXQpJfBcEjn0tW4znJ8gDzyUT2yKoaIlfCj9
apq7gWn90cx1bilp7UndDw61YysLVXyv+0nc9rOY9DXhIFpGPQykxdlVKE4iwMmpNTI7pJhcnuAA
1wvn0XaXgU52UIqhY2LHYkByMgX/aMKn/rM5Dds9YmxERVsqbb07pxiYCuy78LrRo2gS8i32lBxK
VP0Z3LnFFXFRmN84KmUdhSAccsbn4VFLAuMV1MDPZEH0VpQJsvsBFkHpAuzqcXp0o1WLW6Q0CnHA
z0aqdYwtO2sjKr9rkFAuvT5kf2iaXLi6nnF+W5ESCCh6khAhUOrh6bQKC4B9MgM10iZ/ZHOiuynC
Raz7mpv1g++4FH8vZQ888NJMKp4AQN3HRPTFoi7ej2xQUEEw2C5LMBu4DEKrLSfRZMPBNQVgBsP2
pDbms1smCqqF/DI+AFTOjuI7etb0jjdCdhOcX4SeXNSDfea01sa4eZMAHfJ6BPoclS5OentQShzp
5x2nwU5oQTH5vyULjsL0EbWf3KVLeeZvxXUS8CkCnINxTmB/1xZW0Gq8lXpHw8IVFskFYjMxAwMg
dh1pAtLKgVO2tnQCW6QY1qWH69r/g9yNS10awQh2jnSGERptccG1yzlDsRvmeF26ecJVGaBk7GwP
xkjScQaMOG9PQh0vFHDWrOw+wGBPmKDm2kICt3sNAOM6SP65grZSzGx0Blmdzxy8rdRfRhW2StLj
Dxwak+zx/0Yta0g+xfVXISUcJh+43GnUtYSS0y2OGKjmshQuH8PNJalXxR7BugoaJnlDqY7LuwjS
LobmLY+0zYUgjsYKbjPG6mSpbLSZpSL+KeUYXar0SLkYMxYpSmwWtI3RPM3gLRFoK7ZIszHrg71N
BHnRZVa+KJnPi00qmEKW/AaZgWTADQfo51B8Mu7EvD6qvqKHhe8evsN10WZuVZx4iGehup4gkoJC
b0c0yk3SPXtYzryLhB90fdQR9FHsW34ILAsO3UQRFwUkTbk+YokdYeKw6TN8EsiP1g/I4XiJFUCN
lxJxY7OU1j+ceasy7gREO8iFgwKt78d1tuKdc90lEBAu0M5d7z3a5RKJfvakNsIX6p2IRtqkL11z
EVv3tLZJby8SdOeouLc0RKbJ1OHlXZ7W3WBicLT1qK1YOLvQjaJWvb5T13RfJp09ltW7sW5rCu09
XDzyCENeFLGgzqMz8WGgVq5KLBV5UgueR9faN7u2a/vEjpRaJwYbCHpljez7mMwSKnKwu57HEBLq
Qh0ECsmKXGtmh0SABGt37aIpaWNkGSWgIXsvrRMl/YfrZJrosGvD0Hym1SiNZE1rxCETCPPRijCg
ZMI993TSQmZeH2K8FNUJtSB+sappxeS7hBTewOjI5s2VJ++Ds0OSwwNBw46NIgCiptiJ5BiRPln1
TD5JZzO+Yhxw/jT0oW9DgdC7lutCFJC7qeFzqVrvn+ExU1jLrOpQ+L5oiMy+WpWWaGE6oUfZvKeQ
WPV7GLXOc2+3mmDjjslDUUpp8YsBL0c6pAdnUBBO9sCEwvPAVX2Wvvuu3uvFPozTvmoT+oxBq6zO
1IWsEP3jKs+ni47CVQ18HVazBlijHLltR58JUU4NZHgj+i05cEMn9oVsNO34GHfrBFziL9BnKUTY
XZHvSsEg8ITI5enN4AiIjhnuWT+VGmHEqU315tARM1FI6SZubinilLvt2gpuuXnkrsZbql69xsoF
lb/vCMzbMwnotXB1zezUwYTG9uEkbt78JHG86qF342pVbNXX/t8j+m9Vk0v0JOQLxOhUcRe9otPX
H7B4lU+zPG6mC7L38v0Yp5WGyuMdxWlW0HNHMF1d5obwn07DHBbEffKCp6lBIwiDd0wd0IK6YflX
S/It5ZW1zbgy0zEIx11Fkxd9/Vq+nrUb2Z4p+IbKzD5gTkfn/SRtgpgL5O41zHSB9ej57wI4lF++
BzJf5U1GYHZuHHzgJMbQra3eRfX2i+DfDjem8gB48I0H8uz9YswJyNo1M4OYcwElZxpCne7uRNyS
XeKxPqJtkwFqMtQzki7NhnGGo1Cf62j4miZG3KnKNDG5aRiph3tObRI0li+Al80526VZj0ouxINa
LK0lJHBorbzd4R6ZGGdzuJYuNEeRNDMd+3yImJm7/FumI7xGbF80QMgf8P08hisgAzWls+w4Oxnz
kqLEjEkj4m/JN+/MJPrMBWHAQst43Ll+cJlA2jRK/XN+jWbYKNuZB1Oh0F01eJ2Ns3p2DA/GNiqa
iLh/efSh+/JjR1hhM9xsQQ7SQsO/lfpid5hhISDuhTy8FZ1wrupbM3wjemuvMRzk5BT7KrG66Q9o
3d953sPRP9QXgtfZ5OTH8gM018vd6p999bCWv2DHFG2m12Q5C8wSMeiIu9cpgNTBlbGY+lsF35hi
GT6vWuFpMbPGn9VgvXbICeW65/4dslOE6ZYirjFMB33mgXSNTW7M2q28od7ggu22Ysnz/scPNSKm
rlYEfPjc4FpxfVlgCABm0b+hpxJ9YchJvK/jQpWCUmH6tzhkOrYXXtTElEkWw5mDgmC+7rN9ny0T
FiuXwGrE//xRkuJe9UKpizm01RXiu1kbulD2VIMgZXDCL6pXj8B2B5ManWYIVC2c+WDmlb5VyTep
VuNKikqTUgkchlLsMR5NrFuWQWeX01hBVqcauVSSEJDIZLoaF3Ikld0Vbz4RG/5HTgRvVos1UlRy
A0XhokOF2VELsvO3VraNXp+G45NxXsgcuxaZmNnejILUORhGyIp7oQ2ACwEpXCbxd3fcZnJbaih6
ThwScedv5FwrF4cTOFMcE1ZtDMs6GmnR2rlYK6jMTsYzZlM3eIA6N17JKV5QN80LNisP9Mb+hTIG
EHN6thGa5Jc2bnpwSuO97T5kQ+CCgsUYYepAdbaFfksnOJ0EkhMmR4noH61phZwRE4tbfkbxyl5m
Z+MpTTeQXFuLtRQNjkMrUy0cTBZX1CmEtxs5ddk0TmwLLhvQ3t1akkiDoeNJoB+fmf9HT8EWh8nl
Vmxsp9ziFNjzOZFnEA3CoeMl4tKbW3SSrce0zyBgFvKpBpr4ubl9/kWeUlywq5N4zYjKIs/H47XD
P4jM6BpX2/GIwg6aLzJknzTbvFW4BXcbbDM2yVaWp6Aif7GIdNAFl+U/Vily0q62XsQZiGsqkP2C
iM7FJXIyXhdrM5Li+nrrmXxSVCPvYn4BI7hlr9SG9LNY5KA0jObPlZPSHfvkj6oevnPwT+fs3PBH
A6LiyUuxC1KpqGTTT3ZpQtA0XJD5xdv1kpop44gmw+PWDpRMvYN5/WTurtWYhIudMqo3uYqJsmIV
hEaVZtvjzAbHcDTs2W+RS8uoLnMuFe1n2AMgEM9AMH2MVbKHBWvlTaHWH0S4o6gg7nFPrw3FRX2f
Rzw/9Vf+m4Wkh/qNBMp4aS5AHp2rKQzCiz49rEuQKul+baA/vFH19Mb4i7vdJjjVqGKJA7+KUJeh
WZis2sBM6i2eCoe66Bb/xbbBcS7Rb63o3X7MsWF7xUHW4HECIYIK9U10XD5adRtb0Xd1wC0LCoeo
5K8lKpSuG7KaIJ7BH9x1SZn+dFzhXHl5A27dApe4rulmrTPYRoLt7yYxpDuugJgSatEykTSCvJfd
dJayXg4uwTWaUci2fwlWqKcXhu7m+5fPAWnx1/b2ebxn0IWeRFto9Nw4zJLMmO5W3kn8TitOT+er
tsgZ2SE8RDHQAOeCrqBIDIC050E/VZ1+fu5Iaxw33iUcGrGKXYJCPeYpR8b/p4+/ucmWpzQ/grkJ
UZQRV270LuexWlFIb1vvccFbjPgNsRqd0EsDjFFJoxXsm6LdJJ9DjvlFOO7Dm1+w3Bdsx8lvFSqU
+t0YDKfCtyISpV1nM7nEY1rYKywo1vl855YzhUwimKF16lYRZqd8G4sZR2hdaadzEmyw6kloQpcN
+6wUyCfGEPbKwuVh9ff+2Z12eXFrf1UqMpHhAKPQRuB589iYrGE5sv9FFxiMcm1dmAjil3026FXJ
G1FiFe91gNfLfcLp6WAqAzsgqkhO8dVM0ufNwf5AXUC9x0iMk6kKaR1xOUUXYbH/JXtV8XDVby7J
1uHVC8aRWMdfiB2ovJDYuZ0JOVS+O+W061TLIKsN0xe5nkkJr3XKZ65Z5P4bXIvHgzXvEM6TmRzu
Tn9TBJhKaGrF24Q317DLyaavrXvzh3yaVpE65q85IhvsFNEe9V4W3CASnzjuIuRdbuw3mk0n8Ga5
BPes31vq/v16PVEaC93hq9YQLx4xF8m89aNO4rwVRbEeW6Z+AEPouHAshNitAWhe8HYox9Xgz8BI
tHcS2PjyF3K6ENwgtnARRKiGT8NETAWssrwy7O0HywPzWtn8XzHY2digobCJNjY0L12vFFJR2sd1
Qm0TBbTE4krjUyaqBl7IZl0Xfcma3u9Zp0NurLuYal/EK1tNMyaGZ8dJvp0MvympnoXrJTBDWFjJ
xzSYi0mCn/F0Cn5Bdt2pSX/S9m+xCVGHOMgolrWB1JTSyaPOmyK5HFePJMxHOFr7OwJxxqhYxKUQ
+vzhBGsRQRHsetkD6rUbMHPp1YyAMSV6+pvn+3fM+CrUGL3jg6/FZktaIUhy6wzYcmcEn/UsHMNs
rPKRWLO5bCUZjXxqmR1n7lKI4yGN+597jXu6AzurBkN7EJrLj1NMH9cKnA8iBI8+HjnKur010jG9
s/EU3Dvxfu1VbuXijgSFSc6kRjcFglXsctprly+XBW+M/OJCRhg5zYPB0BHFG4Qmn9AJF52sCDSe
7Ms+7oI1jxxyuQBgUBmakvczhv/xdKEPyhIQjuWZLZAKLiiYv2jT/ahfW6gg/vHJ8tce37T/BmuC
9DFy4EwPQdCXJ5Kngkcy2Bsm3OcX63LTSODfHYhOQoOtipBuQZEnAKiQzUVCnDi+J4mTj3pHs/ED
JfWVgENWuvDOWJgAQMgXhHTupN3bjhtRcK1l6qKxKlGdkcDV8CmHdsLI61HttcbH444HjMPkCEY/
HPRTTvHr5hDEwXSnik2/z7x2TR+rwaEKPh6gN6Afw7pKsWDc2bykn8J4Mmv8qHqYZ/0k4+OQr7SQ
V9tkm+Z45w8FUiOTcg7rJwsoOun21UMrbceHyKEV6rcmHYlB2PAtogVcJCvF+RTJ/JuBkHsZgLlS
bmzq2OWntPoFb5yRMI7DpqwEUPBlZLN1n0YFlwDeXCVX0tqgD1771jpNUtPfhEpthvT3422rBY6e
5UH8iz0/921UyqEDiDcG8mA12hZpfFmObP11GqtuX6EfDi1OP9Tn/J3S+Sjoy/kARe5hsQ38oy3y
JeTQIotmtZ6UlyzfOPmNXpaZaaMH4s/OpLJpfgLGHSDYXlIcDlt161Ymu+9f8ABiahO89oZTu0u5
opMNyIKwJSc7aiYU2EoZz3hJNrpvosV3F6VT3jlWn6iYFQwU8aJsArI3ozQ1JiVvwiq7NInugnYL
XAOHDWnXmvItQNrKFAn3iqK/7OneeUMG9CEeuvvk9Gy4vdb9vRa5hPS4I9UNulT+vP8uXO5xdisF
KpVU2G4Yzpk9YXCwI27kk5zk2tOh0MCfFsDWKH9i0to+OlRJBuVvXM/S4Zh1EMn5zYTz58Laa63H
40nHspYMqWhmAfTbPYN9y88fAaVvYKYeOApKtXrlJmS4a9qYQx9fC28x8sTTgT39YHHSXLnNLp+q
QwpYCBOpk4y5dGMKnrL8bpmZVwKOqTV84fSS8ebCSQs8Ces0DnS1Dv1Ftni39YSPOFer2fNAczp5
IbyAvakjeA5CkkwsCJX1r4Cq3MRP1fwZK2ox89xWgpTgIYj4N39ju8E2caxbS0Nv09nv+npVRxNP
KHgmLhhZuvcKZ9UGV0PMdJWwaFqy3hTOlXcIDsuYVC8GVgO9dwFK59tHigURASRiQN6mENE3HSsp
hJAXP87WCaU57BUtlYhywXO6JYVx7i7fOlnVO6cZy2fFENFatXIryJ8iFfuw15eE/6lCj73Dq374
q3dNVobs+NyDDzbLyJiifJ2uODlDbfwqxWAOvWXA9LHRS+Fnqb6j3CryPEJDrzXsSsG9FrLnHHKA
/HCXaAI4krhiGvYtNbV9ulpIaQoYwXa1KC2jHBjGTV7ztOL6AKL+jiT4P8J5V5tOHIkyJ0KbnaXY
Dp9jqZaZlSLoyMQHsJM6jhuEa+qjYg8+qoICv5o13AUXtR5RyuLfxkyVXr0Kcr9dgh3KIa2mUkIJ
dB4gGlVjQ8GloCBsng3TIKhuOvNhd7yNay43IsCZEjxHJ/Dl/n/b40ZnSy4aozFZIi0P9iWXNMO0
l9tG5+2kZVmAd0oymoKpqEOdGnWobD322Occ0Wrr61Tg/u/a6ePJdOK02m5QtgGtWgxPQTCi6H6v
xTk527UuKL5K8Lt/Hy4jpbtLU5vEFzVWcT9RQQ1KTylfQyUnyTmetPsMo6XuEep7MngVrW8HeE8E
2WvBTjmO6mH1V4nN8PipurUaoYsHgGUh0E8W3O/LU6jRsDaCKRcaS1WoSQq5DmZ7iAzp71TLVbVD
9sYGJSil98Ygw01w0Op0kFajbMBYzuEPKGOpabaw9BQvJev8o0aS35lWomMdp8lgcCNDC2QNH2lu
0YZWC5mHu8GRoySbmHcwSTUjXbvV8CPk4NTSGXfQqhyYKDKcCorS1NTzJ7sNGILFzds+y4M+xdy7
2c/D2Intjn3e63TbOwolo2b2tqnVvPdmQKBxx47zb0cigvS/eptwzF9vtAjCx5I/SlZjHacfnOCw
txFKlCpKRv9h4TdlnmDJWGvAFY8lTwA/y6saI9EjarGHWdbV7zAfn8aCVgeXxVHWFZpfHbpcCMka
xW1Gmnjmts5h98lKl9scgIWPSK7Om1I/p8dDZmgpBq/227E8rwhxaMM/1BHtJaf3mqnH298U6zF5
JNzUrq4LyVIWhV/+ZssLPHG4Tht+Cc86h9G5+xJ7wxZdqbH7QcQ9+52AyX0jJGwhdoWYGlQ+claH
KdxcmTiBUezSnnmO3Bvm6nbIX5MOFO8sgPzgjza60R/c+RuWfU9Mw4WtP0v8W+7DZzk5l5K+5Hbx
YfsR9sJNS3VFHF6gXoIPFMBQ0TU4Eh75nL9I1GCKhvCJx+f8wG11mBQUFHNMX4PVN4CCrWBog0Kc
/mx3KdcbXLKP6h+covSsBTHhE6G3EjG5pDAkQ2oPjeMatsvONQOC71ZvX94RrBlReJP2Zy/dhDSX
B4cOe2iHkiSQsmlzsA0gIdfGFeh9LYU4VaNx5/4QAHgLDe0TgYN+wA8wcIJ74wZ1xsZGAWxIs2m0
cJgelViqWLHb7JrMFtuIC5AgDtHZTL3MXU+jk7kAaj5QXWB29qhPL3ZQm7l2U4eFNtw8NHaAcMYk
1frIbZHlcSE2AKNv1PJuX9bUiLpe8QB8UM1L9zJAIBK6A1/jZ9G+gx4a75C/UtKanJWethKNBi4B
vL6YCw5RC+EyMohwURyUUygBHiDcFyozyjZ+1fpjUN8oAFdWKZvbp7y+twIXmCWrKJUIvz4DQftq
eOTxhOUnZF+D3E7pmKYmJSRMxNgXTbIpdDEUDTgCmYkSq/9KK7WpNERHuUO5T6GnAru57R5bBWg0
UaPUwqsNPxXn6nDy8U89ASurpolNR7g6IEXwS4WHkyeb4g5r4gvFHHoEF08/8stwNML5mdbYGf90
obtixTkQ45qkiPKdXbhRoT1pIRaLCD2XJMVF7oVRGAsajNL+wfW4XKVjX4DuKK5DHGaBSEd7zodD
06Tlqr5CeH/SbpCf+JIM2hI8RkDbIU2ZqvpDVmC/VccnVV/XPtq9mr1C1JcygWgq082FXYdIgaU7
dM/2J4YEOWugjYgjr3/oblUPfsGXjNsbK75qO6qk7u+ABuH7csdVQIRO4bHPUL/ciRnSOZJfrMdk
YafxDnWif3C9iriFh28HiGD2jioEDyJv+jyZZzXxz6BLLt8FX71trDVx+ORQTmsl+Wg9O9naoABa
/mfYUgLHOr2mWiSwm8DF6c+bM/+U62pTWbB+nCJJ+JtNoEbN/P2b7haB5byUVedMI/EaX9ZcrlTc
Terv7xRpslzJEn2A1BtvVSy7uzAxSsVUDiTzzylcINBVlBKw01yi7EDUE65ZMMBKZ90K2KFPKmXm
oFv8MerTsl9aMVkhdx6hCwj5RLetwzOO6YTZBmDFz6HDlrIsAynzJHOK7YR618hO8Zy1uHPP+GJU
coFETOKh4+cviDTmIxO9u5DpujXkoRcGX/ddozYX8FnppYmDElTgLwedKnWFFU00wmp3rWAVJh9P
+Us4xnpYaig4tKZgqFh8i65BbF5mHEfuZKmUp2f26LU1ziTGRI/SkNXNkJ3He9zapXuyrTvO6N9E
Uaa4h07NDy/um/oD1dW+5xsmiciNgiSmfrdJGjiW9n/+fgMYbJYrxRYA9fKHptyfk7PUOcDpYG5g
m6+raArz+1/XBPHAVTgI8BwLbjqbgka95+lw9WEMeAa86uMIVUrlCcExGRZ2tsLfZQTM2ThmeUGX
URtZ2w3gUlOm9973GsORhJN+s1iLDkXVgMFP7oydifScz7h1x6aRMWTF255g47hU2cAjdJtV8Pad
lzjERKdyUYzEm+25HmVJ2ZKyep+gYlRDR3IRsa4CsLA+jndUv85nURlc23vdDxXgkdrH8xms8V1y
tiQjznU4QH9zmmpSxJZD4G5xms/vr3gZ1ZVaMgptiODiIxlHsfEQ1coxXqnDShgZg1fOgIHAOLMM
6VnWjDse7QDNUF28z+lyXVBLCpZvD4fw/GZ6XLdEog6aLLVo3BX8p+dOBVlmV5cJJfRWEvIP6kuu
CCZW+W5MWmtgaUcVow/5HktSJLTPG9dan/UjksZzBOqTxCPSKJc+uMPWun6+08U9APCJjXku0qv1
bborHwAvWm9XDe5sM1KEGpb9TtXyhfwwRUF6Blvw1wLBN+lSqFCUXKpjutNNx7+GGEHylxgg4pLN
+dY2JKqoCbo5GI5V75Cb4PrG5r9NPXSkQnAOnk3Z/PVdBJAQpXYUOeN/QrsAauwm4QMiSdbY8u4b
vUHOY4+mtlGF/gT3cj9ZFGm5hfZFcnIL3/O7DqQxMCA5lS1EYL1qGJvPbWUpbAYOSpOHX7/as2EF
x7hLTS4vPZrCH7j30tIvniEM3au4a9r3shjsO6r0fyLbLZElqUsycPOtH4HqOHk3jQLcQpGuYLgR
VB4yehHzH1lsvdeS/Swcw8jrV2dYRnA3iKNh5EMJ5j0YgKCiZrBLgdi1reF5bladUOdLiRp5GbSn
mRFZjhb6PxadC/F4pxAtbTAI2nETWiLb/Does+6uGkxKb+Ty3jlzb6lQ5iX/c/OzUIpIpArgFYHc
MeDFXVAnVYEBask+akG0nG2KylceJ8VxsQ+UEorPI1E4MEOsTgR8xA0zZk5KajaUgHNyVwEe00iy
K2kpRL9Fk0QXFQzBAsKvcHoDmt4Mti6+KSiDr8wQppieCmfPRjiNZii7HZdXuOLlfU4VmkPW7hlt
Kx8wzVZ1tBbGZGCHRnEq66i0gpMyaPCEWifaDnCAloFIVICg10DXq20wtfWjnu19Xn0hZGLgU2rs
atIPxFFhkx0/Y3hGcLoV8M6LLrwyEKS3cYonmeW5598QHPf6vPy0eNTe0lcc9cQsx7+VIiji8wIv
9e9a+rtDeh9Xoh2DwZbv4GutI5+Dr6zf7fG9WUzJfuCuMcZG/vrXejmwTrwWmJ68RbpgyptTYz1O
NkIXsjHgHYVMFf5UyPtw53LHxfr9/i1W6hwN3sh+r2ESPPiSFySGXUNBOpFuMjkmSfUoAked0aYJ
E2fLN/KCWS5llSBSwkIDRm6aHQulr4Wa+cSGEcQsz0/JS9jeJJA6R9ZcDwlwCxKZecOR5DZthO4D
JIUljx1jxHRj0fgLyyVYZrIhPah/pAzMyZ59koYxHrZX9Qx9eDaZLW0czrcDUGZO+qgCGvakFPmz
xtTsuLqh50mXIe24DEOJqVe6JEeB3cGt7BGGaHKTWO1kOqc4KLw/o8DnY3VrVw1cxKXVtAjUkvPA
F4QSEr21VEn0Em6f/4CuCcCSouHFTNB6fs8VEBshq+Cohn3zqfqi8ngEIubv916XqaqGIr4y0g8x
sD3toMk2GN4g56d7pfttfgh/5826U3sfUbQuuloMO1Pr4X9C/8H0pa8AhgHrlerHsWhvP8bHgGot
h/5Ar9Zj0uJfQCnG8TCMWo/b5PBMXSMqmaE5JekrTM13C+z6zUdaYQWL9uRdw23Y7eSmd4hOmmKl
cSIIY/k76luPRVPY5wz/kRPRCi8pZ/kL/igRT/ecVvyYCV2WM5SkYujNlrQeeiyKdVgBGahq8+BZ
lt4iNPPhz4pVbhXwHW5ROt1+7zsc2Rufp1KPRYaEf+3DDFHM0ya4iVHQa9gDL9Ikyy8nYYSpoUUT
0hiDg53gFWsfKMhA9hS7FwyH3jAZQDUohx9nJRGltlA4c7hA8bg5o4FmDaL7t2j8ndcqhsPqhmEs
PJLluWx9m8S21kSDqGIWM+H8vF0ZwxhFe09sjKzkNPJ7zuetTxZqdPGuEvOoW7bKY3QuRF3IGXqN
Sht+yCzFYv7KYftLXZzYt240Ljy0pTEONjrquCXr97iwWP4xF9BEdWUqXu8E/R0XpKCtUVtaElSr
ATZ80PZQyBYvUIXyvEPy8WtRhpnJewqkWmVukpf4rOI+yYY4Y5FVSStoPX2UjETCbXDa9yE0d6to
njp1jlGeIBCW0CzffwuvGO4FEcJRHHBQyLtktT5kjCQVrowOt57D4VKP2vbjwSgJGW6hhhVvt3pO
g+o8pkHRnXtjZiU+bEXM+9b93pFnNj54jYo7K9jALewZsOWrHkzdKq134HpnwjL0OcE6GIWdDNSp
fmN3bDoCNCIh4RYE0pfInlOz/u3YyPDP0aiSWgExb35Hllvyk3q9e5OMOZ/YCeWXDDPTXOZ5BkUb
XBXCBBD2iFJReovXw6wF0IcmmsAjXGvR7hK1AQWfMgwEOFw+Sfh/FXxmrLlTRPhJreZP+JJvxW4P
11ZNFX8oNpC5D4YJayLX5lWcp2+cfFNGPPLTqPDib0IHiErh60rh0ugBCr0JgYpne/+i3qL8xe4g
RAGLIoeNfaxfdxscUi7I2tYZPV9/eh4YEXc/BqiXfVVNm4CLI/Qyq5lkA28+mS7B+4MXGAVqjxLK
glgVXoYQxpuVzLOsyrVHmDFQhBDwLdE8j2sf4zlQ8hPZtf53JN3/HEMQxUaIyTSyjIpH7JliiiMV
T0FCQHyXGA+zmoKdd/mfbHiL72loD80FfBAHhWb42Pzh5xpQtXvr92ZeP20cUsGfu1r4cpUQzuu9
HPm0Iq7evytYFkfZ5TdsVySYSGWBgFKMpoJHZapoSf0PZwDfY4CLdeT+/gUCzpLEIpiUqcsozifg
DhEdnoXvAfhcaFffVpeERy2y8j0VzB4YMn1wF/aarC2JQhJU5RKS4SPAbL0Pxl8QnaE3Eg5MQuBT
CVJrzXplifeliDwKAyOMwrkRr8pgaGdDpsqs9RJT5qj3zjfFOpUSq3LrWWyeZbPxveTV+5RGa3E1
bG8WPbr8WPXmVf7iv+KFNhXrv0+2YtciCQoMmIspI3knNzhzAcxjGWaIzT1BXK3i/u61GGvvnN3c
rjWry7zicYfqmjbbQ07BF+aKM8k9JXAGjJsfSBpKWBZdH2YKzgLiQ3+fySbwqfcd+FORtEFyPTb2
Bo8RQ8TF5+3g2+5FeysW/BzEybha4M7Hcvv/IssYC2+1s0NtjVXU9STtuJ9S4zqSKK4mojEC6sBS
mNHb0G8O9VFM6deUrVCKefrv6N0QAXKaXFLonMrFkUezJ5Om2I4mPdDDFhKhjNUkuoboDbAeH8WB
49aXcR+tq3Znbg2Il8JwZ2bu+7LdnWhdc+SzNOQJZOPgAMSY+D1ZcCVqu9Xi2Mma9Uuok/DzLMa4
gnMcydmblm0KKQsj0YXLLqxESz4Ekm9Ba/biQ1tiM1efK+R/bqQ0619jENEUx6VZDCgxdjQ+j5O9
K0ybK7Z9QfNcaSptMjAkqVinzl1mmABTjWY5KKWKXhovZqqeOy9Qik5WCVz5pNQb5Btdxy54aoC/
gRQX0Y0f1liLs49TNtpSZhzPYs/iM26eBeRoEGGUPT6hTpc51yfkKmVdFKDx394IoqHxgip2BINr
zmQ5pJ73QI1AjABeaZci0bSc+4goaruJcEU+SlQNrgKrrYzOOl7wYMykWEYCIBMn0LHE5clmb2jy
+yYZTF7U7iJDvV5F43UahH6OCqfPRv3XHlO4BXEdCrN2bXSDr4rw+wiEbrTQa0FnMZDGzrHutozd
R5PYkG10PR5UiGSQhs19PsJk8OHvHuOC087Z7o23Rl2t8cpC4cl/TZ4wxwsWKc6b+RKRm/4LGklS
gW2vNF9AoOZvJ8hqmDBQv9sumwMMuqCWM0ks2qqYPTw1nURPuiafULf1F6cx3irvDK9UzkFPovJh
qLuWoeaaK1DcVRML9iCoOmJe0/3HaMrWmT5dpgKoSXOR6DnlxG+yaaBi9dmaJFZW0Fmhbf/vsN5P
FZ0JF3+5a9U89VzBlyy3JI10drL7O5e01kwPh/KhdXHr6wc+BFgMzmPCSyFeTaGQHEMHbj2luLFb
0jTQID4tff9q1/KymXKYMJb9QAx0Ys43d9QZpFtb/KaJEMM7w96W5UdAjtZa/fEYmxd1D/hQ1+ex
DSLmkbrND+N98apKvKwwP5IdnRgNCo2D3b5yMCp6h0x5GpEYTYtGuEKOn3+7cwDhSum8NW+3owCm
tgrb8cA56S7c8+usLohAp9aVT/cNE6Fsp0HdXlT9wfyzlEEp+lb9A1LZzfWDYEKrxdxBdxQExKRr
jwX4iw3LxOr4ZWBlz01+u0jVz64Tl1/2edpYjhqsGx6tBmxbx31mxARftj73WfjH/CBoaO+cG+88
7t3i0fbp7zT7UkbChW2pSyWhjTMT+UlB1wR/qb4CXv1OnFoBGEspFzIrobfAWRJbQiiR1a4kSB2e
+zm2Q5fnovIdaSGIFx7lWYAx78hnf1U7QumkAm83fakWmt90zuVUq49faVPHYHQRKL/zkzZSLfnt
YEH3eDT0GWAJsgTQ/bc9kiBaRhevK10J2dWEbDFODfbF0MLHF9vB3F6FYXYy4WTvqMPXIobVwAjl
HqD6/20IIVbPxZcbIXkbSeMsS8Yc1dIxYsGTjTyGqU7vw4wgkf3kGAB993k9ZWF1BoonbVcJjl9B
Wm3bmi9zm9MXQYM+shHBOAtaLzSKNfUdRpzZtIUfVdDKTcOjC/nzJwMyvqob0/O+wug5OR4o+Dm3
LhwUYUDMLGR7Emw4hwmHsspyQ7zGKeCd5nGbCXJT/Ctor57Mj7Iu6gNYdMdUFzlSnf94u9iWlvi3
RVq30+oSqRjK/QkIvkooNmW1urjsaJoSrnAKJ0prOxCEh0PD24ZGLlYLNe68RcwWvhARLSXhRvmA
zVx7zZU4zebAJ1Ot0edNYFHrqTzZV97ZgAHmkNt0s2bY8PDDc/+6QpbD6TAIPhT9CWZwcGBZWYri
kSO/DS4xA70BOPPL8Z9q2RuoZR/DoMKL5CqzSgwg3XM4j8F3ygAAs+dxA/21D9m3Z79QiUH8q6bx
c6Eg/GN6bfiO0vf3T12hYbwiR4icGElV+dFIXqgCW/WbVsRVpexTYMdX6pm0abUAUaN7YPCEGObo
Tu9Px68ghEgE0kAmL0pPCff2z98lHTrbbvzDlD9LkSeJCOkHgaoWTCyb2le56H2NM5cYEJl1tTYs
jIrmbOaLgjJ853je/D42fi7oSjAkVKAYrKsjk2uhNL6GM5SZs/s9mNKm10AvL1uzRtyr6OzKnY3N
x5XJ7/FUdZuXGxLKVNvVcSlpsMswRI4wM+WHSyx0NSQsQUEGO8z1U+c97oH4CEvWd/8QQDPuPGN3
K1hRM02fqfQ21PmH77icZC28570qTlNwOrV9yvtWoGBIjAzDbUxr/N68Tb9vJUFyvxmMTBFt/Lh+
dj5TxFshtlaCLfWuylO+R3RsOgItqO+ePAixWwGyzf8e2zRsNcV2sfxlj8lS3ejXHSScj0XMxi2i
GYmkS2dbfrauSQZQyX0mOf4w9Jc1y5ouV0Vjb+8HSuX/cnTrrkC1tA+GVXck7fCs2WD7EqttBAbY
4D+AKRXW5qBmqgERz+1/RyawLD2sJG5Irds+cI2kQ/UEaneVCn1c8w2M0jPra50j8SzF2KnuT196
bPkgSTyDFNLzvtuBLlJQ9MP/kEhbFASVKC5v0BKO9ERqgHVunl2NqPK/WxDOcBjmWzFuC24pYj7O
3myfmIHJLqO0m6V3NS4bLWiQAWODwBgDLBJHmPKnsg/ew03H+XWEX2fEBYp404e8HojZ+k84cjqP
CZacbDJEe5ii+tdYjggIcGHi+QOVTBDffbsjZnACSEciyuZJmZTOslY8uD/ArnL637SD+QaQrehX
llyAhdedY27w9gysHn+SXwjfolfS9QPk7QeeSeiBq6Zzt7q25mRctYCmhLY4hRUwCvjU6oYKlwGc
0hY8bGuCwGMR9VxGFj6usE7m56e7ahjQZ1CqN2z2vAaNlulxrvZ+JAjTe8LK95Uky1Hr426tpJ19
rYUEeWDm1D1DnnBVJUicwstmAGvcZAqCQ00fBiGlMrgdXfZ/OjRGphOJ1wTVmNneFTBEhjlltJ8K
lV/XpgsbENMKzHP1gM7/9s3IhrcT67rQhBENW7ZWEf9vCHR3SqRnmR3mbrf6iChn2w1cbIKmNEoY
k+tuE/OeqUlIETIDNbGJsAhpRn4iaSfVHz07xnezjEGbyzk+H/zD2Su+BzGP/kV3krl5BAXWY4mc
DYK51Ic3smFktXeV/bASWH7tRRH7KhG0PtabUl3VtdakdDygr7gynWiUG+6bupGvbjaS7XpvytKY
bojmcNYV0Wuies4dTbDydfBvyzBDtez+eqv9bmzzZq+EQBAE07q9ykQetNtLi/SVXnxTm2QkPXIt
DkSf819KssAZeF5nfcby0b40A9ljWHNUbtja4r2m5TFSBJtzZR64uekqvOgKbDZnYT2Q9VYvuKW+
aBP8ucCPVlhmCgIwApdqsfHz3/eOH6J1uEMiTRabtBkjblsv+xs612S0NC7TYJxK5pkIfKd5nn+l
8lJWikh1gT9ZnzlwhxRxIGy73IpY1zBMMIoX/98CwlVGYkUZ232SGE8stsx1g8ujyg+j/a2j+JxI
8KLwWTpRhbXgs/FKMWcAu1Yo2YOohbK7fuDb5mxZ6h9YRWjY/eyGddjGVDMXMpDOYzJXP0wdKn9N
MqA2BJc6hTJptV1rT46Cd2uQGJSp8j+OHfEDafJDwULXBYnHwvgDkU62m20UinFUOijn4hX3WdxC
HyN8W8nzt0gJcOR6xZS2OTfGL4ZHD3ja4X2ogFoJC9lD5q2pnK8k4bpD2vr1RXX8ujb2X56vbDdz
lD/PajmVW3PkCzH8qjLwfpgTWjQ1QI8GWC0FAhHdo2YMwh9oN7POYoQI8Ed7PW9T60Ehf9xNOp6n
0CEVCOYxpToERaX9LiQyrCZGszRfdjvVuxjMEg8X3Pciy+dOJYaOgHjj5JE5hhwX2ljA3xHhY7w6
A0IZGpl6FFdqrLh3PKV8ZRNwYbv6Al+yq+tUY7dykWScjZ0S0/pewxf8mK2/n5iTYgJGsnXXotsn
kJwrxPjdi3/2xgaPrHV3zGIzJDxUjPEmcxdtJ7K/zq9VX02ipJ0kaS+CLJktbVCyarGaFerwur5f
/Nykb454tvtK7RKQRUyFePu4tq/6Z0O/DfsjPeoGc84PbnNQgJ0Fna6zdWK215JnhdEg2r5BRD0I
Uf0ESsLEwFF/yJSNFA4g5k87Tn22sJ6bLWoEOrfPV4xm03t2smRqc8Y36nJk9sCOenxYVvnZuE5d
GfUXpMoCCE8lvm7tZ3qRwVJUcoOuk3KMdFhvBEMsz23ihJ7PjBiqTXND67m9sh1BGBu1Vm59rDSB
C8K2/9hLFR5WdqrMqeMIXEYGRnled3TZXknZzqlqPqSzePZS6JGqq9GYhuXuMbjI03T1ycfhktgx
K8Vyv+pa1bzCs8l0XM7G7z70ddXzBhWhvCAP3YmKvpTPBJZrMkJZFp8IwqdNeosmxRVPO4N2u/JO
iK//aESD4QjoVgzmIYJOTD3Dg0bNE8wppfkSrEBAxpSkF34RHx/oEdQ2RZMBAQH3UoVzOPOptWmT
oK7Mx6oCDruiUUdZK7PQ1QDFAPTOJRCiHEpgiSg+tx4WQpN/gXpm56PpODcwapUaG/rUKxRwS5CV
yj8mrvZCjBe/+WwiO5VvyzRNnrIvcnfhK6ZAm6bFVJZ0+YyqnEr3Cc0uzjPbYO6X+w0uOZSE0AGB
8JeyfwPiUM/h+CLy2CaJz/YD4mNnksu5mn3/FD15DSun5BwCV5qK7L8FFOM1+mgWbUrAgSF2A1Yj
Z6926Bql8NdsiLMYnaNbcdHRd5Fs5SPoGjxZRT/c4VK4iKi4gv1ViNWFQ5kcgY55x0usUsxI/RLL
URHez4cZBmtUv3ep2OlPHA/41T9dJhJIsJLN2O5aEP+47ooEzSyxmHSGkz2FO7a0HdoypdpYmoSE
jxpA/stssJKrP5cwFHVbw9bSPXOk1nJsJnsJBZoD60A0e4e6DgNk6+qx7eqaQE1H0L6XUUfPyfVP
im6QOONqFe8+MxBxsodwJ7K50WnQRaDWcEe/N13UKLVN/KtJxlWBKfRw7jEbkO9x4+hup0Nf9Z6k
S5ssoJi+hChrDCicQxj7T+foxtdbUrArPLK5/6CkQE4a+1Sli0FA0O8tuq/vYDpk0jsq9BDj7tZY
FtmCaFr0VLxV7GODJmrv6VItQefdQv256tYyHxXJlW7nVB5xxj/jG8TT3Bb7+IsJk3w5iHKPiuxF
gFLruWU6SDdoelW3g+tass+D86ABD91BmTie0UkFwsVF1K3xoGyDKLAr8ZnW3VEcm6Z9s9Sb76Hm
4G98dIM5O6SU4qRDMTQ9K/XZQmAr/ETD/cA3tD8MYByEgTtd5glXVJ0SB9vwF15oc2P5HzHBuMok
Kg/qX0n0hn06KBjUaWia4dJ9Bg7kCOCuT36eP8fsmALSM+JBuxyuxhAVZ6gZ5KseQlqjPys9DmCw
eVr6MuiQDjR6cp5fJ8+4I9sbNtyLXsS6YY9uVwziubhY+0YMNF7rCJd/bmPv8zSW3PlN49B+PoXR
Pdid/86ByGK9kYxpc7KuH1mJEl7JXRdoobHgTtaQiYPaBhN7c0WNfpYuchIY4mys1sqGQIjqmB6k
Rti4Y9acDHTObKSI6kwH0k9uB+lmAhBmwLg1gVdiFMLlLO03VaP0Sstn/2l01+D+m3SSS+6z6J6k
vuxY2ugMaDZIu9t4j+xTCQGAEFlGOkkr6ZZvw+EdpaYksvXrRrtVRZvhAyT9lnx7widVlGs9Ikrr
7GMpO+wZUAMRzplmsOMwciAg2mbbHPbUGrSYFsRVPKy1/Yke8PvrauHsH2DCVRkYUntZz59pOunt
qLn8nl+QJDY54J7WLo9UbJvSsSVC3cdga66SHDC+mNYvugLKlEULDVPL4AcncL4pk5JqPcupbTVq
7jUzm3xaHslit27Ph/VJ3lrspmL5Ct5dZ54lSWco7L5h6HMo2QA+Bfes0fRgLIiIbWW8ywjBFiZU
+YSSfBR0lta8JsJ2/Zqzglr1u+wM++acMlhAArDTuyo4135IyFaXvgqyEx5RrXT+CKqdoXjJAnxf
Sc94LpjmiodSdS6hjYUD8mAT6AU20+iKv7hcR6mnUc3WAR1SxIlB2eFvApx3QDEESVamVy8UlGev
rw68/xs3cTMfvK6DMkDpFLC+X1X/rdsEjm9BfISQEFaVHgVoyf8O0TsemfF72A3LRsml9mq9/qLR
LYjkmVpVT/Jn0iPYEBCaanptuJjOyu4gb4WKfEqkGXLM2EeHlRzsgMgiNgWsJsgjfTn1lv1On+z8
E4H/WG8a5SSgyuULlc8B7qmBe0TS8TofNdLklwV6cDe7LNUBxUgYioAJ9XeuLhULnIcYzkWLera0
ZpanIcnP7Okv+RVSPJ3WEZ3KEJLru/OcYn5WbEBh+W4m084GQKh922MJOgWt4UtSi+PEt0rhrY6R
QVsUQgPdXXpFR2dACuEr7PFQURAOEVotRxOi8H2SyWuJRDjZis+ffq1VxYNHWsxy+AZYailfyihE
nFWYG8S6Dx7k4K9521Il5Fv0IBJlDv39KM60/sOG/O1sxEuZij8wrl2GTN0g9+uGXPm1Aa9thZqc
9HULbwIzd9YJEGTnj7MKvbvGHnBYmdCvitnvDfOdmKoCWRfXRYdO57UCcRRRlU3DK3bCDIHzaB7R
7PN25CzPy5vW/3zUgaTdwqumAsk9sFdBKpoYN2RFiisQGmhp2fROaY/0nXrl95VbZN3ivX4+nXex
9j0jNO+g1qieR3F/rncukVi9hDZWTqKk4jkDxTf+lJG6rKm5XPwgJUs58fhP1AcjQdOG1DmbiBgR
0vFoNc2T+4BdXMgEnUep3AhXbLAegkPGjKp5i04GPcJRl4Ruqdbc7XMaUJ/HLC49bw8RgCWovBN3
IgG3l4JdhKSSjNwOuzYbreh/scsGVKedIGbwYAzSyNgi5p30pF0z7xRgRF+LKxy7Dr7YI6TEdB7X
0JH8x6MyedEKlO0RYErhsXOkSEt306HQhGBpYQfSRMC1xxYQ90yTnD4NxbPN/o0u77ecSNVQX450
RajkewJTxevk0MwK/G/m0r9DgOkqRVwSqhoyU3k+oMJLhBVIB4aQph0NrBa96Jo4w68w9R/0GKdC
WPbWJOZMrDoM2gHod/QqimK14LtB+UAKCO6clSYdTHCSBwFifEYfgeT00K9GGlq/FO4+n5d9sGAq
Doo4PbJ8Co1GYPWtkyOdIDZbznwueTqSQT+ozxLqvdblsR3M+JAIiFbpucMHTHy//QV/mtM+OKlA
FfotNo6cuMqJPXDMIrHcPBz/jBtnsJyWrp3UQKeVbS8Buxx4ZjgZASqsuSIZnHL/2Ay5s5F841oX
t1u45okPFkWG5oOWKYNHFyHpJ9HvUAennnVIVRKER1guPMwybupymbCFUhQBd0qP/8HLS1MsNp8/
gmMNX2REEXvOJIq05eV6S7SmsTFwnSaCc8wEWz6Dvty/IOGLoIEphxyJs/BgFbSe3VC+xp/jOmR9
YyTUp5BoIG32u40RJ46isPn9Zri1DTiRwOLDum85M58wyVIVwzUcOfpg1TznCPcxIvMyDSFkAMRM
RDG7osmmoMRYmyuqUjSPpVr9pGn1nw3oyVrDsQhGKg65BUXc5eC8oJC7G63E+ffqLP5IojOawbL9
IInXmBSn4lPgcsHXaqiIqqPVrcjDyhbtyGdZjzUvaKHlf+XyCvN+1M/9xKNBEj8T9H3IkoUwL1u5
4eGr4NfbdJXMhUyAoN68mS/mCNZZcPZRdP0eCMB85Uq8+FnOHwLhOW9MpGrMAA3ES0PynTQo1nzB
lZ0FhRcnVZYS18HrAf7m9zCLXLBE9rkh50FFrtP1uz/S6r8uUrrwIQ7bIZElsbDRk3veag37NxmC
LwHpvUciNOYf1qHrTNvBtgWP8oqyfVm8/R6bsakChs63IuiiIErGBtlTWIzl4LjAqDx2OqvWxlWp
H0znyUuWmlgO7rHex1+TycwnK6J9KGqHDMG8Xm+v/sDFwGqQYHgW3CmxWwHoLoZD6TYu8Sk0U0Db
bJVjHlrFfTnUGbjedMJtlztyCwoTrA0cEtD/hZjTbhgID+RlJ2KCw7+cJstFgnn/M51leQ5yPHu+
KDAZgAB9M8OuzOxwec2BEyZ+7TpQrC+Rfz3SS/pfX92/DPLRswr+II/Pt2TH0aBDrM2oCxtNaEbp
UgRpgoldjOXccETvmW1ceWv8/friK+e56jeh9g0mkLjOtrWuZBVfgbV73TwvdhFiL1cEgeYrBBBj
5oVogVP9D94gehqqHLot+NKHJJrKwLYIasduTl76SwVFyItzeeyl8y+e3xx1qsBKMLQY4Wfb8xJ2
MfRpHFwHt6IPCbyWLIXewQQ6e3+5Yx/Q+yobmYo/wv3y98oMKZZtxng9ZfvCVotxtZ+MPCww+eXW
bAW84S7BCbbnYjAh4/GbkOvnWtXJ3WkDOlnkl5AIP+KiWzlMyIteB5qn2eF5I9XBVV1jZSKo3QBQ
MqyI1XU6sord7XkKReaQKdflRprigRy28ZYgTvrsg4aNQDq9LdQWj6zgBHzxFNPe0deAN7uLgevl
PTsVxmjaUrCrGe4G/TJRBXOVRmxYUs3g9WeavGbe+HwdyP6LnftCflWT2Vk5OscpcEtcVi4xG+Ci
WhtWDya3XjfJ9t02vrV5cMMaBJCZQNci9smr4V+GKrrUwUatFjNIB4NuzzIJFKWQ23kPvLrJcLCL
Q3JbqiPn0II5cdbi3A51R786rijO8GCKUqFaBlm8BhT2ede6LmFgyCycT6fZ52rmSI6W16cb2EmP
yqMPsC8kV9YxxW1unTqGWc9gT88V/NYtuBxYVc9h03/yFR8Q9kL7ucJWiqAw2tOcyoukazc17T8z
yhC5xynAadKATlCTbdKRx1RhWbzCPZBaxHKbaZjfc4cu9xkjN/RaO1MGAusi8+a3yMlCTu1OUiDC
BFRxUyPE0/hEij/t45ec3/mkUSLlxmB2Ah2W7j/Vr2JAlV2ME6fz18Iu0PHj/5kOL1F18bk4Mnnb
HWC8gENPWxxA6zNxHYW5d47wo++wD8eaUiVr5p8DTvwPqar219WEbVRJ5i7sOobhVRz297PdPSKz
aWrYpxtZDmJR1XejEguoftcb78hdOL+GQDObbT3Tp/xakYKQLUd2p8WENOgHaD8DGU8cC+QMkUhK
+fCerfrbq+CIaL9yxl1UsNtakj0d1/etBOJIK0RBxD41xRXeT+SKqjSgLYB0G6/v/cYyyFB3XYal
YYdnbB1mRBPJOrgl68sLukY99Uq5BR0jEGvtX72wuge8DDNuvu7VDfcVoMqYycjIZxWuUOGhmbob
78v31gwLE9Iiws+uU1287+Dk0f3a3E+/C7hdhukktPbeWr396HJGm8n7QXMtUKgO+gMGRsn381mm
Jcrj/SVqiFSRC9XEIRejUv9PuSuoQnLZt0F5RefUBp1Nk6hJ3gpBXPFaJVS3pdXqNal5E9yX7THT
Pq73zaB6j5ElJ66VD9KFXAF6xWs0c7fE/BpYRrYDpEh+s33RPcSTmlPo2ZM+5zRPbsNlVomeybc7
Cv+7u7g9rrNOmqd5TvU/iAx5RIu1BmZH11uw79lvyrF9QnllZ2hETNrU0AXMUgWQPLFVg/p8b/Wu
9chVjekywcdWuLqiDonGUopf9huQ+Q2NTHXjLQKu2wXmCH//rK/d3krPYoqg/3JvOaYmjIfqyrDc
iVmksnUkaTn6uDSqbBuVx1glFa2fakBuTqrxLmvBkaM/XL3/MmY2VrdNm2xjK9zn1bVpqCvXW8ln
r44muQmS2WlWhG4JMAisTQZSdzMoiGhQmjp2H2GQFQydRQ3WrQswP6mHSVk5wSQVGRRN/GfTWWww
gWJUwF8Urcd81Z2X4bpxzap4aBeW4UBX669Wf4kijcAbZJVyO/INhK/ZscBwmnq8E/bsC21csCT6
a29zREiC8/GDSMVg41EYiM2/DDU7hOEfXVrVRz4wstPfcuc9azyTDNf07daT2HwWSY6fn2Ztc4HO
R7NvQCEfvGMXEewbVudA00UwiZywTfaKYQE+V8NZkmrxKpU0xSpD30a26g2akOG/Ce4mGEcusiC1
j2k99NR5P2aq+XsDpibH83U6K0119H6GYdFTMEUMTXnooogTjBFuHYWicERUvOlM/41HZ5yueUaR
WpfqclhbrOLbw9aKq2mP4h8P4cjOphg3ZMxAm/yXX3SZKstwKg/bWlQeE2Dp92mBE1VsaDtPRrsr
LsC0h+ZhuNDa29qBiBWFf03LxkXUqMswdKKOeVcvDRG8JOP5A2QATHDB93JUA+iF7F10TNNI60jy
y9NhvwNRcsVMDuPYax2IhrYX33e204W1bc14Mc1yAuNG7DaJ5KCzBoyS5028WaosKCnEZMzbbGiD
VIWgfs8B4B0Vn9doxXW00fzOZgfST0vlnrUIQ0P4XVm75gwJz8bBW2R5VBs5Dt/OKAP28URWEbvE
n+okmRS/Wij537sGDUMItPGTV5xGFS0U8v3HdBffijOhUYmcOd6O1P2qzp70T5tKPm5nJArJN66Z
Ocd/sGhDlFyF07Rb88tB/dtH5s5MKiedktWG7n/86nvXJT1BL2kbHUW06Qs+8kCWsw/UvG379Vau
/4g62tayR7IR6rFHA6CYIGnQJIFCIqj4OqKZnMP4OTLTv4qs30w+N+8pyfP27OqYJ0ILpc/DaGj6
s0Mft61bKg3saUNyoGypEnpYQiJmm22XSNdfOO+/amfVqsboEtvL0kOzevJoexMhd2W2PVBdFtzF
dwFgDx0Nejzc27vfl/LUC/yaDqplvoE6xFQWAfTxXO52A0tqlpKNStc1ih4x+LckRjOy4Mj8CF5o
/Ej0zss0XBKeqpZUEf5apWbMZB2646osKdtIjactT+XcVPfYCnqjgoKV7K925mooqCs5nC2luT43
8Bn32uxVLygCzPommCi1JyQ5KFn6gPWEZoTLK4yvw3+Bw6odJohTNuweDOhb1WHODn/pIeBxqoUn
MOlpJVfQHvjms6USQPzc4IXFk/LmHTQnkbWA+mOFj18cPuqE8dVqm54fEP4iY5SGnhTViLuc1N1/
lHPCA6qwUxmJv1ppcX8PDZxhxHmuFOHO4B8p+GC9PZcCmrq4l8g68NsfzeLgpC6ochJX1FgWB6vP
EBc8Pvev1pUyvx/+SykPDVpbHzAZAYevQYFW5ou3OaNmWRtx3I66T/bzPFmWWfV1HNiCmDy6MIc2
e4cj5TXZ6AQgwJocT5z8tL1Q7BAkOave/kQd3riYfn6avyD8TlPe+z7v6Hc/w3mzs9GbySEDcu0i
rRKNAQwvn7m1qDlolRa3lsIYKs5uDLiEZXD7peh70D4SI7IL83GTRfMqho5snEOKnhX9nPMr4Xdy
rYfFKWGhkPETZubOMQMpR9fN0Jxv9rPy3jVG35zdlFnzHFcP/I4I3boNIgigl5gfYj5TL2Clvd3S
Dkw72bZKkApXvck27RKeT22yQFAOYZDCfe41px22Xhp8/P4RNRqt1GwQjJxft2d9E0KtHT39Izhj
hAgEOzH87sQbWpkIoUrKV94G+fYBhq5eGEpLO/hXsbR1r6yYXki/MdJojtwCinvblgbmKPJY3YAq
JJLWC6pK1N1sjn/LuVZw0b2xCRT/mzyYeN+ec10TzKqLISesmZlqYcQ29VfsmTZGd/F2tQT9/Ndm
GcMhpMYE5aoV3AsEzKdCBCqu8Z/5073wg1JLtz2lqsB1quLGWatbtNc3DEbx8TB24jKzil4r2L3v
FX1BJg56VLDHKGXFdGbhPCc4PV6WA9BCgXkLO5cYgRt4t6FKjs22u/M0RxP3SPp2NcO7jJ6NcQT7
ud9dCSpNJHQXId5gitlBP4rN9J40uid7CzFGRvxfuBf1aV7NBFloE8k4o6KwiL2rLh0fsrbRJoBg
w+LML0swiVYPTug1PssXdLJsy/MNNfUm/P7MkCa31MfQ3zIvQqLE1Z+GGLLIDuQOcki56pPVmrfG
iXvTT/lRSM0Bnb5vXb/Pck2XlL6eCqniyL0m/tQAW2Cg00g6nmmf/kq32GxwF1+ke2WabiJJl/Fg
1+4havIny4ZSMUjrS/o/TxYAqA35hcWnqXw1e25dkMg7MsHz3eMqmmMwns5TL5pgMk5Kv1IITkLX
VVRJ7a8+Ipmy62gOEpwxy94Kx0MFXbTt0j78kM7WLou7Evn5po7lPCIjOZrMun4exgKBwPk5wtm4
kjLTwzHbOM5we9/qPVax7nDjqR0TXTW0rrhjcvNLkKQdBM8N+a2gXDFVxhGvq5NrI9CzHGPPo9oz
2n7bS5kvKBRqjdi5zjFqNgSFbk+ZbFnCH9BeGQdXGa254Cd77N2XGhc31e/htSADNjHwRg41T1L+
/AWCtR0mH/0gfge1VMIdj62M7UTmgValGirpIrVVTDOwfTnxRjOT3Qk3H+IPtqKdkBbbB7+JLs8J
CTOe++3KmHGH+AYaIYFoD1/jzA9c/Uk+1vWWxPFJeOxuyTEJUuCKohlTbh6d9WwAzbFTEHhnCiho
iX39kA/N+a1+TTPsQcgZFCWiXwzWakURwsX0kk6WVfYPJVqaxl4PTe7gBg7wmhMmswd/XFJAAgYS
okHeiiwPXAboCfPKqtkP027XHTcKxLd2tTnfjYRArJNta1S1HKBMjCKEEATnn2qCnCdbpSpOgSXN
5zKfWaicj/J6opFsRfDy14hMdHmze6K57fIvp+TvTPLABf+hxk8vCL3GX0vd/i4Ng25Ej5q6yUhP
xbxqKohRjwVp78QgtBg0TW4sqoy2g8gFIJonOyCYWsLnuKktqk9spXVWpUocLm8IXJLproTnplCf
FmsLQD1N3W0t5P0wqEOeyUGWfZZEVteXTk5wLXVBdQhRVkNH0Uj5j/xwTblMp/PoCynb++WYAvFM
XM9sc/4w3DzjAiL0G2aBrVRyVu8knuCvaOmTMP2PyO2lBi6aOqCKT2zKl1a33xO9yNYu7w6daMD2
zAOE+Jflisp8BtrzyoqaJQqCvNYLTa/ZdhQ9wLii7OKhsCfzkqyqLxBGhgCyozohHhV5eU5qs0IO
OZLhLC4e2Xef1uqJDqvkYt0yX1PFOjy3lbNYDMIOR8lZ1gin565Ej8j/xZunU37j0jl32JkyaWyS
Qe3dNM+gZSiRgPwLSBCO/aSpA/AJb3kVAn7wIGODGv2ab9Bj3P4baGmvbq1LCLkbGR9LUAdDVS0Z
TtDVHgfbWAdxkUBpBvhg62erb4ydvZUYCrxzmzrMqnTIBYNod28XC/KXPGoFckAdoKNcBU9d9rm6
fqz2s/Ytg5gTaTl1sbY2UHPLMj6mzCzrk6Zjwxaz3uyFKfAmnhhBDe8GdLmYbAwtTmgjAuw2yxIU
R2MrVa7joLpQ+/ON5zgcjpukBA7wK1OC7dgpq6b1JL+hbqkmoVCvgPMRNchE716K3IJ1KD4jiVXJ
uXQu7L25VqXBIijYFPZvogyPKbWAGh0OOP9HLix6nvyGZyOJJlanow/fharDGijQecsu+rTN1VmV
kC5S7Ead6F1P0SETqh4ReqYz/T7NwP4RQ4IX0onv68V4AlqGBS39zF68p6eV8k4MaF1J2dCmQ++e
1Jpv6XR8aCMVJAU1d95PA0I1ID5Jp0D5iOwpTSs2FbHzQcEvvRw1qB0ndgFljzrEVnxwA0r8pWsW
8JvPjIKxnDF996wpypF2E4uSRkJEoKPMoimeHgukIdK4gKa9gwXVgaO/Qv9FIwxLOspBzx8rzE3N
9P2cFp3x6ly8MaD8eA6U0L8eiJZVahRIZfNfV6eQmzrtB0SVQUNegmNVBJ5gal1j7SlhtUhdTL7R
DSkd9kDxX0Xyv1uTmx8xszYY46XxKdJBLL8LaG0ATa+9rPYURWqOICWFRD2xmb36lPWjl+estoT2
VoaQhdoI+5Rqz6+t6lN8HHQzoWR6uvjEbNQGrvbFG1Ovpqp0XP99qMm99m9OYA46ENO2ntQj2ynZ
bB2O38eQOZ0ONMaqZfeSPTg8vVWK2ObWRKY5yDiz9GCz0Xf5W7YBxIdAz80lHnz9iwZzguzNZybz
EDZhhkoYQtySU2ulDkAfXWCiRcqSFFiYyRLpqDjhhCMwXz3w8KZqFvLPAfv9xySHBfZkpBR6jCIi
0TkuzEtf0h1XkXdC01g9ZyHaVhL8tnpKEHWLn3r51OiTs8s4gFgZ1GwrmgKswWEMWKx6v44rOeRl
uWI5APYseZDwRChdRVhaYxVnjsUjxqNQxkCJqfg08LJhR5wfeeE6HG+MyCGZc/CRYOSzDkouk2pG
sK0GF5l7MG/4CYuJ6HcZ4ji31tzGmJdasRPfdEqk+3Pfr+RVs6jurhQRlrsyQ2/+1OUIyolCCoVG
QOIkK+t2hPRMwhV2lnEUjQBVaDlMex0nENY/KV9D9RCkwKPn0SN5ffA5dzZExPEnRBxNWEmsLjKF
BaCtfQJ1Q9UQM++5mc0yfcGDfvaKr3SbpvNGr8ieRrB6j9Fd290K2N8o2Iv/h/tRchcZp/wUnLA+
Z/SVIfvgR3zaWKbCtJV77aplHW8oTqm4Qt46dblxv5mYyj4XnFEsDXMteepvVXr+kF4Xz7iSyObU
Qnsts+QnXy9zJ+XvnvKUgK77Ohmx+5aMN1/GAjqti6dtm41LSgK1aBRihjoPxOE/PaeIBawm6MKW
mo+oxsYav94wJy2vNhBYMEx7pEwUCK8HONNIn59j7wn2yqySyKaHT4gqX0gJnOug8yCRT+JJBZcd
6YRFmTdWQZS2XxXegny+N5alPDMX7STtyqD0wwTwWqnsZ5z5jxK3x+0xRTkCCweTkxZaTmABQVtH
jx1VyU7/eHg3zQobfqbQR9Yo25Zn0JdWviu+PsRcZyUmcVztsqxld69cTk8tgtz+jPYy9NM5bKe1
YFnYQg5SQcd8eqFaGubp8xTF4vT7Aamwf8s56ZCvtmmWsEc+yVVnVZ0r1a4kPwkWn3KHIuoUQZ9l
hwe667i1HvfXCM9iFDgBB9jQilWrR5Lq0Ol/kFvIzIznCYutICIMJsOgjMmlanwMqUBPGdwrvt/7
O1dAQvWs2IGHA8wPbOuUdMRKAyky9nvfpHDH2wzsrD1k8R3kR35NZXR54sWllgOC5wh5rJqyQUOo
hLuf5OiF/E4pDrnSoQMUi34CmmxB14UblGjXTjd++X3NabHxQJ1DxtqMOCiZW8Bu8C+xHm696O+L
ETZSyTjNMGkeq19hHJK3PYWIYFqr68F6jQJLJFGa54OtumFWxijBUfjx+sYKi5DaObZI3hT10j3P
XWoPrEUFFK0Yv07ZmDIZkmjQMHBlY6fuPOL8Gn0O3jlw8y33mwR2Ur1pzj724YanBqHI2iYKY42n
39mqWneJFji1XnVDdZ01txyYZW8EajOfy4Gr1+RLVKrPayP2m3yqYLj3XtakD1l9wJ39b+ynwmZ5
8j9x1OPyiu6weIg4J8bizfVBtp7S+SVBiM9zLnZFjjyxk5Dt80pmkqutUJmyeaaa4mrPzh28E9bp
/WNeNo0BGC2lo5diFltj/ku/NT1QTJM6yr3gsykMkxtgQ1OkIUMva9Y34cbx+iYvCtPGn5rvtFR6
/dkk/07MRJ6y9NivkyJxHy6YtgskibcPoSZXcfyKknQb999nfUGR3iMgK6N84asy0OknpAyVB0RZ
fNyOw7oJoYk6XCd3Lksg8h4XbqX6iEMcjIIAlf4iP8uaKKtOHEo82I7YExcuNfw/NaR3G1NlK7xQ
18MmFeaGLRzJKpyb6RA/sjNDTNTrW0Qbyc1jfgjSu/nsI0lRVd4TbqBZEJNBWG0DkBpD4AomnnWh
asx83BNshy+qZduA2dw1xr4weRSBXbOR43sh6FHmPtmsSlNlKlqNlmVlQhHUZC9O4902Q2442CNC
K2otFyyaM5pTk/3e8aR2CG9knFOYSt333DW4rpkZZeoyUWDM7PKazbRCxjZquwv96gNDssug6Lg2
uZAOcQGOqowMNNhTZrktT2dBgWx+rO4RpRUxaVIku6poPk8CAI7bvFJ8GULt9TC3SYjakki8Kc3F
tYX3wzLlsgOiP4lv/7G2qT0MY9tQcomAYnCj09LKMAu2dP/ZGiK3Gc8jRP7VvT/SrOLJM2ovecPW
1IRHLZ79ALLtj7/BoqhG6gOJach9EfL057eVynctLe4y01AUeDHxKrNkFQiNEDPmSg1r0hIn2vc8
uRxEWkug6cTnnrUCMdC6U84CYcqHjtxigxL1Ed5Bgnai6NkVFDoArwD7L362MtsokbCrvj/rmW00
HJkSsTkHD2iFgcdzviERnYh6iqohIWFco6TlQS7NeQtSs7JaVIHe7sstmQlMgo4trB0qYqXB5zeR
6hR1InB4QXU3mrWeW6utQ8Ty+uweqIt1l20hXCKduVZ2iXox6T3xu4vgAhsJb5xkHTVsJiVbgFSn
oKGUDrmsdo1NILzxQXHwRLPWqGHx+EQLu+sEUTKbdpSG2LRsUSbRYdFG/wtv87+HS6Rt7DxYh7ab
KojNNBh4cGCtzJlmc5ickQVqXrTuDd9JtT1UA18GM6zMWM+pg9o/XZj2wkIdcZXUPwBnpx0Ycg01
8FefeuF11WP5KDtjT+45GgjX5ieg2gf15y6Kb2YOIU55Q6G4wt42UEtr+OJqOoy8SwZhodDibdSD
B2qYy12L4VKCpz/Yf7qbtw6My+5PmvaTCSaCbJcP/AY3A3uzCBAosLCoHVahSVQBSU7K/KDNfU1l
h39haJCeu3SvxdxAs9SGS3XEqRduFW6gTHB19esTMlaUDtps05wlssvBiySCdSxUCyjC5AtCsNHK
Eik/+bFvbckrhdqOZgUES/jE93Ejxke6AVITNQseoNfsDRtT45ExhRHGfJCxaE8VTlqNHIId3TuM
rbub5SbQWALdg2qImDuXHNg3a1huWubfyLH3ungqKYtZCeNQF1Glvj0hYmg9mwkPu8j2jE17uNnh
FZX119rBLf+IeYtLBhXE234dUD2DT77iCColQcuX8VPvvmECukeFwul7s9oRcwB8vSrDhdZVBzK+
IpNsxegqu75joWAc26ypnjFzIlHAue7Scjb8PK7xpCcWBcPVDMMNRv2cWjtK7thtD9FDLsTBPe3T
/x/xcSe1YTPv2MuRa81ATDnmIU+46psFCiHjt1iEByASx9vAjR5ZEzPhN5ZF79apkpu4yjMFDoaN
M6XZEnm5vqKUz88ubNCYkXIYGXSCeU+LSm3DKJLZNENONBwXvCnewjFxNrvI4hDvUA1ovl79Xrgy
WTO08ESopsVQcfk4BLP2gajtHNbXHcvr9trk4/2x+5RwHWdnJ6w4yYKZmoePRDDv+3ErOPgfM0r/
G3o9J//b5RECLFCtOLuQKLc1atS7649qhaNLQh+PKBfArTDg1ito5M8oMJF1h1BcYtw6+tenrdtS
IkY7rWUD6K5hGPCGkEXInx9y4TH1Y1ZFuSkFkPSA1S6RPLAkcypBxNHjSqTv2ALTWce3ajeDF1Kj
aDQnWMVCcqVBnhbm1s5cOm7TRMKlqZALM2We7gS4HzWpnaCyRtloUmn5OWCHsdvYjFwPXkfDe1AJ
pB3UQfJtXNEfIbnpY8aECRcZhqOasYTapkVcC8yIRI9ULXAGDnLgGasjXTJxEvR8wEaEwTiXQ/Bd
PU7ixQLFKkQq4H0HxX5TGRunyOUYOpFmlu57dhmLWFp++koFXB5YZoTR+/3uG/ONTYR4vNp9jgGr
WoAz6/P1c63kHDHucWXd9/LPJlSQzSWlezvHn56BlMElexChsv9k7zxSYREJ/3WROzonfogu9OHw
JrT2YISnjEoj9r5EweNhduHv1MD2PyekPmC2fi4Ed0glOpojfq7ZhY1CNzWxXpXI3wnOknI6lgJn
FjpSoSUappR6E0p6Zs+3B0Y9rgKq5zWiPFqJJxT9vGmWo5oa+hablzYMScLEKIGXXLhWBvtpIf9O
mDqIf+ZECaXDAVrZLbWI4HrWRlJoV2q1Cnn9liykYoQXlPJ/MwtWC6O4OKe1rjFHgmdgXz26jocA
en5G5IyurtkZduHPOz7K0hle121HyLjn1r8bAJiiZlnGNXhtDfE48ZjOUaWZ9+cPk2BZ14ngnJyQ
2oAcT2HwGNG97f4MAW0nm2oJpMMy8Jj2wB8kNz9xXQ99vfB4CeTvJ4xlcaGv5w2dZq82xHjxytON
JpTCIZmst57DKZXqDlmNNftImS86IKQwPvX2XvsS2Ely+PF5cm6gw9t4agr7Tdx5TLSDlISiyJ22
x03l4q1cXFFMltGeBUzEYCZkf7PFDOk7UZRzm1j9+DhaNf3DVCwRzlkdwTeIQyfyYU/csHQY9Lcy
bINVLqmnpRqvWUGYUPXseNfeKGJVNjm4NS4qhzaGitcIYG5ZDEx4METhJM56/39KequwR0yIl4r6
qxGYi9XbGIzB6bMa2SYz6ZYaUKdNf9VmgASvRF5MP9/C5UTzAzHSbJmblKI6NeSmAf+l7XC6YLqX
4eyV3TaE94UIPK0iuQQztOTVD2zeL9z3gJIV4AomnMo+cnLr++tfbSyI+7SwPwZ4x0wy5Dmw/iBV
f4rDfie159J9A4DG0R0DEhl0b/tKsJI7LSpzjGMqDOmua86YZXTS2qQvHyQ0UhwBn5WUIqG1rtu0
NzSu0ashgobh+iNSM+VzpoC77GF3ynctFAzQTXPgw/2oHk0HAHez9TvQ7IYWuRgS0GLP+4LVvcEz
dT3Ucg2Frl05jz+s4ysmAT31Kze7Rn/i92smJQ8Lu9ENFO0Ma4kn8UsQnLkam4HMfEh0SAd05KON
F011T+dvjP7WoKHOb7W2gBWd3VM0PtwFbs8kN57f5xPApelZY6nv8WGhLRmsuKK5XXM+JhrupQ2f
dlwRWvuVSpsYr+DIckOkETW5tSf3q8BFmhoRYjJwELwkx49OhnEjqnrUO1CQGvZSHyj6WwdGaNUC
RJsnrmZbI6FrQMNQtzSHP5noYMtuaqgZEcAabQy/BIEBgL3rc3jLqfr3FSv5zAx4K8EMGzQY7Gr7
bVjensSWWV784pc1ZQ6JZuoQhZnB29gjY8beRSinN3kkXTc4u7yrIdKrx2yxTfA9VEkDSqxVF5dd
+du5zfWhvvBv4N+hWeMa1tNVsJGvzzf7AQwhqj81Pr/E4MYxJX//KFd5kmM3VbpI+VPw1xcz88cZ
gL5Z+w5owfmYHtf3tpOoWq0ub1pjyTxjSgSJwPhdImvo3PTinIshfWxayvOVPJ7IJ6T/Z1KT2Rr3
u/DyGkNQ1SIg5v5rrq4/Ktd1oCeqpG3tM2aXNWTOaISdqBmmk/BTEC/TiM+qqV4Qg9BMztPXzfiw
Kzl6FdUFGSVwXA8lRJJ9cjAwcGRCwJGt6E9UJUidkLtplvigVXPni7Aws2Ea9uRec/kFskRnzLMa
z0CKsozRfaUesGMIDAn35jkAqzYtmeKkE33+i09MQrlmtHdu9z4SzsTuD4DC1FikK86P0p7NvqZa
OZoq1abwHBPnzRyuaB2jg09GAEMvmOq724RQuWWGfV4v+L1+bYnvQwOzIvpcV7z35GTPpmZkB2Gb
ecFKOKu/uBlrLjzv6Jlasmj/m+kESqNIdJLmP6sk3rgjc/sdSmC0jAX9POZQ0WvdGX5tlafrq/Nk
dPzi5zwQCAwOjscB88mUdu/ml/SIV9pPRv6LpwHX0Fi9BdWwsUAEQuHM44bA59secGrjkt+CzD3d
MCzDYMbjwnhYQ8IN28dhX3/cqjyxwUIl3u5/60MkH5F8VkEt28i+s31OGmq9tE+ulm10FnB2huow
O9c3rAt7rHHUjw0fQMkfYXSceK0JODaRY7ENabi+Ord00Ohxn324C5RHDApQYqQ2svSCea8xN2WH
IFs3lmphHehcDuZY5+pWEXKWwNzbBzQEogyNYKli/luTaj07CeDmOSmk+A2ATKb9Zjb/WY3gRj6h
7xUxPeY1JqdP6BcyVc31uGmx4Ft8SkvOnqpllCRzlU8NQ6Qzzco6ye7ob69P94MoY3uMZvzNUL3R
exS/0ACnIhS83Fi1OH+6jh7iBOk9gJHGXZ5HjOqWlrSOUAg5IojPaGQaBL2Oaois/QN8JeIexHDn
mOB/zoC29QO7lkgRPKL6BL3Hg0rrVAGQl41nRS6AhcQYfE1z5faTHCwb+yXRKaYCkTpcm8j10Gzv
9jvepSEuW5tsnOd2kyGPXTWNciB3fEfaWfrUjwlS7q1pWNvB6dxmWQLUJpK0HnUe53EFyj0+aAen
frdgt5zOnO6urG+9IYxMmEqrcOikqtw48hHHrWnn9XvRoqwzGA1RbjFr7xA/rWVabHDdYJ/Ehxka
GkN6s3v3sQzD2sWvZS1c8PW6Mt2ZGqsGChw8gBol84ugeQ+DCfUF+cwgo11hvJICHI0/90M7fmVL
nC91svHq4u0qqHqyRZq2XcbAHS+Tq6GWwjI4ouCru2LZtI4EpvEmNUT2p4/Bgi9KHGXfgPhZlf17
S4/6O45IJs2V0XW1qfv0sGVOrPsZ1oGIcPrt4ZFa1LS2VdIrPp229cruPeIlDiiCQSjd/RqJR7R9
7MHCByhQ5r8IgTR14JTTzS6cPO3q5N4z78/0jLMWwx9AU7wspFGzv7XDsyAnE89HPNOsXIvx2CIT
As/8aSWdlEkj5iD82PlZL1HA7Nsy/AfT7yeX9RXRyxtrtCh1UFjiva63f8QZlj74CwtCYtu4y7l1
jcDOGPjAiJStB/GFR+jnC19tGU206KF+m/6Jkc7L5N2llrJpUtmm5esiLYwZ9FIuzmdu5v48S/Yp
eHKP77hj8OGjU8AC15PpnqpUVzU6/B3WSozrZYU1+vX2iYPbYyl3yzuCArYI/G9lWL+YIkmn8mwR
Dy+Kpx2RjUzTYihhdNAt909fInzXltmvIUJS/diUIHZKcorWu9uM4D7H2HcNlVyuyFRjxKbjwnMf
gq1uLUmBKuhJLcJuqt7bDL5scw32MQ1jbcOklHZ108ojhVrhQzV0clY3ermYl4x2YePuzHiRhyWO
C6AfVqZjNShE6SE7/GOU+2tOjXSENO9SMI7fusyB6yamPPy7NbxkHqViCic03VjtY9iDGToS6KUQ
VIXVUJijNHHIPN7fJ5143+/izCu2+cexrzKCJFAtd5RJ1ybODouAtYulkrUDVed7t/Keh0v85MKz
/M8dxLIg0Aj50gVA1glGvd1NmXTaI69s4jd4/0i7jn2HZJn7ERdnQGypiDsVGBWCAZI2iOuwTBfo
HDm1LJNaivPF1HltvxBLpclpKI/I6ZU+zG0Ixy03eqFh55Qb1V7sh8Fp81nly1kEyWa9f4F8EXj4
puNnnAfTSwl43ZxPmC8JtlL9AgKb5mRNQp9MvfcAkfxgfFzs8+LcSsVLsHIAeNO0D/rWFkdjhiIK
1Gqj+DeXyPEDGwzuHeVN2giWXX8NjCdn0P5HWgOckNT/w3j1FYMxys+BKY7sHVwjOWc+XV9za53d
oMQGJV3xMGJkjiC9pwmoKOKqnHCHb2zDwSbOzQDZpe6wHKrr5tM2p+ol7zlUFAyopqlDAzK6SDiQ
iAuDhA2RK3zGp0MvSW8Pqx90kYYO3vIRjVAMUxw8ODBrAUEmh/g2KsoY+CJ8JKFLd7nTx/3GcIe3
Clx+QgQ3UqtjX/Xq49sDaKi2BT6n+HEGfL9b86M/IWS+3VbKu6IzFaBlaoNMpSMkDITY1o+c+gci
bGufPWzYQHstRAluU/lSoVsOt/Or+BhLF5I3fcw+ctp+jM0j68VEveudnGgSRLix5m0zA+PUV7L3
HJXlt5MOXm2RgJK8AiNrgamrVQFf3yzWKOQhavloEjyo6ESXe7wwUbReKmhs+JRZ86ep0sYx7zMI
VWHlBssQf0NY/G5a/TCZiUcEq9LrsI78XwaaujS3G6eKM0wJzk6ZBZ6d9uV81fu0bDYctL/X4Gwf
oJGljJ5Ryfge0pktNDlTKdvKunIIDjrnKjzYJB7gG4k/lgft5ci4NCBYb+qK9lDeVVuxyyYSRZ6U
ltFDioeGplsxKzhLkOC70p2m/iDfXcA47nygWtS3Q/AOh8or0J7wttvvjRBZK+AHmXFJBlMQjGX9
cCc6MMUMKjxaHfoZGj8Vo1oWOvKqIK8SpjAVuopkjDIfRriCLIm582EqsNnE5Wx52sIiCwKcDHTO
LJspIbGfPVLB8BGm4kU1wBFQXqNv+s0a713UVIHT398UYvptiMbtveYmTV95YA5JhC94eLMwGsUs
37SA8a+ubGTNshTZ4yHmJXliejoMfZG2Id1SQn/cWrgbrqCYrhdHLm4htEalWnW0tKLQ4I+Cxrnm
02A9prrPiXckLSY5/I6BjS9O0gX8fJrPHC3ma3DJBEEiLoZGvF10RuWIrkpOmHye5xJCLYd+v6f9
UcNeakOp/UYyxmcAf4aS5oAnnivzlKdIlxQCpw7KvLvOkA25V7rt6rpbayP7iPR56V3ln0O5earw
a+wtfiD0cgpuwUAaTVfzGofWZNoSFrvNwhG+KMyo8N2Tvbwj/ldkOkRBmGeSU/HwBi8EXPjPBfqO
0gdVZ7PZaUFagS/xNNcg2SJHIRPAXLPwgUqHG1H70p48NxmVNnuadDnPDIDr1bceNGrFEG5KWfuf
NBaQTSqk2tMq8lb+NybY5wMeGYIa8wQ6ckdiDllaqjSJBdP8AW37hQkJG5cRO+WPXmiQFel8/bKq
8v5gc3HmDp3cjqIm9R12Ljv9dC+Zvx1nEUu7vPNCLYLLXYljeOtx1CUHiMTfOPKA4Qe4GzdDoHc5
u86WQi1D3jsoxDiE5bItqitkSrAHe7yFgrQ7I55+TNfs7kj6Amsf2xM6MTK4FYw9HhAGQapF1vMO
yhe8qXcF9lD21OCkkaW/184asR6qYFM18BdJaJSwYXrAe7n6T2tmnocrFKbZtvdeuNzSncGo48ee
zGB+VKm9b9sJKTykoVjVpZrYlpAkX8dF6BLQJLmgRWkTk0lestrH1sKHcQQ3u5CND7+NIeoBj3Ss
DgsWJ5JRI3IFEm4am2osamsfQqREyEafRfnvMAW/CQAMlSZMxxwKef4cinNIvAvV5YGZ7S4oXIUB
KLw6jdDJ0m3obnPjXbJ9ug1CVioIRXGPKU60SliILRYCEk08AVXId69xJ3vwtFzNYSD6NpHvajrJ
We6oIR8O8QeSk1P9UFvBwt775ObK4dbQQrmPAAKBDX3jdY2ExzerEosyRdDf3IjY4eyjg8rbosgq
ETSZksoUxmkW0DvDdMb2GpnpjyInE+ZQrLLCYLvwRgTPN5W3M6hFbSsZgKPpGWo8erp7Ww0PROw/
y8Kswy7V8SbJJ8gtN6tg5xXG4cW+fnjIp59Myo78jRyzQ5v5gn9876/Bjj43c1gZErdUzTrbTHVh
CGP53dgWyvQrtbaQrYzXHRoDQvTIPO5zbcKHyeqV0X7PBxG1ja/zkzDrjcSN4Wm7va2ZmqqshvBq
I1Ogxz3POefxqy/D/+4JdjPLxk809bZD/PyBWW2ihYL9OHBtIQHiBtwLQWlfZwsQIRdl7eqxP29W
u0Psz2Sz0XT2bw2EQ0ugmmoc4Gdb9XuyUws0a6wA9phKa7eQaChiBe0yRCBbg9LcFQ6bz+AVoHoL
zJRlAnmR+CRtcNaW6vkQR49Zhem4KXOgC546RlJ5sWKVWDa6062pMJckANd45okiM70FXb32MRtl
0fIXtmHLaicslEDbfzFB0JXl3hGN9OrUjZ19KxioFvnvVMecXFIJScdZHio+JtIRf3oSHHdORSi7
6uhpqsfhgr+Va7Ss0w+NJncRX+zQJtIzGX7yAmo6jnRN4pma32SvzOAsaqVDZGAhdbdTo29VWsgH
o6OUfXo60S/0TyDPus/p3YD95EzlBQP/pLuEB9etw7uSjIqcRXtNkGfQfl6XZewNy9jutEo0BZ6t
+qaC4WHFl9TqnUrlPNAEkyDpzaVdzm44WHrs18LTOfUVXuC5m+lVkRlX4EkgiVMoOmPV7z5cIqFE
uZteoa5riaSPUnFCgYNv0FFUE5SoNFSJIyl+KzEgTAg10+A5aglCIu48Ol60IzEc2VzazNesb/7Q
MzX2rjt1E20+mnnEFm49XA+pR8Zz4mH3yTp3L2FlsjcaRwZjNLErEuXdXOK1//+pOaM6rKnfOOu1
9WGwJ8vmrVNWBXKM+sEwE81H/A5fnHQZcGDGrZgN5giYddfR57Haisk4bXnZh+aKkyJoiFPXTnjs
km2O+cpwnkob1X2kyB/IJPuS7ZxX+Q3vndfBnQ5PAR8gTRq9YMqW4+NlujIVyWjpsYztWY+xbEYJ
/I+N2cAl39/BGl4QU5mAm22kBfXk7BID/mBToQmQuaL8Dz8qbSmfGG1G6fo4R4pw+WdjWGpiX4h5
Kmtyj2gGA3XCw7IUTsN7BHi+JshxkuKgbdQCgDJQ6GQP4EbTojbF+9o70VJjnLxrrHMDSZT7bdTf
o/5pFILT/yeviyXUvBb+3FuP3VrIi3+JBfvG35tWCK9cZ4H0YQstiycOip92RHZjdQQCS2gkzQ4f
djEVl5dThtdz03ogulICHkkvH9eXNxBWc9lkziXDxQxWem3Q7+WnMbiro67goJVlfVITpFU/5Fr+
RUYtqKiGoJIw0eBpohMz0tN5yVxVP08TZKp4FDnvghf20+9zliCM7GB5/A27zNXXYprL1xSgXgCD
F8stS+O5M1UIhvnrKVr52wLk9aOR/vjNJzLp8ZUdlJNt/4uLw83rB1XYmAvBPHCegVgZZ3HbU86j
6gurD3snXF7IA97tvWT/KegNq6+YTw23n0ludTL1N7ZCN9K9VmRMKuNOjEcBSWDnWkbajB94cC1d
3hHOqIgeSDj0OvMnzP0U9EIjzOs0tf10aQhU+2Wd6D8jmw57lQOL4cdasJ6FvNOWY0Rq/DLJPnI9
tNxaVgvMmMRZQWsSglFTVTtIOGxCeHPftdSzmvW1yRVMRDtEvkLPTtRr0lUnH04UjfoLI9jRo3UV
3qzC0XYyvFZ72xIx7goodePdoAwnqEICUwIgaiX6EcsEtnsxq3VNEFyw9/zV3m6oNX2wrypqzF7J
4ajvvGg9jUE5EKbnkCm4UZk8gd8DZ/vTBTxjfuXBviRpt7BIWhWOd66Ne4v+csYHr+49s+jAfwpE
atcpyMs7fWKc3LYnVrUY267Z/9BQu4Zpjv8CWA40OMtFgOeddz5saHaQm/9yHv688Sq+zR1Vp0Ll
6dnqWx5a8hs29kzlqbMXQT9ahYTuOABrGUYtC8Ev9KpT9l7dPcxbcIraidaQSTWXkunnQZTGyqyT
HKCGyzdiDGR4B3QwFRltKMHXnk2sgVmALaMSAkXIHvj/L5GmSaVZLk8vyDSXQuyiGd7kdwEYLdrb
KXERcqdrPRfT+OIjR8Me+j5ohnLdTh5c7FgLO+wJkGLxOdw6g57/1o47JIshk7tHzh0QMey5Yr4D
70RTDl3oPAQCKFkzdaOaYKjpSKnDyP41/10NaWKSTY5eJYUaYBW0z/FIZm7riwPy2Tn8Sbn9KrPm
mvjF3k5UBG68eOXfv4tEHeIcPMvHohPsdkWRMWihLuQwybhLBMM39hk/GaDmtgvCb73Thygb6KcV
zdtIsHFgrKLw7JjRCxyG2lV6MjYLyT0fh20ox/VPpizCiOA39jr87tHzd+3jt80nShNzSPtD6Q7c
eo3d1be/q6OUQyXil4oYs+YI4wTnYtIUgrjCJb63Y9E9ay7mQdqE5KIw3YNG6Juidk+M1ppmOq+h
6Rh2oJLkHNaJP+cVmpiMh/wT4ZyQWcVjaFGsHDg7CKbEnxf18AG4tUP8hK8Ei0mBUdFBsAh4307C
87qbNksp/eqJA5+KiPBJ1vqCbgfCUzDSMbOAkMCzQCTldL3fRzjlrDrRFjKdej+9MlOvPe1I3lYQ
YcD98boS43o5AwZHkQpq8Y5jyEQas6GIzd3IWoU2wgRtSWMKt3EZt/veJ5Jj8qReAZ93EwhYEjHt
G/RgFbtBSKxUbISv5f8wvIHpWRnr4dr0iSQSx36dtChBAIGjVk1miGkUsgpIX0Q+o+oUpGcB0oyO
Yw3BGhp9eI9FJhcUMxx++7rhzY0WNbxuDqsODWHgD+ZFf/C7uDbP+ztBzkqudCl4fD7TWrog2JQh
b4R1RVC5/NPdmyKe6FKJ7ffHu7SNbxcTC4rHnQQP6OEHp0tiLhRofk+SjGYx9K8FHgNDZhyJa+y7
h6rKP0bZuMf4PKehWTaRw023Ltp+29GJ12KstPgL9lCkaAQqRKtKaa/zI4l8/NeIcNNyOzLqbOVv
nALCezECr/fN73DmmyFj7+dMFIdeZ9dE2WT7uqE7va5VHoarJLOlNwaYorKBRfvaQls5mBLUTTi8
AdyEQ+ap028y/HZ+OUEXE3BFsMSaMvaLgdBmUJT90ZlTnubGpnnkrRoFdlT04XsnbMYQl/YbAjMR
Wq97SePXMKCQOfYEfHsKgmQU8z8kAgwHZ/pIMCkKn8XT5O37v7B6NJfVknMXg5VVvZgTBJ0wJAiL
+pp6YH30dmXB65BxlAGFATxmamUxkAgC977BXAjJ4DW0S6KRp0dIk4xq5MvzpxGuBw9fyyZqgY+E
f9Pu4ns9pp9pEIfbBjPwPkV6i3fj91K+Lx5/fj/FwaYG1UKJIgYRUahfMgGZvY97HULGrWjnY9SJ
pQE9tFYLU2bFOONk2w2x5haW3bvmbyPI2jtEMfQ4yF6t7Z713S3Y2kQLdE2zmJWCne5BtHbexoKW
u5BRUHJw2RkJ18D/h9j2nseoLM3h7pH2tQSuyAS5x0JzP7kvzjtKnUcPtNnncMxclaz4l+/zlo6d
SBmfCR119ZBn/ZnhCBcDGPCdy68K+3EIyUY+xOQDigNyFQyYc3B1XKk+P5uDMwUD8wZtZ2XE4K7W
02iUK6eWnKxma4h2DGTA6xDSvFOuNZ+XovmNk4P7lRv5nbty1LOipV12IYwPZtadbA9IkaMfY7V2
09B9GXcU3BNoWdbKx0i3ra8567pYVwtrF8j0u+9P3uhkTZ3Y5Ws0XcMJ/44KjpG9R37wse0ywYbK
Oh+dq3P46Sx7T9P9PeTdLJAv9zO5kSD33lbmcWhfz3sk1yovHk8ykieKt/GxC6QCj8+hv4xoFx7p
t+MzS6m+hMMbl4MC35a9qtoBaq9FPdCJOJoCehFyvczXnXintVc9XVl3rsjDA5t+LkpwT4+/dp6Z
ctPaTevnhyjbG9qnqJx05AjCrRLYLr4oDpYqIJEaHIHQxjXouzlDaBIexgnitJbDeAFVqCBdQo/m
Ty3+mclsXPfrRULoBezlpSCDwSDcmrdwOU8GLCFgfgilu4lTEWiYiOwAkul1/Ax5cuBX0hgYZupE
L5dsRlfj2DK3AhGCVyNwGxuOTVzU5MSPmhf+eQl2BhyeIFxz1yd+LRpwgO4vFTG89jg8ClrH4Tdt
GxDRZpFNJnlU871U2FVa4sMAI0Cce1wT5msaqbagcMXYj8U2Nyf/gYe4FRjw2L45vuVsdG2AZTsA
YqDie0tdLuFMkyvXI2sa5I5tNfvc7s7Keye5g2W8tyxrZ/eAZ9SiNZMkLsbDpE+aVdgczpD9UTrD
urHRa4S/DnORhHGRG98aDlaa03WgJJ5DfCIvyPdopB5WfpqXUxoUPTmVpQrj8MggoSOw6uTuDj1x
1f1JXDwEDu0hUd4SPJZtpWRpCOG+47nJQYko3qFvouuD4TAkV1L41FQJ5tcbAzo0UNqW95B7hdiY
cD+37evmb4vZMNGrl1ENiN+gv9EF36s+byULKwue5VQAZc2JnYm2K9uhwa1+OIsMNhq9vP+YtEAU
Ftplaxqmgxx7BeFhDVJFiLVuWpj8f6MRLGi3Q5cQOwMVUeQRYb/b6D2e0HI5zhkUG47A05uRwKWk
muiSQvztnMDy3KmF9O33XJr5+dUFnD3wx3JLIDfr+NSFM2Q8fCox9sxdMLWdpGcP7oyJgzFQFZyq
Vwf6DJSzEwQ5S8I/ORQg1N5vYqbSte43B0d+QTsep8NF8xFJTE8BDQjRYGF44t60bccd6jeHqKw0
DOEg7/cRCbEleB7v2ZED6S4SqPcNSwxAGd5E47K/MnuLkApm8b1B8yPsXl8ghN9s5od+a//A2SqJ
uivyG34XgCRXx+F0iPMiEZUPjYMVw0ZjUU6ZMpaPB4t90EfgXciK0SzbiKY47vYdrbM5FGl15VO5
JW64O48Ghaa2oQoh55OxnCMPwqyPNUyRo0IyYR5ePQff7a0zYUe2Bv73p3BaOwXaL4A6qYb/rZ5j
+oSujlIUjDJWsr5QB3WVfwZRMfzePcnyGF3eep2bgfiXbnDZJEXJWYx9LA9yyZb5VS28Vq7aFjWa
8MxsQrs5VcuVprwZjmNoL4Nm6i6eoFZ6Trzr6JTPFDgNWIpE0ZpbKsZF59L51eOHrlSj/4TMUcxL
pyYXFEtE9aCSZRbiJHVOdcWB1IZwPJ/os27fzNlv0GaC7O52um2aRut4KAX7IMDWblwan93GW12H
VC4j8R5qWPAt/JCkloXxnS1MHpHP1FIBl6+ItwyjhMn54M3/qeOqAvlBWyFnh45209uJzsHskmiK
vDBV3jpv3LuwW6YBysiaPVZQQJGtxjduHTEsNQBMBbYW6dNYF0F8DyI/TSc2JpAEX7ZkoBcwDbZB
w85f49AOKVswyrf2W+4mjx8B36sh4+0GgyUs1cy9thMxtZ9ro16fzc6UzZCIveq/RRlf6SR1JxQh
7gljfFiVfddTJJ8i3CxKDOC+moexYIOca6HHLBjkpBmB5aLbKofetbI474t3osLxX2FHYNY/A6tV
cN17zuo3It+u2MK8zGH3ZMjp7v//5zPEiUkJhkcWzY59WFQqQoYtOzI7RzRIOV+azDaIGq793Xgb
sbplz8dw14NZ2EByncQFS6kTVPEAuaDz0SgU3kDWvnHPFdvq/7QaMD+ouFDpZXG6yBYo85p6v2zD
fBQlttOSsvDKYCnrX/ZbDk8h+v8lbk1v6N4DpYo5vv7+tB0Heh4zwF9Cx9iLewgNC3PST3Tl+o8d
hZT0mE0ocMImvBApeAXXVrvDZSfPGKbDoycncEsEdAMYS83pkhmeW6lCN6TYPrfMLlRRkaN17SLi
slqxd+6QyzOKRXX2A8R3RsGsNnFr/srLzyNTA3CudW7nNtXtJBOhvM3G+WvBKTcXI2iwq5Wxv4fv
FRdvMslg73/GmX9KINRLzLg2AlIABQ39J4EXktd8uBQVfrBnO4ZzOqKBJEgB9n983vcdXVRbcrUA
4r9A/dAl1yvK+cEpAPy93Sa+QPplv4s9aqCxhSMaLu2a/GBd323bLAWJQdpkq7UbddYYlJjF6bNC
IsyvtEJiSceuMIrfUnz2GPnJKwdRPB+i+xP6VcIlQ5Guk07Ydvox1MhCHi7RJqT6JfYQDjyvW3vU
v3OR1uYWivh80hWiNZRKqQYqWHAgCppTF8SHdZHRknnclD11lihVlkKgfzL5QTewFU2mWiAFe1a8
fGwNVqUWI9MrJ9t3DILHyhXPUWC3lhgzL5cQUKa+OdQ/oyEqQAIEMR3ADpgwPKX2ELn7Ms+AMfLm
SlFAdGOFri+qVV5ylxrye0dpk+JpJU1NoqFjo60tLjedjoMtwul6a48W8zRx0XMTOD+kpHrlO0Hg
e9pFMVgIkQ2nJQnf5zb7utrj+PmNeg0g7+uzoA4C1ASAx/iJf++5SLzNCy/HMN69Ot2CZrC9nqlw
8lxysDKSbqLejkAUjoXQfPlm3irqCTmBx6SXhChUOmDwwicoXVSNEsK/y6BgD0OLNkDHG9arOHRh
tNW3+K+o3d5uZuD3J0W2VyGh7kYi6icj6eAoAkPfYKpM3q6pn6/pD0o3R5dXvkUggk+D4bZWaThn
qF7601Uxzq9J1z05DBHvK3Eq/SYqPoR06vZx5VFGqkoMPF5Fp+ZPiLUvoAL6F02PSJs73rxvfY35
5rK7mLMdDM40qCSmxrt9IM8eF/VcDR9+EaFM/xzkqcoOlG6fVd/RUMMBQ2W7jCOspwAEHtPv1WK6
4T+dfF4r0YuAJy06BkIUNm/kTo6075eAmg+sDHHzSskc8V1RF5JAmubyX9xlDpGm9AZP0ONdbI4S
xr+WamX3FOYUe7wJpoMZsrD+aliCLQCwhkAdLLtumEpUbE6UQ5U/Gs2nOFPtClvFTd1IzFJUzBLi
hjdbYJ7dcergTPjdHWtykXbr5Ms6QZ04TCXokT6HsbaGyIERJfGD426aXHNqSlnh2+7ddwl0+Dyt
WR6GODHw8qzaqQhYUXlrmfj3kGvUtC9aRm8zJt57lXk0WruYWSs3q2t/WQuv2IIVWM9+FaAszIeV
8IojN3uIQTlKvUqulBrgg2UwQEVYWWd0roVwn5cuYIyJFJcEjrO4tXbcfgUGglA6YMkjN0mFJQpA
b2TvfVahw6qOpxNkGmJtzWm+ZQelPeJraA9BQiFU6puksyA6w8Vt1bwXELdRTLzpo1QDIrG1iiip
cfIBFCFnSusZQ41TzISAc2VC5qIcxYymfNMUKgLX7RNK3xrWpxL7ob0KLWMp02lEbEPdcruNXpfy
87h3cIp3yNx29WNql8j0DGdNG8gVVHK+/cZ28QIEHfzTB//BfSl5Q3kiXMufzxBlHk/e6wsNAJv/
n9q7Ac/6aCvaFZ+uDi52IV4oJiiHdryX3LAgz3UMAf4eSGTF+wP8GKysrWSEpb3gZQSUpMS23d9K
r38rgsqYKpLUqtta0+z78KrqUW/a35RzF4EQwDfZfvHyyFQe+51MrQWNK7UWCCanWuofbMWqQ48S
BBjFTzeUyr+UCoUM1Bq75IqLuFZpiKSPPEEXXG5qGXGW/x3LRIoZHB6JfpJ4Wih/R295RyvZFcct
/akrjua1RYVicsPQd9GHn3j0M7Sa30eMgp8Mdmx0ui6HYE7UVRugYauq/yCdzRdumxB7SjOUQtIM
2TWgppGGLdyuH/+PB257baQdciIiQsZJvex/Gc7V30lw7PnVW0fP9oHYvOLG0INF33BpXIzcRWna
nWnYqicPIS8sOhuGtrFVfENf0p4PfSjbjOKDkvj6q/QL2+2BuKt2qxgtdq+7ITTnV0ttUuEVkjfd
JrZRWZhH19cZ5aWHbD3K96Fg3kS/praBQ2eIDNHqGHy0E27XE+mxBdNOY5u4VIYsR18QPBybmaKc
k0Ru0twQ0G/D/sFNY66cu2M2jyw10AKh6HnYZNYHn+dSTSTWO/k+ErxWAv628Ww4ZfspPf2Rei7+
gen3qEjVcLuEewhoRwndr4rdDC/tr/wpG944WZlStYHHEDyNFhm6bHyPmrHbCk1ZSVYxWdbaZRJN
jedykOphZukWCMRn/foqOFhGp2U/1Mx/1n0Cp4KxGKN/7xXy+0Q5QxXwyfdpgK0AXqQ5JgH4eSmF
VugxF2XQK5DqEynAyTJ+lFvAihUg8rNarPNmesyczz0/GlZyoPBGIGWSALDn7Uy485iFl/g8+ok+
ySCFWUI5+99Ti353uEVuafnvRAvRcgza0vkx8Tx6QAocqPPZOkfvCKu5wVIJ1rrvEQTjL5OuXm/q
Qu5xo1o6ZZKk5hyiLbjNBQ/Xov0/A6KQ/BSrsp0kMdU7ue20De5VNtfKO0wwY7+yo2SjxmcSd6z1
frSiake6p6X71Pl/sYqYmSvThTO0BD+RaJpN6FTWAWEJVG3GbrL/wlbl+TjHrr5ViMa6CG5YYq8k
dpEQSHFEtu807V7pfsW5rk4yvHhxoHjBWIgIcUXSkurMgXbGeiYWdNhvkJ6kGlcQbCD+x/VqiqLP
5FiP90olhBvxq6HQcfvJU+vG2qkKDg3Bp+83rYm/K8YoLyPlEYsS7wJjqEUNrEju6yyVr/Pa14w3
RsiAJvTn51VjGiRVX+WdsK648xm12TT0Rlt2RattFn8pY5dEekK0jRXzAvRajTo65jEFATfWHdLc
2l2SoLXFVckvkC9O6A+faGud3dfZWCEa5RiG5CTau/7gOR1r1ML7btZWoeN6cSytCjowP5zVyXwu
16Mx9q9+GCkLqlFXxkTKY4cGaSQ5ADCTEUmltKLw1RTcp9mHfMzb3F90/n/YpMpKGGlE9kZkbTXf
zfEJNX283as3e5pAk9kBCUK9WlEYyrXOhBqhDp5/0wyRqA9Drcks0W+yBBsDRc1DSnINzAA1rgvT
qFwJxPI+YvFGXsSZ7+jqgIOivXUMCvSthLE+LclqxHKxT8S9mHjq2B75XYoY32kl3NTX/HtNgu9s
VKKRT8XQhsqcvbYMrGCgUJJW99i3InYv7sKnYWzLrktpHwLAH3SFmSdsGtBUFl/sIuG+aVlCqkah
7EVvLs/Rql/4MZlAdJ+yZ3B1pVeWKPeim2FuMPNy0szyF4f1I3z9sW3L1122nifVL/fotCNSMivN
NATT2ow5wp5iPlntUT20/mImnVXZ53CYr04iuilvD6W6ca+Bt5bnT08ZEvMNibUK2I353iMCOlwW
2Qt1dRkoMaJmQbiAIG1JIjd0msmkBAug4rCpWxZeVlm2wfIfQxRs1ICCm9BAdiBSMJVrmpJMAiry
qxcP0MuS4cY2Q69i7DsKEr0ZNpBMWUOO7x31RgMVHLzIdmFY1b6fr40K7AaarLL415jVQS3cIG08
+UiJwj7sK+BFnQJnFqaeyJVHZkJC1F4qaqGf3g7hmaE6/Z/6oN+bF0rQy6WBjx3/w53c2JADROLR
9xpKavQL7ldLctRLbUmgS9nlO4WK5ge7cQM4opBFsnu0Cs2yGsl8xkpQgYdDU9qhE5NyL7WPlh55
NFkbd/kt4sqMkauMVfrTh9CjkVKsyGRyT+ttDBNal4w8K0AjFBEF6glFo6MwJq0Ffmeo/4a+bCR4
9RavqrKuIX1Ki4b3MhGdrdImCgJGf/V7sMzyH+xmPEtgcdOVX5Ede4ZlxYxVUmpns7O9ogYW2vHQ
9WLx/t0kmUl0EhkNt07Y7BxENJ5XRgKCTt0dVMHC14b0x8zRo1yuSLJxaNzeqiclHK60xY3SLLik
EsWvrDWKOJt4CSbgbo5L4OzWzzYVvrLQHRbfoWN2AUq7NzSLJJy14nsUd37YzfMfZw/V9WSyIlk9
6ee2AjwNh3vFcObuAmA2bmHt2mlyLcaAELM9fyyf9QEcQeeU8YZixFT+/JPRfwXJYxGJYu046t6J
IhV5bRDMWRcVhsgEDg7PB3LqvgZeElVILRW5+MtQbn6+VW+wBD4UCxnnx/ghabuWLloMIUZthLhV
1tOlT7nbOaXqFvUurIP67dZ5mbsKsduDrDukPY3djYy4P4SbEPXbzMR1EngfpzDqYNr5v/9xD6QP
m9uYc+ORYvf8/WEzVAHADZ6eUigYK5e1TSoG9i3gYd+Eekg8wXi9msFnrrBnA/uvTWDgTp261nxh
z8UeG3PsIXC1c435xWLtjiwjDE8lq58vAVMYaIb/V/AqpwqUXi2RWo809JAmJeHBlhQTF6u5ZEdp
NgJF3+gzDGPYHKsgAEYI8sfXkBSMvZasz6cF7Fx5KyKNg8T+6uS3w+HesH030YpzD7bcMTG2p7cL
iJ3irBx30s48mXtWGyI95qNmgf6fHwWTFk7xlE6P0zXF+sY1bznfWwKbuRwHJ8GosrXw9CAxUwVF
2Fbmzli/lVHDetlVLNVYyVXYDh9fHIk4JSO8mZEr2NfQHBruRCqenQ5RUZpfkuEdZdzg3VDpKffE
dMfFum3W168UXHoDYAVTd2N41J0jysiHOfvsDqHxct0T8hHBO/4glwuCx09f9Z0fm+zWJ1y/i2vZ
SpaLNUKZcd3d11iTfW2fw1WGMRJt1GwrXwBMz4DNlP5J0h7+BT/zPDoq4GUZxMKyftGNWRCNImvb
UbpEJtNztck9xOU1wPPl1fN3u00h/VdIlznr+5nLYknIFT8IEcOWfhFcdoWIRlMwF5wAt3lQiQzy
qY56rI48UwWuAy1gqKQlfQHWcVmZChDX26O5ILpuA5KC5wb49AO0qC4Rsy6tdm/NDHx9iD0BnW9X
ZY+BnXR9dMi4fM3kBJ9eZvDpon8L87SBbj4UP/+ZvWrFhLPmjTw1d/zqGCdSbdgb9wFmNtsvcDIC
A4NKoCsGku58jTv1f/BfihPBeomM9/22auSZXJi+uo4IsZr0v+PP4yCfYy9+uDM6QJn3xFtsETOm
wtajpOrhTzllC53PAe3VO9ttHB9NOVLaXs/NzmTvNk6FXq987r5wrxdJbYPjGCd/nYkd5knwC6CH
f7ooX3zsU8y4DA+hNnK8UPoeFsFhjy8OPct+wS3/wjXX8UDbWlgVp/xn7xNmHB5jw40uCzGgkzYQ
kStDCNj9DF9Ib4lK61r+J9LbUqlzlXCJbQNUAHZyyzfeyJMQM6EKWcLI2zkEhE3sidgFrCk1u59x
+cHN75tOOKgsfoFqX+sVDOYU3ibhBPR+N4GkC9meWTWi96Dj4dL5B5Vqy2hwcq0+q7dDkG0v1f3x
s2rZJ4otDZoBe81h9tkfTt4qwzs2uiD+6h2X/d5kTwAaJcTOyFX63USsqWOPXitWJOuj3YXkII/d
5qZx95rrqg8Z5nh4WX3KRvDV4wU9PW1HJxAcze3qHtlBdSyMJZj3YK1tVHh0WXbmp28tOCw7m6BW
IQEm9ik6OyNIvofE+TnW1EuSOvtICFNWwZZYCHVzSYmQesNbQyb6JTjJQtOTlu+riZgIzyg87bNQ
noF/Ro16Qp9nkzW/Z+xBNTOCBlonVSmLDQiJsdqS1uGP12nvvIJ9+hr1Fk9cDY8X4HzBKsFw4dnA
WIVy+GobEJ8/12ebhViLLBC12Ulz1lttH0GuNnP+ZLiPWgHrPptrWQ9XWpkzh8O/zjnN0//CVBLq
QfcyCx1bfRaGxC6ss13t3YcxY38GynP6c6OrdAzRz2Tm3fd9WH1x+p3INQvEnDj/MDVruSNX4CiL
QeufbCGGsEZFM9VEDUdAqqKLhZ6BTl3VxvYGOc3vsnKj5KJk3wJRvsjn9bCW3FDg6+nVrIQj589A
3ywqkOqMNE6Enr0c1JGPFa6nhaFGXUFntRJ1zqfePwlPiStcUW+3lt0iYtVkwurLUSQp+AvWe7XP
yFdarhuyvs27Jnfte4/mG9XgK2Ku7vx1llSZAIJfAczZ0wRIM0Sk2M3tO4uL4TZZFiqBi4z1F96R
Svv0ik7bWaU5HGe2LyrYpqbBSybLuYHTf77Da3SOl/UZSb4TCJ7AWXsRqpq69cGKDlhWMvjYlo0m
U+R99BUIqIX/l9E013vMgxkNfKfmg2xqOrTj4dZvIEZTkMaogT4j0A4MK/RNE7tw7lPennV23Og9
ipSkB2h82UZ0+JMLk9anJBe3eV9jIIXhiOEFzqIifWpzYhmp9yfKRLKfrhjqeKiYoxY9C+6qoQVN
Q+schw0XfgfI00sMusD3JUVSXCF1tW7HxIvkILoHuDqrd8coPJLTCoZYoJicu9Do6Ud4cjiZ59Bk
ZSOLW6/NyuyWF0hliIVUDeU/WS7xDNxPkTlb2EzUX838Cq7FR+eHu5fDQz3t++jlquOmrIAOCsqp
k9sqyvOovDBmyBRIpnpZu3vQVlDGMKXEmQ3JN8VDzOs7n9kWsFi/OG2zua/mBIjKfYq1OS1a7AV0
w2pcicCiJLZSDQDDBUUaaR6t9mSlR0t7t7FbhTX6E/3dJ6DTFrhUJI+glCjpS30YMrlGiiZKrdor
bZuEw0/c8NXKEkAx+ViYqiYytRueqyWtx+q+mN+FODDsfSW7NcSGFtTU4I1m+h/4H6sd8EW4Pq+g
TghCNOMa4EHfQDwgCU68oJkpSaxJ3m1Boa8fZC64S1HlcJ28ZtlIkLnjUo595N/mCXk2ZVTvwDSf
2NewtmjG+EAI1mSTETmMqE0+/4qN2+6C3JgvzsCeWPLKxUsj4sb8wTEwGimwNJ1P4JvKfw5Rb0TX
Tx2B9h5dEsNMn0PvcHNXfzmwY5SOzR8b+55sldz1LMkqT7tuQOg/a6AeRgjw8PLvXImYQvLlVU+b
3Ba/XzhWgkKdoHv7PGdUYuwp0Hh499QnzUfrpeWzQlm/hEJlrAlST3YYAZuikVkI8ctNbC4y/C9t
dqZviqFtxV9RM1luIHGu7ptFlBZq3ATJneqhueuh/l/LKYmwXDKlMLO1Be0+bCspePlDj6l8cK9F
FVptCMr6e2HfYejmXAncjNmDXDi6qrlYZYFmdSEgdHX4i7aeBToBlrqluk0CdjYN1rmDxnRgUcKi
LeWf9xvXMyGSTMjMLnuwg4ZNVTUNzna03pJRMkpvtyyGCFfLdahVH6YUPZ2B0KpGeeL0/1F/ovB4
sRCaAb1vnoKA7xXH2stYIgrAdXoBNE1fKx0bLceirKrXcMgwntMVPtaFjb2X0K2etw7KPCLGoqKb
7R7MrmlEZjnTdgtkbFU0pzPIqA6ZNG3QlScQW27zH60AoZ2UJEG/fNRlk2CMVf+HbhRBErde6gVZ
B+HViRW8OF5GANLzE9Itk/DmcihHvhJO6+yq3I0hLi/p6UyKNz2RG7D0gxnhqqHQxcL+e9piwxGb
PpUvYIRjuL8S6bxMSo9ds7AEydYa4P7aukj0DPldjUnC3x4Kjg2cAVHiiqZfQeQvhQ0T/YmVqqNb
PPJQgcxQsWK5aArHJHCcf/5JetiAS+QMs9v3XxfQJut9hTZcgxy4zS7TNzQaLZQq/n69QZ4eWpVl
vUxSBL68IUOTU7ZOpgL71RhpvUzTCLmM4F9fwSukpr6NHlcGUV411G2I7ml3yl4tTEIia9TOeMym
JGqYkkyZJrsq/DuyOcwmg3uCM3DvmgEEfFJS1XOI4aEMCEjI5jwikbV2bMeX9sRvAKU6/zSew1SQ
q4NOxMRfvM4jimnv9LYO6skRQ+lKyGQR/2GUbYtL3508ibYRPBVXwrkct3wce8NmCrrQuxXQpE8Q
K/EjWYl3i6cSc/ZMZAXs4JTP0OXDWjQJTa04GRo4Fry3PY/dIE3NkDWwTHd6F1mKmaqlLMtC0LG0
/JT7bLgXlixGWNQbRJ2si1NiYQMJNIUH9Kjm4oY99jlXlohAcX5V3hYM0KJ3nR03H00r3jTAKUOM
OwWrp/Px9vX/Sz3rWatqqoFmgMJuYIUVcB90FR9LcBuwlcAu0wpe+AXcr8b3AM3aY6bxraWt7Gu5
nur0qfC/tIcS9DH1YqLyBFf2X8fy6VmHJd/3Eaw6uiJQoG8WRmyXT4ohSmI9e0SN+G+RSRFP5ocC
bJ6k4kln3vSMJj8n0UVEXDwWarmfoGUqD9il0zYlhazos3kf16NHZRVUrd8m/8jwDRI8H2ZSp70Z
IpVNE7no11FnWa6PrUFis+yvZPORfVM+x9P178RqKLN3+Mw6oZT2Go6KjgVtJqZL7nUUa+0RuAbm
r7IgfGq3+Mgxjx+uaWjIGnMX/SP/tOZJFACEFoXVZQf+lF1RjWqoBnudKMYgHhzbdnYEfiA4gX5f
izxoQBfJqKG0eBNHW98Qu7fFXpmyzWYWJMOLQi4Y7qxX2Kl2lhT9o6jSzOGmRrNVC1jTG+yInETj
lYAG3lW3Px3WL7KJTjPgHk/KOP8sMR3pKqSMbhN7VsreCyFjyuw6aDAMeXiocizPYRqdxwQk2zvG
pN/rD9lTulqNc4mcLVD7SRrNajhJqMm9MIg2cllqVZ/aoUcMXCF8YHa02FCRWMIE2OJPHWyQR9rK
aN5ogx/Zb9U99G4Eu4XLRBIXr+Yom9J4r1V8qLoSRfbi8uy+R6O/+cvY8kaj18cyPUcxsMxPr7Bj
GmToiMH5sr3vf1qghU9BoJmTywFUY/o59/jNCYgNvBNAxKIqizlG+krIuYnsxL9vZolxFwQQQo8P
esA/sEfPl/f8YqzyiPALIDE9rmSv6TNVOA9sU3sTLBZIWnOvGi4EeEjGqqW1zF3i4B8OYIwUIjK9
sCnifSemladqNijF/HsERiMCrMFXBk4ooBo7wE3GHbWtSOBbGUWAR7QjibV5W+vlL9q77Oar4HtG
xVWM4t5oLIY0OSQvu7vapm49RtZCrWw3yimw6UfwBd720slGXlvJGcFa87Ttgbu2ibBAkT6essT+
QZRNNHxVorxdUqkATq1IIEX146GBoNnAytO2x9JvL0aUTyJyCeS3f4ih3Bc9OX8DYgsT5by03NIy
4zyR+hbFkXD6F1+MHkS0+tR64NHURuf0YB9pcGCblxm4iRNapgpo630lvlPkg/yvUZ76Avao6Tsw
XIsZzncUPnQ8aBHBh8/s1ZWEirvsL1qTV77yl4V8pIvGZYnB2B2rOhbGKQFsLGfxktcgwcVCxON3
TD7Lgz/WxjrzewQkulVHS12KXFKIuW0mhVhw8XFlHq6+PelBgyGUqjivb/xAuq1hDXX7UfPCm4wu
mCLdzLKvFrERHp5LV6zsnwULszYx++AasGp67Ky7AFovqfG1ME/H2b0d+oxfDbiHeW//Fc4CuFJl
RRWqzk7N0UzFXKBaVxPVGt9fMESheXoQ/YMls1F5fkXiHsI0G6fHhJkZ8xcm5JooJ+SB4CubZPsv
5rhVJJcKqFyPDAM8XETgbh6ElsDD6aE86u3KO2raPDjX0hYuTX87b88+yDV9yCazkJAmp4ecMQ4S
V8wbFGOOzpvhBG7zrSwsx7TxHoP3q/YJS/zf6WYi3rbrYaFWxp9hUKsZa8/Y0t26zjqQ+XRf3Izg
cfHTQaWamOV7+K2LOPUuwBcRgP334W0Yisp1aS0Mr+bd9El83d08ISGkq0/gQ4IuJ5QFrCiI7mSr
vdWYY/bx5izq+YOwcaxSKP0/xtzfxHTD0C04BSjPDnC2cOv+mdv+Fawhfa2M4xGoG5jXOi0qwVxU
fbt7Tz4GOlNgPceNLea845aKq+NrytCkToRBz7g+rkPJ31a4kOdmYm1zqSgaQFUm3xrt79nIH1WB
jCF1Pj6covlHP435hchUVRaept/Mmutapait2XbAHo8KL61+PlPkRCTMLm47TGaCOmZeolsjCeSH
mvdYhB1Dtb1lJmktKpfOFcorw7r+cFBqdIS6HMQJXhh+n9xbXCOfs+Nix3oq9AGTmBXIYKtReLLV
UnFDULORZtXIti8XYPVmn7bopYx/mOdVhwA+AUZpYhbTN/nlBcKkAJ56CSnD1Hfs2UI8TZOMq6/U
xM1DKTSpsxEf7U0AaatuDl7glripd4Y04kiBAlSS6IbS/xbID+owf3jKBuXe4SEljsR9oEAh5D/A
2943MfADIlaARP1piym4gcpXiWGD8NPy/tNnxKA7ssiPHMzYue8Z46xQIeLgV7RieWEy4WqRLVFM
oVZ1JR/1GD3Vsz8OyrYQr0XnjmxaxFeLFjFyHylGw7oqjBeG1hjbwRGgeLqRWV6xanxSsI5YYHh7
0Y4fuYdkjfC7v9lXt/62G4w5gdu1vf5swroxs2O2LeESrVCUCAWKbujTRGyof65uWd+pTiYoFyRH
73Eyvc+VyOLYv6Hvp0OItklpsbygVeLBAkUWKiKHcEn1nv+qPRBA3NPxFdQePDV339oh2M/WsWRf
HYqb3bMm4mSDLIZMBOK9WJRqMETapcFjpCPRxBMQdFyn4d7K6OMEyKsoGHjkFLpL+V6gOTYg+2jy
4e+wJWaraAal2IoYB+BwPfVLU5tiSKhi7w1CSbXyTVQPSmDykzVIBQaVMgbPf5z6d1nQeoDVLpPH
+Vee8rqU1qB73zd0u51NlK23UkY30Ks4sUREX+2JxeFeNt+RJ1zKG4UCF+Zsi43TNchienCidOoJ
6IXHEWneKu3v+6sa0yAzXiXrYIOsQvIMKt5HgBtNE7DVLkdPRw3BYAnY2X/uXFTEYqCoS9QlpKDh
5h6itxc3iCxIE8Urso1V4KWRxa456FHyDt7UzPCcwK7QcysFJodDLRKNC6B70sKqh/Do3wUwNriX
dhSD0/YWP7s+4ypnKfQZMYKC1TvjUMrVClNi2+n9p6Cjtskr13i208P87iJAR3avPBTPHzEy/yf8
YnUecsNIV8u8ILsr8QnS7yGb0zwH37+GIw6rR1Y7u6wmmvy7C8v4wPP8Ef6lPX+HZpIUFnXy9Wgb
OfjCkKbNyIEeT5cAOS1WgK/2q/r+8cIgD7QRuNDirwYMYYF6mtJ95nETJvJxYvMZSY/M7TC174Vr
/ExXMeM14h/exCwMlJLHhBqjzqtr5cTdLbNsq9RpoJxBozYkzrCqFWyzN4VpTEwAzyvSHyMskfVx
pyGwxKEnZiXd8+CQ3189BfYibuBTsY7JH6Z79YomlaOlEhlqFGkES93BBRK5bhQqhJ+0DrMmogTT
aoFVxkdbyq1ZZKRC6Wn6ECEGEsTIUlFlRE6aW3RQxi58MqgRbyhSfHHxz+gxCA2jXyHYK2Gvp3b9
iH8xTdyUlw/j6EVFeuI4xzsmXaNNHHrGb8lQqj88sa2w4YO5zliNzjeBJ2FGcXxDaNP03kbq4DnD
TSqkfpPwB7tkEGK/F6+PDbg8DL8mD3VPdohNsVYuKy+qzl2bSIv+OmcG3gaCA0fF7TOo8dh0OOhn
WTdfW8ojBJUroaoYW6zEu1DzD9yhfPxoK98RMwUgLlmzoQoI7QSkiE83lLmmVT/XWs6NdZOJF9SJ
2hSbPW2vACOn/82K6tVEjcZdVK8K/Gp1+VTdc1DwGFJQPmlXlWjh2TN9IHHsp28BiRpdi5cYIMA/
TfhuqmUDT7gDdtN+v1IoZ0xV9cEMjKc+8yf3jV9Rjwz7sG/T7FNr/Jy5f4xhLIpRqSZDrrsnVLqk
1UA0YRrsC1HoFQ1pLXadYfovkhESeBZLyzyESbX3aGzmg0lOn2rn47tZnG3qRAH55HHn8DLmlRI/
QY+xhv5l6LxQZgGXbGFVIEto9Fv9KsgJCe2n7ATGC1qBFxPc2ZFVYuiaFyu1enJ07GkmJ1msFZab
7xFjIoQYX0rWT4jWbNU4KGPsgvmRBourAMDZOjdfSvbWLKmQxZdEsvwb9mbj8zJCUfITNrj4b7GI
PewCBUArXKMHM0cLYNJHSmbf3ir5tgoiv4aN0S2gKfPD5r+LDbYN//eZ2ACvTSXWfqi+bZxzxt0i
WoaQ8nkzRDd20zclIDBrCbf1rP2MauwSQrJK1y1ji+LR5uMBSNyTCLT0A3PgacsmdpWAtnboGsL1
/knKQeXQFVXFuzp/FeLa527VZWLohaeKi/9nFnWEo/49R95OcL4g/sw3BijQz1hY3dqhSHc/5qnz
TxZ0/+QYuKeipWW7rm1cfXXlqWZhb9GNARfsoCFt5TMKlg5JN8QMkkIY6qNhPgrrVl7kIHwUXoXA
OMNLyCgsxOWyr3re8bMvV9IAF9T7ILdreBjmKcd3LvHb1ClIoyodzMOgPhUkVzEsOQ6+Ld1TxMCT
wLLT4RrFhUPpWfXN+Pqa0jideipK2omQXUPJ/00IX8RaDQiPNtOWrq0PP+e5XTwfsRQYXBm91Bf2
t/25/NZjVXcY+Adu5c+qddGRoXITKK1GqkvV2S9iL6bf9ilsMjfX371HIHCacCrhOPJIiOhhFNcY
UxnWOHB75oiuNFabZ7oC886GTixkDnyf0sYbVtdlIpMNEcTlXAHd7/xCYODXP4MXFTIdI3PNWd17
dPC8s12sl4slr9aRYNTzB7PwDUanYlDNAe+UMX/lAphRXLwQVB4f4wPXQMD1UYRNIbVySMkPgMxE
Lrm+tI+iws4gacmOfBJrRmHM43EJYeG16Daevi4Mi1h2KhXdLy9Rbys+PRy/Th4kheC0wxk6DPvg
bYdZ79CpgEL9sFKtsjfDVB7cq0/5vzsZlagc5cXPXL9TLAGWULGR6qUUQh5w5FrnBrPVGNLj5BP8
4cNxFlkH92IkDNqy0sKp/hkLx8MwHtcYj03n+7wOUa8YUFAToJmzHKulc3FBx/pKEByEfLNzNakM
vmEo9a8I+Wk+MFK3e1lsetNHyTE7q0HjPNDqfb9aSYxYVSIF1oUnT4InOAmihgRDc5AFkoOGTD64
3Gurt+IOmCNuTpTf5i2nO3y6F2/pKHyXVCwJyJRuXfTLq8K6OfyKg2PMZfI6JleeneAVf9MkEKOQ
wHTKykfEWO0SN5oqMo4zYim+kCKO+v43cRqF9Z3XMRiB4Rfd6lbNS5YenjjHi/RimwXgoPdGibvk
99o1dXUBvEQ7lqUnVdXFwvGfOQliAKjbqqgNPWWoawdkZF86FUeel/FcSPwMbuCKM+0VZQGP2Lzt
Ik/TTXdkoyX31auR4mWGHhDzmWAM8lMMuGvfbf/aGqFVW6uq9Q45ZyKqYXBLeZNql2S6kSq4KQsO
2fMui3c0cScLIoArmV6HMsefnh8m4j2bLATF/VzwbwUc/9IhbRIvz2QeWmqfkc7ifhOU6zFKLtmI
lAee8WqM2xasEyFm8AVj83v8CNp4WLJPLJWg1kE3+boGfzkzsETIdtUAMbFK6vxxHEO1d6VhR/cH
KAhgOPmc+fC+xZPYwWbkOWr1lgG8USn0S26w1bhfTX/2OF1Oolcctfi3Yz7K/HupmGDw6fR3E5s/
w6YzE7WYbKBNN5C4Ai63+Id+lhCDqmkukqPdoQYqSjjAArqbpeZUXXPbqEGT4Mz5C7/+P3du6DLY
rr5pZoM6sOSana3WG8gLFWW5YAVdkSMzKsEnmcAHbkQ27i1R86aTLvAueZefZ5cd6dtHafdgrxmT
yRYk90Tz+rwAMtlTwQH2El9BouLcZWco7O/TFuX+JmP1W9MUxOYmGlbWrBbEZ0IZDJ0SdvWW/9dt
+teoFMuXWJ7bXWPUh+gJ41Ii4kUUzHbzFjkZJbrwmoa7M7HkZEyEYQ8dC36YH+zrRrp2OHnjbCoW
Gq1QAZV2jEus5iytoIFc5memKe9zf5MrM/4dHn1QwhBFw53a11fs1oOdzAX4qHsqe2dYZbVT8QGT
azGLyQ5l3B3RtDlH05UJAX0syTtW++yRbOZML4pyMMouPhcuLEiTvP3NzouHDBy1uzJso5H8GYpS
ddbtVMMfp+SMqb9J9FcT8sC7TGLF9KJUbW1Y8DEfJQmuLK0FHRiQR4pJu2Pr4Kf1KS9NdqIAFZ+T
RVfPxMZHtFCDuUktZM9AQ6EegvaseHhsXtYUpSvdyyNWLu7tKU4oNw1ORBC3AHGD9tutIYeW8mAq
qe2T8vZbS7JErxdzJdC1fsbfdx0cpjZCCM3bZHsdsp26ULcpfb6D+WNKV+Yr27KvWGl9sryLu29N
KygQXd97MgybWsjU1cGjbsgj98lEbr4nrTs91BquqmIeSbyPwGYwQ+S8/dGHvUx38bzI6xmYg7Je
E7jWdQyxQeSofePVK+V2GqY6ViwfV7s5bJX3vBJYF1CGWybIYgr1EceWTOFxyryMEKOLmDK2t1be
EA0GtoooLT3gN8dUSOEC87WP4su/B5aO6FK8ysx/dkcDlbyHMTAJTYKVAtwC+LOBLUH/lBIiC0zL
orVHM3etqvcwrNBhkqIcr/8hv4o/WDhYdXbLkN3UZDZGfCTDksp3OD7itvqfA5sukEw/wAKEbBNG
Qk9UN39QANmw8m8XMgja4yDZdx8H8+/EAQnYs3Btx42B7CnzPjg6QA3fN/vnYu8LtealwOdy2QiI
oWrLKT3EBny4Lv7mN3fyrYxShsDwkDMtIcXHL143K78R6PULVHKUyr5jV6W3t3pQ995c7iUyiYPo
og8iFzDflOeEwnB1xW8ZNuRiZbSEvfYLY6Q/oMhbi4UnxpcV8j6eQHxtAmUI3jSjhWnW84PscIdi
C2gzXVSoFOLi+16dNLyQxksc4PKRVOhlyDTdjqefEFmRLuklOQIlabJh5/ORlajBUTyAf696Kf4v
pwygMlEhGMI05c9D768NVdVe3bxnQLNh0xMkuDBLoYZt6ZDvC/s0wPgyBF0yylzqI8G2E5zUMYqT
xqORZ1sraW+XFqt6cLgO6u5mDyI5QqgHk4Pgeko8L59ZCChheVmAq7tVo5zkcc7YC2U/3rh/Fp3C
7Ov8wtBzKcmKamM+AZwh6lG3rrD4gSTiUBsvJw2ufT4+lp+Nu3DovtvdfclfXnNuZH8ZfU9Nr/lU
87FDaSxGI4yEAo6h5rH5LzWvp7ci59i5YzXCrlgBsYXT/DijDAESZLHIU135mDORHFoT9c/exs9T
yf0T9ifS7n8uX88cvoj04ln2VpAHR+MXN6WFeob6UXvI3ijAfx4WR5BszLZRKsaXLZ58wgT1yhhJ
qPX0OR4R2w1uveH7SogHuAOsJfjv9kGy9T541+9lc9FxQab55aL3IyXZh+KEmypj6ZM38d07ZsPv
OvNEE4o43q4pgdRSw9BdEliUqiKn0Qb3qifRWyiJsE6OMKNKbZobV6ZUUtHW10MGEm7JihYgl2CR
1nRdy3oI3ar84O//Sqv2SGK7eCyxfdNjzCw2TD6aXhdecG6lFGA79c/RRSVQTPfWzuwkQJPEKp3p
Ae4FtZKbf3Aq22pCU1me2vccl3mWUA/AdYFjXhVy1XSLP1OEOq9ttaLI60RbuFHAYKtGhHYksK0r
rxNchWWqk3w5dm79cMT+G+VOa0lpLdW13fcW6LfUbUXts/D04Kdf7FD+ycRQ/uWOhxB50M8mn8PC
uOjYH8XzKh4HAm2txO4sg86P4OOyeT0rAV6pTJi/+0l/3JARTATeFpLk6mEO/xHeePopXbJLmnbp
6Z9Rc9g8NJylU52/XPmiXPEoBk06E4WgQVrCiqy2go0fCMhpXvG9mVtqXLztzonr/6vsZNL/VgAz
z0e6MUy/6ve8UY8x8Xu+ClKH5SbZNWr2142ND/NE6h9nPL20LjfiAiHRiUWt3xZ1u3XHlAuU2jTD
5H4WJuEhXqgHV/rIboxV3E0D8SKMPrLfS0NR94i3Pcj+cj3eSOe1IkLTEz74edMBlzyiV28ugvuu
IDZE8kFnlU9yzlLuwR+TveMsKw13xOJWYNi9a4V9maQP9rxeQlELVFzcUCQRQGMsH0ZITo6LnTbu
e9DXX5womdanZlRHv4UR9X40xun/MRhlhD87xP9Bg0y3tuuo7lZEwlooIy4/rMC3f8K+GQzsfCuU
oROVJlYEA8n0srw+FByvMoD0c8zmjUSlv8YqFugp0IuulT6WuiJC04eNEyPiKfIg9NWpGLXepCxV
9BwZ9QO3RSdVzGgxNydZPYJcTcXm53t33bNwFpk0A2O/6pnR7xrDp6DR3I+4S9uX81U+pH+KUxWp
bkDBMmn5f+6EESLnPSGpD2HZEPUYal9F29atAN/iw7D3cxviNYve33ckKhtnR/C1eph4u6T78Xyi
hecIEO7nOwFr7jTOjiOklA6WwBEpQVE77ODPz19y8a9m3qS1Ow1brhFTWFtXAhp0cZCGexPx9kI3
QuEKNjNrqBe1ZfZV0eFx5DFBW2+aWn6jg/el+6Lh1sGwE/rdeVcJ3gt7yQiQQSr4gbIuy6NTiF6S
WUyg+B1N+qI6YASVb+2hsRSbO7wzJ2XYSACPcLfNMOJ7sWU591WEcCWmfphNFj8rn29I6x6f/2dM
pBYpzA4+qHaWS1Q2yb+muAXCW6ihBRyyxZuELGzLaePalbcGFb0EmLx46RWjvMB0E3lVaDTaLK4u
m66P6w4r6G/jGMQECKqCA90yFiyrZVTLRKu3r4ZKPCiv+rUkmxnEzkH+d1uLNw7wMx+e/iMQ2wQb
kjBS33FSZwNvU0ud+IxTX/AobEAx2WAEtRvR4yTNzLeYE6rlAdTyvaf1UyQkqlKV+YatgyJzMBr8
vohgp9mCkL+AhMnKuamIHplmPMGl9iUdRcaQEtkWdWt2FTXR4ESQOR09C+t8prk9/9RNtdWz0hPJ
G3wreVXv1A9aXBO4iSaO6Seq6vPnuIUCCUW0+OE3BQYWHK5eBMyLU9f3fP1MSzynwprgQHmWkibQ
qh0tAEybdWjhbbpiLikyVt0RZtTmxyZjAmchauOe4g5gsrLiMAfH3HchvC2D7IovQs2hLa2+8B0c
DBG5ltXNC1jLJwVAUoqSpdzBK3PEMaX7KdmYxx7oNQZJ+vd31FpIjDR7lXz4uVPrL/0b6HKMb6HY
gYwsY7THvZGXpNLOGqUAjV+x38NtjpjnJPqjWNAMn2VasRCUVeu/5U+DHvQTmCteMkBQlXP7b5gd
ClMY7mRG4pOp1mX119Pav66smnukfOfx3eii8171GoqzZY4LYq8rd+vCrv6G/8d2bzoC3c9D8vR1
aWqk4uJWkO6EdhDP4TmHvSATzLFIcXzvixD7FIvgr+Um0Jhbk4TXJo0GYBmEs4cntlZWe69h/MTi
SMq6MBlZJhPn78dbdVYRe88fq7Iwz9v/2NTqYP1245lJ/M9YXjKjR2j0kCjNW/5aG6ARGLErbpH9
FnjPgzuIK/XUbfSlRcz2AlNgannGXSQ6AwGiZ0E/7nJ9BJbNdgfNBolPDOmRBD36la0yjZbKA7ru
S9yLDoAPqWZz6YCkHV9j+bdUGNU4JaVMpWy6mVA7NgqdXRAPGtmdKxeOBYW/TGHX8nWRMAc63v1+
41A2/klixRWx2Uknclus311nSw+gMYe3abkY84QLFEg2ATPZfIp/4+s1Gxa9XYbI5nrO1qfUERBw
GrwUQ9VCkxImCRsXijR/jx8xB2eiPlrSXtCXDgh//yNxrRsKL6Hbrt/3CyCYtboE3YoXicOddbkd
6LOk7hBGrldNPebqThg8vHvBAbdu8rVWK0HKfJOIONCuFQPwi8wdhAw2pmpg4SfKsbOhwxbxI9Vh
SRxvrwYmRFCIG9/UgexNQlPDPvNwxwI7hbVi4hy7nnThOQmgskpShoz1ZlngQyWFiHpHIiUmoyI5
dGDt8udFa/rXP+AFZs7KuQImB1i084WJJiXRyHmvYTYoqT4ITRbKF6qO54UVTFGenZ+Selnr67uq
R1GhH7f36ACWi35Klw6mCyW4+/mztvwYz7CseNGZKsXkrBplmT34fcY+kZhus1WyMZVc+1O4tWRg
izYDP0v4ALd7W9i4AvNE8+jz1eNQRrwipu/gPv8pnv/+IZvag2XYOG3YakCQrOWF2FR69i12A247
u9YHLO2UBCCB2vCtumq0g0VUv5+d8gkn2cMd/B/2d8AUHwUuUutGWLcGflPsgmH8OXaLGpbQdT5E
cZafynJAq9VlOgaXL/GBJKJjx0un90bm1DzbRFM1jeYB7KDXJxCB6jdeKX18+7tMCRf8k1vpqvkU
fkQA7yPZIBxmRqKL4Pd+yqqH0nAedgoiCmATGeXHTHS5Rf1ih8fAb7AFUkg+621MNTwMkkEyhGc3
NrldwO4g19wyPqZXNrYt/aaVwjInj04vvgbwYjhZKUS8eYg2QMucOagRQ2++fMACHmPK9Ti2v6Ek
JanFzYUT7fqsFlzEYZ4/nF1JZqQujh0N1xIF/pBeF0qr6kQAA8ZN1pmm08diW9WXn6TWN/kzXNPY
+76mCNibK1UB9EWV5uxxw1sgbz6GF8Z7i1eH+ARAikUDV/nipnNzcR2ovT8Rq8EGRdBZhB9K7wwU
bfpNPptvyVqCDTzawiekFMLRvpO6VQUtEZ84Dlne03jg025zxrsIBY3FnvYIje37DRE2f7FleRp7
MNXRlePtRkWWfdtcoa6oSJ8oPnkpth0Labj7WQwToaqjrAmmWngGSrNvcpzNI7SXs0FNi09iJ5tx
1iF3zoPi3UvOeKE/7XvVIPaeaOpEuWCiQlg3DmRkvErW87HcplvN1qvQPknOZouPj6k/Z2mssrZr
wmc1WF3rDt0agl2wPon76ryriQOZDG4lQJCcXGn66SAeIeJCCoqSo3nmvAQnYnJyCF28ew5FvTCR
nzflFCY26GbtKaC4GYcThOYeGLD0ehv2g6o5lxjAt3rjyIobs1WRPLrkGF2p02+ACrE5EJaTtHuK
GdAKz9C8VAMinqgW8LpjIPfuYaWiA/KeYsU5sgZsgHWVdHgsZJ9Cv93RJih24XqOKWxXn/NEzRCP
ORy6nYyqH8K8Xd3pucuMea8QgNVefx+aA1sD+vTOe8Nb+/yzZYwmmwofJEIFaUL/gVW7Mcohpvuv
5Od6fsr9TT19ub0zTt3Q2WK+/qFn4QL4avmUm+wQ8T4VK8mX3rZ76+OX11p5cZpezzP0zvic+sW9
s8eXLoqlMtYwSfiG7dQMbJKCTiNriDV1cq6bGTH1Y3WyRZXLNL5xZtcIpOFU1jk/Y/yPTI0CP0Nx
BX1lyVcS/X1ID9m2XfIcmdFpThxHq1Ds1MRdjoDXxyGSEdgr6wenFStLY0xwp/3+Nhon3+/o74MK
rsqQqvNi4rx29aKMTtfH32Y1mlgzUiWTElB0RsVOeuvRN4TbB7qwKTnTJu2gAzJ/jRRrrePQQ2jk
lQ5ynW+Y1hLbOtBPlZYF1KaIouo+eYxgaqm5rD7ejmrdh95VOjJjMzxp98ARQA6ii0zo5dznhfPi
GWf6Cwoe2qzFxEJYd7vjGgCwMy01G707M28jl30b90Q0ccdqLgRkN1ddRbT0DwmtTFFkNUVXLRqP
HPNGiM4FD8DAQLIGHRqioLx1Qa4wC6+qV/IutqLXx1x6Ohsl+zutCid9q0Z5iPOaRC5tR9skhATp
Aku5bNu+YA3fFPXEwk+sncUNx64Bt/5XVjCueshuvwT9CAdWwIZatcd+NjG+IA+Pf4javJahFdjX
Ft74oPDcCijfMkb7kQgNvPyD3umKBCQBsEh5r77n4xmjwTq2c3lqpSvekzUfES9FtHa0e5SPem1e
CLNwT8hE2asuGttI4a8vEHhAjjRnqquH2klw8cR1Ky0KdfwJWZhx0HfwVRtaUdhtkYwyKbTdL8ca
Os4G2M0zi4Ud5THQ3J95FrX+XtEWeYMLS0wMwMJeBnTuzH6olzarfo3F4BmKdhju2N+IqsTGOb0F
NyEZMlfzdI3fttmndUptFx2lSNv5XgUUA0lxleU8Bs5qkQBXXiOLYYEAloPh5924aOdF3cEIh4aj
OPO9V15WH7g246bustTNeCQlFOccJN1sLHeH/ngkenQD1AgQgdEiIdFQXea2oFtUnHaDT+QYgKJJ
Fd8a1+MOYr/Kp2ruojA98mpLcXZ0uOJm4G3yrXEDileWKZcRdfJHhns6d5g/qUzaOiFZpZRsxAU4
ELlLnyLouKrLDxX03sL/mgS4rHGkacjG8w4SsOgil+sPvaFPBpQpw6iMjCUgoiYFFQX9qLkH/3fD
GndN03qm06MasRP0Hqoc0wtC7Rar85de0btxEPxq7+FRnch5nUdS1sQpfm/t+6aBXnylkQwoGGiV
B2WnH4D802loReSaqMPdmoCZnyeA+e3m01lt0CrAMSQ6hszJM8xlMSErYeMy22MI7PX1Ym38wkPI
jETK+0xVXzf7yGNlb2vGCjIu7j4mqyvJswMAi0YVn96uxmPf6sSQpRxigC0SHbE+Sw2mXaB73uSi
HaYG395YmhSfP2DBmi3r0fQGwxEYJYN0gFdDT2d+6F9kGW9xQaaLKD2eSQ650EhMzXT0VKeKCBzP
ybIVrSzH8GTrN5a9otuiS2F1gGuU3k8mw+RbLtH3r2Jfu3IHgjQOwch4kpPGzxqemcKdTF9wh2QI
Zv9dQAJhNDHUkTriEbFEzQBIeGVB2EZe8iHkPN0/SNgsnyR9ck1p1WaUt999P/VkWJuT9cP+UwyH
4Lv2rQNeaR250ThcXfA0Kr59X30pMjrHFe05l7vBhFFX3w5nUeuB7bSAgiBK6zvXkVi+lb6PQQhf
gIGYidA3FBy/cvXSZYbxbiOI+/VWR4yMib+fUyq3fHSfo1K6sfZ+1CPUAvgDeAcLQ3LkNPhucjq9
Fntdgau/4lDdubTo1JbBlr91KSMwuoQJAi4DAuZGVGcaNz92YPLePPDyY/dJC97J9MY02aCfyfZS
keebtXUGfHpk5LoKQxwj6HP+RDp9PaZLSVpZYdXImukckufTVF7yIhCQ3rs4Ax2kC9xT8Cr6Fxd6
LQwRD6nSYBL9h5Oq1ldYx8qRyaPP5gXusC0vWrl6j4hNJG7YQsUnvfEV9pB/rKpnUS62EDigUw+4
c2nOBrM8uW1OLsAmR1WVSIxaHkLoJAMvvxB9IxLCAN/+BihZYWsS8IUKyehSTCrDBP8PWCfG+MK5
6eyk9MQr3UzFP5C2YadqSiIZEPkGidDnFvOMJZPAJUbygEv8SqRpGMa/n/44EGnbtzF3+cNfblPH
qdLPTZCDOOr+vcwQaXdlTc1mxfY6xXbv7Urzkn+lDxrnxoeE/YzG+MOb/3Y211S1hvjD5QAKsvjc
9CQICpoepD3OpWV5rRXjztescvxOVJI2g/Bxkyej6BpHI0JdbI+rDa+4fNTe3p+gb8iRLHY3HXKg
sfk9sNazd3t6kLRyCEUrIrngq0P/J6DpBpjoNPoHXG6644Lrc28+Cdc921d0YjFN0D8g9+VePS/v
GojsqWDUiUHbxcLllyqDtym7gI99L5RVN1BL5GeRDHpK76mn5LLVm+AquI1fJw8ss6CgqTLvGqbC
1tQAuqCb0qyvwFOI33SNYTKTLCPeXTe/hcyzdwUbJ0DngwI2ENGlU0lv3GYzvwNIbFSkVKPgJb6m
HJXcGpRiRQIUZedm5r4L9t8giuN45+udu1wFNEaLp1zLdfqyKu3+Upz4+Z//wtQbhSD15yNR1ndg
zuLeWcwE+qQSaNn55Izi7p7t46ZhwpkAFEThK0Rkh4BB+CFMvE6+1uB3E/vk1h8Vx6ogIZajNIcE
P6cOnYyt4BL89S7n0G2BUykN276P1GVteaqF9PeNdIJNps1aNdnzAtFhUnqtNwBaN7B8sIBGQLh1
Y9vUENZKPXatV8RHW7TJnKTLy0ptJ7dfJeEGTxpx3BZ1gdAL9sDXEx/pJ1DDLxfu+fWP29FDl0Vt
Rk4Zrp98pvcJOXKSuSLzDIns4ddWB/5gMhFNxPHX3p/OTjBMJJvfbIuPn3DI1uZZnd1HuSDTjIXq
C0BeNL8rOqZfd4dG2EOneOS2EVulkMZkNazWLY44GjIMC6Gw+rkG/cUY05EGVzKRJK0KB8jasM6n
9+Ai5/VbqORIc/UYbCp6WO0iVSa9rWiZyNB3quAmD8RjyLiTletw7iUtuEV9hcPsuCrDEkuw2f6M
gvRGutE0OYVdXQy6YcfPAgen44x+RIp7dSDF8aN96h8/ZHOjmFHMKa3R4aMni15tPoILMBJbcKka
6dqg068GUJSh/2hsAiqmKXy+COGaT2RBm0iej3Bf9X9FcOajGFw5xLryWqBrNDVahVyr40gvwvYF
R+BYLiWnXJVUkocKN7bRdH5SEGixZv4Kq+v9RgBt7PvkgyYmnAOGLCWzZajvfW2lW3+yeslo073m
S2W+aGzJYeY9IUARvL64fhDfJ8sAN1q28qZCPoTOrYA/H3THKnVw2EPt3X3mZnuGlyPYCRZp6+KR
J0Y2BW1ua26kt4wUt6JsFb0byeB2BpQ8uwbFltSoD12q1yjj0Iz5Q7nlJLEniv/zASkCaa5+S5C3
EhAg1M1srNRNRVZInBfaa6K0vUjDqgQI/tbZD/x75az6bNFsxJbsknZnmh11GMYHGrK8t6Aw6+vu
LVxSOZKMM+vi4eLDeI8gAgj4RTee5cTqrVbcR//5v0MnHVgdV8EG05eYIuv5V4cWyxBEiDaq2Ey6
WgJb54kMqA4uHw1vtlZ8Vc3Zbmt0Qprot66VPmYVSsc3k44o8UULB6ogxqDHa2mG3ZTOXtr0YSPF
nNrxajzwuS32Y+YZKJVUjrM6VWks0H+P1rmeyFIY8r/xUGijD7bka1Oqcsizt6sYVyZVXvFuNHml
IH5ApFkb9g0QVefSBW+Q9+N7iB2Zwtf4D31HhYFIp+GfoAhsM1zRLEzV6Jl99mlTmcHB4DB33QWp
4nNiI0HU0+A55bMUJ2TvKZqpV2j9QKzyjKPHcqDXgPl0Z/WjtbpBofHM64SBMVm1isiTRylzNsoo
tf5Tu6NSEar2Eddnfghkv8qNrUVnZhnrtiorVjBZgY8/jnQeQpoEGYNkrH67IK6bje09goXD/OHf
6oLbzRsJhKbh1iNFWIc99RvMI7eC0u9Eew72p+Y4mDIz6MYiFfgsga+YLEu1wJGbV9gxiBpqyyjC
gnolMvIIQLCYrOMKAZfH4CaVTx+qq2oLP39PqtmF9eZ6oSZZglSFAcSfyIwseV9mWX908pZJHMWD
uTw+QNx7fVaM7Mf1V9BvD2tnx39zamyAyPA+G3n60pC8LKk2p4K+uocDwpiSjkO4QFQ9pcOBHk6h
avMJoaqsG4J8ShLhCjKimjrgiNN/lmH8gJ8vU8DPe1VAwoHs6C6RILcpy9TYESDdlFMoPaPn5wa7
o8rz/+svM1JPyG916pUVWQ7jDKhEjkawVmGEXatsjqWznN6HRp9ccbo4G3W6IWBckBRb8QIHUZiq
+TatqDDzws2UC5y33nYXzVwYz4l2Db5Kp0OK+8Xh5Wt5PAbp0DQZDUXF2K8iz0xEjCnCSm2Z3CLN
sB3U/uHR7++oTb2P0USfvu7QkC41xTGMkGXsXs6cLuCW7XezsBMvD4b3QupwHXunJaY/vrT2BsVD
OXaa5uMRx1PSSE3Ijz+MhTLZa7Mk4+9hbfM2My0411Lo1T/9odVTXN5AyIxMBZNgIcUaJdJQuGbM
Ae0H4ohMPlWuz2D/BGYIainOeHdOsqEroMtR1KzjJBwiZqJAUWja5cQoulHa2XEp81krlRj670ns
eG56QFHc4XSN0FtcfY5sPa3qr8bkOirz+fU3Dy8ZJ2j1KPrd5Vc3/5Tc+tcShLNzyFld6tJKYINZ
87Q6gvYB2c+3ydGB9VxXXvl4fqJqz8OldzQ4VdVLxCNZuyi47YV+oLqc/zaIkcWTeduXY1xso2Lh
Zn8WU7Yz4MG9/A/7SXoiSRHguRSes4Py9x3yYjow9oWqyARD5+t0pArXMsxQaovLA27HWoQMsGVl
jPGbgUQPM4UgB1zxWsZtjw8lzSsXEmb6midzU4ISurLkY7fUpIjEVnZMEGJHvmij3JRqiXiKsb42
nkUSey+XdEew+4cArQc14DrSes/yK+Cnv5rylj+zjKsB49/zdno96IjiQnsVO9JDLFW4XMD0ECuB
tGW6azP7yBDLsYKNQwYNK7wiWfUQ7MXRLGIIL+7hWkI4VwexwiKkPJdnbHddfjUyS2FCSmsg0X0Z
IdOZ8XHo43u5tYPFYkm1R+eZFQfP3SwbHjZcJpC3i1L6v07K3bwB+ozVDwIrCZi5P4ho6Uz1Np7Z
wa6DD/FNx9IIhmXaTJ2uxDkxT5HFPkRPSbbw4cqpHIV5yszR6IsexEqxZ8T/r7/7RD93tuyuUgt5
rkQrUJMNUgcK5tk1uTCyItPBUWqT3pvb4mj79SResB7Rltd+Rm9q/gOTtIVkykHx/4yMlhvB+HsP
PQM4kaYYV4KN/IzpQXGvHbqp2kPvOvJzyxV/XB4Xeg3HQKCW4WJzS+ZbzJeHmDCmVxZuOKDF9GXW
rGycE7Z0WfRO1oKaOExXJ/7+x715zL10LVJGobnka/wY5qmKl6QBRnUsz3ngj9iBMjJgGpIJlypo
vOSpLvX4lPeJetBcNjAcUqDQisNxk1MDn2arGBWi+OUP2IMQdYGMr59VIQz8GsMFh8uuJbrBYNyV
pX5u9KmjvrbZ+ZD3GFt91x653Y+2A9GOeI5XYm2KumbeHmBs6UzoHqXX760uc4nC1CG7Kew5lInZ
ecWHHTCxSQly2E2Ym6myMAr37qFRlp7HI+/VTRbm4t49eEvoAgwE9ryGi6m0Lbnd+/GfgquWdUTY
xp1ZmUxxvAT8bh8CikWF7o4FNmc8QSP/raNiie5GeYLvbg3AtrIq1GSCITqV8Z1+jxX8BnMZVkH1
wfPfNKVtuv1xJWk19yZWXEkQVQ2iDGivEWNXdFZJCWwD2PdyE/z5GxfUvl/NmVBYx/lCadCa/fdF
uyfVOZSgVA358qF25t608T+ytuypYIcKkZrWW+O5i3AMEGkY7x6B2x1eVjrV0DZ8x6aHRj4IEpJ/
x5aUMDWTTKWbPBJ7Wa/wftWUWOdDAzOnMXhNQnMJD/FekFYcYVfzvDxzcTPve7TQFrjDznq3U8qI
68XWJNzQx5sZsbE7gawBOYUEFVJM5sAeQRJgarrzqbSH30N2KYcDa/izMBEGIzilLi4IAvl54duv
x+ukh6Shpf+0YqmvMLNIVLYJ4VE22c3iIwKXFoqakNk+xO/n4Kyt6zmbU/hwKtGZ1IBXsXniqjzx
8eBJ6m4gUYnHwD51n/QP2aE58ahie4iSaTMS6xnvPB5FbO/JP7lkVCnCsGdmivWEP0Tii1hafWhj
+gcnqawKFTJbUGA7mPfQB+iSDF39EUOcLKec2fL5wAioycTHnboUqACXcDfya1wkBT3KRD5Dsx+Q
Nnc8D1471Yy16KfbsuBV0v4AejZBB3EA9HeVGY9DQ3rNtrSlrigimqOgamZrTNmeZQnvbJheV1SH
wrYanqOMU2Z7OzbmsYpq6oq05yuDuJNKC4XTs2S76P55EPRZSXnlxELFFnRcdoZkRTjATQWoXsRx
cdXAa9eN52Wyg3r/ZS9sZLpW4fUMOY+FwhK8qp++4dOSn1X3euKejaqcEfoqPjyBM6MyPJSS1PkS
/1g1MBObFRJMafuzWRmU2wPplk9GG1lHO4j/O86ZMHBlfrItkzULpKZ0EBWlBFiIvMtpzpUHglh1
xfftaSciA8NM8DClkYyDO5CNoRgNFc5L8tiq05uztV6GBvbhZWhjw2ETIGB2x/ncNyjmLiYJDGbv
LoYjj6KLCkjdMixUj8ox1HWoHiRQh3vC4wOClxnOCsUMqNSQfBfcJB2Jd70kAocn0+rqzOnOKj1H
fjkqSEDBHAFOd0yByadIARDDa/wQ09KBh1ouRKYrNTW1k+MO7m09jNyC1qCXvscHulSp9+ePIGzX
GiYkWVauSEJzdkl/UP2QSunX9r5rB7kJp4Z1gfzTqMLzFMi9ZFOx3oRtsAca6qb+vSjT5mHXPQkz
79RvgASlG7SmHEbEilvTztwyUBKu+oaTpDdgy7DhwgzEQ8DSM1yLPvjqXIf1nh6MsIn0EQvc7BDM
WxufaoaVmniA1w2se28ghPQwv9ON03lbTFqBEkjP/1ZqOhYHaO+F/kd3vopQeQ+08jfn9HvTICqH
zAJqZ20gRjIm2pSXQBFkPN3i42HOsOmUjCKCWwOAZESMV8tct0eWknpZC+6mTruEwxz03BKFdfDd
FyOOZoUqayQuVG7X2H7/WsgYI8p3a6DM7yMnuMn7l+QB9zRj0lrw/DUh96zhzQeWX4bh2+2yjNSJ
BnymUoKdjWMnc2lrOw/+m8eYTvh7MJriEEG7f8SgokF5jlPfTHpyWebEC3YiVKS5oTHfgwIuPmB9
5ZRHOz8zBQaI/vq+5k4Axdc0FT4e30pzL6jVK9hy5uZGCZCrs3z3Zym0wekDd7f9ZmvTDyq86wgF
weJ1js2wiBZag7wVrnlDjYiZUyUPwcVjk/FWCjlmCLZEZKeg8TcUbFe40A/s0CQ3ZhwuIOXJwUkS
A7qkmCbaqR8ValwJZDwDVG8j133G7axPZOGAckVCuYzztKcpUMZ/ICrjG1xlecXwFtFmGFIT1T74
P/ckGqVubQ0flLQGWohOeWtx5ORdbOoNGYHjgs+nztqCY209qgVm3xbOCR2qJbaByiqmeKmWl0pv
fjRhj7Raogr3vJ++sVeAv2yoottqz4oj9H8RhVEBEXyNJY+q8axPron8yU1tEqSr4hIGeetbZLnV
2cwin9fhApf0OQWqUbNlTLo/ZjczW1+TH7myJ9z3UKtUC0E0HRgOFsinyqg/OuUEr8AdtpfM8eYJ
K8wF7jwggWE0m98SOPYxXwJINidxQcvA9X1ijiCZ6ZjCYmzbHAQKKgUunUA4DhrOyouPM6my8Sno
lf76znEhc9eqgWKrJMxoAimHZpj3l3iGXpyMklmrxluA/8sAqedHH4Q/0eHPgR45ZoUOHpmlTJl9
Gy2l7StHR79PLONzllwQ/5cR0Ohp+69aP09mnlHrjeC1fsWjlojIEhumlyJmiPPlKGfRn8ZB/yI+
E4Obd/sQXrxgGs/SgF6zYECw6tpx56Ns6zr5Q3knxLN5imbA9RtJUh9r/LZTTmPrWvMS/hmcIhyt
r8q5/enkakyZt3fbLe4tzQTqReT19YlqX0/qZLTHynlINR5z5KzOgRbx4s+vLUq44/rE9IdKq/qZ
/AQSrajAb6bgeeEek1nBMPXISVLuZR5cZZNeFi2BRrVh+Hxv3vuUSFmVrK7ja8/1QY2BZ7Rlyh5n
sVHU632YVeL5dCkTOmyJXxiTai7XcNfr/O3NIJTOEWTpmkPcYgz5cD29LU+ceZ3/hWXgNjbceodt
Kf99dyGscTPIOmxD/cng0/43XQhCGCu5iDi+dgNNWTqJ0eF+2zvt1g6HiBJCHw0HrK18GaMJMY5V
lgbTGnmFC4QRyIUrHJ5p7w0thoYhLlnQFGv2oITl3wcvBBUyr76SQVTb+426zvP2p2EHz/O08JKD
O9/kWK5XT+xsxDql09wFbNhuy0riFxMzNeLwSPVBU28ckSxbe3ZkUjwuvvmswUqF2DmpTsZQb4UD
LXCrbCunS/rIOBIDau9IU3baMDgFJa8cAfPa5fo0+sD1MZNOP2c9NYqKQlXLzs+eSJkagksgcT75
bJNRIEtYZA1sf/de3tJGAqGP0EzBAFE8Mcnz5A2/jp0uVG4oWEms81+8zMswelWk5EOTjkSrJfZc
J8Cm93jKsXElvwd54NrrHnNccxB73esUS7hf/Y0FEtcG3ybdKk4DDS3rC3whB0LP10Zwobe7Sy+X
7ZZIPqbFUhe0j6fNTUHAPlrCoxBU8fPhvkpC8nvBb5Zn1da0ftv4KIKSIi6H7MijL+tyvaATxvou
BwowIqY6jUEwcg9Gsd0E0sGKfvtsw2P0DNDXLpnQp9QIPSDGFNFyErYwu81AFsprga3jc7UZwAlF
NtRxvu7ZodrnLY38o2q30KQRP1TGlebP2jzZR0beU71fgNosDxKElALkBBSrMs4cEMmHEfOPfIHO
NmsFlDPq6rwpy3s+0oZNNQDB7XP8c3s0Eq6ztN5j+RViMvmmezVIu+0lKZ2PvzGlmtXhBlgja18E
mTbhDeTF3+XjY9zGj9eoHj13g3X4EGE5GISzw+GfKqcCVVxl34M23eB7XVLl7VlQokVK7gLMUEAj
CouPoWKA+6vC3gOVtLUcbRF0IP50R9A1brjiqXqio2rbQlYBUUMFeOvK6UUHScUbk0qAfmBu65XF
sXlwj2UcPflwiBx7Rz5XjgBRfzE4F8dknOuFLneAdjf4OUDCPNkc2Cia29uWdMRCGWVMzchuM7np
u1WNjLnhMnH4NIznLnt/VsxMDxsNt2CKtPrSoleZrUpxApwrL+Z90b14izcOYzOzITepEpjn1iY1
3+oiCkTG8uUnPwunvcMaWrJqX3Sr3M6GW26+xyaVRokPgRU+kWjJNfwTr+I23y7vwHboUd4ZvB2g
8+lbNXPe7r/rU65XpGDNRertYeSZBPaW1nGG4ptaXhR2zkE54LfIEjvYWvbrSRB8DDA+aVLHFRgJ
FryRDk3u9fV1HdNmXYrbeJCBgty9d8qsWNPLewfyO9Zzuz230ShpuqHh2eIDM592zT3VWP9AuX5E
fEpiKa90UpwjuOm9/DOQHjEJ0WpB7fATM2v2fxGt6Fc/b60WfgRslFSkJgW5XUbEbZcAKMKsZShE
wttLYalk3ENiUzA13IKUnryjTdRSZfrX3lScnEPp+J2IkJdj4guxtT8A5/izJl75973CznR4hd5v
s5ExOMOTyJaUw0i+Tu29JyfB/5IBI6WtN5+iC0btMYM3dHdcYVW52oQJ7prPsS6cXnmOJZTO0M6l
lpU4fH/kqLSmKOZQQW42zBgOX8xe3K5Wl28oZELtsSO65pQDff2UteKv0BXuHeuZQ4KeyAinfmeH
rk5askl/jqVal8VwOaCgpYzmbqXAwUFcBZO6w/tfI3IEJPsrL+75Mjh5WWfGNWgE//5kb9m+Kngw
VPgdiTyB7K7ARVP1cvLeV/jb/O0LElHiWsi1+6Co9GzFQnT1cl3C7MzNxzBsBjzz/IW03EDn6Vpz
h85c/RcJsHYx13uUuT4to9FACkWSAChRmt7s0icxQjNLIp4SJG/gPVamIfH/s1mD0/9xWZ6ufCWr
SMNsjg8jr2BGVQyedGK0bg3+3i+RYDTmpbt5iwVHfPuLOgTi0XZC3k+NQVJzIQKVqf05Cf9eJG7x
mpT/7rCl4gP3aubF6EvkReiAxBkKTBa5GVz0wLjWcPPJ0BtGCLA/W3jM189cFx2rFaTN8nJmJIH4
vfHA1ohmf4evtppkdmVt4QcojHCVT2kax60ql/T+ZhlXLAnu+6/NoLji/Q+tQy/fzSGGvuPw3MzW
ou1lni50U8MoLJohF+CkmFDiaSTq7yd1ABjd8Vcc4i7kqJa5CWtxFLj6EYfhx/akzFttAgwAeViy
sGz5KoR4UIXV8EZ2WOX+HkYQgPmRFrEzGsgsuHMadpw46bYq9NXZuHMY+LdAjLsgL/73MDxudGUg
U+Hn3z7FUlyzQVpD/QIXC6l3KX+0py0fmD65HF3FrpUWn5vT/BNYKIiSLp96xW3+G9LvxccrzgRA
1t5Hr06odTN3rup6/9H4USgFJDmRTvN4QFTEOOU1IigBegAeW5q7CsTmcmabjj5tgIWHKgW73vGQ
msNRws2bGF+2kNvoYQDrfHj3MmtFU4ipX87KEO0w57qCFSThq9RCGc3IKcGyDNocsWVPWiRz8QMC
JIMlBTkHVjfFy8ncxrckiaZ+7RyPsX+refxd4nbVRYJTSdBJQKxnA7GWSkHuyLYOyrf48gQEpuTs
ev9UNlly6YxcBgSjuGtrzmaGcGf/MWdBwv+PRLNMSkohk96zD8rHcnbzyW/p4LQAwBrFoSrURwaa
MlL8aGwQDqGYLMLnMQjjS5Hi/Muqm+TtWCPPQV/YrwNyEM/OEe3GB7MryiuZNeDoeRqkoVEzIHb3
sLQkOjcTy4PgI5hA/WWYf/QW5es7eyZ0uSkSXnFNJIRpiMslwPEeAnGKXdipnp0mzkoD/VbOrTgP
R4oQIKvd02eR8eMy+vxEU2hfavnJB4lGASJdIc3EQAWjXtnHhNCTUg5zBKf75gyl3RxIkMx8rXkK
eHWyjisnscnATgS540WaLuMx8QIMkd2a2NnPVOgTM47y3s6dOBLxO5VnHwAVGoZWIK80OGnRIoJW
2vpb9D28F2G/Bz134rPItCII0Tmk0gxsvvbS9AG/TV+jybaejhbIrkixbZX1upsv6aSBHE7CZxxf
8G+tu7dCqFtNhEfuHcJT1GtkL8/7L7K1UEEGzn9X4i6wfrM2DKs/9eUYK0CwMVFKuDPjC7nTfotW
UZEJokZNMaOwjFXRjUlVWVHA+nFV2Fk5y5F5IJaHZALY09gN5PtuOrOPG/TuD7OwWFcEnQE8BMM9
A47/8lohKsc54bkZsGscDAKiZCYRVt2RKowWDb7+Ljv+8ZaW9hQTcpqFewU1a5enEeje+d4Qt+NX
sTbjzNm46ihMnbDn9sOxPsafFl6DnPU7eBSoPyl5AczVQqAmvIMd/qrER2C6Cog84LXqy3iHxNSb
yJfwZx4jnsO8T+A3H4H0zX5GqmSfg2ezYBny2naF+wd+ng57ytfygL6tDUtdn5gb/cfaTIfHYEUP
t0ee4f21Q/rpW0LIHRUQWTZFeLUNMo1/ymayCZLGZn7jZsFnFNGEcEVMhSqefz5T05UrvkutiWKM
sRovYwkTUn1jrbh9R0bhfdgpXXEg/ldgZ3v41NWCCgKqGSDXpN6NljqSnKDdcAXjQ46O2AHtaBLL
aF9xNb1Wl5nRzPIENHwXkHsBkeTKBLMEVKvuyck/E4qELR7ZwlKN/f0iN4sOn+6QCxtktcmmkOjN
8yHW9XD3dMSw2NW5XOVwhPkrqyg+NjKkiBPOnC5PP8wOt0NSTh0XTGf+ZFK3PMbibYCSL+JKIaYa
AqCHz4d7kNJatDStgYym8Cx2GwqCTCBB9LMp0GLzywpWgI07znHNpZ61bI1OCiPNmy3InCVWvXAh
2a81uJHP20RRzsGuZfo+J+GeoqrXBGnkzU9JhLB2b4niZYZVHT+SVPpevlYyR8O41WlYv4dMQrYe
SpVG7MYIGjYfnYqEJBns7uERO1hapF5jIWexJ4dcx1nNh6NdgZ3Bfdavl8v1Z3Zh8MbEn4iLbzR2
+1xT0uq0ryKIGA0+wk4xiE6F1Oe3wHCn1lEi/Vf4hPXzLKZwmY3UK9G9U+JbVVhGBuHr68ZxS4Cr
H2Z4zfc5o+D6cRV1B/rr/MLtJyNWgMavEloaY5pwMTsIG7BHGwhXs9NeUau58dS83rCvl7pUP+No
4KWcPsU1u4mEJCJ57fChIrBoSxDOGXGU99b9AUsDdwc7lrCWg3AKI6z9MmEFWMiFDSiRxOrTO+n3
HKdXtBA20nnhcgMkaA7TD0LbH/WQCuSmAfb2np0j2XY/HFv5xcUeM7iZdi/7nSoSH2T7OynUa9PV
6jCz9dfMg3DwR92db5PQtZbdvoRClyELDbw9Py9MAsJrYf6U6NRg7cQUPD4AUIAZFa97ML6czi25
HsRXFfxiShJQCkExaphiHXWheWRVwSOFUM2hGI21Jj0M9PB/rsPTIv1OJUNANCh5kSMPjWFnIGaH
C3N2jYt8f6UwhLFTlhoYj0MEzbBsjWZSRytManBxaHKP1vXKMOZlN3sdh8Jtn+KwSFXXk4cjXyn1
Cop47z2CtkHdNTdlCFoV75YXJvfFEu9tQAsOxR1vz3JKfY2Np+MCe5X5hN9DvqitEPXOXN1RPhJP
six+B09IqDZStNE/GyBZeE/Ld2CoRF7cTqxEM6OY7EBGWhbiaVwCDqZjiqDELCoEOFxcYmEk9Xkg
PTJsTXRI69bwoNwBJcssGW406JCOBHBo6HHOwZe9q+6LxcbrJYWsI8WBLHgOzlo0VCJfF8Xmk2/C
VXWfvd+m28B3ohjz5Z9e/8s5P9fT+IZgYRpf9QmKiXEZJa3KVCElrOGlt8BhM9ABtSs+ecldlXw6
uhkeHphayL4WG1zxLVLshy5y7oGNM0KnGBQDqzfF4hukeOEDKshkKGMxMcuw9j/rDghV+8pEtYX7
HzqbEPrS3Y00N6tY4Wb4ITYh3G+sx0dq9oZrBLbRkDln4KKKaWq37aJGVAnGer6fg9xgfG0fgjz3
XZr1gQte1CczlzdOl/H6kJJ6eSNshcCnlY1IGhWlucbJUItvrfN0VyKcJlETbsVwE3YoTTdMNw2P
vUKL4jsevCSNkacZyl8hxlWTKNvwzgPO3EV4k9Hvh+qqcNtjSAVGEKVvuxn6wEGiBSn2rlTPjZjL
TiN26WU8zG43z7imhp0FGB2bi34RlJHS171yXY2m7eN45gMlSV+2EcEThwkGtIjRiziX/NF131vu
48Tz+X/krQGRHRDKH4BiQbBA3xuab28DbWTpwBSqjEHk32cAtpCTn8snMhzDM8q3FDOlvYldZwVo
fFLxRIMQsWMyZ2vhQwU+LqO6XwlM9nbRelb0G+A9aJADCMM+56BaVoNsbgzf10ArGAS4j0KIHuSN
KYnPWI9wSO1dTgEds+DzUGGtKX9GRlHmvfMc1Ku+/pUVdpJgalq0KqaqRDyv/OMlSkew3FHo2PRy
Sm3AExidMthCQCZ75NEMCS+304T8Qs3GjfFHiAhWSqtHS1tNTUDiSwjzxU5jqwNTCjs/98SOY2Yx
ckaX7q6e/jV3EBKMtZGaBsgtntgdxOLYimfPO4/9R8YSYQ1eSsQh57bikneYRkLPTPW33l6WsHdV
MbD9NGIaIa226dXAe1iYCmGsG9XyQGr6st5H5ukWDMT5GFlqKhlWVxRN6rIfTApwmhw0Tbl2Az4G
v8B4KILaYWVzy24AkRfGE64wSqITVD3TglFE8CUIZ9B1jYRWizJR01WaTcojsMU70uN2JL29k1Hj
g6kkKr9tznWz7FYZvOVTCL3+OPkGD3uCUyYei8gGKVSFc+P4Z7twzXBe9/hXGyxdgRe30qnMZ/Fr
Tcq8PlNYwJDaQsNDksNI/XtjXqmS5zd/5Y7W/02E3o336JyBq5v9/G27Lf+G27JGGdavLpY7NWbK
6xrSGOyWoEnqTC0tIAhddG6Rb1pC15/5fFmK/DFd761dTrwDOFCvTB0VJGXgB0HBiUqmuxdhfw0F
OwP7qPO+S91b/0+SGVNuLfmtNdZa+ow39/aiMlkdUmOGBndhMHnRP6781j9p7avibd33t3o/Xidw
KmX0wFmFnPDGCoHh6z1+FPwEKUrhdu5c6FCtPjEmBgHX/kIVbhibWOdVvSpOHW0foIIkYSFQxpFp
SeL1Il27YdeARQcqVXrOI3D2F9seOxR616PP53UJd005CFRg6oeS8zSfnEIthFPqpJG7qskqRJx9
sBB6EMNrw8Tjkb/qejeKPVUnvanIGkz026hMuFfe1wSlDhYAkm4QmLzHNoEm1wTqj2hvdEjbk7Xv
bKllsULhQx5Z3EtTDZMnYHvWymjQMg7batpanL9Y3DN3ts+lXVQPFY3dMjZYYGIv6F/89N1AllCP
Z4hgoGz9+SOJfBoNv6A4D6ktJJ2LAUuOYZBvRJlTD2qIAM7/PmIqPvYjA9fUZ1zizQzlkCr3RhV3
pUGSWtq/DP/VX66xSHnP0o9TZqivCPGlWiE01uStqE/E52S+2o4/xWFSvHxQyu73pO0ZMo9mtsUc
yH8bR2D5BZjKfx/FgAgvTTw2R64Us5ZOuzmR8axZd04Uvp91O/T4sqDKd2OGRP21DBBn569yjvsN
PxEVwpK0zJ1fv227+Cr3dJBakUxQXMIOzdBccYDDPpz2+2AsK6s5S6agUKVllHBLDdrCwt0iYx+q
Zb1+Z2tF706VcM5H9NqopkSpH116F76e/WAckimLiD7GnoykmozGRq0VyD0Ida2Ve3uA2r++0gpd
HBTQbD22Kr/tlyMQa//J3mn1MGI1qEK4ycqcs4CuXzOFKDK6FLvIvha0/IPBumadDC6ZvT4FFe/3
tUhnRugZTpizjh3KHazzVDr19t3s2NB79jzx/zTodt+99BgSNVm7r5njA71IRmdUMIOgtPHShg70
XIdkKNKD3LENTttlFwQhQu31r5BlEDAAb74UnujVwSTI/JzfGDwsD8xbYN0guc/da7wbZ6DVuns/
XMTnQCyMKS5AxiuQdVRnBK27EwND2X0wQUTk4APjmOPTQV9bS1gZamH091igd8HTGEg8KSQ2/Nzi
/Pw23zXV0rv7tl4L93cEJMOBAtDLnOWManmnmTAJ3xSFLgGc/3d2EbYnpLJyKazuTYZ5cXxf/FYB
Yuvtj7UCXtThxNZT7HltmeCOlbBnIiJypDe+G5rSLl965A95KPjpgr0+0vIs4yjBbB1oa2HBST6x
7g7a6Ecg0pQsccvjtA9j8tHLmFOb3jF4Rlur2oO1w7vHSwE/SeuM9AdjhWWZDSCWmx+qHNTLrc/v
soozcpvv8Q8EpHX6awAb/V9gnU5ETuzZZjWyQjBWcDc5BH6eIpjd9IzT+Uocyz7CD41SbSy46G2f
YV6fpeiRNqeEWS3KAyRGaphtzoxrhW5A0ISMIEQ68jVTa2v8bjHR7TGGmrInWknJW2y2NQck5PW3
lVBjymkWtSiRLrifIk/SFVpNHnRmKQSe9LggK/lkgD61AH65sOEtjwCPrk1enrbHTACF1ziOqyA5
cuHPxR2XMPP/a3gr5ukese/+TfVQN5iPjmpXs7VL3ZpnKr2oPwGtuuRMZXUd+vQYDlaP/4ToZs+5
/vLNVpTyvRO2K0Tuu/nn3lT1OIqzBDfghM3pTbL+QHLKNps5AMuz4cEO/OxouG0u5SM7CZUviaOr
5733WGjB44zZ+kwN4Qfa0+wygmoee8YoGfFQpCRM+f11YbUPinZF91Ev11b3rENihYpkzqVCSMs2
Tz2shAe2bp5Wr072VxxXgP6IJxBGIsk2yH3irETUysNjpAevv24KbVUlVQv70d14vb1ld/fyx09b
0+65TbHO8qZB+gHhcZP+CzfvccdURj+WWOVKnlHc9vyEA9A5iWRHiBhxWDW0U3boKtzU1gyoypnc
UAJ7eVa+M5a4r7JvKB0DEg/yPprCrKV5fek09sHavmFz9y0nAPZm6FH4XJeVzaEEJXS9uaSXSnSq
Mbr075R6O4GxE2suLzVM1h13j44ZqSz3KS08ObZW5aEgZS7P0pHQZ7Y+4KlLHnbfQQ4oNqs9J7JO
JsDHQZVAaqvaeddnJ7KLWiE2PuxFXXU4ELdp93Ore29HGeEMVF+Mz5Pz6ulWPnH2wx85143BVare
+Y/1YbRgKXJl5jSpSqIeDnIx5rpjolDsMHVdg1LgXyynqa38eDSEnSLTGXSMNZzAnbvSwvNE/+ZL
XRh35d7dLlnfP6R539D+cNt17KM0dXmAhn9/DOaUovwWOCREfwPCN9Cf24jAzoHGFS1RcWeJ1nTZ
QONXwmnXy01GB2g2iN4aiV947QKJBZ8PbVXRrucPuGMb8V2OmO6djt4b3run2uRh44IO7IV1JqW+
JotkpCYg/3URIpn5X77N+0vxYf7GkZmaOl2OwUN5F3tNRDKXaulv5jG5jCYY104R4VMLFaRew6Yh
V6yavtxJcF6t66GwJ6qHCLgjNPFddlQdu+zQX9UHxGWUEBvwV7lNG8Y89J40Ewbd8JLa9nNTg9s0
kXD2Enu1pebJtR41vhcblA8aon+R83gR0D8JrT9Eb1KUXM8ehOk4fhUImRER4DBSO57WxchOYi5w
3YSKgm/piegS+1oUpCiEvt0Cr0XkRTWZZAVhKTn7hLAu7+f9qkQVvCEMisLvtL5UPLNLT/WFEm+Z
1w5rvIWqEQL6oUggV6w4wD+J75AFRCwtuTc2BBkUQkO8hF8mcGiXHbCaeDOTfUGX5YQfB+y+/vmQ
Q7nERhNxf0sPur0IKUTDHEpqbb4LINvSZqtsq/CN4DNdC/6ioI+ooFOOevMRCErTTeGOtac+/3tj
+8XKUBufomXzMVh6UWS52d6dYh637n3L1W1qshawVWtvAvE25aOfcQcUX8CHGQ/1wbMjVtHlfzib
ADQ19UzlifGQKQd2qpZ2rtDA7vfk7cP5NGuUj6Ewmj2fJWtNPJostyWdcusmL1BFNlz+SaI/k19J
20JXYx3rtqzoyX9xGqCK7wV9h2PkLCmvryyAuNQ3t3RqJeOaGNTkaTWYa2KcdcrcuWXNAKfdQAXE
tuYYIRMqK60pBpX7x97ymoZzx82/Cj0rXoyzRcVj3Fkubsh1c0RkdeMqaqtfiZ0IlaQHzR67ilhq
lu4owHz1ZCStr3Mzg+oRqi+sJn15NDskn9W/QPs82MruN5CRAmE8piHJMMRC+EVWtclwIi7Ud37L
wZquyb5lw42tR2duJ0sSSoC2nxaForZeWrIX5oy5sd1+f+Vlb35w6/x5aqnfjmskj9YC0sh7KGpJ
TG6pr/bqmpyF3yRc1XfsG6a3Mw48moqNbXw1dOCYIZHyaU2EFydSc43dgmuMyRrIhElbkQotrAEj
stVFq+iKO5mJA8d64GEH3RABkG2wUkCOHifhAS0GET3GxeSs/D/WhJoX9hdWQ7p6fVeOKAcn52Gk
6eZgizsdTyoWeNZa0cpgQDNtBb6amQ+na5lXwpcqmwXhJQJR/7MQZGNItPKhSoBF/ecfCrZWnbXV
P3atXG4hijajOH40OsdwMzi4x13lsetml07KFnHQiekDtB6AzFH6aGroP3cAs2y068QjXawAzGcN
qLXOSQqm0c/60pArx54XMrybX/zQrYRNtpgKhbiie5Ws01CCV7mD6BeatCAmYKJOeVOdSlFcOrSf
xGpQCG0j8PBH+MQ658n9gFytP4fqPyxjpJhzbonoBvisfBmlakZZ5Ozlm53rTH1n08KGvANcrSLM
ux56JNqfNKqcy1tqtRU0R2gEJSdJsqwm5o8bj02M2n1qr9uSYNu/5ErmS59MBFhA5lAM6/ci495D
8ZOfgkAZFmTlXAmTWu6KTUN0dT76gWWuKMz4sEZRYMOdjUmajWxKirf0K2uzs7dPTEDOdgH2+OXK
+UCiPjPWMtUxLwmC5La99IHDeaNTaRtwiNjqSUj1qVTHGoWE9mQn6uJgKF+SuKolS7FQYAgAJZF0
Nu8nXvwnxJNUrYmaIYhRPDtfTo67phoFInJjquMGOLmLQJ/v3T7ev7b0kB7iesX1ZORflyeMGAk/
N34YFKFJFpx/e1ftEjy3dFur7lpSZGAEswk1Kz/QLAzk4UtN76kK8FP9xh6BUKomLKyHgRgf6W+Z
ScufKin3nzsgXB3ScuhMiXCSLAdA/G9qJn95r/0t3+urpc8vZPiI0Hg0hPfh4nCauPVSsh1dmpca
EDaBKWi+1plFLySPdztij7CnBTh9gmk6KwYV3FRXGVwiiZ6oA5thaleLqRVFQpRu1cH3lhmwVRaP
8hW3jAS5ItLpsRlS8GJ7WTR3bZDX5RkOJvfnOAtr8nmUcFSatnpKNPJTcUCi5T5dDdai8qIK6Ecn
nrGZtUgbcbaM3TjGXrOs3Njq51W5vZBQx2vlyp7AVJ3Da8EmqyC/1DJw5F/HJztb0Dxa9PYHBecU
bXepnvbFz6vNvFCuR+Uca2Hkzxkpp1U7o54fP+XotD3BIhsLZZUrojwqfw434mJN6TdvxbGLE2fp
YDo4iRNNe4vsFgyUuTKDzImOCpb2ronk+vbcQ5Qqdihci/tuIqOLjxBnUJQ2A5eBztLPY2ALiq9L
XOcXcT53MMeF7XKqeExgRYdtnaEpzfb/f3bWq1L4+/xWH0Pc0jqVHFWgfWJdrt5fQDho8tA1Y/Oc
jOvo49tAjjpkp4FN4cs0gPxxjo7G74joHrlPZdeQv9Hfas2eKWY4WDOJvJ49jrLzC9zmo/Ldo+0R
CnccNQfxCEgavsw5XTrrnSObPnxzSbEZI5oztptXiwvHYSpK8VfQAGrPY+qodzMTrbxa9lEpGnfl
V+Ug4Mx8vz3AYP7RtweP8fZjR2SUbWaAoLN+ebN5oSc8ViDQmezw1Kse8Q6CLG1ujx46V/Owxy2v
cEB3+DCUhbMqhn6LtP8U3PSx/Yim88hiVLI6i5rbRdlR14LQ1MOwMoPcLfpCVoOXErxGisyB4c8y
EjMPvfBjQSR6BKTiCNiYV4qJ8J1B8bDBYZXPXuKj/y1SNtr268rC5jV+A//M3KnhT5xiVXXSxRSc
P7qe1AlBJmAwww1rb2V8lD6EP7UEWJFkjNlnI0UKY4W0+MYBWSoTwbqBUeiw2jZDIeQmqEIsaj+d
cZgDMC6fYILDT9RLll9ioJKwx7/HvH1Nny3/LS40T0x2WolE8zQ1jK4Vhk6+9LMtWpNjDp5yDEPb
JoLeUQjlM+2eur47pTWcnsBpU5MoUntF8uNg+oxJz4ocgPWfAHqvYJ6VylgRKebDMhSkhwsC9XGX
mhnZa47m9S92G9nQnON4Mrl26fAEKkz3BmfbVvXwXm7IEsp28nijXroHLadBlTUshxoldSbAGkxq
ansHyOoDzwVBUo5W3Au1xLJBr6cRQKqet1KpxeYA/KVazPnaAYdpmnECyK5BBx12I5KE2QcZbzNR
ETUXkcNNYWOljnjHN2Neo70pmOp8wP5BTSXsJdCvXNnxBeeMwl0lj1iq0QDRNzwcr7kw0MbXmPDT
Zj5b4trvtJOV7l/tuBJeyAOxpqXTdy3z2wknsNDwVbiomC5x0x5B/U71YlnTvWA91chGNfGV7oHe
soDt5LgC1+6NmsSPsybmdFSFyhO6FEl8PaCUdI0BKmm1JuD7YHeEdh1s3hqxgzJp3xa8DQZZreN/
P4mp3MHzcIHMoMEov3RSoFw89RX8j6COg8KEYARlhRe8gufVfpJFgYq4GZbQ00DH5QSl3W2oyzbe
pYEma7YCjBwAE2Eq7z4yCoLKxPULnCrvB/pJAcDpnRu6km3+y7ImXpggARhfDmgImjaJoYDgZo+x
YJf/JG1r9Zr5RRLr1Rwvu0CEWwUz1vswTetB/0Gf40KQ/5PG0xnHSsx0l7sR6RXcBQ5+hFU3+90v
OhR1DlrjVjdg/XvXII0WUH2LYsgGVsWQtPvBr7I8C1xkEshE6Kx8ZcTEJaw3IUxEln5MOcMHe3KB
SL66RrJqWSjFvPGLGiHlKRs4c3VDvTmqInp5KGv5pZMCdPRPWqaX3qcqt4igg1L8/TEXVjrD4VKR
d9oH5KhKQn+YGpd30RTa02l6R+V8GhK6CjsKmYwbdWRVbUloouxCnjEpRHHYbxTTyS27tLHgNGTJ
FV8zJvTB7khH7XeotLKzIcrIEG7YjcXWvhEmJnwl4Ggz7zE24IZSSQjiNGSkJzU3N2f9Lm3emNZG
4iwU5YY66lSHFMJyQFzjre7jat34kGOX6m/4fF5wlXvFXIa1BT2XXzaEyeOS1i1JK+D8YZFvpJGA
x26p0DqlK3Zq37Epy+NdVAKl981FzMyhCcHgBA++vuiLc5rq9Wn7bhnNy8ljCFBWKi+FD2VZWdJ8
ckVgRV1aP9UUqVB5l/eLP5gbZhMyA2godo7hKagxuq814CQAk3NMWtIFppCosHnuzTxFGoXpt9mo
sxbVwIO9Fa/+0AYljQqCLUcQafB0eIhGdohsdNW9nnb1iF4TPZKYuKQWqoxA4SCZphQKomXQ5S83
zS6MDQ6To01aplR6Cn7YgRGmAkdWnkhUJju5Da1YZOV5lrTMYvRm1UhhB3CqNJCuvi6bsdWaWz59
OHYRqNYJszygp+pva6SvV8j6VVDr1H9lnDCucxFMgUpN03DbIBdIjbVMXz+9QXGo4PEWcQmGVWC4
ixEsyHquFzb/E5htqDFStup5ygiP/U0RZ0fH3fHr484KW8yiB8CLiXojYE1Tfl3HOr7j4/ASmM8b
Q6tr9hjNO+f5sU3zEXgAOdHdOrGvy191lasSSsSydXqxZww3GSxpJRP5YUWbe7eSnjcX/EhqPoR8
JtGF52YbwfwNVb5FpP0S9/2OyES/tIfI75fDLl08G7Hdfz5CJcDiYYIxvdWzMQmIksdNYJSA6eXn
ejeTejlcMH+HkCKbk7UBCgbl/R1pgmsPmSJcy3c+G+SKM2uxjHbdKJlU3Gu6XcstY4CQFvsHzejV
iyK8sLqvyoJM+zY49LLqtzDaDlyeDT0p3R5aSbZqPgODkTK0CnKVvIFqrQgFXvZY9XxAA0m/jmFo
uK+l9d2BAoaTBdWOceqVMqCE9btLp3pDYweJ8g9VXm2F+UtYAPvMLn5rpdlilLhQSHaCpye3qSk2
N7iQwGh3HKj19USG4xJhfuogRA6OTOD1WQ4YK4dWeb9NZil6jjMwQFhgxuPrf4HiZp8dq+05DwWe
orpeVzS17QrgHEvsEg2rzT+BG7SjZVrKRtgEcmlACCUxp6tNRlI5o4ysXKz/mfALhxF1PK5hCoL2
z8BtXFTP3EK7kX2bi0mr0p0ZLxcgJWbmFofvTu4ymbmYTDUOxkWp0+Z7vBGycwrrOc5B6UNhYBSs
7LUBOLnIYEzjHUzUJnnjkrnqk1JMLBM2eOO5J8BDIsWoqlgyTE/puZED8+VE8/tensjNebSwJfUD
62smz7vRXZMnxI24AWRdpiv5A8V3cSoPbQDSpo11YtNpoy4qluSjh3fq7LCvGexESrWwhUacpXqH
6lz6d6yLb7f3MPf+bUmJBHAob2oHitdnJd+pdKJIB7kTh93NYUpQo+JDszhuQuSDNqnLc9PjoU4/
wD2RVz4X+RVHbcHFu2o785TqMzvabLDtvOKoNP+2PcgEU52rrRFdQZpfmS3ZI+LlN1H3T/5Kncde
sio7cbqfURCG2WwV0CG7ZqGfJQVetMHAsmOm/ut3vUbuM8SdnLoCwYBoBuy3btV0NiR51r5Pc1fn
NqlrtPMZeU6sqjLjCsRdd/El3Xg4UKaqC4X84aBDiywKnIJmd6WhKU94TpVx1S054IdFfNXEPq5X
8d1/U6En94t2VRMRlrffrF6slpePuE4ZqYk+92v4nOpi45U47S5t6asVziRGTfp2SLN69RTAxGwJ
kj8vXt28POXAo0GhIugOK+2d7V0Axj2klPIipR7j6lFVVtmUREBTtw5q4G7q/fJ1Tzb6LEQIvP7H
2bdNuLeqL9PkKXjn0s12cQQvifeUETFXJUNy21AyD7cqjf+3PAyBRrGRAkDbPvYatZAjm/kAffzU
atp5nfjoJ3DCAt7McXIHsizTEPg2/qB35tgfSfCAV//3opk6DgpjbZe8zpXJnKNtGrwL5Fc5SZhI
qyeX5lJty4VFOuk44hNyDbByXP/FEGkksgtdtmOko5JbYIC4/g97QMlHPdYZF+5Xd0uhTeOa3vhm
8VNmqQV8rbpKtxBrVLCi+vVmHC4S2jF45rFrOmfRcJP/zcX6FRiSsuHSaNMioTZ1ocMXHF14KZ6c
H5Mg5xFZ8T++UTL52+QNpSZfp91mzSiocM0N0+zvENWzTAntSXPsoleKkyBE9DAujsfpUB80tKNe
Lt+oRgyBWFtdGoQQl9Zu8CPdurmAMBcxupMgkEJp0LwNZItC2/gRfttJdJH6fOUpeic+R0WvbrN8
KeZUwM661BGizsETLft35xNdZBjY3JxYrZVcwmaZKk070PtC5Bnvco0Jrl26ImacfAaA47GQ2OzT
4yzZ3u/WAQtKjYZju2D/LIE+k1yQmXAVbr3ByBkdR5sOLxSw+NN6coWR5juuJ+JFDqNqN6dA/fen
WXLhrix6tQjjN8Sx2vx/cOM74efkYy2MDA+EdhaW4pTD5Wug2xynDLUkGh286lDXYPhoYUY3+3At
W3CzJKLdU/Wouvnw2JeYUhhxgsXfnzg+90JGvHcKWgfwr1tRbmAKIg200O6zXvx2gO+nGsOtREXf
aoTmDqJreN9PqdQ8eV+ZvIQS6bGxyeg5OHnwYtv83jkcbmitmmxXd5rAk0f7evYBdv2C7nXH8Pdu
k/QbbnH5Vn4txddgnLSZ5ULO7zSjJMyc522izFWTP6qQnUZIfB5Af6gK8p0RxLLjNnXkHo6WsF4z
1KNFxX/dCv2k78JV3KqBmqbtjn4+ehfhC6gTyZNBfaFE5AcqAMiw9O305gOJkxOtgrGdmIioPIV8
8pIGf5+0r120NilED1Fpk1F1lzy8EKAURe5ULzyCqcA1RJYtJdFseHv101rJJTI8fhs44nuJNmoL
xUOfpDXpjCcdxI2qJ+CfmvuGodwini6mia8DeKyle4QIqmR5RZ2gdOVM6V3XqXc3Vk2BE70Ndvpy
QpdILMaM2ThVj1qWoa6UBRKYnaBTeRiwmEWKe4aCI/M6aA156Debep+vA7OCiP6XMrXH2431eMD2
D/EY2QhFkIJsEtTooWqnQT1Mt3RDaLeJ8nAIK5ud4DQwnazFOXVuQn3HmRdLuGTQiY+cFpij3nmo
9eLxN1KPSdq7q8fMSkOOTBxeDeaIw+3A/ZsyAu3SulGROrUhT8rp23GiHLg0zgfu+bKP4Kld/DIV
i7o1iEXnuy5nVFlV1TfADXYTcq9UOvcixfXf6oHlp3uVAw2CUmaUjgY6z7DBvVePiuFBOYCTfvu2
V1CmJcaU69cgH5wrVoZwSJN5Oq93m7wFmzTZspjHPvkaA4dfgVqIIcfHiJgr/C8Ukd5sEh/0c6iG
f/A3JsqnK8slWfmXsOEfQNYeeyVOKCQMxXvaH/MskADbZFt624Hc4RdlMsmMoQ7RYn0PJe8loyoA
tfsugT/HigWPibgR8u6+AmqwNJ9GBcUHiFSRlGdCQu4CppmJ0uhoSWghZ7lthsDiOkWi6sCx4w0w
0bawFKQ/t2bKoXnkax4AvOWkGfH+PdX5vIoGvs3T6G3DzA0Wn612ysmkS9P1z4OrmuUtujP7ki6V
JigCvRLfYZ2LLDe04BkPAOymaLcrQx/fXmQ/iaA5W/7j6Geax+DPSKVJXgaWPhk5leP4vB+eUq0i
Oj6lkP+A8s/Fx62aGqqf93BLs4QujkWvPSSyrmiSv1Qg/32isXBvlwi+AvoVCGS8GSk5TI5RXdkS
PZ0Wgd50UCZBy9MVJuVBOQm6eJ4PjLFSdROup9Tv7U2EdKy0pHxvKTRBF1f2ozClpXsetbbI22sl
VhwObsBL+sRm0hxrhKAbu/dNRQrjQ0U9GRmmovnFGSwQhkVdJV+Rw8F0LLjTdEwCD7q6Fs8wtidh
BukpVqfbJJGCdvzcSq7NKzUg99LzFfzRe+tVXyMJwWB3po/AdfDwYy2GzXeIa7b9ytJAcq2U4t85
kVLa5h9tDacKND6naO/sbIhuwysUu/fFyP+pBh3ed9De2kAo/4GyDj0v6wtEH/S+Nd52DDos06lD
2WnVJembBgpn9v+30RZG4DKkQyM7aUHVzv9bADdkFNg176BJYIaRlO7jSC5p1d2PWrO1RWyzqRcu
6gbpR8qQxWFJh+XnzPTN6vepuWFbSymJAjF54nUdpoEwstRMozzgosDlYjS7fU9VElON1VhxemW6
sjQ7KC5nALivOdfMfAAThReTrCrurzYe/+SxFPAWCWQgD/5DkV/GUCKJ/1SaOP67i3JX4S2J37mM
Lqi8uyUbeOpPBSeD1Hz8Mtu3xjtBSesJ7vuPpx9KBnkqaNUyIgXnYahoM+SCf4SEmsA7E6lqgIgl
rsjs0rLtRfEJ6z4rBz/6Lj0+Ya/TI/a4/tZXe2rpqbmJ+QLsExefmuMxP5xKMmEEP93bUFVDvg6k
9qbP2w6b2HQqYCT94tLVmfJhw4co1zbuyAi5HUml5r9R058Ynj2IozqWAkfZjtyZ33/JdgxxAjWD
jG6PPJ/KlVIErNcY1n67UizL9EW8BwDd5ZEAspncH0wwLphAFG01RYoAfFEGuJscw1MTPF6+Zv9u
+U4bq93EzbGvM5dBfOGhorjVDOIqyciKqsYp3n2XSfJIpV4vx3HwqIgI4eKdy8mQ+dcOIVqCyH3r
9j19o+mTamWNhYPBDkmmUJ+kjHZNtSKaiNtWf+k9PvW/vtPq5ZZgxMCxRRuw5rgjdMSUlNCUmcg7
OuNbmjLjqgc8kT+xGbWqc4j5vFf56/CCSFFWNr7U8HGZrej3SDRE/4uimVY4Q3CX/yG5mOSlWMQ5
CD4W2wrLzx1/DFocrVVDTDn4aX5UrzpgzLx42O34CggSE7rBNYQV1kFa4Q6jnycxnUviz/FBvA4Y
a6VaOm26VF2M9qLJvk+wVH/aanlW31CECOkeCPmXi2u6/MrQnA7aaxm0ckjsYqFZMBdiDd5NvHux
dLmg61Q6pSOc1RrX9mt65cofrIFRoZAG2criYFdlAOWVkkvjmXUCmVniIAMq4h7lBzozETrbC2to
8zgGeTvX5+RsDWz5xLWP9C4XiG2hOW9uAvoRFzXlL3wkrFxBOfWc0Jx7H5oWMySnEgaY+rpLGGQy
B/Rj1lcFoWASNemAlAs+POsV2Nbo4bYD3oVKaFINLJXYH7CBYiviPPUbAgIwhftH1CJRGoLAIvE1
wndlA2NvsAa55KA+2JTm0MgvR4I/WMgOkzfwVHvcfqv2sgzz75646a6KrCtJC+NhzwdVkkFnDM2R
yfofqJPZz4w5N2InFvJ0OH7WTn10vDFvNeDcxazBQUW2fFh3i2thTGgg0MAITY99T7L+pjEfAZXv
R3E8BGu6A0hiE1FKA4sFLMyNnrwbNbmfZqpKVURdg8bLJ7aKG6IbItmjbl77dHebr2kOMNt0Qcij
pnvp744czeTN/dA8k1ZC6O9TYGUGOh3HUeVIh7y51PwJvXzX+VN+3pwK8RJdUFXhhotHpld8aOcK
CNAGVCyL/OlrSUNGWzldKnZ6i6fZPf3dbofzSjyuDCLSGRJCWrNuSvJslLPMCmfsNRmN1uaadska
vxff+/K/D8ZG/I4BvdKteenOfgYFEBMGSWWxQfsD1X2pPD5pADk+9D/LTycIPNIWs9rnj2MOBsf0
JiZDV3uy8IUV4B8CF8D3mER0RQlmEiCy31hpCUz+dWz58LiBzbvMT+6m9OxZA+HOCBhHU46+TsS0
GZ5S6oL6VML++Q4N3B/Ybpq9GH1IesPYlcVV74nRG1c0NbfalsKjP6c5NR9NE38uxKRqwkzgCHRg
9pYlNY+AXykK9Git7RN+NDMSTMv7lTafmCLiFN++hF3DDxMEm/Ag4+oGJbyZb87HNXZ/8QIw8lH6
S6uq8km+NLIoNdRBvQV8wnOpU/uBPmL2GdPQM/PZLo5myp0CC35O4VpsYvRyrJIyUOH2Foxe9jyn
TFy0vVmW+K8CBpbeSNhpWCg/dt9po/BMRvnZUpKaezLem78j7Ut7/GC71EuFcA9t5IYhsfQ6QIrj
QqhtLrC6mvyAGr23wyZT+Zkhgu9mWKjjFimCpZits+HYSpk/wuaCt9MMaFxjpV8vv/DLQxne0ZBn
kVtBcC6OjiILxiYgG+ppKvZkA+jZXYguJ1e3IB/0OVnPOpBiobzLXNQd8W7kghS/FQhfbJF1ynlZ
uhFLgQUCAqgimPG1ptUBi3JqeksaoT7mPtj53UbfFyAlccpdci7gIN+Laahy5JmmYJpp7GHnRwDc
tr6vbEPh97HWW3p2Qq2Tq8AyrK4w0viRr2giQNThKPBYLtfdMwIwG/ncccR6k78DIw+O7jeW4aKx
LzDj1pDLBEqFTgqd/XdKTyeO/WmfqqFH/JpMftrWTKcJu9hrvQPWhQYbut+YV26DhMUAKttbVQZT
q5PN+z2PkL6EcwQrAOewN7sDr2UDMiS0ju4Y3v0eiyYar9JfaYI0i3EWeZZ2kSuQh9M2POarbQXl
hq+S4FMYG2/I+BkZCltPormq9U/yyaaulXD5k2XktOIyTMqJbUCcO7fRpTK5/nWRtsqiNkyOH3Ru
G6aK1F1BuSxGC4IEKVSsQkMMBI+tBVzTx4S6YdDEWBLZLQt7d3ZVgiyAoxUU4Fp98cRpWHAGJbrZ
ek1KZPHYK9yOHpT96Jc7s6i77l+Iji9IWN1lTLmaULs8ChNlMJKtQebqpGEdIrmjYRybEZyYwQh9
5osShYo1Bp/6aY2Ptk8NCHIyEbucXXgF/xX0F497z+jkZXnaRBn09LOIXedGcKZposCYO44+k1OI
oiHfFIaHyrjK/xz3plPaFlei7WbhXsE7IJRAmpdUSfn82E7RXKq/uQl53YbKZ9tnbuPhI0O2lMoQ
6FTSMaujRy9wvUfNt6CTmud4XgDXRqtFX5UAaakF2iuRR1wtQj2SPLgMuf+yMRdgKjQeYva+2bv8
oEDF1hTWWJyCSbZbieGF32PkNfJPnzSsCUrt0vMuD0KdVwqwqzlgT7W4XOdBcce/EnBdYpN0ui0W
Jyt2JTO6EmIq486WCj1u9Io91j+7bJQrTziqDw5f10ZXKDvO5vfBLEWFmB0+zNAuwnd0VutHOS3O
uZ1pLC7xi+vaVAfuOK6VHxXrj44bURCbbDz+AQXvHTd48T1u6GdCaRhdYem3CtOv0jovkw3XlU/Q
/1qCqaopo9j3q+rcJdNzVRXFxsuBvKujDtPp9GdUi2blfy5vJDarSjtX2NRAgOfKRqXlweO0SK6p
6r0RWX5Ps62OxQV4NGKtyvbKYxn4WPb/4VTPbB/7oBLHBkBcqX2ZF20J5tNUYtDCDFi/KjiWZE+H
nxmel9m4PpITlTRu3KWeXbCKbK1Yuj7wTfjYRQFCokfIB/GgN8PfKc8QIPnCttphrOYbvPlaOs7k
GL7YlRR5NGQiJrFzjKQVUsYeIdC9UxtmlA+3EgFiowNSQV0qFGW4SfZ0ekkkr0B9MUxO6dLs4jI2
U4OwNZxwZYgClrBpiwIPzc5//3vgrxIoMEK8HirVvFoV4TKTsA3tHnuqOg+nUqjrGq72/FhOq5Z1
SgZAoQgkC8hfKPVKR5HF2aaEEPCvKeLkctEJ1tj9YsWPp0B19lBc//22tqPJn3/xDdggOBHdQsWT
6BdQhbRvbilWdGTLOZXS66s26e3f5QpLhKg/2gZBXZsjTfY4NibPKrJSXoId/RupqpifCwOPpTZR
+IaMt/567ilWt95ZGqTf4KxhUplAD51WZPngM7sPVmR7wbqDKxh1lAjqJmHoYrDnKiELDwos839I
VML8/vF2agq1Uk0LjErRaPFL3f+yCmhrh+We4m+zoC7B/ygc7eM4UCsbnXvvBYcKLc+MtO0gI66q
Czcu5ODm3PaEMvDFQtpWXBX2EjAC1Divsia41/i+TwD31c8nhsjkjpnSFrFXPiGu+5sYR5+pgxBW
orjUigwaeSBE6PuZZdTNMP4cvRPBh23VtUQQcBwPmBofx2xwOx+SfVI7M41KPxBUyhupnafkp67O
EKHDSVMbljqewXFQ6kzM8+VqBk9H8wJLM/jXrzji/7QyTMSojoIuX9NhgyJO/lA9EZLuaHkeL0/w
ivkrVxEKHx4z/tT0kTj/6dI0lvuqSl5qbOTBFOiCqOgBQYDPiGX9Go9Kt4Exoj8eBfk4c9zrSt5Z
Bsj0Q2JdS1Y1Hl4OsDyqpNYrCHjzQWQyj5CPs9+vL9SZoBt+Wga1NZYT8v5pABHR+Vh++j9ZVzV+
MONdT8D0HUcGpS0vz1iqkOaVBRWGcoKjKQiF0XTS7T+jYHrli2YD31gZjIxuIj32w93ZVWUFoEiR
OBQysveyoM1ubR2rTK72j0gOgPFwXC0JeZt/bVGs5hPh4e7z01NgT2nlVJMLvqM1ya95ZsOor28m
iXCEMdlTJlA3M8pwVOsQ17rNhqdNPAe1QN7Fk9463WkkYs7CMNKyh7ZolkszIl3+4BXgGH0u9vVW
KRhAD3JF8nzsG4wbdEH+24PFLMKVT+3QhAskMuJq9ieWpdbc8IYjYnwRbXBUfVJe8p8JffvoJhAu
9hB7IBPKQKz9T6s4obhYuBdhyTeWClPsXN5SwoOa4tS5dejDgEuOrnKEeOVbQ1iaDCKlN1yyHz1s
fyN/iSZFmOvi4wAuhZ0ow7x5V7b2himc2lPem+TKIVaGj4QVCpejSPkii90/FihS6A99P72zaV+y
Ngw/FxW/yncEo/9P9aBVc9LrGPMXoIZY2TpusatRKjVeCHhCQ1pM3kcv2FqK6/3rZ1Har3GA8BDM
YWEwn+z0IHnNdjaabAC5YrLo3ld6dFY54w8PHG1r0kLjpyR5uBtY8e0NLtgXGl18YItmgLFpOowI
DQsK7Hbm6Aivg01ZseRVEJP7DTm0YRFYJ0EVdBz0HnljI/tVZNB8YesYu1AImbxR02BLQhxLl0q5
PGhBztoZsA8zGq0Mtu1wi76kTy4NmJ/S5MEfj/6k8d5/oime3wUItLylLDwQ/6u89ACHX+KSZEIs
rcco1KJiL6g5QzbMsnXC8nutFywLtHZkkC+exSaM+WfMdbY8Z9paI0pImWp14Mowlux/+iHwCgjI
kgwGhv99HzKuRPmSH52okMZ4VTvf88M5GGmmAsrRZRQhzNe887DztaT1YWkr22fhx7hOlbu0hmgO
twqeOf3iO6dPqiUafZaFiFHSQcAxIFne/KU2t1CfZ3ZIns6+vBupu4/5wurQlrU1TXntKxCeF/AG
5oovVszSI11YE8aS3Qb9n0XfxHyX+XR3SOvX5JakdsmMDNqHWcH2jA7q32xX51o6JtXTSkztYNsc
oIn4s99B6mW6e1hCPBGxdQ6m1bGCjeuiLktIiPjZwRRCztDYz8NlDKQZwJxuY2e2tgU8X8szajuP
QcdH+DAAhgpfgcs70fDgzXWfZ3sKGhRXFPJTgcWjlZXov04P+9qSxD6AF6TmcOQfa8luHCLBSbwU
GDBhC8LE97pm074EZN7oMWHhqcbXl8zU7jB9qTQShDuFKwnaFAKOO7pEz6EtTAZOpb6Z9G77KUix
62dFLkmZUWgnXvLAOiq67zquy1ytzzMmzbHX2r8Yus69IwW54EFXMuOdYJf3/Tu1ge8+wNokPJnP
YVANu08q2qSxLxbvAxTTWWK8f/mjNWye778mH8VBPH4M5zOtMbwrlQXjUx3uZaVLvY8/8uo9HIf+
vc4KooyF4oG0GOsf9kIL7aruP0V2wRUOh22IxP33IWVId9Ud8u9DOfswSeWPgA8rd4ju37HUD7CO
wDUCnbHLrl0kDASDi2vj7wdFkrLmoku7XRuYljLkOVLVmpLDpUyZJLlGXQx05Wq8Ymsv7Ai4ZfBE
Cqha09/1cEeYLFx+YQ3Gbchz2SqbMJadpTqm1m23vz0M2/H1t/AO/bm8cg6nZuO/cXbVS3tpa+mO
WmpLI0E1es9HzEaRHhDKVTTmg2+kr6CrVjG7UPEmmXKMtj1BaMCJQxAUCxk1Qmy5YvrIdlkZSDWg
+/N6ltblSSQYRmOI91rWAoQi+obXDMRdUz3Km8VexESzYDdu4z95Rx4HfFXXsanqDeLYHL1L65Tv
y+fmQS4CEBNxyJ4BYHACp7usOnjRuHqzyjjLWo9XQC5+9FSbIHDRUtkD4Gw+atWL6n8fgU3DKZtA
qffqoLclQ6bgykrtsFrDQicshLka49gt8by0TWmFMAKYqfsCzxWHiFdmNYV57s6obDhILR25PDrn
Yipb70xUJ9ubOgNTq9ly0bIlD6gHZjd5yZJkk0HIpAO04FRZqM+bSTvVrVvhtLSEF2VTJB/vwVcY
QJ47YGIy2hHDTWZokG9M/rWj9byrZs6cD8dyrQH2SQM9KRu/JpLLbLVWUOs0bLUOY/iLd7fzBxPy
7K3rsMBUauD66OoTD5EiJsUeCn4EDb8LPQuLPuoMgiZIPAGwr/kB11CJ8bocrZdNL84Qnn6j39aG
qydpRQhUuTeGQhXK2B1SYNbpoYKSJJz9uVOfYS40SsMF7p4MLlCEsvXsktj/nX/y9x0rSPBlWrr7
Z4n8Nxui7RJbpUDfyOS94ts7qxLNIH1O1kmFNZDvcGZnaSjc1jxH2LG4coRWfvpE4EzzIMZXrhax
FZ3IQKgnLE5vatMG0j8FkFiQlAfD4461cFUWvfmF1CEvMKZlt5FESCp/cgfomdVY7OLptvFmjuv2
7go90nmFHN8QDwKU0aEKpkPAwusEkxiqfobh7447Xj+nnVfwzehaar5vVY6Sul8WgMad29VcHM2z
BYU8nNgqcyoYJN0q6giLQZj3JM7q0T9DJSBmRYzvKyj3vWF6HcCiCjz4qly6MOGrtyW/mICyPSP0
Zq/snik7sJvjGLfEi244SwneAv2swo11qxn2r8+/nKlJsNkSsfoCPwGFgXmtIo/ijl3qCcYvCvAA
FOLrOcgZX3Us1vp5AnIswvldsbc+7E158W/QpgbWL62mdcDGUoeRvU476YAuNOUCooF8o2FuIgjw
2XpIiKhG2XdHUUO+qacW/d82ffORigrpBmIHQTzNvTvY7oRbRPjRcBug+0xmOVL6f41h6/sWrSjK
STX03fgD260fVHvGw6/Q4+C83I81ElKkG0Q4LXRd1gqTf19u0Hf007s1RJcFsbcG9YyGJruts8ry
eRctAjymtoVMWLm8xrReVouN9zdKnHPfnmNHZIVkoF7PlMZvE0+TeGPGapCfJddXvQSYkzRN4xqo
3wa2k1doxRTNIrEWZLRpkIeihvURIYBO8XR8GNIcXf7h6pYw+U7u8UYg0PtjXnVVdzHcE8zX3N02
/UJ2mbjzk7ziC7N5KHlyYplgmiRVZhqALmzIQa9HoNP3hm72STMsq4uW+qB2DbxXuji0RPQcgNdh
UXSR+iK5hibSdnn0fj6NUiV863Wc8RXtDTWSuL3QRpt26iBI2GqK5xP2J4VZHSaZWoeDRtRnRQji
ssvQeQtPF9vmx0FxwwZxl1Aap3TfQr3TUdGxj0wT+Sx0oV4/mUgG+ODH4PNbIKduk2rAOh7abuM5
IEa3j2YPy3W2kmYyz0Dl3keIkXqPQzo9bjXLgYL+aIERzCtf+TXw91wAAFxwMKT9/Iv9LEeQyICg
2hNPBhEOLkV2l8xmshozyQc30ehWg/9X2zSnYVGWBBfIUJb2GJs6NJuxKWdmmcVvh+vYaVcYZJlo
auJxF3A1zUEqhxUe3eLfCDeOGG9p9f3PfCtJyOjZ8ce46SeHeOIduNkQLN88BQmQLrCthPPRoQFX
EkZvRqU1/moq8bBQH+TJ1NFSPTvX+GBQ2vF8cVXQ3eHpUevR2QxhgmHWkq3eQhs4CuJdhPgKh8vZ
Jqa1s4v+0LeWgtrndkwtRvp7VXA77EGBkSrxzvpGQEAxoI2gqRJszqPJ93/NW/bsVEaLUT7UTcm9
xyQlqxvWNXuKSjjtbCtUx9kwPSHNAUtMrMTj4i9HtlDRNzWONBYEtuLnIW65QF+eX21af6bUgB2h
xm9kL6rqJZ56c2I2+NEoJP1J9mryuEyCSFEiY8ovRvReJGzyT0XnpbUcY0ukFIh9QJV6hBCd+8Zg
xCZdULqYUJ3yxgen3f0d7DO5Y2kp3t2e8YIHZvZlLf6JufdIenW62eUjJh5XSiSYI2L8rR0TBINW
g6piTTAbsoXNQyKILo5EQ9OW/Q7e4Yrdm1VND/fnWdfhARFtwZbskFwt6kK98GOPNTjJHU/DjCiI
rNI+Gr7NZIDYRDH61WAjHCWWwAzxrqU5iyEzK+VQk8dC/iZ9ZXAKOrri6ebPXF4EkMcRnNO87TQx
TT8t6SAxUsmUn3A+CNE+pZHHWJ3S6/8uhAeTkYZsNyh5/0IBoGK8VGb5JVhH5EWrIl22HPrlzHSI
h/zwvLl4KMt3pnke0WlJQvj05TmO+d0DCcrVPheHYa1uhciwXuXVtEbG9kMjtuONCPhDceLUzlwS
WGwfn4Ox7TkQgATbDN0tTDb2xj0sPBsAwDsDlvqfYhqF32keMgTmpl8QvGXkxLJjYI63nM+JN7IW
EEBsiJTkMfzpfNddmVTTMoTatP+ZulwId/Z+kbXEBsMayGhPY6llqwy9JfueoUB3MlBeDGcFYOBx
j5+1BpMGTXfmU1RMyI63qjmu0jc7bBAqXznoX8fMwxrnKalAj0zBFYU59aXXVPzelljdU9COlOQ1
bC7GbR+7hZt4sZeUT73E1Zi9tTgLcRKUP4cOorextel+Wa4XmhWblHvjDWrzT8CWL2rQrqfepbGr
ybNfp/6KUYc2vsz86N4/Q9FgGbMTeEevhZe4rgy80QBhFPPpMRaOQ7R1UrpBj8WGDvLrlPBjuKy5
MCjaHilHD2QtAsgFiopyCKrkKuyec+11pJrrJ3TKl6rf593dKyI3OajrVeZ864aOCGdamwY20166
8fsqk3mMZcrs4v8NwEDelu/QVhtUSkRPFJApOcabPEI1i2345Q4QvFOxzagSKWnrKnn36VaAkJsG
LLpyupfSoonMXCtImskPlKHd2CAznLw/3eslk9Sx1RGYFgvrbZFA16wTvSOxq4hbe5EvGEjhxcrQ
k+JDNUk3hZ2MI2eiDgPm3QKAJTRsoENe27fWSyOV+xc6p9LMbUr2L29/cbNjkAvLUE+dlXeWwh05
XGzPGvQgeNJN17l6SmGMEgiYbYmfEHwlDDLEQR0ijL57enuoiKxNHRZOB3QRz7yrXejlWnbs0MW6
jK/AeNR/JB3OA3iQLztlUGEnLSFMZMzfKxLvWwLooUN2nM/ehZ6Zm3tHIiWzFdpyOMzvS0TznyQJ
Tv7Px4ZWXXls583LytC39BYFH3vxlzGcnLUhrR34cW7WIHvjUUtKlxzuSIpzK2iwPq44ooblCNgf
71eWC4WH03zZ0n8swXXFUT7dP72GRuakQ/xThzeLDmlxdEjWBradUQNKKmPowGghr2Xen+O6Rwon
WfEm3Z32o08fX/WT3rg1tg6/ydLO+E4IN9YtAZ906ztGY2hDt7Nz5wqhOW9WS4tVp+TVXMC1aLJ2
+T0fKsAMm3mhJ4g+QOhsjImHQhs/WXXAXhT/jM6E3WEKXMKGenmQKsvMAKGUr7/+f4wW3v9rDcdq
YV4xbCnmPuEu0Ueflsh/W5WA8y9cLP/I3TVgcWT/cw/GHCdT+VBdhIvRPH48a1SC/ku8aBUcz+vj
/HmHKrXXekvbIjyPRSycFo8zW029hcf9yLKEk1SDwpgTuCX0tixxyJY4/jdiENvDTruac8fZBEWF
gJ9UVBT4ZSY6n7v+9V1BqSiJiWoezYQlJwsWzPibvEqVAQ8Jk/wIs2MvaY6HmZgB12Ti3rH0N9o3
+mS5xz0N16yEk1fhomP4W4dzkCrp0K19CA8CzVUaNMyW/usaoxrgi3tjp+iYCM+s4zQnum0thpBZ
Oa60kaB7ZjcDhEojB5pbvMSF8Hl2V9hWsG2dn7XLYR+LpvINtmisrfkA/mCr0efTdMi4g9CiQi7B
4xtl6b0EGrgG0yjXBd0qkbW51UHY/++HtOfQkJOtOHn9q8SuSILnSwxRFNj/E16KNEvhum1EPqul
V7u2LzQlN/tfGELuBtyD0s7281MlZoxfPB7OYMgdPjukgIOalF3czmop7cXtJRfTBr/K+Jhfl6rL
3b7zXbzFx+gCrrtboQZ8VG0cvJytohVQ3VDLaxI7cjLPZZvTYW0gwM0T6mywVjrQVrZrYpHWrVgf
PkxuEONc6N8HcaXSvXUUDaIDNb1i6Mwsd7xXSRCqqPMM3blwWvqvA8tIgrhN2qPcN7mnxN8fCOZY
6x4oWvZB7QuxDBFcCFknDtM0JaMVzBr+ryP98QfjN54hlpGMtk/ZSk86hg4VaEJDVex2YvSMQ83Y
f1PrYDhGkPtRcmO2DhQibibxRK6cfvXnSglfgKXPSXmuDt1xilmlDje9ar+hJCMKZnRaxCnv0BW4
Bt5lWkzVMWJ96X8YMcZfahVRq7LUEOCzjOyoFugfOa5tSdlUyD3c52PRf/3O8Ztvd66bxY5dXR9l
pq6KHGW6kyMAUm8P/t5b/WjMo+9Q6OKUw8w1AArwcwtZmVeQGkgregNZi4MIa4k3FebOqGLU5Ztc
6lUBh/+UeuV4nHezyM4MKEMkPWsn2rFGljhryA2HJJe38n4aBeK+Iv0wTW89Szif5ItRE/0tOH/d
j5SoOMv79wqQa+9X/3ufYQ7fNOXBf88a9+1cZEGEQp7v5KyK6xDw0LqGb0ym+U8DkH/9hFFFyOda
U/SKSf4gbnDrWdMW5S0vI6/a+zRhi2GUsLqccBIuCfa4QhZe7+kDjjoixk8HLq2d+ACc5Vx0BCWu
FEhkRJbqGX/WKLW6Os2vrurzQARUiuuyf6AFHlqr7pqhOVV/87ISZvV+xGtawgqSXlZM1LHdUNXK
exkg0Kax/lal6AC9KMMXj2QntTKqDGZjEYTEKwCwtHQ+DjsEASGU1sFWjN2ewrpL9DZMXQYUdYNN
jvhFGruM0W4KUJgPpmIptPeRtbuGW8Ek9/snn06bx5cRcMcHnWpues0D3UuxO+FKmj3ph0FEH7Zs
0gr6zzYNLVJek37mRV2JAmlUNvMZxcuie/g3m6DJKybDSzTY+yG6oOUrIXCOWl4SWYAPGGVLA7Iq
vvLwlG1BtaP6UXNTKbLxhNT9+yNTlbg4VEVQE5/WzUmA2XIh90zg2XT7wwMdEIlcWvhZdPPirD+6
y06wJmqMt/lxur4UtsxAsphBZUjEoawpgUPnuJ3IjFYufh9mEKNtfW+859cgUrwYv8w/VdPs7+Ej
N+64TM/XJovEbqPmym1XpiajT80aQ8cgCGX3EH4duKmPD6cjm36OTQSXDGFJZMGT85CvtNTt14D2
lWkfi7xt9sKPBpGdH6TUx75egVVw4xYgtTEtEqUYrklaU1P2TGWwLCfol2g5n8hwAkSI2OlTv6Af
X68E9ZasT7ZLnnuNlxhVzC1jo/UoF07mZST0tZKCD0qe5Rhtvgg8V0TZfK9kdn3TLx3PL8atbSUB
HH0vpPlqm2FMSPDRp74hfVZKeNJElESevod+hSemfo2SGUwiyDq0K9R/FJvo8MGOL6Ihhv+cCY4M
WhyrNFW9xSppk/K2oiQjENu7u9DsQi1kpvjjrsrGnKxc/0ygACuyWUFKSddzy1iuKwIW+qavhOEr
xmu1e86lDYF2cFeXU5uqmH/M7AcAuuFPm8nePBAmR9pDZRv3j0IQoI3Dg+KHJoXA1EqeLc7iabcV
qQLTsC3xlR0s6a+KgN1dUbyBYa9RMPmqDe2M+HlEn3ZbdLkkP8+TxE9AlOwEZUxqUO0aaSHXRA+S
KRa4PqEf9cyL9Zjn+QFWkiTy9T82aZ1CX07ASL/ZuiJdmLlQ5e+bIPi+cyapWbTlDFeVXJONLwFq
YTWt5N/KsvFw8cbL3e4QvbEfrxzGXAwo5/l19dYyeek6Yn0oZvTgWZalVYmRr4W13CcIG2/6TlG3
3HYiLxAI/1Qx8Yrxv28voaqhodMSz6HfgzzEveahydIRoCVFu9MH3W7P+pJwZPOMO+Y3B3m+eBZ9
jYQ1srdaTs6hr/G66bk9Ojq7cLDAt5Skcvw4HcU4HnjjSGHbFveNwyp7EsLwXXZeufXRyFU23kM2
ClRLnTrX+qKl7fc4LWPAfDWFfiJF7ftoik7n8UsMD/SuT9sBcK8ABbIfKD8+f8tPK2wZLQEJPZOC
Og6cqUWZ6lwLPW86QeQ+gHk+vZq4oY1Lf8CpqCg+xQJgCZrB7LrUYgrIf8ssVLUS2cogBAvABiv2
RUKaInrlRRxCQIs6ydaH/drMig+12dORTiDHRfdRNCrIXopxBSPBi3EVRJTAq8HvqF/F0oXKFdVJ
Wyyp6KuqVeAH7oIQAKuRP1MRQhOTLRqfdWx7S2CfjOW58p67TYwz2fEw+1Rjdbilmi9GrDngBa1N
c9mZ61vaJinWVeR2B3tUL92PRkDz+5vBkTOtkFXupraPbtvDuXpErjIa90WDXVDhnme3K/XMUxJS
EnTlsybh6RuCx9l4MXUwjjjFKSzU04LJc8WDKm97DhahN51KibSBNkH/1Zv69XSWy57gx48HipRt
OLxw/jyP2Hb4vrvJaKHfs5rSV7fvihOeB6LVriPsKun0CjFeuD5sASq1iOjHFZ4QSRC7dNGPh0Lq
C+xHwxKyO4b3x2EwJ6Flhc45refPXIFoUgELMrR/+yC+Zhti8abzTc4EwqG23nHM6vuX+eQm8nbS
rSlTMDcR64Fv75nicNUvXn+Zwfzac6SnRTEYI0HjFU79V6YJ8/mZVvBZzBvtMxuJe99xTzNmlBng
SLr4xHRYFtyBYucTkWO81lCp06t9zpz47MKt04eSHRUYU4hh71CMjb0Kh9xdg9Fk3RbOP5y/uSwr
6Y9FdZri7bwUdg1NqRDJvA2XCXVFn79MaUnAlWUaLcpw9/NiGX3Ape/7w8N6iev/1QIqTYmF8NXO
WsYqnBxB5xfPjZPWGfC1od1AU2sqj+hnK4U9aBEJBa54BawHnpawDbRU5YfF44ifVbBxLoN/JuiK
KhortGuVyUzqrcLL2X6todT5laqee0BsUW/oBXsS99NRrwUoEZtkyinM6TwWwAZRMWlwyQHmbbcV
+E5lGGw+akT4rmvq52wV8bOGcOzVtL+ANh4oQvQqdQvcUZ+gHn+ZI27sKk5dfvfhq4iQaExNtQMq
XjaLBrAMvckdf8B2I9NAQWukzenoF2FiEAfLOpJBsODOZcYmnEolu2pESX3/rUC3V858Xu8VfRDM
DRws5OvdMzUQRIEvUPQFiIcjvtXZB7LzMpxYt2YYDopG0mnsjMDPQTQMmdWtMQcAzRKuA4yMjzBN
6S9oveXu0a7XSrSZi8iaGGokTJGU1iOpHR1F32fEzhS0HVEknbNLT0ymgbx8V05Hoyue7Nxh1mLg
8lCrV83u8j6X2YtkDq6KRPQZLHPzhJl3ofllLghQ0/RTmSXvNKrXEZ3mgJhg5jlwLgxWgMCn1sAn
BfiuBITUgdFe2hn1SBkpR0jD8zAqnODVPYnQ0/hlqq7r2pgnJtN2vYsiHLiQ9OJlO1OOlJmHqad5
pmf89yOo9Vk3Mr+IEImzqXAjFroFAzi85VABVgVFNsrayJGYAI6jadxdRUcqaHC8AHrk59u6oXQ6
41PZT4Ym3t95uch7q6Lqa4UOGRrZKfEJW61a1Yhbh2PAY875VpZ25YxlBRneDkAN3fJxA/xhhnW7
N4j0yIHrFH6BULzuH8vEhKJownZb32Y04F7/hy5w+xyAFChfB1/lHpRgx91JYb36RnvW37vv239I
3K+xfPUQnqoOYAWgU1KgjJGu3HGwma9rUYtTOLGqfwRw/QhZrS8Jrp/PaN7T6I6xzI2t5MdF5EfJ
AQNCXnjNmtCF3gRNyGzyBzaBSC9zy2+sWr0VSn+wqnxjGsAuyU37/9NyYgy9FJdq+yYdsX6nKPiC
mMI7vZaYJl7lGu+rfrT4Quhr0AArVdnDJ1/cN+SH0m8hgaqfY9gnooRSi3Ja2SoIzh41Eie4VSzW
ZXg2lhjrxoh73s+tCS0/+4coOs6wX+0/qlRQZdTx/nOqQ6uW40dhCm5kjxsqESdnudDZzJ0OETm3
9l6TOb/rl4bQvDDis73/hdTDEncEglzydJYre29KKgmmKuze4/4ZAy/l81CuQ+LGYcrzqFtL9g9t
EMd833NReDsZAaeUyJfQE13U7F7xy0/Rn6QcGqN01LZfWS/S6qXsIQi4rZMgScfV8Gzw9zg2+uZl
PzQ/MEKh7qfNZGpz+W4xYJHTxMKGHrtWNKUDbFxuyNEwTHqiKLTIK9+C5cngAIf84esPiTOwqxZO
UtOm+j1fpMdlhPgMt0v7iEWJyz+1VQsLS0jn+TuWCBNN270YsYnOHdpWr2x82HykJT0jtUVw2BVa
OfezFAbwFkYgZVDuxKJoVgQWl7EWLvJTM5wuVwYd9WAphJCJkRVmrr+j2g99Rr7pVz2MKP7qXfag
UR23pW+EIIx1TVRUNkCEnIKTCiAOzGW0TrBHwSN5tGOZ3TV8KfepsbaTV+c8sVmmPOnSt07+9fg3
l9CYyKy8xpLCZ1m1licMz9ZP2MiiVfXjr5mgcOh7qp2oaqm5psE7ydJCGNaoAtoIS+Uxoh1pJU46
aqqQDgdxXzAEheyhQ2okOeaWrFlNXLHk0j3+7qgqh9t251XAwbiUtlQkqErLY4aEHL0EZcqMi0is
TNsIEYW3m36mP70n7MFHzKxVhadcqHWr3XVaBBbUmi05pbtBpyqKz5bCV19o+Phhm1rm9YqB44t8
XItQn5jobJMcT6eTbQzsN1w0n9YvYKZHr8BLNsQq/oCcs5v+DZDONevvSoHvM6v5aiO8v5QOUa4p
EEBEASe16zYHoNB2oeYAhvICcJM4Z5tMsQXcWw51m/OTEKooQUrPHJr+C25gQF970eKiJt+mfxiv
wYMiHinRTPI5Z7tuZjD9YUkfGgdoABaUYudDHXT+B84r+3qvGU2Gh28tmnMcA9MtCkbiOgPF+ATG
zUDqfRBjnOKYw8wnokDMOBaoSnbDcsNJueIspHB6OGlkSUJXslziV1+pg/L/prAlvqDyoI6QYqa9
Ipe2EnLJmizIfVrhZAfnQqsmT5XXQrlEKwN6mHAE9famiB+/4823C+Uv8sgirbOts8ByBsuJQP5M
kedw6sJQGJ1S+yk/a/UuwoHsmbkNxRT2XPnu+K8QMxEib4nJeR5yFemxtQbry/JM4SDumuAg9Zmm
5DFb7od3IQEFTMLwoME+F2Uwja//7poeOqjWEWDwykNUzhZx6l7po2tacRiW5khQ7YD2x6mezBXu
a+B575jcrX88pYkqPmowbm+eGTTemz7hVUvQhZON8A2IqmdptHwhSFZfQSNRv2KDBIc46ciN1hk7
4VO/JMHcKzQPruWMtOxaUZXaNvXfLXEcDoLzqcVfHuSEb5dBTC97tuUWjC9KHxx85X06Qg1Eq5eR
oBpdGqhPg6TUrQdeVpIPnqBbO3jiGPQa4NEiaZUdGwHuVZtgTdz0v31cY41iW4rVC1V1a+w12TXz
WWGvJMzFzLhdV5etv0kvHlJSIQvHeryy5tHorXRj8bML7+SuP6uqduuirHlTrSt7hq8ks6jF65GV
tCSu1u1xIKGeJJuDiJr/zIznvIlO7txoL0sa+xQ8TvlfYm71NxHlR8REtnm8uADfWhw3Y4K7J/GX
cB7Jf3xsSV9iK5pCiKa+/8Se5+Ppmx+gs9IJbPGtbd6LTA4B/WGcUiNbIla/7GStXa2HJ533+7FT
/OHhtQvbVrozkJfQ27xMqAIPef8q78uFFFvXnW4ZLyAf0anfjLfSQHwAAnCme4+xcpO/KNGqP7iF
I4wuuRKLZiVq3bVlLPYLQa5DXqkVg7E/KUTBub0ppyaLvc4P4FjSa0bD1r1I68m9D/ePk8IWdDvy
lQh232RGYFFWy6pOwiHxTW3+6DwQa56ts4OeqIIh7PO9NvV4NVBOVScTfSqthLcVJ0JMXM60hOyN
gZYXe9xGR46xbXIdTzw9Wx8zRfz+9q4g5esTq/34U9Iv5Em/4xU5GjdUNsv4b8IyrnhjHZPeLivV
Hkdu1+tPfWJONn1Q+2jf+g68bRjZzdQZt3iazB/RVbMQ/RzhpJmYzXUPi3oMjWMSVwDbB2f3A4EI
G2IipczMM7CGzdzDPLz8T/rUoFcZUEZoYnXHwvQz3Sq+EXR+Qomp6alpDAKSW0khF3vIRg/ekuOn
JE9U7UrbR+NEJ0OIryFZooB4UCfKFqQkfkZzBxNjomI4paCpTMNt2RVbkbSWuWwuUx8bPz4PfARO
AG87HCL8PU5KsaFmtFphJa0kpIP80SoI9bC7JtxsKL8hHM78MP243CHmbRaIK8DNmYG/dByrAsj4
NDHio91fLVMiVLOrzMAr282Izv4H1FR0GCZ6L7vZIaFUI4MQ6qYJib7ubhmFtECPEzeW1ibegXWK
E91eYbtwklKaqKFNe6fZE0pRpx3dTmExreK5oKLWvYX6dUWKP4SkU+GJBxelstkiTQ2lC8HiDHtz
m+Y+OvZpy6yoUVtPBnsVyyxNVX8VbdkIBDBB5prT5cGt9vn9z1MTeJtXnWlk0ev+LQm127l/hclF
rgN0aKnlMjgaqWuCokujd6xbRsdU8FyMCJX8qNa6IU3q3cczv+vfKpYPGMzZ1+88wiAJQbnz4D0t
rgfSJQOtETLpFR94SJXAeV6GkpqK3wHJ/LP0oO06NJlJt7IMER10chcb/4CcRqOV56jVAOMxb6Cy
vVxIX6fcRoju8114Gs8cFTbBU77DoWu57GNbyb8+aRUI6u7ghFtmCSst7sTO55qCl3UDOt4knkeP
iD/mCCxvRFWyM0La1jheGk6RUvSAvQ2mb7LVkj99QOj9lfC/jVLXvJ72FGHC+SFb48ELyKZWGeef
R2Syi0wPowIKD+venEtrR236iB8t9Jq8iKslTPVK0QlcAxTtTUTOj63h9u2P8gr9AMSQc25TW0Ov
3FEb/PTXgiF4fZcfkHaoLV5trhy7IGe/e0rV7MknhRfMZYVYFMyemPQ7MT+oqzlkjU0JSMVscs2M
Ei82FazRwWcSm9emzlrQewebI0qjdGMBC/bCG3SJNP9LbT2FRWZMsXaFTCHPqHPZSirjDYvaJEPw
2VA9iNZcR8RIwRPCTfrN7NIGFcJ5rCpuX9qKGi5PxzQ7i0gkmhlZB3t591IWV9vRNJSQTUYmZhHl
Oa96RoXR2hk7Dbm7k1pIMSPuNwXBlLjib7H42nCiqYEqpcYQfsfelyh69MdXcOrr3nroaUwRVW+n
ozizNA2J9WekAYSkqMvksaSlFJbO64O5SdjdPPO5XBuDKSQCHIFw3IzgBBtzNII63fKNLIGgpZKp
JwScDKNfKa4bzRnaw1iX0ZPxaxjy7gQH6kimOLAljCcVc82vrKrvdQxsfpRLLxDfMrZO4ZqIShb7
Ym1qxeA2qgbM5gXDV0phqMBnqr/1D9Kz7g07hDX+Sj0TLTRzmhWAz6hnjNuYYFaFTcraySa8Jv7o
a3kZ66Ss7uNq03CmhSMblH3jsnRJpUvSOiNG6i3hCzDl5zZoLIcpjW0r3DXlvmwVZLwcqYufrMEP
WjtEwm+rZY5LNeB8jsqRmZsxDPkZRI2Qf0nhZPZ3sXDlsdrAYLru5PVnZo5FJxGq7KenMqgGCUYO
nzkAsmNL7JJwVmNKvrfq/PP/2qUuwNiofWYIXMFf8+1m4Ax2z+90U/8seQI6lvPZu9FCcCS4i0q5
t7PlHYoO5V0C+UWdyzWuxCQXkP85HyoHiR+CJ4Jpv3MVlamMWfoMt5lkoc2gkw69BGJjJq5omdEr
PGAE8pPu0IRA/6mzS+CqwqmvzJJEtrZI4Pcq30IQ/t66zzSPfdj/T3d+em7kL2U9jcvZX+2a/eAi
z6J/gZdbdW8X0pdWgOg+xtn5gwLmHiRSV7Q8b5J/7hcRZwO6bKCqF9hmABJ9dhs4FxyJFWF1gtmS
g6R5joZRtybH1tt9iVpm2+/4LxTtknH7/uvn2D7SMHw+5WXfBFacWSIw2Cq7j575S5X7cqtHvdSV
Cy9si+hTbb2Qf6X0zidFnAGRT+Hlp6hISsJqMxYY1ZH9hgJGQjcuQDL/YWPQzFSY/CNePdtQFVWN
60X8nmtJPA/WAM1LOUI+SvJOfg64DSUfd+W5lqkm5Z+3s8gd9OFPK8hRZHK2Crc5Ow75hkYhMQAI
VduYqNgmI108j0KQg+UBCQdgwskIPnHsM/OQg6tT4Gsf0LAagfu/LN4Z4zKoH4R3usbbpqW+G3Ij
EA+XUPgKmE2ZdLi7KpIbG5I6uruuDB/JZSUC+XL51/yTE3o0wLIqMO00zm4MzR9gi3367rfM5AR3
LL+4V43k10ZnjH83n+1TsMUzq+IAbCe3wsePPgN/q9yj0Z0w5HLYutC/NsBe1tr9fhCyUr3GFhiJ
MMdC04fn2mNFdW/tBl1Fkw1Z6EuAw2LURwFDpX/lUlHkY7EZGOijD13Vjy5SA4ER1ew5nR6WG0bE
CSjlwNfnvbr9sI4bStWvioJv08FZPIj/bkLpPBVdvi1m1Y1eezbmNzDC64Ci++aWqUvRCd4SnCKY
wA8NRYGq8C7v32FXLvdRqZsAsvsBD2jZ+jM+vJT4Y59/19GN+YSZoaY1IQESTYoAI21fR9o3K3Nk
5xH6W/uiUG/NaH/2SXtMwah9khT70evbxXTyn98m6wEU+QO9OD5fGuthluwO1+DKaQDJV1lwFmSz
upsHHvj2MDQMeAQlwgD8sla9w5P7W62i5+Znv/zdNdpFItn6iOxNsxVcCM24fJ8cYTb+INMWRU6c
WO47kt2WjP/RU9twOwHzj5PlCAIk4uVfA54q9oMsCNfpM6Vu5XwUnqqVKeG7Qnu4LeaBvd82HWRG
4KBc3qWUI6dcwb6F3Q51ntlLTkIy73zoKDNoTx4p0E105fzgTLUmRnKtsytngZ+iJN9LzVnTePTG
Ea26Is4tZ+6N/+JkjO0cnGq9nHtozVpG5/PvEChVtVeKtlb52/opldhDUzvaX3soRtxBSUVrKap9
9cKaIJiggWpexaFuJ1gw5dIouF0c6O9JaWIzDC8oS/ufB+cNJ49x4TyzBIbwY0DKAqBZ+WPc+Cn4
xR+9EWNIX/KHKEpHUfwZxg5EZxAVKaiuV+GY35NMFnJa5CRPhId91gEJFGg4WfvdyknOdZzwG/IL
3QLfMfM22vXabR/wzcljjwsNUF6AnpYaz6sVaBWeeT92AxsZzb7MlQBwmtnqN9pUTiR1Kq73+Zcv
thMjZ5JymVIp2COQaWez5yijsDXoRx7tz83X1RjbBS9rjFxnzvhMcl8/96r5gCcmkZGqeUOJ7N6R
tpjEIMv4gmjCHR+Tsggws3RiADNHYn4hRE/t0S1iLSkwZf8bsqyM+9ScX0aQt+kLnxas3E2Xva8m
9iL7cFCpqMlszIPmBQTaW8HiHhKpHL4mfFXguQcI6EMN6FfMdmLDqGniNRd2ViiHpn4X3gVjqIeQ
LOp2owYQXnsHcHx4zweMZuz8AmWshV8HZFpo5f6+t17LbYq7NfmlRRA1eSaJ4h63iF09bAs7xYM9
JJkj5vKKZ9AuknEF0IO1cGM+3LQ1dSlcX5ejjWUzfReyhW4f/03fyXvD96OlNjRWuH2SmH0Jcu/d
dtdXXujx3s0Kh/UabFDDopRqm3TmIzunVsxs3dH61c+d9q8WuRBTTZWqibcbm1r2YxEqXg8eSL+A
chGZOsSJD7GvRBrsgEwqjJheDF9GRg0JjDpCnsg0Adxoww56DP+2lmPA60ecB5RKItMuQ3YJY9Yv
Ed+J3jiJxo6m/kz2SffmmaSYd6Hosx1MKpdxFIhrm7iuDCHQgVtZCS9YUCjiSHFJv4e0ALXjUL6o
tQRJixX1PK4FYrx9Ftes/f9HJtLIyU9rgVQ1XiuQ4AfTxClxAnZIeIp3EXynGyssXQ28inecHXWw
wjqInZPpvk31TCLFOicMiyueWu5jzjkgmzv5JLjzOjahwpt67y1BdfqhboovzbvyqGqNgaDZm3dp
eCpjGWSlVQ0XwHoJiWGM7UvN656Z5PvC5QbTqK1FB0+mj4hRTIUk0cdKeGM7DVlAT0KcRhcJd7uO
Leb2In+oS5kkzetDHOO2AWekCrDeZoRHUq9dNDF3MboWMf4+Q9eRkJyx1+xp01Y49AoxfYPYJ+V2
mnc2IaLGEMEZ5npfNAW8Cylh8Tz+o4cbNK6/gMiUd24IDEBTviUl51ruxOgPiTukMzffB1PqC5B0
1q/qtpSd5zno5jzrJIxI597kuUAUrlaul+5M/os2F98ogdddt3GYL5YNSjshvAPAaXaTrv9ODooy
bQTv8Ugv3E65IZ0Xq+y4KxXH+tEBPFVrz77xjOOeixsId0wVAndBWhJ8+ck3gCmLIpQIDrjS1iw2
1Db51822JQ49t3+p/6oldDNpdqCo47eXShgJgGcCu/ok6n+AhRl+rw/gIh6xLIP62OU5X4ZbDRch
86Dvfz7P3MjW4AA71KYlyp1PiX9Wlye4ALsRlDcq0sowGPoGSMSzFEDWenGKtO9UCU3m1pm876yE
36dCmF/QmUFIKPROXHdJOIYZXMATOwjwk9vI1KSXZj60F+HwkcVvAUP6SdcdT/Iu3F2x3FzVk883
xynwMbVZD4WzlpIK29joWOvOO49N/Nb8IPwaMiR8HH+CuowkTODSJo+uxUzUa+dL9u/huzZegww/
9Kk/K7KQu4HDv4C+G2J4ThLwT9j9mv/FSA/zYyvOcObflv/YOd+Sv+1iJMhMiCnTKb1cyMugjjXn
7skLEwwdXN6rJyYZt5DEOhAAgDFk0LSxrizxhJUy/A/HBDkFYlmwMv8vG1y+GNjRlOmqSRQ8bUX6
QVpceJ7kcN3r+j1KlwMXlkNKwKTGmEuBRINPhe300hflmd3iwU/UpDB5eLYNGdvLXtpen76gLtqc
lbqoQlfqcn2/xIk3G9iJds6AHa7D/xxc0diUkdsEHODT+KFQvxKNzSbJz9dIba4ILvA8ZXiYBeWq
y0CJ4F3OzUJ8y9itiywTGmZrBr3DvKfthzdKCBHyXRF+nLu5xnLv1U1KAosFettElimDJp48OQ9y
Be7qKh3Ok8UEv7I+SChTQt1yqhebCIY0aoulswnoo2xdWir49tCrzfL+DMUGl/eSkWZ3OsOJP0/Y
eCDvCxATXf/oTE/0f+kWC8Tg1f3J/wuMZ2RwOGti8VCSHqiPNalnIPiipIo/Z59gTVRvfhSsxKD2
k3x1JPCoQPD3qdqu93DLn7CNf3xUQZtTkmoxahxr8B/0GIqb2O1+wLCi4dF+UJLfNx87xHSpVwgj
pz/1wZu8318T8tcBPAqwdUHuqE1k02Cz/WuHy/VrVBe3DEZN/XbAYseI0aApHAkoDdezWuh45Pbg
Xev1aSsS4pmZakP2V53ft3vdUtf5Vdw3ySFmvtXDlyJCDika+A5ITX3UxVcrnz/k5eHN2MfbOCuW
WmuCGo6DoOoSevpXDSBrZNDzXE6x0PjxvprKdid2Lyo2G16fZ9qfAyN6+66z2+idkNECUSfLeVgO
kPYHISkw0L3S2Iw9oqDoaL4R/CAG5N8/N1QtMjQY5MjMEM7J3V3SfrGpJTI1T4iN9Gj7QC55/bL6
nVd9Cy3idfgkxBAWUR6cuSdkT5P4oAzkcmMOdPWMSh++nse42hifzyDpaq+rzWEIUgezzMdn+TxE
JRVaNWbXaIYy4dwePiHWvNwFrq/L1EpXiiPZt+M4TlkNccF8eLZRbKFdy7jFwf+QCFNjVjmcfml9
oUwFSklbdG9kHEb6Mo/ZO8EgS4KMlzBWc1ByDkNL1dl26sRsifekq4eKinvBXi6mYp2wUkeFoZzu
D42xCsWHRpKP3v1KY9EyzADRr0Dq/7utNmch+UyZVuNS3/G88lHq7VlyBjMLfM3uvcn+8aPM0rch
mmyqhLHuu+LSfXh2515qr5NlxaJCNCuJcoC7sYotuR88XPEYEOZ3abT3SK4puefRbKmGx79cq4Zy
LrJupV1NbMTMnK+KCM3EraNXKaFhuWljT535dp0s/qrVT12Uubth01/H+c6FvnENRieG0DpzILwF
9otyH33kEDTIq+FJIJds8zsk+CElyhgHrMbR3HOoNvkuSMHM80vrUOVUn7g+Tbriv+auEhvMJayd
TFSkRqkOwBjUQGlFWnbGUAvH+2CaXMn/xzq2tcJkooLf4OBK+WZELngU1KqPkyLm7S8TNdhU1F+w
1S07+n9xGh1fUfvBKnW5QkT3WUZcVVH1ry0pOX1ndiHcxTupGoejCrORjQJyCbMB+TL+ZZfIE0xR
vzCxSpPng//XT4RjFb2FLFEMDJCYP3+t9VRIogy11doCkxsJK7ekEGA+8KJV3/DRxjg7h87KGiEo
qJ4DXFESKdJTZ295jZeIdd2cDJlV/oejFrcgFLv06x74qWqhOymcDuQTBsuHmSBkuSymc653pMad
iMfLksQP+L1l30VuZNZ/OksGQRjtys2Xz3+biHztZInPFK2P6IbXugffZCxkkaAdy1e+H7si2Y30
HBMat65YtAgPozb05pbhWKFSQOAmVECy/Idcd3pIdtXmWK++lmW3Y9xzNIQyzgfsCzXl8NCTaOhX
k93GiZyLk41P50zwWccKxFLHBURukxgmUR6vk3aUpbkzn/WUGoQ11qlNlYjxB6nc3y4V5X1csD+G
zBnD3GTPQRXFF0ntE3VyGpspMkHKPHokxrDG7h7WOFb794tobFQPyV6lKgFRwfvrUtRoYA0Z+C+V
nDaLJi9hZJhKo6yUzxmw6+3MP7miY6vIyIjk8wQvESXacBW4hN7zmhL9NrBDEYKlk1UMBJy4inAr
/3Q2f+60iWoPlHlwxA6sgbR8djYd9JKnDqWlVvBumdOc+qUku3jho313fII1AdBBt6kjkVrkG3mL
z1q2kJJDpFephvAULGQaQvn31lek7JqDqbXDF4WIEpA0WQXmDd3YGwPTMDm+9q+E5z9tz+czmIzn
Dg1mAPsKh5+NDAr9iPS/0Ge5f/CsyDrESgt+zU1HMQrxFyccPnegBXN6ryRV1HI50J5WapZoTFAg
4vwKQaYqt6Dpiu1VnHBZTUDQhj6HOKmPIFj8CKaPDzn0Cp96ACPivHMr/9OWp/RAl1TS1akwBaZT
F00KZB0e0GGVF0x+jvFPy5SjC+UtNtCzDaB+mB8NHbQ/wFuaWmkaCH3KH15Y5yfNMJlyLWS/nzan
m9fQqSGrXv/gRiiphMwYZY9/UdxEyDnaD3YkeDe19gTi5R5/3jCcVXdJ8j36SsnERTHaVaZS6OcD
EmZrHcQzGo99r7Z5bceHSiwJfWpXUrtdPfO7wrIBKacG0m4scSlmmyvbcKpImliNUFcZjGlgPOvw
VqvqWV/BVVnBmMc0P5wA0wbDUf5+gAZupA3mVhmcoUjBXLKNvLCy5lKD56Xl/Le0FGQjh5xm4AXQ
jDsTr4Co7Mtr6o08MkNP/+iwCAr+NPTZpMNW12qSjNqZe9XMyxaXiZfbF/0Cglc8NI8QaKedeZp9
UPPA5v/phBj56nU8tE9VORso0BaZ5Vh4xFhBdAJoDeOENhOrusmBd2bAvZlfEPrGIcy75ACXXtb2
UW4BJgz6zMBszfbxQBaBEP0+BYYQNumLFv9dlwjAYxPKhFsuc0TUNNMXwGXLhvJdFItb9MwiyP9t
u5iztUzHw8n0OZsnK7pG5yHcF/DV9x6xyEuo0PYGuCSgp2vuoGP9qtvdcWx3Dv6Pm0p+jFe2VEaw
XbZAzGiUbG+T4rtfE9sTZSO1dusOSj8dS5k29NqrcRc2zJMKZQTNjQ5/UkD0s8bjs81W+R6Z9aOx
TAdGdB9lv7nk5fYC9b7n+JSlauioZCyTVcGf/9SVkT98qv8ZFfl/WK/TJC0vDboxrW5KPIHwdneu
vauc2Zcr+0SD8HPM6bM+BvrP0qX5YxOHLZY1Nj2CysXxPTX2+/RcLi6oPcbEE8PMUjlzdG6oGZ5h
CA1y8pxn0546VCS3k7Tv5OhSGWMBPLcoEXZozL7IkfmB6lxRR2sny4eiWwaYeFWS0KnqtOT0KHcQ
ubOHMj6fPC1Nesp9cDGGsBwFTBUCdIvmBjhOTZy9vupf/EZ482pFBoWFyPJ7lsJA8xVM28p51AOA
gdgu5YjydmBnC9X/Jspo9s5PsYDtCcfV5+09ZYbAA4vNDOmKSTIDg9IkeCMq/ttKHKBPt2KoeJsu
d/4ZwA7/cgXX/JtA9XH5NsfDk+/XukQ9zSD9N+rtS7veBfzgQQSBJt6mb1ksJYjRvznEs90Noccz
mgFMbr+vYnyshYo0gwEJf6TfVgJM7cVpNpfhpjheuIC6HEuFp+oe+BbfKUmWffwpTx9BsgirpX80
OdVLy0Q5TnQkunlqGP8NdKmhLHWgRQqHeoWEE0X7j50QE853Fzb1LTgTGajx4mFs20FKmdTdP1dM
VjLWDA+hLVlKKxwqWAAbUNtUWCTaww1wchImga+/p1rzeGCBsuW8nqFp7bDq96HAA7YhINphHIOi
kl63tB6xMmHGzwzdFcQXS0pb/asrxa7EC01iVpzWhLQ/LB/r56zCzOw020+T19udpLL2oGh/wDL3
/jZGSVc9ACQPaRrEzu7knTmFapR/yg+RyLh1NA1cwtBFxXuKj0yo4u3WsSgOwm1tF38+dFqcyquM
4HwCt59oU+O9n3Ah2onF1E0ZLCDThs6kbzAfAu2Ha86RxelXB5TyDaz1L6mtC/zzRFQSn5yMQHNq
mjzgCX86UCUHXYuvSB+81fhqE7BE80n5pGw5MSSFz4LDlZntKHHm996ORNn52jEJRDJJ6UyXaEOe
RkAnAYHxyFyIAMC8zMe4GQWMZM24SInXQ8bsrRbAizCVXV4fr3vVMqx3sIk5g7xO5FnrcDKwfE6n
KQwr5+WC/vkm1V/kdCohKpWIL47pGryGLk617V38GEupxQ7WmE8qcXw1tnRTqNutuAZRKRDW8tT7
Htxz854nbCagTQmriAVpevXau/sj6faoxP/qGdmSYeb1q74fesPVcIPf79EIfJS365ofhVXznjy5
wOfdztbq/Whk8Hqx5htf2TVWsv+qhueGAVN6A9o4v9HFxaNq1LLrOMRkIIc3CkIpxbcKgOHOogEh
tbdFtUJIE+4PjUruMIlTCWXKxh7y7c7xsIaaEMcTOzH4s34oqSu6hpWlrZ8F8Itelm0HM7gqKx+W
4lss9Qf1FMJi1XdQC+tsRu7RZGKa2J3ppM3y9dB4qYBAnEXEO1Xhw0LpjDWCfmopn2mkK4QXrFM7
0c4LYRzOmTl6AqakNKLmv+wRCGK4DVF33TW7nylY8XVkDP8aHQOfE1VcGI0fQ/CiYTcCMYtpAkne
Hq8PV4r/hIHds7aChKIAkAouxhyNMUrrADh9VQzOIf3Rw7/WK9mBqcu34QE1v+vFN6/HZAl4253q
4UwrNWzDKqc/xnNwOQbXmtBNM7WHhICKX6n1sLiYjoCG6mo+FPy4al9r2P7lBXJKyLTkqxFEvxny
yscdAJuVLnte5pFxj6LF6G5wzywnedsqtDn4IbjpFgBcXOJgROYz5WBuEBsTOrLOAR3aFpEBTsbf
SVZuPhAdkvlItPuqMGHDB4U8ClKgnQAmpkIRyQtCfWBIbQ9AsBHP+i6nqopklpBSxo7U1yBd8MCv
yqU0aKaLkf6Qz6UlH7PRpTpJ2wcEE4ZLXIrUkO0B13mJa9DoLcnIRjQun8wYtMYewsLAqcGAQ0zi
zIqfXonlgYjY3LHkk0BuW/Fkzn3RkFaKu288F3dCQiqVWGBae8Wky6kT6GpingeDZ7D8Px7CnBGu
Yv19IXjB68wnS5tV8xQ4jUp8Zzygcy/9Gl8NdQ96ZV5XcTKnCbJjcldKMGxYDxWlnbYY/j7jv83N
1ZitkwKruvtFqup93jrWfFVAQg3wOafo/s9uPgW2PlDzAxWtrCAeH2n5owMOZOX0L28c+u4GmJ+2
j/NnOzb1GsC46qZaJNRznbKP5yJVgn5VluSyRS5qmMmHSxhWxiZQQeHAcZwosqUABd9D7u0cpaVc
WdHcAclHnS0Bzqiao058glLgV36xNvTqo9DRHipI2UBmxCV0TwV0PrtNgjYmttr4NV/o4SViFjvR
O2Ms8DmzqO3UO71TR21Zs7aYgdKD5YkA+e8H+Rnq6CjD5MF8xLFhW37ibioRV0D9Pgx/t8A1ohEo
RkxF/ChJR0q9A1AD5jC2E7atbTl4Jmrk6UdZDxpzklh459TI3rOBFhKY3lYR4dlBiTtz5l71NQGX
t2ZJpmVE6raFaaJR1HA2fmAAOjriTtctEZnrDkRymoJHSi5OMrreBVrNpFWFRMyCLvRmYBZ24tIK
LgaQNNpqox/fNT4Rx/oNbL18oP3VGagE84O3fT+ICtNWMPBJaeiX2+MSCUI7mSfclsmzGcSxuy+C
DNSyiBnGBiJYaNvHU82mtR9qdxPZdf1e+x8jorncVZ9tFhAakC9INfOYRvcBHrPemYX8bpBpsidU
N2SRhSbbkTruru68kJTZWSpmNclZQfOxwV6BgJVvLSAPw89wq1X2PVuJqXhItKhSEZ5N9JQiZohn
Haygm246pWw8x7g/hBhlC19TJUYSvgmO19GUDV57FRVc957HEuuc6TLqQ6sLzsBaylCQNELTIvzn
vqHDq7Kx6x3tDT02VCVc7b3wLENWou6ZLwLboDguG6WwtElil7//ATgiY0eIIvVtyPozMmmYh+V9
Y0M/lgRbsmyIEjFFkhxDlpJ6pQBBI4k6qTuDPaeKo6nhR6oSj0onab5s9l+8VcsEtHW+t95VLZFE
fUmeYGQqXOSLJPzQFBZSHAoE1hwaIVjrYoXBS+NLC/q+VcIT4Xiiy4FKPjVqOodo2Kw3g/eQKwbF
31482KO4QkGag8wPvZ5lN6ODJh1fW3ArssZBegAf6BbE5OujtOsMu7QGgh9mJCUN40fjwBLHM3MY
EDd1Xz7+L2glkysx6kDEmVp3W0lbEmXrjgdbHL1AXE14AMkqlF28XDxDo+KKyExqdZuP60bOecP0
ljkm5heFtXgqtBgPP7JoMEUkgYmYn/BW1NsLwVcdwx8KyJ4Jr6erYvTbNcXp/77vZGLzVdKL1FZa
/AfMcSdE21gSwuylZBZiSYs1vEJqoKs28KtsEHL9alR/T6oVm/w37pureYVyEj1I6vbWS9gOTnme
JGGi9DbUzf2WCuVy9Q4qYBSOROMQOc1/Q8v192vutrVnRQh8pry54Ev8/sGh1MSBDA4kv5TJzKx4
kKxy10PypB+YsjEnWQrxrVAzdOwvu4P23Na42o3gG3hTyr6QQq0QEiyd1otRMDqY7tGijEGOPe78
QaWx0xg6L2KKDUwibNRee0kX05h9TSEetcd4gsbJbavw+CY3vQYU2nd5jOOT0g009E0pPddllL8X
G2J90VvOu6JoHw4nBNNIpWTcJG46b1B5A5X39Gfeo9iB2rI0MeXwqLSnfnelMBPJUqeNW02YXIOE
LYs3mhq3cbsB3cP/k521zNi6vxmCkKPOtns6/9v1IU+e54dVmnQUOPCc30T3qCLGu9aE3YG5a68k
/ziXnFTxb3vUZ0GlFIqe6+XSlqYD8pVM/G9aJVqbUgsXkQ+cBFfS/T2sp2xM8spNWm5nuYvRRdzR
GyhRKtPuFS9b2GhufNVD7VogdRnIBsEm8XnSNuG27NA7puGFXi3eskIEP1zNyLPRNcsyRn1b1BL0
pcBoPzmd97EsyAglWU4yv3+bm0EtsJAXoP8lE25/oRPeGVPV74fWTbBvEoh/FCpb4xq7YAjy6Xnc
kYbl3ctuKzVI69P1/oQVqL+Z86+HRfzHRineMh7JIf1ffARXD1ic3gb2kWnGKRAT20IR9dX9HZxQ
BrNmgzO3ndl8YIV9M+SThfVC0vFF7o7ED+R2AhS55OGTCsywGkCVO5AHLmF5WJZ5ePPyoMYX9UG7
VUY5RfxPJ5B37fBRWDGOuvP14EgP2PNkG9qRF59BBoS5wm7OUnrHntwHtcidd7cOu0bvHWJn7ev0
GqyqauvUXR8oFg5r8EbcB9UxFeBopAXxDBXPYRngs80Sc1aWAkBq7c9zE4JSQfLiFNGmumHZtucU
nh3dBrruRx7jxAT6v0kocaPRtLaxkahyGnTTyg5GVx+o6MLzR7gncb47D01rpa6k4j+eDPxig8fl
Z1KW+NO0CZJAJjBlHCg8J6PFBTD5ISDoNVrZ7YIBDyclYDUklEnqTwRtavvEKWkpFhlkI1DvvEqt
s6UysNoxJxI4KVxCYuMZbr6qflHLkkjAbDUllzBw2GGnsH+chPXrGYLoWVaatXaew3E2lMz96qhc
eeJDK0q7AFpEzCE6bMyXCkfwVRVpo5Dp1eZcuM8KGQXZ4PXjrenhgvcmCR+mGIBl4WMUXlJIkYAW
5r19W8t3gOzGdUyKJA4qI7H+XFhb0scs8KngO5veEwfTbEaDcf3OerwGTdciwxgF/oKBb1LPTxB2
rGmsY9mbBpG9FKd6KM8i6nWi/vxHHCJfXiGSHXkNltF5NGBdwcTIlJL8WDVLhYycB5lFRZXNajQz
vOBf6XVVid1YbHSdlBTm3Z0BCY/afvdJ11JiMiBeQ+01aZs5EF8hhGuFwF1UKn12DrQ2uEcSohqb
O5T+RbY0x9FzbqzsjFk3VtAwZb/7h+o1HwlOC/5JBZuuAn2hc5FDcxTwfeABdzIuuRn1P1SppRcL
e50Du6KtZwGOyHaZqq6roXBfqU73sNRJ0EBZVcbyO2uFFtmwa4fTzn7v1/8H45/d8Vsp8yeIpQbO
yEd+HtpqEv8eAdMi/oVnTbmKVf26i0lCWyX9ZSQsGJUaXcIByisqy8sSC22sy24w2toN2GiEuyEJ
sgs/zh9iAyz89r7QcR7VKhIwNwsArD4gXwWR4bPLdcJl5Y3Vtkt59a+JdKulQoN/RU992l0Of0tt
tKPsxhUC9ukZ1XFWXgnrIPluTmxgGsAEWdHcsObe0GYAPuPfWCQwPVcab9ywGyPJzLogqS3MlXon
1R5AFFn0oO9lyzpUohPlYhoZMQOxy7TY3rpt8JInW+fCeadvJbBe980Ez33PqfXJ5I4GF3QVEfeu
CWBxUfagNdTiQUHt6R2BVB04K2pKGZmmTNZ17tH9SWLjOnF4N4HBL4n9jVLmO5Wpka66TS3qRTF1
3CGMqTIzCYkJDJwjDlviOtQeiVpr+NOfxBue0r050nPy/YTeHLHcZAJ9wFDGBrxZHIQX09c0/loX
5q1cvONtHiMjBBBOwelOFxDX0vK5pQr9VD5CJp23OJlrHCluUrGtx5NNActKe7sQh9r2VmT3Il21
gbeDhf9qm+sjlkyWMdoeeEyHF8hkRJS0W0bShSjWmYcea+d3aKwfrWGSP6maBgAqxHvNKq+FdinE
VN52r55gXZEX9ujf5seCZSJ0xdu6DzQb0zMNQFTbIKVQpPE8IC646mIR+Xd3urDFXaHPiklIbrmp
mUlimsCyDXNiPprGXcUptjK9+cMli7PEdBbqnZ+svASHrm6JB7elBC/N9oDhoTT0+TrXNyCw1VLc
R+6gHBJ73Kb3IW5wuh9uhyRhtKA3viPfYxKPixTEru1NmL9uVeda7G4Ed58Xnn3gEx0tJXK4wTqF
V1uI+ulOfgV5sCsxu8gHdKcv7tenNSXSJDEWt1Qf3TyQ3ZPs0aQlVKsEDQLQzhBQUXrm1yVh+Mm3
rxEF1nYB5MPj6PGK2Ojl8BItmLx0lUSYfRJA7p2SfXo2Zz58LBZ1vtDohiM3BnCuXfXZOiGUl52F
zzOgrdIIO5B4xVLtsAodHsHsI7lvXqoJpF6w8J/IFOpNGe3TDXC0sV/5KSFL5i1t7HzCpulD0MmE
py3iPcJmIYhe8zY88QvWIyS6wb/IjYxx0grwoUqHt/Ln9LLvRmfLRdOooNtgWMA6RLnF7YnFIhXn
z3xxpVgV7wZ07JzGJ+hdlKmmDC5VGcsX91SJXfpLsgscm2x6xyWCd2qz47Ex9UK8oaCCybrcc1WX
+BSQzugKqB50uDEWqobhPoStSO6JNmvy/t/GSJYHw0Vb6HBki1EAmSF5lZeMoAW0xQoSYl1p4d2o
m507e9yxH/BprG3TNUvmYUnE5W0x0JsxQCQ/W2QIws9zwrEVJyEtyvnvHJsU/Zt1ruXofUIRAVHA
Sjwsdds6K3Z49GPW54LXXnH85eIb4CgKYmb9RJmdqOGMWB/qyWfUzQtAE1D5bZaKHXSSLiByGtRa
izye+Agzc4uwUQln7iUOV69Dp+/Zuuj/PIuVhkHCDHNCjw9Y23C8jIyU+3bH/Dm6B13OCdeUJUS9
IOYOI2vEwn3OnXv4DhbxnM2D6zkYSxgnvf56wBwTybJXZFSV2zWQUMBt7/nA7ZETIB7MZBNXnJS+
VKc5jfeJJc2Id0ydXSOJv9mIUpHZ2umw1TcUh/UrM5Fs9x0OHJJS0MdhbAX3anP25iXzgh1nG1NK
znziUOVC/jBJ070VNFyBirdoYtpWDaVcxg2Gqajgu1dT8dXxKwIDtVUi6eRZaMG4yUow4gXClmzw
6LFfr1WqEQkTUpNYYma+FRCyejabyT8EHdEok4D3vXVOrirdITHZZETvJAIZM7E49O0QZb1EKTZ2
M41qVhJ3dcc96u1sgKhYzE3gE4oD/DFyH5RFZv+S3bI3tDRgvJfWD1I+Oo5ak0/B7yL1KaFrQ5rw
iK14lKOmP9b6s7aGcbbUcRGxoLHvmcoSmr3mShNjUJApE/pp8qnXwb9pZ6mtbo89oSCC8paIhs80
jjYTdI+lqGCjCOGihWRVgNL+6E0LrbX3ZZb7yi1ZFHBpEeDohwRHwr6lID1x1VgDhpXmbRKUjHcL
R6oePFglil31NyJWEijdLmLXGSKOUBSKSnog2rsq6atV25HpVdlj1thx1Ary9+UmDqEJD0XyoDdN
/SJpAJ0SDyIUPVbAuZbD0Pp3OU0IZT17EBoIgzc3hTeXPlL/gh6QvRqfoDx8GQefFqTPhQ+Ndgw4
EpaWUgW1xWCmzLpbSx7ZbilPmEVezw7UEPoKt7FOPzAM1d4pYSX5K0Yfxdxo323+hk8/fsgsxRT4
HCvAciLTAfHuMq3jLZOMnMHQXFsafHpVYALup/AonR8EK1ke3wFvIB0c0SRzmNqQ+1YyMVMGAMb9
o+eMysZNRcpAKarJppYGa1+AkZ/l06NDN1H1G4favezU33Xjg7OZG2BsKrwB79EeJM1xaPaT5REY
M/DSb5pLbghasQUchk7cr4RWonSBJXTd+5IiSYRM2dphahLt7btNWclmJgMGeJFRbfPUe+pDYL8S
jN4TwVrMYGHpIYL26bZQtTJU2IJXDo7dF/N8KOgW+O5cxxcWHHCh9qIqwSbdslzJhPf+dXvIwlc+
ghYKNwu5qZShodcPUn499ndaGtQVg4EJjqtFQ9feEbvKRPm7vrBwbS03GBkwkQg/selP0Fiv4QPX
5KQNqTWpV9g4ExIBOrxH+ESC3CLbYgJRh26FeePfhxw6N35ndJUSzS5I82GFBMj2T+DRU14Op+tq
WbbunfxCpb6DY5kQQt8ThU2ds/PSLv4wapSIVdPjGBSaxj8fXDgYlTf92xKA84ghE9EJbLvC7LIv
kcHJOp44bwBaC+NncNxFEJ3sodjWHnog3eXYoGQWEY+rADbpZKmAkFt5mwJX6KxILoVJG5KyUo2x
DKSYobhLLw2bKOb7PEzzchTgkd8qIZ5syYhP44mVwGTrF9S5qJ6QjywXwjcGdh8keK/8B22tH7i8
MiLw0PjQnZ8ZZgD213DfvAXgZ+cHZFQziu6HfOp6j4D17FTJuawtLtTINZQxo7lj7GqJCaYmwCFF
1uTqoww1KY6n9FGi3mpb5RqRLjOsTQ2d50OawEyfyboLcJilHFmW4hEnVVBZaw70nIkKp9bhUMTz
xHabrYDm2P92xO/RCFJzXeG6y6mbtQOMMXAmwJe2Vxm8uDJSPA0ClxUa+ZTW3j/elAZeyxBTi0hu
ZhSVaIuOMpnbQ35tXC+IDuHhRTaUCmQC0pzK2SsN6S3kVDMjFT0RNFOhk3hj5FJGHrKVQpwElJSu
T0W1QoLO53k2AQLpYXFfVeRtzl9G5Y1c+g8rhk1Vhf9DQPU+npF74romB+Nb0zUXuJHjUplmPyqW
QL7FVwJVVQ8FaTKbnSygCjh0hVKb2gJfR1ZSNtvVHWBJWE7Y4ZreBWQPFgh63lj5vd6dX77sqL0k
VjPo0J4mAQNX5Wg7WOF+JWPinCmT/OGDYKZFDftY+Pob0ZoYE3KgFzETE9ZjGcwpBcJXLKwqYxhT
viPDAvs8BqduIwwyhQaQzXrbekAD6TpmsINSDdig4CGVOjG8cRwvEnkaugmUvvE39qyUpiZrsAd8
icykZjpvWm3dgtukw4ImRFouFcsS62GPCgWe++GA8b8FyC39BkCNdvJOaOg200//YUU7k0PnC8n2
fQTivuZaia60kh90KsG7MZGUAWd0OZ/kMo3dKScfDZGeZBfvb2tTVuFDuiIVYzeEWYzxWp90Oocd
BlcoNlqvanDcNVaRtmjMLS3Mmo9ac+OGL3OmJXEePAOvSXheSSYWY3/rX59LI20zllYmShE824bg
WktyzwQcw5Gi4H+f9uFBsoC/qkMXvSB+bY75XBjPo6i3MQpkplYeV/XfX/EZiiyb/UDh2ge+ze3i
1gGCBJrrNd2DoyV5Mp6FSBTZhmigfp05G4RJIahgozpsBzzHV2GEsr36SVZwdeMTWMuHLozA8Ws0
p8NkLBDfkxeJVLyl3HM1AvsxJLWjnNxrknntMu0qW+b4u4U9Hp+LdSvg72SHKXX5K6RzGCUBgrBk
z6tqmFb1Ev6Oa/b/yzCRkBD9i6dNpgU337NSTRROnQFw8jG8UoVBOg0emao89JpKNYmspK5rNVWL
HkGzOfn+6nCTAREOhSyrKJKlZbYs4dQfTL00CL8OQnIDESK7orIOiuuazMfACwNXXe1HgNnpCfFL
2G/COWUxVI/vJRF4NSECFn9W4WFB3JbQJYCvWXis18vUCTKNCBdFR+Dm4PvzSCNmcVK+E1AdEqal
CWuqn0jKgtNBUbW0WAuWFDfSrozaa7tJBDSjY10Vj6WW1P+8RFkKJhurVVrqygsPxig0K+eFkpBU
FTyTlWQcNG4D8AYOgPQfJpQpRkL+A9qGwtMbGWWOP9c1Fx82+6fd6BJANWqmvIgeBWqNP5RMw5U5
mT9hy3eMZq2+hikWjNx0DwFAftOkR83v0VodNku0WZ8UZKAjvx+8FQ6lyIQT+uzBq/xjuzCqsrm0
jAHLLmS502ehPWgaT9SUU3j3nPF3cpW6r2+pY22TnwyaUKWK4qsd633ucegWZzR0UlT/naa7XtC+
swdH79ckku8lVKWmgmbNsH18N55WYFLiPNCjAfcVvKbzPOyy2IcSNFE76lhbOJV1fRPtMvuoxs3i
WyOQ8sbdOC1DGNMfZ33YHxwFiSEkguUwWY3CyzFwbo1rrOHnCRnmBCkYuH7sjEl/f4zylKOpcsfS
qMCC07ctUgFnjbv+/dMj1s1qBDulsgwFAhCqqu5fkLnVs9p0aNiRI/nSKpiXmZ/NOeER7exgvvXT
0KNIYbdo23fmIpCeTm8a/XwhSKV7QjXU/prvz4WRim4b/dLsJSxx35xYkHMwAp08sm6Z2WZ7xLqJ
6KaLFsQDTjWXXWGela4HTvUEdCdNCNxUa2QdZiImcwZiUdrZewSKe6niAbql14bOBgiRrOzij5LI
/5LYfqSPZr2JX4gvH6LZrh6sv7hN0rnKDUA5GRXtCAyrWbKGXrAYeE2xSXkNa+UwfU2fe3H/bkYu
xAIjFumtLDgz1vOcqTdhhVzaGTwl7b0ZHIy1uhpRbjd1Fe0hViFLlitWrkgvufoUH+YxHjxiyRxr
Z3asVF3ccdw6O5n4teqAAUS2XYDlUFB+xV34757pCF81vv9SkSAWlDRWgSaAk+AXq8nB66glGn0Z
SO2KLt44BQCnQ0JNHIEe/4ke/xjR7iqDMKOtuiVo3tFak5J01iA47qn8zg7lz1HSrcV+rapnVUI2
USpZfBPFWrYcMywysxK8xvI6FO1aaEkODKIjcZXwRonYvOUgt2svj3L5ZHoRAgQSzzFZs86e+ROD
Pcghcb4IMFOaGFCJ1Qs0Dw9SEmqldJL5tXUbAiolzs0f3nZpM6VJMGs1FAvsbg9CLafLV06TTxJ8
2q1ECubO8/PiWYjNViNYcQXGG2r6AgNCM8YwVw6PmQbdzKc4h/7jZMsrcvKGKMvshxVRMHqD15Ck
NciIQ1Mz0uWFxB91oifEP8k8vq/TgXsKXqErp80h2BdlyeuSvydBxvXwA48XEn9YYeretjQnHPF6
4JDejuSZuT6ukDwhXRdQ7c4zKMVhoDtwulHyfmEbMw1+f7vOTce49SB/IyV0lt2E11r/Boh2S8Hb
ovWLqETNb9SeogqSmt7ZClNXoWI44CvsEDN0fIWaR49uAr37KOOIBtmOdyinFNtDtUiP7FuXA+BA
hdeED2ha1hc1hOsGGzNyjX4WKYjGQQikXRJz7tGg+NQTzAN7xPVA1Q07/BmbYulidPSWmSy0lPpS
Nw/KoPYpG40yDQAECTVfIdonEeAdvBbmHAWcgbzxesiCo78EWKc6dNHyxZraEkDBNtEtP2aHxwZe
1A+rfr/IixlRCoIydIW8zCxjRRHPT8LGomx0NwmDrVgVI4l6VYT352Mx9MGNzmIewJnXK7IBV1As
DxWUAMJ2HN6IhN2ho9MlifVg0Tje9FYA5aSMUVsTMkBynyXA7sL61iXr3OGRxl+1cXVj079aOlKW
OI1IC75BjtXFaz8yB9+48wGsDQaw2w4OEmLL4nw4fYbx+OsSkhuAbi+Ty3V2DJDkZqGyHU6vJbWX
vIfLeMwwsnanOznwNqyiYl8wLi3n8PNAoJYsJHU2SLdRMl8C6jNBg5cm2NE7bnm8Ml15kjnNPOpn
gI5AG6zoh8ALv8WEFkX4/7i9wUrlBfIHpX39cOmIynMa98z3vzcud5XfxiZVyupACA/i6CnW002D
GNDhHLaIvm1rlX9/NZ+mSDv0Q+r5E7LRnQzizIxD7UtM5uJ/iaT3I4mxdI578y19DHBMNVC84+AG
MbxVSflbbe4WPUMs8kVJG7gg/+W5bHxyRFDvGSLyJHH/ncSW5UNwwaIjiR3WXKqXgUqf0kw3/7vm
qFmrzWTsO32E9e4+XCEUjVyx2J8DP9w8drUvrAtyaWmV8EqGDZisp0sCOvJFpr0z9iDpPlB5rVVc
Yt6XIeGVEiJOPcz6Mdqi3oRd3SWu1WlFE0mpbPfplOT+WaGj5sLnmrAnn44zxDkPZ+UtY3T+ZgXU
Ey+Cdp436l238VUgWaXl1qa0VWUv0SAXECfiZyI7M+QEHk9MpJeXDkwRbghHcUY18ojutNN5wNI/
VKsJkTl3jU7R3eRlhe8wCotwi4i3oXXS3/TiDgOtVbp3FODKDSZbYCejvbMosm+AN8N0gS67M+/y
W1H+oOLFWezPcc4DAIoz38atBxLbVfFMSOVIuMGLlxi5EQvt9CM0HZqllJYcH9bRSvSctdNq6gLr
oWEt2MxnPrgKA34S9wbXnFclpb9YD3FDiTXbuZZfqUxMEwipgGrLMviMBpNP1Q+uPJSwkpAXqRTq
a9Fmbo8ZTI8sA6X+iMay8l4/yvaOp4lI7T7uZwAlye6uaoMFGsODUyJLyctH3SgRC3V7jsgLRMCR
Zqv7st4naMd15TRdSbo69mnHuwKwsobpM+6vl2gnNKg0AhKz87qFH2gNKezcEAoAokU5CSuLHidM
/T/x/wxK1vtRHysKqmFSPjR1thfYNuvdTzQgkO0oEP3S5UfJ0OPZ/7XLrNwjcqq81OR1SLVO2lHn
9sW3sxn4wnQ/in2OMiR2ualY79QyYght866kCGCA+FWNZuouwMFmtR5K+5Mo2xMxjZWK3HN2uW/k
pvFs2pgb+80HI1qkFcQNd6c6LlHSvNEE6VORjQGPD36sLvopgbB2WCRyLVTTMM5mE2CtHEvBNF0G
BiudH0p8/cizrK1ZnV3mwbWL9kiXpM0xYxTQEutwcoygM3tDfDuMlOj2Zhcn2KqNrGcI+xss4yY8
Ds2CvyyPqli80UHDcFWs13mBew+wCnF27592VIXOs1/IDjlpooM22XWcqqTtyAR/Cc5nPlYnCASf
S+DQ6pf7f4OXtgtcab2J9gXGbRUM0Y5d6rQML2yu4sJo4YunuVx5FLRcI0MOri8ozs/VL0lUd1rY
KPYmMVze2GPjcT9M1ifsUruJFRAsNU1hh8ZHBeTZyrjKclWAVyPG4stnbApzpzFRIB6gboa2oZou
4NIOeFgG013vI9HndR8M5sNJDUar7ZqdQiJpGuQPJcKHefVN1mwM/yi+CQpqiJhq0wXBq+0/CPOX
tgSkSTsQ9qcZ4H/kVh4HyZkjwiLARtCXW0VjU+rDkYU+4zlO7fEF5IbcVExCcWPtSTXxjm6Jl4hA
yPjd7y8HJbMqUwSHTTPwkcqU7jLJS1qS5D5kiu6koMkU/qZipjLvndYolEbNpNEyujjzaM6AMRVW
XS7s7t2YomtPQtxs/6vEDV9JPLGoia//HhdXJxdsRZ/bPcD/WYrvDgLC80OkgdVfx5J/3ou/mpq4
X6aRxP7aBnDIfGmLv+t4PNwVtp9yxLg05Ar/hGYCa49mp9ogwUQxcGbUcjGyHAJJ4NI4d68BrNH7
/83zYowDdHY1xNEEymyrWZm0u/4WyHJat9tlruW1Hwl1P3mLOxWh5X8as2pwaShj9l56hz+0P547
yDFLgme9+GZdGP6RoOBp2EwGwZ/rtdfb1nLE7UKqTZ4TEOKzOQpiTVafOwmgsJhZetu/ujTFHGtM
1NJfvsBXUNU8PfAwT8lFyCqS1nbc/EQzGl05+0C2R+GVBgvALHwuq/IlvwULjPVRVT+YX5hWOppf
YM16bIO07260xPbNab6Qxs2uUNN5Y2eAJI/hc/0JgrGSq9qvP/rwQ5amhdo7XeM0GKFqScwzx8dU
XwjH+XsgZdrwzgV8QNZBayrTcEGr9+Q/fLIf13XK1e0FwbGeswZUX0wyAsRswwZN6mxMJ5ZsSvb2
f2AWysWFjWE90+8jiQEU+7V2RD+MXvFUUk3ZMCHD9tWZJri9RAiAsez+wRZWEfhX0ARMpD6TsiZh
V7xaVJXMeL/0noeyMnCHAF1CWHLkoeNi0kyKZQJJDOUIpSyDuDoKvuCWaPX4jlYdKUUtRTjiBdmp
GM/Fh1TzhKZmjUVD6ZkA8f6BIgTx7hpzuLbVRTVYuUB6e+r1XOzzqoNvooyjprUmh8IrpSWnrCgs
XAbA9YYdW2n+eexwjN5LnP6go8w90er//cjJ1fXu+42k+lIC/WpDFcVs5AzHXBdrIu6aSayE04GX
qOMuBPsxQz3dTphyQZoQ+HigUK7cOJxNvLwj29/LCBlBTlPiZ7TcyetnZU3hDAn37srLhfrRLo/5
KiTTzmpJUu/awoK5+ukupMkaNwfCbZrBO4QpB6Lm+6q41u4kP+z/qWK0a1KPyMASsPZqWJv8QduY
9nvWLDsu+iSdC/8bBKONZyPdr0Vf0vh5g5GGYozBMvNfBRuaQSb28jvYfKx5nYAFYryUQVqbMBUX
ULBSPPAWlggxSTGYPN6AFdN5FJ2vAR2/iFVCT2/hw+w42Nc6vfGNeuDI3d+v9JKAGxmcqu8z85V1
tdUvWBF8GZSUPLb1GVmSvR5O+NaSEK7QKrrRxdH4McblZ6C/vrDPu9hM27Fkm5beNviDfb7eZ8cu
Eth5B78sPAQybJVcMdiYUEK1hlr/fvTX2LQsHpp9FW7JKZ6tLCKIZ49KDhBek+vgmYeKGUEcNgyT
7SHnBW/wdAunmlMHWObsYrPEiRqHml2zAAq8Ub4PtHPsD20Ti5ulYE0dHoo++Yy7zS4gGU985/Xc
1c7pXSnPVEPX2fH05x45GHbHy7V88/9Q12gaP9nySsymFDYzaeVEF+OR3ahFOAm6aUZkT8z6lzWf
TP4+jWPQlq73jjyc3tt6X4eWoK0Fys/61zHPdIltq/Nwah6Mv4RT1V/Cdv7KqCNtLoNH9AQnOCh7
KgVj+kOBdBVizgzQLodA1R79Ck/ER4B1kAfUiPDNSDzkb3nJTG50o9HE7HnaKhWq4t16KJlM14eN
HDCSRXlFrZKuay5aU5Gl7kjcexvX3pgsgJFIOsche5K/QJ+Hbh5OaISNd+1tqEFo1PQ87TeLPybt
6zpyneZ1tw4RgQyzpURXd98ePBHx/mmzZcHaPPUV1TqVoZdae2i4PTDZsie+FsfaUfQ3n6NeOvlC
eX/MxYo1WFJhUgyh0Sj9W8kRQ1iLSWF++/eazdQnc4e62G2aPbj7dY54IbDU+1X+J4GyApZOBhK6
es5QARbRlTv9nEWS+5ImvOYSJ104GJ5SBlcvEJTu+Z4vOLZrprhe8v6ItKCrEfAa4d161ITpot+1
bO5UdRXq1YcrLAxtqHcxOL0AT+/83Po6WOMW4yABz0wZMsEY0v+t2uF21D58tPKhQTavP/pH+5eH
8r2ORmYWx4/LOVVqEsCZIJDdbNt2vNgFt6naKPrDUhPxyDBY2UHad4stbJa8hpX+ncU6dnx9yb0m
ntHv3giJPFtnbwl0D/8kXbmEJHnkVFIeT1aPey2NDNCvE3XduJjHVMK2wGaZOyjv77MBOSqpQD0P
s7d1rVnPxstjNQGLO2v/MWDEmNVt6ipz6a1W2nPlxm3zQYBOZTayGGa426C0YqWjcXK7t5343w3V
w2dRSiGDFdgx4YQQDRaKktnwe4VHbiSowYcyGqX/1zZGh9dzuW1MKG2MOspmGyk4f+ekfbFcVsVv
2kFWlNyTVjoqL5eHLG9hGceVUqR9g0gxcoxkjs65w1WKUPwegVZhdw3GopuKZlQHaKNFSHVqGTik
pcf4d5KF2imGlt5AIhqadau7KQx4DI7IGecOHo8chnqV2aG3na2o9EPutL5FD9GM7EzSfYE4Q7Hi
0haM1BWBxOtreYG/GLZbZzVQOu4uFKBDaBLwgSwIEaF+R+3sO05oJOzO8MfuYHgg2rX+Iaxfi21q
zVs7fnp82mi1bPLMIdtxj7Lq79SAlf8pwh3BtvdYAdSyN/DBrYtKVyueOnWTJMnX8CbW4ID6BiF7
yalzO+SMyQmpRBPD0C4HHLxudHCxqLHWNIQe/RoajQ8lu4qCV/DgoAVIUXCx1wFEkETsoYSynN8o
f1BT8yO0+pRC3FaW9cm8BjZlBxpE+v1cXJkggE8T20zoHSDPygGdIU1Ib6q5XeTJEpFqrYga1eD/
l9MKN5JCcMnDivp5Fch66zUK6Hu6krMBORL8u8zvmqTNgynC7hi3sDHN7q348nQTCfYyqAvVxi/f
qCfHW4kg3YAYdd+zyuN8T791sNkK002hkz0VMFXJ7077gpn68CTYafrYNrjTTXffWP7j88EgG6Yi
MHdrV+ssqBD86bAdmTFQO2wv/1F+nmyYpmN96dSVjvvZaA33FmH3v/pWlhwGxTuARGnyv+YIcp7G
B/FrY/0ARLCHSqV9Fxhv+/F4KEYoHdHj6p3IAJKXdB3nMFUgZR1cSljVhBdZRhwQuTrJSKUPLZgj
OrRQYOfSym6jGKwoSVUlWNGq0oncoCev7Afpj2qK+kGDCXf0JCQ0D3a4wN9YOWREuVRUBDo5cAAe
88Y9ySO2b0Uam19BSbBr71t7t8ZrYLcWTVPqR+a1QYAKYfbVMdLmzfS24mT0UTcaPMSyJebBPM3d
BYLUR9AAfX++qRGsbJZ+DSP9Pa9Ok3r+XkQ4E6+K+IBQVTrDpeRI2BOE39YUnop1JZNAs4ARmPTU
woX9NhgZCMr+Nqa5JB3JesBgj6JhPV1IDl9JXEARfxW3ZDxvL7Pd7QRWGMXeKpD53enA1C+aNCh9
KggUsN2+WsG4rWWfIwEsxeT3G/uYJpffv+3z5Q/xrggKb3ItmaIW58lS4xC4qkUGECHeQ509pFtV
tyZz5uae7kL6HYuq3IUetfYLw9a07qhgABJjWLWvF0f8vAome3oDtGU8Xols8ato4ePQCpMEEhPD
zD6QVoTj6/R77PzixpF81R7NVgE+ZCjVohUOm2CB1vRf+h0bEpWVIFhQFvd8dJbIac1kFN+dRUaF
M9wezkuEWK5MhiGtzSJfxUiEevSQpeNCsPHK4vwsyxdk4veBNdK2tFCYNJnO7AQ3rRKejRqxFGEA
To+I/AsW8exD9ACqP5BsjDDikfD0vwukgYvPU9KQvAi0dOw+7PUh1NAJZkwstFbmTU3IegQAd3yV
nW8/1SSu4LFl63zio63LpmLhIKvM9pZxQCm1N4mnBRR+4+tjZL26Rb6ORuh5wKBJS+J9J6Ot/NpZ
nXqWQDJqKeG57apI2JzfyApeUBTSOn43yHKmy6BmNjA/mqwi2ij6xsPB3SB+QACEt6n1of0lJXP9
bHDCb+y+QTOw+XTVT2DYyW1kjB4HT7YvWtZT37+4+gqavM3Wj2lHKdwcGLRQOwN2X2gbeRva7/hE
k4LwoLu2EL4WJMPNg/dm+2d3RjLhO28vV3ZP7RQV6PhahXm5q+0h+hP6UHDPKVmomVUSLmtRw6Ps
EAs9Hv6Go65sOV4g2KBTMGdHabKqHcotzUbKq5AMWCZNOhbfWn/apnoGeHGSD70d6YH5P+hHzGPB
E//cHf+1d8cr1II3xycmkUBtx3aGnVOu8P7acdf4VEkTwa2mG1YsdzwMW2lxSKEbFaxIABnvVKXJ
Gtzu1vR4zrEeXkDwwyUvtX1Qpmc9Xx5/6Yjg0Q5osMDg+l78FX67ijWvkC9cz0IFeMlr39WOWRl4
UiwPtSwuTytBVHpxU6CfVX0jhMChtoGqGhBtwU7sZtHGDLL9a2O/I7hx6HT6zkqcxMHGZbWQfAfi
ffKsDOSasb0D9gkw5klypoJwUqGAdplqhoT4mmhqxEMb2N9L9CTNUy0sFEycVcXPIeo30P3cH4qF
MiW1kFW/LJhzO3YyhRkug9nu+odm+XaNG5k9c2oEQxftnkXziV31wHqGd/14HkkLor1gtp9Olhax
Kzva+GL2yRsN9LM3LZBEQdaLPsBV2SQBi/Do0Ix9wRs+4bT26rKw9c6tHgtFxIcrAWf0kASb+DI1
eoVgfTG4eNCxfOp50lrkMtN7j2HML3siu62Bpb8+DZJG7kZu0+mrGwGWzucnSfVPaf2h5D5F5STq
/aKJbbdbjtr9C9uEAYneZNzujuHiGrwOXQ8sM/dM0Ud3F0heR9n43Bs2fcsYZjEa4rSeiURlAA6R
5stHYYRJ8a3uz4dUgAfsOns9ZldsRIgl3YhawHW7PNsVScCCBbXC5h43fqVhaMyMAZKWQSIMgLZn
WpBOb1Yj6AZd2OkqblYwpyWKq4qOLYOAloZVj9Mys85pTZ5cRs1mJiSrr5fO/sJsA3dMVKzHrB6z
loo5ya4apsb0ZP8vHrPY9rz0O8H9PtlTjKVP9COXIQNmDHcCw3ezU4S9n32FECp7ZvC/lV4TSjOt
A8/o57aAnZe8agXMIc5LJWQauPtEndaI01UFtI0/FUMnQdDFpYgOewoThxI3ZBRyimEUHsXffrim
arZikTBtlKGp2iEzaTz/kwrttHFATb/tOe4LHyzxIrkVgJXGJBAgTQdAz4kBzVwpMEwrewPE0c28
scykt8z93nSS0/a4HGs/ZfQNqQwbAF8cg136MAbckQVRBf1exsgj0Jh5by4JhJiNCB08LrZUvxLZ
FoxWjUhrUjR7bRoS7gA1A5my8LldF7fP3NNcaiB8QYhKlyS/VFgBDI9J7pZFHDF5LxOEiGjy2yrk
GpTQGGeQGfEbDNIWaiwBO/SXPg2bJRnzzAJA3SQsMNAoxHr+4Prf2SJXP0qL/4o4KQNJBTpYLTjx
as0v54kks5tKhqS+P8G0y9u3o8V/2KDtkn+3zUIMr8XC1r5pXK9lEfNbRNBu7fL8B2vEjnQhnkG5
y1qsLrTBHR/aKPUuQ5CTWgDGttmiAfPy8aheptcaBhkjZdfP6Y/Xdpfek56wuojJQ2AvPmhiCn5d
YTgFpsopjaLN7fR3/ELLouceF2cral1rTKx/XcwGSLOysmhwbwXkqoGNQsE6oP5fhyEXGWJQv3by
lZVgBKUntGi4iLL+3ndx6vf1GfOPDlKY8xnuwCI/ZD2aDduYREo1cddUjGrObHvd7eL9TUYDtq6V
8br2ffVgnO62X7/tUffYFzn5DsPnYJtwdkF2PdmnlWucK2jgCVMPmXlrUKT4vGWghFdVwy7hf+Jj
Fkz8IbHE9GxpF5Z7lOHTSZAbBkBKMnqYCVmjb/STSpawOsxqddfoaQAp/+4kLeOJHBlui7a0mo3A
9cwK7/8wZqblC/QjhI5Fv0SaJhhXFyJMHjlKUyHn7mXxI++K/b5+akNEmEDad+B+O691+iEkoX6H
rYu6gYv4pcxzMyC+fYZbSCn7mmIcjJlNEnWNeAd5DvWrXznpTZo7K5pBs2Fa8HG4X/grYQ2Bi5Yi
494GWPzsuMsO9NeBkdc4GEsfQYuJOXLYevqewadS3gjCI+c+QUaF0JskQBjK4p2bH/icT9O2PdAx
rAaY6UHAKzjm13tBhkfgwxNSxfoJ2QA8kpH95Dw3H8rb0zVSTjxHoqici9kd2J/4vLf+Y5aUITdM
YuS33JGAz9GFlE1ZoNhXv1k2Vm6jGHB3Ei0AbDS99Bzogioe06/p969LdCJxX05Fv9oYcCqtxnIs
X4vFzFmARzTFXs5/wKayJhshB8LQDuhhMCWMBu3T6ik2XXc+Oc0tRc5OardeJeXWvTv3A7KbrXxb
snR9iQKjEyh+wdsaIZDlrkRHC+zrKBdXyYbjHk/rgP7BMHeNJRhrZSuiKKKJxeC9GAwfY7SqGUPz
yl+EkpmLBMFMojQB1zC+AAhBSRwPTP6ylvfH4DQMjWP92I+d5sGHRC//DYLXnBHpl+SYY/J1NOfJ
EdYLTbiyGgv2ZRMFZS4R4UTWQ69nzl5RQMM18fl6Jmgqp0m23oilyy4CrNMrm2CwV4EZo6MCy6sl
o/hxwt5sWxGw03S++Rn+nB8giEhKS/ixwwYhRlfwlDXAQUGwGvSlNTa9bwLRNKBiXjuspBoPdFRW
ZzaTu/WfScyusPia94boENlBPgTAbgfIfv7RFOuzcELfNHVt3GyYTH5p2apMdwcjAG/AmROooCHO
jTZCq8+eSpeGxQFm188XpUtHBGOnWKZ8sUVuDAn7VI/Nc+20uD+HO/oSE7k9q+1X7tzkJuBAkSc7
TqPwhld5IiGQFhdhuf/2CegahStfzH4l0ex1oIcgaZIha484apZLOOkOuTUg86rMOqW8hUTytIW2
hpjwvlSV7KMKRsjctxMIfn9j9vfHoDvQ4jwaCb3NyLJmBpg6VAqo1sfuryye+OjI+i0/VwIatG8d
UNZ8rj/qIYHcVUKYtuEw31KdB9RxdrQ7lBljC97hVsSIt8H8Z+SKicQBza8w+Kmg1Zgn6Wyuzi3y
dzYAJENn7VoqLGFQOBnft0zA8kx4K7qFpDKTSbIyY+vSfBYSlti5ZhWXJQvFgwciJzh5wwK6rndO
5q3p3GLj6JX7nQWTAc7s/nB4rERBycO6M58mvAk6PtFVnl+ouW6INkKMpzCI52JxSV9eIleQKD6X
UfSN0nAeXaqE7MCh9OtV+5JdgF79qY/IrYzzk3BsdGCcofBs6zKmJJbP9w0ZaD8pSxxFa1zoZmKp
rlvsmxIEeCmEfohKDQU16xFNHQx9KHm1x2XSofxaSCPoKql+iFX2L10tsweZidgT3HmtgHYqae+H
5tjugbFtfGCbhLN9zev7Knn8IzDi1yQxNoUk6ou1/SXXWkGntYapVpy8metztaUray8Zt68+F58W
mtSN1uqlP8377+YPrv7pYhPS9sJaJsAswnxNykI8ZvwTbTWT3nHZCYjMOZyjaGOd3ezpjMoSgedQ
wCTS/qvMLxWxOtvvBff3EaHJIdBVdvjVyyZathoapNrBpdLNVadAaKITxu23KA2CZd0aRBVs5x2B
ljc3N/rtzPJz7aYy4EAIMI7uEpuEwpqhHo8nVy9o3gWwE+gmEcOzQTu/3JNhYo2iGaRtzhFSKlOf
e6MZu9LmG3rSyCaMU2RkiVv/k2G0T0RBE4T05o2MREkQyfIAX6kAJvitsH2JrLoar42qrmysBmo+
twjkdOSlMKZCbgkt2E1cnnTtaK8uxdouvdKMJNy272el5NPdO1pipgBhW5rrX5vwk5+SjrPXDgjb
vkZ4sdPCmtq9qaUBiV00NfF0k79cxlIR2Y57Pm8H7UY+TB3wZumS6meeijJ3VY/a2BantkR07YEt
G8cs+Qhi/qa1YneuMH+4xi4YYI8lMy6Rr2eXCpexeRBXaAk7UulSD6TeMCz2YvK/I08N7dM1ZSGX
1NXm8yma52Xv2AOtvWW4Zm56s5+Q7AsL1x1vl6PUOh9ZL9zfs8DqBz8TNQYMK4Eo42t4Iy8aI58q
7NYKa/MXH/UvoZ3Z7mH0js2QxOWlhyn1FxPh5pKLFBoc0kci0tDNkK8t/ivoQoD4+DWChhZijsSP
ZyF2Pl/2tMpo3dF9P88dcJ3UBhXLWGLwhvWuUSwDlXfaQhPutYAMsmaUxmEY6piTweP2j3NdEeoY
7zQmaymoji6LMEr20NS/fM94xv4KKnCpd/lv1YxOwcYCp08v2IgBnHVYUoPkwfjZh+727Rjb5u9F
sVr+WsCQ341tqk+JIo545Yn93pSiqTzTZ+YD9Of2Va3F3lyC12i731CU78f7beacnMRI+kdmJGeq
VdbI0PY/NlWTBxNykdjeRxvmYnYdCaclOi+7OEd4IkPSa7fVeK3tmvfdoXzXqLGM7BGoisU150ta
ycCV6zR6beifMe2gAGbnfcdWeq5T7HAe/na0djy40p/pnHwtNKOan8zu0HmRhYIUaM73wgwxjUrz
6bzEGNqZH4mMPMTzWy8qVtM45qV+rMrifFUtL9zSXEgwVEx+xlaxhUqK5GBvcBItLl+tJjFooOgi
jZlI5ZdSe0PlF5uiaLnfbvxMXDwOR0ySWRxAQ4Ce4KOHyBxPtVMB47f+bnq7ubePoft3rrliOF0K
+LfrZf61JjXtvNF5++gPAhq8cwPa8x4OWoFt/V1Dr8MoEGNLFnFaY0zB566wv6ii2zrtXuiFYm+Z
KrEAc08Z6W2cVKnvVviq6Oj9reunJLI6BbK8DMnvPN9BfKXleFZXRMhyiuFVgF9fnpiBFrZkUI2c
gNf2ktuAm66uwDyW2VM2kvavig9xE5j4nmxAxsd20YVrpcTzlGrigyTY8D9CG/E8SomlUaSBdWJG
wMZ+iNyFq0+TQM3cpZdHAycwQVOkIHE7SQYbwMvxGm2AjZ5DSJM4WIBGBb8IU+/iM1Bp8fgv2Teu
99F8sqWsNq1jCjXdyizF3pWgPhjGK8lOgMcfoRm5DMF1+396t3m5G1LTKyLZxMYNF6kTIqtiGt7l
HMW3flsZWDBN7XySyJ6GiHGeafYUCnKa/hiZc+G0aL/Sr2tbDW+grEtpyzCWWvooIbzSsk51UgXF
X5bAFo7TxYYYzcgSy2qPgXBPDDlFBeXPQdshdzFdlM60NoGPo6r1zF0VCf58JD46jy645+2CxYYx
0HlI6TYIqV5Ct6BiA/hVEn3qUCt9yocXmZbNZwRhS20Ag6WOgG2wDnEDvupgg9L0dBPoYGCjmMPX
fgEnQI8VpOi+1Qdh7V/hQOnXY03NO3v1S68E4cw91hygKK+G8uytKWO2mqcbsuCfPx7+J/xPBphS
fTv7+XF0KZ9/1zhRMlISLOpdjHsBeBrYUHeLKx/V4pmQUUGfArUBjdv2T3pZ5ll3nFf9zsEGUNhh
lb+5NmJo509oeDMuxojQQqga/4IWiEJ7w+1xXLfSrr77p2VPJQS+uVOcNdpaNQSVLTn3xZ9ovRPk
Bz9nlf9/kVO0dwemc0xYjHC2PkadOEH5OBobvu8n7iBFezstTLmqwUEOyEGrDmH4/P/SE+/H7HYu
XnXpf5b9+jlkQWXe9V79pHikpHxmvm67VPSLL8usqgsQ3S1CkNzEnLBOi7Vz5KaslwyTZDLEpEaC
rw2ryQxa1Hate8JpPvxgoBngWN+McEfr9SxXfU8bko4bZUuDZSLuDXzUhnd1ByhxgvGRixzc6jc3
hjazg+30RavMDVebrN+WTmFDDjWJHXs3brk278DthsUM7fcFqc4sXko/00NchaGLamInFyUrxg+s
mfknUPN+MmYBjSphqrORzMzRWPTunAQf6R8DuGMQVTsy6tCHO/dOJzMuw346+5ChqrZ4zu3RGuKp
m0IRQ4ShyYdrfcRhSAj+9v77zma4PFkj8vN7sHuRRabyVPX7eukavjmGCyZSd3GCO5WgcLLO3Oig
aIU6Lq7BO0Q1tMzygYJCMGFMjyIMNhW+t9atVNJFnzEqqgDih77WQMK2knGfgLBtVJrVRQHI6Daw
i/DrNMKOa46eV278f3Yyb4yTTGLczaPqFElVLDRpIJahRAoRNXM+O8NWyflX2cp+m+BnzzHP9Tka
rbF8PIMrhfDF5hmQnYSsOELYFOvjlHMMj/Wj5CeabJ9ElliFz+R3Q+EKX7MXcSF1cHXRkHbBHJaM
iVkCjIXU3floIVcXJblmuqC5cI2cyJaB7QhBFvVgArtK4kEb98qkViiH5dpD2UYj3Eb9ft5nV9ui
jfF0MiWBPLaqtRqBQ4nJp/a07jbjOxzd0y0SIHXQSvGJQndlF8J91S63mvFNbzf+lhQ5Zjy6dlkU
9SwguOo5Pk/i0ZM8vmr2BrmHDp+7QYwnH2AbUP18zGTRZxBWZSNJWQ05ypgCsU1itwwMny1+Kb+s
1wcgH3q6/8tqpwAPo7PG/360Uk0cgDruSUGUNEbqJDDDE6bFm72IWE+y8W16zmZP71hWVLxscRmU
RKIOEYIJDYkhAch6uH5kKva12l7PLWPzAyQYpJLx8gJG5LXFhQ5YNUcbl4yZ0/lNRcafpcPknEST
/28n3cRV4Puh9CBuI9EtZi+ZSYfasr6dERB+5r1i4qTUL8XTlQXszpVSKJvnsQ6AxQdxSVryyNL3
P0PYrJ7zFDzs9436WNKO0m7kkfuEGt9nZ3AXET1Qj9hdIY3teTS3GmMcGG13NFxdsq0q0M3vNb2q
h/jblo7uAQ2bLZ/Vlrs/2z5812+GrnXNG2DEQnJfG13wFpMjNnmEFxcAEEQocixft+13uiKPrl68
adAsahlwbaAweCriwWLsuCpUim3AU2SUR5MIeV/uGJQkU6svOU8J71jalEL5tqvLkNroZxTXuvoR
PdiL/uSoo+Bka1N8HngjRrfjQZgqaSQepGziKuEldffQvu7dzN/3sphIXX0vAoBb5V6KcRK7UaBX
ovzWC2aHu8MZg24APOcNNPdw9QY7hOuuMQbI2SO1dBgALogbvT66e5iwIr8XgxQM62lQBNxj+XUI
O6uXsBiCZ/dGJzLhzR2SQwpDcKrjsLQvHtEjGPpBoEl6kYpVV4h/EKB6+Tpmo5zKgdcccbS5ok5k
z5022VWbBK0QVH3Nc/5RE38L+Z9rSUxgPeNMof6dqr+QNlRw1qbiGwDoO70ptOP80dBsh12yBtHl
gQRhMYQ+WrkS6PYSURX4vb62lvCC6iNojskNGaMIk4Hc8KbQTBkmCnIo+gxoaIdbqUXWWrbxjdYF
m8MKw9C38LUg+CY3fFncLw3yRNsEH/ieA/lBCti85LsPupV/5BnYb7XtNW159omBBpqClUdfnTjg
T+/7+YrYnhxRtjOAqIKbiTX6p/v6WJdFwXK9dlwgCQWKW/gJ/Y/8NHxgeUvoo7DwkUO+OX6wOCF+
BmRQwNPTXtzhrfibtAhR1EAOk5E0uwQhvVmYzSRvgtx6PtquorB1p40N1r+MrL1ngYaZgY4vdkLu
MPMgEx+92FANuOCYg01QGzahQL/Srj54Dc97DY9DtEAUXkBpdwtqyfDI+glJZjgonXxVTu7XG0k8
0l6cXj3xI7/f7N6BB8hdxIpCMVj84ZaNd7PtgcIiAvdmq4bLh3n37QY7WUOtBVUavsfDly+WHXsA
GZTxc9ukwSkb6fNZmjQpK2yxe0UqABFEDqWbbsGdC6Y6jDdXHjzNx81u6/kDhJfk+YYMjat1FlB4
O7RXrrJsiwGvRiXqwBehFtrVtwxDbyPJjugezswHGQvgIz2QyLe7O//Llx1v+KwsZX9AtkzYE6/k
HfCS7RV6tny0JIUSI1kkLk5U8smHZZWEaOCMkibH0RfLfaNrYbzoCvM8p9u8UV2Rr+3YFx3/G9zh
Wx3/A15OVPjpsqZ1YX/uePcFhQC1rbalxSgcuMx5E3PZzHz9w3ggA4hJiUTjyNVR687chaJpnd8C
MlUc2hEFTK4WhhRMzwa691QxD/2YocYLy3iKVd7HLswSjnMbHd2YE41WM57j0I7dITme1ZLWX711
kRDeVlJn5JySs86l6pvrWf/59WnZGg5JIUtXBREzrP84bIBJkTJxQRJGHElLjoMYG+mOKGcp2CN1
ST3OFOFW8MM9H0khE0RARClADEFfn7dnrOF2ppVk4Ohpa6LyfTL75R3mP4yf9tioOu0XghneOCAj
3rZj5iPckET6PHrroLtRQ9LQcRF6nkzBRTMTzkCiBAaB4hB1iSn34kOPRbpThAn17Tn5Z2FgH8sO
L/DQSyRpJDXn+mqVHt1KnfE74g7CkWJptvGZ4ebYxFlJWtGL1O5q+YS/z7T4smKLQIr6wx3gEFjp
jug0m+XmNlEQDhUaT7apdwoRwTZOm51ZLj3mW0VhsdEaqWvR14Jx+WrRXsCpxmQ/o/0ZdrVv7j8w
LpAL1eQGOPwqnGTDWcFDOI6cC+PUj/PKNsO26CsiNQF1i1VcKLavpV97x93IOb16sesEWg5fPZ3D
SV3FDOwOknZaH9QXovAiPirCc5TbV4j4HaWCgZQJ3BvW5hQ5TK4vKU8oI8HwNWD+l+KBMzrg0xAy
L+iwqkFZFmr6VgMucpb0YHg+PkaFTxnbnqDCdMyslCMrbvxwggkeEU30Hu2ezbu+pyLhh+v07hok
P0T2Nubf37eVNTDbZvhxV49VZh1CfLxuzWLTBikbWZVD3ezAhTh8xkVz+g3Nq5anN9z2BDomGAhY
FJfP5zdU5Dr6hftQSaFFh97XJoMWLcnUj93aC3k1PnBUyc+VVlhM4HtofIovw69qiv4WxfcZujvO
B6IsqbNW9MaU8nndJh0mAEYGslvA1It3TEdvP+omTMjCvNwE0xJkhw7Me0+5+1JJO5B+n33gLt/B
JUol42wHSFWOzupjH2kLqM/5giMST1ECUD+ylJqR0azneBdWGpkMV6TQ4hoQw+SZ86yKqs1SFPoD
nonSw2nLdhLmRKygMklce2HTDF2o10kDaGGYmzVM6qo1Hn1S9h94DLJaxkwY6gNU78nByowuhiZ0
jPXkelPoHgVzsM2YffjUe8STvmrGS6cXOzXjOeUXz1oJxdr/DS1yvpr4UA3yaD6zXz94+a3BG9gq
/gL+UIx5bytBTMGEvR00cSrEjHGv+/gizZGRiMmJG3FbdO4zbcp7l9VSoA/Uk9blnYEz9Uu5q3fe
C6Y908b64ldvNWePYsuCkuqjukdY4hWM2PUdebiYO4noGMCxMNZQuR3WxSvFqiJ98NViV0fKAU0H
QRQfzSEq0N/0lPSNOH8EET5Shtlx8jUrsXbKMNk0OHYJj5wTP9OPKghE0Z2IMK6MVFwdHWMSSP1a
qOPESyxmGeujOtaFTEvAMxZA6mqfR5DDk7IPm/9a0bjhxMgsDEYmiMTH2kWX8jivfW9b0GFmR6oI
nHcnu+79d2mv95guyR9fBXay0DXUJy5zBWdI8g/D5mNkBvdsOdl+O0GH1OKuBOcoN+LCXeMTWPqJ
8PtrK/GRbKw3rgg0Ud5eLHfadnbk30IBmwgwfYLMCTyiO8kVajJDuuZ/uFhngQ6vNiHa9xHTCG6O
gLJfDdu/g7IMSX0UdiDwLPGFU7IG2wL5PI8GmOk5/zc4rVtkM/pDnLBm7DHAGi17GmVKJwiXH1+L
aGH1TOcvR1KDba44uj8oyImEh1GFuORgwWEEM9NYnrL/eiMR7EeGsrBlptQ31VV7r0qOaWikmgI9
HT/pLIosDA5s6JJuxUUtrEghaqKnLD5G0+CtoSh9UQGo+3G2ZPxdB1poQCZE9iEGTgt3CPJJilZK
LMxgHlUMcBH9jHE4h6K4ZsQB4cWPcD8scJjxTvrSGNZiJUv5bf/ieW8IaiwlmcvMA9Ln4yxd5P/S
59EMqv1QdNNqkwoDk9IBJyC3my91mhuMcr66B7sLFXPS/BJFst+icrkFpAvePjJS4wHi3Ou4BdSb
a2ZDYlSXN3MK7l9wm9aFQ2GJ8+5cM0aCSPHERR7CnQDIjkiR3Jj7vEaQlHn9ln1SLPGu1wQUZ2nb
uySX1qSb9M3SJ1O+wsFoYaOKVD6nrdgPbRY1/WNPLiVe/L6ZkGXEW/6ZoxkyqMiZ9KM992tj2Lx0
K+01iqXcawTqAoJlPDsz/s8882zcwsXTYNPUDqPBw0Nr184xA9JGjbzSA6d5WXRw1CWiBvLSd8yx
tsiX9WTITQe63IGlm6HTUZe1fZFQL2NXPFCn+bE1bEqUdT4KVuBoAbe9/IGw7f7UNOmZhGxGfvII
+8jMb5Xx0xVY0sbPsLtHZZTJHBhO9eyHQ+YX9OYSduvi3X+jSXNfMvBbPb63EKx5k4vdLKITJZ6k
cfj+wRYrHCxcg4SS27BGfONY2WwYA6VgdWFJbYJo9tfndJDmw+Q/ETG4Az6RdiX2RTLRisRDoq48
cJNA82ozqWRZpEV65N8QcUdHKEAQWeO8GDb/dCGk14mNn/0E/KFQuzvUIjrtrrYVDTygZ5k4ctdx
Z+homEb6SVD5aVVObbpuILo29GbzZBf4IyVOaDw3KKEvvh/B5YYN0fClBT+5pU9E4reXRS5j320R
S5Zg9RfZtdDYK6LFd5b6mR7T2djIwX5NWYPX4uqdgH2hhUEJ1N1Z9qb3BbmoxOdvpTpf3gaazqZU
Ds/XKhNBZZnxTjydoZL/qlWcxXbWX6fHXu9bHsoq/46pnP8Y2UG8R91YbtdKUw+HmvRc42KhmGsQ
betjWlCSbQaGa5Ha4ha1sPauBWqNS7hxe8hTo6jvn+FzRYS7eqNU0XDPL+5tOOvMfNJEJRVxmTVA
5UnyZbLrEzPDK9R8KpM++s3Av+e+mrmJi4sqQ1N9dsNCwry1hJbMHpUolF3BsNbQLnEYCSlevLO8
z8l/L7S0p6M9LPfHuv0d5ixCMcwYDGtbkmCQYD0NxISWTwTtBILbb0NAt+opbOOQwVFYly001bRS
GWwcA6qfRAZZSHMWtEcUIVDmNNAgSgjMqGoGi1watZhtAEi714W6lduYVFwBj2/U8qUjndJcUuW2
/7Zz5r6L7qdq3B0mnkAdnzjJsOcAUQwERH6yGd8b3zcbNFyVsU9eZLlCmaWF8q5WO/eA0ILIbRRI
HE5f4aY0BArxyOk+f+IONsYuJtU05e2stYAIpU1m3fNoyPPMvLXIELj7O3RBBGg2ljVLv7IsU3Uz
JF96mT2v8yxTMt8kgsgcdr0DxboW19/GE8f727+fR7kb3fMz0FaG5hBzaTHrSCExIQ3aJ2E1Ds9d
ONsKNWnAB7PzwhlSsAzXtbO/ND9qbln6OpkGQ9hJcm1h0omLng43tdrnSxkWICiugtdTAr02T/wE
CJlCGhPeYw8EHoR805y2uhOFu/AH6jEFmEEWJ/uquTrirYIb3j6y8h8DPjRrnorJIx6ypGmlW8+i
epDpFoBae3rfY/2T3BqmCODPPwh7Lxl+VqWkSLaVHYmrRC+KTdpXBxlZaaRdaaZN+g9dZIAZzZa1
b3n5OJ5GU5GxVoPYlAEOmw7OqZQQhlg0n9KZVPsrL5xqeaqEHqYU0Q9YGj+oZ7Z2XLD3MbJZtyeL
5+Dc0aPpUZpuACha768jlf3+n3DucQIOoVCoEzn7LDfi+tWH5IvHUaNWueqSGjZovJnCxmSmeDAY
hQUOPBve/3/WpFiQD1PUPip5iV1WAaHGEKhPzxip2kpkq+fpXZSGmu8dfpPXIh/B0hnayk2VNddH
EphDjvCJcnOt9OwGNOqtorxU/RWjbl9iPd4/iIraOFG45fBRUMDjkk1n08jDQUY8/P2whGc0wPBL
WsF4RoL4pD6Z5GRI+l6rZd3zFOrN/dNt4Df1ahxyP8MlpOfosSyXNICbBx5L6xxQ/6rqnmB3eVWg
okuYYLGWEHO61xKXb9DP0CGqbATBvbURQ2SUJGvroQF2G2vMFvtxtEBdkSkdc+kcXgDNbh7assK5
o+EtFayPxr/QoKCuOrA10z4zbwgyc05xSUQPOTD10L+WG4iFz2hQJuUzCIxrV7TbYpYLX6WIr2aa
K5cYVzXXsb9lUKUyej9US6eGR2J0Krf6p+MdL570mUsVywcU+yYAus2nB+I/iWBcOlo5kfgQ2CdB
+w/LSkYp7PcXtltyTltfHWSKYbjSrSduZ+nNwzdX5BP9fH4Zsb4B13UdefHglvcKsOcmuUKQNZl5
hdk9HgojSxKUwR6Q/KapTCZ/GPip7h2kjUCDb8RV0LF/gxJQuOTPEgHfS9O0MhRbn3YXOc7L6mFG
7Sjn4wOzh7/Y1h8OgqEvRuirZwEYTEEzkyJ/xfAiT8ShT7oluJDkxN2RS/FSRYaLQsHdpvneNCyn
+dT8FHhoubA+sNa6A8iKIKnpQBTXQnnNx1d56WuV2UFIomN8XdoheiQLRoH33/jt/mtEEzAH+iif
nBKyGkgznommqTR1aFe9os+DjtMSNSVrQnvGE2KEk6vmiw6UC3V2AHOSXWfizinSLWlwC8rJmhmu
MrXJHxws4t21lBXmErskpEZdBNrzJ6lobIXL+DQ+B9H9lMwkkgU0/9Zjc/o0CF+hMvQOlFhU7avm
LwGue+DRTCZxicjp8MxMxPW19fcuxpyAJNeyecgCaU6FlueBG0yXlf7x0fYfXaA+2sCvlSBR3nJA
1LSahJT636DjuJgXyspkTkyybdLTzgwJUD6lN3Gf7y+qPKLxDscSYu64VN23ekkDVU7GppPypuv1
SxP61MoFUZOjy4G4iFAdAIKLWHgGux0/nR5MAXuGCz9o1X053eMXC3bdAC4Vh14mjS3da7tn57k/
trJ+XaU7EdfFVHov3dlkXlJmceTNSnwZGMmNZlB20UfDLCvOjp1+BTGzOFhaenW6X4HqbAP6qmKc
EJHGNSIqkh5L3I00gthLtyV0/6PsYnJJr+cVcwHnoCARsW8NaZnRE7fY8bzENMe1X0zPdtY+Zm0t
FYbahSal//l7v7i3mvmQZDZdRXaadBl9WBhLeDN5RFmPy0pM22NuZ0Zg7Rw5odCOJB1QLFF3lz7i
s9uLaekGMwKiHNqZylxA1vQNnP8lXwhzy+HhCvGZvgTVREIGlUafTlAfBvf9cgIgu/6ijqYGL5l7
rfxKrGg6Fe7VuGqw7kfL5SZCH8ze9GRqSsH6n2RWnl3qUanlFfavROFaU9oRwOCNrax40JQbiQ3Z
r//zvcY/YcO4PDVnt8DAGImO6Soflw9zhHN22NnQifiZaH8QIBXSCOTzupZVoTdVMLWlNUX+ySlf
u9kYt0TgBi73/34MA1UV+MJ/ua8wq5hYVcybt6raJQfT5uP/w6aXMNeH3DuRSj5xU1Sk5WeBiIt8
54PCnMWd1YKyzV4di+U17MZ+hKJDEj8hrl41HJNfbpknv09uoKhGf0/vWoclD2vYFJgPFA2xcT00
vTgc+GnDOpYpYqSZ13zpPGxpziaegjZnJOHLdC5CHK6PBa+Rf6Qg2Y7ov54aLCgbAf0G+2+UDNNd
9XIFCrY7QQs3aYt7KShfCPbLjS8nFK8jwT3PApnfJfj3NfGcuZY6Ns0Y/PPA9E3O7AQ5tfUmnh7e
0xAmWqU/9VjUBVf0jsFv3QAPuiyCsElRJ5FRdlN3Pzoctzc3BBbf5R/5Np+uxS22cq7zEjUIqTfo
BDPEjxhbqWaEsjcJjCeReV9kjwEXFvJpV5htZTiYO+DNkio8smOB5hXDKljMvL2DXt7V6A4TfdRk
wjzvToQ3R4WpL4Ida359Hyt7gyG13ZVYI7sA7avB8O1yiaAmnXwT9OxGJ/2Sloc+S+20LVM622PG
pfz2XVGzD72M404JLkZ+NkvFvp9CaXGQ4yFI4NE1xqfN7UvP6LUFYPAyvoBCRB6lQ5vuqvHJO3gE
q56JL3b11XgOYvANsstx1a9dlcWmByPKyayWjokocP5nburO1y9P5AvY9uBIkttM/GAWRAv4B7pT
J+qwmJALo1eU6LzGCDOffgaiPXZ5GckM+YjOJQO2LlCLiEgEp41DcavcsBqJvP4+esN4Hvp3sorG
MVwj5BGLWu1P82Xg5giwama969lGPIPFdvHyBizFyImk8qzgMpSGYfHx8dvyzHDLyLKuNeoQJG6R
6yiUsOO2i/O39/hE+lDZV/bhPZQvThEKByTDSE+EbgNXV+hJuOrMmIn7cSHX6MjwRz+Un/mrMXno
1ipIk86X1mORDOZ9An9R6HuHKWKBx4hz/bzrm04uxMCNftmd7wnbe8MNIRxIM2Kzhn+/gt6eMiFN
kUMalfx7lIP398fc12g61yPS7nZxzpsNCYlUg9UJ+qA1sbCDWOLcQxAAnZE+ExmjwqdmDh2AzABa
CV4KUbsCeqXkCdZQRkqdNdFb+h66RB/aUgMAU99LBfP2e1OLGBbRS/pDF/LP7hf5nVVGmn+YgcQJ
hjsEaafsfjxeQj3vPSMXoOU1Y7xs27SFnA3YTkXVLnZbCVrHYDuUE/TB62/7F+Qj8Qcu1n64GYVY
MzCVZzZP4tFHloGx6eyFPSqFdH0L/cSoae0yfML1WXBgj8+xvabC6UoNFd2VqBjejNFBImc+GEvo
cYhtvNv6qTMKFqmt4gI6iDFRMYqzz4uHrjJ+yd/GUP1BfaG/P6aiDUPNqSHO1+NvavNdatl+htAw
dVMBPWMmk+DmW1Pl+duHv5NaPNE319JdVCnoE0v1+RlHli16sSBU4oW93kmXbPAjutDIZtL4gJwF
WzNO2MK+rnfF4WDcu8bGSUs0maKUtamqoLL0kePx2C0tviu+a88j9mzaxMq7tRGwVft064hUXnkl
YqVnxw/m4hW/wfomkxeiKouchyQysPjdJePDRj5Xl0fouqwCanwiN0BNO2CVRyZVt4fjgKHYrHJG
YWEFm8hmXaXCj+yU1pS9f2Mq2jWcfpG1t/BarUGbhfrrhvgC4VJosvx1CoXIejBiUcigyHocPVl6
mcbbsDNE+EKK9m+KgQipgYIRcML/cKPnvTM9nhg64ZahxiM4HxcOXQwhlUjGQYns2uBQPQQ5+dKI
LO92yR9oOVK/mee3ViUx74D5ueM6tuTUDAkVC5Cr4DqF/yslwuDnx9GgxlojUbGtfISJBrES1Dh+
3H/E7dPj/qcStyiUAIGgGoB+iw1nl4jiyhMEqMHw5xzIWlk8S3RdCWkwEkgU6/p1M70tI3OyKzyb
TIYLk5r8INIkJxqfPHEpYreQWnKAAlKaaKhgbK5qFuxyPpiiGP6w0x2Yrpy8c5eyfqDBbHT27Kk3
RQapuIbJNFQ1fIsXallo1+y2Jj/NW0AAcBNW5fv/l7r+3HVoL1f75Cln/nGvbrACCmaXxe2pQp6v
VzMKkNEnk7QNSfQOdyBPYp1Q8mRnG0YgTrCSmotq0OWkUXqVjIPyeF/8dWRUh3wh5eLSX/M6jkCu
KxagXwcN9KuVesVDrb7T/z7axHAKgslSgVoIwrGzv1MOewreBgsUil8+rjFxSumMUQMTnvMxXPpN
AruxfQ8hofvWEwECSRsDalpIbZVv7FZohWesWT56Q1QBr62CLDvVzVqpc+3+sK3pw7Gym+nX/Q16
jxpTpshKRe3te8Mn/zPA+jldDPXyDioo9UCtmopthZJO6eeaEUKceLk3LK0+SU3Te0ud8LdnJt3s
EkasGwMACHABFsdxJ6vDLzcd7M6TJwSLwwR2YbOTOQHjEQobWjDXFtPX5yqXgl98aI+Tv1CovsCo
CV4NDtlfY1t/hS/IRTaXZf/jw4xzTkM8jcjGuRuku9mUmdYd6dXogTv2dvXWV/ce7RvP3kHkM1us
NHCkNVW0x9/binb3HXtOB3kprfnZgC1RNbKKrz1hSD7fKenwF/FVAvmQOWjJ0Z49QaL3qrr1V5z1
ncEM9l3y3dJ14FOfXDNUXxcPz6ILtxWw298+4KwPz8VOTfnsJYYBAbyPYrKh0Ql1pE/4PvJWryHb
BzHG2QDZNAII7oFSNFGzjCKxaGVQUtMejmazBS4cEXj/bswgavOrchYuok7nYWBNQ6pjOwIiXZZG
GLxQzkv96CqBUFxSuwFoGCTNcKhFczpV2OVdJQ5pdrPj21x0JwSsxT4tC5EBKDlJgB8rcbWNxJFx
w48YkndMlhYWx2uNx5nITZJ5FP/yDxscAYFwBqTCu4u5zpqRVVGE3krfrlY/gPvt289M/uO+ToUc
z1oo4UBnpJMPzp/sWcSiqTTiM5Cotmx9DVL0izucoymo2VY/tLfWESZ29fubjylweJ/jEGSWS9sw
LbIvoi1DNAI1AiMMhSRD2MYva9pb1SwJQUBv4sIB0K7hK8p8MTXbch/+8hHuk7qambA5XOet767V
MiarRBcdrfmau7K8qlYwXfl6jK/JfCJhq4HgznDNtccdXn52unon8HQGjpu7q1VV46ir2XU0CpPn
vdwI5O9x8agQBjU/AUSA28/Ed9Whhy2huJp2X+3ptWjFtYrDCaTSMjkCA1LJ0PmCuzYxberSYhbB
Xrt5RABMZqpWu2z0MAAWggqk/qQLIh2d9rCeaHdnIpNjPRc12IC6umWnJ9gmitQJYvDyfmZr5dte
F9PMtyU8mr1GH41I6zBKeG/0PWDH3rSDqT6rfN5H7A8lWbP6O+0f3J7/H9EmVJoriwhHdHcbAR7M
kivwNcQx12HCruwmd/ZEoIe6jTkgcrW2/ZpYWBBtcIzopkBV0E2IPduCgdYD5mrGTZc9OyLo9nlZ
PSxd0I3ecJiVqQB2Mlrx2UldC1kitv4MF9Q8LN/2DWpnhxsoO+qS9Je0ozt1jExQG0/QpIhkwx7V
fT+W2S0MpwSZpuuYDLuKW7+CZo8ZgjLwSPjplkfyl8Uwvavs8+mhMKnWx5dOHOqsCd3h8/BFJedw
WHkRXyh9D86i4MeRKXhEoGV/1+JIciyb3v6wDfM7B0pnRKGAt1LqDIgZB0TLSKdjeZZ4J/ZGOArj
xitOiRf+bmj01Fow8ydlukdgaLkL/dswnuoWOYAxdkgYmw3sGbltdSFWn1P6XGcGXzTNjZ83u626
R27BJ7XUnrFPRFk2sqsf251N5dyY+0M7Sk9k0wxWtGSzhD9Fpwlqf05BLhAznNGhgIJiE0/twQDr
zlShdCT2k374rsnrrM5JdxtKIaPs51Bd5Co3XBQW98jbLGLkLuWaSQHNPDlFPcm/fBJdvdK68ahz
DC9CCIeMPNPkMRi3v0md9IQDehknMrw+uX7aDikYvutjgOvRCmfwGc13byqdMolxdgsB7pcowviA
36yBvSZ4EEKy99eVtiRw5IYKTd++mYw4jG3FvrVPYY4Z7Z4UAyAq5Zl9RbUC2uDqDSrPKDDbvuvt
aT4337oT/WIC6C2rv3V9im/C+zX5Qc3pkro9RtsZb0Kuzon6EoRwPNOGbS+Co9X6Rg4TCoJ1OZFG
NEtzyvZwvb5Bl/x/tiJxIukKNwYv0UCdtU9SZz5JFgCnHnEbJkNQHtFgqUUQm5ZONz7MpBXVOBm5
hJ9HewdHZ2CbsVicAcjuR+cGOcgj+y/FX5D1MMlvKQ+XmOWCVILUYQus8j2q/36J5TxSSdm8qjo5
yEzpwz7VYW2G0mrBr1DIZZfx41P7ouWqeWxdGkcpTtZQQ2o8bmKvLwZ8xEz6rME0OtaqaWsqcwlS
JodG0Gtn415+3PdY+9W9adQWsqLtLR//++O1y+oxm78oVRutTi7IxZnHUMouPQ4jrqR+ePwpvKP/
CLs4SOXE093NgXA7SvS+DqpIUhLfeg4eKYNkL+z8Kn/kED2a6ioOiIGVcDw7HbySw9A73tXjhtwL
HlLQUMmYCi948bjmRuGQexDnW5Dh/HIzvIYG34O6Kz7wOC/XvEqQ02LN/EoXPotn11Kyusighs+M
lP+I77ER6sw5SiDTK3NU5TKMdxKW7t7sFyxrGORKb4jquI0/g8S7rwBTcLS2IVkMWICBkyycRfsj
ZnKhXHIq2tk2nrilwNKwDv/5XvRRNVyZZ91CrHVq3/a6PN04/ML8CiREMPYQ3MC1SpSXiOV5tUMB
5mRo6ayHCFWhEy6K/HXfBu1O2hSkr4cMFdxt5d4dloLoAnEQADGs73S3LJJolm5hes/jV8FDITcr
fgsOub7ddltvpKfbMQVY2sKfwt/xP9W8zeSeQsABY+nwKb/7WRd3FyVY5i8hvsDgvC13MklbZhp7
AQTYFOClrgGqyOWkoTzgp601CrV+elr0fXZeZAKGWZ2VbNvYevpijDRGshQC/WP234jvXW3wmpK4
6nuRVMMUJ1Uh2vZoJlGrv8ePkD61ZjivxcxW0q7bu1McIoSpvery+ZvE467tlhRCA2I9xdpihy0s
iL/+82fwC+tuWJOJnHrzS3+GIn2s+gm96kNDDYdYDLQld77cksE9R7ouY0BVDrfCSiTMr+YuhEB2
o8p7DEWXryeyM7slWuswJ06dp+vEyLRpXFBXnzGswFp/cV5s5Y97gsXlxERZFUoNPGpNAXtD7Pwa
F8SZCe1pihETWNGgWi1Ulz8fUDTDGQx8T8pf4po4mkbv+3lrP7w20mSlhZ4QvR/i73Ql8/f14WWK
8Ga2fsYHm+YpTtrES84utsC6pMbA4xLWs+e47s1obE7ByHcgrH9Xep5nCurQ3o9poh2dzp3UszRs
USvM/bCr9/i65fQfSpFVWP3UZWFhPb9uQ9gw7NCVnrC/0sa9pCt7YM0uECbKs/WegRxv68pM9j/Y
jWizAxRimA2yZ2zvbT+ut2I9JwAc49Etkx1Qql2PRGBBWBl7BH8MgZVfM0nOyNX9YrwhbpJKxvIJ
ui27GsAnYfTlpRIkdnqp69MK1txKsYZNsL/uIyqEBRvT7mNqdsM8/oKwRKpvkyetF6MAloLryDeJ
+B4DCYVVKOy7U6qJAXlHw/f51+0IzjsGFeGKz2SZd/mK7tdbrp//l0Qn7mwUPbbGetHCeBRrMJDN
lP9m3JnaIHlyLt+yHCegmP+QJjZSvHgHfkdGro7I9ckF+Gu6OT3gCuwzYVgpE9mK9s7GqrNFuk3K
3YW9wYmz8elS+KKolVuahKFLvpft7I4lPeL6w04Jork/d65YgYnFnAA7VMXE2DfmBViPZzlNN66g
PXLHxchLFQPyiLKjgDEFwZwIUSEK6d1KdRXO9hRvz/u4inpjQ28iRPliDTIomU3gh3msjA3z13WF
gcuVPY2cYJR094vhrBXDyLhzNuVdE5LfVwhZ/bP0kQRRvo21ntFe9c0RMO2sB3Qzlv9rCVI6vZR2
O/7WeeV0qewWBqgDpi5O6frEHBYdD2Uwom35hIL2k7+U71626oZAB/yFquBNnhY1j5pg5qQ/4OVR
2vPt/tfVfwxhfAyzrmZ0bcsJf8cnNmGb6nyJQ1YpHMOA+P1tj6Gt236tbJOGj8eW8zxKuNujzlkP
U4hhWnOln7q1zTxIh9b94V+VnZ0enI7GnaUcjbsFaZBXAhhxHHGt8CUAFDbR//zrb9sBLM7gU31D
Ys7jhH87O69IYRla0WWCFak0AO0mbn29HPuDD+kZER+lSfLvuKDyx7x1Z5qG/mHOzeItpAKGCof+
Vyu95ZNl9m5YX3vGSA1h7CvqCxB0dB5Epa6ivEX2YxPsiLO9pja1IWnFFfnmgPkubFP+tHapJAx4
ogUrR8BaHTTDg4sIgyAoj6Jxfl7ZUFF9DFhLabaxgzymlkbp/u7LDMWuOUvun2e0ULv6raVlcotv
t5ol4SRKrlDk+plqLMoOSKIWskOf+cwZ+in1ONxpiiItcaHeCudBvsqzGOJBsPhYUnoEDoF4/N1F
GzzpEtONqL36Zv9euBpVj8jquStdl0Wjjyaw03zLnyxImgWtylELBy13ZbzHwSA7QvOCuVq2C9wc
3qIYDssbdS9arLWo847eL/9X3pWDjWlhHweRxBg0biMuQuCB1UqynqNAuwXbXiuR7L0CxKqYzuC9
jSbw6Wk6arRS390q/RWiCKKUhP0Ij2Fms25WB1lWVG0MCYmoE57giLNg0+17ZqHNng9V3Pzm40SK
8U2X8IcBNT6YExX7gmLqmJr2mpXZlUQIqQ+XKpDRQWME73bDgASIv5qJZdqhgbJ5ApjLZsbkv8+r
39P4t+Ycj3iMu/7U7W3+cDKLRuJthUJeowXaFtIRPdAUfEhJFkF57R9cg7MrMm3T80fa+qICv3C7
quzjPPGUSlpgnu82cx9axdKNP4xiAiD+NVDvHVfWmbiIxQr9aZqLaQEvxrxLOFvnPLUfn/v1Npe4
IgKa12syWHx7dTq/ptuIWohj0HU04dimBdTAnGn7/V6YSaS/TDplXpVAV1TvbFutfN529MB6wBio
o1eodFBLjg+b9RlgGbNCABaLjW9R4G753108Oe+WHa/MgI5lFH+Roj3MDD841IFYxSY/zdFW+vU1
znmbHvSMVsOhwzMHUh+/PBEerWQaN4Zg68gPArikx3GbXnCMlOw6HMY5dbb3gk48jf05y0IoVo4J
ExJ/BfOuAsZeF/1q2ozBCKvwsFnTilNrHYUrQsHrmKzdtPnyD8dSiYzXlwwaXLJu73+J2JSMOZGh
/OT+6T4CjXY270jDeLogidWeAZuCMMYz+HBFuNR1oRku0gIfVIK6atCOTEL8zCb/nyrkFvjxjQz5
XkKumoK1zr9Idf7Z9CraX46YAOXNeSTK6ku+zfML7DLUGRdrt6Np09EX2i30ykTqFOkd+oQrvflv
bNh47RfzNpSBy8DktszTd9AOHEbQN/nKgbnLeooOF1M6sYSCKw23GycX4UisTWz3gokaK3SDWMtP
3Bkjfn8eRqpniSPuFwlx8t40vJTFIC0UzvGo9Wa6V8vfCY+PdxkQik5nseeyHEgb/v4n8OBciMdo
l14bImESclTNdQPa4yAZOXZE7TPpTsNFnwjrqvPT4Ne4+Cyyr4OOFQo+Zv/48Lq43drwBIIlhSXs
GZ8UcM+SDv9DaXLJpYnKfpXm2u355u72k83w7uYEYpeDtjSgG7BnDVAmrkUYw0TQymCju0rn2l2+
x5amfKAANZL+xuJrMeWEq9/6HuJMwUDUE2XHmtUya62nQ2fnAt9iXdS4at4RFV7D6BBd5JqD4F/0
dACcvlyNiKQkPmF67HaaBY3krvpa7omF3CW6GnrvLm3P4nWdfv1pgyrDCGQYHVwQh0d6+KiFjldD
s1Dxa8TCVJqTIhJUv6SDXvnV+p7wQ1L85ctwCJw46+UNH9Qagar2yNVMoKROlYlmQ7RAzGY6oE7B
/s5L8+vWRAXHy2ZdkPNOvzGHeRgkosvxudUvpDuYDCsyJrQUFeEXUOnzutgCbD2xHk92dxjQXnKC
88KwgfXIi9fiKtOZp5Lre2+f95AptC2nmXI7BR9IlRmNZ1dw49DBiJ5ymg0tW8OzAKiHsHn/LJpI
oavs3GX4g8ICjwTR9Q49y6Z093Z7GmFmoZmk7lF01PRtMT5Zf9h9Fprq/Zdbek0cgMXJJaWGg8MX
NbIoDTsEmVDh4Us2Er4HE4kyTXxPvzEloo/qqUjuEOCy5YgG4YisEXZIsbw/sAI5Ewfo7n+Xs6lE
Oz7RbPURQcqRVo0axAkTT5udEGQUzd8/3SxNt3zR4SOAeWnEJolzAHL2vCCcZlytfZaGu4amBlss
GYCxO+YMRjLEii6Y/K7JEe4NE0zP7V0yyhMKkVVf+nBvWv7fif2lQl0sSAbf+0ENEvcL4jaYXWut
UKiCzniqJq22c4nojnw/xTx8c6k5f1ddZYf7KrP3AxfRNHAhDzD6yGUgTruPQTnhR+jS8elesfZW
xHGSLuM1Ts0bRtk6QSTY2kQmGGmjcdX1mLIEEC9c5MVyfBHLWw9NGmwqhE8RvJHY0GdAee2Ww07a
2cZpNQmMD+Pp5iXsPRLxIc4qicGITDO62HyWLgJrRDb+xEeuvLJVtkCVo9xCyoGdnq8DxdNtsqjJ
16n4CdLbXt/kxmsekAL4zW0x+VWc7lY9h9r9ADwrvRWcZSVJOq/bjDC7K71GunpBNd6QOFfvJtQ6
Mbm805HTEDkNHyTtcuHtTGtDAxFKzhKbMm+KsllRJ2zMNmSIgKzCjsVAiaiI1v1+9o0IlSgcGP1n
AB88x+BIvercB9SGtbnTHTIhVrpCatNhSE4+48pJxkoWWN5yIHDuEOaI/VRLC7CJdE0VhOw+SUkf
NSP2+eAqBQoVHMp8ZyYkKrEhkY1dEamjKlDAa3D/FCl5AvA4jABUO89BmSYOpWRfoo25hq/gMdty
ubuPZWYBSJ617h8o0aWPy3fF1lcMu4zdvJlJYMgpclZ6GHwh+9hcVkLbMRNKu5y9xbKfPj4GAE2R
Y6lbeKCs59Iwe6FOrCaWs43Xw3La/bFsMseoWAaqj+FZSONo3ayMcxH3nLtpeK03rjjUYnwvuVOe
guIaU1sNLCiA1l0Yxfd2auWLJT8G4/azJ+od4UytUvGQGerjTwvnk3qwipAkK7oSaGHnkKt6OGb7
eoS4a+qNNuwaIzSLMvlUNvggxbub3wJUBWrd+Bz/ZTgWjdw3AwTzLWUSdnCS3Ue5zqFc2TWSEUfb
XwlEV+dPrjv8BWXrvfcFENKpJqmhIgvwxi7cqBXkONqnOxIHnkkgA+oaAOI/o3Bhvg39dWm0i9xC
+MdwnVrDLrFyVNbslJBGJJIZZREO3JKC+1/V2OrhiV2PEAWP8oaYMRcWK2G9nxjiB6cJPEXqIpwk
n7PWbQrLDUsmFFMzJVA+Og7c1DApMty2wlK6jsnf+m1TCAl3uQORKni6tY24zTZ2QCNsv3DKeMBj
zHmjVHKq5iHtCH0EeuIAt3xvrp1cZBk7ScGoEAndtod9Haakvy69n1ISQXDnQH4jXcIW1Ku1Xgpb
fqPi14PSxTC8LEATkj4F39pq0oH5fwgPcuiDNqdUljWtWvsbsnsZ0/zucSf6WgSn9hZkXTxSb7tF
hIcBoaJGbI0BwpmBRHpf+Drct5Pd8L/ddpJTKdETp7rnQ1C26rcS+fFy2SM2t1+GX/i+NXtlFsyN
2ZFAqpxtuwCiYdwFcOdR7kTzCJ8cNRoiFcuoYdsvIFsbZqE21k5eMnBrKTOm1JIsaf1UOzjCSMY0
RRgNP5Q3KxgEDDmotuBsIngVrAW8OSl5KhBK5X+QTn8yEMuXOsvrizuG5JN2ezu5npOBV+2uWtr5
98s4ICzaRSEl8C3qWNyd4nJYPZUsueJRmdU/sUQgRo+1Zc4wQYMQnQCNP3aksbgv+0eDdhRNyN2F
2eof+7aKKMrGG+/gYDobHYZ/eMGcwUpaqfPMb3BqAwONHgb+jt98rV3roVRwa4ikoihr3p1XmyIc
qUDw5/OS+UwMHUwDdf8wStK5dSXusjAkWgBI0NZS8gAy8FfxKuirTgDnH3n3sdAO9rrGDQBIxs1z
/8Ot8B8vavIzMuXUps4FialxXfaK+uN0sN+b8WAC6hSrfU3w5+cb/9/xQ8nhK2sNq/R3STWPOGs7
ka/25Iv816DYKVRjbQ4vZIrcPHcNAe+goSIcFlJ+6hhRnSGUrr1+5oxC1gSyYtVeX9FlidKJ6E7Q
2MAF+11XDvxXBEMc69RXrn3oDoKEtjtI6cANeozup5THxKkpBrBS2KGJHRoaVDgpWRX9Rm/XnIm1
j/aENGpRX/1f6pnWK4Yz2dd6006vwtJXeNkWINNeOO9BYYHczumRaf480W8UcCR+bCo5iPcfPtwX
dCvWGGX9XsXW/UX95ic73u+XiqjdN7PNBxKRM/bKUIV2VhCtFGmwKdoKyyr/H3DwhGIuUyCC1g+i
iBAPHeaQeWKGKDBJsWzj3XJr5OY30pH2FYp4WfdcxXelUI9WXSVwbAYQGGYwxOgAWgGV9iKwK/rs
Avuv675smL03pecSk0ZoKBwfYLoGupKKio8F86lSqjSzgX7mmPtFu2iLekZbzOeTlQLI68rQAxXn
HflTSbTqIfXk4eWU9pfQLQSPh4EwWjGrQiMi+ur2WoOsPxDm7nqMZPF/7VPxQjpmK4qyN+qkI0o0
b4HTUp4Ybf8ykFbL/YRoFkOJMyZeVXGBP7qT89fxpdLewVpz5V83yV6o7rHCdaEA2vru4OF9Secf
quqmWr9+ih8lryky7624pTfio1qNoJ98ZpFxo3uZmZFvX35W4CEfkU0XqE7DfyaCu9dlQN18jf2X
9hl0WwP0CKWbSgZRNU/Ck5Y308y1dtA27re+x7XJjhKxM+UKUWawmcbMP7ss5SInT4Jk3UWa5NnC
wEKVT6HsHvdt3PdioJABpN7octJZZ8oqx2/flnP2ZEUSV5cay4bs+aZivQ0QRVYhEpkaceKA4xii
/zjy4tcyIV1o7M9m5nH0ib1gxNc7ep185tTTKN1NTH17coCOP9I9TAAzE3ehJBC3HIebYKeIqYYA
QmU622v1dAQY8ojVyDLlCk7+qg2A/DzL3JypThIqn1iVXDogj/srnlegWuE1FibFaVhgiVRA1evU
XB5zJHu6riC9bsVlJyZ90qADiTsaqqjs4774cH9uR1DjmFLMSrk/EY9NjAp+vLTbKtcrRIohJaJf
qrPIO9MMGTYN/Od0oLCOfjI+cqjP7Z9qjHPg7TpBXGE6Em3BOT7WwAg4lKl+1eDkiXkVvnt6j5/D
xg2hLh3ygUyMWrBUixzwA6/6ZgKdRuCIASgfv0bwKSavPUCgPVtU1XRHYBTn3ks6ggHntIiUIbrY
kUo4Hmk6lCRbROnnxY17tvRGunn6lgmfANbBm2Ddp1QPTYbssJK9QgDFdGO4FeJQBRKwevY5veKY
sCgRC1HebFGVLOt+XU0Q3PzULw2WkMEZI+n/rmNkAkevyw+CHlY2AlnZeRqG/m8EQgzVPEFbHBMY
6vmZoHSkF5w2UBDZCC+s7Fmbu6k5V5JdW6YTfXJHOMxqyERVh31WU0p5EMHa9485vog53QnwPBli
BWxUxqs1NTZ9yC0DQckiKPgwT7/ZLQ78XoCyCq9kmIAEOSREsBm5yYhL/7MscpdC1KvuvqEiyk/b
OpwLG79jPW44T2sM84iOPcGsJApgIJx9FU1jHj2rV7yq4BKLSe/91ZnN4WIvY3lmCETPwkic2kJt
vRhBQNC7HVWtbBkPfL+Ca5OJhHKhDSyJ1UfpvhoK/qvll1iJ+wy+xt/wTs/kztujorgubschRhKW
myvFsYylnCFfUhNWxCTKnepChTtSopnb/TEkYBUi+gourYeT+n62F22L6WUBISBPwVpw2mI3BxgQ
4/PP5XF/Yo/BjJpsPkEXYSsw93uI1K6F0mfm4Pm4YNwJew6fK3wVnh0nh2MQgyR7kCuBm/fVvGq0
l4ZwDk7l+6t6ccWldnqLAV9T3A7shl50C8JsanwoW9wJuCoYN0JlNo01mysNyHe8w4qSADtH3x+1
ezN+xTRO8AelFwVqQZ9Qze7eT5vRX7A9LPGX6blufZ1/IODBtKS5VRJ+08eCVsicwwZ1hkdRFqKr
FZ/aXXV8CN4X98LItP783TlgkJ8yYo3hUdl/sr21wmb8Sy141TFXJwbmA0DlYpP44LEnFOA81J3v
sKZiXINkjtoi+qbJPhXy2FJO9oU1bKGNC2Anb89n9S4h3RhtVTiR2tnINJHmzCzcy57m+tUrlvRW
84ulsySYNzlWz8bJAe8TtgASmlaZDvDYm0WyPP85Y/PhMsyRYMC0s9t2xb2PReNpX5Pgp88geksO
YaejNPOV3uCvYlwIs9sx2ARlVoD1LxEW363GpAfzj765RJ/1ryioSpw0E8kN/oUAztSkX7FYic1I
KzEsyXvyflnHjAH/O8fD6Vin7TqEklRUS4Hlc+1qQQ3TC4c251RrkpPwAz+hI7+fcMSDPsc702CP
ilJ+fMFELOoGycKPH9NuN9KOn7ghjyHt+0a2lRPMURq0z0UXJ1RjViuQoh2iph8RKY9wfW+BaZqN
32SuiWalO0oj41UlR2H2urLZ2C9QVVbScAQxEQcE7SPfgjQdYShYDqSg1gpdXmeblY7hKmaY9U6U
5lPw97gfXJuDTVKkeTgwvwSp4qvTd39A1Sga5VaMxkx62YyzKWZedhcwsxeG1C2Y7kF0OlGUTk5D
RbOIXrAZJ+Lh0+jVqTzi6pacEOSDROO4tNgLArHM6XOVQU2/85GsoGEqwj41KWTZ1ZfiwtApjU1C
Qg4NcZYYVRmwKMKqGju9cT1oJqw/xARQWYeFqwdvZNP2ytDCnoVZ8ruMRh2uExC2kzekte6ebnRA
/xgkjIxDHLpUukzqhB2Cdg5Oi8NWAeLfXjALVMMBhvHNgoVOTrPnPWW5DqxD6HxPMWTCWe6zzwMd
AZejCoXNgdDFknWAKr6P83XA6qhXi3+bPNvzAF5fDAe8PbXSLOGHhijVXz3qjLyFpUVjHlTqiZvS
Y9Xpquv0X+hX91bxC8nkn8g7rL9VyhtbpfVujvU9grViI9oVWdALlr+/uhVnJPNjEDSX4YX7//hu
BE0RJUVeyH/x3vWqC0Lds+kJ8Ju54GxzEJuuwbl79qbsDhl80HzhYsJNuFotrJXZOkoK0Qv7UqaF
krWpLCDulgVnVCYTpvL3itoZ4Xjq9jsR/pznYRX8GYsT7aUXe6FZ6BNZQk0qlF8pbNJZFPJbWTat
ERsKtKGoRkx7rrlycEONJIzvC/ghnvrtEH93E6c9+L98dNtBqGpvRlLhQ5ebc12//aAiU4PtPpuT
Idh7Xjg5tauaaeSM9Q3SDtVbjZ7wX7Yvvwa4JyUqVhznqYuH81g11WJ8Qnw0sgiMWBtFPd4Y4nZ3
V01xx8ebka1oPgDWaqxS309EzWZH48UDuHizl9Uf+QwKHOT0N5RyLrhPkVQdy2tCtSvkw5NizY2Q
L7D2nYZrSEy3Mv3BI7gOoKCgrHP5xrJ1vUa91S+reb1JQkSWjY3ab9zTY6rRfz3/aqzUCVMMHVjL
iQsDmoE6YGZMpyP35/R7MPItTYQQ+F6JiVtIb9gt6pWMH78pnCWZZIR0qf7v33+Q62uqOoE89w+s
GsG8yR7yTRhR5klcKkfrAeu+ZtVYvaa+baAYKbPCwJZ/Y9PRYlWCGkp4E3s+uzzgrHKjlIdQZ3ry
qrDoREfbKfqO+2Q1WX+XohY3fD8zpB3BnHJxbo/g4C+VYMWL5Ig5zZBz0Qb/4b4gg1FdWGlx3ktZ
DyE2ko1OIa7UFCxTx6qZIVF78wHnXsa3mExSgvCdmO3CH4OoLsdZa9AcR+UXg/DGwB5aaJBeBxlp
igb34uUTpzJIyxQ6Bh6cHH0tvd37AVz0YZVn6f5MnS/93FD6BTVjPKupNoMtEkrzs3YkVkyKIlzW
XF2mPqBVwe2Hzj3HMQlMTllhArqg0k6yVybb6CxBPKFKgxZIF0xpLi9BOlPNurlawXIa96WPNVLH
gC9LRRWftVOWqHVrwIgK28ILxpnft2kgvkiz5ufzkFJuSqRag/ZWFYZzm4xHkbukc7Xte/vb9kl4
88VlnuBikFn4O/9SGdsgkwJ/m4UWUbE2KRifvDM6hfjpc4BsUqlXcp9P7zggp+QZ3UP3woB0IKSb
VGjogIvSCwbIAPBy4LADNTGG4i4WEOwDYC5yw5sgmQypMjsw6pi7mkjcnA9mBiP6zxaKAY++YD94
b7qNJIH0dXvIl9XkNd8uzKkcP+fRJMRlKj6dDxS5jcOjTaAkgD6kwBxAJm8dygPvrVEmqZRBxrTu
jwRSf9L9HmC+xrql/YG+hpxlbZAHbOsZHCbmq7zlGUubJxaPf55+o8Bq3OsHfOEjmWi5H+m/hI3p
+ch3/VLw2UcbivUx8NHrN9piiiRmQ6nTroMexajaMAwEdQdjy/rJmGldzYzjZBBgs4AZujm6ATBX
XjrPBXil8FKacqJXrVMOqjl29kWu5rHPrif32THRzP6S7Cy2KgJrgVDjvsaGMMSHpYRuu7tbpRf1
R+bReBbuBnIwY0Gfe5Kvuo4697EEwwQgPVTR0NN9n74M3Kj6uIRnWBVtzhZlxkpJRhYazeppQ+NB
D8INv+SOyHavJU+P5p27VvmwHcECsybL6rDQu/R7OMjQy2qFaczbnpJg+7pq3LWlmdMHyzpXe6jW
feyig2U4tIkoS8iJDyVgTnt5ClJ+iSBmsTBq0RqLKDMhx4n6RUNk/3mf4Yp06J5rIr/VIkVBBDje
xdeo7JvSZsiKObdguheW97/WCw0kfbCAN8xSGUVJKtFx82x5wHtNX6UmwI8cn+QsGnncbmp5Nf0h
xhbA+3RAeAYVsfXWj1wSr9zk6CgSX/KnKByVi6/bXtpy/RAzffqyhoESWwkiTSuPHMLmNkekdIRm
eSeU1WpR4vzBQluRLJ3/U3MitZcq+S9PGaOe0U5mWmM/4pmhiNB/o+raOGSgxGOtOrTiLN8noJD2
/ICd9zrsmcQq7EzmHvOsza8urAGMsTauTVnuH/T+ZbbyeVsbX5gDtFy0wkwpJFNQ80Hm8s/DtCmW
eaGGiUxkKSGfQDQG5QxeZMj6hSUyyVZQxwKjJoPacSoKEmEEeo3J9IN5A1l9xrgdJIXfauYrYXVh
4t7EkLE2WZvkdEQwzuTn0Til7wpSIXPDxxwTcdhZcty/ae4eBYI9Up7XaR1fZoZIq8YuAQ5Jbcqx
PN5o3XXV2QN/impT1+fACZqgUzkxGk3am0UC6sXHohOMjR8jE/CN3ugyOzwyT4yF15tCWSsAbNJW
OWLV5r01ncYALAVP04DjcqO1a02pxJrTOBhGhYQNFVOnR9/XYf+qgXeQll1zyLRVvIAVVS0Xttwm
ob/BKVyppId1vEhEwA1khSIuGrRkxgw5Y8/2nHSYFIiDgaeJd9SwUfpmeqaY6e0Dsn+bJHkFDr6w
syVpbFsbabacH4K4o22fkZE2E+BX5SohZSvhKNlfmWOvvSeLw6DpScKougOdqO1RHhEub3cutA31
GcR16G8l5+MMakdAq9jaTJNvIY2nxGd0D2rvySEZ4VVLdYCq2OspvmKj3wmpLi2cN/743b2MzBcO
NbK+bUdo8uhVYsS1pYSqz9HZbhRoD3wpa29Anrimgdvwv7Yd7KNEflvlS5QBamYiqJfQs01GtjzR
bfslI+xroYyacHjAgHeuF029K/M6mFMblj5M2WC/zT6xfnVQEMlSvOqSqgJpkwVRj802TOZ/vKA0
2ydVczK7rEc3sEnWlHHwgIxnH2nVTKgiVM5pPXWtaFwSUv252HQwHiPpkbMy7OPEu3L3+gvYCsv7
SUBEk7X6Uin0XtSBoDcvjJ3xM0uJgdzX65fPNtyRHWgU0oUeoYZUY3/I75RLGHrETxc5fkDgOQyn
POlHyK/B7D+uThA4oWSPy/vHUvGO9O6Lp7jS0TD10y7/9jN7PK7AKc0wygdpdk8GtcNsXEKqYUGZ
QSIiWJ+yHR+kY5MfMoXrDWWepcq0dyrZ70j0m/IoTsKEWU4YcsIXpA1D18+Ly03VAsLy0dWLvl8w
ipejm5DtEPNcdU4pPJ6OJ9asDjlaFHGvFqLtpEavry/K2Eus4hby0VRmsvrb3LOPj6mK4fsCfYD9
mXkbHZIx0l3pBLXNKe1I5NbJQmCBbvaHPTaYUCVwqak1LPYw4Rr0dM2s3sO0qzhv0Bo4JHvDoGtg
LMMOoWTD3oY33iVI1DTXm44GqSFiGDBFo1AS1+rowXMihW1sgKHbW7aGvQJaI6C3rqFjkBlHKf3X
WLIidA8WXKcMzJ2de/4uofaREZ4jmhynuzqXuiJ/11BkIHthWiU/9uP24kzEadFKUhBmjUTdS4H1
E0RdDUM4sTBlubw2dDyU1vylH5qMMBv3EF0UF09/HSeJCgTSW+zM75LWT+dsayU6liyU/6nOv0lq
/mOOKIOw9G677pFp18t9kLccC1yGK1J689g8UFYc5hAlI1VQVvne0UN4mtluQu5MPcxwY3VQ3YUQ
KI5JnW9+6RqQogtaW0UqlDm9jQemi7I1CoDTHL82m7AnFvh7CHu/lkxeM9La11elUZkvieVN6AaZ
BjXGZ6vHYvOJSxWaVQSHWjjpyql2xyeKaeEhA0SF9GC4VentSq3SWQc/NFsdLKgCQJ4/QOMjC0u3
I3993dO9dlWp17m/ByTsR+5AMue01LHkUeV43cFP7g7Z9EEgig5zovWucJDqwVYVkq5G1YhIzb8b
khvOVIYGui+poH+y1V6MPvk9Ci/CdtSswKch6PFGngONpcOhJTI0dHT7QHeAX5bwnsjbQUKFSnFy
lAOQRruziSztgMfPzaXx+Fo3SxnPlizoUBGtROnBIE+UOrtT8rsxHYl7q75p4Uq0DdbyPauP4+xS
oxl81Xloz7IPQhIWpofYdbO9p2Kz2OAajC2iQGzVo6VJY5lZMbZlPvaXffgDHuGFSqAi7OTJicVo
Ob0fssXz/GEDvQYROOMMJXVU4Sq5Vf5RHPTtK44d40bxsved9Au+FoWw5Zw0JvZ8A8WXa9XVkCuB
D8lkrESLQhI3x6kNGhsZWIP1a0f3maZKWRZ+Wxwk6xkZut7BdnJ9hLuNxk/8MxfxUCN3yyLbZ2Sm
Wf3mJ0Ro0AMjJdY1De8/Brsa58s8kZbV9U3nU6OUTBC2T//QrMIH4gZx7GcelK3ZdY/6ZwEdCFhI
bpyKjkAhr6bPCo5Nfv0ulGaAs1POrklVTxwLKnoOhe5IDr7A6juHV1gj25M6nDiXq7NNAeeXEk8t
qjCyERYpgYbTp09pqH1cPgDX2Fg1ZmrR2BqW+bitAXx1lyeocvd2Vrim/UvC8dFL69O7pjslbwij
PYuhxRxLDQ19BpxwdNf8dReGg7ldjjh0dGkfP5ptnEvcBxzIjFNkhc6FUjnUGjVAqQu9lsXCdu+u
hEML+xf8yHg1KB9JU+DjftJKdGKaOeI+YvBTCAUdvR5OvVMDwXhyCCDLwPVD+Fmi+5DbCV00dkM3
kfS4e2415Gmfr8O1SVtMiK+Q7weo6HS5WPcHIxAP/Is41wWHZki+yArmwN/WR7LYg2d1djOMrpdo
h5Zn5HSzf07AbT1wfuMc0brj4Vk/0LIzTIk5IJXRSD4X3m3qrBt8olUgErRCpKS3nmiEJE5U/9p4
COwmYx3dXsDwVzAqIJeniQ0pTkh8VhFsWMOPgj5pU+NpYS3U0bKYZKCUeXHfyKXZ2h6jrrJ4WyAK
PF+x8jeTGkZkHlpIcoQifzOt93X1x++FR/sGFfFrlFbPJHJww7b3/OG6+hyM1gsqKwIpfXW/6O90
GDijqb0LaayPH9KQ7NJwMg8tIDeWzTO4BYgnuoCPsu4cZ6BoLrSNkC1K23zdK4YCWgF6RHQms+og
H7gp7RW2xImyUB5eWjBmOHIq8kW2VzXwd5EkTVBk3Kf/8dU8+8cE3F3w3wHVJMTyzxffTsZhhj3l
3byVx+585n4ld0kG1x1wmOOQevSC4hwADhFqwGIGLGk/Oa1jgNJ99pWsO9qvOwJn+UiE8My/xJxl
zcXplfvcty8sRwfteuLBaAGEWfsH1wZlupsIMGQzarn55snqsSUsW9hhsCCSB0BGgTYMEvpFSTKm
oVDaodvNS8AnLf4UI7mm8oG5KPeBogHIRiMgZF+LY3Qx5VAZTwD+IcQc43a582yCXlENnD9xWd4b
dwPmoWLBnHdvtf7FYAY1PSh+f1K/4zb75dVIH7i0ODAqVceZZPt/mccyRos5MFcZeRF40tWPtnQm
5pKJg/N1s7uYGxgd7YDpqVvrDKlSY1plFQm+KjFLBknI21IlYGvg4S6lGC9xtkfF7AB0jzDy+z1w
kcw6ZDM4wZBXCk2ttgn4QueuNDQ/UBuNBp7CPKwLfGeoDdM1OnN5z/NELEI66G5QYY0Er9Y02IT1
G9HC0cCL6UWdXrdKXwLQBPqNT4uRajSsA0hEteWG1FhzSLbHQugMz3iQCJlAefKlygHhKlNXcS5v
dRk3I1ZBafmEPl9XS/1stheY6JZB0FAcU15LlA786BnSt04ymbMq/xMO9mEg+uL4PiRZx/0lco6V
7u4LAxzVMOcSYeDM/ASvsF3NfPECHwR9FWmmkcNOo4TRJEL5QSW3RgfZKHYZepndl0NIKa508AHG
T9xMk4ZAUikOnbxOft0xQ/zagQyRO2/6/VdhkLQx4c5yEqw3kIAt586zTxRRKVUNj8JRx3cH5JmK
ky5uyiwmtkI3FK+qv11x/hhSDJXvg8bG+G2gD3M/0BonCBOwLNdvqaGnD7+V2zcvEXOLN6zx64B1
Dq2+dQ2JQNSD/VWRSljDlTT4To016ogeDLO5HxxrOcoLw/Q9agN35KCopQD4ENeauEPmY441iMAA
rdYOL+2xvk7+vocqtiLZmE4ei1W3w8YXVvQf92UzBMzbkRwzFmdbW3iP/ObLkIbnf0s3LLS7ejvZ
y6QI8fdVu/IP3vcTGsMP119mPVF54NbkdjVKlQkNXoezCMPwjoWq/Q4CWgBe/3Q9RAN/OQPf00rn
bs+UVnJqn4ZC194Em5EWppk9pyLZV6CiZHK00KjxUrmxPwoSuH+bbkKhHK8P8Sh8sueV8pLfSg3y
LyDvI+nt6D9gMsvhzGTQjeJt38ERef0VEYb7lA0dRiIEFNIIIALxX8TV7hAD1vZgx3Pr67zJtImk
gdsS5Q/fN+eYK9ai2Y4IyVksWsECn3DI4TWVppyABq9FEetN0nhkA91GhEwZEEfKo2YdKWnDBmBA
x8IUBvSjnGsRqFfBseo4z/gKZTekg4WeYSjHuMU/VST0G/1wN7jdL/SgQPx2eGhVXpyuv1OzpqVg
zBbGDzvsZVLjdDLoIMhZ3LLL0VN3FH82Kq0vv0wLnQXxsTRtA5I/SEr+QT513HaSSO9Oy8F4aPWu
jFM12CKFfNQ4pyI6g/4Zawd2RKKfY9o5TvFPEKGWI0IlPpxwLtqIijhkVHGGq1XzPn+MAP8JlCAG
v6Qygd/uA3G86FOjEsIHKpZszwEA1MC5tXazQWevFUp9gQjQFoC/XEm7VyVN3Gf3dWjIwGvLrOak
wVhC1Si9xQt9YcH4PXHxodxGqu/TTLSX+wIdLYjvxo/oYF8qQ1aCYnnR0MoKurLOlNY7WfNy0U/g
qphLrWYIKkVZ4sqQiFMlobrHK0l8a6qjcueY0lgStMEWp1joWOtutExSejq4+xAXWuBxzSixnHpd
Tns0lAsS45b3POf2WW4ZLxlofhob5yE+8w2zwlmckJem8Rc365wZS9Tzei+hg/dxb9dFKvokhRfC
rAtBJcv9OxMGkOLOmwoWtNseFXTkq/ZCxYnFsRYjDzhVvCkjt2ez1Q9FRxKakZ0qY4eE9CoT0mk6
Akoxp5xPjEdU8Mel4iP/nyNSKbgO46SAAVmlqGxwaDVOZD8NE1lxhGdiv5YwuAIimRjquMsd0gay
NmUcAX1prgsi4DGHghTKlJyXXcp2t4aFI9WrjsP95CIr+XZymDHPBW631mlQrmIDp4y5Ycff5oDH
65oHJCh6oQf9SedV+sg9jSxOKzThUGtDwzZVuEyPXK5SPQ5Mt3CJ3QdxNddVt5ntpURX9I4prMPC
Nkgg1TQkahpizV90VlhMCw34im43qNfexYeYawiRlVvjYvV/6NKOh0yCKiLf41Tvvu5jx8IN5Rqi
pGjBYaxU5VfqjR/azoibBF3voD6ZAJLinprpCRj5jGWNAOU8Z06HV7+pSqw+iUXTY9B9ZRHgmL2s
yCJ001QfLozPkF5PM66cdfRsj443wB+2tYiWFLpiXu3RE4HU6s6YcPv3LS+yKI+UiSZrUgqHBKgc
Vbtx46PIBcT+XZz/35jkyKZpNUsPjko3TUD6zaNAmmBjwcOKeQSuFAaXXP2ZNTGQS6qfJIUgLFbl
B64WMhjBpmgExqx9HcHH8uOSFqSS8WpHmYndjCtNVSYl9aC4114EcScw3zKys1YWZzTIc/PvOS4S
op33Ch9UqvuFOVImToyVy+31wjnheyr8GQVdL069vGjYsu+ISlNTcGOA7xYCRTW5spLMDPZfk7LH
AS9CGPB680Sd4kAhaRGqnlXqMzbqlY/KIVuQszH5buRgmtfuvnrj83aSFpbq3ayvUApHW5bF12dE
IlAToO2LTjnoj5tQB35XKse0wLwb1ePyw1MifQ2f4uMwHCaFfKy4jVIA8FFdsoUoOpXwNXylxrxc
7AR10vo10lA9dwDhdxztoMVthdzUYMw7p2jwhS+nsP9K4NDZOhnuIpI/zj4yw+Ev8O0btyJ28rvz
Ibicbo+5wY1I48Ez4qBf4r76MbOsUFPtmAQP1OFbuhEhb7LY2Uy6ZAEtVXIbJld1fAPABajMho+r
fjCDLbGD0IFKVe9so5MbJ7Wt/T3tMDVbLf4Jg49xT/yZUlHXfAuCFFz+BRz+ekv1JYPil8z8AZ2z
xoBmOsrDeJ3w1r8x40LLeRhIhqv/BDSy+YJ4Z694rBYM+/aLr5e9Bk+4j4/eoXozULh3vIAuBTkO
1Ue4h3MP3mYVU68b51VMjPETNl0unlV3xUyoKCXUtt4etepUjBKMZMIqGpJC7DQ/ePuXrKYmnu5c
ZxHIKzFgmk62lMWjSGcczPQDPTyskU7EAkpGVQ3iCOoVLq3e2SLPf41m2DHg+JhbYs3TA6g2js+X
jR4vBBUCBUVXp6IH8K6F+0eJUQtGps0JYQNRmiVcIhu3PaWyrz5IoMrdeZ7UCwASIsP27XuU2xXi
EBzz1aA5jny90fGxYzV4/Ok92sx6VnlCtSeuLcN8koeByiBG5TdGzKnqX04TcRfTNWemMTj+54ZE
gENUbTCMoc+U5HDxs7uU8VT6VDRZQNyJ9UGfUZVmsGkn02Byu4uLB5Z7wU5UjRt09TwA5ZS5EYxk
Quo81CSVjzWpli2WH8FBX4GQ2IHZjM6XYKlAQ52zy9eD8oG7a7qSOZ1T+ydHxIN8s1P84XBVUM22
BJwmQ1rXsWZzhC289KKacxPkES6O5SLUN5eq/wikK9J5nhZxrtn+R147jofpkwpZpRNtqeraVzhZ
DOW3JnPJE0fB+pvEqa30vgsIRVUQWthA/ODUI3xVbX/siw71OxaYf1AuScsakZdQBFh6Z924XJeF
9tdLDNc77GzomIvA885yczSQIPBlsWuhiH45varZ1AQrcnh/lZLe2Kht1okFI/5VfeK7tPFpSqMU
kL9Wu0WBasKOH/ciS9thJ0Nmnh7vxHO5HKLTKvjo/rELye6GHLwD55L+90w0UEHWT13r+gORCdnZ
06H8l/80Ofkrg55Pv6MWNhzcYmPz+a0RApEJqdch5uXiBN7FFrNaWMsdTlTDp14wF4r9A7h+CgQC
RQFviEwym8yAhzEAW4cPG+yNUApl2gJWdPWTI8X00v9UIOahQVG2N2DX9KZ7jtebL8pIXrJ15aDv
1jraY8nUZyWPwf6fCmgDu+UVjtbbQnnPDGB2/EQHWS0lUqzkSzIuRVNpzCcVLUXMTTyUXzQagJUT
4qfbdx2gZZI2oem3jeDKjl5hCqJvMKDu8yBZoFXjMOYzQKuTMy3POdOzXxdP/SqQ0XJut14+wz3d
uX9kQl5f+g3SdRnXQ3YlWZ6jvC6gZGQ0c+1pNfyvx3yQIMK/T6T49nF74lmql34+BRHR5Qx3+ZIy
VMZQno6v0W00jXxPosbrSy4SKop/l3snfAEtxs/2Ckw/L1tEQ/32aXmJsw60bKdBHiP5142XLwQ9
fQvkofOezptGNlzRzl7yULWbpPhAdFvgr5DqUJoEUd2kO8wV+VC0LhEX7v2andN7TPGGu/gr+7rE
Dzk+iG6v+Sm9UOn8kzyxCUjmKktap/4xkwTUEV5geVZB+3wKP3Lg/vJpiLCjDQXpOpqSPvPBaIt8
KK7OntQtJyGbnYEzVM5yih4K1WQ3DPvrhFMZma40WocNcgtZpt+khy+nB1Vi1R2ihiwczOeA41Ef
mbSyH7p55HndE2wBRs3gUDRMf6eAv+fBV0lC3P2bFhZHqlNFq7ZkYnXFq9Umu6NkHyJStL4eG30G
Qcm3QOrGuJzxzqqv4OJC9zP2OxqK5nbETeQaj5uIZcX1OmTGI0IXnNy4oLRkWmOlAs449vnuivmZ
SS2+i99yxRZiKkPQldR0SoZexKcl1OdMIz0N5uXAyKvIpUXMlIWlk2xkjp3dJY7ElDOwGE/TZIvP
fv0SK+C6tj5/UrFBsyPBjU2kasZ22IoTMaZs8PGEhWutsdHNxbfNx4Jl2MRtdc3qCclMILd+/2GD
VDhCahZmloSMWRBEsHkJOpIWkmG9keq5oRXVxwhwUTQats+B18GrTXwSohiEWax1cHwZzDCcStC3
1uG2aBo2F9SNyGeLfR+Fyel3/XLTal+9X/0S788Z/fUNmr/tOCRinWyJFLEatQCzUoLLOMRVoeMd
q3N79ob+QcSMIXBi9m+rX6sBUt1xxMQtmMUu/vDYiT/33KWAV9eC6AcPlQkw4ZZTTwXFKgon04nR
YR0prYjmQHx4XFCBeXZzfPPlimjjLWJea4dC+VbbvRsP3TWcLjumMOawTjTzZK2FLCd15a/H72+Q
0lhk0RWFvP24UiJ6ufO0fXXyHrP1IyP2lz2HkuWAl7m3dx/Ps+MPPyOm9qFzVzgXIWF8BG2c9q8O
X6+nxucFav+0+yGMiZ/A8Dg0073YUTUazTDbD1sfO4zchD7lT5YlVFi4zwfWXnS438EOAuhkISXf
zjoQZVaNwU/0Gr/wr65TOxs7RViIajkfacAalEU+HfBRjQrrdUmIy0lpmMRWaB7084ZG5Br440yE
EejID+hBKbVWOcqV0O/muvsjDCDUGB4F0uQZcCWiqqr98LzPr6t4M8MIgRa1Xph/JkkzLRXhBPI5
CSOkNcKEt/E6ZFVWY8DcNwUaqmCJAXxvw62tMR4GC0okBIzPhW2I38YpKJ4lUytYXK/tcyzM7vB0
H7esMl2WxgMOxoNtYxGtVBoyjVr/UAhdugmqLMlRpN9Kq2uag7l/4rZvzNnnXKULa+hrBkG6iMw4
fHp4+0yqTCmYQMGswvMjbhdhzlmoy9Ikt2vHvteS8iK1prk/+12nn9WN2TR1xsrQqOCtPoyxAAp9
64jUbxP/kRFvGI0vUToVpCZaK3yqeC57g5Is82Yv8RFJthe7xPxz3/Q/R734tAOVfHW8M6SPuLjy
mKjqE8m4vh+1HCPXYbbqqlTXFSv3gYodtdFVJJZ9qBdDQm2gh7XQMf4rbyP1TNM2KN3I9HyInPWe
pRY8pmVJG2q6aihhBYCxTrtbNXAqlpARY2uGCiVxuA3nWNM8EPV32WBJXev9fUgq8ie2TJ/zWboo
xoTJ0CFLFTWwxzamll1Qiwq3woBJWiXz4ukzeOxUM6YvkCOkBUHXfWSB5ep8W+GFmGJJrlMWjZGj
Hmpla4zz2oCGSnQvevG14i+CFu1n4lWfJB2Y9G1umN9HX0LTLrsefzaMbwilyaIeZHEdFSOU/Udj
u1uOclAXHEdPQ5AN6beKCYYN4oTbXLXb+Rn1PT3nnoBqXDBEBE9kvHpPUzS52RCU7NVOie8oDeVo
vIj4rKX3B/YecesTeC+wKEiNd9R6OtUmBK9OwvAq/N/vC8Q/bRuwYyRVAfo8nytfbxNGuQwMFL90
Q3aJYdHNQN3sEbnP1MVmqN37aDpAscS1NsaSAfNIi0O4FYhVB9F/vOBye64JIjA3cBrp+CiSzWJ5
xmAgqhUdjjt57lh1n8j9dE3t7Cwi+cwlaq5e4slV4QZMestSxiRR6N4RLOJPoZE66mLmuoQ/CWPl
hFy88/d/m0jl8qFv4FPFMl8r9qavKrNOU/THWx01Pz2DQWbcXb9zkLhm2wbjWH+TNqQb9iyjVE2T
HaT5FrjvroYsCgdO0dusTxqTog3GvEHlizXmzmqSuj4KYQkhyGo8uMhjKbK9z7YXMHuGSJDddVXg
b1Gsi7eh9BtbmkLZZ/xzvSufWECV+SDdVElhlV2d5+QfL6RAs2o5NLN5bZM8HrBOrJso4OWm4HO3
PPPEQlBb+Ls8sxfYoF7xczY8lkE7vHn5n+iGGVwj2Jgyo2TEhXkSzWIvAf5ZgEpsFyvMGatYKNf6
YR9eIJjY8ftM/Vmgj7TwN0m27tqx8hylNjO1atubp1AA4R1dh9WZvGeHevMgFn60XmI8x5IFw5wN
8oHWfPSH+857H7iAVFMSn+4kyiW2hy55TFwVx60kEeXkp8QkHQFTyrcDyhMGZkgIlEW8SmEQWiFI
vsQ4JQtlHZ1O/rXh/mNQ6ESGwcazfWA5RFM9unePq7spu4dWG3/RzpNwG0uyvCG0m/4nHtI/ZP3E
i4seT9KGQLuxa3d8u+UYCizp5cWOe1uA7CoWjL/VxpRQ3ws7wK6AEpKKP2piQ3Uy396f6l1Un9Z2
K/SylS2ylINE2geeMnh4Q++f5Mw5JZE8bDrvW26zYvaSe2nTECf3WeJwHLSptuwRP0+UKTlcMXAC
NHvHn+RxE1cKi7z+kK92eRxHjvqXRqV/8XlaXds+eDMEz1AvkJqx1fAoFvxzRJ8Q/036T32mtZVc
WFJGAKM53Hs0CLKViSI1CNN/+4BX3+BsnpVC86BDNSvhIByBloTd8UUdJ1U86Kd8Gt05HoBkoozo
iAK8e2ghp8nlb1EcLlRK88cI42ZCYIQQQgmSqxcEuT55GBHTrrDe8wd5UwemcVUAKq/d3JIDpZE3
NSLO9p1QpkU9XBFWQ90lYVrWvmOcAzkbzpSLMLZ3Bl1KDVwbrIZk30DXKmu5n4hP2jedDDgqcqrn
aH8XSp+L2QHbNyxLwfIIqaqycFvVBwsyeV4fvyj1gvLD5jvPPvNZp+/K0T0hKgkL6unUjfbSs6R6
yrfjFvP37XsEX1uhpNKROwli/sJILgYx/kLnPRnflubBc6otETlhm6wbPtUqvUZnUcbRSDUCiHlF
zBt7wZPBZ+r/hhTiq3jOrkuFD8AHgK22R5wqFou6UZLO/MrYVQ/T1ftF4toeO+seKp167MbIVFDq
maxLPfl0CEncq2zBv+HfYJjsn5T3yBVq8uxsYAQ/2AX2NjUrFohO+1ARAObFYxG2kFWa4OpW2iPN
bGSfmOzJYQ23IlkX13gFz5KhUUuRvxubvX+BcMwRAeYC1u2MAkuj5WtQZz5+Hjp79mc2c9o/i3oP
BbJKdEUtu8GCVsCWhWQ7lyjtEPxKbMv5IGEujNRcOtGhxE/n8puldKbLda2pi7TbHQoPeDn3kp2x
L8dNSgl7vYXykOT68V8rQ9ECJh8MbVLaurCJoJi4jms2k2RplUXXPxjcS4LhfdImq2R5l5tJD5bW
jZ6yR96hrqteA2J746aMmq/nnXlYcBN5TtSLsxy8Xku7/Scm7a7/jTgXc/db4atS+FF8RvsqE9rR
B/Kfz+0uVqwjxp0jlnvzg8f5Fr6jEq3UM56LPWKhyGbD2KBoa+vRrX6hdToXr05hK7n9Lny7JqOf
ODh4RTBzBXUN9Y6d9bAHxtE2B3EgImT465TkPh1DX+ax5NY1XDqAwMhMB9btQkz7bmYCEKiEWvZ8
hoJfT6T+0I54FTAF37jA3EUK6s7yslYhF4uwzC7EuV5crA6GkdYJ9hEj6oQSxRSsEmndFbtWz3oF
vVA0i0di3l3Ww6ArR8DGD2FfFTgCgbEc7cX8HN33q9VA2hEo33LEjjEiZZbm5s52zPxO7g+7m/xc
Gb07vdGahxVkEyN8yH9secpsvho4OejNT1VGNNS02x7+xFKeFxb8kK5suDoJO+Ssbm4zhX0xC/EF
idMzxWO7/o1Ju9pWHKEilpgXRTblyZxpfybjGyOq63zdHIbEZokCrFd/oN8KYPaLzX5Ylr6QBTUl
xHHJnbnyuKD8kKkQOq2hd181/6y+FSNbE/leCd3laq6jLYz0s3dSfcP0/nf3tym2o9Y6DAjA/B/E
xr75qf9pwJbUidJCsZlIuMIEJHAc+rgKEND5VBrvOTKbQ+qX9T/yuoe/i+BTNYLoaNlBAAs7+niE
8fn6AzCOzuAGWcyDlVKpfxGvuv7nRSfkBf9kQHNeXGMrhYyz+HZEBVhvLxJClUBLTAS16dPMACGQ
hLm323KTtx3phsRbQhhKDZMIriGrttECDSoujUBcOf/RUZckX4Qww3w+Y4wH3AR3sw72YVzv526F
EqKpg/PCAunwPLb2aX+i2dtsVeN4kdlOLsjrChncKwnbxRrQM63ZpYuNknvWJ9Bo2AETFF0WGX1v
1NjfBZRPZnwTVxt7egQpaw+B+mwTBBnAuZ9lmCTIT1LVlWkEI893K42NbsS6Czs9iCM+3WDHSQyn
Dd766AvTaNAXdlEoul91pckz2fKAlTZGWo/ACk4lmjjd3r+YTww+TqWVKWeGnD1MQMvZajidcown
sDMZlLKhp69QAovCTej+vxc+27f9slgiHxRKtb0pEJ6Dlz4F8cUORW8Y4TpkLK8xpRPQvmaImrvu
5cjCdHHv0Lh/xm6FNg+znMMSFnoLHCUrVoaj+QLnkxl8PVfh58GcFF1viuRtMUbY8iVRXkdjUhZ2
+t4tXeqYLy1yDNoFqTWtuwQ2xWzeExqRX/qq3s8qmkzK/hZ7zjpU4RtiijY3qHUQb2WoFa1mAzbv
2ALM1vQQdyCpSR3Ja+NNIn/aI9C92AEFxj9kJ37IcBqzCVtRCB9YAp9gTzxLn6cdFc/x36mX2WSE
fTXUO2TZJz34QHcUUBXZaY5gZknXcGKD3lEj7j8MM8AbEX5yV3zZOHS6iD0VlgjbXcN5orTVH7QE
4lSG9hhUW+SidHfI9TEAknGRwwwMjY4B34WTSVd53eRhmzgYAKMEAEFhubcKuHKqO5z+pLbCOCk1
E7ZKx0a+WpEa/8Y1F5uY/Uc4q66vEvA/+BfNVHTyGlcL6m2oEaewjoedGutIUy86ZgQTUlLkQZtC
5jbJiPO62yaKBhDhTi6dICaV6N1cVIsTyJViAS8UA4H5itvEzlTgMKvDTEucA9zsihYq6U7JkW8s
dOctLAcW1wKgLRyM+kMzlVcYl4mB6hQxn2nyn4WEoM7XsR3uhzo7nF4Dfh6CndGb3nUC8/6XjPek
sLps/arfffeBL4yZkw2Pxy0CZrt6q22WK8muu/dsf0nx1ctzL6mfQ5DiJm2KkM7nHmd/ZOravTX3
MAKsEc0OYJYK9WWcH587H37MR82+5EWxRAtNS3HQIPZEN5gXtLD9aFnkeGassivTlezDdz9apypN
XUqtpjGLLzWO/ccZexBu2/iO3YUe20VIEp/WuNXpU5PTtmrwomVicEdL4fXC3c5wqxGqKAtZxNF6
CBkV4c4rQ+exU36TSsF52G1L96xm+ODKmAspqiNCx9d98D6HraYUWeT0lcdMTxFoxfXP/0zjy/jL
AywE1KYaXSFHJMxxtHjmapN0LfT71xfybgjlLSWE7aOC+i1ez1IhPZYS4PpVaMXQWiTF5WtA9nVM
VLu/GYfhjCQXIitKV+X1fib7c1WxmXp9GjHlQPajqPp2BvjhhWNzpuGVpybWIV5W7ofEMRfnKIoz
h7/tCg+BZ/UZmJ6Fa0HnZPX3yBHuaE0GNXReK7P6MzvzFogPnc48ySXCg4DM0DQtNXmI5wDSjIR4
hg3TfBByykTtSnqrcmRZFyzwDWg4y+Z7WXrvJ/ABsJ1Oyw9AQnO/UnFM1wrm3srMvgiNXo24YECZ
5uQqb5wIiK8ijWbsQoK+gacq5lR92gPGlJIHUDZzEHKarHyLEj59fnYVC2SrhXd1MXFNkfqp5AE3
NgWp9jM33jDXb4dFD414P9qFEmVsXyUQTQhVelOslOumSILpYOOsmlqEwz1kscYHSBA0A0q7fOm7
G7jEqiHWoHYCMgPeKUc5qOBK3zvfIEe2cil9siX69p/eOW7jupaxFzjOtG5N2IOduxQserQeF/Hg
/bbb+cM03LKUnxZXlMvfxH6cHXqn/qrJSna7SyUr9lWiLcYaIJXAnoPhETh9DCym/1qyhC1yGSuS
l1KofiZQSdN8l5mMaA51JS/zB8r2ma6R5Ht3ReVCVRF6iRrNYgovraH0nYfGhXPx83KYus9W3W5B
kESGwytIN5agLWxJTDvC2rc+NOl8AXI3KWLNKoDXMypAysKbkxeAS9q31JAbUHpFOfX3qPyZ1YLc
Jg3SWaOQuIT7Z8KvcIPFvdxl6o6Krchr3gFBNIBESoXM7M5ZOmoRalFr+DGezhQiRxomMzH+XuR3
bfv7n/qLXzi10133eSxmXwxpq8K+pUN0FOZhLMWMZhEryZEJzDzUSSLxiB7SUaEvsMDVfF04CDYj
4S3ZuWi5jR/jH/yjyIxPG6NVr/F8cWWs4A+SNo5VFI2u0AgTnVBS1kkaq3B7v5cjsyhTzJ292FXZ
QY9sJ9KqcEjgg6oPzOLan/L1bCShbKiEzLadnwOb5Xk6CRx5qEOFd4P4Cf0zKFKIdcPAtCdD3zOg
lKqwXKktierR8lWqTJbuaYyhwegQB4J2aSLM6bA5KgZiD+03+RCNR4UbeelpGu6TNraRkrMxBuY9
wjfQbMOmqwWJU6K3znfrYygjbfQli94kut3Lywj6C1iRyLYf//0fHbnh7y++RvgHQsaOyXj5qZmT
OYwHqk2V8kRRhK0yq2NfebaEL1Ru+fAf3+bZzvL79byee+l4FrdTLsRLhOcflPM9ksD7hrTLs3mg
sO1UcPMZiOnqB0+ZuSLXMy2Cu1jjYEOBOXOvSTTYm0ZZGChK8+CGaT/jDcy6y+B4qQ1eBcp/7tK+
30hbGxsKT4+012LKp3V4JsgM9d0HxByvQ2sEuHxCRUIZPyCzJV1rsWHksnEVxfdQpw+HXHgcUpeT
b5B9dQYaps+sHGSAmR1IxMlZYIx7xbjJWGXc8DGfev/Gh36BEir9dkdBqJlUGxZjtu9+7cCCJXjf
wZNB2qqURsQ8/1Ujg44obdQxxSzUCqZd7O0SPsZNysPrSlf0cqB3NdSy4Bw2P2oegMpuIAjNtvPN
Sf1HwGnQ7VBZ+SrL6/cd0lOwHDT816QJ65Ee6YdP3KpvuCWNMAD8MP9QjhOGJGBArVbE+MsRpRwI
SyYxzWC69wnpWhkUBA+MQegv29JtybttiB7JSZTTJUKZ+8avgjBj0chnf3b+YWP84dOWJSwbQyUu
//xr5sqqDgZNXpdoTjU9FIZzJuZyINh5kqBmnB0LEbWQEe2x+/326/HSbMv+GDyPX5Os7B8HU5Id
JrXx6p3FXJIuEQUpI2SCJU5Q38WV9pe3/jz2HQ8BWOxfLlh/ocB7UTVAX/C34tsfAeGGglvi332h
zwN9KStUU9zxr6FLTXiBuApvn/xLP6rmtnJFOW3lPlOGrBYNk51LnyxstkAO2BiL3ulbnLCgKTho
jeHGjQknVB99We6SoX9EzkyqSJwRarH8yRaChhyghqkYvNWmYMPpMR63iAys14stx8QPSX4Df0UJ
SqQSFmFnuclzl8VFqH5gbM/BndtHzEaHRBbiu/IF9RfPPRYbXuGFeLi5luNLdr2uAMtLpVEYq7Mp
P0ganCz2bdiOmzd7RPDITGkuzii/tQHQ9SlBNHcUPG3maQ+YI+yuH4O99Xi8frFFldJm/gm2wt7J
0qexcLENWWAzDygBx1k68YIu4Xo7crcE+Fq4KkiEOOgKkYNEoF3unnsp5jtxOgltfWp0T6PpzUZr
tnDr0C1Ebzh0D34/Do1RvOEhwxXzuORsjisDcfrSAwCaywD+WaMk9VhWapZ+eYbPUCAILqGtIrNn
7nN8/zfRhmNeqJjqOOKLj0HYntoFCb0iljb4qkIU8xkTIfw2P5xmZ6OzwExHzrrdYyPCeSc1VE9s
HQYmcEJp9cjERAgnyxmkI8a6aomTl+kM6NyRYBI2jaIGYruZcPWezpKifmfMt2dwgosu42vsOGRx
1BCLy4e36yh215Z+k5aeSbI0jgo7rta7xyc+J/DlsFLq1QCHNz3aVH5rxJ1NwEE8P7czVlvHeo3D
zrsi9iRR+Qp1kwSC5zTsmxtGLpQFQ8G/rx+Jr3m87iJuWBUcwHvVa26P/OnW7GGdmVezZ6wkNk7D
NeZIIIi2+Wti/voBkfN/H0s7f4Q7GDtAkzUE/7oW1h8A7xNTooiZviI1bwf/BUZA5FiBhh5WmAzX
pdSPPx/0y/TEpRdfft8dykD8fERxVBJiUUYc3pIK1gpjegKNgNlEL+ZNP4WdSSTMPG9X8oMdbMcB
7GsRT3FNyA7ApPcpP3HyOH+Tdm4JxxoiWg84zl2YGfGAMAVeSCAWyYTAHefpQ+BYTICXvLQ4LlKe
u4UFCWEzl60Ica+ENYdbHz2Jb/Udmw9n+GxgJaTRTXZpXUJwu3WmfSqKTCvg7e+ua9DeLXwqq8YO
LkKB0ze6rsr6ZsnbZg+T10dEyVn08fgeoCE8qtVnG0pxHySRdAQrYHlFQjgEll7REbV9SkoBYij6
/v2YdQq4eaeb5h8Hvfjhf/jpTMf5jdPbZyjsPKeSjKkNkwSofYAx9TLVss65E7YzqD6GaIEpIb95
iNyy57vQ8SvOBXYCrIPoilOy+/v1xMsXLmOeJZVvWwxpTSBA4O4v17GFoDCJBAgt03M8yNwKhsar
bydBtqc1epWfk2rJ3Ee+wVgBEd7xmLVRk1JbmVhM220pHwpr40ELzZPAuxOjGvwWvS6b0PaCnQcJ
R1wcFywGXAHGtVCj+NaNtrrh6A02JuY1IAToE49m/13gYQzB++KQc/dm9FZjFjnMWLAYKSXJpn2E
gvXaawJwH7dwiwYoBLWSGJ6ekuqe401DWkESlNXzPN5Cv99Dqs+ExAgL7Q+LiIZAlvW9JhCy5k9f
Q4oWEUw+XcOTOimVkJoSQHGhTKHdUmJQnARQ75rxzR8mMqS/pOvu0EDIK9Qe9QR9eF4HI+t/Khib
Bj9FyEJ0WAdlE9f789GMjbhoiXhNFQw5WxIporP5xB9Ax7P8GI+qR4d4ATCKv2rU8RHv71d38fth
Q32FJGGlbNvTMhmOZu1itjrco7vYsv6lGS3L1Uiv/35cIjLBYiFHT2kRZeUICE/CB5b7+clkW0xC
RB9ZLEbSUya8kP0DbvmboLqvPii6hhyAxpCy8GunVpg3lROpb0FgusbtBipWcVvUrJ40VXjAJYHS
HhMAll1zsyuYZNkX8roGX6l1AKr57yeHwfBawoxYWDNxDtEuBQvzqPqUI38wK5BFmjdQgxA2dh8b
mDRDUnyPi0PyS/7Ghgt9I8KNgwqPZrcOmv3+uWpGX0+WTU6Rrjd/ofz7DXXNzUStThQM/zZGKfaN
CT9WEoryNrWtNgsISfdLY+zVt6CbT1DmUo9RymhhX9KSaRbHw9N2OfruvXarkJz7qMeO0h3VZrQv
NYUYruZXiV0wsQflur3EnNeX74vHpLHeLq+dwKoHMQhQ+zc8AGZn2tgn4cAsQLSQwgVZZ1vj+VSk
MrWctkedQahaZvkjfiBICrLF3iV1Zswh9dagS91nBznuXhMVi8BRTD6pPfRf65iDMoU0lm4/2Nh0
TtglOtAI3i1jj5E/3hfBecEjRAc/RDuK+sMY3EBVCSvrXSL6SOTCCGb3QooHLkAWzbtBqRntGn3B
mqR64layRHyZB8mBAFRqxdcFlvM+zJKFU0LYmXTO5CnUOvnXBuWSn4qvp4dtNpw/4yje+oRwmfLu
43SkTp2lCMyGvziQku5PSJ0W94x1NsuGnNlUbGGKaZMuhb3h7PhXdIlEUjIHXmBW5AMAOKjElcjZ
HT4kCLg62XSTsORfCmMv09BDhj5EGbmBu1Ua7yJ3ywa/zo6W9ohCDzFeT1/0/go/yuzkBqFvYiEi
4wAs2J2Bf/MHKuP2gcl+iJXf8s/SCMqlM5d2cUg42/NoP0K9OpgCBa/P2MGryom0uNFYBun8fVEh
3ZJW6tZIfM7rt+d7+gJEEPbDR/9djkfhKCGxgwo1udbXiMywFR/sSzUd9vnkhfw0iWUXfO+WTFM/
gkY8ur17BjmshNjHcVmjeHMgey0dF3+tRif59adFHKSPV3Wd7IpZbZ8dyKAuRKB1GPhMY7RY3h+g
d8MOFGQbYMxi5q09elnuOIWDlZ+n0z7nb6QXtj9rsY3byKOLeYWmCiwejZvGMhIU9sii+jCy5nlx
mgQXcA3sXXOEPLKbwH61nv19ot2tvpGjGLWBdzVWCFkhqkonCCS/OrYyUveCV8FZl5AFJ9vlHsvI
tMGRXpNdspbiFNEseAnhjimSlWI6eJRBYhzvz9tZWk5Z8oqVbTtp9dfjRy0amoIyv1hmyfP0+y+7
RYLEy/9Ncac5x6rGHj9a9GPyX5Nj7V4g5YjJmir9ld8RsdiO6U8/22QYyiawtPTLr5qn9724Q8AB
Gv6B6gJ9dyVnp8O/mHu0i/dcp46Y+ecBij0fqWqbGL1rlGnnVhus3Oi4hAbrPskW0ecOHgCnN4Xe
x0QQibtwJNv5rVTKb2143z/tFXPWhwqZpg8B7LHQtJQByXU72qum/CiZkoqxx+8hVUCZ/SIU9XBj
rPIi/G3BhPXRQUFUqr/ldGZseex0jyLKq2+I9xHV7eNiE1xQgRUH0U3/Zt+Z7fXVFf3vZ2SSx4fy
+mZmpz5fieCQg/M4LjlzqY98hHB7nw3eQcrFHlO4RPWy0IiQ3NGXl+FvTxwskCwHTqywjG0JaDlV
ac7OEIVmR6hMzjTAWe07QyVY9Z7RxRitiL+OQezNKLjOUE1/iZWACopLuNmuEqv6lKfbQSHJPQT6
dgdybwJY/8mLQvumLpmjyEjPltCVIbSvoygwezhGqMpYsYOtnyykU6oKSZ8bLh1xKROctOuuoTGf
dKQr0d2T25R3NTxMxUguxE2NkNwI8W3Zn4PyOEdVZ5CoNp1v7aCO+ygUc/lK3xxcFO/6MickzRkO
GMQBI6COH2TqWCMl1KoWqe7uOEdtHjWZjjiMjMztudbsYtXQIP6WEILXD9jY69VXFpvB/41A/k52
NdxuNHZSd4WbEFs0TSfAcXPZPIAwTQmDADXT/7+XRkoBUHPelut3CfbrYkIWr2teygOOxjrAC+CA
kpXootQWBQv3ixyiN9viCfJHyv1e2Bf8cpxL2GO7+eNyYZVMKVU7IlBALazCx1vjD9JPoK7ADL4M
zYLX99f4WmtgYrrhcHyJ8G3laF6pys1U2SVVcyg5kfgkDKxwC+CcOwBz46eFn0ykpWrpq/1HGVwc
aCJYeuhXkSDSp5yRio1hsDcSjB6X0OgeHCGiJnCDB77JQQDz5nWWueyJCsQN0mjKnmliFLS7WKtV
/KQ+z48iOlH1/TAH4D86KxKLx4lgg/xTWeyzAbLI1QLVp4eO8gijk4C82b3YiN2VnQLoW7bBvz4n
GyZgafMyypw56rrPbGIf4H8lV2hXvSY+9ysmkJFy2wBRwkTARJZVwZcX+RwMKvDqEoieLfM3Rcij
1hs8uQF5YpHg/5PcHnJeFH8Wk3tcGNUaVUC8Y71myRNdy/WAxfy1gC8bQCzHeRE736wovpJ6iOet
673db89IlVzTpsPOQtEHbTNh8WjJJjICSKRuUpKJ5Gd5dcCw57ubKl5Tufz49HKWqeokHKSK/YgO
/VJ5HfPM/+3LICYAQH6C0XcW7XnJvrImNGg/zMW9VeD6uzMxXZu5OwE/SySuzcDg+va16SNBq9+m
QR6+Gy8JVb81q7tQHVodw+YKJD1LhF9yB0x48Y+MHDpzfWWDyRUhwANj9DmCzp8gFOv3fQ5Zn2Uf
aNHyNRLwOVLPGwKcB0YloYesQGXbqazibRC/ahSzAxBK8un3kQwDFOUssEMv9km9VCsTV56byPsd
V+sx3b9sVfR3RK3eDw545dvTygx7S4f7KLzXWMyBMqNVos1TrzcvTWkt9V5oWdUFvgEzfke8rC0q
+1p4gsLfn/iMuociYSk87ZVVQ5iCn0/zdY28+8+CjWCKqe9WCHysYWN8HMnMA4XgW2AJ3kwYeLOW
RCvp94dUgm8FIOKYqv9s/nu84EGoHwLVtaULrsp9nshZoZZobN8ZA7pec3yK0fQeCaUhXoHMuXZw
R+Y5OZ1XEdIJ1Tyk3K+3ASxM7Nyi0VGALxUg0qAEHEAlQO0qQEEYAbTGMEA+nEoFHt2fLF6qOzbB
bFAAaBhfpI5DaOF9DKJzMJ+xDVgCu2kmoxeit5lkrSZ3Eh7kbR/9h/3xBQVazO/zqCMJRog0rxQF
9NoyyiF0yldtHLZp5JV+rsmTz3MecdevhzgVZB8O7ZQhB7OiRgWBs3ZjLdYLBIUblcYcIR54ydJM
bNVfkhEGLiVoEhtFSu4voPrQaDHO+yXpcurKecdW+SuX5i7kCJWsKLK6qRydLAWcT4I6UqCPFXvD
IVTepXzf6uaEBW9TvYECdmX9Bc6ql2rMTrR1kFNCmoC6TAcDueLh8t3L8TKDQTT5F9O5mscSHNKz
C4O3CHlvyIamDEibjwTF8swCEBTP02gi4bVWVu5GVYD45xUUPOJi2N3eWYZtF28SM9vKYcjnaU6i
pZawQqRKWeB58ro/Yn9MWfqB7Lb5soPpGRJhxYZJ5AhPgOJRLidvAqTAdBpZX7ONsa6ECNVnEpBY
tH5LfPLQWGCM5KV2IAzKeinMfLV9kDlOJynH+bak5I+jWZAwB9JbYYX2MXlcD7G1LknioahQWb6A
v4mN+BViZuYh7/fJAZJOTu0IPPrdQ6VdMCTHvM96Y6usOMdNVnpfExN1bzqFCmDTKSvqbyJWAFuc
2vbHdzOUG0wjuaZsHUV+fLgIT9jhvYB3pe4/axOaUfNgFfCStHnhlgSSutXlewgOENjxK5FQK/Oe
R0YSEpnvUGMInVJyEBsyQAoSfZtnbdIDaGh0Q/RwZfq6UxS8BjDDwj1qjWdHu2Q4V9LaO/iJfZRi
d+GGglPoOYCQxubAH0QekOANyfnU3i3dmsuFRY8COQDCNAJOgSsnU13VQGydtKjH/xdJ+dOw4AdC
zz8UDDswE4MtRAvR/bBnl7JkGzckPh1Aa5QtkaS6MsSp8dPQ5SifaQu2x3VMwu/h9jKIKWwxttZx
rytEmpuGHI4e6FpJGmYcE4bl3AGWas8JdXkn+eaNDL8JOw8khZSLWp2aFMj6wYLBHwtRuaZvAUle
gGYT6CqvniDj8jfr09hk+LyPOmp0fiayEpr0XkGQFfPiJqlcJuA7UwQvd50xREiDAWM8YykkynER
qLavNBMQ0ztbYkwjlOuluWw4wEGUJA0rYwy9luFHD+Sn6IpZCEgTEulWYlm3ezoUx7DvNUrxj66k
bfolHfHW13jv2jEpbQJIusmrWuRdZW2c3VQ52k1mUAP3UIRyHVOoTyDxGnQqI6HJLcOZpyF2nVeC
1oeNB37fMXjNtIDUOci9m43dxza72C31+89f9GR4k9z1xD+29bthkmT9rYsXWj+h0zLe2q7zNJiC
cnE9kgeLZSdYu4dPTQvGjANpxwS11Cuy4LxCOcaGQEwSA7ALGd18HUfBUnUi1yvFu/05z+d+zt5t
6Pt+6wVmz53zmjNsF9DaFZ2C2AtGwSgg1WfZA8w+hXxhrlTWAQAk/Uo+SvQcw0KpYMSocdEqHARm
tmYQqXyG8LtTjmf0IH+9rAvE4zFNgnub9e7hLD9BJ1r9Ex/LSTqCB8mFFbKz2zul2iH+xrWzXVEb
7QGYmdVyXpCIrEXutxNzt31c7JISRQiXn8YGPe75Xv4/VE4Qy1G5vT7yhqkPNASn9dj/Vfz0Kn4P
lkD/Fb+r5Otk9RRKcavEBKbPYkrZzcI3WpNjwrLcS/6iVeGmOXdvCxSKtmnSvoKFWrQUK82WHzC8
GYQT61+Y3MwlikDS6wNAh51I/2rZ3TOfu3T2Z9M0m37w6O3htq8ozIrNRTGg/+qKCGQM74y6fuhA
QxbPRUAm7xv1mMLnTAa1M7L5EqEao063GTiTVPkhf9Md5JiTqHervxaP8afZNS8+M3vr5YPNq7c5
f1/9wRZrc+yGaklumsD2B4vVdKbQdUjz8FHBypGrZKlqD8ytdZvVxoxUBhLMSybGcD5sruDXw0O9
Fy9Nvfvo6gW6Z7zntmXF9bveOyuM6+rwNMiJ9kVfeDtU1U87htlc9P+X+VkRRKSL9gYc6qVj116z
ghRjlfYTe9bC4DfCkEFLYN6dr02SOV56KZ/fT0V2MLcoO6K/jVYCamlIqj1+5RgM1sX3b+MJjmtq
XsWwN0mq+8GyQJ2NC3o52deVUeMBSN2Kt0eKPa+a/dslEq2x+FiDnHZh8JaMA78U53DkLMaq2WsA
WQyGsezLu1QpgE0YF4/HTSo13t16o1azoHPNKGzT6ahMtiL5geZf/Zpz5njYGAK0iQ9/q5+xkrcQ
9DVzTZAUzOUts62jR+rC8NggU4r3xqpiqJ7BfUVUmdEsL/ktJg2/oBCCfY8sE065GoqfgPShQSv9
hVY/NdmRLAQO77ouRLFpq3L5FprWK4tq1Dirn+zPG0+HhBL1+3ytEgBCfVm12tkcb9K8+ldckySn
RBSXCZdE13X87e0vW+BGy75WFeUHxpaP68Bee6qHg2DvEm/vGDAQ9b2PRjju1/TSNh+aH/DyjktP
I8ExMy4Ipn2hDv1z2F2vqr9ei5YG6LYpPhn5QLTTEMYcEkb0nJVHXPMTcJZOEwCtYBtKTN1pXGrl
anh/Bj0PbiO2MpJoB6Im3vthtSN+Q2Qt+F3CH2lg5yw4RdB6LVK66NZs5jMsstb/20lo+kO6/2R/
jRN3aaI9fBv9/jShBX19lIl0u8CjAyMwKtLzviMLxeyhpCmwCPMpOIZ4Bq/ohTpuRaEhr+aATGM0
WQWZ7LUYuml4hSh/jcL6U+brgYqI+ghNwhSo46lF/JZ5wVRUF4gbSzoe7tTOgkfl4ZcvhxNiiUIv
+ChRekl9kW9t57EimNvoASUlzXaqID3GpdAVkBn2xuWT767981kE11nsyd1t+g+jXruK6L4o8EBq
4RlNn9rt1DE72+We7bY0376DPo+kjothISXVQ+pitiKFwSC2ee74qH3ObTJqlksrKxHuXWOCf8Lv
Amj6/XzLgIaSRw/cW45iSFJBZYtMKzjV/ejjfaNtA1lFX3rifO0+6uavjzbijcRM+rezvBV8Z/xO
WUKP0oIyR16xNxXOmhykxHueB0aeyQ2IflRicRhDNyLv3sBSZYUYOl+d0LkFlVWClYjBH8wGiXlW
rGAouaKSc1wJXLDIV5+tLMugDxpCINPTmSeZxHtJHCkjEBSgXC5FGJvw0KHx9L3EofE5d24XrXlK
+e4eLfAqTh/b9rawP1sDtqm3yr40IBBmTkXWEykzmPL1PYQeGLc5eB6/U/34QhPhr4M4Axu+p6Qu
emQIuikaqWc1kmMdKdM65Jzo1FUm699AoMzSAnq3jwYXfucd+fGkASPo2FmnhS5nIOpVjBHFjNOk
Fr8dmG24vPhQ9jFEigb0Et3wdVx0pJb4oNydBig7Vxj1fMZan/9l9MLOD4cUrWMUeyVvSOyPWg3x
0r3Y19xx+tcAPxi0IuUyEJPT0aaFMOUurTE7fGS6KKJwr1rHOkTe71zABKQmtdisZhgSU8fBPd1I
jQddY5LCaIjPLzsx3DWoh4ZFVRztkVCxJn4wkA9/Lh/SKnahtewcdfR0jzBl6uATBkcS2x2wQFYK
c5WKT9deTYM4is01nzNONC7XY6LNkJtdZacRT00jeUP8BRTVDRA4b39N58H8yY97PLdM6MEKzt3D
VG+q3Mmtoe7lSTAxTCxADqM2BnQ/1H3f8AjoD/DzPKYi00+mxIeqatRllyg5cmI9oWnc2UXnK8Sg
3K4pqDy4bCW1uJfuYVujlgwf8GSXoRL7HtMysczQcaHZHvb7/vir8yAWmhCuKEKb6xu4V5+JQnrq
1kfqXVPfoaU9dvsb1NGyC52yeiY6ZY3gqp0CUep50BiDCKyAOudnQ26mALeg5YsrWq2zKWq4PnrR
53FKJVfeZjwO3wv7ZCmzGsyHTY0QWtGTehswXgUP+Y04fwz5vnFmA+s4a0HiK2WI53m+S4X6b1J5
UQKPDnhYBnhP2fwj6XSVn1bxZYc256WfHYN+L7SK9TNNiKZtD+dg38xQuTT1jevvyKtce2BvJKX5
jgux8Fa4Wt9Wj+ZM8gTas1V/NRtVc7eg+gw5QWdN23nhMMKkmuYAZnybkgrXkRXYNqpNA/AM54gt
nWumTejTT/zPe+8ojV/4gUy7ABVGuLEXLIOZFdrKxe3T7/Lftot5lVWE1ytrleKfErLwu+Lf+3a1
9QUCKa3NOa9XM6MkIRkoniJs2FMQoplVPp+xXvSTNiuE4F5YeCom2IrZcBRM/jsoFidk2yA6U/Hi
iXOPSAWdIE0CO+ZXH2mhPh8tbDJK51TcM6AAXHPKe0Kf91mySxsAj0bcTlewgxebbVdO8mTInN9q
iGtUqefTOR/Pv+J1JAghy2L5gM/UlhjSotgUbMYC+gbEVzhtkFJR2Aavlsg3L9bWGEe+pJ3sHqtF
wLmW0ZXxiOK1UKtDJWB8qaMhvnP0THhHZawzyobvodCzWccfwE0R15A++LH5HduRXtqJSrCMEEeP
Bz0TkONFZ7EQTXm+rcOyx0vAcgc3WRthQIXcRSpeA4rFRfrUfddbhpu4c110kQ0pLaRqM9eHPyGa
TdTT9ucXGSdjeH5PlPH7za1msOB4PA9wQLgREq+1Ky9Az2uhP/wDcm8QqdEo2JTfql0it8MwLb2l
ntDtZ36BGUOsaKCN/saVgaCNqge7Nq1CA1p6gSXX3pHBXUkdziqh9cccDfg12vdkuyhiCybhPMAP
J3oD14rQSBemj6MMkYGWx7/UMWBkQSTBriFXszweGPoCjfpAk48pvCOfeBeWr11Z/s8U5YAvVNAY
cNQH6riavQG1sB/P/lOOnKLoqVDsSCh17/ptqpgcmRfGv0bU+SAvB+HklTK3TVIj98HrK2J9aCpI
x/9Vo3feINz5SVftMxOt1Ko4XPfPMwglPOUjxvGLUaOnemwa4CQPAW1KJeVNuCNksDLCr4lsS8hq
EXxTLMpPZV/rIgwDsmQVCkKkTTNGxVXgZC1dLNTQC5hHL3d1pELaSeXgJ5R4vUjn6jEf6y1aweTN
ywVAzTsqKhGAFmbVn97egrEQvSTcuD8JTk8Nr/uqw+Lz4GVlJLbkh40FgQeYu5J4sqDGHG1FOGvS
7KSrfrZNtAWhuRXcb/HJHaxYAHYs1ngt8yd1xIk4uDrn9yj/mJz6Zhe9VwYwxLyLJdf/bZI3j1u2
6gHdalWWzjlwzsjodYtZZ0gqc6WAs/G1jf1SK3oLw4jx+mYx4RzeL3E37vxmUFQqF9shMrUsweZ5
fks0PcvWv/BbfD44wci5sl+5nDckrQWERGuPMZNa2mkYbh3WAMkNBZRI9qjZdZcIYoO92h0O7ETu
kMK1sCZiVnk0SbEeyjfuGsFeTI/0jMcKEMTvGrwEunNlpo/SA2wwxUTio8fDC25eBMrYYnVDhIeF
F2t5GimLSLft5wfRA/Tdw8LgoN4BKh+fGSUgs5TCNYfvOAE6S+gZqPcRtJtYlEpj7gV5CYKGMGWm
3Z6Sv5v3SPKhltw/hn7Lwo/XpKvNAj1gl25EK2YsFCH5uwRKDbnpMOf692NC8+/akj1ai02bmk35
9vklBxbZwLHlCHoNKC3NtaQqCixJkF2XxoEHFZlle0+eFEVyR6HH1w9ItGkswcqI8rwZSOWNfW3x
GRFlw+qPE+RdSZFogqOdHITS6Kjr/xpBhjhAug6WA5y6MRXaabsvYlftiqervEWpJIBZ3xmy71A7
IgjVRVanvSkUzhVPPw5S3b4pnaP1XlBSSjgpcldsHmJcFg0NtfYLdvJuyN18Q8H9I1caf+e3tl9Q
wOXVSf2VQlG5PQvxCF/Cc5S6fS2c+hJycGKyja6atWOLX9I9uRII1RtKGOo/GacOQKuhl0cLYP2h
yEy7pw5R0kHF/JjQJUcnDQo4InVRmIbe/zubhkjw5EgoriJACx+jvVclKwhE7W/97vj7BX+Q5WBq
2FuY/Z0jE/UYQ6SCMUaoZUSxdlvall7jIYzn+Ye5BKB/FcD5oOGZ/SXKAyMGlGWHZia6WZLDvV5V
mt7OnnV7CtI0qtM4X8YW3DuXraMYcH7/d4QUacu+w6yIZ7VCqM6S8xys11TTam5WOoUy+7XYdCjX
CwwaDtB9FLF9NXqT9kkKzFP29iN1S/pf+yPrduF+VTMDPZ1zdSbM2SxQVbAXNzospuGZAqDDAv96
vd5W9OnTDAJxi8SvNyw+F2FHs9t+F08rY6wlfMbYTwWapZln8QAI4RdApbCBmpb+XOHt63Zuirwx
lU2JqCBfmuXBMnEWdG5QmRgJfCyadt1Hyi0w4WgCZAWIjdzwip+UoTglI9BAsXmtHop85+W+D4G/
BcqNTD16H1X2R6u9b364diGVP4TIwIMiy5ZZp4tQ8r07n/Za2U7WzuR3vQzVihQByWUmcdasmDyk
vn/oeFhmmDZZQEuWzhfw2VBZYJhOFRZf5hgMywFL1gi98cn6VMd0i5fJS/2JFeRdQoNvOoXl0ehH
5Jr8BK/uAo5ZmTEpphsFZCB3YdNsxV45Ca8eGBLzgJ4NX5udP3DFr5+c5eepSRpwLDFUSPDiguov
k8ueTdHPu3oVaeiEb5O0E1qlKAc6v3AmaM3rv8+FQ7Xdq6zYYw0P1ilhThPsvHXzWz3rmmYDpZFp
o2KaCrncR4K2bkcLvDya4IstehIaO8D1AdcJ7+LW1zCVligWgBpgBCL8XJeQHmASnKckF09D8cnF
nX5Y6cLPSuXxr69j/IBr/9XeIwsI6WOP3IVg6l3TEBNs5/+STb/DXR5AUWzQUyvxO69R02z4mRoT
LqjlnnBoMXDJy3HltdwwNBC3hxKqQ+WnM2xKNcw+7+NPy1v1/KsPcZUd75D1DdsetStERuRj1MuQ
rgg54kaiMrF5sID5h1IpUk/aOx17SVmXTaUObNHpOozKUZn3suE/sCKMdBB3iXqdfJkP92GTLgQI
eMKaTklnbGEQkvziZbViBYNvIlwtWMJHPjS7N5GOpULsxTAVlw3Ulep0Vve0PxbYtbSUbNsmA2LN
2quDT6s9op3VYNutIZA+k+RRF9rV/g2ER1I4NQQsw4hc7p2UGTTFFC9xUrir1mHQpRRNd79QZew4
Yzo5kybNVpAFGHmrJt7uQ4xR1waXqHJGrB7vyD8vECBNrKIn+KfvlRvmpKfLV04CIk7nwVCoK4A0
3vWtexI678k4I7haCX3nj3MIFeeuQauz4pAvXnTJxTx7+vfUn2lfWZMErlGZJ90/x+CWuqD8geK/
VI0qOK7Z2dg+/Ud1RxTq/fZBUXKIYij5OYRyffBk3HmgBkmUbUN1GqbPENDdpmb0T424hnSGa8Cs
3obqW23KJZMlwrBJIn1SJqIVKnpBjGoY7DQahKnVXV+bZWVJ+cIWhFQ7ISzs0pKfE0Fy8Q8ZeYsu
tSEDWZbcckLmTZjPuofcuU7J+cslf0TtXY+4bzpbrOeri2BFdJDigwy7cdcppCSQhyv5Vud6KHgT
agTfJR+QzPqcPkDZ3mVN2DC/nk2J8D8C62NrK5RWu5RSJYlY6OHMZW1fJrK2cdybleVbiRGZLvJ5
TT2PELFvYwsNNqUlJihpkk2XXl1mtedUmiPkHMwYLRMFoDR8Byks2jI/UHQsORw8zMIN8HPuw56M
sbnpIJGkqXdWxkWG/bnWVFDPkT9ATY6mib2Hh/jl7mw0w5J0l6gzBHWVIZ11edUbMkHL0D8BZgbj
5nisOaa0gUZv6ZqUMQXSJ6Gcdgvg8lkHETJdWKmktn1I2Zk67wvAHiR6IbydttGCXMFfdcrbgyhP
b6YFVFD7eajr3zs5/gKtnjP0/nCYINQ+O/D9JPhfW3n+oX54kZf7BrBFAvhwZLkt4TLuJDZDWWWr
Wsiuc3lDsYti4URcXSd9Ul77sCqZGRV3rsASJTjMxH37eceiyJ11ZgFx4J999Kish8O46Aaata5m
fMCrc14g46qcxIl8ZUd1ylJav+MVdgvrspaqM7BImXjEWTWcrVRrUaNP4fAd+ySlmA1ffVDlOrfx
ZPdVE6LdXanA0ZMAwdiTguzIVxjWNiF+QMouxU9roxfif5eM4U7mK/t9YX/PhRSjFL+keEVstXSb
LtzbwVxUJe6vqb1OyUEuamd85Ve5YvHRujEf21CoS4uwvMjH9rlG05icO2KKuJCuNhfwNGeqepF+
VyuZht1bOYQzDhDAdg8URIPXH6rDdtL/0VRGtM+DQWpDXkHTycyQTRnVPlHGciJGPrSBApmNS3hi
TcIhLpgzdG2HU9y9fYCIFHnJF1WIZmQIr2Phpz9f5Zss1IkJ3HICeeM/yPtcKFrTqPOA7/hDmPF9
ibEa1neJtO0cgkd2X6F1SS6X41bahxKVk6XsRjWhvql7pxRJOY5z6TOAM++Tvs0wKHs2PEZzs/G/
zt59qOjyEKR+zSQ/9zXmMVf6/Uee/u7Sn5PCcV8izt+s2RKzTdBzo22fZ2UoOm/gtMbhbXJ30wr9
cPHzLkYbVHJsUUwS97iKNX20QvxmOiC/dMgSUriLfgoFl4gLZiXQRWTQm3EoD0xkQNG2QyXOkjFt
6wQK0pXhil2xdSG/2OgSEVdSX9cTQ6bSCCVL/EboxBftM+PtOVgXORSKHiFeKenpQ/SuTlO2XR1Y
6ly/fCxPmsdFyqrjeqGVVRlF8X+h+MwgMrbW4rn/toc124gWvFA8TceWiJ9J8IVj3KSVqjQ77s4P
HDLbSMch2XlhhyBuU2KfLE0QWbuevhvyTuVFcvcCGJ1GEGza03nshmawFyjg5wY1CFttS8zE/wab
k8ffQAOcCbX51urfr+RLaPy52dRYI37Z9+0Iby2JLJBSF42IuGLRxwjvSg9rssQNkBG7h/SQBebQ
svf9kymiziP/ahkWIuckvSucib2OmFeJa0KqZyrhRNM4QnL8oN2K4TAIKLZTCPS6K7Uy5SQdrSCq
aiz+1Gxf/REMWDE/khp2jTWFU4f2hlMo678vA4EWr00TcLQdk5bUOuNZjKmEsdhdydUL22sKcPor
DtC4SMq1jGaA16B3sAKYjhGZgwWPhzKfoxIcnlYqlKL6nLu1OxivGcCKR2H1oLO1681DD/VYZUy1
HiA/jt3TuscEOcJ3eAsUhuV2KPj45AY+neDizf3SeS4o6uk6Z96V7zwVnOf5PNT0GStnKh2Zk5/4
HmF9nYwYVi8qQpqzdwCqeEc4YrgT6uyrH7I3vUKBOhHkSf4G3lMkAqv70pbbVt4AdAknvo8rlVjD
ByxU875iBzppozlkOz1zpBbNs/yNR+Ilt/iB5wy69XFzpk9McG96EblhFJlBIYG7GctSgFKW4Z/F
1Onx/GoorUAwJbP+nAdbqYubFecRF7K3B9TgpDDABYRjIozxQn+Sddiixx16aPVKynYYyam0LdOC
X3krM2yGxunH6yBEt5w+xIkbw0lMLEDEKcuYplgsMa2vcVNhbeCyUBtjqPQvYOonzUsfbqOTc0jY
GWmGU0lI9LhCeO3+UEq9MBhXOFYjJsZ8CT+uzboCKExTkymCacPLTgSmVOlvrFg0/9zaYothli4m
kamUfTnHJPr7k11UOobSyMWQtAQheuAGcc0Ct80fRhI6ZMHHBReb0knVNIOlzpwaDJoKY1RXVNCl
9+gvfW6QAf5zzfXY++niu9tosVuMKiXxEmADh/jGhZDWNeZW7U/JpMflbP74Goi+ggBozbbRFcgc
sq8YYakIumLSjB9P6HceeB1qNs0WDrx9Rh/q1yrPzuwgVL/Avl7WyC+2NfGdlUbWMvBJBn2In13h
gRl3wnYLEMEuNNKkAJYjGdhU1j3VrHszZbG3sMQTz/SWqp8tS0vM2nyda7emPl5syPy7zDBShsIb
kglpbX0ZUVAsaF03APdCnfg4Hr7VUkSmll36yqi2uE9DfamyAe/xUDpolOk9Iws8mxNy+Q7BZEky
vBkBLdAyDHe+ZA2AFhHOLLW6KpIOs9Gh10G2+IAWycDQL6Im6NscrFjCFLY/GVG/de35VF/oqsLg
B+uHc9PQBwV4MaaRMoXjcinqtdXF6NfgIUMhDDJWtZXFPL8A9gBWiV5+ol+P2XlDeDOFVBLGu9IB
40nEq6sJwTA5M8l1SncJeur5QUC7pu53Fh55+lj9xawBbfmQWUZbrtb9Pu3xgDGc8QWDtFek8fVl
up49V1e9nXGInNeERqM2HstxO6vJT6TU9JpglWQ7gO4X0ia17jM4KFgGGHJMpYaHzBRk0MJiDGQc
UYcdJp3kQVzLqPhB9f1aK6Sgs0gs3oClZb+aDrvkNFkNaqEps5rfvDNf1EracoeB1HfMjedjo+Xq
aYpwTghDCDzd2edUuXwL+o5ih6saV9q4mkVef7ff+8ea5xDNk5zmYkKrm9cts4ZnfZBdBKjLxRK3
CHl0Tgr50xePC5u2+MRyKtrB4dMRMGtdj3S+e2nZE+SyYYZSyY6NHvCCKn72LibTbN4HTem293FV
+HYGLHYFJB50pCX591AenIJOaa/y1b3QommT5zG+V8U5+mDm3s0i0JBIzJIizLpC8C2wzy2wFA15
aBllwjDfFA7uFOlzvD/qbmPpobQN/8IBPJe7hrvgF31bFOkivSMukrMrcLr/y4Iwz+34uL6a3cdh
W/SkFoL6EmJ+NDyeFgG4XVdVf5w4zM74IR751lFSRcTq4jWB8V/Twbe+1uFdpUZA5i9TgqwQ7qZB
K0nWPQfKdoyt1s4ivzhUHDg88ZSGN4nqXzObRGlAPPB+yPkPNNd9nlCcxI2H8e/JPdrkLZZ8Cugq
B5QO2Zy1kpn01F65XN1UX+y9SVSD+eOmRI3nD4/OwrHnC2G47JTpUmLIIgbZDR3ySj2k/1iuXGUW
PzZn+BLzRcUyUCrdzp22/TI8/dQT8JxeO3VcU7eRaxStyRclLW8tt98yh6eDQBY6fKDrLmedScM2
zdHWoae4Bm3OhzVvp+VC7qYEIbpnlubRA+MACgx0JIqMeRmvd0TtwfaxTlhbujLhZGH/1mAyMOqK
SggVpbWOiATF++cf1O2hqb9JTWcbos4JmCTUU7NRNmAUWgdcNsQShcYMszcXvlyP3eYbdeJkQ8Sk
K3wOmWe5dUbDdzptlX8IuEkQsfZJQP0E/HNw1r+S/U7di3LPzte3YayZFKLpdyNwoBkChg5O0r9s
89w/LSx37mwznTLEBPWlQP3Mh3XdDxoPkmJp/PUJKuAZkYhddp/7dTjQmLRPnn/GYqDVoMB3m3dm
xW16K2g6gMRFbQFKBs6vqBmCUTer1SezuBOVmoS9pg6+6L/oM6r6/cr2/AZz/GVXsmBSR6vymusB
G1iYY2ISg35wd4SuOgbWbMdnvdxiabe0hSCK+kx5GaVpPO3bn0CAM+eCv4NZX4LXAeldgtbuKgYk
xhTkg3WHMGeDPlyr09WCiUwCNQF5kqDi0ziZ14q0Ci5KjIsN68ZXZmb3O1ze2P+e7S2SOYebk9us
eLrDsPEfUEnmB9CwEqSyGj8vY4z5T1duLxfuDSiXozkSAy5pec+52mHqBU0h2WGXhGPGga546No5
vKEZXxG/dDvbjhGLcJiP1OzIcVe/aPIiXvJje1ud3MUzwBHS59XSw86ifmeMpsK8qMzoj+EadT2B
g//RUsTLvhd9beYhSJDR/GD3RHb6P1p/HqJrA5lpyHN4su039zeILMFLlsaPWmqhDs629TNxP42g
7EmLns0Dr50SATTu/bb21pyc0T03szf6FwaKDRXoWOqLPEtLUW/f9bILwFLkKiLw5AQKJmxRowgz
22nBCMt8oWBpUyCdCdq0e7YYbekizbP2tUF0XsJzNZR5YU9MYZB1vrkqJRTfeDwqKN7OOgRuaqqb
YhgIQUEAEbCKQqhmM3dL668xOWfgdiOESyM8kN8SA2sS9wmpB87+/Af5CcZNBe2eGQx4R9/lrCvg
9VA0fHC9g2CeVQbcDCKrtNt7r26LbFjlkKba4wbXRhc8gr0GFu7rnI3ycZQe/SfVsklkMjOsYsui
nAo6bUvgxl3xu4Vzr737KJZDE5d3i0jnQ2rorRWZV1MR9ikur+h6yK5SPAlxphkQVoLthAPhYvda
BS9lOhG/7YKzIbgA73xCOtLlnu9Y6iWaxt0ZhqhAdSmsz/eKDFW+3B5+P6wI1n5Wm6IAzK8s4AVm
ejkTuLvqRZvrlsjmMrVZJdnHAP48JHkXbu/hn4Focnnii+kN99iIlVy2Q7YsH8vex+LuGHiq5rFi
Dp2rcDnLvdqlFqxxjPr347dxuFWJ0kRJeMT601g9Rbv08yxDvi+9dlzU0l7mnONSLCrK3vWOIEsc
VvhjwzZWSEg9Y/qilZ2N5hMfUzVc7/Bs2X7i51CSnWPKKiPWiRNw/tRsRWqcoeK0WIdfoAldui2Q
wlTEjwDMzq6xiXaGMq4N2gEFzLdTOXTzlaVNhRTC0ByE6/SL/jlVePAEGzOPDwkCWJnZYx1UePav
7O1IBYEV43QfAi7ZEznW9A66cAL7hND+LybQdyA0VauhXRXKJ8jtiUqlsnYEBQUhesyYPUoc0eAs
IHwai7vD3sO7MuT3HhprLQPQk3rAsck0XXBWyrBDswIoAiFwWffPm4GYdPqa4vJkvpMv5OTFKYbF
vcrhx7t7luvSA7CG+iXh61TGRrJWBfaxXnY3sysS9SZruy7wNGsYGgwTsWh4vMxiHk53UAQlMwQG
ZnYFjdZ86WSCi7bU9VjUpAXG9BIUEejXUJhBtBJmPdJZC+gInUX98ZHqI+Y0o3ns6P1d8Z+Cr9nW
Zge3nyxcFgTNyfUWsix0D1CbfYmj1JwR8B35aNqAu7CEiZuOAFEj4svE1DnNwhG8uSZvqgVh+5Kz
O+B5Rz8bVkbbOS1K+MamTbLGnNH0wwy81nvyWfPSLRleQnHxG2rdxI+xuG51L3tZ/K7Bg3gyJjhD
pyvnUa6EBiV+dcAfD1W6ZUgxt42/qFzymPZZzbovxO1jK0nfv0UCfya7IxhsKo9+rgNGYNk01No+
rNizmhwc73IXIIvzsf7ascaitzyQmgQBQSWIZexMEG0wlNhnKqgLmwRVdeR1FU3rZlP1EdCZaDO7
/wv8gP83uiK9UFUFs88AOdx8QeiOJtIjSBIfwHA5WAcVJD7zxC3QkAG5FLAsXxSeAfRvWcpwP5ZQ
BzM599eygWZVpJroP3/C1ONeLBhItc/AyciTynVg1HCJh6RrWyY5SZL1JA40YQPKbge/Jbytn67t
MCwL9lJn/HTRSWU8/wdD4ANlIaYm+Edj24YI8Yc3DlY2PfqFOfzE9E/1oiZk2ENCsaQrOpcjCVnY
28dvdF/zRjdsZukAWnGldH4h4woqhjFWxWLIHarziLvmcyhl5hHar+Es57WhHcovrWp33msdLu6R
btYYC9SSSIkRrwmcj94THvdRJIW84QsYv5e6cb6kEAuQZ1nBnzMD4594sVhAXY/+zdRv6x044Tlp
GAJ02SblfTL7/y/cRpN+C0LmsHfc1Z2S4PJH7PeVVoL+BB65CRqAK3qOpHZkyIYNiCt2jbGWy81c
btY2jycvm/5LGUBwZJrlzT0WVCmTKn3JXvuHDR7aEepRe6q3XhJO+jdU8cK/vYMWshQjdvA4VCAU
CIY/ViUNL+bcd5mBDq6JhadDyEPuzzz/bSPEc+KMLnmvJKecbsZbwGIax9XKDBFoHXqN8Qg4VDaJ
CIpJqKaUEj+nqbdLQ5Tkz3W6zGFz56ZkHam3Z7jUohQXacWWwnVToGIJVSjCJKBqQvUaSNT/y8Gx
2vJtyHlpieUC+5SUalwpbh1N22OgJWKUwk+Bc253lnYzdFbVJtsJ7vwQPD7uVY4po98N8T3gBm4V
XQrd88adM7Bzk7rk2XUaCRcHj7qzf1OIAiACE7uLFTl4+8iRAJ5dI+MB0QnwBiIk9FnG6TC7SbFu
Tg4xCgdKir14Sbygnfc5jjHPN51NCKKUcCmnqLSLc3+NjsB2QSQRrJ9J7rj0SLgiDNqnv9x8kgkG
+L9nTeESpglLSB3D4t/hzQKlIYj1ozgFszcPpzoehP1Rv/fkN1qWfzD4smvQx8bHkunlVglzyDpx
ApYmDIY7WcXhOVElXGQo3APdW1iNvIjmwGyx89/7mqjxfrXvgUekYodsK9EMIk67fXnWdfOSfRe8
nu+7Y2Otk9byAcdEId/tJ6sykH155or1j89U7XCcWSAFRQwDUPDaMYzhBNtPsjDF+Z8EbsM0spEQ
8hIZ4OOmHOafEQn9ZQ1iuJJ53VeZ6GJC8dmKQAwLqfJWmE33Ro4rFly05f8odR7KndeuJnA7usPv
yUCJJwoQ74LyRNPYj8FTIuWk6BAtI7dMGq6KJhjmlFAvi/n7bx0Z5Sak9QcOcvO4F9y4oP8xE1yq
xNr/rmqdM0tIHeIpnLHjztvKwTNOctfq8m1YKqGFVfrxVSPzRKs61TzQHFPnRhe/Js1huKkxLxH0
9WQdXJU8+w6zMpH30ivQqu8LOGL01qWp67yH1uuQv8Nlx+v2x6IEuczz45xjnBrBSZSYdrFhdHUm
ux3q9iJE7uLz94rSb2LmO1Qzq78qKbiVkZUvC/hLfG1dfDU3XU+zhcikqEw1rwGoCj/Z3igGg8sa
p7JRQvYaUsD35+8W/wBRg97T9O1bCUVsMsgAiriFyHrVwZkzwqvyEfhUs5fXbyp6YliEaSBT+8V2
UQnojb92FTCaKpywYYR38hFIr6uZBGocQj4rqgboPqvB6h9CAu7D1c6ASZWmm7R6smaa1ZgFBKQG
210IFE29aqz6zhnvUkC2eozfKxnCHG77M64csV/u7A7xB/ONitjxOss44+R3+M8aRH47OpNZH59V
r7etlsZ/XkgHXWW7JYpb2vvgkmn3ZJ2ns9rn8fl0URKjzWS6fpGNqcT42J3VtZEyNpUtjMBtgkQN
/xqTeRW02h1Et6hI83OYsWyYL5CN0xrX0WbJeUIy3Z3a8w8sPxHaelO9lJIRiiLx+Si92oJ4keu6
o1lslsP+CufB2piTHLg331mgcUVAP54Ekd/7UDOQaZV/Qq0D46nA0ONis6dteD0P/k6apFGZwcxB
m1T9YomxXKCGpdKUkCfAHlMe0TkjRRM2MOAzt6MxHJRw4oPoIyRsHpJ33KOrx1+8Ol6qngGYw8hM
1Szv0k7NDGeA4+npWmYWMJr7HZpI43mH8A0kwK5/sZlo4DL6fhAXZwSn2j8QT2tf1gOtKOGKv4hy
47sW3p2UzznGfnndnxAaD9MCWdyKrDVl7+EqImyjcXuVH72zaupp5rJaVj82MRaWI1btq8xbCOPY
CmjdgupP21XGHBPV59Bc+rlH5mdtbv9Cfywph4OZHqE0RozUwbA4sYptoN3DJ7xFa2nfHMZhZFqb
dogCQ7lG4ltO9NIxwSjxJUJytl8EvJhuyiBlqyhE4xX6Ov5g4EZrqcxLiU94WCwWDGPK+232FDlq
FgWhMPWjJsWEwfFbWM+OWatKuzY1tvu5QRENNxy4BYmpe4WKPcYpgr0GL3kszL7r11mGAwloPOH7
RlrSN78PlcXYt+rVd3oi5CjOy6rm0VLdjIa/uUD89LsQsRtPo1CfqeZQqFoLQZxYBydfynJf+sIy
f1EGzzSnpYgQFyDXittSOGnNv4WvsV2rOSxB3yZTtks1t+1kRsx5JuWELDEBBCgHDHEpZt1jTMKY
q3HmwKeR+Z33nIkyqo3bj25/84ir/KRkhxILus7Wt7qxeGbFB+VX7+1nvAKrI5jV2lKLcgGDn0HR
nFWlHEhgjLvrQIU4UvcCeBOLCy6dLbnCrpW5AWaawosJafAKr5nI0GckBO5Ve6ZRbL8co1gTvd2V
oqK1CWDkyeeHVq1eYfT2WS1cgFGSeGqW6/kqkEnlS+8+s6cxEiUyH83pbcvDAq3Y0HJbCZk7MAaw
QBROz3ymcOE3BzCKG+/f7s9Wb1VeGWsNsceiuwGbQb/2/RMcTQmnuPeO8oFkMOAHvxuWAa0TrUxx
1hTXPaxRA7KsVqX25m+lz8oYFS+zl4EbqVo61Og32AX8Mszt5Tbl1ZOHsCqM7l/wkPthBGE/UHng
uatrFIFcrkVyxBbEPLouoZOLyx2mqTiPyICFFjGBee7d14h+6lQeZ/tpeWTI46atSdlslvKpjoqz
rbmKz3HrQDJpPUVY5PbDRyXOzQc6gNIMGx7FJSHur82v99b6lNaHdxHc2Y4xrkZFv6hIuXq8aGMZ
kXv0ZvBFuTy5rHA3w4GYhyuILvMXKPgDOPaYaNTShuEVdshqCdaVJHaNnAlWW7wMZYyAMTclLf3n
gIt0uFizosrAFbRwq2iME197BSC7CcXIWIuaOyghnYMaWMql9H4yIUXPzNgYAgk1enaKvuVCYhVi
V3bc44Q0Uc6nomN9eJI0R27WGPwSLYq19grMWLReClyXTW/QsKHWs6vewzyE01OPda5NIu67NWGK
7/GNa9uQ814/ZgptDsNOlvEEuv46n42GkSOtYzLBkTbz0uBRo5DtdKOOBI+dipyMFMICflvN1pjR
r7pic2KgGySotABWrYr7S5y51LrtYws49HJJzAu0sMKFAVLkg+8pvl6aNn0IhTm1SWONAEjnfOO9
T9IKkR83ycQl+9FfJFutDEaTFkfeTgJ6ET90T2vj11+yvGYPslu6sogsB8xtoZQGRYwzStTSHRAa
f1Ro3xa7qMUIMdlUVJmpIocKeos9S4PT6znfqOAGQ799xN4JjYn0FnfVTWT7xoq5wrxNim825uUP
jo9B0bRGaKm5hXRQI/5+O18X4Oblr8MWCnyS2J/6ae/yqjPYNP9HsekajSW4hlfzexsLO7qU4njY
Y+bgl0WJ3dzczaKEIgJQ3AcWyg0hF1ti/7nBpO2pERI1eY+pGXVgZRjNDOfIShRNIQmuNOuiSHJ0
CMghFQcDSCSYKTt2NlJ4OC4lZT/qiSen7YJgPgcd2HyUVyKQrOYPsn09UQYbCnpNGZa2XtJe8nnZ
jlwif6uLgc3v3gvBmcLUCJlv+FIGUbX/D199YkcTfkFjSBCuC3nmktLOCStzgp+Jno+qZ3yBpePZ
g0FSNeICGKtO0uMv3eJXSnN/WgmZiua6Lv8SwENCOFeAqqP19bYdes1hEJQmAh9WNZ8235PWfVaV
RSisSU5bDEsvsOhITYM9pO30fkBatThz5NrkFADfP0IpoiNG2lXyjaZoUkmKqQSGesKhtKJ1Z4Hy
7eH3plgEZ2C5ENoi2b1leOHRjQQvv9PxquXNXuhYgOT3wH/GWwWyeF+QXbzQcqvN3t45tgoHazBy
xfiZ4Pj0iFqrninr9YYFj39sySumcQ90rBj/8HMTSX6zB8iNdzMdfBMWThbXozAklstF0SJktX5W
7sxfDAvpXTVU1JlBfytw5V3UsLSP7mEQXA2DWZr9dThiEqP97szy8x8H83LKY6RiCiSOg8LU6F+7
ShXX2u/OFeXGHDsJbMlpTyDG1wWCQe2PsxP1yEDlPQSpGnC6XBE2dmupx+41ixsGMA8A9fX5o5cf
zf1mBzVnZYX/d4Q22e21xUO0DDkX7u85KBNSPdJphF9kUSXs9rkw+njkWlTgw0Flv0XZTZ+gh7ug
kqnfjIpgBtU9brAORLnIUaYGVFfT8aaCK1lvpLX1G/Go5o1kGC6FNR2V9XIn4F3Ub6Y2PLHCxhr5
t2Yqrgnx21lH4+dyWDfXz26f8sLzPG3z9GfssVKLM+enWPOzXSRSM5216uxIHol8DXdL3zn4syXt
JQXn1vcvfj7P85EUnz//CyLxnlbuSsyUi0x75XEg6jA+Towxb4GyAP8BNLUFfCTkxYIgB9lGlZBa
rrvOz7bpppuZXTEw9VFA/UYtl5renGtt4u28rF6f1Pm5qYaKjme2snL/PavkNwk/tg21C+ktKh7V
3XN7pDY3ZLvDjWnvOumppCeOzUTXXKurjB93RRUBFyy2GJtyRzznDr3MQoqDo+ew7iHkZqDZcqzX
Tccohlt57qcdqmqMGB99en2C4Wm4aaiIVZhNc06eYL5tDST366FMM0eTlUq+fiItRJxxXenWtx/3
BR8GqUGlXf6DekYBhM279OfwgUVOxRz15Kik7py81Udvwbd6a1ePoDBjPeSbNEO2rr1Kow/7oToL
mOxtiKUQahILxf5RumF1USlMAfIRaHkZEnz/9y35jOZ0DFwohFT6IUUtMhmnAwnrOl8CybXo/zb9
V7qXY5lDY/1OJWNvBTR96Vd+LKzzzZiP2f6VnSL6dwC4EpO4ZXKBgtyToC+q0Aw0wb4WbDP6wLZF
oVW9hCvX52u4w0++sE+UkmvSeKD8F1tE2SsrVZC6gF4OEkT8suwTO1ud/QbCyIS4dU7lmEOs6VJU
H2yc18Zr4ezdHIyt6ZgnHLRUSXZhA+LGIEst/69Gw2qTPGe6xzktLfnxXLKR+YKRDaTEwUBc0uSh
HuFaqskbWg7OShOwR+JTu8mF9zHsdc4zol4XMbOwvKvKQySgJ3isQQBhIa2NFiTGPjJUT/TJs3Ry
g0pKW04WRoIlxtCgV7P+GZP1g3xyCAmik3wNlD/yeUP+7GOduB6r93g9nDEc+u29/mvNvC8nZ8Hf
guCU8fVtSunX36XW65JGhoUmckIhYv+Gylwe8NVVZkNulUV+6LJuG+rueP99hnHrG4WABSbYCOPJ
Qtr4i6yYiENriL4+TESPbET1mO+P6FCorMR7KWHam8IXebZF4r++CxjdwrmhbqyaUjwGTEELpmbw
0KWrADfxu4cGnY4IJWKyC+0Xzivr0jI/I+hiTIbMiOsz23WJDdRWB3H1xes0J5eaT5b+WRSbMWl4
IhGFOGYXt29c7Z0f2ooewoIdJOgSW4I3O4CBt+3XFCGalSDOt62gdZI98QasptkiqWUfDuS7mtVC
luP2IYmA6EjQ0rDgAQe05jldCR1uK31wpROeOq1UIlJqi7TDExK2f3r/ShYtVVrmbFu4t5VARqqI
Vw90FcenbLbLDgXQzDK502ptSaSyCMAbsNlJ31wafyYKPob6vvjzjRDWizgSFOXQN3/dedvuEhb4
jwLcLkROx9eC8rZQQyv4fo/GLlvwlCR8PuaIRY5tsRnNBgz5QxZNZWD2uhVX2IfJCCzNG1ztUpSg
eN/TXLpPQuoYkRN8vUalTHbDEwVhdOahIRChk6CvzByzF5bchQQGed8EBRZzI2sQwd/iPH1hkT7x
tlHEFqkMr67a3A1RhEzfMgagNIU/o25VfT3hDWK2EUFE+/a1VFrEw/ti37apleqwGqZ+sI4WKd9D
scwncHgn7fxz+U9/Ftw8bz7SY0Xeadewu9ao47n4pwquzuv3HbG7grtBo0NxY+8pNL5kvuXiTyaj
xEr7eIdR19nbixlSytANO6jX4nsysV+0ofrc+3ZjjrSwAfgmejdZqZbXC4A0D10Pt2W+QiUWSFxf
kpCnaO+3ucfgw2mHTZIeYtpqz5xh906vz732cG5Tm4/pWbi4ZPkfhiA53AkReqr9Qrl7dwrmK4yk
3kdIhBtoNRdHzM0voY5Y/eJ4roJN1X4nZk+gbJOBUorC0FRcakhunCEQQJP0O3mwaaDDVJF8+dsq
YiWb95KI2upWGxPIsGzD8Sc8NIZgqZL4sY+q5mhKXcGsLX+zZpKBCuiAiAQfpCPyOYwLGbkpAYUW
Tp96G0E/9cAt6ueDa9+t0br3IOEYYl19zBXqaE9c/hRelQVtNjk4pgMG4H9rzS3kQKa132RGh2bD
Ss0AfStkgceii7XkJfsV4RpL1MVmKmCyDXCdKGqlO+xCIwoQ9NoZXAWKDmmJU12HN0q0U4KkzosK
do0ZFvBFDLmxl2+eIRM/n+6Hf6l5azZMJTAsjraKL8L2ffolAq5c7M7bTiaZDXKRU8+hEZzOfbFG
H6vvK76OtMFXOoFVnlXDxiL34QJkLN7Xtm6bvzUoHivDfWTtEVpXlpUg3ws+KxknjQSRXjcb7DyY
hjBRD8Oc33LR9cyKM73zC+T1KnJSrWf57laeO4OIk5DfrbQKDnBYuInSc1tiv47glFtXwG35VtLc
m2/EZI7gIEyD+d/ugrjI5/hOS1xQWIXJcKofjjlra006V7jS3MK1Tz2oDqqleYgNW1yhiIBkpZiM
pUldGleHBflWsOHD3LkSZcBX25ZVDHCebG2IxkgXRhGpL44R8qs037jmUIHTk1NZ0azlAQtybiIq
OXjgfasBtuoKUBXkViQFBbIEERUl7vtYeNp76V8hFls744Dj8ql7DnKWmyIZTKmNTmCSkUPk5jfB
nTToou99SlOMUeKTrVQdT0jpE63NQ0FpY1NA1xhfQQvmU3X84TDKTR++ykNSXgh2kFqwzJ59PO4y
RP21lCi85jyDSG9jISNrw1/kaDW5FrZAWuijZckZIDm9j6oG/rgtRFrv+Ix9KgwoFGqijVodVv/X
0P7J+TS2zcyY3RoI4fLEh/SMY/x37+ahH+WXRN8oUjgjQ54ZWNjzy0n0rdVqMYEnnVUPNJszfBiy
VSSOSQDH2IbkKXp4BBdX4sXYkTapKuC5qvuw/RgGXm+CCgyvJjJWfNWgbAy6P8KOhT7SglpSUDZt
nv/qSddb23NXPGAEo6z454ihoPoeZH29rUzj1vuc4t52rFcRA/AT0eeYkoJI7fu7RJURkjLlbfZt
ujAu90GTTOZGn11r27Dedqk/BnmrkyR3YLQYv9zSwb3V9TRWe67EIek0X06jYBfmllslVwvnaqAw
1GZUXFJrDZAwXY5InlmbTiFUP+EGyuQsvFKfPqZSzwIi1m9mvJfLnLQdmziVZRzmVdxXBhVUr8RN
ccm4pobFOmK+rd8sxw8Y+TbFwabiDHGVo9dPSEGHx3OywrXhj5WomqSUNbO/lwNLkETtJ0tdoDjT
WOfTp6SSOEjmE9NZcP3X5vdo1NBJyZPXYDXn3QbIU/m5/4MV2jq+RApeANC74XYZ+R+o0viWGl6Z
iUI/qsyM8r8EVFb+jlh1B+6+KgPkiOcw6PHfQPFIpHIjAuKYtKJYMrh86nyV2KQL02ObD99aIFdB
L+hTRZbEPUb2SB1+rDGLB+eHW+2KJJCAxJrpFak2ZFwpqc5Pp+zwF72LDZQGaxFqEoqM/Co1Kk35
XHfXDiNXSkvyPsOta5Ju4d+KMeHjZ1xeTN5+berQcD4MRTua13R2n5/UdPyxV0zhhjmsxfB+rT3c
YlEFL5Xy1cx67UYPGEED3zGtOmXVUmB0g+m8jNfG2mWSmzw4+YFv1XpjNr6SeJ5MydAG8J6ff0Kn
r6ejx0Ffl06XD2uuwEnX35LIehF/zCL4pKKY/7v62Rfq/6uNZ94qV6l/7mZ9Glr3CC69QAX9DvQW
oi4h3BrQUfZm1D0qx/WdZzYhu6TdhWOGenGZ1exy6v9ruwl5mrrT6N2G65DxCTkdYKAqiuMwOVrG
FsGjP5u5iKkCvaYq6Li5Xxl9brb39F4xLy9IapMfSRYVsWXGeypunsN5bvRTjIuTnwbU5HQvxrtp
LBu8Tx2lo8XoqZtL2peJacc57BQ5BM3ckfzPSUGFuPA2o0kbviMZZEDLSEex9B0vAJoODjUbQvFK
2pd96f7rgSvfAN67ZMU4dcJtWMzao1SW7rB1AJ50WW1Nfg7yUmiPgVvbdmehRPOhrXusx6JMZZbb
DBqNFLiV+NI+JPr+mQ+S48IYLBZFPHchfNJX6MKeNt236W7FqD3gxyq3GkgFMz7utX4ok78DeD9A
g6b8xQu8iIa9/R0+qosgcoPw0o2kkCSqXyf2tKaIJSy+dQw6tdmAIY8wXxeG8F3NNO8SZE33pRMy
4yNVhGpcn5FAd9z3BaM/IKq4fC+b35CPoATRog+PegeslqJdTw1q9MB7CL+u8IyTZFpXQ1ANDN0d
eDCCyuk+95Ls7BwR/1/eoJEBj/Hd8Xsww2MXIvE1y/e0u4gWnh27XfVpns73L8cOkPMkXnd5Yd7h
GZH93qA4Xxd8RURujbjZePV4+dd/GxaMmmqNaQerUpzf5/z8+E18otOlrpkJZAEdnKy4dlVFO81A
T9zPVrKxYNXc5h/kCXldYh+bvd5tdsKRrFE1TCNIjh3juzciBMhqDiHgpG8moZfvCPwwCKaCWJW0
toNhiVM8VLqqxCvAWhW8NTJHsWZXhU8crObIuuxodqkkbU+rWJR3WIWMJFv7HwaMiWmkeKi2CWNe
s8VbfCAlggWsX6iOIoaSwAJbvYJl4xU3cOp54GZj/2AmGlLUymCZNRN10/FyQqIx3bdzaNCAJY4Z
T0WZGAWCBvjIZiD9V4iPTnxMhsb4tyWFiorXgXaUIZe7X6saWbdtJkedWt/McmPABFKmQifkQmu5
XcPvxv+iPCg+OYaZIJFr9bce9lEEKFpb8OByt0lLFHSIxYWRV+EZ/OXgVAJrJOoDMbcMuRbmvvVD
dqvGRfZHJEqqzJTYDSVVKLx8gDhodOX7+mOcqlQZRqq4sBdzdQw1aHqLtx2yUsU/ErPGGMWVyag1
Em4QYChYVHXSWr99CzSdSm9BEYtRV+3N9BKhMCyJqhely0EeLKhBHYTKCU9Av7gWYDjzJpZNAYmO
BeCEhT+BnIpA1DmXKNv6Yx/M2w09jp/UDy8C9QskrNMwtYeoBpWAuCiawqKiTklcYyv1sqc2RNmt
E4ZcmZduqo6ACJBWQmSTa98krmYyJEXJCyo7Y4GT7nqXZq8Ts2Y2Is+4Ezev5CLt28p9Bh5OUA8M
u3UD4MfDOqjs8yPMv0rxbR9buZSA0rjVXs/gejgNwuy3KSI0e7NZDiM9nwzY8ctXLHqQEZOCl699
WIWjMisnGs8n0//GtfwKnzxX4KK9fWgQ4pi2WG/K5P1Fw/pIOcPICBZ0q+rjnsLhkHSqUJP9Pe3i
Snyg27oPt0RQOXuqWvoeU9Qy8LjMpX5IgJ2daTLIbqaDdBKu28qnxQhDZYDzHg7UUXsq/SRU2X9F
8a/Ntm25s57gG7ilySDzj2aWzp2E1aHLRDdtkWCqOrlMHH4mjZQuXemx9C+PilEVhDZ2wZ+9NyuJ
X8y+fD0+vcG9Jd/1OAQyTDADLsLLdBHnLr3dz+OK9fRcuy29f8g9tMwKnNttLN5rths1wm/9eXb7
xPeYCe4w7PMTCOEq4rEafBrjxZ5DTOK7ZMtTzsvbTvL129yJnnCSmOH9rnY4Ob0olp0IGLFDwdf3
l5szohu5NdzlAxlXVOKMDVcRNJScio+fghA4ng6D4MDEK9Bdv3ItEj40V1emxY1u7XDrqhW4aDeI
y78ejH7YEcEmKwmsFDuV83VSfVjV+/LIgjVSvclRSRQr91Oj58QTlFyv4oSmSYOwRpC0B9hhSaAn
VevPEVz9gA24/LVHQ6YdpuPCa66OnQyKQVLO8KaJ9NOPGVS57oJ0iYefZ2H4+yGpEwIAjwNCUCSR
ys4W5QD9eNEFbRiNK24LA2St3Hy0qqu3dI956kgzVeulq5kiLBsZVUJsDG5a+XU1ilfPYLSa7tRH
0hr7SSCYlZFXV7q5MXUIRpmiUNP+lHvTdrlTVkPOtQ1AjyXjjWtSQi0iZxZrLm1IT78eH+QQj5N2
cwYnlj7WtyupmZhFVqKAuIggXZDlmOjAm/8FwbT/YN+197tFhFlL4zG6WH5EcRQJt2E69reNqKxq
Ea9hzUX5Qhx53EIxDeAghbuHxbejsZv9cjl3dicaKaG+UWOMTPsFmDgf1M1lVdK59NghklbsFtNc
mmtXq9SCK8IyGLcxT+Fz/GRhz1z6C7IkaQ/wtBLnQexC+rC4FIr/eojTPyztdcGh7GG/QbQ5y9Dd
dLulr/s0nRfNuYYYWVxH9gK0xDE/LhRH2sRs6JbMp5RedKfZ/au91MXAmjzCIkD0aHIZ9Q4v/zfg
0mDo8VOdP9o6bJ3CzZAOZg45CV+UpzmGYUY8xTHh4/FFcPeuH8wCaF6n1OX60xI3EIR40Ctn1F67
davi/FYmMqcGA1kgCzxglSVvb+JfxxBH4wZouVAH34uVFwgmPblID7fzAXiV8U2iILtwlH+ZQ4Un
k8FWD2BzzNzipYhwAiFtXg9LqDFETdHYbmTZickTcBtVvc5S34LOXhsk7sssZibnryZ/AhxWmDlW
AZ/3mc1WxgZVCVz0gqegSYgxG4uOsezN5fbRkpiVSsUCwU8Znkjw2xIE9QKYDzporQ1Espw1WXOI
2weRzWEfYVKfzUMZyyJjYuMpHV4h/3RItx9ZyC7enWxNhpH7+4enJUxBvJ7Iyd6iR94AsHS/C3v1
CJoeuQJxmGL7agjb9S2zCyBt1Ek7M9NS3M90BRSQ0hC6EeJmbHNFOSxwWJHc050XgXMJrgb6ALgT
R2r06ejfN2ifzp5+a1+Rts9fbJIF2rl9bfllOZ4tgHBkk2iK5XbXVuuZqHQAhK8uQvobBxC4Ggqd
6n9juTxZNwkn+PvOYlZf2RNt81oRDwR5l2mIA/cd+Ev+tWGXkAtt9Z4Y5fB2y3+qJWrsq97dzm5D
GUYXeYOYrPcx3GY5KaQ1SeJopYVWqZ+AhKHhaKadJkrKg6c0Sv7ZpOQRYRuKPP+Sl90ttUzd+I6Y
vm+Bdk7pOPSMbdsPbbAW4gOfkkaQCzHIw6Jf19LahhB8fCAVObOhJxMy5/BX5a9GlVtGWJr1Sdm5
fAUeXpqrHbFNrqZWoexg9/NWlDcFwxy+pRPXsd4a5dKga4/UpO9cH/6ZP88YuIZQwo9fqHBxFuQv
O8DvIZTr+AYgyf++L6veRjAqT9GFY8WVCElYWsvYZvrIRlcRTqHa2JDkWQfKXKb1TMzSrwfppuOj
uPbJ1pfhI3wq9Q2otqPizTlPr5zKAXhrDaTKuQ+WcYdP1c9W9UhbsdFzqIaFKMB0qg4kkfeFJgBN
rh22/+24LS/xlwTCVmL6ISS7tGFSlzDmN0k40Q2pyTPA0r9kG/6VpKRL02Mm1qJtdvtGirOJBm3I
rdAZFg7E2PR7oQZsfyLHkFB3eh55w/Z/syTBgmuOHvowpnQXv4opDRlRXmxlA6O2/7VK1NyMfB1i
RFT27Z7FG1QFxr3RBdpzI+kRUC/zslb/mMJNGa+RYkUs3k5jK2D1aIcEXkANEIrdXp5nfCOiaZko
tqfN89gUhSHpyjK0HjSGPKf1VKcPAEG9y7j9/+ntxkD7Nyi+qVT0w87bXMj/eON/B61YvTT4voWJ
BWA6P8M0ahm9xDMrwiaCmkNJysAQwFsdX56y/npoOtifwV0X/gZCy0u+qtCHesrE8k9DMayC8jZu
CZzNDV6Y3S28w+miS/x+yfFv0jLwQo9/GPPl0AWNgbjnWZPOjiLrdzzMFBOWVI8kWSvhspFkjHIO
6wJpBcfPkF9j3ZRwN5+59e0BUTH4z5swZ2+G9zKOgg3eAIikscnjepgVzfBAgOVb3E1Eu9RcbIzx
hkEAhiKdH9FfnPnuLQnfMJrWBSaaIPT/PArTSn/WpO53sSSZLHsbARUSKmhuEaGfl7CKxpDOV+5m
6d0f/jXzX1qIU83lpTE2aUxHNCgSgdjN6JhzkELX5qs6cKY7Q3D9G1YdXyDoKOPI7IESJ0PTlIe3
WHBSryNBtE7IGf2l7UttTDAFvSghPzjcQOBrluXWgWDq3QC5L+fOduZu86YYZ2fhsmUC4RsSijQx
2HLd2s8Hs8ntMZqMK46Zkryyrokh3Zx1V1vJkQQIHH5w0ZwuORlrOCDwLJvV4IO4vktYkoa6t2sb
Ee7AISA/BtoX66xZlzpmlR40aMuDCFLGOmWyTAT2ea91fnpPYpytCP1JJ4xTj+5yJxx0im0Al5Yr
Q4rrxL4tOsN7mnuUoDYwmty5b4AtU1mSANorEiLPJBld0SQTSiSC51km+JZAN3ZOvvOpAKPq7GnR
uV4POOU/Hw6oQ8osBVLevPwTVjiLQuKRmJnpAClJTAPq2i+6S/cwQYeN600SY+QdAsNwTnk1ul+G
dNMcXORe96zrGhc+zKnknpa8j1xXskBfS6HGsV1LKKhGCYcYoqAorWUCunj82pOUf+74g4dD74Zu
7jgcW1uiGjn+XBVORr+c+qZ8ERLVgNIZH77l1dvMhCnifKOSibvdVMhNt/qJ8Nfcc2SLBKjUoVcm
UColpcBLhfTaz89phkp7JHAG20GR7TqFfMyYfvLEKSAxQc19MrbkxApK4/HSXM/rNKbNVAwmcsKP
VhNyHgYnuqpZycCi2s5z9Me6d6tS1gGQCZi8R7cQc1wPJky3UBdJwfy4R+nKBPGqYo668EvM9OxK
iNxe/CcdDPtFcwSY7sJlvNoDeDdUZfYehxV8pUnviv4nAEQUjkLn1gbhh8gLyjy6M9B/2pNNAsqt
A700af5ZiCeBg0OtfkEylc4TvBt7u/eiombB6tUb6m2qFKT4ShqEyKGhbhQinOzpUlaluzZd39UW
YhDdmQsYrWaY7adEOUsXZ2ymbzw89kZpCABfv1JdKvhgavfUw9aVx6AZWY6ctt8FDQDHHieNq+NV
VhKTvtvxcb0aLsQZ5H3BpdkRye4MZ+Vb+nidHfHcer1m2twt8F/B0QlP0XdALI2GyKOYZgxFJBcd
EOIlfusNb7SSI2FYKZEVBB260eZ5a1w6Q2D3xyqCOgvm42XILMFKGbvbupZsZJXkls3TFQkS0nK4
GUzo3FE8EeGg57MGaMKqyO1xT/phH4kNFXlV/EQTkSOcEr71xkz9S1buqstYEPrYjUjnZzSRhBlr
YyVIoyAcwJxAaWgxlzJ1uFJ0Wx8WVqhn0mr4p90e89lbdqj6OkRqfqGRvoiTCMyMinS3NL5JdVCA
NSRachMoOoCoThEEGtjSqWfNzUkxsOCcYuZvp2LQ8pe3iUR7rPkkjPV69yhRIb7np69kKNGQmnOg
UZsuwl+PEUC4N7DhdzRxwJ8u2Y2S8w+5XX571qMsT6OOBcDMRORd8LdRLjuUvtOmeBm0fkO42FCP
ruzH9zM3Qw8szrYBQBey9mE1o9vD8pKz+qN+UusjHqiKVEx70r/rFV7AUhsBmn5/tU8hDgi55LRt
OQGxsCg6NyuIciXN+Oz+DdQDueUjHVx7h++rvIsBQ2EfoBEgZgtZ94hSGR0ee7odORjsSvh/Haov
K/xghcUk7cdlu5xaqRQ3vifdCGMp9Ejkkrt/23ozpHU/392QJxHYvzinCq4NHitOcrPNlTDzcRku
bDyuiBg/GU8kNEVLH3fGB+J4e0JEPveClj5+45gVfuIzwAGmm8tNfR+KIQHaYCEQrUlMKrKv/VZQ
/ygzrpExUj5vM8LDSO4CWo777p5KrWQ6GIr5jb7Xg4tG/5QYLUxjVj42iinAlZbCap0s2ndXoJB1
5CSZrb1XLF69fZ82b+5dEgI9IG36GZG0bHQeZtvSRXjbPhH+Lrx/+Zv8hgAz5feSZbqaVBCe85fj
ko1jS9ejWBuxN8OJsmaAiM8NYyTpZsL4ggP6A/AQ6gxQEnD3EMH7V0yIF0K6xJuvLFSSVDS2QvuP
MOvLTzGgBKy7/egUb4u6epLAvoKu7pWoqpja62WIqEnNGm5FLXdYk1d0xCZNp/MB55JH58c0fKBk
PV4GZjXH9qRdlqEsoWipOJ3eM+hgFcmRPMX+VQHnEP2m3eEuXAy9kqLufjYHqLX6KjDGJpBng2PO
A6xXP0WBZssi73hZ7EXIkupbO9ApBtuaV6NQ9ceKjBWAOG1tg7ZrpsJRIDGcCfgCRwfgbX9uJKfN
Z7XAkPBT5SJCgweB6eD3hFwq7WSMy7TdESMAwAyodH/FROstJ7wRx9gN0GfmPWrLr7dvZLxJrhlP
PFtR+RMw4u6CzsZ5mv4iu6YFcVpvqiVgjlC6cGk5qezM+5JVwYkbgZpi3fVEASmBQacOQGalRKlC
wPFjhfvgSDkBQ+/J9xR+Oi0y9w0yyKDABWwfWh3OgR5cnugcHmeSr5Ahv8BztlH/HWEIfOkzmoaq
4vGhMhPaKz6BbLe0Jp9rArCjtWqP6REWe5w81xl06T8t67fCLyRP95Sv4AKxVWav5PfdAO9XK1Fa
AKBH1J2lYgWDhe6wNWg7HIg/39j8r59nb6SN/HlJCssBDWC31p5X8jl8zV6A/LH0YsdVDFEbgawt
knaI+ZD9xin1LF6JZkxX+rQ6QWGBiS3YHalF7Ttwtnq5+nVILB8cKWsRO5GD5dGVObv/Xhk9EXMM
pwapp5SLMtXrxAJdXFOlox3LM23n/p2RccymYRIgQdTk99MkClavUvw62m1RarGRxO1erQnWMlck
781u9ZYCoaGgGgilXSEvBwvzer9X2fv8igY/zHdkOb9pxGxvnzPVKlL1Qsd3deS9omDCJDgcESxf
c6eeShrOCLLWoOpW4ul0LVfWYIWXM6/5yqTYblvvmoK0ZzrrtYzg0nlc6MnTgf7T0jgBDd8dN1wv
3FR9wCcfV2c4JvvB9W4KKWCiAV/v/vrtZALs6nH/61EOt80JUxLyc2LpZxm+RBh0lXezfobuudHS
5AuGyCs5inkQ0K9W1+MJYWfgGted+H//sN9w9OR7l/61yL3U5g1waWxWf69y6TnE/hHlh68BSiWO
r0TBdgax2KmniYcBU5xE/goGubcYyQghgr1p1fzza4cc52x2Yx1dt1U2kXLgDi8pTnuNL+7imPBu
1qosEYeCrsS6DJ00/ob0J9OHo8tNHTessTlizyRU8blAFGCUlKvJF/Y39aFXNy0+uJkXoao/LGx1
Kr0cCQCoOrv+E5uyLb3anb5m78umI2bdg9gW8pDtsDH3fsFYvh6KLFb7/Hj1f2T9xV1LA237L9Lk
CqiuOWMw6jEBWfe/WYyBKfg3xtfNCL1ZM56Tb6sKrH/JAydz5MAMsd48JZepErw2/dlmk8I92DZ/
70Dwpn3E9I9adkrVFyQkrdQ0+a4U4oDikRE4Q8StEBVvlDg880CMxTwslnjTUp9+NfPQ9JiujpuK
s00OfmshE5qs4JzABWaQ47WePwsWv/K01Z/3clAwarz0PiPl1nrAcw72zb31bRPJY5aBJNYQoNBg
Zzet3sLmQGPQTHBpVJIJgLWBBQXL3XdtprapNHmiLRunFsLE1i6WlTteWkVnvPX63M+J8lLoOi75
WIp1vt9uVAUTfcMK34zsnRpwjS0TBYsaNk3/9Zmu7ZuPZrgBxomdG7CXz0xcRMIuRnl90vK50vU1
SqBaXQNoa9b3F7NneE4T/+mvAQo67i8Nf5MKdQNufqx7kY3QrxMm3bF03STEOJtoq8sN0qIJHmxk
mtok/4fmP/kDy7JVwHDnO0URYW2Rg+PMuUKeWUBUmJew6k0sWseGJbv1cBvavNVBiQv7IjWCbb2F
R7YZWz70JWyd2PXNKmYUMznktcfB6YProJUU+qnL5yEJj5vRLUUr7i3SwBTGyLTYMDn+lIPmVX15
6OUSlHOeI/5wn7OWnd+xYjVU7IKIDHtIBYxX3TE3arFq8L64J5kHdWLLMIMOEMx8UI/pexRreXSf
0A3GieRF9GNjW7+/k1/5/1iUDSAF+HdPJOK58sRFP5ban+qqlUpd2vQJA8XoXMLjzDBgB+38GUH7
6urt+M/SPqKIU/keahC8/HUuKzEv1Ow4jpmVMmPhABG5TwqbDkv/DQj91NONq9bUh2+nP/f1vdoG
LfpavSKPOE6Z+EA4chcdDMhdrapECcnPQGN+UMyUO0qFpZ99OeNwB+xTmzwoN1T2C2j+Fmr7jboM
e6BM+uKeu/A6nT+mHSXHELUHiCRYH6UzfMuuHMAl8H1JUhMwz4cn8nSk+ILtDqVeSW1vD6s7PqLg
dOdXzYd+zHzE45GJLSWiPOQC2O4vK5xv45/YT5S5VNNJxPwP8FXpnAHhAtOMJfP9lAjT5ef5NxWC
iVRw7x1QxJ7l0zcNti8A1bwXmRjlWRPGHgGFeSOmek9+Y+qtwBLnaT8J4W6qkIJqAIKcCstGNihe
JuXoUNxfqDVXr7GOP/e2ltOd1/1UWO7fTVWAhXXuyn41zyOoOUZpiwNC58TsfnSM8+O2CgJB6VzK
kVU253kz1mp9GS/3BdN8d6ENrOk+v6LWLCCLko9/MVssXq5o1v1FKFBhzVBR3KUQCDHXYsFCbEqS
z77lWI9uqB6kEt1omXFbwhg5tB44Yncsb6G8vjv0jnQS63o5vxtojOxAmlzDzSuVoscORC7bz7wy
oJp8dIHKKVs/WIxsE32jv2vOKa4doi33Y8PvWrM6AdVZdsgftHtP9GATrMf1golh2VIQU0rMmEud
siXFgu78/fm2nP9ozM4RQicuhP/4cdUdfvtLFMiHD4/5Em7A23dyrar/+xC3I8aWVMEwUDopPnnd
mY47XZsKM5S5GzoMsNmja0QV/pVif5vqlcTL1zOzblN/1eZODNkgua0bguLw6JzArRQ0QaloPfza
L1PwDlwcXoZ7yEnnTfpaccDNR+Khtv252GJh/7k7858F4shbIkegkNCDqrKpUxnf/BT+A75sFDz7
xOFPr1XYLINcRxcPrq6esC39oPm4zS6zunH4cpv6y1TNG+5wHIO/5YE7RpOpBZ4xy74Ub7lowpbp
uVXtlZDBsX8QPL/AliCiZRsmNMHsGDKd7fdacbYsrWYkRVRyqY/2oQ+n0WXEZd5v1wU4qWNY86nu
NE1br6G2S2u0nBOfaCErAKNYuDco9PdTfiKWdC90lh0g0fP9esW51sr02FJC73uGqJ+nkKN2982T
RcOpG68UB5/HjTyZ8p1qZEobgv9+6SZKPhZ0cpcH4moiYFm/q9OLRQyJbN70GL6/VxhAq8xQnunG
83UDJATkrZ/YFroX3/VcnTnHLWcAuzpcRlQodcmaPGuppYHc0NQ+q2yCGVCFAXw3ffdnOrHl+LD0
X9vk+iPBsK3PwL+xkE5ZhjRAgGrqAgOgF9Gd+H1HAUD5pV8TAMQFlg8Z7JCkfX3dRjQX6Q9yccwL
crZyOHnSUURILOwn6yP2VwS0ivCQlOfTp/ZLljKWOw7yBrzPLqEvcG+7jVl0etKd1tIbmAyFrYxE
RF/j8Kk5oKItB/RASD+A41o3vkdWLe2Nndn9TZM4TJEpzKzOfma5MJQq3UseWgqTVh+qdXq9sMf7
e/mp7CjKU4DN7pe39RFmNBxTNpYq5pCRaYX/6sAfgIWeJo6OLTL2FHL2c8BYwnSGEpUEJfnv9Cp2
xzwEE7K4wBjKhrRym65b1vchHYkn6IP7kJl7675WjAvP00WjKdKUtZVAweCYtaFBotO0qv0hJtCt
MxFpqs6ZEor/H4Fb0X37If9d7qM9KIz0Z/hUZ4eOftQKxLekWwR3ZV7gGWRK9ElpMr8KUsZbJzhp
2tJPYCPJ3MtJs2a/igA/4FGHF84JRxG30v6qvqor9OTLGVRF/KGrqkCJOxJeYqZd7hKItk1DtJgD
M7xt3MzxnM1TII2APWAaoQCFWE1oXDPC/LaiE5wODGA6byIZlbpBznhPrySauSpEvPQjrD/RXuNg
TJnEZB2NdWfodx5gfNv6gMl5/Th5bEngAhQSmqiBVd3VgzBaCdBp3pbFNCnA20JytFpujfbrAgdR
PLAqSkqGoohy+8rWEYyd4MYLg6UzT7atftoWJjhrs+3PRy6DkpU1ZbVUGklNFTEAKawanpBrCA81
v/e4+5spTRRkewqPwBhg2PlUx1xRb73UcKqm26WBkHhW0ezzhxlwxRJj4d42wxtIDnREp7IcLizi
Ovx5vM4YDuIKyHny9dDlb9aNBmX55c2q5qHeV4LkXSEsseR5/KYNcq0GcQY4o2hL1lHXyjj1TEo7
JX9ClGCU/SIH7Kh5GeOU2gglYaJRsB1gVkEVXK+tlWQEz3AOFT5DwzG9rdiHGKX3qzCdm0gYnZuZ
aYCFdgvCxmZ1FiaKE7W1MNVOwvvH00QPJO4YQ15izxjgqYUqlriUmzOmXL9T0T8Mpi4+pt3FqRwh
y3vF+bHKtMr3lUWiaBxwDlEveJtUyahawlkpCGPTSiKCBoN2krugyGR1K8wYGx3W3ZKka85wUyqk
Xu0w73hqNgg4yvrhOuCv9DQ5A0lvv/J50zle1lgkOmgfo5CWfMvCSKzSwzTsfHW83C38QhkqVUNn
K9+uW8m15EYhqL5+hBBpmF52eoYnrNXwsjASBo7LggitrMkcs9gI7Oxw/nekqW70C0ZNTUSM0M2E
AKbXvwJ/D1c8Z596RO2mkkKN9Zv/2N2HERPKlmz0jiPVEQDRnnfGZJidWzm8Na2/+7vCGpS0jVi2
vEkYucSi93ZOASA1JmVN6/T4+ZGsikXwrFIRQ6zU9wKrJl057+MOsjlE1vdjnH2SoGlx9054xDiO
MCWAeakp6yQMJcLkMm1pRIjfi/Wy9S3zpegCffGs/lrupXoHNTF4bO5F2E5XeulNOsculkWk27cr
NO7wp/85T6ZLYewlc+dncsnRA26EZisDwUJxV5b5T/aU1O0kuv8KOlYCr5yUbXxxec3YGmuSCSbB
etvvC0gsGLr8pRVcVHAVGwIEKXYi7cPnGb5FBScL6KtV5faSH2ppttEtZSDTrHoamGNpT+BAJYYi
GDoim4CL8P+WLnBUtBftlfPQNMuiaOYN3HiVWSn7akVB2dFba/8geRCsvQChFELjTZXX6io30Pry
N4VpdgPEwbH4UzbqsyNmR+nPT7anUBVNZKyf2lAg1RVzU4A17msFlF3c8J7KweRAdFn/VMbKYZeo
3jNeYuL9UI7IyVTGCQu410t5QwrRZQHGo46aTriOTsh5I+kkFImE7fp5ufwqft30KdzcSJ9e0Ss4
GSUaoURm8V588lhYx3wx8yg21hyOy9hTTPc4rp7KQUNeref1MR3XMoMWgkoyEtsFfh42qSX5gPD0
rjZh0SFRcugpDE+XrsJ1GYiXxnKPFzHg9kMjY40JDs9WA0B961cBzXbUS9MiUtTpIH7iEG7R5bbY
R9o5bJSIoDNsEnH0Xb9Aosg2E6Rd6pFgLTzYRVYoQcAqUJpXp1BWEwBT4QfkuC+TutulSyOVgHld
DuSRpvuIbAPf2GyJclJr3GvMqVUHWKVQjpDKvEEH7NQOjkRcXnfp7JH0EUDSOfq1iu13iTB+sWEw
16VPxm/IXWxVuM3IduoQQ355ThRNWy1fL4D3hgaKXpyDYgoiI17vCCisb57kT0nuHZvHdJp7ksb+
gbIYMs0HtP/5aEHqHI1EEUP74B6khz/bMZ1SIU7Fun6/w016zYzkTJTPzfJIbAt74HC7NevBXnoh
VNkg9NzEeS0dOZMXtZg3lVWnB+WkWqvo2M8TSKVr/PpRwz01zpjATa4LYQEOfPrSP4gkuLIVHWwq
iGIrKyksgwPwxiLkPGVKt/aARyvt2IH/e2mB5B+29wpGJxefMwVhnZ6qgM8Z0gqqumDpy8TBfR/4
DuD9jcvWmGmJbxaxUG+EW5ylATWdPfTqh+mjAS1BOpn+Y+cefDyskxVW6PHn2vRaXekGC/meQNbK
sMLUKatXWW6VKdE7pyvsCInOP2g7TgIbUjoRnvjpnYIPw3E1rRvHhFAAHd0dZZd3dJ4NPTWT/Ode
noXPul//V4mrGBWQCMPFRYar7ByUa7u9cxT6g6H0Ku0ok0pkm9of76Zheem440jDf02hNxbJn84g
0pXGHfgIdj5BXReOL2LOROhFY68hzhPmxgVTJc0lVwLIVJr9pLMTGcUY+Ive/nQMOxb+mtZWLo1K
qSROBU43/HLFFwYiUo/OlM+ycRyeRbCCUTZYXfkJ7SlZWGq7nng4VpxH/Pm0gz8u31qxgraTocqO
E/zK6++fXNdtNiG02Fmm6EgFhwem1/T+1CSXCwmnDPoTnZGJcadNQgSQ2u3rv5MfPboq52ZzDQYx
Fusc97RQ54KW4ZHevPZQwM9wSSwWiZnyVD+Pk2xxNGPppkp22Fb62NEu45mUTD7SCG6Hn3s8oqLs
2uDWX/tRGH+kP+Yn0s0Y0izxi8cPxm7wcoLSUc8ij3mutRMjVQ7RP6uK1UhSjzhqH2y7Hab2E2NU
9t1/5SELtZSXdN6d0mVcupQdiOuJyYXD59TLm6wN5/qxjizEIUh/jakzl1wBcZsUpGoFesgIGKd3
eUdZNuj5RgltQIZxuWvjloJNwDArhVbp9+yLQ6QDr6U+J1Wd4zUHR8GW8ZREBhVzTlJ6+gFGlcfk
5qydPT3jJPqq5Hku9PSNDxD6uQKnR+e6+u2kbdTmYrq3KFvJHb4eJ+VFaytbt5BTbxUhq4kwNAoi
6sallv7bxR6muH/Vxt1TH6rms1828m9pZJAwqFXciV++ZaHs+oXVgImTZ2aRS3iaaX8uL4SUd7QE
PV9E07ySSsdfEnTESeBhXGpUKiVKDlzmSXvzaoHajxEOw38IPfc9opXYAl4uBkupfNx5HKIeCiL9
12w8J2GRwj3EI4hvv3CkTmoqSh/mWaJ4MtDkNj4sHjU4hR/B6s7z/4gwmlhHfWbXkcCwkOV8a3VH
fTV+cgwnjHv+NkB7jt9BVE1ZMmFQ7IKh/MQrF9m7hXdOg6Eqy8h9WpcaH9NhDqwCdW7NJ6m9v/zZ
jC4odXFLPQAkcZKyJuV0ZNRJdS3y/prdlWCw3jtqFBh2fpH56gxF4SKAB+DI2JyXp4koVkDuCZFn
owf41Z6qh5lCMqBKOZ2VtcxGFMs+9KkOEBsTO9zE7GyZqnH88qi5d7NTkYf9odG0l8cbyeW/+bpQ
OgLYDOs6xuW6x8ijzTx9eLuAoL3RtPxSMvPZ3aMMQtoARZvz3mE0sUVuYKlcfGcdA7QA5lML7isR
+B4Gv85f04QS7dvjTUhmjQnMeZbpvVi3GhKL2y6TK5LJyv1PT1adX3CVL/9FRM97P+C3wuz525ns
o5u6NiJCaQU+L5pzqvywNNB5txUET2px153AJ65sMQ1ORd6qYiz9YqFbyO62lAWgMGq+XvnLBAQJ
3bTv6rwz7XoYoZ3Vr1+ksrlEDPgVIN8NXvwztP1bSGPktQ9Gd1XJqIG3cssMyjYvX6srxAMrP/Uj
zPaUV0P8g6rz9xCyQZ2kpmcMKdCuCsUKZbywwerxsyetR4qBidlt6e1akpFwqvISXtQVpj1k1FT4
ZZSvQCN0BiI99TsZAy1mUCcPzaEz8vYQ5buH+KI4brPJxEjGA44TBnz6xO20Wb5CfGTolAy3re7D
jjV9AzCvSwnEn2QEi4lnWkpSrvHct5CQ8afkuP6kVUTb1Ddu0FQ6BmTmW2ycoSoxB/bMhJVgTMxF
FarL8O/9uvUKbDYWpM9kHM/s90hPlFX9gIMDba4WjxBJc4bkcaLGzwXprZowFzbJB7kIF2jaAS+L
IpaJBxK/OSRCc3QhD2pqfSuVs04ji0XCKRMtIH4iXcnqR2JTYEvxHpAordVmnz2Rka729P9JLbEm
99x5+Ym5CTuwlzqt/UzD8xtkM7Oma2Rw8axad72G2EirqQvGYIqC9cZxJzqxtsW8+dkgCU+gtKRA
VqFMpmXXf1Xe5d2CdT8tbjtxLSPl7rnRs8w5yDNPH1Il47mEnB4iOehjJDh78MhJoimYJ2Kd1agT
LYtpssbJPlzP0no3Ldwnu0e3S3cJ0RN4+I9kUKt9XJ0ANs2KJ6MkMiYfgshbvfoWWbUHYzddFdeN
e0IMXlVK0SaUUv4Oq5Ei9ErsxogQJ7/Qvtu7LRazlv0zrYIFfi6n8ShmAt5qZ48/NXeWykR6oL3w
U3L0TEhGTQb5MiHoN1cjSPWmKNH3+1vQc/Fjf/tTiktrPcoRtcImsstQnBCS3IfkU+mnSgP961tZ
iGOiGs1FcUUwTKnI0zoPV/c3gapy2ulNSWWm11TyXsLR3cVVCUhwTlQKTejM0CUrXHdtU9EEOufk
m5OlU3tz8HBvv2XOp8ahmbi2yr/avRPEq/X+S4VAxB/kvshc6XKYAmCjagxocJPX1K599JY4th7v
W7JUetcj0ME+APkIyFxufYo5QHpw/3fgDN2dKHdEWPb6da49ZRkmscsb9WiZvz6t8IIjDnnj4LhY
/Db634VSnyKUltffVikryDNmYYWmb31IF9hQ/SHO2JDv0T3eQCjFVrE+L0qPZQ5MagLuBQFbauU4
1UL7yUQizkVeFCfkkyrUcrSrYe++WiRSFUQCEWPN+zXCFfGx5s3esLeRlb1RMjuJyhlGN2EQ3cPU
iAgcV+Lx4kw0UKCigZE9f5pdgoNH7F9rperxKlSOCD59aNI9CPv/WNmi0orCyAtb80NesEJnmPas
ia99kRC/nCNlaoJ/PtoKpdYACi+tJqa27V4eJgFb/5kOqHgFYXYpxCFCNpH4PyvkqD3fO6/0O9H9
Ym1U9fazj+Uv43oAYBQT1zwrYYz5VFPGR83j/SaSK2mN5cbHiEyn/m1X+26M6/aRn1KmVshE5pZE
dNBbJeQW2qy1CZj7OzMc00ayKHs8ZAdeciUCWP5SHcPocv2GhlKO8P3/sxkhu19VG2LBBHPRUUPy
3c3GnCoudvjYMjZSYRcXOAkGBEYseZXmPhrjikbbss5pWD5ZMWkRMdHKfSCAQ+81UBDXS07Xzuyp
XuFuMxvUMOdTuLQGaHftCyG8fQExBVXT5mT5tbrOG4m9CUrAQbbpUBoMN5pUa9zN55/yeduYvY2b
6opFvsd4ajgiQt6czmkIVPVXsQ5xCjxAmpR2Aie4bAMfnZZAOydbLplb5TqzaMsPjrpfzTHkoVhY
J1ZYMcB79paZzPifQMREPDglU5BA6bW7OZMWrWzBeVpc/lgAEF3gQD0usOShYp/RgtjhCbDz9X1g
WYjffhNDlKj7vg/hBtsLGoecUgaRerhFdk1YomkP8W/MzCIoqB7G/FWrMK7AwVw9Xr3OoVD0zQiv
o8ii3sQ0HbsP2c7dzcYplBr29DeC8bMJF4Ep2nUZ72BYP3QjyJt7lUT+NffekaYwCLCONgc1FrE9
hd07qRzvojy1reDSFyTFrFXQAwQDhNrAeXotC1jq3NqhldwoRNMUZsUfIcZNzQasydkXMOD7K4n0
i87OHKQAf617WaLBkSzmxqBNR47FnngVcy2++8KT3apI/z/K2kj1MlfvrkzYJowWPRwQq/oajrdd
HG3xBhVmFZ3+8RZUGoA38nVXKWJzvyxEGXWVle3JPoXJIpzYnZr1e3WQCLidt/8V9CRjtzyMPYQS
54czYm4d277psLEjbMywJAzzR99P4Nk9Ha1SKWDAIJCoh1/kdqhlYcwZBbfrLJ/aHd7ZB9Dy4hgh
g3qo1UwFrwuLfhv6/StxpYFAUKG8ONV1mbx4NLrLB1sOFe39A3FSk1Msh0CQixrSG8GEIQ1e16wG
swbh14VlhrbcZJ2V62BMm6Ctv5vA+Z/bC8nlN5A6tTTohQ9Z8Mj+f5Z0K7xH8muA+pChOE1BrW6g
8HzkNGjaWcf+DumjpF2aYEnuticHEOx6i9CCXAwMUozI+gLW5SRqyUK80vbywdvzk6sHTY4u4kfp
c5IhRugSl6Ed46ZT2R8Wq90ghj4YC8YmILb3f0a4ct22MA8TJx3TCPdtxclyyvudR6ZaqdQ2FfT3
6vtPXyFHc3rWtwI1uNQnuoYqFrxdE5WeVZ9eKKBtyNuprm+IUrN1gGsfij6YeNT8EZUgKIef1v05
PaRSTXBeCE9zNJV9FzA34S92rk/JT8YCD8Bamr8nTWC/5Zn7Ydh/f0ATx95LC2tYCq+gvh5EBWMw
rAAE265TFoG0nN7vQhv0oIPNP4tcmP1PswqhW6tsrTj85UZERnWA1DmPBcOFAJMKsloHTGGno7Uv
OpuRyEVmRgpu9599+YnjjOg4juF0DdnAL1BUPT0THDNQiG8wDTodnGTR2/ej/Lid06UN6A/47M13
BRwybuc47A2ZqAVIIluNfe/6pGtz8oL8OHEZ9HXkQgDUZhrKgJNfz3z09V7vbqN9eGblyBFOdT7j
Tjiq7w6h2h5y62ck3bkVBWfn9Ye8mVb3rUk3upXLM2rcdDrrd6yrgz6XjH5mfQP/fC4uJRkyXKu5
rDKK2EwBQFOwtDJKTDLFNCr7W+Y2s9wwoEnrMraLpHLFd0hm4OxBgrasBeTOCBipkKJ6hd88dDGz
Y6/HaTWUEXeKoM+Meu4kuzjhsQ8BjHe+LhSUWUB4dMfacPHQZxmGhrM9tXD+WfZ+VuEa5VE7C6YL
1qZt+bP/n5hlM4mBLr8BWL3iJ7m3EWjBc/EmO1ZkHgPAfCqtiYl5bcVvlQFgvK/VhjIKVreMfeMm
XGchpnXcJyv2x+TAgKvkcmKXOXX6BbaD2PYqMwjLF440f5SkR7pERx5SWPdwnNnAij4/9/7+/btV
hR7/dtbB4yxpxgEkxMKVddGJ45+yX3aWwSKrmj+xPLDQeiKNYv+rugIz1mrQXD1OU70XpdY8X1iy
yT1fMp3+Pz+Eq0xO8eDluhrvX4rPR8mQxEs+yyCdUOXQa3roPwTjnPArIMZUPHBY5sI+0+3lUJ1Y
ylBE1QzHRMWFwVIy7G7E8t/37DZpZPYs1vJhFKZyPSBx7CdnVBFwwImnVqTcWk1Kh6yUy7zPfx23
ousvcSxW9fw9+p/aIglDstJ2H1XaZXmU7dW6pzajmB4N2MHHzma4cPc2cOmoPBKPk9XTZR162Th/
Hz100p9h+X38iJL0C0w5GJmsKTOBs/pO/cpexy3cx5Oyca4Ozg8PYCDBFQpua68luFS+I3cZvn5M
voR+V7hP5witlfQC4kwxUBPv480jRb9xLz3BL7MiYM5jTB9U4HTNQdQGK22OtJcDHdeaFR8DI7EP
Une9WC4JfGq2bvaLKwEIsBUf/x87A98pgJqGMndVbJ4Ko08e6mwVRLrB+v/McH+MKrD/2p8kkVcw
w4kEoMuFNoLCuPPC3zDqcCJap0VfPdI6fDor6e+nSQVSJYIIYSsQsGcsQ2OSgTbEh6JUrsSc1cmo
ZAdiMC06Ptz2cPwoTAULQl+hG56VcbDIpA/qu34ppweTH/W42Be3njn/NT2gejW+fu/pQVq/EwW2
degoyAz2vH81lnQnTtX1kY68jtuYmVJYLveKU5Bylgu5vS3XwcxsImQ6LjjTSiMLKzdRmllJx4K7
G0TmOS+0MbQREVwRbEuvWK3sthYlkYlwvRwR47zXA3b7F8AzDPKBGQt7wSep/tTGN6aZHNeB1n8g
q3+TQCIWEJIj/bFtIXjJJ4bLcvr9njywyr6GYmUm+ljcHvrISXvWwf+coCL8jW9SsozGda20LwHS
DVDrUjSE7gl9I60TaAhGjCwcrP7NrA6V4NWXhl5Jfm6EChYn3YP/nmgzwIU8LNyNAZnPG0wbsi2J
VbZod1BfSYh1pRqKKRbQWFmP2jivrWtPKW07wYMElqpgheUi8GgGfTIwBCrfSmKnSAJvLmTF04bV
X1Fxr73FnQctmrO2Po333QLJFJ0LOtoUS/R3Bpagawy9YiQ7Nk16yfPNP+MvT/MhQ6aN0jl4S7qc
T8hBCoxosj/jeuo+0VULszm8XXc5fi+MKaTxsKc6aB0vRFjsbZ5LcsPy6FOSfqRZRY1afC1/+gO0
mPvJ3GLc1UAGKJjd0NXRi1SYk6bnrybTbM7jGcoRbEnIoPYBxgijDVgchR4vO4Qmzg4Mvk+gytBE
DL9Ryy5akSjfr9g06qgIzN2z1ZJry3jk3yg5KLM3Ld0BugXPIBqQQNJlP+Q2j4BFVCvT5AIgqH4a
VkoxEH2dPymp+T3EP//1Ht7+ik4R5qRtoZzDLvdx30jCWEIpKE1hjbqvTHfP/gBJrHa0YrR7yDXM
LE2/uDvPy20QU1yObkFkK4HRVIWtoKHff5JCMQqFBKXKY4P04Wa5WWmWV5MXkMJ9W3uFcWEwSv46
zsrt/5Nfff3FxdV/pa5B8Da9S2mlcsAnIWBQMrgDwl/HXZEwX8NEdZAbS2Gb5Pt45uK6M9SuS+3i
Lftw2A4/ov/4IvLm42cMW+BdvVoixxom1M1Wf5ATgMZeowa7nnUrS62DfRH/jCFfgvBhxwtCg/6K
BUB0VS5OgL/UGaZ79T9qmqsP33oZZXxmEj2tcqTqDzPmL5RAnlBwuNB5W8r5mfiBcBCAuasrv/hK
hbxPiTXdkkeolbM5PTkDEjV1yPPEAJUdPeoWOSuiZjSWPDwGPJIJ9AoBw2Y5yvSYnhb1UQPUHACe
QblSJpgUGp5y3RHjdXrCFOh/4/gYDTvTMRIZX0YTYyii4wD4DFVpuDYfUREvMo2UUkjoZrdVuOSz
Dx3qYaz7RLFDSU6/9WmnWSxkklBoAu4W1AFY3IlyYBh4xOApLTYt1XXQ4jUhnWpY10F+L5RLk7Lf
vUxTkv8H+ZwwrQG7LmPVRRr+kZ1LnatpV6QNdBcAgIJb7qjcj8XBURByLSfBdaIo0ABUB99WXuoZ
Otzewf+wJTRdQChzRRXDPpKLT517T33fTM/kcp+wJooZdFGMjBOhTjlysWGakhUJSEj4DIAzyM2+
5ha7d23cdiOjGrzPB0M7rY5QAwMhsVehzZjjugzXrdsxBeEGY1Ei6ojeIUtaq9Oc6ih0cTNbm5wa
Pjw3/uMEmjuPlc8Wsi8h/qN54Ao/1nocpANYUZVZ6q97wGuu08n522UwDDiLAVP35pGRj9CRtevV
dxuuQ4oVV5ew6ZKeMOrp5QlNhQVjRmNXZdKtDGS68MrW9NA+XUVcyW5bH6NoLx6OAPYwPGyp0hS+
VimMTQ9n8ZvLaI+DjhR6kuR8+7+JwtjxOVk5cyODjwwZZ0Sc7uBX+0gyKq+EOYtTk55ohZNmSqED
huFeZa1LcC0yOo6J6uWrNwazB3t0GGPI94rx+Jdxd+XOudrQX7CfTTY1Wa1cnuqlX0SPlD4WTFbn
NVhvjD13ZIlgECel9n2EMNRoGfFcD0UWqi1GytYKktn/6XLgpXQWLQ1teqpuyDaWeCdZHbeOLmFr
J5jJmiqjBsgWrWuXIIUWevvK1bg2TJF+TYEw+Ot6GhN7yi4y2mX8WMiY3wrGkidT4MGGZROk3RXI
mhSX6yXf4crzxFtCrJcsRJJkjM8mtoC8OO5HiAdR2OI/GrVDXz4lLkJT1R76iDjkvD0qpZ+1US9h
6Vuh5L2ngGJ4M0MwpOOJ6WRpEiztaIVmHD6tNqBte2AbU91xxId2WHKud43U3Sv7J3tHVvnLFmD1
8t6vb5CgHkgrk2ZJN8RRu/7c1qKg5mGQNQ6COc+YoDQwe/X6mHiQr9Z1enr9XVSdIMZEnQJ44hZz
Ra9d+s6i5WG+ZlI96K7JFCr4Qn0qaBgRdUgfHgful6090Q6PfgwymcOgZvmlGId3AbyhaLotqTBK
sUwBOHMvgxuBA5lm1S0hahlBIiI+Gwnu8XIZHGfhEipskwjBD2LTwjCsXdjQmZp/khqc3jTAvEV1
8x3VDFxuLiPQMCsg48S9wSSqveZ6jeKf4KpX4FpUuVMN7JG0g0JFRm5ciTiy2zqzHgwPe0vzPrJx
2ry278fKdXKS6Ql+n+vWrYI1uUwLJadz5WohULJ5wRwPEE4sqC2pE/6QLHsDwfHD/Lv2Xfzh9e9Z
LrYqefxVkR6F4o0517aEWNj30BmAteMWLL9SaufQvHSesw5e88qmeOb/uE4KKU+Qh+krk7SGpf2G
1P3v40+ZMw739kCUGgsO334UK9j4JfxslSGSlIm3EHGJgz4kFn/gz9bVhpfJcKBK/abtydelnkJB
bSMETloEq6pu4fmo2PAzosHMx+NY7H7J6JFcJXdvK7bE7s2gZrKwtpLuOy6MOxm2Ply5sZBvxxSR
H1V+sOvPfWOId01H71GabZkBE4hKiIvpBa3ENGRp4KvYezVVMsrs2wZtJw7cH/6WA6+FPBa9URas
WYQtynigvh2cY5dpgD5bjPTQAQWES06AKf/ALtkuoy4gF1YnrtMkxgtQNKTrsSgcz+E1qANOk/Gu
9M+UsP5RnlcJGnCy5QUdxh7/Y0epRMLjEwBaWwaP4XNh0J04dWe5E4b5yiDQ+4D4eXcKifvmEKtl
VF2h/dw0OQxRK9qYUsiOArg3p9eLg6JxINdOUHAJrdvWx/DrYngsmpNlohYi5+ms5kB7wLHQTDgs
MBbq4buT35lcRwVpmFx3eagxCsrA7K8F9TUaRS4SB+wepjCwAgstl2cCTYFru08EnzCFlL/ZPtO+
cpb4kU1pytBpWYhRrygnkZnIB7w9QyD005oVKziNUG1+ioo7p6PD4HckwL3gndbXNq7VnbKDU4Ah
12tPM0ekBMycB/Fk+RUDVx8PupJghgu/luP9bGPoBukAx4bcwl4NxdldrDo2ftpU5WuT/umk/QE2
UdHfI6N3CIzS5KyxlfqRzpkL8Nwpf2iTM25/j8HHkDVTaQxAfiCVg1QRrvZrPYE2qvnmxT6s0Wgs
4JrzNqaFwoTaz6mehtVqNudAvH3uoP909f4BPYuEyg7w7FQQwQdESqcCpC8K5q1bAFtdXjBXdDNn
lV2injvcp+yddRqm20whJwFVJhs/6Z2zL7kgoPweStDgUMgjp0bCRZv547G/lITwgJQaHtPt5RNk
Fq/0j7oeThisn8VA8By3mtGwTil89tsWXkrUG0Cy0gGA5s9EMNLfyvnFqYUg/HdAFBg0mQKy4+Zw
9lyah84URA/nmz1wcsxRckyBJMoU7OsJLvq572vKfidZTJ3Jgopget8jzi10HuQNU9EZcaRWb2EO
mxHHxvknU230OJeXc2k0Lwoq2IW5Q2+I4m29KhGPf9P/5cSL11Y3CqrVeVjUSUxf0F+UsZ4BLnXp
R5lqLj6pAB5o4e5nWYOK4tjwD3k3SsV8RJ8kpPkMPYPf4dk+hzC3VmbZeIbccVbWnUlYRojoGzhQ
7EMFcqAFc1sNHhQ1E8OuIeD8cm7CBzFtK7aqaDK37L/GhFfmFSub8Ae81G4XLCja1qDt9gMLQF4f
n367ey9Qy+g0qO4YrFODQKlx287Pt10I/CJ9K4H0DVy4iOIKb7iFK+wWF106WpTjTN7AgZcE7aAD
X4rHhHNvtwdSPZfFgRI9IflMB8ky9Q7MTSNNgP3nBeMob1xMDmOcyQjRe+fPKe1bIadBbgehZF9J
SguXjaK5TJOqqJHgZr1TYI1CpmZgm7BRMJ4DGdfF7vBW3AfbHmGTEHqY+40OHQ5kcmqV2Unhj6wx
jsoKWZig32HZ+ndVxOY6oXKgbfHNETq3Yamt+fvEiV0ryp9w+ztmnHq3TeM8lIdrKw4K42SL/10z
I943tkDsPw0x8tOuUcitTjzjsR7Ugrz8TwqCyaSCgJOOjXCx9qMzaLH+WtUDbDYD8jeodzp9nCn4
9aQ+I7bX1Yj/tZJo84gxNUhErpLAF+VTxvV44QutaXeFKBb3op83xUcsWAdSI/ZWwGVsBNtw8CKT
8bqUdrM3BPNZ6CDstQ9HKfNEq2oAUR6z5uRBgRkzA78nHleqKQnQVo6zua8FtjqZYXAIRQDL8l28
ScoAY79trlbGVX3NmwD/Bwzzw5cUN8Ys1RjdkH09okorTjZ/BN3dIvWqe8G5ri2w1R45egQlDhka
Q2jYfeez1+kFYcMYOQAV3NeK2Sk8/E2aAGjtTPVPhkcVHsnp9YNm2cHsvGLd2LRW3g6ameSq7Ut5
8wLLVCp/wajptGUDkMolpHxmsWfuecHlUCRpeA9YZln6cftis7T0yi92rAe3//k8jv6IbPyRHlKC
jLU05K+FgDdFeqm8smQEyYyhJp1WoNkVZoJaXmdGRaKjrIeXrLKwAkGgp9qf+naHw60VV2qaGlv8
sgHZkUA8RDkXwxwAAH1KtXBpo5YtB5Tyb3Uq69Fsu4A/Y2Q+40ERMJJmgIJxZv0B84oVsWvECADw
2uFD1qSjjq7hqeEZSQC7i03SSHMhYVbnYTyul/x7sRi2N/NPF6jdSnrtjAuq0VPqHtqMoSEvoq37
Es48KQJfbNmANCE+mKWYQEPnGRRSHqUVVyxsxqcceAd7iRzLgMtqHRSGnTu+RrV8+FXHw4w8oqkF
UFYBwyHGsQuc7qT3sRxxmLL+AcDnH5k7Z6kNQqrGNVqvcqVyJGfSbYZE7O20o9OwU7eEphx/mYLM
AjvPavog5JaFutXvGOPMa4Ulsd8h3V9/8MJAvtIunuC6rZzLEyYr2SmXVQ3qD69dKt/mGC+Wik74
88ivRCCjO0ppgdeAzNbCKZFtmRNFqeWbkIIF02jS6HTMkYMz8zRevuTSrHhsy/Cf5BXF3sDAb4Y4
uhsWV86Sc8JjB1XNsnDemheUTFvRf2R/jRVe2QWIjzOBrHTWQkRHJLmy8irKIuXDolKdkBP1rnXB
6GQ0tpwKgfUJQPdvZrMPsEYoM1lMx6zukf+nimryuI1ONr0HliWXEmbjMhpgKfZMcwTxBOPipQTU
hBTcTbOMCt+US32A4UH3mgdPb1t58OdeCR7/nSo0eCmZkBQUvZUfTDvkF/zY/l/aLLjh22sLVxJZ
5TLiNa4q7lPKvqWhlhQ9Wr1iMWZWG5s/6BdMGuYFlb5JfXnZj7GNk8dUdvm3kuG3iVu10uT9Enkx
1St+q0ldML0S4/t9i9CChvurAPNLegz6q1mCABFqaEXu3eNbLHvI5oKWR/DKCHLI2P3HN2nP1mdE
n8D4a1V22acEhGBSr6ZCtmMxn2Q+EMop0FtZmHjr6mYoK7UE/fr6Mlvn/P2LnQofq+hLOA9elezX
sGhGGiDgVnRLNUdAIggBGzsqEC6SZy8wfYygifvEaILXZnI3Kk1Sv2NfoJVCB6zDCM1PQ+HHOSQ4
nuYxQiZkb5n23CA6tXqNUJWPOOVCTUJO6zDwAjVnG5QDiCfSperzypltOia+13s11+Q7QE6z+EMi
wzZ4twVn9lv24VNUgwQQM77nKCIHZ1S5OCdngs3k6yThP5LIasA2fVJRTdoRwJvFwWQdBw9UyfJa
sHKfvRdYG4NJRTQ5KVV9XyvRNU6dObwGlwLb8udDEVQxd2aQgcrSTnucEH2yWQT30XDJ7yvkyCfv
fytvDyiLCELr7ozirNKLDNGGiLkseDEkN37dyddnlI1oazpGtioTlL6Ensc0EOIOOhf8PkY2nn2E
uZ4qMDg98YVizSfHDYMnlgxBef1Tf02bvIzKQlUmmhD9jjlJwRV4E11My0rnVsSft6PE4KgrU/TD
JyXpBMaFkTaTTdWf7vLnCapCFgOhjUixeopT4rDs4ocoJDZnmiIiCkTQbNAT2G7ml3E08H0sny6C
l3DjYPLytIpULX9nE2XJkyjcBa4sKx4A6nG8Zxb9lTrql2qnbgO0t8Zkho7jMJTQd6vaVIbBVUFY
40TdNaUWEzoMqgfXKopubJtVz2ACJIQBcZ+l5ZNjNFFNy+/3haXBIt/mwD7ZeArquNw7XJ7bfz5P
sQUIi8ehJDqXI6NM49KzTdw+q5bK9Tye+ZPztFcf5Vj1OQ950izRSVdOdugQidBC6AajP57EYQ2t
QLHUnEEvjhwGWrB0csL4qP5WqBYEEPHiOKn0mma0h6z4z9UX3iTE67n5IKSE+hFMuU9PdmsT30LK
6VXh6a0A3oyW4O99vY5po+ZC0Ri7PvOBIy1klfq/40JSqM58M3ywYSur46Nulf7ivVo6GDKMYuUc
EcdbFrDo8JsMCsvY6pGx8NA/tmnkK6Kk/++LVJk0/p+5L0qbuEBUgf495kj1tBGJJt1+TAWJeRFG
iS2mct9ZVRzQHfGuur+qHSTaLixIhUMNdG7f5sQKqSu16ol9dVziY9K5DirqJsoBi0FjkWsVTcPZ
gtXsH1+hZ7Z5rth5a8McSK+P00LYFmhJnZ8ysddYd4QOBRfuqUfO5g55dXw9ghdmoxY2QQg2MeA0
YyAvw65Iuu6nldHpCoZR2gaNkv6PaIcbgFE49zEhpwnHr0ghgIJlupz6ns23DOwaBmTXyAw5SHir
AtKZfK7N4IEBjmtag+FnaqASddpq33nsvygPaKGi2dGrs/nwKcfU2074ABRMSjrTmX2lxUZPzA38
mn3epIPVpd2mz6yy4NU1v2ef8DqPfNVNdPl+GrBWCEhRvhXRL8xTAPPga8owScGGtE9af/15I/Cz
sjfC00zr56Aea1RzUQUi+cjUfCzY001sQFoUFHN5fo9mHoPeSM6zuVfIXTJR0KWgaLNywh8CivOt
BEJVQvm0Tm+8UMDw07q4qj4iiTUSguAuyS3Gn0ZytChwEzVCB09ePR1iNlhzkZl5NeUdQiAmcT/8
3QoRcd5+LIv6lq93776iV+iYaBG+AbodfXorNsLeirHplHSl9ibHTIBTaSdmEGcT3Te/aNc+9QA8
F8UAeO6NP991nQ2OOZaHVl2Gdq3x5BGdgJnrKv/NArrMnYEdznoiQiyCNj71mtvTXuPDCdm5CJUc
a9r9Ytj7igicI1FdN5n7vSkoa5++vUuvVsRTCsejX1UHTN/WmuDtNNoiRxdpvP7SBOMQ8uZri9Y/
rKtwJaquNZDlYRZHMCuzsBrGnkdwp4VnkVaiFik/lQ34VTblSjWRI9FDGF1GCmDyBJ4s4T9Qeufz
X4a6X8jmx1XOXSkPRdKkEhebF+C8326qJQhgnkpxyKygU2vlLNhvO3U/h7kjW7rE4GwclbEwRNSt
diDJaa0eADu98bXpnWu4X9N5WQuq3auYheoJ5Cw1zI2mwLN2zbqpRaxjgbat05lzDdHfT/+h2bYl
57wBAKuQEQ99KSrS6Nf4qqUu4+flNQdTAq1CkXVtWPQ5Wyre4vIZ1v+KCt2V3oQTkPaF/v6NIPlh
N4Mtf/uIOT+VoUYL+z1/WkqLr6DQoHVYhi1AO2AKq2jHsZgM/3ENd50v+Csh7x1pzYFNmV4G5HDR
yiktWjRLdtTUcyPl2plo+eJKaCNvn7kPehPZjJyCekG83BCdNUUhNSpJB9UZyQ6pRAPLUFiVZzsk
PuT60S4gisuEKoeLQ92QdMhpdwGPaVIgxF/iPLtuZJC4nHu01g9wpjI58/WoHV9La4W+rJ9ggrQu
faVOJO5ZE2BOU+fL6BbjVtALOp/wx8nGJxyyl8D8ITj0p8bEPOPvwT+gmXwk1sOFEGHzaxyvgSC3
2+lR51Tb+EGeHFtG768okQmVxt8IDuibqM7mUS7E8uylwCABZ64OxeZPSulkTGyDYfXJD90Ono66
sQ4YWxk0kRLR9euaauYHjg6OuFIkcsFgRGOPlIJHyMzDXc4XQaz5eoi370lA4YLP4tRC3LPaAzb2
q2atXTaSoRo5fHk9AQ+hqEUq3RhjSsNJM9NnGy9FaVdbgd7btvDaXo+Q6Sb/7TzAAh2TtZqLKCrE
u1NAWtjNP8yQZSvf54+gQr0NB7tiM0tYtWJBStAsDY4iKNRz6deCjBZOqlPmYUJpeBLzT9WtWHj6
Tt/crSWbN999R6tSPsh/lZgwvGrnDUGcTtbrNA/Agz+BKQH+fwWNKbuT6wldZVR6CQCwAZu7UPoX
foeyXUqmJjYqwS3FxPB1uMQmUzAdmeBYxy+xOFfnOfNE6QOQB6mBfmXjXlz3DQrFJomW/Oc+Cr/d
BLcTg0c4zPg975kiUdYaiaw0H/tPiXsHalSomWPfsQsUPv5Q66F99omORoTgK79JNh56H8cw3867
r6sHkVxi/xtsjUECix91gD5MxOiPWkg42o06PP9Ve5UEOyBkZ6sR9tQBYak20EzvHIaBBRHA+oqS
e0RGPc2S3aT1PogXNNKeKPOhaLez1x9OprmiFLaBdpU27wr9/3RXQpA1MXfr4Ik3nhph3gjJs9aL
klAm2KisxONJ0i5xMQ7+7AKEx1xJ+WvNaO9w2rDzev2lgdMyMB+KcnvxtissjK/RpnyKitV8FEg/
64ayzOAQBWocjZ1uTQac4C6ny0wIb/42cNFyR9e2bY9CQwnSwWHEWnmtH0YyQ3CCUkIfFeq9Y38y
AhNCc0JRz8DQxXANNoKwsFLjquGwFuMxbvoe/LGIvjZ6wykj/04mlfAwOJNwfcKdmPudV+76WjVt
5h1yxbhT+lGIfCrrlPlA17nzQ8HCx4SnIV7eKlWD13U2Dh4UpZKjiQDriNuPL4coKItG15irqaxy
lnVD7I3AAhPDd1HPLYMnFstrGPedJjD+GKdNuu82BIkQLJccIqCzRkqRLWSs3YivLxBYmf0ayKpJ
cqQln1Ph+Y78RDtuNIjzF3vEImu5F0UxN3mGgMvACkTvi+gez0b4xumsb5t9U7VpWYbniXOsDuX6
c3nXI83OfWpwNg8Os3ZiECtoBEU6hq0M1N+k8HFHBJE2WljPGJSgkgfqjbXdcwQRd9o+g5RnZRg2
OqENGVR/JUD3+bT8Y4WCEBEWEMhLswncZa6mauSqgubnrQ4zMO/qPU7rZYbTfAv5Elmt56aFOP4n
Afad669o1jsi+sotFF7qTJUzjyt+BPbIno/Ou95hgSmAdgplFVWOq1JiLTdlby8HpcQNEoUIk24P
vCDtCBtB5Hm7bYkLEkTeWzmfnyUUEWm3Jvj0YwSRj0HGg1AoG9PAqIEx4wFe4dUHhdlQCTNKLJTJ
Ho+bDNW8DPtR+FQvDE6IMGdgEYcNG1pObt5tnIB9eRCIgGsR+UdxSr8RoL2LB0SqSXLzYMGAUTU/
PF6P6o9t4+keyTZlq2FlM6xtMu5yz+B6jpDqxHJe61hrSftehC2p/3GeCGJJ3vHZxssT+CrZTcTl
mwvqyJG1t5qZxT0FoW5lSlTJQZqIRTMwXNDjpZk99sITGNGeM/iLKEXc0bNnxTtXzvCkaQWVWLMK
M+qCaM7yXC2PoYX7Q0AvjQ7pWWkELcf20pPfYdvKpO9bkiTvxI1fiR35zY5SGija1dpEmhDB8OrB
S/GwDqPDd0gIp8VwbUgxcMQOIVtgRQsA6qDEXYkHzjaoj3r5vg2MuN4OHqZhTnjWTalK8LC5ii/y
dYOUpQqcDVwRy1Zdt9+VENdH/9JbZ2d7h5QcWFJcC72yoAuxG6keQ1X15qMau5rocvQwk6t5LDiF
Lgqx4at7Q9F35YZoXXIFb6LAjNyylBMaZe3JdF7PBaHNOQlZUiKbNi0w9tNFBQ4WaA1Z42mS7vyR
gjXMUJEMANZGcY3n/96EytViA+1Rb3Qw7LgE00jpWU7rxTD5Oi2w5INfUXXmdw7hSZDC6/owcfBc
U3AHuuSvsHA8t/JL6P/bbi+jo1h+oj8ec3ksOLAdWW6KG0BW8V5QHN07hccYy1hSwHp5Mttg5GF5
bsn2vuPjZmd1vu0U0JzXGg003QYhInrZpdP+Klaw33YToREQcgq8ESnumyHIwr4SDZHJ7+Spue1B
oDBT8/Yo6nmH/kmrVdcyRxIVVupA539AOBzQ/zUfh82VPfu5jB2MPIie2Ox9LiLUfWa7gUDA5eRm
nX6g6mzt+yANN3YRxYgdWBx2p4QvIobWyMjSazqUhlqQ19yJcpNlwK6NrRXk84gsiXe/TDLCJrdH
KAapEjzZ9kLp0KX7lRHuf/s6s4PeSpujc5/hIQDt3dYIeRxZmaLW57zqxlmc9R9Pe+vNCEGEtB3N
KWbKnucOX7H5vwzq5hO0pfIb5lR0Q/pxj3qa5pbMLDM+X9tK87g6tszbrAPmIqUfd/G+zkYHIsZV
di86vfv+thuEMXWXhmPjaiOQbgsGwm9QtZ4NKVIpT07UBydZxBCh9nr/r/rGBzyc5BjyHY28GyUo
bKj9SrOojF+NnguMaLS0AwmtuYjKo5kttVvUqV6SUxV1fA+MS+g5LkG/HnTOfaV3DJxcybKZLrUy
y5yNGn75ocCl6pucpavtpRDpcPvXPUyjCXiAjKPWl5wkn5UH20kuj3/R/hSPoNVykMV7T51tGGuc
FasJ5mU/FCiuuh8lnMLsz4eDGwFYq+7YctVWgxDEpc8sdbuwvb8ZS25kUeiF/KM68GoCcOuUMGxM
BkXFXZEPL3/1lEKB+4zEfxvn0sqo1omK8BQO9pSPmsJ08ABznlUxe+kEM8roQwXGy/gthrLszs6+
j3KXR6Fbj6ZrCw+GwkWdrpCSXfyunPZi1lWeMonN5QR4Xa0X1D09If+XrMxJIOh5SJEqDkihZ7Ux
mQmBvKofaynQ4JX+cxD2yxmvS0WCe3U2cZBvj/4gyUsp/bCt7asC3XdZSZVjKjJfc7w+nXxgDePP
MQfPWk1qolf9PtPRJHblKT1g759Jc2mVBA0k1cukTbyYkKCmDZeiEIcJanKgNxP/k8D/TjFfAx1Q
yHlqzFxxrEJo+cDcB9uHZ3I/J5WCi5T4HWhorRZB7OqAA9Qook0ZvguhIbfzN+5huiT9sGtOY30/
hVgi9q0ohBSa5OYSUsaTPwm/+10CnmT23Cf9TDgf84XYOFpMQt0QxFs8V8eFO1cTdOFDbBvdSN/q
iuKk1J17n32VULdHo1SaIKujaprRM0793IgRz7VFzGw/8HzFnmQmC6LsIcdJVr9Zd9Scv3MQunzV
3yQ0QR03rSgKOixWqGjrURkedRys51U/PnRCGqVyMJlUkOyrw7j4gXFvXLzGtRoAP8Kl7I0Ji0uk
HYqFQdKVBayFcOLE04uQbDuNBPWNGBwbQIjbfGcEltvks+KS+qLVaufDRlYxYy9JL8zufWnQgl5a
foK0yXErtqtKacOVWkYdImIEFd0licAkzAl4XNVZd8raYQ6TXACXe9C1KZwiThWf7qSKqC0mw9UX
71unwL4rgkq5Cgv1yzMTNxDwD+6ZfWrPRPak/JFrg3gaZdzpgd2Qx8gooQALJmEA0Waj9Hajpn18
7cM95F1aIUyA/vVDkqCStZdzw0U/8zMFHkCXohbXwveOUMxX4MDWtkwVvknXcGS2mk0mQKfmTVTv
wB8hFK9O6ksAhHfu4Tyark8VzEziHzBmBfWOaH5bpXp1GbW9wUqX7f1UL1VF71boGbxwaI8ybH3K
NKI30KhpP3Z+ptyeKB1fbkrSiDPRqvSJPmokKnoD4DDTDy6X6fS87G4NfpVcqjtYIBCRQFAjxilr
xsk1jB06w8rzE5Lje66MPzuaXl48n1AmslXsbhEolPPmlAAoF7nVy1Q3Vr/bysSP4FPeeRJs9vh6
BfkCWZlBHj5tpQ31y5Yp6VtPt3pDygh0D2NZDz+266Y/2wMch8qz1mrsiduXH1Vv2DNzwtk4v6iz
AXhobHe14aJE4ywEuSBrrRGi9pgJZNxT1vcVmayOVWfnR9jaRUbe4iFKFun6o+0zoLqKR4zLuT05
DLd6mLP+yAejUCk3wA6+D85CQTZ0rAvsdGY1k+QConz5vOUq0EiBxdRPfR3JudXVMnGUW1KJ8azv
Y5L23OqbMXbQZk8JBiNnqsZLzAxq9BbQx324gCNWH6u0nNTGJ7lMYKHRMzoBr+ddf2w2wgl4mK7c
0epaQRUn9GMF96VqVHob1r7yf0zpv+XyVMYnBOkF9/w5qSbLYsWjQkLn7zPoyj1JryORnhZHUpXj
UYCKue+pYganM98oGetwxc9yLZONbRDe2DHvcQ7wXSlUb4XhnZuFEz8tXdjriKq1W80sxuvwbYXC
gJWPiyBICaLiIDOvCtKkHYHyeqKE/Y+yC0yLURnK4WdFpw/Lfp6pG7TcFE3zRbgqX5D4ku4QtFjd
o2j7gGuLG1WxYTEhY/BJpXsEYadmy1r/8FnGUPD5goJ/MPBREI0jdvEq/O2a0A4/dQbyAGy5udzN
BDrfbNYgYV2QmyFCGJWOZo2JiKPwPuw/3w89uUVJf8YyeF2E/m1BiYVEpXjiPF27sEK3I0x1q872
FfqeUt3bb4WmwUGwofNxiCU/v6gKlybujT8NP9lMh2m4GHlGFud/xs3NIefkHdi0AkWsAuDZvp89
c4rXuKtXBdGqFnKgZcv1Z2NYWpSCCWa4tt0liN4KWHHUuMDqiZqp2i0DCQBohzb8UTkaAea1FuND
2Pvsu7EAMoNme2oD12e/2b7MFLwD6K2jiEUG2GRxFZSTqqn1yOfy18g9FNoa2GdlpkyGQCLv54ZK
sU0r4OqFaaOT8qVJNvtkf02mz7Eg/7Z0V41eUBTFWni5Q+Go9Z5Rs2IPGB9TQw2ZoJU4hKDYY2Zp
+lUECwLjKe6zAa0feKKJd1yKQ9XlOv28D5Vm0XEdC5UdNYShrC4WmmiiocuWrI+75vhKET65yDrQ
QjmMlCytpE7JOxQOKWKQZOh3zNWPhh4akzi8Xrg17O5zJfNh468jxT1lms/piFQHTKMoA6OypQm8
6S/jU08VLQK0UlgX860qOXcbBRUof5KoEEREEgMWTp0Ho8GVk3TaRffA0KUBtdr8LpFzHWS0TtQm
cM6ue8kmD1h/I/rXBYoOvwaz3oFBPybc+IIoFD3iWPCJy85bthmWbQALj61Tj0nULz9QFsOoJpGT
rppSoEY0O0Z/wCGl78eGkzkkHYUB+zMki2FCg9nkL8SMndBjd9Tdawkkb5irl4Tr0ptszI1dKXkA
T7angSo71nq+vYnlnrPyk77Qbc4wFdiWyvGuG31p993el3Y1SG58iV+cGvVxvdl1F53Q5DC7pR2/
0c59HUTq1ScGeztWLsn6m3fsHqvs4k0NtIgcIbknfb28iPEgpQuhwo1B0LeyE/MiJF4vjXmt4CUe
z3PlEzefjcO3Q+Blp0qK1PnX1nlaxGwbg0R3AIkLl7DfcrL8ByFbT/vDO0AkMl+l8K/VT/m9cCdS
oFOcmj93g4R8XIVH2h8kdtchQjBxUynwZx3amtGwBDHac3hlDBhcinOeGZ8UyUFHkl2vvx1yfHwS
TuKTMkxWZiIRTLFnCqyXzWzE3JXlkI38icShXMYAYRzYRbaeJRHZcVcLb4t13x02PWyiUZFP/zxg
pstSzd2WiVwy/ZWJCs4A8MKFT/MUuWZ82AJkRu8jOyqnYJV4x5MebNwg+pTj9EREqkMufEvC/h96
bOumduV9yNXQRhazaB9hTcg5BnRc8MwiNpnYTH10zgdrnB1pXPTEkILpDz5KUV5ONmKUlX+Hjvr9
Y5uOAPSy8qXidwb4D1tJ09lAAKIDGSmS8QVMo4GaydDSGOKCgyE39FUOkkvaofHp0YYZcxNCW2j1
Dn/z8mkZP+5hW7KFCmYdu3h3cjYo5PmYbByjb7GaVEaX5PrnX3JkQGQSUvS6QFBw7Em52M2px0VM
OGwRVXJEZdAFvH8zz28nnDsfj5kgpb/hD/ZAYpXw0/b5aITv5WLwSH1KV2hAvTpUiepqtR8etxx3
CMqSieKdPPD7f3nl6EI6u4CGOh7c+l3JmHxMs+kWMutCu3VvgyzEl4RZt4OpfMPeB4MuCHzz02Ah
K4gVA0tVQ3cUYW3njL+FmTHDJ7nFPH/IXD7gxBtimeqX4iLkeeKwWKl86GKXwIwwAQa4/CB67GgD
GWHAWuv2OkAZCTmUcegTkrWL3STa+5+ZLVExtxk/AHZf2REhoJZKBu0mz5xvU2M42PRP4xAk+1i4
t2KVWZc7I5lA1N+7BgGc2ljLu9+KM3f56cIkVwXX4eH86im4zoUoDEhcXSBf0VYv3H9URA7emMWC
TeOd1HxHZ/prHjL2tG8F6DwokHl45I1vWEc2N+clbmzwYnfbumFnP/SslKkFNSPx6r+FdfMMSVEk
6cIMVN+U5Bu5Wil9asJBuYLG76GAHR+XhAQ1G78erDUiUFdn6rHocJWQ3f9Ts0+19nHmLnEfxX5J
iMLH+Jw+rW1EBHMu/nYpI1vZqHRvjm9dLQ+b+WxMCJVemPQxBWiTShCp9FVgKPF5eFwXC5O1hu97
j+9NpCWS1Ox401BQYrWej6zQwTVCBazGzd0hAFQBUc7uKMKHwWzNAOL75rqpyR8SZMznhzv5K1Mu
yRvFF0CmwgJhlqRgnnZRKt4gB94+ZHviCvxuCfCeA1eVnJ4pMhQY6t+lV2G0eVQX5ve5u4uibFO7
W9qMC8FuqPqT8pcGWFrINTmuQ/aCt2Yv9RJ7bjlmgs81rh1saR3ndUIibgT9o2cAZI0UM13vGZXT
0g7ulzIHb+ovXaf3i6p7l+ZivfK22Db1acukQBYl6LFEN+gEDVJNsE1WF7Ptix5ekVsKtDAMRJOA
G4xw+aYo0cMbvQPiXP5yQyMB3ng+OqD7Jm132F9HMbmO3uRu1JqGP0UWq8UcDuHuO1KeNfMuAd0t
EdtqrWpJNLTt8DTmegg4wVZSXsAHMfsGsHWfCJbfSV1iUdzpU/OkGIrdRHqNWI5eQcniwfYTPRhS
zUtDvS1cWlXwlXM8gHHBrV8EmMBTadc5H++mFB8yX+nU+d6xphLDBTsIyE72E4OSFcq7AKZillOb
c0Jn0TnSPQ1112Egk70QL/VPjbGT6Xk7XDvIH8dXvpg5l/tt55SIbnF5KW/kb0I8LZtRjcrp2g7S
RPy7vjr+6jwLlsNweCe7BOVfy8dcgATTcHs52KXUmO+9AOWWKb0kWs2LJbyQzARsHj9j8I6rzBR5
VLzN5EuMxGkWPbRaE+nuS7VRFGFQuoznYqRG7NMLLUf0vuB8123Pj5AchpeKAdrmoRbwJXSP3SIi
wEhXL3tENFLlm4QWuh60vQw737tqFqFjeaXJHRhsgHIZCnTMTESh46vGQOaXHGwNNNpRzFP417AQ
hmWdKRJG1Ez7rzBq99BuWMvrUbKdmtEXjAXFofI7LXH7xS/IIOGVaBS61qh+TYCk+yFax+j6rFDX
DJ7JJA0AyLHZUnuarOogwC3lJXDvxxWj8w72mW4cKnpvIyVFkFcyywEID+MeY7c1M19SOZW+UHPd
qLzmPZref4wVB3akFnNGFAZuCnwF10OV0GqBG4rCwUH3jroGG5fBkPgnx8ndDGineSrNyJ1T+4Rh
/iOf6YTP36sI7S3uRp3L0XbwTzDtCm0RuhOeomFBdMXKcubJlSZDDdAY/rbsRcTmReufIhxTox/a
YP+R1f5tKmlNjNq4f6RrtGSGSweo8sX8pQ8ePQqk3WT34QR8l9TTMZj9JzIMV9uFqxlZ0jqaCdVd
WjtPiuqgfONXe7l/qDfiJZHuWZbvP/9xdl+IvoojX5GxBcrhbTA0fn2S/QiLKaHOT9DiYd/uRD0v
n13xg45upJNzcfe6w0XGaUTsTK18rUvRG93XZX5EY3dBF3f0Mw2fzyQm4h89SRbKYgGsVb92ww58
FuPR7BLlC4qTeQ+bNME5eGTF5BceUcQpsOa2/H32zFzPVvcLnJALWb9EMCh72T4Ip4cal/pfuFOa
62oEYtw8vhbsKnu1bQF96jpoBYum/9OaJIlOLuYyput2imMmy8L7N/XtYHXJ8jGk/oqlGLi8cFUW
ABoHd9gaUktPZsbcyum3pmg97WrmjwsNc+eTT+EeS1SagOMqzDwJ6EFfuO+3B0dAHMMls8PF/c/W
LmDGL+Mlx6huJb2nLYihqld045bJgOPirArtrrPqPv0pEzFzcIwtkyz+0fCEAyxz9du2cULmFkZ0
OJd1FaKfQvd+SCzgCLeUcAF3LwesDhde/BGFvILBpEL3e3P+rD4OkITNRo8lri2qechTjtDfnjot
/5aUkN6TwmCnLIcXS15YY4xDVtBjogxIWNWmajNbjPg5pbtE+MsK/xbE4jBZet2JTRbFbZGyd8Fj
HA92iQB8FgQQGMplmk1EWnBQhB5SaXXPPzUSDc86n55osjHDBMYP7R2QIBjBUuPaSPMr+qMuUEHs
XswrEfBVR0maSXMsVht6pifBZkMtNx6nTWlpWiqordM9A5BPPJgXJ3QhcwEBi9498WAnnBdz7BzG
xqVF16tsJ71VvUorAhY35poAd/2d8LSizlm5vQdlLn7BrnkKbhKDWSeVjXtAjh0nnE8iGvfxabPS
YH5NlxK7NdXRavGUM1s/ulSSdpGTSmx7CXdy9SEp9jUTP5gslDMLCvmr/V2LH3THSj5f6BLasM4z
O1xqq6jQNtKBirFMACI9X0+bG5UEAUJAqPVZwE+YmdrEXf25RMEYvpT1EUEY7d2BKQbligp+tYL9
vjleBJF0jyTbH88gXGOiLjd7KceqUpJ+ua8fKPDA2by8++ErI3COtECdhGmeoB2lVB8XkhS4uBy0
K7GOKaM1AUgWUDGAHR5dEkDWgZqBLKLjZ54DKN1taaAQcOr2lcCt2jDvzN7LGK/2AxiPX2rSckGv
BUAXkbKkwT6uupym9lXqTGUERzaW+Avd9jA9JCSMd8TeIhZcLkeklYVWqD0HNMDbUZnzo0kkjPjy
wZq0hFEqsZjRXzl8wUIx0OTuyVHqCTlRmFWAlW68wZoVSTIR9fp1r2dGGMnpwRZHPWLISrglPdtH
/9VHq0hBF7M+2/DbokS3ebmAQn8ZDsnZALUlyQkIcRfhqY5oTZ/DMLHRnAp7X/4BRZLuEumNumhF
XjSn6nwwBABDNgzcu9lZVZ3KsmbsjwyFqhBWYtyndMopFh4UgwsfQXhHcNRPQZh3VG+Eajs+5/Lr
Fxb5gNW8cDqE2nFGF40nvnY/4mW82mekGLcZ3qhPEyU9oVXCShBk4Ti3GBraRAte3t0gOKj95Kzf
Gg5mmn55LEBvwtjE2LD9Xopfwpj1Hw6nDfy2LohT8pc7MR8zsrXqFkz51teqUuOgbwTS7DqeUpnd
d63oQ+BVb57AmnljuewArbK+DQCFeIx1jMCDQiFS4Wj/DiMQUnmCVcxKPLnAdnBRcHcdb5+WSunf
sGBy79dJSCeYgXBL+2EsZXNXaAVwnAtqxOuqFhVNMV+wVQW3P1chbNkd6GB8tB++de3BwvH8HcwM
ryAXdYOy3/sAWV43PIN7lpTecsYZponx4jPaT9c+zE0b0aVrPrI+F96RA/WkLEdKhuSLwyNkI4HH
TxihY7VOugwe1v2LEe5+S28PMu6Qz5kGjB4QEfsLzLlMA2TN/L3FkQje3mwZovaBnqpYNCLL6orI
atH/KrtnluEnSi0F+TW4yHwAJuNol3TnY+0RguCK6dUqBpFlLB9d5x/azHsIwxKFT8n/kpMV1war
r4OFZq15fNIWxdCRpI28oxorcs9B3XczSwrhMN7r1R5k9QRdVR9YvvJ/sY8XR43B3YXAxbbi1MUw
TAevIS0N0myFVLYX1bRacSafWamPykHn+OGOtSNbwzQlu3LRMtGebtHTqjJkYozvn1TecadUgKIn
XK1IcO8VGlfbmmHKgyqDkyCM/ZbcCdHgvHKDiZo/h45AMtLAxamNWytTibWUSS33wDhRBsSdPJbR
NdQj66TnQ1rMQftjcI07DIUoN7eCUQ9SGe7zGPG4+3/SVqSweOHFWG+r89c4FZDHJWJAfkaW/IsW
isQJ/O007OSvHvFvBx8KATf7oD/0VY3rtpZzxYBResx/QdvWKUFLBuWmN7pkerFASVFZ3NHY5F9H
jzLzuf047QH6NeK5yp0bnX+QgiVLbNnPq2IJV1vPYqRiFeXY5cHa2yBmqmw+ba9B378J6XBkHXX0
Dnc4wv0W+17QD4gddLAf4GZ9wKX8+jdMFPHO1qqZ2KJSPAIbu5GN6Vv08qRj4twPhFpOL7M894l/
z9fmil9MQAKOy+dtCiKy6iY/n4LRVH9IYcjDBv4EDqDFQhDykNk+wgtZ4FDF+Mof3E9N07SvhC4t
wENtw97sTn9JdcRUW6Ho4j1+dk7FNTn6mOLtkJ0LFmRyLs+fqGCVBDJ0mdRPnGVX1Mz5LSv0kuS9
zNUeiQ2jATP6N8eOTp3Ik7Di03OEeIN90Qx6fPlV2FiSI9X/hAtZ8041db9gVr1pBxVqoKufoBkk
nNiUBHIO5Mih9hKZVY8RDrHrmgxIMvjmebEEuIMEaAh7WpTDb6liUgkYljNKyMR8j0uHsrRlGvPA
v8KkCF7TIxmv9STpoCylJpJrG5Y4OcMQZ0F07L5yiOUI/Xvz75iEGi7+DYBlrrRahkMqFNduurHw
XFCID8/rMWsH6Vd2W9IkC8iiqwguurVnN9ucxUF8G02s0CV1ayrnyhXxRp8Yl+nYzLC9vrCnthw7
X9QQwqt2SnmUL/WT5EeJ23MZf0q2Rz9b1lbcYpGhjOKLtOBumPbQZb9hFImqtx+0cdQeNPZrVBWd
uE7OqTMSGGJgOFty8AKpJjhVKjbFpkuHjUyghTYRIouW5JIMQjHrNV0btUSYAw8sJ8RwTezhbYgU
tKOmgJW7fFZgpqoE5ACauVg3Ia/MQDWPjaKzgtCblOPxi0Pz2p7ZBljaTH6hU8OleFN7d/4+WX9F
/8eZSo9nkuBOQUe0iUm5lLVX93sKqqDHzQEBNGE6ywF+JkYhvleEyEt7Mt1bV3Bkq4Cx8+aTc936
0ENWUq7XFjOSkb43wNWjh7mN/Z+AdZ9ORPOTOMFiqPMArVNJcRXcKbF3VnV8HLJwPKsyx3tN8zRE
D8KUdEhSip5KgTPQATNrICPqjCz4MOjNZLGmqjRUBZo2E0K5GeHYMbrp+RXAslgs0DynMh7HchI8
QBHNVByKXoK1kLEjFWRk1JhNhY18OvEopAf0mz90M8/vVSRhpMZ44a/DfQaJ4SF7cvvarloWz5N0
Sj5tnJKFPS8usnbNzVoyPizdoWk0ZLVEiuQSE/Y/fSym3+EiodF7bl5kYWTVXy0wVLVTuWUxIQKm
AozE1UgFcjtf1xkMf1jDMIdvktQekIitEv1XWXlelLRj1D7szaCIv6FYXdHaRj/7Tw3YDdwCmHAP
/uXoVmuBbbd0DN1tKD5q1K5YmBvhunICADsL+tMtq9mjdc9vXXpnWTzQesvWTyhTqDi3lC10xjVe
2erxy5/J6IPyQcRwy01QOvBGntv0pTwTn5KlASRUdW7OvUOrsqkUpnEtga/nqVAiufVJa6BV/MlF
x+6u96t3OLqTYFfHNsE4ZllngGb9EFmKF8UnujT8cU87TYYh9wwki4zJjjS9rfz7YyCGVIm8LgsE
9+r+MIokLuD5QSQ/Mcuo3qWHiQxJa7bo6fB/djntynJc1RPls9vvYGm2JmD0J47Yroeo2lJXSvJZ
c9mD6CNJS7kPc9aO4AcoTKZMJSf05bYhTN19/5eLTajr7/p77Nf3Owg0JBzXPuXZOYyAK6Lvkwi6
5/eZFDypBCKpl3jpoQ1Djz2sKZyT4wbXCxjtofv2ZgVMyoFVw0U1lcLedSCJePYJxPBJS+xWXpky
k/EY2DDBkBxvPM65hoPZSQxEsYPDpDdIRcor0l//DPksoahKHiITPhX3KxFkHb+nUM0YWoTrQiWn
VLrPz3tt6VE56ntgbq6f1eloW8tWIvqkJqf3hLmSA9M3PbVk7lIv3ktXqPyos71QVePOvqY70N4p
QN53CLXHcBHLc+0xL3vQTTH5tXyfhXhfjkxnTl67iVWwz3P89iVYuZqf5G7E1ZJpBFNHaXn/7xn9
6DzEn1HdEArRfa5/GFD/3IVn57MFIgu7k+cS1U2pEJvVL3rxkqH9epaquakpfvclWiMdkFgHoAgS
je4zoePNGWrdeDy8jz/aFA06BQMGLhZeDAkVdNNPnGDx2wl1nSvSJutvDsnAM4acfRPIXr3yF+im
fiYHmkS8hRviaQSph7cExvjNzMHR6DQapbJ7E9gVH7tpLR2HqfYUo57U0tdokm48si25H5qwNvxT
mvHKBf7WbcSKz+bQFT27Xa09oxv6xsiA4lpA2PdmPBvbIEIv2co+eoqlKkIT/n5RzYojmshuPww9
LpRh91eKmgofNBm0UhX+VPu20tBsgrRowOe8BuJ/c3szhnepcqwl7FJ+fgTgPELsODSM95IUicKs
YhF9jAqsEasBxhtiDnVkEihiYw9PZad23APGaU27DUkxYSOAJwriI0iXQYpx5zNf0Z8FR9sNquVf
vu8b4ndy4/gzCHq6jXJFN8Fdbc/dI1k7999LUS+I0CNqHMNYslqhZnTy1rPLqT5gXnHG7nj9zw1Z
HPYediu3eTzlIwE7/DYcEz/OxKirqG+LfZPvO4bGL0+Y6w7y2TantxCpSb9EKgMcCeJtBjBd0AAj
bVLY277l2Ts2/poYCl/q3O7Bk66PqINQ09Fc6vGGabPKZ8TWREGhiaRPlknb7SkmUefzdtG7vJ7f
Mi5mHsw/yQCZBDvJPfV5qFc+ieTbLDbVhGV3ZUfDk2AQiCbQIfI0DOuyUJD+7TEetdvESagFDzRD
4s3rMnB8BysFCXTQBGOFRjHwT2QSVJdLs//yq621+cUZ16oKGniWjEuok/Qw3E3YtZ3Y4xAPLexN
5ZdRS1QIbN2xkVvqJHs+xsR8tH+gdgdYGqg1so7/CM4jYjp0FVU8Cqpo4NjKmAYAzfl9QbbTvwBJ
26HtDYa6HyKjG11F7CFLXZCOif1S0CnSG8rb4g63xdrRPi3mJTgM8RuuxOw+P2PXo2JSPe4fvHdE
XT657j/OqRGvwa8ej2jchV2+hD4bVXZG+p8a8Vjytjh8nThBkeW1AvGd2vAsH3IFgxxFbODZaZYA
5I2xcayV7oOj6uRZa/HJ6+1qNCJ2n5lWwNMII4VwR5LsjGKpIV4RNk8jyVnQ8YHdIYsOkMp7B4hP
OLpmgiG57ba9vsokpyV+k0Uaf1hPRimVZywtTtUpDZLHmjRROBBB7gwF+yhAPwTihEJHXxy1kk8t
XFRI7gTJWVaTngSXgnUiNCpDEM5j3JtqgeUGnjQJd977xdKpG62iWkG9Fncajmx2TaGz1ZjFgCV2
xcaYC7tYVNq5cjzbe6BTWibVW6spoGdugumF4ZyDMlt9rtymVU3Aorjkm4tB0m4J3lZs8UGFAEsW
tQ3TldousF4hzZ4Lr8Voeu0+r2+SpVJSHmCI8zf+5IhcHVmJqylrEoBAQ1GGLnWZCEEJ428PgZre
qDZ0VQYfm7ijBZ8w4LM3e6PhQ8VYCwaR/ATM9YI3+hcHmQcAPBXXP99J4rYWgPZ4AoXOZq66mhn/
QPMzvN9KiRo9gdDaRAaQqw2F6sDGVUeZBBQizEKCoScft7+8fuZQFJHDHn+FgKxVktCqE7lSo/jn
v3Cy4DR9M5alhxkMCxtQerxXJ/epEgD9svjH+AxVZ9WfueVPOOD5uXcpA1y5DDN45dg2FcOhu1jM
EuGu4Ri41TW1PEOMVRCjEwo8rsWkn1qwKBydpnlnvmIifzxtJVYUY0OSvepsVyRbqU/bz4Au+4ho
Y1UocQR8A6HQFR1YU4R03ptTJos+BuD6JYEe6iGis91REJ58L5rRA5HuW9EVcYOhMxVGmNfibCKN
LMmnGLgt1/okt5yMwFnk51o8TcfgBubrlF97xMUemFpUQPr2maGXr++scnZAc3SgzJUGGo2tyFYI
r8WEY3IUK3IWBC9xrMgHGmqrnTmlt98pGz+a6Z4JGWafor/gtGJWJx4hCI7KrM9Vjw6pzV4hGsvL
TFsaugCTXsbXr67qyHFzGfS3o0EmYDsH1pyaHCU6KYCPqMnh2WFWhJgrSP70J8RcdbYLPzyHbv8t
EFcyc+Rp8qqgq+LcZRgoGs8e9PrDt0vBl7S7d1RAy2mC/zHohBZkJebBNWXGTG1UfrFT7UH6lEgu
ciGP8zmPI7TX0Ey496q3+fbMFFW+T13FhMtW7joLD/CLkmGROe3QWRWCW+J2cgraCCPr+QJzQ1xD
jKra/1+YNWQpdOcnx1FXsMU/T69DRsEr9jLkF3CqAXAYVfV0y7RTa21yhBHAmdvAfPGZ4ef4ohlL
vn2edBkX2eXBbffAHyb2zkZ9y/hC4e2pUsWmZ32+w4N3QoqlJ10XeXUYzebM+RTzh2xePsegPLJa
VTTMuqp4SIXQofOB9G4JMHu18iLwSwydlfz06khjk4aPGyUlkmEv1LqOnXDT0PzyeEha100fs5At
KQKWR2ITRr8wRebREbZmvXsC6QJse9Y11B8sk36/xIsoT/4eZZyh+s5fWNG2GtkTCZLndAXZCmRp
yBjHXmxF2QC2maa6ffzSqLIXLirXAH9wrBkQRgPiGMluUub2NOuMGO/rL81NlIX2YGBxdY6C6AGy
itEOcTP6l0D32Gu0igGgGbqayUR+655bRCXgw0FRtaMZDVdNUHs4vCzTtEhRFVyjwKIj0E/lRtBX
CgN+SP+CYrRU0Fs6jWse5JgJ5IAo1ZXAanu1CmYaPFqLTEDDXfs8qOPeRJSxzkGiP+WhGNXUxDy+
pi62POtXxGohEyfOVyultb+NW1rCzNps34j/1WqAYmtrCuwA7HKipJGgz2OTa+cfiCcAXTS3XQbp
+UXD9Jj3Ivpg/I/FIJFfPaetLYONixDYlAzxs7np5UU5azwOSjOe14hFI+p//u8Njjd0Xos2YMwq
KfQLYzNIdCNORCh1jb7StSB8sgBRqEvd7A8oGH0kFQR5EbMS1HIuseYXRYERGQ+28iSwvnJEE9PV
Ts2HsxQFMhYpXo6J0a2EyV13stSqB4J8o+RpX+g0G0phOor9qC3ZW8gd52EF/aGRgdEUSvPUgkXz
drT7KB7p+TSbN5bn0c+Cux1jJay77hxQUK9ksA6A9dY+sHoF8WB3fxdLN6T20GLdsJ/Qu6lZBLP6
ZNfJzDh/heUWUNy7cbuHHljMWjJHNqLHTysTq21Q0vQyaW6ofO6W6M6vn3oTc1vYyfZIsl6X9sAu
7V+RrD5AWeGgWdGmkXG9MjfuC1HzoZzc7Ke2rSJf5pl2tEMWU9GzSx7+SVdAjYwgIuvd4R6JZ8ez
E/w5P6c9jeQHm72hHJBE5kXz64Kw4ZyJbFEaRO/q2D1uK/wUEvWUBmx1t/MffngFjPR2FQP2qOcW
U/iRfrV5jVqqlzKqUFXRmM1Dm0ObwM6ezcwjwGxBXpJQenNPY1E4PEbHOf8/WmaYiajIs7m610iO
uX2pwcsOh5BiWOoqxWCUTPFEOYDLGz4aTM4IXaEMSKWqpuav2vf8NDDxI9XE9O9mq0RhJrGcBJCp
kdF1nDAM0sVeoLCPnkC82+QrMF2dw4KhyYp+qErLsle6bnqDxQV3fnr0plPobBpSStL4nY/+qwW2
Em0NbxJOPV3CZGMWIyN0sWm+uVI2a1hkp/weKxm33WJrDrS4zSPYHyQw2JNVOvpOsM8s3EwUFxqB
JlrLJuLQTRJhweugRkw+PtDGh7HjlMmsjt8FUswVqPfqFWNPYOhmz2uQ8CtjiquHXLYMOZaLX2qi
EcwhlOvmok14nU5yonK5dl7td+w0qW1fYHMkQv3Q3N14lsih35RLB9opqatCJgsoCwcSTriKdGV5
ihDoRkYX6i7WtlSRyaoiuFG0Z0Qbrl3Rod0i+8xAPrtpbqS/uJXD1Dk78AjdORs6dme85IG3NEVZ
jZs1NRWtXMvMsIF2SY/p01KdB10QktDSwMaP20pJMBG46SUznLyaEtB7wVuy/a5lhcJfddvbni1Z
uzBLatDpIhrdU8lvB+hNTVAZvMTMT0/djOn/PN8B//39YLuWMAg76zeEdkeOhrQYqXd9/LrCyomj
1aE2293x2TR+PRVE8U2emATQp4v0q4sFLuanV0hwbeycvo2NimHF9mjs5c7pdDUT9isOo5sYLDaV
YVnBPDjIX0YzSrYhAsXTwO9rkHlCK22goeGa6PcEr6qAnpQfbrLY8Sy5D18gthEtvSIlh5Nn3ul9
lbKr7r5OhoJ+54ocqnvXCrwtmXVmyMAiWIntcDtVgJuk3PXP66T/U+/N1ly8ig5mBjsVIfx+RYVN
w7p5EAYxwqSfxRcRqgK1WZu+1R4P5RuIJ390rRisQyGnbnSEcP3aLQKzoJ/ptFdEEemzGi338YaB
TsfzB8eALVw5EihSAE1RQbNWKXwkGobYXREXuC/+1iv7F6pERD6Hgwtv961Wr8zGQSq+kD2VUHRg
5Mh1MkBjD8Ufzj4UBy0WoTyGjUonZEoh5FAYxXCcPWjUyVfTcL0OIlUUvZUEDChZxXI9/CxnNB6S
8VJODTN1O8JgDZDDoeX63Aa/TT464uM6UHjw3T4jlmnUZ064TgF8UdF4kaoLNct54d/77EAqX2Bt
xQDY+tBu2iGGAn8+RB+zeUoX8uC/N3gRdGp1Y2XhFQz7Dce2s7V/v5WA6CnQRbstTy1uWl2m5bTH
08vUX7t4HzMrcmnbfLdBfo0nbEySPyP1pbg0KNeZyx5No6Ti45v6P4dkjq1UMSEVmGvR3nYF7E6e
TATk569YctflAIMSGc9yInXcFYe1zCFNLJqiKdzTvxvo4DrobAGpcJvXJ6LVy95b21pxFER3h7Cz
E8RMuKGn1SiRoShqI1j566X2osBI0eXU8KoVH/C+3B+WgY5dAwpAqVgt+62112V+60x5lzi4WlJ7
PQQOCONlS8C9W7ATkOLflV23YjZ2Eltd5QvK5nmeBxsFnQSWwEBRka+4ATtZxSUckcgzVAWKIShW
/XLG/iR/qWknReadsLtOw2qwPBTs5h1TP3rgsxPgBzoCaDV/Yf7BGEkjhFRtpVkzMSfDnuOvab3P
Nz3ADgn9SKeZ/kSJyifxmCNGXJkVF9iGLv/FOb8BSxqFEyLOoYH1AfwQg3Xg+L3z1Eu3ZWBcCEv2
0NtWOeBvdYePiAnEKbKsvhIZ9HyTzh+xSkJHYJFdGoJK4uu+s2dfSBikw9VP0FObl0WAtKc0p3Bs
1hNJWTABrKRtgv3KkacjDektyAqN1g6nkNEvMarsrzQpfiIvk/RjJw4b4RSWzHB9plRqIi6AD/G7
lUCtsd18PLAdXGN2459tt6cqI9x2wPApev3u7UOBpGUjxLJr46zZctPoa6debbnLhsSnQzAPUpce
nN9pDmkRzPltgledT393l9/jCN3W67oOhCN6wXOapvAdFCgu0vWuwtLCot7Fsb0rID72jDeGVlKG
jzBvIssyiLlx2n+kgkdEVcuEyBOp2DH58H9rg6+nWzD2pm+KVCor0ZSfXTXAFkfmVFBRC/WCdF2U
SA0sw0yite/n92zoBOzw3Fk+jBF6mqL9MZpM7cuRPncc9TiYE/lMVcaiS0C0ujJujf7q9l2f+Wv6
9ESuzXxRtmDMvdYM9Ayv67UKwXph+1EjVWRIncoDQkGA3bWtpWwfHxRfp7NkKWW+27TbUQ2mYSZZ
eirt4yC/sqmyGB5VXSg85bITFfylzsMAJfxwRlY9/fE1RKBiSk+u9WS8aBuNGl40VVYPEarvRGoB
kx3xk9GSq6F8/fduHjl0gT9/SD50KXygAmpVGNM2H8kM+5FA9IMTA0eLhr0TTExgkh3WfnZacFo4
HOzzFT7QMjvvz1c3/RIbq2z3Mc2Yk4vMS7FojJ9M0K+iGbeQx9JrWRhvEF3ugjXFVR7LGtCjfBoq
g4MvAHh/mX0/yvu9QYbXSjNAo07DQlFktPYvhepns3kewL0QwyX8o1RfMjHjj+8Lypdhag7LiP0i
ZhfVu0/a1K6aP0/CsVLbLKSG6HAz4RC9BY7I9NCCItkKVMQTvwhmHw4HymTis0N7NW184QC1iI/g
dr+5pYsdbpZYbdtmcUideYDmijLS0AzvKTEa9qtreM1EAwOi4KH2GOTDDvMt/95fs5MvTywmCoUx
UC6qJnwBkh5EUH97pzzj9jg3UfxDrd7/h+5fV33jTFqe2VKGFFDwLlW2AQUFkRSqMIr/2bASw3Oo
kkqQmGchwLj9eNfypVhxxknBLsBNQ7kvmPhNTkC6bzD+FRKwCLN/OiT2XPReSSNLS0iZiwgRWk55
3iO63g63JdkJzPCWfsx8GkGyHiHKLNi1hvamj9Q4oFBsLC0Xa8wjHHL6MfiwmevGHsS4pcgHBYRn
ZFVCXl8cPyDpMQ0C3IxofjANAKNLt9uQYp0RTdN54vbLfMvKcDh6dWHHNASIOpqN74JnWOLni42z
v8cYFRYqXfE0T51u0fXTm/nKDcCZMFmE232FQDdzyowLuJpfBtH3DOMDjR2XWDaPS7Qlxpv8+OzA
bk1/NcLzBkIFSTi699cZ16/mshXIK3D3sdWMyoVDgect+g70vOgmOYm+/i/Kiq4YiSxEgUYTPIYE
gcWa9N8UVRy3GURdo9N5o2ZCgbA1+5DkS+fmbmo9w/TPsVttbzPbFh7jVrg/2qpZDyGffx2WqJAW
/B1INVR+7tDhhLpTDjX6w7x+VAOC+PtKrzWmRcRts/+GPvE73kkVXuwnwa90ooJsVFQt75Rl2AFr
5eMWJXK+6RtWQhx7o4pVwIxGDVEb8i67RRBQZ5QeJLmQJF1ZNnUtFkD/Q/iejo+Go4axPoq+EKa6
cgx3djwdlgL+Dj8Gn5VvVVo/sE4rV5McWGxCJjZhgxhZv8rbMdtUug11yjSakmfa9PcB5jW7jIdo
nIfMUEozroy6se4wP8oxKP1Qrfik+eHj3GQLtlVSLcXZqz8OfIqqR4mO+Dz2mdKt69sy7DYCKjnB
Fs/PvHX9TVEJuA1ZItZozDMSSS+14yDcllYzh6xerZXxAL8BV/tqDGPlW3soZyrJ5bRQcykVedjA
UswTSr0mmHt8DeSfUl+GiaWgVVUbGzHrxkLayBZzLGl+4+5gmiubCKftILlBglF/f+Q7TN0q3AUj
SADWTtm08dv32pGLz6fEtYpVsv2x45k3tYibfLYX8fzN04gySdMv0DpkvPVaZEhu2oLKmfRgNq1e
5xhXujvhfmC6CjsScW0gm8labgsRFpJRoQ8iHJdXjjHuUgbVITVfm1iWHiM/J5MRTsSiSZJ1a9B4
gC9MJv7LzMwCebk00MuPpg0BGq/vaWnq5BeB27SoH0Lg173LFOubOWG2xQKXRXKsNUI6OXS97Nxv
3ogrDviLqRGnjMwP4I/CAASem2EeIOhIba3TR1TEd8DNnwZSf4H+xLtno6pibG2DwssF44kcZx5c
+GjaLXR0DdvgpOiwyrd/BkqlWj3cF5XBPeYG3LxcRe3ZVZaRauezKhBkt6QNut90zr0nqCgyQr14
m2N86BfT+U2RuJA7Bfh07XX6/bQzpIa2oRvSUF8G6SQSuGdnLlyli9OZbOWeqlKROR8aJO0dpNsr
EQ4ON2uEmkBF41kcGg1eMC2Mv1jzvU9NQOFpVYOBRN+F4lG/SiQRoVA7Q6pAD+dljdPRSqLwRKx7
XIjfyTGdPWK4CCv5VDd3VNB/UW7JE0Jm/alNiek6wlIHIZ62L7wPsWzX0V03MzFKgpsbmr1qPkLP
iGUpGZQV73jEdGqs23HxbLqQDdbCJWmDsEew5FwouJh2Ose6HoVAwlSkST1JsD0r93PGDAojDXt5
KaayGM64ShMjb/8axYrB+nl57ewbXWBek27mpE4d1/NfKGFKuHDq5WVvlMsi7GQY2mYUl0dc9v0y
KtB622a03Jft2mPp037pFEoDPlBlyCe/VPrsNsIwjDhkG82lCds1+589nbYT0uVAfx0Cbr55YAP5
PgzG2Z3yfzbAOXSlux9KMQqH39MTk3j35CApTMvunzikRn6X0a1zO1SSH3zYck1yKmXWg6M6xFh5
oe7OIB4KKGuxVqMeAePXwmF627su3RgBq/MuwO8T6MMb3UA8yoOWmhEnHukv4qiAWir27lsbUj/C
+h5n7UVKBaKRuzrOM3WL6fkGhaz6pPHnj4Azp0gpzZzxd2gLv8OcZk7cfizM3Uw2b45U8rL0p/H6
qCwKX6zEKg3KecMDg/lFkQ+CI/+/YpEJY36mYJa+BpIILir9mQYFUyPXwP7WBqyrCSlp6hctR44c
JYG8RUqr2v4XtjdWi0DE+DgduRs+DdIwjDIdezNfjSanb1oUzLw3OkELlG3MD1Tyg5xhsig733GR
alKysoPHdNJZ+vz8xamnDbdMyR7CWuzkYG5dvx+Socg+pOHtb3BLoeNaf2eatvLfM8nnSEd6aeM7
I8CNzIhteXmB2AGWHorc4rf1inLEAFDe7t+LJ6lLifdqwnFqxgSGLQLXDsTkH+YYmQmxa3ObR59D
FtIj6D4fwDc4xMVW5jjAHLqmPXSpLipjEYtcoGlLZY5/Zk/KglogALnDzrQyPAbaCRTuG3bnHAAz
1V2VfGTkUdoWvmwkVOXZYO7+Sp5mOJBrJb/NKJjp8VHIeTDQ2ZzFMI79AFObxRu4XK6lrcuGCpA3
VJ5GqtTxTro0yDRiIjBxs3BLOIVFucDJGGCTXzy5UrKO7PNHIgIXAnNey1Hz4vxj8bg8fcaOTbyQ
HDtLeuKc6XVQK4SSVOsNenno/vsejdGg/AJHDReme+QVM8C518PzQMIstw7sI5vQEnRSlBJekYy6
1/3oj7kGapowJbw/HhIdBYaKjOpwckNn8SQeHfz/Kt0k0Jpxe62snGkRkSoLd0uFGU2ru4qtjCcw
gbSGs0lTK2btqalcHUx+f43HJV5PjC9QEy89a7qKppMmwuUeID9l9Dmg8lQTk0Q9g3hw4NKZbyVP
rls1cej8jsG49p7ohk7nrUL/GBotEx3r+q6QnuAu2lZu9IiwbA+2sJs2TLhIsW4PiJyLFCxO1bxR
RcyDSF5lUW+R3tv4EnwFVcLD3yv53/ciRRMDZ/AKmHnZuor6WZdE7iiMakiraZnhr9jGbuljelcl
+WGBslHXQJ+mT4AFh0gf7uQqpbY7o+E3gTERjBEuSgX/6rETqDj+5SyCk67ETUNd2fejeKfTRJyA
0W71dYOx/jx5HIUi7KJmVobRRXngmBeL/cVcilx3josBXT60DxoO/Xw/W7YXcBDJ1F8yQfTSVqGH
dBQ1Ljaj9iN4OsPV3fXGQKa0Y6btfRL0rfdh6GxakXf8tYcsQw7zio2DOD1RzrBrWF4w5b5kGIrs
32Y1eN18oNPXyx6ZF0drVWwahfwbfmO6mXf68ziGZueA207NbxsZfhbdG9W9s6jdEVBCGiDQ8Hgu
CqgeKDDu6BkxONgcncdeuZ6NkSZgTnaYjcASD32mqtnyEarbin7+EcTMpmLT4q54z+ebTZlxc6HO
DXgbHt+Cs4YL9VOKNaTZvYSyFHzPzJJBzu2EFsPpKQeyXtm38yXkIwFGke+m4AuhMuTNGgqJew7r
Rq9LXkFKWJ+1aGiMe55EmeKpNf3H5S1772gHr6Xop/aY2BmJ7B7XBu8tbXAcy33heDxITAnCOPQj
WEU82F889qILnUwxRypQVYIYYtCYra+zFerkNvzuInUMTazi8cDEYIWGyd8u4xmdH5kIRthG6u3H
tr7ArmOWydPWHbenFHGAB5tYGqJjojs35P9ZtqjkFlwmVaq40gtGezOq47DGr8Rn6mjqWgocmEvr
aUxKvgSwccwJVZ68w4yoCxoxyOVsHzE9lbZ6Z8lJR6QxP4rSjV05KUHOi5LurMOVpi1blfpNZAq7
+SgoEdvCfdPSf8uAsg3fP8Bj9ZYQMIvYkH+aPtavqkfNT/5XfFv9WZzq1f2pZARLivpbOqW+4y/j
J9+J04kn06Y/OiIThG/l1QHrTKy4wNTC150Q2/sWYdsMXZXNN+8BAWszCijIn57OOaNkcPTvFztt
AMXopuMidjZD7JOBDI7dGgFJatTqe6MF1pcIJ9qcuHfb/PkEcByHYGIq7CxcZCIpWZ+jNnWNCjGv
JebpLcr9aWZe6T1kqvx99NEO9l8KChkden6qK+j9SxXAuQXzIWNRJCQACf5uLkLsYNF9LAhn3oGK
W/ujzdxYMSL9ddz5BQHxUy/WMp9Mk5WRXP7qKyEWt9E/X8vDfqzX9Mwj0twfzuqHT4CMLAvM2QnX
UwkyeKZGcmOBK5SMLjX8j1JuMWGoX9wGlE3Zto5cE37n687pp/XiGUjmRmzy5POso5QQSH88kK8Z
NhNx9d1i9OuWfmZ4mDz1QIc85MyZApqtKydUHRn89Y3dnfjsDoA0Z0hSMsG81QLsV7naHf5NrMDc
yEX79+1q41pzEvDF1aKdLKWs7AyJYVh7HzMM0NkJgSPbNFXl67ox2Bv3IXIr9Emd4CwktFYt+kMW
7WAaB9CXbpjxCSzbQp+GfvSEDaf/K4GGp5lGo523Q7x16MdbaOFySubwPTgVpPKmah+u4AaY3zpo
nfuFDdHgid3petbDxgVI/WR4eR44t1t5Y/i6LafoKH0jcX7+IPd3ttGHq/8p+CHU/x122T6vDNZP
PmUsWxpdy+iwSPG3JK5eNqrhH3AAOzxMHUQBzg3jGEnEv1LoPZDpieWhNi7IXR6ol+y6tJZ5mH1f
fNQtfQF/U1615SI8zhh2xBYp1xFJFT0PGh8FLDE6e07Htya5bkkCdQ6LxjMcvw0qliJprtvvGy8W
8FQkdXPWDgk7hw2jzObSp9DAY+GU22EvgNtu+3sv50EgiF1HXxuy2BkVLvDQjWYSg+PNeU0LGwkf
qVsZ0O6NrhDJm4EvDXuszxWgptRGjXeNVrHuNDL/vmguzgjphN+prdichNz3xRz41AEcyr+rlF4k
tgufaZye8ZeN6qQ6AUw6AOgXA22T3L68ZRJAthdNkZQlPVDqIdyOUDbsAy7WBfllVOxXvlVBmcOe
WqakXmoQHa2/aBCt4lBgZy+wFQV3WQ7hO9CQobvSfrypxHnrYVeOLLbKf+LoraHevA1T8lXleWjY
l0830O74gTTyIc1gidlbu0RoAEmTHJKeMB87nau287P7JaRmdCCXsG7HcD/uslFSkyxmHKJi3NcX
qm6ExGRvcuyJjcEosQ3ZQx0BI1c5jCnYMmiU3Ty2eaNURYe4hpKMDVLiT+QszIfEhjGKk3jfoIE2
OmCQtE2eYPYDJasI/kuqsXb5IDpbugFl6tShK9FLIGUTsncPAO60dhpPIMkJJAbw3S+KE87hb++d
Cfj6T4kIqVn9hXk13b929S+ZWa32kI3W4uWQDlQx8o1T6A00JXZEKf7dnxyD8AekfkHDrcKn3vC4
Z49gucDRbgqaL2ZLctmge0e+bMEUbpLX3O10Q6yJL+ODmH2pNOk4dY1twvLLMZ7XX7Ym+jRmAJPu
zLzGJXFDcIf029uMwHXDmAxC83+Tcm8qgZcwXRdVvciDdDt8aqGsshB4/gGFzQ06FoGpwUuAuHpZ
rSEuDnPG9/TdMtASVYruP71q9OiBoD5KnLDC1lV5pl0zTdSjpo15m51fdAOcnniHnAq8ohS8ZJGt
8JlYxkte3OXXZ8UFBVoqHMxp/8gek6sGCcJqdCdTgqKETQd7t1ul77MMHePbI5vbFQoMzCsrxjiP
rHAe25FTSOgly0KQ0LiaKB3c/wHmLyTOS4F7MjfpLLnGCAkQWsOootM/K41iXkajeHtTuiOgDZAV
Yi+cANcLdgs3Qbq3iXiG4juf0hQPKjmNX7JU/hBMM8LUTisncD0lTPQPLp4plRgTOryMMeLOozIn
mYPEk44wzcEDZ99JeDUeRk/vzplRKO4HtBNgdnzcoRTJ36SIKyA1K0BWTVhRHpMU3RHO1mePuBxz
7ZYMhsbUgK5OnWd5sesigTiD545eO8vEjpv10VSOXBdEYKQW+g6q0koQV7LRANS/IsHBOmAvOfVn
7kxmDWBQ3EOZcpPTnndoxPo4dQKv9oU5m3rKVpfuXF6qj+cjOwYi35UQ7uu1Pi+KEtwFdxfpXf0c
D8NDrcbfVX8444kqvZP4NILWeOFCO6xhY7qOtoNiQbYSbiTPT5spo+ChBUrrTVYIbxpkaKYJSztf
r00NZ+Tfu0uQ2sHNjl8JLE3sBHCcg3pVaTe0EQ6Qi9aLc2aLK98sQX3aALlqREdzIMu/z0Xtve+m
zXOMOlB/JzIPIlfsCgiWAuic2kBF+ZluUrvl39FFZc0vgyfg/TDL+tq27WXfVvOWOtp77NKDTv1u
QhOgngOEUHmLk7KqNKSLINrioha4oh3CV/EIpGlJ1vZfDNRRBfWLAQmqphUxNgxcQLsJIaLrtJDA
nJiPhqYjQhR4weL/yNga+0b7y4t1RaCx0Jg7zAeGiG4ynDAzhNdfsaMXbL3CYAPvJe5duPAQ3nfW
cEK6rJIPYZyFmExHZHqrkC4G5IY7xonsh9sIYwzniGwqXidXZHq/9+sJjKPUDXh/hoRYSu+nIiwp
e447fe0mFERqV3XkiIADBqdlhDWXwRMDsJi4wTneloYLEEli9ac84QfKxnojlLXlj0C7M5eeKBjJ
x59lzY+ydS7LR+9sH0SKslUZkpNBU6VAwm81Dedh4cIZbohwFxw4GSZIlSNTnsJwlxNeJfgQFK5N
30DJKzTLNXL2jZLjPBxeZVshIqB3iro5+dZZ6/3JANiH0rbwDRvJdTrVhJFjLPf0RzR9dm1iUZMU
W2H8ltIOHXKGo9r3YQr+s69Q+nwpvw0ikbpUBbzNSxXSYrGy7imM8Vr9Cojb4qlXThaCu3rLMHK/
s0wBkmT33nGvoE3O68d3gfUZz+IwmgTUYLdR6rQdwVR0HLacFj+XDPNGsyBB4der4+2clyAn+t9V
EZJVevt/o11zoJaq3A1wxdu00Yukwpef6lZ29+QTOFes79WksYciz9dRn1t6m8C/eR6jZNP/Hl1J
s8TkeTRCe1j+BHg+qy3lwwotjt/U43RoFGVVzrpjQjrTHOUPNe6kD4jc1HanzEi8QNIwWw3s2mw2
PR1UvpkAwEezixc6+T0gSaW3iQWIdwe5hn98huTeGIlGfnCScFZIPu//QToUZjjsVYMdjRxEF7Wk
Hyk0DRGwK2cTfRFQXXgBQbjHg+23x+xtvKdKNj/wlqQI2y8KbJoFOeWCdwXP7yIk019dOID3YA0t
RBMmhB6lNZcrRjlUhZPlszglJAtjHrGsbXb4UUSi+kYC+pgyfe6F5O9AbDNLtLSXxZ3VYRATH+Mf
RtSq1YkU6vqxmnofqxx8W1BeO0X/V37IQ0ZXs3MDISAJa9I6HqgBmZdL2e4LlZIX04rUMhPCniFe
k1vCV5dCmeiXPHT+4WfVyCKELp8SzEHO3LEalA29+YI03ZZLXiXO/AYjSAOSsdiKY9p37Op/DiIz
ZL17kPN8GTCkEYdRftbZ7vYzWQmEVThIL1LwiAnetmq8Ac3PuFpFALLZEhKpY9qxS9JiVdExVLTp
C+IfefNyEyRHndawdenb4gx7iFhNaUhD1uBk8Z0+l4l4E9HEuDExbDeCBbp0iwYR3+LgYaaCdOe8
qaqKvN6fpr9EiSIHowj1ul3thd9ZccTZc2nChOmV9yCzZsp5BYKb0rMJO6hIvdXEQuD9KpOEuUvb
BcGgOZw7bLeD3g98/f92SOJABqC87U2u7Qo6zUTEyTh6S1izXHRb/n88Zns/yeCDjuWkB+8m5iFW
c/slmA1rDkBaE/XM/v1F1kyl5XvDO2FLYH/Z1TMuSAE7RLNdrCU068raGDHOTv7bMpEuvHuzU4jY
T8K2NgiU2aBZolg8iWbUg/CNgEYoAbYMwbDnXkuuUVA3eG59DpQ9zww0tIjXiXTA/cMlZSahBOPD
U+0+OWuRUcZcjhkNvlcLV6pBDoakoFOXOG/6/FIgTdmesP98ETSLK5MpDD2ByHDxjmq/Czowrd3G
CI36Ysb3uu88blhm1CzJscaod3FHr3xBTJ8rlW4pt6sLiaBlneExKzlqiXKSy5I06Vrp9KGF/cII
PeEwrvOx1iPzTIBkvMqNVgUO6u5HxYJdVK02naqFVbL8vDVFDDLxQhNfo+msZgK/Mk6YoqBbl2KC
c6LSVjbkBZ/i1HkKgjM/N/QY/Qqrm8NY0ImZ9w7UDt8V3Lz8R0rwv3eoCw74l4ENlIEXuoMFijaU
QJ/xisrxORZEMVFyaZq73ce4bVBIFAFvAALIDp2ui5a9GMLwbRbUquHrUJT1A8A91X34VquZk/Ey
4pe2Xo24tZn4b9gXzr4wabFEnAFlBnRD/9bVbNl3UWB2iL8JiRE8yc1OmaGSGIzkHBO2t5ySN38s
5K3gM5ZSDUYcRYYqAA6hGVelwdIhjCAbrsSMaksDIi3AXCXbu9SdW90uKxXkjgh8bRR5L8KGJddn
nlVzNmrYejEgqG1IjxoSzun8kzcgBjS7OmhQQH6JoO1AHTZX/NO7rMQ0mDFDc1CeghTNri/T9APd
hEAB5QCyiKgIqMjcJ0Q0XonrsuMLcmjmKrYYa27m2uBo7JnKcYy+YPkmxzgg9ua+mK/VEIEtNRMy
N8Gmcl8cEI6z9eSdGdOw4kwVLAC20idMuy7oI74uP22uczGieU3+gnHJBvc/e5t/3eDi7ARxZQfo
jDC7SymugOLORPIxCwbWgwlQUuhb0AA+B1LG21g10F36tT4Ho+ImzABUZ6xOvYlKzQXyJeoAWZsb
lWNlDYLYZcCkcrc8Up7qF00oJMBdFnSe3TLWk1jet/irlR7ABR8HNR8pZwAHlhmoQES1htAEr2HZ
Ff9n9lX2cXYsrL42qGS16BN8lCdeQa4FOqh62c094o0gp314h7D4GHAHNvp1/X/frRaLUqLZWXnI
+W0/bhcNTjiHT9Q+Y0aOOZLzEcTv5QkVlngducmbMwenC0CiEGnijx6SKXUjupdcI8+91jWeRRpC
igpRp6QHsmzWXhs+kFpEBvHAFiNPYYXTA0XMOFEKPNl4LYzY1HHaeGq7sOKis84WVhclkGOuYnAO
1BUAHfbdxvYfZ04p4auZkjJIjvxGsTb6Vrl3aiggecTMQ2i/KpXfoFjJqM2wmGPTIoS957/+vopO
8ZxdV7pAUR86svTRKPR+CQNzInkKQpDdo8n7rXeTP4K3jeNf0dBMd6wWoqu4ngv4+e4PHDx1t+Br
IrdM3luiIXa5X6tZkLmkgV9zE3SGJnZ/ER6ZOM9Iy6tYLCiF1WOoKr+2Hjz4M1xoUzjb8E8WTw7W
e5EjfextB0NkrITzIKJqADSidKolehvOQqHwbzL5AIeJOOC1EayyI6gpSh+6ND31L3P8AeZzYL1P
7eh9VSUzhXal41L/OxGrYTZ8krEo3sCg9/BmWWeTnuKqn9erBT1Y7GKDTu63BffPb16sr/IOm1ro
y20jjT7hrWOZqD0yuUsF9b16ai/R3uyAB9iqAAIrlOQAjGz4fQ327iet/xBIVMjaGlMtit/C1Uod
ZihQiN97ALp/LDftDua+lohVVp24M1LraGicK8tlL7wj7y4HuFr0L1FqHoj6y52GxpHvQK2vhUpO
15RPY2GUNuBmg9oBZ2BK7NteliaqQ7ADZp4F58LGo1+a99IzKx9/lAq31oPGtoeba8Uxeclt9Kuj
RgBpNfKjw4tcHiPNCfmZw2I664flFn5hAr6s+1HUcCV/+otblSnHdweOISpzYhJx7FvubyOsSJfH
EdO65ascfjllD19SO0NixhH0jgSWQO/fpKn1zsXqZ8QVX5N9r/ZHVYrgGTwADk93I/YD+LnltmDh
fffI0lBCiALm6AKtiIkIZnX3zBcxmPSnSey/L+FR4hEjuSRQzbqj3LVjhteIroFRs46jFvTK9uOk
64cHOQdN6UYVrr1PMB/LwZvwP+jXYDcHkoEyNVLSiPzelg8Z8yMjiAVwNyn8QNGUmA9kJOlcaV4U
YNz7W4CtXj1HXCbTITrzqcf8ebHDhCpAANt9CGAc7ol+O9RVPiTW1+e7Ohdu66KYFS0Gp/PfpqB3
Xk+ecXAmoBrhzSOebUrLRyDUY4d1n/oQRPWfjAfSEY2qJFjNbsSR27bqB/1V683O8fVkXAW6C4dA
wNFE5OCIxgoQ9BLoAy+U/FTcj04kYpEfoi/6xVpAiITMvMaBQAnV1UQQFCVhVrmwBuIihqkA/QcG
aYNV8y6NOiiMb/FkqZCuu8L3kAiEbTNkjF3vVmCm/P0lbXcz+Wyn8sLTqjAJlQzKRlqcDgJZeFaS
Mih/G9h9hdANB3L9PUJDoOty9vflhymnWLZw2PYR0ta18LHumglaaQ9NM0pM/hvxQ2WtvT2ANake
aO+mNB5BPbKybV9VfRqPPyoHHMweFKUpBVa1B2/bmhHcD8oirZEHQLDwGuSwG4StZ5P+KlFJcyCG
GrhqNuPmBaLJ8Q1Gf1J3ilNe+wFb67v6UWbjLq7iRUBkdMLcoDRTre79SB+KBuxRMOZqZnJ5gW1+
SDk6zy3UUCJTHtcAvcQXZzb+IoPb+3wFKKiWFkjkeP0/GYEZZO1eP3VX7efL/uxcnmtmMek/C8K7
lvUKl5bLcCKj0yCSVaDXKOlq3yeksG51ptJS5qn5BzHzVl54MRICsZfG9EQXawzF6rfo5SuOWGPK
eVQWq6tr5gqxp/gxPSswzEyj0ejVJW67qai2c8ItyuPl2WauGf6gHjLg3Z+P34TVx1O5KjL59oNH
Gp8UJfcpmber5eybfdYZsFAq2DGUxm/Srn0e6E//DLNZUDBNi87h6MA+HhtBOyZb+RU+2qQ7ztU+
QxDvRK2eaICLIJ+j8xiUaqgUP9DpE7/MHdlZa4VtIUx+Kj6uIeOg3JlpoLnxKTVgPZOu7f6O3uXe
17i74sEtsuID4F49UgTRuKi5NVWQvqJRe8OhXiRIW3IFEG0X7ZGH9N97hGc1oM7Xk+lBNBv4j/X2
bJVPMpCN2ZAYpheOS0LKUrCh9xL9jvSy7TZnlW0eefxI9H+5chJJol018MwsgllKbX4OIOLhlDQv
9iscwTYrB6BXuX8rIOiOe9yV5WWJPh7DAeP9DML2Pm+c00X3lxByYKVNBDVjUXUcepyX7ZXed4bJ
aOJ6VCRLATuTqdO0t5G1Oh2x5hFwGzjkp44fSO+YDSfJbj002O6NBhK8sDp+v3499+bWz7wMKjdy
SGXITqRzBN3x6lVd+obXdfsfml5FItrlGB6EoY8CZlsAh5pP+VW7ABDHXkCMPgcKZcmf/GUwEo+7
Iua3tSRo2p0Xb4DxWgzUuvbOIkJHSuw7XMjzORgYuS8d7uQV4vr5wX9Yifwc+QAT5M0kpemQn/bp
xK67Uzm+wMhl1dilZHdQ0Qwd/THYPgLzunnf+kBaFfG3YLB0mcYM8TNN6cKCaG1izVypEXG9g8dR
aJj8/hyBC4WUqDfWEJvqO9f2Esm8lCT7wsbvu262PH2q9mnag6/jWlcyFojKoA+GKPabSAbkn+TH
itidhhwTMvjvL4GP0llwX68trnxv7JZofyuFSyGcH4ZOoMPB/HGE9ZOzT9O1Zrski9fyhHcYuTre
4wRsbUJKtfEf8SjZMibsrU4MLwuwFybh38rmtUwq7CCu93/Gkh0Vs3eRRpbmiAiiqR2TsAayUoOf
VYo7cvD/jK1FBIk0ArCoTeLblVFJoS2hrKDykpT7bsZeX69Cr8GM/7Psna5NjLOlS0PGdVObozkg
0rJJK11wB1Yk66LXQntASFcDpTxddhXpBYgOvJArLyyJylKjh55qu2Aujnp9nL3eP2sDBzLundDK
YTMJssN7vwkdIEdxl6nKQ4pmjKM5Fgsb5ioEnX4r2ozQr3CrvWRDlFwagE2BX1Hef9hIke/niHKC
8M86pEHcTyja9DwJhH3EHncHULyljogfq+NTfQQwGEfLUZXT/s59AHms7gFN97pYzVqxF3PY70uC
gJV1w4gl8jMW5CnxTWzEzLnvsxvVuXh6/9nfqnBt/r0ivaTx0jMDIUnKs6J8Mj10PkXEhfH2KmUC
bqoyICSoeju9EijPUcBEUDfCK1HdJhHKuPwU1sR1HPQicgT4vGfz8+7duvtYE0OkFQdrlbl0ZII6
l4FMNa7TuQl+Lg64Tt1RAoCsa0TmTnYDRcHbgi5kRvGsd+1nT4nUDQ9DUCwTnwFMu+lhkixliCjm
3yclSeFrxvrqskC9tLULiPw+ES5KCGqx9Qx6+wDI/YIRSp03OFnS66BFpyMdbcKLkMEcjL+3ZYqC
xA3VH29E3w4RouLssXySkrCnvKtpSqLa+ENTF4k1NdxjS1H1Wk6VQHrc9xsiPPThZcLwzmVAgKNS
YaOYbpNl26Pae313B8ppADaIWO2dG45ITpxMNidaWSqwI72ZtVH0VxUA6B/QYRaPDXRxlwZvqSzD
upK9ZSnMGZFKnkP5q0E5d9a7UnIbL+/OIpCO7J6xVLd1SKYLfsgycb6+kU8Y8UCd5Z8L7k/T2D1U
kQfDMm+cMhHMRmDZoSxK5KSwWtCS/kXPubBubk7xxKOzzZKBmQO1628eQlAFDHbd+rLTwmcTsocZ
P1UxJkfWJspxVbHRBEDyYeKZGZcqb2trqBl5xqr1AZaHMxMq0aNqeVJgZn2PSLS1+MJDGGJz2ZGA
MX9IhzR79xAKJYkJ4ZBgdqV5+7fwPfVBUJYat2o8jnpDoRBTrLGkXRwpqv0ZCiIhzY4tv352/IQy
GyCKbNDza96aVva3dnBhxakPQ8qHPkMxOu3WoUNinbVVXrp0LCmtzNKCl0MXjHrYloZFqO7pQwrn
ZYB6PE2tDmPpPmB9R/MY70k2lwaSikc1Pw4I8ZhVKVCnH5aUMrCeeD0iESv6HJyAY9H5e2f5FJBu
YRu1puTEFSJSq5ZaKuWQ8rF5ipWM1hW/vUvZ6DpExInm47SoOoEQkjZ5dQvgFaE4qMfpZKWYMhGx
NW249YGU3KFmzXmwPnc46axLY/1s2GPjNyVQ6Bk+jaZL3F50yRM14ldCFKKDDMCMjdgf7JL0zVb8
aMBzvsNS6NSi4+PsRYKQrsbF73MVo7qzrI5DM/IILH0IAje5o4rWxS6fAqRTuMnDXM95QTNB7skR
PAd4ZH7qRwjdHNV5x/cIsyRyB5/74JMYtOumgFquKfrWvJjQdC566iWWhDkxiBTlJ17Utv7EZsM1
cVVk2jnR6SWOTVNPKQ9hNm5KtNZD1zFX9rfVsub+Hs05Z8PqcW1o932ZoeiYn4lW0XbsgiS2WUh8
eGjCOiPGSP7Rq8zZXC4ZvtcDn3efwm4cY+o0vZ3/SyVPtcJb1zIs5oNU1r49Fphu+X3TULgKsLWI
WZHH0u3g+l7jRSkc4zMpzk00SYteWR5WNvKeyxNlCWlCmdqvXmO/eBiLL5mi6WIybGWUMm3CLQiP
DRrepANaqP+22fnsmqUFWS4j9ssUoDGGZex79j7i8Ek/uDyIeoylZPbdKTD61yfMF0kIT/gh2+Y7
ZohvbCCGdQIhWSJpDxqjYtnDBKGxmlGbSfcMON/3cgGuD+XhTP8vPG63Jxeydaau7rKmk9S6woEA
hY/nhBtWG7nF69ytwLk/zen3ccJI8H8L6ncXUUviMOceOMnQWCpDdDGsqEs4x6crH3//CFj7x/dr
BrSHbV9waLfXv6bu08qgFm5gWEsaK6DDj3Vzj7UbAWB/AegSTHPzBlOCBkzaKIwpcOZ7EY10LhLL
ksOuRc/cpfxZO6Us/IRfVATNH4Ustep2R0oRKMGgwgq6yWpo14HIt7/ydFJa6hdpNnrqvsELPVli
O2JgkUYnazoydhxgFqqH88fNsHN4uPBzknN7cQ6Qp0MIQmKOcCMfXIZuNtGHCJzEZpbX4Lw3OYtL
6Y3Mxy0NK88hWaBqc6bOpBJw7Wf9qAJoKfMU11lQCCsSwSlCu0j2gtBUtlXSEqGm9PotknJTPlGd
vvaOJ/TlecH3HcUNwhD6JjoSV3nvSpihIXuwdsd8IrbAVp5k0MkTLOuebOitQVQiiDVYa5TwlCee
Z1OIlZgPN6pfs1EcoJ7RlZU7xbc20srnjkCw1gP1hZCt1sRFHGv20QRl0Gl4KeD3giBL+a/UvTCP
mtyXnXd11QzVsBL/Sj+sokTuCYf2hyiX4RQjbR+xgPzNqvFMNDoeUXaUcXc3ruq7HNxptb+PlvTz
g37bhycy1ybG3bmxcGXdunhTOSTJum8aPLxBz6snXb0VF3L7oTYPHSQtgiH3kbZ0unSVUPHE47lN
pkKd+vf9NeEIn13lJDfFKnPTZcfIsZ93uJHW2Mz4mVZaEqePCWLQnMxumg5+XG3zojbvo+lUKsMN
lvTbFgYN4OvaEqMntAbleTGQVAdyKYsP5yU1vk489PK5Tby8wc7yfcHJOv8hc4qPIqlYQCdKPIQn
HnISOAIJ58cAA9Jw+NqHlxhzNSvfGyCkdS+r68x44C85D+IqbVdRZD5fhH68POG4gj969wzK3nyi
CRP5BMYr5Oizd9UktEei+w1yY31sViO0FMlr27BR0nxoE0v5P8ZpEmYG387+879rG6R8bj2MF7f7
v+5atfib8zu/BAeI75Y1UdHD9cFmkmpQRmz91gb37s/IFI4C0X0T00soGyx71AtR7VtLiedzti+F
3plOyVNi0FvwerX9qJjMEWR8+GHbSGjH+p4viWyADSomnHbc8G8EB+86ty6+BzfqVk9VJT44q4nj
6OEyY1e5qRXcoRCCOGYBlAnpqxxjzC+Lc3sQfvZZfElYmoai9qyDWuAF51hFM4A4O6E6r/IL8jrG
OtwgJYx6iuQjTVEbJCbWyy5cq+lCwpkFXzr1ShO/D/0QmdF0smwiyR3BWVsBfV5lfa+zVbJyBczX
jRKZnqh1P/HFV9D320+oTTDZ3Kgbsffd7u8N+NrNXJQ0IvdfiXQBGi8PtgAzkvvQJNAKBwFB6XW7
VZvCDFjaW5FnFjP4BECvT+LOTov8KkcuGMJoAEIb6KNcghj7n5IhoGCBlD5bZbbeJLW45re9ipRE
W1mh2c0/xDwc1QtlwM+IkMHvOkQrpsTeB08YOpf4NoapzJhfI2YHt1IdnoNbx3aWsln16Fz74NTl
272WSXEhJpLrLvASdm8FPwJMa/99fBS2bUqwJF7dvoV/iqkmwjPZx352eHh5Be1RskkKCWtDZOCN
XgTyGRUPfs9vyzv/jniAABckfKHiuqIfyr2uqP4pscCkrTaoS6DjTWr0n5Z1XhsfSEAbRSA9ccqh
ZRwNe97+UrQ8vU8YYYONCkMPwESm7PtultDqMbmIKh3KSj6OYQj2BN+bhYydIxAUFR3ix7L+JxZ7
ve6x2qF4+5r4bq4Mhu35K8DQSvLHcjgz6ap926mLFOlr00dwAUDwOv0heTnhi3GmXf6hqQtE0hme
DhigftVSZaj/zR3P23Z3FxnfKHxnDcALNNxDDlKiOXs1tX7/2UhNl2n4xr+Z7IlY0AO4rbo1vSYH
mk/MLegtLmyYDBjivv6sS6bCNOH4IasO3luHNvSXT+gwd7+2wBqc6RhOyAYFtH/d6lMell7B82/O
kXgiJuY4LJ6NNa5YSAYOc0s1NHeOyvms6oQ3LuUrh4WCZ1GwopRlcUsFTYUS8oVM/eB+PjVJB6mJ
BhLN4HgXGrtGfU5hdQWIG9wy1EY4QucqzDunmTqigT7bTu4iz21638YW9Fp+EfMXUqbWLK8vxaSM
4++T/97CzT7K9vabJnEyZWKCNtsQdHrvgFYVznfiRtzZcFlrUQ1or1WA7WigX/wz+KBTHpxMCqAx
8gU8QQFU9Tl938RT4r/3qiRY2g63XrBUB0LoxBtn1Y0dnInRphR8/zH9YRPBnktMxZCAHqs0tVnL
yJGBfKKsYqwr1zLw2TiGRzykz+hitUm5KEFSPGV7tUI6OPMkbI+6Af9GWDE+lH70UY6wOLC2I7xJ
Zgly6GLYTWrDSzwlIikVgaTk4ODVmXJFsw1in84/Wbev2AbV/6zFY0PLfW73jR6/s2domUcTty91
MqbpuVgJ8+eib19/Kn9BAKRj5gAKn4HgcGdpEbE4/4CzNZMpyGyHKPNEzn8uEeeoeCJ0CXbMhewV
mtCVwxL7FSaR1bMUlWh3Xl4h9/LFc0kaopni7snXvANaGoKoyRW7WIXeDpygQBTI+xMJs+s3RLLs
DSxkCwAIzFF2w6kV6bfAhOu5AfgQ8mkpl5fU+aSv0ITntPpqE6cQ809mjv2oBDHEGIxS8/pPYgv+
ilF+9c4ey24NLnwSS8lrOqq7YKpLeW8FNGBxv2Atne6LVipHmMZgG7CylxsEMxiJwOX7wtTY/cEV
+5pBGL7uJkhCPOhmRlzL8bydUV4t9ARRDqUv2lMdX8sR7ffDnckoh+2cviYQ+fwKZCwlqRbyI6Gj
JuTpOXr5CX2O9ePwKU4ILDmQBy+Ik9XcWHmXeuGBmg6tCTZmM0Z2m1Ajh83VULC4SvOfWYQSiUKW
P8etkZuepF7vSRIu7coH3cCa/s20f7QhPPxD7KMgLoidNojJP0fZ/VLm6oJV2w00QuFftWLkF5J2
QGie9JTwTbYWnI8FmpwETQImJsR7NuOCxeMaO46hMm3QGUp00Fw/mXlKSh1m/8JoOu4f/HbMCcIK
LgbN7dFajPAJJ68SfFks37/YlqfsVFdcCnfZSebXeB7KWFQnbiWyr3+LfibVwDlRhe9jrUieqq+s
BJgzm3OUc6XReXvsrkFk4JC0CR/PdvYUtrWe/nSslMlksUbfdMJIIS99secVOqdYCN0ap5jQYSzv
nuZxNl+vaKV0uGQSeKWthZodolc8asXEFhKPgF+0hSHqX47/fqleDlfhwJ/cdiKPkNDwRg8iqTSd
/LhaS0MxK91Us+24V7soU9SYvorTdD3+6TjLT86Kn5EdIr3cCl62yf4ZqdAnxEUodgMwxUlK3k3B
61dqOcQbwOKlH+Ib7FRDcaNYBftwScj9cmyPEVBk38Ex2FX97fLCBqkm0iW0l23ABRELLAH2MMEq
875eJdlX4QUbOfNUKJjK0T2jEW6dQhWWel0p9wT0melq7QxIKZl3sVaUWzHywlgmPUFhMaJa6M1x
v6PBuDN9wjUA3UjaA+X65wK9drNYOPOkYPrRavGxCybKoqacJO1FaIoEdr+iBWrbd5rUr48kvfcb
q9HKeUnaOLhQDbjh/UoInrpx3LKO55bfA6e4PmCB8abK/eldqQMa6rRnp+ImZBXdI4xPhWWUZhCn
9fmJIdjy8wpCkMTxQ+6U/NGJoD4IMX5bJX6qzmV43mqL30qq/qH3mRl8tc5cwLjhnkXVjI7C8b5X
OgfB9PiOXaguADdmZZ+GE+p7upfH6fBqT90l/VyFMTGiGg7yszNKTXupS0gG+Gv1ygmcfePYwscT
49KC/20pdmZ2Hi0S0mjwKotT2OSP/1WxizajDhu9yaRx6jIlcPfZkzHoV/MB8wgghexqUaUa9I+C
bFkFJJDkTcibBqJKzWFneE+4J3thTCI5BWuXgt3cduK6MSdPm6Ub8LJEDgNliMYr7Z6fj+/f/IEC
A4lESg95wBuoJoHlnCbsajU4tCXYTbyhnpx1/sj0UDab9fuPC2k6fk0/G1o/jYMz5VB0EhEx7Le4
PWRE4+PoCkSbLeFK5zfUdR21Yk9Gtn5c+V6TO5hcPLwQV0FAujTfxryD2x8VA6w3Hln5ABPLcE8M
0jnIohEGRqVATTMXSSa88gNGsnPhEPuCqkJ0yoySuGBiCcjjO12S3kPiAYIXUGEnDj74neZ8tr5N
jKemuqONF+owvf9WSnfLclaTr0v7YY7YgtNAWWb3MoUcBeN2g6io3tb5RfaYi+oHYbjCAz3SAhkz
vg/ROuUcfqBl8nZa6cWLMYvAErDM/B4y8sAAnoob+g11h9ItNHOU0laPy4x8Ma8Rp70XtvYopgL9
YZsmcORsXlzMyrlcAOTjvVWqlLsKjKRoj54ebm9OUmFBk4k6ng39Vg7e8/73McaxaGQ7XOmK9HOU
RRUU9i4Xxy1XG1knH21t4eX9UOejjLqmDAYaWbbFwQsXU08T4LfteUQ6fxcAl6oSTfAccfQO7Cwj
TWqPoVpoQIYF6pNTjfGNaDjUFSHt0mcPdpk6R4rbUvyRd6+fUTmprtAZ5hFjA9WEakW3DcuZACMc
xV66stqpBkMsh9j2T5RxSQLmzoI5gPP59jgnMz/MdJ+jZv/GxJpMqMLu6j8yXndvRddXKHQcZrNh
uyu/JlLuvFftsq3DIWYaYVf0uyKaPZ4TclPtDvsjctFIlHXvHefw5PK1n2hSVexmKSWeNn/Q4ov2
U2i61m+P98GGq2ywUi+w3NV9KhhG9eWxxAwGaSLWT3THlBGC6PVdoX9Vk8Nzp6EMphq8UrScEB3q
lLKDIPiJTTp9cN4J+n9hWXfNZQMVaIcGrbItxC1VQjmouUY3SbBgMpwyG0uEDdiGYBXs3KGCoDlK
n4AFy1Otca2reAOJgqR0zo2TjkXAWJvxDM7RgGAZMfFpir0oyfPc6wPKvtwCCqjkNgf/M+HGeQL2
OdfCdk3CXkxH2upywKRc+beKF7h1pyqs5eh97QmczrIOryqnzUSLIzrlEBPIwjDl7M8uZvlYbT0P
pNuU8duvxWTar2+9fXaGTWPrmoJNrNBlysS8aoboB2iIj8KH2Kq2YqSAKCu8ekHjHj3PnPX0kQ/y
w5z4FzD97geeShGsITleND328dmmzi2kEiIbirs8UDeKbUSuWOyyaqDnpdqY0l+5WVTTfonlSYOo
kvhZVIbob7tpLh3Zch3GMH0mZwT0lJv1aCunmqhByy4myO9XPAWfkOtDbYArSKDy23dabimNJJsM
XWwELrf1PCU87Z3jTmifxslQMzV1FFpThsjTZgSE8SNORHpEhGZX0ttO3mgUt3rzeLwfO+hzH1QF
I+OlWdedFafqX+8eHf1An0vQhgg9lMZ6lsU1cAHsaRU0iwuI72Um30jcEnq5qBUFG7EG5/0yPyuU
z4GcGnbyFBMywnzwZqJLYNFb2jOFUk349vKkS0AFaA6BC0atkl4G6uLJSUNlA4VDMtTLt3O/S0nI
CeK8W/p5CQYKyGVwaSAlTrFPSIDD4Mxc+pO+0nT/poRujeojBjN9XMVLhlSM2kXiZpBexyPMT9v0
Kk2gi+XTS77qK9EjitL/nr4pYrDVau33FUGv6s4LqwC+CXVBsA+FJptrNPwS6OuBkW9a2KT8oKm4
BxLp7aGv5Orr4KyNYixoFuYopprd4DUFwVhD1amP+qYkzPwERitReYk+WSFSE+461Zv+a9pB5Hip
z87mc2zSQD/ZC9d3NmYvCKRO1oQWyTiSSH3yEOUKMd6a1IPbP2FAkA6phCRVmoncRG498RlNADJU
+M0gkVTYLCIWEWqhUIwiSCok+cKDGqjzw2Ti8mBk8wX9OkwD7Z0c97/y4YAn7U84ViZaC67Dqad2
6CdFCLDcB1KcZX6BdzU3vs55Dfy/bimGpEMQsfbwdOv2Bxnms9a8raYf0sdw3kjuSt1J3q0WML15
tRBhfNCIoXA11dS7GRClmLLqtnD9IcQbr1ZjpsUki3fcwjgMNpcYCXe5t5G5Z09Dxqk/OyvNV7fy
f+zcZSaGMmYTYIuzYyY3yIGTv5tGx51q4mzHvIoM6uxA0rL+SH2g97pEgjs6xnONnWn2QihDnYoH
FM8MB2v5v46/LM8DuDKje5rklbmr3Hb3sJZ+dhte3j2N2y5EgPILeq2KfSIlVa+Guk3jK1rQnbil
JF65kCQwStrKAruQCB5byF0L1tTM1L7a/XAMz5KJo/klnuz21aWDwE2qw4UlxkI58aa02URYGUhE
SQhEInUlzOJXFkE9GuLl8nEyQbiT8baxVIAdIqgN/J4LKj3OUKy8EwDmqLGwkFAZhZ5pg24UZs+u
wWR/3mJbgrNTCpj2ZIHA3pmmgmdGStxgat8biSI43lWB9pCO9PVNFZw2ETgCdoagG91b+ak01kVO
L3O9edZ/TxupjUXIy0YT8UC+XRG7+MuI056dFybtp+aXio0lL/3WoRJD7aLtnBEEcKdBOI86Zfi6
+s0PEoSO4CFWZx8jnR5vRyMkQIUYunkOqQlMVK0CwXSVEiwrLV4MVwKVqB0X2BFydVVpif1bl4Vn
C3CvnnoZCAi/p1K2nhJOXYYqQhb5X62zep+o/q1u9jx9EGT8LDwvl59mhzMSQyHrOF5Ew2Gsaoe4
86fqLthK9BY5ExwwpaTaK7PvqhneXkimG0ekwpLzh8l98fhtjAQ63Ym3Jo3IDnhnoHbbt+4GZVb0
Y/UE/Y8qBaugFe+R85XHXMhjRIybhUyufcfQp/SJ9KOmlcSz2FgvSSQdwoadcoFSwvV79Dpn1W6Y
A0pe2IHkhv9mFDbz7N2toF53NFUhrjcvOhB+MFtfz0odA3y6sgSZac0AgZtsJdwv8qfJKfPwhVZW
tshOxem3SsZYQsBICU1hqggm+RT/YBvB+LFkvCWA5tEm3w7P+1qeA230CGfxjvB7Us4Jo5vTOMp6
pjTUyLjEojSmg9LWPzsA6Sh3u0aAY/yIJ8ibL6tydji1MCXFKdGc1HMdBKciRjpdGt6NgPy6M1bR
9eq7ROvFATN7UpIWEJthrwCTexUU87iWq0tx4INla9h824fdGoZDDGCqgOhUxmakKtm2UO9Ne4tN
a45GO+0iFNGxkmxT7KW4ef7s+9DcgmZ6XQP3nJPVVthtWxF8yLUargq6u8SKhdZK1xwTxfX05W1M
rP68o8yY1wqKieWhuMi685dNHxkoEzf9AIjg9Jn2MtdirnFDHRKYHMppYlxR4nl8NR29c+sOfyST
JsgHtrWz8fAM3aI832CVt5MdHjrTbdsRZAGVc3P9uNqtip+rlDHs2+2BqlbWK1irPdk14dFdP14A
rCQV2WwawSMbIS2tES+GBsE84CuzxSlbli6UoKN37/S+kCGx0WPgXNgza16HotafzugNTtMt0069
2P5FAZW1M3LA3F7nFn3O/3OilX0Rw2hkWWWj3M03ou46itKsaLXaFiVesAglcby5xCyAJi5z655T
jaudz0h6+U9mykjMIu02PlzpnVbfdRecxiOTUWH+pnEsj9aDIm80dgnSxtdA2kq9MUHXWLIvOKU/
jlMvznpoKcRq3pAFlGHN9blW+f5lc4LFVQbY25vGQWmgvhBJQ+Fl06CzB4y0i/WHuwijxzUmKiW5
qPa+F5H3IfX0juPcEwguZ8aelxI9+w4EnRLftRovmuTX08rpk6N0bT7PLjYaedeoVm0QwzbsBBaF
9BFksKyq31ORevtxNHs+OFfY4zyXWAQV2VZjUuUMAfa73eXf3nkEu73Yx9X+GPSGluKlV1RBlIai
2qqbb+TC5HSPrf0+Zj57SOX6jSYiobT16OvaWtB8vT1C24Ag/4cM67ld+n3wrGyfmxLWAcZZ/SjD
djFhFHDto1/SyuwqLyIhAKMXw9IvXLH8Ta4OXgCI8Icxj51zGsaOewlEfRBrymGHDKxov1JEimMR
V5aJ77jP8hxcYndg0tWzHg2KMR6nnRrkdhwqpVlDEEaLhbKOYM1n4tf/msFhi9378q5Gpt1/NtU2
MeB8cselx5UWy3xRcS+/xCpKoMACHaa25AjaxKsqmlx4TsW2TzbdUqW3oEEf+ecKgTthk0ewlOWC
2F9POKQAHITiBtJ9cRsvh1ylO4W+8b4UMWSSZNRdQWH90gP/Jfv/LARwbaGipFZgidfyEHF3ivpU
SbI5986/Y4ZbMHSiRteBKSPB8S9vF0tlDLjmxTFiAXa1/fgKuGXwRJ84BlvYwqhkfK5/cZ6DeNkf
Gj19PmOLSKVLutC0Lm9uSte7SMLx+PuNDEzK7Kxr1d5RSLilV4NUG5NNHoKinExzkDaYbFn/YiJ2
WFYa3nVulPhwyO+TIGlAf3wum7cT3Kg0Ywz4l3PXIyevxwF/QJKy2KMLQZxmizSr5b/VVBgD3BZ8
ZvFS04m/9iG1m7lFUi94cRTW0y11iq0nD8z/XVcoH1RK2HjUF+Ow1IS+lSDsjzeyccRLl+jbK7xP
jW9ebmtOQ13WqZ6V8fp+CrPDUIoMP1mIIjIhUbaifQL2KgZnF9OQXJXvf7LeVv5cl71liDgMq4Pk
Adxw7cjbSnZ7quk75k17XmXjd8qdNbNwuosiKubr6r5UyNa8MTq0b43qHpSjW/fHa53JL8xGfe4L
UHqxfLrSb9jmwsTBJ/B4sSve5tP1I3c75oeydIppsJo2t3rdigeSJcaL9peW/wEG5zHe2tV/ar5z
/n836NQMxy+wKXJzSvoKX97pcvo3+xC8Jq9v18S3d7RxodcfV8e3CrKViPTP9+hXQu5NVODeCOVe
qlIxTy430gd8vAwPo1m4IR5FJwHLBfAFcrVZktQBmvQHFwD8wOhkrJsONZuFvhpNWfpc7UvahyhV
WnkluQXJBcmAeSpDaaOX7YZf4c1mmhbQsQmqkjHFaj9ViIbdpUm1Rb8bjNdXT643lsodhdf9piU+
Bx/kxX3LJZIaHyrZdo2PUzFSHuKm9j6MLXwGvTXhZMrwaIaYjnalo85P2pDZy5JLetUdWZ47kCmd
SkDmH/10uRwX8KXvVX22XWNEANpGHW2ll5016uAI9UZytJc540qC7ELtu7Ep+Iia6jvk/R42Fm/l
/SLAKYeAtHcJtQ4suo5jc1MY+IqetxOH17VkZzezVd5RpRMMCBI1GKhhYAAjwk5VYjlfP7adBLbk
7UPIAkWRJPm6U6CgRL89FeGCm7e2Mw6g8tEBcCR6rU4AB9/fmqobBH6GL5nKDmKZVr0IhhfrZ1sr
TirkBmtRUbu17To0qRDtpCd2pNpcW0bMZ1HdZyvL/GoAVv836nSIXi8ltCyvsjb2+bhyd9PYjMGx
F+ViaWkWd42FNFBciDQYirZTjvFMfS6jyGK9FRSogi2iQBsXFhgbbQa+noNG+5/ZaB62oGubdItd
cVpbKfHl7tIM/RXusn33aqi+MAxZ1G5HLPG/RQiE/qAOCqXuJWc7e+KCvxnAKlIImDZPMYDRZEgH
RgNPmgPj1mo89/yn6MouFmAAIBwFkR9ZZouXWZ8EDjz9YGmOxtgDCwgN6UoN9vtsrfA/lIQgmXDB
jVgH8Ps7L5jwjFK4/SuQbX4KdgGGYxF08Uw12cyLVrRreAdUILjTZ4u08kFHT6c+50IJLGqpiuR1
XvQk+ZBAzhrzTT+j6og3zGzUQ5KU+KzX+Ds2SX9tbHJjSzqlOLnKgCdHkDMgrbtKrFfSEjRo9mUE
88Fy49g4z3hqnzt1Jk7+wkdvBnOKtsaA+GJoerSpT8UQiZk4evGegiNQ1kspqPY3tz1fUt545DaQ
u+AOapP9E+i/bGb1tkHAMoZvrmCX9Qubf3f51PCBS1XHHZ0Fql7J+ejvYU8IgB3OeitV66/47C/F
+7ehVzkRn1QflG8GyF9h/99GC6flmUAtTMEShgVn4V8LK+TEykO0dM09WnCTTs7B5MoTEYs/J9FM
mmQ3igxHbVvDZOZF3vkO/USJTj32Dwm7+r1JnzhDkJoFz08NG4I8wBBfC0QL3s44iqipNi2FqSa7
j3rPoKxQvb5hIRo/sj8F9eA6B1sWvQvcBZ3ghI16w6djCosopeE1TL+JGjkugNIeQyIOD+LqXMrm
W1MrgmJh1P/CZYOkcv6wZsMEhncCEpnciVEuLQ0TOyQqv/gyhYy7mwSqbDsC99nBBJw+QyFtMzkg
3xqofwEXJFOcJWk5QzEZrclzgB2nq52kt6+gkuagH7wsNtlto+daPvNMbjB9T9gqWzwd5MnLj3qy
oBVvTANGkSNrz6mCrz68e9vIfXfHNGIWgjZrRf4ZL6lfIpzMUifHcoDtqezP9S6hOujIiOnTfL7q
IhX4X55FDRkvnJDrVuW9iS/OlreS6/OmJsYFFLwjIu2xDeDgtZn9l4WB1DHgMCW1F5Aj1qWsIsZ2
3U+uppcojBSZWN5Xlfk7mDjQ0jgBjQMwmlNAGNU+n/qD4qUkvqrdfa+9E6g8J8pvhTCuLM2woxVh
8KaSQv5cBnbZtC1mxTGiCpSeBxUOoOUZn0CeZWQ9M6B3IUNXWap0HSHsfF5+XSDpQj7hjpLaub9J
6OraXrqMWm1xfMeqtcO7AbOWiXkBSnwN2mJivS/ADpZXjtK0USbWSJ0G+aSrnsXiSuc+6FrcwFUD
LKrkAyITZGqbDigI41yktWee/+0yd6WwsiwTSXNrK673yADKaoBK9A3/mPZg695GLbRJxf6mG79z
8TCuyr6jXaD9M/frQVNIir3tLeQa9XTK4u/kXNRk7WjonkCIoITVR2iIKNiavasxeiz/FtvCkyGo
vEvwsQbN3dTjm5Me5Bd4qLB3JjZo4GKBnSrxtrfwJGZVrYsAODLXn532/fvZCORHr7QSBMPVblmw
p/800L1n7uZ8QpQQsCGQ+30UbF0hvLzEB0miySklodUnR1+/9+zebLpRrReQ0laGPdCqhIE0VAwg
zo6wpg+B6yMt/bxGa9kwZLFA6AQlwn43hy2uZOCkRc7TCYotnfe5K1gzUZanmI4fWlehe2m4FSGb
2V7XCsB9UrT2+/qKDCCSvGJOlOX1cIE7RebmO6ClBaPG//0X4kLU19MEsj/M9ySFMZrgDcyzV3Sf
WJvrvWlBkEte5v40e8LEr2aMYjhxp/8fV0UZPL509QBcBDdOfDmgjoah89G5dWbvoxFhWwPUoSCP
vPB/i1Q0s9WeEvHNrDGLlwaPBH6puUK6fw9uQ/D/0JzWV1xnRIJGpeSaTPEydkMsqHkrPHajBtmG
hxhG8SVOVFfZf9FsMJdCpALauqDPdJ7lW9HPPZ40PFKWTpd9F7l6+DkwvikNZt40w2ltBQ12Qnw8
XVMucsG2mKyzuQtvLS4Bo7TU62zUTiMslFp9uz6w6abB99w7SqOgYljzqPMghE/z08dYFiV3Epm7
hP/hAkkAwAoxI0uxelyA6Nd5MbTDpvm3n2Sh8BR/CAGwfG7MuFLXxBECgppEVBPjwE+GdHVnxLST
gKXGMU2AZ945rkifv7tL0HuXfiBi1ulOrpUDe2SFXSvNB2/alPNLB3b9VJTos/Me2IWwRXcozfmf
gzs7ZHHZmg4fJC0vESGcg3BXsWtEmNXVa8ICVhkUHrgS07jDKaz0a8M2iWYksuKK/WAgt11Rwbqu
uPfZ+bApJThRhytgsclp2yvhi+zg0xCXQm+axK4dx35im3XFFOgHbQGtY42AFL7+xrgjQML4O2KT
gYjGJYxierSxEq8641zudr+4SRY/6257euV8OjRs52v5zBhIVQc5BD8lYYXPqdm+KmB/jgkmGXFz
pKCGt6TDHBq0AAIVpxjkrabrTAhJaZatXwl08pnV00QMIiFPM9VOYdA/R3tKnhBHHqf+1d5FnwAm
WDDmiZDkdTCJnyxDRHlnj2vXTWT07DoQAbLU443lPs/aFh6j6x5IGNycO5ucb2PNkC1swIDmWBWj
0aBCUgGNfivmuU1/ngQk5PXrHkjdLOW8xnWXNSdengJUGAbvY9EgrG7CgdvEWgMukqcZEVM1rMr+
1j2hwNbnSenTFmsq8JOWNVu7l8SKPJC3vTt5C0VM87ffMlLiitalQNTYu6CchbNa//5REY3/3euB
7ZszLoaIWNh+XNtOAykk4I1m9vVBjeB2ZDMlYV019cvJTCE6DKSRr5Bi++xWB0VN3e60qOtKyUeg
jFBmXo5/O4KVBshfLGLItgitgDPdUFEAy4Yj3iBSoNoFS56lcePKIXXyOTafAAMDXHmUpMpF5H7k
Up3cjCnaFGgDG7ZmmJmoVfBX611BpsCXm4ZCu6z3qF7kUafppadCDFBE648bozfUF4JfFy3CKVPY
+mVJX7Kj+KkKmK5WBpvo6blYdqAvzklRUIZvYYv3OG+kNTnlNrSaR2Ewqch6NSj3jTN/pf9Mf+ft
ZsTV6zXF1J6svEZezQNE1NeM46C8tAlznnzd3445m2mO540bhw2IWuaIQzN2OQUXATHQkKkSn2Fj
I279kri82tTqYS1VBisvrVYkO6L/CBa4j6Vqp6WKygIzBWoRYQZAqzgpgTPrIJKhdsWK5eDW7nkP
kVvqhEf8i3aD2h86l3tql2BXk5FcC+w/J+hwznmKKeXIJzGK68HLNbvZ+UIEtisGwgvTGnZw2m+z
9vY3C681FTqGxsTTeeyv5I/kJ8LuYZ3dmpoZvVOSbU3i6xY8p2mpauGYs4YkDhA0vCJsjzldgFlC
WytVk1ke3qpNJEHbpuWdhCMfZ5cqOmdQPTEV/LsrYxG29uZCbubpz/N6VC5ZmftbatmKJwhSF7g9
xMlwcvET6mEFi/BhHTjCy4Fx07M/kY+FOrEkLCEg5aHVjmqSXjXBTaaNR5cCilmuxQCzH1/TSkde
1csFJVp3T0+FYbghITAyMhftZ93vG6mSBkvshBk2JzbINYhFd0+qZ0tz+rC+NGQ1gxrB2tHteFcn
FJoaXPAIH8Yp+cJ2q4fnwCEMaERwqQgLEOP2yrdjnuAlX4izAiHbcMkECSAYJMpoNs4ZqicOuubn
j1PUAiIBCYvrzRYop76lz8XhxSAbxcVgKu4kuXjJLB44J2EQoct/DnkJS2RkyieWvfeSwk+s/md4
vksexfltoapIiHqsQHpl5oi0VnWn/OlJBrlVgRnOaDCOZFParuVO5zaHLHOCrdR+rEYvDyfopwFm
LJFOM4c83/eX/MQmhrT1Nt8GbFr5bCPtYQ0xFXnHnxTelks6jB5YlGTi1p+I00dZcbLDgKNlrcec
JPjgkbmNGKYQxSPSZRCpFeecD2EfshTJLxom14xTfHj5q0RnjazWTBJObcC/fN3br+uYEnznC0I3
lDPPDFSuvwCG/Tfgjt4F8HfBlXEDYH/4Az2fsMrBkKMXx9AVdRs3m7SH9NfbR+sb6ele3JS7g0+W
UoW2swTlblDK4d5hDiu/8KfYMpZ1jWp10IkAI7SmERLvKPw2GVAYVWdfUpN9qfjO/lQfl0HZyWgi
Ek6cn5+bkHBWR24yEPO7ikpUPiePvSgYDfZUkRjhPhsQlwB2yhAq4NLMSRJQb3wakNWsz2tGqBRa
pbrm1Io2gEjVeEQ8XcTIwPyZf4YdXxtyaxAOSvKv+zUgNOCEkS/P0hzKlnWHwq0/cocisAB434Ru
XeP87fqhf79wL7Zge6lO3YYNdswc+u5vCwdeS+t8PzVs7+ttAkHF7EoDlmeWESTL7m1BUmaGmFvc
H2eW1gloX9pEm6gIr33wWRClVxE+mu5h1GkU8vw6dSho4Brjo7UIjrvyjQH20BEIBrJO2kudtanD
MTi/34UCRtf4orWU9eHsGIlVckZk9zk580e3GFumBvXjQkk+YqSh2uPFwbqHoaQyZGoH4Fu1PcDD
a22WlikoOAVLy03dvZ6j8TTLFpTKHQOBNmsnA2YK3aEVHqmMnJH3FHzqM5Vd91KYZAt1ZGj7YmIt
heAjRGGlmuVVkZFqpnDGAjqgEF3PM27uMw4WVwaA+5zDa8Rt8rPqpFWWyzTJP5nmDrLKdC0YUe0S
rnxskfDqIjJ2m6Ew0LktbCq66a+eOs8kzozoMQtBnbw+fhZuC4oHOH83S/PJTCBHsKK98cfig+dF
azB28181w5P7tTJave7uh8AVxGKxTxQdyrSxvj4VGvkFEPNuvQtJBbyMwmMD77lhC2Qhko6DbyGo
6EzPoLMhj1DLnMA68pvUPDab39VQc8e8OKpJzBwq5CFT2LpkMuQ6Gur8gtRQdJIrSPjhMoMo/8Gv
rjtJk5T6BYDvElRlcJCH9JhZYD6Q7HgiDONXQc9QyRogiRg9uXNvYNFRytmRydVgFJgyarX7jTy0
zH5/blA9dIAtyImBM0D7xgqbd1Rno87npWy+QgfPlB8HlBmVO1Y+qlH9y6dFHNs3qZlPvKdOjXb+
yIHqWdbObPhKuVbFNlGoa8yWp8rE+E982c13BQT/5r0H/VrRtbhnM0/l4+WDq1baoiNcZXqzcqaK
aFVJ+fC3B87gZyQXofc8n/S4dnOdBtuPyC351Hz4W4Dw+fRQ5EUH7/UiM4CTeiZmIDmoJWGq8fqL
4a5vlzgtUlc3mhHNkVcBf7JV44cXTKTH0J3po76z9gv8t64N4dUub6fmzFo4vfN2KS9PL91eORmP
3Izg3EeSK3qNtLRgiRjwMvnkXXylTJ5VS2QRTzhgcZiwZyQlgANHrSVOE/m5WyuSz7QzcfdiGpqV
JGcJYMTDmr7azwByzYWsUBi/8ht0VBpyet8u3T7XiYTgufsqlAWwLDQqFNr8Vy/MI20OSoxv8x+M
jGrBZt+EzhoxvvIzlTX234wmYBu5GhswP0kh5lu65jVaU+qkGA3ONS0hzBi1XJf8+y0sIeVC2YxV
o++DXsWcYI88ljGETWNvXW/Bq7tnlaBGhA8icS5QHYmqZXWfqKvi/X1mnb0zPs/b99nAusFlObY7
EnD9sO0AWwSCk9tquhlm3svonhqJV/Q26SpCDIEmPkkTsezTbQV/LpZpB4KNXRsCyTXNjA5ofBp6
sRyj5VYAsLDz7BkR7fAaRXOKWymx3ihcyKshLSla1Bmo4J/id5mcU4Nkyk17lROj2IgbtTc2n2BB
oGxU/UY86NsFjcyoDpj8BZTXDaOXfTtDrXQQFXeT0hIcVBQmz44DG+yXrkj3C+T2F7MwKqyvHxbH
ejC/7Y9jn+6rr6yNP8WIE8NXSkZJkOLSAI5pZnWQ1E2+4774iM5++CrswRHG52VP0AjYHmxY5Tkp
j0v8tkDext05t71DBrtAJX+Ok2D7ZK6bH3pkJvPEp54YG75E/T3+F8lMCGWaW/VHZokr6qXleiTR
lBvNgKifXhcPVvkX4mFzajh6Qi9flRmdSjCmeD6xyZmFaFSfvlk4CY2FBgb01v+lwmPxH/eMvSYg
ZzgGlEMQdVOcujQym38IRKNhHvg1ywGRUWOFyCpd8YZWVs93/pQQwdfSRy1za3GsrVwhwXixFnJB
u1eWDOxbGKt/VKDgpk5Mrzk/IRyANMzXg+pE8V1551CwnNo+ebJt2lEVSPbELtd+416PiZBFyRdZ
af+1hkv5HBop2PsxGyCvDDOFxM4dJXMP+SqkbetP8i9XCZvk43VtHiV5S9bFG4XBvGRkZsk8IG9a
UOzBVssEdOMomfWMMIWQS7KxLGVhpehX6JDNjRN0F0ZHVFXDrZeB5I/XjY7ZFJkxOBqTYQLdghoT
pyUlFWiBwnHweuzqipZ6g0ZdhwyPbIUHWTieeHx+MPApaWrVgITThcN2IGDKJb8luRuU6HaAy0O7
bvbh0nBC9337u+/4LvpZVFoDkNxFcJVBy/A6cKjVV+n7mh82GRAghVDb+5B/hYOqD+LbxoxlVMn6
kH4bzRXOr0SeDaDf0Zu2LnGf7dTxBP51j9qxZVOxKf4c3kmpo7VdlAEkuFTNGBIupEYSdw6IzSIu
AOyLuvSDqenVsz7o2PdtuAEbeuTaWFGEdCP75dXJ4syMtFVdS6RR4zkgnaU03/jJL8oKWr1Rs7uj
6Gt9TJPKYCP7XyWl26v1N2dqy3RSAa2jrLJJRafg6wjBpX4d5VyrG0kZ0GlFOvdLfdpqBTwni7CR
a5hpd/U45gDnSRNQgQio0DG2WBV/v8TkIBydtzNsJDjmOKxC7Wev9lDVhtwYesBccxZxRKjjkLBc
rQ5O41sSy+Qn2mBeC55fPvhKYlGAkYbUaqfpJb3K8a3/eo6pVGDlnfBko4itM7oJNYRoAtqdsd8m
pH9hsQh03Gu1s8+lwM0ZBXm00bngcE8TCmCbrkB25sGyxPuhBA6K/wdu5QiGhYn6dawrkGdxlbE4
zeNH+k0M6sDj/WSXEO9KfBs9+snBWdUZfatMJAHHT24+liT8/BRZgc9eCo1R9uy0gBlJmnWPgnb1
izreo2x/RiO6NBuHTnTq06TFfVozktcDUTt00T313q4l6gQiT7t3YTokh7UxP3ZXgcmRBU/VbDz0
I68crN5IbH96q+tRSMSjXbPMLI5abg0sc0V/QbE7UWCMp646MTwYUbipDMlg3ZOiAx1X/qc+3+7h
JbauMOINK7jRRfoM4b2dWsuxVIsfdJlMbBmGBMwqJv/FyVVuky2hNiQpGwI3yy0pL/UBcnlml+4H
oUF9S9temL6OjZWizdZGSjY4YSqeuM8DYYdCGPDFp7rj/ZZj77fvYliplziFLjoSw0OPsQZz/3Qk
9Pt6bTo+B+EAbyul8WOj+tUGW2VHrFoARSirBRslwRLZtGHd8POfmzot2N/wYbO+oxovpbiABtTW
TjnyeNjAQTkrG3/9C23HbTdl4U+WTyj5ApggreFge7klDeUD5+m/5FrMQ84xy2f/7MgkpQjzVQ24
pI1X2avm5BIYldzAJU3IoSzWhJ/2efsQJ4c1UjOonfpkSdOaLnrFw6VnGBFmzroq7YVab5vZKTrx
MX+Z8MsmWb2Zw66dzbSZO5oRX/awO7ItclE/rRaDNVDv5scG311514WrN5yN/BIrfPy9KauZ1uAt
+5JxEF72Xoiaoz7e4MJ3kfZKKV/wJfjpK7myH7LDjSyU3/uxh7Jlkj+BKUabTLN6KWdhJloAxAU8
JJQpQDELxpMiGs6VW57ZVLIluDsjvFmGjOXgYOwDeMNPA5rhZ/YXcibwMsvBtAc7cnF9RpP8LllE
8tcV5fpsDzvGHIAlRsNuAPbxlXcy3Dc2BJWU0dnIqFpG9SWXT0oX2E2Zavgff9noSlQajMgAjmuT
H1OD41biCfQetkiQPFzjImMcccgrh1r4Vc8w5DtbU2Zql0XhwssTCacB7oO0lCkxqQlZzIql0oPF
Zqh7stb/yVLT7dw3KPf53nnZ18qgGGylzETVdNHjv2ZqLqNwJeeBR+px2T5GYEOggewEhHiDEdY/
banhdEHUa3Lrgj/zFx0CiAWF6RW7mmHzZYUQTUzqBmoXOuTXLhfmexZcSpJYRnZ3b91HB3vIWOT+
BuM9UhlwcMEUjyMjt/xLE9zESzIHk3ZSjNxagsmCuA+FDuBmQULdsTuGenAllJJUH7rgd7DrG4JW
EQ/5Ew8c7D7UN1ofNdS3CZGCaU+5Q4H7tiFmDCL/m3Z9w3ZwZBPE0qOYVUGpuRLIsYuLAn/6NDIh
Q2xh6+gt/z4cMspUdEaQmSbwjrOPVtEk36HpE7chTsbGmHzw5pymw88MhULy3hC1eXj9MR15XjDb
ksfX+NHGwtuvN2aKCaBiHF00tEqRVeJBf7MdHAcLq5+/k5D1o40PdDkEFNXSqs97lfxoI6zqvCiZ
7dSUG6/d4cAnroPOimSX1vMP3hy67Mb48zzj/rreKP869F75NhZ6vdXmP8lwMKb0BfekjfSr8Ys0
/TURNhVQsoY8bq2i4pPrrFY8KIjfkKQZcDKNRNaFElV3Dd0tqJZk1X/q8HQAtlfWC5rypzNkyMcK
oBtMfmC6C6IraIc3h1G9bjnkMeY48jYQuKUZ1qqjOxXtCEOamwFTSnUkfztRUXcSp4E8COq3bNy9
0sGzeL9Oc3XOfKLm7iItTJrA78dGM9A2hD6cASPep+0wd/T/iYpvfJH2qbU3beDGVpOkA31+vmUG
lUFoxz2eM85Zw7GjqKtHVegl939DfTCQwlbcwsVoJ7Cb4TLbADvPpcYZ9yfV4qw09AiOLMUPtoVE
dh9fzYWIMEhkhc7MTM1IO1xLJ5i6vFQSR95f94CX8pEaeBPXYXhQWBN2pRvWJSZmAMVQW9tUtFex
2LjDWgbuqA2l55CkCto0BFM96xWRm8fGrt+9ixRSphMKJuc8e+Ib0f3zisNCincaix/Z1QJy2Uww
cELWQECNyzc3F1KHbjLl4SIprkO4oIYeUGyP5tcC4sLXVV7DmN2+ElzrC6exCY+MKpWUi6YfVHm1
s6V5eHlI56OAX4vP61CQjK276kAxeAZmxXgZt3/JUQuRJPoUWi62ITcPM/anu1qRDlU1wNpsHVM6
WJ7BoUGOYKQrFXNj1TcUUM1ro3bngrj9hJk5Dzjpw3CA/T2DQUnRCkcNn7iIwqblkEu/OBJDkXM1
RrEgcFwE4bLi+8Xo83cOHpeDNm+0g1Z1h3PiB41YdiMWeRFDBgOhRaAiU1Bz/RedxTDtnKEZfidm
27DOLH08ikrPegBndusp9mHT3mmPFqC3KE3JSSvq4LfxGzWvfzbCi7AsX6235b6Pv8hHBeMdt6tY
AXxo2sNEREcrcVEmX8MHXkvgmcZE7vvrFM9S3YI0FQgI5PiDA49Lobv5QIq7xEvC08/DS1nu1NF2
U4YKxJLCVO84gS9Uw1hXfL/TedrsZ5Ru9t//hvjkdByydO9zq2aTh/XZCwrVoa/BP0061dDw6t7r
an+lrjrce639qQBZLrLKzJZgwv3YHdbqG953m+wHwrOgsJ9XeM+3KxgOpHyu5ym/9v+3PkvYX38C
ZHHjWhLhQPcv6CuX94QERonPbh1Rwg7k4IUTAQvhCRgVjVUpJ5sdI2yXkrej8bH76ZyfnzU5aD6Y
qnwLJCXHBe2CcF5pYESpWikAY/fSNX6EVZAlS9BIW24EJqntY1y5BhEv1UEecqFjoot+CM0jJNqM
CTBuhv0LgS9P1o3Aysl9KPj69cNsT5zHbQSqdR43QiNvP15PS/5a0LsBNsGX81P4atbDyLrDkRGO
G4i5i3g7iS32Dj2ZAiRhC5Ai+i/ayyiVf73gCMHnoKIUNB6ebwDiX6L1FpOWHxJnhI97G2xftGMv
sW43upRnSMKUFJ07EI9FknV6u2bCPH0JKf0/rM4g5YPPXj5VtejZ6uPXkjFRfEETuT3JpEKhnZwB
Oq816S1ngVvSu3vRQmrckOKWo7o3yPZOpFW/lz+2ybIjmqTEc+vJPkPU95A2e6BRBIfgUOBYyL4s
Q+qzoEBIa7F5+/KbistB2J2EtlOvujpj4YppU/Y18cFLOrNHW2/bL/ymew8GOZEdRwmKyCYVLIyZ
7VWyOLk6Tm/QBVnXeGtbQnU36E4iBiCXnRO4ueesujhtoZrPp8AuOfRRjGyY/hE2CURUTe4DH+u5
TQDx1fRWWz+Dzt1EcqL8s2Q0sRaMlnMPYBxkpVhWCqo/OVBEcMjvwEiwdRAAKiApQ/Yeu1kXIQdi
L5zoqBzmbVRJPco3IvQUJvN7VKVvoBgKe2zHCFowIaWTyAx+Ok6paOHDjrrVlII9h9sCd71tTN7X
Xaz9VagPCwetkcZBaPRNj7NESLE2RQ7LeSWU7ciiJXTWuBfmuFM3eQhHEwhG7HA207nCcUwYG/wW
TjlZai8B0MiMrl5hJ6fH9TbUu7jx9Fi4nqXsmKn0ChU/fMNEgeRc8EAiCcaAVedftY3r4wqRgutC
h+8LGTT+hfuBdvnbb8i0WS+ONazXNsWoqssEsJJFp1bqpgBdz4ljzE20HJtYWPrZQEoykaCAjNB0
TP3udbjMU+66rfnHTQsg/G1/nbV95OmEIywmTCRofYFqC4KWqw6WVY5FN0C3C+LWkgU277i74cP9
Jt0GOjfSFYiKpmmJXc/GjFOkyJ5J+ZRSDuMEWd+1LZDs9lPOUfrxYMAYQFfYoCx0jDkNIrWIlF8g
y0O81Nrp1p3/eKUUBrw+aoe6GpuEfKwJHD5SI5szcMM8s3fQttxhMX9aHiXFQhzfIbA/EmpZbOFz
IWOAqhmkyD1kDjjg7UDqaMcc8ZEMbov47d2cVK8RXhETgoCpB8Ho0Ec1iJwA3zI1Jh/XLzIjKAD0
lFIKA37Rc1UQxbZgI76/3X0S1Yx9zNRkYmNpXFaGvU+zxMs4L1tdwNyLgusP5LAunMv2/cu8HwDO
d1OXtngXxhczKkhijHwGqcxqljD7lHLMzPzs0zxcWI51VKJOh/p+g5e2GI+ZPm+Luyyivg5KVNCn
8cPyq+aFO/IWZvTx/NEm/izyLW30YH2f7jOtvDZGqgElGCndJy1ytTHmxMiCusn8kGTM7jh69nkh
5bIn4kp9/1kGWbkqTJbhirjKJ5W99O/0lhtdy+JTwKshs68Zk2Crfme3yrBS/9I9KDMNukRt+WML
5y1aIlAJ7ja0b/sbEh5+YB+JW8yjdNCkI6C9joczx5ATnFFq/Fq6BLD9S8SSzzoF4Wc/QbxltdOz
A3ghZBmji+YW1YPg0Y01nEOjW1YBFeXooSxoxqBMbIjdlLTc/lRlwYcGq06wzA1GbDfRCXPcBJUK
AC62RgrOULZks2umgXUlI4/uwcL/5KvQFmSwxX33R8aAO6sPNPHba1Ncfwh6hBgl9l4xC7yKglbn
AF0DeUyf5Gg714wwBdH8RfXXbJ5AIA2mwOARymBUAoaQThhBCH13xoK4bM8p8WCBQ+rQT4av0h+t
Iknymt4kPZFTRTGF0RzW9P04Pa4OyzqnS3NwvK3zSbJbkhHfDgw9skId4nYcUKeSDnKCdevJhf7H
MQeCfUfjY2VccxxIQAofYuZaMc7SHn9Ol+UQXKMTqYNhXhRGvmyYLrCuVXPxEdjJFUZbiS1s8/ma
3gq+KRV7ZpokaSrO+eT7+7LUNSS7bOCwe/0SBLfriQSiKW4IGwbd4rRvRdT2hO81TOMpHoqsnPMo
c+eB/HzSVKiRCuopTk862K7SHKVWt4kvEs5ydtgrhD49GrIBa0yoWvpkjiKHM6peilMMNyE6xV8q
cVwkpsdRb45fuZTFWKa0wxNOFlgafvS9XQLhV/zulz95uCeDxO0NXeg/EdU93uFXNgOrySPlnpH4
Ws2u1tZUsfkmG8bHBHvqErC/lHs08BTzNSFjmAPKd61sAhs2gHxkVFD0ku1Bu29qJhDuJPaQ56+3
G471wXBPWLrsowzfbFKt2gWg2gIpvqm0+Yqp2mRgljiSGqCGiga72v5pmexQt451+0m8A2xbZ69Y
4SLonFGvhQSnAt50tTq+Xjt58tYVF7m2Zai9YdCSo9t5/1JAOXATHrMMJVIvJ0ZZyoof0wQhI1vS
VLKV5KxpZBQ9cLWpplpGO1GN4BZw4HDH0oa9WqfopZSg1wcOZlOkP47ln/CQEs8x1u9zEjT00Y+s
KSXPizWOqm7sFrf2ZXwFYVW/RtPx5BoWN6BxrXVywDPjzxmpLISXh0MTbyxnZ5/UulXqiRYsfBhc
f6YZ9bN5rX8a7/Cv2/QoTDM5hB3/wF00KYahF67sxRcWExcE0+wP4+I+WjhJ7b1nbO97lKWGrZHD
ALJqVOqcXD86MadFTWU7izA/F9vSihD3aghG0EhDMgE8vdr/q8DVKb/64XYhTyRSLj6DF/SQ9cvL
wPKOnVYGMOQXgMQ8MdotuFw56uCB601kwyxr/AgBXmWNwIJDLGA4K99ejdwbmuFNmRPU5cvOUQWY
ZYKlcG4OHS5dBIGdqIxyXJmGP5LrEN4TUzRwY8hjN1365dOFVJ/vl3WFR2zbenib9gqa6xCoOE7h
Om/kp1ENuaWDlw42Mc5p12xMVKRm0Q9moLIEJ5Z0y3sVnLs5AEMW5PjtkJi4LOuoyriF24wH9qfH
I/uiw9Zdwz16k4EdRxtGYaSmI1OR6NXcDbdNji4cUpzgH5hOhk7ONXg5SqvJJ5ISrHr9c4XI2gx2
gMvkq06zrcLHen3xg1HyitwzzIOyVsJ1id4JCjrswn3zbe2oXFkaYAcL1Z5+5AQMTkixqQXCXShO
2C0/aA1WoVF+aSrzUHCPrA831cPTra7Uwx67y7DEJhxYZP+kWoHlunRIkf32kajScZAEgxU2NdOo
46pIuIHfNAnkX/FUrWt+YpZwNi0hm4VoVErq30DJRzYwBeblx+6XeqyPlNPGU1LT9b7OG8+0C0o2
7wIBwtr8kzNc9t1I4x+hkiQaSShekRVIuLZfF/sli5ZmBcVqmc3JTcQTe4LAtRodD7TCrYVrwLMW
14Iev5hPDrh2yHrB+NjHpEj2I+SsYRCQbWF7IYr/VzpW8ahFyE5k9wyoKXPDH2G9A3trF6B9dp2e
rAcaC5UbuQZsgxSxWWxC7EmJq2ZJPZAe990RCnpADViUKrMhwwRngPaoQJz+lonmRKo6BjXQ3m4I
na24RMGKFdKTtfeBLZcEfCpGHN0S4TEDDp5rfYotEDIXLPvE67ZE5S0NKu9GdZebYyFYS+IHQ+E/
jwO6fJKCZcHXCgFGWA+udsn3clqIACuZYJfViGe8H8SU3JEGDVc73ec5iPG0iJrPC39X32w6cbzB
K9UUp6ifX//jFgPS0o8ZFVRDdRl0gxtSA3widIrm6Ph2kIuQCXPy1yaVQO2XJfGrqVBS0Uve7y+o
k5zu8QZY7+XiWAA2jVofQsB3dkskCyb5+lq0LOf8SXdab2D6UYyr+btZknNYUkIHMdxONiJHiF/c
8Wt9kVSVc6LguOzGwK9DH/kLxHY8Yf00KB+15XtdJP/SNR78DANtxmvMJfVOA0itMaxyHXl3Lw+M
m2mQgEzC9nC5hIZ+N/3NMvGxt13K9LCerP+468x01BCd7bnGr2nT1P8iJryT9kvQAIT6vvRsRjZd
SAQeuTrKhx5m7fJIFstC+7R0wd3HVAddRvXDpPpX4gTaGvClHGycF/jBmIPlqPyjtusRoUFVpwqP
l7J1RfNZt7FnEy7A4juP9PD7m5B3YPKDZU9JQ/Wn6TOKPpXBYFPAc+BDepqaB49VugXgvd9AyuJm
7Gf08c3lgVNUkxs65QH+McGRvfaRJtnyCJ2NffUI4ne4I38Ai7VNrvui4KbmOgKLL7bsUzSxqc/m
jrcOd2SQ/asADEp+jgRMTCe4Vp1dxl94VlSijMl18mAGgZhWbfFxIhixNnPNrL+k6HMcOJSmUYGt
nhksuTis7vLAvTxyqDJOL+ckqL/6nrI6WmeHBcyE6UX2I9Zh3OPzjXyKELS91m95NvQRP5TvIdyZ
MdHyiknVRuqEhVPXKk8jApg39a5v0piKYK4oD+1ms8hfq4QDaAGHt2lGCpbLl44qAh7LsntT9CMI
SN3WkQzmtSSCtiXDNUDhCdUMYF3+OcXj6LPoxlRAlmi+n06VaTO+zVqOBZKcQ1+TwmBNKlKj1Tj6
nrAj7LzlkVCiE3TtTkp43qJcB4eiwzwsDFQYSgARifnyrxn0KCDTV2AOR4WW5EJqvF4CBzd46izE
KyflUXmVU9+s5h40wyKib/PxVBpgf8ElD+uKPRy4dDDGK3npnpnqk5rgF5LoY0xaN76oNq3hXM9q
JkGWdpeojJbxX8xJOs0YhVc/k3x//PEHP5OaBZnd9M7mwpfmKOCfSlKe4vWliMGnD6MGdvX/oq3K
onjMCp9soLqJvvjTYwfuUOkUvM20cW3nbiO9WYtXrYRLQXMX5eyJjnGaAu456BZUK2obSXvaZdqi
okFsf/dHM157tBZEtnWMlfTSYYyEEv50ghTdd7uTIB5hm0gjb4rrGHWRTnGpuQWH4CqRyeyN06lC
LCBW0Jsw52lXJ8XJFdOT0W1hVQojz5WqYRhJKepOe7wXVS3YF5SjeudgZjCQw7Bxw6gIR3TTdU4K
DDjktwCcSPJf9+4hiBOy+GwTtA5HMPNwRolzEVXBZzhHUp9Xk8DXeVBnO6i8TWux3sUaGew9UFJz
WTLsvoLTDdbQVNN4ABiv+UHVwhpHW6AkcdT4M7TiuuYRcIUDc7taWqzzV0Z4jHSwbG5O96ghtBNB
1QgWwcOjTyPxgiWtqIhcGNqGmTkD13uv6X7/7lHIKiAnCKPxYkn3V7mPFFf19c7zQBJ+mtpOlVj8
Mja29PuAjMkEVmUA6YXV4qJy67UI5Nh5kKv/KtmFCcBlnpKphM/tkyT5NmlUBMfMn9v37icabodv
XRXh4VZqnV/gzOnoMhsNgznkZm3DQzIfAWLN9uE+fC/kk4Xej7JrnN9a6G78tkKVeP0tcYD28/V/
opKRxY1hAic1HyjxwEX8nHE+ag7KDQtpN1myb87fnKXukvyDJovEJwbY94ZncH4GS6BRIOt7csGR
KbWKg4yPIjmoA83bI2qcVfnwWZPn136weSSa6cn5u8xPW8Motg0J/fS3Wz7zZbmX2TtsAwPa+Qrd
rGjUCoFoBtLicm6WZTLOs98qviKhqeu/wY4nj/tp2/alafxuph9TfgOUIt946jHDwpEixQ9+Y862
eTesDBF0NEZsQpfiXHfDJLS2tecD2Nd1O6rln7tgtHNPvuU+ts6xkS12MiWHopfqwITD7kY29rYZ
jF4bSCxa6zQXiVa1lLamIXrsZO63QlyCn7GylqXIme3ZA+J6chUCBi13Kz9hTPQ6jGHvWno0ClbD
+2/qnhppjU3/+qrnW6r7pmPD5PnWigio+l/5FuMPahFl+mZiVJqoBoCUizLeHhiI5KicE6RCJQyJ
qTGEmU40X/iNFTSwCKXvomx7r1DaUeFYG0VbY+ObLA5oj6mdufwBca/+heFy/zT/FpND5EyUqdIs
MLZg3wDmv0FFhlZuYKh2LQd9tqRKUuVjd3ig7sHttD2V+ant9UQte3oU0DnbpeHHhRhjh/exFhUT
DyJ637aAKqWXOZG8XszE0ajO8E3NUFcokMCi0xFnjD9tOyWpQxtJgeLGZuON77q2yGlexrOo1AJE
8icX/6Q8+oiS0zQ8VuJzDRVuMmuMD1wR5IjXXAU2vWupiyjLF84UUQ8TajA5DZ6wF0rdiAp+Iie4
KQtzLK2Me7GmfYbg33HWDcJNcqTfOn4VuUcUzHJAXijaI5cNei8qrKjusRiQ9y0EwbDkSR2Y030I
MVPgBKjtth/8fIGUj8Ew/1Df2yIF3BMzsRUnO/STu9jXtYZcp1LvXOrVYeuWNNZn46QWM+kUANAi
b+Yzm1A1wkWgblyW1A5aNgFMW/k+DlcEiUgUo4Z6s4nW0qGw/EWFzgnOYx6p1Zoac+qTZ8Mank+e
yG//8pSo//QNx0IPn77yt/2ydrqzgssqbtC+W8+3pSyeC7lKpwJaSVNMATimquVx4wG6Z15Zjr4o
dncIJHCItMArQUYT0VMRjV7nSFRkWk2hsBuDQdP2tj4+3ywZXjAAOurmd8GcoF1a5x2Fhqp16AZL
2h+wZ6PoMFlBdVjQkJVBUSUO7cCRYa1dfVPSZaBtwgfj2wu1mSDTGFtVGf7m4Hkl8/xf6M03I5Oo
dGQNQyPcVUVhCavc6TdTIpBExVxV2HMqQIdQfVC//txMHrVp8loW9cSWjkIKyeiROZyfS7vOQewr
R9sqQHaVvaxRd1IMg3L6eRoWl7KCsrAtsDm4ouoGOJhGkwA+NTeavN2itcAxPkYNssQGgqICTf5G
FdrRw86PDFA5aAqS20ZKncbTe5RttQjLcUvy/57JvWbME+cWX2hjm5sdv9QSyYkb69cBa3IJhPdy
me+hdztbH90GR7sHA6b7YPoHnMRmlq9oBisRoUBOcDrsQh0v4crjbNDjHnzwikHdcvBlpW4G029S
B0SsiRl9V9pcxSW1Bza7cgkECiV2iL0R18qxEdEtsID6Wrf8pB/Pk10eczusZlHVJyV8ijsc2srw
ojDEm+EisQvGxQ+DBCeoqb/IUQV6fxXKxjJY2JFpUEOTnxZLx6B/Y4v2vJk0E5QuJQpvZxJR99HZ
90L7n/McFRyQDU6lNf7BBM54Hq9V9QOZUbBzWYrwctD50NzQl9IDwbiMY5vy8R+wBHvI4NnjFFgj
LMvMWO9+ZEhjQsFotHHnUYmhEBycCU3MF6M29xHvOEdHH5z0yrITForWfPxaCswbxFY+LnYgUky3
ZHHlAJj0vzpRqAfQQ1fp+uT1KdDWHKXHTOqX7zD2stOp2YTOOlF4kRqzR4Y406ldl7MVwnujCXu7
FL/1ldoOUBPHbEM/T7ucJeTSf6iCVZfhJEIgVKZsqizVThlXQsRWw0+3N6cyUzDCt2TOKMcY34MV
uIFuqReJYVFAz14X1y9eQFH2N24eII55waxjryqePWBX+jH0MyZ9NP9lkXbno2UYCuartKSuKdfR
5EHS0Tq0mFZ6rq9V5hKZNFkzoC9Z0FtE7SLsNUW741qCj+xkRN5oInVTARIYByXJF7SInvEkuylR
q5YxgMmBCdTZEvi9wDdUy9vT3jpqTIqd5RBChmw+0plLD1kd9oo0lDOL1uYGUx4JqzpwSDykzYDK
2sj0s3eW9McOmTEijVsmxENRxe9FFlv3J4Rj+6hAsLVjeeviTyjpdhYiR4u9zrzJXS73HydI0Go2
HoJU0m596cfDk2ag+Fnr8h0jZFHSA52TvzGIsmA7eXJenMkuzd+RCm0YQkRX3msSs6bDOyxSVzEF
c96gy1HzToLabBnqqm7ZTei2u3XHonOW5Y3TK63mUWfCJXGbR/WPBq3As2I7oyxwKQKsc8bFAHkf
Oe3WRvgEHm/wdtqkY4ZMAS3IlwbWC713nK92FXOl80hOKb49m4kpG8VOAQaqcb3tXOs3T7/85u9u
79wCATarb50ImZHZF4xbSOSIa++wRfKF3BeyOtuPp9dSCZaM/RYwD2r/sj2NgnDlUgd/ciqisTe5
yXZeQ4IMV0G6ud+TlBbSezoh1WMObDaKG0GsjGIlfP/IWeq40cuV+sDiVKyMC6ZLIwhjtEs3KaBy
70IL+OyHNC6jLnCuzDHZvXBEZ+DeyPATSp6E8ztHojv4Xn2lcFxYisI62m/Qn1cUMJoCCABzvGLa
i3CQaeOLwCTiV47PaIlI8r53hZhMsFUhhSxIyPJp1BpZrmJXZUdalQBUn2PENq5pqI/didcF9RKg
s9syW3ZIluy8TMboz9ixitJj1Tn7mqRXR8jnfCGZRl6djy3ygEKMsyxj6UCMHzse8uSD8eiWbNnH
BKbrL09AU1NZUwn8Nk+uYc+1MKRUw59jigNmPP7JUy1GYfl84YHJcDxTwGDUaJ1t/YkX4ILDRfz7
OoHOEt3Q79JVulFKs1O9/PIaPtb6DKGZAjDPQtkaOS/hiaxFWQ7LA2i9H5YUIBvQNhTT4NVPwyJl
ToZDxmrvGYoUB7vH+M0pNjs/SUh9iXTWhEUEg0Cv2peqJjsZkc4xT5tqNmAgdOeLeZKJHmiGA8qB
VK7MBgua/LHcpJoQ7BgaoIqe0kxVOpp6B4xCi1lIv7iBIp6ZHj41Qg+sce6aklAkQ9IWrBo9ksJ4
qQ0SmQqz9zsiG5FeRxs1whnG5gNxklT7gEuwQbKVC2daUlF91dQK4wMLBX/Zj//xCtJvzM6PsWkF
yAgwTDAV7X1Pukl0JOncIp6/iFgCmQVROKA2B/soSIquT2E01NvU1+Y+FAd8HmWiiTuoUGk3QMVL
xB/E3vYloSXuawdK43VmzTOQMk1Azfh6+I3A4VtjkDRR21Lchut5nzIAJv356QTOWB9CM+ks8hLk
72MSwsYdjZNcsuRCpHtv0wcd9/knrMOD8XkNUkpAUrdbrZsZCi76DCm+ritVLRD0dvdIH5TrAEKv
xlIqt59uIXOllmIBgiKK9hp9K8qo+NpyDc8rONyNfk03aP4ol3P/Rs+sCmGICNdoXgqwwKq4hjdx
9LaWPKkOJOrn9xc9UJTU9CK/s4yAr8ecOAfF1KeTrRFIneGOfCk/2agEfPJ2Bys4d+e9AhjHNQM+
+tImUgfS62/1K4UxDW9GJlWP7fqXRC0WkZ2hi4hprrkdzt7wxIlXff7c2ILtPQVGDI7tfkeQpMig
LidmEzPexeKK3gGuyxtAMjWS3V6EbW73fYAY9zujZIrR84OohbUMMd08jAuDLDqP5y1JhOrszPLY
HkH51xyluzfwhs6TDhTo3u5iWco9AoZEnIUljluzN03Fso7MMOc4MLr2pN8coT8ZLF9ryw8RHEvp
bdIIMb6Z3uWcSpqGw8m7eiqML1knGvCLK4hm7Frt8y1wCktsukQOxRxC496LGZ0U3sXp4w68Tc/G
hz5lAcs3s4tnPViRCGjrp935Q2a4WUiF9t25ZWb/7WZ1sudJSiec8jH0ZmPggHwuTvnrnPztzvYw
aVbtoztn8Gj9c1L0bLBDg1Ur6pd5R7u4h+osjuc15ojfZZ2NwbfYZOOYOvibXPq3OS5osN/fKpji
a6bZcfOR1V08pxwpi0rfqi/mqc42sdg6Fzb0ZGlY/0DhfI9tjmJ/7HgjYLZW58wSQKFpZRUB8Df3
UFh6xIFw5xzDeVNqCS++4fBtPFgmFonG4pCGXai+lpIWhNUbu7eQH+coisHJM/5Qpe2DnO5A7LCH
h4udph5fjLsPnxZsLnzjtYlOrLz8jgK6rCzxPky7lwv9f28O3gb78ovRHTM4yM9LhHOmxZnzdtcE
i9P79it43LIO2kL0VNQCNs/IqJ7ugMJz6Ghl2S9MuOUItvsbu0mj60WgbwYmjEZFWjtSoq0i04Xr
kumigms+0uenxaAzKmlalSDQjtXjYph9o4QWUF7bfkibOsfUtsXeik1McE9sfG1btGmYyrpXtJi3
jPYAAoVLs7ONEv1h1l8IxmPPV6WlPQHpOb7hRiQoVk9KRn7PuQMj70YkWKa8684KbaVW0PJeNfsb
j7/7LpwVK+a4YQhFl2TaUZYCszVPTMzCUHNAlkgKp4TABR+TIvVbMsABg349K1JbV/DnNJqQpfql
1NylDB/A1MOR2Yr0egik14GLVuBo5PVR8z2bX8g37inDBwshZpneHMNQ03Ebz5Is3Dqa6NvePYMA
qCIuNuK5xhPTJtG32MOldOmYefHUVmXFPWmGqJW+hl/QQnTtGKc2y9Dxgcf1t18OmyT9h8DekAa7
rg7ujuUAo9Vst6NLLLQDB4St/8uH8AiIusvFhIHQjASZb6Se5R1YMf6pds9h2lFr3bb+eriECdvy
70BEaXa6Uigom3JRLGw2oCU26vE/JxYcOwq11w+33iAo08KAYoeMYcINxSnwYtJ+G6RRZW/ztObg
LNA5e/Y/4uByktWFoas8725J+zPuhYUQa0jvd5RDUF7pV8/5VEXP33vcdgDx25mdVv9dwtRDyU0m
zgtZXh90Yvem31eCXrOykHVUzORbQT8sH+n/CUV3rij45tZR5VzTJ2UKoKI84DBYpz2Cu4kzHe1S
TXVJdD1noQMsBpA0MjDMZ0j2LJpegrRKdKLBHccxy96Y0d1qjL61JVgbiEA8hzieF9InQi7jX+Uh
iynUrjdYc9S1L620FHEu0GSETVLCs485eXHwvRgUNbngMHsHvVE02/jeLMuJO4Fn6z+7FFds0zT8
oHM4kLDx2Qmn3AFVfOM/AEExNtpeKUWSmPaTAGzJmwmSRKUibHUA14Szlv8V5aAw0oG2rwfcSLFn
/zMgEO4d3HlNgbebWpJGbifkTVnOs6VupRlQU+V/jP+9nWX8vBoXQZ0/sbB8TrtjHVTRcNhe8xFL
rVkMSxEaXlZ+bsd9JRg9JCB3f1UhrjaDFVcSeXFBSDNKcm72+1yKxIq+Ecxu1TCUTk4GiObOGx3l
tg8RXJsbmcadXdvSqLjutcB0DTBnZ7KJ64AAtJ8fBlSVgD9S2pY8Z+lJ7QM2IOXkN3B+E3IF+0Ej
zCBAjvKtfDQX8lt2j88/jcvbgxI0q+HETe8D+HyKWByCK4+EYxBfOEXR1Zb7L79qgcvdIu8vIXjq
TIcC7NzC45ZDl8Y+GQAXkrPgW4AL9QaIqIxRfmtY2t2H2t642EBc/f4qJggDpcK4Y/eoORc0lRjQ
xTPc2kavCfPc5sjNPuPqmd1nQMCaPLE1YgDpUCcHGP2tpJkVBpMRw6sie6JTJ37/4jPLn1mytSNC
6u+GdBPCJoMPjEWBo+ISu8bdJ7VXgCAoFlNdVMV12xOIKpezHV1c+/Zyg8UJ7kZ5nfEllX9P9JR9
FNaepBJitMQHXbgNl2maeye54QRwKvLPZlUSEZc5w3L9N5qe8H5Hg07w4aBbktvIV7AYG4R4o958
vumK5wkAaLgY6eQQxn6NF+GxVbg3tXOxFLbcuDMjfwmqWUsT2slaG2nME8rknHyKwEj2gsVU7+dK
PV0lmCSDtaeh64S+WTaEW0lY4tBwasEzSugTxRpx2SkVN+wYazXB0INoOteyNfup2Vu3YB3E/qQR
wC5RjUHwYmoHbsnrB2TFprX4r1g5r7y+h9R1pPZKOM7iM+l1fmVT2DQEM/5m643bm5WeLZvdXIo3
8i8gmz1cfUP8smoybNsDTQnHgs74acB5TQZJvGnYxiJJyt5cagXtYCQ8ejxv/IT6X+3YH/nJ7rSX
rm8cs1SIlO3b3r1Jem4hkC5wPO30s8JM8Ng+Szw+brLEPXRvgtoANe9qjdlYZRw/UE/VlWpZL+3P
6TiMXg/uC8coYKFdiepCK35ZCaA9LLwrupOxjOWG/DsVybuPacZq4YLAQFRBKHjP6EDX+6ig4Qti
KpF/PB7SOGBBX0QSaq6iLmNV+UIfWnZADySd84RZYCxndICNXEA9FzFlmLEUqAA8Hon/ZcVDNk5F
+Q8DQ1LIWbUQBa937nEb4N6UQi9k2aREm/YbXM+qFMSP8XSR0YM7pVdRebFk9g/eAtVQokaAbWl4
yUk2aRovnJTyrKtVnMBK4n5EjQzt9Rp9wMjOmXCKJZ4DD7tRGjr928uOw4ggx6/t/me6JPSyw+Dn
HoGi+4V6Yx+IaOe3n9ZEKUMv+SNLWWcfwmTddsiCma1epsrN1mJjUW+coJSUBnEH+RjL+UZh9VMT
aQSBiFRxaMWsy8VnnG60UJTzppf0DDPHedyzn1P+4Dz9YYbAX941ZF0BqUsFiu9Tl9hPED5Kaw8S
mIecK700opCZmIKvEDYCXwMGyXI3Sg58qIe+5YBS4PQPR/2Lgf/ajWnTh+yoRD7kkB+VlCwVkDZT
1OXBI/WgpX8OrM2j7IJWPyFnP8HY72w/w9xdurAPpQal4i45dHpvDL5ANTE5b/3KAGliQIrnaDkt
UvR3Mh4tOOMmzFvehuiSWNpPtAwwUZS2oB4x4sV5at2pQxVLXE5Q+MrlvZdborq6yDjgi4YDFZI9
+kb8FSnE6I9FU03hT7rX88lF5X75zmo1mH7htOf0oDkJyb5feieiTBcXqd8J/xUzSc594pR+Ps14
XeUpwqsvpbVhpZRxtLXB9RnEfKxW/kfzjM7oL5r5c9s9QT0v30Fx5EF/qhl73go9ypSLwZXW6KUX
36N92+E8qv/TXyd4fEvfzRv5S/UqVOfTi7nGDheyn0WbEmLRRX2ikj/OrOpwb5OhW50q1HlUlcHB
NpJ1SBIJlT/maph6DX9lQmXAIXKoswf8KiB/uYDQLHHXEBRC0Y09FZPORQ7OpP2Wc3JL30W82B0Y
wIJGdz4YMpMDN8Zmj/UqerSGMGckzPXXqpSSag7EIOWsJY5PEeRQBXE4qhJwvuaZGNAYBBUPFupQ
cEJwt84Ywg5UbXvFpsVUt+iQtrbw3u8tn3Q5NKXNgBfWYQA7jX2dkWvjlNsQ4HNOLdy8+/u0Pj7b
4VK6TtcA+hfC+aOypyV59mAxAbUa4n07RQl/th/TkGHLFcGtDEfi8W4/V/cyLTGkZhNHLyUXQFeb
8/eCh5vA9yTFqqbfMp6q1IiRM/TwVhbbNk8KFHIU3eO6otdA5pF6DSCqd+cV7JA1a3BR4BIxj79C
QhBY7TDmeqZrI4G81kMm4ufxXF6NJMqCw29b780ka1Q6i0TIqw4cHrjVmEeOKMoCRM+2+Y89Liri
JluIWpLk+WtLVeMmyRmAyINxCfG9CQMfobhuc6qK8/Z5d6Rz87Ha2ZamI9vz1voYAjiIVJ+pn8Re
Kwm18YjXt2imbrkAnU/X6QCSXULF8ItATQbvHoyJHkR7GmoicZucNr45ZZ+q7jmk4BzpVnd2u3RW
TPp/6f1oLtxcrqxM987AL4s85b0vqtcP71no5Rsd2JK5q5/h0ol+T8K+mTpfL2kOBZ/Iuy/8Sby8
patnJJ9eXe68Zy4Pukt7w4mD6+qQjyioq66K5PEhHlBR4LNfdl2zMOzkmIwMEXeF2IrqfVzM9wVv
myQOLnk7DzMB06L8rBa/YDJZt3CdRHS/xJXwn+Ij4gpjJh+ivu5cMVLxF5YZQoW6xsp8PFLuOCMh
SOVPS86zf2XG290/XWYPgUF7pLEEIlhlGgDB2O5oyWALU05V82EPi4/QY49a7BdPe15w3r9is1Ra
lz5o2r0eEouTN9/pUgo4kMiTFYUZ453rHdmtRvW+wS3kf8h2AwAgeT3Uk+nx960O2WEBsYFe+GZl
kFKeHiJ26D+8T4VDitvgscTRW+if9cBtPjD5jN2L3aNcn3/gowTGbW0YQHLxXvViFdUbm3b1mca2
n5ZAhmV4AInVgnQ+BK6yMvbAh485Ais93AvBHnalc3sNJ27/JcHRlwBRJUheoej730gN4aoIRPZn
A2PxJ5BorrEyWjalClIbc0qUDEixYzb10+04TjvR2ojEHiBfgcmTilxJsbXY/pBVPkyBmS66Jp0M
PUc+l4e8tDmOHGbIgONR3WOP81rQe78OoWDQipppQ9qxMwUWSzQS1VlOqjxW3Er3Ao01HWuaD1k6
KqFpE+QcI7v+ksMPBfeJbPtDN3nvvvINdhDwnTArwGwFlRvfQT6u6vNEaSLFc+UQ41y+MrwxYHDl
ZwrAMabOF69eyf7HbpLzTQohJpKr/yFGUm9J4ZiQhc0tQe1jCN87w+WmbD31jZ/5Gif3iDQDXiwc
SS8St/XLW9anXnDaiMk8fOmMnB9KKTZZ5TgHByteHKaZmEdJi2MF6MepQt6++t61K/4+EN9ZYIeV
4m4oWCKvsTUf5ar+LaiUxdW9ScMiuXe18vqJYj0E+9QzIeUbRrHzvlkvoSluLlWvZXtqIhQBT0/6
OU0kaS/J3HMjgCWCgrMMvDWRS2oSrdcm3klLvY3N6ju/Z45Cgu9AEpHF+jJe0vR7n9IZVZ61n9J7
nsjYfdctnfJvqApZuG9Mls9ioFgqCn/E3jp7rBVIeFedwVJSrNPG/sT1epfoVRmDyDLaqHf7rfSY
Y/k0+o5yvR0mQcwATtE7Igcd1wVTgNPx9eUHY/qnFeQpLGft0COR+ESQbzVjY4dWlL+RpxwmTAM+
kdze27Ao4RUT05b32Mt5xP7hMguwGIC7+YF1INlZCYSJsfqg4T2igQ2rHFq9pmp9zv1eo3IimVIj
qUEyEFEJW4/iTfHt38Cmz2/lkqNuE3QpUpVxGR57T2lSXa+b7+UFJEy68AxCS1ZBhedwv3VlRvP0
jdqIQvFjKrDhKfLPENNxdYQ3qB0DE557TR8gYXvIdKfqxtqt5W575uzuyCbcpaJ1EF+cPVs8WgRJ
AIj4gDfIMYGFxmPY4Cr72j0oQ4upkdmdeln2YppWBiAwliiMxI7cb7VDJN/1bh0Intf/BM+72uDs
bEsxpQgDEnfEt4Z03RnJdxAr5w6jo2xd76mmk90Zk/K0ZJ+gSUJ++6bQ2YGkoS3QxYwdl23NklDw
9HO8bj1wMtSlKCMAq2qWkltlq01VmI/Gb1i4nkAlFzX48Z5g5nnuhS3pqf6HIdgrpOqiLXY2eidN
dPbJ58spmOO0ZPSUbBiUIpa0Wae+ncJvDRvYpIuqJwqaiiKUtLYXYDDpgDbm+D4NmWhjaVmRFc3d
LaVJjH9lYMP+e/nvvced93KRT7cE59bQsn3/O/0qG8J/ybVv60AaUwrVc2+4/kgFQtpoNYgLVvls
wO5N7nxmFYmmhRZdLxbNNrVrX/alIx3zlJDNdBXTPhnSD9t4C9vy7ptVd1ckgV4xo5AzqA+n3bA7
LhOH8/Z+BpaSikugBpo5C+K35Wtf7cugv16A7IUD+NHj3Ls/3zXPsjH0POgSGzYs0o0YhkJo/JWh
i5xWpgcg0hWXKK/fIJkaDf5yQoVbgSuOwGy/x5lBBAF8IiPJP8C162TYnFP3ZOWp2vyx1q2lXAH3
gJ/uHjrfJcdz9QTTm7dEmcwvZTbG5aWxf6K64MJlMh13A18FBhnzs7ReNta1Ya6GfhWzeAznCd1k
BDcBKIaKu/Vzz9VfpW+lV1yRIL/faB/65snwu/HpTcGQHRW6JnbBoOLSf8lRqIYvAd6Fm6oIa7uE
O4pdbtRcT+sIcb9XlSTzGZFSCfV22N3sxOtAz5pALsurTGkktXK007VqYaLcrEDvW65VSX2VOtVM
ctcV5BeIMi/z0g6dBlAHU7RK50Mbqw9gmJGbdqBMKgp6Y6w2Fq9777iod+5kqMQtJGQ31Hp06ISD
je5s3sU8TDICFFJM5vdWeE8hiO8ZoZeWP0xHPtpTz3tDzDs0XkiN95Y84nBwHcHxFpgMrDJ2cH6b
zkSNJNm/WMieKjzbKen0nn9KVSagjLKvc4USE+wPjRNWMYyad1ZODhjMeCtayM1NBId5yfWSH13l
LQm+OvUvisdMsv2B33XDMxBNL+zFo6HJuQ4tvju9PackOMBgEWdroomQ8Wh4qldi3w7ihEfFFUq5
bvksJV86OYGOs6/agPosdSxu14Tfxt6eV9Y76GRQVq7WgU15E2NItldLEAKaEEMdAXlKREc1p+Ex
CKgnBFw8M151G7OHrpY7Ab0AcxrFBwnIKLTT422iWAfcITtyjonAg5ivFWuxyVB+IxrJZru7qq52
aklG8BtARrN8yRHG6w4ahXVBnjXGQF2d2X2ofEgnuChlKi3quC+8n+Gp1c54oQk00gUPlxCiN+pb
VeeFalHUu97fhySMUUp3eIuGI7pMCY6DcLrc20dypjPxZsWb740tFEb73t4cboKGCpNvlMUev3Ip
p38TarDPtwa2S3HNYvBK0jUKzovH1M9mVv/ZkIVvTiSRpxf9rs/e3aXIC63/uTVT6uEO8/G1A/NN
CCxZGSYPJ9ci78lNs87HLWSPDlq43/ik3Au+8kwr0i6wAhu/cbD0cJ73KC380BvHTYWNqy8xti4Y
MNYQwZdUncsg3Nnv4RyTNIQA+CzRVj+SEx6srI9Zd+DNQ8tZ3oLQZrdKlFxU4QKq9QWRfqgGGEzM
IpfNsinGYLeAjATsFoZMEZqOJ8r3zk0a2XQfrv7gMMw01RvnpWxB+r7S7lSsNDv1dwn4Odeq2StX
fVGNt7WTUu8WR8xMOYKWvAHgeQvBgSdd3zvI1+xsH17QvHkTEE9d7A4wb72+XxRQ83fqHJQrrkNo
N0XmjsfNSWGY4N8DGVXYLhwgxslgxkYQubX6fi3B8xBTtrQg8mr1q0udmbBHhZ1Vl+z7Tnvd1vse
6aogJJajvgH/fcPHHCRyOnwaq47BQ1TbZvHf/CzedcXELPEfQqS0bdRd+eGjXTQfeaDgvLt++I93
KcarNaw9NBj50IOn15Fl+1NGs5XkDhSkZC5Gw33IevsaP0b6pQfSxgZ1NPdVFS5qcGjwwrc3czG3
iWGLE+yu4CH+BAbDcZTKwB7G0QLM5oespqo41cdlywekRGpcboikAD3b2VpH/DuEBogKnyl5k4fe
rLKT5f6huhltK5T4ovbd5kS+ahxoNnYlaVbQfgQ7eEurbjQmszAT+SZJvCHebWQXwe6qIK2r4cOz
u/klcCakGGw/YTpTt4zU02IAY6llrhCg5CaK7YerQTjEtqKXTSEUAxabk6xix/Ek1Tx93WfBJ3rB
jDqKhEJu1e3XlOt+E1NOvh8DwC4neOz3YG3jZf8yc76nJ0AtmjgmHQhpd7d3iavB25FBZ/cPQSuH
/bHRgJ9sLA8xAq36TI/Zn5Gvjq0B8gdC3gl412NYaCDSj/Chlxxtm1TlzNBt+uDXeCdO9q38mQr2
YTVTR02aslamUXYAYwSI2wt5W8aIL/wnnJB0g9T5wqmPbLhj3GS8u0ap++80CRT2KPErW2Vtf//S
K4JV7dJEwVErDkydjmUKeDRI+Gl3oYtFg7KxsJSR14lmA5BzHbIbnU1GwOU21zy4P8GOML7DdZTm
l+HiVrkcO0w9TKlLK38E3A0pVucCy5P+nsveT09nwGqOyZtp7YHKO/2+y4kusKaz8w8tRs2bEDnG
f692h6chBtWEyd1GpLlxMSsFCfTZLyUaQnTRij24xIlcSS9KduJLQ1OlzizYCY0QQTxYAyzpGcgP
p+REHDoegO+k161i3wp17whLf5B/x3VPKk0nL1dnutNZV5yI09LLlok9ZPliu9lKs2opDYSdaXBE
tHkAiJtYhexxXL3nCSVo/PYseYabk5YrMoe5nPa2P0Zxl134dJb0hVQbyv6JwauMkdGKArluOcRj
i95ad8limON4ZRFLXQ3H9v8Sx7BvaPboIHYJS+F0qGyfUb07BcerGGBzh22YOnDZ9nX3b86nO98Z
sWOF2K9U6hdB14ZcqCvC+1DsADRqz0VwfDnKg5n0544Tnxfg1mLe1g2jqOYQqy50MyDD2+pf5cTl
s64GgrsLYAoXmva4gH8ZWGl4owASO0ixe+I33WHlyv/91waqR2ogh74y0LNw6UzgkL9Z1ml1QPQE
QFbrH3c8/8NDZcV2jFoNEfFGqYO93UoGfckZcHXZyINvngoQCeVuTPR6bhBAISmHfK/kU+HuDOBt
ei8W/23oGe6KBhz/V3Zyz3JN2eRuZJFXAfe5RMm5diI+lbCB1cCvVrLzp8JyWHufzZf9ZGS4VJN/
HyJp0wpmoH8XWcyTOjeTZWx3o3g6KuPnxDSCGPsVfEsxF2xFvpcdH0nD1t/YBL3yc13SDm+B62K/
JcrSQEv1QubmqVlVcGSLXIJsP8zNeEd2Qu5LBLpkFfb+aejqOxpfV49AN0vU1X0yuN2pIzn7tokT
JjgrSo7Yt/gv/dKv4FM6Iv0B4sTkWADfLZY2n8w3sE4Aud45dfRuCHDacGPdRTe242geGBfapd2X
cg328IMjyfNPkK1mIlqq92i+Q8q/R05cS0M+jETHBE+O3y/l/i0gHX5n6nX+9SLL+SraLjrussTt
ndLRgyyxRBCBR7SOJnamvOS4VvfM3u+yzL467HyETqOHzbHuFTBDRvBOSKyJ4q6ehvLCKJ3NXiRA
ZZjzJIKitkHyd+zsHMxGWDAbaoJfowrfThly5AmmAtGMFzKnzom1psFD5+8Nv5epEnzW/iXiUbBj
21VvJOEL0GR3rXClKpMzx6FL/XMTILfkGrUh4e5aiiE7oriodR+SZFcE8CXjKBbxti5vRTI2VFv2
pJS25KQ0qoWdwMXVEecNjcI7Gi9XCE7GhR6pPLMZ2LIYEvwdGHPuj/iMtrQ0i42UCyq2QVxqzKhr
sbCgzweR1KzVfRXt1O4eAcrdvUrndejr/Kh+zY7mKbl7XVoY3hoQMeHN8vFQFYw7lVZmoarCfJJR
gvtK+afgPpK/1cx+/SC655llWal60sXwUGnp+0pA1auCj1G1VkzNJMgYmgO/sIrmAXXKsWvFCNyD
Lja0IfwNUwhCT5t8uOqJyFky3E+L0BswPKswhK6ccFDqLmJnwlfUFXqOl45qeJ+cl0P5eHwjlU69
CnWyNQosA1+hsm8TYbfWaGEhZp5t00qRmC21QMaD9bRa+BeVaaMQ5PdTXfojtyvEoKhYhWmYw6SM
AN92Sdj7yBEk4+hD1wUvQ/PI5QlSNitqk8EsBIbJPfVVDDGCJ1ZP7FMGum0uSz2jtjxjF/a0Qcvd
GMubOr0awzVRm+rkAJ4uldXbEpZ/bIHTRkMGViMUKNyFi0ur3aAYaf/AnM2XaKCLcjDjaJu48YFY
IHYbdUf6gm/ZBxQn5kV+niFQVdqVkzQpaFmy47IT5uPp4UxHXML/DKb0fHyyo3eyb9mRa5jdfIY1
niL6pur1CguqGxgx7FPn9ZdmQGtmy9rFAk8aHTsRkXbwUlFYZfXq1isC23j2QpgGAbTvj+p5Arfw
zHgviBsNp9EzkZCZU+hELY6jh+/3iwepokpvPDBFqPDUC/caNrOlZUxiJssQnqgb6sGdStAPc+E+
Llm306IbBuX8XHmiGxnlerrf5ljL36I+cm1Ev2RtBVMBf9aJBrV0F68dD2iVrlGjhZvZIUFBn/g5
141RJDrnN/dVx7tI+R5ttNdT8pX/DyxmjGV+wX13OR0PicfE+LTlGkypIOIWUOXRWIDmFziFelkK
jTOvS83Wqp2mQ95CQwQ1sfNI7gP6jRXEj4ps0NDQgOl2E7TNw33p7RADfpPMsNjiVFtt0DEJgEyZ
og6lHF1s/3Z81tj++LrBGzNkwWkHDpFQ4/mPHcPNCpjAAq7qiDR3FsvxGkuifeyp49txbu6iYUEG
PIsxcEtvNGS1E2u6aEwHmUzi8c8bsULXidks9uXv0t8na6Dp51+gXVnl0xQ3WKUuuounG9auk1Nl
muIGPvKy+ZiYkhngwdFojZbbK8b8YuZqrj14mhMXRMpRkolx9xsqWge3zoAXuC5gBIIEux8ejWlQ
6JZqyaKZFKy+i3sxgw1oEezBPS4Y/zJPNoEn/oN/vRHBGq/5eDzzLjfU2Ja6Ie5w7VeB020zkLHa
TidXn7BVxpduhFZtDrFH7hhXCqYJxMvlN3rpP+6/KsAYCPETOsr5vv3B8P52LuMZT39uTJ9OYVvE
cb2j6zUhuaZJOweU9QLL9F4y7K5RXaqyYZS7CXVuCgq4t1OFSWuXeQDb6WACExxVEWNg+4VejeGv
0cESQ3YkXm3WNdJIiWNOrfUM6z97QqoY/xAFL87gY5pvpYiBSgzD/6EA6MVHd0yw+cGSeFWwSJRb
j6XYLzWec/7Eep8gnaVQxVXf6y+PrVzYD7hP1Gu8fI9MO9kX0q4fXFnt5M9bYY4yIJ7VX1kWsN//
si9pm9JfYP+/qk/2MsMxIxntdniPvhb/ksPWfn2MX0Mh5JRjWuNzPJWzLpHwVLMu+fPhrdp3z7ky
N6pNmytd0evUnKNodWrQhBU23l4CGRV1D1YVR5L5Y29WKnMBiOr3OW2LQR06qWq1tBQeO/c39sXo
vlrOXNnxnGO27W+Ba9wACPOyqdYScOLyt05lz9/XEyMhjUtm2FMPDRFcmHsel9d9d/24ZiEkXDlI
IDo/92/Rm1p5Tx1J41pvevfadenxLTLXz+d0329XsCT0bAaTYe7g4uhorwZs7py0S5PfQLWtpvO9
H17sTPAMwwIR334Fxj8GQm3g/KuoyklqIyiVxsq/HeTOQai/bU9kiUhDQ4rM7OjDEBlkahgkYmyZ
7Ixcc2DtnvXre5dJDFM2qBOaV9wTkpOijXIytXBjB5AIAsvzK7iTvR34qPNCS1JMlSPbBehLFyg0
fzRsJd5vNr5shAdpfyiC2qY4/3x84KpAMlC2ZOakYIH4G5HrL5z1+Da61xocq7spoSOmXSaZdsIR
dgc0jliRT9tVRbxMOANqkWWLOOQN2C2e8bCLl4+aE9OLAlGfSQkZy+OGFYgg9EEdQX/kQ4q7nBHU
InZuJi9RYRTz7E/fr20Uhp0QpBQ2+OTx2a10shSqR20aef5oCWHho1tqw4gx5hmzowJfKIRI5QFp
E1Zco5iNFP/lJxE2wg2fPjTPgV8deKFOiIXNSZrt8AJ3rTU64eOHv1VcphgZkK8w/+9/NOZg7j9r
mGzM/3Szj0vPDytnq4iTDwp/SBy70ITp8zmzhtnltSZKYILJUj0k5LYdcEKx8Ru7caCKV9/APYoV
brTbCjNBWSbrEguQTfz2PXomyuEr/XIrMOnMNMlT3Lv5BTRpqvL0RyioYx0UbhyYM9IZ4vfwNTiL
Pqw7+wN/LGgsDYlvzoQSVtg+6p/HWQ9SB/L1wl/FP3/3q0ciYv+/iLTtEVLJa9kV8BVcgiid+2tB
g46Y1EER8+cdaijbXAUmXmxgF8yK9Bv/hBNj0wS9xh/OMUNhd3kFtTGEGDs56BNlJw8f72OTVpfL
WJMJc/L1sy7ha9E9YX1lTclFf/T7uFrdTt0aTJaHodv//fF+O8IygYgfLWXuN/Dh6bvP2kIhQcbO
QY6GmcFSFv+atIXnj6Kg9lhoLNM6D7Dz0Ar8wzo36bC7FyIoU1ST4Ha9o/IsGMYTbsuSz0Tzg7Re
I+07H8cc2eYz2XgCoE9Bb77CpIMx8juJ2Q43KJnhdx1Xf4taX4TXIntrUttEnlrpMYHa2hTThA3b
kP1rDyRlgozOzhlnsf0JDIzvBREC7BqpbLPZXYH97K7ciU+CgcOfC2ivSTSR6fgkKDihNOpJhozN
a7Xoa9lUHpIBgGEwZFaD+0v8DusyUXVRAWWnAn4irFneKqybAdOWU9NYuBoEHNbEDq4hzotNPJ+Q
9PxjXtjQLQXq2e1mm+dHOrn0y5L/afgDvGoM+uYIzHnA0xhtTZQfZX/OxndmQPJLt66uUKuwIFej
/LtDPZgZfbwy6ebYI7Bt+UVqwV1YpKKtp2H2n/Q1D3h06Ea2vW2Bc4NxE7Ofjj9t5UuuMPq9bv4m
JH4Zz33Jtxx0GTX8CpD4+UH03vobiUCffMoUQNEDIZ6y8W35U4BKqWfpk9m2PmXKZVIhQYJeG0Y8
B8C1J0Up1GuIiswN4JBDTmDRzM+UGE+yZYmcdH24XXdH7WrPvzu41DqzLkcwVg0QvkQ6z8Z0gnq3
EVf6U/1iBoPVVJwMZzVh+tvHw+F6MQKyemv9B1WS1LU6eWxJtHApctjwvBWBbeiUc336iGR3YvMP
zUGDXdBRSjRtNu6MJRPsWtyGNxmD2g0cHUpTnWVkWGPyI/eFYkLPL+iwHb987D0c4hcTHYv5aqpO
0y5wF1ocBJNnlnhDPMDE4exKWDne4yBynvjdr2VXAaCKktRpV/AZnd+KmwOwZ6sbyZ6DHf6Spt0X
PYbap9gyIvaGASD1AnyNH7gjx62ZJ3zVysnlVHXt8Lm2UtSB1Wnwxa2+gw1Q6SxzFE7UJRemEGRZ
DQiR8phyLYQmZse0Fbr5hEd2T1fk07wQ4BdRiaSWc556z+4vrgdbmoKz28YbKhN4cwO2tz8SD+K4
cu0KD5vhh3QJ7AtsikZHVngcHwYi02I1oRfeZ3JYKgiCY70Ls6DFM9Tas3Z7ArXkra6Wo9H/ZMUx
+ETBaDQx7VVH9D+Rq9SnitjSGiT3EfPvFAOl1scoidRmSapchTuNM4VjRgwQBt17NA5MAsPhkNq1
6p3E3Nnq+9Ot2KVIQX6SvDr2vZ00n/BvwVtBy3bDgifEnbTiqFePs6y4jHQuGz5+9zmsrRsl5iz6
w4v1jgd4SNmwOgwMy6/EXIXqrrAGJQRMSOkgbUWuL3scM8dF6gYofaBvfXRl7og1zD7vXBqtpLxm
XJH+EQHVCePhGfOtWPh0Gf3rMDj13/sPLlDzhfLOuYZmfLoPYM37fni43UITLgLElfm0SVP2vQFg
zYpqFBQJW+AT2ZQCjSYlLK/hSHyQ9rOWfeDbu88kBIK/R7f8YJcKRYMx8P2MZ+kEMr6r2iM3cRBD
w4R2c/Mgb2APG4ddmFzYqlUZ0MD1c631iHga2BOFrigLdZP0nI3lryxelnMFEopA36IV6vs+y46z
Q4OBm1KVc8DWCWW3wsdujWkjMg1UspR6i6TYSYZsOB0VJShFEWW14ekSjNcvETQke1Xj7VdKNAAn
qoc8DM6/3z6oDxmp2EDXzc23s3p4nhhTFTGG+op4m+q0x1fA4cwShjtswiK16LaG/jOvKXZRv7UV
+sh16BV5VYYks6cDXNNMYAmEs/GpnkMq4MjU9/6B/pAbGX5iztjK10CzANOIzXAUB0rGA2/MKBHR
rtJmOTiWVmzl4hl2zNhbwxOM+ro023fafEm+HQLbHnXgQNebKg15KkFlZqOAN1XodZkIc6oHErys
9bhEnUQwfUab14UamLqo2dR+cvsSNOZGp0o3U1B/lT7fWtjC0l2PPaFBgir/6JY4aRr4/ccd+VLC
tTvYv6tqO19yjZvcxyGX0NAzjMCD/WN8jMWP4UxaRl1oQIFV0RzSdAAGyPCi537WgseVmuVcRrkB
StSqLFwuLoVgvwQBl5QHurslEbHIkd4npvUV23Pw3N3RvE1tpiIk0/m9sEDDD6Uc5boeAnBobQyH
VbaQijFVZS9fl7B+cymk5eAyMyEO0wW59hPTy/Wadu710tFlO+yy5J/0rWXAtnyCnLxqJQpoh8T7
B2B5STkuQg5Gyc1aXlxegdKX+NasjV8Hk9qBqWXjbNWTXhw5mo425IutLXXXHwc0xubVUpzecqn3
qRfV/KbmcLhXbn6AmTOF40M+GIXKT1Jw0N7MWGESabacWxfnviw77XX7kJfb4o/LplLJd70o5bDF
LxOlUYOJ2TljAflhvHLiyztYD61lUCX2/18ajDSFN9Y3Ubhg1hYWsQu2HmOZq0KmMXAhRub7KxVD
gm0L13S69ewdVBZAQwzhWvyEkWjdLXfalr76rs505oPUwPWcwHmpWW/LjPknUDN0CVpzyxQe9uP6
GtmSoq6IWjMWt0kzGg7N9mWD09cVYtYakQIsMi0pP3+gs4ow45yIoDWK2i80MoXXTn9fqJJRc2le
bCirFewZeS8VSgXjOIh81RvQDW5c0n/6+a5GPr4pA9WJS4hk5Pq7szZC7E/go4vPvix7y1OcQsGD
iuNssISLfjZ4LP/q4JhAMqNBtEbbdPug5fI0HGb3pu9bw4diESpRr7IdS07VD01pMwlVAvE0gb8i
n8PWtMOBa55SmYq5LoQd/nLP/irfwxMTgrIlFETVv7A4LKvhfNG/qzqD9nEut5H0NFqTXKsXG9zU
L2R6F3jNy/TjAERwOoVEd6m2kjptoksV2Z3IEJKh6YXPs62MY10WS1Zr2gOGUZQgqA+s9bU++7z8
0k1PYeos9kPZc44zPk56NzqfgEZdvBaNyeakHvztrhj2rybXRMYW6ad+e7Cb2winxYQcobBzbXhT
kEKe0VcThJ/V/Y64yhkUz1jcrVM+X0mNa0vZdwkDnFkbhlhfrRKC0ny6gSuA165tNLWwGgo8gTnI
l4N6p+8f4ws/lZrNt4hemBHuNAEtzYffiguWDGcXQTBVTY9P1fqXiFD7UXQmEph7TJ/CCYeM3EKF
AgKxz/bKC7KeBF3NidBNAhB8ZU5qBHO51Mg77apMUPgdLB+e4IffvG9fvIdxpLV6dgKDKoPsc8wM
z8YvJIEsEPnTFptym0RXRr3tpaacZKlzjzfzcGRAYkpoLbBzSnMPy8he0m2fF1Qcew8ItZW0i7Gu
iKpBPnQ5LGpBLBw1vbpmeCT10NHJHoO11xvXx4kHHXzJxhioFeQF0Otm0bAgO9b5MEXmhxTrnrNY
IuWzDgd3WtF2ok5vAZZqVVPIVlOBQ397aj5QS44uPDB47FEytWLnKyten4raL+u7t/MSj33nP1cP
mHjXSZKGL/6NVEExxIaq9I55VUfcP67Oc6oh+mwq546Wyzh/AJWsGYcfVwIKkBMWSmDq4/EltyD7
l7UpYKkBcKjlPL66P6Ewr5NYNTMq+l2yGy6Dx8l6S2AYI7rPPrO8vsfCoYZJygs+Ap2HbWUPM969
q4Xj03Vg6U0q2mz0T7GtOgMl652Y5Dk7yCz6tCJYfm6ZxKs8UdwJyVkceLt6I/Z840kuGQlSzhPJ
Pf8DRV2DMaR3/pKkKLFENM66cCjh+0xem1QEe6fEmKfICNjDzLcr2Ur/3+ia4wYsiLsjMH9qUHo5
9U855IF3VTP3/gGgahI4IqWMLjvfR0/W5+awhUnIi20A+j8gufd6sa7Ia5MFL+Krvfy2XPs2Qzkb
Mll+W37uZZ9wI3/o1VlGVwwqXc1120jKsUA9sAmsbJ1FUO0HUXAn2gq41sMb7gRlozBAodU/8oTY
m/rsSpmJ2kGXFDqVkTkKhmG3bI7xtFrm+Cy2N79lYmYNHwZseyh/oDTQhvByvIGQjZrKjqqkIP/p
wkpgJcYxaKF05MSI64qX0pwoImjUmde4h8l+eExsYl/Zhdx4HxWdTbjik12p3NS+NYNHnLtli5bL
9lyahY2H4NkHxzqb1ADdtM7BOWGL44swWz/kU0b4agC0QejkbV7Om6NecYpEQKysLZ84N7AHxlVx
/JksK5QE3Gag96lczF1xj8ZoT1gon0Hu5IM9TMC0dXb4M5VAy/jCR8H20+kVaUbu3buHcCs0SnbY
TL4fwqtxyUfGtoXcx2HnRgdDXWTl+LyUAkHGkRxrKXW6UvIEfhaU+ebNKqlnu7rTGbv0hkXu1kzz
tAmCICznGDUFWSMbJPxUT3MniEk9oHY0Mvij1r0bDhDK8z/B2gG09BEZAuVJTP69P9NLR/vgXgbe
egvXrKbtpBFm//gwtsfb/kZmGuZSGxOxTyu1IxeGF9tFthp5T7vnR7t2lgTr/hU45Odf9AHbKhwZ
Lt1KComyR5YnpKetOpe4DjaJ6EMpvEZRP56hGgo2W+WIEQF2Q1wiLDtdZp6M+CjnMwOCy9ZrEag/
feKNLt+uY62GDT5u1nBXGWw9XADs+Y16Vhmp2IkQlpjeNheAJ5V2Xhlra3Ft89l0x0mr/WJSmeWw
eNylcuCg6mjnMhkV2JeS8qQAwyOXFPLksrd38vOlLYs6XUBKV7q5MipprtbIU9dWTZl98/MphE7I
cXvrpp7cr4b5jDPMJynZejnV9QwZWiq87W2ik4fWwSQHJ2t8mF2I7fDGX/Pu4SLa8WkS2VxVLMWL
DrsniH3xNzxOXsuU0h93Joei8k7nLCc157JUNG7JNLZkA9kKT+4maD4c+Y19cf/CG1sLdn+VmE8X
CfkS4qEzHPtwkenesCnORa2+ESaRib7KdBkR0GAGmzA59J0igQ9aIVJEy3Ud/ml3Jfjb9789LKE2
TUElFXlQVI/8RavpcGYn0M2VqV6/kBf9oLEabuh3p6MZ7A0aut0FVxJMn0qcSeUu8zIGYzvNrxKt
a0lAH/LBXMTJtn5BYcd/0+LF6Nk5BJZDeB5JGUTT7HDqSsIJcgKrOrG8mCQz05Rp5//acgtl/Faq
KUjcSss752x2pz7Nh+3Z4H17ZD2jVJgGLHxTKTO/punec1aOQWO8rlpL/VoPi2Ca5iQXUcB3qxEN
9wnmNULq9V+t3MGwPGs0lRsuEr4+GTjV32/nF/Z5pK0Pyv5JZnCqdYAF5eciREMNWK1AtNDBA9sB
Ni+Ig245t+P9C0By3XQ42rxrukhKRV+Aqgfwx295gT3JSe95obtlQ/XjgtQJEH3kYQEzfERpKQ1h
JoZghgK0SqbHGh+LnwQ31PwKEmpfmq5f9eJkA6HehQbEEGqf4v4WSK/poYVzWfg7zx9/pAg6XyR0
n6uQNwXhMScQC1rB44BngdqUkAA60rmSngXOPVKzbzNXdHGUwPnuy8ehYiDoodNH5NQfARHwlDsR
GpuoxYaxdr8mnI2quxC7j7CvBDKBREy/ku7kobQHM6c+bsjvXzvcIln1IjANTH/VnrJczXdIT9d1
dIGf37+HtvZOCE/pQ3A2VDE7YAMUDVKmpNweYmVN+vkLO4UwRs42GlZwTxYCPkAZ9eIXA8el+gF8
71Bgjk8Y/eIsr2ES6FOhcJfKsSQ5b87UpkfoEI7/7l2hnmuL9ADTueQWJm3LTIrWk7g0UlKZzFEl
CCfx+78csbO3u6zn9o5EKT+q7bBja/gjC4Hils3R7HY2Bhph4iEdKE4QWMFCD5X7LyBNExP7W9cX
f96cULz3n1JwTPUw4GZMmTSdRCikMaHwAxtGQs9H3iM9/HzL08oUTKY2ithY/WH9ac08+pfnc6zO
ybPsjJGPAgaNNiWliXH92+LyWY57FkR2seb/WCX3P3tWTjEXUEluZvFOVk+JeiXac54Y4gOCUQTF
co46pU1zS/r48pB1dLAX3crDwWFteiUuw3A0D0QuSmHVlvGIMmEKbwZwzo6vKic8GvyIe+PaFZKY
2OiaAHI7WaBvQdzbDGA8qjTcx7oYS/amoKUeqCJUbzjvHodzLt9Fqzt6ZkFtryYQSYi+Ez6/1fTv
pvXjc39PVmTCQ5Ym0ha9fnwXI5J3oeIdZ7vYW65rVkOdlCSu4PzJKAZmXmRQnSBVP5sEinuLrhf7
dmIbpOeQyLe6nvCC5vP2rabnV0BUJ2QOtuwtFUhmrPtrq+v+yujsqOwStNmzCgPEYMtx1up3t0XY
zRO5EPMBwFB//DkqzPbD5luSM+ljZNz7LnRNKpu2diJVLd7QawjjckUCCSecSYcwga6VeVQAAU+g
uncyISMtxZagjLL0xlib+O1A1aT4sfv3CZf2nIVRNpHf0t8ZIXw0iW8Bq7eljmpGEreIrQPTbtfq
fkoqZy3AED7NAllz5lWHZpklXBrt8KXrkzcNMMasaGUjW8keTXNdu6ZaHve1SsgIluSkhkfJc3yy
FEcpTcxU+JV7ANHYTcqAvc4mXy1EqQ0cn2jKWu7V7mbNjzB2xoP2iY45R8ng5NpnwuIpA5kdlHRQ
kXk9NHH2VgmR1K7vCoFcMgKCF6ar1a4NYfy6VQyKWrdJbeh7HwEFkKDPBUA9/+s+G6GBHr5Q0ekF
98l1O8B45y/VuNpfk5rJDxWwte7mpI0PPpmohbJtQyX/pBtqc90nukM0BB+m0PtXuObwPFj25c4Z
MqfKsMEM6fYB6wx6uKzD9Fh6zfiEEP4lQt4VDU1Q833jfQhm4Tnl5Yvzgguk3nIoCMj5B3xXRN1r
BW9GIzfPrwvTsi9612WlWXcwoX/ksfj0M+ZffwDR3dWdKgT8WkLjt/2zSyp4Uy1yDoWnGsadTeeJ
riCPJYzHEWrqxV8NGW2UIRUJrFx+brFWGlSrS5TLhkj5p5sFgucNOSEhw0vJfzbAkLeQIQxU4NfO
9NC/ikLyVFZ2x2527wK7wWfxCEl0VoXxDv5wrn5ywOvibsEhRB+m2wL6sahYVhY2r+2OLXJDuMWe
XoaSOHwek8BUEtpRhX97DLQRHJxYoSSu5rfuysZPilQtALRD0+nwWq5f1JLltovIa2bidazRcumr
FpsWzsagg7vRGTLqwkLwaKIJuwxKptgrCnYhKmt1HQtwtc5E4MgsnEfsIxqLvmZx6/TsxUGn1lKv
rnkdfdUg+WR3f5n4PiaW/Y9bbIJXfz2AGtxbeuYiHNQ93Wdp89SGhsTUcbXwy+04Uz5J9ON+6tiW
9xdian4ve1mtymff1MgJ1+SvNYVWCWSoGMWaBP3uVIglD6X1nwx/wIDkrBe+vsoFU1uLr2fWesVX
SbuOo6VrZ2LnIZy1e/UudWYsGk5D4ccn4XWbn0ibJ0B2DjVQqOgqr7zcRLU0PrkhAThxEim131YH
LqCj6lUhFvHZIJayNxWWdHtGz2AkAdM5GgLdyA5EhT1exgyGBgdUZ3Rde56AhJ19P0Brpmsx8b5k
iZuGaSLocNGqHo3acZsvYq7g14lst6M6r71bP81nXkE03L5u9NM8JPRYbV2GM4kzHp7VZlRWceBd
607kCRVU2CrZm2qsd3tB7wURIPEccNzPN0MsoDv+D/aPiMSqlMpNpW1cRKw67/3T6Cg6f5ixCADa
8NJPiwkqgnQZQ27b7YknEIcbQsq4peruYRImDRZBvWyzW//Sw8OMhQdk9QH+CF7kT2LKBgamn86o
NMZ7gCZ3G7vrgnbBY3Ymu+oc66x/4cCPxFKWFQ0nvrVQlPoEBZhglwMKXVHC7KanytC4DmCbpwEM
ub7Ky7oT4aBDNwc+5BTeJEdJmZh7+29JrqdXqVHCyeAZYNEGUDxrJ6HyR3JRj9OdhsJkhotAeirK
szowbTAdiih/kUYDaw1qitkWjEidPDGui8qrvFMYXdgh+zUxagSDiNjdz8AOTCgewsDQaT3o64kb
KG5Unf1TrEOmjtI1AO42dFOe/7DGkc4vdzPmOprmlxy/aOL8WCXVZxYzbYTUoDEoxaYWqtIf3t0S
6OAsDzSAhd1VHC4IynF/SWWTZHkNRc9kiAaJTgajgUVeBMGQ1Kq08QZr56XWKXGJ+pONbhfVFgQB
DsiwaoiPLa+vzCfSbR/GjN5CZ4kiGORCGrew6IyccHu9jZ4jQsZT40q6mpL+yglzDGHLQxoghEDe
NTdHbYaCCOwP9PFre+mpvvB8ohgKd9MeuPJeqBLsjOQMkp19jCn8VzBDHa6DxfFwlMH3hM3nTlR9
f74bvN/cWY5D4x7p0P6N2YFrWrWPsFWr1MJICvUPOVpKGTy59WZART1LMhPdaSDc5ta3PLLQ6rUt
8CjomLuerQ7MK+9k2C+rIyFbS4CxtrBLk/gcQ9CB4oNZW84bOzDCjqzLl+suMzBoU1gK+l8m5s+U
LOnrf2mG+W9EdbNFBDG0h2P38FacJ/7aTUeVoZkHQFw+yb/ukMbBCGQLRraL9AhKuayrmEoxTaCx
miTkFG8/z+o4PYvnRIqqmDz3iM/bJV3JlFO+T31oqimYbRWO3rJ5QJnFh/tmqmT+m1DTfH4zugbh
0yt9o+2Vpyo05Qc5v7TMqCwHwmKWHu89V7RU71jPO4LdUOjkg+PDI8FN9ajmPkRZ1jzmN/H7gdhc
1oMAj9B8mPa1FxsH1Dvn5lnV8dQB7Dz4qvlH7OuAyZO+qiCNFqIXAbtx2k/kC1ntG2VUycZaGqjW
m3nu3Y6UiNLFlebNPS03j0F7v/VEB7Urq51U/dMZOtFjEv71+akRd4rvhwN2MM51glynNWMvGKO6
h1gKhHLuxDgMK1AeWmc7irC4hDhKMnqhpQcY7UQkdTJexlUmfDOapOvCcOMV826rbCdJJg7AGIrt
QpqZIiT4gEYALc2TqJ7aODW+Qmj73sPXtQKygDgMNWjOpxj8QvpohsPBb2c1drI329bQh06VUGGP
2/1F3Nhf1LgZit8FiGRjZ7OannF9BGBAkEzo5RlyUxpbTpXmQplFiEGhiyNSRdhQOiR5OW96G2w0
K5Un8H8VGUi2sq4W45asMP3XMX8lCIwNqJ5cgxh5rGGh7khZFNEdOhiGYKFk3CRtvmA30LF3DdRa
qIPq3BcP1CjJdbeAPwEnyZ/6BOM1VeUjiuizZIhwETdeoG8DWBO6bjPOzw/rvO4JMPjgeRvG5q1A
Wp3eQAhoeREt5EMKFO1pxrOHU4Ckm8RHPpHEJbzAxkohPzoEt4Yydej+CbErcG2YkyHwskYciV/t
BAGJm7kyH2MKny2Rr1fKNSg76EriuqKicuKrWw0tV72gyieIWiIvJ140k3wcMae0eQg9O18tUb0N
rVfanYxswifRo37DPdkO/D5TyDfpm5FwfBnPOESgV/lWW6BnE1eC5SQJFVoJc/ABDZyrX+65ZYn0
PVGtMCyGO5F4edNqerPiGanGIcjAZkNqBlJy71ftaFYRjZ8hIgAB6DKEx0iAtoxR7YnldxZ3XuUW
Ap8kNw/32Ynwuu2ifMHj0UObxpmOoUSum9wArmYXQjflFd9K7xEy1tDdaoyZytQ2kS2km/n6149x
h3XLMxDBOHGlc9p4nlDF+OvK6e1bZ03tE2dRXlQtk3izqvpNHGFZciikGGdu7PjCcuMEM+7m9cqL
dlMV65MDxJbwpdJ6GkFepLAU4eJs3FQB0ufUFAv2/IlUBi23Y3V7g0YJcp9T5WdC1/fQzp4qF97m
bR3AHFlP+h3PgnLj+XUTQI11cSDETwFjZT3c74lNVxgSxdShfD/auifEplIeL8GrjpQwJ50+J+2t
hF7vg9683Yi62ZmtU0IEnBd/yO1z3QQdpMwNF0Oi0vvy1Itg2yAEWR9gRAIwGt83wbBUqHUKMyP3
MOF2PF0BYgmmmEpPwRZ0CKrGPom3YqK9tlVwHXbhwDtSN0sbGjpOj5kJzfjDpqrgWKlh8gpHdNKR
6+TZGe5oMEJzjsQbHDLb0EdDmlpVU/mqkGB0YitHYkkaZlowK3e/B0Vy3jW3OGXRSb8uHRDga9to
3XXKdLrXiXjLyv4KU6gUoyTgvGq6Mv7hGkxlCyNkamsl5gF8Glg7CiDwouYrOp5Zv225+teRu2Mc
mf2Id3ybkT1plg0Z1Z2+MQv38+UuUTxVcJ6vGVuYKCP+4h159j7apwU1+mFqPUTaquseblXMc8N0
AEWObWwWk9LIyBEVqaxoftqjPcBd4htvWzqfY6Ni36G3IgNz4JNnreLT6V074BeCYtsCUVfIDWez
lZjTdmhWMGWG/sPskT37NlerotMWM/1gFKNq9AfvWrICfMF7fyafWhtd4+pNg8pubrivLMaSGni4
c9cuwH0CTlQ3wPj6D6r8/Vivx9XmW3tbdQmUSeu448v6d3vKqrBRVtf7XsorfCQ+LYpGdBTcFpXZ
IUYZs12H/isRt2X82tTeVhJVwtisie+lrn5wTRSgpSgJfehs6ecw7/BtZoPmmCNX7YR+reBpyNXn
LpYYxI6wX8ExIVFHO/11zf83QyIBaoioaFdVm1ydxephAvWTSqVJkkwgwmBCfV5/zsS72h9ZbiaN
wAYEE7doxcWzzVPcWQ7aicByWNr5X21ifQTnZeQTdTbni+AEMnhhnPWsCb3yGR9ei/rwh5bDzd0r
Hw/2rgKkciVeC8Sawbc26c44vR3hcVOD141zkucJFuOrMitrKjbhApG2+X1Nzu3IRM8HnCb+nOUx
iT2QDuxkhhJzlOA/SDosabbQc/6BbheOWpoHA8r2w6QDtnj2cs5GaJ+LWRkIebMuF73pSbqRp8Pg
290GwyIa6161PeYT3ExH4IBdz/Cz5pt6pw2cSizgEgMdxoJzi/Qj9QxQhQOyv15w8rMMT9J3vfsw
CmCHq+oYTAklxbzWdxiUV5U5wBjfMGdryiiCZIkCig45j/FLeW9UKcF15rt5Xa8mXBVAA1LVoD5/
xrR8ya4ZXz8aT1QaDP7uwaqrzDe7akAnhmNfnYMx0jE5ZvlvlzGn2NGbuGHjfNrfpO2WZd4pV59M
UlkywQVpPAl2/0UTAiD3SYfJDZvSWjoI25fyl0DJdAUCA79OALhcyiijdZ2E7PzJzECJEmTDp1t0
UtNkPF6tqkOzM7J1dG6m5WCucz214O1XOqccioP//QsD0DFguyX7g9pWLeYDNqHk5GXzTREo5L3Z
dXeuqodtR8ERYACBzt3jEYf0YZYTUPRupGraKWRbVTLY6ZqeU5dBeTb+JYztVWaNxuklST5g7y/z
vUlN3yjU2LQN79eV2uGG7tCQ+ZW7BRyfnoNWo/U2EWJakDEyjY/7mXbVcm4BXC60zZEXVMFI2nHt
PqGDYoBy/Y4KsgSuAmhAFnX/SneioGV3yvYAwArxpWn0gHZuKChUX5w2md/JrChTpQ7fhii8v6E/
N9cOncdsZ5PMpAassf4XKphkAfr3ag0B8JdGourfYfk849beJX4wsjvXRkpyVtvEJ8AQwtVtSakh
pX6zv0hHSJr0Fm9aLTC/AlJihOhVpb8V21238gJYsK5d/7/kMrdwE2EQ5/SruZBotsO7NKvY6+Lw
ophX7vSsSMxHlgPxQAkSi5fU9VtzJ3i+p6ZKL5HRew2CV7MjuTG+pOiqtTlQ7lf68D86Cqk4QeCU
AftDug5Oc0uqRW1CSlWe4Kwo1ZSTl6j2z3pLZcqLtchV0Zz7+BEzyJcvHO59+itc2VI4ssz29osy
2w4tGIROi46TBmicUCt0Vp8kOG3emQzMKRyjutTra0qYL6EB0ieoQ36igutWg+cGvDfSKOKgedxX
C1TD4r4XtKgpI3/GVOqlt2uTUXZUny2psHmFdwa2UO+3wN+ednpWdMw2wIiwIQqYaxhNapFusL7s
cHHhHiUpWRLoRYPbMdQI3fzSiU+Zp5XC0+SVcbkonjPljs5pykLkQHMXGvXBIAZXy8Uckox18N73
2+29xwJBKVZlDdQpe/SjtljXn7528tC1Rn22qjeJNNPP84ZqLXWzMl1dw/K+BE7d2jApTCghwIj6
sUMhf12bN/zWEz2xIb3bEz55HeO2u+kJTp7GCASR2v2+Y0C6A7sPs/HfBmH6edoGkE22pxSde/KC
yhQZAjOOrCX2ilzRvqP6NxbS3CT4ksrvcQsnOeeAXevpfDWhDVsPgJZgSXQnO5mKbWElMiAHpYLm
8sKnHYuM2KhS8gXRRX5oIsuD3KeqPe1LSeyQdRf1/kUbwaaqrrWynLLzorCnltvkfQUkV4qbpd5h
D7yMsZTXYaCKaPKK0sliu3VHhkBDgqJTv8/9IuGi26SNGPckA0Wixn+vbfUcq4CdmPCJcHCmyRcI
i18gSV/MWvfilYLlL1TESGWdyoKoMlRC0JXNXD57QrMjnTbzpoxleYoKNQermsNqdBwaJ1TjSnxT
20UFewTOryj0b52ZOR+BqMs4Whw8ihAUDLCKjmfUrNUxtDeieQm6eH9rI2vQpBNTOGVM+EHYs/pn
jukV9r7Rt90+DFIhSMXXtuu9ak0JBGGF5IB57DTjWpRYXJbsKqiPQJBH9voyyssIRnfO/8L5JHLG
j7ybT401hvffcGXRoZ2Cjjr23VTOjHteD0qMd8pCYZidmbsdnoz00t9zZyEU2VWgr0oy1dmmypnO
3T/fBDrM0QNn+30yeHEhHXrSsXN/PxuZiZHzKWocYppsQ/WKOwX+AyPXwa7vdnq1ZlvHEvThc1xf
o/HPS1tMZaVZHQjtoweMi+SVDHg0FJRqD1FKvQ2mWhRoBM0cnlfhb9LrMKu0a/x22pN8IbiW7COx
Ec+rXbZOOpKtBEC4fPsI+SEXE0T8y8au/LMlG2hxDgduRpeoDR6Hf4gqndlaghGTW0DFWg4EXTvC
RgH92sJ22kp937X96VPfvEhZIsSIoBrqvZoa3EYQqUTBHCFLTSfULybmeLc/xbj9foOK1DN5etvO
E/dXJpZusAnI9oXbvic99B2xmPbtaGLldvKqIA3HJOcpq4J7U5yDhMKoNZqFH1dXVUGNxudU96hl
lQvZQNfz03xznFNbuuf6rA1XGR1x5McEnxwflHVj2DhSoJm+KmTw+n7Jc0XAi9TogoyxDwcT3UHn
mSfRBoLDxLEVqQc6v/1HW1QQetaMPFtQZurC2cUWPjFxnHeMi0nJD68qMgovZrWgvNOSiZ7/JRbd
lom3UWDPTu6mmHKKIwAiJKaowtzlVrhIIuNSr46b5uQ11+9Az3XVx0LhS4K40J0BGHkrZn5yOD7Q
v3TBHXjjIDJ2bJ0FD1rcjoLP4c4PBkORMELR/Yr1MgBMrABazyniNKF42RYMd3BPs3JYD6ezz+au
bQbqPw1hWwjCcSA6zg+XQRQJ4EUdOewdgf7W3jndX1vYtI2WGnsevBKIpvH66XxkBORTT3a5cYs0
W8noNCj1hYuSxERfjqqBLH3Jnhs8VAFUGCTW6DoCKMefWGeNT2nohtmyMEuGP41Wbowiqxx8gMlU
ZAEAyinRfXdKzzXttvbhzQJL4sPvY6Iu/YbKzEf9JtbanxdtV/urvX3+aZrcWRFBnJYf6K3Cgr/v
p19mm50Gtz1MYZWIMB8iAdQRARsJzbEfA3H4e5X0UUAXdCi3fiRX/agmkaGWOuHEfim5rrbE1h6Q
SFUQQK7D4E4T33SJGy74jrb9g+geJU6hV/Zsj6T+flnm7cbQPUZT/M+N7Xx00CMXBtpFQXpeUAEZ
p1+/kgqiI6O2jpzm9OwTF1vwx7Bj9dfIEpGUVts7E+W1f1bVsTZGRGpW3HhjYOXfmnnA/tzbZqpd
iBQjvECottwN/lvD+c8xndpCmiEhOcYrG8BC2/+wp5fEWVH6KWsN58ejz8rxFiJzA2BkuDUzOZ/g
TmlTBpq7t6GBWnh/DxY0bNmzAT0Z8RvIA1/qgknlX28s2W+94WHUmRCa5wfpdT6qiW294TMSfUVC
5BpTX1ivBGiCWLLy5wfqIDQWTVmRnvUeR/UUgBsOutui9IXkOYwnGBF3JY94E53RAKu003/OTMMG
EryOxJNJcSfiZt2eRr0Pzncc+DJjLHYeMVqOx0xIaTHBHfUJL7xSEjV5pFhupkFUq8fE6x0h0UVU
H/sPHF+vOuKCjFl265rvWWeJBKkdJdujgZGzGtJYreAueUSjQb9HdQsugHjVRYXtw9Pvhokv77Bw
Y7qPcq/VPVuJlRmDc2feNnHt0KlNGJj/NJw4LwOzFNuPYCcMs5PWWpk6wRn/TerwhzzEuo1P4DBJ
00uYND6zWSrwfMvlaZDcqu8aP2G972VHDWhS0oAJk75M/AYEn2f39VFqFN1TsKoK2cI8dT1ZJvCE
2hgxwUKmV6QDdOkgnNAcXUCk0kQPl2bmqSSgLj5avyFI1nap2tYKCmORPlF98FfOSVTCDrLVfP2N
Fjx+q4bc2nlmEnY55luytfBKKoZCyvUGhzjyk6UBSNRZZ1Hw6rNj/SWsFaE3Db5qQkTg99axt1p2
STMijUt3UcU+7oZ5/J9neqyvHnklN0svNNRBKETXkcckV6DI63pLSMgbVazz98nH6Lat2nxjSdbV
qUwb6HSvWB9SvsNH3NlawdrVE9S1v4wCov+8tWE5bBb9sspv1Z2hGg2JCv5q5ApZT9f+okbYXELz
SPGB6azNmcGFdt9oWkXYSB0Nyw3RB/4V86xF5WClLGudx0Ltadm953MrTpAi7gQ3WtOBGRopZLQK
xdzsvFxVbOQ2h+qGEg+DLDuuMGrv/xNneKM3wrGKnzFW31zRFqsFotG9AgmJT4mBZi3qMClT5Tjy
zstl7H5NkbCzrd9+kEgz+l2c8EaQsOMbjQ+ehpSdwWaSSfCWAVm+8MN0Aptxn+8CkyD3fC4ehjRB
wdLkzb83iDCl0Q3TApHIDXi5IAESESeygj0osSBMJVvBvSVzEf0Kjf3h6hmftD5O1/h4jBxWcgm9
GeK5uCVg6QiwVD3DIw4709qa+v1HbJ/7F5wdmPsGgUyVwU0VWd2SNZ4T2oVn4TRgAllWfC0rLoPb
EqtsgMQw8cR1oDZo3uqJjyf4cDj9d6Fdx8hmyGqHhYoXmbO2HdBzU3+egkBTKifbRm/ljNq8OaJy
A+sb6ugyyNlsH1eXv0qvHVv7I5ye3AWX0K24GcgU4r9yjHUYSasTvUt3hGwYzJJZsz726QtMThwi
WYBWpGr7ufEYt/cAjul8Sh0GOVAml2zqosXeoYsy98/OpcdigGzGRb7d4fpKjvzT5TEURCMRjP5m
IrjuWpQBPN8Wws0IUG0PXCoN9eM/IlZTyCqFhDtTwekF0pRV4n640SbpG3z3p5qz+OvP6PrGW71s
okeAAgivKYtKMQ9aeE0V7lOcAJ0HoVluQKbHZ+QTgGdYEqL413O5u6XJ3Cc+3G13VdWwXgmwMLDp
Ts1VwiGUkdW5JKA2+L0HmrH+qLEv7kdpzZFjtP7dAhoy2juI2+7MvGUU0v6EcJ7/mH2fPfcOGMnR
P1SpzDaPPGtmjCtPAHrlxW5cHgJvEWpbfsH/ccjhhCK7xiiA703oWGO/pRDhwxPeNw3lqGH8lsUx
i94OGJ9azpza93uL7NKKsVjiRxqo+AIVsRUNC7f2OzY/uWnvgTtN5XaohlGed89cJ4CsfRdb66js
3PjAEz8ECn12AihSUjAfeAruQWKdwuJpR/AdneghLTDbE2mgn1N6SW3Sdv1KeU57+HaMiV9a5e0s
4VPZNVqmBrZPRO6nbmZfuZJo2tn2L/0IRo9jm0WegkzATQgqp74cYOu0xnlYdg+GMyyAo+CkBCnX
yCVnyVcLJzc1uZHKWayZ9gjpjSKWjXbqWp39tK/OJFnTc39PCOAB2ktDQ9yLYr1/x3lEsGqYhc5f
py8TLb9+liSeu7eOQuvnt7wiMl18Etlk/BgJ6jfbwE1QDWoEzKvFLTgSAoIfyLy91DcZAppQf9tn
kkvp+du35Kk0fFAkeMUUtJ4WiUQOyOnsXmJN93PeIN/6fWuBX3N3TsgQbHQwG5+F4xyVB8vm0U/9
53siI1GnKZfZGyoXE5O7PxmdcioeiYvppz9KfYkoGfdq3B+xbE1PQjaAL5L1obDbCtQwYdX6Ov63
ADVsdayFqG6ADMtyywT56TxAykS4MhsBaTXf4x0Q5mPeiDumbGqutxx9CcB8eG64R2QofQBCsogA
GcdzO9AFss/gMd9YROI7YtSqzifrnHyFaYpICbsXqlZvulmuBUygMKRvS/1xcDwkcLIJ3mmEpFgD
H0tfByrZ7eIBElvaVwbNxHcqf4dEE3lQHM8Xf/5KQMrJ440QTg/VtZJtvZBZt2toHg5U2uuNeEQq
/muaGeGF4rcruZ6UiWujc+FbeTDRRRXt/bbHeMVFYROF9geNTDd7T1qwLeP5zJ4HCka5btEzVCWY
XwRAX/agYhiunMuWTgTwPVjaGGGYL+KJDiylTNRXTEFyM5nbX26X1E7xtRfKqw3s16go2Dr+F0d9
W0inZ/IXWSce8izFh6VfNuk/2hasXTV66gc1s1ydwSB6yShgTHeUyq5Krwl4fS0ZIoJcIuYGxs62
qHCMmzl77H5cFNIfwsSidErb2NUM8WocLEz8xwVSX0jD/eHyppkLATNytgfZNtE/0Gd0JB1no6Iv
avb1GpppuJulA6pZm5E+Oq8JhZuPRwej6iRUfA/UOmjd+HkHFFbrGKSz+wuDDRtI0mtMm0DibpI3
dgQsoWHxfKr1w6wbdQCLG+GPtxIFlYcWkroN0FmkaQyqPzoC34dIU93IQT5bBQwse9lvZBhZnIF7
+D7sXNIak6CeHcvVEz02zCxxE0+Si5rClYoa8dikIFn2CZNwaLGcEB+CqUzvhqc5KfY3PPdRqrtF
NDQe3osiSvnC4W2x7Rtnzcl4Su8vktcF4iPvy2YGQW807ZMwoZx+y1GFa6GLKOr7rqvT1UmDPyNZ
F3dj9w0KIlmcq9ah1rf0JVbgLjC59oV1OTRQ5sCqr7ZpUVbvJ7nyxqzt3Or7AiV9XVVzlFAD4dql
Ti8MtPyLH1m8qExfKN3A3RanQgVacIpUl/bIQ05AmsOfkVCfkcN+HVtc1hCi2G4fpgL6QFe53bL5
FdTDmxMXfLYBMq4u9TZz3UxsTsTVn+uoJ15iNrGHLh2Rjz3SVdvGYUtgZil6EmsXPIRqzwd0gHFr
iGP3kd8YyacVi/Pc2h7fn28rlKcbbuoML6Rvoh3DLiaC7/gKyo8n7iOEJ1lsyC876YQjAExc99Tr
XZVRCamMTgH95aBaU+vaW6xHYWKupZsfGCymanliOmIbQSTj8a6jji6oR2ABk7MlcvYKddTS6kfc
/JgPD6pfPUy7eqK6b0Djozo4GkwjZpxr/S5kXJWRQVsH74ztZ7wyLCTf19UET47gM39k4F/z8GJp
yHTFZD/S7RONu57SK498r8r9xvMhOpJn2pyMXYH0F3TBHDDYOIoXhs+DbboMfxKOF8Puk7inN864
9/E3V8qQeRAbPHrXa4z4N49ujK8iDuTsTf2zFnJqp4Fvgi2NT3y3yC9Xz1r6JHO7Ph9r+i/ZQ5BN
+7tZGiFKvxwEHvagefjDbc3xBI+Bpbxcj3xob5j2qIeMhB/PBpW10pXyRqQ8w5HzNRsbPhQW4lW/
SKqNVcsuOLMyCe+mPvLrGCpiJctuV1IO7WfhGAt0zxd1bjdqd/jRV9xgC/5TsGbNMNhgk2S+Iuy+
S+Y9qmg1FQF1ZxYFWdD5a/0bCymcKIQijXaIx9yxdku+K/UyGIykNylmtWnOv+aRQnL9mhxyI3jW
vcMgqxSoK6tk7M+tjTNZc1Gd339+FETSDqWDGQNoEFxTitViznpupZaW5cUDdBXhJLBESZaBk2XU
II/pnRFt64o5020OTWg01HIExvhEjXLNhIjJ9wSFXBDRRfe/xaVIgzXfy6CLNpANW/WXZYIlY2H6
vsrEZIn6KV0lLizaKWov/UkxCi29BDD0MYfbYmgMzntrCM5n7Eq0pc9ktIT4Oh2UtDydjcZYlo7Q
VdO4F6eLtU6JowWTKFKPnF0SiP/M81myum3yLMVI9tpCapz/eXQ2biY7izvPFZp16s69MGcPLplb
GrJd+TBwxdl2+cfTD7ITVEf++NSowUQuuxDAVSD0i90NRxmtWMw2gTEIFVqGzYSjoTFwuZf0AGCR
m2tynTQ9VfKQs9TX8M1ww/zoSJMVb/PZRkM47KiFfoi9Jp7MvWWnxAxpY7unmcii9y+rLNWnhnMe
PeqZ2kCTy7Txx8rGV8b7Cbb449XNFBAUlVmWSfmMVNrQVtwNXk9IBfSmyYmBGZUb7RqFQOdJRpfQ
W4mVw794oD+qTwzl8iyZ+y8iw+unLddtkkkzJdRBJRYQj/VWxl3d/2P0rjr20xtmVzntvj4KEr/x
VgOnwv1DFy7JbrRoOC2y1TAqgz6rE5B+/52AveDpnbEIVpHzQsrHVuoNyJbghKfT9z1BikYadGMJ
cn8mqTEFcUW1DXBtuAWjeEplUsSzeFHZcEzWyfAPWYickZ77psbhM1DMJ7ZlbTGBxIqn65EVZlvA
Bo8dFJiHOObFrLP+jxq5NNb3co4r7Akd1UBqJ3Hr0VNANJf/d20O+RhcE7t7rc1vjcCf2JeXjqiH
F14wVLbla93oUYLS88SiXRxDG/0Lg8o8SwvJcYcxMLmTm9Xx1S4z9upZei9LfMqeoB9ekpgZ+hVg
dwyKDIdlUIOzsz5WzpPgQq4P4HC+2RP4zntwkWKtKbevO7o+DOhsYJNhyRJkjoQOu4P3O6huYZe9
veQv3ho2jQ8p+eklOOLikERGmlEk2ONrPfyodx0uxw4bKnce3koz//ZnPOgToIctKpQcPwMVl/hT
fRHbFUzBhUoNF9qQgMBvSvrrtmCG4JfFikUaDbZyCAjXabjhDxex7OtOuF5gB7f2/KT8YntgFRDm
bvg2CmeWMqsX4cACN+qSA0u9G1AhPZbCiREq/C8l93xbW+kRlaighkRMMtJbzrJN6Cx0oYBvYjcR
SOkxNuukLSse8eQXN5v94U3UAZssZBWLACQm39z1tdo/zA22pb18kLv7peIv7pREHLIDVzZoCTQd
+id8vfrlbnXGf2Kr351NEYMDMz0q6ghdeJq+DkvVO1NvKa40qHEXEVaYzEh/TF8fQDJXz6i5+ozD
/Yl/ZpbvLMwPps4KxH0lYwsijwXkWto8SBRk9ciCCmoPYkCYSKnuhGeZ2ZE8oYOv+7D8yr/HBkRl
PwalFVmsT502gIJaH/8zdTXwh5imeHwqj7lsuEmXxfhadL+zuCO2Z9dar5hqGQK4wjkiKRo6rE4J
N+CkiFpX0xNAYNXG7d33bifj2WVSlYrIh8QXx8xOYLDpudQyjkT6b/nHIo2ZsvKtHnt1fVka9ZAQ
attmeRpx0LU/gdUD62QUX2uMX6YfaiLXxYMy2HXS0xNi6LD80GNdU+e6+hxZFqwiqCy8Xmm4eaHx
VjrMqey1pGrK4tIA1WPDj19xl05RhIP+Ncq4NVvnm9md0jI9FMJZ+wr6WdoKKSDCPiWSlE+UfS/d
8Mrmpauc5I/59Ax5u1sSvCqhHXZJ9dUQog1B1TeAXwcieFowr91x78fJbuiX6QHg43vN6AXKFe1J
q+Ob5UHHoYMHAtiyfus9e8eMfKwwhMSji6gNx6nmOgYl/B+aD/HUkLi+9k5oDNIhLsG4RuRFZrpV
9TMqo3F8joczKq4ZKCozSRysLj6EIQ2DfszvLN/BcboPeooiiVmS23XUB7f22YMthC1teocFkvZk
EwNGZh9qHR3Xy+kepZVHHtLo3k4u+37PaULXzkWmP7jNDffmxyYOIT5k8NhWAcUQYIgoNzIE8rtR
WWjf62IZB8hj9keYk16YfDjfugaIeObqDC5JE6PUmAlY68U6n097h2BOzEar+OuX9IU8NNK0KPVq
TJxlF4pjX/pvXAptPzmzX30E/mBZa69+ImNXb/mhdRdlPpbl4uHXHUhihbrd4vq5IxlKrd6g9A41
hJcJkmQMVhgyWGvC5K/ci3j6gqQRFf9rfdaYajbA1WIyfU3+5dH7//AL2PXx5lVYNZ69Nj0eFAmD
g3OWmL2kDiPV4opOhglG/4QL4Zj3RKeG+CXdwEii5BRkKAu9aTLjG2tre5olYXs2hihpJbd401UQ
IR3gEWR9UhR6YK57152/gPZ4JF0rqX/3x0GIn6pBCeonb9Iv9GPX644TDXIzsV0vbwA1QsPJO5AL
siFxZMOqiKvOvBB7otZiDURh+nejI7cLvkOFp/GQ8M1fz5xTObQPS5vojbpyl37hpB17wzpLIKSE
UmWgy59SWsoFVfpS49CUPOZQ5QzHC74fOZNZb90zxLYcyk7dkIEDmaZJ6wYEwmLv6E3MZ8HRDkiW
sg3OJ00hwUuyLNpHy7HqhrErmZcyrA6Z25X+/F1f9Bff0BTIq2KoawH5TEN9PLP4BoY5NaCXyKZs
7fbYqixifn3CgOg4eLx0oYLTmpRzLpCBqNaaiEyZu7oybUQ4URwbxSNpnqpJ4+D6yjtr7jNxHIUp
aywL5hU41i8lSIMFZ61fmy7BEitBGehr1Ge2qBP9sT3ZDfRuiF6VpSMiFICAomuN9MI91vM5WSNr
CAST++/ThzUsgRLiecVqTopF47H+gkP0xrfdJqMDGE1RoSPHsRW5Ea9QvsxipYdFAqtQv2t5UhDg
25kXfNxfps9M9rw8Ppcceeg1IyBdLxJqEQiZ2hS6uGAI1aTqmVSWiygrKLssoO380sL9xT8yLSE8
HWHjNlAz37qxK99JGw7We9RSCFMGtSXmwCX19vICOKvaCFrXrqYVEys51Qg8n6zjrjcX3C2YEGDQ
Txes4nKJo6gZSwgUsEjNuti7Yq67PAumE6HFHuaOvuwaDJ5HVCZOuXhDmwcdyUFpsxLsvMq8IFze
gr3x5UwbrHgmOXApoj+tDQK/AhKCMlcb4zvM2bd2Mk66Xsdnm35hTJJ1VQ/FZK/BS+jisMMh0vtA
ZCholHquIbbYVFc98/39O2u2WDzJjKEo6K9/Ei+4AOZCYGRomfBuvif53LC9FWfPl9RujLKQfEbt
cTwhojVzXWCf85X84+UlLMt7UBz7aBJP7SSN3zlcej/izdn6x8Fagz0Eq+6WGEylLGh8i9SBRIGu
tdGoO6OE1SpcLY3uNTlMvDJAd4d0vwea9Ts5uZdJnrPFwkEbNQC2twOMaDWEFgJi57TAjzw1zLvT
vcv2ka5f1CKeNZJdbgA/xfno/TpknntFw47Dul0Isys8EQ1Hfirh/o0lrGhF7o9ZH8AaWLyfih75
oGl/k7p6Wex/LUJogmJKx9O5yfejo1qeejrXQTLNAySLq7l8JXxLqOL26m3r2s82n4cWP0XvlHrR
YGERFlOlpTdHA5p9noT7XblF9LItp6ZRqPnHRFvZQzTm7Nd/GVocnv/wXq+AknFD0kbyqXfbSxo5
mLQYDsRLHXh6fMUGSw4du0Pjyw4LAnUY8sz5AF5pxng5lCGB5GpvmlbH+DfoqgVwRGxyTY4+5K68
ihv32zJR5r9YeCnJB9eie004GVOKc7oezVXo2ArKRuFQ6xybx0I3mfA/cKP8gZj8v87DkOpZNkkR
pMNy9D/PbFHhL1+IgkVnKTJUKLyGnPtPVNvVrid1z9xMOXI4F7VPa3jhHWVfSeAiPDrFGiZMABkn
hzZpFZrdWzAqAgPG+p9hLlTE46+6+8XJIQ3bYwS5K6ISsibLCIYdmwMh8mWeM+mrXEjHR3f3Do8h
Z94FDYb3ixkO2wPKvQD78ENYCn9WeYOQy8+nq0beAmJP2D7KEjaS2v3GBBlf5RNXjOu1nPgarcc2
wNBF17GWDWT9e6YLmBF1hf5lyfuCDKbx2UPolyyMoSHWqGVApsy0SB4h3UjJ5l/EfCYQ+vQUQF9S
06/fXwtw8LZda6VW4kcAzdAuxBDI0qCZEAL3ptA57+RJQJa/dazsVPspP79W0//xkby8g/R3FMVu
dIkXRlU7FNctn/V5WrjMHHqisrRozDg/lqUR0NrjqIGkzsdZdeBXH91ukLw+EQoyH9il53ghAxTl
reZRsIUvYzUPEKK+XS0O3FKaW/XB3fpk3aORFM19rlKphRnUBCNyvbYcgPVNp/HGXK+JcwIvJmWb
s8w+4Lgyk2X7l1xVfJ+GoPnDEz8XgdpmC/wa9pXZP1cqPXNlZbKH9UN0va1CYpHPjk4XwVww61VA
k0sb20SQEHnysx8o3HEPZjlxn1ieUyEK8wuVJp4yTSZLfN7hNIwYEdj8QvOsTaIwJ4BOq3qayDPN
343uFJLt9ry8CaoprArSD48te2/ihUH4VtJrK9+jlO1WRxXdVPYVQbeFqWZyDZBt8zoDpgJf2jFf
z48ax78QTBcYf2WZhdhIl/D6x13h8eyB6Jnc63Udc+I1Pr570gANzA4mtzE6wiUX0zkKqjuzQyNg
Yq0Dzd27Jzew/OwvaBgI1EX5F7sjqKQOJHARGnvf72nAyd6CrR9Ap+9U2N/EaK8hIQ5ATxnsLskS
ezFxFa2SEKPjgBcZR8w91DET8W7jll8uAUfXa2Ss3by+fKhoSlJ89fvLFY5EFB5Ro/4w2qd/qRYO
rcdgEZncp8po10SyFaPINU9GO5rnfWkPJlIzvsMRfDgiIi9eplnGA8ssdKFtEi/mlzuRnYV60BcG
buwLn2lhAccdEIyuvscfE0cqjbanbXCEX5A1fizMcpYB8vIfhKKswVCvYPOsjLWUPxn+jfl3crT5
J5X6CnfojqGZGUons8XVh9VUqF39qBRMutqg6AcLBRbITKfvev7SCKftHbZ/RzyVW0Q0x2pLLlHI
sWhp4tQ/vB+JGrKwuMgoviNAZ/7BeGvwvKq3admSHrJ+Lyo/ThQMEbT58Xf8p9M1AZhCLG0lfX1V
unsTwuJDvu3+rrPezOyA0hUlmKx3A0K9vpf/RK3u1donHeXHVmFZyNHWb0I1fAykFSZGe301pCbQ
lSHsDViDg1SogzDvpwNwBd9qnYiAANFL7iTuBgGMJ0KgfuLjSrnV+JcF2T46yZ4DY56Ax++zDoS/
JtGzv8UqHjofQiAyp8HeczqrymQPFQHfafjvxLl6EpB0cfIZosUlB/xkL8vrCsuLIflpGgEtpcRz
kGKN0YQ1v4q3XYU1wUYKDIaYpVSCLAvfPUa2/mmDKjwalK0zSZrglDa5SZ5DSrJ7VleKm/byaVaM
6ML89hLIjL9qRvc2bS/nPpA7IVZ/k4n/3yyI3S6ck5ZyueIm6I1wZXgiKjyHN48eGQID38UY7fUn
Dg1soRRsQ451y8HlvweFgCSrUC6I4zLbwpfJ3dALlxYn5VxJqnJIzUCpbwF9kRE5AMTLo60F3Q4M
bb9gaPqWF+kNzHIQ3ZAr6HlAKbm6sF+QME9EH0qcR1UGgsFsc+3Jnivuizof5zBeqTFZBcvkLuLY
h6Cgm7ybFzvyEsWZTAjoa5fBIVWQtT/F8wegzM7cqvH/CrJjvcnaaviFtWb3KGLBZAjxt94xjZy4
UELCe5oKeOlMDJcMFdHJ9OwOVnWpi6uum8Xg/6e6e3f79OsnMjSRGH2SrZzFC7Suz+6nQLudGpwT
mQhOzfpTVIGxlMx3z07BgK6hR0tqaYZFDqIPbE8ldwAtyoa86n5iUZXrEkeIwzuS0xAv260+JQlE
gg8WP1nS+azTPEsOUcGUYnBYCmCNf/jwPLGO0p52v1cF5dqa6wiW2+MJd7jpmClf9ObIOATsq+jB
uA7CKpWBzkvbxqWYoQLoeRxvneFDYvu+kWD6NWJbCrCkQjIfkTOXmsjXLv/xvkB2mASiXagzMrAL
FxkhM6t7UWsJXCjEwHizzReXNdIzXEOZxZPW68y8CmQz9Rj4CcbifApalHrKKlK85EAmUc3CRtva
U4TiUWk9i+E6jKMItr6WTZdNzc2MDt1ii7fmK6auBjMa/m3+eFZsDMEig2DGdE+hJZdLV/omMK9a
TNuE0YxwsNmBFzZ/u8ZK3j+XpOrLJj5I2UXgxpwyuIEizWnTj5PShj04k47HLY3GcO4UwQYQ++Qo
G5jgjgV/Mg0EOPkjO+F6rn48sFdM2b8SvWI4fA1VD4vWj3Cvr5PAQiHLxjukbeRfWlbM+x34WidA
kB4Fwexh9U6EvNZTGRbz2dBqKBjC49YdjjVtjFV/raBP5RXZqHfdYQLHAZmlICZ62jb8AiwJzIDm
pMWKETzhEQEvMVu2dpFW11KWlMPnOBG9NrQENWpRvjTtmhL+apcfvbqGqTCfNrzzHOH5kqV0JdZF
LulINxymyNCS70azuwkO669V/c3c5Utp5XM4nUuFENaH2O7V/u3hwsZG/wuAm18B8cc2Xzg6BNWH
+cLe623K9FsHEmxAkSMvWJL6yfp/jjc78P6Mj1aSDq/n/95utKsuu7aaCT2PYRAL8SNYR1f5W2BO
JwW1+L1HoOu7LCZmqRhUAIEJGeiNFkSD8w6y8MvsjIiBiUz9lGgiF0kAxORt2kkZXQ+ZTB1IYSGV
zkXOOL90NYcVIe5FiWom4PHHEyMtXP7+c/NBCudSprKFiua0aQuK8kYfeYtabwrTSkTwvriZZLuJ
mRK/QZSYNWZCHK7MlZq8F2PiDBnEM/xbkxGIVdmo/jEzmFAZICmmgsI/zWlGkbPdbSC7pSBwLTv4
jdCH/nX3nyoPhI6bXy6turKJdw0Agnx8G2rdG+y9zN0YMNkxFiRoekAbikBvCAJq/teFurQnzHmn
vaWW4jp72ijexZL1hCAwG2omAzOZTrH6QKGDMAL5fq7p5KiqNIz0Dm1aYbxeUNkXEpDBlFFR+4VY
ENPrrN6Ibste2zersVKvK9hwxOYP3gpykjRMcSgLSqkP9Cu4X9jj9A/fRtj3FZyZw4gAmLkPU1tr
pnsbrMoizThstccUjQdKP0k5HE3aIQ1BsMrSROX+9m9WUHfCTL6xYTzfN/Me0yhGFKQ3IqqG+62o
a1L2BeeT6aRj6QJ2xm2lnbbNqo7Guwc+Elrj+oIUiifQyAeMw2JLIQMs2G4C94OqutobhbhlVyYY
y2UQ9C2ojhq3qmuuhEpVKj1vGTwMa7TXnFF9gIE7LAcgmkzKlQR548LLV8wXtTrKbNFEZlFOkocr
XoO0OApjG6blLZG4zWfnh2qyYxtN6r7K9OmZI7u5YPk9+s9hU95WhvnVn/n6FYhQw/RLzMl8XYOf
wuCdXHZwJzEOuStflEiHQuHXQzrNMnRcRIcc/Iby9m1W0JoST8oGcg+hzu30j7XhAYw60CAekblQ
wrByZrbA9IKSKWhnSunIsOOrD9zOF6Beasoj4DyX8Nt/IWjRw/Y7fa4bqpfnv+7RdCIHNvV6N4sq
unIwQhd6md2qUxLmSRTXGZaXvI86uCIEH2WR0HoWzlfS4kH3koZkki4r+wiZXHqmVPsAxL3lng6f
MNf+WD7V2yX+k5sHFO0zwF8pD7apKyDWktzCwDgmxyZngUmeWAXEyh7mm1jivty4az6pnxeqKvZL
W7EJex3CWAap67WzgZbPTmbqWwFTBz7tYunuQ/FTTn3esb5CE9dw5yVP4i2fUbSVu+gQ2KuhrgyO
uVXHHNC5FtnaAnGNFzNIh8SdXPM5CTcvcSXhQlmasMpJcp1CWFV6ZiniPnzBHH2W65b96RMcOyHU
FldKRxKR6/FtT4a0vyryga6+AabFRDAOkpdLZhZbj1qA1tg9nK5D7EO+Lqr/5PBxjlPgIsVY7cKj
KImuacEA4oQ1Ky6apPRlv7f+cO077FhraeViuP3RZIZbAaqX8p6kK11MtMcCIOZyLz2V1Uipn/Eg
OCXK5XrfAnVW99lPR9EKOSEUPWAozsRZAMPslEAjtjiOXWS7o7zP/J8xETIPwuXkUeUiM3RZJx+q
mcRyc9x3rOSrL1Bd2p3ir9+Ksb/zVgfZgq36Y4N+npGmNajHweFiMKIXSR9qmpqdz5B60uv4zTEn
5bs22BSKBmCgB3sHw1iIzazPlncpHyiSc/J460JwyMRXtxMSQoCyrdgn3QlbZ3VpYz5dxycJPIH9
7XYl4WW2n2qDTIh/uRNDK6pcpBsU6ebqMgzRfFh8o1Ncdn7F6yUcCem3Wg+woaS06JfCrrXnpNr7
+dWTVHrZz6vIyAXSVJ3K8PLWTP5uk70XV5wbnsU5anu9SL6awOlX2tHqxscxyhn88iLPKNp38zIL
3aiesPiJ14phft66G/8f3qM0XKjK41mtwdkX0aKhQ0u+EMCvWlQBysebt/jku+G9xBRWphnkRlyr
c4Lblyg+ZiqMC6WPqWo8Ihy1M8DmUW6UFSo2CchwXvz0coV8fugppQcKr3XInCDveEtQssRWLJTW
aYEL3Y0IgyZxGvWG0abWdjiI4FtY8ecxvWkYeDYZAhYlFleJ0WW/vY+QqU/GbDDnc7XwC1D9z3Cj
H4fLavxFqXK63p8u6QTfnjLMb2ZaeFtCiE3tPA6kxYGUbC3kSqB2co8DG0M1ueh9ZjzfcEfDmOk3
BqItpx47ppvyUQLf87TlSQcoAiyOp5YBRug9SenM8+OjKKesdEb44RqX3cvNyZH54IntrCaHH3Qg
tNYnG5Y9HSqrkExolgtSEmSVnkDhVUXXICuBEJnCpqUpugXEGRqazn1Z4VywtbfaUiQdqfgHVLqA
2E2GvhxkV2M8i7wJsz6S7qQ3sk8kUxik/yL9PSFDIic0bmR17VQzsjKuSiAzzghm5qINo82CtDjj
tS7H8HG5ZsTlq/98BAwUltfLe0edeU7FJ2cJpPWdFJda5FAV+3hLnglQik3vLyk9+Njw2ePoRBIm
ROGDLlpTXmtdc+ASJRTjzx7r6RYXJlFxP9aO6mVTbYNn2AJC3+SbDh9todqvWmEK9bl17xUWBl53
HAvGsA5W60mnkDaSWqYKio353zlfC19gxN16mbFiQMxd9pC6rTi1xfmsgX1sJCPrudL+OfWEE80p
GPBsf5On8BPWTnjJ14UGCedDPId4Olzqq0J089EgoR2/+ksakuaBfuXXhAxMBc1yTRQz05OokI+8
z35P3q6foFDFKGijuePZGkLoS1vnrAmFKoDUvVAZBI5ES98JoUzOlnu5RiIJhcA9bGpRT4Nkq+rY
jnfNRUCWmZNZ21fFPcd3MXv8n9JJqh4qrYdWTcuiPkAQ71yv1aU8uCF2tyh8jqvM2FwplEe1DiBT
RibnCsr1eul4QiDMH5QDtBHFT40deQal/7GbO+SMKsQZxD3yTaj68AQk4QH6FD5FqOexB2vCNNe6
lJNCvN6fRjFtPIBroZ9jkx5mvpv4DBH1MtVb6ujpVdI/yS7qoWlBip4RWAoo0+SRPHZJxKEWaAC+
EOxMkcCbHfu0xH7GYk83J0SqtKvYYf+eyGZKdY2f5txe69BRlyQFXVyJsnj28bGg3GO68lrvxNW8
+8B6OFU+5HeGt8yPWP6tt4Hl6187KCg+N8OWpEOUymvOUG/mjkkHcaj0sBdd9KLdP4Lf5r4d1EO/
/pM4SGPXvxJM3fLfYU5B4ZgHb6kK/ngLYRtAF/CwsmcPGPlejqMaTM1snUUeQqcbmcnnjbSqKeV1
DGcAVlfNHemAygNf1RpCSptJGpcIA8hpo6QFURFynaW6ZHftHCxjjyY0h3FuTAdZROnJmlTUWrNT
bhO3Nf9MdkpkdD9IGzC31x28oTEzl04ggwBMtzZ+yO8URYBkBlPV2y/MHxiym66AzEHa9Lg/P3DJ
kPW05+7L9F0qemkKn/+Fnei9Ga/sui0fdE+nsSDaGVVjq0Dgk+RqzVd5C3jkdt9ZwjJux4J3b82R
BmA6L6u9HuOSnpSzgxc61v6CRehdhpzD6I5G8vLNP8DNcX/xjqjxcZDNkSyTeC3IbdsQoW6eoQrf
ng/iKpYQd7TGqQ321cEw/afNKX54HFVE9QJW+08nL/83HNuHLzaGVMxZbA1p12RgzM4B8nSJFKmU
/js5imNtUNmYYDh//4tJVZx8yGOlnaeOfT6Uq/OgzNQq3WlvwkLV8tg1UAMUpWNXYboxa43mmA2h
Eqw+FQk5c7dQyl+jrEbLHsJ4S/pt17sZABv6JNY/BkkvdRYCcAopxh7bNEEs7eopDTQxVtFlY+Mm
vA2Cs6vvin8NJeASdHyo1fKHMUAmkLgFIGflWLq3Zb44hs9quf0N8XH0oEL7e3vua0ipMYCEJ5qY
qPHQDbXTlhsLJfXepzZNyUn1JtYu/WdZ1nyflUwoz/+PHVKw+KwdCFXvktIt3pbO6ccD1dgCsi/j
QiGrGt0kI674xRORAV8QGFUjc1c17a2qoW4FJmzSgD+eF5Suj9xXpSu3QpdrLGFgzvim7gNU84G8
36EkrqgjF3fFM7GddvpdWs96VoSNvjfmRLFTqGzc5056kwMLtPHG+XilnrxsBdJlMv2HPaPCnCIk
fIOfKRv1nhnKtXccualT8TeOV4IQSKKxIsqJYzORSelgYM5kzWtkmgrPzvZW0cPvzQbHCqdTMnXi
FP/QSMuHp1A5rjGNhM0JGvJZTniOLEmLQA7KvGolbgLOsse9IVT/Lm1zrQ4S55GnggJ28vKiEMAE
jD9Rl/zew7amVrEPDjthxYl0ISHVDwn14ayB7S2vweEp0Fi6dGWUuqcFzkkABWof65j1iSBxzYm0
22K/4gCWIeZMTpED6ldPEma2C94wv3IOaOJ4cSX/ozMwDW2RVNg1XnUA8gzxIhxpSCOoLCYhfGMG
/QOZk8uRsv03DYFEjQy7+Coeb32plBEt0CM704Mmv64h4NAHdFY2/G+PmIPaTREmLxZs1zhRsrPi
8oomxVx/jv9nxiuTgmeZCyEe1zjGWbnDcSzcvLYKvniWMy4Gy0fNKophXQdQyYpOiC5r7aZ0FH31
t7P+g8JmShtFVeK7mTn8UNdENDE/ruD+e/KQkmxKzwh4KSVwMFgwUKfrzbx+d9CVI4/zIk6cktVm
zv6fFA8EgOAGa49Balv5P8cO90qkvi+Ive6y9LYrvA9/4H/tNErJI90+c0RiaoGNyrmNPhJrf7RN
hnDtlf0T5jg+5C0KpOQ8XwiWLZ3R3PlN3gGk6NRDe1Z1zOSEJXupV+3xC3eFC1FDdg1dgDz7haeT
PDR/xSGP3BM20fO5n9yZfghwR+eIvD/ps2s0Ly1GATun0slqEqWIIAtram4QzFZHnaNMstQGuD96
dNrJ+G8TSIdr4l43q52J2eyJq7iBVzY8gwDB6zRmGrQSCLZ/Q5NaACwx0FKFl5sUDVSateWi9BZD
MFvCFo1skkjUyKqjZ+qvg0SXpebdig2XhAz33jAyPnnSvoFOKkYI+Wq4P4F2gUFVJvcaydSAxLNo
rXrCPAyg7UajHxMFSqaaHqMBONXIWHtEvHS0JHWUI5uWZTsKkj8NGkrkjWMJ35xJtN6JfS7vENzG
W/ujsITFpDkAnFLaw4XjZpsEzoalbg+3jI1TfMDqaHJovlaLQkTj2tYrV0LR/E4yT6e5HU21r0zy
JxbqkdilXCQAZFObwEZK7V6YGlHQAxEWwrCX9D/32aAJhs+8YwDjZPYw411FyueTkclZtgMEQ8ku
XLPqaebew2bI8yGLaV1qa6RhVVjFDawrtgIZ7RBUUCMk7sbq2OJn9mNzxY37LMUJaB7IZX2e1MuI
f939ugpXWTQpdGUfjzIBn5/owNUHhtSwgCSm4Uie7+BybcDI1386IxfixDSZ9Ij9jl6CQ6tDLXgS
HhZ2NrR6piUzUUsMKwAu8Ydu1gzwR3pAdV+v1W+OXOiU7OdoUhuYt8vDpfBVK7K7KO2rqJq4moyt
vRojwcuroJbCzuBJBygGvw+jnJo8F2OTNu7yrVqdrjdlaIsZP4U+99THFC0PCc9m6tij9YXFd0t5
aE/7OM8Z7xGUVwPbQB9rv51jTBp3VGw6KFAV7WpRUDKjxSQu35TGemq7PZ6fqZpenD24MphNwA4p
WKthUST9WMRc5P3ebdM7mUO9PRXtZoaqzycfu23jzESHXO1UCy3IeSN4dy7eOzFtvH7Gb3pVskKT
ZCvzj40idHlm32ORRohn5AOs0aMPmGs3HyLRO34ddIJNmb7o6sGlBMZS2PBl999LTdXnOA1r8bNv
tKa8xDT15hLEP2NFctIlQOAMSwcxRgYuccbRfr9pBAIb8zj2Gg+Om49mqU19IqcdxA0Nk9jbo1YJ
C0o0r0M/QGLgAioucCW3f0hbOo6egP9ZzJkRPDlgC/cmaksZXz/Daq27yqfDwLuUl4ON+EzM0xkt
OeJYfZZDiJ/i6f/Wg2Xf2XTknr8Ou1Jgh10iHwq0jxVUOBN+1JVfyXItzTF9itL/2Hq/SIxsqY1P
vccrTDLKorRU8TXGsKXSadCC1WUUEOVIF+biw1IPQoMbi8C10oTrN3VngLLDu40SinYmV0YcpQvt
Ple6No1Tj5TT30cQtu89DKMsvPINO/QBAl3Puw0XLNKeFz9o04x48HtQatBRVngeFLGX/5zlnyCZ
Ueg9RI9J7VOaGwz+C6i5nJZQivq73TZgvhDh7fH+Wp2lbHuXUk1s5ecXgydsqq8vF3UisOuKQ62J
NUn/KxnNOuFFaddHhig6w/uuucepKhyMLQUhnloMAINIKKvTYQMzAD+zag+Glo7dMasfG2deLNpo
0j+FXDVdsOun3jFGfLZe3OEQR2yGbnwnrppNOhygCEyXdDreLI/qGjBVTC0z1FshPnB4ifA89Jez
GtNg8A4b3Z/VezdU4YKxQdbUyyzUbFVV55YmvWtKdEDKVcYmcn0Rpum/MAiLQbbwUF+68930yr44
S8hHA8rdo2J1mnqGMzwfjj+Tr7oVj7gNJgaJfZDohfkKEgqLNGQiEapq4nl5yjvc0fhC8PagDbI6
mBcgTHTgW7fhnhxI9mKnfX896ykgdcMo7SQCOETnyE3afsEFD4MBlfgeTWH7U4DHxWpWP6uPBTd5
ImJdhGavhseYiMWVnmNFMyswIHdDMHftBoM702DsxQfztit99KaLNrU/ysrtgyHJvEmu6AiSFwrd
y4jTbCbdNYlB1ajH0mN7wIjb3ePldz7+y0gtStkOv2Egr1zzyS1yeydAUEeD1UuC4/unSxJJCQZE
hs6mXUPSYZYXYAoe9ccSFDNuAfDWs1JMc29goYCST3TQ20XIbbHkjj61zraYsd0o/hWA8xMlV0hn
niLBFY+PY+imAS+RIOhZ9D3CrWKK55ir/bLLMBzJpdgx3rE7LHZHn84BkxxcNjyMp0divZGhFOyY
grHgWjLJNvBDr5gnP/duJxumLQ90Ro4/AO3EkEypsC1yeJXkjfa8QI/D2AaBdfRVGN0t+535kxMr
FIkT+fPX1ANfiOzIuP53Ph0cdir4VuJJFiW5xB3cI0E7In/kVCgxjAvCCnhX5XvzV1koVAe8gjYb
NQwI+Q/CIaiezYVZ4ENAZ3oJ4dAApAnA0ul+z8fiOd7mbmhJWz/H/cK40fKb+IzyzyqT+YSFj7GW
2LL4bGRDL5Co+5KLYuTOu8FN5MpmID3/mrlE27oH334+IhUswZZFMkLRS5Sq5mLCCwvkMcAvj4gq
i6ooinGmanY3pQLdnVd1+5p+DUcJSPxldlDZqNRQae5vzKW9C13QVcMfkgGdlMrQ/dwzEOvwDlYr
7ZhNMg/njKhXeezflK5faKqzIXqv7pvg2F92+wAtbKLpKslhOEDvmbz+OwROKZSo/dCnO88Ahp4E
b5F/uZvMRufw44mQIx3ixg8nNq1rNAIuHQy5FJYFSkUWwxPNbJs1jI03Eu6OAejmP9dWJuZirtlM
PjtkUyUVVKkEgnzV1MDg/uWg/WQ+1rvKNjY1j/ktjCwwm84QZGdCO/SRDVShh+V2IcAvuablNeDf
nKQ7foExgjfEyvb1zZveqk+FzFhZhF2NIyAFFg+uUhqAj2cX+v1DRx/8x9eH5i8A3pKkm7xocd9K
45uEj4biMCEK5X2OTsL22Sr8g5rz1dYf8GwlngrFvs+Wo508a/QPNuVrKBWIWyzMfMONmeQQgkJS
96cEfhEVCUVQMy5xx+tnM/KvmIEb2gVQjXUwajIetOEx6ZLdAwo/dTj68O7S/JVs8te1sC7LgYlI
Haulnfvhe9EopEqYVuW5ECBOZjz9WQsMyWa3FqTgWGbKhq6wkviwYfutik/qC/hI4nywDCJ18TXW
TdWTOFssbLvS+TLe02TtpHOWAXdoqfRjT0pBWVPp5uGSLgQ0cLURciaGF6Loi5jf/Dfw03rTleQ4
LB2VZZDkwtpcCYGcjKgowyIY1lWkDtlQKmAJHGGQBgDipwSInIe58RzJCubp7WA5ovPDpITrWbcs
6i9nepPTZhWKuAjUHB7YaIl838AGFDyLDS1GQNSyyE8XabvCXcvzZB6y7jetBuBFg/dFUoau9NAq
5PTb2neIYc5uLihIrBKYstoZwW4MYGB1OYZx63rYbSK/WX6vonykqRlZd2rWMDyCmZR+nCuciK2r
CM1BddqmffgIDDeD9SDhWa08zfsOxgcn9egqxCuQhFO7PBePNiccA8CjmoQxPFCVHpBFdlXsFizw
uGnNWqtfvtztRWaVYwWnlQfL4wYbc7iyie7MlJeV5dVs2XB+TAmWjyzjvoRn7CvGh77qxy1Mwzvx
p8n36PAM8rdhQALHnj5Rsqw0eNiqX/CJmc5DYBehv46SRQhEJIAI2MpfFgCPd2JiSbjjiz/lHP4v
JEmvZQxRROf5sQ5NWISiD16MiMojH6t4yf08K4HvZrGjb5e+nuaPKWmfm4EQYqwAvikwXf7VKoFw
ItjehFFy/cY/uALLnRjLFyyH+qr0QzA4Fgu5nSPW9s02zyXCJ8G7V+GkspOGvnhZm09GghdFKHPv
4h7a1BGSRhsaeZtGVCigFAGUTqmKJ5XamzDnhkTPvrHBNrHgsFH12zKO2zmeSJmBeJ1QnLUus5A8
W92/ZDMmjJA4ho3mDZtyp3oetDEmg+9i1W++7QmtI+nndchPM+IXmk6UNMObgsrOIUAf37AMr2Yk
wZmR36tqeJMF7hX4jAdC00oAimF4UJaND32lz7XmXFjM2vTvZb6Cwq6GprIxxK3ypuJ8evQxVVJ7
QUvCCGJZrvSd/qlgKDjB62WH6EeuWb0GXL0Q8oHEhWFFlDWgtIHiDNbHr5DFDE76YRtZylC4QY8K
eLC7qWGkLygPFJxgkrWBr8ZsEogCAEcV09ACpfjnTyc+JO/B/3Qq10SzODiAi3Bahcr/XCmEXz2R
SQKM4wL68XNSQtDpLPAnSadJSjPT1AiELMDjlYOtaS+16/wsk/efQtPp2DmjWORs0OwvfIUgHlZb
uswTBOmGRv9q45YiYSOhbhBeahqvNe/p3Plu2iJPiFpJeE9rscwU9LmlhrNJIMVTJhwSEJrO7pDg
n2xxA80nkKLVQqd5MKSe+pAaMtcgVUkku1gYXFnBTbNCmTS+76RLX38tMmzJ7N6MIBy3cJNvnzxx
bII7q0j51Usx37SSIOamVwJqcm614PpMQe0Y+MdqYNh5zacEgqN8kqtH2prCdGueTsxcmV2DI1TX
yuMuxRpK/hOjKHFn7rw0o0DlYdt2GjViMldTF5at+/HBosAt980J0A8Lh95u2l50cBMrAdckLU7h
tg4DXZsWz/7qoMA3gd4NGb7i//7N7QG7E5hYcJcYX7AmHviTz7CzZJFnQW5w1EQhNyfiUB80iB3H
vYRrfpV+IC0tX780Na8OlZtIOpBidebMklNjMKp4mB8LWS4UPuidJuWFPbSTDBmlsgVnUbs7JAYX
LminMH3H0XydzKxv4Pk7HvxqosiCrrEE1oiEYnMg7PDYYxtN4V01iaZZ+91iyx4HNm9IRZom9D76
NyhBb3OlpvQMmWqGzGS8mAK3hCRSBaok6mtqED1CP3YLmelbBpbtdP+3Z9kDZQHXyFmZ7tlMfOnz
V/DFggFpegreH7dOXSefNWMGP0MmGyFTGLPfPBVXZZQ8g8konIyTem6/iFhtWYiXv2o4I8XITSxt
8YMrkZkmtbxgIU2HHPHRybpA9/4jFu11qVK84n4PEG7OsuHL3RK1Q/XAkLZDcf7zM0ZUZMzJcwrm
daCLdz2oOZhpLILCDhwvhow9MAbzrsgYB2/Ex7pL/5RBITZpiAUGVtomWIvjKtttLEexUGoIwV5P
Uv74h0fnI/SQk7disybFBnsYn7gKT064iA50bWpCvCZHbmbkBLyKD18/4Gfh3Z+2U77+8zewH6m5
iRhprvRlecMRekkuklhqjhoRWbPPvIm+R8JlGwAdZ678ZyWqpbSWHiUo0FBt/DWOFDoPAjUeEOVI
qndczJel6hzCMx26d6v+VN8JfvToD5hYEN8vMV6iJ2fz5tzZPv7oUdHwn/57gLVV6zHLKeEdwaoj
EkwUIoKHT9iRkL2VlasESdllgfmQ4rKkPqCmw0M7Fzo+V7RKgk8Dbci2CQI8GlIcjK0Ya7Mj+OrV
50VknpVsYAkKwKsnLJZaMO3PoDvBWpR3EKTcvV+QyPbRvd+jWeKjQguVwAZRqivPj6nFsopbQx8n
QoCEWKmErcVgHE6LN0fSLe3+1L5wdFrCvHNLrkQhSWU1A4Zb1XxUSPp71E3N+AsirsKtafwFP7jp
i2RNAXh/fzKfn2k0Kd8RmJVVWO/N/E5ZyOHn7l0wuUKUcIrpzzORiAcJaoumriEl+Uk8iyZIn2GY
bnTxOUCAcK3qrNGmm050vrVPqoksCmIeQSiIqFHlv8Bi2aLfTtGtxXMSSyO8bkRDQwG3ThUj3gCN
X7kJMdA649EmpWofSnJE19YYBaFrX5ElvFzA6FsLgDc1WdZFAIyYUUrrEalz8Y9Gvni/oWi81WdY
N1Vnf7Fg4H6Lj/hW32HnKv2+YAtbDScUokB1+M7Rq4wC4jDqO2eE1R1fDABlg0MCflq0chebw5SK
xFFigcTg003fMBUVddqbRy5V0BrTI2f86vTKLyhu14ZEOiZtey7hGG9eM4xTUSPRAntaZP1Xs4b5
Lfi7ynQFPMhNIp0lw37XI8F9WPiRrOOcfFrX7KE76xIluwZldhzBVcZYfiT75rsJvJBl+Ip+njwN
JVFQvJQivbWwVOn5O3lzkrgyv3DZWWvFn4lSEo49hVN8ENaBErjb8CVkQUReN/IPdCtitNILM3+C
+S3mbEve4P6JVhvorZO6ID3CyBRKb53BF413E9mkCO3GQC9h5ELHKGKutFFrVxe5jR7/CUsqolQQ
G4KJF4utPl3LzwwXET5WpJZgjqAYqrhmP9jVILwmY457S9OplaWt4JaliOrqfDpesPwIypL6L4Dq
3jEO/0z3J4gZrwB+ju4CbKTK2x4QRkcrM2fUMj6v8MD2B4gsT0tejMjDjK2IbxpYiTWmPOlM1nvF
xtLtq1l8OMyFqVVCVH0E7dREIJZ7z0yDgonDX94+LeITjjyxeqNaGQsZCwVTn6fRRWzArGrluPOZ
t1aS1Rhz69999hdr/JRldYLzXpyPRAcfra6LtRwac9QvZJPFeZcGeQzWou2BBDu8jTwzkH3VqJa1
xPuEc9HFpkhEuObtOGgXfzX5czoQRUvhmhF//xhcurHj2lI5538lu0vNNx9DSf14O0bg5NTtApK5
vMbJiARuD2KGXsRazUbFTJzqXRcPcl3OkZ4BO9nEO/eBzKw5D50AOGEIm7CvSFJxrWvyt+MoB/7n
fftUD+ZuBlFp6eLUiDcxBlyY578dqImL11CI/8Dm5gsb1F6QOUIV3564bgYmp+KZfmSp5HKuhFDw
PijWTZtijlagd8ZmoB/6OE3sHdYZpU8H3fE45uB/cMQHUJg5hw/5oHiHuA8gGC9VxANClBo/8v8C
jF01c726RGifF408ernXTzOL+tABf3brvFgPbXnUQEt6aTiz1+AjiqicRwft3IzOsbDo/XpaQxBU
YD54SGEmXrAkqX8v41xDgyHauK2Fym+e2sKbUujvYUY39EBaDRIvd7FEDu1Dzm9DZ1Ag3Y1NVZbg
pV1pdWTe+R0pYPquG1nnkl+CS+snEoOb37CtT5nwCL2hO3C+NP0C3IHPqKqLcW6x+UKIkHUhZSBm
E9BsuEIsd+FNXRY4hp5zSGxLY44D8xSZxD+Fek6tR78fHLHLss1qaQLbdmlsvhsDKJkCd7cSa8Qu
NshwEuskibo4g7aHtDeNxXviJKLVK/OyUg9YWfb918s5ykZ3w82tCGE1UliW7FIeP1K5GSg3ZUfJ
+9IdZwznB2+oTMoZIKC+PfxBnI+ek9/xqQx5edfEYWgRyu2JolWMaXW9wdQiVD0RV9IBUWawVJx1
Uzp30c+UdzHKy2LZGjQbu3UqmdDHz6o8tWfkkBVdH0GtDivh6lljp6QRPI0IfE7/9RqaIve7EuB3
wDGP/EAjoqe68gnvAYs24RbEX0JsuOLTh+sdOY8G9JXo6TM6Dw2E1Km4OBNkeW77Vdpbx4Z1/xtw
kumx80QvW/g+p8lS5ptTGi8VD2ay5Bywjzp9AhJ4iMrl3MaCY6uZSdpNXYgyJWavUarOKMsTEULM
aQyfOnUG0K9cWYrhwk8b1tjXJrPCG7ChNkhHy2CC45PI4YIz9W3g8N3M/ltCkwUd0anq0eoLH1iB
PubhzCRT2ulW8+JmCKCmqmQiDokYGJN0Yl9Y38SJscSAtv9MYa+cNxYDMmql/QatAgovy7bBYxtN
SRY/bOErmHCOQBfPO4KBpNCeJF7gUvSiggvTL4oS9GJ/nTi/asn9iNArnATn/ZI+ivNZzUxpYBYo
WGi9bLtTGaptQxrGr2bbofdTX8fqfdH4wI4bJdWHD5iIZSZPO7BpU1OInDc4Kd/X0MGsYpvpeOnM
+NbLHxh74liAXYTVBXJmLDcMuRhoJ5D8bBr/KTvfqjXShvekpK5SEQGJEwtXNq/pfJ7h76hWqrze
Mo9BilozNdMPweQ9qM3tHegb0EGx7eOM6UF0PcT8p8eIr8VfKhN3FiOpiA18ZGc8pCOCfs3f8HNU
LW8SKKNFYhjhpWrUxGbzwWBuKuAvzBZGZ7PQ7W9VHQ0FkgplugxjIR0dPx8LQxkQv9RDX/GbDRPa
R3WAoa/2dahxq6YGV270NR5BoBEaq7paiKR42Qu1mkdaNj/dvja+zk7+fcrfV+6yrRv98g7N7cYc
M7FG4qf71bo0rWz9QJPxwwCUj20CIWYUTp9weG47zQCSbTt8gxbxzdIs0Gg5YT8I6km6WBvzjdfw
BSe5G5mJekozId61VEr2o2Q+SADqoLl6T/M5B0ezR3Wg9bHkg1ffRWblr4NB9/MXEtHOX+OdU08Q
31+hACcbSbGxiVnn1CcnJHgNruBu2iffbXTlLyA/UWU9bv7JQiVeSoktQUuZ52OYKVpWHg7l4+bp
RSPJ1fEJFbDbCMpt6veie9kziJfWJ8vjORoKLYGZNdiOz/HUVQg2lN0JlmD6IDzHf0xeTQs72fNW
FJ1T3WJaFKkRYvRaNNHuaNrtYUQZ+4diTTZ0tgZkThsrqCUUSqOTm2FRdiv9QUf8cYKeAuoVkrE2
3af+RunHq7E0B3u/cd3gsTfuALRiIdH5j8vOKvXowKMqq1uBFJjCPnwhwNoh5IJ533bXXjzkZHPB
Oimrk5Arjr3FInKw1Up2sf0XWRuFaDnslloXkxI1YlF9GXHlKQSjC0FJ0JsGg537rSK1IYVfqUvU
Lyr9W1ZghnW53c17X2W9QtwIilP+K/A1EpykIOYAshZzSDKp/Xs5rGhJCvroFZj0iEBVC/imWVFa
OgRCb5Qi11L/lZjG4nH0cBJtHKY2NFeMLO6lRMLElluLoVZ8OYhylvfFv3GJFdV7azikL1xU17lU
oZ/IxodnUnMjABxWWEyvyVIqNhcRKqgW/CF1fz3dbRNVp5hmJrY3vsWDW3qIYMk1cE8rKWyMFOvp
IyFcyhN1hGkkBH0k4FG7JZGld6MhjieXRosy1AZa5wFGiHoYw2e/aA+hONDJsh7fkrC70SAWSIY4
VPPSohfudK/3db1v4pZ1rZpwr5ldyvA9crjxAFJWNygmcKcxJS8LjtTSs4124whdxSY+AMoAYSUa
oEDgitMRCs6H4Syn0LO8skkQ1ItdT80R2jCmG7ew7T7zPm4sfgAtHfAuI1y+ncRNnPS270JbpXXf
eAAZ1q1h9DAI3a70ir0og8ImKveWfrXjVbdxuYQoIEtJG4LcXvYAybyLTwwAKtfiJ7Z6aChdY8sJ
bHTTAsAGAJ31EpK/SFq5tAee6ZFKQHBNfWynQZgyT3OlKAoFOhU2K9T0k1GKOzfRWHDjdJBu5YpU
Xehq5Fa/bfSFrs762ZCwH7T9gPb/ag4uAms8Bn+ElIr2/q2bRuFF+OwHDRBZOX4T5PIgwBEaxUxX
JjedHb5kIMmO+3a2c4XEnuOFsBZUTfE6dJTzLOLvqt46NS91YPily+j+q09VozkNjIKGW3PfyJkE
WsSrNGjFXQ7+Eai4heBhQydoY/1QDzsTILd8eedvkKO9vaOXp4ePV3i02QdvC8A9ZPmX1WTydI4a
dXgu58ztis0sgBjx/7w9+3U+/Ius2fObHDZMkPJLgLJNuHJuaTLqncuw4h/cwIB+6ie3ses7+SkQ
Fs2V+8TYR4ACGmDlquWHQiW40na8J6BNXxYG9pOKsNkf2rhcplXbi7HG0DO+fEyg7pvtnyQst4cm
4y82GUExDtYOOfrpnsVA/1dKl6G+GZjMRs07WP5sBQnm5KlTMp6MVAI7cLbyd8B4d7RhKe60cPu7
cukIgw3lAJfyTAnPf6v0sLnRXsJ412DwZN41DSm856BE91dpvs0Qqto92F/fpOy165MPSMMALb8B
MI3DG3xbb3rnogORk0SnjV5X+WNEBRpPUvLtQF02RAVDhaEyqRXxdB2IGN3vnwLK0oVAyeMBqLkf
hkq41WcWY89j692Gpbgw60/FRCch71Qava0SuabgYuJ611zi4o7OFDnNqOJ3tkSbrli8vKOJcjvP
7B88UFLSOsAiWBVhvnMhGRMs+p0qrXnJwvgM0LNDtltUizDuLksg8l6QR+HKHm3YaIO1gIllnipV
aOgqqJbJh6s4LktNJ2Jpmc/U4zeWS+iFVg1OLrJ8pE8lxunoJF2aEM4epq6r4xqnvT4SM4RGR8Vr
AVH4JCbktbgy4BPi6K62+X0R40O1NG/+s82NN+Zpi403PQTnzHInE+3dipgz09r/RifTizYvQvC+
onaXOQ9CWm0wUiAq4pKNuLmhv6w3VydIwWY/g2okx/mTJUaJHLhGAE9WSI+aV4TzsNnmcEsouj7U
be7mAq2dNAawdu51I7340Ndg6+fc32IGY0rtUbBRzqjb9imZWBaoby9xI8Yc3/CZFaAp550ay5f+
rDTyZjtR8BXj4fdYDEmY2vgtyQj++Wu2cyZ3ueFSJXk4NN5jAKS9cZIBJbbQ2pPdHAaalaLrPfMv
OidNCGDs+wJ74Whoyb6yQjXPshdTdnH5WvnwPQayMwGP4EQTew/uWcNVWqMd6Fv15BUZv7Zr5F6y
ReZHfqIZoB18wohRvnr7YsdPijH/++6T0WVn/yUXEl1WwWPKj6G93R1pvarXx/JykF1+FfTlSN0o
FPfV9PFzUnzPNj8cYgVoseI7M1N9iC4iz6OPIu0ZGfmiXIp2EBSFwWLJabRlSIDY6dBasi7hjXpL
tWE1+zfyPCcmZ6WfCsjiNeQPk0FlGfBHbVpeuzKip765dz1Zjx4idjaW3q7ZBhRPKPHpNLULY2Az
/HSnEuTp/huOu3+2pXyn/hqyRaHQlkwenXvT+QlVkBwYXxXnnxJ7+B9VkEuJPMogiv3Y4Wjvzd+M
Iet+9y+bXiyKvlZsHdCCvTkoXQh9rJsKQw2pa9l/cTwAZbWPTF9IMP1hazGEH/4phCG3v3de2qVB
FBcruUQgkkI+8kXIvmURu7Q03WKGW11824ROIKG9wg14VKZg+LF8ubUQH1yhuz6zEyk0ekqJMcdu
jLGGOKn661nJuXoo+dE59uUpqEpwBSW/Rzxk5R94WNKXk3XDT3LqldtUTseNKleN1nKqae2HiE/r
ytXjf1i5QAgRdrB04OF2t4NiTDWhfxFZlq5RVT6Eqm8Gd/PaD8Myc9cbbSiej2NeHuNiN3gqrtud
IHl4zUl/wbTt6GDwXPCTNFv88Ea23wBNCy5Jccv3MsDpCP8ewTxUgXr3O91X1rLy2dN/HlhOZB8C
8FKb6YBXaqBeIs/u1QLiJSVr9h+SbZeNiDKU8Mzmm4d+w2s6vZBmvqapXKFHP5n8A9jfZ0euZ9Bj
QvL0WPmV2e05X06wFUY9Z95qO6/GFwN3RjizTJ2rbBYfZaCYWh9XIF8CPei4u/2a7jJQu69dx/rV
rTBagXt9jvNJjt5UM746kZAfnJb4chvIGdV27m3aixxs3q3Me6OxIJ9MsgsiHeaDaHc0gyElN8zf
a9X59uhd3ey+1Ev/Brme19gaXgxqKZyL16W6jZr/ilbELw3a1IRWLbSWv5Tw0xTVHLUB+Ou6iG8+
2S3uM2SbbBr8ipdKe5TW9sddyuqaYNGGzGFatWT5cz4JRvTgPWtFAFCXQsuKtFLt4Ae+DONrfnqw
2vMScHX3CjKJm9Lq8qKoQFIl8ejfsqJmPYKWCioihn1KzobY684TxVtKAXE6BmKyn3iFAkNSP3lm
1CBXMobEaTZIvyviu4zlAzyRJnMuYHLt7Gy5VAI7wUFu68Yek9lAhl7amE+tPz9C8JlLmryYcGZz
GxHQP3JNg7Fp35FN9Jpg1HwYxjsyk209ape1ZpS2y4Cr1+TXfTGshh/7RMcMECFwnvGVVUxGXKjl
kB4hAVZ9bJp/F6uI+vNsJOvc9m+pgRN1abAKUFSWP6vLo9rjs7p1W90P+TK1ajfRjfu5h6wZbMJa
ZOO77e5FeUgzo2atf4n9VX7axvHbUrrg3M30GEXIc2m3r+bqJzBlbl1J9WBdZToRjOQiuqzQrbIC
wUOTeH1Y4ANFvifm5rDcZfsmwg/iE+feyPubVUBpe81vIdg7qUOh3n1/NGXnyKTEq/NsZy7qiLEH
xvR31uJmitr1mfmKfXrQFu0pB/ZH5mfTNRwBj96rRpRwxSpMnSBtyzPPCTBGtgwIEwTSHqNTfVQJ
3VlhSqcyeU4mgaSMmnyq3Cn6l5Ggi5jE/Wzh7ql6lfoM95ich9gtSJu9aw3H0ZqA6rBJ6sxIC1BB
/jiyLuq6RI0ru4LpS3G407FHW03H6VbrdH19wdFBx0Mgqb5f9To/wWH2+xV3P5yA5KKSgWpC1RBg
Aeln0XPyNtmZqANNNW3ez5u0+aAKX7nBh/ekhjvG1qplDdK1Cpd+h9bCsCsYovrTa4MSpfnpGeKz
XxA0blW5tydMgJBa9tAt2YO2s23UUAVMVNO7XkgsFpPBWuhF8cfs8i/trL2lc6acbSBQqDcLzRWk
ufZC0TgY97bXuB7WQkXvF3QC1Ofq43aDTzDbHCZEoGlXRLdzpSN/890i0AHTjchZf/gnx0PHwtaC
QWoCXdkjd6GR0Jq0FP7CnVi8/h1Wk9aXlp2PX8+G9sInYe3euuYj4GQIk8alqJjkxnjDegHWG8/6
bOQ0gn5qCtZ+dpVIuha5RP/Mwufm4/VQJjvXqup0iatKc+AnHQlZiQHXeTu1XlAZ3BPgnagB83Cz
X2ce8lAZ2LRJcQjMqcn4EdopyRu4re+RPCkqMMmWhhK4ggcLiVkv/nnLeEw7QsJK9sfNBcGIzz0z
28pknRYLMKb5Csxn6l9oelxV9P8hWi1zrNyzHrK55B3phL9sOooIxl4PslcpKtuDEg8uKvRpZe61
/MpECbsKZfZn7mo349TgxYn2Li4QNI0Ovw6tj2vrq8QWiF2Qhp1vwTCMcRW7Us9mJaRcKWjSyfD4
n/B/Ov7aJDbt2O/WA5iyI/JKgx32ngL6h+HcaJ4EUMC+51x+/brPJrMgvGFiHhLx5C3IbT4MgL49
fNyzU8JXjttmBCvSy6N+srdmsdscoyzBUpjmweMhVPVzN8I81rwFaaTZL9XzxUigoJq63kMiIaor
PJr9BEUVYnTwXxC7D2MPiKXONIKWS9pjxzycSCTXOjvXcVzdlq0oT5lLuLqoePn46uDAuebD1LKt
WJC+uufperSdy9BVvAn1dF8AY9oGA0KNziFKtXd/W1BBfxd7DKiuKK3sIlTA6g0sKZhHp+V5zAHu
vprHGWRzFQ/AO9T7q17gs9tQIG8vTXslp/86DmBbdU/5dMQer/k4qVf5qSRB6CrV9PvYRmnpDBCs
CTpalBx+e4e8FUTTwv8gT5f5IB2G1S5xwFIQBtrrRKFImIC8xy9fLF5BAfO3Txln5ktDxio/dtvo
PVdDGJ1KlhkAzwEyjltsUY4vigLlxjIjJitrfJYSbhrE+CPwqbVC97ninK1bDtADb+inbd3+bRkK
HqgznQeBzyXrXXNi48hjZQ+xFXOCIyoaU4K3RKxkEFLF1TW4eCoMeE5Xre3Nn9q+LheGTJaPv84B
+dGO4kveUn4pwVzcoNbwKQvm/Xg3hJeuQfNzOp4kSMYX7CVooq0XjBUbi3+wqImg2CJPbkizwqAT
lqgsRJWgNNqR0sNGg7iMWIL/Og87yEDHguNkq2QywMACS2GySqIcswfJb9ltbT14+4/8YsJx9XIS
I9KOJMnySnziMy+sixfRVdyEZ/+0775sa2ouU/MnpNNOqFmLOzcNRbEQrvsy7qzyEnvV8k9JTLCP
y0yde8UnEuWgtHS+bZzTZDfMteWOStuV1AX9/t011x5I5Umb0PHrAdCDaigQ2oRJ0ejQ05xDMIBh
GEhM7ZXAzCZQhPQwYmeWRCB+njlIxgbwq88k8YisC/4MGBXXhAUqj49VCqqXngj9+miU3fw9JlqZ
jC0Itbj+XrjCwMwDQhSZOnIKGIuUiMiJirWK/C5fGaps7/NDi0MFkPGJl/iZN0FRLJseV7L1ipGc
RwGFFY04vU2Qcad7F/Rz/2xeJdHHY3jqpiXODl1ktI2snmPomqwSNlwkksmyDDFkpIFnw/Q0MFH2
kf3E0uN3NUP3vHROl4+j3hVVuR60L4KU1PVLUn+4u27xITNOeGfE4w2dklKBfDyrne1hHbpZtY3B
SeWxasq5FhyIc0+6rYd9qYHldjfByYeGpazIwawpGgX7f2MUPtIoD2KCf/uYtJe7ULtJWra5jPZI
dTFTKuR8oUCFlaipzTMpQKaHOtRQSFRrxTJFuss6VkIpuEjAItmRnN0+Y3QB4RH9K0tG7l1vr3rX
YV7LD2GXQrNEAgbPzbUJ5OBhXD6NnJ1wRgRh+nZBW7Y4np5hhmnvhDf0RznYdD9i3DbJ7Re/zK62
y31CKUugcvkS9p8EJSl/rKPgrmv25ftp+TOMOv5KCjFIJu3Hv9z5nSvvQhmPtc5ErSFftdvhc3Am
RM+5RAp2xrqKMlo8HEpFEaqNQ3sL2YfzTscE4+XrzO2c6w8LTky6yeonG/NVt8179wQkd1Ws5DjY
3dvBUwhGE9hzFLYHRyh/M4TR8zTMIuLU97rq0N979MU2vaSLq2Mrhe/jhK6bJzlJTXI34Gi87K1m
rG2LleP8eF2P8io6nyM6vFh6yxgHfds1aqc/IGvvxYBspcb3ucbiZY9U1TvwLzAN6CtKoSv41+z7
VRO+fkw2jY7O1J+Pz+UQKRDSF7Ws/PvZpxtEoj+CNKRneIm5jsGe2Xwau3FbLW0hzoplbMXUK9/J
J1dEnqW0Wj3EedcML/kHPzLAWoMxwHjQKxSFQIS9Ie57ewmCw9KvZ95kGRPKs3koE/dt1/9sbdgk
Z4EScdRoOmZz3LzQlzU+5p2eFqyupavgjxm1e2jdgf8Hj+uT9h35TJhCtwuZ5ilTd6QMhGfDwwci
k57xAGhTZOyQECmc9DUab6XfJtDivB2E4cvOueQ8tBkJSg+pGeGKQ8eaUATCYCBcBYrRjm6Fjnam
9uneillehWR4BVMPaMW8CStiF702P3zImBjUyriT7ohyr8g6WvoP+SRnrZ2BTjUN6T72KaKwo4ne
9vs5u3K0rP3E30DxT192kswDlEyQP6p8NV4g1SXE003D8VXv1Kki2xaFixWyHwUKYSnNG4XxFxBe
35zz9tG6G4W+r0M4voS0INLH2LHk1kDVDzskhtJbJHUGK/BQ/ize52jJIj+LRwXNdeUqVE9jFgPA
pcZ6EuQzuC6RAqOidg7+Is62gFLYgU4nZ4xZ1FCNXDoDB2RspTqU9VPtgbD8FM5nq2VZTE7f9P1D
3sqMPlZfKBNWqYTxAI85FIummmdVM8U2pVNCOIBOlqJ27EXNBf/idtGSsaz465wBTxeEf6aO61dT
MYAE/8g0paarROPcssx9AX1SNYXw37e4kbKxZP3iEOKCTDoJDp0iryvk9HR0JMIQV/Fh/C3mEPux
7ydb6gDA8+s0D6/Zt13x1GpI2RSFgkj78Jq6L/+GK30fHqYyV75muvAJCZRM30J6P2YNUIZ7Xi9h
BMMEWJJJZJVDovBHaZywrNwOTIYci7eajDsg7yPulbTnhEoxkeX7/iWyPamBrPqunyiMtxMQTgpt
gvFB/iRWWDjayq0ezjhI2BScLQ0Hji6ePJ5MoMlFm4+54LCokVLsohJPAH29s78fJUXynTX++8sm
iv4w6k/115owp9ebNkxLPb1mW0zoDzLhqPMUxeFixkCjKFWc8+VifpR090wcQxbaYS8FpxTs0i3P
IYultQjXEMyRUuLZGpmAdP7K4WQ8FUrU9k3B7tY6dBXPcAI25hLD0jbAEsukvATRGMZBwhBVVLif
hSr/0nbKVzbYJ+y+p7PuX3k3sE/YRvN+Is7d92GgTfj5jEH/msgPIpDdbkqY0aQBc/I0K3Y+R19t
aJcPV6hKr2hIyHedpiM/NqzCixvrltPbIkxbokfhDzNTIsfspJYCoR9T79hg7AxIBY6CzeVj5lrs
12R95Esh7aDAM3XmGOCiME4ScjmXRBaxOEtYvyNOAtLyeDejOBFLySPDZruapoJTLOt/b1AA/fP/
sg4DXPexOyuszP+7YsrOhVPZNVElR4evLDhXxRb8WVK0pYIqqt3VDQfFKPsgHg4NXfpXGosvsObK
mDCsYHN2U0fIJtxMxnqXW3ExVcjG+HnhFaoqVD8xJNrQrZ00JPeGDmLw6Lof+V46aotdOw0R4CgN
SFit/uq6q6NxUSMl0U6sf2yEWfwt/pnpJKPxfmng99uMfM8DEIVzcaB52Wm8ZsY8uIxzGCF/NoD4
p/KaZsfUNB5ndPRKGmkcfkhVN8iHxIdRsHfqdGf1JX7fbN6ZVoiH31x0Py8v+VRBcHhLFY0oNAwr
Q+Yig8WhjaFqyvNvfVGlEyAGuiYC0MGKOdDui9mx3VfREG0kVgLOPdXJ1ETH6hflvf71WVMekyu0
g3yd95qjqoaRA3tb5vtqJQKs1M9AZxZU5aMGutAPub0dy+INoR5o/hJchYCfS+uBaHBsHImlgfYE
941nJICB+97KdhUOs10PlvDnymTBybdI+BADVT7+kuyZNj9hm91eYkrR6FPZkliw3BOcg7V1g4yb
EuttNPhVqUqSiAJvP76XY9M7H57IqKjdk7eqkajfd33/3HofHSNIQ7z3CVhzcWx2ZHlpsNg9ey6A
HWX7KcP7ciGjEwKAkhTtoMJyPUTjqzCM6f7Lm4mkJX0LEgi+hF0jKxsJklRtTdMwQGlP6rdcfyir
mx2xmkl229VTifGdjh8zs2PDfyP+JBE1Dylz9R4xhrKCbHCL1x7uTrrnyqb77Z5IgDORUHdyA3Nh
/U7+ztZs4ih95vCNj2BexIdAco5bhePp9yPGXC6GijxPCsSuESSgxP+KZZRjaUDwonxAyOT6SpV1
9AZsx5lZVFB3WotryyNKAC6Ct82wfDiuerW4VvpZHhedgGRmLe+YNx6OQB2gJi78Q6qrlP9kEaNl
pAn0NPRkd2+IpRkfyv+9skXQ0rb5PTKiLAosI30HcJz4TK4HNe8zV6XpXJ9+atVZJVlBzQ2ebvta
SBSJJxrhstOfzcTvGdhMXdbe0wkHKPlSPSamL8eUU35oDVeFK0FjrhGca4dAHSBaL5tkt4mmFb7T
BTojVbA6onj2ElJ6zHFtNH43DNPFXLHZIkzLFdQulc5GR+poFx8/2yTskMKpZyTGz7HJN8mHGDyQ
mh+pn/kHeXww37Z9E1zqr3PVQEYv5YyV0CowBFmWulHu1AWE1QpyEeD+xOCX1o/BGKxFW116RhNS
XUcI4Q6Ou7Kr8OVbGOVTSzSc7O9DotO29TkxeihwAEIEeR9zY7Gq6KdXxXidCLlvX1felzKKb5bB
zx5vFiE1mu6tBsZcimkWR1hW2HsVbsimMPjpf+2zFYaa7P93GLQ1oJDcvVcvFi1064jIMO3TJAmM
diGt0cEtFhkyoUvzm9vUko5jwT3gbg++sVFvJuJkdC8iLli2GSAEVuaxm1biya2KQR6bgh68CO+3
wHPKHeOIAUQKtRsMSE6x/8JTJqedVD5FLvb9TsnIYm6yGDFys5if8YiarGBaMJ9v+/Dw4kMuodG9
5DBki6kwFOS0MvIkLeuMpDvy6KMBKKc4kZx7ovBXK9Z0Ro57ku8B72djhZIYtlGzd5wuTYLIcxsL
I9M6DE1+m8SLYHFRCbpK0hZWINHAtdAb/c7Ew8/PynD2iDJ5Z8BJMQmBtPGqNOdhp6cC0p37j8Dl
KCHkbICa5RLXDVZIJeAAx7DiSuT2uAvG9l3dgIbWpE35fzxwBQyDVDO2+icecsAK94bsHn+VhrHQ
HpBCFTpFPvL5RX/QWGaD4jQ7AY2iNRytEnRQGIj8wRu6BVaW2ztJ/sT3St0Cl6zAZUCXTm/TWXQY
YbiOSNLLce0BvyPbuH5AyRvwptauOcZMdlkYn3Fi7zi1WkJ3nuPAm/BqxBbTfThlacSW5cdM0HNa
FzyAFG+WNNcxOF/plaoOfSGFQVEOF33yvE2qG1kkrEWGboZ7X4PFYhgpWZoz/inUbSk5jTv9vkQP
tucnWP+fouDIfkXwBFdwUW/jFxbOa/OWSZm9i6DD6EGHvCb3aIRQA6ArcHd0XA9SHaXTyehWK3Zf
YWWHGj0EHkiNAlWPzEaowzGcoKLsFZUjqcWxmSGY4CJqdjIHAUU+p4jcrpOQD6+1AxDtjE37mbI2
451pKWHk5YP43f9AKJlUz6FZjLgT8OfWes0CxUcn3bnklhhy0Puph4/ccnfkBrQSfVZsFdwWetuc
RBgGBH874M6mWj+sZB+vkzboe6uk0jG4bUsRtHROL+rlXy4ebpYv7aBUvVMDuLqixDa4fjrNA7X/
GfgnFK8F469+vfpjq38HWddz5baKdjHfw2bc1NTUwPd/UOFq3VaHg+cX/igxRnW2BM7OPyk99nVa
3mzmr1V07JnuEG9zcDSDSHzHT8e/3gTzehztHkmU9ZiELQBEE9rSxuoUIHogmWBpah0dXZbNeNdt
iUZLFvoZ/Tez1ocRkE31UrD/y/VPpVFdv66Q7tJ9HV60AtXW7RYbWLQIhSFv1cRnulMos/31dJQh
Hj6pT9wkB5gpC0NqhNiJGVbVSN71YfsaeKg6cLeJoxQIQ/S1BLUhXED6/7Jq53xwR/qQfZ07j33y
eyf73acj3bEVei+fCsk8LJow7UrPSMHQgffxUPZ/UVB8tHN6YoJi96/sL47yCDbStG6A5P+NSZGU
uJo5eZr6WGyP9KtTHE5u1h9auvP0VCcfotEkDW5+a+/ALymH+KPxDI7I9S+ZFVkVMGap0+m7694D
9wVGSM7qGp+CW3PEf6wqMzsVGk+eCoq8QBpt1YYACGBi6pNy2HB/BuCh6X5OPYvxciTKROkqKxFX
1TU1NHlNysJmv/+1V0mo17TzNx2Nzfz0vDEQttp4JoYPb6RvJz2k0AfTR74eFnQZLPynl2+YiZHO
JGHgfGNKaLJNQIYenbVWrjWMbvKFxX2dQr26la/TGa/M03eECQC/ZVlWjgDAsoxl6FsPIGTwBxQA
V1vMabttldTcXv//fPQ/nKgL7oLrqoBaIjD0DIetjPmSlJFJjEM+5gUUybGvty2D6ocUvDVLejuQ
YxkiiHv512HiILCfj1wYd0HqtA7Sw/QWDeHUfnfFY8IcCrhGZy8CeH+88kTyBYg39DDRcHAWpuYI
o6C4QagRAnxbbCOHpPQs5WsdE/3uxkIWyDyYDZnmI5hAT0acqmhtYyOINDuQC9zvZFT9shV5r9Uc
NlWRflB/1oxYexdINjpf745K7PIERP4DPJCP3ws3Rj+qaebW8flqthx9P8fBuYcZkpEwwBYUxS9L
FweG21KnkYwM/e5t/WyWjVPh2JS5fgPSDYmFW8rc7/LSQGN8D98nS+thzApcFyPA3cXLYr4qCS5s
nNppijbSTjq7ply8BTXpImqYgLp2sNbq2UGeI3OjSwlgH6740+1fwqyAqzGaUReOIHkDV/M3lDUh
nU0U0WUZSmTE7R9Muyb6JFSSRYi8UPKJyFQKTC4Zn92mu4WbVG9tDiIF6mhUBt33FopnOfclkwfo
5SfXqU14wHzYuMxSg20kUfQMtHhtzp8XZh33bLHjRCklfgXFtCd0cGUGEIEhc39g5PxoaWg0TNYm
htdsL/qMd8ZlOP3B0CbFeMOZF1FRBDsJIJdxYa11Qt6X9/FKxo+QjfRuhAoO0rrBzu0mFtIySI/9
ZtoW23Iho8AVyUZfCI/cvDSk3LO9nRXpgZTsIsy6ZpwGsN0lJmLaqDHFnLuCxOqEb1kPcXuT6WJm
IwiFvDm7mbDjocwbRl3OshvvxIcyDGS+EiBKc5ugrjfAyCVbLkGhJpFtYh9/U8jx86+fzA8rXxhP
3YFzM8RIas5xHuuMEuVOo63uJ1hzgIpOWSSIrPCGrjmAWqhQqj4ISipWT6f0zovPNyCJ40XUxvxL
WAtNKNKoiDBFwYrf9r+HLK4L6LYMNlu1fh8iDgAuEUsO1h7P3E+BvUH+lbgnW/Qw8hOEIEAkDekE
lrmDxWadWElPoZDwrubZOIC0NR2Poz667qxrKeR8QfgW8O7jNrnVoV2vaaZ+qdJ5EhhiAZHIooSL
i5nI3siRBu7pp3SIVTTfQ7LznxXtX2xpvUaiHHCDWmAD7keBniplykRk+TWnlvQfkOIzEnQOISAB
H9u2Tk/kdMGNtyRTYO9LVQ/D0/PhlndLSNsRtR55NlzPimEWv829j0FsShC8oD1HhQot4Pdr1AJa
e+CYMbzRKYEB5nIt5q+tQLfsaSC6fuwEUzihDAQgI6gTlcGQKBJDq80+3qpEk9+ec76bQq/eg7JK
a72iVnRrnin3+I+YdMbZIZOGwYY2m4O8d7cRABzvF6EUCd2DL6k63J1kXrAoCFmjCdnK7F3iq54u
RDtBJ+VGKnD4lmrzcWxVTCZFNJKtfMUS0SrWDeMDNkvaIeFZLQeKo+HOJtHaM0KpknzYX/xEBwTs
/63oSsHXFAZOUXzzEEHSsX/Hg2fknNxcw8UgK3XBpgsZ3FujRhCMYPUD77clbaEkW9K6PUEDiTCT
iWmeuyVx2HDXottYZOkNtGGl8I2/+TFiUJj4G4G30JjmcocbnwDU0mHclNz3iKOAe4rVMetk020G
mqr6aaSFbDQG0AtcxTfIBYmZBiwlDMhETZZEU9s1TqAlHUQ3E2Uh/DaGU7kF5sefagT/cQvVHxiW
nUQ9+QOcAGhnFOEEeJUqybZCj+LY/P1L/Uk4M3lG15fibp2rSf81ISPZRLu5zsUZFQJAOkate6U2
OorGn9LXEqyBhgf1c0VKq36Dplg0U05Fv0lBIehdeL65pcDQflBG6K0KtlcdDvVpbJQ/fXnLRLoc
atTMY/9kHUHqRuf3TfmbcvrAnLwdzgoYW+DEDmGjejfngZrxcxBdbHSdysLqTQtTGLBX6jgCEcRx
FuIhqg/i6VaD+gzEimGtjCY1vx/KTepf1Iu4ohEGrXDadb8ps1wdTQd55H7HAStrE3340eD4le0Q
w/zSpzhW586sDFl25ebhC0MU2Jiw64pBa2Ds1DVqzFnycP0Hd4wnBzJQbFowFKqeCniBpkGAP7fW
uKSFsfVXROv2vjgf+lBBox4kQyimlZKHEOmN+AtCDs4S5+rlNCEZPaejThOsFGVSN7eeHlS8KIAL
OZ9QODPQ7vF90yv3Is/NCxDo8a5JeozCVdST7+YBmYboeLwdE2DFiJAhqeD2u00IYMQN03uB/c9R
fUysOs2e2N7fvfvXsrVkoP126VQqz38s1ZzNjPGcnEsaUPyHJ3508CzbrpqcipvvviuevCNrqp5W
W5fAnAcQCzjRGgYbpJhyaN9mGnjAtQzgQ4W4Qi2lfKbTtTk7y3z7LHumzPHuoDnvs5JDWzSTBngX
hEa981vG0Y0AeX4EMhdRoibDmdknTj3HWaKFmBowUwy/CIQJ8gb952qf4t2Mp9MtK93IirVv2r9Q
TCkPv3F5Q3VpMQEN5Ym+zQbJK32GmaUt+qVAY0XBNXBDyMKtmGnRcsJIJnf5AB3H4eW+4Wrc7wmN
CG/dif7He1Ec3y9EYlqMYzEqhxc8hvPKY300Nm8LkFCk4NlZyQ6OxopTVkJ/qURZUlpJtBcRjglz
66q01dXOvR2NK+OgzZ/deNGRfiPiFeNxRiGvD7M7N8sqTse3+iW1bVPRX00+n3NAXfJ9bEZvtNDN
Jh6/tPe61gFcE3Pm/zInwySVki4BzP8RVJcrfJP6VeLTzBg3+c7rQbBTwNpcyBn6qbq1yOlcr1nD
hmIfiGQDPM4ixQDe47AvYhvf9qzcaXvtPs4zj/AuhroHX4Q/bzpHrqZ6rdpdL3cF7zTStpnYjl+L
w8jk2tYfMVrN3ht4W/tz5cNePX0qz2NCJ4fasZR83s2zB1XIiRjBXFo91lcnsPQatodNb9VwM1xZ
rbOzHqqAL5Vna02GCCMX1t5zh1RcNsYQnMkUzUNVJ6G3hRMfEZGphwlaMKo+ZAmRtER+p1rcj9rl
gwvLFrxTp8v7AdRKn9H/fh9PIpHFyN9Ido3lXPPmOPVhu9t6lKh8D9HxhON6XzSszoKg1SmA+Jf0
UNSWb9Ht5Qafrw9oJwrVZVyc+rFUF3p24OFdmBTBPJtP10TnuB/vqdFcvLrINA6JNJyY4y4OxI4C
kRU0Z7GEorIWiBL0V4rrW17Rc+HFaIK/6ksbMV20QWHz4GKPziE6asdxJ+cUF0I4t44/lILnQYp1
uvCJ8R5jThZ0nx2IDdmzsM4xfrrGvJHtCa8fMkqlB3pVBmynGb2dqhFzGRgQ+kiG/yt3io+fLQ5F
m5NYKzdxBg8Zysr7rZHYGCEZ958sswuSC2be8bR8YOZEnX6UEReqstosiy5naZVY3/Pl/0UZbkpZ
dmXQidtUvBELXWThkQ2V0NrLSDqdIhX6rEt0l8Wjm7b5ONM7fY18hkzwtMfm5Un4MMBR6PkHVy4T
leLGwNFgq5zMXKiPYRRXQJlw2sy7MgSOkFcA4vQPUjNDBWpPaZc/NfkMGPX7lhynin8Dh4W1Ozo8
/UxNWTwTenlR+QSHBCOblEZ4CrYxirSQIa5afn7o4paT65pdEMW/yGPiVHsK19WIaiRigXjmkfEL
8QYCZ5Fwjft0jVn6o2sZIKnRq9xLJn95cj6dHYXHcwFVomJMkYU2Xp9VP4YhYsOYDoEJLYZFgzoR
L1WhkdpXD32UgGmaWI2K3Nv+SJuB2RBoaUS1c8z1auro9wTHaZuaqcKJ8UVsbqBEjYxmMrqSvPqN
H2H77gEVnr7tVo5D3rHiljnmXUqibV5/ooOBZznHalK9UWvnLbJPswaeZfxmmV2kohOlqEz1NjyZ
BhmAGUFR+83eWek10oGiZdAH0Cs+j1G4zcRcaxubTdMHxlYGnGrU6U1YR3p7eEniY5NOl4mfVtuC
zVLjovGSHMsQZUmjBPflCVL8+nZAY3R9mWATaMEfdO4hXYfzmWoo33KwllZNqaFj3/iCucrQTi0l
AlF8TjGX4UYxt3ZhwuHPt/VXvO0g5lsQ0upwTgLd3U1x3l10IJLQ3wgkv5gdKcLRCqxvEICNJHCU
o/8OkKKRxjaKyTt/mcs4Ot3vRfATCwxokoLTzzOz3LMb+wdVPsyrt4WShphje3S8VCICdaHg/w5T
bb/BrLVIom3vzBYaVqVOCsHnrarcy0xcC6Hu8eSgt9kituK+ivVOWsK7BCS64+/nSwhzo35o5Uby
uOVCxrSLf4KgHDrx6eK7Y7fnHkrTNmokaOj/5rqSEthpQOc0yJJUOoLNoIGoMSF/+6TlolXd6/DQ
WudasQly1IXyGXVC/oazcc7+jLga1zlVZGobeOv4tVHbmYC4g2Oli8Hn3pp8y3ca9d+JnooaFZ2k
VfZZaELVtDmsp7r6qUJvZNff11l70lGMHQhaXWbhomRtwPcgfXqJzh2CJ0Omri0nR3fG1jTfUYtG
waq5sxKiV+PPa1a3FDXrCRDP/PBosIYilgRm+up4CfkHCGDY32fU4TYeDb4s0gKh6z4wp6lPdthW
1FM9JHe78verTXgf+kayt6ct96nbylpJoiVKKcQMFmYODgGZJc9L9Gy3CyGvhyeEwc4fglatZY4E
+OKHLqjDo6a0OwuSdxZ1vjhy/VF3w/ZaM1Pl7JCM5mxsOWOHKrkBuQ6MJ6rq4FgnvqNPiC//bmV+
aHkRmFccWRcCRNYKfSNx9pR8nOvDVZUzuM8BKPfrfUzon1MY7q9v+GDFQPry2O3DRuCB05bUiZmO
xNB0qhz5BNLbmV5xBlID1pXZGrYJIYirez7SmOQoAfIIxLIIp1P+TDsV8bbNBRHbHGhjg1PkeviG
JvoPdudi5iAmzvGKv+DY3Ohw5WoYEIBptAhe//Wbf/2DuorcVUkWhDhhOinvemp57zTG5BbYL7T3
ByU102AX26I+AqMYBBtEdIrxTzW5srkXmIV+15AhdueAuHQYeJq2+hrdz4Qn/uD7zi8Dk+BOl1Fc
8XvHcusvgEHlS6dcAijXIl5+UYLbcvfcNjrAcaKkbhcIWaUg0BjkyK10Fow5Iv8sYqz/F1mSl4qm
uhoYj1aXWKR/Eit0TtQGYP/HWG3KEuO9s49Fy83S5pwHaYggVnwovbdUXOn6gufup+33IZt/ViMf
gUTUcPeGwcLfy0VICW3n5OfnYknTrlXbhie8/3u7kS3H7t/eawKn67mPVR4c9KzMUWs/coj/lTID
91PPk2uuDB3oguK5bdyt/C46xQ/zRA41zy6NJ2hkiVUQBXMYSPqRycilhQI4bREY0tsOV1rLv7AN
XialmJjwkmthalDQX8B5QnDH6io5YA7kR3j46+gMhPjahh8HmjYD+MWaizrAXxqJbkRDfW++1M4d
rcYtwRhbGFdEWB12d8mYyxnp4S7aDKPH6vW9nffZbfX1K+IbZXGeILHeNFpoExTvUHHkar7GVdIV
fMCwwr+FguOZujeNUpfh4ktFBc2wZGmdF+9Jm3d+QIGlIcqbgV6om2YnGP0FwzfT9tnkjCkBFfC+
3cmHr3sNIyzxDruJ45lmn1B45XITL0xjkD3BgF1yuQcIqqIWefVvWQxOk8gUdj/+OmI2D//KlOJR
ljJMcKl08j+otmsUFQnRHKiToOth6+TJBcQ6IC5c6IFgDZKl2vajurHVR+qmXOuaRcutwB462Y2O
pFCgeaZPGZ3tC1Gg880gUt8zGNsDfmfad5qCaqVcrZunpykjSUwJC/CpjcagXjf9CqyaD+TrdeI3
ml4teicZUzuOSvgDNEBP5IelRe9foQ6GfQmNop27vGGJ7I++382M748KNlq/A1a+wCon4ngfNaqL
CxXuUiLxfemkAgKRA57RJ49P8L24dDGEYCeq8hP+kwrEOqEFNzRPgtY05updwYqE94Witg4rica9
VCgePSqPNi2GGHtNuuVBDvBMmIkEi0VkdroxH0NBxtINi44NVftSxvjvvdyR15J/Q0Z5FAP0Axby
oV2Ve8QazA7uTzajmGuxCykzkF0/7KOeQpWO3C14ukDvk02wRh3j13W3SRw1awWkvKB2uzKv88E7
joAWOq7JCqRLDFdtXsgTVWOUKrlOsn1T8mDpW1g6T1CJbYO08Uw3Ukrdy+nYR4YsiKqgsfidcXGR
8v6/rPVJ7AviC7QrZuR0KGOAhkUX8Ns+hUOdmRflHp2+fqchsUdTHjAbd74Q9mXCCoJA9+xiE9e9
itZsbfcK8ALYXhCrFwbKljuLIxH8rn3WTlW/qw0NamrEnB2uEv/JjvbwrNLh02b2bI1Qxpz31qQb
1AepiFOxqa6scOPTOx78ZlK163mlWu7tjAwOBi1MH1ZF/5DczIxHEJW3IHn307WYKbBIgCFHEtTh
JvlpIl+WJPtcKpVfEauw1CVE55Vb2NQOaP3UJ0lLQ76tiPDW82R4xgiLim7XJHDsrnrqFtCqIVQy
xtzAFnQzeXkfF8kvudHGP+i0dgI7qsxNyTibLAXPz4sapVDejYcKUaZI31/JoKcBlVsfF7IG6svl
J81GX0NMgU49BbxcPYRb8yKE/D0zm52E1aRMNS6+6dxTssC9Lua9Eb72zfS4ZTJgaOXgnqALc80s
dueb+tiuTvuc1CKDGFfo8BLBJ5wI2X8GZzWFwBHDUcWWpX61DlPIQY6ugNdgU+S1ZKFlCb9K46EE
toRvzTcPv8MVwP8JHfvq8w/0YHN4CkC82uJqxb/3h/amC2QycoRE2glqQBS7xPhM3v+CTlb93Kn7
HHHUVn41XuNFSmYyUlU633xjuPwjWvCvm06odcHmardBKqEiLgIZqfarmkEO23/FFPhproxlBBaO
yz7iC1KN5BL30E4wKOw+jwj/p2ydVNUfggViOAJt1AFx6W/qkwNKFOr+J06dk5+4GhZ3x1VfMYIK
fSHQiUhTZC9BGftYwGnLT+iYT4YNqBK2umPVy+0M207j0fmLaVZK67bo6O+jg5NdpF6M71jeMOBs
8pK+ml+HiapctQb6RD+xxm7XxZwBgOouWkRY71EevdzYetziUKKucPSJZHdVNQeN4Bae1XvUTBbP
a4T22X1G+k+4uQ9pk6zMm3e1+J7XvIdLbfEAtucPYvCCRDNMwTngeLP78nllSaDITgK5nKNalaC7
PBQnGPC5zwL4YxjnL1N8JrdIzHh1lADqki6I6nrmx35hpJYJ7Wxy3y8A6mdzwYU6oQ8EggJSIBrP
B0ifd87IjPEtyvuNNn+nhQkrAAO6Uk4VTDqm/9IGUvgolcq2/tooaMsatxpkD+V0AX6qRKpG1vge
JImL4YoPVsWlaNYo2npqlw9fAJQhs7gkfhdFab5yUmUyQNuqr5AUkleDf9MG+BVjE4Ly+sDnduHb
mFz6PjIonIDLCoEkeLsWCfZNYJ3lwj/R1uHZyp5zPMQL9vDa52DwVouSvdp/mn0pjzzgTbEA/yIE
S1v772oN4ybCm8d0qiG/ya/QMQnrT9FwXEXuYXUmCMK3f8S3S/I06PvWc5KbJqhGSm4oQTzbSpsY
RG8RqBTVkqBCFba2xmGI7TFfCjDHUD4DkZLuGLjdFGufDedZelLKHgxDRMgY4CgWMNAY6Vdy9Cyn
iSPQyn/XzrGvGJSC02H8tvffhRnxCWpbwNyifI1Qbz+guPY44t4kfVLGhhPzEjfHk1Y9LRZFI/p7
DzOl2ZZs/GXhfUAs5rNOvdJB3lpgtONIZ7ssHz1CHYTvvspXivNhqbbAiYeWkwKCRDbGYkJ7mbRZ
1Op/D4NjqTWN+AFxH9axJlecYEFe2ymZvhs9eCdC0ZQMLLvhfr0Bo1GQ/uVrrGyFvglOSvBGh86w
vZrZ/qo7e6Og8EJa/CVI3sKUOqVd2Ew2qvWRAuqY14jxeex+TqzACh406yCvEz3k/s29MbMaF7gG
oWkukXcEKVStY7R6VtHpvsoMXfwJ4Tf2VpwjbseO4QSpOfhGLSnvjJRz60xIGYZpUbBRfOAu3xdS
tkP8E94/2yMsnmcyNnu+FLaPvjyOu2lRIIWA5s3cewpwDz5aCaFSPPSyyN2cqBJjt7kUP2Dw+Zqt
v7J4Hgz0ic9eJ9m8Nx5FPE92tEGq/78CGJ7qPY9M4+2LZ1KeiDq6aW4AlSY82XFGO8z60MZYe97x
vsXuAIPhSM2ldHPyhBVW9cxGyk2kuhHCpGy4qMTDrRaOBCeqxrWxM7oNvhFEBwxo7EcW28Cs/+68
FSfJDf7Q0xOEApUAhtHbEFQd03yzfqu0P/7g/KmybTxsL4B8EwZMyHj+ONodTI9Ya3aPbPHMuMc3
+LhDlNI2ukt7AAt7rk0iAs3IoozYTNPDddtgi6no5924X5Pj7nQrER0hqoUike6bBwIkemcUV0mW
ZAkyo6Z0Hk0onJDjoF4ZEEt+6cWkPBY5/hvJdr9PYKMs5sYAIl+UWIMPfEbpFWnVePbdRLxhizNt
tEtu49OHL0hNO2UaZYh4tMf4tpGtGF+BGKT7RHpt6FVqV1sOirFD6GfGP1hEcTcgNOhBeZB1gdvX
A0ZZKocj4m8kcWWHvedPNifmBvpGxLWPnVQl6QXBpfxSKznBjE9eY62xfF5MiHymwWWvGgQ4MCPc
IA+hq/6jK0EsAhAgGCNB/lfjGYfbkUv6HwUeWNHYMWh2URnytJ8Lk7ZFT3tnRI+D6lIfVGbapKtu
eOiZCHzJFlCKKHFMRm3OYIWOsKKzxwa4CXu2HHNEw1/e8514kgR4YqVJ9ACdmDIzBsKwSf7zIKel
IOA+qAqMtVpIeOTPXDfyz03ZnBPy9/OECHqBBmRnaiWKRVGCVE2htkzPlR1x2Hp6Ghv39l99I2ff
MsM3AjkIxkDOyc9Y4NkQApwVDadT8X5r4qFHiRY7fTfM6/jircPQV1KoQ0tcztenHVL1QH5Dnt/M
IXLxs+d7mcgEcHDzC2vqb2GPtBbHdCgbHSeTGs5wRJVI6yZfDtuNZ8ttT4pR83yLyDrzfshTbuRG
AEpQtGvsGXBkVbyv/ZIktc8HMVJtPLxz3OSdKPzT48/Oqd7x4sVVNhL8AI1I4ivz6m2Ku9uwkKId
I+jdNdWRuEBE0TsW3TMr4eZyLSWi1Q8jVsA/ENN9bQixThVXW/z5TiKkIQXPCYta6+jYr8LsPDWa
9HEuTBGENHNYGc07dOQx9xGb/zXa3cMGLBdPbzEjIhA+VeSGoC6PXqjQv+qBnRNCaQRfOxvDq2YP
brgxZQFp4DEvbiiQ+OUXqTLQjtQan447T764ax2LThbofskA+qF45wacX2BTtMPtQHfYv1g5G3Ai
8OhNLonDa/nTuJruMSgnFlZEmQiJ1/skR6r+8LIQmL56jtk+C34k2lrkrYKT9zyKScgiGHjwHWqt
HMGuGXyLM6GxR0rwdZknYxlJiTCZ985oVqlTTLtJar/pm2GoEzu1OVXyIa4o9AfOOQZxTz44B+VM
qjB2ERp2D6YocIsimKnDzGgmzVCFYp8ZVy5Syg2FaU6TpRf4Do3Iea5NCCKov6krMflc7ZDmZGnT
Y4k6lcBg6ypPAT/3sCKK+QAP7wJW7munqZ/1PXvrHrKoqCQPAhabUryzG3/wqMH1oSENylbSlRUe
jh2bB2KNbygSUJLBAXs5hcvkfmegzpDKWvUutWXLvB/v0HmbYRPKmjteHOb60NYSsxDYccoCNyLu
MudscGJtPKTx9Y5HBhzOgKP27gyaQWAh9xxMughpIFg1g69V6+NXaYG7kdz3IU+KZzvIDoNPQ8ln
PtCY0hsvEqAdL/9BTYt37ZisIW8Cih2lDf9wMvQtK4kyjwYcjEy0KGSvKNqu6CZcZKBooN4wh6oU
Vh1R09tP4zdAJCvm20vU4BXwWasfmLtE9wTKeHQ1O34nyiR1AjzWSB2J+e+bYxcQdA84i1mXmtTF
b8iIN/bAYF/7DowemRXQqxJJGfJS+kD26tMFW0UvkVSWs1FAqMFywMoKJp48VuUA3IxwgrAfmsYu
RBnBrGm8w6S/e4LaBqGnMFwl76Si9O9CSk6EnhdTogBHEkLFd00EiSxvp5RrO/rTA0olHRAWF469
5lBtEsasZtcrWk5tp7XoOxsmi4MHxH/vJmO01nXKeKSVl3SSif/nQAtYDryDCf/or+XWtgJEzYcS
Dgvg2vbWW3YzfLF7FnhPVrkcjiwcR5sup4Kkakk3VXd1l0yy4OMAb/qZyLW2slG/t9M00xMdX28j
RP7uoIAtGqpLaz8Xz3ztDn6HmzLP0fIUo4jVlg+PtuPaCJInPwRHqpFrXcEFN/Ty05NGV5XBgJcx
9BlR3bgl/f7gqORBe5VMmS5Xwb1XqIZllKzuIHqQSsgnzejP2hMHs5t5jCqbRitJzgBNof9Mhmt9
I2lDbY2Aa+Mtf/BkmBc7Vbzk8nlNCEAxnMIsxZwxFCfbVY/bs03z9q8iR53/2NcKYG4WoKJIpRPO
mmdslkX+Au1xDOvqwOWiQ90gyEa7tiTgWpnQBJpTQblc6a8zJYu+uceh/sCKUfwuBD6ppn1BPFKC
YhNYfgcRSKQ2LOYP6tkKBGRDqCD1ZdEGGSv03RVfEWKRg1OnObeTss+Jde30UZJubRNeaFal77Cb
G1FGLOYDrU519LZeD+9MRZ7oaRDWZIHD90wJyX+NwdWzIMXhbXvNCUdK8RQjGjhHrYIDhA+Au+AY
b0Z8fTmlX+W2YC4a9lhwxFTgkRuf3Zc0YiIlnJyGTZ+yEpy+UXoWP4tE+qAad/JwQvDe4yD6RZkP
ogW6vO/iEarxHJ7TDL6lHH6nsgOR2lH64cJG2bq/Mk3XR+K3tKmsQHbMm/qsTGvcYq8S0YIQzt6O
ab/0Tl2g0lun2SrDRSR0cqZgcTWMN7cBYx2uBZqRylW3Zor3758WQhtflaPAotjnwiOh5gXT1m/9
esjNjLHwyeVzyz2v36rDlArkkvD0TGKJqTNRNpSRNq1CGVdRRg9QTR7R9aqGl2uua35JhIYbpJml
/O2UABAnhrOLWlrrGINkijIuCfX4yij7UQhJJ/vpV08R7JajtZqlheNPDIbKCUII+72SjY9S9M0F
36Y4ItsFw/MjZpe6PboxL/JhLlPIolIv+W+lQUjD6U1ArvOCnmEhhizHwzntM6jMkdZqd7l9xp7s
Ji84Hj7tm82MYiJXuCz6dXzwyOB6mols3ohL2fpsseUhKu50UiF8jRcfAoHL7owyYNhd7zZbCe99
Utj+7L0ErMfmvkezcLTogJVrTFIQaMDZgMU9Fi7zpR4TsqSszM/7J1jjaCu3hZ3qB+6ly2g+/Tu3
vbr1v/XtdhTO46tanVvpT3myMPnSbOeNqDMSiPEZTjZSmeNWleH6xiW1fPbFhXoajIhvMvkVfpI5
2/hGimm3++Rn6z97PTofshaE3501yHqKauXnloPo7u+sxzrRwfXTxNv6iUoXeXm13tV46kFhu660
NCzblGN0jrSbqnjfc74ZksBvasYEtBbJhJjEjZFbojHFHltJlpiOUKvlffmzmr+d0Lqs8rp2LnDn
D/NTLMmzjdudR5BHNyU6Pf3GetvoldbeHUFoz0LUx0EgQz7gdWr04IyfgU9WNk6Dfsut6ljsjkbK
SDW3Az552n3RSAeEvR5qNr8o/9wOcetaorEjwQgvFm1nFa+U5jhTm5Mq10bxHOYuHHq84LDPNvby
YikHoadxO1w47O01xrc+9QtfN0FDVIbCdhSNNUKgvP0O8AJ371lKT2hEBYeMLuPz945xtn7EasND
ofHgA5/e5frDFjMERPug2Hp911JrizCQ368aD7AxkkAeSzeQDpOGeXWmn2bij1f3/OoBTQUEpV8h
U+XLNGsdCuJQqrIg97I6G9DGToiA8Oev9qyQiHy4RHxcMSNA/N8zHWMFw5/aqozGoOFe4ZeoeqCg
VKJtvb3/hbte7bt5+Lig+EWo5W1SNIJaPN5BMfH5DOlV+odxtg3qHNqdRi/nxTeQ+dIANwvIi0s0
WjVHdj1GZKT167ZxP6tD1kCKYk2bR0iSUvjtUFioLycbb+0gReuRRFPA4Ebads+tQd0dylCuxf28
sSyy/TZ0X0lJGiDyZopYQVgT8VEHiYFUaYZrtoKn7NY9e3nKO2YyBJjABNy8seuH0KFDnJ6xmxVh
d7pfpkwxkMlSuR2G1HoLds+lmIwS7J2yE1eiGZeKnJjp81APgWDvhvXqndLywBHfBoki6J3/rXCh
rERUbwW7neD3dYLDRtxXyVFC72FKcpcrL/l/SVCzCLvCua0kQydCFtm0ULrMxceOHH7oGGpDjamD
4e58ZQim+mOVQuyO+cwkMV6LZ9Z6nPPsW9QN2AxUCRMQ06Dx5lRbacXu51EuUel86BxVQWNAe6UM
Hx9OTyO9TDqAor76WXw9zB6kSE3QAfXbslJpUtCQdM3/tzHHl3ahqyXxtXn3Y6UuRKZmQEBVEejK
IrGTlIBrSXhpl8Pd5QRd9CE5tWcfJ11lnUdCSmIIbyFCRR+odDXn9tNckqFlpybBprRfO8eERjMB
rR7kgWyOEgDcCEQTDdSY8oAIkAOYWqWevF62l2lE1m9NyVDuZbWq6d3GnU90IOkP6RwngEZcxh7o
BJMPvo+BtmFoDr2JFXRF87ttmIk743XubsMvO9kjVMtggGDW164D0zj44dWdhxWQOT8wSqOxz8tY
Q8BKFW0UY1I3O34LKw/QL3i5CJh9ItoIiGZpbhrZIQ/hqbWV0UYq2Tj/Y+QUstPEWDlpI6Ah/X45
Z890GUS2U3iocgkFnBAJLOc60LoFrzLnDO57CNe13puIKkFvl8bpxbkd1G/6/9dqdSitNGaJ8qw4
fqEC4kSasbQgrV24VGT14qO0tbKue2dP1Wb97tIXd70X6BBp2qpmmMtJmLXHwMQtGebUgLIFJ6Yp
iu4aHsXnSromZIvXlfWXHk1l1OW4gWlmyHacbszjndvqhOdhvxouOj/kxdAtgVUeb4gbv+M2a79Q
GLxSfFbYwyGJ0qYUJ652OITa10cEmeei4a6NE5Gf7zHoSSFmqkci08cjA7D4Y8d/t6kuPpq3pu+Q
7P0m/rIMdM6eTZGD1MF0lT5tnkLhe1jCwmpe7RJfH9awzvKAfhvyjMv+O1fMONG4vTXwutlNyonQ
U5i55Yle8Zn3x7A6NhW0kQzR0Y/r75UeAf8tP0FsWHxA9yx28jfjdk5XkyV2ww2ev5uc8vDy/MP4
xBUKYnUpD0t/hLVPtZmuOIguzwSB9s5iuWybnT9i/GcZQ8YK2V/eHjIkWPwrIjVVM7Vy6N/jKpZ6
x1nBUrXFVTNHK2N7T4kV4i0PheHLZWvfLol9deA/4F8F9a/0ZNGxPlKa1kuqesi8VwRUW57iv6eI
qwoh+NHOvwiyzPMRwCCAn0MEOEWijLuMhSiMZEZhbTxGP2TMNMcK42LfQrHCrYK+Z+VzLd3xhBIw
cZt2AjcOmk5ilxKe7XuJG9J1iiCStat1p2L+nLivUE+pYqt3QLXwl6iPoXjRCbnaEIXIOQ2kqc5W
VDtxGD0mZsjD2fRa2Av5TNr08EWTHlYtn5mKqjYvkQV06A6Taay08fSzUtdPG9UfhLkJryeL4lrp
KI3kRnPzRY7FEqwVYACumRLKQbV5bWRUqTzGuSm5ZTbQpCVa/988dRgg+k2h0mMUAP3VbvNnfqPj
sUCebvFCMeZ3iY341vtq5FmWHW60L8JxaBf/yeQnT5KFUKL2Xq0Y5WhIRzIErRviFltbeOLpXp6L
GLTpxkN7bRy5TKpu+x7EbZhGay/gs/M8aj22bctKLvzzA1y5C2xA1xUAjjccnJfgjTQGoc0rvTe2
nMlDAVkL7zOpHj/cBhYaZuzPu4UaetpSJjpjzgNs0Zdp/TFadioYI8qdW970M8et8BpHNUpvUemN
rBHekG6y7n7kZDZ6RmiK48iYF0yvKT0liV+0o8dKvdhqNrk7Qs3aHLZHoK8sOGJvAroyWfPe5kMP
EvTx0/6QvDJLv2sL7RNOZeBSOf7Whqfe080cqEoaMvzHIaYAlLuA/NNliCNvZe9icO+dj1Fltrjx
mBvUl6TXT3Je+E6pwXRvnXxYMeCpn7WHCpW6x7hcDueaJYIehVphXtsZiIdyr2i5Lbhiv0GUkKzj
uirXcXVgop8wfATbgnQbxXjWY8bxNS8i6jvY9aOFgmD4kguFSMvfSHNfXeuvp2iQlIeSAVOtYWvd
68+KSXJAPDU+DcDGzZp9aLujQ2CFVGncVJ1CKrw0otlI/lJkdbqNVTuTjJ6rv9OYgnG0Lp9/tJxB
0Sf+zE5sMQEKebcbjefi3F8Bul+pWcnGV22FekVIfJDrbKDt3sntzPHsz5ehpmBDreqYsUHqqiZ1
Fst38aiuYhreu89gQOrKVeFRPzG/xlwXEP0z6RGFnj/g3G8G+VIGgx06fl8ckcvesHd1FpneLzdB
/oqsPbdha3ntb0JVV0CVFnhwfk5xs3T3Q/AF9bWn1Kr8ZTy1TYZxtnDnzENuEG3SwLkAozS07rEs
08HueZn7ZS7GPKraA06txRvVdiHjdDVneRTvtHNF4QFu8oowq1zaeXo6MWnHV2szTeiAGOvGFQUG
myH6jUqdHL6a6FTYeEnyw/7b8+fInRE+NPHO65b0y7zdWsrsQ7MHEEANVeMLmuMzx2a6grmf5swE
uYfnql+c9L8xSfnBaOufx2m89JWiZo+ZSeE+43xLQHWV9Qjod3uCS7GyFd95Ddiav1yNogYrFVct
GPbCvZiT5t4zYJ+rSIZSM4sNKm1cjzJmJD0N1QZCttL2sd7YNQSowJ/ywTsjvzqMZyus8/tjkeTu
uHcKl4pg/pq3zJz/F3L1Jqiv3hd78wV+EoR+Rs9mYxEb9sn4/E3QTYp42yqsBkcU1M49aqQb0MNU
sh3wyGWpFE3I3+p8yZ90uUft7vZh08Hk06uQNGV5BfJtdB828t9I71G2hI4yEFfY5I2rOIF1recT
8KB3qMz8IdH7C/r7q7hxj3YQmtO/TZKHwSjBsj0Hpu41NOQl1jVnyU9lV64hqd/eHBxS5Hclm6L7
xhBbh5m4DtUCnhVwa96gcckOmkxyPOCQEJpD++4mzydXKnRaWhL1Lbc7jTQu5dUSTVgIkWJAq25r
e36rxfc49uKeYLrCxfZCe/P6t8nAuF8eUWfUdQ1si+0I5rWotIwFcw/Gx26baxnCd41yketVI0Jj
IlRxS4c7OodVfiXn4mHZ85+xIYUbMbNaexhkZ3RfQrRZ2BWWcb6GiuSyCfLT3EAq353zNgxQpFrf
DwmWK8P8qL3ll1g/tEHq31xkAo2uR/uv/8tIKEbIRacAhZuTwo9DCwrsCIvQ2WJ3uU4p3A+lI+rq
Xs1bsM3oMtxn5mVoiFOMmeOy19XQ8Ya8hyvDZFL9An8qzSE/cmlyWp7RyH8y4r30eJPeFBGNp4Rk
PgeeCok8kDBDgfG4t+sTxid3nUF9vhnJZ+YZf8R13S1h9cduLfln/IOXS2QJEAfnL8oWaxIVfUNQ
SBxY+lwahvr92pfoByA64ymztS3tYhC0fn4J7w9sPV9hWVa+kgbj7j4dVQwAqENEdukgMCwkoqz7
gUVF9j/csB1Y/+2S/OAcRVM6R9pcmRzqe3En6p5FoLxtd0TMIbCOQMuxa6n8OQHw4JPBTaSbsyN6
mG2tAz28BnQyzZ8zBKU2QqsNMG9Gxo2x8JXu6g9YaVJTvndktYXWfSv05a/ARd4wY2ETuJZbEwUE
PTnoGn3ZRq9lm+H0DM+meVKgR64h0ye/PiCa+9QTQ4Qk5kX2lCb1YjZemOw/BXKIEtqgq4X2109i
FXAYbec2H09eTN8gsNakPySmsiackLury9GpyjBi3KfhYZqpS3DA5y+ZACtW06rE1i7wHdf+qB0T
5z3QG78xOovDmkb6G/LPoHB4Hore9oeVFSg3SbJsML/kS/6Lqiy1vmCbhHpao7wznGcMs+cCy/ZR
S3MWOxSDjssotMKIV31IMZ7pLFUufsFLtC+b9Fq44Uxizp6+LYI2QruTGJb8dZtxE1dDCKzZE1Z0
8qPcCRcm5ZPvN5NB/n3J22NVivvRfju1ZEKiQHGgip8k7HC0e+BgtaFF5Yk7lfSr8jl0yxbds+4e
t3B0rPKPSu5WTKzFXl/LJ6cpJ1ePL0jc1pGC8Z4itcOwSl5QGM14dT5SMc5NP9Hwfl7gpbbZOjqV
uMqFHuI84BoY00Kj3w0YvC0gXvFEg5YMXWElVA3fBCbHC4u8Zsz+n+Va3X00CZY2go9R67YpYU2Y
2C/RCfSsjA5TNNboNnyWEPjb2eulKgHviGWlP5VxihLQWKSSy+g3utfJkUGzweMpDb9g2L1EDRvN
0xbSK0/sZenwAydfX2HDGRqaMjfafvm/vo5pfymDto3DHYFnRF/JaCDkzsjdmO7vsLaIfm+71rnF
9UnhRzyR+WyzH54xXrxUaNPodfkPO1WfyQCz+7GaniIRjGUBYexl5Iwp/sqbleR+dnadrg4k1uN8
IlLpwE5VGeNoznDWtNaBFjRwntSMPYoIOzWk5bj52SY7NlcN9/Ep7A22pwDSbEJunue0arPdDixj
5km52l628c8/8FzDrsvMN+fG1ZSYmnVNY8xGvOwjdPursf2uWjYz6/S2AmQI/a0RvRu45CilISUC
FKbDUdV9Z0y7CPh6SozGQGSgpMxaGGOHH3rZfNyIkrOu5fiTo9PiU+99nrdjb/vrPsRJzlSpmuga
C1iJyJDcOCyA8ZQqmkexMUHyYr9FxRzwVeI2OT6Hed9eZQFf6NLuR2XlgSkguc3FyziA6Cd+U4vH
M37yCuOUuAvvMpGLPoUH972d6iS6bZmvHgKuLFcaUaPaO0z7IGKiYqFHrq//f0+8Y02ujKwJ5ckn
C2/N39+JA7mz+dbCk9YDNLRo3kVYWy+Rnw6IDCGg0ryIw6uZxOjiNwRXIkWtUNcXsjmMfHO1Yuah
yK4hDzmLwb1cwzUq86kdvQ6G2AAkSFuCDTkxpZqnTgjabe388oALg09kW0GAYNRho1VomK2/cIMx
h6IqP1QFscDJbdBojd1YFveTa6iuSMnxRNFNJHnOx6QMznzJpxbfrgCTdeCWFIW+zIO/jxEauJAW
jpNZ0WmyWxihDPHNZm+GpBvpzjghB9iojSawQVeifaC239E8FKxLcQiQYXpMDrI9LrGlpq6cDlN8
CV3wHTbpDPBXM4+Ch+O/dOI0uLCofxA5BHbtFqbu6hX2UhAF8rBlyhpie9s2dI7U+4gkMqDu7fL2
k2FOgXGZVXoHeJ5PdWodkb2tDFpjpfGYaENP5BRS3IkNQnCclq/9Q5YF4JxKj1aMTqKO377KHd+f
tW796gDlFafZ0EgEh/QMVCw6I8ido78LpKUK+TYc2mzfeOPrLZzs/HU8i+qqcJ20ArT1wWIRKSva
dQuu+4fnaV7+OLl2fbwCkKM57ZZ9Vhlas3wjeocxg8C5Xmbyx+vNo9+d5eIjqDfmKeqPg0XvAb4H
GLlNauiMWklstash6pWF8gB+mwsJ9XkBoXy9rRSYz6DcC54H+TK//Mfj54fDDrkRr9khHZe/yCAa
Abu2yhKU2aeLoW5MTmM1JYd/M65Ig1nlFn9v8XreUntxMt2VT1OLFZpE0YR1dEiDO45ODoO5V1z+
DBZEx12u2jB31umQnnqJz9L365wN6yODBUvlN2+2VySGwzRu9ZgThnHHXQKNOBxs/wpyWXBE6EO4
nOiHpH1E6orwR47916Y8MViASGCg1flh4Idz6pg+JIT7FJYA6aBWNy430HfBGfAimW0pFKpfycVB
kbpv34wlXYs7IQf5DE6CqzxpoImmaFE2kiCdMGR8pNVOiqzEaKrdHGJBQqwsiVRCnHFZaILlDR8e
VP3x7L/QqMtRkVmX+K8+A9sqJBrhZb69arzjlPyHNzUsLbL4iZjsGV0DPzMLryE/RBqtzb50Y77J
yZnJXs+j846qdamEjNrXp1z4gnGiaKJJnBZPNZQTBBohYBEPaEfzTMQ6jVnTOn+8yZOIQtKoDEZ3
McLvC2uHx7aWkiNqo+ZMGp4mI54wK7NkcSo+y/hMGrLMgjiPTFHvIWZPJPmQ+feLNFbeeGC+ThC1
emXvU6A7SSUz1HiqHXRAHhVSLWLFvuZWUenNkmDMggKa1tn09hyfMyyLKAwLRq/kQPGZx7rCLY+C
EIjc91emI7YNnwLqnq0o6avazExWPF27NZPBqdTXlH32QlhQj/YDZZmohOURocIsfTZSxw9ctmBE
mlanY9EkFuhiX52mLf5ezlKOndw6IJkzTCsdOdzIgVqjjfGVCwP6gzKr3uJEnrcRCIzB72Za6KHn
5t0+bp/Crmd+/dlQ3K82un8IEsQdcdGY34jr3LWFt3l1DMPmg+nDgFJYEFA0KRMI3LRoNaq1FPmg
S3GOgiKvXcR3po8Wv92h1uSjrBZIddXEn2S2HGKF+VBS7GJ6ujRvulon9a3fkBjsTFi92Q8M7i/m
y1AoHHd/yw9mSpsz22g/Z5Kxxa0XHmLzXNlwfbd2Yk0hKKJgCuYQdebTO4NVTtgj3xpqHFHF8si8
QdJArhil5M/NlGZjJfkWN8eupvE0+dFY17o8ijYyZeXHLxk7izM6XEr27qnWNH2kzWyHt82yZn5B
phinJME6/UK6YIULPUoD72Uha7CDKtqaQ0CnidxF0D4g7tXKOC9z9oRJKCp5DREOh3a42I1FI5lJ
JiIuSxWEBoIDMLQ5wuF+2jk1nDHvlvqkpRgP7tJc/qlcponQ+XiGQlEV/+My5/eG20nr6GAPXAq6
gl28tZ9wTRaLhsqMU8blRnbIltl37y4xYHZR3xw5BlxsiU8XPcEfAyqFvaQzgCliG5ti3FHbMyoN
8nHCllS/Z/X0zSnVOK4MknReiPzj8SF74QvGOojuacNp1g6l53PMCBibDDQeSEYvuZdqlCB9U6HR
hs1vkXKqmGeWVwmi/kQly+kU3/5vA4/I78A3GIMoTC37U5HL4sAz7ZKmYkoFa8WidzDPtH/JGaYM
FvVWaIkdrKrYh8+q8wsyg72Jet7lXYcjPyPTIHe12GN1IY/Fw+uDKpp8bP+ciCgZJbm2b4hbvkv9
+YuPsyvU7AX97N7JGG864XzMOfIQudQsUIol45/8cEKubR+Yd5ysqPlXmZRH8EsQCTma7uQRSBf0
yAt5EZ5BKJXnZz0H179Q3bS5FG3onC6jmy//aBaIqU73m9xmgIxO+A/nXwUANQctuIwvHWyI0S1V
ucZHO0boSzzLtiDbDDYTxS4P2zpv3LV60+3bJe6SdEWkDQjKWT1ZZer+eZWNuHW4iWoBv6/rJ6v9
ov/mS1ZkK6z20c7K4azeUCtUzbVESGY41nbXU/f2poDfJjHX/Rj2/qIZtcL9GooVR9wNGlDBwrzN
8GC0Uk0aUHFnYq+540PvGlmHIitGDkWuNE7vac2xyg9P3R5lnc8MqXhKX1JnFaqvvRtdUCaPVc2D
9F11yr8n42uFoA1gHzoKzuhdJPI8XKqBd9BaYu0sxs5FQJpSU3QXufVPtVQkLAAVkoQ8Zqrw31qN
wyvVLGf2gqs5Blz1f3b4kSmewGF3MmCRMyUj4rtn5kfCpu4q6sJau6eI7YvSmJSsApZorYnaAVcf
f2R4nqhWZOaugZBmvgXQtuM5+fi/c7c0YdDMXnzfo8da6FZDkc0w+DLQu6NixMkAvGc3Vt/YP10a
2mYo6Z4O8EkHC9CRbWS3DG2/jkmyhfYp+QYHtDZ/Z6+93FvGJV81SWbdcvrb+8eNM5wlMiG9m8Er
85nvOkSmySdsuX1f8ikftkI0WLcRPM6wiifjouIKWoFC8G1o+eCe/+Rd/FArJJJKlQDubrXM262u
Hq/nDgjq4Mex6HYxwidF/ffCN8LaQBe52zIPsNQOtVb/OnDf9NEioNbHVVyzF0jYkJ39FZo1vT46
HKffZ3+sBus0As0Uwtt7/P6rdu1QIMExu0h68pfnShy+yE+lLLld490pLAWCduN2ReD9p0p9Ddx+
IP5WARhkJ+qXFmwkC3roMKwj4OYLtnCpnt4TSWdFQeNVlpowngq7XZNhHLg8JNVPYqGwkiYKFn9e
LZSG1o/5QJRIaGaYmPrtICK87yqccBLP6kkYTWYSp1nQG58Ac6A1YksIrFmNWmstQ5CWMXEH2AEE
YWA0qLAnBQp/iiIU/yhvUfXv/Vvl1EMCdowhzXOAUl2ifiwlujSURWsWWhvw4Y1dkUkPE1gHCPLH
znQ/h2z6jk2NrVReHfjc4PLH1WIO5uE8HdVpkRe2RYDlSL6CFl1hKVlaMW9LJU0gkUckKFc2B0Hf
I4exnzqDyoX7DvBSpC6aUJ6gmhYJ/oVPO7C8i+U5bOlg4eK4B3SyXK0seX029kpVJGd1JyJ34II5
4Y1Kq+yWR4w9A7qyYl106Yz6+HFfuNbuFUbT4K/j3yW4kEEYgVIoCjimmwr2hQ/+khz4M6qlpHys
JQ8iFcuV7pclla70fzTiakyh885G7UA10mp6W3Zw/xCJvEsNpNMAMRGElKWwsdoGhb4kWFOjNd1N
/ekQvhklxzfOsgEyjmH7GEXOeOmvcaU+a0zhOhl70nZeJO+cqWMXNyA17oaPIEvLRL5pRS00U3AP
0bNSdqGOaLkkQTvicEy+f5oIch/FFxA+NIammpVEM02J1DFhDXG/yCHe9OUXffi/cvwyYRm7ss7s
vYfFXOJzu4prtD9dlPp/fqkg/WQ9/FyLcDLOfX42szkFpM2Tft9GE0+1Y6hKr+PuVNMalcwpNPdn
sTeGjmXY63BJX5A/bF1GFKZo7dvKaszB75P4IelmohLirujueum/LONvPak061tgVe8TmGvIAU3Z
S+nf9v+RxrHgOdtg1LaMrmOxVMYK18QkNUaYVBXj5s8dtwyr1mu9LbLGA9yTqml7n2b07T6TBxJO
RzcKn4I79WPBXff+EHIiJFAS5Q9kToQR+nl2MlcSjIlyydGPfY5Uy9TrhvgPb8xN7pKIaHkgTry8
ZhmE5Qyjc+Da4nlIU01uFkAaEd2RdUxIT0LNcVS/hULeEcWgkognFodHWbSOF53G3UAC6MC22FKl
Y3wZKyitjOFArpIHDRFB2oAYeOTT41gN5P0KfKr2lsRC6lPFrclJKy6ShItgWZYFM86RcHB0agyx
sXiNQuCqq2jJ9OjcTotH/GaPmXlAx38y+yIpGRfSGqpGLgkB7BPbGAcc3Bx4yMg9WQNdxgBELlff
yrVfIBMiVwyMkH5dCBFqcfwLMMfJa2XE0Qk0nf8Y1r48umbk22GhTHUo09L/9GzVYZZE3rfLiFCy
a1UrEvqxQvE4e6M4vFCkjHPLBzn1JB5joio1ZaVZ5Xaa24aQG3Rf+HBzYQ2MtcbGc8vTBTLxTXA0
VgLSwHb7JpezI1Itaz7b7L5FitMs78rllDgHDhi7ZFrO5Vka66h5t/D3d70375OowNZZukN0/5c2
FmTk130md8gj3l31ernL8SdAiZQnCj6rshczKzscxietPau5s3g774DExu8i5D8b7SjfzxodsNgS
LFmIpfnJUBDNvUOK8TSw7lVlrwExQHblIDBC9S/V/8it23y23HdmFM71D15RmH17Q0NFczqkvwBZ
ywivC79kMdZUfzYBLt9ONCYOZA4Sk+whHoVHfFc32czxiK//vyNHFMX9kwwlAxVtw9RkL/phfryA
IdVgRFSWQN2NJKEDQ7cAWv36JVzeduG4BFuGZdA1dv02ZapL3GGvpzLbWGlyCh7v95bbpKQZnk8p
8Uq2aZH+xWfxU0Y1J5mAICdtfgh/PC8BoSjo+2WGdfbj3JWo9sjxcYb/Wp48N63gmrnyutNKGlKK
T8C9dGgw5U0aZKBsIqCj2FjOd1xWPVfUj+8Hj4WbkF/wtczz9ObZbn8zGUolvnr3/tegGiev6tbS
E+O9nDtOBz/QhnyIr5wGTOQozjtNZp6IIGOiDwcWCC3DurxMif54RMO2+ypubA5Wk1mTqOjnWFDQ
6BXbbL88v7+ZtXl3Ld2yIlxmHTU1pziy1IAr7U72bargMyfv4V4dmptM6fKpuvdVIm1oepcJtXaf
qt25nZq9ozz7CUQC+nXkgb7ZGkiqmGbTXL+EGWuM16MhT2TzeOewTpSw77X2k8JEi8SLAn/kuQl/
tU8qZE8Hbyy+Zwb4yQ55J+wRkOmEXSI/5ZYugPRDPPVSGgHM1S8QLjalBsBK7qgBMSrIpg+LSEcI
vqBeuKvEjsfk6oIDH6VvVuhw9ILvrTa222MIpenXtYOuyh2frpoWY+2+fglLryrItG6XiEVN8b/8
EWeMS2dmAYwp2SIWfGs6W/C7L3tZmB/jkSqYIwlCUP09k6Z3SSXUstWsMVrkQL/Qj/Ntsi91wNBx
RGCpluWlih9ifiCZ8IfNB0wLCaN0yaI9OQ11EEREwhcw8k08aPZbPiPwUaTk/j68xBUVdS9SYu+g
9Ywi+Ob5jaZVuj1l3Q+GWGMK3htDHfUN/0EzmTw7Lbk0eiOVAcKoPjpyf1i7pHMFwnN+x5rqcXoA
5xJQQJ4Rrv9JJmF2DGi5uBcwPS/s1UROwoK8Rkxv8aH+s2bBY7BFyjFqC/l0DocbDFcxm06dpekH
lOMRtzY6qsmm3djizR7xHPByelPHR4zMpxNMR/6GFyb4uYLXYnkaCTEuPAKHgL9cSWKWN5tQGWVB
BTYGXGU/ZNP0SG4SlkSnk84lrNziUlednSHaUQUShdV8hLlZoxR72eDPLHiuGMBGunE35b0S1NuL
W2X9wok1DqUIGNw38JK/TgytkU6+zaV80dbOcbvptPtz1670ngliQn4dgVLbx5cfFt2JPO5AWvFd
jOtMPSz9MqCSJEVzOs3HhvVRE2+6kKXrzKkI8QLs5agFKC6BQ5YJd1k0NjlddFCddcslk6Vvu1DR
YC2VTNYGhCNBrf3sUpD2nXNJlw6M+EJSXO4Ls8WxiTuEGXkMu0SltDgrcDvpF5Z7KjcITqeiWOp7
kPTtlnpIr4QxeuwJLKd7cwKJa6opg0J6scnot4i91ynwS1tbUB32hsq7gX6PhIDnYL069Ca1YidC
SQPfMQ7yINcjBSdMknSASDkjkPZysndG7tWA9xSh0Y6j8qjrfKtmCSgM5ql5uDtzJIj3VwD6YirG
JgYz9MUBEU94jEGvFvCSq35TBz43CncWepv5rFHWiOX/qZ0qZh8JU0nw1DTQJoBSakY+ZMYAsqTM
tiFT+Tr6R7lq2sqxqz8uKUIbnGOAEnA+fpCOF0IzERPXtYNJzCkB2tzuR02KUkotnhv0vupcjd4f
lmGuUD3xotjhyzQ0oLfaT8hjafm51gfIGgFlUw1jX4au/JXJ1NNtvarwJINYfgcjZ8g8QHn9Wg98
mK8egWgS7tM8kTCsZaaUecyX4dDISY2Z6sRETbqO8CVSiTTTrX3PLv4xySkAzwE7BJoMvGy63JKL
DpwqbfJU4WaG5zuFwIucRvFrhQbRdiml4E2upS6wljG55I4meWPh8iMWfIXkJ0HfOW+Y0fQFUBdW
a/KNOjUJfuvD4n+cJt76xrVCHKDje3YmwyHw5Qm/5qbnUiHw8GZ+pRj1ZWRxTKpR2IR2ObD1OhUp
G3x2eXJpROqSzGw2RkGuafhxf2mVJH9Pp9k7I9VpYZN4PwLRgDrnXuouPQfnQRanNFkYKbVeE4l7
RI0DvHGrvNByHcKoIm8ugiCnDY1TvV8D5aJoREjxzJPZ9VQTKxlggOKY8ou3HLWsEPunWoTuXh/O
k7uYh8JA76uk1PmQPoeOC1iVLUbaHiptBxADV8aQW4TfowFuOWvVoSisG9Brmba6144zQYcTk/hY
85H+dtpoe9OY681lJDmu+fP5oVl+K/2wbwQq7hzjY87TOtqVXDMq+uRlalks6cpmOirO+l/nQhYp
1KmIJVqRNlUOnPEDdS/qT+lZDvQwsrRgcHuGdzI5rSLAOqHqkYDQXMx3w/OMbS1g0dERHyMs9ECY
48KuXXPOeTroSDo2u7D3iS427YoK8oTeL7u+9j/4E1Gh7lo5JVlEGbcr+cJHDjcZ+3E114fMXcxr
8GBYwqnJ9Pmyq1IsJsRrWayV7o22pIvAYUIQyY21bVFpPlhbjRZAf/DwP+9AjqnIzEBW9a7scgY1
GgcOz+hZtmaJy4AbD1wJ0SEqOrlI83sVVY7Oqvhu9BAITkW9up8nguzST48OkwRyNvCO+/Mgtwsd
DjMcyvsu6sjgOg/fk5J+q0cGRZ/MHuWc+2XBrRW4Zzv4AnpB+PF3NlV4ROyDzovf5kHbOtWOcNbh
ME+tBTQtZQhxLW9MmXb7Z1eOIctd+SEL0uI4m4OHFtrKkmcKjlBuHm5PTdkJ9T3yfdJ9wzVnquw1
glifNP1LBFYGAb6lia320p5H2gEFCPeM1aHr/MCpy7LwmOs+fBagD8J3arCHpB3nksiwEdt3O2+b
+DDgedZbdYr2kfjnnQmdp0x9pEYMJ4pfxq2VwA15vcvUBYqgzATxAit/nVCtOWPaXpBj8QNf7fIU
c3oIgcD8vQBgJqi22jLMftt1QshuqdaMcGE7KZ0mICv5W5bBsK+gqLpZd5jZhbbC3AulbEqfGtsS
Wk7Drs1XiIyn0GAXBdEoCG1cDsz3PeLOzDJuGn5iQZgTjTdSPH3i5qSi3QZ/FcmuYWXvM8iLrwat
74n5BvBjWnulbYiYrwXbcYPslDDM7uLJFQg18hqyUwYDvt3jcY8AKI4ekK2DYpmmgP05OQbD3Lee
BGXbHcj039NEv442RzT7OY9M0U1kmnQDVi8uHwTEtk7eT1JJDf2U5n0KOx5pRU9iWYapE7Oy6ERQ
WpXS4e3bheciMXwd2HAdqbdtckSLWHJlmaBMbL1JG0iT0c/iPVxfhftas8/2vQtKUFYusih8HI/J
yzLdKcdr4ri3BdMQt8j7lailG/gOF3/2tmD6LUvK6jPlvGZA4ZF+RXxnb/o3i8urFbLmpgKXzNbk
TQXa8469uN1RQRYgDU5IiZQCKegXqTnJChWnBPh98HJ6LiiGCpP1Eh8TbVZwy6ngiuSc7hmgVouf
DaIH8IP6Rtviynvb2BjEiLe2qlJTHjW8UuLDI9oJ9OVoKRABie8TyI/AkxICNWq0KBvnz4YujOwz
p7ZcUQYNiM2cJf1zE3Xu4k1SVRjBBpruLgbS+45wecyyVF7JJGPKoZktayvcYEeBAEgFUkoDASrq
u4rxzCKZ1212UcKhNosjhPly9SiLCnSE/g/nEWPFfrNW5iI+U+uWr708P0o+md8p5ltWBoy4PkpD
imAlyZ/+fwFoZunwtZyvXI47uBJeAZSYHElsnBAChn6y5bOS7scVygreOdcFJ92+Yr/L87Uy/Cw9
/CwJF5/qmSxC7DxP+bGzjuWoIzem+giOiWuogwFdsMSFzKd+Vnm8BGM/jngfMwEGvUM0LS4Lj0+T
5B0u6fVMp0i39NemLmk0juRODGYVDZ5qU3oQXxw+lN6pnXnhOTM2evb1t7+B9L0e/1O+2lDrtUrs
3cjG7hqADwcrUn6n11PFgxThAJET6TYTh4oodMdqWHueSegBNqaju97ITmDR1W0xDX6iP7E3lMwZ
Sz+FC4CBelbomKGonZHe0/7xuC9dCJHx67gOB0UhRv2X+0Oego9r3TDDen8JjgTeVhOQvrLSZTh4
oJnAJSnODjgZzAZkrPayrxOJti0VBqVsZ//Txb3Ce4YxfLBUNZqWTsZjDBeInhRO0J7ULTFFrAG8
k8ZSyQ/sgWUNvzXtLA/UqkBXC1Z2crK7/hDDd5s6sLvHy5zA8PI2iW0L8W3Z6JYYYEVzSMNMkryi
Yy83iLptszBmBGmCxt5c5r0FhcWDQDKFtlytHFiL1VHp1uTvGMA/ql+Ih7r+fPA4Wbuuupjxh1kE
s5NcIDd1pnIyZenugF/I81tUQwtKqfm9UKEf7XjaSFZ/2/xYFou5+mZ9kWt6FVh7q6QHgKx1pbvS
8hAMj+G3K5lsHmiLJLbDWLuJTrmwUJQpBmn1TtX6odoYJ1UyS4GwQttOOSScSItcYmb81t0MZpKc
rWInMZMWsAfMbiI0BImcmxcCqVzElrsW6vTFFwNNJGWTwvoekCRAgAycsKQAUbWwTHPMQq7NNruD
IjNSOIGDwu8NU6gxW5xc9+J/lXvEuLsg9MaIoW8VeZdiIbPxP25vVXynGjSCej64Zp2qWRi8qsG1
DrAXvVNF4JuOTS43j36c+SMiBRKP6arh17tjTJ2c8V6SlN0q/sqZqTv0cfo8t/MsS+8za8fXL//4
2VWoPAu1gUaj/5s7Z4pgPaPwqQPR5vVN92VKbSiLQwUUAHO4Xo6uiIXBqP2NkJ9uN5UlseiGIL0A
jtnxrVPb98zIBEwus+2CtnmaATXQVAvKYbQCwwxl8cWNhyaJ7MN1C3gLGZyQ30HrHyYMyuFFUwhW
QJbxl0DdqmhGfjn5erGP1UAB9duzTiExUhQ+BJvvhPIFnN+5h9r4tsh6S0jEZ9bhxSlBKtEMmYP0
T7zpWW/NHObPT9ZUsqFgqT8KdCyeO4p5qXETc5DXtnAfd7M5kp5rFgeFtOkTu/a5QvUdK8Xlg1BE
QVAd6GHe1FZGS3LAm9JmeWd50XEbOSgj7si9swZiq1J52KwCNoaCdguEa/R0ZXV5MOSrGDmcJQsz
1E1z6CSswBaosoxRIik8LModvWkOwqAlJh9/y6x1hkrx4IgtlVnLAxV9tjkdasMIULmi8DdoFhyl
nsQ8EyB4LTF9dGVeB4d7Lx90yN+SwCEReXBZGhyFGqN3thN74Ka/l8IhZ/qclvpIY1wHwvo8Gd1n
I6PLiennmhl6gFuFGID1vjUfay/m9DI6Tk8Iwe/Ver5fqW17Rseeo0KI1TjyAkuGEeCUu78pbLoR
+DenKKp5rllb9KooFafV3QAVCee1ZWWucGVKFiLm+JtSMyIIkdTu59cNOAUWkKwJd340bbnzdMeI
LYYTyeR1G4FRL2MiKQXiy11c7yO94fkgyq6KRUgcC0aoh8xDzw0oTingkWTxMHnYckjN8En7t3B0
l1aq/TPvOCpfnYaRDAQo3x+O8v2bxjDD8Nv03R0/slSWCPuB4D3ZppdICcHH6Kvm3t0VAG1+GIHA
XI8wYwADM0Fh0mf419S12eRxxQ5MOIsCDYGVwYm7iUBTEVzhkGO7bTovYXWjl4XQCV4BobkFzfbA
NoZ/4OjuTW6sAPG0Ix2T6rstDWfwi1JFrhqS8pVN03wFenLRNyAJLwXLFBWco/fhknRzE/uFqDFn
r02E6SWoadqFk4A65xDMjkwgpsMl4O0ye3awkUVhU8h/j8ZWmHKdbMEiGeMOadxvDgIKU1ToyTPj
uvD5wTSyMcGav1NtfrFqNf+f1RcQyPrdZgT/WJiCA1f7AZq0JwZxmBY4EPxKqbjFfmzIIHZYzOY4
ZcTfcP6XuzR3suz3u7xrO9NK7AOF4qEde0bv6ulTH3K1MFUSddUCEoEKEBgKyfVfF4f/8+3s1xgn
DYYN2ScnsmZ0NpOU67wZDo17LXMlZesKkAky4MnxUqtg92rTfG4NP7pBh5ItgDn8BdKtIchmHQE/
GggDeJC2XzZpirSgn3pas7XmfpD3wNA9IvvG+CHXXgYbD5BrWiHO5VvQkhdAeqRGXEN83Gvr6TuR
H5yRgbx0zEQwP3DuYHM4cAuvwim/C2CW78WUzcHYtOyAvDx33XpHMKPaQ3Fcuxa8yZ2K1JJ7pPMO
XhFuJ+gUOqcJgNmNtajvI7ME5tmeCUuCUR3HctjDcV2yGYJ/FZkHl28Dag7EFG6qsZUYqNan7pw/
X6RAcWI/vvALwJsQgDltOFGDva1Sut91IbVu2yE1/GhL/u4KPP36rst64bm1iOhnSJ2TMQKfio7l
8A5XtBCVkTC+mfQ9+h9rUlf6RM8CryD75IhaVt61AdrAP/MUTZLPv2VamuhptQ99m41wrnWvrIrX
/YHkL+mfC3v7wIcUkEkrO0BFDubn930RrIL+dpf39zPNP0RhpfZbVPZ7/nyqmP4WDhlkHZbpOITf
fl3BORtOlDlAEu8QVI6HymdQviOJgsECn6KS8LGTs7FOorUJtL1mcEAdwpNCHHBbxWPdMutELfBn
LhTGeX7ORTXuaX2qcsD8SNf1GK8kvI8gI6z2jUevgyJIrEHmdiyfQJ2eYBS7THphFs8gh1v2Cuqv
Ow5hIR1Rprwf9/KwPOpxtTEnaLUJHHbWtFf7kEWhgq3SbESLcgempACZWNkgip6MlwQ1jryPT5kG
VkKA75N3dv/y+cITcT/ew60k9Xbnwz1pVt7/KLTiCnCOGcycT2V6D4Z9e2k2IWtFhd9B+oERIpl7
ax+4j7fqgVYdUYsX3ut1JsvWLKOHngU7ydH8uLiShOFQBNNdRCZ3QlBBYLMGjn3Z5fXHn0RXUa1e
ailOA7xzA3pyw7kChLOq+v6GRRbW25h8SleXTjY6chZPAF1vvyPZHfhwspGfBVnNc7yBHNY43ucC
1vWXkqFAMGN2MG/yMboKrNoxLMVH3mp65aDyq4YyT2C1c7LL8fd6jJPT6+bvhV3iRJY73qSn2XTe
THdltBsbTaZoDOYlOOxvjuLal6EZj6xHh7iebwMqDKnrqGdLdcGhIPErM4Q4dHCB2u/tfu26fxEr
PCebuqyRa78aZmx/Iikp8INfDuPdTgNfXLsoCbZsz0okxKJNEHnJP8tFEEcoYWcMYFFoFjAmFzUt
WfJ1vDUXnyPkdvq3s7BjiXcsvoVEseEqXQ7sKTmvieBb5qyBaESk1taizunA6SL4XZm9wA1dDCTo
r0acAwp4plJLvL09fQdrsuJsXgoyFciVJclQ6vJE20uR2flPwH6RmMXJBpjmWO2nNhMBI6sVbHqI
Co6PqacH9cLOm0bkpVHf6Ws2+QOUQ+gFi2azk8v9bZRGJpwirz5PUhadn9VXNENLuC2OH1DPQ0+P
R3Wb9GkNH7V6Mw91KT7f3ME2pP4iJZCBTQYjlBbvoWaWLAX2ov1u85OPsHn3iz99DK/s1R/K7/aW
ApBlKBx9PBLnjdxyYg1JokXu+x+LknkSov/D7cXQ/DtSC/BtQvm+nLDi8j3IcDknRscMx7uKtIjW
rBYfghXg5/ylW5ypRx7g9vOWVgB2SH7z4j077wYEx0DEpr/ibZ0/28MfNy4wn4eWMToCsR2PfiyG
P895pUBZmXOWWfyrp9ksqjobJaulEJOAjfhTiUmgpw02CmuvicmFcpvLgOM+K3ZpQOHF/f6ObMPw
v3jhUgZjysDdtGIeYutu/RnBA01/B9RmBcqg8+7C/evk70D8FTncuR/1jwvis1z4udH3B7VL9dJ1
PLEN04DXhnKN5T990JfzF8SCiWrxY8/yAbm+0KP3LZajJ/4a1ohdQJbWI3n1vsaGkVMwvTWvvDzM
oIK6P045hkcRCFjrJgwG13ZDW6TSqnOdc1NJBOOexTR6M0Abdb5DsWIJlG8yfD6ibOFF9/g/hIkA
MmO74S4OufqD2sfmX9MExSArTJ3Ebpj6kXSsPgJdkul2+0dMuemat5qLRAF5EsMnxnHAlaO/rBgs
KEk0KMZeYiOm8wat12TN5sQ3H+tf6T8snTPIUpVLE0MVXoJ3DKK4GFGZRiNKSBabN7fPhNcZokYC
DeEVzQ1+gwbaqBnrxfQj/pkPBeJx98/a9sOm3d2VzYYMTNItJTwR/h6XXVOS/YJ+FKQFVM5ksfTS
IPjQFqQb+VLbSeOvP8URaAIm25yxdecsUOi9beDkG2IA2OVGCzP8NKPxiMAi1x9K4Q62JNUYWnDg
I9e7dfSWMLA95ywPv8ARS3CA7YQ4ESXSp3iytQdBj6e5GsGG+pfYMvqKwX1OQO09Fm5ItQAvsZ/x
jYKhHbD0dhMHAzNV6a6EQ8YC4QxEPIDApYBWMe9k51JtXbIQH6ZDiESvnFrqpO2eZRD/PfzUP6bG
e/H5snXX9i6DrsT9/STzQ+jb+dghAVViZOLv9k75fVKseIm//rMgVMovlp5EkdKtmIsyzdWVLT2i
rhew7y2k/SqsvyIB01xMZVknUF3DrAxEFlvwakFYQasCzJST2NFkOs/WiC/zDzTsOgWEew1eWNb8
Q8//PbCzXhXWmqqc5kPMKJwhG3RVoPHjFFClaxzgoJ+pAnPPsLX1dDvi/l1WChgzfQKSCgggZ/J4
nmfKzgrd/Recbnw/ltYCv9ZQaK99hNy4BktHVrsL1gtEg5z+jF1MMLAQDAI18EtPdYAlNEklvHV1
ZKaCN2qK9bVwpia4/2Mc0F6cQA/IY4nYGp/6qETtE/lo7z5GYJEfFhrWj6m8JyCuKreo5Um/QbpL
DkJCV+KHK4hISyOt1WNf2Yb8bHY8gy6wfpXgSWym0nrgGFgE6Ol+ImDQ0nHAjjKf5UIdjlEpSAoQ
wzz+2XGizaS5GXlKYwMF7hgFU3RAbr/m05J8WkhGNXJ5G8VFk+/JdHZtSjkB+djhZ0TRpiOZ9gwp
DUGlYZbR+PH2SkFAIznTOLCOE8N0ClgXJPmTC0Aqp+/V6vPMobfqAh84PJLcgygrtx/t+zZuuLGO
t4kQBfwDHQ5iie+bFAK6jbsPBNjBRN3e8LxshPS5WLlEsICvSQWfYzhqCXCFQ+n6Ym7xCyKF00Bq
LCBIDHdQTvlBQJoJ7sCY7DAAOn7vwc6/ck3YIrREjVKVTInLXchQUhDvj7QUCt+yZdU1O+QyC/lg
0LQ46CQNtFDcWUzyOJlyGK6HjR0EoCOVC9wTxLQxUOu8WbedkRx09h8byVFazlsMRzCZmUTNVnZf
M4rdybmLrLqbWQBOHFUITXGfs67wS0hgjesH897QjNr0fT6CccTJM1/OzlhV4c5sJn64mPoso9So
eBh+Ff1IK4DeoX2CSqWE6KC8UXZlXJU40Zw94uMnL28EEfxDchHFXxNd999zy3xhr/9txuOqrIOV
UlewJTv5cNbC8wgKkwQPidcCMYw9a+1/MqW5poSDg3UnIEmFFj5wGX10viUM7ysNeSsKa1uag4S9
+/ZXddl1YFmTY6uJIJGwUQ8gdTSkU3rllA84cchAzkZkUiOl9rFpkR1JDZyvbBsHQEBo0jJ644Q7
QDTBYp7APAACL+K4mT9beROw9YsEdVYsOOgE3OqOQvTLhZcNpMmhGdDPGGwBz6KtxyCTgEmAGPoh
PWKeMOUaZfkWhacN+8c33WY4wxtW8D8UMOohM95fu6jVdHWokyjdwqaxZDzn/wg9XECWWNC7kb6u
kVGgtfUyQGfIlkkS6LPN7fCU9jZbtqLie73dku5LTWWHAs/HftWU0UP0V+VsWKXNThoIAyI05D7i
4tjCtoCixdd+Likb/rox14S9PYeq2U9tgjwa7LM4JKBdDJzCMPLHFw2r5iTLDxR13ML1VLtgYIV3
9mOVTa7J2wDH2rQzwP2OptaYy6eEFVnc80x8UPZZ3sUBdTezmWhDZ1V9qx3/EZNohaJmzs+qim6p
pq7pBtJRnuNy6TbY2eP3oykbXnBtpWptwGP/Et04Y6EfGhC6LpKzzoE81pmtq2e6r/DrnnX4TcdP
pYYluz80wlP2FNUUPXskX2P02tJbqcsSTm5V9EUR4qerQ3m4GRRLwA6WWxCvadZVXtDHiVpfDFY7
krAcXolqWK4YnutrcFS3UCzUl4sQINehE6DtBeauZIFbvbDlHJhqhR+Vlkd0zzKq5kmh9QI6s0Cx
9rGM6VXjyaLc+B65MU/3u9HDmGX8ffg75tPMyBCE/7bah8KoiSbvTMcV3TmjHiqa1NQgj4Basv0M
kw7/5t/FeYGg4hf8CwjtmnecbXNrDhgCsRwCXlU+Y/QkkNOnIm81qDAZdnS8tI7RqV0wS0bZna5o
J/3svxISmJZoJfl3kruRsBug2AqmLLVYyuZIYHlwjtNxqM6eEZY5j5t3VyJfIvqdCDo7Y1yYoi9S
WE6K+E5cQ3PofApfuJ60VLkO2Cc3TlAm2/OtkL8Pg7M9pvVrARRKX3ct3TObyM2iYrE24+4s57X4
OKSbWGIK4RgLm7kq/yyoJ0qYTylABAIikz0iXmkqJrTSNFWj5qmcr6IzQDdTpEX1VP313Ip/hUHP
U0fe/YGtxn5X8dEyvCnfhs2jWUJfcJQ8tHIeAwnVjvMiQkjoOasm80awlEN+LSYLJ10GB5AUI/ng
yudRXGXZaBdWFg4N32NOJd1hRuZVyk1HKxnvNCbZXTfUqm7517hkcEbcZxeEKDcjmApAAKrWCC5C
qSKDpCOcJU9R8XarH43wVW87ypdqvYwWmBRrW9ISiz9hKyXx8c54S1cql435omjJSzY6o5kp5fcS
tmJq6QA7/aozjQNNYt0yDCKO9Eu5xMrELMYR5Gk/Bjp49XOV9STZ9BZms8mWomGU5wSpoJ9emu9W
b1Lr+QGeO9JoLeH0bw1zIP2YMrHvmwiAILs3q8EU9p5K75CdzqBipLWQ67K0UpyAOGTU9/tbcNl8
kQxcDRHn/TFRbin0iEL4ZkhrPG1ekHHINtP8LBRPxyPBwxCPS3uo460TM2Y3oC5RoHpSpCFnCcyF
h6N3EAGKGyl0Dimbo47bCux/elIiiIsf+YAePXB2CSjJst1JagoYk0T/GUFivbEMeQXoc4YdeUwB
WO5PRvenyGT6fFJrZlsIusl98B7iotodlAXy1LnS78l+lTHb0U6Y/4baXsoLGtZBN17dBLr7iTOs
n8xmlOPmwEEHKHblOopt7rGobXAxIqFZvmTFTxIgAQYTIsF8y3Y4NpYVtQOWCc93y7RKkYfgT8Go
voAjevUWWrRn1EAAD0VA7caVwVygAcgro09rghah3xT1TfPMREk3ZhmW9AWr59Ci8FILo/DGo6O2
PhLrcjh7xQKK/0ltCoWSCNiG5QHSmoYFM/Gvyu23vd/JjqErrEOgQNj+VLxR5pxjt7jB7+1caQMT
9RwyaHkQfHGHp61MsnLKIq2zZw3SCXHMcwbjoHidKiJ+6PZHUc2iQc7M0EK9Ul0Z/NMVS0jBoxAp
Gt9gfYIl67c61i2tjv1DFd2yIju7U5nr8O86tkU8n1aEyUg5K+Ykrnxls6nCdrSDezY7uy9iNYB9
pHn4nS8B0jNIVpk39aNco9HAsHiBSVIIIX8HkVpOVwzgUSRa8VUboHTQ/MPPF1CLtnBvTFHv8nCA
qLD8c1EHIPpkWhRW9bluWsEj7zLck2zhuzOan1lR7EtPxa5X8ImsF7g624qJd+MO3kNQhcXxLDwC
e1Z9X6tjzNozKm/BshNAQd8hF8B73otWSQtZM0vHowXrBUXQltLmNOdqWEG1/tpY13leIwH+Zd7K
NWRJoMdJX/P/Z5VF6sDjwXJ4uIyp09ksxqRmmSMd06QFK7RlJflKk4X7PRMf6N5/3kNaiIWCRp85
BpHPcpn744Jc7zNR41NK9+fkLRSkXYq5r/DIdi1URrCfuQ5hehGJ0uO1eWMb3GKyWWqtlWG2GwaF
J3BuQSDpvJTrtb26dcC6NqyrYn6O/aQAOcJaB/VfnSynrPea3yG5XFGmktGhSnhTXgr4+yjvmrc2
UJ+g+Moh38kUxHoIC9bSWkaLiN+sr89HfeGlTTaUHCcH/oxXmnmX5q4rlK4UZbdCuOO4tntX6wBo
3tPx5SRt7A6n0jsOzQu7FAnigSjO1cdY3u0ZecBZPHun5jDJ0E0NlMlHPVNyo4AN4n4NoSrlSsTj
jIsiyEJXZbwDdVoPp/Tq9rbYYDsQsYGzlVrQrh48hb6kQrku6sGdGLQrM4U9qry30j+vBFGlTT1B
7JquZS5tdP3Y9lpl5EmukQxJ8hmK2noZKtn41JMBwnf0xmJwPq7bwrO4N69fTTs4hNAfp5zTK776
7GQk/N7YLEwXQQ3NaNec6f+q7PXgZSq8tz1JrbAZqbNHvNQ1Wow6e2B73itPhLjNrEaKq38kHlfi
5dqa+6iT20i8i7CR7YiP6q3CctglXW7Pz5cm4AUfwMXVjQBkZK0VfzxpY381kmBnPysGKUzUIpzu
phXJJQzmsvlSV7VpKZBBoNT1S60JR2eJMLmcuvyIVCRga1cXRkLVwyw+KsYYsG7Gfqo/XEmN4HA7
LJJ/191DoUI7KyvZHJd16mjxS+ZeAJlwMmCsEOmvuqPzdbCmYN0GgdbciKtxgc3JTdUlam6ygG2x
xtOKl+QG/lN5Qij3mAd9mUs6W4KA4xCs1OXI4UIOSMtBdOgQ5Pkgtc0xCF0SuGZoP6jmF2fqWNi/
/vkPj7not3dP08/bNJzog2noPzDisn6v6Jq+k8yctNttG8JUypwl4V69uDpE+UnFyXuN8l8tlJqC
AFLI0bSoA5A4A6K4yHYVkaZ/JcXOIQSJvpCzNY+QRvv0IXQdNtqCObkUr1ZSZN9E1v368HMfewpT
PWfftf89EyBeNn0OF8BEzd5HZ/FBV91E6mjt4sMDGw5zqXyV0Ntpuq1XX/O0V3LIKWdPwxIZWQg4
wScLYWLol4E3FFXJOzZcOdgWU/sMnYZpTWZgjoUqTVsMOf/Tif8OT0teQ7e0JH+g498ZGtn6YqIS
VRFnXx66U/0S5Ted9aasWerT0yDEpoCVfJb5e8bpfvGcHpCH34EV+DW8oWAsfEjCHbr1BAGlFpP3
ufVhmgYJzXe99pPC9cqnOm7AGzw+WeNTgJTke7DQjqCUApLI8wzuZEgh6lBTTV1ntlZMZ+Hag51d
NTjkZ4bQoCHurQYRFnQ9rUGPvgofNVAJ1INqygvEeXqiqNGEGQQ7NL3ShXPBpb0tjH10ZnQibf5D
fErZ4sav6VVkKAJEFhCbm/6Alo04wC6dzXHtEwNF91r+XUC9lL9Ff/68jBzjRU/6+nDB1/pAwJAR
mSy+9QH3CNRpNHWny8aCYepJMQQsdxgB6CLxTZV6N9jRU+EaYJRltoHfDsBJnmZCr/w1gqcnrIiN
Kay7f9o++6sJVnpg8q1tki/pF8LUHOtBQKt7A/Jzf7lJCqBKoP0hR9i8C8+KD7WdkAlqmwn/s5YB
jsjYFyKFJe6kDbWHcBK1VjVnbtsCiW8FWOPM746abSJeeHc7i/spO4tyFsC3qcnp0oBDp92xkFwN
So1Rbth9vThk7BTIe4Eb2jL4yLuneIuSYZ8jmdglIVzPEQF/ydo39KNBUZTgnwG+ubbE/+VlzZ93
XdHOAWzNK3qgguhClmUhHKzlBAGvBSrRJAfgxfSHUw5rfBjC+sSLTUWWI6VEad/aWI6lfR1OeoOg
+j0b8FMqpfbdsYxlAHDnwPORHE3w92JZoD4sanZlLc0nWm9cL4rtADjOZrLkSCRCDz72JOdOBO0G
AD20TYzv+qMObJsJiuh51/VwsLu9FPugwzOIqForzWJOf/ze2MMYqk/74kTArOIXLr0iKHLcqyjA
qbK8Ekd5f/nL75Xq5Rs+PnF061OPrBct0ZJwKZLdcG+s8U+8TPijc6nMf3EdzcQJ7Oee9btJWgOy
5x47GNkZdWhXAS4C+G6iJ74aJIs/VYCLhdDtiw6vbBlfYlQPaFWlwBb2GnEYrGIj6XBUx9OYaFWw
Chuar3v1MOAyBvII/vBVzzKHX56z5ZyY7B99y/E9jknCaeAN0YEDNh/CpGCxlA3VrtuS8QHosI8g
2H9rc9y9DObs0cYLvJbjc9ocJ4OvXHHXIbpYWyvjHoTVq4AENxFv5XHQPhNV//tHPfRoihspbyyw
IWGzSLyk7cHV9LCTG3Iy5UDRNf2KbpKsByhocik5TZsElvcQvhWQ3zmYI31jttCUjQvv0LUmWEPb
boT5HMAzQClwQMkc3WcPDlH4q/27xUzpZf1aFIvvXLmC4iYAEdlYMgX2LSZskgK2WD4VYADw174y
swavj/LXz5GVFhfqAqZSZS22LuadwIjkcUWCsPb2f9iI4F8M18Gv9itlEI6gaTyGGLaFNXPm+fTv
mbPMqSEGMwbLFq1OSOlXoWw//ZOztIWIId6D6mcjacHTzCWLXUAnqsnLHPkOnZQ9qaYS0hCs69w0
Mp/Sga5SF8NP9j8I9QTOTS0iPPQPMT50AgA7unTxV8tqcreNh8daIlVHnFCwTFuI39+9503vtYF3
m32Eu+V1vFB+vnxJe5A3HKUBtMEQzW8wbXHGGOds/rA4btK6u2MDrto5Wu1id9QYXFo97UJBReA/
yBOrfJFvZHyfuh58xOcenmgONmy3b2YuLt7vxV9GdN1GzFsOEsycPuzyRHApj3HqiLuHVth/t97g
Uijehgf7NEK//s4GsmjCiTrgBuX77izpAGrlZXD5rKKw1jTXc6hNohILBGenFC1H9TVs9mnyS6Ck
33UDDDpfzuQSBN6jYsRP1wCkyUJwh8NTMF39hHgKTefB4WWoZRpLkhlxHv2V2HOeJLJhUDtrCRG7
FxpIgHjrjLNticWSvTrs0tD+kj/advpb+tkwCAYcy10m3PR+D9pJUAUqSwWMfl9qv6H1f6F+m3ki
NU6Ytc9DwjpkFHtKwzkOLhMriVeCW6+DFWitq5eRCwF86DmQ4ZiRYmlxhxTCMJnMzIXcIiHnVVTb
AOGD7Q9lldpGkOu8wxk8oLnIk31VrmC6ipuH02xIK6yio4E/TW4Skb1Rzm5Aobun5Mc/JnT28kVl
a3wVTm2fQxX46XRvaBEa6Z4eJguDVNU1hdSTG5FBzcFWTxnowAgIJG1q5NgZUzKrbKgybz3n2918
XO6+SiLIcaTYQS4T/nmOaG2oTvwGRPyg11aRBiTvivbrsGAkUkkH/z4tlSNB+mfeMG3xVDfCm6VB
ACDaCcsVS3+xROfVVZoGmYt9gJBhjkZxhMHMo9qI/fNgi0qYrFCTeSLOw0sNe9Oxl2Ge/t49VKhZ
Pfat2JjrTzU6Ub6z7zsXUqv6fVI0rt+KH8/LpoqsYBU4GZErG3eD/Iugi3VHiUhVDV4fziA38hBV
6x8/p2Onm4sRJ6O8x9BGYYNM3YLIQFML+ytBVegevoEGX9aZz0xD+XO1HCqWLSlVGlbk0hC404r+
m/m0Y8cRJgEyj6m664sm0ht/BfU3qeJRzIK8Aokxzmb3y/esVf4ls6mMfbwuaEqEg1Gzp6jEzuU1
fBFIgq2KxWZEZUI0qyo9Ui/76GSmqKgiUiCYADpyDTmRpDRahDD/cLcFBlbS4JIAhfxNlDM7bvw+
ZIK1wGETRlgaTU3yoemElROKwBtI1ngMMK/jgCTI5m0kPkxAMaKRD1kz7zUhEHC3dCMseuIISgRZ
6/+vpgEciTAWsYLh5zFqcz3Brl2VQCz6lUMRj4jwmEW2fDzrTeRyPyRwWYEWjeW7vkQ/wuuqLwJt
exk+vkj7h0xeO9H1dJdRHeyxWe1YPaBoN1c25pnkW9q6GwI+CyLdSNEC6xp42BrF5sGxuME0caP7
CEvYDdKYRUvy6pWAIC4goUrInK+DV8LfqxQET4a7+/Til6LsJs/rsBAo1P4FChtyGo5FQk4cV+a6
bGVTAKo3BLEw2U77qcntsvhNnEDLlrujycSLHKWW0N8syF49ZoF79ECF7J6NQFgKU3gJ4dxw20uO
m87sadqpxFiKax73G4kRNWtdJMbOH1LmpvTfkidOvbu/81mW1uVDnNAggLXkw1P8jChMCWEOnKSi
h44YjWvAvwilXA2QRg+k5SAR8i9dtgeqXJM+LOSjFotCRI3MMib+lBE/boCjBP5P7boQvi+65/WW
EsAnbPGwkdHMYLqyAhzGbvGz+4ubSH+MSXQAW9wAIoPsFrpRf3iJNnbAYeeCFOaNNXN3ZvvetbFI
N5RNJI/4+LHJg9sDtcsx4Mqa84xW6HYm3nCHOLxvjXk++g+ZTX8lmnh1L6w14kv8vVgX0Hp2TG21
qU/M7g06Da0Fbk29Jg27LE82YAPKJ/ZjsjM5P9IYkUL5tm9iPaxUTu+ct49U9AbxfQKj5H323EIp
PmN8gCSty3sRDg2gnZM1E9obhvmVO9605i9qO3gx3yx49oMQX6oXjGUX8atKRFfHbyhvPM+k4Q5y
9TTLuhs9tuCHc5+ZdtrbtjqNkiqQkhsR1BFh0McNqWvtup98GwlA79CQSZ9BMAcT2IUjxcuQ93eL
I5WCs//lP255BWlqUU/+AxmhrKfLsMGKIIGjJxs+nCZQcqys997127VEi/zhe9I7IhjzLW7RIFmH
ktoB7X43hlm/eWeZx/7s7jxAsfrZwtNtnUQVGSFEZ5F81RJ4inZEdhLi+trBekJ2EP11Dv/eijQZ
rN2rBh91Sy2SEAI3lfeCXvAOGRWHSN7F5l98+veKBwaFj3rM1F1jgNvATesguXmlBQqnQB/bx99M
EHiFNCDagsJQidWsNiJdjIjtYRsfFv3r1kHfuGd7UP/cVU71ZlWj/KqbsYk6PK69k9fAu5Cb8HCc
NH8icjIp9GUwrulbKCjIg8KKzHb0rC3XOxaJdLljW7zvhXVjYc9Xif4uR/Vz0iqBvLY0qlxPtmJE
kQ405KMrwdaDqmt3z9Boh8v/B6npc/zvVLpEvlcK0n9N2e1qhqFVaOcvkvlL4ken+bG7sGJ17M0F
c9BF6QHQFez0W8Kf5HfKbQvxui9cblwulfHBe91SAGmL/pHq7XnLVELEgEs9QLNPeh3MGkloC3Tx
We7tncc3icEVikZqj0P3BesrJ4ShcQhneK/Bqgk41Q9IJT0hEH7oSLZwpqljrmDEsL/dfNnijAUl
tioXH9PcKn2CU61gmckXCSY1CiyoD9jW/wyU0QreCUSciaShe5313h0etEwug9B13F0mDnfMY6hS
v1G0ywT6LkHitgPfZkclFqAEj1xfxgiUmokgoFKljXsoDyov9IFm+yYm6bCtPGaCh73RaHmqNICi
uxtcmmdjKzRXpzGbL/gya30N4yip48X1cw6X4ueuV6bZLGUYD1Xw52YErAydlXVEn8u/5hgJ73Dx
26wYjtTIiRhbYvyfpAtvava5x/j54+mPCWxDTzmURY83cdR3dWjT2S/0REMxfQJ51tZvTDxF+JRu
dpBBQrBV4Ts84a+bz22olOyQMLUnhufOYb8qRrXx0hXCDLJTgmTSOnqaJI+JRyoUxXttKeWU9lzi
afS5pVXE+tEVuBx/5rttkIY6RLh+C6iXmfziCrwrIAP+zJ1PUaXJu2Fe6Hy/LthO0y94Cy/rAzcl
jIrOpL3GWssMhQW7B+BUINhOFJlzqwSY8e9kYdUx4h84iHIpLHSFtdKvgDlKkOGPfXwoZC6m+jwN
kbPgI0uu3LsqfDNuUlQPl/27tTlW5kMJDCA/fHRZQDF25TXBkqxQyqkZPvWW7zIGjFdQI5gcP2v3
ZjxMGHAhOgy07HDdRNkI1dM9SE8zbK5PV7rC9s5lof7Z8e/fBKZODaOxcUYI3E1DOBjaJtEmQMFL
WtTpXMKeciPotElEW5O57epLXPh+qj8b8HWKdfOmpeWyPtjWwjRFWzwdfPqgz+I85VcF59s6jZv2
ZuiHhljuj2/uet58qjzDyn4RvfRDO8bad1/63smgPquhFzAaaJV7yN6zeZsKQ7wFk7o8DJSirAMn
insoMfaRQz1FLk5N8pC+32+T4lL60LPL4lAk5V3A1C5RRcWH6KCNo1WN7u3F7UxMQrJdhAR/USwr
EAMHmRWSK0NMz4fZbkYq7C+5G9nIPqpGMvDDqLS948QNQuMSNRI2s6Cr+TQFtl5ARLoncNUjFvky
8acwy5DOU772U3aMqXeLgDBx5SrZ//56AzXtFsrSuVzaJJtJEvCQ8TZD+pCEAwTsWqfdM7YMf3ZI
jpA9xHHs6/m3VmltloIT7Rs9baJOsRSu6YxugJwa0Ipx0Z7muZiLvHc/P83k71RLmlkrX8b6+RUa
FvrrRu3lt1NuC8+ixRcHpf5cJBR5ZB6izcvwl9nE/z90ADXJz0DQ6IzRg8x+QcwcHDwDCkE8nfSx
OYYnCukAE+yDnBhHYotL6s91zMexm/qPtvMmTB4soEoHExRHxE1ztqciT5YSJxc6PniutY3EjMly
9bnkJbM5OiFOGECqzF5Oopq6wr1c9lFfhoAJS/80Ypm+JDZkcRsNXiDwfl81eNxuJ/vtyDq5HlAL
Yt20BNRvcNCJwB3pdZlVxcQoR++eAzGI1ECaMO2b4imCjCvees8qfSsyNDgxfqhZyluVWq5T+bXu
smScjw9Btxne1KgeGt//ywJir0sy+6ZOqVe/mK9mTQzer1LxXTPlpi7ZePRlKCvAeoPn90Rb+lPR
LFGMLYpxL150BNVEbSzGh1xq9uoYTRsaX42LP43/w2d2UNNcqY4RcE2NTZcNa5UfsZN9m/xUqIhk
FjshNXArkf2MbtAaaOYKWbU6W9o2r5AOB03mI2ER2hkomv6WZ46YOxTUDylk1Iyov3JegR2w0D2Z
ZyekMpwwF5SeKjY1FSeABrMCmXvc4V07t0ef/2tKtO12+46BZ5eK9u43DMwtpq/+oXlHoRLwbBfu
hNgnfd4UWKt29+9/jTuIs6x9Z+WozwjpZQwoE+XON3p9u603UfBPjoBEO9tvSMhnxfkUlKuZh00d
YLdmf/XWjUISiKOlmiJ3NuvHG23uUkrtr9t0tjUF+QwKPsT4PDhFG5w04/RmYb3q7htzIhApbCkM
5dCfYjPXoXXblJr2pdQ0+NXmePE3BWhcaP+fW0+5UL9RhRpG1mkExeAL3VJTlg6m71Bx5XM302C9
6+WKPY5G4ww86Bvvrgn2c2K9xGdDxCDBq2POy3KwbQhm2RDuCqEP+nUwUZ3f/DZZTjTCs41q4fZO
r4CwgpsTdIfL5v1td2ZrgQ8BKMqLs4/8D35kd10jwO3uyrxNLy14yTbXVbSIsbIa5BjoFawEXwml
1hUN+HnJlfhwj8xOAyG/q8YUAqN9y2XFnGsu2+nI/h773i499LyOdLPw5k/O0brr3cQ9vjerxoeV
m2e1GIfVubh3vuiGkJu398dHe1wXRxkAek36yfo9lEMo4k6GVKIBt7YYDT474FdHjG+5OBSvNlst
4ciUzD2XojDQNlBEAAiGBPkLYPj4MAMudRygrLvigc2I/DpBlomUVZfxL38+qq9yy7E+lopK2FSx
JEwIi8Wo8jYHEinrhHrmqBP8riO/0itPSKlElNBa8pHoo0uHhMidfbyTS65r83CkFMm0oBHWod/x
XxP46nJSQuOB6CR5cwxU3E2Nkt1BGO78yuOFpQp/etDdvH0K2eYnvQ8+4l3ondlsJZoU3MpUXOZ+
ULetBkbzcAt11IQp/Qh5aUUeyzL6ojX9lsRTQS3Cxo9B4TEyrFZ97/XOkQWweKTpB9UjU3VVhQUj
2s3TCAEyb06m4BH7CnlmEym8hJOWeiwCjPIwxPJWRjMLiMb/UMhVGrwhfoW5nqa6cKzWuHzJfKsH
DJbsni0YtHOg0OR/cd9b/lzzfWidriMJ3o9DjD3pFWJvIKPzDG5tKXPeis58TzMRDbcKBYZzqzrX
hRHaGDk47zQLfQTqdcr5SRkpGXCX8Jy33LuTZEpmIr489Nrh7XoG3/U+rhpW2+dnQuiNyuyS/5kn
MGD27VZj4Ohc3t4/v3rUN3hxpRQG5lx1IluZLsc+LG1i8ug1EYQE3wUno8Ydy1LvYtZkLpkL4qxw
8A9JZeXv4uG9E4Qd5VR+218qI1JqjOLnD6YAC8k61M3xps59FEKwr7dRIHKB4Rt6SHi/snSeborF
S4zZ/Ljf/Fpx/BfYbtYs5aNUxzcQReIOjVhXJfaq+lfnlYQNyVIsTXr+Rx0gljsqp48naLt9eKpF
rzhI2P1lOOEwMjzYvhdp+o+MSQVP5y/O/dxa0ivpdQT6aUUk/TUQyBPLEjhncJV/S97y6xwvmknG
NE5NtviUf070GXzGLkEsy9Y41f4LriXX6xSaknrzUiemrz3NVB5B3+ssziuGt6KDTNxCBp3TL/td
tOsFocy64ihs2iEGuBLUPu8xu6u7h32Ols24FVL4SHd8g84fqhH3bQ+YA4m9X8JnV3Wmjh0qOYgn
8hBdI8UcXwLPWXAM0XfUQUBsD6pIxhVl8qbBU+lahncYJ3pXQnFuz0ydymjXEdJjkxz1GdysRO6m
SsxaiIpNXGSF5EiOY+8u3zc//7d2AwZzsWSc6RJly5xRWEP+C7fS4stMQuVsKwOQQ1Xc9+92yBTb
OH8sVsC01bykxq+QSt4m2lG9vz9UiyLCHG3WTFNdbXpfN9KHq3bDtUyQNJjBL5QK9Ug0C84uMAlH
lD56zMpI22dLemdHZaHAVZmn2j6Ss8PZJU2a4UMiRWPbzfnkQPcbNE1qNTBfQle3ifbuzBzqKRLa
VDjswQkVV+LSILrmze1aWjC4RE9pW3fmyxTDp3WENQt3Qc67Iwrkhm8YuwTQmZ/B0uBX6NCcA+AA
z9HUdQQgHNJMhT+wKw6tPDP5KNfuMysf58QY1BN8qGZJvEp63MxFA6dj9rCxYJWyQZ+LjZa9UyNA
b47u8fEozILqll5sV+1t4mwtNquQvL330JkLF5yhDJvilavZQi0oJ9DWjs8NwZ40lZNx0p0MJesi
wvoraLcBo7QgjxljN0utsOH5ZGmT/VpPOXj9ROq+cGHGJHgIGuxRe20Y70IKPuQlV7+Aj75O8Y3J
UZtrX8m6Ug34WKHgQURH+oZWbx0R7yAJvwh48DikcaBJaTD+o7zW6bNQVKeZKA7hDnRVEyYQIQd4
Swfkiz2jNAVmcl9oe/qqdOEkXQL48rW4Iyy0uhdXdaBdWtYA9+DIOdo1qV7m1ct9OhJ6YIyVult+
ohSpKsD8BpXo2O0YUGe9HQqNydZVfelqsfyrVZ/M5WfwnA0qyGlaYFs3gmPtzn1S3HzPVB+ZwJQh
aqHCWtdWaY9omNAA6BrpVoXfBkzjEouv3rYblQzs2cNHceUJSiwQpKk6TuqXGsJ8XdpuhyTMXCPA
ORV3h1ZjhqMkGEpYv/F9kCk68acPDWADwBcKz26mAIvNJLI/J8sVLW4SuSM7rKO5/Jv/rEQiGN+O
ZnGSMfeD1bDbqAHb0AQh7JlEkv6YWsWS1SuQiSXzdO4IbqmMWD8bmPGBBMkVeuPvAqQ4M2mk+3Qa
WtCWfe1Tx6ZHE3T500Zo5me8XlioZ0O/ro1YYX6m1ZqUgg2XqAjy/FLpcC4oZauw2rub9CgAhRNt
LtmZvsoUko2l8E/FHhWWSDcoKfFlloKtHrv2sNQJxU589bJa4FVSOH5AXMcbOB7MjqDPVFhuU5Nl
GVHyH6q51KhHeJWlUse6KsWYE1GtHbK7Xz73O1QnKKV4YTKxT4auexC56W0pBD1j5ovj1BlkkY4q
tiySqei47zubZ2LrOC+5sTZo/WYffRbii3ich9LfI3JNiPDvquHG25P28Av894de4OJ5hib6B9sh
xyba0pJEJ3Kt2q6qT0wTS6pgBHE1AmfjZs8vTdhWLQv3GhtnY2q7sIC4QUi7IJrUQkDsyq5/c5KS
SzQxzfAldpsOYxUU+mPaW1zWMfSTGPS40OB3GUyPMPrF9GPSxLHCP/36+JA78HJQplBKrJ/jrlNO
rEJaawQ8PXpntLWUEFxKyljWeJFLy8O1coJcDF14SUWDtUfLhsHR2yWnoXY9f96MYhA8BlABCvAH
SrEFGtCQpg+nAtdnNhIL0n+RuyoNDgZZJcEmlw7/42IhsMXABwYqV2qrEQIwOXEDMFuKdmRFsuVp
B5vkhGcfKXfzYzUDk55JxyqHOM83mF2kyCe7eB/w+TnhiPInZWapxnoCV5Alos56UTiFG0WQ0r5f
TaOd9zFQSRjrZ0Wr3fJlK+GjHLxClqko6njPlQVX1OSu2W+nmkB1RZ59BmPFb9hbQf5GxbbnJ6lg
w+IiP9Zu6tzKCXKdT7Bf0HaXsBm04Dlx0zVh4PMCSA/ooQ5k/MXJloGKJPWaUt1xRctvsYMEhaz/
HERsLqljOkQ578OgrfXjJbZ2NSMXuY8+UQjMKaQUP5JDAO9VCgrrv85X2bRe5J2Vba7DzRtTrdHa
PsGHsJz0xTthx7wLNwUKW2KPow7wl5LSAcQnB6m6JP+k5hKTefgmZex/feH9oBNHELHgCM965eD4
k0LUeBJKTAuppM7CfUU1KkVMYCVBg3+gd9RoZeiA3pDLE0sK6zfMnXFBg7cDSYZt7uECKdoNiJ4N
OgSjKkm8cjg9QhZdfzof0eBc0iHBzx7v/paeBYiHjM0yxVQY0S0jWgohxtihtSzJ5l265RqCVQui
0XuDOuzSBYxIwY6MYfxrytBEXMxAbNdc2f8nBdoCSr215jRsn1BonWyXZPnIg9Btd3PLLuCo5yD5
jVc8Pc9AZZdW4YSW3/45gb9p8eOGP/ShVYDtx/ozFxqc0BIKNs07+fHHlKNm3HoVv+i7TT0Wvvo5
+0vd9LaZoiyDYFdZrBd4xJ87x0bnGD6HKaGVY4hiFOimJlsFTt6UUJcIK7KR15+Omi1SZ9bA1U6o
PsOxCJxbx6yfvfFfo85r/dFvpOfo4LNIRUoPCFrRp3y8MWJbHC7UI9u0KOP55ydIKgez8xeIwVLJ
Tu/f9fjSiDiK/ZrZly6pTviu8R2HHWVINQN8yELy0plbI1WOGLXkzqEzX8+g/xuEi0M2lxs/Afjk
qZYu4cDycIWEwOrEYp9OjpmX8Y1knuFh75ZYyXF6+nGD9ocu2kSiNGrH4vftJV+DwbI3fEUE7hcl
+9XJiCgvMIh5mfZ3DtIFpfdBu93rS126fBNl23/ibpW4AjQuWrVmWdSkD/AH1uFGo49KF/TNpFVI
//QA/lb0luuP9IzQMgbhVRbcok8sD2playiDgIX50lkVdtbruIhTvHG7HjHjQIECrI55FeTe5S7/
bSbuKoQdQYkODt2s+XrvRO6a4z6kpwbKopI8GQ179uDQP5B75lq0fNdWFeHXMqf/rWTgckTFFyvs
2XfcPFhT2FoXtdaNKxzdoIOD0Ml1/8MY8PwSR6+dqvsfAUvbd4mdYcl49RfwZdCQVh0W1/SDjsbe
74U0JMKCAuX0b1U46TergxPSbJ/pvmTJE6wVr6PI4mPfn3xHqSzcoFBboNpQltecn/RJ14ijmKEz
YT9d8IS36KtuK7bXDfxB+MWDM7gxEjxnv0UNGuVjjgrujZKPrH1jpvb+8HtvOqncx7C5W/pBztun
2BUXa5fQDKWYEquAm5OQJA3xx41NHR3m3dwguL8/MoDRFRYZb6gVWxD5WdkXnla+BwZ6febLCg4G
NsoPxSVzzIuagAvOx9pozXBVgtm2sNugiw/jagidHZDBa4jAAKjZ/Ggy4FEFhiG8zG5sU1rXhbGf
DT3RM3JNY3UUqug+lY1W38WjuxGzHbIl7zvI98hNQTHB2+VWTMBJkAmSfFg9SBl0p+/s8dmN9UBH
ya5251c22LPfnQFs86fa08FJYLuQz+SF6gmsxQnYd69MuyPuwhog4G12Y6yROTZC/B9+/02NxZsu
LK+7E7/03XJKwEQWu/Lu9uOsWGO4d0cgtmPWcqNYF/BnaMfJL+9S6ToTRqFKarM7EluoT9Plo2pz
oNA60i3/jyPN4hx2kq2hVUNxmV1SmCtOtTCiW8UB4rt01MV2f+q35JHJ5Ta7MOn/kxwLSXQdT6GR
siDy6hNrYQXJBhZWtFtkvIZ8VyI7ObNHa7M9pPQXYq8K+3bpNpox9EXxib4yxBZbUpY9f1b6eN0d
rAbhaZvvVZY06cUm25TjeufXzY1Qctc1nTA6+HyNL3NC76872Je8VQAljDNUQ5QbOiGyPYSDrEAu
tZtQw9nFSYUhLs1bDu0nLv9lFrWhS9ngnvzgK72KyOIl8qAG5Q8QK6oCLxUaS7A4eYzdZA6LT+NH
xqtKwjBnK1AeMswcWslBTB8YBZ+pkcq+4lha+aCPa3JA3nmfvgnbweEfaE/zX1PpkO6ovgOfUCa/
aPPgNTEht/4bXkodOX/Gm+vB5FafOq4PGMyLAbbuwsJD9dXSohVBiuToFJw7I9VUoWR6Nk+rEbxv
2YrvrJaWJFSIpeaZ3+v/PLYl2KIn7oalnUlunko5cJ7gHo5ZJR78YIUX0wdHAqXd3hYhOOkOxB46
u0iKqaVFr9JFLJsb9KgTleaSvMo4Vti71aiZkKwZrc955IQcFyayyV1KKGgF5uxq3H5OtNN1SGhU
GkQArn24MkC9nhmLHpv/VSP9PQe8HL5FEWM1aIRAQ6s8bsbW3ovybWf3trxBRZYxs125Fo+Jjp+a
RZqanMgXXJovG4U36jy0SUK9AF68+J1QV/dKpeCbQYS6DD1sOrKh6AjARy9VgkOdaYPUfsaEda/z
sIqda3q2SHum9mqrrAlHG+pakvgxQ1VG9iJadOvA95Hn/BFXg7dPmvy89geapegFCtbDyIA16cD4
rOvdLBqIRWihgn3gFZhg2mrwuflawf8lvFv1JL6Vpwo9viCmYZVB8dRdp6uqbbiQMqwZtV+c5+5i
JW4WIKtuYRoseeKNAh8ey+6IgV+2jQq/GUhRFonJXD8UmAp3QoXJu+FIzulqp7G2NZ2AjyRdMb9s
hDN6Z/u/fIE2lYb8IbqCAn20rRzr4lL8VrcpVGRISTvEqJ0w6E9s1urv5/pTGvynTluG18wEJqro
8CmcjUU8fyYu7lfhJVm62vX1EaBVMmmyyd5foiRDOxscv/Nl7w8J2S5QNLjYy9AhGRUevCvM4q3B
8ah/URqdQkUZ3G2u1t01R9QgmkiFInq782zxFO7DC30WUw+JavwCdTq0SuEhCDBOzMSjo9Db0zUO
aB+kTwRlPDWHEMkQkAwSg8UFUBnP3dmmz36tyhNMc/yy91cyBWhXX4XUVtRBKyqHhBCVTy7UufoQ
bV7KAQe2Wx7xhrTmTmh1CasTfu+OOk3O2Gz5lSmLKLev0FV4BaWwgr7BNtSdVKd+mNTsb3jAug7n
eJhNjSNhw+1g9Kf6mC+xQh+EoxZ+UGbHU4ly1p4yx7erX2VQmPnU0bN71DKLljyHcf5buq4/HZI/
/oWnb5SDTjD51JO3TFhBB9fkq2pbGLZnHPVyMsFLx5ei88KuNeA/ASKMlsc9Gw8SEH5RVChGg2H0
S1otI98v5wqjHlTDTgVY4xZ2FCnbwZlKeUvm+8ZfvAg/5Z+I4UZzsUP/IlVGyy4HGIwok04uFuPH
4ejva8Pf+PCtCIdV9WmOkr2F3IMhQCqFxB+ewh6/VnHBWIDu0mYxPJk+RaYZyuN6m985iDUHreI3
246MKaoNXNvqYQYgeR1XEWk8KgpExgLY5S4w3kK8NJHEeQl7RfhONLDauZ83WB/jhapTWsb4IeAU
P5lyKhutZNwWqYrSEC+D0YTRiKAssmdHo2E01bvSXR9ASMoyDUwuT/9kBxSNbdftDNADChhmJ0Qc
rb/Td5zMfbWLzVC/7KtLo039NcOjf7uy5P0GTgcCbgDmy2ADln/Yy0s+VL7dcy1Tae9QsH+Idgs7
nSfEo3M5t1Jop7cyW+3maTyINsAJ7aYDyBjqXiyriyZ7PAwCkqnn6EJvrKL5eKv6Wc7IqUfnpmOx
YBTI4SRxHsfRqi/SzLx5gvK4u2rQUTwKteTgC/XsELSJ2nNAnNVRMZ7zzYzgDthytQM9KvVmqmP3
Q+new+L9gMi4OdzvRWqE2XnF+3RtiLr8eThL49oDsje40jpoM9AFM/YBalKr3/tRno9lIh8ILc1q
FGkDzhO4ILmg6TUYDcavxGlA0r5akj4kec3OC2MXYYGu+MMvAxwRLzzOTSMOkbtg/4TNa5SCIX/r
wl3pye2FdgJW4f99CkkSn9Qeo9prnxROs0UjFjx5Fox5icesVnQVQUL56VEXqVh8OFJkjwYcUCn5
xK0CB7WL5wsTXLS9B2HBNfcrYAUROZLFtBqsl1DPvnoxebVd15lK1NuvVv8BaGWabK/N7LPC/nxy
FfoG73m4Ctzt97j5c+zV95lwhFZnjh3M6upFVj47m3WvxiKbuGJYC7Ia62syXomN9paJhNUgUyLk
9T9K07+nuVL41JHfbqbJXGSrJs7xG5n25pAID7Zjz9I7YBpmvPqsDSdPM2PR78n1UdZDz8fduO3e
6NwgTPQpB2aQPMNeFdZY4lIZexiOV61ct5PbPihbwCPrtiL610S5TFW/Gl0jLsoX8NMkiZifatCG
UUjes7bGrHV3MFkXzD6jYA1sCaciCeZ2wuUc6GKfz+OVlngr6cT4e8Od9vb09E/+8wyAAlR9ZsHJ
laLjPTR4xhBL8OEJbxh89/sIe0fgZdyQJjcvztAZ38SbqM+mfsBXaFmpXXl4aKPDW5pd6iC0K8we
J3F4uMlDRQVLsjQlP/RcXcdgQtjvSFVE5LaNtq+8L62EHNwvaQBVLyoFd2+HCa46Vg/lYgzhnGw+
R1FlQY43f4qVcZtQJcbZ1d7bWI2JZkKh/9AQuJmMplvRdik6zHR488aazkpeuc3jx45ORVHI2kin
h3OiVUzixgZsDkW9QVPvHD7GfZ06VfSFlupByIt/OkH3ZulNblUHu7vv3XeYjZY9nO4CFT27VHwe
razAeukmI4/SW5pQqoe3xQwdlq0gcZdw8y3i4ds2ueQ+BuvaEiZRfGfn9NKdApjlY1y96uTK4ONS
CwXPcG6Zjm51cIOU7DsC+F2GD6uZ12IWFW+o5vUt4dbyFia1lWs+qmlbjJjlxpEepFeZT/DmkFnv
ksCmQ95WdYFjRo25DdD1/u7gdCaVE/j/38pfsonSs9pRjt1t6OZ8wtM48Y4WjOzbWS+MdeYbQbZ+
tSeU5afVqwZacpALA0E1m0zIsOb2BJJzA3XM39NfYo7VaXH9HIfFvOFGXVdf/LBtWNEiqbKHv8/u
r/OcjHrH1gwRLgAjNXfoWNu/xxSy/NEVQ+93US9qOo6WbZjs0Aps0gnBxcdg8PbqItNT2nBBScZS
EBXinxoQ7O6gbgjwM1L8x87A+WlnEhw7h1xy66VtVwDpwz3qeKW5kDZueZg5esYUh6Bn0HMBg2/i
1stG2CQ80g4ygLj8GLeRwqwr9O0zCfcfApCoKna6hxiDtsdJl8Bm1vTYQCL4/muMNhKbMNkGap0P
BfuWiRI4g3wGdzBLPn/Ea3TyaTPLwLRo/u3eJ1DA8eYXFkeTuV+IIB/KTShlHIWXdr0WCqfzg/Dj
ZJECExQHIvXqITdMsUjCb8Y/SajHAzHnu2Slux0LlusgPgGSswjO0GberAEbEb5LIGpMRR+UY+A6
SP0pedrCoZnc7Lh3Uw0aDscXQwephyouswxl/Z9jUKkDaQ8MDLAO8yUwkoMEf3fl+7wzWT9QFPig
O4VLGhbuQOb1erFlTkC/sdBvTIiZ4tBQ6p4r8guEsuuKYw7TF/PpExF/SCFbh32RZyxHIMIbt0kC
C3zlpTFYaYN6qfQav4sThx1tJCmPw/HkJR2Lnl/An9/sY99vU9ZWkdYf94BxEr9ShSvvYtDnVUaR
0WxYbcI21ZKZO6UNcNDANQNpplPTVQZBDLVyqHvawmLZ38cNa5C7rjb4vdVu3jY95gr6JrQYZoDA
WaYur7k+V+NvD7EGrkknc6drs3cpBrOMe+Mx/DeoN1y4g6Wmnc3kIyyAt9NrxQw3wOURAcqdPQWO
vFOAXkyYxNBfA821dTjLw9fywkE5x7LB2yvK95wIYGpkswzRKD4XUVNEU6M8nOPUYmmcSPlDEXxT
LxQF81Y4dq03u1H24ppNMDqK7dN8j/BBaXz4dvUqPMN3lWRY9jdiCgfp6VYno2D9TJ5AsAl/30Lu
ZoA7n6GoehbbbLoQQMaDdynGPNsEMoR6UgQpfXiHj8/d4hshc9ispPcpKZUX2puTHJH5gUTsYEc8
pMxVUcVPK+gJqbBnRC7hZrxvylLnlSwFp8lxW/JBb3hRWAo03FrbBqS1V0/GttKpsUX87HM++8e3
vVV/f0CZj1iEV2dC5gw5C0RziKqv/PR8DBw/++Sd2KCC1FP4PKK4m2j0dPMLOEKxUeFacIa4WgHe
8PW7uTydU7GR4KAxbqoFvVxjkOmhRGJHlujzNlClHAxZNZlUHouBuVi8vy+7HmsLqjZeK1T5IjDN
PF5cUvbSnNLp2HbRs66cFExhZezcKAUWCedJ7oSI7hn9DfIKuyv/NQXVh8uvgOxYH+zBoXUo6scJ
LfcEo/2cIhB7MXOIHefjL7e0gU9xk13GeLIB9XfjRrEkGUkYflQdOvn6eWZSMQhSSJUYdbpJOYsw
dKvl2fYA3kRT8pcp42EZ4P8lL9L2uxp5gBxz/WuLSw9vyxn63GAlNhg4Z8DirNOPATeBhjONrbQA
TWxZFHtDIAONWQKCFqodJq7HEbuTW9IB9YqoYVmEp6NQswW/xXGq8VK0s5xow8t/IwzuNe6SV7Of
34ULo9SjMwr17hlkK+TeLmC0icCpvuGTwDtj8884rEvQfXXvnnpM+62gdvJal9fpv8UhfBxrHhMO
6ecaUHU0mIglWGQbkcWKjkscQz1nqzhX7UdwJ/NO0QhD+u11NSp8skSSYIjyFuhoN+RBeIw5Akag
AaZXBG2CCoKhmBl1Qv7VZ8i4v3xiSh6CADAYislyuxjYejdBR5PlOiW8MKs6iGxr5JSNDIN4VZEg
h0hVMMoyOv7U2X+o/gj8VZZYWs/3k1LmicOIFG8Zmhb7Hh4cfUQ1Wv5nO8F4jEeCB1UqAVlo3qS7
lsbCF+VlgU19AMrx3gyxedv5Ljw+Gl2KxEylZl44FMQQVnNFo8ia9DcnPiD+d7e7jY7J4SXHHCy5
HUm4C0varjxkGC+AXBalSnQ9eme9mztSzkEQCKFP9XAO+9dhrRIddhIw10yKJIizOaaaSe6QZ81f
wzXfopTJGZk4sftictGav7ZTpQzDeYCuUO6A/IJmJeA/yHun+cQDmhduuHZVpNRC/FrCbZ6Li/fY
3HsPpRFE3PW2tQIjRrMvAtnbJ1M3+neMWe9N501XjkNG42UouGgMFYXNSyzo6+T6qKd6dYaHImrh
N85zC8ZWGCEg2QSC7WuTgiebgerYx/P37yKi71/GPLjxmvHetrBGRczLhF2R+ARTmE0opDAfZb9h
fqfN3lrhkH06FweMAHyDZ3Wz4eOTZNnPW811Baqzfn/Ld46X42vPmAFX1PCXHN3zv4L4Eh7Tj8mA
407TEX2Kq2znpwsCkTP2JZTwzzas1058rkIMCqAajgeA805qNGUQAYterYn8eMqJzYc7csfORFB0
sBWcgo/8OYVHFMtjY3ipIc2UtMZETgOvFTTu5NMA6tkuSsmIVa+B3Ns9hrU9aM7LIpCYORpKmkOP
FGuayaaPCPvTM2nuQNoNsT2/p7zCqPj0K894wknBU18caz3ZamjpsMqUGPNYZsLP4LMyx3fqH3aT
MeCEmITNWZVSvD3dDCrWd3ELHHjyrij5g4ALvHA2YrDXbNsXuUgFvncyQchjYyzJXMqnAzR++fYD
UR5fX0IlBavybi++IhdiiCrPAppbkRw7cZHRAhQZumN2r6g2FnZnMbfcK50CUgpUkkFpUj3CtQw2
0EQ/B3zFQ+N6Vb74WwVsh2fm5f/qUjudzODZQBOikpIekmOjx8Rtl7efeSTxiY6mM6xtFFrNvWMI
mI691HL4R1teL99h+mHvOJD3r2vOOmCt1Kp1iGqjj1qNRKgqVFtjiqDpay7tXNk4K/GTiYB0Gspq
iuGIOgIpYsHgm6mMf/6fbY7Xc1wmFZLZcTgSUwWSpkHCUB1hjIQ4lU54mpCavu4DoX4THLXsdzDV
Nlf/6ohW5RIheX4HOWKhyKZmOfmLxZcUtF5QSzce3lA34yVLle3CWOuXXslAnIOtDXOlVMWuC+av
6iJLWJ9zxI3+jDrLqqeSMA+1FLSMKd5Kycm0/utRL3u4rmD3aj0e9GAWoQhSBtEqCA9XDP1NE2n2
2JWPp/a6QNvAk3Gi9IdNAzI7jxblJAbjVuTQh1G8lfh1P+E5GwuxW1FCFlV7V96SRQHqHqlhVmlb
sBOVKfcl6sqs5mex0AA3qbd6yoHIiIic015PfrrlZPf/hjEEFaUrRziy5pwOeTCL8Mz8SaAkOHQJ
FyMoOQL6cKjmI6ke4Q0NQEgvFawX1ZkfEPjRsZBbnqdXoyn1y/tVUxz8cQwTYHwPyXwzNmF3F+/z
Gd6RRmYd6XPUwcpFUSFrLO+Xq8Y30eVAVsNGHGDq+bKr9INrtv6eYS6kQRQ73NMuFiEgjDLCdWM7
oLOKJt8bQr3zLwwmQ25/AiiUmM0z5/PksOif5vXakdV0sgywn/JpPUBVhRtRSgQbMvcHb+ygZWEV
13ZXJFNh747SNk4iQvWIng0psg1UuvhZlJ+GVqpI+FoLEJAPbmxxxQ4y7CKQdEv98qw98HOc69jp
jqQmL2XpY/YwaGVVpkaoEds4JzzyfVs/l+wh1pUnaFuC8nMH3jYKhLOhGfJq3FBkx7v+6mLsGqqB
ewBKTRdO/lADbH2/NVb438WPVC8W8ZG+7NFbvto1vvfmR/aq/c6UW2UY8r1MRXqK7VdaQLoSjSB6
r1bRKFZFLL7Bq9wbVC8Puk4kyiiEKSGX+1XKldHwYH6ryNV95vUDVP/rXczSfmo12dR6jNeHfXR2
LuexTsysl3+CmGBXGJwj7QZFQJr0RrR8l9vr2/IveoZxx+8AuE8P/7bz/85yyR4T+3gKdq1pUSXY
9K7SwmSxbzO4c8Mx1aKpple/OmCXJU/CK4fhR4mtuTsez98A8/2GM0xBGHmvCZU8qh+8f5Uj5glt
VIQn0hetsmAo3yEDc5152mLJdzoQdrNTQTtbP9BlQexQn1X5MmGpaONPD7QSI/N8mgfHpZRXbN24
uyTYA2YfRgdm7PcKHplKO/Cctj/mFUdVdpHDer/+72fmMx+WbEg07JgyiYwyToOTB0V8fOp/YAWy
k9aPH8WCxz45oMcmahoT32JgUShjc0cWQPExIlwRB9VihuUzh8V2LtM+ogxDr8GpY17B11kT/UMy
XADXXPNvAXxhGQpovmBCtsMxlIBeqTKy3WAVCjdqQP5e/zlvfJZRmoqbXuTtpLBJGRDc/PnUiZBV
0keHCvvFR4jsL2G15uUcMPyVs1Od1rhuMKXNseHTc0y0juq/b/xGHbS4Eewth3GhTcJKh+x1C4C6
DYhC4gbLkyQb0oqHVrWO6rxLLpof0HX0kLdegH+fKscCsEIqRJ10Dlm/Y9uwwZBUdVQdLbooMzhr
FKhFoR8eTqcXUKR3HsaC+RKJP8DDTTPPQx6R0dMifN31S+OgpCjINg1xgulJFEB38XeNBqOoZjBj
WtwmGcSfmOg98tb7jqMtzCOhU/mtvGlAkDOfP3UKizJPBwfjWi7VRGCPLalIhKM/DolIcJNPAEYY
WBxGpOhJ2pqnP0i5s5w9HEuMMWoypWFywE75+JusXX+l9+C3tTQo9XRI55c4QsUTCbxnObej/bB6
PSbrm6NZwDZlC6nXE9Wdd58nuOvVzYzFHOQqah9PGIo3dUkF5TlrPV8J5NsxV2C8U3vQgyFwxCB3
H97ittbXKYoNdmnij3NEWu/gaVrKojcfQnBD85vxzwmBaTCvoypb24+gTeloB2PVQ43C9cCWv5dt
Kjozm85lI1HV2GnwWQCYUKCd07ClALjt5T3egEe3596H+6eYFfX5zq5lo1t18ZONm2tbwZLZEspv
1Ywp9ACymXKsm61ubhN8qXOeYTMvt0cv+HLh7m9ZE5rRskwwIB6q3sX11RPhgjNCnB0iQO0ai//K
itfz5dO937VsR/bBbVYEln2vEno/gvfyAxTuuDW+APVpFuO24VzVAx4A25oGaKWnpDEmOyTeNRQV
IQGW4qLqLCxULtXoibEak5phXq1JzUnPQvUiASv4Qk9eLRklMvpmxa0RWLGXqNAIPAqx2JU67aIC
Cu6hah8h0tz8euQkN8dol/Rh+OWbQuhqCrIMsz+xA1S1KvYt30Bo6HpFnHNyHH78Ga1bqX+gcCAT
9TN+v6O0FkeCxw03AdGST3jiU/Ixx/Xt3spl1Zb5qQA/RYHSQfyk4OxdCwafV+ituJe3+/gvmlwQ
w11VeLz2+CbIJDK5hV09agKRzS6ZXjj3/8mTQd6a4TsKd+0JLMd7mH7fDbD1oHaTqVsEuENZnwlQ
HPZjW1kNjNqj82rEQOWfDhc9Vminl+ltgtrVpsztfFup8ovsS6b4URUDp6wGX3H97tGz1xxkJ6P7
wNIGEa0bkZOb2C5A0kPp7wr6LEiFwwRXD+8HvZovMRdalybYw/iryBXogE1Kip+46GrCvNURi/SX
4TH3SWM75wgA8BJ8VJ6SkhGB1nNIvpBOtVm5yRL01CKzIwrFTVQhuEzwPxkVmihYefpXX6nWxp5O
B+AQ6oi3FGzELh5FyfUrlPy42ak0zzV+zk8DuhsGHe3VJYna9owRwiScHKlK9Qeh4hsqjdNxBc2R
loxy8PJEduNR+stvJUcCcT3khWpgw59O/AFox2DP4CP0R/vopH22k89hFm3hDt9KzyQN/FLABWZb
ShQgL7ZxU2V1i/f+m9e2BjjZAtddfVGz4liGSpKlZOM/+20RvPpxLibN/RIpCITyujoGsNstJwze
0GcFXugN68YhhBARQ+/U8RWwi6skjs621JpIBxNhz4JFS+6N8dcY5p2iTEnofIOySUQWTH6vqcgC
zV0RPAY7I3is69twtNxzePk+osbwoO+bFcDcb+crE1Q4V3Iuv+aZB/6jQeICZDT/j4fA7BVLfwOv
tJ736KBgrDSllMXt/ux4POOk6NdjsB+P7aBuQ19lK2u+N3q3+jRx3teF8Lb/VHd0dSg0oOpsXD/q
PsLe8IB6IgeHnjywgYBX9PJQLw52aOfaR7zz3gYS0SgM637wVk1jWUGyhfMHGC/bolHt9MnzJduv
AI4RDcn1IbARXo6RGzjo5qeqkMEt5Jg6PHbhTdXobJLcahxZmc9IcbdGO662JbXlJyxmBSNab5xJ
Uyw6LyM/2S1Kj8irOpm0WJHUpQh1ZlagOoJZP5C7Hy7Kc7Cq7DYQYFphKDy5ONy+lQRC3uiSjmVn
lcb2vKnaxdAPR0K6RSlwby6LB6tAEn9/nNSfg1ppZjlzZj1u445/VeYO12R1G6f2DYKr6MT467Bh
uILR1/IWKA5c8FPd38FNldXCwRypn2YV6gMZnDyama0Sq0Dei5Z0Qm/ahlDoYtS5I34GQG7EbFq0
pcVKgx+aSus2chROQk+xWlzZndy3IIBlRE/JumISU96uDQQflPvEenSHoJGvgN41f1sQGq5sUxiA
Tf/l5oSYPD1rBleKYUDrH51kEz8hmFBY5rgvmJ9fs5Bb2WCFex8NavA4AoftOQlaxAzw//HvW+4o
I05y+24UtsjSOj2Qd4uwSI2Ko9VlzYW+eFX4THJx0FS1Bk3E4P7O/Fjc4apw4UFJ9ONUbmAZ7lEz
sF1mxLmTF2Aij1JJNE/ShoNHNLbmacH7fZRjGCvvNFjoanxYtBTGEI4Yip2v1uwFw+Giv/IZtI33
9XaXY+Pl6wJMVPsrz7T8YflaQvr2idb0wMKDKupi2QFRKYbjY4zXRbXvHted5bFrpSPO3TKgSR6T
BcktiknSgybg1fGUVT6s080BklmyYWqm+mIaeCcKsJ1UiVNbyl1QydGly6HKuGYT8lFs+V5OPWFW
2NQhBP+ZC8sAbfhT2Ri7iZKUcXtfRM42HfyE9XKgFMz5TqpV+PJjcvPUYYedzqejxi/a0PVGPItp
3QGGaB+Kb5xCDPIipfRluu4MoqPRwvwCFJ9pqX0fYukB21GKD/wdqbCnhOMVu10YkhczCFPaCY7j
gug+mYHkkERkbHKGvhHvUDkjzzGzkBDWO8IMws5jr6eYieZRH4NVql80evyN948QWQxm+mNAvoX6
pNWFVDtiIZJrCYZuZfgepxcZnW5z0gQsZuZeI5a2HkQ/IF63DwpYTuiOAoOh65sIpgfHYVmPT/vg
eh6nINx9fNbHh/raW2db5ORDBeeG4V4o4ar+VDjIerJ8ozu6GhpCHzH7CJfv8URi7uCS/78OooCY
LY12PwMpntn6/oZc2RRKhi8h3LkzROCfVg8CCmI/ywG7gtGBgXJCOFv9SkIXnSxbUMM1EknUpnff
VSFxJSQipElZ9wkiHjXv1ZxQcBZb3NXBa+zjxV0mzPjIpxwMNOgkeSQ+g6ONS5hD+4qUtBm8Mr5I
ww5k26I1SX55py/94BiYfa2f19ETIbt83EdJczJ4sCuOFOvLDLGExMyoYRX04uKLohoqy6OjNTe4
yIQ7u5wRkj7/UFogN0rai/CtYguXiY+6+/9kGWI87REvN1FqyXXl3NPTcY5PrWsvFrHtO4UDVsQF
OQoN6OJ++in4QCEuRDNaADZlk4UGcJFirhq5skGIMHeBlt/SomS1fF4Jo4ctzorlg3tayz5pOjEr
mamSKYQW8sTetwnX6aoAQJLIwIskhVVuXTDEsnmPUB4FPBdEQTt7exHao25zit5eGph3K81AxXL7
g3RaSWhKP8jj80GyLrvHVUL+dTnVJuAX0kl/ttsDgQtAqX7eQSZNo6ZgU6IX2snO2DkPB/DqyOPf
bI4Y2sRbVd1VBRWobbV3Rf4UVrEOj7IoQMg2y5DvRQMHGf4zNgriaw+YoNB8dw7Ksu6fVFNWVCdh
rfoIZWkVQmfxh6j79+ljoEbcbs2jMmB8G/7NDSw/lw+oKxfzLKD0VBeKD8P2laTX7ir/TBlWTEtk
l2t7ngwKt0NtBdZo4MLr+Yl7FYS7h7Q4UwtVwCp2YppERuZapPa5TVXpCwi1lcJFiId2mXVyYQxA
AvuH4ImJ5kCKULVJPXacLRSP0AJIi9uPg9NCL8ss3b2LZlNdQ3fJR8W00UHgeQ+mC9IK7RkKoXi6
3d0CUoQxydQIh4cZiet8ZF+60FnwB79Nvw7Fukc2tSgJDp2PIlh9vWYfOaDCsr8xs4JyjEl5YiO2
o59Mx7pq355q1ePg2OTz7jU84EBpg/1sOfyXhZbX3taNiALGbSTJCnN3kXpyxgKup8duUcA5IONX
usc9pwQKRD51/0R8h5SxEu9+UDvW/oU1wh6DY45r1suIiXiLekl4l2BvcWOWOi9rAySJMGw1bLer
CEboGOPta3Sj0/bsLmI5ihPMHfWQsykuiVYq9hIcXBzalXHh3B8cofVj6Ub8vVIawMuNLZWpjNaE
0+zKMm/fjzki5WeqNgBk/7APmEwNKJlUDbOYleBNC0EgQu2sm2ICWLUxci7fSrSZ5WRNXaPMVIPm
Hp/JwdSNOSMY4LlIuOoZPydmlHNb8lHDJY8M89exetKmojcooqFpnsMGgy07B1GbpNi6xO0/NcG7
VDwNd8PmmJmVgkw09zx6CRyneU+OB4doQAxmn1YzfUr5OOxldvbRBeAo/wBqdKXl6Rpr3n9mp7H9
1LLLGS3ttKAAz7BxoKYl5B4JTvKpRhrztw6rtq65dpTW9FjVR4F6Hqx1G9QHHEhBOLXBGAa6yvxS
gcmjvAK2rVK4fbwoxg38wxHH78dpKywHXuphBBkq+SlOUbBD0mDkcYwQF0kMHqY2qf8W+CD+jeiL
bhnM6/I5Qf6ZerSQEn2DLKoNIAco5n/PigR7WbtTBlPfnHfe6ujxYpZxXvcluZNEEGLXSZwY19BJ
J8e0ZcmPHNKOfXHPOqM3YKy0uYDXW8q4O645mp0jOVOSoCAaxHcmF9WA0MMoz/OLJn3A3I2oTRly
Pq5adLV86uQWgH8CKFlAVjg6jNQqvTP2dO14/sIWw8RcYMplmGnaat7sd8Nz6pcHWe2jcWPcsJIS
zyNAyZWhqrcEmwZ9uwPKh9moFLokrOdKTuG+Yq8ZSv5Utf4HbACE55/Mlyt4p7vqc/XkSRCPA/7a
XWhyEGU2VK7hpG0L6Ddk9YdphSh4IoxVW00Fq47Jv4Cbf+oDF43eA8e2HX+fzE6RsBZZG6rNRi2p
gGCKD30oHjT6cDVuxnHgbHmoA/OgDqOgc6NX6OcM3JhkssnLAJvPQD6fRZ3nMZK+YL34lPFtWZl8
qKhxDYC9PVfkoXfgH7ikJxXgJwpf8FntLQuFJ01g+H9EBgV7oyJNopwDxwdHKOiD/bhZNJsb8SrJ
O7eZH1cTm+mupPQ3EaUsScMkklDYPyAh2PKQVgM6iJLP9gKxhvD4CfSIlquj1bocYDgAmnv1X4Cv
P0Cq/DbmTKsg5U1oUHyms+fY+8dg5YnA6nWq+mcoOfNzZK9IHilWqyaSkSecnu4dOGwwqWxDS1e8
KHdHfKLooA8dfPRf86+Pb2u+lgK+b4XtsdaVASBAgcCw7mi4wn/ZwsZNrh4kQ+zQRlgb8GqTUyuO
w6Og7H0dGkd1Ikqx4cEAOdYx5PQMJ/VMIqLCzPWbTDMV+oPnd4Yqnq+SMBsXS1NGanUNcv1DUen+
uwtnk8XYmPYJX7xKb2hgNhQWS+xfdFyfYoE9NVOrtRPl3NmCcHRDwPCOumHUuMu/jCsDpjau5AdM
s4u4q575QPsfdyzSkNELVRVAdkfqzC/d7YYB/IBFPHhdax1Q2oDJbPXM7YNV5yw+sbhiwSGVtOxr
NR2ss41J6QOZKI/z/fj/ca9MNT2Ybo9sJhlnsBCkEVLFrpUoaZQ+aD+aTaaC93lv+cq26nTt+xme
uc+rQ1Np9ATi3+TFzqjOSK8V/HQe3L2cRQGvVR0NvamSocmF8zRHGPAmLJfyQnyoVtfGt1YNkhQ9
4uOqsnzJPwcA5wDZfq30c18miI7d3GQtwdcDig01Zcvmv5FfMEM9HZnsMzsSjsOpvBzclqG0T7/m
SjkwClkGnYw2q6xCnLkITugJgNlTvm2urYfSZnWxvUgD+NhauMzbG/KQCCf3YLNrVOwwj1VdfDrK
ZGi7DJE3cR2Bkat13WCv4ZpUfXzgYjBjPDQdsY6QRsqgQDuiVfBng4UVwEhmxTrv5FyM9wf3j/A/
MR+TLIOr9xU1dR0eczMWrmvTG3se40SGcR+oFMnGE9s4T1MJYTHLXcc8ftYAfAC73bc9h7MdZe1D
N72RrJavLEUa3IxSK+RBeHk7UAAYlUyDOwpHq82a68wY9nxvn9EzBeGDyXxlkZBITeAHfsMSfWc6
HRrc3LZJYrXhsPwZQYEaq1Foz5nfQ8X7dvSjx2M2SrQ51oFjB9biZaGpncc2h9tEH6k7Lcqq7m+j
fUj2btEWqnDVzZamiFdMJal4b1ipzJWdGNgACRRc9r6lopgx8g0F2ZdPkaq2uAxN8WudBlsMpkGF
HOWuavvo+IzCQ1is9UROPxxchigzIE3qLGAFy2e1nLb37LS/BUmBZwLEjWL1V8BJ8ee6XC5Bwccx
BPmj9ffEfUahylh/78epiQ/aPSTPK3COkNXEiym6HaRHuUhELvJ4NroM0zzON5yv6Kae1dtEpkxB
y/KYrYu7GV64Nk6tNZCLWRjTW7m2ZAJZEqZ5OPFbNtyjoZVpY23Rt6iXzsL6QXrzpc6Otybiu7W+
8uyiI40XeGsRFYJDH5u7vM8i1TyrKmmhiml/3x5Kb+5OYl8F9EMVR7JzSaJhjPyOIJiIRINhgHzr
C6xLVywgDCGWuCa6/O9WvGnRd9WmkXMOQfmPr/HViX3Om5bWvlRw2RNlAzsaRehbqAnzcCno9/5o
I0tXh1Bn6Hd8KlQgQ/vC7S656s7JAKAZh5Rs7rxC9aocaNrcU0mbFPswJWQR7Rj0/renWxXwkBb2
UMicEM1KwwLFtDbppvh1+ZkN03LmYs6yXNh0VqeT7rKYiQ4G6o8hwbAEkP4TeZaeAeD10JOJ5Ggy
52FdWPKbIfGkMCfhbJ896XR4Qe4ghZAqalVG24zzQfvWUQJ/7qXYLfCmBbCChxKFQJr106nCpkCv
IpMb0AnoPCcAIHr5LkHIe1SWFglfUZQ2qQbDcintPyFFyq4sWCCT4VCcl74iOPYh2X5tjUtU9kTq
QaIGFp7irnZCPyeSskdpevkmOIQlv2G80puDnSauiZ/ZejUcxaBwdXuyEMtSpcUch34uMFryrL4/
f5a7rREV8CWxExwnlP7aTKpqnRH9yfRfVZCeULJAx79Bb2srYPMcrgxCGgYOGt0voeGkNhxxqI3O
0R4Wlb/waD/VyKcmvRH5pmPOYlh6/obXn3eTzDS4aX9ShXh9gig8i3xy7YyaOCNj1+hzSLxExv0U
d2g8z6iM+DRHN5KGnc1O/Mdb4ywurQe+wztZNpkHyz8eQqtpm6bFifpr2P6P/ffE/e8aQNMhbJ0K
mP2OVVxn6NcyQmFVOS5BI8assEs3+uYzD79LeWYxrNkiCtkY3+TBDWUbWpQuVKshbj7hozQtn4Ue
GviKN++Kis1O8Wh7KIuQ37JoZQiR3mHzPnhwlAxDHv2DanjaeJt6DLw6QXcOP1RPWcxbN9EhHUAG
9M37BEUCGq1XxPLw26KHSPcLjnoUI7fZ4YPCRkdAPZfx2+rY5QGGkyvOpSkgkBvahkZoHMExiNH1
KuZBCjNNwIw0V+xdl6kkmOOSD3UAbMrBCvyUOVZkznObp3EY8JVBFp+vizCYRdYdhEanuAK1ZVkB
m7/pRMWb3pfsEo74f/gCa0ZlQkg6AYeYZd7SK3S/2rIa2X5EvyA/K0tjHuI4SRwkK0PunIzKjA+n
xQSxyc7P8gEBx6Mhlw8cTzx6AxciY3ZqC7Ev1KsEeBaot4t7i0LgKdX1UNgFWAmpZWMSz3OoMfre
/2kPsfAVOIRo5b+CHCBx0+oBVa6vBKw0s1Aaq4tKD9jMqjlsT7ccI/Y6vDS1/+TZBChqDpos753d
DNuWssHnSINIp6APytm6U9DiGVCwW1EyUZoybff5YfGcuD9xkN/fRfMZbcTn4fJLVjp/f8Atqp/d
nB9e7jPGdBACmB8LFADkN0EOUfwLxe9hNlW6pfDhc1YZ3XuAcmGyRd/FScvt71YytSZR8RksRSvf
a+XmoYm7047LZkU/fjyUGSAPO+Ek4bcEmDxVdWjXdovdKMQxAjdK6xs65k24nCJbEHE1BD3JtRt8
60aJPOxG8TIyxN+lAdINdT4YkcSPzfim562LA/3DNM/YmDxhLew7pk8+sZFEyQlYpUzDfq9z07+V
SE1/twi+uPzuPJSt8EI1hevK6HNK8jhRXnQVmcoDwU373Ks/aaiZV9/uf8tTi5Zlq2l+scpIqr/5
3DRqTgF/891u8SeaTKVJaT+ouMioG7Ag8UhU0NbWtGu1WVI8qe93ai9J75WoBKTZGF8toASncXVY
KzgsJ3RcuQKU+mj4qVdML9LQd/AIS3l4OZm+zv3tVX4bACjKh3FMatwMS+1fdGLSuBpj6q3XLfmA
9J+8QSAWYfl11xHHQAmqSJyVW08+kzgHMSWASwt0eSGGVxY9tRHKtQbJk6LrXaphHMzaeLu5/hqS
gliPGPscFqJeerC2b7OmlsDTyofNh8MKrlsFFtx0ZSY79Mdf6kOB7+3qBsfw82OodRhdHlEwSnUR
d43YvJcs4fvlq4+jgVZm4Q6rUxT/QOb0/ZLoHgBUdQ4veke7C9+M+K3vaHaKWq5zQpOBdLARadi7
BlkldXfz2E4PqBKlrQU0nsqyVDkuFIeRLhz2Y2tBYvvo/LxBlGsHc7s1M41Y7BjiGthHzJhHRtq+
84U+J6AMnt7X6E6gF73FaICmojMVS59QUQ1FQlkdbqkVmZCg+oOfSLKs/ihmPgDmlUEBr4sY+qLY
MEDo4O/tTynuIy6lG+2N6jY/e/QlOB319PD+Tiir8YpbAQjiPonpAYoj2zJfz51Te/FqRK1xg0dR
q3FQVKnXJkpeYqDlT2vO0AoyZNYNZ6b/HoLPT9yuoFmry/ScLyd+/BpckBMaQtxwS3iaSdm2Fl13
BmC2Yoo9JOAnsa8AXUrYkWaOVkgiu398metl/ijGoLfUCJCUeLTAgg8NL74tLV9D05fsjnIk2HcL
ZqLQlYuHHGoBaWKC42PVXmVANgLnoprgaJiTXm6XFowFyi5IU2Pt0QHcYiJmc00k+ZcsQsXrsNcu
A+u0cI83iypqodLkLRN2m3Dl3+0hLTsti2bSuTAhMJ6mDtjxOTkotT3uyyLCN3X5YRlKMM7P3sQM
TptRYFDSqIbun83If97BOToZJxcBTVbBV2nKN8CFPdy2QyQVWPHdG4f3ZRJczmoZ7UGlH3IoPjXB
wHF2x6SuM4YSKv2QVxZc9JO0AKkINgchnNaw1OnWNhDIYtJIf7yllInw/2R+41GUS/T0gGq56QIo
fdQ2pVGWaSOsBB9B3YXVTwDr80FwGuNl+ni4D/ky2NvqXsFDjtD2d4sT/ay4i2E0j8YTJxH3mDN8
zznpfyqsRio9G8/0iB9zuOYUzpLschw8M9Df2bkDQc9uqeVia2rzBkyqpHG6oCukshZj//E5mfb0
vtQrY6770AiUgnwIlg/totLIKXpEJDBeH3ZPjJYsWe2J6XEU0QuvjeZH7heq9qdLdy7KI3stZp6B
lDpLpjEFZqSzRHLfFGdEhVeZBnxdzDOfEyhInTIvh2IKqwE49kYCXka0yZplF3d7Ry3bE6y3n/LZ
q3WQ6mgev4Or+JKnNWdfCIhV/nr9UNwFR0ixMlyuHXvIcDLK0/JrojW6uHje7zmcGhXuggMCxGUG
Dwm0W1WbfNM75/RgAwxPGHWpVPkv3IKaE16DgEESZPIMNPnkCC+uKTUm88MRcVqbJh7ygue+0xOv
7d/N3hVlsSmGlBzKZOvrFbf8AUc4L0/i8TNdBbRVkSDRdPGVHlK8Cmbk9aPsIG79JYrE/O5mdKIF
5Po9E0CY40+JImAIU6OCNvLA2/zQMGPVwUM27yrSTxhgT3c4FhyG9usQkC+6SbYBnN0OQRPWARNF
F1+Rm+zZa9gKRdta540RauD61nGXmjRKKcJfe++DZa7Ccm7GZGM2Dn1IcIVI/evuTqlHqrLC1QF2
qFQJQlAUJHQa1eHqQXqMICUn3IG7wZqroEccXBlqWl7H2NR4WBpkQ0szdMXT7rXBgjdkAceDN0rQ
SY4TbhrBj9lnhcK+Yuew+PRM8/GWtbvb/F6wG4YNmBC1HTB8r5wWWxPJfgxySKRGBq6YAbc+410h
INNKMBuUEF4Xs4FLaCWO6mOdHqFjYUd1soHnWES+pUVy8kFGxu9RSzwTrtR3FXsX9igQR6rfmX+K
fibwmjAyQlWeKi+EVjchUtTj8VqrsYZ6SG6Q6Fsj94ldPXMacLlDQzh/MtF+wazdOfxyxcA0gN/n
mrXQfw30m0FzbAL0bdSEQKPM5yKRGiLUnrLliG5aqOuHMQSv7/Jm4SDtT1EZ03Vn2FYWQWNqadBc
TKkRvRofwuWwK82swChqvb+6B9eYwk4huJradnigkiqpDuKsfn87ip1Ey0SdnyHi3MW2h8Hk1/X7
YqkrDxF0fLzThaeoNPMX4Zuxa6223dZNnqQOi/4RKKRAY39+2rihN69LExTU8LggKeHzoos2KELs
ZCOYwYE7nxS0HO07mhMOqXp9ozeILMlyDF2EfsRhdGEwU4UjwYvKZXnDge/vTJsTWYLpiw8sOpqy
h9Ev0ArekW/qpBtJdEaH2ZfqAew8rKyrtZwvWXAlOBqt+zeZ76VvgREbFQJfVi65/DcrF1g7w4Sn
nmo+Xu2L/8t9p0kZdhWhuGZI1UhdldvknEgy/KdUQCBHUE40TLhzi8ZRQYsRifehKbz8v2TL2suz
iU9b1ceeaS0GMkeqnxaIsbBf2KGu+YDVDb+PRlWbwllFeEY6c9DYgiNp/AYoncgdYhNanzR+IfIu
syhnNVGjbLGhOhMxAFzovOtkcquM9afRc/lnsPKMgVxPadaQpISJE9iSEBuJ9VHJ1JwDA5z9Nx06
wl+b6wCWdvQD8iuX8/BQjLKuD1V0FwcL/LspdP/oxeYUUebM1iDMEVgoPHJLXKHOZAkJwR6AV/4e
LBMVH8PJ2pfh38yl+6a4t1Wg6EmJYjs5Ok0IIfn/0oEDQGsMXDX0a8WH5Ff5St/1HvG1u9PbnM1W
wGhofdLm7dKXnnDTRjo9j/DZSPWW9EIqnJWcXdjxPDJExNMwOhOY3of7T6vCFh/vcWbeyGMSuEAg
Cy1rwAsH3d6fymO6xUgNQixa4e9BE/GkYqkSJ7De+ngsLUjaMjNSqh7UvR9q5n203p5PhfvrCvQR
o1KeOyRk4v3bAQsOnaYuEoaQDWC2eRMsBEGq09WpkknEEBqoEpOTnuIPq/heIW2prdvXjeaJKZcq
K+Qe1xhli/N1r/cJYA7GrXLyDrcDoXhF9AaMS5EHbE8Dvu3KMHasJpjFa74ouD4v9c1kPk6NAZTb
9bo4BP0mX4ylK2uy2DmKzKw0uYZV2tugwA+za4xW6fhJzCSrM8esCe7mcIGcJVjEBPV+fHoZaBo7
XVEkCTDKy5oNn5snuP9iDupKzZnz8zRsr/Ctk0jInCAwzmMvGFgGZhDJMfvRUrzMhb4qT3dukiOX
+Yw85kRC4/0sjImeEA6RNgblEGY+cMeBFKr35tbqMlU+aeI8E8QNKpBVrR9ZBABFZIpnR938vij8
nDTS4O24m2IiO5g2esge9lSlc14xbTZtKSSyz9C8aWVhmXh2MLtDhEzf8ib+sN3QFF/yjLs06f8d
Dx3kSt96DQjcjoNZ5czf9xISwqCBTsXR93dXCzery1n6kVyQ9wJYkCWPU6K3a56aQUu+hkpHrteV
rzqDU5s6AwyCg3cKFXl6l8pp+r30jfa/sIYanxZJTJMR8BC9WrAVsyvkCP2NQDWtPw/gAXIJVXo3
fsKzAdm6FfLXrUrcn9u8tzXrTp2yck4u4UD9vljJLHcG1ssJhwJVmV8MHosh3/85fIujQei/Sbl+
T5MKyVZl0OUWYbtq//LXbrqc+Y0eILEEjhtTw4+Sfyip7emhSrglZG7pbENghmxfnoCzrr2vpRZD
esK6hgmYCg4nwHFuAUL64CIMNJ0DNSyYE05XMSQ+0zPE2aCVMWRvhuK/oEjutMqinrMkvYLBPP9/
iSo00h8icntMjzAUWmi1K72uSGMCZokSYPr1WWMPUONO6c8MAnuzG9NkMGdNqbgHZ95rHpXfIjXa
TCg+X3xCxUdL+inAGhsUo75uyLIvKQ9Co6+tA4jVDaVWnvURMnRcLXVhr7ynlqIPA9oyhz+vprtE
EE2KCvpQOfoAEAOaohR1rbmEu534E8BCB+M/d52viLvq+rkOgHHQIpsx/RAsZALWLozXvkfEGMUz
hWHEcfNK/7oeBqHw6vFUG/DUbM62/2iIiHUoWkZBUznjfwSx5sBqlupDbZvvMDMWdGta/mEzYxp+
K8ZPvpDrAM/M9/euTswZ1OPg4PKeQf3mYDLIPMTFfMLe4/uJpeZxawm1pAvgtscu0q224OP4neQj
eWUrgP3EtllNFal4MImUGHgszJSKTmfNCBt+aeW6YigxegKlISF9D/klK9KJ1929qkGhbsfxK5cY
DMtOlecBE2zfg5qiU00F7UIQzFDM/LXpn3oY67RaWamz1/9fXbYqTTXbuh0WX6Hb3LoXBqMN9o2f
yCK9jPEqjLWJWzDG8Ug348U+HmL9v4fW0z2WJq924R1RweQ7+jbxqYIZDo702y/5id0vFXAy+hOA
q3asvshpm+7Nr3n2VGiWqQ7GaI0TH8hF/OVrr6SVrt0M0YNQeH7oN2A06+tqOLk1P7/GTxR5s7Ox
bAcbd6OotD3nWAGbmoyLTxTq6FfxnVizwnGjZCAv50ymX9i/aNrMqrJx658mw8koYYuonJ1OGm1v
OfqklOXLsz+hHQu4ezhUIntI1KWiMhMQ7E4REeEBJluDvfRZQkgLgpzs93OgwIsgn9JMDDGK9a/+
u8PHr8qelWFeZzC6p1qE8kNMZd9uuyeJ8LIncAlrvZqAcfGcCwzXcMz5Cj+3z/NHPqrytUiA1/kF
S43QeMZPl0KAMNHQz4vu7Z/NSCOSFoDVv97u/2Vh36cVdEqEMsScxjSfupms1fmxYvoseC98UnST
cb6NH9ajF3P0Bl+2dJZeBlL4Hc5jkv+SfLi+JV5KPZ477om0o1VGnVCO0OCK6grWGqLBsgOOrh3X
TTuEi0DaxT7Kn7xVhPzOMB7wwXiUuXUZjHnJIOVXxKxRd7mdm/yQFe4HgEH4VoVQvBLcL0ZCrQhW
fZscFRlvMgp8/Uo2OiUI0k51FgcTlO11MisZCzZ4xp2LCCq6IhuqVq6LxffW+oKf78JtsZbI1pkb
RtnVJGOwVE8DsTDsc+Mxn1MWlzJ4Eoqt+J5LPdJuGsvshScrXho2NKf5VnCtisTc6c3Fx+i0IOnw
KV+D5KIOLDtXUMjCzKJcwUcDLBGkSE/5UKVDA/uZSoibu5fprIG8Abzq8I0XjBxCKG3tgy2FSKnr
FrH4P4HQfTSYh3q692+Ip91DfsfAzqrhoHDz7Z50RqHOsjwgr31ymBAUI4sncaF5Plyqgq25uCrH
UgOt9WTZsxrUpzZrdlp3e0AkVrp6FNaZEGLFymuc85HGkrO+YI28miBgJieuM1GNNj339QKX0k8y
OppW1kxCAuboFcTilHLGXARThX5QrshyOto9aWyXP2S6FQsH33wRHxFAf8FkZUEB8teauORTU6wK
fDm2+Sl/jA5QUXSxijG7O9dLjcRVeDWiQidV8PvH28dY3TuTWIpoqQbicJgBx4sdIGf1Bi7m/dq/
sd1TTFOMwq+651u5H16UY0J+JS4kYUAbP7DyX3EDIQjBVTWVddknrPOUlkG0CYdyS1/8CurwN0tf
F+nUCfgQszW6dAiPZUKRAco9om4mUppEdccp4XwfYbJEX8LrTAoI2oP21+Ha3ZwoPhCtjR38n8Iw
60WPd9jTuSwBvQGvpf25FkW976Rr7+oM6fiZVvA83gKtczIk/4RhSK8OfBcwF6X3uBQfXc3sKh3E
TBSba2LwK+H6Ku9aLPebLZtnV45TVR2eexqyM8i2mQljCHre6PDGQGdu+mvTpd5CwadhvKAZdy3A
GJFAbhWkBXoxelQSWiAkKcOzjwLZNhEC33ck/KbkH9kxp0wtg5Fk0V860pBEEqRuNIZe5Y80pAXc
/lDdRoFrB1IT/ey3oDKcGcT9+qSOKG2YwTo6Ml8Wc5+CGNW82OQ0yYNrViuir7LzcWRLlaBkQvE+
SZVgfek7r/08EN7YOECvji/hF/nQSWT58P/9LQSvcmsynYOPE4vxKiDwN1Sc5N6T9qwBl7eMI55T
YA80NrD6abb1qfG3drDVDwhETJBoqvmO1EGIKC6/+0cGyTJUOXgSgNXM1IcnLfeOiVntSo8D16m1
5P8Xon4GAVtDpqGzF5T2x0euBlnY5o4el0Nu5JyKosc5qHaY90MZDq/GTn80b6RnAdZloEqqg/1P
zVPdIGfN+IRd2ZKJqM0oI5BPp/4ZzOz+1XhaEG7pQuzkparVw84m+vBVEmGmMEtvZ4lBbUlfluS2
0NTjjPLAWF0JTI9r/1s3XXMMLEzt5zuNs+WxBE7keUmlfozqBCk6zh5lUHeNQaSxNSID1wrpf3Jb
N0sMyLiI+N3dtj3/uF4mk4Cg16C/PPZ0tPoiQ3IfOgNEyBNwQ9ZAU81dr+Y5//RXzuGoREj8CxrL
npfeW/DgSeOscljnfJc0GGRZ4nR3o2SErYxOuIVtigGzQNdzDggFPWTdJBmVN7fvoqdvFmgzwEfR
5Adkd7wVJmys+J6vEEYySvSECKbYtFMxcEL4dj7tONiLBPjVueUnGUQaeqnfPS1UOHOf+LgbPzgI
hPEzxaP0h6rusFyPPJEBN5RS/9s3bEUb9zk91AjxITcLb9i+EACr4H5+MK+L6WH29JelZKfqm3Fg
I2WiCP2R8xJA8l7xpInPjDi6F5Dt2z73KKAgh7/RiGCJovT9vLbS55d415fR8Hnua8fWHohLOcn0
s2PSQH4jYcnrRMvhEThe1/qwGbBXDnRSnzQmQC0T1V6EQRrwkqgjY6vzYNkPY68i+oa6qXs4gPbs
bArqrEvFJJE0mAlPDvgyE4qXn6CmtfImZ4cs79axZRxFhvdg0UcxqaE9lCVq4PAB40d33vcm9m1d
7dCnL7oAHGjNGSlE7NX4vKi9WrUx/GIijlrVXHc4qoPyFVFAmtdQCJldrgzxtTn2GASjJOudeIEw
sx29oaQ75Kgnd7ZuwJ6zwyeIY9Cnijxhi7dLLhHIWE5xOKzcTbvRn0YCzcEEv4YAr9bzrFIaVmY5
1C313xLdtfkrRh0s2WIQMq7QQBdppVlgfX2hRfRC3GokTDwn5RzOvvLiA0tHNjNnE5zKbn2uOES3
lbiNOim7JvRnQZ+7YwUglmNPgGUZREglRALEQuhk7HMQIWvHP0reM2DO8q/tXgHkSmbhuxoivpAW
jxk++fGQkrF6DR+4vzhJQIuGIZk8TgWHDjPhz7meNx1qvXwuhcm3MXPRxurqq1oK70plzwS35orn
CmqsVKhNvRby9jr5WzX6Ly9uzzZOMViARkrbn7ihHyU2YB81kF3xSR50SiDBxIpUzAo3aEkSwyzl
Tn6Sau/32z2k18+oGcK0w7Et+7+c4M8AHo6gqkWmtxNHEiuhexotsduYs/0B+Out/G5oaQ8wNqPB
wl1TA7weyGkUau/dODmRpwT6Sk4at7upwEhvwzl5sXMap0qD+2mYWuE2HpaBf1s5hvIUOSmZZHod
L3jY9kFkOCtAm5LvLFSMt2yoqBGsxPItg3HW9h1DUlF/0gSQYfzmISGJ58fE3qeWKJ8IKSllSyU0
DrhI6YnRY2aW5R5icExUp98nQl76xOB4jiqEzjgxlZ+EeXxAMIAAGnImCCQLFx/IpEUlqG56+ATM
6CRWkquyqb7favSOmwniOdB4pr+aSCHnsnj264QOgvwQJGRLaWgVf9Yx1+jHXfxwVvkHZSsQx1j6
2wdtryapyefpT8qabGXCJaekw/zHZsLZNKXZgMvsvULo88jqR8HMZ/cdVvLeQW3NWHVIaYvpTwl3
INDKJD2ITetsqFsi66CYYbcTV9I3h8pGVXe5XkRZhMswJXUVdg5UfBVGzS9sngJ8cYtTtcnoGmxB
YHEKV3k2vAjthyVDyD8iRx57QxDt6LG1FjRxkqkt7cWhaNipqxCGV5bfpnnU7B+VqrUSxGp8+zQW
nae6ZPd2FnpsZdycRkW7Q4axp1lPTGUyzCvshBznrwdBhjdpd/ZY/e28O9nEtmtCrtbGchafKQE5
uTxq9xzByaKa0kdA4p7hOhSPky4qxVUl+7Chat599GoaxpsxrouDNvXqnoxrwiestJd/xTg8BjS3
l2xPbDYwLxGY9aFXK5H2J4fHYaPBUgx34pT66RMslakptIeNyNuVQl1OvYESpZbbDv8vOfAuH0zn
sUcxYipt0VQ7CCHxTuLYv5lT6bfQpCmmY9nskw6nWF4+wB1Ib/be+RQK0tfpFPz9+9O+16AzrFij
GPlxNoqlgkW/j6IzVHhoxbw13CAjnqsucD0ppIZ1IMvWeOT9or+Wm7yBIy9F8nyiH7tmMBD0OtO0
pw0fER4NBLY4eeo5l0IrHSgsLayhTqv5b9eNb2aLbVatHaUJqbOFZiSwUJoheA1b1BvHInRvk9ip
ySMeiz98JBzn2oQRrzmtvzSCTtwNlMnvgn38EnEPWg9gO4vRnscoY6imnNdmbkaScJxuP7jOQVoJ
4ru4aucm0EFMBX3mj4++iRFNmCqF59i3qfF/IaGPpJ8dzSloQyf3fQXt8Rahr693a1o+q7GEx7Ek
N3Zvpl1BL0bYvik0104W6g7I72KX1fp2vc/aTcCYD/LsWBtwsRw9TgAMJ2BelM9KjrgZFcbv4Uf3
qa4/oNIU+N/BzRa/Andqc5HryfUGWBccJD2tyL25Rs6vVjiFKz6sRkOLgIEdILnOWbtau4S1Fsv1
VkmCmZbPQXGJkQlVM2MtnLUQqmOjr4EbSH/VVt3ISKF5Ko0fZfiTnWsik8F2qie7QOhvFyJuTz9i
Fhj/FjFBcwU2jzGNmjYOac6dLPJh7nUS8gNYq9iPCuAmWg9F40qUriTKMZydLGaPDUHTdhbw1Zay
sSbHdv1mCrPM9kRI6w46PvRNlCwZvRXbdJEF2EL78by0Pyw0RqIg6W5H0+QRjpEeYbBEIrq20yWf
TrjhoYhDFL4C612n8c5ugSri1glPZO3ycvLr+caoQaToZoXh3E5XdtjzOAHFybz5KI28X1FYz/Zx
8EwYzuDipQW+fx0uCcz5rDPBAgTY5NssvVOlJF6uDLTf9LnCd5W0XOeqf000gqBmbtjuP8ydtBXe
j2BiHS7dAL7kGTvhhVXFWX+dtvmG4rBABa+ZyPfIgV8Esmvq0WVjhsWhh/6SJI+DCFGHun2CIM9N
DpAj2pbntatv0BrDFkCT1rcqDT5swZf+9A44ff1PaokkuBBlmDtoZu+W0Xl2U1aScnW7h9vEhEDi
NNmqpwXAGkGCroQX40/fxRrRNK0LTwwI0ZJQqUSrc+lKbJcaSFiDY5EF1EUxK/qz/8Y9CANKLJNP
Ofael+YPWw6yVLLlPBaEicrFgLRgATeT4dnJk3FKwoSPJEUgXbH6Di9d670ESU5n/+C6fhI6ZJP/
0iQhpU247vG3OAXdVtYzNF4/r1E9sxP/sYZ3lYL25Gn4zmJQLbMrWMGbWc4obyz1iD9rDJF4Guat
j0GGsv56GdjlOCmNuzFaIRz0wkUJ8xL8JppiDYmmIA90cKCPUJY+meUAAep0gfXVeSvAHu/a1kFM
FWy7KmLk6RNUM+tRa++yCZ+EEuFYrzaRxK0okbDCJCNsFeVefaDzNL2kIZZa72kifm9bXofUpaXc
Z83RpGNEAI0Qe5MWWB0n7gEOBc2RoKewIWyHd5A1F4yIirFQmiF2KkvGfuu5jgLNGjWteHYusp3r
F/Wvbn0Hut97x6064/zxdZixJgW8hBnXFbmQ013AXb7FlkG4ep+Xc43cG22uxUGclJUwUSFlno3P
Sipi0gipTcVkv+QLrD1s8XrWq2et9Yk7QgjXAyhd4VaweoaOJu8OO3nobpEy4U51qkV53Pov3aPL
LZsUmsisWvNWRpIRzbQiXInRs4m7raVffOEWyfxuhby1dkiCbGGRKAZ1lSqOFb3p1Znk0hzfkV5Y
9fgRddu8fnp7RbWZxHh/qYoTmetKeav4MHdN/r5jNkWlhRiNw5yfuqG2dPf9M/NNhqaqaMFaiC2j
aluvRp2fJb3GN3jhtSvYPjqag2ORROeE1b/PA4W8CjypqecyaPmxB4wK9n+FwhhQOpRGoEyhnZRH
+zIyhWhJu5C4J5espc7KvzJORIhxHO/Fc/6og2FH82cKv2jbGrmWUiyKYfi9ZPqlpHwpm3gesR4N
pjTTblTtojoKRZWoT5UEorfONeBfkOcAOqqZWOlFZfpG1GDPjJf+ZdXI2klBvdP4sVDu99oDGjq2
aj90wmQL7GMv/TdHiXSPUU0DEZ6/txUzwVvED1ArHD8/qRSNfjTtrv0SLrZt6L0u4kdZX9VNqyo4
BZ1xUx6Ws/3Aprt0wK+8ty8R4jMMroC6UJQ63qgRcalFEWX0HrcTpceKkMNqTUxVmc84PqMIDRDz
`pragma protect end_protected

// 
