/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1061408)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/+soiblnXFkTp+Q7KTHMuXPz8TFWwO9EMAaret2hYFyPuLIccsTxuEgp
fgj4YKMZ/9j0z9ijrEjbRugCl8BfPhTtnByJ3xDSa4gOZ9vNkosbseC2TaBKbE/AD96VqfmiYhhd
6UiT9K4dVcn1Xe9tqjZUNmjhVxSueUbJvbcZmSfDGc+9sGbru3VsaxFM9ncTJxzDnfY+n1SX5vpE
kCtVvivEUl56hglX90Brt5nWCNMk2ml7P1hMK5PAKX2bSCdBzPkT4a8ngtoB8ULpu+nfH3nOmihf
JgYcJtjZIHuGTvXLcsGeVGr0b4v6eokXFbLvqPdHqdby1K7vH1NKA8a64QzzaJ5RjfSLfOKbeMli
3B700PNKhIviwSpv8b1AjccbljTa46YypMgxsb7XtNAnpFL4apO1qLeORrjKA/MngrZnfttfH8yz
YkuA54DXALws59Vxq5z26+i1qGVsshtGkomPgcn7oMJlgLPNdVGTdEJRghTkf4avU3D0wb/1h+91
tldXNugyaGQH7bGtR/U9WZUsumcc/6T19Kkfp18rfanDzY0Ocj6CcSc+0OGRZEsUtk7paj45yP4o
U9oEjCgYUCXUAFZurb83IF9Fqfapg0oULzppEnCGc4HLE8Lgcw1NdSelIU6o17L44l3ZfslUA2QF
tyLaVqZs3UvZJiikfFCuppXEnGaQc58cmjigMTWE52XBh6jpBKMC1a0wtrJxniYnzv7zrNUcEsVV
r6CJxFMpKq663lG1tUnMlnvNluO5q3g1i7T9E9CQ2kgZfWGe6tzgr2/LbkXQt/Y7zbM6tvw3xfNv
TXIWhxa7MbLED/IqMMOG+5ze1qAKGP6gazXXyGsjUYmift7se/mhJtvf/KaX/Kj067Gihnf1TFwC
PFlJp8kuwAXenOvzLa+ARAV8SCA1fpvfEUw6llNf6COAIhTIuh/Dcp3EXHAtSITIdPcePPRMj9PJ
x8JhnO82JG+ONN9nQDA3XbrLnHYRqjWJRIdY24U3xo8Zly4Sxn0R35pWZKlpdYqFRKqlWSBT+ynl
cShjpC+nEutCQOnaY5V+rAGJ6kqbwBnhG8U9GzJ/bNTGCIfmOJ07abMU3sD5pdYb/+j/n+BJu2iH
aduCPydojkQRF36beeWjOEfJ6xxLOxnnp61D/YyeHG+ZLbpmo9fsEviue+3KMS3x8Qh8osxNyu8m
TswP4KXQJ7rmro0o7rONztcyOzhmAZnFlNSVeeIuBUBROXosuZjDVcg0GpDbLZnNmO7XcOOeIX0G
Pe2lxj/FbPw1U/6rN6mA/Be8jEk2RuulTkQXBOqjXb2VHmoBHdU7ce2V2x8JOcOk9hDcwTfnwqoE
s2/jcgEVXiWQfjKTC3ehAYlL+kfwa9wiQPFhMq7+V0KkdiqofGUBtFHeCGamUzyqQpV1FGKYfHFD
KQlZ/+VzvxMCB+gPYAizp78KE1SKcN8W3oqxdY3wh1UormmRdzTH9zO8UeXewgmdMj1W1w4M5Ehl
A/nWljrPKBp1sJsjtoIpmSnUaREfs1G7XYAnrUhGxe0un9f9TmJNwPQxpNvPBA3rrULeM/e/NnSX
oWvhuHZ6EiOGajg2neCAw6Ls5YVejKKHJUn3XZYZcOWT69jbMiKScnmdEYdhzltfabY3TrTZS63k
69Q5HFDnMqVaKUeVdsFToLDq9zl9QU9oBqVsomXeRpD2NFf7wALchuQk4rYo6yD6uT3sPIBBagN6
VGFRrjHdUTmxlhEHvoHe+T1yM0UTBcg/ZZqhXZOHCSIoG2lXlJp/6XpfOd4rNlEEsG6V8QQEN36U
6TnFLpNHF2CrfCg5gYu6fiBqSTyicqT9Al+gfgCdfkzGxlBknPP9DNJS5ErN8mSzBEjeaiHki54w
fwv4ArLI1fzJL7fHEyT4isorzQYflKrYOKQM83r+gTepOJhKRJsMF/gCtbybIzJuqRfqLPCcT3O0
m+L4yUxSgsNUAIyiVzBiTh5QAe7cg+jZ3POF/wEAgXXghZOHjOA9wdZiUC2S+21Qx+SjUPvJg/ir
u3S/mu/ckjAlBfl7+mYpj93Ra3wad6/0TgCug2dGKpFFsP6eatV+Dy7XbvPylMlkTXRqg2uXjjGy
a46uINUGVhwd0yiihV+9goD9Iuy6oich/IfBrg5JLPr87lKk2LyAMkrRyNQfu9igqhlDbzLC78Vy
QiZ9CgV2YQtjgUT54wCRKtaJEQnL0IxiaLmJ6ndDX7Yzvgwrlbd22edvANVe/9O4GabHa3MmVGlk
6cwXfb5/2zG8SVsGEbqf82BR6dWv6edakpCuy1Cr0pIfLJFt4NENuNh4tujiY6wwYx1BTUtxjhiB
XqwZpHBGVpZ/zIn1kL2IZxdg2H2xEzNh7CNqFkP7HDYXXDoxNZgElpBkjljjSqeeD434Y/OK2+Yp
kruXX1QNTNIfW4JyN6vGq6NAqrKtaOEKlbW7xL3JgeGRY3w5W7z39TwY0Pij7W81bndQssugzT16
mdB2c92jfC2JSvM14/XE53vSyuHHfM3pZAfaYFGjKgN96/rOt3gdTYw/LMd10eqaWRI5Cs3FK8xS
BFolKODpDjlUDjOVI/XsWmxw8PdskuCOGvLCFfvflGNClBYfTmtL+Ta1MklDJh0tPqb+Zi91JaHf
/4gh/n9RKMDTovaEMX28HyUsXLzM2v9DP09b/XOMBfPQv0CJtuNZ8fvn70Zb6KaEheDWglxr8+Sz
R/PPLvM4XRoLMLBZLZQdV8g+XzPPaBRr4fNR9H+zU58lfkqhJ3BhHbjs14UQ9mevA9jruEDqOk0B
Bx5HbK+SBQQYxfGM5mjkjTjdD2e0n0ox6/OIi+KKDe7KctMucSsK+XNgR/L3W7PiR+i+Gsm32w59
0T6YKO6+09IAyc0COdm48SNUz5oqFTT1lRLwLbfZonFJO+wYOdzZE1sHhe+3lH2iPlq0XOBMi3sO
xGdF4928RFAL59D+Mm/j3dgBdL2o2qu5fgfETQTl5GR6gBeKTprDAj0Z4LrBYim9bFM2CfSqpNcF
RtejHTvlPYaQkx25KD0ApKLPGR55XsIHmz2ExH70fh26Df1UOl6UYlteI46TwtzrNZhGjqEfa5/J
9JfkhKAc77OUrCmJ2AMmQAZNHcuL3jeh4DQ3XIR8YLP3TnW+YQphRPKq15jvuaNBX3V+TC2uT9XD
HvYjJElAdOsC8qA0dK+2agtpwhJUt5Bcbq/GHfHKWhX9ACMDDJCdWsAoG9ZE4WSTP+80RLKh8w64
brKPmyrMekeZjn9J/vGejOFZzGDNbq+sb8U9bix8aiXXBDZblhKnz+GKz5UIK0OBz8rifZ5F04K/
HJnCHN8px8s31x/8Ifn93R8YzyqmtJfZK9DC66KNMeiwqDyplpvEKh6jUQesIsru1dc5hSdXJQue
7HnOmAnqTpiPO2+NMe4D8ly4ao4VwO/zXoXObh/5E55J8wXR6ofVPkPE3+jRkb/tf7f/v1xQXTAS
YArPycdDAVkfoDRBVUGLspQeV2r4/hX6OEdV8Hc2quw3H/bnHy4lX6tEYmvUHipZb9zTDtqcQ6Bi
zZjp5HGndpo7TlpxKnJSThykSwppfXHrIT0xA231mFNd3SPo7JYVGNBdVVEcXHAAt/HQfoud3oHr
7za9xEY2sdpHkcTtwgW9XmDI5xCOFmk8tmK3sORBtVHkIQrgx9qJ6Ha3I7E4C5ipx5ykwPd8oh5q
5taIanbz7zwQMEhRtCeGU9VOpk6VyP75oCOBG3Sqo2hsfwH0hg8a0MyA++mbcSZqmXEqrsSS/K+z
k8RPZj2a0MP1LVEZ0N7mse1dEqLD4LCV2S27eI7Ll3/KR3BIomp1OodZLtOhuiU/M9/Pcpaok4on
FWsA/ci5P4cI95eTW140gLdYRMBJ7tjrsIzn/qlivJWoNjxqboFEMUd0QHKo/Rel4ZW063QyYiLC
0r3wlHa2VWFULiOhczapCZ2iirjAuTCRnF9kVuL4Y+zLXX5L4Zc1r07qRoqStooQ4Wr2q88kgQDs
6BRvA4k0y6uciTFIFLjVbAvy34aro/SxslfKJCfpQ7g4EqmbzdNR/wpVE/qmPrruQ/j6G1cGizR3
BGxYGXVFio8EZqajDacwg4U958jBkqbG253fFaEciI59azSxY3vWGNL7OBGk004t8F852bjpIkpx
mnLqioSRz40/4fRQYdTEoU6E3BDuPk8QDnugglMSe/8OY4mzIw/y6WKsXa+OKfZhDtgjRtjJ5x3Y
9xk+L1qmSp3x6rCs2mvQ4/PCMzA9IheLbsbgXtSuKzZuHjT/wHUHbMtSl8u55Iy6xFoJG+AFMuJ2
xH9DXhPi6/i5TJvhbelw7gvrdq5aSyYx6xRhrC5s56T2PtQJvtf1naLsY8C3m0evlO2HV08OiSqZ
qolU1Vv/Bwt1VE32F5Oooqh94SZML5kxW6/883f7ZrFgLA15mLvWLgnW6epgzSaQ1Qjnshp5PsyQ
fWXSnWUZ0MeZhdeCn/JQtA8vVrmnPEKXTgsTT0qIPG3n7PYOm5Av09fVVJbYFYH8LK4f+bURNnMS
wp4ApDtuaFHM+J00DBxVLPB6xT5Aueni+/KcZ0LNvv/YmkvObvAk7j0xCVF37FNEFbhHe9SLKtvX
iuUFOImHCZZa++rE3RoltYAdHPcIoSBZmDX6vDzgh45OT25BRNRp65L0F0Td8iLA+mtAJrr/tw+h
h6yrkbiHzH2nPDLXAIGiO2vHKPSaRrrCS8SBSPTVp0fHwqm3Vq2h9aGNN7LofzNXvLB8JT5VoUDT
AaK7ZY42BAMBNhlxVKlf3YSzjTsjd4V79YAGZsGxf4iwhjiZ4OZf8atw1m2PRJCI04wjjvQDDj8K
xlHJ+Wutes6956SeyqVIxrpY2Fv5VMV5i0/Xw7kE0bFgWjmWHv0c3DOjHM1Xc1nmHWO11bxyvHi3
UB+w8INVkc0HktfRAT2q5IF6d59i9xP4W2b+m/7u3iT7MEEuG+aJ1b4GNIlY1Vd7tI8IoTXX0A1a
rFibge09CikNyVVkdtafh4kTetX0iAppGfFFT/d02fQGbm44ovAV8G2aN44gDbNCWW6oouIGGCu1
IHESkygg2Nmi+vrEZSy8lhyZWWMggQeBSWmLlUpoARpilRYmfWYyZ5pJt+VNbya5OLn8XDOtfimt
/m867f67uKqGBt3oHOoF1Kew/fierQXOnHnKERJCb6VsFhl1cskSwfrxlWWIRUmpAf6ZTT3GKxyx
hCWFG65UNWvyu36tkMN5URUSCPmuwbe3yhNNmYo61rDjTurWZ5CZ+M49QGtljPWMYMfs+irgy7sc
u9vfStNQ9bPAQTywptIMAyBjE7I/mlWY/m+elB2OY6nzHwpe6AxNto9tkKhcevcSkh1N3tUyAc6P
zpacN7NOrNJmo7VRjwVbHL7+QyyiS0Q6XT96Cj6x1q8botjVTkqsL9+G7pZ12PHU7o4/szfByTY+
/2dU1Jx9YiAKO/OBpuk5HHFTp4LMPOgWHka22LN8OyZ6mcZ3ERgWhuUHnVMFN6petYFxQIqkTCj/
kM7KN5GAbAzqrZb6dMlSbdm3LPXN+2Lio58J8x/+DPSFQ02qob43SKUq0RtEgJ8WpAhMPCUEQ1sx
BmNi1lhP4nIXFb7oyZbAoFq4PS2Qlor+REIGALjDb882BTErgo1ctRbrDmXaqy/ko9Jfeuf6S+TV
jJnrKGxCQOQqbv29ISrU7jpo/CYOC8Xm+Rs292btWa9I5gB6u1i2iKOtt2o0eONN97KlwqLPDZkJ
k/bW5DSD67Rt9WoIpIqBAUhYWye7kEquVVe5uTqc9/rIoZoBkRE2qIMEpO3F2/u6TPqOS4i+HfXU
V9AZzxQcAB0po40EzE/lQ5ghgVXy87pEy9IYgUI+82BS8yRdGZKjMPZ74cC6wkvdbwSwGaIvBU+L
vAbP4i0FJVyXl7OifSZUvoVzSx4JDFvQrzaypSKDzU7AOcJDdehbTN3v221Av+9ZsOkd1U4umtOP
wuhukWQH0pR0OpZrUem9F8YVxk+wfKGpa+1s9FTCuq+VaDPHV0Wi+lVZ4G8gFd6Nw36BjAOQH0w8
QdnertjmbsHS3AzgvOjTn8n+zVmxgeC+d/qUHQ/2ko6q7XSDR56Mwb8qnJkSwDyw9E28DrHGQYUe
pevL+cuROIHYlfMUivbv99ad/yrFKQb5H1nBtELA1MZGVTh8cJukZ7Oc9jcYP2m25NsAlgXJUqQp
3/WL2KH3SLqxjVqYSk77WxcFXBL9/tbZKhS+LRxowl98cAC94jqG7/li3t3vM2kaYncJIhv+UmrG
nkIfL5qb5T8xSmsoOqoYhNrdqAfButN+dm6orAcJwjFkaEhFDRuT4FOlPyGXFUEfHVGeVt5SGzhj
g/PlyJHpugxbSTbdso7hQyVvd+EQICahJNF1KmnwGXlBgJieoP9UbDXcxwjQy6ZOfA+Y/eR14c1i
qwvLsBD5z6sOaBdKX5UDStNaMvXycD3ZKOvZiW6W9HNiaIWBYYTMC1A+YRB329Y30Z17v1njVrso
SMnR10oiwhekQ7Hg+GqIe9/WxyScQPbs6LqXsNdW9CcO7s3MfAfVk9j9TwTqzaGB2udCIxpig+uM
G5xbJcDx61S7Mlz7otkHPCKQDGhZi2FmfLBrHJ1Hoaw1Nbvi1baa5oqEqzhClvzvtnPCPHAlcE10
qqXFa38WLhRGL1zWUCb9H35VGrP7VR5jsBLu5Wm9lOpL5gXFcAYwFM3vmucel90M8+sKnxSUoS07
c+jg/+0qDs6eNLX+C5pgP/3Xg/olU3waf4UUmxYIoHPPSunjl/FZ/BqkvpkWrJ+NYV6uR3RpluQG
BLlxSIpzgeo+3eXwQfe/OBLVh5ysPKHPE2IKIc/M+VQty8mCXPq0kFdK7lLET8cqotA9z8eY0P0u
z4Ea88Tf0a4DiqElxLqiImWuDbGpPVvwZZhjLgOKUvTLk5iyN0ortGX/0YeIUynis2vCrQ5UYF0i
m8lSeOiSlqfEqRl3vRr4T+zxKvawCJvNkXxKYBMnq7JGNzXqYeRETBp/02ZNDS1gsLHtxgTHA/Wz
8pQxmlgLsSmGSM03DYsvP43M8pn1C+lAgYpiC8P60Emo+sk1SGenQAdW4PPfbf8v57CKSo6b8kJt
NRAIytfyi4+F8gMa8mU8CnXHLV1E/8X0SObKRgpr/xaCnTxUldb+vj4y9KAb5+6Dwvlh1Lseckc8
BueyMwKWVH/E/RuryuFhVvWyp3Ll9EegKcNv/9Fu9QnM0JVW3hJ0emelBy2mfnvyQ2mUhj0UbfsX
fbB14oA8YQNLhMiIqTuuSGMk4G274Ib9pjCe8hjDcbfj5Hmi1a3HEkD8XdzQIGdKvLnw3cBP5UfG
04IOKNRaz5gatL+EDsr3kEjptKqWTic+pTLz3Vo8Qfh1Xmw6l//O7HhuINrUDFMqknPRzuiFOgWm
F5APCapNll/fj02JA7XSBFr0S5IwsWuCzSfpkRtR2fbiJUWX+if/GCspoHyi31BNIX2cx4R9KCzm
P/pSq/MDtID36f4/DHQJsXtxC1P854W7XBH0kvgRMb3HF3abVAWx5x6LGG6/+P4mxVmJlDljIKHx
r4U+gBsKKJ9XILObMEiKY14dWThaRl+9t8umg1FR7rOnQex55GqfRIngRXorTNDlOCEpcevQ+iR4
GrlGtyHcrZak9GPR8yQpeilJm99Smt9KcMltAPw7Z/0XkWxaOVZHKhyip/7/L6SgSz1RfTeL8tty
IbcgH8NAXK0YQNcAGu5XECeLGY4llf9/f51zPDz7QTu/8HRTaLHvxo6iQ9jF2NJsqm7mxfhPzpxa
54M4ioFYlF0tYTUU6T/687DflTuUHnmiPH67FHerd4Eaq0E70hsG/AVBf2rwtM4VtIqcJJ8cbdNu
L5he78H6qjt3l2+7wcyugugTyb7m487DVvhwFznh+4VQNB8rL7fQw560NGkIHZ/DaMO5Apk3S2fy
Z4pKFbELNNSOvkywgdnOAqXg68RQcSmU93f2jCNfCOdtNUjQy0jblybhcVqgBoVgAdU3NaHkkHiU
Qs0o5i/g9VsuSnbYghDl08oEIPbdqWxwD3NrMBA7G8MSO9Daend3msOD2xqQGIih8QrVeDZ1lImc
5Lsa82z5ZgOUFR7Cbkt1niAk87jOSAav6Ld4gPMVuGPHm2RaNmncEachIEEFJ6rzgjFT85v+fsgO
o3FlDCKBGpJnnB7MBfsOGC02ORtfWKEGteaJxqw4QAkXBNWULZdd7dPvfTMXrpZmMn/4AyrD6wDj
fnUeZ0ZiEdEK3htme+aYPnY5vMV94gC0wRE9lto+eQdbetd1m6nH7mfNvLSlTZB4HiZswXlA5m6c
qFBEA35ww/8U/iovazLzC/wmN7IPOASkypM4qwls93IWTEv2DDnSPrDA58xpt8aNuckrfFnWiXWl
1eAeaH9ADsItB3xs7P7dJMxj1uTX8AhAlOBYIe1J5QW1LYvNi3Wbd34onvd6euO3Od8a+bVv/+t5
TEaa863wigByYYQ9fRwVGt9d8ZjGFlCp6g/izdtfwuqcQXbJqjDeRpk1bni2EM2PlXVd8x3XpXY7
PKFpkPUhSdetR5lFiihP/3evhTnbAJQ6z2Z81fE5L8gFsepx6DUQudLyNeerlj5fEGckx6BBJBZp
wsjXPOdcilzhXXg0cI7Wa778NvLArP7R1jo1mVpT2OR92F0HdTak95zPA0ZKr+vpJLLr6rZfiTUm
mSMyTXDQls9UdZCiSPTXgqvDFjOVA625oku940PR07M0scDP7XuJkpNaU6XeC/ESn9savlk2N63t
eZy3mbPhPtAboF4rsyzd5AO4pkvWTy3coOEOKvIX/lRcd3mxTT28NpDUPpRV1YzlC66JsDMbL/jB
+DKffc/FY/byKE1Y3nIpKT8hiAtQmX6TFnGyPdsT92YYFeI1QrcVUl5+58IhoGShJe8THYgNL9Eo
LYcwYj/NWz668qX4Wg15HTWNF6rcDzcyj64Np2+yhtF+XOKDQiXKCOjlF0KyXREL0rCibLpMtday
36b2RqL3CElV4dyjjs0kv6bMVVQruFUSTknXziggOkBAs19jqXIDlLwdhFF8ia0aUwQy0Z+/62tZ
WMm0HHIQN+EU0qanfWSkbLVUD5Ebk3i9yBDaR5jEmFnPsfoVKOQ0zm0OXWOQWeo28W0Jr+1uWEhN
4gJuuDVqg/049MVkniDJWBYpcRnSNmOkABn8aLsCekz5MzFDfEbaXRJImLBCoSZdZKNwdp3ZuAun
putJU7xE4B/NcYl1gCE5PhFKhMj2Ynearf8ZggoF2Q3UaIkHUDkDcUvCCZeMR0P4As27KmZowDgL
2iK57BPnLZZ9nESExoT4KP8u2S9PnqARK0MFtNGItKAbaTXe/op4I6emalskLlJa9GQVqpEcZVnp
5cfwv1dlbN5NHYmyjTiI3bjcESvwBtDWlgtkGZmRL3XxGsp5aEFi71BXsQgW6jzo9vS/EQcvcZYb
cmwJydcgKCdlLc+DDewIXe06Z57Vdlalf/VNUmcdda8z5t/L7Hj31q/nz6vJZf4TiFWcVZVBgY4t
5ys+h/MbWS45CPMaAemXw3WQTZPSqxdTQGI8L8/7W9v9WH/mD+PEsvaa5rM+zw8h8nAC7MJD7e/H
oOqXFGs01tfackRHcg1sMYMe3RKcq+98ezKkOcNe1W+hx3dwQvhfos+pO3v55p6P5M8zxKVvBiAm
OO4qvPBUeK3KcYyDCivJXL3eoInp8p5ohsTrPNBcWF73zrUcV6i/0dL2WFMW75peD704jBl2FiTj
0AzG01JE34T0oc7WUCoHBmc/xCJX9pPeuwxaUXe2CJCEsYgef/qTuQLdCDy5YsKYW7XniHWBmNku
IFFcCTXv8V4aQjVk44MiNim565YFihdTj+WvafIYrAwcfO3zhVOxdDXDlbN2a74Qn7lM2bJhks38
DizngP8u/Jq7qtLcfgoEVVbvqu+K4x7C5L9O7wxY+eP3bnpa4/EExH1hY8LrIz+p7NB7PNuw6Dph
CTlih/H/ibcp5E1nDg2i3Ks539mgIWOQPrf7VgRXgYDs4YX9fGn9Liy0ntg9kpTflJJlmXCvxJ1q
IhVOqVmo6qiC5D1zYGcanJkXLDawi0Hkp9Jwu4sk+NU/e0Y+jPDlAVAil3D53ZmRsRLTn7DKYnFE
dPE5Jgs3r0wS2/++kAf7wKFrJIC9xNx0xYuhb946yBNmuaFy3lZw9s+vqKQhS2dO5XZuuToafsl5
802vWh6euH3MB49kBycptD6EHCWuWkLL0PI4REt+iIl1Tcq1u1lLRHXoc5UgTbFOs7zBldswFIKm
VLTxVp3x7M3LIj0qYRUtZNBwZKQuZMYzggHtPWA4RabeLmyPWrXTxSy1UDGL9b8b0ZTqKRJB17pq
4MWarvt3uvbCeXuk1dPCy6N8Cbu2VQYyyU+Q9dKJTaRWnLO+/AirdgESd4l9hjmNEh8RArsKJExS
i4dkZ8Yq40talTFHNQwsLH0B8pxfrF6OqFyYpvNV6NQDEgKbjvYyO7FtTD9Bk+b+yJp6/+ugnxxO
evXONu4+Xyg5/Qe70jntzexuXnrqFyolCynv4Xvu5u9PYoym60Yoz46FReB1Pw3g4qRrSZvYgRw1
sVB+NWiJpoGBDvceGZxGZmm9MQFemLiNn3gP12CWSV369WDc3V2sg4CiDz4rs2ZJ7mjX9CDQXHJC
/9PLzX8/FJlNFUyPbRPs3KN5676AI8W1iE3vSiSsqCLkbTbVWwtedhqC7NCZeao2JhB0+X90mQm+
1/i4UN5QV53fqUHOs2FcMhiMzaWi1Z5FoiN1CAgvqA/8BuPytpK3fGlh5iVrmzmMlOsUleu7p7OO
IfrCAggF+TrmGpe1YqQou91pv+m9DqB/n8bGJo87KCMuw7u4aDXbyoC8Jqn3POVqhgHJPTo9cxh5
qak0pO2ZsGNBjrzxF1nCJ6/10SMfCWLn6kU7kUmr8JQ3fr6PY9iGhwJ+bDwWYqWiMfeRIkq6cqsv
FVW0MsCmOV2syE4tQlFbT2ox+dN0AOOEcRb4gIFa53zEYmSOOHvDvnQxbBN4miX7TLiGA89/vnqH
ZzrtrEE+KVXTH3LQEiy7Z52LAuqUcXYQVVr28bUsqyKXOwkqeGHxmoGCSEi/Iv+RvMQiGQXToGkm
NnEtfOt5fCPUTESaXEeRWC0BF1sg6oqwt2p2M4T7BiWolc4pbIxVULhSAxh+Qyjwb1yFo1YrEKYk
EYFgyLSjcTJj3vORzqv8d+Hma4ZtIdUrp3TBf4eNHtANfxZ9uQ7TBoYYeC5mXdf50JZQq/8flCF6
lUGIdwTigty6y2R33BknuHX14J1UclJarSS2YoqBDTO6QvXF4Tax6OO/Xz3PUBkTTGtJszHTsZcV
pq6QKZwiZF5cX9c2nFiS5yO11fMDPKTVjg+RO3bcNb/teob6AIkMMo9x+llsvTVXBZvr6iYxnpbu
Yk2x90LpmSG7gh6EOFJc/53g/Wm5AEw8HKXa6KzpvbEDpPkE+9RVnAHrKIYMXrNe+gpbTeY7ZolM
BQLFKOichH1gJqYjBJx8LbmFk4NDzJCtCFHrYRXtwkXqlBQVQMpU7i2HuFb5tbR7HTfOq0PCAukD
PhaUZNfU0esqDRURJGFqTg30UMvnLM/71HOlLifFR2dbmnKakLgJdnL9WhRezKTCknRWPgNEp+JV
cqnR+oj52w86KgRKmJv9Y9v73qvH778y3CjAMljWOVBWZC6LumJH+L1uWYZvCo/V8y4KMR8XDlq+
wBX4EyYOeRkqYeMGVHkatvEUXTXv6VmGR3Dd4Se3Fawh45wQ4bfxxR1RsX3+23T3mefERl95qDJl
vNCK156MYVcjvgmKhnlXYZENGghtn7GjXRok5fGfqEP4pQO6EhIksDD6koVKNA96T8DYMPhbd44k
4xw4ouMAsWhSOoYWwsclxcfV/ynfxD5PoBSaCfZifbUJCaLQJ4kgY4Ejq/znMh7zHoO9rNGEkaFg
u2fKn9lYsdtoDED0g5ahUb62mjoo73/IG8tclQ/JTbiHGSkW0NU5FgttHlvj1k5Nhd7YxIw0cSJW
I3DDX6Qq/fbNUG4FBQwSyi0n/psHdTf05uwiPOG2NLvSnveSaU3HW/oa7mEA+k5LxC1JMAK2YW6U
6Tw09B3IU4yXFS5VZAMt7rz+Dm8912s+7W/jnjIffiTWepbGY3forWhWoObOryU6eXPzrMCRjVo9
pRkUa7yx4syapD699LkontkfpVnf1FWacsLK/3OXi4xnMmz/hdAVatG0/1HH1GtkRziBRS9iXYnl
ILuC9FG9tdz9Nv27/1/yj+B0gRf1UA0zaSVhAY/axVOlbAI91zsEvCQdsj+PV2uy+CQePlqJSsDs
mqCzk0DpDP5Qhi6IecC7zXwaajZwGXLtQrF1Zp/fOCqXWXe7/HnGQL2JrDcVjPF3vmLi23QY/RAl
fQpC6rC+UWwQvMRA2pBv5RsQ8jCstgx7MzP3ApWKdkHVzVENL+itraPUB1KCWbzBMx75j9tWO8AI
k2MfQKN+H9Rr4rPyC8p1haQ7YVa+X//3DyGgDYQrqpsBq7u9VP0SfRKBn5SmMbAWk6fEGwGnTfbn
wIFjGC7hUEE+g22vpWBd8RwYV5K9JN8luHuwC+gn/oXfIXhjpj+RvO1tk1yFhkVW1GFv6WKm2fzA
OmC5CEvAKVHd08EBbokTEakqL2goexILaZj5lxNsKhPIgQDZ2frfGYf5G0vsIpaWdHO5cYkjcDzx
QjYIaMZnS/EmqhTBdNOLygWshyS6XEDkvGyqS0APQSjBT2VZhQR8ZZhAl6Y0HLW6yQNmCygdwoR4
UfOkQznAOZnMPLOkKVSXYG2AHBK1L7Pqd/9UotDfR4DgftC197CvroOR6OFL5lchirxj3aDLcnf3
TlATlcBV4WZfQwMV/fd9cVmxXKnx5EgNpvK/QQ10BXnVaxDRzKqdaZPuc18SVNtxdMHiNRtxHbGh
s0Me0/PKYD74lBxphAm2hysytIPO87MFU8zG21G334pD9vNHJbtZA7Hr1YdNSIZU7jReQ6kcriQ7
x9Q2mkG7E/cFg4pR5VK4xfKyOgYe/IeE2NwAVpxlG9XLX7RBywsX9wdH3kwwQUq8EgRv3ju3zk9v
ThMTHGqOQB7+hDMGCgkWp/BGwrLu9H8G9t8YnKo9Ak0Urk07C+rm+NzQIm+ZzJRADHwGR1Rt49F0
XNCBFTTTX2+ITBn0DFU3YGFMbuEY2AhO7kzC6EI1G4SCbbeR4ywcTcNOBcljUjz2JSpdyDYrLEDA
lRasb0DAgnJ7FYwjfcWVSznNDqVkK5XZBzYIx6WQr1ckNMlyh1kmiEwotGAFM6vmWVYjae6FmqDo
zacdeLywcGJZ4S7sneRESHnleCHsRYmQdj1RWV3l3Ddu2sPuH4gSZzi/A7tbwHVziieSRmUSYgO/
+TYAskViJBB8cn6r+6JFV6+uQVZ39XfpVavPx8Q4FsNhTVKJAfHYNX1e8Hzx7ZZHLXsZ/2Ch1SKm
PJkZP6CjK4+FEUzH2vhE8cP1h+rTflWFNDEdYDiseaq0OU8KupAdR5dyi4K3vqIaPc33aPizHQ+l
OGL+4d2pYFW4wAGXM7YTES61O/cxkzpHZLRs7R8pQMaS0mhKmrEQbAvX0Rl3yRPD06IlNq/sMaPZ
MYNP0zcnGAY0HyTSFjChjIcADmt6EY4NHz2A1HbNsbmSoUCmwjHp2/NgrOSu0G5KwFdmfv3Utl7K
yQssx9pVaKmFApLe9wZJqFvhF7Y3ENf+7Qh6Cy0cIpM0CS6yVRUHN9pqoetYe0fixZLIhQ3q8Imr
vKn3XLCALqTdut2TYq+jg6hKDW+RknQtua2qboWU5JdFJe0qzlFtKYjUO2s3rLsaUlKhTtKtN+Px
2e6SKK9thVSu9fFVdnuGmOM1ZG6ttqb6f4nm4mnY66/ar7wTimS/JGyYCPWbQFyVmDW3jPviJqti
BCTb+Fl19Y25VWQs2ocidWKgVDsWE7g7jWX/7XmojGSHX8ekmCZYnMwmNuk2v2BV6OwtP/zasQMU
Imv7uRRRkPaFB7UKyhozgvrzFBMgCH/3ErdJ8hYCDC+QtXMwe+0q583HwInegCGpY+Re3I1ypqtT
8nswFItIp1Ay7Y2/jfgNhOQa1XFdedSUGM1zDilZhPgOLH6k24vnL+Ixqc5uYJaGYJztwnq5NX5X
B4bACHoG14Hk3UO/1JqsMXZPrMcCVADHE+zU2D6Zf2Kjj2FQRSNTgev5RHgn2s45FeI5I0Sw3HKV
sZL0vW7VK1s1PEMtWJEuSeWUZILcgXVN35crIXZHTVaqiSXy6Tr4XEhd/mk9/tXwTxK/b6Om3Nx/
ke6TNTMXSaWt5Jtwx5+G7ELrTB4203ztHFpDZeBMGRMZSHgpMD/MGV4GFV1uj6SPSzQPmaB5dU8O
PS0WJ+kuD8Dlj8QsVoiUTtAw1KTIxjXLdubX9wG0iHb0J5bTpM6aClGKOGWaQrd/efBCipHxp0e4
jxFXDaRs8ExszVIDjWUCDEc0CsWv9shxJLxhaGIK0mV5HXmBlv09B+u9dfg9kUrisb+ZaFb7gTUa
D6wsCWsw/QOLuWLMtmcRdU72GP82dg2VdKtcPtaCGtckgYmwuvbW1Lq8jkYxP/MS2syPiSjzkLVP
NJGd1uakyJ/AM//A0RtgJWa5Emu6t097+++BIclUqSIWart7vR45UkhKrFDMiLnn/7AvJtwVNm0V
RQbD6ewy8jErN0EOr03kFhgucq3xBKdCm2+kkwkxGF8LTJ9ZWiGpDIFOHKc6gn4RdR2VP3IeP8BK
VqpPHWJdWxTdMW5RwlPUvZyS4VbtBgXe84CH0eZyhNUn/z+QjnGwV9XhqhWRrNRTexbww5cmKmy4
ku67Ke0dKvi0vNZwwb27UXBa7zjHOGv+nL8GFfUD9wdzPRRvd3LP1XMnnIuY7BvlbrzCw+STkvmV
+NXeTQJiCBYqv3UsMbN7qN5c+Vy1fLqALIY3ksNgnaIY1DW+PEcYrrjGIE3VLSSZ+3db+IGw8UOK
89GWPiMZ78wua4J/3xL+IasYFvt5CIoUCO0YW7tHIFRij+3R7iTH+qUC468b6w/rSeVSdrqWvNa9
EIjw+N0jEBx6j99purdSllytroSOlafVGwJ4G2W5bSFIRe2YkRNtVmZA7ERCDay+nKuzsOSFwlva
xMTlea5uUzu+KCDwDk/g0y7SCHvsXtWnJU9DiNBTJpuP+9Y7vd2gcKHWUX4w/TPnX5NyZqNSHxwp
qFSp8iN0aCOPYfSO/Gv6w4FUv9fBDPC6ab1qcvBtKuwVAaU0xacr0vJBaB1qWyW2zXBzxoaTjxGs
e9Q6AoeVZSqjWwUNcFfIMI1VMK6P0j9wqIToViTGbGb3Uwm2y75xLyYnSaU+xPGePgpueMD8B1W3
fVxGsZFTFFyVsyxKAiLt3A6+L2OeqIxfOVcbCAK0hiP+lWW4rAKTIwf/V7004iaj1D6SQ/GFJqWa
y5LoCfyHgB+0NxsZ1Pvw1N/d5iMVRXK3uJ3DyDNN36lH0KDAMVlXpWhZ+sW12ykS1YK8uLdF2khj
xGOro44qOKMdM4TerRM5mtpjka7o9enDZpe7wMt5b9YB5EOdKByoHNT4U4qeXQ7ZpB4mUnGLQHTv
r8seJgLmUfScJWwj4lEM3Q4VHgk/jeHrNz42u/wusDaYlUA3/fl5dxJhgiaiZGJR1pjgVS0Z3iS/
B5e8gnjpakpWECcNijJgzHgoKHd1iktYNLUV4jMuive+Fe07AiLZ0mh+CJQdIJHbHJo5ecX7deVm
0RCBOsv/8YeHdR4+/vxyODbEfptqhHSmD6aNUyRs0Bo7xm4gfo/YqhvzbJEPlFElDwP9MjfBH0EW
8xpGa8g8va19Jfjrpk6VVFhDnL9h6rqgH56q3QuLcr0cmVwpmK7leoFK1lW3JvjlQIkgEJvOfsQ/
qsCo6o5aDDXG6r9yjcXzSJmOcqjXY5WztyKV9A2zlpsYLuA0ns44iZHnHgn3GnR2+zi7uxgwzETF
Ticuzzub0dWX6SivrF1SnAhLaZLsN2H2g+zBzXQdeSS/JY3n0XfvsN2tqGdqe4LEkmhBdPM3PKfZ
Cy3aDIfVQLAINcq5g6zMTNfT16zaSZTetFOkTGktvoo+LnNzBML3WE7GX1sOWdkr+OmcrWGMOX2B
l2B8J4d8uATQYYlUnhZHQRztJOA+j7dvD0pTTb1WcWjW+2fYICB/46Gj4rZgG2MsF/0rreswMqP2
+XAseBJkm1yzH+1XYcpKg1mU+HeN7sTHBMM9+0pJXQqVW1JjY33IDIXRDhbiRRaVhucTeN929mB/
NaHW3jbCgKdW21hHcnjqUcelqM7xg5OmG+BYccRci+P2EXV5w4TXVvB6VNieNpOOWTJKML8kvULF
yGecBdF1MtuJoI1Zw0RgJUI2FGA5bs9+5D3fXA37e3enGEo8xq+Y0ycEYy8j8Uc10QePPT6cBlay
IU3cD2x0U/DAXU1jORHTr0RLYQVAg+JVmnDp96tuqpPG9y5NNWWn3yEq/2/B+B3iad5eR8eKL15I
oI26x678N++bI4b+8k5gO9ES+85UMiFJnRiNiXSb4bJGm0mTYnlWbSj0NPs5Eh+7Z3JC6h491p/d
AHrJaIKHKug/Zh8HroIkp6gJl8ze4gTkudySrFlJVZTPZt0cwN6E8tjvlf4+wHbTAlGZU1scbXQE
hcqfW34URoffLBVhxv8hPjtZNiwvx6CNCqBj70OBpO35EJbbdf2XXfUbDYr6VLf8I3cTL7AFnacX
mYQtgbtF2rp0Y7PMVms8i9TirJ0q4ZREFP0oXgiv5Jztz5zaxeN3Xk0UPL9KKZHyhhOW0nDURB8/
nb5F3JB5D65NlseDTaVdMp0dyPha3R20+rj5MJUAe9lGYboHmG7IG7FD8+3KbNj299hPgiRBTTks
eGPQudeLbL0SVZwos6kGZZ6Vlq+YyJOHVed76iUsJYuQtQr7kc/bSN3RdRh8xduUT4SPbQpNI2vY
kfpJwPW5Nq0XQFFWz0YKyrXoQaMES+Yf0/ncIsE5yKTyLznYYZcvWXB+oGdcgXoB1aXjrO3GRN2Q
kC1ZwpHR1Xl2fwZen9Et62zfxlj/ZjF/5UYkcTmr29ysZau7zKZp3TWHxGq1TUEqeKFP3CKZXvvl
/4Nlj2miiB8pTZoH3GNfx9KcQqk3Del+ZUWpED8rvPmcHueFvDSA4lq5+d+NtdiYBs9njUbF89QP
VNOVudB308/BLxF74l8PFI8uRlYT7A5RFL8Hc+QSrzDUNJgriVVwrLJOyxsAbT7Lwc8BGOkGBuvO
sFUB4SXx6Avyhg23yWN/h5ZdWsTNNir7E/mgBP6ArLrzeSYxRk3hwRTZCVSHjfx/V5kPrFQfG8kU
PdRaoyiLOpKi2KqViDRKwtd1m5GLXsdFTLC45SsMruYbBHlzSi+FHdpYJ8+on6YuP0t1gZAOHWZC
/qI+tUlaWsZlgO87hc2kEHIdAnsjeMp56pz/niElg9HwbrX+xuZbS/uFnA66DxM1wLCZNopSrZVO
gLdgt7YSjR2yVgxwS34AMgfW5JnnBb4o944HFQiqF/RgGJa8CYlUA5Ja0b2xSKcnccg/Uc6mXk+N
yN1v7Y5TYGdIZLQE7wW1oeQdMKNiEWWBEd8W2N1UTV0W31iLw9DlxUIUG5whXp07bvu8cVuDcnfP
UNpm0Tp4OABi+GvFN24fGLO3cD3mWLMytAla6ubAQevjKaBpZlsHgzynZknbYv61xPTZIJE4Ka2o
XcUOCMzR/qg6vn8tX+Nf+O9UMe4e3eWYO93Ktt8vNBp+z72xMzmf90SRZQsZTXv42zK7UTuMYkmM
09i3ABXjrHF84+9vKcTIAu3N6VK92nkaB0CK/yBkwpDC65xBT5Sh92Wmcvs2rTV1FcDYa7nwD21E
vZOEmnMoTv5JD9hPmbJfcl5DCcplYB2BbjUzRUvoih2aznFOKkjzNUyhWfPGL+OKxZOlAnTQp7xc
CwN6eZUJeS34AbFz3Zxb1D8On9utS2m/FMyms4vSXygIEnldM+EBsxvWDaibmNQ4cmoe1q/jZ0ag
7MhFmvu7gtKCC/0wkQXLkpnQ86Ys6gxxugR/JkcyUf7WqBRlNXRsRkHWmon/bqIzanfVzv6NcPRO
2gCpiayW7VtfiDTx62LFpHpYLAWaohU+cRGgl3sIX9CY9Y/i4BwHOji8HCnbCgZrHQrmKwB3H411
HzU/hsxuhs15v4l1EHtfScIz+5BYQWPCPHN2d6KPVjZkRA4ZhNQzC1WqvqLQCPJWmn2r/gApHGhb
2HabPimbInCP+dIrh4d0074MAbj5fzWfDuqEnVm4/XSqi4R5hPWGzE5oSVBl30OXhDmbZpZWLaw8
FJkOR/mSnProInv5/ebK4LPkdyLuVnro+t6ZHoi/A66qTG8ICn7MfsvuS2EdKNkjdLOWVIRnKwyh
fnf4uYgN0wZ+wgp2QqVn/XMC0o2EgPH7r/r59SclGT2KBYkOc9ya+dD6otuwNJBAMvsTfFxlTVH2
O/56VcpAyiwIYzPeQbK9N0CwVl0j3UCsR9O4viTC9joiVEF5DO+LYvt7jOz90vIdMZoaQLfqdS6O
8aW0s793cSsbFBlfZJ7xsBZezYtJklzEVUUfjIsRuylAA8aXgcJ1KaZjKVpAAdQB7pusDJq5XLnW
x8ncxEIMSDoxtaxQ7nwld7pcC0oKKurBYNIXPEQ+JRz4403TE6/VxPiw1q36pn3FdZ5pgBBPLq0V
OcbqF0a8+y39ShVYLiT8B4jV1v1LjfHOJWDKeb1vlZXlAD6arpsXyPwGX77iQHF6NAZrvFJKSW1g
AnVViwcVYvgznIoJaFLUGLWpe9CnvWKmkLG0ZbT4MH5gGk/Gh5rSBSm3xPqOSPwj/XCiNB0bgqDW
dAEQ0GJhM5+Vu+RuF2zWvLIlWIG9xYpdQEJTswqHGucZ2tvhFIuLBPTWThGYB4Xa977OxTmCaVVK
X2xVAtg71ilD9CQ+Ja8O4rzB8jwbm7yMdHJChvjEGb23jOJqOSZv6wYLzh9H+6RKjgOKzaYwvQ6w
TkUs9+3IboYqm1Y7evmfiGly7gyFXLbb4TBGXzWJ8Zd04dSFzBLsnQ23yapxH4CdXPme8PC1a+p4
Ik81Z56ynqxgus59HRI4xJ/383ieD1YUsIXz9aYZub8T2skDuxagNYm4t+VNAaD+EMriWxBxe0dy
ZjHMJqhs4O2YkYFVwouJFDzVSP3FNBNh5IEzEB/lA/jKtNIxdHOMlFZrN6Tj83f/k7YagUX7OZIn
QZrWrUTnjq2CFVJZ9/JpDx3ntab1zW/fMoR7iwhdNToDsl1kg3fTbZ1Lbix//Yyvj+BK1KDZOFt0
EBgHvkw4e+Py7CSvRUhoix5hnpQykxHhtvrb8x1u87dYIAP+xw9UNki8+Z8oakFslZIBPyxLFzeD
VsAf9cCS5X/uoX7l/ri6MG3oDTFYGUbj1VbiFWzR4T7Z2lmDJXI0iXn0Nr5chvklHankHadiq16f
7g+vmftKEWw41mDuLFucnrH7xubwQ1+nW9ygvv4Pov1iYDj67+7B6tDWQ082M1Vful8LnfzD/M7X
kDKvX9xeCFT+dhHLYFweeQeBLYi4HjVb4jv4YCWLLfB3Oyj52LezY1q3TX8WUjkU68SYT24vcj/f
pjxjhxhBqhQRv2jz3PsYfCR7KsDWhY8YRS0usK3vi/erTlVSCME7RjCQ/wCf13cvqjSncvhQCj6N
+nSndJ6wPxloBUitozNr3uzub1Cs6KVArm3mJnp1REpANDw/obUNlwLjtB+TpzUwd1QeDBwMDqEN
rZg36ho5I1ImEWzFFyY6UcuwvE0FsgmEW+M0QFw9GN4HfipjghX+Mg999WVKzO4Wo91N7MMSsjq7
3ytWBo5ShaGtmatmZrQbuwQd4trTMFhCHFVe03vFNDDh778oIpG/dHKy3yWrOFGt5Tkdr3ceetOl
TvqdWZWCafzP/6Tp+M4SeLp0b6s9th5qb7ujCKuv3aAw1U8ak5H83jQ/XRZoQuD4ZoaIvB/62M8t
DFoKHF4AAKQ4DrWpFy5J65SDhxEeFwPRZA/GKOfNfDfse+4FGj2QZR4F1vrjfXBi1lU0eE1Hc6Sf
gXlR8RIGw+JAj2jv0Gc9zyy4OqKnT6TWCGGVXz1hWYAeQKxdS0uhfc1NEyFF/zxcMMBRvRAzOXOw
7b2MugdhYTaWPVomJ2+7veAZRxyATqK0a9nK8nkB9iDWboF30ao/007Kwd1Dy/IbkMyxuxyDH/AX
FPZCaxemybbyOgQMops2mcwsrx6pLb4+Mpn9nMkZWvOnNeDBJiFn+GO4E/NKVPaAZOW68dcM0V/O
5Eff5BgUJr2FfLDAPgk0dAcDoHq2HHV4oktsWZCGMC5tFVB6XKTAeN2f1CMrnNY+8Rk8KMIDmhjw
R4CqA0nk2AMqlROPouv+hXniM/y7z4LI3c47YNdeAc+nBVb4w1O3IayuNgvUPTTxmWkP4AtvhuUs
HE6SeYUDAJDidhGEIpSkoen+u8YR/exCuIg9ZCznos9V4n0qndAUKvs11WyYM6p6G5CLrkvcKVJ8
yqFsegxdM/7wS3NZkXJwCkg7j3RktURAuKTHFojE0cJHJDYDspiRtQy1odbQooTGHRMCNYoG+EA8
7PlbXis+kEPRlpJo0e08DVToB1szBs+v5jIjfU5MUhvzqltK6PunWPf17tGIGEeGTQqAuKlzIyT7
3Bc/hY7hZlsvK9EiQHnkQvjKuDLLxEetb2mpfsXbItxrkadX93kwjS3cMnootLkz1TyHaxJHn4yq
5nxdCsPBdE+RLcPsEz5nucVGtnZj3N8/jG65ZPwIaihiCmxasOZ3r/4AVmdWm1ISNN24iyVrxgZY
6GG5jeU14PrRKeTEWBXdWs++RIwPWbVcGosSuJD+XpYly/oPk+W/wAc35Cw6BUeeYLimffZV3EK5
vaUK02eHx4VTsIseRVG1pebHvvRnHOb0KMFRiWd36doN5ogwPMQSrilDdMQ2DudZUrsvDY+xKZOh
tiFLV1AQaaynlqMkLWIlSjfgvrqO0U7mIiI825ETRhJzoRkVzSGQq+bp/omsy6Y+naVPNwAWjMTL
GwyCFPmXGlv/Uhy80SsQsiAYfhWAUviHHVoLR6i7XXPFQaH16r1AU4CFdxf1xSTNpJSZ8285yBBX
/OmWvpPmGR92po/+HjwKXSynTv2STW9Uok2ZahN0GJQqlVC6nE0WguHOWqSEHu/M3B5AUZxstM0j
X7QSt8RxtidQXAp7GYuXFREnvhT2Q88+vDQ1Mgo1JinZvIRmfcEfdZlVlz04cOkbnVFm+j0Xrie1
OAymG4wZliKS1++QlQPZjLot2O98N2ZiablXQ6/Rhj7/b8M3EJ7VouyisDF5I5vcf8qBe8sILPnH
TA1EnGjH2aAL+6atI06PQQAebN8KWQRQc8NnFHNk6zjQv2Xlg1R3f2/xa8QJysPQwqrzlK8SLJjV
bwQ6Wk3QHrstXXWB5Gu3SIb7AP84KruNMpMfiOqsy2eEKCQrgJHwNplEfBPeNDed+XK53NxKAIBG
j4Ks0Z9mGRIlC3goJ7LH8q9P6boCL5bEVmJcuoIMHK1SLzABJgTXHDFKZZd75ClFESPRH4YMCrpm
0vQilHyFidP94XwKEhQELsaH/uTQlAXy+HbS6YOEDa2HVv6NkFAGMxABb09Sg2CyussSCRIglXCh
6rNoW3MWeTrnlG4GvwLKJzbsWK5jhVb5m71xldcZCT48Myb+Rdr4E+uY2jfWOoevxHVI1N7AdL/U
nsbftTLIR25uTxJVGeVlrqRq+pulbRHrOBCwyq7w+34+FDa9sOYPPI0Phf0Nsx8wraeiQxJcnExV
Z7TYJjhM4kYGJTQlboMhJmcS+Cn3yZ5t19Y2CftTc4CvjWo77X1X35eAARmFJGWozPXbNarDR5ao
o9kS2yj/bdrqhupdLxeNjhNrFNBiMcwfwgX+I3ush02gqxt/3AK1I25jyCxp/AoDDPcp3UmrPgf+
uoJBYX0HR8dHACaqlho2GNmreFfllyeuchjt3mGVJjDli0ttsESVAYou4BtcfU0WPNBEbDBXa662
10tedcZ9oa7jqAlsDm7n8ZTQzSFSWtFxBSVmahTnB5ZzxugQ1xsSYnJfRxnGFr1bnW1pwN5DO+to
iflIpuNOX3fSRtytBDAdnYjN6Iua/zIwoHd7yXefUh0aKgLuKFUg5EAPJEl6WmrG+StVQ4c2OxZp
7YJRzmQ3y8cxavL8NQTEiMaJHgseRskXO7D49mXHHatrs+RhdnGdu0OjNkmNNV8rY5YbewzJs883
gdNdJVxKb/dg/2TkT+4Sjo9aQ+blUTSc1luGKakiaDz1/DDQ4HdnNvJXu848EE0HoDFBsrVCNLLT
JZLyHWfCfehBsxdQ0Z2gE1kjMvBf9W1P7i4OuyjCQBvke3jD5Rwf2FYE4qj9A2/ZRJz99pTbmUuA
zQsr2Ib7rtwO0SL4xReNZ5lKaISSPx33rGrGL3LCV/5z87fJewRhOsfrjPOfcP9fLJs/pIg1i7GG
Q6oHJ5xsJHb16G91p/RJuqbqMDZ3CRxgMCwov8xdtrBwA1wvPDoX/JVcafB4WLKhPtvq7MkgNTZo
Vg5FtbXMEhRTqamSpMwf7G+Dd7nZ7f6gjrjuRGK0PK90fqkyNC972y1rgHz0vGGIATy5z8//07zN
qR9sXsq9C8C5oV8xeNJzQCHwsVBBWWDlSTkOcMAHeCc4tJfXhBsw3SN7tZRCMFK2TpiLx1FuLuPY
YlZ9k5q7JgEqEt0m8AVNkIA3NIjAyUgcexYSxImJHEg/OlvWhEO7g0JcQC+5UvGJYBYrgpwb7W9u
9j2g/oA6NUfVujQS3xnErtAzMME/sk+WDDl3I5jgsmVRLdPuuTVMxrquWLhi0nEyLp+2XHXSUesc
acZEIe+D6aM0ebMwF0AiuvSi54/eW2GIsQL6uMaBrjsgm9/lN4fhFQnQHP8wj4zi4onpZrItpnIp
he26jnyeNG9G5T/HnQxcSzdl2wRd5MR9r5aRYFfnxZDHEBtl967Aq9feJQe/x3y9ZKpRdpw5vqfs
y+J/raf+uuTPs6V5FAmYRv3/Kw8SKU4coWlvcetpe8VgigajVp7aVdMhAs25xXkNvoH8hZyXrsXX
qVDgy3oev2KGGcsNxVy9nHjSCNP6d7GgNY0UI6ZNAPNzn9/LTIzfqY9dVJj6mQyzzPB3ItRhaoDJ
4Jc3ePxoDk/YRnh9atV5D7huAds8qLFbNj20blsP2aGRhhh1eWlzaG+uCd0NkcV2YykSqyFdz+6A
97Z2dSv9Cy/Z15YhYJ4JTuqrQ+LaMFhsfh5GCRccZawXQcFedKw3y7mSUtLVrniGQq8vDxsJjiCE
Y18j16+NpIK3btIdWdwaCO9zKiiyPOPyyR7w6eDXfWzpQx9iHbdd8F5J1SoPXoS0p3jbg4jPGWNq
OWCZJeJEwIQdubMx6y95KXnQ9i/XsKPhRaPZVIBNSscBHmEfWdR3PEd8o23WgRC3jnDyDzpljiZ4
0ePc7o9CoHpFQnk+zgEXzVy2xqrX9WMVuH5ut28KbVvTHNWAT0B0qeohndp2SU80EdRt50xW4vb3
rfZ8MI6Wa9kK3e6m+F7HY6AlK1DWFZuXd5BRm/KCMTOWq2KjjbrCK8BtgoqTBdMDeVY2mDG0Jv7B
x1wiPgLJ2aS8REwN8lSz1nMhxaejw2Z9i17ln2bjAHq3y0ilR/qLYNwoJatB8UIQBErdHnwi17t8
nYnzMoAHXAgPipFy+QzPf7/KvpPlSZaH2kCwbBPHqjeGvUN1AwrIP1k3OR9k0CM7mMzsh/2yGs+A
kfQ6WsoM/L4d7a/OfOrTnEsmBcBo7cnXuFBYkovvKliWfNKdoGriNxyIo/LBxT32vnmYjBkboeCF
vKMxi2ZqvekbP8P7y1Nel7541eTY/f75Zs94uGDf62V3MIxZQQINDwuqXe19qc/gWUVJVruWuKz7
aE/QXpNpCrSC/3D0p+/G7KXu3sqxmhRfP+0my4hQdKOCTxu2A/AILpmZpCUwZOf6Yn3Z+nFGX5eE
THc8JMwWui10A5KN5GleCA1NIsktKjmfH8/bOf5CMVklizKbTGWHcPlI/b1M3tTgvCBaw+L6BvAi
8P7SkFE5kNG+PFfsmdQnBujMgyoq0+U05Q1QrUzXXrKUtUGDJTrg5UlNbEiC3OimpxonfpPzHL5r
4N1lVNX+OAMByC69fNquDSNCtdqOJM7+NM4K1ZdAMnAqa9Fm6Ow6l/R+biZlwkN7KKZzNvitas7g
fqceAHXj5MezF1skvjzUwWaLYyG4cEAlI6035p6CYq1I2ioJ0djuIRzf01ZbpuT3IJ5nuQNqpMSB
lwmB4Bv1GTDzGVz1+7+JBqpQffGHqjGAAQ20Wi4/DsFtIUhRyPM0RftqJb0UW86doR2Uj9Jd+Yv/
bgqKgI+J/QqIZPAkGmt1Lz1pnPq7EHvjpOLCebsxQ/Efe8B7rzqpqdOsRGNHxGjDuYI5NJPBu+kd
KBMJ7pGHS764MIMvXSsIuKV2AbKO3ALNU4HdBE4p8DK9HLuAq1FIQU2KeHyTP7LVFQKkFWjtB3wl
6Q/zewENgS0UI0lS+FaUqgmfR/NpddiXzHpVhd1qEcURk9A35X0HC6XoroQQmWwlG/oXk7BA1Bu2
32JG7sRQpyCBjn5dzip6EyykvwCfyzHepfurWe45b2LmynUDCuY60tAEOrzQEKCnVmLIorwSsSEo
r/HO2EgpVwFelclZOGZ+lsoo1VBSRn/C87/mbnzwHyHDukUOmDv/9m0wQgs3TMMH6GVNoejXOi19
LZz2d4LKd9tP+jJfy50qVrpBjQbXVUZoJyzpK5qsGhdE2pJRtrqE9160bYQ5njggRsF3CzDeXxQu
hLnxaUMCBppOI/SgEIOR0Ix4gSjrs8R2EDqvDaodMPnA6QQSzaLbuN7Vpc3ZtOiKVRknGPwxI83Z
YgHC5quqjPuGTkZne6pWqCKI6qI8AlW3QMIrBM54grIgP6BT/pjyJPR7Lzh2CNoQeuBl9KPFtVL6
axCaiFNpFhrRVezqoYey/4p6CTsrXWQZuDp6GDsrbK6BNVc5NUqmnJvn5niDluED8QtagMaBajx7
W/edgM5KtochDXMDxzTo8oKLFWsqFNgW0+Rm/hOLYmBLkDkbAjAqqaTCGVWpdytxlbFYL/6t6u7G
0EheAdIWiCPQYHkb61GCKzSVIKhA3fSWT6QrqwflCbzCbICDYjQjBypETHZ3obLRStglSHENMtsD
4fylVKcnadm4qNkfp2y4bjlYDrmWbmROGEHEv1UsnYOIMLryLZzbZz8/Qdk3YLjF8IziRjQLE3rw
zly4yMUFRIwYOTadnYKCJJOD2RbihTAmW7Dota5vYPSOyIBrlb7GnEXfu5zzgDkrTnmUu0httyJE
AwV76U5Xr1/+FVGkYiJLBNagYdjVU81B9Zh56pdrCsCYbKhBODJP1hTXVRvRCKkNTyxMR+QY9unT
aTcjsa0SclIGw5LCXDS2uv4NEDNaFl3GJJvB2TMehtBvuYGz0wAqPYUuSmsnCVzyghwLXDSsAqJ5
2yvquQul7WhBmyy04VKKDc1AKHt4KwHePqmk8kCw4EGa9mj3uPN16d6WpC2Mst71+6ZwGiPJw4c+
eds0Z8TpRHIjc0t+xXveOP52Wch237PQ6qEGrVzUyE/2LqAPmBvkGhZyWTJLNHUEzenh75zO1plO
v4fvDCdBubQPa1pzQVAlN/chNA+PMLtNTxV9l/GzZ814C9UxWRkHgGXzqRY5gwl8+0shqP0KUV+r
9wjxPb/kXMgM0HNtJThvc3/9lirBbR0DD+BQ0Il5L0wQBmNxnaR5F7IC+GpT0+AIymBKTEHxmO3b
goqXyDOW03wtbTHmEC3HYSpUN8KBAPq+fU0FoSr6ANnBGcJI2VwulRr+51JF/ZM4eQuWXH3qfTiS
GPNNMMPdcAO5HxeUkrRf2APzUNFkf0dDYsjrrf6RoPclvasuTYGpGaoGGUF6i3qUVpxs20ZOAZ4j
/lMnKSd3budns0S6+IXguXuYVZCauxNO00hzrJ3x7+9tuRfrDkPNUWsTXmz03fJTU4Am0SqteQHV
de39fSnv4NDEgFCp0HiUb+im9UeTWAsKjXQzfkv5tOcfXx0FWDhxAyoNQktJ2ean8z73q+0cKbt7
Fw8zBEkCZTI1ZpCotQ9EPzUToxNDe9qoXlijfdevo1Unv2PFptnXoPA1Q6KdqyK23bIBVud8p2+8
CEpx8LuaFBMv8D2r21GeshuWKZ4OCuVbntYN5/JVqlSJbRWGS9achUKYfkfow5GtIs1dCWvsnUwp
iqho5STcGDxWlxPH/4f+M/ZF1zirIMWTzJ8xpluRhlHFjjncBJKQgRYKWF931VwYrVqQ3auyGhM6
bz3aZP49g6bp8ZGfEma+/rXCId9leZscc8gJzO724fgfHGRe8Tb6NRA2npIKaalcONSI8QNzzHeM
rq3uvg7vZ9DemdHcWVjUoh7c8K03YQDpWlRFz5r2epxFlJ7iLKNIBG2P84NelE7hHaMKGHFpmJ1r
TpzzWBVFbZnXiMmNNmPpspAgUT/KfP7hHz8w62yeCnjGCtZcgZjwlGSlExrGMcmzHFqEcvFA+Ovm
HoG7ncmLPdyi20jqiGtDLgY4zTPvBUwn8yTG1l3KQGJyH6+n3WdzKRXKlgrpGf9UjbS8ahlgv3A/
LKMtFM/tpoc4kXoKN8UyZKCav7jK4oI+4PMImvGjsSlyYK5NX1wZ/gJZip8U0YdUuVK7OlmavPnT
ZKCiWfAKe/95zCmPepEtJ2fiG+UonTQw3KBD2Jg4uVChgKS2MCVATyblZuMzjCXauVF7zmIbEL8i
99D6PI0I4JtQhJgCsZ1DzmRClm5geel1EiQYgIWrvOv2L/FAyKe/2nzDW5Fj0CL36KR7f9Gjmp4z
SMUAVQEtVTxpCtXCyYAmIXb40E5ZUCHnf/LhOZSGzbgwJdmy0FERooe/nT7aJuuV144BIuaxk8FH
9zBCWdajSFhavuCM31fRzBV8uShj0EFe8YfYwZaZRIdUVYghwbl8tI33eHrco5rFhbgWZ3QZiSbR
4Utj4BtgfU75Ts14HyMgLJmKQkclY+vTLRmz7Yf3cC1KaOvtpKMx5s6DDOUOenzGMareYn3rpB7a
zqRTsUB0GESzJtvC7MQ4xk6V3DVdCBaPb9oAi4VpIzBkmF652A06hIKBJTVFgjPMp9t2S6VOm1rX
WJm5mfz5JnI43+tadd+H9+Kwgfd4eRtGEeSP5EBH4X1e+RL+Fxcausm7KZhKP4yrnM0HgURbiqO1
TSZ9ob549y7Vs2CrXUKWICi5HTKFQB/VAltw3eua5UeO0VE5z1zG02QeDC9x58WU3sODWgNSQtgp
6xT1o5d9F+Gp9uYpDMHMQIPPTMI8+pekWpLXTaz7P5i/NoLmHzZn1teh1v07Jy+J6IdYCX5ZzbEV
0IBfwVfBV4HCvsPUNz8DWXAiOqGhBq6Q9sg+g7NBp52wcjDOnFau1mBNTRqnFctqT0WJiCRiZAZx
1+aI6STrp99QQ9Qf64CNDaRnJYzglV589TpqUXHaT0l8QL+AoDXIrkBtaj50AjR3uc6ucvROmlC8
AOmJh4Voo7MiD4plvMqyzF91oeAMTdjQybqM/PnUE2436+9/FtqQVkBmOB278/bWXo8pS6YJzC5q
q2WdcKNu5DeWV5f163AUZvHB4ozmS92LzxeP0SPkLb5XRs0Chfyg2lwjKrkI0qeOR7/BT9A+a3u+
fIhtqTK9UWZ8qp/KkkOf9UgbiBfTvlaZLs56BYcXygbEFshAL9LV4EdFO6BsITMnqx5Pp/oehxIs
vLjacGd5MEcVvajFaWG4uJgeA89fkqZfhJceHmJoWueIiGrZl+WN4ie4fwrgBClIcKKB/Md8/o1f
jtmnwh6lHkGbfynPvuJGAnrmZq/BZQdaBIOhjjqGxsfpkdNV5RzWM6ryUjTzZ2dxaHjRZ2ApKfFd
OIN86zVpmiromnDoK3u5J5qThjb61FrkY/YqJ5d5iZIaXFJuU+f0LUEgqu6ibnmAoeSO6juBdIEq
GWkPk0s32gEhOyodkiFeqbf4pthGVZfEcSaWgtot1jEuo602Md01L4fQWI1buNMRgofCPv1e5ube
7/CLAUjfodfSQZGjqE9N3+cEi20694UOQ2gqYQyloJLixoUPsEwoFIGf+cnMyQBS45vqCmEY5RdJ
XDRFqx2BGR0uauvY1SHaZjlxjsXShSKfZY7IA8YRkDZpn3Lmm39/94qOoTH6obYsOJBLuWKd/MyU
pNYjX2Fk0cykI96BoOc8+5vHwiZpcKimfPnhy76sr3hD/D02qVwipLtLIruk0w+uxUGlS+0LH7DY
uqYLLWc82RlnQG6xmTDPfQk1xAMqp3H5tAtx5MsDdbr5oGX+277jwnpU52YPWKDF8W9IXdM92aNy
36bH+bVdrEbk7wKg/mmwPUsZVYE6rT9maMHx6A2jzivvJKNxOr/Kb83f9yfshWuwOAs+XPbESoEY
Ns4LttTX+cm7zW6wEKoULTGnRPG86T08qQYVTxibeiHnU0dH8WorQgY+1qVJpkWC3UnD+3ehsjd7
GeH04DU1wMMz4CsYo9Gtypu8r6SVosZ5CrMZzwdFUcIiETOUWY4LCeAGvYlB8ggeDcnYx1pQv4lM
6S9Z6qtHYYwMS+EX2xzBw3/bLkcnn1afagEg99jFovruzNlaDsTeGr9HTJ4A6VtkMR9NzcU6NUuK
LzX6NDOBOvsIG3V2RTRmY2/fEsuFZ7m0g6+wfndI0sP3gv6l1a6zoLsflw9Rq5h5SMZ7IOW7Vits
SIqcnOuxqq8POb6h7Fp+gfBdbH35sZf5/HeqKrxyMNwGcDx+2LBW7B89oikgh1i6rVPeSHT35ss5
pZYLa+CpZLdmtz8wJRuR2nYWMIRlMVr7U+9Az65eALuaAmGtjZhWgnC/t+Ks5d25dUFDRObwtXV8
9j3mV/buZZyZgn2Yqt/5cp4fVohD7bc+/EpbKNAsUX5gL80p17r87+vCmirm4i3BN/PXHBJMiHRw
8J/j0K0QjQhQyxx0nBBSDe+lcfa+jyaUSJVzOujSoYVHzuVwqd1CPN/N2/GkZeYdRe8R5Fz3CLkN
+P4Ea52A/MDWN/d662ZLmDEMY5bYPQQqIDTegAbb4hXHBMWof27c776LCNYPngnoQ/OeiKhoUReT
T197GwKB+4DReGW/xnxFLI8U1aZIBJEmG/ct8ZiWrTDAlbCas8Xmg8+v6SvrVmDcvlAbO+T6/T57
ugS4Nd5yvqBdOxKeJlh6Bw/rbN+wSlcqJz5KDaJQGCqEag1NCuLRM86MPV3Hw1zk0o4Np1jurM8A
hSSqZlhejDPlFf1hee22ceCcK2C+9PO4vRvpcUBdr/NBykc0Ttfj0I/mxU3UMM7ffiE/GTv3KBis
b+lgqdnF1Wtpbgx6A1ztWQ0sxhYY0eIJ+70PAn3ViOqdvlpsWD2djLJrBCUn7cukloQ3q+7wgO1Q
PugEHvu8KbWmGty2gdtn2i1FVjTQjfkF0HfLgABPMw2VzLhUZZP0xbsZ2wIq2s80is67loIlvQGo
TtaLL94fGHzZAsyaCme74+saQWlbWkBOyrhURWbRCB3QhuNzNr6bVVCfWQ8OHAwWVVd9rdYwUriM
TWfs3jaRGqwzxaPcVNof4U/S/PUcE10X6clW+BNYAQ5EP3P43J1Q6LbSOt8RQY/NGN2tk8rduhUn
DRKuKiqknyO/wo75nwQW3yV51ryQOaKyBKa10O6JX8HBSgrqlm6IF3UD4X0+wq7rhSY9oaRlodvL
ZhsSbLaCGwqIe6xka1D8K24scAuaJoe0iL7wyNdEygOVxMx/GGLdutwmmJBa9sg2gw1LWUjOTE6U
YPN8wPdYZwg60JdWI07rro1Mxv3PXD9/rYlSpLMUZbQM8XPm/K7kEKKO4bxEjS8FNQ+4O/RXRaQ3
OKA1R4QwtISxB5iYtDU/Z0o/mD9yVQ9t2SJKvopjWWg/jaz8QPlfw6i7AT9nTfjwFmZ8XgJc2Y+h
T9RkzNfLF4ULysWNEdGn4Cdp+jPfBycfJdVOL3eo7I6aU/ACmNllIx7QiXzDMbpyiKi50i7LnYTF
VUJq0csGKq5MvuOF7xCKlUBXGNTSVWOkfaEtKM+uF+1bm2XNTQQhrCEH4v43RynVG2mC+GDaN6tc
Y3SRZ7X6DRUXlze7nXZBgrJrorPch0l6s+UXhJP6ZvuD4DyNBhYV8ZLv+QV9oC+Rfj7WXTLW9+G2
ywneX11mk4IeyUw4wigyYOsKsPxaEs5hPTgSeXrMQE6xbi7SwRfOcNUAGfP4pXSYZYvyr+j+V8C9
3+j/qpVmbFYVxiAO3bCKWxPnfKOlbBYh07/D2Xaeua/TzQEGro9SIHy5k8Od+sx4wYaH0LQxoe1K
a4JphgBIWUDYQVfukAwwUD9byyu7fPCF7I5PoTDddeqRtcjuCB6eTVcL6oX9+GxDRtl1vPoQooN0
GsFYaNkiRxF69XEDR/GDBbamOk3SxAooF9Xx367WzacP64LKb6yFQSig2dL1Zt5kQS1vJcbhSZlY
1t5heuk7guK+u8Tsk68aX7bqPxnr9FDmMrMCUzL2HxWTXB0nu3gqIQJqcFBKgRDQHR4vT7dDtXiI
zUVVGmXHueWl7q0MbL9gr64Ny1E4onin2kb1JorsRJ3RBLjTDlub3eChdGS3VbW1wsWuNixEWlXh
evm45eeAa5ZGqNOPEeSfH89gN9Q2pNUIePBe3n5GHEPLPf9cUt8wNQBVVxV2VS3uqzAwwRzWGXM4
XddP0pw2kJVkGza4nvCYorZVpM6O8/3ucoavFbvzaKETd73aDGRUKoHzYGZEu2nBS2Uq1aabzSTC
9GtrV12VC5P1gPG0rpiLHiZZBkXqelUOB2dJfdUGJsdmkPH+TjpW2VimODGiK3qNxjXJjrM8qybQ
9B8fCyqJrCbw9Tt6S4ECptrRDxdulyXoB+XUh8ewjhg1gc6i/bsVSuvkig7/rFkz2MZ+dKrXRjL/
5bElOU8num/utArw2vwgfo5gnFCBG6OaOwR0hAlUpw5DIYAzY01911FoH/5P7XHIVfCVo8kLeWed
CaptKMbe4eGrZfByH2s87RAbylZ8NyTWuHCWdd/CgL2i8hTQcEUGcvryZGxrUagTIoIxTbdtBvFV
pqxxOPfQ198aWgbhqbIWyQG1MfbkjsQ+YH+1OhHN6RnN8WMkJYaOxMAqbrYkwUjrVkeY2EqvZIwZ
N0jr2bPqYECm0xMHbTSbigqwv6mCEQgxNLHofGckbpTqXt82StktZ+P/pEtxBNyzSLXdfrh4uJGR
BtJo91rxl8nrjfl56ZegQOlJemfH+5adt8bNtfQLpygfV4B3mZgrFLRCtLFW7mJhk8nhIxfg43c4
S1ZEms8fTHHTvkwwEPxMCqpogkT+yRJO2WRm/MV3W6aWkHtX2Ghf5gGb+8hX3abmDoaAl5GIWEzN
kYX1owNNz8y/kssFot3FcHqBeZZ5DdEFTeVcEtpYMggAFHmnxp9PBOQYjEs3K3Kvt8VJR+L0HK4c
k9CNx8sVjeZ79buXx7Yk4gCxeOFL1qPJAGOAe7n+Y7KzPck39ah5Wp7JZKIKyrzJLRRdTvYiQ7W8
ZvWSmlYAnVu6Ip+8zXvxyASlgqb2kTXauVzCS9Oy5EI6d2yJ3QTuLX7pa3pyldV/OadM3SN105hZ
9hr+pu5yiOZ3Wbo5KphFgsfozYgjN1t0548rAgy8B6ZsuT22UdeFj46ooiAnYdBTdMfz7OsbpQHK
daM/oxR5ElnXgaRa8oqhfg8EWqHMKx4LkNfy1QG4x+PAHzUOJa+7HpIBDbLlLP1H1pwPcmTmxqIJ
mhU/aCKXpfBImj91K0YIadU8/z82JOQBKOtWBL6y4BXqW6TJqv+Kt5/w0sO8axw0CXuD0L1H0Aob
52XBp0CQwmw/1jT74RUqH4zcH41My6Kbv2g7f8pm4ZGV8k1xxT4CQsUsoERjmwflXaedFlFhQKmQ
2eYNPSrQ9MC6yzdyvkbb/WDXsTBYazIM5LpgUqXQCJGS8D8z8KpVj4prlv810aVuQAGBV1O1M1na
PVKJUw1EIaL/2daBccLyfUucaKsFh0OLGDRM/HbkGHbRsg4Lm29hOhstDDpU8A2FuRuf0LUw5ELS
f577zyLK04tj/+LXp5ufPAERmlERR8kaKkMwEuzkQsqnrLi+39gaik7B38N3G9VU1lsGLurIfwDB
s53TbzVQmBHRIRR8NasNRKqt/V+4IhpzdDgaM/L9jK72a+DzRh3OGZYCer6kCNlHGIaF7bY+KWCq
HlWczKtdBOOGLrItcgdsXq0y6VoxjLeVxEB9RDz0CLbT1qeYU9GjDsKFp2cbyvjEd6U5bF02tS/8
ikHGOn8cmzw50vgnbost10OhWS7ynVVkyEt/18i3/nKyCYcHaxUUmU5QgR8nPucStZQ1668Ei+5a
5a8n3X+fhnoDt8tuO8UObu2OpOJxmpPRQ7ZhiTngQooBHC5xYchhprt5kKYOBTN5WmghIr98aXWH
SqWJc6dfmDnEBChVWMVVSRa2ijq0z6eP43amhQdUN6SaPAreTaejgFcYg4dTmTu7nEGJODOYX10n
dHO+UIu0n7hrjTAjdyzOMC+jq9hNyi3NYSyEWsNSv7tioSVqxjEHwhU2pabIMCKqMXw/lCKpIVFQ
Zj8fWp7cEStoYXeJm6m9N0stdlXUtxxUPrX5xyPiWn0RaO4qdr91egDpvZzCbWM3iHs0I6SU1azB
D+nM4syR26+f196A3nRePrcYa7ehsaQOy4fn5QGs5J6G+hf7/4WzXUig/f0R9mcZVJJEB9A29LsU
/9ql9PghbHA07fiPv2Ry1qDRNQkFMqjh/YIg8CCscsKmomIDIB5lK5nlYXmqDNI8o696plbaurgc
7MWA/lVFf8vWTzze7tfMl2uaadpCAKsQY9BBtJH8LV3JYjJoL8YoJLkZlijGnvTH5snaE3TvWrbq
NeKbYZPShniFOvol9PQBf7NFpc3bXat39f7vJg0SEZu42wKn1aFVntCYfXlzUt1iZFZQfZGS3Wdx
JXmwccQ9fHCquLiJcjcdjSSbgPSShGzBJm+L1d7YHcbQmDIibnUKb0yPzEklGNJL9vcaOxTGIREU
S91HUClYuUQptzL7+CsOSWsy7poKIQQ5YIooUcQX2usryQbs5EUACP66sTYsDkQMUi50EU8JFR6M
Ui2frGfpbHTaEw5v3pSpGPi2+AbSvcPC/KYY+K4lXqcx4MjmTil/mv0lvjkyyUc7N7QM/6Wz4+w6
U2s0gwgCYawJ82/J3iiieg7NJm33rUIHESRq40iHHiIn4GRZC3yS3u0laQJS0EL7/J4qdbueUu+T
ZnxqSiAgmk6bKMw2ajVElQqW99XR6J1hIe3kiRGcVxVE32ITQ9GedtdGbBh7xIROFGNhFAgaZnF0
nRw4srH0W4TkPnX7t8Yq7yz/+WCjwQr87XWAXcJE29pbC53dPjbeQnCkNiij3SH4j7VdR2HdOzE6
6Gg/W2Iqa08ObVORETs3+LR5kFU6ToLWstXF+U4/q+wNwPRlyaMpDYg/zL8eV0K8aWDUmxhauXOq
jYDVhEEGwN29YsNqM61rDkhss15vNARz+q2lltSwTAzoA8ht0Rkhhs0tCyIodp26R/zJOOyIzq3T
xZOUQ72OUEAu5s+pAV5sTpN3ta+2JgHpiBOMtgE7dFgGXEKqebVr1M8IAWJScWIVukoqW8nT/iFs
b2wu+WDyvmK4sL3DgHFqUyG0tRky7JOrRSauSlKKMBbu2Tk8qrpyMWaJ545Oq/bewwVl4B6SK4Ac
DrLoDSx2irClj24Eu8hIT1GQmTuPjRuNIEYPGRyArfYFszdpPRIIG69EFTVx9ptNqQaK/fVsPNuK
wZyiAVoa/ltjgq1V9M8rfl01JJRUwX9vfQ9N7P6+LuD11VW4T6yVQpv/9VY8+lNUruLX7qz98Ukk
5LRvKC7EJh7WAbz+bGqoaUGDNzAw02NgX2aL5dDN8Rbq1M4QwuJi8AJAybz0RLASQ7JSiQsnKsyh
nwMHQlYmrvsq9e069PswDrYlrlhYQHuPF92/clRRZfP8DJ83LR+ds7BVAkh4MbDsSLTd+3j3Gbr5
NnhMnqE7OMghYjDRGWiRhetEPXi/AFBCWxddICC5r7FlDlV2VhC9QUg4VNm0yrYDpJffKDpOX5YG
Z+Hz5AboyHEZ6lRrLjWrL9HiQATa2XSqqEQUIQQ9Z+TqQrcEL/Ur918dPNC5QfIannMH+CNKsJ14
bz54zAXWm+OMwMIasVCoy2dJJRXX5EiK+2Rnnm5N6+AOuCWOKxQhfUUVJFs4vTIeztA7KG0F7XMH
bsDO3GzeXxdZqZK4s/e9e6saociO3/81nR/+0B8RDk+sVfUwMvOfE+zQK7dxvSQM4wZpY/ltSqI7
ouW7syLib1NV248SFCg0bUHQiLk0WjfqrpJ4oNL7IaCPmsyfVtHWpWeqB4Box9cx5Y53BHXge0ik
Vc9uRouiiCkYu6Q/n+j4Gc3i0m3xAObXVc4uHwHCe6UPE4MMll1/DVkMLy6382YYZvC0Dv5lhqgB
X/+UCBGYDPri/8yDslzonFQ3U3i1CdgZlaoneIGNJz5zvNXpOyFMthWFKySBhsJtKRONdGHupr7p
McfUUe4ZGfRoB9ifWPEuXD9zFZsWGTHQ2/JCdljlRk2h9Sfw6A6aWTMcgg8bdimskFcs+86BZVFP
X8OnHlL2+3CU/IoKcqMOXeuewPgB1x1daM2WOEjLj1D57X8+dU1XpASegy7dg8hqxQhYsnjPN0fw
UuM0uGioQ51NIcC1ozgyDMhaXnVqKWdbrdjv8K1Q9/oXo//vJ9/yobomEaixvOz/aYGAzsQ+C01/
5939E9Z5qmojg5vCpJo3crZllp7rdamRWyzwh+LBQIoMbzfjw5ZHuOTYejHKM33ig0zVi9ovxmfE
1hO7jmJqk5EVg01al2KkOXvCWiuTEKP9NrfqLGTOni9L0tVZTxguiD3QgJcuBivFmcR2CiCcFgv0
NLbJaZAwOEenYi7kAV+W2RMNFRcyYgR+cnOGzdJy4Z/hrp2ucXNgE3uheaxQTIX/lB6NK64fz1Dl
w9sU8/pQZhYASjMOY+f/6DPlqqJOVUYm7uSsxtxrx2vijA0Qc8mzdJP866Ud9nYmXCa6YC1czGVl
GizmkQ5UIsssen5O6WJ3ocYsHJyZif7y/Tm97TkiIiiNeoTmG1vMgkuwBYhysdEVTZMB+Pp3Waqg
QWA7JVrE9K5fluFviASo+9qEF2iNfkxwMBkXvQenbbSQvzdlStVionn9kGO/99sFtAQdBmC580Jo
I1rA/WH8BIC9akBymV8ThUwXxZ8xiauCYHZuNACNu0FanO0nY3ecU7og2KKKT/forc/qXS8M3Ahu
j2KL9Njo4uJFWkI7nd9pnhFaSVKVVUqDrsYhUa5amLoD7BB7Nbtpb+W8oE2ukVZZGnH7KSZIPvkl
70ICAmUEr9U6KQVK55N2novEt4Ei9irtloUqFmWVNUPYvqeavrTg6zWJ6mYpNHVkTWQFs7CkJdBA
I9LjbXivyI7NiaxnlWCDhjW2D7hV8lsLW93qcnUp8qcZmExevIF5DjE3nteeKrhpa66g/EP0G5Mx
0rKYtJxjEbymsLQDvGdfCcuJTZgT2JmGwNUik6WG0VRf39MkjLfGz7wVk6sQb5NJQ/51WkxASYH4
/4ubpO4AZxj5PKwCGTCWlKs+IzsV7Im3xjCTsTVeOUfczHokmlFTuA8WVqG45swtUDzO/xkwR3/t
ob9m0ue1mP244k5AmooA5BGoh5WNyTvP20P8NSgFzYjQmyf4q6WDNGfSc4UqdysnTTWeYapTgzJ1
iyivVAqPzMN+B3NjNZr/oW6YcqVDvZpskeyu9cwXm5lNYxeEwjgkYlu6HT6/i7v+2hRTE/umRwfI
XepEobXQNOnCkaaYmy+FXVtjxgl4lvu4LwqJcG4DtHxg+ndxz7JFhI2o4ENeLc3/trdrB4zbpM1k
3s37IvSLzVSRb9h2LQ3c88K2jLSLr8JB3uV/EztkhWdCBNdZ8rchQtwMlqgbvoeSDSHlUOFdms2L
mJiofvH+KMhUwlHmLfK2u+sTb8tKfcQl1vAwqj0aomR2HPPAqgz7yHd/9nX+iS8kO5SQogbQrS1a
9/PqXLodKtH3xbWgCvfqULawguX+Xs7t3IFjn2iyvlRmeD/kIWonYUGxZxNmBrqFCNgW9/KslMCu
aAXMFkqY+/mfD6TLe1ov+LU8G3sgY2ruCO12ULjmjDOaVV+4cBPbBsQjT8l6/PfbeP4f2IXXd4s0
6HFsBtI1VH0ux1bBkCrZTG16ai6NNzZRfLC69b5jYUs0cS9ZBglC3/6iif+lcn7QLkugun2SOWFm
AwtVUYZDtGbhtY6X9F7m/S/g7pyBA7dfrP36u6/lQUyvafPeJlGgX/YeLYtsYO8Ndp3UzKiBxFU6
hTsw8Dec9wMd6GoBgwPxSGX5wJx6clI7uO9KV8g1plPQ7q24V9FCybBJMjAckLxhdNHb69QBdElO
2mjONjhvPDmy3QKocTyypoTrRGzSEaMl5JyTaVFjhG1nUei5jvQAHtuEXDsJArJZw9175njDM+DG
07jGYVGWJh0DyLb/8CJthy3X6eEKeL6om6Lx9/aHBMsNeEQ37KtNPehvLvnlUY7mkU35lIRF7O1J
7ldxBNcURoUhkiLhshq/eLK7lw1gazeStkUvbGuQUh/KLLb6ForD4rwW37mYJVDLuHczE8Y5E8cU
C6iJ/tPPx375gaD1p0KMDru49GbTkTBA39FncbXbkXAtsCuaYnJTAnhMQglcByzW1iGk/0Bu4sN4
mXDi5jYMAA0PZGZOR6DX6xJVwoONlUNGsz9NokHqClvcu/vXTWG0tfkQcsF8KqU3P8JMDAxowpTs
qx2bxT0qg2OM4zQim05oUmpqR8XBrscdZaqTmLxQUivtCRu6nMBhkLZipXXVOZs90EqMT+hDFEtB
OVf9pEOFqncdGlfW8hBlJ19jyXLBPJsm87TUJm5CXEBH/wBMa9m8Kebok4YcI1zfP4b2RaSZsi0C
PA7IvvalxakAsTYbTbjp/LMahN5ko+GTIUeVrJf91rbPGUoeU+kINJp0gYatQYwXKkkXYI40qj33
Cras8+8Eqhy6t8KfNs9GqtVDtrawsG5WIpCa6wn/X4J4e24cde4D7U19Yc67sL0tKcP4vGI9TZHR
ttYuDBwjgZrMYCiE5aIGn6duZVEVfZfsV6zPNH/pAVrLnQ/lUpH5y/ks2aJTGgM4SNbuhIl9Ny6q
9oS80UMCT9DC9QA2lYHp4BOp4iPhaFh1wm6G4wPmZ/gnQ+DJQwyQ5VeLXCWosKta+OnfH/0Z3yCC
Fkua/jdWmCZZkhIf6zLg9gIHPp4//4PMtgY9IwAKSmpSg0R2xn0YzlntBMG2AAJ2fiPImcIPAf2u
XdHMbwJm5ffQJmzDcH4nGvCFtDzzbNc6m3wQ73c8SXPCW8TGf9mu0z/m+mmA9sS3FQ4MeLcw7xQA
2EzjFp4Xo9PAE426wd9Y1N0xTFo+TTu+5CMqWscsP3HVzz3jpkyuga4QVela6Y2xmVywaJFMSBcz
D0yJRFZn91o4Ap6gSw656srM0H4XD+EbGqlrekpE6ers35XSSNnvGUU0Ripe6uMs3f6/xmmNSrOl
0gi+QA5n9R7+fs6Wzo4oTsJrwFPRmJ45Vjvh6D/X1wUxrUZdpTmyu5J94oqxhRhBwD/5i1aKrivu
cSCaZM8567FV+ddx2ot388v01A+/XjNPK3rEKt1mSg2a1TDgwGBbZGfBIduty07e5j5rEZC/cfsU
xWla5J0xIDME71qg0jVhOYhG8J0hBEFFhUYakeTxEUWrDT/TgxVA7rq4k8wgghtnEBFDzFwL4hxm
c/khdVV3YYwWsnuLVNEAFmecr/LHpusGwb8BEWiaR2d4AlGg/Ezo3D6RpEbCTp2uFMZVn9DC4amN
dTbiDt2zPrE+akDzbXUDjUNHZzCS/OtW8l1ZvjUbSTmJlTacvJFzsiSz1yBsPseOPX1dRLzcGc+B
xGfQYaffDQgO+NwWhtkMndEPsPEg1399YgK62+1ttkMvS8GZFrO2ngBEJrJmGAol3l/LBfXkUwCZ
MrgY+7lKhjqqhigq521uSjRWlxytde1O1bIfJw4sxoq3taGx4M2x/B+J4dOosY2tX8p7jJ8UdAp2
fntaJezRJhAS+t5Tfj0s/1fiIFNEYE4vTMbaqMn8c1dFhmqa6AD7EqSyORjxML4nGY/vV6/Si1to
duFIz4iMgzFdOeVn3XXdpIF29ta2tEHGt1brCZ/ZnvrUa2rOXGOngwHp6wsgiwqgvfsCLtH5v/Uv
LpJF4L4QuOCrWRrA76HP6a02papn16OGHAHrK9u1PSmz5h8VSpT3jO27G5PHgdcxR3mxk1djQ1L1
uRtcWOpFAMO5CNfm5+2Aqg08gaBDkaBW4jvaOAwkHkNY1DjqpPwLOnuK1TSJathWwcGRs8vWd5WU
47oC1Kqnf1joXSzynSK+R5xTlKECCbMDPag7nyAWKEAvu3B3zcseKnu3imV+1Cv0E8CUTxU7Y3JQ
EEMfDnknUnmmA/+rlAwR6utyXbRyqoLL9FEW7gNLRySE5MaE+5EJFMrHT09NnSLyhVvoEdkDejrp
/O3eW2TyUYnH4SWLr0lOGap3YSl2VgUBo/uI/mZWZN+Nc7u1meeUs7TMdNKKrSSFP+wgm2biYFtK
pBlyp6nvL8gCXVRk+KbvXtzM6HJeg6Z0JigN620I+8eQH2N+MJjDjnCI5L41hBzF7jqVmd6lhIMP
KIboX9kaJtD9+gTzX4ogJZ+ewGj7aL6lYmwHC7NctETM82LN6WtioJnN6dRICZnvRc3d3drOaDmO
y/xA2P3FNXVN6PYzMiXxOAURYUjc06Z30aG/u0Ro3+/vAFKVakQfb06AjcFTolk0Iai/B2IZ4u0J
Pkq7ofIXd7CnipaDyVe/et5+iRZhjV4j5b5uZpWPCBpFGDgKZXMoFj2HQyje0LR5/w9dnOoRN6up
r6lkp5Z4ftWolb0jO2sgJRhCI0uBTpwTFJkqiP4YCE8NMXXvd3XmBrt5r7IXZYvdpo2E68lrxUPt
/yVC+tHv2U+2zLXFWGRmG0jrtLkchdi42G2D5p4Vtx8ZS/GMkO2sKFbyFuayggbnlOFZrjv4eB+l
2GcosTXxX1npEk2B7aC3+vamG1mreck0eBNl20QjR0+KjrPNhUEEw7qhBAkepT6MHoT1hvsfxMWP
LR7pUKoitAcidNlNqydcitqPauYGrqNu7QOg8dho5xBbCmfBIdpstcbcNJQ6Y0FllCQ8tfOiGJbN
PGnEoIvRhdZDiCEKCw+cw+R2Xw2rLUqgNbasMsqbSiTOlmT1KlUrxPGkOq0ebm+WGHCQNqbbLlo3
0U/fd7uMEapnAzN20wQ1qWB/v9BpQ7NNJBKKeYwZugwIftnYNMfS76DzpTEgIm/3EcFqSFFJMDso
3621KWvOVpIusSrTWReh4CDeCxdxWtdFMyPKmVmh3tvRktsAK97ynohMsYgWBbF8BzqEH1pS4HOt
J7mi9qd7PYGKYz/SxTpn1Y/YcuJY5EQW0dvQRPvevfKzL4/RXD5yN+zKtS43WtlZG7//D8PpY/89
r/S5h+NhBx4dMMqLz+pjMQYH57LpB9iURLkxKnitwGFM6tGQn+txDSM1oB/3SjmLGnws2Aq8Z5LG
vsmyVdcoADDb4N3M1uXgsxwazNBtSGjo6MK1JAW4gp8K5En2YMgF7qD57BDjSPJIU6aqwTyse1/7
LZ9LS+wuu+x8IKfaq2jSE6OWfccSuQ3h9DeRW1OndfN2K5yggSwhmEkFYsO/ahJs15aalxlzaXH+
6TQImLrr+IOkUneql98mZM78J1yFgARQ1+GYvGf2aZxF+G45Em9BuoW8iCOGEpi9qfIxo0DpYnYj
7sSS5daEKlUUW/0DoSmGL9jDihxYhD25SzzvK8z6bC3OVOQ0ZTj4AwMnd/6PC2I/9oIxLqjdZ8Mm
OgS3SlP8KcXLR6F5/Wv+lpzA0VaFoomhYYiDxds8DZSP7kQGFgvyFFDtxORoghVOodqEofmoGXvz
6hvJWi2YZH3sNl5EF3yHK9/EDTRd1CNDdvVWbSH2gBFRFv5C1WNW4CsEZEVNWdinlEE+iIn1dIB+
G/sJZ0Fzooh1UGwDz3M1yw5s0mstv4A/p7RzdxcaV38ujGCc6EwdfKOvVGR9dJOXkc5MyHuY7yZb
5Dp9CoU781L8UR+zHCwEjNG2gXfzpoXsQnZIOjAnNiIsBs4Zj3NdFkgSIdG8/Z2cgmw8Ua5fbyaY
fbioZACjFTh1sCe/sohy76hoFoXKjLw82QgfrJNJ3+nZI7YMKCkLPLhPCUoUv7mavAOMJepEA7ot
xBM/KGLSYqVvrc71oxzm/xtJ/ahC55ELU08TCRLadFqV0K4h+QcfXG2JypwV3nWF74OvWFWX5gGH
W5B82FxKHyazFYomKHN/SXAmMvqt4FKaQ8yLco1ZVa60xbMiCjlyuaKkSW7HpMgNxFq4VJjZd1IW
OuhgGPan/zvPq+B6HPK98B0zSjRnz2P6BkhZQp83zPC9DY2Dc+GrNRr7XxKGFlPRLCKqkf1O3vlY
7ZP1VhKMyuz9BcKiqIS1FQxXvdWiPZiLxle5CGUM20N8SeTXPYOm6cym+MBLHKmF7KmoRdT0RkBR
T5uTCgxkkJ+gBH9XD3RCux779dOJlzAI7dI9U/hW8puYuHngC5bq/j6osu+cdylWSLKukkpg/oCZ
soJStFbjtgmgiHxHrB0iCDBmMM/2X9N/Z3fgFKBIA7HJabb6YRguHHqCWYLa1vBGFw3GKQSm/J56
OUOPbQV6lU+Pp3PBb0m4dTmUmEJNaet39LDEQM4bUzVJjf3pD+qmrZNjcprFkYq87sbuTSCQmHPo
IxvPIzYSTkR9uogpLCoKlcHlb0nenVHCLQBsr3D3DhmEavs2AXo/a2xH0sx8fp29XIgLMFcTypv2
o3ewuplLATvvAcCDIxVgFd5I65+5P5nYaM5lKBvcAG2cfWKVtNRAVma0s8LBqXJZyUiWzAzvlrpi
xOdkDza/syvs0RYRT1oDOYSrMk7zMp2EyCg+yp7pDhy5oTTlJZZMeQS9HWyoSlFDNUGsHGpnecEb
mUVhdgybAREdMgvtNzZNNjOcmZN8DNZbI2S7CptCQw1XZ8/EgtjWinnizZL4vHZP6mCn9nag3kfm
dy/TO4t8FSkp57UoGVAXssUvRHwe8Sz9ktZQtwowLLG5Yz0NlGnqfp1R5Nmgi34AvAuKoXBzUSHK
4IBxzHIz+ytSHN5lQzRMWczjkpV63HlJkQE6Dtglv7U+Nh8gvSl93t/QOn88/5Eu2luSp+IzyfIj
ql0OBcQKsO2QLg1a5LYWa2e7iiI/0jB4TgC6qiYF9x2dO1BTvu0uTUDYpEOl6xdCf147bwO4qecB
s3d56brEDgXu5jRU6n4JO3UC2iqIDN2OGuuuIvWI5Bgnh8XaIz2oeS1zrbfXzXSIpdCVUlsvV5mL
9jxq+OWiXC+6wK+QhioHETKd2o7Tl5tmxWHqpAnQ+cOVxsUsJa4PBcvpTI9+TJkdOBBzKXgnNAOI
lpKvU2obXJw49srEixBy0d26NWrdaPvuargHD81+lZzYnA9HpUO+GskPEuyInygoDBV9TdAgz4Os
ZTbPdLpoVHSxwnOqQx25QjNNkWRJuNEw9wtjJhOUpkWGj2NBmCaSs/NEWltNmyhrQGuFLooNXxnt
kc8Nt1BcfumC1lb1m9OaUjrPx1eYke9/SlKS8310x231yT2Dk/NMlkEoRLCzDvmfdT9B4AhN7Rrh
hYox4IKu5sWlYyN9vXZ/+M5WqteYiLBxNmwBcGjAj2zy1pFYvdsjNFrAk3uVOl96ucNrD/cneV4h
oxRbGWm8phad7l2wyPL2g1VsSesrodnhE+N0BpPjp1ag+tnSPqgGMxdYVFtX2tQcxlmyEjdG288w
QFhxA7kLrd7j4YzLVRiWoI/n2xIJ67oke5oVoQckp3/3foXpNuXEgh96ArxvOAXeCIECob0US+ZG
CFnPkbO5w/2VMI910a4CDPjxI00UB42KnUPeRM6oSdmva0DrgrAaWWijMuAg5EAC9vQbOFkPr8c7
WRxy5DO1TNsAufqo2yRDaFGvYgOXrzzHCRV1ewdZ2U5GL4bE1lFNDHDwQQnPq39OIMjwTEhpjJp6
VwislRnEl2Nb+TSNZXxX8OCzD0DyYEnAeBzbD3FLbdbhSNm6Eee3GKR+0jINT64DOhfTdc0QdwJQ
gQ2z3er9f13oCemq/ZPjNEOX6j708Ostz6mOJLkBLjdwNGLdbTRkNIUuAjAejgVqLXZ/tUbKb62x
45rbx5LvdXttsalGoDmTJVKLe7YLXHgZMdDSbj48TwVRtHtmf+oux5pxGIZ2sR83/12Nud3HOn98
xCiYhfgKcLwSC+++OPYsPL1b4STJDr45XhKx1tjn4TDmQKUlZT90YL6wCAdwr4C1JJbxVebZhD9P
A1j9fSkmGRK5q57NopYz62MEoDuKR5szTbOY1XH9n2E/6jtTHkpg08heWWGIpCnLxCDbBU+iajdJ
AaeVI8zRc9z+UKw958LyzTQ7ukxRLlDgB5AmPYvK9TCEMc3ToNwEgykufmWH2Fl08rTsJhGf72YR
aITRwnyyhRh6BxnkKLx+VZ074k7H2g3GU40cLpq92jVByTwJ+036yRCuv4TSaaPK2a3674sMxPAE
zbHOpoGjHVYJwsMyVcS7qOcv9L3jwvL7Tnw939svBvVSh5WRE6kClFWc5cSUN2wGFExVZMgTREeq
YcWWDP0OYbr+bhpQZS0wHsa4im5gLP50XU+6Yu++BLvNZyTDl7vi46vyuwAo/4uA2/l3FNTrrWgX
lOSDsJjNCkhMemxcr/qtHjujTESdjDVSpkdOIeZyOQCB1K8oL+SBp85eroubwDxiBM2CgIMStAAT
FXOm01wjAr6sUEgdBao0TIOskk2IRzYedGi9fSySyXRR/+uMnzrduEZaOwBSXIGTwzNnI2Avnm6u
pIIrT9lAhoCIG0rPiC69pVp/MQgvk3VOv5c5TYskUfowU2LAmuFw/OYu1OYHU+aBeMq0M/bsmp8+
zX1sXjAZsS9dL7bbSDV/ga/55H4rvoazli5pLspA9OgKHQhY9obtqAmvfqCWmMqDLdiclLv7m3R2
O+aP9YBlAE+S0BRbWsMMFU0CCew2zyDaqQiLVUYp8Ito6XM/lNEJZ2eHKur1/9KMoA8XeYXYp3c1
kcy7hydbvpgMWqBay/xSf4f/1LUE1F7wS6ZDMiRTMDsWC7OpbQ56FRVYQ5WGwONuz19nLXg5o0w7
rf7+X2VhlOTXE4geGCSDnrnvFAmXZ9qfnQv8JaBQM7DlF3xlG15zzPlW5ow8EGru4D/rUfDeEGj/
15TKffKRiOErU3SscHJfdlAfq9GSGF9R+dovXL55e9Knzh978B2KZYfdHbxRKKfvwkcxz0zlLkTl
d/l9eUe7JjIoNArpqrYTK7Ec/sx9Ju8o/B5sso/YfBb0mvYRbPoEfTR+TjedinelWz6ClCWRTwGt
zC9oyA7u3layhQBFrRh3vFuobC4YaCRceSzuI5e4L2THvRN+f8qrDZukeUATrl9PVNIl+url9aey
Zp7m5j4DX/kzyxCUdXsSOFh5oLH58Z/Da2RehIQ81AKeScEE4113Fvr2Z5scrEyPCgpM4mElk02+
xRI29KP+JsJNIM3merOSGDR4zJC6hWlSCuS/hFstnQBW46EVrjvkfJdcIQE8wLZMQgMMygNBBDvs
XHW/iaf8dXq/KmktlUWW2UKXkVt6W9tdGJ/iUp5DvNnFkM1UPRDhg8pFSWtIH18xWMHvU3UNPP0p
tinoDNe5Ang8ZDSesWdUYX/W9PvfsxXMj8V4Uo5+g1rtUDgm58rabiFJaZfc6ERu6TYV6xFtvDHf
07zTmnlymPwA0l7v6fHcKJdEbghrdRfW6VpIOPX35U9bY0rjJgllKMJ75eeDcTSnJiaXAVamThT3
Eo5blPOqNGjWPhtV/phpw2G6jfBJIxDegQG3J97B8mxQJs5m1Rg51mcREZBnJZ/pp6aWmkmoiMNI
CQ5uH3ajbZyxocDUMbjEtIfZWouBSGu9+766jw531p3SWFyxyKM2BuqQQ2t4u7R973Q1UI5yiy/u
o0UkTKJK+ttd3mjPJy0uTAHMjfWpiW04njafqEMRFSH1vfhMIIee+2xybiWjtGcNwSJ3NsJ5G0s2
XzyuUKpiS2V+Nnphr8bHAaaBir6gEzAokMgqxOIxdeXzgEbFP1nhisHlAdddl7uMPAje5pKvWXUQ
bXejivU/hDAx65kTgjTSnCOShbo6BhX2JchA39IJKR/XQKFAGgIIQs40WnSMrTc2gTSRx+i0q2vI
b8XyLiNwWLI9lbmo83bKBx/wE0QmXYV1WGgem5MiJ+2YyMo1BmuKc6xkv4FOiDKmyLPz+1yK5me5
M9ORj7kDjh1NsrrkAhl7dl1984CM5yk15UB3h4/ZchvT7Y9rZWB475wHb8e1PQqxyEOdPnnGI10N
xMqBDqomGekCP8c8CXqh2dyVKGA6X2QUpSAhzWwiZ/EPYnooW12jc6qyTrcO+KxGa8HtBhSkBzmN
A9j3Ei2+ASgeQOWIq9oMRlEm+Xfcu/PWLikOEDz/dH0SCXAx5EAdw1knjQ0Rog8vGOXahCsmelpT
b+ttLemwk/NCNSUEJO7+FyeHqmjn+mU0t6hP+aefqjgjdV+8PAQ/DQwy1GDaWCYJN0NfAV0Xxih6
2xbstCGWumGZOAJmx6sYxLj3WvP1a3wrp4H+iLalcpJIl0/md5r6jP9685rz2ftVEynGXmKVuPZu
xir2A4Jqp7kN/B0M3rnJdnU42xf6ZUabIB3e2E1QC36mgix4WzvszmrubujABfrYk/4sutACJa32
F+WXrQRqbf9ji4q1K5OShuRK4ZaQ+oxHNIcDgebaN/e8WPa1drpp+ICiBLMWenkBJ5pGSsem11ng
fKH/Ik78bg2xUjgvAIx680Dv6jWuU4ua5uLQwrlBo+MarNZ/U+vyQLEEJSOQcEwGzk4JArjSMRF7
bKYarMD7coVL5JpiIf6b8UcjGEq37TSC67OugqSumdFEOjAFuU7FpvCl4AH/wFR9fX9z7n76cc5m
XP5RnS2C3zNzTcXtBm86yh++EHHHSRqFB+OvKok4wZmnZh+P9H05asILp6fkOqowLYjTrOu5fT64
DUALdLPGriZouIIP8HUqNH6BEIpi5vvvPgOHbmCxTNBmqIrynyznhBNTWTr8uT5k9Cq9jK9DG2yj
QH/ph+UFbL5cZ5zAnc82VVOoYo8k1uLkhfpMDVlRUtGk9ovnZcYFhyFLHNmD1LuUR6PFtvS5i++p
7vNLlzlEJxL7ipUNyvDe3YA1so/s/vqoDSeZn9b4UNVQiOBtogxlG+4Wvqrid9G0BPzUPErfhfiD
T91kItHs78oFed7TtjNFhBwusyVLmOCDHONb90qHxfhOhFtAI2ly642lcoKtBNNgi2ihcFuG+z8z
dKUzLqPwfgamuoZ6Y+gFrAWlCbcytsgl5uRzw7xhHDF89r1smupEplAnUgfJpRyLdEV0pP8xDeBK
7eVvzO8iL5hA18bv49bWoiv+Pq3IzOf4RZKMM3gUDV2H+Pe1HYIo99AwENSQw/INe7ZfbZ6BtBtW
+qoqcBOeoFz+NlPdjiI9prltL8ZmaId29BwEIVLMRv7RRu0AC8tdiBrc9LhFQsivS0r/JbMWedDz
LZXIX1VpMlXLWZ4G/3+dR8v3gEXeKn0rANQcv0bLhQ1Kozdkcp4jsyEDCnRnM6x+kj4ddaH71LPb
90lRR6XAwRNy6xLOzVprfs53HsNKwG5M58iJp62HDefp8GFsr5uFqfjufGP4/gbuBGAVSIgqEnO3
JZO9VMgMv0jG3zo3ewSbrK9WwPQcMMpXUFA+z3Vm/4k0dRg1J5QEWOKxkEtAyu0+C9dR9vHtMOZg
l1XmNji99Liz+kcaA/3jgdgz6YnHFGbLMUf+AlaSRuaje1aivjy+rwBohSsLp3j4u++IQ2kaab9X
30vZzderzvC7VnWtGn3pEBO4YPfltqbTd6rEIasbkUCkjAMCiTDi6efubtcimONxBDGaRQUBzW79
+GMu9KyZF+mbUnIkKh/EGYsDcR/CT4bmogf7X+UJn3lEXejdP20zKRd9bv3xjupB0QKwFjB8TDTQ
9DAxgiSxILo6/jEpPpEeuLROavxySnWlJ1xJFIYBcP1iJYIjKGS1qLh9tRw5R67m0lMmJbYvs3XK
1z73cJ7qZP7AQWuzpowHS/yR6E1m6tBUUkQ2cMfPhZtTDFiWvJzzTZkg3hh2QG6OPXqnvYUsoudx
DUjxNU7ErSM5+8QOetUbZruxSRGinm2ji9QgfeE5TxzxfEIkoeOLngy+MwWb41t1ii5pL9qG8kkZ
9WDMBJ5kGwlUDE6qO+61yomTfKo8tTJH8NkJfBbCXYdS0GJFMuGmpCikkibW1gZN/gM5csyE//TY
Abru/OSbyHvEhUMMFf6Nm3LzF1cCQ3PF817ZZ31852fkMT9PzUO3TUb3WzDFv5f+1X+h3CmcJquw
KTU3t/Hq06T9WjWjEU8DVlvgmAiutf0Hgm+8SnYZUswDDlZ0Mf1o59Q5+XdTsA6CCGmlDPQimKPF
gB9QgfntdCUKybmPP80U8sWCRcWSv0mYUC7GKNgzjCT+APs0nwD/OUAI6M32PBvNsv0ywt2ttrml
8pdrFxfhYzi2HZqucaFBHm/q1n3L7aRsKOQM1WjPSoGACc0PqNVwXF/P+w5J1cQE7kJ6lzIp0ROj
h6oWpOKxmbB0Xy/LCsrN9Dv3H4cKJctN50wWPXv2GtuyT/5U/1wEiBHuE3cG8KvlyDHXXsykQaDD
nnNpBVlZZyb7tosOKgoELd1S/vQbFXrSJHRYsnCiDrSCJiQlAIAfK+KcyrMzhCQv3v1Bi6A5jgSX
oUoywL1dr8TURPuuO8Cv2QZYEQP+BAxmoNzB88bKPz2TI7TVosjCNioGcqaeaz868VoSWoG+N+lX
ySD0jDnfiWsbP6Eju+/bS6k6AwAdDIHMNnqkYA0Ewdzg8fWyB1zGUzYT8guAhzFX6XrEtW6u7W0e
v51fGfPXOVfGYK658LvCrbDAPMWfaGoJBu+xgwcrk2auWinCQmVh7h7qRINAW/Vg1Cr5ktYT+ldx
0C54gKy7K7+bbGsRvzO4fs7Zm5JMv4CrCHIADgZMUMPbVJGLofwdCWD4ERhF9/s1EUYGZK5QVSXo
UfQL6fYo9vpkpS4Nn6QBwiqSEaHPB5lDGsm4iC0WMdlh1ts40Gqi+c7/+/uSyLkyHf78fvlyssb8
kZHRwWkOc90Gx/m/JnmTkDazrSK4Y6ZT8W7ONtMo+cVXhxKbPTv5hMffGhcPe7qWJtNSRSyHNu3C
NU1KhWcN5i3ZFSCy8LxgLGLm9EBbUIdH4vLKLnJoVfuxslCn3MV0f+x/OVWLR9jjXJ6SwRN+PhRQ
CCP7VdS7S0ilNvZNDeioG7k6QyA4rAdpoXhNgvCQlj0qrFcxluRHl+of8L91fanQL+pnNuGYazBN
lJMdKK5bH/tL/yDTTUIcl9UsrFOyn4nw6nKwd61OVC78hkp1PxBsHI8Lux4cwJcmFNeXxrQAOzgO
8l/kWzXL/m+UrizzNHApzi5rxrUqtoXHapHc7OqP2aj/AKy4eCkWczl4+7p/BU2CJzCdhAv4Sey7
OUdvmSxol0BXr24Z3AiVO027F15YJdx4Xd/6v4PyGH6YS49+emd+7GaWHWrgKpM8CgwAwBNO6xCD
yl8qtWYGcZ4eRj6CKCbfv5U/uQPpcKPyO8D45Qav+I7r/PD/D5Dv02dhsbHtfwMKU/f6bFlr4V9v
uXEqqTn+3/A7RG/V7o/wai1NAm5r+atAaQrG7aL6A2Q1Z0rboc4bwLnMTvxHASOcDbQg5UXlvTCq
ikq3mwBSOqdh9cHUxjVTCYGMlrgV4maXmhT7yv5ylJImXg2TPyrIszeZt3scjyAfuY12RP6awDA0
mYZtNADI/9aBPNk5ulwC1rMFV1ioLohGbVC/hCWKutIhI+y+pls2DxCM3hPMh5htdOqgzcixNHx5
omAPR1O/8Mxz54iK30/lVDGXKZcydvSc+YeKvAOpBy1iK3O3CLBON11rWnAfgXR5wFOkqLidnMcM
mX4tD19Lp+y/l+WypgF5b7Nq5V1HTvF5FoOoFq1PZQLTPdFZwEPGYFzQuxGoNk0Gdj4vayx+5z2O
mu5siO+avM26uWnU7PQ0w3cLKGY9qIODH+FBDZeu8ttp9+E1lGqRk1VrM0SisptWV635ogPe1dDs
HzY6bA3KR9K5eFci55nN8x2vjae4v//xhj87HMtH0RnX2Yn4nz5lKzhU0/fWTwKNIjSSmP0+w1/t
hLgZEbxpYzF7IhFegguS9PmhwFn3LFe+f6nQOXciA7o+qbeF65JexXG2KIPXjeZUXYAFTtdd9RJ/
It2YyRYqKGO3OWKNMeYGjesLEOxFBOpK2k8hD8WCbmwayxsvWPm3ZvvsHvG9DPc/+kTYop8Ff7Uc
I9+tJPZ38aTw5Z851qXwwITYy9E3D/TSFp3c2zIkvS0g+CgUYN7+ZSuyEUrKxr4+tqjAiIIqIkKv
yxzzlPB4mHg2661PW92gu3GxFODvkclGK7VbiWQvS2jl4LsFI/9QJsc3mVsVN0uXcat04IQtRFDk
1wCCGlgpzCTfCSDYiIo/p7B0tu/S+AzgsvT1DMEd5lpuE31Yjj1nl9PiPLW61WhLk91p0z3YoTWP
+oIKjWcVQoyMNYdseJBbhyatJZTPYWyqfuGeB1DfZMBLYN+Oe1Ggf0mfPAE1T6hKjUMmB37zN5Dy
JdJqjviuL/lXA6+3c48QQpg6bXudpvvpFN1UwA6TTUU8q9uo8t92FSEsWR/AkH/UE2CnYs5yIc9a
64Rz5nI5WG+UCeMNKemK6N4qK7szf4GH4HQI/SAeUHiW8sOXqgdnbFjRXWE3BQCTOxNr1G0M4x/K
bY5emZ1INgA1cA4sJRguSxN51T+K8sokhrFGTPZdKCI4rGHVQT41TBzEzrK5OX51kFqO4HumcLMd
0gLFN1oGbfYoDi/ZLSF6q5cafWK6cMEoFo9JDB/6E+B/BTmws3Ge6rrTvPen12llOZeKoQKcWort
4C8tb1yUSYgzByrmZuJKbQn0rg3vvNX3tjk4sQOCWNYYMxxRx6YviP9eOfGJ1OOspKaZ9P6EMGQm
tv+69bmjrrXT8jZKrzVorpuSdehRDGz7LuAmDuFHTmIJgI8PQDdkcfmHAwSGOlJBiYxk9nG1N65U
DrjwzUJ4pK1CH6fFmKUkYbk3EyfI9318pi01fRJUMIEboZ5D05vv3uqLDOeQPc+4BSiwUxCMHd3Q
r9LI5XucGFUpYhC4CgIxJ8OUUKtjpEejz7ehldp9MkLCRDAL/2x7px3qYq1sD35j2iU8R4RB8+rT
NRuWy+mS7HsZ1vKoCW0OnsGJVyRhvp9wK/uM7G3x0sl+twMd3eDMgmOSKLPMdtGPTvjUe4Yy/+da
nWw/7hGNVKoJvdUbshbbQPDQuOVqaM+5hIBSelWbepILbkDPVt/UMl90Eosdpkx+lz8r51TdyBJB
kXr3r57sW//JkVHW0r+RjRIZHEAkhT9Sbj/eDoAW70JEDNRo3fCPfeSYPB6tDCr91PV6/SgyPEAY
WD8ihwoDQ7U8TDyuhdzj0n4m/VDeKQyCTxdSdV6Jspciqm1MBwTIZWWVfIBpC83BNdifReVWFFSC
nil2z714CDN89WbDLTC3fcxeAjvdXpDm+0wzPoFfWLXcOtWccaKiYnjxI+e3UML6oPcAaKeudOKa
qgpOxX/j6x5P5t/9nkuikwfYXjZFCJ90ztL8JzhrFnzxhskdtCDJskWMdw+8WlesrIBEHKGCcvJh
MhKGKtf0zZJyV78rKVqM138+CRLRTAYMGXNJZCDIuJlvjtHq7sgk0/flLilCBPlMUO2hdh6CCL2A
RcetT/K/Dfpi+9TeYveX81M1iIQcaONQmZ+KbS4oFG1dwx2+cHsvXn0fvAXZE8Iyt4upaxwJksaz
xT62zxQ+jae0ap2DgWSwOPItRbi0mQyVC0pFCmd1sD80CWcaDYhAQkKOLn48sRAGo4TmRAQJfDOG
ljVZoQ9s1WjTZMf3zJFz5v9oLpPjeMPwxomB/wKOd4mzsaUC4mRhvRTTGueLMGXnq/SfJeH7lOxo
1KG4fBtC0NxEGL+2C/3/qfqutgEvwc3zRIjhXLxq+NHvZqW9ixTZ9pAjlAUCbHE5p/J7rFNo6MbM
v2BrA1F/T0UNNfjJQAnyIUWLI8wuEKdIikQC/sQWkNyaVs7WDRGSavfAXYxs5l9z6n3Oc8MSHxV6
PziVmRiQgllCrRX9rg7aBmSAHk2ZpUE3lSdrKROpeSjLjr0TWHabABFOe9yws0YjP8gbAz8MllyL
hhQstb/ltoSKiXa8n55GxfCvJH/gL5iaVxHmsH+h/uZoXF8pLnxk1PiTHWKuyrYjz7U5bC7BeTVP
Edi+6dmc/TiVVDaBgmRN1r/Wu5Vt46m9n64NbAzuhzN7+Nnt5Dsx2VOXRf7jFfm4XlP5Tfimca8U
HtSyDKQKilxFs18HWRH/j8i+VDUKIC946aW46fNMbfNtQPTAiwVXSC/VoxLk8WQRZjtTvuIf/m8i
Zr+h4Y0Pj4B/PHz8tfDIirmHXwiNHS5CbLwBoGuB3ndlI5n5NkeF2/9lo09csZ2cVIxBfLdlwGzF
Ok15QgVaVOMJPZOTKmrUr1Ax0UNfGExysdtc2cdbiqa3NBVVwxXLXQ/2Qjp8+tJegvcuSGeferW8
wKR8LMv3XGOinQ1E5zHICKWTgjnCOaBpDd0/9QjoMbtljAosBTodWBvIPBlAKcWsp9ok8hXaKHeI
ZEi8IlQGsIeuse0Cs6X25YpN3wkoM9Qr6nAopxYBqoLNc2cRk6wtLn5+EWxglZUrnjg2YL9zf/LY
j8cQCAG5rzbDyMEWL95jFeDCJKmcDt0tMfPoELzzI5ASdBZPjmLXHaQA32fXMZcsNfWT10oQXSg4
9jYfUhRNoAIvTkc09hxmuiX0WG9xAxDwyuKdpmyAWyRHb/2zNjQxk30jas19+3vasPW9OKMJ/Ly6
+VCjQwPqfxwFhM89nh+/59kXqznbHtSxQ5MWO/xqXuzehY1t6VCT/Pz92/koYonrkhN8G8oEuS9r
yKF1E0/7fvSU2/nYMWNv72hnOWXsqzPliDIfisNNt3F1eQFqaf5xZloNngq7UQj3KgJ9hKb5as36
gD+lk1ZvMTH1QpsP5xZ3iUeHAy3ckePwSmeEkHhmYHSRx8jkFDiBRAplkRMcIGLcvC/lBuoA8peH
QpS+/iYxnm+9TZMWCcCUrJbLIuHhcbDAf1W8+vYKfzMTL8ETvmzTRLfsjciaPoweaedQE3QCIPbM
E1/WuLs9YIO2nftQG3nUSVJtw3lvngSlJRqI4407IJYERnszX15Fk33rr8tnOn8P/iydy43MpYFJ
ow4/AJj03jGvxgVqbRvMcvqdJICV+E7YIDlR6yxlMRB+04Am5eY2Oo5RvAjWkBYl9uNfBFJQ18AB
uH/LZ8SmNHSOyZBzuTERahdZM9PxwujFIvLSI9gfKS6zK4LRa45AcDxugJEXHch7KCkWLHJGFMpu
xTOH6YjLvbKuP9eIsYXqIrR9E7YOybk/lvhUCSNrk3KXfov3HldEawOqv/bmcFv0kyvezqtsLepW
Jgub3F6GmgAUAN/W3HJzz6U+Tdd/kj2eKf98fMvicON7dK/VIMmQ2L6jaei37lyuLMvkfIvDUYlV
3eLEoPW/qlEJAQLTOb72Xrb/gTV3ETuP+57gDmqE2z91shEwMAWwNRI0qxf5bRPSM/dI0s761UEj
4CmyYKnsAKAMN0TNg49u+EHlnVKC/D2sigBvbces5yj8wm2yQ1B4mQc2In5oozYPpTyjz3UJg+TP
IiZT/dAgCFDLVjarz38iww456e/O2N+mn3sCaQ8rm6tt31P2nk40yubXhZUujO1dSQLopeWgOiBm
c4MysXUZ2SJN7SmDIsOeasDCC+5ASNJxPoh4sLAYK2FXq+NFHk+stZfFcsdpnigyRQvu406gomVW
WVjAT5ffeaVSQ5pi/Q1uGxGl9/1bmJXarnu2eGm4qAwzvRpFi8VRvUeLhJZxFm3qRPt/hK+IUmXR
xTO/b5ZshMC7qfVlyFAaiNuhOROoWyw4FPx4Ma7Ye9ijwI+Ougs5tkWlbi4VKypZLhvKqrhzu0hS
kmTdAtmxWfHEg4ReWougnNY1tvSIGQgnqLr3gasoF8m3f6DOCl7X0ZDDVoWUhb/pYixZod0CutO2
UODyxkXWqa15pTX8HLZ1WMcAhpwZIk78CaXdTlw9la8kgQSwazAC2zIcKmLPNSnPQo7eDFBzx5tj
H/RoMHfJ1z9QM7PmHvUcm/kcexSdSM1cHb8CGpGP/0F9n2Kh6yJvM+x/Rq6obFQmjBF/4Qr8WrVC
TWYD4S64xJiRhkkDadkDnmY7LtmAyJLSvG5JPmFxsHh+56hnNNT7aoNkK9Gbcg5OfuOYwRyI2muK
L6amjvGGXPNI3oUgIMVU6qWQJRprPxIC7fTfLHTwPTKYupgxt3zK3fuMLVkqdsweJ5SV/YGiw/62
hpArqoKQPOhE+ZX06VYUF5KRd3WdagneQ8T5BzT6uRzIbcugAghC1FGE3VEgwjH6I85Od7WHEvpm
MXxb5jefutbFeuzhFe8wuhv4snTIelfJR59dtvQg8Os/+2xI/WaFiU7oH2JSOmh078xPnldl7X41
GcGi3AFHzSqVRDMi74R062CQ/EHZWvclYwRdnIIYqQxrPU+hQQ/Yt/0UzZi5uO4HlkR7wpjnMEOI
7wbLmuBnv+bgcl+wXJT0kmy/BWLwov8hjkX4F0TpP7DsUzcsQdNo11qYStbydpPPk9zK+MGUX4k/
MndSwmKwwC5gv7bNswt0WtmlhsaR6vs21QcxCXfYv5ErF6kfxYqf60mTj3CSeQMZnbMUrMnOXWOw
2M71V+eXJ8dTRHeONOAIVp02KJ5gbRv+tQtlc1N1i28zjdFQWRl8fTTif5WYAKrDbv00PKhq3vvl
6E4VCCEuw+bh84T4xUXGU5O1wMzeTy12FZ1F0b5QpLj1WEp9pnvrBR9QbR7Bze086XWZt4GHC0UU
juKaJt0S4Jk67hAbLgW+ARQ5kTXhE5KKtX0e7BnW0hc8EmXlpnvr28FlZD8wjdwcTcBbAd5Fbz4f
hHNuprOBlIQr9v1cKAnputj9owaV94MVBlusk/mNaSHKLMyqLl/AnV+DxzvtYIlSmKrvWEXEIVWj
7Yw0DfREYtbilsT+dwMGgUqibSYT9fbyJmr1bT/3sy2gEDDCp/Y/K3H6g/8w707D3AH4BXBslSFf
BylGzI7jJZwdjwY9cRvdxMsKXAlFrXnbOARyP2rMgJJKst92GP2NcjlPutFMK6F0pSHuHtH/kahB
hnJNmR7NPNu7j9dCPJ0ZZ6pFDMYiWLhQv2BZAwK6stINH4ud/icq5k1kCvzbGFv1ApT5PB2ZyY2C
xVfdzL+hMyT+3FxxkbM+3mh+9sCMGAhj8e8NMUuuTdUOhTLxXgDv3BDmvDzCHeCdPg+gf+dcwFm7
1rzZSV+8+X5WT6Q3XhjarV0eDpf4CYoggFllfvtw1hjem80KAqNYP9V98eAeqomIEdSJg8EQD3wL
PQx6q2F3EcWhUobf/wjbi4vYLI0/b0e+FEUk5TcJpPgGWNeAAfuS+67wTU+/9J8/au74VJbbk7ww
I+BJj5vyWIpB9+h5Rq+tiTvhewv3zIrBS7xbYjsbDaUDghfbpp+fAt8y6gU5au2o64yhr0icKsZy
kbZENmzLPt/JedjVoiwqgT6HLqXfPAMluLqGzVj+wjjEi3Kg0YP7L07s1UWQ+JeDPTDWFSZjlYbz
VRI22P66bpCsW9/+k7kTgIePPC81WjjODUdyxsS7V4OpCoXKPGpmoeFn1Pmm2H+z0WNiBpfkHulE
QdVSVtTPHPXiihPY4jy3iJn6f5IebCZ2wDgPufMY1XAFFlrEHTZX/7i+uq8AMBjibDQ9EYCackD1
FuzwVsqYsdMUQG6XRXzbK9Mh4f9TdJCzakbiyY/BduG9Ko2gWL719iHGQeQf3AJ6oyIFI1ReaeEr
OvhdbgZv6bY3YVwPJ9CumXF/bi1bdbDAkPLE6S5m4n0CfHuJFJiYZGWBpIi7oJa973mhfJ9UQJvd
bXXSRkgorbM/xiFqADOSquMJqMeIUlBLijmxtmMOMtZxRWmlkLGosygRUDFdGvwGsnpwFN6oXWgi
Souzn1iZfE79uN7aURVd2MXwxP8HIwdESpl8o1Rkx/OxVp4NusOxueAU22pzuXRERZsedFxuMDCA
j6lQpOSHT7xltcuwrtvehurFPDjAJXO7x2uSzPkPvVYfPk5uFYFDLz8VZnXF+/5kcj+eIWGkdwof
tPU6lCSNnq4N7KTb3Ua7DBHMgW8NFxxXdTx7C1JXmAknQfT3/W65LEu3s8HnOMB6IbvoC/N9yuOh
LDX/ogeE3cyZpKtI1zRKHnwGYSO4bvoUq4uVfM7EcnDcZ8Ha7q9P4BGOjaNHRbGWqNucJtcOwySj
WVhRtOh2CfFLC3f6wFwpYWKcNx1zX/Nih+1fL4K5rsF3wyI7IzOAYXEz/bOHWY5eK3KdHJ7eZnvw
p9hA9aasmOcDe+e9yjVtj0LN5lw/zcIkvgQrBaknfkMOaoHRSyUYZhc8bAdzdSZSj2/Drzj0jaN7
2hwm7eRuL907U7oDwDmLXnZdaCQevy6VFhXWo2PsX2M8mLes/zvpPJncPc4lHSRVKE7FdxoMwey+
0wc1c29wYrsXK90WkkRfRm53vQqCNuF8S8QWaGZOH/ZyYyTG6EMtPctmnHJ4tnM0EwcxBFvIzVyX
iZAhllbgTcex+qxGEQ9kzayzuoSPFtm4dSLH0fjbVb8G3JsTVtehRT4W1j005NFkxQ1/sfhQ5H2T
Txlf7yyI9rCKGi860EF24TbgvIAF/NHv07q1Lob3/dk1LTG4Zossn5IOa1+y4azVfZR9NJrz1mtO
XTP8gwb1SENih3XtUXfwiDQ0Kro81KF59xL3pxpQC7G7mWDjTUCmWJJ1NCD9WFaiLTPEV9dDRMRm
S2HUq+xbc0qXvk7zgxuXzLJUDqzTVniA3P7A/MAvIsFYaCtCSPzCTnnjHVDQ/hwHrLQVzvRGTl3h
I3E7EEepMAGaUUmo98LNyAu/9Q5eM5KNzby4Dtnz34BUNNYOuQINbmSQQWiQv8foCFUmPCCx2VKk
J746JtDK/baaMh/6roIbJdqqdG9H54ykt+9eWfPj7SatJ3SrplSLM6kIZtIlZDQ6I2siIuJ5ER/z
dhX3JSKQzoXb+24fX2i6LiXKJ8aZiZNQiZAfJ0HKZ4i4ru8v8Z5c0ZcTaPT0zZgeWwXFm0qs744J
JDN/vN46OABDoqp8yXyXPwn6xTouuEi/rl5kSQTo+7R5sqppOUKeXjgVjdCgo9yPH6K0MgaxTUDb
unUNpfbg54ZzcfPS2BHaXu6b2He9Ra3/NYdmk5niuAsXNeMb+/+gvHdU0aTUQ/WtvnszwGivrQbj
ph8BK1c4U8124fEQh9CnlcYj8AmJMpx+8mIrecnceI0LKvizb99nC804HkyLlDcCx3BkZ2g3lUIo
myhumDtA/Cd++vkpWhOI8yagTT66lPFulTZvydkxVbYIMmEmlogOwQAw8ozGw/UzTfxbR9b/gO/Z
w15DhFhzhfYfOgHWW08ft6PRWQwoJQYqNtzu5hyoYLpFFyWNzKT+wnB+BscglAyuB16AcuDK0KOt
c+4c4ht3+eY4fiRYioyiBYoC3vH5AOKw28sNezQNg7jOeQjAFYd9Sn+uWac53caClHUfUzg8zVPr
POQxaVii7Bj3cAidJqPISt9PPj1+ag8IQ/1sb+k9aHYvpwOyWqHI/yqAETRfRDg+Itt8rCyucS6b
+NFB70grhxmV7/w92CeeLsZ6adxdtZp0arvaeJAQzHi0q/Ypn+reaLmXBoDU9xERF0PRQhKSXwQv
RGSG4oTqeqioJZhJs6sJEZyPVJVy+zFOQTz8lIxVCvIgCPrO/PqTkSuP4Lw7fHKU3CJdrYvGI811
CgUjvJvMayXppOo/Y+38zx0FU+KZke0tJ0ZpJYN30KBhiN9FFwcp2kaT8SYamDQjhNsXi4fFq1Xk
KtBgOdE3/KMWGKCYBnfavjQSfx4Q973Qem6oLN/SrgeiIO1kdnMJgbAgA+qlU9h25IxEqOiczfvT
cRciVgKJQE3n1+Ie6uR2tRsLC94K4dt0ZxsFxFzWD/rUzO2w3JFaJsNPPgqvvPTd3JT/HhMCrg5X
OwqvLf3wWaing+5JWIqk7ZpQj+r3xBKr/qOlbyOFjnrhqgjQtDv++IHymN4UJLV/E8IZPwE8ZYGV
RiBPAn+Zz0f/2NSCs2YlMZIkguP21+zjlsEUtEt0jhpUqa/y4Ouu1DKf0jh+STwyq7qbw7CSxgI0
S8s07jNZsIoZsANQTUvOJFEmrJ2IcWywsl2qL+sv2lKYYNDQ0COGWN+bMREP/VY5QhqMKgy5eOPG
/D5/Q1hq8N16CrHQbwyAI0K/w46gVcFJSp7neI+LXwivlsUFzw0VzvHi7y83H1DgCKWeGlDi4rDP
yHCJjbkm8EbFMhqJtYXjOQRDNRji76CWAX8e1fhol0HQtKP9ifIriskezDkYGCOELcdGpYO4bogO
H78sWU0kYTWRSegDMjVc3Ev+jmHPCTlgStZ09MFVmI/3+oADX9jSROLxBhJFfJmemaDw2GUKyHq0
uZOtwyBeEG3YNl5CPu5dl3Q5lukzfQ21fULCXou8JYpMSoD7M8uV3pCXIXlrVePS/7BZce72Sv1a
yrGAylH46MYFg0UX9cVicZFVRkv7S3F6Gs0mZhNlOIhhuaEKxjSRg5TR1IY4IdAWVEIwhgfqktZy
cbnbQB1XbMIZOLHmte/qicIQesNXs00exLRFOCX1Ujg1hLlYLHnot5tx00j9ywkngwbq+RGWdK9v
iKeHDQ9g+NopjKfcKuMEJPhKUThY+CstitmmuwFDNlM+rixNMURaiw+IFHx9GhSSBME0hcpvIq7R
Xzkg31Gch6V7MOg02fa6mS11fHtdoO84tdV+i/HZFLkCiVqXUWnBag8/52SlcFRZMoEitv6Ya5a0
Qpd6jUGXRGKAz8wqDE6cwpp9pxFJtwZDxbciURFP3bmVdXBFewHgbhJoyIErL/nBlII+lbB1g06i
y09Ub1WW9Ps60sKhx0BpjM5pCtPd9/mqrzB6Pa6D/oPhaWJ/E1qaiEcEtwgHX1WpFqJxCHbd4sxl
CjvRcjaeIa1qL/6zLmM6dDmSAVIs7/qkhAaHMqVoSf8zonJJr2zXi0/tsf3eb3KoJ1LxGcAJGWFA
jRgN/CKKvfldmMlht3/3JmEkgqBH23pvV/fdvkAASD4hOAsA0sXic8KfqPfLgg7FBiLM8hHbrU/t
t02VR7eLT/T1sJ8TTj++X7tlWm46MYdWyyEzUB4lf15qYW2LAE5qobeExk4rWlvmCQ8DSz16QJQb
IZpNycMCrQdXQ5werSSdi4mdt7fhDi2Vxuc0jP/V7lnEW6xfNua6zW3cgjvUoezwUX0MXjfDBFMe
S7Qj54MVvKqEX6JT5dxIQ93GQU5wUJQOQzIjH3UPQClATDAkYtkpFaP80Pzsq12CbTSJdcCYWlaX
JzcM8iKNm6AkCNwapWEggqgshzCG1uI9x5FY+prExM5YKi4pKOZSln3DC5CG0Gfy+E5qN9g8NXaD
P6CJpxH6NNFyqnH+9aGMNJm1BLITzQ088emiylaQBXhaX1mbFXC2G+Jsq5d7W89dtL2xxo8ZSWfr
COeeOm2KmJ2IQUagjvdUHL4j5frYOUEt5XIpS+a6tl48BQJyaM+eitU4wc2rCbn6ZloK4Fsv16gM
hBaQgLuyC+sU1yn0jmtJgG0sAvDShjFI1pKNceGUGEW2U1nOqz9na0JktbbZse3lM5DbDHpfyj4o
NxxGQfUUxy6HZR4Gk6RynKJgA6oYTygCg9Y/Qnufhsd/jVot1WuYc1eK2fEYsMDFN0wUhn3gMaDK
MauILUZcwHliclBGWh/d0kXOFkh6iW0hta0824tPDZqXXwuXMKfKHzwvvzDUrLf0HNsT9FRAFxGR
dXbjnrnG5rwmP1rDmNGF7xs0qxob6jxGDxUcsj+gN5yoeCwBmDMbjXBe9X7agiyP1OPJ7pKFlj8q
3ZKzT9chUqdAEfioyAJeaaLw+SNJ+kRlpLvW5BscSwXkkUuZfqjHXk2tLI0LoI6wFQ6jULhslEnJ
Jc0Hixs7I75KAHN8GEitRJ6zQTDvcqf4bQWWFeUxzk6zWXiZa/51IHgwKHhmF2W7F3jsMF2c6qU4
FDeAG58Ay3WIfeY+2nzw2J43iprt63gH6BmsiiVYEbBspvEx7gyzqtkH5ejB96yzmGgQBPKc8ZcD
K9YgJzRG5V5tgOZaFTxtekhKXiuKOfjP5nExXzodkMLzT5G4SfGjzxw4QnWQwE2+cCMkF2WdPyj3
lEuKV61dZ4fGbsXJoW6dUM4HV2sCZipzjvqQW1PrDsCV6cTFPoYYl/e5Z96tH+WgtlPMdATFk+rs
bfBg/uXLdZTbEMWtXFmhoIS9zM2RFet1zEyYFOzBZ56CiBURqOXSrEhqzXOvXECxUNUxTBqlefu2
4OQsee9mmDlmFYGROtGAC7V2ahNYpeKtNY58a3+naFFEfIoEEEV0tIv3M1yIxN5yMIZLFu3vJu9g
P6Bi3ph7R6Yjm0/Ev83LaT1RDkJSGOSPu8uWC9tTtSHRzipJ+3aeWTqKNxTh2xpqzL3ty8k+R3oA
vs5VLFYjH9rnkpvkwIGMT8jHati5zXpB+6TZzrJkph/dx3HzcX8/CBm1qJCrLkCRTTCTZDO8YZ4a
cI4UTw2lb6V9Xb2orn/HBCSOOC549OOENcaNXDhsFzoqPfp6qZKKin36Z6Xh6o8QU6vxLkxkEK58
O05cOGzRXXkX3yGxa14FR/+yJOg40dMMxq8HySU5wvctj2D2qnSVXeNO253bOsOcKcZ9FM5YSPRQ
lmc3eWti3n4wgWPJkzcNtyfS9iGNFc3MfuKyTq7fL9vQ7cMB8amaNTToX7PAT2xRrZmeNuq4c31O
WcvyI/tLk2JZYVTR8MhwcmS4KugUwcN5lEuEUaYrLM+Td1iANDNlhcGe2RHjbM2s/3OWXHe+m4Qx
xmxNMTyPwv+9djph4y3W7KKi+b/piz3itNkOkSl3rMva+V6l2yx/5tKk7XXJIXbGUO8pXy07oy3Q
cVnOsh4JGGpGH248Yh4Fy0VRMoYEUO6hqCUar0p45DaLOyK0a++EFx0sLpXThfhP6/A0L2vO1Vzm
EG+rj3LrdeJ4tzkIawBe8lOKfoYHWjs4kkMB/sBK8/RMvGqowlawuZDcEiZ/FdCgCazbmIIGYFfA
zLncqxNb93QqTS9WU1ZUSwOGlTSDv1AzIiH/7tKkMOOgB7OmLQRzyUJjRoiksD2yudqtIom/nKIb
4/gn3sHYfeJFQHxyj8dXYVU7PGnOPyLJOMzWqDgMjz6zTf4k9rV2qjmZUmEqBRG/4qE5qS0q/xxF
2fXjxu3d7Zi2KdmZ8Me8nWHsSiPr6TzuquCkTOgaySYvAfLM/ue1oPAcwJ7VHExSUWJTEtlH0NHh
HAVZ8gAmuQ810nJGd3y3oKwbmAqvGGQIGN5sN0tgW6Yh4CaJEEVE01dqN44Xqe3iybHgk6TwjmW1
AUZBelCU1QhH1hjGedig9e4f7lblbLObutu6K7mdGd41koaU4PWymtQWqlNl0U/O3Mc8xKrK96j/
ZCYb0cibLXEREssucH2aNqOs3YMStS6ZzRv4AJpM4fE6y9C33Yx65eIO25xBtzklit2plSqzR/qO
kYf2v61pDCXmG5VRBxIL7IT60GqWSF/M3JMyvuNuOkRiuVTKHEeeCy3b8GokDJ0L+DgYKItYeoxp
0veuQVmRrfMTqkuhS4FagCBWMwNNwGr1PtLgjZf/A1ov3R0h7PSMJv+zCgChMxB1y/BfjqKBUi33
i4dy/sxcGXpTkpBKrFq5LbHUnunZvaXucQ4tLJDCbxJF9tDsP+7RRtDFSS8yAOeHvCCA862/xy9I
9v+uZk1hFGOqpiSg79KdlWYncZQt8MXMJrhIlnaVhU7UeRfG+sYKHovpJEeS7lr9RgUOQBEB+LZO
9vXJtBuyNOS6j1/R3G11lLuI9mbODso3rZE+nwrM9vQUpS5/0MG5gCLupG0CHx3lLgcMfcC9cFIS
d1ET0RqQGBTCgXGUyNqupD6MuQA1A+XhBCDWwIhdtt2jBd1HmbykK+7T5xfVilLsf9NU4J0kcIZ9
LahSgkg3PqY/DvKkhl0zAKb8hFzavY+1XAaFHsWpkI7J6yNidma02XQXonkaZhdL8hDW7G5TZHUJ
FJ+z0V++YPOtbS1itc+AORo9aG+xGWuFk3YhLhJ7OGx+RV2r1xxNgKJqdY/sR4fhlPh1Vn13v5rv
OWfhZP9DreFmd7pyFCA1gP5lmb/8CGTya24jJh7D2hMB2DcbFDjEdK0hNQWtNsqqOFd/20N+ULiM
MwSkJzvJumu7ieLoq0cf0LHkgYmTdd4yve/YGd0cekriNJkrV1ysBx6dnhMCyq+12uyww4IvjvyX
NQpo52wfRhOc/HWlIC7BPLfmmUahXnuQMEMdus1h57m72L6SOcglvPk/g4U2YTHEFltFP/OwL0Xq
xCpmV7StJpQ1XY+6pdD1QdPrAXz2k8Z8ktqCZT5PWMntVYlLM0uPbUuJjNmiAeylBGJ0cKo2McxX
NOeSXnBe1MfmEn7IyCtF+1BX2EBA0y5TdddNBdfH1Xu3CQ8S96KL75Kt13hYPtq8rAuYqRC3GLvd
CtPAg6fl0gf9pHevVoYMG+lC/PC4bo7IOXCZq+K2YFUgi7Xu2+wUPCBpbNMS6fWdywKlmlG3dpCB
Jk4DKsjfmf7ci0hM8KQoHwU+Onf3ZxqAJOrUdHgtA1LVQy2Lfb+M76CJ6sNfhajEqyiB1FzH92Gh
FgAUbJjqENoP4mYntBZNfoiTCZOafMwC0lymfOsQeF5yI9+j8VUluSFLpm3Zn97a7fIXzHP05GcZ
RHIZj3m2BPpCGQr+R2qSGlQsrJgp2i3Q6dR76+lPH/iwt3xAgW+9Z0kexbCKsOXenjiDsBL+wddr
KzCRz+VHKGKPSuDllhzvoPDEsG704dGuSKK1bpKJfwji9OWuEC8YPtJfupqpDF5lAobQ19Q814gP
pVVzHX0et9sRKdkYfMJs0s+Wq1zlfTcubVSlxgnPFyKGMDahb123O0Wx5NUm5hOnTYQMj/9lUorp
FtcdXwPlgESYBz6n+0wGEFWxtWkV/hN1CL/IR+7reNiFHKnCzzlWTnB2rZp2/ALjuDBHvNTwQax8
3qGyh7vA+uF/ZUq9frUCS0iCpg/Mz9Ksn84CCG9VAY2U7MQjA6FC+hGn1NwyW42vq7ax4TwaF8jw
7wUkX2xT1unqrFoWfWADD2BT4HBWygLAMURxKVa2r7MgAn/MJUpZ7ooCdWaQyyBcqiKRPokKi5rU
MjCbbM1lO5Yy06r3lPltyp2jI1PpPP7ymgT6rF6pFrFsLqEY8+y2eEAPl6jRHBWMZPSWDhI0rtEL
v4okm2IGlxDpJCfYCARQLv5zA2+IQ1bW/SoQ+3CHxIZ3aO/IMx8Bz6AP+s40m0P7uML1Gmplwcye
eZWz/y6hAR01es1eYjUMRmXaQec8wFPqCIV3pcjVLF0kRkAG6lBe8Bv9ivf8Lxx1Sysx0jHzmnmt
4xZNaKZFrGLrsXTYOCAWz8eZ+MZi865yCqayStEyrRb9I8nHwormjtAk0Shv1ds1VLm9mME5pjrG
CQVEPz1VRKYHfXfb8w/H5SqKl35Vdua2KJTyG/y2A/wWc0FaWiHoRDhTHajYRODPCbpQVvymBNSS
Gnuwv/Bp8jNlZpP6JUW8Cn8kAuMk5N9+TmTaYfXy+IJEcyAg/0KrQkK3VY70+p/HRKb+VlN3swF+
2MOvwHP+ERAK6ibFU0p6KzNBx2WORhRe6yNjs9Nvd5gA4cavywN8mUhr6qWdrFYqw9yqNJ+uucya
/FoDJsYJiEU84EJ/wkActlPMsYy/SKIh6vW+LniKC82pP2dBBFYzi1+4m6CDR1AWqialx+KHfUm0
PfL9OQvchZO758MtC9R/ozI7W9S5KiupN9YNrPmoLfqUFAhxYoIY3Qcx9Z4rJwWXZ/2GY6g5/Q8o
J1bzLoDz4RAfadMbvD4yexEQyYyNO5Zdh7WDAMDvc9Zt7nEa2QU9SuBi1s7PmWReMR5aYdMrdljP
b7Ebf3h/azX8E9Z7c49FcsQL5953gZRpv2G6ioOkZydavgebNCgim65k+RO5634qJdPLcmuRLyAC
JUwFDuYMzAxDpozSXQOkfh+nwOH92b7lvFsYLARR8/wrK4ijM/vuTYoTvmKaTkUA/4p6AdCoKNjj
zUrByyiomud+y5NMcLGl2L75RhTGNB58xHVmDM9dJNqQROeN1bfUq10W0pGvyor76stWXjlJOLkv
+ZAHmkgB/qW69n2dDdaYNDWjHuYvL9e99WZaYdEO/lVUQ3J/OEcNhsg42WrIz+qFjkZQs4mE6UAO
EzbLgjUCr0XTIjx59Wlof/EjEMnW7oChuUelL05q0Jlh9s/PmOkp/OTpFTB+g5tB6G5yFL0t3utS
ENsLzDNRtwPnp3/GY/FlAtznFtTBz/ayOryyy29Zi4YvjFwxlNiLCzQcXop30jE9MTtjktKg0P5w
8EUUyIvSZY00Pz080VUyeIDnfLxutw5bXLdzeBY1MhGgLMugsSwL0kRl8R9TpiqOLCdQ85IPCuIL
isrjk8QIlMqvCDJyx97cuuUu05SwMbt5sWuzC2PkhSO9wrv4oQZq59Gh3KBCVrlbTkD4d4shtQ4n
AP9z81HzmJOmBvLuOxtCL16gwsOotNwpK6NESaneoywD8pvdahkgT/PeqApHf1KwfIi+ZEb9Xe9y
y2rtFoXrALSv9lZcoQ2f6l+Vhlcs9OqRbpGuuRePm+iV+G+wpTZj6KgBfTYJYsaB7ajDPeq5QLxD
CAWkm1hfA0uV3E0BIAusxHInwFliTWH/GT8Imd83bWpT2YlxK3qZk67Mj0mu6683nFRgyZsjnDVY
DAP7F8nwDAN9JCE4T+kZsmSky4y3OM0QCQO1FH7t2Z/GwkpybuPH1KBM++b6Pr1Yq7belvQiOPhj
Ce9z7Fd/sMt65NkfPfDC0w1lT5WSUXU9dMbXLYWNAcY8STlF6pzXKPznn8VI6pmQ7+teta/CAhZP
/lhJRdHOlxpd0sHjRrqNCvqANTx2duGVxoVK6UXyLF+Nb74VOC5wiE8OFn1XiKlNy5MGIlvUTIuY
yTCFHDdDr29YZJrJsQhBD1oDC6DvPwzskaSP40mZMMyPylZsy+gWXAf7s2zkVNsqX/J13cu1NQke
mH8QpFFPFMGyYSZSo8QBwzUeP62EI4u6BlGtMNdkUdrBV0mZpATsPyZZSOVu25ZYjjt8Fd8Fh2PO
tkEwI5HVkKFb77QPksYifV1mp/k5JaBDLn0UgFfckJFU3kPdMkJ7e7nIlV3Odu7m7WMulgjGhSb6
zf8yHGbhNHFotaBHSqV0MBGHvs3OrSyPHtVVkNgKsrGep+hKHMG2PHDBOnGdj1EY3FVyvf2UwNEG
cMsxtggv6Nf3Nng5eGV46y69OziBQlQbILkwW2SWyY2uGGO32lSgEMhHoAb2Jx30YptsaJhSTVFh
4dYKMzp2TJaX8M51QJah6sQULet3rgKmMpUGT3/U0OkwjIu4T4vCPaxslGgJEVWYrVMZiWnsXAcA
eFN75QJ86n8JNoB7/pwZ8DHW1+L6tDt7CsK1R1CnIHTIHXSi8e925h7QQwGP3iz6IV4taoK6fEj5
OtZ6a2yp9JzUCRgBBuS3JZfysXyuzCuEhSZavu5I8/QwmQwNBIaaqPuPNinfrg9bciyaExxctOFV
rHHVIKfRWZ4OqDhphsyKPwseU+OGImVqOScBu+p/1Kiu4ezsW0ER5t2xXoznH928atwTZRNhWxMB
joENY+DUz1IeDGlvYy5n2t4N+qKQbO4UV35045j9y/+LdNR9UaoLyLPvKLoSie7yIxG8jbY1XM/V
+3xoy0ECre54pljfZgp7lh052fUeatl2Q5qbfH0Xe9jMFjgp1fCHH189yBsMKI0XZnEJ8gVz3l5l
phtF1HeLP5l0z8Qou/99hXX1KKbhdUjyI6GoQPTub+j/Vk1XOe7uHQoMIQ7TEBELvLGm4BlOgVHh
TjrSqeEWhP1WKqHOijyC7q4bblAkdZUv3kYAv23GGXXZjxgEBI1BhCnsvKTN5JvGpXWp+WuXDB33
gZLPB8zsMOD9jTGj0tICETfIDTN1LhfQ6GFf0YxThhNJmzFe7+EM8vyKoD20tAb8MZtvnaTkFCHL
enRpHqPGJdzoMcTH3HF3oTeIUDjRniXDrMfheXLgqUofbITm6X7dzkou6IGLThxAaHWU1CM6Wv7J
tnepqb+7Ffp8cLyH+pkc5Rs+DJP5T6ZJ/3Rr5CY7fVQKOjA0xKai+D6wj7nzktISldNEzv3jnSlE
9bGK7G1T13VxHeP5XNlrW+qTmPyW7twz4Zom0StSVX/ag0NtYOYuWIzBFddvyT04l1cBbXR62RBS
twxTgSMTmkzlFKzCI0ey2WXY64jHiw2UFaSrWLaSbcTEdMxguGRwjhGhQe28uDrXEGuMpn2rZEQW
d8g4a9sLIbhPWSfT/JwXq2nb8nYmNJ4FVcLEpfhg2FP82dm6vDZhyAcOi1tDho2Jmuab/hzBOBwa
Z+drhf5ogX5BQhmFqTDVkyYbkf/1eb9vfoMUdYTOym4ekSXX0Dc0yWRRQRc/pRiXT7spmP60SnCZ
Y7/2/VS9a8aUovfwp6nxl+6H2tJLDWK9sYHAbqa6Yvr5NsbtgtGsuuEl2SB6E6FubxBmi+S2D1eD
9PokFNIgi2kZYyq/vs83hiboenGsrMQWX/gbO4RbYRnM0HaMoBORj2YTfBaWR4wgPAWLVjLtdiTE
RuJnWhu9qXUEOP7l+we0+HjdSNlZN81TgJBOLXRuzZYBqy4jVhC61Hk5JPsOxPjJklJmGsmzm+O7
IhRUuJP5FC8xRJLCo4ZNRrSVIPlpHevMLz5q8jqphR/4REWzAZfwRWW0mHmB+3CFL5L+phRThHOz
k9zLAuhhDzXo+TgRiCEsTOUdPCOvvm0vZShzTubq0O+SrvLMdbyKmkmjG85EigX5RYGkURkMhTml
Kp870vHTSFjWpluQ+Rf/ygw374l09oHF/pFi4oKTgkw2JsZoaJiAKAiknOk3A7Y5Z7dJ9kR5Uyvh
lYRT/04QKUVTjsXLYdhtYycf9j6NCGQcTvbgFDa8pX5V+Qq2wgTkPxE6kAcqDH7HDnEjQNf6aMOe
qHlHY/I9o2DHqGta3BHSl2ZuDa1wOgVcZJf/kustO7a9yCqRi8X+84q40a362Vg6+1Jqe4T3lfTp
o96mZ9JCTHgvlu0xTMgHWR1hpR7T4QOSRBpgekeXepBa9wUf2lNV+I//1AwK/iEy2r1Y7n3MSKEo
0VWeKTmmR3vdmXUfyBSOtxx5stMpOzoljm95GuEaoHFw+vmip+1tm2Sl33Q6xQDQ7MV0ZTKkrkP4
0Zp5g9PO8XQVfBz6xnyAHZjc32VykXqrRQ3V8zw31+S7zInT61Yr+jGjX9EALZphjBtnttIlvNm7
C6Cmn86cd+pfp0ZS5G998LOidA6e1WQo8rUsCUgrQUXwXvubKqCrrmUOqWguTjaeCcYturd3fY7B
menyvBra4HOKPb2vz53rrPJSWTconmqDrTK4zWHo0LhyePcAVA+bH2SfPEwub5otghDkWjYoq99K
PBkfLO9+s6TsRIyj3ACEsuMjwUn5LKsxGnbb3Jvqx5NnoOMci2FJsSM7xhPmeOVmPO6QC23kaaYf
TGsJ9P24b9mpjtsWSMV8ZtvsuQw8SgKp7grOWY+neLLtVTkgBy2osNEPj19fDYR0Q+buc7xndLIy
ILbXC57LDm+iC9NYXjyNz3oZp9gWsrnf6aVdlV29818cMlqwYCWREq2OP+5mGb6a9Ikha/xPKFtd
SmUmixSmNNcWB7I+vq0+mCIgWOhwwwp5bAA6ZEYry2J4oDyhiRZG573A+p1JjF/bkb77bBmqF3gs
qIctQEIVFQYtkofxtsxM/OD7pezRepNsp1/ShqADRotfirOngZLi21EI12qAK1BetpjZ9g+RhZrX
ZQIZsLKyPlPliErl1/rCD9+ZrywIu15b5JSHk4xusEMP71lJzLkc4oXYk6tkgetmzhxUFVPpzD0M
VZjJMveZPV4CPZ5KLcsVaObHTEYP6xcShVR/oa23KVrs26AIciQ3Ss6lq54jO0aSzye6DU+QGLx+
k26kJFIONs81RmVzykNvZDHv6nbIxsfflnvv/PWRzfefEW22tufAN3GjPTgCY8BAhNOu5AXJYPMZ
nFPJzdBkbKSndBaV9IDRnQ8K9iQPST3EG/U+ObVfF2A1SFV6oRF9aUTSyNuk3qnuOxeyvx4Pxv10
58ZrBJ3q7GbaN/VrLcZ2E9ugpFYjcXGucph+J7vaHmWYeg0fd3DNGaDNKEoPMlM9wL76qxmkqwst
NDcF3pCaxDCmLA57mJn4w7cte+I7kOUCi6tRTBiKNiVs7wDkP6YCeBlnzQ+Zqu4FjkN1hU7oUtmq
bxQjTHnx5Tcyq0EDUqounUgn/hYssAzDJlKRatFuvT7QUjYmUJNpIHUEE65/rBeK4ubkYTnK45rZ
50S/OqcKeA4OCIdT+Ptb+WmBiZ350xQussWORuHa66HXZHtGLz3fgF9oxRNVeVx3rDuH/aa6JbpT
rTR4+Ds77EaqnZdc6noH1O/HYPR0rVDOHDvL5H7oB4HZrWsPW7HcD/yugVy7Pf0P99WVN7r8dDiZ
lC0+USMJY4MDtUtMqc1/XBdaXoAm97PR2xQPWPc3UcCG/2lStK/AqGEySRkuT1rAC5hrNVTavq//
XQsbvbQ8ZBUDxRfzk0xABbZ3nloWYUsbcEOj9m4JPV5VRyq3Dcc6nfIz59SUMP4H28f7wNO4iQiF
ViTTSkXGBpNAJNM7VNy+AZO8L8L0PTC2GFAZ9c8ElETjpffCm7m74IYigy6bMTZNh86ZCdss1ecW
Zou5NshwIl+24bmjjtL10OAgvh/Lc5yd0YyNNINrFOMBmdLYB60jDSSOLEXtJbH1uU+hdjNk6Rl3
AYRGa+zVyv+x90595BFs3IO658ywy9PBTrrDHaarD5vWKOtgLRYyFlfOiNGwktW1TJDpSBMcCa33
O+e//4ETq2fP+FRHqzEidN3wCufNNlayJfJb1i9cuGgFj2FDe5QxfO5Zk6dR3owrLhQlN+06rx/T
wDbSOLdsidHyvzVMgXigIYY6HIUZxNXAGzln6hvF0dK6ycc5VRLTuPFKLrGkK1Brsdgwe2VIdBS7
A45zAqp/rsLdwThWM1N4EsgqPFsFtMIil/JGtiiB0riTKmd/sytjwrkNj1B3zAwlHBZuOSCpXutr
W0EoVqYugHMmFulG4Nzlrj0cSoD3vY+P2LkvaQ5uXcVE4OlKigxzy7+ZvHIVz1A63jMmRgD6KzIj
BO5LIifVhncxNcqDli1lBRMvhehYilxbZELuyUeI/3JxT52VkqYiN/lcMHn0ZaP3pBiN8DoQoIS1
RYeGlEFwrN6WHDi6Y3LQlepGGpo0hYpI12kT+pOH56mpdI2dVChcFYuwrBHhh5jkcSUwLd3C7icP
rrbm1y1GwI2xniypLpoKE14/an+8VYkTfYeDAOaTGCcQS38yIXFAUW6sva2kk545nRBIABxdGG85
JFr61XsIrl8gyAx6wKqz0OE4YwhfFr61/tyePDnFm448kILqic40CzxOuhy12MTiRyA5jmA8CPD4
0AxDALsbZGlot/gDNwu44o41GReRBEtVlTgYc2DHr5AuXYLHIyavHbgZFhk6A5U/0zDQG05IIzSv
j9HWq7CFhhJjHgVGagZbq7TwhtpSB12JxQTzATixnpCsTw6BmGj74SWszxNoOd1XJtUVXfAgHTLM
5GfLnzz3dIFZheukUC03RpwmjqZhtGc1zhDFYhDJntc6NsDm0B/UDHu3jRmZNuYg3EWEjSb4yqDz
iNhcj5jq+k+suxWgEglVk3WGURq6qqs+M1V+l4VXdY45w4xQmgwOynENc6W04ttWkesmgWsRi6U0
IFs9Hq6sbs9VDOcrX/HlmG552fpOCjIUZdcOn0JGeMEjDnv9D4zkLo6TN4UeHls+M9Y3Z3CZpGIq
6VU6/RbcX79iT3KDHlyx/s2vMow9oFHhgXcs/2mRVwVLzNlRfII2Enyvw64YTKCqHMAKVb5cy47R
tMd+CmK/mGDkcCghgBxTRCy6NSt0lf+UfNVRyzUhkSwWJfVs2TkVifB0sChE79NjFgcQswgwJfDt
2S4BJv6ZZmaMjJRxPrwFSHypm+u2Rw9cdUCufUkQHo/tWDJgrKPGY3VVsF72vpp1s5JsZMp3PKaB
veAWpUcviSbG+Tj4QZLeQo5+E8BZBqgMMO0Jk9tmezflfPzQdtvteQGyjTpmnhHkeOCbqrnhYpmq
w/EEQMqxG5XCzhTi0VD/QEqgUKli2L3ur5YV4mfBWuS4P4I8B78g3cVwqgNv33uVq+AhkIYmDJdB
yoAv+1rofrX5IPciOJXibYQDL0iVZDIKXnTYzR869PzhmqwjkrF4MJtv8K/CFifPw20q5tK7jUaS
O/uaV3nP62HvSKQi80Qg8i+xbKOaOcU9rDeE9gAig4VARFLj8I/WB3uu9O//YW6GPysRemu5F5Gb
xSDaBRmDXDbmv7/ZiMGjWbtYB20OmzgXU7OrfVbs6n97Jds92633L66kTE3W8XB6IliL1Dti1NYx
aBId+4RBQpxsLMfEtswdcot+ZE9fK/s/s4xbVYRNHE/NSl4f2R+JxXvm0DKbfPFOilYgZCtAxrsU
HIOroKcoom+s+yF9b/nuBACbWc7v8Udj78v8xVAMq5ddwnsTcKT9nM1ZIstkSSPdfr400CNfDSOW
/gDfeOdM9bO4wn4cAiSKTTcpPyn4LZATYj36HDmLz2f5S4FZKYj5jNtUa2c1ILjE28nS8kfotv4J
cnExSvQsAYEPfysBUpoUzh2bv9lZ0G2N/C5H2kEGqH3GviLy07P5J7JAO/6xh3CHPQknc/brtbRO
FYCJcQtTP8ix627srhn7HaQk6KbuvTtmNLLfmpkX2I2xmGnEffrDZEgVMsD2701ghs9G1PBlml7v
DJtci0tJL/IZphgdGBfqI22IHTOCUQYo9ram2hdMSo7vO278uyQpgdPVwU1uSKJdo+5MjhU156OT
Mcu67Z2d0ovVAxYfjv/heQ3WxiJVE+DVH85+a93QuMxyx8XIhck/7fTzfKrj+iPXt3j5Pu3LMfiu
lDiEyl0uLLRPSOX1O9cpVmRfHrai6aaXqF2NlzYlzeksFqVIZpWxVZqxSBJZ5YalovvaY+LItdYA
+fNExgY0sRphQXpDZKlgB2rmJqLqzbBkPJxQ/SxXFk5Wrc4yQgygNNOI/uSKP6NkutAyhE/d0gsS
ftkcZx/P9Ptb+CaU4+FfmJglFZVzY/j4z285wXMTW6CCwW89wpuKPWCgziHXnYOVYuKpuX+ifi3n
lD9y5QcTn6U2CTDIz86BreKNarG2KYHO2BcqmA6sEOy1ofJq25sJvYxeueTQgAY1MkRPS/Oi/Oy9
c/D6KduHFZI8e7d7tVmdfFbr+uz8V/ELPW0F36BkSTFkJr5mNGbuz3p1fo4puN5OZr4mr65egU8k
HY17gtYf8hYa2Wi/cYYPIp4GYK8ykPBD7MXoRZMN3hcOwft2/eYaZiJD6L04HkbxXMiIji4V0ZIj
DY9WbNGG/1Cd0Feq1ulGnsD4etviHbUe4R3Yt6iNMCZ8x9bpMcpiafMUKNpHiINthTp7ya+2jUCg
+gmxnSbrMem1erinL2VmIzfxKpiv1d/EzQrcMVniaWnSlv5Qy3K2welLwnwbo3S9NnujiiTuLbJd
W8Q71bb4Sg7fVSjCCFZ+3mGMBn4aIxq/XMRcyshfzzQqYykof5t3y3savhLARw7pn3XScuQFMkgB
Wfo7brLpzIckubaPKTKpp7ZPCrKj94JXFwc5MOg4zVwr6IljG67Iw3LSohEoufQVtkA0eeenfYtC
IC7rBjCzsOqrIJC45xMC98jw2dxsjjcQCd/UdA7zfmDIAwVXzc8OLlKC083LecmKbB+ti3npFice
xbppxMWnoIKuuFLBnY1d7dnTh4nkqrTtR6P473lqgc0p1duSL+yA5SDF0WpltvrFacEcY9/svcbq
PLouXf9wmRywhYOTDAWxo3s5nqGTrDU8V+oSSKSf7VC2dcyes1ijKSJPd2xmdCZn5i/SpdDm5XFy
U7Pli7nhll8k6Yr6S4LmZS68d6DoIn3SwW1gbDZtG/G1LhJ+ngUMigpOsbiJ/onExfsu3/vO4XHU
o00idmE5AEoFZvsA1x5AJaEi4G9CkrkJGER06k4Q9XiMCVL/3QimtAfcFfgX6mB6udsy7CvuyNOd
yuyI7U9vWGbaLczTQvuG6Nf+BNkFNsZueUmCOf2arerYEXOQhB2rUXx0exH2bcoDSRBn53zqwGgp
5LHJAvAuWo4MIycXp3wUpHbGVNxBygqYDTvh3kSG9Ibr8hQ9UaNMDdx497WUDuyieN9YaQQm3yTy
BXvalKfoKf6L0bjCgoqy1Tvh7PdXXB4B/0u+bVAjXd2HTvCwp7eGDy/fBEctQnShTXzMfv/yJpmv
BvHU/7NagPj+ju/IGs6T9oyuhxuF1uoWSL/6jZdMpdEUYYHctL9xBZlC1zxZ5plKH0rtqvyR0saG
xdF67icPAY4A4HDKzfM3Pk4T2crtnVmDbUD8C7GFXe/ifltXhrjg6zkBRZx6GCZalqbkK4uLAjf5
H5zj7hBYNM873oGpX5OFA0aG86DP6+6a7EaSCAiOoSSRuJ0v3IWz9troh+Yn4e8yMw8yHV/ryxZg
155GelDYAwQqP/Tw0ceVzUDzCQ1rr7x86X5OkamTRlLANQSjH0oHfMdk4DaLGYmDHOER5oS7gG2T
pZGg640aT4KtNeMcW5VhWYsYcbOUsIL4FeNwLdR7/NJy9yn0RRccBkRqTF8Np5B0NKeXOQrpYKF8
o6//VXpet48jPIchu09IK9ol0fhKQ7M5QH93tsNliz74JnVy5wjMc7DtuVm8XuwaUE7cQAGQVvna
w+j1iVm/X2Tsn5Sf6LkEytsPvbnU5Zqzi4AeitTOnmEaGdbDcWneag1WIJj3wDg0XVUx2LqmPAN1
iFPSZM2g3PjOSduABP+EerbSJ2heoKEP+Ckuz+zcaY88o+nNyOkuH9IJKDrP2rclo5qbGBt2p/RK
KaN2MTXUtZofDxVUxOCdwGwNtZvnJG2ubadmmGinjZsmM8Z2YZTGKnGVjEiFymR9Fx4J840H674F
ZH6Dp18L04zuPOSGAy90cRJf9As7XM9mANyO08viGKokZmOZzG3ePjq/QOj7qBCec/8kE42Yc5Zy
wT1ZnkyFA4fcfBxNds6I78n5NlkGeK/06yURuA16OIsGGVT22Fzqj+vkRuAWWNvk6q5e6ACK86IG
uj3Y9ztzaX7eYtWB7c/rqq/VZtMklJlBg/X2Y4EfnTTkg3Y5bhMUXKBg4S43kPdRriNvXg0Ujxhh
KfL56yaYQQ88fl0fC+rAKYEtLqFw+LGQuliPED2OAIz6JPTPIxgaMdlQquRur8bmFB3CebhwXZbq
HPZwQO5/LLCGpZDM7FMIrNqymBWlJmsI0R9e88tdhxRZyfm2olDRSTWsqJeyulz2of8PrTHmCUP0
X/5PRf9O+haCJBp8GlAzRwGrstKvsQudH1WeaEenfIoQV5f29ccLzS57Nwrsn46io3I7c09Fvlf5
ljpgSyXcPZwoBuLm7K8d3+7wIUfm7uYrSflR3ql9d43XrFzUDG+6l4DUWGzbxviWqrU3+4QFnMhu
rTMoU00oE+EHpWNMl0ggbsD8+0sjfzWoTIjp6u3QmZ4Hl0tWOCCwtyvXETRVwgUG9GOukQ58rIHy
jbKzovpbfnsSiFP4sfbNbiXy8K55sstA4NIgy30YYgTmy5FBGtTyWiKCbF21YKoW+Hb64G5f9aE4
7/Mq4VkRaEFpIsFeDKWV2ikxWe8/dhemBxlQuckkkex8s6Ro/Q2NInvcLvR6nwgLGy1Ci9JtO9s3
AiWhFPmsaomvp6HwPVX8iS4rtVKrXKbYHy2sOtnReQf7cFbf3KWAQBgXibnYjTlBTEtKnqTHFA+O
9CRlz4mLtzrrgcdArkkmmYzq29xJ/Oi6RiQEwo+e2/FmyUJCDjkU+l7rf60uUwvDJX4qpKA8ybmG
4GtFNSA2z8HlUu+5DA3zAiskMO6Be9hLfcB9dD09khwzNkH9Ch/2L/RTA4stTRzeSvsVSSJ1ydDD
vuotM0Hs1cJ46CTY3h2jyIw4ObiqhGhESvxviO8E5OCU6xEQdvPQH5W20QdWpAd5K83+CQuS8fyF
Jgg74wz3UqCcoykbUJ3aJ4ckOUcKDOODzryA8zbBqE9JFwjdTvtCOzx+v9QhPaCjB++HtTC0QHuI
EQYChAanXOwUUmv0JPnEvO1rPKJ6PZ3hFyRsP4WaRm7gmtB6zcLEgC5TCIxHp7lV71Y+/f7+TdJJ
+l6APGJlZ4tZJ4fu01co7sbplTYT13E4sSG8ETf/DO2SE4kCkrwrz0y9f5ny8LjpbuZCsaatz1CY
7rEPgaFx3KdQMCaObr2t4kKTgw6OZNyuF4m92Gbi+WvtxI72vI41GDgOllqbAqtTmK900QVjV0PA
w3q8ZTLg5/7pdYpZpx7orbHxoL/Yx+D3A2a8gTSuNbjymv0QPdR42oFddC7ci6E0vaDc5DIrAqZP
Oi1p1mhn+gZoQLe2XAN07NJHCFLrsVqPx7yuqMM3cjhU5Cv6m05IEHx8sOnhXjUjXpe532w8Udf8
GjXTW04zG4BQCuKtJgTwhBxMh7wsVKhX7rnB2eZhWgMRxQURQel3yNAfG8JcAeKpeQGIsKdozxwC
mB+vmQ3ecGq0usGVQEarHcyhih3Wksd4IojJjm/U5XUncuQU0LtgOIGrlWPoOSj+Ojof1TkHlFoD
8lt9BM3V5gX/EPny73CioH9plAOuIUW7RYX55Pf61R547/RF4K6Jvb52qE+JURidMiH1lJBYt0iy
6YIJYbkt1hXAPPnCxVCTJKdvgjhGVXQG2gtUKmAhGZZs2LhAQt3l6xAeBfnm80anUCxLUj/ynOvP
2CmQRIRlBKc1qacqXgt2sehzwA1pl66wXAPriYjTO96y0IfXev22L/rIkNRWHAU34LS6tLovBF2+
J/5c/byTjcdVYExT1lKUSjKyNdrBrkeuZRLBma2rBnge2WMOXyOycz/YCIadm+3sWTG6RlNZi5gW
47cW5jO0TlL9UwC2J34i/JKz8JQ164VWMglcq2UFcOYkZMj2n8osNdmnpX1vc3C+o6DkJuEdpVV+
/pQAhGkceApIq4zYSAN9sSNK1Gyd1UCuWomII+OpYXVSShtNM07sF3l9Z3G6ME3luWLvP7yhHyB8
Q9bGgaxgS3CzVwZCt5Samew6nTldmXlYRJRgXfK7KgZ6Mfhu181mPndhdhVCEoTOeXhPRO3ve6/M
UdZ54tZKilW75d6nC3Fr4wId1UVHWQ8B7x1gr1vxVaHh3tOl49Thuh+e6z6uLEWQ0qV42Ji9LWGG
896WY+gA9eMwI7tN8fD6wNcz/ZRZBsji1WyKGMbaR95+j6h1TQaf1nuWtaCNSEeiJXZYf4NQnZea
8JVz3t6au0mY09BqAewI53nFH1Vn7Ol/FVXpwZJATKFXO0qTtTLhbX1n32uRTbitJzGVF8wbwRce
JS+0eD6DQhi3xzaVjbdHCeNItBBM798m+rUuvbLlSkLqkiv0mLQaDFFXE5b/+0Vj7xT0NclhN6QZ
1GquYGtXHPxytyujIVFDaHsxnXZo5zWU1S9N8WIlzpu4F+H+45mut9BQS25gSW/MCAgc3pr9UJl8
gq2OS3JkMli64W7Hi3HkiZhu1S0klzX7oVtWKW5DHXnj/sH3BN3SnD6PRNBaPbBpRioJJbxBk1Az
g/c46h5APeVH18m1G1GybG5vZ8se9otlyawUyWrqJFxi5EX28S/zzsl+7ZhRf/eehbbaXp+1QvVy
Rs7tzMCiITGD4TQLhmOptO9iRGUUSRjymFrKsvkl4WESnJCdwClba+SO7cYUB6Mq+AjAiyCwh1mY
IUqDi66gASBDEqy9nUX4DxWnJmn4TFllp7QYXSPLwtXYUZabf1tXadqic0s27sxuD5TM91JZ+9DY
jykPM5SLjFFIjuP+1DahIpod5/WJeUyZguTAKCPA8epI4vDdLSSIs7+D+x6wq+3NSp/QqwXb6z8g
mfK7B4Qf+Ntdq434oFlP7UL9HkQTzVYkiq9fRI7WfnRbgvBvS9ELC6J2+Acp8iOhtCx6WsUyrjqq
NWQvu41skkjHD+XJd82/jhmzkg9uaa2oUefo+TMzIgO2XOmIGBUpniM7w50LXxEFrEuCYSSqTIRN
hDTHH4u3uZXSZlKAoSS0Cn+MqDzw1vl9im1EIen38ERFu/l2U7r4YCnAptj4JMC8t2GhVmYwZjq5
0RSyli45vN/LLBe3sqyUBMG6SP0Xgs2XCpuKE/nZLSeGIevkZ34hElQNz8N+fGCTRoQteC4IIw4g
Lat7afyMvHJ4am7BptDPFqGrxlR4eRx/pR3Rv97IBezBxV8sdOWK/qyxx85qItYGyE3QGuUcNEyN
afQlaFIqiiZUolYiKA7FZ1XtEsNqqHQDki5lRvzXdzYp7Nt6EZ33F8/v6CkNbqvwYyBoAt2DbUKj
6YbdBZ9mOE2PvpWEbFu5svbhnBEl79+GBKI89MVSk8v+Y6ACoiU3hQNPym00smlqscqPLvs14qwr
8gCCDRPmC/VCnjHgTOv6DP5veIRiBXlc6HMdbGNjP5PGgMIq0+npFvTYhs0cHecvX74P5+h9D9pv
uVSbSKRpy8AobBJ96slxbC6+i8i7M1WCDu4didSxQlSaBCO4Jp+fm9112qKoSQggyZdbgDWxPx61
PYk7K2DMuxFXq8ZU5vEfh7KH7k3To4rV7Lhm84HeS6b+oatuAoL/Pxno2IeLAYxU6S8UzuptmL+d
jnTRTHTM4yvcDyOEMi/Sw8qpjNt88t70i45fyyqQEn75GUhlj9Ma8eN6jYMQaO9rpgWkeUiyMbku
vhTKp1CC4Ccxl/w6dCfXEGvcHT2BpJkyEiSCJtV3atwtUaewqfoDp0nP7gSC/rODB00WXB+oi1kf
zPpxywPe2twADpxP0rBZO1TctAUT3WAewMVXl29Gx580M9kQsKj4jo4D1KvZDjqKwz6d33yDd1Wc
QDDkx99JutDwpzCv8ZQ6iMdBYxxD6ol03H6A6ts70HONfr5krcQL4PlavLXKzGfyawQ7dApxIpyR
0wpSi5eHmY8jOJiqnNJdhXb3rS29+/m7jncb4tzV/MYDCn4kUsg6Wk7OicsE6tRakWaGg8t5bIdA
Rc9g70ROM0a7BAdHWKZwPRiEw3MeE9EUc9cZu5tptmdoS3/btdCmYzgPWAhJ88Zvh7hfhgA/3DLg
xINADFkC5W0S3ZXM6+sdE9JBc417lr+ziliSsv/vBLT13arFwG1T/RICLpDCv4nqECjuje9wP7kH
qKq/gOJd2EoZ6EXIG/1E7gDs90fpYFFhLbg9kXjs9EETs+AQ+MiykYRHDC1GWRlsxdTwkpNmBV+w
dA+SVTLY6DYiDrwBRuMq17f8gtW/5TGRP4XkusCmtzZDMu/PPX+xk/y4RbdnFYBWm7V4yG7PQDI5
ddOGt117VFbF6L8dEsrF4gVtdGjAYY+SYJdsC2GDX+JVrT+cl+sZwpliRN2WUZLiJqJvRgR7yVPn
on6L46AMU/qWmhgeUIg0QCwo+kIPFY7/ofG2byHyZCosDtjf7oUP6opu4X00Rmkauz3sqB5wCzUt
q/dIX2N8nxsCRhdYtdy5LC6/5/4orAUU+MYcKljC0qaU9pAW4bn2gaeLoLi1BbcqPiDkTRUUKRdf
NkHVOud66Q9CrCP1Qt5/4TMhIdxlav/q6DpSmKYPJmY3dmqG87efBZpPwGKRBrj92YpJYV8NfDWc
yCERj3O6sDMj2759ykeLhoBraDpMoeg37QSce+tvL2uWtiE2dF3vTV0vTbA5j0pa1R3THjPzocKB
WP7D+4sbpPK2LvL93tHaSPQkDi/mLooq6NEY5M6YDajy9ksKMfYnXdxeaY1HBSSGKogramhCktSf
UmmSkVRBzkLW4UCEadCQnqynw7gZvaRGzRYXb2tN+FYg/SqM/+IZRw31TZhhKWJrvCH08oOnMPxF
M6Bhj74wMx/RfSWofh3KU8lhm+Wur7oDDS56vZo87WFNlGI7c9nKAT4srapdTGhGUSXcR80OeykJ
OHnCvm194e+G8MkKR95/GqJnTET0zl92iYB+w/5PnCFnhCGccDw8jhQSK5W9cT0/7t6fdtjTRTI6
9oSTwm6m1OTN0Ja2/Y4q+4ReDu2OGjDpu9/Mb6IBkBh/03LVhZ5M+zrwS28R3h5HghNRHiTDcVKu
LR+S4kuDq146dfohVantiXeFKP5rjhScdkoDQ73yQqa+EW73UQxq9LK8gyWDDh9kT6lSRM/EG5hy
sz7D62q6G1qJOfXG9y+ilYRKJkdmr/YqUpK/vl3ktYfTtqjvh/qy4km6f6FsTCtXyVm1QcKRYmbr
IykoMTE+OFXxW8lZf+EV6TGCinFnc+oiJp3UJwsg4ve8dn4vp+/g5RL4R2dSfUmg9LGtvYy4B65z
wUpDK7YbiL2tY66rkyjmFfvN3FPP96XCvIZHz1s8GJj3KLxhPDGe11J0wpfHeuoY8rCVAADp64PG
E9ts/OUpMBBmxLAzQQjnDXLA7piwOOTIo7U4moHQsGUc2h9wapWw1f1vsktmLCj7Xz+jfATbywIk
MgZ9T0oFXJJcP6TeTcJQ0IQT6nJ6pGU3grMW3z0kmUlf4g1vRNIgnXbGMWKnqleRRRkeLAjGIjpM
mll49BVxuZs1wDL8rGm92QhJNzWPo5nVwmxZzFobni9eeluSnHaJIbwT6QAy/2Iy88lRVN2+nLZW
YpqPFaqjaCTvGjQY1KvF5kPgE9MPHX6RgjG1ezMp7B5K7lwFXEL90rlYo73PpPkgQGeDQzIZtNbD
swWxIMSwOs6YDB+rklLu4Efeg7IqQWF6xJaQblZXxGdVAfUFTYmoh6RdBYk8NFRG7FNIZRswANkO
s69hCKW8ic8ueiaHD+pmMbZ1PpTmjYm3crHs1v3/tHY4B2yTyNp/4P2M8uKTz/oKWwuTaF/VlhcJ
nJS6PM4ves4F9I2wAJiPti7u50DKuFveh84Szs2bEYzcaUO3ytZmkRiREb6O2sABseHLiLYP7DX1
t57n6pGY5kBIrWissek3hbnVXG4C8kzbqOaok5LOypyOsqtCoW5M2E/N9HtxsGMWIyfYhQH7Kgmv
uFA1+3bIxQibnBwJP61ShMdwwN5Fzy3A6fZ4G0SmWyPaBpi3uMh+fnjm6DlGN9kRqyOqBDpl0lSr
mirrfahvacIyAnvGZPeP46XbeY1mb5Fb72rzUGP2WmmzkK+Tu3mRtcQYY5KZsYqfhvwJN8WrhXFP
YjL+KtTlcuM65zTtRenG/uqj/eIQOHbbQxfBTQ7XTzAqsIus0DN8N0r4UnbmILZqCcn8yq/oY7AA
UKxWPzwNDm8YX2RzZYVmToMmWZUfXgJEfYCFuqI4LsHKFhsM3i46k13XoceWCmssuYNtrvVVrRkA
tyjuGD48eZuLsqZ8y1+dpcpxnhW/vkKx3YORnYUPFOXAuPMARq+zb/k2R8IANvqF1rsKTdzx8q1F
1UU6mPNl2bMNWQUjDyMhHbS4WZeHS3ARwE4U9wbKD8XpgA4rPVEBCV341p7uuSYaoX3DLTMfoYVf
0iD/eYtCqfasvGZJvBe3GbNN9KSZW0V1vinz8amdtjRJp8huI5LsMgzCsvySYIYgkYpR0X6BNMEW
YN1qusvTJ5fUffLZoIFfhNuKaPVcWftJ4V9Ek9YhK4PIWGlti2EyWcYeqPnnx7F1bCF6V2BkH0SA
7riynN16xR4RzdTZurIIKMZonTp4jbdfifBwSDzYTyKq2Ud/PyIGJiAfKM0guzwz3nY7c78QbC3C
BmDb0HEdjeH5E8gYp4UBkXdmIRoQTiE4c/GQ98buanok+0+FBx4zVCYq+M+0ZhzCQ12LnLh9D8Py
NAOxQmZNJYv5WCTyAPUE7+oD44BVHhcCpFVHcoZzmYnghrWV/nPnUMkri+DIiK7JB7rg7HpxgOUC
9aAbfynZpqkZqZcSCab45YkIYqEbwz8q+uD3mrgFYTAuFl3G555SlxTgOasetuIkAGXacEIL+PZ+
3rdjfppMW49GwHG+9Iwy3OcPjxrbNI8P1zOoXqk8qftBQHFrpuGEwR5Gcku95d9wlx3eWjOdEqPV
PGViN4lT/wpD4kZxqjKb9LEU3Gx0sjeePvysuSK9QF+ppAUv4IA6tVCA6n5Zm3sN7f6Ph1IftAlb
AvMjNFYY1JBAhLf455D62QazUyzt81M1MKUArQ+Q6pPEps6y6OSFInjXPHVG+9EhXf9d2go5A/H9
/ma54H52xZa0iTU9B0Kpo6nmMjOB3+pQ3FjzAXcecK2j8HZJGDzMQXnjLlFjVnjDV2A0A0Lq4Wue
A+kZ8iIyam5eRC1dtFmUDoQO1Kp1IudrpFYM1hukW5JO/DGGEBtwQBtYIhwGQCwKLouH6V+fHcxF
5401DkU9US08LIOGYX6cy0jNmN8wlrvNZrlrB9FIT9t53Hwhzq0D8FfSGXRJYFpBYKEpalrqwAID
yzHdhAvrMgRApHMs44hH1uOEgEyfAtqkh16X387pa1SVmSB8R5B0sBQkcLIxTnS++CLyQ/suz96z
Pjlb4tGCmq8ITDRsanJO36SyG614Sqc1vf8U1VeQWhzYaDoS0o7a2QaixsBgLzqhm6ttLa1+7E60
6L97LFAK5nAwxMH+3qasaAqt6ouTOEokkPQje3FFSEBcfbfFS9mmgXdYQ2vGAn49gff6W5YRYOgv
jDtBzX8fpHqofDQW8yk5plzxZM374JBzdziIDsfBAHBDr1qcxjTe84WwUufgkdrTWZOf1exTI8lx
0BY7GXISrdJyTjMrhMp7SQLp9MfBbDWjKLLFpbolkYH9cB2iRAIUXtHAXa6f81G/cURSP8DVbcCa
lo2OqI+bDhw4MMQrVkiRFn5e2jKkZ0C4+fnFM6MSldC+XHgfS0RDsajFVakdDxN4QxMZhkQe9jYi
EXsymroElCsFhVmrytQuGgx1yopHg+AWdVLAl6zgdT864L6E0eOjaW6BECG4yudnht7ZmmRJl7w+
FBHNXK6RoCVX9GYSapzbxVS+cZDz6PcMar5++TLK1NbEAkhORkovUdJscmCArYJ1DVLMuh0Ep4iw
KSYc9Iui4oYaZQXS8I0uvKPZp6xO7s31KDrMZW3Wkfy+qL+iI7tuail5w6XjxoPb1yc9cNBBZz4/
X2HtNXg9N4/lDgb5qHylZdlkEP6azmjb7kGXAcmNphKmrd+2cjh8hy4nmW6nc3roZiUat0UAJ4Yj
tcM11Jl4sht/7stAhGiyGYzWHsJUu2DGtg+dj945rcfPyj0WeAAFXVszREgejgE2s6/C4+KT9rjM
a0UTD1VDKKLdeFylkRjlU9JBCZcU1seEEGaqBaMslw5bU0PvlhboYzppXJ4d9rQId2XdXX+E000D
MTHGxcRa7Ek1FOK2Rlc3COG6M1pmkJ9PJHdIH7ta6tbqOJJoil6hwXE50IcmV6LUMHUcXJ5yvDXl
nalbwcXh/NxLV3gV0LVj/pj3Pdv/og3dKxPzNegKgRniPHRRQ4W1VVzOAe5mi5gQHgpozGnSzywf
X+V3cX0Qnc5ZSn/Avg0e2xybblKJna/q98FLdAiWVqA5LjPzjpjFmJGoq6PWQ19+GHcRB/pnRop7
wLWqnfJ/6NhDdm8x7h2jlKeVXEQOVCs/iAWMPro/05DZ4+iDADbLjXETk7LTtBbuj4/nS1HZaOtl
7ubwJUHLTbkDSrTTghv3jsuV4V5D6IFB3+fo4oY4D0O9A6ac7Ov2y/hKoOjHQ3YyjOQzbKMQdTlZ
UCM6grMyonLmYGG/QJ6p5Lgbk2gipp8tOv8lqbe6YgkaWvTu3s1bveQXTzk6nK3gEX6m1d7LHvFh
qaLycAQKW+ZIlaKPCFHCYVBrU/KS9Wbapm2ndyEf1XEXXGQjlrR+ajQFGCGPMeI47rYtgZ64VerV
d43FioVsG72m1HNR2/Bad7tIiIcW6Y3vPEpkCG6BjzACFaqptAB5OCs7zTcFyXdgc6zZqrzttPzv
RSZp8SK5coxrOEJNmL2NsnQ7RnVP07N06wwJAwakD4IvrIE6HQOQBuMrBWUgye7ZztxWoz/p3jb9
/IFLkdgjEsuy1ccm7ybfHNAL7jGL55XdpPRpR/IegIX5N6oe60Wj09lleP8hw3t6x/91k5e9LFWE
qAIzXi0Hr2WFZU/l/wJ2Pt6ybMpc9LQOTj8qU9iJcUsMQAAPio/hi5zV/4x7NGC5GVc85rZJoB26
a0yvmRBvMPIU2b1e+sxzm24JOcFhzgB0MuWub0GGvIhXVdF0qAl8r+pb5f0v6s85TMUfcALN5a0F
Kl8aGeJtGBN4FNrie2e1jNQKYimvaZKGrhRHDqF+c0urDtXIZuh1eMBoDuYIBDKj6lErjvWqvxcc
+ISGzc1e3Cc0Pamr/zXfSJXtOuRvcAdu2JzjJaC/G2sqlIUG70ZeIvIH+apg8Tjo1mxykLrJ7qDl
hGsmyRpgmjz7igrb81o0zLW6GlqimDM2gmxc+FyknyfkU0nepmD23jV94vUjTykXPsbKRhYVu+h5
tHqUrxA/mXMxjhKRupfZZr36orFHN1Uoq67u6xANsDdQSI2bUpv40B41cbwz8ur1SVBuggkrWeZL
xExiLvrCDVnkfr3eGTBcBSjC007Nw7M6/9yqN/yNZRsFdDBlJYEqXS1DHBDffXaE3WveZ3MFTl6h
AxGIpxNXbm47Tn7Ot/wTEliTGS3IC+kw+d9DTeVdqVf+wKkJbOOqXJ7v1I0Ba+ibxjHPv1xXLBJA
s+BHGvjOs3cXt8LwxvjR1kJFsWqE/yO9cGORyS46PGlQvmMkUNDm394RL7spCNRRHTNj403h9MfI
wlQmy83IXjPy44DvvpvzL6fEqluO1pC8YyT9SjveSYZZc+hZy+CfPm0VyNh/ZyJWauKPzfePA95m
4SwBMosa5OnaufMD0dxQ8u2r88juKSseZAYskv5gjohUFFy+DEqUGdQIuSWDcWjV/4eoravP8VUn
6kaDjWnX6KPj1IraA/QMWCaYY1su76G9PujSe1RVcBSV6+FYUhfpOp6+w5LSfOgqlt2SZxTFCjxS
Jr9321d+zyv6pQEAFRV6PqxlaSn+8nTjQK8LozXRhdmPVKU1+FcBQx9jPDKr7IIer+Adtc/c3X5Z
IbBTgIocQUtdxWe+tPVAOOVPG8/LEPBp1EXEDUByFs6sXuXMJx+ZXBQm5YLaGHTT7wYby16d3706
tB+wfidZjEEUkolVvkVyfNpIbriS8WRkGOJ1Ksjtiqaysfu0YvB0ONKuuPr9sz97unsfx77MWgdK
gbAdM7RORcW+MLS3d1qT5EjsKV8YWX4kivkMbtxIhCFtivtYTY/cazLxSK2b6EMF20V/9GOkaM1X
z6ERzySJQ9funeO9P5xYBUpw/lOJXrX9HhC0QiHc0WRU1zAysO5gTPaBStGsNxYo7Mtoh6Zg9Knd
zNeUe4D9ZUEOpdTpJn2XIyYi3lfjYI7Fqqp+tmWhYvbcTC5N7PFhAiwAwTKomr3Wk8nnnGe5NCas
3979q5NEdIa0XmM6ubd9sutwcwh0eX8SPzQIFC7r2AXYaMC1Tgfrb+TnxAzRMdNFXVLNeVUofuiP
9pFncdp50OZg9up4no4TNMAvvIwBwWnShjIEearxTAj/YjOeGY4hmTI3F1GZ8I1E0F+HzImIycdu
0/uVh21Lg+CqW/bb/+4B/J+mABvsq9udbidGCv49YZ1YZoDzhNqi3UKaflxVdwNjWLBkK/+p/jI/
+fL8XufFnPax0iA7c5myCm/3GuCwkgKED8rlqvAgAbuFhAtUW2NYjyBgYD+PReeADjMtNxSKlMue
vsDmk7wpnnWc1DOqvIvlC652XaWoOTbiFj1X4vDnNXrl8KywUR9WvTmOzXVF5ETl5i58ePjdPO0a
JZ+2k55oj2UU0kR9o0komzDfyLs1bbVBGac1ylpjbIqBADedQhlPO+NNTH5ZoDyorpARY5rqvedN
kKc4NcRTajGEHTir98Ebju3JJTSBt909yFYuKogT+YBSLjPkaR6PkzGhPL85On/+ODmjvdb8R3Rh
PkkNs3RdkOJlDThim5+hvgPZ0aan0bBN+eztMIwUltawtscIy1KbO0zWQfa54pAdn3rqxtlaTgl4
ZrGR6jbWKNHLXLHv24SHTLhCSfQf9saeFrXkIH3IFRpTHB0gyPgQFqNZml7a4jn4fnxWfq3LK01P
Re5JfoAIEGdYEJ+fj5mc3kTVV+s2k74zc7yn39ot5LqxOT8RUu3eXF2rYT0lZKJRWFDnf1dBlCg5
NjBWOe6vHku729rVX4Nqj2GT36w/JGjOOxkc3LlsVRIkBfeekmWU6ypjFEOy/fkJUHtyO9hmMoMD
baIByCZUmsTjYCwTMIgOCxGTj6J4MF9djUYiCv7CPnYtmC9NxkGRLy36qC/Sqs8RNweCxsmVtrqK
elrYcM9qJj1xpWn6MLiZkLmb8yK96bkfftgk74TH+Qx2tdPxu9un7bsLeahu/uRwxyqcGz8uGYj+
C07tIJlS+23jRbWZp9af2Zi7GmLruMPcAllPTO2UsTF+ziuJV6wdY7IXcONfO3+NHZQFE9RecdTj
GGrZW+dY8BJ+V6sw93MI4Dr3FF7hHO1nuyF2M0pkUo5oke2+GB73CLNmyiB1zA74QP70stLqhWKP
NPcAsknQuGoWPNPqfnHAEAxF18/Xwj9RYGLx6W/j+62RjiX+w1Hk8mMU4TbtRqi2kpPkhHFuLRJW
DzDS7jKSnPF6HW/ABOe7CO48copvsWIYLZL0miqWphhgSJBa3NXx9g2nXlOHdwBFeiGGGlOPjmTx
OI8RFyp5KgCYwf3ml2W4oKRTqOpdE6kMT/4XF/TpsxAeRKmJU/fRIuqHnAtJ2wPWtzAglVy2P7PW
Mld1REhbZsHGBWhvRgrSKvPVGw2vpvqYEMajr0aud8Heio2uM0ThAOR/HVbM0qK1wh9pHx8fm/dx
JBim48evizhNg941eMBvVQpfO+2yv6Z7E8Q04Qb4z/v/25w5DvaB2PgBcq46tZf2LtwKbgfhvEfn
IZon+nYxjFq1uIlSu8VTOaFVc3L0569wksyJotA6xggIc7iH/XblF1pVHDb1OmO26OPqpH8Kp8v5
V9oOYGwYMe92+F4MvfoliU5c4b/35aIG3wRIxbdOyxnG0+Fik3J/+4nH+rFP0Rt9PRdnSypYU1+g
WSlLAPzeR16D1o+WPWzG5wIlJgzg68XAtHG26jhwhfDUC3T7jqC04j615kP12VIqsIy+9LhmBt65
HCmD07Uw3VjmvDrSgPcaeGvGuf5lQrJXxC38UDCG4V0pp22OU8odOWjm9b7MqwZoRqjFDGP9fZff
EdfxIYKfYL/hE/0MdT+N5Qwr/Ob7wh1exTP98K5TyXqwf19F11jgm9K+ZPpDpOfirTHaVs73jcND
+mlQYTpAkCkpN9oB+Jg+2P5ZKNECqGXKOnNOxBrds61BsDQMLV1uax6d7kRJ9afZZjR9QJbEinTL
IcbGbQLeuD79d+Z/xo8+fMYGG0iNm1N1djJBbLs8x3rM3wGQ4zCWRxjxx0M/Y6zyMjqb01xpS+iz
EWx90PzDcJtO1/gXOIjfC2/U8vAxNaVBnhcR6qm9LkxsmwIXnxqoGDV/EkT1VBi/3imzUSrRxoh2
qpuMLYzLxVgz1qOlU7WeL1sxetXSDryy0Cym8pe29nfBNvvPZc+oBLjabSeWlIGoRZQ6VgjXkNAd
bBSbRDJggvFDAjdW0+qb7QQekcbLlLV6fJR/ZfNF6S4+68ZdEP8ncD5wC4ztyFbO0izBOuDZ/88K
Y0mXufegFJnoDFIedM4l9pNJWMgZfRdAkijFVsCg9f34tN6O1qA5a74jqfxDLcDEPdaAZNlc6ZTW
VTIk2gVZTAFufXSirImSViSsjMYqQcrEGK1UVIMh9IkjIAK+ZVLS0AtsSNVmy3zudx/XWq8pNvuM
9Ga31RHLa5VleRWLeJFvdzzeDqxoOnNKPW92nZmQ0k8CLcsNNm435xKy1eWKrSwrV6Uh0osUQJSg
+yo5AzG0lIVyzDucq11zht75rT877mQQ76vW6nLWPI2LYaF728VzISGl4YC+QejBUAtbUaJSPEt1
I/EENbky46j72SvcQxFx3Xp/ypbVMVkrQA+4HW4fkVxumv63fJu83+LQQmfJdsqJAUqaJmLrYmYR
Lr4P0q6yRTIDtiYAqPHzHzwk2ads7UPRH6L5s4sfiXDvs5/d8gklaq5fnPlCVWO0Zgnyily5HghM
8Gk8Gj/hytrr89npb6AMTsB/r/VoTCokEL0tz0NVqASSD+ckSuucCftMo88FvZp3naEcqMbFeAyO
FLLOHP4V8+R3eGv8LyQGb74ghrenxWdCYWuV78d+nxNEhvJoxHh+pP/Q1u1DPra0wX2oHC+J+foN
zNHGNMyHe0GwbHnwt5a/A96CI+MEgYm+GoAa7x+C17wBzRHmWZtCkfOFhG10sSoS74oWGLpoY6RS
tubsl49+xLgdA62Dh9j+OAsxIIejlZSVruxApIc2RWt1n0jEC+3BKLe/JHKBnRsp1WGkc8PZ6b34
blm7kkhEdEm8Coe/mK1Qhjle+OETqObJKLa4a5HT/vGn1/cLSdVJA8iYnePChmLGIolZUN5RYpLR
JDSlidNADSM2//VxJ6KiU8pIbKBsvmvuyBhLpcAkaMg+Zlm0IrRs51nNafcbTgNLXoKtL8B9Add2
kjagHxvqL4TFZnTV5KdxqidV8hOLeUDPwif6vqJtePhZHr/7hRCp3WX5w7ZBFNvXIe2PuG3PmJaI
m1OXELlDcBspAybOAC/CRoWH/X/frEGZWcuIiRdsaI1Hi5uStgLmvJXg+dmgEFgZYPSoQqaGhmeK
9WCy+aO07YbeP+S4ySBQAS5Q204RkHwz8YmSsqXs9OAqZYFEhtDTiJj66KoCMguVFDBChZTcDpti
tmkdy8A1X3Ir/ZzlvzFjiE14ii6q/8O7slrC/J1KHPDYejUn/EJeCEd9lRlMLpKwnoljPk2ebZc8
eWlJFcl/S/co1xteGYRlxQKpwP0/4mkLWFDqZQwyTFa/ImrMzK0NAMmjt27RKf8bW67qFhTVkep4
OllPPURwyXNDzA7NsYL9wengNYNKo1iEYNZgC1pCWNa56i+HfSr/D3zipLQtKWsvsIUsAkgMw+e4
eWP7I+aFqxXEbovdkBprrlUpkdTJCJY6JRQUHWzrPasr7kzX42VYK26xvnGJyAjAUThcqn5QOSEn
Kme2GDjlMe/Ddw8XYtC8kmnFfs/GpDhAvgnzkN4cq7/260mE118gGl8oSzQwNrLUyiZhTWKm6F//
2hkR2Ocz0j64NkyG8m+MdOFYNivPhD4sY2ieNtJRQC2x1xgQ3U7O1G88RDEt+WA7ySI0Yc/+BcRL
EmV/efjb6mOohW1BkPKt6lwRaKkMRzv6bVJ4Q5dLOHE/UYj79ETqylC7sIAH+mxbgFMjCXigj5Hh
xIcykYmcn18ZxdTock5gGPHByqDHpXagH1udB5OJvfN0UTd6LLdxs+KIGpomzojnqHJg7mRPe72F
oxkpIXotKxlN5cPSiQ1UfWVofJTakyY3rmgPIXVWSlzu79mkZ+OGYn6U67OBCVz5jTu+UzXclJbm
TKekFJ+UiIAKtAOfZRpRrZBFdW72RfcBe7nL7FW6cTKU81Zes/CmGEe6tSHcYW6kFwiLgVTPtwRs
LBK0Cn12xlgfvlskyToPw+gSFjHbT//pqcw4WJ39lJguA+hn5Dae/Z/n14RRJ9xE1/MyxsT6U2L3
huvAHPphmObXXJUFczomLqHhw9ETnCX246XjPVe5jFTBgFouZP8jHVpU0BxA4MhWkFXhW5Rk5o4w
bGth0ZfbYUxO9dh7Z714NwgL50xwEq+nrfk/pTDwmmaseVhWJkByVKO7oytOPkXTtyskRrRSJbmN
zrXvuLO36J3P+6Zx8aeoewgcVPn1cEw75M56T/S5a+u8aINZfYFAdhVE1R9Qz/4VMNP8uWk7wqDb
Za1DuenpIn86BYBtPqYIoV6WMqGTRZ95oTkyPr8PJ2Ih7vvjjJqXkGB829xWPnS8bvAG3lLHquVT
8GeJyJEJueKyNe1ZxEqt/aNZz8L7Qtwh+FUlqtuicmGX3xJwr9RdSaDfav/P8q41YWjtNC6ywuoM
7IeYhOaN/ZdG4QpAJjykc03wJdI6mzWTQgujPL7/Nyb7fuucm+x7PYtlKxV7H94eqZa0DUPC7E79
0djW2Hk3w50x09dmJ82RbHwOk7aS/rS3hDUywgltmWSRU+3pSRIiyRdH9DxYvy/wR35zW9EVwuN1
hjyeV8nt0z82LTUA6+52ugm/kE5UHljuOpsi86Fesc/7nfVkWe2Wp9r0I18soLa9uDsecKh65K2D
pTYA8vKdEATfwHtgAG+k6YI8vvv+nRjB90yrLsfm55Cb6UvqqoIOuiWIDDtBeW4uGS133WqNv1uB
0k+6c/068uzkwh1pCnqm6kK5/DIKz7akC5AtcPa5eXt/N712L3ybSm08tf14VguQgaSYP6pdo8yk
ITrT0KhVBM9n/dJOiNyPnBKr13EbVe+GyQz7CWZqj1KBDTjMGNI1eYKMRWzU4TY/PQKi7uRbkl4e
zOWJKoFrrr0+d0/baK9Hhcrg1bVTRUHeTc4sLA24qg8V76TGMVf6iuiaC5S1X6h9DzKNuPYFGpnw
5Cu5JcijTkUOou/Opx4s3dUkBvOPxDuB0O5xMyWe1txbtiPPtvGiSWxCo4Sa4ivVjlaIA2wpYA1V
mELYyeQaqNjto/ZwrGf2Fp1YgVf8cu6vLGiToebqv5HBgUSAEb06O4QrgifZPUVTcIxrueLyilgH
bEd+teVdhMsw7zIhxuToV20zR9ikxrMfq9PAEyDm4bL0vGBFVU9C5UrR2Zb2WfqOjtiqA1N0QgVE
60hwSB1duRdYpdxLG6tWhkgt/aRvImnHtJIbCFEVqexFgAawYu4udbTVTTJIpaQ3h6GnYUhvC5p3
bYbNhieYRHO8VgrFFXluMPLO7ilIM11YLe1smIGfyyaK3/Rj3eYE6RF2VW+ayTbJd1ersdEauKwa
YAnHhN5l4sqpWrtMMOd3Q+HsXzsWsimPES1ksC9pFFxe5rQbZ9O+Sq186TcxYvUz/x8aMyH4lHvy
spRfqahSIc9DTsT5x/fJq6LQK2I1zbn5xMDqMc6F9vXgRIkxReezyJ7gmV4Rk0SvSnebrOPTWGfx
zXzOxR+CQSqfRpNDovtJtE5MbJYI8QVa1ntBMKZg/zJS9UK6pJkKFJDICOGNusqk9yZZa2c+GMgD
OjILoc8NNgY40T8HBf1oije3XmfGBEtf19+i0zd+fg7EQEoxNdl/Yh4fpUC85jiWOQl2xk6lO9jf
SJ4ErbRv/aut6p6fx+yIPXUjaY7x1kh4AB1Uo9GGRdiV9x2RowOyE/2IU+DTGaFSTMOWFWHqp8Kr
JvaL6DEQscYx7OcZBkNAQc5sxTrfJoAfW8QjuERDgV+vQ/E8U1CxMDnXdq+fQZ+J9jAxFICAx/uX
+fR2GDQLrA9jwzJj1dm6vbvR+qKD33OyPQyHsjGpNVF0hBF6qDy3qk8YHlondCNtcCWw0qw7BKjR
1uUfaSOEP+1L0U1riyKEZRcTD1Ez83Kx3yK+ARraUjCsIQKL8/93XMx4rFuFspJyjGkCJKfgbyfH
k3itBqjcPZRWkHpOKmqXI2YRzTTNbmeTdubv3vxo+QQrng/0AoDoFtPLn38wwsT0fIDOCUNHaTNt
3kH5pCo3So0Sj/Zb/KKFMEqOPIq5CdVx/jfCtUA1C7yE/exft6upqPqY9clvQReitFYBmGOZrlMI
AcNKuHIsbdqpfUK4/lsdyjQK1gtXUL4uqV0pcbjPlWJm7oakvl/KoqVGMQxGI13vX9QwYkh0pHhS
jAwFXvguoa5/FMV8zdbObwaFFkvspjc+boM7fNCeM1ncIIPHaxvf2cVaRiPtahNb2rM3giuQtDJM
a0bzSksPheNUVjDv52Eb7YeSr9OhB3aHYGDKiRX1IuM02GFNEGplJ39u/dBY0Ky+c/60cMkbPhaU
kILfUaysL067WA+bEiegbDnIsoD5qk3ZlcPO72NRmhrpy9g7H4Fj+FpRtcW7LRbpPdOjFaUGj0FO
ND9dKJnNYdumrTorym6tC0vwaoBZiiKn5dkhITgifq3FXEgpoJcspwqFfhnO/xl4vv5uFKGRKs4Q
hLkM/jCDlNxFlp8rELBFrJFhUreyvz3H342JecrvCjNEXIfHpY5MR6j3tixj8KtQU8PR994tcg0u
T0HDomhA7AEuNpbzvYLAL7PuaVcEVeDb41ngf3YhYXsqJc1mtQnNSMSueVnyhTxMvFWWzFkdTNHz
r7TNN5Yg5z8uipkO2QhV0u4BbUrY0cJP3sdickj/4rmn+/Qj9EXg+nKLeBRz7KyjlzbdVfiIrFNX
cNk0vAe/G1E40S0XTjWHexop/ZmX7j/gqYhgFP0QxxJLutlJmtcP50QV0WQxj3pshCGYs9Qj9THU
6kH+PeJ4grzKKIgkD4zn0vBgkKk3W+s3xQKgXh58K1xYqEao8tt5rdQ1EkbXerLC8WNLPvQp2eRf
Lh8vQmhNPtKIeCgwCp8Q77bYPHklnl6VLz3SWNaA9S4Yvp7Kwi3sGVzh0aPNaO4I1/Sv93aAIPWE
WfS4xaRU4XQFe3CbZ5V7HB99ey+V3Andx2RH4/GAKtcochTN87H7ptsd3PTNo8GyVQOV4lfd/64q
LXYpf4utNfw/YB2ZSYhTTrrnFcpFy1XWFqY5Quvas0gLaaNd1TbzR5vFejCq8LA8cX10wTN8NGga
UbPKFC53Ho9FlnLvK73iDiL2SlCA7Yk+zby5UbByEg1wHNCPBB5EaVTMM5y5Kjf8w6QRVPyhBGPF
dAgbMEn4fk6bFRAuL7xK+I7dHOPQhtmlijEpgQMYZqcG/x788rO79oXRZbA4QDkezj9P+B0tmZ4o
VV3GoMImiTnv/VvFzoLVOaEcqvMg3ziI9RqNlMfoy1ap9Ch6g1RYKNOm6dLcVJZH4ZYxGvVm3e+2
9hgm3kURSbyW5bWXe3lWKGehSsFTzsU58qE26GgwTEwdrYq6AIhBo3uoQvMrjbEs9NW6NbktDHqZ
7noAAa7LzigR9sMsk834f2dfBbbm96g6KLoAMmD/AmX5Gg9pql4Cy4m2YiYRSZA0gIgVLpLcmQ8y
Gi1eblnSTzu2V3hW133Gz2X0EprExLvfOQXVgIp70dBS/vbfa7bEpfxX8z3SB2SavEh6Xak7z/b5
+Dp+5mVCvtlseEhqjcB4qA8RBfUc9/ohGtNTBEnl2Gp7fi05vyM0iDTF1lva1YvIudWlyILWxKpD
xYhFoSdrvvSMD4PDCJ1c/ZT3HBqOYQ21hZMUDhNTkeu7HT19SBdWEAR8sI+sJL+mNm8pPLtzz4uE
+u73mXdrLFM82WYPdyU4oyg1zC9+VfLiY8kzDwY3ubHVyfWVKsj/bFneVGAjmkOrf5C44I2EJHPG
mBhM43iCgFKp1sjqAnu/kuvlZFKvpvD32sVlYrVD+CkJdY/az4bDnZKENZGt1ReX4mC4IWww0iw3
yGTdaMd56z3ZWqxKig0/2eQ2nNwiT7AcXwVBpOmMooxPw8zSIt1uvxczTHKuabVIDBnCQ1V/E6Ma
0LVUL0A2N9/hzxvPEHR3dkiopS+Buhm3aXHI1s2HCi2rCuSbV003onGdKRwF8M3dr3SsEcOiE5C0
TlqxnDgVt8IrCumqVDhzTUpcRTxvZp8cQetrx8ycM2sccpe5IaG8aIP8gBdKNyepN9qwN8lEmWpo
+KWd8BC8RuoQ8g/b0zry2OuzsYi3IPSN5pAzbHPYGtu+mJ/jndAHpZS46532u0AWZQ+E/LPG2C8M
/0lGRGv2a3KB3i3aqiZ0mtkp8dWztcvf9JNWpJed1U/TtPWTE48FHSzq2OIrJAW64+RUKNVrtcED
Yp5Ny3PklCiQ+L7KSRla/kdO2RzhNCPaHIoT4AeiiRDg79p+WZcHpIxGtNaU7X7wLVFC6aKq0kB+
f1jGUXInq0u2QBJtNIzwHpC/NJwqCXKe3bkgJ8CWTx6WhFRYIMjk82sEqZIQ4FoHKmAW9UE+gMXy
d0mxdVoUj4/r8uq4tnzrSKzZQnqPZINh2kOJnTpNPNhgZczQWMcvnH9triQQEP3cztnZSUQGbHwp
djFeO+RZRzvd9rKeMsEtZK1pUZMcVJSknUHbPQpF8u1gsLuJmf0g1BxrAnR6j88Sm9zLD6fE0kge
mqvfDQ3SshAqfr3EdIFvLga1lHqczxw+GzJV6vLe6ofN/UBWGMc7iZ8jevLPsI1vmMXZIUJtJjd1
Ek07NiMjBkCo/OZylp2a0uEnwt96AijZOZpm2rtC7cwm+RuIkEa5eLBp7+P+eXp5q8o7CO7O2J2J
TKeE05GQW9e1J7+jwrlr3ZzjRdsy+5Fj5l85eqErExusLS3wo8Q+XkQ2kYohmVqCPIN0SF2XAnwZ
WfvqeXfsCvfFbKWJY7jDYkWL+IIfPGrq7igHMraci0M43jsYgJxhQgn40gAe0EE7RfN+sj9ySs6/
ifZ+TMPEg98c3hGQj1CZ1G5+L2sP9YOIaIfPrOpjxDbf7JwF+2i8hP9fmOgvfTnSfoM//HSbxS7O
A7QdRlsBw3+fewoU2HZdTDWZrGci/rntKVndbnh87ifX5tyAqovWTVOr/H2ueHM//H7cwBucebag
4eN/zixAjlLq3rmD8KoZkpLlwu+DswFSYnidKn3TGBcD2Z0plleQjntGa+exE7xWlD2z2/Sed0L/
4CHtYDyJypeuDNjy6vrOW0CYyugdqMwVUCDm5PbcFyOIBAboSZgeDBWFQxLxWsXP9WqZPhmL4mB2
Wy/3CpFIJP28H7Hv+WCb02PbAT9L0J//lZp3j8zuGeJPPc3uD80AH8hR9KuujH4qJSFqpakQPq7V
qCrtt+gefqFjFYkfto7WBszAQhTRz9gbgw+mLYrGvMz5aYHk3WszJIMVGjf3U+20vDU8mY49MhXU
+WcWbd+qX0gikaQC3sC/Z7S5prE/5/Ud8+zu0vm5V26QUW0VJHxTua1oubuTxDIQhJ4guyw0m0h4
W2uTNPXJ8Xue7t5URyYQIsiD8cwPIMeuJmV6ifeqh2dzhnp3kpflvzJU4lai+4co4pQAAJwOuB1c
PeeitclxI4Mt/F1OAYTZGKbDrDgWe4l7S4XlZzcyshjwnsvrk6SLVQ6jD7ih1T+uxSerRxGKwDyF
v4EVqPrwt4W/l/ek80KClyuj8/ae4THmbg+dxCZWdTbJZRgVnm6Vf/VCF0ykBvnmnn+XYGUiHhMv
s0hjiA13Ar8tJkzqaBee/EzjMX5t6qaqARghsr/SUVNw8nck8zFxumbu2fuGQntj+7GTQfAE/EcM
Fd9qcyCeljdym4xZ6wuaWhbJ7Q2Z7LsimAYDQ8SPx9auQ0CDhlicOqt+dSlowBF+LcMBKwufUH9c
R5y3DoD2xPQLT70N3VVgi/kKpEHNYNROEUrlRBHiXSBL3kr0DlJnEjjENhL5M3p2p+Xrt4muU7zy
sBUIK/EQ3G0V0kG1oO+kDXid24Q1jgOZY5Uh3D/T0C4h6iQqQOQcm7NMpuElp8+CR6NTvv63HPLo
YT1K9IzO+MdkW/V6QcPpdNpskO9KbYpMRPGnDlFOuLGbpHjGb0NGV9yyk/FuPTXdVaYS5BZUp4CG
aKaTSYP0dVQJxc2uEy0oIb5Dq/qr6/2qWYlpxpUZSTT9JbcaBy1JgO+Yrjr6eOGA/Zi3jr9TV5WP
SrY4BtY1m0SN+D/IriOmcEu8WEsjGz/KqzNSZ8MpbF8Wiyt25IKMZpXWOfq2EAfPv4w5AgHArGHA
a6zCa8DS0ZGeAt/HfOBh+7daKdDNuwvY8SFmZXkpmMs5wAI6deOAeXhJlksdMREFB6iwCB9YGVVE
AqYfuYM1m4xdOeEZMPP3+hc6RXZbOaWUnc/KVp5t5aHG13FrUgfe7K7QfrHizYFYj2h8QyIfoOjH
dNdFbTYqNYEvWuaxvErm2pTMmFutQSwduxL1UcJF32OOjDO7ZwQ5FyRfYl3rcQVd8B+nwJrpsPY1
oR0EtJGmKrvHo37bjLtvo1b/YmndBLwiJpKTm/Nvl6z0ZOjgy8WVouSZ6BO9onqOAVJpTu2eLEmj
9jUpiwyTTjKLDaBkybPokqtQRB0Uc77pCrHoWTN5iqza9xvotWCtIojMQ8tTGflNMZszD8HMhZav
9NDE/1YMX0Ugu3bPr3dr4kYVG8RA8sWz7k1Is5Q/UpPI0LMmZ21Q7XWb15K8Ugv6hA5t5ITq/bHz
qDD2fVX+ilp87vLqXuSu3kgRrO+rCjtf/fzjfsSpMJOW1bqU2TFjYj/ml2AEjppVZkxtWNtta0gv
dCircnCHowtkB199RMjKXQoDO5AhFRNw5RIDKOkp3MCx9Um2xYGZS+1zdhKP9pXQWHirR0BJiZ2V
5YIL9hD+qceDtNbeyz+/EVxLOY4xrfYR3Yo2jQ8qmTYLCudPq8zP9YlU7qh+nr+ztiLJmOeB8G+F
1LA1RLcw3u7eSO2MZ4BxJdEadf+nR8CPHUgxK4M+bHHVAzmkZYJwJxgRY1Edkctzs7bizijeW4LP
RNtrg0Nid+LfhFRI5Bt/L+AsXVKZ8C4QWt3BDPfT+fKCCOxjRyS1O0OUiuUPa3ACit/q0ZU4jzBy
QkVtG0OrXHHvM/WkVBYOyeYp1rpuiJgNqQ31qK5JbYytP2U31M+6vurMvbXBGzrdH1ezzUfmqCqq
HNiuEH1Tx2HcztPNe3+zMZ3jt09eIxT3fhZXRiSQ0vZ9b0jMzdJmOGLNdlN5DLTNSoQ3W0V+K31y
xdaMFNIOJ3bE+cdkxiicMgxXEFkmQ/QDdF2RToBK9eJT90rUn4DZ+9NtypfTGpqkQBAsAhqHXLEH
MLzcFpdJfS21ehOis5I4/YbK7KtRsKw3PyIA54/I0tc5oAYBFtP7GHQQWST1FVHoD6gi3Lzr8Cox
IceIWCkwBRaiub876nEHrYbpiuczgEvGxB0BwG1nfcJnRyfYbwMKJWGZnUhU57PXze4cHC6AIuzT
QzULbI6PLFpRfY+8cHhgJSF8Bn4Wt5FSBJLwwc+4vkMch/aTJ/5GzeGrhp5F7ZP1rE6dR4FTMVOz
dX6YhDjXvr81y3nT6ov3SVMvjriNAQzIiU0W4rS47mxzxNOgC4SNR1wl6t3jTwo9vnpbveUa4Eum
FttGWiMgwYvxHA96bpZbRRyWQOBx3NBKB0IrOkcWAROqAmDpE41s18vjZUaHqh8zW16O5LGQHeDN
BSVkdH5eJ6URGUKqMaXaNrIROkuMv3ynuW2z1p2doCmuZdh7mp8cWYvdUV7wqvmUqaq0BX/K6Gz1
BRgFY2bCAtKEOKbNv4Q9SjaKt15MfxiUTBeVBX4Vui0eOESnLRmBpY6PetEdXRMFBP0Ymm9mQCDq
p5Yzc9X5U9EgnQo/jvph8ieZ5z+hp21sy8oBk/wktxzVDWtflQI0fz+rzVr56EILUiw+if+7ySxe
5kPyl2laSC+KQmK6RuB/faFjBd0q2Y/iL12/3k0j27wqbxliNXWSmdCMkzVuSTLcP74M8WkWmMfF
gWoV0dKQNlT3ZBceve8IhlB0vr1K4ahPzXDFhPDsqjUQ4/z42plQaWnUw8u0+4vdnA7sRa9IpWvB
Mb1PtJHG5l0jTMFSFCTxqP8o58uMl8soVkHp5oHK9K1CwScPG47bF9B0PR0OR8RjZJliu3eDKyTS
wz5UAkEUFV9tS+oE8iAEdIB4mrE0JiitkUCuMCDcFQFB8coGYMde6V1H7KrssO+P3hHdUjbcKVpc
1irLYAXP8Rf2SWXn4AIyXsTSDtMCJ7yeiRlTQPY+8RzmrDn2yTjn6fKE2Yv/9VSOHXCsvB9Q+fFH
FqOdXMnBdMDK14X3WeXGkHxDTwf4eFYFFpudevpSbVVHHUK9UhwL+0g+YyhuBotzZtVL+9/id31t
WbkNgHPkCBouE4bWtVI5qdGVSoKn7nRh/XvNLH2sck2fLtmR5zzvtox+sjeIhs9eG9LkwuoG7jIa
PjCdAZpWAYRfHMf/OM5o5+rRkjQzZ/JPsxumNVS3doijy6TTgNlAcWqnOG5sVTHMJfZRXMhmpUYw
lRVG6hsyH1XGcwxgl+wEcHR+ufIyhh6ZGcE4HBxOvMzKNfXSSdoXEIoB5B4dxJbs5Q5wv+tu48yS
n/4o3oRgkxhhAXvIYm4KAjKyHFbF4UrVEajgHtjcS/oCWiLjXWeW+fG8PwkB6YBNAErUM7rHFfZt
/NPa0/JZZM/E0h7pcd7CRSO/jDa33H/ksyImm1t9dFPS1fXhSdyEh9Zcx+1DixCC0pyz8Kz944ir
u6U2qkWOAMJ7/3IngkqWqr/QaDcmSwJIwRh8z2repfihY/MNKWYT8lzrnRqWTmvnLc9NGJLp3iE0
VC8Scxvg1/vDPBTV9s3tryAWv/WFN15uveUaeF4XQNipmK9dTbjM1XWnsjfJx+9pDf9zrlFfe5hK
3rsjt0JnkS6raqJ5zDhRn0J6IcAfOK2MARxBneCc5Z7rkCm12dAILYdc6yvfaeTQXgwNcPBiMF4B
ZpngLGjRwhfGcW5H9ZUUy2WNoEneKW0Y0CMi0MECZxUxZ6dAuv4eRvFoBj3uLvMtekMg3UKhv7//
iiIQaDXtyF1CCKxV9veVbQaVBfAHTZnD9RpJv23OiJyRCsMGgN6kND0w6hdnG4N1RhLdpKyTe9iq
+vwbjGgF4waAMGe5y/6FmQZdkTkQ/gTP37cGeHzrGPakMeH/bYpj5GzsvcFFwkhCVjaLtPiWl/vX
ZehoaIBrbyuiEkacP7u6ZS+TUh3ci8CGByosBX6clVGDlE8JSl6RXwVdWJYgq4GAy2ZqvRQ6LgQl
GxdKcOhS9inFrF0qDWf8ESP5cIeeygqtTnIvIREQzKVCLTjpYZ8QNNrYuZKKNQQXyFk43j9qWkQ8
UXmp0Xqjp0CTuPX+tLo1q5bYu7QQiThLBUglOnI5IAPZrbpGdqF9czXk5HIbUCLbQ9CdKGTeIhil
Nj4eEoHm05+gFE6l5+ioJU0GeOKjCo2QKHDkaAP80UK566yXkkXUm4Gu5igUfuAOLoubeRv/DzF1
055TmB9xd4+qhQv/oXRykAmhmhENP+yw4BSPQNVQ88reh0pinrWlUN0ZUibqGIEJ9guZvSCvOt/B
E8z0f7pNkNFzAgC0LnMTAga/FZ3tE/+fjvZGvslbDklKjTxqn2x/BbeVApYnoa7k9kaQRRUOldQa
6oVuhTF+iQHEe+rUTLZoyfyFnCH01wT9Shn85mc3WIqxBWphZkwtBiQdD67y/uCPg1cX5ccF00VC
1TNQ07tewN2ATYAp6jaN4PmqF2JeQmK+dX2OnMqHn57sDBHrW9Pmvtzp2swMyfLI4x4Jgio8yG0L
lUcLrJxVyn9CjQPWsHuQ+/u0ZGxSSKURcZR7H7Orqg0mn5V9XXYaNSECoO9pI14vvLPZQkRwPgag
frRGD7dvwOK7ck/g5QWn1CchdoJOkNCwpdPu0vHWXid10MEci+VruQX4MsxF8YeuS82oI5vm4mkb
uojFpeqk6FqYBieKOpatNR/2yLJOChOs2iJP+jm9+ctXeJof8CXd2kTQlm4ljbXJnpqxIWpo7reB
UQmoedNPAW1aqU+sJIadHVg1iTP9KSl+5Ip1tOeWVVJ9DAk/TRGHNA/ghRTfFEdKFQwp96B7IllA
oM3sW1aWLQ1LO8HjB0fWIxerSGEFLxdjuJc+8SWO4XJNPdH/g0DLLudTTGHHxbgKAkuIgLBoLLbA
Pc6KtoOxbWUc7hmGWbXhy+JeRqMNR2oFMnMSQyCD1XLzFT8LKInXrlBNHxGglOXm+WKAOYJxbKCm
Lm+6GXp8CXvbBWJImwWVvWIq6/BvJh+RoXqJP3xoPO1QXXvm0mDNcCw+h6PHGjLhLg35IHws8Oqp
eXR+Nhcde7WdIs/e0SoVqpubfID7HBf+iDDmCdAg/Tpm/hpJbpa/9wOaYwbPLVHqw4t1ywVsOlim
eOwRl+1p3EWyen9bpzBLO8cVme5zK+ISdaUMKRQ7/2JQNJZllUobDVlTzIa59wycxcXvybYeyLZE
F902e1ApxrvJvRVdenTBbMds58BTw9sY5q7IYFnAXSBBZQQONp+rdQp0c1K+jErA4Id8tk1jdL9X
xIilifeksetAoo4LftNVqaaDUExBafGknjNgle6mVUUkNbWAKwa6sJui0N+1fyTjLqaK5CiBA7SF
AL5zGiYzKJakLLUxtbVRENvf4x79t8nGR7LqJQHLQ16FjLhnuz0tRIscLcBp/TbQJ2jDU7Am4OBd
XUfV5rsvUx+MI8lUCl1rrALA/ng85Ijeser9rtmvRRLclDdr8WvQI6br0uLJvYXiMLHdRI2tjlMl
JmRVmZQBNRbgu7IRmeFCvxfVV3OqG1AMQ7b3QP0U/HSMyMDi7VD8H5MUOtKGMSA0Y4CrP4HIojxc
hU1AeduNXaLiHB1LA7Emohwcsr7iTdkg5utqleFukZRim4hkiVh528n06aws9aBKxZ+0aEqBkFWP
Hmb4pdBpkCgLbRR7gaC8UhjOwyxgUGEFxJe2+NekGhg5gWD0QXGem9K4gzM8slr/0usUlszR/+1U
G7QuImjuY5GcNhVyWFaQmMF3J9F62EAisPHgAZaVJXpjU6z84AmVrq3yY540NOHM3xXbdSfuSRa5
MNTgrXnvFGSuhzKR3iblYRh3WMEd6hV6KPpP725m9HFSrVNmjD3ume28mE5JHoBQreNgZ7Y0Vlp1
hz1UaPmeD1klb9vGS+S/oJwNg/UIMvIj7kPtCYML2ecAuW9d0Q9Qx0ZpLe8TyeuhZETg1R2RVic8
gmX8q8+BvdLmt8dH4Rmzqn200IkvTqxb2v4yVXknWiWwyaCytYD+IZb5FADCr5eOG1tevyO0F/7f
FqLGuQQb2yJ+nvuH2/rCuynKL/3N6GjZcf9J5UHpMbIDYuH1HyEn23eAERxBepNbQ5A5vm6eYSGt
p1deUtvkedxjalZbIyEw7UzvKP5bGapxIL4lJncF4NWe05wN7XwXqTW+72wbMgKOrXZ1aqNc2uOE
fnLTuhBKSW/IZAfOrblnJY+sHOdA+R/hSZ8A/7740FSxlHtnIVKg+g8YcE+BYQqu368pCZEzh5U1
ivD5KGolM3Y2RUSiEfrxQu5JuHOP8QzrNZAdazBVT5za/96ZAYh/BvT6o+wIas/Qjssit1Zj2QFC
237FojwcnXqg53h7CJP2WqK7rDR+XmIVcdIdPz+P63tVIxGsM9GFKmJNJx8b6XN+KGSov7tKMPne
omBMZ7iVzIna/pc/4oV1i41Le5qf4EY4zBg885jenmTIue4JVJYTaIAtu/zhzS2YJ3xRL8QJvlQ9
Gv+9BaHwWBzQAQuwL3usRWv1iSTaVZKkSAdqDsuR8Cb+aGWI2hpymb4ArC0oFZahp1VAK+C4JckB
aBZcmIda8S8FOgu/eROK4iW9LdHoqGaImvKHZCqUhSeCdbXfSZDKSlpd4HzZGeR0aQYNZbvHK29n
M0iz8JQQBmRMEh/PpQGN6JoLDHeZLI4oeUx0Q+04A8z32C3zQ5ycM2OU0NV/XpgLQfyWfYlgQ25N
fEqtH7n9m9TWOB2H7IXEPY7kEMl81PlPXci7xhtKHuPYXsa11IVTWL63WCbLtcTZEniXykifKvHO
zPbV0hpR5rbSgaENxakuSYN8mvhXg/lHamI0sml0sNayyGRWvxd1sILgVKQXaypdAEPwl98CSJDA
AwhsGhqw+fyQTA87fPilDmPeevsts1KlcN0XHDB498UFl1fOmGDPifk2gmefIsd9dTLbLiu2/+OS
LVy0zVwwjuXTU2zNsG02f9VUem3cB+/bIBNviParJaweI2YgnW8ys0KUGCzm+OpvsDmyxgaA6EPZ
0AAYVIqLRgpW5i50nUfjwcD0tILkoL6B96YNeXUNP8iV8OfJPMIfiIx+NfnhHxL9OTOpWMN2yl5U
5wlcFA4A5+UteVevM0N31HMyyP3S7sTGnA9jRY8Wy+W2yMAuczTGpxVATRFE61p3bgfbCXM+x+0K
0pneTdf0YI7myWZhXP6NdjKCS4wk+ZJ9lH2idPZuUXrDzEqFpvnStZrNJmFI9KmnVRZ/wiF8mBcu
/xn9Gh513xjQD66jVxVAeiiT22J6N7cUxJAvVAF7cqF5FwULJSQMBuNgBtkVbAAF+hmu6wTyFGyp
xpYn5ekfL3o4JrTFbZC67UNdTY7gBIinNxjuqye5GS/742VzBO4xMYJqgWt64DU5fvLHYVpXPHa4
B0G8RHXEMeV/TN2CAlPd41cvg1YDt2kq+ZDaEXrYQRntyt0GqSzk4ZfgBSwZlaoQK388qqHYls0d
BWtznJOQhJLri5h6r7+gnWURSYDa5TH7lWWkmmC1rrLdzOZTqE3QlkrFxm3+Oldyx3ceiRrCij46
d60MsCabFm6UOM9soQ/kV0XywHCd1W9mpWHsHpjitFW31Epll+spdvfImNzhRHhff10OGGiNlYJG
O+pyCwCltRXb+wb5i7AUqRQO9gnsmsFfLpDpsJ4RelqfFgpC3Y2IBieq4l9KG8oFuW2ZFlYxb8m6
acWvPIJPslRVFZIGbi9MumTUbeI26KRNbU1o5vD5K8A+uS8cmZx0XDC6fj6hwfqvdllHdA5Gwd+d
KGlY7UukLKt6PCBUfoIS3yF6HWnqSTsTcjHITsCk8fN8bRkuRMXnFucZBYv3tU4HKVrnhyVwRmFL
Wpm5uPkI+30FjxQsEhnMMVYDWFRe/PqvhivWcHxZP/TjM/gN52zlY0flra3iAWGNFRWjGgyVuxOA
LW/elafGkxQiIoD5miXHeoiavKC0Jl9dFSI1Q7loxaRV/kJJx5urR1bNOcd4TPTmPFRPCff7bFs8
Xexq8fwWukPYjqDaHcbcZEv+swHnYecw/qhJsS5Tpr3zAEv1vH2UMLw1V85rzhng9IQkGg5NA4Ed
zyDzreB8Aoi9iLF65p3JLL7ZaSU05K1nt+5TGySEXgaWxy++lrZe3rrcjjYaRhdi3e3eFezcz+yk
0PYjxukVN+6RJ6qtwPNrrre5ksXN7UjWujtfzgDPXvBxqb1VVlsB79rBDO0ZxUVtzwSvtVO1CIcf
D4Y64x0ziKVH5TNjDvjwBUesDncaUatyfOfw/wSgCPTFNP5QfQp5cfOaHpGaHQAYtSmQ0uT5f13l
lod1EpB92Q8Mq4VY9t92JPa5TI2DkTFK7qJeCgGxkz/k2gf15CW48+A6+T6mNLhr4rDQYcGMLMXX
Dm+e4O5/dgMDIUTTWhufYzMYY+MVLhs1haG/0LhmJXzdPAE0s9e93oQAXWDHvKeBY/IszzW1eTCk
ESQEUtdpY1FjqHhMimfVNyBOpa+xq9mdmcvblfViBtBsXfVl5UzHH1e3SUCLD9zpcTjtkHmLFUmK
ZOdqOoZ022zly8+LOECZzzOC5cY5IDTE+F0T/b145RtdvI+dtaHsBx1jQfrkVeVfPNllngw71Bn7
LUkO5nR9t5fhSA9EFbPBSgmP/Pj8t4ivEitXNC79twLlFppglcJc9iVRSWORrwbmVadXx8C/S2BF
XxnbCbtZUY5T+iWs/EYpYCQAPRbVxWUbAWxqOsHQ2ie5vj1sginBsJQybTgSTNeAjyCTpwb3HyZY
+AqNaLFeYzLC2SeUfmp+MWAUxTKDDhHEbgQild6+IWwsfQ26cIQXtz3pNdZ1wgbi5m09yPFaLPn+
U/OqCfYcbeo/eLCrtS50XVe5LY1DZTTwjJgkAT/SDM80zALdwQZMZMW1KL83ORlofdcsJeytaH/1
nMJj+fBBpz5/o9WqRx8FXDp9AC5uNcXluIZwThWUZtVhH/rhrtwfPF6I0BlbK3AA0Y/TOVW54veC
AGRmWkqC/dWfrFk1sS9PUaneuMzpZO+klPERDqtz563mTgzpZ+BfYkwrWxAchnKUIlNZOO9/BfdV
TrEfTdTRh1oEPEx2m7MwRvOoXri+yx4oJiyBpZERmwhVhFxFGAtzqDRCj8DmzJL5GPinNO+0pkPU
hGcfcIMec5tR9zIyCa8XppPcsOP998LUkmHUSMV+QY6HWYtOM2KS5n12EcBw9Mj4t7xEs4vxH1Hp
fgoHGvfhIWcnb6Ndi+eTYV0qtlgLg2lkUtzLMOHbCNaWQpivqB9b9Srwv0paOrZ8T8bM1HzNcaDB
YXmOwk+rZSu+oJ+5YlcqC5P47Jd2KjorVHdEgC+SopMXiNp04UsDe1HFWjKfwLj8xBtY6OEk8vtl
zu7mqt9z273wU0R2rkOoDmp69kSTySEgAmbDLpbXdLFF0wtzJvYwBTftsO5w3qeJP3SL/FeIrC7Y
B+3fnJGJ9/wNd9I1IZOV/ZMtLKTUNMpfHOj8o2kGSBMx+KGIY5pxIM3n1Zu5UrBwdO8+PFTmQsuP
tCjqvhPBttmE4iD2b2iEiiD1gKil80YHL6ZbgRlytYpFONsSra9bJqtNsdoL1S9ujCX4wNOmXPmO
OzRGX9FE1fXO61PKlvi9hNxMLDPLN+N9g9Wd/gZqDfhmhpiAcWJXEcI2svCoaJ6xd3JyQHL0pEAs
7XkBsG0FsvxAPb64RhUXETTrOaXpWVA69T1at+KzospIuqJJDRVQIvOBwZbJbo4xVavNGO9k5lRd
0wj+UhgG6XoasoQFYHM/AATb15rqVu58msfdZ01UMBIPViPfxkypfQwY/OfZnLKwYkhqtSjvTPtz
0fPjADuBD2kNLjIVBFMAYu0gBolJMjaLb+NfesS+w5LTF054dATN58aSLWs4w0Y7GabWu63NY9Ne
p+FPVEOMDdviuFAQG7UQCm3KN2kyTtilalDp1rLbH0aPRcZ15IKB6NCIVn+VG/G8QeToaEW8NSVE
VjxrX7uX8p2Xl7Fx3tB0cq2eyV0n2AViAgwhQdas4JSzK/PQ71UVu/fVq/yYG7UaZx3Cfe8ISRL0
AW6gmNhKhnnwIaq5N0ORhU9BCzBbggdM7u6DD3J/7PjmlvsEn82nmMn77RJjbvxLYSmg4rdP7YNh
b9uNNw6QqoaylhJPfhhnVzO65rGiLxDs+jn8TaFJFAFUNSjvThLp98UA8KiaNNDQGM0jgFMy2RnX
fcExrDT8X3jWEhR0zChmMLi1lZyFRtcBwrL/Mjd86wTYzc5xsaZ4qj1SSdq89gmnOGTjhhjM5wLx
n2ds7syrUW7RFe+LPko+1aAnj+0jKw5J/nzoKvtqAaN4rtXt30bn85gOXEt+BxCs0FiaN2VFeWAS
lB7IHpS8K1aajWOEhntIeyecBR/FPsGtmBr1nIDllw99hCkpImxrc0NfST0ublgY7fCR+OPquoQ8
e6HeFHkE1dCoy9SMx9+aIfYugUCNvEKwov1lXk6ddkwg65TlgEMOdXK5tbjYjsFobZ9gJA7PQT9J
tWoDFJcEvvBFHisswUuDT12RC9VFbGahwmgqMUzET8jWuUcDA1BXjE5hdAe9VyhX1jtUNecPS/yz
b9UfvyMcRe2CvuCRGgL9URKrVKa3WdhDAN9m/veeL8VuRwSS9WbO5g2VvatAyBbpUygPDixvd+CU
1UwSXgUPsIrGdvaZOLKV0CuTSQQjPIttbrtzdVOSSYmg4EMUiJiId5UahhzFg5xa+GFK/3SNCarY
1lKSQqUoM4nvaB281+QY5y36mZygnq5YjIAq5TVDCLAtPrv4KazfnYh+pDVeN8xGPZFfuM3CZjma
RQFpZZvGBOjBEW1b9V13dt6TuiC7HLmBRES197cVQBOsC0uSpZy822Jmo5BwNRSoaN94mL5J/Q+3
mf8kf7s4MxqglQTWTccNFvN6RaZvKULUAGvQ6DVmAXR/H2Qkh7mMRndScbwIcnl3TiZbOCVbdVmY
VlxgwWFatpAh+R7N+n7J31784I13qLadcNxc46GTzrb26swuMXjEEggYVl3HmRJ3rmsFW1e62ucv
1dcst6AvjVNVgJtWhweGMDub7BfyU26OMsXG1MbaI68PH8yMuW6+5HLBuWrkTx7vx8pKVN53bfzc
XCvApMl4M45l8tu2N0RbccWDU9wBQuxYnQNL26lN1Dy80KdiaJ0WY6ves997zpRqkImDxiMVhE2T
nl+4rfY7brfgiIf27l4IrFDxv0vbc7GLiB7qOryUh72nX7kDR5Mpj8jquqAwrKMRr4fK7E3OoyNT
W0kd70/J3T5Kh0O5f+gYKe54a6tQtIVaihF24pYwoIyXGipCqqWT5gw2vAiVd8tp6/hUadtU/G1V
HkksbErJ/c7qakG6Y8sRiG0dCdbb5704jvgJ84Pd/I1kIzx3c4i847Rr0MQTqkjOmmE9shUXXict
JyZyVwoYseIkhDOQoPYqDmEVuT8aERMLOPbCyvjxgkaS4NdpLfri6Oiz96qBiZzMSY8QeY9XA5TB
TBbgiXG97LyTnMNIdTycfsUtOln4tP57t78N44j7/CXwHNSY8BNyQayZ5ModN4yIPqjq3RrtK+dR
C5413Ua30eNQkbMLGYUUU8MAgCfgTJlRoQukjscP2GEZkZgGOjUhu2siXrs2JbDls10CHXxbKlrv
AQ3AlCqka21S1chRcbkfLfGRZfr/exALC1TIhnZi2ywnluraDP+BcL4siO5n7ImJOp0FTDlTqc1/
1rhZvfCLMLFrNo2Mw6ctbLcXCqJN7ym3oCikMezFX0brDOnuQ169ETwAN5jkkhagnkwj0P9gjxgW
dQzz9Ij0I7yAqW+jmdCCMPuFtybvIfDYe+H9ZR5kk2DW3eU7oHIyFFdyk5tcryM5dfOXdBuuZF31
SBqUlDTWEL9BeEhz56L9Vz2lo19JiccaS4uRvY0zY7oLIFqjsr6kGVpl1O2LvVs6uGUte5XVNkSJ
xInIzQg+9tZQLglh5Bdzmt/aoVgjPz3HrVwaOqCIEcNIkGjykIzT6Dzx4lOxVwtTtTmWBNDOha1V
SPJKN4L6O0HAtmm4aF7DekL4sRieNAqIdHMUBYJ5mY+oA/miasfPaW9EVDLPqNK2lTnlfCyyW0mf
znM7VJmW1ccQRGUM7qk/LWvbH3MPBDFCvt/eRO5NAGqErzAJxsQ0N8RjMXnGamzLHiUMHXiwLtDP
r00RmKpL7nxFWc19Mtksg0G2lxUnhIkSngmMLieJE1l88o3WgeRXbz66i3K73dfiX6+eBGrD9cKY
ETm4HgO9lwA7kvhvsr0AcxoyzWHzL/Ew8vK+S2hMGalyquaTeYHk+KFX880bafNqeQXDOP35Re2E
PAhfN8dJv5akPrkCAtx+6hNGGPYL2lbM8xS9vK+7yuClOwELZXROXljXsyb3YcTr7zHyTfC1C59f
e0Ib1Y3lEhmuN6wYiHyyQSJsUIUMVvryMRYurnnqdcvWYMxH073vxJEdhEWBHW/lD6icSUsje3hP
gKhOjRtwRhErxtkpGlrzs3e2WTDhhPE3owHIoOdJmfnyuLBmqCtFM3N+qbvkM7P5dwtjBz8yHNz1
7uF4p8lkmZ0Swc5lSCu2QVwZFD8en5uyHeqfgKFi++J7dWSw2YmJ7fsgTtBzHOADzQvgD54BV1Hk
uAXeW0hPn0NEBc6syMLK7ekaqE4zoKpTojgaY24HD2T8JZ2EHlcuEJjCP+WZ5GxDMdaoc41XjLLl
DGXuLkm8kpdN4LJbKgPuRWyUTT0bU/KpAoJ5BjevEfEFO/M2NIvVMoRfrrVVqx3zRO1zd04S1qkh
CJIcZGLzmVVKyRf7E4od/yDVCnO6l7UR/ZfQagQqJ7oKscORWpjsEE8OIpWOWIwwZIoaFrX00T1H
RMjOa7LRX8W72y8d53Y8zbUT9G9Pk9JGbCsH6ZOYXOXnPPEfTUrs/MK5KjKGJHLWFzFyR12vtiZH
0oWxrIk/UkadWKiEBb2/UMh3mB3gUEcndQ4irYz8N505kU1Mkpeb0IaRDdnMg/oFlKlSGKknr/Mi
JqQt+hFxwT+phpEnFTYIbE/75U1bKjknz+Yv3YN24vhJYW9Eow5Z7QNHo7ETJyrlXKnZbOyblK03
Mik7fW+DNFSf6tr3zywqVC03j1Z2IThYXuOGYkBjnY2X8XL1hz22adTjTfGLrwvBDPb7tO9Oe+Aj
usr31YTOKf/NwLOXYre7s52eWcKFcR98gU5no8TluIJp+DKB3rv2sNnM0r6mUpPXrUBUr9Nwq5Uz
P3cmQwoPseI/pqTWN517fdFQvQDGBY4qk8/F1UO178b273Gt7AlursdKewmb2LssDE+jj3hX60pL
FyF2/yDQDNqNRt73kOpHjUVqkG3Nz+otuFZ+m++QFdvhVx5I/j6934cfyHwWCxQ8VgHx28tWPLuN
FmtmYQdnSQsxNCRwN9LmE4k3NlbqAt0LbcBzSfRlfPEwrYhgwk5aFfDW7TSe+Yrpy77xFs0b0e2K
w9f6CUsrwLglHdLEqj9HcvwB0FdaoG4xKhFRucb8qs5XwsqqUVP7OA2S295XibB+tgjdXL0V8N+9
ndRvpWyB5V7n9hNgEnfRKXPpFhB9y55pFPylaPofU7UHAPTRCUP7ZLpNwnexa/G0+GodiYvlK7Va
XAbaXXNA7T79zYpoghqlnvYG5r65TRzOtgsdxuWnlhUPLM/DzG2zbr0cdaGbbuylgZhjklLGy1ps
nq4cmryrP6Qslz14sBMtfkGkarzDxaGr0Q6qY8vAEdJ5XFmRlwU3VNb5E/58sbC2MwSaWCCru+Tu
obvt6Au2ffbL3+6mRjDudEJEkd/WOICHh2fDoraKNAH9lv4CU5H7i+YhbdKQDEGX9GA1dY6172Ua
F23H7hxAJSfob6LnClqHHK4Ic/4Vg42Aj2kx9U54tx9lZj47py3EeNA4bW42Lirq7Y1dfRdpIOwt
+X/MVRPKF1X81786EsL/yfB2DhBDRzF+7pht97Npo0yMO6fBj1E7+mJvYGcdHDnvEltFF4wJ7l+4
NUrfp6nRtcg3tLaKZCxdn5oHBSSHmn8STUng3hcoIzaAUKwYUnJhyDxJry/gKvYiKFyQ7kOBRo+8
3bq72ZcbJWITDqLWleYcZHgaSpNw3qkot6fZif3DFf3DSKYT+IWVdagy1RYzGFpNa6cB5sUGMI00
fADPqO2aA2Glfk7H0OK3naU+2YRuDWL0KMWNazCmNwSZYKLkUvcSVrQqfAgCVCebFZI+0d5xoxFY
ahinoutwWdOy1082ig+jx8hGzQZFzBMrXI9sX9bcUWnPodjeNwPxO9jJUi0tKB7zbS3jOq2bQO+G
9OGFKydlKMayLsXpJCu5bRevSRk7u0uPqZRoEJmLM11RXUDi0JpjBIoinQDzs0FAFvewQZzH7+qQ
/JwOiu3PkOw+fZAcVi3NE3LL/eiwPrY32a4VIPq7NRf+kIHa5QrWU3ont2eKUS/dYQUsW9M4YjUw
2N6VeJGbwJbwem0pyWUJ4Wlxs8w5v0hIUFs1NFOtZ56B/6Gi8BRU+b3ujIExv+FqrmNIzrWyLo6e
LPAr7KI7U1xhp8kMbw47F7UZBYPYSjwXIPkwYEEUUxTQUk9vdyo1+MXd88GfeJ1Hnp9kScGBi3xu
ni7cT4eNqwp+jJM7Vf0yST7WwLBJmy9TaRn/LaKCoxFh+1cDWVdybIGXeb7OLKWnJ6SbUBzpyD1N
QddSwQ8MDtIZWZXBDxUof+4fhCOdLmjohyASrfZyNYSRUzwJ1ep9ajijlQARmYMfQT9eLjiLhOSe
EAJeGRnv6TLACDs8pyCmHxyeI5PLwMtUgob3C3ktRrMkhVpen+wLQc0RWngItXwbBKRI5WriQsev
KAEHDUV5z/UuVZ9eeuJLmi0yQ8eP4WZwV22gZtWnw0mUa3uWrRbgw+c9f+1q8t640QbiUN1RrYFE
7dOXqvFYRzhaf7vqjJzMShap00Sfb5AYqFBHumnN/87xQXZelk11RR4dhOOYR02j4Rbmnewd0/GP
zJR4vLnh0VPEDBw7viS5gDZRNRNRTE11A4ki3Zi68a7sxh8/6w1IA4/ADc6wYkhjHHJzZrpCFsuP
cT0Lm2nLmpKC3f9L7vlWe4thX3h1LOvsSkQ2hQlNajMFg5uGVcOpc6eCfNsLSybzPYP3iTxSgAZk
fuVDf7moW2kU9IWlVU7Xr5Bp9Sis1ZTxK3PJThW38wxS3qnQZF3UidPrxY9upoWWtvHXPmq0dCEY
KBSKmGjHQx+4qSNfgG1OVdGxMHSAyYXJ6/Hq5Eh+MGJyp2fJtkO//AaiFZKO8PBOiOPzbRmdMf2b
B/v7/5Q7Gxnsf8fhrRK/7DTIpHY+F4FEkK2nDtJM2bss0F9i/1U0z8UOwNBBXM1NKe6L0ay9s0/l
S5F4jX4+fzfrru2Tom/3BmCVpo+XRfeOdvDjijYSn588uULS3uC4KNBJqMXeXwdPVykjOIDPnzqh
xW/9nTw0yhQV7XXWXUFKHUIz0QNt4Znl8PRkBvP03hofFQdyp4CiCSNLlFODp3ka2pnMJfn6xyn8
VLYBg7mx6GQwDO2MmXLLYUiErDtfwlAwxqs7R5wfK0VsFkf0jHJJdUrD8fCOyBM3n87BhFiJBT3A
1gHaY59Mzs5dNl/YdPMJLwuzYb3ir73Y3ViWLz0FMoSX1BB2n9MiIt8ajSOOBgtZob37qiBXSKUK
7QgHzb2MxnlPH7WihCXEbXkaKXbaDyCs7Cq0xL24+JIefRsZGk3KkvirpotprXNQa35ey3/kIAvS
PhDIM+CSlEHKop317ftxNlCFhr43dvPXf1ao9mIsZhqJcemjuNfF9ClWcyGJik2H/wmbQkFuwPge
3ViUlqelKvHcsnCc+kZa0Fk+elkq7C7qQnh7F+qtKt1NBpaMoNRtrNT6VPHV94coYO99zaKd2PJt
2zpW0vuKRagx5ewyUVzIQGg6aJxw/tEHiDZQBuAsZDNEf+0AqAPSptlY2s0lAO+WJOmxnXo6sX42
IWbJ41csC9tTnyB7sU1XKjKX4bXSUx+qqlziExCb14gIQGzhaGp26anJPjLPqnbbMph2cvU9bjQp
muppoSXkKZiITf7+OEs726AsHhV6GvVKuIwhi84/4B8bijUB47OMCXKv2sIjhcjScyNfNwh5dSzi
eqzPvydDOC54tit7ziFjbE0K3kBi9+2YIljYiM0MeYafl2g0h2TsabnEWSkB2fjmP2xupNBy/VX1
0p4san5MB2LlGr1LjTx1AmSVoFbcebb31aKm9ZtcayRwrJOqAtP66BPsfgJNJy8RI9dL86ZFJbJv
gafj2niNYnxYS4sHSz89yfkA+I1ZKX8C9s5jjp+wdoHAHjR5XMeb81ujKN+IvMNDrCSO2zzCAkeS
n2Dcy1zWxRSRfaS86BR1wO0GiZWUCFJGGkGYREHCpYh7Qn6jpxPVF8xRvpMCmgtyYxR6tIOj1+mH
XccwT3ikl17+SPMOR+mBpcVyt1xSVDmjpMnYKOln9wK5B7HnCFKbqB2jqx7pDnOqR5EDVnk5jHVq
VZGD87AomRGC9/WtgUGJc5qChaTpqaXxNW5mGrF0BUuxjXnKGdYa4FkKKRZSJ8PAzAVjPX390yp/
o/6JWoNju5ESAlCnYHutQQ5Lc0fAwFVFD8ISerN4/843ZrZDEZpGaT3KuSsGPhcbi4rVRfM/phI+
w2elt0HxGq+mv5b9qWtoEE5BrE4d1EBR+1MBx6LirkPPrjLwj6YCKG3b8jeIPdu3OKbO2S1I5Sbg
0ZrwyehqD33hHER9Haep0h5uPyf2u0jqPMQFhngr3FPnmrnPw/uGtWf85zOfuw7xt0XO/V0sDbCa
DA1PdSAaQtq/8LO7s0zf2TiOB/nNKE8sO0DPG2/zqxIsDQ+SHkvHVk7dyNCp8tokrz18qaS7x/hh
R8EDFqm3a9g8sg4YT8Qd8/25tN9k5GnZe9CaDFOGwQLEQvgv60bHb+4dKtiy8cpEpxyTiVb6Gl5Q
adRCVjnZh3TRTar9+rHcJ30ldRK0pX8JPAJd5Xbp3LBlWWdHVA6zbct1Lb+gV+ZD1J0pPjO/gbGZ
d5MW8UfjAsYmOhfiZdsYm8NSDwbRZeFffSFGxFwrVEB1bEL6uMK/a+gMON5AYJfpJHYQhv2l/IeC
mT0GJT46sH6hy8cIHp5vF9S/pokh6GsXY1gDQAH8lbny8SjMgCbZhsyRqBB8mnVcif3VaHkag1c+
851EzAte06wUI4HD8hN68OBUjU9yvWpr+DePnXVdvUMI8QJ1pxovqBvJ4KsN/pnZW4rhpI79hyLm
8usW7M+dstzTJ+l3OmgZ5Y9XWyKwz6Xw3JX4B3UPyOFw/iV7ye9T14igzmY1cs/gj03Xg6ZeMCJv
6jMbfpLQKZxxZPUp+s83bb5Qg0T0JYxTRz8fWtwlluXi5lPPM2LIBEcyk7CTBJ1/XwJzoj/Eljwx
tpovjASx27tUcdJYm5kcDFUaWjd0bh7ZbIFVLIqqUXISOPORvIUvxC+2gCUceH+C12HHLxGWBYk9
IK0PsOzX5hK2LvC3BFho1iM0Whe0D6aATD6TwWLE/q9XUM0CZHok8LHA8GNnZRFUez43c3FfSGuj
pF22b6kI9KL9q2mnR5IQjyyFQZIIzs/B1mcGf4oB1VFptLAJcfJSMpvm1kSFFaXnzw41BRK56+Ni
8cH6mwOXApMqNwfD1nRYbleGjTn7AvedTDLzwlyQWzLA8P+61sbuuBDz5csqIDquTDWWL74nCugb
SG6i+cNIWzfrwHWlbghTiRV1GYufU1LhXmxiiDoTK2D4nTaxFkYAotjdyYs68QB8a+z+oDtmVm3G
kcTTaxS7GJzYqwMYz94bONm9kRABzQe6BzGhvUuiEcKSGAGHmjVZFi6E2OJZ4/rdBF9VV8INw9Vu
Frqj9Wt54W8EgxOurtZdARKHPL31exaFImIErCLjimOXtSHiHu+8YJf9tGv+lVNcEpXbMb60TSR2
C6MoDB/zPIy+ZmAmCK9ymIbfqhVm8uO9YsAWvH4oKocirkXjR1QMKCf9/nM0XGYlTHM+BsbXmokD
zcQVssAeYIgsiQuNK1AmlMCzvFdoI38tuCDO4PTmp5UKo2RNG6c9P5WQxG3G3KaQxuvK7EcLFHnZ
vyGUlweuYRAN0PhZj3z8q2J0dE08CGxN+TA4KNym/X5gVcTHuocNId1BXKFfReXY9uoPRmm4dHQ1
iGWaL3h0+GR0Meng4qfo8m0lXUW4booA5kL0QRC1YkU/ZMIxHqWhxHGcJDnHdwiU0gKjciPIw9ld
TYis/C47JfBoe44gNB/FjcZl57WlUh0eJsfslDMuoxdVDqQM5Y/71YH3ujgMFnNDPRp3Tuavw2Tk
YGnbkApDnYMPEHYQ12zp4TCbJt9bBSQbrJzI4SQyYz4ycEHxuVv5yT0o4AqS88hnEdBtOOQdRAt1
+QnWoPK1tmmVK2vndxEbVMS4NsfDAvLViFFUpvO9kJ2+Ly9cBDecv00ziIJEqJuf7tIcyon8EGfS
YY+a+L0N7G4oAUs41CHzMracRVakiA2X7d08CPwNM7EfQe0tad41Imd/uQA14GrWym3xOA1VNE5B
5xi3ZObd3tUiwHA53yhl8YnNyij8cHP+x3XnWIbHyYl6skRAbYd4mxRT/ik4Bmx/iXq2Jt/BqWBN
rvyf5DOCWdYylseiuN5l4d9vVmBWOiS8YcgQ1UgTaxhIxjJIFpr96Qf/qhQYefb1IpqBYTLgsGHC
53Ibkg38ISLiBR7kbS0I6FdX45GXVKx3np4Vp+9WMK5EXgkG/zLYOeXX6Cr7uvqxwWp01CHDbmmW
psUMZWJ8iPUjHm/aeXdCZpFe9Je//IcpgUDKDyOEeUX76f6oU3K+s02jm60Ty8ed/XU5XhQBkYHD
6YkhjkEv2iuNvBvdjldo5JVNyaUOYKOO82xd//+AcRkUixpXxwu8T8x9mBaENxemby8GDNmv3Kq/
q0H1UFcV+AMSc1wJaV9lr+jABOO4lpiae0GENhO3EsCQyCwdmux2FH+XMDSXTq2v8OQUjOMSJADe
q42Q4bfw7uDgHS6fotmiNJkE1Vr/yJXpX2fMb+DzlIhPDKwBsAWg3X/MMYAR19BF2FuCS6oxKDGM
qnreMJxuru0UMKJYu9lHubhdJqz/hgSL0lJB/TlyzUDxa/CMcUA1U/CfjZHYaqnXRBJOuEYKKav0
I+qhv+AzsbQtF/d/tbwXyk7kInVnYWFlBIJgmOWfyLia92i46ubaOoxc4kdre4gr5N4wqFXmw/6C
N0B5ZrmRf02Uv/2bt1h4/Ob5kLmCaSoRyMyb9kGAd4hVDRxHXD1s8rnF55sJRxDruoDVwNNhSK6+
Z/Nl5D9cZKIa965ScHzT2AxAUahvfrWQWp/Eq0BiDQfOugQH9diqBTaMo2RWPnZz/tb9TZg97Ln7
hqND0IUFMAHRtznzCw4KE+vgDGyVZVGuUh0cLB91lpDn0iQ/aq2RbAlrFEQfeD/PlVPN5LVT+5gA
XGZN1LBJCV9s4Vo0/XcOsZLTHOnG2JrfxC/0BO11rq27wW9l9M/gVxDWdGE0zn7euGD24fgJB78L
41pbTiiQeqmlbA+c4Z9jb9UihrwEQeVCIhYigORpcPvYSu1qmTVyT9vY+mOewjD4d8m6yXS0GoVC
B/aroGJhGeYPhqqMs1lF9Cfmedmhl+py77k+rPPtI4ZKbvTddTOP3JIUJKOPh3o5RWv6Wlb03Bby
UjoEm61pizMlQboG4N41IymBG9Z7A5NlLEuasNOO9xexc2F2CGF3EJgKeavfniCSjiV9W1vrKuOL
NKt8FZQrg9xSd/VPtA0MKt4SwA/z8k9nNh38h3q0tpi6z9bPEOAjnks6jlP6WB8Bib6wa9ZaK1NC
OqHohpVsbbFEOJ0TDYIwWHrBBo+B+6wB6fl4KFF24beOaSbOodD/yoqjlu5oyCuSdg7Rfmq9iyQ4
HRUfeym/yreCi+FjWrtsnWbhBxayV0VlQbmHYWv3LaMwBBPXtp1x8avzEd3cg3HqAM/zMTaiZlfd
Rf2eMxXqJAKAK1yGhz6ygUr80bnryHWVJY3MfFr52kz0m9Xd4vum6LpeiswEDsRzAIWEseXjEecx
evt/SBPx/7O51BAFsiJn+JtODjAuTodtqhI938K5yZ0fY8rMskK+BsCfKkr6ATY0lL8MLlYU0LxN
Yk1r1uKQCkT8uv+mgv2A6CzyhAKHCkQWEoZ7cmxxi3NnWNvu+eqkXGjVs/8f9yA2JP/wHPBh5yW0
2cDHiPxLcHQegFBYX94D3CxIfIKe8GA1TGEgSbzq9/bJk5JcEvNA0GgyHUCnXcwivzxasKVCzhKO
67n6age8mPYNJaeGZB2rQDmGnP9fm2MMCwHhqe+0RfSEzHQ9r5mqeB9KaqJG3PMiqXMJaDSNvWj1
IZ5stJk+1c2IrWMiKuTCVoEtIFQ4CPpIMOzrzcKz0UAnFaqTMgeKpSqmt8BBNjz0i96VbxWkHaJj
nVtkQImQB7FcYTwBsaNMcwiu7it29VcZyYqZy2MQ/S6ETcdS2AkEG1SKz2+LUZXDuaHB7uUbahz3
erAoMv5iHmTtrKWNW5K7LfR3u8J9OR/Vv7BvPHKHUgmXASw/BbymYaBeL+SnKMgkMDN0UKmiu0OZ
0z5JXnNxD/4FI4AM6gL+ZbUy1xGhHjorw/6/dcqM35SHMz9/UyWMLOFRay1KRYNVqFSy6F5V6n3Q
+21iw7XZwLOCxsJ7HJ8H/uff+n3/TSzvQ4Kqm4QEwXb5rSo3UgtqHI4fkM7Al5qrmBlpsVzyC9+5
haf0CHLrgP72UX22dj2hRQHGTOATGGf2PeLrlGmDuOt/HibSPnWaL9tYUoHbu3s0+tABV7A8h0D+
RSo6jCELpbgIGNmWRSIX3RAmBrRC5w+PAtLT8XdpLiTe6IMNXzFGOK6GjJSSrkMHfi+3D+H0cS/X
IWDrWlqhwpHvIOveEhSZPPsy/llxrvI+QWGY9LRpsQR64lV2nTEU93yHTuuwUpxl5pzvXym6nD25
BEmPIO0udcrxcBaacwm98w5GMxuoq1eFKekP3bsvMOLz+eNAl/mhL16bX9BEvPx3DdhPiFKUtT3d
3iqKmQ2ubSvVuZwhpsj3wJqdIJZec6cNQtpQIj7udpISBLMrFhBckKe9M62l8/sPlXFilwruTz1L
gdet1Oc8d8Ud/x52vprqujK659XYaHgdq6JVLG8g8t1ZiA+tDPD8MECf/IlfQdU7+fviI+qlpECd
nvCNk2NcW3GxyG2PxTXOw8DIPB5/sAGy+CvuHx7PvayDuKmpafAs1kb6RUQWTyQQlInxBujWWH3q
d6Fre7v3fSSbSHy0Tb2SFIs9lKnUwR7uCAmhUEYmvjunV1aHK1KvGo1Id6lus7DSROUp2080QECk
o1XokvQ9UARIIO6Qq9QUubbdJeMKdNf3w05/DilCWddMZC5gdQKtZ2PWExHnquqvj7aNg97Hf9xe
tD/bqKws8KnYW8inc2Hwr310O7q8O6FFk80SJHMFrWuwGgxNl41dAUd/r9x+iSWMkTHWakLOq00N
p4ZHCfckyH5VFh10MrsL64emRrdqsg6eVcccBH8XTDCzLbie6rINiSQCdqdoDkyYYjt7eA6a+INi
/h5O1rHBu2Sd167ZaJTN8gBrr2j384D31JBj/tMBZ43K5esjO7L5eCLtxbAQ//7sagbRSqRIoTb3
1+n61lvnw2qp79bXBGAqAUWeVAIh9OFHqcCyp8HBIUdm1JhLRWh1S2dV5J1PJkFxfP2BEFjYfHZ8
8JrdEnWx+fruE9DoOI2Za7qbNrAZUBa4ZS2ecph3u87fNlai4T598mNsuqZ/rTWUr9WJOGyDAEQ5
ZVTzEybNUY/uHd002uhqQbD+zTtAILrKTJcsZDVK0aRyq+KlpTkN8MH9319vaSWZVSTtivMS5I2O
MfhLKaHkPlZDYAV+msWVl7uzGNa2Qb07xJSiKyOqScDcRK0D8bAo0x69rQmy3etIuiXXZyO8fwtu
fa5AqF+If6gwohL8WUW7JpIaF4Idr/CKqaStlO2xjSuRi0WebmKJApOpJ+aBWt7RfZ8EpFDQKHia
OCsL8J3IzqgNn5F5NdJAdhTFUWPpzFwgp6iF0/4nWzwddPWhsztmuksTUfJnW4UPCFF+tevPLZw0
FnCz/qku4gGkwfrwSAx8W+ZAb9Ysf/nHdJzPIWJZ6XkA1OxQEcokdvJuxMD4NrzwuB6gPu4iwiZa
F8+E3V3htGtNXbLL4mMnWShTyOTG2J/Xr7C9IIJRS2rKmfI0/Ms8tFMLLs0Y6wKOwdXoGaSoWdPr
gC03KYpJIViTw/jwKUz6wOoaKyh9CGq4Zhf7NpEk7GxzkTYYLnnc+VL5m+FMO0V5Vujg30XhQy4K
T8UV6Oqr3p/7TQq89949A5Fous1gZS/vXjCYoYmgIY4omY55Zr/KAnEP/pVNx6YDKnmXt0e5oBg1
8OMdaCmLy9vMavtRKpDCcLxZCqGJe7AfcdCpLjJ+Di9rT68AxB+17LM03a+HTR0CuC7rLPFbDr7C
oGQs9qQEfU+l0Z75rCo4Fpjr3L7W5CuBQ8IH1m3niP+VqDqEZaHBDRg+pzZ05f5/k/MAXD9DAW4d
CCNFRDqdTgdhmpNyCRB0zyXZnHCfAti6XDnVAJCCdp9tSmTw9YIRhSH+tB7lKvCBimekYi6xiVZm
gD5HAb9nCCJ00g2d/ajC8NrVQWxhCxQ5fSGGLnrtWEaNxpuH+yRU78STTAmYhGtgDF2pTBn6R0RY
U03wzTmAZ5Cdky7ROWOcSER5xm9/qdaHNK4L8KtbwL7srpXap7nC6KCqdVg5pN7I9z05j7gMRcoq
eQekRYVPLTTLV6jLzg0VzeQtSuBwYrsyyd8MDMqE9HsbPDXpo+e42feLKIBBQChJ2BcMsCvMAk6N
DiJjSCF9xzOUbVseCMk2vxHQbsg58yB1dwTEfZZFQHILzeVxDutX4DfX9sAbepqFIBSRugkPk3Di
coR0fhhz1IMFEIsC8SrbiU7ziha+/ogGnVSt3+wxtANTQOjCZmV5TpdSq3FCiQPo3EpqAI+QDnAG
t5rPVLvsXHRA8oLXT7p1tuYKxcv6xbWw94Q9Yk6DbO7z9Bu6rZ8gQ6WncbFnlYulj56XGpXO7yCp
pFEl8rM+BGrltYBn+6DKmUQjBlw0VkLkAtKGVPOAyxBQZY+B109HtCBGBDXn8XXO23JdI40sINqd
hfQwSzXx2iJ2fdBIwPIsj/5u6SE/8kh1bhx4mRqPe9VyFkavG6zAqyJtDjWJ/gAeYgl6l+7eDyJH
CJAfRa1DyduAHGvDx0s2N9oX27r/2cnwsvIQEqr4/OGxMaT92zHxENr2FlbwGnMoDxVmfx47N6C7
djlGr/Q7tp6uKId07O89ADtMwZNGqUbZ9QWD11YPLTUmQKS/5CPx8nJUEdphuNk2tinNBWNWAPJZ
Lww5soec76w1XUnyiucSN1NVZHxMjC/4vujIWoMnQbq1DFebbNccNzJUk5TY2/1Hyhm52Hdis+oA
1qzWWnIyW1uZbFEakATI8/uZTbONe9MSSF2eqt87z5/36p7pVQBpvXLwtTXKJLWtlYJr0Jd/TIY4
DZUSsQhKZqRGzZ9bkp+vzGo7KS2EC6oWIvmH3sM7f3yAiBzcmS5kobGkLRX2jbs+Y/cenz42AlsD
9UWDXI6RbJ83IplexGcFfFVPP8H8MYgo9ORzMkoCTFcw0vq0AZaTw28dqD/Kk5LDxgMiv/niVr74
GX0HjfaX1t5/wOawP2acnPmL7GFrnJJWDhwzrMJGWT3D3HXVuNI0Cnq/qPEF8EJQQguE6R2ItciC
yMi4jovvggd186DouZcv24P7ZZjjw554YQAit4bNxx3Fbz0DbbmmJccV5qOXGceHf+Dl02KCMvgV
Sqj8Z9UFzvKyqNiciI8W9Seyi3sHLw74kEH+o0p4G0WhFVgG4OdJEEt4voCVSs0JYc/n7wLi+eu8
8tzOViowTPAVSs82/POf5/+VuQljCwmzJZR1MfkZ/UJSc4Rk15akyIQsM958LfONGQuN0uMDcMhu
m4UDjBS1RwDvmrIgzqUEyxElemV55S3mk9z1IzFDeA5INZhR+tkxJoVN39WyiviJ5en99zDTeTGb
MyndEnPvQ9zKo/mTicLv/5aFyetalb+Y4d55EAL9mx9rW1Ms9JwOdfy0ynAbgfVxPkjL8+GuXK19
PL4G8bRsnHztXTK7tIefkhj/ffoZgLCR51yBHqtHjf5DsxtRCTxX+xxMuM5Zd/YwwGYxOuPIMjsq
fEdLDaibP3WhgEUqf0Md31M+LCmxjLrXpPTzBlfbODjDY8OxMyGBosXViRi9YGpsmzXWDep1cMhn
OyK12ao4ECYNuH45PWdFsg3qXBQ7wgf2Iu2gJDWDzBS5aM4cWs1CsTQYZS2jZiA7+2nsQTlDBweK
jAbArmnMf1hYIGuskpJ/hgvNlflHI3rLQBxOKX8eutn6CbaOKytBuTFsWmjx3oKiVWzAA/LE9hNK
xnudN+Qs3R89hE8Y8S5UF127vJQBA5naaWlaCYeZPLTkNIGb+rS51jJBTa5hbjvMUZ2xjNYt+ndY
s17zx+ReWHhVuic1iMEO/cBzB7vUpsQuBX7wEyYI1fMJZzoyWs9MCvW09JVAgqXes/a7j6dthDQ9
XK69w5ClwFIh/sCSd0Jlm4H4KctYF2av7LBzk1uzOoE5VRwMca8Wq53VqQAK7Sv5rEACwbIhgTr1
hXZPjVk2RRE4A2tXpOwQcibxo8ovo+zC3udUBJ2HXRF5QJmPpnuIFbLezYpYnDMpKHRFwQLfyfo0
IEvUq8xER14KumvGC9U3Zhthigyi+C9tYMKBhZwOXD2y0VGbUOc1W8vj+G5DHXsIvu/NgsuB0i9+
iqbGd96Q3JrEFdXwzkEkrv4l0A8Rx22ZQBgh3L55wK5gN7HIAP1TNnIU9DffAzSuFHNtuLCkr9r4
R6jfrfKx/gNccNvJv3Tin4LI7au6GtXyOuj4YDYvVL+6wNXMZbkasZ/A0FVgzCpE3vZTczHI7hgT
VDZTTwsyq3Sb3QDJM1O1EbAcvSxX8g5KqoECODU+muGw+PJTiiysjhQwhuKPzGlJ4CTRKNZ06Cky
WTf0go7Ba35jY25UEu6lR5xyqBUjAK20Wso3nSYre8Q1LhPO0XCsONjpjQ5VEyChFv9seTeDdcGY
b4y5DMeJAKUreVCJ8ZDmHokX5vPJpk+4wgCWbl3gAWgoCICGWGoXAODmXC2N8TXt/3cjvZkNOTWG
GqtMpdiGQbCYJunQBZbibM6mbmRNUyiwpZibnnAbvHIBkanmaTlIbUYT/DdmPAHDnmD/BQwwJwDR
A2T01oLWKVxMLLXjKjqqvjFP+n7NpOES34kGTghfIIoRMojCnZgtW5WtZNEPh+aqmYhGqbPfbymj
tRgp/2L59kr233djnuGRwpxPKRHGq5md3x2tGuUt+URY7NtBgUraJLYTO/vKA4GoGPXLM016mO3D
CO0W65RyAtjSYx2wbtz5dVtsdn5fHlGqfq8IQWD1Q7sPltp4h5FQMNeg7juhLUn1WDEivz0ROUxh
hkwqTdDoETAEFPhV81fr/TjxAjAU1ftzVvtxAC3bWtvDmX9KsEi8kMXuUOOG5i6SKwOU9Lz35914
CHFslYnWI6f7vRIXrHuwprFT4QgFLXBv/UgAggFlkGICWl0nF5o+U4HFkHEGXqXLkPqCoJ3Tx1k7
hgGPAk6HACbEF8g1ROgGhrPnZJew8cCM9GbQ6yAP5SxJH8HI5+Qzqc6qRsyFI33umuWYLPu6zbLm
kHNW4w8Qxdj5zFPi4ky6bMXLcvOxVbODjbfCbiBRiul1SVh5l6zzPIrAyzGspH/h65Y58cpbR704
P1H+DdxsePmV5+cNeNS7n1OrMQu40qJDrCRyDG1eCsfYfYFCLCF2YXdNEf8mOq+DIWP5svPh1IeK
l5ZBx8P5Wo8apP2/aFeLtlpQjURM7YeN/2AldYdU1w13rXjAPCcOt3C8nUQT/6kh+8fB+Q3iTSkB
E86w+6wLmkDZbDbKXWDGRm0JC7ju2ycV1vN2J3UY5PPiIJqPr0yr0uU44NxyIGb1XYpdc2m/1J7/
lqwm1PObwMLwf0jLt6AGeEqaK6F2jVeMZmSANWFPQvMLOsTLnRL62t9IviooJuO0KU3f0A3Zinod
yz6je3eJSO+mfncMkOxDC3aOzx255VHv7dXndgKJx6bhzk0lUMhYNzzMqk9jSCNpqixxcVkmeC3k
i5KOb5FlI9qudP4ggI9SQmVvPycA5nZAJQTI/48OfuZaA0f1kw1LT3RN47QxUVlul+Aa1ERaIxzX
lM2KRM0qypaglJAM59RhiWFK9iU1TTINXpkXnEL6k5iN+ei02NwgMGFVebB0mWl8AwGuGsqPKGdU
kAPPowDqG8U7kX6nks7ttS7XTq2MhVrYOGb0YvPrf/L0CB5CG1NK5FwjMFMNs1Hz1VUfsiUhKMNr
3vv6ezsGvKtFLw6lRy0OKV5xdLB5zewxP9j9scpLIf3XrKOMJ1QuqrFgqDqhxzh2wVNepaj89dpx
OdqJvO2Ceg8aSia95Stv+hGpVxnyQCt+Oau+/pAJnknvlcc1Yr9r9L0YiKYQ99jWGiQM3lgsb+3T
nc20GVAeibFlVtHEtSv3GrpInCDaqLEWm9oHtw/HZi8K8qdZLLHhujWNoofM5g2QJy3NvtC1/4iu
OF/Nq3OjbknDeE4QHaHXBiqq0LjVkb+MD0CeBWaqJY1UJUgc8I90gkwQl7x1QFLOhtX/phmkpk3h
FKb8A6BX4LmW9OOrnyqnIRADWeA3AX0bfAVXE6HSj+MfROCkBWCaCv5cTgam+MGdZiwn20kgXKqM
vDVRRaO5ZUnWIoJVA1Bg8kyVdoiNCLV1C44Nvd/J3UbM8lz67Av+Jqr/nO0QezMlPBWXHsaXo8//
hbxvdWJWhKYQpcU8qvmWbjuTYOOe1FRvHKaP8tUgcjgsDftvCBgglyLNhH+rret71ypMpi0LDZnN
Wxf38KRmTRkfJwJ1qg5/xqN1rPl5AqmgaT9Uw4k78I029dg+Xilsub8SAGhA3i7/0NCDFffUlbXf
+PinYjJmKHafuoRXnmmk+LE8/EheqX8RyGTK2oEQ1wSlDqQD2RaqOFDO524i/wtbbATR195vrCe8
kpHBxF53S1R0hHwm+MogioZAjaUQzgxZeYDyEdVU2hMwont8sALMWV7UJGtlfUCbV4VuBilzYseD
YPIA8JEGmtxTSHMSWPv44x74Wv9WSdg6/HUJWtkcFEjfvI7tzfQQI85RVNSKAAXvCkmFnM4B1WS+
3kOFuiVjGxpVvcrqmsYtvwnkPam5rmz9sNv//d2CGM58o3tVI7riuS99gIfJYDkv+rfVglG7MPiv
tzmNeULkY+ONoI7B6oGRvBWn25HaHFZtzsIxNBz7bc0Dq1PxJ3EFCHWNXSM4hi0E3J9ijOT17Kbl
TBVZtozrvYzMKFMtplVDSzifyal48QwiPemuW3yMSoK04vsbzm/W189gyC7PmLHhRAlegEw8HUVS
wyRFLwqaP8wuW9LuyDjvuLccbv3cCU41jOgs3BfAYIt0Bi6r9FbBq64xzcIZpEjx0XLtzYNnwua5
Jr6l1YQzN0LIkjWNRGFMqM4v6+PODwteIbiRvNtvWlGckBrk4sV8c11EEt/6rm/a15RfnXk12vug
qUKu+BiHMGAF1U+sEYZm8tsSmWxDKK+ro0WuSYANYDR2l2kN5HnSaFFVs3lda8hAmedKQ7sJNV3t
h4+cpG66AOx59wfiPCWtmOoIjQx4DpisEspFYuortc0b+XwBjAN1zkosZ+XsLamIcJbMePA1KSRd
4PrrpcwC405AR/DrI9071/PVtd+Pg1zOLVHWsG4iTz3ds4rlgVuYIhSqbw08m0hOldxclyUDLGTP
BdUziNv5LPOI3AEtyoAKXFIrFe/lLo7kthkt71YrpQCzFEAzPoOp5+c2Bnb8hinfmPZXD6A8gQTp
Oo4QPBZlqgvDcVcdbR1CWTte/PUrDLrMJX2ntDp3Eq5Ehkbnqeo/o+X/aHrV6z1QPP1ijN2w/r+P
3aGMvGGZln9ToDjtoZ/25VWDfLSRXTAFPX7Wz2n7sRF2D+CUMKmD2FXNp2S+MO5+qTcGsVOuH11H
XT1MLsx4Frodr5VsHrgo3moprvVATOxbb6cGkPXVkDgTZxD0iHm0d//qTZbpk/m4PSmNj0yixCSa
JYW1maXEFENhi9Y81atwmIXM39UcK2s2lI9+Hm8ogT6CYs5nZ7AwAHpvm8kxy1vU1MuFqdnWMD8M
LYsLXtygeoHT7oI3CHb8S5B4DG9M1NpZzk/80UrY1R4FCovQFqzr/SSzwYR181v1vioWzvt+QVIp
a2vTdFrTwaiCryBYZpFLl7VrEgPMTLHJKFxzzaSDJJrAJ+295ptRNaxYgRibYLrqz/3hitPREknH
7THVFL2SQ0GAMblWA2uVMhkswDSHuDGS0cN6PmlUf/l9fwRNGsi9aRbKYhnJTexbjAT65XGYT2mV
V7q5PLF+uuAqTSmXa+ObRJ5Sk811a2PJuW6MI069NHLynuB9FocdUdiVsnRFfvn53fL2t38BR1q+
sZ2C1ARhVOinjR6e9eh7EkFtI8E3zaPWIafozYqGyYXgFDOuM83hK/dKUboezacYnVSahb0YK7nU
2clOHty1m53CBm1J02udhZtEVOpD3TdfXSTl5llee2+v8BgmDYUeL7WQFIS8eQIqaOj4BwPOkFiZ
RRoDw0NMBVTJubWDeMGYTCpTIc1AOGGOpZAwpPKbYkHVOXDrsKgISnJa+yrHZUmZehqa7eKAr+MX
vAt4ugXCRvulMPrNTndZcCSyBNnHEy5khZVHiXx5AX9sBh7HC/F12mksvFqrPETLnU/bDqxukCnZ
GdAbbRC7tnSKcJyAfPIhQetgwe4mEfaChvNUheVLVL5JVdTonj2TelgoHSUf5A9oEye6Ij38UwZC
+OMQsPi5f4Udz3XYI8g/pZVw8MnPJgiJiOHzPCGmoxt7RdxeJZL3Y1iDf/7VsHg1c3ig5lGBjn4F
owkJ0RtoAxUu5y3fISAnNs2/MDGG2vLBEDXDmCSuAXKUMMnmC5WvdpjdV7X12OfVF50EzezVvKRf
GaJpfgMjpW/uXm5OaN4mgQUzYuzBJy23BK2Trhf43x3psoC4vjMOhG9CMomLwrlbrmg/QjneNSDM
uoUizBos8GyKK9wwoYQTQpF2HbDhKzJ5Kf/MBpCw4WEQPxuB8lPo9BP/MC7gJ5yvdYZ8aUuoLRiV
ZNPTiZUyWk76j2EkmM3krjQ8k+bfWgsDjD7uSMw7EL6XEbYF6NJAnumkQQVga9NEa/GibYsNE4uj
nv5u7W5NgDGe7Gf6xwCdgC64P3wTEPlcrTkzU8DUYl/eCA1ACXLW7srw3njdGQvJroWRoUw3AdOI
TdDFj0zZvs+3nmurUvMEFLCafIHJdurz/Mb6cakqXNcieMUUKvS+fOhSWIqEzUz5w9Z+wSyuhcQu
rssMAJFxMRnucPGert0lcJDi7hbun4xXnyKw+TCcXIzNKDXeM3/aY8sG1ZIbkXazvlzUoGoQEsh0
pUi8axGs3PPutP5UTSBcz/obb2hJUM2vOUFhgXBpHPBAVpL04ldyicjGWB8ftVJH424PKANzzdYk
sl7+eBSxS3R9ygUX1OeGamXP1VFh63WpEP3jYIvtuQ0KA2yKey+SNRreDy5aaqW5LsiE5c4jA9lP
97DUYqJUc11m7LNNFZDGADrNX3ZSuDMhaySlKHhg+ge4iP4EOYGiTp82J7a0AECyEHoLIblHQJut
mwVXwatveMtKc2+NBOI6OM80DAUuzFqVa5YTMREq2srIBZGvNPhkXhcjdCfTterxnOEOgZHNlZE1
3yyfYStIcJnIObjoSBdtV0Mfpb3N/Qd/BP9bJQS+8Q4TFr2e8tF5U0fdDBhs69CVJUp4U4gBjvY/
bnDAdsZWzJv88ENpPSBqABIujMbrz0cwAEsAmM5R2bIqSZIzSw5hZZjOGYZmM4e2CnKgOEwfasEM
wTWYH5gxuEQKVH9FPP+7gmYQY+5LGyptBJBsJUcRSyExvDhrpiomAjpGabiQBuqv8RJXxGCeBQ3Y
9jBa+EeuCcow8UseZ2is4iiCaaZcVj4c21EG8PnH/FP5ZtdEw1Gaq7z1hNnSVqahoH74kyuFbQXh
YwyN4eVnzhxbESuBS344jUSYSVmSz4pkOeTPsM69Qj1mFa63/cAAvSY+Ol7h3CzIZhSZ7//6Z8k4
Vday4BUGqCUqIItT7fKrDotOp8h8MrPJIpA2LldYEGVz7aluZ4TEdoPK9q9t7Pd65THm8P2B83Xq
xJ2YQWutERB2jjAStCQAwj33WAfwclJwDZQzW5aGdrgtMXZ0ZB3Batxu4kxwE2uNlDOTnx9QbzpX
MYVCl+iyNlNtleGF4/lNsLn909fYtD5BAZJJFK33Hn/riL8ovce4Y4RmqBTNJLUzObZaoqIySpE8
s22Rt+mqq3aglK0ae8KDVFibUEyJfmILaDFcnTdm2LaN+e0HPxy52nWHCT5v/qFZa14nDprCIVA8
JK7GNGgCRCgZvkZ9m2TP+YvvElEHsxfXxKkHKw+TCZidVRFVgEvRG68YEU251N6Wy3/LCjwFLOGs
9PuVGX5mwp8Rp4TVNp12RrwF+aw6r0OHTtm7KGf1p5COczc+FWvpIpRNU9xGm2YkIejxPTk6+FUr
Kw+RhuOuqghnf54+IMtrihGbBkRpzDYgMuVOtVSvvjNtAlidXgiu9Z/6Vs5lblVzR55UQDHn3KUh
K97JsoN/N2ZBBECvoISBoxFMI4S2aQAfru0k5GtEhlhLA69hTHYe202e7uuPuOVSoTXAUBWks7bZ
i9reOeSKRFDJKh0Dy0PfkCbYLN/4kYcEu94XZf/iTIGUOYbQyEwzoRl62bpEgFVug8clNuY6KVTu
RbP6aLAYIlUVYtdo7H/JTC6p+VJJP+dxrhJll4iiSbsmYBHR+TTPrZDof3Nj7Jblwyda8o+17oCz
R6eSNWoOP8XWXbGc3SCpx0uKPlkPg8PfNvf7rOgTkVGYlMSiM+ijqeO6prU75GqZ1q+dljuJ1uoU
U5hvqgp7i8TWIehgsZHnuxpo4yrylnPwv+LxBvXD9cmkLuKowdxl3pOE2hJWmfHEK7IwwwVHusZ2
LTF5f/f3tlhRxIaQfNdJpiCzGgRmMKnc9gPk5WPBCtjnB9R72mFzvxA+7gl+ghARBC4XLX0A3zWG
CSziXVqhEf755FJhz4TZTOA8ROigLrIEnbj2/h5nJ44S63h5YiWzbiSc5xCQb+5VoVbJ9g4jHP4g
xgGTB6y4723PGqu74nx3J7czAFvET+z6TuDkbGnBCXzKvf5NBje1X1nMJQYY1/5Wd1jS8chXyTKS
DYoGJfjRsQm5FFsNDBn42kFpALDbcnfK4SkzHmWGChx7VwInFtLqqi2EFxXZnDkWhT8FYkdZGBOl
sbEcAkSjAd2bUhoNXQNdZcgdjrhlAvPYRrdNpMXgMUPOWYYgZN6e+79oDL1Ac9g8DQobVv82OdUw
hYoC8rX0c9QvdwCec36VTbmWWd5OSTinMVf0CLq/q7N4G82yn9oI6m6018tXVpN0ihxaqxH3+2sV
T2aW7LqeM56tGTmbbhWg0IOSXYjDq/qJ6SUXVdkKDDZ0iQ+pRqltj15+Z3jmKQj6c6Gw0RWRhXq/
vHO6E0nJct4vFgVQIUgKHcZhHEC8CxfirEjUIKaNYKMc6vwzhur+fhEGN9e0nIvwrTiPRxl2ory5
uxk9LMdl9qyGlf1ScvjoMZNPYZiFxsqwlZnKY9qwxQAOF4Lc4L04P9tkrT+thLQwY3sm2N5rTyG1
ttpP8wjyuVWETpecwE5XWVQWzUWmEXQF9ctfrhQVsgvEMhCMKrwUuWFXuXEYdstXPDEdL6MD7Rl/
S7+pW8+wIsBFKHdggcITaaO3ITi1LXLpAlFzX0HqJ68n5HIlD93zUdNzEUyNmZ/phloRAoFgWzhy
QUsNhqvDXoKReNKLTEGCcaXxzb9z350m/4vnGdjSQWa+tqid3iGi+CdeaIz8JLmLqbS2JZsHlYA9
JD5+OwH/eohbCEQ/AWRCk6/sxistOiIoA39ENtJwEnHsaSZKKsoxTiMDC/Q6zMr1h8smS3bAcFaP
uOKEbteVNx938nU1aGtwZUlApydMMkAEm70k6elbBr46lTNszsTD0H51JZ8QVTly32pah9nRfwfg
xkY/4+R0xQpUqhbhgBsQH5txUaqyl2KesZ6HtbD7ZI3cVnJ6K+phnytwt1cypJTpTlctbwzDJstb
rAm2NNQ3BsUrO0KBCfigSPgdR53tx3mPxWXhjbuts5935KjLpJEPUZ7yJBLzuEJarxKBsciCM7K+
JHE0i9NXt907XEwJOlfAvKm+3zt+rP2aiycilVF446EEKihyyjv+Wnt9fXJTYcj8d7xaLCCmEOZ5
o0wkvUH2iVzdez9l7fxjIaBfy2iws3Pyf8amB/gRV7PbiUP2O3rxQEgMbrBT6OcZYc1ZmAArUY42
kuKJgV33khUtWAhKgsTGl0d1H0ILJLS8ReRFYfH0RI2V2DyQUtnCq+0kIG69cTsUYXaFplRbGd04
WnYw62nLeHjcYBYXF9To+1Oy91D/emdeVkvoB7hcWnr6YR1BO/maSDIlhZERCswWSf2dt+KxGmOT
qu1REBMOQSoJDW1klnh6zgl6uPvnzWZRthlM2tCaV7tLwkPozSY0crSajd/QyG4lpTC8h+PVauO2
DfjLNiLjTNliKkm1v/DRDLokgYUVBiXo4r+XNh1kaEjlwui2vdaUDoPqKz09VDrlSX6OhYU/Ir6P
uQK4dmCPDqYFyOvCxLp4mLlg+9sroQBMFQOuZKVxinR2iAAk0MA15OXQ/PYrBWQE/4zuFQe5Bc5H
m8bxjdIgbFRhiu+aInWiV2NhAKVuOiV/pPBGDCVa8TmtNes23mA5Fz7CzwEAfil8O9lbUHclMHLT
enFxyJxTVtIWdJbsAizlMTzoeGNXL3VbRuCKDaaozmcNmp/loRQ3qvRM0nMQ32H7t/yTsI7HNBy6
F/A0+nNOgh+1nKVj8lyLE74fAwbWFEqBkXRsta8O17ACzd4oyW/8NH7wOeZNCKuzkkAnYf6nFvNj
NpoGEv977nehSPL6waLpIrWrUNvf71dEZVY6O4Psx6gEwMbH0BKnWsyoI1W8oo2pFBNodIODpCMV
kBsZbeyWun0x0xHosDfrxe6FCJ71PyL6Z2Bnbk6h8bXcYQrseT+DYJo4gvWgmMvkUl3mBjxssr2I
/AMhxva7f2kFdmaURZT6synbUlKO8Exavayc0F4ax9nCH4hWM51BQ4CS8ShajFQz5lttntoxp8PO
g4Bg/xc9mO0KPbHnpM7ytvuwg2TqYJUtU3+N6nLWmNZkjjcZpCFk7/3Wf3DKe5Zw4ZppKhYW3gLx
jCK+PJFEXBdRZcj2vf3q8dnjsdzm00bDGrBjhjE1qm0rHJpQm1vc3uP/YTe/eiP70sIw90fBhdS2
CZpXobMsQe2CFPa5Ev0SOVMN/J7ILmXLiPqhHXMgLzLLv9UoPPx72cgvLGSbseydK6RjnP7l8FNl
wnQVR5vLcHgNx6dx0FMP3ihzim8t/rfpBIluaPFWI5i79Rr0JFyOLHNRGHkN5jgzEzApklol1B4m
XTfHrZY6IgFAy0wIZcjXQa6QuCAc8yWVo2OnxgwOaBzBVBwAxvmJxrmYFqOBA++PWnZ45fRPg/q3
G0bMDzoX8MK9QPYpDneVzWOElxEOwkX+Ma8mhxCXTeR1TTyqpAh9hi+s/9+bHk49fwJrOPAI+FdA
z9oEPneW6I6kQGkK4UUQXnI0GrubfJZGzAjOmFTC8wfLot28VrhPgDr9AiOWn/9N881ywktvGIKt
qY+MXYC1Lhvz78wOFGSSXUqY21v2Oi2mnVJ/hZsW8lN4qCUz/5lVvHu3vEF8hLsEtO5CJJ+LJ/sT
PIBvHAVdpTGIdp6DEPQLaS/loxlV0Dg+lduKLILZ4mPgfdoO9GB+pTyQP1aSx4k5+wmm86GKKaeN
hctbeUHZsuHR71HC4MJLQbCl4epC2VDBfY2ixofk+u1pHn27+05p6bA8qxzfTrsTumPBufD37E1z
ZES4aNsuZdgQe10Cfw2i22LJBwwGCbOG5QasSVCfx9cJY+VDgz04ccgIRxQSTqpzrykcUfZYymrL
G96hEqTWx6jdFbw/WJwrQFyZEAz7V5uyo3RsXKAMl+lNZF0vMnhT+4GkwcDZ9gUAQJYxuaCgFG7L
ucLYSgWD+lek9Rv2HUduUcwnP3x05JMhDdKaniv0ofpz76JtAMygU6tZ7sV5T5tJJUHoAkfwbM0d
JPNFCjipGdQ5tgs0y/6WACsQtSdWQe9LBy8LHlYHc1D2UKHd4W6SxYaPd/Z7iRdIvGWnhWcCK5QJ
pavxW5PgmBqK0WYRKTZ72Pjvj/mDURu9egWZPhDcIQfIvuyGG2cb6wvnZE8lE5V7Z1yqJ99cT1QH
NHQJXaJrJLcARq0VNe6KArVjcCH7yIwjYvv+wJjyG2IA1MSD1RrYmrjUESBKh//P74Ve+YAk2bs9
/m1YSPLOnSaKK4D8Z9MrCI1LoaxRf9u5WdCxG8vfn8kS/V0RRIrsayH5tlO0ujLiXZMsW2339tyJ
XIdD4bmrFDO/yIhOJnrcg3ncrC3oIJnOKTo/vZkXa0NrTQy6n9Nru8i+tKnuCrj4mYH6UDTkjzkg
satPeRdoYYdGnupw5ogm2jwrmIv94Ibssv7dAQ7tHC6RWbfj33rzhAnr8V7h23/eUFrBe+ep2/z0
/YU2fHiNe7fNVdiIQ2/TOG0YW/RH8G8tYzpaBiw3okSyx2pz9ADWxUL+6dZHUtP/nFenRpspzcKw
whjywZTizgMSDUx/YynGJCgAQmhCLJZbB76R3IjTiWkr6k3YlER3SKFnTaNrNXqIfhpheCGaYvsX
qRCQrgyM64yzFXdrqM0s8sFPivpM1JsPRR/dyT30QUlwQlgVZHJBdSJcPFIHWbbfYt/MJzpEASEF
BnRHVWN4sve6yeZEw4U5ypyjHCLRvTYD4MEdeMD+t2gGAeSTqiCPrcD04vo2VhtBuHHie0phW+qF
pdMLGKb/7kqD+7Nt8lAZUxJoTkqagEvN/l8vlfj/xKjST+OBsiK6zRXhhcm2WAtaXT1kvXpNLQqj
06cBh/szbHpxOY/X8zm667r4lzDFqO89USiylJ8USfakoJNR4WVJB+nDZY31pb1uRnDBBKd9dmxy
WRRJTL7d0h8D2oNpVCa7HhuGxqFt97gDMddBDmyxxDIydO49+4C8rOqYe6/LhnIS3NeyqtCysIut
f7YwfHRz8Vh5Ln031u7YKnDQe81iHGq4NhevBmjZidTMtJMFqwNNstOFsyw/KYD96s/MFfkFRt7U
djnZObn/NG7YhbU/1J41wOKakx/XJ/OqAw1SzxlyDZxdBIXd33lRFnd2ot8f1wCuGTzeZPslH9CF
c6rHqMtmqwqZ0j4zKXqkMKyy/csHeA5tdA/sKx3CfYHPQyyyopcZTZXKGt8fUADZJjNgOSecMgN1
9sgXmTwuVbnNedTIWo44uaEtga3LiJZPOzUxQ9LrdjrQlNDNNBv7yS6XtjlnvA388gnp+T/HGUWN
uwor1i8JeCwXZLRPTWvPi2EHfVAW+CwfC5fNe2Y1HC/SXZR9SSEeqnkxTpEs/uk+g+HrItK58iES
PrI+yMdxkJukUYvVZol7ai8qqh7v6FWa3F/ZhYtNv7XOWiPCiBgaYeXH30/GprzLZtXtjOz+Aksz
JqwPX+Oa5DDLkjHIrHQxBx4pJS4xRpcHfgQhkUYbhn6eRdIkv0wbNlXw00TAIQnz5syoGUAOKlIo
WLz2noFRZNKDTSs7+Br4JnXr6MLLdZ5H3q5S52z7F0t5A5nEz3/8sftUewrGNnUATe70bM4uAnf6
gkQZlpxxV1FzbW6GSlUDstoElRuLqq+bfGXUMnHGOssIfLrzTodmuGXWuAKlsKDXmkSagDFKxqkQ
WeUXORuNtA8EFGXkZBNDQbSl815/kSqjYY42NzXhl8014MHERjsYW9YIjU4Sgvt9RKmYw/KSggHb
+wdwa8OxdA/jchzMugo613SHdv1QuVv+ncsxscPL/X+pss6AyV8O29smSHTYKFIrudU73m3Cdd2o
Ek7kKZFeROjSIaTLKbq9q7k2WsxUc+2IEXq3WIs4fe+Xl2u+Ocwz3bzpPC0q47URaTFpdQFrXIgV
1cplFiAURg49Dsz0+tyScKcey8CLng/dtxss3A7AdQXQRilFyYhPpVkAGzQZvl2dbtQhJSJEgzdY
htPWrrWkCrOkPtG2rVrv96G16wLxuBMKBm82/bO4u/TcErowCq/Qf6ayFV0xtl98UFahQJCd1ixl
EUhUwBJ5EFADWsJPUgcKnbOLMdqiqssjSDOMHFQN4iUuQwmakJRxQpTDloafK4yz8OYDxwVQf03W
1JJgmZAXZtjCLF+NuRFGjJSL6g1vHmI+KG8onqqw2b8HUztmjPNpeHeuTOWwBWdaGQh016y3IKQG
8CWgLcWSV/R7JTblVj/HLBRiToWcHitHS7P6syc6FXguIHwtBID6F/yL3jaWe0h1IxWNjonIakGk
DWtOFQd2vIyIYBm6R9w3fcPTnkkcDj5oRdSqXPn5JQ1iidbnph5eYt1dBYQreABIl6H+gj078e/d
Yws+myUDaILxw/Ui29KlinFP6mZReiD6ELGw3tHYGzbmEOd3cdtR+CdlS3lE9Ltf4oOISNKR0WJS
m7eWgQJXHxfFccgRG1j9+sTauWbyb/AxTh07KzwJ/18byfqat0XP1kutyyrRSadn3jb8qJnYAa/6
7ZmM/7uAvLZc9RmpsNSRipGeDCnAmHj4lJdxD5xc4urUw5c/2IiZ/b2vKtXkHvNOfUHXzq8E7ccJ
0EXQabpBJhEAYLPNwhBmQzDawzUCK/dCIO6BKZpafbu9aWrIYlyt7u9ccbMspidtkrEDtIYhlVwz
K78aOC/Xnaj7VtHTCIvyeN/mJl5EhB5nhaGcCBk8u/XFSUlOycII8MIFLDuazhGJSUXG4+8t9gO0
ljy+Rt7kONgkTiOCk9m4XoGH5vJPUPEezz0quwNva+klqx5+qeEzDbE2DD5GZRJIzfpSBBlkFQYm
Ar18yo+n3kcPHvhEMaLIAveTlmmYNUWMsJnTEG9nNNszakuXAY/U6e8MHfl94g1FPLR4r9ArZmsT
5biw92Z0MYh7jNy2xU2EyqZjg7bUUv+LEwElELra9IXCyZzfh3MWE6V2MuJ1HR26kQFE925AQZFh
diQu6ACsQtipSJ3cCLIWvOK2AICivSgzBmkwqyGRp9xhuzOQawWCXgMcel248swWz7sdz+1yjdGQ
Hg73JMxWu3LZAeh35vyt7Z3vVd5Kq4rJbnOa/WB3awTq5RjkxgU7nQwAUzi5RHgyISp1Q0ux83in
R6Tb0NEmRuxqHsDTSreytrg8z2Dse1VNlZG+t5pnP0dkkhYqUoYt7aTmsC0uSZeY5tSfen0MExfH
vBXm1JRbwUYSskiGMY5eRpikc2Hh5ymZpbVmvDXcyCkLa6wJwQFCgSPzCHYDCgu+1CR4zJuM7RSG
DowxLdRMdrD60ASoLqMpxnQWh+bY/OISoWo8f3aFJz1QkrW2AXUvJoOKZXurH3/y9KHsyigAY8TV
6oscDk6sts0ZAz54Qfge1PD9Rvq/V4y68tRpdKdxGvhgZPxxdIkw91hQe47DxhnzqOrnZsig7dB7
B6hyFPB9bwAop8Ga2xm1pw1KIjVLm+YvSDYfQM2MT6YJ3tct+Iv47p5VhWdbyWDXLyHGKa28mOm4
LXR2L5A8n8uvQfj/byEutT3EwcKIuG9r/sCUrfN/NrhnTBjpjhQbzvOxSIoU1vBQM2Y0verci8FW
Mv/VL4KzxbT1oqmruRFwff6rR0fZKIYyXuRPg9g2741oVvOUVVJaYe/X7nrQbGh3/IBjzqoy/tRG
+aopv08gmJ0CVcJu/S/G3DcqWbl2p03gSGPdNfzFNC8wpd6mntX+I3jvbbm4wByut7db/WFCw3uz
bi9ApIS7zfGpdu5FbvucPrldwGj9lcyjmb0PkCDxQhNrpRFsrCR4zR+IvBVrDrSjDGerlDSpf/mn
CWHSJZ2aUMPskkvebp9d/Tte1Wh2olyLmpQ1q/7HRjXGTBn58QIP6++0lqGRbIxEkkficXIDp22S
mGYGOGl8EeASlJlqIXrjSZaa6Ume6zNVqGUhWGBHpxYGMkdUosHn9u1Y58cixKJSTP1FUI92xAKy
3osTPnSO3mI4lamIHG+HaSCKV3J3cQz0avLob4fdB+0KuUidvEOyjYo4+MKOx9c+muwpcB0EWY7V
ZSRhH/clUdi0b5ul0creaYDosGAOhIdM6IGeJj1xCCpqJY9NDJaTrgxyRPV1e4yocsy0kyezisBP
7HfmcJc7WQiJgovFAwUxXkbQnUFN3ASlMTmpel9dUAxTA51us+YzRCHcrqeZ9u01B5XW8TUr3GL5
YSsLwVvmCz1X1+Qb5WRHUKswrI/NSAUORcBHsgq8FhUo9NLzXO9Vue7rcY9m+wnjpBh94Ff5KnMp
m+zUMwQGAjHsmBMy01bvLcGSfSBsgFlOHTc/UOzbRhyhVHU8aQ5P4Vu9wItJ8M8rUtWlnG7aCJ3I
ntpHDBt7F5iPkFdPMfSIzpnIBq4GzT/skdz34fYAiUHLQAWTRVoWBfaq37/lKH/kEEp9eEmRQ66U
YwrTspH0yCV89uoAqR1o4M6nj+Mk9/l7pVmOPyVoWlL9sRrdgBGJKu+BP8qTuyC2it95mVjTo3ri
4FovUV6hOQysFb7vYR7ziOfsGVus9kOXTWrMXhUBfMEKsU8z+kU6Xv8K86YI6Xs3Ob1dtEQepVid
oOrRrwuOelNk4Y0XaMPOQUyj/+ekbnRww7GnAWWI/6EvxXZnVmSobjVqzGvaCN7UobSA65WKJXND
jaZ+S6zb3b/hgnrFraFXfbBNohoBYOhw+qHVJWqAEBroguNEVo1/vdyCAev6pufe1fbmFwpADAkM
H/moYiRPIpJRuIeoSRHTx409RsIsRnaKmcwHyb31q/OFZ6VtPrebh/AvkBMBiGC44AjQDuV9zdfa
8b/mumdHkgxV/Y5bi0E3QMfxQs2Gtf5WYRKiZxQaccu+YphRDwTbkQpJaPii0p6iDtcWQkLV2gbO
3CedCpREViKROO7CfKVkd1QebSsPuFFBgW2XEZo0zyiygM7C3Qt0ZBQeQHi+kUdb82frXYN1hj4R
P+aHZRcXk18yOvX/VJ1gjRbfVhDkif8ETF1b0tOoAk6IU5ml6BB2OlAe0cxwycKPcrgVw+AN2RHG
MVH0c9O9qxkiJi0FLdN4RljM76mZ+BNy9ZtrK6HOqIRF+4MN0W6PYdcqq/Mn+os9QXcYv5uRBqRI
fzwjyPZwLqxoinYeJZ1KRo5Nsyplnjl5MA1s1rLsEongwfuiYhcg5xdLBCPu2WNkUXRQtq/Rr4zG
cpYcoGSyi77Zfg5oWTkUug7MdrEVYXt6PL75avW9WDFkBUjgrvMtot/+YIg/lCF2yZZhxeeAFTMW
EPU744mlotQnsymAkgwBzxk4wOOnRwLXnsPOFRGryxU9aNvAoXsigdPLmUMolEfCArref4L4ysuQ
yMqcEagKb9E/DZFxKAXCZpbkVLlpLflDtxUvogIvSAqGlN24JfCXUvTC6QfW5l3wrH5dge7reyCe
MjZF2ezzk9d1QvwgqwYvIUsUQtDDuTL0IHk4t5NkQi6HK7DpmHUpyW8HDuVIvpPHXvvlGwjbYD/+
OdqjpHPiGaEoottlIjkZLGYjs9w83PkViCdSECkonldMiuMMxBr/tgsXiX3WapK11MHN808OHWrI
/IO3HNhE1DJ87se4P0Loqh20g4oy9+Wc8wB5Yqvgxl9TseAf7OykvlMuFZjnRp26ABLFQC1i+iyG
2czoqkfdqYp3XJZeuHZM1MNz5JqoU3JwvO46+gbCM9vNpG1SawtkkB/gZ4D/dG2nWFDvXNYDF+e6
TMaGZYVGFZOxfgRoy5uYdtLGcRAvtrNcT4ld9up7MVA3djkzYqkbiWY1HT6bgDO+WvrLmEF+4CEH
YyESlUtZG5uBLyi+VToST/y8btHkFTJ1gB+yROdAB2rpXkziMN9jPxWTURALgjTwf+e1jumz6ZXh
Nb7QDvTFdcfQrevIZuc2k+1sRcJ8oEs9HjUMu5Ia3ZYMPnqkeT7QrYt7vA3mSV9XvRBD0F80wuEb
DQpxM+KpZsk1Q/7d3G6se3ru1Ng8WlCFjgHuCIQ3mKn1Igaq+nGw16k8O5e1dL2k+qhPmhqE2Kfv
+lFS/rrHmxMSrF6RQCY7dKmh/6Lgo8rcwW468GI4V5k8eAJ+BGWJW/tfxuMPOJUYvVkay0nkKvPY
icixOYu11M328O0Werov7MlHbD/aZZZIBvVtgE0ai6N/H5TXydxnTp5O9VcmQDdOytw8spw2Q1An
TzyGSQ70Nr2gn6g469v/wmgdCBGuyTQbIlqo8LJJ7Nl2jGQm5Cwh74aKllmXx3dnQ5ckVjw8PrPi
u2a7nm4RqQlcMaQSqP0RfRDW0VhwdMks6tC2uzSLDuUPPjv+D/G5MlaSFuv1/W/9Gh3JOZO4yZAR
MvLtYyxQPWTHduwwEtJJcEMNr/iWb9yZtPCxKlTcvGsgunCfpEONjgVXqkNrsaJlWqLCCpDoahLE
nfj+PSHpCLYFqwr0j7uBrroqTgcne6M3KizH69iPGaDacxefrdaDcE0jejwjuhAFMPO+QilVVGGc
6+MW+Tch/cQ8WBcvdPTgX5ugtNAVpP2bue+HTDeggoY6sJqjxnpb5Pvy9mX/+f/imWcQVGAjs/gF
XxJ0uORfv9QHuqJqyOWJ+CleHxNABEIEe7emxcFYLx7aYEXNyiixxYyL+puDcsYS43ogONVdzuP8
/DiQXvyECadttiQHr8gb97/pgFo1Gn6swJKnrt9n68Vy447KC+wI4fWTp9U1klv346MRIFCMOv94
rSQYEg4qOOftzossVQNjICLR7kCmQngL5U3e2MXPNyQCjULAUJYu77UuOBbUJq0KHx4+NxprKOeK
bmkl6Q5kYNfVgYBk5m4WATv9sN9p1wVjf8zaiozmc+yGzrH8nIDVjfHIalqDnu77yKoOKWAtJefB
wdFap2IVLedEF4pF39LAffvL2i9ow9Il3ynCueA4d8u7ImeEBNA0hq7vkAUPYd3qkfDi6pUIn6yC
ZC87FR8MtEBWzlW7JaW0xHHd4Kl95y30HbLoJ/c/3BBy1WZw2gN4irRPvtTSZrtX9BP9orX3kpAl
79ir0N8Ch1r6AN3l++Pj/s7ZWpdUcGfWjZq38LKUi3m0AA0PylGuMJOr5e5CT6bXdM8TTvuInd5F
PA4vuPFs8FFrfPbW+koJqASB6M9gvEGqHmiIBi2VoVBPnQS09XTYEhu+C1ZdlF+DFTtBaQujt1uB
AApsTZUcukfpCFT+93y4BfrdS+/ai9gPFyc5l4r3sNzRkf0+w2PFs+/6ialyWxrtommLOfnJWpQw
QFmIb+iyh7tELYL4edtE2fTwGue4tqk7SYLsmYhaVMm0o3rr7tEysIiw6qxGAteR6X16EpIOT2VU
ay00UJz9NPPhFbtv1LD73Bnh9C3n5R5Y6xNx/WDhbkl3VOZNtxbQCFELNDW3VYgfDfvcBUB179sQ
iw0t+i+xZ/qiXqjjk4C4CM+Imh0pkW7ZcM71dQ7Bl2ggNR8c3ztG6mhIfUyRAoaAslkOrWCzfJoA
RCCfk4hWUQcpsXy8A0gqUD64mdRJO+/z7sC+5NJQEgEfRAp0BGNwrYjzFARyKMKJDjhA0BKwL6Hx
sCNTFYn1Bptli2XOMQoRPui9iYy6Y+4/IdOzxQhUuCxykSkRhBfNKCz2cZUJPpHs57peNFrA11uI
8NDRkFnWgmTn/j0pi/S6/CU1MxnjJzmQ2z2Lb7YBOr2rPndNznZkKxQIrzmI7qFLQVDxxWViXl+y
dr2kFykCM18wnYScTwbDomhLxaa6K+0DLHpKCsbtuvo+OlDLUGYx0uq1S45yUZrf/OaTwvDDa++X
l1xc1V8xlwCMyKqGi8qmXL+bEOKX02WMgQXPzx0ubLwJdrMmdG6q9HE/xNcQBm6+LK9i72eNvvC9
2iBG+L15irYV5PyUf54vrSN2e9pIOP9NF7QrCgIrPMVUTVUFvv2xpRozR2y4jRrCLXiWCVqKa9g0
EFTSSC7O5eJNhW93dwbxNPLcLsVS932lD9Fsx4MFUUPNjZIdP9Q0HxomRBksfhBuL46lI5YUcZ9D
MeFACh0EEj4wKjMrGAqoDVYoAOhlEo26bfv9AD42Zi7+8QyIdFL5cyvN1cQfMvCeWNkNshx/qbGc
o38DLXYCFWDMxYCZxZr0ZjJ/QvB3apUmKtOfZa5ghrjR6Ua5P8hg54t2h1gsZVPVl0HQvfBoOGfo
kHK/SNmUyH3cdXbgq9zJQeNWwg5VnZTjFPFnG4hpmPR6Q2cBdZVVxEaO4rdAXjJVYTzISA8MwOS7
OPg58kwdWmzdLKp4XciMYcfABvejrrBrX4msxG1SUYnTCxZlkA81L1nWB8vFKZRb9w293bXNy6xF
MgAnMtCRAWZ3ou2jj8O09GqvKZISN8P8v18E9nCAH15jdFbYpwKkA5BCoSVEMSG9oiCKzl4dGzNp
iW+OpyTa70EKfoINhLq9tgayirANXIVE4rX+PUXrYugFbKX4sxMhW2ePyLWN7EYCpG3TNLT4lQZZ
MQLf/BR7U+sFX7v9GTlo2s/mbQnSnkY6Y9Cw1QPKHu2rctrPDDgzz9CbRBRWH6x+Ldq9m98S8ke4
0v9ro/0Ay8F4k/M+86NOzjmQP1z9DyQjZPF/khXRVBkNU8G3le8wPYrEIntP+X6G1JgGMjh7Jjwa
JwzikVTzqKrcTEd9f0QodHm6Y7auTX2UYzQMzrqHNJG39k9Kmh4OC3Pmcw10nV2ix0ySYdRIo+Sb
LMBnT6v93kuhIuZDeex+p/1MWvM1/qF2yhwm2GK6ezLYpxx6oepvTy9qiZPuJVRQeF7wnv8mK3KP
ETsM4epWxy9zSi/G3rXidGewQYN4+F4FGwR4d+Er2/Xe/WHKeThLAPm4aPkd1cnzQNNbK3kSlihd
jnMVYp5vp82LSJz8ZygV8JRPmwS5tEgmruQuaqgtaVkWaMOh1o1sIGmozvyibI7WzFFpsrRTjeC9
ih2sg2Klc4jP+8oYsWv2VtM8PtJXANmva0hEjvUrm6Dedln2uqro0MVGah5ZTr4boYCjDYeTzo48
0SRlazff/pO6Lp3O1A7gl5HtV1a7QlEM5sF9bn1FhU8u1SeQJ8b9DLRYaxpCAOTwSjgj+bebqTU/
pV+639VONzGptIa8NI5iO640cHxjqIrOmKPoIxJKInwZA+i59B9MziliHwqD+sXmkC9om1vsg7jZ
Gewi1asSR4VPFxRa9gJA2joBQy0JC02KHdbc1BmR5YQB4ZGmv4p2e6uwdzG90AUGNxpt4kduIU+2
yA3BFHt0BPbdTR2L5iYxMkvg6mFL1USuSjee9wqFHEZj884HNmNT7i/4aihHogHKMQN7XTAikLJi
zJp1D5SYDYuQaEpgEgBXo0mkZjquDNtTirayl/gIEf5z70u9DtHxGKdU8QeCr1j+TgXQPXYuDrvI
qg4lRgfXuAGZVGFCckU1IF2q36LAV0sJ5wASQjmLRZxcu1WRoEytJMJwRcQqJI1szmTarAPIYRJh
3HYmeXjWStv7VcBFM+MkP9K411coA/cz0dzugirun0oQJF8m+B11Mz/DcIT1XwRMAb+hOHI361Oj
MgQ+PGaitHQMIAB6BbzQb0w61mYWwVHZMeuucp7TM8+4S5fuOcjr9eM/w+1+BiLxrz23BOy2bYbF
rxMSn/y3D12NlAZve2R7Ppf2pMVaWAjUc+G+M147aE6QxpSosFeJ4iiQNtU2G6Sk24lzGTH57DGX
dtlKi+IXw4oxST3nxM+q4HHEgzPeGHBuOCx9Gbn4pgQiWk5Rp/pdfltLpCbZ64fGC8rJVNAhSFvz
1BPt9H6BV5AV7F0/XOXIehzEDxUvo0HUF4UhFBFAccdqVG6hdIjSxovLKq70UvvDfa3gApge1pUc
Y88Ue2fT131XRN2k8xdgZZDNW8CmRjPbQ/NrvPnQReoVvrjKZR1ouWqq89vZc/MbTGnVn9WjbmvA
P3/sq3En/pdXQ/pgFEX1kF+/20q5HT25Ne+h2lJUpAe0AtlJP2UNMHtTFp+//RtwnicskGF32u8U
DxommNCx3OHCo9+CraY9MpaABaFmes16NBfftWm2dsq/g2GgVohsInig47XmnR02ceq1ge8sRTrZ
cAzjMHrkTexfV7rQFDgPH+PyaxxmoxSBr/rQPztSjL6CC9OnQCjMhXFmzAZO95XAzyVQGeKrnDWR
snb1UDtfxqUQjZifbCB4FGPs0v1YKc2gFi0nRXaW/dF/dCvxq32rJ4Z3bqpxjUvUWLW3MR8QLNWY
SKa7Y/e1VuTYKJpgqJqiNIq3u+Hx5rWuzNc2LgialgNesQSa0487OUX+2DFOwle8p9ij1yiuH4uP
aip4O4JfMbHGcjZtLakoehPH7PYsXoMEwcaTbqfbMNvrn1Ravowa2gvy/621bnajYKlDJEE1JDfx
324JaeobdyKiyzSzFZ7h1yeODcV9vB1CiJ5CNh4KESl/Vw+1/NfTvsPUW3gvNGlaXr81flxUs8Fl
c6tCgqDv6xAXJKOYgQydDDQlPmuTwKN0NPiEblC52+AiDrbkSUwbPg7QgMiL6NyiBOT24kuwYglm
qkJTPeEm4Y/Qqj1BwrhETkmTMtIuSf9BydnajyrNhksOeAn3+sV6pBvHp0EU4LrYfLVOn+syJOZz
6Bd618dX086Z+3cYBEaywAxa3YORX+uOCeJR96aFB60XP9AWe8JYx5iCWRHTqzJrNSurMHjUv0+8
T4IMozMBY84gWzREZ4yCQDDhIskTPXb/aVriaps/897b/WD/KZFjXNrG4duKx4sWezE7nIAvK49j
kT6XuKF1XpFC2AwES/PPA8kGswprMbNQNDvS2q2knM62KnUI7y1uSDJqizjjaQzEi71i2Iw8lFqX
stzHQdfL3u/5Ob57P4JwMlfcTX8eXxIlEjSV3M55IrE0yC2m7///gfU01hL5LyCv5NTH5JqH3zML
V7/JEc5TpOZVdRZ1nx+fegR/XB8hGj8CWi/iiQ1+g6tydXUtzk4cZhpeUPwOK8bfpm+sVuEt8LoC
amtT8ZheuSvAmTqWbUvr4iQnj13FFa8cerMwNSh/D1MiTmDiuwALBVvAu6m1q06Xt2B+PFJVnyQ5
uQI3yVa6yxZkNXtsmqv38IFH2XMr3O9n5vqBg1qU4IiSVbDTeICKqht1z+SDj4Qxiq5TTdE48YKw
9nQBLQ9lENBUg6y9lGaQH6Z0FAEO/0esBKcnFNBtNqnro6aKhqJeoWRkaMzIfu/IsvviQraF1pGO
zsgzT8ug3nbUxrCF+hr7B7OYOYlPNNQLAyPoq2GUFVjn+SJhv8It6nkpTcOvk20F+fchhR9mj91m
6LIZMiK5ENAAH35LBW/pXMHwjIckq1HhPehTWhdgi6m9jc4uG9+zyg8T1BE9ZVLYwFMU+KpGYzPx
NyZ3zYhs98UPj3kujrnUDHofX7dcuyPTH7emUcoavmnU7OD7p52PNfi0jMfRhG+NtFFrIpUQHK4c
aGmFANuq5/i5zxuOAca6DI23w/3G3A3OEkqKfVYufDYCt0U0hDYBwRgqJwJKC5Kh1HhQOXdnr47+
7cuRsfiiGsHJVGpAjzX/Fixy2VcR649SNir+mVR/Zc7EYWd74p00xPTVy0uY0x3JR9KEcQWkpoqu
j6aFO3sKCCu5u+us0SINvpl/VsymKIx3ZsRTYKPXcJHSzKzPJ9tv6wnGbsgMMufqeHvZz452dqgi
pQgM1KaIUBgMhHJbd8zjclAJIb8Vjo8WESaGAkp3gcqbSuxmHoyPuv03RF85+Y4JocJ8DHO5kFq3
6FIuRkc/wBR3CxWp40JMABUYeIYHufxxClb7kQgOWaZ9QD/49ikXWvc/91vGLlN4i1hyq486xoN+
iwvbSeMO0CtMGwAElhAPY61KiSB1odMc5KQEeBrVvSroj4npageGLzYXmsStSWkZWndC7IpRb0W2
sasM/iarRbyd2xoHZG5eESTgX2JK29YultvPqZ8j8IU9r07hBSTPgyNCFpDpkw9ffSbJnbze7k5t
rfgCJWascL016571SngG8SGZZYLCkDHaS3X6tIsQDZMHBRnq4OswjRr53nzWO0Z8Y6j90Ihk5jvS
NhrrQplSm+IhvcSKiZWu2ahH/YR9Dzz1SIZ+aRyeckux3lGrwObUXO++49FlpqZocSJDjXJqS/JL
eRabfWhBajbmDwXvUDFCS1ba5xTcJfiq+d3FQGomWoQ0Q+D16ywZb+MUVy+8/qfWlb/Pv53Y0xJb
aAJwh3sMs2y9jaLTmj2gEnt+0xKMZW+3D68lAdEx+YN6UBW5ZLaZ//RcJEK1vysqOrn+ctlZzQjs
asB+WFbz7B+NsxR+XebG6PMwlqOmNwaLtyKnC85/7sRp3m9rHGuhItSJ3yAraHxbAGXJ44aB61sl
idtLyMdiL1Xr2KLUzb6nJ+ZrHADlCK/V1VUk0hwnDYisKRY/Y3e6zA7wBK9sGlCDkY9uo/fIHoiJ
/cRtcR/YOSzeB6rEqCyrQllHvCBqeMTchp92hYXmuWnA58oECH/go47i5rc8uWKbnii53M4mp/aM
w8DQYU0ePObPXqDjvlUvxgosFDPioDFe0ZzNa78l0BnRuN7KhD3i0o+pKsDF4aHHqpshi9Razuaq
pHBHHAcNgMH3juRVVC9w+FWrttAtzzLbOCxTbZ4dO/8dwOEYod8fSItuMITg7uZayfr78mDMSfvz
NNv2jzhfpRA3cdOFAcm+59OCwueH0lHhlt2xudWNusshOZTwKSgRgRc7SGJFpKjTHmzU6nuw5lKS
VVsBiyfPo83NyIX7W/gAt1sFYESxHi0oyJh4lSBPsAYJziudy++j7eWq+fP5N0qIL32BONVBcn1a
jLcnSf8rjsVW8ccXR2H9TC/vTB9126rlOngpb9rZQVfk7I+epSwTnUFPG62egp49j/0XWIdjo5Mt
HWBKARLq0MiHQCN0I1xLrAcjGvZ1wevNLUfei2LOoAcToX8yRzX6CPvNejS8RnUu8odBprVYpPP4
3fykucef4EH7kkQnBv5ZOWNEBMBO7c0d/vzUl5nW6dlXgusERNXsaHTJ5/OpCS5zX4feeqJnewx5
0hmZ0rs6tGnr5EF212U3VnEfuBtTw0nSmgRq4IUCoMbKLWn69ATj+OnDHz9Qu1+ujeSw3tvEh1hz
9aggehD9ugsYgrNKLTjeJCBz0aZwCtw2ga2WSfisecDXV4MwE9DK1XmevBeouTABaZ/IfnuGAoKi
J0bkUdqrops5cnDti+W2C7JjFdJ5IKaq+XnjhybW2ek5RnsIBxozytlNJTHD4C7XjEHa27i9he/f
rs5rGTcf7lTOrzTXSTQgNA0g6oWzIvB+b07Vt0wY/bBbCOI0LDq1HVA3po41LmyTS75S6nKlyvD5
I1ySvecs65luoJFUfNSYY6WhOYl5U8c+U/SjLcQE9lnbD40EjnvvHYkTenLRH0s1bzvApdBtSP+E
Wgrv7zJEA5uE9GZI6Lt2+rOlm1YPTTOW/ULM3gl7Usf0cq9im60ie3E54Tr9H1sZFQrFan60zV+t
Dg7kW+vf8/O1fe/YvP4eiBFL5gGqyNGUnYOswMYwQ2ymbaGlJphs0ObggO0xieeopwJ0ucESUXRC
MbGkWqah5i4/R1jhfCjx9eoD9qUUDxKt6uop/6bPk+uwGNRRGN2zN4uD2pNMFagvwYw+RK1mpDoM
HQfEnjRbEIElY81esboJxohBRxkea5bzRV5D46ws2mRJv5zzw7FQ22GvpmwdD4yuw8qVKnDx1A8m
QWe+o7hVjpiPl+WS0tnJj5wU/JtAcZ7X4QG4vHV+jKblyatx03eWDm42pObGikPXjyZKGSr+YM51
IwdoPyHyIbN+T7Pi8iv3LnSG71pD42zj/nStTQK03TzYur3gUsXYKUZuTEWmAN2NX/bwMRpOQqPL
ULgsD4QKabVUTV/UNtyP/eR8qS+1YoMbqfgOXuWUukjKzPqrt5krEZHTv7q4NXZBJhNSMGcu0uiy
pzFC5TyTF5hBYoLIgSIykVLyaavcPIOIpcHC3czlHxlXk2QT7sC730fHj+5LFr+MaB9MIVUdMKy1
DQU2/iPqbTNdon7nr4siryx49GpFLb/XEJNwSegzzaNp7NN2VOsTsf/lE7IUzNlLbrvqapPcoROe
xmf5NZcv5dIemtuhldtEWNNwI3LaAaae6ciNO1b7IRp7aoZjSezbPZSqKPMM7NV1+DebCYnNxM/X
iajS3duxxZsEaXZJ1AGik/CagaalpT5ZveKvnuNaAbldmlL3kgWtoiuEUL22l/9JB3d+H9+A1KC1
83W5OABF4hscVsAb61dOfcXwcxgl90ZYuyr2qRg2Yx//i02Mf/uhc8TG0ODI5dkBNyEungeKxUyl
gIEvn5EcVEuy+9LereVmVW1sxVcIy/dj5obUXHDkmjoOHIuSgZUqSHaVa8vfmmsp+EO3roRQ0cwP
QrVD2uSTzt5OniFSQNjR76Dx1LN4aDbDvaygj2McgS8zKiup5mejxBQv5e1sXE/3M8nFObw6ydwO
0ua8zw0aNRBBrUqS4v4tOnColcjOlZIqF4gfnPbIqJjv8zPHGXxidlCEJYYSKvngIuxd+9bX06VD
qLoSj4K20/dm11a7HznMYCJELJYTDXBn2Ql3Jx+40f1P6fJMDyHDzuFWkLanP5Db62VKzk4uQfJ7
hVJmVd2kOnUeY1Dmo2trE+OHFijq2G4Wf+5aRHJ3QpLvqhiK4h3CSCKBvHB/GqHSWdOVDzNLbbyi
em3lLgI0sKK/LjAm38fxjIcAEguBE8i4TmKPGZ2Iuz8F9Fm5C0NL76f/5MFeK/TAfpixBlk43j+U
mwjwzoGzRV6uyi8IVFsgnLLNapNSn/mcaHj/KeICIKC0ynlBbd+/aeZu8SV8AKn3vLaDK3wnk0F9
hWjOKeAm41D02BtV/9dq/IyjmoNXlBHNYYimX9QFW+5sVvyP0Ml7RlpMiBcpXGJA6XZIjYQ8ufz4
TXvQOrVGqiuclSipsDVVS/ZByIHaqMjJI/TE6KkXnc/6Y0qgNf3/HevCIHPkuOEUZQ9rdhEcN+z2
mIaqB5bRDIRB2009Q63a37vsUmXD9MobEHX19ZbcfN8HOoxsoYMBDX+XQFGxfrMhEnGzF3qeMDik
BjiCmk4RX1A41ATqmRxjcQtwMKhvmVnbzXH30Htn0dU+59Sp1ClSrK9ZbWCE6+fOgtNvJ4dD4gCq
3ohjR+0LQb+j6oy9TIT/Z/IagadPbRbYozfpLgJjXOAvMg/qryN/ou1EEqwyAsPY0Ziugoqah4QY
rNJAZuO1KWgPbogmQl1sYjkhPVnpOsN034J0mLqk//pDqxEoGfetqS8ADFpzIP2CWH5NfrvK6o62
6uRlsUOA2gR3HVueT3yA1wvrA4VEz7bDuuQV1ix9BNfuh9LJs8wdWabotfZ5+Z652rLVzVIDGUP7
rB6Rdm2u26Bz8J2VsjHH7aXR/H/dArt/4+7Vtxw5QQb/GZuLqu1qfEiYXhSsjpNACv7yZQ9n822p
wNMoszpr1fN7sp6r+7s3IU+GfanEARBmU2aQKEZgwtazokJimXvkMhpyWA2uyihfTbslsyeVjtfr
PijjY7g4pdMmmSqZIfGg5Lhof8Ao/Ml/cAHwJHxt4/wZ6rfN5ETNWswjA/o2ASuXCmURnQQ2j2cn
yCfS64aZucyG9SS8nccIig08jllX7SOImAifJ2WmQ7fyfuldTkTjIirXpASdg4QQ8Yo7uEkkodsx
g4/1cqQEQ0VJlvFL2xPkEpjpMB+oVxPAJZBS2tQroiYEFgW9toQuOWd7bVid8Jz6wZey+CcsUDAy
JOYsXVn+Hjk0z9FACHOyMhvj8+RMV2KMeKUArT/qN2P6VNu7YurTXJMBvHDFNX8GI+VSTNYoLrgg
dIxMA6FBkp1LibwexIfMRnXY7F/e50KvLXDRlqOcwsFzcKT3UtLSs11rayiH2Wmd72OEQ8qeyFvh
U7seIB/gAKtfTn0jNIDFtn44YR5pxspFI1O2oohJbr2nzdQ5c4EIz5xwPWB7JXFgtM8xy3f/AGyW
mhPYxRJkQR9HDh/hoO0kZfYGZK4qIR65jZfAT0rM6yViFOPDK0+I0ix53NCUORQ4FK1+HW89o6zp
YmRe94RQ9vv+6cSGGV7oPSGGBETo2y897cZw7Qh5xBM2JaqtSiDmO7Eua3uinvmHtA7jWmFOtmhY
xCDFa0gin/QIv78ZmBC1JlmgB9GYssMk12cn0q91HQ+wPNhvHthpBOs4x6y3nhR1wfOrgcUCK3NJ
D641gbeslKF0fzzNdBMyOblQhhWh8gTNkTl6Qid8yR50ve5ywzuye8wS1j8N9AQYsbP06wxNawfF
lNYnqw1+AptSQYm4FDJgiEDcLccpWUrSy0vgN7kcjz8Icq+h2aWJ9D3Ow5ytratuOl1OOqorlM9K
2SKA22QTZgDdyKmXwW90qHqIlJK8uDSUE6BBIRw5yS9lBcivJ2Oecr94/UpTp1TqJUrH+KpKfhQe
i82kgwxdtnOalAjKG9PYrSURDUK9kNQv9QDCqIWocS4m5Wgf5+y5POujQ/SmS9D+UNekceYnpbWv
d+EIMMjUdWz6Sa6BrydI26caNobhwPGYQJLHtqMZUviNRP91iykpZDEGqT9ojbURFGZyF1nwdojI
S4mpwVONJIJZYCnr1CKb0XUbPn/mc1+AccvCj9h0duyVUPmEYLnCYBBigPWFxAKnxT51aOgTXaVA
+b1bt2eK2CSF1b6VNJ1lf2XmOHrOLRxF2HqXmx0suwYmCoRo3MksAWq7cDn2LLIykT/CSwn/WkfL
drE/w01UY61msvsxJTex4gOCN3TIFYUPVB9JWJe/4/bOf7zxjNS0uVkKdBYe1HDD5EyGZzoDBwRi
ZuqMZGXWKt8U9EKbxGeXBj9xSA0VMWGUkxaXzwLTp/Ti05bHsYPQfbBZ7cQya5sIGzSVSRu9Ztz8
yfuCZfH9D2EU+S4N+Xl2u3yjzRbGY+Zk/emJyYHKUm9SaLMVWrNknsUtXZFOPh1qbGwZL/wjFPcq
4Imoo7cjWt3DSzL2zdksO9V3CxhpT2DQjRnMh9U8TQVjvvFX3JDrqMR04RB/RklOan5qAbEO+eHr
PxanAk/dGXFpKQuAQ4ejXRT6UjIS+eC9OylvKh5HBuRFgDUipHOwL+YF4Z6VLUHGOPhW6A5zTGOW
gfR/RAIZzj0LzfVHORGZDtbPaz2EI3E3H3/Nrn0BWzxHmzZv8IKe0ey3qLvN4j2X1g5jG3iJIJJM
vqd0C3DSAAFrOHq0eO6K523qehbfJsF5X3erm2/ad7rkHICjn4Jf31fh7NBUwBHM/KCUmOl8AsI2
RDqSFyfA452udgo7W24irOGvFsxeN8FjV6yZKjomS+oDYY3xoHF6lK7bL2jh3Bj+Q3UzIoTN8AV3
7KAvbkMLA2qoiCn9vKERqcIUSHFDNPULz5QXLfC2a8cPipRGpxj9MKBg0Sl8QB8t2xeYMi+Hv1Wx
WcpX0eY/Igo3WBXmX56q7xvYhrIrI63xH1HYo+CodKihaCcKDoVeLKSJT0Cd4Kh72kItCnbaLh56
cRZISjBp+XJLILa8AjHaje+GE0Ikf9MwJn+MXeOdILWiS/Xu44ImOrgCXiO5P2hLqU0nrzJNcRgn
+EG/azIolbJ7nWmvnZlwTNILysF0SfhH97tQIltPWfZ0p0j2O+YYCiltQplnJS6dTIDvQKIoa1T4
nH/NYcgfNWnnSaSuUYnV4J7kRaCPACXTE4wyBN/gZrvQyeoOfW1BfG9CDUi/T6e1w9b/m5J6saQj
nkIeA46naE08n6N28s+sn+YP+jUBMzt1z+kpfrK+KcWbKU4Q8ZoL2rEKRXbx1XKjhqwGwFVm5Psp
IqmMc/TO2S0Cf5EAeca8cP9fzCHDMbmFhY+YIFjR7NQGfxfHpMh1ZR5NkgyGVg5X7rod+00m0voK
qle2M6qfe/aIFQ2woZesDGSDGHP2w39h7LE00fkk7OSoc6f0ARgJVOgP2ZX4mf4XHMFcqHrhojpz
Jrc4FiyPl/gujL8Qi+mGsLha39epnq8PraDUNKhV2KKU+NEWeFPAu1Fw5305G/GufU0SsHr0YbGl
xjHfMHSGPSrm/FI3RXyxRylVJEgUyyOf41xSDTnX3EJae6yVHd/VgPbTCRv3DeCbmymoVhsScx7R
nF6pI/hjp9OyS+p7Xn32uVvNOquMDAdnbsobgsApqEdflaOH/nmTNtlw2svZOum9e4xmVR3YVmX3
NfEVxK+ghB0PaO37sjp71vm5Z/QH7n6FA/3r+EVvP4nokfxYgoiyQAQd4NAx12MxijXhSgcaPZM7
IqggryfxKOEG0zgLQS5C+hlmuoQTsCTSmVqQ1IE4+QgLJwmNBt7b7+16gqyjgw/pD4XZpJ5JJu7X
9b9u1vTEL7KgFehCFN1fFOaDGIB+cgwLaNc+ENEXEOS9e5V0hWyhWcv+6qp4B3xtBRPO3xr92JvD
RN+yLwH67yi0iVbgrRQTSjPtgdJun/KJOc5oh8rXs7fAxRWrrG+dAfSW1i/C8YAEld257Kgz0YtR
GahEUPwpZXiYt0e545S9QIOHwoGCdS3XrmBYLvdGYdgWwe39NyEKOTTjhL3NiZZqdhrPBep2LpxF
TKINZ389f+gHi3t7+YA4qW/MiQnocoVWnINNAsK2ONuA20gpTm2AirKGuvHGhZkbp/NscHNxqR14
rADjK5dqQ9wu2uA2LmZjk9l4Ovd3EsRMvv3UHqOLjCvH/EVKsu//0CBRRf9QRmlbuYiHepw8jQmm
wuiKQXGsEYMFt/JHYS2sdr96MrP2f/1W8bZcoIMyL2dUdgt+v/VXc75xlGdD2njnQ+PD4PMglING
0gHSnp8obaSXiytECJbWOX2jdt22m10V/WGqqAQ+f8yfScO0MVyLVhhweEtkzHjZ6/EAJVgDMsYO
sVznYMY+oQ/TaH4GAxVgYpnUmDEt/WkachDmBgiM0f2h6XwULSkvd0x0KH6qw3w/oSuNvjSd5xuw
Q+qNEHRqg7gkF+u4FwtjKGjfVb3/FiNdDEz54FSo0+/+Vnos0aU/9iCbfAjDoMXcAiRds1X1uEwk
9Q5nbYue5zkUIl2D2BsTezmB7IrKDTl3yeYIW0+uLJagm+NfcBEEGZGTnfVtaFZehQXNNijyrORj
HIkmCbRA9ehKZSYewOluwGGUDsaUBI9TUBaUD2RK0pKQhv/OTdxgrj66EwuQAhhcrJcqFVbesnw4
vrOdRdDXw2D5+xVt2SG886DkMbLvYauhGyJgoGsaEiNsN8H+TAs4jPyT5oF0f+zyzBiBKvoHZ/iW
pbsc7Y71w87RkQh5mk3ynEWXlRUCLmQSGwPwiUbQoMPR5CJW2s0DmGthA9N4fWkOsuBB31ICUZpS
uhahbd56zVH9XbMaodIZ80+mc/Mcpu2a460yO/fQgR2tb888LiBno62XIebMO7+ORL4RIAXWjg+s
J9DW8uusl2SeD5MXME+sjR1k/eB6Bu72oVT7+Tt8wCHWePQkmKyuthd+BetfWCj7wOQKo8yVXWk0
PRbnTSC+dMPpAEgIHB5xDdpV4/1oNBh5Ya04/GQP6d6SblhMEaDH3aw9W04TXyb6z2KYC7TIvIWK
QBjSP6cCK0/ukFiNlwTQUoT+Z0uTIWvnYQmRw8kvhkGeS0hxwHiZaRPBzbYAWeNGyryeYsQExfMX
dTx0rmpItSfDxoB3u9Iz6Gpyk068RIuoNfZNBzW83TQi9YPI6wSnl64RUFmxLTZYOAdA0mvcn/PD
fdCwh1PkTDZBGhiO7s+OZc0vxsmc4m71H8w0IJUnKIJ7C+0vw/TXLPrLpyMxkZGArn6XaegSepvl
juhikuyS7Fl8WDBqgC88aw5Q63xqvh5ASCgt0+3/LIkQzEO0gewH7ScqeFXMzNAKqw1+eHbI6NvC
QBacsORsNoatpbPcbV6QYpSXzGxombZDgC4a5YN0fJUjdHVEHUXuqWJpAkZ48Xe2wbOktVheGSVe
VMhl1IK4SHfgRv9PCVAjE8aeUy2kQJdLeZis26S7ggrEouoUhxB/6SVW37YszxwMo65+sLsm6mLk
932ZGdC4RqyP4unDjpbjqvn8fDuxM74bOJZqgybVSeZEJjY/UA9MsowlYIfvzg1D6DVzUGp/8uJN
uvZ8gAmd2WPTagUURJRgn74VK8e1fRA/stfNi6kj/GdWNVppebtvR3fYE7+8m09hacgkO/h6u09y
REnSxNFwLKfvVtTeOhibfwxWqz+3R9lgQfd/A9WBSEciTYcJKEz4PpwficLSDDc5tBf19fmv5Efa
WrzAPnyBicYIGl9h+8v4uwwGteFWA5UyQvvlqLTEwj9HXTMfHNNLtwwIP43iW4cajr5SSVKsF5/P
MXyQHBOUOljuZnYWVj45bTgDParMO88ayC3FItkmbTJGPGvVruT/23J6vSyITsw8tNfnL73g/RwM
PNxZKJ03HV0/eG9towr3eE3mxOLoE8iIfXGhoCdDt50lxA9Ovrh3+gqa0ymTTTg5HXUjWzxL9owT
UZL3BOP89xAyd9rw+/J2yCYwa6yDoHx33cM9u2axgCH8JsFogRAij6xl7fQuBv+8Kxb4rgV3U87P
ES/u+XLxSG2maObK+A13q1Y/EUSWRXsGmRLKfpMFRWdt0y0vcuERNP6yrOgcOO+xYhauhm/SsF3I
pZMRxKA0ZFUA0g9HrQJiAyRcqoqy+xVzwgMmX7dnjQdNkIDhtiigGYFOHmkLt3cUh4IxHyByMs/W
nceH9jgjZgdpDhJWoVeQ7Q6T02y0wEx3VlNzaPXjpmhgnxloRQO5WtdJBX616H4qDlERKmsysyRA
TTfGA1dvU8Mxy5kH/BQgC+rcnuV0KjBkiRx+2iF5nlOO1wqA6lSwUdvvV+DNg2wgfSoQ8Yr+b7xw
eCO6axlRIUJI57FN9rCoMT/IYZ8g2ZH3Anw90ZAaM6uIMw3XWmzkpTooUsQn2WgEv/iydNuUDisR
awggk7UEzwNTJ6QBGiUi9hu065mB7oNhg9tubJ8I+Xj1hzCze6vQMjT4HeaEbhNMhB+aRMD4NRRg
SI4Yek76AY4HPpnX3ZVWC1G7v16X1RQ1JyyL4Hhf/1VlUozWnd/56upDfbibC1FdusA+XtAXHtlz
IaKj35eV5DgA0B6Dd4DDhZx6vrCnVuFmYvCj6IqTjC02bI3ZOLEzf+wQLGVmN5yOMgfA0BTnY7lP
VT3vyS2jxqP2s8FCFLUsnEaWohJ3mgDyLUvWTUBCYvIOhR4ld+tB+fL4boVEvXlLhn1FkF8HfrQU
EE5kl8KijwpYxSMVhiFkf3Ka7aKP20f8BHXdUW4tMU7+1TWg9pCheKXmxSd5VNWSECOpNCaa2TSV
/6CUChzKfa9kLMHi4HpS97pambA6VIUKEeEgUV+3wQ5dIcvytbcGmEMdTHsjPu8luUr/RNRQWgc7
SVbfp1Y8q3ZO8mSPAaBBr2yMoSNwFxDFh9P11dl8Vfdi006xb/G1Wkp6hWJlgA9Y+5qsbUZIvFlo
Cgd0npEJ4dQiot4C4gp6ZnvaaHikhTfY1dw0Ccq7ewJE0GEw8YzSOf+rhOtX8YdVNp9T9Beq6Kq6
tD3kh3VYiyoKkoFP2Eei3kCOkNNEIM7mkRYRsYES2pZqjyS6vDOTff/DT8vJkkr/yteP6LlVJcGW
BQmUYW0FXdKlkEqtRFOyu2ngPU5sktn9uYR/cfqJS6uCVJKHlBnzDWYTUi0vEVx9pGdp9w6iE5ym
PrBxaq12V1akmWkWnmRmSzUTiIMU8fnpaXpc7tZubhkp1JAoKTNL7kLs2ihh+ALsZxDfEMeV7RX3
itZg2fFwtL9en61gSlKLt5TkCnxs2Km+PmZQ6Oz2YbsbiT5XiOi+gscbaz63u4co+YeXbKg7LYig
rXLH+RRhQJPdO4OnpQG1PevjJB8QD6X7waaI56GioNTuZIIBvWyCLXTMlvuyoxtbzxZ3g24g2fim
Yc8HPA1Di/u1+AfoyVGgMg8IdFjkx3ILPu8RlR70Y85QedWur+xhnfBwFUXhuKc5l2jmBgMhEY2F
zuIYcCWVWzGalqZ1kVXf9zRZoMZwjdM25GMBHsVqul1yPwEnGKzZcKGSa9fEV2uQ6l2GLL0Ooz3T
rgmkv1jQLgPPPVAWUm+sYq8nAStRg0gIignU6oardC/dbnlu4m3v67zH6pKoWXYRJWQ41pKhaLLN
pKyjroYWuuFQ3g+ZrX22TzP65DWJuFoX5lVdn9TmucGFtWEhaj1r27+kbdHkeRvomvgQlKpozh8b
g9P3Gdyx4HQ4jWOvPtzh5NOlIjc6EU1tI6/2KHCEl+/PH71jCUqkxh//rzAaobkM9l762n7VSHBj
5uyR3ubs6/bB+wnGKaR0wIt5Z1Q5suwG4U/Cjt6oB/fAoi/sJOyrDzMpXhlOLT9FkorXaLyVK3BR
QbznZqspjaCtgfZlk2YfI9Qs4Iku7VbsvKBetfMFpSCyiaDt5SmnlVfZpgJNg9xOEMdxE/E3d7m1
WuBtrx1gCCyDa9NZwRHzE+sAzcvjVYq9CHreoUPlv9TNaG4pcibkT+UKMdMbmHC6P9E7lawFjIc6
lZ4DYlLYf1IDxwWCxX2QRO2QzCut6KqlBQxFMPunzGdoYKhf8TMjSvgvi57v7oU/u5bcKDQbDVD3
oNuIFf1VNdaml8Mze+49L66H19ohoy3GZnbOCQhVjpf3D8/v1Om/tOoHKE18rUcKV1fzscJ2utOV
8M/63i2V2+BZZ1H5DGZa0AqxFi5cJpFjCkV+7hy4ynUUnfVuuw2+ABqQ/iMm07bk1a6sjSK5HV+q
ocrBe11dzXPMxlZskynpTHFYFab4qegZWqqT+knYke/55cK8tcOZgX2e7yVydXWznfkbGibl1B5Z
fPl8UZAncSzlRSqmlvrL3Dp9l+yHYk5VN0pI5lD9ezaO/6Y7EENiLDHCcL63gAbJVC0E8BWHj0hu
XcC3xk8s4MQAZVmADqRJepnvFa2tLpIU9SjvsAQLa3wgso7i2GNEZ9eHJgIZxV3WPI1JdXopDgSN
DaHLp5kfWOxUe6HgkKQE9UHCvRI7Oz4OBCTv7eMSaukpGF+fsQ8o/1BDN52NKbZJgT2LO0DphzOu
92stB1tjVulDTkg+iwRG+r14EM0UcBQjj76bWXhpEbVkGwgVMpXFBPrFoR2WeWuKPHrlKkBPku0o
oJepCaqnRP1g06cfvhtdOVQgV1FTG1h2GE3OEMKi8t4KZi7n8K6BToIQd1b0YIehoDfBX/E8vC6p
6MYDL6Wexs1SdFbAm4EYHVu0xp1gae/53uV6E1RcLcFM//CcShaygJBV7WJ8w5kERnVSjgcoZ7nW
iskR2UPg5LrkVim6UH/yQ6Z+qzrS8TRvSTBiwNWOYTw+5kJmfhZ3tm9Eda7IFnI/Hx1cogaeo0x9
P1AQbY9QZSkwiyX7Le99usNVaGpq847tqCKV2v1M43r+RyLTmVUumQfQiAbC6QPrns90n9/n5Ugr
gxSKAxDWf0M/yQ493drniWnxns39b1nsouQU2O9FvuvJdQIpzTvzCNRvmehecyAf2emL9QkflyK6
Ilis6YbFsddeec/CmDV4+6Xa4J1c1sFX0rM5URzzEAAHjxsIqyOJfn0LJSut30BsSacqv55zaMfL
LM+6lkzWWpPj9HoGt40ys8QG9XfwAcm4JMfsM44t72JZL8aUGaEmGSAqTQEN7wF7XV6t4ctO2Bcg
FPRBxslpOpnYNusgikbNpyrdXr/hKgFsn+6Uh8nKLA7D8g/Iw/UHLnccTHkVnzKd7j6C/12IPKln
311kYXPm6E/PzylPYeT/hYgH0hBYuFQJgwpiBuJtSEc5qJ5MnETJSy1hVy5rOmNizgMx6XedEiWk
rFa99hi+SbWYaKkP5Fe7UZrFFO2vi/iXa396uil7nU57qu/5L1lAzxfmZwDqS+VRXD2Lgtq6RYz0
qchPk9/dp8nb5b4bfp37ow6d1wLVK0Iaog5WZrITf3J995+yR5fTXQqNXpt7qFJ5uUus1HOTyr+H
UAro4yduufR9gZnUMmzbC0Qo/q5lSbAR1u/0fRvtJnAbrXmrGHTy3yU7zAFdgS2hy0UjER4mhcH+
G/gJV+vFtED90BB+ZeSdDoxuTOs/lNXrbUSvaRTQttTDRsOxrwOQtzzQavcGkMJ4RaIIILmS4SVF
P1tPWwwHsfMpH2mBMy2b4KENKNcuN2aDXhEQqnajIbQQ75XQyUfdHioXSvNWf4Dqm6OQImvWdnDx
S7nv++qZNp3uifsrOLLWVL8BP0gmdw6zB44cfeHrx9ANUaGRAMTis6dK5U3ml6jbtAUAztwUmBLp
nC+Dz+F5GMj33qAy/z24OLuXk/c5XnsTqASnD/F353KMqQENbjaPUTfDSOI2IqA4IEh3OfKOWS2r
vi3pUeMNyCtLmMwQN6ysyftQwAIjx0H/sW7va25J3lbd2Ga6104w9lmzuf4MrC+/WYlin20mNw3I
4X6clZSd383M/GvCC9jdGAmMiZK3KnqfAlnsjd+YD0SihZt0zKQIbT34ckBE3WDPTyVje55j6GLm
uhExWvZj7br2z5SqUn2yw+5eEcuRIZ6AwNyo/W7+JqhJfzfbqzvWBJeAevLnrhvwIR0jSkhAHhlm
X6hTazwcPdOrAO6Ukt8dJz9X4BdYQ91CozW4fzofcyHaKyQMdwqUBBUkHf9RPAKAHGf4NQe0s4uC
eK96CQZery7qMPXAkrRVDN2Av1eGxLEHf7OBRvcuBqEhu1tuyc0CaPw7pd3ib9JB5S9D2F3Yl7Fe
k//cBpvhqgHre9CKiyS01rEoASzHmlaNekZvYo+1jFcarRQB0I9xPCY4pzD+Ex3dqj5dHSk24qNl
WmtpBgr3vkFCCwVlZ4KCusE0I/Cf5/XUecnT0/zhX3B9fFErsRivptkVMpWH/n53gwGBUl7L3FsL
/xFz/B/OUE2n3D0oIMFQEwWTzv+tJ/fh5YKzljguNMtmxucyxeGEe6XD1d27Z6g+rGNJpiqfmpYJ
90+t5Y4duBaT0uV1GPpaFfHbNEqWrOY+19zU76/HK+dUGJo99jxggBS/wIw+HqB8IK/AJWzduede
bVakKlXLj5GtDMque7GUlV0kepfme/T7yzzcnLSny3I8ieD1ITyS0Zn/MzQApaGHP9uKjrd0dSVg
mWPjrKc8XJ6/EZimb6+cFYsX3IkTOzRtEVTZX134u2oglRC8w9gdYheou6/hF7EW4rwIpxGJjoXB
9GyNxg+3sWT2UJE3K2oKHuXgKPKK5Cw/HHSuf/1UWFW4hm/OYzVmmvTrPeUevLvYtuXtFNrCpuSb
Ss36AU3pzAoL8VPNdAdelelafZfjjxgwjRGqQi+m1OPz5ILs6804PP3LrwzgEXmCvVgc6Io1pGvl
jthcDSOZlKu/6KVTbDTJNenrUhsFvwJrY8+9ZT6NPTQrnfSaodRpVHjCjb/keSJTaWw/tbxM9YeZ
2pveLhKzCH41ISwIxQi1iTRJ3EB0SkM48B00dxmAj/UxtltYx7icEg+4icugjt6mBJ7RDivNB3p8
+Xq16W4pJNeQ61qYQiREyR+2lXY4qSruqmLviT2SYfxBAY/cRI3zfbuCHhIOCTboGMUhW1eIVFNG
TC1cXb/MDrjBjNNN5A806tBKNfQy5jCdhlIqtx1J5/PzUSG6Jvi8ZJobrVQXw4zqeZ4jveDrgvuW
uWd8FAiU3f23ho9RtxVJRWyjYMszC+QMYxXvxZ+3Fk7MfgAlO7HXHlzrP9bqCp9IAsh7c8PCer/P
/hzU3ahHJhgGbLcJ5JXqVlQFKGviFN5IgAzaKhQ1Z1knNYUvJ1P5kW4TGkQW8BZIKFhnLejM09pP
b6sMnHA5zAFST7ax/5m5Z1g0s0BxuDMk6NbK7RueNYkNgGRiXTyokzHA802gvhPgMmgvuvv3mCfr
Mf8KQNHIg2ZtgJelrUktogFt/IagS1Dock3s3BZnFp7tfoRXR1NGKP1j/08SH/s4ztiSG0YtTkxa
x/WNvEWEa0oEHxaSil/vo60HP3WzkWKvKT0EZP7Tbd+bezH/QFFF/79xw/+wRX/oKgUq5OwqpEzT
dURpnnIMoxRjH+g/CEjk30xlRyvNLUkx1npy6QSVEUggzebfBRMYinG0xIObZwzgDlUw8itNhXMA
6rpEupAe+adWFtXaa1BnVn/HqU3euN6id7dqo+jVPQZhhlKREESKdARrw+XhHxnDGP9dCqlvaf5Z
ycHsEtkxIJhJ4vjfCYUdPwDlC6dEG/6dsZhhS6sOXI8Vxs2sIL+S6Y59qB1MHtL0jcTzASyomVQh
2/Y7bWOjyvF34rHkRk1EeDtZIIjv14trYs/CVCsX6wdz//CdI1TNinSI462n1uxi6uR1YkFwuv2h
B7OzlIZ4TKu/0HvdPtv77qIecFl692+tqOoqkf1UxemE1sDQTYw2g3WqGtNQwW56ah4GSUDOKZ3t
g6SDsAkDQjMWmGUcv8LawKcPk7b1anZ4+gqexUeHSxc7aFy3ChOcv5AnTRkq27lQOETvQms1pvep
4qog4h6zYo/4SUkGnAzFE5w/9r1lvbjc1BTeiJmJD0AT+4XWMsh6cC6nUsLt8Leawpj/GdybpxFc
dRQRAX1G9LOAehGDaFrYrquCYMCx5ReH0wac2Jd5oMiH/aItq1+GGTIs1TN9bgkmfS47NwYEDcQl
um15/jZxQf5NOV9b77uRCbqOIHCLy5YznZYESIl3C0+OoZtf2NaFju1mCwF+lpxFIJv3Fvmp4lEp
N761hsj52rvrkLog5ztIwZQa9W8O8MmhEhMW6VEO8o4GjxRmqEjPt+ipnmX+S8QV8lTLOFpVikoO
8rQbtbkJ3mYmmIjbjzqPvOeG/Ee1W/woPpwuUJOBPfq3/+d3XqnnPYqvgKp2Z14Z4Gdg3Vngkz/0
hCzXDIbc1qdrxP5Qzd+EOU3GSkgoKSzS07axUJDbCxyjcyWr6DYhv2DdHTEqD7vfqDq47z0g1GM2
TIvs6L90cSIMqG7WeCOyHE3CVVjgUCcZuD9NrjETGL1GWZHEuawXF937kK6b/QTNIiIRhBl1l38i
fr4udDa/PX6Vbk8fCxZpWK5P7ZvyFk1btTb7TXo5+gJznykxGWaJ7s6EWwWplnZIU0H8I4OpP6Fa
7x9kDwa5qjJjHBx0YiiZ2INIBBUn1u9Fo8TwbXxilFDKYLvZytdBWcYFjiJv+/BUA4sFShXOMr82
mK1hwkfd6ho8rZnr8ve8PbNyyVbj1Azv/pWlEpd0yD0u0tyEY5qG09dFo5f/Sm35zMzQT9MP3DFO
Vu1xBp23D78DwOCbNIteVsJFuFS0oXe+8yHwhxSkJq1IsDqMgOppmHQH4Hwn5xnLjvpJaWcqMN/5
hGN9CTaIPb5+wEKVc3N1xy+WppF9OyhDEGJ86e9cGADFwgGi88l47yIwEK2gs33horXp89+kzloO
M/q5DZ6j5vqPV7N0EcDwoqp8tux1ZurbwJjodsbj1p/slsw0/Poj0M/e6feSBi8s2FH9St4ZqS8p
gnPqhYk5ydTdqD1yZHLygYiK40oYrEfNg+r8/o3WqXEY4zEU1k9KUgadGX8O2eCnByjr6VTNw932
2N0TwnOIJcvnKSLqPahT9xDEdXjYXvviX7U2N9uDUh097Y8CZRLjyKB9XfUQLZq+RmeJx3R7USr2
CnckVKgwsR3NGH8qs/2s+RGJOzC581zJ3Eza4LQVVAdwUr9FeKqyudmrSq2koZDA16TDJEt0JCNn
hA0UC7r85on5KDGVRQdQvBH/3VLl2n8819ClE5stogznd+z5UJzTnhRFuvYtjkyHsVCYHzlWSvGd
DfDAsJVf/6LHZ9+o8BKAl4d/VdpnQvCPKujIBkd3InvmoK+vwnUEj7NVbFZkWJ2YLgtuSx9Cnk9H
v+GQaWuOLJI6KX1266QkWXXFHia7pCoztEork8i4MHW+rhjv1zf+/Fc8cKSS6ef/Gs3pYpVd9h07
5W8tPuSEAh6cY/NwHY/LF/oGhm7XFdLs849kCMa81cObNpVajMm75r9EQaFmMQWZ4J1I7SSO8EDm
4ldL8QV/ktXPRpPj1yKYHmp0uGHx7XjzTC/N4KKhW8E5ggTktqXyLh5XmM2wi/V+kZTYOYFKZLUB
cSkQB8+Cvs23vhUt3ErKLHoHvINRyCimbn5VubpZQ3nL5HGCz1dRBlgrH/Mu2yZne7z2yBwty3HM
qAivMKHf2QsW+HB0jn7uZOKTibZ6UN+iYSXMefRsWiG4TrdmJ2SpriqX559FzdIv4hyIr4YV2H1u
BY18YjCKkD11b+SwQ2ykoRwH1jtC92fx8eATeJHibaGNPMXJEyUmcje7dlMedhQyfVyjhVuyiYvO
ULsyvGQtO4+jfDFJ79Sf5uj/zaUdsBXW6wdpd6j9KCNjdWsiOEo7L40v6Jd2/zCPZ6QSpOyv5Oft
zPU3EfiHeQMur8ALeYX0EECyVgUW1Juq4G3qrM1VKjDdO9vsxvIzdj/V1B2j4+jbArP0VBZFK3na
N6uk3kEQdlV6ye1Pd8QlvTrrt1eiQRGUMxGH8xus/s2lPIZwiFtbDc/gFQU2rmxbj0hqAq/4pzj6
kVbY9R7CJqJS9t08+yXtVtfYF7kWrda0eGEupNZ6ZoEVOJFpEXKOCRdcosq/om5nEJxJJjfjchEp
5+yBeT+0P/Fmh0CNc41bRUAdke/I7Cc4tvP3MFax8K/pVH4xb+bvekfrvHoRfLhx4f254bGkf8+v
SEOcPHpD7sihLV5B5hxmQVJc97Nde6eK50D7tzPhAv9SyoUbPz6Lydxb2FJlOZMckIZp5tiU4tpT
WV3zbKkFRZMuyF78yc7k8xqCEyzWYc6zB+r9jBFadJ3QKGdXIbccXvoczG/wk//pMHm83JZFFbY7
0eH4H1xwpM1zYmGxKl0HMWi0zU7XF/Ji7tc0r+77LlZu47BF1MtmL4W2Er77Dno0ItElIEjXWXY1
xbtThSgSciFZ4clm34eHYOlGKOSJMkfS9w3vKBlukOXmBLVR5kh/6cAQZ498krGZaH5OiZ5SGmBr
1Lx8vGA7gJRtWKkXUc8MN/dNHbe4p/bdtJQYKfNtGjxVFKZxm54bsdWRfFqbur2DuaIlVKiNa4uj
9kKnUepnsJvrzDjcJtMvbVsijI89m56GSGLR752BoKP7S3pYOv54o2smfbs9AaZcHGY2KyYCxOJW
nt/l3297msWJzEVjp7MXGdo70eO/Be3LNW8RarM5PhGkx2tnZjSC+/qODMvD+cpzw2bBi2eHxHxn
PQ91F6K4iWz+kj3kWM/7ONamhWZXJnha32XaP2SVz4TyCCxJsnt1R44EDzAW3RrcbXeAreINPSgO
ybsx9Un6oGkLLE4Je8YO9lMmwOByTqSH4XxNsyvRokO4PRvSWX5eBUbPNToj2nN8SvZR350eYYMi
Ssa4iunWdlh5mtNSe1tuPKXq5yQ1/bI1X6/wogYch+OE8VfEM9zu8D2wFD/DlMcnk2qIhexCR650
Q+EfarkhPtTROEwcMXKBZr7yYQ3N+Ck0g7WP6MaoWS0F5R6xIMEVKNV2AP+FFmKMzgAnFk4vXINj
7+GvjAwFC0VxZXeYQo1mHdJgaULKC8kjjT2N4VMFh0xGYQDqJAcLB/LvWdY4VIayr97ujfwxsZ4J
F4anYnXOlg8bgTYzJ8/rCO19a22TLbn7+GUQ16aAn0RgLfLJJoVXamOCqGE8nYqgJOxoDCvaNPqG
xno3KWaJNWmbDS+UUJle/XI4OhcsAIo6pgEx0xTD5F8zBxMc5hoRnkCxg2xFbINz+pMKm/8Ve3qh
CAf4H68XT1py0hudhbAXfykfX4oIkN4SuYBrOSBcVhlh++3ie4KpTKeYAfAIu2Jutf7y1xylZRPV
KGf8VOOWI+mo5jCf3YXRuX3CH2KtgV/ajaKrQ8ckzyhHUEJPDUYoQ8zgmSyXUx0gJohS+3S/d85g
brlSbCvXgX6IF6eNsb9GYXpc9OPdZhe4vgjGabPQonFzm0q1WGMrndmyYsqtNDffud+/1aJJ3vvd
P+ByTs2iPojRSt+PgaqQViIUytVELI6Intzz6k6MsDdhR5xdRrT5jhRF+PKagpclRM+pp7tR0DiQ
vX/uMpg9QrMo2N+aBgwAtwHNUPzFJ97Aj59dk5roW7ymyamn5ope8JhZ/L7nHU0vzmaZYANxfHc0
Xt0qfo0f1Auh1Ifp184245Tx+HAPqKs8Pan0sfrrMrpUJS9qDKE+t5vE8GdlAmCtStssv/3Az4jB
Tt0RT51+0juUUrfgvK7XOX05fWFurAbwNYfkw5T855z3oA6MaqdQYEmSqnntOQMWfikGFk3fVUny
NRjN22zoT7S1PCqK6H8pZH55kN1Dk6l7uLw6pphsFZEOhuRJeear1p/a3CwXYxc1aurL3KuakxxH
JJJ/9efvXjfsa5DCMFVSF8bVQ3fG87FE3Ub/zK5dcTVuMBW8OmHdsYqEoIUOmi73q7R/Qzw3+pUf
Yn4JJ1xhXEj7H2GZu+u4POxS5GQBJHWrRp6eXRHJFWqvWHa99J6Xtxrs7aqP3a6tsQOCdKwrJm9q
12eYYuQH1wQNjpJibGBK4h/SKXRB4unJ6b2qOVt715liiiXNbaE3SLxTf4FYqBrC9QeHyeQ3LwjS
PGYpucMR57pVzTRGQ34EQS4J72c9XIYMHpxl6KiTcElR8En2ZAyo19ggS0oGTzdlQ6zUbVCq6aS/
IjDzUVi0R8NtpCE4zYX01+0ZHrELzFNF/O0y+OqeRDQOX5vx9qVp5jMI2tB6v7HBZkWIS+kEFBNe
SNYa1EOvhD1XIfghSf14DEPfIMIE+615TRtrQLFcdYtydimRiUDL16zzR49lvcSSPTnG7lUWllc6
+dSZMayQhqeTm8W7xme2q1ihHlCTD4ovdG3wpsw006HD2jmLY1frVl0FFdtHGC1aymorQgpGxHa8
zy4AAzkVUjS1Byot92uFf6Dw6V0ykKM7Mi6UPVCYXPJlVtNQIQ0I4UgH+3uA9LlyFfFsHzSNk+F1
c+aDREVypB/svG1IqrtmOmGxB1j1cmmM8zQxHiAzl4xql5vwBkdlKItSCeLveET9vctQdIEXWejV
QiuYCHINi9LbNkun7CC3SyylW+bupbnt51Bqq/ZcgBaGQHIP0/PaoHU/BYKn9GbZMVCGT1JPfGIQ
7ZEFI6CaeW3gg24LuWhSoIzQGBYrz4Cu65+O5wPXyJnv9vvMAUtn4E9oCzwRiFNYdCdfLiR9CiPa
qRHi2Q5OuA3mB19sB3izEa8qxrs8uE5UOtHpbojWyAHRZafiF4sFwUdcrzkVuzV8pwj44Zjd/OEf
NOlH7f7UgDfFHoiiQ3pJN/uzmEBuwlqJdRA/pofvsfvSSFgZEB4N1TrEEiMhwJqnnfZ9n7q1Y3vK
M4vmlEsFRYW4kB98Kd8uRKuWgfhnlZ7ogOh4Op8ySqJdgeTn5ir4Vyevo0t9tLLZ+q8n3FG8lza6
oEyEFfk38+YbqHAbciGBldA5SQSfk/3JKp8m/AeyXjAePS2RKFALtBqqG2IfirER8+oIFbAw3yFI
1wOfHhaHAdDkid1bspCK75S1aj98JmdUgAXQIhu5yoKcCUNz3QO8DfH8eEgw4g16dWu0hTSqOb0e
x6ci4ixoxSP5hf48sSG6ZvuYnqL7GNXWfZ47h8NnOT3OLZBvLu2unDDFrcAZCZbmWTAONcKi13Nt
WmRrVL2x/Vjsql3lYWm8xf2vWtqOqEMArXle0JPd+holN5V42dxMdkkwnpA7omYggPJSN2HGFUW3
gTVh2Aalv3W2yEVQyw7NI+3xCP9fUR+BxTxJ7zNYuySEjDkJqvsmK4MtPqXmkgAJRdV31HKeAiFC
Ma4xRVKMCRrZMTeBNpHH/oQlhsBqsE74l7/f09yo7Ko3MQrluVpdSvWh9uAN8T1hvnfG6llz4NhV
UtIpOhqpg93GJcr+IwZwLrGO31SHL1PMxX+MYVXSgbPeaxPoNuRE7FwW17cD1eZiwfDZr4X6T+fS
OdP3+ax12aKIBfXe76Zdt514UKeI7gXMCHLdt0GTQfnocYzHjvRrtk76+QSVIa7AY9WWQU7g4PV7
tXsbJPBqCzHv3dgY71LRuzZ09tNbXAgGrBLBJ6Xz0sD6RVLTnjRzRAQ5/UjGsGNdR0tIQleIiti0
VE02ExFDLY2Ki7tLA1QJAEO/hDupMdBzrm9NRL+KnfsivqYQQOckWmw3HTRQyrQDWc0zWKvHa0YL
UbqS1wm7gH+KW2b26x5uAnedO0gB0pklESldklov8lsmPttt59kNko0+vocU5dF1+GeBwSbrD9ly
vwxL/pgIp7NKEVVJMemumVZGYtiHEgi79NvLPe7eIzPh6rjliTAbeUCYnmqFCNOwLu765DXIhg1r
Uv+K/bqCe3AzQRNoO5k3kclgELQALOImqo6qvMYOqC+T4h2yFwa7owXPaPSoj3nf/8YqkEuhccIm
sBWn52F4uq3gp+4qOfKFY3hxckh55NVRi1F+mCWQ43W1BqP6eWWv1gJvlKmPoOW3+4ip1e1bP64X
xUEjiIet/Yd/HhqCte3lhpSxlRxPWmYPCe1D+4pjv6+sT8Yz978xZTw4JxMlWmIL3CkeP5swnchl
fS36FtAp2XTGsvqFAtpYXSc0sdMPsxEaRQdMNTPaDhJejOBJlVKmli6fAdhGxruoqJkupBiu6mde
kmoemhbnyWSPotzfZRucGRQPH9uHbI3MgYN3bwfFXVc9UlFtpfSQC5HfQxNBtxtCJrS2RZ9yuS59
qa8MpeLRR2k7x9t5UUM2d4jokSI9zXZLXUlG5iHsF6SyMOt2Lf6TWJ/Y72lOeZX2YojNu8h5Ghgc
GQk6zi3x2oau06iFcf9mnTJ8Kdza4kDVu89YPLcN7druXzDrEdEYPWqFLWt/DA3fwt5sp24bUlcJ
X3l8He0PSjT0zEGJixKew3GrMQwLDD1tt0r9Kn3e6Cmk06hdIXtptxtQ7+/3thtZrQ7Ej2Fb8NUy
NrSeDxJ2hHyD8ednhsKSvCgDxUoQpEmY27u5rfJNA4ZUtj67jrVpAoDMlv8Gu+QngVm3/K6jZsrQ
fZcZqomoP0tTTr1+9F56yeH76A7JuSMU+u0998AgrE1T5D/eAwhq49rslTWsXPRTJLSxAnaxKO2g
IlOEj+NSiueHGJOOn6xvbAu3ZrI/l8eRmJ2O+Y1eljNvMh2im6mVnqVxV0bsebOyRUwF4rUac9BZ
zFZAKwK5hWKzHHcXZZUzAUj7qOr/eeCDlfCeSuzs/hMHBbwTaQdGGf927V1NMMTHPnECxRGtIQnE
97o9HTFng2Q77F//2acgNGeLnmrqE2QsdWVBcTks5YeDXHT0041yFJyre1iEKVDwzxXprVPtY1C0
2ciGcwVLCEuMmSQcqYC0wwTSSFYaZHN1hR9SZsJZXahSbVkP6IQRhK64AAJ0SgtQair5cEL9JEUQ
Jj5lN/N+jAMWF7HfnCkRusTCLekUMeU3P8w1JWaNTLAfBoO6UmATqkOiJg6TuM1kUEpm+MiOltM5
IJG8M0c2Jbk+mp71PP88BHoKuRRy1MtEa3vDrHgbC2N8P/9uBtWp1Gd3MPrb45/W6mY72a9CT7rr
LbEBSb6vt8qTSufh9Zmk8RYPL0Hbo9hloE4WWXGZ9Jy9sNcG7jkLjgFxw2kRndXV2hZlnbsfWlI3
2oHYYwrldfHgroFAVYFK39AhFlMeemTQ+/4glG3eBSG7K4wiAaCcYBB4a6+aus2bz6bZIlE6M0f/
dwqvrB58h2h3wAV6MpA4kh3R/MBCY24qwWRXNpANQ+BLDkkcE0GzZGEEk5iNW5xJBM0frxaZlAym
4ZFdF4PG++Vjner1Vuvzf9oi0WTJcnUgIIKlysUE0rVIeWNxz9jzVm60QPYbHaCHnIcwCKYiKast
DN7mDfDGQ5oJ5DM2cDSJFBrJaAbm08Iei7P9D7OrYWh3lyi3hZ97VjGCzWeqFYm7asRejFPzthjy
lR+pLH7a0/LlhhzPIMJ6tEMICC+nN88qZpnccrDDGsOjBYiBbn6oUMhVK9P8j+JaMInJGsIQvkD2
PyJJpS5tq9SocmaeMsovm7ztBotB3ZZ7mO/QzdpUztmmV7wxr66VOVJjWtjxmjOZn1r0ffIOSJ5a
VWqVqYyqj4HUP4IV3l96U9PTWgtekBD44acHivdUPxhotmld2L8ehRe1xL0gIaUuqleZHbGgCI3G
tDKFn7opwltxDcOPaEkq3YUdS9ZQ14gFlrXpJuWBJvNQMISOpKKn1rY1jBkJknHlN8FEopgDc4Af
ukN8d3reZeebHd8H7xZPuwy6XAF/Gj/DTk/0RKY8VkKC8epf9Ce0WMU863H6kiJYQuY6u1cWV5bQ
H2NcFGFWnZS9PCnu1XreCMm77wLeQaSeaxzvkjoDGER8BD65rftbW8t5s7sNGwA/2WTxf8E2S3hA
YHH+4VtuhHiv73UR51MsqNeCtgG4WrCfN/qOtXuPVvKINQD9c8LQKbvWDKjgLWbnSsAx/lD2w+na
MJszcNBPKw93IAs5C2qV+X4Oy9Q6pXOSTLwC16rTpis0Z4G9Lo7s8zkak+GLSfaVwKkt43HHYq8k
kawv3n3IjIDFTlIKtssHlNIdL/Thtw2V2f4CmUn6ss+yIVBy0ugfz4lfqQIM07nlACdcMIeiM9SR
mSbJHaanX4ATQ7KVbz0GsqiVrh7OsIxT9twMlL7HrbMTb1rzHIuu0MXJkHMF7V6kPqJlRgI2mjRW
Ww2Gke+lupoFZm8QRblYaIOfvD2CbJdBzaK8o8p9PnObpnG9E/Lczbv/OgQ7T9s0IYRkeUL0Q4WI
qDsEnblRPABofd6kHw30XaHjG/X9SFflhtq/EKXrwSBw/RVeLxeqsf0sJyz73OiZ6NEFcp8pFfdH
FU9mmzbzgF3aXzGzt5pSnq1bM1Z0P0Q1AY3kvz57K8P9mAUVIhK6iluw5kc2n+3ORbOrNWhjITXI
Ri+QTyUeOnYbByaDPn/r3Wapd5kaIJA4+t68Q6LNMem0WQ70Aw8eMkW9WoeCRIY4u4fxVBbaERx1
CyLJEtHmWtQJ2rWtmwiK0x0Ac7qxY9qLsR9Hf72z/85scMof0pvBpkSuawyu388rxBFvtqqzP8vw
3HQqdfZi4coN5FNokGZgiz//38SS7WJ0l6AWLcpfsOp9Fsiv6ZkX+Cc4bcXoDWLYHhqOBXGw2/k5
58w+MEUsGMqiLHhYQtgolgUriJAV9r6V4fZH/idOWk8XMXIP/DvjaFO+XeL494kncf6DykOf7nnq
LRNfue2kjx+/A4owzLGc9axL+II4NY678NRLzc3UgVRUyo1xQdwmhQKvw+KTQz+D0RSZ0GaZe4fn
/oY7KqLIAZ5DL9WC6Ia4dAsSPMkX9UGxqRqm/L3o+KxxraxYWbjkY3xmLO3V6YKdxXNlOGyd/EXf
7a4UrdlwNNa4CJXkX6FY3foPwnfqIdi1vFA0CFDNFhbgxsXYdXvgw3Mq9pCZ6Af6ZzInmfmPaLkz
veOBHRmWh5o69GphzybogBX0Kg0JXwskJxlmVIMcFOQj2kaBWD2bc4JFBJQuUiHKCrZI8Y6gNxbi
/04RE7aRh2FHCOhMf7CmeUPVsjoyzHfxuQ90VGecprhRpwINidLzmiShrgctoN4ct0HRAGQ1Fbml
iFgDfnEH1jkrGIn/8EOKfYOx6gG4mPPB016VVxDk5Jr+WYMo655Z2NTChEWozWdTQml3252IQdhW
V7bu9O4ICc8em0ZluEQyXXeoMoMawfJcgw5IyFJF3AcSR0gZBooRuDU299zkHOBT3X1GQbNpLuOz
OqzwRH5kFr3VFZUqH6FakB6OpChtM708YRsRhpsiXm/WcB9hW/o8XWza3YLfyiDet6VLwJRVoZZZ
grp5PEE+pW5r6cryb936hH0j/Ar9M8kHuqMnTiWoNyj+jrp20ODLfAA5AQ+5ziQYp7Xhi2X+GS2G
s3iGwBxB7BUlc7GOyRYbDOSBZU7uZKvyR02yuVdf2jv8V1KIfA2sheYgX3QY3eaAaM39M11oKA4R
oEOYvp3e5uKr4dctOBE1b1XvQBN6xHPkVkMZ/aXHa4ekUCXQn1M6jbIUIiyWUvoS+BjxX1RSwQHO
sPkhWZZkpSDIfl3Dwj9MeBHfeWJcwYO3F/ljsEKxiTBoaUKzoLXWNoUupuYRjg8f4hIOFEW6b3H4
SkQ+/IcSnwq8KyDGYdvWRFVDRRcb8I6F3n6lACjRM4Zl+8Rh7PlKGgORqf1Yb59Yb62HHi0IL3l/
/iUOIFfH4tAIiaKmNLdmwbUMuodDyiv681f+7ObidNf+QCfEU+N61s77VE5T0LxZrMT6WBw5Mpw9
6b6mdQ755xNQ0eifiseJCofauf91R4vIIkXf7o2K6dFYvmL7ikrobB5sX9HD4rCRKbvWtLJRbTqw
sZ1cUxX6zAs3pnrU4UlO+79uVUiBGJpXFt3Qcpfvcfh+XMQ8b7unfIZ0btW4wxPMeqYWzfi5FRRv
UA016/2C7+97XZkWefriHhozc9Qrwc+VwRYITxdJmalnbCilpJQOZjBjgUJTm+5bcn20WqCFck+P
5U9ajwS8nqLNqqx7mMY2tU4Vko9FCKl9TX7MQEdlA3PnvuIP8IpEN8LlYPNR5OC+WWNIrDXpBSp1
NfFM+5TLQHTGCxkjASNQuRnKTEGmGS4ovXWRTJ8fNuSPquO8Pz1AipxEf4CYTu5WQEip3aTadiTQ
vxiJ/ZYU6uddQKJbqSnW3tJnepjiYOizkV3TLAEFxOYtufy+nQoT2Ej2RcC/QHR60f5qQhqqqRT8
t1hxt2gTYRPNeswLZNuGhGXc05Z83l38AWj6vjUaFa8zlufqnXuIng7Qwk2ekjApXYIxRnVZLISW
TQvfy7FbG1siVn3uzckGaq8ljG/V1ezpN2sqKJe+lmCx/I3aIXRGpOkihYry3KoP0ALnxFHtMPAk
p9dS/aQ6nOVcq1yGV2aB4HjN8YxPDQMwWQHQvjlcWtXNgZJ8/EUmvy5w1sBBqp29bac19rKTn3S2
06yXy9sHErhEXvgz4kFgZ7DRPZntKf72CLAacCssf6gPb/IE5yAbcCbtJ3lOsVSUN4rGuErNiNYO
l/2X3rCSUOZ/m+XlsucAQJwGglZ1ciVmtoY9eR/KD1uk82hkKbkFx9bdy/D8Hcln7e/d6JZGjqU0
zkqZjajr9VZwnrOrH+NsXbKkYqMrirNOqyKDaLwzt8MUdNXH0yS723ughctbvNWeO6F3aBjN37ox
fDvWDJ5eWPvE2D3fymWj6ts5y/ZZ7hP9WeFrKQ21BWW5zXOe1dd/5sSvc9nnwugbFZo6MVpjUzdz
4Z63BvVZxlnGqNIeRbx/4ij+SbkFQbG7RFSWhq83MAELYjZC00fEi/ND8atYpwcVLrqb8fM6u44T
YFvfI7eX7dbuqTLAgGn+e1+/w1tjpKDFXJpUMwTWdWDHsbIeYY3yNH/L+JtrrZHPTqzK6vVRcy+A
4m4K4S06ekNCunyng8fCaPFoW0L078kxwzxDPyp4Tk4DuABibkzxdeaPkCZOmhEnOAaA1chuAbdm
dEqroDvq23aCnelclbjnsyRTU6r3ppBEQy84PemQ3hw7gKW10ScrfXlAmMuMYSlo5/ndoxcWurwN
d5h6dJUwNcK1ZEA7aXG40kYt5wY5SaaQHF3mONCXsuyE827hTgMfZFohGGNnxCkdmttFnXueUTY5
6OfUvs29udpoNkdnrbKRn7YZKawWIeSSxUO4t5sELDF6hxETBeE4Lpv/rUtYPkorwlg7vgXCyyW3
EdUwsfXmR0udPqKKtzNUMaaw4xFLQReOBulbv8o/xsEtbkT5nC9v8DhdhLp0C/o0VOCyiSN9GuUC
nEORoeVU2qiXjIWkl0DDb0fKIa8AVpVJu84pPmA2F7feb6POAbs9H79QILilAjyqZhjireompi5g
ewPelSnMHyt4JCGZXvIEJltQ1Fb7zsorNvaQbCP3zJ4Lf97/kFsumOA+FDRoRI4ZzwEbYN7pEV2K
X6EgHXBmyjbaO8kspBKJZ14rSQKIwm4ELOCSIviZFl4yTZei279GVcLIBsFc64FsUL5XBG2+BD5A
gDaHWtw2oSzYKHW4unNDfqN00NpB/ZXaIcbCVp2crG3IepEpSyYSl85+DJRqzz0K7qnye+nh1ru7
pS7I9NwOa0FUa6bXgRxInE4KPymr+H4juxSTUEPHRPaJz1pP71JJeDhXjrehYWLbd8Q57t88kyhf
exS4oA6GkhBw4y5T+lEj4qb2fgGeFQAsJNDjPgq28w9038bIq2aKzmPnUoq499qpBds4/n95SvyC
t4ZowsN5Pen1GDFmBWmeh3AmChIEhkVzwhZFn1AafiStO0il1oSska1T9x5KVT7HDi0+Cgv9TUCc
UuIZc5MFO/vVEO454jxj0JDpnDLTX/AMV/iBpniEnMSclutp4nadyF9BnWlCaH1efFb0xIfRYQXV
U04WF9bovoviog9Uf5yz3vBoq3e2IgZG0mkZ/eRZ9QLtgi6vJQz9LhK0Rg/yup/yXOCJeVLAfiXW
L606o1Jg6OSaPHYLayTNFkUHQ7I9t89jt2Mavvqehhwm/atgvZQhGdm/8zVDLOQt+3XtewlQ5F8m
e5VhyVOOzYh+WjkAeHzI0R5wFlZT3pNN+RoFucSaQDiZvBnw3SmHpMo9Wi2e3ZNiQigEcYjtetzR
jRi3rAGV7UpnvIuT6EDU/Dn70RVYy5GMdFahhBQpvVQLDzW5P0NJvCKd5U0mJUsYtyE4DF3GgR1l
L4GZ/Mkc/vrDDhxuPpcfofkcXM2z/ablhoPv8osIKGQJCHUPSYmch+AGRgNr2waRNwCm4d6l76Os
r6Yb81X8OgI8DEYbFuj04UUlj604HIhc9Oyppg50adwQUCc8yKtaVQYnr4kTApoyQ9VKqzdQ4LnC
f8372ccGi2iJKzrnZyHAIsGJbjyin7y7sYYeL0VaBoZtgpjEEP7Iwgmf6JGs0EWVbgS/RMV0Tqm2
UyKvtG0L6ihKmkRdxUVTOz+3ZIR62jTHcCpntkyLgtwvnmTXuUGv4ex2WEZqoGD8S1Jas01H7lmV
e4CsvfRzlzERTwD6wF6LzkwsJ6qpvuopDXlYH+Q4iry8KLQFw2KGZBgajK1pd6OmxfVmR/FHA1g6
cOwie6EzRZcyORxFl9iWOiOWjRbzOY6vB9lCeNDjW9ZvM9nQtVMt6xG7KTMd+KEI6hqbEMsQNKMR
OpqMrl6BQteOcl8VWVegPmaG1i7eZuvkY/MDyfxCKrk+fstUtZEo+uk79JrC4Xt5bx74ogatvi1A
J7OoSpdjYXRwSwDRcUzuR6lONJc7KKAYyVr6wMyOu5Qhjek0hRfqd937CUlr/c7sAdNaQTlm6LRK
ixKpqPQ+7SlSgPr4ZmGwHJLcOaXbf3HjEK+HO6ivt8WCxBq2zt40t3Llh3+1ysIoR9XwbdM0aIWt
JA8/Ujq8+5FUVqa1EsKijmB9Rrl4k6yKme7bSJWB7deBIBAd8bZWAM/RdCXLBIuuCzTnjIjf4OQP
kpe+2Qt7wGSBy7dp15+JyrufqweVVHYq1Q0Sf+TTlEZ68NKH+CVZSsQYGredtdvA2GCM6VaXNBSC
NY4odgda6uMxX0IFZagRFdkcaoc7PEEYNId7NEc1uetYOgmVSfY4KQukOX7rlsopos3NO2bEtgy8
D0e+n8KCYDjVdL1zdqW/2suLFrRQMcnQSeFGgK3NdhJ+p04MEbuxUtqqZMcOpaPu0Gees/x+JqU6
niAfKMeZcOX86/8hR1qgGxe2nrCK6mRgc1T7FPVQJ4DmVOAfX0i1fUCHXaUg+DelneiYu18ehwS6
U7jAwq52LmutnVYnn2e3jMh0bQ2jnlfQNBtlfnW3KhoAXa988pZiXwnvj3pgcs+LkAKniG0mGJ9+
R+samlFtWjLegSceJRnQUrA31xd2L2tuPigpc/XbWDtraJUoFSjzzvXXInGDEuPzbp030lE+LnIK
mva3Fio0mJHPAsEm7R13t1fcTMJBDXx4WAv3ihwt8AcOQlAYNj1ilYgn1OzGICqapbk5nVXo9mIp
Pqcz2FD/40/HG60DhsrUFKo9WCAv2WLW5hYJsf9XeCYe7T0yJK5YLNVRMwlZ2UGV0m0zAQ4THLf2
Ui82gMow+ktUFNaRwSVn1Qn0H+KerpMmty+/pJ9RCHDj6nIe4aDrKVtrmI9RkYshjkwi0fhDvSOi
oss26qys3v41RN0sLA7PglLsVeospJ2+iIf9p4gVNmsjCRnFyNwwcev7jCpfe3cViJZ1Oy2hWaWz
6Qo1FcdHpxkLFNrn69/eTfHpLsPwIIvZh4vOqbJujVBvFtulsHFqOZypPAhOv8XPyMOVuHVyviNO
2U4z1BbY8LbL4fLgyOtx9liYJsnGahRLNPn2OW5DaZXVhJUKSZcOdtgh92TbtRg0ydnTD3xC2PZ4
ffmG/waJlXhj5Rz4O7hz+YuREGFoARv9LNtziTMHwi8ihxlOI4pdUTB9D3AbTxQfs/48cbPc9WzB
/n0sg/HY+LtPOqsC65uilnei5SzUFmNt1xftwlqP5ZEw8asBMH+DiSvFsX5/75Fm+i0+IK0XD9ZY
tkQ4D09k91E+M4MjdS8tQzMJ7pK2Ly8zdnVA0VZ2/RAaixu8rO6ZugJuQEUnm5ysxt8Z7Dc1Pb9N
0QUmIcD6peAEqIdxHmFAe7Kr89sTy32nRkUcfKZoM9TJZmWGI3NOZyoIgi2r0LW56HK9LUw2iaCW
bsuM5FrXFb5M6eeqnBYnsUGWuiiNPnFFbTBkqrtoh278o0pE8lXvstrC5cq0BRn2MH+CnpwYh0Pb
F9gGJ4kW3O8yjTZiLNkq9flwQAvuf+mrJGWOuL1RXONo0ALeVSvSSyfjZLUZYj4GrLRPPiQQvzMz
Tycep9rKDHwH4pKomA69+0yoHcfIsaypkB+3ATuGWGnkyV9A/hNVGgOruYMugFGAnjLzibv4fEdz
FZtZBrdrvOVzB9dKLr3gyM6l9HHAE7mfmquxCb8HPB+3fPIaqpfp1wgORtQnjRXi/qfyZJk4gYL7
jWPjmJiR4VZ442vE1+abLjpF9tLsES6547COokVDXGIO1xYwS3QlYMXfSG1KWkmoONdG04O3mUbI
8fgcypOiP7asiprQTJjMn8GH4TY6RW7VMiBxGM3+mayIeeTQj4RwqCR50ZZ3nk/ztn4950FvcM46
rQFMTXiYTWAIBLHhs0RgMqU2nknFKYqs+EA14rsrDCFWulXqGiWWVRYfKdIeveIBZ6/npAdS2HjH
Z4syIfOGrquDHpT05ZEFUA7vu7WRY8ZA+ti/3yaYCu4V1kKxr8xOHcafpMY/tkUwy6Lm+KpSWutZ
n9SLJ7pRd7XChk1a7R/YXQg9gsVU5p3FWPpCqkSaCNaq7hS7eOgcWbMpzXexenuYHtSTeE8N11hM
FYxnUeMBC8Aci6je8swZd2xfu/T90CrqDkMcwLCNhajABhxWI/OQY+dkSEgpQo/uWUwkjA8TeM+y
gzMUIOa4FU2jK9RSbgdFiO1U9kSjbSmzCkigmucpuEzd8tJHRNLkw/f5xLjV1UT41hPVPBH50Lo0
7OS5m85h+9x/qGNijhipuvWqByfmQw6lRAbmGjKM/mX+TmHXPbfYbGnCAZnAVVngJIdKTXBqSOl2
0faPS0HRG5zTk/GsozLXIgjEEE/WZJaWj7RwyMN9ikZkv/fxOvLBJkjsXQ03TWDQD59TKw0Guma/
vHKpqkKOvXPS/qPnZk9qQBClDDr9jfxrxtUeMiVR7QbE8wrwLhzQRXaZvIsD/5CqUESJmK8GsvN+
zTzZHSrQdOdg169ca34Yv0tiogWx4kLZwADKQh593puLUyuwxzvyRdo5gFiJhE4dlPgJrsV31zlY
CvavBByM7zRZFX9Uv3OWb9SMmp36ssx40bL9j8ApwBrDIg+T7KX5w9UGs8SHam1bcZXMC75cCVDi
wN26EtlNPYUu1noFOhnhPgIN0TbBV13x28XVjP9CuFYYj8kRpKAeHAnXSX2DBUfxfBwhHKn9YhKQ
bq+HKZr2nAPq1kLZp1Xw/0ZQOLdM5mAko28x56e6DuEaaenY6jmlPKNR31r5nQS71N8wD2zjEa6U
jG3Mo+CZnGGduMFRYKDNIcJo1b/szZFiH8OUhsZ0P79RaU6XSdRIV4U1/2lBRSufDKRv49QlzYdl
efdgJ9KY2m3K4uBn45WoIZLsSpdkwLhuVpM++zeGnKpuxnFvijZ4SmLebQXyFEF/wRAPKSLl0RbD
hUtYzg8Rup+NDkXMLFNi/Mck+aFrZYsBVy/QsrIqaW1KpqGnEKKLAT3bB4zpVv5clRP9y2K0b3Sd
6RvM29TJMN8Gh+DCX0KRyDr4eXogJlBjyuvZrgc0pg4jhry2PU2fVjoNHLAeHvv25PVOb1C0BP9y
Z46OqFiHP925FBxkYc89lqBvbX0G46fjyL+UTauPpcgLecbMPkKMLZuXOJm/dqQ8418u+PP1AqNZ
S88OyYkwpiG6i3Y9FyHc22UzQ3sZKZesr87Cls85cBU7TBrhu4lykegWX6BtY2cRxJwpfdcyRatI
uGh23xuKB6UDyhHKYu2djM1oZGWIhsdYEToHt3u61ad0sNZ32HibH3J5r86u8B5JJBqvubIeADAF
CW50QCByWZWVb/rH35E+SK9+O53tBE5sUwgIFhP6eNw+DiZ2wUCE0z5Ry/Hz+IXLqERmDfayyJiC
tI1DSwm8qiIaAAkTh9qeafITiw9enNmpJ23dL65C4o34P4g2LopEc0v8nAzdlvc3OeAR3wCETgl6
82i14pkdthMnDYaEAakGPPTIKqx1mQUAIjk/2CgEj6k3BKk2trl2/otujH5CpSaUwL3fnaMBO288
SZ89LWhU/anhtYL9qJxbL8al0hjDMLWbHsi02+grBC2fBO5znKHbjQKumMVoZDkzeaSNrlfy7XI+
yYvvqgcIS8y0LsEGb1VaoecBre71jkqb252EHlBZUCzopeX2+FXbnciEUjrT6rsJD45HKSB1P3+p
JQH9MLiREoS735dM3pwOmWvytu7nXPj3tpvAiBQ3L9F7GAXTt86OorCAa5KA9RI4Sba4wNAjH8I1
3fyv///RIMNd0ptS+pWJLufHdQOdeEvp72Hsh0KoTwOheERTaOktgZvNQQxe/1kgi8MqQRcUVjkv
EtRIcsSyjS2HJAsZ8GOxLGw4Hbz23apoY5LtcjjhY0viLav2CZdCxywczVbWv4Bn4Ezyeq9H4G/V
lKjB6Y4whSkOvxd5m40OFz1UUgdWbJtW5VSU6yY75+PJVaynEJhHb9ipqSbyLjq99ijovsiAty3D
GpCG42yK5eT7nKXW3x48q779H/F81WUAMgFwQQOYWKQaeTVCororkBJ2wKiES4l3+7w7tV7XYuRk
R8JhYb6pYID/lOstvE0l9zNAhzar8cMCRGJmoabP1958LGatjhdCDwXSJqWBZEtfHjLXsE789FSr
bq2Q050Pj2Ua2fl2b1UaCthf7Wk0YvD+4EIl/KnAUVsXzaVdtJcBDzPuHeYvrzodOrqALd2OS6WT
8DjxrDqFcLhRyrcWWTh5/vMiUN6ycUbDXcCrUsqLA8UpTmtfUxl/9GoMTnIl4Dly1xBfN21nR5Vk
ifCXU4QoESiEisdfhIy1pTVT1WA8nPUDptQFgsMghkYbitu8JIlHWit4lnFAT7BRgPdVcN9MMg5x
Hujg9GRbmHWpaSuSQeMGH1qgPtpaJZfmdRpP0hC6lWnDLhsGZdTnuPxTspQDwMBLRUxddq5AC0OX
YJ6yD6T1Wlp6MOgN0j3e1jZrQw1ZBU0tEsjMIFOekhocEKrR4urElX84qth2tElRnx6wk3gsmlWj
vvqNHjbEqERFd0R6qhFppUHzZFdyTPZxhHqFl1eYpxmaLTJ0M8vwIW8A4+NSmnwuEFTa7ow8MvFX
fuY9jgBVbY/iU7rvYrBQ36zXOWxmxmgJIDW5DOg0n3r/ESUDCxhubbPX8bX/sstj4J/60O4kVwuS
ekPhGERQsIJ+8u8Ybc+0kGZ8Mt75xVrpMYZxhm4R6QywrwbN9qv0JCqPqQiytUerbphihzOiuso1
zHpc5Aprr2zxO+eAtQPYEEMeBGmXnK9rVaizxBUphBy2GdFEU2pURZX1YlMfhaQD3lYfOSULeQwo
XO3XOXBYTbleKVduLsIbFCDXV+AXs83Xb1+PJrjyIG/qktq+9QhkfGRUwnBA6/AQVh7CUyXQHPRp
ty8nkHtD0FU/8Ndr8avM9LXlQtiYcqBgWKRB/wyXibwcP80jxMNsHac8dIYJ2AkrZ7wpw/rq3FoM
TcQzX6X6uEx6AJVMnKiEGaP66FpItz+jaJ0vnYZRw4HLBCvz2X+oFEOdO53QaqqYkXWF0ClYsrXQ
dwKpJUqd1lk6LDxrTBgtgRa0ldW0CNLN8lZjsyEG+I1hN7RmCPkHSJy3sVTKKJx4Vo3fk9QzdffC
XZM753TtibJZAYlFFFtMk4hVpaegENkZ9GZgOxiy80APhSMpevWJoVhgNouCcU3DlnhvnTWYh8/j
+QahRvjM1jYDXoDR6eHjzgFSBGbPnqJiR3y+Hyd1axlyGEcxz5+35ZZTItT8y5i3cfZfySisq7Yn
xMBJWDbB60Ihi5jv6F8RgIF+ZOVjCa9ylwrotR2aYdR39Vp74LHGurBaBy37K3s4GTVHv2oNpAXS
i0UxmbEQGISP+WuB1VxfFVIg9Cdu8Q68mt+H4xoa86tTSn/9ZiN7SLnpoKGMqNjz4nVKqUf//AyJ
O9I20xHewtV8oU/BfYWfiOnRhNFdUUwBUUj+8LmLhN16xucoOtIrF2VB5FoiO/q3DrVsQVvq47bt
aYmedY7Jp+6FhJm6P8MBK5Lgqq/YMsHAeAyIPsdVeLBt+U0Ga6u6OxUk38g2EH5XQ/bQHFme7tPE
o6bqQocbHI2wlGpsxywkCbDMkfVmojpc3P4mL23YCg3laL8SKQwMuJWM4sJXGrIUlSBdZXQvN0lx
p2jeoGw+AClMCzRDGMZgCWzhVsfBwndyBDrmnL2QQfWoT7FGQPQqF9tPhoDn8b+UbEhLMEfaHVmc
17eQDkRgEKhmSA+qO4alOdkHNJxRFbr8l4W7AqXSV4fz2X5D9OHNTAE65zOZxGUfLKP86lUzuN0J
USygmVJbYRpgabOuwijiYWv+494A4QLVSZmvmP1ynyiEkQvbBUgvQFOKgFEihy9+RzWEDMbH9bOg
R94KHmmd7V4TZ+tU8jEZlK2KVg2MvdKlSoyPtCTy5YrLhiCIrCZswHdo5aZMkfaNiA3S9+7QWrbc
K3EQAW/03zNe6gP7RVVbc7q7MSKPc9qghmnEm4JuAoCCpW01zlr3WhrzHxpJHh/APRw9hN3oKMmG
Q0pDKJ0nNUgb+klio7BgnOgnCECPAYhvtf93QfRv54ideRqMJ/R5SQl7APeaVubKF+g3VVQeTrxb
U8UTA6XDFCuAasqOhfvQzMwMJl2T/M6cpJKEB+N69YPVXGNpStTE0tdq1LLbGdpb5AloeTxBHlUU
cWaH4Ol/9kCwVIR/NDzy4VyOpLFihifQ8ik79HNgpUypISUME60rYwgImPMe40Xu0IhJKnXdK6NZ
NGu/d50UY8WLRuFZitt6PZNbqmP+FWFx5IqDfzi7F4pF2c2d0ch6OD4XYs0WYWViwZunpSaGRmKw
HQtqkqUrkLBx7/j+OR6KfXC4cxu8hpN6pCI0j8VJvcdzuTR9hINjyfH0u7s+FMKTwK73EfsEfpYe
bJzidpbXWklTr23ubj48ZfcaLALMLmk+pdcke3+bqckrAubQFxd7/vlRA1B2bBZ00S75Qvw2zwgU
6QoJL6CPzNzyTP1vPhk4b/p9MfYIBzH7ZkTEY8Bdon9BcfRkZgQHZY9TAY/h61fKJbS/OhZTyrsP
RbKE9Vr7gt6cdZL3TaFA5Z1KWkSeHREe7/Zp9Kq3DX4n7F9NIVcvQbxkwd8z0b6elB82AY7Ub2mi
ik4f6ioTtr/jifT0TvuKLRcPpXbQiqOgtsWot6tA9tnmFQYlbtkgofeYzj1FrV+h5IPvTvWXPaj5
SVOEIXgxZUuYSkm7kSbvMfOD3sZzX+QCfSfZhT7KjESF3Ke0irdKgb9ifO4rleIKESegZCNkCcnt
XptKZ8eWiXvVEU88ns2uc5s5vwy5MpHhiuqQ+Ld+e6lIPvbAqxO9uYVmkfJoTyAMtPzXh7/tDQwg
qgGSm0NDsv8YdKoipESme2LnMHsZ4GSsyHHVbWlp+ZaKPA1bGzDMmNcymUnrI5NWYoRyK2kRR5no
HsCpzqOJ3993ylk906j5GelanB3Az/XzklbKrWni3Jtwul2Yj9fXXPZwDaw7HYEQ9Xj2bEQdwAkH
Wk6+ctxL1df+Woa+afIfh8GskHwteMoqK5iUAp99XMh31prYH8OC8wHGywuZQDny0CAradzFvOEV
5pptQ4ZJw0pwL6HQkGwbeCBl4+KdNgUm9nxIU+M4D1pZXfgUtRo37pgNL4LPacgBviAluSbQRlUu
roI7qTZdqvgQDjPvcjWqhcbd0hWIv2XXofwU8c3Dv4e4fHUaTaaenAbUxnvbpanAipw+Dh9tQZ7F
21L+QmKNSEn0w1WAGmCUjiLZ0hmOFV/+x7pNgjmb4LHtIRHX2Kwuh5WGzOQMnYci0fWGz+QihgAA
hVeqVUq9FxztUUIpWwvJWpUqC3hJ9ckEZCMhQ+kn5GCeknGq9kF0kFPWKOtEJo0zvjAd9iuU6N7e
/zTioOVJSY669pS9fHovQWNX+KNzb6IEhhrjZhpWlPEJ7ydGd62og6GkT8+mZGD2M/qbewgAIkHu
SFRE9FsIHwDPzLIw5erMjyJ+hqepf5jX09cfuwoesMZQolbY6dJ3X3TE9YCgU8TNUj438zCHCxdW
Zr/MAmTBRw/ZSmt/p2dDkdo4JUFTEFjY9RckSXCpDyvcZoFoy6ZWmedl+famz3EtOWxE/5wgonZk
JkYXeRgWbl8ixFMXn7NNC9onZ7apRS3IQYx/1fBvV/lEml9mv27xTw1gYacvchmLH2EEYZWnAOy7
g95QLy+GiWQ5yQ/4p1mnipXeclbZSPfPSdN96o5fDkX3XEqWNaMp+yuRRMG9P8YjmF2YZkO+Duvt
fUirnjEgT9qQJPR5u/CAxW9x0KilrxAy8A0BmxXenG+ZSz8dUcDw+Gq6DUcH+SSnE4NJMqVPPrVF
EZ8UhgkI+jQ1gO8lJiS2eyUJWN8KhfwV4lDkXAywEWsUvqp75jPwgqtLfO/RzaJDZI33lcqwbW8e
03LLd1IVw0SYYTlpE8jn2B76o5VP8CxBucOy+8CNXtn2jAV3LMlbmAOK0FlFRWa0Dsh8HGMZ2al5
4ugFfg4O+oWqnLjTOZkIs7vCtTVG2MU5YOwVPmpCBNptls+Uzv4Ja/2wuzS/cEmNx4ZUIHegIFuM
T9m+6n6w3qBxLJzR85jxVkdG774qkcNUS4tnBwuEbYYYR287wJwDW49NJk0osh9s7qbaMx5o0A91
4PBWJbAXtBfAHj94Kl3uR0kvmtJlm1b1W8JDA5Be4VFpFFE3c0GTNY29AbsB4wTsSjOvGrx0mJqw
mcRsPaFmM/fbK1q2tUpc4q0wf+lV3vxjtePsduzuvn9xLx38XReq2HdMYJpbjUa5yn213gATbORW
Z6dWJqXaurldq4rMpRBrh9kEMXJnz3Q0EjDeZqVJzcyhjJcNhbIz6dJdMqHbpssxqryDjycuhaIc
aPwOyMADHZEyaHINTHOva9kmPPqycinryA21TmYin6hlK83kLm84Ot5+nKQ/h0SRj5wJ9XFf8wOy
pT6DDpIBp86+Ow1uxYLgpEku3d3iJC0KKi4zz/mV2ML8Lfacr/69j+GPTvd9rCXo39OYY+1UWYsK
sl9X7UFoTmyfz47L4+qbNqgs5PfUZPCy1kLttuULBHh/TVOd/WSJg6mihytCjEGn5CI+lAYghad6
HI3sebI80rj3Zl/Pqz4q2h/IntX3XBKXgy4aWjPO4+pbaTD86cU8K8S/tv4FATUyrQSKnRMwBQXZ
O9N4Q1VYoe6U/Wl3WhlyISOEnA6myqRCeUwO+NYKwzxiMPiNEytwN18o2QH087doyn+w0zknVZG5
TdUZZ5VSVzNI4MOsI9Qm7AnJS65dHV9rnfMWruUfW4Ui2ptACdHDshBNrztwEzE3/TyeQG5rFA+T
sM7r5Ut+huxz5VdHF9z4Et7fBdMxIrg3Vd8fqDnxaN8J3SpZSmHtDo6sbY01OKXiLKOxnt/fupyA
XYzX8Rf21TyCL+ruup+Miwh7HxUZ+GqphxSbtY06fdgZOriYUJ0VJAhUV9/0OTQfa3vafxJohm9/
vhI7PE3nscCFuEbYD9I5oPDZulrnzua14OOwYeSPvK+ChATCIPp97Otrr8pb6JN8ZTB2TgzSsSne
Yzz0HQ6Al8du3hA4q/XiFPm6rB9PRhSdJL46ggiviF2HhFD9bP3nm685iSSGO5sXDfIHdMQOeGF2
fIMTKTC+p2UEe6FocnmeakIuSWL5cQnWejGR23mzzujRwjEtub3LEu2hvMAy/v20H8ADOF6zFpVc
z9SMaGvE9PRuy2ik81vxLpgc0AA8FrUILrraBYFDKlUXAIdIjGKjrO4iD8NyuYqt5T8P7up0GsP9
1WN7QGyiKDBnj5Zok0pmT5rj3Z9to+QvSqoPZrivvztrdUPcu3SYrE6nmwBymlf9N+oDod7g9cvC
TyF1CxOP+4VxOpqpd84a9TzgZW2VwoJ+eIv9DgnI5xgN8wxXfPC8yUHUI7heEQ+Z5mmlC1ZSk5tc
qwWORhjMQ5/Bgu7ltJ8Y6ubGrPowiBWYxiG4qrNMEBDa5bpyWSqZksTUU0IcpCnJfhc7vVVpYn+i
JZytIoa/UU24dZdAf8i7SI9TgvN3hkCG89pflE757kqckVy4NgtsP9HvomS9qcgm+MQVkfZDb+wr
414GTHloZnk9gfgrcYXBchyKyUOUFaULqy+tHc90Epjm+VfKA+B3X2l0GYnON1vsqeJCNAvWE8fl
tHfkpcsk6gNNYSkm2lD5VFjfVskPr3V0C5ZhT6PHAP7vpin1xgWKLnsteLLXaPR4iWh83exfrvwS
7Tt7y1AmKk2k4bxyAS4hN3BxX2U6gDoayuO1gBwElRsDtHBhwqAvigIyoNB3ngMNhAVeIAYIud5I
vuY7hAM08X8Zpmms1HmCmYIiZNq2S/xGB8Kxti3kBwht3DCzNh6N29CMK21qT9FoAftc+9ABbb1J
7gJuQMvVSHSoJf9p1J8QR1skTPJbLKWXVo/Ou7JpIwwgONUX44MetfyUF3UU2DA36uRgD03/qB6u
HnZwMD79JDTSZVcXhbGUvseDhH7ZB7INHmARUW1BWo2zOek2UbZzs1fFGl+SpXCAlLG5hU8ZjlwL
8Dsd/U8Fm/XcFkZF6QzXAjvruMx2v1m6eVYEaH21JAQrUPcI8P4MwSxE4wLEqUrrsVuEtcpq+5Xp
yN5BJv3Hp96NdRmvvRBqMN47ZeiQ5VmWQCr17X0jtGkrykHgoqtdQ5wwsmQ4uXMe3SLN1qaJhCKQ
fg4yHkM4dCgW6tyZl9dy/t++NfJapU+8AkPVa7JiE8vA5WVkpUeJsXOnpxGpjNF7JGAJItQnk1Df
JMvvk84EZr6TfPh7gPFe1nDsRTbh16ZxxcCKEOPfARxjeAW5j33rzt9Gzz0HRsW0uDSebJabh4Qm
jcue5s4AfnLMOOTutyuMmfS5BuaisHnJiTWvGqq6ZY/48sMOvr2qmavmSkH7O12MkhVtt+6TFMz7
1GRKhXKcD5iF7fi6of4XncAZ+oMkS73e03VwR/Px39s9rp7ZRRE4sU2BTFcldgNPEK4WOhQPhjOw
uyGhUvIoaqG5bk3sN3Go/TPXwqVR6qBX8lfo+/1qUzx3PGwMJKuDW3KXQ6y6iQy+Z+D8EDhbczbL
BnNJI90zck+dBjq4ojSeMp0xf1zOpH6udTI0vJYFy1qexxwaXhmEAMJJECFcJzlE0X4xjQ0u4fjR
mupgYO4YZvLPJheQ8VT9mQWyY6ELKo66xtIwK6I2pOMN3tCHJLHZd4q+XkOriH2o4eVOk51GzoJF
ct+JoE0Pbg6O3aDymvXGZHN1rONOxIi8olq43g7OR2TedGgL7At5I1zSP+zWrLbO0SqNUwPH0FZ3
G9ko68ThVy6feA2rvFSdvBOt2ty3h1KlNXIcnaJSdXPm7mUM17ifI9luRSP3W6uu0lmLsV1nku3Q
xESy9+9zB2dgX++k95JaG/6vE+f3jZHYf1yYex+2j5gi0WGaMHmF/Dj0utXIp7wFLuCYtObW/HbV
SXfX2zwcAuj9OxMwFV76PysnuVDqmGQ6+rFMHwupRWI7awzXxLyWj6sADoHhYaDNJ6V1wWlXPIFq
ifN7FANmgSlrNKWKMo9+aQgPO7kUmoopqCq7G7kOU0zz4oYmteAJee223kAwIoEvTeRNy96OWIWe
ENveC/fz7bofEw1DEz7Esv9Gh6du1dNfTrHmMZhZtIYMQJhrGw9IeL0qpknIaXfGwl4VonKwCRFx
PU1vPO5zx6q8FrYcAyLSZIXFlcFz63XssNd4pLsW09/Ivd34zryDaiiTszp/CY1XjUlu8Nx4R+t7
eswl9bbRvoHTigtpgWhiveKrI4Qzi/rffSpiBk1pOFM7+6c8IdKUVuEg3TnZrZjI6Seha0agl6sp
zsadOYM0Izux4IT889Lm9CjaiGYCLlQMsNoPYc1U0iufrSwGcm0yZbNspr6GGzmBiZcKKa+KIp7k
yyo/Hsn0Of94AvfpOzULfDArhBQbwNvGiDbRhkBj76V6uAS5UumuXzMJysSzo14+h2J6IgcphRkD
VySLkOTTsbKciG8jC2V4jvQumKSxApnfAjlb/NQHzBgNKJMTWtbWtMdKOfkU9f/PXrZc6+v9PaNW
FCtbphrg4z5bqXEhbwRHLSK+srWzUK4ord/C/l5LngEAVHm8Yo2sOPq6ZIr54d/tmOdtZ5qaO4pI
5IQh50ModyF/JNq5Z13PB9hl7+wZEEQt4CkoICZavg2g2ymFHlZNIGcYH95f//corr/FCHXXbxaV
VwPkrjdn+VSpKoEnxtLi3QH2Q7gw3bhWfdpZtyDDf/ox3BNm4wwSP1HonTvWkGQ9nZ9gEWIzQADp
d10ZUvkjBGwQs95+sIt1sYvSG887ZWpSxofsel1Gi+GGsfZNITw1QOBy7m7hdqr01+efejyiGZYD
eWkEICc9nfrsj3wdcfv9wr4kYfAWtf6ieABfuOnwgTNTZC7I3FTICdMgG8JQHdB9R90HszkslN8M
cCPHiOxOc2p+Pm5PVrl0YEAG3EZB6FV1hfA/aTxVC3L98Ade+ztsExsw01oygjfZoQiuZIFC3JK1
dye3oPVS+nBUjsXxoqUyxvo7sPqx7HztEIK1MsSed/1lKxM+cuisZNu1kXd0Knjca9zfDN2q4jR1
JnGnA2FHatdetPpbZaISsi6x7vpSjySCCrmN/NKyfmwA0MqeSrUt/wFrXSSlpj1o3uTuoDq3xi15
tzNp94DntseLklFVZXxeF626UnBwBG2QT9pQddEZdeyXOqUtWUXD4T4Cb4bVrtBm4Cq48LCw4SS2
Y2FLxwyJN9se9VI4wQffz7v5hk1hfwjKSS5Qrp0qdzHJCNcyASg+yNJlbTPDp2NCAe96WA7X0iCF
MQPFPKOj5dfR3v/0u0anOIlA2pV4M2nWH6QiPspMZGp/3st9KgyGO7Sr9qW2A0m4a2hmmSZ6DVsN
6O/c8eKk7ku+PhDeiwu++BK1TbYuROaeEEjfWb1NRt/V9I0QWNCJpzDOPWwNGfwf60u+5nBdIR0Q
Azi6z+HwJJZbc1Uy7e0DnU5s+ekke5iREfB0Rb1Zi0E8eaCYtx2917/a7nJiyoQzxVbary+ygzEZ
CWLRmsoYw414qTDls+Ab6OA6Rfl7xohegg3oM0FiFPDNx0su/P1LgaXVSko0IwZohk1Wo2ybJPyE
t8Z4nQwzyvvwozAgYwRKxFxkWn12oJy73eg3a57Rf5trcotwrZb5mGMoLhSdmLoTg8nVv/F0iKNW
s7XGssszSznyalmEAvEhrEg+KcEoLF+sh50K5FKtYptO4oTQIf+pGvYRJ+J3QGuTnxO/wWlpbc//
v3YH7uL0/J7mAA8Y0KWy7xsEUuyc2OvPIfkkdGx1Usjf0cANY3/ujOF+zVRQj8h8S68JYZNTOj43
/Pt4yKCBkLdBCKhme7zEBZwJyV8ZlXRXSKs3XwGcmNjUN4OScx6WKiPyCNvMa071RZeNvj+zX8D4
2GCXZxqDHu6XQYaMNmmWhX9KgsiAWfbWqh1uf9YwqWoKkp9DLfnzZGYolgUlAqRKC7B5k0w1d8gs
n5T8e1/tBYoNhdXbGGRmjWv9xcjrEqHxroN1gdyNFD1kVpHWeoECfL0rvjWJBjQN2P5ozCWX1aQs
wVZIxf4mTqmlcpwU6XjHDWq6kXu/VL9ObvvDCl879TrGk8kz38H+Lj9Od36/X0iXL/15MoxFMU2o
8YtBz339MrHNj06MiwY+V4g6ef3volxV98GAv/phOgGQ0ErizUtGSsTO3PAFNI1eRxL67/Y6ncMq
h2f/tnpNT3deF8K34b0l5nWdta8FdYtvLK2SEyGHTXHZKfCyDquNS+n1czA7C+q26AFRE0ZKzS6y
BVxaHBlE/KGW9ybbT11W7oC0x07tOuuIqdOl5znGq/ty0lf+iq6nM/8w62nFbeK4vO87l/5sXkx8
0NX89lSh/JP237OZb9367MVwxzLD742ZerH9iBe/tKVAPOSd+ZragOmtyf+qO2oNa2OOvTuqEst9
eJCQxGmExjZMPHdrFgRkUKFkTEzrZDyWjzw07wKMAAYX/mnSZRTjRCWeMnwO+oBbXX0PtBQvmpXp
9RBRjFJjWCa5Z+HKrW/Ep4+EI4PewLT3oT9O8hwoNcEs37e9FxeiH9IyZbmlCyDRDlvX9Cn2i9xW
X9YujobVpZqRunjEqWRTmrfVOc2iifPFvPSgXkDtcMdU0GNWfq2WBjPhqz21UFgCDYJ8twqvN596
b+rO6HmODbSm/jp96u0jVlXEtkWzukCfXyIE6Z0bunrvzHFtCLTZmwaarE4HasXX4e6Tt/Qp3SZs
OIWDBjPHt6lVLqGUEYF9onYT5KdT1UTVPbfO+r261OsvRzqTmjKFzfimLPa8MncyqwbuhtnJunv4
fJ8IXzoCHFrXcLPHr44Efb/tHatvCg+lzK0x7Dj3igzIt8fY+YYGduwNx1EZkpOix2XE3lxin4FJ
mNzp3XIKny8ol0YvqnLP5yupynyDw4bsMDvSrMr3NSRfABKxkIy9+xn609R9IWjwX33+r+4OIEnm
+g5Y06DG0ngk74QT294KSxYPuHBGBRbCA/ubmw/H1QnonYx4/FAV+tS/hha84JHlpUCJY5wEX3FN
MQvWg2kwWUEBfvE3c3HEh6yM9oBAqiV6DxH8+k+u1UUzpe23s3UXFr5ORATNRBVoAKnbP3PHxQ/C
jcxOxCGXPRpdriQCyab5HlevdumMG7zQBZ1/3H8FPwZnk+HX15kJnElW3MpIazFmaVb1PCSW4KuN
s3+Y2M76AXN4r6XiNVdMvNRSGTNPsmPdMINzK42JdycqIEwKnOBZzIVx5IEzatWZiTTogg+wLdwD
A36Ox+Wm0TxOCMQSMBhhbWvID342tORujMg4ahVB7dymqLtUAhYYVK5sBoYkO6kNkWpaBgt2QHV+
8SiauHf0pXqValEzgpoMqv68S+TEKsqrsfhL6roYPiF4jAA5jE0DqPoVYQutBbU9NKBRlsGSBu3K
kAuRmIr+F1AC3qIB1o6HNR/reoQ2E9lvtLSmhd36tuO28NSbWm0ZGMiKS1hRKZd/lajQQlK4BO4R
8OXhrcug5W6f2QM3AkqJ+/kFC0bmv098XKCvrErAiBHyrFMQ1PLRMwMUeXynNh6UjrXRsVPbcj9+
MkHdzChsKgkAOERfUIpY4boPAOM67HTKVCqaGE48DreWS8wTHO2szvhUwyu2qgMB9RrCUcEKKemm
S9Y7CxHLtOk6g5eFlxAP0JayWpS8d352dMw6BTHop5vnn8/Be3VA86DN/8FJPUB2OPkZrrUmKOgL
JUbgXPon7VPpmubvLJo8ZvhiDyvRrqaBKnQCB+lMUsn4hgS4P6CV/R2pc43N9wCOSaHqu5eCEMGP
9NcnYYYuTAc2AyW7RjZ3C3odF+3W4c5Q9E3vgupwe5Pz6NsqCVaOQnNFS9Es2YMGyOTdT+VLeR3C
BOA1r5eZQFq4QBcPddGzLS3EhMdOTzPdQ+H3r7TYybzwnmqI7GLXR7oMKFqN05fgteJgkGICicXx
gFGEXiKLCsJVtX8VhpFslp2HUiGl8Hr9EkAefd00seW5/OOTuTvdXGvXb0Qx5KtPh6RlZb+nuZzS
22qoDgmU2BsPMhjjk/fRRN7+ba50oekNgPWgBZc6FZQ1Bjh4zEEDjYxpA+qlL2XIk78lwxMhrLYP
/B55squr24fKMoyEntem3XBasJRg0A5ih7Jke6X0orN94qqvaDXN3iikH8BOq+tJilBPrjZad3dk
HEd+kWoV56ZSokYJZZtrMZLUpWj5oWhZgGFeiA4pjJu0DsqNp6VZwTu+vDam+sHualRAu/BfF0+7
HBMmQlVIO2lYrw4rJ2/CbQUI514/TP9jBiqH4JoCOaT/cVcG2rLYGmYmcLqnvpK9EgVDjYe+eATd
gaLLB78BIss8LR0XYDbu+TulVVcBXfkolod4dYXdD4EEdztq+yaygmfS0gFb4ZuZiZHkQRinJk/C
8Nj9+USxO2yzQFyI4lA6AbQt78MgbHFv3dosnPOFn4bxsLonZYKXeq/hBqnIULCfTXhMYpL3+Z/A
/LWsrFnloHXeD4EPXk4zbzwA7icp3uCQjLn8mLxStJJLz5S/l3a9f11d3o8yFpBisuwkZzHT3yTK
356N8ync3tJfof4gJYiKOvOZB48Ze0dxm2s9dInHKx5ILcMpUrUB/wQ8uNrP4RXZ/k2iIYRTIj70
TX9cJyqGahIlXd40r07ng6j86IiPzhOzPSG8UuB8T5BMP6F05kdFsVXd3OQhuQx70JpXIdm7HigJ
zRlJw3nEAzV1BgtCxTH0b9Zjf15Dp12xKYZPSy+8EIUqT3aMCP6vRhgU3aWBx3YxBf4/KXifLrjH
YjwE6lZyo4r8mvEO3klR50VCQqwY61KGPf+pAHvibIAm2/IBiw3C7FmL84LTtwY6FmfQbQuMSn0B
qU24HQjSIhVfsXEWaUM4FjJ8pGmzSllSypFTsV7YbeRblw7cBW5hL0qZ6dbsMnpplOHqCBHLL57M
8zO3c4OCWDPJLx3FFxc1SeNJQeO/WVzVeOaE8fsMSHZZjc049rly1qPJcttIJHatDALHvSw/Vf7m
9b1cthvYELByc5dSpo1f2Ry7zKfWDttAYh/GumIzB1HModEV8QpCqDR/YrNbTAN/gbR4nj/btOvS
h2JRwIhuCuWPDgMtluL97fRhjJyir9aCIYXhU24GtebBnD4S3tYnJakdMHKbETxGFkyB0f4EIo8u
pmSpvPYM4nppJfmb2m4rDT1U+gST2LIWJUnERMLW/qoIYXzbjTPslM+ybBTIMnE0nJEzC4m3YaCN
LLU48NbL9uZObmpgFDGmd/+L+fnFfIx93jpg4M/iFpJk0PkRP8Ch4tx6fRb9dJb4meigsRdI6Dhy
RWkDwN8it4R0+ba05r96axQBCTI9eiWJRCKpdtdFSHNIy4JYxFkhbq1HqWtU8TsURxuC3/4nYgGy
DwYbvUoFPu8CQGB3If0ajQFSbIFnkZCvD0ihNucXm8iGkaX/apJoeE5Wnysb3ivM+39XgE6dfqkp
zPMq559GGG2gssWKtH9Sz4lUEHPJw7wnVZDVPruONYPMU9m3JyQnA0AYAUT34P0FE1sJSY/Peo7y
xbACQjOV+3RX/80VooZd0W7mxtI/n6PWqdh3Vj8JRmtjZL1XLNpp+HcQaMpbW5H+ugVymzHzx/WD
9Q/ymRCx5Pa+9W/c4UaGTHG2jeM0ntZBATvw7BPSpJslF/SrfWYIJkgzNkfb53GAl9D841JRg2xM
YlTuK9PE8KQ0l4vEkOoYC3xbsnq3ODvdSgVrP4OOMroFo0Wv2DWQvxVr4yV2Tj7hZZtrlWWY18zZ
Kb1i/Fl60ecF+OdK+dMA9bJM7Xy7WvtCl/Q3cdSyPzZMg97dqmqRiAVEviOMm6fQp/6QdF6Ch2BH
gUkx6OrG7qGsaMQQwFVJ6H2yX9NBTuCBv/766aCTqitVkF9PN7PvaWDOBZrBNC4Wkj9pxx0NqAhB
eadizrE6x1JsL50QSlNG6ySNfb+te4URq9YfK0tuN1VNw5qQidaK6Z5H6aeFnm6ndvoC740BxEh5
QW2fmW86z6YmpHIYVnC+ByvMrkyFcV7kijL2DPywIGyL/UpZUBdwGjcJCLOHcui3Dy+VIin7mjKa
p3wsF6QuwDzZLziO6YY2iYMHYQRJ6hLmFQrbiJtbgZ6otjpSAM4XLHV0RDwKIr3C+WYNQOZgvnXY
veIb0EggIqC4Odjo1eHX2UrBcrV92vqybbLtM3S91Z6Uncqn9bCxLQKsSMfhA9iCM7eA1jACsVgc
l/1axuU33ZmjoAC7v/yP/VWmUbowOAfzTcaPVdU545YRzY8Eh8wlKC6RaStZzHvylTomDc5XyKXt
2sT0IW/5e0H33ShVFPHTzBrCejOauef3MtSNrd1e+kB22AbJjfYU/Oz2i5aCwRYl2SxMNgGzsCev
OkfZpAZdfBFdagrLniPD7hhgE0Dbtz7DRW543iwTayjA1VhdYs7kPDPMZlGqZYti/HyxveY9527u
wbCORhgQElqhuFzUfC2d0z+aM86bU8dMpc/AYXZLU4f1GLzGhlFhaEe1bjS/wI7Z4BVxSg1Mcvcj
BRWIHp1INWBe0UELkcYtsVHFAiC5AhM6tUSt329gW0+1pbwalHN/kWNR8ma29yfgA37cbpIeJ3BJ
xZkRjNQHHz2LbdzydkxiXcZJW560IOefQbhwT9y2SE4c6en1lrDIvdD+zVB4F0XV3ZR4vIS/xqS9
b+0qcZ00uyqbGXKfYzqE/BNONChUdzLaYUgsDqZieeWwMc5z05gz6uc6Xajq/blI+j5bqdTLWH/6
s8g3QmvBwFpsBF0jn8vCRHaVyTh+S8s0X2U1JyA08d09TQ2Z4k+fYdxLc+0C9GKjw1aYEcwk4eX1
r7Qx/V5itAFaRBwa/6U0sfG7j+I0pDrQ2pY/ncMIKLLGs9lNxFHq/GD4Ah4fkcnXnojVc0eVDP+o
KRHpaNrzZa7ystSHqBN5OP1XtA22lt+d3DI21MvSw1/LY/QERHRWRDKFXHHjdfbmNlf6Ka6PRPHd
CyUd4xKeiYpMDAB4X70bdOvJfY1qpnFQl++G48hFmlAdlrMvB10hQ/6tRrDz1wU8Uv1nCQ/DUjUh
y0lvgiuXj4NGBXWFTzhrxpcCnxR1ocepYed3HDdWkAhlrwon7raRNdORo7wSkDU/Pa3eVaqHYuMo
KpvSE1Wb+yDviWtbIhJpg+x0VPvjXv64q1QLi2IBTmB5OY0T2i03qXL1b4+vmhqLbfS4vHpjWtUt
Q8+Uro/i9JnVF/DCNamW3celAL19jcPE0XSskpcGF0Mj3ntuAIh7rVCnQIYfsiednJw+QX434RBI
WAK6nRTY/whfMAb6+zHwvCLBBjU5tn9AI6gP4mmyqJvvxaJyCj8eUOghLXjvgbz1wAnUTG1t3Xkd
1BRQBZp5kMQ3waVQJyfJtLC7c3E9KwwBGFE+844L07TLrfMw54qoIE1+5/Tz7vXidHw+pmeHg7qK
93Wk4dqo20+5R7LeFD7pWd7HQORmP7vceyJ5XlWSycRWOxQExVC78MRdBXf3Mfwk83xZYLekvO9e
5fsO/nj7UPjaJ6fo7EkD2fDTXPvTo6JoEkOWYYq8QiN+R7VYE1NsQ0hfX8t6xatt7VRNYVxx+/Zp
3kJLLXZJ9b0MrH3Tre/I2eeJMBGuJIP+99rwCZ2Nebl65yQsKGintVkgJTZmJmiQKTWIMw1+KtbC
3BjV3QbgVBHBT2MBdAa7W6DsKRfq9JpJbWn8efFs1sW4qol6Qxy+X6SgNKY6bHarwdVLNLycoSQF
i0UULCx4B8gbtEpso+kn7Pu2F4AdDCGfMu2i4TQ1y0Pkfv5MhzxWSNzl+PSOHPi0Np+h8esF+Qqa
01ZOJ+6v5OB43r8oOC4tJDGjG5BC8l9d7n5+kvLEyFTkrJIcsX7IW8d8c2kt4X1gX5d0ClzYxjjn
ohS0NScZY3Rw9a/t5g6RJrBf06KUUC27gDXTHbq0L6axn+FGWUipWMjBQj4xf7aJlDne5At2eTF+
GFh6/okawDhVRk15yC6HqOiD3xdqRyiKBA3QoOWgaRJiDp1wlxZQxDAhJhgGttUJMI5cJNndo6gX
vzFOrvr0jU6ceA0L76TXWVBgCC5SZRdb2um4+RbudAsMu72efgXKmpHrsEgn+gMEgo997dGl1rPo
VhjHZIrbXDb3et4JL8zyPxYRmYT7PLDF4To74wW6nax43x8XNKkMgugXyr6WPOOyNIJ9izCgf0fk
yp3dfCwOmC2a8ZLKHJsNxaoSc6WXnwFTzxRod2OVt4VXm0uKM528A7GPC6FcgqA5+BjrDrgEpZfA
oso6RG8BLOJ+CJd6j90en+w02MXGOtjQ/TjCx6zm0ilh1ryVsVDLkMdpMnByaXVn29kU4BpjTF2n
ip/xthEfNtBGu896lwc4ZSmzCL2i0rQuPWpvByltVfkC4atuB99/Zm6ypvkLnbmMORNpfX03CNIr
iezMeyi27YGbWTDdX16H2FSeqPKbyMD3b7ZSrvLiEZQloJ69zhFgj/4pK6qihKJrJ80i0MbrW3gj
k6oSWsllOiVw+QRCz6ehOZj5k9IrHEkiVnJO6Ovgv+C6M/aZA/A7iRrhjDH9IYHgeUZR9KE55Xrd
niWbzoVHeTyqyDtwNkn9WxsDVtYl7MTzkwU+4NJ7xl2kzfnQtKE+x7H39W6M4zlpPj/B4kI1QIr1
YPsT2wleqxdGhhQlbMwCjUP/zTUk190esVTh/q1FPlHdZ/H2rTKDrP3KEHb8brpKG/DhE4UQyKF6
KkqxcQR3CFNQ/QKd4bkHS0ZYQnImpJf6EopLcJmSQdl48qj1Je6ygyvzqs5hqhnR91NsgFxeDQY5
2g0fKfFiBfgqvb/VyXmZ4PJyI3+MXhcMq0BONb/s5LnMqI96MaeEf5r6ykHrXBMS3aRq6lNGjwCb
b44f1UE9WVLb4pq1ttr96ELfL3rbwZeKJRZ+tVnrFiLEsZCwAyuw9aHesqoJ+JUbyYUvNrX9dezg
ZpvXDnUEm8ezidweO9IybLFQtIQRdKwMnQB7XDiihLoPwDMEbYZDqc5MwNm3MmUVTS7EF96BRfk4
XmRHQwyie0UyOldTPe0OWrm7KFkNs1jvrDFD5ZDLsv4/1xmbtSYhn7cHf5d3eRPoJI4RMXbJQJe8
FuJJTHGzqX4kXAMQfd6zBLCiYX+8ZiPFP4ugrtixjKkouVjQHcU7RXRydjub3ZLQsr4m66XHC9Z7
NRR68ofZiQdUqQYNlCt5WGu3PRfkKDwYA/Hy1Wnke5KMmQ4Su/tRGyCUpk3Cnkg5ANwLZ97YIHnn
VFWrh4a7iIEow13/iCxcypcDI8l9ARwfhqiRv3JyfkaxZ6QKGFAuSIDWLShHRgGXAxfpC62fc1Bx
ZUAp0VoSFcF1OBIE4pYIGSQoYhQKxOnrOykYLPWJth2kjBEZ+7JeoyX1ZmRkbLnKbCGFJVgvv9tq
KFxzDIU1FGaG1+e7F3fdbsKI4DGzst3hrC4mcMtG6cHMZKeKPjzBila/t7ieaGnzu/fU3LuV5l9q
KJUMKkkcPM4yv/GsYZVQfiHCc+4QGtq4iU9aKIfLs+ylwbladodVVuKgNXnDYzxOr1aasuw37Xge
/vzw+YbET468295CnHkModCfdlmadBfkXVRQrX+/ebVFccsmqasntlpUxc9r8mJUEOxyeKDn8Q8i
0LYXZai626zcXw+bxMwgzNCWPLy+3ColGuovkAfN2a2YufbJTSYIJa64G0C7aYwmO1XdfKbV31aP
tvp2oDyx90kqFqdGITs7lSsl1FCW+gQcc/YU/f+vHk2g/R4+nZC+wbTSG0GBla5yCZmUf+xfuKAe
FJJeVBb3+TQ7YZorw5krEoZLHPgi7BF3xv7wX63yXE9d8gMjucQcCybuu8QvgIjhFLz4oF32NsRv
lS9U2+4oNHZSxfOwxCcu704nub3N/ArE+nWoDM2gZPCJHxiDVpKrHuMq2tmkazNBDHEQxb0kfm9x
ebK+mQp/Ce7wZcPuHFTdG561pkmvIaMrgaZWCtD4mEWQRVV6dis4VPlEOlXFd2ts8gxJuOArMkGO
9Q8fYzq3xsg8FYKIVQo/YIXt84lIbhZGw2N71Hs/4fgeo7YJn0VRHOtv6Slv85/M9iencMfDc3Jj
i5qnqXXXoeotIJ/RxoHBBqh1AQp/oMxdVi2ZGVII4+E46V31WSRiD4fqCwfLYTK2RTYgjLbh+SIf
sPcYdzzBfkB4GZLIVK4v5mW8YDsc78ow+hDnhwcAzbnLAamnhbU6H7BGfRITcCWjAWbDloiCFWGJ
LgHGVKFEoM1ZQzs9PZgiuGAe0I+jIKdFzX7kpZTa5/fOANB0VNRbbZojAyxQx2eWc7Z7z/t7i2I+
2lwl5tdkP5NZXvxdsQmsHqPtNPOPf6jn916xDoiaWIn8nK19QZHBwC2ljBbuGbrBRYm9dKo3h8un
KueMIhHkvXBMWQA3pShTmnsmfXkfw23x8bps2FoEB5RP764wrSh8mxCUsN+TAyg4csYaMh1xKE57
DNHXRY66JAUxu2Uof9A2e7bZU+Xyt6HXd/G573KQoNQYV31v1+xP0mVQhcriM++g4p2dycBtxi+q
h45mvG98Z/Q0GvCNLX2IRcY0zuFbEhsXXUYdXa2nJ3vzaP6ZjIRppq7eUb60FNjVYFRi3/w5XWHZ
D9JY+9bIj+poI3tBS1do2+eZaui12sN+3KLzPz0iyMVj6nueGGxscCyjFZfkEglkxoChwM2Leukj
zF3g5uHA2XWV455B1X6HlJHIuXd58JnItNzpLZJexJDzkuZqRg30JkaergHodunA0oXg7aGDDux7
NJEYSIYNN54rHyLNsbDiNvkdOcmjQV0XgIaZA/NegaUw/J42IsfWCtVdAwa0RCnDI3EoG4Zi8f9O
4WTJwD0gueTjShT9vWKdsXqP0Fz6KuYVxxjboP9pMPcqEtzRhFs+r3fMxFORSexTLgHa5CDm277f
UJiM1fNJtoTPnsQizhfRME8KGii2uetbKLilSnTRFLaK9H3S+eMS+5oJD7dQOQ0/WYB3u2eD+qaq
Sg+gA58UK5wy2gGQIebuvyB2DxFMpnqDev9cLHmLJOobGGmCwp9O1CYYRnxTUhtk42V+ghKMLsNr
4Sd3OJXtYEzqmAXF6uusfEHUXqrsU9+DCadodIbwQg2bHBVyVM3VHY4ZxLA46N3gVkd2aoZp9EEz
iKfxANKt2u/ZY5aniQwdGQ5TFZooWXJ+V5abC9CJHG9w2J2YfYcJjU4qhigzWzQB03x53iGUHCwh
VdF0PP4OqmbqLrP+nhqJPnklLVaDRHjBftih7h2iGWweClyJZxOlT1rUu2YVy2O6g4hquwl6vBc8
+IG+gLyoCl4YDFpkVhpKDiG22mn8ks4ccHblhTY3JA+o3qewHYcButvoPIzrRVaBbabsj+4wMKHu
ReNQIX1FMCTRmjPzlcUEcpvOuFGquG88WTlBK02UYu54xU+4CsIdw80wErY9AOU2cKS5b8e/Jrv3
5vQ6R6GObhBuqEMpb2rdYQEKwfUNqNTFVOjvuH3SYSlO8pDSB21t5RYrFHPFu5Fp3xSDi65DfJCV
5FlP4XdPbiI9bF6z51+0V7ToEGQpmJaZcL6l/PwiJTwGaztxxTY9HNybf4R7YHnybG3J2u1hN1pJ
ahNynIs5BBkYAmxFwkbApNToCfQQQps+C3ZoqRKFX5xF5g58z2vfvwmiLhh+ugfaH0qye0JEnQ+a
F/0gNtCEpahAk8rEWORPs237fnvtewC+5Pe8bZpjWVtob9ZyThjp/jIiyiVmgjkvS2IZsU4D6nee
AxRh5QCWeDT0y0lj3ASk8/MwhROnRag/ZMi/moukr1TSWgiJaZxjrJhyydgLPy4TQ2cBPYJb78OB
PVZpSKLaLh9myJzGXLzx6C50sSyUfnVTCQEPqtQ+TZZEdHjve1XIzoASGWUnAoEft8K7FbjBc1ZI
CPTJhT1/R3cunA9YVKxRhXnfb1DCCIaUbUPmhIPfX4klvUtZZJ6s90Z5CxfCf1HT2I6LV2viO8+E
DWeWDhlVXFHbIj1oEWx7mvaLMOFt9jk19x18/HMCuBORw+5BzuPEYwpOjpbv2kJWkNQnJGOgfctF
zh1SMoJeHgkZSZqdG9IIjOv29YetX5G3bge75sQKZvUPowUdISSGK+3VHRhD0rTY5Axmeo7wo5re
KbnsmjY1W3DVLYKWzA3XTN2lDgpbmwSUQCiDFtBE12OVQAuFWkyRmB1GVWjy0OLxyP5It1Gly8uN
BDr2q6QoQ/RzmOio3j3WyKONmDaJLWhQbJ3u39XgP1R6rhNHqbQaavBO8zPD2He2UqYG/qcimmhv
gmsBUB4IuDR0crmwnlq+hi2NQpcqT+7Em2PeJqLksidOq3o/LW/YfA2ydYf/MLShqjK0Ncf0zRAs
Crlb2wwET9aPDlwYbwoqegx066KbTCLCEFnolf0iwORINGQnvUzDACNchTCLmERX6wkBA4eJV/12
gp75W3rLFoa96s/iXXcIGR5ft89nd1qaQJkOopdRayO30dv7gANa8yUAwzqpuEiyhAgmAxYP2Hlx
iBcocniawyUu5kYK5QKDpdQMg780jQs8rY+SfQJ6prLDQ6oec43pLYKqF6Wpkel/Op602Ojzu6OO
dyebag7WyqNw34X1KQvDHy5Ov0kv1hQpIxUC+gx9j0vkj8oohVx3nWNZKBtZxNuVHz2zwXtQMeB6
90RUiba9MaxbT+mqinBV8YvYcwZixTp3gnW6CUzRNjjhNDR2JMFJpuUhJg3kWiMrHY70+XFRq7ru
ancqV+onij0WhlzR9cdi6OgfOTaX7exmNGflJmp3hkAjvFUyLu1omA4uQE2+Vuv4ulqstCR9WyPF
u/GrA/2BpEXwGKlHUMqeNFO8D+TrzHvIIvSTHPPlBOOZEwVEl3JPAHZe/wXWieMDfQ5hB/y17zE0
CZpBiFZQVY9P7QEvffeukqiah4U/RJ9CJKtK9dLLfhOMoFwNtaFDE3OxFIdYrVR+GVNiyFz/YxTr
DTymCf+S3GRDW+oTV+wflLW2Rii7OGzC+FqLmjiFHwnKV1O1ks17btSu+npkXgKBH39TnaR66g+w
Kgbfs3g70WE+NVlqO3t69AiJyaG9sQxYR6odByW1gnSOtNLAlbs024KdXV+fK6Lmus90bHBzysGI
1utNmwScZVDhe9t0XM/uYaGuDdb3gNhH5JHYX1pC/mlenGBsMLUkefdIeZqX5+g14U6PWI0wNkVm
nwel9I1h9DZ/htlBS8o8gJdSWLOPkd3CCQTNL/uZvGTvGHb0N4zdjL+LnF2WO07X9hdGD/O1hGCB
ovtWMCbsdNnuMSQQPRNxBW0l5DCznkwzKx4F7gHW1UHsk+XoTn8v1O91lHFOzIcESnNUMbL0CTPN
G3m26jKsm4lTC6vMPdkfRs40ry2BsbLrvby5XO8VpziDViqeQTPpFI1d8+ehZbIaxRky7xayv+J6
AzMktrZPHLYBinb0Mnhy899lC2rYi9X/4JWUkA3DEOFv8qG/IQ94/XwHo5wkG1cNtbzRmerHo7YC
QrblkT/n+MEhTKOEZaBI6G7N9p/JRbJnD2yoTJ4WiKmodeKvIn2LouKl6whHKrkMyEelN7wvqmsV
qrq7RquDaJPt02oEcQq3of+LRN2FjgzAUQKwORFI3vBBcx7YyEeESsl6WnJw41UaU18gQ2MeLITR
3WgDpNYn1uVbGj5Sata24h1dZ7VlkJ8FDCrB0YzzNQC4AOOyPOJbApHYv7X2etpyh0zKUV6lwnsC
0zfZh7BS99CzpIcCZkDP5/t/BCxTapKFTWOWkwW2XqiwI3YSZvRIU+ViccvQHUppPpGeHWtSMVON
MZQH42iGHaRY4vjZnBzLDuyBIeVwZdeMiwegB6K77Ly6JnxBdwHVE2NYjyhAKXufWGqdZcd4O/ZG
C9s6O/Urp1nkS0I79BHHKt3JTCtuue2bNelB41p3XLWQa9AgcZgr/7HloyEuu8ca44O5VBibdLKK
ANjADDwrQ1s8VniWuDnnRctWB/rYRLsYWHT6sUvZtMlDtdLLLPKYeQqtIX639Ojl0B3XTE5vxgI5
W8ccI7+uRNloV32M2WuJu9wGaCmBw63vm3gc6xRhyiDfPYbFg5+vuxiBnX7+o2HWMhDoZ70yFYTd
ixv/GVTSZwmX36z+8OajQR3nt6rAm/Cnwbh6b72MAscL4xWWtu2g4iLlnkD6CjO3lg7Kgr2vtyS5
N3CV9RbbIRS+39VW7ifyFjtiI6hN1y7G+4HZCxVQYv4ooDZ+EPTpmmmf/jlQHVKF2Vs7bb+wwwaZ
PpmajBfqzVd8HW712NvRO5z/211qClVCxH0pm5GtMG80ACsQSgX+bfrf+cu2iHvWTkKb+ejo6qe9
Mhe2CvA6PyqbxhZflhGneptL837W5IX0BfiH/3vYbKI+t/4Dla1rTmPaa1EzK/bn+6rxqlMwypGZ
NxhoKRHDEnEm1g9MLHXZE+2I6lanv5IZHxpdPdPVyNeUQzHHgapGJ5eAxAzfICCG2KJyMmMfDaJ3
+vtMlceQjvgmFJZCDU847wxVP1/CQncqXMe1MPcPYVAWPKtoGKOGlR/p6dVAB2+txjemH6HsB0Zv
UTsiFKCOsUzejVdVZ13Z4cSTOICyckeyaV+xLFPHbfcJFrgmSqwz2nRHYg5FPfCURxqw5vxTtH9t
R+4LDyxhxl8Z1K/PNXwxkzjhpTyAOFHC/9FxHYYUkJvjZBVlStdqb1UHsMlv4Y4sLkhlbGGfCYxQ
E15F1V+zElKCbGHfb4Hf6i6xe76YxcFP9osvHiJwFNT1G0T7/SfOPMouw8n0WHNHTHBiYbmLsM84
wnMPuOsUTKfRvT5fM7uPrq0XS9cDB1+9/8FojsShQBMu4FqLljFAOK1VxKGzBu3Hqx/ARPPk4Rd8
Ml0flk83F+U+8wR6ScrDtLRceffxLAQMqSkHSoFxQfABb7A4Facihkvd23Wpj20h9cYtIUiHEvxo
MVn0qsgVhGhr+w/AeLdOMryQyQ3r8+jF/rqy5NhzBBFGVJl/3PvDLicQklpcQHZVrCB2K9yoDNd7
HZVEFrrZtQ6gOPjKJCP3hQ2pDzyG2XBEuAysiUsYTmxJrOmKXG7GN3uo9dl8jtUtvxyct74O0sjy
TZPL1sQ6Fz6wUEe9f0vQezE0eQACqfmjCxBh90OIE1HzJ0M31ZXnyaRMR3aukSCDKyro91OmuBpv
VjXJlVaA3sa/Lrh5q9bSefInW/wID+8sHHnIudYcT9HTw00W5TtCW0VJb4i+QyjkK1KtnzOglz1a
EJKPslaPZNoKMcz6KAtzE2z06TvL4/pJZBdKBPCzdRH+X4sMlk6hLI0aZd5qZJBjeocjquhhnhvU
WsMCxilK4iwf7uZFH4RHSqX7WzkiXLKBXBqDLRyUe8hCeUtyaf3SrflaytmMvTsp/ou68F3X+gzb
ZtEL6DjtqWAeTSMATB/grZBTAjKW1DWC5XhDwM+j+l7NNBDX3o/QCEAADcQgdQi8MzBd5H3luvcz
vHocWkvvXCmiTChGyU5En8gqHgM//dwLyV08wAm/drTNRl7iLCZNfiaD8jYzXYSUKVkgmzc8DSAq
hKLV6rslOAvCjEABUZZKA7OMruSIyDK+uM6KxuzoVa27vCmQJvT6K9hML0jrfYC4xHbdvA64EojW
8mTLq3tVk0BaemBOvKF7qFcnSHDOuGBGn1puTdm7O6Rkrp2e/9bblo9rgmGnD3c2NgQT8En4aRu4
Qtg2xWZD9OYYvkKq+MIdIum+9/9pBaojP9S8Ku96iBvInPU1MqS+eja/sP7iWvntY7NgKovnGyw+
07VJ2WgEZKUkTdQ9T9UZ2j+xocyNYXOoYQbbYJrRNm3iknyqxRyuaB1yR+pUKnimTSnf++mEdp4J
+qpWtq5tKsaNjugmCwpJyHO5TBnDariU72huU140rV9f11BE/f1cCG7HHdA93vkhbpy1fLhWqJRK
1dNXVz7HCCvBcgby4IIroFK5lhvaNrami1QSkmHPFyVUmPJRlImMu4IYRNAGVBkRvL+XqxWPWzKW
Bz7fpVFWwgsDrT+IhBY5QvMmOlVuqfWgBXYKjTFboDEywCeVcoCF8l3QnS3Mk6nRYSVxqaZdra4S
JNunheKUOegQSiTdq6EwNU26AkKqZa2laLMkxXhgqaquuUXUuaZ3dPUbnj+kirMt4V5lTaeqtWq2
5ZNDVHFj6KToZ01zDRYtUxt6rcNwWHlU6PzNr2Q2Lutyu04COZ29irF7MlQyMXZvlmJqZnvTdkzb
M9OhjKAAp4DrMaOFxHn/SD5pK0jB1M+DHMXjjzpjpUkb7X84YOwxHRFCo+tmYaLW3mjuBj+xMY8J
iysDgX9amnr8pt70JwnRxcTVfqgp7Tqmkof1IOSEsC3jmOv/1ydLXy+4JcisuR0J6BkazwuVywf4
zLLbOjkS6rHys0W6dYm4hXUXlSX5QQp8I0VXEJByep+0ZyRlY3PFby9yK31LRIfHryO5pgpnCLzi
47dEytV1XRZzt8X2QSt+jrtQs3QZN64SSzGdRaZsHnwPjo8OvcrSkm6Pi0E6rBVRAat0Qw0xv36t
Djp8duredgCh4x9ctV72Ocb1Y4v1KVUXf6qJgoihLQO5bH5H/66SFdI0YdEsERPl9SNNW0nBbQrf
etx2KnK1t5ulpZ/hWM5+Ce/n/OXeCg5BfbRX3ImeozZsBQuG7dbxlsXbFWeOBsnkMRirakWZGs86
Zf9r7L5z2qMqP124tjipeoBJ63Ky0CSVrAcBLIwjuxpocgBJAee4DJIHvAvdpcATSH5F6sDoaY9r
+mZqa5OZk+vbmIsJsCMwPKvcDcfL/3p5wfatCS48/JIRK3IY6jLO35tANbFgIClHICPpaNz9OJBn
bNB0Yoi5N9TcZmxMPCkvFNRMiVt7++fqOZiAav4wneFUvNSlfqtnLV0UkOI2KgiYgM09F5jrtLNh
a6jwsyzpptasw+MO+Lm0+LcBzQUDN8B7u0pS1DsLF94O2+5jCNJBAQvE2khYMIorPNsy+NMDlmE7
BjTRrcOA0SqG/HyXYyeQG1f+qRrfrGSK+GiCT60+u46ucvos1d36u96Uo3hOHweFwtEYHbOu67/A
HhhtbN83RyPhiVSamSnlrKV1iBl9TaQvKnj/aBuCaO9rg99K1vRwCLm04AZgtJKtIaaWBjatjvTz
LiNNDPDRAtBD3EDtylYoslu053V9YE75GYDJPFranJdab8vzBRBH8ONa9WObovIBR3QfCzXeTmNn
0dmkHYZAKUmYklAhJOfC3wWRKi8yNLoXrTMuHxhGHkO0yxCNH1TRjs3Tl63HCgNffoeQPQijyGQU
pahIPdxWLCfb2yQ6FGoYz3pIgEBJFs5QUaSs6FqdWmPIzh04vDkjX24Uru4gG8eBN7KWJVLG1guE
Ner6AYbguk2/Dt0SgBTCOejXF8rXq6KdCDxqNrEqYW0UiUwvc/YXUW+Aiw6w4kEjp5DJtO1+Q0tW
aZJB+DwWDvmUL57w7dFi/P87OyJ/G1e8SxLQxhaSo4+6AXEprDUq5Qiw+fq2BWlKT3d/G3tJEXKk
WMJs7/CnruyjnIWQMDEmBulnq2SCxQ4a54uCYNsi6fozvuahbNExTWqBphsPS6PiyaOHZljRILVu
6VS1Ff1qmApZUSaZnQrkYhpqi1tul0UuwPST+0Dv1CIjKBl/jiGdasSSFPefrP41r+gwazKRVyOM
8BhYw2/2DeADnYxQJvhPxlgPqZjSXOMeNn2374YzpNTO1LA9A62YGCTlPDLQo0AaCy4TjCb/cggd
Fz4SuScOHwamtv7swdL9CyXXUMTwusORCVoQq2ndXYMlt2QxWMPu2UdG9VK320xt7UWsBv2qnDFv
9LOzSBO7ZgBsLU9er/jd8m5nE4vf5/MDi4B+R0ObEIx8xHtdvFU4Tgtg52VfI1pMPcjlYxJDyYyY
N0nxMhyUeyL6XhNp8F5/4u9wR2kQg/qu5HJevh0u4L1GgBAwb/ZNpQ/E+0UdSWQyeG/VVds78IBX
tAcWNe+0CQ9gfhlh+EPTZnoCb6pVNQ2G9wvWOU1u9FC2hzfFFQ0mqz2jF6URQfZolw7U/MoemQkJ
0ThChUor7/ZHUeNbARGSRCZY039LmcpVHl2K2Q6b3D3U88DhR9pLcfCQtKVMOKR0+uC2L+X/zIOT
p2z6CIzJMQpRan7jDWVa9jz7C+b+o8osr7b81TkrggGR6CSaTObMn/pe1haAFfPKkzxWpHYsKEFm
iTJ9JmM/ugTlhELsUw3QI5Z2XrCG0LdnWtElNF8fRnGhW7eRFaqEv2wFLK/Ty8tPPBlPz8Y97xsX
IcLBaRdWlA5GQydHEywGAy56BZgbdhW1SxaE9kRUgrmaM9H+vd03YSt+h78bjBSk1YrQDs2Xp0DG
o+OJaFU2aArhzF2X9IUtob9eJG5QVw4svX+iG7CB1K5CfYw3jVBp8xiGE9GytEVesDNFroFcP7Jm
8j5MS5O5odgGLYLgdwS+IepTbansLRJGassBscGPJxZDRpC1WD30hpCF0ZHmOA6ICkthWOUGUTiQ
ngugOldZg8INppG5Awg7omQZD4fXAOusa8fc6IqQXRBjUS0NDVlmo3/qpdy0mCMeKsbfPeZ7gFIN
sJIppVJQJy+hnsCV5rkgr74uEUB5EcgKELuRr7t9l2llfsVHnKabwGkaB9j8/e5PvPbrw9LPCoDO
8s03CFQXdghAVpB5TYcdUfQHRErgdg6cB495N7uFDu12z0L1AaSsMAmBWBoGzw/Q8kIRkZLdiiKe
UssgKSLCbBJfx+3K8EQIanu3eJ7mYJJfLSE/7qfUvH96kJ76RVTBnctYiAexOve1eIVd2dk4NNYX
x9FVQOl6A1rLOTW8wPvlrTLBPNtRfKNEQWJotg+RC6k1rASslmGBY3DB5GMip1zhg8xzcf/sGKr7
pL6BO30VTwfEyyjfP/Hmm2gkms29r3fwUqMcSvF1Bgds5mVqC7wdrcPbb7WbmtrB/jaSrtY7QfQg
9YeGyInf4CWBYEc4WF4eB5UTgL5boz8T76QIf8FlPg5r3qcubraZlid4Ig/WEvEQbsUIwK5BTbbO
hCE+J2T4rWEvaDB3Nj69xUhV3a0IZNMH7SB9nIcvWleo2wd0BZ/xKonzlEW8cDtnoH+nYc5Lr+yX
j1H4yQVmmp/3vCJLhqc0Wp89LaaygR9jj6wWJENKUva8JGUeYKaM7HcGY0U6TUUz2kPh8qOonkEm
2KxCz8gGK/DjFkiOku5uvHsKhB1iQi22wTtj347nq2+G9M440Yy5ouFgwVDZR517cGR4qj9fXfJt
0qAudujbRDEHVOlZ2FM1UZ+KPQeE80eFYC6mjbztPSkASyyTwfMy9/XS60JpjDdv7Zzkufz7P2AV
tDi9QlXz/0XSclnXQIcpQTn31Udb9XqoKfYXUDPpaTYV3DAtUkn6d/FmMIXu/ZruRLmnNvcLopKI
QfAAcgsz4ss4XDiS9hxVNHXc4HzgssmO7gvfpZ0t+MRo/o7QWIC2bjfc2p72WW1c+H1ld5mSJCqa
/NTbehhq7/3J418nrZdtvySypxHtKF3uRM74b6U4X8YVoSxLehRkjP1SI1cAq2JW8ed/0d1i7iu6
2VfttQ8XL/NSQfUsrasj0QvkLgjAi4n5qhuGmFZrdovoDx33Ca45L6LZ2DSh6l7c3oBi+c8l4yUj
XJlQw4IBmbnYOV+XUHvyaDN02s2aEsowaPXY2Sd0r1H8g+6/MSgNRVdKyBrOifmZCHwPyqT2udR1
3tLvOjfk83ZPYM0zR/47N4lEuesUDSL75k25a+zbnHAROzJAMz2xYIazoEu3UXqy6v8ZoSL9xpvv
8X33hJVNzwzYZKcpADZoTiUITguJIw6LZGIq6PqMCn9eI7pTZ25vF4BUJicsm9lG9jyrBmebEtTA
xxU6uJZOrwBX6k3QeYXTlQeenmLt9wvyH+94cZt59p4fsP8eanuw2+6+gOOVTo0sKOplhGw57m6c
BGjpzx1rVbFsn1SDAC3BJAyMYqNzClUteASZQvrcwuCtAEIwKvf9qKDHlMmzAHBLdVlPeAOqSWUm
ccgqeSUtYQNxL3J32LeWJ5/Uq0tLv727RtCBvEJcMLYN2+f0AfLvTebqIXOOumVI1YwCXtHVtwpw
Vyq8+u9a2tTbS8Ec60HlXaZof+Kak6qiYR/Pl+MOei+tiTTLmpPLFwmqgd/ZJqB8x4KRowr43Rc2
g3jkJXUPi3u0lGAvha55s6tVwz4JVsV6MnTsl41I3WqBEWi2hHt7wYlWncfT0DsK8MdBpUu1HFE7
+AQIevUf+rhSLKWW0XevDoUijqi9V9vg0m6UPL/LOiyfwa+ITLpJ/TN3P0g3Y/yLPTybp3JW1SuE
i1F5UPo6HeldrBYefHxF0I0cmcl3WqYCePgnKg4YQwIGq2mT9VddbBamkS7dpJtX6qPAwIV30aqp
VeIroRaekBabcBo41/DQSeIp1LlqWtfMj9mEJq/jA8RCsuT/mSnbGAbG3A1P+B4eT/twGK4888ym
vHB73zLEjNJTyONIkRG5e3kbDyRp3THWLn2qyOhXb3ck32HmDK/HQuEMBSeHdftW2C5Id4Mlf1bR
yKIcUbe46uVfXl9vYzfezWq6oFOg4aQUIb31c81inq2fNHLYgmYMGGm6qP+c5nZs7Qlxm3zNBYPc
5+OO1CAO81NIUvTyXQFV0kFSfHKqBsXArPNjHVPuz9Z+OLiZYhgwjkPiW+8q3+Mc2LfmV4A73ZAz
+0wfe+R0pN3tXgDgz74c59JBdf9Hhlxp4ETV6qgTLZqZFst5RcsKcSvXSMT+OEBm+KNSQKn2UKD+
PJRG/QRvYOZ4hoEiaoCesPXN3GZUpOXJBUK8DWVp4sNyWhMpPhvNJvxeN1K2K/iv+kUG0sOi9LDt
8MKuHtTp62NJYteu7fLD3fU46bkw1l5/rhxXD19Ntpiuwx4iyppoQJyu6gYx1O+lnCdOJfsVCmhS
SvVt7FobZJRK16GX+jGrxsVk0oQuGTUPQTGYP1ZUyRJMzmN2EDfewaHF+Wu0Lvd2Gz4zWoW4wQ5i
DPpJB0gBvOgnqUUrXaz5paBhgp6z/24xKG0QX9lVmOQ8hKH44haKBleio0XviePJDQHbYb4GaSkf
ZQXXY7X/CJlTYeenc0lkIvwaQ7BpGoQJMyOncAhiXy5mViOQT4n/PhxJqSrbaHvCEEIoXr5cmdvo
gP+IeVW3UBRM+ICFJoBxqcdDWjZ8/ephaHwtMDG2oGSDaN1ehcnSu3/XLK/2LTlNobRC2nHBo1nF
xihUEWqoWCCWg6ivEUGB6bIGZGaaAiGp2t/fVA+PI7lRslMT/dNfE/Wtcq+7zBgPNQ6c4VyJRhpF
8BiSnnr3hjchWVKSUii/yUj38KNOwQ7xfiIhESNI+PbSLLprHBGk8nOe6tSL7baSQvCDBj0BYmBq
bScgUCaNlzm0I2xw6OA4cjLti+6QCah1JVrivVboN5D8wMOeIwb27zkpF29xQGshOmwV0DC/8etj
QUZrM8Auy8iamCSKqhLCXY2n36pvzeHbQBIQU7U5QHgQhznU22qUaLET9W+gaA3l6qSVDpgHRlpV
t36a91K71PPqsZZMY4icrcVN9OkpRwvkzISECDVhEIaetJ7idLC9LfDjSptrOQnCjBviQk2uf45h
tYpq9uYD5+A9QLSOXQF34UypnHZSfZIO/RKyOoBgFgLNbVeGHQQTI64djeIfhCHrzN29RiyGq6/h
mqQW8R8koJMnlbBf47wqQHkHgpVM7+kcPCJKpgMFZDWcGUdgC1e+hqBpzhUnaOQILIoPiqr5EmWM
8RvsezFGNpNi7Zu/d7VZlPxo/4PJLEGeC1upcvTmkwqLF+/jKdD2SoB/i0XG313Owqq+uV5gVfSC
su1y9fVJpMdbTdx5TG4AgMXOy0DytEPC4an2mP1BBR3Wa8OH1sH9FMejvxUvJReWfCGVWJxUITa+
KS+/+33E7icyd8kHESlVuNK2Hh4ClMaqNWIilIbFR02dDVYDr0/aeKGOzznNKcGz5HDrixvYI6TM
lB9J0C2UWbMdmEtW1eT7lSsbbG0f6k4gHidobIwhfbMQ6lRA2MT/TngOzp+3T1G/j5zvwNWzckOm
SAPHd39/YO75OuOEMH+QVs3AsdEI6H1fNf1oYvbDF0aNW2fCuR6JZMIEEeiMbAwD5p1zZ0EXweNU
gW+xeR+h7CBN+Z5JaroIEYf/vlu35BJ5IBy4HDhBkwY4MlIGcpxGSmgoR8s+Vyvy/goUB5IY3ZH2
9pHTPgkGMiP92+obyurMYeo8S8Excb4xjrftW+ZUhSElpzLzJj7a2SfC8vxjb4HVU+MzOxM9s6hn
Z02lkHry3DKPGPBrxDKA7atjvGl1GuXIleg/W55IaQYotZVFKRkX4jGLEXM7HVncXFo2xtkPdXIs
uN/34K34cpk94tQHBYTiPjgougcwInut9LIcAq+U1zNHaZf5/kKUgbVvZUSIqb3wSzdTXdfrkR3d
yurmTFmwVSKL3mWVpJS5yG+qPneZfbv9jqVGsvbRkHOpkJ5a285ouNQU3GcSWVVYdLkRqhUNi5eS
bplrk5Y9nQVcmzsQ08BxHiCX/AvHGtZOrPeQlvdIOY3rKkgomgWJsfagfZGwgVyLNrS77T3APUXs
HWwgYTi7FskzWnAnQ7KeDvwPMB7tUUCEKJuoVkX+x5lFvb9xL529d+3AM2GfQSE1t193YeZQx7Wm
gKc1NXYt9j0JBTvB5lXSuSUo+fAsQKXeeZyK7eaVnr3dmjTJsHE5EA8GsC5FWJg0reAxwfWQXLCt
cxNmH7PA/l89NhHnxYWPueEoZE83YQRJEc/eCd2QlKXUfUW2Aou2zaIfd0cDUJWSEv1tlP9caxo+
Ag+j2xYn4UhQCuv42p+HTGgZpVZ7d2cNXGKYnIaoKfEywLsl4rkiduHIUtZHAe8QuS8aYQza9c6H
FdAF3X9yLDIsF/X9AFTzhLULy8ffrgNphSkpdI/pR0LE6Zuq3C7DuMPJO+AKnV01qacXJu3CF1M+
jRz9kXOlTSiO+5MRAtshbcBu2seBzhQGDaHANVg5DvyFCmBhaMCSA/D1Ky6MxMS9z3b6wevy6bbp
4n1eEIRhA9oA9CCxbASufdMTor7P4o9y6N9eaMxAtck4O4BwNyFsTbNMN6oitkU5gXh3YIk5RLFp
czsRvtNj7S6Gr5rpBp/RhkF/spEDABgzozOVyyJpT+riEA7llqqd3SnjrZ1raSFClpShWvcmsBKV
9cxdaMJdFGpP8jHBDOsLRWVyPdOxW61bb+Rk5Z7qx+hcxLUo3EBj0X+0Sk/BbeDwYcyoGpn6ZHcx
1RDztIYtebenKzJi8l703fyoxuUImMyi07/N2agFEj5VPBKArOQsJcmezOPdtHJLZSIb7iEKFVUw
1sfYEacwfExsyinE1+sc5vC1in2igWziXzFa+m7ftDuiN4WxJJEo2flnx74R8KH77E8IZagjypL2
NO0c/tCl4CYLuuIWgvKrESYwqu3fXDRCSPtEbpT45vGO37tKDy2NaPmgkp/Cw5+wLq4bpTCyLIpk
JzaRakBapC0jtzhs1eYg6oWNTEOVnAvq1m0fPipOkp5iYlhCqv3vszaYUK3EbZIvaSw94iMOKE4N
lEiGThKRHkcbwnHafFXy/aLHc8dt68cXSqTw/v4Hj0puIH/HDsOD+0WlLcrcBVmo/I5DaQpHbODK
ElVvhEy09Bl0Hql2/P3EVJxQp7llYi4z2TQgwV5YWNgm2VheMdWgCeiylOpqtow/7g6rLtFyBTtF
iuUGvB9ur7J76MMgztUpdRKSgGjtH8QWq+Bo2kZGVNleG8dNvm7lOsF2F85hfhKTC6Xmp8lviYGE
+KvVF2UJYCzQJ68J+JwdqWotTfPJ9QvRX+w0Ia+GHQE6AhraXS4CvN8MBesrM4iA+jSrmLDbsyFd
TSzNuxLOe6R6isV2KkQgWMcUpSskJcYDOuAk+yk+aPr64E8jEA9D6wvdXDGRTXzQZGwtavvQfcQ1
HTOC1L3TwM6p99Vs+rKRr6FyYSn3juXDIlnfk5cfAbvBYPNJPUHHQaWEzy6LMNU76pxFBqJsHFXF
DUC19ziU5/d9DTmrkoUE3J7EUjgXlnyI10axaQEN7a/VqCuItUrzNhq0vZcOLShZ9ydpy+k6s3J7
yZLg4qi4A9ukc/ECfs486n4PsqeQKvP/iHU2e8xtz/gXN1Rz/teJD4ESI7z3RUWNWmEun+yldgH9
+t423TSL5+XlPzpYa4yayn8IWjapjFod4l6q4V8dIOMvlKa8YV0ymb9Nngm2L3Q4wfyH2jA56uus
SSMGLwxMLKNoYTKoEazGbA699Y19sATE0G611paW6f8ahgXdkQzXtfKkQjkIARFFDqcrrFRnMbFk
xfKuSpGBxdqvpBzLopTXh1m03LGxb+beYwmLGOIjfPQCDPCWKVYBlhUGaj+VjRucRepB8zlT8vD9
JhbIy/ITYaFY8M9+XSVvOq/HJoIaWTE4rKBv8OmHyBi11OX9xrreyweeNQ9VJy1VSuyVfu0V3IEa
ZYZp8O2BTCLL2cIT3VXNSJWmr5InzJhbboJGHZ+CwjUyU1U+wYIl5uemIzi7QpKqLKLno0A0kcTg
2GEBbBWobu8b9sdxK//ZUhtMODWCtb1DrfiU4/DsOVyfjwKLymrRtuQHrsHwGn3MVB18/NwFp419
PNMW+mMQqTv4XSwRl76vK2PlOEKxo6HRvop8aCcGiU2+0SRabx6saaKt4JBkNV9JhqoKMElGhP6A
m/DwAvUz4gH5aknr3F5qRxh0gc90iiQnMS+HEI8YPXGq4unIGKRO1ajrBOeVpjUYc3Fbav5iERAO
hnAXTGoF3kbwlOwSZXZw4unNEhi7Pg7h7eEq7+mzWNLYXbggjJ7QTnMKmy+nbLjISl+3hLIVq/Vy
fxddv7VatLxLPZTmNIIrQxWlZ4jpVQy0Smnqm1llP5JRP3ghBrkh+7qNb6JfiPDigSDbkiUUC2wU
C1D3cDSw/zXE6+59PT4Rw7qGIPODjSHqKTqZ/TSdiNvC8Abuu6+eQ0sNcEQ71Pf9GwlVPlFue1Xx
FuiqwBSCwYMsul7nhPn3RsKa6Xps4inpyHobD9ecUHPDJSgdv7MVef7tWr30n0q8pJygR/8om/br
ko7vKmHuOOsdvphoRtzOrx09dOg+YJaeFDlLQ+Q5RMOMQXmBDF8/iolNc0vdxQUkCGCRDoPHPZTF
4buVKPIoxQAImvxfIcw8N5opXW5nZk7Alx5qmL/triFrqUyT4EBN3Sacbm64IuEhuILHFvNRnPJX
khwp0JOdJolA/P7QYAjwb0GzNiAmdtftbP26QPfvJV40nlW+oxGmcyXw9/tVS1WMzzjEmMT6CMZv
x7UUfvUhBKrbUzcUOOtFg0KCjJz/7jaytOQhPCZA9nLEfwIqmuOOP7gguYsWdpp6YroD/nKp+J2i
U2+mSJzI70OfBkaQ0R3djW1M1/AUHrq7Hu7iUUqaVfJJhoiTHoBEb7p778wpxIP/6X0EyVsY7vZO
+n4+fpasppqBWVfDhc5knjzSeWXSxo4wKdc7MyhZHTsW+ZExE7mm1o4GE3JwKoAElgwSusRmccQN
F/xuo3jMLBkR4mQd7xHs9P5X/95rE3OjMXJGocIOEJKGdmYK5N1JZALFHsKo4bWqht1adFqFYnQL
4xyyqUv+wAhL8gfC32bKakhlo3h6bUkCSDXTSulfL6Nne/Lqn09BDp/cZiX2/1mQuOFxkL0wZx15
phT+WvIYslaCScWbVGtVDz5QHoVSl3yMB4d80dxZFc+1n7lHSdJEE0Gcnxkf02gaQEfucdqRXiFA
yUHkV6EZ/a7Cl90tDejBfEBxLEswLTF4x862RyhjdgEXeHlcBR7W2FUyLQXf14rs0WQXq7nQ8f1u
XSqryY97xSXwkaj5j+w4K+YyFTyb+mBYYe7GNo5NnG3ZGIkGcCQSYp1kqCrFJroukUaphYJ5KbOj
vf5HpR94t1dIf1LnzMFC6WPePIUw56I+hxOymdy8Ofp1/E4/F2+evRwTMJNQ/MVIaU39BOlHQKYA
PbKcz/pyDvlsa2xtSh8iAlu9+x3Xdpn+swCsbE8THWcKoeWXDki4gfKs5eJs5QRqp2xA3QwnxI5J
7WO8+toqce/4zazgoJcwov102K11sUwy8gC2ZgH/TFeqQnqTQqYTVxp9ByXZvO+mG5qxuiAANyca
IOlFzYjnQhSCcNsKM9nYo1jwoGRdDTVvDlkQfQnHVUL1WzxPd5S2d/BsrS+2e4Fq45wI8p/Jsmfe
hBa5wqTnDvU+YgPJl1i3DvAUgXKE/e9xhOg2L7B4O1ZHxBic//B+B8Q1YRTTPBP9AHQ9Lh8X2pet
Vo4m20dvKrxrDWghnFBujcU3oM2JXkdFDwkxo/o6pFIhbsqMN58T6Ilts4ekU7LGuRJ/lAn7rgNM
OZC8ca0+1SEmiMu+y1DzEMXKD680qN6K1HtjxtcztmSLE9W2vh9juI7K9Beduzn8WbJI0j7loA9+
4ivB38Ys874o6m2P+pGgwUqw2pkxr8sIQCt0wJ/pmrapddJpJ6lqX42vJKznSre/6FcLjEgQnjxl
QkJjhnfC4cSWfQFb1oinPL4o6WCRO5Cc163rZaS0iDZWYQR2/zVvGd3AzbAVc4MITeLmDdfapNr0
cIqScOtc275E0R02OG1qd0fb77wdwa+C7BHOBrKJTJkmtCQEP+E5FLJjlH935jgw9KV87MBEdwYk
Rn/IfpU7EjbaEJaijb1x0v41J3pLelgbdd3y0AaFzPln2ypQ8z+po0bDTDNQxTC52WzL5U0i2Khp
fZQm0rzPeLci9s6yNw/7a8Au7e/ruM6QKp94I7E1qCQ1s2lgwwST75Jaj0OYwyXqwxtUz1hAF2vn
mvPQBEV2mdnhobDM5x9+ftc1HMZsjH9LOmncxTlSgqEEkCwjeNYOh1O0OCWaNPcPvoUPqrg9EbJP
zyhJIxEbV8Wb3sIW4/9IINOR0dndHkIbjPT/Vt9BhxU1l8axJnqxHNNMr+RkgxrAuVax5QglcKSg
mjEaunecuX40Z4EQ+8wkkq0bfJUvQCrIM2bQhenh3jLEVyl9vTkUPihK1/5ZKhbUF45rEHLoOsnF
Kbt4qZYKcZRxileDbZrcHktV54gxrgL3049jOuYC2slLK8DLX8fzlONt1uB7iMEYVXGXz211uLcZ
Xafg+NkJ5so04B5v/8qhllwAixqsiPqm9zvQVZ+2pSS9gR7eGPt8NZ0DdLykaJVKlH6AEmi0SEM+
Eu01S4htMT0EwM3X1Rog082UPhF+M5yTqeqwe3FbcYXpG2cKqndIlUIkqLAfp+CZBttSrujvDUgD
MHakESiuRTvUGmP8PeKkaYmOvtGdkDLaP7jFnn1M54SVspyPhRmJS6wflZBx3EVsucpxW/bqaJ1i
TJ3Jp1NiR/jYQ+jj4Jg9juTRlsRCBGE50mk8WrGUb1gdmBs14ijY7RmiFpW2Uwqbnv9JhLacBwIC
okBZMuOiFVNUrP/WEwLjz4Sd1I74Dx/hHHmz9klaCoYeIGYbFHyDhhGL494YWx/dPBp8bdNJQBWQ
1Hv8/cqwGOz+hdfabx97sGSc64DepvadTzLIJ6zvS5Ls64bWnYPCf6/epFDC4p8LDyCA9XShui3G
9RqZU1Df7w30pk791kc2RDeByKfqEMfO0lqxdVKCjjGuy8oPtUcABihtyIOGFuxwGtGM1AvgdKmq
sPP0HA9ijTNm7LUaj7eq9aE4c69u/tVr8U9piGYJxF33NUmaCGtPHALJ6TMQxam6/ZU/lm8gsh0J
KfNRpRWFZJDdYL4HxY7WJnNssqZk03ZbSAjFwsh6wvBldIsv9fNkaWoSBwP56XO+oi5SDZDSxF3Q
LGH19pPIFLBsSoqgkNv1KHO6/XrArkiS9Tbtf5eq35R7FOTggahhCnpamnXsxM7VNy5k5ZjqwQ99
Vdh3L4AxuPAkXPLvNuQ1SAzOxzFge2+SEnGhheDdo6WjYVqYxOJ8SpXWCKYraFBhDopm3F0q7bKi
2q6pECfMwH8gWkfd+hotOOdHRk+8ivY92GxBlaJVliKOoqLezw5xjQzS1sruQoR/UhxekV5RiWOb
0l3EtTeRjdiFYDchZIBfF2LmDaQqF3V9CAG1JKIhu3V1umds41/5s3Lj0qmBqlZoPapka7sueM8u
0wH++N687hIlrjZC0PeICLr7HEbl7xCZGf5w0597GOuQfpLfaxhTGtL88Q+ZLo6LARm4P1h7K7V8
QfGmbfq/Wc3+zjkIoF9dUbj12w7MdnkkJ5lzNlu8JElOxREJj4sIGIbsU77abSjvvaTFrzU77HtU
tOLoZefHpeBSvKvya5IARqfHx2mVSCu0z+UdOu4R0JQ+YK3LRP/PhbZn2UTluwogCh5KU0glP3Iy
xiRX0EfHB/mAlq+PZkZHhLUL2xJEJftgqbw2VmeLmZK2kQ/lROeV/29jOcKL1pbmTUcsf9xLIxQQ
duTi+MO/3FC9J6K4GwqYA+2dPULoh3dyp7k5fjj/SJZe3+pTBazCeNXJ+8PoJCuzUrolRXWKB0iz
de6knolpLwUiJFnYbY0ROISOg6RPjSKWQJaDBj5U2iY6UodQpMYtri7O6+7b/PAoCVX6hWmbJS+g
UmSHu3dAaUWNM3BO9K7raxsGa4KISLd4zSp0QQoYxO52+BCPI2U+btqXY3S7fIgB4ZmLmtnXhfnK
HDtw0QZ/vDvMrt+yoURir0g4aF1r0l6wPzEe9wUXe7Qe26a2/C5No/ODrxYxv93MdUgXHphyd0YP
Y58l0Ka7fOFDgJGPQrDQQkoWBlD/52p2mSGFHijipT/PBsB4gejaKk4V80/RK1dkVgOXaVE5UwwQ
6C9rA020aV4TATT9ppjKOJNT4d+QEBTzLYf1CXuwPjoSVQ8YThH1XhE8Dr5H47pHAfbUoZ+GltgM
QlOPmbIXR85k8X9PlST6zAMlgnODsj6/B7vDFzatdmySoJ7x9odVuDo2OY4AiPfx+Zu83nd7VSHV
gqkUYgjh83LwnJ3Awe8avkXyZ/HCUyMrnKOmCugpWXtlfgJPHb4+bhrPtMXGcDJpkk/zp/g4Ip7d
M9SD9qsAXz2ncAmiiv8WxDlVbM4FHALqOL6mceSgSQXDQ6rgq2mTurX4IyEgdwW9fp45wqbF6nR1
YhcLM1PzJS7hpuFOhotTQ5pa5IPGJ3FbdlCSPURGGHgV135DKPygC9R3mzM1KCqwAGdH8/1XcQx8
dxlOdffv992/W2gu4DVxy8cgRE4972mB++bLqp59UEdmCZDQiRVTQcBX05WDYt86ObZTs+4xAdsL
th2EDuzBvUSZIoahwWu0oK7G1ubBOT5pCLSxKyPBAEFf6wgpluQFgCpQizA0H8AKXhrfD7oLGM0Q
MXav1T6Q2izDkFwee+GZBzkYisuKcBIyMQ4zIqeWrwOW4vitb11kadUrJCsVrb9rr3WBSgRAA2Pi
/ruZM8xogEulIyhwmFTvNnn/2nM/nx4tvdvRwPsSKWdHjMJpmlyv2k483Igr6tYji7NHq2YvfLHh
I0glkIS+FcR35Jz0Bi9c1H3msBmLLFDRNI/CU0NLxKnZWnwSgqEzM5ZLkXiODQGUUkN0BxBQUWvY
BRyFNfIBOhL58oe+pMbzhRahInL9kxWxMXPhVPqvvnL1PyLeK6Axi/VlDUjI5kmr/onIQkkGCWxV
dDlPOocwudNYJLa222/SJGLQRWP05p3AmC0ShgD7boyhTQ4OEUXB0NolOSxg4AHqCuzvumBqvC58
hx4pr/uq4X43r/fvlcwtxH2bMPl6AJkcFC2HZOMBExHSNwoOLg8f0GfAsvAer5j6nod/zMEQS1Sj
DY+beUTeal1TKLZCW+j+0NtH0743Y1ZIpW6wAiI9xf/2+Vi0T0e4unJbcNXgp7Nu+UbJE2TSdna8
3fEHQuN/RqAejzuEFgRWpni/KhJiPFZrXX7O45c5stlLNllIeUKShxLAOnl8oOY/HFl6NwERtNcN
I+qkpR7IfrEC6q4ZaEym1NqgaRAmdipcNBG4yIHPg9e3un/wWFMpWXjKqLMu1nKpmCWnuA9g/JpO
u1hWnFvbbQrRJTtoNFeLfRy882fWWgeFY5Bn+t0PLgEFHBci0kCbi+WC7m4YuvfJPKFjL9l+MS5u
Jehi38mlYIhz0x81lFN43zrFjLRPdZaaFhtg7ECvvAvrs6+DTi835Cy5EwvWqUamyLmPLu17fz3x
lp6KQiz9MWH9rd3zaRO0uM2Wi327cZ+KU4abLXCFRWB/G/21G0SkirjHIU/d1Rbk9Cm8Z0O52gPz
aHqTds5nkr40tQPx1O494zcfjG1Rgd2G3tsih2na3Cf5ckjiyIf2U8z9UDTD03pLP7Yp+nX9EXDt
zK565hbGexakeXGyQ/SpbM1OkbdU0nZ/emq/D7L8Y5VdrwAnuhyGO2PbJZjn7pQS793iPLpXMgkW
Tczt1nqt57z61llCvCwMl49bUUTzOW0B9xqwmKnkwh28yb+yx7QfMUCthfRzFtnKsKmQpjPaF2u2
35cIWep9lgw1143y3iNIT1sMI9ji7tS+Zq5Lt+xo1JZE84MwjNeSjdRPpZlY7m/nTVzAQ1tnEiZu
TeQM9asOGw4APrLNhHBNg3EBmee/SH84R3SdyTK/TZF+9q2Ry7Lla2RaXO9743Y2dDgEm2Ij7MF2
ml6kRv+V1sPCbiyukFx02ZaWJ8P6V5aiABnaOIzsTppAhNdcaaHoMxFbvCkmcV/fAs/5LuR9tXVK
gpdMG+bbAq19E+o8siJH+rn6p6v5DUMrZG3AR7mVrC/7jq8rWisUImUAkel7WyxBT9AWdBgQxIc/
GlpUG5lm+sPRpxWDG0Ic3YkmuA0kIh06Go23cixKfcxyyjw6KtWl1HTB+nrQ8KVNrj2eVXhZ4T7g
2vQzVCn9xhSkP9BqRLt8+/9NTeVo8DzaCiCDsZZq2v2GP9xC6NpuydHwS4JacChx+9jaDdoXNoPG
qHkA+Jkj2uBl/cJpgKzCFohgivyjouQrH81AOFb1cJS2JxCGqS1HDpS7SOOIJ0WIEJk36YUhIArn
usXu19sm7FieA+dKPUygQAbov+2DRRsAKDPvVZCRHipj7NIQ/ZHFD+M9ACikgZCVxGbxB7EoxAxe
8cUKhtdsRl/5XGpK6tzGd4WShjCEzPHkvcSGMEOIN2ZOJ6oegAXW0/LeBo4oRez3/K6qFrDmOOUw
inVCR9XVbkZ6CW81s+YsdYY96MjFsp+iHkJo72ooxDPSwEhg/wt/It5+1HIegI8J6ENL/P+IUKcW
rSiSozO7yb2rXKbYm4t4Tq3AmYRsPbp2CQE+b3U4iqwHZRbJCwROsXYCvnjmcpvWBXEn/SDeTm9J
gUOWTT1PoaWz39ZUhlb52yTDSOIk64NfVytyFnCigwMXp3Kq+cvYYhssdWyx69aPcGW6zWkeYTxf
gjPUuGUAxYIHvYskNk5zv3SfOQ/aZihAJCOS9VKX8ReelzlD6xnGsR5Pd868PpByjKmdJGgcsNUO
XSAz8cjictvev+1hZGxzSN9BG2b8LDVAvRVK7B5rLGi/Ua9ifhEcCOyLGCFHtD2iaEslYve7k3Ho
wcx7rr//GfJHoreN626W2vpd31TjiW3kyRO4WFdoVWGmQc8svKzFZG1hhy5ThqDxlH2uBAXz03KZ
Fpflk8uW9RFjPhipoSP687s4yzPkYhOmP/3pTQZQvqHXHz/wZGWKX3Y7AgnIKro3D8XQf1bQTxCT
0Xnv1Z7e1g8qN9q9ciI2uF0WLPnPP2s/A6GsVd6kcYTPtVQKktXzZpwwXKpiDCsYf3mIRAltYCeC
OwPgkefDQhShw8Cl30Z6LBtQzRFowq9tCCfh/g82dh7Tumw8RnTZb4AhbDJ7IUB1pJ6MkCdiUd3b
YgIRY8Iv4MS934rMIJZAL+xMqbNU9EB0S/somUaOfMcl5pUyqnF1PiZC9h+tOlxWU60rWQrUSJuu
ZPz5QfBj18wm7s+xUgAhxd4LQuFdDA2ZA/Tyw90z8IP4Gzg7NinO1IQIzsfwOi5rsba6NjEUn4Eb
e900Kpn55mm3YQonS+SPcQi926QqLfm0jyWA5FVNp+YlBVA0OEeMtrqnO5lf4yxEExsYkTo34g+k
FNtwEuLoYJG62O6AYmO9Tv72R95HfEi9CiO/Qo7KrB9OGw36g4+oNGqmghF9/lhhZ8esMPPQsQ/c
wxVVFUI3pjIOcvisRTuN4u4ms4tlvWvpaThMb2Whhs4P5Zqtcw8+1c+MA+hfR7dKPvDweocGJDUy
Z6NJUeP49RKmvDjwBxVQ3Yily7WoxbwOBoB1nwaPauR84aEVC3wzrTfwhQ4d6dD2vOkKPpZt43NU
ALbmS2G4q/kTb664g86Z7yytwHw83XcvkJa+s1vkkPfBYCsZ0oKUK4PAy0F3xpz70xY7qTI879rf
6J5e4O2HZF2mK7Dsj8rvsf4Qzf7nLHr5nRewkmigG06KRfnn3OH+/FwnGKpISVql9m9mthftOusd
bJyVbw+6VDCMZj0WlH2kWQcavZCjcymmevyRiS8vbZ/lkg3jfd/YnHpV4VHkJ76Wqj3NZtnjWt9b
WyqXvY2ha52LYSN7HBqAEdOc38o3Zsu8L+YSMwfYqO51Dy9bsTolsOmKyrQN7n4CH1Ejzx6cQE1U
+VqN+FKNaPLs3etHPEa5jPnNlbZdMa0tENKQmoKGK4SP6c0sB9+XSYgj6LpzA5pZ+gYZrDCgY4o9
n0wd3v+2OXBExsIQqzeDbqN8hf25IhbEoaGl4M9JOo8yRlIPvDWvKLQO7NFSHB2ujOF7dC6OMGYa
RnCQXOjXmXpbo4DrxmHaLJEQVWBQEpqlW0ZEzAerKk5Ufnh3BB1/cB4WPkP6xRj7gd2cLiiubiTk
/TaTEr2arPmeQOaI3ghNue3tX6hl1iJn35kebS6MW9d90uGyAVuS55RLy7bcymPrRs17rO0kxte6
Io6oLl7m30CcBajOXdcMiXKAh72FFlzjbW0bl/zJjcRxP4kdnwle62oeo4XHpjg5USSO8GGaOUIZ
O1/vBVTRYxD9tG4oLDEOXq2MJVWTyeRpdB+hsr4iGFiBfhHPcplzSwR3Y+KTYDnU3A93D6M4r/aw
EkbcVmw5s9ZsctyOAcjKE/b9mls0WFXRTSFDdQTuxVSuBglPTBzP+ybwhLTpchnQ301pcolKghXG
gdcnFCxvLHBkyMJPyegHHZqCgXRPTGDOF4BQmuCGPYEiaSWJpL68psadYuDbTuqSzG12nPWGSllc
V5xca6e1hdkBD5GJpvbvBEwd1EOUikRSVXsp5YMS3bebaGjBipL6ooTuxPP3PFkaBGbk7rrbNmZo
tt3AfMs60hn3Lz0BGsLZ3z8uaFlD1GiimPDJCxyWuGn9YUtZpXSIDp4EBoGxviW+QKI5/9yOFQSK
xgYFiLGcIVJGgvYRNw9A9r1Ze+wBEej0GZ2UAv6A8OVPSVB6G6s8ao1ksEOjC3puWEtBs4W6IZgh
q7s/SoiqbMRqfF5GGzg1z7n+LzkeCzBobDmASJuTvPwyh8THuzR0EmtA9Z2h5n1GEc3jhgi5+rpb
zKJdQxiMChrcrLV7nC+LLpQsVICzgkYU1dS3Zf7qplCObcKv2Aq5PwT81UQPKPDfOQ5a992Mff0g
N18oa/ldSki29sxZqdb/fdCNdP2q3Lp8hf07xnGKll1jebqau+oyvPKN/sQtci1QsmUSUx7xdx2J
s7GOzmKtYIdKx1Xk43BJcwqe1CvqOUotOuj7k//sQcyG+nMdmmaw5/dVsqoYoiIkav2GYK0nklaf
umGnK8RwAOsis1lYgvaKv14D4TM/46lDFeJUCPCCCjdS0T5adcMtjPJQ131/kTPEd8Fo8qagFAX4
79qdjRCPIt1oha0CNEKGVAzzVc7ncWveR2EYCYzngMEkx+2xZB1PkAaydIkpWhfdeur7ag5dMN+R
zLWLs7YkgVDfLjUt1aYNyvh/+49id/PBGUUpy02CDNyCk7nuDT7WzOKpfymx0WEixhTJllnwtdKR
3ceR/e5RMs3Gme9sYqEYA30enZlCaPFIw4dDPI6UNHgm5krhMCknJzIK047bxUUNk9amyGJTGpqb
50beerM0jzgWTpcSIt67nNzHr5v4kRyRPbkY0FbtMtkHJCzcMTqFPuES9c44xWksTHoCiFm36Gyo
3pHzAZzk2A0o1qVPrMov6q2u9SvB+Lk0+pElhH/I+zWSDk8toltS7PyQgiQFFeWtC+vEb0jaYOny
L4wIThCUj9CFYC7RSG3sIgWGl2e4p29pJHOAn5spMJG+809TFMA23JgXWaBbysB7dEvOnvb06IK1
ZRxX1mjv/i95XUGZt0Yi5POgYQQrVsl9k9jmNX2kKUnVl9rgfz2eqYK3Uh5JBoVCZTjmCQDJpNDP
CwemuTOIgTHqZlvc2XcaDeyEzOcRcYEX+BnM2yYpjTjU90ahrc0d9XE2vMDDPT6EUbMdLRxo5IPS
V60OvlVZ0Uj57qigA/kAe2FdxolUAjwfPbJaLAYR68NPOvDJ/xhlv1KXFQmPlnTZA48O4CxRodcj
QWq8F23BJu+rJKbZl4B4VEL38Ca+DFgqVnZfuNKuqHrX/tCAwbUtslvvpEvinJMB5gDKoQ4osK3P
nPjaFhS1sJFeZPreQS7ggWmCq+MfAfBgVfuIW62GPxg9rAec6MtLEkPddj7D17eiLrdSJz5ErP1W
g15721hvs2nUdKSWCh/9aKJQLj0xX7TJlsRnkhXmWYftYVks7uaYzYbeWqKAiuOSNcrgdwbKp8We
9SqfbK5/juIowqwPzTinNaYy7l2TlUH5bUVt871CRkzsSSeaeRauYoCGBWohWfr9jLsqInOdCkPs
vnngMRpcsvmnPpWyBPdy7o4nbkyIOKwGWWIB/YAP8ZRlsB1UfkJU3EFhlzXJoxP+t6YQEKcXuBIN
y0zUtanYjoDklX36MLkZY+4oaaC0eCsTwtNanQjdSE5ouBKHWsSGjD+SmiUtCpPAwAxzJ4TdhwLx
Vb61Kii+h/ewpFhj73AWBF2Jk/bCLZ+7oLHIclQqNG/j29/1n/FEair57+BlxS4aUtkh0oxK0RkQ
7bdV0wSS/YxIMnRsD/g4ZhF5+by/qX4dDEZbrUm1YKYuxdJWy3F5POcDRZ4JuJHqkxYoEfN3JClR
FK7/5YGcLUVXpIihO6GDSoQM6hBHodAgXBT1R+q9hU/fS4j53QwN/1CKKPN3+J8D0MwXvoA59p8N
7RSEKvI6CBfOdZCwIfea6Md0oSsDx7Vr6S2R02TIsRDFtfL7gVC74U4YVIsE3AwPPEhksmyWDDf/
+ejqy46+UQObz2mRBiQ21LVXQGBskrHTlHRwbzrGPxMOMk7n3BG6cDfzyI0JMY18GtTsrRpEQvRa
eEUPrOQ2a8k20ePAdGNhDBFsnnC9nkwRVHuSTvFw555bxtwezLc6sUailwuBc4jLyvlJgiGHgD5O
zVDlBz01O+bfVHJeWW/XGJ9m4qw2z594RRTOMyJrKoCqoGohAFTArtcsUQTzqd0lTleP/fcA8787
Q/VEaLPv2dTKnunyPDZEBEMZfNuettiR67GQQ3D1sabKm0kKDIZT/68DQIbn63jlQH/sbdt2liqZ
TUb+1jxpt7gNcx0iNHOoh+oqCs54H2fPuu6aqx62WDGkbgpxd/Vyc8JiKkLkKW0S0s6LiQcGHCtl
xge52FFL7ftB7ZqwP5p+jMCKE9TQUmUT47BnKhqEMpgSGVNWgshlLqq6UK0VLiCCjSDe7LmEWMrw
k2lmCDylZBb08RX9t2eykvkTp17SuUyXMFJhU4awfIM53ubb9i0KicuYf06pQVsyFGQ4l5rwT9IJ
jcOA42V9l/bNtD5uTCrBps1lJi57TFwRXw/rNQb77nGRkaJ/rM3MxT0IJuPZRkw4OGdpRKsHHvbY
fiYjuSO+suXIle2fa4Ff8c1kpw5EGo1TuGp+shd6nPBu74XKs0Sxh6l2nIf5WTrti6DhjDomrfdo
lVRtrq0/NR3i4BJsUV4qx4HYtE4dNehQhSH7OgQTx611HFH2KLa/N4OvTrpo3xad3z+QxLqblq8+
mt97T6vAO3419j4NgjK6lSvJIn0DiuqXZzU1uWAgQjWbpAQtdeqMyYsuhkOivLOKgC94aP2miNZJ
4k/ZdKnCQ2l5fF5/gePkV92FnxzhOLQkY5sACeK95sMTR/gHpILPTPARMWUkjlct66rIsBiZcBHF
9sZ+1qBrh517E9/Y/Qj+Lm2tf2TBgeqWvBL8AjJ2GQ//3flbfHfd5RWlKQLkyNLDZFAxxsWUKPCZ
tRR4b53kVgSLuZ1JHOVbGcnYENjJlHOXsikcPTpuR/Mla/ghoJsAL1slV8shznzSw3rqb94Jjw8F
EhBk4H+cP4KrbJ2TIDBmPyxgZOQFyIrDq3wf8r6lgqphOiEtTrcxZBZ11nTsCrl4RkuoS1I21XVQ
E6C0OowmLQVzu0wsvX06kNM2hMaeEhzBkr9mRCT4JIG4aKaAVxFO0m1Nx+o7eRkCpy6SadSA0/ed
0LOWnDlwbsg+/j+AiaGLn63uugsMn1LLQaeS5FsRntasbRmXMYGEY32+DzvgeEKT0FaqEwi6EGX4
vnXTddacP+aKJhCJ0m8jr0xe3WpbaESO6ahhwKKOOxPzTL4S9rczPE6785Pv+sZ2zFOqVv0ds28b
Bwi2jQJ3Bpo4mSBEybFBSUBqLbesed2JuaSI1gl/pwCtL2qUTAgRbW1jGxBbv7EPy6gdbBOxYjNu
gMFtdTyzO0/XyAwZLOkLpGBaVwpCC9BJ/HogNz22YQnER/DjPcKjiQ6DtCDnm2E/RoDbZy9wgC+H
4I5ijPP6OiwgDBiRjMpasaIob598hlgN37Md0FDmHO4t+8ST/LUKiY4BoEomG6MTl029WmUcAI+Z
JK/WN60xnyNkVMoDi/Gqa/LWQd01GE7DtpBKYF0Ba2PIVctMT3QY+pLHoYmuy5WnA+TFVUbrSdOR
YI41nNHre2Xa2FF0hbbXtWn2+KE0XfS+dfWv1Z8qS8UXWjmKhFysZpY31agvqtW+jeVUhwYBRED4
yuqOT//J9j/FTCqFyB0BnH208aMoWHHkLCwq55HvCwHL0Xq9cEzZ85Pk5Caz9KSFXVsWh70fIOQD
lK1brDOG2FO/AfYF+M5L6GMu50LC7jwNH/MVxtQP8WYSRp3DPMLp7xtIxXqMZ0fedp4nV85Nxi5l
LzGQJb3uTSJrZWg6K+QieloMjHLefoZMPo8Zj8FqjkbjtHzAC6VfAEYBLJ8e2NWtrwZyVJER7XnN
DwhsFWEdDKPxeih7rZUOzwHof8oyvNSvBch1kG0DFRMr8yGbXfYEJ1oZakppEPdtFca1WUKLaS8e
37dB/s9Z4IPn32dIBXJSkFkPedRJDXRLjPGX3oHn7CSJYyYIs4QDgFUJerri0r6ihI1iSlIWgCqr
hRPSmvRNV53X6x0E5nJEVX66WiZtBHfDV2akQHmMgvLjUz1lT1wRf8WAS51xTQw0L0sKMZ5Pt0tI
y0KuOGSQpP6TJnBRJJvBVDAIMOq0nrzNOUAX66F8OKN1TNsLJ4XWWL7YWqB5JB4dopSNIIJadHTW
DNSH0426zQs6+3KQOwIuMuyNZNrCio3ghe+wGUHEyLzbwQsKwaxZ0IvekcpsQGzHTS7Sq+NmiOIE
zZwgacNWgAPBRY2DnCrF6DgEysgodXfxoAxkVT4ufojjj21sUFb/jrs7D0DkFdVfscMKkTVQZ0eu
uscGFBHixVLN9oIAIpZYH4B0TBrVBvK/WZG1Q28XFZldF1mY0A7z2vaDQsaeu1tbTnsvtQ5AC5B2
nwdaH9giKqF+MDYqEKjb45ZuXsa/qfXn1UVd+KYIso9rGP6HJyAJEU6v+NtYuMAwip6JRgOb6ouI
cgpf+Ri06V+HFFZ57ifxLz1fkKGpoF+cFA6EdCSYpxm78ZfkgLiSWZwXozEhHq0EDUb+cbLi/k7o
gsHvSo8CQbKR6acydqH0uY3vYZiOJKEd03Pqym9kuYaodZfexiLdH2Op9c9zcGVifgOqm9UkE+6w
SjXaaAxmkQ6JQuHZCpPuOuTqf1jJFs59oBzMApqSd4mhrWQCyRB2JCORHdX+H3zX1743tQRO2vnB
Mh5G5Ec8N2bYPCiKFlqRVj4tAbxdJoFlGjpzb5n809arO9QV2Q1hYQsEjcfY9Mm8oBC0kYgXGtNc
r/5pHkG/9Q8CzpiYmygQZtLrHEMyA3o4db5D2EFApWuNO5hZ4LVaX53VeZGVb1AaIVQmzy9v2u4o
P86VbPBPDXeaVtt5HrTHFqWkzd3hFldKvywysWZPbpMCxjvNTHgGerGiwsF8Rc6xXCnNA0Ek5kUm
S/Mc1qrxI4h8/xtk7Dua9lPQTs/2eRFWOT0AcfTTg8Sj7eX7JYveZ/eOZcedlpotHy4Wt3RfOm6I
FVemNnhEm3WdQun3++CCktgpxQp1VqoO9R9MumJ1agwJkTLAmYSeV/1zeAeAuMCC+hKEwm+aiCTz
XQr0RRttHN0KQMFI6qPq7GHxewZ7e4Deix8HGIm7IrGqSEYzliXxPhkAVuUjWvweaImjmqSWMdUH
gPbrmpIWyr1V7K9HlFbC9Ly1FYOBItQvMPsvnU79zE3XTI8h6VefuE8bHN5sHQ+4SBmjz/9x0y/N
ZUaVsGriiBNRO7ljk0QWjiGvSbH5qbUOd3K++PR6jXIu7mjt2bSgHeLEbPW/ZZljJUZluS34ycyP
b+77Dw24iTY25aleTvd1RiZLVFsupIlHzHVfe9CKEotbA9pD6XpE6Dhh9A20EB8h7APKLmTAuCcF
1gLARjNFE/0tdY2JklXzrnVthAAw84PuRfij+beELIU6XcTvgaQ7Adtzg8tQa1cc2ugFams2uwfe
/IHbbaJT7Je7oaMI4ZrScrITe51/gz65kT2GuiKIXqrMASipbFXWIF0yi0Fsw1KkjrWO97dHGLvJ
pZWxd/Lz2uWk6GJnSk1JpUqU3f/vcdqkZ1uXvzWVa30WVJDqFGRy5DmwBNG8YVcljqsHg+asdRqE
BnTcnNDR/1ACIwbNgmS/KxQ9LCi0ng/rQ5tvfRbvwKwY1xnpa4HZLDlLEZZ7aEv0eucmM+OP32uf
uRDcL5BTLtkv+O4sObm7p3i39vWmaK93Hyxk767fABvTL2v+dx7Mv4xScpQeEdmZYvb27zPk6tti
ImIXMoBMJ4vT9NiCodjFK2Yo1I/4vKLTJ2TCjNqPhZn+xPxQZw3RYXXoak2HRQ6MI+BugsAhOFNO
QyJUSE/sIqZBuq22JWZa8fIRYAGLuabWZJWu/w6uWjMQdnw1sHFzvf4uuZJKCJP3hwBmwaapzSVp
mfvSDGeDEzL7xtxh83AoZ1+uaJA4pMnJ8mVxpOFOndoMN88kVLxAiRyJPi0aV+o4XVOjnu2gmvo2
Dx0a6bVGBXuzKn5cKYKfhP2+bgmzzFqLWZ5aJX08rewn/nX+PbkbM6D8bMfuAfEpAb+9UhVHk3LT
teHnLufEYywp+unwAB5qpjzGW4QYJGWBb8zXpKSwXuVBr5jA94JlvseonWY4oDgff8CjRBLhnUbW
3j8LyMF4g3aYWMSvBa4by8zhZIVdd4oRXml+ZGzn0PSZ0otJRZ1xZPKXHYtuR70ES0VsAHnvMw2V
vbRmDrDcr0b/79WH1AVJhrF8YxoMyw/mG7lTXCUiARn1gH+s7tmjwc7hMlyw3IfEXKBQdsFVC9Nq
h2grEim8TbYzEX3QXQiwp4M2VtI5y7J6XW/wNmBUE+nI/gsbISMT/yLqn4TdAxdHcELmemggz97S
27rlpICKsXEuZVFDU0ExXql5gQBfYWGqVJPOVhLYCSO5lUp/uyDnqjCxcNcfhgKI9WORPUO+N1sB
7zaoLnrTDeFLZj6C9hbwxkFPhWAs14C/YTUfuOZS/fO+3EmL4pIGKFXIWyvx/GKx+/Og+0ExBslJ
RL7bDMmVlgqzeXozgSamCFozNxt69bb/7EG219A+E4GfkZo7cgxiDHkIUVMB+ftu19Ttn79RWLmx
ubHvaETKyMwU19xR8DAt9QADgH7ur/lB/ZvbTQDRX4pLfwh28pK0iwhSg2jFevtYKc1Gm0q16bgz
jb7M2NxPOVSYyaO5VJoHcGwGzBLomG+i8ZlY3j+a6M9XsJnA/qPpczRu94tPZG/Af6WWxo8w/lYE
tPFuUY+9BqVgIo6hMZX6cDzJaDgrJLjJDhcgAmcqQmXzKgitaj1ip3iDT5f6LeSLPPZDIFa5M4/1
3CGgs+70YCDtS20JZvPMifXDKvvQLSKxiWkWczj9xlpECfXw1nP8+YQzCQXtDOzvu6dfsrFshWRd
gsVGUdp5ttVDxUND/th7kkZm7IDz0Zc3uNmw54vhfe99C51H0f/L48o0l2/EbGj50dPFG8lIM7UU
EftdEQ4sLutD19GfqXXt02v/qpEwW5GR+A5+H24LRCgKV0tEMZMfvbP3CPPKUqBqHxGMbWqT8xiu
qperHaYkZfahvyaB5mAMYFwFMQ1gpl2j7ym6AGqr8iPXZyvJsnqMgaMfZ0Ez2CmQ88E9zX2crPG+
geGKdtqHnkYxv7r5T9cRE05Yt4xmMENVx+2H9CcTrcK7N0ap5QFurfwf27Du3M90iH36fezl/hLk
DmdStSO7LCn4U4CIj3HbBasX2RRJO8uqeObF7EzbOCT09M7qpOsGDDpW5EXxWXjH/X86fCfoorqd
Izv9zVwS4O8xQWK5HoRS/inkVo5s1KSXfQlgC/nLyiI2eXkUOYNF9JnPRtY96xiQzFaPt96disfS
gvvRgwa+xb9AsfXSFg4/cEB1W2sv9/Aw3pjR9SOGP3JcGOr5fsG2P3OYdMRfjOCNxAWU+4kJbqAI
9trNPPY+C8bkuriVppyoqrA4lXcOi54Dh6Wz+3gbzxv3MWKonzeZXAXaEHN+vBkO5UEH1mbeDl8C
KIsKmUzHsy/CyIh02z/RdeAXu6krjaPtsc4Ipshoc7VOzUNMSQAwDN3+BIGk/hx/q5kyLPZ4AxUX
btOG/kOjKOCs2hv0WR/zcFGBmSknBezvIhV9ySlrucZXyS1yYiZhw3VOFzOuoUwHMp2oBufKgofC
dYjbkadAMJLMQZ0XoXeQclXoiila8FQt7x9VrZKXUXiB3p4NMewi08ioUx18kZPvglCPOSvZxocD
B0oOpfhrNH7pPTl1sX+csXlzSu0rlc7EcCzLq8xF8MQndxgh6jQbV/n9qTFHjYUFybfaf0qBnjyC
EIyqibCsCr4gRzK9ereFRhszdJ6wCZxoQcVupoe/f8iFdIHol3abN522dS16DBRlE70JXkTHBS6E
v8XrWKjxsRmqKcDuorv0m8z8Yr2F5mDwy9lQ0XZJloZw+IsG7B2Um4/UKSQIHkOXxoH9pCDOAypk
Rd4oDdkR0hC2G3GQbPDii07xrq/A0XWgECw/mLhNqxwL/tMqjwuryiT+HWUAuedXl0D6wf+TMZYv
+uJ6FwUOj3coVCJ7eqO8yk02wkYmnOLas1BjKrREWwOaJ1kUh1paKc+p36pij6HJPFCOrSbJIHug
XUMEMItgBACYu0ZjzdrujmqBXIAXUcRRmZXN6LDMywwbwCc+nNEfw52RbR7saW9z9C+DACA+IutQ
WNLC7zMSFipfKDD9GX/OTC9FOKkbnkvL0Y2cZm6wlLg1KoM9yO6IgGLzN9w6RtcNl4e4yrvrhXH/
gUJMmI0f51aHAvKVpuUoNmLPLHhzB6OJTjFub8yOTjhEwbRUPGkJ4exUkiZA6xRkrrsPklNv3xks
tMxszzUODTFdXefvjEYUNhM6o9l+mERret+EzHVfFrjdmuMVCMQflaOBNcj8wxxEX3FxuKFKqcRC
Ecxi6w8cL3oQ8bq7EKM8FwkVB4sQzAwmpsVau5gwhXsdcQmn/58gjT/+efZRBsOPoS4krfUMpVg9
YG+ayGKt6x5vm9PUnzKlguEru4GNGswZw+XW2C4irijNVAGFUUEGMURRhg2J68t7eOxCx2xnuj+1
LIOOMS3C1u31XYmoGcIlnNBop3efMOZ67XzDgJp5gsEUo/qLVrIS7xfaP3Al4h2y5Y39CuCHwBMq
zmTOTgkt0Sz69qTKm4OUZQPdJfYV8fR2bHw9ytNEhkDvoLn0h6AlXm6gouPK3dA4P3R00hRYkpmL
wtwBLoa62cAFdocsQ/WGpCG4cZ7ReI8GAupPRjrFe0msFmJWUNhy+YBYyHu1jX866pey/S/0N/0P
crP5aNdWFUdQ9U0Mc7JwSSstOY7GxYc3TPlsO+abuNzvPIqv72PPHgQERm+3Ni+lGSsHX0Ac9o7L
HrtP1fp+jVGF8/Qc83S5wYldChKxyew9abC7Ckvhto0jHKg/LlK3mIPFJ3XdRPZw/M10JX8knGbG
1ubjY5u2y+kzUjnXqh/9uwnMnJOCbxpSk+HDVREa5zmcXWi8WjW+d4HkZIXqg9h4RLwKDrefrvMZ
XVyZXv6SlnYqndOTAKsluyk2KnJuIIuCSvy088SFPEIhosMhuuepUdj3TRGI0Rh+nOXILtk20IQP
D6YDsDXSITTrQwGpDkgJmIFeRXXRSyjIQrWFLOg21xwfcwNTHGE4P+2ZV/5vI97J/qz6m1aLY/4R
6HBl1ln6DJxiUd86/WOM18Vhk2D9lc7Gkac/eAab7fPnFD1NWkDqH10d+kt6aYDVqkIoyaqvif8X
1z3MZzRCnRoYyce74HoNeLC2WBOP329DwAOgCimm6uPpq72zxkim3DaMpZjwXZ0uqN7vFdrjd6N0
NKaxBkhiVv4LVxNONX5/Om+/zrz6iJYqLykJgYYzK072/nS6twzrSfb6n0jYTurljJXCBmnucDh2
0ETHA2fYUE67lmSv3TquHfd8KUfsiDLjDcUUHRU7EEI+pDV1jDcvZoQKg2w68DEB+sk68wqfW0uW
vCwObf4pB7hI+DEFYhwY+OR/6RCitU4WAZd45VUQVfyVDCivNLkg1eSBK/+OFi2KXFS3GlwohD4k
FdawKVSDhe16jdHBHoMTYk0WuqulrKHJF+FSyVQp8xdG1C8ieJo8VEyclQvoQydsIMVaPzR7pUvZ
+7fEBCabn1QZX5WmbgPrR9Jf3Ibj7MwM0Ad+qJf7MApaTc3X4GJsla5C3go2UdBhyRtZ36TYchEA
ipXcuP3Hy/C1tNJSU3bW1+2BYwt6179+qBa+0oGGCp4ZWCwiVlI4/dkZmixSszzDtuY4CSOhv1aj
5Jw29dnZP53GEPkanWPsTeplZD7C9pPVBe3m4GkI7/4E6Ofcslt+oZ7ZcvsbfhwazqQx/V57uDe3
QaV3akX9ox5XT/Bqwh/6g/JUZA7MPqvP9QnRUGCyuVS5s59gpeoLuuzPpcw/kDKroS0lf1Ifm01U
yqCiPeZHO2gQnNZzVLj5M1WlulvnF4LxUHWNyV6OPmbCzprv5OZbmrEyoN3B6tE7u9BOcYIKgcfE
QLBlF9J/+NdCd+6yCiCdUNmdsaiuOQ/EElot03+EAVqEkaMGYqdDoxsa9teumBekZ4L/92ghGkdb
G1pG4/ajINN2oTQ5o92LxFiuXucTSrxCTBiMxU5iIaZnSx/koXosDqdroyyfOtzJGiwZVHhiK1FR
KmvIDecqgQinr92jvuHJnCblIIJXG4gejF1KdIWrv8gYSeOOAC1OzRLY7UuQTkSvab80Jr3W3QTn
BFRQUxCHg6ceWkPRq2X0g2T+Uveaw+9Mn8AqNc0gkzpIFfDvKNoUJUFzG7iejWYBGN2BzOFIHBV6
DVTKEkziT2aFSmASD3Os+sXHUGz/B/Y9rdTjJBO3LwYVxKAANNezjINX6nx8bU8CRmu6OUuw8MQH
xR4cLcR4H79W+KQrKe/rPGqJXdbrjtGSTB0q13MRmQxSZjBfMugSvIuJhumGzS/YQs0nmenOuh31
kkCfm7DONLyduK7d6gwgdLOxNWMKpFEFa40mZwTZ4RppPZ7WJan+YACoaNxo1VVMk936PNqqK0bg
8oV5cFr4Wg8m6H8A5gizVJ07sZaLw5F02E7C6sUZl+IBPiC+Pl5wsxfJYFtPmA5meTDt1kmW3Tpq
04JcC3Fb3SceFVaschej93WYKZtC6V5pua2bM9q7mIcYPklTqvJQAkFbhL1EH8X33SpdpAWynFWa
/5tHQjOLQyC3ucXFmyx84EDrz+dW0Dt5jDjiD+7+njFl9oNfRMWZGP1QUzctxd/5nARsbsjC/ss4
NQp0YsiX+4at8e2HRO3GOrxu02k5mf78N0WYZlbQQTPuRsc307w6Qw2zc8uY5hujYH06tOXOwbMO
WWS5R28aMuExwGB//XVv5qFTyyR9oqPDASmMFbq2YESuDUXycv00Bp3IokOcrhieVRoZRIJwcwq7
kz4b+x28dxPPo4e3YaJ0uXNEhEBiY5R2ibefvNeBA6PN+c//iR7W8WrqLLv7BDuDXbfaNKMNYagz
R8HuRbYwxmVZHJ922RB0rvX+SZ7V8seIgDWwMmvWw9mJO6fDVq30Tu5YyEc3qQswVKLkPy8kvoy4
dMnsPeBDdAwtb4Ub5jJUl3mj5IIl0YGhMVXBOnuYA8K6UC0/Tkq02GaRAvHWFuHBx1lpr8g2vX1Y
vjU47nlpQVKvPZq9SUUN5x8QeA9i2lkWDbvY6m2cgnmmdBHuWGDnQ1BanDU/wZon1wA+eufEd+oq
p7sZRjH3+GEHAC54k8dcLWwgDSZyziBxSyYn1cVTI0CN17jrXuzjtxaKY9f+Ht1TXvZCx2x2ji2A
RHORwIu843+8q/HRwT2XR3Rry9J1I6SBUTTM8HcPCpLF5+/u8LThvixBPmh/GqahK8gNhSsDRTb2
SeUaXiznhGiqW7ni5xvi+z2mCvITaikbu+H4kAY5DPl3o8GPIeMMb9gNT8CSITiFssAWgT+Ts6u+
uDruU56RdQbE6VQrQAYsbTHaYM8f0BrEVSyp2WgVWDQoUSaKJUXsJHP6MyKa5we6+i29ogmjiWZZ
dTwxh0M0JxsGjsBQUXbvc2xWYstL2oudLdgwa06EBmZezF0hzf2todQWtBeEn3IoMBEK1cKYz6xk
CXgCRNog2bG74UQWa5L6LC1SS19oJ1oLjmyXQ+xXn6cABcZW8q8X8Ca+QaHNOfu1jVjDp7A+D7It
S5fwpH/fBWS7C5kit2w8go3yEv1NXiNUSEDLeUh8E/jK83oxO/Nkvol912kcb8cAiESo0t2Qa5br
X7jdqSMLciUwKIKk0KuES8nu6h07T6Kg3VOjaVW/QjzETnHNm4OaleRgQuRhCBBHQvyNWo699bbl
hjAHSzx2gxWdprKLcFMy9EfV4p1JUnB1NTYAp1ArfNSeN5ZRgBuFej31InJ0yvu7KRJf8EZ+m24w
Lz/gm/+6pSnRj8YFE1j6MM39I5V8uhpnqvTfh7nCkIxSf5LXvX8eI2T8V6tsvmdoUYlr0WGQ0odD
tGmlEXGtilqDmAwwF61nvY5riJvoqw3/qJ4aTUjJ9Bx4gJ9cHvcfcsEHoOXfgVynQYNH0z7u7CoC
w/12NdQOWNGpucj6wVZXXfwSBRwhXZO7UplwzxmAdT88nB5E+IanT9CcB9QoANwF//tXMc4a32xy
DmWZ6g/MUIW7Ie3zUgxEU4uu5J1TMkSuyAMrMIfRsVLDfQI81SZ8XYnmGrBv3ZTzidebUH9M5lAZ
vSDPYa3K98z34YVQ4e7FT2lx/39JyndQcMo4qtjy9HL8krXvcZpIyMm96SXf+0CQfgpe5cQVNb/s
tVToHayg7ahaLNHk7v3U6afbMTplTedznKbwRHlfqnMGI5zgIf9ZFMdMKg3BUKMBnR8nf5+xjnTi
3DpmcQ5QRUymPKqfp04bo0Y7FUi1Wcfh3naXwS5gpBBJwF3FmcxshGLn1BOR88NAyTtpaJO2or1y
uNzP43eNwMNZ3/RcCg16d3s2KKurp5V01Vlniv5TzCzJ/ngq0TMNKMxGHMsPvejNE09I5eQSA96R
6PdGk15mpW6zYhnRqiOmA3ATnS+sZ9bazYcULhQVwD+woHzDn/ALBRJ9hueOFycUAR8rTvSYqR6P
UVLWbfW83qF2D7xhAossUV18yKV1mElNuMmh8Qwbo3610HGx4xN4nG3ga+V6skZCTPvXOknXat5n
Y/8JrRecYhGXbK/okrlFpxvE1PizcjsgVEc+nLt1NoE0FjZuIxNsIFaggV706jNKiQJcgRIL+dtl
SDEC26G8rO69kCjJs6+Yo0zg7KBJqLhGFuAnbEf6o91cY3VYt/NeR6PPAwvf1HEk/GmutQdPMmwV
crAgiDPurrqND/meI3Kx65WqhTkBlOi9dGOlVsjlLWBglYo8Dyt+DtJtZNoEJzs4bvOKPGt92Ny6
auhoPYWYe3C7QiklNgo80HwAepqUzTuqu1+bNJwobsRQzz+30BtEK9khuP/Q02m6j6k8g6Ykf3+8
kd7T6zwjNxBp8i0zMqZJB0zP44QoYNfRdlAjDPsIA3QcmnVHMGRMrAMkRiHekCWJMLKIyMIER33z
FLHx4Elb+2bsVyT2xrkl8zWwuop5CMVPn+RTDYmLV+vAIBo74DL8j3qr5p5xfeOlRhb38j7ytfE7
XAOFncpYFGHl22nqttfhQ29VWf10ju0b9sn2nJfoMbFw67H9HL9acbemcaMJ+nKC47dagtuq+pFE
yKhn1f5qngnBFYHnyJL2xLaproM6CbZrsfYbcr6QNfqHgSEHQlj3ktAadhG3D9WGABD/9d6EqlNq
57VQ6CQi5KNiC6U2790D8oaPwWfslGyN7GwPaa4se7iG8wF8uH0+ebv0nnoM01wFhsekueVQe769
9h45qV1J42twskmBvFAMGkSDrfz4VfDMrYhuPNQRIfzJlNO2wUVDyEgrF/zcsISTSzm0HkhhdQGa
O2Tq9SNvqgrJBH+EbqbEQpT5HrFjfqCYVp6Fa6wwxZypFXmmVrejtQhUfZNQK9jFiWq2tai+ytiV
qIgKlSN8VmNVnjuhynNrI7eNQQUVe+BHzTClKowvCUSx9NzR0dl7piV5xVCqeq0F4nLTD7I22my8
kkQV6V+8RdksthbMuhulDKT/vlzyY9NRmZ+afClMidfAwJQoos5bLfnmGPS1fFLt+LtpL/Tcd3sP
Yit/P+FvqVrfTuVseK0jam4bGVEhMtT6S8JQvOax2PKTl73NBT9JQmU4W12FOGtJ0QOfwLoNN8+F
l0i8h42fJzOUxTmAFNoZ+WE9hKqASF6xhCzEdecFK4dORs3cOk+3pj6HEjZEIGqfs0eAY+iw/YUa
iubDAhm9DS86jBcaNRFdRkIU/VV7xaM9A9kfjGfo0Jg2/ed6vrTzL1y/81Z9oM1oMgSOAE5A4KdG
xb6DMqrf1PVMFxX7CD5tuFSRwo/R/vcB5esjSrGYvJjuvP4rF37lo95dFHCa1bZK3HNDimBek5Gk
aQVr/JKJGZgvD6fo3CNiBUwgl9HhaKfnmEpb42Rcy2IDxJE71Hvmtn92EyznnHaLtxwbh6+4qBHE
oGoZhpRl2xEBKGMyKSyIWdVvRUxrOMlKCgRAm0wlCoveSRpwveGh0O6p0mCuCJzKiR4qayLLckPz
Xsi5Dzh1DIRsPvvLAat5pc+vhpiJuGG6pNcfw4eeS+BuVYS5mxmVADfnkBbfn4z6SeEiyhEIrxOp
SdZca6aGdKLY+LjKohehux23E9wMBqgPd4xpv412vT69fCCl6+gfO9E6b0+xW1zvB+LS4B1jbPKi
tU8dtpYf4rJFNujbTxO+DdGSnK4opfEkuizto07TvH+APt4W2s6Sfqe7dihFAFpqVWFBUL6xPu3A
Xdk+firrENb8fS5Eyj6S6S0BG4yc8YyFUVFhCDAnogcM3kXh42L+4SBcBL98MV9ubzG8gU20FZNN
YZyngm5Pgkhj9OGege1jbJwB7XxAGjUUFs/b3/I2J8J+ihFD0TaVAkwN9+CioF27c8mYYHCjIqFY
8Mymy/9S3n8BpnhwJXR7Zy2chQbjg02Am9zwuUfhlz8bt7FU5xkJr/+mh21RbZUgTrXgMYXaPKSH
h9240vCZDRSWCDyv8VT6tiYkSOj9jCCWhGT4vIrflhlJgVYE0jAn2HY4U/ODybBzPBSFFlk4Q7Kk
X/fy6US+ZX8IlcgEAsSu4lkUapectQa/RECXHhvJMlsM/F1g5mgq8cDKUDn1H88pANqtPzeuLqus
mW4bfpXaR6v3AvLX4woGeexFpiRQuZm0yQqIQcbD97HLPRM/Ubp0xr2E8bZutOw+5LAEjCb6l29P
FD/OUGWsK9pI5PB5FLmPGmOePxXYX49B/NPhjDm5LZhu/sC71Ej31kXxe3XdKPldnKeo4iN2xzFP
ObXGAjhDO/8TBHSqF2kuktldlKPzmsDwYqqk2kwEiIvfS7NT6hYswFyXebHXVNQ6/QWmLho+RINw
aS/h1oEX5lB/EImngAvxP0SPljclCKfsnRQyo7BM2FWwi9bBoMl89g0G5bIk5Bcq+AjHcFWR89ai
5TwNg3h0KH8LyUX9S8poRu0VXMQ8lL81w9QWDs60BpmhCxzWBvBTx9nHo/jj8ITBnPjiZ/gtnJbO
n4+rVlJJTJ+UEXur1tNdnsjKCuU9Ab1QishJ7wAL6ZdFn+2k6RlvJjnz5jpFkZIS33muddXAxXqK
cjBurvhWtS8R2hS3Uo9IhuYMFy+wWRBLim218xt+/kM/H9sA/lfriiuglNBxOoRBtM8x/sMLVCsO
H7vtfh+xIxEbLzKAZS9yiUI1HfUNX817s9G/s/tjcC+lmrgL/JezdWbgyFuQJmKOxLSTrhRQ/iU7
+fAVEt/URd0ztEFG9FcQM0FMwL3MyeU/0rlmptmcxE207TxmBdMumeJ9LzAoVWKiz1GOtIyz5KzB
CSFWj21KytMC36wTg15MmOjjpnL3A2pifoobz2o+GTqIZWpQDqcPkZ78SpzxwUsAoHp2iYUWfFJO
e2euzDt9mfWhTEMLwAkHQasIvaxokGJWNXPGtM6MOU/GO0gZyGU4vY3F38dvV57H2NhQiC1LoIGA
GWWPF18uBa7y8nvd0uojPBDpTl8Ydim4+jjtICnVWHGH1dsm0tfqU/h1T4rq8NgjqLGLhUqlgxxF
8uM5Qo3kE+N1iWgfICxfA794zXwBd5All9isaGRV9KFk4WRKtTlGyoWvluT6RaFnZzaIYloztBmm
kskGIdPBGXrkSqcx/iNHKrZYzaovFPyjJjrXj6LqAhYXWOL/PDW0cJzthGSwSVGm3Hx6gxOfXQeT
sjW9GAEnY5EIccmenxnXGQHhvbG9YpVkjzAIdGrDE2/cl4fXg+yiYbwZRwjqunup3C6uPsWEuiLi
Q/mu9TwgPXA7mkm2KLqkBsk1wAR8H0fKxaShoR/PLOQKBE4Vfm8zRLUWABidsxsk+bI9BAFuuEI7
azQIZsYDYKFwBfjL0vsGxT0sZaKqDWQHv47FNI8JHsKf42J9mmU8KX+53W+CqD+IZsAh7niV1D1I
jehampmVesX+JKPTIGokF/1E3RCYDmkZoqm1iiA8X1K/ia+ksc/voJt2Xx5Wl08lTTcVDA/KXRyq
py0LjGs5QviBS6FXjKjtjqYMg9Avs8L4hEc/sr6Umw1XaLhH1XL84aWt8XAaV5WChTIKS7YcbR4/
ZrlvLYM2ylyZCXOOtR241Au90Ug+d0yrGpOUV2KDIT2yLk7jqoH2qD8Mrf9QAF2+3+aDWrX6nlV6
MOL5ycP5Oz5X4akQDA6LvrcCqhvvEFsC19tdR/MS0g7Ea0b4VdoNUHARFH8PK3nAtWRmEhMdiMFc
IGqi5SUNs+OAyLvPsybFTMGsTin8aBEdfk4oIRhyMSlKJ7yIIt8YQP2VBZ4WskffIEn3oXyK2Xu4
L4Ot1TXw5qED1F5llgGnWRb+ZxjrbF6ErRRJ2wFM6iJ5rrBdt3hnJDueYfp5sVEpa07Dq/xxw1ll
fKtrbkFLk9Oq1A2P7icXS+pVdpaEXKI3JUCkAE2j34VDQ5No42JirmFzV34S1RjEUzVo7RxgkIV7
KU0UgeSZidtfDMYlvdlI2JMfSXvLKxUjpQvrKud0QjzJPVm7MC2PbdAHpwW1R3OiVaDtiX/U12js
VuGPhPeI3rtzg39y5fH8R1GCOrIhdiSnxOe0U29kbau5va8HF39tcreGZF7SgCRFySOpEfZfyH2l
+j2V2RUaBcK5+kT69lBfy5O37A4stPFzxil9wa+5JtlDW/VwX6OgP07VKiKJeaO26dCqfPjBJvtB
R90WBhgH23OqYXPochQPYEzYQ+2gFPDgSDIfei1uEr+tllGoBUDpq2i3UKbk8oQK8jU/XGsmrSz0
nVCTsvXdA8dyhi3EQa+CyLZMg2tAUfk/vApuEwyCKVEDuJMHpGfQDI4u6d+FlbH78IKO1Mf12uXS
GOUBxeQPfWFuCdGxVvpoYlmCtDboOymkfEw8cKuM32ywYYhUMDPV3th4zJQy0sj7nbJaW8QIo8B1
TtWtyGgHzSp+LyAlXgjrimZTg4xu8thc9m59G4twFbJ4eGmshf+dyK6Gl8MN9UlZrKuSQlDESvbv
ODApN9YVH/2uVo6TNS1Ge/WUcjlxZ790EgeHzQDdcWbV1davjxJpiNFZAPzIgIvmDXjulXPjdPDJ
YdfmZ2H0R2BWOu5euwcL4keaicszd3CO9VUf9sgUJKXcibQ1kmjjzQhGDZAQRO+9pqIgwJrPFMG3
7drx82kTQZlgW/bmtq5NRDUflTQ3lsvAq/UzMay0z/noHlBxt09A0xeYZFOuiFERlof6DitjGlpb
GUIMbyCcx9ON+LcSEUIR03COb1/WXeKv4rBXTLjjJVJambxH7SApLP7y5mWIUqO8il+C/1KbcHjo
F3zmlwNhjD0jD4Z4chKmJGky/Mk+E+3bA7qPNln6zvCZr4d74bu8Cu4432Ulv2v8PJGtWoj/cx9c
NmklzIIfdJFLn8IIcX1eQ5XaU7kJ1Qs98nHQ6MuRwB8pFXmFPGnNQbj9bwMXkQiJ66GznItinU7r
C7L4u3V+9gD1nKySjaOeGMGVYHg5gz0VhiVIudPtBUbX24J4jG76K/jAJQOiu6FRRt1MEELJfo88
0XKSUuzb9cjD38JqiFwscWwlV2lgtv7w6UuFAtLb07SdW4cQLIdqCsfUNyrJmhoT8gKaIRFwgURb
2S29dOXgdKk/g6Bo2Z4dJcmwL962exb6Bg2gUQZ52j7wwOKtvf297L+0kWgjnahAnhS71XYxWX6d
lD3Gj6iMsOLR4EGXX31JWKj58ujbdShwUlkhfJOMg5u+y7FJTLBNvSQQ5Dk4RN0y2fJw1UH1dKZe
J4d+3q3U1wfsf0QCPJiPi+lu6sLPXl9PuoVLPENp2TDV4mri8ENXrVOEzyWDUU13X6bCkT2UEDbD
JONBanhkcCxNbZSak/LCoZuzHHvksZOt4q04k253nUkD9qyMVcT6CuEggMnv+14Ppw4qqVd72ef9
fHfo/EMfoobEsEGpziKdaxcFC6NBerQvZO5yNZPt1n7BjEwx29Ds2vC8iOHhjt3iez3Qt7YFHHf4
QPOGgQBMNJBi/YkZW0aYfRR6opbtCqGAkdw+++oa7127PwmPPRm3vBl+DxxHyaX+qAVzQMXFGVDq
Sw8xULZoFoe04N4OVu8JXVqU/mfYkJ+dBsaf2AYOq+GFK5v/e/l/Q5y7/zlcj/KtwTDCEXY90NlG
37JOF6aGvO06Q92JeeU1EVqGctkPngny4J31HYWHucTR4jHsgRdRfzCPON+pR5yxhTtuaqzDdyTb
prkE8r7w3GvfHzSclhAeQWMreHhLbG8RFY7u7uIzjr2r5OP6o4kEFUKBQnVqy3XqeESqozCZuJ3A
G7ObR/7LCa1t62D36RWGb398e7/PtH2m3mPM7Ap/sRdvULd/5wIs7ka1nrhV+4wEXBT3tRm5Frrk
O8BU/U2B5dY5pgb/84xgXTA0ht/OZp36d2ug1i1Pqpm6AzxVxbZ2ZE0+PS+rKUJJIWRdXchZacdy
C0RY6Q4C2P9YLbsI7meO6dhBcvyPQ6WvU4N/bYJp+R8dt/itC2h5W+QKK7hxv4ZraH0AfyUmP+EG
1+OA3Fgp7V3V0i+z5De9DTs6Dw8T5L3zwWCJHBvopyEcABhP0sNppgTWw8FjcwlhiJZUwqR4axXA
2jkpjj6+mEnZMZj4VbUjun5B4gzZ8aMflIcWlzyisAFwT/3nG6DV2RrWKlN7hWDco57LfVI49VUZ
LPlBFbKGhFMg1jNZ87Jp19ljgmeOWUnw8fssSFhyKpLWTKpyIj0tjkk5wxfmNl7ZdxCvCmWf/iR0
Ckn2/j9rSS25Pw7I7yUDxir2ycXsdet+DiOLHK13186OVNnf+bu659ziQHxmqILZy29utyH87B8s
eLS1ixhyruhgTXjreqIfujGeo2L1Yw0u9og1gUV6qyEtlqELQ3soTf0oh2g3EBNE5UQHdm0BqYZy
x7Um4YwOQ0edSbGOIUADXI5ZUGuQzU5GDA1WTdbh35+dFCnQMX+N7KDD4zKGoQU8xK1YFh/zOVTY
m3eS7zJtBYp4qLqRMPwI/dpDpOxG3vqiy8bkqnRdFgVyg4T+5pz6nSivRQHuRyi3K9QhVlbuptN2
+x89xYUVfOE+ghV5MCoEuNU4a9pVNGNnQ3wq56Aau50wAkJUkjH7Hx0XRb6ev0+aOJHrNoMf5B/q
OBG/Rm8S2EzgTxj0Y4frQl9sVgXQCYfjvKodgRW58G5cSIltMHAy5SBhsgmXxQcYPqthahy7DoFA
4HROAi6iejXIpN+482LjU3sG1Q5ekZwYXwgidN32BjAkTx509g1JCkagyC4u6oMeWWblYdkkwEcY
k7iYwFAXwHxO2KGLzuHJJqA95QQqBDIbjWLjK8R7nq9k67wsUxHxL5g9aFfoSugjMimLHGI9X6Q0
9mQVyojiBTifCUBagv2UrW0+gnXs11yGuSLV2vdBh5knAWMKkMQpwwn8kysMMhaMB2R/lWttvy2R
563roemVr5FhC7qAmBkETBqZfcTrnx5G807lvGGxHRrhWOx9JjzgRTIOpp3gMGBG5X2A4GJsgkgc
hTA01O/8wJt6go78jWP9IAkd/yOGZqDaSfGPUZR0yv3gJipTzXKmznQ3P9p7w28OJSZ85gG/JpBw
ojE/Pz6HtjYrSUqVzIkkHQhmWpavrw3Q8VovGjJYe7AKhEbCNcj94nrzf3ZvhYlom5k+z39E+d4F
0IbqH2gu0OkgtJff5HL/ykP5E/RrFGh+aTW+DeI5pGtLWMCWvFvyG0oHjgRbOTHIyVkU8a+NxGar
Ey6hSOrPofH6Lo5aKo6BUvIUrXO/ryb69/zRw9kmBforNc0FmuKCTyYHMfTiHEJUXzpQEa+7L6HC
zNrVXC2rKhycL0ekGEhwGsnIf4WOpkkgjC1Q28J0tV6ovMRTNaJgSXaG5oIDYUt1jH7049E/ya5w
2JSX5DEbbyQIOzldg137EBtI04K9RvQCY4LurC51qKzxqB8Bg6+I43hVBHdnTrFBdfs8DBr6gCtO
WAlzAscED6SktTadKzS9ZDYmQISetWE2fGiMF5VreNIHv6i81x5JTgXvNyd7sRzt8Hvmh4vJ374O
Imh31Ao3edlxRawfKMl0AwKFA53Fmt7MVsv3NKika24lF7ED7E112xkgvbhLxtCzZKEOr9+B1KMO
vLNDBONJiazGXbdNPtGY2Yv0K/bgph99odVKEIh6O3tDNEwChLkS0od9B7gni9Ul4cvUHEMlq2jX
1MqI9EdULkP9YvhxpvovCKPoKY1SxPssfisFiat1Kwkyr3lTOow/XhpJarc5q6DDtvu6jA3Wx2a9
v3o4GVcl0w7qymkXFa/a0m2WoCmyaWT8OcsHUiSSoWQVx4sVN9zJvASxZqvJLjZsvEh60IyoIq4n
vlbNIQ7TZ/gfdK/QJTCSUKACk6lKkj/40Nt6puOWXPzxCtgN/fmcsdolDSCwSVDZy47HdcRuf/WQ
w8jwENhkICnsADhB9eqW54R8D/f1p+3xHAkoSMahTGW94vHsWer6wjy2Td5Set7Mtokh86gDjzcN
tAzrEKmYh1j4aHXBTDFpPrjZgbzXGQaNJUgLYp4fPOKIxR8MFt+qYxAHrP+lg2qXhGQJpKStvG2a
F86Lv9ZFdaDZz/jRXVEAZLQhWWBSBDtqOEpeMKJ03ghxVnyuwVxlS9oPn9Z6cunE1DsTW6M5OYBt
ka/wJu2DeLjU8B4qm4821r983JW4V9fobgy43+25hJKAX8MgasH9uusWez/YbTb4vhHKv5MT7HtX
QoH3Y32JLtONO9BPUnvHotRmNjJPAMu4R1XHWYBCoC+TFtJrlHdpafGjlcZ1s+07klGWWw9KbCER
qLxKDjDyMF4IcqiogYlZMPxveLQr8HxgDAY/oobnrHG8Pg/7InBoAg+x0dJq8XiV3sn4vxAkNkfi
113sjwmUkdiKM4+7q6CTO3jALcRASAHHJp9cxt4oGjIuKz/zCNbO9jm8gLiY0ChcDeG3wrxKPqqk
K0Yk2rQy0aUErlSR3lNcYHVwLLVUmiE4z1ffsr+fsSMtGIPngyuwbX7mrVjR8zNt6JRRGSoS8zbJ
kqAnhOsnv2vcX+UA8vgpbSMuW6IV39qBhwcGwuvAhMZ8Xx+dlyy1Rl7rgS9HjlGF51XVSaHIMfcJ
oh5IH3hqLKV3oRA62Wt0zA3QMeKJmLnXVuDbUuBsjUSLmblLo9gycXRc1E/e9FDDc6kYJCFk9HPI
RWwHIZhMRPBrc1KUdNPxQr2pN30L/ipw/QW6C8Pt7N+EZTR42I5ZchuxPiXOp8aKEFKt3laG25OR
tk4kgNjk21tP0/8E6nsJ84BYbatOOkXjLvQyc72Qkdak0rqkVQiPRfQpqfkxDBm6F+mHsx7XnZh2
zULZjmgYsEdAdWOv2ro69+tg5S+IlUoKX37UWZyjAlE4gL7GOrmNZZir5ZjUh4o4nBh1cjN0Ntuf
QGAKZuA5AKgKQu2x0Xm54GUfVAz1BxZOrhtHnzjDRvH1N4wEX5Fw4jjLLBbsS4z2oAcyp5HJiWJA
f47BbvM/yvGZfrf1cHp2rvtyum6SCNyZqtlMxa2/3coZTnJc9b2KagiXIbAXS6PT3OPlwmtyjb1C
JvB+mjNi1zDm11E0JIE5JurTBaRfruNeLWNZAZGCweknFyiC9YBou0Vqd2SUvoKZBasnh2EcvF+t
DCEFt6om+6eK+7s+2O64K38Xjju6GHnXX0t0cYdl+72weJO1riUvipkTHYIn6gURlcDRklUGHGgD
gtj66DMYafkKtoz937fN5ryPn5R64+6bVL9uJgRstRhG2MjDlEzF0EXHZ/1JBOWPtB308pV7nnfZ
l2UKzIu7DqoyrYaXTGVaYDNP+p4JHGz6R7XUaxJYsAjEaEp0Kh4eLwnN6fEqS14Cjk9KNu1Xnt8o
lEaSxqlIaMO7eGOd2+8MDWv+6Z8DOnJAgmI+QZbAbCnSOxQBQ6NBsWIX+mEdNAs0xXXjCHuCH6wz
nkGb1XxsiocNsKiN6ik3XqnbeJlOe/JpJbFV1IiJ/6IlWLtNjAXRfm9Za6Atkl9R2yRrPxwUp3SV
Kim5cMLyiw6S6WEoDa7ZjkGwsqMi6VrVe9Agn7XQtpEZy9KPud8RTTLaQ6iWeSZ8Yfa2nNb4J8Z7
sWeUDxDG8TaP09JZpSdOfjXFkxc3OLyyo0prCfQ5SmZdPkelAOcpPoykbBBw1RnSLWM0TbW7X/Wq
ppWWHkUDK+tq9M7BsmdJsA8FSyNXQ2pbS+a1z314glrGocJj3MoH6b1NTuu+09e3vIjgKH0bui1K
FMVkgRFWPKuDB3xJL+EBkMJBcW18oYz0f9YA6VPHByngxrA3FSGVNzML0Qj/0KuAv/3/NmMO+uCO
RHi4PVeNi2S82Q+Oa+ZWHKGzdPrwTr2AAtZW6hFjvbIx7ook5n5Kds1R7vD2Wxbc12qxtOow0942
PJ69xQnPBQgth4FFDVszoU5ndJeYTykQOfIGJU1+s6XRidABLoICqeix1mvlxMstqVWNVQfV/7l8
jMf80ReL0bPefzpB0kmzBhWvBkvY36nl9Rh7OIJKMXnIW5yvGFmXkmIubrvlCiVo+1UByn7Tfu68
szOKT9qtmozF160tQFqs+RhG7eGGy0Nd6iTq65F+TH1PG8FVg9zNdcfyfu7n/SXJsSp4V5JlNBKw
fkpp1IstIkfnzF2VCAG0IzJfnJunLdKN59r2+vvXT7CaYGu51SpSN0CL4remFmZj9ZN2VHD7vbfG
RUDNzCZloo6BG1wAyR1ACCGJAcQTGV4+rq6KfHqCM6XrCO6m5olHOguUouXx47h5+MObm0Yj+Coc
HY9rWHXwa4wC3g3mycZxlPW1UXuw3HawZ+MiysWzOi+D6yzN3uRolBFGBHBRFcZh6HFz/ghzMug1
HicJ4rB6fcqowrRgsuxBko4H/4tmfYfPzRgBskxRFGdWKldWd1ea2yNPBtOiYzEvF2GY2Lljh27I
LrL5Wa7Bmpp9zI0J7H5hVt9SgRdsQTSK2QYkPmksEVlwwPH/87Gc/7FJYz9VylcQlxjN43Kc4VpD
FNpSsA5K74Alysf2f7+nlyOEp6D1k9IrelKzMdWtQ6DDUUcma9f2QDgGSa4nCqilJ8M4dInHwyVy
j59RlelYBmWPKMMx2gvLov+ddtd34TusbcWvV40W/gmQw1ps78Uz3KAIDbEu75e7whgS4RqP8sHj
sayDTXrLIwB+9wNVXt/nY+baJ9VrevKrCFDNBvgMlRHxtnX3jkcrEMu5ZtVNqEp098LzO4rmyjYM
q/f9DjI04TqFfuATGp0KozupryGYwjWPyXMJnT763/8gmstjYPYl5j3y2tQdcKEfqW3m0nB7shCn
WOxiiARd7gJYxqHpjTgjv6P6IVOstXJ0DT4+4E19+Dyghs1BOq6A3tHDjhCf4ZtZRHFI0So0hA02
Djl6QdQkEAyyfWYBSC1cXT6Q1aFa8BvRGiZq41INzXkMiff7ARYO+kcpq+xb9lJL7p8n6jteaAz2
ZBSaANTJjiUdZ01PaMN+Y611Zu+DhudUVuZ6vBe3kpWjpPOzGTQXl2WHBgpQ17OM6zc53MdD9xUv
/17LIilxNucj/WSUuq7koy3HFIX/891/nODtFp49yTKPLw8dTxyDbzY1D27oVvBTS3fNbOdBLkpt
zQ++G6yRlTxRgtzI5UxAKb1ZbmeGLdtkBVrWY07SuMsGLw+ic5fGdNAYRoL0JYGy5PQHQvRoyXWm
To1Ah0oUVEDM+Qnnn2jAUcUZjFMpAhrz/XJcsbThYLv+cj1bMu2wuV47fZoEpLEAU2VlqJW10yDl
PqPDwQoW8b0YOFZyEvdkiiL1WxbNBfFqwWBERYrqSuYlB/yZwzrB8ZH7JFUNMlBdCs32EVqtM/Yb
ps4AoYkRk49V3AajUmlcoAdQbHEB3F3WZryXkBEzesseEYf2wq+43C5cIkCqGFleta3SmHAnjV9g
uX11lfi5MLVj3lxnE/Ls7TJkAOm0X6GxAzAUETY0RoDKsj5rghP9cqUgyovdcZmCr1XobDoXSHzK
ZyCGtVLVWKl1btWfhEqK5HXGCZ8j3qBBIhSMiqZAA5tjWuGhW3x3kkSo7a6Si3872mjWgzVgWhfz
M935yp/tl1sC1HjItb7w4ISDfzOsBSw7fsNp9rTHwpcENPTqFD2vqeYN7a1xcAdF1k8QcIosyd09
SWXNsh1MvuoKKXF+aTgYAqJh9OrT7VreGRDS1NS2jI5WTcXOOpfl2YgdTVJyzAYAa2Gs3K6QKTLY
15fhpx5d4rTo/d1+7CYdtWVNwWg1q2oFZTpXMdhV6oXop7niNu0CKAkhak69G1xOQXHkLCQotyoJ
KWvpIISqMbpfy+ApmJLHJl/c5Kp3pW8VO6uLeDKn5zC7O99Ma5WmCajMe5slZ/gdeSrYaw1BxYsC
dw70yWwLbbUM7rRZvoaKk4CUb+5NTUcRLM9H/3n1WZZC3B74s695+msxCAiMeTuFxGffKL4ajO6i
V07Z/jqdTsQFdbJgIri7rtIQ46L4gfBrJwds2v16e/xku/HK6HnGtplQ0Qovq2QDY6q+IKw9eAtE
fSxe+WW36+02y80Pekhf7hiyrXSofkL7jP+2vk3gI+BGqilUzOEpDgHf0s9Y+i5DdodwxLr2imRV
wViuBLaYrRB3fJG1an39YM+oPtR3s8lNFromfX0iBBI9JOLEXnM2PA1GkVQiqT3ClxwQq3derWI+
nvW0lk3AAA6NayedO/oy5XFTvcUtkOdowQ4q8Fg8Jl8RKMAtHRSAyZSFTlxOkzC7FNsSmQcc3OIq
16TBAwVMubXDofvFPCLJHLXzapTjFIK0RED0L98t14CUTtEIKjAQI3WOcIj/RHIZi5UUi3fzG7Vj
bErhTpXym8zPtnCjGuXERxtUK/7b7eNy7hQsoWyloXKpqcM29DLqxmUmBRHcr5P6AK6PxNQy6EAp
XYRqqOvyOeGPP4CPgLTZUnNAzFSAbiejZdGYFU00LLGOQj7cW/xnYe4tq53SfmuNukyOnzUXAmj1
XEDB6t18SAjwQLZ8S1qp+q/sK9akCm/MiSp2yjcn4BtL43d4XU+AA3uvzRMiIqIYeke/9DWmvOGa
l/ScOVIruYhNPXeEY9JfCPIiHF7O8dPUDellbn0xioUl0myinFyGnAfbur1nP5aF+NxwLR+QR6T9
cTBDJEmVbxgQZfv+dVTCbOMK5DKR+ZxNiYy7whAwAnMIy8yq8eBGMYtVC3r8eh3jwhlwIPJCL90I
V7GhSqp7mcPHI1Q8maf25fRJ6R3ZZgutV36P/fg9IKZiy7KFbaL7AL8hQuAhx6sUZvXvMhkB31xq
BbTq4DwcYkR2Vhi1zRooqSvPmK86L+9gTc6zkf5Ka/LF+Y7DTOiAAy3FaeAdyRwyQ24TQvXfn1Lm
W3U4W8Gjpe06ctzmRVa6rSUidYrvzQlr9GzDykAAhPnmqJrkFlxTJY06xMg/0FOdOelV6rlZbla7
yb22srYc2wYhsAbljiKnMhuOxCFwGH7g1Vg3CuR+/unru/XoBhon6qiNJwNez4S5BL+qI8UcOc9D
rliu+7/wpRsGy0Hu1FSG28ObwjCWqT/WND14OoE4nb/hp9ciOCs5vcDTmBQEGUqpt4WRCsvZoP72
nw4lkiVBsB17WAUANE/f2EQD30KkZafv5hSZ2t1y33hBWusf0K8xYWMys3v22zL2+RyZLznfkDJj
BszrJimdZH+nlYvn5Fr+I3z2yMwjvLoUiEBMtFNQX+hUyhlE1FOtpjInU37mbJG/nNoMG+CeBzRk
DW33oUYZnIQ1cyOVeeoIBWPQqX8/r/FSHmiZj7wfKnXwdEBTH8U7+uSE4YesjhqvkyP/zXwrqLr5
e556AddHHv8m2vAXDPcEdy68RU3rcghnrcjyd3mpoa49UXqNq+UK4nTlP5m40N8zwokxEKEGFbeF
WK7WLq6JzG5H/5oJMCnGDYEJn0yKVUjW1WXpJ5ohQJ+PR0YjSaEJj+P029ZaIe1WAO+kfL2xaHxP
kTroQ/lu3676qxDzzKbZRZTiTWO26+1G3k+cHVkFI8xr6T1Fp+u9Pd6TxefNg6rM9Nva5oPlfhPw
mSTsO3481MMhTLqprBagwFKs47qw8o41M/BC4YV3aGRAqqzsDg++8VWVHsDL1m68EIH/V6QiRx91
2HyqBk+Pibi9AAIt+TaoPKooDN4+6gIWGmexGFy+rK1tsWSNzuHTjq2N+Nr4FpvQ9N83qTj/y1/U
FLho8Vy775CzMu0AZpGQhniRq69hKOO8XVGWwAAuor+FWDvre4LKWz/2IkMU9LOFpb9viJurLTvS
+KFQQYvBAV2DNdBiWuLd0MI+pFpwBe796SYH1diRq41Mhc/13eDVa5M1MCPJwSjMGBL6wQdO9+Ah
JFTABTP9WBON9klZ2OZBQ5OknuuQrkNKoOXhhVaHIXS1Xxg3566/D6Kpbo59KlUocoCeBCVxZeQ5
t6LFpjw8Gy4+22kNqUSpUmlclCjbVAM9+fKFcqEXWQubx739CB7+3WcCNdPiSJBfVQbfXbEYAkfj
v9QNJWW/XCYq0vAjSWTjIK4aCoyDaY7uuqIknJOErMhFztUhtQy+NZlIf1mB4p72JXtAc+NDGMDn
xPKxnAVm61vz3YOQALHJPB5yYuuf5tu7vsIfqMk5Q6yaeYKeNm1lWdMpdD3m8AktjqThOZ7oxnA2
4P3IVF86qI+RMehU0nWWwMzFbm7H40CIn2CXgA6srZK27wif9Jz3/w8cSlDegA115CePyKyCjUqV
S16V6j825uJdnq3tW1D9KGNIJr2CFuM8hWTsPqGhwjkL6/nlgQM0h8xj3Ia9LYyaKSqTsiAyfaiK
Bx+LJKdQPKNVoAUhBxKIwHUgU/dqvKw1XdlGydgk/P0AFvHH7VPdHF077t5fEejTGi2Kv3F+uI9i
FQEl1kfZZ6Y868dZ8Lm11DjcgL4ixgXHSIZwfBz4isSfNSRsbAuvzCYXkkX/anCo0JZ6h14OuFMw
ALtbZDjkJpp+OoSyryOK4MbLzTladeUDVwaKXY24+SdIjSXp7qaQNcCnxK9jAWiW8xfIC1R3MN69
To2QMFH5FudLVPJpNo2MM+FOTgjVjxcxQhkL0DWaKCjhG0rCEHNtdkLtETdbAHvoG94lt6PzUxuq
mgmfhdIkeizjbvP3/b9iluGqrp8bDiJSGmkO1DtwgJ/5q+l8fNvE4d2jZpeX+T0nk6f503I5ejoz
pGAmNxiXohEcSrpHYavR9/j+F6MpjRaq4T+SM4RffjmbYJyZylhm61YYnBAyCxK/UvtZcNd3TqKg
Z4CkrSE0gSPcVaZ4JHIVzkI9+zh2PygbD0X0s6DpyoFQoBUxVah+4IIXf/BFbDHxQv4A+DB9YcUa
EdP63lvMR4K51naCZYUHSRsRNZuFMRKx08s6qHFgpB8C/x26UIn5U+cSS7RpRvDHUzGRBKGnlzdb
n5V0Nl1oPz14MPeV55EeKPXHWgUrJ6S2/rJJHzM0mdPnj0voFnWUYeqmPhyg1a2gv0yu9E7AHn1K
gy50Ctig60GZxHS6JmMeqG8UaJuGatSVMrOnaKg21sAZynFfSkMlS18UEpTXcxnKNeCnsiM02vyP
SWnyL76CMiMiWhWRjgfaeLZWSGajUqQ05ay97I4yRsbHubbt7R2vv43ZtwL/ZzRtQ6ztM3aPpytt
djs8Eyi1jdKqzgmBJ/MYXu9P3Cojagr6kyiWmPZP8dfxjSb0gxoDV6xQTDjqp+4UFSKeN1K9YxYb
wK6sSWHi4wwJ3DoNmBvtEkvfjrL56OYg9OBaXJJe3kHdnyN1xubY8JYs2gq73826zImlkQgHkQHK
6KJovF0B4zZJGIHV/9gvxNXAPSJtO0mRVvHQ0Dq1luDbwogw9Y5poiTcvX6ORpt9e5bZOl1yA+GV
DRZ2WCdo8D4x4Uh2kYAPLid5CdI5vzY+1SyZgJSezKYJoMPyUR1nTKrTnk6eIBNcFSOR09gcwW6Y
07vgKXJnwC5zcB0eosZXrMwZXw/0dsmNpYT06NsuG+9bgMq4fIYziqRbEnAl8N6XrpQQZNTu+RQw
DGQFqWZ4Iy3O6UHuIngFTEXNrnEZrjLTpakoVKEzhNtWY/ACa9rSV0l07pMO87WhPauxlYugfZJi
jRpViFVN6OP7qFJ7SaTPH5Uhq2N7JwgkY6i4PqBfe/j4KuoUW7aWi7ISubNxeRLtk8UdggvGC3sw
AKLKP2LLHUeHVM/VqEX7/nLY1wpR24JtuBYDb+NQljsBJaU/K3ZBw2shvNMzmAvA9jRTF/tRaQQ4
/yz/pqfCEC3gxLlqo/jnIPh0zZxu2OO15azNmShuBKB0lKXK7ffgxZv5kc86I/ArIZd9e6CmhTbn
ouQWW3jA9G9/d6bLHud+WAvZQ9P7MWr2YlaselwsvmGWMBziIlYoxK/bgssBV20L6mQxtY1+VZTq
N5C3AJVDEJbLcwv5MA4zHuYmmkB4KUx1ZSwBTvCOot8XQ6iZwDn24w93zco3CQrH3ZIhjNYK7oqt
eCJJq8kv83EKhFbdcRxi5W9MuxxMiA4aBupYwW6Tg2CUb98cKV1TAdopUI2vydwpoZMXAbRc5OX4
g0m3L+o71f+OFQCLnrqSK/+TfzVSRPNoWwcJjDlxVLurzgL5BNOL7Irwx8iHrlB9Gi6uLIj28lFM
ljJ7TXiEwS5z+Kjyxu1X0oZro9J1DfVIfZRP3iE8qEA3tVaZ017HktxE3SkWnfRGuYCiZuEjnga6
KxIw2Fh6BdXH66IgUgL4qZwWwA1ekgg4BQHFmsdZXleOn5Si4AtZ+qUkIgpEBgqE5Rk774fy7LK1
OoEDPUj17tMHRxBF4xNeVcMIwo2QatBAw/s36z40fXMqcXzJEndO2ED9OoFy2zb8MPpOirMpj8fI
qg5GbYP3QFasF8eai4mReUdnqIVhZ3eANABbKikt7czfFYc/nNaizn+yOuHGYX0i8GqEgFrN6l3k
UHbqhYhFiXQrnrKprBrxbK/8Rf0SDem4OKG1eMHH0FPoXjFCNRdkULa+4IjGe0sg6j3TSIKi38dO
dWe1Gx2eQXOnkaBRYTUT9lSVYDFWHvKwh50DMXuEC8nYVVSOf6v6cyDw7++8C2D+RUclDlzo9ebi
IlT5DqsN+5+EEifYprZTIH0Ej+DV2+ne9oCrLq03RKKtfYtiPLN1CSKHn/6w3vVTyl9MacOhpNl6
MeCjyPN3MPN+qPh24m/x1ya2gjMwEHfWuugyiCDG0efkbkdkegjkdfk/5zRlteTuP4emUSQb8jwI
EzTAJ92asbQEQBznte4ps8+WCiisIyoohofTV/ETGTvgOafBzXxEXTKLdrsZ8j7tKhGNrd0v3Lsj
FSAq66UWoHluBrUdn6hSZl0dEf26FpBUePub+oZMqyn6aHqYWSJs87iDGTedVqQc+vBL06he5eYh
/QUotp6XwHBc69oH14UhnA5KiVjRFg+Hj/sJtQXSkl2hET3EbJ4TOTm74v4stLzlrW4hB7mLKDEy
QrJaMTNUw2RDdXHJJYX2QJO9R2tL+RCh00mXA/qt1FIB9Hw3ESAEDywL6KMcMp9gDFM7K88p4A3J
newfQPZGK5Zv7KaHDCIH5jiWuVhiA/N0YeyJ6CXjYF8NOO15GAKIHFZ3a5qLrze/ZVbjjQn0pyFK
KiylemnRDi76j4qgdDq1fxiqTeVBamRqaWj53IKYuJy+gzvSmvvcUGilGMyPmlAw2UXRm1ET5FrH
bxqy/vdlYia3TEDeuZEGs8Lf71GgTKqbputcO2Fn0gHflIm4GGa8T6S+iuVnEuvANCrolyjxrxil
S0BTU6To2NqdaDfLQVSe5qH6TMANaxWsxm37XczPwqw3kZ3kF8G/7f34la5e6N3hRgfxmexHPLIT
1n09jnbPCR87HCVduSniMN66kIm4YlQmpMvoybxlFLiwSx1oAU1a4cRXlfOZSTstailqB538zOdI
5nb22rKI64LlJf3KNPcveX5iNMmkQv4oMSb6Oz4qpHPK6zRtVLSEc3+tq9wYVZD2cdAt1mDDqQK8
s09hEB3WS1wAxhyLDLw53pVzD3Z8/5aNkerkV97SsE8JEkDxV7kzPfx6fdQMSo38COlx0eCQJnad
ybGER17nGUKuhBY9Y3ny0D/LvzYA7g1py1GouUvhDW4HDYnhLFNZNVzdBnxYf68wC4iCrJ45FOek
bghsMCiDEhuOGkKhjCctsF6AWeHmxyCscK0no21JRx+7TN0swH5Y1c28U21P6JdtbkXnRqAGAWUG
McTeEaBmg3cNwa9+z5Oykdo0IaYR5hYlom18Om6js9nBDAT47A9j5fTLbvE1csrqywNolDSudzEv
tpOqerpvfNxd38teEQ50cmx/0d4mhupHZ1irvKjttTpg7u+4Q8zLHbEF3SsnMR/VSpCls7BNknAf
CFHhM64COyoaxDmy7/Txgj4skc8sx5bchvuBVbLdXqjDFOYzRXN3bEO7XgB5mDsmR4bowD2Nx+lp
3hlTfe8yA++t8xoAZHWzJXg/mvtKr/n+PB4VDa1lUSC16HB2u9zdXApRNUZEZBEOG/iO3V/r8Tvd
tFOdZAqvNcU8llS/C7T/heeOAfAFcEdCUKAbMhZ5/lWIH5LdWHzAyQNENKqRqVwnUVved6V/DnIg
3+38MfX/94UBWNoyEr72fEtlmbwsWs/A3lg7xvD1K3CX9eWBIbnysTr94UVa6QP559tJujjHCFY9
PAAzpFx3abKMFGRPf0LcTyBhnu/A/xRs48O3y6AjcCDWfCHtwcMLeAWuXaG06SHoK+2bcxJX9Gue
kbiDJpYCpFQ9YfhDQX8gMcW2T8d1iVkiBMx88Og2QtsX4V//jxHTZcWito/71dTERStRuhcmMYit
sMFuIHW1+ttCDqWqXL2Fc0smjYk2sk+mW70qxcFWURff+CfhIvUjqXkkC6yEIDDEbeoVwkChjv2q
3tGKGXlf7fpnzHpHezNEZPY6/k1ThGx2lIcPkpM48xecFRDSE/ZbsS2cUj6/gVSS9BAWDyI4IqMn
kV3fUh1JIoZpgEQU0xNU0ZEQj2UAtIgKUEtllkd65tVu8mHz0tt1WwfUBGV1ZLFHecUc9VCxihjt
CbBlsr0DsDGYsd0pB0Bmv4D5h9AnPtI1zUTEUPsn1ugahi0kxEGYOtJL15mFN6ILMhR3+N+ri0NQ
SY3iKi4klVrnNcE8F7dvQ3N1Kcs2r9SUHwCVHzoR7LRgZE7v9+cYbixTCwgiTGHeXrKfpJc1H7yU
tpVHaMnVc11/0xwnuOa4ZE0Bkr8pHpP54CvMXoDBfQXB8CyHY/TOCWZnmdj8iwTRiM40jnSEmVGx
roBD2UTlTZYX5UzV0lqz0C8X5uWOzvlRkhyuSz3PUq04Mwc6nyFrY6DHo1FzxiexqXCcEih2zOgC
4MFHiuUv3K5GU2Y4mn/NAh4qXYBhxTvrpkaadbC4mmpIa4Qoh410NJxqFt4jLmFx11wkNpzqgm6X
mgVpYCZI5apR7zGde91pXzVoj3n6+b7b9xUZpntLPirUPNWUecZWcBf6d42qhQmKm/dVPmhO/54h
impKn1HgmvTExsWG5MfFU1g32iLPDrRDsT5G1XrbTrojrNisMzICY+UDLm5mlE6542v+KINiTdna
nV1xyXx3YBBOV9ahgKEnxGm/UUL9yeyRt6efNWpcKBfkeOI65RPNB9p9LxfDg8Naj7fNym8AT0Wc
5N+eX38bXDzqubxbR0HGZ2UJA6nDxwwr/DrxAyeL3QAFwRpBetiR9m2kEnWEzaHdHztXa/IuOtw4
sHg72hIuwUERdEtDoZxsAaDTgzhby3A3FOXzokSQgWh103sklNPgvU9waugEMH+K1mm0y7MAaNhL
qect1f6+eh7qTYwdBKPuPBxF4uoHXwgFilaQmyGY98Y8OqGSCl4klINIqJ4GhenBL0G2yTue04iZ
m4EIDvzOHD7PoaFYjaftclgchd3cji+9xPiTfG0s2l5nz26r6BRcMjai/ZmcYw78u6doTZk/dDAj
4+PNAMqmNWMdz5p9I5H+vpxJsMMEe5adkSo0z9KVPmCxyaAjXZkrq4coRqqJo6DssWL0oLpdFMFU
TSKyP8jnjMK0N4SlgbNFwhvMWo6W6+vKpMXzEaOgOcCTnNnnANQTPjh+QbxkuGN3ZSQ4zhm7VA8q
RvtINYM+4Nm6otoZMsLGomHb5yoFJrR3O5YxafhFkbBd/0OrLGlHpdh+XXcapJ4G6w5FXWn1H6qz
d50GhQPyNf9OzfVxHcKi+T+vsLk5a79gruf3tDyWezRK15d7DQw1PtG//soQrk1+ZW4D7XkIkexc
wgTDPHQ1ag03e7eK0pg+gwuX0q001mJUfLArNWiPCjsK5uSvtTi3wJB8Ir+0Rq6Y+gijClDFJRmU
rCW2X5W9V3G28CVgBiT0qi8mxoBRa03XFSWkM5b4HO6MRqtPLPpzsqPeU6iuATly4MVOpTwqFEwb
MSriHHUx63w8CfqF44bscQ52PifJeH5tXiB6BkM92YS4k7N9T6Sjsn5XahRWZZvUK1sndXB+SDzh
oqVp+TLhAPevcYFz4UuMSMjJmxe/KyMuJ2+YlrQMKZlwizPBSZn3ZujxRkgaDNEa9z45BchbR368
38jcFJwPJj4N6n/iGH+ORZ3uJ1vxKtgI39mSGT3m/G9KtTHHTx2mAa/Say1pC0QbwuqH2Tvq2deW
DMkIlMkOcfwnq2h2zUzo9PZqtsQjNUVeEQMOcdpyYJ3ruyUCrzVhihirob/Eewn7kF/zN6+kTwry
obPpBk9F7JEzK4z00lmL0LWNkDGGgHL2r8MzIEBSdpusa4WZ8vrRgX9FLFAhymV9VQbzh/8oDdbS
mCb1HtfS3gwBSyDVdPrEpxeT+Op3HZREz8fHSRbtkn5mt9ZXjAl6LCuEscq/ShpLcHN0kIxWyU4Q
fw/0kZ2UtgVwPbqSy7jFNE+ydJlB6FQ0SLaH60oURCDwIubgQJqgMEAzk+bdM29HmGEqtahIeGza
ldWxczXssXg9Es6dXjWX86zUp4GGsp4/8fP6lGhbUnxLBEyXXuJC7KOUqiP/I1odxsppmlpOTsR7
ignNr2GohudM3kCu6W0gHsLp+ZpybAvlPzDB0jbmy4Aeeb8V0F3oHu2T4MWkkOkQVClim/EFdzoL
dqDiOD8M7uC8SHCvflSU0fwOpZGmz+988SKMnuQ35yW2zFrF4ZMsB6k8r6apv5looNkJdVWDw+GN
NkEG6f6697QamUG0t54CuwbeMMlmeyF2UI2OvOA0LeSJqrEP0bj03qiIJB/XGgv5nPg35F10XaB4
5BaV/j3vnThck3ZuoATd3J7GX/eBoP+4wmNyxZGHi2/tFm2k7d2P2ukkqZ1h3cEP7OqQV3UBY+pD
+yi4mnKbNykDa7vxp1fvC3ZW3et12JnehrbqxVD4rsef9JmN2U7T9t3XilRBh/Sp3adBogebDRKc
f9Lx02Nehm2a1tWxcZcVhvQHTHO3G7JTyG8LV86OfP9EZbre5wZ2PK32yCpdF0zS3llZXO2RNhY8
b4YIiuZ4X+egK87/oWh9tCWzXXSOJfWL3lrh25N69nw2Lj36JuVJ+2Ij/6+vHYtcaDze8b3DQ755
qp9Ggwrmyx7OoWarmtP6gsbruVGm/DKdkwqx0dYc5pPbwiWuNFAE80acQZWs/Zjbf80IQNKdz+E2
C4V+06Io8WaI+NmS5EmoSZcJOzeDpt/086ul/lQYXd1oeYqu4PgDCoFL6DgG3kzpj0LOz8rgj41x
kmsVgBnn/pv8bO1ZyTTajKSGGzkMaIxdrJ+dvjI5GFKNDkoccy0bg1J/sNtR8Vg6lSbFGSMwFrE9
7XC/ZfPZBVSFPiYDt1ZtYxBPMsLkFinfRKQMQWk7sPEezv2hA2X1pckBb+t3lqafUJWlMBCjWGMr
YyTl4fEIE3UovDv4a40NRffRY7HTMtzMpnfqWE854r/ZGsGeoFqHGB2c8IMhv5RhaRn5CCs/HISR
TJbMzx9GjOhfrgcHYosyBpW36bbscbnVYoMgm6gTDBR0mb+cUG8wyaTRHOHxaqy/f8R45gLutZ9X
9fQZUsXDeSTxJZHfh3Xzocvew7iMhG7r68TLx3F5Baf5F2yaApSaazMs67bS4Dk/s7xAaa36b+VJ
wO+TO0dLKkZRDn8kvyqUQ9vrpjTpERpmPA6T6Q/lwT0sngkOtidTdBW3eK5NR+0/QJ4wqGRQM6ko
vGqu36LmVKj9stf1Rcq1822YfxILE+yueLlm+zKGmZTpWRZe3O+j/JT7injHLI1zfvVFOUjQNLhP
7o3VmKqQVTwDslRJ9pwB0HHEPr4DCtAnBtU51xiiPQVoRBF1WSAZ+fQ/vjhMo2dHU3CphB7BqsTK
v3oDEGxwx4HRlUgD195sQPNF/qecsFM3xzAg3dXt7ue0k3NYfbBmMBJDGMfLuxcaYcQ4UvCTjire
DwtUjk827vcoRhYC37WxF5elXo9E4a7cyQ3DwmTf9VcQlC4zk7XIqhUxONDp0i4KcKK4xVvsPOOp
MW3SRKPgqbquPA2OKz4d9XTrGepTCfEL4h9owuBr8OlGaiSa6CEirhr4Nz5KugbRxreh92tLa8Uw
Or+U8q4OJ8POJD1rAxcf9WPeNv9oZ+H63mXEq6xPyXfhuIQslySPMde9PfS3bcITXYn5sOjFTbAm
NKJgjGHdoFMc/X1gduC6zZSKYNp4BGgNlOzU6OOxWyBbHTS2gCy0WHn4jzWD/6BQuxd4HqGcdSO7
EpeEy5oLfTlIy9JNrUCSZQ7uBGG9v2aoaaaoqktks8zv5jkrRCgl14s0GUGOw+n8FjomvRziscWq
CU8eUAG8J2sF9CT6YSBd0K2FnjqfwCI65i7IXkLd/iXFMAcFZPoq10Qp0x0WXdk7BnIsVX6vHXRV
PZH/rjNnYVedMhsO65QVxoIeBOEMsCJO7FE7898S/OWlELCHjHTg3ODlolNWRkgTu5nW6LIxz1FF
W3DdiQKvTS3kiOFCF7UHZS7IM+eE5a5WDOgLX8VsSQ7caXgQFWTOSiWoEXvXSnV7/zwsgwLPTsve
0zR/L6x4m19aGqG8yu2S8ZvL/Wj7zjl9nAuy7kGkdhpQCWObxv72Dc0IwBIymHqxSHi+WBb0w01c
asWlKMEwZhefSqmxXjY+LYyRaOGe5PlKropedcx7vks7rWeOWtAEchEi4HLnlpGuQ0CgOimQJfEK
p4yXO1VzarJpVgxjRNoT8sxL9aY46muluAHe6iAMKwG+Mdj8LMzklluBrNtB+3paqXCXMmn96J5F
O1S1ifjnCA8hEP5mY8dYfUY8Gt6mJZ8z3Bytsjq3BzM5EKaKwezXrtXzOkbZ8PYCDCubD+obVu3Z
ayEiJwj9UUiNBAdbwkFOwsCYDmGivPrQLoJwQhnbFOPQzkF3NUah4YCA+BqTTNBSPigLhLU2hlQD
/6FrLgQeTAYL5mBHbNDTDpGZ/4pyn7J8ustrnZY+KabB1CCPQk5X1vK5NCb7ekxps8h7gaKPNt0S
wtiWfCSddTqKA2lQzoai9e/l0v/GfUsqqHtz3eiU6BLe/LHDVJOLdts5J00n2xHSpss8KKu84yO3
9VhQ1PV46hSMttRZ0AMDvZdJB+XycjMmd5mb2tjq3mRlFPV8Y4DQDoEOCHVltyZ7G+gvmiZZqv2P
YsuQ4yVofun6PuSX3ai2yCYBSyTBszIlzlS3gK2EhVf4EfFx69d1e/Y5MfQhd4CuFUaXbMdg4we6
F4iW9i3ga5UvxY0A9vZtargh9M4qyd4RhIsPrOxgHQ/2kvBhFAFu7D9as67TjwZ63/OS8wDLZDjW
xoZktGWaJpwUXiggSnOF/efym4mLFvjbOLx4QWoq+85mVV5zb7z+R6SNZ0xxsxeaTNVK3dC4brxn
XVj/m7ReH1nZOAAPEaroyit+ofjFLexGbdLrizwHifseMeeE7ehskrK5pVamvGE+EBDN4u48jz6J
GYPO/BqdtZZEumANutYbUrNGM+oP+y3DjK+52Rydo4k41PMuddkHeIJPpGJryvaH+3fS3y+eKzx9
mY3PqYwIgDi/KJYxCxsuNiFyAQwTsXHa+mMBuS+lMuFMOTdhiZ1FV/pgO1P8i9GDOBLmSO1qDxrY
CZU12P6l+Ov6mv+FnlNS9iW1ckZg3pTn+ogydbESZwbv795VIgOSvgCd55rP5O85oXjJPf1p6RiV
MBz4MWoa9mq0IK0YbBX2sdXN8K4GX/jsSBz6EPNKaUNPWxOEJHRd7v+e4Ke0h7AKv6eHhDSesfKa
9HlJQx6FFKAE8E03iA5IfeQG7JICfphzIpsTlHr131IADdhO3bKJtQrTXEdAPWXQOiBnFdikD3Ru
ZCOONS1rIX07739nLk9engqMSjoMWhJtFHIexNSyo8bShfVBlPhkL4e6jOnqoTTMQOew9dwcylTj
aE7NGv2UmMJPjdHOgNIl3j6wCHEKhb3L0z1t6MBalC2f6rXXtZCNetwZwK0DX5yfui7fjPcv20Yk
KWSBbA2DwUl59JTSozlpklb97ll6xbqXKRmKjh8wOJv6EyTIpunF5Ighm6FwEaCb80+8aaEG7dkl
/Q03ZZLKR0Fd+cqbSXbYlRhTc0aag99TshPcA50lucOZY4TOF7jIb/DK080n/dhTnclB9WnkCuVK
rNP310NRgNsyyV5mcLm6Y1zPaizZ2q+d/lKy8mpcWNVZm4H97rmtGxQqjPz0RBtykaoSp4mOqvVj
bslaVkPPJzApHymFhkqTNF9Ur2TGZ+tWap/aANH894W6LOmNqCcg+kZDW3bva32yVNoiam/6UOWy
hjy7O0eg3LK4quo1FS/oA5MJAgzRs80s5nx+7jB1VEfs6HOj98b7pa3E8G8bwguq+DM15mDIwL87
D83NeIwQrFdU6qrxFcErkx5UK6tkEDa6kt65EY+iQAseVga1XaBBbXj4NVzldddCTrjAFaxk9SQg
NPtGnRMESjotzEQ2P4FsB21onE0sXXVwlNJkuYFpgU0kyjQw0HQz5exkA1a/Ft8SWHsWLRgEj8B4
bmiPZ54cUfOV19eTYumZ4LTlegrPfsB8ATLP66PzVjZ0A/xb82IlrOEtIL+ml2W+QBCCTVu4Ru0Z
0qDHmGWsKwGxKL71S7gjGGbibGQTXYUGrUZnbdR3oKQfqyRXIcylpJ7L0E5A1DQ7hxclLNwZfLcb
Aao7sCxyxQnSBl4usgMHiY806jeTX12nrK3jIY5xTid4CmLfb/35q20n9TgmHe1ZwCYOtuK8GjYR
JgEk8SKlxwvMUpO0/RClAwVMTVNNduFz+qV7upW0FHYrlCbPxQuZbr71EiidOS0qTkiiS0HbhOaY
31yWgV8VvFWJG1Dua/MKHfwqvLyUcYuvMedNMmiR0w0UxtHP5LcEcIWaOj5OaFMRaSchFX9GU74w
0Zh6JXOux+RdU3xop/PRcI9LjDIwqejshEGntRnX4Oo1lcu0rQMCSGGU/7SCWoIavMZWWruhTfmN
I5pLViN8lhOuUVTpn1fa0wSPyQFaOaoq02rBFX/yP29OGMFNoA4txTaG9UtHsighSsOAjJ6k/vws
Il/F1sdBdgzCjMnPzuscSgPOTdF2YG4Y678/bObg44AgHlLP01IR+V555Hl5fytcUWF7xr8r4kB8
Ga2zq5Bp45msCakcpiTkqRLFxMydOMyvEzPDAcO3upzo/8ZSBqbtdD6jZrJQXGq3bfYWCg+F0JXB
BY0SBth+2Ec88HIW4UybfdhTlK2AgvNZ0urMN0dqIvzJGzxbzUg27VGKXC0gIInDD12PIqTO7kXR
eFWT0wo3AQ/U4jbTN0pQ0DFnmHiuPpvpCUBCIPr3R6MWEXD5N7T9n1NcIR4TQoAo6qntwhrOCZhP
CpM53po7/E8VjR8MJdcDRx6l2bhk1H4nlxlSDdIHHzorSyb+fWg/i+9d5VFVRIp0n0Pr07KCnEJ3
u4nO4H/gaJqNVyDSB7l/3k4xKyzCMUyLy12Z6IM0iaSVutSXhGprfw37br8l8MOmv9TNC9vrDNHu
L+YMqTcvcl2wOhfqEY9i7HXzQMWIQp6fDMv6lXq7qlOJvMnEIdF8MdhutesTBewuK3F9dtxCJv+e
DDTnqbNx6V5iTda7adJneQ6G3bbzLL4q/cJHdh6a1ptlwq9YHo71n4jL5ic3eEMsbZvQ2g6ur5My
gyTCGbqtQDXXZyTIlTMJ1toQ0Z1cb1onn5XGK7xiisWSO4LuLQ4l3QDWJFVi2E6CTJbmvHu/+KK9
dZ5cL1L5bVCdxyeOeOj1No/humQXJoz8H+l7DvmTFXaYkbw29xMypIpDrZfrS8RvYKxn4aa5Es/8
M0UZiw88P7FB07iFBmHPu3Jv+WQMuGSTV+1LOT+hMA1zhWK6yR5DFJJdX+c7sy+Wo6HzkY0LPG6K
GSmtQVBNiRS2eVr8rP9dBn0kaTkEA0nSyKDR0fEqONmQWZhHEmpDUW668YmGRstMZiBlN1PQ2m5y
faXaQq4rwAZ8glThPRQ3Mv6UMdyQcylP83N7XYKuzWPhVGiKDPEZWMTX9v/s1XsvEEHrnlyPX9fI
SyxtPtSqCGLqZKm6OpL9s3doC6BJP38NCGCcrQ3rln71E8zg9WLJ6h/pOpECjqWroY24eR5e/NEu
a5/U+2xO4+XhZIkXjFwSfGJQ+0mbPZjKHjtKE9fUZ8v06z4HgEqxW06keJsZjI04OwXdoCbzocsX
eib6TSGLXVEW++gyxX33wSE+sravk8oxhJ3FPwjqVyJMjMtZERnUlpL+z+gbQD458NgD5WseIVwN
rOzuisgUelTt1j9I/XqnLREt23z6ywIkbwcQogVyDVWnbv9/ZTvbmB2xN7d/EHOZPeOcO8IPJFEe
yhPDJNqh4Vt8P9ZdH2NmKHz0rRU/e14YvWyMxoRwmPaHxdnW6YSJsVn/l8MXdDPhnMbpO52XoANO
bamH894I7j4EzY0Wh9qbbyHxS+9jvqgJtvLWprnNxvMAlWy9K45tncG7Z2DgxNyr7Wr7zLvR0wA+
7Cw9hKzMcuoKh5SvxcElYPQOkjKA5U2KMzhwOhZUiOi0tKdE5g1mIdaTVpGDf8BkHzJZnLtUtkeN
NzI6N8tYuU4dseq5kx6Jt5vyPoANuLa/eo8KLrYc9QxWGNRW1KT0FC1RW1rZiqv6mNPypjc39hG5
OR9h8QpHYX2Tiuebupe1PZe/fyWGBLIBU1B/7q183nTxtU8FcLSJTe9gMwesOSm8hsnTcMXy55bs
eciDqR+QwwFzxK7hJbkPQ3fMmMXXC5E/9fOWQOHpxEYkbWbXiZBK24j5ElpPeV9DV17yZ0L0boum
/pPMYN41CzYjiI8xqCa9xXm9AmNmlLr/Ee/gHhRgR29P3RetRaIC+k8aQdJIl1JbfyM0HRRkUTCe
HkJ5nmaFGIBvk8wFc/v7xkX2EB/4p5ETy0HVzLu3XHoXIF9DKN4A3pY8wVoaYUA8LyhEqs2sUL3w
2+3uEVIC9VRX86ut1QOUqcm5vfzrmwENvbPhsRKhi/W7iTZmU7D34a9DmgC3J/X6ejX0BDf8eU64
KrFZOzwkZckAfet71ckfNWioP+cx/9oHI1mAGTXzTLriwrA/A/D4qbbzX9EHhVSUnEJfYuFBkow+
fSsFHHYsTnGBtm7OjKskmhUUuqk0Gap7ujFAEFc35612WteyoQHusvkDLXXtwpEWo2hJ+I9URXcD
tEc2WlvKiVTN9ciMcxRH5i4bzEMBmlI6pJtMqZlFKqZL3mSTvyfnnqJ4tLl4jT8o3HLFsWqv7Pvb
atyHinp9WdZ2vzFtk9moKU+aTQlhhTd1APSBZuLAFNkU0zqaMjGsxkrnOqOfv0xpDVOLO6vGcKpx
4mtilu54qFLmjoLUnIUuhoYn8sZPkF9KE9jYYz5A2jH9tan+9TnMKRF9qx8Zjn6EjPRmGgdteKe9
uMDsUJkzneDrY0WEWT2c4KVoKYpYN1DQ77kxbboXXCeWoeVgTrr2ROwuVZB8sufcpK1JkbJi36ZH
XWmv6DO2t9P3kbBONsM1x/KK7ge1RlhHixbdcchtfsJmyD4S40Q4nCqXQbeNYYGGi2s/PDbjZx3P
kBM6zH4Fh5Vgs/xZOzWNosW3rYYv5a2m+oJEdns2+SqSuHrc2y/nUp3VNtfS+XvqPb5OQZOWqSyJ
c7W4pxAUYa3LMuZmaPrNYJVq5s+Qn56eprP0iP0+dNcwxZ+lQCCPkThK56EaWerLJQf13ipn8UNW
QXMlsY8vvxIzJlNRHgPhb3KLJfjCfwmGQqQmE9wae4NRNi+60bIbe6ama+kR0x2W7eLbGp3SPDCj
OKnqbEHwfBpSuN+U2cL9EVccPWUvBVB8zYV5FF1HI+SxdvjlpYwQ8Qm1L8mN20C8+EhfPvmZwhZm
7Va/ZF6g+cbBgCkoMWkXHmA/MqKnXl4h4yQCvYlkMvYcX3qXcM8q1wAZ6hHOg8X9nFPZKasdb4zs
PGW91tZ0DCCjCJVRNUE1ttmpbsvN840umzIR0XwmAaBmgesKCeuX+M7r8Y94q8KnmJ99Fuqu5oa7
kwyV7awVFMAdWX77mC4Vge5c7sThScrV4NOLHw8YLxq8rVkkjeBgPObFw1Ob01hpXeCVOONrP/dE
9EsYmHaJF60c0rL0znQDNueeCBXDHI2sdmZuJQBXg8e5wJhCCE10HTeiRcSvQ3+nPk7slqrLgjGw
xrdT6q8cTnmKd3r6AllK6QuK3mbFUokmb7vF65WAn3JF6bpetFgKk6sdeH4WOpexMFqPvS/w6dO4
KaQEw0fwsxMT4eqA+RnoQzFK2LcUKtFHX0tugtT1rrSDZh+9zG3nawZ9KIeRfM4N6Cyt3C1KGmAz
KGlACp13PsKVCqAw4AkCjE8Ww+9CA9OpRZBofCpA9PQqtvMqU4h7oRhrftBzhQXa9WW1saczGjD9
O4tXwCgWToWhQIVsBgmTMwh+CqjygEx+3A5IQjGZv3fddkvQmbAejySqeX3NSAgLpirX/dvdpOZ4
HCSlkbNDlSQpv+B0JP1emcvtQ7x9xJZLX/grE4DuJH6G4+3JdABktEDtg95wC2LmJ57bo1Mib6Kj
prrCXSbiJ8KEgZ+Vu+NVXxQycGhKkSdaQf45o5WBcm+RXfc9TX7Cxu4sBEz5LxwyaoFmCv1uYHMa
uqYfjcvm79j0ClQJ+9qrLfBgo7eulue7IU1HGJRpsUjg31tmNRw9XuocJa1FjCatahS6Kkd7AV5w
n7KTPqXe88oC2SC2Kqxh0FUshPJIdjipomY8TMYqMzFmAckTOpfhLa5j9WA2qUJGcFbmz10ncTl7
jxqXKZSio3SU1uUpE69CLDTDYlP5VJd/9YsOJdNCTC3m2MkR4qm6mT5JLnl32BvN6OfiV4VKcYwC
0yu2C3yJc0b/71bIsgMsNMA8jiN/9Um11SaZiv9jbRJYsDFPRlFDOs0gcTlln4T20/KvdwGdFX42
SELhv3kNdZOQ5NBqgeLflALAQf57N4vyFT6rNutQBKOmHtQvjOBAPhGm4zsi3ia4FaOx8KkHOkxP
/a3ADH9jY6BTSAg6Nk8TSfb+JvuVhA5jZt5aX73CxmotqfCoV8cAoavmiVLv8+X6ZYzi7MY2Cxga
Tf0ZiQ8lBDIk4yH/P3A8OSSAzihRtadUhRIjS9oajEILQ9G4RIpqAMeQqFHfHb4RPsuAi6tGhelk
YB4dbPLWMI/6j8p/W42laY5e4ooYZWR29E3DdUYcr1qzmhTQ8ghO3cLRm7FQ/PN4n56Xk/HP0YU2
toJZy6vm+itNYQ2/yVu5gnqfSGcjtSmoWLHbVG03BkK/8B7oJ3e27WKmXinL3FElGQS+t7DIB2CG
/LmuisI8SCVULAm/515tVuils9SJDKfJ2YcBySW2v079LRWSEFF8oIMpZUpBDeko4gpqqMTHdjXJ
FjQfSiuTRQOyWIL0cI26tpYLFZQA334Itn8HjCEtUSxVEex1CCMwf8p/jQKGtXARGkP6Ewn1A5Ou
MQPpNhN8SY6FMJqgK/FUOBoWlavNIiLV01Le5XP1bQCHnnC/tIse3b1pbnv6NbQE+lxPOHgcKa67
3H1YvjnCi/0KclXrYFSC0TokwQbv3q0eunIJOmnOylzzp4qEjZ+y6aImf3QGsw3rcQY0HsRbATss
KqD5+ntJGEmOaP6Y13SoGfTe8y4tO0NsIhxYT+4Q84sGA958fIFt8EhQiqLek8JwsQh7+5cMtNub
oe+b3lNA2JLtdvrLI+8KD2AfSYXDnUicRE/0ryW8iDDP6QFtze9I0Ke+uICTTGj0MYZwMq3vJmaQ
e4n5qjeDuEH9CUaDaX2PXsdZW+ADvuz9OI5BtBwQnAJJdpsTe1UZAUU5id/euXGKaAY4TyXceoKK
O28L0v/c0wecwPQmpI6xU8IyDasVuJbhIlQ3tPsGzAgFyM/9F0lVF7UabjBmTZJ6H5kaTvdivfLw
1WqB+UjWRJKgRkHX5GoVoj/zoa/N9fs43IeibDndaJk8hU3Uflsa6ZXPQHVkkJldoTDT0A/3Yzbr
DzYpMn3yzo3HJQHhl4O1VvBjliE5RLKoBsbHVQlikVxf+xjYRXSzST3/9ZtnXXWqcsP6yoeooHw8
+gBUdXSqSyf5wCsi2refn8szIl4i7R9a//gA48AYH2PW8dq6jUmT6Zfq8K4gLs1U4Six65jPdOrx
pjBIwncgdIHxGmCjoBI7/nGTNaWcWW51j66WR9lixL2ezASspQ5r6dArMttT68HgwciBSXECNmVx
+HtBNHBMIOxtvXXgBt115utgWw4ScF8G3XoAsgZIvPboFW4P8BhPYCJPpzO4I5toTZTyvWsLMdqL
2+A5xJlPN7plNewLliXV7x+u3FOcrNHaO+yNcaAn4s/tU3ORns+8xzIo/7PieUU4XDi+EJM76p/u
W219uA0ledwmWPFcXNrEoVJqVo9xvX9Koh2WOHcZud6Kl8llgtpWqW1VbaEeTVFgxvEh8uK5ruQE
dhsWQY50isyUpljzLz1NUP8ajHhIqy99OgXN/JBGkoKYOK5rZJIVyvhDBjtD0MyVjWDRqdj85o+t
zFqipjCsuxXIjnIT1zbD15uRLYZQYtHd5QCQ+uo2htrQTd7WsHI6IbKvS/Y7YMh0JDrYp/bFiUPq
S5P8zRTSdpZHpCDABI6DLyNrDvX34AsymlpFTMYxVsYWUxuad92KSy75/31q9sMwoEV/Lj4inRNv
sjartibvM9AQ0rCaxJT9BQ+q5k740JO5EQ28NHWgfOE80R5vx7SH39kzWIBhL2jAgW/duVtH6h+o
hHgOfMSUaZBrcq1CXIpCsjxceVQPyKJw0r5Hms31A6iDH1Q8tn2ovGkOOw53MMys5HnlceuhHFqj
NxccJyvSLdAjrd+bgzky4UF9wwLSfcKIhXiH/MrB9AODSO90s32Z/wSDHJn7JN0TLxcMNDKeEOuK
TLmOt0R5Hv0yFdIebDXEZHNSuFgdH4deVY94hbv5XXMeZxtMXdF3ktCsCYYjeJEOAReMxTSqm2O+
k+AMypUYZne6VCyOGofAjaMcYN1gHt8YywXEjrW2+QlGSVVBpAeXBTDRYuRErI+IU8DiqSveV7tv
OCeJR2HDFcNR+DjxBI2xlXfyMyZH/oisYzQyOk++d64ZHkf5grVxroFSybi9fQ56dAkHR7wSjs8C
gjGtfGKieHYCmDwEGSulrbq1kV2SUqxf83l3/awFzpza16m7WS87pDcB1kbIgbvs9ZyLMObePIF1
ErTuPZn2Ib8aJkypdzemF5RzTYGDRL1KFx/4IWQivM79dpPKJSVDM2jnvjX4F4aCkSw0P8AiQKf7
P1A1v0LdZxfv7c9O3OCvN9M3ANludQNDiEEG2Kcn3Kea7aNEaTCO8sz47mAyfiL4gN7XVFEE54ZL
9TIQfFo2rHCKPj8Kj9fKB57xUQsDdaOqumHUYAfzvm7Lstvpuw0nq0GeAmFV3mHcA1+CEx/MEfUA
CwfsxCbDuG6jtIVQVORQJ3b6FYGok+pUChNkUPaz6qj8UqBJDVAxHsQpPdLMo+5bejMnbqMza3Hk
x4b78I2brBcUKXLJcpk4Q24WM+nKbseSkT6wgNHq3K4RmTTFKN+5SPkRMsitdE3E9duPFvXLzGRt
W6m6LBWjPI1RR/nZ3yIORuLYsw/LzLE52aPMfXUtZnfYDMtDa3ogdlr2iuZUXTJbftvQXFy4hUro
4sY0OLnRrziInCDYzacmgeNAETEctE39r8sS7EJNdEC5MzKsNlQCFcIWvsCRQfIjlmf+CgEjty1i
8dnRU71bCB4Rr5mFGgVkKxv9Aq3L255XKC30gG+R6qCRhz12Gl5iigrh6XCKBAQZxupVs2aCQr19
/ISDRyRwSf7l4eva3W/UzDiKw58/zw3+j3OkRHuPvyYJ8HA2ABCzPcr/HGmkBm/9cMI2AlMv2Hb1
e7VwI3zMuVMsiAZukuH1KyUFTpLHwycwVqwGesBw/AtCOeFLd+2H+osze2syWRMLJbZxcXCV+FMq
KecieiKpob4YfgmqsOiNsII7KZLtjAAJl4L5LPNKimbAe+jJBsbbPPoA2/+7Mcx3/n9EBnO2NsEp
tHBCk3GF2hETL/MGvfIwPQYfJu2985KR8GZm26ZzoIqF76nJh4y/duG8syO+Sa3Nynkt84qt0vcQ
Bnk4rzQ/2b0lS2vrpU9N+dSAlZWGbf8EgYNcw+fmEgElYUJhNy1Fk3z9k0yPIlXdP9V9xUjLoAUW
4jm+x+vIyIc/+rSq/9p6GoaorgiJJ8L9HUx1D1773SSkOim9p7xYmMrXpAFTy5CrR4ZcnolRdmVK
NpaQfZZcmrgVz7W1YYT8ann14eF1XRs423Yl3BEMtkYqZsDOjjLj5lhnRqz4V19K5ZdPKZpyFzF+
8okEJwuihhoigaKQWzNVik4k9ceshEuYUk3gjCCx/AtZrCrC7m8tqWS9osHw3LlXkMRUQvCZfhD/
ZLFC+y2PDJpeb2dQx+BT5wKqIp09Hg7L+XpSKT9+DXuT/mShL1hFXwKDMz3L0grxdURIR0EgsQQC
BqcMaGpYlX5tOpG+gM6MyXkrMazBtMSCZ6dQBOhWHpplDSRlb9natjS8s0r39xCA+PhYJvPv0pYN
2AuyYw+0+/k8PNiWZskn2tf7uGKAkpVmuL4pwAk1xwPkPeI8yz/uoNSiSmrLR913UUepwGOG5nPW
autQ7VBrFDYx+dV2WMUHlTAoCUccWa1Iov60hM5fcuOvpSXELjJM9aLN7g6042aJfy1otEH2Ss81
kGxwjHHv+uE2kgun8pnWjB4u4OTWaNb37Xdgf4SffdvasiwN7PDeDatNapZd+hlMfS8RvesJNRub
NIramh3mK7jP/wfAivW+5KLctuChuWgKgru8aDQzJjXrUkD628T8a/T7PuPZvqX/F77Ry6e5SmBe
MfgxLyYzu6SEuo2y1+9sXz5aaPIyUTRb/dm0AQ9X3Q12VlHiIBwQY/hlIxyuRfPC9W466OQWKHiz
shEIYN2kNwS45E8TXWXirrU1PVOTdJTC5qHglc+aVjrBwGJn/apBbGtaikXDl25qqKt/o+RRAjCf
VaKNpItgutN6bh7UfTy84jFzEUKFaRMVHeT8PzgpEM3ohXNNPNNT4kMiQj2ASGdg9r5GOxf514Z2
rsAyFE9QlmQrWo76NsoqTT9AJukq9TMLKDyExgN0L/lc60xiC4mPWw0P54pgnsJU0KY1Mol0RBbr
wRLVIPfPEvoKGUJVFE013USbU4lM4bI/7WaHipHI20J+xj1DNdTysuHUks8/ARKJT/EaciqOI9GG
telPLSzKqcs0Xunlr59a+pVzvbbREfStUUc63mFvzH1k7BkIjjo6d79rgOf7tF0BBoQ92huKDiDy
pCIad62knvtEQvIKhsbvAqHBamL0gZJ421kz8OGlazdNVr2MHSp1ow5LKkE5davxqA3uiqmUDqxb
Q75CR10Ff8YCHGqywAMw24M7W72dbU+oqdG4gcFBslwZylZjX3r+K47EdNgAiPEMOTZA2Gil6Xye
y/zVUmfRH9F1Prp3oJ9Or0qWlJVT//X1M6FNJ2zpz1vHBC9bTfHxQgOKDXifxK8iOlahkKEwB7cK
q6llVIDX7Gf2mA2Gd+S64CTnVPV7jnNdXGlKC29JghIrD6lUchm4IT105gm056hu36YF+SHc6pjy
iv0x3nsec0S/wBV7MDpGKbrWh2DXo8yXqCGO2l87+qOx6CNxmJ9k3Vl260xtwt5kUIahXM2Rv02z
0ornCd/L3P+sfZaclT1Zv+zohPvLOOGjH3QIxvULHTNUvVcdyB+533uW2NV1/iVebogVZUFFY9Z3
KEoKCZ/EIAXyhUOnzhYm7QqZK9ZOKaAT+ivNgSdb/AZ0Kx4RsJRmjKtH9LGsxr0AJdLlyAJDPcx6
ypinHqwhWcIT4DKQ5t/Emp7p3iv+oag/Zu/KhpxAul5yogpYD/qzsEAU0NNKp/flsXyIvGMIlY2L
rg7gJFUHv97Xc1wkiAtc/28nrGgwhzuGxgEIdr+CCh1vz1oNrM0iX5mbbFEfN4ICtgKfPxMOMFG+
ril367jb7KJ1/xNt4CU+oib1X6CQe6O6UT9KWhHU4jkSoSU3ibCx/lNZypFF8UErdrwKSUJQvG7Y
r2ERgpxCts142gfkGxe/sby+99bKM4dhQYtlTBYudQZ4bQVvpVL80Dk1nj4cGJGNukenZ5omcMgY
DI8pf+GClt841g9t6poXd0c/XveO/empawPeEYVI7qGCOK52RO0AnmKMpaVm37ZjQi6BZJGml1cq
lpSQ9xadtb8iWVdKlhiS4IXrhrr76k1km/J3byY14KGop5Gw8QDVtdxDbE4C7jXN7drhYG7Uvxc5
z4lS6E6niRy3fiICDtaBy9eWcQTnXe/MpfSUJy58NJCG44EShkJJii1S3k1yqsUeHfn4LfI75Agb
XqO31A3vAz6A+ggdiorGg6LCcutGpM1bJuGMQsZWLww6aOiqrPWQsRKBsRlaciVARXs46eLfQcbh
DmCwKPOg+pkDWfnsFFzIGzEUDo+87xMsWxjTTW+kD2BlfnIzbY8LNpE/1hPG8mXQnHHWhQxKmEG/
7XnYXvEVthmtec2TNkrZFMah8+a9z5k7OATgfnLlu8hsWYrnBcI4bU2JsRW4n+T8UCXtjOGTjTo8
LGPAjF8Al79rlkMAvPrU4NR4x+GWA4iEdkk2l1EMNLwI7evEpvjDy7x3vkJO91TowrHLTDaS+z/8
q6mxwB2tqF7XFkE/bQ5ExVeaneqLHzugJG7Lz31w66HLRMBqU0ScyS3rNuSaA8tky42EZEm6JAhP
Q90nIcgYZSlyGO0DwCZIWKpcjVxc969YkHkjuZRwNnUEr1fkEpbYSZL0Yu55P9L3P1bo/h2LPRqt
EXeKsqN9KXXTvejowJaWHTPqx3z3PWI9QZgDWtT0byysCxNwt/mw2NwqsOjPm03XfH0ytjqmS+S7
mXjo4OOCQ/naocJuPuKBvGmSUPYD1pYAERiQur1TquaoPfzAE3/fyK5kEJCZ13ylhlwikRptcyiP
Zu6JX8x0IYsa3a4B4Gw7uLvi6YEfgGqTNuz+nJI8a/VcG3iSWTQieQnANgPCFUQZzGEdtWEO1oxF
rRLADUFAy4kfogL7bzG04uM3CvEF8xA4E7FvpX0LEKRHQaZBZsnsYFpryxDPoRVUldGQkJh5kaWh
xZ2tRfNeqC6Yl6n28ZdguNns/eWzSVt1g762EP3a/1hUBu0uj6F39YQpfWsDycTg7YSv/VziTSQu
pFQntnY4c3TOumJUvkbf/0RF3XRz04GYcarC3nzFkFtNfVMKI2tREjyiWp0OV1PzZOdtbofRm7vk
t+Nil7AA7w9ih6WDvZZUjWFUJm78YPxIopGvEcpVvyafSj03Dfe2KWrkazbHI+CfgJFfdbk4+wut
xJUqZKKL4gkRrJSIFBuw9nFS88/lUPmgSOLh/+M2gr4kCuNGIP0qX/vdt1pE1DJ/PnfiN5PIxb6v
62kOCU0l+rGnCY+ONsGq0vJDOhvr3TOFO5LVLjpJ1IkvGPJ/itj/rzwwV91/bWZ5dFajKZQuIBce
MZYJy4rgj472RYeMM7zoSMOC2Vx2an6aSvdf0Fnkh5EVxNDOOMLTTvNu+wbgZEqG47L4Pto2DKCf
gf1QQN6Ssum9flZZ7uGnVTCe4DePAqX26GSGB+uGwQClrxCF14IKh4UuwE1UHWENl4OMFg3ebWhX
aovkZLqn0D4Kd3o2ynNMfzpffvHZCzjsJPONbO8KdpImH+W/g8V9Zc8iQ3sOvfD6NP37T9eSgv/A
oVdqEUXOJ7jDYDA7lpm3IRhYE8KocXXawdt4W/VaTigxsCMDdjK5wIsx1fnZvGMmyYHXsqqSoDcx
EjHl7ofgylwallp+qri7udByx4q2ktYSDSzzH0o0ED0Zyz/Uw95HL4jU52yhrLGO7xB0fNM5CM/p
ByDsOMSeohUXvg6Bswo+UzUUm5790Cu916BuxpcaiKE1PmDYkFtVky4KQWtndYsmmP25Df1OyQVS
jYVplqmVnDnZPKPwb+nbosEwaP2oIO7sHCZgs2NZtu7fHPNk62wbSofmlW1hcPDnYR9u8OoMsIt/
g7phWlZ7nhgMyteQodC5jNOWRbtS6TxlVYAuqtk3J0Z6uaIyaKll0o/hwrvGbuCPdNEh90psMKq0
Ui7bftqMMR/s7zB9c3UgF4kmtPO6ZVmi++BxwyNaHFo7TO34DWK93tPxtSgArdHOjxPwsIYoe75W
jCD0bxwJYK1bR7OR3AtxwkIwZoq4ZtCNs9n9rhTfqublXJ4+kKQ5OFm+GzYgwPKggg1tRNo1jgiM
oPhsbWmUYpm9PrablmpqlXgfZpQ3NSa8MgF1EEnm1vSK4kDsJpKXkNsaPyN62jhMByst7TgDUicd
LEXucP2sZd58N0uB+t9VWiq0aDFkZ7WF8UcXiqSBZanAoeJ1JjbiNpSfqz5Ozhm5UgA/TPleWPQb
CEKmvv9H6fDN9BwpeEL1I9cOc8iguoRWMHhB1nFfRidP/tMwWgF/KMCdFYxSRvhqTv53RChdLdD6
64mvX/3KhTlDxIeQ4kofFhV84Smpv/Tgts/LhOrdsNkNDTt2QgnPMYz2OZBjPEJO6e7ydJj0yxEa
O7Xali6tk97ibvBimXfE8kauL4+0sLQQvUkb0pLfwMQ2ANqn0FkxNUsQubeYo76gEwDgrEzRuINM
sHw9vonD6KetpNLCIF/6SbuxL5FFt/lzCqPDfy8/uKTZ2V2JyA3ZcT9xyfXU720rGV6kgUO0C4Bo
rzDWennjduhHFYsxUcIGJgaTwuRcwBBxYF/0HR2VhnmI5Iy5I0qN/tpXo5qLBCmPD6ZgSMqQI4Pk
l2+it9SV0LMMm01XqIEwpZQKu9Nvl0ZSUXn/zggSK4Md58iPoKg3bT2xoQG4jiDkIe9SoyVOvsqu
ozjQIMxY3ADHDSkrF3cbVBLs4/3GUoe7Ej2TfgA6OK32XVdOFUezLAvfPCD1aXat85z+FcKjxp0j
6LSN6egtxyqpu0OhvwHcb4uX8h4zMdY4xYzlwV5BO8f2P03a5DXKpOfoTsPDXsxAJKVtWg3tDlpU
Br80Yx0FfUeIy6Yhi0G0oAqK1gK6hIGWgeKi4RsZKOBvSPlYEpYD8FMncBBG5X/UYl7mJvp/U4Po
i1fPxrJyfKedUm0s+ickesDZlEwAH9U24OGj1FgrUw1UFbitxsogo3nmn2kjV8LHdc4Q9/HUf5bI
ikiaKAmvOZDp0dSrE8U1u0Yke86ox5brpu4UTEQpTCRyEVwYiPhKmIZsTbMkh37BZg50av2On14h
bB1g3BmAapV9oxP4iNOzemHkcma5Sesxj0E0hwX8R1tEhZDYzKAO1mbo8YW4MPrsUwMXkcti1h6d
EeZY5+RLjuQS6Bg6H6qEfvsS1OvA/lqlrONoSUzoinnhloR74+DjUSOh+z7fFMZCoj0zCCAouTKP
zRx6Fq1pxqtKH4uf4a16T/Et/NDREnNHyTfJgVIDaHZkjx0D56UF6YDTdkqDQQYUKjvUzZlSkzuY
MMHhDTxbQg53j1bT9lXN5xWNSCBxKeYUs6KRcCKWp2x9SKlV4ZgezHAmeXd4kWZKO6CplnHcdxa5
K3DNhM5AFlNQ7qgwx0Qy8SeV6qNwLugSfzGgoQS/DnuJm6nSgk9s8Ob7uYjeI65tRH/2Wq/h/Ub9
r7gzxhaCevyx6iO3hDtkWpyzXhZ4wdHwT0h/P3KnKqn5na+szOv5wtBPc9rz59ArHn693RymIT7Z
B3hsnV6IKhGPNbqqEQvDDRNC3+aACbIQsiUOrv8VuWNbPfjk9fKJ0q4E8ykw7hbH3dmdiKBKxEV4
LnHx+i9JL+IPDbeTYqYqXwJKsofZPlU2nmgMH3FktM2CqhLKOl9PiWp3IKevX/fci3kWMo8FnC8I
rHejWHM/aYP+FOQedBDbSIBm+wfrq7LFYQ6BpTxK5DAJq+Msj10+izYIIi3fer4iMoTkocyWC9I0
z5zg6NPxHrXtYKd5oiLbQEY928BGPS0WBI1IsDUca72rayl1MIb+kfz9n17AUX8dJ7q94i5+8WtF
JQgT/sVut5ElcqEyMT81PVJF4BNSzRqQ33RYbeVPB09+M0vUkCfdXmUNGaBEt42FjhPi3/xW/mtb
kL1MvSQlE/da7lcmIPx2i12iycjFG6/TB8EpsBXRTrMeP3kAPB4g2s7HlzIRm93c1TyZFNpQcVPq
eSTulUxU6r0liFlG0iKTWekuBaBrOTnDfi4xuHlmbr3LNnSNS9L/IOUgiPfCjjGUJbCz77Hwsh+W
DXS5Hlo8tqpCh6HXqV2v61/0orKCmIRXa4ZZUyspJEVdom7Xzb6qZGgycpULr8xIEkEYeoagXsvB
Rbv44D9K4ZuAThOKbGu+zfrrFMrQxWCgy330FYI+kl3pRKiwVUYdpICZVebCdhMXebDkD4kd7Glg
5K51K+pOmmZCXvDEbWj7U4c37qAFpsGDjnE+wuJDplXrwpvBN7PwEb4xkhlL+Of5ogP+51hPnn+Z
o6kuT3k5kRN63F9VZ46pfVnHt02mG09C0ougjoocTc3aiHM47wXWwQ6KW4yFj9qg9h0mCPMKp+uO
OfMUQoIknJ/Dy5mMP7pRZSzgJ7D2uudN0fyMyhcAc8FGNtMjryfJV13o16AsTPWIorFq7Hpld03k
H3J1XVrDg07F2glaxx1daJig1BjLLfm6stle3nAFcaXiCmqb9W7LqSQ7PB7Arn6cLduQEo5lWvyd
Z1DO8SECYhcAP5h+Ur8AV9G8qBF0Uany3zdIDa8yFxoDq8AYKbd+N80LDGrrZdTcMcDAT++2Gghk
IrRhGUZ2iQlI385X1oFfOT/9X1LGZAp1ivJcePhgrZp+9GfuGYTbkFsPjnZCFRACR1QjZyDaboVT
QQaKF2mXpdUSJ54dASzO1msz1Gz+6piOcwrS8qrwlJSgWNN8ghJ9voBhP6ntqUZRvqONKwUh0/6b
Ol609jT7Q8N/Il6dIv8cffNByJukpbyT9cDufWZANXhsW82pZI1+6F573po8ETk6sgpigz99dBQe
tGfXeJDADHkYDpRGjq7t6TI9dm6UfI9QEs28/mWx46iscf1CK7gaWE7Hx5Pg/d4RhHiqwQaW/9vg
99pqU2hSPt27Lle2JTLGKv9NiScS0Avanele8/kSSakxviwbHrE43UNYWvWKmUfAR6u4xmXyv+k1
1xyGn3gLW5clXNEUkPpVzSr2hMxojg5rdS38GsSVUn03CBxGCRW7qQ6af/lR3810Q8JdmkItJsoU
06Bup6HqPcm3Y62H4aV/s7wdOp/yufUITBXQdxOLnBILJa4rIYykTdJE+NymztdaHMI8kiqsgRPV
Wphf7Xt81cKuwDpjwZwNGlGmjRkEdlRP3JXLVfayhSLmItfsL3C/QR09JSHnpvTykJGhGe5fcURw
wvyrGRIIG06HQDA135rTaTfN4XX/gHpqJibn3YTZMnbbAeUvdDcxfIOC/ht9TPGb9UUNkWMRenBH
fUDCsnV96djUBktu8mJZbViDv4ThCy2qsMD1ylVGJrupibKnqxeUwJ/tJu0oFP3cbsgpnBoUFgk4
Ip6SatvsxkTs7CVOVREuAeEngBMiTG9zK0ymUeQt3MSimUTVovT9ta/hpzy4zv0iSPz7IQPIBJwT
DjUvnHVl5nu+8bdpLFQKHhCfbIMwegQBrDrbNDPtqdVhvwYMUQVuLp+w56SjwaVh2b1vVQqOxTbJ
adq0uhhuRnXanjo2e/axyoyAcuLDVgMoF6BVaWrg2+wjOcUxOEgpp46l4IwmdLXd95e6wJR2vTWB
S2Lq2uAZbd0gyILlNfELJRew5nblmSFNZumyPVG/DkaXiqvFvrKhvmPt5x/XK4UGo6bESYQ3gOYI
MB9GvQmz+0JdmuwppRrcQ/7G6QB4e6geNdo1OQUrylRD9TQvkG0b/KKm6ZFuSxtvQRRLL6my4na8
TVv2KXvty61m8gE5qndpyokKi9nde7O/6jS2H52+HRcWiMEOFzTuztYgc0Vetnq9yi98FpxCKZVM
l9yMkv3DE25NSi/bLsctWW/IjALVfPw6f8UliQea93U5qBQKjiTK/5QGohLL1vHLNN0tYTsYSplq
uhef5PuH9IGf5X8WMwtBAKPET7nLDnLOzIcvgw1pYbV23aR8tu7+5aV6AmABQaqNRkxm4jNHaXxb
QImLXvLoQFPy6/82omuwtRU4vfokVI0I+ZZYMoT9g3q9Va4qvdG7ZQ00a9MlosDFPBBH2cNGK0BC
Q2T30NJkIDV+cAMUJerdCPY2sc7E2hCAbQs9qHiWCRfMMvWioFOiAl3cSNV0ZN3G7uxId24KFw7W
0b4EQKXg19b/BrzHBfy2r+PeNLRpmrBQP64NxJcwoiDZg65iEm2w9YGYJae67rVN4dgQrEGLMLOm
9jXZNi8ux3G9ry5Cb1RnxRJi9QeNdjXAIXe7VANlJM9PJX9+YnNbAjkroLahhoA6rywvNd+bhZAX
XHCMV29UNp2/reaOaYoRE1HlR98vCGAB8fztYo+zbMzLNBwI8tVGJF953Sr+efKCCcQfBlA4ezpS
aEYB/VtdMybvZ5J7yYPK05EK6ZYUPtM++KDzbaxizTzqVyyHDIaikFB2Naq7wQQ/dk6IDIikaD0f
yjv5YsOucn6h8gVFad+EnRVpzMU3hTWEksmFezb/RvHXrPa0TogS0bMUk88XMBq2GSAibk088jfA
llGrKiag3eThNPExFEPkKqb0EgIOXXl7sVmLFYA6EXtI4wJtp4uzBoFEGcowmZwttld6HENbIwhQ
wrve9KrxzrEHqmViOIz2OMNkeNhJo92e82pA+vPOoYDC/+POtQj0VPiN7KanU+XE/ZiPbpQBjuKB
z6hZ6MTRA1Ddo3j0Ge0HRRMBMTvvBo1LqCW0ceBfXEmDFfHHJhf9YnlJDHYvkwTkHgHXKVz49BUU
luFxO1ETlK++C/dfhHCyT6x2RNMStnpRGibGRp79honQtNXKn7WntzIB+zFz0dWkjKxQxQTTYbLd
XQSlqyeVTqsSCQMf3vxh/BQnOB1lLojlZP9DZAOahS6HuSIIUeCnSQX012xB9xf5SlyCn2Nh/f9i
7gYjs9263sUFOS/rfiE4bM4/vhiyWScvVsetWFxwEBIK/nFJPnzxfZx+4Hc0TYB653IypSHUqqys
VcQ7ELw17Rk+I7rMoQNjsFXeHh4fhtNNH97pgP2BjftizygPU1YpSEuycy5t8IH5DGUpnuU02OTX
z9sbeBbA04MBwCTlRleJKPcMOl+I+HXmZXNg2lcmUsgdRhYt7IEozqMrupKPF9wYgy8fc3Vw4XnU
7STyv9B37MR/uEJZOvtfARX1rt6dG5E0CBHKjTZW2k+ZFxlTmduo6wp9wFXX3+rhPenji2weIdxx
PdAdO3QCqWBzkVoz0rfEcipWrVb9rbtRiOnqqF+HapVdfg7jpXliTHjjknl/OFZXEftsEFvesqik
dogDExG1+tRGCTJse4yOdU/XH8/qA+kfRzf5wicY8hMNIybecL9LdiR2uzD/kwRNhlfngLqoGPSr
Tekf3XOHM6vY05q/Lf7kN8DnT1a4S4oog8gXTRZ+/QrveBCaGniZVFuwUMxUS8gUfS8GODRz6VPH
CeNu8S/eR/ZcIwJp3e+iGZc8JbLjk6jAYYVjpSg0Fvasthpja9odw5+W8Dmps9RKYwqPvl9qMKdw
4fdA5tY9VcFlYlsAa8YIcdm/FCNF//zNEhaC6PlYeADRvd9L6u8PyYX+wevvelb+sUq/+bBoEoCQ
uSpE5ArpN/tIwDLrVbLeI8FKE/3U9SeC/MD2FCpQb7f5CbJ+X5c5R8SnPvgcbSTooS7NwvO0cByH
Itn+6kp5QSdTA6VJIFAHp0fL4pKfkwvDFZPuqDXeYnIjlc0Hs7SqJH9Hr94pM1LV5sh/OzBg2KUs
LWHsw7NnPmvL1FmIEZMToeVmMDKXI/lECpKKZmpSXm+VzyZf1+JhdayP+eZwekH9TD5a5Ti8LREB
RvDARlgFnJ0jNHUC1FjZ+Id+7rjROYzrVL0EvDBm4beLpZcg07EugfBavbjDWQN4yY640hh0fYDq
zTtuqi0MhzIohzHpleXL+VqeCi8lQa04QEHE6vziCRIctvL3Y7PgC77cebw+67JADwtiLd3Pa0VM
Yq+wQBOxm5WGd9piC2lx+cfxAJbu06sqiaUmO9yafHixbdu8OEjLt15YllWhCzLQQ5LGj4t1W8ec
DND30aVx9Gi0gj373kQ6P/Ita80ZlVkqZAckNUMWAOKijKhomjIJIeQxYiG2VQtYmQ3dDulwL/5Y
0wB34edtxpRrs88KJex4vFrI2TAtIS8HLkXfX1jcHbP/MXD2ieHNyCUzwjlmxiLtQ6sJ2qnhh17p
TxnRVsjmAMzjQPPqHJ8NRlWZ+zyI6uUGLoj+sP6N1BVS+4TaqrSec0Ivq4I2JeJeRnTZZ2weXs90
G3aoxP6oNNl8GoWeyEhrVmC2U3S1Zoltihg5rBl3ud+A7bmOYxIBzSMTMpI/sDjqQvsP7X8MV9rL
5gU7XoKIQICSnlLCDqFavvdCaiBgqWeIZdgKFzwhXEe5DVKcj0jfKCYz2rtAN8I60fcea79BSS/+
bxVjVOMGp5NwMD1c1UR9cTMRV2iyZUiXdplxP/LiUNZtp2/W6PjvBjpRu7tCidmMc5EsmvTuZEoA
Qshisl220OXlXrnkvdwFV8kXOH5CjepS/PPeZ5akFJhiQKjcpm3RE9NFCPm/NfQE1FLY557EcmOP
/PV44Q4Vw5sq+5cZDfQNKjIaPMBHhCEzHFth9ydzLw7nhWIqT2K67LdyZQH8tJFlw2t41qbnJvIJ
qS+wWOiuPD+EEyCdhesaYX72NMwkHLAE0JX73KFgws9Ydu3/bG3j+6dR2yhLAJXhwCvtex/G+W9J
jHE4VVFyTruuRgjt2z0kyckir5JNnNtDBVeXPL2SjlSP3lE6YJdnRsToPmTtAdsnaBrkR/z2pn4J
in4yqmhDUhtx3Hga4c8rrzdWbwPqqaM10prtAv2+1ehS7nqh9L9ojkrInL1JmDxMPSZ5zu1JjRBO
Ppp1jd6Hc3V11Sod44cAXzwmp9dqG+0M0l5LLcNuHh1yUYqMEeCNqwejgUrVj/x9dTNPJGLh2ypU
xkr49/Rou+JQcM1dDP+rJ/+q1szSXxF/r3kKuGJbJCyXdHIWj5ywRavDoOinssj/r9rySXGAZY69
ISwQY7RHzu59PXaRccjrFOuUKhgfgNLpiArnh4puxCaRgk++U5YY0NRzxCLU/eL5Vy6TQNF1KWNI
nyhMvQHv3X9y3eaUxpaK6m5Brm2JqyuuW21LuYGkmiQ6lihfG6X5QX3Qx7A3Dlks8Ak/e57LUQUq
uE4oFyuKD/gdEQTtNx7UriajVhyEd9rjaDAi2pQm9S2nz/GYoISMWz/Ncc/6cuDcwDjlc/qfc47g
r5LrL7WaE5oDWM7qm+ipsMYzgDV4l07BWaytt9GnhE7qnSEus55PYk9WWWSCvxJx/RVNnDMxPeir
4bFO44ZAesl0lSfuxwAZQRyVWH5FVAigJJ4h0/qqW43ZC2I4UQ+B3IHkKzl5xjm1QEcbkDH1Rxsj
G1SOvXTvWeNtGFu1mLD31cNrb8hwgj1puVY05fIIY4kiNY7WSeMS562Sz5tAEqGnCnajwFw26at3
1CKM1vwCjKM/kWknltZ0ETye/JYKvIZzm6X+xtv5IBS6C05KFXQLCdnvOQfPCETzYfKXDcCs3tgO
pwcA5LE6adhsb4OuuNdiRFzz5hvkbuorLE3VHwxNOVIZ+TFZzGXKjCspQk42QBGwx4VEUUF+PkdU
g1jr62YU6823PAagfFx6q8cOjJf+bJ+W499LnKWXIL7IsGzwlBZaLrrK+PYwme5xixxi3x83ceDj
wCZjqVwI5TeK1yP5MQH/ftWYsG9f8Fuglv43bZoViOBJ7bRqSIElaUI4ekOxAP7cH00PKoodXcm7
DRfJokH42aqUcIob+fVljR70Ge4jVeClPcVZ6LILy5ZaVi/SPRVONDyH9UDnFIg42+OaMm0sVkzj
bWGKtDA+yYm/mX8Y4G1S96USe32WoJ/yENtnQIPiox1uxtmDP+9bjzkr6x3GoVGJDxWsr91VFLgp
mXWiwN+HbZw1QFtyY57n7O7i/FAVTkQPyGDMFWVQAlhttC5VZiw26xX0Qbkn8L7SyX4P7+zBJvJy
UdGLmk8R3W9iwqTtR5VaQy7TIsjT5FyZHdXHU3kMCWYr+qChfmEGQA1/nFsbDg2sTrgP+BgAZvB9
/QTdvHtT3rZ3jv4hX7BHhzSPWizENyRyjOxf8ntSkIEYP3OrsG7WIYUx75jkNdfmoTlAcEe9J/Z7
JOK3m2JNTg2a7WWrN0pTzcxLOBvcth1/hY3QdAMUROHCJ0DIHU0TRKY5HuRRQGTSBc0+0X3g1qyE
TrUhdKBYI53IQnZ1Snkga89qrlNFIBdQsbOQA/vS83paW3kD3Gj4K1TLqAsouluI/SA417q6V8Ej
UzVZJYISkv6/l8EdYKu0nZ41cNgdCVuvWoNAt0RZxSMLhmbbhOFr7i3epnPn2v9pxEAM3Mic/pvD
T2/Pq0axffzprheO3n66zHW+SLtzDUFS1VS96pofzn2D8R1ovbdYlYtNI/hfliRE4J5wQukML9cw
ClYn9AI+/AUMQGFV2K1ZFagOEsoqJuQ44A5atOl/+yY38r3Swf+FeLX5T3A6FVJ9cdSqcnSqHW8T
PNlFftuCT50iVeubKyrThtals/fCVT0exqgDCAMtz0pfEAGgiKcov1c47udkz8nGIylkf4qwSm0U
zAh52iQZlG5JbkfP8gqRYn9lHRAQMUoJXSph82Bwm644HdHd8G3yBCuu0/pkEa7L/IXYX2IpUqSY
QlYr0UtVSqVHOdE7BXinAfEmSsFgCTEZao+jUG0uyYVmP3/EX2s6Ml4pxlVk6UIiSy7zabGlFWKz
ONlmDfUP9z8Y+QB0tPNNQSuo34xZ4k4M0GwuoUWBi/pycKLauUbi21vSZj7DQ/w+yh4dL4+Dh+7C
bS+vhQOP6tfZbVZAtryx04BCMzI26Sr/DPw9msvmnD4y8y1c2hR971aj8wM2pdAplY/a14Rva1JZ
Qs5VJENsDO9cB6e4WuzxlhHtH9d8Cdotq6VjtgEkibC9PHPFXmyUNg/u+SQvat6emE4oT4A5uSej
SemaetBm9xm/BqaTK4szi8DYkEbMpBxX4ULYbWqaGwMSgrWHRjfkOPptXF3aOsofU9i9JhTZt5y5
s2g1hw+4U7uaSNB6M3oI4R5G+AbO/sKXFfgQTDKnYdNjm40l5dXKY8Kjeyvcuh0/RJV7pUngd8FS
kktt3BF01MtClJ3R3S91YdNLljr0br7v1ztg528tZATzNr8scG6HzjE54uHGukN77TE/gaeZ+3VE
hZQvaI7exypNCO5CKX3pCsRSa/ptS7giccomH/aqd92tgPQupGSiMXJ6O879rtcjWBJGgGoG/aSf
NmMU3ad3bD6WFOTraPNlLvQBDee7fgZRaIjYGoWfCWdz3Q6FYvRTfTFznkAoGNg1xMVZQgDtq/2s
8rosHAmjIg6CNe6HYZhJmxLQyMSUBqE+nzJAK7CG+oJaaXq1LhZDCbevem9+Qs4g8EAR1CXZhOsM
E1aodObSeogX1SBBKYkG1h7RyqvypRJ509WltGfw2GFfp9CpM/VDuHj6mxWFeBDaIS6GF844Jjau
jKfCBMsPZeUvBc9glEd77FoxjcgxVVNWBsKurLpOM60Oaqt/sxythddgx2M1Tdb8/TDCjIkKYPXO
oN+vWf+SI3+F7sPo/zt7Qz7tMofhTE2/gE5e4h1k8GRMMJcyxnKR7+krGnlU/6J/g2/baHaOXEfG
vOI6wq7Zv/I75iEtJiPlQtF23gbE6bNIuMGrNxlUfhmiFbfaOIOLIF+TSAXgANQvW1N3fG3G7Ges
mWHo8/lICpYqQASxzPuIL4cPKoEt8tBrkrld/phxrFWgR92jnlCY/5y8ZVoTqHFaZu6zRz4Z4Ydv
rorryAPfQtqkoNpipM5G97KkPx6DsxNGgdRolKolCrdmt6AA3m3GNAj4ZMDEnxzmTHNS9EJFNbqJ
W7F+ZqRhMkFoo2OzEsaHPoYaP58H/khPeOAIKn/TiHeTNYqnXNZYCpaCbP7XuKrVRRN2DMzDFasF
179EiJWzgYnfRDFXIsqgzDanADbdf/lppGYfU6crz1PKUf1bWm7uQ6UYjn4UdEbYR06LQDkzs/Ae
mv7GXuD5HkwmZVdD/5jlXEkkRUbR04Ofx07FggIMjn2BrNAQgecy8wXKBB/J13kVekTRx5W4HvFU
G5RsNGOG9OZcl1N7bwyh9K/+POFJSue8CjDe+Ud9a4/QZfrEpWAPUgXAHkCJqLQZizTK4brxeEpX
dwJT1q6lOpifOGImCAERimQpA+V1IcnNRrb6bU6z6qnPLgEGxqSOLyfY+sO07ebl+pAeFuyzjaBP
anpO+/5jPcjT9xUhO/hIUJ+0AWd5qD2rLZdyQny9ebhbtFp3NYtS/BlzAD+Tbj51Aj82xvjU6TAt
c9aDbP6D8pQxLEcMKeYVGIBPWXuUFXsSLjG88LsODjoz+2lUtbAgpbDv3V4qcP1SIx4Fv65kWHcX
0x1sKVYyr4ctuLnqfkaxacnFeCXSEfnATahSiWsXjxzBn1JQuGV91hc2dUlV5ztHXG/dyp8ZqtA9
Hn4GTwP5x9KkYw/+EImZxaxvVrycHchmBI6lfhPk66lxfsXZ399oqPpP6c9wGBU775y2Xr1qTuUm
YRZadFrgOHfYfPUwb+AzG2/aSRC/sDLU6Oj+cwyhghP7T28HVi3RjAY1UGcMTGbYkIWOUHR3L9l6
MyMIoszRVwxm4/ZoQL3YAolNYRgvvJ+eYyqGPMxzCvaAJHk6eoPEXTvNiBb1lJef078euy5/stso
/EN+pqNcpQpeyhOMFhdBE/qMGBi9A5UwfRuww46jj1CVZoRBjAK7mgAqk+DHDtF4e3wBT9erxRnq
uKDuknwOpAi8ySahYF00weqsuUxfa9B5QdQT3ELqQr74oTyvXakb93t5OxFkYSwfk8n5pCe7531j
RwKE7GDAKS5DCyIkapBmz515LCDo0IvO9u2SNr+tQWKQ939W9a8PkZKH0AQ6s6tv+wxoRv7Py8Gv
XIzJNb71p/LF/3lv94PBZO7Zw75qLjMLKj1Nv3kYCyegbKX9YjTeOyMIexrGIehN5YTRgAXkk1BL
i/LbCjkjRRSWML/YdNpa0mZuAfErwp1ZS/Tfsm8/+B1JahadUUXu6cGDdufW5OS/v+2483v3EhGs
+e2FfeoFDl+l4p9NkEpAEN8U4pqsaJD6jZrHYSdwrk+0+4YwUgPMSJ5Kl+93JVpdJRKLf80qiZb0
1CSHeIrB5QfXU66CPjZ9Bq3f4VEnmP/V8rTCZXMFuEl0gfPeB6yW4InIeCX1KaRdqQ8WcnyQj/U6
OVDMfcph5gZIVNMBewabd9OJquAm1rZkgQZTaCnl8s2u5cZ3f1lepnZ861I7wvd5ueRqAQlRFz3N
ypehZxJfz/yujkXiwST9+HyE+t9I8zuoBBy61MUMVjNL0fVKL0zXxqAKb/hakX1ZH8tvXukXHgfr
G5IgvRyNqEI6wvanIrsJm2qpPIhmHE/cvzzdwqy753EzpUY7yYHymZEv8NmYaqpw/aZesbrhFn3i
cGX1oSOMUnaQN3H5aU6ii29EXcLu73eCBjmZPnyV9n9s+UC/O3nyRxEQ4Jzlo9CO/5Fj1hZgvLv2
wVUvDUocypZ3XwT2J9KLKZukZ2a1temO2iTFi+x/OW9//PiK1gdlGR5L4iyBSZPeM/jiS1NDBQTv
Z+qLeMSvgGrIG7kp/44njDB6FkvkiaHp59lly8xYOlcXq0ekUNuA9j2SLw2NJXj3dLKnx3weJLw6
rTKl1EkRIC7AMrK4ZKmkKW9IVzGhC0zVmz0NyyGiObp7thQ6oCNDQv1vhj09isfUp2Z+7OqETQ+o
WD4FFoq3MfxLVfo0VrtjSFmQUXlpV470r9ShJrmqy/7PBfi+gRQRdiogV+R5wVIv35Tu02Klg8Jz
2ObYCQ3fKpc5Dg4opSD1IGHuyZ5eCOd4FCkmHH4sjESlADyjztFqUhGApS/oGWdB5/VPCM8nOwCr
M2tRnAipOHCwcl2bIl4ybvAbfhW0vf/54HrT7exExWyp5GkcnXd/x+ZrCBvaAcFvUeqk/mEtR9Qc
Pngdv3V5WJmX1A2wB/y/Nm/M3xzcCgON+NNiQUF+vMjvthxQUxlWo10cdIzdgAP2AodIlAGw7eYs
pcT2rL2wku0XJ8rk/fI51RptyIRpi5ZiCEi7KrhrlujmA8JWG0ZKjKSXQKJcdgiw5gJbyKQWdd0c
ee9Z2yis1yDh4DaCbY3CLH6eF1XRbp1QZVBo5Iw5w98Fg3bCEOKYw3Y+LycsXKGW2MSd/jg7OlYT
GatgnJUsT1d49IO1v7c91W/YPvnmaS4q/QZAOGfcxYylytYOUpk6YazjFn4J878StPTvYw04PFHX
HvaF5E3Nj86h56y0BBfSu5auw7q5wf5qT9VzlezRwvDygPU8kzY+vj4KSp5W9dBbYtMvAXdsM9Ct
JLrDeHbS47sVAUK3AD/+MrC7xT73qdlr1MTcmBX+wPMVOKDxd4KXuu7rbLl1MwQ8jqpRJal9LcUb
kJ62GdnVKwZyAnmlyRU2zp5HkO/NnXGLktgX0euT8pAWf9njnHRW1OYghSJfbR3R1sBsMDArXLY1
+bjEgcZqEKNR+WQYu4ryNHuXOQGCjc6JytW48mt8HVW4qOK/zC9uN9AOD5mccEovckjze6cx/HgK
v6wOluA2f4yYCIndzTymzpZBTvIHigZBL2GJQOe4S/hMZe6J3M71qAVOEgRSsrhDWFSkh6AaXbSO
646jsDmyxLGlRso1HaxNdzGmCRyQIqSL2EQCxRveUksakUokNs/4EaiovgWCk6OefJnM7eTThzEn
KHaoz+jRUJvbI3VQYYVVmDjdAP9MBGMCMfmZIy6ArRjjUCj0DnifEPPxW5w/e08p5+xbfbOCvtPg
RY1I5cG21Q3TVPf0gSL9ldvdk2c+66MeYUiRsS0b8p4uxO3GcGBoDgLwyzPQYnGcwEvGWuEkP/L5
oqISqHEto8wRlVPdhnUTp6DloghjrqU7b5NNZ2PsRKVOmZ365JJXec7eMZ9Xt5ka4+X6L3HTGBr/
GGJI5jz61iSCHjWQBu4Pfi14G3HcKQj1UUzQcC14N1UJbuBLUg24Pcsp9x9R6O9mgqzkGLcyd9ab
VtoBFerDmP0Q0G4N2oYiHb4wXvQ4khK/indifiWIBjbpsOzswavkQrDWEETzYSxul0ZoJBYCW99B
SawU/OHjtI2EF7h/ppsh3fhumo+++HarsGCk8856+2gfBfhTKNW6Etdo3vFDg193jvumfpQ0L1Dz
oX+SGk55LWdzAXQ0i9dgXYcLzae+VO4p2pB7e+Ua33yY9kkFIWNqO10aHayGhIcEcJjgSO5rKBCm
DqbiiT7YA5m62hZmLvrv8j5eA4p3va8B1kek4LASaDrgWjZ0khO59J/rHjwr67UGDc1mn7ACJ/mE
jEqIgKKdatB+KPv5ns9/Gdeo1cot63+HG6hFjaNPHhKIxQufvte07L8w1G3hy5LqGW0WSoGUE/L7
MRLx+IhENSK2Rz9D6n1mZOBWRu9p/mDTPxrFgmsXUhzuzWYm1LkggWc88Bl38Hpf8qdT5a4S8KNy
0/QPk0eIbOOun6K6yx5pVQ42Qxio99wutmePnsFSus85TO51tZ4xxa8zhSoKFQZFObcbnSqdRAth
GnPtME87QX6aFgNSUvTJRluBgtva/+vnTSdhX9nlMmAHWjV4ukWEly/F+SGbfOY0cEx0PfdJdm9n
slzmKSvTW0qSQjA9V2d0BKd5KmrGnRTTn0jVuhGrOUTbujE826ov9uSxFBr4ZoliEZJEt8W5g+9x
dBpCBy+c7A4FUYpe7BfoMmBG/NhBoXQKOTC2U2RcUwK93769f2aE0BbAvXD4RDeL7KgTreGYW8Zp
c5cJXjoYHlJNtlwWdAvG/wOr02eioGN5jYtQdlX4vzLHIKueHKEuBPaObZoJhcbj/vuie+60EzzB
Qv3LEV2uCRgJ7mEUfmJv9ewS8AeSmXnRcM0tM2wCoFCh5CbzEzxbKNHc7C+s9kC/UytVXbJ5VtNa
t1PevjbG7LAbhOs/4nR2jDqapjtWClrIClvNk4hHofcOZbnV/mrX9EWdoobdayGJXK2DAN9h+i9W
QuugmmhDEFlBlq4DiVvWoEWDmjgYwPRa1upAjJlOimdzqsbBtGe4h4kVclwYaAQQfodCiKYR5FRn
PwJH2r+LzaGnxjz35xlDRq+4nMNKLd92/cHGVCRvR11yUdq3Tq8VlhbETm8KreLQLDHoJAh9pUL0
ywSmRfxnaJXEA147blJNZSm1SV9OpOfqzH28758OEae3bJvWzIp52ST0rm2CBwHkgOMEGEqgWdSC
zPlTUUx0T1+3WlYlhTSu9igcruw8jx5kmvNajl3El0fk6FX8njN8T7WN4jQbatsiYnLxFgeRxBHW
9vCQBebHEeaMYLH5la1wOUUaJix/+Gkfq7/cWuLcaJeAP2L1l1CXloIvtzqLBN6b1f17U839P/XB
x21G91YC14zKiyXuh0GzJvbRShwjEoj02jo2x4hhur/ckhuvuCQcSGtwigWSa6JW9Dx14pr5DzBi
komRXyBdvQzssQs281Vis08tjLCUylJO0ILzPtpBOevxAj+VdKHZz4mZLpOqkCnSOXZQtR9/hE+a
x7m3XMVJw6zIo0hQCFjgz8Krpd2seO+Tz/63wcVf2NNcHp7vr7dDU07Yq6GRYpIb90DjExsanCjL
B3OCzUbSD9eWBss73TIrs5XeZpxZG3sakGO9KBBOwRQsJ5hbqpEdPiJlzCr3goN4O743/lT1rY7R
ZWhGkJKX4i1LJ5p/G/qEb39A1PZmqqJDPOyWrP7Wj9EfuEScoqvdO6wykcsix+bQbi7tjVsRMdE/
gCQ7GPdV/4OHfLswy7I4D0fQ6tCeyVjv6cpW8sB6vIbbjsOKoaS/bTJWAWtk9D/XLK/t+ljBCyzV
6YU20CbLnyxYLiEOx539dsf+ohD7hUETtuUrU8ukGadE6rdJ75BAold2gsv8kcYb/6V8+ZuRE6fw
KKi6qJHeszJRZfFMIYyiLMOB50pPxhohjQKVVuesyHJzlAzvsgb+jRJhKAhH+xOO9e9VzGNyKfAZ
Z0BVM5TCNQe9KJk0K1HVbw2TPifMiLGCZyok34VWtJaiDb5AdT4vhSmHMJzQHAMKIub/VEL7qLTT
cSej/pT1XNXRYKYqqfa0pE+Xhp4/mM2vbsDu25fIAwqQ+Nuz1IxYAKlBC9LQOnyn+4tZrjbHKtMq
l/9ahLtnLkUR3jyMLNCkZMakInwznwUDR3GcE5FHk0gUXZvMZFVAZEYe+++9OkZ7tQUP1S1uWN67
hnWGAZPm2DpkNkQ+Ei8EAIyYLEfelD5D0T9J3S8daBGZLncD3VJ88ajtI0QHYwTc+TvHviE2m0jD
1nloAmFeGZ5FLfz/P+drGXZA5lnND7CwlVrm0+2T+ubDRKUOD+AeFNzVDSBN3JBH/BJJM95iXkm9
qi4Xdn8/wmg8Fh03FK6zBJB7ujYe7v7cSk09yasgNIc7uTnm17SAuNn/iT8EQeUWjmNRrFcA3R6K
EFbxw9Z4EWMAESzANUnWnlwQPIKj7ylpguEmb4GIQkzIaaBnVuIVCApGsGz1Oom2y1ysp5J5VI2t
NRrZRm/l9JkLPnneDr/dQjnqZctpcFvg68+UHnBMvNgxhF6Ci1ommGthP5vMc+yAz7ogVQx8IXeF
TqtlyKRS5i8bS1vfYXP+ht8oLdxz+fPGozkWNxuC2W/eAaHLr9qfHF5lwZxSdNKQC0rxihcbBB6h
Ol9erROlLn0bDkq6h2MeutvDM3buuAfTfEjhZ0lDWbsirnG5AYHIpT6rUBp0gXK3BfkUTrlR8sQA
nV3o2AbzavX+ox+io3itV3NfxxgYpnotJ+H344xP3lgVepKQi5DHA8io0G7UlR/zPWGLD8LeQMLZ
xok2i27T0DFMOvZQZvfZRbr+eSL7wV4kALtPkssIBF0Ga1Tc/SHrs6oasbG4TA/20NG3juGmMyHV
qvTu0CkVSImwXttqGvSV3rg7iS2Xe1y7b6q0cE4WlzDf569QLNteUMAZpc5QhCpedNmWz+4ilCEQ
8O61EOJ1eW2eENlWvbHsidAKUwfnPGVsUzUtQPlQsyGvj1p5WL3pIT359fzj4VC5AunyM/d5tcjE
O3IKtHdAkAVeMLQyo/h1jOwjlKB4W0UBkWq2NLWgw+CnlD27x3rkJ/w/5c+R/HSgUSew+fwAbZSj
L7iTqA9KLj4NxBj5Bk12L+/KxlR4kwcKBH1nvyQ88/10rAN4GsB87vRzoBggzG6FT+wLaJ1HuAXf
nEDh0+GF+VwqbYkdX7bpj3oGQoy7SdO33dhOTV9LfUkCZADSFuV3owYjucNNZOfhM0dhqIRcf/QJ
GnbunKd1ek9W65/xpPsWexOBr5YBurF1jpG3CoZnc84DNd1CvSEDu8z/dkcmuLuzUiw1awQWzUfG
80Tq6oZKcT1NzaKNsf+4k1amfekGn3KVEmyvydU/qB4DPomdy8y8A60ETnq0rkxWKiDxjZxBebFu
/VTQ9+hhkbC98VvLtFmCgz3qDfwlx8cS5mQxADHVm1l1ZZPKWwtLU2wY64CUylLFn0FPQO3rCGhJ
aXgRoapuI4J0r9mrP1Wz0URuYXcFkocYc4BTIchcoxub3e0YqyNXoEqoHt/NoU2XrLttSj54Ecbo
4vyjGB7iON5XNj5C8COmHc0aT4SsrAP8v0EDml5DhPDZCF21BmvFGnd1hgrzCugJeeYoxeVEOOpY
0rLpWHLE6jPkzbK/PMKAtKEKa0AFpHgvFdV62dHLy9iPPt8oGRBD+ndHPJFDpOfPte4hOvuTh4fB
3YbQPZEFi1NXtZTvp3lLYOjoSpCuc0kZUzUslkQDvhBvY6QPp/9FsrlePU11zSBvey+RGN4JRTKa
SZUAZIWGxnHGtOMeU6/n1oIQ6szX7dcQMYUW1nMaeIXy/ORKCVp5eLmnMOyAM9/4C/rWm5HlPsKl
wjwT6CSec6tvyOTk1vxbTgmPvKTCIXmkNZj6vpq9Z6gV/i+hv461zRSmrH12V8sD2eYxLMnQGKyL
+FWbeAAOVicbUC0A2ctIFvr8zyNuxYamp+ZfFgU9dNlFPsG/hrzb4eHKclS6r/vY+BMWIlgLPSP7
QV8CO50fK2EGERwBcjjJnniZoe7cadDEatXJW9VV4ZpiTKflVOb1dWHp+UcvsuIIGRhkue0SLA9N
x5bmkKAeIs+J2RTli9jtUOYXbLNUkBA6ICF0ZUykJYY3+puWgQ5RcMm/N1KyYhdPtKbUNktCdKxQ
yIg1+xAjQ4r5v+2dPeeLhDcCM4/xKFWAaOOvWeURpdEBd71WFSbdYdA4blPsItilXurpOk4w+KTn
oyoOHhIzKKMmSLIFE/R7UePLne4WZ2fbcoukRqaq9EfYYTjvzojLrQMXghLrh/EXr0jWfZYwKzJE
p5+7i3mBXcyJHPxgGI73KoIRMTvSPXXZVBsme2C41CLlzjzOSQSolqQi3Vygg4vxZnJDqDGu/BnF
vOZ7NHCR6V3blR54FtfgVTHe45W8+Y7WudX0b0DwMKMH1KvlNNRg39qdd+uSNALzusabSmCyV3/0
yqQ7E61cTmM9eK2q0/uWe+CPluYmi3TMZE4L9ZrjDuqAv85H56Nm1VJnle6tsExyZLpiTH07FA73
/GXUSlI4fveZbjwkD2qNj4dMLDpx3dBTlONQYjvXTVS/QBbVxl+OgMTjIrYROANS0L5/5bay7V6q
cktU00WKrM4DHywk6JWpavHcRSIkbeGDARWt+Z9ByAryPHYiK0E4Sj7EYe0qqc4mwOoCIg51DSZo
sAvV1fUMIYLJk83b5o4b0s9cNlX34uHSa0sMc7WMacppzPsg1PTp6jqLHi0jKXA3bMAxKT8mI2KD
oLgqz7OZFY6Ql43xmATULdDek2EWVCzuM5OAdqRScssANsuAYAGmTl3l+BDNzk5W15VQtSx+IWDh
9HHxB3l0RuTCp9tXqsvPAXQTc3KuEMSlykPzlRtb2MWNnOpD4W61LfGdCS02ohals+XYARlPmHrL
tLjrmop4Qub+Bv4lYqOz4WEVLebW3x2oIvrdX8KM93Zp4fK6C051A/JTAYypE3z1g5BariVzckQN
IiUY3nekwCLLA4+d+NE1W4zNJgOV0bUDrL2DX93ipeJTIpI3bJWCGPaJYSAIpLL9MAf1DfSkjOgm
dxGPLlMMUhQkX6MyUWFLOGg+z2RGeDfXFFAPICFFeWApMW+qqPlTbSgRt7tG2M2r0SHke28qnoim
sSuIDo3rv0a3mA5Lwplf46yP+2hT8FjcgAACEm7N8DCkpoLXw4xsrGM1O1E5ku71fLJBhAOInQyF
vZMogdXBrTp5KsAzx8XmU2YvrJGXPiOjBi6QQrETSYrIkcgM31mZogmS3G8J+xAym9LMU1SAlDmw
v8ECbf+su0oMZjr0/1yecFgTHGWGSTo2ZeUTN7xVSGwS3yjD0i+C/7irAZR0gl4z6TNey6gQYzhi
8KC+0CCVKBQuTTLaprCAVDuxbi5964ruySo2b6UgqgXi035JX/lNcGKYVi1db0LRyV6w39JB+Z4W
55Sg20PKMlnB0YyF2MdPt0NxBa4VwKLdwsa8Y+YqfjKpPjjzypW+qYVuwu6ZR7s4ZR2S6tvyqZ12
RfbxTTCJDrXkh05IafPLRir/x5sx3y+abt7tHmL+WPf7g0O8wBc/JcyANmUkHnHDiV/5aE+W9BIo
gqkZoK4FyPiLRmlCmDqfQQTweYkjxY0oz+9PbyrXyl5txUjNK8YrgT90GbfDBj5+OSe9FSCwyhiR
SZjZB5iaIg6UyWU7hD9tKZY/mvJx83l8pS/WNQCfaBQ0ZYtZHLOGqjlfJh5ztsIOdi1QDrd1JKvR
2cyK1uhfbDA0sjqwUdleNt1365yAMIJXph1zKKBSMQxRm5kdiTv4KTb72TG+Upav2rbQDvhAQvtz
ivXkBW+k+OPdg0fRU9IMyNvHkHX3AdV4VwD12bEejN9a5eKBEUTA5YEaVo0Rzl47qpw1HxEO5ZbU
aX6+wIe48zlQfIPpe2U/UKt8gNDUOenX14xx6WExbdrT3wl0nunqhszVPJ7rbYvPTrDwbheTL9Zc
evrp7UDhOYyW8+MjGpTVlSL9RXxGURBTyQ+2xHzta3bqUjf7wHylc653XwETA/RPjSp7IWgFqDFE
R9seMAMOTwQ1NyaUKJb1U9WcgXeDKYlRTW/Ac3KBb/K9ywBfJ/DHo71ivTRmvh6lDXPhWgb4RM1U
ZLRHXLKay1HCgZ0b9UcAL29IL4OCHCzsKJYg7EDYjJMZ8WOY3lIxBolUTx3BaaQlNgv6u7AGw16G
TZ7S4j2TMQLHqL7Pp3vVlhxoQ5Zf2P+pdygaYiglHtMysAYiWUEGlmZbrJuaBZqXriWdQBoYmmYw
TtX5h0WgDZCgppO/F5tkHvl4W4nb0N9dwHXKM2odcYwJScWrbEhCIWkffDAubBSvU1T5QAZn1tba
IFri6/qHSYw7OEJOTS1sNn+FXI78AUSEo1AWXWHf8fuInKHqYvE+o/IqBhleWHhz7EUJl5FSGOBq
Wm/rZsIvGEL99N5HB5jFzuxZzAOHgVUaCIKh1XMQGKt1S2774PdEFAAKxMwkgcQQvxXJa86xiMvT
IMF1ctUz08/Z8eu1/6L+PfnpLB5gM0d2Lm+Zjp9mfW0NxaKdGLcR+0QAYhIuTrCbzQ3qbzJ38fA6
hy137F0zfSGSBxUCE3I4GSg2Oh5Z4n0Z9XIAQC7aJtWPp7Zla90aHu1Pdd7A8PycrapAfKl6rCxd
hgvSnZVvATUgWQi9BBDdLwhTTsL6eFjRwj54njdkVo2rcnc6O9JqEoOpQnIYEnB/w4PBCFuYw1Q5
Pw1faAhfM2v3O2leyNeGOCrtJvui/TKK3ciGq/Z+WiXu/FAe9RmoJgk+zElRGcWSMyruuVPuK+fh
rfktBI5y1gMm8W83nUzjgDfabTolMTVzEu/l0NmVTn1R0LhOYq9Fh/Sqw9AfVwM5huL+LjiJIPVE
eA0tFu/ldMtuczLPRtuOZmWKWNBbQjc8dgYw+QZzR27mfC5nyI1uTFb3lIh948CyIoR0pZJ5i2HW
1HlS0UXKl8YpztWC0CWzCeQMOuYh9bO++hXwLz9Ui6ZU2lX+QTlXefkwKhTtTfTarZTl13N+Z7pY
xRkPTrEegy2uNt9mozqYlK4Odeh5jis6jNYcquIAU1aB+WbShhTGGv4EYuppEmjBnAZ3jfUaW0zq
nCH/57mBsuQvwFuw5RW/QQwclAKRWN1xghT/gEPU8NG2H3JK9BFiyoMCh6WQ03MNamDfYjZUzXpW
OyXPDRn6Y1xIZMedMjoKJYrFNEBi2YkYVXr4I0DMLxObeAmlt5JZmY5vzNQ6clwDxlUb9euPVAGA
XS1vUBq1AZtw4wAbOjF74OyFcbwwnNhwmJER9KFj2uOSIis1qj7NvOseV2vXDUcKVooBMHvW/RlG
+TmTOTQA3zbmCV+C63GMbcEftTDRC6s/mcE6NY7NaZcnTXRVDCm9/9MBYp37s+P8J/nEJVJmy7ly
glkVkloWPSWd/0uM5K4iKXIpnYlSQOmas7TGWgDVszaBiPH477BdEm4t5RuxVih7hwjwXA0vZkyW
yEEnGZgyM/4iYTb4Xg9QZ44cJ2XNvBimcJhzHx3hvWYu6SBtjiRx6uKzhXN4pF2qJVi2LFldxbve
8oreEHbvU2dZld0qch9OYGPDoKv/IDlHWLN7y0fbsz5cDMu1JXY1gLBSJZ1vCpctyC0mXsr/7a1+
jh1NgYjHqeL79YlQBT/VhK1BhXjcm+MRggX0AxTHRM24apEX3IJMEGEHIu4hlLO0Y7pPhzVVEUAX
njtVWapTwYD0A/6ioPsenhul4MPuhSCpozxJvSuGGKUMpPp39TXxsR+UMoCKfyU+J+Rd2t4QSXbt
z1OE0SuqyHkbqrT3ZTrr0TpxqeBJDzj10zYv4EWstcIaejd3CUWl/QZMRMvWVpvaPuiTGNhcbG+n
r9YZ8dXYPC8le6zcztwMle8oiF+1k36T+R2pkMkBZ0iFUqilVfJ0Ck9XQtElXDUokVCopAWJJWTT
B9R4yPs85ZkAymEYvCnySVEeyUUDcV8Lp62TDv/XW2u/Lf4Lr/QJhz+zxg6ubtDxqdN8MUAkJ/FC
sXD82Hso7JHv2UBCzmyj/r2A2Ms72snErPrz84pCltNvm7e7VS5wnMWFIk/E9wBW2noTxk2EUZKN
Jx2faPcb+NcEoJXtUNd5QF5/UMG4N0L2/7fFN0rT0trqg0fla/O7j8LucLpAgF0Q7yPlblfgsIZH
S7pho9e83rIKPn9afbDtWo3Ri5Xu5zwo2yGRh1EBcrGTiDzZulx+t4LOgpbC6zzaR/+OO3Pg46FX
/C/5h6X9PN37bewWaYtL+jezLQ6xRa4TwpgyMzmjLl8nwt/b7G0mrvh7wtdEwKTnG5MrmrMqBUv1
yrruwpnDLpl1mQDCCUs/dx4r7E7nh39vOHb2Yo3YoTJsclRTvkCa1iBS8ojC2gSEIpOJaALUXmZx
Fuk6MrjjtZVJa+BtiLfhL/3BgiX+xX9jyZck8AkwkKxP80e3hCx+ihU345vZuwR8rZb/SCFJWPq6
h2bnnGdFvCcqtqJBsT0iiRBJbzSsQpEEm6+HIcAiGoTx1aA/d3q7Syf4TAMmvg0DjAhsTi+W0JuE
7V870CU2cJGfPtzfPzRvWssf6k06lPYQL19LNaTELhVtW1QgZVrDsGtFjzNAGfTE2n8PSJiNX6lN
Tw7SJw0gPXREBmD0kVBZUw8KD0VL2yaheYei8z1wmQNvpKTbkh3bqi0PZPDE8U6wAHLa5fTe7lmg
2XgEPanOiKAuL9N5oWQAGkEGP4rWpYw+kAQw940FmMlF6+D6r4xe8nvA8xQDJDTnvz1DwGRpGaqA
XkQqf5yWNqJ6T1RRR6qfu87XViMJxjf8J+sJ+h2B6qU4UuBglD1z2+BaxwqkzIoCvjPRz2SnFpO8
to7E3u9PClHXPM8CDYy9XFNCTXtOtXvlkJKwktdPY3rMgr/GQg6o00+Q4tVnOFgUb9iTCu3za5uW
6DCkfA9ScQVl0ScAKf7Oz8J11hr1Vb6mz0RjfCdcblCErVS/X9K6SU+yY79HLouGQvZ9SVOj7h5T
mrBXBqpRJIUCUNCxorl+PTjPKyu0F6p0GNE9mcDCdzcbC9L+EDhnP+fCG8DsXFKeg7uw/ouRCtyv
08eyd5w+6s7g1MlQhWwFwArC6jJZk2krDHcYXqqvuFgZa5EJmDBv0DjCuYN1pG+G5xmhS/rnp5Ix
7a8wxEKljq3FCe/nd0N4zrC8YLgBTAJnah3mop2cnfGCHj85z0bRdqi0LZdiTIPHVGLPjtv13N6L
cvRW4TpXacLKHMEtw8xaXZ6tOl6VP3DHgBml0Vt4toOMqGA2s5Th7u/zAbcYIPRxA+djClJNKS6n
nYX1VMiCqZc4BmzQonS3eSsKDVqsqE+3IRoOBOaS14VP0RjCJeCMB8I6dcoPYehR98Wmn6VYqVDz
KWu9Gr8s1UL8vZt44e9QvUbSWDKRZUBjoYeOwhzn4noMy4RF7Bmk5DugaO7PJhZC1BmUYo81TkiP
VAK809Biyla3r8sOd/Tq15Sx6OhzOFW9t/mUnAtrNOJRCgF/GN/+8DFvLl/G1MTe7pO9KUQ97+95
bWvWmayhVeBrSG+Zf9dkT46Hvu8wn6RVSM4Pk0Znc2wVdkBqlSYrXeBY3Lhm4z/DTgnueIMZWGIB
GASqxM+bQ8MYcZyBXafhLLKqo4ShchlkNrGqd++AG4wNuH80VIU1gxAFikU/q8JSU66nUU5gA+fY
mxAgU0ttAMzASYoGkADK4LL+d/XULdrx0I2Tai3AxVxCjdmVOGJI/xsed3MkRWms1Q/6v/2/CJCk
5t/GxmULTxQIobbnC6hAdJERPv/f5KH1xR6IKRG9mQ8GZb0EQP21MPN0uvxdWVKkNbzH+/2jLoYD
DIBLX/7HWWNb9tkR+pxhcpbe9pVAst0ltZsIfBEW7J3JnEzuPaF2FlLR+xrVEN/ImxL9Nx6yqa4Q
6weMCrtnrBwbiwYpaj4gj7zQpbrEd3Y/TIEYFKhbmFuMYiv2m2Ljj45L6IqbpGINhiFHQI/H9ZFQ
lpKLTK8TgZTI6infwMewy/RA0ml78HkFW3S8qPKjqSmvdG/eG2V5FDBvU8NllHaPH9A4BS2ovsI2
DbZRYQ8WN5ggQ/DqfahPvOLtTH2g59fsdSVsg5ndgBL1zTY9FVApEfDoS0u1gGTI16rOUChA2Ulp
azFXkwKwQd0C9/f8XcxIvgE127LXN5sgyHcNoUzpQKib28MY2hMYd9Qpq5JHF8x+df9xu7PelBl6
t64bEv+S1g9IeEmPWU7H2woEMVp3aW5JuMfwdmZrkYSRZBSOnfZEtfkQ/jq7BAE1biVeF4w7R/BG
GT8GNCqlwl7iw93093jaEaBD0UdteeciSdre6DxRtxINOZlFlqxhu6jY1ILa48EyywI9c9+GqBtm
bqJLBLXOJP0LCGodKAVT2UUdp/mf6ixzYjaW0ujPo8e08X+2AJCEhpBTCxPgvyNiOmbzeqcjGBIg
hALMCPDZXGCXwz2yWQF7ZVJDTH//98lzAhH5Ia/KyhZDPg6mY/N4s2Tl+Kct3xyViWbaQAlrKoB8
kQYJ795Ide8XaR2gN8+uF2xHENcumTuYhFrfkm4VUe2JMXAtCuKse/z5aKsjiZ2svCuTMKQTkSNn
Nqw3pu/mv0gycUuUDxQZgGLgHcaWqoEue7Aw1Jr0Om3YQhLG5qDoniJTmKkfgGqRT1zU3jhtIDZS
aR6oPewNkZo9XB1Vd1ZuZNR7ktwinSqu4hD8OUs/7RSAHeMwbRzQeO1+UF3N+JChIAXLszrF7jQZ
wNgKLql7Fll0PMctGMVrFG7qc2398WRXOzeS5KBjLoowONQ7JChL+C2cCSqHh4l7g7zq/lbaFHOD
rRY/niMhGBp3DqhCsAzUWvyGRrsQe9QBHCH7LW1ZnHCJ/MfucbnatmKAD59qBsQtxdIinzfH/qIP
m7mMY2Ds53G6VzHhaMwg5aei3gJ5OZdgCokWmAqM+ttT3vx8ZJ0izNFJbTnMquzH/f44R5QkzSow
IeivlCS/0hgQep+AricC/N0YqCOeoBplJL0+9lKzrRgecZqQQ3zOhMVktheNmDcJQoZUdYJWVP/j
TiQsgdkRJjUXUCL1Uucjj2F0elrMfB3bJTID8MpRdH3tmYZhlabWEBxdioZnMCu9azhMKqOrxxrP
HbXThKHwZ2O6LllmGqycbkt7dDpN2+m2zxq3qWgcKdXMYqScoynusPisY4eCCZ/1AcAjGNU+fuz5
WgUPnMIrVQ/jmi+Z1kd3ZV+lSkasqNdf2cd6Hg4gKIOesh/3Zi4ab8r47GaCfLFAUMG3EWG8S/fJ
JGB44yiBr1dGEas0hferKfYz8anlEcmd/vlAefo8DPxvj2TpZ6BqQjoR5949vWgYp6GF5GbHwL2q
m/vRLCMYyRJWGKh5EAcrKxU+8aMJ9whlAuaMRfSM/eqtawGtiGAwLCsH9JwdeKR7BIDkEII0Bxxp
wbQUf/qQdyNleA9LMR881s5xZrewXJrjdCuUv2PcYSpZ640cVQh6pYg7rYWudb00iQcOky11WOhz
FH3AZ21/xBUXUsejk+qyQLK5xmRBjdWRylgr4PYKwt3fWHKbffHkzh8xuVguXmMOr2KLOidlX+WM
kVqG+/FJTcqQ9ypUlDtIGJVSGVIruO4Y6zoN/Jq8ngBd9drBGYDtnqsnxYjZpLFISUzXEaPvm+vP
9DteMl/03MfW02gwspQrhw0gIJQkFwip+9ipNgmD4yp7wF5G4IGGDrpxUMXH956Ew6/Jo4YwV0Ua
vXgCEe5rVkSF4c2WMsK4mMGbKspJ5Mer6li5aXINwNlABSRqNFhZ/9Wv8gvGoomB5JmFlj0BXAwy
F6ZVjTtl6X1dhU/3j9zpLQ7OWEWDbxnBLesgGSYHEwJEa3088tSaykogHHeYR5He+Dux3bIes199
mGAv9LchTF3jPpOjBedF2WkL+A+0qbwg2tVOmz8q0ZodSJh1HIwJ8u8baAC8+esgUQu7cjx2icgB
F8WuW6qfz1Uk45wi/WcpeEpBFDaXLJHzTYLP5ii7OEGBISPHbHGp3caXWk2HOIbRZ1J03ul4e/3K
7oppyX411yk0+qRjye0lcMp2iTpR8BA2D1ydMS7BiKSJoHSDR0UcqlSjM4VENJaVEVJ28oilF6rf
ccnX29wZczDIqDu9VCwZ2QoVBW5IPg+4vdcBJnPj7uIrh1kiLU8tkasQLVv+RDIvMwuYHuchMPWb
AEG8H6p0E06uODVV2zK/wpfkoJv0prFmblMV6lTEfEyMGRzCEOil0MF6xMPxmmJn1and/H+68XsP
yXxaJPv1WOvbdWBTlZMV+fakTSXrTqgsSXKTO9CG/eXpzzYklZdGS7ThOHav9sqJUpx5s5hmTVYW
Zv7rQqp4aPTOa0GBF34m7xV0wgpx8o5hlrh/NtNaeUIWj4zif5zfN/3RTeQltNW2iHuN0Tq2VH6j
5NKQ4lMG3vYvONUfeQrymUN2FCwbujHKau83hP7WHmQ0EofNKOdFkQVVSawn1UNHZO9N1DFHRyyS
O/G4e7wrij2Q21iGGseZrW3wjyKhSebXP/1Y4VJWO/ChWKahDxk8/nO88f1D6qThR/16bVfADqmg
f5FpgSosQhQUL9ZjpEFSdmfoU0pIm5Qm49Z3VkEfDNxxjd4PF6Z2FkkSQhUzxc5I8NlScEE3TNHD
1LYFoxRQHoUvDURIZXbnei1VUmxityDJfnXQ1pV66KHfyKp+Zjbq/JUIQTTXgGDVpl004feoIp1N
pZnohPRqkcXD/hsSJfkTVrfzNeZgggFfgWF3UVk2wUEUYAOzVS6VMA5k6bSl5qLE6G4SPUj7p7VJ
f99mQbj50FU/rLttFtYKUs37tSXAxIF0kGTExREzzLM2DwElvZ888GJ95pk8ASMIl2eODDdK7evS
M+Ra2P0C2g9kuwSnD4M0ME/SvDN/rEwX1zLPRMhzbOm7s8F9sDP56kau27o8tq2h4NY4QJ1KB231
wlZ22PcixX1JVNfa3Y5rEw4QhwEu/MBOOZd+gX89GQGgwRvuSTk0EkXEPQfkM89d2SDMKvr21LLJ
fpgYRrgQ2Np9MaJ+u2YHZ8UG655jCzHNQZcTfgTPk5ZyArTi/dWlOf8DWlaxIDLhfgJXQvLYp4BQ
390K6/uiWt2+N3Fc6AExPDIB2PqHjbLViTWQNIcWCiYWQXRze4WWNf28X4qoRUyWHPwv0h3gKvy4
KJMvoP+lqvL17RpEsFTpRvrzlhKafaKXR+/DW4twRnFC7xSEIdcxD9BFzwGCzZS6S2M64Vz9oTeV
pKoXGdbmVc4n/C3O1a1Ycufuinei1/HpaaUO0EWDkc7FcikOofDvTvx93AN6k5nMO8+R/+lDuyBC
myDPW5QDFRTiVwGQpnTlP8R2SDTqZ3Mr67Cpbwt8Rf4oCpkAQefGVrUzp9xkVFT33RgQCPDwAKhk
naVtHcPumOYNrv6Gqvg/V/70IuXC5ya5eYf+qdWwl58FsEakKWguNf4xcQxRn3VfzeqrG5tcrybM
TIYUo++DSDwlJLp+vp+BZka2FCn3cYe+At5zIrxkpl47sjVkIBF+1jAesu5Eq8UQy3w7G8x1RU0i
U2byUYKuyXJI8RrTRtZ2mpVxZyHaHXuoFPCVYAAoWrOVmyf6vlTpKkJx4JirrlF+L6QStMECw9YM
G6gJXMoUQHbuI7jNwrCGjueLMgYOOqe6R9wQbgvW/l7fu0u5UAxP8gP6C48vuymUGT7A+BzQCU3E
jE0C0em+ls+dWpGGID061nlI1/ImRmvMkFDOeXo/laHuckNd3VQLfrGI4i5lm2ioRSXbqkCKEcOL
qKar9owAf3JwqNtXatmtsMNpR2nKJ3slT2sbJM8c3YxmD5Q7SwX4BDcBb1EpgwE/gMpEaor/b8tD
kLklS0sGNGanJSC9zM5Q14dDFXq3tQvoUXN6wFhzh92dH9OV1QRzLd02gF1/MdOFbiCqKxcq6U4R
heEXh9XqIGQY82aq72uRQFugk2gmhZ/A9fGu+UUQelo9UhbhFQrjQn08+mcwZkJBhPey9fMaVHqh
X3XB3qQMIOkw5CFzmdnuvrFeHxgFsmf3vDm+346Xg0EHT7cZhI7XjXDb6UAlVzLtff5+o27uQd39
Eu6ovqZm2nF4g0crr+mSzWvIxJ918A//5Alp110nGVgPiSe1/f3sxDud/8D3f18MizZZvBvFl2GT
OAMeUgv4K4wpv6P3UwN56Gskq2JVn6pTraVhqgvkrVX70M46liT3qa2F1cLatlDjefNAcT0AzR98
haY+IwxPIia5f9XziuYvTueYYuOBqkUeVh4DAwt3K+exm5e3p1XayV2ImxoSXHpVZR12JF5J/8dV
uDBjaXF6oiUG4uAltODA8RAGXtVHab4kZ7+6C5YdjjzKut28zEAj3UMOmlAVBRbCVDU593S5+Ojw
a94qI2MrOxQh2CWpRj74mbH30pPjcnqDVxr7ZpSsLX51sWHcdzMA2dWCe/94W4vf1SzWG9Bjwf7G
iaFdWXmvhg0FSoPOIRgiencibubKH8q5MYidjp6COfOYCa4t2/yyC4qd/q1qJqjgwQBgZs3Zocb8
cShS3mCRFLT9kqE1FLPTXY3Tws1M24VrC4vs77vZ71A+7XOKtD9VAwGMsDI9SDpI3mjXhFGlUEdy
XrZR8i1xHxDSa8B6lyDVuys0KB85i5Q6pwiU9fCgBSb7Uhvw+8WY+gBiPxE1XGpNnxjXpmYtzJqF
4L0dRZGn+PCzDoxl89I56DeHKSTX+N5++r7rR6stEI/dT7hD8NejDA5PkmLmDnbQ/b1Xb6RPxflw
a2YFk/0XvdQTnl5Zm5wYbKfIdafx2IdoQn5XsrX8MpxryRnnX/tG9znr9L6uBpo6b4YICGOceDhK
n9AAZLCWlNxjsH1bu6DQ5tzmjx5h2wkV7r6s2T7vDZ3XH1eNch57ivhUfEC3kQCIc58xqsLkMNWb
hC5v9ChQzsX45SihB6Ka/eOfxSlQ6FOoKcoRLUP8ReNZulFHK2yWNCRjsILESsUVvpZAoVcKLxk8
QQJjrGbEZBLBKSDdJAriDRk4NRraA/92eysUOJA6GEOBV1+06hgYRBqueokZKKaANwcBrdLH0+R3
VA984YtGE5YPmUajSVZIJSQSwxc762qUxW36CtDl+Cj2a8q0QHb9uQ8B/FPFTznxrgs525xP77xl
WB8YmJcyQGnUDvuxefqTCBXJjtTAZPPUS7eYfB2PW8gdwxrWoCnu1mFpE36pJWpPbcEjhfH/qV59
nh2duC8F857hXt1NCwjyUfgbXkQrM7BWY3YmRZxVSPBro6lVEcdZ4tB14vM3TpVyu18wCOLAz5ot
Mrm5aClPAKGkgBygGZkgJRnWeI8oCH1NZOwbOTQEhyAS8MjBYgQbCVMywymf8h8XaQPc612aUBJs
IrTkbediGvii1gZrxSP1TY4fiIistvrkWoCEpcBwOLCKY1Rtb+eHDaU9RI3rTGFEi/fc3g2hTUXC
0ei5TgacQ8QCqOd1uQ/FC9BJsOe7vwnAWiL9RvfsuCRZAOys5VGtNrjjlzYe3dVpoC6b/Uu9A8I3
BI3H1iEVu8L342+2nx+mXafE8Hn8kZfNw98fW9cm2wszcqEZscSGun6BVeCFlHKah5hj6OgcDJz/
GGaaY/aNDJhi+GgK2tofbRlI67MeFocdlaWvErxOnweQuwPNigxBgLwQF+bQXCkGw0BsD1LS+gEY
uioEN9pPRi6KzZtueQjG1MBRDHTywyOEPVaMSNhjzac9KIpNpFLTaDquEdB7JKuvdAO16BxetstD
wdFgRbkSBT8twfhxOAx6fOA1vVAiic9MPTnYWflmuKA1QNMaijvO1l7TsRvQrxy2jaOBivnUbwz6
3QMFdm8i8zPyg5enPTeNKX2fc0N/oj2PjRVZJm4Marjp+2WoWRBTGygV34Q1ol2qEmvKhIcIgRQL
/bsXKWq5E0BEoHObHrEwOq5lX1GLoAXhuvPaeJK+sVnUh1eDtMycyTFk6qkkOkMNSb0PQRwa3+vS
DZmwR7X/6Dv8yhseyzjI1ChVAskXXfSRXMw5GuY1aV2PDamc+P+zKwOvtS0EBvfFogR6vHgJXndh
k9KxuHinRWd1YvMaBPSENpI0BuzPZUdayAwMr9SIIvpzrsQBJ1wYkTidtoBOc3/E/CUVNV+GbwtT
xe8OyIxVm5V2o7Fod7tSJV9i6Mh80Ktd4kw+3AXmSkUSC+79U3NX224uotVhEKwP/qE/rtpA+4WK
dTVuscpieMO/x5U2S7BOBde1V0kt5iCrb1zSgpxN5FQPRPAB3v3X2+fPke5F81PWHqbYAJjUSs4o
JtZQO07ki3GEGuEeYD6goy6sadxMN909kZTjgdGHfFV0rob8PWTGaYoGql7wgVhdBHhzLR4t9LQN
fjtzW9en03Sj/Jl5MmKwrWGQuhnHm3eqRxCVsPOFVcE5ibMDZ8ytAfSWFRxCqAsFD572gdF9MTFa
DBonhB8SsWYCaCjYDDVszmrrmKEflH0zvVtATWkLidp4gVCDO+hzRnbD15zzP6JlEMpF+aUawjeS
jNX/dKINwsXetRAFNhudLEq7ZxER65QO/gHf+nSONKCMzEv2D5lnYcTFDLzyX8ENi0CfI/F4rGpv
GTlrGXooiFKGnNtYGrvPfhErld/VNQpYAsdDcItulspg9Ms0rToz4lYMl20OtORDot+aE+Q+fRVH
CVVX87tChtNonWpFuoyuiwerrwYM1tWIEhAfwnbq52UY5x5OBPb2D7xISca3OvgT8vXziBU1xnJu
ywxtIlyGB5K1BsnEkpwbtsINNcsKyRKY7/rDx+DgTyO65cjCoKl+xdJMYxTp+1wC9ho1G1ola/0l
ghOrKLOQN3IYgKfdFMJeg1jJlPzeRwhEN9dXwxz8702+wtiV24FWIDq95q4dWOJRcry3spZn/L+v
uH3Fk416XOTUCr+x8AIDD4VlaSvQYGIb4gYDaB4HEvGFOx2UQrHgL+XTsq0iEKyrSvUGvocw8NkY
RfVyi+6UfYaFNQaD8sb4glEtsHHePdqTD6wl7MEg5y7yv+GiQoPoHdrSIcOC+1xflK6qoWjC9CmV
TM3ibUBlT8wOBrv9RVGug8wjaWcrQKBIVY4++qqdDT8XHltt6+oJKjREzZ0qXWEhRZiNbzR9kIE3
G8LVI/2F2A8NkG2N9uCf6XImGUzBveQpGT7QYVmPl/eo7B5UrGryOS9lOk/3Gv4QhqQnTK1Bcwoy
oXWjuS1n8UEX/2OWxX60mTFJ2YS1xJFpvIQMORT4Z39Ip90mWmoS+y/1mtFa4YOrxl7WDVpiKWFm
KvQOmQiXMB/G9LFTHO2x3rCo5NtsDaZac6UDAMY2kAezg3uQxTwIHzkWRtqVRWdhpX+/eWoVbRnZ
EWVq3n44ajfqoJJXDhjACc0adbWZKyWiO3glnZiYt87t1Ezd6Ecd2h/fn/rgOzA3tXuVUEioMdiV
OXklEun8bGxWxjeoMPZukgNxKcSvSiXTbv8SkqeNNxFlUhe6kmo8lFZobxm+M+a9fLSlS8ls2uCC
PYHd7U0xhq33nLTaWdLE9eZX+Q5jvj+TgVSUxSVypfyWK/dw6/q4IrHZyIWYEJ31C7DT8EmKc4L6
G10tYF8aYzyN0Ip2QHY/A+OyAPVrZSQV6YeCWdGXLxwVrGmct834SkvWR7LASumvtqTdi82Xmdck
A+PxOR3jeJJssTvwlOHLhNe/qwoV0qONhMYbt+MfJ/CgCX+z8QgNuJ+ccuaeCyy4Opdsc23tZrL3
xmNi0FCNhH6PzoF2GtF6yyG0aA0E4jREd7s8RT7R5qM2tj6AR5yLFDCe3N8CE63n4GqT97qDlU0K
gSFY49vMRw2YVj/LADMwSWIXO8PnFgkCX25ocSuiWcBGKwEMHS2wPUddYi8ny//SJ43SOnvyArZm
Gf1FI/Iby4cueT3jtGDeQ0tjHCr6TF8dnp6uMI/UFiDcGGR/Xap16+6N/n36N1lyI6TaLp03Wy9v
9+yJYSUFTPO3ZURsaGJ5wDQiTdgSki1yGWyWqRAev5cF3vDgkYWklaSV/rmwA4EZYX9BIxkL0G7S
4UxcbF/FeRlMtcEj7AeRF4xutzR2mEtJtl2u79hvvCX/wtfz56wztkBEGDqE9TuZbPkNRz7k1x31
hlO2ccUvCdYK20cFEnoMw8sHF7x+ykiVlinbUGkudsDKGi8rt+h4fki6s5R+e9qVByB13mnzgo9W
x9rit8IBOKeAQedYH/8o9Y34mYM78uQhpfFcqcWUdh2rN+NgjfvAGtyVGBDlfzUwETxnuO/7ek2/
lNvrAbGIhlIGsgkMW2Ueg9lPXqZ+h1qr3yq9By9Mm554LwaAcu3UdFHGIwMxds1KxpalasuCCrFj
iDTC0Av+R/6rGsHHOcHjf4t5Lur/2mcA5LVCdQIrCu7FeGc+bi1NpiL7rkFXXeCQFQPYrovp6GOx
pwoJTeVZVhJw/1WDAp8vZYjfBZDLXFbrIpxL13wxVBsWT40o7Ei3rp/MRsn9hKJHJp5WI7MU+gIK
QaE2OYkSXHcCc2HZV8YsWcls2rYnyO/CXQkS3QE6avC+M/EcaKXvy7oTL8GTF5kfFZ73khQpAFhh
ZXjoWP0+kObibNXd35ajoIDZQIxuHeMUjPJcTQsKWKCfW8xqRIJElq2e5P+ZZoPenqBxE8o6viiU
wAu1qn5a04++55CubbVakIBXU6zo8lE7auHUhcyJSGAhPEpZRB9G4PxvVy6GVMw0jLIdEgPXGoaF
VwKjZrT4sysrwG6GX6Thku11BMTLjrYxmWzeWXDkwPUahO+yX1Vol1bdTppEtCI+0vU01eCUaQ8G
t2FyRa58JqaLX6Ns+l5DGz7OS++b/7KWMgE5SHyBgJjgmmm6T8ZbNa7j5awyA8WL/EbCJ15FI6Sx
Y1NmznC4ouL9koF8XD5XmIacZUPouSBI+4/jJ+3WH8aj6ieDfz32hU0PwBp+6mzRTsnR9jd5yN1X
8Fl3fbEuU4PdQkI4mvXqzuEJNGW86lSzXNT17r6xFOGnuWSVCueALdEMxRto3x64yEBqtxnniVsx
xu8eX0wZvFhX1ScIFc3VvDMKNogkPGCjaevMpIGv/9LTYlCu7sbqMGrSnMNhBOh+4vJkHsA/0E2c
TwkGtJfqYSJKpVJ73UiEDaMdoJA8ba8oq05tXBFi0YIgsO4JWVYFWgMAI7PQO9NI+2RQkHW04heN
Ch2fRBorriyewWbTRnBKZECfbcFKqk46EXnovy0iemHvJzfJYWZ6cDw3TsrIMZPQoIC5SIxCB0sv
wGObPF1IFCUhRZLOscyTgQvBnGEBvvC54KYas94d9+/Qnu78bOsTtB0BddDDZWU2qWm0c4KP+mhY
E3bIFyznd1dGPNJHfsP9CuR1LADQ4ngXpQe/BclVKea53JVZlLECL5lRAxp0lqysptTKEuUqOM54
TxQKsh6dMu15sFEHjrOrICOx49txFhgEUEvrXzg1/azCO1rOldsq8Mnm+Zvy38ZJehMS80EA9FgD
CFa5LjyGtBvx4EHHhcBmWukloQOBg9e8A0sMmyi1hGxbFW1pPx2+go6tzUx1k+SbtIXGokrOKbbI
qLc3bEmFgI2YIgmqujcrulvw7iNRHRswqMYqhxuCovnhrPTYfbUSdSpXuVid6yh/KS5pwL4Ozs4P
4m4rgquFy1NhzR3IYWHWNkfgwKzxYtU+DgyDSkucrkuCyIcVb95W4HMFquxHTfci/2uPvlt7g/nd
8vBZrvBx21rIAy0r0zw+iF9ODfNxrUT+5OMKogXItguQBkSGi9tL3tuVeKvl8vmF+IAoCznWQ/aS
66nNXSWW64y9x1eZj/Eab2yigfHOwpCUJq0kBNV3hdXRWRooXK/XxldEhP13gyjOxq8I6kZGxg+z
7vogpvTJK27EcmZRYJH2qkIXm6G+DHpkF9tzq8zDjxa7bhvNLWf+74r1n2WHokfi/Z95ulSQ3Rst
SAawabEA6zd5G2p+P+HePQZPtbEbA9Wvp6mCg3K9k5cVdU1gz6/7wZL/VX8M7RPqs7nVpb7AwFM6
gUulIO1zemYceQZjviXAI14UD0a1Uh+gH2wuWoOjgVFRLURfRZV31SUshxrA0/oJBQA94t+C4Un2
287tuHo5jvDkl8IUDul0KDAvQVDdRGEwFm7jngi0LlF4i+vO9cnO/8S2iPavAFHGA1zP659vok35
muxlc3NG56hCFf5zCgmuL8BRNO2HKQdE4zHGgHqj49DmoHWlaG2i16DR6YxSDY6bPmSjfhFSIVqJ
FqgZJ3WYXBZcxagH1kp9ukoLbzs+T+ioVuZ7/fjpaxMttbcYU03ExuOh+faNssWCvSYioCojTvCG
v/H7l5eUuROdKy3E4NB0thbh2ALBXAEc0P87Z//vG9oJN6CjQW/MzxhSVQ3ULMauOneljhpCf0q0
YKDAR6TFVO/W35q8KKMrw08m/2zbSbuhuKpOFNWO4WVylsKHJWilpfHBOHUpgZ59haXBaRZnGTbr
B+kRGkiVZHp7sZ55gOV7iNqG9SnbTJNogjQE8LlDa0zhKcOIgZCEZf/Lbd32LaHqJPBeXbgkzbMZ
V4pwi/xlzoxjgxQ337Yu0eR06WvgQPyzay/w29dBitiDh5x9Jp/f/ps/M0bXm3A/U8t0Z82LBqdO
sxUAipF1NPCZcnU+uT5pdiuaRQFMuOob7rRoebW1/7oteh2N914zaW/Gh6l4PRdGFp9hM2n3ysO6
g6FRe0HwOr4GB8hR32L8yayFcfYC67fHMeHr66jI74VAg6p8LUT+mnIFsL4DCerh3BNhX2W0HeEU
01vPAPbvWC4EnYoQHaikHkoTQaMJkk7MAsQKkepihZJCW9e7G35jPsju88sCPkhXYD2lNr9cbbVg
pfd2YSP/qi4itTRWUh5nRu4NIKqaXEZQuQ+2jJtVeraMku7Qpg8ttXvNT16sJ9XHpMQSVHLAY+5o
HxsbUpHkHb3AGqPyNG2BP4RoXITgwugTxVSSTC4bgYtgvSehXuBkc3tc2j703cklMKHKqwB/GO42
T53OQfdQGuxddqiq3YdDnC149uRCWQKMK2FbwQ6EPAFzHbbX4Bg+xJkZxytCBTGgNNbaViN22L8d
JMOaVQpRN4+J3hanZhvLfoavA/w+Qi6fjQmjT1ntwz11vq4tHFQ8MPGyeej/QjwFH4gbnvBkCO+O
M/JZew4riAVxO1kzaCDxfKRYqWpfQoxmliihkYR4M9OLNqzBrcQAW7aEB/Gq9hG4gk95djYwSDFr
yqOiopx9eToK4j8ikehSNqN4001XPQ5KrI9/4oH9cG3kgWZv1jDs7TQe7Ye1JE3M39nCP4p2ngtv
fQF7IUaJfsib5fb+t4dnZE/2kTBCOEtCgs/hj089nrlDn1iQovJx9/R+kTVqVjF9bbq/nWOJ5cCV
ulMQksceuaCb7wuIbsCScYcn73q6I21IQdBJtrnKGemhqOrm36D2iNXuYDvkEt2xIILvA4PVdLSS
iRiWRBrXke7jrhxKORrCMGKzulnb8AtOypEuuCSYVvaqM/u25Hgd72rkmfRVuKKp6NJ2XjHGZuR3
C1WsEBlhxsiaRCHwRN2pPHDyBxTBf3Z62/3FVcZ9GQJxtFdOFTiHDbUhwVp1TnYe5XhAytMiNnAU
C/v64dVKHFHEgyb6qU/69aJvdVHL0KjcVx7afapbhetPMqkg7znemxjnGycRSG/bXzZWcmPsJ4Ws
QU8fUYvKD5SJCQ66Zxl20kePB+9dct/NyJsKr50Bncyp7rH7iDaKJcm1myBuM7BXNSBGCaHFfXlr
tNOsEeyXJZvZk9BftVYEqhlY24HY/tjcrnouFL9HoLrWd2tTSsJl4/J4m9Xy5/C5TvpD95YQNYGb
3fg6Tk36Mlz14SiZjMLg1Zw3cIKVnbPhuLJJ0+n7fdDEiO0EzKItP8t0Q3is8MMDONK7TxcKbmuG
QuxNvVUx7kXPCjqusmEiKnL6seyjsYwd236S7TNfIsXY7W+HV0Cdcc7ht6shbxyf9qBdIa1e7K0z
0kW34Qjqbc1/JT1bHfJ/GsjLrAOJBAUVSX5yGK1soybVIo4Jt1Jr/Eswf5EJcer/MovbzzXjl0yn
z++H239x0BbtwR+K+BQghS0bf/XA4SMTnOp6L3ZlFGivz0RpM5IcmKijdyGiJf6Wg2xySng1UzzX
3c3Gsd7zETvTCsQFIR0Pvv0DapdhOiMCW70W09F1lnZ8Afdt0hsoMsCrZzalBQmg1YdPAn15nGtK
3MWYgMeVPoS0VYXygDEWpte0hXZnXF2ayGguATzJwA4JIMYUuxDVySJa3sd5ng/KCwNuh1ghweL9
+upciq56eDbPLdkWUj3uukc46lh0qGp3mhHyrLbhXxAgDKeyo7UJ0hDsmw9ZYAxYUmdcn7MAxCqz
98LlLLivR96WU1Ch6dpqmyoEr2DS7lSGlv2e91+XYSIaNsLnwGtYEaWeoOFhJrtmF3kbsxtDpR57
gTc01YUQ1FXpBbwwrXt1K6zSkkTkST5OhPWLC3WFMygjGbRP40aNGIrmQy3Nmng238Pyienmhwae
ocyzWAH4Z7roVWMiw2Md0DeBELTrbNXLflWERk/OgUGf8t0hwfXI5SCRmQS3yWDb/dy6oKupxxpm
Ywz94tb+uoSjATIc0wpiScnnc0vjQtswh2CcvkD+0EfFyAC/zgpmnbmj/kDW4w+tgVUoMnsRDNpn
/Q1iXbHI0gaUSCPp2thcD5u492xJhBdUEC1WgQTNLTVDCA/o3p9RVDZnVl0GVhJlTp4MUi+4BBdn
Kb/AtcW3tNFwnncnkyflUroXsJiYC2NptCxXhKGLKcmb9wclLuK/86LNgEn/rf8w1LqjPyO3soKa
8fcck9bmMsSML29d44VlD5Q8nNxfKLnr7gI4opXMvz9lM2P/Ru8bw+oZnSOmKeLP3R9Fq5RiIqjg
cHCdPoZQhm4h9fiD5wSOpZlhK4FWgePzyuTj7noLgxJA34oXrldb9reipdqn67ZfZ8kB6uFK3Eo8
7QP30YW5Ls0Ak/rlzITcg2SHKnWQxbqwgsCtzyLn0Euao9mPs7b65EjDyys4wJKJgPCZCrcdxf/g
Iq6KHH63eO11YfHRNmE6PH/hiFBVZXdIMVIJ9/M3cwSF3/oVTZn594v+4DnnuIf/cmsuaXHqUP2U
fDxotsWxXzy8mRohAqDNhS/ah9k22eCYi7I8pa1NEiup9uAOXlwuvr0Alzp3AuHCQsCGqaj5e9YH
Dbik+emfpXoRRiXtQHGb3GlvM7EQmIt4LnMdPfMQ1MDMo2ry7SM+aegANCufwgYI6JKAQ47X79IL
D38rmsaz1KBUrf/NmBGkth4DwjfOO9RlV9j9WX61ugJRHyUOOkKhLf0FHPh0F1Gfz1NJG+0EYZRb
lDkWkSVQPIZYTWxEwmJFs3SN49eb24/u5HOpGBVTTTcm95KYiv9MpZFeE2tcjE+zBFCAA9su1jq7
GxGaYoQtGxhji3sO3wvMSjwzyCvhbSSjvz0ubVAtgEQh6xUb7HvLZww+JzRTwx5CCylHDyyTvPYl
haAHXrxpu8T/6ybNQRbtllNa3u7amSoMl8tdFTmeX9eZ7cc/TEYfHAxdVxuYmxTKwWgDzu8kgXwq
V5WXzPl+n97izLEClF6XYnfbX/ICP7vVOU3eML8HYjltL5lBqhTSUGqSdbYfH2CWKJyGWV1b1vNe
qMGY0gqyJGPxOQ/KeZOJY2rxY64AOb6QLhFXei5s7KaPl6kdvnWHSyi5ebg9SV5TzmaOxCVy2Q5X
5TgQTVC0xoYAw7DtlldLBX+O3EldN8xWbSVpydqqofgWImzGOTq01n9p3y6aRvaPk/C7TDIrcqp2
8KBbWdrn79GgsymX0XzYC3ljNFJrHJTZ2zAo/wPje3tkNnCsZdGTpjyNy6AlViB8azz5eTLgxfoe
3GPRP48fxVkc2zzkskPDlOrTsc1kR2GIaoDWv/FUsJG0qjmLuk9czAqVEckfx4HckFcub4UoMwDi
OtU4/vWeJBZvFC625a0dpVRPfkkqk8aJyRLUU9Z6XgrXvZvqKvjsa2zJu+olfNjBOCGsq0AZUjtr
uPmSPL3FgKQ2sP0R1cmw/BUF7N3+meKeYkButOt0rBuKlhxsz3LtNMd9vKXQs3s41fKVsFcTr9jm
InARSyOsLgChxBXWoM4LRkbao0NKd0hRzCqXzO0lbGrGUth933dIO89EP3nM0qvSwUzN/IoqTahn
83OlRBfV7x57/ZPKUxRRGK2Kttc8B8N9FlUBi5LR4jt/DGTHrOIeP9Xj1Hmcq+7usuC28v3W2yXq
bVkK3QQOTFZzVkj2/wK4KtdkvtucmpHg6pk6pyZDWYDCJ7Ky2lLZFHmR9OvoeOSnq+CK9gdvM/tV
4pgJP9sSR7jwCrkJd/cSW2UyPk8/O3+yOSMNo7o2xPITxlPoUsxm9ceC0O68GXAvERZQr+pHfU11
VDJiP6UK4w4M9VHspLlje96SHl3E9MkB55DwIuq7DhkYkZB2dboYpwgka8F+MNueO3ALe/3q5Yct
z5rOVKiOBhSFT3alTJR136fZsnrQkhheiKX+p+AyCsr0PdNy2ihvx9etuyWj8V7DPHmYRQRz3d/Q
OaxSRZ1vo7k2ZNE4pP2CbmatvSsK+ym0ZNvkIiLDgGu4lbMkxhdTLYx+xkPIPHwI9FvJTEfBEGRl
ZjWJzSp+KEoUj5mpE68w1VoijF6RHTa95r+FU9z4SVgWyajDDFM21dYzGhIFLxeqWbAjLhVxdZtd
GCy13CDOq6v0eE2BfBpfor2QXAkvMyrrVgxOk2eWUIfS9GtIy+CXr6uNvCsGWvLRPaazIpKI7cv9
aADmbZm864e0j289JN+r0CYvKuY/FCM97ETdzBBWbma6w3/3/YOCdJ4oLrk2idqiV5MrCueOES6j
3aDjilZSCGTVT+TWbltJhfZS9k0CUk3cCNG/KKVxIDmw3hv1P00pAd04wPts1Eg0UGtErzTyojXn
0u+XO05sB8efvLa36WZ9KJba3Cuy6jEctFkP4+bwCVg8haL4ycKqU8EODRxZgAcll+hYWpahGDnR
EUt6GQrxiw0a2xW7e9JaAWPerq2dRoVft0QzrGc3nSkmuag8GOZ3P09Ujdt6+m8KsbIl4r7nkGSC
s6BAAWbCSCc5J2j729bjJv9fpeE8H7vUJSZcM6tNhr6glueW34DG7DLU6Z5uKfCdM2ITfXATj33o
Uw+m78Vvk/y+ixXpI227Ql9UTk7jmK4iF8l6igs+ipCeUmj9upmTj9Hm7JUbcxek22Yzld72jV19
8n9Bly2eZdWFgPpU2SqtVY7LmI7mQ18z2OgwabWVC+5KTRF2f//Eo1sB+B83mIEhXqXd0XPzs/ih
Gr0gfSR9eU7M63fbuw7U4wtQZLa28gioAThw72mhEPbBZRQ0NPGj3SqKKJnJHlRmzwSHSzO49Elj
fpBytwbM4PD4VQFwSn6U65aWhPllJZx6ndbEjPeP+YNNAhrSgMn9ofM2vPYSP/JTmTBCsFJbaVJd
jW2R0XA5c5xzrnsMbxTsD8MJyqnNEJaCLLQDg+P2yzksfbuWhtmh1S8JuK4wJm+TwptUk5UXBeEJ
fU3g6Y60B0WD+YfgeYFy12a6Aco1d9/JLv+wryapIE6gKDFVR2TtFpxXXZJabVyxDAGhW7WZoo6y
csGTYrrCX1RGTJdmZyz1OiJif4i6Xb7cGSmpm0N7x3GYFdClWAdVqCDJAsBUa8hYbMkqUbXYxKv0
d6nWYl2OOFYcxZVXU/bFm3VBLUm8U1qEVDfCfi7L1iNL5kLVcqsURHwBWB6dZSwJ2+dJK5/1RD9c
/yLhxv9eth5GOEReIpi5onP3gQvFQ4LauoBMm/+oUYMc6GM3tD9n7P8iLfXtBpR8etcElvBFkio3
I5VVOHGKj+7/gGnkEiFCaxAGkptZq6Q7Dpl/lvjElRhbdIcocg5P6ljHazOzHhTDtnxwva/r8o69
0DwxOSBWqKLI717kmKvemjdMR9n2ogsltEFq5JdR+krJ934kniHHSpaS6vBYiDR9ubrRGPIq5a5R
A6TOlR32fiHwJFm0pU/uIFXM9fyNs9h7isSyyHnky2ocTgLQ42tuy8AZi416yICqlgh7icRPS2iR
L4nIw1AKj4xYtY18mnjCdIegLGbcJzkP9HeT62qAo1yiqqTYU80u3qji0prF5rPyr35boD7d875E
r6s/6L0jvgHs5uOGzKFKhXUdytpJ669IyljbjTZ4YWfrkn+xcBprD+d0VTgaVKQc3KWU41YJEL1s
DLcjSeJBungb/kIl2FqlYpFJxbJxZAAxnFqH4RXbfSm2AIPuBd7mL93HwkZ5UJC5PgR7DAykJWF/
tUYHwkUByNV5r6E1zLOWBYqwvUETw1NPBg1vezgzr2ejzhzOebK+smZb8WGU5KS9U2ffkxT77Wz8
Oz+92NnYz9RZ4NS0rnpH6zO4yWYwPmBGDUGfJsOmyJYhkKRV6TohXZnKJzSouCUSmgk8RiYGGn4o
K9JZZ87laxBJegMWsAfceBayW5/UzxV1uXi/k/tMfQ+SL2LbXdWy2XvjU6PXwJugRu+wl7IRNGH/
wzANQrckoPmYfVRN/gsrMBzKvjvVDZky/dHkueUv5mh4ign4KEIIzyyj6vecFXoP06wcMpp691t/
S9rLttCM6L3+DJ9K5txg6/X++lDeTJXKSF/pBUWHL1D7UogWzkqke6x9xIa33JS3NgvaGnnZTtvX
a/bqRgyvy+epCw7XZ1mBS3OhRzehf4j4CX23DRAFWgcv38JhyOjUNkZnkBJSvYo9MT7+1PTHjIcZ
nTz0JWZlExinnjGenKLp+onv26M3LcvAHMIJkibcL3WlXuAgkhrTtlCgooLB+nWUu1WMgWY/NYD+
0uCyG8WlIxeaAd01d7h1z/3GsVZf/DRzsvGNhN+eUC8Ib0axbKMHi0f0wFsFjljfx2Bp+xvVOMcd
DkgzyhYiKNCq1Uh42cvrCamo5KkYDF+EWTSAMOGeMVv7O158+yby2Dx/ti9+RXIt9SNxbinka1vy
AoEsJn0EkzHjZhiAl9ByAdxwh4InkiyvjTmAEWUvIvcBUB+pgpH3WHYlx1z/630KbkEUC7z3KQeZ
ARlV2TgcBz7guXUM26ykDZRPnN5MkvbpGNQXw/JxSRIy4gwyq4SXcXmZj1PyXPm1yIpcMygZdwNQ
RYxKut4gY0hOBAbpK28KQC3rC0uewZZfxYARtTWck/CvRaiJQOunIjPU13kq4fyeniE2H+phqhsC
b3879xJoCGoPKov9DjmEiw9oUzacuGDIV+RZjnW5ALm2BqbqwZ/8T7kBy61Mhx/5CE/HMbZdJcKF
hBZlwd9+2n/tw497jbwmY7ek83U2/FwlTXmRE9MkbBwnAYJTOrVHK3dPFNC5QiLUI+XXei5Og+du
wqhkXkgIjju8tldbcEOWveKJiGC1a2OzkGBWHCfENtw3ItFAr3IEosbWu+vXqPG/9D5CFR27VdA/
BMc+oGqTi3SpcpUZv9ZTHPq9DPH+GV1fhQdgR47LT/tMn5x3+hBKuBat7nLu0rRNlRoO5hSwNNpR
ndpvPXQwttFD64yUg9grVWYSz4qY8Z75EXfj0SaKbS6nC5hcuOZ9ZALnrE57mSuZcwrF4FY/LNTw
RbrFhJZLtrIB+L2Us99akanxPI9Wep4rMThuAY4U7dnBCHS45hxQuD+3pxfEecPz7bIE4UDmwM20
kAfERff5Mesv1hsjb9tHc9yH/TYcI5i3T5/gVlt/S3HaQacCd8V3yrGTOMkFDxepKhSj21wtTbJB
jnmPv8lw3CDx2NflZEPDbV7mvFlmFm8ScqzzaFxGhcQKJQmsKYoHmKLr6PT3s3g8VfSKef7gvHHO
hzllopxOgtkGhdt2kxFoXAXLZeiJoy2iY88xyzDFcm2tH8xfFdfEkwjL5Xasquz7O/wrzde3mR21
LIqFpJusRA6IaZ/SlzvJdYGua6WXiVkL0yI7BVe1ls+F/WHTUsYBkIFXaPcP/9HoYzYwQ1GSkbLB
uwdDeuAOKFty7SYUoP5sJEHwO0qPPJkTGfsPWri9AhS9nDOVfR/n3Fox/eKys+TBVmBKXfxIWCKf
via6FkoofHuvBuvBrCqc1im3/Pa/N7ySekZxJv/ZRkfI+ubmumJQgg4ow/gOcG5J43JsYEtH4hZ+
T8D+6ziqwvNb6x8PCKUvNjY+Yt9UNAhvCb6CglqNJOzof+KXpy1ua4vWmRRRowoFiqHMOc5t6+CW
u9gxcaUbxNTFcG7v24yyv/Ye6XwTLlJF6fQ6EfYOivlaenDY81V0SM8JxsXDRFj3ojsWZerAGWOa
//WZO/nV4bE4hAldFGQDj/n1hm6KmiHCsfgSlCzusJxQxRMx3FbDmtKL56LOuKc/mXghJr6dZSu3
+BY2K8XdsDC28xrRsl1e0+kWZS8Y1DzXchmUpBEZZ0HT9sA4ghZ2gSw0jkzi936w5FGNlKZSSCBd
4vXxhphTg4F03gVA31hl7z083LujGcxJmBjgEADCRx8CZkgJF4LrjNRydvu3r5wJyt3yxFLwHUMn
xbqOHJtg2jJ/gi5ZUGWMPuAgB0EILRrRdSvfkWPee/FvwzuA91FkAsnyjwd6zhB9Q4/hpsy16X0z
Y06kNvcbtkOYP4qf+74AAHsEfFFvL/8gTmRZ5yJM2FOoBHtS4HKI3fEwPKrZYqcWf0MB2RLC4rr5
6DpYpWnufuaREcq4r6m3qcmvk2GEce9lTZqfBKZPy6qMwr3xOpzBqnEhYCfeaFPIWxUg7B2eQcWW
o2zkl3DGrAN0LuPtCa6JTliwIkAHStiHiECkHjeKTl3knMRBTiQvJuH9s9O8GG7k2VPuE+WPRHDo
uGtdV42fiIUm5lUKbQsefaXEZINPkxD6crYrZ38t6/QoFTG1zOisyCI7PTzANI3tjjOTqCXrylRS
xA7lq5wZwQ68HP0tsLCt9n6SJVf0EnvM4+Rp75iXxCGj4n8ZG2JZTAye6SxQBlJC1f+KPzB2YgEu
02u0H9M/8z/SsUwoMt7kSrMgKwA9lrgg/8JaG9XOO2ljCtSxY+6xWvllt5Qrhr71gBj2rO7755Ba
9KokaBCneYnJhj7r2+BNZsjAjdN65tZkJbXUdtNyzn1wLrvNHNpGYCRdPm8JHwwJ6VYn/yV7kH/S
LaES+7Okdrysz4zx6sUvSw7ES3VzvTZ8aSPLZ0eH02YW5dr6yEb2+5i2i7UiPZXXa0A77mOZFtwS
LrOQW/AcvcQ9IYU94X1loxfoFm2uYdnbqu1Swfc6zq+UvGl+HZSIrX9rGrOvhczeuagQfFUvCVce
xk4hsZAKt91EBxolui/Nq3xnMGOGn2aL3GMLa1EXsG1h7t/uguw17yz527xXW2CQOTSu0QI32ras
PEJGN9wOJ58Bf/65rnJlvPwZkL5G8yFgjx2MJnGwXWoY+3GkGlu/b54BHO3OdoDOe/kEnjvybySX
2cHhiEHoNOBoIXzcwxowoQjR9o82ZXgkHXlHcZzDrmY4zXFJtaO2xXXVy4irgG6F4dvJ4BytdCfU
1/g9F07uzbdpO/kaZoRCqWyxlj+Dn2FUZtvMJ/qJ03IpfVXvAudm0ohq+8oKkn/BSoixfv3LIgeV
988cAh6sJRm3Ul/5EbBzRtOF9Lq3JGNMRkmAZcuYx7GXkcH1nYlRNOgqIjTufrrF7acBHpzCKZ2o
P1MhI7eryCUWbFpaQxpPRoL7ZskGfEnL3PhWMLnwgsp5kZpndztc3gD43ocJ5U4qItgbQNqAQ2mu
3KRwA7ZBrLp54qp1ZJg1/hq7JwGySCozfWg+u80URgDi1c0uXcp40PdYAzxz/TRgLuBdSG/7d76J
L4IlxJL9f1IKoGZWxQTiV9gCy0bcF5UPEzM0hJsnvFm2/Hs++Ber6ZBAxMELqayonNJ36N0RAUvS
YcG1iUTzFgZ4MQLc65EN6k+dR8uofyqYHDPxhUqYkSXtwtq5mmr1F0QgDl2sjdUxx5v27kVWZV/y
S2eejNNsRreJScdy1SIjF7MT2oIxGPOG5bKjUdlxLIMscQkqNaYJ7oUouqRxJplAxmhBhgePfEAY
SozLkwUvn4S8shbplZGQh6A5E+Y7BBHw7EdOvAwYrrcg7Leww2iiEOq6TG6qoOkqn+H4VNPP1kuA
9ckO18B/AQoDryVyQ+TAZfa4pnnYoc2EcSudgjqW7POczVXLtcOj9NUtlwQu1F4wcIKzdxtk7uPf
dz40XQVLHbgsA+QuZHbbwZ5q2D9qeUrdD0iZXMoyzKoPqoZYikMMBb/dORo/1UBHt8MrjHjyEwZn
39vllMEhf0tAzyIZkX2B5sc0xMdUeMp1NjoYwKs0VUoQtquhMRVGK8Y6hDLVq8HXfDXa6pH4+UpL
2Z1iDoEI0RMGQ0a0SV2iqT0tqWfgarKvHvcvDenWXXU/SyoAyTOM4EN2GU8B+VpU1aOQbSCmo6+d
aL0flwH/2UjPQ5lYbjA+SScivVu0tINsZYjPJXTonyO/aCiXeYhY8zIuNlY4bmJnpGAPCvbPPsvd
UKnTPjmXtzFD80sI5XcfYg4dwCtFkfBNqnnIQ4sNcocsdWnsKmANNu+EnVaWPYe1fb/2emv3XNMH
wekJmRv8WWvgjHzymyeKMbHdnhAUmcah0AffMAUlNbY1fLrfsroamnpE0Ebu/FIcgZvZ74d5ARws
a1FeXAw+TP6fARKRHLv51oxQx79hTXou4vKI3S5ASe3/sZozYiQrc+FhM76eduWSlGCHm61949Sy
YZumJNUFQsaklf3vm/k9SafAXxzp7Cv9hg0hPzeb78AQArx7wk/ENXCCaLi+IGTcv5hUr1ZCM236
V1lCUBupV0Lrt81DMZTKcuRcWcAHe06vfFnpDWlxytPt/1sOxM3vZF8wKl8+QpAminArNYwjiQMv
5KkHvfae4rNDe8rvVvimOFXVyiNACblkcQbDSNbAi4PGnOpVuUCxP2QL/Y/Kd2ztKvUExhtzx9vY
hCI3hQEZ/4oUPCecxmcFpuAmU1gADGIzPjYmdG/c0s6iO8LU9wgv51+sGOh6IikQKo/ThJD/EOnM
DHP2E5zF/NHM7Mv95KXQBYib8bsFmBOcnlIoB8bkaIelo2W5EZTloBKckGPY3z9vzPbaTKXvOWHU
wmqM8JbwXwIZhJPeyhVLdeXM11djlzcueoYGcB3LXTaDrX07xams+AUhB/O0n1OXxAjDftDZqnoU
grZ5lKvFCXQdk8QiKIg0ZvKLHkP3ySzFPWn7khR/+AUYXDtNnH89W2aq/t+4mxXW8ha6wG/w8Sne
R0PghEVNYYfv/KXKYiHiLo1g3rd4wLvNGANX5frQub+RR1oOn+qtE0akn6F3VAlChc6qj8ABJqEG
+Nm++xBP1dkuATv8cboHGCkQ1DVU6vBlNFwN77vCow/QFd5z2sbpUF2h63lX4tomyqlIJtLqI7Dy
hsPOehWBIvGcr8zUp80ae7elPJMqMTsfenpeyZOurGXQaFEFUi87B7/9ID4T7YKC5dYY/bGDQNPU
6Ab9QQmdx05u5YdzYjIE11togYql7m2bYNFh861RtfrA/6+Qt2Yi1iVISaYraG6e0czo2iTTsqRg
Pfxv2a+TYRMhxzoRhqA6gOHKOor9sMzypHNJokZIlaFCqg7T+WXzWHHeSW4E4rSjeo9jFf6f6ZX7
MMCghJVd0qlViRlmLbvZs4lBHCx5LIQsl6cT7aCyW2TgGsVtVO7vPtqdrDyS+P/tYLo+6R9JyeMb
69HmTc+rUfQqKS7TYzVzcYwexJsWeLB6EplA/KXZ3qwe3Zwx/Sz+6eQmrOgiSdFdnod7EKpAe+XN
c0Wct0xBWj4hC450PUkDB1y2PKFi6qRvrFzkIZpNlhwOf8Ji/ssAehWrfRJVzODscif0NYRoVoXv
mVz/OpLX8AxCgtIH5fZ7BKkuNysNN3ZMLzM9s04IQsp98ebrMr4mo0CAag1Ye9gkzKT9j8xSQizu
NoaHW7pXWlqDzR1msuwGEfbr/jd+N/V3eFyk/Op0OF+ZKk5bIb/HU1BY79yzuHaVHssOnkcM2Tq+
BIoehqZ7XEYGWPU1PmeSaFl93+UYuHuApB4hXBtO1I8mGFO3PPEasDw+yq7+57tXE8ROmy1nhHV9
ldj8z0Bh2ZTTYIlaKvLZWHHvS26bc9fSO7+4T0L7MJDP2GCZWqL1/DOVC1bBBrYWUZKjBZnSDFCi
VEfkQRNdXUuyebFbNXUwaAcp06vajdQbvVjVxpB57T3cbN9j/yu1xI73ROZLKC0ou0vCiPRMbsIY
NSdqMHu7BvwINti7199GfD/4AgUVOw7vLfp9a14e3VOr8mZLkqbG+k9r4hdiZL1TaoYybeGpTwp8
OeK33laRCmjdulQa9fIjfrS0IVI/bueNHrfJJgnbPMpZGMGQ90/gN38bFSa8vkrVUDOOAKV1xpOt
izuQxEhXKCCykcj8QJC2bhlYBEjkfpRGFXOq0TlNDO9hJibz5FvgGVjC1LxaxXMAExpAXvPpmGfD
ZjmRhsY9B2bM2kQPro0EjYzYtla0Vh7qXhcFc/dmqHBYqqMwJzAMWxhXkT5/48ZCBe46LNd551Lp
jKuAlq2lmyrOG9ntvu8irUl8GDKZPy1yvyJMa0oaqqECOKsHQ07M3jSHxMD9UJDA/KYR3rKSq++G
W0QGa7kERQaRvE8ehD9ikEHzokz1XvzQ4bESAUybSq9mNCqyGzI2lTJSrr6f1QNAEUeo4v7eJpup
C0EPZdO1s5sBuopRb6MRkmL0KO/Rasq9dYG7TFBt1/DJiuUVe5bDRkz/xxz0ySfsl4IaMbS75SZG
SwbTkRvBpVFj2/FOe8NaNOg/tmkr/OUCUf+aCm1QyqmMO9EFbMNK7XMvHUzeoEUB7NqGZvDrS22O
3wFSL0TE42WUauplwZF1gEo+S9JGsBg21Mo+qPZH+GJ2VwrQCDb9QINwIL3lp3FPoqoNNuIJKRUj
9MgKs3tCPaibZG/FlWIejd/yc4p12Lznys5hIhwpRBxg6J+ahTP5K4sTQjmvyBVjkQZS3ArE6wZx
uPy/wfKs915P+a/a2e7bsar1LDcfow/1wfBxrHp73jqh6lL6pe2bHhBbIGQ7ltketNUeBT9NQBkw
tL1jEVjnP7CEXoixT6455e5oj7aBPgVMVKSgNj+HG9xl6rmiU0yjMJ0UDpElDnTIP029Xl6/ONIB
5Ivie2g7Z+W4LalYXfUrtNfCXTHulzb6GqPCVb3hIAxKm6wQ1+l5bok3SmNk88EEsTSzU7U5ZaS7
hvkArl+XOEUlQq40mvROtPceZRr+G6cfW8dUo9ZXbmfD8menLF9A4ZfI0lQmVrlOi89ekCfPiIqG
fUhLs0k0o1C1j/PvdQRsCOfWVKaeM92Cg1qPSS4dw4FoEQ1LtlSvboIEob5tMlkA95dIhu2r43O5
fV2tDpxa901BBt1eoL8xaxxTwr5PFeEZcuIN5itujtBDN3B/ZP5GgV7adlCr9hbGdwB9A/3cnis8
aTXX7VshS25b4AMJ7J6F9QRhMuES820mYPlq1XbyLwLx49O7rVYvYO+bZIsJeS0pbfm1BmyWktgW
0L92fPokQ5y2wwTbCneAglDXfhDrAggxMbWhQslhlfZc4ZU34j3DGsJPbaYbcOThwD4w+7Dkzdj1
i5zGFmQTTRedaC/fq7uDJlUK8kORVFJtpt2wWkwR/hrdxpE7SSvuD4lahSisDIXEt2mvOs9ivXFe
925iOWQdM+C9RaOkT4tN2YnUQqb/IPwf9ValXD0qO6m7biTJ1zK4GP2JYoKxZ4cDKBTFfzIWw+lZ
Cveoem58HCnu/8jajyY9jRxxE9WWylqwk9TD/syyezZN1BfVfDV1KzyQKmV3JvuF7ZtF3LlSmf0x
aHQm/zPbMdkk2A3+jzDP9Hp04LYQlhTjXeHW37019ZTAgq8vcpHzR9IqzhcXXDahGa+th/KKBsCw
+FXO0NxFUCffg0tjB/2yNuUR4c9U90XpR2t8UNPjlAWv1PYoNbVrYQ4E0kbLndW9TF6PofbvVTTk
zDFe9+YeO9uXsBRQQkWoGUJiOUPP5P97WPGHPGUJnYlus9Ne6Zht3iHAvrKGlstf/JytIMEQD8hB
c2+X2cqva8faGUS9KYAF31v0+LdpO48f8IVmnb9y5cy7zXC8SchDjEy6sV3E53izEwb3QyFmrwyX
z4HPwAOHe/dYvSY/sORphH0EzP2f0B3C/92YGMjnxQ4YBRUe7Coh8aooALyxriNwQwocQd33X22V
WtQbGGe9wKv5518sEMdW/RQNPMQVV31ga2Tv7VqEmqlQ1qWowzbRWalAAbY2tV3n5/BjXJ/bHWjR
gdFlkx48oq61SQpUtjf49NcikyY5jXGu65tKabqxm4RGjwsAboTNduqkeGkHj5tC2b3Jf2BZipWa
J2HAwuzrN6QaummqVTzYJqh5Zkwm98mdJrPCyudPCrEm+SbdzmPR3ygA40nawMXs1+U3c0BV07on
Hl2bjEMrKheHLGx825NDKMRdbEAbboPox4lvLJZn+vkb3pQjV1fCKJDlCen2F5DPpUGrHvdjKowY
dZAx/P/cxvVQCbBgZSpal4lqGXs80cvplAS/zNT9CV7I/r8iCU1+7jF9nhvzFvF07rflVhG4nzxm
ji7xl1DA1H2DijO6pMIyUe8onl5IW7S2GZpm8cELnk8wiA+PANhyBR9LUxDaA+Z4B921Mp0RFwpu
Ep7hYOdvUsKexT1ifmDVZH5NA2Yc9jgnuYOPFOVCnJmXquezyKRtCyzb4/wE4CcNK4eYoWDWf23y
SVfLGctn88p7x5/ToMTse7NfGgO1sEpe+x+iTIrtchd6DIOo68pPDT8mu1O1T493orhEZ1Lkc5Rz
eDopfHdj7e0NfsZ3ctzlze70teCIJXZSziLTOTjf8NfgQCV8OY1aZ9M8IBdLkhCTN8AA7XGyXuUA
i6qsZKwTHJqV/VvWYWWfMqZAK3wBGGg7hy4C8RsdC034GBrR6fP5mAcwQRFXpb082PERxfL++cvd
0ix5Y2371zXi74gRfua0v+p22XPMWwEIjVr6os9bpkb6h77PMzBYuqMwBNsLF4QiT2BCMCM5bv/a
+eJv0MH6886Sim1QIIBPZtz49Wu0euW/pKPQjgZF3oYls0M3mw6pbnma0EENPSEbR+fKiZMTpGN8
y5wrW9TuxJqRzTEf0vjai7nThZAhlBIA54SdGzq3HH/2o+RPEx5wMDQzBn9zzroCJSrkqmsvyST3
dwcvEzTG+iT07/zUXyzNnwqMC2DckgI138/IL0UzDF+i3/b+5F2IWc2SLs7PC9OQgKdGScCpqRjf
lJMsa4zFILmuEMZGbI58o8dnCZp6wZBVf9X53/TWnCu5YU7BY8yK/18yhO1cfrVGgPVZSz1dD8jp
hKXIRFokhhIROej6v4iSDmD/EajEexxfP7wEk7JRNiNCbPaSqiZlyeOpB1stZqFwZOK6TH55slr2
sYwfg9DasI6vlEOMhVmGpQchQi9M3cb6sEUNUCZiVunG3XA/pTNrY5ZQiEtMxV277L1hJjWnSfGK
9BqeB9ZyfAYJvirVMYP1jtBCNYdM+k7limMGJ/2B1wDO6Na1tRmvqrvRfaCkvyiZZND4Li7CR8M3
rentzwGgI0ls40XVHBQkRV+Ptztyy9h/JE+Q2Te/TjotAfUwZJo7Jtln9f248jtZXCCamtl2upi+
MSWnq4rjIKbsBUmnh7538iF3JUR89FhnOwWfoN+S+shA72n2/lRU0Jv4eKiNubxyT+IDJZB14fY0
pniumQCBM6xvepZlI4E/h39DOFBoHKtYqHRySyyqGQHF6TAqyXR1mcnJW9nokH+JeMMl3igcVk2/
9U6WQSCIbT7ixQxjY2asZN8H4BUUioa33f9FGy6VyLRWuxkKyC/MIoOPz+mZzeNZNFLEugKsz27F
RmqvDfuOgt+YHMojjSnWBaskkehsuZhzV+/zOCnTIr2ubiwe88kqvjMS3cK5WfIiYLkHoH+BBazD
wGdr+0MuS7Dp8cJPicy0qMNEWgKDASw91zM71GkyujPE82t9QX1lJqxwrDPRljYTc1D+l9p/4M/y
8FeJaL5KpITG/mlCw2EHu7FPV6FrJKwpQEODq8Zupm2i0GAKmXjdOVD9+N5x9YVQS3XS/0qGSpmn
Td5y5Px076oh9jQW9VF8RBHZLuDCV3FsjnZWZnu+0dmjRoel1TjNORok8PKqR/9sDRwIvpOhuovH
tmqAFhDcvGOa48SxEWcJTdaMktrHEFwB/FOsikSD7iVuJuqrE4GR5q64Hi0KeEKMJC9cytYqauGB
t35JikqgQklK5D8jEH2dd25WkPPLMK50u0wlyY7K+qEIOgTIXfppkWU3ywKkqDoDPvPdAiq9uuWf
vFjGcxGZ7EENDBYwMJT6WDNuyLtWnSfmh6efprcukwSZWJl5wSeKulISpPG8a+stdusOlBkjI1GA
NKxz4EGKgq0xKAVGJTvaR4Ee4VEnMEOIjOdG3ACi2CxP0yckg0DM9KHNFx6odoCcRynbVARPoP5t
VcGc9D218wqQpSaComfbIXSA6dvl+kJexxdOMOy7xfBLLOtAPw5xpUfFQyriKl1Chh8hN8oGlXQv
fxbZFBUYxCTrauEuEwDRbAv8KHXTotytwSJQxsbvYJt5161WSUOdWRnahGOIAE+mZMn2a8x+y51U
kYs1vKXN/1f4vJMxLYiAEXGYs9xnhWrpK1w/vG8tajfX//+Si18eeLzLbGiAZgLBESr6uEnDLZBP
mh4VWeUeNIilt3pi4sPwDV5Z9CVMSPKYh4/8f+MiqcPGw9TOrKxevPqhizYMpYa7Pf0B38+QYPB+
xKPYyNaIZXocb8t5EIK7iNfcTGPpqBfm7S677j5EkbH8IQmpxvMR+ReZjoeekCEVw/nhjRjtbFEY
8ayFckescvPf7ng0m9W33FLyB2MJuVhr4jVsihPUZraLX72Io16UwmuZEPLkJxkzsUGNwemy/qde
nG4gDCZszkVKQAM4/1dxSl1kPUZasVnLlywLYUxVxpvmRN7e+acMZAHnr9x0CCxKRKMMUYm/vCmq
2IioYatEbi0uN5a3z8D6fyJr2Rgo3E+KyyHBJjJHRjErvVwS7NKI0F3H9zSzUzx8TqGBnVxtRaPZ
4OYrCE+Kafw/8qrmGJ7IwEg7/9A8xKCxuXhWQOoUG8sgoMWVoCM29wOZuyXzzOcwDeskiFDPmZpz
pNeH5ZRCum/JaROvpvQ8sHgAv6KkCX4edE24L4al6fzb31B9kWOZQz5f2aoTYJcpCH7noZqSHLcm
8MYyWNNiWjm5cBkIts66mD4fLO4Tnp+XxzSm+Q/TV1esCyNZGJAGElefqBLjhqbpajkG21Fv6Mq0
ObprlNJbCN3Dz435iNeYFd3JbLxldXn28NS2l8Pj4ZQpup1dwK9jWDBLROR2kmY3ZMoeL2Waft0K
pFLv/n3QqZzuEiPfVkKRchcV+Bhch/t35XPymvjZ7AbvhvdMYZ7ODnnab84Yy8fq0g0Z8Qk2V7//
/BHv1iGI+oUQAsKlRmmWjQr0PTGVGck32L7EX2HqnA0RGo71RggjegwdXcirdCaCsNXQbF8JToa3
uJrD+YF66F5JrUIKz6XF0Hn1Xmp5C4PORyBIn/FaAOfLTLjDt2/+pwNzRe1/yC/dP6VpMmR/iRS7
7ic5NTS7IfiDenQFpb4bQLWK78WwxHvCB+yyiF41OyzU27yvJ8KRJXavnTBr18mUpaG/nhyZA9KQ
6V0EoGwGJ2P79V9zEdo9QJabRv6Rki6NrRZFxqHJPEyLG5xqUfnstmRHMQYD0BgztXzB0J7L+IlF
pOgsScMWxyYYBhJBkGPflGXElQmeIWvwSubp32w7Q72v1Czdch/WO16Ur98ipEOQEnYW/tBeKYn7
G0K6r7H6qeud/QQJxGN5Yjr5tKuX8VrXaE2NSj82HaYqQRl6INyqozS0q6/YZzRdbPt7mzcq4IN9
5GsM7UPvPgeWFAkTzmNWtcBYSnsfLmcTCqMVVOGjuvMv6wpPRsPeFAHTgVje+UTvqb0d20sz7zB7
/B1/NbWnxprq1+s1kPk8soJVrNKTXVkk2ImazOz3fKWE3WuYo0dmfZ2MC0qC5Fk8Y1m6U0tJjmh1
J1bcF5SbK7BKzJvrwEYJK4+mfmA5007LfY98PFylwrRTtTP1Cv2+L5cYdHFuPAkGIANPMdkYvGbz
20ATWNUq7dibjmRGXU6ByouprlEff8hgIQC8BMr1ybtRzM6JbungOXKg7MCmpIz/1UL/U0LLr9EF
+8xe5JS4oCloKjbslPDD6hcpE3Q9gQlMsf3Nnk0II8cJedpnUUvwxZ7PcOO198iZrtCZL8m8bTED
5lMbfmSPu15wfMuBR6W8RtY6F6Clk4RrsdfUeHN/QK7lu1eKIS+eH4EUs61S7SPfDolgdpJJd0th
fRzc1gN39qHr3xKIEeDTMsCQ7PfhArsiPhUse/b7tgnrZfNiDjeKc5UV92F9L4/9xrY+pigXGD77
ujNlPYAccRGaSj1YFdfsgyKOl9jotmTOWgbL62LxymVLoJ8jNdGqJTJSACJ47pxAuWTblhW7fLPj
wfbiuuXayO2upZ5AM/LuhfgAwlSuD8mifVC++h4eyj1j8h9IyY38bcFqKeycBlMIHv6cyvmuLN/j
R65d3AOKbp2Dm9NHGGDz7gu3GtHC4eAbkmUDhOONfxhc06ZDPqIr/7ysyVsEyWTKgeVWW4gKHVY0
0gELdYIX+d4D7zL6Ba0l0VZRsH78NMEJNPEqDFt3b28s4z8/YW7sa77GDOLb72PDWAZMerD2ZH5u
G6bONYtckvMd1Jk2UYcIJAbIzz3JQQjsCOcegR7vz4cZZBtrO4pyGAXLupyYbVREEwojXxG5jhKi
ykAo/kFz0sfSVAWRAFpDb+IzTkpbXhv34KTqzDI9Jur7IYJWkBJhyIzevRh4gHQa/+tmPX18tdBV
llr+gmfFT1w2OKNococi90CrH92KFWuDbY61VqFbBJmov2CKIE6c+wXgdp2vqUVJp52HCRy01Ycb
bVhB7voLvdBdtOVxcb34ggTWBwUoea3OtNcscB53/br4034gLUn3hasGDm6uuzPBT++dvDGv/e8R
CQZvyZpsaZoQ3S/5X0i2INZa5DgBHIJe7gDwy6kAugCzUbnknzUNYvsTHg43mtOfbZvXqTTZtKd/
Xd1CcZ0KaGwE/khTA06IC3SW2eBXVdmVE0aAbETJZfOcjrjIi2dM7pxFtaPomqHMZ8ZVUtOJKqVS
u79Kl+aYJORM9oGB/1Mr8RWNFt0ezAEbUBky9rkbEvKWGgpVw8tkQugMm3a8/VNyRglV/qTEyGKb
GLChopyHkVTpfuf6+bqQCh3NrexCb5QyLLpVg2fuk0IA/J5PShq/5DL7wvKM42li9qdlX7Wuwnzd
nqozaCYQpnOtEWVi6wzbw6PO37hXU5X47+KrbZBnpIthbK1NZQlHyKB/cS/RS2kZc9bUrSt6ifXP
ycvDdSWyLP1r/viZ2v+lwnBBm80kqsgTM7198nckfMLmGli8I7bY9Pz1YEJWqmDqqCcoxDwkYBak
AxiiY4FxbuIWHTLPhQXiaAY5OusGczEzU1qM3t4jFHGGWSUNkHor+UUVytJTHkTKb247u2fvOc4U
pMQ4QCh/41KlO1qCtZ1v/Nm09fCwmEjLNPW9ZuB394RcYrw4V0NMoOrvPincYKRc97iRmtBYDSUD
hqUTSTgzd1WB23yt6Np08M3N6oUFvy+xVbqZqrElFLLDChYtk90aB8F2Yn+/mfdKTkydKP5jFh10
HULIM3JVSx+++s+X4pSHu+oN5azSGqSCH6xy0bgwmdw0W741gr/vBab3qPa7SCtf7fr6eHcvAKhq
OF7m6iUqyDGsFLPBHNLbqVNYy8d6M18V00MUmb3NuinPD/9QAGqG9R8vL3hh7QWzig/zIlmagm4e
2Us2vkmlcEygrio7m+ni5a/QgIfJovrzwrZbFNjvxU9b1UpKgIxigJeTCfy6J3DqoW9yqQX5s6Pz
oerQrcwoLIrsGgDHrVBVpyHC/b2Hws+TrbSaafwHja7IvZuU34d8mpzf9kP7szpcN83CmJCUZqjW
Ug9JWfpDi7xnZaKiuDTPbJ64dY/dUI9QKGfWKBLw8LFTk0a7a5chZoWBGqWam8xoDnd99APRZ2GN
0iQDLFKInPoO0JPSmWwrcKCM58ySKn7A0aXXMKanu00Lpbm3aoTWKWTxFM4KOFWkng7AG8pjWSyT
x38VlSOuE9jC2q/i5Kz6a8AkA3Ff6mb1kxLjNyMs4mkWyVGm+JcMC1MAExKwxsXUC6pvgf7DNhrt
BsMUU/wUilxl0tiVoNCTZ/gqZCeXkLY6CVVVdUCZYKeMSwfL2HgKKFqRa5DEeaz4mLjwvA3w4k04
OHyMC4/NBrhFa63ppyB4qKB070ry8XDZQzDDtNrZJMi2buelYmbVpZT0niO9uP0BCERigdHXM9cy
k55lWoKV93fxYRLLzzgNLPRKX2026YozjF21W/NvwUSuwFaVBnzBOu2YzddH8w+C0USGX8henPFg
Z15FHLwCZAjfLU8iS77cUmpiQxLJHfZZyX697bQDfrkrNWPepGVgdXxL3Dpmfwixcoa6kVQ1hLr/
kB8BDCuJ2z/Z7YQZ+KmNlf6UfpzWy5VkwabWijNu7+J/8R1hdOs6CmoM5KAc4/C7DEJ6FW+qf+tI
/u1vyIIqHGM/tTUs1CZkVULDS+LYENU0sKxyWgMghf3t9zn2uBHCFhHy0ZFHbiAp0ORQFL39aMtK
9nlMlqy9tPyxC/X7S2PYJ466qrgB6XZsXdJj+IeXwuaVtbmmkbAn+EcKl/QStqY22WsO+RzCJo3O
Lj/GXygPJT/Nt8hSSW4OKMkWtZpB63uMMZaUvHswAVS5TJHE+b6ANqx5oohpJ3vvk42tKNmdtnCc
bensrDZtcIyNjYPrPXFrv9Fz46N6W8TUqAuq6yu2iZcCGR9ZNcIIKHJptB3XW7v9fbRxW7VCT8sC
WOYYSAwuhRC+dWxgvrUEyyeBRisGNJTWB5o6gPgK6KpWGa+p2g9AMbCp43TQ9xpdphiQJ/a4D7fV
+1Ut4GE3ODxCNTAcmx1JXh3fQuLrpijkJY94fm/KjttKkvlJQAVoFgqzB36oO+batrOEO0g5b4Zi
5MxInzu+Jahu218GgDTfTYeH2t0cwACd9MByUF7Uf9maN9HDewkWOGFifufBIJG013EOMeCos5pl
BNpBBZI4y2BNCeG0eAeZz9tULI0aVEeVe0eoHb6Eg6RWj/zjELnawikdfzDu/1WLJKgzlU49YctZ
enlU9IYB/jlaGoVj39bYNH0izYCv9gedjF7xFJC8Rky+5JLxZXn3/XsJ0seOOaUiXqlBbFIMpDUN
bPrZSd9G5v6YnkxuSPgOB16etGJ+G7i+iSX5vLfJXcoHVImY8MabuBht67GSRnmtfo9G7ZY3j1lN
+I/7ZFUcTSHFN691rSmNaBiZE2cvRTuUXdSslqz302G6wLndzpiaAg/O/ZN9KYqhvEIpqfF5jd1e
kCUgKGRFE3DKaKSn3apYd4asGWnvfiDrIqI1+6b1BNo70CJ55/962WXfWnyPtdPhv01+jBa5ln0V
T/oZXJGqJ/FWZWgKTsxqN/3yJuX2FirHOCVKAUFIGK8pPhXk8FJItmSETXm+HAwqbUZvw3+h8jMd
xXaM/7pOb6nGOG/7wPPrjZTZHjPWP72DvESRwRb9Na7+JKhSP2ujuwtgXPUOwyM8KsOxQrtQmMOh
EPeLiEb6vsc6a8G8WTQLyJgSfamdgVxhzehVMAA9nnKyUAzknTeUJKBeDru0DtVwPN7U6vTxa1sl
qlPp1DGf5VW084jhDA67XXHdnQyg6RYN78/lHCagrqW1Cy2W/j6a3J3WLO1MdB8GYg0Es/GOb+N6
uELupyujRLGBKpyg9qDqMez/USaPXTK2qXDpYh8gR5OMMKuzOWLo1rjkrkOXc89OJBsr9NSjyUOJ
+r88wFU9tRUlcgS6jZFx26kM2DXS0pwPdZDHC6nccXGj+F21kYvFPwE8dOfm7KlpQBhiseg6RQ0A
Eo+1fmk0fDZcN1bHyvt8urrWOrabjYtQ9kB+OmzWLHVAUgl66HW/yvkwcRemj2BVFmqYjgTCgjua
3eAziTbBb6AOBDTdSTK1LEQrzIcjQih2ryCqNjfAdUpA6Ymhl1I1P+ynmdms59xv7xKbp2+OZVoj
HYwL65ARyWYMZQ/tyne7bTfrnKi7OHpuzQAMm6otCQuhc1WI1NGNEFnjBqXJ6/hBJFy+caIblxFY
TY2sSJ7EN18/rihcmEzxeRh1ntpGpzBR6ww5l4/8gvPvzw/5oUHhnQr2a2a7xYp3ry37KXuZsQcG
M0NpeBIuUiZVN5C7JSFnhEnTTcx3JUjrXfdE4kmFyUdHHHHu81XDxBuaSzJEJHACvTY3BCJEfJTj
X9QJFyKY0aPs74qj1oW/joX2qikImEZyX0/IsD5e/ATbHAfs1otap+LXZdDToBdAN4oFfgihXF7W
UKGwR/Wnoo0/UADkg9V4vDIhsn3FRk+WU0e2MF2iLzX5SpWQICpEVC5CQNN0binj3G2uIWe1/zMk
ZS1SxVwmPbhxG5m0KcasVPJyZ4Hr1FJSSODUAQmuRm64KOvK87hUO0Q3DY5ANgqXpEo80vIzL6Wb
DRqSdNb607wdhY4UmHakoTDcphnnSQyKAaPQWaOmhsk6j56ByAWP6JLhvHICwSObvlAyUdyTAiHx
d0JNzAkWWYBzlptV7CblDSPPq4vjlsld2WrgUiS5QLO7uLSHKYhJYpOaJ1oYZxmrE2UhjOmYD1FQ
iDZmGLA4Pdvopv6mxHUJtn1f/7z4oy4Ewqpl4iRMNbKqW6HKswmy4erIfjcITbRnDR9J38aPwzWJ
eLC+k7Tchi7L/yW0i4q6ysiBzcFEtoKQBk6A8+hiZd57/EByrtDwywCZhNOaMP1pdPQUvIgW0zdg
vW4b3BsSPe+sSQBLW9pR/vZ0JZxI8JITl9qtSiRrvY6aKhwNyJSVbTAm9+HdszFMut8RdkD5bN10
ehQ9uG/FDKRCUJM1p4jvxEpvSd+M7bLjrcNvvA3V8n3wXaeMm8Gn0IYLH+QwbvEAAyylm8MkbjRs
HqM8JDq7CwXLeQJwmmtMi4AQOgE/EnKGsf+AWd78iTX3ZmT7DxCAAqS7kKYELudvjQrpglO8ey1o
RlUji7msgKQlZ8aLIxlnjNfPhu8BXquVe8cJgDarCqwZsKhKUmgzOUGmPTDNHYtXiPIEdfCMtnub
hPJ4uQmvQGAyk7yg30PJsthm+fljK9usu4p5BnU+koxZxBYkBJFaqYGXPQN8YIlN28x7n547esgz
o3qHcny3n0W5GJ8awIDqJ7d8r/cOiA4fgtC62doqGFQny0cC0nIjMMEEZ0nySeSx/UYmy17GRpqE
otegzrpBG5VghgsrDa0iARS4Z04uS/FQeUpqAhw77Pd+GKVyPNR4DvHf1fTvfvSeqHkekPJ5JGL8
9TcBeDQCes5VzZcO4ffqpTF63n2A18eG3Lu7PJ2bx0BRyEXsiZ0AROI8hEt1USijel7GcwXxlPhS
LUR76EKcw8nDvWPfkTOOfeXGwimcS4EVwHO1BM8d1J3xWGP5tv5+l+8UpU1KLwW6P9JCboWbeO4b
vHl0oXk91v5oGrwL4zYsPEGeXhX8xyGIA7AgJvby8CxkDP7iXZVLSu9aE7p3WHWazyyUYFrCGCHm
PYgmE3JyYNax2ACA2Zrz01D5fUl/vrRl4i+8Tu/U5G3mBgi6axiyY2mKDN24bWCjJkZUk9m4cDL/
xvfRpjDj9zFE4Wi+Zb4rsgKZfyvmltLAhRXL9APdBC1XN2DDxpPWch2S+vYwajQ6M6/6LsE2Jsjw
GRmxhLG3JJyx8g4zVhfBTCrSb2ag0udT1ZmhFPMiPvpxoSvQ6zjRU0rkdD25KJM9jWABK+wcsurh
ixwS9oMlNz+nx5HkI7PMMucXL0XPehN4ehZGxQqhzRlZ6pdKbhsHPbxit+1YHUKmgYJZlyRocy96
0kg6z1iywNM4RI4FrGTfSvAgpVKSH94KHYVM2v50dK7AhZCMIfeHYa5qX+AYQIoJHO3skfmSGEJE
Bakxqi2wsdSwqQNU1/S/LRfnbvNnJuJ0qcfYjmXyXf1zsnb//0mfegD4oHhIfbaRy+h+0lWmvDD4
NZQd/FT3062T5wcrmxtwj9eseF6sl5OdZy+qDTFuVki/T8Zs43ugggmS20m4IPBY1Lq07EwVuynJ
5irwGtQMosVXbFe+8DapeZxxA0Q6CSmxLCLzDeW+HbKs5pqtooSX4rOJWhqzRJygu8EZeAMnk8AY
84cghWkeb7XB1fygO1wLA6UiaRcHhqIrOM1iSFDuWXFTqAzy/t5FV94rlHkDztFotdx8K4T7neuY
MUmxkRG5QuGehSeQktOrhaQd2RNllvgl5f20kMRepvOlOg4CaQ3Yhx+zBMcI1k6yWY+jS0vYnqvx
ylHIQpk4rJv+0OcxAin1N5NC2GMFXgulz4ppWY0B0cY/p5NZT2Dakvx8AtPiIUG6odx68xugxyXv
bxX4HnAkBHweRnMeVF4RIA7pNyn/bPfo3j3wq4UCpMPWJywZB4qLDGtgipuOuXjfZXgLHJsJ2lHM
syj5V7JmRV5Tc9/UQUbouIFbT1IGNDchuN4Y7pCFPwukxsciRNT4Uc6/uzbAvRbeMXc7RkNfXiLD
Vz+23bYawwV/imKiUVTEfP6FXnsmFgfHGrr/7tvcdSu9UuhqA7tBQmCLLSND1q7t1CIV8zmlsVWQ
9Lz8ZXm8Y25JnGMd2sm7ZfJfPhSRPmrUcAuhgiHL3zDgTnrfuLJRIFg+fYq02TOU2g1GVJUxikSe
aB6UKBzZWfCUV0T5DJhIrMjXedjUd6fYC0Yl2qvWhACU87hhUfMOITCqbaLOGbmD4tVQn5CaCmU/
AzSuOp7bBzaIajQCTpYhqP8QmkNWnkc3HyO6FWG5/pW1EBhvj4r4ppQH6uHX87HwruAv6lLszORV
y6DKYrVcZ7twZByu05lhn6k2UoewjaUhkjBifop3jbF79TJ+TqxNldFvle3umqHvtqvSgHUSzujX
S0amrLAm2Alb8ikikyrpvggLIFq8CAU+nwDBrPSO8fgCTjuCFgGgTvi2pYClS/VRV3KWd4jNASty
hHN/kqDArQDSYbWGsZm3NY20cxluI/d7gDaBSAzqxj42vQmiM6x0zRePzENrbQ4bLA1UsBkVWzEx
KuC94qbtlVtTwTqGJmEoFhxYoEG6CLc08Lbkc2LSBR1bDqxIqTbN1be9dlkdmEg+GUY5ryuvNH4X
rg1DjvcrYJtuS9TnEnFHaxnDcvE8az6rishjdcLuo1Ncy2225PMv09jBTYuGjrg/142yILobrEgW
ehh/6cl5I9j0RLxmJv8tcF0wcNx4kMgoWBWx6c2/gDMiUqICF0iatd+sGXuI3Lq++/vO5DGZwdMX
0/s2ZfdLXGQjCr+5chM6IxooSBSaid6jN9aJv1gg8nvV/69OKBJL9gH/q6C8VHlQkZ+yL9/gu8Dn
RjnE1axmyAKdxWSD7YUTg+T1+wIfxTCPwOp2X/aCAduD9JUHXKsklESGrSUuq2ST2R0gzkq2HWTN
+fUJD5pffzftESo75Za51llQo2m2gOFp3fuWjWK9QOmdWAP+Xl397Bwgt2+wzIYmqv8r9O2CS6SU
SAYR3BL3J6RKFl2At0/WwHqC8wBzs/eIk6Km7nqRSBVhP/jNlPVdEQC3KhpOFIbqlyFecvSv+I1M
CtJmy7PkxChCcOZZZWRyVAQlh8f/46dsv7PNyZJJWJakzuFDYsWPX1P/EoE12/YK3tnzUXj1y1rt
tuuKxL/icf1gxY5gMR/XljsfKsoRbnMNYC05nibP7+6Qb2Yjh5xU9NAhfJqf94ydWDjjb1SLFN+E
/k4J03GhzuJ64UYLPDehnsCjSwfcZ8tHDiDrOW+uJmXuJ5Md7liAr+33Obmnc7XZ+r6/4Urz7R6k
uMde91znAvx3nwUzPSd9t4MpLgAfItIbZSDq1lG27dmEC7tS6gsIE3zFplCB/bQ7b0OC6Iq/G6sQ
hPzWFKWrHD0bG6DHRGFdPJgb0UT0uGyVydcaWuPaG7thchxGAln8oHPSqN9vcPCyWPJQJUS50gGx
Rr11ywH/JzB/Tli8baLA5h1bwAhSjarORuLwXCEihjkgh6qXHK8V4ntSGkw58cjFPv6tMsK+Bw3B
X3T+XeljmOBV8l0YQjF8PZEHwY5bzIHIaBNUJtOulGo6ZytkRE5YqtMV483SuW5tizhDJXKMYxde
fJn4wMd5dUIe+VxxN8cdAFkbDXNQRxTISj2mGYsvTG0I6oMWAzMTmM2KzawXyZu9Rc5QGsKinVzW
ukchy08iiTrFFKrTe/AX6Itok45E2Xx3Wk8G3Va/3XTJQgVwsI5B405EC26/4Jw6CF4mzcjQ/L/0
G99d+bAdTNDZ3sj1ABxtAAvPoJc+IWeBiD5t48//T5hnRmb+8qTT5uVWGdw+hp5GveDGbZmgEH6k
dSvkhlTRqbjsTKRayi5kBKKVR061D9UmGjD8/cAsOc9EJRBGISVnLdvSnoPnjztUm+hBX1SL4W4H
orud5o2ivWBFjxa4wqJgWUjGl9sKvs8hyPkMFp50YuPG5xwJTT5VjrKwzzBE51kim/aGZga5CQNp
v2dFxRVOPFOyRjmV0TX5m6iz7up030eQDKnnVR9NcKIhC4yFjc+K/CG7XAs355wrIX3ZcibIo4ZM
kCUjKbDPsbOPYthESMWFR8ClC6usaSm2hNesYqdz90FocJvvzzVMwfibK4JDV8uNMjrIV3UZT78B
gwl8JH1dr3guJJDrJZma2v1LLrS+bLL/bsnwtitOk3jKnhLUNdEBMpCCINt/WfMMx7hfhZHUP+Dr
+6IfiaPewUdMjKVFUdeUMumhcBGMudBmcgsELrsfGTXX8+L+UJRDbmwK46ivfV4glOfJTRvs17FO
MSUg9PiQvhws4vwWg1FPRqOT3IuWlogwJ9mbR3tgaX7SG4PZh5UBjYwC4wbmrEnTUE3sNlxuViQY
NRJ+cIuBOCuhIfHd4o4wbp5+qxRfj53BRy1AQrdT4iJQsTD5xbeMHCKSQRAbhuo6WN27JlpWVWHW
gOfve+orBCwgWcfLKiv+HmgtoVfXaEDFCHVnFCY2fdoxbN4GLB/Sv7Yd2l03COj6nyoNdqdSka6h
JvexMjgCDTq6sA63/lzE2kAS+0yFOt97DWUou/Nv2qwudMThaOWzsYawprQWS00H8auamya5k6aH
m6cT0xgxvTDJb4+E1KCaE3ad0+30iNWjNJrAnxsrQdDwbfF9BwuQ9b7WhcSNDw9pMcTU32M09FAh
+83+EwbbFLapeQQJQ60YJFCJQuRMOJG41VN9yfgu4rr6qq2KJ+HuDSg0Ewl4OmBBNW8xofguBt8L
9MSXBpwDqhP1DM+J2DFhxpbq5j8XtjVQ/rQjbmkRVqU7X7zIFO61u2ptxPlV7gxJ3cmBqO8waMRz
ep3H56y+eUhiMRm5nuf9iDc6aU8u/spCPqY1qQjEuqUXTzQ/lE0Ja4MVxbTPMrxHjOUk9DF8E0CU
k+Zp1MfvxC06iAjNu5Yx9ZlIY95wUbtpMlKrc0EOQkuxhI6sdzQnJum0QKwGo6LgEuQPuHa918TX
UVk4oHMJqBHiK0loJb6+DtEJsYv9HL7xE+IUi3OyOu0lDiy5D4XEnesHlVtxwh8MfIrAno+tUyZm
TZule+sEy5cv23tGRlPLIjfpJCi1AGI9gD6AF3FlbDGyhqNSuRTQ6UM5/kg6aXDuC59ubg1WqRsO
rbF5GL8PIHEyO00or41fXI+BoCpO3AOMTyc+Ke5Cpm9srI/P6xbI3vBMLx24YleBRCmFfGlqKZ3C
hYglYsccJcVnrtPAsSGOcU1HtOmn2MbrGjY+WxGIsw/Txwqnkz8nt3Pv3VKOm5Zfd3FBFDp7JAEh
Olf6IQTQWgYpxhoiQPGDDE8f7Q+6UADY8W3RF7wUGGPjN5lyqIw+SPPcoZ2xiEPlG1ZCl3vdlFXg
XhoWk8TLQ02LlOy041IxjzHJb1oo1SmSC67qE3xcWhh/PxMQaiy8Zs1sM8am7kWtE0wRS4EnnkS3
pcAGnxNh9T8btbgkzP0Q0Q7xS/RtORY/B4wwfFyHdwBDGNWQjg+4c1R3n99kOLKvXRzUiWkqYDoO
MjjUvwu6fBTs3Kk/0JDlCtBwpE5PXRQnkSHq+d881rCk38sO8H2xk0Lp9wRsNZCWhlZm9XgYrgYa
HhUGLqywXMTrL5p4JmLc0NoePLSG74R4oqUYj1JCvwfWKNRxs9dZm6hsNvQEP9MG1WZr0SowNmVa
H8Teb8LHGV05INobaToppIWTNz8oaiFApy4oOs9MM1qhsLhCGgWZ2agqdfZI+NF0qKcgNmeI7RLl
spEpHgQYbNsQHH3aIzGk2ng5kPBYLJDd3OGwdAMxk42pzV2dX0j1f81pAJk0mBGeSI7bXBRgRRZG
QpAIO3kYYviZ/ZgSvOLtzmMGWLH4myrqTvzhDdUY/IBTmY+KnxHDWEcqW8twkRJrJfXp5dSrYv1O
1bO7YAtQ3emOpSZwri/CfWqK/1C/f0hi3K4FWwxfVclWxyNeLEfc+8AAQN42grhVg5LFIJlQF6kO
MegLAxRlbxVxlwn/CFPq2IaE8S23aWpjexnhy4EjSNrKw3FAiaMYzDyiCojipcZt2PlPQ5gEzpa7
fE65NvdidljZTRQNECH/UdNujkx5tdWH58eeDqAcfktR0SnbH9iZSfLu7SAsAXi2wptX8mpwCdqr
4PFlDX47fxzqSLHXinQ8WoEwTLub8j4EZMXp5K10+pk3d42myWJ9vpc0bxFSbYVm4fFmplq56N6C
Y8XB9Qhul/JjON+KMIUZEzhV3gnRKF7i+6RYUBW6c0XYrjAp5mvPbeOoDs5w04nCtxo03XK4OyIC
5uU5ZR1Xql5jK2kW1Sv8dUGH1qj0wphqt0B0b2rGT11NUz8IKsNZO2izoqbypS5gsgFa+c9WBPNi
5nxhlZ8rQ0pz3W/6rMO+FJAykZX8dtrynbgD+tCpDDSIbFnddJSYnOiokuiEI4mUzBECb336EGOB
AnzKD5aAzIvLqKpK/s+KGEMsOWz4vIM0FoR3w/PTdpDQGUAU4YjWMoWlmOiiinGcjc49vw3p2OiS
PsM1tklHlUdt9CMwX3uWsCeWdy7oqX2FGHpG9omg+qUpr8zw4W7YEplhRpLZCRoV+RkpM3PajAgq
CVhC5qP1MWRo1A5s4+aTraayNFQ6X29GwGV6ls+D3BKE0ypOsMz4nP17i4R8KP7YRncH6jqho+wE
xopuwJqJ7gV1xb8ZXhdu8L9usUUx1zq8tW+HvzBBiZuWCeBLgtObS6o2h1wt4pZ3iXkFwt8UZU8p
n4j+EiyBLbFvbaYNWOfxvxapOShDo+Fda5xj/j2zWGPLRcc2iRnalCQ3kzKif/wwVuytxb4kVB1x
Xo4Otwibl2XlkT/gDnEqI3akXeG8VtRm2ScyGzCHK5XL3hc1vuKbRXadMi4czVOhBN1/qwUEPokt
ipmgBOGJRsVAM4Ox+8L0E+oAJjfOWu9od0oKoIWG4x6XD/dtOGsvFe/mrxuKOQhaes4THewI1FZN
T2wnhQWaYZVCl2ykjMQ1lr8T3FNoljT0xp8IFCTu4uU9mx2DXtIxLMBKZoaVRvifXA2I8uv7K+fK
2omjaPrSNqzXWy9OD7RUj0zqpO3fHWUDfXcLvvs+cSa7xRpHSwG6vZYE2L5tcCtx9hMJRIz6KXZ1
Lrw+HvF2t5g7AwUL2GPB4gwjHZnPucvY5Sgf2PI+GvznEVL6XUNpaeqwpdfXj/BcySxTxlRYx3wJ
mxbtW8bd6PHoB1udPwK9lpJJzWewtt6NIlTcP+WMGg5m/2A2yWagsBy/YMm6GPQ+XnywyFsLLD+l
m/nXzvM9AVBa6iDaOfSKzsm5BOjC5wBl/bzdH10lD+ACkuFN4dszIkvAZAAgBSxbA7+DUbWJRH7x
1MvvyNgWwV6rbWrCXgkGtbjVjDCXU2yjehZ5EDVRlQf8tEQHodJRlkyybYbAw11zwdOo8fKb3Wp6
wteD3hHkFmJ1TrwTs6JCujW4YIP9hnfQJEfB1Jmlskvk4qpJZRXrxPkjRyb8x30wqyIuWTSxN4cj
3yT+zWQ3twT9P4D9krkkoZOqmb7krbS38LE4XVrXMFM5cn7QsAADMu0Rb0F+oRAnxklYIhq5JcJn
IfZuU62O/2Fyouca4OLY/ta7ZGxHm+rITPaoidAYCbBagVQcD/W0gxVcKJRtJA80V0GAXQOnKtx3
gMo3fbOWPv/IXne/jzYpiTCLEorE4P+SJJpVtWzvjtTmocKr3YTZX2Zx7QtXsCPQhtz99C5X5Ct7
nrGDpAegpURiKhjY+elLc8raNZIiCarDsesh2Sc58Fje8EbpG3+0y3oOpJOMMfRqGZ6Y6fsO/T8A
E96bh7uYXFKFVnVcKFwwGrBlhTR2w1h5rPXb3m/7bEvKFaLQ2WLI7Z4bs4aEVZi8PFM7BEQmrC1D
5WLQj5qCDnPr0bwTvCySM7BuxUNCu5zZuwKBWWgEawqD2NZKsMLa06VWEtZgExJa7kYzhqYTWYae
PNKfwoufLjQ5i4XR3wrkpj1g5nJ6Y4vIkAStAr+ttzNCzB/xCg253U0AX1+KFs+Ex8Lb/zCVFgHr
4UZSxnLLTE0KyAyQhV0R5WHQIqF14PFFQwS0oAgm8EHRAxpE4/7O9LAouxF6iYGnAIEmA23bJAjk
ZPvNBI053/48iMVhBNYJJDOmXBGIkoFG7qRsjZwul2PMGNlREyRToqUMeRpb+7PI1a5WaeGPMeV5
HFFq2FfOukNJqpRnK+bWQXJ3zh+gLH7MtaS9usAGPG+5v/+vypuLiN2B9Um54Du+5Z2ofde74Pcn
aCz/EPWjJqyVuet5IsctsCZELp7QSCSyu52NyzocPSc1XcWGiGecGELbgb8s96oxxrw6jn767am7
OfyHZzXxnr+Br2w4DDr/7y2BmeGESpCxYEH4jWs8xyFtJx8gO3umuzOoA80RcndXdlCSYwo7g5WY
SrzCE0P+m+pWWEqlWOq8UdGR0irwPecn/8l4mox0ZMpneMi24/01eQG6pA+6T4XDaKgOCiThmGOO
TEmnuZ6w0ws7+ZbNDp9H19aQLdxc1Q70YaISCvsKxymaPOyFRfggfilytvcFaxYo/UKmn34eX28N
c7Bqt4sgxVw0WU+ZG797+SBtpUPHdwLTCb0C4kLjod0OBB8vY+Jkfr/SVTkBuch9DIZ8VgYYVBos
xTeJv3zVCqOpqJp+Zv0FVUzbvBgQyBNf/r039b8nQhc4JZmeUysBbpMkKIfe2xa1cfd44aFzrtao
Ol/qpIpDm5svWYMg1uIN3MJGAV7Ztskge4TCuTsZjnHIX5XTwrDpgwgk37aq70xA1iKrcj0LZIT2
CYDZ7WRB4p1ChnNhwVHqmFspdmVcJtFXXg++1tv0nGWZE3+ymavBSez7tz7gGnCHm/fLHMSEaleP
lolh/VbwQyBh6nSPv2h8FrtUWEVc0Ln+4183J524VY4zNABxz56uElw3ffjZA2cTIINwAk+bC0eo
UyEx6gBINXopWiFwCvxg6+uqdxqYnhdu2uxda3Bb3uUnkX0uux8JfocVuyuMnUSVaEmhPCnfB69H
hjXwDk6UY7ilwykoNxSBXOKv8RBuHImGYNIZEWKrcAyfhFtumOrlaorbktsWOLtMW7NTSjVmenbb
FHiSe5qrdkK52gHXGtJOtaU3MmN9PUTrjsqzjeDbnGipkYdkNbyxssv/A/66tQor6pcgj30w7urI
Ez/mUUkRa1QGxxh+cp9FaUZFUf54OWKPhcJb5QEVPQjQByqxYkl7JwSM/0z3/NPxARR02TxxzxRZ
mxO5a/yaPmuUcGqNH9gpFAgpT467jPQyhvsCFxX9Gca7ig2pMXbVEKnXhUpQhWQeJkJhnBMcXQGH
5eInwYct5Bwa3YUBS1IvTDzzYJZxxPowp8Xo0AxKlk+fC99wO2YerC9IVY4/wXt5GES3WVyUhWBM
KZFkEodYYWdj2whoSfDVZ58kI9yLtISW59tA53SOq+thMmZ5QC5/RULJO08MsKgPbrS5bPzO3SyK
jsc/ud5HIH0eOEzwD6kFGeAefxUy5TEyt6L3wi4ZReBEHbEDjYocRdZKbVDH9uRlVjOg/L5qq1cQ
spECnCTtuubUwUo49/z1EbxJbIb4CZKWhSMpvBgclUwo48UA9AfTHCHUoORWbJm95KHSnGJvJX+l
tTgWWPLTpcEdoBy6JWBc6j0s4kxPE9iU+jaxIctiHOrGDsrUbeoo+JNhw2NBPEv2tlCB3riqsW9V
95ZjR9qMwgI83TPp9+k3GZ5kQqAJGh57xXR5O3TriT8SGz1y2RIbqRJ80jxI9G4lrgomNuxT8ECq
DyrkquYPnYn/WYBvB4qdwuLu4boUO3FH1qIcV5qJCe+/X2aGJs7Cl/JkNWDR+/CDKLnhK10Jdxfa
wbRlExwIkJDrSwphY30XTHmV2eJ6X/VilyTFGbiHCEy0auSuAsv0z2owns4tgad94cYZffoajj7D
BWN7DW0m05d4oACsOabC0ME2E8m4KjK1p7B266kKiJ8l1UJZVvquia35w+5cX5oLIcYwytHCxJUM
snsy9E9EXrI8UKbmpae8/UACSrAycESJtQ+NxqgjgF9rZa0fKkosv3lYMnuZbH/puj0lmeLxeu/Y
a4ijsbJAFYxhgeD2EI/H2JBs92EGOxtgT/zZjyLQbTyFZ4ZsvwQTHCrROFaZt4eXt2txi7B7z+qp
q9wgLq2WticR0dNNLk2TapQvMGBjVs+g9alk6+DDQEeY1TOKFMT7YHa52AnjiY8hE9LeZYVvkjWE
JWnnXS3YbVjDUVNEv76g+pVmnO0wKHN3ymzv1tGZwJm5LZdln/fQI618SKnoop34xO30qXI+2xVY
74ZFAwR2j2Mjw+CuVEMQzbhdTOpJ7VCANIK0Q7X9n8gTNpZPBodU0xneE5ctEJB4kp3I3RU6ZCIg
E41TV3Q9FS79BK5ddJvnphFagKZ4U7Ou3Sb6CkM1NJIPS/TNebfxUuu/X+1khr3uzvubsIHAbZTI
grQXFz8zZOJ1YBtkgEvkhk13deDL3am4X42ejwtWypJXrE86Z99Umw98YV2Tzu5WBviYUou7Qu2r
w58EUyBaOG8HS2l1yeuTd0h0EBuIq+lqCqX5zUkA3p7UDgQMzlGEQj3fznoHsBPRGaI2goVLnGjW
vco3XMxQEaZq6fhMVN9eyYbyZ8fffg5os0y0keItK516isp+yqhmZ4yjxDlly4H6pVgovWOE4VH3
UhV5aBaErVqD5I8/mQF2y8mDNWeA7ptZJ+e0mt0C+T+U5zEELmhFkfGxhmRhMIe4SR17xszwvus2
WFnkIRzrMUY6aXFTTN24y6cNhpaBL61jOh/JbZtNY2XMqMmVzAe9fYuA/4NL82A107cZFuEd8KVi
KVX6cQfyPVI51zP+Ve5km7AezUuTbhH3Px5ClW9rmntwJ9yTaGOeM+//1FLem3U/ituHqTggUrEO
06t1uVBfFzOf3pkAiQ1jrsOoVzPIuVv8WRS/aeI3ExGhBFknrPb98LDcgHt3I/F62D+QP7UwFkt6
0YFGsI5+bHejx8bECScfgPWdkrKekB09y1q0Aokyz9eTC08a7EkzuesiggmEkEpchuZ7zdmvKtpN
Yuv4vaHSvhP4uRUzPCc51QFUMYEx+O14T8Ryy13qBj8vQLzzMLRNeTW90Tm6WZ66YmXRyLIWAIZ5
vQuxe2ZJ08kuS04YpVw6j79WN6d29wPKbGi0ifDPd/n1l4FTDZ3HhzHRBIHUe4HZ3QOv15JySw9T
MJR3tLHxeAw3D49a4iIpow+a0/GCGJ78fUzBVus3j1fD9VEVuNBkj6jC5iAZnNT2hJR0/WheVj0T
OdJzEt0QbVEgZthNO39cWmY15C45uKnQVwrlsotWX5n+q66UbmF0fysRNNAd5+D8w5Cgx6oU2AZp
iA5Ixy0DX0K6fujqNZaCTAQlqRuQkMkMAFCmTUNY2WhVYMwEslLWxrsI1KCAyKFDmOkJ12PNy7nH
B2b4mRetbOtKVdo8q3ZJWZuJvSwDxogyjxxlaF5uWPseux40DUCKy1Hra9XC4ibTSQ8DuT9KTWTm
1k9jEV4obeSCqOYcunHZ+jPyg+mYGbIcC24Pmvw4e/RwOkH7hZZN6ylOoVwfWaPI4Y2+JAN/dGxo
+SYdqYqsPKzsbEflfag7XdeJAoaYxZYf1otlixOC+gqfV/vsngC3rRHHyzT/D5dPLrY6ctOvo5Yx
fhXqSvKbn9Zn4I9qNqg0JkUjsJSGnHiPRM2oRXXChythJQgb7fbL7EoEtcg7QHacCN5Wz8Nw++qr
PBbkRRE1ssKnCyFalTN3f8u/HiaBzr4mW7D6X6+IW1xtK66ScoMLpBHJeyxarnWxKV9hEEkJMpc7
Sk2a++1zwzAzpWsN7KMC10HSl4M0YsljNlqaek5QXJ+uaSFipEsdK+oGPYuEBIKsmaazas54swXR
MYuMBpdT5mkAbjiLw3nMp3ODohBP9nIkKJuDUgmxhyrsBO60GrfogTRUKqMcmymZoRVF9/N5pqd6
66oWWwa/q2SPaXqiJvtuQEVweWblNrJqssw0K9+LuHZUvHtujrPJZQv4SCW52a3ApDZubYkXoLit
rzIVzTatAJYVKBF0F+vjavXWGWZBz6g1X7T5Q7AU6xbayYEGHSnfbE4pN5HSgTUpMwx5LvomSpsu
L4qkNrFiQVvKJj7X2SRPK8AxH1vuektNedwgPpJ/VuVBwLmkUnyca/Z1+khZ7ZAGkGZqjRcTd3in
5TLwWYhcXnIZ7X+DBcf5TfY4x323V6odUxYa32P4T9nC3YVIDYhj/uYL+YtgYkJQyUwjZM2PNUrg
7rk3WLBn2052/uzWDyVE1TLwEKMIJ4A56giikkLSdHpvwqMSJUMXaMj5mX5aQIPum22ERT/keHTG
o2cRyaAoQ/qU40bk93qLs3YXg4Z9luLMbnG4jjE0lY1WU2yYFwb92fA6y7fSVQNJrMhBRvb7EgsV
uNyd3n8uT+jeS6wCV7kL8hD/qYOhYUeH3FBciwJ1pXvvVmBZe4R8dRskbtfF9FZ5bkqSfyv7zd2I
Mmp/RTznT0z7hTpNHAI4eBd95OKnSFwN2OIxV0Rs5X2jhAsyfyXD5cbD21IIzLA+dXrqKtHOAcMV
ncOrR2ofS5d/fQ7poq98tknLRsPnBn3Kz9riZSRXiYnzMeImZUhDx13boySOdIrBYWxS5cpcvN57
fvmzSzWMHZpDogyGN0r6uO6vWriOF5upZxh07IbrNvYqSvA8RZk0zmVp3xQNUodAG6A653pg3RFB
+JB3xnaTzuO7K5CmN8K0j0uixBn0XD3tgl5lFwcSD6jqi1YEIX8ftQqLjzwHIyuXKpy6jCg83MQy
gUjNcryP85dDe6BMLpgTWhQJY/tDZTxBE2kuM6vx2jrIASvHOAqfLSQ4y++aYh+xv7K1B08NOLkq
ZNYFFsT4F5Ibi50H+RZH4XCrAJ2mbUM8yTFq9LwnIZI8JgKEfRP0888Z+dyYGI9nL+ZFUqoEJksO
Xh93lnTB/s2zXFkLwbbJK21TtqkJ3pTOi8CR4Mop2uaPoNak7e9bHBBDk2NIg4XKICCJW3u9sMs5
a6hlXZ5FzRyPOTTy5nxBBvCWQQJI9sdqre0Itrz0+XlqiBowj4l3zGQJzGwfNL5a2ibKRfc47mZj
i2Kal1Owp+P9w/eii/IsuUqB7k9mtbnMMtfvTD06nSKQn9mJh0eJvemgJYVM3eAh4G8rDE4Ci5ez
S0AceY3cMXfQlV01dRDepGhpiyvrduYYn8ipnMWlBWXT1/Tk3rdP4QgkQ1TqL9dCU7kAUQRGYtXg
FBTiCnkZ0FhH3OxIsi0qUoWyYjXtRLP7hvB9JphLWDv9Z4QKqoU71NQ2wgKAhiyTjGMZCdqoxc+n
gvlvPs+4kk573xr3Skb35dVKbtKsYk0p2LJ9g/KvuKK6snL0teP1WpdpXX2DJ+vQVLKuFLiRd2JG
9GP2Jycloty/0uK+Ze/QFMk/lpG11pIZG2QJExamQ5rdWsBEgtlWAxqEHkKePPXTA1YD36YSDG6L
bw/iWIGhVVlNu7rwFWZHbfpXBUCuHGEDRExTyMgepKBs1lNlOAvZWGLjlYceWcLNXs1ISXpt2amu
MuhRyTdePQ01pUyR0sXovSZwFA5xreKvsHhUzixmtgkROqnfpyo6E8Gk+rC+6PJlbj17YG7r0Smt
avEEJeGbd8ygnvqYL6nALhAJotX9g5z4MkO4i3gYqXNKJ4HxGN7x++H9wE/WVCz+i1Eiw89FT9U/
HhbocCEbcAnf5OpFX42StZJYCOlNDlJM04362FPZjJajPa9v3T0foCZK89imPbOzxf+u9jJlA3rw
5mRfmC+4Zfbx3tomZIw1plyI8qB4kl2XaxwSFypmBgqPC6Dlt/C2t6FZEKUYonMdMcLc8q5aUx5E
pEZxn/3+u5uWEiPwHM2cENgKbTsGL20/9EENVFr0VudMs7Re49wyjcFPyL43jqLgpBhkl9vSFcJ2
5bKhHX6h94n62yy0jA4lUsR/589frcg2bfyW1GLGVsrHNIad0aiCbUrbBapk+hfSGGoGbJW+JtMs
fTqcYpHS9s3lGDGMQ9tpHDTzZfqVM6u3NN48hEIQ/ky36+k77DKTrgaOoK11mfncpwapsG0z7PRw
s1C560aSszhKXhWrfxcKnbESmbif8YCbnKsm3LB51vPo26koyTeAZaTBTHT0g+gt6rEDBWN8mSPJ
hAENqpEg9hNN8iMpxlzIV0JEUMBbvatlcsTjDXEClci7Qu/I7pvfRC8unVhfXJQoD6b9mc5IxN6J
tKd1haPKO746x8PblV2aAb759F3ICiX0V7YBBoQu/i4+6UomFEnJxZuHlyDlEIIv6OnFfw5zlPVT
cikJwyH8IbwZW7Wdze7VDPahTPw++7nGghp4guobX/kgqjeaL8ZhD45Fu8rzJIN9Zpl5qEwCBNfm
piGzqZ875vPz6IaOHikduAZoYAFiSzQ+vR3TLlWtsSW24ohdiE4iF+mp33LIF2CVZepijD3XrfV4
XDTNS+5lYrqiY+8gahy8b3hrA2mJ+PpnSxmSiMyVld+8DAB2MNC8BGo3tCfs41k5lTAVuQvnMf9Y
2o1xjXioQXUWderolA+XsNDTNRXqWlAocHm87x2uuCUFOSc+8o4x5wUIccQgZSiDbfqLJzX2+qSh
zk5DluWl52fRs0wvjVkv+9YG4XxeuZqgi/BZwv1Q9JK17/bLC+2p2aTleeLaCzdsSlUI5n8erNba
pmGDzZ25ckgWBln9Vuu4QaXmlNF966YqZP+3C/VuH9CpJB7gw92J1CnnxUTIz8CxEqhBH1satjSy
Weg31tLBsgEqjCRazREwOL69KDqU8bOfg80U+2bR4wplCsaeImJzSo+T6T/xNloQnnD6q8xQ1oG0
5S+mNr+88DGs14g8DoHOv5AIQgR50ed5x8RWZ2UlqjxwsNlp5GFn0IRs7BxpumkzzdC9xZmeZpxy
iMvdJovsd1hprCQOIZyIvSrdI/Dg/zszz8BGp2gqm/Y0yrtA7DxlmGVxkFvrZqmO5KQIovn8cwBo
lfreZyrOF7hXcm0tTSBbfqRRf1vImE6jtAtDHWFO0dGDW4NJp51fLcwZmCgD3IQa3gtvxf6gEVYU
GutkNgtfbbrzGWRIZ4TS4EJA77nq9n2t1na9sntftifFHgu8PB9o/vBuOLGNdbJ3Lf5YWCuG3r4C
lsmGZcadwjiZzHyF+CCUMIGBTvWOsrdEPVyF31hdGn70Qegxm5DDN/UHiB7BjQMyFC8I0UZCQi/O
qRn9W28baDPe0QXjPA7/NVu7sEz0NkGuHIW+kJnSwOE1u+ZRrqKwKkXY6PCVvvVXYTVePsVWMQOg
mHD2pWCM5fkSdKikJS35BU2sCn07IpiQPr+LifQyf+82Iy86SQd7wq/1Zll8VG/IoV0WQU+G+UI/
8aI4U5RrSRpfJOo17F6dC4ABUxtcX2rvaAreDZ2f5Mi2FzEEFOeUL4y7rO1CenL1XAbwPXSz2G6y
8irBtwQrAyEbfRa0qRdGBMN27cnmm3uVENMBt3dNTZ0JVHIcshMI24BtzK8kVJPn0X4ma6Tva173
Hv4QiATU71I7rOOjMCVJtzeuxtj4rCwrpWNefVde7Dci9h4f1SxEsUlsGrWw8Ho9jV2nSgUqCsQE
IbxIsa8m4Xf/GnhOfvMBM+BxEawKY/0hHEIc315lmXzny4zEEk2tg10unAxKRmTqWEtMtSVZ6Klu
BXcZq3/FUrPQSOE/V1TfNclaV1joW+2Xq49xofgWz/WN44nkGVMtKkEMxDOk7Ap2bR2a3OyML/BX
oE+lYgPrUWYmUQcZiBkg1mFKXbEQcplcplpbzZwmcEcO6wD44mZCl35nXrXxzAuFutqo1OO+xUeK
iW9E0wnUF5OJ/TCDDYQrsRLpI7O1ArnLS1ajUXJrYtyYJVQ0g7tHc1beyASPQ25g0rUL2S8nhpYm
ZI938mQY5VKVsl8WNNp6j8DImQT0lZSXQNYZOqDOsWzWVFZdZUotLhWgqFKGcwZsZjMcPPKRgI8g
S6QQaK5wsbCyE0HDysyGPFyTJbjJ3txZ3N94nOkqEo6YrxNulHM5xZbGwJZwDgPMkxXrWH3x/VOV
eomgixj/5txUIPg+8hhtBUtYf+BKcE4JxSMRK8i6oBQBAA7RPWRwkg4twI1DspDA46VG196yVoOc
3Z0EW1Pvqp9mIuG4GRMou6EUJ5b0guWfELFAPMzcr/NtRKkHja8l8BuM+jO8gqKg5h7zCmSsxOcg
NdsT/C7B3Jz6wlhnq6WReJQngoEQSEeLzzADvNRIWJEOkpwdL8rrAcRAawRwlRAybyH7ulwhspy+
DMJQTJZrDHSaOb4o+uf178n1jySLEdLIt2FweOz4Zwp8E79EnY6iLr3fYDcM9VouKHdqX321FUVB
VxDjwEI86/O+dj0Gf1y7WWX63qGkjNSli/TDfT6PKztLdq4qxc1Wba1m5WaR0YlEv80C+XvAAaDC
p9lb5ufIQFNjh4+pgVi8bqFSaaAAKaq2xwJUTlUxaDgHnFOQTINm7P1gXFePcvUqHZFxRSjgV6bY
Vx9JJXgfk2CkgRdH3JR6PMwRbDuWNZYeBhNCvwO6jM5ecX7dpXwEZYj0udeTF3KY7vG+eZJc+use
Akhw230BAzVHaizXOCd7lap2H/adVteyd8o8BVLmU/q8i/eiFZClvUe3WV/ojrcsA2VJQXXqGjEK
xHWbSmu0GwxkytTOOHyAU2YH4WqMUcFN3muAA09q4QZsC2ufnMUtytPyDMyr1XXeHyzSOGiOmbUl
JsYw0S4iDeanE5AQSu7IC0C5ZsONLVeA5AMutxGJVplxYg0gS7V6fyQTOZGBp2Bu6RzIqBc8B18a
KPbkKMw0ON/WNyd818NW0G7Yk0APCV8S2AW1A2jycYID06RYyVvLkCzuzul773lOvQ09gyF9ZE8k
F4Wg+DDy8vjUtuAnGM6bWxeV7L1CDWLHenNiHZuUyZBJEQCDQ0bdJ/fAJWjscbDiLgvUDSvjvy76
FUZI0+CKcVh4DsEe6WaNXmmT9xd483bl9i+9Am8zFC3zYLKS2gXerEv23E0eK6/dPsVjDkgrZSw8
uHgIYcb3chjFrgWaOdytrvk4leHOwWA1FcRQP9bkPeDiP1sTEFuxLBsIp2ckQpmmMjees+gdXb08
S4VwCuAb+xz9AG6nxR5gheAfHc+lMdAXNSAbfz/NgSWZzRvcvZuA63SqYYpTzMgJxkJqwj1YpC0a
UKYyEKeI8hVriTOQhwITsz4/V6ZgRpcjmmruyMfr/2BmnIRuOd1HY4DDw6cdu9qzAsJbgCzxwUQq
f+ErrssRVl7DR6iy1AZmzX3MdNFKd/IRVe3w9kNGvZqulwMSnzsWRvARa1pvkZCAsB3VAzIggTXe
hCa5tiam6JWPz5k0+kV2Ixx7qsL29TJXdPT6Jgixqg47kED83cxc4KuOwa65fG5L9aVh14f4kNkM
2dVHrmZ1+K5jCFdmmTsaP26YH4DO7jfegYtKyBu6CHmwTGCaAATECEBwlgTG9PjpjwFthf1g2j1g
eqHVwXegYM2kkyLtN/C+BNfy0f/shfpdRQY6Lg06GkXoTvxhPjiMaBcw3MIOgIpt4qY7JkLZJQEq
FFzA5wviRYxUkdR8becpYdTOKnE9M9BsfYMZcp2JEM/HD68zrw+CfKmoZl3x0s+6PHlyqpfB9awH
SVaExkXnCqxpHOgeFWGuphxmWS4i+M0pIYgAZWXnHFvv/y+KDWVdr1e7l/E/381b4tcEJzIYkaNe
DJTzkgdJ8ew7Fw9aQ6Sho62Cn7pcf6aOc2sgVId6oNwbHkr22dxgcwH6gu6w9BchwrjkerHvsfdw
KIdL99431bsHsIMCLsAPxDmQbgDz8V4lEb6tevp0tku1if9sjkVo0qHg+p58/GDDYWUkp7Lrkl8R
BGZEIgHQwUBmP+YtmzsykTXxD+A5n7qFPVtUxqPCUge8eZ94aUqGbm/5xpezHby+TtrdoBlFaHeI
araXxYKH+zeWx12baOQeABkMvpueDW/qAohc49AfJmpamsLGqfRy5cFNrD0qWkexek9Fizl7AeMk
yglZMhIhxz2iI1/zEzj2ggySi/Gx6fUzVDC0dLjECYU/H7wT1X84lxbiyAb98CZxkexJGp6YQ2Ay
mdJMAEiKEo+MSLRvZKYdPB7xz7AOPo6bTOBZNuxQaodZhcHVx77iplEjjIFQe66AKy6j06sWcz2r
AVaRqqfqernzRFkhuU7r92PpT8uueISxh6ANi2QE5EnWi2KYAmutrcoolGI5zu3WJlePfq1KyqNs
XVza0G+sqpMP5sPpQu3x8durCF5LkiKd+oaEcq0zL2+C+pyt8t7JCwmMnRAX8sdwfeYQq8/AV8qu
EeHs2as9vL5R4axc1wM4ToVoW+/g4KQhdsxpPJgC9X4hXqHHR0e+7XU+91cOe32tjK1tO+lry029
7gOee8O1Jr4yE9EQ4QqpQlqMhrHhYzhzz5kPYi+rCLp28nw87wqEYh95AQVt5sIqxvzMHrd0B+54
0/Ivyg1szUeCKw4fcD4vUPDwOXEkt4AAhZzrxtWwNzT+nhYk+SDQ/rdw8Z/xuYM7K3Uk1ufKVbWu
O9oHiUpQq0bthYI3h9lR+TCUunHtzp1/8bXxgTuEyXWnMfT2QKU8DdpN0ZzujGOr3ihPy34AaFcr
ruJlRxSkriTRxa0Hi1PEcrJm0KbaqbnRSCmALcVjud9Ul3KhYhUBifEcaDap/t4lSA4uz7vOhKdK
YvC7AjQwW/dpLsYN8HWUgopA7tvHi+Rhu5BwJJ1iAN1WVWmjO5tapfEG0NCU1w/9M9EUnxY2nO5Z
bYq7oQ3W1lp1y1SG95mkpBICCwcMVwCTF7oT1mMBLzIk2UaZwbNrzfTUnI9CpEup/tPNO3RfsCyb
ogoLItc9LX/eeKXF8Ru1iqKYJB0SL8cLmUUazKO0bo+lhUoDffu08WfkAFceHS4fS2lKRhewPWrQ
ajMtfPxn5i2Z5CVr6HHIMJX7YDv9/AwPJkjR2kQJLAkz8HcpW0H87L8q2+DWi9RKNCI9CydgN5un
E/GLarEg8w2TTPqYPwK66ts27w8mth6rY5Im6fgIXKODRiCndhnHBJ3Xhlz5ef4RhZLmND4XTlbc
ym8ZmUqrupQVSf66gSC/xub/vO3lpiBEAKQAIA3J/1C4+FiZaYEkuyclfJEzRm6fFqPrgiXVm6vd
dd6XxtUD1bdzYnerJe6JZY+GTtnWonIiddBckiInVkiq8bX5fTiREF5MpRlKkw0UY3msAULCFdO1
p9wh+OYN7+4609XAC0OZHpbq19am7GoTBkzcPNPTt5Nxxz0OXKWUn3yUkUkSZjOYJ5EOZSKI/HFi
aoop9z76qwD3otu//th3uW9yu0bfdyJQMJ8lCI4Jx55pX6RoDsKGBPeQWYwIIfpqcwKNnDm/BlAv
ylujn4iFzMu4qq+V8e3UKvYHeWtnQqH98eFBrKxcrob1EG1ftIRihZZL/Yz6h0bXbBXXwRrFVlK/
h6J8qaNIk/x6xemokoQxkOniEBTjoJsfIt7OY+dxrhHQPjycaFIqNntgP2bfJLV9dpeqX2PIPd0R
TMsGdAYuaSazlfGoVTBs4L6oO0IW0cm8lJdK6VC7kO+RM6kqYoCu1Cxb4wWsuM8+jyOxCRqVWX4q
YYxoJiiif6imuFmmcIJES3hlEjPjKlcvhNkm7R3DSOr6pMs25zX2TaZhg7mTfNIQ/MLlSyLEMCss
MBGIzRzxE08teFN3gN4fAHTomvLWeBqjxM0xXZ/ehhyrbO+ZRk3E+0uec6JzlhkQnX0nQ8GV4Fuh
JmW7zzFDXNfXb1QgnEsQZeyVPUrtNbf8lOsbxFG9INUEc0TuBfb04JKCkwJ+qWW3/PPQlCRLZ0P6
o18s6Jje570lETwSf+qPXCqDyFMOUarmJrdSyh2SCnjrbZOI43HtlcXOCH5Eu2H41l+RyS+2zPAG
6HlB5+C7RFef+8aPssfrT9hNSf4tTTmtc563RdBPiQTh291kX2etsGJ4KEO0C4i+fmaY4DkDXs71
WOPVzmwCaiqmyq7iWDcvl4p7SMZYxbGzz4d/A0zN+6wxargn96GQhaFnBbVLhUtlSoyGc0jCPBvT
SNfURfM+HQcxRIygOd60njT7r1iPb5uUipBZy9kEQBNAG9Cac2On/GbKEKO5gM4xki4/mTAdYPRf
UPPk6AVns0UJAnhL8qUlA8do4ZPlkhKVxNqBPU2odj0NA8zbD4aROwXKz9zra/Y/xWcgrLwv2yyJ
Z0ZKd1jIbS6U+VEYaZyYCvgMSd3Td1aicvjL2fh/oZ7fy4p9IvGdO+6CvQyTT3QI0vBw1xjREt4e
CK7RI5pd+NEyWeygHi52TBSOvphetMcIz8nPGVkrHevKYF53D+7+23QXwclB+jzRycA+z5bL6saV
nege+yVqd9MghA+NoJJxJF0TRReTpNVDJDhO6yKT/cP1TD9RGNNc9ODT8wznhr42vgdWGcrrw65T
J0xEeiBgMF1lwCie+CKm6pEpV5xDg+C2zaptLP7Ny5wuuvNGXr9ZqF28vuFEtaLiB0wA03CxhAmk
EhJ7G67uKbXAr8ZhrTcGrnkXx7bZP+mbVlm26TCjkxODahUouaJIGlrgJS7j+sENj6OTC9mzPEKj
HeUt/QJP5+xpBzQt5PmagUzVfoagxaDHzYol1U9zS/Bmy7iZy1L6oJ1l48DvD/IOTznCRL8Y6lfp
0ZLj3lIIQpr+ORABAdnSqYEHHuMx+9V1UJ9X+Jxkhb4VwMAtCS3WFW7neFl0fiLI5/c0Lg6Egm6G
pjXV6vXO6d4z+5FsDWI/kue7ReT8hKkbY6othE7A+Ee4MdzIbh5NCrg8mvR3VAhc7P18vczQm8IT
tt3U8DbozDdpC11SHWU+TEFRdLCG5CD3o9UIeH0/ArBUlWQAn3HBuJtIBV58/BEArEFz56+/Wud0
vKMrFZodiwIBFd9mJOEOse+uclVTK46Owahb5cERttY5YhsvWH0fNEUCrixoUg4LjAYeS2kSyPlL
TslYCUS+yYGY6htPqXd6HZEd+EkMOTfWhQmVP110/lgfteO2ix7YqN8YJLKjVJuhBrJGxvgqhupp
k0CO/o7w7cyEepUHXk+h63XFOgBQ1NqZzHZjVCDa094tTGfca/HLq3ZukoHZAFWMzVuQa4fR9aSu
yhFrFS9CYixoR96vI/nXSxNbVuRhOC67YFZHSxcY3Magdpp/VHyITlVBOFxVsXbmHfs9ddsS7oOW
T16119DilwBQ3snfA/dDE7D01Cf1bkemI9e+Av3nwAbzNiKG333YkrvgUIgfqGloEnaes3ERp3aD
iya9DvV2cQLZx1aSUqzTam4QlCji1k40UPABi0YdxvXocRGIWK6qO8zQqWOV8xhBQ7SjDH3jz19K
4fLO+yzkmMIpw7BEYKceNSZjHk0kQXo+5pPegxsKsPgl707Fiev4v5PLFuVL//RyQ592Pouxqsol
7+0uguzHecY+2NuPDx3XDb4nCsvjzC6GyOmAwTK4kQ/OndVSSGw1aFYBpUn3uhQd+JX/fFuTfPlQ
L3GuEzMMS5qEZ8nLhFFi/do5eXhYOKoZrXfeNWdEABQI3AhqEsf0I3ltENpgTrjUs8e7gG/GQb05
y68ew+/OTGB75T+1os8QwjNGGDWIjlE9EjLgD/qqAG60hJBm24oseftEtw7llBElr0WYczUMDC3L
0OsNEC56foTEjkfQjk+wUaivcayBxUN6MNc32mkR1t18t9WSObjt4cAjsDHhAuu8jPQsfojHAQTx
JQ3pAx5DWBfhF/e4UNTBSfTBFhRGmwFmJdDT0a+ipcQVZelubL7Z1col3QcjYt15bOlMfSXc7SKA
Q9aqamjBAV2HAhHN7/mIyUMR6bjHnPLbyTyqyoS6uUQ/uC7bPzfUwB+lvKx7WdnUIQhGpmNYy1tT
AHmcaEH4/ws6mnpvF84m4VudVBfky+QcbbZSTaCUm1m7GDquGSO1WC/L3uabcjAqe9SiSce5gk4Z
WHB1lbkLz+nKRr0+ah6yDOUruuKQV0XwwfEkAE/GlKrM6axqGMkuwKkmRBfHg9NZSeUrd4ZbZhk2
zMkn82TtZZeAZ989INCe4k+2mlF4wBa+9CwIbVRSCF7jc7I6+FI78AbyM88c1nR/Hiw81cgP+3QK
rVZtJz5zaZHjNMGBBAXG1fRcS0SnohV1txtfuSAzTwZfPwhxV7u+9PXlQOnK3/+toCmyJ4IrphXS
ojmP0cqIuUfmidTrA13rDZDLj+5yiRxpamV7Vp3V91xx1JY0jDRaKkBUsGSMoT+ndh+rNgsirdKQ
VYwU1qvxH4cBwlvCE8tZVb5GzKPRgoB7tTsg/7ozebnLTWsCg36JQjMWRuW8f59gXwvZtyTCCSqs
IgDiQQOR5MRMpWQkyZ611dylpdd/qFURLo4+Tr9lJk1WHtGj+bbuJCmB0N5WDRMHV+FfHFp00EVC
pqkmxbKI1crswQ7JJmAS1Evs/hjaP9jqcbkArKuSmgC6FulXZWVHdnSSE4Ye1wxRLd7R8pcc89c0
Y6h+fGi4nVtGNTHgkkyK/mGepRWr8AR3CZBzm56G+HdtreUd2AuNfYT8Hjq+s1Y7Iq3mfQJqK6Cr
E4XRyt+UTHsYDRdgXHWMJKJb1F4P7fXImD1jMUu2j4Tdq11wt7a6Ndp52nxG+1ESfnGiF0+XsKmO
NwpbVJ86bcchAnoah0//O6W7rgjFB2ONXP6PQCCWvtuuhjAXOYV6kqT2eH5pn6YilT1MgZxKA9CK
YR2hi+fLAhiV7BdH89ciKpWDaKeKeXio163HF+DNsX4uXDzlFoo1MSFkBbik71rnxjG6WeOTCS0+
lbZpkjnT+O+/4A1PBAEETBLN4bfM0If6G4d+cZ/KgvAkJ9rBprkpaUoTlj9dnrL2SfwE9vkrBTBj
aOcHouLYdvrKMAcxEThCnE4quC6v4xQ0NMtEEHSwIAWqrhJd4m9e+TMCzAoTUidkq3NVrYK4NYCD
HCCuSvfuCJwdtYBEvUw05Yc/Q+KNWhzoQxc1ehBb82nniFZwLzUVQxSp7U7F5J8QsUAxCA2ownAT
atWj7CIBqH/UnOrIKKoOA3nI024gQFY8cWzI5ww+3+/SzH0h9/DUPAQZ4XpI38lPtEnsZ1ODSLZV
ULjQ6NvP5e2AyH/UGc1cuaOzTy6SFkeoV/1MsI2oQqhvCYmSjRIH5fKeFPlE/kfQcF00idQ+n9tu
SZFbM2Nur/LLgMIOzaNSXBuw7smy16DYVSfcI8YSDidsf/TEhBwAImEpH5s1PU/9XmSVcIzj7JcU
TfKY2r8XtSuO6sNEe7uGsQwjnoBru3tFEpDUnNcMpQx6pkP0U1V7B2Cszsa7zzj/TLFqxsPTIA+w
GXlGamZI/y4M3ufQpVoVKzzO2LEC6KjHRI1O1vEGp6VSI9mZVUNi6b4WwWDTbBcbYs2T+t/LRj8I
VCzKPN2SVCM2uGZAVfvP8cFA+RfR26VRqQ4fh9I5BLywaEL37jPaeWBSi29Bq+eUJlxE3dZhL/rG
7rlH2hSA0cKIAqG9LwwZ1gLZ8IhqTwJHXJOkJiCBiQ6Ob9m65cm7AcHYJMhxjtXnxgkx7PrT4UCs
MdFt9NdwHO89JBsJH6vwDFQG3rtjCGq2fNbQZvMRI9gm/Hs3MOLzsaT4hB/EhdNVz95Y6BPPj6Ew
AIgkCPtAYz3UuHK5IGgra1KLuDFBuUzrRySZIALT2axrssV8oXDWIjEnv3qT6EfKKVuckGH1aTS3
n+G/A4mG3a24jx0S0yk/GoLO16E8nzSxyt9Rkr202ZWjaF0UIVPc5x5zepj5WtDpQVYz/Jqf/qIN
KqE3mexCy17XdCVvkiOWKGGPJECFBS9D1otQC+VM5kbVywykRYQfv6B7zMheqaRSL8apIwAwSVQq
VDtschV2vlw6A6QKOR6HnOkh8bac833lARX3n/s1xz/YpTlG1DxQPzqkXjCRglysjnVKVEsKvYSO
yTDeE5mjvIZoQlHSg+VWGgqReDKwg8O05QZweoBHye56kgz5whEhrstq/EVjaHXwnC8y/fQ8L9Df
W2UBCHkzDUrXQUFR1oNRHwofW24vsuYKSAi6G/+4Kr25j7k5g52ZCvqK8DvRjZcBw2c1q3xY486P
zsb6WMZq2plnxpPTOE9st3gAZPDLBwir6NGAwqxty9oH6yOyMmAP5mkmFdLCJ6uaLFPI1I3kYxHK
76+MaZ13wW+fKWRoS/FNTRCLe7IKVkmIQhHVNc5ib6LACnPiAUSKltMO9wPSBt5hsN9epg98jqzj
3vvJhESHPxcGjj3S22VPgf/+lgqp0daCx5A+Ro2jY2fYKRMOETaIANCPESe04aZOI8FuX9zFg3OU
halH8KbGsFdKgJCj203oVjQDhaJeDkHCOOPM+36/z8GQ3yV1Q9ebOo+tHxwQDZNHvOUtRmr2ksYM
RTeH5kQK8Dl22zu67AzC93jgOHR4DrzsL2ux+YO4mIWBG3JLxLQ6rmexPTWM9sJJCEWUbtfa1V8j
B9teIv2PyE9cBkBp01ut/Yo4nk3Qu4iNOap8jfwBZCVbgSyW+IOSpJW0K6faKytZmeOIGlc2P3UU
O4ceEHmmDyNMPvx/Lu43iy6ceZtd/QC24yK3wEF84J/6Tqpo5nj4mGopWp9Lvjc65umkh2E8wy9q
hrst3nXt62IKXhnwSjHlxhKxbPpS2KY1eAgQq8Ps+5F9KzT1Xw3hz5B7o8zLetF9xs8+b+n+g2e9
88uwYwGWJE+1+2UeavD4m4Ia1GXYcUz08wkX2KrMtSnISwN3kuAFByOKl9yRKBmnNioFQdGOYo3I
Oksw18ZjAhZ05DVOZIbv9vkRmk2jiJrS2/uubKNKuLdLCJaAhDqAD835S7SrJHuQR3N/sfK27D4/
WvgFPcaPcCAHmKyLRMEqq2g6bzQ6OuGjiFak4ltTxUBm7eRIqW3Fwy31qCmth2k2YnHr7xGYZJcY
JEUuFqEseXD6ARFs7KLeHz+KMB/55uOOI2bROJeB///i7ySnVHkVf9JVv/gVcB1QBNWzF1104Ctr
4gWwq20UsjDDBLh3Jvcs80yeBEUxc8rGUFFtYvCacW/+wFLUGEz30QDrx5OZk1EzRhYxBD3U4UPq
F+hWzEeGLoTMQz9JFoocZ0MTYbaGE+6nkq7eXQMYqldCMcWcqTA3NCwqBMYmEGFykuCY8MujEY3v
bMCT4QQP2Wahbh7Q48CeeE4Cv+zU2lsULB+PhfxVmroBjGBuiWg1ti11MaunjAg0FnrORfe35f1J
lN0ZlWbd21noHKfBsDCMb1yUqfz4wzAiJeWRE9V1e406rZawosBGq7601su8OjHpP/kCo1etv8Kr
D59jUyQSs/qUR2xxRme+zp2mQjwH9KqTA/NI9MOIRN7O9dEDSrUaNQzcv0iygKnfTuNWRfqAVSD/
fN6iuRbZZs7BDG+wSxVXTHFi4Fruf/MJLtTVwtS3OsUz7aCIPohdrs2Vzx0uGFJkIxFeImbGqjfX
NEoyar5eJRloC5ZUsbO4ny5/Px6Cc8mMh+82CyXjZ5ivxe8flVbyqjHFr16BycjIIhOj8yD+/ZU7
hu8m5fTxfxVWJxU1CgwfeoJIytxEd6TyuU5lWjsFTx6++o30PYbzojZ0uQb5K6bg0dvCecCjv+dd
eEXs7ZgLfRnVMFhnlI9pefj13nO5E8FJIaD2AASgUQpc1h3MZTEaIJUfmDNOqwidMd8Y59rIyx+R
7QXjey9V7zamEZN4qx1PODtccJ9jl/AIm/TeGeyMF2YQasbUcCdSfiaBCShgxbgztkKPjnUHmwhH
SbqauaXRXzM5Y1xkJpt3p0EcmVh9SrZSfH/E0slChH0kCWbZBbjW0KtU+ieAc1hdTij/qdS4E4gn
KcMZFAqNAIiVHVyuX6B/KBSZVl8JU7vQs/OKirZ0xldOClGOct9YJkkUGqB7SJ8HkPwU4p+/sqxe
mhbTL2f+4jEJMuC+DlOcVO8D09sZzsaMXrmcwyDNqBhMZRHoE+tNq7ShrB7Xgg1iuaEXff36WK4t
bkzNMDzJhFmvulfAT3ZerWGeiMgmgK0mD/mguehsvAt+gJeI9EPQxECXFJBiSHPVpWdVQ7dexPIy
Xsila6X3tFR/IC09uXEfk5o11zgZqM/kx9xn0b8m2CKBFdXWR/9XjDI3DTzohAhs3r+EK3zEUUrh
ODjFmj03lx56jGy3EVfGZ78OrZp/iM3ttPgpANr41IkVUO5B1OSsDpS1Ir9ulZJrFO8f52oGmEtp
BOX5+pM8RawH87MZt/hXwxNvL04jJ7G2YPLdWidcEfeiFy19i2MAAHvEgL8wqzuJGLH/CFUZ5vR5
O3a7gQJ/cm1M+WyW9bxpjnvBxMNDFd3N41pUKQEms9Cax+r9lluZgCwZ3G+FTwoJQQuQK8qx6a3A
rDU4D6P4BJZhPd8tXU/nMFvA+JngQ7c5y3gdYeqXtAauRNJzIAOkT0AEtj0LU5Br6JVxfaVXV0xU
31F5GldycdHTKjpsUFn54CZix4iLCsyrEuJscxn4aBpMmih1+/x8UyxCW6ZtSzIvac2WaYkl+3nn
0AkhX/k8z8H59OuADbOwdHtbES8Z2WNiO/KKbpVXd72eCL1Ts6VKOyCZPw0JPMnlOuKpVye+Hlbz
G7SC6o1/Mi8eh3d/ptFxW/20NX7NUFE0ApU1yN88KxY1NM5OBbtvUWohiMuXyjBHmCW8Opwv9Bgd
OoYHGDzQTbDg4wtwfbicCx91v3y0vtg7QPehtODZc+P0WHwNyn0nh7iH5E0/TJ5VYpPQNTl+LEuf
gCEuACG/USVgTk2kuFQFaIAbPU2PpCh0FgKHNjtjVBtrVxfvSpuRh9l56HQSg+HC9pkAM/p+RSME
ngeyDRe2Tn8/Qf8U0nbjesg3r53jeNwZPuY1tuwOxnPQsfooNVmdCX3B44DBfYuigyRtE7+yq4i1
ChXT90Cd1DNfTYv3e0vRhqHdb/6EtVg3FZJX5dI5e4Mnbp2WmFTxZlUDl+EkzBzkK9aQAoRv3eI7
m+NHQT3ommlOE+1HhAKZr07YOjJMaWQ2uGTDTHCA0K8ggGUtFp3KvmXTlwPnSrovMJLgBwEp/Y7D
Am5tcAB0bsFJg3RnzlciBIAJmkydbvBQa0OVJhQyn2ghLYHSA1E04MVJCAV1UTPypNszCzArw8aO
rIhxhLyUP9lhXK+Gm9bjsMfakqvWeptF8b0Cm3dap48ImW4WaTMH4mEOQ92hC1wxaushNyqX0/jp
YGWIQIumZ/gRz58XQCZQTxiLg3PkYfkP8RUPydkgeJ4B/DZ7HnmfPtoxnbZOOo8z4MMf/w4iO7iM
0pOkbZ4FM6g6Xn2yZPWe6UUlaQPMtIDHcrX2GLJE92vfCWLx57q3D/YXoHVlqDWYB/nR4rkqs+bi
hq3Tug/By5L+fL4k4GQ87blGPHny2KqGPahvqwi2e4uFABrRrEhNQjdjgdgE+I+MuXln7loswcjY
dqTbEONZKoEk+Nm9fvEwc+du4uq8Plpj8TdQKupbBKoPU7epYyOwhycFoSfEiCb7tRdj+Je1pt8V
qCYuJ6gtCPEUExu+ZvQAHEfxaOapqKnlw4B7gMQW0n7rbfnIEKgNx4+YaE4GoznmhtqivzvnIGyp
4+x+w5BQu6qS8q5Zmf8yekF88aLLIJD+9MphQhZbLjwQYhUuSW4PzygXWv0IsB/TIwA5oPDpP0A0
Gn76lRnw0yrfOhUHSW9pd/NQyWFfaFvRhYBp9k0JR7Yiu5p//g5mcufgVlwbzLo0e5vLz0Bn6SSm
b+4zkZoEnpYj5vAQYNKTXfBn8HCXd2c6fMkEzhhWWCPs8PMU61hkc/GP4kJvnLV8KZ8vV0QWs+Fr
UHIqBe3Fn3I7OoQdwZcxXKz4fztZCy24+/Z8GAp4ScbY28hmfa6NEvGo6DvjiKjbtSHSP3ZqK5r0
o0nd1WJFLVO6SnJ8yqDhI4t3vExGI5XARwdERtPVLMy6hjWy62IVI3hc3FvHCsaEetafM9Amqjke
RL4weK7wgtqQiYMHj+Es1DbuW9uFRxrd+f6hV0CISJYNY3/HbJ2HgZzrH5lrhIw3APWxx+I5W2lq
aZekIfqEbHrWOPtjfG8bo0A678cN4y71QO5jlwWgAGdKMOZ83frXy2PsQ8MbpgurF+xideR60Fuw
MtjzDt6kYT3loZxD+aGuK0UxUlC/IhGwPMJBCIxggJmDVuMhFK1w7lNkojwLVBODAptu6P9LGs5m
SO81A6h2QM1r0NebHf6NOCw70ltB4WkHu06Nys3WgTbH776bXPf0WIvT+n4D8Sx2jpVrQSxrj0QP
Ru356wxpZj/d65dY+cOn/jmc2Cwzo8NQuDFpo0/69rcoPhXwvskn2IZWpyWvooVb5STVC/PR3mP0
wG/N3lotNvL+t9DZUcOlJpE+R8mZRs73bUTD4R4cfK+rvqaHfFbgmSok9jEaV/iy4bZefnsCkb/a
kSs4K1wPXvsZN85XFDY19tbPotKP+U9Y/MMqW4xdkANSbe6Xk5nlw4zD2HLYRKmeD2tBURzdYIaY
Y/AUP4wwsMijraT5Gr8hpARosyI+x087SLnB48RJWJeYGPR3L9EkULhZJA6B8UTv7bZ6/r9LgSpA
Q6rVdFJ3RivXAPBJeD/huPbmKtmAIM63IdE7SjkuJIRr/1B0sGIgpA7aC5ijxWTAbFApBMPCUsOg
+o82u+KFZflzWs5eIoPAjpxzXMvI3QOH6v00OrGPRtv6OYC3G768IOE9/NGbRIUXcmL65OoJrucJ
5MZ93n/WCJQOvCmLu6/xVVQwKM9fKiM7QT6mIKjTdcgxV9Wc+BRo8jyMZgERGp4zbE5mKAYgaCt2
4hFb+myGGc8BvhhU5qs/z7abxgl1k3ZFPn/vxfdpmxhLIpnLSTbYacMpfCN2AYiWS//ISRrhH2yR
MO/DQs9F1cX5MTl5qupUje+cuSpdUPYyU7xT8wzBMVsot394HZx3cNZrz6I48CNwPSVJnMohSAa6
AyWMAwIcOrw8MMuV7lpmYGX3C7f6eWvNR7llnZ/1o2BMYDB7+C+1/aIzv8tIIbnuaR1AYkLoVGO+
y7ydlHUhlQtwbwMi8VPJx3Etc3tNOt78pwSYkos15jgztPGmd6sietKeVpMT2YDDGJZJ7A8sEj36
epOepZRM3bSVWolkVOXqDYs2he67OIeCbOjc/GZ0NnhEMC6VQLlNg3RrO0uLKt5Y5asazyex8Xto
RrmVA9g8DBVvNRxpbYJzcbkEt5bFUHU5pW9zmMPyagmuScwHNcyC/zxxy/Znk9c96i4dLhKURUrA
nXBwpwSniLPxw9yO1kY91+nzbO9pcJ4YkjfFswBCYZHYIYsThulHfHqTBnaAgSil8dpKSZQ8J5Pf
q6nSYLxKALCNZ8E6Cc9h7mrLlL6V0X6t28eA2Mhxpt94yIsC6CV/DA4ilQaYFdHZsjCOXOgDAO7v
bc1OJIJm9q9oMUuDbYvEKJbP40yFmOkTpQLsJGvp9D/JhCln7rcbIV2ofcPx3VMuVa5+se7EE97E
thK0qSlpWxlJqNWX8wb7xHxJdefjDOWu+f/qgRsUsU2GAq44WMl3XPpVOwVp35/JhPU+1mnJOFJC
KO5ageGE0dmHTXfKltKECiEFhP1OGUngBmp7tRvoF5xqT/AaBT7tgt9yuPj63GDb4lOHC8gYmA3E
BJie9cKzx+wk2eBUeWnLLsql4PpSfizy7jXziYylezpVWo1bgYWYZElrp+d57XUCRhOD/bmFdYHE
lDIZqXblsJuo7cQijk6BgdM0pLHSdLx1hcyyaDcuOGuRiQLbWdjW/0BRChabTS2wFOnphhqT6UnP
6hrA2n+6MTZLCcJpYxHDLBu5Q5+3vO0IbxzOuAHzLvgmA4gw8M76ityvJ7APaApJgLpFCPlB2tYu
cBiudM78Nd3FXJaCM5ceojEBfhAI5KsFqH8hweZkWKIfjn8SDuH+zsNNgWeaAfVRZwcKaIYGgGdi
gWQGGGlQuyucCwAka/C7kNPgU4srHbLj3VIMaK64HCwNEmLuJ5R7sQ6zZ+xdjDH0Rp5A4ECG2XYa
UK7bsHBcA6ci4Z9edWj58D5qxQNBhCtODymj/0u3Js4WBlDYRw0gY7gCVrPcoYZsh9mMAPWd9MnF
znhgPrg08FFHBg69ZpwHKFK8xJ+MiteARUC4J6nGr305J1PbXVq2iKqKprw2B7O5HAf40qeLMCyD
JnpWh2dwogUN/8m+Y/BfxugD5eCXe5k8uHHUortYcspxw5p2DJ8gbQ/7pQ6KrNNHHIh2nSRHO4uS
FH2r9wEmnO8z6/NoAkRCo5Wq4PVZeb1BdrPAsCdb7sC1ehlpvKWmNkAErDPSNMiSaTWdlgep6otY
+lA61eHvJ+z9jdOypEHfHYLSh1vMwR/1zAG9UQKOa+MTH/w+7Dlu3UcGX5ARdY5e2NdV9MOM/Fyn
EnVUJx0ypRj72wRw9W321L/U1chHDugT8GOtk9HxoAc/FgANwHEOAhcmKA9+1VST4Ee3DzWwTXAp
f0TONzZeYXWT49i3smUSD3nXBBlSX3E4g5PQNqFklZiQ1SzLGaHgCe6vPAQY+5LnLCErx8ekbYv4
BLG1/dOL9jsickFkESMKAlKt3rEiZ31EtJZFrZjPbthVNn9Cfy9QD9s3Lr4e5uNG4ibs0+zXjPqJ
HPqAu+zYyZ0o5SOAtN02wAIEa2rFOJHsfYV452AJnXjwzzw8h0CR03/aCAphWyqL+upoI9XXA2pJ
4ZHoWFOoqktbBp+dXgvbQR8ZgaO3RsAZQK86Qcy9/1vK4ufzeb5GpH9jvGkhO4de3MikoGWzCVd+
YQNVNnqPhPpGYM982v69x5G/psvvtNV+Nj+3/Ga0eTknHKWe0pkBIqpNr0PnqoRxAY0nrxPkIPZD
ImAji9geZI2zpFQuJW0HPJ2ZGDBPuT4u3VTH9K7MUxPM6UutIH6h9eNAOnDheJEQp0kUmFayiSAE
5vBwxGRsnCMVb7pWm69YrIOc7qFMzffhynKb/ow7+6y42EtcnSyV7o/cjkl4Yd/L/h4PNQ1h7o9x
V2DO8Xhp2/C5hK5KVNa0xCAhBdQC+CbkkDD438tEqCHN/K58PEA3wRN9E+RLTQJcY3PqstGIu2Si
BcfhkJ3GQEQxC6K2d0AGNj3UxDPgVK1eo+uUgo16dMiLvzmIRyF3Ga3jGs5vBlUiQiS03kiMjHck
TExrMZaVxhL6x/wn3vRHMPBy/ucbiaei/TcFdOLjhbCZGmrOBQOkfCDmaS20qTebuyD1+/ati3Fv
RyxXik/FotFkWGScfzBWFeE/zPOqX2yid0zYgtmvbyG6Dk3+OEPJLKPGPFPiQvYemOZiMoietwgc
CT+nQTrlEUtiSXJKgq9FiGur8cMclwB+1ODiX5mlldRoBnigsRJof6uznmxaiPIGdQfHfjEPpBJl
6odPGlPrnOXOT4TCw+WBTQ04+S5w3FErBoMG5Hb20YC8+ms4vV1QFrcYHcPP01+MC3pW+DvKof8y
aaK8YD9Js4maYGL5CU3XBdrCcpc3pLHtNh2vBW1maKKR9Fdg0qyJo90TpTjP0mROZ8T46n9TSgpv
aWQPDaLNycdKuuAOv792zcAzSQpQX35pFQEm6Wgn21j8BIfWVaj0ZkP/9o2RGB1N7Izk69JGByWO
VyvgOi7GkK4VP72hGlT08uupVnG8jgDVSpqjfhELI3FZg8hsCvSehCBjaNpDys3g9AUemu7Sh8QV
dkc0kkIktGjl1202oI029rZMOeWMhv/M1MEEjJSBZc+Y8czbsJNzuw8WY/BD9ftz/L6H25LuVlpX
UJPk1EwKArXTO0WQw10eseEtLfcUIX6Dwx1CJGKqomvQAiB86FTn189IaLmXNIUOekwt8S8HDO3A
OVyRjP7UxTJDSuJyxyu21bf5CqryTuM4fW+v9a8Da17uHOwhGSqKnR/LBfYosejeZdgnJe6sGtUK
kc/+Ey1F7GmLEQNyXnj1K/5fh+BUeD8AyOUuwDPgrqy9jwrS2+0rqKkkdevq/47WODzrwh4uH4RK
dWcWmiLe1LvB9Ctr/ii7Saft75qnGnY3tZ76EjAyqzdnMnS0LTfUKMEwdvHgC8CBk3dXqMr53qYI
9bbvA9N3fzL/QDglBWMDflre5yrW32n8gBUZJnkWIiCmHatBqLM7hju3MHqkLMDKACZ1Q8zdrJ/+
Hj6/MxgtxivKLmlx8blxjzMNmSjC6q5jpChrzumpbvZAjPlKAAHwvE6RbIEDfuXNpIWbEIQRgmjq
B4uf/UVQedNHcaSfKNDVO7oguzX239LPgVBNOhBtdmZ/O5DSE0PWonl3Qr2xL6nLGSZWw23YS0ps
C0Up3RRJU3ppzXr1thKe0qq6aV09KGQLWpzztnYHS5u7PnwgaW/u92vv5P6tdvAMx6DVdXtiMtGh
A9ZzOsWbct86iQClp8cEqamr2WL56XatfOBL82Wy7dQI51Z4SkMNHutsxBCBUW6tQf36p4C5zqG3
F28ZO0sdNicRUBmXpnedCJFCsGpwCytKKw2l5J2KhQdAT6rr9eP+VI+vgYXun1KevldmdCdZd/fA
zeMadGt8vfqF2aNIT/GDsD2NOikSflbGgtM8h5xk97z6hMtvUGJSH5ce2t6pVJsQE6guhv5i+KmF
qmO60SPc5s48LYDBbnIXF3noeTN2R+PVbohCH1GQOeVdWuasgLjHGO2FNI1ZZNA7lzDOrrgWe/a4
UeSfVDC9lpJJvsDjtb24FqgNXCkY5p9Ixvg6j6HgV4AFdLtEO93F/34GTLZLrcnBnIkyYqTgyazG
r9mTzDEBStHXaH5SlsUTQidgxzgBwa2QSXKHRRZCnb0oywi9CVitqhHxyFY/LXe6kCW4qbn8bbba
TItJfo1kI3XImNIOVpK5tntZwvOcQCz9JxgOgEH3WGjxo7fNSChsVPhKj1D/s/8dUEMOfKVOdRN4
aPAMCH0A5nkMN+3RgKTwV8V/gmCvErItiFHP67woOcUkth98kIadyqG4PKBFEBDfsAKqnhqjGyUi
ALHCHDPgaEQfB77aOZLROuAQwBl09uKtMKn2JtQBTiwh3hZUYGKuBe9djj/ARUexFLNTFaW76Wso
16d8tEkovLNES6S/j77N+RQxe+gyZno6z0P46UMH4HffH8lwfp7LETS1D3Hfp9z704InGVIDpZI8
atL2IQulW4jhSvtgz5KxZgLpFnNce7JXCyWoPzWWaN5Nl7A6OnBRXzTi8G12PHT07TL89l3fEM7T
D3TcAe6JDwz9H/CiQtSkyjRUcC4/t6/S06OuMXxLzFMweX7jbbPZD4rYqRgMdWnnYxkvX3LobGq7
reh5n0HDiLS4u4Vd4GNE4LF0V+tfzi3BwhYUH6nls9t3RiWsN4/WKM6OlrejGbYbpgGZs+xvBpGQ
RCf0pzxqjXK3QTs7q242QkFHVevMixxa1q5JiK43csgErJLN9fyrREAVg1oN+v/Ae++eKjLQJPNQ
81bR3zjmGnhOcnlFCLNJb8y7JHYm6wpd7pRnWKKq8sC/SyZKncd1yKGas+MP6++YsLquxfvfWCP8
QW0Tw3G4XA0dD0MfrSuY4LKQ/IcbMlF04KssabQ03ZEHXxf4tOksnPkPqKlBP7wSIKvw7qnqORS3
7u0kto8/xb/lmTs+l7Y0HPdIk9q3N7X67+a0YR6IY7W7TRyBwtpSp1LOxvJ7atj/vbnAigczM7L6
3UT8mpUSspfk3M6IJaBIAB8wF7FgATSaBHCzOt4Su9vQLJwYhQydHXbIa+xo69Fabcm+fwG21Ix8
AbouUO+Nc3SJhLg4S9qkNLjhJPpOnMb0BKYjapzvLLyn9Fo3ZEMb8plHZBNlG5DdiNUKhoC/N17f
2nae+/e5d2lySgJbtNzATcv3bRz90IGFU4z5sjaHg1nfdaUUeoSiL0hu9O8Lw36c7E6BnZcJI0Ey
Rl9HsplAmc2VXT4FBbcgyiKq+lgMTTgXfaJZzaq+vGMlSKYZHLE0427VGdDl27vPJDGHMUvq5801
+9vaU/joC1MyoMdukngIzTHPnqAmzh6RfURKwMeLFs8t0dmewpRQ8hdLuc/Vv6zmnwJn0h/gvjJ/
IAuRhN76y2yMZZc4ISGWRsK9j+yETgR2fAsajEeWuVyJHmLNHm5/HOKhOyxXSTqebN8GsWEcLpE1
IOxH7DH/stxm/hLCGiqA89Xvbs/BYwvSbLB/4BbmkxZ7CmSJoqq0j3UmRURUgvAtsXDlFKbECft5
XKFJU23lmEUHpeqZ47W4Xh15DTYbDNYtRCLIG8SdM6hB3ft1irvEkvSonKOu1+Tfb2HMP5ZY+Trw
7kDDVpN5JV3Qd9nDR0NsTOCYZ6utPEe0dI0IxmeWzUVl+Na+7pE5+e0CtFlAi/bk4MaUdIg1mKxG
uV0CafHMdHJf8hpi8A2RrSRj71psfN9D36kK3u1Lmd+uVH8U79hJtt5WgZDNeezqOKFrvrAHaJAw
AA3pWQaAWWgn7rkjbPS8kyO4ZZRY5eHgD3xom3m+9kMq4ucwJnpWIC2ZekCQJOCV8YQSzqSapkIM
tKSkPm1DtnE5rHo5rLBgIiqnTKElMRYzWrk49VPd8i7jmru7WHWtA0rJFZcEXMZ1B+4X8gD9xeG7
wW2kVQgEyd5d1xYW5n44+HJjP8BaFpIqYVzBcmj9hvlVlgKeRDJN683J0yTzpiwPEgUrJT+1jB4s
FAuoGTMpO6RPQ/nOz//LtU2UdSvVmsOxsDhcwL/S1YHM2YatWkHnYq2FjANo1egKzdDM3I11HMPJ
6MA2yEDXlUosxZc/atJOPprQmAMOYkme9QcNqdH9RsAu+tul2r2o2yvdgMY8ChYQnJUimsh6FL/R
DeL5IrjMvKEVNuAFhN6zAeHKkIXcc1TaXT2u00KXsWeb/Mx7SGPexFErNO286gQcUalK7TehyAIp
IOaT9uNlTZNfMOk06dZLIYJCV8RN2jGHdpGyQqGBEhLnPVJejBpohpKQeq6ZbTqFf7RHyRaopD+1
bfz/MLvAsJxh/n+IWt9q+/d3Ot8lWGqfRU9HaOhvha89G1+pf56VKaO/XPWQEwgm9Llnne8j8a4M
RTanfKU+VAItO/MdbitMyc89I36nOP3nzkBMLcKjwV4Hhr/ejWgEc95AajO2A11/cirFV9fnUE6C
shJaI/ia42Vo7+Kn4Bi1wIkVwjzRjd8SHGac6W/3Xr9Xzq36Uof7VZJIv5PE3+OoNANk72UVgXnE
Og6aJvYcb2Dh6aB9K3+3JJjDDMOcK4I20VSiA+tz3GYctlhZd3YQsD3Eg7NJkNWLN3dAaEmHcnzg
eE5B+Pq/qEuBNoiBDRX0OAYOTDUijME2EpNzRkDeWsTrdRtIwB55+fvNmMsZafxRP33i1Gfh2Qeu
pXfbEK4w8Fz8s7GIwX2urtiiQN1HKP+CsZxGasbEAQ+zA2RR5yhCNL5AVTdC79Niien5qF3widkN
zYFiwZeeR9XpxqOJR0xM5So5fPVNO8Y9fUujyfUBPdlZmzqTSz9NeLtFOww6P/qrUbIiK23CSrkI
/6b11lGWNVfYl1MR0zTynZQTvO9amh2XX59yH8u7DDqDGl22YXgWazp0l6tNfxgPJLCa7oHt36en
wnFFvoKCVVXgD7R5d3sf1uAZouCj/6HUhIT1c8RIkyau/d6+fSirdQYY4ohcFjs1QLErzpEZVNt/
HtLEWe9d/z5V+/sPXu9cz2FgHy7lMTpzJ2lumOaaOwlRg/60rZEJ/0rncqtEUBJUR/6izHMN0clL
tPzOj0pWtCh8PWi0eSXjFj4hhzGo4MwbR3NkblXz+yNioCX1KiCvdhI01rIqvDJ1S+ctNwDvEtPW
++zPzHmo0iN+Y24cosy92+GQCY7zeqfiinPDJkffdJaDUh5u/F/hnhQPgRLkC8ujor6eGmy7aCSr
i4zptun7CESOHlMtzUICKzFL2DGKwrpQ0ozLf5L5Mr2camUtrfjN2f9TSLXHhvKtb52f+Z55nzyk
NgSicR7C+ej2NjZHE1XPrVtffoy/sZQQeqwOmfcMo3Mwpl0EbLREkO60CRnUA70Bu6AESo5VBrG8
ihr5XwQE9KmKzXouVw66YfyKlzmId9J7NiVlAhcXAe/JBM5Smox1hqhCwzlsh1WbO+C5TFy6mzUV
HVIHSvUHSvPwTNRY6dOYuzZRKNKXpLod3IJ9JtP/Z8dGb5sF9mW2PDB77YGL1nr14y7ZEMPMcXJi
Oq9XO23N1gBXV4IroQ+chFP5UOnbwscueToW0ke95t5bKNBNkxUtQUcJMqYpojiiJulDZ7y9AQHg
f5ZUYoKVY4m3etKR9nO6E/GnvWkvrqJZeGNv5tTp6n2VLR9w7QeLk7m/OkmTwcq4urzUhdsInRwA
RJKCPWcBOIngSf8CkdhJFNnDyxVMCqUr6Zm+55c8ULTHd0/Dmi1dsmKAyinoicwcz6d/wnKHTKQp
r+C6wxo5BLL5xB5BeqOBGkFPxjGcbWxcqo0CZ3GA+BBA3mb7VdL0OpvLglz9x/e+oC13tC3NwvYt
ceeFsHNvjAAN935tF3p/IW5kAdnqhNRsRvWhj4agA9o6dtrmpV9LUOk2QuRW8TpQef2pAfG8bzTo
jsKwLpeOjJtMRKjTgD4+4iaGI6WZuxqpzULDv1/FjTG25Rc5A9v3vvgkFP59doaUxgYq8XGgK8YE
EBmo+SVaZ/jWaMpmHIefiyEGg+iFYRfobXaJ7S2Lkrc62kWBp/3iB2EJZrn7EyO1dIsEC9Xp+j/7
MaFkcRsDIoBf/aRChRZeCFjmxvpjfMPty2zAKNHb+nrtfAfAguJUP9dHz5XvxPDCW+9a+lSa4yO/
8I6xNdwdtH0xiczKnQdXRf5b+8Dz5oYyrPvR0sl59/NqEpDgoshls2HPm8stAbGR8kKSG3o2dwOH
9yS7/kp4SBduWU+kdsedbByCfLhi5eF02EHRFpspneEtyYMDydykSVRqKW97LatJRjaedx99iUTU
MIOBj7DM4IXspnjrGApEf+JS/Ur9eE0bU8PgyduXaW8Jk7FE15v1A7dYBpgYlAgt3dNXWik3FMfj
7QYkvRlfB27r85tYpO+wbC0Td58B15pxbr5uw1TdCYAnIzgAfGi8T58sPdi+FjjGYH/B4UFdyOAQ
qBgwohL/FaBlpseZ3BgwbppN5EzLikho4XCveRQrxS/801J2OMHx+TAhmk3555V2BeyxGXWwWVPP
qwYfhbh1hVHTOtq0SHvbeKJE+axH37G3/4OvOUJBy4WGf7NdJNzq6vuwxGPaYyJwDwyaq/IJu//W
zXNdKyzs3/Y1WHY3QwmKGMpf3EYs6M7wptCUz6Pv/bP5Wv1NaXe1U34ExtKqtM05/170DqS1AcBO
i8HiS4ZbUdlQKzhYGGbeOhf7QOFBMQMcwsBgN6ST8QNyXhuQ/XR2/7lWAe2Z15uT1pQuXHA7u2Rf
Om84pkyIOgK/wQ74aOYT1I4oszk3A3JcfZ2xSMZFI1jMe5KaXwR841/uELknlTMBpyw7eqKfd8hZ
AqY09Pqgo0GDhn1RHtCwTNHKldZCueP7XjH9Od63LWYhTBY9KvF4UYrJBZkmBA1cOvxfMN9A9LhY
P2ireyVC7+W6v47q0vyYRrdRwrcOeR4Iak4urZEmvcqxh9WU6jBWUiNMZP2H6wI4VF8Cv7LkU/qS
9uyJHzgQaFLLtecdRR6JTkUtkvR2mDFLVmCTHj7mbUPGb1zxSE0EgKW5at/B43Lj1H0BPy+n4tH7
yR6AEw+F1kHB7d4ds1PmmBvqNa8VsXqgiSsLTpyTWpPXDeXaNKaLCrIVBHWSiTsPtXyYaHgz+XQF
YqXAuDnl1bMF4qLHamIsCcKjQ+bCe/Nh3I3HfaM5KRY+NAyXfKgisIuQ9rkcnhi6DVjeNSpVhSDC
00+0rt0nyLSKGjp3qEyqvL2Yjl12IQGHfJ1Zi7L3i4FiU07M3ig4U8r1s/zUDSBDeHIl1/g5jpw9
Ww5aibBAT02PAxJe0taTSsxP/0Mt844bURsvNZL+TNNbuy1WJrf60wt3+gFEsErps5MMGyH74LW5
H79K4DCm3vg7QyhNxsP/EFdmL/CzCSkO+yxLw4SwyreQMl/m9raCQ7l+d+HhfbVOz7Oy/oHlXn4D
TiYFGKOmbTZw99Y+zY2mCqj4gvlTXgutO+hWZ3J7hh/9BqeBQsuZApQcvWt9IU7Qw05d9vQUeApo
ai2vBbYTEik5GnVNyuOlHd/NNsNmu+nL9uAzbJedHJaMFNv2m8fvege73jS+1DnUA56/AqcJkaw6
qSOMbylIqmAdffX9VrTNbdWoTkacMAEVoUs5ydCRC8nd58Ud/n1YmJ+J3Qe8MkZ+SA+vDEfqsh/2
nvBXEjIUkR56bmxF8k+hB/o3iEA8xvk7oYeWpinGWhe0AYL6cI8pKoj+sFo47KKLLt0Ct1PFD2ks
Ml5Hn6ElXUE9KzqDWU2Gj6jh5EGuZiuW0gLQH3e/YedWAzZfy3Lg5wVkjMa1dx69z82sYWp8CqQZ
+jwWi4nX1fK0oYzsFjqB+PRfYgj4Y+wIiJEgP0ANTlDvrVk/BJ4vqY5Lm+4IPllEA9/zQfEpWRPZ
E0gWKEtySlo9qPuIXFotuyTb2stNWfR9IBFclPviPLABUTB/B5lKXujsLofYhgfJNiCKcf2AfXkN
e1BnSF4TwciF/kC4BkM5cGSmpM0WyGSlMpfUURW2Z/Tmm7+nfvgqUJVqMqYZmqpYXgCpd2zwtsEa
/9XlWUm8Cv92XbKcLmgwPIWL7/DzyNZyEZ7ibFfHwZYXauQAjm0Eh5D5B/cnoqJugEnL+rKu448k
X8lpMliMmRxfGEYhRRcGfU2Xm8t6wMFPa+/uBAUk3cLjZkzfgl5ME5SinWTNClBWRm4rCCcGTY+9
nE2LjtbKjvcXesyCS9eWbna/deoHXtb3DBWd7zebCeeNIVdh/4JDO3eqMNGzm3POV6zoAs5mYKLI
zzhEEpUmUdvQODWYd6KgPBuQhX27bQEFYcC2uCi5LfmF2mJ/VfmsRdKnDc9YapZq4mLU/BzxpzG3
DNSsivcFKIVqEKKOhjMGU+vCNlf8ejGwS88SY2AmMLGO7lvqyzur0smy25G/vkk6PAUn+Rd9k/Un
3Fqurf+XNn7pnGP/GzLbbUyznWBme4M59gdWZfPwZKVTC0qdC63dlSUjsVPLE+nHqH5jz5iPYb6U
IvkDU8KGLtr3nAErXKCUY5jg/bobnFFumugWTsuY3HYKKxqM8xfWsG0lzJOFn4rEjXQvt7Yw5nyK
uQl1Inw4KTmV2Kehdtg7hRX05aKA8aSa53u/g8OAeN0PVrDh9H2ZAuwWyjHNjTYEsei3o16ZpiyV
Num8F1oU65BN/rUmqiEjDJFNuYj7kKkMeNuBv264sCb06NZVDHSiPjseeK2pvfQLoriggu0YywOf
xjIzI7uiqu2saBiSQfV6UrJq7ZWQjdLPlTbSY0An/l19EZdlj9MIgOJqZjOfNjqugNRb3ZsItKB6
KHS0kuDga4os3Og43rKTCPXBAPF3ac2EocniikMkytsEtijZ1OnLVQSuth73DkRXK9T7ztGafmGA
J8Gh4fFPNKHd4g0DkcAApVdVNssef9XKLw1zDBzQ6235nNYCTP3q32L+A7aH7yb1g649WbFK4HW1
sDTHb4qg8cSDiPOztZrca4qHqp0+xsqfb3kR/6sC1DE8znmFmXlKPEhV+yofLBRMHuy0OUS97b91
6Fi3iZ7QjJCqa3G1/d8rRhhpDaUmlR6llW1p7dD9mnRAD8/Cfo1rsh8CLMEozk8RgXIQGJq4ZTkr
hllAYJERXDXThqIT6rHc0lG7xMZ1bWTVOCDZ0fuO81Qv0Mp+NTNnhtDDwWjecP6tsEETWt9JmohS
2je6kxr2Hby6SVYiy7Kt58k5PgGfaerW3KUxt8kkzqbboC1HIxofVD/rOkLWB4Eot2aCtrkFxCSj
lxjUcAi3C5qOQ4ynbDAWPQ+LdTMqg4W4nLNBK7fWwIANqCOLRA362Th74z3McMIFpSqx7EpmNTLC
Gw7OYf7K/nkHW9hkOFVcnUidnJN8jI4ZWbVsvY+4+a2tdRF8arYdSn7AG0H7Vk5TLh7J/zrO1mnS
fxKDrj90nam+lzk9g97rkoKivhvQfky0zkCjM6ubONIS5UM5JuQLQSKxtIaU3UyU+pyS+InOGC/o
V3VIu9k1plA5+GtAKziN0/IX+YYKkXQmYI4DnLKl4tv65mI4B48G7vAQ4XpH6CafaRdAk2MXGaYG
hXmS9DDavbDD5MIJq4CpEdP6uW23rNVBtIhV+ZJydZqhaLEG6cM0l+RPJL1u3KDCex5w8XrY5Sn9
FaZieCT857ofPAemB+Bx3ceD1RUbP7YZQtzZnI08raFIIxA3Yvf1KTVOned3UkZqq2eHfl1hmdpI
B2xBl7DFb6HKmmiEYQcPjfEFk/s9Xj1+7aFEBN4QHoO7ROR/K44R1FxzeG8FUkify04HZS/YbkRO
W8tRUPzf4Y1bQ2EEyiqmAgrL0+jLZ7c0vaR6bzNujuXzLWSaZFo9wahnXDd6OoJkKETsKFr10EJK
G7n1c0TAPfkfXKNEplEJHc1m6FsT4r8uCTaRu5nOpc6kghXcO2P7/BNphSBG8g9vnORXKMDmcu2K
wXXOQBgd0Oh6PPJ6LzBQYaYBRKSuuQgKEx0EZAnAvVMXR46XYGXjovIfWIvfRDSXXEt7kfZiuRYq
Ar0JxUzNcOyPcjTkdhOsj7C5GMhrbCR8PS1pEQcJ+SyYjaFlIf7Cc32zkcEGGMfN476cu51c6F/H
dzW7DeUUqa4eJg2VMz8kAnAMkfhHHh99DFuztiXRIcinp02WxkdiQqLDQWtIv+UZReB/VU7fq15I
X+uoNts7pYVRplOL+/mXowTGILcg2QuXQpc4Aq3OqazsVgAGubb+6gC4KKOj5dadDeVICYMcRhJx
PpSicw6txucVAHD0zdRgeEdszJ01BVwp3MJnya3mkWSTZrbo8HYyyr0oGXjjnu7Tp9VjRu5ZP6aI
xwQ1oi2G213JaT57XOcwlmvXWoNSMUjJZBrGOSdqFZIkPA6qqoxp+Wm1q5VjZuz+6+pS89ST98Uo
1vH3wV+Az4sy9YRM53n0916rVP8M9fV9n0cdWyyICJMpsjC0Xxg1cyYKNZRAfNRACz7VpVxAn2wF
GezZ2+/viA7EWjwRZd+zp4hl0uFVfJqGaAGDEMLc8Hq5Tj8UGFsGHhCc1EjeRVny4F6EYRLl23Ev
pSbo1z87IfKAfc0c59OO33tcLNTYNKlC6PDI5bcGkV47+tNhQlnbP0W8ykUDNA3XO6Z8U2gcsqB2
nXByHzM4rcX8k69T76Il4cYMHSGca8BPuk5dSaj1CL79kEtLgXA8PeHlVgR9YJfRRYSP18EZQtbs
Pelrpk/V2pwiDGPQGNdREkGb8tU7Yyv0UbKntzf7tllJMQLRmDtnzPOh5Fz5cGriRbozZpMI6R0j
6KBnnUaUdoSdJuXo+JbOuAto+jzMzDJxfC+DJXJG7tUiSEDvXUKcqiepcLlYsw3zw3DgD5XqMKg/
ZMXSv3Pirq3Jn02A4lpUcFa++kTDRwpUg+G52lp8R3+QPPTPTdfgZiJfWo7pnoqs7MEeUiWienLS
CZiHNGfN9LDxuoFLX/UB7AswFcrPaV/OzSuwkY5hM91uKkL+2H6JgPcJnpVA8d7uycZwCOKkb99+
O5wbmIAEYnuslcpC97kdr+hKBK8sD49ibEOKuCxPvg1Az9kr1kh+ZVj3OHQlEmCjSJMREfodgFCM
X3nZf0CdrILuNrElK4/j5dpTKvgnJ3BTVDbNslCDDFz5OKzFTnBOLOwz0dvtO6t24ZdTcM646Q/C
RNDpDPF1iDwujKSB5iZWOXeOw17dD7WBdqn+Kb478/SMiVwepgTdMXBDwAfWGgmazm4/pGTpcpYL
BKroijRv3U3YDmj2MstfUNapD9beheR5ch+WVOvKnBar1qZNvIa8cqyjcNNZk7bsxxNSJJBu/gT7
8LIq10wLnLgoNnBasgbn4D0rAtyIfRzGbB4h5GOisut26jjezvUnre0LlTg4FpvPHX4uCRgFJe2U
MDWveEaWkOCRnUa6fZAGZBIxQr5PVIRu+G7dUJbwKwO2EJJpwgD5NASDNA9b3N44K5p5XwahrvTl
p2LPQQG8/7NUlCmWGKGUvPZfvbPOn26q0BDQBFWK9jgGI7Pdad90uejK3eUGS57HQZ578jDnz6Tu
oo5C+cTPSixN2c/mZmefTgcAnUljMllk3SBuBRcMZkp3UWWlfWEA1GyIwe8WaIXsB6J6HMjLIWM/
zpTEESQnnV7m88vKRaIMZ636B98/qyHkCzJJYJ6xnqLieh+Edniqowzos52co1NKe/hWCtkPySb3
6L/YzsFyoyuObK5rd1J5CP4on4uYpBYRgNn4Bq8ZepYoC0AWY0JZ3AzqVVxAHFybChyXPQ73ZdJ1
Tn66kMBquNPuIduLcaVWA/7ojpBHy1PB8bYv0twQYYHL0/LZEeq0jxrXbCB+jgAIfn5uNch27da6
58TmRkbVv6XL1IlCXBpj0EJMich+0A4uFnhyupF+XKN77i42MN9g7piXCjqa7JbR/oLFnelWR8m8
Ql7+fotmYRMTi3LGPSHsUOGe66nJI0dD127r4XEWxY6nYt9+IV3uPiRbg7WF731XrV+xEZI8B0PS
Frk8D03TKk+qLiJm5FhnbOxxwMBSdOAJo+z1Je8sfiU4O7+4A8BKE1PunqXmoph4jnTnokcrE5T9
4/iiQWFuVOz16CfN4G47YPTHIU/aYs6dsdD4BgzmSm5GcbSOv3MRtoJCBs8ejNTD5fwmtGK8+d/K
lUnVeFKJVynI/ws61Z0nV4rabOEhG489ovNEum8eUcmTgcH0UYw1Tdn+VxWofNyaOvOm3GioXOl0
sB6/NDXbc9+EV406GiNqeGTx3JXXKA3crqN0Yv9ES6SLJratz2FEt+vTozU9EmhCsqFdji2L69Kx
Vh5ZO/M+hA/dBsSfIQuEkikw4sjdeM7KAoJmAvUO4BWKBKJLENMBFHFAluqukeQSw7+Q3CxI+eia
gYjJbLFLIq90WQpa+Lgu4S/VReNbTHvqtoSg3vMzs2GBm4RIE0JPWuubH+RRU+fTbdFjOl4c6pba
tebYtNF2B+IwsmZUywre/j2q45SgwkfBxULG1oJfu3URdqxXZsaB8hSD5t/tOjr7Jm48+rFEIp8v
16921e34X5+KscN8C8iSgZo0Tvak+2+RK4wsC7naLH99OT2R9rDVAexg/D/NuZ0/u0Wq8Gxo6/05
vVLAhDJGtmZqcWYzzyl4Nxb5/jA1jrgZAddgQq1gTQA1WaJjJAPUnXOYqSgjDV4x1/Zj4ygKMawQ
yxMi0H58z+6U1oxV5vDZtVIC9jEECn3uUdB49XFWFni8/BIJr6MP7u0dW422x9r3Df0b8hAc5HRW
cecUBL0OX0hWNT9hMxl3OD492W32snAd4p/CFRqSsS1kbppuTwSwX2NA17bdEHdsHq9xzTff96Dg
vfW43xP6xQdneFKcPTIRC3z/ZYp9Mvc0BDobpbFXWSR1q4jn+CLOUkp1HtTLJkFLMoLK2CM59S9x
0uJIaRNWSKl36r+66i5c7CaJHG2yazbhBqOyK8TTlIaOSnF6sLtY2/SeD6a6b4G0Gdou37EnzIdQ
R7KEq9Ybxpd4k95qg7zJZ/TURwhMByTlI4f67aqmXZ4bQbRLMhGBGBYKQo0xutI5OKZuSDRXUJ5n
+zPdstmDPGrFKYeX9+w7RItf+O/8q9TSaIO1Yb/CTm4Z5fk4QrcfqfBP22d6A8WwhJymxnqZqZCo
KOTaOzeaYM1tcfN48+MKjOxPdb2jTbCA3PR2TLGCVsnW5CqopWEAgHl80TsPRLNjk9/Cx/LAJh6j
I2E/D0wT/X+QF2Fr7vaeiHHVuXvSDBXlEXOsyny/AJ81t0K66oOqbyjv7RV3qkEoJH1+yQ8MKdcx
1srweAzFhhwipF4DNy+Wf24J8C0HSOx4kQ1IUUifIuyZV5CO1qN8S1y5Bh2wkET7iqxrny9CtDnZ
/2HPQi+1qU3vNzDYrkXDWT55rtqUKJ0hejdfp8Ct/Xh+o1aqBgaXfbfZFxHzvpgnykCK82F8X7qp
mDPm08CFu6U8iegRuF7TQlJwjpFsL+B3SSP36iHlMB0laO17Lbk0x+++cRbB0Qw/F8Hi8/SmhWvS
YCcNEXxnPc0N0tgEPSOYfSK/axVM/6XCHzx7UKL3aqLnNAbtAQ5LFPOlfpmmAPlGY21yAHK7Nx+H
ccUy/7ZeR4n5sTyVLTSjPRd1c1373RHSH4HNs+H51DlGKcPvgWIl5xJRAb8tDti0EO0Spvo8ONed
MWMQrxBmcM7qCn3cTbWzVle0vB4+lwXPsVeTwjQRUfo5bBpP2mE3QSI5hmbo9I1GvaFr5sEkO+9q
hlwkHqWK/NhwdFIpfPXtPVJeFM5aAbn9HKqeIeiK27R7T/sRqtMP4w+JcDQLJ+PK4nxm+wdIbMWc
9F1FAzWa7qAEGW/I+V8710CKlQRX8UIZN+csyKCQKrzbsSjy0B6+Ellpm3QNEmrCsQj73rCxrZkU
Irr2ctD/tT9fc3kh90M2dC5oQu89awtJ6e0pH75flbZXbPkrd+h2sh7PykiolkmUhbsF/BM33eCr
IMo339EZzFDxFuh8VqmyWHNYhg9g7O1j1jDYD9sGE4eBOy6DsVq3/0uK/tQGwggRrPLfzZ8szMr0
nf7Vo+uv6AtGfz1zKU5kn+iNNrjocDariszgz1J++D/YsUIYLLntQSTrJX4K4sZBHXp2xE8LUdEL
+pTZoe3c21i84Evarsp/vXasUhcvQgpukfnoNciHO/RJhoPU+vAZWTIPbAarjk7g6PRxrsbCu5tz
LhRsYwYkTu+VvzmU3sOLOkDlhES2xLzKfQt4MjErmR0Galh19rO/23l4Ai5jz/8EZjnjgOKftE/7
UQ3FtDAtZKBSeWMY7mkPsVfzgBPski+VHZXxX6RMO2T0sxsFBfCoZx0Uh+HRr/Q9K6Jdy9Ww0mDb
KE9yHMQHYCRGRJMga5DuR6avseVQJfpPaRZzQ3ujWJTNngRVWe9gkH2VrczHhdd+mVerSgd8jOsT
GBZjnzJm68nXoSPzTOLsqnh0yzXTBiH07J6WVmk+E1Xl/gtuY+w8HhG9tLT8Al1WcsuhVFS1vF2H
Rj68G9GPk+j3p6qjEIl2MrgUedIuCn0HyOGC/6PrsZ7d8/MzkJAU/c8OXhqgmuz9b9UshXjzCRDt
9BXYUpdZMJpAZT6qr5t3MIdrMEewOUFD2M2TsU28yKgahgcS3WQJ2W8ytvENOrvvh6HEZaMC3Ytm
Oxa6iQNMuvatuU4/eiN7vGpdpW5M9bjU5watWEcmlYcKiq2ZpwZytr7P3ilEEuHvdJBInrUhOkwX
JhzoRzlOSrhXDj9XJjKJnPIsNYfMPL/JI9PDvso1ykJtrqC5+t9QW/uY6POCpyiHrTDbNCnECQqD
4x2IiJucPMkjpXb+fw5yAUz+FWYj1qIC0HI4sEYB724cPA/HT1BJ7AEvOpojcCrNhiLDozd003ph
r3XAkMauvay2+W9XEXw2Pixi4u8LzW2Cj4yNrfdejAuqKEVYAeNtFUk9eBwumEfjFFgbewFdTA0G
+S/teinWK4/sjdjm/zxfPYH646UMvMihpJ32eiXJTmoIO2n4rK/wpvReoZXUSbe7sTvFJacPHX8J
PvS2x80zOPKPVYe4a3yzC4u8pHX72la9FVN8pmbrN+5qJdc2V6XhIvRwgF7QUBEZSn5jxFy8L30Y
YmdcX9emV/g9GDfWCcqE8kz2x8PNa/5GFpYOoSAhbz2wtQHsi9DVl0cosfhHGUJHFP96VD/r17ps
6VFeW7WDxckgFhoLCjdiLIPXd+YOzsTaP15jRlzD8jPRrAVdU44PHztAHfJQP9fECphcPCHgQ+BV
bkTHBnY3aQcPhUOyfQnv/lwV4nc/KfAjIncx0fuq+4lbF+fK87qomAzWSX4tJXS2JBV1wlk/T2pr
qmuqnfPESqNgjYlt02w8YluPdlYohPxbFFlOBqqVWV9O9Qz5ODtF0BZFNL7mu6Kkeoa2uPFdyzJ/
AUR32pD6kJ0LhW2uXODb3SLXaqI5VfYoeiCbOtBeYAvI6GvxfrjvUo4dUMxzGz/m52H2NtCWFVfM
i78UXENRnwhTedQ/128EZ2zEx47sG2kvWVH0ITddifhu3+sL6yIV3slcAMrOTsshIAqx/ttpzVT/
kkNrOSRCIecrPvDVR11Ua4A0yhs17jQX/IZeePNRcCVXjDMGUav598az4BmWWNRx67K3D7t/nqT+
RjbS1+4SGtxE7ufK/7eBa0wLZdCiRZbRY4eU+qIvWMdaMeWMlLew2E1rTi0ymea6bI3D1L8TmBqy
Cg41OtCXE9h5IpZ/CgEF5v7BljeDjCn/BAiIHhOp9C43FZqCyZczi58Zzr0zDPH4uXtUeMWkYKAn
qmT9GjlWKPrbgqTOCGmzlzJ9DYSLygH1ujQMiKnfTRvHK3CLCU05F1EtyaIzl2ChAQGoLiYuonBH
AL/j2fwg75ZMAylKGpnDMU4XEtbHQ3vq12MTCy/mCocwqVuUZpKf+aYK7Pemu8JN00Tp4S6172Lg
YQ1tzfM3UmbFxFID1x7/oXBiQyZSdKuT6xmP39YAZ99cIr1j0rQafqltA8+AXlHYtsuOvSC17YD9
7M5zSLooPemyPdbrC+EOQpt3vP5gLnp4C2+UsVUwtrRRVGdSZRx0TA5qoeIfs1lEjOEJENjsJe4P
+Q7bR3x5FFqh09VFhmVYiHvBFg1VLBhX8FJeIuR7a95eX5HwPAHn+poscnFmMXTu4O8kWmTNLzM9
MENtjCXgElBdxMwilhA9XwW0kbk7BbRo6ZeGgRCDewmkn/1ej6f57hZ4Ns1Y8S0vmYAukcYvGX6k
Q6iSruAEKhvDVRudsDH9t/JjQXi8+W5MGkf3ovb+Vjgvg0BRj7ptB3rb3wL82vCY6mcEBnndIuLS
gejWHTwgf7bqZ4kK681RF1e/7f4KyZuNMo09rS6xdkdnG1bSVnQmG4D+Gyv401EgWnHRR5gkzBeQ
rbyAWH5jv01gqdXEHFONYOuxCARihcKYC1hY+dtAxVbGGByBdxwBu7vJIw9NhjmqM7l9V6FIYvtV
BF//EYzjAw6Y/XGQyT3S2IJY/KJdDL6/mcowTi7pW0MFtAGHQsS0G4ilPxK0KCOrqepPCdvWjRgL
FJQ5C13Lp5LMlFADt0oF2duZtBINKsNbzQs8BRGFSXCdzA/3jSt/M8qlxizb2gTDsVU7h9LecAWQ
rP10tX6mtu5Xs0PqGhldZdDOVn8dalv0M5uizmnKLb/uzBQn0fNkTfZWtEq9NSxzjsMAJqMx2Zls
a0fLMOv4vHTg8q0OscyQwOjRNVUe8buNmZJLLaRfDpxaZg8PlU2l3wyZ+gh6stk11VwnlfxAkheh
yVs8AYZMFdhPs88Wgk1E7KGvBmDJCnqdrzofSFpYatNZBOaIdd9F7c8TW+HZC9vC+01cLG1a/SJH
0hltM7TOmT4y4mzXx58s2y80w9Y8ZNva8Wi5duWTxjhcdc5OWHoneDlX42qz0KmyZFSTizGer3ib
/ZrGiBI7xv469usdhm/YUQDPYF0qDAlYDi/0+rmsciJbbTIszQIhhrAPP17CNoWpb4WPb/h1A3Io
kHAw7NeD2PHkhXmZ1vkoGAjaHMvBki4XX6e0KAdtRtDnUI94mSvAWJTW/c95CdO386SYOMc4aKZx
bdUp5WY654gi0Is6AZlazxXBVM8TsiDLXsBOvC68W8qtMxMGqH51tiMdSWOJV55F+9GZGMbsGd+F
0ZPsNSYCvtbNTTBdetKWuFhyDz8gsk1I02N/QRna/zj5/BD+rMDpS24q8hkUiVoZ0fsM2lhmya+r
vQuWSbzwb5gJ6Fv2/fzE/UhofcW7ki4YTJn2LMxf1dZBoKkDoAvxha+Ew62BPmuLNZ5S/86Y0B2R
cTVTCYH4/Uh65nss5+0gx9NLMNgKnNsWssFhUZsLuKWCAIryEJQcwpZDlpplgiS226bHJLTWyBNR
k8gNB27VwoLVzASHupmg+e16ujQF9EQzGBFFcQ8bCYQ6/4IoMvOAhUkczsq7Fpxo/ZCmETXq71eL
iwBSUJaX/Bthavfaa9y64wOk20Na7A5aLmVH9WD6bLJz3qaWydrx7kvOedJeIq5n0Fc9KR1iMsIc
//Kc+9IS13C4a+aBn8bWCD9tPuHh/qoOHLHnLMuAsI4SLRoLiOJ6KAB3tmj/tLWFrPS30XEFOdtf
YSrtp5hkhUK2a5mHPgGpZ42sFlOuzx93MpLXWNa3MFTgLSeyjfN3CL7zR3paFBcQfvALa6BDheB5
jTuFD9zQf+UFrMxIHQTRIsUYjU+MZdGZqisNp6aUSsliqnrRmHGdIeZ5wKYuh24FuPojI3NKP8IT
fhycy7SHORMNgcvEqoc5PZ/F/4hejncM8qPYN2NKnK1KLV/IOpbLQhI7bL7S4xwbLXRh/jQwAafi
vU/qlFU1mKrW22NooYCzgAkI5nsFUR6osLJFLKVBWJZYefxJfEqhM62rKEvsqOMktz158KJ6e2u1
Z09mMQa+aIiiKEWH7KWhmnmLFLv4O9xA8SRz+MBNe+J3TABq+cCCw13H4Fq46HV6nrel07t4r3z0
PWVLe5itC768aD6+h6UoFNpf3wyZUZ4WPbtGHJuK+1TsusHjbogtsMD7eIE3Ytli/TLvKBZlpEEY
QNUsGpYYU1MNVpGsogGMlLKIgY+cbAfKYab621yEgUGXqRZqktHmhf0cKWLzR6aGaKXuJLFwDpzd
7DviHnUj0KkkUO8AdRaza7ke0XwAqCFVDUxfwpqPK8gkpfguD6ClXzzX+VtNqnYPvyP4Ebg9uneF
H9UTUJnfQpWgauWXUk+U7R1c1n45S/qFmgTlDS+ThFIvN548CMTDoVjVfZqvTTJp8vgXkXvRi28s
Fc5Kw8ArXkZ6lyLjVyIU5o5KDI3JJcp0QCX2JsjWk3sjTezrZRSrRwOz5ldT2oLeqoIv8NYJR4db
Vw4dbYUUAYvTvPNZJ/3stUuOVbfPTOIx0LP7NxcAOqT3awFxdzd7gpcNsj2hmgDc5OrprPmILWn5
ul3hN3qYE/5LD9tT0XaT9PeTfI3RMDqMYutr3fSiIEaNsPwZ97Snowx5QPx+9A5MfstFD2Euw1AC
y6rfO3gAckgfjCNyNV9GwIoB0M9/S5vSCjqO0R9mZgCfEphqMjqcshDzbt8djm7onXJlJnhcMYSO
QXtPIzyG3/k+r44C6Pd+eUDvomRcvjNAJ8egxB2W4FKk2LTbgULKAgiiz+qOgeXon02WpTpoELHF
7klr7t+r566v/BPAQ4cODdx+2oaUwnhNbnfxq+EHio+/0/6FKB2ZGkniEmk08UwimQMArogA0Pts
k/5Ufuxoqm9ymFVl+Yrgrb33uwSy1GmRghia2iHB+Oi0pq6GuotGAteWdWL0jQTlR+VcTtKBK8r1
H7lz4b5qYwoxDNP7yqX1oHh5/O1HOyDHB548YJQ4WofL1au7iuFhjw9Obs6i/92REakG6XGKA4JG
Izha+Lbu/zxr+cW2sh3w7VDEmjEoiYqvaKLMpm86X9EkP5eB+aGOBYNWxw1BDlawmoVD3qjbuviK
7dg5hpKLIDo/7BuWRALSAg9UEE7JQq90AfIdI1MpU1VVtfNkIzXiYpi9fRjETK4GmBeO9GdzgRfA
/Wimjqgt5oCKKveVojGKMwEwYuZP31OPqAXSBiHzcHgJxUZuGX02QAoFlEZmA+nV3waJ3Oo+rBWg
pkNCIwZq282mCoXfmEePFRpxYNzbMesuZhXlyfKmDeJ8kBYqrzEX/3+LK9Ml1Ti3cpTTeobWT/8G
AkaJzVhIr+qo2PB96oKtioqgiI61z/Fu8JKXNgpYOLpREMFDvtRFXac2dbcimmXYV4x50ZT+sWa8
Szxj7hNjYCip5JDIx5KXB4xt66KMKHe7tex4l3EiaIlt+OIhIpI5aQickhwqExlM4Y0UTX0CjE78
cY4OlnjtLBvrsyAtQg2lReZd+fVEZfyXPo9vlY2NOEyse80jpQsX+0xvOP/Uw4gIcy2rT5ql9Jvi
/lgE8ggQ6UUDEMAa7TZdRDRQtsgLQYeAK4EZkQD/ALEavcDM80S7i4F2X//1IC6EbCnoD1GSwJF3
FTvfLTumr8SDXrqgcBrRKyPXILNyYuPtns/beZX70CYjwykEv4JfrWc12EUA5tek9u29ugFOCKKO
opDncqKFtZFzw8HD7MGJB+pzIowcMDApvEmpXu6RI+dd48Yt/RpaN3pbWvD+UaAxxIDnsb59/Wb4
4lHGk2dobyq8S1XASGXGeUfdlVpHE9WciG3ILkHNAOxNginOk43WXZACsmlk0uXisOxYOyPrF5N1
egCFzEx68BGYWc95sxYlJqGg0w3Ju23kq2xmGkMFaosdZN6ekXmlduf7ucWZ3Tki+LPrryHe/z8k
TIl4uZoTWLiddUaBwERMRk+p2DchZcpqi5GoflRQEUVSpttkovdCA6b7bmf8DowivvXuZlR8+EHE
VM24KF+eL8mtMSzFyhrzDawUreiZL+SoE3l+Alaf+TsPjW3tgNO0K0FH55C0y6qwj6OB0cVK+fJG
iDCXzuIr7SVKM5Qe4bwenJw7c4HDrFSHy4D9DTe3D4yFMYDtZiCPapIl11TxvKBe9ftHFyv/3B2W
mw3Gdb+ZU+XRmZ7uCwEx4g6NJsD85ds78RMPehv1CEy/VEwHlGB1piiOvKj7BLVG1wzKdfIJpEV5
MWradX5tRGtPQUzYOwQ2N+3z+V2wvdMeZvseyxfElOQhcICf0tPdmoCGS8Cx55ITSKuVqf+JIIkX
kFV0rG7DGDb4PKA3e1UD/yhWRBnNvK8zQriPeEAWDBMk8G4k/hmOWN972DzGt/xop88aDkrr0O4J
1pAdyGnsBKwnhbBLzYeBq090bINAIL1zDq6dqR6Zfz/azPx4knty5NO1CB2dWlU/9Jsb6OQGh3um
KhWVhHJ7FPmlDRYFZndCOtJ4YjTJ4/ZzRG/lxzOB6rwTZYomfwSkWiK5Qk6v915WWxWUXVrdt/N7
GKgQsCDiB5c3lt5YiLcF14JGTfgfpENE6OjZVC+TUyvDnhQrNZ5QPVPSX2+JN/C9eIM1r3LPBTob
9PJcoTCePFEMSmezYUWYRDWbWSW3BZjFKp2bKKjhvKWSKLqnJFD8uxIJUBUa0Q80fkmIuOx5Gszj
HCQKTfSr2ggvWlZcm5XKU0GJXHoZnviVDI7sE8ALLbyVMZmhuymdJVYiRueffXJH0eGR6Qn9WKMH
gGdDGQZnRrwVKxo+gNLhDScRgVihs52dsu/y0Yw6KWdbRdIP6XE80nLecp9h6wBcF5ilPNuDu5zk
69E795JioyWnULZZ2TcaDMxcAIof7JgL4qwKKPykdGFNeY2peCXZMBaQ0eWZhuRsePjNFm856zAu
Cu3vipku46SWGa+gcwCF93RFe4qfC4gzu+Rcc3Yj78pzdbSQMqIvKgUMCAPp9/2P4nftiu9llk6H
IOew7/VYkZChe3RScLbngGG9s80lCnAxLdBJJBNso3rk+TTJZNAiyBhwPH/kHxR3DKATDVdFOJuw
9DuTmgJRUpibITbQ/klJeHdIFnFdrAyh8eMQMNg8AHtgpBjqHBst0wnEYq58GQn+0dvpVYHUahAB
SfC2m87F2rXf+UNJu6W0bQB4FCn3/dE6Dju6WK9DpQ9Lr+iT9hXSHFiJqyKWmThaxNFx91iM15ja
OIedRyu/cjYyVZWhLi1/f5wUKiRBer96EDtLOkiKfFTP/D0RNwjau1CSKz08jgSkrc66qkpi8sLW
cfvqaVvur3RqBUW/OHX6BXe4Zl6ew45gp4hlBpSpo8FFiv9xDKsOwavuFTyRZHtprHZG5N/dqu7y
1KXgKmacY+LDtQF2o5tIGbxPdrB2h2Rlz442KhFt01aIc6xc5+ltuHbVIAwhBhfAMgqpodLMrZna
Sv0v2zk1pE7NsW3tv7f/0NWU/P5bPnzrhAXUpqFmN5cMZ7YA56nquFG5H23dZZJxlHR6LMJlUPla
EJqWtjfIut+vIS8l5SLmpDm4jrwOZY99IcQvhKRhWK/2NB271kx9vDJEPJDmeciLtY8ueCjZiWZ/
LGL49MJTELLyDyOGfiCe95dOUwk8HmdQgKM4awizdJeGPEBvxGw7FHjgTIdJoTdcLQoM3DjlWkdr
JfCa6g2cT1XOlw3y//buGzEsm5bgzRIF5EBWCQ1zpDyn/KIWUK3V6hfiAwfyy2MzaCugZ2H++hMV
SwSGZzDWDSFv7LDUJJnGvBdhvQrlzmypIPCjMwZWKpalQR+cq6a3aNi2wn4qqtXU0gUoW6kmk3XH
8+Vn4JgdHM6cuZLahCRaFzK+qxHL69Kg9kT4Z6W+RJ7+LobUqTbhz+5FKaKv4SqBXQxvGo2nanTZ
JoLvIi4PQ2u7LqLd+yb86FRQlPrKDRf5aIbnil9Wf43t32OD5hn+dgTdLkkhMPPNJd5E5hD3d1V/
PgvZ3eAnTkU2vp0eP19SpQUfCQ38Hj3XQ8Gg05vRPFnVy8DfWf8YQ+/1JMJOMrJcFVX4rqFqCnkK
omt1pSKe61P4Wh4IuKpUT+LDX063ramN5JF7zDbKnb1jZ5wqOMBrSw9eK0K7t31ZTCsXP8j1rNsF
PfXcQp8ntzmmMhGhEu97sKhUz5GiQLLx8QyU5tMIFh0RTsW7GXEkhPSjFLhrxxhRmzHpKWTAYbOW
mj8jF99oFlMnosMpU64SeHUAkiyl/BMndiMGnR8MHbuEbogCmK4NKpKkI8k8BNzT1uawsaY1cCEt
EmIEKDOkf7xV7HVj9Q0SHHGuwD/8HuTyRR9O9+RhIHhiQ2FDF03Vq9siIspHWrIg4rijUzShJzgX
nnYnY7BlgiG4/laDM3OvW2Cmey+i7M218cXNr3tKOrNOu0HIVXXhhnWU3WdIrsfILqFxxygOzT1Q
Ys5gvfruLW8aZKwskSlm/+OgyzTkMa1GDqajq7mj/iOvxTevvZAQK7zHn0MLGF1hYTwm1gBRYZ5v
LhFfRheytM2YY9FFmtBDE3wHfd87OMQnL0S0z4oplzIYjNTAHrhFw4cbxfLEdr51WfKP23xET0nW
+N52ZahNvM56S17uSg3mId0mdN3rO6e1kAvkIYlc9W8SLBV6VIWqtY2R5OjhjSJwfRQwExyd7ux+
zHJOYAEcEWv3wQA207tSOxuHpRBoso0RZMv3ThCxGrohOujiioGZLh2z1XEnIYQnTaDDahQCQMBb
WrqJXVVXOPx0Ji2LqhjtyswX6oL/XfFL5P3kcLoubhJYES1ZzpuqM3kvV7GupyezqxM+epOmrhix
UvbEF9f/q0OnKXC5V4sF+YFAnQfMXlrekTKKF6y+QD3F/d9nm5EWgAfmKF+Hqhzhm4+/Ht958r4q
DxazFXOgkj/BCtfgYnwcFxJjyQlQoyHYzcICJQMpjpO+Xl4gbkUp4rPGrFKkFTpNNx41fD6cRMGo
Hj4rNL4K06CDG+HSXcQmXUSYMb1lBRKz++YVkT/lYaBa9YO1NhBVzRgzHNy6i0sEJsFwirGLYCIs
GHz+5J08Xe0YofdJPp/fKmErsFsWbE4tAGHIBkqAp4ERkXbDsDNM4MvtkUWmnPTJPnX6U8o3tq2o
abgUp/9p3JWwPievAmy0cqjYDWxvXdgUEr1ZWyf6R71WuQc/yrNlFIaIMNUlGb2QQQ7l+HbyWDNi
c8SU28bQRnC1giqPzOhHHCycbfXUGciye2BTgwfTUTuDJzoEGWOE1NQkFsBKWv5K38IEtD2WTT8P
QVjq/u4aQhdZmqq1RX0FU98R72846zCQfAaLEkpbu+DADvhsZ7YRUtb2im34NaI25HXw1z7PUfnL
8+wV6h1pBWez0dC3/TRsgYeWEq6xKd0h6FEMHDvsVEdnpz0drziFenKVB8WJifOHFZkaREtQfDB4
m8JWTLR+Oi99Ig6QCTqVhIBq1SvGRoLxwHyiTbyf4FOc2VuZOzazxrdZTHlFB49Ej+YKU90/lYVz
KIU9GiwxYS2v33BYeuNK1VqorGFgYRtyg03KuG3RodMdFjDj6KelaN3+41TDpXZfX3OE2P8WkTZT
BOuwkYLvLvT8fwjM5LHL8ISFXyDpShPGv9h7/VGEOK7U5kkaW65z5VA13QJrkLM82xwEYefCW3Mq
xId55MjKdPvfuue+NnqKqChaYpBXBXNXp1sKSKA7z0+znOtr90aA3v4Ti9cNE2llGitp7Vnp8Bos
qG84VINtqo8mmyG/rV6mtZEqUnbP6CAxSxHS/0gVMxRZX7XNBqED7FJnHqo6WjY2J0R09zdvJbBF
+HbNvQvEz/a9MnFS00jpy/Gd0+j4BjPZFRIq6mT6p0QbLlloC+zksyD5kU38gegNyPUikPMQ5ZTe
ZRnY94O432L5ZL0N4Dl1Q2088FB6VP5Wfnl9We6l6ptDErasqfkg3dRWiTPnrfs/vQO7z+X2xBmT
Hxi2/QrgOJTHWFdB4Qy2FAkijIlb2bWiWzQPLVn4P2HaM42I0A+2nCxqBw0oUNRtar/WquuVYiLU
sLewyBpuA0/shiOeHN+N3LczgH5z2xxfTPFfb5f4izzRPHJjycIw+DFOC0s0fQni7owImR2QZUNn
xzenMiQyaG0SDZhGZK/sSPPgFVyhEfnICqKx0NIvp13lZ8O/Lmp9F+sKNG+6fycOJIP99pS4Esaq
v39tcg970YPoq/ghcg535hxhy+hiTrsHS7ifs4qr7alV2fLSyLz+R5GyfZTS10fPN3dyedEMNviO
hlcvDZR3z9SUM1gIWJhRmjEccryqeBhoafxKsXxColnrJCxqFbrxDLwKzQUEjooiZ+DnT5WXrON3
adA8kHLhYioT53bUwGI73edwA+3HgNq/FrWpgJVqaABcTRZPBJ+jX3DIsz+shMLypMyMJZClFvOQ
uVSPnr5d+hEddZdAvGxNXkSXGgi5aEHPahPDiuj6btzywlYfHkQvceobfEPnKpFPIBV574u1yxyI
k7Zsnuf8OdRm0SCnsCkGMp2lcdbPMItjqaOjqTDIViEU+0XOBal7uvB7RBHraxFcQZi0zdsBXv46
9DM/UdDZjpr3RYTj5VGsislm5bBi4rPQImJQDDf0dAycjiDMXTRBDWpCItnuJ/fFZm3SSagudwv1
TwmRW5WejFMoTdQ2oOpa10y/6JzKcdaj9PxAW85//XUl2/2i3s0kb87nByocDVU46OHtdBiWIbK3
d64wRe9WDiy1C4nB5dddX4LYSIO6jBGLxZ/1cLyBMp29H0rKxVE+Hu88IbUvKLzlBwdRXHU9qRc9
V9ealWPlkMU23Yjf2/xPobNdGhhG3HPFB69YpMnSj9EZWMJ2DWvbpsPf7FZINygq90MbF9c4PQE9
kwEfHj9eLPdrfSAoNAUAWOMOl1gmClV9GG0st+Q4GEanXdnKBQr4i/H8yV2pLXVHE/XXJVeCJtcs
XHn0azBa0VBmqlkC8+/MppUvpY8Y2mJd5myZ3+uHVMRLquUiC2wkI2hS0NuvQrw9INcJgvPzGZct
El/cpYiiyWChgv1a7OYCyFmUE1KPe5A9MMtKKjKam96hKkaZEPZmIJI8kG+n6r2BiGXatZhxgIk2
F0ZVPBVXvbktlwnHIg2isyXjESsdyOPTTLHY9oynoi9RiQk9JmoO56jiZAB0KaXa88yg4MKN1AB0
p81bA3ExsDoR/Eea4qDdqBa5P3/n4GLQwNdxCRyMM6FoT/xwDB3OhbTCymvhcrnFr8z+NbQlhTEk
qEcujPPFjqitSHsylJ5It7BJS3k/fYJJb58vfA0D5RD2QJMUfrel1OMksPmgPOZkRgwUaR9u0Wxc
InIZ8F9QlOwMxr15C7HyqZzZnOcRzc+YKc5/I3Kq3FIKFJSbzfKuair8KzoY24u++pkdNvOa0UMz
WMqqk3/oohaqmXAzwcjPFkcNS+xDkUhZA1kkNmdticqAAld/R+mRQiQwFo68GWYJzlaWDDwFKe/C
B3KcMr7gGHn+a2i8cyNZFKtyV9j079GiQy7bcC3LIYm7n6PYRVpxgWaWruVg8RNOXl9nvYJk+S3x
fbDpZJ0qFknTar+tQxIKUowdBB4ENfRVJQe5+4xPSp2oSzx5uiZS7vWjKB46pCzEOJpTYUqGKJdw
CFJoPXRMKAo4Uq1SgZErw9TuBWzFa3EqEk3nFy8sM5y+qpzy1ULRZ4bmX8UTrZNNOs85hTSP5HuF
clfAeGjkj2t53KIe5anstJK/IUJuupaBAs0v4iXuwzCSmKt84yTwtiLKxjMNbccky/yMJMKkt415
FP4BI4ZVYizTqsK5Bstm8odyUmuD+pwfivflloDTMZa/Jvutt9vNjzsewAvlPnT7OIc5yLXYqdlZ
6C/f9KhVqKZd1wtqL7FkSZle0K+346221H2xquORn0I365c/+bxxCJuP+M8xD+2QtlyYO1lAjWh1
MyTeZteKqRvu6jfogwP9tuWwIydIMdApVi42pTnq9ZOp8aYVyvgg0OevR6CuhbGAU9LQdYEfHbJA
scgimUn58YASDFkYqlpluJqbyEpmvATBmwT67eGmqdJUJnpsPPM0jgwGMXy5iWuKenWE8GFCjsA3
+HsWPY70A6wk3iPumwBzbx8O1w6psKrEjxCBrx2e5Lg5gABXQPIJa4uKA1mVXSzvLwhY4xmomHM5
XEGADb+sPPw6xF3i+yNTKI5BK2kYQFgOow/bGtdnLmW1qPUZ+Y59s5u5xhBPouEw52GV2SllF5Pv
n6a4js9QJnIZfcwQYqxedE9ZFaiCq+lv0wodOlSGDRE58/kQImlRJEeUL3Hud+3wkV1imAntH4Mi
Jm8kYAgD609rEncHPqqtI0IG8PN16JBUwhjnwZYNbAMvz18ql/hl/n2frmPMayufPLBV6Vql3DRj
OjphEcIfqStK/2LmGHTpUrnz26G/cYqO+lMBJlVLBDZc5/FoQ8RI9nuE5Ypmr3GfLwFIy6d8pDtW
RLXA6El2Avh3LHj/H719/gQJfGkFBLic94V62lD8Q51oUUSM2UzUuQz1Yod4477zn0Hh7OMFxJwl
oYyZYo9zbmO3tkQz1JPSESdW/wzFLc4VsWj6NqQlKYoWCxG9bC9Y8fCmL/aRDvq/4wCrzZjHXYE+
nS3MchpfaUCoj4JZPZhGTthaArsJ44TXw12hthAr35Y5c2PBYRcdpcTkLyoJljaHqN4LAHx/s4ti
ePieihySTKvub3tugtbukIbHcGGnYog08Uqn0RqvC9bplOp0Z1aDvWfazdL1/r2TmYlp9/AWlVXq
o416Plk8AeezLSczOPCKKBqvjadtTMDAHMrpqZxDoFlPMnw/hH9wxE0N4QoB+bMpZ8RzUZaUpreZ
I0muKmNd6LowUcT0BIYBJIUhrLE8bau/6W9ta1jaV+SeUZI2gNMAc2V4Y2uGlRBS+97l1mo9N5Fy
KyVWqVuF3BA441MYtKavoa40FKlRN2wtyyC0QEAXgafrUNThikIMUH4iDiNZu9suPFYYBM9AE7eg
ekVM11qjue0OUVlcptkds9M9D0DZd5o6dxb0VzXjEKlxYf31ihP3vvZSKLSupqheKDVhgaxn8nio
g7eO0FRkYx11XGgf2N3IqOCpKoGH7E9IcThCrZmi8nOkhkTvI14zeFlOaRmUr0uaBYh+9d3nsnQ8
zGV0Qdxsa4az7I7OlcUVif28QKdRBIGO3CyDGgKYk+Igqpli8JxDzZd9TMIGj8vzaF0W/qjKVDLw
j0gZ5LpfNmsF4afPA9oRYxbnNDVYRpv1sOPm9M8cuWOjMSKeZ5/oHD358G1xdsrVMe3AuehVpaML
h43oqp9X+Lfn6d9ulSTvUBXty913H/Y243POr0KiGeKEy8aP74563sC3SJzqgU4FqV30OZqBHpA2
dbi8sbDmHNLzTm4lpzXjZIxd5xX2/ISVvA21KJtXEDWeKk7/UsDW96yakNtRwJwy40CxkkzDLDG4
eWhUhgvRDGBtc5sSAmAgTXrP5LZt8EwQa/8f6Rl3P23nuf2Awsci2AJpRfL5gnLTobwEwDN26PLm
MYhgj+UcEQv5lfP/Y7tteHs/o7aykXfpVDzYJHASDRCAE0FkVGjEzm22fGNUrcWb5LO2lp97NPM0
/YAkLzhhmLpADMPLOj4dCJ9I0aVjldieJetf4ChU9xJHSbgmmxVRcUd3e1YMdz0CYEv7/zuKwyao
qokKaKxFzRTuFO7ITefXYo2RbLEBAu1bMXSlm6Gsk5oPBKrzeUM8HKIMzhRQacrOk/fu29MrjQhJ
rBWOP0UpwRs7qj3R/PA2SZvwdsOpoBC2krserErTbPBmahx5TCjh0xdE/xSKiQEwyACXkena9G9w
al06bX2W8JW9ahOu/3kH5+vZKc9GZkkJP0H0TN/R6yGmsE89vR/fDwmIXKKehBDwIsK+uMrXu/Zx
SYHKUE2zU45LYgh4kEHM3e10VNKOwxfVgdg9M/D/JeWQXb/AfQXwLcN2lrjMA9zwg7CYF9e96k55
x12iyIJjOqwioglJAA7Z3u3coM1o6zER7twBHZtXNZ7DJhlPkRhABne3TZbQWETtF1Qj5wJt1FdW
E8ppieuSTlbcrIh97vcrTa48x2ehR29Aef/2Tlw+2aiyNjZE9QvgtZ/dJbPAERZU0AtuIjAsYIK1
1slYLVSoNVDhzI1fI6VP1LhvgBP4TGdNBdoaTqPfR6idU2yNF6nrbH8EkkOWwoEpGNABOAefaTv1
nCnjLt3DBPyIdTlRcf2q+2KvsLy51KyZv9jkXN/vMHHNU6DZjrtrnTOOi/hJL/q6S/9ynQqaVRw4
h/plN3VKnazIsP+Nnbn3SyW+jVTcSwAAvXRa7YhGB/FfMpHmX8C8dlNqJFPMeHPlZsdv+EbZFIEC
bGRuLoajq47UVxehxKxnDbN5gSpIaaaiPJEEghniobKEVYIyQbJ6XEEG1RVf4FgzgLzxv87JkZON
CbBFdnD/YyR7Lr7uMtIIQIGveCt6EEIHatwaZVYnH5Bu/IMjXZhDh0nRcNrrLftrbaRz54BqXv+H
SnHUdXqNw3sqozGHY5KFSpbxzGb6zzZe6i8Y0zOq4xRskbn4Eb7WjF7/aq+0ZlBiPDTlSUIiuzbZ
aMUACmK3r/GwtnrnVlOCw7znd1YfZb5y17wxEDAByObd1wy2RfFFKMdE0o2DIaL/9HFGubXH/diF
SI5upGNHavsN8XPA17suzYSogWRVIm3OtIaS21lJ4ypelYGmaC59NpXml2k7CZyBORmZ8bDS1Klt
OfG0ZEi136dqfOXpUZmDWhd4w3yjvQGgWw6EZV+6LzK/RODkYEC6IljG6mI4QdDew9qlC9tlQ15/
YyfHDZgZ2bwRWjh8uMWEAbbRJNKS0swCcS7u+1NbJ5RGyMy4P4CatcojSRfzUzyKva6xN+bATVbl
6F9PnEZuF9jRwjZ0H+4GGMVcrURCO84xauOCZ12HE+0P24tWHJzvYNDt1Lwd759yPRTYrE9ZMjdz
jNAdsR4kgwE4/bkSX/H4vkC58v8ozet1UERANkD8mONJIh41NREgX3tn6Igcxo8lPea4YDQd4SA1
Etv0gFdto4hHSsXNfMgSgHJemUuWLUqWm//yMSdAgKFuQr68xHQG81u0NsLICAGUma6AlYzWYpfg
c8rzYgmIWUc9I8gu/+J5WxaEGdZVPko177NknKhwkD7ffBYDaXBb/5wNSgdK/7G0S3AHZ/xG1lA2
TXG16A5jZ+KidwGp/YN/obfgKsmF/gjODvLBKqNNg1UlsWfCY+X2LRu7vk4gjAcvwx4K8zGfBjpF
QbS8xzMld5SVErJBODH0tvSkSoR1mq/w9eTGkNhnpOjfTxeaCq91OLNDRT+IFLYXlh18qy8M+WUL
iZBEQGcdpL83FBpJK+pD+8kqKYP7gCSitjA5T8DgRBWgI2yjrS2BrdChgUcj3jvitILpAifauB/o
nLdvsjqVS0+RYBL10s+PUF7o9FnL8IsEMhKFaIQEKOd8HfNc1AAhehRafrcUj+2yqcbd+yJjVJ8q
CxNVV3fN5Oy/fKkhFJf7ZjlSDiDDEa2ZTJ3kdnh5/LWuZOHAQ4aBdYOVuRCFlFxMqM+TkIKoDXld
MLmQrc9GBpWmZ52zbo3AoASPV3Y0BVHlxSNrCWmbiHeqkGOLoBmOaQJ5y6eLpMwcukNkXgXWy5gU
7a2DYDZyXQbc+YfqtX74my2sdpRTpMVcsO5dASZZcL4o1rlID1hmjzo+ESEPtewDOqEkr8gEj1DK
3bs6RWrW4U0rTtKZ7xBCfD5A2Eyu8AXH9ZHZdSf9a2CKn3U6mAeX3590nIN5LFEJgc7vXplrGiah
UtJBFwD67Lg1mizn3Y8a924uqXuY96fo+DPmtmXMIhUem8xBce3W36JXPEGGDTEk3NHj0mHv9mnK
Cn18Rh8QY/jrZ38Bx+N08gyvBLWcf+FMPCMGGun87WCHHorLwrr7156rpwMOXpirZw2bhBXz2Xky
7WuMG6mFZSYA2+gt1RjOKmQT/E8eD0C9kyICPl1NOiQZdj8Z44c1TPQYlkZw1ynsoLcjc1urCJzw
jVNY0Dq5B3cCk4kHM4uncWDB4LxS22ilvqcHTIo+IiVYvrFptFOFvjIcxIImJlC94xLyXrCzU9P8
BewQeuyoO4rDqVxKyPcgviTkCKeKjGDqqoc+JJDCdSSXrNwf4La0jvzfXqcuT6CJ+k0EmAj/7tYv
qUXdw5TtZ9E+oad6bMAE034IzwpH0NTtBZ0vgwHDpFZqDdit6zMzSLHJ+Jn/bTkrWDePoEAUh35D
gKhr63g7h6uysOQTHWVx74VsoyrmalkpMe4i2m+tJHNH2BcnXSnXExjoO81txfHbzfVBYorBGput
q5uXM8nZ5tTGlhpx/VJHZ/EeV7ImAqhs6oE8IeyeHm1vzpDu+NLZbQrSO33ts3WjLZT41fX1x4Lv
okqKOpETAN3WFjV+Wmqz8NZY/qZ5xCoHuArQEAcHb1lLTu5eEKEXsj/IebF3xhKFbhzBE2KrjnWW
84JmFdfH4Vh6SCW2dkhbHYleyvxDfr8mW+V6QyL8JLLY5THQGmEWDwvIS1QM2jzJcBtyPCKhX/Bx
eIjmTGuDhy6hFToJkWzeeJ1LAbD2MxwDaZUGbBUZhRYkbXJAP/Hm5leGV3kczN9bdaPhgf/inN/q
HqLnYDKJeA9OQR1swfXJtQEkFqcXQBUElkqKkLIX8dbXgYRxqI4gP9+2A5CRZmlAqHPMIrBMy4tv
/iBt7PLj2Qbxauxug9uPiJ2iar6V/jMywEfknWzBhPYa+W3TYK8TncSwi1g4e0nBflEIHItjyVhh
sakxuTAJFV9/sHOWeAQnHMBpFpl2j3tqIqHMNSizQnXm4CDg9bckRCTrWKUmDfLrbToEIkXE3gZo
Bs7sVqoWj6w9x4+oC2hmNNRl6zwfe0WEEh3ZsjwcDqvV++Ne2FMspgeK5AnDO5pdcGXu3KTIFR5F
3FTWfl1zCCSM2ZMjKbg/hpHJ8EDkhME0ljTZnWXQna4IaKA1ggG0zLDSxS7L86xdXvCniGnydi24
2nYZe2vFnZMye4BjABtUGWXd9CgW+6t6tuJXJW7Rs0+AmKQlUGXyD0c3UN1Oq+ztZqJxpRB3YmzI
VGOl45xA/pmU1LFqJt+SpW6P7MCMg+0xvzh9vu2/bHGdxSMxwc7PLSiRmHIMSKtEQQUCZmzeCg3e
mVVOh1BOwu6t4h8OtatYr5Aq99K5vw7YjXE/nD73CPBfx3spSP10GM/2SGmtK4+5HMEbmO9bsxds
x2sTLiosyU/W/SmX7S5ozFC0FMggb+gaUIbeZaHTeE/lycO/H4LMTMqftgLQBFRuWbf2J6SWRsIA
x3Z9CLRgbnD83llpg41onodjZBNSnXGKVhsoyS/NtEmrfYweshWdsila8M2SSrbu8R9n12431YhI
qWZWQQMQX7TgMXCwp0d4BT0TRAbbje+HNNE0pX8BBB2xfQflhZPlWrZdL1FfZ04Gv/UobtwQ+xwF
X4NL0e0vaOk9ZL4zdCL5j3N4BNh36NfHqTJyveKQoTHT3x1FfDVZOc1HLlq7zQj5+PnITyVw+ZTf
zbCiTXXVXn0mmZ7Lwbar6GN7J7CMTXrYathbM/B+aprLQtq2ZRH4MyTNIxoozZviaeLIBPcB9034
ssh/oQWParP3S9Y7iFhfOpor3zs4DzOhAyMlU/166xLGbf8v+w9TxvIk5nOLxehkfRZwJymLZieW
YDEFq6Z85K4DHryggcVIfQAw7bZq3Ig7tmOfDKxWBRWryIxJTJPeLyzkMCSQZgiug8gr8xs8TP06
Ccr0vpmJR3NxnNB7GkpmEoDAKW7bdtLlHt1VGZyj93WSTOr3pdITggzuAQItxxkP5ddFUb47nJ2p
l+jgvSPaHViqQhm6cproiwg6cdGcsN/iN0s4vYITNTpop70kkqQ+PrHHOzPgYYO48Gw+DDKG9rO6
wDMYyjh2Ub38D5WYGAcRrRToNRf8JpuCAcHoytbkIJytARY6e4luo6Ij1A29tu8X6Jd10ci9fGE2
p/jQWrdqSbWOrr+c9wrEwqO2Mam1pHEok4jRTDfxyLkzF04Y+KeNJGJxvYh2htw5Qo7cMmn3Q7S4
AvpwxogJSEVNHi3HgedmPA6vl/faPPD5sJUGHj62SzuKNyvheRq03HCNjC+kZJrScNVOJQeP7Vz6
pKn1+9aN63eP++8ilQGobYM5r5O/erjUVo+X3KFoU6uSmMopJRdsonLjcqZZrGuLooj1kByO/7gI
G7K5scxsdQEW6dFtvUamftUtzS66Wr7VteT7jlMtUN/5x3PLPsLPfEGbh8A46y8aAe1AmmQIVn6P
USqDk2706a7Est7RDkh3gUDEmi+RAWASz/jmDoMq9WBYDeWBwmWujOvDAQ6V/GZYeZNfM/0LlpqC
qrnBg28x/7mZCqbcUK5aT/jVDe3kwJ7Bjp3KdPEFnis9IlDPOES5Q0AQ7giQC13cBRBf9YgLXg4A
gfSZOpkTO4oPctVbnMz8SSZzU8N1oigIpK102v63XVN7mDXlnsPKDWFe7kFxjMCGUUIw5GcJojC1
7u55XeXvHMCrC/R4aMAXpOVl4cynuhTz8Zwv+snH3cOnTvt9uGw5UjdnwqJ8NN39NpqIy7ZELJos
8arF+mhVsALIlSWpK8a1ykfQEvjiORr5YWS8qPUFv8AcpSGGybDkNUZHcOp5XvrKCdI/n2dYuIDH
YYesUca/KQZ1+emAeCsONqzKas9LbUJjv81pVPSCao4VgnIto4whw/MnpQesWlC5XX5tmnfcJN6R
B9H7XHBh8StBaLYSKwiKz+E9Lf2CGxwqyEifvs4MiohmK0Mk063mc3WU9PCVyOu2LzJ1f8M8rB4Q
c5TJoMWCZbxyeCnRdOv6mMJityhP0eU4Hk4a3kq7JV5mzZFDa81nYmWLihJ4erINfT34JTO8VLLT
o/J3XxxyryJbvQmsNXDWqBCQXJ5dv4yNhcceshQbePuZAlTX02EFzfvhAQKsziVAmbOPFF0ZXlOu
DEt/6mQjrGkHB52xM0Ku8QhIzmnYF4gcJTqlV4YJZ07HkdszqZac/yuQZgkPyHEM4GuT2ZDg3P+r
gQgsmnkUX2DuIyChmg0TvnfpGObGAUEM70hkkZZI+erwu+eteVDvWU9y5EXjy/jIc4UG6Kfnh81h
ql9ilP36CWS6CqD5l8f4tL9gosusx9vHjpN3dMlt9+c8bRWNb3NSUwwT+qkZpBPYzYiCv0Sz2YY3
reuVGRMF14xU11/cV5vXyWRuO3iJXnXrd++1tl3R4SYtqOSyh3TVfil+hFT0MVfeLUqtZ/t/Qzk7
kkXmnosQt5U75zzBl+RSeesT5acSKNdkGSILH0H2/QZFwj0wsfXkLVRGpaMVWKfZeSl4kYp6e1AX
d01qdGGwy2SkEes1MF5AqBzBVBRePH+jCWDZm+XuK/z+BQmbrUDMyMay8OIQaK4cXvLL96kK9P8Y
PV3K8ju5Z02obaGFVVbTM+lL+yPXNW8SVUbdncM0ZO6U724fBy0Pbeo3tyvAk42lqW2kDBo6yKuH
IGYuf7Zpth3OQbmeQFHupfSai9wUrjczfkFH8hCRdrDSUyH9pKIJzf/xNbLKvPaDdSppStlOncPR
tpevBMeWxOdtV9N3MV4sWn2/zRbQx3c17OpPdqf63w2PSL98kwPQLJWEqtTwJy7yAhN8CJ04VKK3
7xvkVRVZiA8hx8IdM0xvt4tb6MH2EXsZ/BSrHgVtn1hao8SE8wLVZRfRE4hUEpbJcuXcXrCJBFBM
YDtjVaffEJ2DRutz6Z0Ag6+GchQiGFKW0DRgdaKDflrnKWF+vbPwCpHckPKyjNQ/t/2jECGvw5if
Gs8vxqcWNcOq1vtLVw0Im/Bea9r/UhsTvpiCuoQ6VNgfOwLXeruWjEp9ISzAH57CjT3dmoJEEYQi
lATVkl+gFpQsyeOKjFAOlYSOYT+Qa1fT362PZWiPvDlz0oe35hw4DSRBebR8i/9gBZHhN9rfdjex
f7jgZqgKQM1n5Bt2cErGN3M/6u32K8GxZuV9vlr92EFJdcTmGu51+IoyeT4slAh8gWlhsmHh2gf1
Fg1S0WXmdlYKXnnL+KKUlOHiDoAmhBF0+g+NAinOwDkcaugBvzDpLEMjW2CSg/Mc+X6160BCQG5N
uk9qFaCl3xl7xWc5pIAtKwYrPlqRzz/VCHc7BkTn6LdS5Kc7NjLdnt4EHdtnojODTWJQ0auVPXsG
MWVsBCXG/jLFkbw+O1mR2ISiqmg7EhGa7liJEpYcdU1p0ijIojyAPeYTx2NL9Ddv03BCcjdsHxN1
P2Khii+f8k7+wL3MHp612JzM6FmUNIoF5yqEGyMx4kXsVMrTpoW7txszLGeSCg7kiwpW7CBSIkFP
bRXjdiQOKK6m7YpO6swDja52OcajIcbyFcwynQqh+68tVcEftf/phBew+jQoFG1ansqSha14nZmq
jQ3KAbtHEphRboghdlH16F5fsjGkNDpkhDj1n9GZCsCrYXohhT2DUUH1LU3EtWzbkWgit400wQpx
7TSiaDdxMK8csw3+jb0vSm2BbTvA1gzFnh3viWdSLk0J6DrCXufrHDWvZyygQ2QoHXTxBrUW+jQo
aEQlSZMoOFSi398nhd6oUXYQBpygoGOv56B/p56KYSPnQ3jv1yD8TD76ABXtKfSrFSRxa1pa4vdK
Scbm/O/ZvxF3w4HK2NloEkpAmY3n5f5Fx4WR6asv3c57F4JEgYTsNOcwUllZEL5i6mvKCDYWfOxW
HXQDsOueOdvYiIA52mJCOqqEiE4VKbVQiegxSafibmQt5iGCVHjQidteUWKOMXCY3KryTJ8+IG5G
5cAHd6rDInDNT7FIRfoLoL61qwUEu3ELrAcCY2x0x04EwRgMqWB6i/+NVrEumrTQvYCk+WlOanDD
+B1JvgI3d1HMMH94guRYmcm7oDPEw7+HD+kY+NADP53Ehpj8qtBJJr89TgR8fjCLLCKfF3w0CZRI
4CvTiz4VLLaRQSfidGs3t8EHesUnQM8FxdJGmKEbJ504BXFO3NVmTAyizO+ZoPWZmUMMT0JVxVk8
ntxyawJ28FJuCmep1o/0qC62hxkAiyZ8mZX1cZqsCQv7SkpQqLqhnjy/n22rQjKu3nkWobc98g+Q
h4vMUWQmT+pgTPkuzFVfcxGf8hjBV/7EciQmGapimErGO/zMUmUISPG1UrBr3/1wNZs7Pqz1P2iI
vZnxD2F+lB5szH003iM4fEBH4f8VBP3QGfnldKPvmk57ityuK9fd6Ww2IebyCA4mLpn8LUB+xfjt
IL6lUmABi8+mlY3dBNlXFVpBeraPXqE/40+Nj3eLGh8qNGaZq09gOQmZY5eIBx8ViXI58+u/IDzv
/JeRwi/tORsspX3VX+VmItAK8X3879ZCejOZTo5JQc7vdSqF0XGh52j2lyL1ViI2ImrtcH/UFYLB
MZPkzvNxmhyoy0K2xvKLSI0QBtw9Bq74rbJDsLJ/dNm15fzSXMdKBDepfK8nLWMdBew7N9i4cN9j
iBqA11Tn0MtL8TkyZHkEGWc9lNv5efcfPzOeytYGUD0d0sJkrfzEyPFMFlwgQqSm+X/1iP1k/7W1
KW+V4kUMhhiFTo85tAhTVR0YeElBMujrgKmZ01a/55p31Qcj3W7o2N+LEvxSgza8S/LsPA+lfoGS
T38gdFvH6H1Vkq7H3SspuXoQGiJhzNgQIfF/MCpG46A/DyRtexAJV5e6e80QOv8PDJ7E1ite7r1q
/Wh+proRNaVUr6VqMv2bLSdJ0uBEDTGInGTZUwn/Z9vn32Gf3FiJk0CH60aDvatzGwUS/djC6/Ir
kOsFSgOr+4R0MY07LG/CwDhBWGN1ZhnQpr8yazE6bqzBY4oCNlM8Ycl8kfaVeHOqjYwvngoRk2HM
8K+sESRBW4sidtr8LR9an25pBGfxA40tAYwvVZjoVMlV0/pzT662zl+I8I5uc8MEwQe5ZE9jQDXX
/e+glQ15mcQC/3nanUv8bvwdzu6Wn58ZflsQkoWc0Nx8+xto1ezCReG08MeHFp/eAGAvDfPAGDlF
Z5Ctv6XhTVkH0pQGhc3VpuNFYsC34W4kSfJFRLUOp0VbhqkTcI/wvJJ7kc44ygmN/A0aA5rKFRFp
XDtVzWETJvlHhNJ2EiRHPO0JQuebsWPUc3tMC3mMgN2ArL2sPPJ/F5iAvs1HibtOvx66htMq15Xy
GucC1iUkSkto3v2fOSPadZ6SmGMlCFhYJn9skQL9KC/7ou5HniWhSWgBkzLkGKhWCqHPKccFzeLB
3uzM4y3VaXyinn4Tv2klcUHTAtuJV9gBFRlDwekPXbbGv/iWlPLpytrnEnO3Z1ELsYBhEfFVTV9M
BYaHjbOPTOL3eYfH5wBxRB+MP8ySpyh2dqmVtAEcvqBK36bXCwcy8gWKFYqEbJzZl70U1U+56c/t
5vx6gPfGADwQ9fidWR3ek5/FfFwNcrL8U0Ytbz2ZKRExAmz28sCS+Yi6F+DDuxt79SzlQGdUaX6+
P/VdXoSbAZgXrHNURYDz4cX6kJr79qghvqd0aB3jcAcyZAS28eJAuskhLWNnqkXVZ+sjO07gX7ud
aVToAdEHuzmXPSPGcSJ4PjAodiOsLWcSzNaU7lGQMvcniZ4KNBAbb4RmKczhd5xzljMjYAaSto6S
E95go6dQ5l7m2SkXDuQlwnK2/C90WWWlfg9IPyUmM670mCIfOC0lqGPqyEvHDRdZlpcAuzZUHtMv
WPdbo8qm5Qf6rZt1iviVxrqILFZnLW9LpEvTNaq7pMNIrLRx8vcVMJkggSwNpkSCnagc9ExTZ1OH
w/g321wLXI8N0rYnUl5Pxmm1hiFghGNJcMft4Oxm9npzZSSH0IWcI1Eiv/zKbz3LFzbBNkwoENym
+inBRQD+xu5EIqLsi3kFj4OUevChDjkZku4k7eLYs1MTgm2XydJ2CPpBTzwPdSD/FgFQhhNaUedf
yIFaWGbmw1PSyP2/93uMYFHHYv5XjCEFXc5q8Dp8Oz1oGSBto9U9NL/sgXYxIe3DfG271i2idpnm
oeDI+DyAnyl2dzntvBpKOiaUILkFLEyXeJY+LWnszDlu+wNRyB791CadFgbGU9XPiLDxZZNp+9EW
wboyXzZ9GdTig+0WA52GPrtikKxACk2d2PyjqLhP691scCehcyFSbl3f0cOit12eH2dHzxUKyFqh
+puCBzwxLzElUeiohkdST4tcvqN+PEX/5dGdmzfdtRde5CLDXz70iOuPae+1mZUFcVHINDdWxxwB
hvIZMJ56ESttR4MVjCYHnCxAF6BmyPhMbTdSSt+lu+szRQMy82Zc760fg2twjdINI5jf9cFVIxhM
0jWb9jdT5gFnfV5VcnuKJezs61rFeTuknJvOrenqt0dGNl9h0BtCZA386QtTcjvnbufBi3PyKy2l
FUXnPpmOnvIaAGj8jA+/ek+CL6OpfSrf4efsWdXYOwsjsVHEAWbqLPZ+Vj3O1uSUPqD3x/uFxedr
MgkHJr2Cg75JwbSxT7we8O2OtsKdFVpi5+EsQgOR0V49a8Y2/hx8yOiYRR6HjL305lfpCiyYZIGk
wKoNGFu9eb+PQXsqf4F7YfeFLg8soJC/2qZfaaKRvvd4zJtCV6fYQQMgBLcWZ48PaQ2EEkIIDdj5
L7h90n5S0Gw/EAQ4t4oyxQA/OnkE/P3WlJN9/iRjSj8a2do8jzHFsDeotAR6sfFdL6Zy0XNg2/jo
SfyK8EsMlRsKcqY7DKzT1YQK1bcV2uZZfJE/WdBLGXzlYYEp/mzuUJlIljNsVbij1RN7u3Aonwk/
jI6iy4s0ky0h6hcQUeR/lQ4oYgFfRNl3dwe22tQsu8qd2z/R5jWnonp0wBBYWiltFVvhy4Z24q7v
Hr3uevWIoxd8dk270vKj1VPJgheB6F2xzc94zmkXW2MS0ZNJv0QmMCqADT6ZcIlMbZaPL1xOv860
hsVMrpnNIkQOcp4D2XmSd/UV/K5q2EzDfvCTu2nDXZj3Nu7V9LHtxIZeKezeoKtFW/iaIQzgN9UK
jo94mYR2edOEwT4qTOivbIbkMJqDJhhPlRiZG7dF+E1iMhlWZk/gpMOIS82x4+cGyYvWMeE4wGNG
ZeKCDg9qJ8Jv9ZVMc78U7T7gJMfc4fmLqoP9xCwNDP2TztjHZslGCVmcA0NiopPqImd0fP8nvn1r
/CuBvbVUh1HRjjY4zDuaSSu66AvUGTF/0TVVZ7ivWozJea1qR6PK5g49iZ9o3Kc5tizbXluPYdCI
aP0bZP/3v0ZYUtn7QnCtW238dGImgqs5F9HR86Nu1GlQZf37Atd53F3r83t3UzVvkZHaA+kQZPFA
f9B+xpHng9Ira9gdVndliK8NBOt2r3xEm9aF6CVMVjiZDdIA4j2KmTsuIFyGfa/W7YSHtFySrOkx
Q6ZzuDDKF9Ldd3xzRAI7emeADaFYHCO3s9Pc3bnV/pHOnW2Tfakg7LaQzBKihXAM8EzoAFfYwDoP
7rswhbud2p0S2Qp6kbAiPrQcWnIRBbn7GGH8TXxl4NwtfzM2W1/Pf+/qcQSrs6dX+F23EVe8mskk
SdzrfnMx86MRkXAm2Ac+j6LZrLjJLuypaD6ZKbxZIs1yabLgcXgzPbpWW5qY+Gotaq0hI+RI9U0W
gW5wNlx1s4HM1ti1w3tq1XJJ2/7I65pRAP4XJTSFh867pX8u0My+61QKVO39DProMdl4bHJuIwfW
YwmlK98FInDwrMXIaRLPAROdNg9Q3keM4KRZKyKE199CLZrEQANVMK+aMkWzZDT+r2wdsQe2B+Rf
HrS73B+ZglvRDS92NnL1KPb0pU0I30hAjTMvNOhgQzSYOYTdh7FoIxqxMOP/xUm8oG79J+ZbzrPh
sRYC6PS7UcTIiqrk2A8rI1Iwqvc+82Z7/NkuYMLX17xZYUrwdVmaHtjuNUYe2+LPXybhWRehzP6f
iqLIt59V6PLcMGIkbDnxMDWNdFSZg2lKIZ9NUWzv42z+AhVgxjLk6GM6XypFOrY/+jlCwYen8Y5a
rSB3Hb/2SjvZG+c+zBLhoNExpu3OcZvAVhUfYhD71dBGPpDmunBu15ceIcEpzWGtGUTbFMp+6tDS
O5vlu8+6Ec4gUvZJDwYr6SdDaDsz3V+H4CT6qLlizPoikjKduqikt22IWb7tVFipRrPaMaw4ljVF
PlgB2mbrb6of69+qCMVLPjixjUZpHfxwpbiROQg8u/pWNoYO2rsVDeFoktocoMt0shg9NYMK9jwk
3caO6UcAwYXZlEtSNxZID/044/u2+ec1PnmKjeA+AkmGsMeu2ncCuvTW/yXET9GBakkzqV2gN2UZ
XvTf0EOhxV418UlWQ3PzC3UdAZHS5ZsIERZMFl8MXSZ5ytmhkdKWkR6IKuEtFfFsPt62p+s3DuLR
j5qJK9WdZE4XNKgMyWfVmS+j4q3HORvDT3c3n5vob6erCOMiFReqwtCwbjGjPYdAbWYSn3izm67V
4tOTGRxfXTA5kHKxH8vQ3a9Hrby+rG6+dTGXIDcpMNVDjrlR3fdwD6CQumtxXKW3F3a/RmotGgzM
IgF+v8VNwwXfz5W4/wHTmfhVNfe4sUdXCmgemeXlwXIgKjAalPah8Dz4sJuDH7f/GrJHNRP9gPpl
tbZ2sWITcSpdKcuGmDvwr685lDc1NCAVjmhOsUk6BfXA5Zb9PWpwA8r7Jh0UBg5XKm6bG8ZfF/Nm
Mbnb4AbBc+osZYck79rMUHAd9IyROZBhmvtxQkWWOTxlVRGrmnFNL4BpNbAVascYMC8JoSKB0B5/
de0Y1KX9fK7ynOA8kDZVnAv5F++r5/CtJeq95uTI30Md893vMoZS6HyXbPvra3plNcTgazw4rZsY
8AuRuR90+Yt2tAzhHx1KMjDo1b6AhGovvKtp0cqfZa4pXYGMlxIc6MaFJ9Aa58pHDlQJfM5yNY5B
gMpFnRkEAIAE9uEt865rGjHgaSRDTrsZc8sIzC6knzQqxh2wvzeWLMZnhWKl8zSuutp91M0lKz4u
yRdoJZY8hF7h40GrqxUc9hoIXaOiNRLewKeeGnZ/bRU9tDqoLf3ldklEHLp1PP1fkQY1VXXJMIKh
jq8mXh55yi5FmwS/2e8e1L7eby/Xdo42JBAe2pFZSxJPR9GxfQ2tb72j4XVWnf6BsRfWtsZqSLqu
83o9Zl710APp4+1Jc4oEvS5JmgJ+GKc9RFYi5x8j/9Ycpcr0tpC2a7GNL4nUr2jr/IwY4lw6z+6J
A3mW+uWHQY3KhCEQ3J5QufH3PqxOUIb+ARjenb0K/eeMRJZvB44+8pzmQNnMkRuREmp1nxBOtzcl
u9g1cDv+BNrfacqQ5VI9Kreq09UaZf8HIbnfWlJ9pk20xEBgsdc9WRa4/QdZQXOH5Wp9S5qbCh8E
6QrheWNHe8ZqH1YBtVomHemo+f/Zp5csIPli2WIRBbaRM+qCvWo8ufEYuPsBPGxZ57yu+uYL5hlh
4NrUdRG8p0d44UroUSo9RoqYAPFgOJisrOKGwAPqXVgiac80+wtT+Tl93d4JS9Wbtqajn502wYGH
YRGVbRXoQQely3KR3/2pb6kvJjnWZyccC5dZKCKl3lWOIyy/4Hq7lWqtJ9kPR9GyfuyPaxd8jE5v
TFbIE+YhoUxOGAkenc099P7hkLxHOgIdi5CbelD2AUcWDLRkkk2W9AeTB6hhIV2+VYEDdfYseIbu
l5UdqcUxeW8MBfdBndob4pOEsQ6uYVi5m3j5C+LwImlCBRkAQzA1gwYY0CgyZ9kZ401d/n8EgRfX
MzBfyaDkLzRpPn0CA6/xcSyrB4xk4YolXzs+UPoO0L8iGY4ucfFLdXR0kIucistUYDM8ZABq1KJD
bW90kpIAr403XBXLWvTvDj0EUh6pqy7ynEbsD99HaFZHwUz7MBVDijoSrU79HZ/QYl2bcZSdtUiz
BeCs168lEN/8cgvUSEHPLxNxNlmeubBNBlzYoc5fT7513r5RuGrETu7sRu1OgCPvLxcOjKYTiiml
9DaEo8eHhjTErdy5IKAWzrxZZAivEjna0CmpapzoZfQGzpNKp4KfkyGw4X6UGrVdlvVLg5DDAaTL
FBsCrtzgk88cVf8KoQyta2wqNU4f8+RWTA0J/v/f99+NFAK1Rer7q4iFFLmGMBEFFlxJsGH8x+U7
ycLxOneCR9G4Zpm5wsQYqFQigqA/HQrdQniL58eEaOH1UcgHWqBJ1FImSfBeUrxQx7VBXvV8m6q/
WukFJMCoYzyl0GSDrESHww2uXGQ3fksqiim8daSa4HXlcLjEu4JEPET1OzCMzCHRSkgdyEN+lUan
wtXPXpjqWjmO9L+P0U8Q/dIcbEqeKOubvLP4EBuCSRzKIjohYSvwYKN812VblB9fRWtuFFmq86fz
w0xRVwiQMJTEEdeNg91CsFdP+njV03pHWuTB3dpA6lyP259Dl78ZWfR9oey3pkMrLt4rTIZ18Xmz
Qd+Lrx7bLMBAPfnB59AieCEdxWLbBlkq3nkGkacNhBu+bjzIDx1+eSlZ1NYuBt1TqFzEJhwOIlhh
rJNChEGK281myk+rDCjzXDIrFuqm6EmD4UA3LRqZoJ4rvcnLss0ZzGQI78Ay68rLgdJbDIPbCOu6
ByJpwmtI3FqC6FwoIoGkLO7v8lLXaSalXHjHSZr+HCrU3Uyhc+5k0iXOcxEPZGgQdvQRVJtapfh+
JL6MCgaAYFJ8q6RbYV+Y15VFvwU20e9K/TIiA4SfkEdySAOvqfYGQXnhRAclUGvMnjA6WbvBqZNK
NvdnxS5omv1VlhkSRrqkrNpjU0twrJTeFKzAW2Uy4CpfEfQcMgPWyuoLkTvsB9kvA50ld0VBb1Qr
63GPp2kBGWOvdzEps+2xmJ6k2Ge82IXJRw/omG4wizCC5XxLxCkV+3oihQOUG7bTyow3ZUFNOxZT
yh9HGX9pZfzNOy7piIsnm1MzaUsejolZOQ+0RReYu7cCocjatirz/vEQGqUEWdE/jz3ZSe3mKGm9
5c+5uZd/rHLb58BE5aq3iT3Lrp0NJCYcDgdgRuk9p5cElm75zsIxrLw38G7Q4OnlkPVlwXiMPXjS
CdSQiDBi5+Zw640Nzpv0+J1bN6MzCVujzEcjWs/lsfoG8G8vT/dg8Fqc+m3j3YPmYDqMFzTK5d9w
Mbh1Yoor6N2LUlMT2gcaBnyTVMzCFigNHGlrPthQaAa/d+eMLrSJq8WITFqueg8xTzDb+6lfanqm
pvBuMg7m5sQ+rq3bMwiFDsbI2c3jneX4DUfi6HHwEVvJg6ft7rJmmM8ZoyXp7nKT6Ygy9FC9ku0l
In5X7D+Nz1x15qog0q8/iM4gGRdD/XhpU5kDmR8H1d+nQmnEadMqn3yQw2Wf0xQVIbSV3SdHRML6
WN0IYaDeCP7BLRMabvDPugrfjdJXaEi/CIgc1AK/ynwpyHeoEkIoI2PoWIimWpWU24AlByc84v0b
kycN/vN0Ole+Q95sv1wB16oGbZ1vi5Pg6OBNDmrLj1AjZq1nh79D/4Fs3/4zWZQ0ayeJ4T7WYrFa
yNeddnCv+jl0rjnX3z1XVQ0+Yk/pSbmbtAYrAHqK+lQ2x4qv63hlBBwu3ABFJt5b4aYDQfEZ3q6/
c27oOa3v4C8QyjpW6AlxvyYUAIUr0Le9+RSXozar764GQ0UZWvMyDvPmup4OE2MNtHKE1ZDBRx24
mSdGHOfoBmHqgNoRb/URLlAygdHmHMOe3W8sDenEeo/Kl/Yi+wBWu2S7Eyvmr2BDrmCU6eqYA2W7
mmkJ6i1wF+EKbjgekVHOOFz+I6IVhSjo2uFo4rQD1xluaz9s68C0LnDwzQeSKdXg2XCVfgdUfqBj
GSK48W0FPe8awTKzD4lxBe4LU4hmv/vms1Evf8oDt07FqOQE4ETe1haKg5eeuEEZmICzH3O5b3i4
7tpTjjycsRfe1cy+rIBbizNNNAYBaBwmqyN9+7wCvRUIfpsHTnTNTQqox221a/GId3IhKOIeD1uw
nKNnDBDkWrQ0p6n45czSaj2ANb2fXERisrdm9o1ugaiPOGLUSb4FPZy8wAiC9eMxWpsAOp4GaD2b
7B+n4ZiJDBM2vyvm2IECAXMf9HDFgjJUI81e0fbgTVvZRXUtmXVq7+yPOzRU7Y1cH54fpsRRd+op
R6lvc1JY9P9V1ha0XoCfWpbOF0JJ5dmpmDX2qMvDDv8riGMUWxhXieUtyCwmRqcSeeqpg6fF9Ls9
mQ2YmsR3lANqGHH5h6kkXuTiA9P2kXyL7eWMh0k01Q98Ia99GDb/zuJjHh97/ZyheDkeUiuwetoc
/q0agSBLZO2PuBn4qzHq3xlAfnKnXMvgpJrweR9OHuRejqclAV3FXUF1wsgMtLB+TBZYSsuJO8qO
PSAAsWmNw8+LwPVlesgnUZd19jRz8RwlHVKgkTU+TPn/oSzt8EcGm3kO6qof4nger5Wl/sLEW+z/
yx1yf4jOx0PrGm0xXfBs9Nmn2om3ExrAIw0I9XLOTbgKCAxFLWgedUFu8vff/YjaJwY+XJikF8jt
xCO6nyjMc7N/BFT6aTim+AgSkTI5njFsyhj1AebDLReVucz5mOLsmta5pkgBPPOsYtmtv6XpuHed
xDT28Fgj35T3TTkIF9fmhvmuIeeJEk3gwi489q3znrcjxTwQdWD5mKIgVYJV37CUpZgw43g2TFsm
Am/qmbNoVoNkL3zWldzvAEoGqKd6+VA8ta4SU4h+t0JcZH6IuGj79YCkSeVlXX2heFlpw5wU9s0t
aCMyd+bO8C9vAKRKMRRJ427+lCmV3c6ael3MD7le2WDLkmmBebIqxD41JdOhZrFvRxo3hv3IQENR
fqjoI3EREC9m8ONkO1ZRLuoRH3CMjmc9XwcL4qoewXGKjwKERX/leLs8XvpsyNOO4VHnAhC2/CT0
fRQNtSi86cD+vIcgXWogdxgzYdaFnpp/Zr/OybNdT+s0Mk90JcGR6ivif/8oDGfapUNMg/F4zkD2
+9QBpmjkwmOilL6jPUT9lIIW8kcRrtAjJgiwf4OIBZC62zp5T7c4RTMB/wE1srhYixqGqj76nT6l
5NI6iuqEsd2an44qSbhpuGR7cQ9rEkrpfaG0ABMqXEJELK2TB0q4/K/G+OKPKvJ5pLA8epFEcwES
7Z9TJiOSALOoDj33Y8lV7WFFRvGzjH9JjkUWacJpCbzLxibQSxJ37Q3yUTktZx5NJ9JPgA4j4Npu
UyuQ1DFb05y5UZvoY2qnaFPoM4xXR/ixi8BDRNaP2i1MEzl/cC98dMHgPBqnnoly54/wX0dV8VGc
BULoBJg8iPCie4g+qlbxPdUD6mpxNE8AJuMDqpwUwn7Rp1cfU0kq+9Om0KtGcJ3kjER0dckgEopX
ccUky/hRQ63zy/ZypVm7yD3T2BnDQ+dvlTRYykNOCd5rELBhQttnWjzsMRa4fFzOOzlcOGG7bT36
8Ym9JH7XnRPVNUfsNQOUkCwyzcwgpj0oyHIVjL0jkBdZLqXgcBGLl9Idtg2N1Vc0kpX3R5JtIxE/
CB560cf6dO9nG9vojfbD0jC9YSrP7VrznjKMkEzJZye8UBU6C2Mf+mj1tt5fAZbMTKz21DbsjYAu
Oqq1sliQYEnPCnKdbNQAcgLMIPNTkkFvszBz6kByWdDK4JKC793HApLaPOmoWAEUTQHWt5JGKaO7
DwOpkCUl3GC4gBTC4LiqFF0Mg+UNA3lWnsCSvbQb4awVGTJlwBuQQ7JHP9g0+Pgsx7vX6Ewb0IRw
UKodGSK6pko4cWpL9s53FvGPrW5u59PLz27P6FEAkYb3HjzsgS5fEs478oLkFjVkqMyh8zsX1ZiJ
4FOnCsTGEw1oBLFE3oLXm3C5qBBXo9pHX7RVTzpJ1y+BMXnTj/x9KGGCsqJuwGMV5bcjcPGi9+ca
XNQdyFesXh40x+ZpgmgoD+qtIiZKsN/G7w7ZrpQFHybs+BYLZ7jZLItrkAY6IhGUeQDk3PqGzlNb
ghaom3pSyeImIMH9W3Rofnw4bOqsG0SGo7IIGpZYpka1Y/gmw3OArXhRR21bklQSxbSrsPshLN0F
8GrX1fIsgX/3ty7seZ59Gij6Wy4t51DF5wqjsb4pbpQ6kAMQnptap8l4HXIFwdq3/CY66NybJBW7
m1tDe0wJMPO1cYP052rn+KPkuUhu2LRxoqRc9Tz/d9lebf+kk6rww0FEWsgvFDNiem54xQWdSBMq
u2LkKRkL9K+x5+Xt5DUAsLLAyvsOKKv+tjOcLaGV6KVPf8rkTE+oKkWLgs0GZ+jd8Zf1+NnINBEs
jaTmsslS36sjaHg837pcxYtBFdMId8WnqWAhJLBFgSUkR+e2hy/rB2O9JSmBXRHK+rJNgYf3NH5A
VQy9Bragi3mQG94IepUPeeblikh1en5NR9HVOTL+zMHQo4u56g/yarX9MYYOtQAR89rK5ADWQ/nV
BOw6/ZaSvJgFk5gQrmU6rk1fTA8Xww5wSKjyUocflxKJ6Pi3PLPckB2CIBpQt6w+exd1z3Zj9g/q
RKGOuYKU4qvCBK/J4qJYbwPdXTZC86olbImupVZ9h5HlzwG4FTmCQCSFPlezH0D7B4QJD3I6c667
IQRrMVYq04cO4f/dDsB3ylkAyBa4fh2QwXC1YCGWlOBj6uAkLjLCgRlbGTnjQHnVPdzkE6afFwOm
yllrXZfMSdqX5ALsEb4/bKyipWOBxChjbK+P13pCyEb7xq34ulRDYZZ4P41IOKBMmkvXDuaD0jDO
m5YWSHsGiDNByGwhwKaX0CKqMJNX6ULVSRTulHAqiyl8f6MCCwlSvMSEOqDKeC5HQQZGdf0Y9IG5
H6tw7wIF4M1jJ5xJskUh0Ug8ozcM1a0qXvey3P0FgOeIAaMXaABE/YhuiXITzTkNfYSaqXcd3e7e
8lQ2H/A3FT1ceDnmkgJravvATLLdy+RzeBYm9oWW92ScrILxaJN+yzkmMLdrp7BJ3Mpy/TJkvfvZ
avDBHEJwH2iUOVSknrgO4WQQEs7FHQ+dkC/Hwjm46E4pUuO7i5NDnK4npFwOarE7S/XjrHMzK2Yh
Bpy28X3kOD07hawbvQrFotmsqaPvsXv63OoohQCosWtSbw0YCiR6D/ptcBbJ3AsFIF0NtY69aRoA
33jmOnmTGY484kyQuyahg3oyFxVE67b1D+InawFiqd+gdA1uaB9dtGOj1c9mf2n+WPAJsQOd1nLC
ApBhH4n3sMkok+rCHYirejv5W7UJof59hGjaOhjArhfbLGfHW3I6xY9QOaobtByLJC6VkAO+0aXs
SiSug+jbw+H28fg9+RThyu2yi5pW847C9BFbSedOksfCZuqywtQnVcf2Tv6VLmeaFzuUa+MB1rSL
9TbX442K3h15ZBB4I1XS8IcDpqeHMU+0qtlJ5O+wzCSpCPEDM96S7zmDGa4DTFGWBxNezi0/aXQQ
lZFL9SGOoGay3DV6SgmITUJMRlWFtCh7bA5mbJG9DxYLaCH+er4Ebe5g5lK/nAr10ECID8S0+9N8
DNQ63g5NySEZ3y6wpaab1FsnCcrOpyrhnzcYIwiP0QzN/IvLWI7E3jnX556q9WzRWBwa+Pl5DPXh
gmpY24k3fXrx54ky4gNdl6PbxCwui8qkUJt+Sf2vqsjw/BgQh9YSn4nrDWMksMmf4KE0LY5too0B
4zuJh+W0Y0UrSiJrrxEj09cd+eaX4z6TWdtMlwFZgsaBGDE1knEcxqmDkvMmoSvfz4avSznQaLd/
SRNfkXpgutDvr+BedYrM8jgpsKJvmDF1DNtts7qL4xV4h6+nq8wotStiPmi5T7/1xo2nlfQOq9YE
H04v566eW14Z790eCOdrY/6T6fek63L5wEnmHP9e0mFgc5icn0aKYGq2Vdb3mdrjXVmaM4IeMu1O
sOGWNMXan2i02MP5uC0dn5GYLtQtEyxaTnddt7kXbOnFPa3UAiNS+xV808EcaFlRz70PdiHV8PzU
MTa/egpDzwuqI8Zw8NeVJsteIb/h97MRaE5XUxWJKKqyQXMNam0rtt+SOgPG309DBAxKUxyZkGCz
/LciSaTLy9Ni8e0ro8tU3dSkbLRwSrkEaNwHpfXMe98BIY5CWKkDTayEfrAyRrVqjbfYBWuGmt3s
zw9glEl4D5dr7z+EZJNcGta2txywXCkeM4EWkC2issrR8LirbplwcGtQf6x4qgvZu00AgfZds4mZ
AzDdmKOLuS/AAXtLxghi0N50ZW++1jzw+eNgHI3CTbm078iMLUvPEW7H2U5Kuz9Ws/ncuBDemSbt
UEmumGVnPf/e0XhYsXRTVjZ1nRPz+6Cf9TvUWb8zqOB38AAf5QPuyIo7wuy/EaYUPz0YgZoGAygl
NHDLOLLY1M/b/vjrJy4NTHJDkvo0LkVbqssCLp1MDneSHgznhZvCZxZ/Btg+ocAfzbDc221KnvQs
6Re85ywYG6UE8Y8W/eCsZiDYqmlIFfIRU//v/PgKpVVd5Txd088q4i7zJlpDppMR593S4jxQ38on
ejbxIg9Cta9BK4/M1i+q0qQUMZGtXl9xm2HnpkpEzZksZx8qYcJHp1TTZEQ+uuePn6yhWToPmeYl
844cSiTGcE6L2PAdMRNq60EgvEoWDc7ChZ7LNvXDjH9qSsGfTdKr2FgXel6VmAE/1WuCd8o0utyO
igRFDpLtIePd/6N2p7Ude5LHkR2jp5xaXuWLvOJ4EppC8HlyBRah3ggOwUyiAuC/0ww1rDlDiLEY
JBoiX3bMxEn2uvvnx6WuXIONxZ0ZHkI9gnCJ21dkJFrV+YQYM18Q/DY5Hix6fvGL6qx+0I32lot+
mqjntdW0W7EziEsbfbTw0wCw6SmuoZtII9/9XnXjv9dFuuXgaAUXs9si/aV5uM4kLvkJKXexkESs
h4Qdr+gdiLS+VD60VKL5qNEmu+IHqtiIf5wtHH3iyT7IB45FzRHdtsG7/vzrEFNBUu6WvJesq8ee
k1pvcG3RE85pTUAih87VFD9J1o1KcSaYlmCsR8Rj5S3n7rYtW7A3KGFhfuxWB1Lm676U/Q2erXZB
LNJSP5y7mFYTnejwCzqkD2Yz6VpEWbXC4WxYojGPie6oso5DIAv53OyKbtBNLegIwQrkXKcu9Zd1
OYiMauBReJeslyF+8nGAjZ8JZp/9vWJi4w1RHQDzMdI80wHLmwX3TXioOn/SG0nJkyEto/VanjzJ
tLCwarCc3alcShp5ZszquiuGjSGwYvbdLP2ijBQ1izsy9XM+yelz7jTojrBjtiexzsr48ZLz6Uq5
z4bk/EQhsx64/lw116KCMDejObfiQ5/bJA/kz1L0xkkOWpqkWkGPtAD/Rzci4PVdO9QjxItNfwF7
y09jIUjZNsLf0dOe6aQdff0XwyyR7ay2Mx5KjBbT7Gbi1GOa77McRkOAhtLIpp2zC4FYo5Rw2Q9q
mKRVZjb6YRHTNhDPAVk14G2gZqlGFgIjmpspTmFM1eJpptVI3sI2RSyLn/wOwXLp5HsUtC6eeuVR
GsXkztwuCCASZ7POI8cvimAMXe4ptRmzkufn5XWU0AsJqnmOyVaq8w6toIQgwU5YgccBj1FmEVpd
TWKV+NtY/UKRTVLfErX5lu6GyADSrK3U58uW/x8PMvmn3labAkeYlImO6WP9iiUDQ3Dlb/Vax1m7
cqU9UoiWNgH3TRfuwzSTJXLO6L5jjqNcfFmO/K4q2ei6vWFtaCJyob/9UbCIZcEgLAT/XF3k4Qqw
mOuumvpMrHlE8IuRRkbnkRHtxVvfxe/iFWACmDC4tY2O42s1FAPSWXwyvEUfAvEB3L7jAK83CwQR
WPVPAbxtA7F6rHKkS5LwJbLXVn3DowmkO1hYJefW5Hf8OxbPwt4csLAFIqyLljfQTMmmD2m1dh1s
j205HfShJS0qIIxy5AaVkdD5Q3LvbGjcOcdId01wGlzjRG0DXk67uwVetv8EruOcLFzfdLOnJS7q
KJIHeXUD31pYGrR5S2CfZHBbI5tKC6virMLWjSBheact1YYvwcyYeknLpaPoizA+tXszMfY8ZBGA
lqrHGGGij4h4ynCjO8ZoulgEc5XTv8O0aSDEMzfNLRHND9ubakwiKfogBDGdDPSzvK7sFq/vX86l
j7FRkObDwGJ16bMRYdxxUH0sZLWUhfNFcailfgOCJTxUURVh8WrHbcBUdokS0yCiHpwDSZWDRTKW
mTf0q+5ce35DuMspMXswaNiVI28d6qF/o0RLUmFSXWw1jMTmCodxVYRl5jEYv/6QFzqi3cnS2kmc
9yDYEulDut64S0IqIwlWLnW7A4QI9FJr8O5baACgurtoKClp3oz57/Q6wZCyqS32NeNgo3J6Bt40
pMggh+N9rE3bNBCUdbrLL82AJYuCKYUzoiykCKIthvKGp+e16qTNccVFKi42xgeQhuMBJhPzpvT+
bzJVZAGdGsSuFFYaL56s27cxTIg2PPE7x1uwyma0tOtc0KFGu/VSHxx+g8CsOtqeAn7eto+nkfeZ
0UZa8wFsb6fGHht5vIJFHy1DfY0jsTLajgZp6yDfUweqU4uuaGRg7vxugUKOUVD9QKy7wrwhgCNV
6N+LAX1EHck+Qq3Nlq09keuR0TNjQLrJtd+myLs/Bk8odAP1otZzP5MJDH51jLutzzb8Pou4VjgK
FJJsv7GU56eBDwSVbByDeFFkcKBnjx4cwgmlkDdIDhERqzhPZWLGPymSPdkPB1hUgbjn8iLNO1WR
+8ipiL86E60abDfpNjFlFeB//xhNBg0WuxbmN9PkGWfh7ipMBbrbUkKy3xyOGxpURLwDl3DiDEvH
Fd4UOpjvkW7rWrvz2YxoT/aLIi6dcE41WXloS1sy/ldbaFLkZZ5AmJN0SBfDEqnf8kPOcMPQkGg1
aFLMACGpJqJkKDZbFFZ0qpTYyYxXOets0TaofmToa2piNu9BhTvZq8UcT7FHgsK1oGTeLLth5+GW
+xcUo839wjGIGvXb0uIC0UkN5cQgj5jDeBy9QiYOKGRJ4FZ0FuSos3J0Yp4E9OG3rmznfwBTF8e9
tie4OiY+lh8MpnOyTh4G2cStKhGu8y2Eqne+DZF7VjKc0X3vSYrlsAE8Zu0v0iI1t5S6JlUUfnvN
QLmz39SajCCNIcun8shNRjtvZXZSoPX+PacjhRlJrQl3TZcZYzanYA86LGkvJTD4Ek2cIhc2Po77
wchQzwvSNFV08AWyZsB0ZQf3IrUwvU9p6qGzoyGJzcvzwsRwCixhLNyNDl1afNA0M9tIOlt9LqTI
n0X1QBmV7CeHndlGTirWWw/JN4Lb4bHDPMpo7jPdXiq8g4VOAsLpcfGyVl5I6f+NtQ1MARLFNPvT
mbkB18LclIcWoTgGmPNoFrqKt4HpxKHaOZRBQTbiOXNVMempWv9nXD664C1LEbdGr0zGpmZVj63Q
UpdWBwu3yEXCGdBXSBcQu9OeT5qaq5CCON/b7CwSBmetC0JJqfWy5KaCN949JGyWpJGNZn+yY1Xs
ev32vkRHnPmCa5XgmJpNwZCyB7Q+LVKQxgrvYZYHI2PPw77C0H/UVLJFW6unj2ZNxHT+FHMwEoE6
m0RWkNC+CraQJ+enMxCDCaTSoeZauZ+Z1NyVjFVHsrqnL46itRfb84HoxiwSlR7sd2PZIpSFYKMR
U4UBHySreFcsFT81y5RrP84Ih1YrMGacRDhTmyDyNSq+0AzYHOguugt5J188s+vMxx9J49hJroEH
4rh5s2KA5fZHvI5T60t7Zm9OmuJE4Wgwxj26CJaXyedenZ8hnHdYXrMJVvehJljw0ds8bjrrYQHB
Phl9N/UHnnGL4/S6FZucn8DkT1i3kvApHXJZT0qFk64lcYaZN62cD8Fd5RYCuDEXJjqiZ3GwRrto
73fnRY00HQt7ukCVgy35vjh2Vbff7Ceo448JMefph91wTNTS7JNAnNkPr+6MhWsGLQHBmIrQv2j+
WQiqAPuXkfOb8fD0ijC5o5UsvClQW3WMptnt/+NcRCBls8ZzEohAgP82qf0dwgzmfg+A3f1X2ddv
vYMwxil1luPHxwryVr7ftTnYAvrjHekj082zAePug75DUDvBtdu6tss+wwOjhk9OrPrRMe26W536
gtLt6bwv5Nc8+bUw/DvDfvzAV9uBntKwB+Agv7g1aMiH9ucamnWgcmHBVuLPSNRMvu7gQY+yIaJN
imhy6L0clHU0F+JC1P0mgckkGKXVFAk8fn2v4+Ug79c+vxwAhjKZNJAFBEYqCOqZuP1jjn0PdU6O
/QQ8aWzsaC7SHPCXMCv7J8PwP6ZHfo8QIaoa/izcG4tjshK5Te708ncpnTHsKPCnhtQl14kwyiSW
u+e7WMP1fIb7FuitTm1YgZBNn08f8eD78KVgyBeTccnV5fFfZvHJlmu+25MgcCyAM74bQDFQJYj8
ZnrWT1R+ZIe4sjaCdLFu/awyNUn2b1Nbta3a0wSEGBwg9x4rymq0MOlmhR/wo5HBVPBGoQmnEAND
B3Y52O7Nmy9+scXaTQOrXcJzTK5pob4HipIxf2iUyIkdYtxAXTkEOAGsueNLcGyxj8NP3VaB70tP
RPzo+99qLVNGeIfkCI4XI4q5gvFcMCyr8Wm2pU8fkzbhqAoy6cWAgX+CIdsD/tt39hF+7o+yPReB
kY7RVFlSGhqxzEF/PydbNBELrzDGKZUGju15NKJnqZeQgZDMzJmdyXjikX1MPaHpgYf8r3b5xTe7
Mq0ZnZetuOD7LcvgQvaUaIDhqBLfUOktV7NCadajGASuTDKTlJI0LKebwpI5cCMd2N4/iqtLNEBC
FHLwEfXH/M1NpqAP/ozqN0nZ8uh68Xh10m/HSAe/kzlQhuJrr4EqZUZ9SE0jMYyvGFGTmG/UMt3p
hTinZkW9g0dT2DchpQ9OVNLbjLSYVyq//Q0Y08RvEttP/FgteZHKcXIkgdG6uxd3LxWuNAGW6y6n
SQKac8xL7mFcqGayelUamWpT9kE3NWuPJ1GJXedZ7gb1HJONceueoTRR2BhOT7aY+BnN/PQIfjlL
5GG+iF1O7dCNx/UhcWXoA34jEkc1a/DE1LW2o1097W0IzTBZuaTQAlN23aMbw8GKopVF4ZbRlVxk
PfAyuD1W8Pkyp1a2KADwn57DDtsom672VgzLpFLVWrKlXBscLLGS9RNxirhokY67OndXogEmdV6C
Sy49GsWGHcneMwVP+q1oMpPtUd2DoZER8A+d5EzCFNkHg4uDBt/Y13iRihrs15X4Y5UOK9V3rRMd
OVwSP4E8zkz8Bm5k5DTYKZ+nILGePdEbmPGviXVBrzg8TQG8+38xYdj0hMJGXfmxJxE4nVcLS+/l
+SES0ycgIMhBWE0fhVMGd/cHJgeA8bWYsVGSLlR9ZUBBbZAPnmO/2BBXH8sFp4wA/S1e35AKJR5/
kOodeJalUKxRpesqakxtMFRd5+IpSEePY2qwZCebs7lGphazVNrzxyP+ymV/yulKV+8fIu4XPqJV
5BJMkT1fDaCh1QWpZbZPSnzbnej3BJsjujRFvVvCc/SaoKjv64GI91s1EnvrcCHIye3eE56aowdk
5pBuIJs0MKeTZa1bkmmVluqf212dUC0axbrHNRH6XP9Ckw59GuMJp+ROFoeOnhgL2q/PSqn7VhHB
nG2y4pMCswEtZOFqiTkXSdn+xRmmLQu/eFw2jHI6rCIIad4jyCfVlaJVtU6VKrCl8Brz93V8jzAT
RlNoXKgbgxmlLhKsY7NuCAptbOjYNqa5iS+mufZxXg+45zVdouoXjhTmtZ4VwEr10boznIR0R759
TczggNBybGqDFThz1Pm33kQJFraL7WAax59u2JNQJL/j7y1YMBNULBKyFru7kbMnufJ8z42eDXo0
4JPxSIV2EQbeBgJwBKVZ1tQRvs5K1gq0rYkTBfs5qkejWrg4htsCGCnlvvsn/zTkAUd0+8BCrtY5
q3dYPB6RrsVzSUcgCYd5cJacCTXkzAFn/tdRIPEtJExBgC/AKuAWhfi6ZOqi+I4DAfROMbXMIUIc
nOad5SwxK/cLZopbfFdS93boT6GQFosH8H4TGI66xDJ4PHPBcVDhqfyIt/uSg3PADIe9PfxuNgdt
hdMFQX5iSqYYawesCq2wvREa8+Y0zTvu78R8sNhPN+cbzxe6SYvP45ExEy+tzRLZiwaWXrKX/TeC
kDAMuIaOH2g92W/6CQWFHEx8db4kYBtyTjGwkGhHMtdDz53s32T6yFhTDwqnF8ssg8YNmzcCpNmv
reETzwj/WmDses4Vm+V0c+7+1ruKkW988JbLMtkrMvA7M8hnfy+qn7DnWe6B5pFWkneghFOF1dd7
y7kg//AZVBVZfRhAjCfNID8EBa4epxSaAp1j7uHXoggyvpF1Oxk6QWSloGFJIfuwYHnjXONcrnjn
hPo2xYuzjtL4UK4mm3uS/5Y3mslseoO/h8Re4QUyk9AaTyB/0S4/AJsNrKWj3KTT2G0gG4b+eQED
LmBthzBXeohdceykKHCcqDHB+eYtlSYueGrUTA/d1HqPJrv1M0swiLmSFjtRNRHgFAe+QxBnBR0i
vCQ+Re7Bo6ua0GJUTCVwFseeXT9FohdaDnyJJj0uaHQhNCjS+ZfuyBAM1apB4RFjkk8kEKBefH1Q
cQEAIduvxw1ve7THm8UfpVX4pSznCM+cRqXhdsOtYsEhrbmKixxAEMCVG2RdGN7NmzZZnLr17pSf
tdieqPqWpmPjLZpz0iqqDgPGJIdLWgeFhP6Kf2cmOOyRYoMNwnpSvAsNxcE+tgMcFm0dYEUR7DxW
oXQVjFjpDSfGeV98dTky77HLGobLk6w2e8M1V5oK/hlmY1iRF/k3tyMIgCmzFRQLXaHYlZPvbx5H
nf+1vMvVZUcr3sI//kVBcA9hzuLT58NfJBe0XucVBjAxd+kONaoq2MrHMgPQlMYazYkCJKruV6eb
8NLjvqZFW8CJncwywhaEwzNxMoTBywmaKJSCuv5vUl1t0KxkT9542IcxqSs/1dnrFg9aJujc7UoK
2bRB7LE1OEl4sooWwAxt2qCVxVWyrALcw8mT5KMBDj0FR1F0SJJkyBMcl2fNcFUvTSEEkZok5Qt7
yPKQlErn9ckx5qYS/wr0vs/k1j/SJTu/nKfW+ohcMlZTqwD/jB/bvelgFGo091OtH7/QUefNEqz8
4tYSJiFHaHs2FMMvA1wu3NY+rYnz1U+IXINzQUZg4ZJlyBY8t3gQIwaRIWcEoP1rwJaN6ZX6WqFQ
A+2mQFmfdrzA4uFeNrDuhmvb2KSlWoGyMYLNsdBt7bsN3xQd1re5hcro9/QKrZMrpGe8D6gRq2TV
gaVZqoWH6gk7U8BujffJSGXL10ql4MMEhP6lKCGu2qn2CBTMY5fpiA8ubMxHoCytVVKjvSxVL2x/
PySsvsGoCPqQsI5MOD/Z23ujvwF/dFZxw4Be+vFh7JIWb5j6jJ14aoVI8OcLnrA+9izGG7NQfjfq
8v5bO2fS44bD6KpsWeWHjI8DETtChNIvq5qKVVSKd2NcOd8fryheTpBVUK7+rwKKzmfj+CQf/iZl
Hwshjn0NsBBBsc97d0cYdt/Uzm5q7fiivQa+efPLryhefOw/eIFEe9gqipE2ya9sYgP4jpRnq/NK
nRLM2wYSLi1hdVWtz4GN6jFZfhgnQPzwhFRG+uazZoxOBKEzp0qerWlTTfn6WudqWcT6eTHJXCRB
KO1gVZk+vre0CsVX5J76t80snP0Sf7mDBEdN66RZCrB+Nb1RD0vxjvPi13gCuLrtkemQSeDWseni
UfboqB8luPvTjSPM6pPoVEIlhws9Xij9j+osCV9LJ75aSK9yXEuQQzIc/XHzqyZcz0KAMwpmWxTi
72NtyBMfpr4I3wwZIdsDvJV1wpm4v4bpgKamkiPpi1CO5usRVK5HFrZ3spDss2rQ6LUKtCK7Bi2S
Taw8y8hbg6qzlKQTRvz+Jdz0HIBSAPJONSpHkjWqooFL0xjnxvKPVHoOqjasL6PfDX4hbIvpFGpZ
CvKzxfcPbWQSwo029LHE78xca0zy9oVwuhPPOFCDaIGQdwQQYn6q7CI0A9QqnyQHcSFhTL118BKq
bnpAQ/paZgzCxjTcW1PJc7ClUgRyTysxkAl/891AKyoWswZp7mWUbZ85KobEAhTJVI66SUY39fW2
darRogDij0MMH3d23xbb12bDwQg0pbq+9KQpNB+ZGW/mD66qZAL98ZrLbG98PPkHl+ENJFC3ScSk
UMkXMpfdejYhwX88h1pI/W22ewm4R+vPYpJ77ukrEaZzVLOO8BarB4KQ0nRdE0Xgs6fUN8wEPgW+
PKyRZCC3MTJXAHLiE+XDPSGtOC3aXjoREAXVF2FIpjSjSkpkQLBV+M9xcrAU7aQU6PJizbL71uXH
AW48vEk3lismM6BZ+RktIgqN9FPuW5qBekNAb7MbZQpU4J06y9OwZHl5aK8008m5zSVB57ly3suE
Vyz1F2HxhSsAcaDq17j24hgwRnNyIAYTY65LIENFbgYUiTtb9Os569qoYw4/rph1dHbT7jqh25WU
CGJT7WuilmuURXetNb3VkeQGBWNsJ8jULE5v0cZS6spyCw84AnzblB6r8vanl0xaIvY2OyPUyKJL
mesIqZvgp3oUvxdr7khu6CPIZYGJKsPN9zoGvUhOLvYU8pOc0B/nPxB62+NsOKjernVanN1gC+eb
wFHfvbW4URIGy6jYyrblPdOomAm0OMQAYBfogil4Q591tj0/fH+ndML74fEzkQwFtyfHTd47dhfx
Br4dseUm+zUcz7WYIW73yCPiUvKVnGDXjuGWyKk72+TTmfmqMPDsZjYPv04SqHOZ9uDTHO3HORYC
+adXillFDr6UL2T2b1KpHwmIjUYPOojck0VyHtwvrffB3ZPKuDEx3DlqtkY4+PGfRMiFFVOloPGT
vPofd/AcL00qCp2s5eeho4+mNcwIc8KWqC3GLKv5Cs0XByVj7YwQLnCxQKnu9GuJhKRy0cVeBzYY
IFrKUkxcDfmsKqS9rSm41hciCeD5s1GrV5B99h0NRELMK8XlT7VTUDICRH66zL6w1qd5m/rDpOD4
BvxFukEKsXfs1ZHmbX75e8Wxmt5sdFOHiOfonJxayTHXdAjZQaFb4GsE8UKEoVWHAlsayhiEBz4J
RhLNKo9GpJ08ysHwoxTkHgXZG26BfQuUeswlCpufCjEMDQ03KDXb+Ez9MAAwAYLPcLmxyObg/mw9
tYuz/HzSBva8KMrGfNwhCsgalOjiOvmw175r/n0Hxkc3XWIQeheErIJK+kuOqSzIBxPEbJnqzJtn
/ja1mLW4T1bXsVRo4dDTjIRhveQWuEGieiQ6CJdvsk/r8NPv6wfDk7MwwbPUT35EjtVyOAevMBTq
GaM5OTLwycQhiA3FyaepUCHcDTuw07nhD2Z6lVJNQL0ALWehSW15fG8GtO3U1N49cqAQeXsgE87C
g5DB67ZnpnuJ7kGPjfRSHjMO+s4HRsGNwE+83+0zkTrrrJSlrsRdGGC0kwxUVoMys/+yHOE/QUlj
kW8mXaDdXVklTFRHCoUiKtSVbEfafso5wOjy0vvt5CxArwYsgmiNoo4fLONpYSOy4SXS/6rlL4Vr
33w2NXb7NJM4Uj/wLMVTBujmPOLTzOAbe5cYjAHrIC+Zw13Je4X/PlNbwTbnASeQU77s9ujLlAnp
qctyDgw4dg4iEBs5MShvSXiLpjDVCImA6LmHG+y5DiXxOIzAJfBX6j0Fa+5VW+ng5Ho1cKufbZsh
dAiMNj0ww6Z6M5KPRlQS9Cy07jw5FEShKyHJpK05mxZCne4viRV8ndjrv2j9gh3fblZjtjybh8p6
mZRbnuV0x5KDvh/Emp3ZKFBGnc7kjRIaT0rRzu/ETEJxPg3TeljT7B2Wpv2EFcOH4UyEEKy4PIN2
Cz6ZqHPyN7nVy6sFflYoTHYl4s8GGItMO4omJpQ1MJTPYE2kLlk/LdbC31OwhiFCubXC89YcZIIJ
97k6AQSzDXpd5vF5x6qtYihdwB2WLyYLfHfxfI1PRI4RTQJNDSXtprmGJzd3hmkXG+HgnZgl2x/L
z/4U/jIeg93XYEcO7VQKFyhcECTc6Ua1PDCjpt0fCr9N8/CfMPtNcQ5u3ExHcbdij7d1Hh/bEWsJ
glukEERfi74GajK/hg/4UTNTxUmKmDhSR3SVaGsSRmeoQrHS7exQWcu16yvo9Dl2rIhN6t/bztRP
sptIb8BVIxGBO/qlpGyPOc8+SyweLSKo1Qig85YHxrQZUYSCYU+48vC0QsomjaMVe3SyqGnZ8iwW
hoHz4jlNNjZ7bJW1k63kTqw48BkJfpzswYINdYZYxl6OwXDgBg7XckkwwRFuTXYuP8jPKJmLFNhv
OCxwNO1R2HEwrIJyQulbJRbqIFv5uxa3eKZPCSQ2jTmi1ohiF0fpKY3drAh8Sli6JBjK6aLcB0bs
ckd1xj0WhMIrzSvB4TWKdajfVjAb0LTILocrbr6nGlEau1Jg2bRtuLaaNZwJtJUzwJ461GsLK5yt
5JOR1DJutD4iBioMOHNXJw2Pgy/lX28m8AFt4khMkDNiCRaJlxqwXk/PvWprtcwZ7VntJsmiGKSe
3he9fWMQRL639j3lF80vWo7X4FIgZFTjCsInD5OGU3r+MmvXbYPYGFC3V6aDHhbjVVVsg/UB5Ogs
tQCMvVU0kaabtBKRWzRxG4r6+aLFs9Dvq5bPUUvXU69+VBtyoh0uKnoKsi7Q6y+t1M8uPkVRju2L
6D+dAoM3lvpaZOWqZxjBO5gOLzJLNxw1V6MPk/y5QJ1ijOwwuOMcwDGS0wHPg4YW8YC1wl/IsVuS
saMsHvWvWMVLhJiohWcgb28ZtknnYc/lkxgDkEIzD/iiCH5oScfDzv/IovGS1nmCO+0Gp+iCX+uc
AwNxDtTXmFRkNUBJIzAGkN4ljvDASF7H6jHhv6aNQPg0Izy/J/dX/SHgelxCvXbsB8A6axgetMbr
SZU0GWTnasFnOru1m+DZuuj3pOndr/9GHdzEje8exX+AAJMW5r/zZFsaYRuGK+sQydYhImL+WD4g
hmfyxr5dqNHKJ9yRQvqZkM4OCySW/4c8uiD2Uqt4pAUlP4byj1BqQby5GbPEjEwKBcfody3q2raD
orQL79QowGh0wHJxZuwg7S79yZvrTD71bkcudR5PrbYVXRdzBuNEoTTYqD8sN8IMLWyw7eKPyGaN
Ka1xphfpYlNkcvA/ADGhb1kVJwTm2DOVTPFYKRqzPpv7WE9RlwdIcdKiK5TpRQKEyMC3yiWy52Uu
YuXZPCtNR6XrSpw0XZOQKovAqdnrWcS/Xye3Ow9w8n94L/GBreOOozDn66jx41nIOHjw2WhWa6eG
v+n6f0Qzi5d8LZhXuZUAPpjaylNZaKiEKUIGZLlVOd+dZMtGaFNOA4L35dTBirDNFbpnc7TGiXlm
OeDb3KPn05smM+KkIRsciP+truT5yPJBM0Rx+GGeSq866tH2vzxOU6GaMr/9GMEjhj/aWPzWFW2A
pzYMlnPpFh1+P7YsunpW8IrYVFjabgi22gWQHHgbWc80yQI00BERiTE7cihqKDaRCGtAApoKCd0H
bMsR3DWQglfkhLBYdbE2Vv4NYu7P6SWl9TZiu7G/hykEcUBtgaAo55i/bDsrV37R/3bW6DqEy+Bp
ziaGzL/vtpLSQy2gZFSGQDUKP7uIhjO0izoIqkRhL62XDp54AGrgg+gWcUnbNqBUS0jNGTgbFfH8
E3IVLfJELAeuMGFm7tj38OxRGdI8LDyhFusnWuFMzHHu5a+JaxxDxuoD4VNReO9rqlUQBzIGGDcC
xw5mkfoIIhWO3t8ElPlGI9A6ElaAENHvK1ULqoXmCcSnhkmfsc2/n3SwTflFDbYAi9lEubMYVUUJ
aQUV8f6PZqGTlRQApP8fiqpVXGhsYDRC5IXfJllPFUd+p4k69p52NyVzl6hKBDjPzLvzY82cBg9w
MYAasp7downSmASBW3qtXWMlN+oGNt5klQ/taU7RGOUFpHs9R3uHllWn7iiZCIk7crJ6Ni2rPwSp
TRkm0KbSkdF0RlZkXOG4ZWAiHfSInQgJJbbSF377VVJy6fbeB6oQktvOnfp3gP1f5eMMAMbApnNi
1rXkrAAbzaUbjwgWhjjvr6MPQlANuWaDjFCZx6ugO4+lZa1J+n/8n0tQ8pFnuUq2DdILijayLV5s
qJPQ/CaSv7v1CNwXoagN69ubybvg7755Gxx7jQ6SSX2Ghh5jYoisEim4gIbxf8kflAkW3Qewglm8
HskVJw3pyTus6XyxOTD4FmYb9Jb3vzcNRekj6UrlxGJMsztXq1L20oTb1yDUggA2xiIokinqoghi
0YNvrpQCZlhPS98C5L4s6IOgBVoBMA0+pCu4cf34sYda51WWAFMQn/R3j8cF+04xYx1fJ/qkdKU2
0deTzMgeqWmeoBqyByO/41zgkm8iliRfaRet0Xe6DihMRG2v5bo9+dFtQuzoijbVBnO+Xwojvr/V
+3fHGx4bJT161DAXYA7Tpp8QyEgcHG6e9XlBr7sOA5fSjY345HcSrcRmRvqEhHLZy7tQlsv7nf7a
Jx18DTCtjHEx6w9MZHmpGM+1VLCZPujJ5GFfZ1+aFJPLT8mcvxBe747K3HronZzDpiSdlaroxHrE
qV7grD2VuWCXodRzaOZEJZJbn++z51GmgHbBHUUES0LwYXSm57qw8xrpypF1SgnEgnwffgFY/F6y
AQ1lLolu2aUg+iOfJCFyIH2lzBGYm2XwYjlXH2NC+EIbHpHlPfRQoEJSEqDnRNPN7DsyIf2MmWB7
Z/6nlZnTH6bmOHndiyeJ/d3SyI6RYzLZUU+WuH0wDlNIJl8FV7/Kwj8S9tMOfQ04Jdt5DHYwdD/v
Xqh8QkatsKEpWMVZ6MCNH5PMFVsMDC3GMzUj1+TdnMX1o69Hgbb1uB5EEcGqRR6CUwlhH2ZPd7Ot
QYxz9pqgisI/dJGAyiU7qVpeUTXJCl6d+K4/Dp7FkNeMmt5Owc6i6i3LAlR6VunFK+8NsrFIuucN
u08IdIRALSpLD8s700meiSdoDmuM1RLbb4aT3g9Tff4K69LF8bpMnZ46Q087YJYJIEXa526dZw/B
xco14boU5jW/cYbn6nejYQtxEOf5T/GEACTT9p9pFLMTRfm0EcsWH/Y4nJp/FffZIkXFxNcQS9YK
8pbW359KL9CkeW4jaMLwLWBRHUr81FWbUAXtHVo4I+r2vzkBA4jOLa+hs3z6xLyef0O3N28/Br4h
iDoBs1vC/+7MchOhBXHNzW+ubKCknXWakxqXQx8pjNdpl0flpJ07HO+04oF/nStzf51wNNh3EF2O
RnrVF0k49Wh3C3XDCX0SjwCQgWHo+EpiKpXYuSTo05sOVGZXzw3jlC1gMSE9NvTG6nnwk+pHRkb9
VLc27H01906BDZ36eRTmS66Ry7hrxtQWp2F9KSRiMu0YDdRN6YGBf4Ld+n8yoOxh59VbyenaHW4F
7y7Lig6t8hcIXN/w0i1rkhTF+/GTe9EepCgzTz9KJeL0uuxCE6fCzL+BNbHBTFQEsp8jqyKr0BaN
a7BWGhBWNK2Zpta4hoLKNNNC627RwKg1qofp07pHtUdFj02dd7G9cX8Cn8koqkGURrot/ZqBP7st
531Z7CpoDe20l2BE2cPixQIXX+2x/TBKlivOahNwBISWASlL7juk37GzVK2hPnzUR3qbWuQVqbqJ
WhG1RBL8faocsBE61QZRyUWWKqTgv6EpKTKaBZmaKelz8cRXZZ4VdE0UIYJweFZRZpadJrmOaTXd
AwdPSTJMCU6V3gWWSWoPYZ201UaBqBaHF9Da2nIjbeDaFTyrAxLSBShg+2znzzaDcwaCuvAM9nuc
vyakDAoY3GVEKaAiMHkjotD0TTW77bG8hbJDAK6ag4dupFS84nmCFakqIx//Ke3bRcxl59eDNPFi
Rg1ZcyDlflFn6z1US5TxQo5Xnba4wxw/fzHL8jznXoCh7ssTrYCdGZtMtqeZbf/DNSJkKEIzhV5a
d5Sw3J/yZ0HhSOQ3PQG6UV/aPwmgjHVyxjDq+AIlKPRCEYsuRlNKgL15u4CODg6GEFKi77euSozP
TuTPxZgGs2XL2qqK9uZAf4qkl09Z61i1GjOn9lvoFmK20s7CBHBB9/htbawiMnqw98QDxTb8qiSu
PKEJMTquHACm01jkQEoxwV6Nl8Bm0HVAQLAFQky/QYV7XJFJw4WDyiABtwaDvSRrmw5fU7kxZ6XW
vjOBzdtl0AvhVLikJZt4wHfjulDth66UnTyA8tOlgEiUyASIj6V3VhotE8U16lIfmqiUFe90VA8d
99G5vBFKKFPgccSToDwgC2wpfAIzzlqpDD9hSnBLfIb4mmc1QWMHjLc55Cg+v2bWkzHB1Ph50Dvn
3PecId1QbMEIah/HlgQELXi66vqJGPDaUGpnv6kquDnohIpcQxTYZKKbb1rmBQhkXzlRau9Yggu+
32jU1VtKZ+R+/uyQKDX1axtnu2sPLEebNNQqeYura9LFA8NFXCth9KeXwMaWfwCVGv5vuQUor1gb
83R5PsnEuKYf0EyXFjCg5SakGUKbhSTqidUEmfzSo1CskEchYEC4dtYqLRfkLKzBF617mb6NyOS8
fn6tlruglKwrFJ9FYLkwQHvDwSH9vj4ts7l1qZhxzoPOEQo0a9Rz7UZ+I4uZtd6GF+6j0F7JK1rx
ny3YGQ802TJ0aeC7cX1wWglhW4Gv7xj/8kK0VRItgIzYFGCpNqOVjDZxTZ+38FvISvN7nBZFSurM
tpNKIovUUzvjSljw4wJJLh9SxtqNT5VNF8l4QZydah3qJhKqyQHppOfHWDdMVricB5NfDN4mrAnB
A//wEAO7xfLZwNbH6d9c9nr5STERnIQRXyT/Zpcl69QOZa20dFDT7KvIwV+3S8yISZaVAXnmw7Az
wAfcZEeY2Du0gpgMiXV0GHrfpjep/CLKkZ1UvWc7Jyk6xxVPfWXX8CGmIpd9tSV/HW61nFldvARm
4C2Peob8rrgZuJvH7ZwPICHkwSoqahPf94RfMJYFhgI6mnG+ZeUvInpXIVPcTWB4lXNHfRICBfYM
ViPRPdCMfy12qOd88Sc/BoejvlNHQajAwt025l08W48agk9A99UrKwIMdkN8+CTsECePrjkcBCrk
7VWnfht06dz9UuFcm/izjWU4oi4d3KVKmIxp5W45vtORqtpzs6sJYpvkgRaN1rEm7/Q0HGRPZLQY
a5BFflD9aWKqtpgfwrqfI6Hn0i9tniwsoqzSmZrdHwWcxCgQlpTlpETelO8+tEcsExPMmng4+Ux9
ZA7FumpkIPVn1asME+Yw7+FSI8EpPazOhwFXg5CMBUZRhJAf9pskZkol58G7goJl8R8JfZidEJ0G
cq+yecWPQeZpPNxg8Re0de54ZnDQrwTxNIn0VHK3/vaKZt6AjYugr4iu9OfSVLxAp2voxL02R3nb
sW7X/0wlwAaMXNuEeSFHJHcthx6JgOcjbUcF82KKmhiwFPqdXGxS3RsbuOL8sVw3jCWHD+i75Dn9
WNt/zHXEeq0ftYK0BuxWLGLP5sqGDrA+3caWf0SqwtZ9cRsC8wcs1ak7rCj5hzp8iV6uyJ6l/0g4
EdlSicgeMjFdvc5Wf1IU0N19TVybLypFdK+xeLX2RrsgS0H6TA8fWCz22YJmwni2QZx0yphwvB5P
lqyQbiJe1b9lgso+bkJXxXeF6rdGdXahttK5pXHQwXDCNqyFCy774JAfwg/W6nSnwe1MTU+JxZze
fadzIGeb+NaloG1dxcinfwHhUhieygnYjaRTO0TNKRyyh7Q/8YY7nXVlRSLtV2KZujWdxcymfsbk
tJAeRRo0q3MgPsZ1DCdnvntD1M6vzTHFh243szZKgJRYuW4PQYQz2HQRw7k0Rh7yCCfBEjPeZCbb
Ow1eLNuUE70ul6jkL6GwN+sCq5TbKxeyAYdRDM0JHxMD63V289r/I+74uwr850Cu1N4SYAd/gYPi
jOzhBRfTCTaKyL3+iJzluyheCRyzxunHXRRo6E0qmPokgl2o8YhfYBkRrx2qIga7yXnRVpvJleLG
9NZuYtr0l4L2B68L8HQQV8UdqadUSM3tPc8GzNmUGjPfZJ1AdjCQU7LiWe8XDzNylu/HEwj86usW
eNv47aj2Ggwav+Ru2zI6KQyqaT8DtWTf01J8lrCvND3MhKW5VtJXY7fKkrHuHAM3vOM0S31Saf1e
0k3og1Kz1LhLrcGzZAp76kWO+CuXC3TGUnmJ8Z42AVhcs2FF0f4aO2FNx0Ggfs8mXjQ5Jo5PwI6r
Sh9IjEVXbwCZ0jydTZEeeJNltdPkZ9Ekp+GYGRIjoPrwDKkvI8H8MZGUVfsYrdLlVSAYy8uFP9LP
tCZomsp93IQlYyya1tNVG5GKiZ7CPVGdKUFeNcDs9k9MKxlN5z+bovdZGJx97HMP4+fiOVzdH4/a
MO04SXbH3VUEf/n8vsGhlGjoDp9jeiBgIrP2axfF14830OmTxmxPjUfuJzarHM1TuR6/Xt6b3KB1
Q9fQCCa3rQNtsUrbtIld8QUSt6JjtFA2ehlZhtyUdwYPtqDqExkCDwiOzCAb7L0QpJPnYcmu346M
aGBjj539lTibyR8ds02CheCnDZKbZ2B1iL98jlQNx3F7VkpN70OAhgn8Lj4gWjEmsKzXslwcmBLF
6Zj6aQHktIAWbtMFKEFnjX9vINs3TLe9RTTGS9ot9Kqem8QjQGPlRu6nDhGEcyxYnT//ZVY2WsJI
OnQpMA0V8nqAbplk97KdDbBV3nsTWqLkkByaEi+PnmYayE7blX45BWoSMougSe8DhSXEA9ZTWL51
Fyt16TITIPJ2OcB+TTSmVM8a7xhVaqnTG2gokokK9b9KuAsR47WxBnmesAKonCQ0dpJAIDwrtMM2
gdZU1yZ+6VR7RY5vXxDL2shwT/NhKQz63vKPkyT7TGlaFPOvxrkNHq1orknhl30EpTAiMN8eD7CM
/dZ783TTzDF+ihuXfENgiQEDAvN9jdaeDXAAnSzUR1xJ6tF50iBtbltYwQWx8XHynpnJgin2B73C
d5/df1+JHAKQIFGfuVjLRTZMPMDogCDwejr8aiSs3yu4mXiFzjkZMJnA7oGTDHk2qzyR2nxB4TBt
3fxA6qSbPTuLwvwifxRSQnC09zBV0wqUpSQSbs6GJ22zCBmJAjp/3EVG+q3J/ULw7psugcYjpvlZ
4KkXxWR9bGN0TOMMIiyLqnvogTwEEnTqI0G3MqV9nAnGJl9JZLXue7uKjyzZiuaXD8i4+mmBNGDk
ie68/PmpN8u6BDaJIkvHWAJJD1la5zsz/twWwSlcfQ3DfKrEpNN6hK4xd4ZYShKlfQ8xtgUGCUOJ
ZZAzI71c1Kffhvq6a4B59pUXDcP56jEnp0K7HOJ4w2wxBeTGFDHhdY8Xx9W6FPnwPXmgm5/9a1bU
MKJ5k3BKuAbIK24AzUFO90yClgF6tzCZtIEzB4Z819rrhvrsnwXjT/Gw25eCIQQu9Dw3HR6qU/RE
6R2dSKMPJCzWn2i2eIkTwRccCWqOhvviZxzuzexfBZG4n6X33Iw3nEeKGy3WecTiSIHUGGrUXQxk
Ja0TYl5OjjyutFI8IVp87iUUZlwL4JRIPv/B8eOQcF7hk5TPocfyMVEO9ADLnywpTueOsL+Gs3Ow
q17+05BzfYdQ00VZLxRzYtpJ3QQVxQCb8c/cw4gjJQqgYfyrXzmwrhLBedWp+uOJPVyPazCrLAh7
5PtP16FxtbalbLQoFXq2lDcAcXkU0wcrA6v1CpY2GG5Ragf5BL07BxvSLzIDuZqn0Cxt8y/OAvj/
C9tmMqj7z+qdjXVPvLL3gagsHePRgdQkZL8RzrHBnbkpeVL2IXNMG809ekrDX41N73jHKEoJd0Ht
q+DUK3bpdVRtmDqR76VgTT93txXlM1RlAXew8hR3zAVIphS7a7lj/oe9vtf1ABjf2U7GQzivkcJB
oKVNPWG0Gwy52dd+WGN6TIvLzsfE6mCl74hSeAjjtLecRS9A/hFpMQkgvCi9OTqzwireuOQY2FrC
yaZTqrod+BihrgomeyRigvisKP818oNfQglJwijRrdsc9Tdil9fN2guHwFsNGDysVofrGoOotCiM
M9DZ16PXjRWygSuQ7Ycc8rRlb7rmqYHoEFBZN7mAD/TmSbdtZ0ChmFOTDzHU6pRSfnCBUyd0SC0j
sRvtdhQ5J4Lw0gxAKaew1KutZ2ZYjlx5tyBRAJpYJkOuLI0u8H8CpNK2v5WbN8o1Ur3cG7nVCtEA
AKO5X4IuHzPLfEyLATsKpUfLJqhYDHIAV3zvvnQQjoxpAJESGdBVGUzXvPfY5MUB5ESfO1bqk67P
ke5wfjE8SFxTS14Xada+/MX40NZfFXlbF0yOTqyh/RWp0wV/MiFAaL3ij2AAQ+9ipTgUQFzA6ZcX
gnvBUST4e0xu49bRJ/Q4OrpXtt9iaGy2VeZDpBqbyevD9p/3YuYS7TSwrZ6C8RQV68KW4xExKPNV
J1/dNuh6GAeka2bv3zDTY2nehFIj6Q/2LfPL8kIzAeG6iwJk3BciXq9MDT2EtPW1pc5uLE+BKWdP
rznb78lrVvOSV7DaFTRWfvfhGPr46146Ft/+glzivQ6056rZtBvWOZmfnfJh68S0aF0xn6Y35zvb
vQnM+YBtSDj3c9uA9V1pm0xS/WUoIhwPrRJoCcccSr6s8Krf6YZFU1I/FO3V54ZLEvmIZFDHXbTx
qILPQ9Oh/5VRihAl7A4OcseC0HXSBr+M4yb5m4XwiwxbR2ynSppeiyx+NP26eMOqVUgHc8y6kC/P
F8zGkWowcSuYuUb9u2x1yYlkjoM+trvnAeik/4PXa22EO7/580Pv+Cx8CPb++OzZoLN0TIlUBNuy
a70NwamP92gYnj3UZmf5w4NG0RDTzpK+Qnd+saRA467NXBAndkQs33G3XXnSQAwVVTihyKh9Ztuc
aR3tUJ4GUajtYyiYyFBd1pfmdgYt/E2HfWWhultsev0ObpoYLXnhnVoEG8uVHNKDP9mL4Z6lG7oa
iN0WI3nwBX0r/fZiAtTukpcrmEAaFhPn6xJcg4hrtYQDLNEwZ++zk1/3mgB1d7Tcfp2UkOvhXvp4
quunPOdNR8/Iuoj0oy8YOvaEFE6D5+PV6N5+Ld1dpY2zBsz/+lfWrLh1V2QUspfyFiIRMfhCb9id
M7i6/gnG70ecXngsbOFoOCgVFI1MylbdlmvQq6hI0SBlGclquOZbogxyJG4dZu4YSBOLOry+oIIB
txK2FY/vbk8FvdT39NoDSeene91YYJcHNmdmD4S7qlq8qJySTZR6Ynw3THtjoHVuG52VhGSaEBv7
3xlKYdMEQxVBXDxM7/v4MShvHFI6ieLleBg+g56TS/47EauRPRYZbkfO0VbizNUgSS3jEVZbMhC4
AyF7HeFy02vf5Xxd0gcRsGkwKfIzfr57RAwQBRJhc+UxRukzxVkcbyDUkjRHGKlfnVZUz4CdwWSJ
6BJkunB+ZpaQ7aPLtAD/bm01OjHAJ/VR2gjEbL7sv6DTtmCgTmKoRbemD/GCCw3bgnhwbdvY1ZPg
UT0KSX1f9vJpJ40+Slcr6N/BDZeoYOmXRlNE0Yg1gLVPbASbeCLt5jo2deT22SO/7M6soVHxaVDd
iSWiAJhoW49fL5jDBig58DRZ8xp6jxvBYcV8Lk23QkF7VByS+t7I7vVNkbEMmE52TLIJLPsb0vqB
Aze8OkdSF4t0kDitK4WWQylmKbU6EbHMSb7wMzQeUgW2hv9mDWJ9IggX1exPCCPV1i5ufEM9zs+1
CU/U9UZjwubV0S3eaDTP+YAQjgsrpH6G08883E0Vc56EHbB/iO3RUJnTN2f0T/B3ySqx79OBJ50b
Ea0lgAVUDRAJW4leaO+4GmW1ZBWI42iuK0miyNCUpGOhGTWAvRmORNYO1dxPmF21srEcrdxa66I1
ILVmVWPoVqoZiamFiWGkVSIBn1IaDJlQr26f7NTHoeD0AGRZpHkAPwZW0wyCHKZ/epTFKfAEakbX
LEhAKHziYcg/RmEuBkhhwR3Ma3EuRwzH2s0hreApU3aB3tgUcDRrdvF21Il4xg69lrjxBp/bFoIj
mnnJHQFznQl8aVo0tz46U6wThZBpEhklGva36K+RYLc3LwLXgcuRTw1Hn9MziY08Q2lcuZPGU81v
xJVKsmdXji6JMJ1WBuIAn/KSM5t/Ex6ZOkij2mefpBq+EqfHt6YfHT/c5QkL7NcAwOiOq4Rj17P5
OefexLlCO03lJX25ZA6F7mXmXrp+h36fcJjHG8alp0TNvb7PVChdRetbmP2ST1ZAahBhISdVUMuB
2OPXsOe2QpsDGS9FkwvRjEKTDwP3Yy0jUX6Cff20zvt9LvDN62ML+tC9BqWXXyl37gP3QQCnIt6X
hVuHMPe13Kt8/W0tc2tqy9ct+7sdopFu2l1LqsASWKRWJJQ23A2TUnVLfzWqsexrOGCvIoJq3k68
PavgFOCnFzMqjtWs2P0fKjvRh8O7HcvFHvjwvrO0oBhopO+K13TTXVSXs5I3cP9t0Tb2x99lEWEu
/eQnIE6LeTorjI9W9VRtbBRXfDhS4JJCI2tFt5HxJebXGW5yU47DDFuHD5XW/GU+9HFBKKPTtwGc
0Yoz0/GcDWaskU9wF9ImhhOOPbjYLUdoVxljmzc2awy2z4Mtth/GODd0prz2dDtJgqer3WIsVzWf
e20TDc55JvI6N2qWK9zQLuUZzcdjsYaV3EffNh64YmLa8Vz2ThcwXZ9WVUWP8en8qUjGTe8fwoG6
fOCZ6jxb8Aew1/M6s/xezgct1OmVNKQs+i2X9p+IamzADicjFg2qW46WRCUJwjBZqtsdApTck8yQ
nxUzsVyzgl9atl7nS9HSlo/QnQg8syzHumJjI7bhY5cAqEpEv/kOiIj6Lm46OnMSuPU3rJ6Smroh
LpGdm/GIVjm/ZygcNYTsugVF7JGNl38W7Hl7bY/LnV6XysHOVXy5s/8V1V7JcMIIz1LrinzxIA10
Gi8GnraXseRNQLRVtyNZk5gT24Zf1aQrI8Wldngd9CUEjEgHH8g6DFCKG2ob/Dn0nMDMF/0pvmSc
CKJ2a6S9ePf+LXFs/BvRYrIiLebvN9ZlsoTV4p9uow0eNjWu6gVr7OezGOk0tH4MxojA6uIyXrQn
i54oKuAfbPquArXr83pawEJZiXmD/RXY6F+J7OJfxUTxgGWaCfyUOoOQS3ma+i/v762GHcvxEoy4
dCrhZGKxGuca79HzgIAW/OZMh91cuHufUKwql2AaUkry0XOuHHHqttpDKEOftmt8QY42iUOJJOQq
OMnvaVCuQcho0waNKz66iuw9feXKfVT6aAYjJjzOTF2MbP6NN/5Fjma/+yCw59NTB1luaoaRW5F+
XNqBWEr80MpP8Y7VUgIC0n6l9oPIQjHxCoJRFbqkde51uYuXpmSxQHp4+Z+Y5xbaJ6wMg6oaEVWU
o7vPWh5g6SCegKdx3awPqfP/Ahe23QGVW5uI/J1HLW5zlBBTZidlGGFhAq64Z/klovabEcofzD8y
hC6TPOvUgoCnI9ZS03XQSpbWCD2FHcmIbZkqXTdP/YoKIVWyVAks6hk5Ka1YheSc3WVXWI8Uma/f
zZGKGF7Wvn4sGF/xjZ0JrlcnEZ/BNOT7p7kw32d4vRJCxg3pCuFKdsjIaO5LcJ5XLNjTrcz7nxc9
w1L1uv7dv1YfI9sYMDnjDWEsurbOFhN2ivQKcMwI4BFQJfei3BYJRcqb2r7OTOBIrFFsPBgq9wq/
AI5VkTNd+FeuAF3M/PRIa5gL186oT4tEfMX0zL6SI4hfXKBNkP2Gh1il7fBZ+3eBRD3bLL1kPRBw
RDl4/0tjHq2XaX/8I/jHFm/MOnP8BYoUSzpFy3Uo4mTKJ9mpPUneViKIZJ6xcPBzv0PWDF0CME9z
9c/yiICH/3lHVprOg/UJ76kgZ3U3v3xIqUojTOFKEVpI2Fe6cjfxc1/ioVDGVsDLkRtyiHb5loxb
GgfXTkYcEua3M2/gzIMAgl55hraDfCDFxaqKCsvjYK4LDUWmVG+Wte5clhnZGlGj+j9BsRoeQ1Sx
oQgcgTt4zzVe6ksrT7wZF+46HoAFyCsKqC+h3T/bshfMfpAvwY6HT2iXzeEdZ4sOVqI50bWoqtBm
bJsdKEMwFUx8bdm13KYY7vdvhQGGRh7Pa4fizQYUofVPEuzNDcZOAOw01rxVS3bYq87R6xr+9nuM
GjaNm66BbgLrhTlCO1kjFQBjuRFQ7pe6ht9QaCIMOaHTOSEzOxNUtZf0fKz9XHouACb/HimZLx/h
y+Gw+05DTzM7WxmHFJqFbsHpTL8COL6sDbJxc2vuQyZ2EHVziVi6TGeBm8ge1mJ890v8Hkmb9vyC
g8SEPEqrdKWAxCeGQ6d26DU5OOmye77H+67D+rMxTsgmRlkpqz05tyWsmFoEANk4529RNscIUT0Z
zFD+i8CNB++cXgXZ65ODELB6SsQQJ7QUpdEcnMY3w4j/5h4N1ULgDz1XJat10WMzlcUVEy0IJaw0
7f5tTQxB7xqC/rx5POeHYILz502a8Ff4LY31Ck9wvpJzQ9Y+miP7zMCB+jB3P4UiGaA2KD68rikU
ScnPbPss71voCOq3p1s3REAdWSHEFV16ZG8adgSkWO9vMJHfW16wYHps0L9jl0tZb5184OsqOPIT
K5IdRLfIdHQnnN9/1vSRaIVz6s87JnHrMfUCQUIcDhC959jnhGokn5VDYjeUCFAU7utZCwGHgHwx
Nl+Im1Sm1GMQUR5i/e2/tTkqjbfg88oGdL5P94Oc3BacTqzaG1hI/EZ0PFsQ3zdQQbGFT7zikyHL
OSpAWImAaxX4vqHB/3mrxSCw0oWCl+Efx3O844ahe7RCEeird7tX8anbSl6rknvk2v0WMLM/jkwT
Wm6J3kUQANbHo4P6UkxMxsQdYJNneqvoBiR5iRiTy5Je6dewCaBm5tXmbU1J7SoCd4al+gUuZwcd
f+p/LtehMNGc3O3HQxz1GWHwG26yQgl9AaGsWcRpzrCfJ+cIGmfF+ygQtjurWnEfBX5lodLa2bnS
uzEjxW4Mke7+EUE7oF1YFcSvHkme7QKwxQVnMxjNQTRSlw4dKoA8aKB4HieXKglEA4uL7qU+GU+C
ERAw1kchqmDZDPnN1E/UirUPWios0r34m2kWVw7rb+DPFFrC0cemAN4JwKkICLLY+XLTnVo4SfGI
H2YM5nVmy1Z8lFn3qrf7frfx5/sUkt9LshZfXGQvfKD0FByyYkH/lzuEhVXomnzdscOd6xpyw8iE
a7E9UCG2QxOtMR9HGKNQNhq7kM6dAtbsRoZ5y4Em3QZIxNvoGP94SDBInA+PmoXRqMQW+zTSdxIr
xTU8WF2kWVkziVGrQdRvzUPKduJJl1g4NO8JHJrijvUZn4suyQBCWDdURZWGxLZJ2eilWMnom6o0
Fd4O91rURbKW3+mLPUMwEVU2qwW6QjEKlGPhi3TfOrcH2ZqjDHJMZesydXrAuJAlqGS2JLTDS9i5
o67/V887hGFdFW6lEpBXh4I6PkZFGUYjSi//IVkqZ2BlQNMlbiceLYMZNHuGXrS1gQsL5IdtjXh1
I5TGBqFNbJI9M8N0SqXdK0iCqHw/WOSW95JMFGm/B7zc9c+FgjK0clqYNVItaeK5rHJZ9Gz5UgdR
+iwZVygUR3bmJeQ6gsqwcuiXcMJqYkH8rfMgYzWRyxval/MnRnWufMWnKsPROWJuowfw2XBJmilv
SeYXHC+qF10qboAqu0/GsuIi5DQGxp3Vl9EMLRY/9ApI2+R8IyuJTlLO44m5+HVysKunnj1raGG5
G2JDmESYNZQv5utdGeRy9CZUVCzQH8Cn1Cp+MS4dktoxcGeqaPd9IRIkH1ngRIGlMCuhrrTJGoYQ
spd9G6sKGhoMB99Pmc/z6YqZwrR/DNtsOqiaBo3zzhi5McaUZQ/hjyc3DQO37YYmKwfrPR4PbxCK
ZmYpoH3BIr930Y3DeSXKC82rmES5TlIRxU6SdwE1Dc6Q2s97UYl4dw/dcgHBrLdgmO5/xO/qKzjo
ROufYOtFNzRUbUzCuidBr3hipMh9vCbtzAY8N/2KA1zyUW/evv0Gvm11jWbsLsa/9vy4nzcJqrat
sIuVGULJfPFf4PRgtIxXMnF2iEXhPU0bozTr9c/CMfOMcot2is57V97ysezJxyq503GyoHsNRdZj
x995exesfUxxzUnMGfjhSfq/oD/GCxxR0ceD+IwdzuwEgAhdSr6hFwl9gzhMxSiifsUIwngeYd1i
SBwj5uaU3Ji2goQJb/jyFwEOh2eGGhmehufFaH9iLMvl6QBnRS3HRO7SsfrZ2dfNLRv5vwsS48k0
EhGGp4tLdJc1c7ijWZIkaAW87ZCaPFLYH+LZl0uC6Rh3Y83cMDrHTPzwrLLwgCRLWPWke1lLkAhC
fKxGXqBTWA3jzBJlZlliCXiFMb8L4+UIOl4aybszSkm0mZRJKGR6lG+3YzOSNdirps5RgVb2jhml
487S3OKuAo+0TxnSVuMlwrZkkQaQ94vBJyafivd/p//GJbaL12MctZO3KQJ7AWcRWTo7wA62nAWq
md8+KlIllQgVDClaYEeqbATXnPlpXmFJ82DghYCkARipbpWahJwRpozj6qDXBF6H6LK6pQMf1CjV
xA4UVX5bcSNDyelMKPTnD+v+tw2fpNBZSAJaTJVYs9bike+/rjn4HVOGnpP/0xTgoVBXTfukWltc
JNSYhojIuwV2aSHWAJO/+lbE+kxdGfxbjXzN+3inYzt1vGr77Jmy3E+Mhkkm7P/UOkDbtBFHP2tO
fYKEFwgP0GTyMJAHUyw3aXCbm8AAdEgMMT4/YAid8IXKeQThwYuY7ZFubYCAz0jHfXypgOUpdt0E
sDdESN0AZ6VtjLsugZqmvcv6x7bxVPygSSJUKOHv59060Hjig7JiTJ3ql+2Ga4jg2xckCpZ04WhW
RgVONupC2u4iskNpGgkaSDIfKF7kaOUQckXwQgHPlJM4u7NXkurVtWZ2BQgFMywi7O1A509ZNvh5
B66MvXcaKxdTs9E92JBGxVva1bLJbch13h51eOYTLB8lf//quqBjmj0yXaMVpsnUkrKYyQ+I/eL8
7WNb5ydOpK4+ulSlWEr6Xt+oI0ORknuaInVhrvP4+jzTUjzdOb6UN9V11xEVr9gBc/x1ms2eEpV2
Yy61yWBT6UtwqGTLHP/g3hVsr5pId5K2XB+y7OaNcO/jNSK3d+CTtU3sD+VvzVaKmbU3Mk1yTerU
P0doGWVlwLwlkxTzHKHADsYKn019Aqrji+lPQ4321PSjegtxX0oe/CD+rYCYMBe2KT1oGUz7X0mC
h9D6BEP70MGVB2gEpUBV9bAyvzrYWt0wZUcbRMIXg6WpWN/SgrByD0zYCHkzqQ326GBIoYLjgj48
zaMZF40eSEYGQIfCuDwZ0H4D6bJlCwVx/AujBkOP7kL/z/im2cgjwMBzHsNkOq93uNB0Y8/GaccY
8891EH1TaGIqb37ema3ZL2MPFJtwUFrRFo25O17042+n6u3NROVesDCR2YUg5e1fFoI749c9ehx4
FTs/Sdq4Gpee31gaeEuBavki+zlLok1xUZ7CxlywxwFIbofuvDZjRgNgLBZ+yUZFXYDSblE8I6z8
egSNoQRHgHrpdzVZ7n8x7R9steHipRUbCuirtWD7swrDSMKbwDreQIv2qYw/IXVWW4tgD/R7I6Ck
voq+RgoyVhfqetv5XuKkxcT8yMUaoOQw12ExUnnr5DxdCbIUEOSYLMd3/Q86W/L2zfjpw3NCDxrh
HnZmYcNLryJmhDZolctFrz4qcTMM2Bz7mydoayj8xjIxaMF6Pc7TEcCWdT4EkY9EtBCZm75pI4Hm
Us4oCwAt1iKX6E67/1kuhWWx/8Tk80YJbQJ6yqYu623gpK0ikqWDyTuEq3JqEO51LLhQJ1KNoNv6
morz1oW3Y9/26cJ75meEDuHXkGsMOnehSCfPado8NeItI5PaF5LKBvuIwvtTgB3mi5MVPF+NOs+g
q3AMHEFUmsNzTlHILEBAnKF7fBmRFwOgeGRdWdY5plLbMpK+SIq2kXkoaWEF75bHaJKaaNJKa31t
jyPTLJ5t2QCwRWEyNNneDHNKmEV3kkWfymXI3ksQEnRdtgL2f/LDU1c7u/715b30P9ABM0/A5phn
ogHQQim+8sSk3FgWUKgsQ/vB08fs9ZaUnklOJ9L7gcdm2X6TCcAL2liDZmnGd2/PNgeDmmVUdgX4
V46ZbXN48HB+qJjLfeV2tnTxYhkidbVRIzPcnZB3bo1BCtSBQ/uc1Qg/h7ov6hAxuTV5PXBfwWl/
Nw4yUIX7ap81g86QjqQM7giQzoA+FOe+WCBZ5kxP0Pb0U620g/go9I2rMpzu36X0CZGejeAp+b8u
oJquFB+CBp24UlFNSyGj/IkZoZLlFiRPMKEgs9RN0v+2kzrdpjbCdebzWMrEsapE6WGBcB2+8EFt
s24pUIzGmCpMMOPFgh/c/LfNoA+M8JmyDOlVoFnZBtylDllwRl6ftnrC+eVEPUnhrSVmoY+09NBl
cpGM6kAaKwA2MV+2VjIzVlc/vHDLvr1kllAeqYXy/1runIk50QvUbySUfZ8YdkzuBVDUfYSmWcrt
X4QmqZv2r4dNEJjfl1kI7WeCD+WN3VPOpiF+Dv19OxVy4vKwE4veehMNR14tDCcmuUvhP5hV7DWm
WEUQ5ozHELWanboTd8oOi3JdBUQP5kno0UtIb/xD9LCcGaqJxgL0sPVFp6BgSO1r9t7rnrNb8WXQ
23PxojSQdmeK//6lYDoXvFjLdcW+Er9PKEas58le6121D3Fx12DfPoH3YPNvpR3X1D+vgDURfh/1
bshacVnqFwgFLlcBZpVTu+7WGsPPcOiJdCnFJfNHHhgYGfjZbubsdUBDp0M118CahsxynaV9ypSU
0ePUTWPjsy04DkBCKPgVf1zIG7yCFMFHXVI6n5/Uoq39/Nbs8BLVesWvWMCxR40xlyXotzm/pYRM
IP2pa1wBgYjrivhO2xrLAsWX9NbYHDJmQuPAn+HeFk6VZoGhvjYqgFEtUFxU69qxtgVeeaJjJh1W
+4PpJKu9JxZfhPDNSgqnvLDD6xcDhQNe34LY0zYlCaMBfYOeG1VbNo/OfDe/R+Og55QtKQX8Srzb
+/8ts3wvvU98lgpehCTGXeQUgg+ozV5XrZvn0udYNODMP1PVfCnoTCs7JzFVHZPcucEoTscrz4fi
ut5OKkCr6oLIMgf2HC1NBwQXIRnNnlHI+etPshL82ODZNjZdRX2S57Zn36sOOUPAt3rIr56JRh+9
THjufGrD+3cNT/DFW1OdVmiGXgMPcdpJ1d9lQFF40DtBJzxfd5IiOSkmcvJ4FWX7gL+nandIU4Mu
kG7vgxJKkGsUAKtMrYbi1YSLMLxiTwe0W26R64Ui1wHZ7INS7zt8/48dN7vWajQqtvP3d6kZPWzA
sHkZbXgeLnchXwCGNRrkALnshI7CHk37i/PhgEe/XyIltlry9Q23lKNp6vUxobnkQnSeMjClze3p
y9uKB+6jU6s6MLDuoPTd/dwBN0JDvnsdMqIisfrhAe+pVfAmoB7VMUoXphIPHpFd9CfxDlU+Cy5x
JyVbF4yJw3eqDKPjctel6YOaxxdBQPu70DYc44h2LPyurqMy2xgQ5xMEyP2l7mbdF56x+U1h6mHr
AtKOl/d/uv+XebdXrxoydXrPbppy9597DwpRDNT2NA6EXHSFTpQw+suoFDDTe7UqdppuT845HF9H
nPpefBGeMDVDaTFiPfU4ejOSAB5tFXEUopaWMx2Jy1JCJvhM4n8+sI14C0JiedfYONPHfHVjXWcX
sY5Ozx3nzWB5yczdbHTDPSe7nu0XL3MFGKGdvP563790rsvGeoTFMoGaS5HGSpk7Ftk93mDeor5j
wbtgGZt/fgD6gSBAUvR+hsoUeZyYF+bYxItRUaB5T9x4yfwR25002N694WUVlgogK+XxdjMJRhFV
Fg+Mb79cNTDh4iRwxI8vU8BjMpm3FKbSokvBKwr4J8aY2tKVVOLjyNwhKVLddbx5eLdnlPHhSWFt
7t065gxVmq5Er+B5unWkzRXssiK7W4LCQiih3VS6HI/2IkbMWQ7p3A9EcFqELPY/WgkAbUrWukD8
Z7nW14dDD4iV0WtzcsKPk9JEsEW3gwwgtimpFbgIkri4n2WX/NyQOFQNVcDaJ7CJWP/GC6oQ0a2Z
UL6FcOaldZTo5i1RZxv8hS6+/2OgIXbBanCH0YHa51fxqAMmXE37eroHZk5tT4HjinHc/tQolJtT
y2hwBcIaruS6opJFYJrU/ESHUw+3kAX8xzuTW+Yv3kI08dio5CWgc/qEEFiPZoF6r0Ymt73OwPLL
QYrl/kACPnM35i0OvGvmaNHkmWTZP7sr8kySOV7hwIAqrHYsDJYSfrvO5V1675gpjcZU2Ny3WZM4
8e0xt5v/BMEG9wUp2iEGe3NQJunKtJI4SjWLPP+SaDPu34ZrBKJrWY6eEHMMvBFVgQIIGsmwBOFy
ChjsPqefMCFS49w8IRD5W2Oe+OI7OZy/fY9cPulVTM6dfPHpjdPfTjIBOQ2L8Y+hRp5Jqs5GnAZt
ov/HZk3jDXmf7FpXkPa3m9B73CNN0RT/o5TgkOT3SQQbmK2U4P9fhypzIqx0pA5T7eZIkB+TDidE
5BQnK8EH6LPr4C0xj8DRppZfupfh210G83XSgmjhwWDdwDsENLTzZaw4TRHlXKybaNy0HmqAPt49
56xSzPYiDm/zK+IDvVG9krOo5IiFeqau/CF4LIAlA/KJYGIkKUUjiLD8SJtrE0N7WPuxkceAatFB
2/+22gpuoGpe8XkeZ2hHO9gWnIlTftOQ7EivwW8/OWUezRH8pESu/76z6VXhzokSOFaVP3esEJVa
IodWODoqmI+4qldNYHWKoc9BU3xV5F5xRFI9SzDpPWpgvEueiJtx3QUFetA0GZ4F4VVc8ADlycqb
V3qqqUJFAkmK9bXw024kR1qyJ7ey2jSQfnjvB9pV06C332MAOKeIqtQrcwfLOe1Z+Uq/Vcl68Ceh
gPbGkz27fME8xhXCx0HwOkQbNq0wqfvxJ61hKgXt7rPTzfCXXS1OhS39Xs+F1IwYdhcBG7cuJTdc
Bh5FqYaifM0ztnobyhF6ZzR3p9YYpRCD9A12Gd7T8nA25petpHDK9wLffS/CyxI1jgyo/chE4CUY
L9tEuan6YSD1MVFk157VlX6VF0kn5Yr1Ez5cJurvid7PphsIw8Vo6TNr0Nbc/6/Qne3KEBfHkBLO
RFalDCtED76ISWgRgZOY5tPB4wWNODLuayTCoHiHbjFxmMlpEZa+G21Fu+ctRebPUZtpXwrNDzz1
gijcLdXCZ6kMYUJXcORCf5DE9DFzl5N1o1My/IN6D8S1KiOVDm6o5GVV8Jv8DxVgjrzEz7NivcJy
Twlc8k0AEgAg3cKmIUtuvGSYqHwrrmrIfBCJnpgc0u3qwJmsmYP7uU5LOgbcEla4ZvC5LFZA5Pe5
8oaIZKwlFYbG7YDOEiZUyAy1Eqcp/lMs+LnnFRBSx7DgMCNmgizRfPcpNCl/BQZhymLEZJ82naeS
bUf+QSg4aKPtowXEiyOJkignxjpx9McR85NwxMLtdP1x9zzl3qudkkUoSnhTt/gTRbglRVu9FQET
N10sj1i2TPw58XFI+uugM0HPJY8FIHn81D56rGXSB1UALH/PQll8BN7rFRnVnRTIuVtp82Tvz4b6
J0WKsDecwUrUluXtsT9NMieN9YyRKIW4TbrQlZuEWzrd7ZLIeGijGLs9AsQAa4Odt9oQWYJGbUY2
rPA2YTJEw+6JNpq5vvXNtrNI1WGDNl+XO8FoNqer14vQKlJlam2mPzsYUTrmWZh8RXKZeJR+YtGk
JRbKphbrkj0GFU1W3zM3OG5RWFbYdWu5GqRbO51xlpofFJF05KGAux3RXi5tpbzXTHvUwYqwtwnQ
zGo66HLQCZ/+KP+nBEMfFK8XleYxzHN94Qa8jxufmYQZlVqETW7dQ6QLi+MEUVtgXntgSWayQEdR
FFgyZY6LjnP6bGQDACDBX7uEbAkzU820PMmfQjKUj9Xe/I9VGIp8eRL0S1kqut772Np/VoupxWm5
nvIZrsakZPWnux5J7cdzF0wtl7gjExbbSlZfmYkYb4jVuBJrO+RAUoRNb+PdsF8TlBlmHPxLww67
bj5J6+TBLA/EltC2Or4g/b+ma+KLlBtuO8rHFDpoGX+2mvWq8gwLbv0e537lRfVYVQcfzkHcwpRE
agFScUR3GvYqKgLq+ZFioRfQKE5E4nQ0AV96r3kLB21dFboT3/m2LN1avz/Hzs7jBUzOE7CzIvpa
rCSejxGqKbXdN+9GxBnXOPAB31Dw9Nah2nUDQoCvnqTNTLWCJwSMMy8TUsFYMKqXVPwqJw22btwF
lo6Ndle1BgYYrTTjE0e7cV18J7IdkzQMsmY4SDkgwx2nDwn5WNEg5T0q0ReF7s7bfUqmJgvUjJqS
l14mmNbIp43day1zH1iHWkguAnzCbilziF18Z49QIYFGLR3eeAzI90FK6PkxEIWju9W5SSwqGg89
AVtQvkYCI9BJmQi2FyepkvxKiP85QFi4fILFTcvMPVFX2sM57ReAKd39fHxEKoAGTdT6EE52OHdk
eKzaWvouZi8qyeIhJrVAxVdQk9tz8cv6RorPCLl+Kgvn8q0XhnIl4LWaH2fCYi7wHbhhmiNKzZFM
ScdPL+a/tCV7C3vjCQa2eN+/dJYBMbzHiuAOEvIIzZ+IVsR89dkkll1RCPhLxV2amcCz0xOv67PI
Xe/wYcdZ9LaLCgQoogx3g4xY4sGOf8ZprxpC0zuwt4eV+S7PMnKCNAjVFu9pXSBTj5SFjg2J+dWf
EIyaLbXZIH4tgobAe5ILmzyLpXjRtGe/jjm3tgDwjID4b7D/RN6+kapr+h/L/9Rin+Rlkple3UGq
hQKE5X3ZdbvAShiTodKmBJMM6lQEncSfJivHjtwsfK3Hi+5Pv/jECDSyGMP3KBpAbwTXw1n/IuAe
gf/iTsVoq2EpJ8HBEouI9aoOehVWKK+z6leJuLrxggDJ9k8HJFZT8/kwPovgOxPBGCCX7C80k8FL
O3X7wjZP/DBXWk5whfS9ZsZu/6c6NkCcBD4BBi9I8rOufAHYkQCwSepl0BtgKHoZnsUThCDkwiPO
9jZSR+mW+XWB4Nr2E23/dPgI/R8vS40S9DTe343DCjgdJYh5TCUZvM7Pe/hyVYlFExb6BQ8XNl4b
wdt9lycaa3ojO1g6H6rOg2LKBD/t/WL+IzOZ7UOQrpqDdp7KOuHvcr6IZ8eOoN7C11lVPogXliFw
8KHwiQactGboktbISW3mwHoJYiSgMPwEtFEmEXebhEvnSxSb+9DHD6wDC8RdW+hLT78zpv2wYguQ
xN4amVw12Nrdjye9bYKSEpFLGaVRIw7JwahNvASaTEuugM7eFw8A3T7EewaTUtFhQmfpCFEIBX9k
xqiS/wQCmptSz+Xz8/t5Kte4yGLtHQ0qU+nY87Rzi1Mc1PSc8X/dDb1KMJ2GApo+CcRMbssqYw8P
6MHgjGRDmaLMycO5W6Zy6XvQiu9S5OUM1vj//LEGNG5jipdbUE0kIT0PalE70XyrqFB4EtBCKosN
rreUmkKIiGgrCM425BnzBnGy4pnoejnDX63tOthgIB0H+Os7V376uzgUNtmbSkJd3QSaeg3dHl5M
xOHJt2lcbLTHjwwwLuZdaCstg6LV569431G0HcTjx9G2urU9/7z90D9sSSEZPKKCx/bqUjSieWJ7
v7x29O0Uus2W1J4B8N2VDCjGilqteJSt1f08D7x8FPgAHmCiuVXNhiJlrRtQa/GzuOBNfmcteJuX
4lgp04EZyfvX3cdqkxcIVMyyztVF19ixsKz2auWbk0U8rrH3f5WJdNJ6MTgRHMOfRWZGWKMcdjyh
JOfKBX9EqbXwSshpTmVQujGLbTqcMZAfykJAvG69jo1JzUEwUcfrtzni+GB2IjzCrUlq6p+iTPpF
xlzx+5ZKtxQ4jDvcIVnM43zF7sU2Qok3azrDdXkxvrdDOYUzbxaR2/Mpn0ghfLY6yYqa++mMNm7I
UAfJ+QQp5YHTuFVRG2SLc5w8jByfsoH5O4liYTzEbNBSFNJAqGpPgaNjNC+qQahqpug6OdXjFinD
JWaiEWpRG/ZRUz/yq5ERcfohwqb2aVKj2g0exPhloT2YXz4oJgsSKgKod3hdSs2Nd82Gs/J8JJn7
f+bQ0Y4zlKOvUFVc/eJzmpIWsk7iO90NpiI5Kec2AjKSJCT7rXUGX9qxMFFvpULpVy5W51SDmRp3
h670gfUjzQiABCBb/d94A98tKF8cbT5MtPxmi+Zvnt2nJhlpIxq/FGeiz56Xlv/oNmaWB+81jq4n
OyqGa7nNYpRLiXQWaaBX17xFQtcsUPnipwqJeAQS/HWAs2GImWeDH8hp5esQAlJgMCa4oPGtCZMw
Cquf4a1aQ8XL7kxxWcuilQIfGSHB3dyDfeTbvNVkmtURXPlWWb0z5itbCuWRx1OoinK4yCWLfVXH
ELD0QU8a7Rnyok5/WypZt++nrvv6EEtR5NDef+Jet7W6axvdcymkN4OPca11It3m1Noy4LcSOp6a
qmKN+uTEnli+d3yNBWT6sCYanuMtOddtFlMrWVzf+rRGZ7nSdXa2gAt9Q7aR46FcTLetj6bhIINX
ye0j4yaaRp8GeMFZR8eRlt7JKz9y0LwUlvZvsW6dgiUVaUd1ETXhC6Ps695yz/Ozspe2EoCvT/lm
kt7Nw3oWTJ4Sy00PMbe+fa0Vio/pyhMWF19DSXzreLS2RtsO3kthk9eqKD8gEWFUqe35w+sRNgLt
koATBFbo40jkYPbMOfQQ8UJGDenup5dqPEkElpQIUCS3dBrtShDNXMwfBygqbmH/dQoUzvlUmxJ4
buhSdSqsQuj9Thj2dibMD1+D/Dwf/i7qnca8AeHkPa5/pems9mDg+tWHg2G5ls8GLUFvusK7ctEg
zhI0uHusQvirmrZjmYsQE8SViBIgNuS6on5+Ruy+manj7EuabzZPrkRpJBfKKVhVce0Cc/9blzKw
rwdajhJOZdULLJP8MQTOQwYNZfi94S0/bH6v2GbjxEgD6KbzD39BIITzAEGI1kGO6Er00K75r6qV
rMN/IyCXzeYDu3CH2Pj2gCuinl4Bfe5wu+XxLIXZKhoicK5U+G0xSgCtZBt7b2xprv5EnUGo3+Zc
65a7zlN0NQV+Lgy+kJulJ23rOGbJ15c6yCXTyd4HxTxbZ/F6YFlQn10k70wXT8fEqqXUDYbuzbRt
NxVezAgHQ/nWqJLooDyL8hQ1Qg09pbZGmfTH+CXBvJI8PvfLHghq7DssjXujnLRIGa5MlJhvQyBK
RonP81w4YzP3FS18z4mXowCk4L16d7m75/v5StJ61LNUGCEUms8bQbih1O1gLLIPHYujEAIfGD6G
8X4FQM+02okhzGZFL01I2FJPvx0G+yTjQcCEe6mbQWIXn2LA5+sBmrC3XrOgWFWdPFJpjhvzTPtT
lWV2AwavQltxcCjuuR81WXPrEfAV9md9ZPmcwm9XufuEe/7eoRPTeDKFKmZUd3GzmSLm6StuS8rT
hpq+1+vo/miS4vD6GYR6iSNGvSVdsTqIybrRfmW6dLlI/9E4vkiFcmf963ZfHoF7NLntP0jZs1yG
T0pudZDYGIr88clmr8O9j2WbnxLANxBwBpZctE5qsKFHKmepotUOPClub7YhCbRZ9f4ebrmPPmVN
Iet5sjOFXLafSv+uGXKxWbji2L1KRpX7/GHcvFA8N3rUiRNt2Jbz9rXrXusgxs/FyL+C8dNAyj2V
+M5eVhGP2dCErZS8neG2I1mn5bACnzU+cycwNgHjtpJXTg1HKmpPyBxzoLluzl+I5EWasU7BnZNB
dBg32BptjC1chp8uDgHRRJhZuiHE3a3izErJ2JNBQZK8PEeEkKUp2/qOuWO7pxY39hkIDYRKzqe5
lHstFNjZWxjxIsL+8x+zcwhkXkYCF6vRWISMlBzFLCswVYmIU6KcLpPEZ7trCYK7ZNNm0ezsskPR
xNntun8sq+7kPaEfce3+egR6njKueRI9KyeDN6cO8vNycEl58lw8A91pyCloS+swSTf2AIocjafh
JPO/fWDXLNbD354DUha0p1BdmbwWeG6UbBff8+/UFN+E1AAhl2gdOMjlgzVF1wHdDdIm0wd1b8oe
2UU89mPehslvlknCA/RRjbvYe//5Mg8YugyskGmL5MPj6jRyKaBlGEnHPKmVfnT7mspzKkrAeVzS
ARAsRFxGQ2UxzbnSx1tJPzurX7hErYvpNtWWw+UWPT3g1apG4pYWbomoiJKmgmpmKrwzC5n/wQ3L
ZzReE8wi1J6VbrPggEcIw80ViOYnDWgkVZLjMCZ5+UMsHrO7DEWGEPbIj/dWKFGSkOorGzP9MJqQ
XTls3GJytqOFL6VqwIRzZu8KNiXUkOLgduZmR3mORi6PkPkcSZR/55GX/WCISEt9R/OFebmdD7xk
9emXuGdvk6RC0j6APAmYQcKO0/Xu9Z3tZ6THtNNec2jqWoJfFEK378RhlfKPxRnEme3OeKVNyW35
aaVGRkE6TNlNYi4fXBJuW9bOaa1cBCSQfNVjR8gP/w/ufKSah2tCXena1DZPET9IgUIN7Yi8a5gA
+c32/PU3ytUhXd2o4ek3CONnIZH4oNOkZeIOukENZ4ltrt69fQx3cIxKsvBII+Hp8vOdM9zvcxDW
NE25LN3+xvWQpy7HIN/pqWtapbefcYPu32TlJN9zwzKnSPxnpAQuj5ue8vCpBHlG455bv9CN43Xh
fer4O434TEfFRcfNE5Jlr5x1G7iUEMquDCf6jUoE4/Fc7i7ROJm2rvycxFp/Zb72GgxOOuTxefCj
zSRybmZxQp3hUC2/YjRIIyY6dGe8QgINYa4D2sgPSPS10fjgyBolITc1r44TQn9eOdlA1P+weU1Q
JAu9iiO4Aazq/rPfFtOzc4qfsDf/yLZran0sECgw14i38R7z8SCoqIl/9+NncjyDwwvQT8F3Cw9Y
MkSExggnsChV85ADpzpMeBLnYjx200sv9AZR8l8W91pL7My22b8GHUF7shYxLf9BZhcT4XvIuKzg
n6J4vXxoS1osBton0osi1nOspJh/d/q0+zc2Rbdasc3NM+nf4L8jc7AsKwGXehCHX6iDNn/aVD+k
pzD6FqrTwtjVV+f8t95JnkCyE0XRxtM3laYn0nLn23O/Lx8aJ0T1ATEuEXeJTLNwaYR4yPJ8602m
U1GRGiXpRS/axdSGIfNcii7tdnnyiRpUspYKti8oiiEfeLbNNW0LSdpnKQoIu7xJg7Bf7bdJcPDp
0ol0AEDWgP3ROWFbpIbL6LO27bDJN0kzqb4mwFQazKzXghFEwHK+dM3gNlx6WcSj4ESuekDLbiAu
EQETc+A9A4kBmxnsc9LUTcmtFtJ7LPk6FFo4jM7eRQb+JijDwj+z2lKf0G5PuZadb9QRng6s/luw
lDlAtlk6IGkPuyQQcHvlGo1OMJjbx0PUh4q38XVVVlirRunIvYAxK9lNOHCadCw4ykn5Kprp3F4G
/tI47DsunMCxAU5qB4nZgRB21Zu3uYxQZ3uUOvdOKolbGfnhbXXlpQYwaEEXpVbeLR3RjwdNN2GZ
NzflkJkW2z3jcaJ892fMSeogwxKj2+22f0uSLa0B5qq0sRzdVwVwtHGgMduJ0GLmEqVQ1wzTcu+W
okHAhLynbUQTlPYfTaZmoPsZcnZOEQHv5vfxjYdWdEE9pHk/rFL70SqKfca5PeexeOEoF5zbPK3w
6w0XfHwgZgpJ6WxZSgj/kup5Jxo8Ka/womYpwD9me+N4j43XbLjA4FUACcQ4I2chyyKpwpeZ7s/E
i7wKzquPFVHqBvcoOuyaY0/nSsAUPB+qxRt2J8rHxzbfGxIqHTi/lRALNBT5C6DgkMNlX1yy+Hg0
R5xuWQpWdaYgYb9HQc50MZvHmzu70zO41498feUbk+6CQ1a9kNRaQcQLQQU7koy1GU98DhA24gZm
dwGz8aW1O4QM0B3jvagCcWzjcvIiLQ3v5YQIsN3gXL5oUMACgAzt0dnM3hdZMF1nTSvC7DVepi9O
sGiT3bZ7n2p1/N6mlb0YdprUWZWrCU9TCxkSbMBwmJwqGwKaqYiguRitwwammNe10CXktzROG1P6
FEHH8yQS+5U/mLj9/IseQ7EsIU3l/MW6Pc1h1AKkCc9oIiFcdEfVovXwHzxOtNPus3LQJMZ5xAXw
68l8PXB+ev5AdOzXq/zca5uYETrcTKuiq9byn2JkZgyiDpboG1fjCLkMsAFqZeDtlqRmCO3sM5ng
kuCCIaQ76yCWEFiPJCR9o/CSohJSW4sErEDKQ9FcBH0p+h0Ow/BFa4JqVV0y6yxnk36GMLMIVv2v
nDew8SUpgAxCvFCIv2fiVm68bsgP41dq20Zcg8u4X2A/1IID4R5UUZ7Y14qkdGO8YiTYFKOlWy9D
h3/KSs9F98m3/oMSJPuXmioLEJDp0P0Vr0z9SGzEl//Sr1D4J8ECfCTUVbYMABSAuqADtJD1r8vQ
anAEc8dv/O1ZGcUHsVrsySSHIPpHrOL+1kGJwYAWyG8ChTkGuK/SwL9e2ToJ/h1U0/8kj2OhIbMR
KNDHMvMqlMyPYuaTSQTNFs/WMWohkPy2LqKKj3b3ABqwBAaYNdSkKQuzL4j2prNLfh6Hh6qVjtZK
RdIClxRGhTG2Jexk+undKvk8pm9aA7OpY0VzBL6f9d2oxF7WMh4eHDaDH59EQIqFP5nzHAIHorMx
6Sv1nO0DWGmy1+6YdolFiMdZUO4ZPgfPtE5GxLbj/VdqUQxpxEs5/oYF35Pr7yAL07TuYWYWuMKJ
Lc9DAe8T0lUSFhA/fKj/ExM4Nt8BsCQe9ViR2YbrMhNyb2ugr5zrdFMA/jJUFjYxBWHZsfjLgSoc
mbgVn0bk/OwLKDii+zIr84l9J4pntnKY/BeeWI3OCNkm7AmW8RN8PPCkbxIxI/rprruOSKInqvPi
R5700e0ymtBOlfyxQOiVsO5Q6nehdzEXk8WUmADeBZ50YbWieHaWhkJeIO/RHj819Km+ra/NDIjs
40KsQ/2AKcgIbT9KG7CL3uuZ25PbjEixfF4hvGG6fVkQdwVN9tdxR/W5ni9e3dOahWnPxGMV03Mc
AXxQq7t8qyJ0/QFYSrv48NzXhgJU95jhOxb3zhd2GgcRDOu2JrlqQY/dBCd0bjMxPqNkzwTyEvVI
LbVpPGyTbE8gGH9jvlCvwO9xW2mSYLWCbZ53QAu42NJ6LwU/sqzYEfZ4e/6he1OBL5TS0hSZyS2d
WjqQoFnRw6WlxbIYUyrw5CWxI4EZQ5l/5Q653IqZEXcKgARP27JdmeT+y8RMIZuZWluiU/Dpy25j
3/oktfho6V5WFeLGcyv/ZJnEGcc2ms4gHLY9qip39MZrb9a667UzWnnd0+rC/GwYmypbvQ30xTzi
erSSGAgMxL4XqekI5TAxcUbaEIzC6WyAD8w/6nbEeyTc+sB5utd4X0jJ82LvWwQXkQggIyD33g4H
Lx3dIm09gSFzSHevpJrRKUb48KnfrKEjN0+GOQkRIqzDAO1HQD3wvh9jp7MO+yaFTozucFA4DCq6
ZFSUOeovQUt65JTnyJC9iRQyh11uZN8hQuz4n3SjiNSPmOPFAdh0OyW+u1ij080eQ3/L8WDQmzVG
Pgbe6+vY21cgZ0RiZX+xMW11LHAQP9Us0mO7Cy6uWq6UF9eJFmLj8DJGrGmeQnus615k08h7kRPh
MbkXpyR5pKZd/TJAy0h8VZIXuHZuUFl4WdcFC0sZ7U84iMAGlQ4JnZ6R6HP5SMt++NAvoAJiG9TP
LJZl3O0GGVP0SVrbzpGmtK0ekt4XKgVT0vPrwhpDW5074OViehs6p9rBACliqmO1BaoBeoRP74fM
XuNsDm0EjiTtdbKwExezosZVGWN+KUGv7ZNPDZVAccccAWiBlIK1Svlwbqc1/9/31DlsZE7y6McL
9ySCjjpykCOByB++W4yuD7sdly8rrYpPhVF28gV/vSp79dXxCR8heWNJtmnQVVK77PvNo7vibztR
TWzJhXMdkN+BkD9CXbuRULzVO3cXi4PYpc/cA+UqHVL3mh8bVAvvCdGxLiZOL2PinEqP0m29Y14m
MYBWn6slYzjZQnT3zvDGZcybGzr+MTLYILT3QBNwufW7bsAKoPC/RpI04XwOJBTYCG80om96MZcW
lYua9jMmQz94llif8GrfbNT1+UftoxsPvW7bQW819f719csH1Wt3n2eqKpZrQcRQ/12JMr6UTQrj
XXefvYZ6uI3DawGCKmqLPxQRMsgPgLbVhhgmv54Rta9PI4Gl5oNtHFAP4I7WvGogiv/E17GP+O00
QQM4XDxwEVgrUoDVq/JEuZrATW7qnKjfFQjnfLVFwh/JbrAXEQ7us5WyNYQFUD7TaCwajhygapAB
+8qfsDogfH8BhAzmpFH59sZATfv3F5GEt9/jjkSBPjb6Hu3XaBd+yHvI6SjZ8NbNIGzG0E75lAqu
qvZJi75WucTEqrls6k/5stAP3RqkTofRcpRspSW/0DLegsF/K3NePKtT8padsilK4J5SGFuvUMw1
7EYtSEH849Y/4jPYzEj9t3CSQnFE0y3YU8tXfzJKkxkpuUU023NvdBlk7fD+gx8HBPw7qY8/M5Z0
BsHPOKO5HhOtmYOx+dgvvW6+Du7CVH7I7ojn8sEnY7TVf6OaHEs1aWxzDYP/u828TqbH7uyiy7Y0
idoXU/yUk4vX08e8+cpu3glGJ3c8ZxvyrCib8pbbFPjSyZdHUHbNrPxxE+gZbIVwNZTacb480aj6
6EuIiIbRHTeokThQd04UBJByFFXrLV+hQgBWv+qLA5GZGCd08HIvIHQ1YjSwzYqIcydCcvaLsS+g
ebMdjH3124DhQ0MQGFxdnKLg/o27mRlPEnH5bmGgbHjpRza3kQ/OwOAGiiOCq/BANWozqYpueG5O
9+YByAD3VoJeMawpRRidYBo+Co6NJHbPdm3ZGlRfVfu1gdAGR2ZnAiJhciFbg2driDkmsxGL5xBT
xQHkfGTvjmJdLJvHUGmac/Hb5rPiVB1e255HTgZfzGPovLQuYTmltYPkpQank66cELrbEi6u20xp
afTERo3q0wBeFP8ZgM05x5n4k8/gJDH6AYSwyCwWtNAjaMIqp+Id1XnkEZfG08BTAioL+EdzqMmy
GYIeCmivX8GkBAE8OE/ODE8Ay7hJc1peGXpdUby75VNltiFrj+BwwylAOCpkXjmuipA8rbDSMm+o
Vt9UoZriS9m/XSYMGFTdF9XWe9ZCY3orIaYDJlwKarl/ZQE/2N0Zy9Pjh6vg9d8geFW1G2zEcaeH
H2/e2g2VlBacvoud5k4A119rkMrrsTHTYq6nwxFHWVn3iiWlykICU9OX90llq9kfn9YiZLoS+YjU
dtu07yklwCapVvCiUufWjrkDw5aY9EUrfutZe/d84VGgAZap67dGhtETpj2eXmIUpbHDmzVScZPg
oid0wPLG+kEDA9uVazz96SnIjQ0BXHvDdEJtk7i54PIVANlTPy/ebmwW06XGkAfBiQU4mdLiMxYX
MelqiWOhKnuPAPegA1+6OFoc37u2dL1+R+hm2foDgsZG4btyOGowYq9H472YPQzuKGIzLNC7We+a
QCkhCdHdoXG7MX7mumT2/zDIt+9/z0+eNq8vi+Pi9gaFak9a6uHBn91I+MNNdoruJFR4NLynkbdF
sm1RwfR+n3FXi9ZOSs+AHGERNg+Cw80PmxDSPJ5M42/GoV5iDKpr14LXKTMp6RJlF1eijgttwfWT
GTTljwb9sYVwVwu4EH53h+fsukIF6wrWfwm2yeG6J4UGCBjbpe9F87xcdIK1qPs6tnl6ITuiyGEZ
jSYJbJs0w/wTfH3v5ROBlvz4RxZV+kbp73XOCRh74JRWbLtQ2y9Y70RA+IpCdso9yS7P1/rWnF1M
4nV1o5xygZHbX1cDNoE1x1bKKClrkqk4u4DvOMEy7lcQwq/arDz6XD2J/o+o99CSPkmjvLy0utsn
Q4SHnXP8970868ZQBZ5/1tOtvx6SCcr12j5SNeVQmIJHCnhFsNW8xtDU6qhHHsWA4t7tK8duSGmh
GhV8OqchUB8DnsB96e7g5VYO3F3/Y+fujKwW5/FcMKGrmf20F1TQNCCVNcvXQNDXZ9qRfcJnVcmG
wDxK2hf+5I9AWkBYou+R50Ucjnd9cbqLt7HmU6Ng8RmU2EHPy+FfdqUdcbaOSOwcVWPpI+uv6yRh
KNLPrZcrxog+n8ziQY3x26iacz77/AbzewONMt8HUQplBTEkHuFUOQzW35crhqbgNy4ku6Pwgvmb
qw+D97eS79K6JUa5v8jtEpgvrN65+QKujHE+hvOfOHp1k/PpuMi4QrhS3B7s/STzHjcAqkOJFqTB
FES4UbD8KWsYPsXYQqNtmO1AZP+yppdi2IleyJ/uRqVUO3PeXkWsnFg4dU18GqRLGsxztqvDCjeJ
bULBFJsMp5Rjz6v5JGcCCXBYiCJR+B1IQl/yRIwhzhvR8K62FI4JOtREuGGe+E+etBqPPy3t6XHp
17S4VunBg+xFX2xXxCyYEopd7oKQ9mOFIt/Ahb9RFBmmupVDiTXWJq84Y0L6IuitYQ1vmgOTcAld
iPd0DZMTjXBQCMicsTyCqSzDgnqVz/mBt6OOv7IXSRI8cu4XXmMOLV6HvmupcTWYN6RZyQU/47pI
uP8gkhWHMdlC5e1WPJQnQ0nFOH++vyUdQAnGIW/sZz5OJN0AMsouBS/lHrhcyCQ6u5EDRZfWClSw
q3pdEYQlJTYFQmnP0VGeo/vETkWCl251fW5BecalztDl9ExD3C35xJYlVpjtFRxQIQQCC+efuwx3
g+HiRsT0uJWLbV3a/XVSv0z+nBR8+erVDIGfXr4yXlmMzN+MqjqQgDhTOdDDcckp1iNHg30UfF5S
gYTjfLia+AmlNz1AGLuqcFV1+YGeejtkaNaP98hiQoO/lXqGE5VnyzyVxN7bxiuLbc4PdHQM68Yp
ONYXX0CXntyp/jJmAsTGWruTn7X/tObEt3fUthEZFb5XE6qKt8kgD7ra72nC7KbkxD7IJ4NFhyMB
snGxaZ9cYAlRz1BR72HsIzDsV89fNais3LsoBJq02BxjvbuDMq4GJOsyKoB4ZYz+BTEfS/j/vY98
WWNGQXU+q3obgdF7CziZljFbNyRLM9sW96/6DUcvjbPCeV8gbk9l6e1NnS1UVx46fO5xGEmpG0g1
R376TfsDu8awQQSQK4uJx8ip6b8Kj8qHc3i9wCtRcYtuIQcqim86T1yptZ8+tNP0tXVRPlrtuyYD
dlnX79rtXO+IOTuojz/wLsp6aJ6f43UsDggXviQxDQYeQwEY/DArvPTPMDdDap9rsjE6RoCQtkJ7
4WyodagmChR5TlIwY8PVZWe+i7nd7QcWnFUgQ/YOrqpRGXIkCgmj2YXvG+kBcewv64eG/Fe35y4S
ysmMvZkdFgKiEwR1ZgzgVBIBbFbTbsZq/PRvQARTU0KXvBSxMQS1EWp6MxUlXr7shFfTYLYcHr+a
a1NmPFajLchXPz+kG8JwxhEUAlnA0Q/FwhT2IjD0JbEhFCJb1aDq6D/5eQFXmMBNM9vepL8+VUfw
b79sjDy/+uDbK/QZxGvAwvZnIzz51BPt4+6AaX7ku8wsOWep4ABinAgoKH3/+HYc7wf23b3oE5Q7
CZ/1j/zDB2kAvK8+nojtrZDqqphDB6eekNhRuU9wJ0VeFv2BlFNl2kpL9oTuARuaXr2JvaQv8Yqn
C6mnn2EfuqfySlMnLavKq3xLRwe376OMYff/UACqOgATgR3Ll4ET5DrB2pFC3veWjt/e9fBfuiSq
VdNT19okcicMeQ0plAnWI5LQS5qyd6B6TdK5+gZuJDayPewXc4+MwG7AlLnGz6LoW4D6FxSZTRoY
RHsFgxX+pB28Khcb8z7+wzFc6IyPBUMcgdk3E3nEGAAJNsLUuvqFI+AmaMoT2KvCP8YrBYlaVF1a
5ws+/RXhykBuyn3rbrVdp2OWlp9AiZgdjp4/M6dKa0ERiRztFWc5uQin3KxQ35+fLLdugSzOsSBk
mH7XI9TY9Ktw8+jy38U319rHsp/v1fwPElemEF1RIoOjTtBGIi0S9Q8nRiISap2sBybvyFr1tcAa
fbPPv8vUPltBbRJPTmJ3bfpS7GjCdAWG6Fp5WQOvu4vUZcQOyMKHqZxLNIjiS4mOY9NKz3DuKwSX
cKAnnluSifSe8KQURSI/B+1sPSNJxkepAL4gyNUvahrYuWMWdSQzfD3pH8+gmPi/7nrgyq/gJhU3
1X9ti8FHwEnEkWs/yWHgDsr1gdFFdgWHB0MfR8HF/E03fNsEE67fSSm4W/g+mvKkffigToRnXEOJ
3CrnRELNLO/IUCvVdMTDg3JLTis6uvGjDU/blrT0K7lDo6P+lkDWY29leycsGXSxG1EYAK/5nv3a
M4RGag38/Ap9Dy7WNUDXL6/UGPcrxVuLk59p/pElhnefNfKSTfI22GvqGc6ImHZAFfsG84KbMXO1
jAEQRMCqhQf43wAmbrSzXvAcfEBRdL+9ZZhtUCKd/09kq51RZAJt1MJrjl1QwKjLNgKtGTMURe6t
Gj5itSoc1x2BdpC4HkjXRm3cHpOfKNjEhMM4UO3PdPZjUa/EA+tmrKZKFsUupmDM60uvg9Jh8TkY
ZWUFMV/M91+kb+fTHPwr2c/zRSodeRZ43chHCjtKALI4H8UyZRwEGa0/tOXT5TtflMtPXc7uYljE
oFV7NrqgXlW9JSMv+MDCreWeuwDQihlJyZECKW3aHZlI97TDZgqxeAvPbdgyUI0zIDTTNda031cl
byDCBd2Z7fV09DjtdN7ub8Kv1dMijyy+3rk15FkBCU1mjJ72W+wtHm/tOyQgBDeDJMel0IBDY/DO
iBcbnUsAILGJ1UOJ+YhrmYcA1J3Re+mBSyAAkESuhQfxgpjVpvRUsJMH3V19Le1ZNGMVFvOomC7X
vKuAPChMTx73E+CgIfLhcOLQ+XbBfGpfp7vRGgJhG8nCkxO8gMcjSRgnjpo04orVnCc79S3RUF7D
jpsScx7LNDw+BBgRt5trzuwdEQOxpLzOVO++aNY2wvbuED6stBeruz49g5qpZY2T+1c4uAxUxxD4
nKirYev9A49icOnrPSfMu3HC8mzFCX9JnxLiqzGm7KTRf0kWoK8wvMl0QHFtPknNNMCnS0IuOd4U
z7xEfJcPEPw6F0p3lK1lUeOpXvGlYtF2+AqSHVDdX5LzFHfrVOh+XLV5jJlFvvRpvAnKpdToEJ5m
xNkSMlpc3h3yaH4khXBxn4QxlmZIH3e5dOPQPcNEHp6E3uCHtMg4Ae/1EjR16/8MG88J/oOyU09f
8xCg70BN15S1SflYh2m0NQkG3kuvQjIJlGeGMut/cJp8XJ5s2hUP+MfHHPNcuC6sTeJ0JWGcOQCJ
2giInPLiT8I+iv8JzvfuyZZNnEfX2dtWq3kJQf1AzBp91qN5rcfyyUTOnLtpbEg5HYRVIBMA2EMi
wBLYFqTFFi/93km4dR5iZMxZJKJimPHYIWgZedCavoOecsvQH5B+jKaiiucrnuRkRjhW86Y9eG/V
eyrbPjTunrc6M/5TxnMY2bI9QBvujWhYaknliHahBDJzaX64hXaV/jkfW3sCO52EuqNlH5xzvTfT
rcKY245nNtuLSqLqK9yPWAM6XwfFGFnrZjocQ3I5foRjrJRXQloQZdP/ZO8eDnWninQLfZBz6nYB
I42WMSKeqBtzzQggtR1de/8DCB9Mtl7Exqah4gKyc+Vr5hfWuhSppevuEWEdEW7c6BpiouZ6EQ6d
Vx33AHym4xUE+Ow+fyKlBjiRjr89Tq1VakOZkLuVYAHFTY88M+2vpvuUXQ6kkyo1/u/kMHbHR8Hy
Ec7YuYdgxAl1f7iTfFDIpwLsoDkQ6dnB2fUKtgk/SMkiepl1OuqMBb3qM6QIa1yNpFTs/ZEhO4s6
HBDsd4H+ZvRYKllZ5PyZb9/4xYUPZymDFG0gOHH6KdpVb2icJHwCZ4ojQwtswk3G50JAusdNN+aQ
kpEhdSTVf/fRtMXCcZVXsBx8x4agIpyQG1x5/MF+roAg4Umw4uFhAsKJ6wcLnqsXByHgS2KsRzr5
p+vIP/y2UZZ2y+9ZAVwsnUhrTRVp1I8xPDoAsx1QM2SOabWy1vEEw5OrL7hO+iD0h0uXozu4KJBQ
hLXA0Ck5OugaYXg0KS32aytP3YC433SWBLGmNvVps+LQd3Kh9Bhgb5QQff9s9UWc7ReWy5LQuaGA
aLSjouIGWZf2uhBSCVmxFX5kbCBsmkWtLCTQkNbYdavc0OovvnvoWYwqU0stADi5qjaljtj3rRfH
sCMYzGvtI75VZGxi233tQK006d892k4zI98p8oShBSzHIetqWjrfZOLBuXdv7jXR2ic5N+dulcU5
fMh4pjwWmhNCCaiGFJtKrXuC/Tz5F06vMpRcwonkO8p7TVtpzZW4JZPu/LL/mWFUB6py0A77mBE+
7sbU9wYB1Et2c3ciiG+vZipvk05LlvTtk885+gSuu89RTQUFW3gYHXM4sXfQQLuSgTuGdSS5qBD9
3C/xNv1i7PNn5PfNsUeMNRxz7VDI+rCGX+e6n9X7uvcFIWqgZ/Sy/8X0fa+SXHpeOj4yMQKZbc8C
dvK7BIvhHAW8BKFN7Fq/V/u1obOLS4MClHiAj5UE1gtK8XrmntpnaWh2YpNFvYtM/6+4VYpplM3C
5k9D845dwII28Kv3/0bNaVvpjDf2Zu76QMBs3NeV01N3ykHwJrOyYXQjccVqtDFgqKonKwPkVE8r
ySUXD7t4XTDYLZRIrnOq6tEhWAjg4jtuOcZ5/ESt+Z1W17GCWuK7ukazu59aIL3GZ1gVtMduDIQX
Pa79KII2K/ggjyqMIbcF/hpOBuDFN0lCcNFlRZOZ2VdIDiaHUxwiVf5xCT4SD9YK7aTWODtMg878
kRwz1wb48mkqXz5bjMqvbSEyyztoG0lzJ/N7bComVBJDDUenIWI0n6jFKUHE2lQmP2ta4aStRa2x
AgkMCyXJopylRLA2TcKd1jUXLn/kVODA0PrK3f3A6ogIRTVcTj9bmzXIppkzKj4/E94OJ4vdaxne
mD7TmJhgML3fviwz4IGqontB7X+/D8JX0vThgZTs0K6T/Jmzur1zCCfn+kbLTL3ePR+HfGuzhyAK
WcXjhrBcRX/fNhPQpFywCBd0Ziz9BAM1c3iHiEsU14r51Q4u/lwe1svmHpz4y34pwjd4nkg7BEPb
7ZI9ZGHJzOq8VoeP3INIrPlKHz2LD+0DOM7dyBu9mBg1otnQa2lpe9oZiwL3vcakmNrO2tT8VX/v
KWRZ7OVrRTsytipt5IARToocGUhrjS2jwM3xACQQKBQfbmEvhNPU4jxX9gsPei1hsKeai3tGrov6
0QdLDQmxT/gK6KFmvvcWjZEnPzQKRJJsKbrrIEsyDOgtu3Je4lR8BqZhmFmVEqcPCPKpLMRIGZYv
NDQu6y6cChTtEQOtlFffWmoibJRFSDeJ1SEz7KIGwxClAHLQ89jmq7Jm4NaMKk2fP/qMm8rC/B7g
g9nEgQPPKLFyRfmfqei42R208thmxd6ZZx/2+J1bDGQonFZAdh/K2kZ5MEkebzU/9ic4BAFRgAuB
OMSOlv88PfE721cU/l2IzNZQ/H1yRFL1JwbGsjDJ2vJ0Xpbg3gm1GKGxraJo8XEn9luZhfpWj+eY
GyRsbMP36GB7aVjP+BnU34+kEPSPfXKc+yPvatEh2rJMFm1JRtVHAJdAH5Fi1iAYqJWDRj+8iStc
+Dd7FI/HzRk1vQVbP69hdqMJpCTJgzAgYfIGV2Q9T+jgPb5rTIjrJngIOzhADqJfghQ171DwOl6v
Gs6kGmQoO9uymOE2/5XDS8nLKPpSHC/wZ7fIvLLYjwIxoDcYNxaruDroq7HuB+D/Vopg4LTLoDwb
c3nSw6xdbdNrMDtnB8qvwwtonRRQ6qZlXlnxERpdoUI+uG/fo+aU3YM3cwOIOJydf4iNfbIZBfdr
B6LUssjZOcHgDTjACWbg3WEQYtrAxNuzKfE7BfGy5esVWFGgzGnxrfvkDR/QoA+tM9nrriTtwJFh
eXZi3hAO2cuEupB79yDXFvwHf7Y+HeiP2XSbDC2ecaM6cizcZLpZLs4YmnNgunLYSPfzu1pdj36y
08hn/F3wJJffwM30H/loKSxYNeeyqIy9vwiynCViY+qazl7PhYi1G/y3O1XYZ+z8m+Ffo8NebDO/
1ZUg/MAeltxnsRjZaGoWrE1JocxCjqgJCRP/1V8SvRjq5+MmHVRjlwbe5kupEbVmZaTzX6tuYC1I
raImMnxMZEEklbb1GZ2pC4GxRF6RZDR82Trh1KAitJtYtzqqtkat1UG59pcK2gdRUTPA8YzINT24
KHX4qh9SEHdfGd+L1EG9X2vCJTczGqmw8sXE3wMBerAIzqHwAPrbROythPANxWv8jguBaKvj17ME
GaEV7RaB+cMo557K1EaCoPVmc25K5QzMK3n/yYxussVEPtaQ18Y9Y6ZPhDpADscFhfDJRsdAQWjN
ehfM5rwZ+D8R59hn2SqjHXzOf11PdXl2s4Jbg3kjg/farUanbYsOioB8nTbqEQQ19OmrPTx4r/wo
v05Mb82t0atH1yJu8zAtT65THCrorFpYYuLd+yqPYrhPTD/GxzZnyI9bU/bvnDL+OUn2s/HPVfm+
+kqsXiQYUcvXIlqVHXWHLgHPSV/jiopMdg6Plv/u3NUq8/Gvq9zbVGyCqpAl00ZFgmt8C5f9lipv
wgrTb4H7kqTxZfI4JvTusKm9/WeeVRxCqQt/VYHU6EbtYUsxKNJ4pxHmky+7XmC49v99IqQgHS9o
Yoqog2U6mll8WNfWrll9yDsUfcZTr9pokhi9cyNb6VsFnJHr9Jw5Qd8cL+WaF8llsnOc9/ECQDMR
kmy0ogqNrk/U/l44esyqjbCRrsS0xLcVUi9EA1RSHtP4JuUtIyHM3Bb8kuvcEpOADTXhG2lkR7kj
vy3yslEhcnA67ws7Uf9djARD+BFfXOYh8Tm9TfF83eG/ugShy58B9MBamVCu2eCBwQrRbFRoqwZm
14QQcmUybaKoVelMJ/hH2H6DbOhFLr0+DWQNxm2ry7nIlWtqgm9+koPreI/WJp04D+oVoZ47N1jP
+dGNuuCSk9mLDBN2c0IClsIrlU96wSnfSmNUmsck8BwJIU45ChLz9phzlRxKPrzwIoY+kdb4nJVc
2LK982hJKM9I6L/gn5EdXuUqOjNxb0WzKbftlEfbdOhYMweVzFx3N/IY+KeAdxFYsZI0bWMOq7K9
l1fYHvnOfRCidU17om3zus2HYOv+30XugdZRvsI8oucNfBUDtZmZh7BsegzBA2dOglHTpXYmXkkE
Yi+z5QbRlHCaHZtM3TVPYKUYJuqW7IpHpb5lDuVeihUrWccmMESeeMW14WJ+YeyDP7rNXyj88qse
f9P4W645ZEkXSt+Mi2CrGkeIdPebl960Xsp74e08DptiwdEFa7w//1kS8lqikWhvMTG83C6pyRc1
WJv/+u58YifW4QgKCtG6XTO6+aHYf8NYhpk/EbEjYByMGxyjymdq5tzCDrP8Z98JKhoZK9j+IFhm
PfthryRECr2KC7xkkEtQMzORUZ7eTDqUy3kyApq46NekDMAFPYIuPGbUgoqzz81WRjK+qRI4Zpmm
1gfZ67naSIhB3xWhOMsv0cCE5PhWpmnjC9XzCOIBETxCyrx26V0SiGl0v1bnfsW2LIDDPUyLf7rc
4w79s6wNwaefAp+z0fCLY3Idi3lJZqS7xOIcXRclRBkvVm1U0LuRFHz/BmuBuEkZ7esMOy2CHjDk
7K8Tf7o3YAg8hj7sEeKGcOVl/D/jvvUMAhwwel3jizPv5FLH7JdFwfY4fWTtJndZjh/UTMxng4x3
Hw9Fg+jN5VLOz8fBiTW0UQgQUjizq/aYsZhEDcykw63GfzqrHFGzfzplZRDUkNsPRiPieS1uAGfP
gXBlPxMlhiAFdxVhd4APO6Rabaj+YnZ52EUkojaQKzD53PifO+XTPc7FSYDRPqKP5K1WDes+3j/i
OpbFGk7y4ySTjvTbI5puat/sE9c+Up5mHjNh7g2W922vaj0XvEWW9qSCiQQ+2QXGo5Lh/ckQ33ZE
KdxlfqcUshHRbsVPDef5GkMo9Cz+pVNdGRPb0PbBLKWxV4A/vo2Ca+2+S42v6XlX2nMPkB4kQOS7
4op3rFxY+Ja9+XiM6paxfoOYc91R8a2vpMfDATVylR1VBz6fYqfwvE0IhQUVsCgCkoR6hl6JN7p5
wlAwSadIlWKkH+kYcmj2trO3dIiteiCi59fON6PZElwEhvcWcRjT1M5zRkXVderbBWWj68rFyQFu
X+JbQtp4qcxlbdBb7JfuwM5zOsrj6fySs/9dDgcc1pKux2UX51nwacyg53Kyttvd/yAlnLZrT7Xg
BN7Th+DcyAyDo4hrRmybRrgOAFJ0AEAPP0LFlVSjiRqZG5zRThf2eBrBFZbDODluKfyUZf5volaw
/GPNKpt68TZqgct0+rkr+tLdQl5oR71sOlJOPxWX2f9ewwf04YUo1PZxl9ScLzAlTmhCZTusXRP/
BKhIMD3qPlVRfNrH1EE5eQkx9HLa5VnaxwdTETt7N9CMlQws8O4fifwPE81X15GBS3aRf9X0JAqL
8m8Jn0swZU/JSz5n5c/76QzCoS3/CzuvRc9GDRfPU26ZAzklPBUD8DS3riaHgMZoUUpFU8sM44hK
J5UQmJPQiBEU7m3elRcYSJ7JV8C919Ur5EzQGhir2huvjlW/0OA6yGP+Gvz7m3Y4isGI7Fbx5JTe
FCadlAF8owyYUltww0fF6jW1uZvAtQDL6ZBZ8XlHyfYMsPvNEHNQTgPmIAHSOgeobUkyf+1I4Frb
yJzp1yNxspqtIaMXtaUR51kyWtdGlexJXpJODkvpuIOyoXLfp7m4H4VhXC6k4MrbHWRJdNs5nSzU
rjpEtkrVJul/byUFIvUFl/imwdTBqjolBdNE/CV8c28/1fTxlfAZonaBJTPFlDceuJqqHbRHSgrn
TKbzejZfPsx6ogJ+D+cET8YScOI9obq3ZJDznue8ceX4tLSf+rJihvKOQtvkubstXPkxf/KE7uDF
6p+Hvlw8G/o7n4r0A17JVUAMML9zk1rM8npZB36DqekTwqBUWa5IpTwpdN/PaujAFzEn1vrqRAGo
FcUGkU/2ZjVgc4sz5WEN1cxnDLvupG82Qdh+OG82a20J5uXkqGl2uXNn4+cQSL0Mqq4oLRFqTlp8
hk++M5PYj7vaVdi7RE/JJh/WUOptbFg6KYVMNJEldxN+dzyH9ODfSKcJuWhKxAeS9fQHqLQ3F2n6
O6BMDeNLhXmP5mFuNm1uLdmnzN+WgU6xjjaj2/fm4Bero2417Y3KaAPV2k1uRy6XNw5TERxqS5wU
zdaMmDaevnwmJQkPIw1WsZYNw5U9Uxy6X8DVA4DDO+g58u6WQevgHNIlOBVH5YhsUkvUCp59mYJm
qxiwgK6UMijsklLouWhDHO4Yu2ZekrbZunkmXEb5OVaQUq8DEQ8YQyl/LFQC9DdDvfvBX2r5sYbo
vLPsU54qc/rpe9aZY/CYudNlNPsplVC2jFftMrp0tWSPZC8C6bRlyAc3IctxHThkE2WfPA6Z8iZm
k2R/hy2acKq2UR5E1d2FCdA5qg6ZgBB5Q+Uttb6cAoOR0+RMd0VnyjVw5dgB4vsTR7ZFeRHissgG
ZkaZL5xrg9d+rQybVHeQ+wqml4bcDPNI7a4ruzIPZOAoxc76Pjj3gtso2YHdtH17c8kcDKhvawI7
MB+edyLQ0GiShR8dZ9K/vL9x7aPJ/Wp3c45l/3/c1Gm4A/vYkJzAVFil3yeYau8bxZJ5uJ4J34YQ
V5SxqshD24NOll+YJSsV7apQFVxucyaD9XaBG61OOfG0rAgIJfPiYko9v0QnrMgmoMOUXwUVpw62
gA9VyC2oOcmJqIGuAR+eo+A6VbXgPSZB2wHK2CqM6WHDkvu+aiBJSgn9o6PvaMquz/8AHk75npoC
UUgic9t+Ab27o3sDTury6I8GF5LYQSbdhmBDFfEJ5ZuzdL0mg34ESlJNyvSBe1nZDFIn7ou2rW5E
uXqZCtRsYsdqYJTWqNJy+vZtK2R6iaXSYflpRYQZmyDOLF4Mem3KVELdgPJq+K4DMnOB7A68fJze
Xc7zr46LfxtIMSoE9lxGseoDaJXHgw4q+Vo93Sgm4UziLKKLz/k6tZ/vJhO2+31wBSow4Lf27+Dx
I9aIdm3k13JDc4vdBYXKH7hHXXDTSMdJ4O+LRkkHFCnzBC8ah5tZ0x8ywgSlDoPJ2l2FfniJ+QhW
q70U8yLPqeWHVmwgpAbtNJUG10YFKsVVwwOdvsO/SHnDmN7ecH5/J+1dJOEUflp23CHisxdRYnXs
115rugkjRfi/T3L7aDzGUhUBhPxuABxDB9i7MepKeYLje9KC829bbNfFXy3em9raEpGVsqg0K2as
IiXxjlwbYBccVvR80y60ViSGeG4EDUjKPi9qOMpaY92Q9jfEtGPnDnh8KC4mTHDOK8uMxV+g+uAu
PUR5UTnWLrD07+ju0ftNr5uRBvpkl9a7APxqzQcTKQafUo/mSDFtWy7LKVj+5/dcDRj7CglyO5bh
FnAyNuK9zkULEfZQtp9xT4P3Exripiq2FLue1d8lAXH9KosD/XyhN7TDCrbtywG2hNd7djeEXK73
Rj+6k9WuhJLc+bJ5jzpsaxDJaINIq47XSa+8IXUh5vOpYC5MbXvD/IoylflExtdw04NSVkbKARnD
n6NPCJu87zcHJc2pE1lxSbtjLokZIU6xdC51RjEXXDCInKDUYx8AgieHcPklEZ5hGz27ikku0eYs
zsk2i6H68zYLg9aofXYGWPbwihj+eJZzg9lLuzhmQ0wgSLHNGM2w7cSGvZR8zNxegyVfr0bua46c
euGQVwn3UAUkOcI+epIAZ96NpdDRv2yhKzPuCIQDbyWl4ywFcBYgyy8tcpSNABwGxRu/etyI6sPE
HhrXIAFZqiAiPtewPXvKxX5aZi1ie++f+5ddstubQ5b4WKGKWqp14ex1EeATJBQ3ai3PY0D0BPX0
CgXt7glSxTg5XjCbdXPIOxXQ+kW9ZO0vy5xiHeBILzpcmKCxrb8pIhwIMGN4ajPYVlADiflzQ25h
qhpQaXvQ8/bu1hj0kEHRlE6hzmAFsEQ3w/YNzpHfxvqU8Y/Z8nHs2zCNcO2fOwOCqAiCyxEpVRHu
NSzJldYMtYBlcGzszsRLYmy6M+wSINC1RRc0VznsGNolStd9qTe/+cj5ZA0zBf4pyICnJu2XVjba
Xdp5i93BJMIKK3U0WZ8INUmYRS34mbSgnnxflE78hKICp+S8i9PzLK+Fcf3eYdsgTqeMHT8mgkWJ
HLGE4ZzwbCy6M2beVxUoXcP+M8ivUqyHlVDtjQVNd+2UpWaUIS3w2K4fAAVeomd3ox8PQtYS1dc4
6CUY/KLHiNa07ZO9/Qe38LqTsS/HfxWX+WWR319RqH19ZjPbWB+QMD8mFBwL5len4LDzODJhtQ0e
fNyiw+yQO+jxdaJ1+yGxNF6GwZYCcU/jybLqSDmbSiTZPlSHirMSIxvFS1uEkNtSDzHTY4uMFB7R
gvbOq9t2DXab/t5U+lrd8FFbZIpoaBKJfdwpUHZJGsSAKFWVBNttSfLKmXx7vCK2JQdZLtQGLG/I
P8HYZM9NuJJMRaWLDSVfXaOpiAjLohg1l4SxbrVuQqAmlvkC+wT1Rjb5H+PSaMvNJOt0mQ2uOmtt
sD+XsfDn+43E/4BFZTdAPT4CSZiDsTaude2zLlICaeHrbCWdUbJP8TBmiNP7mMOeXPgzMt8IX7ZX
QTTRuW6ZM6zk/Ycao8SjMm2gXkzDQ0GnUnTAvdc1rzd2mQudUegNAUhSB3e0qRGVdLdc4FDC+WVk
Pg7ZKfPXtEHh6b1jbRpi9dzRmgjRZovAr++U0qLTilcqsd38m5gW2dG9xXf+MN0YSymkKpTRfoJb
7vJJWZc+/WYgBiYJjcu9vNVC7ryLBGkOiswi8LSzIQg5CfXd6e7cgy7Mx8woocRgC9cytpi6erQ8
H5aSXjgGAanHOGiOdjD+qvyVPGjNyIJRPf+aT4LWkgRe1YV7CSnwmmeSr9tUY4J5l5VlCJ3fIhpk
JKawzfcdV3anZQLmr26lxH18EzgfQ/NoYSuT+q42kyzQhfXkxF+UYTb1ttow7suSy2V94aA7TuDs
GS67GlIB2pwck7mLd8qxdelDNPrLKC+DbcZpSUm4qKXUndB7Tmpha0rq2gusDZDCnpk/OwV71G2z
IvskPEin8gyH0MJWFWvAnX6uwuQVNCGHPxQNojkz6kZFczCM9W6Y+kN12FdYH18Yin26IBVttQu3
q4heVH7aHIt0f0ggj2lVGjPdRrqSVnAHTnzMbWfdO2RPq8ycn/j7Y2TSt9BN7hbtSkuEcdRvjf9l
4aw9kpuUr/Odom/7oCabLj0wZXMLJnnkEj3TLS8Sn/zpWe7qooUjotPf1TdGCmnMZ3gkQVFErXPu
5JHnBp3yhfpH8TZgDN8R5wBKz3qYCYQNT44flnJCwzeAqCNYDryHZYczXuSmE7XZ1QCT+lsD5xe3
s7hBTi/lIVvv/C7K8yfQDNHWLsHePmwuSW3g44puAmfa1CqD7Lr70q6TiKGex2a6nNq+5foPiVfV
hX4V3d1PsMWga+/OoozlrNFp29DBcJhRfEtg5asjquAhYP88X3w4iYVgtp+6WqSGnhs6wlAqnJ1i
VUaTycXbSEnCkbA4Xp9J8fs0D2gRD7tea0cVWMEnP/2j3dGC8Ymw+2eXjf3Om897wvYqwGdA6wrQ
ovPnc3Cxd/DTwvNQIOJY1u1j7iMI/jx0C+AW85JjaF0xc5fAV3kHAw8n9mXotD9fx0FU54K6dj6l
KdMnRkRNFyjlEnqRy6E+TQWX9Dmqr5NLlNytWIQwZfEkFnG+Yh98eAh9ITIZKbwcQEnvDAO3yx1+
rMo9TLfNPs1u8V05ddIsWYUzo/unvdAQEA/SKlek75Lr+DH8Fw8hiMoQ2pkvNipNrjq1JkzlS8EY
3KOSbSrZEFYUovGRyMU2hNQMEltVDxoKF97SEIkXwTdl3JmCAYSBvWZm5cTUr4DXbL8CagLTUlZe
I3aV79cNs8m7b2Rh7mJPOSXUabtrQeLCHLUkLL+1ummQiDLKzUZYban6iZvc3+eoX86h0FlU+cvc
wOkc6GqXFvf42GEQemHcbAoZrtILauVF1RXkabtD4t5VXYhiZW89YSmLwUcuXOQjCiC3Bhd3ge3w
3eIfID/WiYZBRArVMZDBdk0ZVeytz851I95TOJvIfhvm1BSBFQ/RCrR0M7asc8L3tfo5uga+0kfW
QROXNMoGmLO0bVCytf5e/z/wZa2sOwwtLTOFqtS4M2x8j8MYGM1IK8NwVeY9ghyfGxDulEtGN74M
BAopes5YA+8CcCaje7jTL62PZsUKuhBHow9vMP9DP9FAnachnFeh5O/k8u/xSSEc4pUw2U50bU9X
muJf8chqmritBT8lfZ0dc2KTvUAd2IBuP6pSBJ6kAMgJ0aVnZyKdX9DxPV4TGBPehnLcxI7VJZkE
ODQwlh0maXgsLttQzkqwBAbD7V29hUYMaFPsPgBfwU9xNciP0zwUpQZt6rumvLKhns0oqyf29e3j
Q69O+n0b+ClDHR7MRBJgmqzHTPZK+GXK7UASQar8DyqljiopZ76ZXbKYTkmkgmjvI0MUEeLTsqa5
SN+bC/sAcHTkuk7THj0hlqLf0SR9Qqgw3Ixxgmbs+tLS23vJnBau5lyrINee48T78KySYkxz8vHv
BaW1pbWILxJQNgouuXnCazaOzylxVX/droh8Vfoq8mzUcPh/KtBDxSR8d/yUE/MnPaYQgXHmNw1x
0DURRxb3zJL/6DNY5AAxXfuet/ce80h7PWUDRr8/D8HuThGhCqDfxFqZo/+eH/TFWJW4iApDIYeP
mn/mhg6rNua+SfgZBKypEbFfPSlyVsyvCr6UGMDoC0V3V2DD3pDmgwhErqxP7nhG5M/QPsdptuAl
7ZB60lTSuWTpwymdSa0sJ9Sd9+QPDyb3ZlgCbCVNRF890gY0myr9zkH4MgcNFvfzBXsZYyusqj9v
Zf32QjTQYBP0/HLxdH4CWqFkvpyW6gWp1KoCHe4ItAWXuBGtxr854JFTIIo0F0nXbyhLKvfzF0zN
LX+QhNwOHUyNValL/a8wAmsrBZKje3VfgmFNr6Jkke4pacu6zZmUCHMnXX5B6I0WTf2vhN88Sxcr
p3BqdqBMb8ahtzpwoJybudEx3/xvE3OZmIJAlO5RtDkDKTHHluJcWmYWg971mvGEnlrL+3NWclC8
pG261CGQ7Cn8BSFtXcVuATpBzFve8Cu/Ev8xiXTtDBToDJlgj3IQCxVF4eQ07REWSPLYL1TxzuU2
0RSB6RubSuqAkV9p4frT13/V1t8x5jamk8WFTKQvnKcRz0alE1O8plIVpUHPeUdG+XiphVU9XXLh
YniVb0q9e2pLBEDeq/DA+C4ByCdVEe6bqVp/M0CGzjH1Lh5Ns9zmt0t7njUE7y2OUFfSNPRW0xvN
RCuaMA3H1FR3wy07l7uPvtTT/tNDxAb9hxONiWtCQ7Z9pwy/hLX/cVEzCsnlDwNdTmjYCo0fpV9I
JFikLX9x+1IQVKOlCYKcuvGlxsp5tDce+3P+aKxbQU1bMnTeoRYEzeXMk0h7RuYbjs2ZRkmqtPSu
SC4ehoDXT1zd+GQ61juYvfXbiVB0FOemyWsg++MNtzOnu3dB6FOKOSHVdnXBbcFJwuVxVQt9yaLq
7TlNCjL+kg0/mgfM8VJHpcycR50QmuklODn/PSKuZx+7YpXAImS8bVG3mJfT6x3E8fUTqZxAI1+A
hShzqr6etuFKvsVm/QVNgetrAtyD4QBOqs2sbAKljH+sOte8ErY310KR78A8wZ3DPHJIQN6sA1Vs
4l/cFwaap/Cxz0lmRKv75LEUPTcGQjV2e8wLwvi5w324aGDCjHRQYf64GWvFiwpQdm7mgmCAWCA2
ZDXcgpWANf7nrsZhA/oZYMiZGF6lkw4qUTcBYbmOcMp+R77Uuc5yqXnZoBH4zwMdGt+KSIGE3K3j
lLA5mbvYRpYgpogEzdmrB3SlLixaaDxbCHbqEwy2HfeWolroJGX2rzmSEwjzL4iccvu3KQfMty1p
9hsAKHFuglVrXDpRNm+PtyIT7efUE9ASyHrouFuqm2tCRGb2rTz2qimWwEOxkoa4cDFA6lRN0lGV
o6D5ljA7dz0CdgDks8Z7FgS5YvC965iMcgTGsPbzw+njqE9gbSooJ32Ha9OlrsMOKNmXuNg0CTBx
hojZlLGfmOV/MiSAbB/rc2J6Sj7lz7ovt/f8j1UNxXvA3e+a0nsocGpja7zIgBOJAdFcOjtbswBw
eOA0Wu7RTRTLUwj3I1Zs0AFBE+VROkRr6ZRbbQ46TPcwPxG2IKEWfZ+gClTcWY+4o72AwN8KIT4s
SQwaSUr8TkwhFLk8YpYkyyEHTTAQ6+QJAPcJn9W/3/R/tHR252CK4UUKonp1Vs1yuYUEWVdedzKi
MUTBY4lnRxIBeBqPzc0pFBgIq2q4zfds40yWp0sUCf0pXlEHg1DnAmlkODLQoODOlKWNNQ1n6X+y
lOqL/4Eq4AjI9TUepZo5w949pSAbFrRyUa8FK1wyXGW3xcTWMA3hlz1UAofqxesZvzHw1dNxBhsQ
8ZUTOZcxRDmeeLXkhKf97GWYEO5qxGnWHpIuf6x7/4m55cTPldBpjesoHfqP+AmQfDhIBoRLOBC0
nc6vxSoKguzo+6vNgOJpfMCXeCxMtPKcmW7wRdnxcljyNFPnl4zdaZaM8x+lHzzYfUrLi6cxCyOY
ILIdBtmr1ZyQKRlqDD9bAXrpNrGJtct+F9j8O7aLAkiCxc23zASYqakjDM2re9gs+J47/d8B9OMx
2Vfk6RJGlHnP26S7d0RRqBdW4aKjV9OeF/nqkDMdCViFTnjtwlZhS/KMfkxECW6uvLQqMifd4d+7
DWIm3lS7LxVj8GR10z6rXe8zhsI/Qa3+5wYBU1ZY/5/7jdUF+bGmdTfzjviE8b12M8PxQQyRo06c
jdDGp2ITshIrWK/4ag0CobtEUFqwbRpK2yqznSfyaxcMPR/4B3djtdjcHqXKl5m2rT4gUeiKaOcY
l9NUtihoeyXcCM3iry6bZKNu7k7F/xW0ysyXfiAwXtZNAffsMMzh1Gko6J+jVdC+1E8dYVcse/em
lj1fciJIus2uJHXY5fqSNJkOqyoo/SW/VgrZZLw3uLt1ldCx7Til9ML4XRv07AO1K4GMVibcvrvl
D9aVGXcgtPlZE4cu5DVP/bOQN3RF7AgoSp8pyt6hdhTRNamXjEqNvr8mZrz7DRQlkU09fcQikyGT
n3/Ai6pHR5tWc6obyMGZQ/DrKHYKzCBYOb+kxuHJLzXWdDbjkJo+n/cH4A0/9Cc9rLY0BREbzX61
agbCdboZwlIkO1g22zEIi18yVMY6qqBHhChg+vDkXXJ84KN9vFv99QByE4yYBKnBPkB+4ui7/EPY
9wd0jye3Q5wLGGPQQS4JAwogj5hd6d76IIQWDJo/udON5kB6EVGjoXt1rg86E2bQjUGWFMMouIWx
drFur9suC/nSmcN4nWfYKBafHPLrwVa+PnA8NiuZG7acP5P/oh27ZqTPWfO89mrbozZoodJyQ+xP
iicj92iKOydT3zEIpIPfVVM+M7iasK30CtYzX4qyMjT0mreX51r+jn2L5fpccu0tCo7N4kLkt5xT
jYF6oTGORgFwJ3SJuMjfzzbr3dVcp6jr4dEl+SNC1+D0EGidJad6HQ8N37mUffdBhIXWxDk2CF5A
iMOEuc5GUPyGEJcENZy916JK6Dyx1EJtvOL/9coW6ValJaYiPukZlZ0U/CgIk1FRACTMBniIo3wE
FEKJpYFhzuxcRfAuY9UEvXARv9ZnQ9r69/xyKYsnPcprvowy493xbvORuTM3D0kr+8csbCSuNX5w
EvwdQFgjp6PEgIRtv4wv/eWeUCV92/uWrR62exKEsKb8I8gTG2lXf1nlQ4fSrdm4Z+6Bb2HdJ/A1
gv5GQ3A5YRb4/zx3anpG5rpNMqBcf7y4v7JX7RZm1pMhwyK17vWbG379JlH54FqsRUV5WwaDTqx1
crtKURHBvtuxUxIGS/Azt1xeKXkoPkJWu8DfRdgqkt6wG2qKhd++6gr+CJ8Z1mtdHJTA3YOAn7Sd
M0Vm3CfRC1BMrrd8p3rkWW/bIuozVX8QTXEWV8lLf1k9YOppzGXcmJnJSGtkWbrLgQhtX6YG8qVN
o/iOAHz6+jidK5UCRhsZ6lfXjCqPuoz3/uj9fEWU+064StztrlFeySL2eOjPiAIr8QClDpp8vEpH
2g+eT8GYGErozeMx+r2iVQrs6VJDK3xbzNBXtFB2S47Z41xnSUlx+Q2oeqVh2GrkT1/E8BBTcgYw
pUoS85aVfvVbbD0DsS1VNonv9jj9nkwGucTNZ4rQDfHSjVGRY/Jfiux2VVchJrP+L1q8JNNV06PD
yTRa8FLxEuxwXYjOnxwDLn3wt7xq6K7fAfRIBNiOxLc793Bpzhp9QdzBEUfs8xMC0zEZhKETIBHl
Pig6iaWC3VM5b6tP4r6fNl7LPDhdUqiFdw16sCalQd3h1AI3LmLK0J2+CEydxUeecpqzY3xgaJ/y
8t2mzjbrZKOrDlJbyHb22Arc/lJ2cC2wp0LTewTVQZL/YHwHSbSL23rRxQS+fb83EsXBSQEb+Ca5
6zN/kbUfbQX1cKY9/lJYC9DfToJV4L/4SGtdv8iJdVu4u9GZHaw/BzWHcJitDhgN+YslgLYa/Ww0
jW9qb9xjTBJfSrE2HAmRWg30egcj5Z4nzvSRzG3y1QSDeMDpDgFZN0JlIq4ZJux7wJsrTA9H2Hkr
fR4ZXUzk56K7k/QScby0bcog2AbbauoHyiBpYLaEbLsQSKoKWbY8DFWdJ+nAlazpyvPDJKGhcR2y
9+PbH5Bdu1B3NTWYH9n6/TQufp2oWZQBdSlrmmkTaRlRyizvzU0NVYCDwHBlRKdOIOG/P+CWbWFk
x5/AVXRYD4b3yr7f0ouRc/bBQqJu+6RZOa3OQmgPzxB2o6PlISoEkYdKIVs9oKyAR9Uh75KkXGcS
y6qNSuOsARL9yg4EnWZx8VFaIcEtsrMWmw+/lw44YZm884+sNqGvG28nJI/zwQwFg3YMu20vgZ28
VSJhOlWSp0bi9Y2LK5qGKhkDMGaulJxR2lCnsM6Qt15OiqRHS+1+gBmkTMoIjDu2I+wKNHjih1F1
gBz+ZxzFR0MwniD2aXPc/ssw4aCpGAOtr2HXy5NwkzlfnJ1NflQ4T7hdCl86vrTF3D1xB9ZsXnd8
YV46iWwgZLXzbIq9lB0kM4gGOKphDAZwAz4ux0nbSX8aDcdSkZ5sdjiSqqdts3ZktbEdwF9BmazL
VRgQNCKl3JJQ3NGcrRJ/TjG62/3AAmIyZnlI5vZLB8Vcj9kuCJR6RkofDXAhbGAuImn2OLmwOiJH
R1aiNBiJI1gc3uFXhYqomOCSzOELmnBPr6LfcuRZ67swHXF1qRQb3zmsw72mJlsGNWkNqShnhQpG
EodMGcvKDiMQpVxXWdzG0PNQNAqWEU7hyGWisvkXPVi6h+EfCKQI65DyM0crsvADFwWeK8dQpIOR
43IqRFMZleKrsnVHcwUNMC4TCtfC2EEtaswf2h5/lcqoDM12fZYS02pgCS/Vn7qPY+IOp6PeQOii
NQrNEkownpTSyDFFOz2W4HueppaUf26iaopZTy6b/f3pAaaGuc7YaaEc0laenP0GvuVD/0ApJDOD
M16ePATBiBALaNRJya/6Z7pxhtJrD0nkFD37iOXcDvdwfJr0lveINhyYX2I6V5nt993PLD5hfPAI
OGBwGSdXoQv04B+l1AMBpuD2e2J4PjACFaExYOKktMLExNvEibd76Sx5gIbaeejaONIrc3X44rMR
2bO6YyDOPuDT837AR5ZEECSDXb+S1f9W37XkVIXQB4CFy2xTnncvsJZRVTlJh9Np/SPKdGPK0cwD
XSI4WdJnGB6w9rwk7+pX4oDnNugfKJACWFhVNOIiQ9T2Jl8FoY3iCjw/c4oMMoMLjnew4maw5ILY
q0C3hGgRTgvYFUPYDDrKf5Ectyg62jXruf3vQm/xKLIYccna36xeEMGPpN404+yOWCbRv0wQueiQ
v5FLsDRkpSIXiN+rbRjw82rFVxm1iOSFtd6+nrlJF4/Yr5tpQK+7aDH7tqJgSQMwgr0mvududFoX
wju+Fj+sudU+QCi1HA/wpTwTsKDgGMJApzNXg0wjJL5BLkfK/Xhba36gVGIxCraeQyMD7tAZhwoS
ytl3DMnGzAF4FF2vFEtuJzqTUHrpmujngALu1AMpnGH3P24OwZRazlDrt9ZF/vKbQ1SulAV6QtmL
gfSPGCzpqTYfTGQE5Itd6icWJcwOMwiDewS0L+FI2HF1BaVqFlUa7L/RpndyYZK7pV/RuMvZ3QaY
Kik5t7Aq/KpJnzz0zARrzCA2MR9WBjqXLAdSIUA+h8hvyz+BPINOgr9pXvl8B79IJG3FMpcGHOxy
/FNKYNJefp2hxmIt6ELiiTZLWNhO/oh8Wc0XBZXCidZGlEaBRkwSIaBBzo7y7KsFqwRpE1H2Em/C
Z3vwHDbQ3Uop/4pB6fYe1V97ODVsMJffoecXVI+KIGlKokqZrTh2d+j6xUV4SNiilS4Ko7K2WU80
7aOuo3BvLk29gCy6TDoGMkUTejhLRIDa8dikHP0THR/Qr4zUqPggKIBd4mGrQ/ggczOGFyaX9OLs
G/vKcPVHogyWtMoV6Xl4WLh7tcb2g+6CAk9drIWo0fU/nsvapGZKndfOoYqyq6KoeE9u66nggBI8
mp5SDV8ez2l/FgCkfRSks48cp51UO1zuiFKsMZGqJvQWKzrVUz8BJQcomKeuDLXMPeWyfcUV7aKV
hGm4lvQ5R0fd5clSWeFwu7evXGGjSsUKCc7nTbu0OVX/k2wZcELQhk2LBxCGqlobevPJpz9zdZVV
iQSbZ3Eq+r7MKPhVntujDqEUDKB7bjxicHiEsL6vmvVSfNJf2fKsfvyd4K85OYdXutceaxZkFiNO
RRUhpuvFsPfnE0nL5eY9L79LC1U+fLju7tPLZEfFBiiAeM+LvHIqeV0tEunF6evgPadJABbN61Ot
FgxIzFynV7NLMXssiLDSBUQtciicBZy79Gk7lp7nbCL53aA68P9FJ6iXItTNFV0r6oWbePp5WR0T
ds6/O+jvD0CgpGF2tUFPqciOi34dsjAyti0DwgJiDFMYHOdp3nvel3+xGxhTIFj/SiWgZm5hz3yi
uhv19dq30ZsQZ8iBpZGwXOUY2dWTgAPKm5o6ChqYJNWIc5xGIBvCC6vMasmqRtNLZeHHCtq3Mnyd
T/B+/DDpeGUX4GqCdZtxmzA/rXYHpH3DG2YQLX+2eXB4N8rqZR3A7z4V7lb4heTVdrGrjXdOiMEI
07UqQI9wCEmCEn7A+y/7CLRmgxoIBYB5XKv65vBSNZfneG4PPlZPq+pzGainqHO7C7pAAvG18AtU
dRBhAWMe+Flg+Yk19dWUaP2cys4i5TimfTjK0rSH6fP1XrvSXTTXj59aU+tVpt4+7DbMKgymnRjY
rRsu5DiFDJrUzke0gtkqOAEx+sz4Vn704oqieAMlSJL7h3Zgq4exd/37rSknaxglkIz2OmJ9xRF4
Jv8pG+IB6iWhcT5exULVbjPXQ6ToIXnSj+A7joL5j/dn7PM4k2TMz8WPN0yKcGEIPTVcYUws/xl7
Czpqq1wNWli/Q5Tus61LiyvIkM4CxuPaAi4WbHyUkfgqqEv/bCF2uDlevX1MAanGg+F9SwrDsX5N
strwCPIxQBEm5ux9EiNz9G9xd9JwVOD3tmoEpwhygZPa5KjFEAPFoNk4A/CG52waqaeDBhBfyeZH
yD52kTCg3aNdywhFd5XIoPf/erEaHkuha1Pw+WTsUy25+zFNxUgtshB/Zt3dRNjGAtlxdlyalExL
qUvqCYqyDn+atbQz7Lrly5Ye2XPuNWfzFmKKOA8dCNsQp452bCmuIQAyx1fPINtZHx2rByZQYAZw
jw7n5j4uFj4gzJDk1Xg+CrBUeMAe6FyK0au8F56vjK+oiXvI+rymp98o7EwvW0GPV+yeYTGq5l4D
KrSa5YadV92uDacDK5QiRvHvFQ3waCj9XTRau6CJkKuiSNtrxZ+loDvBiRHDFClvuIP5TFBknmRT
P7KcTEmfp8V9RKsmnFUz6N/sCjv2SRHQ/sf14bt0dh1753lr8MpunuG9su7rsePjKuoTfewWps8F
/BTgB+FqUbuRUpBGWr0BaVjuod7XnRrTKSu6HBG+xo9MpBE261/nyJBQcYz3PPfDwCbxL+esbNth
teYI/F4n2g27t9Nd7y/CrjfZG/+Sn6NnydN6yeoVvPnc4Tv0k7h5XVAbbT8xx0/bO4KurFsO41kC
9pPuSCuqVus3UJ4xXiWFU+iP/vLJT9b6s3MGbAueChgLkzOcEyiG8ZXIomFXX8raNxXodaTb+SZ/
/aNXep6HwGCXkr9ufECu0XVrvsmDS5iF5iTN1JucPOdAId1O3jW1jCCipLzTq3jKo/PREHnN4Neq
5liLSYyLYIYKGrAfQC9f3vBPKwQ3zdonuXwP3zj68A3IqhJ7ZC26nh0DJ+0R49+UfGEQxgEG42/0
L/fBA9Lor2j2aCkicK1dOMTE3oIOnDPLTr5W/kZk7+kZjko0zsiUC5rNgnMiBSp13XX/V+QCphEx
FDw4VYvpfHyHj1az+it6vn0Om3WhTVeRFK2gcbqDyDFkDfDqaPfx9YoNMhRCNVi7ViCVv21an8yc
rkmhzpnuA1GvufGMAPwbfpUeX2v+I8SIrdO3rd8gUJ0wXHN61UQuW21qOU7N3zakLB6TpJzTWndd
e+aSxiPpCSdfbhsQLtXflq2U8pqhLJx6t8xsWy8rDMIiVtU6iwjllwO3lsAVXbjbXOop2vkAuZ5Y
9dXf6A64qWaXPltfIQb7Dg6lyWZsbCi7JOuIkNlYN1c8JGYEMbBfnwV6IwihLk4R5HilX9rGLjZ/
KBdiWeku4M4WKry/YlhQJ08i5Osz5m8Ckzxr2vy9Go/hkCzaFBcb1uYXUiK8RqezpmVybpEe5k4w
/o5DnBGkreyXBTYHq3DeJAYHPJMdjPBmvmmQcr5QVBynvQHZWWbYbrMk0f+vJCngiE8OhCj79xrR
onMhsJ8BHmboSO8J3DjvSEFiRAcP6uSg5ZOtclO9m0FpEWhKVXXHTynUU9cusvLkN/d2GzlAfSdM
n/du87G9nMj3H8MZhad9Q3hi3DuhdOA7pgDsmwLfDcQ0YUXiOru83Thav98jGhTFDhZKj5yezunX
d7QwPmd1PY81hpD73MtLaXX1Wwb8R88cyuyhJjlHSEfOJL0k1gmy0es0CUSo2TygaX5pMDNuwP/5
qDmxvubDT3wXgMlsbOG+Vq4nK7rTuJeiXhrUhBvSVvAc53SNDcUYfD610JyI+5cUSIy3pdOF6pj8
YDiHlswSDBRLh+PT96V7Zy9HZHJ4rmis6U80LIVQE9u2D+UICTXJm9iL7yL2tGGpM6f18D8pekvw
JN+yxzdDLeWOsoqzx58AWohltc4D8K9j3NF98gOji+IfzMvI2veCUpg6rXj5d/8i6LMA/ZsXs+S5
CvWSfCtbE4TL5lzSCNsS/wpbhQHgW3ucItFKpbGvkCTPwfZOPCNOkbzp3xBCZwme9CfozeaSvKFr
yULwg3goGWAIplw6ln/ahq34ViWFn3iCmjdblu+Q69z7XXdm0+T+baTpj+rWWWuXflb2qqnjCvtb
GUXxfKjIettYiUdZyNPdQ78tkktAmmO7V4yZRAzwXQ+mGb6Fyv8uadahdMX3vpOYuIyh3dRy1eW6
SPdoO8WFGB2HH708qXvfdkOCAk12YIneU0qKATHs/C+Axq+05iigYTdn28mWzVPlW+AoTJ31cwgp
IQuacu88n2SRXOTwElVIh5zp8pncq89ld4AhRHTV5efiT6LxetljgLFq+Mi5RDI1H4hEm7GTTEk0
Tnp+bXwQBe188tOyWzPPXBxDd0gJCfPJXbHHaKUyh3PEpAq7m0CUFNAgpBozcr4AiN5UbgAKDZWv
I8vsxI7TjJjfFUKwqZV3ABerXajEgmZfGOfubyfdqAnsfobVZ4nPFQ8aTQhuW13ZqLUw4bpGiQS/
2dsyBc9KjPwPnrj7BN/xgGPi44hjVVfRqUhZmQyF2vote96MWOuWBQByFYl2GJiL93aKrTkzW6nj
6niegH9hltatDWMgiGZFDyGhZGDPSvSePDNKmlzSiNGS9iivGdcrtzRPdyO8oAJh8qHUrv2F1pKP
Wa8YkGk/2b7r383KeRatHXIBl6TTZDlcDnTEDLpChIfyOuBSRqYXrqWXv4iN4vhxAnAnYew8gk1d
bHYAValOXJmyG6NuS3SXBzkCtPKIyd+lBUn2GoE0KOPN+fQ88p50Q6kzQLOueRSBpy2HPelrITyc
2WP3h2hKxhHEc45fN0hx0A8hs0FKBBMX8Y32+RT2m5gsCfRsSN7clGw+iMLmKmLuDuzXNj+aL7xu
wbkCGtqvA6abSBiq2ITzmSsP8PSHti1DU76wYKzayqmZt7ByzOwYdwva4GnweXzCA3LNZPYUE8xn
K3A4IMXJZcma28kqEKWzEsPqCM7nnVXYZgP5SFy+ltdl0t9ZzrMD29atlgDNWDa4F9FS73hIAaay
zmhyY5bPOyEMM9UDnF51js04EhScUuTJ8+drZ9zAki3Zeb3/diG+C9PyMbk8l6VU0S6pq/0+IBRP
Uic3tMyhGmAAN4q40jm6ti3UeIau/9iATzuI0SXotE4T62i1Qqk/dugZycN+cLMXUX4ULUFqvq+W
ymykzK3PnWktH3dyD6u7SMYkta9+9yHjgvkFGfVE1fIAzrBJQ0yUQcTvnwbTojeTWaCgnzhZr2lQ
Pm+71cnWAVgnnMpNUEHI8KCzomtfMwUVqXLmBENM8JqfaekVpGnrYhtowUbmo3wvVs/SBZuy3yMm
/qTxfc0sCzPC7I5/6aTvlsyAdeYIPBTj1xp4aB9xZQrAf9nx9Y5D4jSdTLrtkmDq0nF8IvcvBis6
8R7mCGIv8pi3vPg4Iqpihrc1rNwLv46yG5ctxbKED5WSBuQ905oVsUDRiAICzl64OrRAqwIcLaH1
ZyPmzzLXPovrxqBIHy2cB0/NtXWVSnVwPG6M+zckYwEFtsgrD8U+ZwpL1qOogcFRvng/v5xpQRy1
EuqkqO2h4Q9gMlqtbR2EMC2jPPhiBV9pnRVxhpOfB6QsSjG55iFC56rmhHqQMXf97dwjxebwCdMr
EjcbnjWpjnr+z87tSt0OF0jg3HhwJY5vt/wUbZzZAzge/CynEbZZ+27KA7nYF9f93IflHjboZIYI
cfzlqcWDvPffhQ3Eayz9vl1UosrwsddxuqmA3aoY/A5sKOAHEi4d2b5K4tqRcp/PiDi7Hn0oucvw
0h2Hqz0TE3sX4xcrDSHt5V1Y+dnGQkghquBxhiJYx4pgg8DQEFnqNCIs8Ic+1Tj8wbnGv+nyZuiU
Dgl0a4QUcdJEbyrXl1Rpq8vw3tWehdkeDvpyegStGr+7HblJfpN1mL6Ti6yTbQ3HYXfoGt9rw3SR
RgowCoMzwf8At5qLnC1RaeNfOq0X8Y68umVd9IQlyjUIrJStJRYYGjSrCQYq7LpjFaq9Gp/j+EOl
/3UvQFymjmh81WqLT28AFAx+sHvceSaVsy8Gncs1TqoA1hsk2ppxNikb64V8rwNBKa05/1quxPk/
hErmcV8prxIK9qEq4Z90QQgCYyWCd9d0MkjYEfUd0mvBekb4/6yflHdTBdYC54dYVuamDTkj4U3d
7n0xHfxoEi5Q6xKgXm2ca2CVBxSTdbpa99SPXphqOUziVbVL7MQkREu6q841uG2fHwnIrZRBLmQd
7x9z9F23N6u9nNfcSdgyIJfxgRG1pR8Qh9+H9hhulG5fmevXOqUl1cHZX5WDrYjYdkeNmtgmFOvm
tmYQ+Xqh0OWAU5XufUVpowmb4iHP9M8fu33fHOuIkz9rIkwihlTawzCrvhjjfBuZJJ6QW3EY6iBf
B2RHnx1LOT5O3z4HbeMnWiVZluKo6mJbAho2eZDpNsTp2CMkxbpUTqWNYqsQ9T4XZznVob1ETo6f
JeX5j7VgGxztPSEUFam/7WCgb7eHnyEPBLkBjMrNvwOXdCAEKFRBIyM7IqRDLX3O9tKPGGSJojYW
nkmk9NvC+PIq8sWrANWZOl0z6R9cqWTUcVBVOZ10KEIoCs3jTj2aVtF2Va22wkDXsixuUsPl8QUH
mlIzZ2ahtNNRSYUuHwIjpJlznBNoIzvOJIVmV8aAiojPOb+xrj/iMsiCTdBwsJdBqJRNHSQM3Pco
jQsPRaQFkUW8INmopUOh0iK7wyTWXy+5cXFbCYIl7anZ07nx80QQKnLPOT4lgEH7fmumToGDFY+K
WJezDb1LlnigtBQIAsmuX2CRz8d9xX/EjkvImKryVdFNyVpXajcRRtZjF/cls0+IR9r23uMZtxmQ
Jh8bkiZnE3MtopiU9VUlaIC9n1kFXrH8sPhH/Kkj1SpoEHHUsgNgHvCMTCo7JBWHi8W0JvcVUcT5
xqJaKXcvspPm6CMPUVGTuVgVOpAE8xdr6SNEo4q17KGyMic3kioxPR+36BeJR4BK/ANxbbGm/ZMT
t6ze64O0Pca8StHvkfwIFr2g1giOqfvvsZWGdmnyRKwya5o+YkvX62U/VZyMGsl6Q1fVFFgqbYyx
TVOVzDBK2taICMrmMwKm5lcYa7HdwuL2TlDwFcTBKy9wW0yWL7zeHNP3jZZZpHSLy7m0bV+AbJSH
crMUJtg3luwyppI8CfwBbWoBKy/K/DwpZruRERpRPhv0CyANR++mm2VtjwzmksFoP3JRcnKwlAHK
rwDZVXXfxGGn7M7/8IUZ/C24OQ4Hk66Pp9hWGQ9xWvMGQXexSeYOrbEdfJUtI5r0yty6JBdkdslP
kR3urj7kQOJWloNQdeNSzsFsePxQ6JWLhsAucvHhTE4A+suDlKlH7lJM8Qh5aBmJqjYUiWlq2Grw
wdTeWkPGk2Bp34PY3MOlo3gY7uESEFz8HLzVjKJqap4MJqSpXTWu1alcQHLI+KlYg3iw05pFoVsd
JKmyxR6z5K8u0CHthqASriN60H+RlXQJTUX647reZI/vX2hnABSMuhTQi2nE0jm661LZXyT+7ZNn
EJWBTg2fHQJhMNrEz6g/9lo6MbHi9igHkapv9V0xvA+HkKdfL7F+wQ3xI0jQCXUSxVKk8eOiutWZ
zNsoXoNuCjsso7/sGp5B0Sl5FQs6Rsx36RyMp+0ZuznDOks7qRUGyAjawyadoVS+D4S/PsSz/MMI
iCphuXE2Ybhmfg50zngO8pFWNn2Q4y0EIHl2dis5WUlvwx2cVIpl2nJBoMGKUssBMwiLUrzHS8/D
ygXFEJ7gklCHdgPjfJ/0VsaM9VGIgxZoOJm1ERT8X/v6ecMEPxAMVVzbp8hfHn2X/4xUIdm+VHiZ
vJHq0zLhywiBI1Ry+tPLr6HLb+i1NG38osSOsasduyxh08unpzWj3oMFwMfWhpJeJC6XJx6manBM
Jl3xEl6xNhOJoGNRCk4ypVDiwYlvkx0SIL3OmsgzKzlyEdEjUvBYNAcAtAOcSGZpjsXh5CuDxPuc
rodlT87bgPhoJ58MWpAcZwpUQOhlaNKJGFZh9MXB28qazHYC6lBM43zzoRbBeFxGLLVW8lS9TkLs
c83AV29uRlJMA+KLFR07NdOt35TcO6/LWwUquepPtrToNbwazToB+Qn2KoJRGqXgcrTwYuiSZ0uY
zUK2kqxpbqyYayQm465L+6nXQxALmy8hZSkvhZjYQUxlAU+s/jaa97DZrFQ7WrvLqtHDATf7qcam
cGkQyQyJ8+ILT4Qsc1LF5yLABrtzdOzBvtsPLOzUa5+c3ag4dqE9Fr37a1z7TCn5VsvsvAP4BoGu
Olr3Q0/1sEKe+/g+wc71xxjijU8vqDgXf2JRu2txzjeb8NKnPHF+QhbNtxVUYCANshsuqFtyjCwl
CL76HMYsgkBdIrQBVmhh5VsvtAxa5XHnwdtcdlCw9AQK71W54PcpAUcnkKyd+ZIYGtA0N7/d2zwf
afFAm1++1cqNNHZuGc+x0QwSgfWqnYnJ/Dw572DE5Utj8XlmnLrp/NRhE7Wj3D4oHFFz8u7ZfXxo
JDTDqbpjFom7Xw3pZ4ME45vf4nxb9BCUTD+n7l9muCUyart/uBifRC/hIUyzDfYApd6jb0zIJPXN
jqbuSO+SvBQTxRJCM7konqEp5sYUBNNaBN3LlwVqTAalybwpVd0IxMRt+SB9HTt/b/g1C0fRw+LN
uLUul7/m24jotmFM0+NRudje7LgtnEPOFUOoupP31X3bjyMb2xMXFl1a21FIMGyq93cde1XeZNNI
pCKOUfYAwB8Ez995PtdQtoV4H/HE49vbyy3b4ZCt5T5BWcKmXwxF5mB5EQeZI5PvS0yKcWnQ1YOl
84NxOM0IpVj6A5XHJj25mD9dRpk1jCHVLiPbHb5MyWjIk9Ghr1stLdtizi4yGQfoMg+A9LTREJd5
nbUR0v6KVxUc+qR0B8epDyf25RvVx7xoic1pqLtn88ghpHmauMdZmBvdjwfdA1JIrK6t60uB628h
EWL9aI/OZrBbrxqhYSkAIwvowZNufWgyS2UE+BHhVVyfOEMiCtb9K0UkDHaVPzMhqUs9b0cXGBDW
5YRTRGXysSdTO6Ly8+z5vHzdbsClyfw2zGwaNf4BX0RzAroEIvkS89wdCmblECQzHqmyhN1U85Ia
5F/Nzc/0/RkPo2sn8g5QwzPeFvftbXYbTCO9upSD1v0RILuor6AzI4+lJKjY2/Zi88jgjcS4CFZW
ZLATMutJ+LYLSNQuVNefHjhwxSHjadOwWdzk72n9MqYZDGErqrsEa4Pt8jtwxU6tuIfW/2gL4hpO
KW6F2HuFU10C/Lof1trRduoD4D9NiYoRr4lqiEOcPO1FyD0O/OS5REcIsL9FxPQFdszv7oO6eNDE
OAnhMO4zD5nj2WXjIYonTviqN9SNMiqisB9l6ZVFW011X6rE6u3vofTpzXA7kPFu2vcyoNQk+2fN
pt+jQJ9g2WfncZ5d288NoDGL6fO3ZAivwXBJOOysUA2RQISEV7gUhiENWB9E8S+PLzS4BbehhmCr
bMFZxHBZgUUhHfJr5a6o3LafRQZZS8zw+yMCcxAhYJ8uUzhWAbunPqQ10sEEq1csSVNrTZ4IEN+6
gQD5JX4NJtmxHCSK4nqVMqDRFrOjA/KrQ7bg0hdslnfdQ/RXRePUR1h27jfEirRPYBiovQ2L04SS
ZUyA10gKZ4zbWZ9tpKvejEvOVETcCjkhZ5zjC5PqWlGVCnRCV+p6a8+pxHll0z+nC1w3TT7ImNjS
AJ49mu30vHu9LAWJQPVOpI8z4jlKxRVwQqaO+qCNEAEjapRtbq0M6xnSu2iYfRt+3pRtNcRajFpW
P4lLESXX45PLPfQZqTbIIA0LtnxNv3WYzKffSPV1g27jHB9dJaocVJjlFbRo5no+9VMHcEBJ+eqj
Bi7sp3K28q2SY5fgzn1hLZv6+y8J8nDBDhCdK9/NAee7dE/3xbHi+C00LdjcFgoS19EEko7yJ9jU
yWyljCssaIOdG5h/SSbgqwpLzoNe8/o+Vm2QsX9DqdGbD5vWOZCsDRh7c23GhBVLk09CxEW3FFH+
p623rexPlsp2LeS5JaMpneO7aQ4DqsQnaA8Yn+WHnmZhNoqtp5a3Hruoeri1F6BPuAS2ZqOvucLB
awlUoaCwRCigdWtc3mtyH9BJGq2RzjiBIWbFap6h4AHDyCG7wcNqsuf3fDKbWBRgcMJdtufFTUKo
NYcjJsLCWw4tDb5IELii+t+Ysp0CR/EdcC7QqJOLORDQTlMUvBPbV1jss1MoilpBEK+udAiD6fcc
iELMVcgSvTl9KpnlW/xnfrBMW8ipSsgxqCviMTVBjSzM+SP4eli+vQV9Zvds/pcsDV7fRunGXzeN
khbbVB/sRsYFiyaQ/NibBefVAndMVnHNabjRfoBt84rSI364A1dnUm2XnPGZFrMFOXsLTaTU/I10
+78fKCsa17d/v/raXbJAQ3Sy/AL1sPMXrV/I9G71sGhRTO0FNKY0wbS07q/L5ro8clIDoEsuTXF+
sJ5kS6n7tieXCOcA60r+xklOmO8Xr/pCO6KfLruqX0Y1Un3TL8B/jLs7bPkHhDoz+4IZbf2IQeWT
dVpJzXlZaX0/qUkheIxV/BNn6dR0OhFYQAaKwm7yK9MsCxECHHn4GnR/Vk4jme6fhNwflcnzlFU9
6mUJvSoZaSt/oeoeAgy1xv6cmo1xEbF8lSwOcIqHBBTxTIo2k4bm3YfpBWYX2/g3wKECqLjrsWWl
JH0qQAFv+G1TfCc/GKEQwsIh07o/dPoLfgLKqdUlLUFf2rjgcx2gZokx9VCW/dFupWju1AfukOqz
wlFvNNr/R3lPw16y+1qjr3yzG4d7Pyf6CQ7s4RGaKhRnWShN8O3l7G/hKeFiryolpGc2bV0GQRqq
rhWYygoX4kBnRcZSZ2ju4Fan6yK3RrNGYeEcg9b7dtL3MbEzFHEU8AU9vg9nhDGvt5Ks5gkHnPrn
I15WKbp9/2WymTUKPJdbvuUB4CdpN/OyeksEnO8KhWXAm9k4ePj1KCk7g6kLI3H/RmgTNOKO/dYt
dip7vlN4PLmoQgj+78yGR9UxgXu7Epy9KwK5rLOu64VRuvTKUQwHdk6pN8zwQzPV/wao4NXIPpRy
meB1lSODpLW04gAly+OGC47+G4ZOaZImOagj2XfiMrk7V208AIXO6d0sT2aW/yYXsqPqsVpchSSz
g5A7sfJVNO+8zCKIqygg4Pxggev1z7urhGM9fKOCV86w4QS1Oe6u8lRQKFUU2EKlbb7Z/mjawDdS
8h5U0/a6U9zvFpME0YVaqWifSzWBMiFZqnKWCghgBi9Ld/rlFCagFvE3F9ZIn17ogeCjzAKe2aYY
nTdLqzIUmeb/7tD/Ec14Bzo0iW3oeWo7nwp4fa/e3phC8UgQyjOBkV2tBcFxhGHZpkfb6f6OhAs8
mx/GqHM/B/SNbHDTGYYxnxK83DX7F5nfe/upBhtNdOOF1YWVTkYcaD9QqOmHWozjX4aZNn79SN4q
6zhMvrubC1X/WQnOXrjqTCBPmICko4bfxAtLJvy1Vn2mmfFI1CV/lUNyEFcVAPN88893lpTx2Eq+
D2AC7fs+dWXVBJxtFHKkezkfMKb9UxlPy3Pvq68qRUG2BapOyv7aocz/Z2uW/qR7Ia2172exaBIx
7RrqNV5zT0D817XD1vhoeH+IseW8Bm3iSAMaLFbPHLEAe73s73OnKQaG9Pi2jNpgukdfbk58n3YV
GrtVt0JxXIHIwjFAGS2at/ZmICAyEV2Y6No8T78prSSKW5KGaVNUSTrlloQvlneX016o/3NFhSaJ
SgadWMxxha1uPupKkNplPCQKsLdZaHAT074l8aLNCKV6obExf1Qu+0aCzb0G8287QeT7z5E4kKJZ
J/u5vVU5eIeqJf5t7f53i7rZr19F1BrKNTjHej0FDTk9BFe61+0myJvtv1ur8AQJJOtqDQwp/HKE
FvP4L/5Hzzm8E5pQcZOkhHENlkpz4K3RKvi3oKBHIN+m29fYU39SU7XQkWBvddEFRy/N3pXghSrb
sRmM4VReOV+AweB+XlPwPXA/4e+ueZlUIXpLUslWEWdB/wvoYr1a5e8kRMphcAXR33nMSsWZPTJs
8FniO+IxQlFu2GmEHT7j8Kz5iVf4X2Gte+YeMX7nz9+U+8cN09tjhzHrLPKMuigqA1bBjhvCnX7x
P3gJ/kl2ytbs7YPP4WFCehy3FWEZkhrjWX8sYrHoAMM+Q20zi2xS+52j9Y2HqumK8lfTCQVwN5JE
oDjsxUJUny9gO34XBSRJEHvycEnYm4Ys/LFGk9Pcb8v0BTrXZkm9InMVKuyDFYQTQdNVnO5WrmHQ
Tx82wCw3epTVysyLlgdXfl3nJBtLHKdpvRS8O+cmZ3bgQGGwmSXJ9ZtXNgsHu9Ovg6XMLtbsp6Sh
qe5DaMOWokfL9Lc7BXy4/wHtj7RkkHQnjQN6atImcjqbTgQv2V5RXl+0sh09G/WtUzI0Je8ZLaxT
GMUbNFoGKqkp7nQxLszq5ly+e/rKfSosJqL7f59v4moYXR/FMWjL1gtVASXrabeyZvbKxtS+dpye
hpb42dd3JsiUSK1fm6dkuA/i9On9YFxvsSG+UyGZjnrtZNrHg2x4ZAw5hB9cEGUh9Fzj5wEKwhpY
gxYuyG2vHmVN73VCAGotcHztwClrd7NMKRt5yvl4mr1gVoCbNmXIwkwrd8AWBFcgNUlIdi7+4KSl
n1TlUKasgXGHlS6ypQoS0YXRK4EPnaXE/NS5GYf5QAy5px4Yu98lTXL99E3v1t/ghAfwQVDWoqEJ
touWysXA6S9MhmZYKg+imq5/UsWvQSxFuAGylpDbGooDT8StciAjiguxqw5/M2CpEN60soqRVCAV
uuHDGG6iyGBot6emhrynS/j3k90RJZuVc4zplHAnahqXNJawiqJI5CAzFoFha4yz5EqFbSfQOza5
vawqH+t4f8g1hOaZZzaMGj3stcEZPLmLS1VWbMlGB552ej3a3kBhWIUc4zYp4nJYC/+uJg2UtRm/
HBC3/AZPkz6yKnLb1coFUZ2rnVNZ0Vklr1buAAgcS5eyDxJXKO4c9FY2Rg0lfZo2YAH1Evv62arF
bbg16P7CwvzKvSdYyv0m1yUJ0GEf+PZ6nZqI1LFhFTMGfT+V1bAPM3WwbAQLwRiIVRxv7LHx4/pd
PtBYt3L2VdPhogc0naYOBLWcEgFZsWvpK7wotR7Eo0ZQWQUkCp74UitGkyEH7uongPJjY64Q9PYf
EVi+9+fFtaC4RQtcA6NzDYO09Tayh/x1PhERLIjchrS//s2vHJtk/tu4w4qXtOC5DW9OhffImQit
c5nUvGYuRbUOJCW/seqsF6gnifFjjK2vZVPONiKJnPjs7O2IW+NBgOJNBSTFsdPOlhZnww3XeHe8
ilHALcXQs6KCG+y+MAfqKxy7JifFSnGchBWD+xkr6pkN+pQSUmdyDL2CqLSDMqzAjj9BLw4/lLxw
sBWAB7NC7rVxZdAXDpkZvg4Muvge6ZDJGJiCR0EIRiviTGA6bi3IZKjLKUt5//I6e85mWPuXL83J
gZrBOIHm/eByAdfXskXFCCFM2+SF2ptoiDokgs4E1PGWntQtEkqmNigUikJZl/qthbWL1Rs0Nwk3
PgAokmrQeZQq/biyivFjQyyFzqMA4qmcSIShco7QgGWGkzV5s6ifLo0hs6aDG2dqx1N4xi8uZH02
ANVtFjFxUDn9SdayYsKjmF5UpQrl13UAPcT1rt1YOcuslyjf0V1W268njwCn8TcYSRHdXuhIpRX5
rAUyru5hOLfZDwVb3qaQZIFtOVYat0y5z2Hf9RZxNoYeN9CqZNXaGNYWl9AMa7StPvdL1mCA89G/
fNINrDBYWTH7YNB617kNVnALrH606bhts3oXPK9KbBzvN1th1FhQrsWMmz+29KLlKRM2Btb8v/uv
Le2ksOtHtn63b7N6321YabOyWVDZOcufVd2Y1xyrH3bjtOegekJw+tquZxiXzdeKVKdTzP6utNFr
pJpgeBabHxkmp0FTcATBYafXdpIg6eDjpFJLEe/8v/1cGj5VjhrJ3ayeeccr5yhAH78lNBUKTWv2
vfuUzY/I3uUcGdwUhgesFdtobSUGCkgusBoUGlVYtgfj+Fwlfe4Mx1ZjQnXJ3uTll0UBjFdxXEPI
/h5fQBA7jKSwhkwWl777pt8bwh2CLurrQpfvxvZErUo/K47eE1WhlMBTwLggkGD8faf2Y1i8x/rz
4X///hVgXpaq1d7OezmFb6jLKp68ouB4DgfXH+375jz0eNdK+Csd07IMqdkboXX3BFQkWkQQr2v7
AHv181YF1Fuc2LD3Dpmp566luIyLlETND4idmZvvqlqbY/qOAFCRRVmYoxWZUEEACvL4jAhHa8Zc
HKR7coXjh67vawsw5Y1wRgmYO8azkbHpVj9yELSIxjuraveBm1hEZcErS/2SA1lHk9+Czw+fH2jD
zFmQMElCwqHnVNq6wStq4wGybwdHDEJMmUxIXDQucz6HjWsvFVZcN9jZFQETr/e/1WHg4sn73E2C
DEDr5RN0ji6+n+5Virm0ILFuJc7jld1NI2B2adkzZ6EvMRDHhP7Kt0IlQ9k8MSd7LeXKl2JArLmI
0fPxYqhTMCLJVI2RQSrS9gXvoLwgbS2mDCzFQFTpMb7jxmm+NlROJIBSFBkBUMCmRah+mu8/IaYi
xurg5Cb9+Gh1o8zOPZVsa9R3KF5/I9JF8N1yKBatQOD8w+P9U3n6d1OkNIRXPoxSHNszU7dAP8ui
QowI2vdBWHcB1rH2XukP1k08Mtzanh7HF/4zVEgteQANxxKeuYwBkSmBkQTSXe5iiVbdmbiMaNhS
ng7EvMKlNugJ4ZHjIlImfNf+O1DpKzwrr8BELw3fkXI3CRxZg0gbg48oxigZeAhKWoHcEh+r4BO8
mGutsGw+1IH8dGsqF7gaekP5teSIHQP825MHqwbGncVKpG9MermfqFfp2JE+CmzHigyS8tm75Hqk
qJ4eaU6VPzR9A58ztPRjFRKW+++x/6QkX7QjBviiGjtkF4tLtvvgJsmnhzUklGPXVYHnIeEQAucI
52kxd/Av5Tag79QGkvOkoZ0+LN4651RVljaRgzyEENwnsdAizomB5vbHzflNr8Tb+bUoZ4VcIAjt
jB2VlnQ+Ii3uL5PuR0sLAO9jtIZR6ka+Kq6gykMebj7ezau0PErl9D8TtxMYNhpUn4G4onGaYT2M
HHh7ecWWt8srErSXCE4HZ+rnVex2mErpa3Vd9RSUrkbHFFFfnofDGxIlx5NWQlzr+N6x9BWc60pH
1JqpTmjM97tACSUiAgmk1QZ9C8G8xTEUfnGZyxAderugASjZf7BFJoqigyWxfnmQIbWJYgCFBsgw
bXkwagNOje2PAIr7WQso1PNJj2rCqM0Lvtukq8uZrgrkRBFOtvuBW4TyrkX4BHZGt1d1uxzePsEd
OfhkaB3bTnDK4b0xGpLUx5Ib5FL5KdUFpnuhROi8Z/OXZ/C+JeGhRT7pfskwrSZ+11etWtTuWftv
J8hPWz6gdkdrBfcA1ODznMreKqShWv5ac/4SAePuJFRCDOdf8MGntzKiutBCwcig/xjL3aVKDtX9
kXdLCmuyG6Y5gpEtL5X6tY7yeq9Hezw32nn1gJHLfk6++dXc5NFzmFqt64fX+EpRJX+pbTKSk6eE
WWC/dmmDARN/vC0gyTUjNlZmH8EZ556AvlyHuTgxZVU2WXDyzYFk779+xFy/tdzN5AoLMM4ORRjp
0OMjOeYcdOeNYlhnQ2iHuGwXdVuUa8/bvh6ttP859eZsLZmq5p6ojpT8U1X4Wpkjz/xZuJBGrYfe
vkxQUohjV/g7SpeXd6sdiAz0LoIOOXjFxRx6ZkCogp9mFCDIwFP+7MSWq8ad9RxjL1a691ugNNaJ
23iFzP13PR2SnPvnJN3f8oCktY5cUGxEGB4VcC4f4sLcJKnvdZeMC++LybexHfQVeBB7fwlt2GX1
WleNA8wuDiAKjjqNKHv4BCOlGDhIS7s6j4GSyfvw6b1uR+JFLZZrBLkNDJfDwi7lLbgD9Ioq7G3S
1e3o6JSDuEl+57xXP84XhusdajrT99QhPryeg/4cIaDNJB0M+boBizM2OEyCZsKslnEnLSj6zVqK
p5YfWGpovG9DYTANXiZ5kt8SET7NT1wvd/bdV62ZPIqr/PquJdiHtRT9i5fRMusdzVl+ghzQ0Zke
LTulb2PBYNzLRkirhRie5NjUPKpgi75gACelCQYmLaJ9oAI7+loaQwZv0Uiztr7QuM7wpm6Nbwfl
2A/+4/NBuoAkPbzkvfH+4D77alBTAtOxLM3utL1YniM+RsTBBNEds2QisWUHizKVB9N6cEBCe7DF
76uIDGSpi90yGtLccKjYty8yggrzrg6kKX7coS4S+VWY6Q4sq3i7dkuD98G20goHWXpPdE6Qjc7m
Ds5aZMGfXAJSUE3mgiNQGthXw9ohFzCOH3TUttR0XbsOUvc4Jqae4ZwmdGubIPndgnP7KHHoD67J
IzZ5TX74BqMKnMwqxe+zSbDLkY4KBwwYQYkRJxeO8/Tj6i156p1e9gN+WStbuhQW4JqZHpUtBHNn
C8byZOFe7ZQn8NQjgA/z733mjVIwpPj5wntnzeuF5h/w9Iz8DwQfJCzBz2iVMvY1gB+gid5WRKBH
jDdz4rR4Jbeeq4YG5D4hSO2XxhCSJmZP8VaJ6l0azea3cNUsWVNkckI1TtLY0aQUFy6DyH8fuytR
2WP48PID3eQzzI2+U4Pzy6wJj8LDS/MkFLg/ZwMMZGAbQfSX0Nq48NdzdLQCi4BOYJ+TQ/mBoCIP
nmHyTYCS7XEqi9CNbSGI1DaG9zoPeMNIN9MduqqFt2UjH4ugV803uaR52rA68m5gvOLDOtdunF5b
kt420L1JW8Jyt5WHwaD05gBJ6TDGCot2gcEd42EmOfsvR87sv4N2SnVazJAQ00RNjVuyy470B8yt
vwa+Knh1SimuiKUiXz7uv0Vci2nlvvJrfxqXCdMRUvo4gOm8pmAkcpXDmwI9YYbO3omnMoht6EjB
9KU9XbclFMuRp4CzdiHZYQsb9FlQV2XnoZJGgZApAhNIjPQidvrD904gliwup4S4Uej+y2dEWBys
BWqmanziJzRYwY+GS/ZzFtJLy93zf9EJABlql/RsQ61VqSvJ7e9pVZIawDUCC3pLFMzjtC+VSow6
+AbcZfnwtptBfYKq+CuykIbSBaaLKBYsO3pelRQZug2JW3TZj7DLn4ViZerDsmJcoYKOJT5XmHZL
9SVyqoFMEDMh35U3FJyLPYy1KANF77lAayuDBgbQkc+X8IsMGila+x++bMtgh20QjNZvXy2VZyDE
dTtHrTV4SKGgodYYnBDljhjS/AZYRRs4hohel+uUSFRf+C1YFRKjJhrdxsHLBYk4nCKbR7LEozna
vxvmdW0lI6H/4UEzI8qQEZo+nRCkGzqt1JqnMixkQYBZTCMFLhok8yE/RVvAs3xossTkCIzYcBb9
D/GRapVKnvbIBR9vLEFezh88ZW/5+SaAZKm8h4oJ6DggjNe+7wLEWwSwPvNy18kpslUhpHC/xZD4
rKngnn4McD8TJNoZuUFJfygKv2cIOV728snQUL15JKTiDkItrjVKe6VL/w84bm9j/DwQX6Vyp/Pi
GVgXYzfkLldz7Nc6GusaJVBayrbUkLAhPXrR8MvaAdbnVZLNnBYa71ppYTsDqXy5l5yoJjJUyRZw
JSvUCSPB0EXGPMdh6iIEyInbGMkImJU3S8uVcRG8u6RvpC5c6GDxEQoKqDTbFYeUS8Y1ZDjhx2LV
XnUQ5cjAujfRhFhJ2SB52cTOSAC0z3C4+1l4hHXyIOufR5yTzIuj1tmm4sYafVQ80XRJ9ooX4ze9
xb3Riio9KKdLtY6YDGOHt7GE7yGwAm3XYDAwd6ZdArZZhxgKEDXFJ2Jotu3q73Rmejz93FQMOzM5
NTaSBy/HLfwS/U7xqC5L0pBLsB9W4i2aCY48r/8qMDj5+a1lOObkpZnqVsF+dxlL/Zq/q2gD1akr
Ru30ZTTo/JDXXgZKdmSQYeF1XRJMcmBrmGKrUocmvS4wKZoGVv8bN+FYv0IfFlgmsKZ6SU0+CpiK
jILYZRkpNCfGUOqxGZYc6B3Nu2L4XsC+tEUY5PLQpPhSEYNuY4zLvt1Twcw9d76jR+y0UKv+BNsg
WQUsF9UCmKlz+wwpl8Y0X2Y6fv1VEY/Tj6MiIMPlOkN1YpdziIDeiNJkipcm237JnFlsr0eSAbPE
33/WT/WOsQCf80bIdS0G0sEoS7Mtsqw5yg24tiBQOJqmcPhnxfe35JJWSUVZXM7RkhLxgTwymnGb
tXTx2m1Zzl4LMf34c1mRdCIZ129uFTkBy1stLqTeYXR9rZhkdbH5tnTKgBIeJmBw5Jn3oIomn5DE
NQg0mAtJ2gAgKt5KhBrp3E4lPpPl1Quk+lXAdsT3g3OZ4va9CuudqcOhmnT8xEhhIl45KFvIRGNw
Sh2nJ/msIuvtxgMxzpPSvItOmGt7I7AK3PECSyOfXl8cs5tN5rXO41xNITrQRxiWl1XDZ4HoRfAW
AwNhlbOLUc7dZu/rlmgKvv69jvQu/Zx/0aFJwuizHl/xxB+nmfppX2xKJ1V+663bOi8m5RMqGQm5
TMmVh+Jea75osldU5OeL3P4fDhCo8s9fKLGOVewpyv3TGSqQp1uZp6WOl4MQlct+0gXXX9pO2Owo
UzAAoeAwLSunDcdO5y+O4ysE//iEcs9NeBluhJT58b8bDsSMvfEmG+cJNTRV5IvK8FCIoRKV2LEm
GETd6hYkDlXsGxLg+Tl+UFD3D2TpSeHsC03tLyrHNiX79i0qCxkHysJUMETCRpn4BtOWam5D1UeV
xVpPGv2x67+UZEcNCTF/6YsOGRY3PASX2ybod+FY7D4Q4o2hVyGEJWgoQo3swEGBpnBhnd0Cz8KC
Y/RJFZuW/oEBnWixIK0eq9Jpt/o7pvl+86K9UgbNHSP5YCcUQ3LT6hTIIdM62pIoBXgC7Srd6dNM
QcfLHihFuXdzMwklHodFBrULk8SI6M/A+RZiewk281abP3zjUvD9PfBXBdisSeUymhZz+PH1IpHn
aq7kQmM16Phl4UP2JbokpPkIFdLYcQcPTDiMfnrk2o21k7Pl+ncx73pdvCO1O2jeJMiep9+JNDPV
oSZdyEilfpOab3Kcvpr7jvfMAWOR/QO4umXQl+MReoas15yirEM5Hhp4DvKJ6jkGhCixHDrAfA5z
vZAPsEnOBxcLqI4K68qpbiK1StEQNky2WP9vEV0RMd5KEuhs6I/MR4cA2m2oXNK31Ubj6+WW5gbX
XUZkjRfzEZJGKqpCUSMJ8GyFX1MwfRS8npALI0UQGsAeV5M/vaGIf47fNESVrIbLQ/GGc0hJkf2j
IjpLYAZKpcda6qtdrVkZgbAaCFC7jPqWH9FwGj3Zzroapey55jadCDZqIpDfVR4w/i5jiwbEdoki
/uIJ7GeVff9BGTkG1irkpcH1RnzszHOQg2APvli3xX7MvUqWsihXIXfkRLRVAjtGBJ7R5MRVxlYi
PhzdwwZrybW7SQu4OI4YYUj3LPHnC8U/6hKq/lCq42SakCihWbe6DZTL5Je+ZlmXJzVKqSKZhKTB
RiIHvafognaRwZId3qk8cSYlX7epcrwx58Mdb40U4ctYSDAKXa8YdZHI0JgCAkMyy5r/sHEjtqXT
8clXlRDq6nc6VwN018pl1nHpGpmNwwXu/l54GOsNttbRjPUHxjMpZvSxOagomR+htN4VIH9qLty2
GHLzPTe9nVSohB/YjjxoWsvnBjWOcpd6rQqR9wAtl6U44195gQHmyCFlhm29yOJrow/lQ+njQ3+5
SWDtA5+7JL7yWRxxUEm3rWdjrIjP7VlKiCccqoreUTmmkEYmDqYGYvy7RCOZq5tSBxFMD8JGXGOz
5LDZFWtthrMQwOKYUXw2gqlGx2LQiTS6MFHDMjyUw1xQJ/OzRRw0IpmkyNnmfMQ1rpScbfZ1kmUy
Ez5yv2giqBbqRGTtEuxuLS9szfaZmtEUBRELp2dO6AC/tFZAXkoDxB+NuAqfJYBRfiVF37S0Yk46
R4QLKQHEy3TtLHf2wrOJ5jx1cxgrDR4dUJOxyLMZg5xteMKszU/QgFpB36iFJ2eZ1KEidCV9bFmV
wKDhQufgYpr441x8Hrfvj+z3yafsuZHFoKGtXh7QaVvEDu4/lncxw4cADoEzkMm/RLJNX0MbkCNj
SnmyzZwNyRxwrXCcu/5Gvf/w5ftsPrlaCYa36J4Olj+o5cwzDSmXKuUAh5f8EYgAkJxReqFysfqr
lRau2Ep+6/6FV8m7UdJrUYoF1NI8gqMQi/LYR9dmImwcjWosXlAaKkes0cxS4A7G1W026IOZ2coo
A64qWr19kI6M/4f3MqrTpjS/jzNwyvpEoWxC7GbzUs2C/HoFo32vebsqwcJ3xujtDbVL5vuuiCoS
/tfLQT3yqmzODtF+TVkPfUwAkMLjjljNraSXZtoKy9pQW7bJe7SLPHVwtbuiAk9yBaswvK544uxX
0N5aN1zHd7SqpIMbp4XDnPrKjo1d862BZjy0qsgY9bYp0SFw0qucUcUpXe0iWungYjY2zyWJAZTI
QQF98/n0Ahx8ofj0GuWY2roV6pDSKtNJFZE3ybwM6F0XLb5t7Gb/Ou0Z2dZCaii7FfnB5BIeFlZI
EzVrC9ZbnrQ4+SDteBYvCIsN0W4eont+pDRv9X25vI5xXsALBEcElaMt+3KMxBgkGTF+YtUoN8Oo
95R/8tQK79hMrEc4k6qREtVFbAnNo8X/Dd9pXQ5n9cd1uddzB1z+KfK9cbVjIoZbp0EpRauH/3Ud
f/Bz5beysUdVIp7xbGQE5r+XpsJd/J7c2ySfnN/W3n7JHzjMtSF/gekcDhuxXnAqCTaM1bojfW1q
IaAI/sj1WJH4JUp6NjF+ykaQfIc0cuFne4hu/O5HPuA94wTRWJ6mA/kYJhFt/RrQhI+NVUw4BHGC
MfStRfeSpXIO2FFlck6C6RIPRj5lISfrHMNYYYEBS+TI8arR33SaHN4nrS4wBQ4Gj3c3A+42sxZi
umNkcXuR8yA5aYRmkE/Y64stx0lO5mbet+9mJXIJF184RyCuvc79vGQ4CdXO1q+O2zVhcM0me8+K
Cwvpsrbgeyy7MO9VPEpAer55cIztB3UEpyiKobKRMa4GS9FZWjd7Qc2sHmLSniJXut7UGWw02CCD
/d/qVETEHziW+LdrwdP3NGHP2AYaKOQJQM7jrhShTcerxZS8069plL7ZmQGDRBg8jBfPxBbLSnFr
ydO37Jo2tFyMdQ4khxrl+CgZJdK1oCBtu1Wqq4W5hJa4R9LDpfzfIgkFt3BlxITDGVVDGKCvLV1C
Zko7QHdMlrRA/+V31s6Vft/RQBWnIy+PyfI15hK/4jVUyaCXTaBhx93te6Leu4IhNju1F5mbSx2B
1S2BCdm/zpZgZneAxxPvattmUc0DuQLNST1NhjSV7n5WY5UGUOtNv3iz6S7OAJ3zMebB+r9LrjUi
TByA8KbLTGA3gu9I/UjblUt4zvqVAYQ63P9d1q1E6NHX5Ak3rlsfEiJe9hP0mXqev57EOkHCIUZI
H7NZz1uS+Har8YAWA5qB82HHOSOxoTZiyPpZXDv55QaD7vGuoDMl3u13r8Djv4DsRh4o50rKEO9e
1iRQQzbs+dnzbnFdbNf3sVLoVgS4PiDnmSmICK9t3JD0vosj59WxRnxPVlhfhDORwuhOECYcTqsG
V1GhYuF2Qw5PXaABpM2BapYEyUEdnmFxpd95/YxpViwlQpY+lPHMWOvTsH78Y1ld0ymjd86fOyuV
7J746MUZJkUnTCOGeF5Txa/aLIWsqUPhAewKsQ3YV+bLUSwDtEhPzWQX5N2X+zvk79eekn2xsGZP
xb4PiaTAHEhSQ8LIShA/EX7lefTn8wXLClwjJFCEYSoR32BDCEZKe9IVaVtThSlZl2BThV775SoQ
rQvQsUoE9+Q0YY5589ygW6HAn/PxlsSGmhfzKuBT5a7ZeRDYVu/D9VmMrPXQ478jGrtJELG4j5An
aqSpkUbgaPtMX2M336cEtg20NR87dSqUJm6aFSUZfUyohLQQ7xo9FU37KFuerG0u9ErvCW+GR1o7
caIqhTTtMayo2W4zIzKx2+FGv55XCXJnls8tTZGwL23piouKHHN+jagIg6EH8kDX+okWQhlR6FKY
Yv49BoHS/U1LYGYw3FMEMLZmPo090mGa9fEP/nU0dC7apXL53R1B8VyU7xoTpujMvd0eEAGbWJfQ
BQs+3x9LV2IW0xKxp8MtQGabbJ2NJk5R1jwcaMmEZCHutiyEXZyQ/6xEmHSA//v4cyDZr1jK31YN
DsPgpz9NMNcM4H/6CkRsCj8lm/0t+cWMjmBPutv8aSBnE7ORDBiDy1mlXQIaWJI1qOYQNPYyBe7G
imuww44pOZQyHaCwHqCQIweFci0rI9BwGUNXpkftYSYVjCdBThVkqaa2Bs0cMiydvipRsKA+eM1E
6HJuMZ4ljtty7uUsxqS9Tb/c1a57BrMvuWi6wD/sqXB9a7WqrUzyNVTgUbwomi1QtApzojx7NHa1
zjJuXHFMKgxYgMyXnPyA+gf62yss61QcKISQ+K8L/oUbnmHcFJ6v/TZFAa9fS33Y8ViZoM42cU5Y
zPrR/8+gsXZT4MnyrVrqh6CqFDmFCnYWFdI/HBHbIDIA1sBgfup6NF2BIHu5X9Oeq2AO0GHbTu/p
qZdrNgGyqouJvBeMto9/9rkAadzCCwCqQh6xncoOOu+JVIOV8HbkTrz7QB87cwSmEfVgSiRg5fcI
a7NrWr6jYmPBwIai7MdmmbFE2ivJ7mN8mH3RcYSQbras1Nm3PqGjgcg6Z9rvC8dDwy3dk/jJ6M6o
ih1MfN+/V1gYTq/m0A27BJoUsQbpPqSRSrR4r2CB1KQ9Et6vI/LBfCFoIgPHBcqjAUDGlHdwiuWH
5pRIxP3hwsyB4Du18ejM8NuQdT12MvcvT/V2+4dyeu08piOMmCPmskZAcZ2qRSwiv1nfVu1UGGQ4
5G2VFNtNS/7QlchFSSdpTZykhqGnK+pZPtGkqyZB4adPUqBitGMwkQm0X03GXDl5644z1VAyMTsB
B4lgOswwe9X4w+knPs6SODNzwYmQo1WClH6Mnfg9Q+e13Xa9yFtYKXhanoVMvDNx7nWNVwAzEYqX
9jbXL6yaya3J1hjKmN68ByQCZRg10UzwMQfYSoTCsnv8pcDxSnfUt9JnhU53xOez3bPO3BDEEuA6
m+KbRvq1gzCXlB33f/M97foiM30H7MkWTmSksGnCXFystb9f+8dRKVfVXpC/faazdKnjzMk/SXCE
nMn+rzD9tlDv7jI+8r+IbfrjWdi+2i8QFN/5JIbSCN47Z2+EJWMwTrPDeyBFR4mj/Yj2yxaCzrGK
LqbX6YJtwqI5Ka/x5nTPlh0dDZEZmfl3DJdZX4BwcCtj+9F5CBg1fRF9YGv4TFBSELpp1Vgxm01J
sBiDuflSpFS7k/4Qw2ArVEt5/9Q48dfuvCmZo8F3WFJU6jGbFCVawUs0dm+5Iu1kzGUmxdcAYYoX
xGpA75cb6Ctv7BKLIZvMQBx48cmEFIBkQQ1bvdmJEFtUHZe0s8BZx7JKYeIPicgLpWajYCMAIHs1
x10TtKS3IsehjGPoyvleVwiX6cHnSO95nz+3ZZhOoK72k/0pDPRZHoW10OP+Mpfaali9KlkqF2TN
JzzF/q3HJo7yjWGgSn92UXZvP5Gu9Ck1WOTk1rzK1z9QkA9hQtTDL99tDmM7omZbSbX9TtEVIApS
93RsYT0KnzdHo1JAPSw3GZX4xjq0vFkjfpuoP/NBTUWMaspLt47KedVJBH9RPqjvxXj3BxDqUbpa
0NfC6h7yr82K5Rf4gPO7IEjYB/pW/YAgghALlRDLTF8kylQyMYQ9T/zf2WMxntjzON66cBWWkJAl
DZa/QSUv6nqom7zw2gpeyqwpOFyWFfU+f4+VMSo/tNQJTYjvYSnnDtcKyy3m02FRLNR5zlSLscAh
m51cd/4iyxNEVu7ZhOh0C9jmcXm9sSt+3CJX76PrcnWnjgvupXMMnx6JoWGoWai+nHLQvi1t93g2
GzUaGmOnrQf7xvbzVeliuELhMAQUoG/fV29l7YRWm7m2dXiCKtvLOyw/Q4AcBdM7rQ4a2kZ/zC6y
GBiveEmiV3w1urYESzhmOPPuHRHhqzRCKgxpizLx3oQi+pFfVgWgEEEJw/aJV2d41pQQdFYRxxcN
cNDCg2eQON4ROrXR4CYQqN3gDra+C+HkeEZh87vcd0NOsTKGPXI44WlMCoAiTRKne4jYrTJQ6jJQ
nnNNYTIX1mjGFabeVl3YvswM77/fzQEe9GhXw4LpWq5BO9Do+lYORozp6Dji0uJUTFl0FxLXvtb5
NWlVNI1xoxOByYOUxR6LOh9e6vhPkyoEXvuuQHMS4Xqwg32h4aZestLGmiJB7jEjHPFh35jzNRtT
M4vgs71e7P5VyR15rVv30EShfefrpokGZwwYUDWmWo2NBosZkxf0kt801Ra0tziClEaBlKYuvYY0
ABveMZKs965zagOWLpeNNbguTpn+XGN0rCzNL+qvenamyZOpnIHUJ8HWgHzxe1wQiZV/K3KsBOY+
CnxGk94vQlgzk/DQOYR4JjIr1qs24mkxKe0aeB/3HTuLQNP3a5OvwqdHYvYL5v5SM6OI7vYEZCXy
afTT7pwbKnNv5bZLCz4hs/kxB8BNY/iSCJFHHwlWvZ4veJ7PbjgO0fGCzjg7nKxyyqnwOce/zyXN
gAoiy6dMTzuxGrfcUfdVHsEcYbsxL/K8ewwQBtih9YUI7/yJ52ZB0y7399T2U1Sd3vt39dUTzV8G
MbY5k3ri7moJsZyJKEZo4bvdK7Pzb6G3IKF+Bh/TpxHxLqKy2SrluOAKUwAfPHXtwW9osCwBV4iK
Uej9sQdwmylYGV4lw1ZVaikyJCn/FsoIpQTC/Yovq0nLxMrXHPrhDkrR3uItx/H4Dmuo4oGvPmjO
Ib8ATS47uh3DNjDlem2j8tExysUgL7QgGqz8PjmkUNr9572UmRd/k+elY7xS5MRE+njbW1Hzor3g
FphFZ2FPNde9znPdDM4GBsj316H6xYpvLrUhsvrD/XAwdG+DOivrS8zL/yLRYqd9F8JB+AZWyItX
8UIhGTIEvxjeYk93t8H53B6B0n65b9CNoSU3646+NcsalBGlErxt5Atqq6e3G4qlOf/AEt78WN1K
/hEfbi8rxekk25Z88/U26rocE2QS5Dsu6XxYsEBVBYcGrmokSYQGCEuBarHrzKEF6j40iofxoP0o
pBwLQC/k3tJ2eobzXyoiy/Z3LG/tb8Uc+5G16HQyPDZ7F0NI0TsKxFtV7E04/5mn2JdTLyHpLrvZ
bPGSwVXHxNPf3EseBiJxRggoTZ0oCH2PsyDGG3zvWLvVpCfGO15xPyQnaVGdoGpQXFrqV48Idbm5
QEGKaA9ggjXUK35Ja7ruasmdAoCG+iDOfrMdrkIWuspv4yf7ySp8ymLV6k2x2pVtTjyJftUL6h0L
m9E8VoUjCw0RWOM9EQcqe7XE83CA9i/ocRxQaFh23GTXKwPza0Rp9dU3xBLCC/U/4tgkBg9pMQYt
/Fvflxyv6V/FbqjlCkb5uXlGbA9oSBcXZ4Tq5fNY4RMuIXO4j3ngie5WlvPkpU9wecr1ck0k8TOE
NKiSqZckvfTrNikxAGdft1Ig7vT8oj9JmaoZJghOYxlNJUVFZdd7NI+Y4niRfIwNdnDpLcoaE7HN
iZoLKc22KHFI1BkzyW+nY9I5Skp4Za6LvlrtDCJihx9IEg0NlDyFGo3r6eD/ZslUSfCx3oq7srxA
6H60yK0G5c4W3xjl2cTBN4snBYYoFHKSjzTdFWezst6wC5ZxoA4VO3/1G0MLH0BIm8ckMGdPBtD/
cjmmCQQnlufCjI7r5TO+55B4pECeVLFZnH/rwKNevbULVdFhcx4K+DVi+ilbdhOQooihtU01LpWQ
+sf1dRhQ/wPi9fHJWPNBeYXFfmFIWdmSeDzpVdIUTugaFbQaQkzakNRoZugYcZVPe65aixefO6+R
SKva6SnAu+0dMP1zDz7lri+XZVzPDaMPyaxVfXf7nMWeuXj1Ilw1lvfUdzqmVKmcfh9r8Um88yml
Sdu4+uNB5MXjHXYzY9BYe1cFMlRKSvjj9CSsGNZ120A9sP7flsC4YmytRLr8QqkYtULr98Hk+5Iy
sTJ4za9Xv/ZNfBnn1z8XejlQbo4wV4falB9ruX4V/wNymsJrWEGdiiMIFFFzh4fTJsfw/YAGq2lf
dy2EEy2Ey0GAhT3TWzL9kNH+rcFCk+eLbmjy/y3OTYyUoiV1FV1OLADO/5Hwpy0fwuz0zEjoXF2e
q7da5Bj8dKBtgx+E0MnRf16se/zuAyLIu6LSNNHxSc/KSnRr4ddzMJsICydCAAdnYyR5yZW/eZ5j
BrlNAn62YOWgPcTFho7s7+KM8SijI3lkWvVymUTyu+HqmVzblLkLVBzNd1nYHpTfvZK8zyxWDJOg
yLQwAGiZtGYvOfTxL/ltzFTiVWTdBlmodcwfG86EQcDEit2tYbUqW9TxY/ZrKWXTFE1WMwzmqbfA
DueO4MeDQSTRSTDPwYym2LNkycqxy3Sl7zRnaT0zbDAuV8nH247vHQEnA7cNGt3JInJwvw6KEvWi
dpJTtWQ+DunFNf2109Q08uUXGHpl4df2Puo9SYdMjs8G2jtj1febyk4QxnjhQbp5ix1kza408WPw
QN4QgczTNkL3kPaO067vsouHouMR8SbJsQ+HVp4QVtGdNvU0fnWVyWhX//CfrdclCg2GIF756O2N
s4w71+NgcfHQY3Y4K+JtbAmMRf55KjQ9Lg5EcecXQqGZ1iRgrKZ7XmAo5SbC5lHOPsuLfDR0Gel/
sENc7gX8UG3c+JSckUFStZYBpt/xS3oAntqE1z6uIOltEP/yV+n/3sbM7Wmuq5vmbYvNtccTaJAX
OMsZqu068nK6bKRFli+M+DtLAQK5Xy7wQId0qS7QlI4P6sN2orcT+RMsLMeF9cLRYATcHi+Q1LYP
7rPFxj+smjs6R8aXRTttpemK9tq6T7Y5J9qP+eE7OvHz18ymuVo3z6KRM8XzQvL3oIKvtqyJcnz9
Nk0yZ3RNQmIEgYk/5XyeERcnaGfBNk1C0ggYmHbtU0mQW/a9pjluhXpIgm0MTfUpxSKaK0RGHifM
s6CUVXkCFcz5s/M9C5YU1z7xG+rshy4j8nmTZfkTAIdRLUHtNgXCvBqXDR43dS3xkAeg7IQno6Kc
KIJeGRq+I/2YYuKiXXWrbZhCEXW9CRgP7HaRhu7eP+JHtCZansOj7CoY1Q00taV4Al8hiyDMXrnL
yJJwBi5wmot/YFpez7ODK8tLHU1MMRFLLFV/h3Q4Jiq3bXV+zGHkFp6rkV7bBzcJcOUh29pz5x0d
pdymZFSjPCjQ5G1DlgThb6ixJKbbfe4TWSYesT1zRsedoH1l/hjmRV6aXlPbhsDNXQC7h5odLWhr
e4zQKXQkIVmmXVIaol3xVcPirIXRrxov1tl7h+nIqO5z+DL4H1OkSvYMSU5scMxRu9f93QXjHRTU
si2pQfAkqFOhtQeX6WpoRfBf1/31MIbT5XQkj6bRLlyfO+DOmNxTCNW34cBbEgWT7JT6D/sInsvX
pmK6nguCieiW2BUqI/gBZ7/0gyKz26goysHT2rLZZRdqrPkOb0+MSpOHGPOJ6OsUQDi4YgTggC5W
z1I2A7zGo/hzbvKzjSQBWVik/UpWC4fLLlQKbrRU1harYflsSMNfQppIMXHp678NwlLVd49uPl9p
JBcOvrqIKbX/gj1tc+zJB7S/jWiMCg/UQfU+mqn5AJ2i3mYlOGbuvIvPM9NcbqlGJ78/uGa1hXEU
qVvbb4wMGPr7R17buFR37D27yXnHk+SpQqL9IW5aOKys1mXvKKe+zGBFggPJn5GpRh1fUUHTz0+K
7wZmTcOjp3iBwkbpnw+XTzPvGakGzI0asoVi5N5j/2mTJoPyvUXhIskVxlz00qADe8Qt1APB4+Yv
BSCrojBZjNcZmIc0ebmRGTAuYqTBklbmaEQA46EA3kzZKFySViQ8ctKf86srgB+9sqTaPZkzwbG6
NMAvM9zDOJv+7lGra2wCbw5pfvN/DOVOoClyZQn6z93F45/K3ZP5OBB/Rk7H0LUxH4UvBWXRUiME
0KXwC3LUZQOJc7m1nfHS/9wXTbO97m8czp2jNqCecAwVf6KzPMq63TM5hrRAO8Zi6SkBMtbcSK4N
NOZkQ4hAoSgqr/y3E77cNIoAS1xex+s6DVfnkzDr1YL/esd69ubMK3hHZj/YCgYe8UDqzeLF1Q2K
qcr3KNnd8gbW2qLsLCVbH6iyfitBEmc+UBATfEIO145LIfYG9XX0t6QO4nHitOKZVz4IwIaa9WNS
NeO5mHiVf7wqgEl7kYVeGFjGfXHB/OAagp3mWLr7XVa0LbMdez0XBzjhFpk6bO8QNeDdmXLYXhQj
cpnupCFITTi1ZeK9dp0UXTIa3KKuOt+WxP8bNU6i5BG/27h5z0Ip+Y43gduo5r6iNr5SrEY3RfB3
8TXpwUzM9iP2MoJrqN1mVWgPLRadpBwmdySdVXG9D6Kbr+29FrWWqi/Ec7JL4BRGaHRvYVEP7SvQ
vwAs23XBpNcvSxnFX52+X9+aE5yGYfhGKrkerzcJsvRXsVDXQTMDrOm0F1VckjFQbVaRODVJLUdA
dJUdn9k6QGjBqYZK/WR/gPBlHfq3dDjNUKBqRRZZvaLCWdlCn/l5kCayiIEENh4RayQ87caXIrlp
uYHcxz8Ky38IqVdpfmLOMJqyPMxDFjc/5IW9FRIqGXuN3x4l2b7mU+udfyAAGOcj+WkWF/aXiZhD
VqXQz/uNa3FuVnmVyrEaYhcTU16Bw8TJtcrrvEqGeW0h5khSe1nvKB5f2AEe8oNRW+2QByN2CHU1
daac885E7wQG4r3sm13wgpJzZJwdXvFWvpwy6TSFrPtwoKWenLVb7k5O9KI30hy/q6f9RzvE3gbz
rqlS3yWrtKLs8RLY4IQvTdgAB8bQLjlRm3dtLy5ElQC564opvRoSSbjLqoPcLw3arxsU7hOw5BKz
ECiE2KMxwL7y4tGa5Mkodd+7S1hDSVJI9SUif4BZfhwJ5ds1mWsGdF10fH279p/HdQR/TsHGbaRt
672ruQ2qaCOAcpft4E7L27o+UMnOg0MDXNHQno46Byp8LcNwLAM0llp4Ci8u3mnxc5NLaOV3PuMN
654ZabOF1fxNpcizVY9Kac05hjeTuIPOjh/UDA8hV+Eh9XFyTe+fMdgTrjQCYo54PDC8qocmIxxw
ArHf3C9WioMgd4BV7UBTPClGwIpf2yCnaREdELQ5NeIG8TQGCVqYH+tnWcjBitkSOuQ/lo5eYzGe
dkhf9Yd44mtruEhev6J/USGgbMMNmcK3qYC28GoBtrk6SPGrjun6vgPKbUU9mKsHSfKYEZQJZW7B
vuQZuB7IBwfRyDWDkv4Q6Y8BgIVKi9mHj2FAxnRthk8eLCRJhmxoJgGmAK8geGzZp1VK7a5tVyJr
phkvTc8K+SAxIYT34MdmKVSq056VTpIifZ5eAZcqrSn59vMXcWJdG8p7BNLyDpP61SxOYl0m/A33
jrqT98dge95HUcO4sx6PZO5s86/2e9EsYPJ97r1hirxlzmbKsvVIlsRft6A2j7WTyI9QX3QLmd+j
zTnvxuI4su50JKCowuJuy+Qpaq4FIM2AhkihpRSe1fc58SCD12mQvHqMrQQoN8CL3V922R6FNEPZ
nD7okXgw5ug3YgZ953wezWSZUHBJcCR2DGgEPfQ1YxOn1O5dZepVYH9SrflEeQhl9OS/eqqsvg8j
X/9SVDp6O6SvRtyGHDXOVA8vwa7vlq/5DbisZX78YLrUm3W3frdcGQlnhBwdtUDNr/z7lA1PfCbn
ISAON+6okjQJhCtz827I9+sbWye1Gf4Mu00qJl5Bq9+U8G9Kpv01jbB9kq9AhIHXUaBGzIhhUthL
UJab778e/KZteNktXAVe1UbEgASkaRtw4uVGAaB1HCnEll1rCSeG/PAj1MCkrLkwNf0+SVvTeaey
RHThnTfuTnJ3BJKFkrnAKGwRgQvtTJPMZdH99RFsVpMHiREr/7W1gN5Jd5dAixBUs21ER9gJpAiS
iugqZeHvPDv+rNyWtmsT5K0lwK2yw1GGPO6Cz4Js+Sf0VF79nGi5Kh6XfKC7z7FZ7vMhv2m4CQZL
5Sl4mSdt/qIG5nj9tvyRK4yj5Wfs/NnsI9yGa/sdT8sE1OcYjzUTmunW/nx2Bmf2S4URcsmlwznu
vNM4L2eu9HuV6Rx+5i1nQVtYB0cakLz70dXSeTbbWTwDCOirEsqM57Qiyj/WQmXMh6RMXcS+dZKB
dX/Lq1/MB38foH6ww9qYYjuF4uvsRrnbYp/waab++JCU2n/Ge4DwREHYhJe+gdqd+T8sP2Lx+Fdl
+pBoKSXr7+IbEZ+IdkLarqX7XKK3ZFAj8nNsXI7npsypAtDSq1JWoEqzFVfGs2iE9G/pjL4fgFiU
08xjEAjuFKFlv8TfYS79Mltkl39Ipblj2GSN/c/+5Cp6JS8j0xRtxJGOqL+In767MvJiIGpaVPR8
nAnBzoRJjPSKL15EJo3c13iS3g0rHlv9LRmRzelThGPt091Kz5bHCSUHjRSqfPvCh4mjEzzTYKAk
P4MjucXmZqiORTZtqXghaQPBMPBZbMTvCU4FdGIZ0LekAwJvxIMQKzEkKp9Jf+DYDrVbEITNjEfE
khV0rouxtxoSphqSlLCQob3QqEJkt6mxXJPTT+eNDep5Fy2aMHwF2HL7YjlCKTIj9gpGQd0fNhrZ
RQY5I+RlU21/HZs/seI4xmNgNpPOMqT2xKhYdb/E0+pB9YAeR9HyZbcu45akbYqKtpXDtx3l65Cs
Y5owfjK0gomLXhwAaXyLy2psfhGbtLl1P1Bf+R41YD8qJny/Lt7CgXm2Bd5HP7p1+4KdlqeYnEL0
OHO5TAVMz5St5tdpi7CCIpRRlQqJlJalK0dDoSgWK62algb0iCude+c0FAeJOdG2k9lzn2d013V0
UB0YnNH/eGxdT3Ftcp70/rqjliEivTFXwc6qYHpk2LtwIeZozgodqAFpr0++oYnjlqKsodDgtOcm
hndFfIjYFbDKjjZaJAwRIdWjieG173xpvu/T9EME/XdMTrELeMV15oXWX+WgZA9KmeP47syhXbfL
FbvnQBRw7xYJtwAmJnGKxmNMbLlUZZQ+Ms7h6kMybhl8uZM46h4SEBdPLCyyrUMGG+lENuATnNDm
wQeQ1Ps47EPN9EPas0u026dWqthtKXvwsAwaxz0xbM0psVf9Fzq6SpP+M7QqEW4oJV70neSnTG8P
zn3NvKAIEgG+ghtwpgk8IPBuQKEVsHH70K3NS9YIgNzjKOuDYQK5mEe/qT4Yd/fZ2nykHnNvd0Bj
GGwswq+ZuTUwGXLs+VYYWC7UG/mBritgPFK73XnJrMFiUYae1cxt39q56+Tgp2RUF/5DM+EhIOzz
XGiH+gGdGL8aCeKSEXXcPYAtiOfhwBZpN4iVf2QOAOTdYjgowcdQnU/SDRYpE5jUixi4zdMNZTl6
rVImWATwbzZIdwnmQRuThRWbn4ufC20nxOhKpC1JfibayEPqbEXKaxLMK09Vh4nwtCGJHiCLIUuE
x34103ZTTBUaNteVlVCamp68AKcrJnshYN8rgIbvWnKrBRjXCJU58D6VyQMToQsceaHZ4gEDOJ5J
RM03guuQBwHGpczObOyOCLbK3r7lU68fLkosd8r+B2zs6ingLy74mblPxJYZKGka2Z21j2XRvVDz
qlYR3kujnKoHznNO6AkRqLohCfCciSOL9czNZaE7SrfcTp2EC6LgqKJ7jJDFjgRmuJEkjzW6jMZs
V7hNAWIxbB3A5tb7Nw3KZIsp8dDJuK1lP2F1IhJnp7Uh9T1g2Ed58ed/QfhzKqOctgUUnQIu0XV5
gLbjynPOek9X7d4jma6vH9dKR+nV+N5O0962Vmi8r8IhQVQVSj4SWAr6S8Z4YVIXaukIoPGwad+8
swnQIr3vwkjuj0lWfYIdpMsbE9XxVrlegwQ24PD8NZ5x1IHS3TdUmFP0QtBxNc1TlczlpFt2APrJ
2208h2nYqtK/FT6M9TkFxNgejQgSghVBgUX5xMHTd20rVEsx2aiMqHvWoGINBWG74egdOxJEVXVt
KLSwUd2qY6O33E22XAdo2CWejcUBaue89DHS7AVYqapOfBScwoU6AYGYUekGiJsdIMpzQqefl8tX
68lqaO1AiJnEOvnHm1MtCls46m3wb2zNb1tgL0AGyL1TIZkYE6xbEGSH9xFQrQVs9xzq/MEo4KZm
FQSbsZB6s6ndajM99LsCXACPQoJ6quDBkiZaVr4mdPB6Yp6ZxONnf7nIWsAQ6ezuEXPcIJooDKPX
aiXrOOFU6bp0bqsoIBmPnwDK8T4qh+LdPfkojouNhFuUrtpz1h5svVeWgf/2yInau6FHM5U9taIZ
8pZPkRamC/im1v059bFLd4i3A7Km5Yt/GHDx29SjGnB2+m4DG4e+3nMcL/RH8xg+F/LWH40nlMCL
9a+TJXtbVhs1Hb/SqZtqBIPXOH/6Fr3k4bxExU1uHXgp9EmimrZxBEEMWFN8gMCl8/IfMQzx1Axr
ySnqu8YxPhXJzqDHB5nNbXIs82SUu2LcRd0W2LlRXDQppM+PmlBS8M4TjV7bB4epq0tG2PNz0MgY
zyQuTw1UCY5pcWGnpSUuxGdbWSLkjhRDtNTqHYNFZvBdvOVtsP0aR4Sv3DxBibY2IG8l+18yl2Jc
fLUSmlNjhuh9uHR+n1hko82mWk6AYp+be9n08eTdJA5pAvvgoel/rMPmPsEW3v52qVuzuDCLv1ej
wfG5TPDQMA1i79hj29ZYl8cXp/EFQ6clakzBFTR2M4OT/2T2AjFFJnL2+J1+hp+y5y6G0i4E1Q2e
kJ8aER6OIJWLLJPTbgPhGC4WcOPfQ7IC1VOJ95uMUyxjCSVMbPEr967l3jd8OUcb+w7fOesWjKWr
U2hKbJ0uQ4OdxmwGJ2+ORDweZsYaP38gNtevYfegeipPZFZO/oHVuh2G+SB1BQLfdimfVqWoFeGM
4ja2mOMc7uTTezR96TqBMJWnulXg0toacESzv3uC42CQhw4uD3yR/bkPz+zqbAsF/HtRtlK8Z2Hz
wqzxec6/HwldalK/bTdMAd2z2nOD47sls7rq3KLGBJ5+ko9PSkunnukNGd2L5FpJPKzH5jeQgkib
jqyCO5DgN7u6qjZizglGl2p0oC4zeLDXgd5S1xWTtWVW6x1l8i9SaCNa9jgt0dVuXW5BQXdhd0UV
XizFQ42Mvh39Arba+rRLKVriLs1Th9ye5e8gcCSQ50dzc9ILwZkNlDPbPhl+HVModebSZpGuJLAt
ru0lPZXqSKeWZRx0YqbCdKovoTe3wzywI85mynT+Bg+71MxhNckavNhWGUTugZD6cfX4XwIRC73e
Sp3li7OWI/hDlxExMF/JVSFYCZ8Q7YkZBlgSGjb9jntkUNoOxmQKtS2abZnqxadby0ieedEg6uSK
RDOc8Hs8ofwTnAbS3oyC/Ku/bl6Xxc4OFah3nE3b9HCgSE97xzfK1ZIhrZ87QJgP8vNLo3hDhV9s
ApUZ5lv/WO9X0Qbt3uDDAZ3yXNjwALwqCQI4K3KCEgx9QMaES5xXx2gOhKfTTp9Wq8CGoBMndBis
FPmqqb0hVQuS+4pyzABxc+Q5QZyZH14G4pN2ERjJBSJtPojyRzJwCVeOeqCTq1iY9ZZJEnMp5NAK
xiNjYHi+Cry6oNWcwubMLumT2LwBsde5FfB/4kAN46VcBnrLH4Q7zBQyRQ9l0Pz8CrI3Heikg1xA
h6K3pWVdntJHVB+Ij15XlvJA5QxMYxrugnt//dLmDj0PbwSD4tyYNU067IFz7JougaT9zjxpWDZc
SY1t3ejIi1mGYn2dohtrkiE7eMShqM5X48FKxBLBg+OH4Wq8x6bifwzPIUKrs/07rqCtQL/NdXxW
gjJ2BWPDqp8lUEECTew9ywB8aVzVgE1/5d01VcFBmlua5HSvfSOhmI11uIDY1AHNnWtsnmfZMtL3
hlPiolIredllSp+w2V20JEOJDZFvIUgjMdjlYvClerWrqnQbQIYoNl8PU0BPmRgQx8PFIj1hthIf
25MBv8BKWGPS1oiSNt1wM7zsI2rqdnra0shOo14XhdTT1iWWSyvjfktoWq/DM9svweM8PdiPSBWj
7Eeze9/xObFoJsX8G60zKV3BEoKCBh6hsrmwaslleJUTaCczXtNANvTyRGTf+mk9FOw/3g8iknzb
U0ZBNtFnzZQd3wNqImo47bBQz7AcFjqRKKp0iqZQHXug4+EOlVz7J/Qt3XhDOv3JLoAekokDrGoS
LcePbpOP0/jdDKtq6HhnALX7BzEhXu7mO2oKnt2o6IeGMc6dzBwwTTXtqJyHjyrUL7CEStHVS2d4
zvkSMMFaO5NBMowogL9kl/r/3Ka9nwaFy9Z6yUfn5uo7ilBryZ4bTJgKcrOzF6AdjBmehN6qjkPh
sKSwGl3F08YhSMiMdiqRbP45oujusW5tBUk7PwhNJ0dbKTnvJ2EbPSbiYNM4dKHXRAFDlOyrnAR5
wqpuvkyfOr01Rz8dxs/ZdrG/9Z4m0id+Tnmyw+Ly0lt34rgWSG/YOWQLBJmbr7liy2kwmFvUVvbR
OabJ3wqDl/osQ7W/Cr0tv3sUdUeY64knzhsTSni44t0s0IGk+i+s6XaCoNqoj4K6Q/JRKY3Xa5BC
F3ljln3O8UXX5QxNs0Fh788gknSNWmw760CI5roqWg5/Wd3OD3U+okeWgnuP/77Uu5fBwYST59ov
7z/BD/oBTgh88p6Fp5hb1z1vesKMm7zwv2sEwZnVa08qC1KxQsKsDH/DgbVM30q5vzP+zHNtcMAA
PiU4102l2aF2NOT8wW3peJTu4yT1kC6qT87/N+rIsRVny5F7xT66OZ8J9ta6jWV1S6+nGDliYek/
PU51VL4V/p557AQXTZONJ3trqP6YJ5hPGpBj18f1WM1TXpOQ0tZso35A+KuniGQ5OHVpNslzIrrH
ebc7l6xYBHb8LY93GWl69qdXiuq3dncC2kBMJTr52BRVtBdDsRamGfJnBOMmO4DXKz4r897JFfsR
k6EuSzwVR7ebl8RF+ioWqM5suA6i9bsfxV8HEn84BujmM7nd3M4aPakBbnS4aWDBqFcs7YcHcRCe
6CkNdfDLlckFB1VBKmQLzZt2uEYrJQ0zgC/j8gpfsB8IZ4uQdxB7AaHZgACnjuTykygdr/4MXPh4
HEpIKuveR1yXrjOTL6RUHIvv3Zbtv2197kYXDQV1pCh+uKoschto+H23XnCAaYpNSNaQJu0QI4ZD
tlvd5Jxs2GoijMgJU3L46I6BSxqWAOOen3Ged5Uw+hEBY3YYbgx3saPgs1vopynVSfxEjsdeW22H
KPmXe0mQ/U46sM4YG1nfmwrCrw6JMPPcTQ3g7zerkd3Uaxyj92oxntRKAbmtVkCa3XlwILYXDiR1
1gs+rFunukdVXVDKs6pfGjHocMzSbr9TmneH2EhS+RJVRBXpXLiNQfNlzjq2iRxv6DzIW3oEL/TT
O3LsthTF255nPQmowJJ810bmOfMiF8uFoOP9uaPH3N7iRRwtefGX+FKHH75NClPk5KIZXwz3WUwT
7P25z76KMCJ5l9gSBAzgMm4kM9vGkaSjsh8bam6qRksxtnQYr3hnELTs9oEKFVqSUdV7ze5Z5uBP
TsRDjVxhyZQxIFz56VKbVIKGNYrj+rtowIKOLxloX7K0jyu3R35i2kbACkJXEU7bxPb9Z6ArWRnj
srGK95TVXef9XbOuQz/q8SR0CUTroA0ITDR9Tx4WG06XF7Dq0TfsmrJioYYZSPyyfLRM/YKeZU7d
/QhCwOOLx7XK6AivfPZL9lZZti7k32C91QyAX5kEaWS4M+pQP1qyOZjcSpx6ShuWSgcycvd1ZxlR
OoKOFm9GZ9YeObzvsCLnC4IQ0QAhuyFJmMziJ4SOLPrt89Z4VXyYxq0CLYLTH4u30AKAUmw+AWep
nSEbToJdOvt01qdSnpF0QMS2l/7gGMgeqQFO1nJIJDVXGVrgejUL2Fm/S8w0kl4rTrAw6T9bI+O3
WS8H0A5e/RPg4dlKTtNjsPFaI6gIjY+PbYs5GOW/ZhAhUgkmlWKkOj0/OuOdbMLdeqJt9c1PaXcM
1QfqVvW0Kz6ItLgcorTD9jb+xY9E2YMc2eL1gKytNp7EjKOn5Miaq6QtxEqleuyhrjAesN8rP88+
P/HaIoHcouV4gJDVJkJVu68IRuhFMMGgv/rE8p3Gyo3flcSTG3J+NH1LqCeFoC9g4PSD6W1ZaqGx
xT9TvHNBrXD132faV9LnOSM23awib8jljpIMNEQKmtrzYY/EuCVOD+Wf2GoGAysmgZFforIuOLeO
dEOarCd1P9OyVBrLSx/b2/OVxRCB+r0S/J9B8OMjOMMfBgVMFUsqHTutsVgiYhImrsuBHIdqUXdp
3VBUZbMRTnEoPtfN7khm+xxwtWkDpLVl36CsSQmZcET/mxojx3R7Sc+nCjVKEgzDXsaPz8oTsdQ3
tFV+U5JTqCO/zKg4oFTXfQhJjABZxwjUxyfFEL4V/Yml263Dc1pqPXxi736a0xN2n1y38QmVnFbd
QMG6QT3nubtcSEF6NGNGwNJhAMyLS3PMZWeO8gMZoBnAG1Uzr3ScBLixyiHA+C6gsFR1OS+GHE9r
mVS6LtPBOK/2uA+BhyRHXhPwXZZr0dD601IrX+cI2hf1W9F5QDMWQiVGv6ViL0rOwjB51dsyIHGv
b7k/8sfIZYsSLsoLYnQTVjWZC75VYj7oFYn97AKpDdiqGGppOlrtaIul8djOIWSV/BGa8gINyo0W
pkKNhDBMjlv8EPsboGvqfK+/v+Q1+grTy9SFmRpMSRnIAUEXZD1Wa7tWdArL3VgRI+2Mh/Q5M4qT
CTG/0FmMrg1jI+WNNzUrQq7WPtASzPdYpAc211THf0YkbErxsmJ+8WajpM3WFDgzWBZab8RUZrS+
rvmTY/4lJhDBUWqT9MvWUVeSIbhLPZvmlvyAGxVgbxatZaixwJxxOP0dWVLDLqoAU3jtn8lssxNA
OuDpFeo9sftYuIzJKf/8SLmgk3zwSQA0+mzPEIHxa+hUP5Dl03Hjad4M0TsZ0Vzy7i2lDSgD4nlK
4eInlU6Dg1l15PfaOpS/pX84HFF8MiPprfmix9GU8B+IMRhSpEUFJmmn/Rf05Ob4NC9rUp0x343W
1V8J0RtWlpAA8/msWhzSFTIXYc2NKZf/T69Oep8bCCHSYYYsxKB29v5CaMHG7Agz0PJxBoIl0nB/
UtX3CpnrJKFacYYx7XVxPv0Y7P1VNxNr8vajqrmTsd6NXJHLayRXTba8/u0ihuXVEFVzqB0GrIJG
wgx+Osss3Z0SQecyw/Xp5/Bq8jgCung6s8E+Yp+vveEcnafC7wkxoVhEshdpU5Si+GDENPp3k5zy
DyjT5QwKfi2MwBuAPbSueKFVt1obRYmbFLVg0yvZ0uq/HsrPeq8OlZI8IKxXCYtJgspuakYaTXMQ
a1U1kmxwIyHlIzd8DP7RG+he0DxogxZrwti8EVzmUDuz/k52Wsjk7B6SdddVAY8gIyFcp2iYcSXb
OG+Jgkv0uGtJXCEMPKl4nO7lQd5IvOCGh+7orENUZwhIx1y1SKnUnFJp0TekZknqK4GFAv20kwBw
/LpcgYcvE0KJTl4xnRYI3ietIIvK+VZVPgg2TBh+iuAnUMG4JouL7YK3RyU9SM0VYQnUy55TLQ+h
CkSABk3GAvW9PFMneu+Ic2uk9VdOky1v+Frs5PQkH7yO2Ckt2vp3ARlw8qncyHTDwmDj+gKRcU1s
Vtvam1K9MaOwILv+V2Zoyz/RhsXsxzulsTAAjb4UCFRWIusmVd/o+JwfsP9UndAL7UL/k2p8T2+i
9LeEO9Nx+P8unfehMLvfIa/7W2bbmvkpGYA1RStFvAw05wYN28qIoVCl/NFgiO2RsuAFGS624t2M
EaN8oSkNqo3WqgHATkLJrf5w7bqt0d1CzWnkUW088tv9y/zV2G+gsKpUBzkMBv9liq1l56Rs/6gE
7OYPx7pdLjkPxBbyPWxprk95azqRZ6dpwcvLyUYMmVfAL+hg1GIftCr5WQXYHNkQaCm/MZsrIHUq
ntl4VPAt9V8sC5sMebb6gkXMNbUkvBmItO28fxzv1Fasf3m/cfSaeMHV5uBoy4d+G84gyyUVEIWv
PA4X9YHTtD61jRuWZeKfJMvA0ZBIGoSDwCAd0PR7HTmz3RcvK/FbPd21B9D5TOf6E6TvQlZxssdL
uq4K/e2/KcDh8YNF3eS032prb5bYlaa/rXCVv345nbKJm7kXGJNxFmn6FWWoV31O538ubuGoK3Q5
vRZWseb/MLZFq/U/5PZ60ulGMRgNS46HdIkuzPksAsMCeWK6iL9qFDEhuFlcpDgwN8Gp/dU3cvo9
9cWfXRgQIUZ5B2jTOgrc8AdW7kgeFHOUt45ismXtOOLy/Fw13L98LsGZmJY8gq5O9ufS3QGm2h6r
a8bPnBonMuqahUB2gBTMZId9TJJ3MN9jL68/ov5ky2tgzHMz60PdS232DMRhbF2FufrKmlaRXN5G
8imzVEYcaerFbMT5HazQxijpKIyNZKAuEC/6g+htn2APU710UmWGE5feP7i73afUJsjEcFpoH1Dw
hko5BdtK/a5dq1HAACgovY1s8BNtewGRKMWNPvpscyod01z0uU2Obectuxq9lYNM01jjRBMogKV3
o0Nf5HGE88EGc0xZqo9Dt8Nv1rB+BmhGK+oZGHY4DQ5EpIhg8S5mxnxnq/EoULy+30UtHjkeHYOw
EuCLPttuLT+39+Yp3x860nyMBPtdZmsgxGfe3Uru3FF6kcfKEvZnP+BfkvqPwRHQqRdg70CoxRdS
Ulec94BpyqIHfQKkqhQ6zz6Ni2PZfOdgVVGucNaunVh766APmmIUbnYmUQbw0IOutfiv7MvgVQAw
g5VWcuP6ZOJZ0oPpXEdcPvoY85vgQ98LY8O9Jx2/2OWKNyvh6ms81h93+c0w/MwJGsgxghTSUe2A
OIGhsmwq2pQP7f6n7EmS6D5HeNsEwTdvQ9BuIB2TVd0Hz61sLox1fvwxYLQ8qBk+yo+VcM/jjCGV
KhfkT6NZ4lrYmg1+zzNj5al0ZEHkIcysv+kh6GqMAjyHBo5cFyDgI1erwv0DBSwYBqIRwYGW4uC/
jwKsyjwk/1Z8Q9K0ApyLSelsc6qfItAo+8A35ZCtV8LEozqBsoZSNPA70QEmUGzVNIV+7jfaVdem
O/c+3Kw+F8HLM1jkOf44/pgHEyxLi01zAWPcAjvcDqAWnIeAolaik2RIfVo7BY4rzpR9FX2ZPPHq
j3vhKdfPHI5UnRd9o5Ti/uSFvds8BOkZTzif4Q4u+1i5DKS5e36dLsRItNVrt462TrxKaJo56S1z
zXXuNaBIlCfJL500RWa3b96QJ1LFfZq0yhc4gqB3mR4iJwulis0bObAn/oAf0RalsCX+AkjM4l0u
YNYLvEpJM4DUpXWIx5wOtRwXuRvfaq70oY8l9wVZoHj424dkhRLt1ySqR8o8LFCHNsVzzPUAhskh
o3f40LC2EWpliqUukiLCb7/kpwFTQeb0q3i3GRscD4CQsij9MIEIgmn5XmzNOThXKoxGZmKnGj6W
FaRSkopTQfeXZIm2rFZ2lYiIUNAmmS2fJKUBvQHKpDRvStvNlsb9AqE1t27894BjRGmZogHWFP6J
wViuoacco8BHbEeF1RBsCwS66uVilCHxQqApMsHhb5XEV43WCAeLFfETYYECNoxe/9S8xFbjJki/
tHGMC1Q5F239o6qUJf5iBLIkTcHcHmcISTe350IWrpAVPCTAY5gBPDFtOil8tL7NC4eb59E+KB6o
fBh76/aYFM5v2ocDwsp3in+OFFWnNHguFfPY74xu34Gmz1vH8kzOZyva8cbJsA+I+MQgbzdqCgR6
C62heqmNtJLGVGEUKH50/xiSLBRCZcz6xi0WLxa2GNKr6q87tjskzo9zS9Xyf3OQC995EBckkHZN
seK8KxJgG1r073HvWpEVqKWZUobVgLY9UBOmWJhaupbZApXnsZH9WRaSXxt46emqfPN+30eqCzk1
zX7PAvbWepJfMMY3Z9/nZ9FjBOdDybYYRTKVmYdwQ2I9X5ZNRfEKlhWDrxfO1lJzjCbuvWveehXD
LjCIkaI/J6/IQcS3vo2X9YbjSWBCga7ROhIGx8OHIwMhzx/gsACBQ/OQog9WOKST0UpYACBtiaC3
3JRhHCbhzMvqbSRyFFzuuJRNYkRrTjh3eLaPpuKUHyZPWFUQ8QZgeg02DDG6CsjIDZQ3SJyCrdzb
2JNRCYiD9AWWowoNLQAU4wCLPzoA3hyJwmlna9RjKZXMrxcKxQx8rWS4pTBW28AeiXWcVpQoJ7v0
cdesGWutBBDGGCvDTpRLBqhAT1Z37VMI1N0VYksCSIpS3bDfzR2kklCy3dijf5jaPz7SRJozUOrS
qeGJTYiB40z11jEquWLoQ/o3ynRXoAIcXPMBi7pkgxHvLHZtd6k95DAuK/0SqY3Gv7IbdXVyqMKI
AjDY83QXQd4iRQe5eLNWcdr3RKR5uowUYBOYKAVzP7Cda+zch+LPiEDyXUUr3XvV0sOAq2KIEpH7
xpK5KW6NF1lXFn08mC26W5iVbl/8+5BiGwkUsfQ4IpNC+jnOP60tGlo6y7N5+uhReqht3h6ddSrW
q/A15Ow8pRSC2HByKdpvuXjv5zoV6Tyrg+TZmwIMwgI99FZQi2ZEZ9zfUUIdDantb8p/+GfKSjhX
8jJTAiTta4eoei7HO4G1t6Qk/qGo1CyqAqDu9qtv7CRi4sex92pNpZUCPIzCEQ3GiBF57bF+9NpX
BJ9hqrmBAwHObN3+ORkOo+8AyJE6+foP899R8zPErftd49ToSR67YDyFUXkjIySMu9ZdUUfDV4K+
0NRK28wEXWTdUmjJwaLLibHrYSOP0OQCzmJLgy8vfSCowXckF769qXbiwq1QqRc4adJ46UgyuPXT
6vi3laXOWdkZIgXzIak9UVxd+XA8e1m2CYyjKwc4EL2oK7w4cL3BrfdP9YiWd1kACeiFPdktGYsK
SzgC5Desil85i1M5rWSRvKgIhIg8GB6lUtphR3UnWw6BdwZY3+hWTEqljHYsdvjHYrmGbGSfxZxs
Md4tS0b+bzk6LW4SsGINJCTqTXfj4Zetu8US09cQMSFlGLABnoCb114Ox1RelIS9RmZb1wkTjYeo
XhjdmSjCRXhre02HVnwtwlTqapjJYmn8YE4iwPE4AcAH3g5X6KVUCedaFtctGAzuidfoYAJ05Dv5
EPwtmrYCUAkHNJNJvj+GjGsXwHTctAHt3EuJpoB7RfRsX8Be3FAXeGaTr6jv+GEUu4d71sL/l93R
08Y88PwzjmFCNuFV1a6JsDn3mSEWlmrdV2uBIlrB8dlqM1HpYAUzlp0iSWGbsjMyBgMy6ZETCAFw
ha7+JwOzHrOPxi+s9aGNchTyHBXPM7YAONpC1yKz8J5g7VhoHzXK4A2chkE7u8WDCf7S/PtJxCW9
RDQTLVp7I/Qf0CpitHYCwKj2hNop9UCxLjtVsrwYdQOKJziYT740LBYODVk4SaPa89B9f1qzrzef
CL9fwuyk5g4oMUwknpsBHP9ZzT1kvwAs6eUnZ3wyTyZAfIO8nzl8AXFgfF7qMNVnagfp8oUxDwTz
/eYQyaOGlBTjxJfW/lkrnwMueB2AGiWeQZiRoKzobzOc1b/lXHy7ggOfqQUeC2mzZV7juQcHIeXq
JsTUOC3XMUY2YBkdrHW88dT09rtiJNmO5Pz6/zjxQHPnzkcZpi+iqHejcaHY0LWkoHyiisWzFXGA
HV7mSiGYh4XgM9RJ5XgiooPh+jQnRBRw4W5XwowhIkGHsSj8n8x3T+qv4MvXwW5yarYI1Rr9csaj
bxLlMRXSHsYY9pOkM1ThDveyxT4msf1YSeXd9zFfPrwPkSy30I/b+OX1NumfFwBis+ZlKirHj3J9
XBLeHrpe2A6lvcuF+U3bLH15tTxvFMO2eEZMV8tQPQmF4UPFJ5aahoRUXpgyd5dtDbXqezhw+xuY
xP3w2Ar/kYk2werDRuMK8kYxRl7fcPxZsf/oiwdWsmCTOhMpjdhlhdccML1I6xhlEcbVypTilHfb
JsMBOzApg3CLQ4pTp1+LBOZFI7+UOy0RpE1UDHXhDycKOstDHkPRkU3k3ZUNtzut/P66xN94TUuV
+BgEl4tGa3cRs9bZGhDOg3vleTYy2r+L9BOIamw9NiTDT5f8nKerfkiD1o9ZQoq4w0HA6JVZAksd
fF2PY4cUCL4MYeMMqB4Q5ZUaiZ59Py4UrKjwAvynD7S4SdZ0XTYbf0O9y2X7q7Yu05ERL+yVIwuw
+3p1mDDCBT97u+rTlHfGpK5KpIBXe2x5OClYiUGlv22iN/zxk/N4CbkLhTktgDf6CHmgKWNps4c4
FKEFCnEYxOM1YDsj1IIEiTpdUvzbT9T9UqVcePfBsZc4xoqvECC7E/u9P3EBFd9OvvsDEhuuUbAh
bdUxZ2FmB7amu9gBQV8rrBdhs1FyHLvtA+ohWFJTqTEHMm36Op72OZ5j3CfnU5J5qrZiSQZsk8ho
si1zdHMT/YeUazDc17Q84nLo5HwuWZQalCCHCDonIf+NDdzPkPnuCtZsvO8fzmULaqNnCwBaLmix
rCfHuFcCtMpxyJZ+IwVtKu0Sf28f4++Pyy41tQiuNhcWdhycqWnVgXlw15Kxd7/nFtMSW0r7Nnny
RVeTK1fSJcY4g5jfD0X3s9GandqWW+gOI0w39r+S7AS0Xpi13TcVNOmFhP3Cqq0IKtwy22hJDfnS
935Q2pzzDkRZ+0seTcneV/Oddq0OzvF2w3ZMrn8/8rlr7zzdEVinvSk0q7Hoh7BH7mZantz/Cnjm
bVVQibI7c9oALmwEnyF3MmTKS0e1h1oHh9KeOYIWWZ9gXdhwwLwOJtjPhHwhnXkOOl4srNpkZJqq
2t3tkpeaVJG7l/Ov+z4JLYpFLD4jh+8OdWT1LcAF7ZRwZIjTI2jhmRtX8hVmgv1RUhuHQERjlORK
7EAfrkhpulfFk6THeQwcOendAoIWxMzawFe9Mek3CNYBAo3UUvM1D4PhBTvBwixcGA6wJKIGeZ8k
qQGHYHANxImUIjRVlyqYf0B84F8BnWUdN1euSxaH2gPOpYGt/8haafUPnFhTdnsmfkZuYbyTKTrv
GG0es+pay0zAuI6T6HZgiUe3k6mlwCgxO2fmaNIT1JNw7mD4XvsKOI6vVW/CHdr6B11qcnUpWAA/
CZcsYM6LxU6IJS/FZG73LYmInVY4DnW7krIzKCvXqY6etvg1qmhMSD4iS3MbA9D+w1Fg3cGZjCh4
zz92hWDRKuV2flRKG/Biin/4Ka+g4WUzbY+rK4tWE/xMuYElfi8+jR9TpFCz5o2N8L+75vdasuJB
5x00HFuKPx8h+Vml4mJToKeo82zOTtNHRQyCTRjLkR0IT8r8cDIvdAIcGV2itWBOZh8aI5uLjqsX
XXFoju1zfQq2bxQe/k8vpK5eyes1igf9eRbParKqh/sgxp5JeO7Jetp53fUI6OL45KMqe5JyJe44
IUsiG4ov876hvkAsFo9+uImosBH8k6hpqiEfp3mr5VYkDXA6u4XmAlrbWx+U8xOCRybXIjtkZIpG
cEFIM+xVvRE5jwZfsCw3HDNWs2tK6carEj09m7cRzMVwCTwIKWGnAlZCI2IDu67cw3IFo/a3b/UK
iBSRzXb6cyidnJaPGjnPb4Mn6ARZqlcPSb1SuhtWsAwYgjGsJXROx1v/o1WvDLmBp/um7EJNutWY
pA64plzhNRzLoL9gb8CMlWyQpLjlYk4pjG3rQcK3Vwwks4rW0CF5w10G5xY5N+mVtntyYW0oOFzj
ou0ECbRrvskTVj/CNwroMWAzA6AWe8YoLCmFqjmRko1IEzZrm93lSmYmGAEaHrzA431Wb6pSeB0Q
/ZESZNlSDzBh+MJwjwRq1Q7B110eIodzFA6Q0RAhlBOw4XSratquF0L/YwCsmaUQjCI9auoa0/VF
p2tvUI/9pU7XErt/PFlpR11xoy1occn6JvEJZ/83um8rNzK492dTFf88kzieDsyrsURKwqzy7jgh
hfPLvZg5KORKbyl6jzojGuptTg6tFsoXltihJeLUy4qx+SJeJAOq4rXnciMfFNGJqQWeLX5tWrht
R5g8olQybjsus5dGdLD8QOA5urXYfX1MsaE33jL+7gOAypPPZHXOTPg5pPgoohKkyBQKtXaescmm
+iuEnpq3TB4DHTe2n9Up9E35tkWR/Bo/6fEFEdclb/kewlVPhIiI7oD0mPcaZdffBdtxAbNt+mQG
a7CVdGxIz6cI/NO0utCIRI8nqBRF97j1XoD4AHIHSBM60dp+eZ9aGbrVI8Awt2bOypPGOJSp9jQ1
5bgDuuaRHivPnQjvvsp91w9v+gkpK2EQwPqoMnXburOtc6gBL/ymwq8RlnrAZ678MtcMzq9KzJcz
hslQ6vrzQaqu8yCxxCtEGgt02NmbR/XagPDxtsQrURAPwsWzxtI3AmcuKFOMjqb1hS/QJx8cs8bj
+FwKGqzFIQtPuA8C2+PJD7bz4L977wxQ4xfK3d6jQZHoA9OGX4YEUmLCUAWFd/0HK4rtwMkKI09t
ZiSAqJcDzWhYYDAnJwOFRbfPsWjito8Xdz0mGS4C/fSI/CoRBNz/ToDWzsxRuwLHp9rm6onKfU6L
3IV+PfFLAkS4CYigPJlf+57c7y5c0IMVlqUyuk2GFWVbQRvS/OX1Sk55vVlGfUKGuzibWlAU20lA
IwnGrk3H+4V9W4nujLMmchjjtc3wYeJYlrLESu1Ybzf2UNEFUamskEA7mWE7MsB0+bPAXPHr5ZMf
MFL6zoNXM4ua160yDUY3WpCiHalbiI+rfk2n6FfgigKBjav67N711yqX3dBwiUi1MKS1xQTZ32h9
tJNS5cZLvlJKlGTSL18t2CRxAiwyt4aBZeuMxqJ4sHN8P84HrhYmNURnHWzqhMuR5B21kJltE8/C
cr0MY91T4DiaQAERJAmsfn8SrBtCtzWlHsHJeYeziNgNLl585doLkTVAMZOSINaF5AU0MbLQqlEu
xSB3AAbLDE7JWojWpapJf61fBSXwsQHPYGa3UzbPmSxzjD+D0Huc8hndR2sLaz+5iSlIk05rfLZk
E8aERsybpBlWdCtDZ9VWx0JELUkpDQSI7luHmiZIelLNDEv2Fx2GKYZ4PE6itClM5g3sb3Fu11SF
ZqZB5UTlFH3JTy//15/RnkloF9Dc5HLs4A52it9fJAVpU9rE/pCvHouGYQhcs9tJagGOt9YnleJb
wPDNQ8AfxBrk4y313zdMUq0lZDCbg9ly3vkXjWNYgfA1iQWujMDHFsXloDCfjMpCbJE6Msks9Euw
UiCMhv2PHRGdI2LKjCU3BShXO+PMlTkelk9qDQ+uMyUUnnwTKSZ9Ke57DRnT5uufQPrTGUXBB9KE
f5k90BxTDxrMhDMozG/R/BIMsYzmLbfirK6hDVcmNQ6qXMTj/RgXUVT/1hvntzB+q49Q9lxV61KU
3gKm9AhJjz/ACs0iQWqxGv77N1uBW+4YxYgy1xAFbhqELGfITPrAvbJoqHX4uACE9pqc53GNpXtw
aOiFFHiWSrfgzNsQl91/NgJT7v1iie0rW7Hm1asA+BIXF3+0fYHMLyv6vq3ee/wedvV49QeRyGI3
MfjyQBD6nrRI+kqhawK8R50SvbXj8m0tKqrdRqhXzF4bkRTMs4DoJv1w+qE1T9H5Mx1Q3m5sXw8A
TaTDmlAcW3K3fJ/gU7qd2CNsLczc34YKnN0L8uwv8ByyJi3y73ldFVfC3TAHx4KJ3cRK30NKJ6YJ
bZfBiy3jhpk4IzlNERGp+xT2azHmRC/PWJQU0xWAdavkur+AZkD9LfK1JtZ76295uJHr8VcbbqMW
3itLBoMdPOozMxhduBLohZhMh2FS6Je3jY8Yv7oXe+1UJp/kUtYTeT7zAXSerCV337hbrQluQ7iX
Ml6u/dChkQ11rmVcqABl4usCyvWWweq0vnAkh0YYp+KStspLvtMxSYkVy6CiLMwPbPOdgNacSan8
K92X7OOtatm39U1M1lIY3mm2qKjeFtYnNy7hIyqgPXCQ9e/YJirecK3RF7u47l+/W69WuUn54VYU
Da4C/k+AUU5QgRBGsqK79GdaAOshRVq+KCF8sulubR9ZINlMSnkQaIDCZPTRkZvRcRAUiIlCcclA
SZwnx5twYrc7JLbVB9x6NveJdiq6tsaKVM/DXt9usytzeA9maCLktNBi4/Ra459nbS8EEUbKlh4h
2nGEGRRbpElD5RP6jni95lL2a18zna/NWvajfDjjxbRKhuDrMDrmtaFPnJb6vGAPZhjWSUl9h44A
RIKyylEX8N9eAU6VPTojD2mh1Zsl/QTjE2RM7b8yxyKXdtA56zzsjA/QUvW9p/Svzy9a2ML4PC0K
fQtPvda1toQ4gz5FvpCJepLKIKLjney2P52m4vqZkf2whcqL+ocay8f+iZu6gQqn/qOIsXwxx+Mt
9aKEoypE6Swim0RCJWj0yFMAU1IcESHg5UwVUvVgyyu/+GtVO4zCU5Q8+81uuVP1p2Lr8r0jplLX
LXKd8WA930giIOJ9UXL8sOUaxGcg+CTEUPDGREr//gsRhuykNKPD2NapM6rLolpYpnzeMcTQWeiN
S0w8ZhiqvIwQz73dm9AkVwAIIQxVQSEqCyKST5kG7TqlIhJ/k5JTz8ibj5Lw2a9UmpCxOVXYc3Dt
O5Zm4Xev5qnhX51WTVKuRdFqfGErYrkFoIDfWKb2drS7jLutLxaEU1CMPklaRc+uIBwgT9XUgWep
wMB5yRrjiWUMNjHvQ0ZQ/e7WXa1lLO9203CV0jZp672Kjf7lzxyXHS9t1EpHtIVn0YOsjfJjicBd
Vb8yIrPmL5pyHthn3HVJDu3zvQew8ShKZoPuMLJvtVeihG7YAMLESvmGbcb06psSJ9hl4lig/f6q
14/DwvRnGKZ9cGc6dBCTtaWasROF69tfkIVYCvRDqrh2m02WrPwkB8b8sbh4l3hTtOXv9/5kWesR
FzPGjcayaqqgJHX31S+fAbVcKeFc7V5ezh7LRAofVX7XsFr9jCA4HzsmtcC3kmguxrLYqo+mL4aB
bWS5se4j2iHojnZwPCORMhT/qBkvYUPX2YQlE20zauoGqoxT3cWCOd50LvRj3/t4Q0vQj2IJ4/si
4vIgiRf+9nZGzunAYYtYiRma8O0BixgeheF9FujfeFDE7zoSpCbT/umG4Fr7OTbdyp3eP5sprTOH
HF8el9K0S48uuuFiWUUt19QLLYc3qqTzhPvpjaElr3cKEArGyEmJ8/ISRyyTk1MfR3vSmp5yMuwQ
oPwC7s50pH5Rvm6r+XP9+Kw4ZzxVac1sFRMd7JgiHIEtNhq8Nwd9oOOepk/+y8LsHxSFaLMt3d4r
F4N6ZSGBBAAjCi6McNe9RbKVxhAY8WZjEEkpqfODNpfgkOdWZvn39/ZqshP8yfZrkMtapocPpPX1
JV/Y9q1kd4FL3tc0gQtVCsBTpeeryjx+pzXIOYkV67quR/hqzGHvzs6fAxitE5ZOjbmQr3gCc4Qe
JLTlaIX3nrSNDcheqoW5sN2cmuHDxAIe9W/79Df6TvPAHStM1pWTiWbzAAk91qA5XeQT1ITG50VC
gYDFEux4/7pSPgOiVUuEv5LPnIqMFpx7mA1Z+8mY9vbgH9RF/RxlVn/q4sUc0ok9nojqnDLz/O5v
KLE6g1YE7vyPUm/CRIfxH7N9T875c/7Q/ira+Eiuyo5d5K0SouuYogasa7gIhmkBUQ8KQn21uHFu
uBXEN57K+4T6R/VKEH9QBo0+NnK7hC9rsflVXZSe8TGciNuAUkwYgYbX8TFcABD8NBZJiJgks/HK
xNzdVexHSJBGdZilnb9wlIC/qUqmsJE6kmXpPbRQ/jHL+PnydframeHCOnfgEXRtzhWfUALwImkf
Rp19QynEq8SU3sV8nG9DL4PI6t4J9fVSs3+HvPP5mP4Q9P+tX+12u/Fzh1JeJm37GuORNlTifmYJ
RH/yPkg1jVSpWV31/KjljeF4b/Xq/A+eak4nc7hoJPLuB/qdF7Zvz2AxAE7mLP81PZCtEE6RVgHI
KA9cyfDaonmtzRHNTJEMknHHxOglUwxxESIpS6J8y5kcmO70PukA5so0uWVZ59xXCsdsCZOxG1FG
HaN8NspeyyKhz4h7ieJGdLu7YPiy6yjaDZQL95ykhqpBl4ZOB3VY1MgOX9k2E9ni8+/YoJmj3SF1
vBnr6tY9FHFp89qEEVbiXXB6wvVOEP46Uy3ggtKeorEU4pdbSvgiP6tles/CplsoLWhBhkQZSrB3
c+dLLLgzeQd7G1lAzhQgxwAL6AVzbA53AsXSqrU7WiZiVnB1NJyqrbvnCXcYR9x+HSGIBl0EPAf3
JsPunoPqdvRXUAjh2umS2b8csx3jhZRx3qZZ+Dsnn8YGtVqikedJ1sgCwsu095vOSapvOkHqnW86
FGnttFPEeXZe5s0/Y2se4MX0kF+3HoT68sqLwYNj62Dqn2rMFVxODJ+G++jN1EUqNIjcYycfqSlW
7FczpQgT9L+sWjAcmssXAY18ej7H92/xkNRRdPJ+yTwoxVkXvGRcf6Aif1JP9APLlVzKbP5pr294
Jq9Oq+Tm/LI4ZLtSZ+ZtJf9WG4JdpSA9pvDf8l0qM3qZysXOHnG+/yjbWHNtIv6mSl1gWpYJOVU4
LbQ4n1a4jLrzvDjv9rZrkrZ2CXZ/W1No75y7mA06OFWSUKJk4Gz+JfjMSXiEkkToW5H5q5yG7jYz
DdlkQDjjFV0LXGe3NtiC8CrDFiF5NCYQQ0qlVsaHbKbaCGzzafCJP+BEjUQKOqEXN+3uZiaixVEM
e9uoXCrWsFqJ4qVBtsC4Qr0GNZUzE3jPoSPyzmxBRSnfVB0hrvJKXhO9BbWP3aJupaqhpkoCwfTq
QbnVUHgLNZ+ZA5aQEhdXSW25B/YfKoONNRS2g0Lrldm99FnJJgNG2+WrBtzyoMrpPaLJYNgZOENJ
2bx3V457XeGDErxCcGURJND2tmFdNNstixw9BV/NFoVyVl3BxBtqA+O6sKp9z8saQVpCHv8pBvCE
px4n0N+3mi60X2ULPLMA2Wo2dZEsHg5c9DA6z37dFOt/Wyg16jENkBWvuJY6SA2tdGUr6+zSFB+k
raD7V8p8lEe0vM86m1Fiptxfx6Q+XDus21H/snj7MkU+VIO6fPkLGg94RsmK+aBoxkz8QsQljQMw
jtQGBCX0l5cBK8o0BXCmsImRAXlEKhH4EkX2AL4e+T5Mzl2Vgl771XZmRWQ+MQFM//Q0494QuXJr
FWPPiftK0/p+RuToRF3UEUkdnSi6/UNAYoMgSSh+KnXogcl3EzgR8QF0CDh9/GbPUACMq47E+4hV
dufGpQ5clHkEYx5R0DT6FuZonw9DetsNPflcTWAmJ65DXY/CZTJkkLgUQPDijgUNLddDDb0J3wDe
IroX9Qhy24NQ7YErjCfKbHTigGd4Z1KTz2MH3IDG12shfLEsRkUqtTMaInigGtOdxmGABplg2Yf9
6k/3SF+dp8h3+CYJcsYA6qk/Uy0F/4b6DxPwt63CsdCq0YzFO76fy+CKdPXejy3HD4h4OiTHIEyX
A0NefM4yioFzBRDfE2QU+IunmyBWs5nxftmquCGyfAlviyZRKbjeaPc/85H+5KHgE6ifZ8uzwsPA
ZOVjUgRezQ+xfWj6Pu39sIfATFe/pe0nzQR5m58gPrzJ/3VqcRaiXM+iYc16C/IsD21+IDAM2e70
bRcTtpUHdcCyp8W/mFFkRZRB4t7unOd17z6Gr+o0EkmZCGwYCt8Rdfn3jVLMtGomUriWGQvaWv6G
uNUqWddla24rMB2PaC/QEJF9Keac72/dazreocwBW6x3cT/yce1sgZkxA4ob1wPsGNtvKdOR5twW
p6q8AJQwtMf3Y4KKGuQCrnVWVhb4i+5VkG57WWG4pPlsaVasdENvQhAY9L/4nm2A/NOcu/VjYdVo
Jep0GhWrolglY99nICkooDEUe/Emo/FRszxqGdR1sNpithg60vB10KfvzDeVfYXUz0qaGcVPcmSw
nYRl2EiCITjwGeRWsD48ttOQ3t5oJ/BRZ57ninG6hkBaKpNK25Ty+JnkGYRo25xlPmRpsoMR/HQn
acJHOtD0DjiqkLgQRP6UV3QhYaNq1qj4g81VnMa9SEzqOLc81IjbdHffkIMFU6gCcm5eJkHJxnpn
rDjMPN47XxRdTpCQdl6s9Kd0yy6zpC/p2tT97KTLXgaqlr3k5W0tvL3iRvIOAbnQzvCYoPMa7FLz
IDB8DckcwCXWpXWcLAcXtv6jjrGWk5MKcXfj+8K2YaO+abLUIUwQXRoE0DTd1Y6bWFK0JK8+QYKJ
0B+s8T+03AaOVfTtf+kxtANMAC+jeNlNYgUfv2pKEsKvIyxmw8ZSYgExPdhl7e1DCk/HQWJV2xfZ
H638owBwEab15JQzYqOs7Pi4qllr+I97JMDBXU8G8xhpklHc3R5pZhkusOAlk7cri12pzVC2C7js
IXBpM3WJnWrs5nXXMigbK5FDLMh3nlawojcMenaICyQXbJ0E/eGeBMWjTCNXvM5AC6mVjyEOe8st
ZWENzS+Zfrnddej50izU+TqNI9hSdiNgQNrGusvkpkbpVr/yRnbOxQXF50yeRgsE+NTB4AaLJWtU
esUiIeU2CqhLmusqVLybibdG6qS/tUnI9Co63mBFza3HkdaGP8KdBJYuoO9cg62DEjVPT3pIEGYb
YMY8Xq5RMWxs4jAUcpjGfxK7J9M4rQ9hbIgbhpLy+B0+ULrtYe0x5oiux0AiWC7NfBLj4JtwbKqP
Fg/drz4jEa4io8YFq41cWjmB3d4CllSR7dRqgQq4HsIMnCPd6oVmSAwFLf+UmK6ebC1afNXNWlko
uiG5prOLDAW5sECDnT9DEg3fvheZD82fCLTmj6vhe/dcnuaSbJ3oHCKzFWnoa49DVCkPd0p+8ijs
HET34nTDgMFA0XsatsSGHxm3rcr7yAK66VwdNNr1R7w559VOEU/oiFPVvGhNY6XuqlNTUvs1QH1v
5C1Wd8412pwfyou3c7tV8UnD1x09am7kXYzcO0n3196+jN9FkLzLQnK2JDmp6k9viuZjfjZI8E3N
dP36jsKRZuOH7ZHwgjuDvDx8WLNlzbORcos6HsCdUrXX7I0LzDjy0DkS8koLdclCzIGjzB7v3x/y
YJnEAq89dRTsLfd6QesQiNuAqETpg79I3QHM8z50/HedUEBW3G4iWvsQmrbNe7AWJGITdKmoHf32
oE7wa4vkAqlU5UaO8enEH4FY4/JLGBn8I3Q6A/+g09Mi1xnEBJNBwOqnxTa9JvwsR4x8dWrb0bmV
UMHr2u6sxAxcbEMNTclDHawTf0wyQy61A1QI0G1JbX2fLs1QznlU22fVjaF9Mq4S14VBY7A4dn/V
eoCqgCdfSrPRbv5ztYRJK+AGsHWF3w1cWj6K0cacinr4CekL+lhERWKC5L6Ioi1b9ubsI+CgxcX9
g1A80V87cBv4l/ClUbO+NjSdje/cMODHZJwdMcDhskGnnrLTBer3+6mKHc0zT2GvvI3Zm7zYO/VB
sWfaSwE5DZpgCzG7JpVPq0MhX5bmK1AjFfwlnl9qS5dxVsxFwuxiCbg0byLaJqas7zz9Ik0nJa5h
ZTDHXzvIzq63Cudn41FnbXVVlSNnPrSdGV4LCQeG7n7eeI/dXc/jxlDiUEr+Qu5dRT4ntJFMrAVY
T5mEnDC7ZYBJPxbs4YEGHXUUsLw/SGOFdvyJESVRIeeHpt70+yw7xp8mmGB97MWYAX1V+FnC0W+F
rKnc91XTcgf3Km8Ojo811TEkAM3CGI38+tGzLGoY5u3avYx1jswtI7j8i1WmevJkK1h+I7SPLCFH
qjX5QL6DMzhtoyPsa5u0tHuUCGEyd5qCJqKoPp3Y3KYCwL8mjXwedx0ZeOM7XMvzXbKPSxoaKwGX
OHf5KenRNx0klAK/dBjXAVlwk6I0GRBYswLMhmA7thru3FDVKssTRCOzh7U4PylJ+9QdLG/nMo0B
Ah3wDZ54/tsIyZqtpFadwxJi7Fdck2La0P3qCB6BbZldMri6xrT1DmBB1Aw5vfuDINf36vyXYY0m
OY38OmNzm7Tg/J4ih61x6X6SeA8B+vd60p713FKfvH8YoDXDZGQHoIGnbhmvSm4zJj+VQvEDNq/y
8j5YL8tM2qPfwSrfN/Y/m5FyYia+UVFyt/PLXDT+wcdi0MFfB+NoYrrQK3KXo54LVTbHeyrvqRM2
VMMMsk7vMkMIrT3yL+N1TVl1eEN36J0v2edhktf8Sl1DPfno267lNmuaryIuQoQPvi6+ADnGSLyg
AnTb/dQJuIrQhREZEuAgxtOPsHeFxd23GrVpMYl/wacFBF+SfiKjTDxOipXSJwapxco5C5f5Ul28
MxtItgYk9Zw5Ek2YxV9FgJiy0LUnls0MnxvRS7QbevxU/nQ6D6VmZ4rARs6ro6at+opvdCaADsNa
eWn1LUhzVx73bl0V5CThvgMrRBeQoiaEiPygRKHeJnstn0AKfRfjsw/27QFU/NvDW3VYCW6NX7rJ
YPpRI6ENXfS6SlkgUP1MZu/yzbc+MIuBTWmD3wSFAPhB9G6jqVHnhaFhEQ0W311S1JBkAKCZ24cN
UoOE72ndSwKcNobOPehuaWYhCBGvWCcId4RQ7fPt1ya4z+8/6P/UEZL2XsWR5ESqifg09g6w2cWT
CNoVIrBHPfOhpXpn73l2NruvnkjdgE86ZW9brLIuk24+pEqPktj0LwcA2qYWynGiejboE3oZkff4
bTEZOmtwTEvqwa0HDhTJSsSGKPScAFKVQHopJEx/JWXu+gsNUjLD72+nxy/MwoUV4fVBtUDrOt0Y
gAsoqgmgZze6R6lIKnH17iuJz9d7rfnn8QJAuBZW8ylhGMS77rCCzUZEust9hn1paoMjFGHSSpW3
C9lO29hPSzavAWHkZnweZ3ZheFwN868oUbbDS9Uv7qMJSo7WuiK0UlebxT/a3QFtJIskDg3myQxK
thz1iqJg6gVjPFvtgTJN0eky3vZ/2wjwcOzaKH/3r+CmabvsvpXyxO65EwAKbv04c1L+incoZ+oC
5DFA9X41Kn+8zgE/wp3KL8t09329IziPBUN8qFsH5vYyymgsDnzbnBWLn2Rh2KaG6hGL3cbJH9wz
K+oLXd7ktwu3ojwybSwjqStDjF21Dss6o47FHof5tP3o1alGGwbGZQ/BjIJPXobsSSUU3s2jyLwj
/omZjYO3R70CMicPAIsiuY6uQST1tWNbp8n0JAEsjQTKaeHw2WvSN9FGWlIJb+3HoON+kDqpFr2z
Li8V8EA+r+viCbudi8KnMjk+74HEUqZu2fIvmnBkWC30Ckzyu4pBSl5SH8e7aKTVve1rPY6O+drk
KRbpBUWe4b/VXXIJh+N6DEN0e9Nrhm3Is261wyzkfIl4FaMGfhGeDfCem4NsDamyPHpNisN0PEk0
UYcbqMMzRARzqRxbJqqOC1bCFD4OIp8Rki9Hn7yjUsMbTX7rxFFvFNcrTEnCRx/S6nQUDw2KeNDd
kUiJCGVXkITlInDOvUQOjIB9wbDaOneAbOgKOAj3cuDKxuhMU58P1+RdHnOGijulDWZckubxLFRn
cG9NX3IIz3hIiT/ce7JNjLNyOUMQqpw5Bcmo60kkn8dbxtDIgwrp2ag+GjOCh7hQEsk9DF7P3G/i
0MY7c1rihg3ChZVzU2Iwxkltigg2cMaFnyWlfqA1tvzodvc/Vv4lFia1XTFyeu5PysQA6UxDKjtr
MKoc+IMUM8BPjBJ8ML1BMm/srjMxWXxGAOxdv2LxlYtYEh611S2ArWlvn6Zvx+gmcwjFOZMjNJKI
XmNTJrSAdKP3gRFNZthZlyPYVHngUMSHLx1ha4L/Gy8RGkNKbI0ul3NMM0zMdTFfTahQI8mdDr8Q
Qng/1HufPrt8dlSZfhpRg1RyoWtaHUVu5MYtsVNMuIIzFmrB5GTEXcvbOaF4c7Za8vjK/U99irlA
vMT/vgdUI4NArMbhHaYImwXogOcrjbwRPBxA+XmPNRSChfV6AcBlAow7g3eD7U00SuEwdqBReaUW
blkP2PT3tVG6l1rs869LWd3WtnCjHvzbtLapZxQEVIBhZkrmfv+bKnrRs3xWmWUKx2warpXNCWNZ
YC/PC4UnJVxO3yYCMpZG5Wy6WiNKqUD7Cf2orVaVsWFwQ7FfY+KuaKlrJOPswmKD/LIoa0gCU0S/
NlIAXNckct5XzSmf6mIhCTyT3n4nIVB6LG+dp+WNVind+jxisYKeRtCLyRq9dHtYYz0R5P6hJViM
EhgH2F2AHkFLIn8cQINeFT/xsV0XS0MD6Y7192r8NDeIJtDWhC4u+XhmDPjwv1xmbzsaavy80dpH
Ky+GKxKVRb8bF7fxxvGwzdEfxqGiQtKdCqfuxV93l0mEV9RVVzHxXpJ4rF2xSFQJm9pYvf34++AR
lxIpPBh21Q4REOXGeb9oY65X3zv96T6SrJJHkNX/yg0LBcYN7L8gs7khDk2DpEGObT2G9tSRY2nh
gvbx/X1s2ZU+vacH6wfT0tgKVj/kvJv7DNUGWvzJABG1t/YthaNDZOO48JMESdTdAz5HI5nG97hV
LYhohox4RjJWoXjmZ+0gB5c92/aZzGiTM2btuSwlgX4az2GJwYbYScRD0sHTGOgIG7YDtVVq2OaU
GGwRkVA1/DCHiT9zPpqkW85IkJvRaQjNWfS1aU1MxAv7qJsV8xMFEXZNbQKhPBQT7iI2GQIQNtp4
bxuGFR5gV8No0hR1vRH9fBkqJe1T5zJDLXhakVsTxUSp/NaIqEyFhK2Zx9RBCmIzZ02/4XvktKTx
CTfChbxgc59AXMKzg+rtPf7Wdubp/1JZqZPl/mh/bDrzrSDT3E5MVOQKB93waibJc4771aliZpoq
MoBnyp4L1pZOgiSrB+cxHqrHEOnIC8gbCCwPiXVCWw/YC4cELKNR4GfV1xIp5euJQgE2ROVxSH63
8rRlfiEITD8b9H5wPChIkEFalMvAs8qstoNT8iiCX/ZFSg5i/laFoFOPq8dADpo70RsjBIy+wKOF
jgExYivzAiZmAJkaJT+W8fQwtVj6azgHoZRsXdm9EWo9XX2VjmZlxRunoH+uVKf1CC54wU69DT1U
MT7mMj80RHEVz4Sq1cNvXxh7G4oZ1QymnQmvT5BTQWje/7Mf0qOwVA0QxrlCicpr43Eu+Vn9Apd4
uq18jubTBTEncxqg7Re9Xtd2rIlZghQ1kY1HKd6Ao8jjDMD/BBhmEI70rv+vtj59+lnkFen0O3M2
giPTymYmefpLsb6JYppggJzVzPjuuGkh2yXCZPMlh3DBdP3mroZ2cvTl/uI3VYJ6IcFgwm0c0LFi
qR7IJIHugSbtTkQ75n54/oL+lr/R96OLxdL23UGvNpDuwwPz2zLmUrgAeTXVV6L8DwQOvp6FzZxV
FIFwmp4eYn4eI2fySbQo6DVlMO/NRNe2PcwcYBYqUFJ4MeU5N9t64vx9pBPqsiiFDlvAD+j33Hh9
OaulD+WbOzm21+TU3jwK2v8pZYbEQvSAxhzRADgKtFzT0oWT6zQ+xSss1gYAPpB7PzjGif6tnyJf
x+ENcREj5PtRoeC0vhkJqwlXUGeMTIY18Rtc1SE3FqlLa98s92+4goIZiC5dIiyw0HUuK0/+cQEc
kfkQgilAzj0N/cIG0fc2X9n/336ew4SsSYKeEd8/5vWi5yoY3MvSELC5LQzppcsxpD/KkbqMzNtE
QJ7g4vYCV4Ci2IqIWnNeT0gqsGHXkuNW1NM8s29kl+mOA4+hEVncLMD4ao1gU7dros8C1S8qEl6X
BwuirAK+f2cpBGhydYHFLhfVkLmbSVmUG5lXkUTuuSUWcGRkBcir/O/HE6m6A0B3SJdMDzeBwuQH
IrnDlzupsMxZ2A9B6P9tNcwbFGBn7pm6DpgQW8LBbug7hWdYFFb9bjpaB3twFaBkinuMBujxsXNA
PV+KUxvH+8Wp/4pxAKB7GVP53Fr3+q7Q9YpsD/gYn8ZaSHMRctwy2kCCPcitDQnNJYLfQn2REJdI
e2P+0TQzrupSNklCt2s5jQWB+IKmyFXXEBzx2EdHa6v8xnllq5mYbnijD89gcgnFzEqsfMMKZVAj
vtqZDxad+ycoBkdreHJ0ESdPSuTwUwvU+mGfOoTy2xor9C6ox9CQ2dbugsFzQfGU0kagqnNfCgzw
Rj8fexWvVyeDjCVMXtCPTq+rE9f6svOmKegmtCiRP+Ij4nBn/axkgddTa7jc4KTU/1f3IIAlcOQ+
QPa6aYAobjN12vMdlReXmY8XtOYzZd4R1ObvDZtxqJ5D5v+Qxh03e3RM6yux3WqcR22yD6B+WFra
MkIhtSOFwOqw2Wc2mN5K/qaCr19ImfYy4987T7dbwJDTc5QOIpxpzgx3XalFY/braenU3f7Yf6OK
VLYcDKoIVRS7vcTl3iwTOTNT/z3oONmXUJtGljNlD/ylycu/pLiGPTe5h05ebdLprrzK7/H3T2Hn
gWDJfJAKFiwtHE7fPSEfa6V/xs0Iovd9rFkDYWKqk4/1Tgc5BOe6pKxdHRzuqI+B7dwUyQqGlBug
SDEoxXFdtHSl2TQaRu/rOllPWNlg+9BbUjmb2YB21rZRq38DwYrMT9JG9k5ULpJSi+pzZKMffyqU
uAsX4BKvr+NeSGeb/+oEeeIyijG0aSMMJpemhkivoCaU1/f17CqCTiYed3ETwb+kITu1d9BwS1YO
IKHiwwee9kFK9trL8Tvs14tIQcaNsEMP48jtg8jPvZIsS6/5VzDAJ89hP4GQIvAEwkhYH21WfDu9
0o78Z0WD3Daw7rOIbw0aU/2CWcMGY0vaZnBKieZ0wL5ZcWsAKCybhONWCfpQ8Er7UWEkpv3yE2AO
60BMlg/OobeWzHnrDrUfR6ap4icTawN+UJKfQ9SWUAZN24CaXUFdoSL9jVYxXa5EW0kReBRqYI/A
JIScSk07nYjhNDSi/yPb2bKr3NRSotc6GhfA8HYajvlKei1gcapiN9Hoq4bfbr95xpRHUMOsdqrY
N/klac5jFG2S74La/ZXSQiZMUsVMndZPZuAPxt3wAS4QUDGpVBnVFoeCtluBER1HjlGX6G3WhwE0
6BWJH7nG1Kpi9/1N4OjoD9tNbuvFjwd9pIcM73vAJy67z3GMYflX/hmlb/lLry5aoqyhUWQknLFf
LeNX0WSqFaBMsh9XXWnT8iQoKcMI7f8/EFjeVGja+Kzru1WTw/DpHuC1bQYJCi81WuX4bRGTgf0F
E+CjV0ay+E4jCtaFNdODOwvNQ7ODx2NnTBuMp4Sn3iY2giLd190qrdxDllMLqNxZTyz9oiS+esCz
T6U1qmB6o5o0kRNH8NLI/hlS4Hn494RIU2dergYwzwlqW8wGYSYdHwRMjLr5N6MUnfY0abLwlAlz
Qf+hHSefkHZnuodgvtlgoegtK1Nz7A/Wd1AVOB2YdMJYxFa+e7R6XBSe8gDozs51auH0B1GAUhyI
69Mx/wEwaq1dyP/FQXXRjv+1xvk+dg9aFHRhHpDsD5LfJ8zfExJlX3uisdbIb1rC/07INr7nZ7xy
ReLePGc2D0Am6sRkPx9OTubX2no7bn4I7CROy2LGtIP7AL8F7U2/ua6yhN5gJcP0Mj+IP9fb7F7Y
WQksAmOm7qSDOsvHBs9q2Anly2caqSd4oBwA1nDNmkVKlA+7YyPIqzHLKv9Qd+9l90nUrJsUrstc
maXwWcmtOuf0e4c2+y8Zxrl6YjsqVQtntrVCng+gyww9xvZltd/I6ZAGWU/HpG2lodwWVfxPZw/c
QrLxzSLruDiohYd73alwzvubeMESNnpDtJz+AqLOeQiHvFxtZ8rDXKA6b8wYnywWA/IGISB31yKr
VML921/qIt/FY/KZk9C8ypgVd1Y/TzBppl+O14y47FbFBT9iE3Y+x6vCD1tmSIVc+5Be696eSNUW
V7/PPgNDClhddWyAIyITYMHrxtZuXl6u9onPefQDX+KRb3n6Nt5wYvGYAP0IUNtFa4GRtJ8KbPuH
+Hre+ZyKejxUDH5NxTDwjlw+tKuzqwePSnZltGdv+611XeheOgGKLEddZ3X+2/ttiRiYTza1W8PQ
pM8p3SQtYKh4Kf8TRQIJ7oSknt3fgS8vk8OUQmTHbcOSI75wHNELJuBT0vKL83QzLmeaMtQK0u/2
MNGoFy4MveQk32nWvNaHsWrJxTF0qDRILLsTlyEhQKFcMJXbRv08SpaKVSeLys3+ybM00CBRJ0Ee
IhwGT7rkhuZEAUwaXX6o2woDdgvix9VFFJi4IeXgN7FrDTKPGp4TB58x3GV1GKnhyu7TDmhDdk6a
DPEGWFlnX3HORvrqug2L7kNFUUIyNSJ23uyJ8425pker8EJzCxrGefLHMATpYFXeTpvhG95E/Qn9
+gb18i94MZ+eafT43aqfQ4sc1oY9W7qoxQFHmkb2/L5iOuF7fdfgSyGBoZj0MtX/0oR0d6GKU/Sv
etpglfXFwnr3qNbbdFBbMAerSPrSouUJXI1W6NBXOujrK2uXKPoqKuFNFjHPfkHeJ/ChnOfjPcMr
KZoPPXTUSpbfhAdQXs3fkc9vDQZXOZ+30IWlgEuEnejcQQVWOmTdgF9i1fQEoiw38O79Iu15DBlD
FJnAVz8blXEJTVjhr8QnswGwFmsk10arKL9HzJD3u4BXQPs/GjHiw6Mjti3vMa6YWhYQCneuL+BN
qUc0kErtUgSH5STfe3OynT0esjS8OdFCOga+vykRg8QXo1DWaUfhDb8e1aQTNvvyZiSEt9Jd6WbB
LzEVJ6VWeTlrv7m/QzIBiLydWeRLdKv22/Tm+3RiyROJs690ujoiYQqe+gWaLwKWQDW5g90R3Wkm
B16fYhHYeTS9cw/CTRszqti56IZtk+RBkWvLOBrfn7ZUzlCT1VTTKWaF8NUYviGRoZ6KrVhw2xap
BE60KcMy1nkicv7WWGBz9kLn/ySdz4BzJ8MWftF309W2k7Yho2KwGsuB4VRsLy6lhp+kvG/sBn4B
T0HwIFQg765yJcoKwc6Sr9Gqja0+7Y2EkdIwsnUdWJYcRXX9cUA02OudYJ2t01UfaMyAlXsXWRgP
U6DCi8/Ho6Uc5ldI6I3yRmn99LmPQlJ0TxAp3c87Op9h6fg6lE7qtiT0DSnVqkLroajIYu07/4kw
kty02IEoFibSTCvwE4uG9TaeEloiS/8pKbVapsCKobdY/KeYnIMZVU14le7Pkm0En3gtqI+k+IQx
RRj4jl22hINiNFgZCJSlbmA7RwNqpuHW9O7CzVVrRn8itYSZYTz+vlRZ/tztds4St+dUwy8wXCUK
KD6P212dItrt6RaP/koP3+DfmBv1grS2RedPz2Bye521kshMZ961l0Ybg93Jk95KW48rX+DPItfR
co3d8ZYw2qeZz0oGdp9EhZDLxWs/2adsezI2dEbdyaS5JCiJva1x6S33J/997G7jJUhWdKrHVfyH
Qg/Jm0bKCNPkyG7fdN2qwTQoeN2/fL6GwAUS7rP7LYrynEM+rhDLVfRmMi4WC4GEVMHpWlKafP53
zRLUZCd3tCRTNIiHhE9SZlP5fHeFoPjeSFLaXmmPJrnE5XMWxCmKHsDtRdNB5HtcJH+Nde2LUxBS
oNkDrJ5UnFU1Q0+QBBYNpy3Ne7ItEsbtP48z3jwe41KtmAYDpfrn6hWDFL5fMr8RZA2kJqyq64iE
1FOV/ZWuPnclRNMmp9HVo46zsOqY/sIJuv5fpyHvN7acmBa3U6VC0XUKwi3Udf0LA3A6xKcjJ+Ni
AT9vzkBkiuIxKh2Hcz/Nf/Y7RJQH0JX3T8C9SRw0fKZ8ib4uXzv7Uwte665pU7QLngz5Z6z61X7y
w/ccy/Q0pwAOstIVcecqXPoDVd/oRz79SYOg7M8S1aT/ci7Bv8Qs/XaW9WSplhZwLfYYCDc6vVxZ
vYuzT670nThwtIN7zO5Rxh6LmbxFjM7f5n47QnHe45loD4VGsw6kh7srzqjpWHPJf74ePvH3WxSX
b6LVTHjgx21taX6VA6NsrKUXp4PebQAy9JKApqJNeLSVOx+rSgRqpnBk8XF76iXxYpMcFseYwahO
CkfdozNaPJrco4A3wxCEsoRtzyrvzYaom3KB3yYz9ca4cRQRZqNznOxYPKKEzQjq1hmaioiYqliH
L1aot2hf2POZCLr2TEI2iO/rsdfwrP/qHyWBwPDTLIBjUNcquZWKiHxtJ/saoScDB0bmQfB0I1t3
Ljowb4Hk7Xf+oGjvFszdfm/WG7RD2vL/bFnX6ZOVOkotn9pCJCWK8rgE65UO0T1TzYgGD75DFYje
IkByxWGixuLlHKdhiVU4kgdmkjosMZ/XdctO+4gJDuaMU/tXknoKHL0VGl2xccEp4L9ilTOTpJ7y
pM/z/J4nhP2SlxK17qRDEezPNSAKGqpgr0I+o21KgmtqAevELulrUY2V67zNPDwHOpBPDBvnqtka
T+32jodV/bj7XKzeffYr1b+pjaiSFKaUsUZxdAI8g0J0dF3gxHHgAsW6ne5xeNl9Ei+68K6xvoYm
qR929rqvunA5QUD1IylopkLDlt53Rmbg1luGb3tKkjNWOXlr0GLiLZgfFdyKmGoaJuLCcqfcmbd5
QVsIxCsWB16ycN78N8wlVeJQYbBM0B7pmgM8Obagb0dSjfBqwTJsBRCggcbyYgSZulfKfGx9baoD
hDojWJuSAKZxWrZS6TVcSRBQk1GP+PshEQutoV4aOWHigYIBZSHnVi7joyisElClXgUlvOukNorb
bSKXYt8dbe+vsziIVE4+xuocwQo52GyVV9yTVgzJAT3kIU/U5IR9nKarzZdfpFUNZog5EekjojvJ
lb4njgJE+AW19/WP0UnrRJjSe8a1o00c4qjZY0K8pEWqGO8ypVSpgpz4ke8lGQ16qoPa1HU7PZrP
rCZnF1thg+tbvuNeK2/oRNr3e/0YrdcwtxDIHAwH4KmgnvI80+RM5MrXnPc2J+7tCnA0xgohIF4z
01D5ulphH8tQLVS+U7zOMwnXSjd1dFtDv8sBETzYunZls9YsWpDTFEbHXhEQJxinPrmTVInrh8Nj
XJy9kGT3cxD7PUBMwmf/NGQuRChEMNEy2KCN8GWjmBcKIeTdXNs1FCUHZFIV2J/ThErKDO6CZ9Bh
KP9Wz1MzKRgUlwe3d95A6+9SZThp6gR1LuOyIPePv/TzVduzgIDD6+QwVjbTtXk/znU8vCAa7tl3
UNRmj7ATewKjf19/YBWP9T4a3XSIRGDn/VjelRLHBuLHI3lMR3Xkaq+VzgK5IC2doJA8Lv9GFp18
I87Z4JcvOvQZURHyXDfkEhVRdH9pItbTnpld5KKwoine7ZxM/4FGt9TdJ1iwq/p5vcmdACLlvoW6
3oIcbSh3UJsyOliY9ngMupkDMxxDIJ398l5RjWH364oKmAg7c50ys1kjlt1iBdAmQgfJmOfFGJtw
ypGc6gmr24ZwZxlvJQoKqjHm1MAStIuGsvvHPuLFRAdpWPhYm5U1zX6wx1AzqzFv7EG1mB9Aaxa2
9A4g5hNkM0bKpOs5IxDyng2e9K918tHXoniVpgk0pYhiAHz42WEIgMwvNubMyZI03tio7ICHJ+V4
85dTwyZwKPzocuVRDFj7/oEP2TQa5K5RLl51j+LoEfkbvOUIsWYcN7kt4KwLl327gNg1gfLBpK5L
6ttn/Vo4lpB7j3oKUiIFxTdICCfg/rUxEJDDNtO7TIigFPZfycgAfP24axn7ooOhX602v4YOSDcc
PRDb3mEk/ngy8tqTaJQzHpUBgokgcQ7uWX4+i7FoEj/gBgx7dzi0hqP3DlAynGbx07zYBgXiQQW0
0ogBqfTVcaTsLKDbodRpTisvkAckq/i2jaJ89dWKM7vx8lNliF7akZvKTHJqVd7+AM+/jkR1rcGy
/rmVp03bYa60gBTO+lkkfmuq+cIFZ8suEp0U62g2eBZL8Rd7lVc0Qx/Ks090kvfrCeNWLUO35dR5
pqPdUKia3C6d7SJDCJS0Uu7XZl9MTepoyAqnV2+Q0KSAaowNkzNdjucQX0Vfz0LYVWg9s8AhRNpS
FdKEBYP7hO0sJs2dzcXlVs3Dzr2DPhp2Wdeb7kL55U61e2NzlJvovulwZ4G9FngmoSY9FDI48eHv
K0U+RljbsLVVBwJjmp6XRIWfBDbOdF6RSJgafZEVE2nmlUd7W97TAC8bRvFKIHDfqkMfOsPKQUwi
GFUiZ8VJUh/nVRYI3jqNn92ducywtWH4M+UmGLhUu+JJXqsGqJn3PLhvcI2Yn6dd30BcaSywa6sd
rZIdVaP3m9XLp+C86yyaM2KHEGFXCplc1TDU6C6nAKW6vBiYUnFmfJanG+pYu/GFahxpPXXFlBMC
M2S1m3b4nMmef0f7KTnb2suMMcY5mRP7UjgUXxo4vUlpmZfU5u23lC2Y49cXLMDrs/DyhH5J+5/Q
aY38dCco5vMJazVwRJae1SFGr9//RHSoPgwPCbMQJUbhn8ztwxVZBcJbq9VCpvKYPzGMOozi/Bfs
oa99njCRMuTiZicqQ0OcCNxt6eTG9tpxZADDHIg0AFDL5cPubJgAVP+v2rbH9vJ2VCoXuNsbicES
js0QFuuC8U0TZ72XE1X7FrdF0K82QEkxGpcfJckvl8zQcWOROIurGtM3Cm88Xe4TgrrbRzJDw1ts
Uip236TIzsqEmKmsuP6fiGPJkQ9W8ZXcK5E2V9DS9w2YwmC37/zG32BkDNB3jE1g9DfMItyxDMxd
LhtKObzYR2hTIkGmWlLqAeuMU6cfkz9JsnBo7XNHVcirRyvGnapvoJpcLvtGPRmJWGwe5uRABmI7
Q7+28/U8wyb51IdVLlj3ta/sClnjJBWvU+kII9BwmEBD9E1C6XGe4THNAvE6OTjyJBxf6wLesIRJ
xFpXIXDK2EEIqs0AgJy0GInEGM2VbURfvd0+mVylmhQfFIjKztP0L4DbyyxhPZ2BHnNE7AY3FZ4A
b+utRdJA09opn6HVpEma88DjnfCPhkyuriCb6AYzN+FfBEIEGGBTcxK1XUMfBgo2ylEzSjm7WH8G
Q6Dga9WLxuWG3TN9aeHxpAi+rRTAP3Hg4cxMX3TwWlaSOGZnbPXEtlxbtlyqlMuUL/9mquwdOgsn
yt8PHpEV+t7vkH+BAdStywS/Wh0po8qN3tFc+vS7jkDi25HIPNmi4u8D31i3eIbSrKSkmRKEdBpP
++0IYGePIUNKm1RMJySDC/uqa5LcV3NcKMadVNcJbetR6Shz0gCAH7BRinl7v49MikkRaIossI65
Je9O2ARCnwUsZzaAhryozyQPeKvLsiFsEJa4L/gzXMtYlqxZIhIa/h+alMpDnDpu58MqgVGlRfOk
Ass23w+iY2ZSfmk2DYaleK+D3ivJEgGG2WHyNEbUwqKCJGA3Xv8O3+hHTv81wq1MU4wQiJFseLBI
nd8FWMrVBKH5vQqZ3wiO3B43QhgZ7jZpZlIaKQ6irL4ZMWjMQfHv+m7H49i9UEKo8rKzEecfpXPS
CZHm3Ni3nIGt6q7muyyNi3PNiGKdwCPyH0CcGyFEXziE0DbcaabSTqmhKVe1sg7IvmfUIsDMoIwi
sLQuhjOIEqBizTvp7311Pd4Sj7aGTbO/h3NBwBvrH4xFO1Q8nHWesUw/+wknjCLmcmVn7VxPGwxq
jrDYxMVmWy+gKf7FO1vdEP+oJbLR6vz42tDnbhCtwcf1z2hHhorL8yO+j3KMOcfsDV6t/P1OzFe1
uln9p4Qk+8L2WmkSUnlMnXfLyIoGu2TgJ+RgZHnZwng4pHCFbKaGvkndHfYAuYE+ufmwDNH7q/EO
NOyVB9mEKHVkHNlV045S9XGqgMHO6HREc4kczHTNpuNUt0sWEJFwbI+X/6VITVGyznTsjctuQ+BM
yMhnc6SMadgplvy95hNgL4kI0CO6JJTv6X3cu9lUOdLWDZeqDfM1CRNPJztMiu9yiCNjIXoZS8Yw
EhND92Uduax7YkBmGfPz2mt/17/+MBwUHDDHXp4UBfG+nF+smKMylrqUBJufLx0mnrqtK5Wv8Y/0
0Q+4Ke2A87buooRdtIHal9+lLMjad0pPKtXD4gsIYTLHITyNKkdHW/RDVlBBUaQUTSnxFdSs2vGC
+xe3Zc/jSJ6wpd3B13GCxWl+XdSpotswEM5QX78qesRoraPMh35CsNxheCUCB9FL6RkLWpQrMYRT
DBJvTWGvA4cBx8ZNFNe7q14Jtyp7CiqKBpfofZYc8i1MN/iMQth08U5iyp7iNWsw9IlwLAfEhFr9
vQ36mpPpKaPyXjrWpDAsZgoC7XDQodlRSzOvEPIvRqmr9UAuD/U6lz/Wj5vGj2v+aas7uf45dZNL
LYFZyx4tAaVSrR+irrKZ7GhdlSW/EWbtL0hbTDDUvNb4x2cLwrokfbIMBirOs+ewUse7tCBSseKl
b0/TDCKKlAwGiBm1EvvZ/Z0iXBovy8Mjvra8a8EUq5Md2jF2AMfJXnhHDQ/bG9qr0qAs0KjHwxfE
HXcr+J2uwLkcohvW7euU5yCp2xUX/BauFtUEkbe8pA3NFdnWpXR7+8fjHSf9m9q+9jAjNieZpEcv
ZA+vG4P2rG3xFcW/0u7FudwPf91WDu8RwiX6n4zXJpGU9Q03rmL6Lwy4AeCsMXyxRVfIzkUy684W
Rqpv6q+2eWzvhstvyU+fff5hAadp6ndQAMdiv88pXXtmTn61ZUr8rsGiPi2LyJrU0qOF/OPdn1VO
Hca6cTZLJLHwstU6vB7wRUJFJqZcFgjd1jPS9EuxbMM2bNoDDmrsKzA7L9dF7jwdj/Dks5vngviT
8h467wCF5aGa/IDNdxMMOIrI/QvqBIM8Hk/yS598r9S3aql2S7p8wpj+YRniwvKv0E3kef6SykWe
fqCvIM+GrpGjdrgUouZ/6CfvrPphFAGr6HVskGzBm7IARa29ajTiB5X6QmQOWlRRMNTTzU5QEnN3
t2aX25LWGzfbYpKst6OrykrSr/JnRu7i4p1yhaj4pAkmkT8szqO+xZtX5BWNglW5/Z0FuLIAOjl8
ujgQgu+djefG2JzP6/kEdasAFA5cPZvbA4j0khXA1TLnnLnnLLblbw1++J/GDulP1kOghsNxWQwV
iwWCQ0h68EcCtj6igAZno+BTNQvrP9QwdANIajYdlAZo6TBQS7a57VtlFe31Gdb91Eybb1gn359I
pYl+keWQYedh/1j8ArohPTnEjnyBFkXUgKlSN0xH/hfAjD4LfeLwU+Es170vTqs76EeRAAG5vU9H
YOJmmrj5L2q63DveIRMFDCBA8X2Jof8VrVPxzJC7pNHvzYxOpzdrAe/riRzNMadM9hAfaTTGM+DU
yo8aKls4XJ22PegYFUdPJj9wBhsjKHg/GWRD+FPGhmqeMf44vYu1DqvChTSCfUkbetHQpzw2/evS
vXNVsM6vsCfZmF9rQzNm3/7oisS0oNvNTuFj9hev7pgPTs4o2joE2ZFd4nvklpkKWT4y4ysdDcb6
eM62oQtlhoKd4ole5iYi/vlew7hrUbqNIENmKhvL6PZ3g98OB0GAUQjVK75sxSsqoLBx1ODBFnWy
LwqiDapl1/v2HPrTQ+//DEFB59SREHCzyzls4nk3uq7YZzBrNS8YpNdoyfTJ4mZMhr14CwFpbNMc
11lBuQy/MgNeTICvqhwgjAduEP9bDKxQAV+LJBulBW1J9n+X/khNscF7vSgz2XchYTpO+A364aBE
7YF4fzntcNAHZtWsW95AUDTMRZxy1CvX4ewSDdFVzCISkDlxhmlPQTjD8ujLdHAOswdkP1JnQZnx
6RHSLftKDWyZ7rqCcC31SNFPwWdzvzdNCkdIm3oAUMcfTiXjwYrccbX05wjGHULPPgc2XL7tVsnC
Nmqmj+WXw42Sk9kRi+6L9/m4Pr8biW8kbCUBxnttYOMbdvYSCXL4NMtlXq/t+JedxALuGmb7x9Xa
WdMUJSYnHdPK9XgGZP1+B16Vp9T3vl+cg3YqcCJpNJVVnM5Z8w8sqNgbD1A6EzhBGLasUEC8htOc
J82CJ6UKV3xaaD0+o9zrtCvVbVomYJ11mgSyqctlOtVwR0+CF6rT4JuZBtNQaCYWIF0ckrbM8QY4
BsQxVdAH8RgDV/5s80jhSGYXbFmb0ys3F+ITgmhQstd5RMqnHxnvnIc4d8O4YXYJNnhREzJJYv0V
EPpQtXg0lh1TBtzD0MBcBH+J1zMySVLUDoZOzgK3g3LWAp1CFZrbdoX7f0y+nUH+DKnZbyaEDRrb
DpoY73GPzCMQPIleLBVN3P6KeNhDQZlfBoIbvUIyjjhHh1GS6QMo4pNsFTyiy1bnAoSZgXJUSQm+
bNJFQtupMKHM5gdnzev+eVb5XXo4re7zCyrQmTbKhl745wnFiRwMUMfQVn3hwZEZ3DsCY/ju8iOe
pkb72YjyxQ12XwCtePli5SssTQxn8dld29XwAyhhwTWLBGaXtGJwxvKENs91ZbsmKJKe9rHIRiFi
eY/6hc5NtrNIEZgFeiTaDQWlHnSQhRIdlJCUGmXM53sfpjMwyBTQtQW+PL5iDl2t4Wayi7xDZb0Z
5FUpIY36UR83gJ2U+8qN9XnKAe2ukF44PidwbTiVlA//qkjzKGWXNNXcY/FuGgPySn5RCSl9eYUA
ITxUyeb0dFwGtxn0vSl6YQP1JhRHZOCuQP4wHRWPptaZMDCvNElZ59iYxO/nM6t1XD2GODpGGyer
9oP6ykdcJ/RRZVjvPKqTtcD4tZUcNUdAGid+jx8IkJ2Qu8anueh/aOe6vpMR9SepT/K4v6yUfxIC
OVRBd2Oh76LZkp01tXzTGDRik6tAnXL/bIMCeKdihzianqOYulBMeCAx00L9SAR/09iHg1vEuBmg
WOvMkDd4P22/BNQ/nkdKdQRBTuPIkVg2bX0O96CjzYQk9stJWBOdGhy5p4A3aendYrZattXNKHr0
bUWCPfuBkES7ryAiOS6LDrcwDSfHEQjXC0T7xLVEPBRu5E+CT/RuTDFtMSBKM/NpV/gV9wvCBVAd
tC96o2iDqWCGs0doOy9ET2NdqHdEya4GduD8FaGhpOIpPYszi8I0QchEEWnJHZ6j/K2nyW+J25fo
3P9fAeekgESgR/Zt0Lwm0dS3wmMrdU0rFu+5i+JjYXTWFD8NQM1a9GaEVrKRpwhIEc+04jEw6X4G
4YdYjhWyDip1G67kFR+/tMsCFBD1MbGpaFpTtWScbo3qb9o6CEknDuhzhQ9Jclh+kQVk19ayqtnx
7jDnpevnXdv0ZGmSuwhEZl6X+2oW3jwNPzEETgtwv+qW4lh/ZK9vGOrEou4e01vc7X813N7H9GaH
4bA5oL0m/LnQ0tqbceea6f7y7+M5NE8sATT+kBZdK4EW8meURYIuOsYVumgl2aBy2Pj208r9aMsM
xE17WC30OwOtW6ODas4TSkJvJz8zwTTEYwveDcv/ewvHuqLWHD3JLPwIOCSKZQrpzE/AYyalKK2K
u7WnR12PTfNKKoRupa9y47QvzKXUAC4xHGgZT//5qnQP5i75hdVIqbrBdCMHHe4QRZfGajZWIzJJ
2GGjkSBDa5HFr3OXAxOXVQvULvvEXLc/1ygjTUOO4Y1gQXxmkg9Qjna9g3iluINTGI70rWSjbUd5
p5BewlwgQ3zhklCP/f9jd//F6STnK/+hEt50dfygC5DNcaYjMiuRS8M8/lQ0gOgLPTOjha5d9G6F
bV+ikiDvoJjGLbXy6PLiL3x77w/8uLnrCshOaTRNPfzmBYQBGXmbjxJoXgbHKLZUToq1ZkuxUDyc
byRtf7YprUfIpfE0/+e/GAtkU3euh1no+j0pe2YxdoQnnSNShuFRLpbDwWvsPogv5SXT4FuadFVM
gEftziIozQSliSHgtfg/MQrQIFVhpMspgQ71IpIAR8TmXMWITW6SkRfy5t7zfcQYZMA3RBbKzJJ1
pKnHzapvsT0bHb5xY9MEY1IcUfr8ipc1rZ6oLIlMoy165v4FecS3X8oV96z7AN83ibt/VCk7+RfT
vkweB7po6a31b9N5GKk1h1C9Lp/Y+jdwkM+mFTrTigFtMO8Tt3+fm1wIERHxI4RSUQ6T0Jb60oi2
TrmVX68XiL83pboIkvF0xIa/G/2c2CWH0dBECviNo1qrmZgT1jgYtBqBTtF8sgNVy3cBtbcMljh6
WrBW31xBTzcDCQ/EHAvFMJ18ERFH5oWSVhcwbufrDunSPA73SUm8wpxk2ZjTLoj5sKA15clISWXP
FWaD3CpAdNIbwVKsQnWfqqOEQAcDnj9tgqyFXTRfQgdyGlB+Z/OMMsW4JXoUJpGP5wfLMdFCTVI2
YtMYT5qrRThlM6zx34E9iPtrxXUf8Kp99JxbshEruX0DKXAlpTsG/VFDV8J/bOegeyzkY/AC77nn
esJ2oBJK3PzSo/jNugHTBBH6nWdcnp5tIuj7E/UlEDqM1bM+XhXHjY1Ku5/Eu5uy5fq+lqz7JbI+
BatGuEknAH5ugEIzuQdrC5be5IY+8Fo+kMSJkHP5K9+oPkm/psJa+dij88hXZ+C21mAMFO2uDzQP
PyilvrVgbg3MOA4I445a2QiTIoQeW2Q7jIJw8GKcrtJOAONoleFvJeBrToaT8PLqgsI3os8vTXYL
/u4HdyqP6ds5upYaBqhol76YXvWJHYmN9Z2Zf5/Y+TDmbVl271eQcy/qDjgr2QHm5sZn1UJuoRjN
GI2YHYWrywVlHJiy9+LdvIKnIh+h6aXBR7pZ3k1sPT7/FIEVsm1rYZe0IyPxl/tFOeme5gwzhc2g
01pLpkNu0nkFuf+tJ0EsQjrcrsHiqaYb05sgtp+N22iJUnP+OOz+Niihvj5zcq2ORHMEFK3KT90r
X2NQokR9dPw7hvaU8mbMWQwHf2MbCllwTMq0wlZhMN+11fjioQvy6eztvl5A3p0RjIp/sKs8QqJO
2zBG0h8yTOdEGPrfVvHpCtRceTrr1WxvuG7msXgRpQ4KNF60rtGGTmdm5ueYhDp98Bl4cuNmcAU6
PN//lmcS5NYUyIH6Cym4mBq92/cBI+DKCO2GLrj6g7TrTu9sOA8wI9FxoY7nAfeSPKlGcrhi5+Dq
JiaZvRsVKSB2f/w3RZ23DJtZY+GcOHfSoB7f2hlD7zHgDyj7vCPrpslBznN4IJH3hlvef4C+tuLw
5i8XivmXj490gV5tr+YgC3/yX+KxekSsnuJeiLpMDI2V3ugv1uaB9dBgvSq3MjeN3vWbXUYyhCQU
UuzHngbZRNPqEFYmF4HpkTwIrg0XfEk8rUL2PqoFEYH9t1Mf5zgrrbkkh3UzTIjNfnQqrn1Xa22a
TxgjQYdRDzW+LuVsEldvqkOaEHHSMXsuFWl9Ui8adf8jBCnxdZhGomQ07jVeqO4P5anrW7kdczXd
09vx4CZTjvWjTkiy0WoB2GZRJN0FTP9trd5h0EK9+DcjsrLi/6ykLvR+TqCv3a4S7L34d2nHh9RR
K5OM3C7dQrduwgvBefgDQ3zACyH6TxkfxqVU0ijdpzEjFDLBNUo7SpUZFPdDJt+XHhzOA5yYbCF+
RhXo7wkI2GmEAJConSQmlPLpHNUwz+ICw+eM86WQDGbzRSghrdyiYTF3ed0O2jIzrHti8cWJ9u0l
NdRwiuQTySBi1pkEZFT2ya+eqdsX/UU+qouB0ePT5HcuXi0hlGjRJUSgK01Sxwq8V8q8CmpuyR+y
udfMjJeLLOzez4X5/oc5wOovyE7iHhCAi2aKojFHHUs85/YH17tiz4eLjXbtF9xzCpqwfsBUlJn7
Q8zYV54LkAdHuDLdH/jUDCgrMRBRGBSYkqssCha4+G+yBQw7Y84gBONTosJA3dE4MqbhT2SAmfW3
WOC08YBeJwf6YK1aunZDAoxppyhWKxnhsNdFM0a+6GT6XMuA3OB++GNo/+7PZqqmhMh+Y0dGHl3e
BKGnoMb0HqpMSjYmR7Z3wyTOn36kl6fQkovi2D36DoJ58kL0W4D+09MQ7wR2guqwfTacWXXI71b3
r3cImYAHJWVkfCrbrS4kNsdul3p5fhE1A68PQcTbm8jzrtM93FVDX8m6uN7vXgLsCh8HbKzr8GO0
TzDtEJj4u3lfrbM03VdDPo2unBOT6vQ9YE+eBskG0qE4pvyBgYW+EI4wYmteWYIyVkJ1ilf1nLPq
pzQ9oQ75L206h40meUUhQQZufwu5NWKZrkLv9UGDXFLE8g++PCoepxMyogteNelgKm8V8AbTq+qR
TQ1cYxuHl+/TsVFZtr6+kPiPAd/qWDtZaB3AmcWPmaabo3RLxTXVDsKbG+bOQId+PCHFisCl0jxP
RHznxGYxt8iBQa0kOewGJLDr1zmZU2lBifVmd1oCHAYu2mSyH+wuK9X4rZQ1OrSTxXFSKY1nYFej
YwW2hn2aoFT3amFX7gDSadS3hh1NeWFXxKtJ8p5lcp0+hUoExF2vgpRPF2CGL+Aur2WogBjPwmpG
BQpKXo3WGmLrDBNyzp1PYraqUA3pHYmr1zfZTwMK3R8PYXODKX6Fc3/tiYu5MvnubSWStgsa5elf
oNhsc5pYWSuCYCSsuIhjS82lN33+lPSM21EwHEiU7vk5bMlMsNJgh+n6kD+dhz7AY9K/vRP1U/GB
c/ggsJuY+NaJHOrfFBf5qFocn12tdSZvIoOoTuUJyNWdDUgccUbu2Jo0FqK1jf/lanoA3e9z7n5G
AXAJnYdEViSR1qU18r9CMgDYNTKcUzYA41aN+Hx/8i+gsodnJ14zYyxtKOCVsdqdirFEHPhvHh/C
RFiIgDVfwCYn+MIn0AnAmuK3nMLJcPIQvIP/PQgVj1s3Ad+lgslBLJ1DK9mOILLb5BPtsqiKbOKU
nn6ctCYSTqsSa9ijpdQQwNmMBSSu1IVHkzShOH/BK2scln+tx4v4wUBTet3Nn0EYDMZjX6H0h2Ly
YrLEcumqXmaerGJlnPrwxjNhShI3Y9CEZiYgwpHC7pi7rSJMnK9LCTfAszChFaEup4ca06RdoYYM
ODXJvci43Dplc0zuYYZMWJz6HmWsHu3jDut/Wn/JXnbA3JWBKQhDuWia+eLYL/18A2NvR9PUNlQy
e6WjgQdrhDx7gfT/p6tRgATQLwdUyj1ODJc0UW2EhtXo/eRmEZY7SdfFZEWrXudBWDShDCEkvGCj
D47c62CvRoW8knEBkz6Ps6a3PKUN8duIrTsyXPlX8mqQUAf1Rmiw5JGXoczOTxi2sHluzZtS6IcW
2ZmWBg4zlyKPV2rUT21r+eVG5m3ndTBXp52HIFSgP5/PMQOg8VbWVj8Uar+pPGUTd5LDvWIOeywm
C+1ZMkS/2xHsqxd15Pz7Jsjpb/+ysTixJA8sy+Aj1Kxsvz7LIC9OjtBVmOQQak5ts9i77iRbAG2l
RTaCy5ReDNvHR5v7TmBMOCfBgkZeTx0wGeO8/i8rWaJvEwo1GOfvf649IUJ6ZSj80ZOl0eEFXuN4
IAHwAuxRsli4sfUjF5RLrPP2yhUynENUtzyH3ffkg4+JyNcpoqlqRawmvTJvMRsLt23L9BlbplVs
RJGUzJJIAiYV6qHloO1o4/14eAaUi6oawYD7ZVVDk879IJpvM1Bi9FiBEnCw2j0c4k8Bc5omaGVz
1DNWwDdw4+q57WyfoaJ+5tcomRuQGUauMsGikPyHuZprA9051eTcjAHF5CbCfTYojH20GUj3uBbP
iuwsWDv0ztCpecdd80OM/WGB9+gjuKq106ffIh7fHs9cdLkTF4XaxJ2jreE6sulR1yg9Iu29t7B4
phJpwzEwMxlB51OlSWj6g0Dm8TSr7Jj6IsjrgExCm4xjd0Kv4hLzZEwF4xLp/+CGWajzU/ZZcWHL
lR8rFslpyLh4sXJBIs8ijcPI4MFfDDBD4MT0H/2SiiVa1Bm6fHKYUK4jkrjGg6tAkvMQMY0zxatJ
I5rlMrdQzv6nYn8SVGbxyE6M7vwDXddtTxBqxwl95Lyci7W1zt6cZjU1bjvcLM9ddbnxyDz6VN0V
0vmqt2YYs+VVcRHxfax+rhg2c/v6wADyqR81U0AYiPC4mT6Yq+mKFLW9/50y3ahnSEbR/OpUmRUz
mzYuUbpot8EkCp1F+l2NdTxuenJmdzJTvF/XFVfEWY/tUCuHjQzEufYg/EQMLkdHvNvB2Tjw17YF
cfSK8NuZ1UdRm53wobflKO44T6fM12iEMeRc7AA9InPi70eWmG++QS6pFcC3DUV+o4/EX9br6s7X
NbKY74ugjrp8o1KkUPbfWFmYpgmI6ZUQghXEYtBHAYJshocAMylQz1YUqp98bf2luD2QWIyzGadu
XKbm6wvOURyYPlmYWC5trbrDBPdWKnpVdQfYM0NRNhyL+82qF57skRV/IhIfXjRhnWBBB8idJvvq
AnTlhmfeSTjS6vIcBFeAXXLtTFeSDCDIXbgNNQohZPIkNzrSlqAL8shRdGshAGwmrsrUsN5I5HoS
rGEmlW9JjPryjye93NZUUhDn7YVJn1UEV2xRJ1G3c35Zmmxg5Iy/LsCCtgvNgkYz4KAXLuJGAaOG
lk1OilfRb4ADQ3FFxyLf6tjy8UQOCxCx6zZrQLMtCXsHY7JH7WDi2f3PJn2u55QNAc6ns/Ym/TVc
0SZtZ1ZBGnMJh9xMq6T79qMxEvQNRU/YiEPPJecaPVTxYQu5glJMay8EhDkbLByaiHnUfd2Fjpco
zIuX1s0Gm5iNmqvuI8ipes9VaV9wZsS/PvXoGdWKburG5MsuaEaKukBZbLzFA5qqSHQdt3M1TV0g
eEr6+hoIefpv6sD5u18ysRGYW21libN2R1W/usMw9nvC8eO4zKNqqc3VAmK806Y2FAlr72Wx/kxh
ns/rbEj4waJxuFZyVKPiPbUCfYrnOczQ9K4nCQykyD6hvy+sO76b0d9P5l9E91AjOMxk87uXdsqM
MHUjCaK+Jaras2Qiy+r15WfnNql9d7lw5Nv56otKiP1yiKG/AwiQKlfWtCEr4x2xLuyvf80N/jmN
WO9lzueGI5NnFLAUgnVREph5ePi1YIxff6DmYaBdSldoqbOMgEIEQS/rq/eMyRJzyL4c2RtzyyoH
gatKpm3yFVTXsEztvl5kZ4P0ZUkpT8WAVcOdz8qmT7UTK1Z+VbbfMjMIkIA1SpXfAwmBtz4acpl4
rnLlLp7Y/9P+thR2HGEaEARwsVy/SQM8o4n4XS7qWHfBXMTo6esyGWvPlWgLfzaY3M2erI2hyGGR
8aFd4SbxSO1E1z+nwrFkKcMbVU3Xjo2FSdTsgfGu5g8AX3osDbj+/BFeSGsBEkKiW6FoxQm6vPTA
6Nv1COZgKmsbZxt9EHW6JV9ft1dqrX72IW/UEgP6cOLt4vMZOGwu3cXLe5PqI6HinzTW22ikD2tp
/+n5Vgrhyh93yCBpfStm5fECXMb8eVu2VC1X2AtRI62ubb4N1QPB+twBGNZ8aO4IPovzTnDuY3v7
0/zXah47Iog2a0T/T7Hew4d5M3V7xNtgonVgO1g0TYhSvh4vCAdUcL8kw+ZW+21WgSaFwzjZDC6H
Oxt4cqr85cO3LiBExTRCaxryrEkFKEuvb+bJFh417T/ZfIyQKkH4urkPIhk1H52jWM2EHSEpGw3H
M+jFZs453tFPuvRaLBaoRoUzW81o6/xwdnG+qAG2vgiOMweZApT+M9Zusk6AdVFfnaaciABme5Sq
COTREdHKTYno6foEl6ZKiEJgSOrzvqDhowYjYi5uyT7tE8bklk8cMm+uKPVrN+LFy9FNeGnV8YSt
9YI8X7ejYAYvkclF61ayRPQRkHJaixJGun3DOY6tlJkapRKXLo2iKkUxgOtDS94xhpt08EDPF8sz
GjT5jZTTUMFfdfgfCE/dUFGVC3uvbN6BBSy2bRhYB0INSVP6orWXXK8G9aV3xT8oVeR4LR4+bOV1
RryLy/1rDO2sfxBS+hH4BnEk9D49yvVLeE/1zUgqbRYUqKt4il8ubRb5kokD3+f/4saAVsSQ15fv
NkVMaCHk69f+8sLaJ6v/Y58rQT5SKK/iInB2MSzI2F/vhpN5rS+aMdT6RDyG0JlXwo0/G0Y8fCHZ
GQLb/s4pN/R2MkHzYLNrBKgL54ZMkU04Gfa2S7h4Yspdtxlmms7p+CoI1kwFeVEqFwXwXbdotqDK
344S7NDVtH95taHgoBV9TZCVccVMvTJU6iXpIS1Gncj/nHHrwvROdIrwK3dfUH/0+dInL+qX3H9j
nOMbDxvj6Qy+09CN63mwUQF3Cf0ef5lRX42zE4RrcJFB9LR9KBUmS+pDHddnyTyqTNyh21G9lhHG
EJS8fywogJu4HTpsG6iQFPCgQoNijN2DftAN1EriPwypEFk+BcWDzUF/XCxqzwcUK8rnIjs1OGPa
zhg//kg48xfDPmrNpISV/yKDZ8mSJtonxF3dBylWpdCPXW14SayXjSptgWE59rFvTZlGsXskDYcY
6bgYAo2Rs+QITX3Eq5y7NXdyhiU6TDAsiwvLDqMMcReNnOpgJzUh+es/hMvgUT/eb6qtOHY6QL3y
r+eMmZgePnSuFx+dtPqcD6OpRL7R3ciTdarN1p9g7YpvVEcNgCLgXMzGOV8WsKq3hOQlhCxAmWI3
573oWu2pz48iK5VKFbbUVaWAQolW0YIx1HmYpOojlMozQV7f9QAzBK2k5bG5Nd2AJXHSxWvj6GGQ
+KVEX8VjxqWSTD/5ngSHyHTJw3sKBQPtd0fjaGetZ33xg4Hz6iWHSB2wDUUQXtrG5yEcNcnSc3um
ijcLErg1v1MHxMF/GmNPiv5ZhNuMV4GvlexpLdtTOHTGQeKPIAU3oGSPMaPFM7/+pu2yi6VwItod
XSkVDSn6RhO1+0vMzrl2pgfbQ6smc/SapIKsoKupzUNxM7XGHIhMLVK8FSAWpq8yrAgYLYHAkOVv
PYlGv5d46cir8s/Tl/wnHgFFQd5vjoHcZBJc5J0K9u3YKhqapn7NzOIrVVQiCrdnn676MBt/VHxW
C+R+rtUQ9lYXJTumDHMDa4WveqQIsetmBL0Nq97bPLqcHvLumX7LNV+CRapnh3juGXAk0L4w7YBM
q+Tv6qTA4Y8ECziQB0Z6r4+8WZNZ+E4noKXKyvYz80YHVLlb/x6FkGxiR1VQm0M2x9bBTzNsYctB
N5R+j0EHzC4DPiYct2ihkJ/DoHKx+gRUghjUyEV3aqd9DwMA4lcr2H4+8bHvKdw2Q4ormJgLG3Om
Re1q3YtfJPgYRU/oXnTSspLRan7+aIin84GH97qrIaiMWI0NCf9voMAb6NA3+oxQkl9qL2yDGuKR
CDqN/SLyNiPhTgMU84WFN89FZOgKgFzM5Hoi4BQ/v7ZWslqLjo1H9HOcS/lqI9WcIoWjEjz2/AV4
nj5q9EyxOOMRta5UzDBr4PxHnR9qrd9RAcOYldlujx2BY9z3nZTwPzdFgV8PWd5YGB+AIiyov2PZ
/SUECuXhVN9eUAmjgKN+JwTpnYawWVAL2aj3t06fTPdr8a0EQqRJ1jUy4kJbckxGAAwp6EXwon1W
CUvAYN2WV9NR3KWuuOJje5zPr5TfazwyuFBYt0Ta7Yp4LHFKzSS5ihnO37PCebyB0gogi1Dqre9g
PvXLHj4zongSh9exoqeg7oeO3IPdSdUDBHSP1prdgJAyzPcUagb6dZAu75n+/qx/ul9TQf22DC0V
WR2CPQiTiT0djWMPgVE/p2fq0QnCE0eO7dJLHVk8XHyNWIzJuf1CB7HbhpCrFjWjL5XpdPmz+xvQ
pM2rfPcEXhwQXAc6erLzpGmqPqB+/RUYaIxhRzsauWO2NJ0gUIO+4mKvaktTDbct36x1vI2HJXSJ
tJtpPWL1ZqMx6VNL2bcfTrPme8TBEiGXr2lE1thWwpi3VqurPuaoAJ1j4qJegKPJWV9kVq4oMF5g
sX/cxwWFy8j8VzXEeTNxv3yDYo7FqzGwBAHuVGsTCQ5Cui5aoKJM4eP0MsXPyCPKp2H+ZBrccTfi
B3AAB2UEqdIC5m+0WsRqeNMuAGD6Hh8HEzXC9261eJQb3l9x2Gvn8yy7s2bnCucaD2bOkKbUwdi6
47wlqC1AbEsjEMSq4TPdDTfncxjfHnG+2blmQxoBMiIK5Ab94YSNhTensWAI+1q48iK+Z+qk29KV
YGkabgOv2/B5d2crww/31hyMk3ZdGNp1JcTgBcrskxP1wZ8+Ms/mh+tCf0zRf3LFjUQGR3BvrgKY
DeoQwyjsquFsnN+WsHF0cX4MRaev+o9K+oPTCBilrjqtqYNG3jwxca/8j4VvGzWCZLrnOy0FuWr9
9VWPXeGEjSx5FvSnCKeZUY30ianx/8X5rem3tzNmL/zaG1NH683YXrdh7gw0rfXjxfA1mmaDjrcv
e4C32Gq6ixz6FmBycOMJY/x4AxSp1V/mqkC78GJiVIQPP9l25YRE3KqgQKIht5qhOf7Momg9rNVT
ZU/B+a9ngTOBj0SWrXQs4ljxY9IBJpL5QdChaip6SmTbLNO2MmC1+e1sgYBM2HEZuY5AgToK7TkN
YCqnLPnSFx/Awe+LATgc+uNmEb18Z/gKsTm5xHz3FSD3xn2JEF/XJ0a8y4SwzSN/ywqmip/BHuXb
e7vw8C7sUgcJn0y53QQnFM/HDyFBEhhOQushjp+Mi7pGPTwAy4wsRTg4+cgyHRA7BAwyyPytDAsp
lRy/oQDZkG/6rtmb13oFwF+x/lmWaoG1fjS4Q9Cbs8i2B48zmUSBhLgQz3CsloE5TNRIP8yz5Olf
1iC115YNTGW58mipkkMHSNHpoh+tYOTb31f9ogEVn1XyQx5aZfjlZcTY1yjeXns/SusoshqvcUMh
Q4Hbls8JRa1+teJJiwBzDmeFp/mKTqZkOAiVWN6PC/Qp4n9J15BcLheSKD1JELckLc5KEMQFNvHH
9nqjcUQLmDy7H4g2/tqSl1VlE7Tt4SPGl/oghrQk4jjHQxpABwg5+q+ophMamdY2zHK4cImhMjoC
gB4uexAcImtO9AWE6P8/6ZUbSsaBghVxwmZi3IecNaISYsAhVldzp4wWpkz77A4+25rb9y+ojEbj
Z8T+WcY6oBMqMCLNiGB+LuPBzew/MDd2Qs0+8KwTMB9bsfgXtaMw3IbxUQQlxFliCShgD0k6cLFZ
ofl27GmkclJRQD4ae2pEVn/5h60l0GFIflN7+SMyWMkLslyVCNOMkBJ+mldzBZdmOy4Z7i7U/knU
dF1i9o7opQUI4J0yPqaXA3yiwzWuPtDW2LiqU1Gfovs0aLpOj7bNAsVXQaIvfieB15/UwyEFDMHr
Ou780x/iYBlP5XQKdJzDvJ2TITa4u14pf35Gef4jPtFIup8AUyMc0akVjN1W7EScpuuYEzhYsM+w
YPCg+K33CH7cSf3KdDl/6Heh+rrfi865CvrMjEio+9NlR+1+plfNO0RQnfaBDKwTIPn45+Nqt71x
94rSi7GKraUJjt2pgMJw3q3slDrNYZmnnLQwGdDHsa0eHRy025eyF/+nuBz+HemT29df11/mcMl6
ofOaXTzNOocROPUM8EaQm36jeajIMVEc/dINk20PGXYFon6vpLXExbDefwZy4aselKNbK4eD1UhH
q8bMpLU6C23pUA4yPA6oU+gR9HZfIi+Y1g1z2eDzvf6mwBoKu+dU2ualK42cT0C4DEG0I9Yuvdd6
0k091VnKDX/MXrCleQDS0ruVbV/P4J+ngA0O9ql4+KjOr4LwNXevg6mOP/WHWXWiPyOebdq3u7u5
9I1OlX6lyzskQFhMThj/XMCnqWF9qhSmdOHTOqEQpOo0mP3qLnMNdUzT93/OqElZ4R3L9RcfQDgA
u1wqPnZRU4NpcMtYN+XpgMWe8wcYWF/uAjJzfVx/TwqauxxpMNrw8AN3fTTdgGG5ERE0fiNugBiI
6gZgga+49raPf84c8bgpoLzPD3mbJ2Dd2KhirFxbwk0cs4GRyjd9AT/WWw/r1bGBWxvo9TG1H4ug
A92EiquhongIzBg7/6Kl4k+oQN+XcWJKrNKsKz5Lqjdk2MwVlsq4wHAFWzkGXPY0Dg6mxMN2Hnth
LWhaf+28wveo/yDZYj0OktYoDl84qSuSUMdMAYC8zp4wbjhzRWFWpb2tLXhuZ+79dxV1U3KSkP+5
vibwb9RID9q2yiBELF8kvigsVqt/53jaahqie7IXAjQxpxJdYYCmDHDeow+u5TOlQpV+zMx7/7F0
2wrTCb8bZCgAVCwdVyFXyHFP+xUGkx1uUJM/UL6OJTgRwbIBVyAX0cc1lv1mbouLxn9e2nvQLyP1
3u6yj47XCKRRKGJsjC0YGuPHp39GNEk7ao2NRi3nRn7coT04ScaMg7po8OvRfB6jt3i8FYcaidWB
N4zeC5x5BMpwAuvEf2YRiSe9/DsLPjZsTVh7LDGofvKzNBJOYxDV/2gdMMxE14FlKCNU9VJoorgj
/pIHAId/Nhkr1AgQdN4TzZig6s1VGuPVOxQK5/BsrIziwC12zPcDc94sCOpq7CuzRA4Ixp4wIr8o
pS7gXBPRkOjmo/Hxq/2YfE0j2bsnaFAD5p+cykVO/F4EBL2gnwfAdoH2Bc1B/grSZGlbNl7r3WkO
1foIyFArwjEs7cPcDrofjG7if+fO0RdIiHAtKba+7kFtiPDYV4UUZ/+fCOcW11ilkY6hlCsafkdZ
Dk8XZnC1GhRfgZKiHTHhuuF1JCDa6TU9TlijRbhdjDcCi+Su/WFIG4RJViM0YqWxM8dBD0nzjnHW
wUq6k8fyae77pq4EwdmFYBYu9IzYvM+t6ljwEqI+Ob1SaJZ4zfz89BggaV5KXJLB88c+oJuIS/5e
BH/m2a/eINI3GIibFc11E5XuqLmWB/+plT8yLNuBKDIQ3HvVcDpnPzq7MBUpscZEapD9PaJFerir
E1ewAoCz+PFvpmBSqbj8RIpnyJDe5mj276pxdLLX//Fe49oLAn29hL41yXRXVNjLw6z6i/JlWl8r
G1q8dvse4OMfEyZq+qmZWjHs/GhV9FyPk3Up0UHzVpt6c0fOQe4m8JMILLA0IJRFHcno0qA4fUR1
xcaffUwCwdqJmZYLcnZVOvLp2Q1BcmRp3Pt4MBPKoYjmv0SFE4WvlC7nqPT/EtXduqWCnas4KDhF
fjjAJQ4UvA1wc8FL9/YnT9LHj8EEciIj70XfwQQUuN5aXciDlB/oyYsH4Jf9bfHs+1Nhmu5t4uf2
cBNlyVH9njn/ySxA67/Oo8vUURr7qvQnuyDN9jIdTMLxTI1lGxvk7FX5qDq1LIjnFwDy9ZQ5JJQC
MgHOFDOsmohUAWZPHVyDdUjQOb5arnSQFEjoZaTeNUZUTy+BS1P/wY+dvyxh4lzQTxJU9cCpRptk
Rl7ImnKuhLg8fXaYaRbX8gkVMYcCccW7euxdySxHOdrtMPYhSvktBFL1Pqfwd6rQh6XlD6h1DtLf
Z2ojYmOBwUgQ+8Gp6Xq80iNVy65wylrlUX4bnI4aK+9tRu22Jq72xKJByGG91WKIaU1+F5oCpmMt
BX9DHx99FSNOQ5fFJpPbc23SZAvpGROq5+zfOO1RAM3YZ2NSiV3j3e2E3z7cBKanCrFYBY65LMeB
j9aKze+NCPu2htO8W+DGahalh+KcP2njV8k3lB6nsbgn0f2tcM6JbV+Y2mnY//PJu6ceV05LSAl1
NwzT/lyyIsLS6toL82Q/W7gwD++O1mXZiPGsPgSEpslWhOBNMZrBhPcPMlgYvkLqLOMnZ+V/g7uj
QkGvIzZEHukrOg8I8NZa/WY5MF0ywS6morjkyHSs9Yc5BTaO4biSIsN4vuCM9SnflEtW8s6oZkLc
ZOqjdHii8saAFkV+1OHQIMVp2mBC8fqN6U745KVmx17wzatX1fVjPbIENaACfQhU1W62g7i7TYtO
lYM9HpcxNOCBYPAFHBhrCWlj8BK8ULfk63hhKm7o9rH3P7YRWwe7EdLbDZqvyeGRH2IZE06Shrao
07EBqw+LCDcH2CJN1ejKH2Ji6UzLUo4Kv7lfEBTJ4WZgUzpW2sCoyyXEfSaCBjx+yvnwkmC4WxEG
VYa02xd7PWqnP+BPsyxRtQy9avysPuPkfmRSItkxtefeGY0k5tvD+gDmkr0wB2N6zA6JEI1ljz2+
cbExDwBHhHgrItmvKMDATnhWLJrIamnHp+JUisA0KTSfIU+eXDkvU5JzpooBlKQC1PtDn9gtWfbl
eVIc9HPN1r5f8a+kYW+74lHrJNEpP/peaKfUh6oHHPNqWu460qCaJa5g+6JtfWcuxJrRpa2W97AD
EFGzt9NiKmRoPlWfIfrf+djwYQKU0A/IilddT32tYEggp3r2SqA2qE8QRUNZaW/HN5rIBKT9gWj1
KAD2z4CrK7PSItWnvkY4I7PtjKOF3saHzusxqTma7U69rAxkGRTlhmkH6LRjC6VfkulwcPvSSFoH
8gOsjiC5fI7JAebj9bc5jIeiRAIHhVP5GQl1tDKGmulNiu2WHZaVqXrnLy27G+XP7ICT/7eLOWXj
H5t8myneQCH+oXwHkhU+I/w3rCjdq5vepAoJ4u19I3S3GUGhxA53egK8tWG7OqIvo/VggJFpeUOh
F4IP0B+jamBLaafoLyX3iLixBO+qHkhiNKW/e595EVi7xQOobzUY3eC5CR3z8oKbE2PCTy3YoPtm
JyY4dv3dREmz6dzrVGP8FEEX5pTtXC2oXslT2j3durG7OkDDeQ4CiY1pPTCcuv2N6vrfldjIH2uK
soN/ADd231GUwFlMJuaJeGNTcHLedDyG9Fwj/bdy+hxK7zHKydJdnyterlFlEPFt8HWmz7b7Xvee
vpbr1irU70IB1GTuZ0rFaNf8WHmYVpDjZ9HFIi9HoOJaiiP3V0jCV40yT7gpGa5tkdC1mo3c2sCc
MS6V29tife1D6QTk6lx3j4PCEnoh81IElFelPgO08uiW0oktzZfW4TEV6H1M+AH8AfEIbonl6Ivl
eyCH41D6i+1ZILxKMMsdF206T39JqKcH0T4xwaHINUlBO8GCG+UyV33fTuZYJ4x5eHg5lInHOPLx
o13RBo1OPIWD7093lSCBQWwSWnwJNBdCfvJH4mVABka4zZfGmXRYko/ugSsdml5FwnnL6dt/YBbQ
XuzHp8d3ObcBJ2SGNAV0e8fGZn8uMXOiWWV4G/x9Uj3zzIHwQuYRGteCrIRdfuT3VTU8sZgrWdzw
H7LqY76Kg4YIw/YC5EthyMHnkY768Q0KcFXv33BsykJqyyX+42/Nf96VaFc8Rc5AvlJdUEE18kML
qHyR8FEZ/vZgpuHwIYO/8jpsJGo6lNAKO1xRNLLM/J8TIa9tKzohLNzdSrlXiwJHUnIWkFck0VaQ
PmNYfxMklFjVRP6pdqP2FN4hsKOCs9rEA2qsPefawW0iyDs+p/vqHeOewHEjpjU3Be+sgYpwqcxi
MF1HcpXVPFOgUl9HZt//DOcbHEOwURP4ge6GK0S+4nBQOejZT3N3QhxVx5NDo/DyscoGeB7YAt4i
kr1ADx0RaOHFuhIYVh1/8TYiTPN9WHYyi6pJGIrFndFVsja0VL1WBb2EOe6B79rmPu7DzkZUH1S5
A6ZnqWqHW2T+5Dm55YZ4RydRuC2OvI3pOZK9ACFN+OGkqZu+a0lgZnpdoxSJeauYOwiYD41EZApd
9ZcZIHJNrgNG6sl+dKh+hguOAXPAM1WUwYe+06yNkxBonXTNpd45dN9VcszUygYzdMLGh/oLcKrj
1MxQtS84rW4IYu36QFqvhXaihxyPJa2ueyjcrVkT8eOD+5YraxQGGROXpRj/EhD+JQTuRh5EMtYY
yvPxRlzRyzutvT/NT9RgR0MPkb4hU8qKP/mPojP1oGx24yDrSbN35L8s/8bGV+p0V8rJ97jOuagd
qylr0IEsqIryXVKym76t4rRdQKxTZAPDBoFD1IJfRXSgOsZODHeepJiS8lRwUjz02XiE8yfXcgg6
kx9TKMFNsQcPDGuuMZjwyG64kLy/eXABNgbWAAKtCziVzk6lGtJwpZ5r8ljNUJSmGoJVc3pOAvUI
w6KlAvMPL+bQgyH9mif/CN9/wDhQlHd/rQO8Etszt2VfzuKHA8AoPrj/qSPOfA4vThGHlPHlIzOR
NtDgUfHfDVbjsHfmfAVUOFcWDVw0bkOcRah+zd2WnRbdtdXdo1cxluZp2Ow1ohMn/L28YNoVc+ez
SP5husPGNzlu7RM3XtnZoyuj/pSYkSqs4xnTSaZx7VyGA+5lRGG1bv7wNEc+5naVAsVkxqsR1oe4
aEEC7FOYCLRHiLXT6bRo6NYWJitCyKPW7lwy0Z0JwzAVp/yjpAEw0v5azYvb6DdTXxC/kMOrUMq7
U4z6lWlSfI1Jo2Jr0x45CPk4KqwYMJFoCWIF9hUB9xyyoWEIs8hw3J7YuB5kzC+Y+KYe9JpuwWrf
0cBSZqN3BmHZHT867yuu5UkUXK4iVGHJlXzJ12Qrf6fk5NVrfaOZ7aP9uGPkz/jxRqjlrC4GYn5D
7U2/P4Rr0wxqtEh4rYtfSewHDmuARnlCqs8tqaPoZ/acopcTwIENh07TNpoH/o43mtFzhSGkURTe
aZrf/o7bFAoYcZnsJJyEPc0uCVg2Mn39xW+2I34DrhNmvSC3tJxYVJDGPeXDvAzP4IzchcLmzWSt
JlJQH7Qxr9VpRri8E+uECPWcqgW3CMLul/eBMR9Tzn9LJKyZbdnfeMfYFkL2pNzyCTCfmFUnx+ck
VP5qbh7HOWiN+qQFs3dy/MSBqgDCzaqxAP65hr3tIpC+X5f6lSqyA3c5Ppdnl7jqsmUx6LDFIOA1
ermmkeT46DSKP8pPNgaD2m9KOngVhq8LAWwEhj/cZNhz8bV4YD05aB37ZUG6JBOBa2LgoirimuyE
6G8/NLSaoU5Pwk8hxDy0SMLnJa1QwEyfyO15QC+HXYq0lQm7fHf7c2xbW9DVoj47369VFHJMWO1W
Yc80mt8xF4Tn8V1srIPjx5r61YbXnRhAeKsKaE7BxYmoX1eSGWW9MpurA4tlWp4jmCDAaF/mXuPO
uNFB0o/EtErc77t2w5Ty5M6vx7N19p3q/ngMcrkjNNo61WMR8Uqeg9uOmRvxSc+oWgLNoHXAZFTq
dUUQ4G41d0dZlwPzuxM5P5HlU8cRuyNnNk6Pb3JY9Oo75u+z9LF4JuCkUiE6JkpM1H08zil9DOcp
sZ1l44wSKPsGNDrEfxGbYz7sVqzgyzY58ljX+SZBYwpJcxTrqaLZabzZITqg65f/33H6zAaQEn2k
UQHOuK3AL1j6AanCp6dvu0odHkhAQgUum9AzCt2I4ByloQ6ktgmU/HrUL1jySsQYdWb0nYdNCykl
7fh9KyJpRtDfAPJYh4vedWL7ogRdLY0d1HTH7GXVrNTLk7WOBlLmdmeTFwFUHT3DZzFMsBeo3J/q
f1llfqR9UbWtM5t0FOptUbiCat7HRlw0L3mHtW+SK6d9zQs7zE91BdCAXsp6+zpELJg/SSbo73hS
3nSA59gcNZ1UGNQgd7Ese4ufKb+TTJP709RMU+P5RFIedHjxjeIIMX8oNxGY9RRlAsp7T3WR1b6Z
F3HxucfB+AoE7VS/48HadE9SwxB1obUryQOmtZTpbT1Ar1fdQvMQ4UyVZRlrz2EGmMJ8ZaCkSLXv
lFlnxgyBng7Am7lzSAwZoG8hFppD3NJg52rhnMj9vwkToQlcLo+PtVGFSXI1HIq23suqtPFdqdxy
0EFjk8xyTQGAyuyORhCFTyXr9482/N7kWv/knQFERShPegR8OCkWzKRiVA+CxNlLUmF4Lr4q02N0
svG0ZJQnRhLdk/UUCYMK0KAOsai6wNDm+LBVhdtzS0CbcZe7X3n+S7x4fx0VdNNFJONS6lmzO41N
MjZQXrcig3TbqlC5KjmXZWLgrS28xxFVe4euLSWEw3x2VjjKiXJUZBMZRECYt9zXqk2qd6E03gQU
P+mV8liXy8CytA1O9JnnkE6dgT35jF1xAmLuxsO8nHBhKhByHn0KE9QQJoQzECgxUgYTX2DD6MDH
Q+K6avyr4J1CChlcd1QWtFKsj8+FPiL0BYnrJUrj7IrtGZO+TiWPFFuJ+yAmMf13xiT5gnnngb4F
f5Sb9km81MA4+ofC6ww4aTFGQ1Wh4E/S/Hvb6n3z8QpGxS68UAbB4jCwM1oIkuy3d5sMvRGbRzX2
yU1svQdP5+wDvPwTlGgjzco23sXMoP4VtC35OtU+5LUh+fzU+r1jIAICxkV2btwAIJFN/iYJhrTc
2AKqReLCLF6pKwCUQ566Dm34hlzItSCghAnAo2ZFkCNi5YLoLzTi/v9mvIAwOoAdAl6zinXYC6Dy
RO9+jElRKDUG/zqolvkY7QRkhF3YCuWHhhcjR2OJmUj6UTyo/DUkb+ovoiAMmCZGpViQsGKwsI9M
rFMU822LjcZ+CnioICa12TuFpdjpa/MdIMC15fufBDHREfpjn8pBEzC+5PCW3Nw04e6giKeYE2BW
Wrok3tgUkp+Kfw2liXWN6yS5KExaXQpRdCeTUuFk9/yFVvx7nbqpMZMKqLuaWZ3rFIaQQ0q/Sw2w
h3v9zK4H1f2JD6R1Ab8bEIjKKl8YX3jESgEYiSOZ1boEgS/+1kdoMocBp8e/SKyrs9GdPDSTLxsc
Jg0AmgfjF7r3dM6S/xg9cRm8RezbmFmMhxdFgSjnn+PSr5u91Ga9rx14im0BLkaPU4QtMrZzzQqr
/3rA9iONas+0wJzQXdPkz0RmQj8+mwv3KvXjWA/0ojeykv29B9Va7r2s6Eq5SO+u/bKk+EfkEC9C
uDCf/ZgnNnk9PVqhm+XJTgLJ9OS9AMVOdqnkv13Cro5K/hDSB+w2tklFKLAdJxE0Vm+9xz9GZPcg
AgSUiAvxlUq4FbejofzvHPhaX/utrSjsQw8VLiZOQ1DJ3Eru0JtFZF4VZCDroUvxRPw2ObO81Prg
Tl37wL+L++NAOUhhk3bHxjgd0mFdWlM2sTborMumMrz0d8auOnLaldoOGWEKfjuJQHrAYiK+Gxj2
qC0+OohgDEnaqRdahSc3E2nO+NzCVuqP4Uj26xQHGpd4CL922PLS1CmDb/3jxSuSzwYLt9yciFhw
WvHVYokusXSD3WzoSAWZLRLZ5dMb15IkkkrQM/0kX2POG/ewaE5HIoxOFx+ecbGJKc7qawcExtmL
v3e7iMajieCePJHif4WzgUj0AG+62rYFisqpLIzZInwuLV2vem3iJ3iLisLcxFaQvXFYc7an05uG
ujNyFCsDppe1bjqMwgglC0h4MfKiE7Z2S19JCWkiJQPd2FzNUt2dhRoDhB1po+uDppW15d6HKRG+
kbb3dxRNxIJgC/O6BByz20zHk20bqXDUh5Yev73ovoTlvJZ9TIzSYHluHRzwtzztVzDo7/5QMSj2
QuDhkFOdjhoKMPElpa1u4QXSxWHYEW2KSgHlGqew2G9QbAzKWj7CPUN/E5viowwWZXuS+hu1+wyW
wDFuBvbgLo3jYOWV2H8aYPvhPZmChoMdTvPeph2WGOTZC2+FgrlG2J5btT6xMMFkgIeiwWhPHsS+
Bvd4dIxaAwxOjs6VOtouB1uJwDhPDjhs5vlMyLD+0KMqiq2kTlYY4nQ/fOzzOpOK5lJ0JVj+RYzG
SA7p/6vMLav0N8K+eZ3X3rN6CDYMI1tlfOxsK+NXdDWg8uA2l54HuARdLJ2vB3kLGjdFeEeFmVYH
1EktVDTYjiF/mFYqVdQKi07jFxl6cFWPY0MxVGc5N6waXk2BEr+lmxdFmNp0e2WrHZbcatm1A83p
Y0yBh2jp7Bf7w2lItBpM9P5lS8VB7FAlrD51F6GbKwS6b4VeMA9ah6R9m0s/qV4FJhlQK3BuhxeQ
sn4mj2QcVZTjZ+d37nC8MVUdWJZVripvMyrLd/cjRmeLp2OosH7oYBboX0RBLwLVylETC1ukzppU
+2VfmgDt7Mo53zlVOio7zZ2/5iqttez1/KsbqJlvGRo8FKI8ANnv3uxNdPiZn4+WbKx+YS7Fz9Ot
Zu48jMCf8vqAn0WbLep0WTgBzVJ5ZjNBxhg/7REANYlabufz5G6t2XABdK94iyEBBUFToiQe6KZF
YkE+H1p18y1oh6AHbifuo+9XLlvg7V6bwJXDfOVv7zv/PcSj8wfIhAONHkygbrb6/Ofuc4O5lEnR
8lnkucJ76cq1A6+9dBjpn88skczu0uARswZeEskJhNNAAynHKNr7OuFz7QRSM7LwSvzm4qqY9sbz
/kBJBZX9JLiBkn5+4ImDjjDPfJxB8ve/itiAA04RfBtUwOAV5CM+X9o+vniZ3XUGuHi98KSMDujI
QriBs5Os4i3AZHTgy9wm7jZumiRhmxcJyM0/D/SwHrZeheQS7JKX3fIUP5VZE4/tCoGmGhS4nGqv
KAZbR67wNuLcp4ZQwGFBfsilzVQ8VRUMgNWUW0TvKCyO5kCdd2m0aKraIcR+Yf/oJYKdFwbHM36u
3CxnsS8MRMWFmMp8rtqvg2WPyw7chdj/59ncvRLFCHKBAHrIEwe5C6UTvb5940bH0IDj4B6NAArj
kWcRQS9KF7RK+5Vs09CWQU8eV5nTdmcYQqi8y6hrcXG25weThCHRX5blosal9aWzwV/THq9DegNQ
HEknwKy2XualjxegkhQJ/O6/+8AwyT1h/l2ViGwDN0RqDfxP+I0N99GMu7wR00gyl1AhOGc/kMM7
al8Fm0Ead3Ayes4h3mY+/FCK6zRMZ29aEpra3gb9+B4I/TxCiZ1UT8aWdtz0rth/b+emyZwYY91z
CIkIHoj//jJp5KFh1iGbX1Jnj6gq4YKiPEhOts4dSjmoNJZwqgGGFdeW3W9/d1HRB7xsVtKvhrzz
ueoqs4IR3mn/rWEUj6jAMXHQO6yqaRIPfef5Y9y+WtTm53mH4dE+Kw7YnZZUn7b33txPTq/5bDjD
I4pWh2iAGMOzmOYambyqE7doKLBulRW8/jHABzBlhn9XtXR01QBdXRvKejTQ/aA+g9cINljk4lMd
dyMJGkx3Ycnztb0StagYXaLRULw9ahx8hTEfebMaDHvG1pqxMrWHVFToZmmz676OQFk6AfrpYpOF
EaZ/857Ss//VPyuNnNUXXa7cYVXLcIdhet9/sDw53IX4DntfYFQocuFH/YRW5VpzYLC+JPIVcsTm
j9U/9SfDBzSGo+84YlPpDnLFAtUZHaZKiV6GA7it2vq6QzyGY7WN+uEKtb2VevrdeASjNOL6WMoc
H76UqQCHOqS711K3jyZ3hMFEJy8RWe1rAGv2A/8Ll5tJ0eATRNinc4P3nMVNFQOvCHP/9kuV4yrO
GUVaOMXci1czudqNJVgVwf5+eYPaFdIyU7rHRHOq/X21ZFzPrp3M7m7gUzGkuEmOlpCKL3nSoOW8
/qprzxFR/ArJfx67OOG9DmJJdWckcAK2XbMQxKvhsC+Kqv64iM3A6TLzk9zj573dcU6FRfQksmzv
l5fbdfg1Wj+Jt6jIPNAR6w+xkIQv3dxyvuKua1ZrvPrci8ZvHF0XseJmetdo0PBmI8HndkeoraF5
fP8eondFsJBBxpg2fMQKWMG0s6qG4L2v8JGf3qY+FEqxnq+1rGhrnjn37y/f32KCqhpqWeMbf/v1
9w/mw9iF7LihAsXLvvIQi0a7rZYykUSjfoR47kFDd1r4h7Z+169FpFd/cOLAlaXCn3svVUhGjbCZ
eQqVTT/aqyvh3oh0HFqd627fW2fQEfHYG7j+3kgUfoi3uhNk+Is32Rn3niGxpkqPHPlT72JqQXht
Bm0xb1E2Y5RKoWD6pmKYUTJvreldq9Pi7mkQ3CaZFu5ghb1z4nEP6lOhJjalUNJIrMoZR2ot5YC1
Zhq9cW213zaYo3zpz0ow4cJNzpsWuTMn2j9vaY1xsoMYiR5ElSgi7naNOUPnjIi3ZeowBbgVSveR
0llM1gGDqQpeQeN0QCyqhw6CFgk5ieEWunZk0ExUQfLoLgDdLJwh10ad/UC4mWuSI88tpAOIEPnq
6EsA76ct6vTiFKOEvmzRwciydE17fuIba74WFc8Fv08fRQOVfxd1TcAw+GDpLbj51vDMJTOXLTlX
xKOdfdCKGfFGWlg97yQq97cWl7tPuOl0VdrVbSYjqXPiNjByLcjycwGYqK9rmtgXXIjDUvY3Fx5y
Kgk0fYpN6A2/1x3YXAJ7KqQBtvnNZ6EeUmINyQBHPpISqS19EVAJFaNrGwA8MwH4sakKBA3uyB/S
wqNbIB9XJib2PhnXrsTpWfDzun7a7j1/F5U+ZqvaA/LSrdQSqbB9itJK07xwKHRDLo3DAZtTg05V
oHVsVmSVEpSJ7soZ4yVr6C+Cj/wono2Wg2FKBDf38gMCu6GnrOBNld8FrGrQTjMd7zEMXW0xzYO0
YgdOBnzoZdueGWMBUsm7kwjGXrzUHFslCkP8YxNIMcJcqXPQvPF8TsQFe+jyyvNRWhtlIgp6MQQa
b2UalYn/VWxcCChzWkeD/090D8cT9YcHEIeS86yiHcu3OagEpEyFJpYwrWs01JFmfwGOiXxapcBL
OHFcUx7d9DOmjqW1jPsnnDcxDZu4NnSJDbfqX90wBZgnsdu9Ih1MDvE6u9aWGtyfpBfG9IGyVAAJ
JLrCCNf5gof5NwUQvx4MBLKgrGHE6UeDb1DBOLWnH1ZD79Vjtnp19aI5fhccYSTQGVenpka5X1+g
5rVAbO3ExuzLLLqjNqDYmW+uFl7WMoaal6z4JjygEi0lxXo2xqhtL3QSkujQou6EnKWgTQCgSMND
PPinbSTj9QrGFM5O8E1RXqNhvwS8m17SJfJZ50fdaH1/mmDGYdSKCcIZFRd8agBzMuh1WlS5fzyL
7/4iPZp2JfOx7nD0KqTJcJ7nglAXv77XduXvdngN3KjhSuEFc71b5l7SvAtwNKLDI1uA3JdEQoaj
RvkLbTjxVTche64j7uv6I0KJf2NwVW5Dq2jogi2w4F5/ODqld65576Z8TC2q6xS+l9z30kx5/n9e
FcX7KUPq8OmBnlp7HJ7y7lxnFEt+iuscBwmGSOA+AaVtSVPVEW7USW3QQM1+9Exy+DFTy5IVGkTw
NMJSrx5WGsbaW1FljlakWpGRS3ThnT1+aGeWSfnpuU7hg8I3nsmeW0v6ppCnUXsPFlJKTz7uPn8T
wDiz9VQ/EeLJivzKIIxpF5jDXh0gc3x/vhwgNFY9hcs4tlL/5Hs0/QoQgEWZ8f9ZL4lp8Xn/XAlD
Z/txyTQ7vnxBkEnJc67BV9jGmQMQHSM+OQChERUCAbP2bYpRyn6QWqADnQsEoY/m+9EaUaGW4zdV
nu1yNQvHihXL8O2YURp2VYdZFNfVPlmV0/Py0qPNO9jeInQcwSyhd8FKElHRzsAcVYjgzQcTx+xe
frpqtk3SVrSNMXdp8kySekOfJkVOUsSsqGZO0VnnbRmwjXbeAYP6r1ja0W2wbx9ycfE6av2wgQEj
d8oyGEKnDaPEqQdgbKQ5RiPAcdovsBPrZE+g/6EdotMe0iYcdCS+uPgRyvOjX3Z3CG84IBM9+GKS
AjtfxzLNdeTSLXMDdK0/UhkTwXTpDY3AYM/qTTW+BXCwjioQ1H9VPoxIaNr0xwPcG+6q+M3jFbxO
mz5khr83ed+EkXywkMo2R9x/omkh1Sgj9bUP9fEFZHVKMdyLCXWvm6eItTiY7wQhNi9CTtOqWn15
QD+h61QUFRwWhAuiMLLsMUnQUqS/d7qvWqv2r+SFgD1iRZAXMfEoH9pIq7TLLDzmi213BOMkbEK/
wGfiY7xyfANRBQ7KtBEcJwWomHkl0x2FZDMgWXQ8BK3/iq4ZvmqIJOiPIm5YEDqK0gfIhU62Mx3S
oAIylKDRzAG/ZYrp7/ze1ZgESWDey5fRsr81g4XX0TIThBZ7g77XAXXjdAktY1TTemUllAB6rcnC
dm8Ye4C4Kb6XrZXaVDGR8Z1I3ZX7QrlKAbfxH7b1xPemlvKVtHO1AtaOWwVeJkIDwMKADmcsJCU3
1Nhh7agUWb/KyBE9LqAEE8Ffp0peswwSCFiPI9xwmMLiIExBIWGnmTDiApIVyt1qLaQPPoz8/++K
xK/tlACpD+HCZWzD6LC90JNlhKJUA2KpTU7G2/W604VY5XtTHusT3OJbAzTA74QBI0Hki6TMS5wD
+2bVL+5M8DvvB9wMUJwVOcFIUjRv3tzQ8Wk1ukAk69XHnC4ogszJWxg4ATpSnhRIzZmPq7nj5DO3
EhIfScAdeGuMtZD16eFRQn+N1yH5ZmOdwP8+QcB2vw3B/t6qPDfRiM5lfsYtxdzGiCrnIpU8s6m2
TCppKMCqdfiQKjUrE82Wl3x5LTM3c5jK7WTpoUovLezLPdW4vTCLv/5UZ+g7jqKpdB5VOqM6mdfQ
EE5hTBjblgQi1sl4btnbwJJE0JUAvEnhfzE4Pfi7W5vsEAZb33iKnW/iRwRP4jB9Bv4tEKih9YJN
lSMjctteOSFfZdZTy5Gia//E9/EGT87Mo7Dm7gbVFaNELPwScgtCaSwR1YeCYpWg8nUTMdD4Z6ul
Fz4btNUnd6XgcGZ0b1ctGJRtj2o4A5Q1jp73VCivezcPqoVTMHZry2uzNyI8Gqc+BhyCxqerNB/V
feJjxqGgps7T3alhRGFF517NzRiXxI8kwloMT+Eq2fivlRV41tCRF64XVwViB0VS57dCRaHQU/mn
/Y7QtW9ZdE1F1MUycUSatYsw5tQdseCVP21xnnacqlQP372ug/M3Nx1oG8mn1iIzL3JWoECJUa4g
fNkbano3clZtDb+9nJLSd96XyoTOf29mIf9vG6QvS9YsnWokkolReCKqerCgBYp8WLQvMzFIVoxr
N8kSzdqPDbYS8DNv9YTxbhHzU/Q4zbH6b7ssUgJRwA6qYFSPH4+/vjVlA0Am3iZZIfC2Z2zhSwnB
rKrWiKCaBzYc1d+AQBHTQQQggqdmO38mEdpGILB+GZeXh5Xhip219yLkKcwiWffYRROmTankSHfd
9qovXpTQC+ACVZv2K7aIZJF+sjIoc8xMFeR1Stxp6Ngl65vNbtYoYIpVPtenU0RzjyZa+HeYtgQm
F+sP19O/Ufi8OhrW3gJvP6Ay5eKTfQY+c8CicV3vbdIhbrPdDXl8P4xXT/OXaiJ913KnTlYZlohZ
hE5hiIVD31Zs6bT0Zu2OYWDykv6eIfkJTy0rMMMzaJsqABba9yBJiLp5SfI8PfKGHZ0MCkkoT25q
r93F5iL3WEkgc0g7geJUJN21DOdeZh/qnaPmW0POYY1pOjDLk1/+bIc5b9vitT+Mx0U8UfdKbqWp
d1MqFTv2cAk6EQOpq1ooWJi3ZZaqwxRwve24d6RUhP3hRgGCgY1X8S1nGQMqoGVF0El04LqDdqjk
2z9026/Cr25PmvDZ0ofUq8ZS2sd63pK2RozZYnYbzUs9RdDDtGD/tE2gKU5dUDJ+bwo8mbgA3BgO
Kk3bIe5ixGmgYpBrYJTKjVtAgoG+9zl0CPwXAk6Elre+8mP+wQgLZsiir1nWjX4MhZpiwnf1UXgv
S4mDGl1skhgEEfMUNXoLVqpcoBJQo6k9PTlkh9GLgnwl7GdA1LJcaIvi0qUnK8TViEpE3887Qg/u
UpKgnaDCtRARu44+Y4nz1XqsrzPlDm+y/BoNdBGEsF5+0J49CViYIMfSa2m/oHg1FF+9o1hWSugl
IChEZmOFOxhLoC7caZp03cXv98KGDRVVMfLLXt+EPKHqL3P1GJy+rpVmoAS0sI0cugQZu3aze505
3Sn+9cf93Q0amYL+PkmZCshcJfEHJ47mBI3VnA5+21+Sz35p7/OPGMND3wiUZLqnlozYzWc1nkoS
5DnW4EsoJg7jin4YqpryReMEEkV3Pmpuzlk99wFqWfWBJDsg0iiDhwsHPluvkdluvn9JuAQPqkwx
WbOy0pu6OtJbOPOWVWXPRz/7BID4J4bJNNMRqdI2/9iyMmNrrC2+Ai7kdLcdU7sgDkEvQetiNyP7
oCapgBzNSE1ySFSccxk3sErLwI6iLWSaA6QkHjcFJLqrmYO/3IPIyRwsID4F06d2titlOdeRY0dj
LnuDNa441K7HLGC7Gi7qPuZCCidjuiiBqJLW+Dv4/rpDsh1cTDq9uuWM72w2UmxLwcu7SXj+Zp+E
caxRli89fgoQfNeXLncfEbEU/nco6Yds7mC3DrDEtLoQEmz9ZbQYaJEYM9YXwCwvBsHTndwSvOce
UcNtEK/cudkrq8gPicH5NbWiTwrMma7SEPq42Ko3SxR77dFS1JjKKegvh7fo8jUDivXA1z86nwga
jDYa6V0tC7egazjYf8InyHXw64UFzMO9SgOuGvAyGS9VQIaaYHtRxIgtRapFSWq9fcWlLNV+WLHB
rpz6/ZiiLtFhEbITSNpG+0CJbaLBFcnY1ePqlI5Rz8chgtmgEMEU+Oyt1rVGxPIvi+xxtx/ryvhA
6rFsIMBhDs/fSi5rLPLFj1p2owN2AJTS7bz39DUbI9GAdXKTr8i0bcImkXVvsF1ZvDJ2IPbiN1f8
xmCWTmWLGI/qmG8W+qRMtUoLxmLA3Fw68KSm65CyLJlU/0emAesAHqTWZF25lEHBK8AG5UQn6M+9
ekU7iX3RnI8AoAH1P8Q+VS8R88fUXV56M3DDIN9ssPMfZbHB2ZNsbUPvsj67C3msyxP+G6nJp7LY
5mR4DiscZDyXSJWy0qVloIHrRTC7qPKen7r7VphLcDx8BdHzjN6vS9x4cnZd87wBh8KQm9Ee8qBr
DFnWyoWsNl1MbayfUAjaoY7/CShzC7cA2dSNB7SbWuBqpFc4fu43RLdOi29VI8uojKdfqgHeH50P
y3YLylzXokPaYfcph70F6wPBYKLNrZjwFJou1D65s+q6RftMshocPIWFZtRjyjKds/XyE1n/QA1X
7PY1OmSxfMp9q+XOzJ1TFybLwUUnJPGM6hN1Id6YSrQgI+lJWV+D+U1wV8DHIeYmrZPehZqUwn6c
NXdltRhheLyhONdC4vy/QMOpfUSyOKcrdqYBeYmN3IqKw0ukFDuIkwyqBavfmoLG7ncnKXwKWF+S
DfDWkCpTMhiOmGSgSgWB5XtY8GJnNTBXjvOQ0/l3O+PTdGaEIpugaM//LaSfr1yAaa57B9CugRFD
2OEodzyD/S5s1QZwx804KZY73pO2aNq6Fe4pZ/wNV3rsDfepEhLf0vPkoEG+Nns1UHmj20cP+i2Y
d5ClklCOgOv5KtywX40G1bCmTDN9Nq0+NoNZnOWrESTHwA48KAE+J5dDFB/3sk/H3A9QYB+xI/p3
u11pkx62flbAAvPLjJtjSYblmyAekV+wo9pRw3fVwJaWK9SJsYQ57aSkdxFzob/qC3pkoeA8RBOo
TkvjN6TqZpi1IQ6hOi64HHg1TYfGes5fRr9UwIZKlYKZaZRMLehDzXE5m4yk1Zb5IhZni9NlQ60U
SZERb6I068L5tLfCClOdsHbpO5YwczbA7AxBFinyrQIEBSzQF1Vst1emLlIk55uqaK74qb3x6jy/
OkJ4BCmV+usWFim2//vEcQmHtr71m5/sAkQ/+5Tgl11hORQ8YMMo8ru8yvossegGxvcRa4YfyXg6
zxkGoR8VPwC+jsnNjRsYo2JCPQz5w9K4ttPXxi2K+Nv3V/7ntxYyaWLnxblHOc8jwmCjZm0vaYMg
055i1fYL4zmJFrv0Lojk+zZlh0hj0FUXrGC2FHXihqaWSp+SyhpEIWw7OdF9gDL6emEAHEMWS5Vq
Jpc5fflU6GCjmXf4b+43iF79B0rNjRjTeGnJrA8Le3iAp1QIU3JHxjMNikQl7IIDl+U6TsesXhtD
VtKai+74hNlrNDg0KtQpueLcoq+VlHwdXrd6csYLjch1glTLVD3oM0/XpsCVG9vsxgVJdv32JcnZ
gywnj2thiwwBcd7ho4TF1ezuTc1xgwGYHP0fw30kVNOBFZROwxM04ATSC/bgG0HV+IlHdlPckNeY
OXdTDpFVmC9Gw/LlJ5hDMGu4KTV91Wp48LIHqGzv+eUNOo9SdfV86weYDv+0zQAuKf+CjZfeSqA1
3oUNCovHj9+iEqX7+8Zk7iF8YxNPAIyuJZ2xQb4fquZWha5X3fENyQ5uvSIHeZPwQXKr0BuYHrne
UMN3mEerLjTz4xdEBUfz4+X4dtTUkP/ebtV7j769mIlY7DPxZX26ViQzylc8nHqiHzMOKIqomsjU
u9txnizHJxIjjSALR+mJOlHQg99KvLGN6V1M6+ZxvABPVPEqacMIKTORgaTbSPqOPpvX/jUsIykM
RqhcZiSuZiSJD+6o+3sxaK+LCxYq7RCSpHfCIzKu9nqCwqCzXdigdIieqDLwxnedR1jGv/vLoHOD
xl0Hu7nFRZwQm/bQYdqQnCr2n45U3QpRBhUs66hsKt1uUTl76U0EP07VatUat/Tyv9zNDDqChKU3
3JscYE1TgawsZ61k8ciV2oM3PlGGtwoMvyR7OWuS+qlG2A6cfbTE0Hs4Iz/g62At6lE0VC7L8lFS
O3eb9Q+5RiaoFnteq4nRY/sJcaPIwPbmCk2IvoYS6WMe2IIKAKb4FYEVZk2FX8j5UI+ZmQjmj8RR
1LBtnqmZUu7TNVemkrp4k6a7xe2OfcyUzyNQjEbVxex7yYUjmCMFMYvpifQgMXdcPLqe780HTGBq
rVFq4h33JYsXlxhwf6vxSx5yM24zTMqwx2Zg0cTf8b7d2gQesztrEgdCnhWdu2AQO+xBTKwwtApW
UXiV2PhMzO1p/DwKqIBRlB0tE64iuyHUvxGEM+H/JvHWJf/yvKgfO15OaDfehLcKVpkZ29rLKYYX
Ogl/k6Z92fEEcGimyzrg8SrnSAngMwMjSk61jApDHeX+d2iZFUD2xjzsoSQ6qyeFEa3GgofRuMen
WbvS1muWclhMgP28I5ivAmL1iGx4JHsxthqgq6YLMhzyzYcFqhHA+3VSsH0sJ8pR+wLMtO+qGC/9
cbhrcLggn0BLN9yaXT55Lc1BSRVlCzhBBofb0lIt+95wkMDm36uVasyaT6BqDriG6k86fel5jSZf
fS6Z5HmXpNwV/2h3qxkTGsftUBkp2Iu3FGpvS7Baxf/NUcoitZgCWEEOuPmcy5iC2kmtz3wdPrmV
FtXm2s7qIT80sgYkEVKsOpfHm5y7hsUh6t0Lp6K3jvNeFXJ4KEQuHirYRKMPwVb9IJWIeVYvDqG0
fmewhdiOJ+6oONPEMd1QBvMODr115b3ZQAuO72Wi1H57jvg9yWQTnslzNtH5ihjHjlB8fSDBIzCn
IZ6ydd9N+qGj9WFKbkJDyff/TFYO6SgNw5zxCobn7x+JXYNgeYQ6z2Zjb3sxydIUQlal0ukoCHGz
+rIpiSMWtv3rXQhYmPy584CHlDOzX2xSd29xc28Z8NuD0DY45kslsHC1LhYotIQGdZo9CA+bYuAF
MQPlDUARjw7DkOzq4bgQxAstFv7rNYoCkpcCdKvIS03SZ0eD+qeVI3f4tgAuWwGhwYWuBa/2CwS1
blJfxTbKLhX6FE5tg2AWMwjFDB3D7OW9SNrLrAWGLxz3XXY4X1WqQ4knyCVZxv32p674gma+uwzz
wOYKlGwdFuisl+e07J4J/ei6xa21q0a8L7pYSV6W/kXpJdzaRJk58X4rePFFz/xGOxl0SjEoYAKg
fxzB6oeZl8h20aZQTCV4L82DUdUz0t4aOtIuRY3fxDW+ffC3D4okJ+fqEL4HsfJCSACXsNAFz4pq
O3dRADo87TxhMRZPPcOj7p2bOSEXiSvMaY6i8n6haZWGyg/C65gG6E26DeEyuYm3jn/ze0aKRa8i
TUAP/2YjPkG0tNs+qlAICG92KXXpuYJVwHpzG1MoOstKJrEqUYmEojdzuD4py9KoLlTHsNMMk1tU
NPf7NMMR5c+KtruDUrWCmlhqupgmr8wQ64StcvNTFuAkRHowuJrvdwjsYFT31/m/DySoX8jC/kzI
x/6Az4/TlMAp77MpD4J4w7xYnS6rTVkuIiUeNzdP7hC2+8VAfOPE6EIqsiI5C+yNFTofibLDz1QB
fglPnBJEY7NW7ohj5oNdBgd7fmJEbqzSIL1nKFEZbk2+3oxlbYSJvGU0IpuQWiWqLWLvmx4JFsQQ
LxoKCBsruFxc0icmMjmG/C3N94Y3rAFdN1tvTp69GkpufgA70lBeVs3dxaXmkMUE5QPwJLvaGPHg
lgZFjP00lbMp/8QwsHWheJfF2PgMZMvn7Awg2wDflArnTlvI+BPxkTHaW53dJ08CaSnWo+yNSUTC
PEwqGh/XpshaYcw5rUA+ETl6mLvMgSlv4He7Bb27v3x3JsshN/ao9bLQNLZXvyAI0qg2OiwD/UjG
DtL2gSZ7m6n+rbesOOmBStoo86qoiz+8btnEnH89LoyasmgEfjI5EMOeKl4mJlD5fF7lMPJJbu2m
mGO7HcDkdpN6KqlY2DrpW9kVLTISjaU8nC3XJuvsRNNn4BA59aRo65BMz8TZaBaLe6mzJBV/vsiQ
llN07PNzhC7aZI83sspcEs/AiU9p9Aq+cVVFpJUZiGWZXkWNDCVmPyWsnJu9CM/BSyxp+d1fqt/z
t6VG+WEZQjJ24FeWo//5JK5Q5kJ4D+LWmVAlc6mTXC6TPtWY7s0yOb9gsMjaqVuLDB1m9WA7cuhT
FJbfXv6LK/xSDn48mn2+9fKEoGBcQGyGDM8BCPrXv+QnicMuwhkL3QgDhqIBUyEb3A7n+bFs3PWI
+x2COfy8d6WmoWoV/6nvXhlDbmVxSkiC+dkilOXROWXz8U25PzDaH10k8radIl36ATWATiw0eIow
T5MZpJzRJDe0EPBIRfVi9evDJDBV28Y3siC/L42CMyczbddyFB5JeQsjWor+Ix9MPWXU/C2W7Dcp
y3H+9faon2MH4UdLT3l+M8fBZxXsV1VlfWWMok/npokvYaHblR6jg9b8IlIDtSRfSSObLBeQXQ3s
pIzsM4FDF/ZbOz3c+5sfP3gAc1ia5+dBfArA+khGGMutJT9SHdHuhRw6zvg0MFQhV4VtDg1QsdWy
Molh5x1Ml0CSYFGYDB6a1yPZOV5KeL3YsbKPuSn8odg54tYFDteornoNVR40ZP8ow1XsbFeOOA/E
XnycVRCWBO2fzDMxEYF0wbkQmZBcxTaCHvbBPyXa7wKoUI0Au/yGDWwWYy6G7hBymXkF8uj3ZyOW
2TmAr8/TkBHrAqaiS8uBH4hrQDW8zFcDS8Qdz7iJlZbJlBEiYFB4dFBC0Lyyjo6hWzEktAxatn7H
uRO7WoZtn5Wljqan0yeXkv98i33ttFMHGSJF4S7Hc4Ii7Vl1Q5L8gLVbVHAi/U00nV+qJqIE95nf
Fz7UBTUDXqRL7dFciWcAitCycwo8l1NWYmBMENmy3JvDcJLfSpAfs9TSpoBukdT8ipw13b7/aw8P
a1jJyJY1/FYj292svhiCScsU5uZBSnJ229WilvvhpbRtsOSxosbadkiMLC4W/e+GHm8NM7AO/f+7
YaA578DaPZJRcSSoCj64wRcIsnqkyCbEOkm5VX6DVQ9BGC7qmRsXpO1onvAGzIrSRhtz1tcZc8EO
lS41AQBm7R+vZ8otwQ0RhELoDqypTSTVgy4hDjxPa/ZfbQVqh8WPkkwYyxAgZ/44jIRVwadI+MfH
1hzEaMf8PEhd9BRGGvB5lXKdjl+7yEwq8Cs+mwsZfxCLNX6aMKec/b1M8VvUDvq13Krk7SoqQOZw
e7P/GYXS4whNkDSJwoAAJi4xEcsnaGFcuXxThENIDdMllasn7E32B5ksHCG/a4P9rkxO6VvXS8kb
IUKg8eNUrxwp56+sT4fLK61HZgQfLFMMYXAQZKGZP3oXSwL2fBYXiElpiWC9x2VI31jV/F5CCm+4
S9gvATmhWRzthvj1pzMEWXVgt2XQZ+vY1hOFLc2jvDhnkeyd/EZoZ+KONh+xOrtC33qEvQOK+32j
TqsMguP1qQTsihRgbP+tAHFdQYJvUkRgt0A8on297dSFg2LDNQ3ACOALhBiY1XL/T2ojrTHJ45Bk
+i/AciZAwpNi5tqvMmE/Q3QL7zsz4YEXbhTTnqY4HQIATVO6D4jPsZd7euItf8u4vYKzspFb4Nra
94VIBISYIr+GKT15ag7vK6xhRj1PJsISfNXzgl1T8j+OSatYBNY8IrvbtigeF4Xj4g3kvu64V+Rd
jSqqEKO2pbYIKjV0qTmAVSob6dEawbYsJI1qcYj1JYSmcF19ihiETTHWk9bIE0tjN1fkp+obyAsR
t6b7RRtVHY5xpE4BLLTnZ3gDAPLM9EiNjkDf8VBy//aVA7ZfLFqhsE/QkJpIJ4k02NnNtF4Ij7Dt
gYAU9/gVYHOWHMZl/7AslqCaI6WoNWiU2ge4kOqfXwCtIg3NvNPkF9lqCKH6D7ZVBM0fNYqvr2SV
ijE4csKwc6SdWvhnWZ5yv92biB9Zi5Cm7vIo05UWuy/6Cg7/VnUsAigUbJx/s+l7um1rdbigifZn
isLAipVvebihqk7Rtv6AAXRyRjLRjA5u4PLb6kwNBJJR9JJPfT+oiBwEXElyTDpRqVJIvfc67oZX
/KCivY6BRO0MHFAwOxhskQ62oq71yCY4gyrNnnXWk7ZMLHSCUoExXsXjfuPTdSLJ+wPOy9eY6R+D
Sk0DErzADN2WsPwbPH+8GNWy8NvhbMXcv82Ou2whotb+omyzz3LuSl7EGg3LAjstUYp4dO2jM13L
KR4rFBQqmcIgTjYdlYKy2rndc8gQVdY5FBLAd/aGHgBUXb0iN1yldH8J9pkEBpOcnQ7aGiWzHlRf
eoglewxlvrSqx037JtvUT3F1pzPA0jkkOVeVWMD6jgo2yLFXuXc2dIyj8IlIc28eDVm02CJWfvt1
ua65XXF/GlaYGLrThdxJKaXgnxrIbi8KyffaNab3R07eSh3tKEwTyDWxC6PWolbzREeGf4j1LEDm
s8jvWDFME5IYiGxuGW8i4VrNo+4vdrVP7GR8wacC7+oJ1UY/M5e1iKgbOYfQOCQ/DB3UvUh4Re8T
Lv9Dc9xTWpU0gUuCLb6y05nwIVEEWxUG3lgCsI54CMK5QNq3WXXaKHFZGrbCLNhYbFOzkWj3mY7Y
HFkYoyoSGLA18K3Vl31VbcuR4YUqT9f7xv4ZGbctR/GkUZ2V0Pvrqd+5Heyltxv5ZrfqKYusEdsb
QX1KPZiyVYWDpvr8tRI5mmYPvclXU9fH2NFTQAdhETp2JBD3tdcrPjDIbu4/hLBRz4E6DRlVti+o
FNb7T1u8biDnpbjvBy8tr87qvbBjCDEZBMki6qOLr/RYFphYJ/xttJ4bidoeSQoqDQ8mbO6BTyqQ
nT646ghQzYIMAjqJUog3MqXKrZmsC6T2L/r5Efh8eQgmCsaVuhH3hFoZ+4pZAyLrGVeQ4Hn3EJJR
w4x4M03ir/kqGak3bjb5CWT1SZ4czp47PUURxshpBDKOy5EwP1pjrEgEgI49EjROnUUj/K86pj1P
/qFiNY7SUrBd25LRpwZAA3OyjgJij+UThpQac8gPbSxSIue37Pdg+kbAhonWoAXu7GGdHtmeiPe/
c80HDPusZjJrf/TDuxOBdzTGPjRYTgtGP6htUwjpkcORWihMlGEqQHs1jkyUVBalXydOgW0utgdK
uIaFt3tark+ksbTqca1l/Cueg4VqMfDaVTibdyPSEcp2lulPe32spkQim+PsIJWfLKWLqq3mMGKT
VeyCUyi80tnRt6JrZW7OO+Yw7koDF+czekpa88GQf0RfqwnKDrAbvbllO3YMY/2Be1m+kgj4wwNj
lin3HvdK9rBN/HZLRLLHWIoUrIBnw4Cj+uyaOTSEOD/eOjtbgBVJlOsGnK2513D0/9Qc51iuG7er
Wc+KAiGdnCdb7TL4lotouSYsK7JKSPMe7jUUz+eRHrsGDEcct3dK9v3LO7UxsCnBaBf7fRcdF+e3
luMM1qx8NR6XnBiwHIUKMb+rLJUDMmZyx3CBE5JqzHhRhHOO05iTVgbmDR9Urxrz40hAORXeVz9z
c6CCCBLlJx8zXQD3iIKIMHKVjOasN2eYYKCbDH5eSs0AcHAHodqGR9UrOQcSQUUhfgEBM8yxKlqI
czC7v41yaPJbK6ydW+yFYy4nNpEhShwQvhd2NFcxYhO4Wnk1cfXrhkaoZccsXEHgXBm9u5Zwpatg
r36pR9vxN9K24U5vKDSi+WUbfmcqzwkgSGKB6Sbhavk44dkuehlqJS6xPMN278h24ATHBxRLwzcu
hhodSMyy5tZEYR12l1NfUHtc5EjitVBrsvWd2/Vi13U8VBb1HaGeoI83k8v/DWeF4aWF3/UR3lke
shtRqBglaLuIiHoFu62uOfKZ/iyebPYen9M4qNyx1SZuXy/sOwXQd74SiGi6RFsLf809hLn16j0m
CffyjQAWuPaRuKTzA0642vT0MgJZkdLydqgbtQr5iEHnugQqAxqO++KPWwTSC6u1YIznSwwjwinX
DHI4WVMXjKzrElE4KbP5htJWHvL9hAPuWWRnwyoeKpUNCnqp9vM7QoG80XM3QakmW0ye9dG8d/wN
qW9YaFMYoZuekHm6at0/KIf+w0YXdRhxnlNKeX2qTCeKfvgxOeLhj979VWEsklwMMiuT6EEUKizU
bKmVGfYdFfw1ldosqdrsYPrIr3R+BGF+8HUoVYCc3io7Izt+dFvFUBNfYTDFq+RX7mpKULOVRl+6
zXfkR7qEJO3pXZKnjy8EXgaP3gl0WtIWpHlhP21voXoIZ7uQQHwZFGBx1TI9aiNlMA5n/qvDB4EQ
iKmWVwSW2waEQZBg/8b/5vngmk5A4xMHFftJUOIj1c5dKgYqueIo24XjZ6py9kVTeL8DRV6DsC7s
CWoru3jRfBNZHM70EBe6A7E1ZEBMeAdKXppGdczsIAaKOj2NOGijNWagLrKP+0nZVZSK7Xcx5KVA
E/uNd2g2lXiSgMl+AA4dobNsqIivoZfg3cm5AAfJZDIayxNpiEhXD3tkx4KxNaC2QOUh6MRLmvk/
yXdoPcduS9E6fZyvM2nW35Yreyt/oQHRBBuII3/lEZQoopJKHtx3vtyBAtIVtAtMQRrPIVv0hz7q
SJNtMXCrFnLk4rE1hQ1CaV/Jfa5FfrZaNj9dIjOxZbT+a5EEpGUJnuDcA0txx3dWCZZ8VLgdYOcd
s+q81k0s8elg1YRErLzLZAgTRW0y+rgLz47Hq6tm+3UKydKQ3mWQf1YK5zMiYbaCeUK3Ld05vMXc
B2cLHrQ+FnHeqw8GkVW92AL8IIQI6GR0B6ujIL/n98mua8h9NmLn3YRfwCZ5QGZeLQaAKFBHrsZH
1JCv32IZvPLrcwr3cfnoD7mXD4kAhDkCMHBu+IlxLbeHJ/7bOJR67W50tP/JZ40R6EafXDa+zmNq
5bl7ybykrbFQ4kd4Az+EHwvNeBmbBHzqX2qf4v2ib/aIzXb/iXOw0wbPgULbzJ8Y4PiFZgyZOWI/
JzriS67hOD9ShJvX0DYGGtlkHmbeEVAGAVHEjnFNQ1mohNbUehJGt+jNSLW233LP+wgLlBg7V4Mb
JM7DBTtaCR0+v4KGlkwA6fGyc5qQ6ummtQwHsmSYU80GlXi/F5aRWusm2lJv3TfqG9TktJycDXeA
JwD+FMFVMJhDwF2yTu+MaggWYJUydzccGbsRz70XhQ+qa/3+t1IZBBgzoc3X9QTpezwUTcXZKhSJ
Lj4j2VwZ+UFpwMkJFTm8lYX7QHkrsqzAWnNZaOBJ5f/Kipi1UW8YsFoPfRNX7NCLwRyXEp410bOg
N1uCSvulVLh3MemmksP4IfQlp3eM4RxF3n6uW6n8h0XV003utr7yDcXMfwURyAi8LdF2ELmzomgi
IYq3mHSt2JA43QriA3UY+nJDoXfy+7ybFoIvMZtDe4M2ynj9YazwvexcDWqzlhAzKOzI4Y474OaL
i8zrdKQwioiwHgVTiI0+VOVE3ID2AfPfCZ4g3iVH/+oUJqh9ZDVtVRv3EOsFF/o42d7717aPLLtN
LVt6WaXg6YMsP8kqg3XgZX7byVx0dUHMt8ZTz3EajvxTef0+4u2d8pbMmCYGmMFaJOpOHhEFsRyS
DThvKkzhuiM8n1IsJQKMDFUMvoQgK6a57mM4RrIhdZLRZs+106bxoE9hKjnaN0iHoyj2aumwlvnQ
cu65uawe0eCfSKxhTAzgLpQt1aFTSAm5X3hDfdJzqYG0W7HH+hCn2EBhwg+ijje/rpfM4tcKY4DW
ReL5KzKzFi32pQ9PbyBN8PH6Rau4DqyjQOfVgqrHpT2S9cTrL3ikFRnbsQxFv06lnKXioT2uxaQa
DvwFH48K8wB3RN9KRVIibNsrhWbwALrReWDMCRe6TSZPsOsZOqO2CyTEz4Bgu98eA9cBgJbet+Vj
EQkN/Fm2jK2uV3sKT7cEK5V1vJYMG+xK8YuNGETOWJSEKxdKxr1YkGpf7TMrFqAYsVDNTJGpgXQ4
vE5SKFIzzyOxN3PmLwXMGpDa9OJOIsy689fOU1MVMjaz7u5xVgh4ZHLkWRmlXbCW+1ufriCgjxrf
y2gGVn1g8jDwhaOW1pBKWI0uk38/YfrOh3/DKZ1U4fnuSj6lHYbKHTXs32ohdh9annDl1rBuBX7n
BsEnlUcLZm2kDhXbNyDJ34izxTIxDPFoCSP/s2qe50wpzb+9FLTTYcK7FUzh3Pej2NEx6lRNabax
3NCs7aJaQLoloTZpaTk97EwkxaJeY+JSFHuJkXHrvhuqdR4rL8J3lJ0VNkpsE2rnIALMe03JCTXv
6U0FDaW3PQY2D/TsyhRsbjUwc28bBhAjp4yWQHIIxd/+bw9dVXOEP3obNbWHDXbpIHkXBlVlFTLb
7mO33t6ZyJzlo5DelsFy5Tdu9S9495CrSgnWHIgvdyyG27528LeDwUaFv1kGpONfeOKePWfqaNA8
NuUaXlMCzz0Wx+D9WtedSxL2E2QUQU0H5qfi3MrPLzSYEZEsmhnZiSDGavIVbebGqlSqgARb8G5O
o04k4j+9UkqrDzd7dwKYj4NFz6HyQln3VbMXXrr5J4LCgN122DAqIOdZcGxTXM2r842lRCtgReyo
MkNGyhtTynws9GBINkZKLk7p+RcjTVl7lQ/EcrPt87mn5I+BAIIKyh60ZGCqfUo0X6D9mc78w8U4
By6sVAcg1it5PTEAfdPsiykBXXtXZqWr8TZe6Chqe8HCkqV/rLkC8XLuFtx2IO368yhC5ZlihALp
IymwvV0qpb5iLsr1+s9tcHgIWADXK3j3a+YxENw/c18J4n24rY06/kQVSdqRbVZjBJjZqu/uBK9H
dMxzYoVzUJmWQoh4UTfmAOVCFAsDF9O6KbvFeLvBKOynDb4y7fThwh/BwjM3zTaMc7V7jo3b9gyk
xi+mQdNZ4qLdvFxkQ02BFRiUzAuPYvZZ1RurfOw8Tfd4A3pHAPP05uGtjDeNn+c516pIc0LZ2qbE
AkYR/swcfrY3iSTrWyuUjjJuS4DK409P1Q5U1+Vfh84r5u535IxBWQThSa1yFLKAHTC57HzcIwC+
n/84vlqfkAC4LhznjNfopDMretqgzF8qu7JB7wE9e/kijJYP2hDk7tjDEL6bkuPYLguF7LsqJEO7
lvEv3yGCj0YwXBVUFOxu4NOB9F+HT6I1jF6hgCf8aijroFJXLcYqupiuNW0qPwhLf7f37Rzq0NyP
BnKQvrq58RzzMArUQXimQd6lLRNlkIRz2VU7a+xDhcFiaZZ/HtyQSoVLtkANH6CloVa5By/xYmfS
zKvnj98sUdAcV0ACBqtmmoGlkv9vblFt6GP8IRlAhqbs6f/5QoWfa+L55GqWEoUD5JwLEHm1A5TA
KNyUe1eVuS0L2Wgi8gFK3QwcxTHIuh/vTSyhm+DJHgCY3TxaGFpTwbaKrBAj9K+4XkuklPCRD/5H
VYqzRAvhnj5FC8WDYIZYQBCTJEdWcjzWvbQ+vtRyZzVh/gy3GMupkuiiItzTBa/5QcQu+aY/aD7b
MgoAZD1ZXLpxNd8XfCuUFqPO0K0YHXwv/lEJarNdcLl+LleJf2ofefrP/HR0J6/ozIa0jpaEEaEu
juBwJXEh8LW2GRF88AJAyYp4FzUkeE2fQ4Rb0B24daC2PiY+LHmKraamH3tR+S/xrL3QpD//jylC
SjiPsSldvFNCxmw3GQq22/+O587/7Qh6zUqKH+KtyeUIyBr7YU+rDz5D8ylG8mpqm5KJekt0gYbT
QwK0hHNmfkTfj87KPuHm7TN9tWgOBrg22k2ReTEXUqGtJ433u/YG63caPRQ9GcULDmVR/FGb8kvy
ZdghYBeEdi37J1gc6LhjgK+H9Z9IWtDKyW4j8YElb4Yq/PDQShwniYg68VuGlOMZzXuL+pSRU27j
RcTTw8A/hNg3OcKRVQbPWt4WqDJAc6Tw1HdRkrmhjC1MhcDg09rL6CMOL6vC9frAVt4L+VzNh88i
ISsOtj+ahoSGvQeTeu++FDPdTnNTCT8Bu+rGGnC7LtVycdInWesGhtlpZFyAwLuJ3SzMctnyjBTD
3jImk66+Z1Ntj6iy6hvX8xRSBwzjGpwhsYyOvzmo/XVmMp4BSwb1zjGeOielngELz7rNI0fSDYrp
cPIF0hs3LKGCn11UO/fHlUO+CuNB7/MQ1GKmYTaWM431TDBEh8aR+1ISgBMdO+JR8frJQ1Sx2prJ
P28kr5KCwrFVMA2BiXW0DxkODdYB2gxuciArUwbQrIdXA7crbKlQNTZ7HE1/iqtXQKktEUkdXdU0
spRC4gMwYP46eXMDTA0bqWDiPsP5TPufTovL9e9PBjVt+LJfIcpxPgtYL9znSB19y7QEnUB879cg
xYrsBmlo8ppyriMaLghVTXIRl9jtxq8FjG0hF7CpW+yq5GEd89MK1OSL6T/B19J38OJuR9SrZbw5
BkKuW77NFjy4rd+gAYCGM7QmTotO1jSvHNgb7l7xui85f4iBdcjfNFWijwC6bR0+8CblJs/F1YcS
lHohboNcIdbRlzmeqt60Vbe1e4u8qiZOlmoE8L1Qq6tb9K8Vqe+OyStX2wxd4cSg36slj+boUplh
g7IuG796Hbu5n+Z8iwc6++gKze8U/IRZaMlLfazS57JddjDfigrFmigD0PoMcQCuhbUGdWyJ4I50
Zqxi06Lv8nwseX3oVfo7gUU8tH/53rbYNCWcQltXIG4SUYoK1NsKCSK1g+DENZpDR/0qH0lMLuse
JM3A5XV3ufCCu1AcANirNBzSyU39cUfVQCNQf4ix7Ea6Oqko+Y8dvEJwb0gbDzgRILwTrXqAR7+n
9hMOhEn7+dr4/GOczo2EhUHHlBvQwYtXM0JIkeAB1F+WKw9O8TAwtY/LqoMiF/zsAaimyEMhdm0a
fb8yCCu41P/SG7xNMzSNUZCmzO0wVrHAQ3Jo+viYShKK1ojxkIdRqD1iX+pY0z05D+Ltg3FXQTKT
TWZit730vcFOqfzWE2SSJp0nW6Ik05IFMqWBRj0TwwCq2gWGgPcAyUKB3rC3QSEG6kPKhRAl2iUV
A7MvWpNFb5YO9j3OmAdLUkJ5LuMQWSDcCuG5Q3TDjMPuVuQnkcX18NbqMmjpR+d8ad0TJSfsnZ3n
IUvoSeOFfqJ3MiJE3F2sZvus/quwoxxbyejewxMd113MCPQ7/WY1Mb9WDhkXiNfEX1wjDelJ1Eim
XV9wgfoOwpjVLs5C2ndJFY+Ld4YdZheRLDHFGP7OSZwpLGhPttiXw1j1fvWsDEDQ8aAlwe19/RWa
oZ1csKqh1rjBgkILuauB6pdZETNRdLC0QQ6C4bJslHb4TqCAw/uCxILqZDEktE2BzS99+GHbRKdn
eaWO0A3na1EU9vuMC9dKWifrVbaRZvxrHwRTioWTZRphrzzF+s0DOI2CH3y1F0J2WB1eLtPJM7kc
qIK6g0ATguILyltD5RMAvKvl3C8mjWwJ8RxXO1qIVGSCATbtHMT/cPsxPcULQYNgjHZGXbOQM8Bd
ScoOkSDP8MlmW03Ihdapxe9mYy5LxSUfJ1QtWK6P8aK3s1MsPBBQG8DOpz7HOWAKw3LOkNWVVa8+
u8Tphni3t0JqNCEmJ0GwjRglt2peFQ5bP5JSeesSk3OXFePIfM6k+mkWHwqa8r5zOTqHTpxkxSw0
+tG1JI6fnaLsclrUQS3aOvxwa1+hV5szinXFABgnz8VSKRJ83gUN7dc/oQKFC3oa8jZ1Q5lEmwFx
LbiZYKW9A1vgGmSxAw1KGc0Sy80aIG8Tw6Dp6qFCnqY8Bwt3fti0b1pyiwmATYlrBZ9Vbi/H4MN7
bZGlcvx/L733mU5LIudlltJCxbll/WAvmcExipdVfe87cbNez6lU6RLlfcgRwyhTj9pA/XtPTL+0
KU+kNNuorRjzGW1xIGMLGJdOOQ2t22GcXryVHsQ2InCV0Rg4DFc2j74tP5kSAlIFf0Fbqn5G/GPd
2C2D5hpxlWmmne6aiFkzwAN8cni23AFKgR3LHmKHwbPqqvxVTILmrvzEnA1wBMLv/sBKRIi6hm+B
8XM4D9I3QgYsMuapmwVHqxhK52S5E5WRzCDNC1sMrntfX2+WdAtRlC9ElhbgUXN9QWLfdsegJn4Q
B8/KVxQOnlyOVI3lBkPt1xHhvegyZPlsPQY+myvHCcjS7JfAiZhwb3qUXIYJpy8Q77KxQtg/+t+T
Lh6XKl7TkEj1ZP18o3W2TpNrFqvNzN/Lz00va4BYg6F21Ah8O6t2X03OfjrwVEGggcP91v7WM1fg
FpjZ4lhKvAJY1y0JMuUehRQ6fZaaj/GtEKcDrQxhodURkYFLoyeMKEea43VNJeUZa/ATnpoA9Rq1
41V5fAwrSSY3eEINb2IOdXMXNDFxRpypAQSpvBIMMNkuJOQ9Tea4yNP2rn6SYYaSxQUrhADzB5IM
1cPBHdcJyvZby2LNR8tQIyEEyvzG1gb9TTXkLy4xYMjiDWjZ8qydv9Kl/80qunbiGRY59sNEijqb
K89cKk/bQXdSFmilE5Yg3N0S+Gq41eZvOtbvwcIo4bQIOV9vYcmkGkP95JUzahEKHbUcOKN5/e87
qvH0SA0PGgdsttMSArCJQQjw16Sw752Pf5eM4AzpJQjST4LoJec/xGiNO8RfsvjDs4UnD1UibID0
+w2Qm6DpeL3BR81Z4GHfTqE++qSxGIju2VGs2TL2s4zmvyPhlZ3OZpD5s/jgtYEPqKDoNAso4hjB
Woo+sxOVb4szOGHRIkhihrpVP8hzJUA/1R/++ZaBbqzQuywkpm5LE4x2xtQ+gwG0p9YgpTlq4grY
B6srA1BVgcrKTjE/uIRYqUq91HiVK72PF4EYPV2N1I4ghEW92UjOI+mkSu7L1B67aGalNe/hpp+G
IzrQ1KQnmqHgVUH4t9V+9fXM0U5yALYqen3XMr51T2J+lAJGCUFb7HawsA7+ndjMaXOPuZSZ8lVD
3HPzusyFRMUCxspXQ9IO63Z+ynE4TbYTwY2A767kSSWfGQMzujyazPMtCF2pXnPHOlTt+a0mRm1c
1czSqKQ59NcMJTcd4I2K/CfFEB2VJeokOVo0obqA5bP3Fw3bGXUKkBPl8tbEZKA51tYWieJgIJKv
KZbGvXQjM8+SIsIsTuJSrsFK/RIZmm8/oj/oe95Y9I7w3Cxi5suzeYwRtoLs9aMT1y5yKGiWLs1f
w5ut7EkScjicJc5284eQVKOajUza2gYXMj3HQ0SPuqGqVsa8oACVFWt/rw7TwmA+mO46pxqhZZcP
ylpkYs6irjqfFCfPA/qH2Ndc9CHq7/YiwW2hsD94/o1XLXq6tVLUZGFfjHNFn48muacA7dJHOS91
g5TkOV+bVwpOTmV7FeDOq8ZyW6+sMQaolEwIUNnSUNHLGoyRCn8dvIHw9QlpuMsoGdEpAP1kM97H
fZ/xm7XNsEnVBoys4gHT7c7ps2L9obI7QOWnd6p41F7edy5CfqM5UyZpd+sHyadBwPeITRFAr6jT
2/cnbTJEP9S8owK/ihLi7V+9oyBU4anxAVU7y+79vifLI7Sx3qwnpxJFKnIKxOGCXHx7941DdT+A
9Tiai6CEAbUyqmzWfQCxZMebAxkxPklhuj1uLC3Jg59vWH/UJ5YJdlr+tQ82wTMgnXqjQCD2caEO
F9UjnC/BZPsT9B0WMyiH02zsWc5f9xVMR2frYn6i40d3AhbJ3zidly8or7ArDrtHdVf0YgepE49v
E6MuvvSBqBLs57+ibwcC/6yDY+L3R592fk78SCCQ4VxRAchAPuMiACndf7C/xoiP6/SP3RdeYoRC
XQR5YCGSsuHC0ORf+aSjlGXdzhSjFKr0Dd4a2/0/N4dU+CIAk5mTtqrZaZOJ8vYbO/M1Fuqsso7a
h2a7tUh53VhKC9RMJW6hlOVVrhYFjxMbLVSOvmQoxV8ai8C2DswO/TfhCS0NcRujC/XeFs15/5xY
Qn5hcH0CaQiXTVKE0dYjs7whubH+VLZKDCL/9ezP3QXztHM8fo3XrUHuBkLQh+jCcHpeEkP5QPjr
Rlr62QscMH2kasO4x+NGN9ZhNPqNvaUmlVz4ftuHffQ4zcsqqIN71eNoSyZy8O728pyn+rYcj5KB
8hKCMcnWiVOqhV8qQ1SF0HO4E79nlvVpk//ujjitnF2cQl1O/etdsI6aO2JHVF9sLd88AVXWOWah
lW2QPDjhJWpqU0o0vxt1Uik9MPWD+juYyXxtUHLhA8UYQVXB4ht48wtuGaGj29BZyIGcu40IHJGd
Hf2HVMz7tUf+A+M+AoYKWbvVPo/qHdz3AvMLhFDysjyGWAd9dTVNBUyHD56EeBaE67ndVjI9lqiE
3JHk2jOJg04bb1+cm1CG3c4UF/bIXAITXlkbpDgwB5E71z7nLbvO5Cmr7q+mNzkLKjtkjmpF/b8d
G9hqaiWnk00Mn+cV4Cc4+E4JYcyCgqgJB7vAG+ET3olV9qWnapA0XnGI1k3LtTVtEmMDBVsX8SP9
BivfrbReVod+Vp7Pl+ZiL3v1mhUxxkrGT4a7hGerNKK5VrsucN1juNSh9vV8rIhdB+IFA/qESe/C
uY0ZiZ7o43BXQ2uq+W9Zn+rfJ7Z6tiC1WPnbYHN20hSNS8/63ANMjJpWKZqF8NHUYcI1pIXz4Oup
OWCYXkKQoeVXHcJ4yr+dhAO20C9kp7o0S14v+LcyiCfMVVZiaMOjZqVkQbTMqFxkivCvdZQaC5cU
oQBCzLmGlUc/y7TVeaIJpUBhJmufr/l2POvQgT7UVb7eOHsX5iXbBHhm7CmL1TbLIfKXof8YkCOo
ObncEQDPszvJBWorvycLCWCpIQWAe0yMk5RkA30NCpL/a94+8bmaUx3NPaqVYppTEUjDwgAau65I
iOQu3xRUmd1JRBZUNVCQ9d9h7xX6KqmVgyffR8pU4fcyVDoIQzwmT70yJpOr8OlQ8PgGt2FxgXTi
Ohs3ZXaYAbh8gWTwTgdz1BjNEHlnIl/MiAh8d9Q8eG79SrG1/QDs8UDbtzRkZeQ1x86SzJtOxJx0
V9SNa7+oij7s6nxEtAGJGoJ/VO/Qstu+c/ioBSJwmsu7dDLENi9Ms0HrQ4Xcseg+MbhQbGbc0sFD
xPswqo5go5LzSGM0acdXW5VffTVnjiNsykXpbdNJGWrscUOG4oavwRbjgHtCcvT/0L8YVacqq4sy
3wJVWxafxDM4l8vq51vOU0axbEQns7kM6fFgM3mnOhskPlu10K8CuLgVpBOiMyfr3c7GQsk6e2e9
3qqqWICLDNR2XbL8aOz6fUNNdKJBDsq5cpDCytRClDukYGjz5jGkKih6zIUcvyj+M2ZtQ7TwwA8P
1i3Q/Zm6bWQKolVg0gya/4PFPgMIoKb1VTD6xg/cwtAjQ3za95zdOD2g/Uq66/4m01v4nWfKKL40
+DYA9TdLvnMOJWypfPgH+R2rqr6qDio5OODaE8Y0gXgbRnz/0JxXJ5cSJ+rmCAhatGJ+CWLyqbfb
lMldJVqWDH34pIChLXphv0MeBU2kNTLRsGN4US8kjDhHk0dnH9gu0ID4cljcgRZIlYi8ACDBeQeZ
/1P8/xfcp2KpN2nyiKDi+4Ss30KrK6Epa6oySJuPgaapW1Rv3GhfANP0K790Kep4bcOpii7A/wY8
FAa19vEKfTgSHi5lW5yZQwho/GnKQTUJMPb3uqHQRBmOZySd+U9N0rNwVb3gbat/oUKgnKfIlrYl
eV2FI3+hUu/GR62+wWc89xvjIt5XUj8/x9gH8wPEXdCJoXHZ2fli1QhC5alUKXSzHtbPkCdkJedn
6obHBjcomnQmK3NBs/fADzQg19JWiAICk8oHAHhqqRmmbO4Cyn6fu12MSHndKn/3Ms6h8/IsuvXa
4el1+m5fyO5Go+Df2qSNIdYQWElYGEBLk9o89ZGZQjU59yT0ZJoEHgGN+TvnjguB7uJU3a1vpYYP
7eDZF3Jt2Ujphte0IVoNCMsMZnZZA1pZZ7W3uXmzXJ4LrdsUrXYZe6I1Wgn7SZSLvXhx82JITFDo
d+Y6r8sACrvKjOLVURSUNXpmvlfpb8ZQY1WtMI0wPJRAl8rnCtaEadMzY9ac96cYikxWpwqpq7g4
HgjnFZAcYYNdpKYhYX58tlPDLgEEqqfCJi1ePQ8p13QcSZuFcEyi56MYPIipzPkz6u193V7HSzmZ
a7NdQaf9b8+0ESlJmq0LqRc1YwpmraElwomJTXj04wKnSM9516xg3jIj1EEtUxxfMJRhSv8+6RnC
UsR7VXxwU2g73DJc94EhEOOTcLJO/Ai9RqtRe98BQndCw64z+W99i4aAoXvqMt0keoar9T117erU
bf0YvHhxKL+OKSa+MSofn3phktnhzkG+LgQ5XIUook1iJBHUBm2p2ygnrrdIfrQifNn31lLJXhjj
MdF/x/aB/GpqVwXwsqXcWZ4dORFIoqHIZcTnMODsGEh1dEEYrga5hGnOidiRn8Zt6Nrewbv7QoRe
r06y966PG8YV5zP0O4hqsP53XfV8u2w2ibetkgsVR+OtnjoGGAsSN5vFFLF8wpLAp0CuZ8bKhKDf
zoMwWddVjRAeFd8BIzS5h6GLjWUODwojSuFbioE8xan1fqmWcmMczyOS+cj+R2GBKVGE1R3Ae3PY
qaaOrz4l6HznEsN/RlVvUOfFAaLGevec9Jv/EeH+f1oKzMrMaRzHoWjWwFISxLJ6+PQTfRD6EUrZ
NatxeDiMttAs84PBlUOtjCzY+SeRIeDhBpr55Gr9w1clMAOLKsjKidVWGUIZXnGFd74iRPJroPyV
SZSDQ3as2kzO5rocQhJIztD4ng8VYiG8sPj/3GaG6xrT5HMZGn0rqx+TUDUYNowhyWn2ndSv/wQK
psCHg5DimfXrN3n2iIR0EMdqIxTznXHukz6hDFoiKP6fOH9pU5t3wHQ6s0g9uvO1MK5rRnGmK7Pl
QoMODfmAxaFXMopT928sqMRd4YtkztxwNEJS94kaMsBs+nViQh/BTT4B7DHM4fqqginjGpQExsPO
ozdHtnnWIX9a466ftiJNltX4IBKuyMWB899rCk3gm+m1dnFqjLimRCHE5/hJbsY6Q+Hr3OIcBlPP
u9DurLrTVbM5hp55gZ85TwPlwzRYZFjrsja3KmnQBfQI5c3CPTUUMzmqQKOaICZkotAX6vtQxhV+
/suZ3SkKQigjG9l87oxG6VE2muNqoCSLaL0iukB/o49NsDc8xyfUrPKW20Tq6V4AJ5OUrAAa9g+1
fB8kBMgFOOIO4+lU0A7hFz1T397rrN6V8FBVN9W9lEl9Js6IDXJZQ4r6h2qal6PB0UH17o4HGLw0
/Fvy6trMVtBjLOzKy2y2QOj7UqXctBIjsJ4SCnYHwdDJA5ZNpQSPnpULF3WlMk8POqQpm4e7nEO8
ncQtMHEEmUf8rSI2jk33IlNQRFtGtur7tt/u7KTCPwSb5VDF50Ot9QMwM0VvF1joeHS4REjTrxl9
gXM6X/Zmkra1trv1E+ecWw7MVDcHDcqWt+NBakuRd4TUM5cHOgGmewwX9IhpW1z6aUrLfpieiTHE
TyP+6mbcjkf/TpHVwF0VudvbQcncmCudLfiI8wbgnJxA7K5poHJrErhunfq+xIqWqplrukJ05Hqr
xZOksTIDooypr2D2BZ7DjsAtgZQ/ZVjZ5fIeU27avqVnt0BwcIY1oBplF3ryLD+ltr5alREbv96w
DMUokcyvPcf0KDgnXu8nWSKj6fdtc+hatNpssbrRoOtZBH8yxOSogBreBgUBLWujlxKH96xSeoun
i87RquspsdvaXH4DTXCbNrwNJNA8oB7ooIozIq3RraaW6zu3z6etkvO0j8LsFQCANx0jPkeuzuU4
aAl8Ofqrn52qcVEqHEcvuIsc1xAQAUmHTCu+lArlvPw5xIfN6lz8r82csewB9j59zNesurAS1I85
SJXfEUjJWybwFWUqOIUF191zyx3xYVsjcY7WWoFSgZhKCm5vFDskFK86+4UafyPEBNaVPvQzwHSl
ksAbIkKis5xxwAA3RdQovz7lV216DWklsw/1nuvYRaUhotY42Ao8CH/moopj11aRmNuPMUV+LQ1A
nudG+1uRL6tQNIqsqLCV2rzVb/FN6YHdr2myME630I2ZUYsdQLhZoE0yIjKpaaKN3xgZhTBE0J7k
9PueAoKyF5pkCb3tIdN4VL2tsKIFAsThtQw1qoGGmARFnsP8M5gLFHmtkUA+xWw5+IHVng7XkLF4
XXElX4Nanvz82l9ltCvY1fzHv0u+awwTAHNMbud/5J89TmKjX00dqA6B75zqAqt76wYBdXWNIDXI
YQCjf3xzM9CImXorGhRexsp/HsLEZ//cir4jMfAN6jNOaNA9RA083Z1j+utDkwOxTjUHl5B1nYG/
sN+PdwZTrV8Aly7R3v82btFhUDdYJItBOefNK1YOA8Q5zIrrkqmMFFCHjbRTyiV1eQKxniYqEI3r
yIxkgqu5mPGsjdgdbJhWTkPSbIHAnxAvpmceOAN+Kmu+LBhnX8/y4kqZgwfz5BHRK1jnrZ3GFqUc
GhODyMzRiXlFZpkBhIKPgNWVQdljvgXaadD+GmPIpHIEorG734u+4Fpp8HQSelp+BLSzn20g3AoT
8Hn/QRsYJ4rBA6zOB++ApGrpZXjAS3ZhZ7y+24kniisA0Tl0NDOnrYWFvPz1M4kbTOuoT6H7AC8g
LQRlkr2nEg2cWMRJ7tPtw+3DugG3IyN2hHbaksDgKl+jRRb7yPLr63RQP+MjYlkwZ7Q5E30wD7NO
3G9xCI+DdUA3BISLsF3/DVhcVWbywjzs/ixoEN/qimXUTSb4Pfv6BaIGnJ1znb6eKnU1va+L5Y5R
u/oJjG2MCy2txIrVCNWEOmsgA2koFew7e9n8ZiO5ecwIQqt6uPAOKMmBmHY5w8czsQdEZVh4V04E
CXUvnoY6b0oMhngTn/5+YrCXTnzm7Uu+NLOenif/7zPZ8Cb2GYnD1QWLkL44X3qv3Hzvy0iIN2K+
vOarC5mEtUHaJnxWeIhD8kdEmK77DpChnkUIv0i3EvQnU9ododWZWvCkfu65/8o9UKygphaNzdNZ
B7XRHKVQDh7OfCkyxzqq0yn0dbedU/SepDWVTSPkove349mU7P3wAfh5iYSK05OXN6prKlL4+kLg
/1mZxpn0YzSf763a2fb4xpWWi17YmTWW8fXrP5J2CNKJY+bXoRbs207aCwqeoi3bH351W6V6uiO3
IHGjC2Hsmar3IBDhMPed4CBK8fv1aMrgc0VOanaZj9Ra13zMUDtHvGy9OMNm9Oeb2kyShT5icoqy
xSsnXaOog26MqeTLrA1skcrboZEgoQYlEt1KTCk29MyEoXZsVoZ5Z4crpoipX8nZ3O8/em/vstn9
ozR3rvtO1uiY7/gMfMDS2N/IQJWUYtL8C6m8TXQKjmwBk5VLT9m78JLLffSd6SEQcINB7lUzQLM+
Y6SY9Y4KCRjyayDmarPyEmYtcxJh9jlOWGBdj+c9JQP2zRb/rM8jNFRGY4vewdbJ4ftYSUXCaAN7
VIgtLqKKqt/dOohFlw9NpMAajyXiWwo/8hCArVQlrxOFx/BUWDoLkxcgE731w/JRAP7uisGQX7zL
JzLT04n+1ekx0dkuuCm+cD5OiA0NRR1mXzZLLEP16S0KHq87eq7ZmuIGAEIVVPXRAT2SUHNvOZnd
iALqMFZdJVvc8FQLj0c9JpYu5a1eazc3+5mzYTQugTT9UrV3/bUgwWzfuix9W8PvyZGW5TXmFH21
poSTnNv+9MWZI9s7V65AhYjhQvBt6yWIz5kZNYThs5ZqJVe049wLQMOekNuXjx+mmd84iSWtVV7i
O4RzZ8aC0lAi0CmGLjPsc1EZxCnk95pOi0dv5tZEhZTGG3v5C+P/84HcFMBYoZ3vW/YpHi4fGGgj
+IP4vjWTysyuXCDEZK4ZBT4/rmqfu/Yj+6C9zxEmzhxdw93nEbrmElNf/WwijQ6L9eIjlP+JkIOs
jsZwXZ1fSKyP9o7YddFNjHQOHTps3Z0fwTRA6XJI7h5khW9N4KRWv7lh+ewsfUrihtOkizXrDBHi
GP6NI9GTD6lGuJHoelymff1e9VtjbIk3BioP1Ut8LBUojiJHL1W4TQMNhOB0qYL3mrr03XizzVPy
WhMJF86uhH0xCD/JpkEBda8TpUOQQ9Hrur8+9WpOMVurNZBxfA9wct0LSMbu4blxu9uWU/1z2X5W
PiCC3KEwJDggCf82d9fbGhgTNYw6+wBFk6yTh28b7HWJhQtr99i/8hgpw9Df5yyavWisLVoQx0tD
pDGx96Y71PAsocCrsLJ2agA+8n81R/lkUgViMB9LW0MJS9cuL6I3H/UxWKLnxgd7Y5WasmsSLaYD
LQY1frinbmIz/OBCJs2p8c3XTTRdqBhujY9w+pHsVQppNETMp/zRwp11p9XvZGVh1RiLrnfoXJWt
wzVhpYTX0Q7p3vdpweXQFSv1R8pZRBT420vnbdM4/nl3cgX7w+41xNkI1kOXlLRwFBvWwisrVVCH
WVUUVeX5OwlLZOkCBiD2Gmq0aN6a7uyTJ5IsMDJcftkRvd64ZEf2/6Kn3AjdhQvI1EGlakm8T/a2
iC8Xcf3DDmVcnbyUOsTcFpGVQ1SgFuuymjXOjDlTN4ikyed60yj4Xq8dL91zevC1kMoxvEZ1CdIU
2IxgQWmgGU51hAH6tGAHAxgoTg3mpCQ/EaqWcx5psxAnKLeG5/wlL8IEGjT8SSwf6fiwzCIHZRnK
0CDFx+EaN60iZ7cKTbwhOW2GvMI6nr88X2Y175cYjp7xUrB9mwkkMIoOjuz+N6R4kx7ZRZBAU6IB
ACtEd9Nk2aq5MBpqINjEQW97VLMyuCTs4dBdI1ikx9HEleeMTglRftvtKKc6PhSGfK6puHRXcQAs
cnGwCrIKrKz8pBy40r8Mil+kFE+XMie1h2Kkr50Q7mMuZ3ogATD6QLZGuyEeNzwOUcr7Mqku9zyq
kc+raNVfCaohCpouDbSKShzZuxdYVF/DEPKRK+ASTk2BNT/c8JfsHJVrR2UahsA/P5kDkY3UOEaL
EYMQTcGIsV7DYUelVz+kWS4SS5N/bCj8x2eebU78jg9CnKQazm2tEyldI3Vl3dI0azTkt3f4MXGZ
zdtWyoM0GOQcqZnyTb3CKGF1ai5k+YBcWauB4mJXmk7Dnq9pUuRLn/0BKbtyYOBvC4nWf+y4h8NQ
PYlsmzJHS2Ax6oJ7Ksiaw2LHdePlCCaChCjfOkd9fA6EIRhSgAOdpnIzAC+Bd+sFrg68ijW86ZZa
NW1ptSKt0Cs6FHb+lXNH7TSQgLjFokLsuCrYwnYBo9M19dN4hGWqAT/RiJKNtZfCYt2o/7e8LgTj
zQMCNbgvtVSVFLOHu7AA/jxaesoDLJmbl8wtbPuvurL7mUtWxEONj7oRXE6PXjxkkQDv7ylQfP82
1+tz/WgZCNSTxIy/9YRgqaZjoZIeGBO+pX2iSuyqdlQzyQZAquQG8rZjPx3nCvcViL/9FGVoG4et
lP4r1OFB+8IrP7YetnvGbS5wxDmvo6cBOwQNMWkQpqPV3hJwHpgRohaosDXOKuRU8kXoIfkI/q/O
3oG5nsxah8BpQtd0aopMZbrPiOvUpo/vM0fb/pmgbYaZWqgO1dNyCnorfUAxj78ow/K+wQU875K1
0BW0dx153C1HXiWMqBVpenQQOLwGqJPpgdPyJgiK8LKsVnNwdze6yIFM6J4+jqtCEqYMWsB6tZbF
SahLLb+HvjSsnbzOEs88rUWRvA9IS/3dFsm1/woOCi2+h4kfZTEJBE7gp8gqdJn8nWjaTyf8xUOV
yMtKAFew6qU6Jn8xYtS8q3m2zGDIMl+vLFWJWWGadwwAn8jbHsaQtVc0Qf8Wz9saghHoUDQDCTEn
o6XRHWQoARhMM9K5Dpz/aF/dftK3eMekWazmQ7jIsSx/YB/eHdexwmNFZFt0hqIpebXCBxzKik3y
I4yjCV6crcIUqrKd/I8R3MRM/XtO9p4eMvaQZPI1gPJoZ8cL38PrhPmHxWvEEkr5MJ3VfVq4OAm0
MDeJMUNQd/0rpKBrzQyDvQV19+Nldg5jwwTX7Sar8zOxDGa9XXQO5pSzxNd4aRIThLr+rguIH08n
ExhsoNmjjY+QrToS9tXPtyfUdotSTb3JWu0aY+fc7tXi5q7M9SBA5Skh+dCFdaWTI5KXBHfg51tq
B0XtCMiVwXhuKiRPpmR6JJJRH4bRBPKE9MeTzfxYhcJ13NiVoQTeTABhW9VYjHvEJzxXLQ3BXKw0
uPwYaQcnCUpU25RDMUgcm3MA0E35Q1OVEYeJBjPxuKjRc/qPBKafvsecLpl/aJfRPfrWxp5o1lmk
6uKKy91vPC5gJAVj9VwB0GBGizFEHmUGdddUyoIEXBZaXMzZzYpgkn/7yj4cmcyGaidcgSuDqebJ
Q4YD6NvISR+VTEBL7hpJ6egBXL8Yyt5GDgNHINaB1SmIDM6XknaNzVAGe8pgCTHCh3hzC3DZuBSL
5O806Eyxf146PBuvtnwVPEu+doPb9freJXCl2i9a4NUJkHa1aWSC970WsTYu+7igWWXd16PwPage
e6pgkX6HFEGocBafkbvkGKh5T2gtLKxpWkJ/klHN2IjwtwAp9hKEUZLG30EXSJpIMqoE+IzvFSCv
6Oo01afq+POwndtzZcn/tq1tsQjMzNNuL1ez/Yxf6qsXHwcc4CnjI3JKGWfKpIU1ct95cpDgnuZa
brbmLFafGyOuVvpXeLVBol9joWb2o/m9HAWKYaFiF4CkI3kmxryUvxXwhus699nGAiiuOoaY2ojt
ekykHaCF6D+wrcm0JcqfShlXbJbct6IFxel4MuIn3Gx0SZhsY5eGIYYAm2m15KZd8swt5K4ngA/K
Qmb4Xfin/R0rluVNi5hUdCtAAaTuMiqRazWKH6cn3UIgGLd49uDB6S5R1TPczlu/wNuWtvqhoB5R
nbaKD0dUvh3W4AYL/XwCxrcBBKWfL1PPGUF3U1Tv7cXsOcC3+vklUVxOCMqDUbx/+EdkPk4QTMzj
uJ95Cwt3M28f0xUugZp3vdxZa1VKtno54O5VXvONnxptL6FiClY3xfKebjtllDfuSRkUA5s52n7Z
XQd6xRnBVGu6FVwbS7++XYdt5ifqDi73n134NUhGOewAu+0o5L8a/5TSs38pjkXLvP27wde+xvey
xfqnREK3HaXGaFKU1TproyUbzW8bhEodx8SMrXv4UxjJAlERu6BBozrL9hwa2VaETbFU53NJesLg
R2BxInOPFIj1B8rqnlGWbLPkmaRuxRWReuWeR5pHxy3FJ2UM9Colz0mSVJynvNp8z1Km6vyHk9Z3
2lAoi0FzCuMDKSXrf1/QOKxJnt3LoPzkT+IzRhlrQ6p1C4ldO364j406/UWnPWJiCUn4CDWCFCSp
RV0htafusPygylpGaxOAzos+33s64LmXFM3c9439dT6AbiieWiobCbPrhRVL4Gl0ExJ6Ku941qqG
yvI2lpnhvzEmbg/r0obDBRfqtd8eQmXCCTFucpq+tc2YalT7ZOyPpq1X+lZoMYJ726XYXTKsI7KV
WftUIhB50FFih/kprRu1rCZOI6SJ24jtqZMryInfjHaM8HltFa+eLZhSQ5s6MdXLU+N1vbScYE0x
IpRJ4kFJCsb/mPEgNEBbrpUcRzpcnYbBKt2c/VOYZY2os/SXrol+tpLkXQ2JQRrDQXMeyVlHgBJj
K4q7c6ovqtiw1DPo6uFQilWxwnWCfI8eA28qUJdxb1WfXIcKK/kqIMc2kaeGvzUUdGLnrmBI3UVL
lTvBqNXVEXBgypuzbiLdhnvhJyG0dLYd34QXZ1daVpsxkyEf4Y+cQSZm+wbI7NbgpzMmkoU5D/Rg
AozVJYzI6/c+5x7UI0VkpFRAZEokEqFOuva5+3N66EFvXreAeFyK+uoem6b+KBClHzuSQUpAHofk
pbmvnZ+WkP3wtqeNPr84KDgdkHLfTvqxrB6ol35M8I6XBT4UUHuRQbMZy0C8c5I4NEOVf935Kdfp
PFG3T/kGRPpMEumnRDSMEk27gujIRJNRAZ3dN/m8PgWve0uvoDmcL0JzQ+xHwQae7dNriq+9nd6d
WOeutLkIwU2C9d3E2tuKupsGDNoYJsVdMxaApJMS/Fl0fGSSpe7MtYmSeXRQFAO5/9btP2Ldd3jM
v2tOVVH3Ccmp9QKtS7lxaOt1U6Ufu8eI0QZ92BAPNlk83NhxrHxDNP2OJ8UIN6vn6yTGN+fnJk1L
92CHamrYIxznHm7hwaTkXK2oBNoshGwyOABzgAUHp/bM06i6V7/jqDgNVoTYkw+NZTJGxPQNm19y
UQoGKEHPTV++RcyS25mwp5s6UVZ2bmc3bWZ9GhSsRjcy824X9alpNjljCXq2BYW5bRQYwAa5itwh
1h6L2k0c1PEVYUh+3zvYV7eMDVbNkDwCEO7bVHbYDptO8kWzvIxj/omU5qoNPfnGVmD/54t/RvIZ
y4PrEQ6dWLD4VrI46gs6iIW+5HGMawJJCy2Kd1OvqFpDvIB29Owf8XTc6N9rdgNGRklNehwSRikh
/Ut2mGyheODk6Imn31lY+ioVZ78M7Ajl9hc/1aL/xtjwMZZNyjAfqjMijMO/EjQPpTvpsSGAsTQu
Bm2phREKPTdGgFTGZ6z1yOD2Ko1d6Qpp+1y2DrjsTiY7eTSRG9VDSXBGVXfgEp+gQvR1xoPAaGI8
anEn76hMLGE2zhkSdcR+aBog9b/AUR+mJLUPXn+iEGdSR/ZQywRIAsyavYw9StUgYuns0oSATY96
tnlTknVYS2giijPc3IehwgXiTf4X2HeNJRpHQyUyU/UZ4arLBuiUooVtkqpH/KvuYfShVB5LCnPo
/63DOfu5iFpZ5oDi9JKL5gUP5OsFlf9dsjKGgHdLUr3l7RT66xbxrcsU8CiMJDYEBm2uCgW0SvXV
bbrWq3tLM5opB9hGciGf7KO0t+izR0nBVw6p7KaPmlf4EK85lWj3wLtaD4mIB1Z5EAIBl9MONFLJ
frP+LHxdY8Zbr5GUzuxm6VQpCdpmISKMgO25XDSGwXujbkdoj9Y0axZERcATIUkWouD1m4nSkqRx
Fwsg7S7581Oow1x9bqhUoG/jZoz5CL3DkNguR+EytQaM7uSCRxdKnpRAx3GkKEWwIvMhlDoreFSq
6dT6vitPhXctpAXEplpLW/yw6CVem9ITcU8TcX7l6JAgSfogFVktfdUUqtdBaSLXAs2IExLdFSFY
xQelx3m2TOsufWdJ/IuNzpz3Cy0J/70e0cINnHmLBqNR+U3ZlBXfoHqDhzxXN9XTQMRX7mURwwvG
dw909ovG44YdtltVUeGwYm0JhNYuHy66RVJc7p2XDOz0XQyUrnCm10AvnzdajazpKHuiMeV2oG/z
x4wrD65SZ5KOvvRw3w5E0N2mknBNJujtJvN6867GG0SwTTcRsEKqQdkYRX1fSOY4lv6AB93U4qdN
aaaZ2uJlhbjx378zap4p1Fbf1uPVJDWbR6seIsO19qbJMqJApY3olPEwlNkAnPRihErNV9XTDa6K
PsfAOJO6NcO3+q5SUMZWZHjDFYRS23coyKzqn3r9uCt+cGLFA0iyd8vbwhDMFF+8KAaMiIOKgH2C
Ceh4b3NEEHFhmga1A15WQ/3vgc7/P8/SdjYykolDou/k8vNBF/EwrCQOMgXaSiwCjA6X4lMQjN/v
XPEb47elnNN4muZpq+e/r3aCLFtTA3CQ9cBrc7CwqVENcRcOAB7NJxUMzb2LMuL7fSafHkTCmt7h
5mo6GqpFfaMK9mRYKQx+5QEBJkIkU2OuMrl9yzIFEsgx23FMQbo5paa/23lK/RraoeS08r/nyOP7
QlAKHf0+Hc2hioHobIftdDR+Ru3J4EceK9DAaR+jMkgSJWN8OGFG0KDaetJ83mSI5EGa5H79Dgxu
rsbik5VIbVHXHyDrhhTwvf1R45437ipYK9eAQ4lsIuVbcTJ/CPm0j3Z8ZrRLld79uH8KyJqY/XVr
ZsKWW7famTJxV4Bm90GUMyyT+gzjSLrKDthi5Ls1gokz+fwVvrD4gXy1KWaITFeX1FpNw1G86aN7
qULBAgd5geR0FaQ6nu/ZBdpfJAR057vkavkw3g+YZuuuXUvkvrlSy46KKdsRhlBoWXK2IPWlOKwG
17UgLE+hznP6NjTpqMovOxUwm8pkoh9JCpUzAZ/1XQafjWfLUmYE9ys3+fRyHT5zTVy+BInHNaYY
jouSIt8dIsHzBtEVF0nbBgE/Z8BJpxP+sQ2kUPvahzMSQsTBz+WToDlz2ijrKwbt5/9K5y/N8PTY
1J4epH5Yhw8M+CsTrgNFnumYLuYKutIHeYViikl8v2a6n5OhPrt4vMI0RscwYkuQETSBBTLpzGl4
TlByfYcz+UXtCaXQmOHn7KNnTdKWjeeclX71D8Fvs/tCU9sxNJAUIcjuYGKzAbU3SDsm2OhxdzSt
78us199ard8xy8PUiuSa66EZwDT2CvicLgnes4vPKuvhx+sIGC4ZEWyjyDpDh+UdrQUBGWbsRAUW
g4XaDLthDs/lwVR9c0R182Hc+GuF4Ba8Tn4TFmrEFsY4Xi3PnT7CjOfgzeVF8GC8jYmZPVy8dLar
g8wDZ9QIb+npDuddiDYOw/6a4IG2Fn26XGOhkQGbwKBDJ8w47+6GgJ4o76WbqJMbeablLQ9WBPpT
KN4Yf8cMAyL1wpmW7XZc1J9R1Y5Wz5hQcB3/uZ7JTENS1niXZrYDHZZO9rePH+X1cKE+h5E/JfNM
1f+lALbktMR38HFlrDWzpE4FmL2ASUtpvy9fQ73JQOxBnhhLbTgIVgUWS+i6ypSy6ctfT8A3BVV5
2jcUTA60S+QJbVGsBdiOnQuW2aYy/OlYYNJvNvFRqEGDYSUX/kHyIv+EGSYiXxW3RtMXl0cDfGEK
R50ffrEY1pOTKVmBBMyhZFogHAmCMDN0Z3bTOjHWCqqBgDtlxCQGCapmqYKnZGAzAIhFLoV3schR
37Q4POHC1CXNKwbXB/NapftNp2iiVLTA0lRxcNN9fQSPJsFwAMVUqLT7o/q/2AElmLYHueAEtGQk
fHi9+moFGvpmPmmBEA9QGmVsm1ZjF0wpQpGhlrmJcWSvgu8buUkQsloUH9kMRa3f0Mjv2143tUUr
k5ZwkseQqNpuyzvs3kNYAXlW/WclzciKWGYRGw+cRq0srapImf//odsYTcXjSqxYUxhB5Nb57Rz3
NN79x3eqL5UtB+BAPni1Hm66+sDF5KMJANeLHvDADdFAhAv1+v0mZ5SV3ZS9Y03wdslt+5mvpFWp
95LtfvYnm05k0LJQE3sBpGviVtpW2yoRKOb9ocOWNWQr2qEW8cEUCVcgt8swyOBz5h5dsL2+5EQq
MTMJH6ZF9LqptvqppweEy4bAPj1Et0gR2guG+tqpeZXuioOCY8i4Vbl1nLl7S3scCIbGCtB7eg7W
9JPqwhdJyhQ02jYnnD2gb7bllAlwm8m7m54odOVjE8VJpbTc5sAz/WxZlFBe8jeHqiQYQvbsWHVu
vetCev7DfgqNNV/EW4BDZ3wzQX8Q66KkkpEtf4tPgiylggQ0MUYhTiP9VRoXBPQa6Czcid+WaqkL
wiP3DQhHdSOvKwOq5e774ULtjOWgf8TOQXfSjx2iwFOgo/kjtJQ7fuwnoqQoujYWRyOKI21I2wpq
ycpLE9JZ9A93ubu5DIGNrcop3dmVhhKuoITEsGs5fTfM+1OFAca7WgNcDDj5cBtm+ZOzj7a9Yv5Y
JoXPD8D+b9v1C6vu+Ye+YZecChdwtw9jwKOK7hqjIxcG1TTavjI9qGU1IDKuB03fX3W4+3GTkx0O
hDYt6xzZHZyla7V8Yofoa4mkrK7mO2ilwVezysXRSm9BM+dnn582A6ADJZyOoSmWN0JUKGOCuTob
hlWTIUSrJpXur0jLdVr+CGOxN5ejjHc+6BQffmnsboM6HAkjxspCFjWoERMnsTbr48z+trLzl0Ty
M/McLoSumfQ7y/8IURKGHk4umLmu22P+6NbCcoOU28JrNQ1KDdghgAg97TQXAIw1TAD7k5nXdl14
wQwhUHTGKJoKDBTRGreBEHm+z1P85S9XGjoI7SSw6WKSc8CJvqJxW5qnQLtsLTDSNb6EtvET6BSK
dZe4EHJShFB48xtv1woPDFJhK2pJXGchMGZw7Wjvj7h4OrgdF3t3u8GFu3XQTEJSWnUbKGyIjVQ4
6yQc3+YUq8wQKbT6b/mB2F8WNyhwPfy/8e3ZVVsUykREREVIgn/Ml++BCKjfTWbDTauoDxZThs/P
r1VBxlwoxRZVMoVqL9wYu+QzK6yrtMh1SehmvGWr6t2mOWb7soIt/BSPnQ8vt9XIq5JHmJhBFgpn
Vz+sZ7iIDMBmCWlvl5jclbj9Cg1qpeAlUHPUTE/3o8ampGl2bNSar4HxqJrd7+gYbE52dxlF1kF/
xbUnsMV0/fcae2S7UfnipT+jCnfizZJgn80QU/ywhoAGTzEraQMnrJKCXgDyjSI04JtNrZ3r6mRX
6sYHig/Shany5YvH+WgM/BIMiCnls6L2e8dGY8blBSV37lbDTfRmAMqbk9mY6/6m0A+lxAfqFOJx
iV59dRJfbohsMiyOJyuurmkQPKUfYXE2kZJioymWNvn5HFVHqFM+VQZP9zXEdtfaDU6AwNv0NtMH
DEY04aRum1xvfO+ozruhjyevLZ/pB2aWOkSBFjckS/g1nYyZMpw5Y45Wok3ZngRWKQfHOFdoES1M
Ox/n1RLdIo0P5aqI3gLjS+k/SzDLJD9b0v5i36bYKyOkNh2vkEdHaL3khnzq9a/RaneZpd52o+bj
fqbRGe8ez5k1hCshPCdo6Upd4upoRQWAkBR8/aoAMb4YgvKZXtjiGYbkYomVH+vv84+PkEMzkSwH
IxTD0TXM3FupXNgH+TgdUPkqQlcagK7BB9V7IgYRSi+Y5R7hZRRNzrDAjcyQ+9P4KYWW+movilNx
XZ1SmF17py5Asj06iv66BwxZNnv3TqoHefqKXe715WFtVQHXjIEEW2xLH/5jrr72LhQcbhWk3wYb
OwM9Y88JsUpPyk3ftKQrueUEAC73Znwr7x5TvxNyz3RtaEG3wK5O/ybm6iicY9YXs6HHipR8jxTe
Kdj3Gsa/t15V72LO0vLqFssL4cd4riA+TabShK1eCSDTbxzqPIY0YfbHncjA3b7wY8TJME1qTg21
KZuwAlewbTW0xEe/D7shCZn+bd078gO13TztFKBL7l6u53gEz85ENi6kmVBeL3cLuE6RHp3vOeiQ
lur4JVsqYZlIeWHBNrTDh7aDE6iZsIceJZ/9OzPFkc9l+qdJ3LnuJWnM3Yi3kbJnF5xv8DezZSaq
K96u7DT8e+c3P3SZdvMZuk1vv+3AN3xtDeYEjNzPt0ON74HJ67ENtb/kphyHHHzXwXuH6uwn9pqj
jF6kMLvd030MkB9gOdfVVHeeBrSVfzxMboa16My6i+8o8dC0Cnok4LlznbF/eqzQyrjc0oTAvR/U
o/DYoPmNFwsxAl9JHaV5WnhO/WMwbiJiy7lqhRxGzVsq5ixw+Dzh/zt6DekfSj64+W+3HbwzhzL0
D5axBnrIe/T4mjRlWEszNVl7ufipfVKMA0rVgOBvu5EHF3zYKIz5CyMzAzwxDZJ4Z/+pTXIXUYiL
nHYEQl0sKy60w8juMti51ps1AYjtm/89GJRysJYi4x3eNvuCEQArxYiq8pMe/ViyFtKRidUY38MY
Ns5v0qvk5HYGO1SSNvh6hA28XivJSNtE6v0iD/J/XiXTIqqXBuvBOO3YWdIUYWs49gQ0du3Vy86b
g+tGme7/+jgDidmNe/rDwtOb8t96Ya+AAgDKqynmI7zeCMS0keuCkqPL9CpMXvWdsvN8wPm3tRrf
3gLCzCtXGK7bZfiaHhEBrT4niqPQnrp9/x6S+3JgBD8lR49udU6dUhV/CM7fzz6ap4sfH3MXaDUD
iDrFjZ2Vwj4iRM/0cLA5IHXDXX24LkuU7oC0O9tpJlSVe/MbjHuKw8Gl+j4lIcSge4NyrCAll+O2
RgN3lXRQiFqGU6SJUa3Ru8GscFe0k30feLtfLVv0IKlgW1ZXvcSBWO49mKQMyyC4Y6fljWaoBfwr
V8jDKfrQLRSgdvGHFyLI/VXyCj8F01cFXzRjpzUwzkDGCc2N/T33UazOwvq3bxBLlF/Exvom+ZVx
7s0HH5jIq863T6q3mfxdvcWe5zT09IIZkXhdxnVHKCHpJB6l2hrXVmtF2yzEaEqMtIYWAdwzpic+
+cNa4ctp/UfOAKkmBbAu2s1Jlw720CTCz7tRMAdH2aBtNc2U/EwnBuXgUqXmecYosGMFyUx8uY0e
uyjqnjw6jTZKNWpBYobgFridk9ZLGH0B4Szqzj027UJ2NQfC6bNwj9o1sWBdt1fyFMONcb1tfvXD
Xbm1SRc1IJK6mV9EXCRINSmvz5eEo/0lYvQ9ccvcaSj3LOsEofHddwXTd1rjpvgdn16QIJ9+UBjE
VqG74BfKvVnQccwYMfKimCYXY3DZ1taChbtOINiY8XGBlS9THSWO8arAW2ac6wrqXV1SMi68/R61
D71P6AEuWTER7LykxVNiuaC0JaGM8SmxBA4mUs/O6CxNJhbU9sShGKLVov6b/HYWvKTEu0zx4Cfg
FkDPOhQtgU9Ujs3dMbOgdBjXQ/iOQ1Dz4OXDJlLpTZez3CeYEZ1k3Wg9rulbBWHWf9HjXqRIncxO
l2uE+y14bS2FbTqLel3ITKFhumBEoH46dz8v3Hf0sec+VEC+9/wNwJPXJN70Fz4kJLvmuiFxYQf/
L7dfeGqSLdJd87mrRDARHk0ayjCfyD6Ezu/ntvt0hX5d1R/jLccvFAoBl7iMAGJHDOPQmUAuj3hW
Z2GPZ9KWdSz2wKNq8+ixu8XETMYQCs2qr0HExLozxpEMMJ0CDfXVsHxYn+Wgc5ReK+efOVTa8Wh9
Pc2ScNPZy1fIsB+HFA3BNbu+oa6ZnAKKRREkEHI4CCYqLXWTBzhMbDhzkBT7z76kbw7inZp12SNK
Qpq7pcu2UOfA/X9dR3Kkeyf65aaAblqFV7ycIHiJT/JaynHW6LNZ48xAHYzMUFFgefga8TtlQ50k
eJ7So0svJJjj/SMc4Ezu7j1Bg5JgrPJwO4JLbaZ7/xdgrw7qIu6iSAMr190X+3isfdEgYuzwu44r
w1+z2F59AR3pgX/WZL6nC8dRXfKUZ8I/550WgXLsEeAByDrpq1sZ0LLLh84Uxb/Uog/1F2pNDPri
2C0sS4h4jKzanIgOPZO4FnKWMqWnP5I2LsxPtx4e9Qs5rhp4FBmocXXcPYnylgQ8zWOZ8AOXX6Jv
Tnrv32x38k29S/qbnMqTKrPGm+7uZZEzXTAnZEwuRptnMxAhanW9rxXCOGWW/t9uOwZwoGSk5w99
2Otpt0cLKyORpccBoX1DB3o3e5e/fvtlVuHf80mxyPctJOETG1bnecI1z+z9NdVWVvJ9abgTRqSN
sJ0nqpw1oJrAKH0uX43EfEe76CxU1df3e6CqZNR1avm2G0uccuFy/EABdjE3Vvwtodu01TnET6ep
vrKpSqs6q3Lqjvr8vPH4pMYjFnn4WOGxldbJO87+fjcdVpCkaPtDTiGfkIS8mEJbwJudzpPGywNM
xCagHK42ZPQEMAhvZPCtkNPw9dCbcoWwodz1C3iZs3Ws6Lzg1J3A3htFlbBAlZaxWgOrzCFqhvPF
m8rdi6npoUhuc2ZkF4L2kD2N5j6FfisiPPf/15AxHLyJ1lJcCJ1TO4cUCoaMdZlaxbdH8FWqWeln
W2Q6hP3OIf/v99JqdK1r8Pk/KCchUPels3RAapZTNnZVT6gu1SvE5dEtIPigupgLN46wahGBrGKN
0eCQmt//RDGVFK0sQuM7ESOCRUpqU8qU+uWCA+CIyieXAudRiUXvYy9O59yyfxdVcq/Ih1KUyZsX
zWg2ylSaV8ZVyc/hh7qgrOWjX5rYPLqckRnnBz7lkmnDQdMneEA5Ugvgi4i+rdw8h+t946kHcRUL
fjO/wSSGJanEmIsoeR/MS7DW6Aq1FNsqnFptMtnQxTdqoYPqPBgoQBZHHk3MbUjhH8NI2wxj9GYL
6ug/S0VEsA+BkrWWHXMK0q2MYIiggE+EHUv6JTPCR2zH9BaroML+Qyc4cIeNdjGsjrzr62WQlLCg
gwyOszKE0WBy0mIGMwMG20kwEf+bEbV5B9E6MegTryCJjije/70p1YBzbCA0ZxxrRt4O/HCZbYmp
pj/TYnLnBPV7L3ILi13K8wBazBjcXwQib9XtmzFgdQDwGGWywsx6HwaqfFDxJO2EEk6+0zw+fY2x
SmEdmvRSI5EHuTSGrvgQ9sFFU2+zXCLNubMs6OzUP7j4B6ssoJaSjDb2L6ZY6TnqIcKemeP0M2K0
2GQcrBK94QvgBYEwcj6mh4e+Lw5OmuyEq3bQhb+4cl0zQdMlN9jD9lLLJ/gEKLv6yJ3THWZslWl8
WetV1xvIET3kWkMsFkRrE4GbDNu3wmoh5K+MartB6SOhDK+oUDOrmg2Gw7iPnjvwqUtUCY25OyYR
GSoitl9MjY6jgtpo+TxEwAa/jjkC5EzkAcc3nVUJbu8Zqp2coQ22pW1svMoFUz+JhNe3QZQZonvt
tQT8F3yA2eVcA277M7OtUKEmP+C/VcWliHrCTaYyZB4VVrCMaas5M1/6Atdvh/OiKW6NY8aeA+GY
yn0P6XY3QLgrWelEOAgqBUZv02wwo96sgTHeGQ2wpZKwedyO2MVKvJNTJvpUKQGz0yx4V8PMLYE3
kd3EE8tkfz/gwiWii8ZNVqWc5FgPVUeUgBQW12/fk/xZQEJlwb4mxt7atrFW4snaTkBofyBrC5rT
SYhw8OjbtdO6xRzrb3jbSEcArfLN2Sx55ZfVuN3T4UVTaxjv58SxKq1otK7oMVNq7oUqpYIhWCdn
xViRWsutFpf46Swt47lszSa1Xu7aZIANZTL8XXMe/2uCEqmJY8NPMBQYJOQNon5VjdHcTd1IBnVZ
wo2dwJHT5cswL8iXDiCeRN3F1LMT1KYO2CkW2oLEIXS17mQ0Mk/ViZuaV2NKywhx8eEC0+lc4uzU
T01xc09cOFP3jIVZkW40lz2P31aGMfAiwGUF2rnpYqvqE5VcFoMo20gab5iKmutonPBqtb3p14UC
ncIcsepwrrXoeAb4hScqUpc1HCnIMRj8EaqvXW+Rxim/aXtsJEqeHVHtBbw8XgnayS7SmuB/XjOu
RChc8mJCXNrOtqT7VJGST7JyRq9feEnaTUcPow9a/Wp4STX2JDQsVgCXykRRyM7SWbjBJ07Nurg0
X/QJCqF4ZU5YVQ4HEIrm9AYI3eHkcFNowoT8JkjwIfs5/TISVcH3ylM4MjYugnfgSTqqN/VsV9ln
beZJeY9AhGyzOhPRT6fmZ+Xyx7Oxn5xXampPsHmgjflnUIzYW8P1ivIcY+TBkSSJiTzjdv/+3xHx
lnnStfT9d0xr8TEPbGV2sNFJmrM7aAkgJhMmNiVd6llUVqVmw0eM/q1RTXGywCePIZk5T0IEv1y7
ORRg4MN7M1I0YGJcyuDfE2Q1eqSIJJLhQIWNT/OGys3kf2ontdyJ0+zTkd/a2r/rWUpwnBcpUgMT
MCidi4NPkxF7kWKvk57Q/c5PSJbXW8kLKPko4TaExZrDPGgiQPVtkZKRdeDpXPt4qo1iCEegd4Fy
8IIOmtjIBwa/vrtEwDp5Bgn03KKh5PKlXc7q+U1yq6Q0lsfr6l69vfCZQgZektrXi6DGRTth8pe7
T/ddCGIBrQprZVmPI1WGoCnbZqRRz7Vx/dyu3tucTtTkVOGdjKgGABi/2xtqDqvZVSLcsaSaoabS
QsSG943b516KhZCaaoFanDqOXp+Uz5S21P9aU/R8yTvckOXIM5DjwNa4f9KCk5R/qe+LFdsnm1zI
/xVgKyQ24shQvIWbd2PQF8M3J/Gn9JtfRnMxvmJ/gR82iRYvx1xP8i+tXxdvIkTz8HdsavXUv//i
/cIt7Vfg4upRZFSY+HjW86niBhB6N6mzFylWBtQu1+RQrewMFaWDClX5pICbDm3aim+rPAsSsskf
EBeJtK01VsSMKMtdnFIhWJEr03xqzwqQJ3CCVob/jb0qaxfpwx7nb/fyFPe7K0ThPiJEe3v1Gm/j
KZV4NRewG05M9Llb4mUL0nUoKT84yuoL48XAFCRi5w6p9K+GHjdHdfesaooyCJ43CyhTeQK89XZf
sv+FmbnSgfUM2F5/N5c6/IuoTnK36XFTnKMfIF5YdPhk8L8zor2E4w5XDSy8iwd2RlhI1UMn7bRg
WRhK/kB6EYSYDKlm04DR30c6h1at6q6sW3hllRF/Dh2Q36Qz9Xue6495jZ7do9jTnwsv8jHoJCq8
prZSHe//QGk+HHgE2H3iDuOugczWd6zOWIeuMYPGXLTUnO6tkCh/sO4jNPq8N2I2GBvWWo1cjkfS
reZ21XGP34da4jS4mAzsHUQ40EIN7gk9leFcjsS+zW+d7eUsvbl7RvdYoIYMkzJzbnpqF3Ho31cE
rZ93ZDmA0CXamrIwuEzXSPOTQSlc3rUetqfqiNhFLHRlMbS0OrGLaQbzSpxFUtTk8ys+u/Tv1AQ3
q5MRhw1thTab8LRc76DheMhyga6L6aKj6P6Q06OaTz8OOGTDdMV7OqqR48tKI1dvS2mEyn9sewFq
r5QmHJOeWQCN4MdaGscC4JC5GHMVcDaI2Ws3qpu7hXEudXW+s9ByVcO1eYzXvody4aOwfM2hdBI0
zy17hweqKRNavuu2ODgVLNGhMXNNL5MeMDsG5TVLMyWsVIci7Uxqq4hHcXPvPmjVTJT4WZqtWue+
SRvyTXExWZErGUu6iaK9TL/mBBYHLjauaCWsHUjffy7kurwddYOk65FbUjelX4GorZsnnklCD1gG
E4N7dynPtQajzUf33u4hWDI9WJssaLGptvrOdL1U61bbSHUrMn0fzmmHI7ujI/CZxHzSxq0yk+eu
A/Q1JUJF+7Q7/jJ0dv5v1aZQ/A4jIjc5Z/keRTJDgUtT5VMDIAi0NNTHotQlLQwwWXTka0YGZ4nh
bqKaLogLDk9xNDMc5STwxZuJ3VbqRuSeQxzUFTDMu89kzoqSBzH25LaP3FTKBpEWk8yap1M/pjsa
jvQvw9HRik9i4R8luMTJe4xfyq+Sq359lRKxRgJOvg59nOW5SDJBs6SQXwlfrQPOH1ZCrTo/43P0
3kNTTOR6edTb57l6a9JB2sSKsIEzlkMk5gQadE8IFB66gnOe6vOwBQmqEnrAACC1joAAfcXi7iti
o8CI4VXcuZoWyqcTsMGqwfeuER0Yc6tXAuoi9c0qlcYDhIvzIRIM5YCxjGQytcbqZ5K0PKFTYLXd
TQ6NwUfVfDZ3yCWgLUcQca09tccMyXD7W+CJ4qNfTokZD5rCPU7Y2jVtkcNjU2PPilvHultcLEmF
O8O947zbQ2DrX15PjvHrHt8KPSYPGpKcoNAy98ECQwAcXPblxBHTKWAi50vG8T+yIEgUH/yWf0CA
MhbAZ8EQC+DdirrJxFW1qdZQJ7nK+C6XwKiuGnH0YpUvWuoMjytezat3Wv4qjwiPqQSfddtOm7g4
EIxY4/s9l9J6am47FuPrcKOi8D50R40dfc+dyU1NZhc/pcPtY6KQwkBpImUqpGEudlwD8ulj8n9l
FfMXS3WT0xx38WNrI0AubYO6iuF9rbZN/PcThItwwyfNlRA/dI63D0XZvZg6sYSPUXC7x+J4rbtz
Cr43lTW1APpG9ZHQJgfjq8GfuvUh8w3atfI47MlKWmmBvrI5WU9dJ352vHbrxgj+/TX72mAbzHlZ
J8usYGAowgj1TT5fUR7NTYqJeYssBHEtqGbfdShux3gziqL3xz96xnYklzs09EiVGEtDbYrXcdKX
F+JAKPvbf4ZPSSKbwSBWvAuPZp6Tlch3v0TKCMQm30te8r/91U5mYy8pGTJ9ynECp2hgpDt4Ikyd
fJV8IOQWp0gd6MAfHVNzoS4wvOMiBZ+ZITcXN084jzSNnQb+sTAKC++kbDrEUt1DPrXCsIkd4jJc
U+tXLb4eL3wRULvJlpWLDp/t5Fwmz+10GXrR7U712yUXOfFb3s8Jm6q1I2S5Q82QQhOfITL3Gxmv
I2jLt6+M0ghbVArXL5XhK2+7lo/nXmDI1A2agBGkKYwJ59s6eFpRWIyD5L6SPw+OV+yz7hnmUaEV
2+RimSBikAeP7k89Wu++y+JBCKD4x+RU9YdM57tEHK13kS7r1FtdEL7vLoFaDU6RfBAzQrr34NdL
TP0g6MeEgb+OrrzMfjU1FetcKJl+9lPo+SrNSnb1QaN1Frlh0HHX1/SlAWdw+Dgk9hAT//jLZkcs
W2Y1uCCCZ2MLz/PvpQAG7h2XCcoma1BD/GoEVEpGLP9ctLjmHoVWAKnWyRgKgMaqhip0xjb1+L8g
eD3804KgEyVkwezEEhcceoTb6e4GP6Zq6y+dqCLVlDbNfccxZci/v7rXbF6TZ2rpWNIPCtFikYoq
FAqtd1VKzTPLNDj7mrrWbZbVIHf5zlWMKiwHSDvr4ZtUJm2I7tov8oAyYIjUvMUKyFlDY8iJYPu3
qAQPoQ6mNnrsM4WmmYkkmBnSae/dgSsLqJ/s6SKNoZ7eq+cmlsE7ZONxVVyNZgO4V7SqrBMaYTTG
IrPAD8vR39w5jG3UkyCfHCYTuvv9kAJZU1+xxhZFzvNBLbWxJMS15F5zWd0b4nN1yolt8QdGXs34
Hpndslu5dBy+1U5OrOUroRUtONUo2FGtWVSF/5JhBAuRLOa7bV643fSSwGV9t01zM3rP6Aze7sGB
gilgNYg11dXTAgKl66LD8721cJAiQNg0PFTI8mVBycu9pUU/YS7yHFJrVoTSWBU17Psc5JpOfjcH
VMSDKe0jMXdUsyROCU+ZM3DHGHI7usK6MIgsXF00IFt7aJGGZb0RPdxMvHXZUY0PJGP/49n+wuYn
yu0hdzPtoYiKAUVWAACALQ7+bXJRpUVaXiupNrA31iDO2NF96MzkX2jDxmInNhSBM9VUiatKg/gd
IL+Z2HeQptNoIGsNmSmgK/LCklIDd7Wqkk6yfldFNo5eEg4bldZdbjCz1d1cPZpWLRTm3eRW4nnG
3C1/jZN6ywEHw9wfNqIZfBwiMwgMYAgH7sZPNQaRSZaJ8AIKfbRrz0j5C3g2BkncBHHQYiPc7dlz
KLhCdiwht+wK5xepTPPIO3ujI862J+N5HTA7zs78D488CcXIQ+pXR331i2Pst1B/gKNx0qkicbXM
6PKpVCb4Q0pLgeXHhWl99A4rWmwCJq5T5guLH2y2dtzon9zBSpQteLwq8E6JHU/zcie4JoY7wjjM
oIZlKQ7pfq4uqKb2f6UZUM64U4BU/c6TdVJPW8SmZn1MBmE6xqOyvccLAVNbxaSd0gyNz/w7+1mm
r0HjAIxXjOVHEjIxZYEmcZwERbc1UqOSdAeIlXwhjlXGggg8HuhWCqYf1KsqZMu/yQUyj6MbdjO4
yNiCFq6GJOdTFkEXnBHjojqkOROzQBAtn+GpCDzt1/d1Z2mBFTSLF/lzjRvHNj2eGGsUQ7bS/tzW
b809cSC+XPZCWeh297oAQa5/Zl00DNsJDvLS34zmPqw60aKQUWO7xrpxam2jbVvCVQcklFkOBHT/
/uA0evVnqphgchAVluYfewz3KvLKcpDqqw8PEckNc3wJCQz8awKZSZVNX0R/PM/larlFIJO26fb0
U/ntJt5N0gndSSUccH+azwVOGYYXIk4gnjg5PWOXb5ix07QnCOOvnHHT5MWPzI74lSFhUT1QFVYE
jofexQ8RuuhQBpjmOFzUemEMdHe6/WujWQppCXXyzSs/m54e7CMkC/uX9rvt86YIzNEhHpn4x+SL
f84DM0hDep2MPr3IdOg/QUpVkAldv2l8IQMqo59RLgTUzXYIU754uNrO8jltrGEs7A2q0recGNhl
gkMjTNvpTdRPkIyNcrV9q77UQPBf2pEM7Z6Z5SxRVvTVaNA5k/aO5zP5fFKkM3CstjZPYc3yenM9
Ex0IegLH/8MmRMBIQdphTvzGS9rzWqYRgIaabR52Uli/hxBoKwnSUswzXJdnnjpreEjJqSMZcpv8
gCgb1MpLF45w8OrOgLlkib+k5h3+98rhqH/gHaVNUEJfIgg7K+4WJucm+ei2zSXQlA4DM7kuNMwp
d6Mx3axnKJlnWvTLxn95yqXx1z7zQ1r9brLi9rrOgZdKRZApc7j8xqIo2CtfruqSWWjs/X8s5mTc
8QnHGbWra9Rz9Vr7WAQxl2nD/oRt335hjod/hJxMkf+FPRrI4mBdVnA2lpc86bJ+tKVubox9ixo8
3cIDaBDC33ZU4VfJZHw0nIg+aQUjyIqu3D+lmP5Ea54+L72mP5/oFAPehVyojq5Wu/IwXJJNRKnm
Ds7sizkkxvg9FZR2XezYmyk00lz8vJg/p7Leky8h9l5iHTppAgE68kxdPO7jzJIdGeTln0yuUQiM
/wsbQnMTsZeSBm4sAD8O/NQgso3+3ah/BMuVlcDyKMAPi+cS8OG7zoF7+qlEummi0UHUrZ9TdCmp
HKFG9+iZZq0XYlkRrgYF1L1D1MihhKV3kdeI8JS5WDHspGczOC9/DSciS42n0jJ4X3XBv0N9HqW3
gqZtaZR3mO49+/F7thGDKScR0HlQYjuIXGAiaZzwHXtgUJmqFK3Zsh+b1dFYuyHv+WcUrw4iSGqh
kpL31zfEX8mnJKJdXmlqPPC3ur24jJNKq9do/tVOyyZpboy8IHCxpSc+I02EJ4TBAMIqkl1Qvo4K
xEJ8M7ZBdntJfpGgml0Br7KHXdMaAY2ybY8xxwa8lJFLu1aM+O/52sc4zejlc3GLLNvxiIdym5ua
Hda4ezM2ywN5tJ5FI0k+X4qUj0l/V2Pkxz4swPovgEQkSa8QKNaQXS4MQd/OvfB5VJUvfIaChAp7
0HCTjbnT7ItygXugcWdGDBk2aTSwm79BBD9xtRu5bdOfN1pyd6sxa/Nr+xIVsgX0x85Oa5aeuRQU
mWIFCYsHXhTh2sZHd0uJ3KXhtnFrpiWNsOO+TJ1YuzC8DeiItAUQqTbfTiyXYs3Q3oCuNVLYAV2c
VMAZ43pYepPGp4s/hSCzyqHGTldc9cRc4nlRYIoqw2dAVpMNn0gua/fU6HlPcptfQRDGlfB9rC2s
xpbjcbIaePn238UH/ZdnEX4jxYQVXRrE+u16oLwMyH0V9u/l6Qxpkrp84YCujCe6J+bWZWbyWxKY
xMIcaJpm0Epe6NYbiNIJrvYdTQvBoKnk4YMUfCvlN0nmv8X+ZAmU76KGkyLT2CWZ4KuhO2LHuIdf
pRMvAgGc1ud8KPdHoPk04TuddIim1z7Wt3Cn1/JdnmaOfnB2IcJ6LZxfqXS2GZ+giIJSNEwB0uTg
Yqfo+hEewLU7Q5WRXKrLktxCnGXRajwIoaRpA5LpNzPbC83XTEu3DMTIfKN7DS12i3xuftPGXCTC
9yHJJu4DMIvKqIo2W7nU3YMv4kqTM6hp2UdCtb6R7r2PBmb23XbKqIBnSmApSHQ6XcITS3hC3LT8
AXKoe9pgNsUMgI8kyMowUTZZ9WREI/b8ddA6JykAd9oF21I96NtjzokJ3LQ1Iwqh2HSDHHvbBo+v
KVw09Cg4tvHtsC8Z68caF3Dc70wFpY3nYBp7Ynin2aqZBSdS+p9VDa1sEMCOzpre80Rk7yUQhpWi
G985KeXkU3ChbX7FIPOvZMXoOlL+t+tlfMCqfaGipI8BEB/xRLM/FNHCNJzi3RNoYGZZd+q3kiNh
UKV6XUSnBXzHS1oWwFgPJ5uQ6XtQ/YUqy1gnEWfx2f6LafFgborXLqvWsLzia5YyzO3VQZfJ7HYu
6wEU7GIEoZZVpMxN+kkFy0U2HWarYbMWIi+Zi2xXvAsaUp+pmTOcbo7fDymVVcAocMc/p5QeHRS4
h0lcAkKjDQWW2ce0SBuKfRwNYoRLqoqd42BGzKoruAgA2dewDonAcusyVrDYG2Go0bIC7o5Hj5Gg
kHnwr6S6Rt6F3tN40QZMFyNXk3Z5qjcylr9Z9rpBieG1tVoqNkGKxawBZOXnTpSv6tK1GXp2/fs4
nMZZzBbpLZkLh6TmRXMeIIx4kgR2iCZAslSAPsWjxa88Zro5zZychi1wzSA4ms4AHxZusI+VqnMm
kmsdCogRzoHw1i0YKOPvMevP3PWPFaGkkTya5XohxIgpCyfSLWm39ltICj+L77Zlo1VzvItNfO6t
BG3vIU2l1MHD2wlHdELPEpwmsCm4b76EZrZMKIpXV4zIBZG8d/BSM30xJWfP3cydpw9Fkx7dbcBA
8tgYsq1Zzvgk/KNPRbcKhoofPaX7FU2x7OlFa6T2rSZWtz9AwLh/JaMdJnQDN2rSo+NmmlhifhG3
QGK8joYLZ4GKU2XClgK4D40tm0z+gtCf2NwSYskZjVksDbYW4XAyI+EH2p3iBI3V5aac/VRoYQ4l
dopOzDrvbzlDJAcAPU/tClfVWwht14IxNqdMLl7oxr8Nj6e4QotxpuZBuQIp9ynBrr4ZdHKsGLLY
Z3OuisT1vWlG1NmgyslwcYc7VXFN6IrXgwiKek3bGJZv2YPTVegbYYlwRQVACTBlizTQWROj0p5y
usRiL8By5rbli1FkLaB+WfWxKdmK4+Imu/B2NMfe+81rgzDZKdXtduyVgf28W7+9iyTxpBpwDadH
LgIhxFL42L0A+OkxqulXlxLoxqumMAVbvgALHyWiLwqlKej2GJvfJlICLlM317k3H11rwDJJmlMo
UpaEQ6cDRVINO3B55mMx3UYU+rZYcmOO6MVclnqxJIO5pQYOoZG4FWrZNDj0Ej0KBGtvJTdsOK5f
XI0vAbqCzPn+4w7DcbFh3rqb+ouzTKmjYEYoXjP/aMekk2cPDuZIl694ozMJO94tx8nJgfKmlnnT
MJ0A+WMingR7GBcxJeRpVfF3dn4gL2v3oueo9bBVSZrqYlJvOk0FcpW0iCFHq/K9cjEK45i69bEn
1dn6zx0mKE4tRR/D9OHf2/a4SOS5Gyt9zB9+M0xFrFlxrvTSwrDjvifR/swFqnyJWw7NBp1qN6FM
VCQtmgsIx4hXfdUk9w8yKJLxrhiMSMUFECdhcAl7Jm+9Kj9aGb/4FwxkdPMojHoU2hTsIT8cj3iQ
EmzMrrZlQKdLKuolcFNbQPfcgHMIKFak5gwDEaRg/Q/ZTIWDIo87GKYk9JGVa/Fs6P6unkUx9pLD
ZbCJI6dPCgrzskKneBn9tZYwxRv1A/nav4j+GXvfNYpnaqHHW5C6ZITz0PGX1qpra1RGIe60n17D
HHzuNHfns7YhAO5hXcBdDfv8RBtvAi7FcmqAGMYAGy79+UhgNMvekKs7h8yeWSx8rq5mh5OcEKqx
0+/u5FJxVPMBhj/BVzbvWKAo9lAlJIMhCLmmwwvBGiDswpXg1E6iJcIBGYuTzW9/JD/8e0sSQXzd
yqiiLJw36Ly1t3q5hXXFz3ecXZzQF6+uEmJAf1nPsOjBwSWP1MkgXQqxeNrstcNtYLzPsKjHpgYE
fb8hBDKA20ugxAKGoE2s9yz0HmEFrthdCnDnd/WXtcT/ArYJ3kkIvmRLJIWqpjjOFUCK3Rkp3d6m
jGgGaU5aLMl+RjP2gWsTfDRNCcxi+gbqKuyDPZthH+eWeQvYA/Z6h9qu7HG4funhnvD7MRyepN1c
NJVeDvH7xw6EBV6gMu0NKKIqFDa9wDW3dRl09NOvXbPkOiPmb8Qg+Y0ExzEsHxBVZgBw3Ph1EJ37
U6atYZgfRW8LvrSG/A3LtBrYpjtPO80KH0MwCjN1QMRW9sNtKSNujhjB5cDg201a20pjPLLhEu9b
B877gjYImnpEA0UpNITESxkWLBKLPmRbw4grnmf19trmiHn6QqNTbMXjBFB4g7axFMwfYR2gn2br
m6plBXSWTF2Dy2DHtAsW8fUWv5hjzzeXM7TJfijAGtf3guBWneKOJs1kLn2Z5Dt+9Ygi0+R+oVQE
0Jkfgxqm4TEYe4pgl4g7q22jshTKhZtceYH6g8SQPly4d6wVACC9Kf6GRbRRMQQogGsrnInGRQZp
NL1p4/Nl7pUCObSNjYuo8YnwVXbzp9OhWNcetv2VmuAvHZzPmKCyqR/eaaTjdoVAoaUE4j+HvKPH
IKZmT9Rg59/sSruB7ZX8HshGKMDn/ElIcClJYjldivW+gbExSjE2xOs0pR1uLVe5rCTDqWMbFobf
p7KxKyZihybeqrdRN6EEL5D22Jtbl991M9BJjg8oqn31hJqV16cSgBdVHAITiq+w+EWv74kqB5Ut
/yCS/c2pHOSVj9OibJtW2xqvgRpiE1eMGnpipDjQrivqf8DJFg7yN9KX/46wqxR3LSQHmsjShY6b
2nnh69Eby993CE8jI9HHkiApiZWaT68bvE5z2+Dk4Zgr3SNwZOhJ5PZqyBbjK0wfw3SQdPetrkZe
iCoG5n0HY6szSYd3sHxv1G0pWeNvo6QLzmSuBt3gfPUCFOApGJnTCdxNjJKI2kLabNFaBblzT4so
7Uq5HjIb0kLMI7qLo8b/QLB9JWpbF3dDOf4QdVzbJ1uUczjBXxp+gVJKFtLtQ2oZJ+w719UoJYqp
Qxv42KihtXDwveDuAg79X+kOF8aKd76EuzfgkW+eoBTgCYCzXGIhVyas5KsC0pdffqTQN2hsfLkv
/0ED6r2iDc8MJYhsBkYUJOlcb2UUHdnYDEAk++odIJkdvXt1AhkdixoIFydcgWBd1RcP27oFy/UV
jTuY1SIv9APBUnkgAjq3fIB13Hwn9+Xc20Ep6PNy2AX/WVaqzafo7vy+RKr7g9RYht9gYNx/weY3
Wy34VjE7HsAkQ+SxjmVTSwnxGFjIJA98RPyD9hkszndwBmZQQ4vwLiTE3CR9vpXN6ccS2sIAXJcw
Uw5PpapXnZCMvSWdqVpyxxZhLOx7bxIalJq3WW5+yOnZRFIX4cYpxH3UsgTSWa3Mr/IxfrISX1QU
edyOxSwpLDXE1NStgZ8PHn+2OKjQ0iZQp3y3VcJSnQJViJST43UK804tDY9+prlp38JW7kREcv+d
l6zPOVVlpPZ7RnZe5dqJ3Nss6o6Z29IXcizkqNBo6H1bfU6EdJeb4HFELn67Nhg46EtbBWbYGyPS
ddRJKsx3Ws3c5AeRrDCgunBK64v+5ORvCxtirEwL2MCk+ljFz0ycQu4MerFvMy0JroO3kIAwGG4U
fwd/O9qMCTZtfAwyYeXTY4eMzlqYbB8LiylqXeQUykTS5zGiDNeh10nvjrCuFMstAZ3JNQnjHTdM
yQXYgGI9pz454kf0RmHcxG4dVShDikY7XfboyRl98DydOyRXuBhUhSV71Zl+HpZhSy6/IxSGUtMr
Hzpr+4A3N9jq0onA7nOUh6+125rLX7BHxgcbWcn7mry/3ZnnUoBYABaJegX34lz55rgtbW4HFd7N
6XBlEnTRCyG13zmfPzUUKxgBTaJJlLpTO+EQRBWzwFn4qahX4bPgsnRBgeWJ/bdmOj/SjngJiDhm
T6VNo8OkKHRxU2E8kpOmD/Q4pUGZdxJGzZqKy52SE7NFWVjFxspcY5G0S/dGOu9XLsPTj0t0IA2j
VE5aMvylqEYVMeNF0J814AtCcY9Ehw8dmwVDnOBCDWXvzn4SMGY/LF4r+YrDdRfdxSWwqYxxLc58
KOW91eSUJgkvvErL963TrzhWAaUSe5WSRVXaOvuopAsRiApG8j43QyguYWgo0mOSwkU8/nPJCU4B
a8vN0P+7dL1htuJmrVUwzMFzgaUsebGkuWDGzO5a9kVMkv/zquCFLe7T6nDXB5p+fcopWfiHS3DR
6DPKfOA+nP1mWdb0e3zYXDTAyHwNF4pDLPXFpKPgbg3VDZ86TV2T/zvG2w0u6PlBdG99CXomBpKF
pOMFoH41hNYOh2xGHAH4AECSS4Mv8eJgDokpKuKAynSzdnve7wpGkA7DBf2ndByAgDdrQkypdMWl
P/REnlTAlW6fZe/xZI1P2u8ByFKHyVLJBnwiJOcIDtgFaxz6/nIvtjOl8RA99ft1VDDbib+HgB3c
tLZyfncBZvIv1bEHGJSSrnsw3dHwK5CgzUwaSg0H473fFnpHGWZ5BrrwsRgZi4Kt4f0M5HVNcMcJ
jGrEANWLDj4byPqaTRE8JY6gRl0puChrX8e4omybLaYf2xN462zIkRrq9TVQzc3gMn6xbaV5B1nl
w6qJFN01Y5YnSaxgemmaABU0/vNE8LDNsy1w9I1+s8rgDcb8yLNzPEQjXeVy9cj+GCbhi4uB1pXk
rgB032XUl4tgg2Nl0s6Ksytq4gt1lH+rZPjCYVLQ70olrTjGGH2WqHZN/wQ9kvRc4eqt9slDJY+z
mxbkIi1SiaMYxrXeRVikrYg91t93db1V9WO4mf/73t61GR2VRzqVh9Xg8qcr81ohMm0wYpMZJQKD
T8zgNtQa9zPGEB6/9rgnx7iU8vaH8pcXju5Xoz58wqnJ+9bDGfycrmTz8kkflgYMtDw8ITKqzzrp
7dltO3CwWSwzz+je5kmQ4pv67gEd/+NL7aH9+sFAt/HSiWK2yjA1uqVzdtg65G43gGjN7kRs6/Dx
0ObsbZvkok1ghDACI0Vq/ZJy16S9mHyVuBbpjawNp5gOv/0NNTiIYmr0XqoIGWduiJ79UjT4bsIJ
AQV3Y3+mb1JXy9Hvw2aH6719zdHHjHc7olpVyLhb6y37KYmrKtmmP6TmsFsulV0e6r0U3rEbAN24
keHbrYQijGyODE5lmIe7bUvoJv+P4i95TkfEtsBKKFRQr2/gHCQnVtXTz8dIbYERGcHlfhZgvlQ2
RpukCFHPZbbnFMAAKO5d8nHN4hChiRnymnsuQCFILqnl6UcuHYcRXr5P0aBvHHDdnvDgUrx+6O72
Q/ZIiQWVwdN4DNFKqEEF8TEfSPx96hCJk5mA80FivA2dO/+Ij/WlCjZPqqBNW2NqsHrTb/AznT+p
RDGqiLmnRx4Nqu/tr8T+mwV7YfdvyDlzK6jFOKnt4aSYSaeYt+50wULJz3s9hOHY86Usamdf3CSZ
KhHiAuMbGxB0e+cJSYJ/qFv/aZq5+PPrU19oD2KNoxg61m7tGQ7Jw/WzPeDK47ro1pe/S9dkC1dJ
o0VPKDe97GC1x9v3zewlTT8jF3IdAbpsAi9+/4eo1YH+X5YmcF0EloyFAQQWgo4OAIzHpnb6oiEO
V7tqD2/GjFMi1PAbZvrCxkEuR5B4V+MY+1WFJsYAnUWEznLsp+K8WKiok5+HPKMs75UPZTf6n224
3hCsndyWyde+WDiBSbNwSZ/Ax1nU1z8jrWsICUtaCBYJ30qpPeNbadTfR3Kmt1OoLuXqEZkJN68A
wNlG5SdJbB1/jSbdQbJLp74mkODzFrVcJkLhRu4wX/Ib+vtzui9KkhZcLxHa7xeCHEMD9Cpl+jsL
bFZAMTxz9mtn7zArYs3aucl7YQrgvXImKOb/MmltkzbietySsARYmoalpB1HVZ+MSJvZLoGIVjDt
e34K7y2Yg4HOGyMRo08U8m4KNeEkcU7C9IXNLicU/dtpinfcgQ2+l6XxJMMSQJehuMrSQlspJFDS
3osFkDyYiygi4oys34LVi/Il1adUIEahmR5mAr0/uPWDuAWodyeauyy345iyVM0PGQpZjjHiMn1a
nMglZD+Zo5b3qqE8IW9bG9KbYMyiloGn/1RjZlV0+tADUPJXujE2mK+x1dmKUZdnLumjSjZKOC7o
fHwOe6QxW2huJtsPh/1JE4daObnRJ3MtZYzLtHB9T/7KQSsqNhEeGK99YVqzt8zly0sT+Fnm5zmU
1y/oeEywf0T01sn1+O+AH9SeYwkAdn9fRedub4yVor1vL4u/SHd9M6Ih7C3+TA8YFSDLVf8d7UfZ
5oq8b11msF4iYfOhFDBUVRQrChm4Qnwr3FFES3CSkdkHDSmh8G7tP5JW7uVE4qUoh2nEnhWpG09Y
iE3rl6J9o43v8PDXkjW496JP9KNQpzNxqF/zWHs6XcTergkOrSAS4C/OubaKC1G2miTnMV4OWCi/
Adf66r3j4N3kDahZFq4cVqUg15MudcKUOWxQHl2kwaPfRIBo2LKeZsnYLGCf7PViYyQcQa1inF8X
O4y1KAnuNF4Ml7CrNDO6S5LI3dgKUYf7wOcgPHe3Bz+gge8/Qbws32I44kMdo4OCEOG+xLKVcKnk
qTjt1jXSH4uoY0VGH5L/2W+ygEBYFPMWX8UXsuVwPSTb1emQD4N7RUVr4Mdqv+fgCJR694JPWF39
PQFqOKXDzhX2aI04Ru1ULXb9FVbgvXOiNjzBGll3JDd8UHD4QYunfpUJESN55vDBMJJcLmCffpEj
eFZ4EX5heKqCjveSPywEaJwJ/nX5PnD9geY2k7jJT7PvsZdNwt0ZKr7xHv/hHYcUNy4HCStGtlX+
8u6kd6nZ8f/BBXINkJ840HlWK063DZeAM1VCdFqYWmR23fRf4vPAMX9cDCY3WlHPSIX8Rchqoy5h
lk2cdLdAmI3t7r91Z5gymKRBuZIyKQfJjtbmCiVVFoJWbbvLS9rzyE88FaFJ8+3FGGWVwJzUi6cJ
GhnAl/A69XkASP09ju1BJaUL1xT08yAngOsSonYsmamSZ2b7LUv+IPHsJbDf6qUbS5MbYjWzvcI3
s2Ur4k+/E0ExNW6J00zHeCNBK+UvRzLkbYLoa/Y1e2fzo07rDdXzOmdm4rETHEBWvgUbpcHH73y/
lowKHclKs6eTuP7ZxkwmjQRuUGymGw9uQq10ZXZGIWeUajAXsbCi9WN+oUuM9OtQBn/7uxpg482p
PJL5zJhjhmtQPql2A/Gfh8wYbYLbCgmToq5KcYGrf1swyE6Ur9y6GL8eRdKhlR/eHDIeRDC9itWF
rwzJOLuUdqTWpTayL7Vp7ZeXO3sYw0njQuu/GMOYhkQc4eLn9/UuWrl36aGB+CDjahYO1HAiFHKS
wsdyDrGzX7rdQVwwVqLEPbGVn/gZgchdbvzHOUrFrMGYMIgZV1pYfRtY1rogKSFbMNBVVZweyi8V
00V3kJnlz+DCRMuZ+HtA2IfzPNDujkf0dlNh35Tccr8jJgclfJM0Ug10wLv18oQAMItWrXx772Ss
Aq4ElZPfG3PwHiemfNgW2a6gnJrYa1iyoVH6EAnGKcDlccYwk18d00btpHTqPM2sujzTlperdnuu
vCidQpKGSyPTkQY+dr8X4fZ6NrpVtV/7eFa6XqLoxfxjbRveMprtX84paNh7+sc7cTGHseZ15fAb
wA+xSKVYofcSfAEnlzyv588mWK4Pr7kaaGjM+CTcIojEY8y9ECeZ67HeIfb1wqCO6BiybjOuQiox
CDJ0XN8SuDGXN+kGk6qr6kVHfDzUdULhOwfOb5mLtFfuZlfpMlW4cpsryqZMmBrlzC9VC2COKbvz
Dw7DZvVEEt3t44LbIi9EuYQwxVBl3kVe/5qZaa4ADKsCGoGjaL+4OIV6SMLB5ZkokRizkyuJUKNs
rrlBMOOY6XViAqyVcYZ0LqXhPWt9QnMqLQAsJyO78xikHhsHGMzdtEVbwswofj/oqIn5lYR1CO7v
XBJMnG8fYMQMqlUWJrdt01HQYX6jEA3fU3obgxV8GoPnCRFDzZYVrNpG4+k92lpLhxl5K6eP8Y63
WeGQcpE8E0ymFJ1vTIK2ALfrsoc3XTZkwHMpVL3//HzT52dzZuxWZqLpgrMW8zTMA4PotTNl8vLG
MyLanjfl7CIv19eeWWQF748YS5V5+0P3gkA46n6AKDsexf+EH1Fa64roE+pTvCOv2ieQQ1hOekJ4
0DPdB+6o3tSPTCdCgTdXh/i5qSNyyZDgLVyuVGoWRmZjajJa2WmYBQCFDyS9PhFR86jtp61plHEH
rF2sBgqyPQfdunMZYXFWm2yxBe0A1sHSjxDuSIYm3nRGvW0rBIL4psj8jDhagBarfnjz+03VWd1o
T1AHgPIRjnIEqpwmvdgJ3STd0gJ2KDz8yFhOGeRfnvwMiQaUZ+mQPxMi7PKHmwVD3atpjHtt7OjZ
RNwe/YegYEcTAzpPhipivi10JGfwbv4fIu2j0KjQW+ZmUU+Usofz8vmU2t9ik7pub+evriREtZrT
FpRwuhKVVUHu6weiQ7j6P2X15z2LFwzKiJHysA7km511vFzs7rCfCCjJk28MV8fj1UvjTXlt0dKf
uK7ZTfCLSAM7NOUdFrBRF4gITdtLv4iATre1oTqrJooEOwGOla7lg1vVEJ5u8yP4UkUuXwcOY1kO
DS/OAeUDR38mFN/64PMfaW5uxUg4JbTSfsRSGoBPsvGDyXy1OzuA3336HfpO0oSMtFdDRDS19k6C
21pEr2Ftni+6B4pI5HjdAMmZOykfWGgmr9fSIiXuPip+W7Prsu60mP8V22hbktHpyncbS5OqGlUd
/QiA7gw9ZnfQGlG1i/4E/YoaGDvktc7fn0qPCRwNB2SxFARQfer3tllGYgOV/RUrCx/81AsiHSfB
ghrmrMDRDAA8Hw5JWnQkpA37zd2y5zsk/3mORdRLrjOfwiGCI/6uP4sosWkWCXJ8ytcg/+vzXHlN
tIErF7k1kwwFt+EQWpkugKZ4npkTjxwLZuINaXDhzn2tPbg5r5vrLKHwFYho1Yg9bW1d/LLBa6lc
hQy8+ZqnHJSTmh29wIG0a2JefXJukqafZ4XgznwXvXaXQId/jGWL4DnV6Kydd+d25WsSwv9f3iy+
Pj3Bj/8jIFq94kFOs7Z6hPKfUCFhC8ur1ljRZwURfx+vzTHM3r77Z3jiz0D/frtmxMd3Z/DMqCHX
tmcL4TQI/MzNFmcu6IXHMwFb5l3xc6IrGeDwZ6hYSFsSnfJZWcRYkwVzuDu2lfCD8Cw+WyktGr+o
CgqqEg/h+Psd6W1wa3TMtQ3jGD827Wx3KlrPQSX+LDVgxS2DY5tN0QDPDCs5WdtUxsre0pXYaFZM
ZFPDLdmeFAwedHXD28BTkoz4vRS5HAeZKNBG7lZjLStT2wGHKyLdfwVlnn87UYQN1dTSHggC0MK9
3XgE4FkE8w1XJCyjvE/eb7OowVyHiqVixCOyy6QiFBtkUHMCAkP6vSjGT8sXe4tXDn/m//F3udkJ
bDl04RZJzuufRQaE2Igr8Ydpi+70KJzyiXFI5eU7dYaYiljZuz5jH2tVq/4iBa5Q2WPmsADtkZcS
OJfLf68dsHOeP/tTFaysmELHLIDtATIUhita0UMAuWlNGP2HsHlBErKcjIJ7uh9WYhoycpDyIyeN
mhis3Bal3yo3AfYlm/87jCOE4Awn9mN5+IxpZdaZX9TfvaGOJGsmV8VG7CehIAfozVvKfPte0KaU
19GfivUE/BwijW4SjkheV2yLbqBqrkWwQB1jIPWMywQW5z7TvvIrrqBNksP2d9G3A+UbRbqeGhPT
3tigHA9bfCPhRsHvTOlJ8eoV7+GH3LWkFaPi1wVVuLoOe1+0eTTqVB3vZla33TDbi1Qb23wfGx09
TIf+EW0etcR29OHSdWJ60SjYy7AbCShP0AhNtXAD/o0PpGwi23QbTx9Lgds3BRbpsDLWfVZafiia
4qzT7C/JO+Yam6Td5FiGQWT51j6OBJQ80I5zZ/Y3VkM3XG4z5waQ1aWt9RgjSKLwjr5It+BBXA6a
JBQ9Ioc7IYxLOxrqT7bgG1hsERqAU7Ijzij4ALG2ojxjQ1jf3iiLiAJXKKlHbnX0/6NEnZyyfGSz
P7BphgJJvWg9U2vp5emHq6VF7cpYBav7aqp2WP8T3BlFe6gdbcHyozzm1+WNqLe4ZY9nWu3JJeFV
Ws5MGRhtwUe5bWfzeClhyTrKDmEIvFqImaR9CfQgLwiTRALhI65I/LkX2KLrRr1wu6/FILlXzUzG
z/4jLHQR2PzAQv0a5424Bhrs4MG6DYkjKwKksjEhM07s7b5ZWBZhkpyCJGDjFGMOQKXRwWujElL2
EhV0sSQ1nqFa6yg/LZd4RrXXXZn0TWu0OWePxXsCyAfv4DbuDB9gdM6IEx1avm5TYrFH4M9ePcGZ
iatG38Ka1patu9IDVOL08CWWohqVpwdNDOmlekhC5zW0YzB+POXw6ZfOdsmQjg08t370yHVEbLhm
lPGOLKb6h9kteqNTHmpKhgkwYkd5kZl5u6pe6gOmKR5zf9O+7mRZGAwA6BLMPVrBGEfobD97Ggyu
qiYtECsg7bG6eyVzI0KrRqLxoASRI/vOb/wnbRvo9XV1dwzw4BCnAPWfTbXDOIOGX8D2LxOEbwBI
Ye1N7chz+6ZWncJrQyaclzZ25E7rk8qx4Onflz97RAoyQyqlx6pGBqstzpL8P29lv3WVidwSzF7o
+ZWJCYuGXtMS/FA8HgCbViqw6daNphAqWXTEm9fmbAi++WJ1N2Npeb6FxGnF+BzDwu2tdaxLkqTS
RO6NQvaSqNOoI6isnkszac/ZsG4JgjG+ztt8vCVU4mQPHEbIXDw1+Tc/0KBmalnvAuE0Ri0yELgi
LPRQqX+BCM1Zc5GUeYUwy9SyIi0YdYFnAI2hDmqoXOHKubdO58olPZQ/9UWUszr22N0y0bi9U0P6
3Q637+d3LUdkIGv/2wY7amutPi9j78lGn2xLC82+m1JoDoon+lZqIi+JhgddNn032Wwhpbgsg9kj
kFHRNG1zQWqkZXuradIMRA/Vab6pxyB2pNJHZlxdGDz/XpE+QLtZMvwiywsOnXOQnd+cmDKl+B9v
deQNA9r61ZPUHJqoKrjKHl0nCBgVSBbLdirx0zFUnNRAcCPndU4too5UWrCjo7aeCeG6CGEbof4M
B/TpOW71ewgLVq2m4E1bMYbnA16dN7wUM3KdRcHknIchmP6eSpbSQ4VBTVBnScykP+TPUpNYof7Z
ImCwpVwoeHiAspmM6wBvJ30hsOiAuS8L14+MYGFkB/ZHesghz381LFWsqir4GVspxeRFvieGq3w+
fj0Zd1/ApptCgvZwjoz+Ki70KGVieCeblG7lr6SBujtSnoldi3QLicKTtx2vI8SJv5uEgqdrt2Mg
CmYhB9HnBj4r1KZUdZQXkboDzeMXDI7WNyx4pVkuYnrJRY2fRkGBACWNn97offgwMBhY/c7YzGuV
SLA3QqU8wUA+bBAmDCm2y7CngOVcGi9vGjgHEEivQbrTNilNepTj/ZEeEJnb5rtpZexIE6RvX5Tk
bJgD1PEWcdv3PZoELY5C2oQTPwVtvYyrdJ3ZfPfUf+4+xIxCdM3eOvT1oClpxmQJToUBKsL2XZ8r
qK7miH9nCQU+d8aa82dk6Yqwf2rnGS6SIBjFQiFIYfJhHcMrfp3k4uuTEicqTScGZGIvOYq7hXwv
owQd5L+PV5UQ86477zQBeylVtJB7C02YfjZPaQOO19PBsIrnbf3xHNhOjjedISPBvwARocN1vu74
YLiskbEiavuPzt6xXoEwiTOOS7CNHJ8wZV5hFsPEMs5JwD3Gls9QxvTUC+Jjq8WhxU5ol40G3SpM
i0K+vPQR2J+f3AAAub+Vk/1eAOIy0cmzdOpZhJh6wyAJnAvcXaxk69Ke2M5gd8iMy3JaWcn7UDv4
fNiVp3BrGSxxywi8CpbpqrwEJb6URR2qs8QS8LKj2Fcu64hozxznlvs9f6wxSbpgvUXAemoIvt/k
SokT8CeNMgipsZNfOfpgSsbJvvpAmyXPyMzB0syVIYKwQInopkaMSHFl8wOlFU9h75qHMwBNviXr
XbgRED+5WCD3/tsLBJXgfBb+285USIycfsyTEmRRGwTnZNbWWEvj0dSscOhvqmQ9h/i41T+mlTsc
jFhq1KeeZBhe5BtbNXcAVIm4TrneW6MXeSYP9G3JlGmjfVJt6o30Rkc07mbNGnR3i5N2+nyHYam4
/ZIijmOwJATJ574K/mWJt9CR2niqf/zu8O6vQVB1ivYv8Ijv7KlgKC234tXHtMXjMPHrFOFzpvtq
RYGLtPJ/tFLz4lvhAChcp6djHhpYbOq+QtE/fg/EQjyIVCLRPkQwtGv8pZNOI5cRRsfYKaKVa+/E
2MhNm98MLKlDvmjct0aFKw0T/YJWrAyX/Kl51hgfrVId3oXr2Nvzjy5dN3fEGGJfBa53rhAoCfgK
Dx+QMTHFbFIt4ZtQH12cO3KfzCPOnitVPlIFHPElrWfaUJxCYzgoZ1QSCeRDeqluCe30X2mZdGuZ
VRZ+FkXRC1FTmlQj4E676JKWFxdaGl8KZzr9w6y+uhHZ1zb8EtuVcrxNSdYmMZc2+F3BWQRQwyHz
wvT0JeKgxab6NgBkkt3ZUvFMMhMDcw8XzbEoHp28w/PeHVSWtxyWOXQkgr2PbVmweL4P133br9ef
FdF22dDP8FWsoc/3h0ljLnrJcQJpO9XTW3ludqIN04YiEk56buSDsLD2zTYE1vB4jtupUJOEgtjX
d5M3SFXEQUWV6LqHtnz33Z0KVh1GlNTtIBC+LWvqaniuXZytRicEzcZ3szzhg0nX6iIo+GnTTdS/
eiy6GZ4uAZiiDWxXnKMdChIjShySqf/wPfdlCULNOl/pOg9S0fdo49hTrSmgRdqSZJdUU3NSAkH5
eqXlqzCiJOdxyKo4iboxVgDV9YHo2Cj5y639RdLle5V+d2HiFvsdRLTWLfnZ6rmXf1O5GrWeHZFv
X7R6XS3eDF7DeczjsCw7yunYPwL2Q5XvTrkbSnW96rAwltiWMfsGxv38Q3LzmveSAE17auztZzkY
KQegVC/pzNDaW3OHQ5vrle6fR2h+xlF8Q6HFoUNzdUGdOiMxuY+bRAbdQafRKPw85+BqBTs3hCl7
jGBPu+MpogFpQIcmNkJ0UaNuzVM+DY3ZzdURAkFMw2w6VYnhOuZNCiNb45VrWXhGri+FqTBoequX
P5neCrf2JDDQd7L/RW0gcEAC3KE5xbUm54Z8RoNNVyEidI8r9JkOjuTv31MhdTrIUBKht7HmMc0p
lQKu0miUTP2Bkzw7fSFPBefiWGo4cEpo3kRz/8PWvv5K1mIbRWWEHm+rGYuLsYb55H787FtJqDM4
W9wKAd0bzDH1Pxk3cJuSgxtktw94riIsU+MT1Y27WIhPX1ISQ3gXzuf7peYzFhJ/SDoyFPdmvlXZ
oRFWWPOrgaASiakuJmpnBHgnp2M79fD2O2iHgUv4qJq//X78Z1gibwCh1iZakPR6YTXA2F6lZpaV
VwkK4YZ75a9Gg/X+g/49XAuKUuncBogu8z4zqDoVHaL+JF42kIFadjcNn4EmRYjdnw2Ma1l3yjDL
1oJ72rGwzTy9MCIpkOrrvMZ8pB4SfTu7gemNqXEgWWyz0vd7LjjdB+1Ir5XVkAuiaU9CQDnyUweh
qwWlLKHKjilaP3qDQqIKjlOsETOfaH8WJ96Vaefs7DSoecyBBkCHlizS5/riuDH591TaxfPCKV+C
h9GUszl8xaL81dLx2dmb74HffN9nei+V9AxS3RDa4PX7Tndievw5G/I9XWD/JCOwTOx3SCD8Qqxe
ogin5lETYWgWJtKqp0owxDbhjQcDqLWuzMDF5/VolV1g+c680WN5U3zEnveT1+qe8uXdUAY3zhu0
2363P/BphPeRYo2F2yB7qNSGmzpoVrnxl/OIV89rf961ifQEyTOczZlkahJMYZTB9cxljs1802OJ
BYatr2pm04dX/vE6L5Yz6C2QjSYkbj5xV3474VyaymfWftxkb6eg3ew1oF8viQ3Rp1NOSxcjejWr
gYwZM/3KK0oxC7YnwrH147k+29BYXpMc8Bb1ayASAYH7Bo/BL+D36afm6rJDnxTrJg0hsu5giZtS
R4Kbqp5J8ZLJaxfXjhevmVFrwWYt995G0s7Qw+Q3UsRPDDO1kJYX+mmmAtCxIXqau1ApGA0evbaA
DOolwx1+0n6cWXl3uB4Lx3g60ZBu1uwfSLyaHFYUnNImf3K/zritXMRICxnzP+BVSj7ElEpU9IX4
Ap7bZiqTViIOsMZ0JB3fcbILMEmn8BGfh7CWL0nKrxj7ZrG7wf5mBeEBXh56ay5CUFn9jq3aq/3J
vMixYzoYyjwmNFD5bQOf/bRZ2bCW33UPHIEp6MnfrB2RiHyPuchVQ+/IaVbzZkGpt2Qy313+LAXV
sWyp67wStW+MNb4pY+P6sNp9MtjkXNaxYEaiG7rIQU2FTpHNiiHouTmA+Ubu8wiVWTWPTs0l0Odm
C8+wlK7Yut4ZVwdkYqhMFJgvKLvkvRrj1j+qr9IIeP1lz55sd12mzIjBDPxc+48/I5wB8s5hlXTZ
xF577Ki48OWqxO0qls0v8WcwO1TVyyKtBuugfLQWNCNJiYsm1pkuFh/Io367SHC5pBseRxpLgXs4
SDMB11kxNxJyorMS9BaYNCp2IfpYsec860iI/3xV4EXXtQ7IgWZxtzQazQXTyA6rrtV0m/Vur0bs
yf6Omo57LQYVFSwvGXuTOcE28JQqf9vGgrZibhF+YCZ6sh5capUBuFr+O2obHG6mR4YaH7jmYWvQ
IOQme6bPyP/RWRbvHkajwpHoAo/MwEW9X2nshTD2BeoakI3E+A20fKurzp4+3OVFDyEMfsQicZoA
FgQppEM9UvHS3R3pmX6FwlfdMxZf78tTYwPXtWg+lHvkJuGcvR+YE3M7z5lqKXsD7pDgAKe1eXkv
zMXXaYP/uBhCSC9bqeLrpt2XNMi0tyQOLp0AOB/3yW4uM8hJVJxvZ5dJRqMjfiXRj+8DnQzFjJwd
lFQVN8ewKDL9w0F6dW6hQD+85T09ThPDMD0h3Ww6DDfS58H1i9L5R3Skx+doGeJs1XM7A2E1k2DP
tnjEoVUnT1CCBYC56H++nqulRlvvQw3qru0nts9E+kQSmTNyeVFXlVBU8aJ7oMCtVe8Q+Qw9v5aW
Qu0/e49tQe5TSriKqmAGmOQyd4XQu7wdFwD001uZsmDxbiWzYSqFUCcbZSD+dOMeKDdJi4QEFUVV
9YqWotmpEOJq1QPEtK8UZCOFOF3j3Xnt721kFlEY0N36hqzeu1zucVGz3OKeZLTOSzwJGz9a/aed
9TCd2X0LqL6tycQsULiI+5VlD7ck3Lw5SXSml3MAbOXql//KQZOJRRe6JUZWoZfFAyEi8SEuIwCB
SstTTL6D8z3ZYkYs8C7nu9Pz8h1/B+NYtL01MMaqskWJsHuzE7r/qdneDY7ZmmZsEHRUafh2047C
tG3dKQQcYp05OAZ/2O9XM8fxx+6BqQHIfINVU5GkxjMZGDG0EJL9YzWLJdPhxsW25UT1644G54KD
zE58bSrlXYN7Qmt+Xz7vobZPzPBJj4RO2/mo5F1rqKmkEgvRblQduSkw+lArSKODXs0xy0satZ7q
P0vE1D7mA6pxYKET1m8M78YuSvKTlKKrzoVgqVrlD8tUo+gvJWjKsLn95e7QXVNWqxn2qzhOqkcJ
DoPr1h4oQ8uA6ogujdAZRtfuMpmdt9T8FCIJNfUHcdIrgtS0BY0+PJK7hq81sMX3AhyDBOgNzs5O
VEg4jiy1QEUxv0OeFCtEyHibHm2L9qTkP2ce1IXiD+4NsuGCF8QyRQOJ1swMdT8ZvRuk1OluK/jg
tCEeGZwTDDG50NKztO6ZECBsamP4DcUKWQncf8Bj1t0X0hd2sSEEgtUOiduq5OgpvODQrguHYruk
KfZVPdGmpb7074yLAv2ojilxUtD2kX/4PKFtu6ialezsDuwet/Tg3QFJbATVlXybYl4IQtm35Wmf
bTcphtho/jpYkd093SmkkzWMT+El0bbAb01Fd4mrUbhjXrCgq7Mts8itohrxabq6lhrt/qJWlRtS
751z1hpqr5+dKR338/a/Ykxwy1XxwbdyicRLtwsoj71ekn3EMOivEpPZjNi1AXratyir0BK3Y+SG
YEz88w8t90NHEv5YnYPgm1c5fU2ehFTqGSOq6CtAU2RZ8VlH5fmBqLUkXCiVB8VjIm1k8Tf5pcQL
gzeGBhSpep7wLp0fAa37HAhxBY3zBk/kb0Jk8/L0OqW3erS+8qpv+SvNpRR5r1O4ZaAqrZfdHEj8
DXHQuw1L/4K5S+NNCSxWVEL5LIc4opPJz9AFAF3zxD4i5YVsrOLNuV8/P+NXu8vxYfzZIbf4W7CH
0EXpsGi4+uu6uUCWWM0Kr/wACAN4kQ8B8JTHo4VHq01N6b0dlFErzc8A5eQnQu6R2la1ZP0jR1jF
aVWSezD0CHJ21AhJ0fExkTxbTnvkZIkcF1XrHnEE3hFcerGPmCj1w+sGq6eP8BkauDGDNruIdlFZ
zhS7zmBftFfgc3I2sussmZeawbvomCTK/au8yLMXh+MXUHhi8YA+C5dZMObE0HfbLEhc2BTJ+slK
8BYQKr22FSxikhuSSmsjOZvPvrUyWMZcGKXgbDJ6CmqMvEyv/hIPw7C3z8Y8efbtZIszeBZuL2m3
IUtXA3XKEIEC6K6Rbyc8FwzWgTTN4US4L/l05g/MNrfjmmjZcPKhxa3MHb5N+lgtORqFtNiz+i2W
9qepIVRdfskO4I3bkgNsE+WDJ5EOOvwnb5nieCFikHISvY7Eo+5NMfUNyekIGG1V5BHbL1ZLtF/c
/xYCsMtNswALzz2soh1SgtsChGSssCPzJt6yRiAITk4lDlSIUSYEVA6jOTRJN+m1YB2qg/QyT6lg
T911pYpuaYEg1eaugHmW7jXz69X/2Ln13SnTG9hLMpaY2DQ5cQx/8oC66piLH92dU4ZpRjUqHbyA
sc1jQ1yRnfKwmyYj4G3bbYR2c9z/DXuQ92CEDYiUIuUpmcSyJgq/HyROarcPuX+3kimfJxxrFVRu
1RYTC9sSKsLrHVtt+N2xKGWfTAHu4/ViX3dALQ39yzf5GDgo1pONqMi72iv08dJyFy19UcdOCaBI
JE4Sx80VPEXkP+Wv1Oh2GI5xJNe0nDBrZ+Y+W3KW7ksSM6Up3EGp/sWgLqV6bRdJ5JxTs0I6Aivl
B/s0QIosSmexW70oZrVzLM8gXSuO7ePX4cXJqaAJ9gAoAIfxyo7UAvNbc98bx19Mao5w/qOYBdCG
JXoPktfzHcw1RH64+uqasFKFn6/91/wAqcxCBNPbcNjRKAovFYzstPtxWM29wXy83ifiU92iTz2u
hCdIpAm+XYJ2K72Ui+tdNk0BaF8sVaT9iPyY3Fl1uBDzKcmkXW9fp2FCMMkDIUZp+3h2uuTloliQ
BOdUBUbyTcZQaMQ1Bva03cCNgICih9qvik517155g19L39gdG1TDwgjVlDcFWzcYoPwrqDKoa6vr
xBb0yKGxlFHplN9weglQuQ1c+Dwt65y+Wr4d/IslxI6IpCPSnrXkGHm1D6dqQPkS99d5YDn+qxgL
by9dzlFd1jXRnXWy+6eP6A1+vMTqGCX1h1qT0R2zc0pzycsgV2xKoI1ax3nfquSnM5DfcDckRX/u
La4UeHserxwvhT/gIDEoV+DkSRoVG8BOWz8XxpMYE7Q1w43pxDBp6dRiV5BVfZ7ZMcI8y7DiybxP
PCr1OQg6HKbLHujqftH+XBtgpk/j5qkvEYTN9kAGKEN6xcXLIf0RZxiyiVn8nRjYFmC06C87/TJ/
F2Chx2KKjkOgYdJT6hqT4eJ+0T2uQGaCxp2/cDF6nWbvJahiPp9q/fXCzQ4KktmzWR0ABFXtLGDx
0h3CKT1Vgk+2F46b5xDr+NRVYzQoCl7TSPOHEs08Y4uM7s2Bt5WHPbcv7YE/sKgxCe62b5Nddsll
wH/yUWAEyQS8RszxgkD/Z3onwRbwKnDKaScPNDoQYChpD98bt5Wi6gWML6eQ1caTrs2Yt757asBa
naKJ93pRxjKePfpxXtAjldjqOAZD+w73ol9H33VBBt4Udg098Dn2cOzqQWBGetlaO2d9vPZ/4lsR
BwoEKyNErzkuB0nTekm/OUoZnQoZT1erTOUlvfY+S9pA1bpTks9KPWg70aatRqhSUsaZn+MAjvKW
zQgdagKtuuUGk1Xixm9og9KePPStRQq71T1Aw/rR3k/5m3yhAMjptBMq8rG65kJD+yYJhjPzppBu
/KPHsy6amhyuhT4+pQIYx+jK5ow4JNDkMclcaBWQdVOGLR8Xiq6ztrbNBA7cGbSKuMCi6MXOMfoE
+oxsUr8y9aOGjGvHreTyyeN67hn34JViatbfwQYaCzYFMuX/vSFimLC4Zczx2n15zuc1g1xeEIlH
Yfybhj+UVx3E+aB3mmLYZBEzJsk3twt6jJ+J7MNSl4cYXeasIEgWoAt70rvZCekYf+J/LVs6NiLV
m0ohTuB9dy4TF9WHe7HS0bwMEMGshK78DuBAIulsgQ2KfAtRZzcTEQiqfok8jPTZ5NkHqZzrq4gG
QRmfic3Bw6dD7l+mJ9V5K1V+GsZMPsqmwcjS/MPy1vor7hjp0YmAlZ4K4BUESDFCfyL48nLxk4hk
Jb/XDqFGsBOFKGWRau/HYY12hhbN4+2A1uii8X0+KKnmhXPhaTE+V+lUuKbZLKaXm0FH+pA0JHeK
Ww01aRTwwlL7eNgImTJVJkzLxuEeuQ4cCoAZfotp4SQJtBtZPhx/wHb/xpqQzzoUfq5qc2cf/AML
0g3g9cPlVOcIqWEcWU51Nph6sw5r2VOu5hUej55jYdW5rr4+oGs5eyt4DruGorBdTn/d4LHLsO3U
D4Zn2FYLKfUz/jpZXGct/3x5RW76DCAZFXmB120zgHbpDZZcSE+O0HwN13Sf2yN1bpklmdqz9tor
THbU4dJ/X9K2kzJ587eagGbr+lDEQkBx7xynk8I3TH0eeoNlHXhzqaYMvtoEJN2d0+hyqZEZsRJm
dKnCroYN8YzHXlC5EZIK+O83UVHR4ElXOr+pYLCyQgGygoe/S1c6e3b/PBgPKy5qkKha/dyFvt8p
gYg/qy5wPfDmwhUivi7SsUXRcfkJOYHxY8Njnb79/gMcVkp1C/JgEY6W7KKGVgbqTdO7pk3SPPPA
BXTv35uhRfr+IRPMy+OKrwquDZwx8lS+QtFGqoL2cMdspIxOUaDoPvrBhKKOBRqKVoO6a4kIxCg6
aVJMIhAuVA37F9ObQqCSdf3JpVix+8rF0iJyn0Qt5S260mWwkEUSnVTa6I18YBWjckZ1lA6bSuII
nCNHswMQRONH7pVfUBAmVwkR+bmpDIg+AMVmwlIESdvSBEJa4kRHdGb1qjuUj7/65K/1Ms397ZXM
3ef8ZGHizCUtUAz2FsukV6ok1vqsrsS18awv3DGlY6Xw3DbRVNInrrKx6QqNq2poYXONb934hpp0
u5wEaS1GsiNeGige29HjmzTyku9PaQcGp8Vfy4HORrLEHqYSb3jPSBq0Z28UeXlUPWlY0CR9IDzh
UCLrV8/8WJQP4PbHQ4FulkU9sx8LF6QM3IPUA6Dqfv332t92eWsBPxhPkCSoK/vsQDvdAU7+ddqe
mo7W7oeVBYVYP2ElhwoeWYfs0rD9KSUkbWDzfFVlUsCb1HqbQ6DSCrqO2j11TgUOmWjYfkM5W/YW
nkemFi68Zey85XwyzpNVPunKu0hS/kavIGDllxBOa8XO/Uvw/M8Ga3vwYolvTyIEtd9nhphtMobM
V3ENyC620I/PBFBP+6I1OIkgeS4AQq0w8HKFczlxOqDpTMifsCof78l3bSy8gwm0k6LYR12YmqXV
4wPkIWsVws2khDNzDMGR+hy9IciKTA6o72sa0jEtMai6Ea5RH2QL4KlKCXbrxVJI409lxmA8mNNU
I2PZ4kwT1/4cbFeoUQUmwdtLN3K/bFczb/2NOgpqukZGBQ+M6aM7XmOT1H2+MRLnKihVyoam+/lh
ZKy/aKGoianQ/Rtde6Pr/vL7e4/23ylMJcca25gpDQq/noSOrEVh9WmlxWq3ssRyCSibALLr9GDZ
kY64eBJmkjiOKGXeSwjhMP8ZMn8RAmHMtzhtXi4tQuQ3anFK3RUzpuXNeQa7qSKV0eFg3+3jm1du
QbFScfdEX7G1DzAe84N8TmtLaS63klvNr2m61iRQIQz6cC5w4Dj91YkQPhpZM9KWGYVXWXiEF4j+
OkuRoN98A4hX0XmOD0zOvRDAFd8jP/35j8U7KYAKxtqjAbONYp5EW4qSBGeon3c4C4+vCXg1DC6Z
e97UhIyWchQAShOxIl9GN6ELByIYrvAq71x1LrVqsI7AY7EFq8j9H74bIBoRjawTVcI8U9gYmqka
d0HPlBq+MKn/pt2IBsYewhmMPcY6cHkro+1d6sKL4bIIbsYEVGUtzkZh0kvTrxjWdjVebzy/fEuW
/K6XMOGCedOljPHluqDacIuIxyVlOMlAq2/f4v0J6HdlifK1Kv5IGGfyIk2yybSIWUYD7ImB6PiB
glNChEdKEfeEDZoYT5YscTvvRRSUxBOMwUlonNHrPJqholuAYWCdzuYCXp9eO12xBPQQrWZ9LUHA
BIGfMUAGfbTf7i021sGdC+RllVf2QQCte0ztCYUdZZNKHyd3+9InPlXgPgO+mxifjz+5FA+hdEes
6ZEkKSY7kEpWzz1TEp3tJDONtmpv+QERn3TrwrxgCvjdG8ORoT5ugycTrTv8zNEhI7T+z8YqIzYG
/Ct+QWmAkC3T5hWdbe/nhtVz3EhZL4ObkYRb0lFKa6h2tEKA+dRYsVzxhGt64xguukgFtpt6APwD
M9uFC2Ofqy+vimotgI05KCTbDIEE2jbBjh38DN9SGBV2SZ9u6eI99zFpBnocbzNr9k9sRPBKFFaL
mN5qwsaErU9W5wtOa6Wg4rGLBF5LLhOEmBY++H84oRYQm1FfLub0NIoqugcMux5v+2zHpuZRfjZe
OotTE5hEGhYA1tUuO+Wf9EsT9S04yZSE+P26PuBR471yn4jOywkb/LZm6Bueo8AoRftPsg1JR2Nd
bwmYPTJaQeLbf1dtj05vFcw5g/a3LmBHM7OgtRvJZ1dKTVroDoMVsRy/iGWggLYILSrCAVQAHjoX
k8P1OEIws2phsXqJouTWtX3Le5NGjKd/gwmGufVOYmTmmBmCK+KWrmjv/DoZAbJqlohNCBty5po7
tThbB+o8AEeaajwo4XDzrQeMDNhDjJ29F7FCbyK4tZ0nia2chrBlfVJzExRVeU55BskXeaLJAWBr
ucTnluDuCmtyZx8coEW9+UPELHXpaZMUG50DIkc5VHzS1u3KhMg3tEHLbg73RgV4KV186KrTwKNV
ICD5NDj9urqlXrKoOkfx4V5jj9ssV+R3G/2sBu0t9tCfMnC2G/fGWSTESUw0tYMYG3Bby9elGGTc
clh22bfaZoZfXsdAAZUtsa0IuizH3hMmiIyxZ/5b21VeGY0k8oPhnK+co0Ztm/6Xw+oDTv3OwvGf
H48cKjpTLdB0jP7HXa8jGzfe018UqH/Q4+EqC5B8fNl3TbD46cn1YByZpwOQyGUC5w7Rt/3fPmgB
oF4jroiHWLZvlbkU5tmGytwYcg1iC3PgzP//rCBPW8WSALPAl1wq2x9A0vjcm7pX0maNDVHqxyl+
R22Q2PG5a/50V4R/mt1NhVQXWwdbr1gpI4Osj+kk3HfVYMsUbConI96LbhPnL2aAgboKQFL4ZztF
Y7Vqo70UbRcokSRF1ajBhV2q5eKOQoumChFgigAaSAPv2I3gUnWue7qVACmtl5TPdsiG5B6CIT+t
puNsRVQlTSdbHctMWsAAfC63hhknY/HLASPKydQklFtymY4Fr13DITgpuAwm0jvbinPVuO84nbTz
wjuU10uuzrcz0NMNuNSwH+TZwDQMdeocxCRGeR3mof5iJQ+STDs2ypXqLBkhavYFnWxS+wRq6Lbm
9shpOfJ7iprZB6uUUFziqrscV/oFvrd2mlxIxALevxdkOCtjFSjTVoBo49fL6lVCvl8XyIwKAqja
3G0jpBESKBWMjb7Fv6lW7YG1hAxD3Wf/dD0jbwagQrLA9Xjd8R5jZMcUbCrNE/CzHUt3DGtggvc/
s3//L8hgMqrQNFLwJ9eaVdYfzHp2RvjIfladjRqnIItw3HfDc+Y+ZWDZ+DZifzuXOAmB2aIQasqP
ORjWJRMeBetNHVfUwZSfdYr+2IBco7J7uEuZiGy9J5qdfyHTgeKwvE8CFBYMmT4FarI0RyGjtHK3
YMlZlDRWiQQoSrUsZpe3HxpARCjawXOPQhFnZ8K0butYfx6Jlu6vB5mE/y29I0dXDnHBPT5FNFzM
1iQ7S2Xl2yZlWkpqhi66yb7VKaw3zE4aokUIVRQNiYZ5t1oiRpnKhjLxTMzP4s/PYyNGUvNUjw71
x6y2JVgFKj2zQQ3gYhG+4hysB/PsZQQjLG2Bm4HEElYqZwMr/P0EIB5LZfe8Q9R4oo/bJTGYFQd1
kDkE8HPPtRAKUfdHIDhiiZkgYM29MAMEcRt68SNLriUG3QAG4B/kq+L8Une3XerQRxbty4acbTVB
yl7Z64BTITjvfpzHY+QhcA99pLkIvmxlAO4f3csteMqSErL3oiJr0d4vbD0bWRD2bHNZ9bVu4dug
k0zLF4Ciq5XIuSNQASIAP5XJGsJ21cs2Naa31QHRx27wVDvIsu5EnT0Gqzl5oY+Rzsc1C9wZHtR6
12NhSZLGO/QzpFk9dshY5An56w6F7WdKbUd/QNXwL+2HZoY0iimJxtgf0n1VAFZ6/vARNfpDiO7z
P2y5g0ZKx93Pwze1eb87wbMJ3LlorFCxCLprB6opPhOW3NPy/uNsP2FgECSv+HxXdI1T6UWArNM+
fVK6VLX2DWm3RqmoOFqucAC24hPqXYFnB2UnFr8boivB3skVRDU3hF4PjMPi5LWWn+sVo/dNLpXt
Yb0c3J4CTqycYc8rRxnCAGoQ6Pd1/lfIyAbkZHuvW0xZz0mqLKsTPbmsC7bnoEGFQTc8gRUTd30Y
FjiorWCG6wFFwv4HTdIaFpr82nadLjXjjz9EznJB832oW/6DgqGqdaUIfUyhYy6BDwOUGiXEOikw
VmjGQtP7f9Mj/0OT9xlJWF8mg55DdbNF7ndFBjso4AVhOdvSAUWkdeMw+Zi7Q8uVkCQWHXtZL0Ru
phCxZqTSCLrizn20ysNTRX+2HET4mm581JcgZEPcRuuxnPoD2p+v6HkyWFvvpoPQkIIc1KgSzItx
ZKzVefTqbMpjQdQXAHRXDCXh21hNY2344frY2lPDDTdCqZEWLd/+Vzn3ui+JjXIYJJG5m7mD/FZ+
NCtuumDyY0LL2ZC0kLkAc/V1eUwqel5hZR3vdWF0QRpVuesL6dHjdFp+6Pr5OYTElVKj6H6PveMQ
nbUhO7jEBFRTufAUI+Yf7hl6szlA5X5GpFdsWA3UyGPlRkW7jlVDp3XwJoLwTmE2ZdHX06bh5Kxb
nWHu8Qh7reFpdF0GetG5gwIHKfkDmWW9o2qDFMZr2rgTkAlPhcHfPUAjPx6bAtPWl+/CcGaicqSA
/gjoXMMLNswaMLvADxPk0rHHGz0bGiBBwegFJRDCgJlgRtswZ0xcmxKlrSzWaa5JVtVg8dYxEKka
yFmdwdiDx/aFBexSWvp5KdgJHCdSVbd8Y8Zfd+4bgnwf2gp1a00Uxbfqj/k06/FrDEyHy12hSjJ0
jORSXw91QAgV0FsWCD/e+g4y6VNJWpMP/fwYD3LZPRQNAv12++BdNVxBnmT9NloFc6HIuiHzTrHm
zLQY9//gi3la1DHVUV7luCkAOC8KL7pK9eSs8B3lqBtqysQglJdgNtz+EBz1676So8wisz5QC7cI
tP1R4IQFIo/T0BGUT5HBKi7fCmMIEmxAghElrhrmDywMzjhWM2lrRb2A5Gbff16a2WDRuiL8+NYA
yXdmzxGrisgAVgjV+59vM06eDx7mN70Xvtzw510mqKgaLlvaIE4xtUjrtLSP9U3LE8H3Kz0ShWH0
hgWczmvgT9FsMUoSlk1MqBJMqEbai64LhCoyU2HKNtRZn28ZbWwLM28mRqJD8cCxuCDVDZ57Y2u9
uh4pZVTR/MVN+7GrM4g3pC3bDaaaEhZFYo8JGi5nt3fnZbNBRaop/2iniZCXmYXWLFm6FLjT08/Z
WpBHOL7MVs6NgpSRa6vKSN2s58dcuKyaBEQCQxyx0vm5xAdyiXzMtI6cl8jwBjWie7odTb1MG5u7
XXnFWfnkh4jFdLtUmbh8JGeGyripwIvuPf3MxBxMHdbnL46edUtGSikvKTrzikNLg28sYLTFkXmY
Q2l+9b1gqHjJISHVqSs/yZHhQCEcj5/iYgY/eI51t4+Q2B9CjRYFRqn0VaybveJwXdypql/qK1Fi
WinfFzwBWs+uBIysNNx5BuTMyj16/Mc27AKXckVElCgwLb4SSxgAuOSohKDpTBStoG+uZ5Sc8D4Z
21vFa3WrddIfq8iYrrrICgh2kvE/gkv1yIyrtsHDbRBCr5Aixfs5H6rtaOx25SO2aP27FXIkFyG1
bKMpe4cKjG1g8mkn5F1uRiHooyOpYPtyk0CBaUwkLVB0H5u3kP9gTFhHOtASf/LhglmWm6FAlP0A
4N2d1szYQJuQp6mHWT6GDrgKx2RGgftIBHT0qcou9i+gRbwpe0PeHwiVzN/LdyV9Y7BKwFhVrRuQ
ooCvuHf17zS5AAeLeeA9yDy6RX01vF4rBqJ0t2LKBq/5jNNAsSgycqzbijfFw7kL5y/eZeDLlAd7
PxI0vF6EURtsaOr3ln31L71GuqFlhRFFseI7t5nwH4x5VvHrGCiArjDyZXCyzfIMA3xMHm6/wuSu
mlViAS9NNkAoXecWKlvu5m/xhcUbKH0mbl1bkqUXQB5ilzZc8kzLcb+BT3c6SReQMmcVikq+THox
P4Llzu/kU836vyq9CVj2ErUQLfx67xb+GmXJIenCdckToCDo4Lat3aTWUOuj/rt12nJ5aPeF7moW
1sZnNysbPghmIrbAkeXq4qoKLuwLhdcMY7qAomp5Mg+bZ9EoaG5A2RpiIcQW+aueANRULKUM6GrC
XzHc6dcxs3K2l5CraxXLuxoEo63sg09XM7dIRaYjdWDk7mmauJj56oB6Y0I+6jlRIOJKYEPyD784
7dMg72oX8I1CYPAEgpLcxQ4oaxavjdg6tYYqz12eGw7+w9RoEfZhs6ZQn+1S98JK9iFzzl5YKkJm
2brlQrSg3sRydJN1EyBpEbDR3Mu0PC+ZUvHFTJ3hGAoKmmVGfZ7nQb35M6vX53iRqRdY95Vude/y
3fLsp8EF+jPqWHoAUg2cOdDmCUGY+Iqwi52J6NuFgTkrxhUp92rNQZQro5Ndu/k8OAUAau6W2Tbm
U2mm0WxncYoB1fxyBL1PchSy+y9VCuoVqbDjbi5BoecoY/7flnDvrcUvmRoIIYNxEGSUZ7NnncQf
5Qdgz6qyFFJHn0uSkq57bSGczh1lfyMeOcH4KEQKIOIsuC/T1TdQ8eDapfhfZSJY08eqwjqKmq20
sw1NvyGJDzguFyKzg4pi+DXKlGNbOD8PlFXo8u2ayW1AvZCD085K8/Z/XFpiTs+90352kTAtTC0Z
84SBp13FCDXP7IpqQ91OTLozFJ0I4ZI0rGLR6bpzzOdB0CE0lJ7+E7xRGEa+pr7P76r/YTeJ8Fek
Xlrxsbggxu73SN/QDDDX36CRXKICXuwLyGI4ua3VddClWa4T52f6WTS20ww7ENhS7JXpTpeuH5lN
XFagOHqPimrsnRCJrjQ3N1uFGxqVmWdDEKMZP8+68bCg7bA8n7EDvXUeorIivF+gp5Kw4pKq0WLl
WD0KWQ/n37hleE59aL/2zRd/QyfsyrJIWMtIl8ELw/G9IxpI/iuhFDU+L03kJQHSoE0au0UAnvAV
5j3mYd78tREMrMwdsFo5Lsdg3bXIAT6sWGDKZbjmN6GqOKQd9R04NefOm6a5p1DMqkOQCZ51mhFH
yFyVSgaJQe/UTNZav5cU4kv+sn7dKwm4ecs3CuJFbodZn491zH4djCuXa/DEDUP/aXoEs2STO21U
ya+fATt/9SF+1+OJhe97cew7tFkSxdObnOdS1OvZSBRpzgLS9QecRXcWQ6GAa/OTJ3GPZ85vyrxu
9xd9vatX43egql4S+nI8Nd4P2h33aDZRmyHleIepyes6cMrc4xJpd5ykaWv04J+sq171Zdt19wWg
O42MiHFVCUJ1O+LnBugssnwi69S3wXLzivnnc8UC7sYV8TCUyiyifXraPrcNfz8YjhVJL3uMpeJr
3MvTB7bmcpmmYESw5KSov6DuymWSICfcKIajKN6eBe+iflDl/GCRR7CTt1IHVUvQZPmyTZ2NU8Kw
bvHbpZ0s6jWgsQkUEg6QhORFtDxciW9WoMh5xPJvxGKatGR8N0UYipLXZNH2vJvS82jVzFFbiWac
58QRzCbSeDH6+iYjsIUXfxx9DiKD1FfMkluMPGzogN/HY4FvFURHBu70524KAO8Iscz2bR4QPVuN
97gVTitMmJNlfScOGykM71wRT835qLdFxGe4+IChxcU6zGggZ6xwBh/Cn7ZD/VRr+/Re08UMP1xs
YlBNflawXjkkgAvf0hEMKH74/2hO5hz1UlKTEM7tQ2vzozinTg+YicUcYZ3v3a6CW3haya10c3Qd
p4O+lxQ49w3BF0lQpvw3rXkdBNkkVgJCHdPlh4CpbwMaKBAW4NztVLJWDwtD6vIh2zdZYYBG4Gsd
ORlMGTzzLjyAacW3EsN32yDD0TgVNr/wRGpNKsY4gQTntqeEuqF6l6aFCFrmH6WOdcFAb9D70qV3
LBqdfzhgY3iJMzOhaLQpJlaU0ZGE0KKsTcO+yTW+TTDphAiTixtDXe34Us8io46RLfmQw2KWA1Xg
s4JiKqqGi0rT8TyhoZeKR8X0d87cHlhv9+qcFnhXczrgkJSdwPahuByXaknZUHQw93uLOa1mQri9
pDieFa40d3pXEqniZeMvRyzPyCHvORDAmeiIEsk7CMG8F8YFqO3VsKMlz1D49zPFBIA8s56Eim+1
k/LcDo4K4aqI+POHs3+Y8U1na480G8582fvn/aZqd/rkbU4ucjsmwSdqhEi7Yr2CPjAKAB13c0sP
wG4rDM8Ret8TdtibEQ3N0qe+oOIiBRmGi6Dy5UQwOzZHruQwjyVVmKuiUVFy7f/RCiXyJdqjkaJ/
x5X6AcCcQdOpc94ijuT/zYCl+KK8N5sTQQvORLBTa+B4vAKOigwYGW8+xrmsVXsln7dE7T+XGnLP
GgUnjTAw1vRw2AHM6ulIxZ7vOAx/+p1qGpoBTvNM0Ceiw+pQBgyyGpxrHgjI1V8tosqc9S4Z7UMS
XPU/SqQFYHadmT0s6HUvuXSUeaB3kYPMySv08oqNZtWPc8NTlZjoAC1fLsigetMfWlIPC3jbLBDe
2TN4EQYRS6fn5IzDfyPMfL4vKjoPxomK1jFE1RUA6iZQ/Elpe0Mc7ztkG9wz0WhoV7afGv4iWTPw
UpqIqAMRW7LGBkGq3el4fEOl0EDGM0dox/6uLi7ryS5B9HdKVjD0SotrE7JpjJfymzSdqBVrps65
c28eEG8GHVv0bX1n9QvNwxyXsHJbl0VIO6wQP12gjY9U5t3FL7MdtZueWQmvAXhswiQAZB1p5+Qg
QBcnJdPZdboPE0eT//MBwreH2piKygPwbQz1fHpIINfJ4SmwHQ1UXAENLmnT3NbOGNP7RXFcg1zK
0SEEpw9JrvQGX6+kNgu2YowUSOKO8YXQBhwN0wVBbwLkTWnxpYIoZ012p3cxHA1cjG8Cdt2V88ES
+o16DNfNMH1ev9c/p57eMN6lvzX05or58fQ+lG9X3lkLCamutABCApj138Gs7N6cu8JDKZT1jiQ8
IASf2t6wrWVrhGd3+AZQc7hmSJ3++RvAc98Y6IJGY+JGg3SDzbdRPOhtjZ0phJJ2TITw4YjlG4cM
7RPSXBJyu76R9adeR5N1vL0H2mFBMHZxly82icGZ+jzhfl7b9LJo+Hz0fuMvh3pqrDpEY9iX0Jw9
mkfdbyw6nQ6RZ1ExRtSxjToS62DVpVT30J6z+yWrxAvrSiZjd0Bygqy7t/QCicci3QP8+/PjGakV
dT7LutfkExeCXL/4D7Wx05jpqfqQ5SQKuk7UECJdQJ+Dm8SSvm5VunPxCbEuwcMZ5uXxSdKA43d2
HJ/fWmJHWuYpYfl3JmSrK8NITosWL8Ii+pk9fnl9UsRJh63WWRi51x0euj54297diFY0wtjzYIqA
5SoyiXyYmCgX1L7Avuds7qUM7O9ZG9KL8VURGVzNvLur5sIzBPHkIvImV33QXGf+ywfKe3MlPmwN
6J2OtBKcaLXGqdhkVdZ4PqrkI2Z9xM2YKoqcnIPkDloOw+DZSdRwWfIuaVHf5hXZcocZ74BSZ5+N
p+9cF1t5Dcmcovv/6ZwaY1jc+f97sbKwjtyAFOu2WK0LdzMiRwYos8psEZgVGNsGB35zrsbi5WAM
i6YZH+IqL8as3sTGQINK5EQTXvpfHXuNzuhxRVqQYzdSkZkLUCoiOAGTqFuVRaczkCpsdThyszVP
u3F4IRMmo+vPVGlorULPFvmkV5VP/Ki8Qx6eIO7HeT7rsbvMwKPgkziWO9JbVfcPUphKFbKL8OuH
NxwiljGbo8hj+PtqQtTUN54lEFVnMv9gmuF14RF7m4wG7txvfsrb9jg+tnmzw0BM9Lj/4s8f66dX
jPESiI4IVtBIfficLNRncq7mZwA3r0q/I8hCI3oVFQgpbj8OKshHG/kG1uJP3GOnA9v+fsAjP/n9
XQQZLPDIDHA+HzzkfEKHwtbPzFyu1wOi+8Gi+VUz4sa7+XwNpsRMZ4XNupon/A0ClHiMxGBqjtwO
xhNJdNlpilz7d8/4YzB4FaGDuuP76fHVazc5wS8QaBs2MPDzP4uzTnPuQug5p3HkJi5pF6qrEgkx
VW/X12RME0SPFvw8PT7bI2SB0FZ5ze165qs3XRJMU6Pufa707TQjyPNkKk17hwkycj1ehx+Pp/jA
hQo6raSbIhvQiyTNDXyUVhF7JEcb/gbcdxdldmgVISDM51q8MXWXcxKnARc0m1kVH+f35fLeU0yy
gh08hencvryXmBIcGFcvFnNrVthG61wzkSJLvBLVecSowCS6usoT/9tKaVYMCOMSR0a/ehb5cEXJ
rChUemsx2tB5l+KhosAYwUyM6k4/ZPkVu+BTUGHLPLVd/+LY/YkLsaY/sZgXuMZg2pCeFz8rfZjk
cIbCbTj/kGAj3zNZIWuirj6DtmgcBPYlWcUrxCNrnQTOP6VAbR+vCyhFZiJWwD3fBy/2J+cuGTVe
XVG62qMXGhsgLOVcb19z3+XxE95uvpaicPQlEhFGcoh4xk9eankUt9YQPTN8x3u1ereaGiOupKt0
gbuSGhO/gGBocbPhAXq2odRpwEGm6iDgCBTdVIBWi491AlLu6YghpGQmR9ruJ/UdrQEjozauLYPY
Uat1bJjnw8MlE2IDfOA5bRCsRqu+dizRybwRqmJzKJaDo/Ru6rQYTTI/uk2xkz5SRd8G/y46TtUi
iHiw40CsEtaV9rslDTC9BdYMVYaKjpRR8g1BzNEozvfloPNtOV9KuFEJRYKbrykmr2Eniif6B/+m
B8jfZyDHoU0vDVGgTxUFaY/gqIg3FSy5NTpGd91U/3vuC5XpY6P1oEwwCW3B+1aAxqnvwcZHcl/g
87QOQSwxTYtOe9Axz3Y79C2GgPgw0wfqYZn2pPbfweUz26aZMTrmbMl6Lb8QhjbP6yCyXI1mLLWe
5gz/YQJhirSCBlHYNGOIqUTsKWLB4eN/CRAEYTYaSzuLixMbJwQFqxhposLv84lCodJiGzWZjLLz
h2Z/T66ZbYCpFAnJivN4TfIcCa/Z4aSnnsa/HXdN1uQ7mVBEbnAHULZAkVuQSpHDsPVTGQCa6tlv
q4qxvpzls6NP0/HMw5uRjoYhe7qYKNMKpAU6C5u9LxSKg0dkdSaeRdKSqCeUHiTpn+LDs4GMbHV9
65ZO+msR+4WePOC0r0IJWR0CD1/ZzxN3SnkWefZuzqLXJXA49p7QG+KdsJtxkf3eXZgtjPXN3eng
JtUw9Ko5JNfD+Yo2YR+Eyj0pNNYZELVC1uDj/bgW0fzVMGH/dSBVUrgCMrqT5/HAUyaex3nz06gS
6W20wOIVS3M6hJNa+TGRlbsjg6GclK8Zte805bXKfcGyXJ60hDIktsAKLp/GeF7AzlcUROrR16ar
yn9eBU8NtHC7AGMF/b0W+QasZdWtaQSDLxT66eV0zOh8MViEFrYhJmj8sBUnrctgG/gCkHPVcv3E
4Epn0OMZWXoU2gcdVYA5DB66EKlkMJCsFDJbqVH5sqPsXUopodDQQZ8FcI2ykbb1jJ17WR3HfXuJ
gpEI88TQESZW4PhswJhpjE+V+g9kMwj9+uIEB3Q59CuM9gkHiA45vJSElVm6JjczBuTkMndHQg1V
u7/Mb3sGQg209Sfi84KCb/eV2Sqq2UWMHLZYsuMtcYZzM+SFpOAqOGDf/Wgxsih8aYJNmNUuqZbm
W3oavWKnmTs5aIGgyiFJ0ZWF0K1BVdXsk6Whwtblta0NHJ5lS9mYGfjgMPAXWX9EvURHNaVGGX9l
MXO5yPprbkMfIZpGs9to0YV/sPL+NDFQhG5vScSQi1EzAX+TlkSVOin4ytm6VugS0ea3yXL6YHXv
6enMbKXBt0NuvrMTyY5dOW9KNt5zJz8xE5LzrtBi6XaJmXgVa0gqR6dB1a/bNk9DQjovGBeGDcfR
Qk8J1BXe3ge5gw6/mELwC2rKHyZk6Sl/S6CJTR/7oCzMwkTNKa7t0sXH7RIooeAQhokFtzIZhlVX
af+Uz+6jIol4NkIzpHCReuFVTcyOlM9wMLu+6kOvWrK5zab/8S6CndOnlZ8oX9yw4SgDmUn0kwPl
ELUws3NWvmfVsj4R3u7rf+QT8giOECFlopuPI6sF3qgHIT0++k49YvvAEOfHJJ9GvGJkyJbPftTN
MN1Iog+/A0p0Y24XWzeV1JVZws2+HIGeXXJw/4cdxe3uCJ5BV1RUYHYprxoyFMlAOWKz+UG9Adxv
EJsHxM41oPpe7GSK9oqaMp+4Z2OwN4zJa4WDwCLACXosU4fkS4PHjtI3/keFUfuqoIUjlXKuO7Z0
OGXLrEN48oxIgA/bryEjnZ0af4zzTEcZnHlM0toaqEDo4sBTszwZw0a7Y1AsAobi88ZJHRdVpwN1
FqmawNr4TAXCiNH2+2F/ZNpHsyyFcIjUENlU1jghql+xF9QM2YGVsHoPPjdQbb4vcF0vx3BcQuGU
Ktz3N+EU3e7BksOd7hrrvxesO7XLXY0O5pFItEIU2m+ld0sYkSTyPtmFL6qM937hybAm5SdAwkxP
UK/Hu5hz00NXPDXH84J9Y3lpCc1hJ329rxLza/ITorIILp9dwJtA+763Vj6+1bAJvSPLFnwjgacZ
4RD2e//qe+d8mb1PYlw8obWti+NV+lpF3lX1COIJFfoHL66qEkYPDqb41caWPW3LbPgRfWLBtAbb
ZPWMDQ7tFsgZJoj5e3hvSVkFWtbOTVdGdNBg8v8aCaWDbYpvsuOeWKLFsJxEVME9rPCeGwHWbOFF
pdjzOrwB0/+CbmSEV54ykuwNArjmU+K0T6+Fw04VVAGer52C1onbSo2Nvdk5PHINo56AOeeelqLo
nByza93WEFgCN3porCZn1lGrdrFhDOJvnuH7Fl1Vk7Gp1KlSOtjXgqe6P2fixkO+tT3TGx8mvVbs
TMnZGyivkll9hx35b0ot2AVix5cyK9S9A5Xkchp0+s7FcQPnfT8gTmHn7oxXBpYCyEkelahxk2Pg
Dsy/OHz1yHVLrHTFEVwAZKg2FkDrlq9yzzwIVM7uaGKMKI9I6wciydXfvJd2FL3W5yYBWpwQdlDo
cOOr69MyHEZauRHijtq12L+8UJd0g4g0hPg/98Wv3KZhyem1Njbr3MVwhQe8CQobxi9oFL0BWUyE
8BZta3FRU+EJ2egh/CUiAmzzH0J1zNnrxWTmcfs94/EpYWP5YCS3nULOxuhAEGvYustCtYuBrq0Q
ByD1tv+g5uUbLH3E56Jz1vNIIZKazXUSfrplFYAR16IwO9WlglXoRhOKyVyEJgxr6h30dudVrpWf
iuk9T1D8Q+MIlQdC6ohWLOYLY8nrOe77XyAzLWtCQHYpqlFAiKVwpp2c158tBvoAXAv6JI8YRENk
5MVstHMyQbhB0KcziTZ2zdPFMPXxfYxZ2te+E2z9u2qRbWyxf/yuZTx2rPLRc+gPQNWDw0lfleN/
W8UzvzwpSE9iSXmr1FmMvxRpmWGuYramNZm9YXvP6dTymDxgImoi5h41OnLCEIwsYsElVOuj9pyG
EBp4X35SgrUROZLiVvIFCtnbyAfPMO82+fbgUgZnoY5r5knA01AxyHg+POhxbUDfqQPylO2ugghK
vIhRe7mRxJAnmLQWW8l4MgypXz8NJjZCPQNfqNYY6MEHk1tm0HI2gnb3k1zZPV8RrdWR2cBZQFL5
hgfQ6OKYgT1ploxSZieRRtOs4y4yyEDMXd9P1niRjbJ4eiXdK16Ghs4t0e2djuN7bfGCPIohDFo1
31fkNJdpxDeweGy4Ununm3YAjMPF0aYECHAW0hmQyJZG3qTGv8KPzXFyRdWdaj5HAwpl34GOsJaE
7oxB5BHdorqLdutFkHXO0IS4+1bAOWJWb51tovGvrDOzokeQztc/T2xL9sofzOss5fmbTMHGzq2g
UgrkpgizeNDnkMvzNoODU+ofUGibBlHyrhI3/eqXQ35PNEqn6pr9ZvErDCaKyxEcKqMRjZqWIy9v
7jqbiNc20ZUZpaDKL04Vnqhh3wAN1WGzC4KvlvUc/5+aKn8t4Z+IRxvLsPIhzZB8iQb7d0w8IzB4
KEw/Fb6c0To/gk+aOdvF0LwMRJsUMZw6hGYUSsGad8VD8rQW5AvC9TNXwQBhOvkj44KF/ILDmaIf
R+e/0Vtb2Q0lYRIKWtXqOpXS2Nk3sEH1LNFSrmyD0vrPutM64DAix3hwlp+4JRREbXc/PinsNotb
RnAwPmV+YERuS8KeCeHXkpGlQiI0b4IBiKPx6YqRMvg14gj/4IMwAJRcqdxhXKlFW9r/kyp9jNh9
E87KkyB3HdCfQQOCFqDyzuz9BdqJMBOqyOTeOKhcR+M2I1Prz4xGZRhvphU8+FT4y3N93iIx0AUO
RkSxA7HXL0UqQ/p67z98wFUiOSTZMv8aTzOEO38vgKJVdzd14HV5tHCLI9cxMWPaTP6x/xgIZfM7
SpqHMGzJsHudgJObByV5TrN57CWNYguLrOifRwKUqxwpZNam8mgjAPh0pDhc2dmVMXL0ALQv1QV2
WzNPeRRVMzgPkGpTcKb6quPrdJBPrOHWt6z0yQNmDFbDXIaBvSmqiL3ADlVt596e9CaRXplKDoDm
R8MXME7oJ81rmU/RuUFINb/3jKyPnKS/AhchIuVJazYknhU0Ho/uXjx4Tgq7OwQPzorOrK1NjIRZ
Oq6ixSX3FKqY3ZUisuTwvPqxQXKFgSWKOhD3iJLbnROb+Ib1HG72a9EoDsXTeAZH2470CRV4vNMY
PhwPp6FppML6yQgwVPxWYEOokhChmwbr/VKxdg9rdnbn09lirMA5BU6BW6Hn53xQIi5E/HI2sCHk
/OaS4Kd7369l8RJKl7KvPXHh3TyB00zDO9lokMszP+AhubFT1IrfKz7XXEFNpEWYbHU6qXJvyVpN
t6lj32QOmklIK5fvEkaptuMD2lsxcm6xzXNiTwEp73Z1wFUpYCTVta02T1wHk4tiXhsSqS7QPa/4
T2UmmosZsYfp43YEvmQyi2GxJYcuD2Uy6V1k/fQjhijlxFp0CSXd9eopiVlh9OsVhsYZycGkOBKV
nizDRbyYp51Vq+ixj9ymMUluxhnZ8TCSUIY6EEm5iM8zwoi+e4p4bFKgMueA1ura4QLNjl0WGatI
OyDmd3pqzoCrQY/8sG8w40V+DrRLDp0jPvXgAw1rGB2S7apSGukUUKo1wqFJxFT2DPmwp665vjpV
AVKE0eJzsPknqsIATyOGtOBcpRTisoF0sExmLSTnP+Vd8T4/SKH0duFvRolz/Gtn7qpnDNnHPjw9
x5bnSnsXjenBYUAoy1AWM3Bd0k80H0QwvMVEshzFkybPPgXL1gS7+nMxsYCyN32EfmPqqgaod8Cu
YGhT3xmncvYow2i25o29RNVAS+0wJInEgCUHz9CD7wazVIXrG+y+7pZf25rSXHhZkhaIKrixu74W
+n0NOuCO832GFlDcwXC9jFgHHL6WGP5N+DocTjri9SSHKvggMq+Dbx8OlSEUbd84aB9fAb48CS8z
ysKT2pSGH0hzJar+4sjBMs2vXSfTy9keEFR+Qp8nyde5mq7a1u4GTubfa5xWO61rVIX5zxW9p5hS
TY+7MCs3st19WqTmpmlsq5Og9GS8QTaj0tdWIMh1BaOSDhJJZbbfC4KWye4BdM2yBTDffjM3JjbZ
N/BZOhuDwwUrfx6SQyNksYoOnY2dCEOri8VB0hZszmI1q8CuAKbcrWW6Rj70HC1oy1BH1FqyWgJF
I408+Qmzn+5UD/3GHOf6rvjU929bc2JiRC1048w0E4Y8FC0OAn2ScIakECIAv0MAh1TirKItU90r
sZ/2Lb2Q3FeRuwGQJDvhj0wkM96LpxERwjHZdp3n7h4DYeE2VOow+lQmQ6IdMJJXNQgl2zTqj+gU
G+OKQAH6QbLdhM/rKB9mNxTw2dlGbg/ObuAvuWP5Q2fyg+3Q3wI1l46CzcsI8aRjq81SxcLd3KW+
EY27wViujw1JoesMHiwrYhyXn1tR42B7qc44A6XSmcDjDCpADnSRMJB5iBSiU3dBND+6v5umm15Y
gC0NYAWP7FHIKUMSObwMXGX8w0cxJYNF7/uVBIokCmAGSAvO0nffn+hPgXmrkpCbdCV5QEVzcLQw
bJiTWBI53my8SKhi0JOBKMu3r9sc9D7A6l2jyyysOtFbWBkSs1rF6fZdTH+j7S1eLY67m6oIa7WL
s8dUCUFs1Qd/9HEuqWWFKfPSb2Pbjt8eSwwqZfsBroqibxcFJpihGU565CQeFh08VwCCUJsDf72v
jgFTXSjc00b0rQpyMrEUKb3MHAF3ypfWMLndFVAHWuPNi6LeX8nijYriqYK0xmxmAGMf4dpFspC7
y5XzftteRqug/KD9zi3JqXWejg7h11/Bg+7WPQp1wyNuqbcbiMGhZq0luuX+0pnXDLpl9UX3tC2N
jZzoxTRop3U3sGQ/W9ccPow8HS7E5SEkt6om6u3muqCT0mG9GkaogYT7z1r5y6CQtNi4tlVsAjNz
Xk5tpMJfxFBY1N7oN5FxcHGZYLGVHy9SSsIKPJQMPlKRjOoNXZqvPtnQ0zCo3NpTembpRG4gOEtm
1SCm9Eq763da6saHVUocscSFX9kHZdGRFcrDIg5xGrIkVUMRtKfN/Km24fsw9hrAW7tDiem9HHdS
f8zcTYZiWmwNrJAickZCnJlFxjwGp6rm7xv6EuN7k0z45Vlyv/QCkhc8+M/MDGAqCMQxT9sefLw3
TpXJG23e74NHMIAhJoYHBaiZutTHcepezUG+9z+ZwuzQNgd+9ZQ6FB+y0/FhB4H/qNdJqUuT2HNp
Wjc4vDjlg+93RcAyMEyKKRhSGY8ATeVjY8HPD4XEQfB/RvLDxYJOyaYlLmmZ00V6uGrjERGy9gbw
pKyFbCHMC7bYtxIou0eUDbBxTbr8UlpNUiOpUsiSz1jJJNAPFomiFl2gOuPOSgEWG9UeXSmtt3Ul
LpydV0FPFlfDay2Er02bm37V5EqJv+kAKBbPTbmPEtgv8gnyu7qk8+9RbDzjjuIa2zEU1zZ0XS13
UEdYWJHzftZq7Hmdx7e3OOC/DhJ9wW3RcHmkf24SEgNK3Z+9RWrej37Mz9iIG/O2w2y0bKyKO373
KfXQMS5Zn94gSZEeykU23OFf/M3sPpMjWoNW9s66jZooHPRRR0N2MVa7FH0XQ0vcS/JWiZ8h0vn9
ibc++CYAFqAYtybgCbk/bQ9mblsbrpV8W6wwfn6nhaHDWP7TEMbA5Nx3PKRtpYtYGJqIqDLJdScg
Lc56a7/Ap/OdApvkv3Eg1FB61A8Ejv5pdTOpD62rsQGy2FB3u6zhxY1nnpY+P4snLJ26cI+0P+nk
2+w0vCOvAwRK1BPGU12ALvNsayd9ROvHOE7R0evZhSB0pnvgw+sk75XwP9zlffLkP4PCOUZPfScO
R0Cmb4Qi7wFguH6fF4lL0bpXAgQG47JmXACJ6VemxYzz9t4YvGIY3RmzvvgWX+fxzAakfyoQpp4T
YS4k3f8WR02cLJn/MQSYhmhSiA9C/lcSuD7MOQmKKNVqGbRHLzvplumcDPQYV6kNwXtfGY9BY29o
YNTCY1CE20u5Xq9XdsiVeB2GHXnWFrVBiOjH+1p4DagxKLldWBrvDQO7dmRkYOQxopUhlQtlP87J
Zuiuw+8yDDjT5wWDV62eLWI5IDq6o3GavX2N5NFwXxFUMky+5U0mHKUc97np2NtqpTEoJvsJ+XSu
BmpcJwIysSVAmz/Emj2Q7PArndlqPRYX0vb2SYErOJYAyI6zY8kr0QLe4Z03d0Eintr6ynocqW34
JCMuSBFAPwoNEc9y8YvljpUF9tNErBmqT202/u21co8bZWe8yCDETkiSglyqf18GTHwGSoOBHUkr
5h/SD0M/YDz2cEjX8z1yjxiYp99m6DXpA9q8XHnyFnRA7vgEEvG8vvX+Api6SEDDa9DJPfBbztzv
/eicJbvVQYP9vrueiK2swfnc4TZnaBNtz87kQqF2n9iqrFkWREXLtjblJAFCi4edqYGnMSeIrzKe
wELmsQ7xj9tXH2ZOwTooZ3cYM+S6Tsyb0Y91rnch8YzTFdVMTmgRnzaiIb6T+GptY0xGCZt1sTfr
HVjZlakkYldGUMqxhpumNl040DInpmWmbTqg/j5VKEGYAufprSgJ+ezwwQkt+wzHTOdGvWQMEUbF
ng9rH6XRpERBvbStqoHY5vIpiFV2Ae1/Wgqg4sYq3791P4ktKBvfd/DQZMyDFOhhLbveIxHtjHHJ
k3Y9d5CkbAlSbarRVmo/tjrxi0nSR9MPABys3SpXfXmKekclvllEP2bR1hCDQM/qCaGMdEWwuiBT
gR5UypRjjvBeLqXuenBkNtweDes6p/JpsKhwkIH3w+TdCW7CDz57oRurev9+Kze1DZc/0VCr2zRz
u6QwRW6ePDS5KWTjTgAuIkFK2F/Q1MfqzuceQl4o1yt7dDEQzYnjL9V9eUnFrpRS4si6oaoU9ajh
wtoOD7LE0aj3tUsn69g74sa+d0e/tYJ44f3hH8bUV0sL0C9pVgkb5EcvBCPr/nWL0AUhZw11WJZy
Nk5217FyvBB99coFNhxnJw2cTEuyhLNixzrz6FpXgTYJUxtFYw0Yw+Wp4HEyPXCBEjDTMz+Uw4IE
83FeAJeuNaCJlW/W8e0+Ug6ANn/kU4S4rkntR0Cn1FCKtJju17rjcNnY2c/THXh7b80Ax6A1o/HP
EmwTpLPXaZ6VDg+OfN61OGHZWO1gtg+kVaNO5ms6sPGdo2lmKRto48bIjP7OMafWtA6Vmee3XbWH
kgIJ1xO46dilntkWC8spyUla+aJTvlwEXRs5kCWKYzc/Qh5SueRkl4knZnPh4wH8qBLeNQb1wEZa
TvmUIGsm4lAXy75RkhtB8mQEfEwh8emnrq1ZoZMaMchlJl71WFUREopqhNex+/QlAAVUgu9bBUtC
RtaUbd23IMtO5Iiz1OrNbktvjHshd5NpTEMlIRQvqePJijw+j51talR96IwPzWgjAEgCbBgxE9Fw
IjBG6vCXi9Q0SZo39j5yN4n9LR2NabQolfI1WIlIbTQBrKYXPaOpGUtu4JzC0xrsqk/0YRXaw/G2
d2tov/T17+I55jINUugMxfHS/kdWJzI7Ntvj/aTotRHUxim5g1oyPQj3oKzsXoxfcT0EcnNdhqwg
1qENjNxao4yOW2uc05NmXIZNsIeV9Q7pPoq9KaXqRJmSfB8pTletJY0OYqmOPNK/hpr7JiD4xdS8
wk7IVUrzTTJy/7sNW7CNkyWwxmMMz6vMyEgV/l4efrY+zFdHlChohpn2GjUflgeYJ2F/raYXYbA4
mJR6jA90xm7ofUmuqqN4PIbNTzRB0UuukonT1S7NdhRThYcW8/NvJF3o/klCO65Mf9o6kocsNzOZ
pZkqakICa3Y1uCvexF1vKdp1/z7SMKz4xSaoyu/Dc476WOi7/hC74CbmqyPs0DYwBN5PAL3tgrCU
B3VEoAuxyhEXIr1+TnOl9v92T7vUm8HnyV1k84CGE4NE+rg92uKFhXSrez4BXkNQTvwwxemjvJ2t
KrvjYMFY/PvWVu/AD/EAbnrvVo/FYLmGR6GPoCmzRCHHx0Y7bQPIHQD/HahX4U5pjT5pYC+4bJp/
bMnfOvo98tdzeBEtgQGOindcY6Ve0BBL6K5NH/DH4DaJySOc2qt+MHeaQX05PHwr+FTtadsGIvX8
VQHbNSPun28PK4BIxiZ5EUx+r8TIOswa+lUZgsPzoGPYprt40RlH4PhgOAHij1n6v1sOqhd4/W01
LPIXCHfSBzfRjLw2JuhozF/3tKnMxNLRwzJ6xGpgjtdLgISmnAyi+8SiPvzLfeJNmSOrh78x3QW+
Lz5Bq3SKLf2+7MSxszq8L0RDYbQ9QU0rKaw2zwWJprbuwRTAvst8valoF8qztU8hmpBUhSdvMlHt
oY63h2/5ZywoQwKCcZxK6GEmXj/xh7xFMUtcOqhO5ZOK7t6DkQTp0DgepwG7MEbhknebhMa9m2ig
0SysLfYIwWSm2p2u6Elew6BJXJsaIuEylCkZrGWHHw+tZ9tEwIELw09bnKTatP1O1MIkKxP+l0F7
Q4iPq96aQ0y9gEXQRdSRG0NeLCSbaeWyFxsKR8RtF1MWfdvC/O+XaXi9ZudewEROOvo7+NzHs5ax
oNbnzpIN6naVQ0fK2qOkzS5u4qqOGnZQcL58juNsbeTXDCBIpRw4FLkw9LSxfOgzG1s4tm/7CLfx
Xw3npGM3ijwbBRdHGppnMesH3CZvNjwQueka3O1mPrgWxJXo5n3KxydazeVLFCQ0a4yhAaat6k9w
K3G7lYOld3wTPVamxmagJ9N7bsIOYbjP2nHOBMtq/D2QJkLoYdMnbcU+Vt+wtOl0znNNE8OQqnD0
nfPJxchqwy+FXjrYkMEzIoRe0kMyjqk+hiVSvMhAJNefx5r7/Uel2F6sGnJLigXHw7Vq3mmB1PXD
4Fgt2NJR5Upq6V1TAVRqlLck8E87yiRPrBghZzLGPMhfQUHzBYE4xvUYlVtYU2qGEZByrw0gERsV
jIUCZSZ5re0oqi5zhXi2rWuLHw9/dziVjiYHARJvAhnz84FOm4Ywm160ly6eb/0XISpy4zXBMOZa
GZweqgYj10uOxtesRq8dtcKOnfoTbmO+i1xY6J+XQb8C9b5xBqjt1lNkU3KsWFHRKoKvmijiNnfQ
6HqYP6H4Z27V5ny+TPLKW3wr44Jelx40f8769xmGP84aDLni384QNwDH6VmcAw3eiRF83WgKBYoQ
zoEHBBxX13Ma6pbutE/Nr5bIcJA9qKZ+CxIDtoef2nEcfv3WMmvJ4Q5bijBrFPeFy/AxK0kjSCp9
yXKMXQHeshNlR9q/+vT5w2pFbRxUIG2E1RhQ5bRSJxS6qBLmhW9AdKG/FORpVwJWMzguOI5Rq98K
BKzp1KxbA4v0Oa4YzhlSCGwEjtuAlPBh1iGiPwD71rz63Kmd4shWgbCrLUP/9V97h0K3rfAaInIf
eop2E/rQBSMPr2v/F3bWWqlv/SOtX5rp0RlpKuWVwRzxe7YSlU9fWMdTUf1SK69KK6asr5BtCxHu
4Hh9fdkzr8wOcvOfien4jiYo7+UuHKCPzJROs8FF+/Jy03r3bNpZmEKkwxqFMkqyVC8YkEeUT4Mi
bCxqbs6LSjBw3nLlIBlABhJC6W1KiBrge7wpPS1co/0YlV2vc4fKkFROs7LenIDAwf7rmE0th8kF
9Vs7niUaWZqq/KMB5+gyKI18kWZ4qZ10Q3wdzlbGdqHju5nYJhdEWfGEG5mQ65VD8pz6eSoGeEDh
cETPD3u068nZDlTZTApfSW5hUTG2NZJJTp0R3DaCeYk4B/y4qS10sE7BW+f5B6+wkBszf7Nrmk/f
z4VsEQtTQFY71cli08wthtRVRL1/kfPc0f07k4MWgwZ3QinhqunAAMXrH5gbx0Eb9Jf4fMoPzC+8
dx+BliWrwoW3e8CZAiLuLzc6+XNV1uvA/emJW//534DVkZ06tm4eSX6S7M+USokyQqlICXTC9YVy
lZsarJ4FMJKg//UUVcLqbNVAn3t9GRwJGvBYiEk7bE0g8WJj8xd+itE2EvvLkfh8HvtvWJSIqp6y
LG1+dW87+q58y2zncOEbskecDcIAES0qgDIUdw+Liy2YgyjEaFWyit8C+48rZ29mz/3YajaWdpnF
kuCreLMyj+K4HScObolngi4OeRabuvQTpg/kXnxzV5raN/lBR+TeUTPTxspy3EiMv3iyAnjfYOaW
ZRnru2F+e8Pk+gcImy5gxclWZTbqeIRb/umoVRsHms6bA5QzzTSlWTpXr+1kd7ZKBurYFrnNh5sb
8xj3CX9OGiVttXMox9ELRlEUaBHbLmT2zoEvcHVgTEkkB8QeE4Ag3n5N+HTiT5fa3xbgzUUmU4nB
lmeAYp93kxm9I9H7r1AFrN2BL710vHNw2SAs/+SJn7XOccJSQjrjyRcpH5aXiTOSxv4rCbX1Zw6c
fO4NvsOxTSg+lM4/8T4KOBqipoltqDn3EPT1acOdqXo0VC0BJ2VbdMkmWur1a2oJyfdtdqK/OZmS
zx/DJOrWxvCULKP4L10WiWhbbHEqWE1LMsm7pyJwUMD9yYSZ1NPeePw6BPFe2TfPgtY/vOJWQs9F
lZKydxP87dC48mKEc+UvjikVDWZGpyPjhdG4jtbBZicHh/x+AExTxoJnbJF8OIDn9bM/PX3J80Ds
k1n/zpe0iUz9rtS2NQqkd8Q/6M1lpdJm5Fhb2Eivd8VykAikAMn6fPDuFljLpeAKXokN3mZAJ0tm
gS07gbeZ111mn6LfCNZLpMmOuHmEjgfb6tHXfzWRoSmLEUTvQhM+sCytEzYlNBB+kfSTi9vDj9u5
qBCkV6VYE+zI72OfyFkBK4R49cY26wtQz1JCNKhR2Cn0zVl8oy+15959A+FS2wbssKAq7NrCyZmX
oS12Be9FJsLp3Q3DYZdhXgbKhLM1/meLeEh9jC9AYXgbCO0ejvbbPsX6HKyGo4l5RKEPnSaLTlgi
rQcdKsMHch1G72WYPy2oU1O5V5ZUn9uIWDDbt8043NfzCKOOU1cnn2ipeqIWyRWkKrjiB9SRR8gK
QT8obTxTy98HUa7CV8UAknqbCqztfvnKvtEDnVXNg+QwgK2Ak9m9l0GJQuHE3GPZk8sWTCWVvNx6
XHFfwD8TkyhaicOvtcGxgFBw2ECWfjMyEnA7BK9kVUDYuLSVQs7TwYHdlvF2JwrZl2CLKPE2/Sas
64NU0eW/05y8U+LOGVfXxWZ+8oyY3tPTC//Fw5gGkJEzXFiRijNEBEikdQKgk/RwJOVXDnfPhXpu
68wehLg7kzOAgeA7GYyalhQnfqDXNgpEGKO3nfC3mgIUvZj4WcVHVlaCcsNYs8ab9NL9FgBgJqbA
IJCoC9wXXhZW807DeQb0zFX+fYVFN2iXKr1x4Lh32WV/soAJH6reYiq9d7GoqwAacyK6dDvyDrlp
Yy0DRQEBgEyGnp3tqHjtvWcnQrcQJEwkb6B1x1cXENqqbjcNabaHzxqsJfs+vnFQcbnd1RoUG3T8
AQ/bztIIWXnid0mBFFwhkNkIfQmVwWX4OM1HqC9oKehMLk6lxVjKgGeda98OPHqmP+vlgWcBmCvo
AbARRGyHWUnNopmaEpp2tqp/ZXB5rKwMhxf2NeZTqLMtGLoGKg9fmHqMtnMp+7I58LTxRG4Xx9Q0
8VUplCvGxWu4s+U2bvPejcftJrtnzYGPtjfFSIHejjG51xggY+mV3MPXxzp8ZhFa+xBRZOMmL/9a
fd5EnA4/fs7/Hb2FAptXP1XHYwNBMNGh0unmZctivn2s8QILBQRg5KQ5o0s7HctTnM3ki1/FeEyi
/ICsXnOWL6swipad1Xz5e0hKdk4uUVQYVQSPqvbi2ZlefFn/2HMon+GVJgidfa9y3lIKUrZSJ93V
UM/PGB5iNrbeRVvqTbtWMVv/jp0JEAfMNKAyIfBrSeAfm7qmwgENPqWJ7M8HUULkFKAKH5g9liYG
fnb1He2Wv7ATX+lALkiRyzcx3UYUzG4mCZgm/VFvwAljSW/9MgoM5+LkwDOXLaSRRltBRKwQcP85
AbsDZV9ZzsxbFQ2X6+PmuIT9zhFBy0pl+nrN8sWhBRo4hZiLxd52AI3Olb4b8Hj6OMs0v4TdhmYj
FtDRIPyZ94gVH+eNli+GwR2+cm0RoTAf7CIpFNeOamHQ5oxo0FgbK4QpnSF9qZBmi1EtDJddfZf0
yrtHMAISwcUymr8eSG/yjKJMTdtmYhWXfDUC1V0cSozkfim709OFGZEyHSd+YkQEma9IrBVsV/Zy
OcXUx6ykIjhq2DIfwC6v1NFj969Y1gxFBbd+EShXHthzQQBUwOl+egeGMkE3GXXnM4Yc3HNHS1LC
S86piVZNqeLdOjmIxg79kPQRDt8h1idFNb6SfGFQAdYSmW8XVuqHDYz8VcAI/DYXEJU17JMUicab
kJBCJQCQzOYy5qkMYEFiKk5S2T42fxSEfj1euITKviMUbUifPhSlQFCGVLhKV+aRYNCvq5Lgw3uH
AzFZTiOZSV/4j2lMpynYrN6T/NL5AOMGvYR9f+GN70CgIOvEFLO9Dr+NSaR1OGYMtTq2XjxEamXv
rbSzZPWtslym+Hg/iEIPpDYQ8eI4afctr8IjYIpq7hNg9DN7/yjI0rnlgTjYfBgdSP/P1XKcljRk
93wtM5nWHKR2zMUGV8qSrZKKtiwUi5a/p7assaRNw/jYgjpTxQkmlvyHL+Iz6fRcAKJvSJtCNBZU
gSOZM8hlN9N1JXWOfs/YklF3sWelSNGO6spXDdHNM0RNKUdF3yHnwo61PBkL0Jzz6zaE4ZcvT7TP
CwLIALygurKkakf5a6RmbePT9MTvNNGjP0khRiwU74bwfZ5xCV1QrWNOWoN7y3x+Df0U+eNDWyjc
zQCn3JUaD2E4P+SX3a5n3Scb33U+wH4UHmfz9iTIIDh+BiDTjPo2bIUJdglQImZNpEMTtnL2o2Ju
lXcVeIbGSHxHJzUN/6g5bEndt4XfWaTvCkPin8X5oStR0C48PEVXN+5LMAS0M2ZmS50CqFcTLYMz
D6J7ozPwMwRNukBCy7i2xchwxkc6L4UNUy7eRszBJ2ZECgzy4yfXEwQonKUdAFEltsOqrY4zfTyP
PATWixgFuS5w5t29ExF7QfTLI/dxW+YUwh05mCpTQ000+VbzPJvPYqbmSqZ32FtOjsq1e3g+YyXs
eMiT/92vYvQfTEN0zvWhoRv9eTG1P3l9nTKgwQGj7YIdAaC50KcCGt5f5uzBidZxK0ogOaKVQyOg
NIP9dxU/ml/9oUYCsNyJDBvip9pMyEiP8o4kn6Et5gI4a7YGxyDuM3JSow3CGt7OokbcCwovEfOM
YIrkxEyRyjyh7W9wOAom6IvznMbrbfq9ksm5k+C5F4X8Ss+PRUPW/iRNboT+/AyrKzCVVdocS1K1
2zco7DSFT7cjJv23KKU9nHgTiCjktKBRgWA77ePEq0k/tdjK5vJ9dm5No4YG1QttImL4qPOi5YOR
PqEJbojjdcsZnyhFoWNXx/we3Gr+pc3sQ8fy8M1C+FVQdO3/4UlniVu5EVshtvXQW4HCekmH1A6Z
mInRjz7XtDWrF/0kxiPYcjTJcWrQR/HFZ7L//1eJsZX/ytqdMYgRv0ahsqy2yEF7e0XQP4fyG+bb
vlsuzvIfWwnXfn8u01I5aFpD0Z1x04yI+/xfKu+U8Yhmsci1hThDSmEJKa8P1MJqNMqaEBdgNZmI
oqaxcH/bJj42orYPzkIFEJW5v+WzWUgMN30mayiEaL31bzRgdPZZNVtJw+H4Fo5jclfZmy5o7Thk
SM9TaaxQ9RBEbk3kx5XqUExVIt9JPYl9RcYTZkle8lqx/sHcnnb0rRrMMVcYZloRqm9SeGO3oKYQ
lBPIQktB/EUll8WR5ZkJpkIbI4Lrep5MA7eUkEK4E9NefpXqnPMVjAqwhGUQj82Im0rru1kVmN4t
hQBJoLow4cXS73NR78OvcmsJr295fEawk0uDaX7m/jKpjg4pRMaDSu0OgepFndqIZtaUsy2eM1vK
QdriE5NH5y822yUTtE+m2WvmwR84rDx6DxRVRmZKADAGQaXBLm0tpO1GPDtc6QLBvvi0sRB4gUsW
ZUriJRlh23aUGBDL7iNHCBSap+NEefAeVEM0roHyalHo3I86th4hDXOmKaQUY2ZGobtjzGtWG3UQ
uxJrKOHKIWaaWHqhoXr/rDZPX4d3Kq7sYI6glfhx4GdAxObYFwvTuFzZwaOGld6rQWNJ4L1G/i3Z
oonTmgZ9hH8Rd7gGgMcVk+Nezf6eVlaHPre5vVESzDMLr+9t8n+4gzxSVRpX0aODr63+UJDh9U+E
iHAKBZkx0GlvB20IXT52PjQH0OriIxK80NG+EnVZPNMXAtSwMz1WYQLNcKWlAl0DNbSUdqd7x/aG
j8nl0tAxiOvFSGPsP7jSypbMcQaW5GHtiOc44mBFM+/9X/GkQU5QasApewfYtvPs1OXim3V/4QAG
D6+b2mD1CokptSVqGvL6pdczcI+35alwypJep4hvEYhN8lFP5vJDrwGEIImFXaPHPB8gxs0r9+Wn
uxprs7slrAnaK2oqdl422LQpq19obLehOfvmFS+LQNfQjH7jaO6zDwG4QqQ+oi9ON/yKrqyQbdLJ
S928Z6bVwlHcT1RTAZhl0CsgCo3DKD13ESVIgPoVmN9SO6BcgSAK2rF76g8bC+8GUO37EhkC4yIu
8ND8vJ3W7FpmoRdKYsJjcVtYM6pY3iGumIbiKmxYRO9uTSaZGKfylQrFm0W8jfEH1MS4pny47dqP
e9kEjQiGpPVDKv1w16WP/WaM+XciikX24/oM70AkzEYAbNI4mRieM3YzVs/w23STpgp4wviWN6Fw
OgkK3paBVdYUOLneXvzbPElqo+WPcSxLUUGj/FblA/fh+JzZkA5A/v/hJeOxO1V866QoPWxdBMTV
7xwmjBGWHnEdF5cs66MwzbAQDKDIbvnvVC8Cg6vlmxjcQVeybPMjmhkuV0fPcenXAeMWEhboDFPM
aBEZyrSfiGmwmOxpepRhqWv4vmQXtU5B+FHgsbPGuqn8OkrsjPCy0Towm0r47By5IvOfWqhz6Vf2
nohs4XpPDJBWPRzsSBtBemNAO1dBgfPLFWB6mTGGWQB5H+NCCoh7FojWyiznuHf3BG2xM+/pVOwk
upcz/a9mVDd/EpE6ythszQLNiL/Kl8h2vzHnkvK1VCVT+m3apkKycrD6Co/MvZ/TORAct3f8y++x
xvMTHVXguVloI7aigXhdS9I+jKBPFQj9d/Vs6DcjVEj9lAEhWv06IwAA4duy6uUx1vXjRlok9K6u
Wx5Gz79bZiSvL76jf0mYa496JCxk6TWxV0p0dwBOBhnL3hpdZ+fBseMbeYbplzSNZopIO4pI/Zk7
Ps7RrL3MU/Gig8EuTK33ykJovvOjGovtRKydCkIMZ56hbCpdoC8nxJH2fWGHKA9un0eddgu1CsqV
4TQz8yUjL/2dmZBRJ49aVRvt2HwIbZUGPz+60mtsGaAJ041K68LufEZ+xRyhzFLLecQCcAcKgVBx
P5i3yFAU+SQs/wRPfLiGP9gsctNyyWB6VdCQie+XPhk4uvgP2Q/6GF9gPfmYBwa/jWba/j+upb3L
I/bQuogM2ACicZkkm4xlmkwSehSbDXHMn1Lj91kSd9IAtVN7U52/jMkgDn+mkV5DKnvpqdiHCVqL
t1ZLIAvlv0vdBR9lp74HdTSy6DxTX2HsrkcXQHIHsetH6XFKSygcRgzccMX0kFsnAhTEzd6HsQb9
FAg3QsXUb7LVKaCRTYR9lOqjorGoiVMsW6VfoLxLEw2l/CpVYCXqYCilVeNzB8QE/OhmVqJpgULL
flMn6LIGqO6K2809lSTZyLgwnrBF6S/5WQTMgcN6M14sI8sXx6oSLOeanokBe7xtD7cW2QMRtHIj
YKsDgreW0/+AeIph3tVQj9BcpM7O6gjP/h1DfZ7MbzvLBBAna93iKNRbuUtYVEPDbjLJIgPwviqW
SPIEXnrjsjXyXIWPBdnTTMkindWwcsq/GEwauBu8EOn/ARfaKTh4jW1DVtqv0lte5rLcwORMdJUe
WFz3M9ZCkf/2FkQQvmFhQDVMdJSvobh5/csJMCQh0bU2VVkSG7rQxUVjFrGELHWzW3EkMIPaAf5A
YyztCmG6x7j1moDwH65tdgzWJBOEwNKg7nSY0PhIIKtIY9k4WOIHvhCGd6r6sw2RywDxsRNZ3l+b
8xAXKomJsQLth6BkxXYdV/UsRYpziRdLkSLisVpdBBqNZdS0yTSFR58Y8iNIkkMlbgwfvU8zSMkr
AA66V2NGe6Ll40Qrfliaw+0xtkDACaTRqXK6atJlpJglhGJaOMlR7FPPIXvRskJAIxaZt7p6/3sj
QbKZy3H5O7JdaxRpbpBjX4klnXQfT+RBir6Ey1NG9lxvvfS3huMcuPe7/1ATeLtKt5PUNxeWQfdE
JbGlPdvpvugdSfApYCfbfXLF0lDslHP0ul37aWY83T0JlBx+bbF4kQ6fe7HhyEmL7RDRiN4BKj67
Rek7fS8UUbDU05maQdg2tsXh7MyOv3YLQnqgQbQnQsm6ZpN0apFX9yZXoDgz7ZELnwclz1ZY8MW4
atlYYZDUZZlhNTOFLwMQ4SdROfYuMfU3gaKCy75KMbQJ6jcr0Kga4PgGu+RxblYGPgTQ2gZ0ZOK7
7oM9UeREj5N2uqArsme3xky3/prH+ZTBYb9JHn135iGXXAdCzSSbe/f3p5hXJ7ClQbWmLSPkqBpA
wVRQHpEgI3CSmdD4zFjTTt6ReEQ5iea1WJ7dChLOH2HiHiwICiQVP238hgALVhE7lAGdibETNQXr
jWKzaG0+Wc7hKv0YYl2RpZV05eJQB+137jNGbEJsTBN/pRmmk4yVXKBZ9tak+KhTfURBicKh0k0j
Wt/uTmDvxMocebxU91nErhIAed1BVHGd2OI0c28S8aCY2a+GEl188PC1genrGN1gIPMksJj8DNgx
NAv7Ww28tAXwNb8Rr0PONWxxrBM4geXPcRbKqyJCZweo2E9U6i6ckvYO13S+aEd4liGPSBB9mdX4
atMRt5DuDGXqkyHeH6lfqljuxe2pXuERZlT7yfPIeQYaKG62JJH7U2P1K8sg9wA+HUB4Q1OI2hv0
U3Kl6Bp/2xyYvSarUyECdg8pEe9v8NNzgtXKnV1j2zf3QtgKtdm5tjovmgcBZX7q7bLTjJ8MWcTn
SZmZTKrwpYFgQtgcl4AxYL7oaXEY8Bq4Junwl67VzCxtSPPeJlGGiu0t6e8dsXewyq7LKIK7xUSO
P4pTkrk4FZAZZSymohMQFI7eQNIZs8gR9N1mEvtyf9NeqGfTDsSdmBoMxAJyxVmRP07VwsU8vhE5
+HTKPMmyR1RzKmHY3Ran29JMBH4xO3Z7QUOwT0/e6IsDIIjHMUMhx9xlYQqPbsiP2e+UP28EXZQO
t1LVi90EKxOjNRbZ76CfzmTBSfDnz5K09Dk3hAMKk8F/gaYkQyfV+wxpSWv0OFMq8xGxqruf0pv0
AzE0Xh7QFaBFbZK0zJG6/Th3UY3ZtM5Y9z1BKUd6mIb4J29cm/082MnI6b9BJ34qdZuAn8tXO0mo
GxZc5QSdNoEMTDeYuHh2V6JxniRbSuOsv2ft54WBN+nYuWDoI3yp3wCP7sC3OvkqoIJsdVwgsU63
O7r64VLqyj+5an/mVh82ZKJ2zeW14loCn/5QmH/jNFBNi0sxtdQ9FM3qH2IG5RxywuysPz0jhGIf
kUkcmqm/xIIPOmYfCXX7KyVJkJqB+JHcc8/ykugc1MJKirGC++rgFJbx3EHqLywuH9FS5BdO9vDt
HGR4q01dDzk47vGCwsd6Em13r0ifOtuZ8Q9/jp0BDa5vl/jvhPuNKgsFHU0Rj1QxR4y5jkvdLtj0
LywRyuV0dTvcT0ZR/YRq75oULjP9qxtG3mHSo4Elq1MnO5wIcG3ZGctlTmm8OY87vMXtsQ7jzfrT
tu8PYj9Syv9AAzqnyDhkQm/G8wg+Tv+aMyfesZNmtdX2ElaVWFyK1UBVhvJQTuFP5xdkdNA7h4Ki
IkKJSYr4Oe0bXcUNU2JexrwZ1EwY9xMtOraQGH1xTNxGOTiDZCdoXdnKe45MEeo5E1g2/OJ9RkKS
vfmaUZ6b25wIUBpJ1JYovbRM6PIakyi99EH65YowIo+Y/D/g2onySmNuEKsdl5rDhiOj5KoWos0I
LgR39i+2WnahXDnpSW8K4kZ4uj1p7S7HsF/DT3CTCremPWBPK3XBpPYqlURInIqjE1LNu5t5QG/o
fDdpTIXzPz2AIqiH/qTMDy6Sd7EEU+g8myrp/+fBdUROFHRmhjiZQ4UTxNVdGDG+XN11cqwAgcfX
FJljq5rxWpKja5QauePtAjQgsz4HQtPRZkH6EkxFrcFCeIXTtiv2sYPY3n5iolkB8HWr2kNl0UBN
8TQcA8lkPiJsbd3bbH0LBPn+vA9fi41YO6S7ApqjeqdPIGC5qAzfhP8Ju3Tc68xa//I3dWoQyaik
aop2ux41Mrp33f5h5p6ujWAN7exlqZdnaqrONj+C0ThrHfueInJokYR50eO65HUG4GjSfAJoyRPo
WhYFRBDaTflMk+g/6V0eS86yjRTfk1W7VMHNlHaNI6CDenx6IHTnl6ejf/zhFNqcsemku3K+lK5Q
5IhpHyVuJBAmtJvky0ms36G7C9yBMq20CODEzawYrNHtT3vC6juUryXMJU0GjUVsET0BfP1LJBWA
BVw9smOBfgcye25KoY2vFAendIyORCyz8D8RwAsXCbXfSG5ZhCbi234PknqrLmcUW0YNvqEn3BGR
kvbIzmYPiVg5JxvIK07ZyGCeCFKHhcYWbu8BbIG0br8GGZFvL4L9maZuFgOrtNvuGdd21BjsBRlG
u5H8C7o+L559yDmh6r0ZhWeIp301XQNTwKWYngPLu6V5htd81q0vTHpuJ/HQUeGEbytcF8yfn6M/
g4MpUNXQyxomn6Bgk2ghHL6bLC7BIiWUNgSu3Bk7QpgPdU13DeCrKDcfcf6EmH1r20J+IwJN96G/
G4lkiIIhRuBnfZ1tHfowMC6SgSFiiMlQHRzD20cbAFCmeQcmfYIKbf0HXkOv5KwV7L6hLAQ7xgEP
yOEWCWBXMuATZyAANS701aY+qdJN0+//h/CcSFw6erq/8aEfmgCq/1sDSi8neuY/Uxt+TWe4aWAn
fwga5nKnqRumaV/eMRTHZbOn2bvIxnTeQCcsv4QVEwdbfxdZgiwzsG1RY5LohHmeM2pB6ix2m96n
u2/uoNE27wxQ7OpWfaraBtZgRypxfiI3nfy86crZZFiR/8bGQxqyp+DqD067xdzGdWRdDsbsAYmW
u9RGrA3MzPribhltjjKWzyLE5Da0n7+zT5plhCAeIuj+kiFt3MJI6Ik5aQXfanmyC8X+u4Bu6rep
SVur0DxYU+zyElK54kxx/ogRrEG/UqEcYR+ZHTaM0mIBZyW0lfcskFf28abHBOqj3NTUpSOXX+fv
/z8t/D6/n5nIVT0XWO6Fqbo+F1sp529Si1cPx3AmY34rVp2/I4rs7buBFf0EqzK/Vj/y/2b+bx3s
PXbsrYoiVeW3z5QG+Z0tiwoya6qvn3sFfnYJAQLpapTgd20EuS8JRm3C6XNmwBE6Y6XBB8nWpAAg
SvVfaMa6B3WLc6h7ui0bVCRincui02uBVU4PWM1tH4/z0mWQ09d19LD0f13YuuXWnRu9TXQF9NFD
xQdOdgzJcWRYLVhrxU7Ag/zwePoeUNW0EX2VMWP3BIX8FwOFUvM8LzHzKmOpU427vOh6GQ3pDixp
59UDWsVZ0WRIHkTD3qmRu7ihg/t/XxF+mXHZhijWtDf3wTKIhaqxzdl53hrQOZiyffXWpWLJHhC+
F/p3C/IFbCJIx8N8ooJLxR42joXpVSYZ3VJ12FBqKgx8QK/xP/4z/WYmXPu645zKCf09Jnl5Q8iV
AEIBF6DToDmIoJcTLWt+/SgmMHJh0CNxliXPeUQWyvsmcDHbooY+T8JSj6TcdYfq0fgKmDKqWM0N
0qYOCWjhhZ71mmoMGZoi1XorgClD1HlYw833uKpaiy6xgIgeKpL/c8xnQHHj3jT/XavVj+kXt9CZ
TLFJYlT849TNgCdgPGZovloTkJdxf0lLRx9R9yUSL30uGbh589xrOuwfnPekFd3b9SRazuTCzT3x
qGBtFhhGJBtLp9eR+5UQe8cldBN4pAPSX+ynMFgYijY/Ad+i9pClX0jf9eiX+59awJ/BEfD2FdEf
OTEX0C6j8NLUO8Rsl7OzlTf+5kAvSEP92fPrePOfAEGFQOyB+RTjMT1JJTeiKBv5YpFWagr1RzQJ
9thyijoVOTcVwU8X6UzkWX1ihImCd9PJU8ud45PnWJLjIkeBkFw29mSf7pfr0qFe+l9tKts/9aTF
wHa2h6itRErskmofd+DIiu7S2yocQvwiTPi6usO519it/TxX0bNqVvCIY5kk2xO8Z0mqCmWsUUOK
RFJLqOt/vw70qR9ryjHLbALP1guoA7WNZ98hOaMC23CFS4/nVd7L4mPQJyYctO9gVYvvrPgKOt7J
Hnsdj6WCgD1qPcDuvt+SYI81Jndv3II+D8zH2m5ZfRPyJt6CYwuTE4E+n9IRLSt7tAvTHQRLH4B8
5f1yTADbYgJV/ZmARhJIcXDHj5qBr9cjm+xo+Av0Ik7EAYuyY9sQTsPOiZzdxeYd2yIXSeOXLkwd
Q5BfXP4CngJEwx7ISoWp/1aQ4hmGLyaiHbLGi+1uofPK8DjCn+TEnyQse/5NzfRMPL//7FuBUFKR
X6klTKPxdSfiv32jN+lE1NKY7ERAT+vvzdYqedrVEpcIOiAqGMWGUyOin1ZF/QFDSt88vccdEuXg
+k9qMsSdV5nDjC6o0R93Cii1b+7hbDLyW6XyeJIb+f//ND1Ea7nSGpm28PJo0WeQVGVN0g0GIFh7
eLZ7Sw2BknRj19ttq3euKvVZwMNP28cdkHXn2cGNMkKldNTZhf2u48kwPgW+JNDR1CnaHQc9Hvkh
jUPE9jm3aruZYJGHKA9ELK3ffwLco1dkgb6UIAmOSaI7QE6+6FwCyKGsmeWxP0bRl5E2CfenAlYA
b+Iq1FAB385O68DKglBuJthfNFonajimGEG0CVrd09gUjInC4wUzJcRm8riQAsuqaTgj3xsiE52U
SXQuybInSBhk2IUHHcf5mJDUsue0VKXNZuK8uHqqiwG7g1eH31vIhKBRHfpXD91T1JArF5ASK7NL
AQ8T+vSDA/AqDModCXbs5QoAUMQ9C2ILGHKVbi5s/JH5czrGzRbkerheZ1my1bE3Cw5mQ2xoTWD2
PVvHRDVGvab9OB5ydmfDZcTGljd9hV4sDhEuBhzMQjwpTwfNRZslbrRcghzMavqn10mi+btH1xpX
rJuKtd6Cj1eorEKmupy6+jL5zt684BVgaUIctLd5e7XQx/7kYSimE9IF33gn6QUURA8XHChNSFux
7vsRfRhuGtu09QvxMJbJnYoaOvm7WiWs3f/5JJYh2smF+HxVBrFjtBnpmZOpP+lTersZnHRHR73j
AuCHrYgatBIK+36bGO0i/7EB/kV67jFBLCEmqTnCA81Ws/8wwLVcPFmW1Ig+vaR89xx8e/hhSQHt
CJ5MEsMDSYG4fLPC1u7TDaXRkUDrKh5lMdrz2RsZM5sZwj90HuSLLyewUHI+gFPghbRs3t+zKam8
Oo4qk4GDPnNU67TuLglhsWLn+VZDtRwuc0UooN6XunyGzaMxVptOcBoLKU4prUESK5b3gQHFHMq9
G5JYwK43mwqbsCjjGTocoRTnqc9Y5T/9XRZGc79mGYDJNJKVgl06UZhuzDe5c1eHzT7B6sGLR52M
fKR5FIYT3nni9z/wkf7zJGBFmzSAo0+3FHfWb7Qxs4F6Zx+BA8msOY/lHdM/kXF3G7tARavDJlxv
FJGHA+HfgTGLYw1/7DZSg+WvYTA2sT2gm9vi+JS+GEhJJ3H049CmQhohSzXe9iURGMYfmQPanBlx
tZLI2C2DnP1l7+5sP9lo/qkJT6h7kBLi2cvBfYwP/c1R9tphn0oujA5hG9erpeENhOYtxTSB/19G
ufdvtO5oLp8Hel5pkJfQO+T8liyHtt58hsSvv+PWKPzaPnrmRfEQEalVKGerTQdbVMF7SpSR+w/X
69OFpb99jYYTBax+/V/+xKMYFo7C2edQ3Cw58fVCL8oe4y9qWbSBM4aMItc//LhX8s60ogKNqx3P
PIuJ+/d3mr+tZp92I10gqqOZ+gnI1PKPXnx0ZGteczj8YLKz6SlR6tOYdW8BfZBzH2yLac1/j1Aq
iaQdv+G8ynE6oz1d6BiMJ5YqxBCQObQOIDFWk2tQYwepcg0psmFhSS2Hn3EIgk0zdHcFKTZsx6p+
uSH5RjFqkSQo5ytfnVdWYwcHWF1+vSDOW9pA7bf0NVOXgULAWDVPPd59yA0cP0uVdA2jpU5x1uL4
8EeGSiBoxTiu1er0cGR9+iZgla13fOmdekQkB8TnSyhycIy08NUhDgYU7D04to/k4MSRR3y3gMYm
zs+oT+VCrX7OjWbVWmlGhv/Chz7dJIOKkLhvr6X6vorWbkkPtCmUFgEaSAb5hwvZH4pCac2Mzjps
roDw6k+ZjJbI3Yl+GklouHJLk/+YJ+8cQgH9ungOdA19EI/W+Rr1ok/snfSTfuXJ1DYKrbD7Jc8X
9048zSt8hPj2y8U7bX/l6cDcPr3abzGycDe8S7Q6WV4l1sa7NMuDAuutiirpw/UOI0zlrq/wlUFC
Coowrn6mikNYGdl3zXA8Bx1zyDJN3KB9oWau/V2vEyh3StfEdX3rpdrRzmeQ82h2dMDMn9zDT3pY
v5Cv+Wqi3DVKyLNMTyNPpb/qNxgXstnjKy/5wfX6fCztjJ9XzNDSJgustSfykkj12qQWUBW1WHdi
Y7Oiv9xVorFzRnXi+T7noW+dtoc/QEmEqyn2rd6mYuVC4hsxc0VSGxN0yauPdA+MvNsYRZAsjagc
AuAAzT5jwcgpNfx/InvitY/7EIn1jEUK2yusPByrZMSnzDDiLDA+TxZdevfybveOth2vs0fS+MgW
zWL2Nt8ueNp5Jf+QVbWjtVOQE+7/63bJ5frHXZ89fs+WGiEGU7BJzFhP8vwvwOKZO1hzUwzRw5tl
cK/VGmUq9/Ge8q1InSAMIeXSrlrVVL/VMu8N22CxZHuqo4yhODeImdQk37uGSlfVPtWfTf7xs5AE
xa99PzsHGnWmSkz4EWGdddHhPdVA0e1jU2sXD+B2cJ3QH7bQxE1Z3L3Hbmy9ylrv8ZdiihFt2SWC
5WHlb07NBTVo6K/7PW2qmfm9Jx/OCtSM+htMGwAah9lpiAIg76i+9FDLRUppiEFf2K+U0qqmaIJ6
/N6gsmYHc0E5brAUAc9HnmYT7dff4UHnxkmYxG3hpdIddMAdna4sZaOHYuSjVzAb8eBGGNSGsAsf
8awWTqwPaLXzXN3xo57XbG9M84otoupenVbF4SHSP7QN3DoN/4r3IsYqHVQas9ChrjW4StXubm37
MMPwXt+v+794cF+nW+0cCAwBRvt+K3dBXHaC+kKzF6bW//sD0ESsr1EUpLEwQNjYk0zvD4J7bZKb
1tLNLKYVopCw5CyQ4hTDmoteTPSlg3/+EQCdd76KCKY6SMU6ugnPKvr24nNGG20gJeH3JO0Hadqb
KDTfL8ViVym08g9gVqB47Phf3b00id91WrNToIglx0RzFCoF/wuIwuo1ZaMRu3jtdpdc1tCXWqs+
ipVyxKP9n23FMonKbkn00Ji4VDa/X6mgQqJwImvlIvbeg4Wis1SNdSD3S/Te6EJxc5keMWpzEuos
lBdv2JUxDWJl/Swd3obiyKX+ogCqSPLTPiGxj2FAC94U0ENQHxSZUs0+dqJdT4/k7LCcsEvmqo0q
6Yv6l8xI6Rl3MHHLMohB/f4bLCCeP9ACzlHd57Y7nCLNrPK1u+PgkNvWy2ErPNdUS9JfRR5dmBHc
qgJFLOm3pOhFLTbCqdLdGRVhDdVdvlHEIv/H1LP64Ck/PGmZKJlr7xb/4n8whzP0UyYShMJ7sABI
rK97+axYs63twmq9tR222c2uzIWFL/Yy0IsvqR9LiutKuvtJ9ppM8PMaUxN8gtcpt0ygIVRAOjDK
Nfm8W2iiof1JJECzQx1TMH+cuQQgBLu+Dqp74ymbNMvCU1pQscGbbyaTw58OjdphAIz0rvIOoD9L
H34nyKwabzJsxciHSS4oVurpGvJ7a+xVWtkBhH5BkGAJNpJXcbfML9Xj+om6bhzGvWkwd3MaYgk5
2HzyG5/OwPjeW/8LLk6E4zKJDhjue3GD4zW+bf2bJd6SN0jhUBFhPvJ+TIPTbO2Gx73AoSu0FjWw
vaE/ZK6ohs5GeWu8SWcaSsOubtHmFKL5dwHRMlugC+C7/sgAKFGPe3bnsQgm9dtvj3W67CB6LFaH
/oySbL5SmEKxbR0MXhIrZc5lbopLmubKqsAdjkp8zr+W8oeSg1qoYCSUMi611exzKkJs2DeqQSDy
Pzxe6IQfd9kgDRQB/SAJcQEC9HRHbuglsOsD7ahC2bNi/5MA42OanovkWm/tKlKiRF7Qu6+i2oop
l7ym3TpnEsCeeD85PeeTMeXHbEdCacb8QoNFvaMSWW+k18zg+v2Ncg3HSAnjWxjy9cNwQhCIfIjU
hPTmTcxwfqk7rhtrxoiTY5q5+1C4WmKgsC/A1yz911sjK8fT7REGgtmZke9sTSGPHxdJP0gFXQfd
4aYjb4Eiyxh4XtYHML23oQA8zL9gZqLc8UHURGy+ScWy7NsiqJ7rv8mhXckPabdog4tKsRLFVPoX
GV1i1tdf8Nbf3T+jGhGXITSyObjWAd+mLJ6XVW9XyI7Q9rr5JcADES5KQGNllEeDDKsrS1CcHlZx
Q7pUUVEMpzQt+GpLYfaUrhBWUnmYsM+n1K+B3ns3abxny3aOwu5/i7VL2BR2LeaZ4ESEjHa/Swum
kbzKZCBCUoD3z6I9SNJCeAW56dDJpyD098ih/ljrUjAzq0cElUaJbSn1a1ht+rJ9YG+3JS7vEqU6
QNx/aSQO8QNQEpP6n8TZYBpcV/9XxcRHxnEy9jVEapSKp9d4YxJVBMgqQut26FLxheTQZs+GONQB
YkfbxPrf8/XRfAzEAKF4IFTfXXVL9iI/fZJwUEZfRmUhgi5FADHapnD3AVXS0U75IpTRDYkUCsrx
PADy7SuYLniRrli/RvAv3trrp3eXWgkjsznmqg5eU+SFc23MFN7zN5li+x1Fi5SBUlB5Hg+GMDhQ
aIw1f2v8NdN/pTp01GaGvCVDhe1BPfYO2qnCYDnhHSJH6PPSlpNckucc5jrzkkyKUGWIbk7RI5eG
fRWgWUMzo2m14Pczc2NlUljDMHeumU8Q2zAobkhyzUV/CGaIRCCnlLEgKd0mrQ9cv6AmZmh84HZ4
+mNliCniNMGa+zXFtbNv9acNcVxYcgjIZN7BS9kX3Bd314W17MN793oyjVKo3GXM5dOXiMbVKqkJ
1xFgkiFr3NwkU5w18sDe34EmfkmAbTIcWqudsFqdcHAR1I/9Voe0F2Yb1czdEEtrv+3sOzVXfQjF
ieZEVB+hwtJigO6MEUFFfYCTSLQmJrHR7Ct4+OEO3oLVDbCvsAgmZIquOoZs1XDMU0LiHr6muIeF
mfNwCCbr6gLtXTkMfJoq3iCM198FPudiZA7jfFezCgcFzzzf+nvZakkvj3D71F/BbQGgQ5EXt1Rg
3qKUUeLAtg5PK2lgtN/5vw62lY0FAKjb2sgiqPhyby9pTTmUPVBkkWDV0xT4HhCRDOgga+vei5t/
IARHvtfhEhFvaAdPtKK0Xv9vSzMPQTQu53V5eIITv3Uca0cWk9Jlq0/Hc9fomWeQ5PDEzw2A+i1W
aJYzU+P3chUXvZ+KeC1GQwAxolc08/N2nEF38hh7T4Hm2T7YN0kajmiRayqX+cqwvUgpn+ItiBhE
Hlozz3Sb4IKy6QcX7gyA2EDHG71VBAmCRSdNnLno1yIgZsOe+QgzvL7EBhiPEI8cq8jlaPZvgPVP
5Yj9PpqtR0h3G9O9faNHj1SKJg1DBcFx+b4pKFONhAaAb7TokSD7j9L0RvA00OczGBPw0akpDX9G
GBWRgecgUGhpMOak0Krwzf6PpE6+Jvvx+11SfuxrJEveRlJ6qjbN39QTS9/T9q5UhSc2a3J3IeEc
N7pU9NeFCYbRlJE5vhf51hHHPvwC+FIdz0Dy3QQdwWc12DslP/knthyCs7Ucd2y2bpNmJT0yRDmF
NzDJFjWhwvLPdQ3wdLFGxQidauwoqJv287KY1u1WJjhcMD93QbtVFmbYUSazkOx2tZbmL9ZtqLfP
wDKaON1spsdr7a6Ikut5jtMou/CJZsQNHX1IkpyoZjxrz9sKvVF8GozZiEnkCdD4okcoxyZ7mr57
gVaBlg0SeGl/hvXCDyNBqqYiYSb8I7shEPxLxbLn3nztPInV4lgHHgujHvUW5+fvEHlX2h7ZgsTR
9twnmZ7bx0qIdQJK4LSclxRE84T7UE0gWRFpDI/EkeCcAHNXA4G/RRMsIdY5MzAFFZ0q5MKYjMcl
2+0Ts0o01BwucKAtv9d9dyBX3azXEvGxrdFFPmxXnQmwIcPfpyljDcPkOL90Ay2b/Z8HDw1A3JaN
7av+PTq9nwZjdvz+WyxJPiPWWsQ9+D7nl2fw+p3yi72aLCX6WC8+1oCUS1X8nnz6vJf0ex02aPI8
Tj+xAN/PnBfapp93/4UGF7x1ULmHHFEMNIFDBpGOkgthVwKtflRKeKUzXWHHXD3jFhtJYhSbi2V4
4hYVpKQFicO1H0NGl6b98LXNKk8j70g3AVn4TNLXBRz4v9t8nap8mSNoWhS1EewQ3ZEGIQNd2tai
4F3+6eOWUADZ34oQs8ggd405HZ1yZKhBKLCD3w4htK+yBG+HfjIxY4rIs+gBBONacqBw9IYVFmFa
7o5M+pmGJaNkG5ucyx3O6HKJly/2UKJFGEMYOjMsB9yngOtBpX/Ut26/17qhGrF8p0slpei8STnm
hydzBBxwiC1PdTWcKe9FBIU5lz/Bn8bjuU0bunmpgm5w6AMmQbN8BicNPng04hjHkOnnR9OzueZU
IwbXo9lcHseovsRyhVIy6IiLXsPsGxkiY6NcjO/1QY0Yzldbu26tzf6eTaADFlVv7zTUHAj4gzmd
AH3n/69qz5pm3DOphsxJGNTFF1n2ZvepCPJriOptFhWFWmo9Zh589Fiqt/VhqJ1km2xEKNIibiM9
I7RSK5wYvwr9RjmknvqH3hk0YbHn6e4rJPwskH7lMgOzGgQ5aK8ZHArDOMQiEm/CDcwsM9oGLgSY
wTyUaMlKwwRLWCJIbK5cc4z95vVCj5BE+xw+MWbU7VYJNtXKSQAY1j1D8KqTFKldnja8dZCRmbPG
kqVjBlaMoCkNtg+sAcOT6yA6NkC2fQBg+f41z0M6whzWQp+Y9pgw46jIPaRaLkIf948sxRzsd6NQ
TmdkEtVlUpZGKf2xUsGDGPevv6O+JORtbMN0xAuVQGK6W0wRxSlyk1GpAV41EbEMc75BYP4XAnR8
DOvSYR0YpHpNH3p1UK0+S3sFE6HiUq23mXyXBXWgSTC1l19nB4cOJml6yArQHc+BlKJLBBov1bvx
D3GE5isFtg6m7/g/0QP2kV5iEOP8BUp+q5lBwUmYcNB5izHqkj7/HaWf8EQDF7KIx5JW+d8zUdpP
234B1a/Kt0tO6mrgDxvyqz0qFQOBmlpBXCAz4PQZ+fyhi0zi/IDmA1t/w624adRw8xCDA8n1lbKB
AvLFYAFYxlJQIj8zEt9xrHBkj6fwRn+OpbKFvBxyWQ392lp4+hc/oCRoH9BR2RZAwdaPyOvUrG6O
LODVSEbf+571NsSmAlNrINYz1LlEb6k6W7DIO9fjwfEMVJEeV/Y/IRCQE8STEb0yn9GhRbx/izhj
eFUOD8tnTAlTyUAygUtuA0uHf56n2QOV60dkV8d8jUrO26MXqiyB9G3T/U/FNoRcKNhJZ98A+nv8
ld/4NlxU+A93RGHTI+pTPGw67+oHi0bqHujI4igGVOzNmj4U/JxGDiCYT+jND1Ac9TKDdHvLFt3h
KM+t51fbh80awPnrqx+JpB9dpclCw77qjEASNKmJ94KlKr5eU8oe7WCc4d4KBi7T1ICk3U7zVVd3
O606r2LROV2WLzL108kDDgkNIzfoFGBV9yDcEmHqPOwpz71WQ9nDYv9jXcoKrTCZuABgYLwnIxi7
wEa0jfsgtYleWcANZPAGNNYH0afvYuCM/9RNBw5iYflDq2J5v35/OCD2OO5GmjgHofKSI2ezZvj3
7hdGUO5yGdHUYvNNOo396jylTF9pTkMOQTfe5G2fd3MAyunOVXO53z2bLBWbzTXOM8WLEEbES1GJ
7aKJqS54h94SOu85oYHE+UwLNAiCM7J8xa77OZsuFg6ODKRtfcR1/Kr2s3BG0anM5LMU53YFTBZ5
fnr3pr4vIbFHII1JqrWzIIOWVtEguO++WzXL+BiFFZC7vUz6kT9mBxrXq/0xFWL+CuzlGjHFWeD9
gtJpOF3BqX49JAsQJLHmZGv47KwTwbrNeFmhH4ayyVxJkAVN6gVI6kjYS7VKD9id8h98f4X3fmZw
S3LWk/6BJZHhBgPSmCX08t4yL3GGbwr7KA3/aBiW+YYV8Zs46gJZz+GtFLVxp02OBTlTAaB2YjOf
Jxhtv7y+vQlZGoHwn4str3oW/8dUf3W19pvSnLeapgtQ/F4+g6JZ0ct80ZjK4ssdtOtF8SAvsjnd
Kz1FZjTrr+JUgtcgKvZczqQX8wBJhh9R72a17o3yXVbq9EVplxWJoIudVL2JDuHY6D5tes8pmtJy
XVCBt+pklJKf08xbNH14XIY6KV7RktN8CB9cxyDpzv2xcrob5ylFX+QHOLyWb3hYsR/6/iEEOrVU
FP+i5AoX752Uhu8vMzkIOIMM80yBf5yegFiPx1Jo9V8uTi5urqGvquiOCqa/+GWsXttb/VD66N7D
8qdTLdyuRZ2zwGphqiytOO5yvTi0a/1vQL+ilmWWAt1ks0p+Sploy3OsOqro0+eOhK4rYMGmnKwr
0Ny7FYO+m9tqBhNy6jjpbHleFSQ9nRh5s1n4ghvCYbK9sKONIKVGShv5hbd0LV0UFEkeZ9IkSyTe
nH+fRWDlbHZevgkAQ1XDu8lpSMpAD4ZjCryQuluyn3o6AeNKPhKmeBXKbFGApwJCbGN7kG5IP5M8
zdaz1zdwFSCNT8khWamuMJQdbo0Ef9UQKBu0mfam9AD4oMJJgT0oR+Dqp5zGTcnMNUcAhsFoPR/b
OjVrw8y0lat67L1U4YOl4ktv5rgcjCyM1rMpZaZo6b1qxiHr1mhg7Y4Z7qku76d7KYIZAnCndptA
VxF1BTTTzqe1hjXrmFb5q1fvaG6XXPwGOOxS43BBaUcGtk9OlZDEn4dNuRzwQeLevSKoz8KEkb3G
znowcWZed/p8X8oIUJkN2eN67BRBdTui7m8x2FCLVXbuTiiSj6P3l8IntkOFwf5JyAHdYaHxswzY
f8Q4LErHhaJ4aaup7J/K6jXZJ/Et4xFxdEZKvajJX12mDqVrGI5PKAPDN2ptN1q1m3gJV5ZHx9bO
DVBgPrY3FHCpTUV1qvmmyh5PLIpPi5Jvl2isKZvttwcujgkBdk91+q+0NVJuPdTcaJxVUZ4fx3bn
yRkTi3S6z1QQSmDo0tuSIJI22I9zAR1DvpqopvRlGo5TcuVsucH++nzbe3V/8Dpq+9Z+fSEN/UlW
1E688wMVNY8yJDrlNqYt8s/57r8ycw22DsxbxUwUIMrsVEMc/+CG2X7e2QyTSFJKRmmyGrVaMOCG
s8Dai+7sDdk2rumYzEgXN8jmBcIQrRZpZFKk1/iFMpcHRFaC503z/JM9kbzY5dM8BlFQ+YlOj/+Z
7YzNg3Ngfkk/Mhdt5k7gPemZtYIQ1QGHPDo3Z6Ih1tNfs6uOKJ9EqT61Fj0jDGuV9RQi4W/n2Di2
9KrQvUNWV6s+vPy4/Dx7Km+Vj2okelHOaf3OwFk2OCtwdxdeBxjjCa2DjMmmVgWlajqEav9/7jMK
VtEfc4JbnRDAxK0cYSFz0+T0++cnBUb6xSPlN0JSIHgzJ6OqIPwVLnqTOEfGJA4iiiVqckGUr25x
4llfIGX7jw/7tWdFW8zA2bOa72ActQHEd9XYDq4QLU0iy3PqouD/7PAD6cdukrGLwb9lgkZZGVHu
1IET23imcT8zz/JRlTvds/K+GMglK+y2nCihLhkp6grDb19HY1FnN3Z2/4sGRNF+46gHy1JqscJz
kJO9DZ/vu0he3ot5Hlo2FGjEHcqltotARRSH05+m1oNcDYTKnMpNahWeBRPs3KSawP+sV8xyTYag
dRH8zYgUh2wAhU8oC9Kl4KLiKQ8EkIf/PkIr9X7qgYEbCTqL7FfFTYfKNLljR34FR9H32ed68Gc1
JOVAdODqhlqxwmH4tCWFdBVKlS8X1lTi7AdvBCwSjDRDIhNly8zb5UqBz8tAJ8Dn5FmqA+26IR2A
9aKjRaVmfvoDibPrdjPwcJ6ZL3ek+l2kB1zT6If93UI7yWz7zxernHCK9jkAeCk8x4p0AEnf+oDe
1f9y4x3HDIJK0SXFl78IMfJHQxomnn4Du2dUf6sKHWsZXQlQLBDRp58m2jBZ/GrSij6ov1CN26su
t6iDMYTp+YrlPTN5PLq9Joli7qSWo+Zgo7cDslyMxbShLI5+XdzCTv676kjJvsPX6eTkDinMn33m
uqyNBr7z9KlldCTqobH3Naou/PrzC3bz4ovOJXsHEef27IC8yz3Wo+tf7nY0xFTuuL3wb3PcFKcH
f6gOhujgXhRcjL/riPGThis2hcVo/RMMMZjt2tdRCncCAl2aIfHflynF3/mcbv1Cf61F4bKnT6C8
YEmuTwP9Js4p/7QM9+LN2JCCHtxpi98dIHLWLRyDFmywfJEMi5WntyxEVL0UnuZJZROHQ6DNiX5B
5rKXV72MvVhlrD4lyMK0ROh2ZjrTW1Wkf1iPi2682qg4csv1/nb83Jl8kKcdYRVsRhj7IvuZHwwM
47/Y7H6bny0tmjSWjxSQgtbLAH+s+IKsc+ZWtFyGCtYZdU0eXAKHvq3Ty3IeWTReTltSjEzAJ6pw
4QjVXTcveRnNWkxWZ//4/BUcrf7fq1mtXWL3vIujJqxO0iDVQTy7IYp/2dSnMJxltikkuIKNmaaa
vqPnH3iLRAMkSPL8ST7N5XEBCujHXYLFM7WFgh/PjOMg/4sBLfrr99XlPQFA1FAFBDFeNyI5XleX
ZNBqkO7vTKNbZUdxkg5D46uJlpz2UqvbkvAOuXRHyUDaA/6yFM3OB/W2ZVrpt3/NqRGUKFHS3iWc
o9iSGhJCfnn51Vx9sMlaS7ssZ5UvaCN7konTOHvVld4Kb0XugdArM0QL5o43b166g1XDVcyy662k
MjbC/Zr3v5cETjnmdEP26IcFe4zwR/8nYb9jq4VkTdCahLHyWmpHn5Pxa3gHr/CfK46EicZCKKEs
IDMmb5x2WGrJsQcmWHTqhxgeXSG9piUTkciHBZ377+bi74cTerlLaRmaQRtgj+vqy9nGBzCVokHv
OdTr1yhJ0qa3l0q9icYFWpI1MUPIashnW8X29s3raDqJZAflsBbdfmvnnsI1pkCK7krbWMy91epI
BKWAO6p0SpJCGwHUTpTm+S3ZzasRucNheQfaaq9TXHHAyCvDtHz33zthaNP9WY1jRB99kmyRc82e
eVkqdfAnXBESx/CTk9SH1nOltwAt1uEXoHvU0cn1PaMSZ8L9EtJQfhRXHQFdTvO46QzLIjlLLIeq
tqjrAX7Y+BwJmZ1qnezNoak1csH7j+eRAb8xQXRdbfnCYWHyu1Wyz4/lUfqDOwYUDYFQMF1gZ+zC
tKDXYhew3Dqo66Pol3hStANgeEuIY9QQxBfve3iOwI8egRHDJHPY+kf/TvMDQpDM81xzHmEbH7Ym
wQhjCPCptoBwu4Q82+F8P+Z4Ez3L9dQGlB/btBqMaxMAakvPa+3kb9yzyrb2k0xZIPEafNW4B20W
B8s6HBy5wCLh8RhZULvSkxEsii/5+KVNd0VFaS4eDTJ0IkCAEcTQK9Q1vPXsq5VOuPyHF2A+NM6K
7AauKu0ijEgdr2E+q40iYkWEwgJv7QdDWyd+1g3GV/4wT/s/isfWAuHjjrKuwfuYgyGVCJEPlKzH
ZtgZ34/0uFpxMSeH9+nBh+7grROARNCvM4BloacQiJii32gr3ELNqWtYMTjDbp1L/TWavbh+JDI8
xWs7uTsMpcveSU2GW9cXxPK4fQ+Il12ph00X9olHivUK1b5NyEBx9On5xBA3iTHuuEgl6GFL6FGW
yEJC3xAh5/1myXRsoZT2OOMWVigJS0sDFQchMXXbwizzXUDA9StIoRQJThbEuUZ5hGV4gTOFmmA4
daNOWfVRwcEX/yLw7Scz/RGgKLUPkSvRyyPFo1W5OKNli6u1ZhNGqOuFvGWOE1vW5lZaL/0gpAQo
HBHNbzk4E03QIa5L9GdLCwZh8uRkuJ44NS/at9GF7DfP6ZRVpn1/BqoL4vUcEAxOT84JgQy6MB9j
WDB5KawibQNjLb5HKeky3kXzommfu0sOJGFklqJjJdTY3xRuv5NLYNosgZ5dzQ49o+3GvySUUK4T
dd9rlPHEE03Q1jVqvT91P3ne1roGcOmzewhmwhW9VRnntRoficBkKr6lL+NRyZLxsY+FfOEXkhem
06I+EOzr6rkZ2w8p1GWam4FG4jfLNnQDxxTwpyU1ishZtXCMD1zCBf6ZUTRCyJ5tNznffPXhtPhY
HTgNMdCDpVCsmqXJpdulOII51IVU61ubIg3d1/d6cJz1mFkHY0oArZ3dvsXGrPAmq9g1CaHATXjp
x9xlXwiDkEIlitKfd+8yezDLDkKvt8iGijVQS8KCATwR98XYi1cM+8kBQRplPg5LLTl7fsDpB8iN
+mGN3vk/wsFfeuCcoWZMmb/HThhv6nvtOWACNwF7m8xBH/b6poSKx3wjeJFyolVp+9v2bFZtA9dD
6ETeWW1MkGq5c0B1Yvw5gbtQxZahTFqP+/F4cp2vYdlYSA2+IsO9tk1KqqNVEqQ2EPDj6EFIHHE+
ZAXVAsES+ZBR0diM3yLZBImf3XMhY/Msqr9T0KeSUs19kW9QqBOwlPptFNjC1168l35t6AgqHDOs
ci1XSKIv6RnUN31klHNu6aa99JEuYsdD5OIaNsmGV/Xz2nzSy4uMMMJAfrc6xThjRu8Z8uFB6Duu
Ywr+Tu4SUAsiY8UjmHMcxjeRewn/quCwnyqJsMXK/nIqt2P1v/qfCyUc6E0WkWB/dH/P8bHF7qpV
AmFArJC1p2y9Z/u45VajIbBPYvgYYSd7OaB/cYb1JJr4hjdW3gohpigvHtQCbY93eLC/+KgYmRjx
funArQrFYhacewxxaeYQhHG8qc1QOFfCt/2OibADlysGeQARZxwdcugIcrpKLR1BFlqi8TyC/b/p
jruoS3Zyj7rJuUZYNHadGjW+WKc3B/ATZJPFjsOEKIHO/K4Q1hADY3VXPfLJDzFxSnwtDdOeW/uL
+025Rq5ocelYXqYDnrDC6XTuD5hI+SMkc0cy2PUHXP/BxO/PaG57jkQO7iT91JyiR9kKZDEjnohd
bV7tQOU015Q1oOwMJnjbFELEAO0xSomN9vrbDTDCmCuNv08eK1aeqyRYYdMN58m98y0pj568MBVh
RXjeKzWeTZC0cRVoRoQuu1OurdsXQpi2oZ3+yGM8tXyIfRJFiwVHGA57QkfUv97rwBzzVMvxf/Qi
kVhGpRxc5VzsyW4uwqV2oMLoy78oo+OyDu06r2j1izFqNytYY49yZqx/D0UGevZidosAGfTetMeJ
VjSCCYC2iGw8nwhp2yHF9QwclSxQM5foVeKVW5xXxHVSOoTcbOVLM4hVubTGBtO4VXbPI8EY8OIL
LfSyf4g6ViaQWKvFIMN3Imwx/SDHgpy8ohbQ1f+f6oTAKFP3cqW9Jbv9pAyw15Q4T+z/2reklb1R
T3Mm8uxssVNyRNkgdrRNcZvSWmPbi2WqmG5IULoWLx9Lm5i+tV+lb3K67LtBM4j/cJjyAGJidQ85
VsZgJG5Nj/C3MzoraE5IdkjXTNPfoH0zqB+OJA+eHFy3Xm9OZiaXn/rwK4l8NvsVeha5PvmjhBE/
mFmXi+XlH1V95p3GdwSsKPttRroINhUe/oRGX34XX6P174Ovc9YZG8feeFV5FCg4Dvbwnl8p7yA1
Xi7ScZPeWbp8Ix5wHY6lsP/oO9XMvBjSQGds0lKi2iD8iGFQqiHlRIkyPW25sHtsoIrfzv0/FKRa
sGkGKIGiKPgh7cTDdTQeI3SOUbd9H+UPHvHQBQFrwaRMqEB8xBLmrTkptKoYW+zkLfAk6GYWcSTz
Q1qRnSlFY2SMvGCkVTBbTCiJ/36wGnQ5ubwF9YCsyLJDvskdVLvUeTg7LG7qFAbGQlUnBJBYdtec
vBrMjeWX+64RxtY0WRLlzbrNFLEP2JMXj42HUOQjq2UIzcDAP17wCTgB/tJa6NMenOqB1iWjptIk
IxKntgg6zg66eQ311JtS5kVaEEDHHz41LCJAZjsJEHndcLLFLOdz8v65+ZmSlXeRWmSHQOgsVirZ
Uhv2fSFMXzUxTI9lXeJuKq1zrky/Ksm2BZFRW4ACoduFXqexA3OMtfBHvwkvDOujsneH2WTr5n6p
T/akSy6VwvAbdXIbtSWiHPT64CgdxjxWG+BepJ7yqoFKbEypOk/91q8LHRNREBcVbckoDGsTcjk+
1jEfrnoaedmnz8sBI8Q5NFLBFy9kgx5udK9yUShGD8VecOeLxuPPrAG0KppB4ZJIx9OSMNu2bpiZ
hkgt1lz0ArH7MTG/tZxn1ROJpp9BFi8WYDbbnNn8U9vwbim+NexdXTaFwAOQj8rurGQDYL3Vm8H3
zCX7+OJ1sJkbPc+wAlEATU4ArVhkKgZzEbRiEvTJRIjbrSCkgKNTDjWn4wm8XfRcfNC9TLHVAvm3
j0LAM7Ij4PiwmV4SS4+6wKjERTL/Lpg+NkK9PUlQumBqLpLVlycG+vb652Ob6Su0cCaDTev3MQri
C4rgDIhhSJ6y6u4mmmeBdwBYDRlSo32y2ALifiA1tcAAtx/c9kl9YlC1bExyfJFoTdbDY+Tbh4pE
uNIxnOwpdpVA0r6ifjExD3LJ3RJx5+HPmURYXt249clwBnpaEQU7FgjAxjAZlvwl7bogY0+D6U+6
K+Qc+lANcr14UNUqSOMA8OewcAOPAxxzLQsfx3/u2RGa8f35fC/MaiXmF3F9r8h+Bz09jzdAjtZo
vs8ylET5/0M6zW3eGoiASoK7C+7c+VoHOTqS0lEysz5dUkCfZBdcYPk0hly1RMVS2twZh/WFGiib
tRweD1u3QSh6i+t7VmXcFG0xWl1BRJOhRUApWX4oqAb61wm6SWPLnDfSkAEPCWjjvHa+j+k55BSB
t0DDFdnGVe17tXqKKI26FI4OkktmwGdo+2oaX+qcIUlVNQtJG6XzUh9DD/rz6oMRlIiWBXtbAuUT
dd/X7OGVtCFxhaM9SZGkqHrE8YOvjHNjgob2IBTvHEmD1Gu/+oMzASjErf/9wQHsVFQFe7Xfx8bc
Z58eGN66LsOeLJL5wX7i9ipNpGj9SrXPCl/TTjvQhteVr0rxHokCsHfWPgrkv3Qu0iKpanYlBcdi
wk0v+UtFI8HMXoI2yalNlNtkK+YDBr6ER6J8pnhhZWNIHvKTVkFqepahr+z0aY+0ItGIuCnisvBE
VobbUU+jqqkejdxZbVU42qwYbvXrs2F8hoATnuxOAUQuWZeRz6+PKyoXnO5h+UQ6q2EarkWoaLU2
TSi1hhoMtrqsFz6wGHzKhhgCpmkS/6WwdR33iX/t1mGwQa0u/Ygi3COw0GYXZL14ChkMxA3TAuR5
jyidLw+ZmWA5SVjCYkAkZhTuyz3C1SSLMF3mLuB+yE7z72K8vzDxVxGoIyw+Wae7wNSzqQzSQubU
CeAAKhdzxsVzap8NCzBwHf0v9EcbTlrhzm0UYrYfWofduuFHLzK6Wx6gelzsSAUFX5zE6xIkCLZ8
zwh4vyII1Qsr68WNBQeLYwLBknxXcxuzyfxXlydFsmSMNWe9xff+CANJuVIrONNgNV73WqiRLJby
SKPSAKwuyNfuObE+RzAozmEbguwaFpajv/h+fMtj2lfx3Ku3xYs4k2qme5ljB2MMCOkf2gUafRWa
EgDUkQnDb02X200DKU/JBPgu5XIUf0ikD40M7rwtVSMmPFAR4nVBsBPMrF+fs+wJvLvwklWSn1lp
1u82I0mmsFOrKeijEMydxPb8XFV4vkGlXf04Z/xeBOphc0PzT2PNcOtr4YxvNPe2kZd6SiCt3pdH
r0+Sef//TJJpVJXRly0pM1SqBM11qeIW7eIYGaZfd8/Kg0fdpt4zvxR1xwlGEIx/zCPWsQ/1FRO8
h9wZfntMY8xF/245cMp65qCsIWwbcQj8nJqBxq2VZwqnlapJYeKxuSeEOAetchqhhvpTQypR8bck
78/5VvQ3ZmUUveDtjqMuim+6BoA4SjCFQQblUnnYmm3Ct2Q1gclTwesTtcQ5VOpCF2lZI6bTydGS
Bf0NWCrQcDzPMAXSst8Q6JVj8ZVwiroI8tUx/0EteWYa2JkyyrswZeVXzLcvV8m3hP5EBYiTHjMh
gnY31soJCsxhBc4fBLJp3l78TAK3F+OPORnPMqm/VgOiEyC3mnjoHvJnkJXK3UwySe6JSTc25Qih
AfF/hc8+no5ovCAsuXAeGayEIjr8GU+HjW8sdRBBXkDCyRiruzu9N40F4s2UaTE8t3rcScri1oDo
8HkxQL7Jmu7CT2iN0s+nSIrA0ad8f3EpD7KSQj+aYfJAnRXvHmhOKbb+h0JW3LcVRRCV+Uz+9oPY
Dl1XWyuuRCuq2Qslb9NGIndF5iG4eXELetDIEWbxMvOye5AH8FEz14O2mZ35mFPfRTIvfFNjNUbo
WMoW3wFagvGhkbH/bisP8dA+0rxBtNOQokdEYXOzoriVt09iC6g6Td1K2j6JEH5GR9wvmaPhe2zP
LFitJT1AOJU+Nnv/iDw1TiVAI4V4G4yEYUuDzQ+K06sTKV16cSscxhryByO3b3xxBLInSYZRAbey
u8pPGBj2HHDHynx01/0n/nGkTKZ0JjSUFp3dIMkmchH8jWnWTItYDblds8b7Zxu58KXFvvdHgnH0
S4GMGErD8ls6K0rhxfNN3/dReajE4jUJEUy6yOIhFBMQ7kHZx1l9wRFHsjJ8r3HeZsfsV0wbPjz5
U+f+rWKMA1IzuAT5A23zURPjHk1U+XPxLBO+hyMMprk5A1pxAhs6s+0sWLP8E4Rzs+D3SxgWr2Zj
3kJKBp3vkC4S0GQCPjfuWTsyCxC6dgMqDP7WZq/Rck+Rpbb+AcBl8EBJEx/b4eWCzuSwJ42t3Lgo
MS5ACZWN8PMy0bYI/JetJoBG2DU0uIe6B0avg4dyxUUzpeX583l/0kJ9sp+TXa6n4zGgSc3bEx9r
H61Zl6JN62h7HGVcRyGoQtx6IRccGZ411f0KyG6/z/8IUEfyF8c/ydaX+r27/0si7BRPH1f1ndqL
B3sW8tEa79sMVC9a0eP7Sl4gt7yo0PLlYoz9yJJzpBns0rK7u/vix7zgQtdrYc1fYMV7rgXWZjW8
65PZgKqQOAmkQZvscLPw/J7hpYAW+RkuoQ9fJHSE8HFsTxZxNi+Oe5Xb3x6TO8HrQF6MuMRXWgIX
jCW6VnfEn2+jORA2Ccmx0JMwLkVhjyLN5jLG4PqtqM2UTf4BHwH0uNFSLnOeUsYcR5YdKFqJu1Ry
CsgEvYd9ukvQ8EEeqvg99zYe883xHd32k75Kb8x0Kt8xJzgdSt1wQKKqTecbwm/oys3egrlQpAl9
S/Uwf6o7IkraAtHBju27It46GXapf76e7kP+9SwVeu4aqwLpiga0NRxE1ZAvl2gEsaeIE3BdaMxd
gXC0I2LquESeY6sxi9+iLoRjd5lMsN58kvcWjRPQTtJigfFcVRE4mKqJkT4Penb4AZeYxGVaRsUQ
NBEBWa9XBLtoPGRopAALrMQL+NE4Xt2BhGVrdECEMLA40D+8EA3ohtcSHjVAe9ZcivRgiXftkAhi
pCJPOEI/QoKoHujZAGIEfm/Si+ic5MJlGKUbGnHVmPGb8hnRIllejQv61GjcEThZfgExqSqO83wF
1u7BU/3lvjro3dragG5s12mDdRgbmJKjl9YgsgUvBkMZEljo/PDiQALGPH4r9hp9AqefkEgzwxrW
yJpJyXXUciLiiUH8exPs8srAU32fyZTZCl9qrStIeAO2Wx5jyN7jmFWWBIsO8tltWDqxOJ3oRT9Q
dn91ghuOc2Rvi2oTglEh6Wl3a5zmdphbMgAlN2b2wRpsZU9O/rfR4Pwc2jaD3tgMiGL5NM31F0eu
VuFykKAgoIK4xXAUW8QXbpZsgyh1zDmS/DtOq1kInevWv6udfxiXNFQSpN+rVZC6YM3h06p0l4vR
qeF4ayRZMgCww3ZATrB6c02LknJH372FiktPu9HASBsCY659iXbe+BsLj9CdTQbs3dDiQyf/w0n5
KrU27gAMcbb+F0uT/V+ZOS0KUNcdcBLMDxg/ZD0wTfvw46aFM45+zp1rrK5N/hAMBQRExDgUvMSj
MacXtz1a3ZO6Bf/d36SbOkSiBvQZrSD61xerRuH/Q8cdqY0lwNqJj9ErST1RvWh2Q0QlLtu78n0D
gtXaUAr2/rh1zPcOb5CJCTsef8dVeZbiM99wh3XKrnck4EGH6Uc3fRTFmPH1ADkm2VfV9yHEELpP
Z71tEPJ2ihwqCCXQywyvIruUZdGNzx62ZmRoDpjRhgBsMwihJKnIXFdzEALXmLm+FW+Oi7a0JyXs
gOszpDic7od0CsO4mrIb8UBcmdzI9kzedPrNoUEaZy+Uvcfuj6z40Qg2pETn/EN+kP7L5HISx/2V
0Dkbq2pWV5uvHtR6WV35Vxiu/2VAlF1WY9JH/157UNSGDkZQsN5QWcRqN41cD8Ueh+gtCxm93cwI
HP/lYTYZEvjp+INjBHstgNK9/tuBYZJs2lnjUIBnOpj77frYyPxlTTcNvSYbeFjY7dabvuSR7QaX
bF4o+G+WEiyOmZBfXVpNbk2ydhuoPBC4DaLPsPWMkxTjxZ23uJJbifKHFJpiA5eyWvCQJhJxKH8d
tUDLhkBps9e8mZuaqo5fhjsZTM3GE+xMMg2ZsOhUYH8Vw/zgm4TDwT0iIQfv4suhTp/2IsXOmZae
L3Bhi2lYH2tivhUXg/rj81nsB9curPDJoA3nUxwqkkTN0SiqnXjxJ4DzciBEftAOxxDG4UwRqSRv
uTkHvGiMhWfsstCc5OUrHRig6IJqAop14N9x4pIiQl2RonJlGvMkevGVNn4wrMr3slrCQMkqRDJa
DFVxErLNzQZ92ZvKfaUjdhZK5rTgwpuL6OYU5cfF1loi3/+05CtOCzAWkWUwvM9BL1Yim1QiNt8P
pxFD+cMukQ7giw/9xLy3uiSCnNLoTvOmtDMOkkHrH8rJtreEqRHVjLLp39Yx3vwpHTexT5X1mgIc
uFo+Phs9FHeBqqPH8KPH6PXiRpbdt9L1SF0lJH/nlaRMaGG3xxTGe/gYCq20/jQ9pQC54EpHEnc+
TxpQft6YDAOpB4+mLMoIn9O8+pFiaOU92f1vVKmtkA0VF07/fRBqM2PJVaME6apwl3pgFdsspppz
JPIQoSX/wUkcPHQP1S68q7/C3XxcepUgfCiFYitG4W1UJa+cB4gEGp9gPi7r3AEnpxAcstsOR3Aa
YFG+adMh+9kzmQAdsiFifXhPwdDqrGlpitKTKohWvP1tMwgDD1LwI0RFqfNfySIWm7BcLKMP8DNH
LoxhecdFVrroYjFr0ssQ/PeFrOwOLFDOJ1wS2AKl522xTTsHels1aGAFAt0L2ifCIdtLuZ5SFZB1
/+ut165A0hcW91LubAQWQZ1lnYWtYFkLhT0cYfLPejUaISdH96mOXa4bP546dYr//fUMt09i6laK
nKMGulJVb9McVJBMx+KJ0NMdpouSBd1+6ZGU3qqJwk/cDgJGhgCoVjg6Y4it4aQS2Mi3USkZei9R
YcIwejBvcdVAavwcHFnTcYWlpuuWzJacR07u7p6Aos79FSRZfW83Hvn+pU6KUNXHQbU1Dxeg00Fp
6eUC9Nypnh0gHzCdMkEryVn0OGvLx4UBJ3jwkQribhPhiD1rlj/JwjStC9mJzJe1kkwxbh7NgwdA
eQt0ykaKTjke2zx2jlrxZhHqYby0c69ut29TzwrNhh45432q3sw5vPcD9pLYCY5pPHd/k026HuP7
dDu8/ws7su0adgaIpa6Ejbzj9a8lzomWYIlMADflCrzkxxraejMDPbYVw8ZQfatETd6o8zR6S0VY
ibaoMXMMmUOWn4H/bHSOMzy/cE/k6ME+gPF+cZDijLGiHl8632ISEKTOe/eiV9hVIkIjNSw6SgZr
94xQFvNmRv+9Fr5n9E82hrcwTRYfF7BCr8c6xHI0HCvrGmh1MGEV/k1DMTufW20K1R9RMjWaj3qU
GF4T3j7vc8Merh/UXP0wdAMeS7jxWAznfiRZtPLLl7z5XzkYX+YQ110Yaz1K3QDV/GfwwJUby6ob
Plyv5rg6B4D6BLEleEmTEZIeh4nRI7k+WW/aNFL2Nov1Al1EN3QdUZdC+t4rB1huAvmQOVdl9oob
4f+hqfbuuBr0ll6r2+eGNvHovR58zD6wBJCoalsMTwkC1qAk9JQM6xZNaEPwOduM7nNxgdonZkXA
QTteiZ4TyAGy5Njzqd9g6naAjeMaithVQt3adptGNBWUb0ujwl7AoYkdzB0mK3uA0dyzBLjEPrqK
lhiM9tyg6MC7mx+ihF0U1l1yd+u9uNHH056QmlHGVn6AH2jtZltqQRGe1gNZtAisrACvctVwplsS
XxvqKJnf1IQfkz2pDmHeHq3LIm8ElWhmFtjhqOH3BLxR79zE2rk9wAIsgjJ68FT+o8hFxo8DDmof
jJwBgIku/5ZNkz5p7/pzgaO62F2Xig0F41VnohpgXGc6ctuJePaQ5ZyUCm/RXyBC/lLnjJonZb6M
9/yuzhB+SJv1OZY4IguwKDzDTD30JKn6KqtrOwZLCNU9rEK/mHrQfaOXzZJyPlwzF3Bo0BP1wZ5s
aGHE6PAqlyDwWAyv8mxQtc139xMklqk+hyAC1YXQy2pGo+CdMjtKrrsWrz4ImmvtiHQLFa0BzFGo
JbBPGN+3JQ8awRYvbuPygpeXtCb3ml6Nvq7IEbxNlNke1yEZRgQsmSkZMeZw/9zCiIT/UFt2nvVp
dDFu2HSWRLXXPglN+bLaD1YASpvoiMr0JdYV0krFomJnY87bBb7kUVASt42Yz2EAd1Uy0NmypMNX
92X4XD2DefeKBhdAkC9yLmUDoL3gdhKJ71KmD6xQ9HBb2UDOSBDefnFMv5pDPtgf+bncDlKNIKzd
+M4lumC2R5oEtVP4kSqdByZi2+bChIzsXDq6jRjaHzeONL3NzTRQ/ZCyqdGSYVWvc1xP3BWUw+Rz
HTirJm2/UbHsrH4HSZMUyHBkuxMUQpBhu4lr2bdrVBg2hgANL1/mCDDHEhfkIV1k+CT22XbkyEZ3
zglMn00VcqqKqZKW4m4vjyT3z0NLGRTEeElz8npLulsZG3xj1jb/J5D7T+aA8HxmtMD4bD8ykX9x
8IxG9umWngRFr/oMCOvUhuvDv+dP00MyRnCsrVTrFyn9DAuI65Z6viLpyyJ6U4RDj2Ken+0K5Ae2
tx140vB8cF8c193tPHOjXlQdkkToAGG2H0E0evVDfJxcpZHvAY/s8m9BSZVI4vYNAUOFID8xRudg
k8GSXoCfk66rq5csy0BRntnc3L1JnaGmdZGn7h819+29h7tN2BQn+91Acrifadh4J0r5Rfuig6O+
vkG/vzy34DzFPH+RtAkYMAeZYlJYgECTZ/UazSRCjUzN+st3Um/zw3YYj/ZbVWBG+oc3iEcs+0Rw
9q2f5EoVkGiG6piDWR47eOxljr6KpG/XefI94ixzv6/zqR2zllrNMt5I9IwOTVETrLotjcOCHaUw
S+jAwUPZZjnxlvSX0PKk3/syYldolVOTc8TSO5f2K7EpzQa2c9hHIeCPiRTbO9azxznJJiEGQZte
B4+aqWbpsZfz4af/5+CvqjMZKNIVB6vVfDB2ldZ7fQNSVKAjfS6fjEKg+0CbuhurKWD+yUjCcEAa
235C2f6T7LZ3coroXxKdzsFt9dNPxXWcrDwdGqXEaI6di8QwV6n2YJU5Qf11hGGiCV4vdC6zKivx
FmYCJ1/6UbpotSrxd7rbrOuFvj/JHRf5OnVXOIIcVKAaLYsVtDw6FQ32Buw5ni0h/Ic8xgS9dZY0
y3hptVnpw4Ujt/2KxTeoOq3FzL4E8OQPeJSRKR/ptFJk+tkpHwt+sSTAvbzh1s62RZKRSHbqAE9p
K+TxNnXQnGPlejZBNzOoQdt10HWGhS0tzhT5gtj+xuc3063t474xpD11Cy0pRWEUJgXfx8vhN7QR
4Xqnd4dJG5bft27bJY/pBhuDmRxMmXcXrE5Fjjzlbp9uFi1EAqseauuz+sjVBeVN8aAn1nngFYyB
0pYxOD1MMXKwBSrtQkRytwYKeHJ+09TMaWwS3z3p1s8QDdbdxT1FEAvv17eePB8mzlYHDBvpzTzv
fEadPm7ADZCAov2wyIPa3m6hKnv7r6aREhc8mWDsjy74erffC1a6oew0k8p6gaNwhG60DnfyA76P
xRtQbYP0wJvoMUd/gY/RzaEeHyNScDM6/QiZ5QM4mzkoqGXsLqYCt2xDlDeXl9ioZKcqLGATs5PY
IzFphSYmsCrldh6ph2zQwFVato2QAQaZxuh19Kh4xzzhkEAlYxcaHmM5aFMBSubl7TaASrz1H5lw
vqrwE/b48vEmsJj+GqLwkOgLimp3yOhFliV3NjO23t23dkggPmg/+DgRT2gPNuCX/4w+rjOfS1HN
j+0Ma7gzf0pt2pmB3QB9hCzP0Y859J7C0awF9g5R19RfNl0p7KhQteUDt/x4OswMP6KjZFSDa6mI
NsF1x7F+Oh8x/a5fACyHHwOd+4PUCieFx6WwnD37zKPji7J/ZahaDRCuAYVsHaWd2p+ZvcWQ+1Do
EXg0fOxTVuYKFmnr/21Wu4PmyeS4bcXzVADS2rW+DfAuUOA+LjpGIfKyudTs4sePow98YtZn4W7V
n1YsTtHWgCcIshni+DvfNxwGJrpcsT9IBpEIzMazbqbmQXyX8u6VqJALGjHO3cDGIuw7JB3Gk6t3
RzbVSYuypQFVJsvUtiMjcThy/sXTD1NUSlgbRgh9AQKUgw8tmtRAuHqIG90EMcmdIRCLLDfmm8uB
EXkg5GA97DKcI2egQ2tsznjNd3FIX6T0XcVxJCpdy96vavsuuzZYNof75asUGzYGkwiIpCTiRAWP
r2GmUrHuBc7EMqrJ3PRySmPTqD6NWXzw872og0JJ/4vZyyVhu4o073JC+ASD9C9d4mNoIHJ/Ahu6
s8gk9b8LKn/2NEihol/xoFx5qkpPGVvlqwtATLHg6kIDcn12EKTJCmr78df+STlw+IdtOW2CG4WH
9oCuJNKA6yVFUj9o7b9y5sSbHdZpIgE1xo4QYvGhI0NQSBm9d4n/Eu8yJ1rXMX430J84KPzRpSTr
ee383A32L7BMvuOGKoumt4QuDrzSM93d6Q0jb6LU7/SMo25mx6lW8HMpADw0qwi3sPfZ1VdR17R3
oD9SelrYLmEk58LASPZ6nRjjtWv4BQ4+/XylpaY/lfRv0IYeDQYt6Z9hzvwRk1REbgLWs76MTTzj
Dd4vlUwq9o4gS5YXw/dlFxpuwWUKUtjub5ay9GaMQDERZBuMngn5mvnS3ZJdyJ28D72EDle2TAlD
zDXvyAWQxx0JczG5Dj3UIYW7dMhr4a+LtkGxVAPh2tD4QzUKoeUvv8vnJT7G+iEZCiVrx3gSVCL8
RkEgWvCjNV4/vfeUlHKt60+hdzUeVnfKVAudJxdcDtEmOyBu9F2QFHqkOGcXD4m6Ggwzo9KWuGHg
Hxujid7+e3oPLT/sWsJu5xXo/KxzXW2khFFjFdvEmKgL1I82W6ZU36720xaRIAe1vFOvqj3bBeYN
WrUeVIkkErQo7yT/rxEJ582aZrOZwWgomXa8ITonLUVStXzyZMDiRUB7cTgAUisVLPT7Dx7cqFoa
1RA/gCCOos56lhcn7dmrv7F8tq1xK8SZPR0KzBmLXzZ0AkugPwz2GYtGsByZCE8QY2X1mxkH6QDw
2thoz0g7BWMxUvpsdTpePEtA/Swo/KPA6N7+ieJ0xNKqONefiRpviME1jAUDEywUShGfMDLwDlUn
3gD6vKNNo41AN/jrHAhWprClI1Ha8zGhVRpentDzVHKeDWM9UxBqrl0M3dNAVPs1/2a02lyUtGxc
qNV5xZXhXVP0dDMTCn2gFZZ0C4zufFeVN09ICIjtfk6AVcCO16FhuBGoFSeUeSSoOlhDbexUMmBU
EIyFVGH/jXQgYto2Bc5cDPrYD6xKGTknJwzyL7cHhI7VHG4oOHy96OUyj98ZXOxwRxfQ9C8ELD8W
v+k8uIkXn74CrFQ3ymJZ7JNMfGtfIOHTNKKMMMOQywzra07ysSMP/FatLhQTZ7FKXu1/aBpnEqlS
0EqShQWkcTrUzI8ldjHys0Ecn+1nQxPr2W4XYH//d+dhQqUF2yNSRatcPWbG8neiwfEi26HlMAY3
Vci6+gKAp48R5X/Sey5JTxPtbEywbdHsYKujRtNonUBlR74k95EQClEr7S2Teg6OWOqnyHsSO7Y5
ZMNsj2x9DKfkip54bEVFm6EuHk6IIwmiXQvTGDMTjZkHrMr4084raCb/Q5kmwnbOezh+ADFpSdmP
nTIoxyzb84sdx3gTsFfnOC+kZSGcKz0yQFreG1MELej4c15sHrP6A06Tkf8kIs9rAcNDXGwhjRx3
nlTZAman6mdr9JXL5xWWvscbyCIKwYnrTyU+mveRI+Hvu8k95l3JyQvrpqHUiYpOoGnShjpOMXxT
zYiN0ffPi+JgCaC6qXCDtDow/8TxOSZqbAJ5jCv4Wfy8XuxGfWmD9CpG4uCBjxn1XK9YrnzIU9xE
/feQRY3OI5zc2SpH1Ki5L8WvUUZcvWrn1CuqN5RS3qIqlhsvlxl+PNfLvgizge6oi2Ga99nx5O2y
4o8LzJoeliTsDtez6FgN6tcKi6m9oTyDaLvws7D97NwWgKGeVMy6Rf5G6D+XDNKkwwzNUElRPhOA
/Zid393aLZQ7wQnM17px9rQW0uQyT/OTEcF5UUg7zhh03D06BiYu7MIMx3q/RcJc8X8EfBwvnb1T
WlfsyOHEeXlDh88X7YvYaFEmbFY7jlSh1FRcB6Y9K2IPLbCLy75Kg2rI4m5d+pjT2UZMXQIUYsy7
qEEAUabBmD/E/hpYmq4ybNIN4m7DNfMLoAv24hDJAVBKgeZ+Ai9W/EBaIIh2hMdzdFkVLi54LYgg
OG36gzBpKy+FLIJ+0G241AfSxypKtSEk7yKH6TIiVNp3QmJ38fQxh0MHNiOzMXC6OX87gKUDYynA
Xd0XzhARphV9vve5NoLF/Mp4fLpbiOciLKm/a9+z487/eeHHKcESX1Ku7KJ1egSF5NBbmSJHAEKK
FMsZ8Fp0oIOWk0XmD/+TK09PJR1CfJoK7rZpDG2Y0XP4mDHtTPPKBnOf/i9fpdL7Ybq8oel/eP34
UL0A2gxNp2XnkI0Qyf/lHmKXxyJKkna6uIpacs5g/B+Sqi9lNKabTZrjjJlCYHVnnKqBbtxIjDVo
lkFwl6/6ewp6Z4cmr7CDs/WGlS7QvvWd85vUhO3bJBcC7OOKJwi8OqYIsZifeCRpypolDHA+9ESp
Rzpe9Nm1JyxGnIZdWdUHqhucqEviOJuVMl0ZQr8mRlQSGtj2n+B0INe4jn3zfSIcCiThlf97L2HG
9QF1FA8V5lpHFBVvzlN4S1bxd20FdHSrUH3rKH2FycmjKbGa72Y7j1jO8hRA0fXNJp0Zgh/XAPSj
CB8HWV6cB0nMZ99uenSQGVJXmNQiIV8sAaG2mU8Ni3hGdJ4DaNuWf+FFCJnjp2v+b62kvPJ2qeHd
plmlu2zzWDF6zUoMdpr2xc4OHyWukoBrXOtwIl3liSEpWwc4GeWeHGw0Pyxjjq4RFH3OeHC1a4U3
MiV5Z91ikNGrUCDd+5suXwCKTLIqNNNimNMMOnNiA2Fks2rjYYLZMhFIR5zg+iIDsGr8ByuZO67b
DqmqRdFe20SbZf6NdfFokvCWGC42TsO6LCvczQJw9PL2ylRL+OcweyfnUK1JUu5dtykute+P0FBx
at1pkRIJLxHgtJvSSoWEcXtOfMpI8x1YS+1n40kiOouxZZMQcU1HpQdsWN19dyiwbndisPnmfakP
rbsVuHKf7cCjNz9rF7Kf+Iv1PK9jndyQTLiPnBPds1Rn5OXoY/nvSbsz7Y9G5CdBOkP78BzsmleQ
nvzQgEzQ8DbgQzuS6RadkWMKA2HftRoWZb0U/NmnyrqsKSHSOPX+WHpl6z8FyRXcLTEc+XxDvmCo
kq8dOmSfbqYUDPtLXECLNHxPs9ZMzbdajVDiEPqOR8bku8V7n+7O/89Y2sYRnNz9KaYOLmf9rXW0
xcfanEm8ReeOYlWkqCGMhxIPN175+vQBiJXhP2nLoXr5AFZdc+tYFO7dsftH2NwcNqEGDfqhpsUy
0QKKhEKbeUpwEMDeZssJ1CQXv4Zs6OgxDYSlRW+VcJlJiB7QVcZP2rc3GfOvsqhBYm5LYsJIIN6l
Hg2qjtcTLhBPPhLDAG1PxskXGLuOW2MjxbAXcJO64XpfoJTbJxSibU/9i109Cn8xz1cifKyZ0mOM
xtrRYxMyUUI22pK+n61XnSUpfTvDgG229qTxShdp104BMfXZBYuCckwhHjNrllRKOUJVPMnsQpz5
upR8bCiChjMl+jqBIr4LYJj8O9aB01et4VKzCl+rudi1M4qBLbqQQaDaskNQkbsMw4VYbRP27g5V
sdhjzP826nUuTRzzwpYfXcDw2NuEAvHy6GroRam6BudiB4h3bcpWyO7f4xwLlAcxuSO6JkQIdpdF
CEqhAnxrt3Oy2w0/3JVpMy856cy/t/Z1XWOuqsj7FrfQcjKgYWb+kwxCvWm0uTN6eCb2O7BcLXYM
rOOld4uvnoOxcW4N2N+naPVscURWEKhUneAB6hUKzaU3SJ2jPD0eZXs8kkJpuQwnyg2NHVFYmP2p
oKNb5E1doozn616yYVSuainWErEGs9GwIOmzM+LULZGaS2JHMUrc5GIdwkMGt+AOo/Df78cbfsis
ZFjCw7W0nZsyED9YHaU+KocGsPbHCL7xidGDGcRP5P1xthlM1jkyj+Kaoanq2+8JukAZKE9X+p1h
YwrEhhJosIfALWSrzF5kxU4Pgrc/thyYwpMq2jW4daqapTWGHf1BRH/zMkiZLNsO2++ivitLQ2/M
BU6wGWZTUCn4HZ0p3ngIvNyFvkbyE+mKFHNOZkuxJOjm42QIPmRpvm/ekNDoMgqRIPzUYYGpApzq
/NTStzFBAtUu0tq3GtsMKqvjdQ7aAkRodDAjkmIevqUK1waYYMo54lzPITijLUdAsgSowACN0VRT
sfswFcAAXkjFGf1BjQGH6qR9+kSOnpmMBhMFKcbzYbNSfwDRB7ukBJql3U8leQMalrO0pZS/N76q
k8eAGNxkZP38hq/bDeXe7G9dwkXRY5/HuieU3M6LXagTzo1YzwfpDRtcgp1iTk5iA6WxOcdlnN8s
O+MjmzWDkdMPFu7GAA/ugkOVogg71WMcA+5vmp/vlyArbe89Fp173lNBJk+DIvZN/rLZxrfNdlU1
n428yi87XnQCX81Z8jtdETWbWkeTCbW7aqo61nMNKMe3TltydjFGu8MFfOC0IF+4VCLM0N+YN5Ir
BFpom3b8b13P31OGYSoZnTYlIu4NwpKN6UqrKla/0r7c9FSQy5yVs6DZBTjSbtvDckdkwlGEgcj3
ugqXkmw6XZdlszGQtD8ezIAwzComATd4Mm/81r3Oy8cB1JlEQxszPfoWMw3xuLkxTXnlPedmL5g8
7nzi30bN4c6QNiBgeLtHTqRDAHkZZKya/PsdpyJcl4+ygqC7shnxQPWmeC4vcVgQRxdNwnoja6XP
3+6+UOZVPW+J/12cc7iBmSzMvmXfMaFHu6HyCihT9foEp2K2oC2vGowUyWWm+pdj1LHji6yzPrQH
nn8a69kJfm9n1eOTnp9nZfzMy4YsgQEEA0vLTfcyHuQXNz4o71izejdmSwfNwuHJ2XFMF0FB2Qjc
Eo4nXyXGBF9vUCbTG+2B+z4eaR5UWrSyPGe5TlwCsaH1p5wficuPHsf7+w3Zm8GHFlBeYrF/dBtk
Wlh4n5e2NWBFCuT3w/QQw2q3LyEfsdXmXWLdP7MI35FdCQvvx3sjJhb33O5NoituKyvH5T4pK3ge
bWf8b//C/9p5xgzSz9IyaSi1NIK745vQ13w6Fxc85iZmmeXH3mO+cmdShny9UAnU0iXsqLdpBuwt
db6fJk7cQvgM+sDI2ZVcjWh6/AsZsJVca8KMVulxHEWI+/kgQnE1/THP3xyBjaR5IXqHersRsa3L
F0ZxJznV3/3azDJl+quJQNfYVtndLacx5/eV0GkiIWjT/ezgnCP1a8APVi1yheRQecVjGo6UCcoL
0TJ2l6mC7MNR3n9n02WZNdRDRXOeGB4AhzVM6fWaACo6diTukBu0rksVnxOaH2LnlMt8axcnZp8B
EyK5ulONIozzHCnjTT0DrhOf4JvXCaq/2awJgnM4Eqv2eVusyYWF5ox6p+8U2UBxqtldx2ufEnEm
CFNaj1n+ExZR0CWq6f6vYoiNGMS4Jbj02jwwUe7E5Z3MBrEqZyVXBW4Ii2Ff9nyNTsxGDppTOHV3
x9ChgLuNNlKDz99F5unCxHcY8Ut1rFunYIcO+GgFQUwKt4k1Wd1LoisYMFW3KsqlnpzHgHWC/qp2
LKdRJxcTnOCr209sV4lCwWAl8CWfPVkxwyz/t8HhOlVYeKKO/oTq/B6nYi1MtCfEmsv/VPiV8zya
Ftm9zT0feNSCfHaC5f2drNw1XKRUBevQtlkIoGj0CrhhobinooFoe7RDNt/6HbT+KK+WXpSOXp9L
H7ct4blN2jgVwXMAH3nxVT2y2kxPUyC0xSCISih2h4YYEMvH83HAranZcpVtaEoEsFqYINwI9gAo
uTp6/BcrzM+w/42DFzik93ldvYfisIkHsFtgUfm1ZE+jbpAJyX7vK6/iIRM8W6gUC34E4fU2A3oi
Wy56mEC9uEEfIwGP8cHpuOkp+gLXTZls5/idEXjInivZeoNw4wF2FNHAeHO0+NQyTom6lLB5pXm7
XMMrPdicqyOvoPWcTTzsTgC7/zvVnLTu5oBAULlEB80HtbfHBIgGuC3S7JrMdTRmMk5cXp7QrJPC
hZTuavPJ5L+ULhbJkKB2LDbyCSzFYK8myxpt7uEcTbcVQf2KtxtFXPH4ZOK+6BOEj9xR+1JhqtKn
Ikvn/Sz25I5xaToh4Vw+4TIqzfeRYxPAuKNwUlVTMEcAcU1TAb1F2eI54dGH+ky1LXjouP1rWlpc
mBJC2IRC/Rg2klNPIWqoxL8nN0/7KexZAh7qg6ySDasSioClGKQZVsDtvrtUBhqL/Wyh4BRacjqt
tk1DRWgtdy1E1eny2s5leuwLAke8al0RdGTONDd9voi8AM6uNPdR/nJC2Saez9ej5HM3zp+uQOhk
L/9RPpJ6mZnptbhcCC54tnY+8fU0m7AxsSQPV1Hxfy/0zk+3kvd2gcipnvjC395as8IOa6tr2VW1
MzGEeXYy4o8Z5IKrXFvo2z5+Qa1jdvsRBVcu3ElE6d7AkCJ8vRGKXe8Ey7hwoJnmeEGUAxoJ7hp0
uDXi6ubg0zSt7dYRyXSbyx/Vx6f7m+f9zzdMRoPngiOmwZ2VU9Xxa2kK/SBUh1kZUn3RpFcRnNKH
Dm1XKqPuSR5efoDugTEqgdb2QyCngazwiM09/OMTzLVA/Wa+qH2OJlZBeUwvkULTPmJmgBrC9wqs
ZxFKHaVVqL/Ion4goRseZiDpNmTt7mb+S3R6UQzG670dsif5JVZWUw6DiLDUyH3yZJaiOC2bgmtD
aNlqV/HM6NIfoVI3Hfhu/WfVcb+vP8GoAW4c5Jr8rx3LxXZIc9S3+7Cn/bB35XVSRcH1vO2TU4Vy
WiMbSnZMMKZtVjxHpvQWixEujHUbju93AvKQhAnnkriPu1xc0QxY/IsLQPHjKsI1Yy65uDS/bLMb
562ImoN3XTLh73y8NLlTm0GD5gcJlpt/eMlIiEYasOi9J3T/uJhOJ12Wa70+ktAmIj0oAvC6B2os
Fwvxv1g6nFu84pAMFjSs55yobf9QnpJ5jO6r0vt7RJDghkv8b96NkL5lfTYG5tBwdIsPcqyXM+u7
sdXGrxf6m8FM3E+F0IRly5vDdCq02CarkjVBlHUoaRzRf2oQj0yAaje6xbJNdJRywHiB6+rTigJq
UrwPmAdT8dWrJCUgejD7ufVZFJv0eo0l5FZ2hSycAbYLU/HXSsn3x7iIeiGDtP5lh06Q/SMNfmG1
idgE9dzZ77DsvKvbKaI3B/kujqvLuAjkkUSpIpIs/RzwpImLozTbu0CSr/+vrlLH/iFphyVmllG5
pmUHZPcTg9HILRLtpASTLRqj/mTj+2ugrxj6ZCaAbGe4/2p7bnbSGMv1VQMblv0ePfiYzx8SBjdn
pTmH71Yr+rtMT+DOEg192WJyjm/I8Bjo9ZsO7NmENKjyDwlfeTa658vohBc7bCzWTou+Kr+vYA3L
tvMil03dMB+EjollhgKW0Vgr0BahMvomLi+rnQMXNCgcPULW1IsFImwtA6JBZwdhPPrJOLNgGzBG
HVJrPvFwMCGOqrMgFEgGg118yWKZ3MskL1Cc3hgPcIqaD5z6dvWWUaHRCGjJ4dOn+rZT22tM2n/U
CU4hbcK3XSevR3/Cn8taoCDXd/MDZTaYX4vYoA4vppUeny0d9FMSf0VfR+/auH+wHhQb4DBmhqTk
JknUj4EUsBwmddge1eUTGJhleKIfrf9clMd0nC0+S97fcsesroOuXGWvc91AnmMahMESmPLwJYU/
4qPooVP6fmNJodrSqHcAn6eJx4gIakKuyKSnXIyUK90uWOkf1jjmoDWqVWMDB13dLEMmWzzgtVC3
ZECkKffzaVkaoEkR0YXogQypedidyY6qfC0jXfzlrN23XFELxWOUsyaur0ZWWo00hcSSBQJagxpz
lykA++pmvRJ1vpkOX5B7xRz2nuScJbiVaCwH+VUCgD7Zry5d2p6KWa6+p7dl7lwldjhMKFUFXhPr
9wckWy3BBx7d1rO20avn8+R6RQmeeiYCCMMsArprSkWZfK3wh3FzHvhbdUsIlLWVUvG8x4LQmNoD
a3h0bsBj+r7BgZidgBiH6PozoYPGsfjefTTR7yv8eItGzD48X9UwU2xuE2JKIjJjyLOyJrU1pLu0
XmzKprkkXQeL+o2EasO3hksGwn/T0iBWPMoHZsN+8vOg7OOeTUmlZ5Pz+KJkaaUsQ8PA4OvvwjQY
kFngZ/lxQBQrL2f5i5AgckN4jf1ZEuqs9DH6LHkn5hUUjUMgRCvKDGjX11ZNwiL/RVa5///wC3AD
lpdzWuqFa09Z5+BTg7RwSH0Nv6CutsJDXspdHmcEFYUa4CPvVNzixwENyT0WP2+PFtCyIPY1EvDX
z4kkQNlT176CltQNZmQvbJ9HCmkkE4CF9Qw7o/wr5ucYrDTKXtdLSCePGip2JhxLmyZqlaLEq5pR
Dxy/A1fs0G56itFY3qlB5Cpe2hwjTFLgnNrWb9FzXgNIiwWGQvMtFLgkvhCu2kdSZcTAaky43lyp
/tyn3Qe8D5lY1rG/vCgooXHrwpUln/TutHcDEBZoHX1AQ/5hzjcjE8RUqWAbPldoVv15aj+a3oCW
ZgiU5mVPsAUdG9QqyG2yMPgLvlGdquy7c0rkwlAP0iUBIOWT0CCkcWQYQZk0pa6LyhitpUnc4oMv
l0yYavmc1l4cxPklCM46ZIn0qg2XHhMsAHaE6E/1Qs0Ec/cLyc0FGcY+OFgrOrn00cUiVRsvtEQa
3eYg/atFJ6wWk7fMqKh83O81YdJMWQSJRF0G3IYTMa685WJ0/gWZo8FSeU2+MhOhPoVmNs5t4KPc
6fd7QobFzuGDb9y1f5OsHSufTI26FBnISXDwYC+Zg21R24qMO51YGUAZt29S7HYOp/60Kd17qz5p
4e3KyzycttTjaHh1Z9QSB9/m7Qgk5PSLkRPgTnz6llzIsrjRTl1eVgsfHI70FH3e2izUEq1+vBCM
3nTPq3mFkECUObzYOLk3Uys6wPcvDrqkbZZStxettHct1+RNcGGAXL9NPG7boP/VvmqLa1xVr6d+
vYaoqxjswWFIxUnUfeQNM9CuMg8vZM9hptaS9e0utcxDuDk0kWosuma7zXE1kYWue32fab0dGcog
NECqUrSkGoSQtNDIDNLLHK0RUIMD9sUXLhlphl0yWFongHNwBcQMzejjmcOngjA8RtlHMkIuPllx
YCDM5KBDPHwh1gFvFkw8+aBIqC4gsHBsaf0/o4RfLHSBpi0QHgbhY58tfpSvQd41jKDsWb2Yw4MV
z/xwZ2fNoaYq70CoNKYlZ+O0qrorM4fCprueYPrykxFT6nkabZ7t1utMQotThptM0z1FrIK9QfWH
PEF7lQkpwImL1TIl1f8XnYiNcccT2WQhQE7hPeML6JYnL9JtMo9+ZRrnHZHG/OMG7o5JpY98mjn6
o4cb51en8HN7Nnlw3wutRXuFpocpXFVGzK87Dl5SmH7K7ftRL04tRjOw9XnU7yeEy8ibgYXIthzM
hg88WVwJ1n6W8G43hXhdGCDJKbh9bYgOF1Sh6kV8Gp74ysUNcI1kmTPDHYpiDWCNM/FxhQlKbD2H
sD4xeh0i9hoXoHGEeTzBPt7EB4cdI+3yEjYOX3/855miFjq2CIBaDL3WXV5yA7SYfNke02eM1r/w
CkO03y3WgP7ekqtF0uNclllP9xVREzwmBCCgvE/npWD1vx0jQvVp9ybbkLj1DcS57M9MpBGoqa7Y
xIdHiLZrLHEvHctHJAiuHaW3HV8goZPc61o15/A1olEfxLFCU2Q8CnvQmxURoD6JcSvlPYjNEOwx
30KBncBn1uBtoC6LirL7XEFn38xm/uHTHm3CxL2b9kFxwNn2UYgTsCFoDcYPF9zK7pMznkVKnID+
xns/ZhrKhW9PleKp48f3Y1BRDYx06uEOLLbiCEW0jVcPcaTVpkOQ/kSDgqI8EzWqHHC8mMXlBfDn
YX4TFW50fQOw/2Owfjb7yj+yun46bBq5WCkbF5+pi+MBSOe7HZTCwNaD7+RoPUpEomBwO3guXFI0
YBOBciJn070uBocySIeF2vpY03wbFVhDIMu/tPDdVjOzhHkovS8hJ6TiqpEzuswCFnU3GBzhhdq8
oJtcmGh7frSSiv+ConWYFkanOSDoBsgjfkSvyd+zbUOXqaHxRgIcdxSdQODECMmCUY0zoFUp4EBi
gEBfAXfJaLvlDc8wupSZ7v4SaCc5zjTzRtYWD+6oyyahXRRabo655GAcj3vr5kGy2FDSqmbYd+Qt
JoeCBJUDtH6BIPoCYL7wA003eTtL0x5uThWGnp3vi2WMq/x4ybMnmGVIZmLmv5HJH8VystkrVm6W
w/sBCz1Au5uVoFbYo3MMKC5Wsu2d/GGaVxXgZ0r+vH4NFoxeJVOAFwnR3+p/ew1Ad6LC2TPw3F4L
635kaSbEY2b12TaAkRajjWbamAbHNUT5gYtmGT4y9txCLX3ErDlkBD4Lz9RlSvOW/xyslXgHMlhK
QOJpQu7+inx4t4qoBhQNyDXYegJDvQpkTokGJb3opyuqZIFgE6/eQgXMbk9+Rz0CgNC4I8QG6Fqg
00ng2suGYw5SAKAYvjP1C6QweZqfKjjcbJbgDGmmftQa2EWfHs0mfqJuM10DUpfSQi+54n9nMN9H
5u/qIxRLAxvKBOjoSuHde7Ai9Sgsr5HOuqYZwcrK6mJWrA7zXZwzK7quJ5XtoEW2tLlhsCJLAMtr
yXQunbGy5+NCWX+YZB3XM0djmKLQSW7rnh1Ar15gyHnBMjMI9mO4wV6q9TIFXZLqeE+ltHsaFDoh
It3gdp4zDbMerZJ0aSgHTVMPyq7ZxCuRXbnCehJFVuK9x8n0Q2JaPiWFHE5rzETc17pI/Hd0CD6S
WpB4QdAgksgdezZve+DnD/zI8AIAciqRulBEh5p/FBYl6BF67VNDCP1sMnRIGkryNAhKVmn3zcxr
OMVZxOq+LjzfoWkYFLOwkQCYicFth83UJj2cMUl1s8MBhRIo5ePq01V0e/8dVxiYJk8oH2XrVy7m
o12LI1tDygega5dXek5G0CymAftFcYfY5vbcZEYYNWrBuAGpgxy0fOgvpUnKBXHWP2/GpIF7x3GP
ymDBFBumLyNmaapTgXawdMGI41Dh8LMhQGoQh5FGSfTjbmj8x5T3wjFk5BXetfe6lp5Tiyq4gzwM
CGOtuhGYRbz+wuNMwiE44VnHxKi481JnpvFi98s6XRAYQJRAyuJmvO3YWSkAppsLD4YiZLSIES4k
P6yQ370B8wUDtHSHZzx8GUEnkY6ZyliYDHmQmreAfTOtgAweOUpCuIoVsVuwp0q8v3M/hm00shIv
5wwhUJVvEpAK214iZQVpW8/Q5ewKM2WmKewxuBHvYb49oqmBp+LcdjxVOuoXjhDqsuvUyeIZ24BX
l/rBN8wu5fWU3rYipyJlJB7ODkWBub1ZC3a36aJJ+7Q05nFKRm6ZJfGu9AloDkcmdydAdL1kmnUO
JvIwKI3l+pu0NpydU6M7K0ztyUoopDLCbgxVBggeCq3lmvySnx/30w3evsWNi3uRLRKX5SjNh1AT
JvLZcYf+WOjyJVTpyu87vwLvoHWPNRgwQNd+qeqcE/XZXjNydvuBgZgnzOngVS19bS5mmkcegaWa
U5MYYeRB2NPuABrqK+cp6B7YOPrs6JlzEGfTBbfnb6EkqFYz7MEqaDFs4Hawe7lN1MsJrLvzWcE2
4wT2lE+Qy8Uue+BEWeYX9LGBoIvC2GmLtJ4+t8OWuiLyq0woq0SkUkvZUqv+x5Yi62Go92iv1wOX
GNNNGMWwoFweXvVQcmsXMh9Z/liYJOUIAMQtJ74DFmAc3jSk6V3juHfwheM+LP02R4zEjAJ7PsIB
Q4HRhNn0TZbuM5w69T/E/FkHxt+RF8x6+1AkCmGzRn+Ry5f+xR8EuyumOWb5SrQC35uzgRbkhnV4
cXtoWcUNoDuDdKMk6WrhSkrDBNI/DaabE7zxSh0HBfBcjFl0wRXs0vCCE5tVqYuIgHJq461xxUhH
TP1AIjLfKhXR0urxVgw1/aPl5d2Cy/wavwZKIA+G3LLf+W/TIOBKVHkZ6FTwM8sUYRMPrv9Mowr9
XazRh5JJVzptYwbEBogaVOTt/rq6LZK9tpD2mRUg0yXF2QalPAbE2xcEEPTZGxK8s3pyR5isd7uL
Cqg8lMUm//CgAgdpEkfgJ9rODrBMRT9bWmQFuawmGc95SMC6JJHxBR63iT+NsVq3cdSYeTllxsCH
wR6XAD5pVXo+IllqF1oYDHyGpSuJk3y8krCpkHZohRva3iIUbl/wA92giNAiVnW2hiptU/XiGqha
GMPnI9CWO+SM2AioIA+kPSHWJgWfH2V5DpNKy6yJ6Rn3HuWXU/qglir8IiG1WWZF/IhHtUXoXz1h
rXRsXcJ43bHzMJvg2jGu9Z4ypEUm4AWqgJqUDRxIi3JoEHzebOniSinLxY++c+3llJei5twjX5W0
zIlLeZpdmCGTafhKlr7/seQLUNjybUOz8AgtnqRclitxsEME5Y4gCa6+TJZwi0z925gPnxSfZAHJ
V8WMlmJO/DzHWUfHtGH9Qk3qqNtxuJqwkorFFahAcpU3HrH64hGoCZO44jSCIOMH3a6fgpRAHFTH
sEbDNZPDqbkHKqVkWLF4cao5LvPp/HUD3xTwYkN3PIt8MWrcMD8yIyvY+foNZUhvq8SlF/yRGAJo
A35Z6ZH9+dMCTfySzJYsYxJ1qhH8VURY+EaNFCYZqt2VaMyCqDv5oHSf5dfTkqqMXcdv7I9wpeNa
MlYBNJI+xtPgMz4guVDOuBf4RCy0htWfEKuXnV/kOTqdUikrxNQ8MSvnHaZCz+fupwWrF0vv8yle
2LF8tAzfVRayli1+N/7Q0AjbE9xf0JIiCnuJbSVpYfdnPR2mSXnuKlFTVnoK5k5biW1F6wIWoqyQ
lQEmcj6+hlg7mxEHAGFAceyxvoYVhmGTWCwJxpqLOoI0MdGy/oT7aLUh1EGQH4xr2oI0lbBQKVAc
SKE3iNuHDKABHXehkqIMPzgfkGZ0bs9bti8BNa0UICA47dB4ZQV8c4W+VmhyNeYLw0XxeWdZm665
0feW6krYGaetPF26x4tk3l8woHyy5q4aPyXmq57NKmblKb9EAJ4oxOqfSCMCkoMKZej4BsKBsBG0
USa8FCPtO30+/f0xk9soygpfA6TAglntSjxa0CAXnPa4AR/iRnVi3UhKU9OQqsws/MJQ9yypuPA5
WJ9/gtsi1ZgNlQw+HU+9gqPiwU1+GUaOoKvJgBhHkRsAE1/3Wh9myPUlzfyoC3o7FdUrALTQT+iN
FfXYI3zqSpCP7UO3jF4/HLJ1aqHZacVMPooDjtlNR3sBeLgFfPuyRsl+HfHtJf8PrvPYXBaraKOD
0NiQlULxWoew0W+uXj2O8KNtmRYbtID553XYBlT2WqypIrhDvYFMcJ3axdWWPCSBuESybFqAjSuX
jhmIzNypqBojnAYWmYtIoKl3JmmTKUwlIMqud17sxTg2GzebpD8bYdWB7hoxJdPpru/NIX8QkQLL
zT0wF+sYOq7kPHJGpIr6mRXk6cmmPviLaXxg/9TaB/w7s2jUFHREHSzed4zlhiPh4bh6Cj4soW8S
gpPjgVUYMIrKuzpT//4FyJNomAENmQIWYjQMyGKY5JhuNGxNnF+K+NC00aKntvLCbM98mUCmSqey
p1T+i36xH7KZtR3fE3a8hmdPC9d3DHP2OtYFerwl4rDNE44K0d2W52KJF6aqxm7D4lqB6bYkfAQo
+G/2/g1O69EBpBSK8bQ0fYXeuR4GmrSrjJbG+diDxubzyvjTiEmyYdtLW/b0oFH6QptTFP5P/HKJ
VmZNITgRrFiHr9gfyNGxzwze9fQ/vkANRMdXKqhJjFz7MhXolbbRQlN3dbDgC5z7lg4MPwONMyLu
lN4FIQTxrlbbr/qEhrFiR5CvjFzO1GRydua7scqgjqnFpfHXxFkjUfxcc2a+hMIWZtFlUu6J/VOy
T+n4ICurluS1nFR/DMbRFwVzskxCFlUeQ/jmhaabNauaF8DQt9kKp+LSvVYLtU4LzAyVNj7TTKmk
ua5IvzW8jRWMusBYjxLv5NrN7iSbv9sJOmOMSuNv1XJekyzBEOXBCqjdJLbdhMJgSjax8POmIUml
mCh/Oyq5n5T/2MamTARKBLgmqP8joRrqyUfgIp12Lt3ri0913tvFO5MsP0DyvwZRmeJOMwRZ3lqn
PGAXa3/dDWqW4FEakv9wwmX1sHvvgrridzRyG33VuAT+6yx2tLhqmzXBqYQXkvwV4xerXMj/cyyz
Ozd06fPKm1sbWQcVlXi28jpUt7SyVJpp0bRY2oppc061jbD7TCjUteFjxNEpTFSsSXvHdL0eB0Q8
G1DQBF+1VsOR9iAJVwJkD9PEwO2nicvV2YUvYhZ/yJikkJdzNYmq1MB1VrsVpf/hwVeU8Wu4T5el
1b2alJHg7yU1gE4HBLVCtXeGJwgzxs91IYwRZG+NQ+0hFEzuKj9iWMZPY/duuTXwwiCbscZpdrTz
gngSIKg2+Lnae5vfYPjYKCdYBS1u3aHnQhT8RTUTc/6G+sYsVVYDYXrA6leHH2E0h/JatfBl6AMU
iP2LWvqiifNcdYDlfBQiFaNijaygUVaHEk7KYYIF35iXekFEca8eOWrLQI93rfz1ycWQsXOeQu5/
TgXcuIDJGnG8BGWhMAPqzlVrThJrwYNk2P2YtRwObL++xQF0owf9IGQL/4SKy/1Omu8RCjTh4PBi
2p+/FfZln+rDyyVPK02mLYD+EduN58R+BDic1S4tCo9LnwxtEH48qSqicFq+WDKehy57yDbMU8DE
u7Kllad2mF2k1xjG+bfhXuIEhmE3Ofn1wKc35HEi2XJw3j130ellAzgZrZgOsBlr/bGs/LvXslqo
KxZQRn0YxnBWpC8MTuWULkV2hn+CbZCGF/tLpRTKZLYMb91lAbu6V6au267cRKVSjmpi3sfLioZ1
6EeMHcQT3mA1GkTGMcsvu2lJnhnTEr+cs9dY36r1Yb/SbYkqpsC5NyPoFUl2r9gakumTjvjVwygQ
wrmDRpNLPFND4ny4dGsPNkHs0mC42bL2tcMfUW/pkelNJZQbhchwLGIb8NAfQigmcuuxtnD5gumQ
GnRaVohGqtCJnEYr+tKs94Xs9/N+ZcFzvv0YTvbp9RBA47QVVMbWVT8Kes/q8mqt7gBL/TwAyPoa
WRa9oqYjPd6c78xvEAqJzfD252a0d4qVRNvOfA4V3UnaAzyElLf2nKxe9j7ocRu2erjtwmDVmKfI
RLz5vbTrOy3TEMd3H2qLXXQCCtLfx0Q0T7d39eONuabKtTQf/HEqiyme7j9TKD69vJn/JTSH3zlv
sfQuyMriT/xI38wDVLL/KrrIE+ibszIXVblPrehWOSU8O4kZrSOIR2ylbCfps1JPf/xOiE+2/QhA
WzucgkxBsN5f0Dr3vcp6aZrBcPIKrf6d5fj3FSb8k4/h7saMmFAUe2OXpcWZSy6g8MCVm1aFuc9w
GF+iAEQ9NxTTXYYnqC1sfz9i9z7WxMR7hfS0HVXbhzBByBxXd43Oz9x5lSLTgP0jf135Br4KfWaK
rm8Bh/+DBGF0oOj17oNxJ4e5/EEJkn3w19CQwA9c2vj9SPYeSsXzeG+6C50cGv5p8RnGR16KGIpQ
Bb9u3pr261W/wuhY7eE8UsFA6uvvYq4fhop8MkRvpZky7VOL0n8bIgjz82iPxRPDtgJzz+2azhIs
+okKGhMndmfmQdsA0MZ2bVJf+7vUzPb+uK0ME76RnZDo7m+7rvgTYt4PMUB/hWvnNs/b3nG6uOwi
r5Akh9JQJ9OtzdrHVBlxQYrpiX4DFb/XMdstfuTreEMfMCSEiGgyjUhcKPES/dT1tQ6U4fssKp+D
csw0/dz59Z1GuSsz0f27by7AwXxcFog+EOtSur4lv7qxuTp0WsG5Vynzq9eMwwTt1R3tRq8TP08U
Igqi3UxPpV3TJxCib3cbhAhGJlk+6c72XPN821rMgDqjclhrEblwhhPrjtFys4U3A3vAoZcNUARC
FFHjOndliZpCu6G8eFQrGxfcxX2d18oloK22KyQ3F+Pj57XH+gCMjuqgy1/rortVlG22UbeBoaWy
p5wUNrYYhkdSVi42ZZKNSJcafPR/HYRsycT2UrpQM/DG6ehRNpj3Q87ldiidTqb/fP26eWrQsvHS
MtWHnq8K32lDQEh9flUJ/QrTvPWn0Qz4prCmgee0O+QGu5dbfkoIoysDa+lEga/O4ZitmViykyZZ
pQUXLwuuOoBYlXuK1AFfytHSMr5I+6lz9gZlgjMKDChV3nOA/gLK+jTzBlE6Ip9M/nX+K9rskNzi
iuM3bPKnnqHqHHoNoSWrZQ6dVRwUOQE5ObVghmXt8u43/aT1IQ2iSFNpVSa58NTsuuVJZa5xxplm
JrWF4ida1vTl4mDGHi2aHg1KICBoGZmsMqjkj/86Fi0DqxKYE5HDxT1qD3xhNuLAVfVZfYNDfmz8
si+VBEQWN4ezmMPkQH+JlYF9Bnl79wEKj4ZllAgG3F/NkXE7NkJNrFhlXa/Br99SOAaRW/eQpkju
i+y49n1ffmsjCP+RC60he7tfQ7/ay6/ezUREncLdfkHxW+C5qmN6fG/ObWZb4f0lHLqh3LKdTVrS
jymFhi6Xbd6F7xiLWhhQIM4cJHwkGTjErK0ks1QKH5odkLBhSq8ilzEXrPaB2Br+3f0eFMYglylm
jm4ymyV8QjFdEWeFQkpx2lfls7UZksWch8/AyTGq6tLEcgULUi2NzgMKZytpToIs8nlpGqNmIbRB
7cr47DcAYOQWZOTuPNq1zx+ReFqrDgsqDmlL8/mtAaE9J74YQFBQHwU0DWOqqdekC9Dln2kT7JNz
j0+7Nw50bxykvEg6kj7NxblK57a3YvKNz6/62wGIDWSHYQ37kloo0IRxanmAj/kErs/9WHbTwRgV
mCZ8ZYxaxbk8fL5a3bTBY2nV8qBQvuZ8G4C6iCtzk4/Kuq+TkSOmhF2QIR5Vy+s292pxWSkdo+68
wUxiUOY0M+wpi3B/UKOHgZHhG5RRRm2H0w+7RfZ4/ysdIQw5KBLt/hmjGSYn9LZ+w3jyL8DtvPUe
1nhq9PUhHf8o0Gjv2Wpxrxt9W9UKlWStu7yq40Wgyc+5nWwy2XO/FkccUULmktHA23nHU7m+3+mt
9S5bTRPKzJCwNbBN6H4YDPyphZGMytiQ7zmylHe/rRCIv5ZoBrqJVruh3cyF/egFW8wcoE2kfrGK
7WW7aoqfP3SiSOHNSIaLVDhQX7JtaiuMEn9F/MNdhooj5cdDLxjvNg0G9k0x3V4bV0YWG1sEu5cB
mBkJ0BDJoHwiKTzl+vzBl8nNjd3xQhwYUzl+l/Ja99t2ETwDmf7uB8+zDqLpiSc2LtAcpwMKsWvw
jx2XleZ+V1VqH6X/kioEVCHTVeVQM5K47vzUP5lfacXg2w55nNRRXU17EdRpTMhd+r40CaXOzCo8
VczBQ7/KX6//3Xc55/kdDyagvcuFViv9GUUELEo+Mc/DcshbZb/CPUQO/Ja+FtzMfRcLo5w4UzNo
JliOjc3rt1zIK+3fk/cCTbkqdw+6MAz7lZBLk80mKp5UNZiLn5+GcVu4IAhIFf03wtdRwy/gp44l
Te3Up2EsPU1iM/QO5o/APpFPnyUagOBON2a76UZPZktymOcaAsRnPFQbplx/j/KWjML+/YmZZawr
cdp6s30CXRNUAtvYH5x3KO18H90D98PKySicoLaTGsTQ0qFiXcXzPCUPXFc9PMWuXeENqvlZr+YF
8l8yoEqxMRoeXDL4dOc+nVAnPJT47i6AOwHxcLWBfUrGalTUvIpZwDJmPdUsQXsTrS7+jFA4OHFS
7uUzVifXpxkUYIipB3/LOImPJDyJ6X2FRWEtgk1en8fqZ1sjrdoFVuFi6qhL0TvJhOq8Hay1A+ZZ
3IxvbYQYk5F3YOaokglyudfGc7m6yEeytOHVIPPj9mYyNYxdQUIzVpYv5+Lx/amdhz7OmeNjza05
9kLbvB6+IuYeJKDdxnXJkRACsH1dF0mClmTgR8CMOncy5aMjnCLcWYQPL6vdVzLjFSM1mYFo8gPZ
ongK3yi0nrSJo7F0WxECUyuuywPWiHGpP7fdw2ggyxNwMirH53qwU7TEwVJxtEM4NEPZJmEENqmb
2QE/TGRsnTcp+e1jU/NWqY3s6eOePaC7xuagNUUgy50oA7owWYXrsHnHU0vzjJxVTzaM2bsca2Bh
2HTpYKKJI4P+9U8LUgQzSnFrC/lt7BS+DHnGryBezqLESnhS0DSNgPvdtVxJUaSR/BdiukEig3yQ
Kj68sw4OvYFOvLq9GkxZQRiL+7si4tb068kh/AKn1duW2lTBbU75WvJVaJq8kvuhkCPWZb1U5MJN
hXUE+C/qmb4++v3O+lwSlm5F81QyXjRxybOrY3JwQ8G6d4mBfrFeWDTByQLp30ysGyqb0geGH30O
ZA/nAHFgmNKnFa9ASWfpAHjdo4W2MklCfNCNJ35GoW+EjBRit/jP4RaF6BlsFblzE8Clmvc5Upu6
d2BzlNb+5PcGx9sD5gh7/hN5BRQsB8QSjvPas/I0PsrsAFZAwduNIDyTFF5U6y2NF2YdSmbH0U3C
9241CLD2cRNEcmegXlWhM+b/CNwmexFC6kp2OoY3C1tumvzYAiA81U5NHkfzfekxTCacgsPKfNCa
UF8dsKYJOqk78tS51VtrH0wCXK5gHlFeOOpHnwBwRxrpuSKMWtV4lqIexGDfrIgY/yOKfHOFILr6
lCYNdiVAy0qNxklmvu6UDPPoJRSJSK6uWQlgskpco1FvFPlLk2xBtMWmrliH/nP02SXwXBA4V615
b3zDir9QsYBc9aVmnh7I4HT1WF+RaCkiumZ3w759Je0O4Cn3400MLnnT3Vt9ea8/xSHu+T3cGNeW
Nw50d4Fr+80Wta2S1tfvSGO81bs5FIxzgmLxy1N9yxfz6QElTY939VHxGldgobiv6rjBcf2ePsR2
HEqW1smV6vCUUd4IZ5teekTmOF7/kWDkhiaiFiAGvC+GHhXhNhasTKUbTiubCsb8/LpaCuPba3jb
jSokI1VEO4jPkleDFTownDl9d39yLNFNU1NKYgQ5KuHZgH5Fk73kx4O4bblSp9Q4CbhvRy3WD+CR
lWbomjpuYqDAqLMbGd0qXyuYdweFBkzxgTdtGG7g78uMIsJJv/NmWNTLoKH4nsi5II+FdApzk4P5
lP9joWtn4uAlVEbB85rQloHIxJwx6JjS+vjOWfK5wGkDz7VKTr6g9lctHkHW2csoGPjJ1MytSWWZ
ckA8W52z6DP1G4QP12K/bZon5Jc31noEPK6f5WyoiESNb8HUK2TaCqME+VvD0G9rVpPk/BXhNVjx
YjfXYPkA7mSRWkCh8EkHUetH1kLalea0qYvTn+wbZviNE5J6sjMsI+HJa6Xyd/6Wj52BaI41HsnX
nNHLme9Pjs8fbYJcMP8eMarbh31NE2khA0vBH3JhGVxEzlA/3NAQJFyG+bYXMvF31qKI6oz9kxUE
cldVpgXMC8w4As7kxlClUHPTrwLtmfwJN4SQXc2vkSt6qLP1Uf3VSqQ/5B2tEL56j7W9LPL61JN+
w0tPOG9mdCdmHcc5FNBwhN3uLbqdOTU0BRqVU1POh6G1TvCgYfCe9PwSvGc2eO2tfM9OT1SbQEkU
u7kBMrrDibbN71ZzzhY3Ze2rNMtfGodwBlB/PkieZyI1ecOyAYMAIbxK1U0kKFiYtuO2DXHBU/yw
1kxaALtxQfbhXgVk3hp11nDQeg4/VZvvflUIM3EkxSvQWneuf/I3fp1YSczVjb7Oin9ZZs77idPu
KtYGol0IIiN2a4CR2EI0IuFJ06mafb/FXvylR3rzB6NcB8kXte3dq9FQ67SQ8guS36fdzgXJRpt5
7vE872zP84Q4oeo0bs1j0Bcl5u00qHPtxdQ5oQ7Dui6nCiCLwdbWUJwLH59ujf2Ng+aANeWWEVU5
aQa06YkdbxafjCWaueaZzYqtSiDOQx/5PDgv7FJ/6aZwarPtTC1WCtlZF3lPinv8FVnZO5XCTKej
fgZxY+2yTz+YW57ngaCUmAt4KY016xr6huULkKqy5Ku6ZnfzXcrC1EAchOhKvsMjVVSJ9uTAiVWq
LLFfwGzDjEgUIcD1sg5jHBBNGrI/4xKdDVQloKnvcfkfa+/R+Td1glhuz3UBWOJsn8T3xFUJVxge
ic3/CDqx1ofvNnkNbt2tKfafn/iLIHikaksS5AMXsb3Ux0dicKeK2vxUS+LZXaa4HmCnY5k8+DKy
QtO/VGU8/Yqn4p/cYRI+GwmcZCPq2STRts+sCEHFF7ZeiN/H8zQZtB0bVGgp5ZdTDEPjYhyhmIP/
GH2ohFUH2RC2zXBCws+JyDb1J903kuwc1wJRY6NiGCY95PEFEt6vhUuK/tc1F+K0ZWiV5SgSk56p
wZc2uhU8wzxs+j9F3y88KmO7THD5QOxeD5s09Sev97hte2CcyRysTbf3N0qiTO+cxunwHP2hhT6v
lKmzB1aDZyzpqq6ZtjBDqIFgvoTsoUy7Xe6orGzT+2rUnZixbQLmNh4m2/3ruaDj1yw7HuENjg4j
unNQ6CXqLIdlI0/XixEHKzF2OnYsmPpXMrotxbgiFwkjLh1nlKBM3s22gkOzxyyGDGCaN2pGYeaR
zSNjBWXez+M9PbZ46cB+h+4tDXprlFTL3TN2scR+qy+KtYvQffbSvMnvmo7J4lCNogTqpL145avf
15Mmye4neq6c+DNUNkTj2FsL6J3GRHOGEbIjque056rFReiDB5RjL8EjaprjEt183VwdfWCsolAW
txLobnYOQ94MwFS4yGFYzNI3UEKoKvGltNdUydqoUfivvdsnmwwLjw0uFqmWzyxfwwZILIwwoVwD
nkxgGGtnAuHl//09tp8vbRQ6VPqGF2m4dWriHXqHtg4kQHjUs/zImTF31i8yBbiLkAHjJFNLcp8Z
HuEid40SdvA1xD2infzG3M6kLJuBwRLgIJqCiqrEwR8/oFeiAK6Oc8CX9kGMUGTnOrR9wcQ/lxrc
n4BBxuCOTukO6m0zWMusv5VHh7nfnXt1DAF53E8suwwwUOKdXrKkLIxM2Uslw5CnhhYhFfxgQB8Z
CaeLZ9jTU7NrLUgyrX3V9LhTQh5xcsJz1NUmzLQoRQBV+fj/i2k1HxAE2Y3g4wRBHjGG4QPlstJE
pEyiebep5SXeXkYonNtgslNxhG/3NWSLHLq8838vMYH8+v/a0m2MW9hHcjZY1PDtHrOlaSOS/Xzx
CKhA5DNwXdIjt6Sih9Pc6l90k7u+aDvfv3b5ezjeNUz3BSzj3aExY5OFWFnwbbJrcKCaF/aFETZo
VvWRZGx81gI2qtUOinW6YlufFQJuAHiJtiSmr9s/PNh2l2OXszU0RYkyMDIhO78px8flFOawivqg
G4r+s31Q/vjNYu/H8FE0NuUE3TinfU8eTcqFnoBwso3yAIHn3J79FhhjTE07loydgnEBjb4TaJjU
vDurg2ox4g9KUmv4MC8GtdCJcfy/+BByqBxmH4EvERpLEeXdiLp7dIxhVpPIcPCb7gH0sI3SQGUZ
I1lVBpywzeIqHPlHkaBoQStNAigyZaZTnaQJZbtq2yyvgqmPYdVc2xEkUuzvp4rXkIERwzrSwEuk
c3gjej3kQy9MmkDUHD+L8CoP8sEE43SoX0iC66oYtmOUfb9Ulh9qxiT8/fMj4me4xBSf5i9K0NNG
vzqwkg0VBrVxTobOVYVTWXC0SDx9V911LF7D7ko4o08szGOvTJrzxhOtjyJbL6aLLuapNL5qS4lx
b0Wfa7ME6OAjtMzWbgSnyLb2OSQARgo7OWhX/V2WqKk/m9vMGka5CcZ/pv/27PSi/h7DbySWc9VM
nKR80dcvvHoNealKjfmUzwBZiIXLaE+du9ayTc5xOFyBuS+9mw7PrQ38cy3ge5Y4+gK1zI8Ksi3g
DEzOIHBHrEJfe/xp0qkUzhEeqjJ9ZwBZ2p3VHRmhYf8Sxl2DKsXaqmFC4ZyxU8ETxvD4qZhCDCQ3
unf9ni2xWFiscQCXorcOT/aoSDhTgLJs6GOjj5PhO4rBTYq0YwFABbMZ7Q2TSsZvyHNK3RfSOBXu
kfjBjq02GbaR4KyIAhWQEvt4v1H1eHNI/nNm2/e+QpUeKcxFOSaceoxTNd+5aP2SsPVhK1++AtAY
cQtFizpOXgyxfPy2gjWg9+WzceJVZ/C+7s+oMUd+B76zl4HcznQaha4TxltJFCFun9iUqMD6SlnH
ZTKaR+cnXRIqp+GMn4J7E0ag1gGuvC739H3VcqBUrkZQR2T0V5D394inxoF8lGoQ5eeb+txWll7J
1GLlB0OUrUKLrBi8llvSHdo1ERCa+LBTwv/AuimZ1z1/hsAKOwlRTYll+93VXYV0jH1hDM953pWq
Ao/ZgIE2p2mUrgoj5jSBo4sklguqV1c0Vurd2oAJK/0O7EqlAeMO6i7mti78+QGHcZAbZVssksv7
+yyxxHm07f+nTDwFxnvTWhQWKb+r4dI1qE5LlDdBbolxwe3wXRGS+tIxw/7h2J7a8gNLkNm6CA2Q
OWhwa6D7adu8eENuV4X23tLEw0SWMylB2/V82ZtIe8MBetxEjrZKkX+3SuYy8ZaWwJfxgJH4Znwx
bDSJZD4V27sOYOdkv9UNU7/2YAbmTVt/ExcekfMezSCgWO2N+KsEXjqChFQGD4FLPcSl7LDjnp+R
kFFGb79wSbPZIEDG2RvJnWJwxNvZQ5+yIRiwYJYjMs+aepVW5CfmKT1gPIbpUqHYa4oy7k/MZShC
xET1FUImJ2pzRR9lwD+6vrhTQ1H+2Vh/CFYhRUn8JzN66lD7K/Kaxu6OvuqFzFY03YuBHY9SjhqQ
85v7ZSKUMOOvvqMYhnFbXwMh1V9esNNIWrBdHWEaSWDRCdXo+K9SCBCygxhmznoS/ifGnb9Mjkn7
13Juz6Fqc/TuEPDBGFMc8A8VxkEzDpmWEwpMJBxSq+mU4FaFmk76gp193ElB3nYhybMrfuDIENAn
cJUgLu0GSfl0KKZdQMrq870hsPKJLczUDzs52RSIh/sHurzE8NRYYSW7ux9CU39OvNQSm7vE24er
9Q2nSBe92La/LvFTb79wTRBDFYsYCxZVNihUsACCxHJHroHSbuzsjXePMoPHOaWlr2EUr1U3/Yz5
MYcaQPp+sKRdQAYEPc/9YoOnf7Zc3OnXdTWjyCYA+pK3bQUXOoh7/W3iLtE4m1QeF7A9E8TpS+z3
C8pDTP1ezSBvxAgRSsa6UPr6mFNO8O+C7PuQJwCltXSI4kACYedumeiUiBaO5aS9S4olwxYykl7j
y8j4sn/pYNNoeIW8/pyAg7fhHD2413uSv/3i+RWpwQm4FBxYS89VLttk8G37sjvjgXmDvFsvB6xy
NkyAtPDPjBhQ9DZSkgr8Jebh5ysTD5gS/5ldncrLEQuOCR7ZV/QlxcNeAZKSxAYlKDcGhHf+7iDR
7yqjNNi2UZArFo9rivI1fLlv7DOw0yedu/zVONpMjgLl/j/lY7WfjNvaRID1zHZPcIL6uQ2vPOFo
Zs0D6ldmycmyNMssuvM1RoMVWA+1oTWqHI1TIKd0KvJOW18+XSMZ9ptuv2twZ5tOETwjrWSgB5v3
T3jVqazicztGlzKNdcle9qI3MV2wUNOeXCZZvKbydSOj/ATF5jPJwp12Yj7okqxofpuDAIiIvX4B
eX6hx7RcA5lmRc02Eof3MPcOu65dSe/WpKWwnkExClCxf4hRxoU/bPBHaxT/dnVvNNSUArHO/zCf
tnr+C/EzW2URfSq8aFUfC0nqP1Kp0+pArR0qFwjSEVoGQJCRt9DH+gM14EmmZOGXqnDzgXY0so0g
IwcFEkkTZlq+YSxfbK9w+b5U/964+rMT2OcW7qlZdCWRkxs8XF10bj6RuCoB+Of/QESQfYa+VrDw
n+NKS7R7e4BqGT3EDP78YQB6p+IRwg7bodL0+x9R9gYGRPASeBHZH+DYYhs907Ctpgb/Q1an0wWj
OZ4XcDUG/ttwl6V5A9Fik33gyx+ayB78ThnCPON4yDoI4pLWlDZLcFZBYBFdFfJXWiCAvx2yC+JL
KZ0BvXBqkBgbpw2nYSyLcTi512XL0OCjfXtpIEk4evuSjo79P+4SmbCvZTVfk/BL9KnU8aMjwN+e
OTTjVAN8g7EtSQSwg0fhRbWEGyz+hJ4pEzydTuPmTW3v2AhKs4BQthl+BKAKNKftwWoi7lBLbgsu
bKxvIykymazTB1+r7w2B/UOPaaHchFpkZXcnzR09Sgyi9L4IYSMzua9rLYBP2ejF/BglJ/oG79EA
nGX7MMwUq+tAzFN7ALnPYhJU+Z8sw3LUu7ADI4xJvKS1lznKrYri/Sfy90s6iLQQ1RUUwEw4dluf
rqgHwqmouM1w6ZRsbsfY07DGG3uIIvBiPPwfZAWUsKnPKhM17JwTkDCtFYAYO8u5VpiXVxywon0V
U9+AnN2e36/J+7MEtLua64T+J/O++SL/F/ZhtZGtHo5LHcdSy/ppEFtg39wj7Y0IXQaaGA7LhYDa
6ckgVvPGTrSEfBFP/4kLyDaeWMY/lPqQvTgR34qAeYO7ib2xS2eDs/58tW65j0HEHaTBUiSCsqt/
LkVMebPnBhlRirBti5FxYucb7DchG7lZhieHogZFhxRuCjPk7I6f+I9ICSz5H8VtAsB8xYyg+Z8M
CoeoHsOdLCmBxeiKmxMK3lDumEr9bEursT+H62t3BPHbjNlXZmgAMHqR2aVVZnbIcYY0jQFE0Js9
x1NV5wmJKXrDtoA57RSbEvHMGMuer2Dzs4JC4+htuBYhV2aOuu5+xM+vsa1/8sfEvpqvOHUJ463Z
l6iKlqvm6+242RxbC8JNEO0+HwY5xGwfOdiuC4XmAF5U0VtIMwj7HL9T5II6OLdBuVDzzpyzpLrA
cyIYF1LofJ7ipf5sHZi+ConBitdGsOjZdFkXJhVIehdwkQwbUG68ybPzmeW6ii+adwmi/ZXpc1CJ
x5n6ZvR28MRig5BYV9GcneOCGvF1mKSAOlixj7D2W6DfCf4KrY+pTfo/2u+vW/SXlKBQZY/Gf1LJ
QudjpKmd7Y4LtMdCgm9Gwq+tX/UGKz25Zhf8b0PFr0fxe7+UfpWLNtLUQCT4x38ybRvTU1RDVxat
fEmmU+mqKrXvjrdJ23n7CdaGQBp3mVtJTTSyiL3JhymPu/PrfOL9ZG56ybrFP158XJ6YzJ7MHqNT
IQ9WdJ61ajk5lYC+BoaCl79EyyNDKd4cx197nzsx7gQa9cU4BXdp/wDAuj+5fa1nONM3Co+x6CWY
FOYxVeWNiXrvKyJEEinn9l+OjSOG8AUUAtL9oZfZg11no8blHzCHaPLNDWBg82xs0AKeiUprshyj
Veenr+AIdom4WGlF4WRz4WvW2a6u+ln+HpY/9YKKySU5bgQXDyvCj1pnFVxRMc14bVdWJ4Wui4OV
P+g8XiA5B2Ct9z4X/7/etLyJYr4pU66SdXSRgFRvDChu+hu1FqY4JZoUgNjUpWG6R2gtBrNOd+SO
iLAH35NJTjmbWiwpQxggetmHOiIkcPBKSgcTpXg1RvuDV1rslD2p5HcTmrLBRIVB81O6ifvntfLq
lOSFcl2X7rsjriRRUKNs9oZG2JNAl08ozwzM1o0LZG/PwKFbKOVID2GQCH9gE6k1t18QqpeC8ybH
sUW4D1+6xUz8KyK5WKAtvrv1fAmH4Aq4z1EzePLTT2d+L51xN2xpxK2nxX9IREFwSMj3+v97zk6E
o+jlVJR69I28dbTdOHYcvQQ089I4qgjDay/D1EIk8/PeT/Q0m+4BQUrcq9tfixOpJ931bJ+fu5F6
CSFlzf9pJ6e9YhlO4LItrde5uzxelWIakFC1q9/+sV1776OOeXidGp+t+JEphQxTCg/l34WZ6c+B
JzzjJG3Xf9GyyclGvGFGnWtWlm+lDOaf+2S2rkMvGUN/PSKamQvYl13M2wuwV+zklAcpygr8O18J
ld9rHGpOmmEdqtifR0yLiIz8Lbk4Xc8WJ4eWNYOBvDRpDds5wVpzLG9U0f0A1+SiXY7xxhjFh0CI
Rik17PgX1elrLvzLNALOMR//XDMZasQKJygW/WzQi18tA9FHKu/B3sAELuyVsCymYl1tEfTFQKw8
MKs3gFnsehusHbgyZJg6GigBmm6v5HWiKwzle33egCLrQ881n2h+kFhEVi7TqAwP/C5XvWawEnx+
EoeDY3wVb83tdZIPgWPMfvrbg7g9Cxjnaepgqd60TEKF0XIAVOUZQ6S/E5MesD9TVY5cnPNzQtH7
MmpsXeFH7a1Tcg/lI8heX8HcM07oYTcYJPsukcPAWF7iHQAfQYkZDn01Y5FI1SY1faHfmpi1/BFU
wWXPqmYiZu4E0AQMQB8JuTOLyPkhorwKitJPGnzIL8RJlDAhCi6tg3RnDJxQPYida1YCzXL4J5im
qhfByeC9Z8f7xS0n1s++Y9oDaEh1xL7Fd79ixW9gzn2EBATry/Y8iuJMPe+PNGPkGF8BmWlP0CHD
A/o6/DJq2GDhgaIrLdk1J86mGKUAs3Am6o21EbOMdq7VqjKdqqgPiQZ0kLGCqp3n+wwZQBuWvrk7
pv5tTRjx25Wmr4wWbvQ8y8yNDLu5Y2zWp+dFZedcUbPUOwXYupfvuVh5+hVjkPA4lJSwFYbGyDjr
eUEWqOpx9OoVJTQ1J5Tk6G5fe3umIjnWnM7Cb9usfrLk/vENb9x8s4VxtrG3s3+o/yvKHXAPm3L6
u4AGdNQg5giSNKl9CcKf9tC4zxFwrME1HZUu9IWXv/ml5Si7zL2itQ1UvkHhyKq9EWHdn+1D1fYw
YGsKFwN/8tsXbn1H3GXBoxSltFtRFQuk7fd53nuu9cKbpoXXdWbdPkZAhG4wdKnviXdnsnLhv81M
HyP76UJ9dgt5zLLfvpbc9qWVJHoFvzW6MViq6TSfwpmq1aRtWcIeShR5pQT1dAKdGnSGANMw1Wi8
AvTWwmnXqj6noBnrjh6MpOAd/x5VTyBiU9DKighNkwoXtjZUlBlXOWOlwSS9wiu8q5TyX7jkS0OQ
UBbTPKXBcN2zviYqKxtXMZ2lcNZj5jJuvKwvWDT9UOovw5QO1QhsVjXeYrYyi+oqefdboWkoGa1a
5u8UP5/JtYdcmvZdurj4tG3Jpc4N25Q64/qcshWSCFjuzBK85nOgeQInlfrWvIy6i8m0J19hnmOg
EInWnOOH+dl/yEcmbjOHGP3Byl7PZ3s3uFHwHZsnupA87pVPz7+bOWvfG1a66xHWRdy3glodKEfz
on4wunRex5sPCSOOydwRv7EQ1nkRlOqyjS6kR2RKC0dXmnrIOP+jC3LI0/yDLL5RKFFWZnAOxQRM
vN/O7V2kV0NPTS5zSqhaYkAsOlwzmFkLSRfNs2V+UL3jogokI77EatXfwzB8+F9s2hhKw1Qhm598
hzPZTLPdy9aokmkgvgu26TF7OxnlhO90+H5zm0M0cUQ3Ig+8y5ySHZCaeyRpVP4wOfjuFN2uePjh
qoSXzHTLDPz643MncNLabcqDRFTiXePeJZ096Rp31fBXUuybtuE53Qs2TT8LqtfucIjlY4ufi/K7
D3qFpOKViGI/GdAcZuTkg7e71Uyft+ecvMmU8RO11lmlf5PfBAEFwrfJmYVTFK+LdjYmUS5G7F0b
DtKMHBphDZHUWikorTpH82bd1ZOTs6nuTUYoE/UXTRiEHyWQOFNRgUC03MicVq/gNuyZMsGf9XCJ
ibaydh4A0lQOsqKLhCwCR34VDnvF2mb9/vxQ8sUgZEDNa32DfAHvOJTXrWoskUGgKewBBM0jz63n
DpuRVm0SmLGjcR+6F++moHrWz2rxwiSGUzmw+DEmWPMRvzUqHvmM4XW0ZCrtwwlpznfAgc0Dk+C8
akrfPIqz3US51yfOG5AUFdShBokjf7Fp/jCHbozw9+vgCR5EZZMTqaXbSDpF0zyoKac2CqCIYPN3
Te8B7HjHsHnot9fWxwLHcAR0yZFRsUh56jEoEFgepX0omboLcc7FkKJzlcu7eAneRbnH4dMcMPzS
GPKVUw4GNZq+7NPTb7Mb7QCgafgep9IA75fY0SGQn5PbIJRuhA2oCHvlnm+ZXeUw9/c897PBGwAg
HaX6Mdtsf1Hc5iawS5XRxkONdUa1iuImR5Wv3aW3UJjX3iVu87/PG0u5AcX3vzo4IHoZS1hEHUo9
CzyHCCocPBx+3O417POUQoogefmHXDcoX6hYF5kQ1214C6gkFcxjf4vYMfr2L5aDY4XZtzWyGDfq
Oj4sLp9OhUe8OR01dWHMBLWokxbWW028dG0RJKEltod4oukeqO8MQ9jI2tpifuk19///g0Y1t1c+
IfoUXohdal5D859HjE3V8jGFdwgwMdp1iWGPUxfTduC2Zz9kk0S+iJl+RRIkrT+pZXblSIIFKkXM
xlUJA5fiJbkA320hiOjaTGTdDudeoSm4MpacWgWpQNyL5bx7JVPEOZOUP5u93Fy8HoE/EPsxVF8f
Gu2nUU3oDqU3SLesCbjZwXL2oKxUVq7MEI6xJQbZl3GVAn/j0GZEEZQ4dLIOr/paiyK+R0m8A5iC
wLtZDcx9x+JM8Epzckt561OWGEY4DQ1LHU36LouVnwwZcZQnmNCi3kK1pxuruf7rog0qNnhmM1aq
QffqLV9DdlIHaqTnXAMOiluNidwd0KCBsGjOG/cDbCxwjWBvoNy8FJLNm3ZwvH4zlWPkBobNYJSV
7s1qtwTy3+4bJ0sgU4ec5CROSYyZBgdTDNUPMHWfCDl5OocUSA68z6mR5ejoV3qOYDrRRkOCRAVV
yn2z0i/u6QKFuDaL63kX04NSnORvgRa7bX1sZVvV7AIaGrKW0deOlON7IaRueWB0zHAmWqLDBmD1
t4JkHrXpgq9+dbi9NWtq2SK0y/epB/Ac1aAo+V9GbQ5izEUsv9BnWFLHtsdXXsptNDEsGYji0wdm
mkEQtkLwFYyxcqkNjjIQxwHyuqzO66LPO/V6kk/ENJ6fkjUHvf3LcE9Gar5VNdRZJLZjYyLY/xUJ
4bfiFudW9CAronb3s4rZW6jUH7IinKQwS9qCaQ4woIMrbWM9c/Laxa9BH6U3bvrdO5hN4/7Mp4hp
YSsXgidTmM5gAImz3qLf3thy/MWpLlrdi+nOsBJ04flYzxi3tNJx2zlMZBfs5kqBUTtplrjtg2Nf
Af8SK8lPGUgMMa+pOu1spDdecXGlhlmA57jaK2wHvqF1fVRMZy3RX8IwDeCdgh1VfaAUbo4gK3fQ
rU7cFrQ3g+UhE2BPAW9dNTquFvV3N5x2uSL/qPgzk1NwSdjCJXJuU0qlUEKxDMjsiDxBcAJbUavw
+rMEoreWkvfL7v1havBgy26kmZX7NyVnlvS8sQc5fDgge7X8UbvNf42ujrhgsuH/leHMm6dR0GXy
NPHdcOatKz5o5DnlYeWOaDg8DA2qUlpCaXK9Rn5ga2lUrrcuTs7n/HwgQ8e0rGfxOWOPTqZRjn7L
x0NwHN+j/8JAn8LqTD7lo6zeFHHLY7PjjVbPJDYeGWs+O+dLvR0hikKK6l5B8XwzAo0tgfW2KLwA
IvgbVTBOfG5VZf7JmtXPjjcfj+/fKGQQrHJ5su1qMR6pJQdfli1v9+vHoXMQ1ROvuZg58WU1ygkl
XC8pUARhJetF9shaakxiKY79AvtfYg8alX2Vyug9SfzTLfw7grlGMb21eyT2GWpIkZkV52Xmf2MR
sV+UDn0gRXKNJYIo2aomOVxN/ctOLCooEgY3BU+evaUeqqE7MxmntY6PvgWgD906S6c7D7IaC6sh
j0st/P2au12oI6LAS6ZvJVri6shnH1cqdD2de4M5cBBYZ4K0/lxD/EExpwQRr7Sgh97nU2J1DNB8
KLkyOGCOqj4F7NbpSHeDzCQqC1QTiVZsi45hMhBvlWasCuT+Pv7SX9PyP5cOK2SsqacGzoXd+YAV
kipw6bgv0XK+Z0pEPtitrN6IsqWwTxVBx2dT8LDIF4CEv0YZrIfAy8qwCiShp3rhbOIvcnETHYTp
KMFiDkwvzI1pLEssmhyXYek/eBpWEmVetgTo/FgVOjflYzIgTor43WD7NwNJlbrvTcTWczA8QSDo
5q7O/9+ggdxwjinqQEIKaF1AbeX7bKAK3lTEtty/2paFXH7YEv7Vm6Eo564cN4VjYJ+024Vf3JQd
wTUJKEwDCEvN242+AQbigxs1qCgRnkeJ4EUyd9+AAhmYrBYC14aPpdfp0FOUTIqiZ9pGTLHU4zDq
EH38L93TDxWj3z8LtWmx9FMjLoTFLHFpzb9bHv9n1AoxARXOyUjf7X5qZL+RGekXqIyCd21OKkwN
TkPdMi8mL1hKZCW42uSqzWTxn+F3RXOXxSI39ng4+wqL0FtKu2urqGrkm99kEWsiissGFs1enPhH
kwV+Slkip2OCcO5IoRGZVntfosZprUEQ7y9Xn4TOEzvyRUjlEIx2b+EhSprrQoo1G/igB824sxop
/O/AFjjeHPBcUDZHD7nBLo7ZVEmBPHM+Wj6PuPmkRF+9Vw5JqOarV4/xZVD0B0bcdPKZAv0inI5W
Tpizi7Z30+8tcF0VkHqBM7pWVANJ3hfsVlbvsstT//BV0r5zZ2v9K1ltwgyLLoWkZUkGZW9c2/Vf
KYW1ARDqRLCzi7Dr/ZQfkxfv2eYAgK1aLJmGULSOSjmRCoEMN4O+Kac/IfZekXUpQUmyoerdqUt3
JwEaDF7FzWlqcq5ev7DC24LoGleOxko1nFDQzdiFPlIjWjp0qsMJvNmIXWrabdy5TzoKnLrKY4u/
NYfr5vOG1Fr0UBHSUqIJ5KUa75NchDJ8YxgOiUHunWtb241PvBRNtX6YvAeqqj6sOlWS9eE0gtmN
URc9u4dMIRDvxmn2C7Ue2szQ28UWx0NQtp/cbP2MVN751x4h2mNoNTvOdIIrg0nAaonrrDtVEE8x
lDXxsZXCCcSxkqOxHLUkDi49DYAogXTCtPHqumldpOq4MTBxqWzgWWFf1VOPtJScprySODjKVver
KpY1O0EU4BdV+hA9tMEmU52cE0jWUWln1V42VHUtvSrq2tRMyhtjQTyym3AN7xIKYdR9OdGJlD7I
iShfs+tPQlVWR8bf4BjYXkq9hkcM5TTv3WIEIRemdHKC98uBwODXFzXPrp/y1lcOWtJjf9iAd9sP
KGa5C2xA19i3UfzvFNdCv77RByUCC3H2cAkJpQeprHL3RA/zbyuixlhVjHzCUnVdPILwe7DxZOYx
5d+6VswXNrzgGPUDuU45/B/59C3GoTyl6JH74gnOhnvDYwycO9POV3AJlDXMW1sx9BgWf4AO7ISj
3f8OHXEERlANz4J31wZHieBCOfC/CK7yJHiQXs+74btrv9OGFKb5JaSN+vKdQQgPcQKeVtGeEi4o
59P1jOL/TK0XbKMxTlcHWVH26NdUyOOSHo3OrVuoUkRNIziO0/Ocvp010cuF6bayzCNSwPBtOj7S
Odrs+Dw3AkngXlyKy8MThQSj7lL2nD8wvL1ZfBylXYivVddeXU9Spyzz53cxZtmfUA89X8G3Nge5
gE3O8X1o1Zu4fL7R1u6QaM0KNjG6BpxtaGb19LMPImCSvpQzXhyLX3IMSLS+acufCNP+2YpVqpA7
K/BPDWIyTG2vhAnfCXohqruNJPJjBWczsMtX6gJPkD4VOCFbxgaesGBC27LXS9JaUfuFNe4759Vf
B5fEsLA/YkLiN7ILMZQSuC3BbQSLb9shcVJCS7mpuDzWpTm74PJ1dbbJmeFcOJLzsiffBtjdE6y1
fnjr4hZuf/JNdeAxSiLEcbYg4hletYH3kWLBogVRUaBoZ8rHGUXCj5bmmexv7l9Kfjfh2YK9ieng
ajsklH6TYm7ZMq8xnfcqfKuLCyZN6SiA7e80mUBHYV76wSc2PoGw4Ybk2bZbajsJt71pktlx4scU
n2wmIiADy+hCqLJ7RT8tgs/kBxsxRACUVSUhTqpxtl5c4DFF1/dctzTxs32oKtT49YopL42Gyr4c
f98CfCoaUir/odXhewVmHgutSdGMfjL6CfWKPwpm5GjokVj2hhV8xW/CWzQbRRHiKcJDg0M6nr1N
mwCRKp4UKiLNTz5Y2Uw/2tuvtQ3CJ+gD3CirdywIT8zXFz6avFmkfegWU8HXIA0AA9M1XKDxmYvU
p0AzA2ile4d6YL050Cj1+Yc5bw9VIn8sJq93VklbbmSwTIFQEAT1f2f0HXYAZXqu3doYMATgQWLs
blYqTenymRNnhZdacoqJI5Z39OsuqPzU/mgf4h8jcYS5q6qCieWM/gMAy1pFfk5NyXiTamoOIK9u
vH+H4mcFih8VexSWoIrTiehfILRMGp/f+X+E+3asDkF6fcjT6W8w3IiaBoS5oOyoI7W7wa+nqr5T
3nGJkW80XaDEtImmuOltbYoU4/rS7e22yTLaZ2qBt9DhXL+5bB11567PmojtbUVL63D0ZlkTlLvM
gRQjNpjQd0tGjEI8f3EL41xnLpCrWyecqhDkasmWvIS9c8O9ugqUEFUabkuIlTWAkEpPVLXnWld0
ryRnqWOFDSSGy6c2fI0vZ7OafU7CMaCdIqQbc3U0C1/XE7LNZ90NnRkylrp/CzRJWWH/VIAk5wuN
+czHpv9hrYohcxAAvQAzsThguADj+Nqqp5GWvihm2a+wcoPJUoaieDa/j0aFcpSi8+isXQw6h2I6
/dMODNimVJEQhSFeb9MQN729UOpTE/oqN+wzrV94FWHlRzGq1TQpr5/FRV5B8WwMZd7fJryo2SDp
YkO000CCBikC/PyiGzQgCOwbTt9msSK/NTIiMLOZv1KECgiGkTbmMOfhYNalhaFjqLPXpz2FJLO3
+PEZgWBUBcdtUUEnrnhVRd2yFewrCV1CXqIlaxd5hupjJoySMmMboCCJPJJM4tRrQWpTYvj/j1n1
vE5v7dMNukXAYWgBJH6/5SV70RxS+IGNp5wonm9s+rPtb1gKkoO2FNlRST7CtI0iNRI6zqAic6iN
30etTMj7OjdC6/q9chbgu7D2VgYkq5G7jd8XQ2bDjXpiq0R3CPqWjd8fADnIWtoxd4xilDLP8b2D
4x8ZRtxEHQEE8rnKxo6AR++C2GULUSpre+NchMoQSMetNXp0q4qiElNHPV2hBimx4CO55y+zb0JK
mhfHL+urGFSh+tiCfhR2ST9GfnMr/NX5sZIULHfnWr58s98UUPpKhdCIdc8jTP0G9bROhkLQeKYE
g20PsPylp8jERRyKLmZaMJpAgOIZWafv9aovf+Yvf0OWpG//cuKgMqusjOJq9xcSasNNjgnXnWNl
FXhFIuP/RQLl11mkecJsNGHEvcFraN4DgYvSrMRkb7JjTXldCPEJ2b3ecj6Pe3LKuLZZK+IT24HM
Yz1UaxjaOvl+R7lr1x7Kbu1ftmlQTFaTawKBkqy5BwU9QQhtf0/8RrD6V3H0Zlr3SZzqG5mNm/gF
oYj7OaQMlKJq4UM9t9roROM24ogZgEEquq1DLaR7ps5v6i3SQ1wcet3of2Qp4l6Q6+4JqewNotbd
eUyYEfWSHeXcveyQ5Dq8Qn4mFq8jEflY+s/j8nLwYx8W7vGIQ4maC3GfukxGWLyi1G/KddzvmUhl
dkuEjvMsSBVh24vTJNPv9YRZXp/7VlVk/pRUncWg1SnMQ5wuc3LZfuYwWUW6PhqezfmTQeJEungs
zPw59M8xzei+N9yHl0I3bmFuuR8H/9akrUh//f6PAX7acCR1X8Gj7ni2THtee8pgFmU8rb3/nf/E
l2zl9/GSAgr4h1MGUROY5yznZYB+u0yNtVw6XNnkgAuXciBW3N8FC+ijJD08nfUcgm/CAjL/SpPC
wz0VWX84Q+tnHrfkeZ6k+QnZWaVhxqhTr1CRt/xmNYG1APwNqz9MZrLu2VeEQRwBQxePucF4M549
hfS/seM6butlde5Q5EnHVET5jC+kWoxy4J1E7DB5NRBI+qHbfrIAox0HPQEjYOi9zTdUjoTsk/wm
CC2GUNfFqia7x3s1NDBOhb0bhn5EKvYSqGY9Ke4nmuhDb5xXr2gX4iGdQVKP0x3PF1lXO7Pusx4c
Ur1xdoxdzZ++HHiGUNpS47TizdgykYhFKR5iZ30EcCBwNauI3Bi/GZhRz53WllciDn6UDKt5Ks9L
YsrisvQbZjZJ5RxNXNh0SnhnLLIThdux+tPlr5OncGHxygs/43NvYdvUuo2RgfLrMymSIq47oMSo
ea36CvWuZkOGOz69rrtMD/OXd2mJhSaBlWv9mU9wZwCxT/2FRC7mtkFT8zSVfMqQr8wIbZDHiwKz
FQZKOfESRupQYgmHlGMUaskpnezZIPL6FnByGuQirLo5V1PBeRnLLdsniAWS/HBu+DkBJ4voBDqK
u68+6X9GSIglvEVAlOLcf1OopYv8YkblN9Q95kMqB5zPTfzQ9r5c8rdqcb1pe/b6hQx6FDRkUJU/
NEvA4VE8p8UzpfnWqPn0dmgb3jIVjnJx58Xw317NfLNqTUWLtvtrF82QvnJRks98TlhKUldUau6u
HQyvBNybGhGPxgkajYix/awJym+nj9bFVbNVy0uQ3/7qkl2OeQwk+hBql+ASn5ZrlJBqeyTW/cUT
/46jfMcNMtY3lR1M5zNIotSjMhDQcJRGoQNpZnjCZyGKZtnnfCCo+rgCNd+aybmPjhiJmBT5T4IJ
gzU1c30WF7LgmKPLGzaAbTbWBMMSWTCXBB0Who79rS0odh730fH0OWd6ZQg3dXF/QLgh0LGwjjiD
ZcWud0sPZLQN82dJcBHaUnK4QF40VpipxEQrlhi3i8YcocLecCSaV4seeJnPcJZiMJEIp8pdjdsL
IQKQoUVOfmoKXIP9Osl5cq1GbsruZC69xxrLYO7s6CZtkB2DaBCaoIqNIpGQ2OQDTVdyjAhIpxzw
7LJ6LebNIKUOIttyno8dnt59IP9J64DJ84RcF2CcApr1gehuq4HahGWtkb9gWR/ccrEyMAmvwoP2
z1q96zSqJbNALkx34Bd4lhHwEIZl9CEEJ+dSCU5TyLbaFsgXUX5L2oEcW27HHwItsyfjUAcLAdzJ
+wrM3VTHwY/o450VNkWwTvoW/i23JE3VhSKO1BtknP8nZywxHRWe6dI3knEBph4DiP1mYJu+WqqO
Qe0Xxw9Sz0c77ym6wlUy3obOLmltfSgpe99S8ahGl+oiBBF9bCPgC3vNnG1D7cOVwYmcS+fqpSYj
J0T3hecN2zG/+0UeogCcxd5WFSeZZmlkUYVT6ZIDTRfZEjYEGO3oyE4ymJnaoQfmLe04DahlcDJY
miH/HVQARRHoafC3l2gkTnDzWqi6wZOr8lg76gZR+A22qzWO68Beg2ZRlY7yexfRGNHWAYc94AaE
/JpVRv0aplp7O7/OHDa4SBwpxKjLvBuJQTOqXz9N11yLp8RVvDkfUGkLD4aFWO/VZzIphNrF/tQ+
2RU3mRu7HSE7dWh0HWh1i3F5BmnmQvZStiCzBaOCix7q8HmPbx514QOqvCW/1kLg92e6z15y+RxM
Gl4Eyu7RhGxEjDd8J2e6WA4rJqv++gvkIP1QElmj3Jdl2uhKwLpiWc+28U44rGAWyfU+NhoOeY2y
MoQatExQMbKBrBt62AVMUolFNRlyFNj6bkLjinIYmck4Xtpi1HO7Edm5/XUTMmvSBV9mWZZaWO73
VqCUJZzVq/5zMtOhlrBGS8TWukpR+jwortR3slfDXvUgJRfjPSVEhQJIVv8/R2m22mVzbBZcLac3
7flgePLOqlyF1VhM07s0vBTQ5MNiuM2PqUe9eDSi9ZCL1Wiuk5ZuJv5GHMLxll0ksBko1p8hChZR
V/kV9cH/3vU2YBq5gu1XLsbyxocbxrvWn7rKTt3U44S4VowhybaivVOqA60nAmLfTHjaVLKxOd6M
QNBrH8+eTog+aVTII6UNU7ZdefhR1EBVGl9IcTONtQbIcmaDK4Vlzb3zv6H/GYTe/2Fl/AJ/fuAc
uwDhE8z2OQOdazBW/UtAaJLJXmIbrQ5Gm/iZbU4rbscP3tBLCxJCKVA5BW1AVHyj8GlPgCxoOfvq
0AcNpXzRz5KiOZEE849VnqRx9IiYFHOwQn/eYLUJaPem+mfRlO90XxYvURdimxHg93qRybbmI8pF
27zAKjf+GHFqp2ooHRTMb4ofOCWoLFtXUssmzr3P2yT+kHom6UT+zP6psO2gS4yI1Kcz23ayRiAK
oBv/URLDn6iF+kEiFW5IiDwscGX2aayIL4zoGYkpz7YPAN/Oc2BBvQveEkEh9QCIAt4ejXnWAgbf
hYcYZJHvs7i2qHKvbVomZy/O8l7/z0E9LdSXG9U3WJFJonQvrwxqHGcAcX5YdAsjxpsavSa62Ie5
xGxY8kwqPXt1tA7f2dxCcPBH0U8KYYVp3h8K5jmTxlE0oubF/TtIVr1dHV+jFAS1hfk7T2uCyqUX
VZIVDmnGL8Sb8hos+GX62PVjjUplXHm64TAHlyUExwlqV3+5m/154e/kLbltFwMjONghTqj3xtJQ
hfxVZmX1bxnH16GDmKQohQHHaZy+u1EbD3BX6dDRVjKZ3IK1OYmdGUIsOLlP8cJ8LmGZvfvHIf6d
S6u5SiVVRQ857IXtm3/SbfJPPYCgSbFBJfoCmKlANEffVk08Ms4TY1Qxhb22MBR+1PpT+Y8hLPw8
wWH3FbQuozpM3X0M+H2UaP2IW8OinGrWCi6EuCUaRKaDFF4ZWGeL1bfKusfSMJeYi9w/t3lRb2AK
Ukh6VzWT7PP/Or5dwaQAoksYEJjmNgGVhjPGEexVqrWUsAcul4sIcQqixtKvgoeM31u6NXJaR9mO
I/IfEFanpEIpPkE8yC/CWrsKR9ZXkQoYmfHFZz1120fhZzvFn38n1VrErrz+AA9rqN6YuHb85nJ4
HHwxOh76YBOdAZ7y1ekMBc39DDvNMkeB1vgXVNn4Lsryb2ym7PdOwwvZZYaz/sQQvA9sGLfLsl+Z
HPZVHJ8/DtTn/GPHNZVa3zx5YKilJKLTfz0k/xZYKhPDlr9UvP6O2X/KMNY1rv8Nt5mcHdJZSdjy
bseV7pl8UCniCLKiDtqHopNX2Lif1lf+Dmw3YTSGZHfD3OVHmWeKLJy3MDi5G6uCO0YLIwYDANYI
1UCqbKOkyCECsuScJwRCML0EfdWkSkEzXNXe2ExmQxGPpKc6ppJIgwOd0oqna1gLOLY0/nl5pL5n
g5GjXww2cscWiwCFcbOuKD7fY5MCpSv6Uvkk6IwTyU261uRlGKWrkTE5zgX2vZBkXXTUSQGoOGL6
noWBEbuZGP5Q97TbVhUA0ewl6fJ2nbyAxIP3n/IBg4HIuhKGYmE9rs/fdSS7QZhh65YYG6h4Z5Gb
2Eer0sfSZM8/suPcvcQ9y19FXzIC+fn8jtBvIU7GeRaHa2RgMI1xDSLB8dWj5880yD6fUp4tgh8I
UkjMwUjBrfnJaz/sxOEz2wWJMYe+Z+k5cm8/rcdDD8CAW6GM00Jf+64xJntaJaL4WIby8KUAk+rz
3iVoofN1Z8fWIbOghoK+YZ+M91OE9uGVyfr+fEVw7HLF2QYU4lxkmvIWToQaQ/WYp89LQ9bP5xEF
2vF93yEv1eDXww8mnxvQyjX39MgKyVGu2OFqpX1Yg4u8WR2tzP/5g79ZNQr4RKKedPpjCN5TzJ8+
FeHmdKjvbnP+GowoObB5ZQ8OrtzL8bkNSrKbRELfYnwnEuOJMALYE9bM6CgVq4FiSUhQjBhWS558
ylBngKZKXvVnMIBZ2S20c18gHQWPX0RoGxjhnQ6ZP8eT7yPup2yz8umSYnFkCp1jPFT85Yix/88W
v2yPYJs5F1GUTELbb5OorY+FOkJ4p/FnuNNATkoKjZqKw+7FgAPo+4jVKp9c8Fn5+TsVLhG4z1q3
vN8bnQyaBrccA6BWhbD1OkW5vUFo2L3v4xi4O2OmiGf6xhE9zjKGnM5TPhxHxdrcYtmFSC3x6obE
MiQrjgRcodXLKMIZZVMeTJFwbCC3ejVxWYsluK63UhQFmPfVZsl4kOJNK2bdrOODX5TsgnqgNEzf
GJyd1PGK3EneNcuzOa6GbE/ZLhaksLVk1WRN9ib7G3S20uNIibNPHRIv42oRy+t0ZRUBlH2nDBvP
GF050X9RCZtO2Kc2TH+fniEws1mFmDFXiWLeCf/othQ6qMjLGyKWzOeORGDTSCYMP6EMkJFJZDmR
KIa7XUGXwQCqdtr/+3k4R+9vWMB3IkgJgsYGKv6WXyjYoluplzmYISQBtmIaVQy1IF5xtjRwHKEZ
hOzIGmsS0T1VokJAX59Wcf8YxG0ltRD24QUEOqz9I7/R0/uew3sfY/gnFloc/xBON/rF37j4nfTn
x21jPo6gjCaPgUruQNrhwEjYjk5azBq2i95rO8hCAtOkjAkhQVHkEoUtOeiifmGhd0YFPunxUusm
Xm4WzLlb/RMJs6DEq+ivBnv4nRZfQMIcSdWpdQX/JNHHPuMGML4kgY7yOCUtM/rsxMyH17+NLFQN
hJIKL5xhJY1OUTnHSz+QeIwrkhH9MOHwWNO2RF4gsAHJ5JmHd6vL9f5jB1gN8ffZJX6BmQNpl54F
MQJPxrQ53w+jpCGpb+Q1NJVap9XDYH8/aGuRx6axNNcUfQU5Kn1HkVtORKhConn91O6snaKYIPXk
XGH/U7/IvnET/9XkJmTy32ZR1h2JNpwi4KJJFyjv0rdKLH+oTbRvAimaS8amhptt3keyl3PIM/j/
vFIVjpdcFmDGBNDwLv7it1zOS6ng1mcQIctSfWdSmnLpaigVtSCPp2tINSQ4Ey+IMpJWS8rVBFPX
A1q/pofQimPc1w+iIb48QxFayT9OS12DgT5kbFg7+xc/nLUL3R9GDahlyxERkIp4kFekdJK6anCv
j7fQF+lRB0eAMFEpc5DECjkxtI8OMhv2qZ70xFTi4EDPkjzGEeD9Qx40cGgHpnds+PeyeGpfOqEd
gpX5ii0lmyiPHh8KLYIYRqUBN3qQtHW5yFtXzDWvkUGezp46oGnSeHyYS6paqi7bWJv5SewM0P46
Selk9Wgej8ZnOfytJVydW13VIpoQ1425DkuAwu6FI111RG6jOeRt0f8MiXXkaB5FWS+fwQnzQaVu
tc8BSymVlaivDzQvC79Vp9hHTd5PV1DLKTGROfh1zilJNzBts+AeCYxfxwfEM6uwHr+CHm04MHvF
lN1Yx43VeBJFR1fv9rGu5ECJjBeljp9by6onaOFOtwcYUyeAFJL6AF8nnKKovpCOhzpqssZQiDjR
XoxZdGLY7yh7yIQjY8HGq4ly4z2G7pvP7UZMLymgfP33t/zw4dpekKAAfCNUg5gMAik6B1+by8m2
Cgo/Z2Ur1bEJNKDkkZg0RY/ZaCgCXPGs7vHHDAxqhCXeZ4V0nmOGMGzlbYaijZqIuZ0K0JFLSeJH
TS9/BRtnMVgE9Ev8S8gPhlCa1sVLue5Qi/Ba0pISS5aHX7NN9xl+90iNKVQpiHlgkkbD7ZpAaGaX
7VL0MxPw4wD+V21YHmshc96QPmd3nqW52FKIVhl1vNkjlbHQ6fiVdjzMq9tFiUId5Uu3xZIBxt1M
+E+rT1B6paFbAfz0FfMotT/rRxj/FnlvpAdWU/D0lMf9BwNuS9pbrP+6soC5KqOa8a9bZ6yzcDmS
Ki4m/8O8dK4rgDvh4wG4ms71u+lP23a/ZZcANPacc7YOkIZr6HbIjptdMMsl+agtP04is1JzrXQG
8gpjDNgI7c6QEvgdlFgsqhcw2MPr52dmT57U+ajPRMfSSbHvKdi6bkmntx8feh/PXMmJnr3mdJFX
F/05P8sgTWuiasEkNCRDNS8K/Mc7O4Lk/K/1vPsdBbuEjsSo1L4y465rHUujYtO1JreSKPRl9TYH
HhMQ68WDyJMYqJUZ2uu8tEF1n88pap68CquNt9C3DcSEpqJw38AE581VErgSE/IYPeffvINqSGLW
tJgVhORB8o7wOKrJjauihtKRcA9V4nKRHzotmsTVZ0T7PJdZBt4vdBqNL8sUIjM4a2FIPEWV5yoo
OGUdAfC7BC7S9w7NtkJx3LOOo+7XnnO7o0MPSeO5SUPxiVWT0kuTfGAdD7LYdSZfdt/UxXRt9U1j
jxKzQODMp9Y3Cs3A6OP+KjSvT9ErAnEwOJM0QcxCdL+VaNPA+Txgnu/iCMqiRc9z/WyAkdcSWb9Q
0d+HKdogChdKIFFbpYPiz71l5lWQalcFyEBbiUuNEmnt069OXsnVio/2wg/2n2iN534c1TheVxMm
Iwm3SXbmDlozJHL0tFgESEHHwpzCrb6UKbBYBSLkpf/RIaUEZ6cpEC3nKw7+DuOF5mptiPxCS+wx
Jp4L98irJumfw2k97ES5G3ERajfFfFwOwtIQTgrzeV1CRxyMajFPVuf7BiFdnaZtA2l41k8SwNCx
q4RiGVauHyfc8gVil1SI9A2oT9G+Fb4qcQ5GzkfapWER+S8Hm6MyyXaG3ZGeHzA2WRzJMnJtzgOa
qQHDLkARK/7GVMHELURXcJuvH525qQhDKaNbepbzUCYkv5u6XHOIIa6eGQnSqnJJdFhQTMTWIy9v
7lJrm0Nqb/0IxKzvxZ7Ct3aVfGBP+YgdObO1fHdl3g8idyPu+4NV3xhpFcUIea0TWFaRg0sbFfec
yFQ5tbDY+4oC8Tcqr4mRB96JnPhI4Q2NmuSKM6UyccfAnuZcQaLRntoNg/ekng3nCbEbBq1mqqOp
xC1QHIfW8feP8Z14iOgCIzMBZiWxUo8S2X215QLcA2YDCtyGn7ub9M7xUCWxAtynPqps0FTPVG+S
YiJNefK6a76tA3Jf5CPxBkjdWAXQQF+ReP3gtVQ79cNxOomi+5UcZLJZz7P1c6p+DuA9VkNgiB9t
mLHJbmf8QrT6AAywl9LbXtuDs+9wT3EvGhEGEYhPSQkhP6lVqTey+dvcuJCAO8mfq+PmOevYFIcD
zr1f5LTf3Pg5fD03HQqiriOgKQS0mly2YR7QxNReiIeO3sHoGXdaBeXaLm06V/qwP1/+6sT2B2fe
rJrSv/vdo7nJB0azGBKX3Z/GMKtcLbF04YWHpZ/qTE8OBCIbN3sutL4v8nAfXBtczvJfQGA1wQHh
LzADnSKVzvOa28FSraZv5nHZDTwEjonxATrbnsa4+If/vhq0l0UpGdhI/7paHrpBs8k22/goUSeo
Oes1FCzdsR83ErAWBU40uHUo+0kptuPyzxBvpeiDedI43SsFpAaoyoadZT3IjzslkrlA4CfjVqYx
180RrP58kYFisQEYo3SuwUgfDU470uSmPn59HlPTCpHtaHia+3nmpAsBJg+Bx3maAstkuvz+Be4k
Wbqyoz0AuZDyS4i9ZT6ukP+KX7PLidizsF/Z4VG8PM0kVj0XpHuEZ0jy3+wJWysT27UpBTQu6cJf
vvSIut9dKoKfOnRGiE73MhT8dfa+0GJG1Nw3UwZKUO5grlWmhlOl5hpOH72uLipGmmoxWYLaw6/C
m9lMWOfgnZJ7VB3TO38R+gnX4xilXgw0M0Sxnz1JHzm8kJv+UJAFORjEk4ZXBZKqPgShgyqQbWd9
NPcepTUTtWK45AuHs8jYldpzL9qOOwe7IMGiHPPDI4AVnDqC1qA5G83niQrENaWeokQWTo6FBXpT
b797L47Y4es3Br/T7QJNsZIDtqAqZyvbagnBvcE1ty8u6W0jPhEFpov9bbdRdMjnYEm1ytn3+Jnc
CN1EOvzsf3lfQAdjd4d6uSK7quQIxQD7UNh2jyXVKcPyUYd88ipVrwaF6kdwM3mpRG/uWgp27IwK
V6ZIcLk+weKQRwmagCb0kLBybxoeyWbBw76HyqoyflE+51jHGHNR+u2uhoKSMS4bJ2p6fY2KRFsk
gvVn2mb1FHpJsGfq2A5YX8gg++zQpCN9S8A+R2Hc8rgPePQiVymSl/7dDdn+91C3bN8TO6bR9ae2
9jfTgcbYpr1gpNPhNSYjcCrAqTLrV6L/mrPb8tPlZCcFR3wT/wyWSUPIR4M/NTTPwWGpFiUBU2wX
DrGfYXjupxW+7Fiyjtvch52sKy/a+VBYQzv+crOfMjN5MBCpdcfRS0EQD9++MWKLeJY2rRnXVjT7
t762kfkuesVxB+h/etZDWJvQl30o6xBSwzxKp8UFe1CT3nUgIf4rtOcaDdIbE2Nkz2LD8BGUBAlk
ROqCizd2ysTgz1bPuOCUG+coRfhWIqAfWA9Zv5m7uxHyEHNnWXQdmcb6hfkmntcDYZZ/LEh21dCv
2izHy88+nkUNNKDbNR6n0CxZjJHecIo+jlFpm/VN81S9JK4fvO/hVyrTIvaZqt8Oe5Apqv80ERYC
0ErJ7Hm28hpUe3mvkiaFIVOT7dTx5kDKk+FNQ6mX9w0uUNNYCE2u4ynxBytsahcQT0HmcEDsnlIH
X0PwONtWwVJ3zSFJO81sOKdjL7FEySQR4Dc1uUCOJcMqdR8eDBtLxpHE25slJx7dzJ7wu/mlvV2f
3Z2W92rwmUjYjL5IqQBw8mLgPZkkKHoAHh6Z9XnNhmRxh70hLXHJzjGGkaZJJRwtR8+YLRKTUsFx
ceXzFkqj6hm1cURYzv4NGL/jh6bHtYOAkho93wxx3ZnZlkKXtgepJMRDL4wm+/6ps/+lP5vzRLAx
xaTSNEbub18tdVVwFN3RSmEjuX5fhJvWmnxMN4XuH5DMEy1S9aoPWQbGnyO8ZCJn2vbGQ4j5NeO0
pPZaoDe1nCnRBUlSJVPMXKlboAbhJSc7QNTpFR4WfncQMINJlsQSgIKqtJ5entZFcPshShjUhxxv
YBaAohiL5lvZPsvb9BIBaEqwOh1IyoAx3HFhztKT6wb+mQaEnNy5hHhcF7rB4paLs9YDNWRjIh+t
KZ5fzP07sGpxKnA8CtAwnfEhR9moVxdinMNdShP5yR0J1YwPJFM5JZSjo68KWD1l9y1p7Nm6OwOp
pHgCjGEHtONCF3AmO/9hxTFnlmZrHCAW8iN2cWSB17O9yI1dh60JGmG9AgSEJIOt9AlmnZHXwjXn
rPClswbi47qAXGu8IWHMexTsBTZsifexp4VSP7Z+EEfVBuEDdbheZ9byWdqeZhQw9zST+pSRCAM/
/aemsSjahXh5ROBPto/wrDdOAMdFPq4ZUOx3YUq1CYr5k9FTaYYgONjx5yHGl6ccWyRoBXV6+Iqy
uNTdoHgAlbJzol5OG8wEiExnZAJb/4nK2q2FzpjJeKZqJfWwk7x26A0xHZdkWWxKWTcZQ8UPQrOO
1ZbqPnPHNaRh+xDZ/4jwQZ22aNgFJKhzyuNj037677ttusinachlnDzctnjmx8rYPBXeqUIkCzdP
1TzW4SmWkTq5RU9Zv0tBAYliqjMYUVXSy4/upwIaCXi4YqfcInzzFtbadcS/LbLqzPyfxXxwAk9P
izPVbCd3aPYdbEIf3aj9DJ2+hwlHkuvod/rrreL2N4FJ1ugJx3cykI921/5593vMSP+Bk1r55UIC
VAUOGQUB4IIAGAr7fNHm+8MU8vGHGN1KtuMjwVORmso7MiB2glM+Vz0AWGafznedvuam3kVR6xJx
UHni0qpy6pMVmGFZomIfg3rJmVmCbeHWnYDu8h1JalTmsZEIclKHBa8RTQNzimvM4ujuCwB0GoFv
OHciF9ugj4G4OlbDp5CNcGL+VbwboZUvOV3MJCMzra3oJyCpoRa8Ff/9hbdYBrVXUWSKSvAvat5I
68lasTHrfSXIYtuP2stw6VjSbReau0Uy43IEcOaTRlp0v8bFFNFO11tdiCNjhpNCjZb+ZBuq8c9w
kYeCiuj4SB34yU7iirA2uw2rrfmgEhbBawVqdJy1yYkXq74H1SIXvHBDbIYV8s/u+uFra+5l37EE
LHVfWQCHSHk4U9Z3r6X8qparBZEF6P2NF2IxCrtTJzbM0pWWjqRMui278boeBh0n+ejMHyhmJ20/
N2iGh9DSE+KAgP01y5Avln4EsCRLEY9gmo5db8w2tUmnjHplry7wxu4TCh1sH1/QTWHjDDxqK9Vt
zocVkpLNW+vnMuJYYjIxEUth4hUytBtE9LVRLc2ctQzyF320xoBfTfnUOF+tmP2L5mucBnZccWMS
CCRyo01q/Dq3i5FVuJ8s490T1jyaBlqTvUajnjutWYvg2ASbRRFFfR0GhdmnIMBr4hKqxV7QbGxn
7HeYsdOQPB3zW0zEXCLPHRY4x4mM8HxCQtMs+2KN8bk6SAweU/0z2uwTv9nsK6foog45jyODugGl
exRKEFQb7edlkFvubXYZc+VK3NGZBuwUF2FtTQAwRn+e1LmIXF0ApjxJBhzuZjY1twyJ9qGskPw1
0geT0eorGWkfuI79WQ+QXC5iw7FyHoU+ZpglztykJr3yefvIFpXkhQtTaUGDnS+MUJXpZGWZT82J
NDT2+WEy2sRCGuP14h8tyt11A06nRxEjm27fkeqRJgmYSHilTA9kGAVMv25KVExccdf2rdl9eTXb
TaRTC0D8zI+ijxwEKPW1EQl9JD13diDSYnIeyCfxFB8vg2wvzYGbkazlB4212Lwrh2XiZ4Pnnyv8
yI6/s9rQLkEtt6VP7pj9PBh1T/+qfq6jPyiEo4J997Y/cifk76DdDII24hmcMEKzpDuiiyFEQuBj
SgaUWmfWCOK/93WDt0DffPWxsw4OTLiI5MBrydl2AVhPVPfia/5ZOfdnz3zw8FKbDkNtw94hwBDs
7CPgUMZTxuH3i/s7/tAXYd0lZU3oUA57SSTbkX0XZrBj2opzBIDPiqbC5nnk6xwWUJ+uQgcnHVUI
wEsl7kl6grfVQKDVRxJLPMGV14n3jvgEqQu0+yqcC5KP+YMy8FbpdKk9R7uYc7N8hyzOBthZn/3P
r1G4B1B+XH7q3YemkLWv5C99PIA/RvUjy66NpWyJJNocXfLPJO/FGMzHfGKHrnmOTtcIkzJtQhIN
dNXpNgfgIM++yU8dC1AJN27ZrdLA+dYVsjEqGnLwotAYz5y2J7bzJjUok1A4uDFdcCmDLDaAQ0ip
r5t+6aZffFkYb/GaK5oARG12sUfz70L/rDiHRG4vXKqeNyM/n0N+RGv2+dcOAv9xd5ZWQW6Cp7NX
eebob4aaOrIWPEPUcu2slSYmZckxlFwObQCSkFh3aw9YQgoI7qk2wxVx6TFMwAj+6nqZ26mosMdw
uPl2TqjFBfvTps6fMlpmfuePkQ7fyAhIzCtONafW1PG46IshQcLJ/j48GyLEFYvKabaC4z8jpUnt
L4D9fR/xs5HqiT6+8ThejCGrE3bywIUcYFasFYKU15RU9rvxiZIP0C8U7mU1m4aiEhs7VVtKbYAn
QKXwxYjri/ogkxwHQSMzts6vQAh+gCmponikeq2ndnWtuOIsJEw6WZEDZPLxcn8fskUhAuCN1U9r
YQry0vhKUKWBtyhp+tfNMfbuAiIDTNUndB1h2X7pEPW7Suk/cvNPZMyJB2t4pZ9+c2kG4XgHXrQ/
FbIQnVjN6u09B9XahADJgZ6VrHOhLn8SZHifyrqbzUkKfcu4XGPl8BYSoP4aRNF84wOvG5Fwi2la
Dfvm35cxOoycxDCwEE5eW8V4Z6RnpTXP9Fl0+3nwnGLPPlV9L/EOIOfWu8UuFsXd9HqxAH88BGeH
NnBuGvk4pVSdd+b81DSKWs1Z5jHjx/ErBGFZSQKAm3Ku+EzFWcEH2wWqUodslhk/W1UcDmmKzdIJ
A7EGxQYJIQ8aq0beBvRQwSpVJ1naoEOS6UbwqC7Ohi1JFmF5s03z7CBUKGjV0KHNzOAKXGCKP1i5
4bfSwgo2+QtoZo3L2HQYfAVCt+QHHiIacGnlJvcpP5mRmCFs1syfQw9w+ULwn99viirBmcwtKPPP
ift7NDXlAJwzXnrzIOWoO+9QViRBldyJXifPahxEU2KOgduFv/0QRJqIWyX9RHe77jwBsPgCRU7D
Vrly4l+PlpilyIj2v1qDeIX+3yxTtrKMuKUeaGFbDvDMu+U+wXda4SyLZsAHMmde1RqYIwCQ/zmh
MqteYmO9PNn7vdSMQHEq42zn7Lk+qLYR63OvB1LZoaDechEUy6BMt2/a/EqRq8mBNNMnHFQDpAUU
DM4SakEgm7Wz2ZOOfBUONER2DaC9UtxPwioVqk9Ghxoc6IhmTaVByk4wTZJtY0hPAbFqNeCSJlFz
BxMpUZVhmYsLAUwVz6N1lbab9sNiHpICQgYC0Hwk1quPiBkMx6R2rqlc4G2POCi5GXE80CceWSdc
aBlnNG27D3d9gvU+k5WTOti6j3zDTlC73/xua6WxH5gseFuRkQxYha2Ozq0kgpDvrDQL6UjU/4a1
LywDAQQtgI6focCWOAOsNC/2N4Odn8s6HmntQSo7Oe/SWVTMGXq08ZGFk/jQ4I+zoEhWRU+/zFIk
1GHP4DcXN80QUkzEqvNLZqzAIpUT5B2rCR/86rlVHgaUpuKaH/iIYW9CeSW+X0T3fUyNWv5e12zE
ZbFNsuRvjXhCEduX7Q1oxc7gPuems+W7g5FvGixpblAbCM1RLxUq6mg6P0YO6DwD8Ss9JvKO0EgM
4OCRi/oKvN3UruR/KkgfEOlVu2S5yokBUVZY1HsJmWBvGqLMRKOqZu8Lsx7Q8VkLB9/RuU0UJVKg
VlV2FSGCSnuKbbZ4+g8K5nkH9umGt4Ohn/wXBR5rQ7UT6Pk9zwrHXXrpst/PQXBX5uglsHgs8oS/
++Hpiyq/TMDkbfTSEaZNIEYph60qZX0R5m6zjobFy9jmFF0omkVMLWbZE6vODV13dmMbuARHIVe0
ZwPaZ2KFKXmfjDYD18AaEl01yIS0EONs1i4D5SRY9Z5Dqu7ky+ArGwnVSi5Tfjou1PwzgCuDrCLI
0XTLOFIy7jqljNFpGxPGYGGmf89GCFncQPnb7bA11b+a45WnUJtJhpTMiTbXt8ax+cckXTM+ON3r
hgQU8SBYr9ICD3d43gn12fALY7O6hnBIHMh0khlFHFvpbTWkWMrTiYhe7cmPA7T+Et8LtzcAvUyC
xa5kJlAhfpC7p6/2iNbBsTnCtwYkkqqCizKMt9piztR3WLXlP0VSyw4sun2lfyXqZskYCTSi3Vot
GUs2OyuFKHIUYqLp7enzf7UnN2/fhE2bxamkSXazR+h+ietKUcd3xdCV9lIRkovePIN8ipi1RdYo
RP8kMV46KkIuoInYG2WKuXdDB/jvXOvcPxql2ItywfVtrYs4IlSMUdlqewdZ6BjMr6Hi77Hsd8nD
0YsTA4UaMNDuyQKXMKu8u6CaxiDHDsjKdLGaS9fJXnBy+Gl8WmeUPC+bVR6sF3hkJGROAvtH7Ecr
Bv4QDBijnkR/EpcbRBx9U1bHWr5TQ/RorrBZNoCWcapaLJPSri1TcIV7sG3wrxRm6gVrusOV1UdW
j+FROpYZUOgiQb/7qDcSK/qCW7njRIGYrBDbdhazpDPx/i5Rlm6/e6ytrwbU1VfxwagWumceLBlq
1/ovF0ffiyr3KITu2LiRiF83pkytXnKpdSVhXVbB/F9O7nmgkZ3a3/ebGf3ILELtREZYWxLq9frV
mlqFz6J1PqpTy80OTOKm2Ls2cIs7zM1mC7VF0s9scWGjbuva2VE8cSjHlMQExzvgGyCFubG17179
BqIThneJhHiGF2vBFBlL4cN1ctwmMuIr0toHBTDzoLUlE2qGkljSTccbEwyqXsNeS4kIxHh9AQ24
FxsfJK8HSmA71F+Kxiz8y602dUVSRXCJ+4JaYv5wRUYg6OcSIo/JSYFrl08VRC6q6i9P/HF7ylt+
SNYSu44zPLLBnF3hZRXXIlg+vcehnxBoPct+uY21W700H/6DtTfK33HMoaiWPA92tXRnh6daC/YM
iksCTIWf/GbefHCtUwBJtj2TuMdZQ98W+UxoPU0yp5QLCucejHT2nMu0DrOxMvxtaxjwo9bW8Qs3
ACjypgnj86SElAGUL4C33XrCP2/Rokt5SJdtEVWto6x3DhV0pivUXZ00szR1en4X+vqCs1a4HxFk
r1QNPkNROuznPPjwINdG4eelCFroQEyFTh7Bnzk5s5DBlM98XH7z5Kl1K6AwaenB3/vKsmDfyyn1
iKyNPwLeHgc1N0qc9ijHgk2lqSddGZ+ou5Ng9ddVEy6cbIiPzIfzWMrrnBwgWfes2QuU6NDYJ2Vs
LcXTDblUuGE0qIR4GMrybfei4Vp3+SuXCHQ1Yw8FSfSWRNZdvWYXPlFEK7LxkE7BZucONZtZaLsh
0uXYqt7YJscV7K1aTWamEwZs2Pj80fxQcQy7iyE/timYALF2lmIMRkZ9aQsUWQ2dv8KYRpffNntn
t4V+17Yxx4ob5PpdaeSYjCI3jhOahAbbgNc+BK75535iKXAcJCS9qJX8eqRLq5+Y4iH7yNxLZQkR
NscEuOmbdCTu8UxalZLAOVM/fY9YQiYwLdvi2kH7Ee77bAcaSotkNWpnpf1mO/NFLawHmDxmhjbL
x/WIhV3CX1dVQPk3unVqs6jsJGJAXjSqPQe67BepWlkAzvNQcyKPPZyF4ok1EOI8Es3fOXTfR5cf
R4BDp+VYF3qMlj8X05ewTCflSJgTUYA5uZttOyTS98M2A5NFPOVs0jzzhg/tAIAPsmx68UKOjXMW
aDwd54rhKzO7/bV9TgA5MCvBteente9E3ZOnvtS7orNLWx2tgMaJ9epPIhrRUgYBj+2+dFWwZcIH
QNs/Biv1G7Ryga0t+H3yEgQg7sjUpSiZvzvjKuvxmUUW4o8YA4M8TcZE3mGRxCA/ZXRJBHqMBXEJ
f83NGtSeGoO2Qn5ZMBxVNcfBQ3y331xWQotZP8ViXHr9weiXN6reEAZReomQ2msOgecAMKslnK8c
++Um8+2lD6fzJ6lcAiNmkK7XaVRMEuKM4601DgX/yYHlf29SeNMJJi6CTL0LbNBrn4vjUgfpWtM+
6ZS8m7l9YyC5vEb+dx8VJxWhWTmxW7Y17bZh8TFXQDYjkBa3VKgVc5gv1fMjveMRL5X0YPf4P46a
XENgBvx3GGz7vkQcQLw1usafaj0yzx6FJ3nvWCZ0HRS0mbNwg+gP95qw/JG3hE8U/bVjuN9SDS+V
yXx4hSwkWd3fONHJ7+Pv+QLcc6BEyuIOQ6BELJ0IOGugTYjEthn28inDfHtzm9sRdRYZlJFyxL/4
faICyt2cgxJdIbitaA+rtaIkh/WhS2eWorYMHtUaFltQLbn73QuVxdhYtnZT3OsQckyI6vVkJ4+x
8JIoeC83dDM9faiOw/ZaFVCo9xFGBQIoOZdvwrZt+Ap9PBrWTEwA9MY2xVjNI5XKy7ADCAOMJTdb
etd1UB3gYHikEXBeKGXv1sJ6mLjdJkeFkzGge06yZnSJYCksfCQbbZlvovTYMsqUl9xYYuVLTKCo
8OaB17A6J5KibdsB40jln4A0HBQZjjE7BDTkAzhvFkJ9tL9ZSBi3ex+EArcp5qm0L4EZ6wcMdSHw
XqRYzEx2LA4dNngio/bQftJnEcbLh2vzKA16CfcFppapCH5I/UwX866F86ed8in0kijBn0XFyn5c
2ALj0AWWQREAGPD6qX70IXRcK4OQu8q5poSjNKI12IAX0ppchhTkdX4p43AT48PVqMGbzRnHq/qA
dq7zmI/SCzb+zBdQACUhAZFHaWnJeqxf5bPNed7qp5aCy57xbImR5Pc0jJED00L2BJJU+f20Thrm
1Bpqwy+v3U5VzS/PUjpgJFypV87rY1V/XgmBeQddDx6RHBgn4D0d13WpAMQHqsG0chUdYGyc450y
Wf+CXTbQNOUslOl8FOqhH6bo2rWMQXZo7mqMCA2c951/2x4osqWzfEq3FWh3mqMukFfzbEDzrWAh
zM05G0nz1H7d8s+90sHDunJPCyYKWJoP6jyW1npolBTbFHVydk1er21+/XCet5Q1Sn20V+ZUbGaR
Hbp70BYyUa7EWDxgjNt1gYvIClzIPGkcQD3PcVB8LHaLQrU93zyr3eRyxjWu0t53UOEzVd2QjaKm
uV5AkXSuLd+tyNZXEkb3evo2ZNQslW7JvxHcxOt3CVhIvJNMReAMyznjiUlatUHzKbmtn6hIblvo
oA9dJ41RimwpM17hxvPuzP/t/Pqwfqp4zuonr1LlPT6XiA5Zln8njQB16LgpwhyxgSp2quQ52Rvv
0V/jmvYBFhObuygr8gf9ancUXedLWKzq+WlGtu+KJt6LQUH1WZdnR2gZ5UG3s+DjEahpUet+oYPe
6K35EkvJHjk4eA+RUGFnc1AkziCv+mkCCDBIg28gQKyxs629v+dZ1X4q7WagE80eUZJ5+DSs87n6
5Pxesvd7rQX9mOyWzZuwNa5h570QuFeCfYBFaDqQFt6X8O69gZpVnOwXldcIis/7lPomhHoYpMA7
dl8jmUW+9Bzfv0i7xinEvbcaNsduhRyNx+0kp0ftxr598TvkU4qc52Iv6HEQvOsXXwbYA/eurA6Q
QR6XlKEZR+AfI+Ia/66zfXncJig/I+SxakDcXcnozhOxAe2CPvM93nb9UIbIbkbivsLOGNG6LUfa
Wk9ZmgrftDfQQiLUg+sgshXMjuqhx32MU4FCpMrFQh5otue/EwVE6JXoiiEbN4ndhFXqOQkTuTzg
KyQYlCbSpUZZ9expd0C09iNVUQo90W+dNEscakPCj6WLtcD9KuynhAXVbo8CDX8WSAtt2xR04GZl
8StIS03FP8NOt6+3D1gd/DIhE9XxnRJnP2ADnuIqDSuEXkplXKynlCieHOA55dySUc2x+UyYF6Mp
L13icd7VPYyhqefpUiqB4jRdYSXBU05vqYbjnQitC+xkOYNQ1EYOABufmncRaHkqSGQDbELBF/6l
dBAHnrmKxyUD/95Bpo8BEsfYAvrLZf92EleMT/5wprkS2Dto3wLRzPFQxVj30/moM7DT9Wpg2iyR
rTyThP1ZfxQ3rvdKtf1ftZgMx08Kiehu6RKPKMgzN7ntn+M95Eh9xI4Fl5ClJaoqPCvnIdnEo7CA
pMPAdXjoJQ1NH+MyBMxuZ7LhRq9zj6Ghv4Bgu3Ppnq51sj4FY+n38ExGr7nATOV1mIqP6XtRzyd8
QxOQHMDYi44wlwXaqxBeaR6uRfrLLQz7zCpeIjsS+cH9twFyPdLXithds5QRYbarZ6chtgSUtLbR
+9fhG98/tXAGcn2LHiPBj34FER+YzHcjA99IcaQMAqv+74PA22/+sJhGzlZ5rD57dYArApyIc/+y
9ZF1czz6Ab0bZIEHKFPyImOGsytWgNij7SuSzHYaEd5GKCnRctgomtqcuNVtMZHerB9uTJ0jhFXB
v5M3YJDwOQAPPziqMdSNYUK+P0dRPUFqjoyZLS0lijjSml1qE3WmjMymlO3seoWjcdCTxcgUr9Ui
/654bIVBZCPCfDE6rcfKTWaDW9W+Y5d3BNinCByXpZquxSlSoVBFOYsXdfNvnaDpxNUEDN0LotxJ
Cq806Pi1pQ3YVVytXVk4bixXFgO2Bi3j4Uitkl8h1wClo0XoiZjhPPH7PG6whazUM+Drxdxd5JNo
CZiIT/aDXUOPC6hVGqXM4EmYs+4MXLaLq2itm4ryZsKKaa3ZA6FQ9Qmbqm/hq2EnuXK2+L5wsJhh
18NaoGv0k00rnyn0vUIcRwTXqzZPVt2AxxbGV+X3e9IGDQrYAZE9A+F2j7twe9JdZtqYbx8/xiYK
vKONW1T70fHgeywjghFN5ktVl6IgWyOqmmEIB4KfogM65O/Cnv4jgh8MV2xIFQff/mqgYcHkGx5w
b6PET+nPD0MRAsgQr0EEHuwxalAWslsdhF1Lafp1V64+HSQJ1a/9ji9C53vyeRRagZ/iSnIPisML
XaWjxNGvz9EL6KmUluUP7JD/e3VZOkocPOLyPIlWMJaNuFUmvZGB8fXMhKtjvTyT8dASixD9R70q
xzF/8GHlcFIUNAGWKY8sMCv/Hi0F3WPmHKrB9n/wklkR+LoBSXmm9NavdC2x7CQEbEzwSkUS4Olb
lxEQBeFbjsh0Vnvv84s5YVwOlmnoH3Eb/bX0wndJUth8bqj/pKkaS6MCMfbPgtWYnv+436S9Dlod
f36csSAaxbZgUQ+fytaqsNwQvZMm+pM7LQBfO5h5eJQ8lVdegn6Se35HrJAqYOOB3uS3CvlTJntz
hg7k3Qv1gGPupbIFbGdpe2aEJlEVvZ4sEGZzlw4Cz2owuiS/wgSuWMl83xyPgu9DjiKWXyR1BIjX
2Wak5yI02DHZ4HQzvRvhZhlY/KgNP/67oaz6EZ3T8Cl6tg2jb1gRryHP4KFKe0uBLifBwjxCk0+r
x53ne63u+4UAt302a3OVHddw3gNCHPs2CQKulNIfPihvrVry0svYLiQMtZSe7PXmFHm6Bfp0WP21
bRdkZIy2VxcnF/NUgMPM4lHxXBTKEIDz/Ii1TCrp3edPpZ1gHVo9zs8EnLPE7679E2mpLf9UPx8h
iS5b1gEnbGHeU5h4OVcehxbW7fATSfBXrmZKLz5YYTeQg0NP8ZTmBhfTHq8AYZa4r0Hk0vTelOaO
rCXUpZg0OLXC7zhr+JKDH2geB/zTT3mO3B/GIimroaUo95BHG6nOVifrxCycNHLjvbWNBgmaUIqe
MflKw8HWHE9ydg3e1WcZAJ2aTAMroMc/YBOHQ+i2cl1tMiZ+Llcu2DNsZN0kxRtH6matESLiDSvb
uIOl0tk0+xszWg7NntsCqYumsbnVG4xCENDaVwytqbjDe5dR1wyHDN/qwIr2mY+V1ZPgLeX5D0V1
/I7OgEsYY0N/csFRiKvPEccSUdcWOvQn7yh179BLNTwH6E6JDobdB9coCZeBIbLKh0Y9jGgw1/Pz
Mnd0Y0S7xXOuZdoXSCk6Nt5O7l5ER/HsHqqbiNs43u2d8+dWvbeoBglfrGmUxQv3MGKqiOCLNuZs
fvV1CXZRKbcsbvdm0xDpWgkrwKU9nH/7uLs0wiDNxA9EGFwgs2D7taL/GfBLMqv3RSmMcYl1rVbl
38i8x4jKJH0mIM22bf3KPjCfF+XRIilwX0+AnwLBtaVNObn5IbRfpPCbcduG8QUUz+9PGMaHBJSY
yfPbftslOdYWJDA1c0ujHm533A75xkLu4M91YbAKtieYd5bD6y3BEbXbrMwFcRmdX6+ZLLXrx3yi
HZYOqbVGZxF4gy6DXwiMdzFlAUB1GtVioXEghycqNaPBiuKLRcJTfqMtOwGt95PqxarYXlClOLc/
7PDFTrwkX2o/LJzet0Z/FV7XjdWwJ3Ni9ituPxhpqcNRkVsv/iMlPPK+GvG2sHzOoxyRkvmOGhh2
aCwjS4kzg3ON1StLePvWFKYYZ8lL0rMYIywr9BodJrzHzkplk0PQiV/NISK7/soNRQ0mrz8sWgIQ
6ptxmHIsEw/V2blpcK5HW+O+tFAFk2vVuRqPmX8hGnp812xZNlrHVyosKZAkG7CylySDcYs99lzS
tsshoSm6zoOTQVddlUedN+k/ncmRVA6feBfxkimL+IHqu9bQ+7dGdZ2DpBPF8i4Xtq+pJPVac/c2
ArmUPbS0xPRJLaaJK7Prxm40SfUWyKEWy/CbZ8VputcO9y02Ah+2D5fAmk1rLoejUqeLYYel9Zgt
sdv/0XaWLd0DeY2N9KzMWUqmh9t67cFuFKcDMi03fOzTgN21YoS6idq+W6m0P48WJuir5qyDpVDa
WsEPR5xHgmZsvpoz1hiRTib7kt5jgJN9AOcp39wKORHtqB0e62n8VQbHFkc8Ubn0gTMr89LUf2Q1
wOtlAC3Eeo9+pu+DeU6iqx43gkVUOSYtupFjcQv1vJjitWY5s3cjwryOORODhpI8HLrWhdgYmD8o
pNy3FVE6PGy06ZJGDvdTnT8PH0ho8gE//SbWCGNfQdpkQYTl3iIYra5OEw34OIcjIQ6LlyYTW8uk
fgKFObr9rfXkkQi/zqXvgrcTbLbqvoCYjOrfIIOLgGbQ389fNkIGMPdac91g1th/tTxmVCTJHCJe
8IMVSJthBf3G8jiST83iPlWY4hCZE79RtuEdre/whOCjx3/2KKAtDLSbZNwJcjECuOxRTdXWrNXS
pbyFDg6tWm8K7i8U2878AIYjLmPMjVUCA71LD+uxEZQPlxXXaukE+FAD99xYqJGUfx04vaPiqgxf
mvvB7WmAMjQeVW/+25IvV64mDdo1Yoc9f1/OYXFaaLa8NuI06ktDd/1TSMoP/O1Wmkxx+fE9CCjK
lpZEXh7Rf6U184WEbXMeqcEq9qRQUAp6u0wlkgJOA3PK3fe0wBNjJlVaWIirrrpo7u+pA4j2kGou
8XaujjJW+X3Y5MoO4HaE1onzxQvAZwKb6hff/PY7bZYehc7J1LvNjrTSAo3obVEY/tRcQWrEK5u1
hg47T0WxYZIbRdWn5OYMMfhplz9a486fe119hnzn5PUb9MuiBtneInhb9mWQAJe/f3z3PjWRuZhF
AGI4dkhJW8hrZ6t2BW0oM4NOPuuH3zClAyuYEVKQ4ndwifQPxxaRUA8PYkyLShH2E73bGmBaAIbi
QgsxkVEPZt6nVkOC7zMl1JhqsQydTYWoaApSG1LGhYK1Vs/5iH+f6Y6TYXVfS79ojPVfKPwY137H
P9JGwfMR7JciA3A0QrGanKSUQGHqYiGkgwQIGJlyb69mUbo8Ks+1v5lG5VH/GuBGGd+oJyXMy7Mn
XdTRwtMYPyaQLM30LSSeqPml0OFSt5aWtCaSM0uzo34BkAefwsfzbhUy5J3TlMDdSQ8NoGaNkuq/
A7Kj4QiLIl8ieGvv1P1Hlyv5QqRoyOIqjfYl3VO5aXJsn0HxcAi6ny5claVA6SY4P2Np2o+g6+mI
RFzvi6tTQxGLgxhN9DdxJ2Ad7hUWMZl3xiRRsuYenRt4Z/y+8Fkh6deYUZp0YTbLAbY/+jnsjfj8
VL5LhTPRyeUsFFp0/CUK7D65IGDUz+658jxWzMQEuELpyHpIwYJbtGz60Hb1MmxSkhbFjtp5Mmj+
WeDOoHL0oDiqNc7NwfaLocZvwJBvz8Z8cBJMBLSEk7YciGw2SiDNTSE0HlZkBG0VD+UMDKNXwD+h
gHEX+o9R6OJtaW7qyN2X0j+14MjqnAIx9TVXRs8FiTnbVvKPPUlhthqsHdJCJGWAAHAZhep1cwMe
HczQOn5cSJ+HQ+fAjTXKXp3FKQ70qW3O09KzeqbooVW1oaWqa8OTN6YqcIj7Won8vPJM3uEIvGiP
pMzZmS5AJItsBMBlWLFG0f+bDwJ3rALDRBomsF54w53FUfc6kb4M592FBtdB4Dk7+fod4JHaJrRI
2IXyMnqaHHedtkU9DgEWeshTY0thzOqPIouKIWWCI834c23WwdZ1Nh5uP68/4m9ePfvQRG0G+ToP
DnZiQHPptU1WtqViTe7AIRJzHRbSDdMa3AEkPWu/8D0mDcpWLL9fUmjfQhcsXLUy7tK930pWOMuP
NvgEKzO4truRXF/xFVgDfmjDu1CWsdnzNfJ28T0+1JooH8dsW6J808oaBw3NLXHvMZMV/spBtWv7
+vxwNlZpzjQNn0QwQ31oL387SuO0ZsQ4QS1d2OzPeOhNNn3sTGOWsYpbxEVYJRjyylCjjk5uVnBT
90lEFmrgBdLzj3lhtUkBky8r10zf0QwQ1jBGypdRxUDqX1lGybZ/TXubEUba2dvwpetq1D97upA7
54EVeAPyzcPrAOi41mqXbRTOZWHbNxUWbszg9iFacx1KIKFgavHcrN8XlVWH9GGtkscJ0Yhmep5B
paRBwHbucmdPoqMbY8JlEU19ctDOyVBl33igeEerKRuIn1pLsljoxysq6a3/xxq66azHFPc/X5+i
kICi9n94+J+VULCl5r2JsRKVeE9ArjTvlibUorsh26PLFtttu8Epm3LB5OVkXJ5nqm3FVuDNsy7l
kjzQjJz6C1uRxo+gqmjFpwODBAAaOxA1nI0lBn4gXOiBA/IGvv53f1qLAuUdy//tOUCq4JGZIlWS
L+M4xWQEP0QSNInMwR7lRFV7VnIh8FLc0iIBWaL6QVS+ctjb3W+j6y9ludYWyet7FUn8lsGQ/5qy
3K+Fz50mT04hfnbNoCdgae1k6OpzsB5lSqlFqk7E+fvjSHiz8O7pYghkwbPi127qVZCBM1972dlR
40TSwIIyYT2JT7WQ39OPDuDseyHxeW5mfFHBp5WhgihHMp5q++nALbdtqYJ8n/Mj0LfWvf+QfOTj
PEYxPTcONbjsuJQo7e3WvCXN4nn61SyMjNwjBookqAdPVcIzfvYFQ3spSyZGlBKIIpIvsVTXN5ob
9yEW4l9PutDuMdXo6KZtkhFTHVYu7dp9J0p2+jdTFXtZiq4PfqsIYY/rRirDTXegJpH1FQJJDqpa
Iutz/86/X34z5Hnr6boEFJLzY3Ln/FDk5KPrjGIaAY3MjxVb4Q8rROCkZFjYD8gM0fkC6bzO6icp
nNSufRsWdn6BQ3CFPxg3RbgneuvzPqWn/mOCsLfi12u4D/dYEd4zJOS+l5HVvbzWBAxbDOpsUR83
NZOPFSKpOsVN9iwAG6TDv6EoIGtP3vMblJ9PrKHZXVlWF79ImWSzvIIjCdwHO44PsaXVY15Zuh+8
h0a9CROIiqrh4PSjgMtyK/E0wCaJLIf/dFl6U3IbX9j2zpTSUowKBr85vitC3lQUNAsxmQXZhg2l
7iALt3q+0CoC+AtiAb5nKs8LHg2Tp22xET7Yoiu640QdM3cIazmQX+DtK4ed4sL1qTujwj4LHy6D
bByLRMclH9SrH86iqJClCinpPuvuSvITu9a4Uuif89J7HrrVMgg/wY9SR933MYwsYwr6hN8CKwgU
WbjaPSy7379Rvkw+R1P0n6AvJkv1bgX1Jsf4iy7TNW2AOwFAexYRMylnn6ZwzoMb5Tu6VZcdb0fb
Lvnbw8n0Rx9RWWCMZrc83y6yFwkyBXJFng3s1c2WCuRWpqpsYDs/955oU/5ohERu+egcULhY7nAR
eGc6JUwujXGL7076FyzXoE+tppTb6VjrVE3jhLWH+PbZTZ+5hdsep0WSIGBHU/wuqAA1cpDc/yA6
6WkVYfxKQOdL+KYZBF7sgmNZ/q+GhTYQ9X+styALbSKHcA3ey8soIbmWW4qtRlVJx4EQueJTaCgg
X+souzQB5oObLJCUA/jSWlNtg3B7/h0MRXEgoD2zBoBAyNdZarDWRYyu6UVRZTSi9slx/e4lDbA0
DP+dQtOsS+ZgCnLgZGbbuMJoibUd7qPKyoGxJrbQYqq3Bl0hNuyHklM7u+E0aDvWOH2UPYCKW/NZ
oU1o6Z4NvaOcDKd8+i3tZYHDJhouga7MROCCzVkNV+Khfglih3zOgmlwemUf+QluFjyj27mgllie
JJ7Vz843wo5R592+BX5AExrPRB71fNIknkNV4njPt8e4GPdYSOOdyBruK1tBvDnj6De3o2Tg/5/v
bKk902rYP4cLoHlxLJWs1LJDya5PNK67jcLbATki8QCseBrQ/tRwMctLaARfgLmq6r2+3zM1CH6F
qQdYCa3ir7X9xBVnQkHCq5qxBSml3uut9rE0FN0aooW6Zs86ov7M2uYTudKoCoqv9Z2JHHAIwKwp
zHdzaYZfbPOwOHcktu08oTWtpSTiX52r7x9PlEDnJRYX1iDOPdKfWoHGgh777nt55GheX4sG5Tzs
JBgiOJEUDTbUH/UEgHjaeMLBF80VMg8FL4oLFj+Uwi2Yi5vdCDBPaVN+E/XwzsrKw2QW55IjgoSn
+C8dEByWe7rTItdvVWxE5/xK9VqMvVuLaNAQkHOmSzq2SisVXzpSkOYEU3lDT27xBGdj+fHcVMjc
P8m6t0aBV5Gphs3Z40yWXmYPlY5cCFkxhJfAi8FdNs8Co4kG4MZw3h4aQRPZ4B8IpuLt/Xrbwfuc
dFSQRmu+oB55ijqSZa3PEKEmIdsu0YLdXT+/eIrze9c5LFTj/niY/OtgLsL/uy54yyaQI2MRPF2R
ni2UhaAAT+GWm/0umbj4t/uSC66YpWJnCSWF/65iw+dtYAiggYM1pS5ZJH7x1/jJwm+t66mEXOeK
23C2mkcnI5ES/WbgMuXn4mmNznsI5+28LPKB9+yvLZuWCJ0/rur7wtkd39vElMjbtiNlfg4DVdPd
PJwoH48e7NJA9nH7/2arvoqXKy0tfHiDjvgpWB2zxMHan5kirJp16g1j0ut5DlxluJ4qSICH5Guu
d4Zv3DHcJRQnjX1weGcCs+yfaKzYDarusTA6GhcUbUXWKKHWFpbwYwWdrf6XSXDq4vncYs7TfqcT
ngVDoEi/4CzIw1QaKEFShr85CvGa6brlvSdR9ayWteTFDZNKBC+q/Ll73nk40ZuIFZBfz1MQ7OeZ
/XeLKUqCxHRm8Ynn6MxSgW43q3aOtkhAmIOJHEOHNZXn5JEJK+ZxRxVMybktYMQhiKMMGPph+0Lx
/F9mUcB7mQPVm7Lnt7o/DwGRR7nxqvsmycVw5UOLu/AOM35nEUTkPvabl9xSQHsdmQsCrs8j42yn
nxQev5RbONFzHJFOyVL6HGOuPiaueFJiuG6NHDl24Lg3+TWdBnXoAH7r/hI4OvT3fqdvU5mnBmgb
bfw1aN6G9At+MruZDDbtziDLgd/Q/4F9yFciMk7lUSysZHMLW61Qv8vIzkejV7K/v/PAmu0igSCz
qaTOgsbfryuLlremmzd4qpUPrmWt2m/1d4WMixuDgtukqdLpeqQIVHzLaSKmr3iRkSJc+6rTfvxA
2QZv4GqHs8hOCNJtpOQYOBkFisEcmb/28ASmUlC/n1uMQ+0WOn5gnx2+nvizS8aglvWyox96wamx
leOmSKjL5TsY0HGPWdsY/U+hcDen5qqAD4s7fFvlmuOm9tWNpluJysszrXNcLn+M06SaA00T+s4R
34YIwBc8fdgWpgfyZv1JtOR1tuaz5qYibRWAH7Hj7Au7Mzu6l2jHS+mQuEqBiQibUJgYyihcpVEc
ICo5kI4u0lSKFpnpOmTbQAqodIC9NkVln0q8ziYWLr8Ba5Cuufx3qXzvzmSGsOs2kfG7RhQa4mud
nUEdschFN1RRdHMQUXp81MVukewPtVt/0eCw6jeozrxza92hWA27gZ6+9up+MEeG4lJlp6ywhIR5
TfxezX4jtm1hJTmPNefSpgPTAuALmSU+kcdBfiTFOMdtgR+3lBI6cn+dbY948DyjV0o6qWuIOKgw
yHTcd4wZDjui8IVQwt6GA6vgzhNBBbZSZqhFoPWYwLTVFqEFRV5v3KRy9rW4UIpwJubXcDto5HrR
xHPOaVk70/Juj6ut7W/gISroKIJpfo4kvclRccw15mpBv6w/54Tchhg9NbAB3V65sb2Yh+nIxsrb
EGDWTED2mx2W3dASPrR5XzaXGHBrtnHvRfCPN/6XOgsvaJQgagT+1yYCXHKqx+c2EtQoXIPG6l6H
mCkZCpfJqHEBUT3GJWf26WRfuyW/Qf4Hv2ZJHIU7Lu5iFr3LxsYz3JdWjvc5af0h6gD9IoswGhAs
UdacU0SEypvdA0/l9zPyicrPKtDCVbuHgUzLPiXqdH+sUXE7yo5LQKMOzEZbIv2ZdiYpzD3qc8ug
EIDBat6gf4BqoM1e/ALCXEtz7cl05qixY9yRXPQR50qep6SE7h/ptrKyuIiAqM1Kp4n85mPbWoX0
8f6WTnyMc5h0t/WliX7W/dW+6IIWVTjUsUA7Ni/FarolcEDe+s7n/AFIe96vtaua1mF7Ofue0/0W
VJOGYxNMrzS/03wgHbQ4cwKV2f1/X9NEbYSnvM7BwttC3dSRd1hrIIpTGW9CVqNOBHS5MxBzwhfp
IzWiSy1ZUtg3Xn1BO4RYvKXiGKnofU98LgxjkEVg/dIcRjlNYr66dtxmNydCGZYdKh0cyi8In8EI
0dPSlCKfzMOPPQPj9Xnw0fnMMvPVmvRbOYis0gEOtK27rGNnwwNYRD8Lw8KI1zIUgl//1nPFWaBD
LHSJa7LArp9B2RtPxL7o4LFD9WRWHoUPDF3mBywhbRvUogpcbM3B8ar4ykMhUUOrtjgzUe8ocvnI
Bt2SE3eOnfHHPDSLadEfQtsg763fXHPQQriaiLzjkSIJRRSeLtbkLfTmwl+3xfJNmujCEvMpgzwo
cNF7M1GLxWmnBfX/D2ksMUClrblHaMlV+T9zg87V6eFj+HI9fL52DYoAlyMhCHhQjzMNfYZ2xEEv
pnhHmZtStiRed8fkVomGhI+d4VMoxPQfp9FF8gLsdRWrL2EesyoPo/HFpR8vTaB/ohzHv89+yVQ4
mkMzKpRoIMxTXUJO+M4vLq3ZMgkJ5RyNFQiltVL0N1Y7SH9uQEG89wp4lvMxgKUvhYtHAySfk12u
NVL2XD5qwZ2/yhmHfiMMlDFMKGIUyQZdHTWHCAfxCdqFSbfORSabAYeAHaGtg2ukegk3/lOSeLfE
wHxTABqeGCo6DQUDPfdaBVGvWuwfeIdyzSlUsPoVMNYX+pkaQEFx8sID+epWcGNSdhG1KEiAtEE4
6jzrB4QDJ5wlz2NjIiV2sQDZFiwGeRyri+4mdsglzOPewA2G9V4yD2ljE+QdUKSGHAzyWq52HHzC
e2+lWZFkhdMzOSk85EUVkTVcM2J3Q1KBe91yeu8nF9btVAOgyJiLh1Dci2tsNTasu6K2Vy9VcDOK
L7khl5zCMSLTtZZzggn/MdqvEPVwgUWlN2F5fc4jW8O2QWCOPaDsfJgkvcLq/yucx7V9GipgIhVu
JdxcyFC1XY1+tQ/yY7zOGStAreEo4Fg6rfXcR7RkVqY/G7lQNiCYlTroluz8Uw6v3Mgj6TZ87gaf
GJR6+ZyV3jYRbmo0SIskow6vwPUJmLa82TdC4fThXLny1KiE9SVKbB/RjYsHaU4yT9IQGbMY3AWG
pKlz1bhD0/BzpiuCAiuauTAMiFhTa6bVkTWjQ48c54bFxizV+/gHYGMyBe4zLrkqVAKKu/gc7d4x
0rU4Tggv1CaPS/x5k1wotmGDykAzceefaOJlvzulTEqOkqwhM+T2o17w3EN2E0iuGxIJvBSp275k
pfXzoB2+ZePIP5a6DbXE3OvKCA3I3zFy8br93DdHEAsjyfhLvTR6K8RAuMyaOU1yAoZc3lQiezvl
w0RkPOwUJpEjGU4dKDrC3JrstbCJtgteyrD1Q3T8/PJ19cXGbNxXYeSfgvn2dVMKcuqJ8P8gksOs
AYu0c5+/OA/kPpm+FCz3PjrbngXCzJC2Zo0M+08W77B1xYzxQOY2FpKBSui1whMaMQbdS1f57vfE
6QkDf8ePM0B+k8B9G64lZsB1wRPa+0Dw1LPi8oSG1MmA5AAZTFl/tRFK9MmGuoMBq3VihqNgW8D3
fLhXSnYDCVCftm/a9bjR9sjSz2tJu+joBg+zfvQVlzFPpekMlHsM/1lNlIZ8UbcyuvdJwefLts9X
OVOGp+Ppgbs971TOjTTz89N6WnmWozDm9gTkY6q4EjIaUigLSXhg9fXRdWfytDJ5g2U9ua4es37/
L09eQa8X755/fUvNUXTGuw2vmi+XEzSNSVSA0TAWD66tehgRqszRxummf50/f93ZUqX8uVqWtaX/
oxESF9surJz7uY2hx2m/LlrEjfJbJUrrM6D6XwYbOCPUqMnRZ+RmxbzFqDZCxfqFEqlL7SgXN1fq
Y60o0HHwb2U3p6N3kcXkbxDK/bAB9g2SuIJbggDVPc9YUpiCQ2VuAt5G8JJyDWZUIkQXZrC7rcsM
04beixuPlWWkujsZ/1WDPMDftIuAPgtdlDVSXxmzlgAbiwLs3S5f0VXTMiNyNAjF0qzlCK2bVR/k
zjFXeR5Qs/WKSpmATG013OzKXec4w13GwpcY/tvFXtJMF5yQni1+B7nPD4PkpJC5WSJTHObxCq/m
fi8Nja4dK2g/8qe1XN1bViw8FEPLQWYVmUAu3r5a8T/uhHuC14cjaDIOTfB19+Ok/k1lX3VtPvOI
l/qb52dgGxBIQf7muc4Ull+Ld1EjJSJWMVK3wE+5zaP2N+yVgnoE2L/Sos66SCSGHNoCNmda6Trb
1/PmJ4kXw76gCvsKNGFgTbSb5YQaXAu5V9CbMVD55h3L8HzO3u4FmuCe6FKq6FidDiSSYoGruy2U
JI8Si4BUjXb290kgivjxxOyQtU7LlmQRv2wirns7RwJqJQe3mNVZCJN9Pbba61NVAmkyLscbJ2i+
rBqOMPxmJ/2FdBONoXJuUYXXQg0OMkvNhVlhpzVQvcV68kaM4lvNbMh1x+14lSxtuPA8aWqA6imo
bzUF9L0ULd/dJOQthrUkHtPex3FTJ33lBl2khmDb4jCnknqyUv3MbZDfK3UyRqejxH3etYv1NWgC
3xTsdDo1CGHB9ra/JwaQBIxGvBcg1V2WJV2jWFXx/1ZLKHUIQqwJKzh8b2njGkxYxiCJ7eb+UuS2
95ch31bv/2BzggkaeTqjI69Z5r/BCDKe254wYiI+nwEgvnhSdCw4GXLEjGYcCS1TySZTz/N/xD2/
V+1sTs8w/A+BfBywSiOKPJYqGp6z7z27Hms6IaOJ/vHygisCMiQBtBaqW0cW0aRMEjKmKyLDPVE9
NLAU2luoCnetn3KmttNVHOVmJQ7CVjfk63dRLggX6Cr0s+b8r2nrhSWRLzQ5QUc43TJmC5ERcoyE
bXvyrUxGs3qXXKDg/n/Lf/ttcIf329HIbr0BA7S+EMo/mck4onDBS3V23k1NKh9RzFojaYhR2BMu
cfghFrMWrNaKm+sns7PWp/WuYhh8m1hO0AEKjhVVtZreXc6mcGJPaMDcqVfWVE4aUhAPmcJyequ6
4T+usP9rH3I/3fmFqBmJCqNMAAag3eTL9ZPuB5i54hZzJcMaeyEG5MZQ/QLNgDCsY3MyLgpQsdAz
vV7CL/Zw6CY/aVtsJyf9wxGEXl9D7JaHnu024cIPINREPraCRusCXBaHpTr4xM8K2RNP+C3CfERP
VMPd+JaJrv3aJkYwHzbhky0RDo10kauAjJ6eH7KXn6+jkqRf5iM29TXX789O7/tA+cser4Yvw7aM
QDYi7Acb74b9z8nyBfidTo0cyC7IJUxssAGt8ie+g6NAXNHs1klq/YHm6nM8OkqD79UuG4LOjAVy
GZGjGwSkqXaXapxFCQ50nnuTyZtZXUVP3t7CZy3S6GS/vXxAkDn4L3aAV/xDltLRWlnS70WGD0yD
oITIoLaYvlGQxEqUIjvyVPX/Da6FILROOgG2CkWp2+MhvhDLD3P1/+HLK/sLTCVi6scgT74yOgSv
y8lJXGCje5+C4dy6CIm1YfqwQuuhDNyitK0W5FWm5IOqeFm84fECzQS+YElTbyA7NNi2RNw5ebeM
uOWmT55hU4SrIHLKBfrvUsQdixmTzD/V6O1cU1cGmJDNG+Ed0n2AzeOE9OWNWMjprCDDA4GnWOoF
4xK7deQvG3CVrTmA/dWXQCyN9K6mQd6I6kC9sHimiz+uL1AoRdOLKALv4LJR/CbgOvwA43bojN8g
XepxnOitwQgbl3yH0QevzgaW4o5GLIunYO+iC8mbtxnHoDxUZDLZUyMXTeksKasZgjw20pe23+wg
1lkuxg4r7y9GcilQEUT8ZAn9J3yqfsuRjzDXgN2jGAm7lUQ+Kq2D05N2ITgGLMo/+4nbsrIbV9aC
zhVhVbx6jk0i7DFHKMAeMrANdhojHo/zJz4Ax3o5z8PX0y2nYAAGgU/OvWvRh1ym2mOWewXYymlG
Q7z0IJopV5BKvgSELXz4a/q0xaZEhnNLw1vATx/pREG7jNbAo8r2ylF/+Jw4o749kmif2FBWRNjA
7tjQJ5LFIAIlUlAES7Svigo/hDzFRP14Hg85wJnEqhmnBwgz62a+UqtmdPzMZOUx0XIqMcssPvfU
AWwzA4+PEoZkt3CzEtiLkAQ2xx/f/w2D7S8IFMtIiLtNRPgktGwN79tJAAW3pE8OvEQeFYQxjtd7
HC8n1SE3CaqyzQu2bvfOy5orMys5Is9MqPKlI9Po+2hvak0fuX4ivL8VYEFZL6CKV7602AxUbEs6
c/5VFAkj8yMwn2E6PE6wH8LksD4JeDll12ioTKn/1nfWaVCe6mUhhualBmD1M2+RHnazxefXAlUl
g9a4GfmPTtQcA6hLQ2jwX1T4syVvhWwb6NmdqKkdbwVARcGwltraL7pM67/LfhtLXPMD+vEyjM4X
+UO9rx+rBjjb6rIYD15NPKHgdIPn3DJSorhkRwPR5rNBj/ud6Ea3wvoVhGmWbH4qsPdifhp/YY4P
odSZ6xVXnoTActvG7RL6DUwuJBXkepY8XmZeVoGVdizyIhc4g8g9gLp7Z9Q8MLTh6h/SP2oykfLU
KRnU4tjrBV9T3immOFT7xQ2vKRT99uv1HojFAlyMYyUOK/3dVu+U0gRwpD5Bko5BqedL5sXRK5n6
B300qrHdIlyh5fePUxN5i5Szt7WS6/kQHZt/CHua3oD6r4FjV6pYWaN0m95XZCzRPHgJg2dFXIUn
Um7dOzTFahi9xlFVVw/QP7pzq9/eDsBy3MCG5+1rrunVuNGwUXkGQOcY7f5cpNMdSX78uNE0TwsI
nBVBJBZTRJZWukr7W0UkK9EGGI5h7vNa5idfWD+az+0cI3fVVIddRQHBZt4CTnVfTqaBRJPYgpkN
7DQhWkHR5uCljNHDEGIa2+hg9uqS/LTstubOYsFzLEy0akk6EEoM/ta2IJHecVOCen3pfXxMrsK5
XJuyCJAOtd+FffhxWpkLfWIE5LIJ/SaZHd65gTA4sNVd1Xm/m5nvuGRKKVcWlIY7/8e3iuqWS98Y
PAFIRrxfYcIt42aS6RmFDHSrCoWZv6s4LkzzltPFUP80yBo2sXaheMcHbwM6OeweWq9hu5ZST0/Z
ZifQu7Kt7r0Nto3NpKa8mgGHvOr2O2oDmvwYXh2Fua60ezg5paqUGFeSQHjSe+fg/yYJD3NM5ggm
eE9Sz1zuUHnwQ2m5/+BxTIGUgo14+Uy9M+QldMNedjmDMd1nLA4kC7EqF6REoM9jUZG7O9gcQjYO
IndKX7D0PFzZE4R0/Z+Q4t/hr6UBpvKPvLLy6OnASG+wmo4yqCxKHOs7I8OmoborCNDSzr8fNfl+
0+8/zIcEKncz2piSABiJSJ1yPkl/4CLfN+CsOLsqvzyrcP1gZvHlVmc9bLBR+xt1MJKUB92pAxYe
Ju7r6hW6h379O1WqxbnX2AjQR4a3/nDNlbTJtznAmbE9tYcwJH0GIQf1r/zT3Su8WyTio1nt0wRR
N5w2EzCq9fGsJxrZoSFHpWP2tj556n84Gg2a4ObNmZQmRChvZAwMsUnskpNwDjzt0RKZwg4dLL5N
itmZTRsMT8ek1xYMimG5hjKqdBVZuEmXY8IjnnDrL3h31/3BUc3lqm55AWn++kQ/p56GpTXTTN2v
OqQbxLQjdU9VJqM/594Hmog33SPzALjatmaQi8yhr1k5IZm6J+s8IOgWVVg2c3sxRmrO9L7pm2c0
NzDOTWoooVQDdBnyUn477J9/Yx28BevBZe2JsY3VXrdY+8+CdPdnKkVoeuYj4Rj5rowvbc33nWZg
Rmz3Q5+Vuw67dYJ4EDHCJXH+abXMFh5FvOa77t6EN3EUm/RO4Lg5NFseHzqdpoenzV8AmR/Ulbs6
z0rV4EoBgW2XCt8ACLP7sOTS8XqG3ChJWn49j2eR1fYq+ia1iX2l4Gby/GzMXoJ3TxTyma54V/Pq
OphPoLFoqxSrSiSnW/NjC1N9Tz2BrYafBspTxy/sj2178hUwtOt18Ywyjgh0vUReTQHpho7EKEo+
SBV9O2bAzRZ1f/rupFqlqLBGy+zGJt4t+C2TlP0xy0nEx1s91IohMawfNgnKgjfonCRifKg/zSzc
QVe9Qr/xi7NvcIgi+5s8tukUU3obJmmHeMiFvkotsgatL374dwA8AaZ86cpWZrI1hc6wKumQ4r3q
Re9ZAJRHbYUuvj0n6zD46mKJevjKcFXpbbmwFbf5AMHspkkc0D3CDS8U51ONVU8xaULUakoT2J/9
zp+9ySYrUlXTUenMpP3Q3Wx6oX7vCze61+JVGQG/4lrbxBBXX8I9lQMxC4FXGx2kjeb/L+40B/64
Wr24O9VqiJqlrrdoeBF0v8zkmHZHice+J/m5kFabJWBA4oZPNWCNVn39/q+p0ofrdCLqj5ESz5oz
1bhtgSvwJLj+K+jAnV/y7ZmWGE8wR0MI13uOr/Ap0mfBCM0me89H0tVY4K1uNndTIeJFUkJ5JKuS
D7S3OV7Azsg3uGt8tXfCdTgpL+INm248vKonq5Ub7FNm9i6H/LVHA2C/7UZ619M6MpEbCn91LNr7
Fcl/O9HROqHa/6SzPGL1cqSxdBRNMSCn9BnDEtsWJqg93GjUAi5LHGzqbg6ECbCCDGZw/e56b1Df
mGsE9dk6V4H8USf/ImI1dQMYEGbGn0OMR+xpHY8XvnqZ25cwaLilYhIYbIpARKN8/zvCJnwSPBDK
de+DiqM6T5iJEel46XSyPseR2PTXONdSi4QkQ34fe8j4K44ttySMYgZaBXU82HEUrAWspRbISowj
EfthU5NzR4ehpsSOZkyUw4aBmnRAyJBdvgC/5dme/9q8gaADdPmOg0IohGOn5sy7ONKPb1cnuuNj
L3D6ANDQuyWZih18a3KFRjHdAWkLq1Pmy0HFHtZYf8H/ADNNfmEsPMUXdxtfOcJAGOCLGOtFmAaz
fvGfnllPjLKKv2Ur85VfELsoUN+FIIA6w6K6z74NAmONaaPpxU37GfMJcj5J8rmP8NSef1qK1WkC
oEIdd0cbvzEDo0iSebPsri2wtbVjXtpL1HqRcwPB25/vjnuxaCSeLNMShAhSzqtTZEv3YreO2XB9
t5+aGFv1Z5DKprdwXZpy/kY9ENm9YeuOeds7SVtLFifiPT0ioNZsPrd+lwPi/Uuu/YxxO0mEP7J3
Xf/pKzYvU4LJOgDCBVFii0M2wjikkemh3GCEuHb5VeLMkT3+0UXEiwpJU1gkUq6hkYHJWi8wNT+l
ORutahU1Lzi12dscsx1X10byl5gcNND/CBXJrgTY0EBpYV8gTlMe66+O4H3hHeP2bNl+m5MFX7jP
AAo92MC35sQgbEQnFMKURVZ6w5/q9ITXLbC3FcqD1ChhzmVd9t3pQmUNeliti4SuRYx9kUMnL6/H
j+KIRb0I47LfaHIjCuh3raVWkRvUHIXDSjzhg9JrnA+f8HCeuVTdiZGuiuA4uWdDt/eECQUO3/nB
6P6/QgB9KKkupxxVIxsKOYbFqt0fHAT9+Y8txkDTV1dxyYpGLC/L0Ef/KQDeXmXM+yaWXXmSzSXG
sA80z1q3GatwEABi1Iz07fNWMcwlpaQpO4BXAiBafVBkDY3u884YoDDV/3Wh0XVinv0wxrgZWKdI
8KMjsLVLoCVN6uCkIYqBo2nDpqHaLQ4bPNEcL6uS5hGq+HIai8cA84SZR3YKcmgli1vmxh8CNiYP
mwDKdtR1KRlt7iv24+hKQNRXSilPsYqXVGz7xD2eu3AelYaV2jwxiy0J+YeYvxFMVJVWTNuIxIla
eQvzMrxOWrFjfB4hdMxbXciRzCLYoPB4RELyvxk/40k1ke3smpSiYiKJHEuOcImSoz6Hz1VMkNQs
qLGd3zMbHvqH9d+ISsCp6/RDDgSgeefIqiyG4p/gjVBllapre3Sh9PmbYVq4Mi2LZ7irAqhY3xy7
un0w4Rj1QY3SifZ+PpL8FeTOY7kn2xKjCPsrU81HC/hB78OsDuhWt+w1SNayudxd14Kb7YQ1ttX1
v9WxorKwQN1985rpqwUAPsbXaJ932J5p6WlHnfUqUYRAKfi7ancmZOoLReRqXrv8Vk31n92++tjY
MX3JWUOeiLd7jl3Jwmnay+XAcw6xJpzAmF+YeiAl9W9FCK0rx0y3r0D5x3SJTfqFmc37vNi3/6pz
CqXNhY6VvhS21aLV6E2U953ituJDezNAuEsbLCZa9N8SAUY1AUFmybrmUD4oqLmkbsPd/dXR5Dct
pEkE9XFHxsxuMK9xbcTG87wetRfMGIUZChnd0rX3Y7VrvwvBSqZc6dkgrbcf3NDUYZC6CUSv3UoX
g+OLA42iSdZmAJrZAzVnuZ7fnTLPaVRH2CwgpHykYRKg3bZ+cMqc9h2lZyONdigmpbWlpjzIXLNe
TTulygQ/bF1lqHek2H96q/Rvy08DRWdag0z3tbQHtSAB4Z9nQUB4NveFL+PUY8PLZZoy6UZi0uhU
RBoaUvfA1LnU4JLwNdYjEaJSECXwcPPouWc9K93+k4yOOppFhc7hP8TKfHGDtWl0vY9rWU3hHqDH
GMVl1JHakNrXxNd5j1d98hpXvN9X9Fr92/YGkEK0UGA9SfieJA52NP7Mko9xPpSegD+9LfCzKx90
KiV7y+xO0opLP2VRFuQ/bNczoOQxBZ6yS4Bv2sH/xqIUv5uvIQqML+Wu21oBgvTOBRemmx7+odxp
ojWpgpY86/nuKSgzPcAITvin0ViiYStWQtzs742xosWhIZ7GHQNmzUdW4WS+FMzbs7jFRjAzJ5z8
a/svN/jZzo1Rq7K1KOwuP6ViKlIemWNh89hAdoJ6XokZv6WHKRHKtuqEejJryN0uXJV4JB21kCxL
FtluUEeLRbP7nnhdqZXtJmXUQB5WIcRAACmOqQBuJDbAZgxlcFIbnwJCKW+3xj/i5tT8XxVuKaNt
YeDtyXTgCZk6lrNVPtZv0GKmOWzt6bXZ27XZD2sUnhtMf9O58Xs4RoKCT0U7dGyQpfwD+vePVgwL
4+gTFJrhBMl6byhJR9MM4PwPBQCrCwAk8pLaeqBH1YrshTxPjisFsrr7jGYvn0v1gUzz4UEYh2wY
3G0kzx1gctGWlzOreSObrzt/Yhze2DZcf5tON6/CgMCcBsGeMLoEVn0Z+gpw1CFC1BzSGATyh4TJ
0K4u6wk3ZPZPfqEBJQSAUZCwURuG+cQQKywf5AknogrpMqmjz0ZWj+PMB6tT9NMsWJ27wNPZx7Tg
FWFfpXOpE4e/d8DR+irigRbcwl51RJv+2QXwp2ED9lmH6KLKJvXPvVJCa2EgNVSmTY5FWUwJdMrJ
XOLdBVystorUMs6W2bwCXQhheLNsZAWkqp0esm11zCKdX7W3SbJ5uI57cayaeWGqu4G/SAfv6MkG
bueW2CzJOGgqT4gGa7aEwiG4WcjS2WVq6D5NN3oMVs1Obo5Yiy15sjpjbriWYy3gI1RyqFxE+5G8
sGUPhMq18/znJzIc2Rmh3EuqiLFBTvgj25tD4MuySAyMdUPdhBvDFAT/0ii5xeI2nV+f4Q9wxOsM
L/ZQX0UrbxJbH/g6+Xj1+f5cFdVOwPC4dcDC66culP67XUeQBYXkqQjGdJ74W8BRQtXi1F/1OBIA
fEHZweYIgC+Zv2+A9su97DuUP3i+UTNunnyuS3/iA1Lti9+Eih+31ynBJGskDh5mt6W/CSMDXhqR
W9kzzjsYNYbmnhSCokDlalKmcHgae1S8uxSNctspxEL3CGPN3GtcFzFyUraoVERE0XYkKKr0YD0X
IbytiZmcmUX852FfmYTP1VPL5aUWRXL7+IgWPSQMuu4x1q1gDmQxl2GGwKlu9YwnFdLnMgrgUAho
p2IVNYS2XPqXgtyNBjDAG5omaM0WQIqiNRfRKDDTo+4kTbw+GvuanqMXI7TNI66fzIp5Hua3egXA
T/dKujv6r2T2beWemcz/O3ZZvPymZojmO/b6khYwvctQPGCn/6tRJHHO3s65BAPxqfBO0uG0YtLM
sXPO/JWLEqU/9iU9ftzS62YdVwQ70HCEtpxhTdGdL9fLXcyIVMQFQpByc4twEw2x8x2aNsmytmAX
Jjpgg7zKuWGH4xAPlJ22QeToHfkEtvGD2C5kixkahYz8F6J+FL5GINR+ucRsa6KxrxQCRMyv6FkE
Iui045YmDhuD9++aYAIyJqdxwWBn0IJpiv07TDOtiq4RS/yfokv98v5KuL6Co6j9ikaLCG8dGl3l
lTiPQk7t1mCf+UeXsXb4j46kORNb5gvlkfQpFVwuf79eusjtkAxncVyuqjffLZcgjoF445oNpTDm
h21tkPDKI8FfTc+YCbM0vEDpUdZo29QJKgB0F/BqrYvXXKQdJdSk1ghu2lW4CBHuNqbO0aIsrPD+
wzLMo9j8E3XQjY2IjGKeNQLB7ASYnDqfBT4rGhU3jbPBJoaPz0bRvT7VBKjhJMTa3JyIilttD332
Y1k9Eh4aK4Ol5SEVDqOhmcnUODAgK2SZ4FMQbVgse5ofW+yc8G6suCMkqIJXKM6HqchcqBkc0Keq
7wTWZ46SGJUBDvtQPbDzhqRVaACG9urBiM09hNJ3zTOkRWICu0o9w7dqHRMfbhz57Hm9cJnA70Kr
v9fmuU57a4w59MwylWrBEerGTZdbtKU8sGXHibv7lrzApMUEfv+dXy/8L1ugRzfPYjQmjLyZq5pH
zPFx/MBi9lTekzZrdSXk4rXSFWKd0PeYODO6rNjri60Emh223rxtVAkv5rumpWhCxFZVbm9AqvZz
DVdI+F0muHoce3AQfgKb0cTcLF/a5KvJucY7/lmRaDCMUgdelowIJupOwICi/p/CC87Ll0c221RL
PuIhPXn0BvD4GEQoDRTBSAfU5uBIZvPpXpveXwIpzOekOd6fnVmQvkcW0j81oBamyfF02pMFy4mB
f9EP0qPaCIrIUPc+UfvuryvqzTQHRN1l2Hi/PxWYaGhuga06EsVtdihu7nwgBxOs01vpTTDFhyV9
/KWV5uYZ71ABzCgC+bgfnMjEZIPKoYSbGMF1VXe/DLCNo+sGNruEFekcxmQbTyu5KRoCiKTulv15
hCvdDE0lvO1Ab++6QR85R1sDZw4d2Hb75wBfAHvdiFwzXp7OeXgy4z5ZW59Go2I/sqxStqsHxfP+
fR08Zzc87YqwOOHhUtZ/ABHPX3gHZxU91Dc0PIyIcsQUL5De9Lk8fGjuIQaq+kacN2585kybiXPB
JccuAdfLr7GUYOirXg01V7u+TeYadWlaOZS6IluuWCSLJ7ISvVnbcPTeqed4NxDAw4pTqVRMtrCo
r5qv3O24h84OaDsdHCADA0u/08Ch+i15Altp++2m7vVNyPvznI+tdtaGUQd231sJTbCctPx2LwCY
bGgfnIP41C+J4FJ+xg3/TFoNm2wbyg9R0zTKO2tGm3TT3gIQHKP8ciDKixCt/I6/FbOg8b1CNEye
iXd4v0hxiDJU6P/sqBqXn4BVJnn3SKxZIjlvs0StU5vCSelZFqF35pzbNc6ZnPQSgarHfWy+FLlm
XHw0IGe3/hZHnyv97dCbS8R4deAu0UzxiSh9VKcTJrPNP0vsHKlxa6fsNOY/GD7YMWkNFnkFXQwm
LqqvBYalT/5cVjlfMHGLsnd/nj2Rz4WUGWUAqLmKZMJ4MuA1yyebPgypj2JLNMZTOD08+L8gV/G8
QmC4GxUJkTImb0hVbldL8SyMUG3qV2aURjdpDmUB5zfh2v5+w5ThMwlRPGQ12q0wrJeQ87lgq40s
ePj+DTNQITcEaWa7yt9fWiM5KS4DFN3pTNyZu2jAoKDAYqdvfyF9YGsCG9DFXlVsnCRhVjlZUmhN
ppx6TTTXTRvn8F1MJHhvNxGgfglbty1S3TnhXxEoxf6EqI9u5OhppA6cojbe7/wg/fg+8gWSIxkr
adYLIAuP5Ugo7jTjybg4zKdq0lTdVEoweQGKoAHnuBOLCCmC/Ys7Ihm6eizBHeypA8gtNukc+IpM
imE5i3OwVBX7GBfEraPjy9sCn5XlUbUlt28WpC6bjOFGr8hcrQXlU2HDcNgs6RXuHs9yMTa9kApF
RHRYTCvuuXVHk9U+tpSflYRa37r6ltw6GkdcBTC6ZXMYtPAniD+lD1kws/axeqqifH9jiHn+aZ4y
0IdMgngBrDBdZi77wPQCGZxOoKhkb3yI6Eq2xQf21MYIRDbgAEuGJr/OgjGbU/9EDLKqbczYoRlR
kBUTNmggYe+uVIiPt57lNAlD6pap3AhWEcFdhXWIsB+OXKuj8QTeoHWOvmQ3aa0uffaQG6MP3l0t
dF47rqFpN8SwSNFoe8LbqrGkcaCg5IWNdBDHwdfEfk46s+df/GR6aXRrl/nK+/IkOel0slZsCzP4
al1x3qT07LMHxU819pxhqivovsB4yxdHcbr0qo09HsElcBvZvIjS3L8aTQIb20SMCKU5OY+/a6d+
vfqcO1k5Hj2JISpmSbwmGnZEqWlNIZ32gWdRfjbABB70ohwjz12+jtoxdRAG9aX8/8zgqCnJ7baE
3SraVTjus06or4kfoA2+FVPpXcQS0SuKhq1h0GV/zr2klUnaqobN51VgeSmIq+AVhDBlO5AlIm05
Dbi15UoL3G2/Gqs2h/o3J4qFbyNODyHENonkTIUaf9mmzdktb00OD5h+f9I2qZt948rigYFFZX/5
imuB7dTNYGbQoO6QfaSOuqPsjFdz/eiKcp+GdJ18HuxbK9jkFm98cn5gPa6Y9TBlbMfnTGBc+OPT
ntKP1RG29Nw7rRnqzbRQijtBHEuS4Gs4NZK+cxkeqUq/jVYgv4Wpabymnm7Tn5/Mcz+JQlJpW9Lx
gho0wuVSsy0O5MzknLkRJvulKyIPyQCBWyIYesHGW6rIf+lPR5r0qtx5BrOq/vcz5XUco56G+zjv
5BjHMQV+Vnp5Fw4rsWF6tZgMeH/1NU0o3CGq7sbCtezG389wf4MS2yYi6fG2lnjRppWT0/BBbDx0
SQ3ojBBOHWYbsi3pH3P/LHCsNg/x2IPZ1yD45Myg2/QMC3adrDehaiwnlrsCSqWdd4eEEq6G6c6R
CvnKk18h2cM74Z+bxiTsMASJndt6LmoA6B13cLsjwkoqqOWeCTfz+TG02ouO77yvdcen/oRHRgwX
hLk4zHhj86wcNACQxwSKNXmgBebEERSVJQ3OmXMQV0xlDrFjtKD7q11/UnjBtZFGz4Y2SAPn04A/
06/ht8vYO2584wBA8GoYJfb0+3p0t2A53IBgg/Zr17kTccpjE/LUK5Rc/QumdS/iOjyvOWGFG8mn
8jwkHTuUtB52jLVZ9nNVJQXyHmI8VulrJkToSBfNC4kJ2BNxkAwysVuCECRCaGC6iiUnvzgI6wZv
sUJbD/WxcWdgff9YiPPAu/bCOukulIYSZjgoYmawsIB47XCXmBhZEjo1Uf9K4iLlXKckT6gGm3KH
WiX4Mdm4v75/W99QwXagUpeJg2S1Itp3oro89Rd1OquSAbCFgEeVROyeAtxu8lzAOWLK5lZ3+fH+
uRVLr62c0IbXMVatPrTOc1cuvkF2TvlIKkBtjUhmm6Q6qjUuUl1Dp1KQD3l8+icoVMwkFZcFyAsN
TTQ7rJ9/i3Tc+PR19ep/jus+jXCpMuQDAfyR3mNqq974isH8HaHdNS977ras93T+sJ4mqUD2gm2R
NE13NC56GDCL/jZkhboHDSakAjeEmg+gHDPADoEd7aSfysoiOaVNa3Whg5R6j84dj/6iPqneWYSN
TR82d1NVoKJ1fu4dmJT0C56RJ8uBC/tAdtF8oB9nIT8Fis9EFp8q1SC9mJrUbq1Yilom5sTjnTNc
KtM9CLkv3+hVb2K8ACZr9DzVuZaBVi0H9z/rKbxkgu6+yeiaYUT+Bf2naIshq+iZoJUj4zlDfC5C
LTQb3587cR7AW/sWMDcyxrSuR6iw2g+jAq3hJNHLk/swMFZ4DTpA/oVg5lwPDFtbAck5WyTXGxhs
x+05YKzPuvppbLAiHyadxTQLXDm/Wkx5K6aatnVxFTtGx3k/ebDAGBuEPAy4zodCj5GHSAs4rr/W
s7ymV7yONSD4uLcaHJ6zL2Yne1JVc4vINgDDZTNgMZFjt1JhMg9eUuusv6noLMkijUwWxBNP/yPk
O6wja9YEU9LV4is0sctGYXCfrrm4YF6kkZwxqGgy/dCtv+Eyqm0qWpiyDqckL1RgQDRjpFQWwFP+
2y/nzv45XrZ+kA4jw4QEKv8GAC1b9EDMqNllCVM80dNYdPWLfxy62NO1Yo7ixZ0tlprd3llgmXYE
YVXUCfibdnIRHOEF1kkmwMWSjxNRLIYW0C5RP5W0Yv8LQcM8laHDA0V0vD4dDYmKU3shHkeyTnfk
iNk0Z2L6sq1Nycn04L4zntGC/Bte5xXjyxRrk/FjPVVkFuVOWRBGJ19h5d5RmTPph6Tzcvmw0Xbt
e4pBcyzsdN80a/gRxUTrP9TjOeSl9rbWStUPqh2BMQWqDyNgUhCj4qNSsF1Md7EMBv2x8QKCM/Fz
w+20X3DCVsEq5qwkmudwPg9ANnHU3n+YtvDjIRJBVnFpUAxr0foyCnxDZ1moUqjx27oK8HqqXgtL
UVmCow8NYsCQ70r9wZpt6dglOSS6nomSDTw2mJDY0nWhZgkQzocnDDnNVf3DR+OL/7SX8jRgglVi
WRqazu/GdcN+5fDEXydb4EzzfPGZIKiTXMmlsrTObeHYTQB7gZera7uYPEGgkFll3qRS1yNWwx0b
yH++2l8s/P8w1DA3XwRi9hlNZZvrMFLEc+IEVLDfY25KMbpthRcjQcaOqL5EHtztJhGRrINLPDdr
KFIbcHulTpha2B0vDRyV5KK2NY18qA6HCSlb0fQiSSocOTS3wrOhp9V2cKIX1WteaoKEpSCHz6Sz
qXffnGbdbXKuFEVihbJnpSZisHcdt5bVvp/ZVK23j75oDrek4mih/vnQnU330gJCFtWZ9k66+zrq
6vUuYBJsspXW8im6pV9fd2ymGLE5KBe1+bVdmC+c8XWl+SkmFp0pLybPt9NPyga9iHXJDC4601UF
WM1/utSz7eAYplhQH3wcg+3Aa7516BG8if4EGDkxgiY4Gn2DPAPC7q1LS1ya8qK+KikaVLUA3y1a
2V6bjEtkUARIH2xlZmWDAjU5BzDLMe1nkMNCtZ/71jYIHGlGPc75NwujcS58bMNon22XvHpZcbhx
oGH1pUeEOxWRMPLFe9z0yYnIzjytQTiqwzPtbEPrgw95xMhZynB2BkD2Cz6xYyKgCL0vVoxgVWNo
blV9WjXPjOXi0DqLBMqnHuqTRijgXd7NUfjwIxcpRvGjJNGAPH5Q1B7dcP5XJGX76mD6nR1DQPc7
QPOtvV84J+Ya/Po4WAb3iWRW3kubNm8sT00L1JUf41KSOde/BcPOx1Bzy9kfKvt5u5UZezuTTNOw
wsP986jf9dZ/IRgJoHA5AD4nzF/pkfX4RTmZRjMYzNgNc8hcCJ2nqw6AhwK9Jb/dVHHFUXKGC9Hy
63ehANhXtTewHNZdCFjrd9O2mD6aY4g7Vo0KA2j84HoSTytyYca2h3G6ck1TYOSWlYWzY1cV1aP2
bdjiGjxjvL1VzjkhxTw37QI3C4mhy+JsqKV69kPjze9MvKV3aK3HI3V2n3OTPWn+iQf8MXOGgI7C
3Krftc8ZbjhPcR6krC7V6/EjUGj0zCuySDEu8VdJHIc2Bu+VHazsGYHGpX+fOY7evV6RPQcq3DpY
yTUQL6RPS2gIR3DAIhYJAXP5BBZqvc1RxumgqP/GHH8A18ZPAbium5rFRh1eD3YolWSifw5CZlgh
pCjpAyZxpgbYyuq9r2t5j1N6OW9wCIdJ4Z15ezkofT9e+gIzcIKssS8S8N/N861UBnK3U/UvPQbO
Zd4qbfVPaCfFd/G+XauU2xYs2vc6eWkchYM8D9V8G0e59ZsMif1aD6XPVS/AFbkZ262f2fxfAV6X
eFp5UZZqOJYrodVepWF/adkD7HayzRfvEoeGUelXB90M0FGRdVk58JUrq0egOre/FtyVElnp3oPC
0+I73pmBOt/22GWxhQBoCDvbyQi7NB2Bh6ihwC3Mglp01813nVZpT8ddMN6Xq6gpR7jvDCjwNtcF
OJqfj9NyHPzX3J2IFPJPURIOCM7lr+l1ZQaXdYSppHO0WDMjXeI4bUB1nnFvC3TPVumfAqjvd8P/
HhGglifZ4ed/OtCGRAH7w3iagROE+9kvxwttHCDhhiDSoXabCw9clvWK+esc/CeP/EVs7tgIkrsz
/EPfsLoQbz3xILdiLVzhWRBqPqnofNGyYUlwcoKsW9MPHujORjH6k7Z3EkKnJWCSNBfL8/B08/vh
dstPFnIB80ifdTUtyFBF6ke3nShfAF1CVd+rK2KLbZ3PMMFMbSE28V1OO5fN7IUCuMRGVTv5k+p7
CMi3dvFrSq1pjpAhfgTBQdVSdXnZfiweh/Sq2peZ1POwWzDL80VdGmwnn6O1XUORWZw1xlT/UYUq
2cqUYWXJBbwKK6vcHpAn4TQySXTit+ahArHk9De5olM7NEBIou/oHQJHAytZ3eXt3m7K3assqrjh
qZqThdkwpYTMKLSwBMyZEHGcKS1e/uZLrL2xmYkVzp/k1VZCkPW47fOg7IcpLYZiOMJFiedS387E
yQcEd+UIbH19UaHYvFfKU9JM5+llnRNyyZpMqtMOW8zKRDrYJHZf3FYNUVBOcoeZk7vSRgv1aBJH
vFpdRMaeSFPZhEJPdkxj4wvzsiPEJxU0j+uWMIHujD7460ie/ALNVBeHi8vdPAwveYo6xH6Aipg9
GuDgqR3RUobZchp/QzhNbWnfHrdQGc+IpgcGpd5o38dKCk04tAUv3Kd+jyG9Ac+33wcjgSaMvg6m
5aZF216/33vXmcsdeVW5W50jDhUBuEwGivWusrLOI3yMrhFsdzPpx7LNArB2I+biYknPdngoHXF0
oFaW53EwHEsNciBjcwcb33p0Z9xuMOBvsIj3WneA1PMJW3n/E0BGYchFqQALusg/p562xbguHmI0
B/wL0yns1H7xxYi1W1015BhhJ2nCoyH2U2VjXuzXn1Zycg2pyYWgIE8mdptjGk09gGh4xbM2R8Eg
Ditxvt8pA5fUrjjPnoZOD/X2xhcCuRBry5ejAQohcwCkxgBdTQHAoGWL2HfCVdCq50gq832ct07P
WnWgp7Ftky9mUX3JlWuE5Vlxw7KGCxc97UkMzcxyQmcYUvfuaw6Us1qUXHhsO6FgoRJqpRiHTfp0
SRGuRJ7p5vMXX3oirN16RaH+T8/y3VvT2Pi83UEnUyqd0rBhsdf4cRkn9n4FN4idyHKlUSp5R+p2
rYNLDndUxrV7s6MK52W72kOiuvhzOvYeQJpm5+OyKEGh32SHetl6/ENeM0BKTXv3MIPmNPobyap3
mRukjpYjwauQJtMp6qV0FFC3YZWm/UzARkwKnI79WGs+aveF4OCOZ6QTM4jIM+CdWQpraDLUkKEI
log9pslbJtCh3KnGgLYN2cBbBXcHyNK3XjPqdiKi9BXGajsydzyojeAeNqAtUQDLnvQJwh/Z+xgE
KvGsQ9RtQmN/hAMNzXSH48zuMnwr6vt5KxnqS+86SWRJyX39FHIbja+Em4CaeoFNQWdN4v/v0LZO
4O57Sb1cZUzXNJ75yNn8PJSHmuRVerzFw9iGAGDBrdA3kULck1zqJ0RkyZMm7/FpLABngcO5eG/V
WDq2SZxxc52n3LWYAuDtE6ijcxAKpZzD7xnWUPUReSbGVe4lYl1tmH61mVK5bhQ4GpU1hZOtQ2Hu
bgixvuQ7hpGtt0I6XIpamD9pLoogrAQPKrMmd25a+RkxjO8IEdcSIx463FBzJ/OknYkALwiRsmCT
t7GnABF7u00ZZ9TkX7LFTkFlD1Rm/DW4DDQiuCrUx327LduhJnwvVW/8LFLsWNl/D7nlnwLEOmuM
2DBOmI5RfIDIUlBy/PohzjEcHPJVUbze7Ai3nh6L8OKczynhwrjzeuukuI5gaa4EYHjUQW7EdZfn
X1qJpn60J2KOLbhKfT4Cint3VCqbIRdZEtG7eOc/u/5mzvKKHYEtQ0AFSj7Aj1abWI7quMzAr94c
EkPlqzEF6lijgw42xRSddjgwInHapqkk0Ta+JAbazFvCVCtRD6utvM50aXLBB+83dMXLPvOPhn+8
6eD7Egj6JqyQFu+mkc49Gsj+T7LUfasvS1WB9cnDr27sgKnNceeB0YfEro6GdbE41xzJmZACoq2J
t8/kj23t+H+HdmXuFYGdeEWmPm92ocfFJE4gPCgjTi2TQhHqtpN/pPpDMK5zLo7zVaQXblYKxic5
NMykFu3LQgz63X8ieXQhnEle3FEyBHVsVrX2uWK/PPQ2qQGHGfBQJTExumF0KUtMEme/MUhuibi4
rAJz+ngOyWJM77i7CYQC2mtMNWWGhhEeSHVS6ciobM0o6i7//dNzzmABdwX81I6SsmIc+uymktw+
HoXrZ42zClRBMBXCKQVLKLvazDVAdO6fHOAs/ucJ6zWvUlqYVLi8gqrzr9VU6tIp/XKORsPZJTdn
gj3073M59WbSeWy/1gVgxN6aomnr5MQ4ynviEqgmpHUxF8OX+t2qb6qccdhSxsadMNw/E06zEHH/
e8h2/CPpaMbI8dEGuFkDD3n1LR5hc3qJN2CjyhFtrsZTmUEEXQCrbEMGUq/XAaguPItF4r+i+7bb
gbRD6Z9IWiKR8/pNVi/VzOlgvZ7b1foGQAFmS5R7XJDcaqtY4v1XnHamdxydIqIDgztjn+EIQbp8
3d/c+t3G9J2KuRK3PMcZvWND6O1AdZ6UapbZol+H6caZup0Nkah7zhux0RI90omYJAu4xoq1aIDh
UYqGqPE5qgmY4xcXmC/9Z3ni5IQoG02fDS3sLlWn5gqGd5bqtPaHQ+jcKmYRyJZ0kdTtR7RVCOLQ
Og9ys55MQFdW7U6osTcGcqfS/c0V9/bte1dcIi7TQNNwUD3SGrkwAMj9EpWLlirpb+HwTmAM5Dnt
/iT6x3175/So/2X5VvKF9sromEoOI0yjU0eNIJWC9aKxDeiKcrBxSRUTZiwkOh18eOLbH5VIobdS
rN9Y1D6xP6JhgMeZwb8IuaY8mYlxqbUj8t5ToQnYw4ZAVZ9u+kWUS6qomip0UPH6TdT4ALqrVgpH
R9iPffDYsGbqJtnfVTmXDoV2V2jebRKQzlD2AlF5ujEHC4HN0f1is4tJDnucx4SRRJCoijQ7JvDX
4+LEu6YmRRGR3qQGLCekG9inOst6XAYcKspJ7ZcRi+mQD08NhF3w36icRrcc6v76U5xbTKJd/OKP
IKfNYz8bn/X2RTkuB20hn2i4APG2buR4I0KyOkIjaijPQwBHUKhLj4jUD3/3TEFF94vPotWqjDjg
xmGLOYe0hFx24vTHKAVYVcsjGvVdFg5+EehbqVQEse/p6qn3lMotTBFyt3MKAl9dJjaf2BUIFAcY
gJhSI0TLeQfcHI7pykyvifJdk+t6wduGJgYxrxJlwbM45W8pnt40/CIpsL2BwcpExfe5YHUELRcU
qR1EcZ+6GVAT8DClyGlEt2keyRZ/oUCajikn0N/2P2bRW1yT8vFEdZmakNE2Tja+aJt9nO2E69dq
3Y9eM93Yru5DKScRBeLhOsSWuvzZ1gEpQRS6CIBzhzPlo/PMRDJrCtJg188WL9WM+ikNUZs72679
7YcI24FrTaCNmnKdvNaHivWC0OzMx6xxwNEfgMyqX/PqYju41D9S2rodpolmc+5bXzKcXmdyDEsC
95hL/Bl8X31ygOkHP9OE0wbIjw9eM5H8unUSgr0/4+jOdJGhf76PZYBhyp8slA4qG/hBjoDQcRix
FmdVDcULrxPX1D1hpqIfvOpkOOSSzWpxxxpE2b6Czr1M4Ju6rlQkewV5ZyLThzvfuAsg3yRWZyoS
loeqWiT2CDF9eYolD/VbE3zSiCSfviI7t1WQ6vISpgXVSMOd/L8GtOkL+8pwjiczPpwNJb+B8sX5
D4RacG1iL3N8w0CL439S09BtqcP8SNYLs/W4MIzjZN3FvhCaeP0Zg0NWYcAX8qDWRnkKpfWFmLLP
XzTo5rfrdnuiYXiQYXv5SlrfVREjiaAbneYc2YXmYKA+IpDKVTWgjELLodK8PLA37qFLI2cvWteC
rfADYcSETZaNq+oWSNnctwj1WCRI6CjqO+mhklgF0ygx1gKpTbSTGzejrpY1IcHFqtrm4O0zp0Bu
lpXI0z2mtZglQ8uHQhCaE4SYPMu1sGgC4NL27zKQ9WEHiieoGm+tOfQgYfgN8yTYUAHkId7ip001
5gDGz27lKQyc4neCxXT4Z1B8Y6XrVQWJLBcYc55QojXY3/DBGMV9T/0hY0niFYTbyROlXKTVcNod
GzywG30Y2gxeiOvK2U6zSnFhEphISEi0cVvRQzcqifXQT/s5VQi66GeEghOce5YyZkCL49Vd/jEm
nZ2JsXDzwxDfqawOg3LDgtQaBGcjr3+8IP/R9S4HPRy7aZfxt6Q0JAz/9ZNk/uE1+5RL+IkXNKZJ
szW0S+qx+Hw5KvGckaNkk3USGHhurUDxSYYNdR99j4ymv5986IP2JiDUIDxGYs2reBbDXE/OEuYY
x5lZKxin0ynt66WN7RNbVUPCrv2FnLlki1aP8J+QcZG98rQynYA1ryEQM/CB/nMBL3x0cu2Ncwpn
RnuZA7QCXyCejlrlpI1t02x6l8OUY/S72WkT5qwSoo0zfnQl3Of69yVWVAITVlHf+bmqaNE0ZMnE
7/8SSyP8Dwsur2KbhmsZwS2xmzL4iiwdDqvfzhuh2c7p+e6K56YycbJMdES5/zREYI9+q1PNKNmB
AiLRP3jU34jwHOAlajCgQaK5yYDXrhqjBBC5lNRCnVSSMCHlC5960QvrucIKPSFl2Y+jnrYazg7U
L/vabXwR45HrtT0bqvgjJX3SOPMJ/zEgsSOi1c7F0SKhOMtZWm10Gn9h1gIHwsFUNmfwOswBTWWc
9ouUMJFkZoHqoS3Y+HDSzEsxp9M8AEoQWtoCTpdl6d4xMxsd4cHWYrfOcNzoPZjmj252rz1Gna/P
WVk1/bao3edjsevGVz6HoT7vib4518wjN9L+KGMz/RksYTa7y0BKM2699YX4HClBASJU5mH+cKeL
NtTQaXTrLMUfSYp/h6e/MUfwhKQ1ecdQhFKfDlNv96cLZtmJaVRkPKTwnWB1tdfhwxa0FSU6LP7b
lVT5Hxu4B6SdOFjZ1u7k8qvOlSf/IB60oEqWNpd4OlVXb9gu1eweA6ce6bclV8UmangfkINQfgA2
b3mHXrVxgA22IDme0oIqqDPwMKJpCwZxcDAy1skZkgvyLfb12iHYtjKxxeJ1L3GMkhZjTIpCpVKB
qGhrZdeQbQupXS7djwfLn7pTLlpf4/cU+ZYisQOpEGoPEqvoKAxc5HolPRTjecp85Ov9ayfRQ3uV
N3l9sIAikU7eXsu4NH7jxaecApbrbAXTUbxCSF3S6GrXHlxpLkEYladXCeg+TwuOFE8HhbMvRpTu
1Oyi1SFjoFdJFY5ZbtKqbAvyUShrL4AyqSNT/VjlL4/PtGbFFFzGJO3zKmjRGubs5pKzawT2P2PJ
EtTiHCOJ2JXS+aNAY/x2Ji1x5/wbs5w1kvkAMRdc7YI2qBJlmVy7q1ChkmVvlFWgZS1wCutLWalJ
1NQPOhgBVlCkMNCiIq/MbCKXCX4gNGq4HETB+vSheuiL56xuSjauTVbejgVOzxBkZ/hmY/hLlKce
oZ5j3t7tmKZWTDd8p4O+GgcsALwhiQWhnY/Q9e3F52R3f2J7WjA1muwfiJMLicRbqZJRBmNjdXqj
rwdv/CF+7ODABcxj1VZtq/NL7thWKIExNw9nL0UTI8J89txn1OS3rZOcJwh09O0UXtafsTKMDy4/
royAX1RrRhbY+mznC5NGlv2uCIZnVtdD/kfkzhCre7MXn2rtpw9JLYmj5K3ySgeSo35p/UqcS7Pr
kl4AWZOzvdkvg85n/RIMpw6h8C0PRCa26+lTjC1rBosHHhJiEG+tPo5Hlzy+LHpVZ1b/Ijwuernv
2s4dCZ821ttO4H627hzBzUbgP6S5DPnB7/CR79QPh87KLE76SnY+RBVTa1NWvZ6QlqtE1L7WA+Sh
X4XTayORGHq2ny7BUh0XFq87JQd44yU6EAgaRek3MMlcxd4AT8aweNyoERitQ9Ab04FAYBoBJ2vi
/GNXvSwKlwjvrSdi/kRNd2U6PhlHv24hixAKarlLotPFczEpNANCm9o4V/Jpm9+Q7HVzWoY1S5lo
6V+Ns3t0pVkxYXlMMb1RLW4uUZpPc6e5XVbGX13UQkrBfITMd5M+jWoRUdKyUDt0j+ryVotwf0fQ
40K+0RUSLHUtK5tJX3FDZAbbkogD/E6xSEDdzorMhdTiFHQePlId8DyWtwzx9XZPo9us18+23iQ2
JcsURxiaX1Yhvkoj29KaI+0R28CRx8akQ/BpFXjYsOBDU/xCf25j5dWGb9nzAgId2ccljlakYtTl
ezQUo3U0B18mgwkbRfHpKU8+sWWL8wb8nqM62/wtOn2MTwkqQJQ8xVd4A/dILm09/VqgvBc3lIQO
E9wUZE2M0enuTD7QNTs9TceYXNnb7h4v0dxIZu74r2iv6JxucsT2xdcGqEaD7it2qCLNT3m7tB/T
Jb9+kuydt6YbdnlX8dORKSydSi64v9oJMeA6h+MmOSEZPzA/M8SfyTyY0UM9FVvUEJmh6MMF9EMk
/xn9GSkkfRgJPxlWbWh7c7dsY7iDNstghL+g7Qz/yis1gin7lylqwNbQRwHLh/stwHselIkfxI47
iXqJxpIvwjYHKyfVI/NzRAjBBjIomQtM5jifXZpaleJj7YCMgUpYjEQEENPZ+ZZ/4uM2BrQRPqTT
rJ4WvcKQyexD1ZvNCeZ6LAK29xp1egFlKVpyqdssMFnT8oAtN2llhZDHNpvIXBVmwLSOZLor+pJb
2R/kBzvCQFXeGcdokfkMqLeio/pdVUdoHJi6crgdS+r43QZJDrlRq493ugOXocPtUaRk6u5fkbOM
6hG3W03s/8ihxQ9bUebJSPdbbY5KMzuMfSLeuwmyRVZfmxJY5d9EDDNZd363hvD/uV+rmyP8vUn8
AK2w0X4rgf+ydMakH8B5rynvW2VqJyuLH22L+6L3KEYDuvvLw98tNadjw3L1+1c9PbJqK0eSyVq+
kCQfCbC8BVrKwr1tvAvkLMdfQxjPPDWbuvxWdUdZ5/X9MjHXrgjOib3H+tubSuv96IqzlD+GKibg
NLPku2ymOGZUsOWTZIeOucFzLMxwSqfvfvGyrjcAVrACNfCzAAb5diys68RjIlIZn3VymoS3jbvQ
PNAEeVWWHNLN3XmipFEjTxUnRkgJg+h1iMFGjJzuh5V08vs6MLLfTlPc2lzEMAWhtbgiX2FtbYLt
S7X9y28Gpem/e3imCIMmcmBoOK5nR7Bo7RNBYdyN6jG+ZdbFidzd5bekBSOSMaVesrfoAkKh0OzP
e+mhxXWt+I++5tlLR2LSnAKfZwhPNYMkWJDY4u0PqkWCNoJI5REq9o9hfmRyo3Rf+8dkuoLFGt5+
EfkE/PwymSN9f5GLKJ+gNUW8L6//bFhlLmllq0zoWG45vJ+P4bx2qz3oeBz9Ua8hp9lmE3Dc60sL
KGsC7HuwfKTeDIju1JCtEFS9ihP8Qb4GVkJ4mWUKn8TeESbluTUyjztpmqvPK/kwq85jPsAICMUu
aRxr8KIFTl3bKeEW7d8N8icXja9iFZVa8oaeZxTqzSRZ6fEX4sH5nZRh2K+5P3iL+E6zIr75ASTn
1yxuLSz7T4/hi30KkCRq6pkyB8lBSm8Fpvt08PuvglTyOoyFX5xwgl4vGFDUm8RHvq6yKxGRNZZE
JOg/tLyUAKibVqaf6t2vZjUpYmBWWpXuyF5DaAfS4IYWUz5bIetegS7Ssw33GTamPT55lDMUqOHI
1qRm/T+j9smc+VrlqzF8++ccIx3oMuv5j4jnx/dCRACHzsjjzxfVIT9Ljcmfxci4YM8XsnCws8oU
S/KsjtES7QHn81WYRhKqkdSP4cKCFgO3mXeJd3uqyUhiItgu3DKJx0DmF5zFnzaqVOaCMdKljqXD
pSjB/EbQve3Mixl0SLd5PnD046Jn/+s+EExfQdUHcC/dDSQC2NZvprh8SbGpPVV8PaQJiFWGwwZi
eV2i9/tPMD7s1bjLyNRZ7PX5WVAeMB9nGHUfahOSf8nCAgPV9ljkqdyJvGbE/9S82ozqjxroPofk
GpHr5T+Pkuhk7alr8Tsl3gY9OL+8rg1zLMCvOotc8853EfZkaaJekm50jQTqb16PNdTt+Cz214cZ
GXeeGw7nzQfegOorTHZr63f6c8y2YopGwtfWUcvuHZyQudVoFTupBl/SA+GI6jZ6oJZnnNC3L2Ys
zAJrY0OJ1opF3OKG4G05iUwwMs6qprFnmeDBTA/kXNWz5xyGx6lwigE4KTJeKyNupVXkdkjm7RIx
ftIOO4YAEgH8AZwikZGZSFtuPBj1Ye+e67oh/RpWinuu9JWwfbiy9ZUiuQONOfQpvg9E+liqsmrm
9io0aIf6SMDtA9pntox9B+pmcJ/7CMHt6UUPV1Ekh5sAYEMlcqjuUrNL+2ze1pGPF0bGcqWRHiLA
5paa5uPfiBnbC2sly5uSIC3UqhEYSu5dO32FwazT/PVrHQW2y4xr847R2ASBg2BwiVW/0QCGjXpk
aUZG+4++TtHLpYV5u7aP0lIYzrG6ON6ZuqQdv9reN6Ungp34r9kruk51HPvR7DkvnAK9ptBCe4Zu
lInbaAxeKYc3cDK7xHq0pRXanoU2WDRcMM3jNr1mHAX5DfF659rI5RgrS3YXOtYBU/omFSP6zh77
aUAA75OPZQOv3GQeRa2jP2X+Q+JYjfFf/F0DLn7OmoyC1AydNLLvNczXEChnGaPba6CiXhEJFryX
k7FK1oYkRdWYSgComYnjHk6vykdVOzUhB10ySQzLGGAg8O0iEo8tYZQ/rBjtk6/289FNDh3FGPDW
pmE3InPepkud2Coceau+LQEoYZOFhs9zvJvnqpqwjNQDVYzr9u1HnXrUoVpCLbJ+WcfQETcmfivk
yqsGWkXY0JCfJh7YEJqegwFUeQdFFoxGWEnd4Tq4XlGSIhSLoux6wxu9Fg8NKGkwTH/Bo4ZrLBMm
Ol2mhDNgLimJ93jZDxojhC7u2l9ggs3nR4FjcbzFkmnW7gCvEYtJUtpcsLgLfipTZC+Vmfcdd8rN
ow9NEwreUzhqn+4y4afbwsv2nSShfoPocwmcGohLv+5NM9HbZjJY9HrMZwxzheFoFer29WmFU4SN
hpOvZLQmfl2aViRvMSva6JDburlFQzvzXeUpYB1X7VHBI/T/rc+p5oep4v6C6zyhVH8bh/2VrRKg
JuQnDfugc02icvdgW5yKZOSCPSrk+pUJaMMAVhdsR3GKFHxFq1U4eb13hQxNEkRiXLO6N8naf9ih
XwWUEuPdrCXlRtDiYNKOy/qvIg1fBDswcCoPB8emBBWRxT79tZimw6L9jZ2sJAVMcMd9EzqHYuYa
vx4LScuUz4Z9lcswDmiu4xOaGzH/IUGO7iM4IC9m4cB2Hg+iEljJoB/fj1YacVIuSq4I1Bd4oK4P
MEs1xOViO33kdQedKmYOD+ffBOwretJV7Jtu/qBAiKeRD8J0G0JXcjTH2aG7L0QW5ZKKHHaE/Xa7
IDLlMidooGBtpt4r6aNwbxw5YecI8SqTENky7bjbxUUW4mU9zt6ACOQCMU47ThQMh9pmxwTW3MPw
mevrffZ9Km5zACb/Hi+7mdX4JaZhZeXkQVwDJuHv9RSYbzcl69gWLTArvCQbnejVT84lJPOn1t8h
36LsOFfxxSQYErr0C+yHHObvgxYmpIBAm4Zb/e/mCNrqXh0KRZZBDgvOxbidtzaHjylVpx12xeKg
zgR/FLZbqyHt1whA/Ekm1VSJbudy/yioS2PwJRFSoQD7YiuOiBLeyiFSYja6iswlAIuc56bJEAB1
cTgX232XALVmgPy6kL0WWCy55EOOa+QrhqsDepaUTDz0yH+xcGdrKS8IVZ2NAnZOw0/WAl0wCdo2
G91r35ofvx2soUiQxjYu2QjztyfvWR517tvnIL9bUTlEsXUML15DOPTfe/xXIcxou6BTD8/xs1im
ZMduPvjB32AFWDueApiqOTPo9+J/KkL/2+EkcFBdIf9Bx0s4A+/fYGZSekY5OV/LAmVohjoJH9nX
TmtNv2ifFWXrI2k/pBDO4fj2mVT0u3v/H/c/nLY+iOvbyKHhyJpit+8wZmPZzZK6HNCREbkF8teK
+dB9dvqjZ/mI69w3rAwEVMag8aCevq42OoVOILfQH2S9PxqWfBblYHHF/Zgc0vJeT7Fq0PRhbw9L
LhUPkjAmLIk0/ZDoDLfxGWkPx283UsWZSlnCSLiB96HmJV4xlbndfeJ6RT6HOyCcBFkHRxhRNa8x
Q2HcehBnlF8uJ8//6SaQ2P9wqtCOiAkz9sEarkHrCJr4mTuphc/2sDh3mO5OttR0lFBVziM1rvxW
T9vhaQOF4RBYAPr7bi0SJzdR3cQHKIHdf/w9YIFEJfSf2w9NauN6oxe4XwseIWOs/B3Os+rwSX05
KvzaA6qbVFxTzpMjwlJcP/BC5BszQTbeaJQvEp+JuQQ0EpBFZpxvAy5wfoK10WpZom9T4RrrTW/C
ZIlk0mckip1/u1wppwgEWrlVMtoQkAw0eKaGzSL0dR/G3szjkNofzpycqtNncbmUm+x/nAJFT3ja
g8uNHN4Cd9qKjCZoAZOj1oStAW78WYs8Imm2Y/zOVf8XD/2X9eBPYy9l1LSv2IZz/zkXpInrvq6N
Bp+KYu18jrF67C9kb/ODgWjfA/TdgUPabY3CIO5spaIrWypZX6no+08jgWYBVy+IMvXAISFNeXrN
w+OxvpqSXDpe6mOXiRAGFdV3Xu5uSEk1XUQwfx204Sds+GmvYzwtnOX69X2w53wULtMd72zLyN6s
932IIyUYVi1EGJTVKI0c6tIObNWbmxn5nDz4LsHWMJlop5S2fAlw+GvyUpFBg+LKHhyWN8l64dIP
lT9RdLEUMHj7SdDLnxnbhN1vJ/DmjOETEtR273Z5b2hRHegtLNrW8aunUfM7rovSc99HK8QX561/
b0JLcCmdPcbuVSB3Yf2sREmMs+tIQ00G1tCeK4e2laGgdOPNWldxcRHhYmYBcb09Rz17CfRsZ38e
4UkqlZ+w0IvDQYK+6tHaO5ieXcmaJi1s+/Stesd4wOw64cD7mLC4RnNv+jwSZmNbnA0J2ePRhjrF
LXL+ECDDtDAJFWLdgpEpepHdHUMzqBjULOKlokw6BBqb1T9wzGVFRTWuojuBhUOhNMxaCYuRPdiR
VtfEouVmlRMxt2RHyGje/hyuIE9Eg1rs0yOEiqw1gDeOzOgFaun+Jp16NiajjLFxZ8fNXZBhZJ8o
p9cLx5CUzpnczyogL64JPtq67JPZhMJp4RKcrR0AwTPaBRCCNkTDbSnJNwcojdLO7bueKm0mVntq
53q1fW9IIvJkdYj+YykTnnd6db7xxy/KdFkeDbly48Ng6nDp+swJOsqzQEsWZUTOfIWldWVZQCX4
Qr41dFTRwQkUbJ6yvmrVqwKvTu0d25DKFCiJnQaiBStWJDQpCn4LObH9duudB9UlahIv+3pqR9sE
w93Q3qw1X2hfa+pgmok4tVb592a99nPy8BYkt/gFNxmARgffCfHBA4/+Pivo9VQ73JR3Ks4W/pmC
V/xq9Eh1NXD6IzYCWSqn3vOBYI1fvoLpvtRpRZ76TqdG5xH3VLsehaNYAj8DICpRJ6fKchFSoxTk
u5Is8dnRtl4SLhlg2Dfoh/RamtpvLhS0ZNV6TfzQ/A0ZmPYs8jjoN9TQcKURm92XrWuzee0H75JI
Rv6qq0qMHFws2/A6FNbMxBbmJgngOMLpnLa9w1/EEvTxIQlAbim/ri6QqV2eRf2tZLNRKy5j0MVW
eKy8G4P27OX+KniAvEw+KFPZrGLJSTkTHiuLell0L8DGI5WetFn+PLQCfbpu3BPg45Nqd2aBBzSc
FcgavsbhLENgUfn5oFQWTcVijr1ox2C9Ow5Tm3rWbI15k9XOmdjTTPCZWZXQnwUZD9mTkRvBZdAx
xR6yHyUznsASMGrRa/XeGV1ZoAprHrxlso8IaeI/NyqdJ81qwEcHzes36DBwL5D0M0hNHgvMwvzb
qo5UmAUwnLxG8ImGgieIuHWfGuViXNY+/JHvx8w1QnoRzfau7EKJcaUPof+R48zwFdDmMesgOw6v
EV9p733/nLtl9pmEkfXSYXAs5mGPXouZFYpzWtzf+QtzltGz+5hLpfXk8JmE5QS1+00DEyPx8jnX
2FVrH3nqOHwn7GMJjxUMwpbCrGP2Q3HyxZyoN3aMzvRbxdpXAVRe5rYgC9Gl4rsAug2oEcYSfeM2
Min2q/uNOD4M8s1k8qIn7Hd5QzGdgYZeTezC5DDg8TOXe5caZiTn3ErYY8cFUPmQSaMqwUltiywO
HNvZ7xnLwPyKh07bk03RiOSPN7BEjBy/fSWAmWoEEj66HCr8jydrsWReoN/VI93kTcOibcqbqg+k
GQQwd3WpDv8K/vboubIhp437D0Ve/TocpZG9lha6WytfyEHw9Kpku79NIhlP1SVOcnfm1RcghyBC
o+MZuKRR75F/uE8TBAEgTf+fwkrRveRWlzSpDrCtwEbOT5W9R4fKP6f4PuUdy4YgRKvek0VenXni
GDMH9zP1H6nY9nHogxx7t5JhaKnjTAFZuQNi9oxC/fotMkteSh1dnxebMtvOlkEY0y0hqG9q03tK
QvLsEUN+5AfHUkK8QVath2xlMt6Pz2eeMUzQ09mGJc5BbewnKEfvA4ESa73/aYsj1vWasT0q0fi7
2Qp53aQLPo5iRo+Vn/0qC6SSAcmEpAkJ3cLaytxruTDlzNsir+Y+s9SUvtF/9ZJwqhntMdk1qVbw
P3ANRBD9yGj9JSi+E7zLvMGSxpDUyPSCY/2q+L3uq8edpYTGMQ2Ezom3jjvZBTCnPis/4F9vPs39
1+U+zebS+JVnZqN6pMu7wNUAVXMYPNf/d/x+4cP586y+Z8QJw/AJzdU6SwT721TAbvM408PwlTfo
vXaJGdICMftq1expbjNx4uFriqkuT5uIytOPYBIW0y4z0L45caVtROmYVZ+J9CW0HGTu1DXqsKz+
nunugU2RYrIRSE7NhBkmSWK3kC1s5/hR+5MO9rxqgL2UvTuYfUqyNb8qMOpR6k6H3DxhFuPeDr9v
YTCc5dD2wIN2Nyorp331vr4CejvJ5EER7SAmYKLARlhNQumhD/RWGXGtXyCly2wHGkgVtkRXCgvM
OTikSZHjHmlOdney+xX9FnJAC7kEJl4q5r65joTn+R5V6p2wtdQNwYv+whGC+dVTbb8v5wYlZjiF
Wt3QDsgmkynjYyEZLqu2GSGEz/WMs7VuA1snC46dU5Cnt9esx+6E52w8nsdQ4viBXYlRs3cxI9Uh
PGAfe4i3okLrQOvg9f9VL5xT8JpFZEuaoVqoNgSetCwGKKTgTVQW/stbRNnpK7BjdzN2lXfCFDn3
o6SqgYKB/9KwUoQycX+tI9ZRi6Zy6p+N+KtYHRJjK1GB4DsajM4CSiahBKGIgBVHYlPTP6aOmae8
9vZo4/9ZR1jyLc7SSn2Te90IPFhnhnR6rMvomq38v0GePoOgmfN0Ho/hQ47K7hLyodMzGZE5NyJF
me4XIZhf9i+EwHqjr7Sv0nHuz+PiIBNe4G8y1ePo0OqfP8FaPhl6Fl1zDrjeAWc/BsfbhtuovF68
3ERnPEU35kIQBuBMwiNGZy73RRVR1X4quYbbvGRD01LvaZXlJbUl8lw6vcwVOC+uopRiDYYUPckp
lar6SnCGED5oC7Myin1Qy56DXjYTf9EnjiAaxo2Z6douomPE0cgqMLx0g7/YOzLnAF7CRV7V93Ta
BsKy+mhqXQhAOWuERclaQTQUpQUHulJSbsgmAQwCNB1GqaaWfvhFmad5SMZUy+Oy/FeR8tOHRPlG
/wVKczyfaNBRypLhxHZfHVwTMazlPGfjt8CM8JFBf5Np84Ucy5m7LYdeaXWzs4e94e9JIwhlrErQ
1/zBxyDOlW7ejPHMPH3qdPDfKFeJ79R0mysLaTgcF1cLLxhocDv+Olkw96yRd0y66z1RcVu0YA0i
UI3czyTga6FQM8JwZlTJDnhORfNd0RDh4ZrZgMYtpOb0n0Leey8a+oorinzo3im6WjKwe+O41XB1
wJY2WxWGbWsYdKEA8Pco+5NmiOV3dhmAXnS4j93K/BKWjjlQxwLQ9FtGbJVWUZE240osyqG8dbOO
wPFwrktLJmClV8kuJTX5mPCV0Z4TXwR+JtGkLa9C5VsVFHnQb66dx+QAMEnGGmTTjtmtglJmeDIn
STpkl/ITLmtOYbZ3zofg12friWtNrttiUyvXSLGZKdCBXSQa7OibbyPiiYTGhfWgMst3Lz49B9IC
/8rtiseVVsnaq9P/V3qvi3Q/PD6hjuEQlTTxJDJw0fhpydihW6Ci76E1YTgKqeZ/kStqaLKXJrws
HYUxNfgGKmNiWgDfzHMWjKwpkeJFtowdAD1Kux8zEHHNH/mHW/SBPvZ5paMYQpVMOCB7h0olD/x1
e0DE6TAMj4GaPVMvwpW+iqcc3rBS13izpPfebda+KrbvZRkX/naJSzQTh4Dy+66tXvSN7lSAI3NL
LOOsM+7tI4VC28gUHIZ2xtmD5SHlq2k49kam3SR17ao1UWj4GuPU/qNe6Kdy4umgAZyq8UgOqihJ
MnjLqHKxHfwu6TbxVVphXT3XqdinyvJTifkDkHcSN2So7Lhppkd3hYw7NxOpeDVT7gdsPMttyUWL
eEpgWjKZAYqQ77JQR+NdTzjx72YSnNdSkj2AewSjvmUXNgrYtviXFsTVpLnCHIReB01P3cuUn+NL
fpDJtgi36DBYIT88twQOZJg6jnBkJNAD0VwVy/J20Tey42/A57q1ABG4Rk2zDPgeAnSAER8DTFMI
c/rX/jrgTqQSJJNZAWZAfw3CtWHknpwo6gq0yslPVwje2sLCIWyVjvotPRcoh8eaZgCKt05vOOfb
9x6pq8EKuNeDH87JtW3f68+7e7l9HPBHlZuEUmpvW8jBwyeVcDevk7SYvvX4VgQGGDoGG1v76C2a
4/zJI/J1jcxTj+rEolOICd5RsK/k8sMPpgbg1qzUWetaRH8+ed/bAg/TpS8WAhOITKwP1hJdtYGX
zvz6ylxuC0ATnCk7VkFUV28hDxxWK1RRRiaFnZmtII8o4WX0ZtfJIzUlv/tnklGvVQj/UPr8FDX6
gKy+eVze0BXwcQgutcISqT5M+SR6cSDS3Am/fwxYlhjcy9sMpnSJP0DARhKNMx5RvZqljEO9qKUO
Oz2s0khT7WWib5U5JuWwMyWPk1eR6Z3pPFj8cgDd1VQEMzkQ5xE/jHH5LaCR5rXX9X3RHcaI+nGn
yejVhrX54mA+q29myD+0VTBdIQ0qaGcInwnURgLsv/VECtGmsP6gG0tXbAQFa8Bt9oVW0pf9gOZr
id/ajtqNaiXoO0xl1VW3uvYg3mNZzvCSXmqR/rWlYFy/TyPQ2EkODMecu8NbFESZrffm4xZVpaBg
Iz8P09ts8Wv1AZ9IMmXfasLaUmAzY/xmHEMVFr7oscv7EPc0RY/qWuxHS0HFepAGdbHMIfGspdrL
P/2KDv6sHxgo2sjxPCi6ZZvnvAnlBvQnauGG9tN/DgRBYYtzZFk++VSOXc/tgWtHL6dGkwpFU9L1
Yq8ZHG86RrZeXRKtaOx38PQ6qeCDWeThTjx3eIT79qdBX7SYwSqD/0XxwCmRKBIo+UIGoZV7dKb0
FwnpCpFmCC13MIEUoL02grqfZ3jRJgH7RXofNAS/sTUkrwgbEgXmble8Zll+IQmwrdKAeC6VN6i8
expgVfBUGBFcekzsIsA9pHWMVE8eHF09LSLODOd7hFeK/vV1VCEIc5yeBaF4Vf42d/sZSOHP+E3o
7VCUERmzGy2IM2G6afNIF0fO2jTDu7H7hcVDBhlpRAaIcVS3UW4kRGEQggOlgC9yAU3SUX3CdSon
jvW3m6brSnz41mmRxVJyhrLl0mQKs7Woi9qTBiqL2pn1NZt4vi/+XTmZ2hnp0z0DMbmtDXk2zTh6
rKfJJm2gBa4BL0gA2thAwzzfzELlIxh6iK2bTnGFjPQRGVeh4WDaAc00SNWBu9B0Fnrw5ODtF0/t
WnLaYHlmdVhpu9oi0ikepkQg/zKUhto5g3jyXdfFXj5Giba5F8HrkeaV4oSTOapRPDdd6tkB2bQL
sy1VeL09hvBI2K6sfg1F408Y9CQuuWLZLWwjIM0AqlqP+8l957GdUcSv6m1ip1wcEuNv8XFlWMvm
Jx2wGrpy3805GYxzB0eRtwE6Kqy678zOlEV74BslShR9s0JSjWlusXzEny27ucia7OO/Ytu1cpfT
2Hua56eNpnl9PlXLkyjOn/Z1lAuhTMWCii4Mjka0apt4QO1Nx0rUpvUT6H54GUVFFCtGeaG7Om9M
o2+PJvYAr1njc6UNUTM+O1h1n0D6rWwSlXbF03rury6DGvy71QHrH6ZVxCw0FI+PckvDLAll17gw
kJ4yvWrZTJl6pFjJRQ39evXShj1d5dCTBKUs99MSABJQoQi9NjjK9rWvlkuMLb3fF2AT1LuQU9sc
ZDAgWhqM2Jj3VjTmAZByFRCxu1nx3GNlqv6/kV0MzjKMqWUahhvSzEjJOT+nxjgiJGxMk1KdyXvb
jI8th6bplFqKFR20l1vjblJhV5vYeZPWsy+YMeuSbl42hoPYjaDGdSskJ5JBgu4n7O6IKyMg42j1
pYOU4PK4FTRHkT1Oyry2XChTjDLaZkPXjhTmH8kvQRdNyUvMbMXPUBLNIBIhizmXz4/iaNxaLN9g
ksgCmS2CuC5jyyWtNwgXf9fQ5xQxVmJaTLzkBlJjafBWg4VK82EyIG4fO+R0jOtYcW91miGwnyVn
Ctgvr+nMA8INESTF4nk+nt4UNWIgj7UNzanH0Omb+KkeK243fn5M/+RneZzpmiqjh3ttUkGeBd4d
L0MOUDHoDTNorfzB+gk/zakoW4Ph8M9P2E9t2Noy2LF9ZKMg+yy36d0ssZbQHHf2KVdsscTRRgRm
ncXFwwRHjoUfCzbUz8UWFzKKmcAVNYDGu99dCZGLc0y3mXg53tYXd9j0T94G4CNH2WEyVYIGuFJs
lITfJZosyC/eZgbvN/sksHFzNU7pFgFCmTMvl0DiYBy+fJ/i10QuCtCLs4qt/j4NlP2SuvRTHmNe
GGvDmmJguMvGX5b5VD0THjVdd8yl6IPVQockXMcf+3QyPn5mHSJyQwtOITAnXfumH2kSjJUEDLyN
yeVuBDGIqxjzCJWQjyKRciO5eEpCgal8UbGXjBJpAXT3lZgVpuerBJLiz2ggxtg2mDZOM6Tj1YJ7
piDskEUz1gj4uxDn3pocznMgn4CY9I6c54ZZ1m5c0bO9FFBeOnaa9Ob18mq+Q/a/TXkLVjqO61YA
y426bMcVIcoTpQGTeDy7PKT1zy/7XB1OLMMVF6CUV/wNpuHj6lYNyh4eu6pDfFUXsWNkSBJjJs81
boKHtFasivreXcGqEy5SH8m29fryq2QSw66iXKiMx4kWPusQh8JGe8rcTgc716k85zNAurP3ERW/
G04vBTpmKFmoir7Z+TRnMe1A/Y2EKKNy602gq2WYdb38uINdOKrUYAlPMgvm9qOLks/vPz12jsoc
onhyYvfYviZiytFyovBQ72Sv5jNaUJNQwfV7aCCSCQFjlHveZE9raEzAKQBEKCnTcuLBaw/2g/G2
6DbG1KiDqSv3TFsE6YhZw8r5kYvH9F+nZUesxoi9g6zIX+Yd4GxYw/It9eKX4lpXH6hTzRZtK2tn
EX2I0X+YmgGLjRwN02czfVytDAxIbpcnXxtWQCDBNDdpiXEBVOoKUJQbfnA3vHbYaPxG9ph6ruhX
/YOKakprZAKMNshfptNAOu4ursAAPLTdDib6o65wocEQ+z6EQar/4Yts1TsTgpmHJbUvi3pMz9Kb
vnKgtIc7M3VGPTWv0nHtDN8zUhF6bjTmV/BkxrgXKonQYmLxKJw+z1te26EsS/BmDek0x/ViLKfH
vxhM7gHB74ddGR78vpmuaSzPR5npC47vp/EdruFu85VzLBHwMV/mAJyqSkBzmWelpTEbnB3NYiSN
2Ho74ganD1EDzURdMca+5RaSg/c4mJQ5dbfpERI/Buo0+uhWkis4quF+ZH8cjJ1OC9r9XGpavqTz
A3y3r5ggEvBNJaZ0NDpo4v+tD0HJTT2iroSEFogViYWgZ6sdbFUr0Ka2ogXu0MpapCUPQqjFBv9N
7Pcu8C54650taC6Bs3i1+nqEIrRJr24kENnwuUUizxRZraV+5vm4+APCenHcc0DxrU+ucV8/rZSt
KDBeI2hstzfSsqWxWR9FI/qicgZpSbeJ6tdp0gXy56xBEmLjsi4YNmNVtCt8NaYDoU5jyf/rI7ZD
PFqquSNq0Acq5fZz/9eVS5UicLeYNdDLW+A46asHvnaJF+SAqY9viWDO4M70VGETheQxGay+3jNy
hzeX8HVYnVnQIUPyh4NpHQoD6USk3JSL2Sbx+c4cL+xTkrYi6g39aWF3MApu/uITHKJEtzGjagTq
l3iBSLvc3I7BpW5ViiPK/TuQk+SeX5mVqD30anjPmJH0cwbsUjn7GDy4pLI/MjZhs7S5BYBUnqoi
NKaTcSNJeznP6mEfU3AA1mntcIUmC8W6OdeCUC69WJ/6V4wvfxwX5J02K7qwmVo4ZWWVWwGgsfQf
np6r+CHdBZtJwkr2L1KKfCzzcLV6wUV4dI/w67HBRVTDmFNfiW1GjaGnPqMQqvdV+37JGJwd6c9c
vy9QVq9IRNaV8fYrv8PbuXBaqua5MEmgEa5m6EziihWMrHoZzpXmPqfCfDN/LdJxAevTiMPZDfpt
capaHojmRTLLmvBAFGmeENobgdTZuHfCMFRXm14yUKoOkpWnDzbmQ/vnboLS3UzfP87f4uK4AQi/
zHPZT6gFZF26yZ2jZTVVQarPHhsbZ1BsBkL0n29iASczcLhKR7QZrVgm5oriLkqW4/pYhIoSLQBD
LDafVt0nA71qoRaEEbAMsVDLD2bqCiMSF0jsbkzIRno3uavvPuOX8fzZDsSW+4SOX+hESd+PqX7z
ZR0qIOcOU5qjC3HFl+Wog9oAxCM3GElBgq9LkYKtaLcTNVGp1QPrzr1R+rCgeKE9VDg7evkCUKss
e5fLNdwz7vjIufQ9uSPlmPSMaJX3516ayZ34yABpRTx+dwZm7f3c5sHFqUXz6WwM2u58IrZPfYoH
v3SiFOLaOBpYGd7onWMEzNanUyYkJYPqJYT5lXTSXZMwd5v9M78BGVOJGR9d9+jA/uw0ep0hIRob
uwefNN2VARj3L7OsXp7dClOxLtPSDe9MAqjzogEFv93qZG8bnbwnKPgAfnrIEKyQUzQpIlC4wPwK
TUz6bvIZAUDaR1dHPS9dsb6LutHPKFsUj/TDswRhGIEGv1GUJlLgEQk8uBd1B4L3C6366N4xGDWl
/R4AdxY6ZwJ2oPNg0yNwALrsevgCUIy5YhHIibpgs13inREEccEG+9dXAW8a9OPg6OjARyS5WWak
txL2NFzhSjOjlH9FKR5ecxoI7rJ2+C3hhTwMwpIA/z0sW2o/FXMQOya3K8sphEV3a3Fd4HTQfEIw
z7e9ZZVQVqEAppGo/HQTWMg+3mqufU2eOgcg4PVcQiBDKvM/4LqRvPkZphUApSLfU1MMpAMhoZxQ
RC8CBbsAa36OBl2ebk0xP3d4AI6ZRE84ye/L3ZsS2Bd80uLcFqxeXsBXrrNCeiy7MTsMy1CpzR8p
7Nx2fdv6pp4RUmW73bfaJO5jCXgVTSWVMsqcidhjdaPR13GP1JC2UcHE7sebl/uoxLNxzeQgA1KK
hwi/j39KcNj6N5nw05wXJ++BPFtq5sDq0s2IF1r3sDM0A2XabjYuLs1pBdvrWhXK2CMudxQhOMaE
PrR1av2bn43IPbUfVSSqfFcXS+hWolPOYrMdIvyerR/GYiPIyaV8DOWW2amFlBVvyC9/+Y/+jpMW
mFMyawxHyNKfhg1iIEKRmBg7oeIo9wtAYCaHuYT908IJ3rTxm1E4Omp+SZr7X+V3m8X76es46sHP
3R9dZZ0UZcun8+ii+IVJEjCJqVZhkhWTA/K5brljlHQ6n1DcyDcgySVPeoISzMn+js4N6YQOQYbU
Msb3hnSvymGlhEsRyUYDosZkQ1vlvOMW3fCh4nXHpSsgwM9fCVgL3V/I1S4w29HiNONOStI5Y2QR
gvXjkNtWrnZezmrF0cNxN+OvnqVyc4MXfOFmKSs488GQFK/2JDWKzvCj5GMrF2jZFXjNcpMN4UOy
EZpVdYfeAKqcEfaGO8lVzXoMuX2ZT4CFB3VIgbJ0BSVqFx94xKc2YuHXHopyn2mwcBp+z2N4vxaG
kD3s+kfD0pdEVqhTIaKGUClPky0iveq8ZV+vDRYRZzTXNnpJbiKgDU0AxJ1TGn7j95ASIIPGwN3y
8uEmKXlBPiM45uSmlMAR/NIC1Lle1d9rlomEebl53YwzI9Jwwcuda3x6N2lWPwbMRH/ghnjA3Xx6
Ogj3Xo6PX0uwwuA2owpbgMIOc4U6XhT1j3UmC3Kxp5ZNzFgoNzroRDTmYuxHqGI7KgWleVlesoIM
/2mCxnh88b4jSLCo8MhB+kdgR20PO/nTY5njeuA1xo4oKTeUvGZWkZ6HL18hYK+7IqTTRrVw8RbP
GtcYV/JqPBdigQotgOpGmhF2LlTfK07Edbuo3ocZYj+g9aFI6iPZeWvbUGf2RJ0VnPJwS2651PyP
14rEM3hN+JxS0FkrqYHrLR4gArgmpV/4FsqcR1HCfVvw5rKeSUYMoa8+fzD59k1DJJ6jvWLBrpJQ
yqEcD/qdakau5YN1/b+xdZzZmuW/E14zgXw9iF7JJcKnkHXGrGMmeofndWvWY5szb8FQaW6ovGZp
UIf1D9O9yKiLqkbQ+A0F4q3v1QnLrGvneu90R/T/iFTZ5gHiKaRt+eys4cCALmAYHpJuMSBcs1OM
ucpJ4ddOUBk7oul4Rrb0zjVIBaTVYbyLWmQQsVZHiok3+upB/Sh3Vmbpis1vUwD3oDRcYCNXMREE
FQfpPLoVWtpoZuTjaPTuLcsv1bpoUQbuQGHhdhiBfw5HmFioJAhtt1pObSNcYr7dAIiohv1UXm+b
eFpzMxlO923U5wBFRhC3T0YIcQYE61QQgRho8G9a10PILy+Ief8OS6nxQ/gw16hgS50OBb+kE8ln
yAqammhrUMBQSXzN6BCZPNKA/eVKHwn8MaR4L9lO09uQvFYmhxxNwv/3wI50OjLjkhJFiSHUKhQh
Hho2r5TcWU69JWTOjTqs9RXD824vIrOzt9dxmwzzZoDpPLTnFhaSp68NoBfU42Exog8N9nkw/CCN
N/euKV6+hL01xZUluufZMOoIwYhdNLiY6PlhKjUMPYTYw5r/j9UbW0eFKafs84q5+czx50x28rdV
TE3qQSobwDO1k7YqxUh+dW8WKxBI9KntAsfpJ5ihlMQw9KcPO48MS+WdYCySrH+kyVlAfOuSrgS6
MdTfUwkA3c7vmEf+mE7mW6Zkcwjwrk3JJyQpClI/OHt0YFus7EIBTd9mTAXWgv0Sh8IEn/yGz0Js
P6WxWBdKNA6iMlGUrenhfU6dr2W99BsYx82UW7rZ3Ur/GTMSdgy8DW30ZbBgOuIyIO/WWqC/LDix
jNK0cBo2c79XfQd6S/pWOxeIVGu7GyQAyuxUQG98IC9uihJ4jSg1DmqpNgyIjN+mT4kM1At4tIUi
XyMgTQrVRedkuL40XW0vZXYikyPLwziGZHH4jZAfbxJU4VfNjW/tt1tnKPohhRLH+kYAY4t59EY0
9K7SYG2wOnM0boD2eDJwu+2xua3oIWVI8XEO8tXtpIZUmWZj1UGD+wIGfmR7tAVjB3aIAWfmz3/V
0OJOl7WQM9tkri9Ti/4VFgGg4XaWZUj/2/tooXyl1uYNRaH3eBofcOdYli1cEDYDJS3eWClw5P0o
lTdZQJWz0gryIVGG9hErTBJiODuBNiK3u5I71hG00cmq/ZRtKbv/UVimCF7sS1O78NsIyW3wuuy4
gjkW2ecrV2Fki6BE7K1V6WP9YTiMqPtUoHKOguHc7vIKQKlZm7AnUsc/5FSvRi9g+xir9q9UjdAH
FnJdishc8qmNP1garAQMcrtoizv7+CFUj3H9tq6YtaPDQhhZp2T9cUnaRUyeueu0n2TsR/QEWyKH
HBryEPOiVtsdrARzv4J0U7YVo9h5D3AsaUCdl3xM0AWTIKpS5f3xaz4HX4rjf95yKh8PZL+ggJMa
Gj3zHaHvsXHIQqNjBsAO6xXsLE2UghN0lniF79LcuqmSdosocxjAi3+ARE+zyosnDbYtqd8qGNjF
V/8MwncuJSPlZ6u7Qcg+rDvlgN33jRf4X/2PD6Y2nPCCWLjKcehBTXCmIPBJYdP/JzIx9RaBPx39
bnlKMJvW6b8jeHZsLQV5W+2/3GU73sr6BsIABgTBtvyIEz+fUhDKIJjxUHTd1IxRI4VrG3MVbmEF
BlhC6pokXBle+xf+MZ+k7BGLFdVgcpqah+TRMa11i1AbgLwKCg+Rk3KJc6Hwtz3B9OAFM0gNmngb
4g5f2mguba1OAxAuSkG95XZ5Our9CullQerVNBPuMZ6HsR9WT4nuQ5kSlp+5k9SZ9e5ANgXaxgBn
UwVRu71q4QKPkCZJ99U9aVwR2zOByeIv/i3k3RY70AhJ67exmMZpWaHHVlEdtQMDZ4aYsy8Ism1A
nxaFiWIU/PhkjgcmQi+4j0f+pn+Vi9vxn3HpbjML8i6NRYrwhmfEQD7OkQ9lO3llOfBvR5xYo4rE
km4xvT6LE6Tkdiy6vmyxbWOnOOl2tZ6UBvTfu7YWH0qBP7bDLcgp6sn5PowsUk62jYqAO9DWLjO+
G/c3mr/sInhQrxZzeIfbhVLikV/8wEhqifwnVKOUTHfwQ7RcJHAafkHUGYB/XkNhISsa/9eE5WA3
iT3Qp71hKdhflroLJxjPzhxiYDqdEhsc/K1oyU+LeLC45NDsBF2vEik4WWWrqlE9l4ae/bxtSZLN
ohGKwTsxLQvZlaa2Rcr2QPJmADz25W2TCgHlbEIvrOVUo6PI9u5NwBjIohVerf2T7yFbxAbCjpqS
XnqRuovMH7v1bLDgb2tlRhkr1ZB8ePKVbm9EEPQYlZaBYTzGKna5fus0rPpN6uhk9Y0SifaGlqpi
nKSVbz75bn7/gt1jQzMyvDFSP9x4i5ftnXzn3Wqo09t0lvWP9NZpfQGG9w3rIpPOy1G+VrH+L+Sj
UaEtg9ZtT6bPvM1CwGS8sk/hLz564z4jREsq4jQG4O54Gk0SHjCFBEn5a3rrqDVrjW0CnAx6hl+O
td7qT5G6+J848tryf2x1KiUGSrnNcTGzOFXSKB7BKdoMUS5n6jnQ/JBpl0bgsQ5QW72tIlVQqDFM
lUHC8+AfAH5V4bjmqFmPn+UPFF5Hc8RxUUo7ldnfRbAmpye4LfbuKHWNiDh1cD+mjcIAQ313uiS9
Hn5LSQXqCs2yPxMPfcnn7aXtT9e9cu0CpPhZSEzJjalxwA5YKQmUrjk/1WNRA+Wjyp3FHHioHYdy
YYnhNGvr15f5wQB9nI+4ly5wM1k6dqix+WTkIjU1fnzKTm+pI5NvP0/Enx1YuAC8dL1nQUvT2Cbn
pM721s7VbukcqFkGnFRIsdYu4jZ1BJmgCCjDgBcg/OPI+/BceIivHiqceaw2Zke/wmWHt+Sur4qd
9oLo6vsh3gIdtC/GH5gflRrwWKhKDrzoaUlOs+j4l18+ZcsHf6QQasUKRvUg5yi5E4GwczpwbEf1
Un6rDPXcQI20jyzcGHjRcCsjHp6PG/lVSoHzRF4Nk7jTZj+BsEkXmyxENzM3F66RXGSNLDhOHeQR
XeAX0jsG5CT8VOdpQVs/h2kbAC2CeC7tNgdzW1sE6dqZVvdQcoodebMM4aw6ONjEpx/8rp/89rBb
8zC3EZDozkRIeUZfsS2Unx2Qe0bPrL810ndRE4HUlAbfnsDuHlAHNh8zA59/jw17bSDV5qky4kNM
kdrj96PrenUF2ECNzSXtHFXmnWUkFf+PG3zgeSvs0Lxzb/Bb4CnahyGqnWc6TEr4j23Xs+XY3PiZ
yR6201KnoOfbApyMLxXdnqmDRFBKRXtb3msSveEva/dZvgtYety2hOC1FXEU7/xuJTrggKj8Ya8n
+OOQv3fQcbmyT2ae/Njrpx39pzttfEOnuhXmWho2t/RHbNYK4I8xOvgYNr3DUPhUJOeM3iyl9OVm
9EMhBnMjBddLbtfTLScxR2+F7WxORcJ5RnV9anqo+tnTQ2oy10MJ+xLYe0c4e18S9Su9DUbBreeL
EEvhJxa9FzNR8d1c9YzSAIO4h+xvOHbcDl/+l/gCrpb+yElcMdOhu+GtIX369tMTQasMtCgAckOe
ef7aYJDkrwmVCNeJhwMtYTuJpPYxIKkbkY0YrF9GAEEOEzCaRQaPppfMk42nU+PfRmOWhYMTajQf
0Xdj5RVKyyrR0Nt6wj/z25gLJTHXJcngf9WqFnAZChdLTB0ZufK1GpQOCgEJyU0nSEdk0bNMW5hk
xCpTSKdTwFi0IjFKgseqjk5jgBVwIBKTOUB8po7XTb5W0VwOJS1j/yaO4+ucY53T6N0QCiuFqBfi
1FNpcsiWNHa8hVajqMoMLC7KenhlnDIZtDPhtPEQqijQSrdfKA9dSIVOU/JHa6jrM7q96RGpPiV7
BpAqIugXPJR+Jj1Jbh68eEYdfo0XDgE2DDD7k6eJWAor5Q1z1wYKwmK6AQOSz07agXhOIUxhncTT
T4rkEeUriGNjKPTsAj/LM88LmMY2ThzI7x3w8gHyIDn9UnBQDaLx7wGZ3qJenFt3Zj98oykcDdXH
Zric6uZttNWlI2UHqqr91mNZUzvFSfaj7pNAZtZwB5O9rXHZ92c2cxBpij/qMh96XwG8LnsXLD+5
uS+fWFu2YNtHhY+nGvUOYlqrRoEw5JU5FrNOUvunX9sBBmGoq4pzcMnb68cO42L5FsH1JONpBjum
P+AtDz14/qM4j29tBcY20mym1S5QEIV3tYBE0mfJBYnq0B6l5ckOfzpyZAhoW6TGJo1LFiBpYxSR
LhKgFYMTBpg9ssrza1VwdT9jroj0sqVRYh7+SPD+Y3CspzMyH3IJ4X/j+BU4IKsm7OSU0aKLse9N
LQ/IBSCHcMZ3OUWwU+D2ZTqFInFIgoN7UxauJn3odZr0/f1Dpo7em/7eqNGFbeAspL67Q6wg/O49
J/OyA9FpHdSANeGVLZaF6lB0dWXVIy0VALYfngoQHBUXMCOaXty3Oa++XHvSOfjnSe4x5gDD5MOv
KiNZEFeZdHlSZ8Qy1/SrC8vBrqaarAJZRStUiWNHIsh0eslMHzAa6cWiLjEsV0xCynq9IDFbttr1
FTDLatDgBMw7kxr6t3bennpJOwJNjr3wljA+6+WkFEx1qZX3SLbNM89hHGGr64nZPVcnqUSTQ5ct
YwUj2Y5kJftiOrOqbALcQ3gf7YX66xUAjKVXGIoF7X8BYg4v1kmeGNXqtqsZWQT5uoetE5Ms6v/K
kUgKXC8PHqABHJBZUzKWzmUib/XYaptgXLwX8PUhQvp1rvPLnm+adxVX9+ew602CNbW8snxEn1Il
EldTfuoKU5OSkoA6QZ57S6YxoA4DKe9oEtoe/YxYUYlgOAGTSG2MviAJcdhW0gLxXR3Mf4rvxDWa
xT+glw5JVjF4d9UWwJMzEpUJnE4VyC7tXGdT6b1fK2u4O+aN8wkjZdcE3pdWRvGee/2FIsvhpp5Q
xnnEA/vdP1Fa6fNzT7aXIjJV/gR4+V5PfMvAr6xAQ0X9EmnroB3/qSCUPQQIfp7l0K7/g75J0Zrj
lKRDnLMDK0ix1u5/cWMRBaXLD8ef7L0x6aqsJulrrTk1/bkf5rvl40Ph/JvQUOpzxCJ8Xwhwg9eT
7wc6j6QB+SQ3fHzX9pVQnoI+z3J77fgPslRgaPKWqYE8WXb6gvoloBe1nCC2Zr3YKTsCAslmX6wx
ojjiQWlfpAJu4JReQgTlLlO0uJaziIKCNE3x7qQVfc3uRU33qBJcoUwEx3fpOLX9r+REQXZoYK+G
vk8SG1i2FeEi47sNKGw7NkCpurKpg6rbWvh853CL4vALwgsPTwt+Rw28pwB4r4+XWyMmE6Yyah1o
MQVXJdqKnym+U6cMXrIbnYO9KSeB0nXV2Agpm4DOIEYEo8BVWWHQV12BQIqn5ENiu+/MRuQaBGLK
TTTCvNpGcQejLptJdyQgLSv2Vir8POHWtfrfylJv27qfuz3U/48CSDTJOGWFx1zedXQ8LBtM1wbr
Fh3BNJUDQbpznDGSx1MTMkb6nhGPLUQuw2dFyOZ8NpRLEGYRwuQK4cUik5YNwBJtRh2C6Vj8GxKC
3SC9tsM+zQe/dY4KBoktGhVeCoH/2zueL6/UhADt85yZgP84VuiNvtxAxQiE8X3/GqJHTMITiYad
K/cX+oVBL6Wm8r+ELjR/Wc2pZ5HTO4l4sKIkj9MDrxfwWJVpDjmqfsuCKpfaNtt4HCixcWFlA84+
zJOhHMZ7sDJbuHkv5neoGP9L/TZB9dhyMs1U1BeyQQ8pkLd4Oq9Nyguqf9jhzrWDWarwfgQD0lI7
G8slR84sn3W/tPVnQ7B5DKDLq+36kOVN9W1XiLbT3C6p2niL3koLMA0lP7s05bhoOTtAXbvAaY9b
jMmVb3PiXwBOWuUhymcxYWiOLUop3BKPfMszyGrYHS5d0TLujwOYvAlNtTf+TvhdlgaQZ5mZfEVr
mPyDYTlLmUJJsjAiYcK85lCWYrkNlb8CND/WDAkDpGruPcsovqnqFmKRmzOBOOzykh79ZzfecM++
jtpcqkrt03Sx9Ed3EKtaiHHcJOsUoTrRVEgRhfNEsIEEHGhCcZaPfaeE9WYF+66GGRU8cOVeMetj
yGfftS0cQGQPRuQ1LXUR5k9DQ3mTzJIXUEBjooNAMF+HH4UHS1aJttxNT+yW+Y1IZwfRVTOSMcjs
EqY1C8AJUI3iCJu3c+46iOZqJxkKBUkiSTCcbn86jTQ1SIR6utZERFsxMkFdiuupCUvUlql4Jbub
82hVRX5fqL1YL2mETHKCZXQZUotGz4oM/aSGa99qSYBxXiaYdnwFrYRbZbt5LTD1X5FMfaO8+cpG
G2ohXSsV5oFafx9RhOY8Hw+dXEKwxDjntkCa1J/Isbn9Mdl4BtfIJYxn4HPwPV1x7EHZ+B4Di4W2
5sYuPp20aicuEaM0SKUxJdFFaUb+XdiKoUTN3ZnW2tHVu1927pmBf70HzYdhJ/PLQUCaMzjAFx8a
nmU9F4BahyUmXcVWMLrd39kH0lHWcib+fCV5aCY+NDXgyufR2SkXv53V06yZKgVdqjoNES7jtREq
0uASuibjlZbfJ8o+OebKmK3wcxPUH4WCNdrB4wTzBHF6nuFT3NyTjajEly4mhIsPEsi5HBOJVUz6
goUlTB5ND7EX9apLhL4GDonbY2CyZgtgPD+bD3VuWkTcz+iiQCTJk+OShuFhjD/goH/1/MiDQ+Kt
8kmqdrsuLGyqUgJfi67YyL4b2Onxx3/X3wiDRFeetl9QCLpgp+zi8f+AUqMlpRTwMloSYs7ThvTY
KuneUuLd24nKdYQHDG5QTl3herXnHBPSUPG1z8vrvwd6w6JLkY/Z91L2m9WK4qp6chAM+7rLmOHV
07KWrRbai8iE3xhxBFURgk3CMdmmqtn9vWJrI3P6fek06pKcKIRDe38+h42jrmYGFzQh8n+pV0y8
3h59vZiHA/0Zc9mXDappyx9r4VGKevaQUs6lptkF4HaALOzoObbnn8PQTyMHrswLEtJ/gANo70xN
AGB5HRNDYVcaWgoMuMebLMrKP/nAVSPdTasZ5SoeuNi5SbGyYkEcDbhLopK+Guy2RTdyh4qPx3qh
aoYpTVFJvXPfT9QLqsb+21hPSkWezwlPjCXI+oWfe92uaWty/8fL3En7oPfPE8XI1sm+vyXfr4n2
tajOvnyL7Da8UX7EHKez2MR9WZi85F5MJPLKyGE6oF3besdzib2ILrhw2JUymMmiyodTqkjX0qAR
mxrUSBXZPmS9GT/kSgdhI3/HqULQUEzQ9gQEElW5GdwS5+ZTMGw9eEMw0SADmf8pJuiFqQJwfqbs
dFNVN7qTHWognmZWkYfwQhxp8qdTk6VGV0jx9c8JhKE3Pr1dxTrT+FBonrt7nFeiq7CPqK0xiHKC
h1XVADlSz/cW6RfP5mgy+ucGzybt8iF4rcRhY41jwOmv2SdJcJMbgN8sYYp7W/6TUjpcF/34iqM5
2hphV0sy4G8Do5pISxqnr0eJ91kxffQrFxQSn1RgN57TyML5v2UflMY6Dpw0CQtHxszvtsfTBEQb
RpbB46+y1xbNAqGbXXWlUbk/3t2+u6m+1WSNSjij2jFGXJNZyYLSDcRdNLw++LwmZPu22VIfIq3M
r3LcxRCb6xRZ6IMO70d0apWPGcgYzzuV1SLU38J3gWSWSTRI3lQrXe1d11UswMq9eFIEp1tokxnC
LWLZhJsX54XOmwTpLW9PXJxeDzaZsYFYzMuymX2w6jC/oARzyJrVuJGkXECzGbH95qotz4CMKz23
sR5RjPWyyi8h/PAi5nulJXUXra3PjZ3GhnprJ+KsJ2hO02a/9pZ9rj2fmDsCUbYtLcoOjD5vtLM1
+wYuqKCcs7JiTE23fRSYRdnVx7vRupMLTpvBLL/dAF46H6Xu5TayJAEMm59gkSSKTlDjESiY2WSk
6ZnpCYgtLB3o4sZAMNozDF2wVlBXFEgDFUsdgUSGnIFgHuKd+JFdPCCzcGCDl8PpebesPn+hVX4s
yMkgjESS5/g7NQ0K6C47R/Q15ja1CI18K4iu+PL2mrNtEsPAWBi25YvPh1UPx6rU57cPTUjQ87GH
6vTeXEaUxzDz5UNK8qwNNmT01LLY34PG6VeZ5Ev/RnHp70jXiWLStPvzBJCeiiRXTIHqoNviqMSE
0+Um/yc2Nc0n4yml9rQ03uK52sEvbGMvKM9L9VKTCgnSXi5kb9Sj+kpCAnDeNxgpjSdE8XiUps7K
cjIM29nsZkJ4DJWR+kb/kj7ZG2ASVIcWgue63JF7xu2dw3LMrnFsffcjuKQJX6+fAuUwN2hoTQT5
9zTRU1w22yhtCN8C4ZupcXGzHTVx5PF6U1KcsXTfVVDvd8gCY7dbFgd2Q8IH7YLgQjjQo1qq/VrM
Ri2Na39t64P96WE4zxfyeqT/XGPOPiG5U2DxFM4uM6tzLMueiHhwm0UHHBk1drLFBV9Kjrr7vrZ+
xK17qMN6k2GvR4hJEH1toboLDgnB/sDn9B9BdRBTinCKOv48/owLnImwg/80MjQ9zW6GZdIlo0Go
sRFcoC0v43IQHv0wvA5bLJpUTKBmBdREBFb2nrtmz7t2a2fwadm1/ItO+4kwjtoXUxvN4WJsLH9h
CCFPj0q9TYkVPPFXwUDBlvvgL+ZxHEYIoej/Ik6SY0wkB5VkIHr+ErwaNMQsl2mCoagEUoERZHtJ
8hVhf+gRUD2MTz8XLaCpf+3ybuTCmCSatILi5bigcsiJVCU4CtWh9+B9ylIG8s5FMtLjIqXjkxWn
ji8Lb7Vnvv3EyEsdHD4mlSBQfNX7MJQCEuWAbE/kaFH+q67fnlm8tcx8qdpykwKiOvUY95NdPZzs
qEQOZ5eQL5dZVq9x4jOlkhZdD8EJRJ8m5WOS1Dw+QmfTgQg4yaoZVgvUQF0fHZcqaczO66Ea34fS
EjDY+8DfqyUaYj1WXRuqdAHStYVoXTT2fiVb2691vf6rKsybsGZLyfrRRJjzChtSf/JbqPDzjMb7
gikLCOPaXjlY5y39qfRgOtdM3mNuB5w3UD/J9udmwGQ2QOc6Ap2/OUZtfUw3sNjM2MiYJtAmdfiV
Mx/gsKA2iwU4RiJIWEGZ7z/k1WiGqISb78vZY3DwnAYcUDHvZNZsWgcTOGWAFwSA53ARPlwkbJFc
oX0QJqdHSF2/svai+L3sISR1pl3f0Ti9vWf5HQRv3JiacmFjih1GmEpdqvvCWeCuyeNU2ybe4s74
/9ybJJcpdB/rQZmX65xPBg3qhyV1ns1UM/LPMcXGitOeRNtxJqcN49opowzcVFvuDWUTn3eTGfhl
M5XShfBggzB6je3fEqtPaPNoD8nzVMikQHDKzhZ4JWOq1qlIjuFPvmr9hBjVReKcEwiiI0edGnvT
Xsm0XoPfUzCTLVjt7ATfcnMYw9L5vBycIq+AG/DVnh3On6u7rzpBpfmy1ttROEnZLtUAzyzH62aK
wMnCIuZZvFlwpJ/STDQ6MU9rMIwQTOfQj8cz5dsV+zYAuLAvzQbJcUhtYOmeTc01eBbHBrCOPt2C
X4IFtp8kkmpJAuTQol91KythrFbLofQHhJN0ZhHJwO+B98wfX9U+UZP3WRkkUvy7Ae4UG7wl9VME
blUMQrKd/YTU+LQX2uWokDncEbeTEssGWOaNDlVddY/tDB+8FoXc1ytZGJ0wlCSFPEiwmoRkebbD
kxlrzsZSBqUVpyCBogPnGheyKVy9JUAiWMQBb2GEKwQ3Rp2c4GaAvjAhkDCI0TnMWg2RmxRxjRwZ
cE/ELfJu6KLm9uvGXP5cLE8UxRjW6W8XNPPW927IhuUhiR3wEYfVh7Dbp/DiQC0H276H1qfA2H9w
bI1RxsUELoC7wpejllI2RTkNVV9jdmBuDt/9L4ruO5P443ZF6YBgWRmK8Yb/JcZ9a/QkzBGPkEAg
x8R1kaDfdJqiAvxOcTb6l66iiCUFbQoRFSwdnq9B556o1Fh3X0UoqDpKBrpHXTUKFei04Z0eokrV
0lOWOsUiX6TWOv2tHr16JvUBH6yLQynj3LVmyqLQzde4Jy6Oz8rA86/dDeCxrEoG+7sywHb+sIEx
T7tfZmiqoMXUEpE/5Oar18MBsQ7jVaAKu8nq4A3ItiXDqQpThW7dp7aNZ4QZKkPHq6sOhkuPVG9j
+m3mRsKt9dvCny7pAGvenoEvhnhbOoRP1SFFsm1CrSS+ZiNV2H15DCwGuqVHA6MuNuafW61HUmpV
k9QpmUZv274Ld6bIIoEk0omQtxA0CjyNvIS5VjHBMyPgO3ReHdjLrbmWu9+gj0wPkD/ewvlafAtL
LeERHwH8WrYz7n4na+Io7AMdgQ5KDxoi5JXtg0DxoTYUrTzaysc7t+unEbhdNIdbxBF2223ZHgfv
GMN04sy8rUdaOF5xyKOj/7IZaZKUjbP+nOK5JD8MbgG2MOsrh8UXjRYxJemJDo3GFBMpx6C3tghS
kzFMNflatkIcGuFxMrqCdSQ/LbbgF7fw4hpwx393+epjcElUdXJfgU+q15zme0yfPbZXY9RDNxqp
XYkdJ6QVrK9+gszdAhxZfkLIYasICx+O50B20dHoIMBuo3XYe+AgjlzRIL9ZECEDUgUmCZ4Pd6SU
+gTiiBbg+WGFzxw6dggQrXf+fS+Xlt+IP8+cuX+Nx/XlAybOC+/THiWSjqEnSPAnWnQwKlvBB+bs
zIK9o+WCRgCZfZszzqvfGAhY+gx6PxqYV0vzWZdhad8VdL1MKzZCAKZ9P2hFvWqwfBAcVls5pmUK
7d7j3tTwbGEa3pm45nNtaK+Mxbj1Wph9dhAv8qDa8opbvNJWic5SzmHKE0baj7raZ0Ud1kis2tHx
QShxKI3AV6l3Oi3oAAEt/odSW4OCj1Z313R4zvVx4EuOwhYhM9JNa5lSd0CZYubaJwRaacc1hjT/
r4WCXyeJcJu2P+Xl1nFh9XK7ttH6pI5N/d9upVornppgJ+voGR1SlS66r8/YlCOYzzmqWhSemgoV
+PKgNfS8TbWv8klgVhfrfjdJLm/8IK2Y4xY2shXtX/v3Y+0AV5TzVUtoY92+JZ1VS2HgEnA/fNLv
L7Oz0ZzlrPq78P2skT+OmCesCA2KjQ4felS6AUWHasLSW3ia0H9facLNtNLnvDPgOvQm/JFo7ZNs
6tdxbsCXykw34Ik5S4rfwI1x0DomXK4QNvtEg2kktM3Mq94M0y5Cow5RVYNh480E6KssN7L69bAF
jAHtx41u/fdiNq+qeqqan6Sa4V0q4u+jIHX9LKebw7AOmrT0Ho4CT7GowYJpbyucLzW5TVEuNFyV
RsZRGONgKIc2eqEtkAgxl46HgFNCLe1eQsv27HFNLS1u8vz/6orSlmjhCk11yVFK7lQ9tRTU8Oyx
jK3v1EoI3S0KGjNbh1gYn+fIC6Ce0F9sZo3LTVc/V7G4GD0VH85pQQ00IFkrIK7VZdSkLbmcC6p/
KwR6h/edG2lCe9W/FmbQnam9frFbqldFHt0m88R7oJRxABTAL9OTVoyhxNl59pyjrXFJ748/91J7
BC8baEagOleeRcomwtLz37iBS0Njv7h/fzTQiPjfmpTWBfhQ9W8sYnOQ7xfu59TxtV5cOB1Fz/rf
pSQDxo/xycrVwUMxkSAjsgmTZaPYTjpuW43et90HiQjSxIrlRv32YWlMPBfmoTsom5aVG0VPUC4D
E9/M36aRhG4cYvh1cKDH4/fI6DZamwdhUKdUWForcsD8vKOagerL/kgmkW043l8yXgfRBbu90ev8
suioYzvlkrkWyL2KkmdfkBuaQWqBuDxPJDkitTLysliD1RHMyFmxjs/fNTfozYtRxU2TN4Z/m648
KCZ1MX8u5szzS7910PxTpR/aaAGCgDY/HDb8a9bfKeyAMvKtwJaFMJUAsvby6R7pnjNqXgUqhpsZ
9BeHnvSJXb9ILgHfnNRSfoWLkwCrZdzAhRWGtwvMt764GsWrF6ioBfKXoMYht5CMdWWUkZxz8I1H
Ng0q+6W0Dquf+iXR0gwOtbrZBgp0f5Nd0iyCnH7Vc1Yz6UiNOQqG/oJppex/iIhUNIQHHmCwNVur
0B/ksqXbvrTg+5OZt56RekwfaAXNGHVDe1xxktfnbJRXehK9e64nseE9YBug4xUf5JCOgQhKSuzY
0+lNLKTU6TVDVV1DK0MuO3Z1agSd7Si1hXOdDMfJ9CCqP1gikyUUEW8z0lzzTN6gUWwHbncQI2H/
UfDAI7tOoLm+fMc/YrEjYq2gOShJIXl/vVcRX7NzGWxtHRk6PbjHBvifpnnSPQebIXmClQOaT4JN
ACG8fwtSmqS7rLBIgsqbPBJrzFODjxOsg3q4aHq94z+bl2nWIXj+scSVlhdFjiKpEfg8iEKqsaaL
2QzPxpL8ExBQL69Gfk22181HXf6wh9sa3FtcUEpeYo11Fj7MZ/opHQcovud8rkTL6dpbdSowqXbr
n/4gfJWfRD5Sv1RkinOjfqwPHpdaBgHD3qsVnGvLSdoo64u6pLKmE5Gfa3FCJMQ5nbFijuSBDecx
iziNedEchvE1+21ldj5mJOKu4thmZQHNu1FtD656CpPYzZjDVYEGVScp/5eF/fQxXXqg+TjgMOlU
OkDtcw/YWUC3Y2wVnLdAAWOax8/md7QfnVjLCbUCj9XVAVs/h9oWRf3BZcST5HzAqdYihzflRXhf
aJY9jYDE41U+SJKsRAzJHohzJSSu2VPYiMP1fNKZ4wF1lp0HK1qGYeyUXe+EgcDEUdU2AwRCbCdl
qgRZdo3pK5p8+2XSMvwD+iY2FvaCNOrKjB0yPW+JIsbIABz6hmP26Y7aoAeEpGra/IkzV0TW2hHr
/Q3NIlsanEsEFskNvCjXmJWNWkTYAhm9g1Bc3+oFfE4Z9IBX9Cmfnj/AU7qi4hc/JwUhmPjjF2SU
GgI9zIlIxucHluaDqzC0KlUGp74bZCpM0BmFJhp8PCTWaIf/SRxpYZkHynMUFBnIuGmLAMplNsOn
YHSO9ELlN9DKLHIeAP6UtDYckOiu27DcXlN8mqVxYz0VHTGNPD8Xv3wwQBZ9INdxH/7pYY4M3BWT
94wlBn08CJQ02z/dUdiJZ3mQb6K5QESZhK2+ZFcRAp2EAI33nyY8tdZdPBcPYMjJBt4I5C1KMi4E
+RhiaTH+yImkxSaYU2rub5YYNYzOJPQT6NMByqeuo48f4WcH1ORU6e1Yr8LewAgRAUnP4WEZoiUv
0pbcSVOOcVHdiijTPsfC9FYzwZdI0g/IOU4rPFE/pVsioK7JF+NZfHkBI6YU8UbCvU59793/NfvV
VYK2mnLiheoUl9sogCM2eiUquq005n2OGyPgfUdzr5t4x+isg+X88Lsenl14IctpEO5AuA3ZdC64
fUAk4H5+l6lsxxicwrPj0TH5kW7GECg9uI3YaHqFY8V3KTkvmdivEqYU4cX1OpRNjp5/kQqq9xIP
XQ0vOc5yD16+B813WWQPZQPw1t71Ll6StHOZOIKTL3nvv8vNUDg+mdGYnnEkK6DWOC9vuq7GAiUf
CG/Dfqq+rcwzh6TAmi9hatkf50cQVlx/z4ZMc3fRRrti2c3ByFQ2Z9Ay0v1yRUtDKPS7EVCCriI1
uk+OGXf4Qfgm3khnxAkqZSDjvGr63jHWrZHDILXUwzBrZFwLEvNp4D0wyKN6nUUlaOC/4e4lnaau
K08j1KJklgdzMDjRWBJetrEIC6OutBYLEbeGDDLTOYE0dSGn/zd1dhHt9/IfcuFGMO/M0G7IuH9a
noxcil3tcBt/k6EdF3eaLIjt2OpmJDHZHpjMCpT32LmJ4wO8cIetBDICyRoa2EsBnV4spNkfV0aA
STlE5dfLrfLrM7/o0u+aScJMbCLaRDTUVAOPNngJrhfZmqylYCEqDktN6/BPSqUqG2dQJE2cymUs
sAGXc1CLpsk7L55pwHssuZTw+cr+yg64PQWLw3GNiT407Yx9Lcta9u3pl3sNJ0n5Eozos526Ff3z
9VA7kludJQW7xPjdE598kzy4fxjbhRIFe+0ohBIwcyy+hMiV5hBZE2RI5UDoKp4M+eKC0kDp3qCG
QEtQJposCiSDP4Cklb426NnDNgsnm3Ok5flVWmYKk9KBLLDPkLvjDdEOPVahu4tejh2KjLQFzvMW
+kb6Moi7KcdfvQ9gUIZNncS0LSWyuwJg5UmPachVg+qG8cV/aDWj/K8mlCIAcnflzvGnHVt2DCn5
zd9RgEPb5F5rGa36G38U/cFSqfvSvr/Bz/+2X7Q2TTxYS2YQ4wIRB8ft4U8wm4yQxhsLCDGQtSBq
UrXg984OhBVcTANT9SqyRRZ9CNpcMOpq+Ds1OEjGnXqpXfpWAgASlcwrf1jpIbiyGs+rI10vmxQD
t8Qnwf8kxzu0kJ9h/JdUNDho7t31tWsQ80W5TYhIch3G9tSvFmIOeP9+apYlJMFJ/i+T/ZtuCF+t
57T1EnlaO7RM21snEHH7pZMbxgucfKyPCUyuZ0GN7HYQDSmhxRbyqffxp6yDgX0dGVA9ANG5aNUz
NsCtAF3ns/XfdZ5/3XVrPbuhBHYl95LmxmB4BBdWzyN6KKGni6PbryiWWvCDJUenRihGrx5icQgC
fsE0mTh3rYyqqmfO8EwS9DxyJcer5l/q9es4AVlGyEYBQLTLgla4b7VTz6w0yrPiEBJF6MLUfgsn
VwbVeU+OZNXeJeX4QSiGUzM5i50j3q15wgOmuT3EOctBO6Qzr326n1IJQ1RWPQfVwnsmAusDYPIR
raLGfoMQVsAHwGoHs4F90EDI18PiVXrlpZ10XLquPXbYEqH7VaFL5pxldfsegyS4oIR4kaeYmO/F
d+tdjfQ6ANzkm57k7gSr6wNKdrAZNk1/grNnWAYBrGR0xRdL/Pv9DO+9j3TLTGcfW31OZLmF86oI
Fhs8MbFHJf93cLRcSIsiXcd8pKf6NMIdxgGK8p27Wqg/Y9vmZW89aWnsb7+bBC0Abr96siB3PDDS
lxfDBtxc/T8Sy8aP2q9oXDTExvPxdQHMlacKK85Wym2RrLaUUHFDu2v2dGOhOoRYAF2QbpbdxsiR
f4DsFAxro6Y2p/SmmXG+t1iayXR+NDFjGx+RA3j02x9nADnOVKevyAKWk9U4mjCEWuVjEq8a0aAS
KvExTWOwiFV72e5gVV4F8/IjH7ukH1f2kP6Tyiiw1nfgxzcfyawsiydHupFu5TrdeXUFwQ4X9cQ4
ZYqey3rc0hE30Mv6gNayYx2orGa8WqnKHGGU9P/uz+zTNsE1pt0svUyuy1peWpiyx8AJV3KDpw/x
gFMPgMWjhyizV9Rs4IKPvYaL61tXzz8v4mi8s+RfDIbRbU0AhKzHSLf9OGKItLMlD9iaVolXnMJx
2RiqWpau6oIgaZcuHFP/Z43XHfc62pcjVlxR48ktonPAmLOWd354Ev8M4zQ9ZgpQ+llAmvNGlQH7
ehADRoO6BZDVo/ytmVLx3cF89BkihnVoxIhERPzOm9CNrx+gfOWQIABIL0LdS2EvprK//TdLUWw9
PawLbxjq58ePqZnG9l6Q2uEHYyYAZmvHrVPl4bmm74y4c6q3JTNOS2B/CvzP+tYNxh1UVbboOFPV
bEAkXvVWaLSGOkfgV7bOaddY7ENjwv9fJajkDxPHBDUqWggJSClJ+FtMBNBf4dCWYRFxgvGHpGHu
VgV8su29hl45Md2gSJOeExaRMa7iILVc1YR5JZo1/wqI80gLAuTf1w8/SERRDUKBaE0rN2dH5rH2
L3y6NbqAZugm3aqChqnVcqzcPNVyIR44GmsYDVbqVC8whjoSobGUFSrZT7Y6e62LqIDFCExXNOgJ
RwqfS5eJ/IYTrQlU0jGJk+PNFVIm9epytPHKQc6ptgJoG43DEYEMe9jmZS6R+112Ssuf2YfckEtZ
6LWc0KUC4CUqCIUHrf8sncb+ATMvdUvlsqr4Qc46jxKgX26z/rY3226NwGpj1Wj52yxwL2BRGp4O
CsjdSLIqOT5bUpu06NYIB0yyQvH6JdjOkoeMeoxvtbyGH+NPqkCoWYxyAmrrAwEdXDHt1mP2fPxj
lml95EzIAsRhttHqz+sqbkfiip6QQaRKv/uEqZlyg0KbM9TwFDSSynV59Il+f1krejxLnUAnS4qq
I/TljJPgLudkMScuJkvGjNqNXlbZcAU4Cvsf9qVkj4fJ4Um+k7/yoMWxmcNC7LIzLcVG/athwk5E
MhOgRYT1cDO/dpiFx9FxA1c4r1/AC+Bd1Zbbh1ncOfLy2r5LYbedPYi0uiWdqCyqo/7nX8lSYfcH
wlxEw2DitRA/w+1BOaMAi2XMA5CIdQfmCdDmF1ItaqojF2Y+/66i/n9P9RDSeP8UuXOJexO6yhXQ
jrRDcbQFaAMafv0t6i4LVf5JkyBEKleyJ7Z8saZlk48DKT3EOmLCBgos/aQNvmuBie0VOebjW0Qg
2GLA8gF7s7jYo4wehU2KpgEzFuS0VDgx3A0L9eoAULv6O4Vmp3cX1pEcY7ymkTnr8UwsoNyHamck
D7mLv4o3QQR+gUVWChmzxQNXBWA6Gac9u7Y99hasP4Vu6FZRaHOdBESYqHwblzsTSEWg4WtvdX63
sOJJxdhXAeccjDL28iMOAupgOH7hO5GWBFfLNqj1Wq5RIryZVhWrkhfPi3v+txugHA8Alii/HyOU
pxx3UOBMC+UZXPsGlKpVdYCopHgq3DPMcsYoUSBjCBYJvoYc+A99kXQZuNjfcPMyHFp/zJk5t+wu
00BZPrQsLO1cVVOIsEk6BMyB94BV8xPiw77BRAU7f3+3nzDqF5FILmFHEwDPxl3Y1ySpALXXNQh0
St2HfcZ5imE231cENZp3cOynMemqVWUXJ/rXDskv22bcjEjwfxDfLaAAXfayHPAcCtwqOziF1Ib5
6x0SEF8/xs0SCXxXYATgOwWI/j7o/56j0BvpAbbLo7Y9SILxamPLrVm9RipORRPx9GKLIFu1tErd
g6ZGhpybLFHbeKCbeNlM3DGSdTWnymQiSbrQXjqgcousLogHmgH8T06q8IV+j1aEdFd0YvPbJXWR
LRysx2s11dHGtK+dLwJuM6okx3QXxHcx8BYy4Ypf4mz4cJnuFGcZpkDvT2WqGb3OZAStlSalkkph
+Losya7Zc7S8D/6BVhje9AmlvKms4TYRRPLSILjtLt0zN3SeTX1roM76itr1b5q/c5iSSluw1Hwa
XIzxp4GAVI0u/Kf1OakfpjhoVOGpqgcpz+4OUux5MJWJtwfyIPSl1Kzog/HlBzn9WHsbbWPUKxQK
qBOWtti8tBuNgT5h1i/u+VApT2WqpleT8rk8KowxYKNVix5iexJR/HYGd7XzdDvSPJXhWitqjRQV
iKnwa1tfqxW9EzQmtCmR5FZGDZczI0UznYD/Etfx/6z7ix7k4os4X+Lp6fnA2aHKzRtRzBrqWG1l
ANdOi4sLmGrumOT1/nOd5nOuA0jAjuu2tD9rvSkUclS1vvndOzT1pPaFVP915ewgYsNcd9W1q2Tq
mHZ4g+q7fJQAhAbdzo85JpH64WBjKRnPkXZkmcGclJCQXBKXlkqhVczmcowXYTA0M2kxujosgvmh
yvrQria5DpL2WK5lJv+J0KPg7XvjTKVS2y5A2tAdqOiRAT7J0KvX4/cybSTAn3KBaG8Vk8n19J32
wyjXP12SuBDO2lsptI1UMRfIJlWBTF7MOFecYLK+lHiM+yKxseaCIf0n8R54a2teSan6s1IyagBW
XQBWYHc9zsCKUSI2ZlfqNEdDnimAVQHK1J4iP1e4rKCMkfOoP90H9n9/W27hyamNUf97B8+hhxgW
+afB6dSbesqucgVkHwa+uWUpNBXpD3WpIhoxnsJlPBGdggIpDGEVVU9cDnGboIYAPSLXGy5+KjSR
AzaP8P9ReIE2biXN9shaoP6yz0QAlYB29xatJUQX444vjsmucui/bdzSfYQv+QEYLnvpf9M0nALe
JumBUs6cKuKCx4a0jW6N557RYB88MKS5Oyo8U50cbHH0sDlvthYksDx3Q44C4mJOmx3EuhE3nrP/
v74UqcJEwpDZJNTOP5ntIgeti5gI8FYJc6AKEAgTHB+RzZs26EIuYQZWKBZ22X7QUFf9VD+8AxkG
2nLWwDcxrQT36hgVZZDna6JBAvOmGg83evFkx08Kp2PZ/aKa3g7GDKyrbfAhdVCQEIiD54JidyGT
vc0lL7xlVwziDFhgo1lBjuPGfS8OUVDbFvyM+twJo2rt03dRlBTKnXzFjxM9FHCVXwo/MIGp0qGP
tDSV4U/RdCRob4nn2TBxzWENVn8tUy9Gq1AoAlTsoHTM1I7JuJ/Z+Fk+8zJIhPUTJM9T2I7p5ZPM
+MDmW0KONG6Y4Vp8eYvM6azS52bz+5lO0xQdPR/t8zHl71+DMWV/85PCDrW92uSnBq/SnW15YOmr
KfAAH4SG15hlnhETaDXT2rpiXDLowbo0E3vlZibCB9lg2s6G+HQhBW5VCaJl/jtSPUcP5vu5NVAh
4oED92H0TpNU6G2+SDIXip6JwPxC96z10tztqyyYaoxaK48b9kQaNqyb1lCsTxSMNsY3tcO5akge
8xR5kd/SavC6mcYmDAxpPJCy/fbqq1kdZOZwN5uUH+nJDkErT96CdGbtjUZsB962m6l7JkyzD/kU
FSM6Q4stCoCOipVpUDmIgx57F/0FNUL19+I25NYjMuuULDktv3zxOUSak8Lgr1DGv+qRLzrbGp2H
xzVdo+3CTubIPml6eL6lEqb1SXfK+iVX4nLn2rjFKURrnEbdLEcttt4GfTIwi1iWxWfcpLHvuW6+
2hZaAqBde4RpKeqp6d1mjwZ2VRNDdtvTG2dTodNO5FjrGkV8pasKDbyZvB2K7lsAENFH+6pE1rrF
DB4r3MGUzkdPbM7BOzQNLMI17zqXSodxNNym+TN+G7qXWdOrUupMCdWF89lcBaKYseq+KUdqFsn/
3tGx2/tQdhpC2MI0QaYU4GEqRi/imVEulgiL4dUA0Vl9+PVHVvAqLk8aRQHuygPE0VrjHDoUOiys
3axYcHWYw5DCSA50UzaW0cFsAt1hWOsPVQoRbk2N37MgFKS1sh160txum4t6vKuPFejsAms+4arX
fpTyxn1B8LE0uK6WUdWEUMUseRzYWPT7h37S21nPGFSGFZQBDHMgsZf943LrJHrFaacjvh7THoh3
chzxawZi3eeJYZMq5PFaZIcGSBG0/HFRMEQc+s9k552jMH6iZKinjc12YcfB3qqNiRGEfoGiXrsk
Spq94+blH3G/GJ1FhUoL2mzNtLbrb21WPcEMJPXKQKXEv0w7+1IJD2aX9isviSaIxBE7m7ykvaBN
bVh1aaP5zc078t7ki9G5aj2skrnj3JVnjl/G14DzdnOkemOcWUPaLsrvLZeLgr/kB+wN1UecWXgC
NgHv7M0eZScxrHyx1ykVl/ZcL8tOgWZTubcXgkB0P7sPZ8jCwQtJZ1GDJsS1eAqhJgsDhtviXnzF
/E8EZ08kXFnCw6FFdQgvCjHEqXuRmyAwTRXLAok7ND8xzTv4bLA6Mp7HxEzFd++aUHswaEdrySBM
dpCSjMte6anolZR69OSenpTNUNcW+n28mlcyoiFWPDswp75DtP8sVbFe90Lo3yjqtVo6WwcaWDFu
dYw+69IKqrC636QKJg1eQSzDltNRrPx73B5PfaCLX6B1TsInbSUwbaDhfH76N7QSUtTToURltbKc
1QAk049eledYWZxZZ2VOXl8EakLqtuv6sROU6gRmCFFeORG2VxOAlXdVT9c51+SHulCWXgSUg+/Y
bprtXspxWyRCxOJXXqHq6ak6WXYy0bxZR4M0McnB033RwiS+RC7s+wWv8xNjS0Y8XUVuYABtRoFO
Xxb9rCNuX33Rg7uktz1Ln9pPrpX1+w/MLcAZWuX5rF5pB29RTUa7rgjUTWAxebuV2eg1qpvL73m/
SzT2ZJNWo1kwJIdv0k8lvZy4FUOEWm3ukrElCcGm15WnAaCzgxxqD2LDKyP8le75pZdwfOJNbKmw
Q9US5Q7GQrYLBZ+uSCblCTERP56GrRngbz8OnBCg8Ebgf7uxoha/0Me69K/2H0FXM5yKBna/4TqR
fx1fswhawhMlgywYb1KRwLsh4IMU2YUBP8IvyoFiPDlOtc1HXmHcpqBLM3jl2mO57SUZi8oJbqfw
Rm/5/3V0IVGvBxbOaF8ZR17oWc//wf5rvdhHR2v1VVaCOCoxjo+Cj7D3BnRVhUOv8r47+l1bdBpd
72rtWMnCS6Mk76BSRUGhpt7BdpfCA6PO1YoPjN6wVhnE+SUPBoejhzbryHpe5UmYbcjSypTjnX46
wog9lU2J23lL7zPH1BjMo21HnBCtz7Nd5Xv89w7iULt4he1F9XKXHfeCGq4Ojz1sruU0BYyenbxR
NAmseozhXHBwTqknrzOhsPkGaMl/mDcid2D6xE/W/bl3RIO1k7atjCp1LFEP4bZKPoGm3c80fA/g
0RRaNzMG8BscQUbr0fsJlp985aTAbgisU+DHhxRYkrgkUFZX7/6CETvnYDvDobcgCVmHu8PD/0vs
WoLTRgX1TaUYZdxlMTN915DM4Q31XrmBf14OMGrQ7QxKuzHVYpdkNVluDZ0LPhH+9huFbMQ4IlmH
992CPTuxyMp7AhZqxWKzr365cly/ts1eac4WnrZ2uNvNuWlsvYNO/fdS7zKhwOXbU53GMxM0rpqd
dc8lOJJYQMBUS/9dvDM1BDhWoIbSqY2jYR0QOEtv2UBEJBPY0kdC8s6BV+RZM9Guon7m4POJHXzt
0dE6WNP0xvl5QOAP2lcv/YnYuVWNRd8PO3eNtydSUErlaCr7CYjRbyf6pvH9AEpK2UM3iheMafEg
8m8KNmOH6xCC/gCMLXVJP6gsBdTLKWcYgpyFYuSWdahm51AtHIpmis5xdMxRGRiycNrm6nR+il2a
tWu3P59c5+Ng11gy/yn1Uy+SxdIUJdI/ZTP418ePXoFdKKtsX0LS9vv3M4CGOMrn+6hyKakrxBfp
AsC4r4XVBmX0zEtj5+Ju1ZGAgwPeBBB3E8+2z9air14YDxu7lB5ynJ4fyGsJwrDIBmOf3OhEMs8i
LV4aOaWmR2O/+piRKM2q4QYmX3Xe/HyM63r5zZ1WIIPO8/xMFu6lf+By8e+aykxdF723kG7pKRwG
4NMJy9v4QXraSBNLDapHeJMZtHg07KUqrpkWq7cgi2bWtJgcNq5tR5kvk6qYnsJ2hQv3TjoQjWUu
C5l3/i39ugDg8jzA+Ais1X37Enyhrp8GVVQFRCjvBjMpxZ2jWffLlZpvT46mo0u6BUUJbseBo2Jm
qu1YVwZniuaFIHfNhb4JBcKFhd4nifhdMTj7olRNHYI1oV0TM4PGiBBM6CtSTeFibHeiBvcnp8J1
lZoK0cf0ZgBL69o8U65DX5yVvNtbhPEzjmgDfRTK7PNjg2pv4ZD8gNCigW0FVuOwxM+Xt1O0Q0Qu
868Y7VasmWbU9Df+hEBiTuu+nZ/ak2WONlvZhbPvxnTo54bu9zzEkCIIBa8NPL9BVfRQsUXZO21v
nNwFoCUWpeiVhti9k2NVDeV0glqm81pkbFXgTzlBZllT694JBwEfd2K6XwW4KP5S7pOyn7sKtH3O
lnZKmitXEwU7FNyrKM83Bqwg+8hTbOP2ex16h/dFrhUIuUWVC5nTglQRN3tYWc18LIQtUS8nisym
veSAyE+vrsGYHq4XefNOa5wj4QpwFAFX1IFB44TY9wSch7dtOlAPeA7csCYUzQ8kyncbKhB5FyhO
Vpq1k9WWfEjNDmTOjYLoPQwFRcKPgAulaRYxFW4yNmrMGYs4x+r8j8m35Xw1Xr4VPYSTGpTS+hWq
a0iRYCYBWbdeMOqN6vNZ3T0baSJFBKQ3Rax4NoOhAlGpK3YloDbsk6BX4FPFr0xQHxq9vRcUs/XV
NJmMO1qmOrMmZHqsZLqdZSOE6+IAmqBv33EtAfMJVuvG2vcrxsIWfroCZQ5TF7HlN7dqjsulXJ9F
SasEQuDXeFuXHKrPlNZZuPa7KHH4yqRSQcbdKDr1xWSTxS7lkntYIYfPfrSGCVp7D6nmiO1Xmp/u
8tj4jgF05x3ckMNj8vQGQ8KrLS9v8lZ7nI38OmH85dWzkXfpXrse0jW9eV6x3vtYGpj/Y4x52WXU
EzgLXQ2Ht78ImJVkATtWVf2xBYjDLuPjkgxDkUJzi6nStk/YDFTWAKwBplLcsRinnrie5i53hGjT
KFHFMnlM3PAdC3ZS6W9Lp/mCyIOvnttrpTF4BCodZhe1FtlV6k+jMjrg69RnWCc7+OsYMN0axdBk
WjfAfmubaajk6kaRQSBPKBwt/BMSUGyU4yJ84kjnE+DoIchIyruNDmr9TPmUDkqlMI7N69+Pm3sJ
3RQ13mrUjDFUjVpQauqeN3b0nTQSapUMe7Jq12YGYTrOX5bCn3+8m5MceqAj5h0J9a+w7+qWWhOU
8EyEHWiAnLUy9MuoqqoWSRH8M9e2ESBopYQixak6Hplk6lbkuR9UJgNuwcBwxw6iJVB9KKqjDh0y
qWcRh34NDCjgoW4YoNZT3QbNiq0vgxL/AJ2Wheeu4yHLlZi4j9OEp8wLAIvVwAYIxI2BzifUbjZ7
ZzGfUpBFYdDi5dtvuddslk05DhcF+/E3+p1cYLUA8k1xM5EbRDllKUmR50+zrqHIEO/kujQjzwm0
2mHFffve1sHJ8Fa/F57dLhAiN/UCD/bn++d+hIYfz1SL7Dfy6H0omNpmhNY5V4BivakSnPYJdMqv
EjhcRpkNyhj+H8NYr9YTWAqUwI/5jQFxRMPcbiJLaUQ1D//LdAXA3Ay+5nVM6mG1x73l/q3y/h4l
nkLs0Ctc7j/l4vpjBz5sDAe/5fsEB1IfsPuz3VPynJvH2lv6d30sdDcBGpCXpfB40r2Y+zvlew28
l/uhNgOpXaT7o9f2+8QifF/oGDlqVO9w91CP1lXRSfh9NM6+OI5cIOYDnQJ0m1QiYONtnpTOhncv
gq5w+9DuJ6YuTGIP9pOCC8vDLgYKBgZjowFK3uE+QVS7F7AP6xJGmw5YtYWJB/8o5LzjR/IF4KEU
7rJLvQMEjHBCPDDts/+AXXVJA2eEklt+9h6RZ+R2Jcs0GVaEz6jMUgWvcgHDIz8GfCcLQCZhsUp1
2P/PdORw2Ozo/va+RLLNMwpotwxIRjmvB55KhdxDwRR2enyrQDUV9jNQX63GS7u2VOv0Viz0pYBr
dWAeYXZoqon7Rp8akteQDU/hlbCSgtsn35jK8WaUAYhjPnKHL2wRKN56GKXXk1ifqRIe4ReTBl1u
7wK3cO2+mEcdtYFBs4S+qn15Bdt3QKCm9tbvO/I3V0SFAseQKB23uSTByVcqdipLjMX2aBAmd7pM
/NKxj6PfB4YJV1RJxcuuc8R3hLHQikuDuVhOLKY8NtgnPjF75WWrkKQBqtwsWLkzUkB5nuDb9CFW
P9bd+w/GdqTG39mU/YQaTjkFpukxjKnxCBqDGXocCFGRt0Fj4kdW3s29vWJ0/xyRmTNfBOt7VVAX
ltUA04JCSdoN6aXAhoYXYcKa30AWZi2PC9LCX1eZ2xnchecMC0I/LU5tTzBN2Pr0qH3KpBeL4WMR
DX+BnOoMePpp/MN3qNxxcDfI+bZqo+5+B+pbzRM/suhUdk3WaW9MGRIlwvWL5HcCgoMgzPJLVB4e
9d1VtXnEijR/fulCZynBf5kb4ZP12/qQjAgv2WsuYx5PdlWSOqi4KqDQ9/koMtKVa/xsB8qWKo5+
rZcBhHSIBDTaXEf5xKUJQIHyp4vRKoiX0VPInoth73tj7ioFjai473nXpr0J04/q4odkozINRVQc
mYq7fDCSdljYcok6Q14zXbauAK3em0Y4x6IsYCru7/NI3khvDILbLrRS3egE6GhP3oA1y1ocd5dP
Bu+OnxNmj5cCDOybpSyiY6hi4vwVD1IY1cuyEtKmcEU4dpv8lRbuQQGI/7Hq67boX0s8eykkVVXE
zGjGhJmR168ry9wqySbtbPbBSntbRRiP0LgX7Dmzw6BluOfxMyIyPYi4MRZ5S/BnsFx2RPaAUunV
+Veh0bBRlUkwC1f/IuRAL9DA9AfeveMidQlO7YVafb/U3cn1Gg9jUr12sRbhAvuAgD7HLggGaA+i
Aq8vaIWf7U0nnMrOt8XbFdgS6wK16jjPWiYx/CA/ebPQAmn8sNTY45qjUou4yd+0amsTNMzYDNWT
Oa3KYAjCoWETOYi0FlJyld1IRgoKthOlMdFwtoKW7CGKEF+ZwYw+85WDvEET9L6kZmPs91hXOlDl
GcEoedUZKCsgNk0nylmqyxSlZCqoHI+OmAQjOv8a+g9NC8RSC+Xm3+w0hUr080Yz17v/D9QtjecQ
MXEqUs5dUSyFDpIgIe1R9845wP/D/GDim0WeC3g1JIHo+LSGqjb8YEGVS1BjxQII89uLg6cT1Ezp
XcxDHHitmIfGkYEI45GkAVwrLsTLvAdRgKx8e3/UH0nyCWUQ2dhiFTNx5SqWzL4J1nfMh1Sjqf/8
Y3Uju4CDAUiiLy7PSghpticqji6HVEDaVunMqx02Xd8JGwERZo37Vc4TxMlItPXNgxPiAeEVHdeT
nRn/Zzp46QhvXsQKP6JaR1sHbkr9/QzsieUU4yTrPJ2CSd1cts3zZj4XuLg3yDeO9sEgqyDIzGSZ
UuVxP0d1fHwYCBjeyrQdLsjWk3JZQAej2dGWXYmuQMULznHkgFEeBSIZ5Pm/1gCGywdqXmozRRAb
MmBESs1JVcBAOvAnXbDRtrkKaQTjAN0RKnc+s+5Y+iyJbQAF5Vbniy4xsLzslkwJoHF2n/fFWYFD
ys5/NFeJcsXekmdh3WD/P0P44Y+LqFxv8hBIoTdG0E3t+kD5EklD4n2t/AZtm4o728GWlUBQ6EOF
jmeuDRfngGgDJZ+58qAlRqy4MZUMlXepYnyhusdw5MPEQYRadL7/cNLb0Zr98XZnB6lOOLU3zSQC
ormbhZ88ec7ptsdL5dEWDmSa3c2gaLYMyNVDHtLAdi4asOjhH/B/Wx6HQWsk2cTBcAMH+ZwucYV2
n2zRP09gDbNCJC10BKHCsSR1HjKNdUJBl9sL0IV4J3l74naZR01HuUPSO4Sw7CpZG9LAdH+HHIf0
gbTBwgSBuT6GtSF0M6RFvTokBkDdG0QcjGKMMwDQ3fOs175DiLyh1qijBAmNsk7623E8n1+q4qpr
CLKMVcGL44nWS3MaJPHBKtDX57WQxm7p1IaaTZj1vSSlzUSfeH9apPt5oescuxcw2SL5NnrvhlxP
twchvWO/rDR5iBqbx+DT+uvEpUCI0Zu/gTXJojdAHV09y6VOzTTe+gGETNHhLP2SwK5j3RxDTyLX
DosPY+cz7FC6YCT1qIuvFrGCcexDcnTw0Mhu0nvg4wB++0GzTlfGcOHgtoOuLzwRfkNsrfSYAEFh
5ca6oSROBuiLxkn8dIsJs3PvDN4ZWz0nCYvy1mdopRv1mj3hdsg+B9dveKU/8rG+u8LKLn7KewsW
QVAGHII9M0GWYaCcTrCEChwLoE34130tr1M5t3ZKqp8GFeDnivTdx/JASruCd0+7Y2eTR2eG8Gp0
MMUPCj0RxSlOSb9K3qBKzg9eIIzxeV2iHXiGH124uYUv4zVvdM5PmAOyYKqFYvEByNTOpd1D2X5f
eeCuF2StNoV7CLmeyC6T/tJr/HeDlTjyfat5YjWZwA+r52W2Y5WA294Gu1195mHkJPUqzRdk3QiL
eI2EfKDc5A5fWV9EZwHpkBQb4buXRP43d8H8pVdNtfO1uAjcIdg4MHImHOt4hYpIw71BqIfy2x6g
9vnXUNacfMqqHTWYI/iwVghjalaWmVYTe2FZSOZypEhntwW6lzxiDL14thmYjVNW9gaml8jLICpn
VD1ooFASJzHiclINxlpWBXisTHCTUicX6EFPbKm7PnwFZETW1nIDPCPkws84AhgUy0S8aBxzI/ua
gQxN8tT2iTmUI5r+NlacFMnSQtHauMXUO2wDnMP+ibrj5QDe8mmzcKbuegkVMTwoD1K3CMzmerZN
ggpwvlbhCLsbfpNung0ExGay9gR6wnB9gY4ToPiUCCNmvDK3LoTUwPvXP5JglcKS/Pvz8b+haP0x
VJKRkxQbLHJ/gZTof8wNOzod0i0r6qOLAh/+34UsdMt2NfxCjObPwb9F9pUtjSPaE2xlYtNhPvmD
YEMKdGU0AS8XzJGnRRI3uGXgMymcPuX3VA0ufNL59v8SaQ0EYS2BxX8yxIA2DqWksrf2/HRdbcis
5QogafInANCn6ISw7LLuWuHsDbXJOf1RBFo2OzxmaSUHz8NmMGAdbLRRg8RsA3mHrkTK7OV0KCbu
M7JgCOq/CBUK8eXqCmvAPx2OV06xp1qPgZfE+DFPC05tFKOKTT/QFIFx2+X4ZH+IEO5C4iZYXR6O
KS62HuVDL4bJQG/3rRZdFgfO8uhcUkwd6E8xQHRVTq96ZRyNLCH0tw0CjMYuUqakcVObExl1EHXP
NRsLsEjz060yErMCdGswrop4p1jZb7s8Ex5a6qrmc7Le/nzM4rE+27agHWoS3lXNMIzKzwoLBlW+
5/09kzKij3qF9uf50qCS4iG+D6BwtmAAFzJ8TTcFNNbivXX/heAAN5cHk9oEI/qRJxKwvd4BgkHj
T5Nfrnga6m5bxeM5aeMgBb8UTckKYTdGaG5p/BfSHH5PLSpNtyhMhhcmTR49oN1LehER53k1FlBS
z7XYeZpCYWCKyt//ODlmQGY23oOJVE1KYQFHauvIKke6+gOLGZezFCoct6hvD/9IH6QaV2l1z2tw
mi5uY2h32/a6CZySx3Ec2AWV/aBJ9KPRXCBbkx/J/NKl+PF3kQ5UNZabykrjc0JxZNeOrlVuvuv7
y/BKycSX9S3EzIkxjDc5arsYVV2XS5aNSVbKHsGD00dllCxo0nqb6wP5BwMNOwnNhGknkS87wUI2
Mz3sqFdbqtk/LGu4p1ddRt5JbcTLwFoNlojHBYpiKmT25fXphQqO8BAGXr/TnsWUVa0aLdoxgp6c
xQHzM9TUyvlQ6mN8eTltL30QJ5/NHYsEnIF2R53JR+e/Xi3q6nbpny5EoKYddd63rfX69FM6FXk8
gMz9ryQnqvTRg4ZVE0nrP5H+jbT0E8G34hE/adJPNAlQuS61GExMiKLeC7v/HFs0l1e2dQya/m/V
ltUyI5lzUn+aayLMmoSXqEQkDpiqDU3YKScEPQ953hLOJfYz7eJNAvnHvt0xxXonL2oy047trg31
GzLPzLKDO+V3DClONNaJTLnUGSIrtb6kpkZpHmtwjOb9qu2Zww1ItLG+kyBR5JRrUXaBTXW9WdIl
/kYl2uqFT4XcX0u3EqkEFHOXDCO8MtdnHzoP1mGrPO5b+PZo5eOyG9plfYurLNEBQS9/SUW6D1zj
BhzoMRPDis7/Z9JDGlPWhLTkfpgtgAWf0KhgpGGmkcrECGLjinpDpJ/UIqi2/sjy7hjevQh4vd2A
C8FH23TcgfBB03aAAdK8h1uiQYTcjIgHzQy+PyZIz4ECbrcvWb7kwzW+8faaW1jWjVX+vIdI6qxR
pA8hMSTkJbAro69njvFvFz7nGgBbDbUZ0W40uzaBd6TmIUYxreA/0CryVeFabNKKJLn5c8GWIuhL
Czhx1PcewewCFh+BB/ANAhkNUZnfSIWmc2Sr82N7ke0hpoKDZDXxg8Ci4E86OyzksTzeG2I5rhMd
5ZcLs+RqqPwyzQc7TbItfXxpTc3mXTkThtj2ZrmMxzsIm5txEPvzVTkjNF+nhMd/uwLD2DpWwemf
L20xMJADr4bEG3wZojbuR2/zx3LUQ74Ts4j7dsV8JHaSkWnq4obiOo+5R+COwredETwkAyaQGOl3
iuWdxmv+X/xcZSGP2ZMq5AI+21YA9BOtbvZJ/Otp+FR38EIuHca42CBEp9YdOODmzIULT1ChkFzh
e7RtQeQ2YnDhRw3PnR3fcSocFLiUt484J5QXPLFdPf5Lda7PTBvJdk3GO3Ifted+W4LykQL2sWGD
xLrS+nZ8iW03SxOkNJeXL/gTVBNRL57HyI+6ANwttTI267ZITdIJD76IyduiF3j/uNPLuF/vUrMJ
v1ZsnszSEFHRJE1DQE25FAg6abk6FBF6ZLzaQqVn+rQtCDB92HjRUwu8YIiclojMrJ8E2R4+AUFE
8t82LOa276aYg1hp5t9j2rc4ux6EKXPnknlp+a/Zs5DBbWqmZh8NssXSt3WI+SZUWOW2zytRz9ai
M4YNMLsDOdQ1OUykEFHJ3j1CSLr5hWMpaUCeVi/ICKSl7c0YffZYuvDUH8g0ELtlyviQ5RWsic4V
fXV33iB+6xaKu6tvC/mbl49FMvTDiwWpDeG1DLo2RyFwQ33UrC7jSx62pWUUyMoHjPpQmDyqm61l
U52wh1hhhhl782DeOb9ziFaEhdKcoiMFEENAFTyr42+RkW085XlFY2dlzAHsOS/lxHWmWwvY5zpw
Pb9R1dLHQyhard+6Tv2Bnqj2udYNAturvSAWVzsUKKU5kEo2eSrk7cN8PA2EMLR1ArA9YKWIAphr
85bQorakxdwb3izsWeFLbfHoaXLmE0n4fOQDAX1scYOwImikTkc2Lz5ucZLTdFy9Md5HNiPF247l
Ub0yCDTb+m6+ZR1t6tXyoNMBrmoQDUrp08upt1MymQpYGmwgbKXog70QEH+tt5C0EzgV9QWFJkqR
N10Fx2Vtyy9gUzO04sEM4kaZQaIacnN7rcz1Mt+gNgc8TLsc29m5QFhjpC9PAsdEGxbCHLKhTQcL
+iJaYpG8K+ofnrOUZo8lm52wKME4in3rFS1Brdc8i/gyJ1mY+tAGxaYte9x7jNT0XMSiEHKS50rW
3OcNUZa9LfQJS/fUuPPUuaBZrhZmtFa5ODp6g/coqU3OPpbXbO3e0VRuBrQNQT8tjvJ0pmlCSGaV
9mixXBvRyeUrAhPD2Wpg1vg7aLo0bcYL8J94zU+TsO3lXwk6555WCpyJLLyqRfYLeIW8HYabJ/jH
LSegSios09A6ymkn45Syo6cQ5NsDgDAraYGKlq4Eg6cxA8/mgAm9VgveiEKCM9dY/7AsgMP93GGL
zJtIOSXkcR9+Z4QvEC3sb5gSJKtwFQdfXX75OlaMb3XtBCTtlrVJ0VZZaBlWyyD00z72I/2YwZoJ
CdLMn1G3zbt5zzdkw32NYEMeBAXS5XRW0KOHka4Duc0bUxfoInQYPWhEkt+EPFskN5UxYmWQz3eg
dPPKe88O3WcyRew3yuIok/8U8rXfOaX//QMq/VrrdsdzJWflIlYWfOYa46M7ElEuRUuVX6cZDRZq
WjXMVp29sWn6WY/bg5Iu0VzJJM4Q4c3IQWw9uqNLzPS0+C6KxUOR+S+kYLk7Me1yn5yGuaEl52cL
P6kaRM7m/hhd6HuXQQJ0v6H32AdJV10eXFx0VaYJ3MOvNu4LZFcBsHaxgz9kFl/00K+8Y3W1GXDn
3GypQXGfUJfl3JHRakVb/n3zDc4N5mOCdzIGUIjubDWHYjrzJvC/pByRgseB3RiUFItkBf1tKoRe
P4L94Tv/cqh03ca+y4m27Luc21Xo5tVdrVL+Sc0CBoRzKX4soWltB7Tk1gB3A49eAQl8tnluTWsN
NWxunaHIBsssbKoJjYHj6H+m9EQI4hoVe/V1LFmLletGKdHNEZYSpSBevAXN28dnclge5OrkT5Zq
df3SdeDkqb2LeK6g+r6WuNTUll3DT8fVVT6m9NsP01BI5C5jOMGZOTesI96c2t9MWC2pjkDemHav
6qjQ2yluCCufF5wMVSR7egwVlTOowp45Md8okzYo/M0rd3uGYqJo8p+YtuNdSbUwLCMY/yUTZSTr
S2Rs8GYdyceBxLUT/vEBh5qUhFa9toVinIWLFwaw3O4qr0DBouwFxSl8FFiRDbKp0/85L9qH8rwN
JzpCCF6lrfN5V+fnOvZbvGMi+2AMCseeSiMhT7H3n/SJDXokWAg0eOtN23n9A7wtINeNOsFeWHYJ
4SlNNrrP0iVqAxowK5mylNKgF6LeYvS/+l9wqjL2HHLLsEs3IZB+1pm++JV6TZZqY+nwDLvMyrtl
Vduz20fI9KN48fDFIHRQrty2FQlNVMXP4pEcC3Qup3CoSMWeGkcrgHtafdqFefPKaJprz949MUam
Z1grCT+3eDY6+SuoROF8gUGWbqJmXwWrxQC6lnOOVzfMYxYsAttP3W4/KyERPFyoYRIQ+EokOrkM
FMFnEkc6Y38z2/kmbFGgY38mzT1ccmSJRoNE0q7xKes6s1YXRFz6FJAgfh8tvYSPVohDATxh3oa1
yTzsaEOvnb9tRzzN39uv4ZePkClBx83QEJIq7f9rRvs5nf5Q8zieRNzE/cwdWIRwopBv9k30ybQl
AMTOhEZwcfLxX5hfzCceBhQLps0vP02L8TE17MuZFzgLKCSDFG2GT85qM4EA3s2VwrGlChR/jN62
unX+kP5UsND4f4MIJkAm8pRDh3wHXZr0QvIRwzVz6XKEFw3N3Ct0Cdzg00l6Csy0Eu4Y/gGiB23D
0GEqtI64qWig+/QOclIxypiMEcZ+9WBi0pGlKe5eEnUFnR0HQZ3bA5RTxwgm6ZQdUL8q2solmW5f
8jMYf7VBwSaABZXv8ZPofWRxwCrdYQBEh+Pa1wkW5wdxM2R9hXdcMcoe5NHq4hg0QbJjxnV1k4Lx
3m1VyEA58qd7ciP87UNKLEzYwMj0JElbq78vYBwIV2BJPRrh8SzoXjjSSy+w5R5dOFEX3fqqPOzR
qk7nGjgpPyoKa1mb1OcdIyCRPxwWndyFAyLNseUhxpzjNATEzuno/hj+GKS2XVO2iP0sdE6HQT9m
1lMnfH8lZ/mbYve25MI2lP5IG22f3ARh+DfFPhxcBCfogCqLBHdHhiqxDCRRxjMUXxaYU7eMCxll
mor3VWEdb0i0rPS3X6vMl20SahIuKm4lPrdKBLAWGVOmwyYqHpBJ6beTa3BLeGl4MGmU9Cgjpp2j
GWCuwKmH/EcFSYxHcABL0J+TqMKqAsD+fvyijuj5aRsT6n/4J3q470Yw8cjcyQvUaYK6CdFZYh72
iUEDZin+NgAfF2e9yOZFj26DH3KkKmdGnKnlH7MOBc/Rujn4HTePiwPDgq3ruTZNjb+3XkVbBJ2e
v5RQjSkKxCE7CIVuBDILpaRx+hiyAJl+n2+46RNduBw26T8Oykb7R6HtnZRHnwUaVu1cZInrPdK0
zPRhsATDoQ8LnLejSGcG9fBFLVN8p7EMlOWqSG6dFwKLyB4n3GXuutuVfO7q01ZhmeTA8cJTArFS
mvkHKgS3zUX5C27at3HWbZiEBFXJPLQQfhSlJsNtcvyk5E8G4ALaSLrtSpB1fnaYhT0rJ8ZRQYOn
CKoKuqYEJfzKH7so+/tG6glCUtoOP75GlglehP7xMWqaFbfBALV4A1wN9L0jIyoOXMYinRSIE6on
J1OFufakk9OCGYksPXeQbN4TyvB1Uq5HPMMAgZgQVulpNrqsW/i31vFoCGlDRncjmkRZt9SXWF7R
SWrS7y5y4HLf7u4MnOpT6funZsVZQs4UCUyJh86+0xsmoxvvgic3OZ9kObcI2zHi+3aSuatjyYR9
jNvCYyebvHO/iLrcdvnbk86m7RWCjI615yZ6cu8xyn0NVur/xK1e4CqhvfP+l77WhIWFHOfGdHut
VADw2bhQo5FA/b13qaVl3d1NXQmGEPSp0T4RJCdRQ5AOqRDIt+iFD8Su8mjsS52e5VnCNUYKFoGq
BoibV3+hI6Q9FM0IfUjlB3Um2zBKyx0LP343EXeLHpQbp4uGS2nPy/FhEm1DELNyF2Oph1nhGFXp
8LHjCFx0KAFcinVmcFaVKqdpbcWSXVIbUynjf3E/wdomAOlOB9CfScnH877C13PcIwwjCD5fyRnR
YZigqyz/A0xbbBm+RT4yvCKI/LtnBvqliNLYW6V19aKA852+VD3NZggYWDc52Nq5MtAES5qcLgSd
02xY7Vo27dq22tYXIXCoHi0YOwCMnG+PHsf2idJ/rVpm8naIObEbJJ646n8W06Pco2+8zJsyQ5kH
mGow7Qj+F/RgVtNc3kDPpDrcxoNP2cLyxzCwjFeSMsUoOBJ4fVx75sVEU0JzRDEqu8ySUL3qSpv1
XtGITf8EphAFXAX4qQxgb+aj+BQ2MHC4l/HUkkvENe3GcMWEN9mai04UWZkcx1KJZhgBoyWEhr4y
gqJngNJkditrudqAcfay/AnU+goH2nkv3sPJiK+pRYQsRMqIsuFCwZ1anQZlQLZaU9gI34Lwxcez
eLTtvEh8s/LN2GEbs4nnDV1Nxbcs1fmAF63Vr6mRFS5Vx5NVDRAbyJgh4wnYme9U+p1UMGKWQmvi
RpBXP1owsZB0KMrIXnF1xv/vmOY7bPZzubr6SUGFw7lvmy1fhLhFuyyeTuUkJG0D7qe1H0BndsQ+
m1eDhP9LQiE722vT9mv0UteTMP7SInSh1j4vO8gFN6fFPv7xm4s5AshAhlbq7qPFK0FeBgZj0vAe
VEhQY8+l9nfr0f8gqFmAs6QRCTsD8/FdPPWNa86ctQCn+EXouniANm24Nf+mXwZxkWc6vYYzrgpT
R/RHpBNT4KxedsudNF+253UIes+0f6n8rivjgxNb2PWYFPD8ysR6rmMylBfQAXUt+9Qm2ol7i2Vd
BPjoWAG65ZpUZ+sknQ6I5bjRaDJUrlnNf/IKiY0REWP+ukGM2GjRLehGkXE0AbjY4+2nLXkQgiV5
4PcmiCW5Ndp4cNfa94/You5OHDMbbylF/17lpBVvZet7UCyHmO2NSCUmKrZ27RhCRLyMH+s04FB8
TFESXQh0arunMAtdPmqXvpMSMW+4ZR3mr+tgpM7562yTiS3bbOvIDQ7eOPT/8JgA58oCG7vRNB8J
OT7sYqPNxOlh1W20bLEOyxPT/LsOF4PxYOYH69gpzHwTztV84oj8bGs1RwzQ+pdXJXaVsbHqMSeM
fsybm+MRhkA3A0PpqAHfO2Yz5HwOrmfhI59KKd+TLiwqEUglqEFyYJz1c+Ifm6Nhg/mvE2jVcbiq
6UuR+Lveq1aiSfDiCwuTt0i6+YS1yKFGnWs2r6T2G2A/FiRF6O2hh2DJglmzu+H50jhBsdRqZf7A
tuCzRfGaIytNMUAdEgHU6wLJSpnhSexG3dpNJpQPqiXFQfCagNwam6Q1iDquprT1qObeD7EPHSvi
0y/CB5NEUbGo1ICD5yNBMz6s1on5f6ziJHPr2+3BRGigp3LFoS2aRLfO0rJAMEbPxZ6HMFo3I/Uj
I8YmVm+CYKu1pxoKxdPcC8MjR3L3jxwjcHY4RvNbmMr7u0w5JDFSlrcjw+JJfHVOT9n1swsEp1bD
hzhd+AM3uA7Fid9xMbBEDTqStVOWkbCoEFRPivwTQtp2ft/zLKg/e7jaCn8HQab7bknglzpC8WDV
Ud/NDz45KkNtDJPKzIL6E2hRPpECy1vnDbzahADycDuSUmFffPVxZz3QEBMjeGEEmFVNrzVl4Xtk
t9cp9qHQ8BzR6z+kngM88+MnYxk230fuH9kSiQDfR2UcRQKoWPFuGbFY8IKFHZdTcQb1y5OatUDg
IXnA91ovo3cCTeCZuCsINmZX+Ebzr2DMkIovNADeo2yJAU3LTx8wnoJHxGdCVr6owmFBgjVQBHZI
1zAjzLe177zngwJ+tL024YTkQ2LB5hQEBH3oH/tMgfsqBTd5mRewyfVtD5DM5puwr4hHWUg+edmD
gZU5KieSgsHQ8SHXLbz3+F1GrijBsArCx9ykDoHQVPqfbT8CvK7BfRtQzBP3mbnewFrKjnBUNgvG
I80tR2m1/osAhCR+0aEysLVQXksMh+vPNOA+cbj5bBpw/WT47e1pMYO+VFZQVEmQSJ5CRLXvNs1W
ZatDJvYDSz1qxbVQjNc8HICa5dqlyBIlpBp7kxWOArLRzIYdrDtLPU43zuFBOi5TMaVI0ogjJxNe
POr0tGx8ICiuEQAqErk4Na0ljoqYIFCLvF0xhFQd3Q+vxjhLRrYm2cK7cXL8Xg/GmmsgaFeso23/
BjiWNJsJ+/m+vZIVym8u8STVbStRSxck/81jV0eLQJri8YG1xoY1tCk8oXFtsoha83Vy/aRR10im
5hdVFdqbDYeOK27vkWoI7mSCYe4/CFkClK6n81jT6Ax521hL+oW6c5Be5XcOjzA9YKxTbyA6MjEE
hMbC8LsEDdGq9R5fmdZFmtXX/49hW0bSdxTCWyA9OwkXpyc68x2kaVSKzKusMDl1xt9Iwet6htKQ
seb1gJMH8QvlbKZZRuA7MoJ2CiznwowAR6bGA+AYHlIGVAeGhA80N+Ceenh28a3vFztzw1ZCtvKr
U9Ofm1NO9fV7M2WHRMrbkFKeSHXUU3pB8VePaqjOroxaTA+SOugIXHHASR030BG9t/08NdWL4G4t
Ibx2EGqSwWaA/GtqcWBgSIRvhkud5+3mrQbVkAdOyEqdSU9M430r2367sBjWjx7ad0YoJ4KUsiOY
UyF0vh2eFjjQFIQ1mBxv1z5lR+IVtzwkmQMXoD2M3XkdJAMVFWXiinHtamKZLnAHmLPoh5Fip4sl
SuYEbI8DetPAD5fjX0VoP553yqjQvk+ye7tBV36+lZ1sY+e1e4JvrqDGivNtgGaZm3+wFfRxA9TR
9BKL4YYQ6DWHnaZkiYMD9lc3tMVNB9qkXBwlB/9HUR5IVkjbCeaKhvSu+2TJ9DAJZRZvKYXuQ6JK
OFKk02aIKsFRf8XmunyViduIRCopb3idPjMMrm+nNas0pEYlqL76JgxznBcgEFyKwqcbbragNBcT
kzhoGxcQjHuogFH6RwJDBgHw/Zume2wNWA8UA7ZVwWYzFJOvTVpmu9iHjR9t7EIOEEPz7IofXWIv
qMR6pXw6oue7dOZ/TcsjverefKcZYWfV/WYPjwfiRSiTKclvDdAENO5H7pyoABMR8wT2464nUsPH
dlPJfEhZKbJAS00wXO++4Ao7jlvcb7/CnAaZPqcX2cG4lDKHpAY/6Mq3bZ/X+WBspI3M0dyskAGM
hBfL3k9SxHVQuun6WrKD5/tchNG0XSi0YhocsSa8Zs7OOz+t4Xr0kE6eaGaEZPcYm8EHwRtPmhW6
JUYcyTah4x+Bt4cScxBjfhmzP1gJ5pUh5ggfnkWOs+H2JVhZzs6i7z04+hYbxNxcPziR/JHdO8fv
Tpr/nkoKmtgyDQ5tv7UtlW972TSM/cPC3hZvBXvC5qsorv9bXGp9M6bUagTHoTtF1RJdJQMqDDEO
56yvMtJPEJXcvZaykuoqhFytyTPsXjbmP4m+C55egsSFiT4jhBgPjwOdnb+ir119wtR/v/fnQaqN
FOpYubVufTYsO2KiC+xYbqEda3sPS51iJfYPtZhIAU+ZgFrWpuQo124aFw3ynX2MX5hYTnnoeIPH
+YHGyCofn+7FhaP/zPRJgsmDR82O0H+m0NP+DN8X1erY51Oo7I5TmHUJA23/Qwe4yXpSiLyqF7rk
qWdF5DmlcnyC9PSMvr2oJ1X6hhQim6oWxOXu51ooDWQOD5TPHXpOh82cVwc+xiiODfPLggCKrrx/
BAZjsElgnwtMD2WBexhwxiJ6gf2sVzEiCGt441vrPKypTTn1xeIHcFCeuwzSFfTsZilMXjS33VY2
YLGl3Ie20HHsg/AwBLT0KK15kodpMqrr3alHm6kJyW0Y0IC0B+1J2hm2CW0T8jRAsEsf8kIAaEhE
dvay7AsZGLQx3rjn4VPGnfuiabXNk4a6kkARIgB1HTxNkmOtM6sQUjs67kbaRxUz63eL8/EnYWvJ
+dorGjsCOpKaa0vU62ckTQm5N0sUlArgvPo+YEAkM/2c0qxsvhnkrGGswCHSVB+9pSffJQtqxr/T
Wuvh73a9g8m4BA4sOyKZ6ltpZBnOf12QfLCd/CmyDGupMwCFN7qr05aq8RtEyzH9xkjmbQtsxlW6
8R7dixyRGstJP9nZUYQR1XQbtjtYB91vuH29MqgAQ6ukRhWmJJkLkO5YYJ3VvLFPAMz0dEgpbS2D
crXLLuFHDGzrUkIPUaw0CgWVjvA1FiyHgVwMbEQOo/qyDkVlQnJZOSHGMI5SkDCPgsKEt8bQomj4
5a2cOc32zoEapjxI24K6Mw+mnokeA3Cfvzm/nKFlu0BvUsU1csZwyryJrXPrdB+X2+hcnkWAOkAq
Vg396vEVicCkPGYTPSv8k4TRUXZ9zOxak1qN4xK3K7bp3QWEHwEBEid/EUVzHIW8s3TPJAmMAsfJ
JJh9DTX/KceOHYsArGxD5bAcIoi+K7edwRVvNlHmQPtj+5WCD0t5KYiFbR1C7oceS1iMCzTQodZi
hT7uqmc4DKOdRPDfun7yIQGi+GNidL6zs9Qpxrhu14hYBFKSsfzVcKVWh2VROKk/dWT0swUNOdAu
ncRsN0rWmvnpLNm9a4TlGdPynXzr0FRXEXhxbruNGMS3AToFTq9u90PrQM3pspWsyWa4btqWQxt6
2RvySmCPwELtkKWWz5PBLhpf/pxKFEod4qbTtzE8/nwYpgn8MGMOjo/ry4bJ5TRZ94XmZeCsxUj7
YF3ifGx9He2lSAoSL8Nu1cVRA30DSiw6Lvs2B9PQbwqnvNv0/SC9mnw4T/roH6yZKvJ7/J1uUieQ
2RYtxR/YX2aWORog2BOJVKdwCA1sbkiYSyzq9Mno+Rh5FGXXcYDgdVOpSOfbu/9FYssmlWYj9qKj
z6s/27PgIT16P970mFitsG0IPMzroxqAyyMXuyIwczqSNO4e2bXolu8+57ib9p9i82kNyE3VDt57
z/nSC06D0g4KhJ76vaWCKRvp+MkGT53Q/h2XeEYfLZb7rikSlY4yE5K/L9+QCzpiE/OEGcvkvlTK
52vX5csj3jP51FUtocsXEVpNFgnTV5NsPp2EiEUDszP5rGdxmO7Pm5f69br7tAN759PZcZ2lUs5g
mh6wOkdLYqMypMq1rOCI5bEt60uAY9Q88/OYNlZ4aPI4gsmJLbDVW33ZxehOVITL2xEdbKKrzwom
1D+vSM2bNqcWva6+u7cLV4ysMjNJrqMEEymhmFasSOQ2nmTQl/lIQP8O57Puy76CqcSPX57YAqq+
Y8+hYXtpHTdSI9HklfHfiGHV4tTcJQ5QQVPEFiUSrFWPonefe0dTB6W4bFVczrFfrSYQLcqk7Dbu
IRTfUdSYG6pv4XBkMmZq8mC8Jwek8WE3ijEHHJ5SL6SEaYWIp8d6AdJ0nUGyAOBoujCu9J6PJp3r
qr+tacyby0JPCixlZ4NkOn+DeSZAdQutZR26l/LcFtjVgLFcUTMGDPj0lPdcPD9sUDX5RFMHL1SX
87fK7ZE5yngRtSDm5nBl+svhdgXxchzrnEfgrIhBqz1q+CSyItT3YguAV8qHK0goCj7dEjVK0M72
n89oUSi8H0dE4a06Jt8nPcgA1BOLzkauN/diY2X5T9vvh9ETWP8oFXd5nJ3MXSDFRfV2H0V+NRfs
8BquO5rY1vYNi+68hvLuKoA8c8G88M2diNkJeSejhkKDAUu6ieVIAbazeQQTNp3K3YyVf8hBdcYv
OCyMMDkF/2Ab93YdQ+M3P4IQ4xADJMPqkkHLLTzJmqISSF12XEJaS90NH+PX2i+fOmZClOOY0BGf
pDul/7Ii8Q3rL2FfFcyt9M9plT9/b/47PgFJ9JXXLkPapKhzqBa3hWRXd0cOynSrvYeVwssW8bWi
I13/CkScjaRNpbLLediIyL98UreH8adGZEWqT3eu7dF60anUaw9KleUmo3btrtbmxYRbpev/Iz6U
cZ6CoDrg5uhn++3RrmPWEoYdc5T00c63U9j0PIeQrcFPDEz4OUivB37EkM3/Sxbnw7fd3xc3M/Ru
450kuKuV1hSsXYrIQtLCUiCKc8K+U/wjt3GoUVKnnVlFm4oP+iFo1aRKaPJxuPp9GwahbybbFCLG
4GifEGkx8s9Y/KEn12fZxZF2YZf6Kxrw+0UDvSBOsQRmTQxUGtpNI8Wuqec2HeuisKrGpe2P5dck
xy3/C1DUxxRCuk+r+QrnjMXdz8gVMSzGz2KBse2mSUNWO4l/CiVfGZ3PG5WvSDBvF+TNPyBDrJA4
+2qab5cNspAoXv8sfFCsEmcWuFE3bB6ms9YLTeTeglHDvuBcq0wUrmqy5fP0Vq8WfukQ+hJUioWz
e0BtOYsdjNXsDUwYdxcSmKEMVa7RzPif1hBVX6F3NCVK/SJcyrqH8fXgEkOVRYxFf2IB5/agDJeC
wfJNacN8YzetVpQrHMthAsjTEEzB0ZL1eh5RdBKIUd2LTX5DuU78YAmBdqaQYf8lBXzXwWqMRhJI
1nhoj74J3QDTn5b2IfxSHgXl+fUWkZykITovFnyjVvIsGxCwP3JH1p6LZlXsHj+CR7F4ywmVo/96
c8tuuH8LXzMeMESXh0RRRVfsMxV286a+xgBm5ByqB6TwHvZH30+LuQuNLOYzzEP8tawA5PI+yfGI
HognbXgKOwTMSLQz8zAJrHRrvWXT4y36e6Gndf07wfRkZCFiW6YHsqWiIWefyQv4vXWsLex4vQsS
D1GILsiT91yEsdpiYGQlLKWVGSzw6hJnXt/l3s7WI+P7LlIXyT+B1/C3QnQQSoJ5b/k8Mmkkl+/R
nbQniS0ck1Bl+Rz9IK4Vrfu3CTl8pHTP1t6NJKCE2YbfyMuzrefXTAGrYI/T/YvBMiMzgAWH3M+O
NsxPGn/J8WEBwk2F9hOoI96sk2cD1xI9sIQcNdxSGzbulw3mvPD06dBpm99ng/l+gULHHXhc0vhn
eSBWe+d88wRjQaqkQ8VGUzZbUXLYig+4YVIH2WxxOt+XtRvw+IKkUKlCEl9gTNddmASDL84Mr7Er
aHAQamKEpNDVqk0FZS21kuvw+YGJ0axtojnuJQQPJ5CjiLgvHi5O+ZyGZpbORHBdZ2D4tufLvrot
BgPXaQL9CAE1z3EBx5DpY0ZrNt1q80N2CSrULr0oHkM8teGY6kYU8znq9v3GYKAnnJgh9o9sUWYZ
kaj/y4O7PyHDcixJXPkHrz1HIykbettR1CnDYCSlxLs4UhgnQ/HuwC9TwqGro3iyQNz8uZtpDSIG
3ARR1W07muaFA1ZWc6J6K9g6H09toPEKeHl/7RmtzCJPK5Zonm7TZK8TD8o1KNH5eBF/fkMixnJp
+GTUoKAz4d3lWS8rJpDpLfs6a8q7y+9coQAv++FWak8zjM2DwVfhjfKv7nO6c60TLarq2H8Jm+nB
Jz5b757dYaZVRVbpAqGK8GGDBIaIc7xA7HM9FpjSgStP1UBAOMAU/xfwRaI4qHFTqaTeqCQH0iYA
eP95HLOv4+1HxM/LtHDHpLyumgUkcM82QdTIfNQmurS0hZ2y/O3ffbAC6QeewhM4RyWzxLSJfrg8
bgQECoiGjffDX0uD02OfUGsJK1Tw8euGNa5EgQZxVHAH7a6WBMVGqewIcQYGX0laIX32DV9nMbJq
pDiyttrGLKSnm/9BTp8PritRHA3GCWMlJHmJSFx73GRK3b1fPxUthORZUa4sPSLjgwRJIXzwmheB
/Z0LHun4c+8jv9cu78jVSnGrXZIlMF3qsDm5pmsSMq/RMvnyrLzeZlA75mJ55qb59L4Rx+0sm1AC
jqM5FeURZl6dhnyPNcUiT6Bu8nT6R6ojzYMwDkQ9g9Jr1rqiIRbYYKA1Idmcrvfsmm2B8wLzB3Zm
c3R//YLbJ9sY71YPnJ9ariO2OEt0SVTr23mzge2DZBR37v2goPShXjTxUVhxrjd1IreTIKhsP8V7
UJchYslTma9lfQJZGlGNJ0oKKl7kpdCaDqeuRK9GSgZIl46SCvuKJ/wcfYYozepuYe2OPdAjyjJT
aYSIDYPI+w1Q5Na6gNrl206Ij3V2tI3gbxXucB2P7TDBmSHMd64PTwWW77H52g/WC1irs+RqY9vU
y8Z2E9mylJ4wcJ9V6ZhqN6GgNNzheTni3qQHHM/6OeN76sV2eC+UhyyllwwmubmfvgLk0JTMnJQR
DQv5Dsju7K4jRxlpkE6XzGBadoCLdnyhC16nMUwU6ULSAisb4VIFgsZTck17jC4BHdRZok/jE2D2
aLc0/f3CVUBz2RolDC1ut/HsiRIain+Fh8fuiirDZAMnyIRUvjZMabOKemTSCy4dvMGW2WTzvgOo
89sIGEHk8Wz1gHLCnjnmTRcddC+HrSbVBveAyiiYXqBhNvUe090xZ5rt8W043Qln55SycOVzGFRl
WvGrWMAf9MaWVMhCck5kktRHbQQWQ/V0ZuHkj3Gr+BqrZQdUTzPKLVzR8c1esk9HZvIzgV4a5d3x
POtdXcgXAhW4JIuZiF4Z+iv0Vg/2FglLxXcT3T2me2LSCWsYMpxYrl6mGVXlgxULLUr4zEvTNpGW
EMa5hIy+hsn/3liuI2OaWVHosnbk3dDI1WBsg5OhieILgUmHV9V8UlOUE8yk4gPEW47ps36jc5B6
uJ5PJ/Rn77JE0LXI6jP1EUuNJBWBh0uqd4CpR7MnCMXLtuYZtOHkEgjsWj160B+mwpbREppwOq23
8MLEbB7GtX2QE/J8oqYeYzCFM7XuMhWFCbRanH+rmLqfszkOvbTbJ5/Yw9WUSUk5nAJ9y2zCVDeU
A4+21q9As27VXw1JnuDZ7bV6roIDHoZ9Rqt38xAyz0tUX4FUbUph/sjwrIFuTzBvqoWGepn7OlKb
v76oZoLu/816AYWLBCR18V4jTE4ROImQZvQc2is2Z1sXKhGUKqj1M27kyrIrve16mu0DxuFbfhnk
fU48/0T0XR7jo97WYFzj4U7pSBRbwVbNd9mqGWEgxbOW8WFdTBdmS7puJo93iWHT4dE6SIsXJUxf
qIIYNeyYRSaH6EOfBEzD7YtIxoBb5BT41WfdC4jUI5G6HBHI3MIeU5puZYZigJ5R9tRN/RWgwZlQ
hvH/XeKfKXP8zvoK3Atxd6Yr/kz4PYD0qOSRKRudJFEChL2GA9YpwPMANVFDAvPcsywgpztOlaYP
E3g7HgfJHNZuUKz7OHxfOuYbJxTrZqef79LMtwHZvcjx5Z3OI/NnS5SGvp9hdRaATXnQhapZsD1o
cISQT+7vHqGOr9LRkbqfSy+vVM3YyDIjUWJLwZgRsAex6XTDG07Yw/ksZeymDwxolQnvepn4O+WL
jNclxiNL2vV3RDjvxsq9t/xe6OTUX8LkVQsph7Pra66u44cC4LXobnaU2C9/m+LfE3uTN1ue1rlG
d+aFT22No5ZitHs86JBdUAPl+1L5pI3kgLan1DzTgziucB13kEry36QHKkadfLy2Avj3+uyS+5Tj
+bqmrHHH38E1vh4SYLsUDWrCkOSKKxx3x0I6n8cW8f3S3lEikZbbjMLgLc+rasvxpX4XxnQ+oa9e
sEBgUMCwHgH2xu3UnZI0lV28Fw0Ihpo2RHQhZ6mD0FBS49QVdFIEtZvHMRvlW79MlH0gEMtpORab
cG59kBV9ViGRa2gYwkWknVxGjZ0TASbrsJs6MEhqltnkY09vfSPmbBx1y+gj+y6JRdoey7k3T7MV
C9Wf+uI9CR9/asZe1hxVEt5SAgCEb4tJVcwUK8w5uB1EYuLz2/0V9cVPmQQL0Xazztq+50A1wPgn
CxiKCGE4oAzBQMa/UMVqa/0WMEVgMUWigzAKO4rYLPh5CJdEKJSEAqFz80TsSjv+VoHMOIHpjx07
u5KPqgg2znPR5eWq/I//nlnMZqomjnfpUgxmqmwTvzZVGF4Ff5QGBD0YKyn7X9uDI9KRatyk7xQN
f8RjbyZaehcaZC6+yFn8vf4ROWRSAeqwO5sUodNgjXxW9tcxsbRnVV26Dw63+n5E+mIwyvFyfpXh
xnngnAxzvvAJiOn2Utb72jo55HBqdwvhjCdVnV0EP3m+7L5CPW2R00Dftv00+asjrpyfkJxCfstl
+nix2Rk0pFrnCbkPB65xM4TMMcVNZWfPloaL8ghDVMK+zbWeR4ZFW4xrHwLNUEJU0cQg8eIbYpr4
pMT1GjkRpDyhilA2lk7UOYGjwFensDhvKG/ecoh+V2xPItK7A4d39YEYe9jgA8W3O7nuK5dAl6rt
aIU3nhJ65t6QCmT8WB5bQyRjWE7jmX24wx74Tmv7NuYp+jmYVOF+9N+OaWjof++ihfxYzE0/Le7L
2MFu8Pszp9Eqe+3ph4vXyxMXSjzYXYnP2I11ZWgOvxbNqw7WG9aU4npWZDO5/yHtILFLa6UWP/ll
K2oEI3pbgbd10PL88njj/0pGD7b1/uHL8ULI5U1cI+3VrimIF2TXn0oqc7ypck0ZsZrjOn/QeWG0
gpl85gaqu9K2AGYxY94k9QlIPEfxUE5o95Dqyd2CnxXc0xXvWIiwrUPU0y8WVouKcAxXuzlu0ZvZ
Nxa8oOYBlQ5WP0cNtonztBhTbyFsveYcmLyMAYT9dIa9hLYJzfrNnzGRmkLhwDfibz1uNP5RgJyN
NIMPaXU6gYK4ak8QnW/R6Xig8DHhmznLzZOIYFWJRbuzfc9PDFzEyEB0Efmm0PulDCyu2n5WgIYV
zY46DNwqP5w/AOGtARW33E1jqLMdMdCBJFxLL9oyLh1Dsbqa08x8XsprfLRkiGxDBCdYnE1j5Our
HrmivDYrVwiMy5X5rmTou17kzlvVA9fQadI+GSP7kTewrFhYdtL5vufZtD9fF039PRcMD+oyHdN4
lP1GvNMXZDvQluFA30btrRFs7DL3cdCwr9XrBn5i8EVeJRDynsHdtKxdrdJ/bAOGMEMSrmpYF5VW
GjRdqW6y8fsQ4wItpqLp/Z965rIJ9TAHJw5I+6fgN0hKFpVLbmtQaBVP95ACjEx5gvCaGV/B4XRN
oBs8Vkbp4djJvG8NowAoYaYArt6h96LBU4hWD3moGG/v5dPy4mBc9HpHrMIX0DxmQOWBRG4+DfrL
fIAmpivAKs1s34hvlSFqQXkcS7nLcfFSyuGHK0HlNYIl2baHT+6oO8GTB7/4Z2ityL2/E9MaO42p
+NThgenbmBRmeCgKtGLYMtOzlRQegNHsn5ThLate+tuPxEzyDlNuY84GR0lxBfEwjSBzX1y2Je24
O9NLGVPSrKi3z2QE88xGagB3f1ZBlV8HAduTPBFymWQDtTFfIV3rPQ2ACX+lFmx1b/TxpiqY692s
oD6616wfPsPG/KqGOpLamjHqEim6sOZuC5wQwOinjv6pTLcFSJCZ60hUZ0F4g2e7XzR/FCE3MNc8
Iqyw3fSTUCI+KY8wo+zD7/6wP6i5k4L9BDFhH2iGFXIMaNHp+tSTmWOIlcJTtyPrkklgiMqz+GgW
Ic9N3vSdp2iEYyxzbOXc3FzuJyHJWcmsiY/ruBvbyzYB2eMD8H9YA3O4aGvirGzDwV+ryU3qa8X5
qMjUd13QQj6f2jwc1Xu1jQAUpJH0y/7D/ti01rMVnHY8Tj8ydLWWSElby9lA+V9jyJDWsVwjjL/K
rLbnZ6MhidK81XdDIDA9Zr9jVUA3Z+o5sPL8y2rcQySMHaH7WsArdWBw7vPAM2wfHDJr6nJW9i/f
iMyeg9yE8GpBREQrGJ4TIxinIViCYY1QFv1REZ3NYJcSFxc7yYIWBRj/fMN+Y9LKjM9/DkF/5hjl
qwD/P1+mxniRqFossbK6FUAXPk02PCsUm+Q5wgOHSEFim2+8JG/yA0JgGzzY7LH/2Nk/PCC71vmB
4eACEZzFDRxu0p4x7roM7aG153A69JtYxs8uIKfgWNYsSVbZQTR/T7gcS9laqnnQXLJ7K7fBoBcA
2X8s3D5TTxu9Jf55GSppr5wiqFIJEGHWO78Xqw11/iAUcvcneFTvZJONw1MScWNA+PQ5H34phcAz
/dGCiF9cacwiBoxCRcdDgIAHGG7p9TqSJHwpShxCFBkXNSZOVt3hZ+cfUoXgp7Fzqn1XGqGhDb6v
fsFTdKNRT1m51dhF/b6hdyXOfYyjTtjGTRRWUNdWOs/fD7wIk822zQmFfJcAa3wWND1x1oCbrLRy
rEf+GRtu7/cjeqMp/7iXApnvexErwqRH8+ZmPBermot/PbLGsXFuEmwZKrrs8BgTlnwEw7SwsUwi
YluGejeejgQzpMjxj1o0+11kERPCOIURx2jNNqavpne43X+9gOeDusutNrBkTbhndO/47icsAGef
Z+0bJwTEmEie6oMJgpCic4oACbrCVe2dk6thEzSt6FKmNWGmrePThtGT6EFwcnoUawIKhaeKKcme
9Lz0LhV/2y402zRavIUhnJk4owZBQOMmulBFHhelnxkOtz+7Zy9zsmFnsxbg56lVZbTVowqZPPPU
PLSwimm2Jx1WVWu/OoBQvqEMVwwxOKo+CLFf8EBBoyT5DEdOwJ0FceBBHGOjSHDEWdwScNkvJ0F+
+UAoKMyuA8zaganjgL4ImGskknBjef2GaO76TLeAqZzyZNRbUDtFufT/TaRIPLsKnJx8kX2Hntwm
RI74cTbPRDLZ3FnNIPrUfUAocMYGLNrgSJkem/2/1qOSzg5Uzzse5s7YLCn+Fx8v2zgYJxCBpJNb
nOmANAZhjC0olX/JvAFkODJT8Bjozg22vQKD3WZLcVXJXn4hQswIm06/lkXwBJM2DtjD3Ltdy4WQ
yEjDl+9im2jY0V60nnmKaLPKv1JGOuGOAa0v0AozDAKEkS4+tAn98XpwGQBcP27972ntkeL3c/Er
QnKB3G9/onXecxV1OblZZ61P+LBu9ulzHDXieT0ST/VpFQWydr9RMMZsc6eg0l7ZLDzxvliF3dtN
w9zl+bZ094jkNMWQNhNjvEDPV0Klk3qaO/ia+IBPUcJXarRNe4ztOPwZ7NFFkxgu40oAgMHz89Qo
u9ZrSVGSCW79Ua8vWhIzfqykUg2mT0Fcs2r606FgBPT/Y/5ZktQEKJc1a0StObznU1clAC1LCxAu
Ti16s4IOe/j/VQoCe3c8O1uv8m8tV057d2QyBErF+GJZOCYlL3cjp1rnXN9sxWnObo3cus5Jz02w
LuuRicUWpXXiDotbehhTmN1FkSDIbmc1a04MZJbkMYt54GNr+e0Yfe7nHnpncjp54kL8ktA2BYoD
WO218sZuQh79zTgHGdW4gQm2I0TSIKcGAHcGOiBnOt5qYhp/QvoDlCCcEnWFoqS+2hxWwn/5Njp/
MZhy80agl2sPytArXvaIwgOg7+M9WxBrfqMbLn48Txf7/9p/8pi2f90H2GE1qHGcK8PlDB1b5X1k
G4ZBNQKVpjDZX4qCB5C+M0ZYSSFH5hxl9UOlMXLQKR/4+WmW4Z5+kmmgjuH2f9dm8z7R6GJDMjWQ
0Z61qvfcxaD64BE+ApyzGK4ssnU46rGrmtp/0q6g4V4K4x/eQUnLkErWOH7zM0GjVgAmtxuK7po7
PiELzOAS/7xSXYQJg4TPi4eIiztNB7DvZZjGM1Fm6iGXfsxHkcBgafJnExDBtqpSG9Yxn7J39J93
E9OiJWYyr85urOEbU59G+ZedPGPFd3J1WTfFrsMCHGNL6VjR+J17p/LO+EErPznhwRYdVjkJ0+bT
1HpZDqRLq6hSGoCUn7+Z02Sf8QSCy5nH8GX5tHhZj/BfcJ5NkqjzFnDZBan7jq+JUvj9jFCj2jW9
PzlDMBjaO2nHPHErdqJdCz7WwFjlsW2XmnVE91jQ3x5IYFJu0/aNIyaLOpNynU3JqsgGpAUzhifV
yRWknYONEgSeEQOSOpoI2Z81+tbpy44EemWKz6BNw96PX0yvOGWY25ghJKtoZK0hJSzILfNWYsZo
YAMg10XRlg6jqsCvNexqLSvzn6XmUGLHBcsxtUreJ4KjLqbhtV8M2HVbi9aECr95ATBeph6mouPW
XTQcEGtl9+FDxVs0xeZALbrqogRY53ExURSCdcFGdfXJLAae3q+EJNCT/huOT+otWC7aBMIFdY+s
355RsdlG9vp7dA2qqCzg3BEUGceQiPyqRQ2/GVycWVs+6zf6HlpNMvp9G2I0gYw8XqNSshbGuAFF
vTI9hrnkGPLtQTfrJ+Fy4rrHbZFY13Ekujrs5NLaQ2zszzpEFzEXV5oHK4NfvKo2BYifWq4KMt5A
No1YfheyL85nuRQjJTC8EA+iz9FXQ0uWsnBp7//s5MiL3vPqKMekOx+1gudMyXOmisN2um9xzb5q
T6uiOVjUl68/2/0ucccd8byYxL226Qt4XVbl0jAl2NoCFICHyM1teehsUCZUwwOyxs9rlsxA7rN1
xw+WJSwNuzIN7xFLN2ZNE0tskvrIHkL+SxrllPWQ/nkCAShd/VH+Sn3gjgcWMnbpBNgmO/VLl/iA
cVN+CP9DHrQ82wAGfprOGmK6Y+ODXsh22qF77e9nB7rpWhq+MkENv5PdA2qhGGZx8u6UVziiYk1P
7DH31Jg8a86FeKDm6GkK8vNK2vJ5rl65gTkLWd91HFwEbB3QterMv5bZI0nU7ZmbfzfImdoGW0LA
KXIKGPGmK6Q2+XyfjkIyXvyZmynAhuFYMmKCbbrswb4kt/sTzR5LC/W7rVyi5SF3wsriA885Qo07
TtokXUD2zebLOIUJ9LoQ4spxzIkT0tLh1oefaIidhEfvRjosW6zikLWcb8jUh8z0CQBcZmgHmCG6
vFgqpem6DRZm5KoyoiEU/TfM2o/Bpe2aqH3Iw8uPte6hcKSSpR5Fzq4jwz+XhrtsQ0LR9xhVZs/x
jNs0XXxBj/oZI5fzr0nvCfH1hjgby3xU3GZUdMxu92ylaJZJooiPv3T7Q0wJ4F2Zpvx5Ju/Nh0aK
de8OQLPCziVRsUG0DeMFle3cfppk8vitp13i+p0E5vD2NNQLrenNB7CWbRhhUXJcUpAn5br9oeX4
oQ1mFx20wGBlpamW4ss89lLqJ/f/nkkqpDlffvT4S9+0bJjzRh6i1DQXieZ7DU7A2eOPGjEDZkXu
Q1ptSisP7Nbhb8r3tOkeaHiW7WjDuQk9LOws9KrI4dVhWWI4YXXStrcUeTceTp+2R4xClYC+Vb3c
39e5Eko9dhq3aNPp7AJZRYwlXsBfmH91ziwcwGAlYGAlMeyAZbdoxDsvWeJNZBqE2ASEjMeXbMev
0hYTJ8o42hShp8nCSUBoK9vuuzhCucvkaKoaWyoUolbzLsHj6XYkoQDvXGiyW5th8u3RVe1Yu8q4
YxoPHrGyM4qo0hRVL/NjEl8b6mpU66vJhmOTrhDLOOUXtAGcO5VrkZwMEeed7hBxO3/kE6gMu679
JutFBuOSe/+/55HdM/1cGh8PDIWp26U+z+nusWOP79tsqWiJK43s0FzyFsUhb/SmlevcTb6Noosh
oHCS6E01zlmkXQag8nvdQXZhp8a0VMlF2ZUyUL53iibtAL4pZ95qeg8tEEv2oyQpH9B5Z673Vs2i
d+vMy/VGFzbM4ZKFjuItd3HcxymybalfaKOCQRr1O7hr5tGOOllZzLe4AhYoIQaBBS49Rn1UUp4k
PsFc/g/6S7Fal+Y4AaUaoDheRcfftJHFzs0stJcun8D96MjWgAyNrk66PD5F5E265Ngt+LTTdMKb
/8orIAw6mB01BKRPezhreur+sJNFoRv0sPpgzxt9/gZ/akghdLooziHyVb9lDJJusYKYMTVZLhDJ
Tas16l5YmK0DfkylPf4yEf3yYpwKl3OFQ36YlhiTFltf99e6PfqyGghD6sDgpYr9qo8jkuLjI0s8
n75PK72K6rOy0gqYA3My4B1lUSAIRnkReFOn452T5Tuj1btPiBYA09bcDMsvYOFQHKxVZheSll9z
Es9u80wka6KRkBIMesW0fCo3mM82PneS4D1Mi1P5HMfY6gd0b+xrrPoRbUYiWojzeKs3wACZXmZm
WAsjqZ0vPZXyYDV9SrEu9XtNZiDe+JIDx7zKN6d0OOcpJRKPRsNGJWP0UnUTPj3RtIQNLulF1Qnc
Ld/0hVY9MQERXP6ePnfixDaigxyPx/I0Ime/EYjFIhnaR+zeiHtonk0TO7Ol7bUaJwtKTSSVa/Jr
klysBsvm5UVI771izkEm0526ZDIyrsTGaF5baD+g1kC+sD6mRQbpk+7sTjM/ISIfn+zKHxy7tmLy
EWtr4S8e7CJjX56f/H40fRlANzdeYicc3DljHq/mOGLvQ39LoqwK9vVjniGFihRQA1KUPMpkXBKt
KHGstbPetFO5Q1MWDQtV1FGyeAFumRHzM8jvPPBiYMP4cswvpGPy4Sz1vklTfOxwKW9o1itMw0Pp
GlP0OsL/r3Kyg/zCYsgnZhdUaWjF4r7eeL+vUaNefNiSDCth5sMJQIL8s95puarDGK5hO8Lh1uxE
RQJN0NXyDv7mKHxVplj8785ia57AyErh4+dpPK7Ukk7lQOKibr5U3jw9JPkiVJYWU29ok/hv7bvN
baWPR6LRHAn48VlJ4h/ZhhoN+LcPqYhCUS8wo/4CuHDqgOyptGOV8/yu+czau7hl83QXpNmeUlCH
tw1tlV6jNR0QUNNqZ/MBHxVvOfkneeAMgqrAC3MMTh1NREw4x/+MRP8f2OEMflHr4fYy4t4rHlHv
fNtvpNOWR2K4RHRkvlUQrEpObxQOlO39CLoOTsy+Py0RRvSkirOxyU8Jq/V08WMmnryXY5WfrQpB
KTSd3ZdZ3zR9Te56CXbuA9D7Y1hRgLMwsWQFgx42hB3X41qpCidmuq/TuOy6QfUIxR9qKkamT8Mz
hI3d6C1vvMED4EVpim+CjRxZ2/0OotY+CAWWpppbvfimgSHsFT1P+FD+QZib16YakmsPSw4OyFmM
O6r3z3yc38Ad04uzqnT1TE7s26Z3JkZFnqmB9Bz+MVeiRkZKMcYtnOH0x66cS9xiFKQAzANZeTOb
IBtTiou7RqQXJMimKPbYGhx3GS+GCIFOQ/CvJlBjbHVXWXEsosNlVsYpRaKy/VplGvysO7FJ0fq4
aR49V26rUu/D8qOOtN1gNjFOhTkGyK7k4HUH0zsGD05WxGC/I7l23BnW5usHrmAtQFVb7rOMEMGg
C55KP+JzKAYu4rthtb5WfxQyZ9mfmnacd1zCmBWCvF57lFCKsVJOA+BTYihMLYMqLjoEOJwHnTgd
1d/MLhWpvRdY1g5zoU4JMklhX1+bRiyGe8CKA/Q/2tXtdn0W/aIfAknqO0eZJWAO2+hUTF9/av02
sTWtTY2swHP8hc+m88LwTqgkpaGNdBRBRbYlIGm58KxOVVD4MIOIaXXzPfd0f3lV0b+M4dS6FsCT
pN/GTWeabgduvYbBdnbkaSASlbJ9zWAZiyPY/BxycqFdwBHKVTR5NsllPynWmK5MyZCV+rRO5CJk
yDxN+g6UaLw6KKfC2YKa/VJi+L6YfCc4/os+pA9jGCVSa9F/fggmcGClW+rmF34hELvQH7kabxm5
0rTxFFMDcy0DASrdzALzxudUKdXsx9jQK7G6VIA/21PuC44Dp3iCDBmNwHofOWsm5M13sHGESVZA
QVs5Pz+hoktp2q6vA1KjS2AhKqC+i8N6MWi4FhB6hvuRyr2NO6U9nu/pk2H4t/U5aL8F/iAkcX4h
vQpzwsUw3TgpwIfyq/J8oLVS+OhHznkVAJD9hmRwIJ2eKXXf0pEcpMVY3Y8p29Ly3x9UIAyep2X8
u7UvHBlBFthTCzvQI1QZRIf5CkY0Lva+GYKSqkeE2hvWXxcY0A+IlO0RDtV8L6mqYv8aYWxfgcMN
Lxp1wXbla2XT2JdyDjgEyIJeFBPHkwKE+NLKEg/ifaGLEUW0JM/8fgNRX1F+a3juYW6T8ex6hYc0
HiA66EB1kn0c1dTm0Jmpx2P6Zz6O3V1jnIgHVWVlvWSSI0jvMtD7+flhGGABOFlIiZ2nEwycyBnh
c0LUL0eDlwX/X/vBFdVXP/htZHwObGPNhSTlf0JV0n/yr9iv+5N4KfmADvskGLkceBEbB7M1umkQ
NhdSntbRBLIMBZdmAU8FHTAxkvkUvEsnClJwMsJkBNjfAAkOywriGkTofGAv5LvueamoyceBeZ11
XQ67JLRNyZQNASWeLYKkvr6AdxaILyle5ewmFCUTdjLmf3R2BC8rNchq/6q1FI79h2r+VGAVF6YI
GHZOB3+FrzfoLR+oPdN6F5ojv8C1fTFrJYvquOexBFrGftnFBCR/0V43l7kGr6d2SBxKhIrXq+ky
Eyuy9mEXY5iLUC3TUOIJ+WX91KON2/dUuLLFqffbwoqAPI2d/1Gc0rZnC9xe162fy0zFMmYjQV3t
mzQTV5soEDjM4UIpaHtjcCKrfXKZrk7jA4w8BGkyqh8dac9MIOstwM++8T87uaIgq7kEZjCDkUJg
SWfqadgdLOztaHxyOunO7OQ/QNtCaI5MaVF205iXRckxa/vX/st43qeeXG5EssBrdJ7Fg6sFwmNm
wTVrxJ/58+Ko1bcmuZRcVnmXVdwZDSRDcwa78H5V9m2toMBYMrJqQGDoZ1joTgWbVpdihx1yZgBw
QzJ+aEySyBzJf54QZCf4fmUqEShXoyB+orR9+YYm/2OUKRSKpbdEqHmSUuvbEK82qpgkqRkk4TOG
+3WkJF3+PlHMBGdUPNGCl1tYICHbgmpVY58Py/wo4bSgEFr9hljuiKMboMofh9XWgD7CqWF7x1Bo
twuXOLudHLX1HuBhuzpx/9qW+Tsxp1WtWbRAKrXjGXFaqGyxHpzd4T+loxg2CGH7NQMLG2Zo5aPb
zbFIH5msOcei5ZMQZdvvJU6Kb3MkwSWHYYeRyj/fhdzU2p9jGjhYC9g4i/VdFSYxDkKhzkalDNlD
UrYowQt/ifJexQ5hNzDfiwPbLq91IGRZUH5Kq5AkSG9fbXTrGSTuaCz/s2V86rRbP5vkC75vNRp3
AvgIwN0ONVukTbjwllROeyN/I4PTsZfaORe+Jc91U5O5Df7zbJrkfdda0KSlQW3L0eG0UY9LUytM
KI9v3ChlImWaSeaNADA9hqkZSD66YHLmp+ZJaoDM9YQz++4E6hYm60FFlHY/dDebvZ5ER8bcblCY
EhYJhgOqD9Th4JIZwtYcqE/ym+FcgbL5ESoWwqa0xfe7bjCB4ZqPN3gGOH0b5pTWwsglDVCaEqIy
lfNOtUKz72sWGJN457D2Q0sRteropGLb+bLjy1aA5PHc8LsxoR/BJVE5ej7VWjpRxHxH37div3N2
yOutdzNhFFznVYqNVmQpWTepzW39wdKTKNU/bPKK7jAjfLe7oj8k8EiYpF84wVXicK28Ujz7QV5a
41jIpR5cWckVl4rLrgZxzYeFDbeLkA30CeGI0OCviR2RiwQtj6Z13SUG7ttr/tM1Reg+Wk+jdT7B
R4v6zLQreRyY+t9PMOIk11J2JxAD8fN3QabQEC6fIh+tRPrkZC60YwN7/QIrBoC5hBduMB2ukIZj
7LalmsN5+Ho83ozFocQPXU+DdJy2LW2tVRXjcDpC/8r2wD/UZ/PqQATkxqOLvuFZjvC8iLUJEGKe
J8kbIVLu65t89VKNYeFCiN6bNnn6Qfjgnm5Zi1zVfYTteCEEvEUibil1KV9IPHFXGAlbU8bsdkqU
+YRk2mMLKALIVP03qwxLJVljOfRSfOYLtd11BmxcWO2SYL3fhiTcK/ntke0CWP1SELS2XVDu4uRz
OoRqAft70QXEUDTmNIeY/coEKL+YFGbD/Z63arZi4WkA10WfCp46OoOPsnJe+u53aps613YMC0oA
ZD5i7wGn5DYIfEp2d6qnno3+IhUgDxmX6FVGuuNZvVq4bNDaCVXEYKzgMV9QaY+CFM+JjAuITqWm
NGgnY88mmjByWIIWupj1piPv0poweulc/oqP1rRHsoGm223YGftsowc7XXh32kvNXR+ILUF0mDdM
PkctzRvc1dsgSS18BNEyQmnocDUcB2dLPCABtcNAO20MFBPQ0mmdnazuOMg4Q/C3ghAWJg8wCJm9
BD8XamR554UfDxygLyuSPOWhVgq6ztURYXcgUf2bqKPYCnm03wU3Qof8cyfXULZHH3NITwmf23dJ
dfuT/9tn+pV6mhp1j0N5a0/cpdcadj3FG+AW2E+qwB/GbSauvJC04GobnrLgM2BvvG0aEoJzJBdB
zuNvTHZuWjjJsyLNl6vG5JqehjwUUhVBGKthNgS3t0NDI8G/gY2kbRgmGBFxwtPfkyKeZngZ+QZq
i1K67cIdenTEHcs/zegHz2QkBsdIN9uAZh7fDM0yoi79tS2ZaRGEGMiLDPyItMEcAbuM9Mb51+k7
7dayAu8bnNcji9tBCQe+Hqvj24tg+ZGlnIgqXV2VxaC3o0ro9tEelTZV6RMLen9865tAnWh8XNCS
sewMN+6eQAOEfCauKlVy5WsXg5ZDy1MNpeA38XSq5gMISgiIcf8jv1AckwsAhu5Km/rVmqi1noIq
N2ARv2ppXHNpTRJUMVvGiMXXsRy8X6hBFFyK4znOy2zVXfQRRvX3Tq3dgdl+LshVjQB9Y2nhOFmG
KK4cUrqj/HWqeREV+x60yvGUvZ7NGQgDa3zPZYH7sb6bLMd4f8N23qlnpVqS6Eb1QclmL+Agk+nK
zvrmhuPGKbz8qt9Rpx0dJbGihurFT7uBtm6za9WBK73ov7fuSui64I+NdnBKz74iByrAY62jQF0U
cCraihyQgjgmYsYESSCdNuGaPIbVApjSMzuqwtcaG5ZmbsBaA76W1UHJqJfWjW+2g3dG6qGkQ286
11SryuBRzPplb8w/rDOeGHnUPirFJAW7KVyvpVL3afOIsSTUvfpzXkUQxJPZ2YlxwV99dztjO2pr
3/lVLSYUGuGlaYDGRtsyHM068SmwzI+nmkmbj/WwjY4YYR0gxZYr46trenW5mwrZBYCXAGQPDN6f
BXh4CFrLeczF8C0JhWU/JZxGwgRZ6bcLPsq8L7T/01n63n24BD4bJDYmyP2cIJSl1Pr3smnfuC4w
QvC5bNjzLolFans8K6IOW92jeYYE0ooYLsS0936npEMaX9Hz4lrckAdQMbQn/C9I1sqzjracAsvy
neRIuFyYhQUKCBWTqzguJ6O1mQHYlfz3SixO9rx0RTfLC5ZymMNUEtor+2jPxmEr8CklkatvLAqA
ePH03J65MxjgeN7osHGnwL+Xrz7+EKg0q91xw3OlwFxD41SC+CL6og6ow44a33TQg9Kk3IJ+S602
BgBZebLI5InenvSzn+Qq+ZtBI9EZ7+53sFvNG7DiBXnRnx2mwfhK4pZsiHNwLVI5YR+sIwQwGpum
C0miu5+jsOqvj1NkeCjxzt2m6gj5ZI11nsjMRWL9xvH4d5iOdpSygioiXBpbQgwJCEcnEO3B545o
2mSDhdhluyzfMdwO4lD94E4lOoTnOeQQ0BpAg3utqcwFSc6vDsckChScmd38uR/X31D7UbOtxRqD
nACNcr4KDWlSBZdwGiDvriUd1xGK8b4a0IgEe45CQrHab+TEzthWJTBP6casDCxZeycz5HirS+81
mz+iJmoCWYGAvm7WdKekZO4gRjo5FiQneFKvL4hSN81ZatmtOLTAkHTFPiBKhJ+TzCbfbkX0kK/0
XUTPYKUeRHb/wkxru+shjyI3gX4+K7wZEgvMvjyuj1z9YWTzD3IaqoDt4Wnu1T6aGGNSKnOZJs5G
8haW0Fzywt7gRopmBNEhBGCm69X3RNNPyTEy6oLKnmwffFHEI4BW/4m6tuCRFGZX0Dz9v3N4VnjF
Nj2eHHAPZEN7fjobPItgyodlKzoQTSW3ITfT9REvbIBghwMV2bpoAxo60R/gDAY+095Qmm9oEFlS
uluexPMxJd+dl0m4+GeRDGpwu9dm2WxgEVZ/ddQJAJlfeHRtMb6yj5qOzdASI5gbt2oEsRmVLOFR
K3oxDAAik0A9f9CRguwdnEOtfPcPFVxC5RfTY/V0T2zGGf5PLDXnc4VkX7m+JMsIPitzdHN+AjED
Y3SWOgBo9VO+wcIJg5XcD3Fvh3BrGhdTf8F4ReVlq639KbmRwq932FdYjBwjoVeV6UOVG0PgOLYZ
9V755fSN0w53d4k7a9PBCAxXln/ztC/yR5urcGb0bItV0GqqtmanydC+YMS4pH9P+vhddwbxVEWE
GYJaVZ/GtqcBWjmYJLSuKuvet7soNpz9dAz8DcX/JlNa32wI9H3PQqJ0caQeM6U6hBk1/czuFnfX
QBBcFwTwCq5uh2HQsgML0z4Yn3u+HPjIu3ywN/+U0zI7s9zaTKwmgF3/3cr/3gi02AYewx/iTrEp
r0B/EsNh5vDIfemWT0RVghs5RHjvxEUHcTgfSMJxl7OvpcSZNSH7q9kqbzyIZmTjHwFaJeArfH2g
xZQtxT3eawPsUbq8JpHDdb06h0t8Rt8VLODLGSXWEyLa94BTC2MPDQD8s5PzjmjsQcJzI27d6hMO
9L3L7vxuca7Ays9z2vOpiTEng2GwpHlW7V611mAhlUi1YHL59sWNdzkFLkaAc2eD5CE3BwergZJe
9tPw1Bfd4f+5ZVK8iWu+r6qCcd0PmXVlrdO61/GHeu1U+pg+no76ijpS3VwzfX5OR08WCHPPR7sn
FcnSBAfUFraKFTtCzDCuBtHnBQtFd9XVWbgIArfrF8UtCyOeyzWr5+ksnvAYNnvj47icvwQ0QahV
WCYpnjzWMwPXNHxIfEQYjlRNpYlxACThiDDFS20K473f8WNN6mkviMiqDi0yTReURfsDfVilSY2p
A66+t/o+o1Bw79AtLCl0o8qRO8crEPCyEUSubZjjMXm0p0EWCGENXUYGzydYzuZbnMapNy4en3yF
Ve98gHUnvv/UkCOF64unh4GRFDs5Ak2+f8h7M6EicWU84hCeFGuKma42MQFq4cOWMIm5cW1oMaNS
5zR9xBWZx8iC+FYzuBR3Tbwe/vwuCK28tK2AuCzZ+J5VdTbrzLnLh4WgPJBwqmNHjj6Pt5ChPMCs
qhekQOCgHKl5F0vfMqIIccHyBOQXC6CDh9NededJW1BcSKWCeg5HPUC8s3RiVvpdKe+Rn2CqZ8sA
el8i+v3RSx91Cog6mEvdEjrQXKlgk0zZQ+yjbZMHnD457OiXME9qo/QleaLhKuKdWGkJTJA1NP54
sdPnxnxQEgMkFR0tfDHQrnRcYXYuC9sPFR9e17+T2IF4+JH5jYF5DYEULXl1v9QKHx5rQ+wd0aNe
SJ0LuAGug2kLBrZgzionScJTvL9n7Y22c7jHgS79UJkS+yHi9WieHUmCEufD3FfCZOedm4+tOdR4
THJ/gCtb5gh/nWvJzpgZmOh0mKvrZDsmxYlIE2Qu15YWyQWvp3ND9LFXGV/xApOBxRrBUG07C/dS
bSFYh0/2jbopNuFQTdNhNk8jvvz6r+pkX38wuT2tzBaMZmWt40QKmaL3iZeggVwxkevq/QXaIija
viJbLXQl1glJS/hBHJSQtpBVRWiI7zRVoYb+quAPhU9G0Svl1vtpvETkKRnrj9uX6ZCaxo1C22qg
zoBjLBlhobzBE1AfHn9p7p2XxGqVatZFCj+ksKBTEirdg/go8gCDrukolfDUHBUsAPh21ciMv43Q
hQv6y8sYwl5e9+YaJSFKQRGQywB0WAcVv9ED8VNp0Do3C/f6wNqZcgTH7DbxGnegYnY27xQdTlMy
864tvPpDx+RSHQ8B12fWysv5ZdfN4YnBDQ30cYuyAz1rJvzddAlMEe8FdP70qkSvk3+j+MqD3orL
ImMP638CZveo/eYgYV8m4t//qS6qWZ8+Cduyb1bcjqgQdGjnJjyoiMBemTNaMPn3NRswVvT30SOZ
pBYadjqPLA/U+A2Bzt90KH1t35zwWB8a//TuyMa6MJ4c/uuORuYClsnGkoEytM9PmDMbumEB0YV6
r5TYwsVcPHwrN/s8LH2paptkxlOUxjTa+H8XtA7TIXPAbESwISqvZuXAexA0V+9eoU8M9C6+KaPD
AVZjdouUQxZKYor6StfcFsc+E1hAe4HEF4r8lhJouTH7WUnmTcOXxhNZy1qXP5mDLwEMZlSP9Gc2
g/hdVLvYoji2U5SmDSOn3qk1Rb6qoL2UWjR1zORlrDI1wxzptgar8xxNFW662JAhfj6aaZ3EaB1D
erIl2nZkDQjgkqw8N7utoyfgdCSXxU3lNe83nc5Gnb+y38VYu1WhEP03ZnrqQDs566bDGaMWdNEI
0J+05j1Psj1GF213Gw0QUm/1Pxrsb82xcStFjOQheMBx9AvegeArkZurydjlTFSFfzsHQQsyKfXU
Xgt4OnafCbAK/XqiJmPQ7E83KG5rBbvtMtHfqf85aUME7jgHOYDf9UL8p3V2EUypic30ic0wEI9U
QjE0FgsGT6MwXsLmX4pOD1Tkk+1sGw6ARgCl4PeoWa4+3I5I+oQn+PhnGIh5qXiWieNvroyFwEjR
1sYrezisw+2QzNX9ng+nyHbZVGSyoUg7cfYOPj6E/+E0PKRjzAJM5/TWuD/EnGCoKsHsLZe/Vpn1
OwCrlzO621L4Ye3Y0gLzNxcw9Om4DxFx3kFwLOyEitBHVXiw3i2Dn12lCel2Ve8e6gsaBLR1tvmh
KWPdySDYOtSdn95jWO7mp398HUXwKvznD9CopzX8CicsHycAxcfEN3abHbq0mhGspo6ZL3AtBz00
SSduZ7dj1RMkS+FqPtNFbxyZR6LglIeHu5SUC8s5VmqlKh49pKWeeqkDQshG3cjI4OxJxL8NJx/D
NSvRbO6zXu2tp4BHSvSPaBbet0nxxyITeFsWKgHFhv8nk5UwCOQcXKD9NZhNUd8MqUIsvhq7DFtr
UpnLrIEyPbBq/iSCBvTS78tsHkP0k9ycXQdZUePxUtvdx73cpGpBMczFFozN/dvhrOs6FQ8PJ32w
Z3qrnsT85XoU8iz7GdW2p6eXECLtUac2rpYDjztetFK/OJ22ayeHavH6eY3SlBeq2QaL8D3CCIJ7
qmC6htR3xRMLK1XdCPcA3KAsYT57b4FR4Dz3fweb5lTjHFkNk2B+eh1r3mWbfKuNTHLbIJ2FqigF
3oTclUzBh48wLWhEdrqsCCZsL7z1ZgU5AHrVDbt7BVbNTsOCkL/OcQr+MCHdIaKmNQSFwPPkUGlH
q3B9wqc2qlAddDILdSCYaFTsIaazEgRw8sJAel2j3gcLGeXpYzVIBK3chxY2cRtlr1AdFCxpAlRB
Y8I+mr8tzlnZStunQJolwxUfjJXW8ngGnP55a0x+ihV/KoFnrNq5UwfRns12G0tsWx6S5FuaYXit
P/6tTpLpLh0lifOEQD+sTYATI09YphB/s0+aOOpTaEctZC99n6KyhphsJNUwi5gu6kI8tj8NzIjk
Vp941PXBf6RwOrrhHexB4sCSTrXYp8QgUSMZDkpPU+rXl9Q0e7Dy642pLq/FYG0u33h9nAvAReil
RbljaNXXSQV5lJkDPl/dp4UWdK59RW9iAUIEr3wYw+9zmEDeOqAwvs28SKEKK/2IxbcpAviMFELK
XruG91zRC/6SoLDy5VSwfl/Fpoze8VKs/I2g/XOtyz4S1mYOJjQoTqkWqvo1oEWOsyrtNEZ8TevB
tlUTkWtJ+suniiYvsl3jwU5D7topDonYElrvKq0dlTBXpP635otzRFxf0RBp9zH+oB6c4kAoezWd
FPwh0mr3/uyxA4GKdMsxLzoFCodEVeg1zI3bvSIQAc58dkFeRMsK8SAM0kKTVESkeKtEhgnvq/9k
EbfE3YqUmjvpIH99dwIzgqGe2Cvx44+UVnBiB8MnuzKPNLtyYTqwTbs0pYywm6IKHEnBkvrs9qGn
2yG8DvKT01ieTjMk9zb7WpqNOHmRQPox7/GCgtZD3fgPsVEFK2drAPvYOeNv2qo70zj6j0B21UaP
/MFxYU5LjyOAA88WNaaSprNTC53xvwm9IhUVnXM8Hfsg9N9R3xQ2mGP5XC6JQuiOfX+Q2SZmMMua
3p1A7vBQbxq+7Um4M0rFzTz7A8xarXR0EL5hNeWI0aO+JoQHWd9RQIqjC81OKeCula9MYmemoWgR
1GiVRuD6fyfhkR5omCHA5bqrQN4D7XV2JBdsVgkuCvI7dm2OteQZsS18fEV/mjucL5pO/tOPzSCY
4fYfOtJN8X2qtFhgExCBW2atv9ZuszEyGDEAPs9C2akQ+K9oPydGIP0AGHjhTV++xUrYjIlFkNnu
+YV8/fUgHvyDZze57y6gMT+omXBKGTyMP37/ME57ZYdNTSme4KI+Pxl9pmXlAVKBkvg4QrW8pv1X
UGgH7Hl4cjvkQBPLsqQlc2IE0joRvEH245owOcgPrS+ZjkJDGKaoyvCKuR0Wv5RzXL4iMZzhOwfw
T4jhM6wjvdfWUOEqv6TZAW4ownKoZvAQHDD6rHbPU9gzn5166qHmH7H760H8FYUvZNa+b5rd/dc2
62SUD+q9qK7wAKuWzdO4bjQlkRNDJIbq4KSMd14ZmyIhaXNHbTvfk6ROcaMMIUn3+JP1xDr2eIye
RonzVbORru24c9pJuoeOSyiW6e1cF2haDwePNHMMdSRKwEbwuY8zpymxLPkcbvfP1JpN6X4ruCuj
pOL1BW+yGDle19Km6lg1dV8z+pNrlhCz8DBNovrPXZ2/cs6IkmLR6eIIRULtFZSfeQjIq6x8808B
R+7hQY3KXdXQ61PEPCXQ0O+UIMGTiZnDxU0UAPSdDu9lfc9oHIwkXMRnxp84ICHdGENOnl07VaKp
p9TOzNzTxgdTnE3n3mxYu+00hSaWdp7hhG6CGGzLC/3p7o/TeDitjfdZVXqiKe/p78aLryk4CbJ6
zTiXGiA3DHsgwYBapV5umk5Jw1+/rCIk8WiX7f8Rt17dh0Q4Ea1I732r1Trahyj+9v6JhN0T1y0X
NpYlOTou7vpR0nW7o5fe33GrWvk0FUhnz0BJiVX+kexe/qznD8OsCRsoeh6GSXW+LCIQCuV+rBrn
O2+EShaEwW/VanYkUoLPwdrvtIfBtWSWfEsUJTj3h41IA8e3hIJHkiYEp5ew3KflETBt3xMJeaXa
uwONZnlTt3gVO9mENHuznI0qFcsxvWs4xZSiZ9B56QhYx0DGp4JYWS8BoxvfEJHVL4+yZHvDlSaU
29WX9F7FTXxhZe6pI7GTNlxkZXnXFBte06RJRa6oqmdxqRdL/ZcDNr0TP5U+gpkRasYrjHTCqALA
w7nRuuTNsAXdPnesI2CC4pEcBDVHng99bKiHWMGq/GOCshHBKzSVrNZBI6hOA3VNd5vFanqH8hTV
SMZzKWFU/rKjQI4HrSd7Q4fqNOBP+h0TqeAUrCMs0DKwctw++j4shSgBKvJWnzz9Tjg2cKtAVMTj
MJz2FvcyVULxSR2VxrnltBEjJuA2uWYwcRdwixRU6hBbg5FteMlQyfthNO/dxGAPKns0s14EFrdS
P3lAokzxQC+0lQFmpGc4s//hI10TlBAtcaSTK3PP4nCrob0IR3aCFwgNhb2Bcs7aX37CwIuIVggs
+F4o35V12fq2CwExoHr3TcnansItJ+3GtHCsv0oMqoANAQVk78d994UQI5jKGmf4uLfDLYsVdkP/
hy09fWbE5sgi1iDmaooKIb3cF7e5F5gXXMh2URZGRLzTu+dq5nSpPPxH/w98Fk97HDqJAtiKTiU1
IVrDWBtMIqfZ1jpTC5dGdqqZeorrL5A9xn8x4saTqiwv4CtD8IDzccs26FUeo7sdRP9FivgNHltN
enpCdkEzUIumbPTPowTQqQRqsN6N6IaJhw33F8La7HF+q0owrUb0DinaKyl1HNzmPDWMwFX1qtMv
e0p6dZCx0k0ae1kksHNLjxvKkaYUqpOnTAAjP8kyZ8WQazavLqAR0fR5Jsvsc6Eb3y6fGZaIiLgp
hlCM4vUoq1aKoGzzvcZYtTIfTpY5BiAdkv12qfg0ux8No4+mXaIAhq3nVZRkRVAcLT7cVigwf0ZQ
FN7ETrI5QaGYu1S7VSjfp8RkUcPB4jFkffPhLm96+KeIc5fXuYZsGbyEK1t9o5oJPB/HPdAgxZId
b38BOuNoxVkRjPOPmIkwS/90qlHSpXSQNDMYo+Ab3Hm+Pe77UfXMYT+FAA7MrDn1iUMixxXoUs8Q
sUIWkN+wmh38o+g068T173gIWjK0/U2nujw8qfK8T4jPlWpsWV1TXTo3RyRDuf5v1rwCSYCW3/nz
ydo84OCXBSkO56+93A9dTdZJPI14iRkRSrumvEb1Ld+9napgyiQudS7RfKsR6lyTrNWGjHXamrXC
4kRKa2RpeqHv7IPRdKmJtKfAVWAWJrqdLuTa39fMM3UHOjkg0D7dVMFK+WLX1Qa7dWVCkaf5JOGl
WXgyuEKNoh3Ovdgzg2bQeghbzCsag1EC2bqbjBI/XzWXiluZ+ERFBfCk0d9hwhn2I7DbITlKxpnH
CpSpDVdDQ+1e7dIy+el6dDaPfB+6ypZXwlFwzlsDBRsdWwWgJuIsg7ob7yezZ/3YhdPRVAmXnmzQ
g2Zcaqtg2q9UfDoNKd/JOcxehFIHwXupt1OP8d8m0lOimykNTozPhBKAa20JmFd/+V3ug3KW1jfA
tpdCfo3ydgFw/Rjf5xnbbT3G1/25N14wJhMl/dk+P8CbF9mDvdNMpflGxbPJRtU4uAW6YZSRAhmM
EQmRvUI5uuCZ++m2kwdKXPMtYus9BiH6+JGq1Kn+vZMocZT2pvF6Lj28WEmQqcruIh8fuOsqvlR6
fopzodBPDdZ7AMjCY813dgBH0mVGII3rIJi3V2gXTViHfptJpQyrCaRw5mguxPGvXDBQ+JlYAO3q
URxnEC0QWwvkAya0Iy62GIxs/fCaFg9JmfGakzYIhhLwkhHYNykSN8ZYpH+W1cnzrCGIx0GQ7wtN
PQVIQtX7Y3zAr6v/oTRL9m/tfV4qII9bW+AbiKgMJOi1xIQXly2QpsMtNX4ewM+vdjCxGng3+813
ranDZKCaPsDsF1AJc9u7XF1OnsfPdICjiok4NgoF25yDbxz1kVtaTlhDGf0+3G2AqmytexRICWcy
8Z5QyaDZlJsMi6obAjPLLOhxe85VUsLsk25GFvXixXxZ8Rqh/aXhKoxDXPsjVJ7QeTIMr3/LJ82z
JmHs6qdeuUGQD4W6rX5w6rQ25+6Hd39GNOXJtNZ+j/cxiBmi25AuPy0T4KhdV+iiMuuBdPeDPrd8
eq0ft6cCLyJq50TcDBG0JFuoySYewExudxiA3xZ3XpAKSncggRRcK89r0mmIx4WwuguMIBeIKX5C
tAHX9E+8KEyVZmFBoll9a5gPr+0HMm6/eV0AsxSFAuEsHSLYZTCjprtP7wEBH/H90TP7X0iJ4zh9
mWU0bunWtAkB72SQDx9b7Ainbcyul3C0Eg9Sz4lXQPjfCtnlkTSf90hEs8JsVBxl5k5L27h4jr2K
LYvBXU+EaRmrQqtv/bmt7dXshhT3G/+ZVFiIo4V7d5XTCejWzU8GukiSDQKUNzAhCiXWe7vt9++v
segVnr2QYQChAtZsVEkFTL7a+SZsmNzUBh9TExn/+iidlA3wNkGsN7lgddaF4iAAdWwfD7ng25tb
Gycod/cV8eiLViDfgyYX0HFvrdY58vJ/bsEHjvOsjj+9OM+ainZ8864OuPP0OJDRNmeekGj1fm0p
sdOtDpewaMhky+x9o2B7gOMAJJZ2MSEEgA1k296HZ4PWPp3DITptk6yGXddE/yq9j5ew6UJvkmop
QHDHFB6ir08LxVC0JycP6uYoUatHluIq2K28R+WiQSBpzH+7FopdodgUJy5pvQCQ/5ORI6xxCaE8
+99gvN7Xh1IAvXOxcVV44zl3aRbZESGq2iyD3qZvs2M9mr1r/Gb8uT9oaFDuSG/AY1U8K9dyQne4
p4t5pIXc5Pws8rjcJNASZfw3ESPn2n3vwe2JaiFhIP3dUa/gEX6A1qTP79hCaXa9Kzqc/yiF7tp6
oKvBeYK82+legzjju+I6LX1NIjPPQKMLv37bij7IgfQhHuJCxII+ePCb4Vp0huMGrcBZV4dC0vu9
aFSvayB02u8r4MzD132YyBDWR0IN+n+xBKEfCNU7Q7onelQR5BVRfRS9nbASCM1oyRmM5ALk1B8E
FJsn9fqozwMhOApvGwe3rEUDC67kucc3MAGtLzpl6J3hBA6zPCL8iNU836F1rpVEJXJFsWhIHSVq
v21ckYJcvWxbovtFSlO8l0bu/ldSykSJ+WKkoQ8h336g+V8DOhaliGSYlm+5gfXJ72pnCkeApo8C
zD3s7i4oRUzMjp8HWG056S/v9UihzytGrhnoGKsiCl5U+ijm4mrX2jY5mzCa+tJU/RuOTP/49WUS
cqPQACy4ZqfhMHE8MvulrB93V5dKHNoD1OlEulr3Nfv+ePGg2PZ21OgEGc/hoCaEW3s0/NQHABto
DIio+g6MNuyC5VJ6WnT2KuwvAhlRFdmab4PZGIacGT4A/xyohNchO3d4HADPekhMdzEsVx/yhSXz
DfuscovkaGkwWZ5/1rGyuRurNiB2aEPQndfJSnO2je7ZJceYn3l+Is/mND3CP6OuzZZrASm4V9uT
HdXtdW97h+OnRxJO6ioH9Aprn7f0tHVYZSqHQvGlJGY8+XoKTzvTKi3vEZA/LwzH4xnDwEY4b2XF
bhJOUF45ssON3tdcuAyyTKtT0V15GMg9B3xc5kJxOh3BasN6dJXp65aC9bLCKzIEvmWlIyFymdOA
bWfdJUNqVsoypswQH8nNZ6faYtaoAiwJoWqVNuSy+DNQi2zGAFxrao1AM7paAZ4m+7W/oGaDhBGV
W3uojQrI/4V2x2YIv9cKZkqL9jgdI9mFA4ScJCgX2EJesh+RrM/c8YcFdtLFK/lIMA7T9NuDWX+U
z70zaXfXjO4VvtlwdeojX3DIi2VkAccu9Mlr3n8YZYYk0Ec3hzlkSGA+JtWITx3LydAwu/z7YAFx
mos3pDbvxVxm+CqdXVbYKEY5iBbnLvkuv4x6Kt64hS3VgoW8AgcrVw6FnRU7xXnoddNOAiCDqJyN
BZ+1JJ3Gc6gbV9oqzVdEKp03wWghG80aWoB4hIbU27aO5ER7VpJNsgYTCfQZUXtmd50QjtEZaeXQ
n9YuEVtfBbN2CA+14Lqq4+X5hX9y3whkDD2w6moDjUsn7zn13/otoyXv2GmmjtBLom1Uqg/5WAb8
Ou/ZWO6T1PJ+O92JW6zeiEJsIpGNjijqEpTmxY/9V6f1yBnDYCEFluOg2pTwFyeehlI9VO7VnBSY
jOnvWhlktimSzgliH5Sft06npSURARH06Cko7Z65s2x2d+c2xOsMOG5HuSMt6IAV3muBu2kdsIMj
Y5v/Cm9JPYlSKHiQJk1dwPRmRfzkhm62+NCrYmSDeOM4bZ3CivyDI9uORcaF3dCBdmgSkUeIepcB
X7TCn5blWZoGhNDXR7X9tsHsTAyvqMhrA7g8Ttwelyz8G5xDc2DxmZ0+9nV5Qe/fg6nJhVI54HrF
5Cbebv5kis275XFogwfBjISpuYMFMhk0nx4qwbqNU78tmg/RAii7B9UZkdO1abO3xWl+FUzJ+1r5
q8CcnwTCDs2PcUQcLBwhH9/u6dvm1pMg0zNfKzPXkS2H9twA0cNpREeTpp1PG4XboAF1s/kQFdTJ
21EgP85RhnmtLk7gX40Sw/3w5N3cubBtqRA0sZ/CpSmPB4gNjwNhdQ0u10q7G8yo0tt0eAhV0o1i
1fmRLiGpjmwcEUwqhFI9jpaz/td8B9VuTuZ0HkEtIT3qfw+yHb/x7xYgjyCLlPDk74TJbyumqr9H
8+aM6KnHyHs7IluChVp2BgAf2IN6xcTUVHWIj+EFtj3TeZpVo9SkIzlg5Dyu/KgXy+b4Bx4QBDMs
Fp+eyUbxM8/DKYEriQNKipk7s07lAJPXIK5mTw4OHeHjJC7jhszd306GlqR2B425+aTNNWUQd22r
++KFl1cTQ1uPHzPb8QcQmbSMT+y+9YNEXdgGwVxk6MYGT7uOa1m3DxdX6TmnvzgEsUEco6XANd9c
jbJ3ksBd5M915AQpbUDQHXz3GYQh10L1QddnBebQqoh2RvP81euve45I1TUCsrM3afDpJWPg5Qlw
lwoEgNt+xfv9sPZXIPJN4gG+GUHmdAh/RirTeUmDhnNOz0QnR5sSqar4q4OSZZQoj6ZbN6o2brF6
8NilW+Fad5L17JnevprKBnnpW59vF93rBlMp7IuTmKAj7G/lu88vAWUbB5UUOF1Fn/myS+EY3hFB
7fqng9WgxfxESia/e0mTJtsEK30M5eFle9djW+CxX+WNyz1hyRH8t/6WoIKUGU9flDJRs6O4jkSb
FpVyPjrlWRkrbh6asRTXgedNnIIJDtEm4hNDrD8dKEQYTZLOiX7wGfFEOab8Hh692VCuLPKcLZR3
WMZ7xdnRdZOePmE2pTUjlTPpMBUokT2TsCeUipg4eqF3Rwsos3Yeik5/h81HTRR1vFdtWuFfSYGf
8/KTuw+QdeSFEjGohCinLrCWDxwsGrpIYrMcWMpMrKKWd8+FE/PvfQ2OT41D3tpJ3h0dCivf3G2o
nwlgfZikVQDi8F/vZ08c7JcvwJLJ00dMRlZuA7G1q01oATM030DOG0BFkTSnt89/HFJ9qRk3oLXB
oPFymhBIuIrwwcCXd1fJUUUFcSsvmwz3Emc9EEsPiEbi+p86y9k97V1cf8IeMjYZiSXhJHr311wG
0XaSdJvSYGQ7Ub3LiXYkzwhwJqAd4gnnY/ctXhGpiWNhRC8lO52SysuZda36qDSyRrEXkh3qeQiG
h2rXWeqVK7elFc4dL+D2JBjRfbsG7BIeXbYuk4J2wMkkaBXkg3DHGRFDPJc4FsfbDvgyw8J+K99W
QQxVtRItUPa0kC8/C/yQoxd4X/VCFJ47I9giNAclFfyn1gkXoGmp7P3JZpbboZnMb5JcCkApgrgW
AiTNq14c1kMXoKKnZ9l4/xHPv48z+xP0ITOx3jX4BLOSOq/5Irx7nSo6zRrmKkKIb1ZiprFiAWbw
266p1bZApqenSw17I5DmB3fuY+gKD8HMh/AihHN1R7iqh/hgp509InTX006XrYHtqIcxH7g+BVzX
LYGH3k1kNdMyxyicfiPezPI0P4P24vyOfF/SDJGCVOWM5A0t2q0njpbFqqm5xjSwbU7qtJqBiIal
Fpt3gjKav93xenbcWmWT1KUDBnTXvGCKEvxICqYgKvu2Lt39WZq8eK2vXrUzWvwKk7eXgjXvO7lZ
1iMC9vhQ69ChUx3n7qeMvVd56Fv2FkuBESa2s9Lj1lCUI8IC6X6Sm1tpuWXfMwt7dtqmv/T/4LiU
aLXdTRT76c3GHen0iXC2PaEtFIETCtnFbxq+24wqS0g7v3Aim5ZKWtg7Pkt9LoShZImevSZrqXYn
//256uFUZqdQVMhWg/hVvcZKaWMh4J96NItbu4Xk//ZHsQSCKwOFHz+lHU3NlZOTwf+LzpL5/9rQ
GBZeTHqMn6jT4G61Frp2D4XcAeygV2gAKbaiYyZ5+wx0XMteZpqL3kmKbOZ0qoRRfv4ldfKKI+sP
4CmWGsTqtkG9g2BBvc7KJjq0CC3mE3gIXsQ2/wNzo7qK86x2+dcA8FUIJ4Ia/4C1ya057cOt4WEC
4dEDEDyDAbcp55Cp6+Wzefd1bZeBZhvt7r1UBsF4H3mHQ3V6NF7WZsY3gL6W3EMhTN0SsglqMCij
Iu70jC3wH1TJP3LtVKvR2DAnL96FQ/Y1OyhGFRtt088QCn6pYE1/Ciu7e+OGZP2zFHFEdYSdes6D
9Zo52GpSL6dZJredYZVomGMXOoLZshg9Rb+cfLOYoU1oY/4/nfK6SotNBoL59H0mLFnZ+qHm1PRL
PvEhluh7tbJ25CEJm8VI9njnIugkD2Mir6n+xa3uGPyitCk/zc8HPKITj1hONkBZ/EQPv7uPZCeS
TIqDQb7WHblCYH7zURK+Ih5Vl9IgoSJFlfMzliPS6RZ8P/iktb3U0okUZk+gAzcvxoONaxCv9yDq
SZT5laWt3CIpZo3cNZgD0KGdgjhZnrgiDYYxgzBSQMwknn3+pl6mVkaiEJt53AY9ysb409zRVMSn
xhLcvNBVv2Z5AkDMc/5vudiKOQs1R2XQRUK/iiu9Iy7k2rGNnWMx2IAGSGcs8Eu1WCnbCmMSZ9Xe
pGyaQjYijljIKRiQ9e47xas7TfTrQczm38esKCW2+uKjp7zMjPzVpR1LBpN1vxTZSqdT3LZ2U1u/
wnniJFXGijOlmXYCykpWfjtD38TMv7920hbYxI/t20h8QrEc7biN1FsbhZL4nJV6azIDegxJ6bgW
0jf4vCGVCbtq8y5To8ne2i16K7sLXc9mP3Qh0IjAqKrRcCpWUSfOQp4gxCBi62pea4RIbuUSOHW7
ujNI2PkqVA1hRLG0xZpiq1/NUrQDHklnlyKPPCzavLwQb/kHCRw41AkjqpmeFJbxNBNOXqYL1kZY
P2VVlYrTmnrdlcTyRtjsRx77JSyIJK2n6L29+AcKt6xpBeoIjNGN+a840HMRuo4FSAbOaZcaKhKe
JfGkWVNfMYJH7/XS6Ynk6MUSWRzc4qVs8wWcMr0yItRlnQtbdufAXXyH1NlKnlnURVNoNxBSUsEp
IGCoGKAUKPPIItbGZbhRyGpkT+0iVIRkqLNasEJ2J3FWE8nLyijB0sg0JUMuKlZ30kDi6ITwFA6k
vhkAtyOq+XZ0E/QRIhYtU+AOVyXOB9HDF59PHPlR7CGXZdMoOMvHLk/SIY6ajofPQWQMdM+58vz8
/f/tcgYcfS1CpFKfElUInY+JicVNsp7b7fK8a1LUVOkD65zNWj5kMqK/SPcG86qS2GIxLKJ7ipz2
121cPLT6oWcMOdIl0n0n9cKbKek5qfaAoFmVL87P9DZsvjLJX3Hc146i9UUYCqb8+2wwBmY8gTBm
AtZ4+iuQWWAGXlLZ4iECU4nDYxsW3eLW4gU+4yc0fCFPwC/PPJboSpDTHnEm4Gh8YBypQjDUKoig
kKQR/m65vGA7S+sHqWgckFB0EJg0ot6lrbhjdGLNNX2cS/mDeAq8rF7NtUAYX2Kvr/4cgrqSfeRB
F201i6WE54lrvMTmrRyW53BNfnKtZajo0rRYQlFiEpDdZr0L7G8DdoF7X2VisF/HqAY5c5QROgjS
jNH1+gXQZn45rbB88S5wUGbnzN3YpMmYNfiVL9Btvp4OTf/SFY2IA2+gY0vHk20XkLfH7k3DqBXW
bz9l65XAHR8RXojXPvF4VCbM5tcFT1TiYHifQ1OSvlSWGV9FdbWKs6Wq5fINw21hekBtxeYaw36N
vOakgeJ7bfQvbdt+K3BqmtnCfesjFB/B9ykDsEcHaCUzUQmquHHhtTQjr0W8D762QK0UuuNZwgcW
uJWQxIGLfiIwE6FcleMRLGy2ahE77zjrpFgOmYVDSR2K9RrByyR+yEnfwwxNozNxiIM8912l3iSM
qvQSKyO5Db/g7HEpLRqOEXuN/JnuomXqLxj8RMAjz5md0Dr1/T5NJ7FeAOvWhAJArIEyeM8JKm7i
97rm5SxDUj7+Ls3lArvwL8bkSUuF+YQa9ilME20g6hOLWyNt9wJeNT3AuwEIWr4bXtdpIfYcIDAI
emyCqexPOlYeK8jWmBskImq/Yxl0WIj9N0CvEWh3guk3rTHmdhMTWFk3q+94aLzkH45DlWnaQQEw
P9k9G3qFsp/U5DOVJvLgOLQgJ4x+vvQBJCEvcvdd+QEKCqJnb07TlYQ8zvmFB40ccF7Q9Yd/c1yO
jRHHWhJydvT6+fpKPfgg/NHAY2Tgk5e+dhZNt0WQdnnwSSwiv6QdT4FSpVv4rvP1OP9r4UymxZuR
x8ODV53eX/XaH+VBRvswI97FSJ+/k2LtnVVLmF+zF10YijlofBdIW+tT5zi+Htf36QTjLQfFPbaq
4+fl81doGj/GduTEBSjWZ7VOfoFzqe43IyjqPF2VMe3/D0+KIy7IlB83u5SBd1YuRuw1JuDemETv
KgNvfRLfVGBmqKoAtrxzxALym7cSWHXy5eZeC7DKaSzWlH8JdxtY64PAx6XdJOHHQn35TTtozG3L
ix9mdxNpXd/OcFTgle3Aig6R0GDC+88oCpO4qQMRTOobOQPwdQO1PQuyAjoppt/YBLwMMfug2nh5
Yn923kJHZYXfa4MvWYXTC/fl36E8a8Yxx9iQPOTys/HgG2DjIPIRsdp8Zo28D2AOTrsQSzQWA0WN
TZcEnda2N01zCoRkFu/hVz5gOIjJ9uCOG7lVQ+zrGGdU5NZEGNFXdMFQKb1eTzyz27bWZnad6IaY
GNrSy6FL2F872ZlgEfgY3twy22EkBVaUVIZ0HKkbiOfTOGw1Zs3LqTc+LcvNnHkGj1RUdda7XCJX
nhhjz+HWfZFmb6P3/9tLVi/KASuRAOxs2ahjiuY0LcEEC5D3OkYvNJVK1xnzwfLjQ2DWxZzBiFg6
V2awJwshroOp26VeNfJ9igBTVgxtct6elscRMx4/6zC4J6GBLfaoNz7sFvy+lrQ61X7XNUDzMk2N
eNVs9TDSmFX3pYhbAkX6BaKdq3Pmzxwm4jCWwn53Ww/o7HgET8fkZHfNKFLZhvT4HSefcJ7W4q5f
dpLnSafr3JW3BMx9sfWTWXGB36Ex6m9LTGJuotTxZbT2uOP4mjC+t0Ml2ChGYlkkQFADQYCGmolJ
fRwpd4b97dDIrSKZJhUPStG+hYTyDSuY168nKsX6amR8lQ7rS6CZqb8zs9+zGARYLqKnbmkHr0DK
CyfoCWAjDUobonM5wVHb7YzTKBaHkDSX913scMnTAU9xujYDFe9oHtZbRe6F/biYOppY7koVNoTi
EYPh5krOIC22H0EnI185zDuA5Y/1Hb8zifH4sDsVPaJEmXHwwuwEL3i36vdnqosiDW7dIPhMM6LS
rWpTP+V7TEhoBh2JgSguEOWEHJtaznLTmsifJ0fVXswrRcsu8o+x/yqLpoKlweYLb0Kl1NYNYY5X
SnhYjzo+o1HefilAz7iVqbWNv80lpU+u7dnREF3tghEMKp7vI5s3pXjJuLE+zqwSLtyg5UyBOAEn
IFmiEUI1jgqMlg4nmCc+tGMFzE/7PxqzGo6MQrcm6uoVh01QXOd+O97nqxdQMYBTCKEEQin8igDE
7JbpTxoYrzWY3RrdGlp3bAAGWP7f1Imj8iHz3VGovBVHiP5jyE5rxySAj/txcbjMRfQVia+mUlNv
hmoO34NNgpy0hK6xgD+4VqkNBclnH94sdOP+O4JtGJ4XsLxv68V1NMBT8+ZL+o87gzOIZkdfdbKq
7f5geg6KODwBv2H4eFebhTeaFc+U0y/ZAwpOLOyR9jm0zHQhc6sZZPtVLHf6iw4CZvhYQzJhSldW
zWMWoq1lMGLMIbMwnYh2Xbzw6WEjOXzWiTgAhl/9v2xuHrnQoJvw1hyTQWDAirGZvxlhCpVoC/Q0
kJjcvRyrvYQUp6EGzmEHXTpPz//Y3mrE3mD/MMLcgNmona48glS7qegKxS4C5Mym95FopEs/2kcW
qHQn413/aNo0TtEWRcWERUGDf4mtKOFWvgSvBvQud1+PJavTVrqcPWpHelw198gT46C4bjqxhM0g
VgnVPGK8+SO6GAg5LG4u4rtd3hXxJp8dppy0uF7P9GKA5Y8OkdKfomu1MsYkK5uuC3AnwSxRMsOO
Ukqkt5K5T5uls8kTUO7wYfVO03DRGeUEnF50urdpawReNXYqlVFjjXIZZ1XqfeJN9izQ0R7j0ZEJ
KMRZF3j0FNAktQIM5b2ZKnRzlLFyKyga3o0rPuj67wt0J3N8mwPlBh52jD23ZePcKTUO6UYId1CB
Xu6vC5X6Wlnx30pV4FwzqSB2VgDdw4H8KmL3ABV4RN9CpW+LrqcRcUbXVPGvgge+ntaFZcfbw655
grL1OqmybxiMZ8qmldRLtkqSDXpXyBW65t8bTXw5UKdhIwqR1cCmFix41uky31TQ30blfGSfpQ54
aaN8JrpP1rjWPsHMKOaqwfz630fwe/AYBUxjg71A8nG5Q5ipNsL93Y7SwhT5Ow7hA3H3v9pPcF5a
syHYYA5L7K5Sqmxo74KSL2U0XKJxqCodoDw6blpXORsZ6wpfi4H4bEBLa7kfXUIChYqsYN5VrMBX
YyBj+B7jq/VsfWMGZDRB2MnsPzxCCOTkn+Zs5hTTzndJfsa8vAp5zXHfHaXSb8brP0fHYZTCdjBz
RUBIaFHZloSD9E6eLdyGc9LSmsGL8ZSsqAbQHPHu1cfs2l3UzHuYG0VF6pyaZVkTovirMeAVLNrJ
GsNk8zijX/PbbYXmfY0caKttTBL/gsZS6Ve37+13XwP7Lz3Li/imdzfKX49nDCuZeQQM0RxvwAVr
Cx3u52CEBE2b6nrANszkfQSgEgEbEeuD8ZT1l4QuxUU0F4Wgd9LOU0OIvmz5buzotOsfpOp40JFP
r+CfIsGDCPPyuHovWqlJg3yz0eP1nBJEGTg4d3rPA05lDOUx2d/5zKv2PM8YGSEpWPkJzRlr/MfL
0vqxnF53aKvvYAWKgcIvqsHG5Ss6jUXRFmUd/FxgWKQNCitGwiSzjvP4LUVM+MpDikzrLiN3naB4
KTPdqTo+6/98OEy9kDJmcP1aY5VbzMGBuphKThTVvgwSg3oirVR4uey3uyxvRhR+DpsFzl9Hhyy+
glXM2GgdQkB+Qyy+/XyKihZqr0a+OGw5z9Cx0Z5CT+8qONDjZOlxjjRKXEY5Wsi7V5NDdyB1XiBs
DBJwqXq5ZT8dyZx4hYCSgs4ADsmEJHBgvmCcv8YGrhpsMz4nFmjhodbrLRyODAJDVCU/JUeJ37VC
v4tErQpqZrfg1BW8mqFJXZwjJiv8NE8x6Fpr7yBoDqOg4xUPQVruU93kgHlVUQbK7Pfs1RELulCv
Efucvh6kn67qnm9OumhL/ig15er3aGTmxMq7ea15yPiK3UAbrv4yvAMDvWn+HQeTB5IaCvQxKefZ
UsIh8Gvw/I/94RwFZVZpGGKnxkHOf9Yx9LaVRbFNrAr0WxSkm2SlgoNOkjnVuvEf1vXkY+WKzIvs
qEkdC3Jvjfv9imo6absBZwqBI6SKGy7jzSixbIM6QB5cm74pbd5i6OC9blSUNjibl2aTIVg/DPCR
yOxL6wRUXxnUh6dyjAHGEDVvC0w9f/UZJsVxnYPYncsPhz2TucwEnn9mmOerp3lWYLyO7zmEorMf
+JQUAocek31RYB7EfuU/HoQo0y0ddyMljn20xXoRlZZiOyXuiv1zro507ocToYyopNe9NeUam3kg
ZgVjrVaHaMorA9xIpjJGxpnMIIn+kbPXuGzFf/0IlCTLlO949VUpzpWi9IwbXoY/XWTjNGhez2Mw
C4mmuH2z7BpQvm9Lg5/KarQZYIPmQEOJvq2EXy0S1eFkG0MYCdqhRg2jwW9pmoj4M9gR425qlnWn
g4QpRtIw//sqv6B6A0wsIM5jT/0KoOSsisC9AhJ8TeqAW/gf/ayVFQWc5UogBHlznf3e0t6l/HGw
Gpr4tITXvColqaYlEGa53VDK6d6yjNzCwNuPEN3qvmHHNdQ5OsCkRR+Yhs8c6S7Nb3rVv7XTWgI5
TTio1kNEwN28qO18nrsuux8dY4HW/NUUhJ28GW5py/RGw+uFHVxuyNDkeWtTun5yqhoDxHneEsrI
s1FdtV3ffBxX4/Znf97+cUbcsMKKiAZf6h+GKR8ODgTWoI4trGuUXdTCbENYT8e37fR5FhdYBYbV
jnTpigxT5p5LNflosymjHdLOhETLuxz9WjHhW1pRrpd5uwbVdzLhCWIJX4S92JcfwJpUM0OZ29M2
jzBgbK6AxW54OdCWVbN0qfmoank8TyTFp4/fCK3rzkkadbHfiyf8OQb2VgKYOLPuJevO9hR0mcC+
b9bAvt65JgmfsldbxnffpZs+btGeQe61WV+NOO1Mx3UAj8LtEF+pGDaHTDWMDrLyyiWCmys3Xgbi
5jaAcTQNWBGo+y2Suych8M85nfTIIpPKOLyvuXV7YnPYnRLaG73F6Xuf+8rqrjJm4F1qZRaTUsCA
TKHAB4L4Oj2C282DE4+6mvJNWUX6wS/CBasj9X10cEhvV8toVIJux23uMfUOakNILG/etDRwDXPh
2ymi4W9PZlT8akw2xbqbKf1kswAgw9jXyqG+Khpz6YGoZPxk2ZclNUQw0HstU6L1nqyHe08BhDsV
wsBJNEx/7vYnMXPCBV1JiHN1OPN8LM+QtSObUbrjyLdk7mYWZZncqJH5MuTm3Eg6fdA/dMfEjA1S
kRloN0cFnGBC5pYvOd8naBR7mrGYsW9n3rcaPYDpPBGsQMntqfhnS/Vpnc/6BmztKffmWZidx5gw
lO/MUEL2akoS8lXVAdZFpBiTdiSWf0y1M0g94k2XcPI/msPcP1wUBjCXR9HUnAOPaNS3JxR94ndU
l91kZCGF/rj75yBI3KlwE8MRcz0ODwuOLtA1aCcpOmujF5u359fozzslg1eQHiQxMe7Q6OUwTHhi
B3BzKws+i/BKEoHmvBxSHfEz6rYo5f/LubTZ4Do3OvFYpTyD5Titi1+9n36n3OA3O7TukKM2P27B
NWFVyntwS2ZzosmhydbYMgx3nRNl512F6SbvVDLPEKooJijPDv5qc9PtoLV7wwWpUvFB2+ilud/g
j5t3Kx6LKufKwLJxXbG5ZFFuK5a5IsoGo1ARSSAT8Uo9rGZ1/dE7lwxvzHjaoKsu220YA6IyCDSC
B72vnHVZWohdUS9jkSmLqOUAA+i5DxpnQ5bkA0r2MkqGlOlg+clbXtmnECMtWDEoC7VI7TEj7lLQ
+n99kt/TDE6U1IMM9oO9dlBk1327wM0k+wUelKvxXWvJKghdzEiASzMD55X4oVPXpx4oKqiBljKx
8xfJVpU2m0Gyiyaqae3UiwAQ/JdiqUWyfAw0/FUEX6jroE6ATEa86m1xpR5PCj07YAaivu7F2Kka
WbBgCCO1AjLIBmj5CoNC1qfiIBt8eEwtpbFFfOxtcrRZ+OylY4rVJeINMLGWm+hW/5oorAqzKla2
qERrnWx6RvSlxuzRprlUg8EnQlh7HV5luQy6H2hS1yvB2k6QM29BTwWuXouKMw9ai+szEOcirLYK
Ga7wO+88Uu6n4Y/TpoIGUOP55XChgWpKd9qLaCgfWvivuT5gMFt9ZzwKIS2NgiV6cFErb5rMaUAH
GJ05sIjW0u6JX+RIlPp0kw4A+Cnv95OTx0JxHvBbnQDoOo59qSENgYRzzyPTrjSh/n9zj1/58HEf
Y6FlIvAlwiAEJJz5KxIVZ5l4xOfhqT/SVrnMfcb14qg0C+/T1aTgwtNamntnVTDxnMgay8B/SekT
DPEXFKMpB3NCyxBWrUSnZObohEUTEpNuVycOVfBKwWp6GZ/4CFMAj8mzjcrMTx5l8K2rZA+xsl9n
jhvZg+d/b5IjvBzl2dmo8J6S9NBFF06F+OPzEoYdc3j3mE0KbziwoUQB3BzbIjrTjaY2umeqNnou
npbLSwTW675oY2dBI/NYBJa3XW2iNznlL3cPbCPCPJZ48X7lJwFzZWcOBe72unseVlPGAA8zNd4Q
pmS8MpUqLWJm02nUpVRewtDIV2IkadfMXUBmz7xQPyxnT6v7TNr368aLKs0yk20ni55EUafp0SAK
ifOMIFNP7WnDp5j45GJkPaF3lOQXuVND335rtDn+mUO0TF3x++Qywlug41VCQTV/pyzaYw9qGk7i
LGdYnJ0vxKDZvsdkZxGRruavBdiNMm2+Tbc2b6c+bQsaw/ra/8eQoOe5upcupG54M9iuRq0Y9keU
mmuKxi+135/gMF32mz5zRwsdPl3rty9KOLItANBAOE9qheBibZ1ODQ6sK3DXNXmmuGg1k5MLADV9
5+Xj19DmITYJWO3kqKnTUKN7SkORfyO2vBxPqtKKl2oPqN1cSxA5nulLOhwpxDcylKd3SHyl6DwN
hANezE4ymNBKjxyP0y4jkgRjCmls72fcjHwKvSt+G9pG0kRCqNIv0I38fF7Kl6nkqqbh8tXEl/Mr
6K9WnhCaBVrFfG/l2VvJX+kWOwmvDrkhJ3ZiK/7oNv8CSuw+4Y2F5In/jLXBVewcN7b1Nk5h8GeO
PgSsmZIBdYwe7Nb7UV50A1FH4qaJgGzHrf5TG3zUZVt+jtRO9qTvp5MAiL6hM9K4zSRPwcafPhim
ZeBLsG1LTsxrfMgiF95Sax2n/WxblZha/wfot3c8EMJOQXasPepC8bwLkaFzQX0cKHQiaz8QAK5T
EbJL4QefOmU62IohN10dRPa8hikwVWXBOKWqQVhFEuqanWERJ82GY3bqSp2e88oB3zrhJoY+Ma4y
qzWY6/cKtp5Zgx94o4rYuS3op7THWURsWvxxfyvF3F+UrBk6LrDlZC0BsP8T/c8iE64UWYzOaOip
7/qbIK4wDKlFAgX8uzp8j0SLL+MMbujNRVh1emibcxWcPfqwHQIKxmNQZtboCL2OfOfzYX+QeJN0
BtA/1M8dj3GTC2Kae9vnQgRTwFzDehiRPlprnUbx0/q/hhdvjPADv+braDBNs/XV7c8Pz7fzaz9k
RvgL8pT7/vEUHXjUnBYGKFPmc99sZNhLl6j+THQ+x5OLvS9O/m/RYuf3E0B2fqoQcYbWoY9ZR40m
ZOQxKHvEz1FX8q6+24ETYwgS7L6qGUbAsI2/bk/IlVK/UgxOeDUICIInuKX3Zg4id2fWcdI9P4JL
ZnvuW0jQmFcw+dkYcqJN4bTqJu1dSVdf/307E/5ajwEUtAqpNttuZ54D2DZFjVcMd/q0BA9FOZSn
pbs8YXgHCHS9e5iA7NxfFbAZvwV/KSGJQZR5FBc4zo0XrE9UTP8Fz62TAYR+Cew+OB557rLmKbCg
SOVlpPhVCVQTEWePCZjhkJCotVSG0H8hZ5+IjKYQ1Z+F7Pr8Zhoe6FIqIPTYcKzU/CtHsTXEnpU7
7cndfS7R3tA3yUAqu+CzDkI9qTo39d4bc3U3N+tSvBWII4rW2Kdi1v6ioale017jQZZ45k3d+RTw
uIMu0Mrsvb+WmVUjlNPDCmZwE7VHzld6CWcLPCvUCHtdDE62a5mzHqVkNi9c4g4jJzp1Q5VWOAdm
iXTs3OVQWYKajaB893v6Dz/k28xsdDDzZC87RZ9Vm//At/HQNUQ80FLjKE1RA9IdqOfYRMdszycC
SHJSF/NyqxCGXo1+CygNfZCovoitipdACSZcevmmDj187uL/nFBALzG/bP5t3RwfbmqpqDpMCWLF
Wmm9ByhSkjdyAU2MC9y0hLrNRJgwK1n6h+f1tUDllf74HLUOhbcxy/7sWDVrlVefHrawyNQq7NYg
6dhSIzqbhUs3WRR/L4Jvs46EVu2BjU/fvLhkH3+C4vAJ+66cQ/TuFsgPkVVit++ONLIyRtvzN0t0
7Po8D7KHJpbmPIC3Bdgqwoj+n9O4PxEvtmILUUXZx5y5FgeZB8uqzeiUqIKq3nOiaTbnbkVNXG4P
nRCmUd/AoMKEq6emQY/XU+m+m/h6T1ifDvgw6q5ygdA1VBv47EZcln1ucsBeO1t9J1FnHWXhcBgG
2Q9XqqrXtus8st3XFKxjWIhBY3s0n08hZIWCgobENOGk5J1dd1xpSnQKjguNNcVXkShJl5fCqMNv
VH4pEozfJspeLjFxnDuDJjbSphrhqDDS8mZ6CD+XKYb4xz/cqPYkcDk+jrmjy054D6ys/1hcNVL4
jHqTMGhLMyNDjd/8iTJ4ng9AJgAuit43ITsFLMdJOGTDvDobkKGtO2+9djGfzD6XsDw6zEtfg+Hy
CZWDYNLOkT3MzK2WwcSXI7aPsc0Rj+E7Q9nJaJ1bwUdhrdppV065ZOl5XCWT7v2FsjGPObzjvChM
hLFRn2qfFMAdiglluQyk0uupMB/j9OM8MqGrCBPsJbL+0pmz/VtqvVMEYBYeKoyUPvBSh0uSTSJ7
I2sT4KwrUW0dUNHfO+wPo5f2I7oikc57SLe4NrsMUuaASNO2RLN7c+Vblyb2QspuPdoe+hIkEBAf
zwv/di8R5Wwb7iSiLUXYbq3Hx2nhvQQGlOdasIe2LZDdPBOG01dd47NtQwqxCbwRkpZHbH3K1r4d
MnwNhP4JLxaqKHNVoj+9LC9Lw3oMOZEEfYNfZzXHDyCy/XXuCK4uANl7k9+o5xzZQOFt5AWl1l5Q
zBqjuvjewZe3o3C3/FlFcmGQQZgTLYqKUudZJ7/wXo4xfFZcf1ecM1pUNDEXXJKttmMh+oOYGh2j
zRO1KUsmqPS5cQI3Lq6htp0aR1v1Jg2dQDlSUhH56ksujTCL/bl/6QHuMuKdp8nkzisiGWYJFJ8A
oq/NiLx0kaQPAvDLBNpBxabJWhBkf65XtXaKf7Ur5UKlQhEZjxUNko9pNX2B69QaAx6ZzE8dAYf9
2JOrQqzvJf3rPbjx5OG9A49shZcWyuyqd90k9iWtz3fFli/KZtVLvemhFzKCjb02K0zwnnYlN94G
UoVDBuhP6uyz0T2H950GXdzs0FUZ4kewmJUenWDUoMViKT3OLzhTeDk2SJFb1/ONKpyZ2O2IjWrh
AcvbzpgaHpyUBgbcvziz3MHNLR97zhfVSfJcnWzoSWRW349FiNmFyKV8zMSEMlOtY1CZNU3M4DNw
lTb9eKYRtnH4SKI++EzUfEVWWoqxaAGNBRhaitwNHv4QPIkbuQD/vc8jU5YUoChNPNDN20svXiwf
lPSt2r77/32jY7WtcE/3z48IixXeWYnjWC1QY0ChHkh4FJB4+vljPy8xe01Scj5R+POv3jYL9YrS
3KpBPV+zbY23twSnUOKyvp1NY7Rb9HwYLxqvMu8CQbjV2DnZYRytGKvEkaGSZdFgtl8ad98ofhHw
QSJpi3WS73n9s64os/mqgm3y3jijzcLKoDDqJQRvxG5whCmKyqoFEKGSo1ZALzkkOZCaiVXpwYQs
9TrNggMD1sBM3GOf2egEdBZnFklT6JVODHtrTZFz0Z2S0xkuyhYMpo7DtbWGHa7vwPdiHjiOqB3x
jvxiCMOfVQPIiZNqY4kc6OBkUzINEf77+Xo3/jkbdJP1KJcR7HAVDJiXQbdU/hVFoipb0P/lvKXP
7PBtJiv0lvNp6U9F6zL1Kbz+uYLGEExqDmuYgEWJvZ9oF2RqgngCtAVxLlIRJ2om4h9EGTjjsFx9
hUN4slqZAlxgPzcvGWnkIsVkGyUp46CzKKs5VmeWrPJaOHHPwP9dvpR+hnh+FF0LG+1SSRIxftOU
tf98wRYSPpc/KPwRXEvJRoOAQEOnDcndFBsJRkjuaPWYMPZ4A53RN9zepV/N43gh15yZL/WPMmDS
lWYMGUkaXkKQu2P8QMzL0cZtdHqMIB7Vqk/r/4pEI9N85wd/JeeSpAqgmY0RAd486aAKnq3GK0Td
EA9MH+w1CgqTL9VlNgtMe23g+H5NcM7tMmPKF2tX18jnItIhqPDDQ3AdpCcJnEGg2q/QuOh1sASK
TbDKLzbQJxTt+Iq3U+TqcgVfRWUWObcvEjUIfPKiTKTL53ISFPnoUxBvIShgYxthwW/KAm9u+d7n
9DRs9WYp0TMHMpyV2aY0EAq3d9BAjxm3Ef3qoK4+KRcy4XLSbWpDjAHxnPS56Yg8KAhN7i2so+Q9
uJcb5j9jW617coukiY2eZo11fvQNR6LbYqjzKaMmjS6U/NhPZ9fe+BgfeUw7Inbzh3co/+54ei14
vaEsLhoaW7xrg3xn2WEWAIy7fvuaLNUISQ+yznLvfkwy6n1BdeuS55NKY6uJ3PGRi0GwRaBmqwae
mD4Itx7xD2ezsoY32/p8x959/TH1RgtHnVJC17dqhJfLV8D4I1yE1cDipw1XzrmkObECjUWpBiUk
rQEuQXvgTqwDMe6MBanJVUllqq3hOi/TE4ua/nvxwlv0+fHLpHDMZdhcHF01pZNNDfbbEnPbelk9
HaLF4OGuPIA1m9eZZObc/IijvrgL3qok0C4kaZi/ao5VWiHZIv/MGzJAsRlYzg8PPJRdRmrvQI11
6t/lmQSrNv6jmSFkgpF45iGTm8QUuolSFPtvEgdLZhHGcTBMsYPY/5IQ2L5KGm9o2zh5NSwOh/Uy
EUDn87BNB5iYa3acLSiZgS69WO9plecdb8SSHcTDIZ3dqu/sh2dfoB9am29B+E7Qb1CEnu3caGgQ
R/+viPfspW70Bhim4BFtktv92BLxJeo2Rma9GqId5WBmT7a7ZIu2C7G7ZdQPFJFlXStBmjCk5Vzt
tDTecq0mEiUq3eNxQOcG8w27t7tNMRS02219SrzxHXqzznteczwZEYvS7/N+sQQUQiHojdJK+Og1
UxuVGGoMV81n4+osRUz8cmJgiPFu2GS8UtgvD9A5Q85yCljwd0FXI7fpIUyU+O58PVcI3dY0xEfp
xb/4sy7CE3TrtCl6hntH/m2nPQAEsLbg5RYs2hU+shcY4EML2V4OaRiONlpiXrsBwS/BDYufNr59
o+iw2JTzLEoUrHVbOCFNF72TKvbVivueJtHtispZMwR79lTwGnflEO1jl6adt4AWZQd1ZIXSzvex
IslFks2SBGQE2nBqs21VNxShTd+n5JW5ang22V0N4gZNYwn5yA1w80ipHuOdkv3fYOQ8FuX1CQ27
LTFBtmsuY7rXAnaTHB0w6iaKMBguV6nJLSDz8YuInw0TGi8tUiVsTykIYMPA5tB90wbGGZq5pDXz
GicfgDT7ofuWqo953eHCJpqL+ssjyfrh3zZL/vdesso2pEmAd11/+n1TZrbUY5myFFpQ44tb6pWH
PVFqPpPRtGRlVropQgAxtN4MzitYOwb6ojQGtkbUzFhXEnj6wQjW3zIHDR+YA+WcwrS/gPSUAqKi
aXJWEXG7pm9u/+dl+dGrvAr9okyR9XSCtnYSI6iOIeF19NLdGTZczgcxfyzYpOs/6GWkLSMCscLx
jSU0iLQj2hXWSJZuV5E9pndQ5HKCykjtA35dbAef7nhvC8dGVkMelLng7qLoNcLLwebhLB6EmIEL
FOWlM6jhCg/6M/TgjNQCfo6IF2rxZDKR/OfaQNJt8x7Y8eXrh+/vKmx9oEdZzzXtGSIje87rMl8f
Icl9tIjwHj1GCs1JTOFCNiGn6r9mAardGva9WCEER6G4zET4rhnxLg5NQfkXPofUXwPr1yQE2dAs
r/eLUIYpdV+OQ/jrOTfmSj5OMR59XnlP3i3wWuwBObw1W2m1oTIABwpR1FARu//2mvaQKV+4vy2u
ODjot9TvNVa6sY8AUN9/lf8RQ9ex4LfRs+9Gwv1+EcCZ/tLv0foFxhNXQuAwh9i8rft8Hr6oyXDL
ilnBXDU8P6mHBhCZNRRB5JUDD7jxtKtY0kt8rjECo7Zm7F7U0cAyNOkiqDeWtdDbNmoNcmEZSXDA
voWkr9nflPvgJgajtorGfvhPxDMJ3mqQiPcbQyw+z1yxWGR3TFa2nyXGnfh0T/W0Jrd4ptxJAeyH
T4Xx8StjoUltumKnfqkr7IeO/1yabtJBrogEsm/4nVNeJv7B47F14cWwYAbKs+GbX2+a8BjOpRlU
fjZ+dAa4bGBb366AeZQIFcua1isP8JfckfyqPAslppob9Feww5jkzAnmfQ61ru5KIpVoNRbvapuh
spQWwkxJ5uikxpW4pYCKDQQJtxsqHleTqpTk0u+PZrsHL8Z1pDocw/AvJZbEeqo+pKf5s+3O0/KP
xmKqTQe+PPwgUlXBFrLxYuTuu8J1qbGxQiDimPU3QPfGnKI58N9oGr/5FVXBQmiiERoDR7G1DGpa
1yz86vr7hIZ6pqtBY3w0cNvSmpuBXVGu2TgoCphN9FkBj7bzSFvd0CZ8qyoPNG/DIzrgO1u/MhIt
dcaFNluN5bEAi/Z9ggqVfKEiv49LLUtXVkpVKm1PgkomiUEVjgnz0ptHdt/7zC9kS0NhNrCD0kRj
AfuJlQNyoYTnmkLd75eF3MBLDPnJpUeg7wfOnVpshatFDVyonuh74lbpuGTOwtyfw7EuE4pPw4RO
2nJBWqh8BLMtdPW+9S9EmuZd67BUIkXgBJMqyvsjL4WjdooKWgsFBsAcHYzUd5njWMfp8zj0WFk0
o7v5PR6bzWigDcgXaV/fW78O8FQYrgNJ+G2f1NZ4YgXtdICGnBZv+LvH5pwhBQYFNZI++kw9ZSxv
9cIMpjJU/e5AkQ9bxOCIhiejD+5uNz05ei4YGPClgJZWJR3PQ2Qn3bq9U5TkUvUwSsanm3/vUbjC
2T5McTYNNkRigplhPKCbNyyFfBlTPbG2F7YWxgHeUGv77BGdCjVBMMSDheUsUGnTtgyyI4PUnZ1Z
CZbkj7nZadc+o/VPiivH+/mGxkp1gvGJzdbudm+DPX4yv7nThNG6evYqCu6SjBQSnD17LfMPSkGS
2zHqyoM1FMPKASoLiTkERf18+KuQ9xzndxVJYPcSzgta/VhrwRa3kgM9B0n0g4PWTRa1zVWNHffW
KI5wXmoX2MifDUBIg/jHtwCTJcgsqzwmsujEmxHq/4p5Cf7v3GU+heoeaaymGqA7ErREJWrsNzRM
+uJdjYXEYuIPT8UQWI9ivcDAP5K6A0rqG4Ibe9MNOiprmGxY+1OXCPX4xbRi54M0Z2twno24kWRx
IaY9dSzEbe/gIl/nE7fI0xUvNPWk28v1b4RgxjWHV/sUw5gJ3U6mxf9yrtE++EPqt6BrM8J34vKi
/TlM0V549FIW2BVZuEbThrUXh2vY/uR7eB2t1EpZ78DQ8QyxIuuAgptN8jBphnj8YqNtwjnd/dbS
mNP9S3d6UEaslYsRZSDhcevWunp12XW0B0KjMs3vnWeXwQ4isYRyZAyUcGst7CNrajG53N5PEPl4
bIiRfVf9pZaRZC3dUM/Pl/U21SCnCJLKt5Kc4//7ajh4Q0xXrJVpV1tC9ZMAl3PxSHphVD2KLt1S
OsbFYOABJIyBLl6w+12s9GMdmH/gIKb//TCV88V5yqFKAxf56aiWVvqvgDTdNDgOPQp1EOEUwfXq
9Vl3wqVV0ZvEniXXf3xiM0hXhxUwk7Dc3iLGZJ3GoSLK8faG2wP7kAz+RXnbP8sVq8cFsEvBlqgp
igDR9QjAvrOGZOB8Uu6Fo81AJdyWCdP5WxSaUZNsga9DbKX22mmKvUB+7RndXJIY0jbIYmXUXXSy
i+/5d7xkDZW4D/Fn7wzBMIYUXWzZdEihBERMHMA7uW5cCZb7yF28bHySlZSxjTw4Udp7XmShNZzg
1OS9tbwCu/pUOGzhDw6+LcN/Vo2BTNC1Yum673FZZh5nB/SXAQBCH0C2vb2hwLQXMfEXiN/tWyPy
j7Hg/U5U49s48fgqx5d/aGsPu5LuqJ33OZ3HoqFrkQ+hOg/pyVo+7WgQ9kOqrIOrBDGw3Ufk/Q7m
pQMZG9fhOqRoVJckBK8OfBJvzJBcCYZJ1x4Kg3jeONxWkX0RTy9v4otX12Ch2ceXYRpkmU0jYA09
ph6GvVhv7LhKM7bk6X6vOZb+OGlIWnMP3y51x830lBNJMpTY8tbagBqh2huxfQ5EWedsfXPCOnDr
IlsKbqc8XWVWZSQA8sFnReyoZqyOuyfyouK7C5bUqDkm/yVshCGOt84Q4qk2APVCdCHfEaR62+22
zAMwtOgeMV7CTeiiLkbhI2FRQYgFkpniKTRJwJtLCg54vKRhyAVd4ljFaGhjNlx5pTNbwYMdxD+l
A5lWWZhVai8cawd55skge42chQiI/zpdzsK3g2rsZQqFDlCmyYh1VLjJOzDTYASD7uemacx3r/A2
WfW80Wnhl4QX8eUH4hiFl2Z38ueSf2uIn1cqGmTGwqJPvz/ycNwBwkRYJv2VgBwYv/zj0KPxscuW
utCK7xKyNO5CS44/UFpmOUkh2H/zSklDcj2cWje/NmH2W9NNXFyde5hfngM1FQrEgHW8vVrEFOC5
Sm8cWnTLL6pQ4XsBtE8RckvqGG4uVD23Dd9zHXoymrvkwiJ6HGbFg/28pJJqXBeq+nVsoyhfTvX8
Hq9PhPldTTM+mrQgY9SFPaPKHWIpGZ+G91Z6TIB+1votVrpfJNWd+uaVwhGVxEFvq7o5IazakyEg
tvC2K3EoFkIVRY3psyy1wea6kgs7ZwT/5v7BJUMtJtuwe/wSfOUgmr0MdlHL5xTPiv1GVSzMTY9w
HkahE9C/s4bZVyb3P4Ml8KHlrUC+Krh3pmVGRFQTbD5hA6KpknU5KKZ2HmSYrhpVXjtshx7kml4e
20Fr6NeoEVwHclyaRA39Ryd5RiwCGwodQasSjoJR9KVGmTb8DpjJtuLqJjXrlrZYurEWE9zY/Dy1
h9H/nIm/tqT6Pv6hwBceTowHr969aeZnSoGtPHJx+dJ0oqUO5VRqC2s+/CQcweGDwawSdgmS4zHi
7z0amOqsd7BM6TTvVOkWi03aG7CooekK0LodOfA35winbOijhgUDr554pCmDumuxioMFWVp+1BO8
+YkMlhCn8WwWlhXqBRInwbzNmdJ6h/OLFCmOocV23gqxMBKhLvEwFAaBrzcyLsUvI3wpaaSewJwo
AHFN3XZmV566xSTk0Mo09dwttpy0k4W3mRWzsDQc9dD7AiVsHVcr0zcdUDiQQQTJ2kmdEwQskU7j
eUR6/B6RJJUr5VCHpMwnBOcQJIm9Yn82oW2OULio9zJJzxZr/GmVvwah5orfmauUgFul/Kt66fNi
VIZDjZVHiHpF7lqv40Y0GgczJFlOlaGQcYZk+dnrubi1qI/NnNMQhqEyzPje+AK+0hKP0Y1OqqVG
R/IK/NSiX+CZwMCoI7vSYKk+f3z3rY0mWxa/8gzw4d3zxNBeaTKlLjPjxhEDBrixSWeSYKoWcJmw
pch9YaALaK32h8Cn1rWTzapVRiK0Z3aKFydXAuyba3kkC2/ew6LlWuAw/P16b9UeQPYJ5j4+rpua
FII3HSEcrh5/DHjTHy1gosfPymUp5ElJjuzzx3ggT5M8beJ+7zW1ENS06I/vFLVUBqYcDkLA+sdc
9ZsOgVijZezqpnqKIIxTbdi6Yxz/I2z4IZkURraACsdkf9Fxha1JhMD1MgS/c/wLXbM7R594N5XT
4MymQvIzfdeyy/q0xmrxjY8CpUQSTtBSyiF5CqUK891DESp01F0iyt2x3PFzrEvByP5C56clML0M
wjBwX9K112/T0N7URA/yhbMXrTuKY9XxkzgdTRAWExR+AIpKuoetV+DhdTGCU+ynL3p92PZV5dB5
t+yPLYq3SkPrny7sTMyRv0He2zo+dIHp/thexd9XM0QVuPA2mOhuwmWaXBOvOiojVvK3geMrbmqB
vwPPBLG7Dt0nK8w41NHGAdI+jchAwOmUNOYgyJZzov7du7DMOn2ywAE7OYNMqhs+9q4WuABk5QdZ
y1sAiCcwZV3hG/syK7Vhmn4WLMXmllLBKZXdtqdrMtKVEzBDebS2Xll9+AVgHKODOmmr1OVz0Kut
DkQ7Wh3IXD2hk6LKznODWEgDwywvR1fXQfVajSKQM+JGY+EGq5n1AF1rzfGNakdZtdM3KRy1uX4D
HBGbEuT1mHzhUAdNsoUQoHmcmvGDCI7/AQdB3UFIAQWZ8glxiarFhzCiKBjrAVfbKrPJTEak8sgN
Uc0ZxpZJyT/dSZcDHBF/9WWqNvYYQ/SzWjy7wYCQXKzzHJyxJcCQ3nKMpB67lDwbg1TTTzk5yFpm
Ce1HFu5FVMdTYRjCP+WhK4zl7EcH2jU0yYNg4tpM/czEfTwdcIbinUz+kIBzKsxSG0rTWIjnzJ7g
l6HwKlHqWkbkJPgfUH6ItL2yIrXDSFhlPmENDayakWM1M7w8KvF8hNQQiuW8d/RzY/plFapmpVAf
4f+wokype4TTmaV6bmsi4+Hw9QgI1ZdBdLIttXfMrSCi6UbWO0TaAN9EoVfQoxl90w3KOe3TBKFU
S/AAESAFjsC0fl9m7Ns64LhRO3FSW3GVMnB3Xgc8q82cog/H8mK1BcYRcIAhh/dDlevrqQHEPLNU
vxN9TzY5B+zaZtfUGZznO7Ui5H9uQ/5x16RVSoIppphSPRch+aX9T7P3AKMjIw0B2sFe/mB1fR9F
r2+DnVvF3XO6ezyGshiYvjV2qaswgFzoG2kHqcfcK5smj5H2c1u4ysUcmFks71OGCpNUWGr8uAP6
tOzY8yB6IFwGHsNNSlDM0fJih9J3ounW+VBRDdNFnHD8YCZCSUa9LSjlgg3AH0woOohfXJjvQ3vC
HfBE1E7vUE3b6CWxad5N2xQaheDdvqDPxDyKE2xE7/hU3CFjms0lHiVYDicdntKPEIfpk8p7St7h
SWAeK4Ha1+gghrnd00OWLeVvHKne4DiRZ4OY4sqXe3S+vy+uzoyNYJdiD0GxIHpxnbyHAqQkxFcd
wAVyQ+ZiJBEAQcKcIJDGolVBvCVdFIG/DNpWGWi9FOnNP7xDkb1jX29aXLrv8I6V8SarWXVHPCXW
Ennj/rfmv2rP8hqWLG55PPbsdd16PTPlI5egjo0rbtfiwvBZXj+Z3ZcPH9/BLzVAA9KhVS6kC6ga
KSDFB7Tmtc6Xj00dwmq8K/h8JAB5hBKhQu2aTbBcpIyxth3fqnYZjM+7TuwM9qCCSIaqHyp4QLPx
oWM0hA7zsRfaEISuMHhnjw2GGxpsR/BmNisFuF4F5RhCAipOdSDkWzJ5bxVpDebcJXx+PcEeGw1I
2bg1FclE9QQg4BPFk7YFGJPYherbexj5CAWR/uKufOcjwMPVEVrK6ZK9xwmhYBMcstlpNACcecmI
ISsL24cOCxuUBByag+fqc3GQQ7gkfbesiNzvxfdVA9IewL1k1z0wUAaSt+4ht3x3TR0RX8XiDIWn
1NCnMoEwsEoK/tkTs3e5mrx2eJimkoHWHzPX5oIgm647wa8CWu1hK9p536DR3uHpf5sH0Is1oaVU
MMWRr1IZw8cWOHiybnU4NlJkcHYZEw3ZRti5QOEapNaaXui6MGszpXO9P6XTLuyouK2tD4nuhnB3
2kDu8sA//OXdvvf71I5ZjDBlvGFfcbkrObSb7jK9JGrZbVAGHgdoN9nmKj5DJHwJ7cPoEd1XheFM
3sULtKBy8ZpRKtvXKs6+lhMRwSBAAleA3NRlFR2NsSdRc6OUr88xok4RBu/yItSobjsaYK+B1RHO
E2nhOCoAcgaeNJqUipip0erlWC32wbAZnVKJ44vsdYBUgEHHcqDMJvREO00KLjQ+LCT1Bad2aIVy
V37Icn6jZTbuAwUEN7JHeQsf1gJVMseqDIYVS0K9ihxFQSqxtLuTNeWqBH7wMvYi8jd1+yzhskb1
iDdgCl33Nz5EqiOgIWspn7KxXY8x8kqeGm/GKqLA4/iV+OEUG3NOVA2HWITe6PDw7iWRndQ+Xrav
gomCFLFUG8V45+IU42/g1RfnVIJDMosg43z7E6iVL8PwPD0C7fz6Z6+zF3PBLhhlGto8lEGzttLX
wAUP/mnq1wzjD+V6APoDDnxLYa8HQlm1l/SQk1AmmQwGKy1ZfQNOxl5Jij9ToxZ4x9FI6PpOctnh
/RXHBynt+xAl17UYX7cQjpKlz65E2FUcN1wQR3D7GM0aeFFR8jaeTQysCuJ2e+SXseOGVtzupTPB
c9yvwOfIRmFBabjv6HFhJ8OW4VcQvHcqmTLn+JyXpH1Us+WaYFLKODOsqwaQtI48M5ONZOorzilu
STdw5j7sOegyKfHqxYKN9Opk+XU53RhYPrurAalQU/XGGYe2VYXW8OQgqojvcy/YvKNJti7izhZv
fuPGy0ZZRI/jWpLE++jK/McLGYQo3gOPWNrL81hoMb4efSpUmsRHlqY3ebyoj/0RRGruF0/qY/fI
lXUBdGyUpvCReu6+AIEU51d1auA+ML2ehe0qtXE6v9sME254yeNUQpHKI4FJrcedbkb0U5LNlzx4
SSrBRCpQv7g6YwyMmqCX/cXWTpiot6uuhJ+3OySHjKqxAT2tQ5VKl0hhO6wRqdI4lWeWIQ3fIxgT
BMWeNCfceK8xUH2LnFUidczRu0WfKw4XtsQX8moPlUC8RnPiCsefGpmf2XRNEEqL9DJFzgl2HW6t
oMokykhJZFT6PGE3taxdLhF1JUvVNW1uKB7Ri0Babb0uO+/H4h3eZ5a6HMHHRVj/nOluiPh7AVgr
LWG4IOdNsadkhREy16IwEKG8lo9LLeK2Cn7Avc3qyn6wHyf69Sl215aSk13a0kclcAT4EgIa2P46
wM0WNzmqkelH+1bXBoA5ItkHkuVqYNmoSIK5h5a0zD1I71GhJOkiE0TaiYhGqy/Yc0K1BqJR5xfN
5iHMMpPFwCSScut7rIfmhwKEl3/dzXUHNgL/n42sGbc34bRy1oCMBu+AASieQOxXESWGMKFADRxE
27YNU5My73vXEcgbIn20qbIDnHVUC1F0CHwuU1OKw72HM0y+NfgclVbAWiLveWxdamCGgMWR2o6i
I1P/LRh2ThrS1dWz7PUuRcYBlz27MUvE84CqroPDUeIHzvedgF+CwggL3DeLAj9Q5N2Q+SmiWUIL
o0NMBldpiDoSaMM/J9dGbM1GG39uEbUYpSmi98ohn10Fp/pZYFVBrCq6gmyZ2ICrm9GriF6/PUkA
Rx8aCwcd9SPdl4gu56C/wUEMxXxPFOAV7VSO54cHjm8+cIjc1m5/j8D4ZbKOVEC6xTtuHe0LQ2K7
wlPlTvsUfF5pC/O079I+VSOUx/M6m+kroN6fPOimlwYGJXVv5RKJF3/eJnX3JL3PyUP91eIKGbc0
emfnQs2QqAst0kssXfB+ZFMT0pke6iT5pxbHUMQn+fb+xpl846kVBuz9yoULImr4FWsnQKHooiz8
IcSlYw2Zuorkmu8TFWkDAWXTSSwRIdVS7mN7lDqq7C8D6ZPUj0zX80Qkl7vbWSa24WrKyhEDeeTR
tUkNS27vkpJBpEnL9kT5Pv/X6CxEGC2EouOHebw/P/GRskoPucOKUjFVHE7iReEvULC+e/H0Qd3R
8j/QQzLnexcR0nqmv7nJfY5Uxx+tzCSycpwTc0jiuOlnaqL9smdydCCl0zZ17/5od7RJuLmEm5Ti
1mDxmZzQ4A29QB5N6knI8mMC4Dq++gaavrwFmX8v2h+6w62Uti67355Ot4yUDMFm2j+9Fzep7yth
bFSKrAEFknzFQ5QVkiflLPR213Q4lj13aYwX5wnwqlzJHGyu/N0ksrf3ObxIAwojMJP+hapWqJiN
fcqbQ+JLRRFJdeQ5ppeLqn2ro6K4lrWVdj+pCD7CS8l77TlfomkKPQAD03xwMnmfhxBzANxwsr5y
QWovIpYi8GDPRRWy/307oEr8CzD5wjpv1SuLBL1vNx/jkIGXy/EfNWGUIgIcD8vmEjIOVGva3IG1
vu2QGPkbOOTk+PSBEgNmtERj7XHwwpmXOKmMCNqhXWSWJ7ZDDXChpvXpLoFFlOM2JBwjBIHy3XqS
eOuaiF5wBNKXThWhbdT5yvXHvy4sZc2SwDqRNDYfQ8FW6ixVOhSorBBAJxt/ozCq3M5+yrqMJ+Ti
aJs+EpbLcRGIFTHAb+BzKBPGmdGPiZWeEumWw7D1sJ6jJALAVfnK5JoWegpaFtTDu3lwWgZZM7lt
n9xqs92sieBF5BStuP4fbd9ZJAGNgw05witDaTHNEHXWifqjvTsWlrUWy7JvTXFRHGiYTtoXSqHj
CWzKTAux6ksUdr/oBlPi+i/DfXWpPKGwxkxeE+nr7GkMs+2P/uM2TZfNZ0zHA43l8Okz6JEELHKi
sw/fwdNAobzWefA3OmLx3o5ABAFC3oQ21sUQbLYph5K4RnOgspWXLbgZoQTlb6HkaQYPz5vgqhiM
WJ7hBVqHI1nEWDm8D9GRGnZnabZ/l5ABaLpl4NHV3shAFoElHnZcsNytgW6LwhUDdT+SQ2MrtB+e
WAYJcGf8Aaqg4Ud2ySvDA0pzkZqQhuKATbarD2SnhvZMe0FmiG7K+Qoa0+dM6clHx/vZYWErxmyc
sY8HUq5SdT34jtxBp7eV5Tw2gC54z3ur/IpeSvSoKR+Ns6dg8GHOo/yWppmkdz05gbhBjUHlEzPK
tOrDECk8DvFY6JvQjDd6NWAnjKh2JCubRG8buzAZ3bhx+BLzGEk9BpvcLFukHPFsMS1sin3GLHoE
lSpbaQb8h5xsnr7kuZSsYSHfqzzErT/ee3t+bOgC0U3REDPZ61+QZlzySyYlbXjsiWN41O0ZnYE9
d1DwxAxjp79av0ZfZJg0JVlUIW36lZSOS5+wA2EkLAfexace4zR4NweN7YgiFxyHLc4ydeDUO0d3
V+0jaCfBz/8uDGcCkrXk83xs6SAL8GhU44V0SjuD0LtyzjqNdcWukUrQHsf3jCD6XRnSvVMaGYlA
b0nlZNpB3o22+8UBH24tPHNEn/lAZO7ftznYAq5WOUxMv9bzrLNTsnX4viSUs2ErbYEYTjogFA5e
rDZo9sg2UnqTlPrGt/uY2Ud8lUdo8kEM5bd30Xl8nbeTaLbGZTP3eI40YbTp1TsqxQFElvZHUj8W
F/eZ3sZpKRD3pxvbNYl1GscZHNJCHr1guDBZQ74WJDk/MdoGfY7iU8H6fAryiGLbVsMyyIRZmTvS
aAoC5F+mwofcE2YcPfNtZQA5nCbLmbH8gpF/Eyi1D5qQ1uKl/Q2NYVdv+CsCixElG4IUADHh3tVx
RQtgdGkDS4NH7VSt6DkkRKuK6pfv3zZNTJd2MdN289oJlsEvCOZ2a27CbKb/btYYP+5LpbdRWAGb
SMf6LKAXPTgUtYFd6qx55BDitZnxe8+kgcy3ABOzCjOYkGMWqPA6NrxQTQ30GlA6Yc7Hv+DF0jKM
2Zfso5wCXlUP8ZuNzF0M0ncpEptMK1I8zRzbFEhyvQ/lOF3n3NQE5v5yEzTil33JMWT93GwbRCW3
hPPp/O3/uSbTa8+qeKSfDMELuW7UOfGTGGxRhRhVpYYGZfXqutJfwglRVKUWaXs5sJ8TP5jwJ0TQ
os/ExzY2jOmcT0FlolhQ/RpTImYmO870BcNE3+3ugCFVk6n8O7+yTPtf0gRg0aq28MDsp3V2P3eK
9RSYN/rhzOqjJXg6VesuPkAMSXXx2xe4Tciw9bJ6rwQACHI//9JQOAQJpziaUPOzaiaoJQ6uVqf+
dJbYfj2DkWu6JckhrFouzJla4iqQc0+570T36Qy9mFQ24+p2w68eY6tJ3MRG+zYhuqtHMYkW7bYK
iZ476hEtyt71BmmK/OU6nllgxoFiDAMH8lktWvfJjPQ+2NgHdr6FUNswknDbMGdr9kiYcTBN79wD
/BN0uOR/R4pDVDdZFPzvh6hfh/MnuLqT7n2SP+NDsE51KAIynOE4dr7ASC9d+ZWJv6eQ0x4miYc/
zBCG+P1+XjntJZ4kWjYj9kIZvWmIc3Gvdt9RvPTX2QFgT4z3FMnBEFGjMk7IGw7QgkF9bBDnI+xV
p0ekT1TeeNO90nM8eB6iGwkz4PkBZUpwL3yNZNgSlFJAz84+9ncdJVe4ARmiOYRraf5YuBXyVunW
yOCO97fK7vjc67Q8xHGxjZCe783HP/AuOLgDzWZMmb1o3qqEiqI56my8CcgnmT01blOitlrLwgu8
TMaInIlm6wOtmSvQEqXt9u41yTS/d+lRVhrZtzJhSn5as13ubqVBFAAN9ImffSNWFqJ9h4dWpXsY
CIr4ZYVCmK+U8F31JWUJjlaFLcLIwBo+fUUfhPmVCcj1kcS107A2B9IeFd0RWe3iHkDphSzM76jN
yJEq/CgtkUHDLKHMlsL1Iesh6VoF77zG+DC0zsoJ2c41JbhzOhGm9s4jWtV2PpXD0E1f2CXqJ74V
eYYlfJphjbU8otYKGE9niGr2vjD6ffcdi/vxLQ3aStSou6pBtToFhivyRtGxHnfMfO/nGzBWmRie
kXH+DP+2P4brz9pFdnw5BZsT1ExxeRvmkKDUzihs/JSh9MPJmFxl3RXSNE7LtKBkaqgc9OuAB9p8
0FAP5/Lc3ZAiG4UtNzH1CnahyTI7j3v/NqxG5EazrMcVwCB11ny+pCzWI5G2nQXsWWRB4N4noaWB
zvCcQBRpHOYat8KMwxa8HqCZriT3L5ggZHr5qY/yGtRUQr2jwVQM9GP8SHnvqNbyXpNvHqhmYmOz
z0F6Ef9Pg/2KZaO+k/GVN9KPGXOzzfZ0sPaDP+5crzNy2ctE0cut22WXMP0YNbTtl40DytyoDtrl
whKQnH6eJgUTtFv/wlhZW1lB41aEB2zxsapIujWqVHmaPb38CKN+ZsCLk17B1MzhVcR56cb2zR/u
4i92wqxWQ1XYV/4l4pqP0E2pN9MJ7NEOIPj+IJLjzyhXvTExSZYuVc0INkzeF63lbBrGOoAjBRBi
xY5lWBL7Fvu+v8/UVHqxMcleuGADeH0pVGZaT+oPkVUzg8+NQmViKIv00CR9BsjlseBbNuh4khtO
uwCpQNtNNpUPQX+e6/4BMWXvQ0DV55Tt1ZH1VDkWbxVBTRXxOHWy+1TS03mU8yrDE1wfH5HYIQoV
fN+sJFkyl5bEZKuK+wrLbDeUrEHzalKLZTFOH5IYJLtTsANCaPE7ns4GrLqqz3p9vsEqnoHTDJ/O
N1mlt3tkHEo6/DRHYBFnqTX8wJkQ/2jbthDuTebovJQLuFlU517zmoHRYYkxgue/bhTMfopx8enT
i6xpz0xB9ci/SI/yr/14+5v7Xr4xb2VYOGeT9kbh5Wb3e/0MAodzD6nMXa1AnOPv6V+rVguHSjET
Qg8GBw6BzRq4BYs8UGfBWk32UOTsuA6TQHm5nUzlxGxdwoDr+CWd9lW8wLjmVOyclLx1TMzRdxG1
U1X7abE705dhal/P6oXx81SssO1hFNWXS75BrajG4P3FkIddu8ccQ0GNR7jNBufm/G7B0poMO21l
27Ut8kgip6Kr178KkAiOesUcyAhlk6EGxtE/oWpChAO3rYwlXkod79EUWdeYaMaEKNvSFnlSx5Iv
wbWxvRKhzNzBui8PuNqt9D3A6PfvhBezwgufz63CnSWfu/Ji4dR0aTmE/FYIFI6gMqv94e9YPAPn
b5dkhrupSGO/xYXrb5wYcLpNUVKW88kvS+sseoY2C6LE9AXLUwfjZ7m5DN/bqKPvI2Kp0CBoQL7i
4e6iEPP4VHQYReHLLUIrx0XaqO8QBxYjlgCHGyzHCRjO6H4aEirInh6qgtucKgtAjHhdRku+idn7
lb5y1JPOELCA3OmoaYM9MGH4XgQMO2giLtFnPOjm/bEQQiy9kOQu4yktY69Qz7nWRijq6Gz6kan6
uEZIBPHIEjuQAuNdQwF3/f1BKTEnR1UYlyxeae3ZjgME864QKWp4rYel8CwI0fv+ycwA0hFgBSwL
+9zTPRs+ioKnu8/LbeyK8TpQ2AqfE7cLFe6L4PYFxn0KceJhDXFK/RBgeJ4udiajAU4LAMjIufKL
GE3bCg8JBw7syZ6fBy/gG5KUJ7opWbLLtNqQdZ+VA0w+ju10oJKkIVWdHcnt1VtcQHE21D4otq+y
r4P+fTal1QNiowm5/hCEsS6eY8kdjl4XJMvguyqyLJ7clldV145kHdtXSxd2un1U/HB9vriB8isC
KWFPUkxeFnwgshnH+Fr24ka0R/iTGqPYDaUsmvrRXnxd9lg/BkK6EmBcNxU8PfWJsONMEEcKeIcK
3uAlkgcDl9mbP+IJUWh4tZ13/AQLWjG/l6NBYoEFK1LOYymehZJ/zpEj/9s5bYZdwMg577ArJXkh
vOTenxl51RLvYntyNxQLEsKtSRWWU5H4mwk7giEiBbzW5pVNPBwXODpsWgg6s5FxmiGGyRhItP/z
JmxJO+Ycjo9qrL9QAB6AYM1DMPtFrdUiTj0KsumTOWatlg3DGmsDAn5o7lKNrQecD4Rp3YASGnv5
8vIkV9puk90K77SOmksmiriw38c3odyYP8PahT0NBHuSu5vP2kjGdJoqFVcTQvBgNYOX8fE+QyWQ
LK/B8CMe6/C5uG8/euIffZpiVzwtsBlBajP0ebjxIIbS0/XjdoHygf9BZPKxpfDnXVyUuUUvIfi3
3xXQBrPExCtHyxJ2urJNUdHELD+UHjZfnroeNz5jqcegP2vj9n8h52zceOQw5Iw/C4TmkI1GTjG7
VQFMWiPChlVqIGcivKStz1+5LWChSBFvFrfLEsYxWVMUwI6KsyXQebGvD3oLc8CAjKEv/v8zwUTa
piFh32i2resM/Bzl3NYlOLdvJ433UIhn4pASJ02BAKpkU25eX3OrAxO88BzGvnVCeeAf0LfSaPFX
Npi39fvWviH+lBphzFRCFb8ImdCk+9EKGhv0RJ0RlxEArlcHks6Z+epUHLWbLgff5huG1cwXD5SO
SWXRWbqpGYUxgOQZSsFsFDJqLoJR9/QujCHGwKBzekibMXah5j8w5cHmISdrpweU3cJJIxi0ds49
CSc8RWXriXs5bo7tYhmVM5A2o6qo0HcQUlv2o1kT8DdDDyY1VMz6A1xQkK32vP1LKOZY3WR9ipDj
SwzfBy9/KSDGDw/QV7Os0HZPXiXaCYkrI51XW+aB1Qf3gH0NbqdULsiCNIsoYELNvM7+1saJXwsS
Zj+gOLYpa35TI2EVuDSR5UyZbne1wNsgIGHvfet/DCxPi0oe02BRcFpmhPphCBCgEuGFKXczvtVP
UvEskfFeDO6QeKXQjPpV/iDDbcZagOZsKPCixKIy8nBmPi9SRTxg3CvnG2u/cWWXgdaf/YC+woW1
l3Hfs9ffxQltyay4/28XxPgJeVKRkzY+FEyTbstwk5zsDBpYGX0NETMZMa8M376qx6uTf3vFRLv6
gUW7bGCt2kvr+tqO7S/ph/kB6e4zdWSqtFXGEAvrTwPQlk8/3RqsoPUsEaNMnxGw0U5Y0Ip2mwvA
+/gokWjpmBzyMBu8raR34mNcv/sMCE71xxEhQFsxkEHNhjVNftR4zAqeN4lgT/Anr7MeGjtHJ7Fd
WDnZ1/tjTDRvGP6iC4pkf/tKBBcxJQ5aqf23Z/vHa2c900NAOOQd9nlXApLETsJ4yIRV1lSU9Ums
e0K6Kw242YqmkbFnoiIeHud7RBIdO86zSI96TBi7TYlQJ1EutSF9jw/itW6mGXOH23R0kDKCTo3i
wWqZViWYDY63zdlf8yjwuSZybjidPcD3KQlqHnmHuVNuLO+AasknObTtvAa9UKMn4ErMF350M27+
U01yu8vMjFEjrFNykt0BnRdT5U7oZH+IgffftOLO09eHFqsPz9cL0j1NuvZKd74XHKJCr6PSEGZH
Eb++Z07rn4+V+TH+t/mjNNvztrVrAjrFmvg1rPoWhWCqe/mO+kjCX1M820xCsQSgpYBtBh2DB5Bp
LcnA7jLtOy3rEZMnG25jWbJCxn9lXn/vB5/7pMmBTnSr8ppkvWcqadYcGJTZF5DSF9Lrl3lZhpDl
In1XByB3Ih+HlL1ZV0AED7/RlvtTZ7q131y4Mbg9ZXDPu6VrnELLIiKXbRoYVC4gL0FksKMyk6Tc
Rgf87Y0Czhi8djcpe3/+cjAQyOlvY+3SK0E/pjIbybKno6EpEaXSS7ZEjUKFSou7DFn4ylrDzkBM
6eGukDFvd4mCEs29ycKCDv8bGmsrRP9uzH81Qc3pO0sgn1ZmdodchbJUWkOeHtHF/BBz1cnfQzM+
bIOGE8wLIqPGzCRr1rm1K1gOhJT474c5I9Rs4gNddiiLrsHZfKzCKGH3C8Uo4OKQedBUlwFpktUV
Pqbt3K6QLFiBQdZQFwtrr8G2xMOP3CT/9gqPpA7xi7bvDeYygOsGH4VDgjcsx2Z+gcx6FVMmjgsX
zujjeEjiCnRhICPSim7DOK0bz6zt8rgP1EEQcl3bEm2pDJtjp4oxHdAUxVBy7l2/QHmPzCvKgonm
1Juix4lDXt0ZkbZAmnVpHkEyUVoUICU7WnPWO8PRu8r0IvY5XF2BZ3uoJwe7D8uYskAfvKySp8gE
7mnRp3x9OLe/KqvGLEgOuENaaU3Iunq9wqB9wfihl9mR6ztA2qxe0eVnEbjiW66hiDe/5Jr2U0Qo
HzaYAJUXfXTTSOG0fQ1QOqPweuaZK1n4ijducpdAwKUaD0avgp3Ls2MruNQUMia2CiKe8CFU7C3h
hKOiwuVXiJCUmsA+HbhbbaWYV5dcEBMLmeuRISWes0bg+fix35L4ZFsAvPYfZtTops3+JE1wrAsA
uMfJvHqjCLJzaKySrjcft5NOeAi6g21SARmtL7bF8eEFZ/+xSo2VlAhkvKXZ2OkZyy8NXKLXAaM6
DkbdUWoy2prif7WXb45dciBizb7UuwcIfsHecGQ77V03j06T5METgHdE8YsxxhBCQEW8Snb42TXH
6fQIebClk+ppEdiPA1XGu3vWT+cxWtSCvH6AGm0tN4Cx1Mnt/E9PogKebWWOe6YbqBbrKYPilT4G
YJBl3WHO6ndDbJQn4/PRqpBAqpr+fFT7tqhhtK0aiX/XUVn2asTs6Kj4vF/B/pTGnHxx1xfsmPAm
UYhm8z8rLjFu9cdOzWFypWFLxb1ejrP+3OEYhzFMNCXeo8Xp0Sq7poE+8BDOpUEo5YgkvK2kSgG3
5d+YIpQt1Eumq/zynnSztWH5/10UN/28fEf2nRiQGdxcLIsW1fiu8El58Llj3QdvewvKc+Ebbmht
0GiE9Ca1yDQezWUbcbT7we7gUpHb+v0fBQxZZp5ncokeFddc7UTV5HZ/wNNBzr0De82XKeO5napt
vLo2Mr2Eee3CQ9mEBdvS9smk1c3x4SOouIYbzP3qe42JY+LwUo6s3NbsyvmwAmIJA4mXt0jOXU08
yERWYV736UjJHJWxccFT5ip4tFcOK9n/WVfTp+1gOLy1XEsbZIu+ipEqgSA+RPVOSSzX58Nxn1Bu
19a3wihLepEVtm1I9lN0NJrHrGDXTwkXTIE/jSNKeWmnJJQda+3LBqR2dM7n1E2bqQB3XGRLTW4E
uR9b5h6MixdYWyGtJFY3iE0We5Ua1dAJCX0s6nOE6mBIYPoOXB7fTYa0Xh3QZHGxEgDpVC6Bchii
G9qUvwO0DZAPnckLqiD3oiZJGZ3ItnTfxupRqnlJUujJYu+eLkkcxLAqzRZ/dJcBGnF2o1bp2UaV
e5NqZrpFvQtzg8pMEkTSJU94BDt/HGGJaZ3Ih5xWnGSsJiGFvdyQeKsowaPepBvDvb3/H7DUZdcQ
4kLYU1RzvfIBAHiYAfz/y2QCtUElFRudHGg7xFDtcM57I4r8Dv+E1XB8LkKXgzhPh89DxjJG+42R
IWmOXyWOxqkejHSNYhE1nL8qIuvniM9mIMUZn8tFCljl8LOLduAB04+17QtDOTIKsqAxg+2q9Ims
STSDNThC5PnGTjsI0r6Saq/yQoN+QNY5I1TIgicYhqwbRJJqF1SX5Lp1vznJHJ5PfNxyAq9Eak+X
TS1DWgLjaQfGF/3tq8t4Oug+yBs+Z5u5PuDgALk+wNshE/vd2ezsQTNGgU41nGB0FBHb1UjZCVQz
rmYEPgw9uoQr733wz0ScRlBJLWxSf4BwpthW3N35U/+w2CgDmiQiI1jhY2jvrYGqyJ2osGppSjHD
ZW7SnbXJI/+eZtMsq0gEuhWtqziQEQK6iC9OezxspR0SX47JOqkozP/NwA2MBBNP+I6ukg7sLdE1
l/KmOOp67q6mKrlpSxL4az6DXjm8JKHg/B7uMQdgrvMAR3yxeknUJdUtyd+CQRdRg4jEqBgKpAdv
XVUyafCOglAIOMu+47rqjb8UOiahXVS9T5XWFSz6cTOj3OCGG7SAhVxXPao4ZcpJy9L4kp74LyPa
mh2824LmJd1yV563bwTEJi1t8i+AWeYCsgelV1+mQAsOmIKFiLhgOZWQ41iCetxVcSztRWjHRfWo
KvfsWMj2i6kYmbjqHFjWVrHPZVaRk2S5CrtxlH8Ves09YU1ctNYlKlUMnuinLEuDFZs8Nv+EpEuY
3FmvUvxdhepbjnvs069ooLZBjPeJ+oDG62QL2jmSpjLkZOvRKmsBGMFcl6HvEcUMF0cZYB8HztHD
OKG3kTF8oIbn0UWvlvulVu8ZATeddnriSdBPN4w16GhCZKsoRE1hBoc5PNBV+oQXsRlKoUHg2BNz
U9Qk6u0IIiA2fCmrGcCcgjKvGoIf0TNYrj/lCPE5BXlurPF03jF+oABQiHshDNdP8sCpx91d6yRm
0cVaXtw2RJ8GHo9Q+TNV4LpkTlC9OhghG9nDKellI5visJs1zUJy0I905PwrM91eCRzAhmUmSg/D
KFeEeTtU/4N/XHtv6gnH46WqC3bGozEeCMEqpw7AzytMk7pFymVdWQRWJOXYbOtyFBysXK4iolGM
4fQEvflAqoW9YBDD86d12hzYRtL9Pu839opr+a4LhLQsfEjOZ+1KFV/HaeC77nCNILXqdGvGNgEU
bA7MmDhV3gkXDxmoHnywU1f5HItPe2XgQdkpb/EV2oRLtIyLZhI1bEfUeZ4Ji8E7uGrY7gULLjFA
sv3GqqHH4Euqfd7vV+HhvWGEDLSc7mB0ErVayuUnJTLNy53/mFZXzXxAoriXbeu3UyRuX8SXgxN2
3jzj/dZzZD+WWowlevYWaK5R1IBmiT1zTNPVMVjHaOpV6eLIR8CuxRpX/z+2RR7UuS+aBQXxirTo
7s1j6W7TtWLb/YvNoNn/bWQyz+DjaD/jrHrWIh5sGd4DPj4IkO18i7XQd6FvIhkL24vcWeT3NZ2M
ZXC5/6RKvpk0pWS+GaaPcNvbKpLonCrzIUpn9LshM7+6CmUTmyyVdYpjFW8XnSW2BeqXyCDJUj7K
EyhRW/n8eMXzPE8LirVGIkry6ny/2/pQ+0Guu+6OnEZODnUQe9YiNRXFtYpt+C0Y8L6XkuEI9YDa
pxUbcdHTR5jB/nK76nU0ZmUniw/+x9F6Wu1CtZKjJmxRqt9LnXqPsfKiBlY1fVssizu2mXGR22kX
IPJ4LykfruFT6a22Fb8g5yBV3xkYzCbvEOUl1cxatazhMdqEjAHulxUXbPksyGxhXacmO8cueYOS
aA3JMLLzBak/Mc+Rq41GlxqMSRXbEnHZ1H9JXTR+t57ibLTCzXjhEg3pWny2k9rS6+iARnQUpnT9
qyEg3SihqkwpwPeI52ThCp9Z+epyCG+5oayQgOCa2ySLyUJvHBVQRRdDRvh+Hd3Hmjy+vpTYSlDC
zu0vCD5IRiayeq9ZqhgoTv4eKJDASQyyREUPRTwo+h6tV+yrSDlWkKtgcix6DMTVtH8y7YIuyhhO
2lBGlM+Emx+IFtHkOgrJk1EB24MGFi/ErUyNRHcA//T0MQsV2gydBIHtbLFMpDFpznELafCqzEyg
G9LtBFfF6slf5w1bA3CMopNn0rsxgELY2g5aNEXGxSwvummY59pXQG4SrfKVsf+vZ0xp7vHcTAN4
i9cOVi5mL51Y0oMDltTh3rJmwhsgZHNmoix2vgxDEYv41K07NlGimZ86PiRBrjQJy5lJ9KA84rIL
7GPhywort5AdSxE0ghTcvcLy3K5xquw2/U8r0DvMZABnUllfRxl4u7AFdvjyeP4vX2raDhkpwgxJ
21l9OPOv55Er8Xcc7/UrnYHakI1kChqC7UIq7GKH6HcmKDJVX5VyfRR1vrodbnBzHPFg1jQgE8EC
6ovRU3OqkO/o71Rt5Yc/V7ELGpHq8qvlLLD8K8rzGRN21th8LQYv6OMycerGPzZC7zl4apO7A1eu
oXCnYKPXypFboOF5PhIj97BQuYBKTa4MiikeuT5QQkaQwvgvVNForkNerwx12Sq0OHqpRErFOXt4
8kTQvJC3iz7MsN364HKkr/5ChGNxVbZJZoGBDI4+EbLx4QoBeCzjd8Elmv3w7weSy2IFxIAEeCDq
S1WcWvBxrB7diGm3efP80j4DZbgsU0xCMX1ejM7MeUZmvYkzZK+1zdFI3K03CZ/zYa71gXHr6FyC
4lMsE78zWjOQBNU4NJI2FlQTbo3SWSsMOsZKvO++noW2Xs3qTLNDRPOTn54FXeLfjs7nHAx9EAXd
VO0vN59rmKJlp1Fbp89VHCf/g1v2KuA3Aa8bul7ryrDvmcaIttu54qy/EV+FfyY21jWxiBegZC8M
vuPdh3vKoH5XdSgpY7YkwqbKrTpOANFwcN+XJAQ8rnOXzrqMyQHHJLt5eWwlNXRSmtAXKYKATR2O
rsMK7MNNdcDVvOg5+ocHWkMuNGKix9cSHm/KhN4kkSVLjbwCt976AfvmErTGl12DvWnFOBwZssym
aYyqHsq3Yrw8a5X0H1WBbnMyAQ8WN3odsQn+xIMH03dee01Fvk+1CUOv1d3acGtzd8v5W8zoByIC
9ZVGzazyjpF+ZlkhcE6CqdkXvzLHoE9iGuhisOGt2Zn2NZyTrMmJmHo93zghhLLjdGpyBo2grF2Y
onvuEGsQiFP4iuP05JEHxxOS10QwUVOS+9r9jAN+DctwESOo4kL+wTo0W60TkL7VccagKYcm7X4/
vvE3BJ9d8WRDdp+gMIZ/mf4CtoDEHADxU5jJjZyv6eiKQu5qLO5VbgoZdLnewMxQMEQlSFOk0b9X
FbbrmwH89f9cz4Xzc+bQfz7lf8wtNfXj1whssEPkHOp1JCj2VbstZjYtPqRkzsm8RpiAX11HE0Rt
CEmX8+p6FibQXk0/sA/K89nYJqISHINg6IZTq5kyle+gKmKhNc/joXnnnQKapdIBAN2yyd3h1jeH
0s+vWd4zbaeWUCa1onlJUKL0BsiKXf3OBSbcjBEowXMe23i0L5KRwnFi8Y/PRXTUbqiKccIbVKfS
cMTE36lLsOj8p2CQcvSDmiHlvIpea9JwB0aV4sArLLY2t/RiabQkydQ5L58uXRW0gEYNQlQIxkyK
AEe9JmwNhCPGXzXt6u/A113RoDrophDRseV+Ymbq9TL3kv4g5KUuB583dhCPHdZGtzZvgUeRJBHJ
zmMAtSCFSc7YCFd8JutHI7lODYUCBsyTMcblRcKIBCG8y1Fl8wvVbZQWWwDxr6NEp/8lE/2F1AA2
JxUPOlRnX6JLyc8ZKEUSh3o1/lT8t8jCKXiIulAPgYxyH8jFHk7pSIyOoRsWdOqjTWBbHDgg/+QT
+sivvp1lz9ABorg4QAUitcHHDyCOQJO4XPclrm3nvzMyGFINHJOeRGPVyvZCNRc6drMqCw9ugCcl
vVdBD78WcRv26TvClcDzsUMQbnV7isI19LxFTVkk/NE/0N/xBEQ5RmzuqHnAmmVhbDFG/t9Fn159
xrRgXJo4eOG2W6bFSeTGKOej4R3Ch8H3l7k7HE33XTWuPUFylui7Erh5bbJHFJhTiHiIEoiLVZIc
4Z47Wn/lm0pDV3MRm18Jl5pbX+IhzzfbqQLk7FnGy4nXqLcjJvzJ2vbZlxJNJL2CesZcdUbxIWy1
/d38xLrAamg/TcdsbpsvJxERBOCemDyLaBRW8eu443KVSJPPqdA2kHor81eQAyTg9jYBL2tDNU+2
Y1igEEh/x2lOKftV/szCQIuHCtNDJaZH0pbDUk6ky433HSFrz1LCZgGfiAgWZQhBHF+n7aathXhW
ghxmkr2/ahpVOllnraCcfzDiydyncgc1Xm8PTDPzxUKy8pjigOy7rvSJ8iXXgARO49OUAmEyBCui
9DGrKpZzhG7juv9M3IBGOPwTnMOs2bUn7NgT7IeWxr0PY7zp9qmbGHFFGuVnXUJDl+jDij46gkrV
/vK6L0e3KVbYmqmDRnkza4kG+hHZO2U52LWrk1fgIRpWTJYRaZ0oNLnHtLAu5yIG74fKMGDzwUnF
I+odH27XzI8/MjV3zyAj0IXgsr+tPXve+a3huo7tEaEHlWf5/2+fo7qS+O83z0xPBWNlV+tggR6x
hhGTVR73HYCC99Y5YgQ/lLbGCAJvY8+SLASAM8vlRkNMkP14zbwJdZv+gAW1BEJhMk1eiAZFWKIW
HUNyQ9fiLMFpAps0uI4dWKLo5vx0iPNDNisdtknWqyxH+jJuZoSez3vHYbcCnfEcWRPQznQJZDc+
bPvs9WRZprknnGnvsGOnTyu/C4AnmZxQT+eNngXnxoo0/kKOMSB/roonxZVZOoBrpu/j76sBPZ0M
7zSwFCG12yLlNTQiaEfqqMvhCPqoUzF9ziUhzUut19rW0DCvjgEFwKwhS0ZVEHzbla37K0qrS5hD
6PeHvvZ7EST6NtftTXBF4Nu0T2r46nJ543B9Sc22TrAwhhCDpvXK2wlmvGH8Ec1czY9ljMN4ebCK
x0clM7zBnlJjUHwvVwGkf1vMPpVLSNTalpzeutQuu8xapZrUHQwWYIkktyw/qy584OHHRYPVKcGm
zTe/b8K6uDdWGt2X+MskDOOk32itWtLgt9b29pcOhLfR0Q4htfJrLWa2fKsB9qH+mCez8XQDlscc
3M2iasKm1mjxQlKo+zDqzHdQ9HzIJO1bgskJuK1tAxol59+Q2MHREj9mv096B9JE1JOSVvaZdDPp
Ql1jirf/aUw0aFntzrb0CtTlFvqcpvqJUuazO/09Hm4LF8bLSrLsh+0TjSw5C7LLMxJwzDRmEclP
z+3U4v+EmLGfw+IaVl9svAhLDHeeBmtOuaqbzZXW4j5GBJ4WLaSsSNOrJ8cltwoEMQ/tqwGDt/uB
OmVFkAQrRvaeItGssnW+wJ8yakM/C+0oZqCztJuRqVa335gTIZDegltLYTHo5TE9arYObYYzbpm7
mF+DloP+2Y270aE+Vmo2fG4gFf7kDLCky1guJiIeYx1/ZC0sQxKw4CKZACQMjBgj3K6wMlNUBN9x
FLv7n8uVrrTkoo6C4UPlBkQtdRe44+Gb5yD9xXOkQ4D7OBYAkLQXvh6/WA1o3D+7pAZhumd8tB5E
WNlkJJzbvx9H3cB5JP9Ql10b7J7KUN30vK7hOmq+k260wSW4y5iBAxPSgK33xIPcruopBZ2h6VKX
UFZJAXiRdKSYyBl0Ecy2g+WR6WW4ZWdFsIg/4BDqmupNwlwvzu+cdHfcUbc/zyGCPt/DaO3/dvtR
8lU/f3DxNVrgNpwkUTKQBaxPJ97iwYn7OgSeoLDHqz8OHoMAs6119TfjiN08LJRQFOEFKeUYghYn
ngTLziFIBddjSX3VxO/iTvpS/rprLaeY86KLgadcAneCKg1hW/d4sx446lQ0/Db5Vfxsus7dC13G
O1u3edIF3DrtFr2dYr+ceebyEmA7IJzk9l1oB8TEgyu/0nVvtg5qaN7iqmeHQTULrFAPaOWb8AJ3
+TODN767Ej1Jwn8R4VbX9wY8rYv8sKUqYhp5fGoEMjCHjq1mLROD3ZFZ7PKyvMmWoeA5YmDpZhD8
FmpUllTpFppcQnxJVb30aSUy+PA4LRx2VM1GOdsh6a2ZOXDuXZdVnr2qJ3sriLhCc/v15OqWvz8h
XcMkQJcnqecgUK9DHgvsi2yOQACo5JtEp7hhzjP8MKH57VGwAyUf6e1mvVPXp5Zz6EV+yHb5w+Li
NLDf9rWQSPQGKlj7mnIg+LTQatrJ4X6MLRMy/gbeEXJXYeedies9FgEFnxE4BGe9wew5eg2yydk1
Rdq3aI4y7iTr//L9j8nUwcvmz8Gc2A7MlqLQNNiD9EDz1fPbL4xzMZo9te28nLwabE8FwuJH6pyj
wcYiYxx6cqB6I+hxJkUq3brhLOufDLOJ3RLN50LjS9ZBZYPDS8sWaafoxPF1sPPN/pW9uEI3phTB
J6xkHU5mh6X+GmatU6CANrbRJ47EtkvVj31tqinV2k1mXGrID0Je0dD4rA/qqr/EXdzcrWRcL3D0
+gGfF9UPqvIyJG7w2hnPzDmlTNXfE9pbGYMbbsSdlabATRLIctSLoqMNKE6I12LTWE3VDOYIvdCR
m64FUAbZJPx6Inp/XORj1CqOiS4qQksyhmLSaGiDd+AdzO+pRwaoNbpR/S30cmx9wUS3a44TA15O
i46dfuLsJdJLKgSYfOS7nkZ5GGh2U3TppjIgwtlScUBZmWOq4qGD3Yp8DuvnuN6EAWZtXpxdI3Fe
t9l1l6zKJXVHBb7WWO1NR4yAc8PaWh8H5ZJMx57TtsE9ejrzM6GvmFfVlnKTSx7K1z4OI3qrHzD8
USIO+ii9V8k8l0KGHTfTpzE4gVjh6IAHbY1c8XEmCc4Fa0+kFZNkEY5ed3F5G/En3lGyU9PMfYSn
fCYUDK92AyjhwIAATMZ14DsD3IpH79wjowEHz6BvJ787ge/V9cZsXHDEaIEITcxCC55BR2sHriKi
rgFraidv3pJLRoB65v0qfn+lu75lJVp2yZ8MaHXBuB3WnCS0zekmXczHPs9Lt3SSUSL/D0tBceWm
FSXApOdcmrJ00rD53OeQ8jnrT2HFmIfwyvLk3xQY2ijdQhqK+oT5ezFPaoRXHCCwyrTKRI8eE/Xo
WRLQqHWxPAkQkLBfeEINzyUCbKvOoXLkNRs5q6ZH4H+sEPE29Kl/iQhvtOLoiWP1u16GMiM3mDiH
OFFqVFT4TjNdqXYdmE7A+0y5yx7y3F4I1l6mDnoMixGj5OSw449qOxruqvRJSZIfBSMigiz3hi2o
rfABBp356o8cOZxGFdLdn8F8IZpJfNJRW/jbvfLB3Lj/1+fF38YW8eS4j6SD01LANmMNDJYhS+YH
N/ST0ErHFx+LhvESeR5IWWV3mbJyMVwKWmtdK9Q8hYsbetFj0tZs4y4tnYMmswVNwL/y30HZyUp1
D5uHFrhJgWouVGpUt6/uUtMLI77bPRBJSwwfCitJdD7ybBAKPc0tAMVGDeGv7/bHFIQuGmfk6pDv
U0uiBThjZ3taPTAC9dk/2sLDXF5FEG0LO8n3Gdw7vmwbwQpER6QSVuR6Xdlhu1X2m26ltfZzBvtW
eau2f/t7wSZlmPYzMGLhsl11vjY0XRkOrfrl6BGidezh9Xr55XC34Rnkk5cOG1JJCyDRxi1Y+6r+
bWvrhLx0Stp8tl+0bWYoh6cQXKAofRLwc7xZfCWcPWbeTtMEYZ91zYdzphzs56hmje2hL+6132yd
jXVsFvK2SLKXj4JeIqfkHqKolmCghJhmBcmnpEhBlYwyWDY+dzRpk3SY/n14Ajor6BBWjpGCxyry
UrdTlQuybPEeK5zFCs0vF0kM9zjZ3nUPBvyjnor7YQJYMxjB7NzLjOUy/bG4xdW3FvlUcGKxuTq9
OvUuopE8B/EmwFOHM48rnPhPJFxtCrRkv5ymI52iAnEWecOMA2K9b8l8pd83mZagZ5A9H0IfQV2N
nND+99rlXLL6SnupPYmnnYWd6yDibckQyRDZQGc/lfDEzQQ3nPHetiNPdF74uBh6ydx4Fr4ULvkt
lXa/2UpWdWKCkHyS/LM5t5FJriQjj2hqhneC2NfzRaC/ZsyOtH6nEtgg4/WISDgOvnGNNtz/l17P
s75YfTiw3pMt1xjtyuTBPQN2yEvXKdh48i4g1EFXEf3bCsSpgtVZiIwae59mwyrYmWQmzy3AXSy/
Nfw7sisIu/BWNLosu+Gi/k3eCF+2PH9BIOxa+H4yPvoRvZtp/gwP3nRJguw9bXQScrfO60wDRWtw
03swD5YB8HyHXMhRNeliEwGfc8eAWvUItbD1WbcFcJOezlUP9oxzuw6wkNqni3IHj/ISGPBmAKSg
iH3iIr2ZDW7ItiF2gn3TuKtc1Gzv7eFrkbG9vHOj92zpbbn77nTvq5MxQxHKz1BNlZXOP3bVVm1z
yWEiYJAclTJEIOE1xFRa8H1i5jWbc8tpw8kZd3H/OGoHYh6wLpmw15sxMDBYw1RoH0VV9yo8NPTZ
X2JnzfrFGf8JRGp6YtKFFDujygz1l3nOYv/LLMdNyXv8rxlXejWge90dIeMJh0Eq7r2YsYbd5puR
ap7abh+YETQPwkGlo6BkKhe61jeYiFI7Kr0HuvFUqfMytNoAOn7RQtLUK9fZQ2eZQRk0ZBt227yI
8Kbj/kVITI2Xn2tsRhHNea88F+HyCs0dIxM7zXqReFLDaXgiL8lLfPFCKKMjWof4xMPl9TO0eHSl
sTlrJYCPTR/n4yEzrMB7xppfBHmS/Hy0tvN4jU+zfXIit5oItjef6bPH2I7YXPZfhgRrpdIJgnIL
OWAEokU6NzcbZAzK3Dfl4qmnzF+THa0OOSZqPQ9rNTiECp2CgXvsHsQOcAQF5q6Dz/OfbhPAJe8S
9Hdm7YFubgvyMDK21gGkH/RGktJ7okIPuOz0XQu+uAjeEZ/PCIQgJM9oss2gAWRBDTdcwaftzh76
WlRW9Ngda9Lk3vn7OifEUC+VBDCgi5adUgpp1VOEXkc/ph/gdxYLWo5W8MmMhPNnQGbxVYc2qBAu
4pF1DF3Fw/klVbDOwtv+GggsGKXP0ub4pn1SMxXDZeSm9JZ9yAJMjzjRwLso0p+MX2zmdYWl06JX
Mp5C5qj2SZ2S3iXOZ6vLQcDvjjp2MXnJ1/BCCwL3AD2rwl6j94k7gFf94sg8csLo30BMt3p5TvkL
+f9bsjgT/9ZA+8s/GS9dOiMhpjz4nZrYEvCLitops7BHTyvbv3l1wUPZ3HkICsi2d98cIgK0zLxW
dfV9Yg11PnW9aBQ+wQWNdq8yRSnhqLVaNuTiMRQqwmW8E6Gp50wAV+s14FfASJ166Iq3IMioF3LF
EU9Sxkta4i0nvBC4p8tTeTYYsReMe6dILxVaDPihSSRB/GGGqHCFROt/4vp5BdEvEJVO55HEHSmw
0k84026672q4nXKGHZn3dk7hTX2lHHCiVxRd3EYwNC8av4P+79r2sqleiQHFRMyDvlSoYqlIFQ69
GNMdm+aWacaqjmIKoZCLWbHVTYqm3jdomMw3HJZcQcOTePY5jFo/VOQx+KwBbZj0rKLOCvqkE1Zi
Tpid6NJbmM0UL3BYjO/6AN26jn/RlS/9UDfnWlAlKfViKPulntESPrn+6belel4s7a2J7Bs9wGNQ
a3SF5uScWUtPgKJhTctm2FhlWbvlEPH+doW7MEUfToRc5rVfsBOqDxKPjsQ58rMU2Bc3Sv+sCise
UsmGz/uYeMold6j32/RpT9d4UU7KDpfvxGAleIAYToNah9C9p3+1mGEKa4erSoupyUiOvzyisfog
0T7pcOZr4Ve6JBMZ9co4uMZm7GWpqW61BiqMfBycoDpESiywi9s1q+eqGsOhY8YQH+9yypVDx+RQ
wf+SeCrJLTkrsz6+alCZa/olApPi2gJ/xv3QKVnBLNkXOT09oaNKBYf9ZqGqjtBNONzUchGrlNDv
+e72shPtZDWhurWaSmNhKdpCVme9WaOiGns1+58f0oqtbgElTyVzbROIG4URaMLcehf7n9wpYsRg
zOPkXJXOlB/+3zlPz7UtEBuWySUCW2lGpKj/Z6yP73SXQf7unHvj9ILURUvnc414Rxb8ZqWrL2ir
LUrGCzhRoRfGyaIj86KrLo5Tlxqw8z3sY3CHR4BGQvqK1vYg0FkHnX1yfMv4WwYiryOHpQ77yfqm
FXGTsIQg1pdAo+zSWRyeaA6arU2ypmt84fPXnLY9pSCPh/cqcqXjCfEBPZBdVpl/cuxt+l0TzgU6
akanMwubnAPykETmaX8LkaQyen0HGMlWymW7JEfyEblWFRHQ++Ly/a/T/i+013MOkZZFteb8ikyv
vxCLDdTCnX3/WOL7k+pom5THpEd5gzJxw6uE4aUK3A8h3ttPuxB2sPqjp0pLccfX75qEUyJ3D2ix
jociBKI5ZJ3l6Rskr7KiiHxsKl6VKcpal4UENqKKniDcYbADbxqzvAtysVhl1CsJMJjrvic8V60O
uYeI+ukADjsSZIMU6qR7lInyYL9sXA6W2A5NAOk+do2LPOE+WY5cJptnDwwfcGLaTb7e3fR65Q2l
AnAw6RZZqcTsjXlTQfoyCY8z2ODTlNfAqZirmjwRpW8sYcDMQyCieD4n/phFVfZ5/GC8kPnhKvAK
s/mqa5OhNzp1gFaxVWrDLoGi7K1v1DFfUr85IKdSyfsOuTr1TpAJ9nK27m4vrY/k43GVm2DbWXZo
8lRBLZW6oNQEwkZJWeoRQhGHo4fwtytFUwiwnDvewoLeDZgnwQDwfskbKR6V8daLPyklXW5Je/cc
HR7sNqEI89vBFiBbfmJ7pXAIfKQ9TlZFyBXkkelI/SQMnfisNYHbFx/K4YCNg2GOiPvdH1ZIoywg
8MZXl+lvEQKv/YQQSJZgkMieNPekJ+zYkdent38CAEZRdgosBrsLPXiQBQdk324v24keCErMicTh
Isq/jzyEnGjnW+rZCbaz+ALIr7ADghmSA0MKtfxTFEiAtb7nqILiLB0G7pyQ9VUqH/sOQa2HpCeP
mcGYEO8F5mOr3KBpgTHZMtZPxOUI+nABd5E7DenRpSgTpvNDeCx+Mczk+QPHlH9noltmQAN7Jp8/
K3MWkjRBNNkk5O6k84CnXu6Py19y9iTVGI5QLuzb4NF4guwoi8pO1VCV2XyUrhyhrjgEI0HQm/do
cG40atwVpN4mfnLHpZfE1b2SyYUWLk7SM4KobsLmZcjdA5Xxs/FP/NSA+jkCt8AcwSGZcEAyGmlY
Aq+qVYU0830K1nFkFA90sRkvlGEyTNbS1FTPYYlbRVlYlysUMBk8mHiBQN9c+gm2nI5U1xVqQ8NJ
272PyJE/mLuOsdhha5zZVa0EYRsnj+fJh/01QDzgfftRLjh/AloH+tOSElBKW4wDrdzrX7wcLZRq
gptdGLP3zeL+LliNdaJDF15GAtzFGcISg930dMzX8ZBvHTXXuqpqcnBv9PmdXotpwFsNhCrdnc2k
Eu+t+OBSOY2+2uuyFzMmuCsGutfyXroQ0ry2thuBQVLSXQMBhTJipQmx0JvyZPGAz5xPSV7g//9H
tVRQhbDfdloUbBn4dFW3M0gsPXWPncCr6e5ctvZh8ZZZx9s4dcAiby/VnqI6u+hUH1bCTHX1iRWo
/QNbsjcOS7MrzsWvCIw4IzFl/u6WBbQkPzcr3F6Rf6N+6YAUDzGUWczGUJvpDVqSONTHDovT94Q+
QaEbD6YjeqjIfHrjQeSjTqXWJEGA2cUGMZuXCbDmfYcMSkYE04buQnkEFcYy0U+LI8bMF4osQ/mk
NxiUCLFTCbye4R+g0TjCSy704Ysj5jZY44L629KhZQUTFnLPBT5sZOLk4nnmmN04tJ7ZeUb7XA6p
ZW9AmQcMuwyKTd3kQC0kFU0Ow/fLcT5+vH5yht1sAro2u9ozM2IvxVFz0/ofRrpwVX6ldqhqW55f
pm7xH0aBrEqqlKO2Rs2I6SkFJm109k2L7+V2Z81n8RXxMBC0EDhs4zXn+AehjFVmnC17s5EDq8JX
LvXHTjMX+tstzRVIQb5ealIkRaKN5N0+gSmuPoY//ZmiraLTMV8oBF4ibef1hE6XN0u4rNXr6694
uHyQusXbM7vDdiHZoEaQ12DxVAiBKTKKEAH6M1fWtlRAzfznSaXzKstolYPpRfM9238ZB7truJNd
61OabKkqE24+8gkn+lkyM2QvIR5OKZDNOAjO8RelM7clRx12kxf4uPGc+gehs75eD89q8p4KFUX3
k+9ETCOj17I04P7fJPUwR3sRROhlZccCmv1Ly9R1c10U/h1xYL8rS+O3xWcg+YxM1ozIyh1WtqzL
FLyAnGABT7ue6JrC8aCJZD/ZXiMdrNa0s+T0qkU3yU/erY+UXzZRA/BtMGoQtc+n5/6BYwKv2kxV
K+qLVqI3TIQNT53Wp/94MmLMwSciGdp/mGEwAPEyzz0dbeDjsyDIU1s2SMILLLPx4dpDz71kR9in
EqBKe8LX5kEmSyLbiSlUOiFpO05G9SZOWKalFJXgKaoxdgHVycItzd1h4zCUMhOy3/+naLY4rxBg
OiamgxtPo0bmQzj5CT/VKpuZVCaaET4mvnURkYoITO7A617P/yvNJ+ufH9ionCxnUQOsQzEHu8Np
LNelwCxESrbiCicUv4NwymX/K9HDQAIPFnKTKFqBSg8cmSdKTITr2UsHgSy4fv/8Z91UoyGa36y9
IADP6ZkmjtJzzOAILJ8R/pAPBF/Nj1KS6BN2y56cEI9p8l56o+rEchdDgJf4ydo9t7uzsip01yNj
VKJsCiqZFT1XkdTJurzw72EiEZAQLrK+hgvbXWEYtUn01DHJpxJGCVSetzzaOkCJLQZ0QpRj42+E
/Tobt4UwCckgUb4xECrgfKgtiRJq2StmrpOZKReJ3PaKOS96xmItdBN7zKKkAdiYl6MUUy46QAzS
D3i3WfB+yGXaTQoMm/TdSuEF/zf+dfiLFE6mBhOaZQv+/K1sRe4VcpZu7miYdbV5YTpVwy3eIDha
LKm8k/AY/GGQDL8atKoOlNuE4sKynFRvtok0Ln1+qGYhV5ZEvi2NRxxtMlTWPUorXz3pIVEsr9WT
sHSPsn3IXRnLRWN/EcbS2vfoPIRYp42NguKyLjlwV3KlKH5c1y1bMLctheF7fVy6e0UG+nNJS/fz
mCLoF10fVbD7tBdQWKOwFqQi5TrKHpqVaRSoTYVahqIpPnBmmc2G3A+7SXY/Z7VpSoqEDszfu1+q
nF93t6WX//WFV83k5iEJYfHrikMunwv9YpLVQMKDWcfuJYICqpJdZEm7VEOuIaTgRTQN6Z4ZHsEw
VzRmpjy5PniOrxj+lfhXKS44+dSkKBcqWjOnblYULVRxuO52eOQezGOWyaXYU4ymo//rJm1/VQrN
X9QXZvZ6Lq5hcjImCCDmJiAaRa3BiGtFrDtdzN5vInz2vsR36u69drtmXapDGLuK9s3MFHUudBVu
KO/Zz7XCI7/3KWUKmo/TbOUhYdE7U9k3AiWR8Dz2kQjgEExQ/+2Yu4tkcvkm/2ov558Ja1VNfzqy
REcRMfLsaWybcC6MN3L4U6GvfbTjFjQ1YAteSe406DNkECSE0IWJuFHo7UrV09b4PEhyIBLV2IBM
MNPpy6s8Pe4dFtnOzhqiiuh38yYWs+nOFKOeWGUcuxqdCcW1zlueJcU8HXL9taGE61PNMzO/AdjT
n8fmkrZtt+AikG0GWRuYSa7IAbbXHw00klUeNNJvxlHGrWWlPoWrKtXo1QggNLV3LTKe9Cd92LGd
T3zOfKwlQefA6g4Er121zOinP8bYvhyfiIC+FvrHfyZag8nqz7FGgHX5R40AjfaGXKAYPqkQBVBL
UwpeYe1FIbRiHAXAMYX2c/OKJBd9AnhAP2tahfYLy+xto+g3Y7VGjno1CjCzfsLoYkkUHNEX47j2
wV7eL9naQ8O+kbDt24Ciu+nKlUDRxwlwuw5vd15lEmv1ZHO1zOWy0mUPhowdwDMRfK84MXocOjXB
bKtTSmzVIOsTr4N4GCtyWvhLwIndmznxdyrqSKviQ7pId8Elpn1QI5OjHtqfFwTVK5Xcfr3K254X
OVvWbJfSFxW7tbfr8vGbTijOaSb5fM1NCMHAApG2adByFt1d00Cz+1P2AI/G2X3LRkHMzK7qerv0
Mc0fT5dBLXNubV5pVZPa3Ltq143IU7ztvExEm9ryxUtHMExQjiyXOLqBxJrEO0OYR/N0fKQyFK4Z
S8JQCWot6UyeDMswceBTmTh6PWTl+c8XajEE8mPE2+LjlLa28BKPdSlhByZWbzS0kndCrqZiK6vq
X3mUtDCRPjeo2rV6QLxDY3m79GLf/NMw8alVC0sSu8UkR5NHEGBFnXF2lsklLVvCROmQAl89fchW
5K/r3SsVRLthVF2RQutSa2EX7fOuSMr4MD6NG0vAMHNuuKMCMRqoBuV9VJgZZS7sY0AHDBVOmr3R
RLB/Mu6L8p7UfHQ0d8l8AnU29d2nscLDNCNq6ov/EDpAIpp8RUUEQ35qjJ5iCY9GWRWgyCUqChE0
R9ew9SGlQ30WjQ5hfyudKylb1wRHIjUyg2bct2l9aUoZJzWsmmhSQJN5GnTchq/S0Rfjke579yfa
EmRfcf7m/rNCpCeRteVYYZhDwPmjVrqTkNdTioVcA3lpjTBYqScApshhKHIrZR4K+OWSPUB/3ajD
9uxhnxDAqORb0ltCZJbWDV4D0EkQil6pLtOrcBB60UB2FQKawYAzuW2jXrBFQjz/mEetZRJtZ6HI
VGM/P93IOJkIVrpeFgMcctWAuLlQAXn4QTutMgQr1dZ0VKKPkhmKWV2HPlXPzQ/0o0A9kkqrmi/m
XrBsCIBYfWUS0yIdPvH7fWLuBlZoHxO6eGhQka7DnlnZukEm7m9+cF98/UsTMOEXl9K2Zq7V0rNg
3t6gyrQ0JRhZta91Fcs+0D8ISGy201wOgNPvDAAunkYhlSlp6q4VnlM8l0XhHYW31etgD70yDQEm
ttA/qPnIzT5Y4XkLoYu3433ZyWmSH9cGR+H/K7PvyTevPLZSMOI/+UBScbKwyioGmSthTfBs1yB+
uYuVZ3yJkmZA15LyV/SMVDZFUguPVDi9Zt7nVc4T4TPSGEkVIo9D9tQsuE6xuIp2H90gYJltmOje
lwGGigrGd+Twa8OslUSfTs4SYWPgW93Y5IUlvfpYIF8HXSenF3P/awwDzPf4OhlPDmnuq9QvNRqW
VcJpyHJkWGxnbEdjedIT/cTqxgRxAumfkwCnadmgT7i1u/R2NS1KfsMRoOsQwLzy8h01Ln5qPVjK
vYoQfnM/MJ2E3RoSKVYd4iWqXIaZjSk+fBpWsBEssKB2Aeb63BvrExBUd1IWuAdqpkRcASGcaIpT
50AUq2iKVaW9dq8DmXGCHUoW93JHSIN6nwsM80BfFIGTg1DyrUL/VZiuE0lGVn0s9nLGfAFClkxQ
M1IvnxYToGje+jeB56wZeYHcr84Z6crM5Z7zRztsmFSWMGvD1U/VYX+g1oLMdhwC2ve5S0Ubvp+P
2ovvhe8eOVSyM0OYukt7W6Hb1igV4VV1xyX9AnfaRhEcV1wlczKyCuRWRBLhYZjGs/nQ866EwVPE
ns+eznzx4ixehSn5Cdoyp7b3J8aRvNoD5m9pFmI3h1VpnKroxlx0jTn4RcZLvophpOmA3S0xZTHQ
4w92jyiOLqbjg8EfSChFULnB4qD5a8iIMY9qCM/aox6Fdb43l1ci1OtuAum/XTvZ4v25CzxvTzl8
pi3KCdyOo4q08NnZkjsqXXhAY6SHmvAcSlZx02Oyw2Vq4A7hlwVWrNDkUjFdowFPZhuId7/43eNq
SmjJTi4UsDQCBDvnrUR3hssjzXsuQKjLQ6CYitysrxW+0onhb/h+rW9mwOHwloK6uT8fcTwwJ/9O
lwBLExwEF/tD9/YBLQTYom1wvO+HebnewP/RaFFnEHGjOUmvkz7yC72coCDgMtm4MY/l5iIoEq1c
HbCSec/Jk6rpPdvlb1OvSXWHGLzvsA6P+ninzsXIOlJ9i0tzb4+ntcHQ3zThEArLoDI3QJRXcdPN
AeM7L4xKSTeufAPKgZ4hBgHZXjhUo7kCMeYYY/ALhkapzpAZkT2TVEDDpsaILPsJnu+O+JE7Wioo
s4/4gcfs2Glhn7keCE8PN7izXWjHYEm++F4d984Vu7/VoLq/fe5hRLB+4HPLsSnJaW9bafI6ma0m
3yA8vxPG9YK7g9jJuzRqaX8ucAgox9UzInJGdK7IlNauB2u3Tc+lQDgutV7xGkb7juzo03wDUT9l
dvoF9ZcyFv9BVf2aA6oTZIoAjvJe7wA0oC4UkBULrEAG/rm2MTmmLXWy6rI9QxAV2AGF7nKueIjt
LS0gP9Jo4GYQsS3ws199mkt3n8nHLWGmExg5KCFEE7wVLNOHnjNCIB4GVm/522LjTOtpqcQt7o0T
tN3NswXP7vXkzeFH2HLFXVnocyKr/MvCtzagxISsMcmygNenzO01eCV5XZ2v9TCBs1HdJ/hJQbqJ
KOPAJNlXrTqZ3LrYZ6lEP82GqPg0zCQ3Jm+a0J/ceGReuq9zu+rqj4A8ARwazFbTEEpMtfNKggEr
j+K/mOIX+TSRItEoLCcFU0SVudK2ZhwEOUg18hi2Dv/jeNGjuofBdiCXVmTjPfTU4yk3CQt89rlP
LcPA7BkvQofenoO7LwKbUls/E5eb30TWSfbfvlQ0Kp+epl9CknynbHas65RcldkLtSXNG+VgQqqU
x/2WL38SiQ+XLtFHRPeXgZIguhxJPDwAAIzaPXUyRZDCPu2lykB07/7o1ZtZe9I6uA43JruPZVRS
LfbNrA47BE7pkgjNQNni5lXsAGyvGQcEiUr4cMZjunF+h5ksUGJb9Zd7CNzyQHbaPoIZgn+/ej0c
1k6vlOwbI0p9SsOyUCqxPkKrbNdcgBRM3aJcxN4L0bTWTImdzbAnMDDc2VabomTlECTvyhdPlnKK
kojqBVaBM0oMAs+tus8YnQlab5t0BEtGnYiWJSHHDNoAHhFzmtgmm1uJFwFq8Cj2K2urAZ5lAvYj
ErIijy6zZZFxs6DZ0SwFhBai3agGM0LiNUfP3MKhPbbaHemsK8IFpf2QoaXsoCUAP5/XlW/bfZf9
02r4c472oCnATAYlXepMoWCGqMJ7sQZJcgvz/NXFYmvmbJbmTdaIf9f8EhEKP3NVAbXdf2jb1FrC
xtEqdBRnRIUty24QF4NUZESzt5KOgvEOfX+x2VCjzsih8xpd/Vn7MloEc/1WDNGJP4RHmA6Edbc1
Q5eW2BM2NpmO9JOBTWTPa1zUdFbunX0A1hXfWT0dT/cgy4AOhLv+QKcJv/i57dcJkCkJXHy7ol0S
/HJEzoSWkYqhMk8QqnAnfB3OLxn/BUj2EXHZSHrdE8ZZ5jPs79n93XYyy4UIEebZbFfdE47fS1i9
tixrRRZPYNd+gLw85lEtlPNI/4G8pIcaLYi7e5Yfn61aCgyjDAvyW7HT5EZxoJhcR2kX8pOVp37o
h8Qy69hhgbvBobwK/Rz1ZlBS1cqbjlscAeyXkUA2Pvd69iYgqiMtR7oTViZutMKt6YjfJHCq99F6
9izv+fNqsRznJ1uZCuJZrQOR82FZVPK2NtBxQLPB1iVX6J3qg5QdulqrDwglXVJbL48S1D5virh5
xd7R7zlDP0Jp8gjohBzw8D3t7HOllyvp7kWQgqHtFVFORmmQWD7gV7ix+Y/T26GTahbPLY6k2gCe
iNCuuQsblD6JCYTJOxfE+XYkM8egLPhjXns8OMBeP/LsSdJnm2ZFeSdn2axZZDRBMAk1bbHly4bW
QpDJwyItMLNOFP2jXbb69MaCwlS6vvdLVNe47OUNC/llSQc+vpasanbmO9Q9LkFQoVQkc58XWuP4
uXICyrBGOq1QPS0HWocvz4owbZUS/e2HKTL6j8ODH0QEFcIlOjQ5zutMCsJgwRiSjaQP85rOk8Cc
Hs65BWsIIAMrN594LGo7FVnrvqXxFY0o5foSzN0WEl4+GfABRu82zkB3mgCLc7IWJB+sSiC2R881
U6ct1cE8LyZ5zbIBCOz83s8eWuwnI1gvua4hPqwflArvuqyFLemFLxGVyeAdTxivuVjHMax7kkk3
nUcOVq6WaQxUNAJhVemlMoCRNuQoI9yf+Ns+w7dYoNbJjZnUPL7O0ihvaQYTj2VYbjpMT6ltkzE+
ZTvDdHjJy3WgaRG/50d7ko/6ESbSQNjBJ8019kzBHjKjPoeNxi5txUPnXLw724N21XOtJcIA79tr
0tqzcNsdF7ljPOllxRQrypsRQvTppkIgOEHwjAHmXKuMxc95y1lii91bUBpVpFb9+nfwD9+/5zEi
obAJ0hAcDLYwoRECBQg4vFKj0HkSVNVjj/tgfQvSEC8HLBpCIlYIm0YnCqC6lTkc9DBgyKHL77eW
z+1EIKcfX0VHL2jHSUpyB1UFiJeCmq0UXwI+8yiX+kWT1cXb4HvbU5DMiCWr2FPz06t7agUg0b+y
pFUAd7qorREwq5sfEF2xZpplFhNt3i85qsmV6NeR2w+0SpRanC8FSpSHcwBJXlOEjix4C7hVJTSe
PPTVzdH0hDCflRNf2UZfL6U7gchiTmjJEvasxYUGhHO71igtpW8SmryNFeQVXOfvpg4PHLa9GPHL
WAGkCfx6TOFr9xn8pVLMoseL/EIwyaUsa282KW5NjqotpS1SbL4R6g8VuqYJrMFM+syw2uNPvaBH
LK7jDaMSj9aXy2r+6b44btX1lo62md422pFSl/TyviQp54NLBPM2c3eKYkfaUaxeP7Ke4Hs67LmT
eGA7PVOF6ilTCpriVBfoH2bXOtNfk2ZV9gBhcTaDZuLjW1MMwIhTnz6TG5teaLQd589yKmlZc0g2
2fvE2i8YmnfWpxCcT4jabu9apoLHiC3vqgNGgiPanFGRqoo3boXAdMMdqwO3ElWXwN67CWfycytl
dblTW7LlkzNm6gax1Ovo2aOYwr9xI+JBgMZZna3JiDQYHuHAvjlmAhEOquY2j4uud/tzqQcLy5h2
ehfXWemOhRWHmfQK7OBSpzZr/XpcIzpQcJMG86l0GczYHnvJc59XG9KUYyMcI1Le1nvO5UDLlgCl
w8bxZj+yqJDcRTF/66ZJ7jH/si2OSOOwdypL4mj5DV/KKQMQRk3rkt0w1irL9CELVrf9q7uwrVJ/
4YqYyvGHfU7ClqPRNwJBSGTVgRhFkKGWVogJzQN37weKEHZMY7nWzVBjH2Fp6Ubo7kxQDJDVH/id
TNObWZzMIe98WYWrvltT6FN4oFqucqX35SL+JWw2rALqf8d2Dag5Vebg7ybIq5AVFfA47qWVUY76
gzYfm+kxgKjNe2hBlauukG09e4NwObtUQFhj53iLPNcdEjsdJpiP5b6rfijLgKjv2ErzmZHBsxPH
+l5A83lfPKBFrg4S5Q1gSxePTGn8yxhBnPpeTIVzzjvaN8gU9iC22Muj7KsOLJ7JW2o1JM/b69u2
5MsG09TFv7no237wECiflnzQvUa3Y6NNHkw+kzXm5LBXspKbYCDdJbhlScgtdQ4IuvDR3GnposKQ
s6roztNGZ0ZSNPm1J5o+0zxUMzy72ZGlch/YjPC2mwBtw0RO2FBX+YdNOkOQD0jyjt0tFzdRfREs
3yJKzt+E3ObezJo/aEgx0PdfI5rkJdMhjSjOCFdSu0s0BWs8HPStJmTWYvk5H45Xv5TNEALCsBZO
ZgLoLgUZdjOtYnI3LZkR2nERR6Q0mVGg1nvOP3GKNM1mxy3L0TexNbmyETEy1ClBYay82IQ3/pPG
atGyYLslK0TCV/qiNpKbeJFTL8Qx8cL3YB71EkTwfR49GwNQSxt/HTw2QsszAbi33KYgQgyV5alC
YD3F6z4L1JxHvPS1TV5v8eAVenlf/hIN3eV3Axln0XQSA3goOeegwwqaF4EpNlxc2kc4+dTUP32X
dPlmw3kZ6WZYt/lq0cJQHsKyS4m83DHYuvIJk2DhxZ5D2Emp4vc5Gb8Cn34H6HnCo4ZDHY8mH0QJ
JHhiDJsHURbWIjm7NGCfq0sMcIZdR7wIz2WMN3+M3NTxxu2kvY5bAlLZNDCwAlKKDJSko6I66yZb
zRKAO+X9VzcW9axHJRwzg8N2gkJKw/OQpyEZLQ5j08MFTws+hX/wWOInugIOak1UI5jUA1jip1xR
oWUb4c5ALExIq3IxqHrz30TnTuQxlFqlnLY38OvE605WWEeiPkEw5lnUIUrvzlN1E76+R/DGv2Xp
k5+wCCC4ByP9XM43/Tp47PuR+m0mJ6M6FD6zTENZ7tKg4ln308aiUrEUAGCQk9ZvNtm1VMbmMWwz
3R929zVljzzqmLLJqlyyNCxxo8l019XOZIm2/UQ3Dcuoj5YsMYBlQ1YPFZK8HgXVca81veJ6TOQb
tKmOH9DwaW1431VM3KO7hiz9022brQ+LmO6Y7HG7uYbCE570EyzEXhjUNPeCOQ55GS+MAr7pkEU1
+zrR8ZwzfBhhTY61hFGAKheGA+lSPw7o7VGXx1fPR6LHnj5VL61jSsmnhRcM+V78aTKuPgJWqxT1
EoFeYRFvBxeW+ApU8Y8OclcrtSMvNSPngZnfA4vN4p2CGlP2OxaGWtIFD0fwlO4nnsF+Orjmxqa3
oi3jZFdYGjkdA6SVQSATQlXcVfLwLR0ZPCOc4ifdxTaV6lh1kdprDqwEjA1tdqwoQ6nIGw4e0giv
iL6HRm4EpcWck1H0kbzEQfoeotElUz661M8CGXUpAwvpXpVKLBPQgMORKFAdiBSiu3LlMpv3op0g
m8gzFvfxssKiIAkS/bf/8A0ztz1u3+ewHscv6VRhnLakJXXjZpen9eGBBmX4kje5LQSOnoFd5Ev3
GdA3EECG2NwIZhC943ZGdu5sDb7ugyOeGmzkNjGfln7J6+xSXws7zCGEbmVNZhMW8LtdvYsIxf/d
8hhKBs3EdZcciUF4hY6CnPAvReay7zVMucj0C7jE7O0F053XmKrSfrO73Dh5UE2TWbuWjD/e6F54
UpZ6/um2upjG3FGXQHdTCDVioGoI+obBzNF1TnaY6ZJokm3RGiPhCS0DrmuOI16/ktpJLUxAxBSX
wosZIwLOnmrblbOi/oEbBj8zHqDOdBcDaiB0rfnP3W7KdDkXVlbhSoXdB4/Me5xQSfjNfUnr2bWs
GNM4JSi5ivXL53XML03BzGggYjX2DwXKBEcL7Wcs0qth3hyLGRApqMV+MRbzWPIFettlizL8yrhS
jVfGVUvwt7D6zhlFpSkOkmjHWE77ASsko64ZMDNdWw+zekdtbRmnjNtuXWlV07axNHalcWWv865c
Yg4rbqs2E/4n9JzwWljj0R1gx/HN0WQKFZFUbl3SH37ckSYDXWBuMWsmOSLM2DC1LtiyW6rDwblX
Phx7xS6b+ptOaRaqVMg9M4B7AZzkQgNXGHD9uyrb0VAPppT/cs88JL5oOo7FpqqDLmtGyZ9PglUc
CzEcXbW9mT7gbikdwR9Z8aele1U5G7dE9KFXXzTeaytU3jBEe4RAKVJXwW4DPR9WsLlIuWxiKtlD
nU2Y7gGmN8Dar1CMrPV4mw1DSeYR2V5JVnctxmAWHNY8yJSYt15z+JuCnJzSq3w4vBXWAi3uRRKD
vxwUk0iy1TETG+lBGiChU1ysswQcZ4KMOd6ThDFkFiUvM6sp1ov8/o3Q/QmnvTBL0gqRGeofZAQh
rbqYjCamp9HsaKQD2f/Fx4NaTbngIQfmQGv0PuhsM8Dn6tAjOrzFHY/93tSF55YkfjJV0dKfMTX5
MECoksLS/6O4qdGwTaQd+e2HTOfW7+7W7fZEWASOCgvtr/dPV5F832G9Esp2ygmTeqL4W/U/zmnF
iUSQK4ugVD+0azxRh3lAA8VCYbeYqzkuEuitk93+owZtO6zVM1jKcfTMoy5eH/NpGpI9ubwVsVZh
QFUb9Q44J9llqnYlAi/dqzUoFoLwknQLWjlwZ67kyOABgrecSTqu9nTlSC7Nse8TIdW0yWg3HsYl
KKdE2hl4VZtEMVxRz+3gv9Mm+5PI/BZZVcFMlSvibxcaq/KCkCjg+LR22KsDOdg86hVZ/9kX++bu
UO427R4V0S/TwUJgVLML0qLDsDfLBzke3sMr2jNkBIiNisa0reDBt1RoJlzu+30SQ5ObeJFoLcoz
dfirSKU76G5IBp2WXvNHCxegx58yFirvIj91krYEB6B4KBWv0gts2YdrnW3eIvB/lYlDhsFKu57f
MvxlJgNgfdmQ9YGrcIv6VQgAd0nQXAgmBpKytjyQVCnIDGQKkttpKU+Lvka3nSLFkC7CFtFDENlI
0htY6HBOO22mbjm/od1Mu7mqbEXe8C3uI5l1v/lnh4ldEJ/SoUsOSRpEX2uBYm2p0RGB1S3zjtw0
VYTfiHE78WB6/yPLKYHfIgTaN8i8nFQu1NhfttPeG4eXRgbnX//Q9d6uDn64WMqhq8Bz6KT2L4/6
TUeiLCAj042F730JjdJyRr7Fyw/ouBq1JLyeDquIyRDJZZLFGTrBuMmXooHk1pFgnPD29x1Ukm/g
Ee9gK3pS6lYA9Qn6MTdRYmAGVoY1IITUQCwsGG35hc8bIruS0/Xkd1VElgzCZBgJmyzGjvDS07Z/
M7Bh1xWKNZ/h2Ay1Le0pLZPjUYMvL3b7YWJLCft66nQjxnE2cVb4vvTR/ELgG+5RWSsv2hjl9oJ0
H6FGZ2csn7LMxQ3QLp8jt4tJaqrSEOy+VfX00rNQJj5L1E3AtUt7bq0TucfJmB0ONv046t07iyfO
7gsRTSvuNykOdF5Aozl+K/Xt2dK8NrILFxHzdVz9O8add3uIS1XYxoVbajOIKjXwXUBgPeGHATEP
ebPF/i0m09Gi9krmxhK3t4QX5dxaZz8PS+ssFXvhb5nQvkC1QGS9DEJZaLTQFeuBXVY8zPf1anB4
lECFN87tMjXo4cSvfbNewpr2rlsHpO6EQh9l5MuY2Q8UGMcl9VNerjtCgLeekmNrnIUcBVJ5Sj5x
SEO5rklD91KFRNA6231n0dcMUuQsqNIjg4xJX5dNq6fUreXdymlI5cw2W8i0J9PFiaBiDqNCs1VR
/pFifDoM/KI5nG+kcJiTVu38MlbkUHyhYosCyEg2eJA9oBESNKOiMrqblCR8ixMoMHxCkBcwof4P
/JQCl1Lt6Kia/yqq4imvTH6qr75Ax5HFVMKawHQPcIoWSc+s1saJFTwJee9ZpauMD+AY29GkMyIE
1Si6ckWctMsSp6H8cwF9GhVdjTB2kaS/ulUXp1QztAKW2GKAl/AnAJPbuz6pYc7N7OU7gVyDKlOj
tEFQB83Z/INt4Wo5uuB0OZvXw0mm/9WZa/J2nUpGAs86Bggru5AcT7nFd4fyJIu3r+/KirK+qNe+
LylPlMGM7RzAZY9lT4CxRdcnPtqzhO97rwA63EPOQdIpLzVY60wXGRQRwYvLPn8avRXkNPi9AFnc
mB8SDlcyyt9XEqYgPERbrGO1PwiTYi5OTFysuXFawUDai2luzYTm+6CFiHylsjdYoUYEplvOU7Nx
6l81g2Q0LmWoQw5GlF5Q8j5Wj12kvH69/oiZkqjGjnVgowrC2oe0yCh3mJH7S16SnfAdnfz+CYMn
Srp5aZMxPFWc8/zt1BD2wI5iWAa6j1XX0gAcV771lTK+42s/uSmL8dEF6AjXJj47mQLGgFTtfvK7
1Lt0ab6j9O5fBG0kimMusMpwbJrJJaJ2qmqMGIyomb8/YETJJOzPeB3zatCeS1G2E94++1GTEkPK
/mu/c2eLgmWThoOrey0uLdxeqVp1X/i6SmU/BQNRhKYa7PuxIHctS8FmHqg9dIkJA1l/ti4TmE27
OsIl42kXhMLAqwimr6C/FSUqL0gFYxf8zPGD9G1IBUDm6R3TfN0zLx59WKCFpIVWPl/1LwEWW2JG
e4eZBMwRrJ9X/A8xnXdcuP7gaoJwjv66F2XSB5o6MlUWfrfY5W8pjYgiron91Wp71U4/nssP3q6Z
6RwOTXx2y8lwdDzS21snQZJS/qujh+kAv13JUXp/JTPI2Csnym2/rj9bWxQ4JGvHqoII1GaqzjoV
yh8iX5MhWpe2YHCJ3ak/qIL396ynSd15GWbzWPIzMMHQo36SUYom/ST60trpPyiswqvtEFEAI38p
UTSkPzCbzWHwjZmVRqB5lpmKgMcBUphB7kpuwZPcMSvAkB7ZhGnHFqSrprqODGEjwCfGlnYSayOB
JqYbCdhmHfQ72lMpxOFNT5bnWCYshyYg5avDcmRQh6p+uOeGaCHIKfDB18qfs/7N2RE9QYv3VU7+
2Lkd2ujIY5ieUOXj/KwBVrTCF6e4GaBpUO750S2hMAu36MHH4VmD+KcoQJEANkI7HcqV4lgb+cNO
0d4nkA+C2sS5rp+Hu+GTL00DiEm3fWLRzXJhsMcHgn1qzK9qLSl3XpKROTdt44VG3ml53ZhpFn1m
j4flWFDtUXVuRaFHlza4h0nkJNg1iyck1Qv/By9j33LAi/75c52VmRa6+SiwThaCO9dPApfGCw28
yapVyVrZ9HXBO+rvc1MhYv/GsvXoeL4JU3byyhwJ/GbzHW7gNmosZMSPjRE/Rsi8L+7ILtX9+fFz
F9sMCe3Ufk3u30qMlV7nWU5DDOhd3TQEhzN91+37LsjEsK+elT2Ml3+7s1iDA3X1bNqiUuLm8n5+
H+Wjv+ZWLRjkFN0PhNE31MonD9MM/ClghIlMU7r3I22601eIu2SProPFTrAct0A6vaA88PXA5pb0
JBDqDSM6RnPhPk3R0MgvRuzBE1HK5R0CgtHNlFKph7BTpb5aJxKxRs0qUXo9dGtBc7QnX1OxQ627
c8uFIE1mEgUzMSIAx+pHMto6CsYJtCkkxe+la6dU8ZaKsFhUs1fiNT30G/KwE8ROawBZej2McQup
dTqjgp6u5VA8oPM6AlGJfh74Xy7wuR6IxhSlvAFR7JDW2TIHESDy5g1J+EQ8Jc1zkFunMUaO6tOJ
qzS31nm1dCaLCEkH6Rl9izmVMeJjNm4OvJ7jG863N78NXAtou8h+W8CIx9YeqR+BWOhMDJ7sJ3va
GG82IWQEUtAfr4dFT0+NMyCrO4VhjLcmHQ9Eg6tEsQMyvpyftnAzzBXhZlVy9172Nez35Bxhy1Jj
DriOu+FDk3UErzbP2mgTwaR4kCs/5cFEU4+jy9hFdHtP7lh9LnI0riJPvA8mH/d7DxmJRffnEjna
I4Qnlc0mw8MpHIxSdgz57FMdcywkdnI9UlqWjJcgD9Czw5L4tZzuXtrHIFXQO32T9ljx89XSn92Z
nSYYFtBlCEhTgMro9SY0gILZjNOUjS8UfvCdrdeoMfaFHBS8VLbeFeBQAcM/7FQBQi2Z57irEYrx
Qv0FEAqAcw2zXMnco6sw5slsx+/PW+pgHyJeTXXf66TSb7M1joYqpsOR2TYC9cV3ki1hcwsZb5C4
LsAY14hLMP9EaVHEkE7yva9GzesFu0lOWYvbr1yeub50gNGNqEjumzqfruUONfTYUbdA3VxodjN2
taltW2eXT/Uck7ty+fmpS6Sn8qKm0feEUqXBFUHBZklRWR54hvEO6yZFesYgFNiY78pkzlPDLK01
jB23wWtAjP+eZWjFDf2xOCzrFQ8xsRVQun9n5FPwsTRXKP6+Bvmr5kVxo5sZ9guzJYHoSky7Y2JD
sQgUaGf6CZrFqm4Cl8zKm0AKyua+ZGiNF8aBA0kOK4BjJpOMeoqT7kS4vSzp2GVZpakq6CZpt5nl
7mVc1bPqymN9QuxSGmyEdKtWdiXw3jdeR5rNq8Kk1OSPPuejG3GziFFirB4E+y7x+8E06gEalAFY
/UYKZY78R8BdtD+NwhrTPByTqEDJvD/XqRHtNO+cD7Y92mY1zNFkc3oWvNgV7xKGd8nN0gDNXhAe
jBFSp7dW8rm3VDIL6umoPf24sNvpmysTQqMTMeG9dgCn5XasTqDpqxYwCOOaKorfsHzpMYqtSn0H
JZkmCUEzsbsFOxUTn7+35Jq8h5txaPeAtQqS6pFI3GtMT9ppXJ40gezNYMzJvocYaMTgePQXSw+i
FJH93GhfuyNtl+gchAAJcqlW6iXzoKkr3uE0vAuZ9f878ajkSpcscdH8qg0MBhrYU8koSF/tUuk8
gI0oMx1vFz8sZmyZaygfqTTXXvMI4BlTUdGokb6izdhQ+eyf0adGFV0tyUB4I+N3XLMzQ5fie8NY
mQhLsyLJSVsFXp+2CMNzNHywa+/dMEgV/2WXkXmPFNamURjEoSKbsTEpDJzqxhBiGI4GVZ0irNrY
fW6kc1WmA00iZtd8K0x3anb9QPI627u8NU+7gV85u2StwHCnMsO8pnoWFbX3qf332e7dSK21P66m
EH9ycJH5KcSUj4TDIj0Y3J1It5REDVLlRUFJgEMm+JhBY3FoW5YRrqTrDNP2lPFso+BJSECKOqfr
MFlq8lcSyfj/QyjQohm1rgHXoNqZLVEDZ4il0U24houZzDpbqm2moyxa4vNJiagEAQk04XwS5lv5
csDPiQwiJK3gXMRLYN7zphjkjsyTqOJfksuxEBL3uR22u0elnHssW7ksxn/62+YrwhpYbeeIYo2X
SkN3ZQTGm1zuxdQ0am8oHbxrhbNjWuoob3PYsQza7UpX2NgoOqJbKLA+MlJob6t95f4K/zvJjgSg
2sjm7I7MBm8ToaXm7J6RN8+UcWeHtvmoSpiY8L6tIAn1WA+Vw4PCUAHJro7yAFbwzBGg3Bp7UMP5
I5EcsRNDM4VE2sfYSIR0ZskSOUgTutPs3uA6/CfQGkHvDEKJ1uhQO4KiQr09KseE7yeZfV97dELM
s0eCv+tq9bq9glY3LTd1IqIX/eWrwdn6E81VKgck2sJ+za4Sy8Jb3tzUTWorWKs5/XZWEo5kBnw+
T/D7YSwZpt+rIVsniTMIbBArsynZa+ESxy93C6Xw5WQBgFGiPHWBazr7lSjaCR5pzJEmjO55yxcQ
BTgoZDFm6aikmjcsB8TjTn2yUrM3Mo4PlyrS8BhO3cEgFi6m4r2IESW51LSED6pd1jNXhFkii2bQ
Bhe/QGQTKK5UhUxpjTGpPBqxp+mN70jf5LE80NRozhG8cvPnXZSkkt+qYSSqPZLTbchTwdWiOpvu
IYlZ3ffIl/8Ti6ObC1zKFVIxfGJd0qfr+eJdyaVOHx5zk3DTC9DT3vl64IYO34F+7k6AVrfJD3+3
hkmK75iElcFBRw0nrGuEp/Wu0UYbpdZK9qlFQSnJFvnpoplTwUiX1ALm3XXowGI5I1Znya9k8Vnn
fdOxNCZaW1DavfLRZo8xu5IYrcoCpmbgAeMslgjzq5vo6fNmIWCkIZrj+liXKxeJGIyvgXjubRJ/
qyxgWFOz3LwJGgma7pZ293UnW//X+vOPyLUpwltEMa1vfUhfyWX0LUhp73i6KDzLeuv+zrHPFBrN
0hjU48eza147WEmZkesrAGPlif6b7ZfcmeDgY9q82Li8isr8jKXMY7TMTq5COEVulF7DL59+ZQXB
VVEC7fHsqYD8ULSOvlQYtlgHMnsUzLvBb7QSVjDgBniUNfIY4gAkGEaNVbsee74py2YU0ji0+FbB
RG4O2bRVN/vJpz2aIwUS9KmY4KFQ07tanVJOwkJqdXt+NkvreuxF+TZ6u6ovQSNjCevzXdol/WDh
9bXDdvUQhGc5nsTqdh638Ywn0wqvEE4T6qlB9gEL8GGgwW2qZ8FkR7XC2PpQpNuQxd6IG84LsluD
Z/TiIE61YMA6M7/Pp3CcQkb8TGhS5LfIsj84Mz9iA3D3IY1iJVfn11TxBYzmX8MIM6Rt5VNGYrCC
RfCjvjw0nZflV+9a6FxjxmJEfPmGbUADGxYy3F7Oe2Zs23+9tEvYvWge4VsW/VAGQI6Djrp48Ope
4pOB6q3C8cJOEBTv1F9hWz3Q5ulK3DfJtCRag3eXohqQCIbIYwiGEcRFIJNCavnjQzro+x7ytARR
KypVi1YEYtFcoLiVl3KQQZScfOXrBS3lVeCQviHPoj4BLBylEBYAf2F6302JHixjParpNf+NiVx2
MSAyOzbUklAFq6GipQg6Wx1U7lMSVqolSuKwDz3+1trMcbMWzb1h3CQwxPhttayi5oiEcX+WWPb2
lwSjbcnLBoN4r2vbvcMQlXToji2Cw73EcwvlerkWgjaDLWgHqA6hYIv3OEaO8XtZ5ie7BgdTugSV
IVr8IFVDXhkF5C1QQfN5uD1x1bygF/KjztnN6vxmFsi5ui7Z2ahZYHd8c0iQjk6vmH/JXV7Bm4Kk
GnOzy2RyjfY+B4sH1rQAjEamsSq3SvQ0c4G0OVryMjKPH7ZIQTqAIWovHrK6e7Mj/aUJmO2/Dusi
e14zCXZCWgsPPIMX+aC7o3gXzKQQDjsADY8Fn/vyzsEfCazN7ecurX0Php5qU+t7u9GdK/txOnrv
1o1MBlyef8S6PY3ndIa4bxtgNL5ggoTJVbbGlN8UGAh5iPnr9Q2IF2tnbWtxjyyomfVONEDzpQ2I
oBg11o+fiKI/M7HCvLjPkv/aYF6zAH9g+PrRu7TjF+xU/butrz8h7ggF1CnrCjkdQB4xlbySv3i8
P69Ci9l9RU3IJh5MM59Lbk6s/YOST4hFUVnyoX2AqAJdjBPCOHCLvtTUNsq4isYG7pIYyp2cMScO
RF5HZytLMXxO/E4akDCmF4Xovtb+cJoq1EAxnnSHwB/Y67aV5wcjWIILk90dDQJUoy9R3IMeioEk
NpNCmqmr4j1+N9kh8LSCh0cOB3MAEVErGhg+geEnGXQ2Pe9SNsE5QVuffOARWhItuSGtDvv9EqT9
ej3jxc5+jHzG4HESM0Rk2N3FEvs63UFMfqLPFApRrx95BJupSYGlSHo0WRppzR0eo5SokT/o7UoG
Nt2Dbwpd5Dlcmtmfae4Gsga8U2qK6zOHwmRUehxdBoJ1iOhJDftHVPAexSIKRM5y0vcM6bDgmqep
XlwQHcz/xraiwvRvgJAiSVXZvZbyVOVLTEpUZN6enTAPQBIb0R8pmUSbRYC5r8DwTNzZhGkPRCRc
fey7eyy6++swU3+IPKdIwIzxe7wATTV/DpO1cDOdu29jYfwk7r04pX5lcu32R6WRVNysicpHNReB
1N14i3CiwA9mAUMY80GKYxYBuU9FXObed5jYA72ftkNQ17iSMVvJEsmYVcpsgmYORmwyimQRYIOv
bSqDiT9f9Smmcgis7IDtvclFBPgG9iyq08EtzZ6ZxOMsit2ziYRdw6rMmR1VwRrxJt1LZXMHrM8M
8JCePCklNQZ2FTlv19Yt1NP+ci7+8RrUgW1zNwZglL41Dg9Yno1gqHJlxJ0/+jCgcQzrP1O1ce2Q
JmocRMYLcLgSmPtGCAgfveiL/QE4gr1rrZ2RTINSeZwORfymCphZZGK/b7986VghcUDz9N5XaF57
GkbCURQywgRzW0457JA2iMkr/j36RSSS4E1JSVH3/VZI3ec2WROIq4F46QACGC+O3HZ0IWmnVnq4
en6pKmF0j1joBJqYN5z3GG+1haurEtqRMonnEYabm1JBBlnIcyGjzzHrw4vMjtUzccGo8yk6/CDm
3frryRhXPzxowsYV1WMH6P4OfHtzC5GVbGjXKyT4qfHcnTfU2RjsxNdZ8NXcns82gQaJun+0CI8w
GeWFzredFWHcy7ZZqgJd4tYz9kTYUoYZdGWJjQb2FOvSQGpXTGGLpbpf45Lrptv12izI9iAIYlQ8
MQ9x38tovOIdvCFcl2/E0rqQzhIt4r6UU3qXwvzb1+npipz/f5qK327W/0fnrxuNRffsOOt7v/sq
y/CJxrPmQd6m/5ww1CSIu5ubbQ+j///0T2w19clJkGuIQS0jnuR9T/OEOZFa15hz6uWsrIdmWv9I
s62fxGnnB2BD/E/qtk8pD5u9+5Gd9rkZGI2wgvITjBQ8iAVueey7TGStTAaHAtlEkS8FYBoRNUs5
ZB+rSU6Y06q9JQgEN/xXpsKWdUDHI2jMh8bHMdWYFJX1nknE3acUI+e1yYOP9miY8IpgqGM/ToaV
DSGDG2RJZSJwT4S5eihQk3VAa0/hEA4l3vFfSmZLltYwWQTY88mqAftd4ft5B2kR8eFdy68oSAei
6l2Wlwk8yse2YM9FRYrO4gSkXqxzpYCM/+ODI1r5HKQJ98f/KEc3yOuhYmy8PAMiteTJdlTZLBwn
1baMbcWJE2Ei0W3Z1uclAvTVfRgRAm5VfKe/U2CU0cZSQWWfsq1dKaylAkjIq1ndUIPHOar2cKiy
Ut4QRCTY+hOOay1MIMNZskl5nfQarucS8YkG/uVfQHpQjRgC+wWkGvW4qv220DWj1LGhfLqydhFq
sRaqJLhuoobrG+XJFuJ1/r17+VhyomShG/AZz1hEs9c2He0ZQyE6cQoQ3FnBDFmaAhwBnbBFOpYE
OS2ytOsabcddajQ75OPPUkXou895GV5YCQcO8YEd+gtE3roEEpuzUWXsRD9QVuavVsXJVBEfRVqu
GtDsqQWRkjmYEmrCvoW2kNMKSxnrO6kmM6kDoyDYgsDpN5fhjvE+VoNDZiAwcgRLHIiVB0GD9Y42
KQ6MvVGS4AS+5d80bjXeU4TMuVgXoo5WWJ8RHPt4Gc1f80eeBQ8UnzxyMax4AYG7rGMsto9f6/yI
a5IJC+ZA049zyfmYO+p7Hu+uW/qnEhciUngdhMRPLAPs6vQkoxDW+vyKJkWioT+EBmt9HCFsTk36
peMLvPWxW3GFTAzJhx47/hwK4F1RLyk062wZq7BdpBInau01TPKKXqIn/dCae9kgwXel8QfDbgBn
IIimkZD+aHWcLKGfFnnLJwmCpBRKAJfz4oREuStyEUrDltZlHxdy3Ap6wgCE2Yf/aLMed5Kqd76G
8ceqmAtoZfTu7qStpXgLPa6I/Ju3Vdr1nrLQi1ZsMR23cXlq8V4l53xa5TVdr+dRuDg9B8B0hEou
o2QnMSdBYO3UmOzf+N4ZZ6O+pj+MoKPDObSg35AZOWL+RXYdN97X8fGUqeVJGg/rYnVaGNAlId3Q
8C/h/3YgkVEGQ5YtA5AIYEUV/DIK5B01citKXmpXNLqD8nJg27m70l0gQ6hu9L4n9FNGbO3CgwG8
xmPS1j03VpTtvttKkIlkCvTyYJnceZAi9MAHdoO4nAH5rXmKd01dXpw+UOqMGPrlPMcVzOvyrcFS
41ZZXhMr0xcKqEChQv0wfXGwsTK6bORqEBCHg82yuse1SVSl366xlSYDclaZQEsMMqfl2LYn4522
VmDBS/zzSsJ+9MyBbu7Ejcs4Pp/nfzqmzgHjuzS4qluyQHEnBjkOQVo3uzbuwCU/k4HYdJH8a2Jw
5YHRSog4wko6LHMSC3/GOQRZzTrAT9D6InKAUq8z8sskr5WtHCga4Y0W1P57zpVwJ5X5NGpVC5if
u0lfjMZqwkJK1AeGsXNUChKHA9YiPgTEWFxaMc0y8s3HpcyC4c1oxCQ3RZnQRibZ4kIfvIaXT8vE
6RUkTaq5lBwvtvdLFo51uuQIrcoydcgzgtcl9Vtb6RTK8Lyl03626jJw0FrKmePMaFXXiBSiPe7J
Ut6H/PhtbVipaN32Y+oJmfKh6PkwNjzqJ5KlAhNvis9sq0WmGPuMHBQ5fbOEDtpVq9+Bwkn1faft
rcVhA5kKSrr5KOEYzj3K+mWEwstL1wF/qqR2vIVU4FonIFceD8AvKBFMBWea0CXZ/zhT4kX+Ozow
mAU+wkYobS6FICRmTKqZP/qaHSCU7ujpeAwGrY6QSISDKa/nLMFMoyzIRY7BG8HsuKTXSqZdMDOn
G7E6SjCf6gCFsDvDkq4VN6uJeKSMyDPuY/OLEwongP/XAg/9NIq5lBhAmM3XeBoIizVWKG75Hf68
/ErMpdnxHDgBoKaU7TOjgSLPZcp0EOzFqaABeIji10zaI994R9sPj6nX8XuhHtLFRbLQz9HsJHYg
eNRSVoICWEaJxywj6iSs8msjw5UBb0jDHYo6dSqpdp2pDwTYhA4iKoWCBOXX45G+lz1Id75g/ugW
3n2sFTmP58MoYqhxAAqckdhBNfTCuFcS8BlwWodeBLh7Azb13VS2nKseSQ8W71GIg3qdqS1vje8E
6UlSZsFyuNlLotBlRXkS+Zydt+cP54lUx5tLIbzMBNe1+jDMSVmX6SnkBMzqdwY1VDTIhDbHYcKL
K+cvYD5oY2NRLDU3sz0aYBpf/u1a/6r7j5ANUBG+us4uDLSscIy9K1nfmfEPGkJSy14BdMX7HSTi
kXS6zxd0bcvVreDu+20Lr3Wuyhm8s0LNaPsvI61cNHC8gCKexPPxQmR/z2Zrc3+dgnOPp+vV1XpP
lPfLuRZ8sqtylXj+n2viVhBUbRA4kR3eBzGb9dQJfCYyNb/JKvBCbtRcZ24DCGjX5YVfdnp7QgIq
5H4JgPv8BcJ1aa87jWHTmJNC7AOXQ4T5QKBGxugzKz+5LGZdjpAalwv1/tdAWqb2MlOqIpi+8KGS
nU4P+vK+WAyhD2B66jgMgrBHkSidLTpcqjvzOuj8/JPs5itG3VNJl4DhyVeeKS0vIA3W7CpMACK7
b0fMf3t+m3WAAGjkiNt9mcgkS2hv31vdm1UMI2e3U6gnfNwMJuafSAV+dZcXJxXpah9pM8hFq13c
RAUw8GBGD7I1uB7D8DSiObTU/cmrepMFlA12nm9Fo6WuHEpHQVp3Gi1laEpLDCl0TmNdfe7ZIQTh
s5GMDt8mmciqPNx/PbXDC8swHF2lASBrNv1TX6P2z9qIadugGKYrXmbZuKUBpPT/2gGnBrvVrFtd
SGUILaAmm7nCuGxF6HpQPJMrAtz4VKntWfW3bV7VxPO79fQC2jQtzlbjaMLJRI9siabqKYfgkE2c
1HcW6AlgtSPEFwtGnkbxEix707UDc6+W85bOloOi8x1tna+fYnaOxXdzz9MiSfdE94ru/hIL4o8V
4MvKdgKq1aaZgv4jBWI7tRkWoNy10mPyCFEEERv5+Af3bK8HEnQ5ME0wUKXOFzZcbafWt6/W90ej
H/Ln4fb0GF5XAgt533y7bDZlRbryU+nysCaPbLULvFl42s9w/IW3VGbDUYkfE+BmZkSGqa+rGqhb
TTtDJFg4gZTPJKUnhBBhIlbU6FGgltC4h9/9v0n3LVulyseI6P7t8mRy4OGDXA3pcKS+Z7jwwFdg
b5synUwnYInUcqRV3uFytda0HT7GvU8NRPSSwYLvtf/UXlv6fSZdht7IxuA9ZvHD//yNq2FSZSpI
ocOll0kB5+kw0+JJzG4r/fCuWIt8qH9pzu+0OdfZw+Y8tUgXtT+AxMMaLRwetO7x0+ZBhoilZyA1
w8hgKoKi4SNLg9mjt5sxVGh89kgRNAkeHus0e3LwZNGpLZD9OVXkl5FgHGjuCrGHNQ8FLueai9DZ
H3D/U6EM9fKTYdrrbdiIrrH9KVsUUyCsOmO6GKEv1spBueBz1U1o9yJx9jOXmumsxEViX2cvpaba
iIkRJNEcknA6baRvIdOyOxTYTcuOsz1TrIliMD3/U0GSFXs3bleQkXZm699zzeQ/4zk6CjuyTx+Y
ot/srlu3OqyRlR/JSwp3Ni6iCivZqCJZDqfppip093ek8Mx2MURJB7r0ymi8TtiFesPleaGy6aOf
AHEXz3xl8SPfDlXTuNhYt5zSFneyFLoqA7Bg6cYhGFA3/QKGtbyuzJTvrsfSDy1fSLuOoaxxnGG8
twywJLTXOPk5lWh8qiXrEA+mUvN9cJr5596wyV40A1I7EmP12uWg0cJTQxO11spkuWSkqJ/PUKjs
VVnm3MyzO84+aXFyXbx3QYg2MfR5OikGUSwjkNaHXnTgiXYcA9pn6N7zwuFg/bZKro+UsbOSEB4g
ZsWI5Qiz708lpTLj47MOl/4S1jL4YgIFaO5tjzDEFKLMjAyAA28lgRMNMeFpW7DV23ejM0xx3SS8
cxOfmvuC1JzR5cF1o0DBt00Gtt8/kbbSRo7C5rvF4hi705lFSGyq3PyEk55NSddQGzTnLlV4cIji
glzpKIjZ3OYXvAQkwS8kXYcpn4n8dY92zLMYsNjwgIm5ZSgyd9keNzLhn5OwqSqAW3acBw/kEe68
MPMi0M8HT6Iv4ZG7loPTxjU2Qt0fR5t6qHSHCUaGUSTJcqjslqI/fypqbmy2VuNZSLERo9wWk305
FOqVT0rnTnSlC1wqXjX+01yXhb4pc6BSZOkdrd1xVdCQ56n6QxUufpIeoCXFzgS0EtSuLzdq7l+T
SwCy2HZPyqL43x4ySY45zGDQoQoZmkfidu8Ce12rYHgsU48VX0QlN8IgY48BeQAqUwISFY+tfHfk
my6rVEG2aDCFqCY/PfIjMQEMw1Vl6x9pmKumzpz966y8djElzasb5juWcjPE/my7/o39nnxGDkCf
WagJF0f6JspfSb2mJ/IUgl1h5Aa6qPo3vDuMnKzH9WmDzSkOYJbWBpV1U2wg9t9qDRYx8ncEjPak
s5HeKuD7gh5JCvowFz3MsR120LTqB1Em557kbMOeeQaJGQm1VyDwl4sUrZbLv4uXlzZqh7JasTH3
3Xa9BreWqBzDA+Mtr08fy1eS/q+to4LSdaZwjrvPuqHt31JGILlpwKWHOm4LBrDSfyara1Y0z7Y8
FSYNemiZIV3BHjXAoo6wh9g+BfQG/51mfzlArK3tOldNCB033LO6u72UiGvYfV6YpXruFNdzNSVl
EaAIc+utsM/1ce5KUYETsmvLNyl0KkUCkgk+KTy7Ycaz3XruD2hgA7Uzf0Mwx8XteUcVIWMpjpWO
Fc3w0cUx1iHk6wYcpLJDXex54/A4chq+cEyW1yaGAPeaRgQYV7CsxQA3JuwrmHQkOQ365E3++2fV
c7btaNAUcyQDnkUG5hpHeAdRn2c5rU4/WneX+If5vdidk8BzrbobiVUqsZEO3/mhLaQFFbOihGQi
zUIfJVsCfsKQAiM7RG3Wpu9YWpzfGnOvMLqurD2lwpVmaqNyvsyGlbOBKW9ZSlKLj2xNbZkL7GzZ
LzqLwQ+ju8izpGWYRCOKtO1aidR250Al7z8Ai0KcQV7U5mxN6UGo+T+v5xjn5OSRFrVMV/ZXxS/A
+CFwe3ZuAGfIyOz9jvcootqFl0jxCDWHzKZdUC259zm+/4tD/MORj7LRYB+oCAW3Ua63+Z3enATy
Guzw6VhT832vJMmLh9l1UBMBOzIYMlTT5TJ+8Gl18gCylenJMMDJ8PGstIMmYfxCC884SkzMa6XZ
4db4cki5WHlgSAWEh0vlJsCLHntSKbh8bAM4aWyx26Lci6tt5EBqSwHBXDeb35iTIKYYRFyWlCGT
MnJZ22fPBhqFcH69MljJCS5HdU5bADO8h3DjtBwL+xbOf54eQfSmFh+GGtIQHAvbopZZ2nTN+TZ7
ymQws64OkZ5e03TRLUYIu9/IaLj7DM4nWa0pAWyCiW5nsZtAfYXrj6IETNyCYoN6aUI+7lyRpMXu
PRBP/G/PYzuMWWPAhd8Rh/uhgwKkXkLhhIlW2lA74PMaOG0Q1VCO8k9+gsyi6scIBp/cidq5pqod
iZbmAOhAQD0wNlQcr9ZzPuSE540KadyI+VO2fEfCOWpcn68br265wGEeHLyxZ5zafA4T/T/gn0EG
4yQMsrX6bysfkv5dEj3g80HnyXYSpnQRZFPSWhitI0TR0adptV1BtJM6iyYI8mIlAIJnR7wZE1I3
X6OYxPQivJpgPVKh123bjl7yzV5HIe2Azenqa1NluBrbKKTzna5JOPTUyMYmnjBwLYm/x83Isp8+
orY5R5luhvs6rmzxaHn8R1OrH9CVP2pULnZYCDYhW+UQgohwKBUgZ7XWDz08YoSHeQnGUdS4NEYd
UTTuM9+zkovfTU7+q1k+wkvI7bY8z7kwET3YbEFef0XkTPcx8rHNnCPeUbgmhIEPZbKN/wOpi7x3
V3u2OXWIeuHs//zjxaNVpmPxu7gz41dYyTFf4GMqi9AilQ2vkSm8r+U9sJl2e2KkV2s1uLxpm9Qj
uOvvz4RBgzuntELEEOj+BfGoZEkKJcCuYTLaOZlfqMWAeR3de2nGR6k70OCQXUKx+boxjmqrpDxx
sRFCVH0E3q8iwKy+Ko4kzmHvDtM3adGO2JqZDUEB4Sct1k4/rTUsiEvf1IlPkJ7MYzDTCWBrwDrm
4dFyUx2fLs+zs+OtUuuzrwdft+j2AtXXhJcw+NLHXmd3GE5VZZBHzXiOxqDqsF2ImHb23LxFVYuI
s9dae3LE85udZSYkoOrG/I74Gij465v/I8JK45RT+njiTZKERakY/UFyzY4no4fs8kzbkdESeZ3U
aBBFphLNmrl4nPAPkhxzkmdUXg/fWsr+62kDEVjRZoMIHhgdNoTP6b+MXdz0vWJunXGH+IgIq/H1
0up+7Z0duviL+RFy0I3fRczY/MPwmCsmEzowXj2OpNLBPRwVu8N54zIlsDYN0hJsIQ317OhMByOO
u4hr+bMfmpjdEOYJa28zRTBoOgfQBH61nbfX4EhIsOXapgkBmla8TFLP5YEtNv4a+X7Y41Dijjwk
lg+EOnWBPpinbPvrUr58CUPES1NKJBDOucVITlEm8WAE1pIFx++lvlX4lzfsms6LnZwN884W/itG
NGS9dPSnaF+2uzjt7sF8HzMYyA2gtWIML4zz3nONNhq0JaXXp9yxtaI4MaCiaeaSpKf9pNkzx1Iw
nwQzqV96CkKK+wmgxB+y2m+cvXlryNnIuLwxVd8fTw8TfTfwR/xqrejwBpguAFwTROHsxJzQBZR1
OPMN3OVJI+A6ecrWCPUgFA8/5PwZXDNAqTjK7cDtnuYPkYct/WJ5h8tqgqUAa4D3+MmuS+CNakZH
EpjFSEjcYKn4LcWIe1r1BrFZ6k7m/Pg86FD6nN108dEX2lizNXedxpJ74DA9qaaRk3YqoL3kXY+Q
ZwPYHV1avJs6nlpnD2xBG3M1KROOVkD5VGrvpeoteBOyUOJoqd0l+W8Fd6ftf17gXsXCQeFLrRyx
NjZTi3k7i5UlaKRBW3U0k4B+0k7uuduYfZnFDOW7VYeB0oqJ8AydmhNNwGBgaxBD3WgzQ2aqZcMW
ErpaCC0nQRPmJuKyRngiB+cAXB1JGhrqjFCzjkP+sGZ9kFBsuGkoW1z02f/pFiDqUDUeIUKRF2nM
hoZ8NgF1TAfRWXCYwZCFCO2zlcsGtjc0bvnLS4Gz/hmxoSbHb3Zw/j3HLuH4AkpplaW0NUgrKSsD
aiY0Sr3dPdAOywFrkIlrO7Pw+/HC3nhFvXEEW2VtE0B7qcQO4A5GrmgDGfGvHoUaIUxRsrD3B+qt
QxF47KMb6UJDTyTJO51zAA+BPTabS27o9vNnI3ZLNTfRZOMLXtMRrtVN6lHC8RmPYHmgX4ML+YxV
5/etd/NPoh8Jb53TzEbp83/OyJ1qwlfTozVqHSmwGhdNDD968+PDG0g2qm+WHYJ5gSncLASLuKea
jtaOVhr6hP5bkZ3vM8NbGhsNazT0FtubSFsd3S3ONH2VXsngwsyZclUKdRzgYoZMb8MF38A01JhO
mjqGyALvuBAyauujFWrQoOsAnP+P5/XVwnlVWpYHK1IhzS7eSuBomqJEjrpeQjqpGJ+QgqQrJDLn
7lQ9wJ1xJiZkApJhJY3kLkdqf95gVY80eTTDgu0ZLwKfcgAVnhFvzeAETIIrZQrJK6QxDKrpS7IU
YLklH5i9VKm80Ikpu8QM2R4u2zRpi98lSqoqDuToaEhrmRW64as53luDhkizkTCb1jxJ9s2kJaXr
t7Ep4inTPUlCMbS2rfGPznwY9UKz9O1mWuPuhcKweLRR0vj2/kzicoS9EuluGABsGX+lmBbexanz
5ZG9w0vucYyuatuFFsLUfPXw0dnUWNp1Cu6TyxJNvS44BsTgCRdKgWKF663oOK7OimrRwNqVt8I+
RZS/jlkRiHWmvLI3GT3sKRDsReU/afUJTaFWwrVhSuYg+c3XYnHLCZKd3eVh2AL3OU7oOU/1Wz4G
ViDs/r0uHojzmM5sjHMJIOWx8KUeqp7XX4yJpTyTp+e1uQop+6r7+DC8t4L0YJ8Hs7UpVoAJG5sY
FZXhF5bh4SCE4S9AutU8JGhIDG/4zutJkaDRyB4Jjq+GBsPk+j1FSn7WIA10esKvJftm3INxk7bT
VCZQR7Adu7JHI8FYGdRkB4s5H+1gJkqLJzeRyAHOO9QTc5HTgBM2g/bqYlfgIAR6r64wGvRq/2HN
pxraVKGaRYBT2yolDCnbZLiBPsN98BpD7Gz7b3+93HLQm024/NmWdK/TLXvVF7u/qiLQexgBbGT1
gFL/9zGCfnYMgB5HUhK64wGY6cRbpUSEQaNUj1yWm9fxMnsxfaLJNW6bCosC8s+G78OK3r1s6JoF
LwfmGDUWa4AgtulfL0uyUUzqfvwUcqdyQcKDpemtpQW0Il6vo/DXTr96HlYG+mI6Mp+MNPt84I4p
udeW8MqgGhQL0r/HOFKiuTLNcIzM7FN+2trthMhmRPkO+b8LrBPLMd2n0KH7Ane59AjUcit7Vl6h
FIquF+cgcJGLtkOeYI+FhBP8zoX2FZD664+QmUHKMFbwUu8nmE7rSxFXKy4UealF3frlB7VeZFdx
kX1cTf6tg2+WwDrEctci0k4FbhfRmRV+oUemSyIK1AD3JsGTw1473fsrr4aRrq4MvsAcOmmDs863
5GKTG/G9Ihx8AUm9UNyw7cs/M3azVhGFL+YKmsOOmUjXcHTMyp/UTc4Gq5Gub381xJbjQaNx4eht
jhTCyNpHmT0lVbhPDctOrfdpdb2HIscg5Ff7GxJyyQPK97L1CMRKhmca0L+OHztuIonM1LUMEOcl
T7ta+vy7N5M183hQMvjD4RapNFUjKLo25n9pRgGoMzrFL5gwTA7LPdg9I0nDZSDraRG1BsbLRu5u
P+83vVzh2E0hqBWpApxYshpTL+X3TIElFOlJjqYVMqs2CtmQ0ZgRkzezcqRX/m/rQSRswhvu1g+G
bhZF1+c2zXz3ajfIxfSSRPYFtukBJ/MVms5oodY04KVcFId8CXtRbBMwTRkbCfRhezJ1ugGmwIEG
M5Fsr8CtQRy8qMPlajxxikpzpR8rAbfttAOlaRG4UDgzlTs7tVzcFzbodyU5iXasV89wb0MoVWvs
YQtXWnbL0bDlT5mglbDxXX0qy4p0qT3a2FD+5VTLhwldCho2AwSL95RHcqIKYGI0Dq6Q5avFSk8z
pe/YVfqbyUnp8v7wdDmnKrW3kKZV3q4hj+diHYMuw4/ByWa/9Rx98lUlJIBk8zzH6b0ruiUAjL0n
mOZvnJxe3wsbYtHfMnOI4W4vRB7JlSZWyo2EeCh7fMJGmviqqFq2OvPjagKV7BlWafn8LPiJ6r40
LSNyFyVlGEkszH3/iPehl9Ade3Y3zzoKdNo+T7AdDVw62xxnAjb66jLi5NU+l16g9KERRLz+nWdO
v/fcjwxlK28DPJLtxU8KMckDnT5ijdvSevx25535gybXc4YlqEeC2donh+kamgOyL9SzSbRpnWn0
dbrXYEFw+Y5sxcajmkEGPH2guaojFJCh4MH7O1a64e/FsuaDgqzB3c7WjkBSMauxHdS+afDYHuYG
CpAlUBfh4TTqZFh+kpWCI/xktOOmAKhgWZIHVXD8AH3Jy/hu/qgltFory2neIMyCPPFIJ5Mb11CU
2CBZhN5e7HXZG8Ut4Jw42OV15jfZMStEdpV17LH7V3pZ7m3WRWo7SurFD9iNU1sK1OOn2krDTenE
9tJC7fKshHjMKDrrLJP+UQB60uwKZitxOH+joxriHqRZes3U+4Imqr5GcqY+rKVVCnnKLSqILEjh
xFDUCVR8X1krgtAswYL0I9+m0hsXEd9RD813w4d9P9F8ovrlAAr7aqS+cG1oRqULt4EAXmHwQH2g
VlY5SF8fk6xWRTw4lB+kuaHft+Bhirims+9G0HUNjR8Y/90mpvvlfK39dpSVkjQnCbTqlPTHImXK
g/SVvlOvEZvDn5OewkTWfFsgv7cc9Q4AUBj5gvoWENULJPfH+NyPaxeyuqU3iJZGctA2xTJkwv6A
hO7He379SvLy3M7Mc157pD1OOYNMNu5s7D9A5XzqBW0T3wu1huG8hl7az40xcNphZTd+uDNrsxxL
GvsUZtDvDYMaNacfg1MI9gB13qbLEAKawT9Gb3AmbwurSiXuvMWRida+0xmRgZHWm2iMX3mZyL/G
3cyv92S8zU09TbsItHxNLHnAhZ2cCNpdndNCCMfBMr/Nd1w2xuH6xa7zKvxD4OH7tQz/aHYU1pm3
MqRXOWy/r4rgUt6LGUPR/nj72aFbFmcHYD6FJrhOLcjtknAvedCu0Qqyy4s1ZKe+T7UMOu4MELnN
pkh6FZo1vqnNBgnkmjteM/XYhmy9mMqlQBYS3Sw5N/HJAK6ywT6s8yhTkgiJ0XHdQVICuI0u9EOm
SfY23jtBDTX5ACfp1LoEY3pAi47s+6Y8c/J+3/9ABVi/mSz5bLiHiqreXjdgBRfnIGRIhrhB3vJE
fHQcRhQKJPYWxR2k1dv1TH+ywrAHX4TOJxjnc6EPdOlK5qLcx1Gc8GqGIVk5yF8LvujJgGCj+Wne
83hRZY6Nz9tz0NoZLVkQEnm9f1MD23WH4DF9NDRZR94SZd6pf9OgbQf4nZlJt+Kz1NvKkbpxRbfu
vQIX3my2zTg3FlngNAjavL8nhL97egIkoNTw13TghqwA725zAnkMFWLFwW6x3fyYGqBP9x5gMK5i
tCVjIugC74j62EnQKcLSJgjgQCHPpaYphtECLExzF9QcIk99wxgNkEvddTz9suvFeMnm8fRlX8Rv
ksbCYrIXqaXEeoNECkCpgFN3QAOAv9lc1AONkfY8jgJxLR6CH2xi4IG1KilpRR4Alz3EMLwJ55xx
2LVhtV4a6wS3a2JtiTFbOH7Iq1zrpOjvbFCjhlj26IXr3Z8CIaaVk5/AdLdYfGrwId2MlEQmpK/s
mbiAFoYlaaEbArvqTnzD1sP+2e8avNzD4kJaFNdwPuj0IZ1r5MwpRT0VGNq92tkjRCxY5YwpK3yC
7955V39STCjZnWE1vKLUMG678DsaCaCuWgoxGAbOduY9E/HtUnkX+KTnbYb2twRvfD2DMjUMNLcO
CbZSWEdpA63Huz6LYzQs08gQSFuu211Ynq1K52rq+69v1N4rxGP0uaZoPJWY5M7V2zpxyQoT70Jj
1CAWr+BKvZsAWzlrUuZ5Btals3jpZUw5GmDBSRH8qXKyxB/iOoOSyzOk8rMBMVF71dKGTZD9ryvN
UzeTVM+QXHh+6n8KQbRH7NOR3IziVfpBMH94W6wfSovKDdY3a1U3C9qOZOajS5EBIx/6uDIrn6Sz
eBaKJQtkgEilMBiS9erjayCfAQLKl/Vv0f08AOn5bSD9qONYns2TWLYVa9G3/n/Ntsu1od2molTv
fdW2pSfEjD5NZMjIWtV0f+xkgQmaajjjoO/d7ZEJUETWBIW4yfWDRZWhPOREO16CihEBS79gsIQO
gOAh3bL3UCS5uzG6sI61r+nYJLsMacXPTlKedrFnmtPK22LP06r4OXSzOhSgA5zlEQMaTkp53Jbe
gGRu0/dXgykI0JBVoQ6hAS2dVMsH5XKa5IZpAIN0BG9+OUrumzbJ4/aXb935Y7kCn0IB1hf8SBCr
PDDZ6UDa6D7PtlrbAg2eR6x+wBo7SQBsOhOAgUX8ZpQkVz0vAgZ7fv7HikHWEbjm8hdXVD7sQMdI
xqhjWFsq27Ne6EwBU12yXMA1m05tG4mtXuoSjrf2rpLCJBsIuiBjgV7+Z67kgfExFxo0WxNvyqs1
tgeQj/g7bDXu4vjxKI1UItPBJBvDMpzGXlDE1+E4KqgPQt4eWh7uUVbPa0oD2bn4uLShktvMFOKf
Hdmg3yb1N8r01aF/0UgQwiTeE4ycQ6yS+sJH+3pHVI6e3007yrha9bpLiNhzPh28YT6NvlVcLxjJ
c7OHjlv0zvpjoaBhCEGvfV17bR9MGoS3xW1aMbWJ1iExaXDZQJCTuO8onNQIfodzN3n9E2884nnO
KbpC6zIrFM5y2pCqx8FQgdf5mcRZeO+UWGqTtOdwovh+0NGGFVqb9So8fUzP2PMGP0PlX2hUPI+a
z8jLcXv8KSpqOghM229Bky9XH4AwcpKIGq+2eKmRt/M8vfnQRd0dYArdZ0S7jN9+O6b7d2002BJc
qS8kATpdUVuEWofq9uotE6bOzDOZLl0bV2Ajx2/u4SuPkx3REG0+dkNT6ylU0kJAg/pTQYeL9bJh
Q7WmGI5zxinadDO8tymtwU8N7CFJ8uKBM/A4rDNT3HbH74APbv7PNgSlsIFrjiXiNe/bLMBgreyR
9qcVDhLBODRxrfv81vvh17LyipgwG81SqpMzrTYSq22mP1tGHDmPg3rfbbOqpBdWHPM95T027Rk2
HcAXd3fUhlVpn8bacT3Be5kCxy+A73hWOKFper6A1MhedduhYsP3ft5puCIXWa60oJbKAkAYxyNw
peNc1gs1WKzg4/F2CUTLgix++znFj1jp1hfN5XjrVG8H9kqla4ZUN1oqEXpIf3hTJjNIMDhdN14G
sTd/QLl6chOJIKQ7vwQxbuN2YWY4tHHDP9TMHbDHZTnZrqQUVOfUwR20wjYhIIudgwfl+U1TVxYn
Z6LhagDlZQAZfUm462bw7bRnAEoQHXLUqKUSGf0gpueExwOPUY99ywKcHhoADAFLoDaUhGroBSqO
PQVQke8ysGy6+q87+WULfwUyDjgLlw14b8lwY9yti1MkyLNmW2u4rVtrjv0/5LySWAQyNjAULYhp
pvQJGKEaB0TGrHxBALsHNCbCi66lLlq2AkMSx6UnACIGTLd6T/7KcGaqaSXo7p6KaXON3WNWEKmP
Zm39Z2G0+bb6L6rPhppxWsk0QbYoHdk93McnakSs92X6OsySsuO/uwAyodgMj3pqffOkEc/fXCgR
qsokgJrP4Wi0Kffuxo5R7FYAl7NGRsjlHtFwk1OPfDZDNb+s6T5+IUu2vTtdvQ3KsmNxsLIf4Ilt
1yU4iBcAfVo4t9q9PegKcoaTcG6MoEMVLe7BTp7huROquREECBz+MQ4yfI/qv/peB0vWs3s6Ki0m
X1ZQXPxwukjcZks6OAiBPkSFrfG58dITAqWA8zHjS+E24JaiWJLewVN+7iyfHq6VWbGvvMf0c98T
7PKahAAII4LVzAuPXvHGjW0jGDUfvBPnQCTimcFeDMQJWbqaA7Qvor2/KdX3Zt6IietxOQGd6eL0
L5ToLM0tkB2o3sOuMXGGveH2fx783VkAbWDx1+ZAp47rD+XaxvWoG7KpteUbSxaMPZgQ4sYQzm3G
hNjflzR4X/lavsJPVn7i4pBol80kHZuXZJ5GYzNJv2OScRGFsqVOELKIhzLwaMgfDJ0agMYkSsYi
qruV5n+LE2XC1lPc7xEHN7kN8upd5QIuvDd9cEvWewnA5A2TU+AYTgU0ugqA25V72MIV/Xbjv44G
JRIQ7fKs+yUb+aLs/daBZ7ltfipHMvbgVHJSVcqfOfj3uTeAChKOLY/mX/k53OwYtaVMxwJ6zKSZ
8fAVOVqpj2hM5wozVZpjxs2QAqEtfJ6EMrHWUJ1BA/Pxx9j3hBz5XctEEur1DR6CEL8LUVXxkR/k
FbJGlzSsEIIG34c+P8F00a8WdhZ9YZ3ghFHoq3kmZA4DrAnexoZQZaFtZNBvHBuA7h3Ghov8ttJo
XAVGrc0acSOMkXPTz9i4SwIbSOGUImfNOwbj5LnDmv1g65M8JO5O+haQlkRuwQDk5/1GiJ218WBY
qSa8OB9HfMxvLEFOZza35gWYShPPwX/9A7zgWOmACHUAU86PTsulhzPLkButkiDl77+Qq8ftkWug
PTXhlGosoWNnXgToJg8NQEvbjQCgCrgyuy7TkuJzvJ73t7NF1hf5IydZ0ovWojwhaUSil3Pl57Ji
OVHIylDnlB9dXc51BkOYrge6ILm620bFDf5Xqbq1ir8hjT6Z1b/RwEuL2KckhpndccBILxdU6iyj
atzInbyj0t2VyA5bqXG7XPdA1HUtO3poDKJXR2Fvc9lpC6YUhaHCJbN5uooIeogGV6WfmbENxdGG
8LX7QEnQdQCk51ifwDdcXRA6hyqStqzodIMsNp8v53XvgoBIYp7PV/eEMB+mtX4aiQKKPlrUtTiR
IUr8c7cmhG6yUs1T0HFNJ263KRd9IZpxhupoxboqr/ACdbaVznHMJ7oMhuBmZvFhB/Cq0q+nvR1q
GM0iOYVbM925b0htN6idxCYiC4YZGHm9Th47S2SXefW0MxKqZbRMIjgjl5IjpY4f3HUjPCA948SO
RC/F4xjjbH2elJ6FsJRrOPuaoZADyGY9RtQFq1JqU3hPx2aVy76Q9DIEMVi9Aqh+mlRnUtyoDxhH
FWfV++89U+ZczXJHxHFdZhTxEiqEP7kyIxb35i0J11UweVyZG0BK/y/4RUjJI2nxGHwE5wsL83CR
lqwqNtOIgpoXbhdVl9eQZRPE1C47oBTtshlbmQT2dE+d4o+AEVfSLJz+pfi3Dl18dANjedTOJr7b
WyDT462PoYz4XwgB3t+2kgZXDMsCuq+WJtysizlCEBm7S02IVpVcCSEKsyVYsj4LbKYbVfHpODZw
QhFefBnFpRtLr7T3I4mADyIYpOZPu2DaR2oG2gwUYdsC0AXSUGG57ykkZAjVyQSrhj+/OUKo9gRH
7jlrHPsydO8/O6Kbxb2nZH1GRmEsBitqzpbX9cd+O7EVpJ7mQbXrii6mzQ1RRkT8dj7iZZWa3EUO
mTJDalxkNXfLKCbhTCW67Ui7BkPsicaZEaUDpgByaNpkac7PoRlj48WfZ5EdyU2rudM/Gdt0N2Yj
Qgyc3GgSnkwbTmWpQ1ohboL2d7nAr9CQy8tJU7UeuV01fyoHsOoAIJU21MERDGZ3R5ogiQcqRAtw
MeIhLN5bfWmw3pbh0R/ShB3BxMXdGB5PgepUHfZUwSYsr5aqnXus2xSsjmtJRVvgidHBlWRoE1C/
aqB/d6NTazE+5/+ziZxRDQ5IIiW7o5tZuNC1EYxup0dxeE5yPbYqNIDCBlOhtWzehoL4IF2pp3wy
kWt702S1xRHNWJ0RKwzR+iM37IjtRRx2p4Eyy4JOt8ZyFp2ORHTr0uDgIikgWlr/kj66szU/pdpb
O3nbJWeKbJYrVMBvkJ8aE4PXY50a6ziZq6iQlSQCRiBU07mRAg+qE3Zb0baAvgmMgiyKJA1Rb4kH
/npZoJHOSE32o/o3aODAYLvJ5L5OtAm8PHa6Xk+VSe9uxhilySvooyEji6DIFBOe1Iygu+Nyus9M
NynZC7V6WgUbwUtByhwdTEE/iaGSCYU3AagcVGxCEIs6KrKWo3IIjiLH6CaBVIHs0QKbmYDHzfGB
ZmmVMM7KFnjSpt1wrSiOUTVJeGSkVPtWjscAtmiHBdNe7oitDEaEs8mSdo+l1NbeeWqea2MxcYlr
DsT8cdqCCMUc+3X5fJtqbmMmmKYTZXyjwtwT9sJKQyaINVx4+59rCf52K1Lcc2xO5EmoUyT7VhSR
S/36Hf2rkpQ+wwNWg2umuUHHO7Eg03cjJ8x+NpOrKHMfjgL0lK/Ms7a57SV5lQfBITUgXTFwqKnz
21WyCmHVlf5zZ3Wfw73qHMqd+uTvkcSX46HwU7LN6GYu6pv7nrqXGQQmpcSz96/M3lZ5ugM/+cVI
7ich9lPSX0YUGppnRcAR02swWHfeGnf+cYJigB4ptwMmJqg38oW/T/kVWi2DoHR1PeEKfcwGcqJY
eCYZ7DEMpDge7dTtEmFx6PUn6kaP7Yek6xcn1FPrWO66KUg4VjnAk2VmYxVhjYeQcEdpXn3XAbE4
rkHatpb+PnM3AWLvsdjc8YNwb/hMpydOHTng7Y2oD7rxCr2WPSFF/q6WTHWKTVczO6tSX8qJ02xQ
Q8C/37UX7mA3vpAdkL2XssuUij1Maiavz8SGgxKC+A+EPlIXlWdYWt5SIq3kGv6GaBy1OSKZOC63
9R7KFPF/JUe6JOraZMfjqSM+84bGjKiLzFyLHZbBNfZJJCj+3Tnycm9uIAL0iz94eRbHY8oDWw6A
sLuB619BZInmhBIERpi11n2y5UkJJ9m3n4Q9wl2vxrpLh6r24M2H3BKsq0GqZ2oaijUjWF9d0mng
eWN55xYc4yJkyxWSQlzDoP5SLILz0ax5WXJMt4yNp4GW54Fjyf7swjffja/uf+BAjSqJFLb5Y/Eg
cmKhNBAvcduJWgW2SIgTIhFrEk3m88Y+0y455W3VwFIfiEPsNTWuZ6gapu+uZQ73JLbRa9J49ke9
hTv5kF3VryqzgahEgKm3lmwkHUV+ynFPigXkSBbPZWa1yfd+2kN5VuWSgMXglMlreiu+ynhpGtVf
zYMU7XYO7PkH94uGnlNRDahZXkjgZWBB5I7uCX6obXywWZFFGqn14NrHq2H2e9WB3k1hqVzTpNyB
okSlLhM5fL6jd6kpot2OnBPVGx1jJ+iHKTNtDQFiXcaW5Lt44DtTvjjEUQG9ikaTXIpb0jRNi5eS
WwqE5648cR+KQyH2ViF0E3iYVq26fqOkLnbiihxV75zcwRoTCg9XgeaLt21F4DqY8JcElFjAbY7Q
5GgT4Y0H/sPdo+bRDwe8W1e96Jgnbu/NJtHOKGdX6wH0K8GC7/zxgoKRtolAZr1w8bagYssy8vRo
jHO9KOQy4YPoJ4R+35lEW+Ca6OHlJN+mw92EVq1oEkWnY5FI5geyiZjGk2n91dIu6Q15jfT2Opph
fpdcNhrCqfQ9i1i939Tby1vO5hzv65QpBw8O0f/SD62jmUFVz7jxdLJRRYwkfhURtyum69Mtl3ZH
V932qeKb/PlTVb95Ac+Jfu3GRZLRzseUeNMA5MO9TdptX9bcJDdr+FSW3e+aNHLFnNrc4mECr908
Mo6tZamiPuiKubuYX/VEqgmSUJ3XqqzECUo6Q/Pf8qMz+15RV2xENGHQyAJG2/Jw6Q5WzEXDRj78
TlNZn9r6I2mR0etTqcZkf29Ih+CMUp6X0G7tov68IdtQJs5ot4rp0FgmL7WrprRmQHqoBc9RjeWs
P4+zZ4oxziZ0wJmIQCmzH4zQKjxycr7jzT0bVJdTXfXcskOqq6XULNgXF5HpVcGpXiwV8my/oR/J
LWiSy2Uure3W1K8dxyfwWbESd3eROM/LtzFRLpwSmwfD0FT6Z/JfiTRIhm+am29Yag1sLaKoBNtj
dLgcFSK1kICEqbciLz6N1r8eNbkcTaawx8Jobt6L1H0u37B1xgG3r4n/d8Il3mGS0N+NbEawhHw0
PNPmUFybtPPQw7zIAKSuVc+2pxbFWy9WlY6hcZWUhHTbE+tMdRKcviht6STEq1FJhudzWybvobZE
V68elXJuiWG0t2ymDh1emwQy/gECC7oigkwDAmItyPeM9DTEnQbmKgJtZBAmQOf4m482rtI1xIfr
vr8unvY3HxSThnea14scy39zo2oxCqfXsLeT/dOzgBDx+xuJwDZWiH29AtrMKJUU3cO7twTJLw9p
duXScTmCRFdFYhsDXMmZ3bJWr3mNav+6w3w4NiSXkK4+qna/AtW/pFZ5MFKYFADj0JOA6kVIBjcF
bfmcGKCNtSMVOF47rzs+iJqLXea08Uxrt0al6Oo1x1NHNMfu1Safl+NKOHm+G93zLTkK4YMi+SMV
3vFZ19RssSrxuz8vAJpPb/GPk59QHKyPFixmNx45x5tlkxqtgScuI4LCJcJN/XL0Kx2rGT71QeHD
TTCtGYXRuyL+iuRSPDySfPy6JbDQ8VTi6nAyET74mPLWmFj/gLVLwlxL6m5V4jbceYFoKOdBtjXx
Ph6G79lqkGSxeRt9+6kurDrlITb5CE4LPgl6Nzz3NxAm0xMnPOXj9u66GYwNCqVI0mZSHlGJtrvk
theHQFDY2ugqvI7O8CtAbuMIl4PXMIduyac88xJOIi+lWXTqAVZNiLvEpy29EE85YZNqVbY2mIf4
gKX18nv9It/b1eet4fSlxAvjpHpwTWb2Ke08Gx7AV+Br8pscqMDyJ+Ron/UIU9MmsVfZa5ImYYCQ
exhSP8BjCekEU3KFVE/A1IvSLhyCpUNBwmxOVjod6mnyUTPz4T3HFDjSO4ePuXiHgowcOzano3f4
LoIitQN36pq7xShsJRCtdnrN9Kri0fVLu2u2KLw0DbbdsS+q+wYvoz1dH7wHeoy58iX69FCt8tgv
eiOsdn6rkcTlPX8OPOtZGFoDsGlKh7Pk8AqZjjngKjUFXTaT6iIkfoo40Pj4VRY60mtCv0W1mJF4
k1515MlglFy4h/2yqzSLHQr8a5UqBmmd0XrXWlMm6zQ6ib9LkaCu0GCqnthH9j0sHmJUSD4CwHhV
vqagbJFNIQKkSDv963mbpk/vu2HO+F/jqzJjtvwtw5DDH9lmH5Xrdupk40Qwbg61PRxOz1UbC2rI
6HDC7RTKreQKVaPyZpS81UfixeUu3amAeyQB8rk0KzDJpW9woOcpbYntMv505W/a1bgrXN6Pzt0m
mElH0T92ReDPfzIDy7h9pLJRwy1aHyg65sCdABDb4ys6PTODt1WFcAOMoeIC2Kv3xK79Y3RkVKRQ
32q3rE4Cir63A2fRXOpG7BfxRZ6CNpKMq12FkFztFYijZDnJsUZKyPSqWyN8y0n5QJgSN6ZElbKF
rkBNvP3cXSVJ9ZlsqP4zoBPz+gepL5Eudf8gUNH+EEItys+rECxqzPZA7DhpbfnTuyOrdMG0O3AL
OeKxmJcbSs9w8rzBUdYCs47hNTq6VoT8O+i4mfPqJ7NbH993tkkHiWSEbZfk3CNzFHInWAJLmFgk
BYIGDfbtAdL/Z7Rnf7ohk8gUaHby+nKS3/vPK8uywGFOuWMbx6s72Wi8lpmXNNwZ6AVbX8z/oHFk
Gz8jPYV/GEcEiFRRxmN7fa1cmas3hENJV4fbAUqBv/NfSWVScOHPYIjU7LwNLrRY+WQQPShO1hN0
b7cS7O6az8M+zEq4m7HQPxJW1MDd2XOgMtZ7LDJnpJjToBG5Xnp97MSvc971zEn7RFj8k94CT9qi
1kJa9UrgIZlEHCFVuwDCsOPVO1diBtl1RiEVZ2CjAw9aJA6jnRhmioDBFAIc2ygaJbx9m2Fcsw3r
PAzuukvbPE/D2DMQ94iY7/jjETDJ93RE6x6nvGItr4vm+QAs3rv/kcT2NkT3kSc6CailC8sJUcyy
oTLLvDW26ZcA79dBbYTT6RNe3lp9uO90k7fh6pBJgw4aj8ESg/1H+3xV2yZk1fiMzSLyb5wgHcKg
e+hF/CYGvt0Ef+L47+TxxLd/aID1fooCRcXqIMbksO2QMmuI1f4aQjKeGCKAa9xq5cZSetRM+pO+
dGBfJHAELaEArOLI/WDILKd/mTnED6NhDE9zdhld6YIZsUV5IH9cwrrKrngopiPb+Oz2SJ3uzwji
G1WHXq62J9s14dWZqCIC/zMvSiregD94uxiVbugCjtLuvffWOdh0QjCYQZh0DPaYwN+411lOfZ3K
NQTMU8cytcSbI6UzQsWdIp9MgfP553m1o6+I4byt+y4nkEftWVdXiAF0z2pfekqCo6l6axIJ1mCc
kpm1lC6VdUkmtbMR0rRqRcOVP91rvnxQxQkMGYJFU6t5PvOBPiGbVe1h45AEUoTHz+Bmgb6vPIqM
2HR5+PrBQzwz5J6yM0VjKMtYfOyxeiLGYXNSCK9jjsMeJy+IradQlEYGWi0I0snzA/R0e+euTjgv
BUurXPlVAuTeueXAennFAisA0QiAPc8WbAKJxf1cor25PK2fikt5SlXb1uYxoP3bEHdcP/xbWf1e
KI69cSY1wx3CvWeTJ367R63sDOfdM4gQ+uV4LB7/hnVuqLVSXTUXK3d3qkHAcOw+an74kco5wgKB
gUkLLJmbgkXNOesMEShnK0xyqIz3r5gcQv2s9NL0EZcNTxvbHzLgYcqh6n8TWNj2wc7MG5/qCdWo
JTCP6FMo7auSNKm0d/Ng+VGhBa4Kli2+0nCUeXUl4X8aFHvnFRUBlQ73nGjKuMl1y4DtZ0H6x08e
JH2YF1jOCSO88ofo06t4h/MZUFXxGFU5Cy+Gbxem42bPqRmLwhF+gwxkbLbwd44xsULf2oO1SKfw
3JPdZwmw3Vfx+BAnMfuzRNwPtmA3lB+/hqpq/xT51m4LKz0tY9/3Yl/kaIG+ig2MK7gVFORJCUem
n9/85BBpJatnjhj8anOeaJIvgNc047OrqKw+oGXdGH43Tpu1GqKlN8GBTMcjuC6upQr61ysfrhiW
kJCgfoIJeflN1ed11N/ZjyCinRrd0ldT89tGfztd5LzDMSgSK783QWBEyKMRcfGlBB0hFovKAEoS
fuVnqApnnZghYatJ3BZHEq7G7R4IF2xH5Q8CUXHDWyjjk/H3+ZHEcjJaexQ6w4MuFbu1cQBNht9/
lSvB6LTjlMp671XPdFkNwYExlkDXGXRnhtnmGmSMBBq36qMUs8ilNHqBDKlbD4fiGrTzrgI3zIC/
JNq6BmxFb7hTVo/l27smYET6ASqLRj4pT9c6/mNl119mZYHGKTAGJzF253h2hY4gwzPeEapcBUm/
SSjI003w50Jn8P8NM+sGwuBbWyrQaBoUpimGt1pPbOtS9DugooC59pfUYPj15CYN+xFs3X06uiqX
jFMuHnniaP6QVNQJX2ey3UYw81po+kuPEni/xrs1D4joiONxN1ptG2xcji3PbXKrfuS5+P12eZfU
6ED5UuHab6nzbeRAJopbwsaHpikgpnXckkiJJsEG3ZUmjA7aIMPta6USWRfPCtlgARlAdnyvSsNX
tGQ2BKYD0cuEyieHA7EVQv7w2nLd2rkk+Kf36AbhJaunrAp5vLdCBKNzB2NmzTBm25Psx5xqydze
yQuOay0nxhyTlrEphemgEdNTDT0daNZA+i/W4k4MfSu0gaosG+IjDqPeyln++1XgG2AIFPp4hCkd
nM6m0z9i2EIL6NJC0PWpfeK/JNFRhd+KYSAuTkjxYKuRBBpuZmqixDqS6eQkyU3Lm2TlK4fyWJYn
T8tb9lu5zlmKf1+6OSMyLnN8I5QoE32u1vzDe/+6uOmHIWL5z7nOQJRNwob271nIUknJWFZCRGKI
p0SDCi4klSo4P97joiUR0PYc2mXoV/YGd1TR6Mlq8s/CkvtVd+1/dqOZ5I9hkRfL0CymI2GQI1ZE
zhz+m1jZESNat5aNEogMHbLTb80Tkmmw/mXmjhQTpCKfppv+OXXRqxmuvyLeWJwv4lOlYioG0Ed7
8iN8ogwJOK2oN+PRuwidMPtKcOLUrNE0HL9xlivnw9P8ruyMBXfna1XhhiMVF2WG2l3TLYcCLVYr
Bgb38eLweK9l02sIiq8nDfcvu1IotA0ZH/BvmhYPvl9IUa+vzn4a3UOgeyTxkjyVTqpZja9qAvJI
2MUUYn/BVz1oyLvQhIfxUCtpt7VZBHUBokfAOZbLWHJbCPhXYoYdSGKbJBDaX/rpjG39FQu0/GO3
UgROFK8PZohG+SMkLdtWO/UYgq0bd6yn5GtB+Bjn0vUCzyerXFM9rPVB3P2XatiPEQX8/V99ffnh
GISo01BaCgDZuhbxdhSaXFKy+joAHBEAwbnHUdxevPSwutewAZ7MKt6JVDfF4FGga+V+wKiT9haB
nauEzhF8ycmVZK76mK8H44Iw32ehnbBP0V1TZBQI2+AzPikLmRmkLKTD9YkOsqI/QUdiefh9dvmr
Ks0dTGrhzPK4faC+DV4ox5MZNWZB9ifRXxtG9hOUIh9KrnI7HxoFR/6fD3i0Rngis0DuOrjsyoU/
74jwXs59P7BsgAGdXPG0ArNBXf79ebtFtBjYcL0UZCeiJ01gQLSDFY1RCnG0sNvJk/AkzeoBBrH0
lgFClBuHSFYrGMacQW4hxQqa4PnSKcZ6wynmmBBodOoFgmvTjT2N9hOfQW0OqzZLYNyv7zBpGAbE
i5eZV+KFTJKNR1u7P2qO9v6bZWf8kVAha3Xo4LLNSMSdEWjGxoZTK98zjvoFvAbnGA3655o00nGi
ZknACLD/03MxbcHXguwVtJkE+XSbpjzK60MFhvEHxPlzZdWMCCmAg0+10gO+pjleQbRd8TiBBQVt
kWJpfWjuriEvB0mBnA6NqkAlmw74FIeZ8tt0FYvBm2210iMMNjUKI5obFxl9g7cWU+Ga05rcW2Ef
0orwHw4gdFqpwRtXO1nKSzCezj3IBgTsdKGHv95K0Bk9mOumTTlRxBMp2lwRhBns2q4QhlUA5MZE
zIezeygJPWnBA3QgFVR3SQaYe1wiL5qAAFmfwucxoO1Zm2BAc7qV00pLpusirPrOvmK5r6HxZ3m8
1XRTBoyMau6xXlKbZsfv57IDL3f2O1GIqjCJRoVKGSSOZCA0KCYyLwVKuNzDr0EB5ok7H0gVrEpI
Fvgbyxqbu73T9CMCHBZrDpAdXgZ9ece9ECP9nL6tMce8tFcM3Vbr9t0VmvMCvnG2esCFvgE6Zmfv
/xrvRZKMq4aAWJH13w4WSwQYrXOSSShiP6ljyvvLt+XgpBl39lJ893kUv8eFie3MBl23S4XIEigj
SPMZFll3zRQMdqeUGtPHuGNhROePwf2Bv8pzeEQprFyiP0UAqM/iAgs2fhCTy+MDasG6OfsMda1B
6nNTnZ4rh0q8DUPFvfQLipxxi4QgPPDfntZKC455sXdl1TVzukUYlxaTx5p2xSXhVv0Uk5lQ5Swf
TIrnWEsGhCuDvETqc9BYzcRvOnQzPkvrgfsfU5O95rzonEvhXlTXUIBbWKGCEZzomt25nOW4WLJU
730nKslI1/FjOqbXIFxK5Vn2ZRavp9FZgPzMoCzpGKRSZH0PGnnohxfWsTsBWoDXWjwqCBoY5ZF9
nrpK6Llb2LI2fPk3VHadmo+KydVzJUGBEaTPHhgmPWI4V/wwZCMEMN17YpNCWv/uF8szKrglTKFH
VKyD501k18WFV86fCC5aCV/wZbgsw7xh7zXkl9uL5zgkmSafdQpH5DsqQ8qieQo6+xjjIos7lcB/
2KSMKlbxBvFQ1sV/rfxwGlnuFbqBXdEQRb/T8SzkUlLUK7a7kkKQ3Mn2DCd7q39cuwU+yoLq7ZH8
/7zhYt9hyzJvMyQeCaCi1qYHkB7WgF9k+9OL13jAY9AMfSoUZXfwChXg2rrGjcZ/w+fxRojbM0tR
JFIs3gXu05oX42dyhJIq9ygKSncW98Ghffs0Sfk4jgWBbIVhpAUz1n7RCEoCtL9najAE2TQFNPME
4iRIfSbwkHoMt8sm9W0VkVONwLwEO8A7CbdjtOXx37kqZCt5YtLYuQZ1JyFLNE6Z6UE6ISwwGQVo
N/FiY6jop5Q4jBN3ntf0tCSN8OaxXHHA8XgSfmL/NhCwhAZYw3lVVm78Sm3JzD2fz3piXe8qjhgX
7ZF4xD0x6kDe4tv1mA4l6DjuHyyVYTvl8UlEcr00wOg5kyeZMUT8Wkph0rh1Mkhw85KDvFxT0rr7
8boCYGPqQWN1mh/FHBO0QcXJNF/pp/GvySU+rWj3nAO9kxSuzmCZr2renFNcr7lnXSpjYD1KiRy7
OXNk2oL0LcgL4dNnDawA3T6c9ts5A17EvKmU6B5Jhs6XWN2Q3u4khH/zbAcCsna6/A+ijstyVv/I
VpUNN7Fs404FPsA9F1c3HckROMgylcWKnlCTlPUCG7GrmKZcnHFrfeps3VV21y1XD3T3OdmKeoAU
97nccS6eEx92DvXFTE800PKQR5jvJIuFrlKPaFTvPKXdHO+wesrBwJg597ARKGkDLZ4ZcT68iFp8
5pyg7VUlj1sIjes9+GDhtMNFCLJze5Xgt7RQG51j3r/7bGyx2azfw1lIzp9o6hefVCyU1ffAdk/f
lKYy4EOTgpBUk1MB9ucE4Bu5YrCNgRFJLvcOpp3F6Ps9bsMNB4w558nvGollGNdhrm45YMMDW9Cx
FKNq7wuVyINoPW3eVIdrPelFOxRTI75zU6DMltuUY4kQ+VSa3prRIPE0+v8fZ46Bl4FUeYryLQtD
NTUdv9YOUaZtbd7k+0r3i/PxkV3SxgSvwchd0JnI8uPTY4jrRQl0hw6svc31QRYP5yPRQwCIjve+
EFcxGvbk0s5ogrEw7OoEq8ra/ahHIQyzN9o7vGk85iEK3ZKSwqqkPXx7tp9lG7/csShsRmhsKhHv
GewxjWwQPLmyOucUdiiDDDiWlkNaS0LdZSC5DRUsgJMjy9Lanaj8Tmup6sl4g/JFyKJTa9eVSVDJ
+Iqb6d7CkA91iYPPSuXt2sHOdO8OddvoM+6QDy1po2JxM0a7uKdNLAYyz+SYLLehaPJ8o2OB90iF
d7KBaJsNyEILFwYLxJgKKNNSa/t2cvOpLfcste2NKzFyBax0UDrJILTvrrt/aSSIEdxn9Klgz5Vn
RTsAuG2aiaSA07hConKnvno5gZ4ryGZV2W8ZC/srwBjNJXK9TJNT67kgXkkdDM2/KJKlaz+XQZyS
4W51LyBJh9k7uEk5JnskQAelRJslmp1VrOTTZouagIF7bQrtIoa2SiFzl+6zGfF67LHb4xR7Gdbz
jN6aNLWl5nmf++23Cx69lG5vVAV/g+Y1Xk5QcDDTtEOdk0qyo1f5MaSekIJer1f8oEz7FMYuN7TW
4gqZyJjEOrAcWAhPmMZRBHP1eu3Fd6aIWgWuwd6IO7nng2XNYVZHATwTUfUxXqmcAOD0JZUQgGQz
MqVzuEDKn1ldgV6O/Jvo5FyP22ca7xvaHylnxrwF6i23NHxhYtRkTFJn6H73F3wTZdCvyOV7L5SV
hTDAkOx6rMbDOxlt8GMEBiKcda+nwQI9nYg3R1UJ7kLZqO8ouNNlQGwQF3vv/zCHoyUsMb65+AI5
/CLcmwJ4pEx6eH8Cs93OiClneSQDLkzsTEqa/RpDMl7HzsrXvOPgDcnuWwE96gyOy2EV836urdTm
EcKzhEWXwjhfCHJWTM/e9LHeLiW424vS9h116x3ks4P+Hk7Mf7dNNS98KaM6MjYTUkaNvfCtgsxh
7AeGzx+UZ/31MMWHXycBP2fV/IupkypTeg3JAnVqhwXFe+XRavDIzauCrynhhjTZ2ImKt55HAI6+
ZOI9jHMeYdrpcLoe6ue7qqIFrUCWLOAFfTVTY68T74mBg/RWM2HTyxg/+E+0AT4yeLfw4tgFDHvO
wxqddQ76wpvL36nLtZ89pFO5rhg+yuwLmkCOiRGQbg0+MDUWsmNdGyDxNJATOYT6HSFkV2uuZ4ES
H6/bfS7siFQyAyL+dK8rJNq5BNYFvWMNWfFUOTJE0+GjybkeIZp22kR/YOPXmjge4sWzF3iyhH7I
2hvtab6/uFSIxADO/7H+/hEnSbngdYDU3LXtlrLcqwYv+0BWRrkTnwkd+LY7Dtqr/iQbGZMKzIW3
mzavZazxnadhEY6E98gYUGo3m6XqhrqH+kMXJ1tUC0DJDMTak4H9tjgBj4s3kU6NgZtMgMmZp/XI
cfUiCRGK+N0tPba7ibCYCFOLmzyuBHOTO/f5d7RmsNjl35Lcnfo7wI4bAluGoR4G4Tz2nU+v7FIs
x6l9G5VckVHgHYVj2mdz/R3uLyZsATc/JxIExm0PiZshf+wAA0YGHCXYuYA1kAcUrR3uVajCum2y
PcOXmLmswfL59pV47aZzOtmG8ZQj1zW+SyzbTlK7r3ydSd1ziz0nmIAYj2eWsB3WRKTLyZInx+Xo
BNuk85sHIWuHv+jUtwy/iJa+1rt8h+GSEamNfNPDzX56t8yJai/QRkJ7rftnCFEuxW61tkOcIhDl
thKCN/hqguP0Upkum/oNAi6sKWiuw78azAAjLNWb2NBpWqNSGjq428Z4AtEfz2v2EOW8hUwchLid
OjHcIX7vzUi9CUjCRjRVHcYbtMmtL/ZXFUcm8Of1qpArdBXBzuhCL24g9eXykyhipSu6jMvzwODe
MSAgjAfSZk/IGtGLO+xoyrnUiRSPbO8XRUJ7Y8lavX1KUItxbErG8BG1GM0ctmWvNGqRz0IxRAKu
0HbQ+HvvNTTa+sUh1elVB+a4OT5O7+/A0tyh0B/RTaVR2yU+AbFxhuF/SGJxQnhIGeb7vf1Ql7tO
q33zqli7RPU5urpV8UZj44J3KFlRiRRGwKVlvKMHG3zOTtfkwHn1kwQ/fiG7Ot9Gqwu+OW+i9xHy
fAsiOU8IvbgFrUtGAHTWUbMebdAOgvLo37OBdhVea+Dy9cERNXFkEa91SQiwqjlAoaHsB04i5sne
TBswPJqDVdwgqWYTXV13gsU8qDvmcZXJyVI285FW8eHU4SqBWSZ6izLNlJAO8Jjce0uB4TvnsNVH
tm9XlEIKyQ7ipkFmG1d8hWe7fcuCYWn9x+PgveXCjbD6R0Oi4SLfDsXMAajrS6AVgoZuhO/PS5gZ
fAdZ/0u8ZSWS3EK2OmYIngwpcL9D8aLRf0d6qijeXFM4x+SNkRwhTIFTKzgXsiLY+fIr1yZGTjdk
umCpU7nP2FkYI0wORkvQzZig7QZ1lNO+dAXMO/plZ7+diuQY762UGpw1nWa9iWgbqqWi+CQgmkhU
LgrvfqvVwwWL/a9hnngywBTS143aQrmVPyPrbUl4vL4DyJ2wAE240gM9F8P9stpCAcY9DzDSO+QH
RaQOsig/e8K7TExYyrRyB+Lapw0l9yRyn6vy7fsbnhPD/YDh9GISXn338nZmbDZ4BL7dG3D7OD6H
PVd1plrWZPG9Mn7+ljWSq/SXHKQd7mchTcgSc2qIm9goLlOB5bquepJxtir/mTl7uM1rOJ/XFBN6
vjvLZ1xuEDI4tkW6oaKyaXUaZnYfCzKk7pqKbNwA83onxalp2pq5/6VW0L3p1hkBtcWDT4029xhX
YmKxMirOjlXVlczPVyg3y9NbFjJRV9+HC3U04O6FYdpLuYSEhsSqvCf0ug0uq4DjuADgDqXFjxZl
lU45G/sVMbBkDdEqfjvpJwUWVX7II833shAAt4DFI2X4cSjui9G2KSnl7V/GnApYE41r8OYI7xrm
sItMTSnVojwXEnivFgV9xMZnJygWyX6O11sGkKPQTxL7b/3vP52CGrEiw55UM5yNH8IeiqnpfcnJ
MsP9PBwZKQC0aMKk10aFe2191NkMxUivX01g85KLMLaZZRF1WlUYDWvkT4Gggq6KxK3OvHh3t7MS
KiOctLwI5UpdC6DhdLPJpFJ5rFqefA3qpzflh8k20O1vpIrnTH/CTSfiMpnvQ6pUh75z5nA2p9l+
QWVESzbxABmYdHSztXmcwbpnhl37e10lM3UDgQHY4ElVzwaI0ydRazwaOd5U5UeReCUVqV2ip0G2
+EXRX06DWcV6CmWf3jCz404/RCwhUp2eQVAiEVwfMPdDS9gPfr64yarHENjYgIiwZ8tY22NwPr1K
r5PllHyyCbIMrF/Z7Ydm3zglTqEL4LipHo6oL6+pgRDCTC0LCPs54QKB4O/yups87uuKSSJeVQ4b
kJ90kA27JUcaECvfMSZIlB2Zlsldh9l5NlQBDOr4CPfY/+FP4FSKOfshtGroB771X0j4RiExgfb9
ZXr9GiI8dr4+wlg2B++0FpdtkSnfl92StNfRsDSN1Tzn0+gdwsLSsVkRIyw9VysOjNZupflK7V3J
2cT8aJimYp8DrhpxzdR9lTyBkheAUoaAwOOuHYUjdLZxdzNXM0NjpSYosmaEM5cnlM3v/5wg1gG3
EVEMjqeBEB3ejSv7Uj+tbEgCXphg/VluoUmOtSPwsl2BwGOupzmXhAdLR8EGDEoQoVDie58gLXLG
c+pfsWg0OuZfEs80lDyZON0lC5NNar14/WgsO0UXuESzVl6GrqGNBKxEpvKYrhn67CKS2uZvZPmc
1ezl5dGx8sLjezHGhn1s1/yueZHa1DGB1h22nx6HlNkJ2UGLKUA3L5RmjbAGjFZHtxYAsPIFV0Fy
8HwykGUn4Ud0h6knrm9sobIoycFhCvG8IpiWyXQbaxjjONg8axwBeqXS0m/37P/Qs7mGVgTMG2if
5LanOfcP/ugssE7Pk3P/VI4wU/GLmteAVxnnjdSOfXMlAKN0aKIMi9KP5/XC5F9t6aXO8qfyP+97
7Q07DOp+lKHh6d8CNlatxyzW/38GokJ9Lml0gcYy3iVq7okAS9qkrW7qKlkgz0sbFu7ODzBsjJcR
EPsdLvQdEfsT0sxDiCOfMjx5GcB2p4Vao9+8ZaU4QK3Hg7XfqX7eX13Pgv9fsbqRQRtftJ5fMB/H
zx1/N3aeZV6zloIURVGdC/iHIJxSMS3srpZwMMSqPHJG25VIyLXWUmI6UKhrBVF/Yc5mp11HFVea
K0CxnkcPl5q2mjRhtEacgJ95xCNsaKO0ZIOTRoasCoM00fOZOQ7X5ID33JjZFATModT4doGQmfjE
vSnxR1tWlaTftdhQeZ8/TBmzsUywuaEKG6VM8NRbW1jgpA6SPIqf2aEbvsjOKSWVBggRaJl28xqH
XrYQEUYCUvFCbQq0F/t/X+1ZQFv4ByRPHt2VJ62zz5fo7k4FSDKYmIKLYc4Er5lOH59Dhqk7x1Qp
C4JZMQV+8T6P5C4S3TrW99NCCFdW7KU0yowNy7FKyR0dAFRkdqmau5BdkUDuXBA+XWgG+RQdrcFp
qlJmdPLDQD8MO1zVvKNvEDuy7eNwyxoMiAdbxfyVe0b0iHqMHkCKzNOv8AtYFZvviks12h7YyFtI
V3PaSxqIejedsp93A/fOvRv/Nvem0E3kcRtsWgNO0B3LDsji/hiQFsk1PsMOWGpmbMPlyPRMMuj/
BlUUYk9GWMceZ2x7Qe7hAKyZEBV0HXaA6mBGCxD5/BAyf4R+AgcvD0J2HIDokSSo9DRQhiCBpQrO
CIY1vv6C9ZwvnaD0z4IzMX3yxLgn3l8XMTZ2Q7lQEKCg8/4p1M+1JgjxAuhK7sI3DvW+Zqctkxvg
aiiqtvbYdEQ//jzKobFJL7fQ2gakpwIdj10wJNsYXwWpEmsHY/z+5a+/R8GIX+IQ/0R78u/u7t5B
Tl066kLZWVCrRWdZ9TWaqbkXMzdpf3pN9NYFRzX6vIss2B0HspJLUH/+syrvHJ2m1G+kPmg4GPdg
uGQHH6u4zyGwxjzk4CRzOtDa9UeU1BzArpox+rPGiFN/+7iBOpSh+glH2Y0e1lZwAzShXjrt0Va9
8a7GOuHjHltInNGWar2bV3E1RU/prXFQzJEjx338eqa+VJNtWsAey7/vGmIQ0FxmuU1Y9wJWX0YZ
3Cm9QKpgEhWorbFQnBL0yEwrI40B9DUHBTh9r41Qk34WmMIPhZwlOylKdll/XfU3pJguVTdCVh7m
PXuPV6t4Woq6n34fkSMtKBwhdlG77GaMn/9RSQoGAkcgZtMyyr6SPHMbyt5s0llfAAEBjNblDddh
2R6360E0lnTEd/i25o/iQwqWW+XHN9po/wxzyQs5fq8ibp+oWKps/6U4YOy/ZIM1uvvtwK0tU/5w
kQ1mZFXISb4vTgWvKFli77NOHdE9f50UPpDTmg4bnNkOcb1Zt8JM4qGnr7xcobJn/88LYMi7vsEt
waGFoVwUaS6eBaKqOZ+IG6iOD7MeuMCDX2pTHZSOKrCazGl4uYz3iLjDVir8sW2DVpIlkIoDYtoF
Jn0ZGC/x0SeYifUleMiNBXSGN+iOMMSrlvQR/n4vKF0lMtzeOM5y8wrhfbADYia1gh2rxJJmtUEU
ByfxKuHFxzDKeG34cgPow7i4MjCnbBURpI+pemfLrjXi3YJFLMVIF0Cf/dNtTfTBkxCkxX5ZqfNJ
4q8oP8CiR3ggVaEi8Q4QFAB+TaXpFkCeGhAnNYQIZzDL1RdqS8WGyR6Z6sKw74ysYpgQHM34NSK2
46kKmgRHQgNa3Yto32gIkWr2/9oxiHEBPo+X13Nqzg5AGtaLYjrwqEXdXUEk3ioVYY3GkBXeeqZ+
z/YVbtHXVsV8A3PiP1t4FEDuhY4BuRyx6smP8f/HrH/O1I6/KBm8+coVMZVvaydaiu9ek4LbV28x
4o0B+otbEb5MbtsFnIzcEOFK5dOfjZyBorR6xmoeZ2zhctQfJTu9bNrl0Iy7Rok1RLomxUVQtNgs
ZXhe5bVclOWyxi3CPc4TGB62UxHmxvbUMLZ2BWYiBSZydQTLpqtzvNmytN5QcTygOAq/CdCGMWSo
SYTk2UHKmkw/6yesUzao8ryGs7Zkz0rWElNM/CKeZE+X4BUHkI8jkv4d8GrMCo+zmpVUXUvB0t//
E7ojHrQ+ZA4WVfGPhoHAbCJ4fGzUSGHRfYjYONeySOow6rIVLlm782yMB3LQ9XjOVoHJ6BWDDsLD
A+03zA0QrD6PNbvn4FzwgGbyzxvCOPtXT9tW/dPba9yO+AQvCupSdHsCHxKr521tA2k+DdvkpWFo
dlz+5A2nJ8qwYhZwmUOzyLYszl85JHmGqb6hkyUEIpi50a1gvr1kRrlfwG3nuWSQPyertnIq5vhH
EIn/4xbF3eLbiV73FV0mWXpI80o4RMyWN+dm2/OJHxV4n6sfc2LKs30tbbb63kGaUX8ue3Hv22nE
UZJXGzIWn+5SrvhM/0Eb06I9MZkMg4J4PYXXGuEn7AYq4LaSGYYr+fRs1u2Uf6dsrZDxq6PGSV7k
kIcxJFRbI3icQMyK3hcs4yXT+WnQnWRn4cE3MOHvvx9d7L0+caAOpiG43A/fXyBVjH8D5V5LGJWS
GKG9nwGduG7Vp18lIHS117+xKuOZfWiKRcNvrrKmIF/fnaIXHpLvd5qLIN5nUtzJoyr1vjGYDWPI
M/xNKj72BW461ONDPpS2BFsjADs9Wwp7QSUQn6ur8x8KJQJTDoFns8WM/efO4+3+iJ9P5ei+7qHK
PLrlh5woRzRDxUg7fHNyQZVLXNYYykf48c7CbYKY6UoGkClPbFE8ZYYBd1IxT0Vc8FAAJNU0jSVh
odZjl2ayXfTE//GRtRSy/geJDEVwHzGtDZApNdjzyvZewOi4lwVAaVuwKsUosJ07RK7LKuLvhioM
W+qg90DSh/KVoRYzjouOKN6QNeg3Hxb68gFLS1uil/k+0IhGuQCg4/6YgL7W2ldWaXpgM9zO7fD/
X0dxF67d3Phwfs/uhwbp7k89KwfKwSIJxFdgBltD61lGjW+4LCHc1uxvJkv6iARoz5s6dcXcyEZg
n8QntPbMg82WyImw72v2fzubCmxMnJLzqpIswnlIDXc062sZqg0VrB8mFguPmqJhPf2cSjnW+KiD
3POY2rPB0fLciR8u7QCUR+iY2ESsfcPd3znquhRMPRMMsmHkZq2lCNIB4bX7YKh4wkSFESDiaTY3
PszR+pSzLXXpMfZE8b0gWaKPoarblISY5l7zStUXQiWux4P98gcvwnNtwk/4WJv/yeEv7maxmNDj
37pIqKKQdTrEQIIJhSxbTvIPpO41eneAG97I+eFum+KC/ZFM3Ya1kOqu3rZ9p1YTPFAdDnZr70ld
fDtnAtVacJ6ASwabO0gpNOllak9kLedJDmuiRLbrO7RPojbqBKTD/qjK80A1eF27WKw6b3RDhwm3
WGLArcCaLeoLYfDOyL6mYf3ZZKgTCmjdKpxvHdEE+suwXAaQFA/gL3Qg+0DZ7Q26Rg5ayjeHhjyZ
Rzbt3yFzIkKLxvrbWugKaCbo3GjxaMdaPxH+9REACEZ/VxOkjSmeWYUWJnIc/hqB2XI6rp9SCL0a
aBV367s+GIapiuupNGZTSxai0aQUFscmDCnGUw/J/m+dRL6WL0/PGG/ObAGmsSy61QY5u903Js/c
WZ2lRTvvszAIyz14PuW2i5Z8KtMFocSv1Pb7RaY4/HbLvFz99ZTiS2w0fOnXSVhH1H9AoOEMuSzn
HsMxVQZH8oi4vXimaAaMwfPcoGT0W5l5aRSsH9yZMUC8tbTYlcqYpyuas6t8FtA3w77SQ0JgTv/t
8E/H5skKsYttBwQxgiytj1I0sK3iMiW6YQDZNHCwqjo0kbSoHD9NC69QHhyGJcNiWhCXuL6SpQ+4
DrUNm8/wF5UVLFtAbI8EHfieQ3OEhVD8QNtLEp1ePdoyONIQl/KIeEJAN3+L8TeMdp8JnIpnf1bI
iCz5J4oLcJA+f+HKGcSJfq73UI1sD6cA5gUPIgpOg31YSBjYcvqyaFfnIFUkalM9xBGLLeY9jw66
5RS+mO0feOQtdNTq64Hwnjlp1VKNQTNpmWAZXJ8EFE4OIvkjwD89ypzUbZs4Z5JmNDUQwa1J34gJ
n+GFTAlUH3vm9qd4NncErhF7xjkKjkLww8k8sAwWnk3OCZEAZgOqeB5YJ1Qr2Z5amBGlN96qn/0E
OrcSOgGjH6B1Y9ilfIlsTx4CzXkUdW8N1x8kyP40GQQZoZqZ9IIP5Dj+tDJMkcvDxgPYVRFIcdrc
Q+tG7PImU2hCDCkVfsRDhrCA8g/XQ0gyYiRwU+C/dIkuvuQYJ3PAaTUcsxdsyxDvmBN7BqPCHC4l
7m13UHFxMUniSUt+EuBmgxpAu/nP1bZAs1cnYMFo0NaXVRk9Lyk9mES50wuQPj2d4nY3kvGimM6z
5GmJLcAc3fhn9BQziHq+r7203doF+3kbIdTZaQ+9k0800UDo0UFh/mNtIPIb13yBHIE6oyIEDLZY
MNkNqgd3pKWFdLFjOzoXCmrkgQahg01MzYC1Vmm+AcThLHywwvpNSIPAI4kh4JobUzx1CHP0X0Dl
1XbNSqJXUH8PFwEzsuEWQYZCdF5bZ66wFOSaVJOcrpi3GNrkrGTkcciRRLDQLJ3pPM8hWW4+4Sz2
5pgRKx0sumtdjqdJ/myi1+JFB2TubuXuecFxceaw6acz/PsgV8fpN2jxCXxQvu9MZ0hTqNankCGB
vebimwquWya4rOeUxoQmNE/vqUyQ3rD9tXdh6Ky0HxGduoSO0+9Ha8nlKSXVB4j28orYF3btqDhx
un05PSH/SC++Zo+P9Lgo4XYJ6/mfuZHlSzTbALQO8HfX+xUL6DFN73jcLVSODlLKTfVu0vFO6lmx
ThKc7ymb+ip9UCwTLZuVTtdTe8U9Z45CoqMvUl0UD4YExtozfQPfuHqZVax3iU5nxw+ZTut2xBNM
NBOMdCPQF9XoSFza2fz4SUWeWJzZQ3Az9GCgz1IpgRNB7bHndlQkayY5bPN3q3u9iWyqtHyGzEh2
HJDxfkHzBhnuqcfwDPwOj9Sv8Sd03jQztWcdrgIRPHa4ZyNNi/X8Yih1gsPSEeNcVS+K03u4H6ee
sNayBks8i4FuTYjteXwIz2vljdSciqBt+gBbv5UQgvllPRQt2QW5U40SXF0dajmCHAUERTTJcckG
43lkzjZoGu2lq+00Wf7La3cB18CjeUyaesTG45baWT6J/Q8XDKfke0MpxUESzdhp/wSyOaNuhVq6
FSZCaM8kptGuU7UAkwOUdykg34Uet86qzHu8bJFBgkcaZSSyCueJ74oQDpN0ZcIumbHaKlTSzQwG
VFrRPdq146x+cCH1ZEGOMB3+CU7P4W7iYtDRrIpYkt8PNCBtvI2Id8yfkeXi2Q7co7l+O1QtOaMm
pHmiQXADOp2kmYy1Ghk+Ib/KNNEVm85XRZhzWr79AniW8P7gVKKCEgIwRJjGFXZSTR9md06tg5NY
XPaA5Kil9t7E9pEMmg8BUVxWZn2A2lrOb3Oy1Oap6z+0gTiiwZ6wErIxb3DB4Y5fVw3hS+3g46qe
BOvctFrNNEbhuEGsj56jBy5wa3s4ip6AEjlHkwQ6hawaFJaKHjzqF2EcI76BR+ZqE1aKeTucrQx8
n7QxCrvOLAyIJiArHbf0yLFojhVUFxt5Kf2gTNQlx4sTK0+d1h1CAgYHaCFh5fklPr4be46b59mz
3W7h9ycARHzT5hbjuZBoO2vUh8JQVZj71WmgmBE7OQQX+4vs/w+/WmAOqh+l4+j/ajr65gvZVF+k
4CYrokHzEX2yjBN8X4sfW1ibbJz7tOmk4fIHWh+o5HRUkEVsLZSTzAyiky+TilWPqZhzNRjgm9SK
jXZjndyhvALIiOc0haW5gjTqOhdjl9Li22KTx8lA/nNkA+ol0KUSzYIkBm324AHqsBLrsP1A8XpA
RFQoF8KgxvPqUe+TWJurMuA0WCUNKrgPPRZkzyfrPMiiD5ffqYAXU0Es2Wca5sXKyfCPrwfkeoHw
cU+DoE1YgnC8bNFikyH+8EA4k3+34UOM7vkeS7P9sm5s26MyfenxVLlYV4aVFmtb2oxRu9ncff/P
z/Ty/AlB2RY7HD/Ned5+ozW1SSHkHMZH3NVVdp6cYRmwbtM7krpOo8uaEGLp2h8D9mBGq3PFVVKw
KGwys3NIDGITCv8JLIWbuI8ZtFU2ptZhfbd76HvI9WKRNsACOrHeMgZUDLjoKgK2hATtLczTc7uO
IxVwHUPZMBOXkx01wNYEHrq+DMl1WLnN/fopRALBOebHsnpQ2mvk0K+7LLkyyxDnONs+xDN9KN6B
swzGU1YQprLd/pCQzTAD356W6oeIUZv93s7crtaVUyjXieHFZ4p9PwqwFGspPRmglsAmPxCb9bUL
9iROsjM8k5gEOqLnpG5I1H5KN2/m661sqGdYpy5m+1w1Us4DBi20Cou4Q4495MO/CgmI7O5z4mJO
knb/8fjx2gOIAMT6OgCYI4CLJUTVUUlRfRzIQCGovbLdd9SXQErxiRFoBVZUmoeFggEuorRUwsNb
HYurby2OnhPFx/sMJHWgGncuYWnmUPVytSKQgvLwhVnk10mTY9J6iZPCgYmbV2PKmfQS+tyCb7en
2G9Brg4SoUZtGNeNrgdDmfZyXD2HAxy7FTIYcKswkj0K63hGbHLh2yPYlimSJeRHCP2OkmsLYDD8
CDSqM+GIZO90fSDDwxhfwgBxyrv9D8G1OogpL8w+9e9MIWbYhXMbqwhCPlGnHrtFkmCOBZrmAyRg
ATkoe5KJkybxht1Uh+itaeYuSzs39Qi37sRqDLOREqUl85fHch2GQryWOQi9x2aOXIFOOskNiVmn
OBNujPzS3p8HMTdNEE6eXDBL6nNh5483jw3Qpq9HgJjL3zkj3k9+WuEjKfOFutwyfvqD67MHN39X
UeS0VgJ12+acTxPg3GOUmcs/3reXnLO8wTejqPAaRdc5WVmD71sekj3XL6ZPFn/IOa4Z7bejBCUn
NsiTiyHpUeNfewiZCRwsFPXbH5unBFS0UjsU+WKLFBUyMM4z9nynECwCVbGS+aEtEEjiVgwazb03
muKsQkPFcC6yq2MtAEH0SFwluUOVgOxmxmkq60Vcr1cxqnfZrkbHL6o/Ob14XbT/X4jsPcL8DgkI
fsfwUmjBFatmPeA0Z2ov0eyrK4Y0zIFcNe2yCtxMO/On9ZRYUaBVCXKrmauN/H0TfAdURsiqMp6X
F8gw9aapoK3sqa2gzNZFaNOpDevG6yzF4L6X3GX4+6Q8A5BNR2E10Z1OJlaE+fp/rGnfL4F4yTKW
0+oHoB/2uKJTQcit3R7B+k9QWiHpOk7bmN0tTjyy4geBXCAnxFjRKIVMzlbQz6xm2qxYCXwdPmCo
ZAG97EZrMyah3PhU/5QN3kdXwPC1VZJpDHOwm361mnFIAPNcFrAteC94tC5aSqUdGJxflphjs/sG
W2sEaf7EAgrkXTy28+FpCb4vcq6o9pvRjzSxgjPEaOsgAQSwPCOoCgjuViTBX0fkjaoTUSuzVgFk
y9zWkQqaB6THtzeTJuTRakeOS7IrQOa21odBElQ9s+6FvvALuq5SOwjvUET9V7Xz34lP1WzsJqzx
gln6IE8wADai8gRVIZc6neB7dhr0cJEf+Pn9YOHy3gx2WGHoGp1pu1NuWTctdND3EXHk0CS2W52d
Hwy3Z2Kkn6kQAq2Y/BvaJPa3Jc8cfeeu5YX43+caQTe7N/uRqltNYP+y/mJ/0VO62jzyc04ZOx6i
oV783LSoVVYDAyebFUjUKlmopckGocf9mqH858/03sJteDN2CNjAWWVSLOXE47kfzWgkU0CecE+T
b9o/FuMHkoKD71+Kgpqp+9G8HVq8cZIm+tsDNoxlVDzk5Y+djVDmdYljO9d6bUBYnijuM7Hma1MO
U9o66RrR2IjK93RkW2Gmxou4kY7vTUMFb+q5i2+g9kAtnqRCaoyG7ix/7NehaDiwBzNfSv/Bvn1S
fr0PzFzuZzeOTPISGjzCLe3jjKg7VBWpiU4ZJAcdp0VenQRnEW0bkxIfB9PJ3cXm2NBGCqNGUGFq
iwpp2gKr51hA80jy+j4Nd4dCpOW96FQyQbtjQtiSkc2Mr4qQ9LH8MERCwZaS9J/jdP0ppWthi0W/
XwkV7EHM+7+Dn5u4NjiuuC//ic0IJUOKsoTRnbHXkXDlDQ1/zW1dOOyiz43wlcO71CuHzohnIQGc
f2qPlL4n3ykqmx6Dl/npC6sGXzZVwtojKTzQ++F2mmHJ/cBaOTr7i6fDJH+8LBdPHvZ0XMdDW+JP
24vZ5LeIADjWADzOu7dH/78gRqdX9NPyCY8FXU5qMEMnVRmr4ecTMmVVM1P1bi/uQelQkpPG6JMP
0UN6w0oxsCkJipjiRHU2PXizO0sYTpCIdRC6tpsWCMAcDVeiyq/Yc+TBzblwfL+SBcR2vDN9HhSs
HDRIEPT3FrUc3oSCxWueVNFMSej1M0q/UIT3BhyuGc3DdhoRNQbfF7GZEL50pvgtHbQtCDbXrgnm
rGgXNcQ2o6uPOhSN9Zo+Ih0gUKizH0ROIOLkzSOXrrSssg2dgaVXtLhNzexO9tgBuP/sRX2x7Yvp
q6vOSJFCn/ldjrT9GalPIrAZr+Ovca6MKllpZlLjchOzLkSPajRPfkyuK+VKUKpkwWkdoVU0i6nl
EU6WPEawTBd2bPPlykWj4ixN7WIK6RJUC14dCiKUy9aYMzD94ymFhklwH8fRESkXpNykHXXyP0ui
WBwphTgMpwoMET4yKqU9uO3vf5tppcVpMYvis3fJvOnEC3o7dCOfOkqmlIaUCeOGZE8LPQR88CEx
On0T+RQu751ahqRaaMPhAMjUof00bDDdSaLHLbQvnIuiuxZX2EKztcLLL7lzG9eGKeoiKvpqInTo
EEG/aNVYLRqYPwkk2sE9uh4xkjU9LW8wZLxO/uBclVN0WsEyJM6ygtz0IfW4aPJmHEZCtHuHxREI
tk2pqAtNzkLG+GPKqRGHDZi3Jb0dbfLbE6jIPTBjv6+PyNf0jrJRcpWNVd606fyNFHbFfLOTGRXc
u+HFSRRDyBffGaZloIKffuPTAi0uHzsJDuQhAWkPJnKAH6wtRN1UbqFqA8X0vhMO2u9aRue5LQlX
VaQVec3zBIE1TCnoL1JI5ZZu8dTA0OFvfWMuQujQmlXp9Pt/sqC+SjMK8SmjK+42EnljQVanGFd1
cLzV0ux5nsfOoeFSN/DyF7pJJdsQjmMbPXWcuq3wm8fQTbL9aO/AKl/nQv82SHtuEowItcyeHxHm
4rX6enhPdD2mjoQqaM9lHDHbi/SbT1D9brZnVUNgb6LvRqheBghNH96b6E5bbBdg1xD4yZSftzF1
ALn4sa1sf9c/J3oft3MIkWdOa6YHByijP8OK+OE4AgGU5Lwj6sSuBXM+DmonyfJ80YaQj4ldVXLo
5KaZFnozjumV6qASGv1j51aczl13mdXuTWzxu+jqQm3uK/cD3qSlWM06MGfo5Gh63VoOo7pSY7uL
/tjCgmiNknm2pywLR3sh4huLgCdcQJQvhzSebEZ36RUOX7/30JmTU6MG82KxOHLCH0N3i/Ahf5ON
vWiiwB8rSLZP532tnHPAh5WaAIEV4abN0wHhSnA3LE+y15NtOZOU2IXzf7MzCtwAIBt8y8xy9qSi
JSHNGLDiDcUSlLAjGjYDi8Svs4K8V5H6dRBmk8rYwwY5B3nJxdGOGsGXnOg+KtAg2FcRZJow+5SZ
2/hXrwDP5CEJ5fma36a3JUTfTRMci7nTgWoYuPuiDgfmGd1NUI9K5YARf+cl8imiVH2C0lGO7NdT
AUQrAzg0FlcfyuiAWNkBytzVJ5Jg9qSqpuj9A2wiGZfm2Xy7+SEA5U/eJ7clDSG8dyIrix2ITm91
HEzFD+rtCk+F22rASz9MdO4uKsEgQkuvYDMwd7pXqslhiFWjaiG3ennxMCQTBgg1ccpo00HYD6V3
tmSI64qGmx9fepVdETJL77Q3fESQbO457Xl8PCDY//FdYHte9neXCZTT2KC1M76sM2XpdpHXDDi+
+cRJAoI2NiUIidCYBB5VhWv8HqkxeJG3YkBK2cKVMRX844RSKxT3UxFbjRMASojfgeVWfi5erXrP
w61fkeYpdWfeVRlwHRQYbsToEmGau/tJb8nfehG77hu3exwmDbAlIQgvsvBkMlwTh97q/bObIMHL
Z3ygVh+G/KBb7VdMau6WFY6JlBFB17R0WcMwyzsPoVb+tbHF9gM9MpXDncxIIjmNr/CnYRu17ynr
NRe0vMqHaiKJtFOx9dtFwcnBqsDjK9cVoNeezeGYxu/e7ScPJbFNH0xWBVJK8b5Qj0zV92cJWLeZ
IA6KPzKqhfkyHpPeFI5cmayvLZxHLeJcG1xKsEC5fkhh8pTtYehqyNq8RBamzE7YRhMrjUlZwLge
I6qcNK24dyfAXtn9PTX9r3k256oD638pXrt/3KqqIt7hR3vulLmN19y9WfcqhcFxOwmJ/fQVCizO
tr1bnSBjbaUrhf5T6hmIyRLjJIBWj92fbipWiZlBi8IjgRXaSKH1IEz60Mb3577MUIwCdSm6V4oe
NzQXhy+27j6Vtm3yQUjsM84WamvIQtMh1LrdBqWMp6gtmKA0q7B5nAvvyyhBXiQVBfRYkv/Cfl6B
uc9P10lorz1tL+aYEjsx5DaeSsLqRH+aARsZ1uoHiJ1Joo72AAdZFyByH5OYmld5ASOI/7SCCmYJ
DN3ud5BTLuyOe7vSNAFTX8GEn4eWZeWWpVzhD5uVBCDxxPlHdTCmJh/LXI/bZYy7hFVg7JfagnBO
7+nvsX+KTsDab3fMQELqEqdpG+FiridUz2K7MOQMctt27kRIzs0xcBwP1BuyFjRTXGVCc99dH8nD
dK3fCBV69PdUhFbprKdBKVkn1yn4h/QmA8iG6uprjcI/QYfLrkatTCf2n0VUOJB2kUUUqUL8U9S2
LZGXYAQMBRn0GqwaErYQqknxFLfbAPrzTuTotf/NpvsBk2z2zjGTdjhFGFX9G0X9Y+hrYZVZXEuA
nb7ix32mWBZKxcrBzuFIUD4mljCdZUmaPOdA0+7JQatdAjfS9yzXXCQdgenl+slMWKIWBHjeNa/a
U9mLYAKmavw1N4smKtIb/yDvVymKO4N0IZJTNEgLWvpHWQtWWlTfm3iI0q1Ew5cBTXvpjRGY8kPg
05hpT5bqN49sC1JWMLd/6EFnoXSUcy4FL4z1AtHuGkdMr/8tEnt/jQLBAK80vlSNxkodIwtJ1Zaf
FpzOOE4IUZSr7wYtkxQsbOWUYH20D0MolKJaX31C877z5FOgZbFbQG6+Kehhu9FJ8ySP/Azeqh1J
RW7dlA+z22m0Yrr9TnxpXPrafG/KtJ/cRVTu7wP+tOA4GeJ1qJoS6XjCmO8mwxqnpY90y9CaJly0
o/P51CKqfYWX+S0p84RgTpJi3eEE2+ItkRH2q4RYCGIixkPQb1jfr31aFrzt2Qlaot5suyJKVHCV
Ah2jXqMxiuv011APVsaFvC60S72LfNCEO4cr1NOfgjtyMqAFGSjgY3d26VVMErJUMdz56FrBm6G4
52BF230J0FUrGnwDwcgSpp0a9k3r4khwkex/qZjIH5rmIE8UFinroVZwte8bcGSva3ebY3k+575/
J6GQzwPm/GVB7vsIlZbi8StpHSyqeRy6x2kX9eftKsOwGpwwOcKmq8P9PzzBpWIx4iUcTJHYuKLZ
mlx7A6BxrpExHSsev/EAEz0MFvQGHmLvpxEkKC/PasnoCN3ccH6ewqqEPoE0+GpLH6tkie9JuEAl
CzyFZ3B9t95xX6lk8eOfugaviIoKF2FUC5AQFAL0COM61j9g8pWF5nfvGV39vjEmSMpZ8zoBGBKC
++GXeau5+bThXkXi010CG+9stKYZr23RRk3MO1W9KwM+/ubE7A2YPXF/opwM66/1tBJKOWD7HHPe
P4G7t0XGCld7znYfaBZsoNYn157kD5iPs7Suyd0EJtp6TCpuzKOytoXR5BiMzv9ZN7DarN7PXrZ7
Y8+j/BCCLYyrSlEfnt673VNPXoO5+Y0smajfr8h6On9urOXZ2eonRD6nnzx28BTKWhCuTwJCOZtz
N7DWuyOPGuj6ce0CfGueqJtMdE1lQCCqo/0UB/R1Kv0QezBsHpaln19aKCpwP/26CZii7APPrvM6
WDCUhUPVpVb1O27Kr70F05Iqh8qru9POuv8lPKjKSbo9Cg311IPpHUyhq8R29cR80AHsmqZcAU/O
v15lrtmee6MPI3P2cOR8t3XxmtrrIECqtmNVnYcnNP75x8JQUKOeTCMPJI/Gc9ZWN92xMI5s3A4u
9JxyosBKS2ieo3q5nRzqrcU/EmuRXTgNhgb3StYbXiGesa3JbZmaMqN/Vk3T5CrtiOzANN5d7ciQ
HpIqQTpRUNKi3exlXXk0cuXpzVAkN5y5AARrh4/N9tZspvx0NCVLL71vTCpZngRO8aWllL/t9gvE
zRtPxeXVUFJqDaLJlDsZSJLKDAYn6ALrEkvGVUzR+LvtgVNKv90ZxD6Bzyfsk4Wrm6NyIqFz4YjK
oNVsuCnVKNNzjTj1G5anlvE7zzP/bpqjipQs/rkUOSYdzOhadMEmdyyIhh8Z8Ydbe2avrFcKQHBQ
Zc1UDW9iAerdKt/9PIdNnpfTFKWhrfcJ6ewro/yPAhZEWZazjz1dXPjldRPAoiWFfl9cGa/fR+rf
ifpRbMSBdFkMC7DIlb0EhCN37QzQXsrazYr3me5HdBrWCWfZ72FD3Fl63zqQYoAWHvxOHwCwGLNp
+Nz7NunOzIAifCOqIbtp8+t5UoHOKWImG7h9kas28S+Menn2FoRGIGuRjLGZ3HCjGxhFqyg3ca5P
bFWlIfTdDSkftXfQ/vdAJfarbRzMz5axTiuAkcmsc8WoeG/t6PwGznJBJWN+jO+rY2ZFyCwNpV4p
Bq+qJZgDEJIcaCmSJjoXZ/mp5EnM7ASFExZuZgSDlTvo8D4ZCi7YVoxEnfY/tP5Jfz/0Cc+ZZ6Q+
HPw/PVhYknyPJDcE2aqnFpg/K5BGv+WacXfsk5ZHgLYzku3hsqs8R2CNF8Uo2Kd6Ciy2pVNe6fI0
eWmDW8gGBxQeaF33XpMoTZCTBEpSOT8UeUj4qtXMGboTjd7gwLUn2JuA5OGQZT2Pj9sP/Pq3L9Ok
gy+dCnutUc7fpqIVtnYyrXL3NOyosvzUkhd1xaWoBwCmHpsuZKtc/v/6WMUbruWNns5Jg9FWDFPS
/DKEAZW367umIAu6+Q4f4jnQBO9QwvDRRPVKNAo9pwhSxGNs1a6htrTofOq12WfTxFP+4Pa0XuQR
Zm0kG3e/qkVQG1LvoCcWlshB2aqBJ8kFibW+A0tLLKTl/maKwNvdry0qlfIUnQbGhZk5sVuIaQ9n
Dhem+g2Z79lqUjEtDnBJCYDnLr+XQsNu0/FQ69LqT4ybHm6Xw/WAF/m+FCff0Xbu7X9+xd8Cl44q
hI67qSf2wwFF3qkLzmBiSE3McTMGSlL8ku2Feqv7s31fYH0nZD/KiSb+J5B6e4sN3mJR3PQldy8l
BFWqHf+PEiRt5j5zzGMIXcN/MbzQbs5/o/vngkacWj0eXePd+4G9TE4WwlaYAyW3Bt3XjZM9LYW4
SpALLKuJhYVI9pPJJkZuwZZP7dKDAeyQUVZ08uP18ZS9lZMz1If0DDNvFyKCWpOjf4+oWDPr3nZb
qEPkqtah68nChVXjJmAPxmcW3MrO92nnwlVmvY5/m44jlQIHU6CXfstB7PZ6/iHM0zI3RixuLD8J
RA0fX8wVHaAxECQ3A5HOjgCAGphH50XY0Ybg4exF5q4Iliw5M6Z+ye8ND1wTZ2vHa2v8rjXeeT+X
kHa8RYEsSTxLFLdzbfIIqzgXu68h34em/GVSGNWOqQh5CUAcjnS4inz5wHlaPYV0tItjP2JS27Wa
HR0/GoICICMew4J8bfBdCjI6wZJFETpAq69p2cIQyPB/KKHPzmSsYovr4DxgnSX4bQK0oUiZgAc4
ay1KL1jTzntF2S9Xo1v7Q+Ih8jO3vpU3P9xl5oYArAMtZtGntlyINp/i5m2ZuNUmYSxLaj9WUsmY
uwDjPouRw/nxO6QU3uYYcsPujiJ2qYqJMOIAlfWr0k/IjDoJpijyBi4A/vt6Q3iOypi9gVvktu+5
Xg8001TEeNNnZNGcrCKRSvuNUWKNYC05wkEdcZ6nYbhKiFpPy2GmE8bXzobDyv7GmvDFLv/ZPMOt
n/dTDpQy/TINnnPc/mt5iwVtPmwm9+25lu3/NkVnDeZA0oYrTCggct6AC1I2++mYf7vPnrKXDJaD
W8MrXC+dgtrj2ZlZS3M1C06PJfgnbntDFLHeVrdVq0LYQnunbj/iQedF4g+m16LkCC+7OcLcgg/Q
NuzQtN1zwd7CgojkJgywWukCqvIqp7D9gV/mlGfpjQ03apd3sAMmUsUTWGQKUkQLHdEFb2JM9594
D72HAlmlQwRHfhdJNxP+N9P7uD8/p1qLs7zWPI5y6GAJ648B66ZrgXuKtAWhqidozU8kbteINITf
g9pGyFmlJnYYGO7zSXEMleUFQX6mFRwITfFfBBmtsQxgt4DPa3/MoteC/Fjkne4GUq2j1V/WcaJL
tzBilOdqCXqy+nyXlJkFA6af5r3HOk/YX39vFB30IrA2A9SfacDXTIozYMEgdbMx3mDBLqcetHq5
6qSlgEB9IYIwQ8v7/yZL5das7Sj/LHx2Qv00iYH54KNxkAG/Lzuc3Nplyfrd2qsCcnbQU/HHWOqj
Qal8DQwLUbzoaNh586RXoEltlgXvFTMRQS6R4QOVpbRrhHUECAfEfOZEYQuOB+DZys9388UeuTA6
JcSJzmhvc99F/QjFJJY8B0apwcC4aT7K8RDjl8TO9GOraywzMEIDN66bk72vpH+6f4aq8tQ9wa2T
lSlvEMv9acuXSWvmjR/FjIY9ee0tS+CtQfhSVJN2RmlTKMOiru/HDLoFWa0Bk/zgBeMd/c7ZXaFU
hIz6Leu6Uan1APdwkf/Lrswdr9X+LA8Vg2xrZhM3HG8KGlrpmrw2RgC1ZdQJT8t04pVfUE3p1MiB
WMq8IrB5ZyOGoOhpuKblbVsxf4VxXp+H91d1SS7SGnZQldB5GOqvgEy9eM8deBjsGSuViac3T+1R
4T2vkiXLDJr5c2vtiazX1UcH/QPv9P3pPWLK7odB7aw7OMMHTA7slKbQxr8lmmqXQHi4DWdPTiPX
LuwYVexu9BiPV8qBL+cb6Nbx+ikH3HwmsVso8PWzSBPOpfkVP0kxKtgFJj70K6mZFHWVXBJrBZCx
GTwGTJYR5mlqogF63/z+EP6gdRzMK77TpsScH5ThXHtA02UVboIfNr/3+JwXx2CcJBBccjSAfytm
7uqlTpAR+b4EE3arD6usgf6B0jHFhg3c5xWViLzcGf2o4PQusd0I55v1C1ABIzYikrQ2gdyCyduO
SAFRScIywyFc9OU+Mo3aEMY3gdcnvCXtHcY9zAXBfH0AcY88NwDHYAMyUXBh7qg5a8klzgBV4FS8
ZcdO1+2H37FLjsABFF0QNmeP3UfKCkaW+ba7H7SjJfqtUlW6rfRdfd8CaPiQF+L7A8nZIIOalrl9
sMR9k/5WztRXDhJxYA/UpJTMBpZWIR/TBQgBoVcHB+7hdZxKOc8fPFkdZvmpBh/27nOmr/pDaXpZ
INXA4/PeFVveeNhtNGYIlNSs6S8D4UBfEwdY3faYsz4iRTVDFerWBVbTuqyFAaIwfjldNaV2A+aM
R6oIiYZ0KOJervWrdXN1/ZDg8g0YFdhPOfdy2kAoavFpIxiLuU+/5TFbezMwUFz9pWn+3c2pogbr
RYsHPAzcXl/0+o5ub4Xjo206ZSwjrrY3v2O+YOm9/+gCUSQ7BpxEhUGySah4JRe4pTjYn9hJ+CUP
xjUq4lZhsckjfDp0oy6DXzMZknyydk5ATk28aS1m6aBkCBhiHCTQjB90yoLvdbAWbNNE7/6HiIW0
yZfs2KijrzisfJSK42LrgskY787s+W/yu8Mr5rdbkQwzFBdq9fD5UVfRFFvJRSnVYAX//StnoSfi
LwJBflKPphu8qKGx4FiZ4wbqgnh9/DCWp5AwJWesVdt27yPxAb9M3IMR2Y8scYRGZrdw/KDuKXaG
V6jYUJPigBbZmlpCaVnTvjlSJH8S145DbBZ14xHk4HoHfmPq1nWEDxopnIuRd/d/EFMzrh+LUo7l
D5KsGPfy34mdllXnioftYMQC3lA93LtInQN1wKV+aOqJmBbyyQL8QE1XJcbaLwkf1a6kS2quT1Hz
rOnHSOFwqiBSc6nxdbvatD6VXRyTCjc3+QqPh5gB8XPg55YtyW9WQLxiG/ZlsodHEyB8rgWN8NXE
mQC7m8UO5/VWK8pdmDAsnL6t4/aBkZeEsLEeaH9mpzLDh+B6IBmYGvQFCy868vpjr1ZtJ47jggS4
TV6I41TRwvNZWlFZcRopA/8tSFUEgaB2dg+JncGMVT9cLwvGeWH3brGOUCdrOzUELLLVFS0rP4JL
pcOAnCyBzFUniu+cKLJr+7aBrSMFXGJUjsk/4Ptws15YucBYbatoqD5u85ZqlZ0GPP4t7NkFic3W
JwAQ+VX64xBqcNgoJeGRSwkS++qE+MJmCTWF0VtH8GxKx2T5tu2yIQ7ZdZEpEnTbZOlCnmhlLkYW
x+z/i+W9rYEkJM/NMCLbr86nxf3OVRdddEgvsp6NgKc0vgxP+4CIhiaXwtH3mzBkEpryLRNI4n6T
GE3Bf9XzUbp0VYGt+XKzKsRoV4YVlMIeYtzkZo4zbt3v3L/Y7qEwRmWHAtle/k5cOa0XYW26hmqi
2+Qc93K9pzlaJ7O6SvhxJC/xoQkwzUjWW8B5jifnNGs5jor5ZcmJA9RhdZSwQHkKNIJHAQ5+KwkP
ydlZ5OsNdnFMavxWGLFAbmv3MCZLN6G0qnsi6C3q1WRTKbyU/Wwpd4Jr/wEx4cFKBM6R+YMEbS0U
UD2JV/zbVNJLMGycJxcaEyqw9a0ospdoOfAha8OjdugeSC3nPoU56xheoMvUdHgPW+W5B7mJLZ+c
kzTuzQdM4MpW0ecFOD0yHM49juv7oaFoDBKHNqm/IEuOgncVoGr9MWZH7L0/a2cOscB6R6TxGxH+
b1IB/oZSHebsNX6xQKjIxQ63N1sC3mleU9C5fZwy3P4ciWvZcZcmY4+cPPnKhgFHbij+d8/Xrgvf
MM7PRdYnwWax+37+dmVlHfQmJrmJGW5zjy23pXiP9x+4rUVgYsUaqQ9bTRx0zkQ/QQf1nlXbJhsY
01BWfboTPXuQIOWlTiI1cwxut5pq/c7ipAI9JOeuyo9/358YSA8SDe6ErYU9VtqOdwIV+gXg8smL
eCN9K1KoA9OvrY7WOn0KvtYr3C23oB0BaiNxx1lcsZVecZd5FsZE0eTYbWGNXvTgw765VN9+aUx6
wCdQq1yCaOCo9Rv1OdAoQpjFHtjIPiR7LYEfym5SYlTiEsiqYlrqzL1gH4Gr30/fsIs8yQYl04fv
8lQ7Hqr1AHy3oJrG5WDFt+eEPERodGtxKnmoBut9dvm5P2wv+zp4G4PJjgFrjDTRXHZrqhAo/eTm
3xOzqXP18HEXvMB3dO8lYbGo6lDt4KQeZI0AKRqlnO8+fuSwuEnmXeOHY1vcZMppgVw2FzcbyBhn
vGF+wyN18Gzmm9YiBuwzIEDjaHmJJwFtbj1rNPzTCHB7PLH39AFFvH3+ciy7a4j2K1bQn1OjV7+Q
m7lBb1d0Opg5XOIVPjn8qgR8jeHgxDH4sDXcbrxahnh9GolZ1szEN75bNY2UzPLD/AzmfkNEQMIj
FbjSkjLq5sjCHNnswHVYmOhttzWeIQuseADtW68/8OiA4LuiPEMdCd2EXsunK127rhu1j6iaJkjq
mFT1kyne6ttB1egvFnycy1iKdZjw3uPHsoLTp0geEZ952+vWCtSp78y3eCFaL9FPZ6H1t/JdMsRx
87eQzpqdHd741sHqXgUqc0OTS4nJ8oGKYFUnqynpRRfWRQvYD16r5stKpAuPayp7nJPndZIErB3N
P2wUtKzCar7+5N3cKUBQdi0EKSOM6Y4lMHSq7alTBYb3rn42igRkpJ+WALde1nVsJYY5kx3NgkBP
0RhMJV039R8SPubeHFNLys1ZlNJniuRAa8fjGRgtVPZoJhLYIPEKxKE8ivyqzVIrMl6CjVVRxir7
MxRRr0bCAG411zaEXTdecckCqABW76dLlBtKfDpXt3sLVmZCCXTCaUFlkDGdRsUuVSRWMYVsMvxh
JJGa8YbPV0CWYEprHevIHWYh5lNNDCL66AtkWYQ1REFIlOviIhztY2226wICqi9aiLHZb8NsqMv2
9Oc/JAC/1flX6CpCAAdytdPbw7Z17NTIxvLdpWR66l86Eek1Up6QL6RxGRzUw/SrWj0QXt0AIyGG
jaB1vQ1l0dCS/JoEFwmhPlsypM/l4fnUZmtmDbv7faQxsFSa3uB6N70JQYIXzG3kJIdTYpVszfAh
2/s5bzkbaVCUnHe3/QxTcqEQBhY+1sfTPFvpwEDBvLqGSU/zZODDC+vDLCIlrwbmqzmfm2LkqHDC
7aXtqNzqstoMKBouPaqJFgbDaluS5UWotd0Pv9p9wvC5siZMVlIRa2GRB4HSsNHln5mJTyBHJkE9
P++7FQWArxPlB7O0lInaAio+kqeanrsQlM6mEUPAD3btPWB+1M07ankCx4R0bGANBHw2hIy3j7wN
qijhisOUiIOObDebLgvapPW8eUEgtyTulPctUReIpCPYgRmEsg0fijcooAf+qwi+OJpIgKQJKlda
DmJdVbSTOD6FeOgbLHQYNaw0neSU7sFrr+luunkzrC/+6mJW1Jg7TLdYfTodFfETL8eJbtv3LKcR
fOJwooMPhbh6ISO06P/LAFQoz+yqfsDPggTEQFp7TchQVIyNXBv2Minh2xHamj3932x8YxNd4dbh
BsDz4o+XfIziBQ7lLslQL4Mo1jX/ng9XOYIGl7SnZSwSay57JZCSC5dM7Gj08SS1npwAmEqWQYFb
B83A4JxpoJAeLmu9JLVnSrLmp8blyNCecntzI+uDjY7fVD7S8UiMYbtF68M2POQVqTih7tDTSRu6
J0iDhHx5FOzUN+CWIDQh4jZiUcd+kPWlG15SFZvziUAwzYjx6QeuAS7XSnXI5eFNPhACEth65Pg4
56jEzACPefUd0TDM5N0HD65hRlVwiWogK0Av9kDET2CwLJ8kv9gXFxMrHSlsKr82QYiePgYvnkin
fDF8E0os6NYQ2wFoY1EEm0/EzRI7NlWV/oC/XKAGKfVGrE7um9N3NPTDDbgzvJZJrTdDUB7Cxn9F
e/cx78fY9LgBmkUkYj2vj3uM0VVgzC7HYF1vuZdZStmQyLwVThCAZbiqs5hTIUdbFJfD7qrDvb0u
bp+rpdgjR2kaG2nSQrSIYAsYEdi6XLGK+Vwfyl8e2dj+REOR6mF8A1uI9hRgcfM/g9rQ57XCuQKq
EbwJUoa15HYb4RZcvZFDkduS+5k2PjQv8nc8FwKLaAn1V9fjB5VXVaGOd+2Q0nOUz+tVDbHjl1lv
SyqLN6kNtH5H7XG60LN5h8JXpbWBo9/4r5bHFOylhKbCbQc+24B+UdMytrBPrBwSXtCGdNgVDItu
5Oc5p3iBIDfwAKKnWbMWl9nlplUplTtB5xWq6XDECfnqVOXiE7SE9X91Pt5ExgMt7hpNvDZNWBiX
3BlC1yvo82wr69QZZKIkyD84z4AbEK/XBSZw/f3PzdMwcBpqZ3MmfbfvCsvwEYo85Mr04r4qjfHZ
M7wbHmXPx7pXp6PevthnOPe2q8QB1W7X7tz5dhTLF7VRvW0Ge/byOiK/LyV26ECH7O6/8xYVlHKg
e0hmvagkFYhCC/YLCZrPx7v4gBdPu8bG83ilMq+CAXbRdnPM4E3EnSQlzfTA45WoXjqKBxWNaTTY
H5+WkIaOSSFXz9rlIfE+kBuRM7Ajq8XjmyT3uPP5wtFlFvkogDp+5cckAQNaEUj5B4JIzJqsbIjv
kj7KlnvOadHjfVblAHWqG4nU7wbkgXdTGN94+V4DGGb6tP36tCOGEKpq8nrAxYe+TCrUQ3S+Nu/w
DH9cNF7gDQAex4sihw1RxE6w9EKLcwYkAIuYqmpU4F8Wi4uoQdM18BceXN59randcqIng9XOYaTw
aF1jRgistu4Y2VYB2j/aZb7ABzF+NwZc7TLDXq+5I8W6eMtckYGJ3qhprS6eSkV1sppn6hF3lsLA
npBYaYGdSx8tQSplpRVYI54PemxhMV2y5crpzmdIKAtVXYXJdX7EnxIeGFbl0ezDsQlillJFVVtl
Loga2xEOU+uKD3qW24Sa7PaLOaA4LyCT7hrmBi3O2qEWbladmnJM9CAwYXL9YKqtFqZ+h8D4GNH1
/AEdcBNtzElckggaXOt955O8hVMr6ZxcvgH53rOQs7CE6knKsMRYWHzuJKkxHSZM4fEfEEFy40g4
UFIMexOKIPh+C375ZxnUBJzcipjo0xPWpn+/9QKJxO7MGEiVWZONcjS5pJ/d1sROAQlaQnkLp73z
OgI/DYIdaEtZtZDblkKkTOJZd2CGPu9xjmoezIRGjxnhkRy7G5jVXRa0lfax8BZQvThOleiW/q8k
YVNtW/f9G/qTfs2GRz4U22L4J0U+4D0RMNwnk3vr4N+dAXii/HobDAamYEbT/JZBsJvNqAkunpM1
W9Mr3vFgGOyIDohpb+6yPnBCQpXDV/F+MYIU5lIwzGrXGb8BkklKHO4yTF2sHwCu16Rw5LmtnmT1
XuMHmvHae8hFkrh/IR8U0RQ9Uv3Ph4n7XiC1xNU2j005MquakUa4aTEtlo6pmdxct6i8ZRtDTFyP
0TI6DNG7oT6vhLi/ZkUV4y7yD2uur71pi+FQNwB4K4bPqqLMD1dRrHFqYJCZhundu/XTbZ7YtYsS
sPSDK6z8bbUsYquv0Nd3RTcRCG48rcGwQZlgrI3iJ4IKniJXU36PPew/mxPhQuvFN1C5G1meYPsS
yZRonUvjDgGhaaTJPEB50WF+Qd+Hb9TfqOKqZ2oOeCRoWh2BI8wLJkgvp8vDJVzwjnY6vhRTp7Jt
HSupEroQD0v6rqt8GZ+15bknPLpRraMFbmW6mevYJjbUupOJDAB/YAJuZZTN8K2XPpi+uu5p6lZp
isl9+rOZejuGxakneTWWdQtrTIV9H3LPMBoEBhVYYi3/kcBbaQMKWHL5//JRY04++b3KXeNOISyH
H8TfGgowLD4TnR4/2Oa1zsZveeme+bnAt9AbkKym9S+5gKLbHOY6LaxxiB2PcdPlWCILIv6Z5o7y
msB1ka/+1gzRLk88Nw8H46zRpLga1RHkuIwNZ6pmM00iUrsRKTUqSh7pEFy9pj8WCuXN8u9LYW/B
fHBlV/4xZ20jFFmi/Sg1ppEYGMNDHBaKQyvXtYJyoYobjQDaFJw4ylR5DVVh6bLEc/SMKEHO6h07
Dd9OaG84sq+WsV3p3sZ7y340XJRVonl0MpqrjFV6NNfzM935xm+x9qFozqVW3RDIb+q+XQDeEHfr
j/jHFElUrWuiEBeehA3fXFkxKNheNkiWgDkql37DGXhOpqIXKqJ3ftLI2j7yscxRNDQUi/4V5PEx
Ew5QL/RtZtA6mUdoho7sOGH9zq1wzdvkMdLzMV9i4wtydOtigNIa2P3UVFLkzwtBppksMlvG7qfu
hxGLGNuHE6Xe1fHHx5jC6rz43SyvOKw4O9ArGbM4bpp/TlDMaxiyupdjCm7RGd+S7UNhEfTKM6su
afuFi6r5GPFzFjvtbvTYog8ZtdWhvt0QFhHEmjuazVvuik5Ve9FLCm+xL0TWUppS496niW5ZbfOd
jpSA9bjjb7ziw6bDFBtwlFjVXLUhdsLretjMWfkoTdyTxcnZRcIi04rm2t0UEjmQdYeWOnsPOq8Q
/ZYr7/6nTI15i1hkqEga5F0TUdqVq5SJ//GUwUfXAUdgFrfVYLhjCVqQ2JacnXFVZrosePvbprX2
jue3krITaG/p74JwPRAyI3Qq/9b4lxX32xktrZPvDA2iSUq3+j2Z3sJS62nAtUdgTzKa2ItVZfLZ
EP5eCSqojA1ohq0dMlladPKiO7psZwPXf8YEIDJH/hKIoT9uie83eF3Kdp91sy7GsZzVZ5mQj131
YbCIw7BjP1bwsvKvpVxYpaLo6f9RV4NuojSKscVX/wuIwHVSXqCnyg+n5U7nx8Uh0FKd1bAGcY9c
D0fm1CmMEkuv7vVdAZxUBMCKzdR9YwGnSvwGYBQzwW1YER1yqbrk8gOTwElNMYGPXLrwti3W+dW6
j37QrkSmtGKUFoxx/ZrCzG90py87ZCHMiPd6V14pCLmZsaAZwEHv189sFxWfvwbsR+zMDH3Ubnp5
W6HGBTJI32tZSxC1HL/1WzFvVeLAU5CMqlcxoJ3cRotNqg2gFmrKjVkIthHjmqtrER7um6XjAfgq
pN40Mhi45Ovhuhlx5lHEoUGeB5KH8K17NLHmHRIUi2aXh75ETSxj7tnPpX2FvEMfGChKs1Efb/sj
mgVKIkPECe7oquFXFfpvyPoxGpemfIOCXbU0lpG8T0n9LRNqXUvmtbA5yhaRlPNH/Lmd7DR11QcW
imrQlYkfzn0zfLmLBpcjgrbGxiJGPlz0C1Mn9oqxaNo4zMUTu6NXu9RJavlYPBEqVKu2E75Gw8nl
0cQU7YvympXL90IVBA8cbBt2g7VHxZSz2Flx9Is0xC5w940NrfHHArJiM6H8/2HhUOxctqrZXEiE
5Pn4swWwP54zj+z/u/TspX/Y4UiMXBRj+7F1W6ygebIVLC5P70H6F9TkFnEX6xi9ac02UomyaWsp
/MBJPD+7P/zSfGNrcjyUHQaBC0g7SpNoDYjwAyv6nQWs0TUfFO0JGVVnTd5PE1NXEqHxPkFmKC9a
Wy8apYHmzfnp+F3pLuMvpx8ahRUQhaP98HzDSy6rPGlvh4BUBYCudLdD3XAbR85mk71hARFPkqnl
aHMbGvBpWxiSh2VOhcuywOdhsPUyAo3Yd9JHN5dXClXbxBhGTmXihpOMfZTj/BQ4RyEePGN2Zj+0
hQYtKzBu36NjJDpL78rwYSJBo6aZiK9lSisjcsMqUwJpFNlhOOic+hUy4sDSlUa5V1uw6Cz3KMBw
+H8nejzVn57zm2j2MaA0gGbqmQtL89oVwcdRYfWVRIsGfQJeKHrXxOVszX5+vEy0NsOcTh9eQlHN
yBKetGRdJsQtHBjYOTQTM13NwotLksFyMLhBHLz/U9Mvz/5OyiqafRPaaTnkD2K01rVXHQDcRNUa
BWfiJy8af/zzsAMkCWVulyhP9bxNnFujtrRnP0g38LXY1RGOaanIJKytwJzPPXZZlGq3aB+a4xhL
qZFKm4MIP1O6Dt2RlxSI93sq3dvjo1CBNtRY5DkWh/pi3z1UfszNDGmcytvNax3scF6lwY0VknLe
qKr/8c/NRTkYl50m/l45sijCLQCHQC6Zs9efIGaO1d5KEMcI+2iWKA1P1pRzRY5m6JHthUqQoBjh
FofGC/DAocH29ITKP39cpV3ZMheF1OEOL8F94hVttvG95cQWxPH5UFOalM92fh4SYrFRSYRFAky5
9o7Ckl2QXt10TjMDdjY+C6hufwq25EAGkA80AVtts5UCvUDPp1RqO+pAAj3D6hgfRIlS6/RgvuUj
VBrYe3qnNQb+Bmdp1SE1dhpAVbAZH4cp8p2BjT7NNY9Dle5DECaSErNFSzp/xkAzzlZkRq+XDYho
AE8fb7at/D0X95EagVoaj5QSF2bQySH5kEYHYxvhsamf7x61llJRxb26Q+iLlRjo52ilVrhSYsGh
sszAYZ+jVsr7d/NoWfFPjPAq4H39NaigtRB5EL+v25PsX9hDEIvkiIaTj/9JwXfb99dc7eAU/N93
cJvJMP6CzjhyHg9wtDHpvDHmbAM7wCvxHel/hJNHKO8f86/IsLrPAwHKUUJLYkMAfOm6Hdz8MHss
CZJPYfGZVua1ka0fyT5Sy9Kp3HcPeEczbw93mSCWDsU4FdZr0tzTETUoer6Uu6Bz6U7ElB7FklgG
9PKN2r8Mhd8TfXbuBwvX6qINKkIUEt2X/F0HmvmKFGq7QTyQr/vFhJ3eQ0G5Q1z4ih4zbDRwVzul
ona4AmxmFj7DVA4AHAghWdu3LR9FoKV6fXoFIeyWGQCyZ1DgScZGUWv6j7Ig+hyn4acxQcJT6fbG
tvikaAfSrU011usMTxTAGqR8+jGotm4wiqUgdV5Iw1qZ0yj6n6C5J1YYqYLOGJDAhy3B5C02Ss+P
cAITosjE/W9n3EbIH3H/LQVh5fvI/dH0eMg891qGJLMVXdAJqekYcF81qd2niOP9IQdXs8544rPq
RB5gxh7lxKT3AEPfGwzogJA+T6K20Tctb8EyKANUgefqh7LM6ZRQbldOzUiFOmm4g7gKBn6KBtqQ
7DYP/oqQB+EfLk9AGvER2RHmb6+GSI8eykgLC/eBZ5kd6bX6MxCP9l0154dQksZHypa0tuPi2v8I
KyTYSbA1FHA7DyT9b13evGbxZUNIumpsPQiPRP+kIwJvJgpk70sdix2v2QE9dPsqzgNm42VbFGkz
6KWoQ/2Uvxf0xgJ9V5OrWObPhkfitDhiVRO+yw4ZX2xjlHgu5qfWcrxY945JvEsuncr08NCL6/H0
nRpbgKxdyKLCSFEkB7d2gzjqKjNOj0GKwh8G1tK1UwAWgicf+u5r3R9ue5wR//Xp0w6Oa+lXKH15
VvctBU8oAXCppA4UhzybceOn+Ya4qQxfpRJoIB40RuNpwUiGt+kbFWdOkRNkk/T1BbSWYBnQxQSe
OOjKMp+k2yXDHBAeaR0Nkc0+5HCtuB2FD7bPE8nCQiyINzv3a/G8+M3BtPpgjhpk8uuKvEHTPgCY
uC8Sb9gQOBMaLk0GWy5QcKpeyKRd8F/d2RfSCoEiOGSNRseyl10S1oBkOYL9uAUTSFRJNZSMe2gP
ui5UQFpYM8+Ix2ZTU01CmSYx1LLbikeBP0BWjXDegyTVbWMEmcFM6gLevrI6Cke6nS6GOKZAS/W1
l3VAMYxiw6Zx1Cz7sjc6+K7+dO2/mukR4sx8fwV6lUpnYggxlwZ6pfMPS7Rs693zxDSW9zS99mZc
RoCRGh2g6Ccl/iOgQadc41q34Y8nJ7tlCkYdCW9glca9VJEBQ9m1EYRnUo4EYELb0aPF4I3XFrZg
W++GA/bgPky/w44egmumHokpbK7AUz/P2beyffwB9zR/hgdYQl8TfsexzOS5W++pwbD5OJuz8K04
8IZqnhAxi4jebRJEJ2E5SoqgL8cGY7lvrbdKFyMLrBKAU67HL26l7aIUw0RVQGUOeYjWI47kWG2n
Kjy33qabE4rt5QCGNirw74PzVQ1fSjE1f9Z0bsiYZLmqTwd0+dnWxCOCgVDJ+/h0/FBfZkpAA4X8
kxT7N5xvuYKO8/+U9e3XXlIdx32yxrh30n+vID7DGMzTx5W78P2f8bcaonVuSS9a75tK2Bnqx3cs
NEQ4gK7TQHLpIvd1osDE7OWYIZ9AOdUl9rxqOLSD4owhLowVtiBsebb4qijGrVqPHWWnP+eR65mr
lmCC2lMzcgGJipeyI4NC4JEG9g2CREMMlPMyE2l8BI5MOm/LUvB1Q8QtSyJje16urZPmRcMDqRIH
DrKA8Is8vfom+VI+pr+hiSnfqXYQIow8fyig5SygWx2OCCen1RV2ZjX1bt+oreFC3mfvtWqx+1qa
xDIlexufCL6DMyu3mM/ckPLrsG+0vqLFEdEFcB+dzdmtsMGKZe5/SRPnnA5v5N1kObGDOKXW+FFj
gSopOpPaRQhZlA4v2DWWMQYK1DWDpH10jC/uVK0Ls855+HtGAnHLkFCThdRyaJWXkPbqVlzTr6vP
Fa12dzESFr/1fEJDyTCQnrte0xbRWYdR0zq3j101+eeevZYtLgR7InkLv1+uqZV7wbsa+z0E5KJi
7F1vhsYFrqClw1BmSC2xMKECWyq6ktZ5ZgnnbVTLy15+qA6COisVgIi4JB4jJKjWYRwwrkqBBAtb
n1Prd7f7MXMgw0QSzpxoknIjG4WaFb8DaRPz/m7fZc5vtA8AlelfBHBiBEXSAoP9dP8gOSOXIohb
b7BJqTZESupYd4G8XtW4WHIE5BfWZzwfv7A2/iYw+HYjmnmOrHZH+Pw9iu0QOM2sDKh2L3QpMCn8
9S8UPg5MIYcvkgPyPehzK7kAVaHoNCt4Fo/b2heqCrvd69pIHLBdpL8jWTQ1FAvf3BxOC2COycxT
CSf5P54e99w5iQRnPbg14yoEGqVGrQNqIy9LPduua41ustNp8dD7WB97VLCUb2cS44/arFWrRLj9
a1WtMmghQ1lGHJTyXtwgjjHKPVvzAafNu+6Ujxqaqxsn1FKc4k8PTtnHJv+9Gpv2uTbt5mZ3e3oW
Ip9FWadQ/Xppf/YXUR9WaVOAEenfXSpKJ9sGwcMUtdQGvtRRmObK89W3J8/jTDR+M2b6nfZBCm2O
X9f+3Ov1SvmJNUF7vrBLAMyNp2pgPf83jmUXatpWdBdZDx+Q2AQ/U5pP6LE6hBiWBiGESLG+Tk+U
czMdBDwAx5n4PhVhmDxTCpJ24Ew9YZn6hGjPoOJgIL4yNA0A4R1Yc3wfRMzbhlNHGoNy9vpY5yQO
MXcBcddaRNHDX6wocTikObrHYXWgX7No3ay3gVHQWLsY9BeJ0MTztlij4RhruIUMSfBdAVfHs82Q
bQ2+KO1pBuVzoi9rEIRGi+iPdkLvr433Csbr8Wsgi7xcWr7WlSC5MugLG2lnHUZx+Lbpsj5daflg
nruEbDSPQqhscgSnwwzUQAn3FTWgL6w+SHtifuDlgqKmB5Hu8gUaF02BfKPBM4NBOna58my1JX/N
aSVuiYIt8XLUtxXKCNymklKJEDxXWRNkfZ/1T6EtIdttOB3Ajl/S/pTTA8is7fkCgUX3Fo4SX8tG
7Faw3hG7BkgY1h8mivHgcCBgBRHcvWgwyixeF2p9bYWGlNQ+j8p2NBcNrGpURPveN6OP7IEIB0hV
KxiadanmPMAEPYsNiEr77xei0+ZzAzGokZ8KiPeln1GYvCtk7IR1Dxp8Jpwxe09+zLBod7Yia2A2
Bi5FNkEALd/vJqzJid1G4yrqYHbDfyzJ92ts4WyZr0lNWhfEJLCY5tztuQbycbfFjMznRD/GM4Kf
goFUwvoKMaMG9GM1+STB0dQcqp0MFq5c8FeN0IMKv8IKKthVVKMatmyblQuqzBqjgijSp8q6vdfa
6rwDZySj92PIXOR2NKU9PeQslpYtdtsA88+aUM+f1sqZnf/wGjhvkLjJl8rKZjF2hD9SgHGNlHV5
mEAzPDH7dzbtvzshF7nvAjsUnrPTdXH1+vxUMcMagPrMXW4CDtU26ThRm6yhMuvTNzj9YRr6F7yB
Pvv0Y3kul3G9TINxgEBqfpyGguaL8io4V1hSDFJ+7rCH5KXoOyA+48gZoOwX0DJxbFbRXimp3/hh
zGNwjcLDuc7mBuyTBxNdeJCMrYM1sZVIbcwYjal1cGzGpFvhJohklhcADY16vcYUxnkdar+1M0q1
4ZFYV0ExDoQTqotrhQvIrDBODfvzKiMNU8jNMTz/9qzfMwT6drOYPbpe7hca0RU4sghHXMn60H1G
8NuUXOj+DWn1Ujvu6sX3dG4oKzi/pRv91O6SgFELTmtTNTnqR9lrruAIykaFU0+sbM7kM5bh7FRY
n6Z6SMY/yBTgtbuz9OBLuyFkQDZURsGKW3TsCdO4U4nldSBIachFz42nvnUVKNoo4k0EdVrGemxc
JXN/tbt4SM7noo3XnffzpRFZCSPnYZA4xbqahCmYqQeIiaudWeE/Py73eD8pN8JGDp4X8a97RJ/K
a4k0R1vXJmHRFJSI4lxWI91jv5jhDjIIA/AjYxFT01TJ89MDth+GOhgf0mqgI46eqCneWii+w3XX
SCYKq89BvzGx+3T79hSZzyAe9vOM0CrB6TRXoy+xmVAeFHs3A/rnnf2qowd+ja3TXFkuk1FtLPUm
MSgKM0u8XLtqfy4Y5fK2gk7VmyAfYRMKD8EeWvCfeyZ6/MtTk9BFRVEm0gQMySarRvmDl/88gE+g
h/iWOYjAdVjlIzXzM11XDdu4vldDWW38i3TEBFVMfio+r5Ka0JeM0CJznHLU3QPHmyMqPPwDGkdB
ZOnR/pOrTTaTj4wcN44ezeeXkp7qIhpIoKTkzlFQ6IxfjToWjKIDVi2j8Lm8ebqPePWJ6Qr8d8OG
XVR1tgr7PXpUR4hKNY+PSHtY8UvLFzwCHd9AxTwIvTUeOo1rn9etJXeu04IjASWMQzdSqZTUbzfO
sYWincAB5FVOLmy5uTRWRNEq6KF41kadcuERq7bqYYlEoeI3iIa86Z0KFa/+GY3Tz4FW3NoZUg4n
mi74TBWos0D9tO8p9xC1yWYYO5O1LxyYwTDS+7S1UHOl+Xa9oKlp8Z6UtOCp96ni5VR4WD2nl8nc
BlohqK/GdywJm7NV4GN9ucNbXS1Cbb2/OGO6g2VtNZjjPqjZZmBgi1TX/S01gpFETBadQTDb1USt
JsMNW1SPD4/k/OBz0i0SYXG6NgSjAHLB3UmwOvDaJ1cUT8aKKEQcUq4duV78KshzRxTG+lySEMB1
wBlB9qPqQQ9gMEsTHAx6rGtt2NVtoZhP74HZL+/hLdqfHUHqJfqMBH3y20E5iWH2ReDVGTkg1wgB
tnsgzTskxt7ahqujGHoJKRoMWJvZ6DK83+B+8NQvS41nO6r/dtUAAlxKzhYqaoa8QVRSoLH8Xh6A
H7qYcTXh9zf6AEt14od0x/uLQSBQV0FRCEbPksiVfKCJYu05ZPhwyhWthvVF3znCUm3Q81gwTvwc
8zgvFnYA29oHhTA8TfZNl/X+Rb7qaD4PuqD1gf+f50pd678eN1+YtutqxRqoYjPVXjNcGtvvFP4e
GqKhzvdPasNRdgSj4KN0xXNd8URc/6rae4mtEOPFDsSgUMdOvT4Lx5cin/la1bBmGStz/zexXdLG
mAs1oIc0p2y7KL7LZtmOnA93rxjieJ2orU7gGtKkX0E91jQ7TyvHFbvGD0L0EYB9evyMwOB9wUP6
dHCaQesMxM2MqBY3q6Lt+j+M+Srac7fQFUe/F0Z566hrGbkruyO6J4yEb3Kk5Ox95lj1S2UDV2r6
MjqIERCSoZWayN5RHp1Ulp0VV+5uGOBxlQdLxlOWkIzRAM1TfCRQxjcJEycM7WaGlTBOPvNOgc/k
m+H1rGEf0hTwai7f69MpLv9autaBE2ktzgWhSBm/0IMVxShY8L+ukZ6x/d6ddsX3DRKbxQjBY6/7
ehGMhEpzLZ+tpTABXzyd9n+6wqMtBL1RJimi/yLF+1FmOgQ9RD1x7zv8QorMapauR7Y+Vx8ePL89
WZd3wSrIzcZ5jmORvxZckAX8wcgKnU8tqvnu1kp20ifIRIp3wXhsuwjAyMidYW0646ug0vnxLgNL
gjvLRwafOKhgWfkm+ynvSg4BztbAuBMQ97uu1SwwftJb1B2Mssq+H7Rgh4sX0ZKukVzF8+mTh4QU
QuI5C1f+UQBaDnhUY6/+oxUYDPkSD6YpQnUUU4/s/08/7inZfi5EE+e9IngmX6oI3Bl4ZX8ORxKj
y+y0zeDKFSwuZXiYq3L6V3MhDrjpuSCR20iaxeKg+l+M7WtDzigouoIaf7a2eqGnBzaUuMHMpERz
LQHryAejemgyPX7TRyF/Hdk7rvGFweyWPZ9u8HBa0jBj+EdIr7quGZXnO0Wyf2yDvTRHReNNDigG
S56kNfvIezI9fUV6l30cg8cnG8Z4k2nRhElDYWPioaw70hruDPIZZSUQ1XZnMoRhDrz+DTxHznbR
1m4DrnoYHjgiRCMm+gIuCCrNAR9XPZo6fnPLzj1B/9W/7ZdK448aKvZPcglfffVtUHJm7MecUSdx
7ocW8IYd96Yq43k5tt4N1bM0wEYYgAKp5kGH20YEPspbuqNglovEIwgIKSfimoMro2oT+NfYX4Sz
g0gPD9wChj0HGF+SstrfHDqDyhQA6bpQxyLwe4v0Yj9Oc75GiBwU6Ku81is1v3QiTxkKKmE88nTR
78B4yKpF54+hiWmrQa3EmLzNokbCOYH9VCK3BJkLuDHD0yQB+XskG4+EW8kgt7q5UGQdzVyddyf0
ivTNXBkiooUiG+ZkQbHxdZcKWf/FYy0DhdBxx7y+/cz5aaSXRjYzFJJXCBF8BYo/om7DHAWbh6Ut
YyuES+kIxwifcam6YdB2HIcTYjbg6borrlV0RTbS0NFVSaDhJyOWm0pCmXjeNLjGQTCTEuXtFXyR
Rb4t4fGGFLeL0VToMZxBBmgvBZyN0/d9e3lepJN9ixBEwOV052O4ffF/XRD7TtLp+XSHVoSiUYzI
iLDKvAj7IJo9q18zva/rxS8A6OzSHGZFXUfQZ/ZKzIRj0sydryLNA0wbdwXvJyOTkgJrAvwRfkk7
uvjXymLluaW5LC7lqInb1u4ckzgu44mKDGWnEwV65V508ctiAOMgRF5FBdVHJMKR+fYkwSixqTbj
22l2tL7vsIZYHNeGqpl3807B9Xzm2OSP7Nm2/NtxQpPH7f/H1erA1PcSKJVNi0lBMHBHrwjcrhAu
Aq4XMTvVAacc69paGYezFrplqDa9Xi0a81OGZy3pX3Y8tmmKBW/BZoPzoAqW22G2fp+DNdPGxkkh
VdR5PXMdReJ8gVSLnTqvxT7uYaM0CwqDga44HoPdjEYnz6/ZM0y1mPVpwPhIEMwMAcckCrdXEX2M
Gk+zpTNBWQ3H89h/20s3oDcDuRrs6yFbceXL5LMvKJ9qnHZU84KclSsInoYuTJU3XI4t2HVPqgT/
ApUW104riJQe5B/EcH6JnITojr4ohZB+n6ChpylrSE0zy1y4WRA7aisxB1cObT6VQA2ZWWNoGdD0
k0kOh5iydfSAqPZt+thEL6Y6plNxuX/maCCTUt+flecM4WVE0/gP8GR6x023PTTkFanum4wCvcV2
egCYWzkM2GIikUxxlqUjwvg/P6LomC93lfazJXskgw/vI3O9oHP1DqeWKG0xPR9aCqxYNfqczbux
h3LJFzv7LgsM3ugibkI8BuEUc26hiQwx9ONrsK2wHwMlpAAuPKAJUmVjEkZCGy6aRs6fh9fENuvl
lFE66sKP88SLng5Ht/BucZQJUeosvWiEnl02yCXO3TMsJjWjZG95zpHd//n564Ks1ZLHusSFIDzH
e7Qf2bSjllTvYs/ZTmmFRzkEBQGWWVEhf9P+77TRSkId6E8D3cHppNiy4MEUXFtR2ogjkPfz+ZS5
6dXhsSNtaEYT5FiMeUexUozRu4MrNQ0/DJbT77hFM7KO5BsYmdd4sgcGY0wCU69Nrp8i8RJzIoOa
4OgjjYbycM4l832Rv+MUZXTJPCd0j1nI+sWbdgenRwtSlvuHtEUrDMvwLBNFwtSbwS9w8eu9EBav
pndgRYbPTwJj1Tf1sarNsSDruEjW9p0iXM/NsV/DV1yZm838dMPk3boxDPr7futFenS3ob5/UAG9
HO/xgFCRNkU232sbbFYzCiC2pX8nrBDZ1beBbHaaYiay8PuIHuuonwuGUzj8DazV0aVvlGQ/aSvl
ymZWaqZpzK7/mveHWfQr7xvZcJ3iGMD+RE8NcxNHihdQ3Uv69Jyp8So4JZGQJl1kjOGCCUpuR6In
qDy/OkhtK8fIive2E5QvftJcFJ8tFHO+TiPalIx7/0zZ5KOA040v/hAmBKsR+sbQ1x+A0PmLESUP
vjafNBvoHTxi8bdrJ2k7naTuLcYlpsjOUgmWBnf+X38uksCqVeynlYdXoSA0wgNtqUsQ1HhOlfQ5
sfXWcL0zfiniY4kC1S7mVfcc7bOGsiBZh3TQXwU2VfB91uodyz6aKo/chtx60IRiDaCWA29pEOZ4
VhRxyu3uD43COqvAzm9ufdwsqZ64/TSI0glDjeSz4GixRsIA2dTsRtml2yZNWj5ToRYWHo+wc78p
osj//QHz0UtL7whEhjxHqwICTv+Bs7BnYrD7WxGqcErcjJZT3VAoxc89Ak255VmGUmdv+3VWkHgs
jgQDNsdUmF2ry6kMLY8FcmauHfHJR/ueQV+elu+Igaa2sikkBPCMRgvGqS6SQvh9R8TBZzMystM1
6RiX+tcC3mAhmLbMIFjHyrLo0tPQ/oOL3Gj+1Q8rMiHuoZNp9f2wpZ7WhRedsCQyrbxKWjkvtwL4
RU06dI44IZvDIaXmZZAfGW8pmmqAE98g1dhbIdOdVDiN0CQ05U5XlnwG18IUBUAtx+cy8CvMJajZ
llbfDGeDCyjdEOG7qb0hfvKajNKB0WjTAk4iLZcUKAh7cr8jt8JPUKN0aiKXA0UkmVkco6s8v7Xp
nO7W2AP1tLBI3LTP4+XstPpD5fBb8wYzQJj+RHFvUKgpWMNxB+WU9KrwOwQt6PBleRolOf5X3BIe
U1EUcEeqk0jsJ9mIJN8LJks4wiTDYeixDnowubNBwjg6sEs77u++MC/FbtmRK3ZXCFugJZrMcIk5
1hmO/4q35Mz60zsZnMj57UTy19HZeaaedytLhNlRWzABM0BUeJFLNkJvJpgX3qWUvEZQZ7UnrvMg
6yMsB4IEH1S13MZQwKpVoayiRUZObvvY62F5eK6ayC4uAQpqIJi8IgzcSnnCc4xlAEJjzVyQgg7n
fxGChC2+NjcNo68SsENAc/uF0m53mDiB3qmZ5ctoxGE+Xpdb2DdRCqR4VNV8Lj3rXPOvV265LFk0
z9iMovx/2/bWAeSx4MD4wbUB6JrEOB4ZQMpMs9A4sS7dmNqI/rC4FviETiCyQ2cxZodBI1P95285
DxG0nZdFTL484wiwi8hjB3XBMU6vqpHba5Jp1ERbQ9te7JDtejM3fsS8Hz9UALea8YQbjJakAcTW
cTfTV6VuX73LlnBQnjQAqYBScHGuu4xqwwgE0z0WegNz8lZLcmgMaRmniwvyA8aQfeT4tg24N4SD
VgVZX4LlWfBIk62V8deMHbxvA6jD2lUiOBOod9HbUBF2QskrxC00QxyGO9uhA6HmfTjciGTdyYJ4
L2ex226ECmkrffNedObTLfykSobmGa1uUMe7ajGqVjkQ1zcGaBQLrlbdiU4MUGbGOfgIAsFYYC7H
XbJKj34DoRWlb5+wmDIlOx+D6W+ePirP+p49vZKJz7t/LAuPUCHobSB5ruNzFcsRofmKKxmQ30Jg
BGWTge3Bmc7KVcT/lqV2YKhAvHMb+E4un4UHAjeDS5jdcVsttCziKTmdGPmZQKzMrIuwdCRkzjfu
Bcs5OJFDejwuLNDGRT8AcznIiPTHxVbHlxiwU7SXnhKzwBR2mOS1GefmF9XH/Xpd7WKFrch6l0eA
bVjo/6x2uYQvldrCxiAUvi+NeSAKKaESGqAnjZTRMUWb87wX4EUSvAh4HDjXh2swExLdngo3b+b+
TVzJj9paYWncJc5LnY9WU9JYnLwwEoltni9rOpv0S6ixZ53OUGUYUMILFp6RGmifWAHbEc+Hafe2
7TTuY/5Se7bUNQsdsDi+BaRX1nYylM8mRF2dvpkdhw2L1No0ljymBPCU/qUcovDicqB2qXkJZSQE
n6l+MaL+RBSPWiFkS5VLoeuY2CMYJ6586/0RkfHuV27C7QPXY4fBzQh6rEN2abKnUGWYuZo+Vr1f
bQCLCbpXM+0ozx/lryhnPM/O0TCEwFKyicwsx6g8oEIssFxm7pi4Jy+jmawFVLG08hPkbip8NsWa
kq3TLkTdpq2jXY87Vmi8+6caOgcQYxFuKxSW+JxvA2tSTwV9rmhBbXmH0zGYTTDwC+1DRIiA+7fL
Bdssx8N871YOjkHccsACM5fNImeYMQciSfsWiEKJZcspUG1SaY0GuJ0+KXX5+adkp5qXmpl8Tyk5
nJEYBReKaZfrL5hStcY//FZEt+NwxyPos+xqOlfXvL12GW2hPQDBrclIhExeRPVdgLhmWMK8vzha
8beUbXfjLGe/AvU6/EW3V7R/20qpV2FYsPygk6EEn9PD2/A7G7FktarNtKfOgSaj1v5wpdBrhMdP
wib5rK7ujJyz0w04kAsU6PoWqSon+L3y3UytSn6mO9SlHe+k7pezPYgxi9ACAxctzG56K/uwcO7s
0ztVsCFqJwt8gPmPqFYcrWtNHW2KVSA4xn+J0i0AY9XuOz3wKXYye++FXwBk37+HR4u1ku3DzuJU
kN0lQQZWdldR7Uztu/L6hc8gJc2P30aMLZFHXNhVr2eVhYrCq2M8Apl2uKXfptBeHFIVhIzUjm3R
jVxOQPSOY3D1doTY5g3TRYxA2FX7bHD8/ByUrsYOpXBm4VIzSn0kvrwWiIlzvtNdkWRLnuXiCgKp
EER4/YhlVDMW6cGaDBjaXseMXHhaJq5vw2Sth2ycvYRpwTRJulBmt535aAEmAOwHNnfJrmNn5Yor
tL8i3cmQvOi7gyUH1m2JOJg7UeI+aMP82N3782F2VajH+qu2Kv9NG4iFuer0Xj4N4NTHRnH7y1To
noHCm62cC0eZ3DK8hpHorRnJ8bmIEJSFvQ5uL4fnXr/7e0WQkGKPbWwBFgQ8jhnbSP/IzClfeFJh
jEBlwahhdsYlW/QIoGBACQCj6y+bnQcfEU8KAHG8lAfNztS9xhHwPjyan/jAznjTOFQr0N0l0C4N
dPZBfaVsD1WpEtDmIvaCXkHhCZXmvqUzPZg3cSwVVta4gGlk8NVtJHpqg9ugh7A6iNMUe36etJqO
pdkf0M7UXfS5yFlUBlGp3p0k1V2sGO7r7RAxFxIg1zKRZNdCS1IzUEvgRk3/ppd4yaxO1mdDpxcm
ji0GGejxV86WBXguNXf+vm33CqTUY0/GFEcozElCS3NsnTSV6dVm1V9xlvcUSPUPgdoNDdqltosy
m9jSKpblFMCWC7UfSu5ktk+ukO7N+u51b4CshmLeobwjXxm1y22M+dRA2rVGV1zIndorAq1le9oO
DArjwjbusdp/kJXp5V4kWZ+/4qsim39Kh9ERfpzbAt0KF5a12IHiXKz4qlR25+rFuit9ZYUe6MwE
jkLpO9Grb1SJAfWfuxvcAvxs/bRCPq6T7UZqez+Iv8uBe5aQDVqYHo9MmL/NrC01iq4KHdpposuM
Kvbec6P1WDBaqwwOfLtp5GchepO7kvTWrBtBLRHx5Ub7z4B9alMovkrWKCvgfcpZAKLg7fqNO2Yg
OGFwYg8bUYez95h6E6idHkBvvji2ensBxRIfpPADNQuSerdxES5s36WPQtAGaUVWWkNhUEY3GLgO
LmlBL/lHsr5+fLIsK+wrFkCSTgwlRAUozmfPcz/2NzqGHcVARYApDtzTvemM0tmMg5PtAeo73GJ4
GX7ghrDuxQc3/buSq7FVrhgF1UMV1bZD+s4tniQ7gJnwWCAYhvp/CpmU4cZsluW0ISM7eqedhPKg
pVG/EBfctZoXkXyKdNlTkZ1n6IjdWe9Rl7uhkI+JXgRkbiEMIGn6yUMbWmGdLvfB5QIZJtJoGk+s
h9QQlQm7WXv6tIApUQjtlwqUZEMZG5y3Zq5RqQxw7O14QzE/7fdPjtGcjPeA/NA6NVqx1SbGCL8j
1JBkxDPNl4Va5y0ixbgAsW8ewwqcP808nwtnaU8/lxjz1s0BFF08ZEoyaKYNUPiXR+8NGRY+VwSe
Ur7I6Mq2RuoIO4SZ8BWSSA7dEa1qPWi1H1bRfD7lZnmIMnnj0wp9WxgQFRBGv4Qa6GMtF2F27H5L
ZXZ0O3YTYrKri24XDN8PZBVAaqtJ6HloM/uV5ITv1NeJOXbmygNGNAOXpsPbOgMag15li7+H1EIV
4Wc+38tPnPI7Xu849fJtcFX/eHA3b00fvR+XBJCn129z/TtR/0/JqiuYwNX1VNMf7e6JBHB/9Zfq
ZUrItPvssLjJYmiQUyoQ6608zVptr6oi5QanCTnH0uJ6t09JHyzszi76gR5ZwfzS3Y3GYsfkmXl8
AODcCpqg44jQya8r2dS3bVobu9mpetj88mEh9K25mTefuzEj7EaueUvUtj3Y4neOzrLCLbqfIHn7
gAyUn37tNaVSaZh88y7BAU4ke49k1xdT8J91xJvozkeoS7QkV4FzEnDR9WWetbQhgSWp5r5trpTG
TGy+y9OoUDX/YEcgkZPo7aw3sIlxVtPs+oZsNP9XwSmFwnByJbIA3UoCfmaEgrt3+JUisPuRUWy2
U9sOxX0VtwKKzqx/ZlIX4VE79BkOxPJGDMvaAaBikqzqGsKm5vXAu85Qn5qge9GkaJn0yTCo7Q6s
sy/mVsmUWvRKjFITmATIDWnGpY1fwPnovEAFiiy4jCjl/3BpG9T1986L74p0M28dutGF1Icx45S1
oOj2lmdu/2W/1Le96ci1iW6wdQa8tJCERMpFh02Rwf1RGwV76e5bvIUUiMY9lLlE/twxS2YfGDbe
NOYT5RJ01aVtlK/oY6oYPXmwYQii93ZrrhNz2Z1kwtVeG3W5x99i1LL/Xp7OZQkUcm+ABQtEGh5P
b0zk7NkFlGg+0lHjmkmAA++g08Jo8qqWNgz/H95swVjg7MnzXg6qdmZBo8SC4ow7nw5715TJC1SO
Uzj/AcM6j7EgpBbGIsj4lnx3PjDPFgCrHCVlz3W8QK+frtq6ws7dN2EdcrXxFQ5pqpjhi/odScKp
B6AUVzWyjQkTrY/w6dS6HdHD8alcfYJc+MWsBwF4aa2cgid6b1JjvL3r25hGpyCpzPVPMI6DN1Ul
fZBQNr1+H6o8fUJHjh0iPD3pBSwSwP4qcngq9/nSDSFzqU90kRT0bt1nC+iSJ0e2S0UfhkSDGrBA
ZsbjKtrcIURGl+VQjtBr3yVdzGx3sWsbz9pTn1BN9BeJR5p+v8lT3LUKdZzIiZMxw9CumHMTVk6D
sMZxDZwvMCfNpjLNvRc+82+phJD1lO0iw8OeFvRNbndSYG6bVfozkv6414+aW49T6djpPnmbnsiW
XAj1CbLA3gYNrteZPmpSY8xJexHr/wsalfxIQX8uSag33QiaL9uYOuh6X4XS6esNBMKSBHDjl+Bi
iSoXLZGvws/DHkUDHZRcoCUVzjppn7npnJTbPsvxnBuqH+vxbNgYxw2SHsIe291gY5dgv+XfAJr5
6mqgfRvzPsd78DATOycl18aus01AcZ31D5zZe8ctykIKWOnGCu9rH6IeDGid1DlRsdKDgBP9X43W
jp9jTpBc9WXlIixQImYJZ/NkLgtx/1GfDtrq85K+q92pYbMnKqbH5pW3atxxDQrEuMALvxdA6ScC
Eq31KygC2XjoPrQTQx1pRM53OnQNBb1X9YWMXdR2MisdaPQoQD7Wzlv8CSQoyEKiiKA24oqZCRQt
n5c17T594mxpstQniICrZFN6/lrtTfP7yaabAd+HEdRMXVYU2g2acqzg+GMDTPnvGo5UyloQuPf0
OYSD23KyasSsg6KEGmsHgnwWvUEPsSlD447VThXYQY0aYEb6KaboGDm4mJal/sFNGp49y7+gH4TK
B2pdLyNNTDWn+5QdnMhMes8q2Q8ds+5s1sjxr/3FXMrgk8gdajLH1C/n0hWjjHGpVMJF5MtICXsg
CQocRsxgGkiBHssIVJbT3K9P+ZqYuTuGNy9kYjGwQxQ1dr5fOuSjVj21xu3oIep8zDw0TBdoSq9V
wEME36XZlGkb0XAgN6cDyAK4JGj1UfCsNseb7PvMtoJnpQVIZR1BGOTbSRxMytCPwRmheNsUh+wI
Wx/33xrcGWl7wE+VdwTEa1QgoN1iTo5up4poJr0ltoOWufVvJDO3YNSFGzlklX6c9YSNmIeOYcMf
+KLkm7vwCpRvq8KGhtPK4H3hhprSGG10+b5d6Yuy71oH72dhb3MpSCBWsvwm1d3/TAFg1HJfXzYm
E3cT4FDf5WpXC18n+agFMrvZf7rF8dp5VZBwsHWNeYoV/7q5puTjRCFdR8rZtaGprqr2ZH5BISUV
z3Z40DhwstY+v6t/8R0w2eQV1XYqXTZu7+9xRx5SjWbgK5fxFqQVZ452GJlUxIKnc87/hG6RWSVA
SX46j805MQYQXtXA1VZ2oQnM2Wh8brpKkrV75LEXeU4zzTGJJxrvUzBOaQ8vfrFC7EjsPgSa/m0S
Ur1cREbaEx2sMdsMkjRvain04mv9MQdcxayqwjqAErLFYrHgFUinB315juc6IVMJk8M4CcibD7Kr
GSIzN/AvKzzxXOosh96oI01pkhlJhTQwoiXUYgtqL1kKU0lMLH1Lnat2nvDh1aiBmKOSaBaTM9+g
UI2tymwTDa3rP1mznzxFJwEMwzKZ9LtK6yc0hOKbGz/MBzFhr2iK2dKIKlHSFf/fJ93FNL7h0Vn3
Aa/FFu4AipMpS7KCt9vTaN8uNASKKO1m5k1V2//ui1ASJnL2kUg7LyGUp2rDPkyj7zgCozeaXJch
KYy29xfkZdD78WtjdJQFyKZzDnZ8/0vB5UGvqaGn47cn+n+KxSBqNjPRy3rkIhIdy+/5ncSfw/vU
jB2ci1/BHjgLCI8Uwv0+FUXEgDxbc70xs0VNMNSUdTrYmZGnDTqr4jcMaXL9nGSpuzJYAOgp5K0C
m1Bn4H7yE9JNIyNU4+LqwG9IQKLNsoz/6HXAPvpdgtrMDwctIyPfD8pFs7LzLwTDEgpSp4AT4b05
xFpZRqWJF5BPSsC4VVK8Fvau2IitfeWNytQr89wIokXPDUeXpfwm1fnCz8bFGMVze5wW78oG7Bxy
fOGgBd8oSWNBoKAWKgcGME756XM9j4/yB0fEVD9oCfXd98Ev55zsyohQWOcKnoc8ldgxe+bEMlQN
uotlvGtybC6kGwDjo31yFhbalLbCa4fcx8ZlvP8ZOYOcd1kopVJkAOe6vFVty+cY7sj7Cdmq8Ve2
TXGGQ8ScKZFRxBnkwPOpyZpLVUUj20/SbrMMrGD9Y5sdcwtPCHL4wIOBXbAelZlb7Nx4hd0lwMwf
rnqpOqR6n81WpkfNGsAymj/MD9vxr5woly+vcJ5sTHx7TU3eI8r9NYvwHjqNDLKxTcy4sBQvIx7T
G5CZZandR32FTR+YQzxAaSfMG23BPh3tVzKo9hw0FRMJ/XSRUrDw6vHXIgTrnWTSVQWSKy6QH9Vw
1Uca3NR2CncOp09hHM43GfoiSZUZ7jx0Cd/L/8RKr9WuM4G3pvvOS1y5wW7fsG9aU0RDeLEjaVts
xILLAGOtbAz7OiwCymNWfOI9hQV1uGkav9+s1VV7Ta0QpflFxXX6VxYyNQ71v7HR77kYXSqE3/GA
z2/O6FId+egsQCGpA38fuGYCu1nUrDEqg6nBvsTQpJy7Y1BnrMzXjO7oihhx70FF/UB6nGJ8mDOL
c7Wr93PwQD/n9KyBGqZEWWUeeARvLBEJ6Ay1zZnep3pCg3tEd5xXSSDMm1/GaMaCe4sv7TPVvOGM
QXZ0aRYmnvf2d12NJQ2bovbNo7vlHEYqd39VcGs5IdE/uybmDcEPo1D8lXbAXTgVJSnYyTXyKtDz
WJE+3gNhGLWlMjMjZBgp31Yr1WzXYuto8Emw0JagKFu40hN0O5i6l7Y6IUpF2OIo77Eew6eMNc9s
wyKY8jZI3Bmv0UbvehPmaOXa1cbfZJgcZGrMAi4dGx27n4GLzOFUT8iJ/5V9ojpJ2FbLSoRQiABq
ogBFDv25rNjX411a69nuFGXIrUHnJ+jD339KGQajW2hTqgMUMRfMrHRpW3VopVsDEi3OyFE2blqo
iPMB1jQdGnAVTpsGRyQnkOeZxdOkloSFQY0Wuos2j6gOnYM48K3Ue4QDr6W8G8XzVY1zFVxe8b/f
y8SKWVUKtI+f3mVOKMSudVaLPPiUNrcikoQEP4HX0KoBlXrLzr/jNRwD6xRZ/YQocZMErx7JsTQW
dnTu1SPUBZoiInmASlMzpRZXueRV4uH7s4/lqBDG21s3xAZ87FLOCTpAV+7z9Bpqadl8JcMjSTPX
+4lwp3hsYbXGenRWpeaIK47oFPQlj2svHMkDta+7aBB+zlK15F70m4lHGTa70kryKRqno3TbniCV
0WlWhdi4gByucr9KymOj/v+O95iK6mE9i7+uzEwme2UQCsfGFWX8zBVCOJ+w7SF1SfYkJEXa2dNN
M4hbo0Ck9ZarQsyGSvlpG2jnmrreN5wHB2HmcDW9mLLzPvvEM73fXayw89dG9/J6VSUfeM4I1MiW
fO5B9vWH+1wS3LnsDMYLo2R+0D+oWe61uL5fpAO8ZVZRbEXzgtikaR1TXErzmiffRLWoCBivwPnr
5w0A3nQ/6Uyg+k2XzPrr+QrcYUPtLUVATfec0BHk+n/JxThm5l7tM0kSf6QPODisG3qL7s6IGJY9
q+uMNwTaDXsCE0tfgXzKGk7fmxbU/EZ1w3KfzML50H6ofhVQq/F0YGAEnZHqEFj7ngPDZiS96KbL
6NGSTmdm86krmlOn3QRu50gr5uDLvyPjB5142xrYdAdHgIsgT8eZwohmah/nwajiIGoRUPsibLiU
UmdHU3TTV5R/3agF33QKtkdlQLXpo108WosSkZIL0ujqbZtno9bl0zv0AUpoJJ5uVfBMPisTj9rw
1vgS/f93h0VW7MbvXkP4fjzK4RKIqNLrLyxPqqO1/QM7gmQ5zdYdoPP5Cp/MeKhI2SCV2RcdDEnF
djW99RNez3umDx6xwbV1S/qXWARH27gFtmDE2fU8lfbkhJh5IFh5AKumu8/CzWH3+AkVDZgjFCwi
xSgSUZvwtNAevpVhM9Nd6bHjmG+sygaay2sU6fKzA8VFc9aXXSDP5+WdMpOM871M0CBns57v3V70
loeY0AbTBrNMyUuWZuWPsfPSzasb123urvBQa38JBJnWPcSIU7BEZcoBYsJBnZYFx39bJxmTqud3
77xCc0CNwKLfhw0ZCcdV0PhMfVhTd9NgcNGvPp6Lhj9vKsyiLIv+BJOBhQAZ0dIpYpXkw7OiVdlA
CKVl1rBu5NuVuPLGcQl6RRBoHokToKDgwSokC3kjHfsIfR9XJv+Y90M/UGIumurqGwl4/zo+wTlt
NlCjZhmmYwPPQXWRFUGxY1rVgTMfVkcOmq/vVB2ZKpX3vBFY+jDYiNKmPe2CIrqZ9MQiz8lB/fy9
XFDuMk3C03rwD8uh/RrWZz5Ol1lcZ08zSnuz5L1BEPKXnIiL+fuOgWlV0/h+CdLgpcN9R1i38/fh
BeKRxDVN/DBAWFB9+8YmcT2wFxUuAo3Gnm0heImhz6FCJ/m2Uwf3Sx4WAj9PTwULjOR3o8u9S6QT
qMnsKI8t9sFVZ49a06GxtONb9FLBnIdI3PbD/GdtT6g+StIaH/xibsOAj9BZLT2G3V1kAlXh77oc
bcKlkKU/CY/q7Nimb+NU1i8tLGSkcdzAdzajJYNjr6e9ZvNfsteAn1iVTvo/KFQK7E5kDjTQRPik
0LZ4NqdMecycqYqKU5GaVeSgNKYGdDfKPXwx1GaTt2KEunGaydFnuI4Wehb73JI/71TITO0/J6ie
wbYCNZwCQLVVaaV0XD8O0gGwS0hC7/t3J3ZczIDSOO+uYG7HVDFIJ/bsQZdASh55GJzuf0Hr8BOZ
qeuf0nGiUcMIv8NVI1r7jWj22eLq9ooIYf9hp5tlfk5gauq3KbxU5/B8JqeouxSgbP9h5QnD3CGO
3LaMAD4q2Qx7mKRa0ZIa2wxTfvfOzQE2hGRDVEXi/f35tCc5FMYy1zmHhRF/rCfQNwSdvvKO6hX/
dIS1rUCrMdtRIKo/oSRlSbMQyWO/yG7KGg1aYL3zk5q/Mwf+L8SONV96YQDY2k3eDC+YvifwLSKg
I2gKf0tnwCUtQ+E46NSsptwL890o/D3MNRfG/0Qf+zn9cF3O+NFIPrwNRz/1NuZtB6kRWkfQdHS+
LDM09QUOs2Vc9cR2BMLwu/DpjPkvjQSkyC6wy9x3pB0aP4FCuSZyApLHAX1DpMCKxgOa0VjE/qUZ
/1qRX9NjPQ7cVWBVkS8ThS4b8/Do7FdM2x/4aA/r/a9As6ayaMdGIdvk+i/kjtowspo0iXRG4d63
iAMuOZs7t05wU7Qn/0+8umNLCFg2+OLjgqcNd3n0ityxFy2bOrTwoqOUYdlUXRV9sroqgHd3CutW
ycduQu6EwsA2DK31dV2GF9wHBHqNgXdyY3egcL2UMfFmybIpqyE/LjhVIIIR+rredEO0EDDRjEas
phNUUZX/iEVEmb8toYVmlgekCOJqJ5ts6pi/JFrDx2ZqscnLh1nlvGQcyOdMcYzpYWWd5YB/z5k1
a2vyrmJbMBMFdU7s/MJevNpQJjPTsYWeX1dNsiD+NN2ZAiHkfFA1qGTYRdWAdu8ghWkBmM+heymZ
1R1+UbOoKc0h+ry+X6I3Soif9nNks13wtZmY4uCQkh76hVGYfqN/q/wCROvkujHq6aA5vaLL6Ccn
UMbusWK/jtaRNbtW4KZTni/wT/UiiukHmbocJV45ZkHEues3qTR4sbFBq4A1ScM1kUwA6AV5nt/Z
4WTQUqLMlx5Og5AW9CCxfykloM6MOsSSO6xCNv7Y9gmtTmkAGVeNANSgtnjWrLiDI/m2Oojqu839
/PHUnqRnKpwZyOV20pg44/odjHkQks1pw87ao29Gap8eyK+gim90uUzRLBjF1CgwCPDYhSorYUUR
6UypUV7Tq8GZb0yRohlNOwuQvDt0gvBPJ/2VwOxkQHESXr5uXpFjL7RdwbX/0hXb3LbMaA1ta4sO
x1uAszkr77KqbA41AaLye2kIlmfDZR9p4Ce96fNBVxuiEUOnkBJNDRb8keL9f5KcdnCftsilE8xQ
nXJ6pQLkYh5lSjhxqmViDDhkKcq7aM7pWpHAh/ojg36xgGvnH6sS+r4QW/uXAQZwxli33cGXqfKH
BvtUYshsItwC34PhrON3MUQlyR5vYdLfgyWfyfrGYhyeVfOmlfnv0bXlZ1YBCZYESeGVXBccZLL8
SpA+4MdQjQs7qbKZi8HHmyjx8a0gBxm2rCOraw29TDqQXxxE1YgXcN0bzIbDekKKp7X56cq2qMUG
gl/xgwOa/5DZZDiRxUi/X6RNtVv7fZTUpGTCDZRedgFHqJ0YEGBEOPEDu8GZgxlaQ0pW2NLBiT6Z
pgI86fFasRJdogTu/894bo6aI+aoJ2DE3eqgcJjsdM3d7IOuyzY6hOlYkboF+Ir4gq3Q+0g1AhBd
02KUCkVpzMP5SO8aLpSJpBWbqarRLQfDM5AxlH07/SyYidAL+p4TNPwIT+YZF7jvDfjv5UcqBh7B
SJAKX9JdrZ2Z7hrztS1i7ijwWVJIGNd4jYjd3kdVuXZxBX/B+ggYSzPqOL+NfwWIgi+Rbz7acPz5
wh1h5brNgZoiHnwt8sZMXNxo3rL14BUyYfLP0Yu7C85n2UBzLGuxJCl0rM2ytyKp3oWXIpTzSaJF
tB5RF+76PXz4bzXFBhrGwTw5CbrvAvMyX6vRa3DW1veFJSBDt8qqbVcugUAME0zyIEO/1Dv7kz/n
cCq6TykInbsW/f59WfZkhEitfG9N6asOSVbMBGEmFcSjlHc9Ph58JRiyUqBMhiILMaHorzKlxFFa
hZJgajj11zxWoaE7rQw/pQDLY2WX2pqGLYD2ZSiSueJmYPZhd3swstVhfJU+XCtclyz/5tFS9qo2
ynktYLn92sBZY3mQW4DD46fGbsYgZNZweCy4KqRP+xeS9RnvjDO6F+V7cnCWiR+tsC79JPsEIKiU
t7RBuYthZIkyU0rmeiT5A7IWZXHHyUXunC3Nh/oqProkpNUupyKWAQtXvzPkYRtkbNX3siEfm9Ka
HSfzBBldqK5HrnYQqUJ/GcZ9UzVwdv+6q9W7FbFaq5qkmbbQ2FD7hR0CaWZ1X9YrU7RaLvRll/kc
X2DdY+qVYtRZO7ieGQtlY+h7hJN1bEk4r86tv4I0THalsZtLolNzWSZ1YZo3fvekGUalAyofxiqS
SSKKAC/ysTcxn432MGxWHhtR96vghl589wewchRy7Vy27ngmLTsvq477ZH+Q8UWtR/YqoIMlKenk
vaYegBmiZiiRTJHqGt4V7InUQDDGS+EAXzT8WVgBvIWiR9EuN0wRkh6tPM2ISo3TDc1hPlbL6PkF
Ki3DQJ+fg0S7apQnZUPQJmF1dEPxYNE/jqNbsriJI8hFa1MyKCmnxNkca1KIPdrhVt6Og6ta7z4g
Cu3txKmGcttYSzQdF59cHibxudbt9IQXmxQus3wAp7gBRQqvtEerj0VuqbsklQFMQLD8Ij9DpPNu
yAbGIsVLn/YCzkBOr0RZJnmbPIJqu5TnBh53F2UiICrWG8iPmDA4EaDCFFMXIAv96RljS4ojKjdq
Fv5Srtob1QGxLQ74AA2ySdmH7ex9cPxLUU17mSlKVKJJANnGsZJUoZuAjjcyYfAApPw4NATNjnEW
Qebuj06+y9bfCtjF+67yjRIprRDWlfL7xI2lJnES8lDJyK1ufqbfoU1eLrHlFEWOw77zSasasuVc
ax7mOoCHELK41jnD/W6EXbWCuZaJy1yABgb8nIxSQzvBPz7J+gTFD3ycmnfPGxo8vzIcK5HuBzO7
8YQJviyfPVaUXD4L3YSj+YlJYd1Df9sgNttjUmhR2UCJxHF6fCY0VS7ogaYwjnzTBZKTbnixxiey
rUwpmgN/Y8QNy4Ktid9cJ0HxLWpPvxVpBGqoGNO7k1qB3SXTd3ZdniDQlF0k2yYWJo5/NsW3+QXC
77CiiS86dydNZZyDxBixLj0kFobmy+zuNd6Aw+j+sCcgyWrI9Qvmxg1C+Vjnr8SlLIQdx+YHvQmv
BlcBS3cbTqLviVC12iUqaaJ4pN+zTMhO257OB5u8JQF3FKfWlUh1iB36P8LdAchT6mWo5MuirqBN
7ucG+wCJysMmnQJL3bL/B/v9lk96sRsY6dQN8CXjw8gdioKbvJxA5TTUMdwspm+pOp7XV0XzCyz9
pGxj+22Nm4gxBTVPoA9TWWSx+64IfV3f2LzOaGTSXJbAPPzUdb9nBe1i7hq2HMdQ4dBGy/4XwHBO
Bz39E9UjOPaqrX/odA6OosoVEpuBWi/FgpO1phdj6O7HMsxZ/mEQJ/Zdgogt/0+3ucLEq/VsRDTL
qLyKvxpJo/GyjClKC7rjhvBDxw8kVkvyzdE1sFlybQuAKpafHQhTvNraSKwK7Nj/1+fuyZv1ZyjY
6clwAQnSN/wVY4yrw3qusA3g8BlYh7HTSN1FbQBDqTW6SnfNBO1UBevYESPCV8fgCizY7aUSxptf
Eh2o72kHWcQ/aggVq3ONhwoTCE1XTVVt7GwXqD79JKJm0csatBKqazkIA/QN1r1OD6ViUWw2b4eE
zh0Qz6n7SlwMnsi+/eKncUXfQklBCxAaiZFlOWzpUjGIuxh4PjVoZbAdTJwpOsCmJkCamOqD7SuZ
ZDrrkczhtuOg6miSwfQK/jHSVgSG9WKsscljcFsbmLh5b+RCAtvZ2muRYIWpyNibmq91VsqgCt6I
vvo4iXzBlWRjczdrISr/RBlOS2QpLfWjYi6AOw9Jd/lYbx9QpVs26oCfjSTA49fS8MeedJXe6K7C
FIUo0V+Ubgao1tER9NPXQpafd9sz9FqOSL4C44gsAmCLV8gfaKGMwB3kjdz4G+cFp8sq8Cj5wKNS
bgl4fsYPUg0XP9kvKQvXGzKsAum+7jr1Rj1xtfNTKWeaPU63hK5213BnQ4Bir6eigWphC6FqIlfg
JBnsSFPwge8C1k1Obo/hCQSr3C19pBLHHEs7aGpiKVaNbSJryMSQcMFByXxJpRGQ/0X/IQKZ49ru
FLobm6dZx1VINllXOcR59f83nThCY0G2Bt6x4Oy0bri64Td40HP1uzMGEYdBaRFknP6dvLS56tUk
QWsWR6wJrzKU1vy7NJtfmBQxMdYLxZoHO4t9C7eegNuczuCMyFhb4w3Zl7tuJOGnI0oXjtcBMz5z
KDe9XgO2OY63VbeWTpEjZS0HNMZUJyqsFIIp/r8wpwHF82s6j9rCK2Cc3MONgum0E6xI600uBZeG
ZbWv4L6ejfBR42vRPI6Uo1oIKwAwMl0fUeJuj4yBWL/tIqN5H7BnIv22TKNluzrJWDnc8c5W3MnG
R83t8FbWr3kdxidlYMOzO4hguT5/7KRNntHaryp907FXflDS0YkgOQPoOKPaULVLlXRF5Al6xNgt
OK5javJ46uuLueU5IqVsbJOwRwjFpTvPO/bq0oBWYbUgMFY6UjSVG2tgiXJflCRPJosIvhhKgmHk
ASeQjamRR+Qbqt7QmemLebmz4FpK33b0ixA1exf4TGqJuOg3tlgJpA3oETOhD3umam+IEfDt6muM
dfLnmr2OlMf+YoDbPrSRC12zJctpmr1kuFGCw8wQbReQe0vdIrA1pR3uyd5EvQPVUve0jWpDXsT+
AqBMfIYP0gmKy7Rs47z8EhM9cxb67uf+lYU15zQkISxqxiNSJpzHWWGS4N9aA2MALIREMmDFfqsw
fdXD9V5a212uVVJuPYd8O5t66gVOGnzrJKJXAl3gFDheBxGV2Mnz2N/+Go/6uWjMpXlsnOKvq4+K
LSolfurBIQkyIVOx3S35E9l4JbZCVaoYnXkIV4+EMfQO7ecg02F5q1gS7RWU+B+F6q/MUA2IKTHq
f4Ja6WKHg95tS+4VAXvbIYJlxfVWQkmGlJvu4UE4iL5NVYB91+sF6o8WLATTkzt1L9V0R8C/v3pk
K15k2jVEg5AJLUn+7lkV8FcPk6KZa7aagcFseo5jKF2tB2UirXclP4/EyjRbeNI+96cxprB8cy+B
8lg1s3HDk0FMOE73nItxgSqg2/oy1sltGLMLgsRspRNrQDf102JOK3a5HiFO3RnW/qF4QCJoE6Ps
oeSWPJ39jju27m5+3CfTqLJtWi/8N+4aO+wTYtIngI98Zi5P0hyo+fbAMEOwu7Vdmjle0GGtXDK+
iHPM1MqqBSJ6YnfFpWkSnTnPTj/uERuqlhhFsOmPv5SQSjb6paIQBYzGNd/H1UpdLm+579BS18Oq
yK81We3qiA5WM/1eFkl41IthCnH4xgrHbSobU6l4GQJ3RPNUIQKG1WDO2VnT7IQNWbov4IGVgxJ7
v0uDetwICQ3v+S6ILuxDczMAKp9rEv7+R9Kd0vDq6M/ZPh6ntesXw6LQ2W4UlTY2KmN+HwYyoqwn
GZCs3wwZ6ChNGKljB0VyPxqUlwGV5QB361rz7385qFkMq/E/46tA5QQmswvZ2wHHh90QdxTuU/cp
yjmpm4qulx33ZFlh1s/KhdF7SBYRGbRoSgGNao4xhbzXr2Y681/cfsiLxMzDVtDytXuyNBI5AlAh
zoCN+ytnrYrBnofn1tqcM6QiSfDLiHRXU4WtFtc6kUBcqH9hhHH5qkfWgXLr9+MUbroPP97hwnix
bNHvi0iFyDil2rkPlAK82unBEw/jyUbT+jGITxWAbOHV6m3Z1TiAKl8M8ahZzodbaCHB94Ta+Iqk
/6E3oWszZGj4bG0Gilfg6uNz3OkwDFqC51Mhen0rZk0ALPcD1CMbe7xHyLLBgdibfMUKWSYYaxzQ
eIK9wIpgqshr1KUSjFCLnnrybnqdvALpbRM1pPl4jOTiFKsGCLi/IeuLj+n374Y8Uv2mLvHvL6jb
GmeyXyE1hnFhJta6cmOdqTybe8n9F7VnirsUgryu0b6O3lUnGY3r7dKA+fFewDFNpnQyOIyrrBU1
dsymzqH6tVzFFv4iE4leqNMSls7rU2eYvSR4MgGhQ4Y+RJnfgLDFoFEOdFCW2qkYUyF2mFV51Zbi
H5mVJYcyLBTjLySnWqCbuqdAfSt7GJsbsmli2ebxoXVGZzOcbuf14x+ZBPXEQ18BX1G5HCNRntIu
r//Dy1l9BOYy/6n0EzM9NRkCNpU2CmU1bx91hQIZsH2L9KOtxyfmpeNzuzxPyfT9RfjtNE2fJSBw
OFvYsqC0zI+WL4qTiDvA4DVS1UJ6RYmGkoHHviCl3zXv2Nh+V4nMZqBI1u6D6jAGZZj4RkCJv+j0
KmCmtO0Olfp2C4nWUrpUVRLQ0acQocpDJ8A/mn5+7QOJU8JFQZm7BO34O4JPeWwTm/r+pCoKRILG
VPyOU6j5MSqKToPggCqENAKvGCp62RM5RKMwWUMFJymKrRC8hkZzNrQ33+YL2U2Yk8Oog76+TlEK
gd+Yf8CQww62lv+G5VUUm0idXK4KidOusJIuNZtnx79iRwxoquDrOk3bQcXIQFQiMikn0Bl42gjH
CV7agTdBdvsaAVNv36Dk7RimNlzHn4+cMrj51CskHRRIcthequYrTrR0sbyEPTnpVsM+R2z0BK9B
ZcJHwoN5+pniAY55MImFTuA99UMOP8bCXidiBBXGGL6VomV6XchPYtwohiFEi1lFdjRR1u1fe+t1
hCqrlHd6+ukF9rrOS5AgXoQNVZNBaj5c/yC23Z9C6KFIUygpo7ToyWbiEmVjhTP0F0vriKYGMLyz
Q60ct1BcfWUMlbHU3LAmyIerQ8IYSVCbDkBx5ct7KJtj2ptnPXbNC5XxZaxl0rlusOd2mCNLl5Ad
m1SVYuldLcM3HgcJIXQnk+BADOU3ietHpTBlLk1Gt64Us5EanDYCMgbk5v9+6BN/MhxmphtAnYHF
7Wsi4ZTmL5i/D8lfmdV3Py0Rc0uJuHqp1a/05AY2e2eTxY7t7Nm+ArEmJNBuYmWryLeQvR3ojYq1
nsCbfMm7B6fa3cMIofhEox4RqR1RFwNsxdo7B5kphwfxrnc3hGU7K3miGHQCnX0bKBrjIYx8RRcV
6OCeqCcNRyc7YQYztKukpQX/spENKXESQXlHn7V6jp2GnlWp7D0gzeqmIk5S9yem5wdSIOMkJAj0
dnijqdZRwsX/4Cq8Xxc26D5bJlj0vgwO6w9KFtkhjWVxuhRHUghS6P4L/E60zBMS2l5NuHh6RoRM
N6R7ceUG+USiH2Jvn3IbX6txolt4MV2AvZhxzXOQhX8+L8BLzhx4bK7OM0oM3l6EjlLa4ZdLOP9N
NJVYA3pu79v3BAZ3c8gWLwsbfr2bb4rjSb83uNOibisy+8I2Ga7SZm02nDq2JQEPdAUxl84nz4+p
4vT+eOzzDxH/RCjaEwIl30avX//0TBoxy/xZyAkMUTl0oOgHSabDIZXouE4OwlAEd31/CXVlcpm8
UhCoudndtfL7wGiz6JPWa8ouNt1WNR7UPrgdcN3ykB8jsSJanuVS+IBKbRRpuzCIfzxtr+61ei6S
mAQ5w2ALKuIIIzobr2qps2YM7Gr2ee2KbFICLN7VPrjEvO07IF8fHfXSlv1muTMg7vSLuCP1NdM0
u6DJe4FZRDL1NVZuCgaPrMHm9xMamjTRm0UHVknxCuwxOQxfUDgNRmRl0ytNMuVyzIhhDRkcbXst
D8n6qZiz2L3R/bVg55n/P5xmx1dX9WytTk5lIMDSInUARlxgYZPayeo1+wuavAzxoYoD9oYG2USZ
3uQBNzyf/g2x3twS21HQsOsZN6AkyoA88n56v23MNBFsoSu0X8xuWo3Qh9Z2d5QUzKLvxbzzBuzB
Z4fUqiejkGIE+PbKDyhCb5kvgnha1+QpVjevrs9q0rlGaYBY2ahf5D58VgWs+hnuiw2Yz2xQLzhF
1rIZN0RItOl/RiwFhiFhwhUyMNaIOYQeyU8sctfYyRYNmFM3KVwhQp3Jy7pbmUDGLAjhvLRowniy
qBmlCwwMVL9zERTQGm3dHwg6mzQYgGksijaBYRRFwf/8TOf6UXWtItKA7Ay7UmXcyO+4reO2fhGP
pP2ho258u66jDqj3eEmdQg+mKNwncnsLVzTk/f5sZjNcbaW5z9ZKeNu3SxldL02gN0F6JP08JUF7
EPrAlDGSZRLx1VQZG4axEmEsPVFvlFqbdzmXZOBCY7kdZ27i8pHvHSI/EMNlVD06pBw19TZwQDxM
MQVR76LH26n90dh+S2EhiVvGfxbYu5DJMRLlaTOrKQiIwqyhddxdlJswKIVNvxhizvdPfxd21cji
WYsDVa1MF8gjV7fe3T/8kcrRnJ2lk0V19Y8Jq4FGmpXbv0iUrwozhNqaiXHSCu2BDLtIsCaqFc4r
P1v4T1bDdtKlcoDUsgcAnGtj+05qvbSPVQMQwflaFkASszRZCiNT6sBHarol+D90vVMTM4ctu7F4
0l6dtdfXsXaE4MPBwwmkTzJSOICKg4rD9KqrIXP1UjF6khBJfZEgmmH8WF+JbJQ0ict9s0aJXNIz
vcFPkFtbocI0Clf+8pfjeUdaIXBPhrsWDzp0x5yBo+EW4X9Edheh/bS5ASLz4rgAIrgJMoaV3e1I
nvTT5MZ3tiAM+8F1EFGSL4OY1TbZbLF7GfO9F4byL9hSk6ACnyPjTvSqi+QNulmu357d4/SfRmb4
90p4Onw4t9i9oIMWh6/zRjomSz53MlLWD89U8uQg/TmN7/jwARy/3FxNt/IGnSKBEOiRM2YUg6hr
EVt/GkeFoXaWs2ZfHqu/NzVPobaRP3K1VVNLPChvaJ4hp+V4y/2rNS+wYVDJ6S5bX7dMjQSzvR42
WeDXjv8TcEht2AbWpp6HD2Wcao1I9/fu1USk+WuTIhLRsa87ndvsg8+rWlT8y2tYHer/TRy/H1D6
JosEkJADZ15gfuyfVmru9saluXDRE3xkJLMZsiozHHIBRMvqW1tIZvTbvCEqgUGVt+LP7jFe9+OA
oG31+465K5lFEwutFaS6X3bo6du9pTQjL9L8F+KZGCFZpsew1VCMWLeTEJDlrS1wptrpnMjwchwo
AxEcuVWVrYrCH/gG6uqmk/Y4hRC9b9mMt3R72yok87yzZxWpIDZYKIl7IYqiEAeejAsS7N8pgHus
WMHW2RiqIDsW9klAI1Cynb9yVDnKC/yJ7+oN8xVozTmVx2mm4x5XlbkjxSEGhZzNNKRQzHZ99E/0
qwf+Z9oPAmnUlkqHa5gke5yP66cBmFvMC6HmUvUcg+IF/5Qw6tWw9usjWcF88HLXpVjuWYp57GCJ
rnqdEJcZhf/QjaJvsaf73RW7Kmw9XpSI2u5r4rbcm6vkI9M4sQv9VKuWabCUzxw40wjF3pfyNO3+
8RpRfpX+mj6XmWQXaomSjJYc/5cEauBT1WM4NKTdOM8qRVixNgolLJTzFuTT91B/zX5TeOkr7YhM
jzXsvRaB6SmkNeHgPVkoyUp+8HEiIIbk23XO8DpT5NF75auODDpIzqcfgO/sBIREt34uJ35dWWOx
gY7mFKtUD5qZLBlXoxLwwgMntmV+OHpNSIGQAwyIaIm1USJo5mUXDTltER+fTYX8W3EPZI6+UmrF
fuzSL6WzDM2AfeYS88StUpZUBrmPSMVTe8chk0px126bGmmzEXchkKcXO2O8X7pSqo74CPV2SCpz
zGIQgkVZC0t6M5P8LBxCLTL/biZ5qgLE9II+90gY5ssBCTruW4NcSBV9YwwHhd+rwqwXqDCeAaJd
LGQ//0UJimlrZnH97DTVOq6baLRLPlZ0kcV2xxkXUA2oaTB+RzzVpCrlNsv1tuRQkgR8W8+0h3Mx
ATj4QjvI81b4l/zlhYCTTxx7srXs5Fzj53C6+w8SKFEdf89Sf89eo2+fYhUXULiokby3v+3fZP7o
y7xtFRfZ87EBSjCCEz7JMTOMS6VDtSdF69nMG67vJ19zcmH0QnIOYgOs5wLGFHEZLypQcmeuJc2U
xouC/DUhFWUgCaMKdOGGZ+MNzqFolEmaFE2oMmy+/2cezW6NEDH2sQqRujdw300g75Gq13T1Jgc8
u5G8DFa2nMEh5Q9Ao1GCF2l00BGpeGQGSUjlk6xps/5SGnQ/mcv7z1tlnlug69967QTv7HfCCUsm
vtWMATV6AZX3QK9fwaXiSe2ueZ+IlxZqYXI4iTPuJGmvtS6Fu4QDqpn3Nefq92YP5mHePItAwscJ
CYcetUbrsi/aOY1Xj6MoqsJzVbcRhVHXnouKUuPS+szIbLNO62bf7L1Zb92ge9ob5nCjgrsNYQbv
n/q5XLMOJ4MkiVko9Ag21uc2yWmdRZzQcl7rveS2efZp3DPDL0Vj3B/pH1ScDpKvuPXU5DuzQpL/
sDcVsoGy0Qg4aM30cBTp9O3qdXWCkLo1ckY8jpyBv9F/zu/50g0u/6gcOBNLC7RlQdSg5rzJlxfC
xgEnb+OkifIIGbBSqjYZhDjGehjk7BwgW5DnlDKOcRotPPpAs1y03azlijR4vPczT4ekHJpKGy2t
O15B3ff8sNBa1y4ENlby+mYJrLntplrthqOy2EN1lJ23MeJXGKA5lgrTHc5oVmzH2p3GL3iJv7cq
iZHK9x+vIZn0O4PxxSCjoy2R6vAKIMmmZEhKXQT0Tm3Vzvuz2SGIxzd4DrraV87kuteF4dl2xQPY
fSq2j9da7MxDhAynYNwgFoVkw8O0c1fY8gu891ITuQ2EVFF7uYcfQPucCuz7UErR/z1NW3l2qcRg
0sZwcYrl+phpo+XmImDsS+qMCTaITS3UdLwjoY3NJ0ku/azvqNeUA/6PWLn5llBsGCf3hV6B8Nju
xuo3kfXTGxp0qxXOV0Pgg9zhVerw+fUYvvo4K/u/W+aq0dcZ+f9giLe9RP41AMvLMTZfsduRCu4w
z1zJUaidroVbeJpvRdk+vNjwgMyYOhvzLmTwQ2pTwOT3SElB/eGrzHu5rsFzePVNs0PpeXOpjOoF
7zKQhw7qmox/5Ug/ix56MSouM0CReb0rNoJ9HGNuASa560sb2DT5hbJm219JfHtDVkt/pq0NYd8b
UGeMOiPj3imFyGnHz1CCEzKMpAdwTYdXKwF1zEuE29Ed7/UR9A1s3/7nbE3BPzSP+xtDN9xhm4pD
2sMmlWNB3T0JkHZ67YeDLXMVdV8Vo8mIckplWrCO1CI+HaxBGp6ZeNmrU0MvuI3ugNcEhw078glY
zYZMsMoSpvy4IXd3xN1GplNXtMtHzdmFYtWbn294SPUbA3cezEaGAHwt+dmbQINoMGiY89qrZEch
F8sccWnspO0erJNMPj/i+wUII9ePoYaZNfXHQePgDjcSoSNK85IsuKUBdUv60+9tZFpi78oOnGXQ
NLDtDkrChxIjO6foWPFBNTN8dNUOwJ0Wln0CqJ3+1pMb3A9jxu7uvxjYu9Eq4tRpU5Tc5O/gdB/B
fcs5sJMSMii815lPc8oVqgaVyqSE6gxi89w9XI7iuyX41ckpXzdOZkQV1W2RO2eZZC1qElKazQ7e
ReUgj793RQoFDuP+WcjBzx9iOhkk5ZvycjSf8dsoIit0vi59Hdhaf9RLaLv/XJYkPyAzp5JkaqFO
CgKsLiJ8mzVjcmv0S6AYzjF5ZjjFkK6c7/RG/HtAm+ksptvOqFsPuWe/NLKASsSaD82dfJ05DbWh
Ht16ybSOHRWAn2gBUVTfnWMYrvHNgMqm5Esjyyzw8h21gtfaz5FL9RsGMEz2uBzjzyjPJmxcO4y+
gGItCJ/h4bBTTnboQsrL5fdwqxAJEcNE2CC71mh89tnwnMLWQ3EuiWAgvLmeyUIgA727m+ngBheG
yF/XJgkwhwSIxu/JFOihxl14QcsQRG6ODMmwcsHUR0j08SY9fw6Tb/lcc6jpoaEvMofuREZ3zjfd
OeAEGxskd7iYCkui5DLmKx3TkOA0zop8yznXlyLCCZbw2yWJpBf9lxQkahOLocmFQMQTfM8qmzmw
4txX/RfB8NXosSlhClAzBr8eFs/LUh3bvhBdhl5KpKgaFVla+dDdz59wyUuCzy1wxE+t0D3UNSbh
TCgdUJI6kDWV1iVSqnIao05VAHQ9ntJUCmAAVvyuA+GBWYZgUC4Tck5t2WHMIP4jaT/azYDRe1Ao
uaaqCsk/R9wO8kdCi10uoTfmV9KugDL4iikmgGzva1JLIpcmliz89FEAqiO5lBY5MWVTyE3HSfo8
4U8ou/GI4AXT0gi1gt/vvOr9S5P/yS+xpODRPrLQP9p8iL8hMmc5zoxs80+E/gQxs1WbYiQ/WvN6
J1cxpUWJ+Lq3RmnaAkBKUtYWBaMgm0NsrmnbA7tA7Fj06m7Vge316w111hLsJRepbNZjxMNH8+s6
sd5n7Gzw0mQ2pglmgU7UZ04SBJ1B0MhPv5ZRcoF67rugsSKjVrZlyvKr8113KOO2m7ca4E3wxBRO
iOShEnMIfUcCgwHqyyfu2mes7QDgfDg4sfHqDZGYd17DYcOPUK0Zo8S3IK/zn+ESQOs7I37VNNbf
PoPH1sM6HF9lKglwSUPtz0aVvFMPKlYs1Z4L71F39AaE0UajYBWMK5DgVDBIQNr5yy2ZvcKgWXBH
VYkrD4BhQnQnGhdZ6LwlDRBRG2ok/dnIEcoUiQxpK0vSHIg0KTpUOC6JT5WHuW3jl3eXwqX/qemb
zi+KcmVhFxYXC48LMD8NnL0l83++8TBOtdBr1lOLJDs07pbZPvRaNGOA/P8gBRWq1jGQhDHS1Ke9
GikP8y3HfuLz7vEwVhPl7pjERPWL2GUXOaI57yitWd+D0jHyr0hZ/GrqAru6BUEtEgKE6Qe2WGhu
OBUEJgZ2v8XnQhblZUF16IWKnrnXTCAfj1dR1lrj+bxesnHLQsq8nbouLXxYkoDnpNA+k330JEvL
sO0071xurlh0dSDqqJu8kI4Q1tcHo77fYLSne38PNXJNanQ2Un2SdCVZpNp28lysm1FtrQNWgz6P
iF+9K2eoY40X3Czz+RTRERhqPJzzIWhlWDyfv76PoISdUSGxHGQneJWyuhJBj6FcIu7BvYmIHPXp
RxCmsgQGZob7N97rtvGkdg9FC8hS7xwqjiM1/P2lE7eZITNqyJNsqDdQrIDYfpPpWehExmNVL9cz
sLc7V4iTiYZRqy/HmG1pKDLRoWct0u7iB8/gdi/LyxRx2N9hDc9eLNjJbRGSrUEA0vCGbkaKrXRy
npF1pjQwLPT/7gPpWFmm5pCOh/A/GF+BqQ/8JsQ+YlTnHturxOnEEwYEi+3G+RRdA8l0o6IMB20+
luLpiR/O1yBlyIK5jphWmeKQ3jtXurcIyQfZ5dnvRzI0loBYbD2S0HH2b59RnuexX6FWtXUrPHYl
I31/K4Pe1wW6N8QTfSakEV4w0fFo6TZiHzX6YGkinA64rP/20ht+eqOPBbX0O9fdCIAkqV+1uGXu
HTspn9vOa35BlzBJSjeWqrEx+IlCvgeik/iHEcdkOARay8nNpnd9/FTpTb9xipStUCPpTJ5JzkeE
uakRF0oCRgqjCUN5gOXYuD4LBYBRarPJEg+00iriS6gaj7aXhGb2y+G46IvxaFw4uKtwnTjePNkB
xQx4W/IjABZq2D76Uov8dJrHBsU2yLYxj7fIe/cPArXgtB3YLQdQu6TJ4EzANnnBPTlz2VWv6A+R
8KlhS3X4jSCtE8wBY5r/dJ/NTt//L7yXLRmYdRgid4yvAMBh4RThGzZojv1JeFxu/s2pAtzXmzHJ
XfMQt0mz+b0wl0Qc7AO9TCBsyd42M2Aq6JJLJPIflKxFAtRJ97AtB2HK5vLkcNu8wKNO4hpQWjiR
1p2XpJjO5bxioRcHi4+2Tn4UFiJ1fSZJ7NQ7OtgWWBNliYQ2CpM0EvIP5QJOtLvQFciNLix77hfV
dcqAxtLXSy1W8qjQNQ3LLzEoSfwvH2Btd3Qwzuq1Hf2v1MhYolAl0op5jErT5ipoVjkeEvQkgu78
Q/EQ/BPsFAX03Vbe9ocefpXcRFx9XJ3LKb7Ix1AdoQRZKEnU+BcJhWqF8aOPYsJMZyvU9U0E9ozx
yZDbcc0xnLhAc5oGokn6s5Bso4V5m+YHme3Ugcaymd9zHEiowY7Aa/4u7yZUcrB2dKSrM1g9VR8D
DTHwHeKDKiKMSIkb62fu6i9yS5Cq4WOKOvyAV+7a63PvlhoAk/dyylQhXCnMnyBO4nxRgYBj94xp
eDMyr3N0nci3p+WIKy8ypY+zcqk8nwC2UT/71yknCvP6daapEtGWB22hCw5LVeVoomKi1LeysaxI
jYerg4OuIjNJ2spEYoF/KNbogkiaiTaDbvziK1hc+91Ht2ZI2ByojUv7aOevnuZwBA/xmd9dD/Of
PTyONTyYAQOS7alTF9Hz9QoOgSyuXYCx7rDECb0KQ+5QAIkBRKsOQujdwmNx8LlukgwoLmjGqZ5F
Y0H1+6Y2kvXb1niWwYx5P7J50cVz7pI+RpFBb2pCTOF6/dCkyv7z8r9vx8j/nEiYIRoNPopV0lsc
58PIj9lZ2YgRwdTjqzadSXargsTxESpu0UhM1z7TyH7645tyuaA5X2CsLFes1PVh3WEEhVADZi9l
muxZzIgsW6kdnNJrY72li16Em0+cbiJBcesSWgQzoyCmSjsY3xTsMq7JbI/KBZwNGyCphtCvPl9X
xMSfxTnyZXz8ja7TGBYaUi+wRQYd1npxlOaMdPcvx8Wyj0O1A3UZ0YPykDlMyOiYyxKNFuZjcL/9
d/daEuMkWSgLWaPkY5KGZVQvl5omc2CuNBeLoNMwJ4wu1UmaSizG1bYES6rhkbsV11wNCI2NNihv
WdYXSz833f2FGDlYk8rCcUslZ8dvr/OOoEXj05YUz10HznI6pL8aVStNZGQHNaglGFLo7YnCwolf
+2HHK/ghQ1CpIEVa0z/AvDUpVQE7/khJzt+gncQ7IRaY1sGPmwpVgTUhq8nqMKhh8hmVLzEJo3aF
Utv4oDjjM40uU41UCNevpWI9W00+SpcTDFU1rmZ1t/WWzBf9kKQfxZxny6rk8AC1bldX3LjCHTRy
mwKkq7PgJC7C3Jfxmhdc6lfyzZ4jJXWm9qNy5XUT9vyN0gI5QEb9oD5GDOA5pxh8hnCQ7CSti8WN
s7RP4cQs+eAGvZ0LkYYUm3q71ThK/ze55gvxBRwr9vSf5GL0IbOF6nicaZZ2S+ZJcdqvdIw16SH0
gZ9rGnlXXcMLuzso1DEYNckhWBXWtyBPyUnC9u7h1AFmRo49KShdDv7vLF2kEXDDHMAUfZeBh1fD
GdG2tuTu4RTAxfJ2CgRfvmO+kx9OsTG8DOmmGz/ZIYA+A3Qbe4eADWAm1YQYucxuS2wne2EQHOu8
H/cMa378WVDDimcdo5q+dgZzcwCDmfn0EWBirRVo2VcpqCR2rcYlj7DX1sMQj/RpNq6gERRLjP9t
IUJramPbdyT3urt8vD8CoqE2ZqYs6OfSq3lER/+elh7idoYtH2o53KCPcJnJSUGVdPd09bmD+gyL
JNkNqjdbxPVPFT8NojRcaQZ9jGJ3yabuMc1tY38FrKLR64in1bIXdwkwcmPx6yVTmcV/hMiqjNSc
GToe6lwAdHzlFBtQafapfVw5yZFkJMPV7A6qdD5DVfC97pFXMUlBKj9Evt+jlf415aLBXGrga1bb
HXPxhdoXD0aEx93/Dcj4lIeq4hW3GPHxZ4SHINLkAovv2qiel94x9PifaEHEtSJ0x6SzD8U+QAda
J0u70TUh5QLBGRUd33e20w+aMx24k5wF1G/g4m4Xb1SIMKbC6xTjYsu+GeCsutfkrNGGIJ2b84Pc
lGCfgE6OZJPPs2osGRSwkZ7ep0/pMEnojiKsgoVaM8qfU9MALb1MecXTDqls3weeIVAb9kqvdNym
2yFTjXj+Z80DmclpWdVs5+I2hMFHFpiJ5HMXqnWYOQyJQ/NaVKD9pFzo7oao1Ai5HHad47O62/Cf
fbA1FdSnJ4aXwiyAiO9UAOHwQsCDhIrJJeonQpMSAmuSkpFX+HvakUwzvDW9jO5kYNWsKlbIafcP
BSjXlnw/+gt7M5bQzOjDNrri9ZVxyPmCFNn1qECYFdSE4hp1h0d/i/FwHtAFS8V/mGwzONuy87fq
HZAws8Na6x+79zyxy6ggXtLotMC5enWYL9BIxub97AHKkEkfIE89znQux283Iy8GWPRDDjo94J08
oAP8cE3Td+svEhv+4+xWcWP1pXhxW3okyVnJVMi38w3k8BwOloxaeDo0l8z/XaoWBhsj//jzZkGh
OVrjwf40aFwxRiNG1YYedUenST/qfijx+eNc3HbPNmkCp9fNiWPYrOa2bHPY+CDFWTZOenVvwaZ/
jE3DiYL6z6Z40UR41Ty5JxSY4yUEhUISkYxutKOp7xsiv8tJZilv/5h/lSbiKfE+qusTu8fXcZzw
sNkLmoFI6DgmcWDRQ2dqfKHT4SuShl1fMUVjk07vbb4C/t8KgEyvkJijuNBqwXVr7VCoNRRpZrh9
7Bh616lL2dbAIpX5gpN2plzSFRVyY40zQgQjP3agVFWCJMvP+P2S2V8fUXwon/7QYmMfNI7FTw+S
Rc5S80iFKDWjB4QLdliLSXcBWGKNvAtEgy7vMbAsAu8y+2iTq0FW3+IA3WAa/PTGTfc6KnPWqEWD
tBlmx30IOge7PZxB89Xk6rTuc/NxPZHGYugowgPoI/T5dXVsCKaMu7xGakTEnJ2uh+AHMzWmFMkx
16Qeh94rnMuHEy8Vcf9K3EhOCoXdgYnCnLbMDuUcpTneOV9u40k3rp+PyMcV2UINIJAyr/qCrdmt
sUPkv4knvldLHpZfxykJcnD+y0VLbUaOs7rCw5BRyP0CgTaZpakhoDCYUU+8CRbVffWCdfNA0rM8
Ntddf0Rh5V3CeFHsn+uOi3hGs34S50D/PTlkcmNGKN+LvmEAGZxg9s418pIBWjyTCCEhsuPI0u/i
vrvWw4IwF9p796sI4d6yzvx7B5k9PGB5WOq9EYknF2B1Nwy1vbRaj6rGzQ+hZDkZgpMLMyoWNIoG
OyoML3LK6MWBYO45vGE3/ZNBXsoml+tKzTk2qcz16TeTDnclxVB0sjMgPYP+QeODLE/QXTNKi8NK
j26mBYTGBNVEOODobrZ8UINJs4VmYSyfktLM/aTKTWTn9urUIRpOJW8V2EKQm0LjHDsNIpL25TXK
Q9F22TGPlxfU4wUJ0Bcf1SO/SALt32hUh5ZHiw922AmUQvtcfVJnasbsC5spqDmqfH8h+TOk/av5
fWtVp5ttI7IIZlDUErcFtsF8lQdDF+McL2d2w30HU1Ws7IoUyWep246S9SffO+QIe3P7Mn2CSFYt
Ywq53FCBV6I0GNdKPjnOgqcfco1ihH+mwkPRw5KAHNOlYVnv6azmRoHQkDG6eH3F06WJE08DxFYf
YeQ6Eik3E3MaXTbcASM5Lom3KR9OS+N8DrdmbAXS9S92T+xhJTJ08LHnBigz+03i5JeFzl2REAoF
vFmkukZkSRNqarT+/Z17TBbO5ScW2c0eijCaG04efvuGasfaYY/Cr7IDypgadg4zONrAhZeWKIRe
GfQTp7kL+DNKJRgMhx4rCjS+Tydq6wz5zKk1qdg7RgsbGxF+caUBlI/AMnDDzo7LxPjoHSy09PgC
2qZdKhKTuz7tSXb5O8OzBI55wgGaw0NoqwCpWSkB2jCnsm4ewbCv44Q08xdi2yb4I7CExnAAPrCE
Ap8vW1I2w3PygXmGCMTCzj4sgyczHFTm1pf6bQoY6BsB1eUX0QgD6ZH/4FwSldYJXwIKRmcwfDEu
StsUyAVSzSsNQZP+7YA/X9aLTlod7UrPMuc+r51lVJPy9SJhWbwfW1EHyyP1oj4nxbDwwarDs4Xd
pce4dxn8f9vx+bUYHHBA5XGE6Yi3e/tmqzFvCfQzduXWLkhoty9SRO1yxTOx91VfS1RXcjp3mvft
wHkS/lLZSUylkpTxsxl528pKcAF3Pt4SK4WfB5Z21IkY4E4qRFDvNTwevfAdC6XL8OrU7TgLYj5U
RbnnRCaEICqrZurLzZI7UlpG7q9OW6cdyqm3cx4cYWDWyp7I1wEH+d6FvKcsKlPNVIbSpGneC0Ds
ffG2fY+oMa0rsi+TjXU6YhVxusTefSd+RQbrHDChZcOYXkoWPleaHBDi0V2kdFmHSgc/Ze9aCJBG
6KR/aPwMJJ1GQroXLDN5uBOwAn2JILKwMbyiBdGxZIlOpL0lG6o8UHqoWlxdeNQuskSrH2jt8o4f
TJToZAl4xVl/pieptpyGFDaQFGNK9GnfZbo7umjcvv+5+cwMszU7SnnqG+o8wwJjJsbJmnYuFwHN
KdLWA9DBuwbnnMIIeDR0PuXYVxt/eOWZUd2jo0HoWTpjTY688O+HHNRHa+gP9at6oM1pUL7S2SA4
sMFo3FdSssDlIWiycgu4Z7255xUb5aOWfOKJSnm0qpsDFitKeE45SPkGgFWE8yOsYFaS4bjkrzfZ
JKYO0gUMMsR3escBfUfQg3NBp/moLY8I31GlDAfRK0JdTFQTSiSdKBSFsLDdW+7GSdwCUCuI4d2G
t7TOre4wKyixNna+s2dXY4sMEksgOrmr2mjKnuVirCF/PVrwyoRCIRlGCpBc3GINNwRp64iRguh4
XQ1nfIh8NPPsF3AyrVUz3O14aE2BCz0ujlG34kI42pw2VbOz+8uAWOx4xtNc+3vgijq2BZK9pPJE
xj6TwoSRT2zD3CVtyZh9p+Pe2N21/EBxLiqLL68dTtT9m7vVPELyUXVeC1ihlRkEinWG1N0gHS5s
rhJZVq7aGAbwbFLe9gKt7BmzEK42yA8an242EODaA+RhjMPazok37jlTxtmBSL4BPZRyYnBryGaV
Q6XxlugR9NPMhQI1MIgOBjaDwDf9MTZtslmv77GFiuVTAHV4oNkpGBhddhghVoUZAlyoD7+CKkLO
69EV5qym9M7f9oH9asPv5jX7D+ejq02pTVJ76aL0MUSUIOWW46lsoD4ddSG7f0xwwZVNGN3JflwD
uqBvzarBM5omcrgDKDtf48Ta3x0ATBenrNapKl989+8ShqR04YdCoidtb6NfvW3Nd1MN5uFEb/mh
NOyLFX44Mf4Bc4ZnfOBDKkewNjoLsmks9cBv3jI64bicqRwccwzqWVP4gxRmkwawLiwmtG6B8kKu
Ce3FfUs1UqD6nRnTGii/lKjBewq1eImt7Er7mYOvAKFH/uTdAn1Prdw/HeLdEMUWQDLkjqiPQ0KX
M5u9vBNnxWNZLcrfjsW+stv8ssg268SGtvUAGqrjl70mAboISnsT+7OB1akVQWPNZCsXfLzuCAR7
FQAYq1V8oMCV/lGvZ4fHYebYGf9cIhKqNCQU+ptVLqWKMW0Aca/M9kbwsjmxilEvygXpUnWdvrvC
pJqr7okRqFNsFtTFyrjUKV3vYEY5ryYWaISmAyig6oT1QsrfcUhUHaf69EphJNWWfwLvidH4/1T9
sqRMOxPA7I8zX/NOfWX8yW4S1rZtpHbrdr31hZMZMS2ZW4HidPlaqFeo8vASWp9TGAPIntlQ3MIt
43vOapX6uUleQhAoWX2FQvIq8+1zE+V1+S3URPdxva/3d6OvYNmqZAG6rs8GpLSfTSO1SzNupXiF
XMTAMadQLinXs1kGl26897oEYMOzoeisobJL8HZZOMq07C1ndgGMSnCbtZksE+EAXHLu2lCnlzim
M5CDibnF1cmEOET+dRtkOHHwqpfRn07BIGSZVzKyXDwzQFs6TgKCjbLlXkxIOpzECWhVrldsga0O
T+BsrHAwaVf4/Ppj7UGQpq0RdBfmUcv4OJIRThjt8vwK20c1FGcYqL8W6DO31syOCx8IRmFUzYan
4C45HW5y8Q4kgLHTUoI5o3qwomRbkNZ3g5NChoaRZGoq87oKG3IFwII0SJMPk4qdVtm09KzitkY2
AgRXCuIhgUP31/SwUbo2M/M2zo+6SSnA/SQbnaJPC68OzF8piaXLRLKUceKjLA/CCRSxpeRJphQc
1lyRFiXn3V49aBX07GgvJ9j/MBRDtj1Q/xO5pzsj6INQ+8l/bFT3LxFCMkkDgHkrAMPDbnDiePbC
bOZtK2Vrw1W3vvc4xYS50NSL64agoNK56X8QM1OhS2C/7JqNkXM6AFlDtbCJ+58GYVBWYJCWRFt9
B2ky8lNvd58eDE6HUoT8JsZ2NdbwFnTld5M7WOYJgrPiw8RPiwoHJs0kAb2n0TPSZAs+OJiIyxHb
0byQ37j+qBHkAE4NTJK2aUPbrpiXVl+HZjdWImrpqC6BDAM+uTpDmSDRf/wjEKDdTAy+djJUs1ba
tE+NmnFCTji9tGbV7h/pI8uPk7iqBggT+khw1vrmsGJgc4xy1HmEoAnmqOkl74lnpcnCQ5qwQzEq
qC3UjZV/fsqzES5BIsHvUew/uAWv+Wgv+wgCJNodrJ9xHHcMquzjfltTfJVrQuNBTSA8HzueOfmT
jsVnxRM6YD9DbTZib65ObssDGBoa5QpEjccI8D/c1+FwKwc3hfrUccO7CFRT2UfpQ7dTFUR+9Awa
ZFPZKW9qTwBYOz8hIutPlNvybO1SfQbU199rfoh/KmRp870Dm49Jqiw1o8i9HGlbWC1HfCOrOFRU
orZHixRFCO/Io6YD+NNj4J/SkYFuO+pzel9Z5t8Dp3mi2vAjxwnkaj9aEwu1kfLt/Mme3qhzqD3s
Q4hV2uuauXcHP33caGnyHIWihxrVCSjUyPanlmcg3uGbo00fBFwPcT5nPX8diI+7iJWVa4bqHT6Z
UGU4EX97qgG5hUYs98AqJd+Gf32Cu9ecEXEQU31y44JvuJRr48wgUdlbET5URzlWfisgQH1YWLG6
DSu3KKyXSu/dQeKhbSDae/jVwhCQDtixSE5myFAgKa8B9RlEXxJfZ4xS0JMHxMF+m3Z9YEvTUYYz
5WfsYjU33SdIQJYVgx3qeCKBdNWfTPeJa6i/brdtDVJML6SuRX5fiLGUFDDwEJk9I+PzA1iaL4a2
JZZjMz5DXXuIV6/LTfbVtvyPO/mUxEXRE/voZ5oDt+iiQBAkeRrR7eygiO0hU8a04hQhXZYB4y+0
emAP423HfgGkhwKmqcqKng3c+Z02HKfiliUGxs9p5DZ2MFonR3ml/eIiZUUkuWHHX2y4S6L+fhi+
dtTUiFPbBf3mz2CnaSnC0YveWv6cZPCj/OSU7SaRTz3QqEqdeffF221f/kUJ1XGLtlcJp7BVrH4D
Xg1FiWG+JglDUEb2L6/MNVPjApb5uPlA5Yfb7VY3Hq7KnlrnbxMMGW0oaKgVmeb0yTqJpuHcxpY4
bEVHjrKfdI+5ZYjuPoQdIdZh98wzIWpuPQQl3QVspD5opyJWcXRqvqVHShMMpSHuOa0lzOLGudXO
iHVmOZE0OzgICrd6nvyys6SmfDA10qD6atebfHiCyJ2PKg418bZWw84o/8ANbN4GZp4+lZUggzBf
+KtGps7zCGt7XOzUWp1wkB23riJPwrjU0jDjqg3bG28Vm9fpm6Yw6autB3x4/qlXyQw5HH5gtuow
jI590VY/E49rIBepdQCTLJk+bCKJjgPrW8Pu8cCU+8dF8kSYlsKC+Y0tibPVgO/KBtXdHLkz48AR
0NqG+9R39bi8E57FmiKhP5VwmUxs/i1cN7XmUUbhJpfA7+PQoSIe+m0YxMuMJE905jEB6GRZeSqy
4i0kKaJyF/uCKmNivdJRUieVONAQF/w7lVZpv4OD0V/ZpaF3DPSMVAqrM0lpuUx6h+EDnlPcx1qF
z5IgW2qCt0wrM3GJRqC29IYzo1ImeWZGPvPxgH20QSv1U9MM5aHTZ1qfU9EEbg2o6vKOEsgBMOmd
9DYCQ8pmYgM/2pakgLUnO6TA/V+fx0Ag68mp+A8OtazhRRWSX2pPPORi/t7XnPrzK5kAWrIbutDv
gXJghry6w+/GtucfbFx5wP0MZL/J4iyhtGUKC2FkvuKHSVX24TldL/8wGvLd/o7MBUHk9AI+tbw7
CPWR0lwtbMny/w2MNniNghatMpRkmxHewSRCjAmzlKQOAGu5vgl9OSqgytodGx1rOpl+E3GttxBu
qJl1g02QpnfNnrG9JrVzAm7//zIHQmxlhGzvAjfigb37WM8Fn807LdRKEVsRn7qUZAuyF+TpbSCn
MklG2NV33SpuSQfSSAqaEjG2GMCLMDh9b3dsy6PzYzwcd1JNoUWAzxURcO4wosuQD5lP2WidFu5B
+FPRVKe4HsGiLNV2eC/ZH1cPTiANkvxEeHD/+ZGq8KK1je75RvsHb776G6+l9pjEpNryd4pGzJ19
QWlSGR4zOICIOG7++jgk7YgfE0bhij7DIOrxRV5fFTC9wxHXPK5ayEqVQzWJ+65FmXimE/nNBhT8
ojeSOKbjAphQ6B/MVbmSzAyJ6tu+BiWwwdBUIuPqcC4rao66jdaagP1rtGwAdx02j/uANM93gx06
TdVLprc136oY3SqVrP2vNqkdGQVxHrgXktQPOorMvx+pJ6SQTtPHu1utWNRnsyqtcmocy6E2siiK
sZvhJ+Yqnii4sN0kaqPfdUgtA6nt+fch6NyjP1HAUNllmzEikBVTt5FTJhmQg2ZzpP+zMJWYl+t6
/cstPRTa59TtEDHg55+LqRDcbCz38FCLPkUtJ84SaSdx5zhYlmYGZGCFPAwSolznlnY+iKU+Gf0l
5FYGMWdOaNdhHyqUTxjTya4FTsc84pUGEbadCD+0+/Rzs9Cl8MqS9NJ18ZnNY2a2u2A1yFi2Bpjj
mZLuOkuKZm4hrsWKurczckub6aShXxBeNYYeazvp5fT621CTICZ7uavSOhuKog1LSk17u+Pgp4L4
eecAdHN1+T1OrU1bfMm7k0K6vvPq3l7c9CACsdVIiSLu3fr1H+0lGeF5B+3kNXPcpDW3Z2g4pwIB
7bg9xnF5T18VkdSlmqyrmvc0Cmbz0Es8J7uo28ETxU9rzMyihEBEj4iTKyC3MoBmC/2/TbIqmlWq
CaYg0cTHYFInNYC5izq6j+8EcbKu1bVx33cXPoHwQuBqif/phdKL7qEEXlfGWF6/+1RuZL+LElGl
uO9Ny1nQRtH6IqLVocqfr/mvG1vuIgJify4m2dW7xSQ7oiQYSGCCSEMmJ6w3mLbuu7+g+DLsFPtx
MUJg8hD1pyz2FNVYAi5F3P6Do9oIO2lGcas3bbGP1EB3cKC4TKpID909ymmGx6AyxkdpCOtExozE
D++wnRTKmrJbvyUtPz8s7J13X1P/UegRyvhBjvOxef6vlh+A/ClOTxKSm0rOzVPRLb0UiYKy7qh+
HTzR73Rot9bxXYE58rYPbbIEBg1YdbFeV6cBaGdLsBbAH1JR7vXxeUmxJKNYjrhhGcTClqa6lDXG
cV+RXJV7xuCUzLLNjuFgtLRJGWIBrBdLU0y+LM+C4B8FFvinqsVQ2hkSc3gXIeJVnGbHvnxmLD0M
tDDuZqqeHDiBQFlFUj7hdZ4yHw+sRSHKkXbDqM0h0HK2HXCO3HK/TY3XXsF2upY+9Mno3lO6ClAI
pEgV6hq5MXcGC/90/22Dh/lvcMSu4O3vJBDy4aORwwm43MdzXSPWBs7ahtFOoW1071JaZLS8Zx0z
3ZyJUf2aS1whRwrR4m3E4W9RWDmqZzTwYz8hVc/NORaFb5MHVhjH3uIFN0MS7MrtEgTdgKjpbkoJ
avL/Cb85Py55/aNBqz2WQdPKFnkc+Yz1mxkJuhM1mZf8gU9UAltlvIc8fGXglowizqhZ8PNLtVAJ
+wBNbmM3RriANuXkwfDgNzbLbKIPIgroDw6FS1ZMXSD14Oiw9kHfSKd9ErBENsYbRoU57JSoQEgn
m19JXzlJa9hwADU8Lb13TnLqXmE8fiJzmjcMw33NrMn7JZIyNrTbzTFSACZ5H2cPYKimC0N++b9v
0LdHWmeR6WyUC77AkLNupoGxxmZ+yYGtvcbkQCEPEAJ8JQUEY7wL0blPYtUChoCGXmpUwv8j2XuW
3fayWpA5De5iP2urp+k17y1dxOTF5/2PAiM6enu89J07dE1tn7bBac35RxJW9p0Ec9QazLYOwEBe
iEuU8QaEke0X5sL7OeX6aUkxfHEaBpTCURTWUbVoNU09o6xBGfg43QoL6wih9Ocqq7DhsvxdWtqP
PjNnR9s52RDSqp2ry4PdvuM+ZQIDAHkEAL5cVintceFnSzxxMsep9JMpfbEnZjzpFD5kQ9iPKRr0
90mB+0Hf7GRV1Q1V6IsghXc5nq4yUnXvhxauXuzKZBkblHKRMHLAoHhmzYGBfM7mU5tpFi85qQ+I
eHnpOHXyWYP7cG3Pww7frkE1dZCC3ccYtES4jfI8QLwwcVIa74Kpzy1Y6G90Koaz9gLJDWBYhXv+
vs/BOq4XwQoJDEePL0zNwUxuUS7lcwuLx72AD9LXyO/uznsUd9YPpAFph5w1oUiWqk/YAn8x9UiF
gxcjHNaLFzW59AKycBHeU9ujOuKSNEwSBZLBXQgR8fHTchNhhBDjBIIfzjMDCtKrFSIqfUr9og3t
QKx0OgESHyS+wOE9xmnfs0x216WZEH9EZd67AyHsAqfSLOcPli57LskJpkqp7fJTTXULvA8C83Re
/gZt77X8R9PPMbe/qa9ABwAecGe9GJDA+11Eyx3+wn6lidY39I/ado3WEfh/euSe1DM2qZv/TGp4
ciQ0X1aN67Lm6MepEeCar+vKNSEJG8bGepRwq57FWL4sfO1a44x4zZgeERg/TBZtHQuIDB9vEuv5
XVi7NhS+/9KXY8hJK+1XkcqboA+5eeGpdm0IXknFSWgg2FvrJbwDWyHzbYuAJ2lWl/C0TKSvPle+
3Pj6YpMnkT97CQO4pKnftpBq+IhtdzdUO5ZJvx7qYGc2ffUbDTYXOJWiUGCSQcMg+A8PDxUnEctn
aBgqPlF7MnOL4cX7bRnOuSCGIlEyXaW/q9FNBdX/4k92L3VMpWQu3XGs2UQyjPQUf77PsBEw629u
p+4y0ioGUZF7AFjziZvDIyJZtOoVaMzffq2SPZjSOhFKRc/zY8d7QcExg9L7YZ2iONykNrs8hs3S
zJUpCTNGsfZxT5OezZHcF7ScnitnxxG8xaxBI2PFuHym8PMS/nHhIVx24EQ5s8gM45hP9QiSGndI
Tgyj5exHs8B5Je81SWYhJMyB9SERangWNcm9bCygTB9oJtpEFzD3eaz+hBCIttClsmHywOcanS3P
MOZatbxpyOvUdqKEDmHjz5svmnLnx9WGZflMnchf9XaSmow/Nrg4aRs2XNecqGSvfQKCvUli9Qr4
8xlo4JfD37ImWnvmplVU3/SQ7LvA2ps5F0nYDjEzLL4h2S9mVLayk21XoNSAfDpUOWNBMnzMIe/W
XawTa3BYZ0Ymbxju7b5Q1lChp7hVtwpDd75xWsxACqSXQZbspapiNJmUEmu7IslKqmHQoDYhSftX
/5Xgs4hIA54Fa2VuUqB/LM6X4PFsrPyq2Z2wz/LRLM87eiaL7xOEszVvpgdQ7sylaUiGxly+jkEE
U3BuHz40TVKUAFKm8SBWD8QavZLAbUxiPL/TDCWvo/XeSF+6QolSQ8yVl1hncPNfP144awHknuZz
Qr+cH0OSDfqVQXQvcFOPWLrX7cqaBWB8kQNKWisLIANBhWThlnJUBO1goSgMfotSVxUfqGqrJc5k
7+0UlqIE4187zAFLXlb7BMAFLY5qEIlFslPZNBlUPNFNqvwg1Bet3bOMwJaSvYTxj/wid0PEd0N1
2PCuEjXG+L6+udH69zkKlCii01BNjKpa4BkKHkXYzWJnmTMEjI+xlb9zkMuhnDGuDN2bvxxsgnj7
7b05wCHEmA1Kn/1mXRshiKdAzr5xdJXMGEq+TbeH63ngT7SGJea/gNu1j/1iw4Fq0d1URHjo5Gxk
p5+hpumsrfITLfAfdtTNKCKNPiUOW8bNPjVZWzkLOBls+ffjIJhOwlgdHLoFsIbLrsJhixnzq6pW
6u21OGKHeX6lnD0JCe9W/lFoovO2xdsX+rj3ul6dl4afYRMTRwmlYhLzVfW0p+rhCjrOI6TFz/8u
sWPhCE1O9mDiBMkj06VQBqBU0w3ZVEII67LrmpZhFq9JS31V4ZM96BWg3nR6xL59W9A1ABXd+QLc
yM/ZRVpbOq7nIRNHvNVW6JfNCfZe/0PskHkddrzwyyDo9+LFFjgv65YGoBxCy4Fb7U4xk0Xi3f3S
/9cweFMgSFaUad8uH+mjHrHC/GDVa5HTOj2u6TCx2vzPGi94u9Bp9jozcPvo6GuyHoWPcy/cvNEp
AxDQCLKohP0P8E1bq0eDo7UeQdn4FTHjytqCVN5MeYtu/sgvGLoA3rQsxCCaNlZi+Qb9ul0b2VUg
XWJb8BcpXbxqsWZuCms7xLXSkA96CGQR0L5Wb0m/IhKVZbV5evNrHAIqpPZ92kBdIFKLvzfHoIDQ
TO8mSSL33fPmlaulUMaFd0z5mLaEEAMZxxeiVjeFdrIaOQwVbDAJ0ypSyn1fbNsmgG+gKZ+I/1Px
fnizdhMxe7hAwe8T6/l66ywd9st56B1twdiwkF2U4hc+4bN3Rf4gtN886WGqY7YQ1b9RKouD4l7u
Ewur/bdTf4ngzG2uc1VkCjBGHfLjhKjp3aQZda0Z0PI4t3XyaytaesaJ9++AUbsd78YPpVwLkQaK
YWGu1onOfKtyzE2RfuF5RTX3E3jshfFHyjn3Zi8Orvm0cQNBP9wMdtBtbg9o11mhKwGaPSZaTM+7
rBpvvCHYw8ZraMwCFeObGeQECPop0TmAklfsz8Xi/ok+nS+LOIhHf0wFH6RXJeedqqN9OieFJYZg
lcX7t0uEX5PE1chTvtLZCAS30Chinj3cDtuSW7I2aj6na35p8lgCXYr8t9i6ShSUTi9K5t6bnzUq
Sa5hrNb/29cld4t9McS4knNQRQA83ezLj+QhmWIR2m6eaPNRyGwz8QpJHT5lqId1HXXZ4j278Nva
2Daatkuf11KEZgFnA83xuGNO+JucHPkmFCwtLz7DueBJPsAN6YtVptwqgHCgrru98IkaXDbkeDH8
pEWTqPDoWoocCQSx34t6okN5+siZodqo/GQtANGWpkk9K+NUAItTi1z6S4B24xQp5vzwjp+CvfAr
UUlgv4nU8tHUQgscJpQgbPVViy7WP/kl57U4KawEnVgCO0kC31leWdCD0A3WQkBLEbhxw4aISonQ
0+R/mhHXzpWX8TrYXw1BH1R9aFpR8Qbinmye8HReKlo6Nuvrzu5EkDcw6jLZ6YaisnhjIbasxn8T
Q6XIgWpy7IDH4Xx5lhBoJnyaObjvgmQ790xKlEcF8WPRvOkBRXNGiDhQ4UJlJlpVX/to/U8zKHsv
gg15QwEWGMxJiIkQZkN/3kcLErWnFfcSp0AcjF44foy3zKcv6T68yd6Zrfo0AnCAmdBKSiqxvFsU
J4bdrx/WSxb4wyrK7gVRtmfQvMztOfFRaUsLSxthiTnPCVSRWsqk5TcxuUybUegoB4wK4QRWQPBK
Z/bvXGs7wRk6pzZ8ixLeleo+dDFEEpwEGia9SuwG3LkaYtalaL/wqdG72CLmFs8mAuC7yScP7IPm
wRK4FjWDr5EPD7bxFRqjVwvAZ7jqDoH6U4V9QuhSflO6wjcbM6TtQ15t5Ajjq7US9f0KmVqsNl3h
UAuH43HSEGBmyeLqCHYAP4BcnfnDFf9nogn9Q+rQDf7ICJTHdfUQqs4fNr5JGr4fcktMmaU8YALp
Nn3Hm/oyYj6donhhXLiOymggfpBgFqNHIhYRUzctxrG7uWDJYO2R5uN3jAGg+sUZgpbjo30xfEAY
J++O41ooHtwKLidlzA3Q1sY69lGSjr7wVGjhO3B4EN7HR0ZODOUFujBzW5KqLpfHQFI+tVlBbAlg
lvhsaofgUjO2kG8QJnV7HVn1Nn5cpHt3PrXNDRz28ShxERlMvTzeOPbdQKTN+LgcFKG7ulUGvXNA
NrL61kqi8lippJFclYhWNwCNNIBZ13BOntuvvUEMh79fe6643EwsLGkj+aaBpfYJjbe2/kSDkrTo
+zBFwsgSwKaCF+/PbAcFkwtp4Tu5MX1MEdiP37Gq6sswPk85QrGAoXyz21/3dA/RSHa1YdzybXLF
ZPKX7kRbY63V7HBkKeiVdLN3a12g4yKshWzduFGil1RVh0o/x/0up9UL+D7NkFmINh91/hWSkTvj
z6hE8/8Z6SX3cxsybdrx/JmxeKTZ1WLS3R3r5xbWhgB88iZ4g4fwcwD67guBCeY7Nc4TgGKI7lYD
cuLnvnSoI+f++KiYImv5kjhUoJGssaaqf1GCWn7xGR3gcd8/MId9UmaTFXq+KhE0rgXZOY2qMj1R
HOPTsKQ0l/TNq8f9R6XEfBHpwmElbi3WeVgG68uOY3olDldafplZsFC8Q0B9msKGdYqQK236nKxj
vYXZTS45k1OMJ8ICt1uufq5dvoWQ0SFKrj4LD1qCGxubkDl07yInoJmkDx56EKEJZmIYM8tRx83n
0bj/cHpl/sFDv4NhYHImb21JHtL90rLgWJIou7hLnqnPGkWHPtJSIAvuFw1KiAw0SQ93QI6BOMUC
sUc67KwsiJUwN7Cyw8Q/LGSdcTpRMR6Tgpve3QPA0fxrdvSs+div9zqQpujquT+RzxSnkrG/nvnp
Y5ZSQwebTywHeCCt/TAm2IjY5zAI0TOORtLnLZqbkQx6SyKeneO9OpC7CHGk5SMP6PWHVj5gm4Ti
sqV5NvxHgrx2iTg13O48JvpTiGMu3dHbua1sgdpeTTL3IX250AZ+omE0aEjB4xU2pvCluRgW+4zG
IWywbRe1GxSDL8B29/obEIXqeWBUku3tEJG7gJhgNX3tz5x/NVbiF6ZSiHINMUdfuCAvHYDbmOuv
mE+NcjkCPjJOR0iD28tHudEDt8Edkd6PGmekSJVau2G23ULvGrrGoUP16HzlB30btYVfnfKeD34i
zS3QBIVyLJBpvS9PdRGpodHhnS7jns7rVU+OJi/iIxiHdGLvKplEYHrqWGRukcGS7bLKqkB1Rh0G
gs00oZh0vPj8nsk8v41BvSS9Y0F6eLBYrPXxoXpleqLE5lowGLwhVrUvyRhyQUg3zFfW8VGU7ATZ
8II2NV+741KqyVLGmcipoCzvSuIgJ1Yog1crqkdbGcuAJVNI4wvXC8WPdoaTJzsddpgZlJp2Wg43
VKE0a0+htPPtMIM7C1eSSEX37lBuc8e8YblHig/8Kv0I3kNa1O27lxzrlj/kblkffFAFiskUzKDI
Kh/dGhgm/OsIw7to1GXuCO4e4+rjv2EE0fkyFpWpw6eymFZPcEFPz9hI+OcpirNwDONTAsRoWLPT
yZIGXRgBxtDLh9wkfcIuMMZ/F2VVKGFbhsKSED3mmvPlW3D7cvbfso7MMxRLfAsWCKTYk+JoLuCH
as5U9EtLeyw8kuy1+ZQ1MngLAwxO57t22s0qEJEKvHktnxQ1cArtbHJEoeA95cz+Fqg+9azZz8Qz
8XYetjB7vSQAe52pZf9ZT9ijYzEfcY1I40s8avzzQt8seBMyXJXueTJbFOSJcbS71ZdLj5CYmTND
KTWLn+FH+yBNzs9BYYRFZ6nOqilAHMGDaUb0ulp61wQWZrexAs0nQHYYKTc00bqcXnHGPV4yuugo
wcRC3EXJAMdrKZp6dKt/ZgHhca9jVrU6QgpkZcx8QPyhmx1E5wW4Vqd+m8qTp2obvkCzW94GesNu
KKZUc93dDVNYgdTqVLou+0kJEDtTkwNjeraeNixo5vHKs3KwrRFl2/WECdR5d3T8jyH4YJm1rDBF
wf+y9PgzlOmfPogk4UmzMkbOREi13hs77ZjzyqwZkrWWm81ETehuY4febYz4JvRf7wQKN8Jv2uvz
dRDbKdop03bQGGHQQEaEf2Ovjs/DzyjabOEp4ZDdLs/+Gbk1BnUPTu9AFWHgpl2RhumpdaWqffDa
ALhmjA/tIB7rlbMQMbuj8F0IuFFOBo5XWFFFX8aiQIvVrAXyIFQkvg5auXrzRXamIuE3son3feh1
jcH/qVs1Vg2BD8rGj8MJ5Wbi5LC33j4nly4iyaB0psGeBaLpgR/QxWbbe0eOzy7vBduJRDz5ZalO
TLht0/42uDmow/L5V+oHRyAOCW2W2XaxyDvLIhPjzYDuUP3V/oChRETOEJpSMuexhbqZqy2YYsk4
lwRe3TH/cMayhYTlHC9uNHQjrmYgREuf+nlfMenfs/0mfrK8u7DmBi1O+IfY8dClDLyFMf5lxwgD
1k+EM/SfIeAiZXOg2OAi+oyyIdMKzMuphPeudoPbowAydyXq+L/V1W/t0sbLLgxnuTdEY+xHDQnq
CchTOdTbbHsTnAGoaag3zcFnorNfkMjviLUNQ8yvI7jelZNHkX7NA2usP+eAE9OEQRW1XrT+lHEz
3XtDH+MBfnhEo41bcInhQKzIjDyWFrv0N4atbe5Nyo92Mu3vwqXsxZAyKtMaqqg9Mef7h1colCAW
MZ1OmlxrCDaknnKw5QLUyKFFwwQY+eiEZ+R6TPGRsEbKIZqLfGzZzrHiniKfH0W/MUg7AUZQh9Pb
sd0ef/60/A9y+EfavIlqhBTjjXk5OUJsAUju+OcfRwlpNCvFshU3U7FXv9yjF/odTd/MAt0KcJyg
7VVVpgJAFAsPMUVyAwMdV+3FS3nyjUiqwTSQRrsMfupqg1Y4amtHoA9yQgWJyT2xcbMGn2ugHMLR
bMUPJizmHXkviUMT6JEcq3ZDxYFAzjJqa9p4846+HOS6n+iP2ziBMO0vokSFQF4V3EWQBL/5jvvl
A20ZTDRwgSTCQ42fip4DBXlwId2Jays84QesK7TlzBg6XRO3K+uuIirqPY/Z+ZnzeJYhTFBDI92N
0+bH/i0JBUc3vH8JBUeWw5ZMfmSrfDj8cHm6dtTY4XHxROck9XzXdSML18JbwqMjrxOmHN4ZZObd
r6cq8Xvc/Ad1SjnKG/6rofa0I/i0PxmLS0/UM4cHulsSUyWa+IeDsYDkTvysQAyFhCYnpPmk+9nM
NSNyQz+83AJNosNOWL5WWW6MGwmo7PF8G5XOrRXnPWJjEaaNqVTbYmNU/UiBTeXI6yskOoCoAWv+
cS9wFwdGgb9dugqniDPdNhIqd0Y1cbksB0BNTOZw9yssFt5bkDGsnCO8qm+86zAoUCZQJq72RmdQ
h/BXGDIllX/YVLkvNZmDbc8i16yzL2DVL0dyG/MHFApOmAUMQ8qagaHJwUJlTa1qviitbd/Ryx/P
iansIBubqM7kpPdjgeB7uZn/fJblIpsJLYCYIWorshsR0jK4k+viIlRgEGPTH0wXJ4atqhLDopFO
WlyUfluU2Lb80ZK2tgfzNh2rGjyahi2lyvllUcG5K8FMuEmxwfv+1PnpJVt8Npz/jTYRgNdsz2iA
anytYOdjunEG/1DITZv0YgdKPBwPCp9Gk1e+mCHZ2S1mULa2kGm4FaRsO8dgtuc+opq2HHtt9BMs
qeXUYFl2fDsbjG2TJvTty090SG4V5NjutQkkvpAKYv7QbVE14cpeWlYpQFbcJ4wn9WKH0xa/Pqia
SOFSmItdSMiZaKYtBdYnl2mqX5ze6naqFBTk8GWDhZqGLVPrhb1xlkQIjV7hyMFw7s14Zh/NBXvJ
aVbPyhUTLqhV0W2uKFG96W6OZgn+KEv/gowBNgGwrwysmQEWv4nPiVot7A9BaBWgHaPhDOfvjT6/
6oErWgZusawY6NSBzjkiObf1XuIL3gj/Im1RBdJz6f4/UsP5VeznpoZHiFlNckVaBNk9707y2TXD
Ln8HqvNem0RHZKkC62uDr9Nj7h0SDyJkaPaWcqj4LvhoiHsrHD43ijHvgsEA3e9QbwgBuHG+nGvd
w4hs7uSgz2lsnLs7tS+u2JqS0DsVaYWag6KDXVLSffFJt+fXVS/FA+m7F/7rzSO6K955Hb4jCTsc
zihV6hiECOERtaAJ+T0qWdXyGT1nffHgoexvnbeEg2Ho6EOtACD+12DVi6pc1PBZdae06OOwtVHh
w1RfAgkovwOAvplw/r4fGBymleFk3Xl1qwbWT67QkOPEJoDzdjCr3pj7JDbjqMPcYxed5ZNvOvJm
DC4ZRdI3XjrtBDMjAoTRem7YocIr2oUZljcrkfmG17D5xzOH2B1EF5HIMppvGnTCExYg2opLE1qJ
3fZddpK3mQuuL7T15JMROUcz63utsKICoHj7Nc9ss+6esw69bP17P8uIOw/Elr/vxX+wZseFfGDF
tQUZVHdDA7YicJp+rCs6XGB6XIHY3ZFZziWTFcP872aSkja9u3UEK18AI+U1z7irY0h3UIia5nZ3
03Yaim4KSMHyaLX+kUPot9/m05EZ6agVb2Abjvt2lW7Qq3nniEbwoUHFWnIF4kZziPBhVvESrWej
JTOMZwnzczykZYaGubzDvtNuGE8VpTxeudsak7GS0+TciyrMXfhk7ACopbjbYvZ0a4XaPLik/Xmk
EJf/tL5e0rSHmOccrsCiW42mAEVzO8W5DFNiilA2+An77eFeZC/4EEAc+n1MaZ4hb2/u9Dhol7oU
Suz2+ph0gri3JX38dzpz+DYgLN+uR886pT6Y91f2aDZeeJVyrBqbqnfkJSHTsI3XHcaA7BQMz5Xj
GykmPEw7YLZ5aEyI0FJZX9dAhIHZvuz+HpvDQ5dtEPdiZgUR6n07Pdyq2tMs/rAz2mtrx5eJzIeM
23RZTqMqRCKXejbdOx6yMtCkEYRTiBQnPAOSLh7IHvzHThlsH0aPbmU4vhfDs51Zn32wF/uVmxKG
cdk5g1sP1Q12f8P4tpAmekNlyGYRd2uQNOHtzuXzv3pDOUz4DyihbdeKBPysqQsQGAJWVwC2M/Bq
ERDBAumrX4HQ3BlKCBf2DTmoO14IX4uOdzEHBnPoNaZ0a3b62ICJncg3BdUwlPWig0/6k0Pvht/K
wXihcCoF6du8LkV7TiXFaVXBQtmHcBAHXyC9WkOsGuakj7zBnHLqBEzy5ndejheguhn82M5tPe9P
oH4khFqvq5ClLWA5c06nxol1IQMKADpCp2W785HlB4UFraNIAr42OpPpiZgCAnIylv4hi0lGT93k
TThbAALFjW1uNB9IT6vaBB2HBlMtRtv5/7nHS4ML3DoWstlqcTVpcmvyzoF/alhwzypDaNLfcB0H
hwR+3Dn2N9BOhK+GnoKiP4ziPOdoWKRCQkp41zp4qdCH23u8k4n2i62Bxak7RjwkHMBQwxQkLFgN
c37nps7SIrc+HeV8xA6/SUO0k1qHRYCX6Yu0dePbNGsWUFs5zSSHEX1FrQ+KmFxJ0sfdAzMBdxKW
+pONNWUmxe4OXmSDvKvKq1EUwZIBsqX0/5QehDNnTNUqb1OH9qHnjNUG5sAiMhX7VtIuX5MV1J3g
7YTo8v3MfiEpVKUM75Rcr1soGBr26X7cRLROFe8fSSg8A07HFbICqjCFJORiXFP5YlWTCl+iDQZv
BtM3iL5iy63RKq3+NKCzVtEWf6tcu4ij16+aq03MuXPVxwuYYew0PAHNeWZoHmXcsKw44uKzlhyg
3yLavoeHEbJwN+bGQCR6CITTWFWLFIp54Yc156dEDnNyl5X457SEdpkFxujZQAVK8kjaIzktmyIt
yvJf5qoczK3zEMCHUvDMXr2WG+2BPrhx6io/o0AcWsvGcNljj7ooJPqnVozGo3Ia/FUdJ/nMiBBa
8v36wRwDYJs0O7XsYBJVOaYTer/vi66p0bBZGHXBySIJ+n/rdr4A2V3TXje9aEXjTsvp+dp/fG17
XNECa0ftwvdh7X3/Q5p5+x9DIiqrpZtP4j49zJrizRFvdGe6Uw6M+8SWsz8/iG6NyEU0J6/tyBWW
NfWy2GcDKjX1bgp4WHKhh59eLj8R962JYDYUagfrSasf+IFycNK7lYtyfH5cKkpiNUCjW1113fMK
XNGqZXLU75/8HrpepMhKSa5LuL6U0rj8mYXWXxh1erliQBvOk/IpF3wPlvtZv+il0cKYTMZdAr0u
6ldo3vzDNrEagprV41hNXpe4HCAHveXVFH7ZqZK2B//NODVTJPi6rZL+zC2H23+Os9EwLZKdoiGp
kzSoTqHpIr0T/bkouANka84kZPDWtMsp2xJTAp18v6cGJADkdc/xceOtFcT18vQAgfx8MVjYojgC
rjLLEQnsIr7pVYoz/LGJK8eG0pv4TVPf/Lsp9cq7uftJCT8hrwFo0ViQ1VD5xtAgZFfg19ujFKB0
drbxs1m57HnpWeodgCqbHQxbOXeQPA+Da+4Iv2IulxS3l70TPhBkoMf7/UXz2CeMXeSZY055FIqU
XOn6iz+wQEmgeYdSXWNpFhDaOX3unV8h+kzsTTsS9jvp5ZWvQXfmA02NG7wSi/hn96JqHMnQUlb5
W15Xj8oqyEnVa2c+/vpt/xltzKDSnpUVzUMA/U0fAsTpS2ZVPlS17DuLGfTvbIrdfDGr7ufoUzNX
AVeCnS/y+z3h2lXFgX4myGrkElBNAnoVD+aQtpr2bbJWLDlnqvb4ub0jVkUpImtuJ9RAZe89xnLl
dnV4/KDhYbPa+YGGsqCY9XtPFGR8LszxmL7pHd4yDFUG7jmOgzOh+61ZWR8JOLCeNa8tpS+EdOe8
u6PJGypF9rBPQyOUCshgnmPPFVl2VrPHvD2wgn61RiO7rLVXoZ8l976126tGs/CkSLzJBjBhRljb
lbZDhErCHCrWw07paoQuQo0zfv9ZSsIeSoE3FW0qOEJRWxa42ixGxP66ByVqsGpe0IWBjhQyig2N
MWnO96H6dKrBTwZmBIo7uQXYV3cX1Jzp9vmpEETuGzkUPJarCt47JYkUyc8d3O2Q1LhLBLFpWCm6
Pxw/bGE1xIJkt/2/VT5p8txUgblfsohdn7uhiojH5DbP/1VKvypMZD/s76s/9dH7Vy5Ly/45dxlH
+fa2MJwb3SZJRD4QvQbF/QfhRqervACqjUa1qQZjzHAkNY2llU3WEUG2NTmObfG//H8yFagBQjGk
GmG2shsMTwz7sD9qYeOL3QmlSHrXW3dKUrudaEWyLp4n37xfJuZqUaedd2TSh1GGQbnoshYbNSMf
7uN+ZrQmJnXLVJ6xxnLVHGL6bKvmzz9E7WezcEjy9kpEAJ7DMLz29bFbEmZJtCyCKd0g2Wxv09/6
0msSYKIgMC9OcI/sz4cybdfFz1q9ICLrRVtjT+IJT31GX2HUbzNuJDfUJjkkKzZ6C8qIU0PQOaeL
2roU4wtQ/Y+gbMU/X4rFjsKyMKzhg1TcVjlg2pLgOELDSIibBVjLKwNCq6BJr/VJ1PU1lUThhKJO
+3P865+j6lwsJMZjREUap4a2II+It5yWjalfoD/5ooZTUm5UiAmb6ukyjkfR+/wSZitURbjq30uQ
ZRWtx3l28QFa74cnDOjXwDHxOFd34i8zTEzFZdJobmckBxdsPCm3rVJov+vBGSyKElhpjFj1vy3y
vuhsAsD+JTihbZtmabdOBHVaG5iHiAHTxwPyG4oIscjWPRj8Y0F/+WB/SSVv9N/I/WZrMXUF9+so
xotnJNP0GvRWLclQh8Wm231QTb0mn5d6svcgvl9L70aaX4BnGrIgvbXKcE0NP4jGP1XjcYGw7vXX
xoO2GxaxcsLUkYyDKElw++Zn6h5bNjJwenW4rPu0/Gb833kSerO8oeCJNw10w3dbW0BYcV+9z5YA
VRXOC5mLVuzedP+BDAw5xThMw99R5OsKFIHsqIGV6/LWKCs8OTCGeXpXClKxqT3ktrIl0cQ6Mh/U
rxz8P4u5hCOlmPchYjVb/+nDCqCvoqdF0bxskqzo+dqc/osPnHyiBcKxbiLQS7cvjfZGF0w425BZ
Rvr/Wxnjr6n935DyKvjobBpyIFLSL58fkxu0W1YApOamFRSvqYA0wNhrRVUBZXrziaOo+WQLpGEu
+c3XOMPtGFNk24xgycHY06DPbgOXasB7jci1vFV273qU4IPBFv15rwG0K33exBmGAI5tKiJRY/qp
+2BDrnEouPFIVsJ9mtWtydy+0wxhGe9UhBIeWWbT0IkhAJB4xCFSqSBgEemUia0oL25b8/xvH+VI
EZj0LZC7AQQ3dWYw9mVVOiLqnY4X0vtHpi4fUlM2tICoMmJxG2ZJ1sHwG+BXdRuiBh9p/m5b7Us7
DaIPNHFhFw1sjKLcnB1ziTfJLWo5jLbN/PLnKcv/qpuPK7i2NvAXSu+i0mz+qb9xfKf9LYIyaepN
yyGieqrgwCmor7BOtHaFOqepC+XJD2qAkESRYOEahoKNSIv+fFh0zSv+p/dCc3ZYonzY3Z28HjTC
tbuZk5MtyxPT0tl+dMx0I6MhV5dY1jZevRncTseuEJno9yj57mlC1RFb0RFpgejKhLnFCTykYg9v
MVmIREUkA3jRud6RxFJFPVu6XXhRSl+NtC72pHoQjvUDGAV0e/P94FZG8Q0DOsB9sArHSb3ueBi5
GOlNOEu2ErTW1UFmU8BRwPgTniQDLihrBGFc317pGCQ8q+75erPJoOtUCqOgot8YPFc1pACagWZJ
QZF1TLz7x6wzB10vwyk9aXHCBAzPf+NuqCPMxM9KR+gLOIId39QBFNL+Uc1wyLnULcsqwaPpj365
Ue/Wa0T9l2/c+0xkJtzzi3nrhFbS/JauT9qrOgf+1MZeoqGuZvudSLQrMVHGWVuOrKKN6nbum2Vx
GMF4ccKOqSmtTxQ4pZ3Kr52Fz5tuZScae6wsFrjbkUcmQvj94aBeISCBU65RC8oos/7tGu4vgeU1
xqC0NIG1dP32K/DoZyxe1u1JIQxxsHfuSBCLeJIb10Of9sG1+bpfetOVpdRkb8ythFkSwABy/19m
h0F4D4iWhBTDQmoAxXs0JC3kYY2rEpuVqiHsLjGq2ke+kxDYsd3jGeykbPDlBIBfyiLu6VGh/RGx
uJu87SNOq5ANg6NPoWG2Ia0+9RAPcoqBk7aD0JXrc5ea/ZAj1Z0AL6LuwHZEfxffm4brdDlORKwf
+Mci6/nvsHK4D/1oJys3RI8vnCFKacV6umzgWcRfvuWOs0nLPhHqFGEHBO1LMQtNS0SzzOzZKX3F
LXhoEWD7twAJfts1cHuDCLISyYCbLP8C6W5euo20YZmI0SfGwuKt3GJTcU0npe6CZVhY3jMaTOU3
wour4/uTos5GfXYDev5huL9yW/Fn5VuNABdoGZDzaFTqLSg6tLW0gFGqux0GER1IdjBEIfZbWh1M
DOgz6IECsssYQxrfgngy1U/eNpMlkJ2b0IbNqFzSAXX54Ws8BDlZ5uzfMYMcMUl2AmMhPJ9y62kh
JKRchGQZllAKliPybNEsFvSYbeEF7lbB75ykkjwtqDtT9VK3qj1EZ3t+lckoG+/n2Qs4JA50aiVQ
Sa/QL0GwT0g85wRwxy/yTvQ4IKDlC8RBfKTL99zQt4lr61hdx93oDPvRV0KRe1/NBcm+YJDZ7BCF
NqFhHwX+25XVQ8ZM76rH0amVgdMnIgYGSztwWIZYICuynrkwseL2FiG5UZ07JTIsD1+0lq5BNT9e
kYV1hjbs60HXfnXbwRjtbD0RW4hScpSh8+hsXVmuHwRJW6qcEqNRlVg0v97kIfc0BBWCLIxTdgr9
/XqROEb6Q7gJZknnCLi7eCC2QFkMuvaaN48nrZfMYUKYZsKBYZp16y4UWTR5DW3UWt3SFiahwerO
NRgYU1k8hQjq/54IGDjZTh2Oj1PaJRtipK0rd28GXotdHyL3UgBxWH6kZESClJjqjFxB681VKctC
FMRyI5Hd7QzAKnt/CCpsIngxcI4G+OcgJvzmHYk39unzhTVzKn8QzthxlDV9XoUVSD54ezH4/M3V
3TcUPod62b1aAmrGo5laFoC3I0wom7f/yNMrmBz4yJmK+J7NZyJqC5Xs32EHw7XRtkjjcutI9/EV
k3ZsffyRS4A2UDQK0FAfDLKgnS2Xx88Pq+D/b8x0DVTpbDi1ApIIVcAyOarZs384+O11COuF1eTB
E9dc84qvKc0tS6tp/15zuH+W8nPpSPQzm+8qQN6tdzJiC4N7bBWK6ekHfOLTQ6ZU3xxt3fpZ5Tn9
6cn+ditlFDBLKpnUn9PW0B9ej3NHHKdQInzZjtTZJVYYR8ZzmlIofP6UWK4OM9gKZCsR0XPxCZQJ
j5aQybhF7U79XjOqTxiUviVkbrcxQSEESEr1yXERYcfD4DliYO6x6drrTgGuyTusRM1HdDHA/Np9
qs7yfzmBC7WiJlsJxMAdvorSNFgEV4rZO4lPEbEb3usFGCqQzGjA3+Djj5ajSl1LWm/0sJWE4ipr
9wIIzX996IpXFw7b2yhcWc5Mqd/jIPpcQ7lBGK8x569JNs+cEHQZfXXkDHgj8CX9m6U44yT2YG/x
zlR2rnKVNtErZr+dFbm0kqVcldHRqA5DpC6wXp2wzNBS3QAMRpEGO2lf6AjJAZiGRUC1ylRXF2u9
7KCSLK7tkqqLrLAsRpW1jtcEP0bSzUj4oBRO2+k9Nyx8PbR/FkEfEfZxl/YA/V/xjT8U8GfDWwwL
YuwTTCHBJH6Bn4otqCnPqVJ7lsH4KzC0Y2fRc8vng2Yj3x1afovmWAeCihfoXhSn3p/e0boErq4W
bmQ2H/0P5tA7bzgYFSrD6XuhX2QNJAS0xNgXa6LiE72OXlqWS8/qV+bd6wXln9aMfTO7gqhSxqzv
PmLFyXZS7Lo5nBcBfJgK6O5YqRf7GPk2+Mugv8eb4MI9lqQRoblNgtUp3beSwyFQ2319Y4zbBQse
QN4d0Vxu7l1mJa84zvjwef5Xo3t1tlquVecixKT50gCFJmra2Hf3LJM0jtNOnvQfPtCljBuW+9Rm
M1x6RW5xKgEc0NMpHcKMYoVog15yWTmQvuJM+ssrd3PpeV7v/UEhoITuBbZtrwb0IrJgkOYoD7k2
9cO5jJEytLMrscv5+13D1arqrnnCnH3yshPuJh79hzsuIZFAyO7JI6mkZaIHO+l2w5T+tbbZWMeT
lBwZNUODFQaA0hlLL/BRajNIFmeAFI+QL9IBAzGy3v3+Dcxy2TO0WtNHT2WHHewaLN2SZHdkUheP
88gMC8aRM1OpHmZEnHWg38ty2uaxUB8I4OsFKV+AJSbatQGYEpqtvcfG1gQqdx/FsJZEFSLtyiVg
hIL0Qb4X/oPVlhdk0hMP87DXNAXhJcYoUk6k72/5S3oJNrQyzCg4TaJGUSoR5g6KlKfZb3NjubMQ
APyPiAIJIZmeKravy2q7u9JYrQ9ODSFXnqYmhkS449G0HsBGyJHJQeN7jGNs5Fjh+/W3jHwt59fZ
pIISt27mw7CHde4zlwLqkZSquhNDGLNESX804LaPIGRAngjI5gNs19WBUc0TP0UlhtRm6cCkGqGx
Bck05E390Ypr1xjA2AgsgzBg6eiyHxOfHrdmp0SbVUh1LfzwQeyly4atPAv6/zzjQWnLiouSUwI4
Oz1jv6JGYWeW4azWIA1roquKL2qvsBKnskn2vPKcFhGMY6rYL+8RZJ3u0WCfnAHp4Ckg4na8pDM+
DzKpaV9anC+yqRkIzo+yVrVFOttXBAqaGHn3PhAt+k+b5xFj9lLkGlFulW7DpZpJNuLG19iY3ie2
hgvGWicVUtR9VZ4Tmod46CRzHZQjB/b5iU5jvryGp1qTYAUAJ4dUMoBBr9K8M1DkgUKZ+ki+MVBc
wPn1n13lieyGCDCQI1piOqYAM8nMGWx/YdxTXvGrecLSNd56LcAY8b99+/QxxVHrnrrJYIF/x6gI
/AUKN92qqX8AV27KobIMBcJKEgcrnRePp9R1U+xRViCaiqFDXr37NmCnuxF6P8U00rfoDOYFBZlC
VCYPW5Oe0eIUekKSLoRaEBkAwHJVYHXM4rwr0NvqvQmMawLJ1r4i9NV2vcGlxMLB/VGbq4nBguX1
twGp2VtFYQsfxJXpSdHkVBM/G4/unQ9+fyQTlDwv4JWE5ptCE1Fc633IigilmLfaSLaj/Dpp/HgI
YXHuqa/g1BmLjizUnovFmDFZ3QMipYdD4w2J15jJJcS9rmG4UXO6HM+Wxvt9lWtORAOZO0N7djBj
Vpq7R3NPEGsuMbYlBTUcF/mo/djIV0m/FtfEj6ibf9Q0RdPgGoN5YYbUPLSd/GIGF80ECVY4PSsX
gsQNNN7uKKnQ9XxWyJmupngqjL4vOxSYs0DCCv0lOD0M2y1WWlh5l0zP9hkBgGeslyqPLL7/53v4
akUHYEYtYmg29VOVr3S2dnP37M31sYHxRpcO3ND1nH516FAhcxzPfgACF2Q5etAe0iils0auoeWk
sAR1Q58ZOLwAXW05sZXAG9SgawzGRyezBNeuagsmWgVfYOrgs2i4Pk18fiml4IlaVx59YMFS3yMN
GN7+eHU73uRnG9OplkiIUMrVWmeg6iFDj5BzOAozatr6FZHjh1JQ7gQdrf6hRSajLqxzE22YJpTb
4wlbN8RRMo6uOMgdIN6kedGfafhWdklIeRtSIYJ2+oRQ9HXvs6/7Af3wXekGsPNApod5bpqLNt76
Q0S3wFfCcKbw4zlDtX2/dvapbD/WQPGt+8NkZbpi7doiM1IWlutmhTx8JJkrQ67W8wb0bPp1Cf4K
ZJLcg0Q2Rs6vWQqbQI9XqDqGB1wZ1ITUFK+2v+34RPf2iKCQ4LyepASjhnoTupqa+QFEsIVfVa1H
1thT7hUr7qtsOrwfAdpNJeyKmlUq9ecK9VmW68sEla4xvkC4dsgnpWB2xkEsDNLweHmwODekGL8Q
pjXdHLjP89PSSWF2l52QK/vpQTXD073aOr9UNX/LukWVX0tfg1G5DspxxCmqgqXQj2o1sxnChRpA
51CF65H1PqUSP83jTRmZ0dqiS5GFm9oV7AIfDULi5o52tygmuMf3CYnG0ZUtPEqiDxMdXfbcsnf3
zjcVs6dD205eHAjZ6Y+IlN83yUKAcj60o7njLNlkgeG3t0fBl+1CCZ/Pwc/pNjJVfL+k1e7ICgRS
G0Uhtl7hbyMOtQ0TmXW4kvbx4PHgZgZsKVBFcRRYvqfe/B/KxWSs+/zNavpT42hIOxwA4FfRWPsu
odQ8OFMDPWB5JsE0v9B0BkK3FQvBFfGpUVN+RAx70RGcmVyGcE3ZBP0pBM3aLTHdl0ta+eJfPgOB
bvOgibkieF/dKJRPvVabS2x6zY/yPdSKbOs0Sk9NtzYapnp9cdfwIUpzou8aMeiUPavkbVW5Wd2A
222SgAJeAwek4gCGKXEhqHFeKdyYlX7or23tweaFQc17rhhKn2tlk2vUrGUyObG3oCPv2WEoN4dr
inlvuzAq5iclLMplrbirW4x1ctkXqzBWYw90Y7XOmLR68dHiUReU0hk19vRqG0VTicBSKqoDHFnp
EwsTl3ezPB7pFz1iJ4NuSDPPd7jOvwX54zixDAY5I8q7pkO2z9hRzqE0zvIkUkSpLQALKQDfaOFK
SW9EiX2Y/cxjHsrn0vctsoNVo0CwAcG24jD3puRRHNq1rRiJsFyl79ijmfwU4xi0TGeCyrDRV2Oc
83pLCUhUxvWu193E6vbfcYTugVidgbPiQNwqXQRuFadox0veZVTK0ZW7nsDnfbipsVvC4EUGCvxi
/sjVAM/YUGcATz8/AqSuPlnkHoPIjsu5Ug/U3XxQpGIqZo1nq8s3+vvaOSRuU5mRIuo8BQJCY0CB
/dSBl3abcRQmbvYrmpewrFGDvRFherE+AMLEmcIveUjLCJmOk/LebFSOEZtIlneL1BylpJ4IqGNG
Wh+cv9eoKWJxs9axGYSMZGDf5H6JQdUgGgI+6+kcHQ8iIErWjB2+BoUmKHQIyl8rGp2CXa8c/CQv
lWTeQjfGvEi9kPmtcCHRDXXQvd130jdNgAIjx6dyndAtwxpTiwrgktq8JF/gVD/SM6TW7/mMQvUF
em1xLlM+K90ZvNea1DhRmeikiNUA0CbU++Bbnpj+V8TnSqtsUsxPH2jp+ZKm7wo7c5JSHAGpcPsQ
cKb6vOZZ1bIVm/v5hDpZ37AJAnxvQDHmEuwSG1ix9EyYNZT1HjrDOTLgqAgeGzGz9MQ5h/0kcPjn
2uHu4gjwsLLSODlMPb0ia+6SjRIct8LSkM+dHKLOgNaJyEbajFYgHbhqu9Ug60ZV3ffgkDKzKZAo
vl4OokyU5rPPP4sbjAiIDdjqWjPeMNZ9ThS3QYiYFBPZtsF/+aSpknlvAMBUNEk/GDqpxvDO1mn2
Hy5KVZPQC16PKKyJYFPZlRaAppDr3wSSwon3KiQQKpCXeH58eQvmknI+DDKhYpXoEpt6KQeOfJwT
Az00kpBewrMrcPcO7OTuglr7KWK9oKJ/yOXyIngonS6BbFn5D0/xwhA7ZHVkF7Ar+a54NztbAzKd
cjXcK+aaZBOPa6DwSY8TTY3GeMxwO94UWmhe0hh/WxhAzdskcqFI0JuMTeK83KDOepN0co9PwAKy
99WW/mcbkb1W6srHEGbJ0SQ0eHQh8bCmbzYh5vhwkIZTDN7/S9FxXxUyQJY/slj+bEiZT3Jz4pmL
s8cszuIL34dcUogMlAMLGEHBkodPDVLVk+rxlmosrJIIR6lY2Sd0fAd/KfAVbz90yxs7NXWvXXRn
vmYtV0JNp9YKqueOGRy84MPcbVYUz+Kiiu7qVWfBQZRFElVW+Gq2kxRguZyUgEnlaoQDwtZi/6cE
j8Qg9c2Z05DILWz8wSIC92Xyn6SnlpdjpvvxahJQtbnfsWdMv/3bHN7jfZ6fGUePYYu8iiofjKHG
GqI/VYv29ldkQKi3ooWc0SYH4GpAQbOjvGx+SVh6thuRt1Ko2RRFhApfbIjW7h+masBda/1upeRx
JX20HYW8qeWRq4g7GW9cQoCHfO0Qv84DpVVFxQhVG5WVPIGGSC9nE5eQQXmZZn2oV8ztU15yLYVp
PpiGPBs6qF63qa3g4BmDB/cF/HGrOHH7635Dfb6nhHogcMIrheHz1vYODrs4xjH0QTtyQjLotCdW
y3vFPmzqD2EW9xu3RcQM/j09IhV3MgVl8pqcWwSEzsW0uAk45txq/O3QOTarHw7vqk23/2J4015l
aS0s1ArZCt+fen75KIiDKn9rbExGHFLjfPotlyK0cOaBy3Ls0GcUhHMfdxsLq94XwrtZ8MFq70n4
Zp3NMC6urvz3DBbm8f+Pe/IHeTUfl8if4t53uzQBLCw8He3ii72puVKeZZ8TgorLx7++nYeyow0I
eZGRB5M+YKlfsh7QtQzlfBlkxuDOGzo0qqUuE8OkIpkx0CWx9lnAZAKZFwr7hvT3zFCvmhJGy9hh
NesahR81QX5EAtbxOLK9V1ETaVnAKp0lO4AU8iOQOw/mJs46e92dWP5w/CaQGiuVJcxOYeA1Ze+O
XJMJGCjPU/P6DRNoZwlKPXxLV5DVY+dhExNahUxu2w3pwYFOpd+fo7c2h037qcfFyGIrqC4tQiQ4
ahRvO1iL7hcgHDaZ/a4LaFM+2XL88QenCvuVXYq/BWmbyDrU+CQ5lCzwfzwxc3YuGwHqsSN29zVQ
TMNKUqz5uALzXDfmb4ZH+hbYB3U01yOlqJL8Tybekn4BmCEPki2iMr8qYA8Hs0aU4f3YMGQNRKve
Ji0GSMzm0GrHJumUKu9EsnZGnyiBnUwy90ildbGJZU4TEAGy/SHLbg09l3qjvbxEWl/kMQKq5gxT
9UKvEo8YWoQLaq/XQ8DyudtCum9KE2AWlUJNKODzmrXMLqAmW9P9tqmyqEvLFQ2fTHOF+9itZWE8
+sGzlZ+2nzyBhi947hhSVkZfhOSBHmx771sPxhp2ZonhG8PSgL2CRpyOZzNMvscdDEm0Olj2Js1v
rURMZMSSMLp8FsukWu3y5T3NlQzWNV/GWiErUxqChnuzVBsn7m49HxPp68OusFG4k8GJqq/qPcaj
fV53CROeODUYMAI9kIw1nezsLkeIlIXOUUZAR2rUGYyD1X6b4b5XQZyB8iqwFzlClOzJIgObST0g
TU680iiWm8xa0RNvp2JRe7RdiPvVVwuJvgB5UFQPY4P+WnPUl/apyTpEwTf7L9293A6S/dievdjy
67NMgIvC4b/Fcnj5EYvhJipiwSPkB9iuElVaC0Xen3P4KHa3RqoEu1F74nMy3lQAvCLckIlXrkTu
R6u0fqaHOzPqBEY0m3wi/JumbpVL22jDI+nbSCwy5FPSLlIZoDBuJ6fD3lO7KTwoqjSMEzztD+wu
6+ed7duqXhL7WObtx1E5/l5byNcYueI/PX+3ZV+Ys8DsgMjGzKgtBDoQNW4b1ebHwgrJgNyBRy2S
Brscin+mI7aOD1OflE8wr7vF2YisCoF/CRTBTAQbjL71/9iSd/ly0qfOOH1e6tkSQ99ykvKWV6JG
6xqlVMZT7i7HAiM7rhYf8eKMaC9usVqZl9hZFDgiKHQwLq0hGJ9T+sLJuwwnNao0xltGsfUcbVso
02YcOpbRhYQUZL50uedImmVYa78nQ3LVcq6BKapK/w3OcT5l+a32PDfahLCP1WSL4ir+2B8Na+va
H1pLi/8ILpNXHOgnLrLj1uYowRMWxkl9PY1PJPQ/o1gf2civxFh31r0/6nqQwpm/Wu9FF80TUqQQ
mEwPZ0dZVqk9hykYvXxp3fJ7lZDLJFzfTiZBbYlF/Km2fCDdFI0/ddPRixc6SVyNJnDmg9AXtCF7
iCy61o+WAyhrek/qMyA31L5h1Vmd8IG7r7UlAh+CiFN+JYU7HCRq8vN8nouccymKSoWljT7OPK8v
wcGJXyKhWi5Sca//v4XS97uPgPqxKBVeBkfXvnc/sCIFAhvh3aR/4qqgG1cuLJXhw1It3cNbUuJC
1crRgmVhO+C/WyNq/I1QY7sIMS56FAhHRMRSHG9HRIOkeEchayC07VSCdzxfqfhrK+jrNnDmS/P9
+ig//yyBYuPDG9CEimepxgv0TfK1FDQWlx/od/SCoRvu+g8Jkm4etRiy4BNp03vNQJkDL1bV8WlL
fuOVWsirGREzy+TLeMvG+e6cMFK7KS16PGSB4q3kq4nSniw/P8vJF8f1DdyRwYI/7jxsHI6gEDdr
zEKqM58R57ibZzHRury4P6NNIQAnamagExFj8dac684abwqDemedKPdT+96B1g3TckIBMSwSpEcY
v6Sd06wJYDzBByVKax/tLYluGRHrj91q3Yk7n0EoN9J/iBW/xVNosq4Wp8AxskJ+XyWp9GTXZLDD
cQuy1mR3rLmIns15CxRlKxRnzU6H5tiw8irqQc1IhU4BgMV6rD9HRsqPwk+6zQLDxICSswIdnRUt
lKBoOos4qSasf20gCmc7E2CCFPb9SsoYBSHq5lPOd6plOonU5GTCLdvdpGWMlX5crmaBIJYrLnA/
dDBpM/WGDxN0MZSCksbjsidxnDwBY34G9xWGj1MqIRrdB9ZlYiCEjTNnR10l9n+DUzAItSFOGo5T
jnoN41XKPK5SouK28JchSseAY346wDPPRm9wKEqS6MJkE6hbaCCgiuHIUGcPvOmeIyepySRlurY2
0vO4269eZ95dvYe4ODesfY+7pStYuLSeYMheA48v3Iy6/MQsVx7HTTolp8Fk0WaZdnL1B8OGq6DI
AvpZW46WAryoSXEx3W75EcayfT4229b9yrIWe/22vjdAdcZCOD33EHN2UziDDdbnIZ+ql4xxU6vZ
R4Q8Xi5swhOCoFIdP1FfIhw56V22k3luDXFSF1rPbiMnjDr6I7S4wQ6H4mVLESNkFwtapeoAtqzq
WVtS7afnMB0u/pXPUbUbts5PILJyQKVHlkB4UKSz770PPJrnahKHEewGk7Z4N58YqHGsic28o/5J
ZiPc6ZepTrtdK2uqhE/5HGC+xLsBDpnculiyYgBKwT23Dd2bu2UmFnNPsQsGIdo/IiaiXW9oMw8H
BSs2nyYii+QZdUJSCgk4qw16qNsYya7nMpJ74yIFjYfaUY+XyHBxJxmrttw1UmHzoL+o5HIUNik4
SGZHTracv9ucQQn8T8pIyqr8T/Jrid540W0Ryi1kr7iZNxrVC2GqIg1jQCcMjfhV+L99dil5/Q6S
CALDvZBcUEuQGBXJHJMfBgSrUAadVb9y3f0t3dHBYuDezr6l/cjA4cHRDYOBDLoxY4+8+1THaqjH
WgzOkOF+DO1YS9svS0L34FxGpJSllf9RvCKY2sBtRruOYzpB4ot2oKTVpp0fRDilvDeAm17ou9bc
pg1ysAhQSyEUhqDAat5OoxkZQtC5MFsvkTUnrqor9eNNrerfso99AzeHqf3vGbR3KeymT8RLAOW7
ktt18jXVmcwK75dOxhg/sTJokNayoO/7lp1gl9Yvf9meUB1MhqwQxWqvI3iU61YYiN2BlEEO+G2E
i6riGSH8K42kay2+Oca3cqSImtn0ijngSj2koCKjVOCXyWYGDZw7jOmYwLxZDjtnrfknXDLRh2Qa
1k3Af85qiC/p7RSvGNxigFssPAmkqV6H2SXYTxJDnOLNpMWqTKTyRdHbcswwWMf1p/0uxprFCUr4
qDFPCZrSgZbS8oJ2a/rFOPfKEbk7ssL8Wt3+pvouIjM+x+mxbuAczCu1p5BaNiqWTwa1jLFHfElA
9zbhBSx1tW7zjEI5qE7riGMQEEdaLF1pjOetavpV/nMNDmBv4pLJ6lTaXLxU4O4MVOOpFxDvEhdO
UvFKmoznffmXrW+XuJKT7Kthjl26dHfFaiUiMloNA2OJlzD2uxHqLsIRuXj+oEms2wQUFmdcreZm
EJAGx6KcMJX+/cHW+A2c9bH304zR6YNO1x6A3VcI0MQheLz/km7SG++ImXkbR3Z55euaC8XMRQ0i
OD1/vzEkXgHGC1HGOGP0gPzSJX4Rz5SSc8IW1ZVuDAL60aKA6EYQIQlei6ZyseW5GUzgzKYK3RDw
9EkJ+MaWL7TlopgEz3KZPGLpcFhVUmv6skUFNI2YpeOvjYKHA5ARu9jsN1Gy3mQBpW7DeatpfKmO
Xw9q5WP5wPcvaL1fo8GdfjdbCVXi5qCfEH/W1JWw3s6gVsA3pGxFFF8JCbwBIeFZbuoJdIM+92jR
PqQgfBmiqivX6eotxR4ZUN9XLGArUT1p/tm99dNnAXVl/jOV3ps74CgBR3kDHrErdEotDYxl/Tcv
6Iih+mZtAx0zlKX9/MX9u28R3nQEuM/3bId3qMS5/qkAZVu+2MGXUHDwNjPfar773LmUkb7oVMAN
newHDnbOurY4k+9VOCMYcDZCCwAoH8t3xP4CyIID6KvdjVzaM03fJaVeWfKUZiwlAGd2bwT/Vgw0
2gjhM+MtO1qFYsi9GaZAj9CzQp6yfH9QfGYxxYeAdb3esGsvSEsKFdJDrB5P7O49OJJXKKaA2z3L
nnHmin/waNRGwm2qLJCar1tHxG7UmmrdfMQgKBrK5WG+JBEdqqi+CaGa4WQatEN/xX4Wl7NKsgHq
8Nlw6tgpw9nECBXovg8/GkCzFTSuFtlWC7Wm1gNwTGe7m1ZS6J7PZKBhU75HYWTZFjpkqBu/2Jop
cjX8Soe2872B41xu+UQ6jjc3BsppE2ZFF+zxE2WJRE/s4Ah6ubV2E+Z6QfalPGBhQF5LZJq75Ufr
TxVMiXnoTgKmvz/fXplutHjyhD6gYrVBgB/ZO4X/gh1pgUJNu8CNSdB0TXDPH1lZf8aAit618XWH
/rith5XEuOgdw84Ga4GQW4/Yy+HnQgTXIhA2KlcIjy/c3cSTMg9F/r0w+4TfD02GNr23n/OD147m
egasoH/Fsemvekooss0jF9dJOmTwuJbnGcv7vy7Hxm/RWbR67lx8Uw3FULTk6phYv4ADqZF7/z2F
+Z+x2s9xcs1ofmjkdRFZaaCLHrXsXPI0fo5jGESGqmsuza14KdG/v2IKUGjblh78SdYC08v0IQSL
HHOgZ6tzgBIGUFKvAtsKmgKL30ZE8RFX561kl/0o3pojyAYzd4Ca+JmLiByk/f3oCRxMejCQSmj/
7BtHLxMX4sJLB5jqWKJ1q/ZNA1RsxuR0q+YI3vlHjuJyvm9g4x6S90L7UQRbySyuerpEuPWE0RL1
t+Hrqwl3tT1gVUR/N7FcwU6yAbz43WSSJum6D4sPuggpDzEjgg2xvRbmJSz0ldn0q3lwa+HdZjCr
f1h2g0WSVbadilCHIWtfJZ5UaDB1IrK/3L56n2ihY4qZYv6iLdV0IKdlb50rJfEe2daw0NiK//kg
rutZZB48dW2goffz+wMr/Gqr/oLdISvPt/o1Bslb8BPORyMi6fAGbM7S4c7n3ShpsimUIqaInjbA
UH5aZO6AIkjEBvrpag1MXEevDJ8twWfL1AP27MjntcNu/kaxOjzP0pLL2tb2nuU0DIehkd1cmypj
bh5fgBnjHJzwWcYBjXfXKQLoxBYoiN8sf8Ss8sUZsdbA9oZqF9DCTRKbdrfzwTTDy4gdxJbauatK
+eSr7WbLdGFKgxy9x1uLaMhJGZ6WsZjTZCHn88zRXUO6nQQSYs8M3/MQCyA28wCpp1T8gMZRJMl9
KxCU5o2NxRCRyVKZCidV5MMuuuU2xbJPWpJXJjFMfS/+XH2D1HAFj0zc5TIPs2HAnU1pwjOM9khK
IUms5sR8bVO2/kUgRpZnysq47J5do/VNj01BxnD9MQpFzY3RvCPU2EziVK/3n9tFjg0R6BiNfmN0
d59G9DXWYPEAopo/DkfWgf5gjEP3/panG/TmbYrNYeZTmhb0AkkQpWYktz7vRigt+fqtJdKRBJyZ
KqpeLxA4LnKZZFaM7BVEF4o/GTeUty78CmdO9T8UsEh28ijNHRoBtKSHgtJVZY0UCi1JF00UNS7P
69TvJ69Q2CCTMcbo7sI5v6XBQuCuGx7YjGnOwKonRzZlQ38niGsLr+EMzddoo7whoOoBNsb3KUHC
b9W3u7ShFk14U1+Ser+OfuXfpxR2Y9FtP1isJkIBQNDFjFnN637zTLbez8cAkgbiWNZZH76jxvmt
jLYQR5PHeunPbXq494Yo3eyIca/BRbMAL40+JrpuQwE9Y0hVCuqbXhdyPETgjGE+SA/FAlRVDcEI
6BLUJtvmXG4fhhEme+REUkIoJjV6K60Nz9PIqkZxD9vSixnBlIpaQixHUpRhiFrTpALiLRjIqy+H
jEMDmfLCc7Ep0dkSVMxKySey6Y8HygF4gIcThbBv6c15WiwkMM+CNx7UHLJ6gsDDnOpQUJ1r0RCr
ntbf1Gts6Wqt9axRyuYBIPx2SgiK73aIeM7Ww0Li+mlELK5nUnohydoLVPR8yx+p2FotjplKwD+e
GfKAID/itc8SXh2jGrpYWYcWAgQplXdBY/gEtS+0X8DBFssK3m7cc3CLljEmI1tzNXMQAdsw2w0K
PRlH0kz4o9lJHCZ02tB6LzP/wOXlv1/L/LNrAhUqpGn2eQlT1FV1VNx/EXMNbpDFX+m7jh1aFR6H
aGdV3qSKVtfWm/CBHW4iFwNZbLicu/Qgr/lvXRNC70r2lCRqNgvrXHHtuyfCpt0bKX6KbmvOhQtW
9CIENuG9qJXzjdGyOu4LLYjY/rZhR9hwICBPmsVMBQq/2To2stLEBi7eO+oYBvMoTtspfNuSRwAd
f2UnDe8GC3C2Ae8dgLtP5EHdKF128UPVvEX/qqYrGOp1jDwAECbRzqiUh3OBR9v7vhI5A+jFqfM5
r0gNrRCPQnQNmBVdcDffjkhExrWDmBXjm4Efh58ofS0CxA2Fzc8Ngw79uuoftCNNic7ts0mRx1M0
CBvJ+mQsQyJVHp3opCqfSbL+oZq7r7Ft3ibcCFQ+k72EVSuaQj+cZETHj5uNTFGq9/R5R2yr+t4g
OLKCdF14p7ZgfLW6zJy5TQ9FN88Q0LLR8isWeXz9PeMIHl0RmN+f2ffIATEMybSnlLc8te+NxHVr
6bIRrNw7qEfKnSFmc4+1dXnqxMUdEmfHo/4IbW1x5rUs1A8/Smn27peNMjfqtbxHfJSJaQu8cpn+
OuSuqNZk7eJarHDLEWQO26B5Q+4OhnjvuQwWIuUge9FcvHvMrvhFCZRN+ck4wi9eJyy7iwB1V0Hu
lw2rNW+TI42nM61xrxaGsrxYcRys+SF6n2Xg+EIinIX29JVyDYAGEfPtbbmKYA9PmUBt/rGli3nd
3v+JECYbbklJ0po5f8qvoTJE6USxczuBCNeWIjpYiJCRkx0gz1Ink0xQa1xPvDmadACFyp4wCH24
ufYvFHI3BfSgjxqGPOto5hLLZVlszZmbeUFsnGoKcqmje5Qq6y7ROKxHiXDCVo+bw5STJKT3sr/8
vSbGBivXSyX5kYUVUe57kCDc7LMFeV/NNxlZFT+e+Vr8yY+KnTgnE3Y7yguguaiW2Z3g1IcJM7mI
VlXsuysGv4i4FyrwLAgQsal4fnlbwbY8QuoI9n6lT5DZEhiwcmSUTeY+IldqTcIMe7+yzNosFjLa
+kgYQfhG98dvKIG9B8L3O15k+dMD35hnoQU8ydtUYLIjJrdyGRIQOsH3Vfwwo6RTKqgx0xDBIvnv
j9gxO3JrPTj86UwT0TfCG5rJ5u6YQOo44s9eo6iqJpotRmuck2xUxlQ9+cWuTYKSLET2C8WVTxtX
ekhzjndGQfVN7E4Jy8LKwqUycja7OtqEMeZkYoGXcaB/MioWvI8SyZ6jwJaRAirdmEj/J3SnW3N5
X/AGtd3O55jBtoF27dwzHbD/LQbqrNr72RXroeNZa3OSaLVmD+cvSp7BVUxy6Z4GUA2xHAUOPKcy
XDKnkQRqakeyrXlk6HYnqUswNfCN/yKPw1zP1vxB3LqZ132aB3Spw/J+wkpDGrbGLlWqTclBK4JB
WPXC/zR1G0ywlmnr/cptT9wvYKEiDEiLqIgAs7LPeTYHzCaxt/AA0ilZZju0ZJpixOTVtKhDkBj8
mrrD5L466C8Y1PiJ9PxsohkhLylwwxnQsMIWyYRI5GaIPPpDc142/4v8c1ZzJ+YYcWa91UCJGyB7
S9WDh3/wYgD1sXBK+3Ih6yB1BMxM+EobeW16H07Fb1Is9hkzVo5cauS25tq2V0uhcCNS0h2Jr72+
ktXz5WjdH9yMhXVGuELI7ItAwo9NhywPF1Wv3qi8zrF5Ht2JjRBF1bea6pTe5Tb9aLC3MbBgJB9R
FPfyC7Zw5+KnB/CWQ7HIsqihUdEHU8oobwmM1dDT8ufkEQlveSoQ+kPeEgPZmlr7tqCQrMzE8ep3
EvK5eML8ijNUgkNHRsMk2b5TJVzQY4yNSQ/P5ORQbfRiNcrEv2YTvUJ705XpdEqCz/RStiRHPhw6
edH+I24eoqcTmGOoGaRQ6msbhDQbOqBsdreWbQnTprNBWk+oJnwqgu6P08gL7rbNpGtDeG6aSLwR
q93HHHg2IGA+ktNW1CF5a44UMC96LWGKehKUAsTxw2HKs8qU283YodO7lUBanvGKYrf17x+FMdkh
VnFcdDoX+YFNIIdvh5IkjGUerd4xhOEziSPhOk13MjYJESmsF6Dg5Exo7CwNxpi2auFqed9EsWma
O4bxxNIvuxo2D6mDwRp8sBOpbewZbfxr7tHE9jb1ZbBdoD4KfXJB6TPADINiBxdhJgP1tDG9xbpF
iqlRndcQBCB/kRWPv2pgM6M1Etzq8xQ2EaP+Ag5kVjMn4+L/Q1OLkxH03t5PYefIdS8gQLXgE0v9
eiyAFaMfxWG0mpAGQrquqcOvpnXFUqTfeB4veRaJ9ZZ226a+jL0nJuYetyrk0TY5RJH5i1vbd2TB
XLKA5eRXWfMFVe+uwN74tnoqMVWQgce57/fBNFYY1yV5sV8ciJwAUpEi1AIVvVtK3T7HwfYNjSeE
zNd3x8Bt6L0EiVqY2627NaSKMOVqzLFvFDD1Fh1hzbeKNF+WLS+bAmQievDqjrOHl3aUXgZrEMnP
b9Si5wtGiL5VJd1B3y1QpY/rEejW6wJKZr8KX4di1GcEV+ULWNK3+SH3cnR5fbhVW51lODchZnGQ
iUAj+6sjxSCIkrnLx/5Zc/qfwVZJjCme25arZjGrXwvrxS8ffRiqb0NaYK7F+jS+6P7nKMu0Vccb
o5zc257YxHoE+/G9j7njBDZXSk/0e1jurXG+YrGj1uGHDVy1jRP1cvR0i6KB5QniWqd1Q85xJ0d9
/H8aKRfVCjQJOgWozpcsXIXozs9hfdZ3y/BTyAheT0dd7aqeGAhM3NBrDIzory4YoPux+uGQQL8s
oD/lQa9nLABV8NOKDFFRewLaIw0nsqmcRrfNWq13gAQs7ngOhpD0/+/s4u4tqm0EDMtzBA8fMhDj
I190H8fwWUy7Epq0J4+86lyAQw/Aij+cwY56/CW6T/AXLl0+M8nYfuUDrW9GQLOK9Q47uTltimcv
1g4R5pGKAmQzzP0oroSuE7V1EXuETp4K8VPLOeJOY2wIwemhnAILST2xL9MLF6WgKiWZS2y2o0Ab
uVrIuRSBttNbVSiiWIUObepqNlnRuXC07gqZOoz1ciQTnz/dOml/LanAmXKs/dhrkFVU0B39/xUb
0xYIZRYCMzPYg5sfBQllEkD5ltEOS/O0cb1ITxr7je68SWImmyDXrXvu8h4ECBmWyxx5hcsh5poo
O4FoaNzxgiSNJPwHtjNRFtzwYdiXSe1Lr5xdHYWsezujnAqiNDi4Fs1/wDsSrUlvZVcnTkQIAJWK
V51LKFgRqoDB1Xwcp4mjxTL+rnhedi4hbLamFj6P2qWPVK6qUCYLYXGExeIZQYVwP59cYvH4j9oP
POhPMp+fyi66Gdr5B+hzHAZ5tTWz8j8ZsGwtwUUPZAGE3ybJveq5ZwCyZOCxU5bIPxlLvfMBDqNH
SRkYorNHNaoIbOqMS9NmOES+v2KdnIAmtHZr6pxJp2YupgmRUA13eW761+ZjsUCrwT8y54YghegE
mx7UtqhOXHBWbESQwYJdgr1Hbv+wXKgnPGxQH/hPrbqXg6hsMjfbzctSOVyrDt+KcEw9now0JWYv
WBWzgHgiI4g7SeEpOeZ40cySeAWz9twA9FBDaCKXK584I09sEjrXWSOoTzBFsdztkHqM6QdWdHOr
9KfHlhoSx9VJ5Ie0gZAvKLCxxV4WKToFiLjXdK02R2du6kXM0SQFFynv20fPNSVvJ7P7+KCS6hpo
PbPYyrwKvavXSQ89UeRIpwmcJxkEjp8QcGuy+TudvzrXqf6ybtO2ZIYzNDvywEtNgA7KsmXBhE/M
f10gJ9Aa7KpRj48zGQN/0fe8Q8EgZx/HlCxBDksnebIFppMkoxxlmeaQabHAwtQrD9PEDOkZTpaH
rR0vhTlsPK4U02/JjbcWzyXeGwPaPgUFdE8Ouevx8UT3BIE0pkxSEv88WumXlTmXGlegVXzkX5dA
zsBTfznDsNfrmw5JPOwxpL1d7TY1+ngTEBV68JE+hON0rt/964OIGJzYpEEHmTGFCU5IXsyZgawp
+ALGNQaDp3swQacq+IH1+vOdiqMXHDD5vr7TvSZeUObYaN3PePZ9jORTFHr2wEgC3mVaVZBGMESb
yKWtGH/XjUELglJpd+TR4K31jJ9rDYpAmko64/QOT5mSvHf2dErVNZk0bNbC1iSskRVV7aMmfBL4
NjSrG5xm152u4JVG8szc+FocuToWYbhoivadVIUqG+uW0MxSXFSFhgEzSrrZCpXOcxZFEDm1Mlvq
CyFyilYGTi1akAfcybqcD1RZ2QaHbfYlti/kqZYBIp7UgD/8FZ2scbkhFEgGT7BxI5dV0T8qQdEi
+2JnDCPnBN2olUVIs1skaxq/bNXCDkoOx1DfTTV63kUPRwMORJPb08Onz5og6kqgFM7zKcxazLY5
ZjjnCyvXv85jvG0i3t6bfWE0WVPUNNidH6JNRl8vCJDysTPKVmc226kmHtKogq58ULw6f+wPlkFf
BCNwG/3BbvviFhve8Uxx0AQW9TXUbP1v0NVcU76CNAYKGuOEnbBV1rAB79zubuYIZmZRU+WM2d6/
D/FOLgIEEITVnl7G2LmNhYNpH5YPDMBzLc+KaZ3Vwwg2tYEKrpxH2HS3pIomOgwGdrYJuGVtiT/H
7BpJJXVAEPmyteHG/tLfK4171OG3Dx1obLKqaJSZQJkfv2fRJwAZwKXVU/gQKaQkY5EejkkM1see
oxRKs8vYZfRSqCNvgHeeYGcAd8xsxARHD0zhwMfqxAiEgP7+1uApOpquh/5zaKmRhV51qJHNWN8B
gjVRRnwHT+NnpyhpijTBPhcdg0HhHMSvbJGSYyb//NGVe59a0/Ufm1pzHTxE570YewmKtmA6uX/k
LNYRt6rlIxxGnrhQYNCE51f9k3yW+4nzVpxPy1bN+BVnRVHD2XA3bCormRc5yHyFsBz1D+G+RQtH
lGoVopZj1AgqHmOpElNSOqS/2Pv4hYy96Tihy1p626ZJDi0GNxfZVrlWQ4X/poyyLEFt3x0aYBj8
p06M0qPL6lQwfN5DBhNQ5dcMq3hskcyMs6sv8ThiDIUCgqwuBGRaI+a+VRaU85NCT049fxdsndol
uOtR619KrN8U7anzCs4uG4yikMWNVSX6nSNytACDPKZZFF8GdAC1MNaINhmNiMCAqzqhdAby82qy
7F4/ckUUn1+0l3Q4fn20TnM3NfpO2OQgHAW6REd8ZXWOfABxGtFP9ib37q5oaX7X6l+dZOJP26tt
/SjObjBnKo7otL/CTJuyR1uZiu/nqGOTAKXETB1uPOGDJjdWciddPzSoHkdac+JvXnybO5gl1/8h
zBQcDQhwUaDiQ/351vJYaeeaYzvJM6I+Z1dmtmoirDWVkh5AxmXbOKPMqZz/hrjU2y7vSHSNfpR1
24GeaMBazyalB8vdJAsk5/M0P9/oSiCbdxgafngtQBrDrKdY9VMfcazgC36sIXH9WxAn10NJ+3oO
q1FxfDUgCrpjJg7MQkNO4lwVytdeIVsz++fId+Y7YHU683zjmeqzDVwOeantvIdJ69+AABRHS18T
S+KeKQwotN+VyX9b0RExrmKtU+N3NOGhoSLPXDZjT1AM7l51xfsU/Q44few7LhVZWgLJkGG3GJF8
qBKXf/vs5nCv0YVfb9I3tbeGNkKNs8ORjiUV1v02ILwO/z6JDbCulc9gJCEF27Xuz1DX1ctMd2S1
SI5EG97mj4Za4loJGL1gyFKu4s54+Bs9+rHmFBaMY6dwY0/dc4r2bCVzD/+i1Q50fFskZjJt0YJk
viEz4lqs5Uaftsf60cyC2q1Hvr/Q9Pdpa1zQ3SL//wfXpNGZ3fF4iaSYlsTCHCnJ11UoFjHbFcxe
2HiS1eytSN7DF4ijmvbdd9brvUbKOcZB6PjRYu/W94wXVocHKYN8/WhRUHJzOAY4pclLiX2ocve7
zNwL15xU7vH9LoT9L/tJABUcxJQERFusCa90l+rS3CfsQ4km36yhElnpsJpc/RADRZoQ0LruDLgn
6m1wt7IQsMEJsSYSxusz6bMIQPksq7jG4YIFPdu8l/9V9XestmxzvLChver0CWkmCNmVmG65dVgB
RlT4h9Vh+KCrkTcstxO4b7aJ+OULxE6K9eOWKd/HtCaPv7vA+8cNVrCT86ZKJhgo+39FTu1F1mEu
51xxvHMgirp8AydTu66y52NFlbWPQXDtS4Xect++ui/UeTZuWgrZVAnuAe4iZV+GypsDZLO0ooHQ
Jr+VoWcnSUrHQYWkP6ZMzyRHWxrzYyRnZiW4XNzro4mkXNAB2TAJmD0SLe5TtL9ZB8vsPwbWQgN+
n/d4XxEV0aWZWdXSXLjR9tdHfSP3lCxSISJUCk7GKc399wJVRDqfTxcu/Te6UfquAlAVYOzekmMe
mzhYYG5yl6O9NBO95peaO40RU0Xu/ks8hEPUuAzXYaaidX6D/xfdgT+555NBFIALEtNM+iYIG2Xw
1NRy7rvpgZQZBxcZGYCHheu09OXtwu1zMzVg1iuzUShPz23jkhPzm+aido0fNfQkBt1B/dvDYC/q
FT/Gzyj9SDxczFnuxjyPZJuSd9KuR9dG0f3Z8gd8yQydVEnnNZnCXJmEmNS9quRqyOtLRPhouzYM
WBmMivbtms3qEWepska3mDKFuAoBXLp9OJJrnLwUefD6yQp6CFMRuvxKTicpjmgXo5AMgEkKENok
gR15Fr+V05L4WqJ4XIEZ8FveQRyEYfYY2eX81ygpGhHupJpd4olUghkjd5u6JzjjmXRlrLblRv/e
epIuqzrY71W7VseCa46vQo6t4nNSjKYnJRS2yCfZTJqh6OZM9ZuJ2H8+lG0mr5EONuntLxqIpmys
KQVKqo05LiqCIo90MPV0Jp85yYAZ1jcWXLVN5REZVQ3TK7Tb8DcSuHJhGr1xE3bQZrK4/weoedCe
U3j0ptH3MDtLIWLd0ccNjjq9E1skYfgaBVhPTxCRz8PuNH89rqTQDbmQxLEQN072vKg2ykv7Spwq
DIAaMApRcSZpk5jKR/kWqiNMI5E1K0gkwT7uAIuZFkMuiA0gsi8XalTe78yHjTqFXI16UFyx20fO
Yk7J9rSMo0X9IdM7HEJRLVE3oHWqRowty6ZBCPqsv8pSaOnSh9PnLmmrHpJq5xIWfua2uZ8fOwa7
2aSF1W/b6mxcmQx4AmXYdzOmNTVnSCO1d40I9LcEO+EUuXxEKyMMUhEADGhnkrJpYa/ik1nPqdFb
kiGAtntB3IxccwrOrHTNM7N826Ij3CDmnlMi5zHlbKk98KgBOPA1lf3psAEmGZA9xtSMECCynB7E
gGlLFMb3A5JgVfGyPLsYHBFpx+1OMj0zifG4wCpA6B/NMA+P/hd0yjyVcI6nvSRp9Hl0qni1gnQp
YzJgmk6wnCC0wevFq/5AZy4PhGdf5EYgz+/ZQZsSfGQzq3syDfiZPkN23IrjhFknL/cWgSTgAzWV
xpuEvxFBwT8aabQKaLkfqhtLztxJ9mf2ZMS8owgh+YUlVaxSqI+h6C61yQPy/jhsTvkylFuSSRKv
cIPm9cNeCzFI1IGJo298/q4R8QI4WgTapnxfjlQlMpDhOo6br9iMi0ChupaC6/MbY014685N6rEl
x6fJQFE83fsKF4gyBmWOFpUia5EcYWFV+bzEwE2ZsdEgngibJTaqKfFE1vb2EZL9FHc1L43kei2Q
axapGA/r6ELAU6UCA/TeEvkDmYQIbr7QyUDc/wdhpspELpUnK25T1mrnEDmIENd8TjMLvf0AnkO7
H1WgXaC8ajR6hqzprl3u6tZLGwZMgHyC1dLHHpKSRNxtKd2Y1Xi9s6SOHjUX9qKOir2uXNxdOi1g
GRUbWpR2WFu72jCmR77jpU1qYDPrheE6/WuubO/AxkOPHg2/Gxg3I9ytA/CgN+gJmKmff4CuY//2
5gGaSg2018d48u9DqSPkiTLXyiRvJ/LrQIRofoh6GlVjmX7IixyAZ+fVS7j54iAcH9CapUkWMIKD
qhoGLwMKWOvNuGhEz52ml9A+QErVpC1OH+DvY8NVzerwT/fc/gNc5ULgVER8z09DWZJ4XA3IhbEr
igd9H8nL9gaWXfDHP2w3Q7nnSbhpsB/ODTw06mqoSJzsJkOcVEBoHFkTaLErwxqhyegXctYMcfsS
g7S0tiNCN0XvYlocEje7/hnhJuPBzFihS6Y+JavrTbw92I2ipwbeM8etu1SGz+Fxf8v7zeuQZAWf
fgdnCvEZ/H7tBlW0CL78u31FmKeF7dTKm0PQdJ9OrUOnItjUKhvEOcspr7x7LFj0nereQvtMvLUz
U7y11aHCgCDWinLnsbnlNjNEs2T0BGeJoTvSpOnvW3Y9RtMPbHrH7HE1GWMMWE8dcgzlASBpOI+A
B6XwW/Hh1SRBaXbWEnL7oD+dNATXfcMyIdKcdOPs7kBU4sKU3k/Fj2iBdQqwjYnIFP+I4L1rOGI5
6RIBkbv6yz6Run/5NToKMNsx/liuiX3L2yyW4loNzUVQV5+a9gv2yGNwhGzAp7jkXtZL1jKP2qZm
I0iyEPIKOCTMFOI8vcWoZO4TMXqv7vXC5hwM16DK3IRvKqtl+wrJ/XO1F3uHwlnSfBAqTL9MOfXE
NdlCUoBVyp2XwL1ix0ZtMa2kI+X9m8IPBbLZdlFJhPQr7pNtls7ZpNfUzqF6fTJ43RNRHLo295ZL
DwVegViUfWotBnEgUbAmiCY2HOLfM1QgPEW7vSXBHU/e9786dCLKjPsd3jDPdnLGwYjEjFdNWY5v
UXG7KklcMBNUMhZBw5dv5alyBs1Vz4osMW6khLgY/mtSEyrGH8v6ec2CGVbeYPbv+hgCKEjcE2+C
pL86K53qL3LH03Mxw2nQdKMOCZy2F5eVJ0Zi/LLIUr6iOBjj67QTkSWPzXMjPGagP2d7X4hAL8vZ
JyND22jQC7RQvzQRdzfqbvdKbfbxH3MND+dMiCClj8A2Iq5xzt/L60us/U6C7wAdtXfkUcH3/FcL
nieCQEueyPlSZJfpJcbYyGTFZPOOgISfFMVRFUZCgK/CfazwiMaVlwr1adIi+VLDP4NQ7q8XVxS2
kto/jMS+i7inULmKasf+1VtGZ1Y6f9m+gbqIoPwsMay2f4cTwZLkoQL51GXnU/ECnMSW7oJQZVUv
xJh4gUfqC7lrAElo6hcN/Ad4KLnQQ1F9LVCjvxCnaYcxD6+M6mgh2eezzp/oK8JYMmjsatG16Vha
+jrQdWgn3TNq0Sl9jHtOyGQslEIIKTLGrsIFGjbTi+bQ1StAP6SkEVzHv9woaE/HeJbw44GoMmuk
NAvFcdU7GqXeGtq2H/U+teSf1x253Ujp/Z0YeIshCDklakvl5+FCCiY5WY4a46Y7dcTOW/+7q7HA
frikMjxQfeXu/vYq32RSJIcfOx9CdrVgxsg0mCvqRcRMuO19yqfjKJ2FmRpNP0YMWxvpBrs1no36
Ep8XT1q0vhezvHaMTpbzDZMm/TLZ94fHKpdoNAi2qPUof//0h3TGZZUhwHCuil8zbdOrHt8kvQft
POf+lJNi6KHp8rAEseyV9Txd3CobyrhbXsO1KIWsCaFYlzSN11itFh4SYkknHe52W0qb6zMRkdiU
J74uLv4Rf7xqz8E5LGCTadlzV7I0luiw7oAW14FaFTrFGMODPMyOX1LgXk7YlkhbMzKQpedUd14z
VNxJLRn8xO+Sgla3ZEWA++0x0B0pUdYS1XrdkCX1ymSDm46A+VsmYAxF/3scvVTdbWnGz8+l1xm9
iztLlFh0zKtSSQEybICbD07E9Qo/4JvbtFSzgCZtTRn+0EAfrVEMO7X3ScpnJQpVSkWs+C2KH/JD
88jWkViqMqjVLmuAD06Rp8HTEq/s6jGo1PQMhWuX5KL+zQBZ1YiAQCOuIlzChtX5PZecsD70GpBd
9Uti5X+PJZzPtTc4icDJirIKrsNLmKPE3XlvQiM7u8UOAuXm4HJbrpefX2HKRO0tzJjqUPk60zlx
PHAAy0KprqQxL+uU88h151BaC5sed+f1p6TSty4S5H2LLvpagLYnuYhMbV9pmqhYBAWpxX/VH8bq
AKY8+A4Hl2yVDNY+r5UZK1LJ6bzDjP4SO41v3hzp6500ROjcq1Rgp7ahr0/+jZNpXD6o5HtHrB5i
5/JfZAfD/2FCeoxPtK+Ompqgm9ev5MBKnx9EWel0Bad71ZqQEuGV1nnv50wDhQxoiCl8NwkugtbU
ausOkq8BLpygQBfMNlBMLvUCz1sf8r+xhQSsVjNHwFTMt8GRhEBTrtTnrbLBkd2mVQbDfih5Czrw
FHUwHeBSwpj2kqClwYB9zNUCUlBj0J9o7TELxI4+bsAXg4gWBfmr/RGjSWbdhQ73Jel1cnD9g7UY
oeAWbRJGG/ZxwHS/pFT5rIPH6DAMABt4lmUYpNDT7xCi3aGeC7f7HtLJ9Ulw3tLBofqsJIZReNjX
ILKLcmlW5jxHXvld3uY6ByxquRiZFFsKRw+1sih7stT2T5L5QCIGBHdxwv6ITlpNu/0Eb2ZQHhzW
Abe8Xp1CF/kvvI60A6bDCfRPKkmukv9rzO7bS+FhVkznf1TThiWHBQvrIQwhCfS8YXpk7M/A7zNF
+dBc1VOwd3oUXjDynmWaamjeHUyACfzYYSrUqac+qDBSse4OkOkeVWgAD09MIFF0ooQMIK/HGGBf
etGFus9fA4JmR8+S8eqhtDGuAx8ITubTJIGMlrJMYPppG+qnNOFB9bvxXuCTBMzkYjfcQ5aHCTSI
jaS4o3RzSFylOmkCXibm216lCuleoXYlrssA2ys7DCwzB0ewlA1sjpf54HmQzU3FhNiaoB7Rgq1j
UqlCqgLbea/WqVYXB2+/y82NV8JdLPgrygMqL8gsPLjvlWReG5ompWQjfElyfs2shOhOowdbwo4Q
4bYn6wyD//TwvHM09cAiGM+eG/qqe/ISTjNNyo46eoEEJOcpX5s7wcp5IqFmpHylTjxxSnswdmfG
xkygRahqQPxiX0ewJ/nT44HikmyBQzeXan/jzGbUoOZGysEnwyvX2ujq49WW+uNtLzEms3U9HaXJ
DVo+mimAByD3bvbQiOHP9JaOw7qU37Az2xxrhtG/qn6WyY6tjsJr7QD44cC1XEYczeaEEoDUfjwD
3RjvhGRl746pWusRKMhKeyNha9ReDJ9Np3h3r1RItu7mm10uQLJNMZkYQGUb9LC3H7lk3/DlPj45
V8f3od06O+jHGJJZ/px47g1NIa5R1IK9Rn+d2rwAgCro2RXeIvojQ1J3GMFkNBSLWjCEIxIc8w58
dO0eOmPlvCkLmVDxKsFZaZmYWcaocoQAArvQ2XMAV6PObFzLoJj3BB3Q9/OXvJu/SBNZbQ/fr17f
RMi2g4ibA7OY81T4H501bx9xXTrQ31cU8sHJ7EbE3HOWW+OV4lVxmhGLdSsuDcMHNcyrK9xMacre
+23+EBn5kXnvAlZw04wVtiVZ5+R7V+2k59bHcEH2IlQsrwBF6q3r3XY1uBCcsAJ6MapBNjlIEhKJ
UKQIrLGaEQcO9RmDTcX1ce7+mOnizE6vHLGwYKiUvr5lDjGeBclG7nomPJbrRPZUhmszB2n0SL2X
onw0jcUA1VOPOZuh3paY3WjGuGUg+0n4JBAJBcmaS4M81VTze/jShE/8pNO/lWwsaIP8WST0TJKp
Xf1PEqrmGtoHxOh6CzSAzY9A5LiImeGc7duYYJFUMyJCACu43GlofRaG3sDVR8WXk6hKcFfEM60j
Q1IFvo7bxKTsMpVFr8snI7gUI3nCAF57viwevEFYMldbAcBM+0Eb+mdiampO72gw/Kb0f/MydaRP
CktITRKN313l+4/Xky0ryTbqhcOpyGDkzPK9K2iZOKPvy2Legag9CCGpXOHr1L2cv9YKh/URSbSr
N0jIqPYKbj45eGSAQOzL6N7T/tEysGcDXTtS9BYav1TTv4fGYvUsSCA3h4jIq+4iztb4iIEcv1R2
RhtvB/qC9/NSlgk1acAli+odI0zeLyDiNSAAPLJuTEVTB+WFquj4D3BYJ++23TqfCR6aYmhqUj7c
7LT3EJsMkDZlhaTKSFnvUsSvTcN/DpI0Zo2hO/Y8MvaLyr09s+2xynV85p2nVu0fqPYRJaUGTVch
mlSNVKxx3sioTwZUYnoBJzO7B6Nj196IMBiAhjlRoEU0iCkVg4o1fGt1J34TlLSx+a6medMNVta0
awGc+7pmobTCO9HytFRd8cIYnp0nNZDUAT3HD65cylx4rGY7v/9DBnHlZs/4kwjCJyUi5ybFBRBO
R8jYv1baomQ7WRNYti3urOF+5HYpv4OtwdsyJ6KbMdhNE8DskfQsg8fKZAY/HtkWFJu/tizBYTto
TfVnt545UICA9uosiHwgLL5hS2Rq4QyHYVDeksbVh7o6Uo3hLr7r9edHXFstKjR1gtV1LtUeZiQG
SBdLpbYSZiGxHapWxR/miyQIo79pZtLDPN7X+Wu+ycBIQFsZf7WylTCBHTNIvICv5mgjLmreFQjc
LOaCye4Y6B6NbNZQzkJE7tqYeEZPBOvjgi0pgCcvuTQQvUtPDtRgkMfS6tN09MvFd2TOnR+zn/qY
7m0a+hpqRbGCaU2KXT/g0HFDJWrlr8FfNgwHIbZ6J21ONe0iZsfl2Ks2/zYWjCaE6V/555xwp4I+
LddkhB0fR0YGYtxFLyp5h4mkZgJaBqdeAW7/06ibLBgNc/JwrMHcsOxpNJyErRO1Wt6sBDWUK7Y2
V8XUu/kvgEW7DU/fBD3e5jBtKQgMQQ7S8wufPdaHOnsiZWM/ui12d+cVOPqZGH5Nnhpg9Zw9RuSO
mkmsAvzQxI/NaLvijA/VRT+qOFuAGHHfkwtpJx8fICjVocaRAysoTcZekkE3ZOoyIPDop4AcO/m7
yhnmVxtm97cB8IgeB8IggKklbG5+Q6+gpfdkVUcoHe4uPwll3UpKv39W0zCgzJDQAwl2wUM5Vwe9
57szzovd+wqoi3qea7uahNneNL373Vn8A5g79s3mlT9svaZkIPpRxeXDYCOLPB1VyyXuJ3GW8/jr
tmkYVgZO76TCTJX41Ivy8fLVOPt/sJPSZKd7pJV51xFf34zBcItOXYLs5hVsx5WvY5D/LpI5NIIT
gkhZZ9oInz2dWolEbM8mdWx59wAqkBlnt1gmsgvM6ybOd2PaqFgmzVpu/G97R1Krt0eqpKDfdi1Y
VzaZtZFfjLXc56trFtlDYrZbA6Ujtlam7//pL3FeH0OxeXzcaAJt0XM6/0JYA8u75CEgi/iAECdS
uk3xViEkzB/vCcpLUprXUd2YbHFpt6vTFlw0T3sgzkJEb8jG5ZgaKDVc9lOc4CfzMb90C0687ywm
IawGEDPOoAKC3YCsnggR8/WTmQxO6xQ/rbBf8xRe6CweLEaHfFhfEO0OVT8uAAebbh00PO5NVmpB
EOWdSJsNrqw3pe3bFq4G+oegqu9HyRAQ52mEELOViWQK1LoTZJaWIBSMZjOVMuCHcg3k63SoxW9y
t1IzB8GivGcRhSCu8lol2Jrrde/Oh5Qdz7qIgRCqXrjq8IZoMyfm09kqqgISbqEgj6IMrVcast+s
OpCNyYxBvv5CL3rMf/MtO/XFHGCTxBmzE+Ou1M52zkc2rAiz64LCBs35lkehE5cPujKg4PwHNvRc
veYGBzIFp+HFMkefpyNpxLUR3n1HUyRSwEw76YXlzV3rZ4lY9yQirZISqLAJqx1Ecafy7eUNv4kF
JeaHEmEAywSfAF65MDiFJg8/K3/DCI+8jij7OwGdc+NA+JGhKIvxOFeUH6yGqvBWl+RIEUVqbvXZ
Aia2LR8t72XS8LorLZedEC9BpH1kC2Gc6o7DAUjEs847Ka4cUuwa7FTXuRZ7gdTFrBXI0pYqZnjN
JHFW5hE1MuQKweO0UXYt2gAo2YnaESkLwrdnJkwNjRq+cbrB+F3Zg9OE24p3aKAWSf2XxF41yxPt
ApeXUUuoEgQUZsIcLxrzGMcXXsLaDTqL3QM/Hp/snYIj7fBfHRJLMdERmX2HYzmgnz68ujaummCs
/s7amZqDTa9g/txW89MKiNaANsrJ0H8TdhvEWVu818Q+QCQ7YZOnOR5fpxbezcZblesdeYAKcziT
n8kqiCsXnVWznbgjqa3V84x1bOOqdptbOru+SRp2//sFvcEgXS+X3qx7UFVKbWPIYT+QMjSjJxud
nBy0JZbnBVXgm+1lx50WxN9E9lcynTp0WVWa3obAcWREoWSJH7D/HWdCL1vX8O/vhzQ6A/3sjHUn
1ov5T1EAQU/aEWUWYAIWvR1IpjcQo2Vh+pNQFkg0XnzxV7iGEO/VdNYYPQxNxa3JALnuEkk4W40Y
7SUyDYGf3GT+CoJkNlZqvrh+ITIXZeWC993T/zZNMu4dXaEOhOyj2mz9tWGeCLlM5LaRevtB9E1N
Mvna3LivRPc/i3F8C4aWZ0QWs6Wg1MBcm/vu6TLHXLXuyZ2TH8Qaz4GnhmaghWmD5LCl8zx8ekYd
ydcjTYhUR9PZmZuKxhG6AchUcrQO+/sxpN4hbxGwR6Yn1gaWrGtFWlTvFmgqMMby9i6ftGTP2J0N
NrF86vtOxAQC0FiM3N9Tb2bz2y/NZf4LfpQqYs7A2lGlNxCgZ7Wd+uEpK2MbsB39pTIoMK0uihNy
ZmErT/iSztaqndqc0TJPj2R1XZ5QP7vMzzrvGdKFcmAuQK2VgdqX2KVqGK2GwPQ8gYTEEQA+kdFD
avE/VdClcrcHbtGg8QJk01nXs2a5p1aFdBdxkGbh7oK7iL4RHw589mbd1fFhTbdGwgmOohdiDBDe
5tzHNV884bY9TbMAWhikYM2vW+M701VlpoDXWcIL7N4fJxLXdcZqt3rCRT/XqUkkS0rFr2Db1BX9
7ZAAZVMtcfdY0s1IHNuURyuzKpZrb8yuEmksm0vLMan4YwlvN/hj5EfgYR9RymDBCvo1izqRqv7x
u0OVuN7tqqoUPMuR/IQMxnWLoaQfP2QuwhX/7HGGorwpCQVOPGdge5zUAXl+dk94G3uZ0iY4C51a
4bZeNaBC0hbz6n+pDpIk8+6N8wInipIhcgmAs3F7wNcin6txRpccrfps28IJLwRP1iF7G/9fvvZJ
By3U0glVesuZaHFJA4ehQliGo85ucDMScomCcgiiT90XjB3Lc6xbx8Db1ZKB1QHRwBT72IBSeCD9
ESeCxxThBs6n8tzDwpfXbdwrbTvlnerTOYFgmUNIO/pZPOPyDmy03RNpJ/5JwUYEiijFlBLmFoXE
HjvyPP0GAzxbQFWepuAQyYXr8tRhKIUkMFsQ+FpnLuZJcn0YS3OFAbp2obn/FF+Tt8n6S/lVRkSF
k6O1FCnr8pzu7uP6Cx3f/MMFAVOhfYK9wxs0Zi8ChnvGrvz05Zg46t9mJEh0ITquKZpeLwVaSA61
5Lx0ai2SnJQ2QVTAPNX3XX1nW4LMHFFdOdHEvprF5TIuYGRiAIV7jGXDHL3Nz+iSKfVCDLMGkaC2
QAfUGh5vl+ja3ykWnfXwsXkJ6fz02Xel7U/Ga45fYfhvZVxXlPyeP9lzxStoled9v8LKKTzO53eN
joMHa6Bmji/9gJmA/szmJ88FgTbYWZ7fLgK+K4LlFPLIp7cDDkkykDR7IvFWNl/RPaVrUMuFhv6L
/+LEzIgmVq6gK2SWbTSfcipOR2k8WHVdsshv6KJ9oOV6dx5AQHmNqk8RuOWvlm6nkdh6GJeoPl1e
N1cg/YZHT9vrtPMT8cmHf8X/weMEeIVoDAm6vMj72XVl1QPQfaE6GuuuKb/veYIzjvmysfk/ZEj6
3RJOyibPG+xVCXMgMNG4t+QSNG8RTDojw0d04hS3Z+Ve55XUaL2ta+EuZjXwCW8E5MdgAWEQOKfp
ylOcyN1/GmTnmAeu8+sMP+rMhDrjb9izTWEk4qPiKCSarfZrFplgIh3tiPmjLdXq+xUeaWpYE63z
A/5Wom37dKU41NZi6+Ds5BUqM9f5rrFFzZ0DGn0nM3wnyWTluSHyDaMbGq1ZeeYNiE4bSFDmbsO4
wbiBxFxQE4tSzQmpzdokeYAo/LSPIqaG2rGFMHFbMUAhtYC2DRtYG9wo/gHZ7DlCfBGI0xyj2mcv
2ZazWJV/JICfIIpgMRuXiTXuwe+wIIXruBjb00hB6P2z/HfJi1MUr683LuM59ZRfyV9ax/GHHKUO
To/xUWR1dnCrQcV9Zp6SCTnz6vq3ME+4iaCA2llUnPxfUKRWrPHxSvdRx4PrHFOCrOjLyyJQoCyD
QD40mNrC45ptw03ZKkCOeOQuxIzglnWQHfDKy3B6FHibQmbJQKDqeQZifmOXHy4oB77SMe37WnrE
IQs6jR0fJTBoknFiNBuq6xHrvYMBxtAJhC6vjVODo+dGpkmHX04b1/UX5AlHjbVQaJb1HF24bTdr
ATnnB8MzLuBe8xCFTKOiPGhP07a7oe0tGm5Hs5NfhwADEIiqR9h24Ud5bPGvj2Ybdiewb0ffI5yJ
tRWXYZVflH71fBn0REVK3sC0uPJtQY9OlDR/RzteCNWs8XPdL4zXqJ5ZlJ/VDhEJlsibB0P0KGaf
fRV3hrZSPVtnozF5pShn2ArMv9xPcL264Zap2DMVCr2vVViJ6FQuCnAkenWht1H84GgMnZrA2zZs
T/tnz5E91FUqECidiiYb8N52Z2vHavcqtwuMm/V6/UYJcvoGA3MMG5ZxfDfsBIvYC0lEkzrOJbmZ
oa13b92Scl7TM90HC0x4o+Gz70hNewVlAMryixvJ0Or92oijrXaQSFPCmYj2nSaN7XLwj1vawEer
H6W3QoO9i2Ok501JZtTqN5Bn0Vs9unxrssdh9FCMEF9cv5IxwGRD4i3qsvuT2RGpl5lidASN3fpn
fG2KmDL+U2kp37Q5A0VPM30EiO2o8AOPPA/oGIXl7lCpT2c1ZFBvUs+Bacc1nidXHY+EHSc6EU5i
8xBJXodfTYWBF8PIaprKj41ZqsPX2thywuJuvswlImcEIevEB2GCQA4sCMaoS78WMDFzu6k6JenG
IOnt0z79eZ4h2iVZFHYW51Hs1p0Y6o+6IoXWv3Ybaqt6/+wjqQjN+E5eiFXWjTQ2z36ru7VoJs40
acdPbuFg0zym2LRdelovah+Bmr3Q7DH3TjlTcPmP8C82bwuP2Xy0RVJ3kM4MOl1TO1AqEaIV+3zo
x9YAzEOmWPCz+/SZY6cmRlDmIQZz4hw1pA/4GTQ+O94Y8XfF+ycAQbuxNDCWI9VVChMc0seQi9kc
NfYX1DApyexJT0xQy4ZeINuNy1vz6dRM47da/RU2rz66BmL+LioZtN893c/X2TUg34M68muDBLoY
3koRCW2XHHqcMUxZYkhjIPFfY80JDC7Notq9rifGBp/GaQYV9/0iJ6FAsVpa2jWF2Mmt2on1FE8i
UzRqTUKeD9ygJ16NZ/NFu8kFxFhS9D+MaqQUdi1w625vnK7pwCT8q6Zjeu8cDdk87UHtQVcv8fgD
a/sE6WC6FVwklG1UGuSA/EBGgcoTY20uyk9AKzuidceMd+6olp2aFk8C4UXkpOlkRidFvoWJEBMi
55kZpshAEVIELh8csSx177jPMS1stGIAb4x8JqlmcuSyVnqQQA2z81cB4ubEuZ4ZJFLjrsatlPhK
cCJzOIfdk/Ct2JxG5cl3NZDloUMhufql6g8mlOfY6uBFkeELYh1lrQne/nFWS/tVcMVWVBQXOEMy
PLa2eMl2Qx0CAxKInViHsfd3Y/3HTVLeB/MDoRNIdCKURkpMbX3JqBy1oGWIhmWOYDC33HXQGHup
HAl2ZPxe+jErh1CxhUFMBjnN7X14TOr0AeAFNtstBVMmspCTeLJTFzF+bdO6xN1bnZ3S34rq/jok
yG4c/B7tKUhy+CPXR2KSoqMO4MHqIeTHg5G5JFj5hqG1fUpBDBXSYDUKDfKt/Ub2h3PzKxkD1g5C
o/vOCcGGmY9pByvueab6on/+W1HrwL+JAdb67FIuaNytm8r+yRtk8r6Qki+QOqLa2BrEfG/US5X/
WPo+k4USDJgsYJ5JY6zPrtWb18Z4kTjg+yyoWyKMUjpw1CXAsnUw8VQGIjIEVUqBbQ2vfOPX48mr
csSAGJ9uQQkt+JH2EBAwZjWXjW1f0oqEOSe+BszFLdbX0f/QCBd5FWshXuLHt5biYRTBOaAcbHjG
WbL7m56v6PzVsOe4GqGwbObjaEDnZ1NqTk1CXoNBxv8RqyTH/IE4JnX71o23VUlbxaZQesy3faOF
qhwNCyqF1829ppQrf0k1DbgLXsIJqF1o5r91grDUPkb9laPPwO575NFhRv2ZgT/ZztRJfI/m46l3
bDvNhIPzl7D5YAwu5sjTm+5Z8oyqqwhaEd1HwHZhW+T84Kwy1QZdjh4BZGOjva4onOK2/XfFDIy3
xxrLWs5XI+EYeIgSzlgdZJRtZgjAVts4kv3dK76CmR57jc5C+WPzM3B0rQtcQemUpvjVi7ROXVZQ
kAj35oU7hfooVl4mxJ7FfjGp6jKzxuJQh1X0UtbK6MvI6+NNII3QtCYxUMxczoQQSXtfIXdH5vQA
nDK1h+T0qv6t9omJXeP0vt5bFhy3feHrmmAt6evOsdS9InrWnJbMJuGK/B0UjSXz+JVtmfVf4SVT
gH0CpvhaFRvPMDI8n4mOZAjVUSHbtn/R5vvSKaWpIQw2Sy1Jkx0Vm/OLvU7PYk9sp7sIZ0fOcRbW
+jGH69PUlk4M2Ro5eITexipZ9Lc7Xx6xNeLhcDZFZ/3YuLD/ChURJjcjjX16/ouGNTMV8xgDuKDI
eQDw5zP6rYyqEStZ6xmL48i0BgcAFvFhYZQQNLawgY7Qrk/4oRf38/pOkavbyKMJ/tPoFYCXhSht
gGC7Oma36SamkP7qwDrw95+Z6FKK+ZMpNqT3rGAEwcejymcRGb6/MvzqEuQP2oT+qKtHsNcF6SUD
TXC0c39bqoBxs+HeMUMFtlA3HrqA0RDyiVoh9c/PuDXZB/egVTNMjKtQvjSZeFC2n3tdrc+0862W
KwP4QpBAEu5+xE85BhKVVmpiW2onIUEP2RbRkT6+dzyDzx1LTS2wQ+cNtBdtdMLKaPdCRLAX9UtG
CK7Albou5odDcJPbIUGVcK6RXJ4kssoheyNdj53Wtym+qsI+7dri8QGRO9rZbFHeyD70FLzFVg9+
MWrOUAVbyuwi4Krve4/UbHtuAJLkFUdx/jFfSvdycCs9aaERGuo6CAD6ux0/U7lDmOvu9RXvss7W
NTVQw7p8E0KyoDSOnk+Gh5Yjms9tCTsy8YdGRNyNXektRM/8ZDSAt2T89vQLuqn47rMnPxmMhj1q
xFSMlh3HvaSzutHJ8VMYQf1U/J2x/uTkEgrdpESY6X62sOY873eicR4t2jQAIxYbOEYJIlY3+FN5
NVOfnmbPjCLz8wJDNSU5CAKKUIe+09d9f3640xl1O1jmT6p1D9FEJKcLAACKBJXZKgECcSpENQVs
XQS714icdIk2/nh6zvHrLM4O9WyLlrVHZKawfJhVx4Fz84drMFkv4GK/wjwCGvXKsOH9cnDlDeUy
P726wrGTiNcW4N+cqHA0z7Rv8CJgeUZ9jjsxFCEh45uP360zJ3p8HH1RoYUj1G2xqkAycNYakbbW
1Hq660ZoIudfFWGXTZzJnlTmswxex4nH81G2UIOvbTMPpkF566X3Q6SUxu3WoxQDPJrQrK/VVd9R
kssNfvKX/MxfDK2x8CDtdzkCX6B9VUKT85ALrEFyTa+kVUuS3NdweU6R5JzRMFexv42a21okpdIZ
Ei25dOx7SSV2j8gutRqi13zXVQXHptM/hjm/UJyq+TN51xhxStfNccTG1xyfMXlHVXU56RKNh7yZ
wkAJ8rOpYvjMpMEwdYjn7vs6B2USDuBp7FD72h0Efo172rOLfGcyCFfCejxUOc46T9wX4M2gMduK
yyucS/qlr4632TgTsVxaJezE9TKBKybStJ+vP8+TnHioHuHslaNttVqhTqTz8+9+cqdT6tbLVyEA
kUOYRAh4wYsubI37mE9Q5CMsM6ICrUE9FHAk54Ugu7qoC/TCmx38ZL0oPNher/7WrUGtgY/nA+QB
KRaaBg5k8GLW4c12eCgbPN+OgD6vnPUut/s5F7pUXypEQLCPK/nm+AfR7I7JHysMqHqs6P+wayPd
Ac+x/4CdiiAwIzQ+lEJz6QopgUHdbkzXA9+u1y5BuI6Z9xd39BdmnuYgFAn73Gpq72vHd6ShD6Zy
mN7Mgm2fCzQCgyTS/wmvamW0heW6ZpTkcPJsZKImy+td9fk7qdFJdVpPjbd5+MlzS3I8fB2SaQ0j
AIdKqg3nVfCjQ5FHYF5XGr1FVXmj5QK6k85HziG69Eb5hV/bVWoBvO3v0LyFWi/8kxmPYaSpcwmH
SNU1dnEL7wn5KNUNwiM3D6t6K8KeyFoV0C1zWd0vJQw/TkTQDJe0HQoJwRzIKbGI+UnY9o3wpwVg
Kkdl+ey7zrzg58NuVUCQlnJ+vWysP3kz7RddgaJ8l9gAiseNpojHPjBAki66OG1+g0C3UZCQtud/
dLU7xt0nuTbZ4tTIPLIS2BsscjvrXxx3pzNTQRkmBiN1Bffp6GfutEgOkvGX1TW9dHQklqJm4asO
94vlJir5fvBb0BW9PT6tZvWsJA9P2ALX33Vscb/cUqnPi9TeXf88Os0j6hgZYvQxZnBt+j/WluZW
atvqkLv8BLlsEC0kM9nkvCw2WZd0vX+TBsrVBoCpWUSfNNHAlOSJE8FSFV94wqreLBjCuF0WJTFA
Zt2y943/7f1jVqflLhBwh+Ry0hyFlauJmEfUhwrLmX45nkO76CD2nlOV/95mpO+p2UUZ152oXpuQ
2Qp/XRwaLfiIx89qzXe69oovvisyetEa8kqtYvHlrwEnsTMmDISObRsNKlUclc9jHW07zXzbTbvC
LSikYDgwqbluwxLqqoNjfFjyIWdpMEmbSRwh3X5QdNv20rpEHLTL84O+szo+LgFgikAP5SS7iU14
ut19qyt7YQPxmfpAbZMwIHhZ6HV8oCg2rmf+TfwTR37vxovLQ91bl8quruCBK1lStYXYr+RMSqCg
Vr4NF6RgwLY0FAmbgyVf8lxYRUQn6gsVaUX84W0F3YgVzKSF55HPEaRD8as7II0UtAnZgeWS3gu7
XwbfyMWQoJatuMzoDl/FKBS8188jIOOwhQSNA5jgYZ7nWDL210ogeYE2HK4JcD9QIJLZueoFOTTP
RnzixPY1gqbcpPglnWJZFHELap0EV3rKypryG0wObJyy0F3vYtOxIlQzA+5nhN4/hpdPCno14rdX
o6N/LPz0yVCoHIno2Shnnz0Y3pYKOXGtAOERppmZWNP/dvE49UUW+mSBOyq+gtu29IQZLLvO+0kO
9F3oJ0PZHurC1pyIkobH1Cs4PXsAkbxyHSvwHAFPJ3J0nHYVIdmylEvadpx3A8DtDS/GWoGzQUED
XtQocJHEHfCDZfmfMSppZ5h1SAxOAGKUnEFoxSW/GRxJxuCGDG8Shre8bn7ggle8lqP8LFG3/upr
zatRoe+0W54HO7ytOlmy93pJ3uGgWPDPaEP3OKCGFkBWtqVRRSUW8ZI0FXCW/Nr2IcMSwFe4JM1j
ohJoeB7M9etHubato6fpDZopbMrD+iVmG7UTA4UW3mcGSYgJmrn/iFRyBL5zEnsMnyuqeUU+JLGS
CUbL8MJC8P8gzceYwkUwL+Wl2ty49TEkvdnUFzgfMBvD6ryP2SyltdSYUrDCaT5ub79j2Eu6WvgU
nxyDmuZYGAk6hDLmhKR/AkgZ2RD7FY4M3TCSU6ki/R+HHLtZ46Y+gwG+UJiHjHU+ATf6UezEofiS
59xE+skxtR6P5TuSm6x8mMmGieFFH0SIxlVoI6dsIXewQWrIKyQ9lAQdGVnHUwUpRPXd9oMzTbC6
gAzglpwbhSsmnpIgh60TqzJSViJdp0+EGkD52m5uZsGuhnNmCIdq1Q5c26FPWkZ5YHbLIhv5Gdge
pYUEX5dYDgiwQNDnuid00YAVQQ32JuuCFfpw+AgJk8a+YXI5gnzYp/YKRCxTJwwnyXAM9w/TLEgC
D/CZRjGEeIzGAT76QwCZ9o7dY40MTrxN30hwszHDGNhsVzJf6jj+p8Jpj8Dm+XcvjMtveHkUCZ6S
/tEl+OXUxskRI8SKTemzYHRsAeR/yms4YjWp5p+wBJKPFmNnVSHcyWpY3KF//EM7vft8r7X/r+ya
WQtPBMkPaeNZphHRyMLgOpsrjV9gvSwKjfg3q4AWzrlLcv1E6T+3WGBtdrv3m0xulXwLGVFdV1DG
M689nZ/PF7FNRguurGszymItys4teCh4WXAGO7cvo2pQfo87m9z4xtgJOV2uuKdDP5cFmaBjmqIX
a23L3FT/u7j8xTWcQ0A+TazRwJZ1UWcRc2ZIj9S/HE9fPlzpPIMpubsVzQPf4pf1HfLVg0VVggrD
papqVZOYbX8DCozwDLj+PdlXp266/SX+hFm4dIFsx2iiR153gyvgQ5/LTPT/nj8IIInkFiMDXl9T
GUPxZp6jUmjFF+7jGfE7w8bX77Y7tpZYJACfXbJRlAFu4q+RD7lJCSh0vKBPj19KigCOQDvTNZWC
0tFtDYeFFPwSGuk8bHc/ednqSmFNPVHCR3czMTdGPy8jCZtZSfhmRkrz2TapbamiQkCDbNfclZfT
d99YE+C8RFyP7EHRLl7DAWT6IKTzFIAOMLW2RjiVWS/h8vyUkytNRjSA3qytu4sBktrzxIL1p1M6
pasj3uX2bdp2aRIqRKhM4zzKTXAmh7ALzlWnRXHJxkNuWETUNoFMiTgYNzN24avyA7kKV6Xgsot4
7FF3isz1VvJMmUw71w2q8iUsq56+YECOmsWxbou94Fz2V8eLKc2k4RHlS/40uF7HVUPYkXd8tFxh
J0q553tdCxvGwMaeh+1KOCC4cVggwfJRLlcSVHVKH5jmBd7ivEfnWV/JfT4aFRqhpkAQkXavC1IK
jNyHIsWVbtNqjsZZwoAb8HTotmQUhPtREQS5w/HE9O4HKY9dS5Sucu7MZE+68pqUymAOgXJV3l4E
IlxF6p4u9G0OCMVyA/QJZIo/bLSS1udh34W7vdN6Lsu+iAYVOPEttsXmGEDWOjhNYh+S7IWn/99Z
rgMLhmYORI7W39oLbEHxGJMwMOdscKZyzDF5Gli5OOKY2WC6TptHGi0dUcTX/jJdxCZu4dqXJYO7
NGfMhHG8ncKY2zB4PFfploADYnj57vIPVhViE5DU59It7bCaFtQUJVwDetV8qWlZYGB4jcxJlecx
M7mUC9agnSpeSx4fJQ1HUuybat9nwy93KpVjg4MX/wuUNsb+cn7ldXvctYVHjDdF8g30TwcGYPaF
KT+WQH24xQELQvLH+5sA3bmQJPyopSiTpL5rbCvFqxv6M8MNTSGWf/t7Ib4Ap2N2J84Mr2vgUThS
lNRLCfqoMrBaI1XyQgIQbSN4ObwQ5tZVHHvkIGLgswXAiHCLA+ceZhrHTMdnt8BM7dq4e0AnaJzQ
mwBaKpi+j2+J3ZFLt39fydj2R5DSH1O7f0rUVbLifr2b0Uh4zSujfyUEvEjiLlZGgoEKiXQFRXrQ
5ehPGWFZqlr1rfWuH+/uS7yfUWExnCWW8tS44yCJWPO4ALlZlh9WnPzVkKXMFhlzr3e45THaL6Vn
lFpwt9b28UGoauIIGOKgIAhLFhddg4ZWQ1VpxdVeHBcuJlSaU/WVzI540DyOOIRhT/3OGDqEgdzv
nMsjMLo4E0FB/SsH/xQIjn0AAk6ZSux0ckF8VMCid5H2V3b22XuDPZl3FvU3m1GIfZ9fzPy/8zGj
SSxRxgxNCeMVgIqz/iKjqBTztP6Be6GQ7qznelQmqZE/kfeYE3edcCvnloFVJb+9+g/NnM1lE8Ze
LH3klJmBoFOHQSqNInLo4MjSBSJvOfFtfoGDFlBUovhO2WwT1WKupzsDzWWrcVJ4cdMc9W5KR6Zq
BWZXDXR7fQY7DWccLwe0bGnvydKMKLsvOyS4SuHrMy1mmpz0v4xXOAjAnZjsrava5fgURY8MPaAA
Zt7sNLVMvOtdm5K/ro1qF62vhNxkGkL7rEqXUdjFnPUQJjuB76GzBF0C5x1XLEZuwiesdbZqLJ+a
43DcpxejQDmQCCvBePl/FJDRECrLNrGECB0Q9xAy77FVirqVM0BcIpJyOkDXWJi0ZMak8EGTSOBZ
u26NfiJfiWAZpwPjvJy52dh8hCppplxzIdt8WJC6UwNlnsowRrQgkdfFJxL648zNQ7kuIh5+zWmS
jI+gXjuYosPbx75MT8fv/hV+B1Q550r29eqYniYhXR3dcoH/bBenaT1PGlIJMZ39baR5PNwoRc2B
MYBf/mOLpLtWjzQfetMbMCOTA29GOuOwIAZl0Ey1h2Ya0nsH7tZxTs0vZ+v73XvMkS9Pgjhs/wTW
xrM5sKwrweGEKqony83T1nNzMkzDhcfyZHI4S/tHzO7Zvqr/don9kfB8yfzwG/WJX/qQK1zBmpgg
AfSyUmnAKOCy8yEZ8N7dFyzubyJ3RLSKlioUop3WgZeVko1p7Zd65daKKGmMRUpbL7WtwvtNGkBH
Anv8D+L6JZkR2l0W/+hGpc89pY21vO2sYWNuCOYMKpEFE/oMl9gvS3SNJlEfjp4Q8apokq8ujKt4
c1naYBOzxeTdGEqy1zZGMwiiDJuT4KD8YAQFDFkSeZbmBhdU/kT9ZbXqeMsM4gXI8wiJlGctKkys
RnuGPGuZ189WTclcwMP96BTHbOQDYo5qB5kmL8LVHz/Yml0yCt0ss832sRVCeGomLcGo9Ghse+XJ
DnowtP4qDYywYPOhuAf2CEe+WMs/xkW2zJZSOYEqXF4wiCUvGEb4NEfw/a889Vq5kLHbpCHweo30
zubnBQ5Yw/zMcz2N/cG7/DXzTUFVZo90fzGHun+eaug4HxMyG5B/dtb4Vzn5Wr7jfSJB7XG8fPZz
wNILlGkvAuMPiT8ukONLbHHo+YJc7Z+4SoXaH66XrmOJ9mtYSqB4SziuAm93UYI3LsGx3DyiZaRJ
unh3TDwmd+gKMPZKVhQ1z/nGUid0PzbcNJA/JIL0qF5p06oIirP6mO6XtgUvbj0KGy3MGthvtVdS
XKqFR6FaicDYJO76XusE621UDSo+PZDvknARajFUFoOZa4xzqR2k6whIrjKv9s2mFVV4sfKpSg+U
Qu/9qs58UhODqEhXVf5Rj5Srwgk4z5BRn/JsdhjLtKqGBqFhDoGvpbR3Ir6jhmGY1/lPtZByqCQs
83NkFgFBf+qS4/1Pl3expwFw69ecCzKCvs+rFbb8XxBjM2UuVQm9Ldp1HRzGaiTz5/5nuo48gK4H
kXytRWOYlZ8XP2flzNfeowKYnzjj1VEv4NE7gaHodvYgGk9+QpsFffdQju4kYp0B0p7XXo1+BFP5
b1ZiNVGSIujaB5FMKgKmO9L5ArcVYksjC3YemJhuGZGlj8paLwVa8P0CPeAB2Ee91ZhkYpx7VU2g
rAphcbkKIYNgTXhHggyepRytKSvzicjGbuJOssffpWqmdj4oR2Z2/40Irwc6Dpr8veMzQQg3MoWV
uZxHLkAXZAYS1mM6oGwspWdH5EiYFylOA2r6AtmdOIdCsPPd83iQUxK6GCvdGiT7assyo2Jcs0DS
wqmpN6GfMe5u0XKI2e4EfjPBsKsyeV9siHzWTWPGNfEZKyYsWOvDKzQRiVugg8uHfE11fSXP9/ym
R/ys7cP7oxbdqXXznC48zV7ODYjv5HT4+VLk+tlNQgF6xV4u+DHLMR5HqoMIr3JklPmKUesLqNjA
wJUW5mLYYyuGzbonVAw26UQAvaeYiBqWLLA4gUfoyAsxJSSHLXfeeMRgdre5suW8bTJ7ORwRsvDZ
Kdp+WHY8M+nvzjTcTDaQOpTQ5XgRqldGa93wgTjOkAbu80t6dddOuOxq/rmzYaC4noQBxW7h5fCu
iF5P+Z6fqqgThEtGkc3oK2sv2Oku49livP8E0uamA51jmYowaX/ot1dvfCzCGdXmPz+F/brorGrE
DnwMsi/UxUd+sfZ4EfQUW7ytJGi9uZRd8XD0iHi9haPkF4kvpAwEFwIvB4UATXuiD20OQucIPtPw
Xc/jYMqytlKTZva9yr8XYPJxAj7IzbLj4Gx2itoMzAVhge9j0fyhJEx/CTWOXUeuDtpPCuO9Eoqv
Vs8vFJm+NMJS0farUGm/hUEQoUN7gLtuwnqWL4owvH5sJF1PoHg0QfSssgCQrjiKi8CTegG3+2Mw
oBZzMzTih9o7nol/3n4vuorkTGIULXU93sk91WObXBJnnyJ27ZDRbwT+guNsjBaQkFhodmgwCgAc
K5uvqpFdNTD1h+XUQO6kDd6oWvOs3Fbcl7euNOxCW5MzW5LnKMyu/4xblNoTLsdlBbJKm5UaPlvR
YFt1lYf1I+C8ZbGG/78Aiu+g8ajr9R+2XSYe6ZMUIRIp/kG/6uilhN0home2N5aQAi35hfnHgKv/
bdC0CLvmaNS+4kWaAyYV3/ZMfohg64k7GpWgLbTxoAuk0UtQXabQWwiw6+cQXWl5W81rX9Sg3f/u
DMt1OAjBFj6pr+tFZNhB0tI3zF3hZETusJWxW7QI4fBy1pLb6A53ze2kekF60eoSM4/wTByruTJE
Vti5eSQLLJwyeocHSzMsQ0eTElwfWU+TzSDixYV26GwZ5lb4XIjshWSTzW20D9lrNeYHWQXR5pJ4
xkYzyqkWtq6eGyY1xjuLMgtSFsEfljuU/peDCGQA53GR7ZdofUoGM37hY+H0iqteS98aoCt2tojR
z326dDGnKij9K9KBcG5bVa4NJI5KPs08SmgDVKIS1/c89QCXkSgVREM5hWbfkxL2X5CVmWqYWrE9
K+jk1WL+hjGrkSp+qk7/GbmgTihzuFjQE0os7VbYqXiaDL2y7oaxp3hOYfTBTHdyc1wbpySU2Xca
S2HFb/ZTf8YWxmHTxMY04wNJMEaUxcQ+bUSsFvXOOXYHwBUKNUMDEzCUOJozdAqZ5hhQb1qfV1vG
27YBD8/TRa0SrFkpIEBWD3mpj4qGPyNzpR+9en4DH5Pauotsj5gViFJ7gT7EUMCxAciutDXeLaS3
V1SazzR/QmpgKwCD0EcDDmPF+EHVlCMz7pc8mQpNZ4+pK9Q1CvhDJu/8yyCMdT47rLDvGd4fKvYr
qp9ODcZwUtrBXj0ti6UWG5rI5HbMAVfkM9LRA84At/DlUDHcYvFi4jGvnKXHp62qKDYT5tU6K2NB
96yv4WnsJUO8IpovLT9pZPR7WBNhcKRm//+I52GfzIR0AKZfr3L588hyq09UP8yC874lIBBnoZOF
WODLPZdivUAQxkTlyTSFwPpAC13YeM0hfy1TxyqNcELKtkHAzC0Q1CNQXGwDHU2zo5BA0wIDAkIE
ALVlrNuWnnd/OzBmrrRQWaLdBhkpvAhxuB71EQ87ELlPL1eqNLkxx1uiI0vnrdwML8m6r0uy+Fj+
BoXDfijG0RHIx2XSdpF0G/pkD/1bG9WfI0r+2pH7ZwQ5vBF3x1eO/T+ewJF0nfYqVPnyD1Se65Fq
ICB659yRm7vmpKc5TUX+JpJlxUYQJGkJ4N6A83wteoF2cQXW0Qoj7OubiUDdqXCx+rimnML9CwV0
OAg+bKbZnUlfHWs56fdyk/tvtC+nx3mTZms5nwOPr/o0E3WevmpiKdCxKze7Dv1mVxfLvJaf4hR8
VxzTwEvKVsBUKh9bloYXrLEexsRFJiyxDdKCHe/KxwEdMVkueEhakloXwYXREVIFVPOM9vNX2U2J
V9ZN3L9Y9sAWeFWSiyKMi7mwdXtpI5zTGuAOCf4XFkZ5zXbWAInLMg33RIazmr1+enNCxZ81nLoh
QuScBa4vpoD0jxVLGIuo1k0GjHc5ctsw2POslUnIB3xrQBmMzarMsKK79EGRRLaoMFmCLZcWND+/
wbgCKvG5GLQQYJS/SIJ7QfAGb3GOn/7uwqJz4ZU/dYjJ9QGKoKni4eLMf2nfmQ68kG/QDAbcExgB
Qf+CjhQ3tkFA0TvNa3jwKffM217u22GcxAgBxnN+NW3mmIkATV653wJRSq28RljijVGFMip4uMw7
h7xDaLnXx+qEGcZn4UFoN2XkvUhYqWX6d33BSFQ5+XdFznTqaPbPTo7jKObXWm9z4i0GNWQY0lGB
rrLPeTFBDRje6YVwUvm+iX+RovTLecAn6Kzh577F8IxkKUXXpbM/spUOiB/3SWzMIOtyKrjex4G1
jJClST751LNvzTbUfGef5sZTzlrS99pUfLo/vDst0+0i1/1M3UyXHBDdqHzkL41g0uimp9/wsXcv
mZ9kbsW8/U1ONMSDamP1RpC4QqW7zOGFUNAo9lh32rpFbn74RvK5U3P3wCPO7Rry1vzXZ1p7oNKQ
FFgbrCE9j3OHstE1qrn7fJ19vwKGoZjj8rLhd8x+qJodb6Y0Ut9vPAmWS/jtV5PjRb5hALH0/OL7
SbjSwJ20pFWmKBe+jl5MWOFgMAbu+gnMi0dYOxaQW9GJqcpRVbFaX6w7kO4a2hGXVE5OXCnaF2Q9
d8/EhAQqS89of4NrDf4LiF8io39EKWqpepviiaq1t3X9o+VMqbHzNPTHkgKAB6tHAri37YRc/Lo7
Pssmr+8Nn2qkg3gBsboC038oXUfdmO/rprgSIUhrbGZrQhKibsQxrMz+E7LzySIOatYAmab9bCBf
z12RwpQLnx/P6uezsOjJXCvPc7eu7TJmbvHstuG4bx6Z81+LeGh3P6BiDZgd48X9f2HoI/qIF2DS
XWjrC2nY8zq3nyWYZlPiZVF5yxGmwYFzM+X2FSxRyTNGSH8GmInf4nKLSej/lR3Nxuv/M1XG8PXb
W2J87DIUt+VJLSn969B2aL71h77HDkIVatNSroyEoB5Un0i5JCMie49aV1yvZVgUXxPBmWsn4CuS
YQuSzVFgyMDOjQ0le2Kh5ldiExzF5Whk/Cg5GxtTPX8LzDOV+q9JGOIlWrlrF5tqAGyeFv+VysdH
6rUWKmKNk4Td53bJ9QE4nbxeQLgyT+Oiorm7weZQNU6QBXhQfyzTqt9O+d2xFe9C7MsogL0qh6OP
MYBxtdeMo0ZZumfAHjpNMEcmuSCrMVvTYBmNkgUpQxNsj027B4dl/fQDH5RKRyuYKqCyVQ3te4Tb
VvvAjYt2bf1QMmxGkw5sve0fdmKN+E1cYIz3bPZYZ3sw+u1rXQiMQb3fMsGBcwR/hFpRoNrWbf7L
iWtigQ/ww1CgB+aTIP617HjBGpNadH2oP/RmezPVPS84lrnCJgkoNRVu3gy0fjutjgdow3SJRJfL
Fg4CRmJj/rSle1mKe+sy/h/Io7Mv7Xc6agjbB6GtE9vrmPF0F+zxGURDnOmhWrA1yatcBCvQLhh0
Wmo7Ku2hJNEkUzFt/eLbMPWtDHq7e9xvVJvl0w9kC1W1sUEStelWuKlnUOC97So7VVB6mTAoAu/G
0766rPWIS4rLkA2BKLE9urU/jzlQFPb3r/V2rRlm/zn1HwSVTc0mVrPClpma0HH99K/2eiL5uhal
5pfXiYK80TpAyz5papHYcW9ns6LkLKvN564fz1DCnKPMy/ilPGnUT2T78gAWiC5rJnxC9Gk02M/C
Bz8sELfSUlkEOV1pDrPz31bDiHP38yd1QB3zBvbzAWy21O3t51pzfYKDQpPuOEmzUxBR5DaXjByb
hgh3sOJhlWF1ItPnjHVJHyzommqzlzWd58mGokkPpHYMdBy8e3KSAT5n6340g7NJUCT1VEJ5WeC9
TFhPvPxw7z3tMEIcvY9K7vBsA0p16gfDt9JoZJ/BAzdBVSFabv1egfFztwRvi832d6I5zZQnJ2xS
ixvs1Oq5jNYKJdYxG0MNChdo/3lmQARh7qobVhXotuLL/bwm81Gcyc+5ChHNJ1VsMR3YzMcGwLIV
8XW14Oa8TwITnNtQdr25MmYIIuvCSD57QOt+6ZwyvyhJBHDJ28Fr/SKrYU5khmKuIIZbvx7NVdUk
aNZel1sT0YBCEtAcetLJAkDdtrI+UI+oBveNSxGeUB5w5xZQ7I5NOVJQdyfuyOP1EBJ2AGhPESCZ
uG/Y8u8ciAggoDphpTV7p1Gda/Yd/zajVxuuGSht6zwVQpY9NVVXxyALoVuXE/ivJpf9W2AuH3GM
dUh4MnSHdibL198ShmBGRd/ULpYICxYEadA8apleVhffkaMbEQn1Rf2tx9WpLBH+3W5nD+EV5tSd
R3lXdSuR2ZclD/moW1sotarGZfMUJOq+olcxMPE0j3UPNRAoFyG8jOCkalKQ6aUeuE1BNUPwVpCm
mPpdhCJszwvVD0MtzZJOxkb9qjRgSyOF+PtXz0p2WlFsGXq4hT5W/xiaov9NDY8gDQsA84GnS73I
NAR+qCPkrO1MWBVRrJJ3tV8YzZQ+dw1f7NaibEk0uCqmRfzXm3iQd6P3k8iQz2ssnQYBOicLyJNY
YlF0tv7BIdSVzNDDLVPC3wAQl7WI7LtnIUUfzmPTN1+TVGMiFzDg2ZL2MB9Y/dbNkbvOr4D+KaTY
a8TE+EnBsZVrAcWYQ58myyLbeVAVvj8yv3Db+FC0QtIf1ruwRSLhyiZV0e42Ns2QzW+evJ1y0QeA
6Uvh2UKj5Z6z2fFFniPad4rmb1qrIE30IQZwBVnE9r+MxcF/KZe+s9pZreBp+oGeSxTWGYGjmBHl
0cIvvRrw9LUK040n3QXfC/FZP3sDfgc4XQo/itD4mer02NZTqg69NFj9NkvfZnNAe3HX1OC/Qxly
pwGRfQqekAJAWHiHZTG67X9/4VBVREitqer8FE9DVfd2+XZR/OcgLgB7eBaEepJ/qH6uZhzeQFJG
E8+kE/22oH9OjnFvL1wxXQFobvQ5uWtzTrt4eoruLBlBfmIznl2tzrETNCPhj1BprYk1guRbpM/S
oRdA82oF6QLnbCW10YtjlJSXPsmssVjwWr9nGnYcyGyLfVLdP7hFpqgewgNqDiq641HllScOMdMP
8FcuTOX9zP1/b/2w0B1e2TMpgqF7XVt/k8L38VMOFsbYqRzRzAOnFgYAxHRyhRTiQ9WR7657IEVj
hnRxiTYlNJbzmoaAImsjyN0PCiyjRNmDDDeqNRjY4s6aeN7r9fsY+xhk4kjDpXv7dFh6AxcdHh1G
BwXd4wL4CIp7kArt+L6y/LzMaG6P5chwwkVOrJqde7Y3lEeCAhlBRrtVRZ+Lqhp/2fgoOwTo4odB
+i3ij1IJmQZ4juZR6yf4oWijBmS1qka6BhRYa/PTYj6iz9ZqX47Jwg0EIpNkFLT6oSn5NzjQ0ivy
IvAtL+GMRY1LZ7sKhJYISfTVCwXfjdBynEQ0XRjUdaXW9xMxJ2ubvH9fJFLPGlRdy688HLIZ/KUQ
ZoETVXKh+28lX6BWGKmWMa4ZtkYWeqPpqeILVWKInxFfLDw9JcfhUbLDyQSi8MO7uDx0hFgZZAJ+
k3V9aSvuz+i5EltfKIl6zFLN+3wv75EAsuk3jexc2FQnn57c/+Ywx7Gz1USCmF3//pKvTNRY9XOl
tvNt+GiaHIjDS9Wedoc3phSjHjtOcWHlsHpP4a2thE4tofdyQgRFBFgPcuYExiM3mrqxYO9nT/lt
+FChFmG8csbDnity1nwwHiheUOlMZbkQ1y+K3L4AgR1e+mSaz3tLoK99A90IJUbLeZKDBXZjgvvq
zisEeu9OwY38A5pxrwv1Xg2o9hdgggl0DwXlgqZGDh0h273zD2XDjkjW7CNr5ADhwlF6tb6enLvk
t3Ji+Apktl6c2EDqje4kO+CAh3UWHdMTVaOUlcYGwQKZz77kUeiMjjB4r2xPCEJvyFkeZR+bTNI2
Fgq3gHbtKIolQyFN4tRFqixxTinY09dSbtBq9YDwGfv89azbcFaVIpBbcCeV0nQARp1/Pj8JPZFB
OHt6Ke5PFdNuTCfKWPX2Ae7nTaa9m8wHA52Be9v2nKp9RyaqUIBVN5NvkGcEcfLTSFfy4yyg4oZf
WSH1/Yh9Q0g8hXYwqktg41MCdb57zBQq3K0VdEiBW07r+9eWVDMo/eASbV0JwSPsAABhx9nqX7FH
SrLwJXXLwcJe3HzOGXVnVhcHCntTs1TyPdUKFlmoIIdDMbo5J7SlDlewv6vdkOIEpmK+oTTtxICU
OuaycLFaNCF74YWXlmg+BGuv9nNh1BwwuHU1r/zBYgxfwJPeUx4FOPtoROFK2FGqdSeDe19Xf+rf
oeB+vJPgTwMYsmmXbS5rFDBQnQv+37Z57EjIz9HXSKnN5tnznGkBW9dvRXlz9mRFmVebjx92Gm8J
GR/s8TgP5rTkchV33LBauomMi2PtDcgfD0fZB5q6DR7OADAXryp6R1oByUDqfVQJ5Z6vTvxCn1YN
7Rtq+93/4SbGJ8K/yjoVTD0rImZoncjLX2Gyyv8zpyH0mPJPHrucR9Pk+szPWWsUMTvpl836PYe+
5FSDyWHLkhWwq17Qb6r42anrvbg3wOilO1jlcRRQZDTpqMjQ+M5jLZ1nBf3RGvWaifPE6gcjbIyr
r3OZAEJ0W+uzhYJQw9+BMmGIneE2VsAr1F1kqqnt2px3GloRL9PzATzEFN3Q9QpL/dWPppuUeFgK
Mkjjy1bqUUqNqI6uhWoTIMQIFBe1p6xVFnD8hKpdZgABSEQI3YGMXig90N/olPfRCcq4AD0xs8WQ
NTMqHgXbcZy9zW0ZExOD91dnRQ5t27jH9POr1/6Dt/ZZ2tSZd3zTGCs/loSGYAyOBYJs5P/mRbV0
xhzXlAXk5xgJP+EsK9z/+Gyuvp/4HVPUQGBxlk1jYfpi47HbjsVherOd2wyud4cTzX6ey9j7x1QP
L3XLVxuVOTIokb0xDccCDW6Be+ieeuf222vMUMmSvhA1hgdeNgwLVZ22Bq0f80qkvkWVWWu7ic0t
2AB4oy9pnhfNbSHOBtU/fPdFCHJSUAkUjs9DP9ZJNdCE6fN+ExGjmIYURNyqdP3lSGr9V8v+GAd8
XvyCtMK1GRJpzzda44/D/GqFFMDDHyAXex17Zq7h6OAymUuZhBp4XrKaCItMqX1rCbGtqEGueF/l
scNbOTYhwL2ev3/pRK63eqfT/zA2UhQSKv5yKW0O+rw7UDg+Hpvgyd1xmOexgLmrW2IDHalKbGOf
aTAbE9n1T1epufTaC0FpSoAwcQopQzTr7awQ09eoB5JihLSHIQ5Xdl00LqeTfZZKuDaXo7RFml+H
rtTmGmsF5/2HB4WTMM2Lphnbfq0lt13W2BlRyPIVR2SDKeZQNC43+pDVodiii0lOMUXQ+KGrW4X2
Zpqth8UsvipahyxO+vaPkjq8De/kgNqxmmX4SAqOJ51vR74PrRHz2QqeLe+54wSrKY5HQR1bPdFb
EkwSMwHFlWRt7/6y7KHRf6WURfLMmA8Er2tTQYcjN86bnv8RjaHvCsnLhI0C6VMsr72kui7jGX0O
5PSGNkUA7aYFHGxq8F8shmQ0C42h6aceSPYnpYkZBwn64xzj6ewT4wHCD/FpnMeyZPLR3ViGnMGX
xNSsu3qLEQzrPWt0O0GIgL1VlWTNlM905UrH/gBcna/dDVp1oPFNn6eRNTKRRBSTdSoi3kEw+cmN
20e1sedT29lMLTScyMS1SP1SRgoNuZaVU+7wBHDHXKrvnXM35CwHl7WHbuWHdLf8m69bQgkgpRqQ
UJP/TAoshiOvPPs9khzdXxKVlu36BgO78/p3E0oUuZstvOgkyKflQAw46baIxHJjX3epGgFAICrG
8K4v8cUK1RD11tguKopdVQevPRMexYdGoGhnOJqeiXfPH+t3/iyBiyOnLGvDmxUvGtD0snF5jGic
JmdwYUlGMaG75U2EJI3Ydhge2WssE5+5N80lkT4yY4j5QvcX6o/sMq5Tg6cw2Yf17PH+wrFmAzj/
p8sYdzIq43yAfkbOV8Ftnxov+uo2JcOpIG94pPR4WhdIiORY27R6+9ODRJFxiVtYPCTU+2dBTdxb
P19zGT47yjvp5vwHDvukgotFtVkQLiRbY0ByWN3q9/bjFZCx0RfKFJ5RmMY37SpyXt+StijA02XT
bJeM3JIXQEBN6mAehcjJW5cTFsqzsEJo7D+4kJ1UT9D9m7hquaEglquNQM0SzAm/Gh6WtlAyPAtA
5wwykEukQbDvhGTjv1ddcMmMJzaWI+bAQfwOfebDis4LKYkpIhttztbKTj9sRcO8ctK/onR2+dw2
zbMEB+16Xr+ATHoRiG0ARymMpktJLgTYHStI1PTKkeY3VsEwoZf+9WXZCWuM8YZ7cUCbyLXi3cou
Xxy+jEJ6dBO5jA/eXxDu/BHh2VFRvkt79IFPvVeNzCmByWeupIXGDV9tTJF96FvL4Esi9uDcUMPC
X9x2AJzqMlzJ1Shcgsf2sxL6SAHA8mn8HjBeeFMj+9fipAMeifcShWJUsBZ1MmVKxnNlMt2gpBU5
kyApbJcknrxJbbE9ir/s7QUhrksEhDTYyyGJTjLxb+22wqYm43xzP3g7VXY4JR119AA2QrCtScr9
YLSo7yx6ABLQDFAb3PFiL4qz2PX+MTK7TLYDvAxv0ulTMXJbKHuHuaRLCNqWRpA25wobL4PFCktT
dpy/Jj+pwe7iSwkPeiMrKFJ1TenBUqLznpNtrWiefq0915iu+CGzpfqjw9BGvcr8zdb1sB7K1Mnl
lxADf6hjhqZug0siOaeJ9rDD7dBLwMSrJaX/TOvdwvuiNNDh79drgarvgBPQuP3oKA038sXXClJZ
fULTknl7sUYm9fyNTWY4pErWdWWRU9yvYY6mz+2Itluscr6/snRnE2a53WBvHdIy+i1+12uLbX7I
f8HNg6h1qF9l4lmglneECk6esOD+Lc/doiqOWlGXWpjtWqsjPrHLC14dtP0yBjF3li/aEAUgBV0y
hIJno/eDFkbFV1zFqIjVEqmfg7YQz65qBCQpW1nNDHy0fjCKBRWQKiWrsTAI3kGQ94XRsldUjboz
SmnS4Ub3/VUP7ocULNBplHZUgaQEuXI3qAt56TFqU+Iz67WozUu66+lzfaO3sTMIzZXoshZBPKGm
tOlxhOt+HVNdotJOv4I/45Qo+jIM9h236hjsVRVqOuVK8mB068VF8W5TQ2Ql43oBmuwwF7/ZA+Yf
gFbHMww4FTX6SBulpfyGtmHxJuxj2Q6hZX5VdkcUjS8XzD5fuKrlHDk6mlf4tyaBWimeoNhCnK/z
tz1HxndbhSQfcsCfI1uLyEJHX18cPfw7q9W1q/mPQQEKDbL3J5Iuowx7uxuvGtb/TVJ04zRYSsSo
PCDM5u0ARA0iVtnd3lTVsouZ5HZy5xmEe92dY66LwnP4ZKovwEp2NJq37HFXcUM5IfnrL/ZrUD46
tBAhv0owOQBSiKZEDyOLPCO1/lmblX+5f77AobTbTJXwNgg+WvGJBohHcGS3lB/ZpRDaQjMc/S9b
J70DRg1tD9mCbajsckCitZDuc9H1Ht7bJDLMx5rCKvljTuBXN4tOiISL0SiD2PDvMCYtxH1/Dy2x
0B/nOoZqRMtIKdEV+w1jk9l9V/CTVSdXt3jKpP1Z95g1T0uV7balPGV2EK+vzC0MPcZZ0RJH+2WK
JKHCDObMmcOSe3FvbujD1fPayUVMBDh5GZIpCBu91PHDDLU7u1aACV2riqCguk/00akh1+B+JBjv
N3NklWj76QwKuWIsI9mreiOKTXCuGdHUEAj2wmezTfqnrKyZlMKERlbdCt/AkGi4CwkVp6WgjF5y
llXrSvSEL/46A1f9RgDOponxyDXrG0cwWjsFezAR13OhOMuN7ltFs01yqtMBayuD8Edp9tDD/g3b
Gxs+n48gSlpIXbhDMuXrk6iPF9JO4Tee9alzM9oWKp1UlFd13sBvYeCdWgEi+MuLtU2/HbSKfd8l
htwbUTS3rUs5sTl9Fos8X+pBdc1f18saAV//v1U7gL1eJFNTusBk19wj5aEFQZsEnHDuMTAEf+u1
IaLUQwSBwFzFUMDZTtRcfVZvEtJtw0ASoDyz191TV1KPOhKmvOfb6awOuSfeFJSC0m58xT01iPf2
dxDbbGbKZAk1p0OOYHTyEEOydgIsQ9KEQDRMpmfmcX2BseVMEOzLN/ZVzH8UY84SUFkdF+8QH6VM
RAhr+SYwPW9K0L4NPZtY9OGJxfxVoclAMxhHycW3Xz4NfmwD1s3ojBBOPxp+swUtjN/2EmYNp+zY
YvtWgQRrAAUG03MTtqqhImnngRLcJAVc93AEtSIWmYILeYkaeV6l7pQrpo69ANo91UZdmyCBtqvK
JQ+RTucosDpUh5Bvf7tJ1DHHvqur9TDoc7xh2QUEFddUCdQzUvNtx+8GYD9rK6uHcyCnwTlmBZbg
7YAk0lG6d3yITxG48/ZhGD66SaZWu+qupif6RgQdIJjMZ+PXrCht9lSWIMUchcFJvjnqQtNYbLbZ
JvCvpd67JW7mBUwOXZplX7RnmjMnn1JhKdFMhZTGEmPaKQKuZI7gEoI9ju8O2b/rdsyyEEDQnbYQ
uveQRiXJpoYXR1EJcY6lvpdQMi4cn5GagtYmoJIK5U99SZHoHvf61KFleNUF58gpR+eEKDKflNOQ
Hd7xDYz5abm7bXHzzf6ftg7it5UjtLrXTaGuSvGc/vEl4erEx4nL5aOn32wKRJAb6loPg93m1DXE
LcL0ggaHKj7dAHFo2caojbcmdR+3kUFCf02ytqtzoUe9yeVPgHVXxnXwnsydObyD9ptfRKfKgZJt
ieHtMFrqM5SS2Wd4RldQJk/7OvsW/neSAZk9DLzKXOYcyUnlDDccP9gOX3GNlufgdPmvhBOt5/Gq
m+Iy+w7xXW49HRRlNlgDp83fPPdoW/O+iY9VIzY+j4KhR/3C//BuATkmtY7cu9kZLYZZldpdpccT
448W177x69hBk2WWacXWLLieVXp4L9ZyxnfXItOjIPsgXxLCPys3mHKKNY2rAJu3oC4RnES5GGjl
T+9P54EPUpqDadBbaxB3ShL8jRza6Lk3hDWG6BzVuVMwr8Wqj483HmmALTbeS9341+d+veDVGxsU
rxisaCE6C34RqLSChG5/MLROmvy+tX3LyfKrw4l4xXwSbdv1KrPP5C/YLMrq+xDcZG7S7Ad/hoEo
QLlC29mWdS1lgN1rWRUaxhbEj+g5R36S8At2NAODxhrmpClz2OM/59yjcQG2swkctg/MglYs0uvP
P6Tn6Cl4kdconF3K6hCGnk+F9OD1BzSAmnULNaFMbt+gAHxIL0SCcEzx0/8egwTq18knP8Ihd3yG
7HKBItqpj56CuGMxGSJApcn6Hq3Sr4qZabPu2ScM78W/cDzf7iQ3g1rzrSzYRUZgx0ElxgA3pxNb
VXSbQrIEF84ucg+kbD+ZOdz54MiVctTCw1naQdt8YNLUQiyKKxDE9+tYbvuwje8szQ3q+GS5831C
D9954MOZnnFCupXtjqndlWM+TgXlv19Ws/fmzoM+bZvNgFnUlnUPVQRUozxkGM80U+ApxI+/udh4
+2KoeH4Zb/AYj1P/PS0Uskoxdv7QW2Zwpx0r0Ei1A2yUxXdDPEnOAldOFKncy7dmbAsa0lrQnzSp
4m91Z/UGK0exjhPOuL9G0fI1rMImLjLEP07PrAohVwwZuN9E0uZ9LH6UhF3YDGshYwRA0wnO/xAA
It53O3uM9JS5jz1BJiKln1YrbLz2IkeGQsHTFLWx3bDW16654trAhOPNhlV0XDDRkq1cIGj6lniZ
0zcoT2zTlOpjohKvB3z/twTFoQAZEB6u3rTmlL1vVxaruiOgK4EZYWVnfxQN1nxxKzi+rkRi1LlY
QazZAe6W0Rs2Fy2/Cv548BjSTD5KnECbdrdX09oWhZtHVY3+P471oROh2tvp3Ts250wUzg3R4XCt
10yyzoUgi4GL5BFYCjOmV7U+khW9i/63S66/XvZdvINzo0eMzJPLiKsNXaT+tRTUpsSGo9i1Mb9H
kYkRQYoRXJM+FPxPR3v3zS/MMnwtvCcjEoakR/tz7HrPzpV7vflk/TPqG2yVG3FN3507hqPttjYO
SEjQLS0vyZuaVWkITNb8JlHPtqIpCe78MzfP7/v//fU1to7xSVKI5TH1AIdJy8QqR+m3nKe6zgXP
dzEY2poKt6xBrRAWcOcNUOtc8HsTslvoOdief6COusfITjUt9ylV6KfqiPVBtrts07yTBd79445U
tkfhDIQj2n1CvPRqFULwbNZat7OkNuiA2zoz8us+HlL8xI/ncCvR+gnvTj6xfTZB3IFYQuEMl7yW
NCjGlYBaOpOY6tFEmWf2Sv9BsQwK7gSDbnDY36mK93CpdZtw7+BbSRJuKoe/kfe24njC37D8c9FI
+KbHkbr5ly7rXOUpER/w/UWSQF2fIdVGzPVh/NFkia3UVz6NZutXFZ0Kn3tqXnAkbVHsFhgySjpQ
m0c+7xW99xUxav3aK/6yxbmVZLPcpQF+cKfrIsv4W0BmUsxLcfxGl9A5EaSg9eQiWm8rGIg4E6LF
eSeOH8DX/diivXOcaWCDC+Tt9B5DGJSwK2Ea+/Jv0kpmeyUyY4zJb2dWd3ADMFGced7P1NoUdcou
WgJn8Pa1pJ2bnIwYl8OaApnwZKWc0QWeFcGwei/huAXWDhHI70trGjPVRtxoO7tITYbRDg4UvTtD
BTxZBKRJfoqrP5aCl1oIBeBS4SBDwLNdKoEctfl6xkdn+zJEqyKN48oHlglF9BUXUWBQ25f5z8og
mVeGKhT9OjnaAFfzBcfLztIRBqvafFt1VdsFHbIHupKWyWDiG0wcRivM/JJVnfrJCM6L1RgYCbRt
/JPQLlLhY2TUNbuQgJrGZWkS04SZtn6DSN792aXHoa0u26igPgmnE1iMHgyk+s9A5xCtYmVARSvY
iNJJzqpezBrJ2egcJeSy+FcwCVkAMAUyhiDSpku1Fm5VHtcI2WCcfclqZCSvosPqqkhWNaXcXGBC
KoYmhHwIRomU3AHTgMSwJHpTzV8JuBph4oE3zREQPl63u0lCtZxEOLD9cVaIjndqL041NSLRdYYM
PrQKBqCupMXgQX9o9wMpt9b+liKaiaQHzOvlqtL5WAwEkKibYBoHMfsOMCE0p0xrlTb++6yl2QSd
cp/4rkwVyKuCtmyy/Pc8dlKAl5JrcIFXWlyhIJJ52+EqrbTS9XH4AgQ+VccAvW/4yhaoC5Sj14CM
4syGATGm6+lr7KSwWbodD2a7wYpuQggFzwD+ZxLeAsD8n4s5A2vOtL1DR0Pta8iewwI2DfAFwGsZ
LEXClvUMNBWtrzyLmaguZcl5/73WYmbGf52dtsUEHf2+xkjhLHDdPPuxRgdkJZEXsV+lr1g4pD3g
E+rEwFlZVczR0GkpAHVJtyxPtFbKuc85psRn7jhvA0RlFRKaIREMmmMg9JIaF/Ls5cn24wvwgiSb
3ur6aJjp4JG0em6lGOGLQcobpQtaAB8oddX8zzUGLiJCp6EWBbFKkuiiV7qVhYpZeeGo2Xv/KmoP
F+ekL8mxwsggDyzUdVGS8dxraNE/cxbnARmwT26KXYnTLXRutv5koUtXLHu05HoYhpbCEPUuj4ii
YUKvekE6zNB6YoFDJesKG2zGd4UTPt6YuUbPlntKrbWvxR57RO0wHJXUuoeq5a+afNs/cu5qpjaL
AbtoL0co4hDMkvMRLWUiKvUpMgB9Y+F5J5h+ZbCWGDKq6II7VpxZkTnAd6QDK/FnigDQ/tT8BFze
lEpFzyXzesHzu2VZfABbjKcSBIIOP6YdilPuygLHcd4F4403TUvv9Cp6uYypGBTJaY5X4ZOxzxXy
gx6RvB5jG3KjQJIZjKTMSZfMfWDvxhhxlVAAzXgkz2inAJKYUz3D4UgNtGWegJgn35BFUZ7zmIY1
fRmnWIsfLs9fyq/6Ad6KEKGhguvCiA4oG7fEPknHOsf1jaW2BN+6FK+4nKDFn+NF50vzjGINHPAu
7maTGGg79+HNYpfVRKk8bCLmb40qJwtfwmZ4ik9yon3eeGvnnJ52qs8anFKqIz95tZFcthbwl5CD
tZtw4dekdxra387EkU8/bHAxdUPmdQSHRg2dzm2pWLJVbry/RicuEbep2FTgKLkRmKcuse2lzAQZ
GCcj34Q0Ck80F/LMED1BlZXLEE9+3G7fmkjgsV1aM8VynvZj0Oy7lUEwZMD22WYhlibwQXjOsNEe
z/PHsWj+5qXp1Tbm29yGCxmrAVxdSEqI6bESRKtS08cUhb9zHH8Cq/hBeNhxW5wHmoxG/JxmdIg+
I7mFyaia01OJbDQi3yvJ4xwlrMHg051lUvOoDoa7Iy/VstYmsoXHP7wvfUDLiUhOMdvU5vpvRGfm
MOxuwU8RRkGkM20eYH5LYY150nMJgB0CaCmIPCA7ueeX6oTaBh6UbuWHNjJXAQQywi8OyQY2d1mf
QDFBROiU4IGApARZqt2ll86fVjbbUR/fO60Lwdt4hHOb3Kxus9x924Q3oAxSTLqtrvW7HZ1SazcO
2+i4fFuiMueKLcOG40RCFbTsR6m7FTVTIawpBSG6xQud6H5RrEGBFsBzVtSA2VYxUCKhjwPz/ysl
dbsOLoAfxDdlkkjznnQDuKwNKwlqx9VTbiO9CZP9vRu353jWPNhPJ1dfuxk7yprP3m0M1dmJyKI7
qoEEAzKcByof+tDxssa++PHsFiCOFyEjB4UiR10eyBIPwejKt04IRZmAJCHVvosGHcSKguodxcgK
j2xdMwBzXBSPZ0zoDBe8KC1BQzivBZfe4BGTQkInwMgvb922DRXwvglrxVsMEYG7yYZQM/xRNEHM
M86yzH+e9+9FugtkJb5TMr7AmdFdH5iSPtxL6DsE80XgOiZq8AUvdcwKqiB9HSM02V63H/8zPzRW
2KPeixwQglELAsLVgN2myNmxNAqDWl3Y5hc1Q/gC8K9luXsCAwFSoVIYlVClhVIjn63Iw5WRqVDe
Cq0cpBaef+jMAPlOQo0sknFMaGTYljvpwjYQZ63p1KrypX1xrH0wQT8hsiOU+TTIqBzlwiQRWM6/
xl9Y6r22H66lEB9asqzwxGinDLoseaTmklPvdBtAnIXcD5BMF0kVu8Mw+5eHVVilK0Y5a2VNEwwj
YteXSBQdT8OxFzb2OUTxx8DVxMbbIvCr6WvQyKehKeKXooDAXzwDzA/5Yvm91xeBqpi+JWeg37vP
aSor0k6JKjzZMT0TamoVFNUGD9tImE8eJ0Px1v3YYELa2BcnozBQQpqG9ue7wHpV0lBdxC4CBJgi
aF5w2t3ze5zJyPptDDRsBpVcHilVsuK2THlxf5zeTfjTN4Ys4p3LLRIsdRGvo3v67UiDNmX55ThT
MniJVix/Chd83jbi6A202YZeBxh12ypS/uU3t5YGwIEfeWszzeaJQstAWKfGJCoFZkPvEeSG5+Gs
0xuKeuyxxWI/zVu9WeAlzIYlQuseL3OFbcO8gJqC+Hokx4Z26AIBb6pweTH9gmHRE5cne92B7rwY
V7ezq7FCP1gnDquOXaQFEDLT1zY2fXEfdGEB9VLBqqxDl/D89vOLZDoN0vmUH3ZTX94syzkZ7liK
GfQAy4z7iDk6F9XNgvz8oTmGVI15ASR5YCp/zqR2FQci3umyNDw5BEv5Ljtq/pyzhaRFHKIC18AY
JUcYwSokn6WcNgYgmTUVX3Uhyn+WPPmvw4DazMqgtB/4CH2lSv9vteySxE6hwEchAfdnLiNL6F7m
YTQYF/U7Ce5blCx9iC9jVit0p24Sdl7jWQ/So/ZIPoXhmbqZ+Y3HKzkyy2J8UDtST22rcpR2o4uw
2vQM3o0TFjvAQuRB6hlIVwt9RopgNIyCP8GytnOQLArAKPrZLNfdCM1kPrXnjjOQv5qw0dH5vIAO
R5u+eDgIz5kIL/fJ3vQjNsFjM3q5DL0zpN26TU9uVcThuTq8XhLIzEhjJXk4gty6ELcCHfyo1hpp
8N4ZSJezTpL0QOShQY6WnBL1DyKK+jCJaMdQhidi1Xk4ziWnuDdsACkWm/BzoW/NcULi8m5Rlvzq
0p7Rw4bonJK4AvdL0Gn9/yv2wjIiHZyX7sTfR7P/fyfl0LxEf4yzDIGZCdkbpn3mKiYBaJupooSu
i8VffqzieiEiqULWOEwaycUNoJAAua6NqiFG81CTYB/6dG/pycTCSMCG4DVWKdR3V9sLmjfrgAkp
i2aqiinfjlakU8bJ7woXX/YXravfM9yxL68lOShlAwFAMhLX/kMm4CeHk0Avk2lRwMvr+Q1O8fsv
X6tj83AZApWjHuZdiCMmwNCIobci3eXvVL0A5QGK8qWwnr2oNTDYM70NucknBt6vV28B2gedspUw
i+RBguwxfGBXbpLLpvtmQwtxa3wOhAPrzQnMUyIllqTj3ui6VuNlKxW2a4yOmoO/TihXyoUB54ip
z9CUpx2/Qg7soQyBzB3bWWCIpsMl2Qq3Ay+OsOEWnaRR8v5ehbYuxcJBhlaTV11UBMyQhN5fBBp8
EsBFSvWPfmkqWILhOs01WwgbUVMvhy/WcK65ERviHo4Wgc8yN/cwyZ5tr6lEdqevcAr+OgKJ23BV
vtlVI5nQkX74+p7HuALR22TS4N8ci5UJeuIR1J2mL5I7k8vJJUShovqaATGdmDP2UlmxU4Nbllaq
6SPYkCH2wMG0WHXGWtzKNvkQWYt0ZWFJWJWa83FFI/BgvEkh4IG05QL0wfKQE70OIYcKBfOxg9sP
aog1+VSTo7ZKUmcMb0PBZkW5d0jhnY+v29z5IElrrsmtbyUdi/e/GnLN1e1EuWseoc4fRvMm/bfK
DsPxKExpAfFKLxhdkv35HqsPYhZjkG8aC4UF5uCFtjh381GWbxatzxFS2feCVScUnXb8dZi7mPnY
M3YKO8kclg9Rd2KluiWLNFhQ0/cpEAhYSqtzDOD1zqFSfnPai3FXc7kvfdcHfUUeMdjXLSVsXyQ+
HhIeWtJE18Nr0VmGhQPZMfPVc0GDO9JaghpPERgKLAwPgkpYJZF8YGG84pz+VVt7MdR7CUwwpnuN
tQWQlc3f2otIe9rxfz/o6IkMjsy6YTV40sXJ1glw5KjjKYBe0UKCIlJwBPpCZLVp84Vr0rjc2RwC
wgFovqt/PXncaS/g9MA/Yl9PoB570DukGhqxSyNvZ9dz7vPQUNxi3smB6JCeUpYlij9prEaIbbBB
MfvWAXxjKGg+ihLjLymZebzF2aGk99qyOXiH4ePdF1hGrABa/SjyGlxnL2hU9cREH2dF1h8bx8/Q
O9+r/OWAgA2xtt/CuOIbMNUVChUi+6ycSw2cfcVdn6p4MF1NIkFa+tY84rPvaPdbqVKy2j1HPoje
0vOWlGn09AfZcWadrQd1a8OOjBiA43qrShtKP77Ln8qUzd239onlBRs12CWVIr/yPC2stl4NbjAa
BGT3pTuva0fofsA3u4BNsDUzDIYp1t6rD/LCXrcq3NS5byk2fr/CY2StlH4KOiZDc7DUWRxZTw85
4+YQ0xEVWSkcQjivcidBzaFMe95aDRZFAD6Rcd8pfnTSbI2JQ9xmOmicZmuVguy6rR8q7bJn9tuz
PU4z/4wB2kezVu+a3OKWsH9TLxVTsucXUDiH1CL6WlhK4ju3yyoQiV6pQae40PE3EgKy2fK7YgVS
BXMucy+Cgfcv8kXBBrP8Vh+Tlpk9SY2gXECItPaZMQug+ezSzQ7NFcQIXxbP4kszxNtDeM29HVEU
vq5D40j3iG9J0uFxlZzRBc8eyvto2gg9Bm8+w1s2o1C0EZOqjPJKQgJtEFKlwj+CZfX5YNwha0ZJ
MDro8KBhvP18EzKXviMpCnrpuRLQTU2nzjZXpOxxzE763IDkkGNEIewF/OAdF3QqIuQm7ZlLVHFt
a82jORC6oQQQIHtArqIaqjVSoxVRSZBMlL6e9eNilVPnoXwpKoGvusg9uyh+ykNeqyrzT30GDhsh
73avDBgZ85V160hXtjpmr9YO5s+8cFP10EySpKjSNljhlUNCxrAvMKe7xeLNL/UuNf5x6NxEQP84
ik9j86xCDCDWgxpWwbEZNr/hHBZ+OGAoaia1QqQAQs97bGfoqn8Z59v7j9RE7GKyK75ttQ+ODvMv
FP5GkTqm+e7M/SD0MY8UfRMVO/iV/ml3UO7Li5ePXhyiYLZWrcB/8QI+2Eo1evgQCiktEKcvEH26
rEI21mDwhJqfSg+xw9Cq+97Ht0N5qNs6zQngKWVNtN8XxtmZggSwT0im5Pz+9rD0KQwbeZVtXw/x
iZx+MfpXUg1TBHGceV3kSbDjfMyFllT7jepn3T/BO+IUW+m6b4IdjKB4htUS6yD1pgReF0t4Fs3U
M2FPC5zTtlT5ZJfMN67aB5bx2+R44RAyy+LJdqzgjSGqA3WVJCijIFXp+bkUtsEEBnInbPEBG1B4
yYybKv7bo68PpEq+ZyQWW/XOUIqUa+h/3cqmoqjWnrYXUNUf8wmPMSoc1tTKs5Bu364DJltDSaON
S8efK34okEtgyDQNWWiSLt7eHBIC3KFK31zn16jfqkQyt0xtyznXa5+5Ey95z/rHeVkHcaGp6jO6
weLXYnOMamld87wJYlsR0/kljnK+n6Yj9CgrL16YEQ/L/FkX1NEJSXHeFNW6wK+FDND0iCshwiAc
os763hs7QjZcO/OaT1i6uWdK/yf4oIcCJIDSAvNSEmAZo2C1YtIgRp7vWj1po+ypG7oi99H1wKbQ
zv89T/0Qd3+kApwoyGSYG8e0qUKmzYRAoyanTNE93ifAHg50LMDVQ85nFcTp5oodfDqNJh0ywfId
kwEcGpU6nnMBoGFvjMz8UULbOFH/PzyN5VPA2xjqOTNpRwYSfO6hkxahvNjbAJQH3b67ra1d2lbG
B7haw2RUoxXeIJ6/qsCz+Fx7gJ3QOvKAoW5ghkwu5v5hcWnSrq1oB58z9kqdO958YnmovE362DXr
xHwXqqH1Qxa5+/4XVyc7ZPUzRxpmoJs1ZzyHc+vcckdtXJQksLlsmDvZLi7HreZaOX6Vv3yPA/Na
3oG4b/T6QeEGhKKedsSIgA1vubYLNexOPV1bXOj5d4FucDFxJncMJI+DPvnsZTH8nKv0uhsdNy17
bGKxjlT2cpwYTGQMklPAtbSX0mQMNxG/HDdx/Q/y7ahP25a5x4EdhnGsM5eAtdVRJqtjV3TAck/j
jr3bPPOTnLHfFCug86t1AtU7brgvb+RciAOX/LKdra+w0Y0KD2/soYNO1SDnwzyUfb8sGwID01Y4
00SP/7EbtqF96zEf8NrqdsSE7lVS9gxSBpUWDJS9d4mXcvfgEj6n88r0FS23xrhk2EqEENB8CsY1
mOKAUg5oL/I/UKC8RlhEba/xDoEXdwuXxwZcoWwAiFaYfAG/+pBKzF+KqWbPptFUbFEvAJEButVG
gHaME3I3oTheT7IpqI4w0PFfKHWHXcaRcDuztuCgx0kxpOcJbDm4a4ssZoYlk8xXNo/oJJBOViXX
+vY/iGqz0B1sLbIYkRdOMVKq6bs3bM8vZ7nftDk8bcuXN1jf8bXysPBrzv/lgZYBtVnYqq9YImRb
JQgnrCRZakzV0mvTXFXGYPvQ9fH8ILqCJMEiG+MX/RZO7lheXJQF6X7nUS9joGtF+zh9ROVlEDDq
C+tRx9oxCXwW/T/2iwqVNu/6kVIvi2/wREqvN/J/kiszQ8JTHHYdZoX9cWFnGJfQZz/SBOvHppu9
2uz3Q0XzyqmOJlGEP1xL7ojYcmXJSiRo94e8og8cWeo00FrOB3KrxHU1gj94q+DKuR2a6L+leJHW
CnOPJFnFxpfVmioAkTaz6KJvbu9V1uY5Jd2Gl5mabhSp3HtCLXpHPpXzbVkLv9eaRZX22ox7HeWI
UekNFnXoBV10UF3Zare1f59Ca0xv1qCEL1o+/asfLjvhhqILbzi3+1eVaq3/DWr53vyMoLIKmPhY
THuIXQCR8998QdglQqS2IcIeGoojzTM2bIqT+r1N4B79xvoAv+4uV1jbE74EXdoe0Z/lTONEKQaS
JQ2HkgVEJ9C0IFGvg8UjHmxrvIGFbmovK56ItuciddaoMOLYvTROGB+duK+7RpuHgHDwQuPJ9sfr
2yuzOaK0AZif5hVOs7ViibKeHTv03XA5mXbcCQgQZ0JZy6fJJhXXOX8TYaQALToPX8Vl4gzi/Qh8
twOZDIFGeioGXpfVtiz9GIQRbjWOo3l/cZqUZnFp7hwZRFrHFaSDFH3Y530uXtjpsBh+q0Q92Em1
sckHZwGl4zW0iUZfMYvCXOn/oxYDC10BP4tHHITQBcF8gw3Q7JbXYkYv9IXoWyNXeeLko2cxm7P9
xFfH9o5tRCpDY3WedCbQA+LHe5Ci05oiCVl8wJeKg/1Rpyuz1zzBucaBtG92NeDKU1kwBFTse8iM
0wBxnWhJeFSa8jKI9HbrzD2zuoYt4q0+nNYxRxlOH8uubV5GSiBpRxJs7gTYt86wgwVD/OHKrirp
OV3VrF9XoQeFYs6hFz41ZvPs566JKID2nFwjIW1VkBSkETtC+kr8+f4GLABJDDNO57R1CMJ3O4V0
Gh0pQAJ4P+M95pUA7XDoL28+U8y3GfozREcaQxZG/G4SOfe7404SPPt0k046sGk5dabrBvhvRA1A
RoCdF6vBLYhijLtpcIY0lh2ja8PtFNmcaqODvEAVn1/98Be0/8Im0H1Ms4CbhFACAUDKyjQ0eqOp
UGbDv2eMSbxuE96McUySAy5FeGpqqScXzeVBvahEMVmW/ninjVam9HmN/bZhVQZWKJoQlZh6Uo+v
gb0oxNyDV2uF0waFLkjKmgMyhBP/zpVAs8BT41oU2IxhCqQYIzIgcz1Y+IXetqxUCZ5WOWDoxUnp
GqR9iwO5UQm3iOsqvpVEEHZN1Jedd7/khgYASWW5RQmmQeY0/RfpQTnoJsdzH4dE2DsL8BdLrTKW
zvfRR7xMvVXwar44v0PfGk8u9nW6lvoMLMF6fAtBgQa2xQPdp73wroQPwU2G3MY1OYjjS8DLtz+b
sNSKgvnA8HT85JtfVqz50B/auinW5Bojav5Uisf/YiJfd2UHVDOzPyy/QFLy54/VqDOd8+MTCa8E
VnmuDYESL+GaftuOLKmrqxbM8Da+wyInvRuNE/xIpmtzyzqdU0wHq8ExXYY5fGrYvttDM7PjQ90w
khJP/+ZzqlxJSAewTU8SOeeU+xA68y+boXYr3YJTmikt5KhA9sbXtoBiS839nsR1lGalwyTjsWWK
7TaEJLwr1oB30um4RErm+VzZ396ShNzsfB9zSzXFYwsKLvd+3tnkASpR0SdUeUlYsUyZs71OcBeB
MeCU1u5YEhk+DxVgAcG+HuVYWFcriA4ne2GfG3HEitpuZkxSqpxMNUnMk9g8eTjGbDPjhPsy8BgH
3CTrQFtIAOp6f++WP1mv5vNTGsTH7NAIa6wI8UOFKrNKF+Cfvxk2XyrhF8wpGEjBOdXEA/kadTfz
5KUQTH/gaESEondBKlJseQQ5ih/V6T6DFKc97wE6AR574UNNvzM+t+b5QYXBopwtw+nKzIBWEetb
p9+42GuoyyGlq4waw7bPD7Unp1ADh9uRRpfxhxFUDHcwfHpAJCifnPNN6mOK7KgrtHNGH+QNjvrF
ao6LoTHXZCAu5mPTYocri5RXG/JGsdioPE3iiiA84b5+s016R4sM0BmU8zMa1PimIwEYsog+7wiF
C0hTkS6q2WMXt1y1ZgTGxlvoKBkfkPrSbcdMPMlYtnxlrQnB7pzlowoR7mGOHWt4+c7B3LbcNEs0
tFHJ5Wtge8arx5BTvVZqrSvvOW69GbCylsuPa/6R/mjk0dAdqKOEnPfnhAx67zFnXt2Pne3oibE8
89BpeRWKNy50slWrQqjH/LHvXsbFjpM8RSEYtW2tyZ4kaKEJaR/qr2077kSx86dvTVEVzrxCBZdo
qCuAlvRkh5BZlsKGomR9G656+hYUzm64Yq5jeuA3xrsDbrxfA/w2GONB4RtH9U6DClv2xRvk0o5f
p7n8zi1I6ieZ4M1qucGq3hkGDhe/MLv5hI+tlxWzSyZwh3RJSkOYvnyh6JAVvAtU11flONr4PTqw
UAROXlsYh9AMdbwmLbeI3yG5q1XTiK9JwWcmS1/Be4e3nj7pyTsAAQjMhIrllBPvZvknPxBZ87MR
mgP+xrZ+qQ8Ojwg5eH0aYfNQMbq5iOuIwsWtxgXPxu9zH5lJv2irI7L1CNjCVIGEEK7EjsGrc+zB
a5CC5t0EuKkwGnMsKhgiBdESsLq8gqF3XnRSQ9qZ9v51KWYyHeYXnv/IftEYgkBKl7o1xlQIRlSs
7QwZ1zXpfbBtjtFX/klVdYuJETnSidK9VKHOX9oBqwu9B0pu9KTt6SVdo8VDGrwUfTJcJfiH3Kpq
C5WKxkkNS3Y2ljJ565RM0FUvHTWrz2Nm5M6dD1fy0Z18whFFr3BRUOi7ru/ExllHsVIHEvMqoYsM
ULcaSb6MtrcB83lz0+/ruH6AMnIHsBtHFmTkGk6QdJTZ7QLG408dX7Q2TjC/9qRriWWcp0ijhph1
xc8JlnFyaJFkxXlaekknLv79t6CC8AgyJLw3fYXW/Khs+Yn7MjIWS+tUVMbXwnIo1IMZ7fwUrZoQ
hFqxvV8BdswALbFmnqrXKaneIuM5K2NI1WmgEuzmIozFzqaonDCrioHbH71iCdKkR8xTCnN1ywEk
jUt+891JSclYegpGBySbklMVN5jGf663i1CAeW5ILpeC/fsrJa1kMy/IuC4HFHJpZjoX1+Z0j7YC
LeSp41Rk+a5esv6Wq/rxG+dgbZ5i7HQ5Tf8UXOI2kqfO/4UY50Dma3L2n1iStNhkdD7nnJoc6vmI
frnPUsaFsGthlyniTpYDmZm07pAsl5zpfySij7mXLr4nc7UHDZaBSiq1yJYI/qG6pY1AIzwJ81fG
MNICfBydCkPszfGebD7Ua1xulWmW5b8Ta4mAAuhzLtFcb7Fo9lxuWtiaIiY6YkQZRJtURvb1Vgnn
Ti7xGR1fEsnS7QtAXtw0ApL0xW9rUp5iX4uqr9nG/bukaQUuhf74yRR9J+MH2fPlsJCSe2Ge9K2p
o8NBkVJN9uroxF26Cbw5Djdlv1qLAJ2GKwgn5JwZNV3HjdV+MLSszDgGfcS4KoFO8pJDSDm/3LmR
ih0rTRSbq5+L8QML2Mk8ylq28nyZpr7jgeF44j/dbNrYwZDbIlI2vCF1D9D4rRKB0J4B+NrNB9Sq
XPnU7HJi6tY+7QfNaxUpDpGgfuIzRobK9pwRb6qXjLQZleYU02Bb8q42pqNTQbrKyLT4uB/Hadqa
k4fnBfNhIIHsRU5zauEQtglQ4F0MSMCpGBE4ezKcqQEyDeHy5KfZwPE+pHwqyvS5Z84Zs9IjGoC1
5NuNarNQxb5c2DQMNsPrHftJyEO1bAk3tTjp/azGVtOqIjGIkzgUJmse8jQG+dzwIrYO+2vqbimP
e+/HqclssdiXm0HYJEMvdmTnoi6LKr6BqQlV64R6pXb3lllg6gXUXqzOkvXsT8g2kQDK30DlOPDX
qF+oHxRnR/SeZv/OVZXLoA1kUn0wpSJtDEmnV5i14EcNxt+ZjfwAxwdV6dSmGDtH0DZ19G93SUCK
7gwaO0XCJT96gjTFvyu1Qrg7GBHX/xO9dgxMrl4iw8iswnMc3uafSPTzaN/UdQk6lL+P1g/dRBPa
+eDCo6mmwb6HqVKxvUI7v0r0T3NGbr+vpC9zhqTJ3drzWL+L2iviGlxoSh2H7yHLEecF28AT+OgQ
sAg51Wo/RO1GvAJOk3flzPRVSoTILwlYFEmx1Jm9dabByfaJG75ZYs1ZykAAuxk93Nz0J86E0uHp
jIJc3W/PbycS+XxjC2v5eDjU/WDWrpBJ2p7vd3Pds4SzKXsbfGcTBloXZ+zx+cFVo6XC2P0+jQzh
dkl009/aqURrnpDe31XS5ddzyPC8MATDQ6BX/YCun14JeezdcXYKR/5uTs5in7xRU+/b0FSVa6xA
gP6CKBIaRx10vG+sbVXSQWTNZbMPGMhimj8KZOPidM5EXsLoTvPBayCGTpKJpiPeMTj71hUZqYmm
aIKPO6b7TL+hu1L9aFYnWzoki96+3cU3L3VsuFLEacuM/q/beFijQVUQW87B7cUx+IuVl3OnS5W+
s+iOYTLGHXsqdNVrjeYh1ZzRbUCneE499FW+fd6PfJebi16nyuDZnqzsDOV4sc+oYSnfzPNS0SZc
v3DJxXoMvO/cd83aqbEhuDmflO6oqVjmbF+4U+OVpSDPynnCmzNVoJTHJGeDTB86OTCFiRqion2L
CcgqjOelocKBH3DM+axFNHamG8pKNK6eRdAUUlnnCFe79plcZWru2S2VpEbNlD/QzUgsBV45wzki
+V9XhWyqH//UNHRWQcjbng7Pis4W17RD6IAWOlwa9HL6KXna1J9W4PtialnDAyKgU+3MaQt7xqlv
JbcvMzKsxkyaQTo33/YabZoe/35MAPBgZmVPL/jdRyz9nJ4QPmfg3tGo1B0Obr+mHoceF0lmmjoh
hGsA340HN9UzGomDKsKKn1uyKzrVTjwAJn6SBWzFjEl5cgWmGIBRnUcMtAgy+5OxBwW/M3grWAXu
t6ETl3+fay48vwktgRtsWGEffSU9z1LA8qEByisAWS+a4h8+7L3gIfwDoKs3DjpsiEeHqgAOdWXf
cyFdOMefhVXippj+2o+wEOIWTD8y8MWDMjYWIwytqMHdEEj9MnvfIgok3NhLCRR4mfuhPTO28Jkh
KbF/Kay2GT8jwin7i/WnUNvaqQwHxYxocf57EozVFR0dvF18AILCt7xK7qglx7Clvi9XtCN5USX4
NgTrD8ixo69Xu17hyHMNziY0fah2D1969j3yipcZtYJab2VdLs7IruCcLa8lacArwGYCM0ZqiY83
kSllzq9wU5fYWD06ebY5Ioc8fd3753WBdjWupq2i1bsWNicdiPEOneqJ2je1p4a5DMaemb/no9CG
lundJ2H6JruhPmFclgnglLEPyA1dEyP9d+yykTdRd0nTnxTUyB0N+WKcN8ILXA+yflBzRO4TeUlX
tsxVCjRStOFWbebgvBMmzZCcS1AlSghvzfps6lY4kpXJIzSVcds1FgYMK9ewPuEGapoo0eY2KvJt
kcP5jsOmuSQZEFNMa6HVWqW/MJbYtbn9vxepJawn8llEG9osssKCYLRRA9FcHuZRoxYVuhv1RFig
OaFpM4jIytgUrOYVC/HNacMA1yWum9edVQNgNtOMJMd7tfF2xd1mLoIkrqcPzzRE3JgU1COOMzA7
jCr2NaQSWB8gsLTD/rlBkOYGy+/jcW49JdXixcT4moUp15Br1VHeWVoxhEpRezj2UkS6qSsnIFz7
slmRZbbLd2Qqaq7OJDzztTUYzsRwm1PpjyIl2fK+vApESX8w5IeIMamJqFWHswv6AyoxbUFA2Y+e
heNrvjKdlfHCuQOMAOHJSJWQFacL58DuJvmsXclfq+wDHcQOUtyTybYoue5KDkOzzPOJy2z8ngwF
ZnRBWAn82IPECdeg8PtK9h5Y/PFfw9neeUrRh91Wmmdb/4ouJ9bPMFoZO8ZK5Un8gL7cIUvaTbxs
XIaY0mECM9k8wU8/7muzPJuSLjK/4y2QupSTnLiwIDEPx5w2plNPKWZ+p9SGDwa5oSpzBUf43Bwa
4O50kury4zpVa021MHdia88NK1mKnOxGfQFspERn6iRnVqwJ0IpmJ8x1+JSKfAVcbxpvrjRl89qw
NSG7/AWKpkvHi/M/9bTv24mUGxfTg5eaDsJU3HIHeed5V+j9jAO+KZvx8NMXIJmE8hy6jeRmP48m
FYzX/tF0VKq/YFRgRYRPydgWYwp5vYGFbrUcA0O5zudrZC28GJb3zyaH1G/RyltrLKwDlhfEngvD
RGN2wn40LRYGwkm8VP1ANj4R6MiEbiya5YW287tkAldcnY6t7iBhDgRkyCYXw+rv9E0nqNGmTk9m
4QaoU/vEbarZJ/SxYbirhgV9aO0fDXZ44hyk8+EiovHY+pH4tQ3yHhnjhGwSeDodqrhWR9aHsBgj
PRzlaLblxDmf2QSunhy3srmuHwb5RIVF9mIgl5gTzblOgwGvNGN7uvZL2f+jNN5J+RCgpXOG+KML
yF480g1r1UCEBWrHZQYJAYNZv5lNY6Qge1i63R6NIFzDuKcEVKVjLPgPzptPACoNGuHBv9msrSVg
XrhlGrnfNupSbf0GM6ebE2DhblnYPBGcngMxpDsDRQN7CfqOsG4tslT8/8rDxe4Cmk0lF/Z8mLc9
zjmp3TdhPqa/XxkR19Hpi3pidlAYCeUn8NFx7KgX111RowdK/jvhBbrPCFPCUCv0QD1Loh7xFCP5
NaKUQyn9zMAJPqI+QmYNUfXxqLAGOTl/6OOZAZ93bdty9PRO9pZqduVfsB4d7shy7a/CFbbk0KmD
xeuVfUfYNvKG8uWFRxsjD2xBoEMHdHLvk7lYwM1sRZAFIJcTDRG7S3xWguLJGWtAmRaQ4dWi1F6a
5gs727bDVrjqW7E8xo+Yx22MWrnRZMicdlJA08NZhJs3M8J7u9Rh05amHaUrZrMnl009G9xBJMZg
bnieGUPoarrxymEMWzQ15cfa5Kd03t7b4G2gMkV5pX0ZD5TRL51Kyz7md90TVGTQWpOLTnBXldEA
d/GyVFbkseo+Eupz2zNX4Dmuq/iL6ZLwrky5iC/velpT6Yg6SFzleFDajemfsZ/b0mSkXaUaVOUJ
SUthipzASp/UG5FaUx52I/LMzW9NsUBTf3Z7ypS6O4qLjmNI/Lp1tQz862+OkBkwfsbsyOtmtq4M
NNUNuExCmj4OOg1kj+axQuUTDyIGqpscji1zjQ2cc8jiea1qzdnMg1shUMJ61wNyjxNHA4kKhUmY
RS6XFdUDilaWvq9ok7wIoqtjNs7jkAHajElZHylUftN4wgR8WPTQYNxXtfoHgQku7ik95upta1vE
fNlmD8GHdUmGRv1fKSzuMQx2mAJcivxDzq4vxrhAUcWexv6T9j+Uhd+OEd7g9f7M9T2j7/jFTyp5
YxR2ILc/USjQa+BqPGqIf9JGzsuxt1FXRf0Lph6WUTho2yKdU4GaDUfbkVqTks9emOTWCpkR5Z+l
J73zAPG8eqse3HcxOGKkTbZUBTl3q7Bs9jvwXLgmAVGyKLTfHzrlXhBtcN6hpdHRytZQGxy1AXWG
8yaAKwKdMlE3o29pvOAKc0d7pyq5Sv0HS1Gs4TT5YgeK2SulOBD/x/+9uMvEpOgFO8GCu2ZRIAKL
VBT3LRicyOoMCJkJbJ67w+SEf0ZRcrxl6D1uZ416gm9zF2TL6emoExI9uAkrRkiJRJvTs4Ggfjwx
yghHUiIGHu+qeSBkJH4TRavTN6mM41zSK7K3QBDyE4JnM8ovTbSJrx3rjq/kajqRlewM0otoc5Mi
dfgbWgTwKhLjGRSO7cs6XKwgZLELMZAgYmenWg6ocJITEix0ioan4/21+YansVONoPpNPhboPNdH
gaB783W9Rav7Ti+5SSv5va0tb9kSt4MH9wt43WSV04UINuDiFP4BzXyM24XKSZIKehC0Uokr0KtG
bIr+124lEfDPMGrVWMfSax25PKIC3z2QM4GiAt9CpsGEA1n2zgkgPwWnz5PWRnks5jOBwUx9AbZR
qcR7aa7bYmzqc87llepsBHagf/QEtY5n7m8L/RYHViz7dr9ORGmzQi5zoMo5Jn8eb7jtCdDLI1LI
LTswe0w4ER3L4WIl9+rsHStNH6vp4g1yyIB3NpTw0vVC+w+P7IHfemmAhKzJsgjDQbtTdU4q1S7Q
GJ4Oe+Hy/pYhfQAebPQCVZO1re5JVdSPJKla0b7u4ojR6K966q8CFORgwfC1exV2RsZXODxR6icU
qi7ytfl6nNXEVK9+nv259w50Z3QwWS8Utfq3CuUwEsTANP/fuq35Sbi6C52Te4uxsWb+jDOv/cUc
+l2dwM4UE79US5nmJjtvoqRN8KmsRIlPwbzbJVZrrQZQ6+QjdHAN2y3GKw3trJqm8gpolTZ5Po40
yDVvsy0/fo8yJA3aoLdIwOSfln4c/pCIU2acEjMTmRN8eax6+4CBzo39SYsqsD/i9a6/VGLK52hn
3uaXbbVRwHMbhHb0sZWOQBIOFomIE6OiNy6fJTMvkipgjl8FC3pBGYfYNE3IoA2CJburR0Xdyqcq
2/YB1YVHFS5KKzSDM9uzGLDGw0aFOq/DuinIh7t8m8m/dEfhkiw7xV2bRJnJj6p5iiWLTesdi7mm
dgT9Dz+HteI1wyn1fIGRUsqejvTM/ZwG5dLsFZeXNLHzBcRmLpHgT+dHSgdDIKOB1UkutykCJoqM
LiDam+E20Nr9NOb89D9mHVL8ztR1m+BStIeg85s+vm358lem87LhZqZe2iyh0UluwdzcoBhUaUwz
/lrojlj7m9tF5Ggh+Yemb7ecw03Dbi+MgbnFt9/wS6R4+cwYPnyh4dyn637ciwgrXTwTJtjfjMCB
9E84DSrLW9WKJkI19S5IWSbNBtIJdJNijgNkp531aXRLIsrZTY+vRSY9bG1DSxa81o6Q7dePT8YT
QKO71Y2pC46VG4zK9XfRe2e3gdh+Uifa8NzkOIl0w/b462hBuHzAq2SHc5x+Ru6a7q4gYn3GudlT
EZCuSHZsdFGW0ui+bEM2xCAR65kiLNePUoTatkmk8fqjQGvl3CmyIsbzPoPIK5GH7YxDLiN9dp2+
YBPakgU2wZbrCqB+2XHjHYmfw5nHzbrsRfC8nZH8aJg8sWMEFRz3tmwpyZsK8mO5mXkSmcSf7aKy
A54wk3u+sLR/NNpNwj6ClBV3eMA4XuCuvVQIE0/BGVCxPRmKH2sOCzpjMHVHvK0ltOQO8GjB3i3e
LsEL716oS475U+FlxD6kMqEs0mbTdxvCBDXGQ4+7zFDthnAixoQD9+QmN9Obpr6pNJkfo0IxoISn
lMtWeHKrLbQwq54ntBHwum1c83vBSmN3mjmOik1kw6llxMe54wmYN2STwxaNpr6sOLzIlohb8n+1
yuwOWTgdd4GHPjgm9EthqpDmMt5Z9cDTiPZGAOGHzSlLj4fi3lm8gS9hNkcAuIh5HH0QELyECtx8
Rn5FrLySbxXS8YKMWwVv+OXCVRQcIR7wrp0LMbHCOjGG6Ge62Ftknxdyh8il4xfbrhPXJ7BY2iuZ
uyHmuvss1cMO5xVC7aiDNFfKDZsAeZxb6hGPHW7bJtrqkzFOQWCX6rvRr3bz3ZIcWFF5jDRDQewS
pJp7DnzYK8WRpesTqehwTBG/xQj0vJpOWjKlBG9zC5kJzkBRafHg/VDkLB8rbIN93GTiVEsuS1al
UXUIo+TiTJGFYdc8FvMfLZJKgMgHOORHvokK9/z3ZMFEPxkkqa7g9zPiNAV67g6VhlEXGLwuPg0I
Iq9aUeQVoo+tLJenrSzZd3yXpUUkQcgKaL62+3lKSaShzVc43WpM9uBlUXHh2BvHmT5nK4dAVwQa
fLyBP9FWqbJJqpXrbCGDQFzKzYl2xl9HbYKwSZ7AceIsXaqG2NM6+MwqEelPkJ2+krB+k5omKT8N
qgejRaJQkVVP3IcHhG5hqdOkeD2EhJrLJnhNtz8a246Te7FbbJcc8yjMQlftyBWjQHqzDWCwfVJC
XR4B2bV5hbQbtA53uQ9oKFWE2H1UlOzt94HSU+fB4qGvZI55q5xWWGUI4DSevUAoV4o21gI8uY0f
Ns2YZrAtanvOsOXwlZ2JkeL+eRsS/dct2xCyfXt+Gens/lCZD/8YGuf2mOKlnxIZVbjiaUgw4h01
yA2/okumYb/lMIbjDuuLSRkJ9rq4S4D11HSbYHJURKL6Nft83Wi5OA/OoJfZOQZU9gKstwI8z9P+
IqCGnK6Fx99VRTCctdW+hTW5b78o0zgGut06n38zNPqnZzrh2ItCLUwRiKki6p+qkmqQ6ATARpll
b/7ofEZCGJaoMiZsIuoaMNMg+gso/NQDlsD/RoScx2BfQalrhMtGopZNV7xlw/8JYEbHNO7ZnxqQ
jhLkwaf4Akwi4q2DPFVO66J9bVJk1CUh2cgd+ZJyS+DPKshwnGUWyC3iF38PcvRKOoroclombQaz
ArO4TTpjiVTUHv+NBcWVUc27CIz5cPZh9mtDrLyVKqlIWOI0VRlWn5ySrhM94jBuzHO/Jd63w6/2
T5KiVW2sbvnFUcTZkIhTDaGi45kDApO/9Qk8nnMiwCjQeWHEUP6lk4y9+IErNXVbT2DCLo2XWJNA
jNFjhhBA77Eny8w1CUpD2nKKx1mFbfT4CTHsUq/k5b6D3Qq5lVU/Tt84glt0955xJGGnxRHqlMFi
kHEiAPetKTO76H+286dflayWozwOmYNtyutkh8Lw4NHjA/QiLcseq+163G67qLS2c4A670D7JOUz
4MCm6Db8WXwmwTiuLsHuOteHRU/Kkw1/4L0uHggaE0XSvJedHJQt2C0exMO7N6vfiDpNb4r+fD9t
7NeU9fiI47r6sIYfIx19rxWCLGDTkD9bU7P+ot2P+LKFpcQBttNf8Ag7hDmlwTxV9WTvEIWNw4Vm
dg2PYYTZhur0/k6pNlPTQwBAJaLUsE/2wYNSdoWI0GTp/Q83qcmBIhTbTdbGzacJVQQDSQ2pk9zr
tTWP2covjcswqj7GqMyo+Di5lROxhgJgsa6zY2HJJu6Eoyv9KOPeC8W7QDdlFat5cbMLNw2YEz7j
X5D/f7cw4NagfvdVEZr5lRfyjvGLW4A9Q3a5kHGKRTStN1J3KSp7Nn7vZrk1Tj2EEqdXJ2XI0FSt
Q87HKMHv0bqxzjs+cetXc38X0W1GmhskkFerxQd50hd28c0qJeT3/yxfD4YfJyaviYv996q570nS
lpPaDcadzmOQv476P0MtYiEiEDcYBdQ00OlBuHr3vLu2bNYkNSrDlzPyOUIrAKiEBhpFyck2FCbY
buh2Eoo3JxY3MO3dCgQcmcmmJPAw8l0B5lNurEdAMpI8hSclUFVJNZK8aGpniGL1ZtZ28AFDqJKD
ZGGc58tKn80wPY2ZwVg2tIJOBvqJJ8mrQQEQoE4MQaYQ5Gt6NKXuCNQNW/8UQVJ6tgrIEpWAZeOg
/Mpd2tYtcSKg0Jr6USoSax5QgZpfG6EdQbUk4S3ZsNxfHDuxURYIC9ZW9pNlVRtFhQEGajixGCPB
A0kcInm+jkyW1yA88wgfFWFO35zb4MEbCuHwxexrRaPPKzv+WwJTSQgKs84DsGn7Tj3cnM2cNz+n
eJPU8iKe6uHDPUpFPsFbHrfFmc3TI7w99eZ/c2yLwBMjIUeIGtbsyJNxT5+a30dFA4w/YvtaEnyF
uBM7xxIwyU2AbFjLwOfAs+YG/p5A2E4dazPI0oeiJl2tJFNDeEEVe6NT1sKx1ERaYfP1eqoGV+iS
znXVUy9b9t5J3AsMQfAfw0UaHSmalQY4WMW3znC7cU/crn6IVw+Y4pabILp0UMobHNUO/ehL1CqC
xM2AiWq6WgpoQCwUTOtM+Pwx6QxWs2lZjwmbiptslQ16ejNytaNXQYd6xQBw2nRKGZex4OPI9fjS
onSyKkg5vsdYoN5ZFj7i0tOlQk7tuSmr97jRhwj2svwQvAQEVMnkUzlkkh4lgsIhhJ7SDIk9aX3m
u7EOSrKmJeyCnE26dGanVad3/1qyvmnQEe23VCBDicQDcUR4SJAupM6poTVX9+ZSk5ab4s8Ohayp
MwOxOpznCTPzAMC6sxvu4CHQPoQKwcCRFjW6SaEKWckcJU7jqAiNFcJ4hoFo2Ib6M+xXit3hOqEC
W2P6HipeWbeeAWsmjhaVDxdeYf/Vh5nsHDezZgKujc+dcD9qs/BuhzfpmNqmOtQve2cJzhsopFdb
i0gbON3PKcw3ZtTtEEATnl7l1bPO/U9U99yk6fqh+0bQfejj5qy0bRabh/6zcjcyQXFNOMLGzNhy
HAQyXunBM5K1poEA2/Xc94PNId01rb330uNtiX5NlRZVOA9rIO2NJXPXR/O/hD4lUzJUGpJlBuY1
P8BFwFVG4gpKYq1bmyow8N0JUHoPP+zsxlABhXKKGaAASmeJ2evRHBvi37Is742uLirl3xkolStL
3d08i8IMLKSJuRa7Sh8iWKcF3rl1QfIRIV6coTJ1k1XSbm/PiHF8pAz74W53NYXoumpmfO+itcDy
rMJzI0Fuybr10cvZLCKM+JWmDgMg3TCAAvSd5lnM93aGmoy6z1C8KP2N2Y/csxiFEiKGWcXCPJLt
CtyzhtMTbiGbDKGwRCJIpxFvZYCau9737x/da5JlzqNhjT2NJ4lHWLMFQ9KOcAzHB0epsFB7pS0J
4O9BHRaMzn8ueMVokOAwVMF/NSeGleFv5H+QVQzLbvqncNmIhizUiSKz+yIUr7lk+TpZQfsxcDxr
7g0e17BnT2eZfvVxEJlIA0km3fs2J6/NJ5HzDRZooravjtZme0jek8DoUT/YKwg3aBjqcJ/CkvMF
vvtS4Ql2G8VKULWSHyCdGlUKXHBqqtGb7R3O+YYSG+81ANxWQLxmUmOf1fgI11PtODqNMAD1NzpE
lBDdyetap11sSKNZy14fjLBJBPQXVakbusjahTBsVsIZpna5Dz5gTegmnaX36+HJdbTOIRP2fzHB
40tOFktDPY/NOpnpQHfSh3sDSHhH7kwMuikNPS74Bg/DDF+c92bXYu+99Rsa+KzeLmCE9qWTzCFs
1F2bv5FOdlArO4ADr5Ybz8XQQHdcyGZ5SSKpQgvTbVtsEyZCCTvGx0f/3scMp9hDjRMz4qKF2rKr
ZDXgzH1i4lQw6sw7N3bABdClINYX6o6IWbgv+0szfjOn+j2TjNgpSOdfMrN2C6ib+zHVcFEts1ZY
4Q75tFkQ+1qSBlX8FkpZ4zp75uC7bO1r0HPrbAP5iGFjp1YXr97eLoHJVzUJXqnD8hbjRNB58iya
Ko1h55C7CQHrEtRSwmhvz95vm7mosD3dIVkZhChm8JDqT9KA5simak+JIss7ZU9rI7e1DSsE8iRn
EJ7C0bFtxMYILaybKsO4SJeMWlAMC9ZQlmibOl5kowp987XrSROGzBSzwh1Jyr73qYP+ODCeDfA1
WBG/Axj6mKDk/DHDucxbfu2mm35UwKfekNxQpf90zMCh3B1a9cL+u4F0CiidySydZ2jM6dsqcIq/
QjLUosqpSot5910eSd1wv1KTXDo1+98J73Urlwj5ucUaaxfReGe53DsnNX8YCE34bixYxauZoD32
LPMaHirCFoguSqAONsk5Ei/omJGi77TjQkMurtfu50j0ehsKOMtzV4e6foMmG2ZIiY7gIjCWiulK
PvjjNyFtrxIA+SDnSbevJjkBvN2bRCM0w8VObQfEODXA2xy+Ra+5oPSkt39st8J7HTwZpMlR4Z/s
eAr3YdECeZUYXdaCgqGUsAs60+P5Vyk/C6vxkhJXOfxo0xOQrKVj3LwLA5G1yZ2CnWqsrXK8Fr0u
kUcjRxXeJsRgWF4LK09Io7yxyTVdHL5VTsr0gylwWRgHb2F534Pm/4gPZqWbhUBBsHZudqqr6icp
go4+tQXbgJISldUXuOA9AWLZZ5GYxXaQPFO439cWBGVbvalBM/qdMuAzYBShu8k+yxRTznW9fMP/
xc0DzCQJPQny766p2XNy4vDNHvgQzsiSC/rkZ4w8yOm+E/c6B8nZk/o8DTtSHjFD00JdljwlLFl7
Y8rVD4rIqHw46eBJ8i5mqclg2Nwk1ope4SxWkG2rLOzMt45ylg7evP/Mp9l5bmFgpkFNhvw1DIh/
m8q2UObqAziKAbRTKR3w+q0iBQUnkQGdqQl+0FJzIgSRS1mP0Akj8SvE7GrTQUvjzDUCvJNuMrrF
Fk4e0YnKV5H2wjUXPrJlBR0OgILeJ+rl2j1Yg9NKtOPPZk43sKUoSfi8A+v+WR0MwVChrcKJ6rOI
hwZ4syb3AioPCvWui//HycqyzHc61zwDSNPzoxDpk0hHrEYFRZMLCJEWyC3e4wQTlnbtY0MoDtDv
PMjeo8zvd/kGepo48DbxOWp1PhcoFXuARRYTUJJFPyuPt4koXamSHuFYq4t0U+3LV94M3UIETCzs
YbjJEDNyd+PIPXu7JT/IDDIDh5AgMylTS4Z4cCs0EEucNAHWYcFYDWDMrg7E9bFLC937JbTIMMK/
e7rtDCVHMY6tzrBSNEvhaTsTBVAEFqsTjwPo1wbSteORGAajYdUj5oTDiGtSNfMUqtKK8RF6VPE6
tbN6+tdqQNflgYoGP1vVM5oYUk52K7fyhFGsOBqEHiVo1MOX0j+6NDprn1NBhjaezR9hcZAiY2Sj
TiPTSJIfh7ZFhs+WEDnNbdodZWHJ2cNsntsr6x3udGaZ4IVztxtO2elbEkwxTyUvTPOru3HpJvTV
tl0gONt2vNEA+NGmwQCIfFz4rdoz48H77REO8GNY4W/8ijJ33mGeMO2MJoYBlBTfvy+3URUKPeqk
rgi1aQHMl90HscmEEJeQPi6RbFzOcLS5mn6kVfETpwjBZw9iBufjvBiKfcYAbAEtHEGGAxqLHKDx
yKpKDD07DDsVgevEdVffo9AWC9vvwb+v08/UUncbFFqYLRmNnfIHTUIOKMEYj5E+9f8xRyruFr/R
UJ9j3XkdrGZEhcvmCEMyklGuaTb8lBCJocx2ef5kMhQylug48F67GuQkPoZJJPaYhNZiQowl70BL
W9MptmcMqYZoAA+yW+R0jJUjInukEC+k/OawoX8dDHXOCvHes6f0UF5wk5dydvS/pK0MgQ4bsX3S
Vti5In29heOHaO+KywJRFQF0bIvev9pbjE6zFEmMcsmWhyQ2bYo/PfzdrzHThV69jRscpLTCpuKX
qRNUhJnfsUaZuo1rhxb860wCyI5+GoEDieaAErg8+GTmMpDl9S5l+LA28ZC9V8qeBWgG+HYr+1Yt
1SXZVt57qkLnSSBZqOq9D5qPYmfX9Wp20zLBjKCcZLY8hfTbs+nxaBPkWOWImutYJFpKTcxmB1/O
Wss5enGNIWg8Iy4cz9pGBCfPdNZI7KQkzpCUmlIYILiCv7mHK6EFWdCBN3xwultVg5TOHLhHTVi5
l4jvkqvk+fs7yitCGizA7mRdgOrhOEl5iMD693AUSIq26Z8QadYs5Byx484K8OXTyNTwlAcUWu1t
nRbamsZ7JZHp3YU+kGgRxRw8I2cvsIZ7M/EyBIDcF9hOc2OmXdwHkPnddOX+G3VhVR+iSNZMAk7D
iQzvs73/52kbY/0Rh21nPKSZ2RZffjjWe1Oe/snkANRXYgbRcxt6Co2hvKkXXifa2Bg0N/kdd9aK
aiIxQu0FA/afQXMEx0VbVE4q4lO16XKdoYrU059SCxY/N2yrgtC2RfKUYwekBMEElnxCC3rqrNYs
olYdSQJhhpmUdJy8cQGnEAeA062RtRBm7K7dSdlJF/Nc6HO1U1R+QBFm8TICT7forcJvLnZZV+fj
boSaRKHkxpqYfnN3IkbjNkvpTrlqaZ7LqofYAzhJl0gj3qU6GGhita3/HvWJksvh+u88BJTcuC6g
UC57dQxniAN4dfzScgYMXVVCvGJg+On7U/TqGdIWQFTdfOZGyDfMdmpCQjZ+MlogeIpTyd47FBHc
EkLu1VvGaNGN5rdxgVk+2dMOdlz6wFQaG2p3Fd9aS1gYRHT4V8bnD3yFKUZn36bgqHI6Q8s9Z+kL
TB4HaB51cz+s40cNXEJPcR25DVlXuvWkikPBVQFv2k2icggHcaHkDAKuqOnAJ4t6jR7lhFshjQGc
EQufdP2cPdmR4GB/TwJ2mN7A7BADnbfoaAtA/eWg3Ez+yyugcYCHxDhR/AioUfRwefKlPTRhVXz4
zH9XrWbp1sqWTY/bvcNBz/WpbQXI2NldWOdcz7cXqj8MKW6Odl70hRbZdDYQs/XzUTXvb5MNEOKq
LWO+atkSZ0jFilyY+mAjweJ7m8z/ds7DrVPdos5iSl6gdBWAO9ynwQxisDbEXwdgdu11s4CESnLi
6upcp3lXt0vu1bN3bZpw5LzRa4Qcdi1lR8KXrFezag7nC8DGfVpJ91nbGlL5Uurir6WB9LjPsXjm
MaseGCanrFAIxJbm7JIBUDGrfhUEhwtcSBPI9zAgKcePW/CJnX+YI4GZdGWxafXhpp/Zessmt+vf
hrNGq7Ds+rupLxWMIp9VDl8vFYAj6Tk2EdZ8WSYE4ss+t2hIHcfnnXGJ6w2roe+ZxWTh+dmFEXQH
FJobzKr/KzU8vDdhRS2PQd2LssuQ+zdpBXgLSIn9/P4ZPPPky/jB8anJ1wVcCJ4SwxzL5DxBnafN
9l+CPUp3o0PwJx7PPgjuZyBEMViauliGjvDCD9YfwzJHLr/bBWkY2I8En0xcQviOcvsVcAKge46y
Da/Ew4zrBRn9CklkJRpE1suRJNm3pMQumQr+hf5g3TM1AK7LVE5ivSJgnOOsfod6HZcTznGmrSIB
ASxoDLDCTSkkTjtjQVsyZtokuxNbjV6o/YyPcKg0100ExhiS6IDihE4Qc2dgEHjiYf5Wg9+KJKTu
Cef+cdmkSNwUXF2WUWqI+FC5mmt1o8CtrJtz5h4lD5JxsDf/1PEcYG0OAsjxLFSYo5SS9bF3PC6t
PL0yR3YiAobLEhdwrsML7x5otDGKSBnParPDJZANVq+lt8LKVierK7t7dWDD1pVW/s0WSxL2DJz6
vvs58uqxtLMuDNyP79F8NaWLnsaVJ630UGmV3imdE5BEeoU9bC1gltBVxSW5k1p38P8Lvrt+xDuR
/k6O7oqtQ5COjmbTKfOAGrhXhLjTlGr5LEV5AybSYv/Xwxksauk4XHupe+78908BhJ8s5QtthHSI
wgVbiJngX8pR8MwzB8V48vDbtyImm0z58Vu7BI1rjCV57CpqZtMezzLqInvifkXduqS9M/KNz3KQ
Viyf0/4TQM6eTAnlJpmztBpt5kyzmp6/mzrjJ1tbtnUC6UDDrSnGl2mUffAV9Sh1ESWf7ZCBzAOV
fsz+StnUjNxknamMQ80DVnr5hFnxNzyYm0ChZLwkesJ++LaBBx7sP65ZuMFwlGJOb6yLtJ2hdnwo
Ic1cY4SkCCOZKA4cutSUiCrPBDCmsGH0wUYSSsJhMFCe1dc2HPtyodhqfdL6ADcGqwH0tcylb8dl
9mzeyOMpLIqb4nYNcFnTSYwaGSlg95lSsicarrlAhzb1FWW7rjfo28CgnW1VxXrlqAEr8fejIhKO
fdbLbEShi/BDhWpB1VHxaD7afL6WVQtTCO3W/dua8iHV3A9xPg4dUGwE3A2lCyOEubXxvc3b3LHy
H9C7PNzGT0aTxHZOGMqj0nOuiaPm0PVtCRv/mduTahOgsOL/PxzovH2r/MO4gpmp5ityLelH/hMq
uv2a8tjMNiMio65OGfuf4hd/EjRV3N7xUuLJLo/w/OXw23j6opC4qrQanDINmFljdtIqi/+peU/Q
9cnF7dlHWHscIbm7zP7OIneCFh6MneNUVX5uJqd6SigJGTUO3vum5xoTkK/A+gTpK19frjWJ9QMA
RXTtUf7tzo56SVuJHGLxQYy88R/k1KxOOFlv9WPimZvgVEd67C6I9kRI0GG0WJ9Alko9FAeCA7Pi
Bv0RzTLycIZtrud7USpvQ1l0xz3hT7o+dzsUxZSH4f/bwFjboDyLEkeYlve4usW+3M2q4/6ZZUH4
9seG2Py7lF1zZThlhtGWrDENX2b+oPru/PkYOivnzcw8ERU+jVSKmZ8Zi8zviQWqlb/1CkOokdNk
0447iODYgonnc8gDvg1CQ7YZUtoyWgsbN98XTUlTKW5izg47dROGTwRbhM/0p9QOOTV+VfUenT7+
igmslD4HiLMmqsmtnDSflZIqXYnYNQbtPUIFTqqNXpipimmF38IYJHxW1p6Lt+ZNOQy3m5ZxhcRB
YY8rujYOnzDCY3QhCiUxVEXL0wBstC003tYve7AJ9nZbEhfVZ/Hu4GkqESalDI6je1cIq3zuLO98
xgC9A0s9Za8rTdwGNrsLQvWwQ7UAQk/BM2dXfI+rjvay1DwhWsObe6XhKB+ivMb4jMIwk75hnbco
AAc4z4o9ye3vu7OZhkHkZktwbcCo2jeC0YSV36+yGCMyysq2eSkJOoxpm+3Bs2dscFp9C4QJ+1vq
Fpfy6V8k4ro1m7WgWkzaeRXVYcDQ7qi0hBJTUBO5ee0Lsog3Jxw/8UMhqayMUj+5eW2y3sJNLW/t
kpf1CHMjk330U8A0fP9DxDBwzNPpCTV7zJmGQ1e3vKNxbqRqSdzC3Wjlg3KTn91i2hjOJvBPXm5/
3vXMGPJOyKkBa7Kul8/PqvhUsMaGo3mMB//jruf5GWRwC9WTNl2qKqdMbHV35kLmvX0dra2AQ7u5
IqPD84nunsuP1cNe8mixbfnkuwUmM4VQITGdr/m2ncw97FQk3XMhTJfl+YH0wu9Os0lg1lpunGiX
qVijm6ZgvM9DycAHkVmqP8105XmyQ501cRVcvgsZVeXR20TU1CBVUuJTUxh4CGxExaF5VE82kl5J
C7PkwQhkYNB8PuAoIRL0ISm+MebiSeZg99Mv1gn/3Y3k4ORyUaCUX2jSz+di13BEDkbh7iOd4iaN
9KFOmHFKWRMo0mgwLJt+D0j2vovyzSXdaB7CDIQuNy+hCrqhK5RUkg9iI7bpSRJHcufTKl+Fixsn
eOtd9HbqSO3JXS5+/IznVZg1JHtxgyBeQJMLn14oHpcGsUkD+IoiM8yOfyquTjqtJWJokM3FNB9p
2qrn46k5l5B07halGDv8AOVLxzWFC7kyAW94DVCR/BushesNEh9oMl3SVGsxD8C/G2Vpe2RCG+D5
5vi4/WNKXqNYN1AEtVcGdzGovJLJiP+P6dPRYSX4ZlqVL6ONgbu4goUcPTwVabIGouEzY46MJU1W
j8XS9zkpiOt1HtfFH15c05mwgAm4wIEamm4Xd/hF4ylD1DVsFZDAfR0c5AdyBex+nLghNfNsr780
BxCMTm3OycTfNksplIWYEKw23/Mu5O6XYCculGHnhL+XLKOQylBGi7EY90hVb/KW5XGuJ1dQeciz
/SOeLw9IvWFimL4sEhdW2nAeTnbkMHXnAzq6YgwAr0sA8fyYaIWZFKscdxpYZ7VXY89daDkJDXzU
dByjaNP7RHE6GwKEdqgdL8RA11CvEPsHKYt7cSNfuRnhKY58kFyWupe4vUUpwg30Xn4//Rv1kYuJ
/HsaRkXL/kZRKTgOPMC9Ffhw722lYGZy7dDeptGA+l35MzAgCqVvnG5HEag6vRbyBHXidHWRXD2i
J3TAkqljztsmavVFpLh56M99GHOkIeQrp0lbrLr1THXr5c44MS50vTXY7oX9Qmg7vTS0YtY/BIoG
url+D+4tuIveDSwYg4kS5lR34QZQp4YUKqapaXjG3USffTyMMtQjMVOap5Utywy4KWOe7eCYQyxo
Gz00dq1IaUP7yqC7affaDoZcntQDXKTFwVoRQTu9M3xP2pV3QuowzniK1kjXvIHaYqORrp2ySOhE
3u1RwuDxrbS8TrfpXoCkks7QpahopsiMiwQw6KTVZdq0aFpKLntw7t3D3QV5fcyHKSz3c5KLdlx4
d/4Rt2DCDyTcORJa+8NrmQJYCaPfj222CjqITDb9iYcHWQ3DE3GiucENywHnmfi38bZVTnorhM9e
JpGz4PJNGDIoewwnNv7kL828p/0hA3jDIpilsbkGIZIE2LozSBluD3dwy4fSYaafM0Um9BrXwm/c
jgIEFSP32Y7U+emiqUwL3k9IaLZWibmjYWvwvfaYd7QUyEdVCUQpPVqqDKO2+js1HqFRSMrsYy1C
VODkAZCwk65LnswKVuB64VWt0h/tdNogN9+f+WjLBfxYYEFjz+uVUqbTlW8yVjfzsVrj3UVGoGCz
H7Id+wiJocDiNOplnaTDWrJGBRSAWssItOtilvYi/1yXOTK/Tv1BEmTMpfHz8UM/Y1Ho8AyeyiDi
t1SX6tjZJLZjdGWUgsc+NCf3M01ftL9FXG8IhCUzt2qjNqzm8gVROwUPSKQzVV5lfmnK38rgfy9q
HhkHfxF4af/ELb6rNtI+5PB8oC1LoEPAq/jSJAxqTYD94TcFI2N4zJTFL0kOAcZAZt+jxJzAOS5W
37x7NeD4d4E82rY1SGWzeR7O3fAN26bPjpMsim0t43/OJYOMszTF5YXJ6AsxB/+RTS1NdwkRnlgp
Nzv2NgbcNH1AGnGR5okY1SJiwWM2pN0eaI+u+ie+466Ym8YqKmv/bN6L2pLr3HpLHAzzkSSPSEJ+
Td76G372xA672yfZOdHkXntuONGci63KgnuQLFkdnQicYDBHBhBWZHHNPXYEMEetJXSEfrAe5vxs
FkIdL+tO2zvkAsaZ/KowfRTlL/TV+xz5sOVm+OQ2JM4IWHkuDdNt64RdOYBjbTe1h6aRvlKTE25H
VE8j5kcNqNZDrRHcJo9y9oDkzRAisYVTSK+PNCA9EAv29sC6+z+PbIRDDBJsHhtEdNAbq9GHuLEL
7ION3F+lbLYvmWIuhtyApea7eAxdKgsyYP0R0baZIx02OVBQ9xvhjJYNf3N9UNDvKatmsJWcPfAP
7t8auNHWu2OBWw2Tk7m9U913De+G2ZjmWkujFx9+NjbGytmD5CDqT6E+G9BdJgi9gWVhJHEk0uJb
IkBRZH/ILMuqEtlHs5yvphMopO+Yd1ABbz88J7nXv5ZYccAKB57KdK6LE4gFfXStdE11xCj1qqoc
STYSTiXLXsdWS30CzQoOJ0iLA71n+6pHd9DEKyyG+8dseHyEBFPtcFJymziv5qOsSZDOhTxoH6i/
CK4fEbQnuy9/vqtdA0I7F1B0AU6GHeBW3wAHdNakqt3eXJdn28fNGCdQ2o+5wOYG+OyB4LkINchT
e7H22S+a6zgEaEcgCPfSTektugnsEuUjkKJn8avQFiemMidLlR6S2mwy3/RlIulaLCMuk079Bj4+
vOGzIBu09cOft1xIoPWA8iBOWu34Y3X6DhGadgK6Ckd7ts91MoPirtmvDCGM5WZfMMfY40ZEGgOd
/MWsCLN60qNvr4fL66VWIZlq/jpVsXhMh02sUaqYr6vFdZET4T8P3VTKU0CexMJ8PqMHEgCbDRMj
IAoURzkKemetNPYQX3Na3dNcR/74NbvJ5XIhrhMNiSR2Hn5U5kKWMNYpC4c1xTD5CitPu6k4WYyV
aEZy+i2dZtyJBr5cJischLh6cCEVZa36i/0XHU1jjFW7j8DRpdqc8PRbghxJKMroVXpIOlK8eDiE
+SblcnyQr8DQgBnUjlC+3FNp3gGtsgASfuB8gEj6Z5B3+JV2h8XvKPQFuTT9ztMOkMkctE2och1t
FsucbMMzsVRghcCZLmXzUSYwMg5riTtXLaEmlk7pVP7BoNW2VvybhgibtToTMpS2vtUtVlZJKS5a
u8Ad9szifdOCRXbp+ZgTOpxwBnw30S45DdkRnv0YiIQzu9lNMxd3LJa/fjEPzewk/vsxR6TqxEzk
zZpI6s74chNlLbyrC7cRFnHAmOwJ57Zn7vMCUUuZLCAElW8ajvJj+bG5fw5Fc2sa7ZWGdhg8nSw0
v8BQ93UH9ABMUUsqWpj0GNJ04TSlTe1PrcaWfC/rHmxuZZJqk/lfzN2DMAOoOtTuIy/ivsBbN+p4
Pmj77iKW4yIxuy+mfivDrAOLnrhJK3b+nOLdTWo7hDYV9ZkCi0jubEuB70Gqx0m9lN2+ppOxQKIY
9RZTfL8oK0MfuqwoiNqJRTjek1uRCRs5HDhwlRNEsrsZsyauKR+XiybbHpQdZOWeQqaTk/3pYKZs
E+QYvRR4hoUlmTttw40kdPX8O12P6k3tdoWlpyMuz5uDo3+OvKQaGKu1m79yA70qDu/MpIPmYD9A
XqRE/vvUw81mBI6lIgklapJ9USj3+WK0PaMH8Hr8zRzgvJ9hUhvTawldg6Qt+uomJijj03KRIaUK
cRkw3vQCCQxsJfWXtyWPBWHtLBZwWu9BwKlL2topLSl6/6TFp/CKl4cLCQ5sBVKqTji4Ej+RiXB0
A/t6x37Ywm0n4VuTO1MfLlvh4pxxiAK7atvR6Mb31ygas8OgGkK8JVgjN+8IVfB38zjtBR8ZtMMa
YxsReQq+qHE0qyh7Yey/rY+g5FyNg8Qw3MAdgSkslYeJBZZGSHXFhwwhAhdLJM2kozIRvt/X6eyp
kIGUFfKlCEHAZlaOnHqrQNZzOOf8dBzd7qusEs4jr5KOVOGOprCaxaSAeov7qmpvugnLncVVtH8o
DWCK8x6rHff6tMCHAzoPj5GFp2TwOFtALM5i7E4hrFhkJkDvyGNlfVzjxbyKpvXC4KgnJE6lvzPD
i8TdJ8hhbS6sP1MURtBAOVzvqHpDeGw6AbDxNi+qCc+9iMSQVoOmoX1wxhOMyArsTgQroUaZCU6q
9kCX7uD7iPdAc2xImpdwshg3yy0VLyX5gm5Ct81G1STNMaN6uNIzOdDm7pb0KEk2vp+qk5dw1lCE
PLlGUdXOWAbnkl0urH6IzeB5+yLRLGUwGTAam7DP0E78WElzxSks1940NfldG/7NH+12+psoUbnF
sCR/GqDt2WVqve5GkQrbI790iDG5w4dV/yo0J+qv6kncZzOqV+nLQH2FjUo904VXjhZT4m2r9JtA
Kco8kiPzIO2fQdO01Ngt65pcNWTNbzK2Ze+MVPgNacigaxEO7ER1JwdK+W+XVQyeCRUtR8v2c/YD
Q3kVp2WcemUgEIVSQ7uUmuILT6vVNBNgOjTUR5OfZo7VbSP0iGT3fP5hAfCHHJOntn4cDN2K6W+k
neGDg54z4L5W8eCHP+T34URQazOhzX6dQyGtqt168w5s55eGzpQ5DCtOiPE9m12Sncq3Q4hTzOCo
eBcMJuf06W337nRPGNz84/codugQzG3O7BjPOrKIslFQECtFP7Qb9UjMlyQ2PlZpPNN2gGXHgEPg
iFPaVhIjOa6Uu+t3sCnQodQpyEP3oC6277iQyeDtaL4tYNnVCsiyeOt42Hw7Ry99ddUsWwFVY7oo
U2tT+5zchzW8pyEBOWA4Z6s5n9nAzZ2LBkEg55SqYsR6lt0D9rwDaUdodfGdLZFz5sM3CGDkGcuA
yo1J2cuqT+HHSlWgjIz4CosH7AwTqUXZMwC9XVkAjZEOIoo79xBwp+25UhpgYiBlGKHsA/I8HDvw
VcUZzbLOQej20JaOglXTWrNsexgq8PYEdZT9G0o7aKeldt+zli09kNojdfeZOevf4hPAbtzhjLob
pMAkOAkY9s5NosfS6sW0pHo37NVGIrCQNS49Gr9sISvs/mP4HnLupt0dT7tBieERk2Gbjik2sM2t
sBmLrOgqr/SO+L+wA4Q1KTeq+7hyd2AzhYuRSXGSIye6Rd2TLc366wqpDaZpRfxhtDsCz38z2A5Y
w6cs7NpvvywkLHr3msrFDQFYYtNDRHLh9fP1Z8h1rh3J6v13SGrpG0ZLi8rSIbzTPRfkGMVMMZcv
8kvXzB6DTpWsHtrdo3noZfsP64zGWgiyA1Du8DWX5hb4EpKeNCxMkSHaQGWHkM1q4UQ0P7J6inhp
CHtJDBod/diTKD4pJvgYFQp00orRXIsoU/SPrlEWoFlyeiUrWK6XBDNkOZC7v8vtnxO8YwsQ2Yrh
Ad/vZHmy6wTGRWyUgzMxqba4IJeNl6+ZuAjGvTUn5fYiLQmvPU1e6HgWnW+BIBOfbnX+KoNY5NN8
M3CntdijMt+VPLumkfR4QGpHimwqioXdaW7aFm23fQS/p/mMLWiuQ2gyJVgP4J12vuNNg/P4hrGc
4tUaFCjcSxpXszUVX+GZn8GAMtMN16Rncasz5rYBlm3TK4U6ayLbfdGNeSX4xahDiamgzG9zvMaO
pJa23PgD9awRgQWo/p51ymM7fZyp+j9tD3CjGrmq948ASS6d5JuTDNajr+cl/oQ9RkJpz8MJw0cK
mO/p0n7LeIPh0dnSl43lCdFWwB92OWBbDTZQLyCaWJ4i/91uO+/JGO8VMCiJwLgtBGcCK46gqt7+
4PqEPY9/fvHm0fLIJHen4W9wwyygk/zWpju30WkNxSTu7y3c+heKJWts7KEYHuztLqqJTVK536oC
fh5UtK90E1HdnK1Sh5y0X5K90aAQt/BUwQ7RSgt1rU8llRnKMHdjzlcy+/tVedtS1m27D+/0dn4n
WotpX/14gZm8mFP9AfCUctOLKxYGfzkz1IwkiR03ZTEJ5FjH/I/8SYoia7g6F25RFIudsnZS1Gna
mBtrYpn/MTzMAg9F6gDo6Z6B6Nqmye63befdKLwya2ii25A2GXCNCreZ3pDGxWKSLeDLUZzYd9XW
Rr2b9JdX+NX3aE3vGOU3c54mVxExvt+o8P+iBGuZxUP5TCHK0jeVQb39xdk5l0icxauEcYrBQfWH
YkjLAm4+AXpIqKYTtOhs4hhoOaN3nbJuXEh7UVU7/IGkCT3NAC53mWtomvFlKaszcFgE+lO3x3Gm
tewHoJMxRxfNo7oKCZ/QlrCciQZAlthDD/IgaQfNf+DmUcqW95AbfCr/Y1sE7dyJDPCdAMpnxCs5
6uYTPptOkmo6hxVz2Q6fpKhw1LMvIrIhpXUdz/4Uj6dWBp6cRVAwm3pgb6LFJoGk6Cqfq3K1GKv8
RWYh+Rddw/IwmEzrbB6nC4mm7XAtGkpPr/RY00Wo3HX/hCycu0Vo5/6VXBYh32jMgcFGEYZ9bnXK
VsBSWTQiu8ezcmQ7A8cfp0bYFFmoPxNjhYF22awSUgLEurAlQkRAQSsEM679OULfUpzIb0aNklBW
NNw77UK/NgDtvThprK1VsHOCagLOSWvYpJhnRiixqqNEdSCZuUUJAxF2Mv534f4x1TLdrF6PzFGC
6gbuydBURWREVEuAvEkBzevuseG2AGuSiwamA92dYr4/TFK12z32jtFdp7s76i3UriWJbMsbeD/d
n8GctXC3s7UjwNU0H0U2uGPbX5BuwKS3ADJYYFpj6nXPCIztkvswMQbA+bXRKTkSfT5qHSy2kpws
F+u/aVMpkWvix/N9Jwy753JGPdDFjn+id2GgFD6dxKD67ru8Ty4cEdiO2n/2E1wdexRlUhiRj/rc
ZYcdsZlj5EO8NhJc3jcBE+sHURfTt9l5JtEETHpDE6RVvMAxyrvEaq3HLrkPoKAll6biao2WBD8s
17Lu7yPrP1KJI3YwbAlaBDM8pNwUchvudgomep7/g0WV5uT/04SNAwbyF96LFYwmPUJHGRKqdbVj
RDWssZfttRJ4Y4Q9Q4P/DOq37i7NeS1aHF05WRDWXOUTtmAxQO6h2q1II7MqdKkEmDSXdnjBFPIv
kl6yxUZ7MrLjojjgbOgheEb2OgMNoPz5SSEfKCinbG3CIRjUoGBBEwUH/tepPoIXLT9paYYqZgIm
gJ9lYNwGZuGu8YVxHk81ce6pAUBetDlPNuIZQXj2DFt3jHpp2oxNuAPFECKJbWNL61Q+5/wPcd64
tEJEZ9AnvWC5gEsGsl8CU1hnsW6oRhc+iuT1GHvRYETOz+oFua7f7XZyj1sQbk8XSsMJLhnvlFdA
rWb2EmOvhb5q6AE8I1gBXX1notEilnZk/zpTSE2hqitPq+ZUBt60dAY9FUKCD9s2o7CgCuz6EkB5
/lwYJEP3T0Nb+OQbSAsxiizfgchhHIO4x2Hra/toHQjeeibMVej7TTchcwpCut2gBiHTA2GXbTrX
mEe7CRfl8cRkf6IYX3oMrUrCkYpAXClDd2t3b657NC0obwtkB+4OUxy0w1g9J6GCtSodSeXnmc5M
Rm9QNzWMDo/AoYN23aFAlb13FZPUSTmxrdKJyls3q6DukrxjKmsHPitpGQz/yoEMtf/CzcCMCDde
1Lcj+3Ogu9cghOA//ZWex7Aw3D5ruxly9aALbQAsxsZJReNW1uXa9Zbhp3mPLf7GrS4cDW5IU7YG
dlEHm8mcCPo9EQuVDc3SN2tJwshfM/f0Bgj2x0h50D1qkMT61MNtF1OjUMb7zqJIEbMuwtFy0pxR
BK+2MQvP1LJmnX4/V338PZcwJTArWtuSdLfRPwoq1CfY7ZOQrj7q+5ztpyD/aYSsXOKREQSOxy/u
dyUIym9+gf6nq3OP65CxBeCMU8P/V+gmoe0J8kTW5bI7LPdmSlh5zVTfYGqEhHDjQjPnxTcXmev0
dCBzfZaKJ0rhzKYdcoM3hidPxczDVrcXx9a657+tUyNVOWnCHhHl9bh/Ly1kctr4SmYvuWvUuw9o
QDxmDigvIDXlIsk+LBNTSMz6SiUGybRrNCM89ANsfoEU5i/FQVXSYiC6CIqAIO3rcGMGYHMV2HlO
gnjLApfWYCnC0OPJsDBZ8r+5Gqdbc1moV60KSNAhhC8Ke/jJVNOoh6NSlPD+oqmWITJy0uO4OqSc
kcwuN77h9Ir7MmHLGqFFVBGFMLvygaJVqbrpA/f6z4FSvMIZ1E/iYE5fN0M7Udtgb3KmQARLq5nZ
C5ZPA8veQ3OJCzCKZeZ8KqrgmY9atql0yqHhIFN14iTQI0lp5eysnoDqVInylMtEq34nd6/CK78G
j6EAkLSRozmGg8buAdJu2OmxyZfWpZZns1m35UqxtHycd11tkMp+7H4eANqJvHl3do+c8/zBjZPD
Ye99G98ePm6B94FkFgYeoA2syw4k1eAc5ldFKD+QdTjZKOheYbNVssyOZ6Sp1h3ZH5iB8/pRzd+j
gFTRHDnHLvwNHCHVlfNh6WRiSJUujUtSfaMgKyxIRPF+PEW0q5KGvs3iJrcNta/4i97OyNKvMnq7
pQbAOxjdRI3bpDz8TUJihn9oBf/7lNUNi9E5D+2TnMGI5rArTCVxGPMJmz3BcZj3d967Ja2rgetY
9q3VFeGvV2KnBENGb9q41AbbVWGzR66Y+JHFGK93+GAvyt+A8gSQRETYolR/rIVrO4jXqytfHiTn
AtozpRfxc2c+qzSuCkXeT1chCBVblW9fpEtfvRzYax33E4yiHAsrsAkWxHQN9vH45UQckbl7tdXD
7lRDl/6AA98FhCs6LD1ZYb5JrHrOyBDY8gBQp9PrZwU2KIpXXx+LlG7zegW5HbupkIXmI6mmLHw8
PxkaFC+NVib9o2IKfIgs7nabF9n1Xe0AgyEM+2rcV0tSzgsT6CDT3SPJA3Y5hNe62LAUzij19f6H
2wBtg1UakxF86Bt35Ld3DQ/EUgvCJ1fIMnRFfSq+xWb9tfr3vCjq31HsEg80dNgWtnmX5584tn91
j8YGthZks10Icfu3cinOpBJbvi+c/cgyKgX46OXRDER8uG+aBrYatiMvxR7rNPNSsgpF0TS1x36b
mYaEPv5jHr7aDDrCbT5D3s5M35vIL4T6wT+/lUfa/WucS0/1amm+9i4VeBq3NRM0SeDlv4R2vl7S
HQyZ7azyARkaLR7dQmNxN/uLt5S5qP6znkmyk6RBzp7k6UIKec8JLMw5siTQPMMdwC0AbMpuwFGX
TJelTzlC0TfRRZJ7ViotlX79UE4qwadkDsen+NCUXoPPlFj+iGkNU7EKWAPo9WCSkplS2/sLgQt2
OX9OkNTFn9d/YufsvD6uDgyaNAZS6JknCU44uIzdE7R/7+cX4v5iMY9Ctgt4ICFxZq0I98Te3O6a
iTgyhktfYxegmEzY9VkH4N9IhCqRsoRaz1jgqJCsOIZUbR5PZdD+zFGMMBYv1LCxQ1n60fAy+MuZ
ywQkwnSya9f2yM7XTmohVC//Nps0faxSsd7qg8zyZnCe6lgGuLHz+F1lWg9SrMxlWhIS+XfcBTO5
8cM+07v8ZR2gPAMWCMmeSCRYed7893sZAU0R0nPWGMQ8fqmsiHrxhgL8Q2sIpci7RyIJ+VFUiqUs
kB+60T+MqbmwlKSsQ2jJhT6o+LVmbz7dopmi3wl3AAh/XayxYh+bA1fh7+p+f/UXe7CLBPHtA4AO
HQGG5B4di1x/f5gHuZ8D6F2pD5nXQ387AaQyUFmM+woU8yPhjO+G72OYA3iFB+EwKsggModSGIz4
Cn8/xru54C+htG0+X2BP3Js7FR1ZBaJ6EcP6dQcwywbqPd0XscmArKfkM/aVlcHW8MLzd8pyqwz9
lGKqosWAfh7yG6zaKiAbQfZmxyLhpf+yW6aRy9DvprykKYokwgCt+64bGzzHpxOxpsM7hW+ZiYl5
67Ca9UcMiGhX+hl/NLdOdVJePvo51ZE0d1se05G7Qa0r0nkA6U25Ks0zX/XmP1WY0InsNXwoVX7T
kq7bVTL6/tsE7nLu8Hx3/d0I3X3ruQrtUvcu4q8A9DT2nfsV2pAUmRRlWCu83aRNDeLKifEDRWos
h69Yybc8X3br6htC3k5zn/rdQI99B+KW5iPy6RITGdNsPOk5uE5zE+QoaMYgzfGU5mF27JIy2gnt
MLt+Dzfe0UB9KPDmKD59cUBZoJUUSp8m1DIQbZvNnTU1z4n/lO2CoaEIz3yZ855XOuLyF7Cqcs12
wLKVXK2OCLsUkKgUhBiymH/xKXycxRW7NbMlYcntbHg4Byw9cBR+On7cCTwzEAzO+etHs0+lo3wr
l3iZH/3BxlYC7kmCDEiHXhOuaVI4+Xe/K51HF/F+C2vdxJEjaL2/sdh06/5CCkXlreiUw/Pbo1AS
+r3YmDwPd0s8J6nBSUjJgM687Tvvg++h8Jl7ldHz1gVYnsTmWi+1UxuGWlgW2KsfcEijoj+w5tcz
o/N3Sgfv3+LpS9w70Dm9PU0N2U5s/B8OO1VhzgR6nd21Om9gSRq/lieJWSHLoxh3fc7mA2+SYNzd
OpRg792+7kk1urn+6AN8Gzctvii1WAbBH8wzKebyGIJMpw/7quHmBL1YrN7O05xgl76lAYC8bt8d
dmcCO9Qr1SpaaUYgA7Wk6YPCqW75nIeo8rOT8F+FQV773O3lvmzCClsWqbi0SvwtfESxAuS08h/x
YYos90rkc2Bsag0ZQ66vERFEfSZcZt6mywnMP4Qk7wZp9AkyO+LwT88iia6/tX7GhZwbNsKRIzMb
tDKfy+wZgZJnePNoyrkez9bHU8KZ/zBhT20eb4Qgke0TVr37egNB7d6zGku5NpR9fPpo8tqvgP9J
hr+WIPbBfUCVZf2KIvp04KhPCgrZkLKsbiUvFDka8YrDeRtoNMyfd4TOYiyuXzzwLy10JszB3D5w
dQL3pByg2RXNgoICt9UnzLC6mHkDm3QyF/CxolBFSzSvsmfKvJtm3Yiap30R/DhwXmI12u1q72QT
6WCJGOZ8zHII989O92Vn0ixDBfmKc0fp1sTkFhZqAqCRGgY01L9eR3ZEYpvftWi5xsmvXSPPRAXd
A3Klu0m31yDfpPLHytD5JUSJ1tyNRxQXhSaJyZQC4dUsbMObP/Uz8W2x7pkoUpPCVVlUa1GEQI6e
nb60O7IdOtzZK22LAie1xak2NqBSoz2/eD9XowNlG7CnO3OW8O1Og6SphG70r5uVxDoaVx47iV6B
e8BwH217KdjDFCbO0es91gaUdlM4UvXM1AEo6YRBo2joxLjV8ClJ2ORnaIZzrYok4Ej4gLlcNLoG
oK8TnLMf7Si9vhNaHKwvKksoa/1iU54zUQpW7GeD0nSJgUkfYqxJmY+CSA9n1gc/uIN9v+tejaqi
9I953fvSsaSmChb00D/lgUdmbibINk55DbmY2ZVJn9iGQj2x9iktaR5dhjhXtefHo/AtTqjqsJgc
i+zPZez67GDkaNA/TmUMIJHnzUGAmDepx/6abbV/Zb+CKsT0J0aLsWv12qBYN93piYTMniSs1bKR
QaVsGR44yUOT5yS+L7oURKv50AisuK5tUvwsrE/SXBPGXSMs30i0XVOMdz+YLFsRg5Gz5plT5Deb
6/CUrOQLi3DqGL2bDrbUAJSqIBP/2wvShu+yMF31JA10HYyJRT1Bep0JKxyii9gKqy1We1WiGWvc
6garO/4RQhetoqSun1YAybR/dMw8nkBNFRX7jdTHFJ6Fbhu/GahnGztWHXRxiPm9g/BYHSJo+IUU
BVWjNtSftM8ChlCTs+5gyMYRg5Wua//a2rHrqZyzBu78H6b9I9plk9X1hf4FDS5diJxfSExzLdaB
vvCM9L/9EraZMhbogN6Pz+OiXlqRRjwlNne1y/ROyfyVYPll6yGSqwQkFaRI7UYKR4h6kzuVhcg4
V1cxpY+XF0nV9Z1K+cqEXtxs/LwvQoKPZFzepqvTYbt2faNoF8wBL4SGKSlHHwMbCPOCokuC/xWt
NwK7g1LRtZH2vyj2Mvz+rT58r6N3u9S8EJW9GSGKb1DvfR37fwtzNd0IyTitmalrpmdemHUnWao+
Xdyh6YivktmjvakUVr1ioxPT2iYKvu6UGH/R5IRvEpgGGH04ajD408kfw5oOTXqrzKNKm7zsVnRY
PZu/GMUiBoZaDD8Epxzgm71LTxqFLY6cv9jOmvnTSKH2qVMUa9zGUeAAj9y99gK2g+adn5YBZIDb
L56bnEh39K+eK3CediKWyvi69sZj3G2x4gRmgWE+wHtg1tmSSXxn+HAitx8mkAJYVUJJdscGm7/s
bar5oNgNeNfflANAB27dglVBOUlgzNtVytFSPZ8+E05rmVUfpBrlhibeBWmpNHzGAJIFihND+PhH
GQbhTmQgySkL+SfOP4DuIHfcbtvLl46q7ERkcApIYA8HIMaBOK8UDwGWS6EkfYQuC7ziSajkgmiF
DUJKvsCuC49w/04XUmZOas6QMqWyJgEr37aTsORfo32dx0ziM1tTQ+6o4FoDmJvRKoQ3M9Z0nc8K
1jrRr+D0f7nJhd6HrjybRAbOasbgGg/q5O6aRlktTU5oJFBj16MWiXkyzo0sbktNSGVLpWF0AJYr
HNXqaY7k4QdVlj5k6GYMgKTt9idHqrHj+zfETZ9WXhhfFUZMQDrg/mZ+tasolvMSSbkUF/JFXr9M
pB11gtOPkJODThQkr61/EVSGcjl4ys7lS0/icIqTG18gxoP4dlmJ3RqkbBJCOX5RxFmjHLd1ekYu
Rf6IBGMo5H9j6nKX8uxDo//IyPtduJP1fNbo5oMmLywh3QrPxYaZt39QrM86csI/igt4BNOibu1J
rf7Tm936v0xmk6auLy8w+wyJUzGU1kLnTThHOHGrPK5rgU5+5J9zEOCE71FOYLrm+y5/xho9+BYw
KAa1HjArtRYjznyk+4+mMd4GWrC5RTtc3y6lJhQlGip7ROBXYIAeP19cy5AiFwfEInFpR/6dm8CH
2FoXXZtTLoHCvLBWIWZe8Hs4o1AzZH6wJ7mWHxSKLQnybnQyCwpUV1ZA6wKUM7Ngh2SINo3pzuXZ
EVwB5QCTiobd9/UhR2WExEhXS6445n1t2fzlsuGrkQcIAhNKupHZHq/1zhvkmcU2uqlfZEJE1ldn
Ytx5KUT7M5AwR85zgZHoETBDo4Kz87UbnOIGMKOA7bTnAJ07hh68Q0jQe4mcq3sOPX2Uj2/j283d
8sNy4tcRDmrvDfPQ7Jsy8sza6DNUu2RMQex+ZPwvbBKyMn4R7QLsRls9+7O/OzHW3b6NAUjbtRWt
RqAw78L4sahUxSHBm1rLJX7b51V8Zuq8fPSGV6iGQPuRim0GE5fJN9OV86otaALr9AMauIbe5q5V
LfcebggwDhlAy+rxKtw3E+0d6cpFbjGBkkor1EMFQSjw4GmJh6iqWwq+6rs4+FWwL1LCmGicFOJp
hvuyJ82UXNHcK/IBYsth0vPOBc6Gaq1WEIGKQFQLiAZDJycUPzgMYxWoyhc3jciXSwlW+WiA8i8I
Qi1MSJMMxS8uiSdKLzHItFT96w1qKQa6hzH/3CVdd8rD/hdVM2c0WWE6QJPzmMK912BG3Q5GWc5Y
6guWHNlw1uZVhCSxdUAMHyH/T8oPrFMR+vcvSLjtPzY4jFkTEjol4U4yDok200Zjg2Xb4JDaxR+U
EvADUO2lIgu+R01lnT4+8qY33znWpmW5ctLFn6kNLaFycsHuS8seANlK7+mwDHev8EYDP7sFxlpO
Pv5BmWEolVOgMybo/xh2V2BJwdeiTi9WkI5DMMj4S5WClC1zNFo78Pi+AMMfcDW9vJsUfGHm4KUX
NuNYvoZ9stIwVhvrIcQSwepWBCJidhWnDAvO9qGWyen9YHuY3AiCC/ulw+5sMskcIWAJY0Ip3ie8
g3J9uosnqn8q5Ea5ViHGGFhzj1Pr7rI2oKaRimM8XuORpvpPtsExq3FM3AJ9nQz12wIRHBCqs27q
DhNNRzvv8yEmsctjLW2S97Xm3/iYu51qx+VpM6fL3y8WGgqnYw8qAJpYznCnN0Qh72EX/7VOHct1
tLXH4XI7V5nPsKH2F9Ua8OxcjbjqlA9xsgYPD83ktBPazUffSFuJJz6fzNTfERR9EwXSDCovzMQ3
i1wBAI7P0LQiXYKEr5QGmDFNW+YoPMm8Dk4+0cJjk7+dUJtnuSHKP83rfVKAW2frKVTRRSGQIrHc
JdmbQrIFxWznGUFrBYeIg/FfiwcMxFGiIOmOv0rJNbwVBhTW1O3E8j4yX8BMCiRfMkKXVejxxc9q
UX/Gfy0cQikHQUygz+CN8CfaktEHBtpqZqwoH2cilU4QLzqJmCZ0ltNWavTy2gg8YftZW6jsTb33
XWps8L4x6v5ufiWd0959MkksPVNke3/uOynrpqXLGiQKcAT1W7qXnTviET151FtiTC0E5cgpI8QZ
nC8c7oqUJtxrvQ0KVbnK4TFSclgKHTqUdBGk7nYsFxiqDrfklAznDKyfmy4TDiaUbeCQhHwh9cKu
++kboU3CY5fLgwMTOOsKTdwbIQLpCS4S/WL1SQtpEIT49H7biRFazvZsYvTrdDimJCt9c5DPelwC
BvnRLWbhAN/c0l8vLu0wDiOA0iXgtIG60HDgcTELtd8dIydovEuYDAvQz4+iDgKPsyAuFcueAN7A
mECxC0cMyUqp/2wF/eBduWg+hyzU14z9wDEunV7XOb+CCOyFOOZIPTZHc3iK/t8PvJanV0I61ibD
MB4JW6k2AFB25PBbhEPwp+3POZKYazVZmbhlNDck4l8wuClnBS3/qqOagsP38es+Z7VeOseKVVB+
m/cIWq4b8o/AfWrWWSguH+RXhmpIXy2SJwTF7EI/VyesOkcgMYOYh7y+K82s9X+3Ca/+c2tFUmbz
sl/IstKcyTkDf0607j9PfDUs6q2Mdcmutqi7r+wAdc0b/G8DQECE3X7NPpfjQgWDCjxn56JQdmxT
JcJW0mPG/nADRGra2QqrAc7e1Kkd9+3LXxD3uawOWjZUpCkmQ8OEUub/J2HuDvp8rhNh3l6av40b
B9jYCO+R2/ztS7nV3LXUa9piyEuDAEXZz3P14urpxtqD0Ni8L9TUjTC9pfPJT79r4Kc/WxMO4+s8
JPMLl/S/wdq9cW2GYsFckNo/Gy4rFXmRZLLSc4rgphiGvPTYEv2bRM8lwr8JOWQoHoO9BeGtiM3E
8BWTwwaEr1LooHVwK5SX3ml2HqwT1SjjRUvWSVOV3kcTEP4ieHhkdY9KOqZ+5NkedMa2j9ecbiA0
ZrEDJenP6+sDLb4MgIPIP0lF+iohqY0p8Z5RlD+BNyZvKHcRGLMQ9XTWyrL8wAyZY1lvHlDf6ww0
0553tjZnaE+5/PCBsKsaZY8fnRlsDg3sLcnRR2uMGF7faEg19RfvqLoslHmyuAobAsFA9ErC8EvP
+B6ehG/umVPB578RrjsVCPC4TUe+rgozaeqzBnwJuP0MiQlOPkRturXpRuglGxfffCDbszboYUhP
0iPvxZTqI67srYeUyL5b18Q4zJ6q/DPmneMIZD+IYU/XZBDmNMpxPoeTkjeRcWXJG6b+lS21iNrg
6EWZhmMX1esoCmRf1Dhg9a8KXpJPsLLNGaS8gAXcWyMW+p+oXDDMhjyKpegisGUcU5QghxHidLJr
htMO3IXPfEiFKLcL/zrottvNIx4aJ0FceQQPGl3KK++o1mtCFI1RE+Yz+Q9idWKzkXwEfs3rSJQN
cAqTNY6az/B0iXOn+kDvg4cX770ludLqoQ9GHtj+jpxCbc88R9mjE53944KMf+2AdNA1ZZs/4DaQ
ObjApvSUMvKQDPP3xBwT9Gk95sMdhueqXp4r46X1qJMD8ty/6u0b2lQEoYoiNHKSSB3GICdL1rKa
ufOF0dpaJwyNWOvbErzJcToowqc3AXSxhzDo4TSVjKhLs3CbpC6h4RBH9iBRJLr62fVEzA5P/u2E
YvwLae+f/6RMAZuk7qAY4WHfZzfelcHFEcvyf4O2oanXLdGNOr297LiQrPkT+3rxQ3hCVmu8nZKU
36NN97crvqIEAMIqbAgZ6fTOkHxU+WLjIbeMF8bKxuik80xzj8JRuV7anaD4Vy2CEPtq2FzrapOB
mh2AVOnd1uxPIpw9SfkSqshidrEc1GvDYBVbDhlDeR2ocWxn8OII9Ka0w6NplLWBtvW+xuhUphcT
lQPhtTe5dH9ZcSK4z9kp9kKBY0ttA39ZUd3horF2Q1uDyTRhdkJ/gtN8QySMYr2+XywzbDI5iEhS
wMZKhsMU8AxJkVrQqOwkoDVf9eiBPwwKJwyZiAVxgR1XIR7W3zF4Vlpu4WvIZTeLNaHnUD9e5azu
hP8Dmi9epJg13pZPCkqZ6X/IYFIpr6MOGagC+sW5kIoKDq/MgVUBW6QtBhOg2Fw5AgRdP8LinxW6
DqpoOky5voT6C9O5omk3MN5YfsBSUt8iwes6W3PCRAOVqk9sYei+YTsYoGUycuLdoDSqai5rVc1j
neraGxTQEvTFptopLQYAjVAHyX3YXFSxfCYh4xoJc/I+o7A8P+0ZjPbxpQpPCG1ZleSQwLpU0SEm
PyT19SAd0sMZfTSFINE0YQIr08s6rY/s/SE/c8JVLjbot8FPMvrJUUjxI8W9lt0ULFpKACRIK56B
u1Sxls2wXQ7BU+EAuBbwQMJTFIzkAWLt6YLyjid1FupTuniTtaVTP6TyPt16QgkLjBzLvBz+Dfjo
7ywmir2kL8E4jgTwzVC8tSSpOmGLBt6iw4FpkzvRQAhDY2GhC3tsLbS2DhRUDTydOD5ChaQCjQET
gmrY00EuGOYNPXI4A+q1JozRSE+2RMdZQuqdNvWU7QPZwOrX2lDFrG4w4kFDG39kSdJokKtTzUBt
EeBvH6OxgwBF+KeI2xnqdgA/0ECWbvmyyehQh/6DmdPADUJGJCfUADAv5kih5PXsl2JesfSJw4DB
Nxxa5LAhoDuPY0tRu9bobqgBtbgLqUt5iCx8qko/WI5Ox3/s5dUlu2TxspqENMkcDJSvrmtzhp+Q
GEymG2mFblAw/2/MNmo2iRd0oP8PHwoo53UtVju0N+NLZOe8jpU603eUqSNq/YvlcxDTIjM73bsb
Sv0FqT2CbsIOpNISuukJ6/smgeVv0vZO9ZOij8xPnd5yjHcM94CSquhBG++rATBWSNSMd/5IaVH5
qVZAYQSWU/smTQSj9/23vJk6Vs6Ee69SfeWfdft0k/FLYSYTuUUoHQzj5iUCIcBY/hYPExEg3PXr
RokRlA2Z5LTCT2QHtHXeE3yDQNUN9N3KrDzToXsGVVBQVDppocyIcIQjRq0WZKkfKo/WbtK0ZOaD
8S/fIBKXFnw3/50206fxd+HChbNRY440SUJEPrl3rjkRctydsLLDToGMShKWo2DyHH8jF2669ETC
37KTsSBMFJKcDhMSPev8UQfuKVpl1+yreAYtMp3ZM3Ic0mrUip1Gq/AHgn72twYmjX8suDZqyPVW
DZzSQqxjqh3mXIsNFR3HihRQlRsOkPaTH2qnYQpWGsqQtoRGzNJOswyqlA6FM1q9jIwoXtWM0KYQ
2WvNcVySNnBiVoFOZPYliG8aK+ASa6N2Cp6WmSGlwEfsRC7csQS1slWFl1RgtkHjjALrSBrlZEHX
xjUmewVVYzzj3sI6UftgbGBvPA1iztz2ZSDYm6bcedlIFSWDdoprHLLuk8df9kV8esSnmITYIbpF
b/mUsbVFjQeZ2S6XIcl8RqXD+XUdDWKCQFJeAcywweWwIuLoPgkjA+rMTgIjtQEg1h8sAiRJFAxS
5AGsjKZrePM6MBaS75ZPtaCPdnX25tkSqOt6yTZxGmTJFiC/UKrh9K86ImlxmYO11LFPWt984CuB
5FmV7ejwo0OfjoWZYkRceeZjm3n5Ni2Bf00b3qcsTCP4M/3qKxT8sazMWizifgKTGAQD6Ktu7UWT
94KiZ4no0bHvuh5Ax2gR5vsrR7XZwehwp+X5jKCHOdM6X+cA656kc25q4f5KodV6zc5hl/jL5ILD
hCG7wEchATPQUUzfy6xUi7mSjYu4B6qoXooZ61HFqPCsEngUEkUQVwtlPYYZ0rFN0Z+AbSLfxZ5k
ZDL0Uo+qSrHqGGeASY4Kly8GnD0ghtGjwEW0LoN1wBTki/jFWpm5yOHR93h8L5y8yr9TkNj+GNqY
ATo91d26Ts7GtPcetZysWP1p7XxYXUH3i0H19ihh7EmqlqOTVbpLTQWEFr4nMElHhdgGKFmI/bq4
Al48iiuLVxNurcwSqh+OWROHMD4/gCNIJwGevQKQrRY9XorRGd1+L/k1WwRSiBgMrGF4GXArUfAT
Zo+VsYypDPXnp8bOmqMdQRE5h0AXApSYqYPCanSa9O+KR+xDECUBwoN6M09w+qUQIizMCyBTQSmh
MpildJhQgANRl954KV/U2eZHm/YZsuzTEl7pB74O51etsMVeFp5cp8W/W6Z3L6oFK8hJuBkQXHfQ
Ok2mYBAJyFs+0B56R5bbf/CWDOBirab6NHEGSOLJJCZ9fUW49Xmg81h/02hvxiNa5ZXFRfe9ze+f
XbTf3oxaPc7FzwKSjf6ZvTWAFL2ve5nVRQPP0rFgI20ok+RBhWJQphrgWjfW50jtF6Stc0dgprnV
rEZWO9r93WqLYXyDpKJV10bEuxaTrpD9KrtbaxPah5byV/FV1mF9Ukcloc3asiTRuODfBl28RRw1
fr918VHnDlDTXeUkDHqxGQeOkDNZR1Os4y1N2jHVLHDMy6grgDTx2fGfKKhWBa+/IZIpGjwrTFS0
whyLwxdpdrWao9FCWQsrkkZhM4o0u7HsU11HaIzeySGRrp66cQFzcVTquMYPKBcRRdtxhLjDHDLR
ah5Z4+aodvw1NU7Tp2XyZzz8Iwiy1+n8OdA1T1CLWEe6G8TjdICzm2pd5QQqSt5IYzeXgJu4uvqv
Gryk48/mLvknsEepWvDHH0OyIiayddltMrcBoy/ZKmro0mL5BZvGbFDpo2HMa5cH834NC2wpZOaD
2uuw4CIoNo1XzueLtmK8SOlM7mv2etp7qQSe63YbdAnFCfHkKcscqBy7HJZL91hGS1CvHwbXkdkX
4UAFHn64TEkoF7rHpH1O3/NWlHqCf0kbwmQTyY39n2hzWMBUcHEnKZKvgUGfunt4AaKw93kAWqMz
7xRFVoU+be55jsoeLkpQF7KRC9kb9xps1A5mfkwTnvWs5mIaCwbBSOebBGx6arUZYc4J9ZLmrV7y
QspTdYh/EV2xojpb93ukX9SiWEeU9in6nrCaoaiznPsKuuXJi+GX1yKDWD89NHuY4Uw4oswMFqlD
Jc0EQmrZvl4DqtGsqDNkrl/Y3DV9Ye8eqXLlqxqJJQ/08AnATwuY72V0Jk/v4iYX5EMFEIWsl1Vh
ArVp+UB+Z0+nyvzwtxfsFZ3NydyV3OLQQDYweGwtpsAOMKOl+K40gFGFKk6TO1TdeClT9/gk0q+e
X9rgfsPP/5cyOC6e2RyZXUvopGJSDPSK6VnTImUw+lsKYEWBFKVyTedf53uoGfyAhwPfHwKemsRU
WM+0r9ntsWHya1tvAvJC65U/ieCmpDufuk4w7uliT8UL6hzASRHXfebbOBo15zEoesxGHuNOHpMM
x8XNBhW+Kf/p5LYAT+2v0dcRzWZHyrXnmPPTCcWlNKuyTb9ZxkQTtf7IluPEvmw+jtKMvyfOZlIL
grgNqiS3gpCQvzcTgps3OtR2BY/vSS6nZ9jkL54el/2zBc/uiURBTv87eZu6/fUb3qREINlhj03r
iiYvaJqfLgAkJsdXmtDBzJjzFrMb7WBN3KYgkTMFIfJuhQeXTgUPjlcYlzFipsQugB6LmEENEnmF
NlDBNVYSvE9A1wiysEpPDcwZcoZPIXn5AbAeZeiAoTQLAuhtTCbFnbuMfrxBsvkObSdi3FGg0H/c
Ng2cganz0XiUU1XQbl/R9/XO3+xbksb/0XBGAWKswYmiZakfU9WQtP2JJK9BeKY3RQp+2KUXiFHp
wasEBvMpHusJDObSJ+XRcHMGj8FWWnZe55HA08y9qBQFqIdDn5BhqKsRWfRVOmNd4uUOC/hMxrrF
n8kJpTyndAJ7o8X8zcSpp2YqI3KT8WpGhtdLAoPpjKQf2dGfCyMWjZ9FuwgNuL5T6m1X95MHkaHf
4t0Tyc7kKTiW6x6zk/f4/+H4a8QF2tDab2Ugje/OAv/10VqAbXdqPSogSxuNAxsRqDSbOYvX7J3n
zjcPwE5Ix9DPC8x6dpEKt/jtS8m9JmhstJt9sCIDzkW6dwKWuB5qI6YIzX12cef3BuCcKnMl2klp
wYba5UjeJxsElPoFeZnm5PXkh/SxlG+wZgkuGs3h6NOo3/6TK8Ysx6becI5ajx3DuIkfQNhd2wXf
LHznTkGnqICUSL+iXf5uTy3hfkTRWBcizCZMRDp/4plh/7cfhfoF3fpdTkcMX+M3IbKefDIUlSiN
2frnANHPcENsoue7WYPyNq5SuytkZKT2XY2FBrVr0urWEjW3T7S8lsbXygIB/9w70FWM0Q6PiWoH
k/9dHwQVwEh4jpaXJYK16f1Q90e+FdeTUeO2YVLK20B0BXqSONJIE1oG2r29rFOSbQGA9sifwOqi
Ue8/1L2bTvRgtyEy2DZK4jPXooQ3/Eo3KxMqrzd6ugFYs+wGeDF3zza/apyCa5NczsulMFZ0mxne
4oi2Dabqwuo1SxvGUMhAyBY3wiMwHwbG9lKV8A1Wf0pB0JMUSL6DEby237bWBU50ii2J1CP2n0JQ
SNNP4bGF32bSUFPcgmHPyCWT3QFwXp56f9jbKg/DowStsY/OLC3yQXjNPJ8B08wgzYQjPWMsqxIj
fimm7fxT1Gvpj91P4B5FjnUIMPZIwdMJTU5H2l4L/iM6k6S5OAfechu5WJlVjHIn3NgPu4a7vMO3
Y0S03m8BOJHeL8d/hikVMsk97bHbMGYm5TdQkOWleR0vAF7oEPIyBGqE4jb7q3wFmWgtqSYixUdx
DhbU3eJ20+D4uKY72ZEKSWwt4LS/uA5H3+VQe1z72+qZgK6LEOyp/vAHMLYKF9lUvB6qSirSIjaa
MniIxPNqK2707nUL4uzixPvgeR1wgdLll93TftWH2LStWCgcF9PQt7kTkC+Vm5+dvIjHQhcg1ikd
N5fTYKHToRejvrc7Jd+80VF+AiLe1rg5uwjZ6zGZpS8IG9ZdqhJejDTk7x7js0OahbDDbG7qxs44
Yh4soVdWPL18IMrz1qBikOKqXBw9BfMuJF9+m9BEt7dxPJMowBA5QhiZyL2E7C+PjkFIBUdB/jNb
a/QEhLiyG5Mfrr46jO3FDPo9bQDlLXPHT4V93Z0IoeWs2S1rbconJZIMvgFqmZ1gwsc8UFPcbyuD
SKDp8gnKRYGLnTXCTNcmaSKUFEEApNuqlCidRdpBw37fcIwynC36QrHZ2SdW3OPmuoa3gErXFccQ
rTajiHYkVcp1fzA0z2kMHXmT+wZs7R4QhUopekohPZ/RiTWLhhzQilH+fEpUfKW8FjxKXar9QkFO
36yF6i9xAiJtzN6dR+hOSXyYduXB3Dh2iF4q29r1xv63FDbMvzNqzIuilL2yOj4p/HyR2dVqv1gm
o8mJty5eOZm/CZZA1olcRE2ndzO6GE/Lt4dBYr1yeGZSnqM8QteSyIF2I7gxDwpw58U7dhL1uBoe
bEZmThoYbeGdaBOTMbsgKMBZdF/fiGXJeXHbDcxoToigZ+LjqPVcw75FIAaON+QazXTPgqI3LyJ9
i7LIr7nhFkTahkGAUEwSYst7nGdrBu+wRQ2Gz0AyWBtHLbYg8IhAaEPsEL/RVqn1p2oqXPEBMd/F
9Scdsr1K+YtNb3IDg5SWteEPzIfgUp8wqO4KX/tcrDPKROjBhrq0KgcvUUe5RYQmY+EtitjHuVju
byJF93LUYH/wLV9BjrCaoj7jCXldLbpM1Wm+L6sOOgGx9DKqb2z2OWXmwBYZVB21WnKiwh0dduf7
XgyTJixpRNHo9KqG6FKadkLo0m8siJppjvp7V9WgNvxbCzd5iV7O0zfKDT16PJL8vtEbQUhQAFSf
E7ZGaAhmn7+Ubju5Eu+RZmBERbzBDpqsV9Nv40eVs01GJVAdtdKwQ/Jsc+pJJuUve+8OHHQAtLkB
JwBrtmK/Dy3Sd6FdqXPYhCW0u30hezXktKhTnFIZvmR0fbu6AFCcpjcee2I1fZdFPdDEMP4XD0S7
zeUzsnK7mQ2TgSN+5e38ZFXQQEwFb4ujbj1V8od9lBf0M9d/yuZmsutqo0CE6Mhh4204acrbfUgQ
TVqSsDRb+Hh1sSfgzNBRroHP/MWlbaPV4gzAxOmQsVUBSVu5JMLSs5lImmHAmPnebB90HaCx8qvj
Ncku1X/a1rcfEu3oCObWndKlA8+3EKJo9N5z5H84Zw0Twe7PZtUJXIdw6/dctSkvfPZMmsVeGtrA
gcISOIC+54to6H3qe1RDVZfUQCzqiBWB1vU+fdyRGg/vzmXYz8q7UeADVP0Jh73lZiDzmk6uSaFo
4JZBHtwR8wjvPO7t6U5QExehtPLcq18vS2gvKvJ74/MVEonAqVZYT2c57UQLd5JeKf8hMQtjtOW0
UREGykNSfXwvGVRoVO8hCQmN4wNkAEVVR5V/1Shd3eh2zsATsIXDLq8PkSIxLpgXFu7o0N5666/N
DYxJI9YCE62C7EGm9MjySPvFoXd0X1gc/Al9aj/2DA4Ups7CGZquBl3eA0/muqvMiL54/ugsXsCC
I1+619lzg8gY2LBXfeFIAExpd9DEYqw8e8GnDXmXlLffNlAZTlQE9BOGXInlFzU4CskYCcCKz43E
BLTNVVbWdZ6JywRKmgi+bpl27lQrnEJg7+zX9Mm3vvwmnPKz/lzpXryGOkoLETSSco8m3dVdEOEu
cIDI2JQ24iZRYD30KdeGyRd34Pgc/pXUCtOa5+4hEpKpx19+DLiM5cRbiHTesJ/w98efnVTRTfIT
TFIIY/APhXHqyaqSLqOnuL2GjZzU0Y47sUpL+BR0wXHAeJOn92CWBKnLitSr6Vv2VRA96gBVBTH4
Zej3L48aSc7FjCJKt/8Vbggj3rrRIVHVis7e4C80uPqkNoRNq48ZL6kD5NC70DKEL5vmyGQ+gVRR
IlwmpRqpOevXG4Cke/s+x7pm1PoObQOROKs7REwLPENMQnDaiVX5zmuCwl9oaKJBZ06XhsbDHCdJ
0JNu/XU9EWOzv5DtFXP/1ok+KQ2lAGl92i25qiKOOMcOaq2pCxI9OEFeS/ItuOi5TqHxQZCb4WDw
XCa8P1YTcr2uAU9ne6d8pvcnF4CNikS8mIHc7efCnNzjlRko1pSec96IBvC464TRyZeGBn2eQqXk
zgOuFiAbbU9oBdefRvTK3AZa3OFt8B7r4ULnI6lR69c5viGS6+KsJ95URhy2+UU8N3o6jOlorZ/e
9WFd1vzHA2tLQFmfNvzqImGwVogPHv68S32rIN/8V0dBfQMbH3KK2QVLYXdv3SLINtVmHPjVqyvB
IZcy5DT8uYtc+46MMud7E62DquSWwU3tLyj6Xz6CADkBXtn2NajkY+Gx9HT1+D/byeuYMJThRH5w
Sg/qdZaQq1G4uH0vb8xyTwcU0IUGAAjCWOv8wxhyRlygaHsfS4ez8OUrk99KgxYT4XUK5SjwaU2i
ZmJMCyFXqky/Xu68n+E8O1P0jDFoMm1CIcjB+yExT4Wpfoc4EiaHvHUmzxpWWVJgfUEEIaW97lJA
UcxbkuOKljICYuq+d1ntKVA5NYkZ+Tr3UuTFI8WZ7FZCwN1zEzUrBfPVnuzwaUXob170hIRSzTOm
nY5vaVwRaPZctnrSiYReFhb5jYkwBlTQ18ivYGwlbe3w+5mIr1fl3ruQ+mtVqi5Qk1fH3qRLlpOj
XnLodrjmwcPBA4LvuKqHo+j7ruJ17jeYF2bRLGkKjlc1Y8IK2crho9uQfzp+7YbkxWD3pjknN7Ob
iae3AywH9/4b9RIL9hI5CjXmWBY9uiPBDfzuGdmHFE86xxDwrfMh5mipe55VeVs3x9QiKrM/ndwq
5S0STSiqPpRH/0B8oKhCstf76SqUlPn4XRS6m+yxra+ADwiXfnwstPHoewp6/juuBiFRjq8JhcRG
Uzf3J61w7wXeypG8jtKwDnYFba/4ClHa80D1HMVfVL+Vp55UWiYnVQml8PpbtJ9SUkXJWzSFF3WQ
v2L1DxyoTRXgtlJscUz3bomuHvhvBBwQsDEG0JfRPchFEsvteAbQuV00YjHAk3FFVY2C/hFrZn5x
GUhE+q6CLxMDUzb/1u+Rs+vHrxawjbZ45zYb+y2KCfOmntTdo05rW90Nt/hFPa8endgCquvDMmqy
b37b97TmE2qP52gJ2a1XWoZYWbPOeLi77RzR8hf845VBa0tC72ZLLm5ByZ3c4Rg6O1EYXDfSlo+Y
ytXGkx8eKVXs7Xf4HXg2A7yd/q33cfFDM04V/wmRLZqL2YWVHu98UjXAntOcXMSDMX7+xRabbtBg
+7jRrXKjgto7VseO9TTfxsIPrxXAyBZ4VEAOOw31rd/wlIRkArV/sy4UcwPZVJv1qgtjGaNTFagK
ynQ+9fJcIm2SBkirgCQtmrGvBZGEc5WEJnceE9ixUlvj5aIB3UjWBhKIM9urbVZhlS1EkiVGQpbD
OZ3AszEcaT64hRpqm6vCd6EXGPrJOyszJ513UUxlqVVR71vIzTDGC+Dekx2AEw81w+EdC4i2yXKO
s3QO9oCDybJ6/Yq8EZwqG134IihItuXR9UnnZHOA3LkRKH/zD/7CZu2VsZGaLBmM2Z8nEjTyKA6r
jsWPFYMubqg7k9wC7R+7GIfWDdC7HAuJ6+6pWA9a5Mx4L7jHSss5Io0+YMgTGiRVxPK3VUdvJnfj
eFNN3oZr8sd/Nt4chXavoqRukRbFSfRvCUkneNbSgG4CaVFQgnlTV2uXbqJg2YfD6TyS+2ge/0w4
BfgE59ujdWQm8HhJYrVTWbYMYJE8txo3X69L0gcy5NZJSmyVjn5rY+I2lXDN8xBWFBKYjGMTDGgW
RfqaZoAKZGYOy8uLp02D6KnuNW6ooeMlGlP9uopDLMv6t0+W3XVzGFP0GrDHzRi0WQa98J6KdS3n
5C1OpdhEKnwUa3CnX7jKrIKIqq0GQgnzPO/mTsz1zm5dHDriyfeO/ID9c5Pm54D3+IVPDmtzwlbv
uDx04BIR8KDz4xnfb3sS3JOUtgQekKRfSbV5jaGYRH2ssbjJo1MK0a3rYyjEZdmYQzzwN6c+Dssp
RXl4wEgZpAjjkd6zzofInEGSExlsyPBZ0HJlRdsUILKolPhc4iHof6XIgHBZFCR9nSgP5oefkPCS
lt+cISPsbB3ljhx0J1bSRhLRJ8CCVSBu7m6YtPykQ/5stiOONCDQrFnftVvnMhd9qgAYCBoHTzso
UNMnOd8usoiUDOc4S772lDfOYcOPS0UTWY8YiMbWOkpJynJ56wvmg+mHkGSgSKIxh33ZzWckptUE
IaSqG+KLYJtWatDePY99PWc6I9kmq/wT/lHvyU6GqbYtOgptYEpzuXshco3hcYYy7N6dzN4MBXII
tSJDS+9jgbth1b6J3u5vVuod5cgc8/ho4OpqQKp13XGJ5e958DcDDTWgCx0ZHnDg2bji9MIY1rgu
kEyccTRirLbh/yRIWREOsK4ZSSxdEaA/DkQArLdrtI8u81Pz4DgU+HA1Vo7H8sPzpuGjsZijnTaW
nkjBhsch+Lp7NBg9uS/iVXyqGsTHny1aYt3A8XLoFXInwfFmSYZ6a5gY1e3j3Qhg+ZdhaUXfZ2T7
px/hI72/ns/BkIp+/4+rS5RKqLqlJ9VpGMlEG5WyaQNm00r4hRxqGMQISXjRb0n0bHsFy2EoOwJj
TWHmMEz99GbUiGEedaMLIAJMzgkQxyQUScBTN1dQykJi+Tt/a756fEfliHGEu/s/g0vuhr9BpDRv
nzo0h8yqxVV9kizrTOtN9FybCDfq0bYvdcayKhwaseFyW9Al9lErguNyRdTeDLhQE66jjUJrwLXB
5w4C/Bm3Izb1+Ht3N590BOeq0XEBacsOgR4H4krx3XJ4LeD6AguNaoaHgeinSjSGBletL/EWcphH
TaTSTGQ/W5w+AEy38PAhilXsRUHt3+fnSfhYLGYz+enrYyn8whFBEgg+mqyHu0t/T6/KtARje9Zt
EADDRzLmutynW9i94cM9jY8k8IFHSqcXggn684WD+U/FMJ7O5wKftF1z2jOVFXXbis/iYUF+EnG1
LQMfBd7i8Eus4vo8PJgGDJuVI/q2+wngphfyqSYrCDZlxzGNjnbftxNIhAWKnFsIvB2twcy1+J6G
EGqE1LwCz1+fOrDjROHxnyEDBZ6Ykncf6W8HGIAx9trUb6tGUFVZ60W1GVbrPncacnwtsgjm+odf
uSxiZEbe8AZpYSbSNcD0vgpWzwAtM0RNrRlOGjRMYB9RY0v4q+W5a7oqovjlMv8tgPkf3KmX1Ms9
LtLyca0NssjUNTksgQBG+YUfy4viv1FQVZZn1c7QanojNTo4WeCAXkDUstGdEno6yefn4bL0X124
MTxSSpxMiQ5r58rw1mLWBrpsr+mPp3Ak5XbnmhD2GJxZnAb1OorAjASjJEyl5bC3WVx2LFsxMSw5
nNd3+4gdq5YdZANYaeHt5mnPcEQ1yp1M9/6X1Ri8ySS6RpN+lMrZOEaLU8pu0FiElBNKlmEBTzT/
y5IJYZSQrX97js/NcKCJ79RWLrWnQVoaQzRR+oA6WTgjkORxLbpuqBmVW3P7iaoc4nwU0T4IYFHo
wEe8RhHX2E9h+Kjve7puTBJWZ3qF1yGOooKeghMjcxWMq8WYh1Jz/CUOzWm2MfnaRwSJ07QkjGds
c51H7R9JrLUcqy/7bGjgYSy6Sv/MloNW7QpLd/oraWnwmCZrrTVGH6D1W5esaYfTO5idT5z6XrAy
bBkjOytiY6gDtQ4ULz/GHH+znyqXg5yH3Pqbh5MBXn7t9ZP5l8XA82GlbsHchthTwoSRqunCLeYD
XqVyaCX5P9jvn9QdfsflT5Q4qOJg2KCDHXCReBTFErzqrM+5ZcRBM0Hn7BjfegN0ejpW0t6/VOWC
GrPYIsi3qbebigBbTCXzU+8AxLeRbDjj3F3LpGIcZ2qI3cHvrH2uoVwef/1pWV4aywMhxzAWsy5s
UfwAZkL38VULuDkijUWJCcJuAgn5ARKOHBLm69UnWvORPafeferW26rlijCckW4enAx5Zh2lUCOM
E6CZn5FeWQM4lfFiPZfyhNiEgcSyk3HzlV3z2LAEAdzKmj/UNnf9NGbxHpuCrrcsH/thOqP61NVG
6S+GuFXgAcDauZeHOv8xhcSJmya5+KKIKoIG3m17NhsdE/nRXcy2Py0MUu2v2azP9xQgTMmwvhRe
hxcS04ZKQ92hRbcQCXEmYjooWhYqdVNJtvuYtNVA6wkF+yxrSZT5bqrg37K5lZzDYGF5nUzqv/dL
mnjId9Gy9NF1NOfIUg31lQTnOMwV9uF/1yGrcloYFg/lboxD9EXInKCKyUcVfuSf7jHAGz8nmyjm
Vh/diulwl9vXCN3o5CVctOK8GFBdqK+GVtXtfNdHqcyPbekL2jUuYZSYU9eC9JqP1KDdgwWkVCya
/WOvlj7XzEVeLfx68WILIWnbT6BiDLQjdVsDLOa4o7v+IPzZgJB5L4z/WfMG2hNEc/7QCcYiNqzI
f1+RyWcNK75jwDoytz0L9nusQvCzV25LHh9HOcYaQI1L4MT9YuIoeQEQaP+MB1ORRCn2dnZvm4zU
sYJ+/BasXI5aq+JJQ4P+b28R3uaD07f01uqOgdk9jna/ThAWvBjkKhzupbCSX7WTgheE3nZgaLtR
nnkEadjoqwgr/2dVZn08LXD/033LRKeVTMzMKZivrwDU08SHZuilFBER3xcKKJmb2xBfr5eewGIL
mFI3FUN9jelislRWPBVWTbM4e9i6+qqdnQXc3a3mYa2WOIBoRToxSdo6n5qrZQPc9WvlN7p+k9F6
eQrZY9abn1i2ZkHpB8QVH2R/YxZ7eiUkvuQdOmeC5RLUlfq+KtbUSbl+bjAHc5SqtUJKf1slupBk
3QvIIttp2Ladnc5v/IcbsxCv1GPyCSDSFUjqRCVUedA7c5Y3VcAdDJbcGvSrvXjxhZ0V0bCN5JH5
AcRDlPvUQdmXUoYeomBT3hLEukXj6xpWpfYPWEY2MQza58+twsF3dkBZ4sqodVWZKzMeWerf/z6X
Mkhggg7OC1iv0t8phltIba0tl3GZ4iSXDYXLeWK10QC0JjyCXEn1TWRywY8w5fxF/d+Pkuvgp69m
SJC5sfppaipYASp5UNqfI0cB40REc+WkRkyTwh6XJqR3DWCl8BHXtEhc/Il9HmVzzh0t8pFRUiXM
/C2xNpZgGCU3FVFXeC8Sv74BNR1xb5t4xkcllbBprxD/knjeFwxDOmOstLsqwjUnh029PNGIRixJ
/I9FIKBOcW+gkgADAF+qkDdgBnq/zoIKl0G8LnMImNpUZPr0Huq7d+UL7HPwWUhmbesVWV4ZjBxE
Iaz5Pt1BOtOClVWKwU9A5y+ZwXm/k1WEBC1YIXw96UNTeQ4yKJdEMbeOMKElyIXxTnoIdWn4cApT
lEcmPo8d3Z/6U9evKi7efzWwhEqA+owVdQ2hcpmIE8nYOLd/GGU5UsKRqhG8lbX0EFHD3h3BrFQP
bF5knobCViQKmjwwqy7Y0XfSojuobFFI+MUFONSs24x0Y7VU8wGzRCWdEq+eKWqmpE6lclnhQIq+
iSQSIx561O5mo2Jbc8QDV08evszwhbgqU7uU44jANVo8+rw0Vrtfg76DSo7Mjc6c60Kg2MJeMk0C
J1QtsUJoAfL0DQmsRulPlrHZaSmGTolHlNO5+mHobW3rskAB0RbCdV0OhQ1F1y6jTGhYLlEJgJOn
cAxPbq02ASdvA9Vi5PnjAGcdEVIsVVAcLZdeqYJ3mqNReU5QRdW02CVyGFdREqc48+Jy+KlOURuC
G66374gMPbymx9oIv7zrScY3JZtYsorm7JNpHJ9YxtLsw5iLdz847t1aswbXg8Lb2RSQpY3d7nJw
ZzkiAnknEaB2e0W6MdXbiNrQfyv1XV8AggEsxDX66lae2+UmAT+6PJE1uE0abeT+ris3kJmUCgdd
d2GLC0cGY6jBOYyyf020F+RAnNq+YM6wMS7ihDUO8S9B3ISei4YmGwq2SJfMrw2+N4JAb8IIP9AK
ncNVQeoKMGD37+Wv1MTBSgd5S1shXblZIkaDm6bec5zJ9QlVfe3hKvKdN5dDyL7x7FJKiKFTvnvw
zIFt0F1YsEA4VPxbcDXdD8ifCzvXbEH61+gbBvGNHfenXjb+yPbnGNefXo8l7UpYy8MSU2ZH43Rr
d1ZxeQpzlvCFDfYbN/rzjml9UvXNMe+rbHR8+sCj2OqE1CFskmCR48HSBg6UKLf5SBrdh4tEsdEn
H5kUfxQEaVVyeg6xMbnpZbD8coi8DhKQN8vBAue5fdWVlOLZJS4b7BS8CrnWauhKsQJVNTZ9ajP/
KbIn3j+YC78YOBBlWNZ+DkSybrE3ZbSaPuKS80uJF9SwBG7rGZSp3tjX6oJ1lsobM02oztOaI9J7
gsNuX0iGyjE3X9SIfubDye4eqq7coGiE84u4bYso4HNSWg9eA4IOStZ+hVNcaMVpsJkBL4Z8wDxR
9GmiJozPJdaItF+nAm3zC86kuZuOZJSOmWeSzVMkpa0v2DvWzLgmJAQyVVBUk0DcTIy3Z/AkOvYS
81bposvzaqZylKlnqMXDb1BoifgTIKEtYLUTc4YR7fI+uRqP7LJxsKRTiqD8RaByzmFTrIz+LwVN
kSSNaoJTPEFhnirU4O4n25FuKnKrq9+XHZPrEjo6qC2mQ6tE7SiH1cpNH4Y/XoJ9yfOkKxyyd3Js
iu8uDn6LMFRUF8Yh87gFd1p83sYD2pjlkNTR00G0tyLCUr3awYRToayld1JGnSip1R/Dd2nLHwOB
vzXlu3LkPdCOlTsmekDo5/HYzWvvKRtDdEJdrZfm4JSyxH7uY1HV6iZb0YRth8kODI4Uau2gbz/i
uj4w41qly9S7REAJiNUCQQPJUy3uwuMpr3Tk6a+DMvVCYePfJ1zrwD8CjZRO6KSP3k7bcTqx/ASr
oFFZVEnihOXhb0FxnQv1XoVaa8Jn+gbvsqccfzQLCkYk3L+1m76XFE3yHKdNtgWEHNMBCE4UI3yH
ecRfjfSzAbPDJop4KSDEgrzvGXdECIZ4wHhVs7jggo/5oP+BMFExsdJsQv2XOKv02w3aF5QreZDi
OIoXt/UVg4Vi5QtYOiF8oV/VsBy5myc0yZ9Upyfu07YnbHSSerVrDr8F1gOeGPjUuzq0ny4tqlHM
d5LUrC/MbTCYDMC9zd/ScC6On0OehLT1tZyDtRTmzJr0OseI0wg04snNaGoQvrUSMiyoJlVAIyAa
36UB/X1RTqhEUA96if1MXFVf2NkK2Laly6w5RGwtGOY3JJiPKA1A5plNeAuLArIz/eNWi9AUSyqg
IiWxGxbzH7HoLh996q+3xThVDMV5O4tQKEdVPdDjpluXvC60d4OYf7GW8RvO/Wo7McrExsg+o6S7
Iyjv0kWI8BpC1Nmvm0g+y07ZaKuYylY5vxGFyPBNGEGU/GkH2eakqRLcg5Ov7XaM4v9ke4T6odtj
4nlue1meT4GQGtY3w4uLZLgnyj0NMs3exX93zDhJpTrkw21JXClnq5+I0+EroKrxe+q76rSJy1DZ
y+YUJxW8cqrmaafJl2nLVpTGHyv934lmsO5ZPa2uNOBmbaiwPCJcPskx4s1rK0L0arN27au/Je1a
Hu9UXbz23bpXT/hfP58pE+krxTLPGz7HbHI6FBYMXmosddi/wojfrzhU9Kt9AwIhcFI1awk0HXFQ
keTNt5BH9A4KQKW3fLQn1zbovGMCDrcSaZoGNvozs5FQkqCD8TcWSDE/BXTnFi6F8fuvOax1vc23
8Kp4hmnreX4b/RWIiJiJcPS8YcWanbWt/hem9MZn7yS+kAQqZy9aqbKbaF78TL0gPzQk6M27kSRh
QcWqEy2GNQJBJPpEb+yxKCC0TEY89imzJANC0Q3XdHa77Kg+7LJ66MIGKsaNaadzwSod0mY5hU4h
k1Fqjfow5HT2BgogtcxYT0wLr0AoDTnJ9gjrAQITyCfckxkXX9ktBhMrWJjJRDmRYP9INWU+MbH3
J6wDd1pnoE7Pqu61TukhbZZaSiORs8PTVts//G9IQFE117qRlw4zvY5CY9ILirr6hIRUSukmO0we
H3KNW5O/yXQhSSGTGfvy+DkDMUorrqXWPCyu1oIIa1rHYXLZG98TOUjcmwFa4gXQlrS43z2LJRGU
+0D7Y3p1zIrkKLcKaS7auYZGdtiUMF6wLti3OjfBeSurBsksNYgjMLIGLJfii/3lt/JcZKDSTUOT
bv9gu1EvKP6p7Z1V1ZaLoAmHSDjpbmsvvMB/GgaE9Mqpg2SkrTMXqrcSExZKysdBnyoFuhKBKBHP
pAVhRythKT30Wmwi6j2mD8Q1OD439ozPcAIMdv3aGE2ouCqxDv85iuq8/EMOpkPRLlIARLdP1mo8
fqbR5oB9CCgRNkqjtcyUmikUb4pXjbf0W0vR745PmbLSGgFqIf8UJkkPgH2K05A4HL18pkNdSi4B
eBK4DqvOUJQ9dw0205le25n+/xnH4pvjLsBwRk9S+pMNi7TUTMLoC0l+SuWpQDJTXlNyMA2Q/JzR
rW/wk6cp7kIjG9Kr8ww+JLeW/TozDC3NRsWYqjsSmA6VVziF3zZspecluJ/k0D5O5iExRIzyAUGx
clXZZQmRlfDY6rcuUgkmjL/RNdVZE1SnI3DM59wUf3n811G0ZwqJtdAg0zZ6TjaCFfwVtAKFb2gJ
Y4rsgLcYBvlsx5Wyu5Ei4dC3msxcbK8nQaXd7Usd8aFRV6XClEPX3fuGc4Kj+ILR8cioSgZgR0+q
y2hJdwsCpq/FRMmsUQX9SRoh+enuOVz8S21R+6Kb5UwbkTcWJkFzQuX2cjRkM3b3Eh3Rj7yxTPbE
UWC2TETtMgpM8+8HCsIIbP7ib5Uj9py0rhlk8Kurb60lLiWaGdN18NZ19MDnvTQBqpm7v/udxD01
KN8TJa4q2gshcarhxlwGSiJooJmfe1GnP6Q4t63+kO1vf1566GmwZhXjceXjT9PS2uYP2ZTlyQp7
MCMAK4HgC1qAIJJsiZHVT7Q95tfnnVUf60qGrkWhheR8oXWYA5YXcwDsb5UJGOtQYvWymSN9lvUa
ybosn8lNVm2GJBkhw0dj9uEOO4vo02wjmxYutMrXccVVTfaFQ17KPgJLWmWP2OyfD2HpAolcMFqS
ylt8MtxVdAFVdATpqDl0nqZ9Y3Vp6lxLwEOKcM5c94SG93wSD7oqpV/nx2IB0xXAcnpaegi0xAlD
jL/YyDUwvNqHHjqLwBwxBFIulgSFwMIULjNN56/L1oPX3rxp2xpG7Iz1InOp/GsmqRnY0IL3hCP5
CJeDgIAXmsxdbSao6+0VYB10mH/PWpTy3wRRpyPXQrE9Ki5S8EQ5F2f3WjxnCbeKobyc/woQej3P
0uZTocudTTDCanC7qAf3S5gmSwWQ5/j0jG1FzCgRrf5EkAB6X7Gfq+khJHxrI+qdADNYGWSyrZiB
YtJYhUHLWqLUSsR5KW/0loZKjAizMPuZQmLF6/A+jE5ieEYPiO5IiFnmTKblioLJiVtzNieDy3CO
V0wLmfweygrph9Ysvd47AI2uxT/wZW59Mr+Gi6QmS0J2hsE22I6bM4bkRrazDU9TeGSMEH2D+68U
iRMj6fT+fm9p79Nob2HNHOUTE3R89G7489tbcUCSc04LM2gAwJipwBYiD7d5jHvmqEwtbNc0N59U
3ZNZSR3pQkuIBTxy+oUUxZr386aEY791EIe+8UfDLh4wwivRZ10YbmXpalhI34MqnlT1MQT+Uwb1
0kpZg2U54CkQYdVufJQabmUPrsF7zscDflFg/6gJxVyu/pttHtO1Z8sA+Y7AoB4/mJJev5Sxm1Lz
da83vtZJbWn9cAfKX0mkVPPR2no4v3ndxA6r7Qw0DG+Ua5B84cTsHe0880Jm0jmPxz5I2/DTSnUS
MQkuPpivBwP0oFJjBdLqIv4YyT3gVYRwLQKYDUfdvKkBlhGHmwIHQzOQT735tgR4YevF1ryH3tM3
WmWQpRttfXpDfHh+8no919BQP8zwD3Rdjk2xM443yMSF6vss2D+/I/DOVfGJkUItD2LopRN7ZJQd
9fK7QhHMdfOl1Dd9JqB1sKVBJ4A4esb4Kwt5Jv7yFVImJ5e65d31XHMXzpoAIO13WrTLUwvgAx+3
uNj2e+3JOOp+Si3sySlu1Nqe98JOJlL7W1JabeBIVobCO1riLgp4aBJl+J8VGpYxmXeYoYpUp7Or
zpOHvsfpjfn7fDqqTuuXx1IGzU8JWTqBBUOJAvwCKfdwtep3kwkB8G83b+jSMrAOvAHjoUJfFwka
2FaaZOsn9meIvONg6D1JKaXXL1Qkm1bCtGjuU8sH2vztvYHvATfSTofIdKb7tEzwVD0IYxLeAqyl
L1eNri0Gglq8iB2+H/ioWSc/tipj7MBVashtquN5QsC/TsAyY1o1QSTH8cIR+wSc+5jfiMv9Uoqn
ORcrbPqjOYAm/AHEoA6b2vMiTmEfjefRlXO0LBRc/4e70JpKxV3wfhwsKGLcprSuVt8aevccV8fV
sZGjSCMq/pyiNe0k8NQKaLtoYufvrPrxDEd3oWz5EKF7ipD6znI+tDZGp+2u34C6fAJBrDofmzaj
Ou7iTsydwHVwcQazxVijyYZuLSnQMhJn+gNqvRzMVcrW3TTLLaFoDADZ0fBx/l5xGhwHjTN6Vzgq
eFsFxrfZe8xa5VEUiC8dD7bBFK0wVizgR06wQuyQoAs4cChULQ5PNVcg+pfxBwmgVKyIT/9C8/xG
8RgIOtgUxnxRm7R0kKQmZzUqmTwjmtpbqCh+a6ZOKvfX3XuhUHhC4DEe10IatU3tZ5neDI2f5o70
uRN0pYJCn9BqWxIV0+HCZqW5CHH+MQy7Hhcg/dNBIcXK9qY3mqHTq4xJ2dG2EXixrLP7TM9aXsWu
MVVRiAEX/4g/7FM2rG519hSMeicBLuBEqdmQobwdGcKUn3e9wwu+bDEoQ+65+BoEN37TkOdHulsU
FlIETJVJbNKcg7VKFcgWuVFbEL9i1ArrIfeynsVhdsrxVhqMkkSjmuSBJ+jezb4PJy+5R2H2+viK
gBhvqfo/QIcTQsD5Tv7eOzDM0LMhMQ1aVBfCHRcQuuc5+soSkpeJDokKqd08H+M/+byG4zx74TtS
Ew/V/skj0eQYYvlxnrJcVhcDZmyFVBArjNaSvWhqKmSE5GoO0fEI3Tj27fkSL6DkO0vFkGiiJJ7x
R4RdiB4FZ7MzIu4xdHHLMorph/imf/8ebWRtzF1TOeQkIOVMySyoe3phZmYhflZe6DR7Bt4duyVz
eLhDKUcjqZ+ueN9Z3LIfDOqocOkzv2sf51xQbJa19igf0K5WdJLWkbiFYZyUCnkG4R0G1wa8IJFt
bWbSl//1tzLXFy7xHLThJT+H2PsMkaSLiZhxH9prGDOUGovRZTgNK0JufSjVdvznBYHcUXlAq01y
HKAY+jtNWytcaA+qNAo+2IvTNlZE98wPSM6vLRlysd5Vg0s4Y8ShlvbC8ZKVJztgf/FonTXpiyou
SmEcKBDspaVrAHIfyMoXjD7X8dXh7h/2MbSZ7vh35SIuMn8rDyth2eXJTw89aQg/YwVya4PYx4l0
Pr7BYYJmf3KIzdRt8/hlEOmxIfHbRlvk76hHMBOlHz2s7DP76fipDLSibSQ+DJMDwwqQryHt6sl2
o2cunwJLMpc+SKKQHy5xtcG77fZgKstGcFI2yX9VoJz91efTjD+Oo6mUudDw5Pb0rIjrzExJb9WX
vdm/EYolN8IjGhaBFzENgXaUQjiwHegJnO8lmZ0zrBXNmjbfucYMkzh1QtoSiFIYSzHEgNnDasRt
hDXNeCBzP4aRqjlCjfvw2TY9kNx0C+9+P0U6vvkQc2LvcvnY5rgr8xge4IbfQ/eDuN9NAON779V6
hJt93AQdi9KpGJWYgPSTDphFJHeJNiTqhXX7dcVVtjFmIkzn2UYbmX0ayTwmVmkPL+5AAy9vrwKC
ICZNa4lOiwRnRWZ8LGPsJzjaLJzk4RPK9gNMK24tEPx2ZARCcFZCVa15W5sHRMkFqCRfgRxn5d3Y
zAEIV/A5uxC56+xvYfMxX/Galgdx8MowZqkPc4/NT5rP1+56vsC0DuhRrwiZ37XWIpE+bBiETQhl
/kNrveL138qO9u8GScZEbanPtXHKImrUhnSXUDkLq3UdfeJIURBcOTf60rHIpno8JeL67BhYt8Ej
EfAALHZLHBa6H42xDKt1hlXNN1hp9F4aBigbO3XMW6zEN7yZRbUdTFXWJHRSS4jAtOdRGGDs7NwZ
LTo84yzhMRpaRduDau2s+Ck6hBAvgvcpf9rDqqwEavQY2e292dKt8GVLMn7r+Ja0z7NhrQVjDiBu
IUEezP3MyQU9LeKccWlmm04eUAc1pk/VnqM0Wv9rh4SxTQcwF/9mt24KHdDQTq0I0R6+0y7MKdCN
uGoiqU8nYLFZHi+ixdl8fIO2DPGKVPJ5ge2ZCXJ/Tzn3eyTJU+3Qajm9kKBOqptP3z7ugHlRwoWV
F7hSLEtaozIdP3bDbpO1/bH1gZv3z6eDeWbEvCeesdkZFRVy91nY3utjJLlN8IItt2im6sKgwMer
OemGhcSjTRoLkTSupnQsd1JgmLa73pAkQ7TltjGJElWkBxdll7UqwsjcSQhoacGnrVeGyZX8KNDc
LCbWWHbMspQuv7Ce2J0A+fIEzTCOQggV4B/+VY37KDJJlo5VZEbepAmw64yx1bsOzZvKsbRRFb5D
KQqXJECsU9o5yhlfO4GD0+PqXwlzOFx+R47QcNWCgLjoSig8LjGFXZlOn+xGGFXl3kdCt0aMYTHO
V5Ygqw20oWBZUOguL0/I6EKIdj52lAgAUW56Kx5MShjYY4ely2Fnp6oy2t5VpXBf56VAuUURMI4V
eVqDxYdRTwACer13PB+TJQnUr6d2HjqqFXc6l//4mqceNp8ysmSO8KJI3QyrXD+YB3h5sL39Zy3z
XEh+wiWMVqg5eMSIxfkgFCdqpsRUdxSIyc4fmXVBRrk54SnqC2lQ2z0WkKaXS/Q9gzIl3n7mPmo7
2/9hW4sOQ+znjzHIb8sTLeS6u+egYyphmdHGsKrbQe0MhheOwcNksmmOW+V79E5RsIrBETvK9Bz4
OzuoErnlnzcFRF8/NUaUozPNycN7NnXP1TjB+nfgsH2/NryjEAsf0IqX8EWYWC5qczXTeaFUdTwO
yzDeAgrcqXK9EMaq4oAUEgfU7kLyKlYguFeFyYsbmaum30A8pQkMI7Yr32D09bqy8BhvZOXxIBZY
xb2vEtKl+RjKAY07mQr/2OUkl90PHkLsc9KD2jCsmZxJq1IC3N5P6rrNnKgP3jnzkl54l3a2HE0N
+xD2udjEZH78x7O0TZZ0MMeZOwr1vE8vCZHTAVGtzu1wyikx0xCHLTVkmYWBiA+VAL2aTXK6ejQW
iTg7VoNQy7Aa607Fqt/xGNIvYBTsijQFTnxiMFDq+cJWMAFviO0cHVRwKwos25X5gKyp/6MF/6ic
7hC1gEaUE9f0f9CzuJGvwPcypUx3i/zW5SjNQyTnETkLkz4ybWQimqQgCp6fjWQIQkhAhB52CFo9
PJFvP5SkpJuXaxGy5QQeRL8h2T+gCBAGkEef3CXhY0AoJutjcUGq1SYl+BMC67yZ4A6baSSqNLMd
BAbglROetCccOqIpZ40EegsnpDtG5MbQKVrACYNxOzBoSDg7m3lL4VKP9XVcUkkWLVDQqswv0tp+
ooFMLNLXcWOAFhK85F3aYxj1XaXhB+VYny8VVX0DVp7FCsZsbE/WAyelxZDVWD6/81a28rAb/70X
Rxrpalt0hHdgSg0a4B17GbZA+0UMVUcg8rcT/CM4g6X/rHJIo2/SdxZeax6S3ud76yadclLxhU3k
Xl8/VZXsvov1XU2Ebu9lKUOjT5IV/KgogmTzM8uL6uD5stHwqsa7796YvXsh230JkiQZN1extnGq
pFzf+jvWstE6Gt0WUv/v3f/OtGspRs14g5fwtLZKnZlbk2quaxQiEOkGEcjNFF+PUA1exrtbl47T
3D4h63uDAGyXjciXX+utNE1azkgr9oG4U2JPejgElHimLDYtWD1Js+B6nJ+FhmGMcEIYWH2jfRF2
N7u0/gVdue0/fuYm7AUtizjasJtiu/CvUUq8aARtcklGaots9oYk3/axqves1o02Vxs5eHuj4oWU
4cAFob+7sOLvX2+27SvZ1P8KIxxB15mLhBRVr8j7CInUaSbYWlAv2NUkFhIeym/xM1wZP6U0yTiA
E9Sq+Zz7TD9quGFlQZalUFYFJCTBTGVyvhoE4l0iRljxLSkBfrafdn92HfstxDKq5iV6u/rsVJaz
LLft6C/8rp0px7Nd8JbZ6n+zlxaISjwFbFPuajE4eXSDr3d2FpF3XqQuI7+OFYizx0FnvCJo1Zta
raNI6OvNRC4Gj9Kxrvp0vIBXjzwCrj9L0V+f7g/Ku8NumrhQdUVipw/uj3hKiZ9d3abotWOaCyPF
O3byoATCARZxAVmoupjTZFQaCKSyKQqH8eRHmSOXZuwBCJcshDFJA1HEovydfwieJU5Y3d/flwsH
0yjej+4mzvb1F+egrRi/HNtJq4DnR5Cz49tuZUeIqh7/RrNWv6sE3+eQB4p/TzrgY9EQRIexHNv1
T3iKwYzEILkdaRCwdVZawA27Ak22lvWyzcW/X44PC1MGvK0Tz2yWmuU3AqOoTCUCfrVHImrC3LLS
ZG4K74bAeTyIuKfqPWJNwneqcJWz41aUylgfrHYC6RV/mVRkGjv8hA3kMljnWw0Z2zOx551az35D
+PO7/do5WZjfPZ7DnNSRneoykVHFjk3yEWuz+Sl8k2g8lwiSeH6ze02kT5m0B/kHl7DdcHZQV2jD
+kVv7IYerWvQ5/OUZHXDddGxkgTLYe4gDVB7Ri2DCRxCMKMd7y5dhyJt0hbzOE5x1pGs1P1f9ZKZ
84Bv+oWg/N1aPH8RkmcERN2XgylyAc+N5jR/ZXastiaGVwhxZRwW26S47YpfeUEsBtqvsj00LJ6+
mAyNXJPSyxSW2AFhVeXTvWxzbJT+Vm/6fCBXsoSfL6vMU2PWiKfxElTeeIqulcaBXPTTpMsMlJEK
QFeQdpI86vjmv37r3J4zcayy1qDQB1fL0dPt7dgmhEN3fXMPGtffPo6z9mWJ/E/RBHZdukQnCAay
HLY4rjhNf+TVMSAVFTvuLQEWMjoC4K1IMdQscSrbfL5vmpE6jBw35UsYIfuq6NGYTZ9LoCLiSpvd
pF8uf3CRLUJAczmVXEqdpIFb9JTiJnnXmyRbE4tM+UpMInGRPpUP2rM22W6ekXjVjWeIEOXuytzF
KHXxVUDihRLcGOD/NJp5gGICOuHbS/uC/kdKv4RNDt0JvPHUMFJAvgwPuHF5OI8OPsfstY3WOK53
pIDKT38ZCjAc0U5ijRfXyJ7Er5E1Y2mzwTYTwFJqKTWT1MjD/pX+D9PxFpnqTpWgpsA2a9gKX/Y9
Iw8IEldz9vYNlt2gaiFjRKzefyi+aNkkxcwYKFUKDh1ZFVY5FdF0+AGvG5ogD/SJFNefReSmRD0C
vXapoQHjMIbIJDSn+lOlKGrYcYbmeonAPFr/45uBPgcCHgphlXFzjdjtooRaara8j4+4i6mp9dvn
Yq6rw0OjgyjOHWPVHmLSq1B3aJIaz9dd/RvLBYogAIhJvZEp9gXa19U60Jhq11YxsGjNRqWBHhTc
wtw+dDKlYms/O2Os9ybsP9m9B3xtn5C2eCHTtx7ISDFuZcceFK9Vdkh5nZOT9rNoHAAL2mjsmarP
yqW7nTQMRy2dw9cHHuyeCOVRqcxrkuELjiUbRihU6vXTRYcZXCmv/Ck1mB5ex1mnZLelsCdFHz48
jv/kYtdYvbTRnPRuvjZU0VAAIaAoV0iyx2yovqLxdbZ7JZKS4l4RCxLqdO4J+Q6ma6nrjQH0V4gn
JQ+uOUUAaUZlnGHmS0Trr8fsRV86RQb7sXn5XOYUSzpFZtWqJwgM0VM8rjD1DflBxhmejVLRCV2J
DoWpsoTxf16gYG6dyVdVAEu4uflgm0RGFSGGJ9bJzHnqDVA2MKTzjzCI0QGORTR5CWIa/eWVYu9s
3VV3KEwMYTurvhgksBpGoTYvzndf+FuleSfmhTc2SyQmjutQsOhCE6VQLr3WYeFAXTJH9AEsFwcT
1eVIsCi21CfF+GWvHvpU5FVkIiVZHmw80synqtiAjQtu7bBs07SHrGoAyde0wcLKiLqXFOyA9PDu
YizKps84GufxUdw+bdHntmdDG5Mg4bCGs+tIkmt9RZxc5FDq5S3hZmdCUd2t1TYYoyrXRAIx0Yqx
440xQyH2jjjjhUuyC3H8RYCV8NK8t4TgGHKhE6BJ7zBxDbfL6aemF/rGWnu8vHhYIhBrHib37DNM
CjAuAefCyVNBsdqUxOyap964tcMlipKdXX6ajgl+YFUpJotXZZcrFyMXHPbiy1qM9uItOwRfl3Zi
BGs5dZA9aqUdl4KAENQYQlpnah/92YrIl5aDxEbLAf9Y0kboA3/Nkojzn12HlFjnhkwmPv2dFAZd
XZ+ulH/HgUY3W+9g5jeHOdtcyKJdvvsbqPlb91E+GeF/uWJORU3g7/Z2sVySk/vBaUdQR09ooFCm
LF94JwwtPpaISC6r13ukM5fpH62SZuzilyzEMBtEYoJUwenUsjo4bjzF/6tDcjP8OZprDbpuKVK+
O0g8S51KQybR86QS1RrilpGpVrEqLWllyan/xpNTYaSeDWR5MuESOweq5zd8evaq0mEFGwoIva/E
PsC4uqSHGtRLQekg4nGg9Y4EhOPCT5LD9j4yJp/7hR4eL4zs4+zDMyWQanxeItAtHMc7VXMtYPVC
y4DmIJmsN1xzjInEgKGW/ohrBlQKmh9g0B42c8nlkuGRg2oWgKcDdel88oxsAYi4Fyk1Uk0050JX
kWTu1T/XuzFXVb+xHhEGel8K8mwkAZWAFu19dcj2BM7h18Te1iuxnuD5acN4O8cnZQiLk6sCaRHv
FwHIV6EaSHEd/ANkyCEK+1H2iPbGP3rIwbhogGfRJrpYpq526fyflvivlFIjpXPutL8BLgUlqfZz
UWF0bH0iqN74xT9Fgg6U0Gl4FMSjERftQSs4hKBYaJL5bco06uPHLap8iC0r4EiFbkWSZe8Btqa1
/nDUCvTQ120Jl1oi/mQqxHlgxAQj0CpcjQBpOPHlFOrjy1afd/b/efOdAGW6cJLeFaZ+7JAFDikl
ppPCIijLSw+OiAkYCa+wH3oqc0Ci0Rezxtv9Q2kSrSER2qgvUxOz0gJec3YluPw1kS2DOKCA9PSO
FFdlIAB7h394+cMkDvO/8NVHNc+vm5WZuT3LmKVfwxXVLx9V2THOVHUZXG2BnZlhzS44RQ3T4uCA
VkF7r4gX5I+TCdedtbPnjc5Zs3tnW6BkkaoRRj9IwDQ3GRvnlhC+Zxry5Mx09GZYxxRue9mBYVB0
d0xgfFDjdkm3jnzxh2L1ON8tjx4APAUE2DmVtEqWO75x7YtOE2ZwwEPZC3mSSd1nQf1Y+uM63wAD
ALmGG7J/gbxhBHuv1olQ5bvuYcDfoTocd+Jq+Ct+s778X+qZnsN+RrdQzWwfAwDypaSsIl93ZTrj
b7J6xRvPdqAmTUs0ajkLkb2htnd5G01mpjrZYtZsjQx7OyKaFmFmd3hEGUMs295RewV3b/PODMOY
NEL1G5St9ORs+COp1m7ekFfQNRNdp8xkgRzTN8VVE5V3bfo7OfcaCycH6yhBAaNqrcQtiZ+vRsEV
1IsM9n0kulqpNKC0uSAEbkHExd+gMSLGjsnprqH1p8J1KAcO4Sqj/8TRQq8vW+J/p6oeQmc/yqCZ
pjekWxj/ftzuWYBCNnlpyAAajeJZsj5cJM1ccAOteb0ZaOCC7szp6Hrfa3M3MhqEnq7MLaQogLuq
+yD8xH5MFZuzdwqK5f8c4tLxUk/Cu4+pGYy1aYARmchAX/a77BnzBLyAE3iXOO8yHQFSBQzpLGBX
N/fY8eEAHiheKgCpxw3usbpVqLyXYJCHxpdOBFyMJ6RgVpN7+bhI9Y3gN1Noo+UiKiaTG8w/rZ6w
8xMgf9h1Blgz+nrolXUvOj4+nf6RV86KRWkfQuxgCfqoDwEe3tQr7fb8f5sRaYKY/z78DS93bWKF
pbr9Rk4ZSDSrvgekSinQzzt5/hLFVBf3Hmcx8xYIDXZRjpdRlInZlOmJC0mvBtSZLc1mNuouPK3U
Gyn11LG/ux0L6+XEd0HJAIBlchYVEvQU+ZrA9F9AhVI27nJPFFS60tzkXcSM3c8nKbqLlie58yKO
dlUkoRRsG0AkoerHhOk8wzaNuVn7yRAQ3EfqfQlrO1M8EFh0F+8qezB+TJcnotiH2Br/jJU58oeJ
8XwqBKXL5RhWv5/D9mZ2OYstRkOcs0Gb3BnYDnQBrjJffZ7phkZppC6eaew1kDTAX3/1TTXAD9He
C7/H7U+bL87rVZdXd0b/H0a3bFGAq53MiOFpYtx/mvzmRH79gQHnuly7twZn15QKUqRMcbAOEALF
rtPCSxnfiyh4muOHV2Ir3wAFAerFGI8y/p8YsHTlX3V48tHQIRaAjJtys1iSe6gTKICTItWW7Bur
1HyV46i9nxY3/XczfYJVwVpP+9ppjloGvXiduxFlQ/GJ1OLhoJyY3Zi7N+5Iy2S97B4yASmBs+ck
rU9RwJjN7OB/eQEDpNelfzOYLdohp3D01xBdogsykaB0xSRJe3AskFBTmosCCay8g7OsL11Uox2T
EqUtg3hYBWv+b0wGK7eWqT9g0vjHdeM7q/KB/OjVsbbeWdNikSYop8GCW3FJqNAok/90z7jHYPc5
gTvkAbWSOV9VUonJSpzk+QaNeZQHot/xL+EQ+VwMUl+MLQyIjxWy6KRL6Jae/frj8QYAPksbL1h3
/awz2xYrShdgVWY40b8V3hNc0c5Tyg+/NWpSjsIXUX+LnTg+SPayNb5jBbSWI1L5G4jzRTC4tdeb
ppPXyXjijXuI03K9MZxmE19wrDuF2pGOofWxaiZoYn2a7Jvi+Ggx5SmPDHSWP1SbG7kwcQIExT74
maOfHa4qwHMR8+JT2S/G5GiUUbc80ZnfavK5PdPaCFEM67x1ZgFVM5T/BM/9l1mLHDzP/TGqVpy7
3O8kmvPxe4qrWoo0q1VOHyjiWOaewXGyxVwRCGn1OA1ODQVwpgb162eY9I6lhBIdMaoihGSCquuJ
CA/MgWYhbk/Gj/evfvdZyLPLGcgD4NUic2xgjj+9RPjLfWBX7hX2+v9uZwW4SbNOjcq7Wcaqctan
3pK0PZdzFwLsbPmz0p84X3zGY27SY2ZKlSvNWHH40+/QnvYsC6rE8KbUkRzXL+ZpKd9nYKBQOnPD
ANFgIG1NN3S4q8+C0PTw/+X8DB0469LiUQLaoHAza0kOfQgb5UeV2jIlObQL0AAI1IyF6NxJHg90
W7EHQhaewhcjYM7Ig72llKEUjznhrHlxNw+lQnlNU7iaHJdIHtLHkk6DKTAYroPR8047lLPMHxe2
4dZd6bWBZbxD2uDEQPNGsat/321U2NG2C4oUQz5YE0/O3XJxDI6g2NLjdqvD9wbKPS4UEYJF5Hri
rWxnWQRNj0MZnzWSWCqZMYsHkdFcsvFWkWHaG/9V4zE+7E4wV/z3K0lCUDpM92qmnvU/Ufy6GEGZ
UVIftpZ0zz0+U7YA+8/5kI8687qEmTu8RJVjZjuVo83QQhssaB/9QtMXV4wpFV1SkpmBSa2+XgsD
dh/mYv2yCA/t4afvWamNI1rLU6WpoxBphHIxvZ5C+xVsUZCaenOrlmK2lp5HEtsFedjTb5th5RWA
1s8dqJDAeLQxWpuLSOvcPyvJzl5XJJYMV+miI7EG5xTobSywG9Px+ymob9tbMNhl7VyHblUdGRJV
lGIcalC1FuGDrcm2laHT0vWXv31iufdGhGN1vcfhR4zPps4QjeQCaIklEt+GoerSUW1eQnytQgRt
gVqf9FjOzrIr8hMO7+52eGklG5PHETaxsiOmkVybk2tvwC99udS1zrCkoIrSBc4JNI7ITBTmuEz1
zk0/ENYb1wk88+uqjK90eC22EJmzbqRXRTIso3CiuzEBpUVwYQXu8+FlrGM4+WmxLnRt1TKAQ7Wy
5gCCzlnXlDs2LWRUwzus7EeodASHSis74EqE70HlXqisWI3iQ/BaKjK2IhF6uSYg/CdJf9KCshfr
fEu8d64khS9x/FHprCOV9jP2TvB9e701x9gvJ9YbONAMPLXF/UDpLZPRV9sk6Va0S/+rH8nuAlWM
14yQCC/MgoBHvA0OgfI4Cho6VrUovU3Ce1UixRpONmh31nIuI6RiH44QSU3Tl1c2ST5z15/bxA47
AjvP4rTtDHx45rYdnS/JNqekB4m0w3OwFXJe3GSiTXllMWYiJlWIUSy09Sd+5VPqbhOjM0v7Rxba
HlgVyoyaML9y95yN3ghLML/2H+VGnPUOOWcr5FaFGga37xDErSb0QyTvxC09UMDOuHCz/3kxmzWG
Pojgy7aR559mwyldDE2aMgeeJrb5pNoUNj9R6fUVv39D4wdlKRUUYUvAVvZNW5QBFd3p8XpD3pOJ
THg8G75ogqCGZjHQFZI5RmDis7r+kev2ZhF/1Ovk8xj1wKdyoWtXv+qyCWYcC17x2S2oXaeiDwHP
yxQ1xJ96GToCuVAW62NJpRMdpZORQ/GYbyhkw7aBy7BZWkitYE5YkN64hLj6WIJFNju1Hrq05qE6
LREiY9UCjNwXYsT/WehEDFXGZuD0kZn2KBh+Qb5TlM7gSh4ZHjOpqlHVc/0ibBHA+8ZMH8D88Unh
16o038M9TnR0Lq6rYqecxoLQeTyqSs0qPeIzrQRmahMOS/EYT19dqoJwOLgxXFlF7Di3mQwcuVZH
nKQn+Id3dao3c9DAL5AiEyP+XjmbjE8fmRNTYglUkj9O4vz8Hbq4WdZruCh1Uo8GNNSD8/dhIhc4
EqYdmOjbo4QDXCAUMLH1r1SFIQYx9ro+ousVv239+Ay2RCbzbWt6tuKgd/pNzqigqvpeu7tUWOSz
sAHs8tuQalB91DybrFy5Nx/8LeGnbkmY66a/kjvhK5adogH97EpPFetTDN5cN65AE/x1AOXvdtBM
vRiYy5VWrzWA9anG34RdF2wsD14mA8urISwk2k10V5eQYqK2z2h4BZ5XNWdAUQp/+i2yZzsC0hOL
X7TnRVfwCnWQfdnLifZ5pTqDs4QkTX15X6qWl0SUYmPBlJzHuflWIpwqiXX/OaGaOQ9230Is2FLa
4fUCnyoxOUof9d7T2B9oDlwx9x7mujDsv2ixmY1AwNwrcfU0cyOofrpy1WupPjSHychgHpEdphQf
52R1QsAKbvE0GVTWblkfEL911SP9b3ha5rby89q9AIfNeIzVDR2Npl1amQWxlzvEq+C/Ey+vGuP9
U3N3xlJEx/72fsMOAHrhd8DuDQOeYPiw6NtAkORZZvSf38pLqPbDXsGTIkoqh8jxuJkh+BWqKBsg
wJvTLFqRrIXgNjumcQKrR4Nd1QW9TeCIFd+5R450k6WYm9WIeQ5BQYN2nlIhadQF9cbok3B9ULic
vdBfMb6GyEURZBUheuMDbxmKR48KjkBM1rIEVR6iYg7LtjMaziLrrBT8ZWyoICdxiNhjUOZJBl7E
c2zuN1itljnx8rxL/panVddQ+AZG7bW/Nt6+N9fHhFlHtjtnr336zkP+xqMaU7hGiMmcpnYX8X4Z
wFEdpQn1rl7ZGi96niIecgXLyxZ5+e9CwqELN14BbS4ItLhb5l1/y09bOR5NM5rvHX4qFnGZHKAF
hPPrllfBXjM3lwhMPPLpFEToSoh685JmBt/GxGnDT5SxqVM/QrgWopgq1SZSiQm1UDhObCy6tRVW
l/3uTXhfz3wQZBZKayq9Te8SbcS3T9Lp2OJYF0XcK+YxiF8D9fJJWTaf4CExeRJ+SOLess3pcvHl
xNhEHb6MXxbE8LFBe9rMKGj9CcFPmqD1k2T3YTCrpNcLVe/44Cy5t//4fzg4B81jQajTUKgyPTc2
IEVoRl+gEScN7b7BIBgIpBmI3OYnC4F8VtktIMs7j01JrsbvyzSKJURJtTfQIkJu3X1Yej9cZ8Cy
SXj4hr5ulKXemNBhQL4MQr4rhXRswpfijWFv1EOo+YqFj5eVnAl+LENQexllgHb7KULXdfWXVrMx
LuWkucZUqW4LmeVQWVT1QPHNKAjLjpYqjNoB8DxKZEpwMUbqfePeEdEVnvFfbEJsOYDJhXguED5K
0c8vnHR77pgC6pJEzg+MfJve8MDKI+xVpaWkMSyL964kOwZOdpmB1coaZZGqhHp+/48WLFJvxy49
43BJG4FX1xwLwk7UqYd8zn97c8LxDn5B+STU43psHs2uKxik2mRFhvjb/xl2w2o+FV6zur+LXCeL
gTw8vH2qohDu8UKifX1A90mN5iU7aL47buKu69YM/gsjyF1nCfVrzQD2D8bc7P+vppwUCN/lNMNV
7hLxtAg7+H54CY1mBmWdwFJLe5+EEjquCX7+89PCXcbz0bX2ysHUcXe7uhopv/Ugbr17h6CAzU2x
KaZDFcdNwH18Efn3chae3d5elAkjDiF8L0iEVeoWJcliLcaJzHybQSkxov1pnKnALKnYggIvjIVO
L8oIRZ1NTVvw86/b8fD8Pxnpn2wQA6f+YdIOhrVvFQbA0Kx5EaJGpFpgX5pGxCGSeNa0w+vuwsy5
c8F4qZNtWg4JKwCwOFvPV6Y1bJZtSFq3AMRxvQEe1xcVef0rskf8JDFL7CO67zT+dLOZgoymS9MQ
nvhU68xnPuPCjBg+yM1fS8nVTqQxYT54EW9lxR3FbmWzGdDHV5HP7mr2DY6DATv9UL6aT9hE1Jdv
oXIlilDSk2UD7EV37vV+ldIwYMmintgtWha2V055fx8pHt9OEzi4IzMLlmSarYJWq+CTCtx2Ud4M
zfu+x9in9+KUhokiJssm5XkjM315tl1ga/mKpGztyG8IizqDA5FAbTJN2O7GM9MVzodvZExlWUCc
45innsDVi88emI+uDbvMskpUWRghNumsofdX3cIhBhGIo5ZxZjFJvHA2gA1VXJOAmMjLV3uH/jRq
fip2DbLLUIxNIW2uKIOYkY/ygXjdRsFfatIm8fJ8rZ7a3jjosNg85hTjUFb0Rx25zg7eKg+FTUJ4
aFEQ58l778oK8e8qyOgqAYR1OMKP0Y5LGfRRmZJlKOXnHlZnyJbSwYz4jVewC1T5/4lwfW08r8Vr
7JwujsWchUMiU86EgaxOZvMhToBZd9FU+VFIxvDZHtjmOIr7RHqDdDJDnB5bzcPTDOzpZkkOFnet
ghQ8ptngRTgIf9LRU5MGU2jxmO1ubwW0VO2K/wt2PEnaI5Hozf/lfZPSWRdTnAn+MPpDkj5saSij
5b+2U2XbJ+tSUYPPjGNXXN5OMSMgTCbWmuq5Jx2NREZi4iaBaU5xvHCoS4JkxrZ7NcpO3+9WcUwB
Get2hLlEVNhREJN/xNfILvJifw8rsoU27T40smVtfXFLpN4hAPRfGYZTchb0ME8Xp9womzmuhUtU
dpNs6fbzRxkq1iItA2xKwFFg9L7pRaBtlOu/PA2EWoDSC5LT8iYLOqyPSJZa1Bpief0Ac+fuBeYK
SKFuvfH9ciJbyv1rn8Wy+teoIeiJEpteCPblMH0BEEJnBU8yw4MbqGYU7QyMDp9i+TLlaOdfWsQa
XdxUsBfU2jUBGWw2LvubU8JCaFCGlGelBxUwk/gpXJikkcYO+rZP+ir9XA2S4fNdeaPRNPdVU6pr
5O5PMLco774vjNZ/D7DzS1qz7v/lT6Cq5u4yFbxm4q7lk28GUlOC620b7i98EYFpFtB1UZzUrBbC
/xxV7sTIsz7Yn8aM9Y7XIT8ctj6938Q2v7/G+7z/wThQ9nXz2Y3QTyTu6fFweHgWVP40URrYyObG
fXfY57gZuemeT8yHs7VkisAPMD8Uo8xR8qbfrTDWyJVR+uiMY/XblEuqFf+g2K8oc4nmLgllKWFH
IZ484vlGaTksP25gO77AXfzLP0oiV2R7beNlQiUQRqoEzoR73oRRKDF9H5VgbZpFy1q+Y4pYHrCm
d4P10qpgKyQ1RTofqSGYsFSMIxc8qNXElsakLNYZExMTslY7mL+ahcEdgBHCSzJmLvjy5AzpIXEm
vNEmHAf+zwLtuBaCYxNm4rPRZcH68njVPXmYvnjezreC4FSNKxsxMaPrShTreRgNzar0LFkeFXBA
71luN8HLfQNwRVFZk1XDFzVLqej01IwMwYnvhXN8E10vnRXlFJaDS5/b/pW1ZqUZCpgGW/jCZ2Bn
L16cRjx795nFSHXCW5ZHOrije62LkNj56px/fMdwkYKNbGGR4GP4Y8VL8EOJIIwy1Xb3Y0z9jwHx
IIU1TJIf9Py5q9WyW0Dc37zmK96bEQY+LNvZAZ27hQ7Wc8AiQXf3Rx6F4MjdEHCcidr+VHqySMBN
y/aPD+1zHMPAMn70RbhkOxNVo3Ncg3Zu1NSRWF5JbMX1df40KbGBunvxu0iftmF7+AaLaRYAltU9
EcUeomGlcn14zFDkJ2v3y7i40btkbY1Nxue99Q3UcWV+lnAftkgnHmlGlagrJqli9oalvZXiZiQ/
/8zoCymVB7fcWiqkPAuY+BnSa5hQh8O4UXB4NE064JzPB7eW8uGbGVqOcoKAMPQ/XskgMQfzZhDG
KCGX5mI/H0hvnVGPkQjvjGkrJJDyTsl3rZjYRpjspum0fAK1CugSAAH6CQHBDTE6eYJO5ZXB176J
rsUqlP/mySiwrHmJ9yxjhJckCn5QQz8kjMWpXirCWE0WkQF8oeBkLOxcSZKABH6IROM+D5TfDyUK
+DKsXp/FB0AZ4lRTn5Vo9sfcj7fU1IOf4zk+OkdBSl2DF+6XFbmjUPFvE3wS4BzsdUPey3sLTlNK
XLgh77ioKp3A3dUWH4GP9siyf2xcoctUFcFmqO7emgr39k+qjEhyHBkTBuHiOPG6IhdMVyA9uO6L
fHe3voDHIXcu+Rs6DzPen8rJlYN27gsly9zrhwbD2ekYiNXEbjHm+pQGjTs/IU8VA7AjCsJRCB26
HbkUeOhKbpRH8w2p/pOZU2l+kGKpOBLi21FX9eTdg/fQDvTq3/k7V51OFW+Fvszvk65DfVFUqwr8
wuqj/cGfhMSU2fgg2oz/f6YhU4mqBC4QEkEeAMgfOYWWWQDJzyUcnH0zjdeAn9nuwkhOmdEEy2Zy
mwbR8OzOJfE94IXWA7UCPfDaWLK14rW6wCDV+kg7Zb8f7xDZ/Hb0UrwVColBN6nxieBY40E9+zBt
ngQlCQh61gyrNCmxYZQZRz6PYHbNy1MBXoj0IKVimSnH8+Htkox3x0I4gU40+u7zYkmmaQVzRAU1
wqAJjase1tHih7/jJenjHZxzulje6nF0htVSCysRJl/QTr6j1CSagtBOVvAFzlPvhKbvsmduonAt
2FP3bhK1xRyPz4l1PESg+Zves0uy7Qq+kKk5GQJM+5mcIJnCHsnYCum/1n1643n3E7Ouil7NYvkM
EArCqPvYjj29LDW551DzU47kbY9pBQQ/x18Guht3ZoniuPLULD70nqLzqaMpTngf5VaFhN15vK4J
w0afw6efJQ/k38gyjiX9Xl1AHAs9TJMO9YAD+J+54bm+x/6h5zR8q56TB5LECMCCWQ9VmUvY944Y
Ik2bzCJSpcUSC5wlrScsezg2t3p6Y/BXPyNvG09xqolD0I4F0KHtFQazQbY5rOeBbZLrUYaOvS3U
qacow0JbeMUvy3ez12c8Vl/sUBCeKG7UF+j5TvPGhZUfQDzeKco9YjpaBOZyzX+D4vIVteIY0S9C
ILtQYHKtaES3VeiNPvU6ePg0sRyNWoVViyEykRFYp/GjrJEyQkj4UMtTzs3BT6RDW+P7vNEfc8wg
Uy2/NHMJDEFEh5JCM1MGaaOxoYEsObcIf1PXydPVZxpN3wmCWkO+JD033ORFJkcDRWpCJ/ehKC7B
txTiuDgYHFiYIW8GeRlmkZCgoGjPd70ochidunVkYytrn4nzeE8D+0tKqFooujhNX2Jv8aaaCqw/
SIKIr/xmRU0LCt59k7d9iFdJprJa2kzBkNo1/u+XZchXLbp3OpkvHHwYllMSbIv1wcJ9QZzuW0Tf
kqkHLCt689S87mAVau2+dZt/qOTN3GW53mVuPmuPzZzhoJh/dfUITni8EHpj7SnVvyM93dpBqH2t
8wglP4aHKlzVWV7xcTFmTldh+59P8a7aaOp0j4ETJ/jNu+bzPiAD9A7AjFcQHMgfSXtleA66Aln2
Qm6aJPkZ3Zr/GA6OS6EcyEG19DQPYHtu4/6ylxwzsig+Gr2z6ImdLKo8Ci1qzTQIKegx8Rf0ov+P
mKbaPQoNh7FQ+IfGaBpVgBc9nquyV1pbLV73IaJlj/HdC7Gz0wBVNJR+47tVhRzoBPV88y1JLtCU
JukZMkLk5l20SfXND8X9lbjX461BquYzLomEfsVBeaCAXVgmosWxlIwLEDagBnNZ6wQnnfZ5k7ai
mRWEPT/tqI4ak7/Q9GiFqFobxAi5I6NVbCLs1QRDiLlBFPWr5TT1qeZ8/Ihi4Il0CGo39GUmgtBO
Bs0Ei/TmVvhV37BPImXEXSVHMqCFYqTCRavcmBfXntUSNHASOvvGig8jrFIjvR/hEvQc9IKiPWYQ
sPShmbVVvgGmZOI9bmBYfuXfpWocni5T6mM5+XtNXsEUPVlh0mYNu/be6P4u7W70kzkhvj4lnKUf
7TyC3HsraF0MsOMuO0y9URD1ZFTyzOUBhSlVejcGgfcmUpEY1CMhl++JZd0N36rV1r/UVySiQDe2
kDT2xhOadz4LFdJBy0DwcxX3KmL6LtQMrqWTiwwBOqmeu34hsG+5EFVPN3RWz49mus79PiK9r514
l+6Qe2HwDqTEZeUwdF4X7/zsdL9ycFc77BcdH7n+chV5QSU+x1L+/2eABlCX/hLl0EZ0SyxLGgLS
9sw7qZdvGuKuK03yDhevvImS7UclvKdBto5tmBRGwDPuV6rYxr1+EuD+byoHFdL2gXcNGtpTPqKY
7HuD4k6y29Z4oUa+s4aPXSHg0BcayfC4nt8ycgkUN1PCaDVlPlOwyxYuIb4qtIg/U+zM+villDat
p0oTuAisW/ComZR08P4hhfXBkNXB9uVM9mqD9Zs3pwKsrTX5uoBESUHvMDMKHMBuwJHXaXE+CEyM
SYEuEHsnRhuXPn57QovfDf77lekfEL7wNlNi8z+BjcTCYNPDxc6r8uwc6XMo2Zd49dkan8MBHLsR
YAna2wCjCRHWLPypmiumXpOeI4FNHywShGFUIauzMKzH9AFpS5OZc8SzEzBdNSj0wNI/qG1A8BMz
CatYtxBsyhVohfC1a8UiOXdQhvmy84VxBYKhLSiJuTqqATJ6XTu7lthA4/ZcNuZohDNPzPFqY2D6
hSmLJHtz2mGzT/YipiYswd0DIGyXiQ49UOMS/wMOm/TAo4HZWMvQJE0qrPSCXv1tIBng6fvMnvg5
fhqX+UR8Lzg3I00xc+gC1gBs4FHv4SyHN/6y8P/Qw0wCucjYAE0UnnyiN4AN3wYeJXM9rva9AlKC
+UwM5CRpajdQ/a/ifFC/7kTCgVJK4wDwad0FYojNf1u5fAik8jtKlZE55kkgGRMVz/sqVY4YaGkI
ZhOUb5nkYjsv8+UZpxPqlTGu0n+MT2tpj3cB9fgIqQaeIn7EmTEjL0Fs5JRLWuyn11SN75amJ5dT
+VaabCMo+CLU1pQuUGFoLKRxP+0/2bvT8hMMNJbEg46eCfs+SgekPGNOJ0A7L4rq+qgjua/tyzG5
dgZD2Q8PGfH1DGfbge4kVAdtaCYGUJG9yZW+bLbZsgF2pTWGkKk8MYPUUPBRL/4Hxi5FvJwHa0ri
2DahfCycsB3gRDJGhimwDq1QCkP0sSyx3sjWwoTF1E+OxmKQ8c62AeHiPsmIl9hAV2JHR6WkGr/Z
/jIFCRKpyYdGL7T/GgCOQYoGcGGIA9iM/0lXCHxBsKgBeZ0mjfG0SbvpxhEhZOTSllzJxnm26gf+
+G53P79/KH2NO2uerpgM9AXCu+BgHtXjgMX0WZQeYidXAudYd4vOSJTV2TZcNUUXm+4xr6DF4xls
yW1P3UpfS2d/C1x8X46YiqeGzkJlGDQrHtMnzA83+Z9rOTNx6xvbOsC2A+iug+Um9tallDt3l45o
KtkEJoLlddGnuayX/vQMRuhOWH8Y4okTybiLQPkU5FGrpdVSnQneJkw5Q9W1ErIXkAVe1eTPRoQj
+wP94K4AoS7F6ZanDGEySQXaNHzuoHKW6cMJzBRykLO2RdMrxl1I91WGFgVlkWbBD8tZx/Whs/FK
2D72Ar4wGRPLWGo5VsWZ6yVw5wHA53otWE5YhtDEF9EVag/1oVTlZ3Pl1+CcoUL60TkYu9T7L8wg
LnNn2YJ3HFg5FLSaNAmVb3RFc8yUTYS1Gj06WG0gqaAnXGgo4L3NIXwbzrtaHsH7SBXLv99eFXlU
tRSGv3X2mIsVJwu6eMdtNXRX3lvbQcQfpoOao3OjT7g6N2pMamlaBLF6EQXairdrxkbmveZDh+zg
JGXv649Q+zcx4ex5HOu/wmXf4xQvQOPQKsylZ8Xl58PodLnGXDnF/C862YgNJ3z1tdier+bfmPN0
9j2dNIhtHXrMDPkk0bHCTzvjoTHGXGbtlVb4k2Ut1cE/0XyM4VZiwdUIJiLCPhrn2e6F3oeKmxdC
fWZlALEvemFJ8lHepN767l7AKts0zUWAiK/x01fKWbGN35RaxBYeY+NpTn4L7hYd1N0EHQtMX38n
7ImdHkomSxWYyfin1E0PnvQIHmDlvnu1myQ2O18jHoOW9eSRMk859bSoPTLukwZnlV7LhzKlCIOg
lfHCzOdc/AkvQ8bDz4KfzEUDvVw4PRvT2R3mGBktLOmwBeT0ofVYsYnoXCORhiPyu4X5Y7TVZOES
cZ9kY1rQYUeimd1dGtI5AGByvx7wJ71nuzXkoJMDWdOCLxLVRVyxEl/cWBg91ExQwN9OyTCpdzhP
Z4BA3bVkk5AJON5MDmafCQ2dBfnCci3OLVGUG4vK+PUNuqeD24fo1WT8fejG8kPLZUQjLxlYPHMY
0+Lf0xN9FEwt5Jkzgjj7/hBmfxGK7TsVvwH7qXOMwJcouLdl5og2R+pfk/J5XKUk1mSM028ti8zC
8kcXiCiYJ/jNc50WKspasBPFiJ3YDtP+3m4eQN5BsRW7OE5D2CwfFWAAmNx3PhltlCwzXLL6zUAl
aAYMieVdhVQ1H87KrRQTB9xwvjEAWoz7JVZHHD8aMT66izm3Y+ZNlK/IAHMvOtY/DnexylOEcsz9
QyrGr9v03M4RV567q0Si8Q655UQ+PPY2PlEBQtfE2B7qsXg06r40u3BvuXjSYSk9wV4w2SJfLwOk
XKXIET9rqIvhRylIpXfVp/DZW3yaxVXCyDqLwn48Q+6VHhC9UGILWnFYuYWzPzJiFlT3wLQmut3X
bkEsUXoSVnHC7HGEUushilmrj3xuDO508J2DjW58qAlMSXSqgyazbD2VU+TkNAsyOZe+HZBkK8r7
z9v+Q1fkuPFrWPe0sdTFGs94ZZxOSqb/kwUHNajweMLA//Y6lN+c+F3/VTEHex87xnex8PbH65pg
gfSjHsULBVvV/Ydp+vxReB2Y7HoJN00499IGLkfvR5b4ZFcNq37FjOJ724gRsp1W6hVe+wOnnJER
ld2vjHVXYXVo1uI8bi3lto0zRLiYkZEo00JlNMOSGPCpr8sToM/uuFsdFiw5+2PfN6ZNl6UE5OIQ
lQmbbg+cjUoSwjA3fL18w9HL0cgDjcxAFT/3/gXn6DWhBHH0u01V+ZXilgtv/rladnXBUQ6Jx76v
ODyCbRmcLzYRBjEQ5oeLxqpv5DZkBDtLz1RdRQVZoF7gDhl3t6DJ0fiAbF3gNRMKD7BqCpHYPT3s
9nx6A3TzLJhy8xT3ResYC9+vRoHj1jhrsBPRSnyYF77GrZbmXgqJMdVl7dFN45XsYbcUQ0/7cvLf
YryD9VLicFFaP1x/km3RagmIqVWq3hzCzAZMKD3t0JrBKfDeoyHiTjTQ6Vi1t6/8XeUWCTTTxnnp
vcGPeWJXM8qxPKn7KEDf74FZvlLRLHB9yOOfRHQK3q3DuPgriJWvOdCVU6Lqw9vQF+hybG7jH/9u
4jLMk0AH4aoqMNbli+a2j/+TyNmEBgXShK+pfLVMpESmmoTz4+T2RM4g9uxRWEXVTchCOuUwHU5s
0Uh//7Ked0fFc+2oBaIeBHVRYMGwlha6qMxyFxAevDapE8HSLoWQ54fIOexEm757D711+E0GTmGN
h3N8ATN8048oWsNNZ72nEGDqL/QGLS4RlTpAY/AvqvCvnkeiMmTzWNWhIUmG/8hBFw7ys+azyI4N
615m4HTFjU8NW1lpn+3V53IZKjK+J2fWMPVgsR0oDa2G6iiWft+EsySac3RIZexG25w6uGBtZClh
TyZ9mJD9FVXes/VgS1QdBmN5jntaBaX4N9fM7lrPjJMgxtpfpTLcH3QhBYnTyUBxCdZ4Z/4Fv9lc
9Jo0BA2Ybz1jBoixsiNKxZtAg9fm1L9q1Q7Rq3WcHXSguLj4X6QBZCwpoH9ONrZni1wu1pQf9Vu9
sAZg73q7nbdDrrW0epRvDEaBu+HXlj1cexaJ6O+oDaVumkZnK9sWEVmQ1cEdjhd2tCMT0xuN3eR7
ItpFRQZNKDkEkdUJk9owuemjgUEBvQubfsW7jmbowkvSoBba/g4rVfnBt3lby9wy2OXo8H1dP/J9
qwIbRGFhS6TCWI5oYkxdnI51Eacp1peb/2w4gMbhvYL4crQaNRtvVvRm0+tX8oXD9kmWRtFJlgLT
G5iSG5cP7Z4TaY8RImebuBreRttU9kJYn2jp8TFles1l+42ARHNL745ISQS7jjVygv79ZMsfSz4f
IpPvUKeRtpMfVCabTaQzKtWFEyvZaPaSGplxLhLvzx8ETKwQDX92v0z/i3DvMSgAfvinQwRD2Ki1
nSWaA7fRmuVwXf6mB6FKCKPBS+EC1Sd877jv2WkOpWVMuPAhmojDzpxsiZqwGmHCNkAGHLCjdcZJ
EhWO2qKZ9VXY234jXddGmOFEkS8fADTdGQspbZFAbR9vp4YYJr1QhMTsbzcKSk2U661qS64rUjPv
7c2wdrZQmvyYEW3vE+v+ZwrIuCzbYSwaFbac0HiHZVXJuxCUbuOT+bFtm+syffsCannduTzLNz8E
M/fhBiYkI1Djj9FPEQHxnqLqbmdlaOTToCW5IeBODEzu71bUu53K4GmuC1SNHikFu9kYqQ6w9XGX
SvVyr0rpT/Stjg39B/9Tzk6xDbkqAtqM8Oe/26/0HQDugfMjWIwxPFmwl9rVulWn63CBXmpzecGv
81f/PbcLVgf5FW/u4KabFsGaZz1ia8c/yuPg3gSGdtJh8Z2ghH92i1nsZELBTSevLTNJ33oxabVM
wG+BPHfHGmwV16K9HMdgPAGu116UDlDTDNmx9rKqUzqypezxuwT21x8y5gONgfk1E/Sa94frlcxF
+bHB2h//mccTigb3otB+uRWJDi4UYqVdZB+qpBV1HJbFLeOBUg2GXNSU7oUQVE5lxXWfawjBkanl
h4Kyi/d4lN9zkDMOtx+zytmQxk3cqJoZr6NTcyHoYgqsu0IxBr70ueFKoJVeo5BCZKhPaE3u7I0F
MbT4BmtC+3epRF2NEB6Io7QMPJfn9DDql49AkxPLkd0vXRXgEXccDH7xRvUU9ZpuVWOSklDWliNZ
sn2YLTvyCdQNOA1StoEhLCahltOnKtjLq9OjdyI/GXrvaz+clNzgGiGPLMWb3EgQmiKkRLoQkQLM
z/gLz9bhyTljuQHgAFyHUsN5xwItbFrxv/oVT3sadZhywxY/+PE0nGJCgHMzvsUvT7Pm+8FOj4xx
KLWnLHsubgU5QtLqWIVmHB2vcPb27o8cE1a2exOxoZW5yeBdhEKFpnrkKlSgT6yG0f1QGVxmmlhP
aU6rC0p8vRPN7qlmQWB4c8Qnb/W3wsI9Ml1QnPhey+7rmLuCtbmidH0cMphelR4hBq6MTIdWr8BG
5FNUAcf1pvD66CG1JAkI6IvrVTVs/eW/vCdFyZjb42kgM+bTcQqMJ0t0PkCQ5cXYQMnfX/kR4ePr
pxisimplWj5LlH71FFTaepRMZI9wEuIkOXzGCv3FakGwUBW4L+fU54yVCzV/vHAwNzfZO99d+PnZ
JaoeC1YfqUNeZ6gBeEYqqokXaAul7Hmgaqdi9RStOebrmO1rlz6zDGZF1w3Bzpgwu+uduiZKqZjX
eCnSR192Y3CIjJq+SFCkfU7qp7vBPsx8/5y/tBW8/Wy4zUJYExA5ptPOzTg8Q0EFEdanWXHK2f0W
luxEGc/0yO0RN4xBuhNWLJEgtJNDQdZncObc94Ly+VDvmMINjFdrb+XdCnYKh1/+VYNuN3yn5PiC
Q3Dobncng2Qxj6IaRuvInlNZhjk4knhJ6GeOf9DYJV+qTb4Ihmv0ZHafW2XNS1ORBr+7Hmvnq0n2
Gav/r6ps4PmLnrLmLbaIUy5uiXmUujp660BUP7Obvl75epeMcnowUNW+qN6xTK0ynaZFcxAPNRVn
mHVbL7XxO1d+uP0jlt1X/iX7BTySlvB2wo4jDI5OnHD3UC3jpRMKgdrXrmYxR2KxvgbH+G38r8Xg
OGJYbaL81ywpeWfMkt4ACrl5Kogqx3L0chucD8aRTGRQWzoQtZ3NsOHCmAMsB7U8qBu8ilYR2y3A
yw2ejz8mi9/BNx08eP/0xE4iOGIvI8kvB2E6JPgIthcFVbtpLBSqaWkRWBrYjSvlG0mTGen/wJuW
ND+6z5XEzt9yvliIlULOwUuajN12R1he2//SyWBuKr+kkbOs7ZIkc76Xa3ZFpP4wtOd7xKJSYUGm
mhGSX8lN/Itoj+0fA2gKXxTZeXPCUKzyZd+EKhm5MWjtim/4SBzcGfDb5y9QvBMB2qR0FHEiPGIh
MTSoXYNjNGzKHbrWptuSuwBb3l2FEtjeOjlh/wyfpS1INZyC1HCWiwml65vzWo6XA/YmYHZ10yof
kt1dHVXCRbyojN2q7UcgQ/TjBmSRautfN6c8W7P+GkW2NgO+OXNMJwlKrSj7Q/OdxoCPgKIETwh9
W5PqqVLjXHDhnScrOSbWIFB2Vazc0DVihV1GVvCHnZDdZcyIlFSWtHb9Hhcg95AvQ1D7YqlPBzsk
/2b6c/eJ9281csD1KXh2Cl52FsV2yDM9+SY9icuq6IESImIHXKvDjzD6Wl9+rzQUQFhT0gs/davf
KSeL7GYOxvfux+Fr+LhWrgfaz2AUbtTyBiJoJi4xdGsyvKSL41N0Qt4+tVG5KNqwQT+N5jm+UPJL
L22hQoymVThrT4ohD/fIwfkoOVejNkfLB12Lq4fHQYSTySQx8NLxdq2vEjw6ubdDsKbkU3RseR0n
+OhnH5+HVGIzen/s8m8pq9bMsbLrd6OBxq0qjuWPiT80MZcE51WLSaA2pNRLh4CVIJG4YkFylZ8Y
qC7FNtb5o0mpKxx1t5DHHF6Y9yTkSp5ngPGfxEEqgkKZtO+/wu8coUArpWVBxXF/gsc833kCEnD+
EZDMY3Mgv1gSz1+cFrzeSTGlPYQTaDAIGy+hou0pkGw15/vMyr+KYqFjXCE2bb0Nk8JuhpC8I5ge
6Dgl7yuzXzwGj8kwjpq45wbBWB6o/yHTJ+JRQ609UAQ9Yd9915oxDRKiVaDmM7Y2VkToHE3+PNYr
lth+QNdRo+IQ1DnUj3JGa8uzlov/sXEExWe6TWSQmNGj25WJsyTAcFUubia2S2CJBrKEIMyHC33f
nKqfawOH4NgktoTutQgx9WYGJZDS+WXubFAaPfWsGRc3p7GDds/Ei8xTkqFhlgt1TDiT8QIxNyYv
C/5HP8iXg2aEjy/ptTkV4MwGFX5UCJLBcIXf8Y2tEk3ENL5zOYYx7tmyEiPaUIBE1cizp3p0modc
gfejjLe4wp6AjBSBeDwQ+AGDvtYkeO1VTF1mc2EQnuJIqdtDKhVcIBCEmEuwppwIoip2bmGysmR+
AkpPLyOVay9z1f66EeJYAFiBStahjRwGZHZ4WfveuicUcEF7mlQVF1XfowwwvBaGHt0P9dSuoPqL
yqNIOvdrLEoIhXT22Nd65oHuskzSdOvpodqulUPkDy9zGdvdQZ/Hdh3j4Qo5lYHf7r8aWzdzfftB
Y8DoL8yBoKe6FjtpudfkJAdtT1rw7iRVIRGSneDg6XtnU6ojrp8gkns4zgjuhkmZqVqBhMPDGFQh
o333Elymra4VTU3HQKa+mXmZgOogzNWLEEyrz5Dcvo6CxYTp+Y3HEPl17vz9MYXamcMAqak2bYU8
58K83eDFYyBC7cP06N3p1E0VdF6ZBYnNZ5PyUnLBr/GXZ5fyz0zR5yEWo+sbVc8BUrGNerQrFaCQ
EvkG11u2wDuMdiN0/TqV+JmBupqmTrwGoUSxfKcLARoki06Fda8h/rDEp3TWPuaIK/DvIyqYGjXO
LgiCoOC/dNvLU7FxBxUbcdoFW30gN0Xjrgr6lneTgkXb5L2qXNpXrqhZ4mabVKKWN1Mg00xJE3CV
zdoQKatWmISFM1Ekia3OtFEv599JwsS/LTY6+8SuV+Lgyagg4MS5hir/MWiB7qpn5UF+jCHhxjGO
YHCLaP6mmUDR/47WmoxVtaPfD4C8MtSCB6LrzHT7vp3vT5RBlq5ueek/K3zBQj0oaf4Ywt4C800w
VA6crYRXRszKMPc9etOmG9ZRrrFCpolmABUl6aJ87UdXcUiUrnExFSYTek6YFGwIfF9pje40STab
Z7V3vvHbu3YQQ3pKVuKClaxcT0WUl5jQnQKP0FdEILbBKfhQiN3Tm7Q2qJ5WtfsUy9r825YwFW4O
rcKOJRlFMWjWXFKSKYQceb+sHEt7fjfSwOv3rj50d8udnT81bs0vW9w5rJko2pb1tDQUQyeCK/+c
Cxdq5/RCN5hSv53V3eiu5EAveZo7wUCn49tzzyoC3pCXrLCvPrjsgFnqwV75RkCQgG0bLIvumclD
EeX0kXKRsO/oJwcvXK8XvWY0dTT6gBc9ug1gK0PV2TFeDmlsvNNDu1d3g6ec5Af4mJganY2Im1PA
1up+URhuafhQFn+Pw2EiDUbDcE0+BozPJFdeG880GIJSZh64CZ7aZ2IyEBNxtNW+cWmp3laxdxK4
jP6ImGznAVU/Nj4d07M3PMfcOqltNiN0Blub1nwwYBnT+fHU/e6hMWQ+miCtBg6RU3vSmiI1Kg49
3FQIN8vEhaH9wpozagC4PHYK3LC8/YoSbZO1htbVJfPCItKvEnMJf3S/2m5/JRP0eSipJ5S8W0cV
sF6hRZbNo9UG52gI+ITB4SSYcoTqiAW3supCM5paqTJv/XYxtKzrGsr6a6F3wtnA3/oPRv8+xoDo
4XjaxZMytZIJZjpONY8Q5Esz2zuNCLK8iKKSRHzkFuToX2mjzNxI/oUC9J6iFd+vNHlu3GICWOHX
miCR7FyLRg1EOjyXBp/eQ8mt8AC73g6iL0JrAL6yQMe6QjqnNZ0IT6XD0YsfIOVCvbh4IIrg+t9I
JkYtaLa0IkgSEBC1gfwEJYXEkwqvUhbKR/axQ3U9d+tXKufOCQkJgMgsAL5cuqWHHcFZR6DrKEkq
dj+dF4L2SChNRWtfrMYHO4f+S1SEGc0ghItUln8UZZhv7KIf7qZKlrLppsARw+qJ/clb30t8ZWbq
b5uzvjhkSiY5VrYztRLMZmJwLj+nUdJQGCFTYfxHBFvT+GG8WA7eGvAW2d1qjrPaBzuO/yb5LVUZ
FGWfVMVntrsfw9LhC3YPLDQv4+LNmT0LbZdPnlgU9J+2BOpQ2puEj6S1Cuj+4BArFOkZqx95stCB
xw86pXPwNGA+VDOFpegh7B5Ax808VtC6wX3meu9wbzY+4yloQvpXzUY0J14atJvyv763VrB3MxV9
C1B3DvzwrU+70aedE6th8LyTG9nveSsSyMMf+oe8GndQLhv7f2mRxvUIC9JhUqhcU6ySS5Bl9h+4
pIVqYOSbv1K6VBQBfju5I5f+VkyHxszTm86Tz1fL64znldnyAo0+avBqRaWY78bVqqVoYe67aSKm
YzQYGXQ6nB9uNCuQIvKL0MQf3bEnnbyV/eYyHEsjBA2su7XK0fBrLKNC+IJmhx/Z0yubnNeg3XFO
Y5JaNfyRDT/uesUEFBWTu7WWTKsNusangCGBMQ3rOXrS8ARea640TRi1COda6vT/YoO+rVye7Bnt
TDKLqqDhSAtPtC6YD6HSRXuEzd1cocS851YGYlLHWQE6VUNhXHH4BtJRDn0vz5tQSXnaqbQToeEl
X/q1VD7VUq1REua+xXtVJ4wScWD8/QdKeBbLeaD4fdG/UONQyg9Kmb4l6I1B2kA4TgDipgVQmibm
V5wh4CzaEwwzwUVAe8DcqiIk1VZT4RnBSdqbPe63kCAxk6v+/rD1YAinprmvxLmJx7A1MFNrYdna
5loQxipAONgca54SSk5eUFE7uSAv7nUSzRPYugxps60fUJ+pJTcSohssUEco/+9f/rHS3yd4Su6n
zxzdi9tAnbanjl4l7yJJWCK27XHeqN0NG3tN0l1jEAQb9Nz7SLPqWHYvX/+nbomn+JBTJWP1GNZA
u1rdXz4q3i5OHgJV6cNzaGFYHHsxQp9LC4PssV1kJ/sJ897XnXLJcPxV+Uz9kQanYxwT1aNUZOdd
k9lsfjeVd1GtRxSjOn/uCTdHp+5+a+iV93Kwp0qg//HfHF5OuIUcCCiP/xVMy5MlAdXdVbw8b3pS
krIhfxsg+h/1ySPus6jQMHv9MwYKmJIiB9ib7ZKkfG4y/GZ3/HH7txRlS6rCiFErQanWybn1/I81
A1N3mKwm/uQIsLRyqbXhZtBBCZ4Kl9AZ6QJqoCNQZUgRZWlgTkN8gOTQBwihkIfRz0+AUEmO8cSw
6utIlLz6Gf960/5H6coiyNjOCRy7se/NMeOPaOyXzozbm/ytOSHWG1zYXEaUqFqw7s/Q0J6759rB
g3h+HbQnkbHxdINZvrc5xm4H1EfJYqJnCiFX+J76yETRfwwAJ3HmL6SgMsGsxyFNybjrr/NdLfdx
1Y00jqRnMHjkBpjUp9Xv75Gi/5NbnYUfp8UE8ZHuUgAYUSsDZBEdORt3mq72Lzyx/Ub5/ps6X/rX
9w6HDsGcQx1KqNP+97NaZovGXkoSTcOFTlgxjPRmT84FBwLOnrKPqM/bm4uffCufehiHuaf7lj5A
QukZQlUJhlxvTGtY5AqcOqHyTUyEl4Xs3zTbAVbDIQDd9GNur6fvP6SMU3MMrB4tzSrpU9jenXVA
VgfDYBLVFxJ8R7YblAeUrPa6g9CBZ235yVT/vhcE3o1qStcaH6M5Mg3xDXwyHgzsnygoiIsRqQUh
yQh0F1DDFahwChfzDMvgT1XRZIs0p9jU14vrOQ/gPZOzs1rCchbhSlnQMCFoTIHOArlhTcwoz0hH
1MszV5s/bzR47xGtavZLIPoEld1v/KdzBMvYOabXsntVxt1FGJV424XzBxwe65SlcFWoGZ3acWvP
FeTjl9tQRiqirvYXlrRJiBP1TwrQ3bpZL8QR9MaWylTnRWfxACquu3FKzWDD5rejCLO4q+oUcAZ3
ct5LftUJKqKsgDi45hHXHPJv6WstJY8iwFcOD98aHTvgDBbCvP8qZPXhxCL32p1/a5XSsovI2FaV
WXK/PBRT4dBCtuusTmNCHbxSvI7maYJMRXd/YZM3UX9I9osT3BJTjNDixWS51r2m/WeuuEqWjmxC
u8ho+B2MkWSaST0hJBy9epCW3xX7Z22hrxqTfyZqr0TWfqFPlh5tKqFB0tJLNgeScp/i/q5Gherf
bY8OzVSRjGNzKDWR5nhljUnGZrfFSO1Ljk2Hnswv1Qzx9r6s4yGzY0GvBbb6sEeQ5NOczPwKN20r
wV/VH3rKe3OGoeNWI6EV/2yZRwQbiXNndMeIJdMU6oDPvTDO7ukiuERc6g70STngZwcpVSyke80n
epnCmccnCFQmFuX773+Nq0UFptzq9h7OU77b7Dmj+AwWU4eckjc3Dd+4tf6CiP8hyViG7lHDrpva
nugj1ivf5mYR587uSUBU7njbeo9wtVX9SKKKWLBLr8GyhFAc6fjnLXO5gZa02CO+u4B7MtOL3pc8
NlL60XQNbMm4axJ+B+1Up/jjPUh2+n8G6DC0xao9hsz3k41u0uwtr5BlM3rDr9k9UfTj51mXdLLD
WQouR0K9S/ypJOa559LhJI4aTcM3huzyGtBiWtO28GhO0wKGCtkXkCN/89js2i3aUUxqM/5loug5
tikRUPUdkcvcbPwjcIVVzfsgN0UEXj64NqI6RPsg5XFzZDWY4KdybFsZDHQDoGGRXKIn1NdtYvFa
nSRZ2BZHBq2B8KR0MgPIqKieP1zf/RF2bRCv+Zdep5kBkFDAIZJmsEzr7uRQtLALUjJBUmA707F4
L9IYNbNjfFczIlgY/50/b4xzOOwZ5Z1vNsEnMw1XXbp4zMK9twyX8XxLvBX3QP3Posp3iqz+krxd
omBS0M0YqGILh0vr/rQJVZ0r+vkNOzbDyumVVl7vIT16tVn56jFHuKU+nDgJwrlTgEZ+w26E6kNJ
bcj2MYC9fQ+WhKI3vdG/+i1SO1JXZjVKHsW8sUqb6k/Y0CgDyAYEvnan1/OfjjJLDQzWEclRDLvi
rE80f6/cdiaMhXH03DIlBYF+/DDTBooX7ej46n2m2wEvFirRb4yiRPkZagBX0MUBZnBDqUUtJXL3
YChyzepm5keoUjEPY7U7F0SeWw7BNI1FJkTVlXA5NB8fHaw/kyQI3zEFOG9/B0OK3yGnl6xpF/vq
vuHYdswhzzmF2XceqRvelDTMuMGYYfPPyvGZ7KGtE5GBKnxaUBBYaUpPuZ1GuikqAxdqh0oeMcn0
XCfzOhZ/RboNv1ejKd3oWqAvrJ8L5or4pkhK9EJuSPujNxBqXrkbBXy9EGdv3QcJ2uGfoc0DdnYQ
OG7RCJvMNm+lpq0j1+xc3xbrCB8lY4xk2VwP+AC1kttHXdO2o9RrvOexC33jab1qFTE4CkeBcOOA
YeZtMrXuyZoy8xcjqsoDnfMhufjFi3HPkQXndTu40c21ZTGCDeDd57cUEP5vVYXThcYz+OBb32jr
L7flQrt09Mf09LObB2NQVu9PHCQRRduMFiPVaqFAsu0novp3W5kD0LvLhd/ApgmRZ7McGnRKPuHT
V/XL0AA5Xqix1+eiKT8T241qK1YC7BQuIvvtJdEFtE8hqB21SO01/ElLcoFOafRqrqPDALLLYGfo
muJb5WOyRbVlCY8E18EYQUHgus/jmkJ2KmRm+R+tNX3pCzUA4VgIrsWC6/hoVxZV2L7Rs2tGTpxy
61B60OT2NgHO4GNYjVTiTp2jdElSVzevwygdwc0d6gFAweuGOwAkCvTO6AmXREpYd7VEgz4ESN+l
shHezSkSnlrtynT9/T5zkZE4FfEh7UC6knEI8ZZOi85ZIGFYBZbo85nOAHOw1n8cWd3KsjeZhS2b
qOxRD7bKKqEQnMA4/jjtgBKwxABUU3qklt5FG00CwJXoTmL/vNw/wzBQZC7l6TS0Zs2ZNaC08bNN
YoEQ1omzoNB3nwezK96Ye8s7pusysSV0ZwCPMBRbaMg6x5htCJztZxL0XziYLw7EYcwS6+EkAT3A
IztwyphsMasZ+DbP+0NpGeTjkBkqxUsUGnv7VldY1ry6DE6o/edFjfiHTgqF7EpOPqWit2VHTpIr
MJVZGdIuHW6/c8J6eZYp+IrUpdgBgHCbLZ/3kMTaiShFgfluZj2AHEwxd7TOnlE3LyHaxZw4x0K4
KvmOUtOTiBRbWNCppp4CEB7f4hY6ADIvweu60son6cWBfePOnAkHLtBonkuS+ZbxZQdg5/GvEfbd
M+n2pU8wOHZQohwPiLLuzZ66p1ReyJKqwREomp6+5hHR3Io5fiBy02jeHcNlCwDxHV656RGK5fc1
2Zmb1dGoCpBmRCKvJSHFVwoAYcPtd9OBEdGniGZ8w8cRcfAP0KCZ7vCb67M0aMZo1kLYivqLrbF6
jXDVJ0MSpPtsj+fm1YK0nWp3X6uJ4UDXxedSiqXs7dOXGhFVE1Ppv6QDNqtEUP4gNXnpOXf9QFW7
dL1IetPB4XZkkOcsbOhbgHeoFhItEOGPN1Ysl79x1+lOdPQIXUcxuB5m04GwyxPWUjQRZNzgSSPa
lamRGwtOTGVeBFHO8KCsiVclKm3AL2s2II7H6ESMp4QARCnpq1I+0YPhOTqhI8DEtCsa+sRmx5kF
NlZreaumWWMUjmiyU6wX28vInZQ745ytcK5CSkPApaAaLrWMylbrAXAWiT9gtnHzh7sdHDPzMNnw
lyJ6wHwDXDrxdIo9HS99NQLTyK8UKUbFagf59GRNlKYOz+G7Im1ALPmgeDHfn/L4Wg0fvuB/l2oq
AaeMQ9riWmtVbZ1MgmsclzmAQxPesT+2iBbENYmRMWFR51gYaMWxULPNx1Ff8XZeGq2nhwRN9MB4
HP2k85N17t67on6HN28YSaZNju/E2ndgXVo4U9LoO589JEx2eQmbreqzEq7nwGhv5wHpVE89TNok
Y9yvdjI/EZNWF3fh1WKoHZrLh8A5bzmvW6UFS4fsf2ZPz9uL5AafmeO+iovioqSq18+IXVJfHsMe
CeCevmgs8Q7w655SnBnLvTxlY5JDIKUJHXECxgWg54qUcM4InfZIVfbBLIMX9m1LMP3lCE4hEyP4
7Rs/xHPld6qSkBkRE0vnXfP6+01yCijRFtaLBjOhIsyM8w0rCqLK9qaviYAH+ANKGvHcfK804FYO
3lkYs+GeW4Wn1VTZH3bxKewqfQPZrPaL5nY6eUyUfIj1/2t1pQt/Md1Rxk/zeb2z4402TwpjZT21
u4BXhVIe22GJw7S0weALMre6RYCQkJet3a1LU9xtu56438xHxoAIzTXLWZNbiPK5OUFeBN2rUfaG
xBDX6AgjVoyaM6iS/lwg61vvwx5m5hDG3iuXtwzvZMfFpfMD7m4JStrg62sFj4ZtLxa2cRwE7+SO
UfI1o9waVLcpST5Sm9wf8IgNznAoJhMNxxi82g1AQcwRTS2V5nzb65qF4PlavGS/Uj6PznVM40Ej
vKGiOt4oIMbyqBgTgDFnRe2buWrWj6LxomlCtYbpB92QNgoSrxG3rAt9vH85cWP+7AkDdnPqQANB
QPQvrRV2nzoZGN5X3e2fz/e/q0t+6PvViplEXmIxjaoBmfvegY36SaddzsnuM7yp6FL9ykOdL7lC
R302+/M3VDLAmFHzSG6by9qe5e9OwNOu1qNHUd5w6W4Xq3jaJWDNSFmpY+YPOQiza8QUQQIIhRh4
/aR5bV95oLiL4yj23M40o/jlx4e4Mlx/nMM1Ulh4LKPqDSNDqiGE7rQN7aFF8DAV1Lo4wVPOc59e
VQxXoc4zy3nIhKgRRxW6xGslXd8meXyNYMgYMRNr31iVnWBh9HdngshxW1MUsy66wztgUQEp/TmH
7argQfCzrhckRKB+w29sOjG0BjX5v16QQLGvh/XG9G85G1KnQn1IK7ddvCaidnzVkrCHLu4yCGYY
6mbjpbE1yWlI1hv519hiyjAvKALMwVOLCFvsHuMzDni7iQnSVwuIaeRkFQsQ9xhTR4fXRNUYvlYj
U589JKMIopg0DyhVjO3co394zTo6M6uBgY6rSdU+3xPRzhq/yKlckDbltDXhqlG0IRAQrCIF+sQM
5dS/gTxbS5zIOYcjz2ZYvpoMAxDSgpeR8+rsa0F3ZKhq9kGl+UGSWQgKvl6wAUqXEK/tqzhTjHBu
tzh0WIuwIR5EUO4w3UePODjg07LmyOXMY3tOzOgEBIJCvXOlQu4kQFVUBmqp0qxn3fdnEvyLSkcN
WLsWliyksaMtmt2veK90/zod2qnvxnwn9QPVveCLaekg0EMUMAAV33FuAq+z6sjzMbMUXf+WuwXV
M5qy4oqCl2Bj44msouUbrmiJ7nfFwZiS0ZJoPH6iRPjWhT05Qxn89wjIpWdLnW1CN8YdVnnIVc1M
hGzPMQ1+y22LwlstTsHDcaMtagtdFZkceTH0O6TGo91+UPE08MLVsXojHp4lAINbVHhMypzUQobG
lQj5LJ1qGVwDPz/26GsDyQU/k/zSntcENtobb9dQgC1MVL8vwq+9yy2kqaRArETqPLmytZFjJQ0H
BYUATNrhTsrhlZaVcu0aKIdikL+QBuYef7I/IGFdA7ZSLbnv2LH9hnRGpa4K6GXONBKWUvyACet2
JykQDwF/OlZBHApQIDNAEENCls+nkTaX7rtYxp6V0YC/CsXVQOIRs3I7Sld38rYjcq3I56rw64qH
zZbrthyDyCb0uXM4STR5nMmrWz8u7Lswnf7Hb/D0xD5TM3Ozf3e3+0V5bnsYE4j9dhOzZ5dRXOPq
T9yyvzgW7IIsJg+UfOWKnh309HTs4rjKFqV3F4wV0o9RUadXXL9GynmBO+fuNbDkYJC15/uFO+02
GiVac3h8FqAx2FEUrJz4m5PrC6UBIiBPvaqgaGAfwgHnFTN84RAY1tZ+vfn5s7SM+8ww+UgflUMY
+Y9PA9uQOOfYNlurAamv9y/wnz3ClBJPUYeAmlQaBPJa0xuhklp5erRFtTSNWlHVl9vMD8IAxuaB
KVXMmhjoo2rDWfnMJXkRkxTo2hYuIvVVeJCccu39t7YUdqZt7RtvQiibHyozHiUBNBULBA5OfCja
LL01wv5U/Rq1cgQ38nU2EFzKU0rOow0GHr9jkRxrDzu7xeKQlVzsF97fw2ugEZE1bICG1gN9bfW1
y3bo95ZglLKDhbuDWvXBCCMBnNSbkd8ZnXWAqoz2u+UEnrUXIh9kU+0B+fMKOjNOOJO5OSbrHuIZ
JYSitStFlLtUgFtnSwGGLhlvK6qs+cxnt2XhHsGQv6xBES2IWqFZZ9fulP81V+zIz/++dIzfh2BW
/kUWF53Ars6buiRpY+/sYCTOU4z9FCDfMsiIoMAE2eYYswEWHuZ/LerQ3Qzb1Td5i2RgBb8PjDDc
Yny9e47Kq47QjRNfwDlnSOSXYgMBMjZf996cm2CaF8WpUsK3dvqsDlTjYPS/tgIDLBi+TvVoix+I
FIZLv2dY0Fdxtg7qXRKJR1zazk7cw8h3+hi4xNACrGWIx+nH/ivLdcjsBf+Sq/3CzbpCCJ1ACp8p
rGUW/3TbHnZGGer7cou4eMmlW9URFAIlO1UAbRrkz33zPhWbAR8oWe9jgHG9KRviqaEK+PMoabPS
QjXXxWfHHMbCWMpX0pNpRwLNkm8C0B1uzCJ8mV0Y2MEQlg9eDqAy9KbbJjLPs3ThjctOi77HVXkA
7RY7zku9elrwSl2F5qnkzejpqH3w1DO+xbN0HT1THnCUd3OkbhU6GK6wXiIGLR5cG8n3hbJgnsUR
ze1cvyz60rnzeKOJbRTt0efM/eJU8OSFFwH3SEXHOsuKf3RQqsVx9BnahPnIzi/zM81x2X4aVUCT
pYLNL/ls7gr86s3iZ+yVSntSOEu7KnYJiblH+3NdIazKKH0THNDDh7uc9+9wLs3CoGciZtIo2CAE
I2vdhxLuOKEXKkcNjCCaRWxLf7fAMi5u0Un3nmRvSvRlWqa1BeJW0ATuXOhnh+9iP6267HrywHzi
5Tt2HdlcpCJ/FoFhzrHADv6b32YbD+kHt8VxI1nr4QTrzp/0F3PNry81PC/KMU6rQJtf1IjxJs3K
yGT5VNlkR0gcaVycROZ7Sq2eD3K7ptZ8VpjAGSfXvY7cgx8rjvAA55HKB0paBvdd5pGq3tEm3s8p
Kcz4gXYMPvcIMzmHjAEH5iZPfROQng0hZ/HmQ4kHfF+YsyB8RwwTxKBLkbwiu0l4UByxTJU5i2bt
GE/g6uv4XdPZXlVUR9YBxALU7uf4+9LKCFO6ZWAS1o1mL/LSw8Bv0+n2LSTS1lY4Fq4iadIJMvRE
qh3xdeTGhYADI35kmw6d6AaQTnjuoHNI9IssB86yVOsVY1NbqGrQGGWB+FwlVnWu/9cZv7rfraw4
yQC1ibMghNXh9KcRuok1iqzX2WoLOkpikMKJbB4usnRKymRz5nXhp66LiqxpRjSF5Je3pzv/4GSw
HHo2i6GtGQ/4KA52WZzpPo6+kS+RXjUsElIEPg7tyAgCHsYpyz7xSLA8KFEJY6/4wz4xuNSiIPX9
oGtPVhoxo5gp784UlvBWlSZyZ8hkvfF+weSWArJ6t/dBW+CiVSRO/DL7gn5aur6beRiCADIjTkbS
jqhCV7b2xyDLx1LQD8Tp1/rInTeNbvrV6wysuSaOkJM0rSEgX7d6zJq3onVYptVfy7A7149/nPvw
LWyuvZ5eJqJVt3crI2AW93qF6eg+ftlicix+3Cm3rfBLYlhgcRux1dGnxMljDQk73dTLc8SatTad
wyCE2DicEFVe0vITmqGFrFmCBMbRSrx5lHPhdOph6SOf23bcYK6C4cmg+x9m6eV8/YO/YTdNrx0O
zzycmnCRThh98i9VFcLxrth75nKUyujroTZyktL0DVFAu1hzYi/guRs9jJ375BxEokE9rLaSKN42
sq9YkoFF63aBOdD6Ndvhx8m60sztBqDmAHhxBxykhaiB9Jagh8FILiatjx5/dFI4xSh+1HUJMb3+
MqQChup/S8yUWGhztbtBowzSzsNFMcjNRAm0AAdI1enUMrdGvIP38QQyIulygM2rpUuMtNrAfiql
8gciVVrinUfGD3zQdHqzxDZGM99agAZ5Wd3x24L6HMtpfuBd4OajoeN6bvfODvPiR28bJwBUuQB9
ynuhgNM7vTP1ySyVy8r9Uxg5Mm5u6uluLUBfoSFiSkrFsF3vWjoo4FgeDFFAxEoabDh/pNJfCewr
GujRJpKIy8eKH5cukGAqds+HVoPgbx1eLTJPzV5cra6qm5BEDOQPKQMYIb1mnjBAI1Pezv3A+9Do
cjahp9czlfweIydMnfAFhVSJCc7VEN8wBvsPSPSLUwvygW2BPFodn6uqsdy4pi39fMrSavNfcaFJ
kzE9ktWQP4Yae+uvSbIitbGcPhhFqJAprC1cpHBZcU1y45ljAJqMsKrXztlheKiOOZJNYGWvN3J/
GjPwiZCdmPLz5yHGDb0kbUH8wU6VmSLcVQXeNErpIrvIdYqZeJgBPdLIitcCcMnKEuNXBg5dHx3v
Z37c0GDWyFb+lMWOye/fFxnUGRX2NoslbQlRLN1NIvbUm7S8kG5C6zOxF2s4buHTtzbpQZaxtnuw
4tqKUVIzOU9pd1OYBNTDzsgTZFA+7jKFVEj1TagJC/BUIaG0OHqd4HheHqpp0yPBOxO0YPz1ifwr
NmOtSdKpKB/Cc1Srvwz2PzdU5kAI/SWSYwnw7QIfci++x22Kgyba88bbmEXAmW5pYmV/aog9LPh2
T7i3lQQB+hh0MyXsms4ja6rXNl5eVf27GFQRQ+AAgL02L94hZS66nAi6TBjxY2L3xxTykKvmEngf
WMxd3tG0toQ5az8wWO654JcPnHNJX+Y1qp4ovmy68T63Yw3myfIPlY48brLMcE0e8qTlTOOXZO5D
Q+Pq+DsB3lesBwIx6nkgdFrpInNgLpVFhU1IyLDOqq5elnNAPxX6DLacIeEZOfHYNTPIcCRfWauZ
XcfT/SzLiuPwHprPR2/Z3OyvCTLoqz7+9ZllZ7SFqqDRztBzzJZv8XSdAnwcF0G+GfWKfzDqrjaF
oJfqmVPCmzUonIzzWqpRp3jJ/MqPrAzOa3GNzhTAu8MWEBW5vSsVbzu+OOy21SB+W1JPzf+L4EVy
3FETfMPEqa2ElYuWewBXW+NhXvCbkfnydBqUe57xEY9XqmoSlDuMwPQDfEx3lYe4R32jYHVVh4jg
PKBu7f6bLe7JJurmPMyo1zLerdk0WutMiSp7vYxiWIf6cuIvw5e50PsgBQK+PIn/vW1oEDWnRzW8
LqUG2h1Fj7J9N0Ik9yrP0T4ao7nI5a4Bsu/yI/TheC+PwlE9Z1MTtsAkUeDcBTN95zXbtPi5au/j
0EvCxyYaV3X6vIvq2h1sUt0TycZV0FpRgxcsW/lVppgfhBFSXeLgtXGbIa1iAPkItPshSxDoalKY
rKNI+VWrGHd1OMvWHwIuGgAprLlue7zN+PEjBSP3J3so3atckSIZrPMqU8RbESqimF6L1eDiwT08
96GVeiA49uvNmSRZCx87Jfprd3JHE2qoKev44VFPodO+/2iNdgqhvOqwOA7lbc1O/XmrQWj1KNUA
+7pB+gbzHLFQGMF54pVtfbkE7PMX2hnjUjMAUCquqdBOwivVuySfZxR4UgnLzrSZigsGN7Jj+pHq
1+SH29GZC5SCHMfJ/dnacu2AzB7ZgBgjnb6bzK9KUMT+xbvvhBMxOa4iYQa2vn7gsjJfnY+EbYN/
hOW3AySI9ja7zs6a/eWKAnLwxdrGLt8jcM0ao0yMwo+XRB33eEWqDenP0FWkEQ1oSv1Zioe0f8kq
UdHaz/wZ6sTXCnJs7rmTAXYiolKvK2acyC+QimnbCYHwUo8gJ+ppWSqio/cuHLgRRs8AAQknE6W+
wsmTvVwrbe0GcYcOr9/eFfFw47fBTqfyqTf06NyhDxUpn8hXyAJi1/Celssmfw3i8w91r/ztGkmp
9SfC3Ra9p3+CSwmk0sCrKlUfLz9v0C/8V1c2eqhPUICl8wx63/5pQkkT/qY568c8iLUYHnSpMUJ7
/8TgBBkSLa+4HEDtU4Am24NOd4RNsEXiwsKTuLHK1fu8veUCxkkZegsXfEZMRB9c9yZ7zu99t4ic
ISdxg1d3TNlUMi9jnV9SQf9DQmvuxl+3V8tzk1B3dUSXjUy0YwnySlpcQafJ9CuBrPtZPRAIfs/T
PszQCuPpE+eBFFfd1bDFLYhcuKfqSH8PSXe8QqyBrQbSobzLy+nZ9Nx7RS/f8n58jVv/ONzxHq0H
GL8IOsnr8o6hAVHRnsf6mW4CPwKzP1eA/q3u4qQoNe1sFJJ5XMDRMgqycSrWZyIHQ0YxFt8w6OA1
mMDTZFDbwoa0gLMvRvY6NFj4y7zdqJmrjz5D5Z/fkWYzbmjUDL4n/gpUEFHhU3fO0ZeU0QxPiCWZ
i8iQ/0NFLWy/+G25ybFZCv1yXsW3tbIXGkwbL/y/Xwk0EI7FxIt9h4HK4C/Ot5+Q25Pnv+SgyqwE
ZhBFU0uZHudawzXLcuaPP6JD70WmH2lVWeJWt30ywoBDiBfzdFhYrv+sVo/ZNgoABH4CSMR0o9Kt
5/xvNcNKneRv+8vf3tzb3nhk2Xw4U1ynEMJpKPtvzs1Yy0ShDhtg9nX+20BgS2VpxSUJ+nrqNZ4P
jiPZKHfP7MMat+MG6ksptr/ZTy0TZuCVyWC4U0GVcR9InqbZooCulvJvlmSV5vIAOKbggqnjzQAO
LYR/J9zQ5v3A++owa9hcdrxZQ9/w+qDiID1AecQMRh3mi/a2mfn38Sy6aVyPLyvcUGwqccS3SxGy
tbwgE7nohgF9KO0t+2hCiN2pvrVSklsID2TKEahj93poN4zXiulrkLTJxe8czJGra81DY81Q1GMN
MZkqZ9BTsepn9avNmm7LkMyEp3e5Cj4LWXpuoRNH9FcHisivXauqNwrCLW9zAAs1DUZgA/UPRnpb
xj5GIRPRLRxbMdIPOT65wSMWpG4/OzOk/SUV4+l/CHHVrLAMiA8qAju5ifbALclyfUZ63itZxGWM
eFVuhdBMiSsLdCRnAzkGOclZJwC8e+ahGlDze1ejmd9me1q+IH0A/RnP5o53QxdhGvjtx19IAiq+
fxFJLeUPPR3eMl3K7+cMLw/YXCxz8GMsoYY3r5Yf50fWQkextSTxBipgD0cDcxwo2BlX+kSzdy9n
MFqQ9p0VwFRT6zLk/6LJ6n0MO7l1eM/oLxfHrii6USnzN2Gs8CcghOBWBsINOKHJh8vvTJC7fWL5
LAsHYL8hG8r1N49+Aaig+KRpAqQLTgU0qHrDeTG69eaT2huK2tdjs3my3AwglSrNzyJ5vCR8PjRb
/PYGKsPX1U4fjjNmM4N/RBBCHTxRd+a8kphrppfm7Qfw4WUjl8KnAfqE9C7gHWTA71XXagbfdWci
z5gBX04Aau7JrVMoq/+0B9TYW/xdYOeEiEO005GRUVBcZjXy2zN9lXG2i9is7JndxCMLn7KZPXnl
jiK3sgAN+JzxMtQ8R192UahiZpAcLDMDTdfp/8z8omDhC7LspjFonMb76ggqFdjb+uh8Ptj+0Td9
FwOh504EU8P+oRHkKrZ3hWsWIxEVnXFstBlEsow19yO9EfTFB6XwWBbDyeyQp0hvAK3MITQfZkqi
j1xbgK/sVICnkNPdoNyFl49tUWtyMMm9oMhavd3Qc15+NmA+Rb972QE5gBwO9V8pZ/NvKlFncla+
vhXTBIcKDne6f9helT4JhmYh4632y0brvIww1XiHyji2nTn8u/VN4H+sUXg/4MCmq8pr5ZDBZRd+
6fWyWfrz1U7jdXMOoO4CqbF7m7A8asWTi222RXaIBptpzQO/EvpMKMVGj7hWk+SSqbT0I3YBh74C
P1IAPCekxsrygnsV4MEQH+m8l2UL0GTQcQ6cViyWi8UuTg8axwK/Crkdw2aoerdDXn63JI1e7zW5
acs4EInGD1jrpJmG1AOvMF1M7gBLhWPXS5Fu4f0GkivBEDo2edaOEfrV+HBR8tonAcjKMNpmgkyP
Au5RdOyQvGBGpCKUIgZbd6KteCtuTfWBlN2w+cnWTGj5515bVfoc25RXmg3H+lTRPGFHvB79bAdJ
005ytOF+lPCbeU6dGuaXWoJJsrB8uVvvRkdXhbSZA4qPvD0oJS5X/iD9zgAOtlV2NKqcZewtuD71
QBWwQddCIazYwNtKjUI0tL0YifiTUWsfQbhLemfPsmITyoWMtrIHvfeCOkjix1SrGB0TOgjxf+6k
UwGpsiqrWwUpLVffzzeQO9UfJlVMdXksbBorRsmX9qvdXm1z6H5swckKjgWDWiI7mHIC+YOA3NfJ
DYSuT41JxHuW99Mn9zsQYztpQcqIiZe3oqs2U1UBQfEbWLRIDxlnqzkTt1CpAF3neimYq1WlCaIW
SqNfgOXsVx7fay4C/nNXb/bNGfU4U8Uv6XyDdIoLawgkxbNWBYbihn5V3+40tP0JlcQt1p6ELq0i
/xPD9mBk+ZTkzBcR+0zsgoy++oNY18o6RllM2ogXNYqUOmNJw5iYKVyxZOMESvncHzdXiH++deXC
UdRly8M8QVyfLgHYm1EtR3EpKbhGYeLYxXVhyE/S2T9DTLsqUnMdrgGL0I/4Jg6LP1Mfp389pO+N
SCwb27a2xgXHP+kSWVmBEo4B23Idl5dryT/gGeOauauNisQt+tPGzAwaAdvphGeSmZ4ToqWGIPb4
INdVY5D8AJvg5aCu0TVacsPEmZ8xEyhdLl0L7Ni2S7S1KhAiiVvTz2jQYYJHCu/BAz6O/D+ZcU6u
kdSjXMod8+iCFI0sUS3lzsC7HFy3ZyA6bt52QJHg2viBfBVb+iYqtJ93KdOpUYFZqMB96zzjTRqI
w/kNutpUvOb7VJYPqbCiU+E0nSjeFSYTdDKls7ZLMa4t4fJH3H9kltCjvYe2+OHOUaILkiOsZEir
923m1+cgfqf4fxYCXNOYbSO+QzdO48AR62w88zzOZfuqp4MVATFn+cFfPgtAIXBaqy6lgYqTR2qF
Ke1VlJpm+5fAberTm0P0L1jEk2r/qniNBlFjk8L6bjYfmry9BfwzBhSTYtVMJJI45i/B1im/VjOp
gwQY9YRiCCQJys1u2R7meki199Irq7DCJZu/9L8BetyCOlOHteGNDDe8+ejYhSRsrz2Nb3PIH70H
+IVq6dEBx6+cEnr5nU19lDGv9g6Qe6JyKEo1hykSbs3B2x6ICHPsrXCLXDaNsNhs/ixnttH2GThy
rKSI5D+KYYhms8h6Gwxh2PmplqoWBf/O3izoKwypB6b1SMA6Jskf0aXvS9BZk22W3romz/6ya6VU
j9spLnHfg1q4WV2/B4x3A9Q7IylvkjVtKzRZCU7NlMLDtDQffVvfNZbRrXTLoDxkFVPUmnKxaEss
h+/lO2RaN3DDLo8qhdl22wDr3mpuu0+SPkzwU0wPPrK0NNyWpF38zw2Xv1tMk6l0EMdmIlfgAEHX
niFAnjG3uh+uxdNveJSbWyYzkrXds3a/TrNWmlfhliTujpzdXf3CbEYZl/HAttUUolPtsdbUoB2J
UsUOd0PAUYH2Jp25AGKR2LTIVkG66O3/Wt5XDZPM0I19DKP3d52dBMCFBOaEkZxVIzx6PtkdJGCi
8rbiWBwraf5i2aqWO/q95qNnkwX4WD+ooyO2rZjhaBWP2WaXNvqpF6sXaaYTkrnvyNnz3xTngg1x
QAMHbXq52lFmJcVDTTwFuXRJsfD01+BJTVI6W1kCilTmCGXLyrHQX7XRvF+nshah98U3TG0hKFqL
mdynZ39bOGNAPzkhMDB14xTXlDBuu1m8J+y+ta2/X6KCNWtENiBN4rRbbZYeZ0Rn1pjPblnkIIZo
23GhY0zqEWdZEdYpZXgPc3z8gTrOlWS+o5L1wJT26yysQJU+IwKWZxD6BGzmbvLSrgZN8cK6hVi2
cfRabUtR3n7VwfWgxyTSqnXzCv/ksp1dFjrGpqDjbEu2b3eiMX+KUllr6N3/VmUVPoZkjqObeZkh
8JIBxguNibB6cADG3eqfaphacvdPKcn0RrfYnZpsouZsA/3Wa3/Iwgr5c3nXYJ1YUyzkOJNbagoz
8OPtJJUqIrZEiwAmDgsCjSk2EKc/Ig+wIYlS781cQUXBBmArIN0GuBLErNSW/Ck4NoYKnshXPKov
AQgOlmI5f49eUMZT93xjka+qmMq2dsYyBl1G7SLhYMb7zkPk6Bxdlt3lOQKPN/Lz6uwINf9sL+jP
eMvioSzRuxnWrCpskavCKc37dgfujPL1SHQzSco7cnvXPH/pkJf/tiVB3B2aRNc78zq61VhF1yL3
01lWN953fq30AI27RXFcNq+nkB67yTyAMKqwkPGdukCaKyloxXblXSA0UzYm/n92UKG3/Xwmfds5
NcQm7fwOvoQi5yQai3bD1Q+CvZa9E715mhiO38OfbdY/s7PwMSkqSgb8e+zT92mDUiU4K6MXUB0+
DO5QSpFTIoWuxNVi7tRUynevcGiemNn9beIcAVxpEo3Y0LVXhRoFtoqgSvusN0V36a5CMdD2urDI
ydkSEwlkfHQQvVAYdutAlyxZ1BFpLH7SVmi92+KaJl0ZdZlZuRjxoc8SlPK5uF2RnjfrbmvHCd7E
4gFHWwjUKcDbA2+s0AGptpwJnHM2XC/exMni8IVuZSMkxTG4Js8rp7tGlFx6IbqSbVm0Yo2TsTT5
vvTB7SrM6fN1bEyQ50oVLEWOOMlhZyebIDCM137Q3cjarr4rJWSS7QYYV2k36juZgkzzb08KmXoq
lpEsQ8TCdCnrrpD4QFdIhWmvPpG7yXG/tYfDwLVkul0Sd3zDie/iUI6tImSzRRH2k0teItclicdE
KdohCD1sZuk2Z4Y8v7sKXFWFrJzglDnVYzM6rYoKgPDq0qgh8T5GMvV9b9JynyXczeKJcEWWAV3M
+t59USlZbE8gEhKFzbtfXBdpGv6Z1/+uf4A6Z6h6LUjB0KMEQverVTITFtx3vF518qyfSilU8UaD
CtCKq/9ZPpbsG1fuTfDxkQg0PAmAKkTqW0nMIJ0AGg5kok93rPG2v7bF1jylMHxEh7n49UUUvQLS
tfxyRbE4mz4kmqFZD1Zcc1pXlkPplW+4VTa24PT8rN6RL7yUthLP/ZVBEr3TP4eNNzZhxbKLzxLc
Oz/+rWoDcOU4ZtpQluGB8DV+YRrP/NM0FeQR1SCMAThKhpEahCC/YVWwCxXzkkiM7EjMH3vwMm07
w2tVoKnG/PFOT64gkQ65OzoSfoneOJLThrITyMcpAE90LELsxTbYjEP8Q4YxWJdDMRW4bWj+TurF
n04pee3aqKNZul7wxuG/Mt1Lp0q9lTNqWonMxa4LXKMJ37KPg3Iu2Uf4FfiX+GgQ70Qvhudl/Hsv
G4ycOCBeQD6K8oxLfG4zrdnSrDGxSL9VM4J0iObXDsioQDvoRX+HxztNGcGxvWYx8Iy3a9MehoE5
iOy4Xbl840RISAKpOAM09L3iRlSZNjSritVFi9CdBAhGDIdDvFf5K314aNowuHkvETOY+mj6mevH
YjTUfYw5WocgV3Ts01BAyba4eixVpG4IWxS1EHZxvs6oS/Xexu8enIEivtOCG5OyO2Ad9t1CSkxp
IGBjlLsToplpFU7S4rUL4Z8AqOeZt6h/l5MGEdr1eoauSjFQVf6GOc/icVxlhxg4zLbM70saIOAo
6Q1AiWxVD6DaT7lZRAkb5A8jx/e2XVNZee7Hz9bvCZs0VBEDr6ms5qNSIFbjho131wtU0WYsUlkv
DWOmJY5DDO1E5RQeVAgXEfbHq2MlOQoh7g6j9W9cGMd5wJd+Ut4xmq13M/rgB9B63csfERX5kruH
qw0JhFPCZaB7mk2WDTuOGTH3clazN880WYk8dFyepZz3Mkp+UpFZQPaFJCPagswEPj4WInxd+EFV
YayQgq9NnMdNmsyVabBfTyT1RTTV+ELXFM2hHtXrCdAhoI2jVAMqJhoeHiTxc44Pq7XUm9/jhay4
KMuDScKdEnGe4uYOUzQomdeqbOTgBzsf3Aio76b2jcXqKeiaKEsIyrfi3pvWuN0JJjjIKCztx+Km
zBMzCV6PnLzZO93VoTj2vX4O3t2I7SmB/s7TPJwG2nvNZ627H15BKNDYzjMmNvkBHY86/XaRJbvi
A2nFiRr2y9LO5SxsL/n9MTwjKHgAgBCPipZ42Vm0JqSEoQC/GHKr213TGYFdjfpZinJX2Sopc/9D
O+Kii8Wxr1p7hzFu6AVLdKGVtrEGaC1D1niSX9SoKZ58eShQd1AACr0Nc84AcgUhhye7S5kw5KX1
ga/uVALsWd2lsoOozE3KxCQ38Bv/sHplN0+DKhK5ICHmeEktYJFeWD7cwBM2o61D3YZJHvELi8Eq
kW/ZYB8D40vWkbi+3+ojaZJ6/AcMOhEGQawftnxFATR1QMTRkt4bgKlsoFlduMdMR+Jjja0o7FmQ
qX0ciIlQdCMcFi86+7tNNTwozCbIN7HbCR6LC0jTfc4yXR3UgNyhlCndXBk6QOea5KM1aOJhjuG5
zHLlH8VnFK3JVwwcxVyRtr8CRYUohRFyubli0M6WSa0r6haJJidICWfeI97s10wBQvZHQKjMfsY/
L4qBmqdoJOnHwS08DeMmpeW0v7nhe/QMuPvkmHotXuo8Q6J1AY6lNxbLY7aJL0aPJ3+RAyoMTJpj
8V4lsMWAVe7wsOzzh6goBMIsA4lu3RIlrAg+YMCmCwvI5g0xb6hOvRqQb97b9H6jnuwvyeCRNGjf
9QjVLzyWrYrsWoYuE8BvV9o987f/sK5rXZUiw4UPZwRT4ZlWzrkLnx0myoS72HIwnxAVFNBx2Q/N
g2NQRzDVq7FHc231ooMdUjAwKWJvh+DuJJJj5+pB6TUWa6O5rLch043O+pC1N6n+UsXBTYHg6cBD
ouNGRN+Rx4PJkKzECGG5LHP6zwhBn8u/4ZHtiIC8dM9hvD29yefgMc+p1SvNI8qXxgdBcg8zVzSe
lVn90ct/kSiyUviAy5dvfAoMinjBo1nOsbjBHbKdevA5TqHXOkA5aPr+NucD8K8WvKmG19s5QsyL
xG7wIin/VH5gVC1HPqLPDuMYcBuemXUSoP8CMndlxHLhnLUic11ZvSjDhxbxwlh+20V4Zfa6XelS
0JlChRIG8T+5MBz1WLpp15ji2c+DLtV0y7RNCUFiGaeOZvIAhqqy0qR5X6gtI2jp4KWKDvxYFL5F
ARfWYTsJL4UdQHfMcW2AP1xF0LqmLYfRGsop1aXJwO6KJLy7IaWeBDHModTsm0acK0QZIOtXqcet
Z4Ij5NqUrSozNwjnQfD9zaSsz4LnCOF3ZqBYQz2wIADT2wris+j5v7fIsAeffOXivAaQi4/pHKag
NeMMJ1mrhAYynZL7JXwrRNczHzA+vERZfY59rzz1xNcglJhl+6rsCDO7sVC3oZSOPomxQnZQC8xA
irQB8u7AXTWhrVq2Lrsc/FdOBqTjuc16LVQTTDfrAYeopUaN/1rkKp5iaZ63PUEwreyyB6VmmS2O
58lRlVgKSdZQJBDbWdNmOk2FHR98etRm1/OmVLH5jSlwAL7gN+xG36kaEeR2T0EIgut+kQwEVj+W
UzAopHPH0fUMiRNO9gUIxXQPIsqgqQbFpCVXVHlq4tYrdfr2P9uZXSLW2kJnm/Frlx21U7OQi++t
1JXDOhnTKA69Kx2CgvmmZBDsdKzLWfgfRPiwGxA3qkYsCKzn1/y6O6vf3x4ZrBOThoOIVAv7xB/K
cOzuvr6MYG48CS5nFL+OY9boZaJSHmWRtERKUY+P1d1XdnS+Ncu5d561axmXIr32UPhHWeaKhc0r
KIEH8Dtdv5GpdBTNrjs1K4pPTRnXhv0q2VEI230izMB5TuzykQYWdgQ79FnyaELQbSFLGDp29B0h
WyNCi3u49nSGOf1eJhBK4bU6NZa40jPnat++oFtuwO+Zmdt89N3YPiWxiEB6HaY73PmK+HjJ+oF1
kPXuiuIqRJ40MU0Fbailej+yVmEubLWN3drtmFLP7qre5OqbVv7RrIVyEwL1Glqeb2Zr5oNjo13A
dLJMFrQL34TEcA/YFEX5plFeZc6dnBoPRrsD4aNea3iAdkL9760mnje5kRAcaL/fhiFUdzJspjmu
HGWjyzs0s06jHPXMQEawMkrehjdYBEs1UltjLf6objcMlmML2763E8Og50qFeWekNaN6Wutx946b
FMbEBwYAsH5QdVsPLIHGtNxYY7o2XA0KmpMVrVMPRoZ5NJx1jIwzgisjF82waQWQGh42vbpxwQjo
5HG2rwLig39z+cmOJ5vKQnXd4M62ogOqmG/13KGT0BAeM/AoUty6cYut0qfV5THq82rz+BoKq3hk
CtUo3XA/CgbfLXtdM2824zOZndaGR9HFWvUbBQlF/j9FOnUnI/n+qv+OqpjkruzUdk3gFUeCqfMO
2wDRZE94SYCuE4YWqd31/XR5GVXSdqKO6ktekx26sCs7ZZJtNKLZXknXhqhiSfmID1oloBEDZWWY
AdnB6mviPAADuNYgaJ+pnhAKjgrU3R4/54FmxdU08YqqDh9mugjH+UkAl9gUvI+xj7QmnWg/FedF
nKitR3MvqjcIN+wReRLP8iC6y7GZP6nftTJ9lBt7N+/NFQ4bNIznos/W9htvM0d4R26SCerH5FUj
iYSqhFl5WZwcGpfAwUsPynE8nLicNUUae9a0smyNz84F0DOuO6Q5mfmI8w11z/YJtraqRlzux5fA
FxWM4yyfN0REYwkxz21HGHKgJhy2cZXkVn9BAvDU/mJn5HLOZ87S/v9gHXA1mVI6xd+R3uvQ3NRe
MeY7fPHZr5D+U9bg+Luw17dAxKjMvl4eX+BScTUyMeXw45md7OraI2F/8+ynfjJ0if7/yKxJublj
2xgfZyBX05uZE2rFFFI48Y4c+3TmNXWG9DQSPvGjkul8WqeQStZMLVEPuEu6gFX2d5sc4w+CbOjP
6RutuU0SCwrOhsAolrvjN2pGJ4wasHXA72aJOMpBxAtHp/tGqdjIv4usCIhfKA3m79YKvhjQmw6M
ahRsrGdFhsgrw4sRoz5KTSpNiWf0EFPLbVaJEUaamZ/VyljT1SLsqPVe8sb6NgPq50pLLD1ISVZa
b6WV6uVq+lo56fJvpuiAF6uTWte7YdE9Bj36MIIoNcZX2eVHASXxkaLSX0kZA8T6N+8RUUDHBCb+
2RLUEaENADvgqs/uJxcERGTtzl004l5SdsX5cbD3tUn58JonP8pcCDMh9V0GSElYOnU0ENV62q9i
cgJRgKgYiw4NLxP2H+x0iuICv8aFB+8EJv4XCWgAyWpL1WVEsNzOjbMfCydjA9G+iG6myZcH1kh6
EQKCmjF0t1of1b99g+dSUZDLPAOf+mT9RVFknQ846uRXxrR/QwKjQMwB1jUXeKJZlUZzBauZxCQ0
r2Ux/y4sXCsjkYdfPg48dWplsxLxEsOrCPlB/7t+0AjBZRvsZkMwEVvkTJGEYqR4q3Z5tKK82qNZ
ENJJAFouw/LgTqMnvU3LcXyJwobuyWY4i4UIGX38HqmCiML/j+dhoRPKehCw79d9kQkTwpxfa2Wa
FTNWl+bf8iOgPXiSD35xoPaDjEadde6uYWwgZgDZ1mzNJ6czmwAwtSfmi0esYguKUrn8Q0mIfIPR
SetQVcG6hJIyEVNU10XcHFMTKN1K7lzQxudU9Qu8959s++wvVor++EYKbrRdTcrXNpslDmtRuZrC
yNMquQdKDdb6ZgL6mwcmjYTJ3EIYvjVwPJmlXwrVum7NXJq+F0j0gtuVUcIeIa1Ba3ipAQ3qdKl8
nf9SuPzTPb8+CYRDvDy2OiZVl5CSQMbQzpAMYkrPbIJ7PpPXmcYjRCN/zbhtV6oUJjsdOOxqgI+L
0fPWZShU+T03WxMlnVaI+fCFyrX/4pAbAZ1UVsK246A1ndqC09akER3DJhVca9/ZaO2whoVN2NUU
pB2XxihYk1NWAPfn+lHembOQdGrDSVBRyBDLFmhQDJ7erOqqc4HsaKk5GoTvpy0sj3aYZQb0Yi+m
XrKP1ABlKw8doWAWpcXjCbIxG5FVvZkH7gKiooJcxak60tTl0d9vdnyl4PRdECrf4oVHVrS6MdSQ
VgzkPkPPjdp4mGnUQPhrc6nbc0YuNdnr80eVJQLE9Up2QissItU5mcfw6vvIyc+mt1kfrXgZoMRU
P7RKZqxoxOQtD6UJlaE2evR+kEuCgwDCRyOMR44K7XQGxK6vhiRu6JYbxLp8DERhWTCQvNiOB6ai
hBQ87ao198wsJ5f701zAO3IY0zbW4t3XA+Pb1P6n/wNnYD1ph46Z/k4KMGJetdOrO0kwsBsrbcIM
WZFjnwBjpmaRPykGNCFkkZ69+kCTrpAt6XJkZDVe/NX+xqmYnEDT04CDlm36FCUOz8us5Dbli6Ad
LizTIRTTM1Yq/GfeoZ+06dpCpnaEjdmbRPAa1PBwtIGoi3qOcPsK8Ax3fAVwVcs2YgbcE4zTFPh3
eYqefYf6XUbBKgdcacgIjW7bNcAqCGz9bUtNfBXDCbqxelnIcSKuDWBz0b9BcTHekpMfSzNzIXpm
E/4WPcxLl+TyJR8xgVJcsNuPy80WgdqCwIyX804IwHqDu2TiE/Zky+USgIpm2yw2sqEOvhgQPCE8
gaaDijd6yLmgLDeO/sMLn93rOLMze+GXI42KDlr76Py4tYhHaM2w0wjCp8uIr6hHSLnVUnekCIkK
N3/q3QBXynVeFCFV+vgCcXY0Eg3AAD0/q1xLeas3n+ZDiK89mk2iYFrri8Y6fE73Wie7aVdOrxJZ
EZBUQwrTSqUSr5fIMCT8/W9MpBLg6wW5wTazpJMPOHgkTqcTOZRHFJLRzu6gw2fzCydKn+244C1c
K2yCAB7eRo2q5oKT8x6Kmjfa38Pjpn5iO0jllUUHNakt+I/D4v0d3N0rumrBs8N5J2S/VBHdsSDE
7dMlLEPUXrlvzXG9XmbnVDCD0RwrbRFMEgh3cPYN1PwRa1MRR95LKOvbwOIyLSozf+hl5UXAJ6AO
V0xkOvcNnklPqseHQ7in5p5+ql4J8bCqnIMZCJd54AfUSeTmgdWxPqVgdVUKI/FVHyCxQ5G22txN
NnHE+ENVFvFf2pqalEULZkozIFlF6xFeau5t4zwjAXYRIxhT0hYH/mB37jtdiHK8sscYxNt7SauL
WHtxkqBFqyapCZW8s61bmuag//6CdepjzrP3IB/WQJONpnWhwIYNEkBPbeUfs5IwjyAkuIWth7bE
wMzjW4+jfSdyad4UfUTuP4iEnT9DRjshqp4+kGOSnJKSPSC24myHZKefZtphS6mVOv/cvibuh2G+
Ar9ZsCh4K5TygBCRodqgrXRucuKpGhQ0yuWqmTj5GHylkdJRlJADlbiFoNXecrtu/kzksnFdrpvO
8f2qGfMkBnEfcivOyb7QEc+SVgXIKqR8yPa+aDncJ+RKoE8rsATjW61Sq0elaDBUyS2rHgyAyBk7
82jpojPvOdO00JDEG6/vi65NLqEmQHIgmarvlrA1D5hNKT6/vIxDi2GHOhji0UcJbSKy5s6CfEX0
QGDNn3qLHnjDT5RM3/fYdq/mgSrGZVLLWdG6KeLezVxY8u390igd4DKLCAHwEAc/yshc8uORzyiA
3YczOD9Jen4Ol3/8164zYarAWkGt+SP7bHDYOX/xFBtRUVuGVorOiR5Bgtf+d4GlUk6cnPhh8cST
x/wlndJ8AyDhvJmXPWI5pEsarSppLE9RVmLLU5Mn9DNi4oXU+irNNUInfRAOsSbuoNR3TwNYcnSA
R0ubIrIE/5A0okNfkVEqBJZjXUdpEIdxzDCcQcsRJiMPYaXndpdI42aRi+BAYx0xChv8x6+N4vXH
4CbfjN1JgrZxCABQX+8wNamX+dRzb5wCgwQNQTpKZnFcGe7y7BduxSzQY6e9SvM9Fva2e8Dli3Kz
RVGvYq7S5yPSV9zj4241Xnr3hZ2p4qS7S5QtWMg2kqMCGzz5IWbrW9PDXOO+SP1lTg3gdXGPm7KI
m4t+T8y2WXG90tc9mZdV6bOTfBXcr9BGteQtP2C92Ah4LAzQbrP0nHEVif1clnSFc2oHrghY8fFH
25VlxXXMW+f3/kWV+imih8U5+mrgg/1L/88t+IGGU2xIG6TSGVGFBQ7vwEjj13WJtfYZq/9l60th
3HH2zT9jpdgvxN75WpipjNIsureGL3rwIJ90YdUreyv6nJCVkCQvSIiZHFYEIAI7gEDmqxfNCH07
gSE+/kwHHK+YOYRi7MBHWymJoKnsZT+LvbUNtB31G1hwIUqIR6fphJrMx4A+L5tf7DtaCWyaasQN
GrrAlLF6o143g+PjNLcH4TdqwEmGmrhW3YDQWrWmlsVTiKss+D1rmGOSCrMnICpemDOJnYd6MC56
hIZxcdoWSS4pWIeCQVqgvTXgnU6su3NOQFg2tZmJv3xtDjS80s5l/18QWV7r3E+0/bJWVagpfmu1
j4rbzzJfXGLrA8XNJ4tRhNW3V0gmhRTIJ1oCV7BwMtpl/ZDs3OEBQmvEAOsFKwf9Q2VO/8dW6dMr
1zr4D3np3MLpLEZoXH8TFNhuY7xZ8Vu5zqKYEpSjd1Q3F6cTmKoi5Y6nl6ECR+rJR0/UpL3XxZeY
jrsNv/ZuH2TO2IiBzMOfaY1a8ujThliKsci4BDO8L7yCf2NFor67it+VI0Cu1GBPIaGv+TLj5nsb
kobzkxCAwcxLSvtcnZOAZNiJAnjU3J4dLZsAQF5Fyj02oz8MlU7G/kL8HRpUOqW39fDxlRNrkAPn
i+8Sz6RwReV5E2j9Qht8JuUXFgxlvBMQWZ8Tn8jtRayha+5tKXAJlLXKUJcn/u0jj8YL3iMCs0BW
2orx70sWfVjrM3Inu9BBvu1aHe1vNg+2oXF6XoqKXK7tNgaXsteAdvNrXtSKwV/sO8fkbon2tOpO
5YeIfbothjWBLpYiYyez8k8GbJbUVGSFOzEPjlF2j/pRXB5OTB2DT/fgnh1epjdfwOSH8+7PUJCd
6uY54afJnkD9MQXVgioqCpJoqIldFGBmN8vrF638AQNXLkqjhsSBmzwrIAjM35qJINhBAzSDCPkz
UEIkjYyGaScMo0wesmBl8zeSsPKyOi+g1I+EBhqkMGk5d87nXAiIlrgCK6j+YM63e92UpkOEOdP5
+NebgSDg75ERPcBvBPiG7Tx2eFZgpQ1kyeLhefdPFRWX82pIb/sKi+JK2xAA5FZMZDfVw70hvFWl
qCn1QMrhJ5aGMzFOIDG4cmZmCrvXiP/ZCQ2l6h7akRdJYypLvJwJvqjj4/tclZ3hFPwYrQVZoqhm
Rjvp/7EIoT4AnfKstltxR/1VinmOWOEjOnr70dq3dw0GgfIxcrB/VGnz4CMUrR+qAFImLRJcA2oR
XPM9PV8Va81OB/oh3Qr+hsug3IiR7WXVDHyBEIankL/I56plFuJwWoGU9YHL4k3HEk3tSnE8ldop
oAwg7iFhaSTRC9NixvROV7ycB8Iw/jceQkOLEztjZDYeNgv7wDPldeTVBR6GDHzPGaqi0jOkgsIA
Yx7PkSBjP2KomNMEmWme3VmDQQ2gxePgczdCxIU93i25cKuScC6Y2wUa+4B/NqjxjxzIzVVSLjMl
JR1FBOBE3vyK1zLRGsoEtuzW4JozmdWYcmRcwrfayb29ea2ZHshadA0BH9bUtaZH6wDOaGY4Tmyk
5FhuCGog6v0poCEKHGwcvPzRPYxwjrV+PC9bbwwlQ8BbN0fb71O0HuDeQaK/AYkhyjKCXQKPVUq9
iM75zKIztiLau0++rbi/NZwrRRVl3dUdLLKSUc8I/2y43i0qM5hpn2y4c6YXJ2mmwpqHEG8xe636
U52JhCIGaP0ts/vN9WPPg7/4KKNxnnd1oXGcRVR9+308OnEh0kPFVK44UoN1KfPLgrZTNxZcCc98
wi1c1ZvnbHX/NB47JuqU9bgz115iRNQcX+SUkVTtVtz4QhscELSPBaCE791pJUM0YR57H4U6mbyy
+CFZeK1vG/qe3YJrkcj+D9b0Oq8eBQodKvqMJJsczFUNLQQ6cHiWZDvX4fJpYZJ5HuNlVT/tez3v
719VkMo0YYPx8GaDexvw+ivmI2fUPiCpGr8zAefzDziPczYXTC31BnRbm0yaCv5fB4TDzE3XIXui
Wk4lQj5JPl7QenpWVMmbXnx8lABFHOcGJuKRafS8iCZs3xYQWG7BiR4z5yK7hZxDIvmZbQmFi1+3
5oDfEel7wvjiMsiIBxpqnz22vqLd/5B72ZMBINGA6Z6O8IYM9TBKlGnfl13TJKwbFIerlngIBZQZ
DKAkB/Jj6Ei+ltF0qEL5qmsOCbPB11w22HFW2MyKIy6xs9oEnkKlVqi09zaSnszRdKueR0xDGs5d
fF4FaPFU0mbZpWltj5P98mvhYgzwTmThAhA9DZr7mm2AFl+UwpJuRLh3DEtzGMYkXRqbI9keOBNg
tSEJ5/Tc9o8YKOUHBlTsMHrTpIT/psBnWW/O5NrLnwqmYvetoRURyh/BfrjMxmigX7Vuk7Fj+XDX
yBri3iDNxiswBkJvf4Q+N0A/bkmrHZ133Fg+fkCO11OkS0NmV38TAJE33Pe/FeSIKbUoq4XqBUX3
eSqq979MpEvI2jF621uebUFNGtYknsPF5Z7mMqC1WM6loA9himBdZwWrICaDJiVwqY61xKRyUKnk
6/ucUcEndBkbEv+HkKLAm+sI/AHy+Me/U423qo9F2ceQqXYafUv3SYYBMwg0mRW/XBdhJ7tjwf5f
kXkgn9VvNBeAo0oAWdHyQOt+Sik0YPIdZIDA/GMhHkT+cRvYaVs0pp6L7ldXPX+t97m12WoSpcIF
gNjUwo+FrYMqQnJa7xfCixiGR9SnfLGk1lDuEPcvyvqbwPEpkmfpUUzXopX/WGs2zHlv+NMBvEdV
/gead8on8YSSltpKB2LBChm+lzYFpfcjIirAYqX5xhXQNTh60/4uv0NtzDXi+63F4WD7BR35NatD
afStzvNke5ziMfEtlcE5A2nxY74EhuIOW2qTD6K69wXVNBH201kMaW3Es025rLWMYgC7c89xttoT
TvqJWx0OdQ8SVNHbtP3SoeHfYed60eDgsU0kBDNpEDXtZNXDL6wlMHrIKdMrmCQw5NajjjKBZ/P8
kAC72WGiz60Ux85AUb2B8zy9YlbjscQpwrhm+0fnG7vRMrTMWjx6HDsIWqonkjYkjReGZ1UqGRwn
Eiom85903adnD/Cp7Qg6iEZxuJBkfs93UXEKqmX1d2zUm07QSgCENFvlGoZebIAI2W/anfHEKCCn
OYscDC7zdv1pJf7DXyJFUg7BAuj50/OSbeAqQ2tDEZXVuySLBmIOp88nTYnoMt2LH4tPyHGk+wW0
8nlwpLR6AqvAwnRQYZho+t8mxACNXMwbBXR/Aa4HO3jCJp4sgRgHiVxgX8U7Kl0YnezI4yVSY9Lx
1asPiyyggebMWHb3GLoikNHnpLMrdq0YStE32rXxzEOS0Z4uHPdFIVMNuSUgr9Nc7KHkyAgoK6aS
fDLq+kXDhv/bMqf5TI4eMg6hgmlxocwhQCyeN3Yab6EPms6tQjxhDzJsa8cofXKGROK3QBCOKIEh
MSNtsXI3cSTYcX/NKf0NV3FOSYPt24rw+lBSkos3GjueBuUpaUhQCdWRekMGqIVA/wavRUSyrRz+
xxY/DAYv+AS6le8JJjGmIFWxVmexG5TyBKZz4FDavFTrx+ddCy0pDSwDpzcZxnCATeJoEJY9U4R7
7gN+t5X4l5FGP6lITDPMPqjqHeZjveXaiVJuDEYY5l8Pmfz2LRPfL3Xh1eXgPAHAXOY6Y5SOTI8B
LmIJTo4Xi8BjIBAZKiMPZf/Eqez0Ruaneg9TDx2NbCrpHzI72HpBZ8uDfAGi4nodsgFPYWF5Svss
7EeCd+heu2Usy3mtrX4XPJDErflcpATUd3sSS5bhRkL6q410/HtyFN0Lgf88eVMA8eTYGTkSVcPK
grq45vWj3GW/ExuXfYOuk8dJ2dDSjbnVSGC3UBUN2YlQqfBiAp7lVSoJ3LxwAphbGCjEwhcZGSQx
vXJRQ4U9qkwLX+fIoxWTZrrohMxgKYcour6TL+NpNtzY6hNqkdS78v47mZSxUsTZ8nO9nTVQQcu9
sTUXaaLRt/JymQpKpLqiJ4aKSHZoZn4AoAiTspZ5jK5YinWnip8tYT889WV2xFuNWb7iiYWl1Zqt
BdTw+Ko7ccIgkl/kd8UAusP4xLf+vo9pXMv5ogW5MR3clQFhs/+HM4jGUi1sqqfSDMKwEpFBA9wA
WvKri3yoKvVq6Umh9Wp0YYvqe4IvEn2PdbLjO5C3mNLKxrvx2s9Nm/1bWtEEhdL54VInDUTNqpG8
b/dSV17A6mynLCcE5cJCVjQqCyPHt954+/wct9OjtqWJROQPhPVmgRI0mZ2CNQw2QUsFsooHSRdU
QWI1Uc/rrY5E4LmNuRBMX2dTetEDtKb+63KyVSqX93C3Pss2UcGhqvrAbH9hG08invzM0JOTsdAJ
eNcMRPFZesfyHqGcbp50O3/3kc3CD2qcCrDur9v0J2jp4+Hx1kgVanjTZQfW5UFocsRsnlagXL7V
XvYCVL9S5IU83qUujzSWbmJ11uBW6MuIkxqE7AoQ5NIR32nvH/OJtV335e9o09MTCeU9+vuRUI5e
sclzF3DsqeKEreO9+CB76iszVgDnV6k+MZuh8hfhwle+jtseo1w/+iTYd2sO35CqZ2s3Ova2swPh
0gFrPCESioDT+7PhM5wO5Ptf0e9SWXxnd2MJV5TpH9Bx0ORcKDHGLrGQWiaZFiTUFysyk/LuspUD
KKrcjNwyxgCURoVaNeqnA/Yba/pgQpY0cTkziZoJ59DCswiu63IWplH5BL3SDiW0TCaF07Lff2Ee
ueeotZk04deAJd+QadiTddR7O934uviIgtf6I/cCRdDANQH19HlmGW3z6k0efooWtbChJcHcTetK
34nnGOyKcLR6ye1PvoTlLWPZ0MWkCUPwbS0W4dI2VTb5KBA603uAMBLQySWo+UXd55+sEoG0Fj1R
lJev/Dkig6b++fGkK6Sjbp9M2o3Qd9dPKKE99YpJWSeUvcGYNEan5FHIHmZy9QqEbJ9dHbDWOpsD
gLwD5dAzHIHg3Vl1dElY1Inf9+18XiovjxKws8EbzprL2Cx2e6I7s66NHMGCeDqCKAQDFUYmTON+
TtvtQb6mucqv6dpX2QtREjVIZLulaQ/LezyF3tcXD3R5xEdneyRvp0z18b9iYjk8/ejToL4jbVXA
VRJB1nqPb6TDBuGnUspuG/Md23QsapOce8m2LI8e66n3TAdhrVBzEg5H5z4L3EDT8jhGmHeDly1U
IxVEq4VXVGEVR4KcLQB6Op8IiZUU63Ej17aseUOfy79opDnGMLlbwBUWGsDK8rFh7xqwxKPImWL9
SmsXeKs9eplH8afHXfmE8LVlX8iuCxyT75Qf2PPs5xbGdEsgXcNqkBc7OSj1v6JbSi7Cf4hBsGu9
fSqO/K6VX7D9YRVa/LTQnm9lJfFidqhvnhZM81qbdDbk7ITYAhdwcYr/dsfL1sdKKO60IwLNK4c7
mlU/f/egEAOU2p2JeLOxQxbC1Iu03ut4Hymf59VWpleqWu4B83onTvmlERQGEdQTM8BgCbaM3Qs3
oiP9MKtontdTBWiYVtXLpmHt+oKOBiFt0pwU8Z5NXb50YHgMQWcFKaUkVoFZD+34NBQPfB3v0VWD
JZ2Y7hICfJIpsQ0tA8VhE0FK9BfLREhQt92NC0uRaeJt0/bvoRysN4SOJFR7Z67+RtMX/6JFKYXg
ybGF8u8ghYNB4A3VpCeqDw/iXNCK72CqrFbpw2NmEnDDaPnizn1eAu9tKkJgg94DYT+DKs+NckiB
JUR2BDpZEUH4VncsoeSzx0v5nIfp2limRb7Kn1u7dyOtbwT5/4w/ptAXphlqeh07bBOoKrHdwZ6o
YRg1Rl48BpCu3eU74cFnxcmBkKcERi8TD8mhAVtFVTG9LR8jxhM9SloA6gHsyTIIYLD/iJfjCXC4
/rc39GWVbwjXmonODnWLbRCAjYZoyJYamgOYoW7uFGJPzRQWdI4aRa14I9iOFqj/FMRJg+tblv+v
UWGWZdm/qQNA5Z1yPx7X3gVDItq9ZvOj//0EmWqawnA0+WLOMpZI3ywOevLLW59xHh0u/ujkojJI
Q556iFm+LmhnswiJwJ6spel1IMGGNEBCJ1gWJ8C2AuYkWlyOX/9gkt++/v2axeh+qWUusQBLoXm1
d66D9stoMKY2mnLdsKo6d+jeHuvzjc8Ca+XNVDZEe3X2dYf+1cZLsCza1FPJvw76ijSHWPFs1pgU
To8q4qiAmLBUkuHAZ9t/UiqlBW4zxII15mPAwgSBCjzq/S1B1C1IYVeE0QY+HGVT/QZ2ShNM/iYW
n9e2GnLtwGYNMkcSIswsZK2yeI3aYINmGRWzWZFKwCpe4UQjt8OVvX5gYvOIHfo1aOIDiNO1yKt6
D/3R+uEsEqdc3uzb5442jiIIbNCwQ9SwBJMzwgx9hC3wnGicIBwCzTNHoasFlta9YE+MMCPhfHwL
V1GC/6e5dzjKjHOi9xBf0bexPTHxuiyO8xItOafeeUyvoiPVG7Kte8SsLAgP1Z2YCYUDHiEAtt8+
u0uIw5TCds8Xj75OY8rm0a/pboT4Xd6Ea8v0zK6WTqI0H3WP/sZVrx9AdLMVYzyERS4Qxt/nNRj7
ltKP/Jb2CqGMn7vvBb6oLhEqmfMxjnU9hPnGNZDiXF1S+PLK+kZZN+T6sD1fJfphsPxUr4g1yA32
QdH3i9QdUIjUHy4s8wdliuhbA4+aMNNTlrse7PnkmPf2W5UnEYQ7jq+zjl3j1VIF9Ta5+krFqwtY
m/icQe83MXFtpHGLFs+T4Lrgixfsec9J/6XrdI9AXKxidlpN/zeUJDBujWYU6/Gqqh1RZ0RECyKm
xttlMS8A4EWSzIwesSJlfdBOWTul6CCiFyg+UKLv10h11lJvDsA8rZ9cSUDk4tzknWbmd49aX55j
+fq/rxS91SsEyj2HqumY2IuPS7sSc6Jp4fk9gI4ZLajLljMcd69r8z/zrhoTSJIEkNjqpJ3M4s6b
GubODzAXCuBC4M4jMlm/CNTzlgq+0Ze5KwlO2ODjX13I9oH0PPnhU5uaYSXzS7LeqfTugFytw+BD
YAOVqfdm0HcErcbtVOHjxJNzTtEvW/j5dvGq31rRqgBjtz0Q74ibZpwL2pBlkliLCbnBgozJviTV
y2+GWOt8a73IffUwJBQQjSiCO0d+58s0VM16EAWHNx2GcVGTcdG95kgDYmPHEF0onZJWYnAhBsEt
yLLG48rfz9QhbVA9BajifDZPxCUBZneZg4OeA/Kcfwf+SUkBDvgJ2K0TWuQIYZyoEDlAhWtc91vd
2v6Lbar3qUk+jDUUkLSXhkhZPsccB8tTW5jvq4m/ZrKhH98WarbGkvU+Uug75AwNXq+Q63Q4unqX
jMzmYxZ9b9X8MpuyGEh1Vy/CClAZ6Kqx3CBXLrrpUyXhdN1q7+1OqANjXNtRKQNcXFZE52MA2ZzK
lMjsl8WU71vPQDDbwqxEWGiqg8zckWO350/VEPUwgpRubCkz3ufz/AwBHIZh5mrHNeveBNnaMKkl
Ej3rf46t9pHBc6Gagck0sN/uk5f+5OcnJciMegrfM2tTHzL2OnTYaBARVQDVor6M+6M2zmbwgkKr
KrWtQUQ3Kku3O1Vp0vd8r2XCtQ3ek4TUJXSPPbHJQWx8EWFNZyUcfTYv8Gm6DVrx/NLAcQLjNgTE
VxSEY24oXhAtkL8tUYeGAI5QRfnvXkkqLaSmtXt8k7iZOQz5Vrjdj8AskUcxHlyqjCSgPZeiDKpe
s2yPvgGrs+o+hSlRFcPVMDjEv+lIWZjqa1HuQxeD6B23y0AL0y2g9jXQPF7ksaKjs2m7GKzvfz3J
IOBJTcRcpG8yumKKjfBEH+gQhx+vOFWCXZ43hSu2dg/c8ZV/pRJ9i4LBqltEXswau0VYzXHxyDUS
zGHqgWvFQEj25nWla9gtOXU2YLudHae9DCJa4dyQ3VUTHYN9NQzsWTlMiI5Bp5vamdmFyFthWuNH
G4F/wbdceLxgHX2zQ0xAVhF9ZCJbd/ds4rx7nuEXC8BdLTILhvyx20Wry5zsk/BbWkhgC5+ZEQQx
NjUrYABep9D9OUFGYXl6WWvilPGwC9pBfG8hbynwHt8dd0reDZPd1PPztPHfLudHNSwCs9Emp4ZJ
yxTs9W15Kc9tRclSYhXZ2b+1d6lJUWV19UVqm7QXbwZiIernY2OM/Vg50VaRlqr0tyDfqL1lm5Fu
RKS9G3L/ec1VQ9hX6r7PLqw4OI+zwn2H6AZl2FAVw/PV5CmKk9vx1woRpTwbNGsVxEZLh6YM3MXh
PKwN0MTKAIaMdG/kwiOQkqQE4O10UnRSzkvgvRzqGYKu8C1JOZZSrrV/T8TJ8ESOuZuwPMOp4JZx
VuX5zVF9Gg87kXfPnLWTDCMEWrICGR9aFMmqiVrpDomon8oOrUpW3IahF1/DlEV7ZE4+nK5ndu0D
oBo/caitO29NFTH2aq9l9N8WG4Wy0gcUTee7sYcnwysExiVFi4LS5C68X80mw00x4gUVqwv5KLUj
3L9klbdna+rcYpWSoomle3Zi+SuGn/7nqACifZvOB+SyJuIzUq7f2ql/Ba/Ja4lZKhn7IySWTVuz
JRmBKNsK2UfcvLrnPSQxldRZJtHTPK5MNMtsK0+4y19NveqMZVRUxCGZJt4m39kTVh9ZMPiKI36Q
o5lshJ9yb7etv5mL/nJRd04OK6F7GB1mTQwJcCsqxZLhBE7Z4VQ0daw2exyg++B8XuEVcBkYncvQ
oBRurWaeiootpj3b2Q49EFEI9VIkz6Mwuxf0HPeU98m1q6tyB33qSqpvP6PnZE9fd+3weBbx3rqD
38xqWxluE3/2KxhfXfbbdqfq3T9PO7Hcj+TRzAuAJLB+F9k3Td9Y+RcCgXiPZETODJGz4TNy3s+G
hQLYu0QA/I2aFXiqc0BsfndcLN9g0RUZcqFDx7zFVEnkV6BNaIAYrSmEFVpdmV8MpaZYVa+efwfx
D66Rc7vezPtMbtOaCoFSGjkjCOgJ9DkKZvNz10Yxr+ifi1x8LlUBerBK7yKEsVc4Fib8GzNMxUiu
2GzHONkCEOVKZjLf0cCd8BObSHLAEF4NVFoIr0t9N1quplOl0CDe+9PEaP4FsDiOM77BDwsZwzdN
ebCxnqZPKdAp6LCTyqb9Tu815vUZxHrz7ZeHw6ky9BpL9PtV2H7qT0V+/flUmmRlkwKDLDg8k0H5
1n+AX+ReoHFO4r1Un7mD8uIQKxlsMyNTV63YYmoPPLwVZ3/mDoBpI1/f/Oq/TiONVvzf8ewNkc7G
tMItKp1YgRYQWOGGkIXFVwHJbUMrzMAfAlp79shLkW5tAC/X+oCwx7oaZPJpG2yHm/zFyzhOKY8s
aDXrIyLRkxeJrwFhOA1NTzgHMjsBo3kF/aNRUk7kY94F/sfTQTPue0aSfkBnbH4rxGLcHUPFoPuL
8/IQN3Te2s/vquMZCjzB4YuvrT0uY4iZ2OzthUNqJShOWOruRlwhlxVbcmSbziXwut42Grlibe6c
pGhJEy2q1mrSboM9MRaMttxiCucI/q0yCeye2kxcY3N1LhaGN057QLBaExFtB+vdYaQGvkv2Mxih
LSesOTFPSiaeUK5o+1VdlnqqtgOGupneB5QJ90ip1nd2CeSeRjL9jRzyOzYnFeNUXtvwAFm13yEc
HbBEoiSffCZiiTfQBbJ19DEvubaAG6NgSwSexp0kQgNj7q1lwhVQsZPnIFEb5U1icB2pHWrNP3be
BGm42/D9f2cde3cbNn4Sw6xkU6qWxf1NJatxVPkc1RRBqedoE+yAkt9vzlHDfBR6H+YBKQ/NLMtE
Ard5EthimWl9C0AXy9QZjMLao4d5Un1wHBMRxgaBhFkRuiITC+Csnh3XcpL62vr+zNLUWuEq4sQ3
uW86fEU1KMdSsP1pMyqRC2FIjneKUDsIPUgOfF0LmhSwIba6HLeHDy9wfZuKarY2Uo7yz97i9bSS
0Rn5InuuGAXaxEAPfLGy3NyzQM0EwKkI+u7H3hNXL4tIOrfeBhIWTTWtE8Q/wkHbhqt2gSeGELz1
HpOJHEm43ThYgrle8qOn5XtXPHlZ75/LRRp2xD2wyq8oryVPsVveqAEY906kzBZL2Ofhnl74Vy1r
DxPB/i0QoKStKNHddYejCTCHkjm7gKA/lYg1XC8+ttXcMxP273mQNEtp5jeVRc0tC2JuQ9k+o2Z2
4sIu5CVT1TbFf4yaafqPZF9dl9QuRvP/Y0UIiebYoI19xjNhfYc1inj+Aopm+Ht1qDLdyOU6nzBZ
8fbEcgnN7QnMwJ36KjI5WxXHHAIUe4aVFYWwYgv17+fJ+ik7O39x37dkpsoIjE9BEMvxaBFlQ5Of
h/c7l50raEGgL/3YtA22HnUccXtVJ8KVxCbXzm37e0PSDpHb++VBCiUK4l4F2D3KAX7kJieTNyDK
6UiAHHrq82ijbuvKkd5sRuoFaMCqgKUwTM4ishSJ7hmnHA7FbLxUpmhpPs6htIVflwWwA+Ee1mIO
18YvGp34Xw2NEy3aHn+ZQLhI17UUbSNhMuoN93eNtYpP4SL0Y/Hvyl/MTBkgK0saNi5tZnjpii0R
hVFXflOhgREmF0DZlEHr20j8vzBiwEFfgxnxKXwbbQMrdXlKomfffPwowKXTncR2VI6CIrtuqEyp
vT50fkrhlxfNLTQtnyMqAVHd4XxejHsm+hHLK6x13j6eBwuHI3zNGvTaQAhSevWRcT9tWeQwPhoB
BAKrF2VOfoM82Dw1tmgPW3f/EHm9oZZxxJP6Ng3T6Lg6M3WJRqYlZzIpTUQ/bowGiJYlagcA6t37
Zlq159d0RSU8oGQVynhItiEWfi8AlPFzGpFTqY3IWIp+46p/pYb7jCpYDyAeZWbsQTAYyVDE5Hcv
oshF0rnIxbR75hjtnO8/RcVWm/upgve9yUJT+ZiEXLcTXu7c1sW7toRIHOe4TY0SrzBdPm58ZeYh
M0PPQQv71fCYV8dNgI7CZjqbTYhl8NENoHKe4pPtSdcAL2MC8JP+s3ZMa+QKvT6q/UU6CM6p4P05
1WlHoxshXYzJSe1pFOk/6dUuJS/Iab7d2n8ZVxFrg2AgbPtzDOhptldr2P+iLP2mis9HFsWh5WUV
Ldhhede6KpjxZ5iHaguP48/uXJlPThLcU986H4PdOdpUs5FQJvEdKpdHhcw3oGk1Zm4qDf3PwmKH
22w54yXiNMC0zTsFTePRKOb6+M0F3I+u5cwURaIO4tHjPnTwgcIbqrXjwbrkNEjuwVklOmlT6rmv
OBwFgp3zmZeB/EH1ZznzZHV36zE05ojcW8H1VpUXfhjgVm+HU9xXi469vTOKfL501wv2vVTAZ9VU
7LTkQlD4Yhz94GYOERI57t1+Z8wi11j/4mnUEHw8KJcVDwZW7H9YDkfGIhkvVH2s37I0i8PTC/Bo
bwktb6dPPDf0G6tmK2MR7Uo/WMIfGDwKTDyPAGeVXPiJWrxqXIEIEn8jNsjuCVDESEBodQHNjRY4
940JpRUh2Z5G3NhBPLqy1E8TIFJL6CmwJtmKl2HHwbuEGqndyoPaCdtzYKr1/WqjRJiU8Lo2jelu
JRzAhjH+ACeFL1+TORscFT/BIuujCEMdKt7kHYLsUJO5ri7zhNZ072BJTn86adjl/WlmSvfryunq
BcPiF1UG1WH3RjU45NOQsPFQ0pfXh1ivSDh+HeGay4XjeUire22nnSgMXuLylFHW3bQFPBcQGckj
lb52FlmSht3YKr6U64rfXtq1j3uDAOFHGvpJ6AYI14w/t9w4juLr40rXBt0N5yXS3nlNpZNoME/4
ibQNzHnEkQ0CdfqXtWM5AUcuaZ8Iv828echvlDtEQWoNCfhaI8u2eSpdOnoGNXANBkwbWcjh/xiC
dA0VCvq/a54gXPhDJq9/+UxC2tDjB0xWLRP3JTXRfjy5Ln3QMCoaexeLrkaEeJNBLE3YnGb2CGhM
e1nFVD/SfofGH6brko2tWLlI4tXjTdZTKYQFHEYFAODC7cECs0VQdH5fFq3gY/YFJPkjMP8j4nDC
upEh/u1a0fAT6SJMPx1BOTFgDutWr4LPdz7yC9QjcYROwLg9XvpjY6Z4O+LqbtgggQrSUNUI0FE8
xNZeQSmJqzWRSVBIcgVWHBoAzvXLB9ArP7aKp91ehTX1EYYABN8S22cTbqej9BnjYYuQR+34Q2Nu
9zHGGpsBrqvPVQsxRvajs3cCrZJCe8Uy3i6SffnAh6duDD+3S7xbXas3PzygZXszM9MXAG+PvoqO
f2mcd/2oEmTHyku5k3ATRIJMK8wHV/5BU87LY65n/7AFik5rxB8mmNmholcreM9DG+wELT1DvBPD
3TKOMuLn5dv1bnNaYISChUQEqBmbGex/GD5vT5fYWge7WhZzqxLxXZLHkw+7RUQR1EcTN5s9H8Aq
gBcHnqZzToijYlxTjfvRnIv9JMrV70G8/kCXnd3K06bV+beUM0nkwDvvQsp6sjUzL7An/UExr761
19Db0RSMTM0qYKsaE8N5jxw9SWDPOIzwkdse/Ry691/AbA53k7w9U9BLZzupj6KgJijXk9oW9G6O
ook2ohFOfLqzYe2m5kYw10FVXATL9GWFmxUbUZRuJMO4rJWYn7RC18JRYyc7KC/VODqHubQudf1u
KWDJ5olzZat9Lpn8OlfiJnJASwBALD40pfk+t5lcedCNLYQbMG8y9Q5a6ibTMk5seGjGrJStB3oB
54EQDfodIUJmnUTy7AVLFp1L3ldXXidDBRV++IvtyXeBLdb/ewKQGU6Nfw+2hiEJOw0pw2PNzRpT
fIW/nFHJPE9f3ABp6/R69GyC/oHmmjL6mQW+uq2sl4EECfuP0T2Ti2/NLqUCDUs/aZU8ASMIIZpz
+RyJ2PIPr7rH1KekmUdJMQrbHZbjyg5ntxCI/jViWSUjS2IkJa8eYNXNjfViI0bNpDxey6svDBV0
x1UUvODeDxyzDcnMT3CHGtT9Cw+oqjBdD0VL44M4tPzpUOjtFVg/mYSGW7VFUrbH/LXziAUzNjaG
wE4h1UiVw+mBzYNG5xnNf6U0FED2OdAaj0ahBVCcpZtsDWFKXMD9dJSnwLBstqpsHnpAsVPeVLqz
YoFKh/WzsE408chU4Bs9wnCSxXrCmdRSOfycaaAo1/YlOZbgs74WkxxwiarbMGpiu5D6Kl2f9dHv
6c8B6Pn85i6K9vCXsGoDAEZzg+RSvDW6Q7RYkosE5dOh8IqwQz3X8jbCSUU5kyhamvD3L2SIuA5g
SR7HC6/qUccy/ycXvumQWKcqKlWhxKQkaQfpc8sbM7SMv13q3dy440H3STjMEZyQscg2zgwnchaj
Yb0CA4e9BDbmxc8ikUKX3oO53nKh7oyd8t0+GAkRmvT4DDrzIh1OCjQe7KWiiEXkBBx4+qA+JQKj
mUTtQEyIWrCG6s/vAo3cHWTB4e25o8jJwxNIRKMlvmoRNHEOETmZHbSHPHIbWpcyXA8cdPzwlqMc
25r0HpJL722OkkzCarhJ4bLhZtNiPdYgIrS1pNk8BzD+QFtvXvP3wHXCvVl1ma5qvQErzmGWlnd8
AmIYF8yf7oDzixDdRFZDaI5qyspZRfZefd/XhDU37dzOjz1DZ1aEtLgkwlrYO7HZ0eiAs++HTdoZ
oKuPNrFJp4hpVP+0zLlLVnQ+7fMPBzuB+kGg+9bwLoSQSC8BtF2Ky42oWCmlOT8kyajBkxNIjssJ
mQgmfGq2grM5m5MvKZ4tNo2uDGhxfEXvDOieu8GEtpJ9Br9GBjTmzYm8egEgOGm6FRmE5cCLfuoe
SQcdLCGdkpjE7jouOhDVapQUQ66qh3hEl5wRSHbbP4AoW23sPPNQNcXYBNjoSyZOcXHmPu7flWP1
5WM+my+T41jvU8oUXna8tGaW9SPCzVTSOaBnVJXbIFHhJ+BBH39dpE7fL4kJR7SLb5E51eso6DlI
2dQJmfoa8nFCzQigscQNHHGhUPQIV+e0sD6mK5UvA07eR76YEccEEJdFTxV5J0e5REe/bvNFrEUt
j8J3tnkq5l2WQgBU+ixqi/XF0pKCs69tYpeMS9rgaM/AJbkhupW3duRlilxPWRa68GVNiKwQ9KJv
vJE3HzR8sZa49g4zin94o0oBWRqNK2QEKMmRNfzViQqGYbVPNZ3IJyoT2OKOJcynSYF0IkWLFAKv
pLxuvbIj/W82R4WXB/QzTD1P2Q9LLYcqnT7IFJ+XTJEid61S8BDeRXJuZOvH9z4OK/mJHvYFLUv4
P851AB5gzQa2/3ckO8iYVuxkUj3U64LDDtI0fb1hz9mTj67LYfPEYzZ6Nfp+L95aSVSSbGqchQIh
72AkfXQq5g8qCgyIck0cwEDhSv5uqxR02kzt9UsgV3bLC02eOfkc0gh2EV9Ju+nfCZHYaQyuv0Xh
atWpq9mv26eVSjKjXXiIDa7hFhBz5qftubNceziE6eQm4BKMieaK/fmXgFArWvYbdw7Ed13rXRS7
eZwcFkFGA+tjZmaUi8mvp/iCtnxmg0PykXBPq9khl2DFA3vfyVkWjTfVIzrdsuxvm1HM6/uvvDtN
tM0xI8qPZ5ihIij1C3gETlk3K3PEe2ehg0QqSewgM/dF3wGq/y9k4ziXlgWkVWzSRxBm2zNafQq6
qGP9EBjuHhokMhPnPLrfpsvJjY5ojvDtsWJbYt1G5RFZq28rGEvSPpcwrI5XywT08VlQVyCqG2vv
8PtXrDi+FbDTiZETqDlw2c4HY2KhXqbJJxpFNhDfFiwAC7KGkwCZADKyCLHjtlPViVyTK8lfj+a9
+4wj0rbInuFKV+y4dwuBoSSru3DeZvmGFJLOHAnPDsUIDbQjxSZj6WkCBB0qrtUXQdz251jPj8tf
ndbdygdGVEx5OZknhu79G1O8Lzp6YkYlxzIJIl+Wxx/OuEIr1CtWSqeFIvzfDIYBptN92WqAIFDY
EZqDtRzCJqBN3InSc+XpQFdqCaAiDnG1fD76qnJD65UT10A2jxVesgENQ9pHkztNYBFPez0V8BvY
NJxxDUuCUUa50Fig1JwIqRmh3EWMx7+s0Lb6cBrdk7heAcasg9RrlnHDJW4fqsbRal0j3wFWitsP
/8Fvlg3M1lmJAkA/GvGubWdzd31az6gqCMSOmXTQhMrnPf167q+qq2ZOdFpeEfNw1iCr24caIsys
LTWonukSoYNMbF8L7BcfHsBWN3gsGzntjai2zntexkokYqedNUZNfnUAW1PoqgnW+ehLGCtK6PYU
qunPtqYX0VlfrevhVGQlE+e59tFDzCXF5Ye8W7nIFumD2kLPlRGTc6Dn9rHu40wrfexz8ZoMGaF3
5L3ND3VPJaGq1tJ+l9tXX52eQ2PDoN56j2hHk2CmXPnYCatLW3xraakwMr5eTuIwLjY/QOJgX5Ke
6CC7C79vbue7YM9+xaW37QdiHu0CoMDAiYwE4AXik5+csYLsnGZa+dhawvTIRM9x5vLef9gkWmJE
Gkx4ejXdWO+yPL72HVCHerFQ2A+whMR+moD64MEYd54N3vvol6bwkskHLUYw8N9FEFKRSYyr33Me
IAW6c6KLfusJeIMNMCl8KF0GX3CHeqBrHLaloYUuSiW0qotPox82PEhH31py9b95piJMgfUZFSbn
1KsIrERklN17WK2FzWSEh8HCkvFm0guKPTNJyDQDEHtnZc8nRO9LipjoxB07KaUrtTUdfp/YN/K6
sya1+dP+jeX/1WPOpRp7im9wPVo270OaBnSvcZRcrYFUdNl8IHwMwoR4P3NbVnaRAvy4PB1Xxvgk
kwN+WwRjT3CLUtn6TpJ9zCQu9aBBmHzGtcFfc7+Sk8RNvwQoO51anP8WhRS5s91BHK4ECuwKzYRP
qMZ6ypGWeDlTEMMNfCnsmis/YC+37Dgvt38+dBYlFKZ/5i3GOkQ0GUSz2o4qrBC23vG45FnunR66
kmRdj+QNyD888oeEyaVz+SNZpi/w9/8fjFbWDCSTXSCrw9/xUmD7ifa9TW/8i8jbZQRwSAs4gR0q
3lraztdM5JnQMN9A6uYboWqSOjiBjNfZl9CQa0LH4Ruu7of8iHsd/GKqxjlaF3epMFqEMVcfzyAy
5fLmG+6eaLTX+DtUHN2vWhgbDmW8NXyU5dnu851k3FFySnQWSv8nJ2Nhtg3U9Tk0eeYhEnS9Evll
dM1xNThrQnbqFbkEYU50YZEF1tR7NABRH+dHDaEO/mKAEZ3Hbm5s6r7jmgqjRzAq7h2kblY6eB+g
wH+yDsTtCpyfbUM6f3sTaBSvH2tHxVRjak7XsrffNucUbrd1lcbLSLgp9iVzB2O6BjZu7IfkeTpS
VMdWdcgoVnakv4KkEVdN/fLWEDPIPGDJXes/M1z8uxWtmIfChxpCloS60nEBRuFhTuHpRbrZ2Fsr
A9nW7z14CbsMDIUpckrhqihwYZKDQ/r/tQzaqA28LieVJaXaUjligAJQY09H8uB9+DekjhyfAHm/
9DPFMPVtc//sZ4TlCyxubVWTcrwSQRdtykzUZeu8eGrKDqb9PcKcnx5MzoE9+ShvyyMMzF/TYIMa
Jzqu3bZ9mYtSZ9qoHkC4bp8n+qBwwKT6HOcRV3GfGOv+X879Tfl2GQ9Fwmmlaq4w/dBR7uX7wJqk
RqDE7qnvSocpWu8psMPZ4e7ygGbqZ60NWv48l8lbs6V3+YzjMkL0m9O9LDMKgsc5DoS3F9TlIuGl
EWqKjSZIDWc9NoCremO2nVr8jYxnWEqVhmPNn1KlM6/xl1uRifN3rY/emnhZEvIhTnJ0GhW7IctO
mMHS5fUiYu+/YgfjAmhCBerqn6UHGxsd+Bs/iAxil5gClmv0OEDdhcvDQpXGo+nsAC0f/1eVSnda
dbvqUyZr3D+vchcINtxywn7d8H0olBrPgb6ytK+ZOzxIsMevf+J0nBDqMpHHwowEVRJrE/8AHM5b
hmjcMXYEx2F1AxTWZBRtidRpBj+9KIOZpjCh06VtQq8uRJEYXVJF3q7gK8NMMPGu+PYUMkmXqLei
bQtK2DhW+XpsS6FXwwsQLhFX9tji021ID2WXFHW2w2GmpEqqtWLois8P5zLBxsHJXyqo6MKuq2vb
2QywZ3jYmFKlETJLJAnaYeouPqdb+kIxMxBZg0G57hYRIw1X3tJyrox8iRpj0EaYPkVA9hLoXKpT
OrMfb/jxJngpKEhyklG4Cl8MDk1J3jm+dk937Y2j2Vy9cORN48YodN92OX1AwKTVzhdUTsh5KYhK
NhZhlU6BveBvSK8akPE3iUpDJxU2p7neVRAbY+y9nZBQm30pLTj5MRU/XieS8QJOLLMG+Kc8zEWS
skN2HQCx7Tg7oLuo8erh5uDmfFSKsEqZX9JlRMuFLPSw0KUFfHr9hWNn8zblqzIvjjqFAntP1T7k
541wEA7JTRXkoAb2ihWApJNrXOFl22BGeM8+crd9N1kIJAKf9SJ3v/hAGZUI0+KR+2dawWR52aEW
2h+rrXYqw3AGknJhBWe069tvisO4O19aR5tsCdLenob/GPFW4q0+rtp4zQYZtSiIBuHGURClzeVm
V8LRefieMZdehQlBHw8NxuAGCxRfbhQRK53N/iVBcSVGm/8kpG/jGVn603Q+Oig92NQlhJxiBCDZ
LBAmQ+Cz011jdKHS5SE1AisenCpnsZKlTpOXM1jBOq62Tlaei3CbpEmccRA7UwrBnbwuzD8mpnnW
//eRJYv74OjOQdI1l7wJWiuL87Vw6RUd/zd6slbutUL2DzegnZyXGpwuAf2+gZaWCbCvpJu59xua
mlNJlNDVFq38eREuWq4F4XsCvx2qOVGEdDNLWiljLqNFTbHIBflJJ9ldRMwFxDB27LAD+6F76Mx2
re1WHD5PBXLhcB9INwxpF8ywPBC8oU9ziO06IJXez6vD+t9h0PP0isXVmaMbjsDts/caQrpux8ef
dVVrL9rzhTUjm1r17/DNba1PnXE+wy3hDE9UdfjMEBjFPVG3kkUrMXnknyGYYXL/w7Mi/808Tni6
qkyXu1Im/WAF1w5HsIdfyPmWIDj3877AtIHHERfK9ooZ4z1xb6gWXmxek6zwofMp5savERIwvBKL
iDFef5pLH8pv8w61rcyeidHYaOjG0/A/g75rCU1ba3c3p1hVopIqhounLUnXfLqj0QL62UoRjs6M
P9Sas7tmsyh9o65AFqpbQY5KfL7DzDLhBmRvbTQid2cDA9wUnUFxndrrjJg+zIVSVoXvIFzMDT0m
Qd9tePMvq+AMOycpH/pYzPsRHrj2BLtiHTK2GWKQMi+d5Wtvvsu4wJ8yN7cwFhmt9xhyv5MdU6q8
7d6wlxVje3RKLnKcoLXMWjDDe2vIOc7o+EArm3Ly3/mH+MiOKxFTpX3BO8M+Lfn8QxeKkO3FtTL+
btVqZRoY35AZCuJPOS7HmWsHzRgQq02jcqQSFDevhTsQQoiFQmfa6CeHJMR3nLe0y6zW4Rlq0NEO
NkhjW7eSUJQH/DLBYiVijOBM9IrZeRI4fCJ+D+Sf2ficUPO1wnffJjHM2sQcPWHyJrrImn2exUhS
rIbqMi+F0J5mPJ/Bvbv/I9Cc1jQKHsl168t0N9KSgTvWAqk2tX/7JrK3EyMxvT/6PDQFHv0MkLQo
TWz77GazCzbiyh9FjJHiZAGYOST6mmnYCrahS36wwcx9hRtj7FWl0TcOgfKt9WTAv1CzZi8xntV2
AgbJbkm98fKExo5WJVmD9rrwUL+AAnw3FUB0sxoEqrAYd+jnAgUaUQ66K1tfSN4MXUqc80rqR7h8
zUvS2qI5g95chROfF/iuxIT31L+/Jzp5yExF6FEs9OmPbudCRY8ukh0UkFj2ol/o3VwiV58c6DrA
s1mB9kzxUZukAtk79fcfR3XwbAQoAu09/SWa9rH133W1rA65s8X5rpsIntHNmBssNq3m/rhaUmQs
zQSce88htkuOl+xu/27+yf33WQ3BPXDPSkmhsvVN8IyAHSe/oI23CL4YP+bN3FiBCQjqP6X8yLoC
CnveP2+c3HT3wFWzwSaLLiVOLjOQmBcj9Q0sq9OKnlv7epZvW6PuKb9ufo5FU6I+NbU3kmj9LAy9
SAJKm6qwZuLT643+8exhTocUfxvFIvIQ4ppt32X9v0xBAxHjIfmGKPtCJLca3VRgYeQ+2SZhLQ7E
PYBpkIbbBzjeiJ9q2H6WFJzT2I6q/gHQF6LGkxSR747B7BR1QxbnPhkcydfqbct4At1CatVA4MxN
/W6WXElLpGjttsPuZ4hkdUSAxg0yWrgVA+goHIVQu3caBWx+/QXsEOUl3pj+ue9qgKE+Mj8EW0fs
dYAki7ldVamLWG8gWwMjSabBLVpefnchEjTPNCraBDOLjlcDuNr70Jk+X9x3IFoVCVF4kFWrPvJF
HnSyGOynLZ071wdLEtjelaL1TTd5fx4nPWVUra00dQ95IN8vxuSf4QtcD9k7FcGK66bJNgJC8OGB
3lRxLOI5UObPTbW8JyaKvKyP1ceINFhxGI3qmMazDRtCgyRAAOnxwWmxJSQQvGt0d9wGLeZF+Axm
SnXQ7OQoXtvkjOz4Xe8ncCg9WxEFr4b2y85ACbCm4BC70icvdSab6IaKjxzawkywH2US9uHc2ltI
ugYGlF9AcmyaLQCEFmS0RKyd4rdPtKp41qU9kyIuqXP6rWZPacXumrCOcHtpILPM52V4vpkzdDMj
4rHeAbD/fr2olLmuIKuAy+Kxnpx1dUVZHuJN7RJo2EF1DqPQNuKkCd9j7VebJnNlcZvdCTgt9W1y
EHVeIA0VYt7vUV5LCIpLvTg4DlqoqBSfBfV1JUkTZ9T3I88hOANc7/mN+Bq6Z73da+y+xgiNkN43
K5mYptyg/hrJBIr91R3a0YkK5fgC1d3WLfLLwKomMce8fzWbryh0Mip4sZddvRZZkAvth1bgOy2W
+akr7DQHlzGZdO8IjvkTQywCd7umBXPBEvDCtf6aryDGdgXpWrUP4cUEXtwjQjoDtHgxzm/6X7tB
tnh5Y5TcQihsqOfb4uc/eLVpn8DElMoVVzUmDOAOhiNIBJpPJ6xrZlfyOIVXUIpLivHg6j8l8BQz
Bo75d7YF7kY9l23exNSKn77CrK4S6zRXJJ7xp2Ax+wgEXDVIsl4XX+HR+FJ5R5WuBbBcxMvAbwg0
5BHO3y2977Yq+ONbJDA1oCILKSaeWMD2MeZtnDRXjBrZB6jrpqXBGBVVn+85xlLAxb/heNyXJFtm
Y06CfVIYu7G9s3LvA25eWk6hAmMe33zDdCwMPc5l/NH3HFHYFp7199J7e/k3sLkIBOKB/YZSUFr0
A5vr/1uGd5W06Z3uSZ+zZFCcf/oDG22qgLTWLqSQQt8CYLB7JEUKxeDUhdpj8J8m2jTO0gi4eWzt
ZntDKKYJtDLbw8Y6rm3wdPyGa/xnVthdwrCe0y7cTWL+/f3gTAJuB7PrvHEL0vtxYx4zwI0F+9f9
9WuIZgx1kGoALf8nUtIVILBGohSoATxots/SJf7luQ00J93fK5pu60iADT6nSO9uDtOE43fNjm3y
EVwZJlbizBUnt3Py1cazAh6BHj6G94tn6nzG1gzOZUIJBXzu1QfQuPxYhSMWUKa32VgxZPm0lGmd
rvyaZTW/3ARq0VyOQ5OtWIQsxUWVVj0LoyBbp6TdsGKEwwkd7qhjCZLJnO9RaCW6SNzanqi1TIBO
0K13YGQZuON+qtJoM11Xu8sK2A4/2+JlCsHZmCCIOAPUcby6UYA0NohKbcUKOmi7zLYL1ino2zYm
sts7I/7u8GXcKCfYu5NdKhg7VERXAAfSQfLs5zL1z+DZrcA+YFR9qZmLDgMLDQJqDVgsBqtNWKTA
2ewE23syU36/uTkEv7ptGNjdHgbVSr73Whcc8nH5OhifOJpdG0U+ut8D2MYeDBcwfDnV8gyMILOz
GLOItYvbgxBSI2R899uvj5WV1vtQS3Lt/aBGpefF5CkBJv1UpDE5fzgncRI9EPkSEDQlxCAU7CI9
wCmKiDRgAE5aSaoFU+UePl7LfhqkxnHXRhfdBc5r3yWt8FcG6E4i3hlTq87Ld1+OChoYKdn+Rqgz
Uy9qQy5Rqz1BgjFPsangDOxUpHLToVQVswCrKYwizhce8ByxI0ySjEiRGOxQAjCtxMNT7rTIvXvY
8VP+NNSTuusbse8SIpSSXxK0c4dmb17rcS8SiM5SCuHmsuvi7HPzgAM3Oz6Z3Jlj40vNVHrmpFAb
i1NRlperFE7Mrxul3Rt9bM06jBBUWNwrA+5o9z4XyOfGKREdiV3KE/B15ZTjiQ5g9v9wE2ViOb7c
xnmCsI8qnFfkBwf4f9nr26kVum8urbZTM2kU7UfkDIJqewNWTjHWKfzd1+iSZ5ksTME79TWO5iu7
CCaYo22/BKVY5rGY2JDkWwUrENSSRGWtE6B0Gf17j17m3SdYxlSg4LhJjJ3FSbBIDgC2mqFjCejp
4CgDbc3FtKm1HPXw82NwjCsAjLFx5hS4LKC8F7CAzCE7FnqJh3yOywkOpaDTcLLMaYWczlnP/qiq
pgddAj0Trs/73vymlUZsVWTyVflAJdq+c9oYQ1GNaFRXDdVjfcudneVUCP9JkQWUeI9w0vAKVBLe
gFawb8wJN9jY1Xlc5xgly/BmH6bWtTUxcIWR9dKwfXZ2ASevrA3lE6PPDJJvwRzrYjI0mMuP5pzj
6deknl2mEyFGEo4ak+zF0PxUQGb4LbxWW9B5dM2f3JAcd1IHnyQIg5Zl+3SpZEojBQj5jpWyqDHL
lMseh3zLUpBxzybVcmzo3azSi6cVRaFifMQMfx1RtnelwgyuOALiZDartSkyBQTzq6zo8XEpC2q8
s2Ul1Ppo4X+1fLnx/UvXddIckfjbBOD4UrSovkrDAmlOauk+fAoMyVYsOPATyBcKSmWpu2FZFtui
goCUKtq/xKnEx+709SnlM5S1OWPUkoVErNB66zA2Ja9fwENJ5pIx0IKfjcRdn7OfjPh6MESo+ZAh
WHlH1hHEC1N50YN+w4VYQS0dH9Rj7Vzuz1Da5L7ISqe87rUfgYR8sdqPsStzTtwTM5Th5EoVPLL7
W8fBt7JZjcze5eJunaTClE3GG0NnBeNxdvvOaPlH4ieHd+R0LyvtlIaU4irwT2aeUFrLUMpQc1tI
btFXLud0I6yOWPUsZCiw6qil/WxPYh/CuqLRzyxDKbni2wamnkqftl74ct1vhm5xiZWZPkTlzQvk
ITUdXhwn6vwqvLEyu+FduWj0Dj3deOMXeCrRPWANZMnOLidsrWqYH0VG+xx/pTVCq3cYI/P54B6y
A/TlSgV2tiZTKfYCm3rFX7yXe+8FDclWfbaKg59nUklEcOqgVQa6SHNVTCJ6YRJ0eCbDGa5r5qlf
t6WSMxYQX8Kw1816rIyofb8+zP5nwCongjiSdLMCH+24v32egClRr0cZ0lLU1esI1LqbfITqoL0S
D3fcLggW1h9rlZGhGaGTJqigEVdIdubBz4ctqYwE3l3mQxU93FUYyIBqPCO3sz7RvOnWV5eA0aXf
strmT0CVYS8SMU7e79nqLYAMcmX9UrFX7TzhjUeDlXenjogEqPcAl7m6kIkX8g7AOt497HBHY/3I
2dUEknPa2WnT/wkfg/dJ3W5HbsLxlsTB2+cF8jXsVSASYcU0nFlnNrEZAT/U/KAvOM9tsfExXG33
TlsbTAiriqQ8320VMWhlH8uSiJ0PbRM4WJqibWBh6MVnRX7avJZuMRkGBlHdSGiVPKlVWa6CWBLe
pD1gh3q5GyspMTCTgjOPLXhS9l4c9JQ7UupqR2EA4esF4JSHwNNAKvN+agMbGCoEc4GVwn8f+Lmw
MDZMBa4C77In8ecvPsKK9SAqIPiUl87j3nkTeh/JrmL5ar0mkwPmOsmTWk8Z7Huw4Hw4ybrrFUek
EwM1keZ5sduhKQ4nQDBFFtsc5ecPtoNONJJemH5kdUPGGvCVcq5HAQupto+At3jK4hIwSePlocZA
tSlFdUO3wOFRpP4yKvWMvhDUu8ViuECYXyY1Tcad//D5Yaqkj1AOzN2Wvt1aw1ydUNUhwy3gO1R3
zAdSZj4tY6V00EnTyeeRDbnqocIgdE2zWiKMOQH2VIzH9JvBj7s3DAOJduDISqjf3EDQ5rqhwDu1
Qa4/btLJvkC1JgAMGk599ErGZieU9/unVJQMuCYhr3zPCTCSgebovyMb7RhpP65v52r3mjzV3gss
4HFx5qZ85W0Q5TFFVqQ4v7P/AmxCTMR5BjMhNloe+kELy9WTr9Y3uz4UL32p4AiQ9x7LDMcmnCIS
eyfmAhTVHy7P3pNOeUeY+ibHufzJHCLz4adD70UJpeHe12DjzejjwnonwG9xOdj0u/LlbDsQrc9c
kuds+dqnJSQnlYcU2W5VcvxXCu2URooix0CwTPOeenehvvrHE4vJN1AMFhxnO7es3sE7Y94xTDBz
oKXNl1BF9LZPIi5ahjR0I7UbJCd/tiwknlPmeHwEkGAJHoUQoY1OPmwaqH2rCS9wkqx4dwuRPtlg
4kWUaxSkaepWZhR9YPLTNrgnvxcmORzxKHcSZFYMPOigGzqR8/KQrjzccvPQFvag9a2JkJ4h7qfz
zPja8Ayk3c/gtKF9IxlcRCAe7Rb5tUBDsWIH7xsinGsrliyj35kK9UDHSN048dgC3+oBtzPe8hNz
64lr3i0EUrc1C9/ggerrYcPQm95nNuoPnznZDftHDcJArB5Xn02kn0ozNZMr9orAy41bip+Bx0e2
5XEDHQeB1FCSjncGxmF4jiLdu9DeBC+aeP5076Yu24ha7t6URyoK5H6EBQzpZxlbZZYogmzR2S34
vwKQWTi8QfxzZ4gH5hLW5Ux+fWqWbRUkvqqAcxeKlhUznPylLTNlactxKimffXMnzOjkcNKE5ZQx
T3OlQv1/WDfjirEM6LPsbUfg8WPF5GCniE/gw7fypANps7iDJG+mqVRYF5IVK/CEey7cEphrHw+G
Y9k22Rc2yJTNbaUfaj3QQqD8xlWgUIwARFNK5w3devORi/zZ3rCK2blFQLAvWDLkwXjK4MN+QNCu
c7d/Ffk+IfZVZaI1XbiuVhobeCB6EdDmBABVYN/uVGCf3JiAYuMXi5lDcb7Wb/bs+nGHM1mDN1T6
3Q57gParDo8xpqDa0mxuFtcGOERWH1fJQ9XcAixcHCbqvSIWNmbIz+13+OGajCIlSckOUyYGD2KN
7K/yMLDDlW3IFbzntdrdX4JKBOp/p/wdfNZAvs6oTXdvrXlWadC1X4VEgtXNzZzUjdFJsiuFei5o
BD1isr+wAW9MR0/rKK98ddAxKqLLT2gFC+NBFTs9DvcqPMJkmXab/NLsxGoFj2SZLHVwolHqoXxb
s6tPYmDd/SucRDqlcXnYFUpx8FHhQVhohqGW6A6Ke2ND5cNM/VJ29FDiZq0DkCWv+rFm5OVgwfWh
xxMg929Agx5qqzH2t94aV0xTrjzLFwbHtUn3JJlxd3rzSoDlsXJZzOnY1oH3NCdrxB88bTjpq0CJ
E62VAVGzKoYFb74lh+xRPrDRu6YYcXwrI8jvJcN6RAGSR5ebsBG6OGl5GQAp/BAkf+6aOlOpvKu/
K+JP7OOtHAeyFNfSbXKzUlLLSs0QhvdkvpVkA1M6WmGcyxRd/NAIe4JFtFVJqpnLS8wR4Xra+fqt
CvT8ox+JxCmBUEfNBxgR1h5Kxc1dOa0v1SCjvkdsEHSje1DUcECOWHQuq4DZ8PzsaUwPkyyu7K9S
Z8d0vyHLtTbTrhRvg2Y8gWypx9X8cNKpxGa82Asx2JMEuV/RNgaWsnoG60SziH7zwBmJIW2FnoN0
D0P+FSJpDiyavuq396vCoaPF9yaRbevnMACUi23GyBqSf0NTmk/1hgFu1mLE/BF63Fd82ajbn4M+
xgxGqd2onaXw2MHbFG0Nw9U0bw3X3t3dO6h24sUJP4XaU0xyzwgIVvZyWTyulzXEobbINroQb/g7
9IgslGgED0VR0Jgrb0y1xI83UPFHYNyf9ZSVedLyuj3FNy+kcsNJjWsW2hZRtBTtIeBldH1yiISa
+XSY8KxSDvx7YQb9tnvd/RiSv4h7HsrS0XVi+Y/nvgcWVmvzOdHcnboOCpLQt7dfSRsr5u0ttiLu
8NvvLtW9tGnwinMfqRlq2UkHNWM0TY2s8/Wjs5qZ2sRLFCAAHoJOHJN+vY/c+Q81OerPbDOnuqTA
pA6B3agNMuGETxE6G4/0D2c1iQpp4HGhnc704fdVWhi6OEZJ99nk4hBJBR3DDUYsnJt/HYKX1rsy
ywp8lmA5q/73oHL9l3YdgZt7nQ9IG14o+5uT1PmYk9Et/3NPksFBcryI8KhKQwOjGGnMozH832J9
Y2fM/VbOHVmiJv3KyKt71iXx2IMg9iOc80YkxvdVc0NF4lqM5zupwuma56kl8Sw0XkaAgPycmKVL
b79z/oovVt5K9QKEFHxHRMLBzL+XmHwtNcUtsrtuk4UH+J7RqAWg9H80+qn0gX5QqOSdWlIS54Up
j2/zbnxQPBqkOZkMPlBvXgnYbnnwQZkgCzgifTmL3YKwZKqbbmkN1S5bZ66k2LlrIJewV1sQwQ7m
Lz1wkWEwdg1wZP1fTZgQsDOWCtc6qqZojifvp689N9zNQh4apl0AMmW7JdJNdSKm5/+blDhiT7xW
VBW1VNk9r6+rg/1ZgSgAeYz2QKoaC6yl/8AFmDa5gnfvtpTdzBhQH5LoMdIumhYNi2er5FNQCHHO
QQjN2+vjJUeH6LPvj0QT9M4ds7oZyu2BJCS11RkBO9Pc6Jh72XoiAQX5sFRjCOimpwC+7JgyYXdm
lBH0hCPdAmO8NtFWxXc5f/AFjANoO9FYv0d88dxn897tgcOQwvkydQIuY1iqd8kQjdJ5kO/kC5+a
znRABhx2GBEbneHs3OAGExmzdjAGD898rIniDibICcJL2V55CpxmDzDlIce36wKnq0Iidh5euIgg
gza2HcpBVdmVdZx5x6rkWyRCvJqPRm4rtKlxgpTHMT2B3mqHXKfEW0KRppCBp6/0/omQlTYJ8BdL
OpxzD8UpcKRv49nl4vzmNRFBWMSjD4YV7JOmJbW5Bn0a4rVmx/1I0fXqtuHWBW5wWcRydE7Aq39r
V0VyD7++KUJW9EzYrI3dYEBl+MyVWxHlMYgEHyGhTqqoLTEF5YapiwSBa8qJU9IZiemIvy/fD5V7
lD4hjhpo6+oar3cHkoQzw6OOcgxxtV3UBeYEYt2HPUY/YSdcmJFum+4pLs1fSn4r2xFgrtVRVpb9
3+1edmvd6ZHPpYE/0MsD4VA/9ai/hn6/nODeto2DAV1ihWdbKqPY2dFQWW8tnDTPBtnqkOLeysRZ
oEE2qF0ycC9Wj/2Zj3wvTlXmsUFDgCaywnC84rN6m0v0ocLM2g1fEyKO5T62Mv07WWooMZF8lPap
BQGIpN8KQJN3jd5Gi0Kxbiis2ynrLduNqgdo2Z21ZCVwY77oYoowu1Cqf7G6F1FQguMHyJgEX2A8
9dja9LBxrLGtOyKIR7vUBoe7h+FHPQ38VplHWX1UbTFLWdQ3Gdm9ByLyQTe9gcQiBlxdTSUIeLHm
maSC888XUCB6Lwqris1+wrAGdaxQz6cW0AUTuq2U1cu9KeNpJqM/a3ntWwiDT9qMu+8vf1BmHfMK
4JCQKucAa7nwg+7xd1xd9b+WTp1rFOIK8PS9BD8/2Ck+euutOIloF9UGW7w4PwLeZm4q7ZI2oHTX
wWa9rlgr20WIRWs13Sxo/AaYPbt4YT9vtwYXU+sUkVWXE35wwXKSQTyW/uzs0X7mIAfGYJoj0ruL
aHnpmA7W6dCGi3IzRtfjYLX3BezFDYQQaikmiwMCoBdG9mR/x+SyZHABCvjzsPnVYsH4gQIGl+uk
z1OrxpFwJMg7ZZEYGDGymhFTpbgeGdSUUbHWstK8f6O3agViHLLatBR7cNA5cOp6nWzaI3NhH9Kr
jpwy34pHU9AugXBpnI5XZlo4Z9eVVk847/O/8YZPRe3oQmZJUq0j6n+OScyD+Thk0mAxiCp5qKnD
2XNu4Y6NftFdPzcepTJtiAHxXb5/tyl0A7bpLJmzeFyCDJL7gVi+Wt0ElrGgU0fO8n/BvfbNLyIp
mBAWvOgT0czQCdervg/7IlIoGe4poaewRnWvjoJHSTUAVePCMz8WheCijrJO4kFuC2+0Qt/58Apy
rrGRNpnxSRt90qpvdMPz64v+w4YgOWB8gRFX12IbJ1HRysX781Yo8IYOcoiKoUf4pqFsqqS+XKfT
oX3Hwc1vEfPy1OcYoqrWUKF1uOGCHIX1bnou1c/dTv+QjGRzwhEjdSkgK77pcGbvkKL2XEn4tyH2
k8PQBXiz/JeEiKLBXNfUWTt+1TU7E1kCE4+yFUNttNqK4FyipiOGulNWkDesiuF09AxvOJRolu7V
U/m0PenYkVKYfcwKR8GY9T/QcOVmE0SjpBC+a786mN4RBTZWuRSXkyGyueMRS6Z2N5tV5beFs8L9
xGJepiuLO8A/6fFSfd0enFeW9ZmNb3lcTelm9VqoB68e7jlz2B+VE9uJqBgbHQ1tgkp+1AhO5Sy0
pPE9PKwuP1/YAffmgksiJxjNYnkW52Q3r/OuMMRH0/IWZrfzvwDlaU2nJOsTkOfqqdKQJ6pxew15
feYSImxBJUUbHkSqS33KpeuqcnincAmuZ1zQMnMLA3+DKuYJDx2OQouhIwwUwVRtwPnt+sYodYx5
7D/li/oZZCQu3pGD49rd3SLs2YRVpBQ0Iui47TdtsOkZ62UE14dy3IpcZqt4BLQ5KyN+kzh53T4f
s3RM3xRpj16AAZHyPDtvqjyZCIn+ouPa9NOFWqtu1nI6mZ+LGI2pnzxQNZWZh+uGVx09oM5LGEdm
tY0WiI3usWUUxp06IP9d0a6pATTg9bxfdLsPZsiYrAxDf3tjiUF/pRTIhRhr9do1coaJppUWqzm9
ls/6E9rVnR+ZjpD37LcFSdVZVvxbu7xcYVNssBnvVong3ouC88FUY5KzbKh/QGltwI1GXtluOG84
jgNS/hhXbebLsCsxOw3w9Wqfu/sLga0Uv37mTDwjbWzl2TDquQofk0z8bzN479iuVzztRj/G4VDU
vxjv1h6yH7OSGW6AsfLtvIVFMRDNxK5i/SvrGoMLczkOKLAnAcZWJcS8f73lwnUTq9difPEayfzq
Qzib0UaLs5OiQf0loIiu+Edc0E4tNcgF+LGuT3Cp41zug/KRksffXcpEd1kV9JtpDC3SxvUn9pyx
P6heu+akxeOB5IgphndnD4D7/eQuySROMYdheypY2/iFOYiTOiqo5iFK5c6uY3/FAThIDeOyF75S
H8WPy+Hr4fZ2GJNntClJUm/ig8gZeyePIC+tsHczxhTToZ5Sq+D5B/hNMpDmK5w7lciSbEAlY9xH
RnHA2VGaoLynXeFNzmcQ0fmUrSTLUZdEZQPfOEOLYll2Y0Wo0g9NeKUsQZvggrcsyffTOCPmGkQU
i1be6QM82UWVsS+0Ccg3FDTm1AvhjSXn6lDHyLMS3Qglt3qiTY1Nt/QRDLFQGGP3HO9ziqzJ1oZX
KAd6VJpyDDqNS3mvj8d2z4tWrkXxuZDAp5sDiKtfnxSHbXC1RQLI49j5q5ZrT1k/AmX6QBGo6Rg9
0BXKC4jTAxwF+Vboh2dWZvx1BxMpq5i7JVnC9PZsKt5+hPqiwZtQNLnYGgCxKoP4jlfoP4CnbwKi
1i7JVXWq3u2NdBRJf1eYWIc8Vd+5K9zaSZDYL8BVoxlkgSNY3xurzLA2tToyb6CTBeAdMTGSGevi
8k+/ZzVyFeX50gL40nlq1R31x0rUuirH1NuyjL0DVIk1RfssGR8SICOyTDGLqbxcIWLcyyO3AO7c
orqFoonT9pT5hJtKaF/QsHridZ9YcljANRic5SUbV79A0CJyQ37OevpjCFfKypHr3ftMfGUiAsDc
PRoLfavXX+ItnEkKa94C/O9Kn8mN0rtCeSwS70/yldUaqWDuffDVTipVvlJvS0xZ88fIY2lf2gZ2
xM8YPieOAe6PH+yGZqoMI0OgVJQfMqIfcYvlEIPppiSJPCwwP4DNeVLOaMJZMjIUfFIVVmnOu9Lx
WceKpOTxu1PJ3knSWU0AQg7Ng/5/wJqJ69X1owB6NpoQwjMCknV/rfoKdYvi4/CQnUF++p/nol15
cqcKnB3D6bHbl+w0eigF9GUwyNskhOgqkioLIo1vCcGtD9A0vzpe9611kGCB4AIqRCDiwRBw7CDV
a7kuig1Uyigwk94B5hMdMNE16Goyxg5RcBP9ZqvLD7xiqqeXfmTfK/xekHBMUByg3Pqogjuk21hU
kpeQxfrSU2Xivg+015fr7wsJ3SG78+sgEP3RncINr2ygU8IRPKljX4pPlkJv6/rE0AWeAQUHr1+v
NJP9lO0pCugG9z7iGnIxS38fYVcK0yqu45ma8sauX+GhilVlO4oKvdKDvowE8GeLzJYfVGTdsaJJ
j8bRLNTgi3o/rv5lge7oivgDJABNcGdJn+rFrCgW7jZM5oJgL/V/EWG2G3Pvd++3TazzwugGxLHC
q/tGG66omwABUjEgn6qUDg3Ibrb5QuKVgUpA2oXj7LbHrLnz6Cf5Bln+omcC+ulMnE94CIZppyoj
R2BFdrv7XAHFB6nqlNjQvAzC1RF7Zi7Dlrk5yxjFrnYVWSbmKOT8hhi3adMgPrafORZS4Won736P
SlQQ7iVebOwqhS9uxusNciV/T/RBUYovDIWlMzgq2j1187IcQHAtYBoaKQiN0FdGvdoWlfPUXB1L
jGk6pM/4Kphk2lc6ZlcK9fh9gfEslmnRk7eHACyXYWfi2lQtb9bJi0I5a7/QeGiCCXjarAylRrs5
pgjJaPvtRAEAPGbfwdM944BNJpJ0rAvh3pU3N/DVCYCvjtwMhQj8edj5pQiTNVjsTyltCZgMhepb
4W7WG3pElcM0oMa/d429ilRqdutpm/Ys41UomkDstdZi8epW1LJ3w6ZyFDaQerh86vTYZ4U3gsWW
rOzDehMw7iTFsnsHbrmcKiy7XbljiFoOC/EneCoU5qy+yNen13BVLEFuZ2D4vY3wxj1PaKF6uVd1
ScHJr6Ohd0NxAhv7x+CxmzuRGaLxnulkDZps7dTb/DnCyBzctpVFEWfUFD0TPqUXkW1mT8Tpm5Oy
4UQaF8099Z1tvOemawTCQWwYSlZNLj7gYMFtp8lX4OMAfHkWh5Djoa6YA5floJLatrKxp0USUy7h
uAY1uQjxPYWbEFva0naz3acYIBmEJhS11BGuCxTYaPZbndFwI/jI57ajdlAJIIAUs6BRJQ6W1CN2
sPaIRA3byXC7RwHhTpkgcRH5Fbvo6tIRbiK7p0H+ZqyEmnjZRx16wvDSbQfJfwhscFhD+ilYsQFJ
Dbh8NFi9HzlUz5nnH2y8V9gm8G2cTjAsDmkozrgM5jJN52ktPETYC/Rq7TWEtbGQNvG2LfJI+qTU
Z/7ZOp9l0UqM+Pwv9XbmOkPu2DB+dsl3dIV397HAXHVZ4b29UEw4xa26oQhCEHlNCK1HVUx48ml8
F+IC0C+nDii6zegjtmBgoU6ZpoNvRL16QrsK08PmzUylrRD1qNU9TBcXjODQO4q7VgpiidXiu6fI
Xohay5KBGXzNwWI6b/HDz3+x9j+Yg9xyEzwjhm/wZSMh0p/7Sqnqm275ZRkRtv7SVeHOP0SMrExH
GTtiJIq0CYvhV9We7puTA3K5fPG2mULOi3xY29Dg9dzyyc7R3hBKrr6YEqtstmtlNaxxChUdR4xT
lLNOj3hcJJ1uzbmtVR5jGasWhG5+96ri3Z9mWK3JP3Tl3rxBLyA57palolhlEZEXP0NJ36qdZGsp
cmMg444B9/iByncF0bRQPHMu5PIiXDUxr7StwPd3kgXxvX41QtnBL3ceHDcH9dS5JzzVz/E6VI6f
nVc2BEtycXvk9FYfnC3KURtoGkDfBqfAWHTuAGuK5bYqg+5J5oWHPLsnr++8Ooj6+JpAsaglCpti
h909RgFjb89IbydpjyvriJiSHzjag7TX6kB2ToVUP9ppn2yXdNxH0/kJweYiCGJLtWoilDf+LIOj
B15gIV7yckjIw1SXWSVQn9P7pbPg8weD143JGxdsR/1uxgiSCio6DTFtG4qMRXA+ZmIjCEOn4twa
7Forj1b+xggGbot4/kJr/sayouQiQIA1Q3VG0XeFt7YlfPk0ccliwh72YgB2Mbsl1w90teCzllE8
FFR7w+yF7tmGbWI9FpYZ6hhKNUB3uue3ma8MMNUw/sGywxzfm9F9zAiFP33TI4dGoMfe0C6BNytk
YEY3z9ymYgfwfiH/rdFppwaJM8E1b1XsBQCVlfnq0ulleKJBMMiTJNlrwV0DkxHxjfgHBHvM53vs
4GSkPxXHaRvNGPzR+B5nkbRRgT1GgO99Hgyh6sltke5i4XWs1QI+FBNikK/8ZGjZHSmHovHRUGUa
auK38UTUQpwfvbhq3B+/xZ9OLA+yyt9yA9k9CVdEiXQ9SaVtSi023BJTNr6hvsH0XWHkCcQXQ3lw
XFBikaDh/bL/5d4LCiV74KsW5q7nC2HAggYgspzbML8wL1/ahHsXVAi8Y4aOJ1VzdS0RBbLWoGAQ
UbBr27Tz8/Jgi7OgXObF3EC7RTSESPhlpgbgM4jaoJyiGnDED94FLc5niB4e6H2vl3RFGS0eJcWx
Sinl6EcEFScEdzTlGiD8TqK3lWw9GKY/63C0aRIPz3p+jG05B/ND1bDMQkyUYINKiEdqGVmao6RX
OdYyzyVBKI94ASaIml4uTXWZgBwCJSZP1foGW0l4K3lfdcOF1KgrD8lBWkWA1w3tvt3o2j7EdMx5
NhwMgRMbRN4sGin5ci+CwSawANJOvHiuXXLDioEw4H8e2fNh4qOpjNpaIF8bKsv3TPY3acBL0Efy
XcHihOosnxCK7H/yzJ3lwowFpdrzxZ0y71Wpb4VCSP6q7r7f8+9LGz6cKPyOXzmX7duyhU1W8Dab
3t8iUTiPZctw/pj7Sl17xmAT3z8Alz0T6mgX8JyiqRtk/n0Eo9ZkB0GorHKqintM1vRNxgpmxZmu
T85lqumCQf2L5hmhBQZMZSsQsPeuW9Y1SYeLLo6blHTTjg0L0jlgDph84fso08A0KBuZSDu2QfZ1
l6XKVpq32GIeHOh2i5BnQhll/8tCXq6JLrhqSa5RNFw7htWQ82CjHbzpYN5C8geiH3485QZOG4Zd
ygrgaHDnWvFtJBtuZJByV1TwmDnwRDD58jEJroIzvvvORtuXRcK9T1vc7CingA80oc+gNolNgXv6
CInFJxauHfu5Ov+lJXrrua4hj1X6Q9qIVJARVKLf4khyDqxRb2mi4ZXkmfSUiSWV5HCJmXn3QXje
qUOaGxwIE+6y+VVivi9S1weurNsAA3+rUbECGkAhgaiu0zinTEgODPekxzHEvQJKeyNl4tt0xs7Z
igmfGtN18F1svxbzJgjgK1ddopaX6nKOLuTNUmsGHmRrgJSVLMckF8OLZ8JWpRqsSKtTmPnlRHcb
Gv/UMNdHkEXDt6btllHbMEEsJIwQ2MsDasPzPvjXVlr190D4GYaLTOeSt4YjN64Z3LZis4WNjItz
nmw+ecU1zfryAFZyjdOAVeaiBYz+gWjFa58qmMHfqbaudRNqzDyOsw9LMd+bkKyGkKKGCAalKL2E
ybzxgYJXIPxQKFwAQsHzdiBVmmgTY0mWmc4j0KE0woMlQbo0fH75U5D2/9q7mitI6J0cvNbPK+/1
TuVBa2HkV1dyXXYbTfR3zxY0tExFu7InKJOA75kpxknL8FQxFTZjR4C9wLs2ruXsXJuKf5ByMxUT
OgWnvYUNx63liO/vhY2xMx0AWi+8yt8RQ0ISXC5RJ6rx4seU9+d5mcrdrlx6xHzfkmPGszEJiEZ4
TVgQohH7BvUsbj6VlFozIEv8+KhLB2rldIE12XAzqd2LdxdRJB+imy36JF0kxNo9MJ7PN/ZLD7rk
efKeLhP+HW4SOIUK45uBYP5WzwU4s2y3bXB+fhpOUlUa5Pbk01h0jnaAKlGVd0E1V8b2NTk0LMjm
IaS7UI2GgAPVEGliQS55pR//afxO2X55fVeVM/vWGL5EgBMufu5BIZb1j2lXhcc59M2OjYyGulq+
B/pUSPH/tX9aVMT1pBX58n2ieFT/2Vf9xHQ4r8nXJXFfT825QZOR9MaEPWezcpUiVkkexafSKU3e
4DPQx/9LnGwLpTBtZThoNSvlMt5zMEic1s2E+z2EHUnYPRzKr8gEDwfxN60ezG1icTbH2NHcZJJK
FHGW1Y3dLDbL/oIjfAUYNcfwiPnxmk5EiRDJ+Bl0cUd4cI93p8z8MtQWEulhlCqbj0v5DkSaFjll
DYlSh48BIfZ4Y0EgpCDEYAa/gW6nqEIcSpZ62Mu7JBCi+Fgbq4rNek+NWmL14gqX9/J4SrzhRyyy
VFvIclt+zX877ZpAP1Xl0DEQ0+rGDjHLwBzeneRagWZ6v4FNLV+m/sGa1PccduykWuKUxI4dVsOl
3iCnbSWQqVL8w1flqGX8ysHlf1MU3alAZPyowmLl9nmJE+mmuHP1zHD8SpyNs5kV+8pcTcAGkndw
MnT3Vf5KgXklF3MzIxXfZO991IPz5eKwU1ZvvmSGFwPBnZY2f6dKfnb3V7ywBDG1RdkFS/49CfK+
MX5mIsmdno3TtUuUPGzjqp2TJOZYIT9BXVahl7f9kOcDeDfBHSG3QC6I1AQTMDZgpF0BrfXBpJnY
4eEg5ktahcuTPh5GlZYdkA3SjfZEIPZZ8x/m8eaUy+usHVvjfLkwgXTTpj07CT8nn2HoKOrPal6/
VGplenXuu0oKiq+KSYasEcPe8M42711R7bYZIPOsx4o/q+aQ3CHa5dm4z+X4C3OEj9DmL7yg9aGp
fyLMwxSkkglKWrScNTQ0FNwfybp+g8sPRbwYijMe8DEIHkI5iBHtRMv+rKa++aWtwMloMhkRzddq
CsQgRfcoHXH/C/fsGaC/Ns/4wx8WY4oiNrW1iH1he68K09ZZsryLL3BrHK6ZPBNqW/ebHfBn8apj
v8epXSloej7trJc1R56+cb/25EmlS6Y51XGxUyh+MV5vWPO5Lp6kNeAMdEypoJqNhyHDNzd18yFF
D+0a2d3B3RAighpr9UuDkRZIGR5BSfACZ6wMwS7xfOloympfshubMCmCVnUIhvsCyswcRtfBzIsS
A/QY0YxNE6e+vBoOEet0yMkv0foRmbKIpOW7l6UMCR3qnvOoEC9ozQ4VJfdb49QTaQRt633Odtiy
fvzpR3KwlQzoYSe8MHyFJtnHKhfwct7BMQl5ceCiwkWpCmAR8qat90YMB37ro27tLo3Zsu1fMkik
D08ziSanO5Tq4mVcwSVSLDZZPlwqraYvzT4mZ4Jh9ALv4i2j76d3tRztOewZuMSTuqAPYAQ/TEEk
kmtz4EMoIug3Uj8Iyb415Wp0b6yIRN3n+frpkAnTGrWhA1UqmiesQbVK+YGBTSqmBRjYyORdT8/B
z2DJ5Xgx3kUsIadRYIHaWYOMRljB9/dk8tf96ZAYVIc8krjvAtjuN2srL2hitNoivCvhgZwXm6nJ
QCuUFu+Ac1njdpHHTOwd8jAW8z8j3yNmtWNFBslu8Jc+sNt0Ml4002nyxgM/mizkFihBNz5VNqtC
k/zAyK1I3nNWELm03fSdPkk93mumUKc/nT7pDb0A3K5fSLbdj1RFLCDBci906xWYjG/A55ZXP6nr
wbnL6ifMYRuaxKKlHl44phCRTVD6rkAsmmnTDtPEPJ4MiAnOIot0QWKtjumtMWsHqIe01x5+NIJy
Qol8wMmyP6dcXpl62PA7D4SE2ECT0AuEgelClHSgxIbIgHHQ+XJxszRFWjH3xXTZBHDE+WuKUDVE
pZZlX1muNXUIpdPi6sZbNTWvBN5UkDh1dGYPMDn1rCZbXI58M8pY6a7uSBCWak0EZrW+UYHL0xKz
hK7+Ku970NEEOL2tuOn3Cq6jxrlr1uVBbbbZMVLEZRARBlBuPUwfaKklm6zu3rey0+jV859rZEf/
3tK3dLUxY8dM7hCR5KgWgGWW1cCbkuEYugo+CynhZVijxYWyKi7qB2192yNPU7L8MSM8zLy/zVuU
8F/Y4RHg4zNbGzf8g3p4bXSzRO1zOo/ukiMKCdNmWY4NBkfV5NHGAA+IAN9lVD3XvbuJz9Kdtj3F
cyhriDiVT3x3grgu0V/f4Y1pbSonPtErlAt2rJ9mfd6dxzV9nR4nuDCFpip7hJkLjMx4wtpFNEJd
HzU50GMXKN8Tgmca+Eh5QP/aznEQjAIT+qCotjZCJiG5WVzgLlRWTr2Z5hqVvSnXHVHJmxhCzqHe
uOi/ZzF5LNwEl2KyWujvK1RnKQD84yruib83X4ErlLhnoXZdTsof+1BirREMqWEn2W18LR4UCfue
pUHwgMmaShqKtid5Afw4dtxjD5NRa+VF1Ha/jd2SLXZww2daPLgZpdydL2cbXVZTw8Nyi/QnUONk
k5ZrCJjx9wd7asYaGMHG4Mak7y9yAwOB94laG5fgP1Dg4Ne43z0kShbDWPZsf6smr0rO5qPWrKBw
gOfP+Q3bYvWpdu4ELZiC6cnfc0Zv9sm2SKLa7sJCoXS997/wnKyigGlVhpaJutwCsvaUj/mnx4m8
3Gur3UPvsbv/W2+5pORbfj4aIfoxQSsAXfb7a5Zb57mCeocV95JdAm3LHExSW7wJco2XT9gYCQ7e
8dKzlpCsSO9oVv6Rn6nZOskYYwfRQXZjlYpUt6fKfC49oKKk/i2m05GZpCEmpPkO7BaOaQdFc05h
xt1FTYuHckAqXqvlreX8oWmhMPYEG8pOMma9ptnzCMdBgxNCrXQTVCWc25pGE+Ck9f5D1+GwN9ag
8y0baQW93lSTzk8UUCgx5uMs2w0vwvvt18zC70V60vLwF8/1cyBSRuqBNJRjLqaaPPYUT7A3GrPG
NFnkvY9eNRcL8azHHCi6y/xjjhSxnMh0T2+Oq8CsMa65+93iTrTRLzz+FPGfh/D3J8jQfR5U36/p
RX0tZDQRVvBwMURiMbiNWolZiv8m55bTeXn2/BhxyfalkMZGjfxHyMqmH8puvcxhK2k3ezZOhBLr
5x7dt79vEQlSWi1i1u86cnsjQ3cgbULr+pIDDUjRHpChjWixodcdZGJxcMzvGWAq+b2xyji6ivEy
q/FoW/kafkbybc4mceCoCOpJufqibqL3g6cKSgoIBaGci20ptQ7S5vWEjNeMNWKSHeCfATJuTsL8
aLtiXFuZ2nz9ZPlurq0kE9FGO7OF5uOQvce+Y6VomLvbsljVf4LWYWMcnsc88fqtSAh+TKb0bmi3
AqvObl/NfQ+ikYMn1H0cAXm/4WZ2qGPbRGST/Tl+W6I3mqCVba0mV38b71GttvvL4YaspEtMW+41
43Mq4Tqi8xm8jt0GHpyovYWGpr7bqG1H6PfsnmglcX94ih4xeH9KtLw+jHsBVPWh3Oqb+WoeTnY7
2XIZPZ2MTHK8SYe7GsEAYnYGZJfEdy8a4AQTKBK43VgrPt0GBTuYMrnwh05Tw+JKXm/qs97MPAho
KQ3UhhufyFHokbjnKhnLSLzE69O9n3h87govgyzIQM/MC1VMvE8r2FqqxgKUxrWIWV6yCV8Kc6Ft
UTt1ss8vNVzq9QllHRfiSP7ozHOZkrmKQ+IRRd/UtCZrXByaRe3kmQQzBoIyDhFKBo5wxj/uKdpI
/DWHydmOUMvGSL0tm+urd0ZrxYGET6ywpUeYbrhcyTE3blzF8rR1JcpwTsw1X/guBzM11Dz+d2Z/
4ccAH4CGtITakHbO9Pue2pd/R8Rr+PIlbBoCATZ2JHX5qaXAQS/12rmPYVW7IyNu47YczR8qagPh
Zci3kmnmXEMtkJkinSfr9JBc7VbTlIj8cwwKr80Ng/fxNHQZ9VVNeBGP06P2FYOUjzNBl3s8FTAE
0MjYNlpm/BM6x1tlHIt+ehwsPMjM+r7yqQJRsX9QCSeeQuPUca8i8MWvzW+DT2JrXaTdo06o2eY5
+BOOzCy8+y6NjTsAOvcwiAKMS97fRJPF1H8YV+okVgrBlqw9RgthNmHgIBs5mUFF0ITiKH7/H50D
2hn3/OaCGJmDRGdXZLvHkcxvqutUsm7frkWJ3RVPSozX5dnNvvSYoyQ9f2j/jTK1w9dKotBxmt4V
5kO+GCvl/DZFD3ACODXyAVnDrHzgwrMNanqoda728/xEl7f4klgy2F8fnWkNqfoKSCykiG9xLNRE
JjVWRI/vucbXWPFaaASPjwKaj4CMvvppCsczO080agOsYvd4HImpOo/yG94UwuAmPjTyMjMqEN+Q
eDQU3DHHSBcgJ7b581SFjScgwCAtcn7CF1Ha5pOxcReNEyusEnbd1X7qMg4nTjzOI3pHp2FSus1n
SH1TuqEx58D8lnZCoxlUMuYIS67DBmrF2HCqz3DvRNTGd1KBnWX28vV/2sLavX4f+ANzJt1DV/A8
nBADq//ZjaWFU470BTB0K1Q/+ZtFT7Y1v4m3uWn/hbT5SpWKxM+SPHpc66X90cw7Robd3dy/VzWM
xJtzqMv9DlfVsiFaU8HpYDdFk44MTO7/177hfVMo/paTEsDq5GLRTK1HW2j452CYJ8SxNJeAR48p
rtkYpryhFsWo4TgwB1QjqIg9M017dFYlXkFDt/kVE6T1rA/W6NCEspG7wcSU+FWIxOpMp3U2gyXw
WgIH3FblRBimYukCcTN3LgW44HZ8LEr3Z+BPI6uP72qMTGQj89DTPgkzBbfP3hhVWe2GGUirS+17
6Une0KEeI9rzLxSl9SVaH+j8u9Qikcv9b3vjaFpTrNf33VVgsbItKEOFBrGU4vgw4OqJT49oy65v
SPbjNPtbiZI5v6P9VNaNRHgb252M0IsNUFAOZhtUK6zCto0pY0WE/3Z3PUX3vn0K+RdRd6vSVKtu
bHew1ULB8C1rRAoo8DffF/gpuTLVPucGrlFUf+8/zfRzL8eAe1qgtmwbloEq5C58hBBaiq+zKL09
AsghrQKLM098ec3bFt7SRWieSAT26LSqru5KDEhadceYprhv5WHtxvZM1Wfix042gGE/UQAt0Xcw
NVFuxPbpzDjx3ZsUhlqkVCKGk7LccA75hZzTSBcnfDgcOYpKPxVARIuBJmhS0s7NczqMNI7+Wt9l
5twZPWSrUE7mBqCaY4jaaX4Co5vmQCcWddDYWwvbaDOlFA1h7gJqzPWSHz284LLdCcmCFxTJbwsB
MawhtVwhxCRAs6PMxiBKj8S5+k+WJePZ7D9ZG/LoXOnDh22pIC8T3MWwcqCbe25vpevFeWKQvlMC
EYBFOo6KSWqFmhic70DNHs8THcRjKWgYpfRygq2X4AGRIa5tvq6AdKcCzSTseGVgR5OPZDglWIAb
IoQ+kB/W20fB0IcElSJYYhtn9HTsx9C8lMv/uvf+umq2zDZL4C5zpPrSTRsWwWVKNNOIpC686MFV
aN2s+zDNGIbchiMCZEDsKTKAsQWfWK4g0uMQesSODZh7AIObhOMXLPMUe4nhf1ZPeXcEGvHXbmSX
J8J/G4fHKg1ZTQuGH2oXvm7WXHOl7CPSqW+BAREenWJxEdSRFP49Y5yrUAVwLOB+Uh7DmHIChn+s
QKbwozU8DPBdbnvj5W7kXabpmrqj7VIXTDR0uvjkB98U5IzhHgfWrsXKIQ+tMJfOonJBBBZt/YBz
Sjm4jH37Ap4XHCXooxnIRQ72hVci8Xc9bblDHLmF7G9hn1Em/bO+ZRAIzylP3xWP5Yr4xEQZ/XBr
PHmlrCnmiqsQaepr6b2Ijy+YIAC8fiBcDDBjvljrb76YTBuTPobNlJHYmcjhZJLkjrVZrE6RHRQ8
eq7nWZhbMXZIb4oDC59fVIf6cWEETh3DFpinBbU5fmNcWZK1lTZwLVQEtazQlMPtwXP8aGFoOjhb
+XkeAns0KDvwZiW+oj9mhvK6Sag99fV2Vip2nJb/ItJP+Pc6o+aepLQGBrf0Dxlo2H/qBkT+2xl9
Oj70pZWtnthi1/2UbJ9ldkQxFPBj8sUQsoj3TcMpe4Uyfuff5yGdcaUm4Y3vvGSCInk6q0ag1Qpz
bAcQzQYXm/iw80nWrjS1VecAEW331dhPs5cgXGipPGTYm1miydkxJF5okyrNN1SgY82RZrnL1BYc
z4NiX/BSTrrPR5lvJba4GRBH16CWbFnLb8fXLHC1g4gC2c6pFyBkMBKAB8uMBOO/x/R2VeAPzzVz
38gwqBKMCiAvBYOVZgiutRAmyCoGQMpSbfYvow+1Vj2ywipj8wEuwSeq/wewkHee4VGDCEYUYvVL
HTnEMH8c6e2a1aWa/FZU9y0Wi2H2LZdaiW3oWP3lujFaGNGNxRcwlyHm7uOfwRmLbOpE+3yHMKfW
1pUbEGcPSq1wM1rW6MkBOwe8cayWd87NaCzl3kKNDySn3pvMSqdeJbkM9ER/wuDyRcOCmbom3pWF
NTjp7YoySQMUUgPbbxeCvpQksJ8T4Cc9xuTkAZ9dD+dkXX7sZ94z7F/rq7Xrdv47J8w1SjZsWJXL
JpBTHva/bYkOiINAmYTuYziwYiIg7UEE/oFsUYJGq6VeuabggjGWIl8O75KqgwY0cRCdbhqEuKbO
+Ib8rbbQ5VMCB3/1NXBanEmON0M7o+vlY37mVOFLV2CKJC/2qjQrQSv0DYPtRr9S55aBl+Gbnu98
Ci5IQ8Qp3X7c2uwJhsAEVehz5uaH4fAY0MRtgbZJmGd0QM8NeQ+8rhkpij1aaXkgK92CngFZRQgu
PvG4GcNYIbbvdBUdiZIIh78X0cWRlBKIl9T/LReAqIMBal9vbcbEDG+ME8DWbxcqEsHXgaF835IU
nOQLZ8gUd5QW2ZuclJ6CZpG7U2AQoD2qiupUS7AT3XIgA9555EF1WpA27XPLpGplrOsj8UuuL8bZ
qB0umEZQcwMnPcYNCzjSh6PtQBTnX/8vZi5MvwTKbXssXWWLL2kyO0nyNRuaV3k26RBOq5rSKb8H
xOUfxrobeSjN7jyaWYCbzAOcMZpOdw8haaBSc9aRll6ZTpew4QPju2CxafFlgxufy4mal8uOyIf+
bBS+1dSId38vSOFNpSPrOjsTTBexNNKGYDP2kT4ZhsgQPxFd74h06g2FUfCuTVm3rRnjZ1SDppC/
i6+AEhuzuP1m4BUd8W/LqsB4mGwUkHjcN/6LSQd+uDA7jxx5YQ1bSFutDBDtOLT25tph8eBnN+l5
Il1bMrn/K15fgOa33D7l3a7jmtKQ40h66CQJpEa60eXbJQtwG2jzwQlyk/gbG5TEyNeSjXk5kd99
56O5wzgzULV5ONs0r0JB3Wox42IHlWbBL6uKbb8mxSohFgyw1EeSvMBhA7sVu8wn4pL/QP2fvRHS
QeWIapOVew4l5/nFBv7Fzeh3cu/RnUQPOxRNPey700JgItcD9ORa6O/WIxmemUjI3M//+vA/HJ32
PMstkUUdkPpbdYj3AsA/c1V7+5JMvCKf6Yi/1yxqRlld5jFaqHEVNVuwAhpZRhgZUHzKXhkP18/6
qWy1iBW4ZrGQ1jKoqqPueYSnBSnEhDxrhLAqPeBlN86s/UEOtkJYnp3Q7DQ7Cw0r1UZrGgN6HGEA
lvYx8S2bqm6BArmMGK7cw2xelO2E045fsimBMRLlMrwes7Rs5BngFu3EIhu+R7/w/EbifKJ0cvqT
VJ8upjuHxvjCqD4kHIBGTmjBIuB/6/qFvGJurIzXSlexCDO0vDgJmO7HZpH5/McdOOsf3nC2w3zy
9soX/wOYf5PtKACXQ1m3GTjTux3D0hh5MVhKxIFhsM4C3N7qy2+xXB7nVROrWrZ751kZn6sTySW4
po4/XgmxofDVJHVsK7ZCQmE7ViliTkZP72RSm45j5UT16talp7Zu98sHvCAO4qVcf24jWBS5uIuK
SqmXpEU9KdeMgZxybzRhuIS5NUZBu84MKsMIO541s2koS91/D643Lsw8n9tYV4cGNahghZsxpe7s
+W9/vYI92M0B9eFJPFgtSPmcWcjqta/bTz6HBLReeI2dsrNkiqE2ajvWZ3A7cCZs39zGIKAytSEj
Fc2Aq1IW/ewFPc2a+r7UbJDY9twAWTUgdDpggovQxjtlykZruObDXiXHjFjeFoRn5Dnf5sD9PGjj
JPS8qk7/F2c9rhNhUTBUIaTVsW4o0GdKX0ZmqukjIWnHz3L/nfXlupBQYMb5JJOmzRbVTP+suXUY
cXRoNnLjyH1Zb/rj30W8dFZlUILZX7BXzMgZ/DlU1Ey1ep/BZT2iW9RRKhSGOntCDulG5jltXHQZ
Tik+GxIMiikNApzi7GdATnZ68vCebpXLZ32gRrkJi2Qo1OW7uc1VozqvANGatGbUEvoA7Hsiykk2
7gRuApNkU79/RrhNd6zVB+ZJESgZVe2SPwzIF57eTkVljuLdk74a9w9Qe9KPXsX5UCdulOyHDvUv
AbgsIpFWayY7lKCHlk5SpX7S8W1A6RmfmlcnfUcJ0oKL9QrlXbFSmscZ6K6FauoRn7/+DGeNeeRH
n8u/Alwpro+TqwSDwmDFp+9P6fpi3TEt1lcf/U/A/bU3iLbwc39y55hcdvwx95sxZvaODGoJ17tJ
zAz3DwxcSPsnIdq94UbDzaSdYrZ1N2uYVqmavRPK+HEP/8TJ+tghQ915zlTtW/aYknroUvWCEDhM
i3CrvvLXpUs3OtijjvTihab64eiLs5L2GOzLCfUntDwvimKvlKTdq0y9S3/wao9p6pFWAsdGoCe/
jCy7sgJUzKimN8aTHVX+cH+S5B/A9sfY8wkSCJt31xNIHpymOd6DSos5WhnLTactQ1vmDKoGubEe
3hqZBvlW/usA2i7D/JvruZ9IePGU16r39Vg+tR5hLUxGsZlWESkRC39Umo/20zgO9GNhzZLKYUPu
awtE1ya3zMAeVFYRUr69Nj166VL/Dv61ePIiqcWNIcZxjItsPi0Je5p9K8gbqUpu4rc5aQVWPzr1
50mZiZsREo4XxGVQ2KoRvg84LC5Er5JsVhU8xil77mpHWtxsGOfBJEZbl4iYYu4yA+XNBjLNEUhX
efTmxRvBlWGr1EYOyznQBb/PoFXCKwKXORNkPMAg0cVb+Dk5oiqKKIdttn86ZvtJW1zBHUoAm4vi
m14r4bg9SldX9MPZVsYv5LresbOzcbAXeNb8gFdoiDoqXx2mIdPNocebM5ySuM7Lmsm1MULrvT7T
RVkKDyJtSAMmFiODQLSUhji/xZMSDCHGoncIno7sR4gqykZG8FB9X+jLXnPSz6qHrAGwu3ljYgjL
TdlstGvLvtpajoM4F3FET8+nBIeaIFtg6Hxw9HpP+zZX9feEM6ibsuEvNyFLIz+Z1OVAwXc5fnJT
Y+KHVt08yW8GYeCLnMGiX9GO2QoRF714K7BCHdDtdfHxCAWFARwr+eIhoEaikKAsnLUYHc2b16rA
ciudjUbS6CvX+6IHxEKipRn+Dr13bAsrseCElmYWpc8tvgy2w0FoMj3BiTjw1waCB4j3b6ane1TB
wt4iI9Xzn+GGhHn/Czi6gIhi/91Zt61mMK6f4pAvYGW9if5Ayk96oJP9DqSSTQIgwy3WevL5FvyW
ioRpiVGY4Nd2EdvXSHGoBrzpWSwbeI67BVlSlQCP2ZVum81GlZorQWzKE4h+RXpl0FJztsgrD0V7
HI7sBxH/CGSDEdL/bw5RNXCJItH1qnWjLsQ2Y0auasyPE4/2Gw0W0XhjgVdRZXauYujMNVwUEZLB
QYizKUDKZj5h1L92vIyRblsZQ609Qj4mVlan5+DgQgJp9B/rWeAOTAyoE3uTbaZ+m7qAbG00bhEi
gdTVGY7Yv9R6PspzTo/VEbb04VFG1uNgDeCx5hbQ0toeUN+0nmrCO/uXFQuCCM+volDD6MgKSYHF
ZqyMVRKpwuNFNIcMxY2Ib+wm/UlzNLt25QpXkzDNs1YrjjG6xqY4H+QaHYBe41RhpmNTwWhrL5jK
2B1E/fLREZ4Iu31Vb4PaTXhNOKkzBwRb+oJhobNBs4Y+aggXv9dFRfYpTT94Z+/YZsX9OrYvoU+2
oauz7159VtlDR7WTNKx0voyuffeWN1OTelpX3El9m38x2tMsKBeZiQUXF9AUSvJxubpPuAP9CfnH
Gxkzj+2t9prmrr+Emgc12hwPjLcu5tQfQNKEiQ5HWHg3V5u/M3dQyThecWz/i0UHCnnaLpE/Xm/J
JisGi19fTiXs6lH5Ca956zIup7C8JYRrAcj+iLaWI+9lWtMOnUhk5BF/b1r05cWof4yK0DEen1Rp
euiuFukeqe0bgiSk0r6u+Q+1UtBD74ti6Aw/j5wGewpS3abjZ+8OXLzpGubB8oPa4AIc47C7xwBH
V6pO1ecgum8k28nhO7QKbdEV4hSbzbVofzvcOAXRcmdxXlh0rWSYlnQWYGlaHBk7ANXz3A47HAlq
TtdP5X+/ReNgpWuZR+ZErF9mEFI1uHkLhBZ6+b9/jCeUXnUaIca3tNmke5cqw+iwfy4BlBAoOxgQ
dOVjtUKmyU0JzGlbSYJCJDnkRFjLFpFPx8YApHs2RZi8DXrUjRJXfSLbIDJNlKoM5ov3rtgq5iBB
PgxmnOsICj6zQXZuFZjz1n4eR/0ycsnCsvfU1ACUU4DNIbCCizpSDQ+iCCmYXbsIEZEtd7f7Mu3h
OFLCTbHq7IjFVdIzl1qIvciD69cr+l+XRjjmqQrAq7ivxPIRqk/qLrZePIMThwMAq1CvEcBkfg7c
1SmrtSxlN2VDIVxa4MxF+b/3oSobDwEVnCgqx4Z6z08RxRwCh2+ToFwnH+VB7KRgQq4Ar2KM7zYh
nx8MxsvgtSXzVRwnC2TU4Z2hgFSjiBoodVLLD1+Cjts+DVifKr2rcVfJnbAdGI9qNL2Dr1nt/8eu
QWsV0A6CDqxj3wOoarDV8g6p3z5MIfNEgw3uGOZrke1n7Yz3Jay94jeyrLw0jeHZ/f5w9SxrMUNa
pL/FXfZNUMTQd/F68ZyynUUJmP5C24aepL05suzXtEITZV5d6M0CgdKJ5a6MvzvzNLGk6/CHeKL/
cqPbFTOIkEDWL9xrNlOPAyFhfL5afdup3SJ19eovTGRe0rKQ1/jsXXS1MxDOe5LItLyXa4hIwaBV
eIKKl33cEk+HOIftJApwLY82ULZumY8WfWyi5/5svaquswyz65P/OoAfvQcxvVy7C1Fgpius8Ydg
p1ZCmqQ9BjbAEs+hkbjLY5vuSig+XnJid7O7sR/rbasJOsw5q0cQiIkW4sBxTybcXeSuRFQ2dmil
P4D//0S/Up9oFmXqIL6SfzRvWc5YOrk9kJZOIbreIi+Pz9QBmgBhtQxo60fBlY77g7e73c8zoBgW
mdvVm0KHIoCSVHN9SxV19E7flsyxLxA6CZmNsv9y7nuRHrTNti2Ny5MYeQ3uL0QrtahcaY/kR1pQ
I+lxkrpK08Kan6e0Xeh9Sip0mC7sgpuM3J3zorIBoiQJsUDOZo3HiUyqbRqyk7AAAiELOeCsN73E
FGTsI3e4u/A6leAQBg6RscDVrmL6jpJZRvY/wh3QVLximEBbKaTRoqJYBx3tBGxnTSombooE4roW
URwcPrqrYunJ2LJ8cbZ7LsxD15t0OeDmTTmF36uaUhmzGy+nqfYnt6pCodINDVyWuZ1CiE3TQxal
ekIHSaKZ01NlgaCPuu3uDVaVjzD8cLIviIJ1kqvALyQGfg0ej4jo2krlRe9NJDNT7Rx9yiIwKMi0
pf3CmZJR+HY9EnTm9rnbWIK97cyQArGB4yG+5OiV8zBJzWXZ9XXL+t3xaaIBtEytpgh+xQHFGDTj
MiNQQQjJzuWuJfTEXAHBTT4ihZN4BH2922z+7ieJs2PixH9YhrUEWu6wbH6DUCA2ZeZsMA9xVJH4
OwUAK+HFKMytF80UdEFNY2AgUb03Y7ehZB+7XeMRkdw7nBL2k1e9zg5EvOcByKifKq3oR5ren7sv
kA3kER9Ke0HNvGZ4O7oUfT13WHpOlW1AvKIJrxPWtXkpT0PN3GekvCZgvbdPWO5AFRAYlMuQr7ag
cWgnnOexNM+G55q0+8/kQkZyuJTQHl1mdpOUUSRR2fQXwBEzNP3eUeXILP0i3Wl66V9rINCh3geJ
GnZBa6WcuLgCS6L/KFGmWZWkoD1oCu7j54BsIxKcTJl8UlasoncyuaxLBVnMUF5CcxfVkPTNZHtk
y1xeJSgTBl+tWRqguooASGw4xrDP02vSY8IyXhCu/rQjrBwv2isa+8ws0Ougv0ajGkzuNXl+okDL
mwWzytC8BPq5kTjSedL1Z2JnjpM1IJdcH0nUZADstAjTNg2eP+FmoNAaze/ppwCq0lD2g0Xhaqst
qwPGdXtjAu3MEwLq8Vv4aesS0qQc2jMqocUrd3C0Sg0b4iu2+5+BbfgMdZ5G6q7Wc+jKUdP3jJPj
15smWhfLCoZ8z4U2VqTfeZrN1ID8pRpTJl0YD7Gyto6HLzEss/nke9H506PjmSltk2ShEsUnXvxf
hbJs7dgpgNyaXP1Rcl+wGYHbWwWHnPwaSofhCipzRD2dtb2GPDaE4WaSb10XcBMRTXtItizr/ofP
oTbteQ1n8jIU3zvSqG92G7yM8ckKprUVlicPqA9Kikz/xw/gD+l3hKDnisXRkHcLyP4yGj6D2w3L
HfnNPzz8bIFYPxMvzS8Y1flrl5TSwwBeasWZC5dhYPu2Z81NQ3AJGDipMwXLnFZA/02TCYDzVjBo
I5AATBLq8+cr/tK/kCvXuxbNt07COmn4Tk0l3ZQvgTRlNo9fPYqTZ26wgl0ocvF+gTvQFm+kK41N
X/s5qEvuOPYqAnMT5tktgTz8Ip4/XCxNHKpGaiuB6cI5SL1rTVCA00af8htTSORkJwzMSf8lgu0f
GL2x9pZZWsq5Td5RectXo7qhFNFNMgf3T0joDjOs4FV8bk/Y64AdQjmKZ/FBguJFBOq0VGgL2P2a
TZlo0LiYsfA/9mWlVEwej3kCsrqmqJW3dUaq3swnGT/Tnovmx1qmByy+v+44FTaoTd3TP/3sMDXL
1fuqeDX1r9229BCtwm7YRSuXMC4MDw7dgSjleERdUrt9s3lm7y03+DCaDpVLyis9GKpvCUg72Oxw
thxojPyhRn3pDWl/SLm5FLce+04zu8XwuOBUQ3+1+Q5F1Wdh4xDdRuROSZRYRgy2UjpC9aD3Geqt
zVpCZZQx2HXJeeYWNMPp3WXLYqFVQjEN78i8+VJUlujsJeUZjaO99pCQrrks68cgpU2ge+L1Mn5s
FdkRazedi2WzFzmgimbXnbfpqJ4N0I9+DZi9DLHMHLgvM2Ey+cZ59eStHtg2L0MthRje5/Xvuubx
75AWHFOz0sxBZ6qFibPwxGpZpnlqVGp+qhah7ey+sE/PZJX8aSEQE2ZpwQ5W2dFWumaFO6bHu+Rx
xuGeI7rPjL1wySLfojMxdc87qc0KMKIeZgwSHOkAvyv4HkOKAYn4sYkH0zq4hIYNWPv16XVm8bEl
C6otyNPFMGOWG2cX60iTlDMcljUB+sPyRBLjvYKxEWq7eMcpw6/q9YI47XCvqvpVPZEmEwnN/iQv
0MnaPz3kkoBUlP3gkChcymqj5KCCFKmy970VEIixKWjfarJIJc5w5WhV5TJacBSpDmgUieNcFiRV
V6U1fhjkeRURzlSJUZ/pOaXe6i1Le0eW1E6ZBWL7Q/iLc4DMTyqhQ50ccnbDyyLZDciQY2R1RKxZ
g9e2rSzZUSH3mFCr0Mbw38GrROw+5H3Zh5EO2HoVr2TYRmfSN45xN3NGZ1MVtgsQj9OoLBB3BuCE
X5HC4tz64bjMJ4d+zYbS7tPnwaCCpRAWU/wxFeMADtJmZXeWx3DVNIil6qxMEO9yYkIe2rLT/HOi
TT3CX6gBfQuiSaCP9FoyCsasM5IWyC0PUHYv4jpudt333dJSzr105Lek1CZGJKNEPuGXHzDMhWsr
P1v1KxmOe/kVEToDx9TtI0GtSvdTOzLtekgvkf69ObadSwTKu7JIRlHF/zwtdRo6xLDhQtcIkHZD
6ocBlUktzLZyIqebtjrQg0pImZ9xq4dXOdubnVHEuI1SEXL9t2hKDjaMeQVJYj9423kRhBMNerGs
es+O1VPK193xxlsuK52jCnjf4TUBzyRU5XHmxAi76FRgji9ouRDhSlTpXvtb3GzBUBngNBUlhXiu
qPWcCHuL5mEMuqWIcL1dk59vJJEcpjcqnr4JjXS9vM9GaLjmcErR+rGSW5mgeV3B+HxAU32lRpAK
Xj6ZZEfsQ1JnG0Gv5DbuxS0bvd8YU+KCtoDZSww5AcfJatg2s+VgksUZ1q8h5Tx0XMcIZC/Hyz+z
wov22FNBH2TuEtALozb7hh8MsjRvBkZgind9MAL24fQH9C1cMZ2R7L1Z+J0sgvGoKUzo3maJBbyP
dRDDTwICrJejE1SmO+Ko/xo64xL2A7M84QNhTEpqHK5PZ/m/PzLYzwd5qIAQf14TMYbpjJs/0LND
lFxyhWR+O0IpKe6EzurXqJFImyj5aVyNDlqKYKkqfETiFAIPlIr9XiAVYITySDGhcKQU8m3JrUjU
kdWeKZ5cBvpfv7kBaqbxhA5rX6355AvBFqzNu3LPSvC1w7csDiUKzyh4dYo7fYIlcZA7Dqpa7iIJ
74Rs2YKPIf9d4ONh/HGcYE+oz3/nNGlGCzoiUmgZ5Tpegt7MZMWDn820yWOTHNCzN52bsVDBYblq
saKlgNeY4TcK4yMqNfgj2X39qzz1mqN7/PQQcOxzO3mNbuyjwLAHtTI/3q3Jv3dWeC2C8vuy3YZ5
PigkdXFW/VUMZm76fZ0Y1UBTjhPBSrelA4w+eVuQ7tk7Rp/nEIR+X7uq1+9rCFmNIUyYNS7w+UAo
pXZzrGSPaS4QfmFKNVZ5QD39EDtexMwrzYgO2lWRdgQpzeZYxPfw4O9MvrGmpYBSBLKWkDDGCvF8
REMt7NDYkD4F5EIy1yV8VGiusHOYxJsq4BrGbbRMQjaKMUEsKNNSOnhG9H+2T5K4yWaTcdPOOYVQ
SvkXMF8MNn+c7TAy/VEmFPZTJO+ZfmJxmCi0fTCbpFKeeeHjK4vVf/meCEWX91UFNuBPlN4MiPaM
ZIirp4h7kz4vAXy4uuZuVm1RctSPHffSv6K1ot2Go0zHPWp+DVBwFVo1Wv3PxhuTeeBAJovI/TKz
pOqExE00JeFhVKGF+VP9A8HBHDIL5XkenrC3R0eWo8Vi9PT18gfjibudTPWnDtd9gpHzKtcU74F1
6SJdnMZ7hbKJWVCRK1nHKHV+NoMQwSn5AU6ywifeKWElwSadaGPk1tp4Dsew8dMJd5ZU4Z526W1l
xQCDutH1Trtx4anGKcVBsyDS2c++wVlrP/56h9S4swM8STfFtKZVHLBVd2X/RQlvp4CSq03m7qnF
5svsiZujwSpAuqL3Qb8g4a3IcwD2d5272IiIUfZ5S12wXWg6XYDanGhwsLkS3Oj1UmTkNI5Ukatw
gwbt4XC/vOou45dNgoBA2DEZMG24djINhZcxbKY0wzMGxICemEoOOK3mz92aPkFZNKZIdg9Agt48
nIuqoGBu0vMLbGG0kYpn5/ZMQuzOvqoE0SDUO7f0WNURM3e5FTztG+mSKCWeBm/udxB8I6rTxvf/
ONK3c8IwltLBF8PvuGR4YXeKoYo02+VORvOjSQuSKssFczKCApG6sdVmBIHFZLny/ca0UROd93ai
YApXC5ADrRTD0hYvfrmzhbRKOIjECYYbDfdmaqqCtQmXjePslRmj8NMiOyk+PFc/8MrNmhBvy7wo
4mu7eeHtGZGWJc83WBnyb76B1vHlZ4UNQzsCZbiZaK3aFeVKqa5wuFDyibrHpKvDhOzQUNRRCgRE
ha9e1vBxNvGrhvh4c57P8dIKOW5REfq+d3j2K7qWyyBSUj1IC6VQgb/juAPlnR5rEHR6g6oeRPNP
+J0gAAiac6Lk8rjM+XxMKQ917tcEIbLRjTmNMX/Qu7q6gR+1Ul7vmn6sPkhC6accOruqRqXPpFjv
i20fgEf1/Uh/BKCjYFu6IvhfaayFZXc4V7CVoVlyQJpaG08A3nNsYlsQ5x+XCmhd8tFRztC++IJD
Qn8bApv2hhnHRzYY+1ovObXAegNryWqb3TmpIJEz1QfnEC+t5TSLYdSXDnFAPLvjJVEVOGbdOA8T
4HIYvxfJm4rPU+j0xkvZRbj/xMfA21Lg21YPengy1a54Isg7HMZW6AUsGuYiF7o/73K75Wh7UUCU
YMetIPh/j8OoqpRp+BCmus/N/8o2bO+qGiTSaEi+a1Lu/xF4K1YxHUHW4TGihV+LNh0s6RbNn12V
nHqh0DgwbZ9uZzOH3Mvx1hlKe2ea/wluOtBXO3K3W9U+rLxOdDxUrx1rtloMgB8j+QZMVLuvGN+a
MLUL4rIjAlKqVirxbcNwGR8qqvmDPIsEOPXY4KxI14GoX1/+RksXDLrhHSF2kRASYmhamcbMdHjY
Sb/ySKvCCTZ3TCoInCUCoeZwYzHVyASvFAeUCfRWRtLC7Ih5fSDVgGjz2v/oHj+ZVialUZ4sn4NB
zF2rg5GzzQP7TVaJjsgh21yvykwqIOrYnVcZYU2LLetvNgygvVhsXQPqkY0eBHiYRaxc6HV8sjXD
XdnYIpmIQ8hgeBMLzbz+qujudBAPaSK+eeJmSzZHP044qUlp5H+7f0khlW9lu8F3i6nRd3nP+ZSV
v0sL1KNG+Yh40Dhhqv8unrlR1xRH1jqrsuNX36S7NjxUpHfdrEKfy1IAaskcQILsg/SNbJtrUSbC
6WUFW65VTQ8jDzSl3g1EnaGJXiSgvRtZJ6B10/52R+xqV22bYNX7g8dOIyZI+kdorl/tuju4WXid
E9kTKeyiNTC8isK0HktMtS/ylGSJrFo7JPhaalrZZw/Njc01PnMezT6FEp8qKA5J9b6qlFXQ9Tsr
3Cw43WOgWbpv+w8gALzvkVtuSnPZsHPDfN3IVd8dZkUlDIxWa+4W09GNuKfiGXVeV432GASvWe+O
AmEADfdM+LSHS+FkJOgCstucuwHi3MW2wWCn7Ybx1aoJjMPO9FxTqLn8AdRGDC9qwAc9uGmIgZnm
zp+Aadfr+vJCyxYeGuxWrvF/MbgO3eiBIySrZZTXA5GIbZCAeYixu4gFiHTJDHGbAj+LSRTTzG8s
WyTGjBPsEQYEI1ighJkSn+HMfY0jZZujujloAavBxxQCKK9HrJ2TgbgeYVwd99W8C7FiiCwHii2K
GjDUGJu6JBtXHo78lUaDKK+tT5/7YWKBTKjUUX/r4xY4/1kA7nY27falb+Ed+sgqVRcP+xajUuzD
PJJjadkL1iDwSzlxodU5bC7O3OFNNgr1zyKWIwxW1T8oHLVNsWQhORun/DLNfSdwwa54myncTeZi
KLkcCpCs7ht69llDRbCiKa0nqsFnQGuSedhtV2x/jlFoQqd4wKDRv7opGdIeCrLdDCLqoIiC8TsM
qC50WRxs1prQ1Hl8ZHh/lGyvDLzNn2jikuXHc9qE6UsEiA+vzKfkY5tX+VqZZv7iU/72Ee9k040/
dzAsRIIFPjOdtI+Rgm/4Qp2DVpoQnDVjJT9Du7/DwIiaUTNBrHJH/6ZkvCr5KWQELu+W5D6zNOwY
22wxJ896HMwdqRkwaTFQL9NABsLQulGfpx+sKuWPKcBXJAP6NAN2wtxIfYnBmDkIRJXtPwT+yGRJ
OrQlha1Kqyz7zfB85TnxevevxEKKvnn3XMytOrKkUDnb306S2Fdet162v2t9rgZyF6sk2RmmzQp5
3FuNw2hGgHwkm2FMH/dzbwST3I+88G4PyiIf8LIiQSCws5OggYes/cFpDIpXwzmU5BLohvUnqP8A
JsGjERTidk/VEWlwAyZGAd1ZT70PdL3zRjztflH01KIz2U2sZHt/N+6cM4+6quwPgvJJXvnAfxdO
hMkVJqrEBmLajKPqULvHIa6/rgtweau3PFbt5tIPunbZtT/aGw50VHPrJT5pGwpUh1XxLjyNi4Xq
/lDcnHDs5c5rMvl/mguAniuyW39KJs7QeHf0JURVVZ/4uw2Jn4gQFYgzfaGseLTkz5zuq8ImGLEF
9Xxpaaf4l0CTL+Egea3ORx1VBdsDcBL/eQENH5Kzd71f9Ky8hZmKdwvBDJFsU1obRTIxXaVJuMx/
xSsI9XP8lcGd7e7+3Pm2M7uml64thJ2f7rw0Nc8yxI2z4YQEMQnjWD2wZj7uhEvmvOUJ+sdNufDg
L2FQ81II3wkDIWHGQiaL8WJZeQqXGuBLSGdKpvB72l+nd3GplKuH3Hp4ojQNwDxPmHaZBCtTpK2F
VWXx+tvDszxtfUBGWTZj+0ThC0APtY4v10YJHiyjX6OrKLpS5egKDod2aPBMwGdmyQDJ5IIHcjni
4vWrO22DzLHDy5u/+uNQmUOcmUhQkBVa09dprKUWDM/U1nDHpggVhlSjOxIHYLKba6tRet8mcXfd
X3a7KQ1fyzuOoGFE0M2kg+mf97LAqI/WW5tfw/qmLyyBpYIUDys7zfuwYY/OnINXQOARSYM0KR3f
JCmP3pI42nqDiQDFhIjUMwX4htLyI2p35Op60acWN3rKJVRGQy0lQ874NybE7o5/6dVzmuIt97+Y
QCjdZugdU9WoBov4E3tSfYAVGjNdjCT9qbABwm2Un5IavVlm833I9QEFTMeOPRm17RJsBzmGExIE
0uNizgq3Djz59NpkDcibMUk+gBpSFhtwX1ptGdgKooRBWXooAfWnXCaJHHeRcqqeTsgr6trxMXfr
6BGHuZwo2y4bqOvlNtkmSlXNRUIHEPtVsoxdFmUqQdynWWsWQFr99GUrMJjsZMEnP0loDgKGwQXF
KefkH1LO9iR1/TUfatFoqdxfcSECAnWqP7whRPLE/qUknwAYJjtB9EtmfCyXVLIG55c7jBPni2/I
Gy/ydfgk5ZWGDEeiT9sGO0zULeJFwLSN6g41K2Kwn2zVRfNr8yXFuPOVT4BLRO2u6RK8Vxu+FbWh
BTtTRQiHfejLjktRY7P0kdiQlJotNQuko+3yTfvZJPTdHzlD4QFPx+w7BqCwicS1bQGrGr4/+sta
JXUfno90ZGxng2NBAUzxJNYzIF/Ihq6idPnSIKEYm2fFxfVeFgUcwlGf3ORRAPYThYikqMT+aWrt
o885s1dZwSns7hoIj3ROHQtiJageNGv3fkgmcw5PxVq1jjQfFi/MfssNkvzOjmRslchH8vNtbkH0
wwjm0+hbuFlfvLtK1+pA6Cz1HF7MiV5g/zzWJSBaGFmnfZWrsRYWNCv5f/W6JwAC9BeS4TLZc+LJ
ZSjnbnmcV+zGIqUe/Rizm8JvPGtupdrhidDXEHc6fslkW0QqN3zL5K8VpFsjsdcbZcyfFrjY1nRD
qfAv0+rGeMR5hXd0W3YNqHhySy49Z+uXW8qJRwRLrPFASPkl9zl7wn2oNwS4itUruDQswsoOmEQ/
YE+1HqFIqVXqQwzA2GPeZj7vnXjvrOFjKMOROhOWXtWJkCQ6JAhZT4B2DeCvD0AKcUKK6QMmBsD2
IVEZ+9iQ8nrm1X1ywUbk5vG9xpg/911yhsdQLXaadwcRri7rXcMHUnXlLD3GaVxI2CHbre/fxEqJ
uhp57YYWRPHa5U0CEyOleFWvyfjQIAMZzaLQdbA6LoJ5DAgqEZByPDIlq43YfRSyeSCkWgXeXnkS
YUWOBj8ve3TB+c2FDe+USjuPxiUiJX0VrPNfzW9r59puQ4OXrU6WYEeObEOCRqqGH2GUXNjdQqsL
SUFGBOsi6HKT7ml8sxlbFSb4nnjNJWCbysKf2xlaDHF0xEndMuhbTN2nYu5KCKqLP47h8tiMY65o
2x5xjtRsVydD9J7aI+l3K7ENF3Ce3BlL9kc9HN3wrFN84o3rcAv3EELeuzDIL0lOXoKK68Ddl8yZ
DwudMim6HzkWPHXNxo5O+AO/TVQ8R9D5lBYEuqPIiLH7xb5OxLeoUw7gZNy1+TaOkjVmV0ODlEwF
V5X4WevV8lf/PwBSn7lxu1hcF3QbgxSFWdmiPGNc7veoKTkush3J+A4yWJyWZQCHcPsJljIo7Mix
aBcv12Q/vCJEX9mbeJv8Pafjvs0wLs2Mo09JqEVtELjRhhLKJjFwg/O9ABbvcQla7x/C3eAtkLgG
ejyxE2+8bS1xDlnkYECHyY/9SqFSNz/euuUnrzGsV9z/mF5aNIScWsNR3gNFOd7sMHi2W79nfDYN
15vzj9ToXcLsNFPMvWNgMb5C50C4E4hC1XkDw1hTkB4iKWjmcV575J/Vdy3VwEQgIEZF/CBt4j8f
os7yQj4MJqWPBhN5ZvN2aVGYoO0roGD1ZwNP7MHVLbBj/SKuaeDp6srbutDMCT1f70NQMCX2Pxpt
eCLhFrGwuvKh0CBwnNT1PCQPXrPPPzgYUlrUBFI907NiGvNf5kwS6fP9rwX6SsQbRhbk7s37yJQe
qIFWrwMPGG52BWsfhUt7qljJmxdC8be1Zi2v8dUNXLo9P2nXNObYb6yuYuSnY8v+wZRvsw50CHNo
H6yNMqSsxiOpHLr1AgWD5ABCMm0cV7mKF3mgURUNZV43Na5RK3cOviWB9uuz7pNfuz1Gln58ITHt
3ofcWI+NAF+KRIiCI3CeRSfMKYnHnwinFgIn7CeHvQ+HjWrjMjCqo3nAXs+WHRD2VpNm+A5VI/YY
2B2p3Yla+Yc/1OqUBlL8PzgN3FKxrI829wCSEqLLynFrq7Kd0DsXXs7bmG+9GMc/rqvlPiCoeUGs
mC1JK3k1wpEHxkqGgCYFZ7xEM858NiByhRLqiXd3V+0PzOnlbDrn8ehjIm49WmVnjdjX0UIh0tYt
soaHFp5AOBx489lerWi9gJAQNVrtA4WFQxpW57uczzie4lBVok6rFYiC+J+fmzb/fxdkuYlq7hsX
9l+2Xho694RYprLSn2D8aIZcwPAftJThBUZNQ6keYBHMUYttCgwnz0ZsKej8qd6RuziO+h+Ur6k+
sVRy96uFTwr7thLSQjGC8rs85JgXpox3fnnmUwxh81Fw4SxjHikMM/WcM9z9rDraK1DKgW9T56fh
XFQkrz6/wJvUE4BaXQQkXnGiDJjqNI+XCIJQXqWTos01DGVU3ntolMS7LcsDOVB06Ft3fk4VdVDu
eIX5NcrO1yM8grZBiVC79I+3gYo12UcnICEQXEQOTn7niTgn/5Ihe8DZuH/Do2Io5vcKPbrKu8dC
B2GjHKS1hpeGGtcJB5qPpyJpoRhFVSPIPU9P++LgShuGxXqXiApbZ2HV0xe4A1Kjg/0rrFfLyLIj
9egdfyhCzpxdYWTAGEzClNpRL111K2SgyTwXHNO1pJmZAyEEWNme0EgcWxvgw7P8zSBb/NrvXSat
VZEyQ/SnQE2KzRSdhDJ4eeJ70Mef90rCLLm8G3OHYeJEcWKPBJT2tvHsmVQEetnFJXaWhtQK9lsp
HL6OQG9mmfozXemAlB8ecxTwilhVvJg31DyMFpiTSn8d9PEV/6Nbs+R1NuAO0HdrR2xiTxPA5YaM
r9V/Df/uUJXNa3AbYh9rex3IpVhEqork/MZ56XT024geDkR5HPS1ScfPIxMRdRYQk9f0HS+hmpQX
9wFlPYJFQA21hb2KGmJQkR68AmSxFM+PP2Pz4/yvQos8/P6Uo/V9+DZBmk6Gi4iK+H0R50/n4k55
J/kwKE2djSqHcNZ8TvmJPLeqqqnORB99Rle3bTEhAZ3Yy9S3NJIL9INSoaBG/2Nkd8IbrxLuytnS
0BLIXmKDWdMOOeqdUGDYF8NUwbc6gLBhOT38Lds1ukJmVREzY3Z1Va+PLzgh6CKuaFNPEKtQePp5
yhprIv+zfGBG3wgFNlp6PM51/UYFCyRyfRO7/UCXKsI8bCbDOALffw2KlH21lfRY/Yw0ls/c9P9r
rdyFQD8R0IBK5Gs+S5GJP+63dN64AtXKr4AFar+3ynBW2J+rBbT46qOGuhax8tgd58OQcAfjDBBP
lxtrgmXlJRE6kvATrRAbhhQ0SfjT4PpfMzyetNbqOeZqddS58tNpBQHon203xFhom+nrJJT3vgyB
M+W3Ozo22h+2D57enK5T6hGqwfv+gvAEQEEmUdD6HpfzX5soYB/SV3eu4B36rzT6SVZbuEqegQLi
hNyxcw4zVtQ+ffZvutCswA7Jb4Yv30CO2kUEk0UysgoKuEtgPEJsdS5P3GPlg8YIJjD3TM0PMmrw
VSmTvno0LliHufqA2gTVV8L5GYwcLD4AX80E7F21wEHEJTCS7gVvxvTvvIXSu8uSxIYijtmC2hry
rTHAGXvjznCMhychJiN+Q1ESnu4Ch+Pq3+EssBaK6X8hfQ45cf9PFiHEiaI5RY2V3whgDWM8MOoG
3h6q9Fom3r0hiIwMee1a0eGFaBmGvoZD1IB9Z5/27fR1ubGZ4t90Ykva1FCIQyCKmlvXzIdY4/ip
7ojME7cnQKeq1vEEYrSnGP1iFRAYfuBGZutnmNpq7flznEgOAXS6d3vb/TlwNLBCcOLr7sMnVSIa
N1UzAg+ZDZR3Iri1k940ZEserjKUSvAjAm0kJVVBXI/Qks1bYFh3tVa99rh1Ymh1w6zZtooRy4VO
jQ8X3xXHYPu9vHa4lW8P5cT9A1/fdWrkQy2t3FQtSeB+eSpc23Txj5As3GGy1mT+oj+QN240g9Ce
wFtqRWe38Z3LHCENkl2x6357tAAOfvRQ9hABqF/tt2GJ3PirEwKfITtMcj42UjaZAKBd8l566/hU
qgU1TGoduu/feBvEfqdT9muhpmSMAPNhHFkUVwyPA1uBqQn1sjCsTRABydmtZlbBoZOkcytFFL2X
m+5bGFHOOEEOPeWLoezanzF+aazfxPYfxeC0Sx5ER2nvjxeNvqkthPJLUvP4L/Z47IWejs9cmuBC
rh2GxeKPd9wjnOwaGLp5EYWdtftjwtO/Aub4GWtUZebtyKF/SuLR0T4bejOFpErMBiN1OqOb2urd
Dv6PMArDFkINOshf40Fq/CsGCMcgbyudE9wAqaTIzApsLOlGX3SY0FuHBxYPQnzKeynszT4TJKUk
Jn/RVrJmk+8pcFloe+8dsIZcl0h3A8/E+WcUSJvngWd8sRUIfv3wBD9XfMso5E5WEIno/J6CbEZ9
tRrWKDo0JuR6oHaQQIkSLFCQ7x+9A9NSBQzF5KtUBXPm2hFLrPO0ZaQ5eKjxnlrLi5gy9LGxQsm1
DfK/qcm06Ui4iRt8nZZ3Ir8q1AFo+zX+8L+ukBfMb7TkbXa0HICn4y6fdfY0rsy84qcM4scqsBr2
u6dfrNvHChb3kyzjYg1cKDkVxzV9IPmcrW6yTl2yYEL7EL9G/m3Olp200MLPy1Fz7nJbr3wSHfzL
U2Ap0CqBBP/9vWkAMHUiaHHcJ/WA7ca98Hodb2OGyez6emQAVvkdqXk8JBced5Oen9OusXXHxXvz
zxhzNLOorcciKMpeqJOIgid1HBDz85YQx61WWGQ86bNgBS1r9xkJG7DTt4u8fPuAmgCqcOFNCCLu
T1QfQuPnurYenkBHO6o/yWXBerIj7YqgLWrI81smIDhPEqUACtrktab8HQww7UubPUZFne5w5kTD
yxmUoKXF+A1O0VO2/qKKSUITZF0WAGwo0irU1aXYEFinyVLD00I1+vXWzT2rKh+3xAQAT0vFWaV1
A+UV4DEMDytsC1Gi13Mvme2FXL0L/2ZUBjTBN96AATUEvOrmRbBxblAXiMYTnH4OAP6EGCCckNPf
QaZIsTvHKeqCOL9dso8jzYJtsIEzAmK80xrff1fVEMMjrg0hVuYaqzC3wTPJqc1qdNh8ggpaoV5J
xCLe0ShhKpYr93fRfnySyQlB+Qa/Fc/25EyT2L0aL76cUVMJd/oMcMQA4gN9U+LYNZ/hgczA6Ib3
klVKS1RaCpl74ghIncOfocRKTDfG4+Q+0gLYQHn6syuqSz62iyd+epwoEahtjjuURfYTldPAILCI
P/WVCprZtKmF7m7vGnWJNYLBHp/IYDFGNbtT4EYuguQskU1QtO3+83MlbCWoP9hMSWaNGu/IsFEJ
dXMdty85CgMCG6MPk76fFcGZ422aHeMbna4HZzNqkOX9nztw1Zc5taLcEg7J0ZAdgr4GftL8BlqI
0L9hL0DlhbK0gUpCn5x+ULPwH7xoIBWLTfjG5EJAI/suUAuqQDb76Xg96yALs7P++L1BgBDPVQiR
+MPCKGxMOXsDk7lDEfYcEh46ryMe2N3HSe6Fs/4YJt4iD/xnz+bqAIu5sYMNsXl0nEsJ9Uj4OVfb
TAIhVIuKBZKDXjwSvHQ0h8sSg3tltiqhreqnbWWNCIOT3v6BdAmOKvE34SBBx2t7QdEYeyhW1XAm
Tl5ZrNKbKkc+9iqQujD+T4p9HAQgpr8I+sv2VLQojmUcsN/AXTewHeS9Qkltd1M6bpa1r+k2uunN
/X78/uzoNwnLBp+phKxc0Bb1/W7FJ5meDmCv1NTDUH7lGY4WHvbcvO0b7xlK7keezpCMAo+zFYzD
3Dol6bhfImatw/5j/AuwcRHqUBBsO3xSwDw6Yq1GBDTX4cb1HnHS4iYJQfRD3kdqGrKPNZq+0hxk
ltOqs0174YB5RWpE2ydUSdujBTp6dEJgT2LnAQScUV65HHdHEghuInyrQ52vg/qz+IPa1ZU27FNz
+I3av95mfraTzw53KGmHtsFEQ346W0yYVG4Fs19iA5QzXiIdab0YR3nDPtZvZvUA2NBYTQDp4guW
16EmYwWS593P5iNkW3/f/IDna2Ky9pa95KksF+/VvbrFjVMoAg0C/MOoduNCSS9rcgB1lSwFIVTF
g+ZxM395ZSaNkKr87q8ql8SayipyOhDg9poiI9mrUsaZiEqdouwaAZbEyVEJKsPJ8v5uIoyUo29L
d8lPKRsH1Ic1FauI+zmmLoUB2G1KLmxnLIeVLg+2HsXBrbqPChUK4l3bm/+g0vQqHVxx7C/2fViZ
ax7W1yp+10K75XxyPbRDaCJd/u1twfLDdVGRlXbjLRGni0Aq4l5/GpfIyfbT086JXvgQHL+EeOgy
BWMr5TRtJHosG1lJ5DeqIoQ2Be9584h/r7aRabA5wJAAbbesPDXCWvCwBXgVKQ9AJy9wmPQcsIbJ
Iprk/BYKKccqwCRccesrA/UyvXZq934rppjsLo8wNjtvDMdP0Z3/dcNX9QgGlX2i8kS8T8gfEi/R
C1QYSyNz5K8ClBATCqSQHMt+ET0kIGOalxy4tGOLRREh4CSai+rxyQYTGY1HqUoGkGXtF3gi1BqV
miy5Wuo8g3gwApkI/zEV1cYYlJr/81cixlNJECmx/1ozezIMMuwbxtPhow/jU6ydJHweggdpVj27
elpa0yWF5Fgp3ozZFGMDxga7IJbCO5hnb2v4kbVM3r8ofXngEHSN6FG+QAY0N2Pc2hT4iYNGrFtz
wSJGhs88K/Wn/yGYZqy9aPglnmu8aihKM/SeB5dDPzCWhQDRKui4397q9bo7rmFICU1zTVt9dGgF
U3coBVbbg+Pj1IgdboCTr0rLnsXeugM1mG9MxJSxMNBQOL+g/8k3/1lBzp1g38wcJlQztbnlfP/d
kGQjR9TwcqpujSbftDJh7o9KCaAV0lc4z496vCKdh7RH1DzEH2mQ51hoOxo1HCtI+EKNy5KFWyNv
7Sl8cbdI1MHlVbO/xgHFci/mvT+ENqkBPDlncWMUmtCwFvO1wXzNsYrTFw3icNyFJisPjkbbmHsh
8XwEG3fRhJf851+tCD4/EM9vEDhZWcDmrPY9zY/Xvhs0TlF6Uy16swqWQoV9PDUMEEXrjzROg4yc
/BW0mkM3Dvm5UMhXlgmM80DQK7v8hrY4IDs5uoPE+sZcUy5WBdHZHgACZPNzhMZ78WviSXBmkvby
QpwzjW5QfI9PXvbP2iR4DIAU0NztXPBWMq2iMyvfWe/kTs75Fr+UHGwBG4CmC6pJgBUDwsSAaeDa
2SXnyPXW8l9YBZwSG8LKQCHUo8egrRTcat+BjoW4TWjWVxhtMAtIYJHym+lx5X2+m4aLkZ/PcU9s
4+Nf4zprdb8m/cAvwixe+nkfNWxVCO8VVtu7ko5YjMA3ga7qLUBayJm4gvUVBY4lkRnpIRnlOXd6
hLkhBWEY4DOyWnFT1O5i37ZDNoTxnEizxpRrWYq6NYSWZ88xXqh3mdMQ6TC26INv66M9pvW2qCCV
MiwQmO7Y2dXKxgZ9Eo2GzJ7Wl3C6Ioov/pzgYgWT8nMvXIGLDlmevGnpfowHt1BoQTf/KGvx0Hxs
lSLRNx39WuUeabGEvo+SjWexbp/NjwSWBSDMg6/ACzUGKFw+Zs7byjj2kHflwipTUySRF79o2X8K
0Gfr9sG/zMf4QsyKWqh3nkyRf+QC3Z/SqtuhrziB8Jd2N2lbfmwYGhGOumqwqKsmo45KpATXRfle
pF5QWEo0U9SYsplLc8IDFRAWxenqO5dL6+CSGEyiq+VKtY26Vb/AFpZ1JUCXfkMPhyT2/U07N71X
IqCGl6BR1HTUl61wZo1Xtn7AH8dDC8Pp/gkuCIf+qoK7nEkomgG7JZjNvW8Z8GEZmGYra4d3iag1
x2X7DQ3VYEBHaYX+T/nI47K1cTlPUWHuFa40gqa4ynDa5JV2kBpHGpK+HU7qCmxvLFqQcgOYEonK
2aYpKWJotZiBDWqPa+gF8vH2KyZ/agaXsK+QAK5wHsj1m1oc4dFkEPJ0w12fBCaeTJQvylm6HFiH
6N9fWfvvGivzT7NfPteCLx9LZH8bvR69MkEP2HWQ938O154yodlPNWcraApQRiyALkTvEt29nr7D
V+nD0FLAPtskNguTzZLO0r82MkUWFrPqYeFV+/HoqiPNOqWftIG24wltmI6YDc7rZ9UDwjtaoM6X
N3/tJ7oZa99U4Y+k0+tU3Z/hXTI+nafQj5+p8yXCIQCL5Zl0DGhINpbcUPOIY0cowGuXKjggkCbj
lGgX75q+A2JkdxcU9xPiGNOzFRAhjHzCUrA9upi3ELGSc5bZjTZ86by7sGK/QXEE6Fd5JJHo+8MC
iA3J82agHPLNwa/fn9uRwUWDJXdGOug5qmGOAMTRmAG1azNau0ch0nuRYWCrOqhJUujOrGBb+j+2
085SsqnV9VmWkka4IZSLOTsMaOxmBuVOyVvpqS4P6/MLm2y95EvODbhLa0daJva+cRRfa9tFHyHv
ofoywsSUbOYUEMBjSAQhykJcpcMR9S4qfATckRiUN6S6vlewfFY7RiPAX78jVPDT2p1OSOAbyvkb
tGcQX3H9HjX21HlFaUk9N+stW7HzqlskPhrgZj9pJ3vmJuoPULkysIr4DZ2fDDcybg6N4bM9suru
ppiSx/onArhXzEYY79o+a8AM1/K7QlmOODEhJcX0pRYhCFPHDWpX5ps85xUh82Jz65mjVV43fKUj
reWDksBRFTPwA1BHzOhJiEbc61QVT8jyTrjGevRnAJGXqNaAQJOQvNo5ECAApOzrq9fBeytmE5c4
Lw+ex/Cwq6gFOMObf0NvpvMu/S+rOnBeIdUhFJfOLTir4axdzpyeR4YiqpbrfcBooO/T9yvOvD+y
dUR575XygF1X3raBTGq5UCA+7A8SKvT6JAx4dJkHGSYBsUZeQO/AVQbzPuRKiFGlChlZteo5Pa3t
6QWUk4XS8uoMSYFLWpOdQD+1rOCj3pbujLaVtJ6UgZc8+K1jvnum0B9jx0R+WgvSYDlGKBmVAhGi
PCgOo9xD1e6LT6ArtWxfDQmI3HnsVXkdVGSFtwdvGYQaoYm/o6uJTWnsjmhdrPitrsQTjuITHPSi
9z3T8Ds+ihECpvoFztheCTAzjU/Tgt7DBCnLObp05oeSkVg00L1q+MLrnTonT5RE45EZyqe/oQIA
JaYCUkcOaF9GHLFZ2XwUVAmsgeJfZOF/nh4YaWiJCmJsrW0a8K+SubZ8p4EPGxH5NynmHS71nOSa
7l1DWUMnYjbjVMM0WrUnSV5o5G8P2QlVq3Ihdz4cWXGWtppqA5b53aEYH5j3fwrVj6QsALrIdnkH
KPXjquwtb/UbZIOAu7Rrt5KkCa2UJsyB/nZRJTa8GlFU45REngslP7JiWgzIPBuGNP7Q+q6iFFz6
kL+zSkc8bEFrosOUWKTrm7JFl6DngBvmxCR4P6u4yesBjFwBdC1qnKFggrUwegQMMCuJUoxIh1m8
3FiWJ2CDqXZV4zcO+M9ck1LQnyl2r3lPy0XL9sIHjN6kzu8UOxw7F5ZZXkdNOIuBkPbVn172lC/+
Oyum2JjJUZe+8ewKJAjj7q9DodG+Ll0l7uWZEuNPLeepJKKXy4hfp3mo67Nka4kUwGOogDZ0NyVA
KD9+z6zqbfQeUi7gdQwQLRRvCN8ge9QEXU4S8vt0ntz/JqIOQqWchaoeKKJF+VlsQB+/0YHScBO2
FYftxaxz9If0IM0TMsGcBZZ8uiUx5/aV65bqRBVI9sZzRiYnXFN9hSwtHsy77/+z7YBvCc69PO7G
5UF7t4ZHtLsrk/YjfxRCKQOOcUDS25jS7C9Ej7eeP/57nzuelZMRFjDI363FW0VVOtoDn9q67Yq1
wXZIXUfh89nxF2tPybndygVBwDrnvRbrp28RsAv1Uy7jgWEnz6w52pxPDcT3FEY/Gwh1bIO4n0Kh
INdFyyPoDssk9WPNekOmdY1lKbkAsgwD6aWprhF3Z4YvwaxMCpf0KBHl4Ur/pBKcxWAYM3WJWjp0
KRMX7YdW6+QcgBYAsYvhghwamKrcIpuoqGHp8ljGxUWOyaIlMdnGbGdfd4ZVut0PLc1LQx3af4Zn
nX1ywqZNbwhX70xk/pT9JJ2ZqMUxnuKNyVCo2w1hIVpJZNK+9j79FXPmEscmQgmIrm/P8MnOlkPa
VA495YaYfHJzLwwKdfCVfiSg51aKInvetceVayMqHBCOJAD34dFaWHxas6MzudB/InGR8/QDizao
MEfcRqCPrdQfF77boJwPEOYi3eGfF05/l03o2QAhu+JV1H+4slDWn/HgoHyApbowvbO4zu8aqsxg
P2sX3Ui54AXBksbyc0EpHARb9MqQgr3/MGi54YAJG1RLz6Ezx08or5Lh2iKm+Cj10g1bqeYnpcY9
phEzdQWLZQCI1RWJcybbWMwwyW4VJveLnTKiAvGAjVG4XRYxCWWbi74IeaB87LqNoJ8QI4uUsltJ
Ys1Gmqt+X5pjxlbwaRV0xVcjT9pwwy8W2uMGRbgiE2RRgxTTg9sZ6Bo7vQB3/MrEjCsSLuojDWDU
LQUBqHwnEiClKpu3p+cUKkNaoJWN1om/aX3hD+irGpMx74aB3OsFrxbY8Ui5J8vkO7TJhg33hIBX
lyTppCLs6i7R/1PWLw4XlO9vAQFxqsjYvBetHFyv6afieUJX9kzWjcGpYkohY4Y80mtt4jtsufwB
VFiGYVuoCFhHxB08dx9zM/g85MNjbJMEdvG3e0R9mQbRYVSLoUIAgZr+BL0YROJLI59YmfrsWLJh
6ouilT38DYpVAD5580344s7lYxc2ZlXs06ne53/EVAQGtqb73XP8oQH24YVlk74YXi+Yx97Tj9aT
7OQFgsBPEv9c5Xr18Z59Yl/XlWE7GSb5SDJRYxAdJXZV8gd/nqWb32LlVlcNP4l3L1MUCfVcyUKk
igvHhY+sVDRQPrhzoUlP78eDH/FhrENu8BwPFpVjiYV+OnoMNTU5Yv/oNwA+f0RrP1RkSIabpa/X
vZJqohrAuD/sR0nRjJjjQyORP9BYynvsiGykHK2iGYOHaHL0z3+J0xaC2igAgJSKhthgaMBseOCK
lkhmPWMZ0e8D0QkeIGtQHCNDfbqxPQW5Ru9v1CccxUa2bvYKU2MOTxMBZylr/EdBOVgNnkQZwE37
PDykO6UdpPrkpLXWPi2JsjXWbXUHa1dcBbBdkCarWYi94C5aRNEDRLO/jSCzUG2r9jMkE8DBK3d7
9vra/Gex2EpKZK+pD/1Xfg4d2ado1MzP3EAuCBUjcxo8Z2S5Ox8SzCrqwvvuKHZzVQJuvXEaSbZO
h+JNoFZ3oZT3Uu0ERCgGXGT30Gt2pGXJAASgHxmykm0hYDe0m0vsWLkfDkdogyR0wWtRV9mWYAAp
rwBY9JRCMT73vkA4FzAkWVXwwLYaA8gr+tu3e0nSBkt/iqv1e9HTjtrov40FgFRkGGVQX6p6sas1
TFOrwBfZnsSXMWzl66qC15fkqJtQ8h1KDQeH+XyOBUNat+ftzLj3yih+/02lrkNyljHGRqQP67m4
JwmBjoQIUHPE6IT5rkaGPCk8iS1p4+ajkiFr4VhcNhfwZW/Kmqam70WHl3Nv8eTH+MPX/r+VoZ8e
x9bCb1eq8iOUUAt38yfhT1jbUCuXGbHA5rJS09wLlH+KTzY6mSwJ+DltuKAx9uBokALCw6xBlq/p
QXBBUNDqWRh+PL6Oqi7mRoN4XEGLUZhMCnBCIOTpQp+UvbJ/pNu+u/Y08SGks6SCCzBn0B9gUgHj
x5T1UM3s8Bg4caXXSPo+Cgge/EC1Nd+caTNv6l7xwXpowHUpc9rBcbeD71xoLemztYNRZJUeBWGr
24VBI8AnAD4vM1LHeq5vx82DYud8/cLV1Q53YajEfNC4H06m6G6ZtUIY1zN0CX3STw8pWP+pBAZy
lFsIAaCu9KO4CL7YAh4jptsjgByCTMmKaQAMYAu5urAn11L0ofhdku416R9kZuN9m/Ai+VrYDuWB
eK2JTH1WN+2i7ipP9nukmW1ilKu7gn/HDiRX1xVF/7ZBONWfd4V5vfkxL7ZX62hGAFLI/vuQ1HBi
O6qiCGbqm34H6asJoERbVYoNWbfX7zqeqz9g2jlpG9d8jN5nf7S1ug7xkIE6N6o3CTRPbRqFtxsL
zLRGuiAmChBdH8rUSVoHEuLkAI94q39IBqvNabwirU88hediz4Klxh/G6Z5Kkhy14hjPKnToj/bI
VoHnp1xjQ1rhiknalSH0vBjzAKEbv8+pY+MZzZy7mRMQHmFhmW+NXL3hhqWC7NylQdQz5/AhXIQa
6Qi0zEpCNyUj/6/ypqcB8vIoWKggaXbV1PJLwexgPeSrRN0TkcqO7UHqqC22oGm1yYu32a2dDbea
GaCSVY6uRO3zguVklS0ItHY9H1zGf0GWqzrUU/KjVtitr82Ze11i5YCrtq4q9s6jvPpaqGXWPyy5
Z0hsJGOuuppWmAVuCB/ISMBX1yafZT5UGXn58/Kye+GuHSCB/Q18zPK1Obj9yITF25xlJ3hzquEJ
EKohkvPpHtLh1p7A7tcrnop2eEAB0gB4rcK8KZ4NmrRhxkqEEmf0pXOaBtEy6iqzkxSZcxLGM/sA
VWGF8dFvnzo62T4ThChEiuZgemDhyoTJAURuIa8n0TgzkzHqJJyQ2Ii3KR8AMece0/DCjh3jtxOf
RXhwPx2laIAuI6X1BJM2+9MUNMs9CILrVpzurYiiwQRItkW/Z9ELC6GrUVrGCnn51a+Wuv7JIuRk
EL3DlpHGcNJpuQzxe45qHPgXM2Z7Z01JWkJmU9OHIPQcDYAnD+ReR/g49vQxRQ+i6aE5na8GwP8r
6yZD55vUhNYBDlxY2MXqSANZSoHwt7PIeB6m9X8oXKLNzmxx/s3f9YyF95kJD1gyag+WaYECrWzb
Spz9gOpye0VFrjre1L0DjQyt7JnKndHOYr0IqKaFALQCbfFJWtK5TCtLbnZ8pvF/MdPZmnDxp80a
2p9PATYFVMFKP2SSr7wVbNMGmBG5+oOQjYNo9au7z/tN4VTTElrwFe/giyrroFHqULlLwBl52qH5
a+jWBRLlWXTrqAn1ChsriT2GCCKpyFmu1EvNWKAc5wL5tLhh+g69+zJ7HtgMFSB/FAYewev6LOKT
kTKEv9Pe/W/wjJgJb5FNeGc8cKiYJfAFG2lDEb1aCu1WC0HAAJnch7aVyvrRZDUg6giaXSBgatAk
YkaLDigHxDfsqneZXgMT+7n9CRTRePyODLyjKrqxh7vQFlEZySi2PagI9ErSMxMjVs7YiChi/Y1W
g88eRZ8Hpz4JueUI1AWWqGWHWHlYpw8dxNsB7vYUHsH7qAIXeDA2KOtWEetZGGdGJC+qu2ibUQ/m
fGSZpI0rJMhQTeN77wlldl6aICj3Y6szHEL1Uhp/MnA4PpREKxj+xQDy9N7+uNDpedGkBr5xQA/K
tC2rPDpYIf9bDtOf12w4NjZZV3BbfDETntemUS8baw+ezppuMliwY56bdhYPzNIDcdZgMrSiY0VG
AzK0PrQX42KH8sQmm+VpDfB8oB8Pnlyz3qrGt8ec8cpiieKiGKb3Aa8mpw4EzkxVtgDevNirGwQJ
uoqMxUhAOVYkI8O72lugaU5c98AaVReUTsB30ews/JOccw2q/bRUeJTgKSoVrm61KZFwrIpMcHLN
0PlI1AqPYO81w9JcDKJ3u7OLCKmmzffVrKtsngxotiegZ05o5p3rijQFGUamRCyDsMfpKRK7pT3o
gLE4jcuGoCTBd6pPRn9nqpWeh0rfZxRsbI9kipaXLm3VmbEXVtr0yVItI3x5ynoUM+24wYlzprGX
M2U2AbzkUn+U7KdxC1aaNpD9CfE2La/GCG47beCFjLnll/LvzHMMT1o/qMT9m795BG12/a66/5jU
4J1vAOS+ScNCgzphXPmdXt8FqLIBl+Qe/U6kqkPtroZuTgTPmRPLHB5Cl1LNItSauS3TEuGf8qWY
nLUbPbQy7TtXiJi7BO2u+wiKP3+6YftCguZpah5JgGkiw2NztuUrcWnuvlSRRpm38tETDXS8OCeg
xprW/SORRkktjy1tW8q54lNbZnjpv8WoDGH9OkE0kbWHEIlPTdPqfcYS9ShXzVbZMle4A5BzdvWN
y97ru6yQHONpj5i7tU9RnMQ1tXY5SIOQzfQ/Gk5tRbF+SAjXQuYaz8oBlelnZ/VEgDuFAKipChFJ
eyr8yPsGNDH1qiWax5OJ8C0VDJkuuniYB3pKeYL0Lk3OSLWsegPrxdyhu7ldmpMCK938tKqicFbT
QV+tlaDm1sMZ/eOKOkfvxXgjwIiqQJhCrXipBNI9BnPlRDUtGDdE/7gprg0b8HZ1ehajlepVbIwt
xAQJXQmUVvYEqkmcCjvI4B0zzgtkkE5YHptEPcW0QynSZZWDEvah/c/g+4QQxKE+/UdEtDLeaxkB
r80y5aaxXIydDp4MO2Bk6bqCtXgq7gy4vsE1XrYHRV1ewjywRY1lylADkqE/4e9qM1CPvG0c4eJM
zqACyoSxO1qlwdbojtRD5ozPS/VY9iaT/49RdPRZDIK3AMssUIYjSG41R7aVQxlZnwrMTec+0wY1
pUOascyPkdiE/qm5zVg7kXYHkPCGWZlOx1X74VVvMSbyAIZVsn+GPl13WsrqFMH8o56pWVvACwYJ
IpjagIcgompcnyGCvdQK+Qeyvf7qnzC5qXE44bjSqtIVVUEe7von8AFpIeQjQLmfgiFRavzg3vkb
X5HJ7zh/nBeKxJJVvcwGCeJWU5fnO1A1MvsTN22F96tSU2pDyVlrUvqmZVqqobl4rnfl88xAjrtz
POfNogO+LX42jPprB8z9dAx3Xua1hvYc0xGFO7qqSUl2jbITcbrpQw0FW4eMLDnoWy1pxGdUApSL
JPSSXqF7kI8zUd65Dt+vtAn9BKaMpw882U3WnTZpYOaJi84LpuIGpzdguSPggs5DpS9kRA/yCGI0
DsYexmgGj+03/CIsRTdk6kBo7P5lhZdYGYzt/SqS72qWXlDOGRKSh8A/SFeLxemya8vANO/FOvyV
nSmEIhgDRuMC3YJ34ghqY+jm1nUM39Z2KXft+aApH0/5EGdC1T21//P052jk5s7ruqgFU1x06NuL
3lN8bwvnprLv0MBHab2ufwlu1AlNQUC0+JO03U5i7af7sPCS4iefyMYQuhaqJqdQLN75GG9Zax7z
BDUFqt+G+wgUkA1eRTcQzXWWt3pnZ6O6bqfyt1nC2tMikQZfNliA8hmeL2GIP4VIJBesKacQEORi
rm6A5+i0pxscYl1aYjlKCKZEzA8wpZRWSuUNtpTWw3nZExkYVfmigcB7aj7qeaLC2xI8clIzvyRO
6//pQlHnGp/uN8T5TbKwcSvJXgmnbDmkB14a/oKh5fNDOY/ggRTQYhBPr/RjPv4B++cH1O5ndpwj
PNDo5wyZVFOn2yKFsXG8jnGjIhZmtzSncMqXcisqBpGKlq+wfFcz4PU3riY7PDIyq6K4CpXyxDZ9
mjDbAHpKpnW6DgdP7uYRJNkE4DEI1SeN8FKUtZpFdEqhewIDN1/coEgEXyv//3KE5fleL77QXRSh
ps9sol3oA7VAkTk4cCYP+IVnZZLXTqzBDg3oEovpoqSgf5FGfjHa1+g2lVhmzHVF0R9YwETBrO9T
TcCj9FF0/kBjr12taaOSWTO1Z+18cqtWTg7Fzq8qbqZlTCk27vSpRmER8NcpyP8oiKRXpiIXznfV
ZYQslNx4R/68gJFWhHVVTFy/g87aDh//BiBKcx96AcbrirC3qmw7EOeV/ZicbFbDs+hwEwM7DP6c
BDXkc5twJSGd/aSNrW1EwHw2mXCExfFuOxf2ZrMX9YjurPJPgHn0zeZ9Pm0qB85iG3CdUTG4L/iU
S9v5AS7RBEHbgpqmEZwfbREMzuQT6j6Lql9XgwmwtwK8MUnhuS+MT+qPQZj+tKlWHA4HP5Kk7nL6
5YqjAZX+F6r4u048U6a4IUhJAcwbZluHW/V3Xgx2V7CimBKHoMaIBxaWwLT/sONIjsncS6REMu/F
cGNEVL1JpdQ+xSxWYl5DQVGICpXNndA4DJOMdVOnT5WAQAT16evswynR7L2dSNZGESlYM4O3Js3c
xeFkQiajicAShVX33rPYD/Csk7A+u+0MPgo9zKIDh+QMx81YmW/oDqemNHMCnsRp7qFNxwaXODDJ
P7sU9uWUGAwRHLxiPzEW/4cwuG0kmpHuX/zg1Zn+WcaAVLSv1XCsY86gzJZkjWTFG+f5vmwkdzYz
OtBK217nTwEmSzw77V5UnhxcPcBRJfY1FWNryw3VuII44IRoOwjHhao8wrswGoqi9LHK1wo0RLdO
y9H3goUNWw3B23TQAp0l5zEZiYX+AODxX+GSAmdH/8jty/I9/3nx3qOJTDZ9rykIFnf30MSr1eiA
Q4s/KkIHgOo61oAv3I6ycMHqzZlWZ0QLyv0gfWn6Ze+OwfSM+6V3gl3bdXOPb2s3gQ07Nrq5sJws
sG8wR3lkbNOBAb4VfaKuPGomj/mKKvvRlJHbnIU0tf3yCvtuPe1RF+HrQI5zzTW4EZvsnle4K6aX
Q2Y+RhLuorORoCmPskTco/PW3GKkbubuA57qgF99PNdwBnJTp5uc5+6cW6D8Ysf4+cX+5zqMhE6+
05oymoB+sScrmCNQF2c7OlvHx/Gnn0jYu3LQvIc2Y8AfUW2ayy6ppwD/i8NN2nseP0O1lHF/yH4z
2J3sn1PlDmhDhZhhrqKvg/1aA/XyZK9OG+b+lxcwH0Fo8BYI0n4rK80EMbh/8Mlg2/Cuu/Xhb96/
yMbMK4ctv/SfpRd76WYZhyR3DgeRX1aFccTQNONZCgXJflBip/qlODy6MXZnajjHnmZVxnZfI4xo
qqao9JD4776n17dtE6f30nzv74WQdgk/d+iVl+cH4RV8iom44u93pxje9+i76vBIwqUFVXXbOuEJ
Z7zfYFrrbMnYyI32VJjMuXW1kLA2LttnMLer53/oL9Iv38TajkZsJT3yjSyXSRQhvsrdah9P75YG
vYNXgLvQ19ecnDwwvGO1BxHwE8GbZzxAgAcPcbkiXMAHuM3bTcYncswhfK3dEMHYrHJJ4bbFSqww
qEYu7sSGjgzAIQvwEnz1IBTOh5HdFYia/5O8SNrSurnFQVs24Y74d5ZFcHLaDbWlXvPYQYecrVeG
EE3ZrkrkW9QhAtHohaHTpOgLwuUixeOT9/JYc8spO+fwtw5EXNvQQHsMNCMTpYWsCYWXj9K47I+l
Lc2209yYSUu9TYyFqmAnl7Z6KlGt/wDzWew0FqZQwNvcjPlxA05U0q0gGxlm3cNKPOZr1TnxD6np
M/p8hisumarH+MZC77PXI4ZEbZ200ISOGdInIz9Gbgs0gwreA3JTdBy5AmhGo3rpY877OYEvS7wq
CJEO5KVA6RToikX0/e7YWfjTIkzc3ZVzrBnhAuq813GBklnhET8YVBFYEhARCjaIpxWFGzKMfhnQ
jul2AcvRbCoxd+ogWNXXSSdWPi1VMVSLGGqOOxNVdYSbDw96CWflbjGMHzpJKvELp6vZLvndFRKW
7mHGR5AiWJzEp9xQm9dMnWIvEG9sABADavNR7v7qS8KUZglDMcBgtixAPesePB7PjCsb07auXinm
adhDrDJKahfe9v0PgIXngiasry5B+gYrb6C9BHPJl9qH6ghZGTUBxpq4Z3tgNEfjlBMW0rL+q/vO
UFS6f7OyExYL38VmM9302Ef2lZNMotkmNA19Yjof0cCWbDPvw0xWSr990RyZqSzAgx+DL3oyiJO/
zh+rggBSS7xhInTRC48No3h9TrZJ+jmsETFYoUtnJ84pf66fCUhYJ29Kbo7vlYLsaB3lfquBL2aP
Opklw4hBs6SvSL3BtXfkGayfQqIFY38W83ApB2jFQrnIf/EjMc9O9UIexThMjQYR2YnxzKpLjyEI
ytZMOv3ge+o33FqWGOffCkS6Nluc2bD4NMQNAZP09eMug9fy/0VSvN42lEdClEoz57x6UL+TgUWt
tUK6p8Gi4w/Fe1klLX/FSN6zZIxcqXrJVTtOqYO7cwUYscWDnpRpyC60HxCw+tb1MDZKbP/djgMF
KNgB0t1D3MfqEnWI4y97usw4uX9BuWC9ldT9L+QvV7HVHU0DLqGY1Akj1nbYWUEEIBR7USad3CB3
XOAHN0gW7MRqe53twWBO43qWVzZRaGiQfCwis1mLYUEwGZiS6poRl0nmnRznGkc8x0gRtMr7UuEB
L9fLJEFabR64I7vDUKljFh5Bm/yyGVkpSdUNvy7o8sjdUr4d4ymc/68w6f+DoanFTZAw1xd0yETl
eN3nETHsIoXvjsi6UpM0YkCQYRhY0o14V07f/m3lwbPfGwYEMCGFtv8hiEiBvDpOX/O6e4hvWWDR
guATutcpy2+yp05+R0DSWHvZypM7Z9KyezLJoMD06CEuFy9fKUwsf/2Jbc4UrDo8ccNTtHrTwCNU
Yzs7ihbr/1coZDHf9cEyzjfxoZ2GTVoFl+5VtFFNtH4jAqECyCjRkOmMtBniyYFRjukOLO8+te6Y
qqe3DKWu0qyS8jNIKaDDIyrEQPnPlfQkJ6A0B9LTI+7qmxEr0iE6OBfM6E8VVKnh/HASM5KiLJqZ
/wjBsjskvQqFgHZAcIFjbCk7XZNGpi/iEm+IlHZmm3XpinFVmHU3w58GOmbq+NNc7MppWSvb2Psx
Wj2zIEfZuilv0G3ccwh1cWwqWdqkkv3TTkBjJ2vm5N1N9mV/Bpp8R1Jnl51MMVcaNWy4m4cakIEh
+qLl/IU/vhV1FtWel+V5DNRvMFt/z21/n4cDP+wFVWszvZFOyZm4H1JKv4WVQRJUDgIXa/XdCelW
r8tnIP5OKWnAC1E9Q8I3LGsoy2TpWli6vewufTsAtrX5dOE5IeIZcb8GWed3D2ePnes1ddrrEd6L
j5x3wdxP9Y9hq70MlwQgC/p1qtbF1KMlnfX2sCd6C86ON3KiFNfFWHAISWJVscTJHtTTGoiQ6l97
aJfgSpR/Dkd2uvCHbt92jI1D7NY4M0uprGZw6PYWTKh+4hYi2SAG8Hn4aCx2nfGPV8Mid0e0Bgw6
m4xnlyWJTr7+OosKQ3IJAz0z+D9yZvA0cDNPuBDtsQG44JIZjr+TgM+DzsMEyZsD+RdXdWkRN+tN
6X+/u4KxWgPS1z4LUiCDhAcpMyUNyBkaLnmc4yRwFS8rdPeh07dyV/MxcEt9OnvuV9Jbsbrdsdqj
0WLe+p+EUWUZ7d9u63r+WD3Mcwi2ec84f3mpVSCjLQxquXY5BxQECl4hN0B8vCrgG8ScKO2rg+4/
upPeoMNO9irh0H4yEyfojt6Xj5NSXffUb5KKEPkDzMsjWaBPqvz1n3rCWa+wiCT7kOe156Utc3jD
622l7F29Fy45TFrSCoaD+revQyjQKvz6ETr+vf3+5Yw/Rr5Hnq8gNTLKP9XnhWunAjr+j4owI9IJ
/8Rwi7uHpHAhjpFxjgpvJNXxKNaRuH0ok3RCWJN0URfPMnzGPqYH2EVf5YUWVzSC4LkJObJ1B5cN
Gfr9/eLE4JNtMcEU+Had1Pk5HObRh2OzSEjLeVjYGreU9sOXI6D09DNj9kypk0rrIOB2VG9+TKug
vkISgOSJMX1uS4zCRCYkI6B+RJkcBL2IQ41IrLstbVhWC4yh6AQs5XfdatpNXB9b/b+3TXFkZJhc
XgYqfup8og1oPiQk/pEishRKwwxA7CCjEt10zyE+/eC9Mrs044WG4bO8ydQ8JopyD8cQc3kOD2uy
6EWKy3oc9cUtVedgpKr7j/gvKOKYAB4Bdr4pjoTXvqssAZPCJ0WsS01GZEzzEhUyiOlGLFy/AD1C
DDwRJihhfI2iLZCs4KnQshL2arPqPV6RJvDJ1F5wycbWwXxhggiyLVGpinzEdYRNrcMJkhBavAqN
jUS6YvbgfRS9o5vRVz5svI1ft33Q/bM9dvhkYRreWVowkfvF2KIGS+YevatfDdbkTURVoZj+BS1r
bYSen1PHBWhEgNrd5Uxgb1KClwo1YhhxC408LifVXpxLr5YvW6I4MYB+suGUzZQOenpFuJ2lwBn7
5fNBKnoHui3S3jujJLNCclOw+63fxeBUA6PTq1STqu3yTErKk0bxMoe1/K2KkGDyftC+vl0QZm5H
uPykC5oJxfQTrEk8K8qTNTm66/5dQj7Ye9+CyXgd3IxKyarC9M1RyaT5EiYjy7mdQHUQ5N1bC1F4
6HPUZY4TjG0ZlYI13519pnzo8r6i25XPBFvUnYK9mczGAvh01BMzzLeerj1KSzmut+5K5yczVw60
MfASXcEI6GHrD5LwHuykpM6/2ofMMDucirXcEPB4VYcrNQfWVXkG27d2A6hg1JWArYN+/QPPxov+
WxDrRgX/6rMrvFPpZSuFj48tdu/xlmGlGyF8THZTaewpCkbGhcNZX2t7LbBdjczB44o80cmoU9UD
TlxiXmIfVn6anbhoKxmyY55obvPgQiHbzVZEkAGp6c+rfC34tfALpK3q45gJZAuk9LZr6mCmcjI5
/F8ZdF4qgS4aeYaY+s6xbJr/7mV1t71KQIeKeIXmbxclk8f0w4e+/QLwQOjfpZvgFLu6TFmzO+Tt
E9nX6vVbgorucBCWjL87hkcLOjg0VpYCfTsxG7LLKnsEAj0++LsVWFCedQq7QHJXj7XNVIiFa4zL
7/YE5AjnV7DwiwaaAk/1ROpmv1M9OVHIXN/j5nO5tZp5wrx7I24EtVRD9dnG78wr8bRpYx6UAxyP
zW5/I2UjI8sU/8SlpVo8GsgA9c7CAf9KGEdYuGuonjsejVsVwoybLFmgJf4xPmiJ9y89mQCJuGWd
ztgtFNFwP1Lu9ItshY53FI43m81/+de6AYpj724MfSjyjqbjpbOkQ/IIiUY0jUvzLeMoiDYBZNDU
arl7rJMO+W/M41FWJSvkuhNg0KLNtoE0N7/mQRY8jxlZRPfpw2TQStX/+IWCuyj0r2GVnwAoZzzD
N5EPWTr7x1qsHQdtN+iHR7ITpUOSuNPnCXd3i9L3/4/YrXSsGzlH78q8ddr+niWEpixI8nnJjUbO
dX9SE88o0//pTpva9xzFbB1JOwbMUjC9+xGTUk9xeSwCcYtiYEs2nImX7o4bg7ZmJqnRcDU55RK4
fciW9KSEt2fEHg36/hkxxDlF+NiGNcthsfNNKrXh+MvqiYvQEVm4+ifMdB4W71eX/a8D1uV7YmVr
+Pt6FeBIFE+wBGpZR+plPayZwiYUnuDGY/aBHiPi/iSyYHpZTEN1XIOETyzUNEWUAjOCz5dQ5R38
LGctCbcWBdZ+kIjvREsvakbaJrp9zC6gefqc4mUDgm+96Qkh6R0kHahuwEXDAS6JtNlCU+DG8tOJ
DhQtLPKHSppYotthpobHQDzqLzSXUbIJ29E2wCftLIsb7eBg1/jxBNWIOrrrLShEH4M9fbwL4u+B
4LAjBmhAmXKC63mbY6tzLmzlLi5/DwtJ/oyP4xMIbgnQjVDRYjSTiKEmc+++HNlUn1cHf9H60Wc/
hF9FPwfw0DZPSYtYYTxBTOgii+xFywrFFmUORNtgkCJpiXtWLSycHGyyVgSN0yNEc1fBrVO30zGI
kAecQHIxF+w35ayN0TgdC5Qoron0+sC1L5iE0U+I+6IeTITmdyhQ9d3Lu4m7lpQ3LGCRd+fVtL6K
1rf5FVb4Q36R9uh/CQyTIkuhWnxgSVJSnICRcLDSb44fWpcL7nIiT5XLsTemo7goZJ+gauVs9e1p
FLNbkVqI96fxnR8MTHnLP3H7P4GLL52cIKEXGyGR9OQAYGOMUg+lz/4QOsg+jIlkN5/MhqKcUxr1
1kFRKVf4d1ASQ1AmE+eHzzZEHJ/Q7CbjyMy2swSn/dQk2Fjxinj8dNMB/jvFa239OVcps35xhtX8
pPaITsAqRhM8E+TAzbcxdTQO7CNt4NcGhe6+Ovp8ENFz+eFVMv6AFn+3opPFt0eoYjuDpv2tPyAS
zlbpEaoVhlk20RhixlHnxkF9J4XTi48pEgmhzDeM1PIsMWkUPz5ty8OZ0NkLvEtmTaYnIc3Mr2Q8
TvreNHDxqlEmDOPkp9uLPuCjFblhXkhX5hKXKX433YzdWZiVwycb2rdQsTvV+mBF9JW72y54zdoU
zzU3GzhMV30ZCPIWMKBDhyMEJD338+cvWCn08Uux2OoHRkWvMslVF+k53AyKT1OHz3KjRJP9i6kd
keTSRKx7Oj5yZhmovOj+MxrzJLRqq1dsqF5vp84VbE0Flf5mXGMXzPZEZkzEg7hVEdUAEaIwCNdj
0o3jF+BIdKojBaqvlv4rF/X9WSrvB7owNZTdjfx0Au/gim8KwiTHuQ+GKg6tsds2KLOn3rKBKqig
5dDY2oy5M/yw3npezl2IGfqEy1tY6QEYpo829QEnrUEyPPx6WDzN3M6W7ihLf2P5qjifA5eee7jg
r1iot/Zw7Dc5xdwcj0pFPdpuXHYhoxOk2ieyvpa+aHWScJc0HFRLSajQsNufCKI+tA2vnfK0MvYZ
fIAzrNs9RCyfGJnSjXIklTmFmd9F1+ga9vmpxNItfsuTqZP7rJp4snXr2dHRhaZVrDBNikz8rudx
TV2+SagVl+kSftrTF1dJfh7VwLNfiqiCNqURplfLqovWqX8bTOmdcsGCn5Oyfp/1Nl5hsN+Uij3d
TR9dmjaIEvuoP903ljauf1OLyKwkxFs6A4Ym5TxIBEaC9def4Zq/LXu0u+sizgznFvb1KZasN5ND
fF2+GP3RmiCiQmsiyoAvJNOuf/6+qBkJrba/F/h5n5jGe+ROKU5gsv3zxTPYPGOU61IDGuOUI/Um
g27Sc1FdF8IE46N1l+5EE5ctWlVilxDzK+HyXrT9Ob+WhdUhlmyL+p36gpr6oZ9HDTNExOPUT7zm
twcJkvBVIy2vrL7Hd6Gbkd0SCVDVals8SWLkJqJ8zpigFnljCvUVQ2vT/CpJk21x6jsUrxUbuLCU
zV7eYHffTOBhi+ID5C5ExKWzO45ZBGIfLOJ9r2/a2DNhD9yLvunpGejejYZ3CCrVM2TYJLFJ8A9t
UoFdO5lGvLI7DP+6HSp+ncwtfccM8jQRmcI2wls8MdwEhD0wm6ovOOyKXGwZRB6vYijOKqq0TN5M
fLeOuhNTzkWeczfkWPZvXZubTdrkMOC8c/TCTHX1g1SeuIJ26djuOmPsxxTakoxJgLbxhpsYvF4B
iIKCotRf7y1ssbU53avsya6ZCBZYAiUufNAbXxYJvQfCuqpxzewhxw454U9pV0obnxUrs3gsHOHK
xq0EfcYmShwdoDHTJOAhnnct1CJLvPZZZLgLoJFWkwXzOL/UZzNZqz0RpYefFEUk2MRWfTeoZfmW
ene84TA5dIgW9unUi59x4Ml9Od0BFoimDPRYsUrEbToCVos26Gy54oRNL8ONQADfRTWSnr/YjLG2
Odh0WdTBpKHH0HoQ4y1vXE5Tno9Fy7JEE/LwxwLkGPwKfpdkXpG6j5MOVPrK1yhrlyqCvRl3dO0v
tfQaRoAvX7E8TAxpc5EoWM566ZyF2jNlhdVH6f0NJL3pHIR9tEgVHE+WuaAmdnTc2DXXycy5Rf69
P7VHZhZ55qvdU64NYTj5WjJp9UHC3iW/oa+ZN678IvuqfIMW0FnagMhQlLCaxgPD1rBl17zTE9zo
F43edXcbPjuhd+YjzF4vLVEmtjo4mX1e92zxBXpx9YRXYqvuvoypV1Zuyr5eiLLxCUQh1NJkeZzl
DV3kTAwh5SJ5+VRp+Hywu4GL8KO7oWkmpg7Nmab0dGEWiznaY4XsFomO1yWGB7X8+DgmHFBc5qzo
L+wAPr+8rOS29yXvCMSqvfhtM46CkDIVCvrTpUk+/lLIljkk5PNf3xBxMXO2Fvt665ZAwW8D+fHM
W6eSvjvMl+DMJ4xBfXcAMv6CwjESAEX+HJ9ULgkWRxP3ejzdyVXkt2Ljlh6Ravk+Uj3b24na2Kc7
6QEOXgTohFu9BklfTxuuRyOICO6YYANPluNXo9NNL7bwj5ZdSlzIM3PMggfqis4gDTz18hv/shJs
+J4iqkPEzTmaCALV8pOcr/8yQhXDaM95NeBBJD2yGKEdPhDCQom0Qm1c0JQmF0Hy0+GlKOIoVM/d
Wr95ACs7nGP5FDeilDINB3HhHGzI4/PuekV3D9bR7rZO/DE6iWUc88xic5I4Bl6Nm3EQRMOmppLR
7mM+2Vq045CmBb6wA5s9PPzvKSVAPFioEwxFaTofqlSgH9q5Uo4n5/aBHo697UWA/02wWNyh4LEg
yDU79hPk4Hb6VpuBDWGXlNF2yHYUwITVRQOveJ8h3dPGhLx3cTDAlUFY50fNywdaqQxS/rsGMtz0
7OSaoaMGqI6TjxuqpGothKEv244Z4EHeAAgKexRAk7EuVIaPnYdsTvnTh2PgLfBWHo9XAl16k7QZ
FR7PHzR5926mjLwaBKYsSH30Nx/1hTaYu0D/MyuBA2n7ZR1CM0v7NCt6BvRo49tjqJ599aTNlWpl
thct4ZNbeLzLjU/U1AJ4bhlxrGvhTW8s2xVlfLHInul9QrN0VhKD6oX3O+E4W920aGzw74qtDc3u
0v0g2HzKWJ+1K2znRu41YPuIT0UDLcysSELNqknuhA8gOyh9ZjpEW7++wNzk1sdF2CgF1xuN9RgL
2O+zi964Lzg6qbQsfqUAUIyN1pa0HaWqJ22KOFj8NI1rKiMHGp0ki1FCa8HBrm6RML6+ktx7l8Kb
/adEMGd0cuwBEHfd55xH29C3KmDkAAIjAqUfTcigmcW/+tqypH9/P5lbnbJ+8BFEQx29jzj2cgi0
dlgyfyKwOk/75AZHJu8Fs3+hJDAKI32WMtuo1Ex3C3e2+PBrPJL3nxgIrHCr7svr2F/4cvLdfV34
sIaS5055Rhl7KLRH0APMmPPnlysEuZZccO8fQVtm0m+8C1WjN35cHm3PEIInLiEujuRGLZts7/2g
4ufGF/picgLYJuUdcu2c7c3KVy504PKXboMNgGVrjFY8j8cbzEDIaHxI/wU8OD9KnYgo5kYu4oB5
KRBKRQ1a62IQZnpJ3U/Afg7v3Ejy8OvdxYMcKKtwIVOmaTiNjJgtKWa81zw6oM2g9LKGwtI7yWa+
m4NT9aPiyjwgH8TqtsEQQz8O7UfaVGhvfsd320tvitEP+oNV/4MO22I3Q1E4fosebnITYkYnRhzB
FhLXLy1O22Mx3CWO+RJXj2cmjyjDovwQAK28ZjEwnv59fPTZUSgnoWn2lbk/sMGKXe7UzrbpJSPM
lPGGhwyIP5Tp/4TqE21aTtHvLN+a8UJGuz1YtzkDVGl/wjjb24JkWIPtioK+4xaino/qoic/7rJs
Yn3UEm8e1AEK3dyGScdptr2rsMKQWaaPsUjUaPTUWLRKbLqlpMFTdzFVvPuFLOrP1tlg/3IJxDOc
/kNmktBHBHZoXT68iCx4D9d/daffdM7NrI1s6+50XDlprVcxM92hJjpHF0ky+nk/bgpdiFEkUz2E
iR3jcUtlS3DqcKqecp54Dxl0zNzIrHIAZPcTpsPXGkJ+4teIoLmbqvNcapOiHqECJ351n+hCbOSr
S11WO3hSZmIJaIWFrcT/6yfM2yEAnwQmomefpkatahO1p5E+ykctOXSJA+4pLwiGINriIt0gJrkf
ORijnr5WdN3ODx062NQ0JbVKG06V0kmy1fZMmawkNqgFuBmMaIrPhBpDJkrWO3kM/axJ4rgQhxks
77ZUj6siisRERpXJR1en5C8xwNmATBrQBFivkp00UCujxzfk3SD/A4q2ja1QYJEnEWJz/Q21phZ1
LUstjVJ17CyESNMH0/cmn5dOmnL2kDIy8g3F0An7eKQAmvGwS19vr8BBteTW1z/zb8sD+lfL+TMO
oBaTToGnSDHJk/+GmjqhfEP9SUYyPrp7DPkxJjTSRV6wpI4o7JeGVluJq19Y/tvV/x756g5IVQHh
udvmYNdN+JlR77r4P3YsVvwcHxef+agCkLlg0AerM94Ce3K9hXJICLgjkxGvcuQHKJ52SvV613VA
LjjNoX7wMYO8sbBJaUYMc3IDw+KNdGr2WhF1Y29gcXgz92QM/CHtCGIQEcvp7JOwv3vmgTd5xJEY
JPBykQMKfRpr2msarlbNxsncc3pFM4AVGiQFVzkZgoHOiBOPPolMO8G+6uhMD1CZUEM/Ua14bRab
swDv1fNqklZ1sDJ8vFgFSk1kxyhMQLrRofkSdgIswgHTXfs+ivu19nMCbtUvzSISs/1dqzPU+qC5
fiQe7Xr8Xz08u1triswnVmue7ybuBNGLFGm1t8dvqOAK5eEGOUCWVPO5NYiAQH1c8fDs9uWT5Zqn
Zdc0WbNXPst5OADxjn31uWJ8YzhQFL2DsdJbHp54OF/TcKEhAPeZhzL39buUvV0m1WgtOOMLdAl9
bJWZe6behTqiGrNLeKGhTFo/LphV7gG23Vs2aNdkNOgOQ1Ss/pAEuUwD/BnNlRfQqrYmPYNtT5LT
bdV7hizMpyL2rKYZ8XRl0Dl1Mleh5zpRYbQA60b3T2S6FWmQEqGqqh0AvAMoibMnivSB0FIGsaQc
HelmXIMfET9XdCKnHcJ7hBj+Gt/WLITWmQwhTIsezoqFyD1U8F7TFe4diD84X9MGi2jOMVYUzruh
5mGGVcn7HdrSWKaAvSyKmYBAN42yiyjSYrIDG4XVHXNQ/AI7Xri9vOjCwK576EKRCnyomY1d+fVL
Kwalq6+TRFruXsO9QJrV/8HCVDWdLgUPJM0kS4djRbXVIF56P1M8R3s2SRLtHyXVya+udcX9t4ov
daRxn6kouvLgaP2QNOfGs5wN+tRFpYQ5SdI3faV1rRAl1BjY5PW5mDbo+RtkIEFOBAEqPETWGYX9
qekrKLruH050ea+Ks/vulDvPFdPA/ggvNFYr6CxRzqpoEBK6q72EBDw0z8mpSrTbTxAgc1lKq/sT
izBBCvdwKpORHFXtYueBRJPBBJ16vH4PZtHXEQoLLcZsAyx3voSahm+46kn+Ma8Yl5CLCBbY4dwL
u8dyBdKBqZQZzfIWsexzZ507W4mC/GwlgiVD8vOrp2Lu258y9c3QIJp0MBB3qf97CbuhdpYPVLQL
gtjK6L/+2Ph3auCYeEfHL7Yb712vxo6aZyuzT1cNd0FhxlZXXAtB5lrxf7anO5DxKMyObN4GiO8S
jI0PPwiPtnvOM/Le3/s/AVcnutmi0peiIkuwamVzD6Ige8tPGLMk/Bt41pfVHXuGlCn3Oa4jHY4+
QrDlGVuGB+9iist6zDxpYZ4qRdBRSv+bd6vGu6LE5jZrlO8pXrU0VqE4gVVzsAHB53N8/jxcrpBE
5ajk+mcpF/KRAoqQc13IRDDcYZzNcEy39x6cu5hVZIaq4vapYenEZJRLxMLjEPHr/OjZqW0TwL2k
b+b2BIR0gMkfCJF9CIzmOFmCsjWyU9USX2Fe0UL5LFJGYT/yLuo/mccNLjRuamZ3sa28Ke/CiTR5
jTce2m85WtvrqFO8UYOV8QvFxp0x1oDtsq5VvFfZrTI7wksyo9Mr3ROcn2CZxzt91AHQWvZT0lED
CzIAXFMRen7hZ2OAiDVX6qwrz5rUJalbxrs1jmBDylZwFfS3VHBxEfzhny3vfNqlMMrKtSCjrqC5
50sOneN3O+J1UrRIDE1hYIBVYebE+yCwRoIrCX6R8XKmmdOdjk6nLD+2Ba1afqCFbpvamr6ZCssu
P0VIvDk2BOJX+k5dDL5p0N9a4WGg9ixKnWxBhADVa77fYpBcnIw+h2XwgdOPPpdFKLkGGfEveTOf
bDEX/9zEuZTRLXFdQd32AEVgb7FA8X13DYIXEL8dzDQq/fMfbZ2SohEFcK4jFtY576FIfdHbqOWC
G3xlKaqGuiz1x/20R8985E9h627ahvtD9QwQKLqTvjgRWmw6BXYuvLKJT71Kxy/LQZwY1ZYtIcsa
oGBBCR/sJhvc/ImZsDUpOriI5AkLUZcVl2oUk3kXJaxYbtcz87Inxer+EA2N7qB2oQ0FlEJrq91W
L4d7ZQMdHBG3bb0KvF+BMUGcNiUlT8gQecocW655roTdb3X2dIfPzNEitZqRxoZUDZx8BvOEZ9En
mkulk+EWWOAJHqDk5OJtfXXR1ZBTkYg6OA1M3zktEZxnnrERtFHQL3srbbmuZPwl9tRAtX6uMEhC
4IHiyMbNlf3Q6CxfYtxoejyfDQmbD6seHLkNvtGN5HTWYL/JUVnxdZDQmZ3D4fFlwpFLfLZ73zeL
5RILpTe8C7pu3KphvzaqcTI2xqpn/0U2D9qxO/xsqtPW7I0YiPsCupAI3Uh4VT+7ZSbNQU/1dJSj
q7WkkNJjCPeYsmM6Uot6hzWsH0E6V3wpkemtBBKt7ZZZBIrqW6qewdMzOvN6p93eRA4H9HRaB/3d
w+P/J6nQpkFfhVbo7Ob86fHLpzVo0StHNJqsz2mwjv2N+Ultp7pm7drl7vO3dfgRQwieOAXKqEcS
IXbD3UnqMusgZ+iugA/tOwPF8FdOgL04Kc2P5zK5mmfiRQS+FabLmPFDh3OQlSLgLjTzkDAyta0c
9S6fE6IxKfohmZBVtUozH9phtMQrTaCnILQXSE0dDDDx/H3xuaeIUXR+cGB4ICGNuv8nHJZwDNcT
bDisJ7cXm1O50J6mcIKAPhjxKFyzkJHeFy4u2DWABfBqv4s8tJsAHcwPwsgDTbTuowu86wkwUOfe
fICUaVfFeyOjMsfwmf2WapLURiRma58v3mgo3t1vsp7zkHiQa4dW/BKjwvQBBIqhTc4GeTWVj8e5
xnBKUZFEsau347jRReVtVa9kJV9OBcIljrsmh4n9QW/OJRUYpnVZ3C/X8zCCOJ3/nLcv62g2e8bX
VzNV3pDnYiAhRK+SV8jTXBbV/mW7ydabVifHo4OlbPVaqGzvr2k72a8LZ20cumUhpVwLc9Ptavgm
QT6mf3vT84ZX08OQxL+w7UloTFosQHj/b1rjZHpi70pnOo0oxR8vfhP5B+/uxf94Az/LKJdk29fG
Rz4OOxxRuHFEPPV2DEReROTP5vfWwYdhiKutsZ9DhT1nESW3P7mnSUsw1FhPGY4c9JpBV4GC3zCj
FTOpXl023zttqyrp5oM8sVnoYyk2JayOhjj6LyAEKu5bVJ5X2T6kVHiMIVj1w+iaLkDiSe8IgWNP
IItzr0282/1+Jl6vG/3hNvDHAsJWyqdA/0SccRcmPIcb+BN7djZC0Cge8hnM2FU56HgjsCfNdwRW
TkLZL2wqYN8N7g2FiqVdSms787ZC3iIE1/ToGgtzyPKfMhoqH2JaAXOLUOL8j8sJYR1vClA5yxjF
OvU2XnvkSxTWgDFFkFdNJBctnzsOxI/2dBePNvWB39f80EV+PPtHrsSe7EeonvW862wHEAiCs1a4
MXpWxbmNlhyrFhRnbO7wX6xaM6jnLgeSKOg+YmoCiKlYxXzZKwTLs8ufx6aLNP9TDJY8DDzIoESD
ibPzu099ZE9C+UqsCu9cTbs2/UavwZFyeFSqbtns0dKXK/ducV/FRtiNlr9iwV/MHo8z6AIQE9Ai
lBGrbLVLQ1loac13KPj5knY2BYxdejYV38nU+5UQoVNAMy1jC4HlY6vKsMl2lAbX9OGuvCVzoT4v
qCexmvchYLa3UoCgD6nvqzKyo1/OjUw5BwhXgC89wEpTE01LEBXxnJbj3GanA6o4k7oJW/W8LJ9y
bk8UegSwu3b6TS50vzxZECBrWfEV08HFPEP7/mFX4+rJdqH+RBbK6AculWpd1kRc3Kw1c4v0zKWf
unSCBQzWTTmbRhvXXkLLZVXUvfrhDoGhQ/3ACp99Z8BG06M3dUwNu3E4rkagO3YTYY24e04mKwOU
FXqemKHTcd/5Noue1qZVIBY1P7cssP4P6PEu4TeoCjobpnXy4Asm9OjUDw1Th7mxm7xYo/Jq3UJU
LwEHRmaDkkoGgT+40g78x2eFBowW3cC9MsC3JzCswAiBEZctDsVxljgfJmW4+nV+u/R4n5NC0YB7
ivCIFfvrVPuAgMnDCj2X0kepqsVPB5/2tNuQ8lDdlbBIvO+Zb8AYcRWUfKuj1A8tZSx4uKTQXzwG
5yth9FwwkMpb/gNb/gfDKzQ8c5Z6onj3HdhPopyegGP/T/w6AJtUZnzua6t9PDaGVuae1tfgBVxC
16ZP8pBFyToFx3rGb7HGtuyXLMePYPPgNHDPX4qwqxdyOltsi1fqXVMkrlrNhF/FK49IXJlkfL4d
ht50jduKaNhjoPiq5y4tvbrBtuQEsvO74kWEC8uawDumL6NcuD5StTEm3hqTXcIi+861o3HoIl5W
dX+r6ALBP6eRKrLloqY5X2FQR9y8pJV9aK9iaBiFefVsZ2pG5/gU2QL5e0/jFIxP2aJr14IoNKnK
6RBs85z2xlZKJflbrncN6JNiWA0S7n8dshKnbOvPWtrpzz5NtmCLOxnTJlvrg5ouezgIDgeDOwFk
20CsYnHLFZmmmyTM6NXDfbzGvAfiezgUHWEPviS7q2OWom6+A1L0/Bf9o5PaHbHFIJiC3zygQXAr
hhNEkjbGRJ4+JzaexICdtR3/FxhQek1VDt4pVVHvkL5tZlj4zIKKMxqCyBHGxsXKwEv9N99QcZu1
M9fvfr/PnctuDNyansVpBEUPrBceiJc4tfTHu2hbxX1T8NlnQ4eChaG7XYN2jwAVTGnoBISG+d11
2vAUAsXeWyfVcX7gKQr5Af7XUs4LOLcMWyDP6AcsU60IXOTlGNK7cI0+Ey0AZ5qt5zVausN262fl
iM/f4ENWlCW1KCo/+ydsHVp61CS1WbrkwF9Ai6qJCAA1MLqksX5SMwfnaPdcH4d3kD/5HEqK+/cE
yOlOUuRijbxNK1iSqb9WwPK5X+axXdLeSWpMD6w0lfxWO/87jSDwNY2NOdsJjcr5TqXDW/mB2Rcj
O5VzcuO2KGbFGgtsPaqF2b+cGt6i6z2NmnHaxLOFhAjDuMy3ADxSU+FK32BwbbYogGQvkKm8ZtcG
cn11Ty33Z7AR6iGQIrbqpLw0lOSFs9zQSpsH+zZDDaHTuAtqptlAvV1+xSprTeT1wtLRAnj4w4uA
MkDe7BeIttfiB6XZrXSYA9p6QDcG8X7S9XILRqhZ3mY7gNANp2Sr5PCrloFK1le3TzanCDbEX9Xe
qtlFgrmIgzg1fPx5WceSVDb9a02aSrJekUYu1cIZABtroiNIrryFCRKVnkxw1/ejlnZojOJyhDnj
/CDV14bmafmyqBF6Wu7rtmaCyEnOV4NFs5MXEl0L/LElvBilejKsjddvf59mNTA331z2TkWH3psy
mrEy13nOvEm1Fv2h+T2gDD6fy3lfzwtKlPe4zGvr3+VDPxMV3ik19vthyPJjURcmF/YHPd5SXSjF
hgOg/RQF6uBXMaCYXIA2+ZlvZduy0968k5tk27sqE4IuZq6iywWSYYmxQw3lrkaYo35GcyyDVWPp
/xxobCDZ8IJJQvGbI9hxxV/ZB7cZMx+rpyIIZILGHofOjCXiBvSfDAuJjTjxxMhqGgmwGa0d0Bbq
UxxPgfpAimiNVl9OdukRV/ORQm98mHBrx0lftMpz13QjzPp7Z4S6q22WgfNkp4g3IgCHTGpxV4AE
aNogNxiIvcSHPlj6lmp+k4KpHwpftVOfDTAmobH+Fv4MkJPr+dNa3V8kYADSVU/5OYOpe8ZTMJN7
JXX6nEjXqzruapDFE0WVA8FoIZkHwK6U/Pg/8oQBV1i3NpvQ0fgL+FRYrqOOkI1q4gR999v8232y
nyvAJNRfTOeMxbsH764996VY0ASja+q97mMcpFVdQ0M/NSHW1eCoHZ5mlkAdylYw6eINj7LkTxii
Nr12Qceg6enW/zoQPhOFKTV6sfuXbQTMnfPW06viJ9ORCgrsR3YLIeUSxhbEugBmwXaPsWZP3cB9
+RUiSPkON10bmjRzLpROYR7ZxA2k5fftg7OyGU2jTSlXE2i2HHzmxCzfEJRWWs6layaG7RPsAlQT
SAcP9LZ+E00oLybYrCl/cdbkV9bjk72be2Tmuw+wS/ePeoPERT22eoTyKq6eTeNkBO6JfLY1OrPz
pvy4s1uhBfOm8D8cyuh70HO4ZbV1ssUVOg41mAHxMuM8CiBAXo6o1PzbO3PfOv5DPt1Wr61jR/vg
ZqVLOzFchMwb6RyWoBmioVudyc2X6R/TH+CXI7VcwU0WwJ+bgxoxWC51BiKsNUUoQJJXAJvxD8+w
DmzZ5Dpr8DUixkXuaypTCVlYtY1zAptTatz1+5oYOHmqHXNqErpFqJvdMLOFupLqRu2Zopa8KfLg
v7Zo8j3uFTpDUF9zvhvnYgZzaHG10UP8co1yL49LBanYFtZ0G7E7YbgzogtXX7OMPASGtpV47Jjr
oYTJfoamLcx7uLTrPTaqJuy/z57ob+FwFIAVSuoKTi2s5sulDsRI3pIog86G3VrYUVD4xVlbNdIi
Sy7c2oxNbEhpi8aquYPnwNp9To7JE9iiwbMhhLo2RHds1ery6B2s4CUHT2mKzcFC+qwNdxgTw+wd
psd9pci0NRlrHz6SadTN94lObXUJSr7B8Pbu0RPzQr6QCHwR6pis4sA2tmxCQ3wvyrKRR9rCz5l6
9pnJVfN8+HFkqXVm6vZuDe77cY2xP+0NbQQ6SRZo4F3Pn15F0sJKv5lArkj44IQYbP0Gwe/Zi9Rj
uaiTbQIa1MMx6ylq70bCgX9pzzKKspJ39NBQGcK/g95YqNviJbxv3BU8QeKvZxH4uRriGsUVQQ5H
zKFjQKKbvH1BJ4hoUTqzfw7A7HtmOuq7XlCBaKNVDA0GtaU8OgtLd+HKhy9xgigrQtmTaZhtdkHq
sSA6yni6uZN+S9GRQTIPBmbbbR1I0cQWzo7q2r+nqna0i2X2oq1bPW+8+G96Zzz0rQ/dCxxTSXyi
q3CD3xNNtjjB29hOZi2ggEc7E0fUZPRXmkTe5OFgShugBRFlWp+DemoOnHmlxfUTeLJUofTL//sg
1rRBgDeJaGLfEknN5Uttuwg2I7bJf8WQOkTjYw9SFHFzA19QGoYWQIcMGiQ6CjgSyjshMeZfZ06T
pqFpFYBjkuRCKaZoHUy7HTVJUPIPTa+GcVhot85sq2PllNdQFFef3CXz/iZMfJ/8HpHpGtaMgFVv
MU+swNxob6zUqamhI5ouFmklKs+OmWthUXccWfhsCqsLW4Vtd/4hiTazIMfEy7BcUOWHNLn8Clve
yT5bhkVxuw4QtKhb8AY2i6CY/5d1bL/EyrWBkxiS+9JzoUKlTTC1LF4kk7b8h7N9TNDu8qvSzwy3
qNLEUnRxKKey0WDYzuHjNlRr4pG0g/0LM/A7FxgI82peO1EuCaIoQeJ0DcJqGpH0Bu1ioMZFAlIe
M2xN6Rhhqs3vPM7JESt0J3YstdtDNOLs4YqZ4dwSrTNL8Vz0SBvaoQ6mhrdEuENMeKA3H6zN7IFm
qdU2z4JCpT+sEzyHjHQXFYG1BEgFyBPZmnMyVdW4exvsKO8K3gK3hRuC7QxVTSr+6UNQy7GgUGCn
/HRdnAuPhFSRpgVe+845pwwocTl38iJGyHXpO7Lv366bBgRW7cHKKl1CrV1bweZ0WsreTr0ctm/m
RuVpaIh9c6fZ2EX+tU5vCghuLsXJQmXNmfEsVXOHWvRd91hFhnx05MZf9RIlZfNY6FYg6Xk1mBTb
8ASyg7gZVsPc9ecVqzuxoqFP5Glgnhh1PdUvgmUK28T7svkvYflotUgwosjj8atSpml8hLdNaIDM
KqSdl4tP/dayxpOtI8kEXm5TZmx9Fd+X+U/lYiJTqQxrdJIAENjhX2Jv85jsoRv9e3bSjt5KQB1T
QDnUHu5TILo8dp1RVER1S0gI0FXVlXECLNplxos3+wZM3zc5LkINFc2jjNgipq3UrgCICHpjCptz
ikEENAujqJ9fSIHKsgi4aCFscbIwDoI9rHIuAxeI9VXMX3WvKZbsOQ4HveEJTl6l2rYniYG2xwAq
PUctVTAb3vNg7d88yEs786ctrmSZNvWbGyRGlASepyd0aDvVgXsPD323LDuaUTl5KRY/ih/kwy2c
gF1fYz5WUu9uXDG4e+cLZowja5NaOb5ZUgOLOyNhj2f+H8UUOmSk4V2aI0qwV3oUbaSquaWt2Gm4
5lwIdlN1wWHzADkPbS6/lxJvDao8mfe/bZ217jjOHziEKnWDRA3f6fTwVC2Et9yZbPQnUAXV/xtg
BNHv+0sG4UaBKKp28A0iUj3qhfrntwriQJKMcpZShqnTL5UAxpV/ShOiYeG/sgeFhtDQU5rwjRlf
XArL43vkX/vKjg8eLqXpI5hU8YkmyB7TFHqBi42cAuTj4fzmLmUFXMVSdpHttdibLR0rcK5WruF8
CgeAUdbt5cC0HfA/98NehddRj3EgHWMzLpdEXTv2VuLg5+atDE7I33cDERa5WiWQR4L5U179Aw2F
H2aQC8ppL9XPPgGX1ZyWM70fzT4S+zRJKxv3UEbH4fQ2mNN2Y2mben9yBwT+Wozt6bei5KsRnnGA
sINdOfSyhqBAU0MrTQJIc7CZW92MBR4uIZpKUyeuZsfYtyat7NllP347N+LrJ8TsfKZlmpM1QrDg
MYkRlIk/HIl1p0+7Ag8h0ZKwnoYZg8koXILaQeOn3UDhQ33XAqVEnJNVvHmbgMAhM6WVoH7ILo4q
aj9LGWx9bhwJZm0jQHmaM9+8pXff+yI+d5PxSrwIHgbrxdbkNnaQIRE57PzFnMHMUCZFzS0G1n5d
QJp1M16KTt4vaKjpoSZXQILbIBTFqRys5N8kBXZbzDOefdko0op5qi2UFFwxI2+DCebX0NMknd/1
PG0N24JJY3HPoweQZsYcQAeiMABK09sVtl+uzds8dzaambNNNbdLFmCXhYRQ5uLMCGxctkGE3xv/
nFFqKgQ2bKBNzL7Dg6K7/jOUEvKjjfRu5MrdSkYbPhqZTdag6dvnos+XPNUQIhEqoutzyoSUSevR
tQzSdNEF3t3CU2Z/HFNWNn+qVySQryXhR9ra5m5Zc0aS4PelidlvpFsZ7wBcjMFvHZueLE8Kjf2m
i9jbtMXVQXdGUqtDsYALq59MehjEdmoEPQnXdQGLut9PSn5fcg+niP/C78wicxiS6B42wPs5BOAT
jNCuuxPy/zczajXjxgaybdBU2M6MBHr8mZtRPqGR1LtJ0P5naTjRk6nISsL2GfrPNZEf1oz0JiHm
0b+a2YfyYkAq3R6GEgRK4o/HYGxnNtqvSeougGZkFJ/zuhNSrjXoVWCiAcslYitpurAYEdrVg/Dy
YzI25YtmbgLF0o/gDdgxGz4qDefddSN3AHGUjb9C2PLBURmWR/rSB8Z0fBiUxIBWGCb5uHO3HQ4m
MjWXG7PuXOrA4tMBJzc4VIfbJ3Sip4jZgwvzNdCM0AOeWoZ4nxRSsNKbSUMemclbejfJncVlqV4m
xL4G3sx8m3iq7DfH/gLm3EZHVleCK+wKoIhyZcV879ybJ9yB50aLp1WcmgLob0wM+tBDUBqHzzFF
ZNyrvKKKQOgFR2NlQAGrskQItVH2EEWSStpR+iLqCqaY+5jAUNSw6CgmcR+5wCfgIuPnvmOzhzGz
Rs4Lj+Oq5PIRb4AqYgeTYw+4Us3WLNTSb0lNlLjDjwewKtU3d/VXvzQBy2no2eTID2V/9WDbwarN
nQQDpc/Ci61YR3r6u2uFBxRahPi23evgVkjtOH5bFzP/N0onR06BlExe5slVgjlDQe0RJdo74jrb
816yynVL0OxmOd/FNOb6b+2xS9IoaZn1EpvYQgiOJOGv+rQZy2aUkG8g4yaSP42IeYU2wjDcVHK9
Y4lHQJU8ddUBdOo7PTDeUbbFFKIlatEgMtERDUXFwzogeteXDdm3FCoz5kXqIRs3fGnJ/vF2OTLf
0vka8Rto7jFBJxTIzcd2RM/YOXAhmtrX3C912aiH3/WKBlIeh6KYWYargB1ejVn1tr1EAxnxQqw1
FpX9NlAszLuJaVoYol8Zf1P9eEx7s7QCh90MioYRzcy96RvgL9M84CRiTukBjfDxXvPgN4+kbt/m
Ha1zkMRkMo2O/JpZgmoIyUvLA3NmyqViq9qVA0bbMpjSH7xdRd484+tMWVNnjLNwCNuody4HiQZS
RQRm//tzcj6QCAv6KE92Fqj1eLBMBY9dLqDG4LqZc33b1rJ/zFbdz8w8BzMqm5e4P9RixP64/HSx
1XtcJ9yNrbDOxWgKfGbvD+Liwejice2oZHnMWfcMKzjsD4e/OZuBov1Y8/gb5GZqC28JfZBie+en
18i1D6FhJArmAhkES00arTo4ZQ8BtXFulhSMKLSOBcrMhOhl8ON0ixY32vfijlIUCL5El9QiUQh0
iE77a98aaxAD/A0uYDA1ryenEoD6QcIMYZvOok/6qa6vNVWAMiT442hATZ3s8tgHGGdtNvmsG/ZT
AU16PUMgRAFnHtAHndMKWmJ4b8JG3BbawlyV3W2Eownwk4TlXPWzDW9bX7eHa2iVizRiukgQarJw
1sJ0iV1KuDWwD7uWUI0r1OMry//uETGYmo/7UU+sXOsrVETydL4joQpmUkHB5C6cjmDdxkhPvePz
I4L2nl2SWdHx4DnIvyV63kivrjZqNsJlD5C02pY8aTB6pr13lqb58ZOawyWHmkHhHtx6jrC5cFD5
w3bOYGEXwYnxZhOl1htyw1DZyFxV/GZJaON1NYbHdgA4kh/TXaDKGSnGTR9bd/sz+MRHccsGxyu2
0h4jVHmj/MvG7eNMWGghSp7YW9wBlGnm4rCGF0fs/Vp2IS7q3IW7xQfMf3TsHxkNt28GBRfUMAen
PtfHLHilhv3ukMNrGfrz7jVRBAZP/HakgMNhnjIkb6XKndI2VRgvLHZsk6m3nmus6+wUaRg4Shz7
Slq2v/AltRJD027w4xk4HbnJMtlbEE4pY7JTAEX8Gr8Jks2WeyikuiHb/gLTikJVxIsmGjzA9E0S
ZDLetHJWx5Be6VdYwVE5chfpL4+AE8GkkrbA80/EUVvVnppQVZSw57jAnAHGnzCYihR/TyArSHQN
98m8Qv34gEGjuHWBIiMDz33KrUrgSKbg1D/KT9KilOFZ3DVPZ66p2UO9pqrqU7bkSAULty7knB+y
N+6M6FZRXav2uKn6WtQ/5bLOf8EdDURzcM/W3PHYgbQm7E/PPlLWDLvBIPlLQA/qPMHjvGi1k5g2
1yV8yUJC2Z/b232c1iksbZ/SwLoNComyhDzZfIStbQ5Md0GHoaWFLZi1V43YeYer3FMCItD2S19C
HzKEKnI1jF9wRw7WkAQgPF4jo/B5Kkz7VUSBVRJ9zzk1oXE4PEQqJT/LsmkJDiPfQ/BRJg3NrDuO
v/UHBTNUFAOnfn7coWEgG5i530C3wl2vey5zsc/yTPNxweC+l1pIpQBbNzjiIN2tIb76+uJLRu2R
auDMjDphFANwiRwu4VPfifMVmEZiz41QtLIipOoLrxmDMn/2w2CtkLlS1x07L52FTzZzxMvEjZ3s
CTVg2B9pGSoPTsriWGdAzYYvxIeH7mU8wk090V7yRTA2HY83BWUV6Pmy/tIIHbZrH2aqpb/v5ZCX
r6E8O7J0uu/0symkEIWw+n4EdO/q1rnMJGhIoITSVLqbpiI27s9/U2CJFhGLQQrFZlkiFWMNTcMy
t2S3MCbmjUT5IHZXaAy0Ripo4APee1/A6ZHWjnaxbg3nNzsmDvSvcIan1K2kQi69NEpL+dME5HCa
sjK6KC2p6NgUYUajzvwZpGT/a80gOSBXM+xPLl5SBvM2eoNhhevNbb0t7RTlyzupdHMeloN2Rk+q
TSN+HyP9czH2NU9UuYQQtHFIGmQKQ0a+WSvOxwTWvjdnqWMLDCByd/OoQ1nNNVZgK/Ql8oJpzm4y
Is/v970LjVhpVqEzmTi/nTTEgku6VJvn9uJ5+uxxmnjul0EufNP37/EVhHJzijMYKrZeBbtT4PVV
TZXhU19Vx6inV4gzUkxOP3vPGenvupiPECWmA080/7Ovf76Le1C+yMEwAUX6MjHJSZh0s2c+mRfT
pC14vmEJ75Hju4vDW9TGYEw3K9rJcsVvN0Mwb5huovCSZdN6xnRR8q/SXyfIzgdiV8BBCPJj7oU5
HXjNKCeKZP7+39ICFavNOfCZ/piL06nb9l2zCNcanGGw+8fEsWOMCRpAhrDtqDO71D5sEQs30/y8
8NP0SVrIwzFmuX0Tt6GXD67p0V1+i9K3i4kNWC+b4ElTg7VzdWMofAH7SR1bWTqJykRk+T+VCTLS
hVpb5UKP9k3yXcHowsudz5Sk2lmS6fptZ71QUHshd7R4iQFcHWUYlqd/Yrb0mdI5gRrO4Fuc+0Uw
ovNuafG9XZJFSRo7pMHlPsM1rk+5ZkAuiiXT/7ub0wFX1n/rlzpjY31OnnewFxihcSFOKCkZeMkk
QCYH/JDW6kdyQ6rS7y6Ih4LsS8V24d7In92UddV/F0sJtkCKlwWmmjt1MbkldKDCpaurutQIpOHU
+cwY5jljSB5juiX8po657n87hvZvNPn9tiuqsTzDmJHAi12DFvbASvhhRAvymGuSQ8RYwVEWGqJz
MfkwRC8Q4aWrWzU3EmdCEse12HvoLutYdZgKp9M3oeJKkNparMN93wuhHWuJcmJ8xNU3linirkuV
dd+DIY6abK4Sb5vXVoHWG+760kfsIr1hj01wdxPux00bAJDiicUAOvboHkfrZCY+yzbiXhUTdlpx
P5uVKMPUClV2lH96Yw4Z1WLFSS/gbhxpO1QpF28Pt6XNYlG+r2dX9esFwBy2IeKY3IfELpSk7MFQ
g9nWG1RHtgxg0eWuTv2AA6kIbK8UMZdQoOwmW3h9TlhUX76H4Ldp09wTF6vPeMi+KUNv5JyTT6TT
d5On+44IDpITRbynd34tZJO3UetJiKFnjyYysEduYEsI687CPOihGhSy3Innm5Zv01yoeo2FfTe3
+ROtDkHG59CcVdaaTzd5t3zBnwiO3Gm0Fz8iO4qmY8HHZH3f0HWWn0Xa2rkOUWRx2F6us80wW6E7
ISmReLwLkgOlDChlcjEQQntiuc9mL6b2WGMD6LGLLQLP86buwli7DX/zQFNpg0zzFuaWLghyawfn
gpN6Gi8IkrcDvQiijGUW7gyUAOEpB+waT7hKhtAgi+XWGgd9EiAg0iCvXVfzv5Uv+4JO0su2mYh6
+ldd7rcASjwCQhpc+YYn5fKQEuguKMHUzvLFhmHWcQC0DxUgrlygAyam26I9bj4WONzBoh3w67oF
En/dIsx7ogtErcGlFBvxL4dVPwUcRh6N4eCFNdyiuY5+ZXaguicP+T9va08cc0COvPlwN1y6Qjhc
/hzar5/Fm/e5fHQZScLcwWBoNnQdth5Z51frKqZvHqf+jdHsivuv3XJCr+85cggzUC8U8nspSKPI
PDVXFfN3vM2Ak6moZPxVuaiXwGSEF0XwEpxMqz+hZozmRSoVgbXEuz33yAshoQ2Ky5fwXbTFjZMk
La3RoAP4PcnNwSHoaOke8kNvN19keBM2SUZjRLm8R4lQKYfJb79CJwZXcSpYOLx3f3yBXLfXZiMB
7S8QOj+z9IRwg7swoewZ1yhpM4h5FxaKbYEYjNgp1m2YFutg5i2HfaGhPea2mTW2aTFs3IRy9k8u
NNYXeGPSAzo+/mvtQfwGaZiUS8hOhA+i4ybTLucjxB4Jf717fom5m8neylO02PDpBc+zDK46UNVr
MtE40QLLTle2JC/OIq36qjGupUb9t6JyR11jXcLshrq2EjpKggyT4navZULqKJB5D7r5WuwGKAIH
CS+sfuF8sB41TpYOL3RSGYAZEkwnNSjYzeDBj8MjNE3qhjMVGi14G5ZwHHQ3EPL/BZmtmNqNmrph
FH1k1ajbXHEEw145/6BoJEJ1deP5sG+PqsmvPZpeouWCYGTm+fLvCbHoouEXo99TJ3BvzZ4Urt0e
K7mt2aFtuS2tEYBpraB9nfE6dq0revCFh+RvRXYPqI2NHJuxQz5LLAK0K6sTV07alW1oDQAOL6VK
H/RoeL9A9XYbMyFl9sDxOiAkf8g6qv4w4TfIbIEt9+xOodaCRVkro90glJW5EAhVFJViUHAV6MVz
n5rIO2HT4aGw0/uSGIJXpZCaUGzSKB3QHyJcZ/zmmTd0dtQa/U7C5J20KMi9hXVVLeqDNQckj0nF
h1NEVtC3/y0rJeDW13A/DG30Ynzbf5YSugJcg/wXOIYnTkXo1j6ciTb4SRTrJ+XGj3ptJvpnMkls
uGpNQahTG7Y8G2jfsm8hSzO1/9owUkgv3m+fg3BoAq0+nZcYP5ZisVgIjYClhKzbywRczYbgJ5NS
0KML+Twk+tFKPEJg2THwMLcqzz1yHmsNEFj9Sj81h2QYyNzJUA6lcUgi8HXlSkKPkgdRs+bXHysg
JR2as96qL2AssgZ3BzrFhh6GkKELy3pQWxtarjq3dDLuYLx+UIVFlyrK/hPoEATxVlNyJyyPP7AC
fyTvI4ZP43et4Djz1l3bM3s8j+wH9HtasuJEi7bEwgorJtKJOpVHVrrwBOLcqh4bbgx/8bb12s9m
aFxpKKOqQlXf4M6zBjBKGkRB4oCvSIxczoUIcMcz8vM4gtPn0/JLA4SnDPK6LQBczokfT/4Etn6E
Ek8j/9R3gUINuLpFlIKyefcxXaqLuwQa4IXBvtAJsDLVeFA2Orb5xEzR1Wj2W9eBwTIwPOzt6FlX
NGowsRsjqUgLsoHqsdBRMpz7U4xb8vBby++h5HDzEJEi0Q2J7Dsz4XKBjmgWedIENYHSWZ9OFBES
TawJqaW5TSVxhuD0S9m/U1Jm0bnJK+Xymmuz4qAmx2voxMJC238Tygo5g4vBdLiGL4e7ULW6dkN+
QKdHlKvCmg1qOLYPoIomCqhtANWJzXAKVOrD019Bjmwy0NiLvtCBs3yv/jwBXqpFA1IR0A0FF+wf
ayqwGSfDVEH5hVuERm2Hd6bAvwRIcFIxKi0/Pc2SbeELdFU3KoKurJwh+rdVZaoIMGppUfKk+Aam
E1di2sJ/Y8sC02guNdBD+NXULGDOQqsJWfUbw2l0dF2d4AEUCw/gN1jOPW9GARuj5VViJll01N64
iNvgJ1Og6hd6/4fIxunyLJ1qn9c7rYfT9dPfoJPdHkDxwX1GBScr8lnRWHcyWhTl6Y65Kh3t4aHd
LeIfVDSXZBHtQTmDMEH1Yuez2320Z2plaNuSgeYU1HBF4q6gUL2QeZkA34ZU+22wAuBGinDrpJv1
OwzUbm5GgbVx0ieVzRpOlVc5E/7f4nCpabcABRVsaVq4uAIvQIURYljP0KZEnUOgX8gGikyDHf1D
NuISUrRTToeGvfD3ABQeOtkoU8PUwWZYvwGzKVw1HikBFZTX2UJuGwaoSnFUw9w/2+gOaieHjeZA
ktApwscImLlTFP0IrK+Uv5TdV2Uw5l+HcDfJLvASE5iC7yqIsbvZuMtFxq8N1zdS/dCq6qzAw6ds
LzjZNPFqz5AvUc7fMwp7dnQPmKiKpHtE+/quMjPl81DiiOrCzjiOFxo8l/9lwJCFDCWTQ/qE6OrM
+PDeLcIn1bnn8WZm763uNLmJLTBFkH4d6n18pswXRTF50mymT93sHGq2HpVNDyikpV3/9hrFY+L5
QAcvmJ1N7vpgcqKIe69KMwiNLdm7n8ujLxrhiqiGdvvkMdn8G2VFJcdpCFdpC7shrSZTsXrPMuxV
Trw7vrHoQziR2ODifRuhaGP3KNnKncelTCXnc6ZF208JdY2ZJj/4lUyw7RMEbcVTSfa9MplhfW5e
nlEQlbrGp3GAdhHYk+uOuWVip9Mb7cMnVk1q1tgvz+tjQHryVG2ZECj2XsifPpimhTnSKhr8tznw
jR0WrIZHmZAf3KfsxSvm2i8s/2kI/9P6IhKUYJ9iausa54nNYbjo7KPxkglXdh5LN64x4La9+5oX
c8b8izaJzdXfVrssa4aw0kUkE0kmlzqj4H59QuQI0DhBnd0UTlK1Ex9q/vA5Uv5iq6BKV2RZizrF
gQ6WIybjNgrQ2QFhkYyK9o4KOhJnL1Av+BCx7v0j9WLpyHxRlvX9kwH9RrvxJ/eM9kA6JWG9wwvj
cfi3OgFjbRkRF7OQk3DL+ppvON/utPJtj1t8XLbCdxDPKKbmYbnxJkoWZHXb5h6WeBteZ29COsFp
n7b28Po5fmm+nFYoR6i5OkQLiCUsZYMs4sdH6LMTK78wtzKQkogxG0KX/P7A3nLoNYiyLItjIqrG
Puv8TZ1JxDZSaXhbiG497yCccPBORnTquXgnOPOO2qiXQid08flMynMBppQBeyTjVC1+uavMk39q
2qSvRHMeM+9lkOKXsyKkZjMBbg9guC2hrGhURVZFBFwgPzsE0E0vKDZslNwbe0aMvJD1yVW+5VyV
cnnGMmKDGcmAazV1Q+AnS+AMN33+49p8hkAkL7Tr1RNd8lyAFa9AMD+qsYWBXT8tIGtdpTgHzR4r
y5arOA7rb8kPrdp5mRxvOM23/Z7Jx3GrYS9FlVoGrO8P/XsTzm+M66TIoBLRyNzIf0WhDllBzk8f
3sY6Q04cYocLWJC5afd7cE967xVrPMr9sOeMvoHBKTOswhVFK0cCW9t1a/w0qMwUk5XFtMzMDlR9
sdxyMxwpo27Zm/QDReJ+JIOnEJ5OhMKMEw43xjActapHtjA0E70HVZYPIpiWEAEzjGEpWJ4vEQGh
dfQnfmHqj3J19PncyN3+/AmPR6btmIB7iUuX0pCqecMHWU65We1zUrGoMPijLqvK7t9rWuouNVvF
WzC4GIuolLnMulpjeZk3fuvFiup1z8NIdybi35TN1TP6YafAfcxNpme1XZWjgdQ8bh3sVyMn71bq
JtgJAGBTDFnc1iVwwxcJzAkekZse/nLnPKOqecrhNUpjxwU0XYqNV8qfPHA8snvqwHERDtBfhj5X
qfMD2FSzBL6Qf3JDI85oqr3ZnT9EwlFcyhplS93IJBkPTCtB6GBSEwO5xJxFji87MaNdrjZo2sYN
rGUyl0rIxWOuesjS4ZPiPj4Vn+HkhXgJ7qN1Fe7hVGJNYVOlZkV/C0psPsR+LSoqva9W7GOvk3mr
JKQ/JSw4v+4Vy1B8Y6c+lI8QlXs89aPmIaVmL7sCt+BT1ejsgC3C0dggAOUNqQ4bKYjL2A5pYsUi
IfYbRlC1AYs/mZneCqdavUd1YbkGfYViDE06r+9BGSrmfmOu6ahNJeg5fcxGkItfWuPny3ubAXaT
S38fJdBju2yJorSuV2anB5RS3L8TuLwQllOVgX/FckUHnE13BtS1cMbGaQ0Q4KE4tD/3Y4sSgFeA
9B0rtLzGy2FRZBiK5FXATKVTssLNYbB3Y4iCS1YPYrADQN2JT//b4rG78vguQHVmfnKrkfOQAUcJ
xX5rjZj7cyWjDx2P7pmFINLgEeX9c1ZGnc9bjVwedbExCF3P7k4UzcRrpp5+njAbo9JT6PbXLw+u
cKFmoboHb4lc0OpQhKDPmrdFirxcuiFzSB0UK0p7gOqV3GXJmp9MZ4Rc01MppuAdXdhXnz8ByVtE
Wp4DmSG+RKxV0aMiitmKdIziccB8j6U6zXSxynBWATYpSIrXKF3/RARtYeRpcpn6tze6H19bvs5K
DS5G1V2mGLGEZz5GKV2AZtP8GNCsYDUjDxhPFVtO7fXj9EQW7RsO2SF/0MCgSn6cw6salf1sLgBF
22vmrCEtEAdNs/FAYklsg4Q5eQoLtCfTz/2rrgiRdo7SBVjhIyM8gAKXFcWzfbWQ8n2DvmQkNJlN
HdHljxdEIPXChaHgqHyBAgMUP7OoAS0BiolNFrhWPdSyfZ9nSG2UkqsYhRGflifh06MQxkNLhFTW
WHiVod9B1qGpppxc4BU9d2evJj13RS0yROtCJJRLMfSDDjB8OhTX+rjqn79rE9ypZ+HuH0Ruxh4u
jwtWRQMWlNzH6IL5TtRiaX6RgS4DEWDVbQDVjgSgWrOsddHdVMRCN/SJPS2k0/mMot4KawFY7vYD
AqJkL2ukL94K0NP7XONfCHg2MAyVX7ZZttiCmsVPFMGL4a0iatENubcbCRzCOPRrmnQHajqF9rBc
64e5CXedcf0OrlT2Z505bsaBCTWWMMs2cT2s3G5rzxPou8gdnYLjK+b/06/O3ZIXjD7T0PFcdYj0
pR1epeK+BZOx7E3Biju+/re3SUwqA0OTEKhSGzLetjBjapqnXWJPJrMH4JtB5R2NpZYuNBbh+dBu
EoxfttFhnDZDVmok52NppICvLSjNcGDLTF2vHotj/CdIbNRM7BgsqWAuwJdZqakKTIcDJCKQtY9c
AX2r93/epWOMM+jsJN4gPwWdGN8lg7YcSGwvwFifk4rgnV2Y9SmjYMBxL9loBOY+P67ImFc1vrgS
5wqCrexBfQBdnEpBSrYFexpixrwDNdh2WuDvekdgq3xE0qGK55zN2uaECaIhcOrn3G7Fpc/oIUHY
iW2vYErqzf2wQVp5zL4p2vWta3eK1mznP06nHpQQ9f2ghV4pG89mCOBs43pRCxYri2OQy77OGGdy
+zx1btOsfa8dBmwd4HBjYi23S7Q3gKAnGkuhyefJ8cdyXeP/FUNs+V+Ygt8gOjIZ0S0ACkzlcBor
Om/aF0+XdZLQ2nPjX7X3qpRmIRauDETedcY/iEGzKKSNhBKrlmfJQpFQ825yuPXmvJEHLOsThWLT
h182gNmyPf/ieVyCK/O8YZPN6VHPfdFbRQQesFTTYGBqXjidSoJ7JzA4RFaP+Fh7B+iIFFGqafpn
MKTfWz731LM/3Lt31PfFhrylt1pUeLp60ca2Ri57YFEQLN8IUY8XHOHsm8sXExPkJbygglRdATw0
AR/2DoRc0wg+Hlfeq64cOSnRwXTJA1XsNT+lKKfegOgtvVrhaWfahrF1nN8P5JruPv2gRjJ5ZEOR
7R2sGaY9z8eCvn4XGZFzUedRD+TmXXypHq4R681FN/kD/h3hjAuVFIq0mtxDVqthy0Pr5uc2CVH8
TPyi/Eqs3PCazdpaGeurH2olBgDXsPeTCxLKKU+MTXbGySS/ujR+7oUgdMWy1nfgpObD00AoOT8k
SI+RzM3lGiDPODOgPIzW2mnlnw3zlQp0insfUXP8JY0BNpWuuY9O7bZJrlUtNeNXs4zGg0uDIM72
+V1yQyAYOT84eQjcHrEcw+VDa1kB4F7nFAGTFLx8kWiZPr/x9KaL7JFRyXMwGsT3nt4iuBamw/hQ
7I9M/EEOT4E2PBy6vf71KQk4o237RYsYbPqLz8jByXqb9mcGVBbmart9/i7cTdHQyAU4Kha+R5hF
jAdU/RBIgqu4HbQol9GJG/J7XBUVZI6OH0vz1YDVuVLhtCKXE+nIVjwgqvBSerP4QwvDFFxk0/YS
vr45zpVy0Bm/OIouJI5rKKs+7pgvyw0pyp9Euw+Qh271Nx9QsdW19EYUznDWvNxXOs4wiDkFynYH
rGOiR1nnLZzpIxOejLDS+xsT/WJrECV/+Jhckcp9Lh+94KJzpxlo2+LWfbakrrb8LcGsMs9bxocv
sd7nw2lOyPwTci2mgtVOi1e95xuWGK39npHsRw4kSkQPbk3O6Z+/9fpyAbDWnvaj0iimbI1RjVIl
jzWJZAJMWuZOGD0yaA7mp0cJ4eNaT6OZ3xF8xduyEe5lXdi/IP5WDIyRlkkuVxP3aTonA5BROZYx
00/crO0phQ4vteqXFeAESx/jRYcaHmajI9RW3L5P9gvZlkY8D5gifYyHPVK7jVBGDmLiIpBQqM9F
NjsJm8dKTfO4mYN7Mb6aymeGgHNTye1/XYtprY0jGbPttYDa0bMkuiIjZAIXdOmY1fogk2ZHnZda
Lb4b3lT3uPKLXWlnoXecpaRIrgbFgFmumU4B7w+QLfZt7h0LiQHxvk9oReV3LdEH4bar3yr3tVEr
5hA18P3TwkJqduR4IdDduQ0MOAVoiUQEFpo7wcDiAPKGa7xJ0LvIgQRKls4qQR/PINdAik/84b3E
MZ/X9BDesLvR0i/ivCM9Bvc3LkQAQn3BuLYcX/Qo5suzQGnx1vliVe6A70Mi6jXKXO16I3Y3syp8
z+2e5ysWYU+5OBTjBI3IrNj5PR5LeIa6wZ8e+9U1nyvcR3Xe80kPhRDTBICw7ePztET4dSV9mrDx
vY3y9WFQoPbrfr6hPagMe9CkUMf6CXW8DTVo5eglTRxU2RGUCjaC0GFaVxiuoPUJ2QcHEgJK3den
P7dyiTi2/TlQsSNLc3zZmvWzmEm/XokfYnCFa5ylJg3QHuCnqcCVXqrOyf33oOlbB9K41WWJX54P
DiIGVvByXViMba9MVpY5h/JbnteLpuoxw0w60y1L0yU8dGvtRQ0zpWioB8kGF+cp0rONnOqq9jZD
bAnkmBIxDSrUj2U9NTg2pPAzz1Ov2VdU5v+sLuDShb46r5XM7nv+lEolIQqgSQlTdGcx1QKTMPIm
qiAGh7niPyJ8Qr2Ez2rVukW0Jsv8bU1t1e1wEivq/36MjO4L0B7XLDyDePBLYchGZZ5qSyOwN8CW
QmO6OGDIeqkuNmzGD4triZTW4Wqfv5Z8FvoUMpG8Tt79Dxvj6tBx73A6/wx/kBpptk93BXWlHQ0s
4wjDEy9o50evvcJf0btF+Kz30sB3THVkHhhVAwbVNT4HppoVJ32jWrOITwqL2ZdKie9XZRJcP209
8FInh3vGbssVJiacgM/IVsMUa6wocWZXN95CRsIO1GJbb+kJgR3X6mdBnySqp8zU8k6ic4kzLYS4
fRd7e2a9E/CHlCdtVFdrT2H0w9KeW52nAqqhNEoLstwaWxQ8wCPQ2MAIgU/5gCkRh9nux8vlqMd0
FSXlL51OcvZJQJyiXqeVzMNI9tB7NYWn2IMqkh6FlHjoy62qAcegp1henQxaEF3F6265BOO+Fcid
ursF71K6HvabtsTCpgvOknC6bAPvWkZgyC0Jv3fsxXujm7p21uxLqXSMSG77RtBnuo6SaGOhUAD6
89MbjEghJncqVkFCZbmfrVEKY9SmI6nx4rcR4j3hZ8Ro0ol4R3j1pEaD8ObZTHYkJIMCGOBzGbJh
On9lkq4WocWlyQuS1uUo6ifZjMP6VBd90nNrozOxbAL5hpmunBSy6TLEa5Bk4r2vZtHrue/hY+og
HmGWPazasGYBwikNxayqBCXtCk81lhk4cgcr8HTS43p++MgbsFDidb6DG+IPDHrEY7BcKnuq8XSF
eA0znXXkHN7j8tJRqwT+BRWKeKjIJ9Y+kaYak+zC2uyOW2/Ej9uwKbBVoiklNsgxin8YLSrxPKE8
DqNC7bdel0dIMHu1MFwo+Pnr/qEBkKiDhT+avDkufli8Koew5wA/E7DZnqNcLo9UCULArVa8/bQK
jflREmPM+xkNC7IES3byRPSK0s5eDtN89694ivLHs7zpRB3q3w+9eEbogNMDbuCtYoQO5uOSKcjt
GONpY23XYtqrJRvFDXMAGg1BtlFczBBHNAHkEmmgdq3aGvX7YOaN3O4tq4mVkGqKM+CguRaI5NvR
qXLPXMnjeTw9zWu4IIwQaZ1WaCrcj36Y75OiG4+eWmItfrC09y+NslNYs7pcwHRJs+T9WjZH1pqP
b6sqSZWsz+/1q+Z78ZcdeqA8X/OETT1+9QjRUmi/kS0zG0+D72jLDk7yQ3BExPM0oNVCxr23Rdgi
kJwzv0Qeeqkc0Lr3AWoTgcl0fOT9RrTrjofIB/05w+LRiRBsB3bS8yygQWaGtF3rqEY1SOdozm42
IIpoUZYNKLkZuvrdCGMGqX9T/0uUWyaS+nl54EBtsAlcmaJkbcTmDH381myQc6lat6foznS5q7qO
Xm9uvq8kL2jAFMjFQbIxhpmXvQMIsLq4KBKrOtHVqCu5E3uEWzGNTF85qeQ5SZwO35n/XRiIVzIK
B2SF9hGSuL3RNVnqiQIrVuK+Rx33o32d7SxgMeaUsojooNBDAoqL7/WTAiXJODRK5GK58Hf1BY+C
Dc1Xcsh6PfKWJ4J+QBQsLaXv5z4eu48/3Rgrv7sk3e8I6WP3McNpfT5E/kxESWT7e9S389h2rEds
NUeQzG10TTMgjgoKMIRuiiEOFRXMSiG13/EF8LfyBS3A3b61PN388rsUT5NcR9C8msLjl4L+l7/a
/hOYAlNBBM1MuKplEx12PKq5yv78qj3MFw4Z4GjlJY54FfdTf+Nk7H4xd4g+U5vAtsQ5uJwKH79D
j0jam9nEV/0qVu+v249NqEouxx/+mdQkRo8WP8tiRl0J+bUj9k48FVZuZo1GYjB6/5el5HWGEYLs
JNyjbQM9TlRc8Pms6gMbjYkqiQP4SOCMibKc+pWjZcTqC6tB559r5dCQl1O3jcJFVz43ApkFHmJR
X/6DTBsaQcqFkBM1/R9s4LCL/41nMtjTAiPbSasKE2A0TpvaFtahDQAOInOeif4869t5vo+lx6V1
hRO1xTIHrx9RO3OuE+JAoacDVFUvKpzLwH+IN1IswLeVOS8tFWMPnr/QJZI40/OZWWAFN1NZ+EL+
gfMawqbmQUOmpXtGtOA9JMqnsDhhxI5m3rwdW3hlEma/F2oGJJw9hbiWiwe4u1ofGUjVEYPpJg8r
axqOsu7bqIOt3Ltx8KFA0WEjfHw5YCtoo0xYoJDu43bIYxbuYjA2rN8THpGEvswGXF3W12PNCd9z
MZ02J2qc/u5ya+SvEK4CFAwCVQI4VeppLUGk821/zNhdH7fKWR7M1QKUP/exundaqUqAf9Kt+xfd
rAJucGf8S9vAymkBDSMFsnsaV7ZznEtz3/0yNLgTZ5qSDT0XgAABikCymDMzmUkX53Ls76L/wK7E
x8CxdgdX6y3O+2ccNYdLymMCBgoiKZJo+d7A1duQq2A2KgIGfP8oavn77jvk0zpB3Ihi5mCVWTjx
E/rCUwl4yAVUJznmSczeLSFrk2tPyhBW3lBmr/H13Z/xfaY3t/95txfWMiJ7rO3ry87vmZw3Fjk1
tZ5JGhCAYuthvR7AXgUgGlTZys2wEBO8AZ9v7/2FD0UCPgHChSmnVWJGXuK9s58MoM7ZfCHzQH5G
Yh56J4Pe5HjeQiDBJTq6LHSRgtpyqqDCArr74EXxlxQpIuNZzu+BW+0VCqVau+z61qiY7Mbyfeho
ZW1/lorIVm4CDW2FV/com3+oyT7BALvT8kBZ8HHsEO/TZAwkDdN6Subkug1okOXfXTX89SSVh4Pp
CtwNxLEYKLSz/Bz9tjjyyYSlPcsIkbjqtEuEWw1cfr9Ho0Vca2ryfbeX7qhifNH+hw3IUAIqpj1x
cbJT8kL9pQSmAyD9CwKi1vKTZDUPUmksrkSAfgLkeRCSg0ueni6tdax7VS4Xr2gTDyH0G6SJSyPg
TQwpTU9xHFwsUVt7ucMlwe4u3I38YVqJBvIr6qr0pv9j5HDI6b+2bvebX4tSuMLnQS96vJMcp37i
HJtejUo7T6lP+32g4bsXMhLwy//raYiToLwHrJLcBnJDLkkIGS+7DKubfo7I8vlgHgIniE5Mk7zC
FtmrRM8ZClFQrn0KoncwwjCmsTjkgd9MCF1wyxy81zPwGMh1a2JFOH/SlHnFPTznRGB6nRgjKOEN
txKNFcaFELAo33SSujgDkIPhasAL0roTpbbZe+BpwU3tl1wJSi+j92JP5wBjMJjdhgSAUFukAKQq
C9uCNcfioaFdY+NWAMwnlvW+4e60w3umXyiY/MWWAH9sJ7e4atQAMGX4sP617J0NMrvVmSOth3aW
33S3prj0b2XsS5JTl1UV1WYhrumNWhgmV6v/1/McBmcQ+manyCwNo2t2RbNLNE+Zahi9g/MUlw+g
gP64xCWZzvL1NNoT9QrqgzeQMbwkegR1Tb9t0pvXFVL7HHRfGjWWn/58DVDfmi+VJXbefNXRjsx/
+X5Xw9j12MhMFnqWKiMG/t2QMmjM2xAQbVl7KaCDtni+GjTkbutyBBMBKRumhTv4aCHKTCJNXOqb
pxYi0HKID5AgymdeYNXGy2QgCSmLrXC6ylj6bRXy9qpjgYo2AZuAvtpOIWV7zu1MShaiRCf4EhBx
M/CKzhSJirKCTRHnk+NmltHjKFD2z3attAfvDNnAs4M4enMg0SHMKUnOpkbWniwU2cyjZv8kqxhS
mLf2FzJB2Xjo2LPso+PZMP8dXqjpmM9qqHxhKrnO4AXagteIp6GkUD3+YtPfXpbQEECk3ehqtpm0
uFztJenOHhGO5rxg7DRQPC95kkZAk/lHMF8vlmnuKAKEaTUNn8UxMJMJjyPaVHism0uIq9zgEods
o1DFzBn4Gmal+FS8iK0lZJvFlvbv8g44W75Z/fpd9dnEvB72FF96K6O8cvaLtfd8F14NtnVYTal8
S78+UhxWzvMhfJ4clHtCs0LJ/Gu/UIJKcfdK/FOgienlbTzixyp/rr6zBqP/0sySMmME89FK24wX
F7abGm7JmuPj1fMRCB555nKhbXT+TKvX2Ah8jo0sCmTbUVBZ/bEuXzanMcJogqjFGqk84Nw6GfzR
b2e3kigqqdE67TQvL6cpY/NQXzlpA9/GusEkTjcwP6ZUpqioCmBLS2XuXlXLprH3bhoNggSY/Ybx
Ol8e6ncYy3zu8vFccZjWldFTw0e7wvDq8zf6U+rKx6T9dMRM6xFWZvC3/9C8B81ymjHLy7BhS/sB
+bU7okLZQAlDsJ4Wpmuv69nwOMW4wqrqf8IE6mAd9sv+jBSTTaGu9ot+X9TkHAqvM8eKJlPji9dz
fh3Qyu8+PTM9XtmIJq8AcWFJ7MSqAWpj95QLFeiUTNql9sXBhUSJEowUletPjmscgGFVe0wJAAHD
NCJ7/y/XQqoNvZl++fd9jI2Tep5V2csv5j1GSiSkDP9l6KUpg2FWlCZ3a41SPjCySUaq/YexZ9US
Qk/qy5DENlgzGb55007fB4dwjRAuEUwjxlerkFb4MIe+SPNQtz0013BEToZ8iY5rMU6Se6kDbBT5
mCMUtFIKB+UwCkuDHx1UyoyLEcmEdr1DBn2OYMPyl0OOXXRkSRJgxfiflXqVy/kJOS0H6DObCuKs
uAxaS1HGecNhpoRlDw6tOQXaphEWh45aslQxzdY6SvuX9VEmUgONPQqYBoRZfwfAshw8AGVEaYRK
pUUGWlcb3XCuHvtLn4AAOFnFAGmVoACxhkHCG6wVCUrqU6GSdNVAsQw4pP4vewL4aGxbF6fIyl+8
XJKPXU6y2rNAvXCx+Fm65vV3axVRQfm7IuMKVznWoVi6EW8uILfowYk1O/F4YjsZUjtbCV1haM+x
U1UKab3MnbP4iE8zOSARjENAbnn8OZTye5eb+YK9hVD2Vd08/PZbSUZEr4J2Bze+fl7toYtYSebf
/8Oe8AZRE/kzBTBv72Pi6eV8U7LyovB9V/1fP+Qn5D/FvHs/yjywnjNuuJ2t9Oubrg6p0X2N1RDT
9wfO6ukYANLM0Q3SQDus55AUfxoqXTPWqwOUTPoegX/lL8d2HAoutkZuz29b1e2PXM1YleaE8HW8
Pc4gLSQILqpoHGpTDYgiMtrdfeyY/uCcYgFfbtwEGs5FKatbrPkHvx74VhPmK4se+rXpKwmz5F95
4y8dGUlW8CfkMaXWiDl3k3W05+7FRM62/du/4xEx71Xcv+6IHCeJXIryciaGcGQfz3vm30cxOgBr
khsaF6d1CZc7jDT5ZxGcged3rpoHm0n1L+FyZfEunCRCk5wDfIDIfhKF69+P8Co8IYR7De7DYzSF
elIkZ/kfo01ZINnPh4nLEPctMJH/LMSbO1115Oh96YPaF19R6R0VhjXla889ZRfYtbdCRgRZePPP
R7J0eQl0jyvflUkuab0qI5y+7SqPHkcsHvSsMKnxZEulbAMseTBpKozBmp+/jqDkZoW8FaPcytzq
kZdGMhea9bDKsva94T1eo5nYV/ozNCcJfugN+11SNNY37TRj2FBDNIEBnaDmIiulyyW2s/9nUOBo
Zca3acNfcpiEQzfrK/whlHMXKb4Rx9xH0zUVsBYBmwtyZ23uH/r0y0EfNPv3Pk+yLJ3sODCv796q
zZJhAZCRYxrnRT6h84Bw2NYbR9ik1XjRyO21H/OTIC95MIbPggpQGAXLgtZkr2UG6WkeKVTsJPEk
F7mCPXSQSDt9s7vFH+dbQagYEU+V/eocqmfcYdc9yovCrI5O4l8GwbWnl6zq9O426UNbpdDvw/cE
7G3JYMDbWtNdBaQdtN/osF9sdvdAkiaufBdRL3hWRLr5G98OtBWhs7+IaeCYzLR4ucaUKyfn13HI
tRGIa/V5JGWsdyKpYN9guvf3wZiNZcFY1/JUUAQU16JPL69Oc6ReAtbmbDsvmU1fb2jVLK5R/mJA
n/d+NG6Eds79p1OLll3FT28yHq6J9moe88Nfn5rSV/IU0hf75c4VER5VijxrhOAO6jVJ7CJcwLTm
mP4IBbe2Lj1tUhKE8bPGlW5YQYKFPoOb73SV4g/0S06zcynbx6Rm1ijxKN50LHURy1FJ1Ugk5ekh
71cAKOAcVWgGYI3yUdiTTnnx1dU5h+H97VzdIvZi2utdo4qIB6P+MqbUehrQ/JmLwvlyN2LrQ28P
+OhcqUsNT6wnY6Y2fnavHB9QuXMuuC9j861994LOy4f8DKqaZC/G2A6m5KgkC0hc8jcjmrTn6R3T
j8Joha7d4pjo98AfiSS0+P6vwHX2G29T7sNFIqU/du14SXZYqpLwPWEgKL3FvnAcG38FouJndHkD
jevDy5lLQ0VXhVI7jGJa2tH8uaIN6Y0N3Vfu62QUetAUqO6QvBxiV1uVZgozDTQNL3Lz29zut64r
cAzFravLMFWBjh3e6H30jiVk9aZ8RhpH48raJbIO2/fuzajo90oR/U/eQu3Yx3PaTYlivOQjtpYe
sFQjvUZy72ADiYMjxGt42YE1XCdWNGQ7htygOM0+cs74+vb61pDT59JWFbPPFVCMrXMFP7opv4kZ
NRL9YH1Jd9HdFOT8VaNr1O8B02vag1qcz5TAkv3GG9fSKmm9XMGbRoHhn/8t03dbgshZJu5JOavi
x9H7kCZK5rot1Yr7u7rFBVyY0e4GN8Sk2VEDPLd2Pt6sy36Q1R+grls9FmBWR1LudGOFcijKqRpA
/LehM2q/NmaneCFR6AVo1FuwrUFN0TxXaVQWslTf9htTSFktz2FqVSNFi8Pl6qF+lbAIf7kChje0
fpzLXoo2AcKZ0/jWwEYUXpD6UEDucvy/6FviWHrNvfG/b9Y5YCLmX+WYeKs6BacKCi+HbUjzz6GY
QuOUpR6uxkdKyCvcultItBIDwaMl5fblYodVy7HE9cp0jkam5Cydpq4CXzt10YbaYQOzJYYQ+F0r
+UidPJfySibyH2zSkVeLJZGzS4qoCuV6gxYxtAQ0cjuoE9r1Dei227JoaEFphFF9bVq53l2cbBHT
B/IZ5RoxypfdQW8WPJosISZgDS3YLxq2K9gNBZ98TEWWlpZqu2QuC/bFsf+bKj0ChwtDo0z1iS4O
KQfLFdp+F/SMb1p+fNqViODnJgo8/kNaGkolj+2yiAaXdKdgHg6Ro6I0ZFcxNNNECaTzdrXgum/t
9ykZ9hw5NSggHZC0yj0pWF4RdyXM06FDtCkjFG6nC9024Iavp2oXgCuVaPbRjvp9+xoEd17bJmT3
e4xbcoWuAfk5KKwADB4Rz6V59T80Hs+jV8Qi6gb36uPHVVSRrtoF3nj3cDnkKL97MENWhj7TzI/4
Wz0w6QzhsBf8s33AN0OFtxU2vB38UNQtMWDi6R7M1CxV7VrC/CWptOP/FopvA4S4ToSaz40Dmfog
KLr/joV03ZM0VItftueLtEGErToggoqYYt1ry6wZICVH2jKBmTOCIYnFckoCBTZjwveTXZtUFZ7a
LwHs3/+1gauB+Inu5ejY9L7kG4YX2GPcT+02ulXsNe8n1d3M6DYI4TGDU6t70T8vJqYHkEmUeJTM
s3wHd/29G7kbaIH90XpuTGFTXH0nqWos+RxHGUW6PSmT1hfXNi8OV1QjHwwcyA6UxsFSnjsIcVhP
flqPwWw8MAGH/VA8LRvJ54QCzkq+0z6U1u6dv6Jjs+/JgaU34iEjTJMrC30LRB35uffilAGfEQMK
b/ZapqgXjHLrBkzDD3IjqJpfk/OUBEqGqzX/2JU1I6WGPBeGK7T17NT0L9elqnCmmainZRBQeaa2
jUD80A5RgxxksMJ3FAorct1JmhZWl+3NaoRpjUJkEJIUZcnNlQV8zYslhimkdeZTBQAlLEw3FF/h
xxYsVt0rDS5dOUD7qDI4AuTgtDgqQYkBBtm8khvEhL4NjTf5/CUBQzKl6JW00rZznoxcBia01Swi
YTi9rwk/rWPbx7LOjloSJbOjjjYPQwa1BhwGu0lS3HI+PwCknfSU00L9gBf5Ow4LCN61lm/mZHhr
9sGeheLP8LGeTUHW4VNVxmV/5Hb4n3e23WIiKotXkNHnYcdXe0yNzRjSYvkCTD/zoaPHhtfNR5GT
mtGesex1ROgCyFdCxvP1oZa78/+SHP6rAGojazO4C325kR/Z1HBCLU337UJ3lTrnSGFtM7C3wOEJ
UtcIrkKoC77Yb69clIzVEh904S86rOmPfOADHo4HymCvURXnRW7ezONP6Zag7idaZkx462/RAFfr
mqPKWpUPB/nr6J1F13YZVFHuUPNd9+z5GjIsJG8CplZqc7kgD2ckBGRLCJqdnRk4r2b6x9IP3BQe
f2kMZm5MGdgOirl/cG4Kkb03CLqYsZkq8gTqg2LZ4yTLngXsYuJnaizHy+zOUO95SKPuWBtLH5RE
uFgO2csL/3TZwUGKhGtAERQgGfFOreVbQoux9GZqrdQXzrIFB/R4mubLfSxZw548zFOHS+HQKm2z
Gi9Eb3bWntGNX2c7+o/ZATZrifplXIw5rDEujeF0IUebqiXEtlVLS0Q2JjPBps2cLemn39NeSHFk
d09M2XVH6/olz0zYTtK438+goRB5vcOM0Ghpii69p21d0L0jax8YNpLVLZktTWnqePNUZkpmAeX+
T5LssM9NmXD6QFbmKRoVvWY7KHzwS9Gy/K6JNvmcG1qav11ZOS9qTdgrr8rTWh2Zl0Xs4XpKfu4n
+PK3yT7kvjuGkXkM++sqQIZiNhyECL6nQbLFAvsejXphly//ruK04VC3x63pQsKiYGN4HkVfUMs+
7GBwVgcqLW/swRa7lBwBSRQcomUodaPaZ6MA2LYRQ4PB2Z1Iqiu5dWH/W+G3sIC1LxUpqR+WLhm9
FHnM0XkMJXxgLNFtXcgRKDF06CHme0snITqq71CoMQstTE58510EyXhBu8Xr2vVML2g7LeepNw8X
GCfyAk+UBxNz2Ng1rO4WxJlOiRN0kWVd3vQwawh3IJLSJguK1fWli2u7nffa6hb2dHTL5EacHC1z
YxkNhm3QpdNG0WS1kpAFM0WSXChQSN+nu2EXvxe999Q3oHHGNjILRnWiV/Ae05/kkGQ8eHRG/P7w
KpcKjnGbPqfFS9BZUixxAUrpIB+G+fvm2oVeEZyQ0p/HfS3df39TWCQmKXVyFCY5tR5vFpr3rczT
SFHf9X92rxgmT42GvJCkjiaFozduCQSUeYLrwoie0GjmS4NtQRRSMMiBPnCz8juzE1PS/3F/WByQ
z8CaVDoP++vr95+Cb5u8HK3suEYTma5AIxKyLuCkdHM/EiAH1O6foXvdx6MkSX9bzsATrCMjGe22
Ty2XcQB1oiCgsEY4sFrxYYPiDFSqFluyhJMxJ4o2IguO0W0uRtdcI37uwlUnyT0GkQizTHTfmp2u
nPYjt0vtZG2mKsOR80KmX5uaeujJP0vl3oCDyL1RLNGxCctxOS0XUU3QP5hyk+9/9/2qdUGHnxGN
PwNTcIKnMtWXlDeNWtNoTe0VOdWtF5b/JnKOQ/WSqFQuZuGCa6Ysad5uGkg/BAT76juiyvXPY6OA
tx3LpdzOrEV4QvmQq7wDYNuLLv7IljD8hYDriKBc5Ur5D5okN2Yk97BLDwajiUkqi4H+fJbaDjc7
j5yCqKrLOysUkY6l02YTWn2BcDFlGZzwYeWslR7hV3wPqm+Q5WDv5CN+fHMP/tdz4G7VdscI7qf8
QcNQfgJjTqZKsdbQNLjGtwc7JYpHBUWgbbvXWeV2vzc1lAdFs8P3qq4mODGth0AyWz184FFXCl5g
3w7Amn6EDY11EFeiEn4S7AXTwwQWkDF1kO2rKEqHzlx8ZxJYcMrndFYd52PqYHDd9iYpM7T6y62o
fXZ3mHKF3SqH0eXK82QqR7Zox4pPppFBf5M4a2ECg9LDMsA1MIIBAyy1Ae2/mmQzMHgzRtdx+4pg
q1Ucjcu6feJ+u4d2ebRWcrfaJ9t0KWulkCnSFU5NJ4jNQWI1VgySvaDi+5aj24KapR/6gxwi7jUq
z6TRA4SCJPBHbH32EiJ8abgYY17z+hOT6Qj3ZDhhKL+p186fGzmczYBekzEHO+PIFRP5j8GrF0MQ
9WgYL/JU7dN7EgHgEPfB1AXQktEuBPrT4xNIUMSKyvnYoukgDzXJAFZG1swSaPEx0nybvZtw5I9a
Mqt0/uZcpTGQnEGvraBPSK1OcubzRqNHlKlQRnQUBPwUI09E1+ALsNB/YDY4mOTvWPVZCyiB5gp7
BUB9XEq2d9kixAkA86kYrCtxJqE56QYflmGH/+lGSMnQrebfDBfAENY6EQLMfEIOFYSXlL1aDvPg
W3FXnYSe3w7Tj/fHcC1xji/dmS3rrLZ052fnZHlHTrkUfV/9MXOO1zecjPbhUBaFK0h8c1L9SLJR
G/yNfE+GV5HgoazM5QVwXRLVvfQZbmFVhEpTGFS+N4/w+cQ+GvDfnpQDu8ExJts+pb7TsCxcPmTy
Vl5vzEPFdrWXS4On7O0DWIapTQSZoNQ8TCkeTL/hLPL4vNnfa741JGMjhL2TW0ihhpsXB+63bIui
pc7Sg3F+YhOd+ophDcS1deHMTLbCXWLw+hAS4+c7ljg/i/rY+wxREqp1hqBBrJrYrddSbTx0G0iQ
5AFKAI4xlnICtFSxOdGsf5hWjQP37leDElyRqZXE1DPOTKOHdkvHok+nf/YZSyVDiTAWK1WGScuX
FrXpilYT5Pp6GziPOL4fGhn/DSVzR2ETqif4IK74Js48VfrY5kYnRHnfKXCZyP7xjc6h/o5vOH4C
ToGvKRH5K47Xp1OH0tM34vWLgQCHMPIn21Qw9jhTCh+GTELIsFcCNfZMyeds5u3sxI2otJGE7g+F
1xsEi/lfxtcZSreFftVDuhj0790vSMoem652USiKkDxGVgVBBX7IO4Q02ngKDMPVc4IzVBxftP9d
rx3KLRrjSi7R/v3r67FgLwkiO+iYOezzIBVNp41A5ayOAHb6BkQYB38d3Ut3hN4CO/DQJbl3Dx49
RP0QvkOMacdtmpMnhEeh9SClpuVK2RO2Bqvrjw33gyxVRW9bvoEEMdwrOEvhnhNfrZQuHB+dZMWF
CXqn7hRStBGQPWX1HAN6DnD0fGsW9EXoJFaK5bYuhni0S4e7Wy3Fm7NFfKAZYnspjwuZpK1if+Vn
TvEA0ENaXXppK2IjtdABfsUvmvbYRNogmRvSqWeRgJQjJsDms8AYXkmvqMtG5WKiaMtZo7z6G9Dm
1KlgbJypI0Wruplq+K4iYXlH8dWHhy+b5nUixBPSmSZ+KelLihqN8yJQ1jma4TG1O3g+Mk/Wi6XU
sReCfsL+guhYGH7zooVlYyuJgHDWsIyJ/EWI0ryUi6u5flS3uL/lePBAK0wFBicUZ8FjAwO9syPh
TXrEiqmZdN4CNS3zw6FjW+ipVYMw2b3l0xnntI3Jgzr2GdPFzLhsN6SgOlvwcszuCBx/3jfJ5oOO
7zoerd9a/CMBfFsNTmyp+wtKw/2N4IKJxVHX+7wgfxGn8OyWqrbAr+FPFjscySMovtL6vLsidxJA
3Ys6wssoOBl9IBwJf4/GW6trmH3gzC4hzgNA5m9YYQSJj5nPY6zx4HKiO+Bt4ctesETh5Qd5RmNz
tfCvlt929FRvUtac7nH2oR2NX8pXFEQllnHrm+TpV27UdMh+ba+OGCF5iTyNZNeqQtnW9kMmO1TJ
w/1gAt7MkMkF/2A3FmXW69QuK5GVjwtTS88/6z9nYEpon+XoL0JwJIrvzE+GSb0qPvT8T9Cq1Nlk
GXZ9PgY+Yz8qJRQ2Vg8WASEpIJ+oAWfmntEeCddmAKgFYUXE5vBWho9A3i2fOt25eF4S5am99W4t
dsjnqMeHqs56T6w4copWbxFaStv7u6gJgG6PbpPBropFOQTzpaQXKnCRzOonWRgMEQXcV64xKHqZ
ht6h5H088i3ShsQGOno3KXT2gtAyunZQ0H1EzSJDVS0ZcirhY6J7q3WLwyJ4oUcI3LOlrPPmKl0W
U4w3SFsN1BPQ4bsx/Pj+aMhyDo8Lz1ZfOV8as44BwFFtxwuU2AXD1M7xUS4Kc4SylbvevuUe6SHD
Ksiu+el5eqyMZs0NOpje+mxt/u8eLtEhtUcn6neS1aGW8YoxTq9JAgFzCboi39y5xZ+2xj1HIgA/
5mvgpx6fx/NPfkTFwVSZHzyt1KLCF+hv1gVJZlQitBWH7+vdFtIdKwfbC9zBkGq/xG80YDJMeEtW
lB9lbktFf7qKTLcCA+LTmrPmMU90dwt/sJZY+3qQlF8kJF45qjbfxjJ/E/15XWh22pCucVgjF4HV
S607CinYeC3YcSbJZCAYwPgQr461/02zCiIkQluvkToW/RqH8vUwWlilSTFNniQKbIsR/bDwmgPJ
Jf8O1NgPUoAL1k5IyMFs7t72WC9YFNzUynPy8FU8sfRYp0f+5GkRT/Xuh7JN0ITZ8OxXMwK1LGeY
+Kt/rg3FIzrJWD2h2f11fm+4ap1Kpmtmz7z67E6sjIWdfq5GEWj+ZYfaHxHCTOWkNE0wx8xOO7h5
qqbsUhjz0gqwOhH8cXmakS3uIZxmhCBZYo26hNSgF9xmR9IAzd/oRker33S1r/A6YkZEZUz6uqgN
HxMijxqjtL9bHuQf8zWaFe9MJcji7emTFQZA/Q5OyMx1VYxRFYEfyXj3Eb49taNG3AyWjeNjpSv+
tNe144ykBtIuGPWVnLiqyujhrlKna3MbT2GW3kKow3xlDkr3M2TjrQS2YFOW8Hg+jbZhXmCKdc3a
U+dvEB21WXJtPOEveex0rCM7rzIuOwL6r3llWr3U+7pgKRGGGNO5UIZ2ceSFea+PliBf1Ifn0OCD
LGaaShJZSFA8VKHbNDbQ6ZOsde14KJ2ih5O1fAo4/I6w/F/+qi/ARR83glgSgS4RVCFeb6ic13cY
DjqIscpVcW9JNgCzjwrcES0NV40bemRIeAkyREhSRgJaSNsKHroIF6ga33fX946joNB06oFEEiWe
KR7VZCw5xM0Ko43bHnqNpmlIGlFjAuYXYwA1kx/9DYFCe50V3pJBF90OOQyAnHpcd6HUgVCYpS4G
XB1l3wjsxCTIeQL3wypeewTRi2f8Rj58YaY4PYKJ7Zwie9+KCLWRReySCmU7B0O6s5N3rkm7zp/d
WV4oZnJcPyjmQqhoWbT7UePfD6noM+LYnT8oYx6QDBk1EYCTNEa6eSgZX+8Woijn2eLDru0vJiId
EgoXwFeeoPr5aEGBohASdKs+OEmsAePl7L/EIIVbbWkta+voMliWFCLqX2cG7Nge4Mo8NkOC4Fee
Y6ZS8onGupIhxCmTU2ASxEv6Rp+wsxJ2DJwfCOsuURhdceBwPWf8QY/plXwV15BY91YsDFzQXwzA
OEfovXUxhhkAREmeUn97Yp+wsg8yd7wKJF5SlxmEYBOQxHBYFRFbHlC6ZB5p/L1Mc96lROr4odwf
Kar/Hp7PnoX/JOWg2RsnmAUb7A/+SHyF119Trqack31Ju79/R1cROuyn43oETnb9hKTZ8Q2H/W7P
qkYw4g3j+7qOOMRBjAA6To0I7/qXQ5bB4GgTVQsuyi5llzECWJ7/6iYiAu8G/TM7mbhLNbl1JKo4
JbbhdaFWFOjpo2dUolub2maRCF6AlQxdKbvaLEvXyDOWrRaBTNLZkvYMApn1+3AeqysA9BIZgUTD
3bej06nwUzdfrluYLrjzn1AFTm2lnuaSkMB39smS0FbuEATYRAE2yQetN+fNDV4LFwejwOZIiJBi
sYNJVfarC6mQe44F/ShG+lxWoASuXnSdA1jhy4bfJSGW6/PGRPASKiAHOnBpIVU6BZEDPfzwP8uj
x3FUSnh6NV31u2BgHx+6Mg6kELi09LZlO2SNQfR5BYVzcI5pSG9ec+uMf4kJT9EhEs9vqwHKNKGd
qYY3EMDAOAK2DkA36eMruRaKnr7s4f3qUyVW49yfubF9rCdp0nb6csn1ZdcK1Memy6pdaviTs+6k
LcqqhtuR4MlmvGiH4xWH/kylIPTNbNJLJmLvPyWHRLy77t/RVfWlGCjchbeN7SKlUjKn5x/kcveN
pZ401vKiiVZLXX3r4br3la73Qa/9bxO7sQCmlEvFNEfSurDmiZhm+7B44YpP4iZiF7YK1/EgxxOh
SPwRevwdst4Y4eleuPKY8GPNwgKEMl/XogiUBaz1PNztMW+/0AuigHlX5HWsNaatPX5zjkRv3Zhy
drrcFb50/Q3S/Hi0TG2K/pQPw1CAvP5LH145wYiEyWJv6C4SzrOrOjhJGOH8qCWS0z2AuZALrhv2
6TiwbafBAfitKAw1gFo2Xw2wt5TVYlLetc2zjW/65cNeCkhxUeopITxVDUzhEgWZwpT+OhzNm7BP
P3XQCcKnqTmv27p82ESUOoCQiCjOXWo79c62i1YSlhbNOyg4hZnP2aVulGS1JeuYMDfeVo4RzvEL
jG/IU9+Si40J8+d62TyJoSE7Y690iglOnsJKffsULiKRuiRy/gsX2JSztvV8rsIGGPQUgYU+W0Ee
SgsfXo9fgHElPuNuyrokd7R7qg5P71rL5z7FuS+pBzAraYJXu8O7imhitfeAlmXzytBhxDrmxzSg
VAyzhG2zdJA+GR72EK9BEXWWlWhy1Hruc18u7ew79lIJsBe0cUD3OtlbGcWJvib3IyDX11v44hCB
ItqgCtOJnC3a63zZloZH8rIjtPBW1ruLkuSiAsMzS28o/pCXx7VbwrdZcy4nvSY9qTNmt5UR/6uf
SH5bsIEGEArOAxnaQ2QvVuzmfCFr+HKl6CtOROJ3OGrJydwGFcsCL82PkGDPPTrMThnJIYbNO6J0
2SwkRu2PeZuAxCd88Tq5Kmgfq4b7K+f9sWrxcWa+jSI3rczBsB5fyAtaAXJI7q2bnNIjuEQ7uhL9
S9/9vIxlRULz6cY2nVGzjh2ETqPQzNaWCuFFacnda7UBmBCyelSfNO0t65CJUdkobgwmRt7TMHFt
ufCj2PNkVCUU+CzcQYLF/TwQn26NCO/0uQGg/Uts0pPeR2P8ISjNNZ2F1Oev/bRWXG0wNR1hXsjT
0zJFbBATVT72gpGUrUWJ7PUYUCr3hDyY6PeGrsr8oAmH+fsYlkHzXQO1f/+qKEtyMvzdKyHByB85
WLNZ7+p7kO3y/yLqPFWgsbgy87Erf/+dRK8H/HakGDMu5+PwgX7JApNu2UPu+ZCdnIIcCQLtk9pe
mQAHlnYKK0Ko3sHL00HnLcnpocERKjVBWUcU7ejB1a8qs/5LgZhgCpKEusZTcmSfTDcm+WHBZDhq
cx/Ru2EK4IgZlyPiundOqxiYSSobm0fbfrL9tSnm79UTkez/YymSn1k20kCA35WoLPk3B9AhFxUD
QoZBJoFXFlSvRFIKvCo9dRoBH7EmfLp95AiqU3yt7PbAjM9A5dU7fUkmMjL/O9NOy57amquX3fU2
I3nkRSpsvUUf8XskmuSDn4QH2xqXuEVka+qaSRMydcmr9ytgyLbKuiejwephqSrlk2yixlYJsjIH
pt4XTyIKTUjpBN//w2vO6P8QsjUnWcWbhuFgj3VTWE77B0AWxET+cTGes8YwbUzEKkACFKn0hlSn
i6G2p6I3nCNh2cEjZV3fXcn5xep7lx1DMzNMGmjZAuROYRqY7G6BsVyWc6zU3O1FPhj9kRa0yBdR
sEJ/PRnLEjc0Z4vlggWAgeRlUuvDdiFaPCgH1vXMX2SCW9rRVB0vjmU2teJBpzhBXpTpZN1Eb17p
OZaoHEBD7WU6eiZUnFdCLjkDHuXoD10mOiVXoMdQMGFK534R7fQxICx5dfYqXVua6HQ31KnHHyC0
l7tn1b1AV8aYOzbOfJHoZ1wcas1tC8CYdg5gkmHK4CVSfkrr0b/4YZa9XeVNXA5N/goQgCNS/EFM
q+OOZS2kkz43Ds5MdE8U1lDKZrvr/nmwqboRRYN1lqUYgch/qRQNiiPxrcfM8IgU2trDE9V9ZYCz
akfGXfzJpnuM1NsMzmwyf+xd3Sl/5ve+AnCwdftXucPC38hHC8DN3CDKcMiDjNZkPkrvWmr9vase
oAdd5zC8mQ6YX0w0wZmserGz/5mPPj5+qq7dIUeZM0JlhWzECtWbz8TEhwfrnC5G6kgDxE9Ytjkv
zhAXc07v9+WIKWFQM2A2m2Gd8cqQIUCs+Q9hPjOiRiQAFf4TzDpbxyBwqkfKoInVHgLUntOTKH01
yhTY76kxPsIzsTdhzIo4ZG6RfL2wPifbgWJwFo4HqS1cJQrmZmrSPQJSTxTF125UMvJG0ymzouvL
IFJD61ZZZAIeQ6yDgPpxTraJ7V5dzpp4PWqQ7x0xCL2fyIbtCoxoJk0mlKjXSWrAZ+TSHFTf+wxd
lt5FtW6wbUla7UH/wIOZ4WWaKViI2SCk5NOVQZZzfQoUdYfLHtbHfElYrvbrbkVijglUbdJlRv2S
BR+7lPuv87o9trSFpmUROo/kwZoReLJf8NstpfFe8mJvnMVk3YNiJz5AXUzlOVV7P8uXDGCWqHiC
zXydkdb4RKLqnbisKelzsMMEu6ZimVrv/Iy5WV6ENThjiSbCLPWgsoAOMMsuwgsmz7BWMnVMf1fM
YUl8JCllpuT55qNL1x3ZAy6+XJaPcO6Ft+yg/a1xg48TcfJXEZ/hYc7eWGapINimHfFefl08/195
34RZKvS/ddCad1zZmFlUNxU5Hv6Jc8Hu/S9/4/O2BBBkCvZlZtKelTqhu6eHdUggr/LG3eJBWz17
X/GFRjwVfcEEtj93cStxexTBQRVjKatU1h4UYKyoLkZ/nGVBuR6CibHg/LxSRDBf16ttYDL4GWz9
fvHebqk9jqV7STGcp4KVaAHI1x1XUrt1e/SxPme3wJJyyautdSQslDLgfMlu5whrR7dWbH2Hr1Uy
XE3i9ED9LCPALJFhJFVexM5LouhsHhjpo9oUmugM4aGvZI59/QULU4uaFRIliv7pc3FYhJJ/Nsx3
Grr+nF/TBq2QGkKLy9DtdncqFAR3sdrJS/Eu8Io8mtCC1Hq/yBXHeNdOCl/izMPTZbZARRGAgmKD
qKhBXKNIrr+vSTwRjZ3sSLEObgeu5eMU14OoK/AsgHEDqjzku3VYRPHB/R8iYaE/nEwhfhEhDdBO
sVbRePXmeZAYLTevlvwwnQaO/ezPRoO0jpsw+xOrDEkW5q9fBxf7ba/AIrmWFgJls5cST6HvruI2
WsZaAoPp+yw4dq1RQlr/FlbFIoNpogO6RZUWWml49IiHJMuWWf3PPl6IsEblDMCQPDxYUJNeAGBU
00EJ5dI3w3RnySpMzMhvT3Ff5+ZOjDCQhmfGBiAdeLPYdYnOkb3VFa1sq4iCuyP4wuDCu59wPWlt
d+F2YBfdkqirXMv7txQwq20Rm2LGDU9i6xXbwEHfM7rLYxxWSp6kFJXyH1MzdyJPy6VQvaijm4bC
EfOs6hn9NB0V00ilZS4PmmKH5XOWsGkQodYi1w2RkNyAhNPG7ZKuzMqtxiR1GqpQUkOode6NyDV6
g6tG7o0+tk6eanoAqrkbBB5bWdBczjWTWV0GWeTszZua/TyVIX1lG+MwLGaT5deCXgV5jE9r1BCV
twBZ2vzqCs2rUFAfq8QS/HSmiLOhrUQKh40OYrzQAJxjcJJcBYs6fR/7xq6COdyFowcbZ2YHLdM/
eo08FTUtKtWgSOwpsweiA2Ux2kqfEcUgjDLi4wnmL34rXkUICLCQDXkPxxaFX15IzXXo1l8WJUDW
8kmCG5bmORI8pkPb1qWsXwU1CGQ04y24V7P49DtZAuNx4DQv7vrZ2N7JgiN7Kt8TELIGIgVH8uWw
zQj/FHspSKm1rWJ/O5x0bCGqxHCo/34wagdi5o066WTvnNT/z32q3VRdfL2hmmEPi0vkTHhOWw2j
gOl1Ru0d3ssEhE/7ErS1uyBdzQFGbju7brZl6r64/G7d+YYGMTJpK5+d3Zm8ZxnO9Frv/fwdUdQx
atXFTRA3QtOOmaK0qw2npK5m7sSquaFdE+Ic7LJApTXnwzUjaam3FQdwBR6rRO/7RFUc2cPDPSvq
VT2EX+EIvZbvJdeQy7M3AJRyfNFiIOFYhKUlDfrOeHb12BHp8fpbXTjpU8DoSwyZpF++UGma9lp+
0C+o1KDQ2FmwVtGsVdbvreQH2/jQ/urGk661XSWrBreroZpr3wN5GaKF64TsITOMQfYk4+UpGd8g
E05m1bWvOEh6JEc51DQZd5vSLEuTMB315xnmBypUMw7hVJx4veI/6tbGkcxccJnyycUP0wvw6LcP
FUn7QJVPU/0LE70DeDPjmvwaBWPePIjQdQKeTepOrK1RrM2VD90D9uRHmHNFhT+pmqIL6A8KDBzu
/KE+0niKYIbeJh99TCW2vwo25Vh9++cRlSacrv60uw40MPR15U/u4h3ws9lpGxSxBUBuyRTnXZyg
09daKWs4B6QpVQJPJrJpm8RMEENDCheZCnASIr+XZtF1ZkmDbDITykp+oeQL1us6xpg08bfCkjkz
fOJvLIARMAK6RhtjtAc9PrzJWijddyOafJIpiCU5j1XX9s9j/55bzA2YBsnpP2IZXk5ujB7zDZH+
LfUPs0H/KsBAvIwPm3YGLiJyKYdqIrwkyFF3N+BJYuxiD+RPr3QqBN8jDL5BqJD/HNmuByennkMP
X+stGw6mGdbCEUAPKSVBJWXiY7ee834Z78if9+5U/jdDcwzmIdmb0M0ZcFuviXJ8V9lJYT+kiMTC
GDutOJMkVtSaCqOlNz30fp4i6ihQDw1GnK8hwM7zpEOqSW4BYrDoQXD5grD+KyPK0Is2Mr8KzEDs
CKweo5z+kQtHQZMBsbX/utyDgeXVksyCqDxPy/BV6+NZuCQTKWlvst/Hpo7dy6r3KLsr/fysyoyb
jTwdHHn8lkHnPD1PPdpcHRSwnN6APQSFKPUhMJIGv7O1U4Afu+jS25/8CHiFaG0MPhh2R25ICnBN
shF97GXDMO35eBPDYK98ls0LaRTRVfWL7AUOQh1oxqx2B1+egiD6D8riz1tLWoBASZX4JfmXmldr
1na275BqBGwM3jyf+kBeIt0xUI+IVQ11xFaKEZZYqSSGU0tkbn0yVkvLJ6XxdhnGslBgTlxSPPKp
BLRzAGrc4E0AqL/4O3nd+CigwGXN41wrFbJPokIPwGK3LidyOCE8aqUsER57r5yr5MO6a5rrCO8W
6BhlgI0S025eO9hdiz0URsrFe8lEOQb3xM+ylf6oOYb2m61++yJtcQT8hQLizRT+WwZswMIwfhtL
5NJrTHo5WLPN7vn8bXsljKvpZUuin4jgQ7eLD6j1p0bUvNP+wKVItAAGTkQ+Bb0B+stP6NQhEDNu
7zfoK3ufYpVQaHtoGnlKDcaS4Br6HMV44QTVbpyh8jp/QdtOPnW5TI4/1vYBbegkCwjCeYriv5xB
5b2qr6LJ5LZCpRMvK97WTgFcyiMfabGNSIDWkntsfD0vVy3LNICwLBrYw5YeL/AxUzaiPogb+vUf
EeOOdl0JB8rT8pp5NXuoLMARxx4xkB8le1WkUSB1Z/c/EDtOqNXWacTiM78EeYZ1bECVSq9rpJj6
Sa8Ug4Zeur/TiYqmsd49JUYIkrkT9jRECiloSUsU9/r2Yiq1a+33QykJA6+NIrJBcBmV97aqSAfl
eoXYS8HQ8mCL7GIW9noKuZ4fssTvbDICPsjX4PUBWk090PkvOtVHWJ7hyiRZmCUrZ2f6tkY2UQBn
ajPCh7/Xo97E42WpzuMiUBbaZmJzjR3LSwkl0JpINJux7hxsakdOtUDPqiu5wefefrvu5jAWluSq
KhEu/uL9UXbp8wmlLPDe3QennPoEuRs70UgzhBaI/1XS3LgJVIKdoaYYwfuCuZnECMuSp1/JCath
85Oo8dxIYEQKH2pOUAi86lhVzcB5P47rGH4CsYkb/hbOuXyizmlC8XF8u4WyZ1EDIpBBqhICxcMo
XKr/Jb/ZGpgSpIgjIcmOGSrXRBKpIaWTmm6k65w/LUSJHfPTAagBW4PS8WkyZz2xINOI91yMRjMB
d74/ST/BG51IDQH0sUq64pycXU2bh5HOnhPQoLNHIAuA1/kkgSvmcIH9TiRd9ANXuJ6nFykSPAh2
JTLu4xr1m+KV/hU2jFL7OBmpU/rO352sfYnYbrEs8URifgaxNSlQxKLl/shcwXRYiH8/okC9R4Ie
jbZDesXXzEUvEHDtqRDOkBIT/kU3kk/x2gVEqNW6XKFJZDV/qABMbtoFG5ThDPtUP7Pid7OrlevF
czBfjBcOGu8/MD7eTi7gio7whjRYBJz7uj4EaMFKk8J37JN3fN5dciF5wY6fJInNB6IB+BvHYU4i
w3IXhbI1aAfMBRlCle+4SYqKhOyzsyj/2rxS8kRmVbNQQ6CFg5n6xIVUQ1mnMUBq4ucUVn2E/s6b
oN3/Da2cclt0vw2ot17jnNeET9SCkSqTeDipbZMLFCzbJe3fdHDkIHg5DTVA+sGBAsBip+QdXwB6
y0gc6TwHWMH5rm0/SbG34R5hAWr3iXIgb/oMfcqLY+IyduEUmataFSIDrOvoR4QjWU/7KEXy/lc9
KXV5NkeIAbqhHrjGPvgo4Pg/Gj7Q6/7D4Snt13pansBjMXYVRLzYtGqekfB4dUvF88E3zCwty9x9
RbHaw7uBdRrWitIyif3eyTVBXt0itqYUROXOUJqxCSwjbK+rBu+ZMowoxv6yBDAdd92sbF44rp2C
CA7DE41yQYhQ5STDdkhgBaqjJkZ492sEM5TqLN4GjeKD+PBRYQ6QcpKZWKimQnIrCI210wHgU+5m
dwJ6iGc61mTZP8YsCCCV7ng8h04grwl9MqqJZ3Ty6m2xCwXlRFzyXOyhQGmYoNKNwemTr8HuhTjD
gqWWY9pY7jrVPE8aQtAVqcaZ/r8SeK/fDfInX5K8VbzCm6cqDKcgzRw1aiRfJnzDjj0SalWpoaCm
yE67NZ1azLubz0ffg5xlYVkNrC0eg+AWz2zC/2JjCv1Htl6HtjCjKUmYA7bxVbvR0jMOMjYzZhkH
NFcFuldUKHK1hyf/pyZqu/aOs8ikYM6OBHngcoalRgAGVNrL+JxfykA+vMY16ghaJP6KlCpsYpEK
piT9HHRR8mhz4BsK5X+tdXgGax5VpgOVdVgBcWrQbXHq0WSciQUCyAjZ8m3PhgBh28dDy2b/t2S1
WE15BdtCnYUFTcAaXcMMef0egkfg8ATnhL9uzSbLJQCJpyTOVwFAuIJ8qUlKPf3EuZy6vTSZ6M3l
upm28hdKA3HRawBodzXyPLUtjEZYGSaNWI5C+IhF80LgUefYA+FlCYPU/Gquwnd+WAcpnAzscRVR
P+IijaJEmlApqwc/4blltgCLgLg3gq+9IvA/hIdYg3czNoR9XlmdLWhBwDah5GPuJqejr/Qa/LSq
70PzDTX/M3aboG73a3XqWNVAoX84p99cDXP/oljwYZd6317pT3JLgyJmFP523zx6Bd8AWZQWJTbj
yotzquAxzBUNVaUvTOjIYMC/1TT7lDq01e2vNgYgMd8WGQ9K0hWBPmFlaSQq0MZmeC8+qJebihVR
dLUmbPnaodywurzpXRHdjE+KYIFF3wpEhYo1iSZO9fFq4xHxfCMtAVsOfV66bTy3AeuRI+8/jbmo
Gx4VXLqPcn51ELkmpTVh0tX46QAJD+IxJVAQrWwVvOPQvh04f0O0RiyT2MtySpgbsU9XOSQQxFe2
HP+4LiotsiEXlTZWM6LTQ4QiFtbvVE5ReNhdMAV8f7qQMhPY+bLeq4/Gzko9hgYzUXPqRVQcycP0
ALnRsN6KlKXrX4BZ0eqpu4up0ibOsXUo44VGjfQA5ti/7xvGDIOr014+rH2FXpvoCyqOT+F5zQ/I
2MOjh+Lc226t229mXJlTzL/NQPk5AkLTDy0xdwHwd8ViIeh8N7RfPSpJK9aljbIbG0Jt6ttBaSJg
7l3ycDiT3dSuNqGVOuMPSpgwDjMraQN3wW7HvaeNXfyv2ovXOfRo1UQ/FtQ/+3OxDfhldL+rPw0G
+knTusnQirP0XU0IX5I6xPpj2n2Qq9B/z/2OlGGieVsAJZvkeLTXDY6NRFzmIl2EmjBUAVgslTux
lbG6ZYKDAilCUXZkeJ5bNhBF4decYyX9E2zyt+FwhP02tnglojAsqVLkJpbUR4hrsENGJ0xMzuAl
rZXnLML+TFrRPIZfFn1VAZbjC4rm+nPu0kmfn6nELx29FlEYDfYY2q7aTelvRCpfptcjfeJ60xJ/
VudJO7FqVaLClt2Xq46WM/SC4Ly+h0DUhQO7xJvNk0nKlAZ13MiE9BLwwaWO6/qfRqAPPM/So+Cu
6+Gyp6wmP5amNUiShRE/fgdmMGpB+ylngd8sEEufeEvQeGEuEqSx7cBkC+1JGK0F3qzfQToQqpWB
ZlPXqSKMt79h6Z2A7qnZs2cNVjdpSew6w0SCKBYOtB/wB6JIRsv0XG+mcNySCN+dMo97JDj7A7Re
mmxEh7XnDcYUJ7ezmQf1yes11W0zYwEc7aWRH+8LQIlA5l5DAJv6vVQATsU22PnxmxYz0Qh11crW
DB3yMHksx97bEQUt7axCjQ4D0ghluGNJL0MaruErrsJzbi/GgF/cYoBal15QRox28uhcTRmYL+ZH
rNm17JnqhAiakqNOiIbtjahjHpsmpHG42F2iUmAYs/pAXmIgIwt9f9XsrNCXgzvN9yfFvXsJgM6P
foXFe3iU6z8UOWEALm+G24/k5jxrJwwR7WXre1x4TZmHA35Hf/5GUKWMPhprNhwbP46oJwnMwg2j
f1eTZhSdv0p47YJR+/kGtClA0gCVjbed0TRDbMPWkwDMV8EXNPBUi3DNczruUhiSyVRXl5TQxZK9
rs7pTt/my+MCpO9hQZyKsHNCY7EJy5r6SvZqOmgoFKKjYscLV1oFOlDTnojEXCvcfsZSiYO4T24W
xUaS+RGC2t14mH6GlT2e/nIsCwNd+ha3y31rLOHdG+j5oKTTSOua1llt3QlLVnav7RVPv//ARVwc
O/9wO5eRJzP40jbCmmGswJNJ8UL5kgQy3DvKH8ynnri0wycQE59gU88GnZe7KOGYtaHTsw+FBIln
ohRzg2U2Mth2ZJaXHTKCK3rArjjdmoXVrjYWimi9JO3uFeJHHHWZ4snmy/3ZdstO67mR2J8j0RTo
JFjdscUv4Kr6XbqX/uiqFXiaADTD55J0nnIzW1Pib4xz6XaiO6HK//eSTw6XG+eZt2FuvPmGq0MZ
EgZfNauEdKB9mpMn5oaS0nDU2aqC2PY4haiGVV7Av7FYs8NyDtIJDJF0aZiN36mYV2KjN4Mauexj
PfLC58sDjGEtLDPvV1FjXVAjjaklKzZocPz/fIbdscavkE3AI8UWbWIVxhXVk2o6IG1zNrxgvLGo
ss1UOCSg3D1WEwdOjnsmmyubQmO0A1/XAiyGAzuAqRKOJasMhwihVhLmhv5PZj3L+BE1nDYdFOUv
I4bAikTBBq1LRvLdD3Gi343UwqXPDmd6rQjTsZ1PgfUaDLy3N6fcJvsJxup1YFu16f3Byd8q95Ic
nAcf6RvuJjFyEupYloWSH656kLDEmhqEEnQhvqkx+UoryG9flb/WDct/kyLI0ndYcv/guTueGbvy
A16R3cgiOQCVAvCjMNZeQZdeBWFiaCy1TaMTjYemstD0LAjQuszh1vzKHoTVj/hQ35TiI0h4ULcR
maQCTd0pDNcXASL3Y0PgSTDuopzeEZDjea4E4bly1Cr5qQNpGH9UneKYihejpE8UGGabYGY0egfm
q1VsZIxH2/gUwgvvsZxQvX0Q12gT2MTlJFFd2b1a6JYtJJpxOfAOf5GgMJ/QBPWvxHQRbC3KQyeN
o7d5NFzLLu651HC5Bm1OX3CY5z7huLFV6lzdsOtYV87E891bpGrXn9SjmKE+VpZHZLYXydAAwzGq
PmAK01uBJIZ1/J/7044kea1NwbgU7FhhCg95eGrV1aVmOabtfyJtoEEnF2SqbSuBezBZwbtXjeIo
v70NxPNFuFLtNP4O4sqLa291eY5RrHrSI0XOobi41AU27fmY/Gi51W8hwK/LduePE2BQJTEAy5ck
UegnMeygPGYBqU5Q9TChpH+bn3ffNEvYGjwFFIqOczbgRbUPFTXNdWCYPMCGL9sNYLz/89GOl3V3
WYnSeAQ0iCxgDyCQWZdhhyQknNLgoJjEpgBtX/HEvR4CkkVp22GkIeFgv8kNlma1D3jSLHzZeG3o
dGcLfg5STk3wN91+xTYP++fGVtdFd1bjYMKP9VmQxXEvvnv5dCwp4qwggitMriySykoslBlfvu23
EzyqYWdHg1gTA+TI7pBHb/z/qpek7tammFxSCuDR9iOMTJY90gZCwP6TQHNEbdt5TLMbeG33vS86
8jay53AW6Pnqu/cCAKkLCMwnhAcrzGAezWuJULuEQJTQE0jN+OWufhErMjShT6VqHFJuxns7o7bp
Io3rw3/O4TnCUsh6EaFxv5XaIZ1igGYXK7OPr6tEsYFQTwanKwaVcyqwT9ONDSXWuRJKAJb6Gftl
h/eXr665VCTyOXkbWzIH0SVHiFkCAsEch2tIpC+lCF9mlRAwe9W02naga4PABI0+KVRr7wOj+92U
c5OFor4Ot3DzPp10e2QYcbS8qIjKhAiBM8Cw7BxcrHl8oblbC4mOcz3gGCEtigr0iyORHWOmtKho
egx+d3oSefubdQK3BcyFEo/hGZI7PSvIa03wUqT25tqCZm00S9Xry+YWihs0fTTQ2kUxOEBkYZkL
ze0SawkV6pAIVzq/DpH0AoS31IWKdnlbTQE8JqjB8mAIGL66+ETlxF+3h7v8JKfzDSh9fiyCvPmH
V/ZnrlCHIFdadRJGFhTr2ezBrjGNGpwBDibGlzTHZVDaY5FLw9hZsLMotocQ4CMJ74i93Bs7NLXP
mrbw5k6GOFenjOLSKKfnjeidwjc15+ZhFF1rGJZAqVMuYb652oleApnTclT6yq/Xn9i/m9hkgyAY
P/Z+cRTx5rPpKI2oERmehMmb/W9viZjSCnFxQ9RjDH1oDUjTlHUfcHPUKeSwIYpSGr3vtwaqrz3b
GGL6C1D1qGm5gP8qY8/4vtFzU6gXFmKe4YYUCA+mJyVw5Vi6WqbiKzDS+Poo24ZGADtsb2c8bsOO
755TRBMJlRkX+SYkZ3glAS1o3ttMKiq6f52QGDMLtBhlqx3dnFFsYI7nEgOGKHBdZDt4+YxhLuQ4
mWZ7MmOedx6tSWC426zg0Ve7KzCjeOj0WjIycFbJNAaBtaVMIW21qiRPjnrjHOUuSaJEyXjLxM5R
UEFdcM7Kvxpc0hlzJr8Ce/N0XZ8qKAE0YCOeAFX+LRPSRF4rSm1R3nk54VFfqCxirQunhRu8TeHQ
devsWaFC5Gwk4pGSJct7015d9ZNUf3HRcxXiQdXshmjAyvoYSd9cgaDRm3cyr0SVZiCffgv4i24m
mNRAf8MGiAqDGpgslDOowFEWA95vE2WmLFWpsY7BvVXA1qnQcsHkkDSVfMo2izUFhM2yfNbp/jEd
De3N9ExDg4xxeT2oq1tOc2E4nuryiVElKhKhpl8EmJvj5Nrk6wsQHhrMvFB0b53kdhW5RVFBR0EW
haoUbKjgWo/B1z0kSxxp7+2Zqpnpt6iaEyuFsRWN3W24HBKf9Dy0ISoYaKvWI98dqd+2UVDnnIBi
VRHnbNatc/0J8Bzetc5zCuC2gtwox2cHzr/yozSNbHVYJbpPm6oK4jhhqjKx3y1T1/pgTYONFfRU
jt8nii5rqnDBPaAacDW5Dtry4DTH5eWAXrt2P9zFxQRx0+PT+o1+UMPlpboOlqmvTmv5rfmvZghQ
cHQrW/foYP148lYV3EYrUrYqU31sDWrAPeOvkajPCUlwPSOYz0CmNSD+DKy0IPTHSKCfF5YUTNPF
bchHU35vQ7bN5XLBOG1Q0bKg0oZJMTV6i5Kl7UKFROMpzDVm4Z8ZVzkNBFMRlbBoe6O4QlsAL/Ak
5ZtHohEwoYtoMs5UymtJiwLZXp6zNhKTFR2i9scbwLrAwgntj5bbQ81II3qx+r9ADPeDE96NE4NP
0+PqeKZTUhH1k88comOzXo/Wd8U8zVDP4dJMSLpPirh2CCuw+MBCSChfVL6lwpze+Q9UrWMF0XXY
cxFtRCiLZNH9F9/DU/0P1aswvmC++fjmvIFhd0l3Qpj7gt+biBm5mADvSlGPy/e+/8aBgk459edw
NBNn1b392KLY0UEuBufziYnHoKTuIj7f4VCKQcNM0hVhTpQf3JOgK9IISJqm5I/sZuvFmjkpi07w
mMFO0igaOJNFmUnPKGFvgJwTh2CwOZHKiOSRcry1Fj+W9Oby3I0V3j3OYJDA6Qy7xHtJ2LpxGc72
ELrPhluDfM5Emy6PNuiko8dox2w9ei65LlSvKdAW//Tje/QnspIFvcRWGf6go7W5UYKGkgOWSV/k
UBZfCxba4Krj4dHs6JJb8Wc3RhaKGXp3eVuKypntSDKMdyo2Hd9gUiYCTRTDkOC9BdmOHvbYLLPY
5f/4OV9+FTSnnW4rNH4aq5icwiHqAXxiGJJ4j3RX2RoOenGpAK0iWcHc7VhMS+nzyfqj43tqqxpz
cvOytZRHga5JyCg44MubYtpiG0thfNH/45CbbC2VdG3bIOjF46c3OAasKIryx+rPHyO9xU7CykT4
lk6sN3kA8UOBMb7f2lTPH6EUSOuCLeJhe0EE7c31VyrfcSsMtQKie9OuG4gVcoXxHCQ387TET2yj
A3TCma8pCuH+tCmL4hVmlVgxS/HFMixqmQU5fz9lU8WphihkWHAPJJvnlKdRGj0Pyv0GKe5UDQIK
Lth8x/yWcfGf+zxumqMQneOh+oPP4jNcySjVa0LaGnoMXM/2O5TfK3R6Tc444s2stfM4v3bQ+wJK
bAstr9qH6K1RzKx/S8yYa2RK7tcerTZnJ6PKhr2xuYYGSOWX4Z+47Wzv16h/GAwLxqvKk9BcpdwB
hnV4/O3VUA7kgDvRLuNVuWW+NrXiu0OfvPd7mfOtdbYexkB21qsPm8yJrWp7Di5QsrWyr2uQEPbg
frvaunmAWdVjtKrdiQ0+Q/mE7mkTKt2zOz5m9QPrRacje5zQBNw7eYlsk840xdn5DpCuiglZunta
M+vnlbN7YBdtooymdnrfAWvNaCjoomiAY1a6vapuXh4blQR4D/g+gi5aMsiXiPTU3B8R1VAtgv57
6Uo2QxJj+k0rUbChsaos9IkXPunAR0jiO1JX9y2zY7s377wSGqm05UdUtxMSM5j/0wdkTfBMIIIW
m2lwbEkxnpmpuMK32o/JoKwfNd9SITvpUr5f7RU4eHizwSyShWIoCa9XQapmEn5mq3JTSDhoR66G
O1i2bS5opzbX6QtPZFIl70KhmiAxC7C0QHKXOhqa//5PdZAS9NicE2v5lh2SWEoMiddm+mRWtZLI
tismyasJD3e8IzGtVLzFLrPQjOInNNaw9otZ+Kmkk+cG57BRtQ0skcLT022r2bR5kWHAuGk475Kg
pROAOv7BvXvdjI/Go6bS4+Gf0SMMgC5XlI+tdmF2Dr+rDj4r1aRrH9hrjceezqv5L2cEWYZt8rmW
p0JYG3eZLxw1NINoVKQeNsw9dWnJefnOSKThuvnrXsO+RJSt08rTFJFgfqCuciY46vQHT4EXnUPx
V0sPRgQub4z6RMZaL4ToPUN4vBSGEMqRSYH8Z8PK5C+ZLql0HQ//KvQsXUqwCnvicKyDDcK+D0k/
B0oZ/0zenibf4w+LMDgRZgXSbZCnrM0BPFj7nI2eapg0XPk5jOgKMMvIvhR3s5NzQ7Nvm3gzv1wA
58kQTgevBTDeTxOaC8/+cRzzMRA/ZQaHggrSotuwhcMe0pRsKRjTiq41sLK3e6wsOHd17cC1CmNf
tzt8FTnRxCw4QWXkKQ4+66GgS/gp4B7qVGSbY/p9N3egBkXK9X+TvkpGj/eJfIbRpfr5jSJlRzyn
hLbQe41NvGXlMBBs5LODf21Rzi19hilhnk7PVtDsa1QGYMYR+u8iSaVOxNxw/ywmVBh3f8RGL8/H
ujo6kFCFunWB4xsHebdwy5rMWamECZCpuSnevVKy0WN4P8/m3AhmBjGzKptaKAlajglPhES4xmb5
F0LC6BkuG/MsS/UzJKDCgYwfNtkIleQmV3yfZUCPnD9eNEDGHB3sgcQeIOzB2Aics8jvLrq4JFh7
mgCsF7SIldIS8gWSRt0ILagbgAAhr2bXEl1iaX2v6qIWNQ91XivdLprnIIGbDFYX4Q+DVpidIEa2
wYnHQH3qnCn/zps0Jk3wtM4IXrc8lurX4FwGrBII4ZPz3u7kbjXyzwFdMdtA0G4RPEQaB+Ub18xL
UQxvce8suHmBp1ff99b7MMsl3IlxlMxhipevk9WZGJJfaiWZ3TNa2jAzWT8SB7dz80kxh28IWGKw
q3DUaLc16J03jussOlpWJV4dfMaThmaZ893NXsKfIhyoUNb/jb1MPxHf+cGGOx7DFcueBEOCv/g0
XWAa49rW1kzpTCbAAacrSZvpniy+CDWmx4LiFuCr9GGmEFOwHVoAIcOQJ44FDL0eFwfj0mHfCQtG
2k14I9lO83vwYS87sSKnzdd2talsHkU+u0gl6zo16m9AyZ1eny4TNkR2lq7SI1jtQvzLfOzkfP6s
xXlyUZybVuoYpFYMfKmjL9aGv4XSrSAGaeNI1XQiuX19GshnMJVTEaa4QdpLygT1hDjjRKXgy7TM
2luZ12io4S2quLaSFJOCJ0WA6tmghhVz1dLbzolxQQ6Z+n/Q6xyZe3VBdFARiT0uposrjaspxlWT
T955vqkTdpI16E7vFMYSQmNMAtjaKPLrIqFuNIl7WmzsA+v7k3ruF7wfs2Os1lGc8JLei0YkqTVX
L6GN9MPNq4By5+DkCJmfQxx/7UWhrbm4omBjAHiN544wsZU2dzpm10MP/mMajk+BmkE2Vsw16/F5
soGdbyXZ11E/E4k5omkY0+ncfLqxu2EA2jfaU7Ux54wmc3p/UUPdWNjt9MpNyJCfJ0iufk4AQJYY
QEUzPOqvjLfNmJ3+qQDE/SG1h+WK4gP6ECmbXbWnuyKXU1Hys2iXVaLb2Zz46VDPsO/cces5Vmo4
OXLpMRVUaddRfdJTCpCZDo4+OIgb9iPWXSkqdx5HDkwDkpT4cqKDgoPL8M4RVbUd/jcGIFujK3oy
7sUUZ0OnDGAPHu+Q7QAOnyIcSR1ATBxJZnVERKuJR6YOz8PYbZfyjVrgL38tTP/BqedojSA/gAGx
cBhAwcMZfh+isdvIpQy4HH9+nTknehAOdKKdP4Rg2PCrIXMGmpxlpFdO9sMagSBQwmtHusFnGONX
HZ5mQL4UvSF3e9rruSKUqHYKeQtPbBcM4OQ+zOZOxHWyOgCd8sXpQUVY0Udfz/z/XV7eqRbSJmaB
43MLTghnbI+JL9iUHmB7GKygyKAnq2IisgJzMs53unSP6QXNtORfiPtQ3uAnUL3dTOgxo0hCl+3X
JkrXgFvmQ4zCifDQD3DuTHuLlkxuM58u1Cu7SLppfIKscnyWdnZraJVjJlK4NKzwCAO7wpI9Ah4q
MPlDB5B6ThHwYHGP2ADB6rrjZWyIYIlU5aBM/bKMtguNe2kM1we31e3AiWVAp6AUqVWYz7FJssnP
Htd1qutI+mR1yTwJ93g266bt8MWqIfW55cxnmToVkT9P6rySwwia2s3cFCsxeCtJe9xR4Hntx9SL
/11O8ld9OsFE+gTxufvXrSOAMtFXz+lRUXT/u40d2txIhKGA+ULQf9zSktvII+Pq7QsBeOsy5r4K
VkSDvpH9IJpZEm58u9t4iFBDmBIL8Ckp8qg787tyhMv2zPXFhoIaaJ+HXBUJcKyd+JU93SbpImKn
bDBSNrkbpKT+Bp73XBYIVoY3s0XfJALI8B9K01VYepBKndt0z37gLbiS/He5H256+CDkamGWAWFo
4b+9L01QzqKgcl+1Vpl8laAen+5zmYZhNBwi8LSpr0OOIUhAKCQKkWr4NVDz1KRtBLobm55Wcp4+
dOY4CGHTGgjbUcEBSYkg6TMw4Ohmc5TE6ezpTaG6I+q/0/CsOc9eipIU/ynR1OyTFGRwe64CQtEj
fbk4CFg33Q4xkj3b6bv6w3lVOsTP40BrRGZo6Oa1MLkiQowPCobwXmd5JKqCrt+8EUfHhY1Augdz
6ABLpxBWIvM9JQQqEpYUOUu3orMk0Y7YNgHx4lWBTPV9rH1bZQ4fFuqQ2K4r/h8ZBw9PL3UbqNBx
sJYWaEC1oxZ4LrdMAqIga1BY6BhA5xEtrG476WlKNSkgClYCfQ8Q/VLiyfErGwkLzVaT8dEfbxbb
7kdPE/rdOnO7zaK2gTRtmJobh9rIrRCijsHQ3b72g/s5M6KWPIH2QFCRHOkKE8/WWpbNIQNvMIBg
OuPMurn252WVa42dS+4/WOzHgfk2U9ig5P1N6Vz6p5niaucqB/9Pwm/4y29aUQcwjh05cXAogvvV
Kv9tnq5wL+se61Ue2+afunpo6ZIWPLSm7ULCrNbomwhzknVcTF7od9569HYcBW5FwP4tz6LMXJmK
+XkznygNa9fvzZY4cNguAlUjK4HqvOZ6UJdSx0ruuUXxC3uU0LtNmTVezOrN29x4Yx8fIpWZdcek
V6478KN/co1ZhKVrixItNtJrqN5yMC3BCfrIsvOHpyAg8gvuTu9ajzjoelforGIBtOIu9tltxoMg
jFPvm2qPYKstDpJbi7WJdiAmXcZIY52dbccHPi/azRefYNqvQOc9CgqsUbQK0LR820/p/k9zc6a+
+qKJNigvpRhTt+JxvOVeaIutN7bXuPJcEb0n/hGlU1Wmf0QxBuGSFdtwPvbHN9SSLVzwvz6DfERD
uSyd2twoGByP3ysg5XU4paJM1hyDT+CNezANiVDkPMGy72FCd7BPyZtaTTzjgMf+R61XSS88cawv
hzkx9I/KoCe67tqM+55JgjcSSPVVugAluYbRNl6O5k9lAeZeL+HqFc7ZKjEwPKg0h8Oclhvkykps
Hr1/sgQqQ/vnyYbdJmDte9LKGo6xtuV20JA45gyQlrI1pZV4JRYRgcnTXO7se8bC+/NSO78lBGKh
aWWNkJIczJgTHK3KuLNKEGEsOffw/oar509kEGu7JgBcThSCeVQEpdzum/vDUd/p6/Y5hJ/VYSka
dQrAscylnKrxNHQb85yAEORsyw8TKvg2bRArV1cMY3888TqEp9GM9wqUmheBQNNvkaa3xKXgvIay
4Suzr+RnWVhqzXR1dcjWWk9oRVOUc+k3jFeHcKVne4sPP3LtJPfy3U2EZTR3qZNKINFSsiGYiPpY
7dKzhV3hRs2nwmjRGz7LTQIfPQr7208Qtg6tKD7MYJQW4mYHsZx2bNgQxro9LIe84S0Y6AM6B+bp
hXN1LqtNIyoZOoo/kha6XEIOn3OwsI1S00S8g68Ow/bXSDuiPwXtzfpJtUMLOQciR/5agg49q+l3
P08moV5GwSPThzCpi8X+qwYMT/ffd/y2JD2AIslb/Tacd4jzQlVcPHdAXJ88JKjVBB6Ewf23zvO2
ge9ReQqSdKtuH2VBDegJ+Kk3WGMxkhrGIrqi8fb6K8MI/l8nwYOvfKGaiXcoFAbEBoLVuwnz1r8U
3I7PmgSFm9PUAOqlQ4Po1WjG1tCW5RSTCtwP8/EP+NDSIecQ3PEipIYrMNxR2usuzdZsJnVa6E9j
G2Y0y2LKjM9BIOxLc4Eh3sk40MlEgG6PWO4sNli6MsY43Gf7v9sUmULxSk61CQqhRPt0vGergyMp
MX8OZsc/dKW9bfQBj+4d2ArWvHPI2TUxccumF3f7AD9Glf15Bd1R6JhyvqxVklYo+Jkx47+Bsifp
vnpNGLcwAa5vUq66SKeyl3+6d+++WD0+9wWjpfcelZmawdFBwXnB5lPhmYc8PzAaoPAo6aB+zDey
QjdKH11CSvL1Ab0P109Oy0xgUc0yHt/UvsCm+XKuBcNSiHwvTtI/CTkXO7UDUmHrWJEKPtVKkdTg
1u7XFf1cU6YgT2piymXTeo71bYS7HdY/hDM/fiJzu9Tw/d8QovOlD4OOZf1lofwGMMrl2G3nesrO
XAD17mgJ91Vxfk4IHTyJP46f2EzqpplZM1rPD2rwlmXZ0Z385z9W9mVDR3CAQqnZbX6bExs8XcjT
Uk5bLEzOoe0POUTMg75SKg5k+liHAUeVjXmZVaNIYSGUT7kfTK/fvwacWGB7G6dUnnn+EkqFlXtK
nfLOak+iS7iDE4hsS6HN3h+D0aYbNlEpXEjbRAyXY5CRRZUk90QkY0xCzeESxBcsd4WVogl+6zsC
N1pAr95z9eMDLx1seisjMax2+ZhMyzI/vS6kgmV9zC/+eS0G8yUcSJCngnzQd8RJC4aZh3fnxgzv
CTbfMc02PUQye+oyFWymG7g9Zygop9LshK2tX/PDbjsR21DR4+gumQQcsHnQUZTouiRMDahEdhTe
nJblU0vpt4vgpP6rwLduKWye3RMUhMnaifVgeeefrJnIPMqb894n0eXqVXCtxHMp7HSBSiiNnh62
cZ59DKLqpohEymAHfjLZA0d1MmWWYCM8VH3J7MYW2r9YUmmZ2aSpJmDdsemmAizTXNP8kk9XtdjJ
qBSdzdYOf41pzWIkT1u6PSpI3/+HsY7lRPcUDQE4Y6xevM/2ZgTVlkGBvZpyBfWHeia2G2LKi6VC
ruluOvPYI976WkG18gVVUPal5gpfDpzGuorofyo0Hk1gRBaXTI3SqhlH5zW3QsiCD7RlpJ2ukTen
wGsDYYkDZby9MUoZqCWEmDNNoN3e94wE5QqRbXcM8U5CA7TWz/qwDVHEeSXitu1IA56/0AQTS5HX
EV/gJBD0rI+xZaZFSo0HU9sBBPIOPSbM7yjYTllLytq1EbEP7w2Qjr7Sk0m9IT6dkl4qSrZ7Op23
v5l/i+Jcl06gHSNW1+ZDi9Ck+TjRkv5v/9ZD/C+oldznfs3RDYljlWZemKqlrI+4r49E16482ItG
aZlz3xkHMo4mFaOLcSn/zpw4TY9zAwaLTetnUfJp1yKPEyZui2LPdfthKGyv6hKYZLufowTRmZsz
W+QEZjV9wGw5rUWGgED8zm6iALQXXLgMTFk7EC7MdBso/3NOEa4tbSMbaPNVsGKaR3d+ssr+Ifrq
GM/+JFG4GIauqwW+etaUJOTM6v3j2RXOzO8/NGQ5ri8uuf2eREnSjZ/WH0oaSiRqrVFj6DZI/0RI
HJDCjvG8b7r96k1ypXn6ejCN2mAK8d05UQ3Nv6Tq4Tdced+4PhcmW4G059OC/723xw2+lUs+S1B3
zEOnjyL8xYtvObZp1e6bUoMXdEuZAMkKT2/2Xka6KG6cDUlfY/f+JJHaAfXCsJOv2s7XXTLDMqJm
eTWPoJGF427zMqheH5kwAVakl8opAV3lKSivtXwzqPLsJf5z3iL5/iIblUmy/UWIFEYew9qYs1qO
YkgxwIBXSxIh0OY3qplhJkOIyyp7S0oM43Q13iGAzcWIesePW3HIZh06SVdbw7B5810UoQPyPrIH
SdeF2qsnxLUkrng68xV7aJmw9a7fqZ9z9v9q6bXjIxQ3nX1WfyyP4Y58MvG7px4tl5iFQVP7sDvV
GEjK5rfq9y/gBuhJ3JynVRdC7mTzeGdaXpBOJFCHSfX065+92IombOkZnvTytt8GagYuKqvQ30r4
r7GPMAh8By7x1fw7OJ2ihUOv68xwzt18GvvGMv86qCNFa5wnxG7tjJJzlOTy5PuY2237rzIbMH0m
2WL7ZEn7D0WUR2NlmZCoKa+KZrrH/4fgVoXClr0t4L5FAdKgFYXWmc9qchV6TybBltY+4/rF7hs+
tNa8M5pfL+tEcNKYsBcE/fBq9ttdWKlVcW5ANauw+ifz5oWjew739vUQQnfYERsxv526t/NvcMEM
kWHXJuAO6ZRE+7AeVxG8AcdApVMdYQpSjcW38WM/hQM+FBmqLDyc+JcTwEXumRPpB+RWp3NAVkFQ
5tyCwWb5q5EQz25BOo5tMA3AIQ5A1xsoEAfzflCodaVEt+I4mlNtXdsGUA33A806J4POAQhctItX
WHk1XYhLBw0qahCxoLYZ0Ka9HvcpKMEBn7okXQwVSe8EBH3sve/7PpncgKcz+fwVVhQk2Atwk4HM
p1RJwJ7E7UrWktTCYPqQXnbS+dT1pR1RmyTbAnMH9gsKMfnci2HxoSfbZ3UztdL4EVjEzDQeLqrD
MFDgEasrT0uODLBxLZYbx9tn19jujMcQcQqUzURyk+DKAJBz72CKl4gtJ/GYuvJAaQjxFfgNLRH9
NoltZe0cj1ZQfS3kUyTPVRleHHcAbLrS8TIZB3pI1fGTaV9gYmLHsMq3Q3X8n5bGbiuAKkfCaTFA
cAirMgXmSj2fLtBeJnBTt3Vfl3rwixrcOD91sPsRDmYK/yEQmVhC5FN9+/pQrtptZ2QgVfslWLJF
EtecLQ/XVT30fFSOmGB4u5ZQHhrs6720BtYp5OhRj3j/xuZKSZTwsS42mQkBSvyEHDxnLDMTdIaf
BFFU3FI/tjVWgkllC+oUr7ly52YOg/EgM6MaVPzzQTz95YIG68XGsxJFsEjFnfx9Z2fLzddXXBBj
IlDLdtVmw4G0MvqHcHeAuIc1EA+xg4+eeybsBdHrfXnOPOJejV+4dqD3gP9n5ftknR9kTlbDBY57
/UKVKZPyIJnr+r7UdmZJwHaYDwu1x+/BtzDF1oFZN3VVVxs6o5/vKjsBD4vAaWl92+QhlI3Oe54l
Cnqel8L6uhcNMac4jQo/zYJ0gsvJ++G0xTmr9ZZUPGPe51+jgF6wW5utrqSTb4WjPkZGyDnK0XAn
TM1A9OuIxTNUFkVJYY3delkTtpaAzthLNsX2Fs2/GFTkmC16gqZw+SQfP30IRCnUCWbGsw3jCTIt
xPi4x+a5JSb/IAYOv2tI43DijOtTDPm+/31Gf+LcLc0xMK7+F8exHsQeeb58tUdNwE8Tsrw2174N
Q2WNlGhOv0dXukx6UzQRmiOndCuP8sgI5Krr7HWWuz0icizwvqek8e5aSEUR/y71oyg6ITL0T0gU
ijK7vhTGqoQtdr1th9dTwdz/ZseIwedodmt0OKewO0nUYbJ2BzxxOEacZ3J40ZDvivW0oW8egj7A
HTJlkIk6QZb8HwfjoxFXQhqSLx63JMx9l5TeFUoQCvuont1FKFPMn6hPVqh9U6ttTejAfPd1ik47
IT4k2JWPRzvgpLKkMND/GhS9Y1qocxoUDORKQe9bH3J1JZumEG1pyGI/tkAOanuBiJCPUNn/Bjg9
M7zwFUKNE9UPHwq7sDvSZC1l9MDSe9PLBpaS7D8bY8m3nuSMOpFhR3j4e9ez5YuYB8DcrfTkBjOk
/Ut8yWfNJc2MkVh6DHc0Za/7n6JerBY/DISL4Vp4fH4jIAENJV1rwbBWVBYwxFyfQmlM1cUvhFnW
YTY8zWSVEESIIfyw1NOx9ztMrK66c6AUuCv0qCVFDgwIFVu9wGHZzNNDPfwIzBTHnavTZbm1ENK6
82kmK0ZpjVHuoWLGquG8V5QO6meO2iOUudwB/lyYIpRdQUUfyj3M9NA3MgpqBY5St61T3/E3KWYc
6uRO2HwZrekshzSSqDptS6vXD2jPc53wwdb15ag0XzEXRNRr2PhOzGm0+eOzo6eiAXdBmXHyX60N
YHaAALz3CavFGZk9HaOsq7CkxSZom9kBGPfDmoLrRyIO8T5gA6s7wnl1L1O8gveylOPmLdffkFTP
OL11dFWREzuebxbm+yTxfXvxgyoTsNsESMzFWy/WK/opI1euQ1VK14V4HxZkjS+4/DeuBnCRtv5Z
ryRoU72Y7Yj0CRVlCjvnJmSJkF7l7LrjNzqDEX934zzL3Rawn58IN5IpiBufHAndqLZgjaOSEBNf
4FNn0yw/gwk70oA2BOlu8hDIglF4mEB508KrJ7Cz8sRoYlsuKZIQCUnWekaHJ5i7lNui3nmrqhaU
UKkARWqEfIoQr3DxYezQl1hmdF7h8RLYGlUrw6bnKEKT5DIWLrkioh9stnZn5aSNauduHaXO3Ryr
D0gVgr2V5VU/b16j1Vpu+AlgyJG47KcfmMsYByFcbXwEima5vOLLEbmYNMHIBV6TzaYPZ/f+jaQu
QIWdikyTkz+TmrBmuImfWYnQPVb8uYxUq2Z3an4HuzWAfFMvxypDKE8vLMg8lPk9nXPRE0BR0+z+
ydr/LiX9C/imr/KtuHqd1m7Je76FWTLx+VuFVDUT0TpTQH1hkLivJjAmW8BD2rBCxWzNxL3Gdm+j
IVBK04Rg4xfTtWl0X24VvosTjLV6R2rnbsElHdgvkFZmdpNzRtDxm+sTI600ZqZMvzNFEJeMQpjP
pvG1uUeHVYcoKwzu8yS+F/DhfLNJN20aScTB48EAvl3xOdn4eqUapgCEnlj5DgHZGd0aVYjaiV3f
vp3bDgOgM9/xSnU7C9LXq/YpZoXcvNWd5pH1vzK3looEA7MF2N5P0qxCv0X8kdOSPoUEwa8iMX7a
ybGD3Vc5cUX6RC/40MdEMXvnvdQE4p1WqFKQFkkMNQBmQ9w2j5XzARKOSJn2jr45oWxD67Q+Vvsz
c9ZqB19knFFNhvJoqHBbx/XmvWWdPqXjT8L4RceWvAMZuAD1xS1cWH5AATgcPnYTFW61nLwpZFZr
kje/Srp+YVjAALmd+maOFUT7cAgMpHbCLxY7DPoJk+54lboEcfj+HPh5c6xJCxPO9aVu+DE8nktz
XC5FZ8OASuDelqX0NRsndgqfjH5n2P9jVEUrX6rOYwdsiqe91B2Th1bhIY5n5FYecmxfNLJFQUVK
6aUnLK+6++o9PqDXCPEh69RPcuiirBYAUfbsEzvyF/qduyc0QrXbHUCc8lZBaucivPAL9Z2XH+gR
5sEa3njnK61qbbEBSDDn2Ka+jWHxDcNrJVxA3cS0NkSy4cjuTRlkBYbB68NJeX4LHoGEQQPe98x5
6XtCoGMIF0VsCJmHJzdj5iPTD4aWGMv0EWENA/OE0wIP72Dr6SbPqu+TG2rTN6XdzolGyjv/2J6W
uOVorOROwMscGSzZV1zf9i8dfe5GhyLIcsAQKzjZCYrUVCkouBBDBtYW0CqwjDVjiORz6JtLcjmS
1/Lh1Kt3GO3MQmsUY2SE5lf6P2H5AeKVnaKQ6yvPAe02Xsozb0wNLAOirg+dWJhTTlSrAn7g5m9q
BFe79yPP+MROlj4AodEyofmuvLWkLmHLZDAyjkWk3VTZc4kMESVDj/63XpQAEAYhaRqTlJY07zi9
vVfc2boswlPIR/0BO0SG46DxJHA2o4Q7/oTU7nSCtsqTcJ+A9tqO5Bucq+B1Xq19WwXxH8/o2oGW
iqTTRGg6rvUXl1DS7uWMnWbCV2OWPX5OXLex2/bQ9z5mBFtuh1AudA2Hn4CRTOIrrINalb/FqZ3+
+TXgWYGnpFPUFQTSP2HTazKxsSOPxIcsxbXYIrhzoNssnpt2yFrvEEf6TPMrXeN9Oq/VN951ThKt
1YTO0NS5ql4fhkomDxq33o2weQQJGNzarX+Cnzt+Fp5a5MbRocJvGkB9FanSic/xCbwcsGhAzxsR
FPF/ohRcoofv2wNdYDNGj6VYL6P9KSls4ThzWvhZs8oLMKnyGVwyJClqYWxAoPcp1yuk10pnvW0f
nmY59V10SNRGe8q6vzfEjrEMj3fDQWvQj92Eh+f34s2a+EA4uucrNLe+BgNAL0MiHwKTAJZPodzI
3S4qAHYCIQomFTMfiNzR0dIecVE2W8pL3uZyFgp4uLAPPsEvav2Llo868LVE53Cb/8yHXdrMMoEJ
699tNcaO99MWyuIVaoSe5PKtpezrjdtcXolEjIaD7J4WsyNIsYW40MRoR1Gt9+YJ4wC3N8grpe4T
H01LyRtU2RvaKQ08mRbYX9UBrYfkHEg6M+H3ZUy8BKqbkFlnXkFfE/7HEnCa5woVCftM3JbXh+5h
0dNYEKe7OgOjj01qUX5QiiWGAwXI9YzVvxLT93dESewgRyFVhINdH+sH+yTDBYnzCHU9iwuYpzgp
zqGLxm94GSJFg5oeW5u8L4JqDjR0K7p7t1B61GR4rz2VeQB5metsoPXZmoJrNnx1nRH6Pz5wa3K0
0nzu8RiTjlZxGfUq2WGYrl4ZZWsoACLaNr13nj5JHCQUUp45gP3jIVUCRDiUIMZl2G7xAttCDeL2
PYWMli3x96vQ4Xg3y8K//1CZTKCYy16c7hCVGFW70sz0lDTFrsosQJiY0XoqA5FjtH2tk8iEblla
MAmoAYuSfcOwtJK3S8sBXNR6EeXuV/CUNc+cixdyYrdmfuh0qUC7woUQHxZ2tD14mx0JX032vfo5
mZIb0mVywYN5ImkUcOidpzcq8u/We8TLeyCCS2cvLHBHzMTDycojf9tcdZ8U72pWoSsYBQJ2JuLP
NJdVQVAFvcVbi7tL7vL8EAAz/pepsatvTNFSj+0c3f2bOIG12zxYXnQa2/Pi4FdHY+wDDRE6N0Mc
Pl9HQIZU1r9lfsMXSdE5/uN6DFzo3EfiGnrBI7P2sxAbB5G3piiXkXKls7E6F9V3euwWJQDCAmvB
rpc/z8WEPEwgtQePGZxe8eL+SPja7ArYxiSAt0UeEZLccvOWfJW0jys6lMIRAoYOy1re0Xdsxjh6
oEtpYGKI+BCLEcDICQz2vYCR430lw3J2Y17qOnd+95s8slK8c0z1PYDwoBj3bQTNd3zlmNocWZqo
0couYwujHwZfGpM5/H02mURjNDrmXwwGRNMk2D4AvGnD8AXtQWgbVO0+krZcIVG48h7JBp+bwfVu
pON44M36aSuc5UHgUJ6HdRpmTyq575rWo2RvaTh2YSRKiNyT8L3NE8JdTTuiPxZj44yF7w1IYzyp
pMyWkGRPplhhrJso9Iy3fKmWZyBtC3heNHFwFMHLEhmrC/Cf/ef4H1+wICde20A2cLBWGKxj5PTC
AsaQRfnVpZzG3jwMDN0/rsqvCfpGQUjxqLQnQGap39OBD+Kg06R8yGLFJtIVd/GpTO+bs/+Uwp/Y
Y/z/QUJt1N9TCl8tzt41pAc9o6IbsB21nPQxDds82L7A0oPdeIl/7mEe/PgxdayKQGtOnijKB4Eb
9gGcwxesi5XSG9hP1s9h3MAB/3YpShHyk/R89lfWfGF6o6MT/TFMANxNguq2oZo3H2Cj3YjvrXyC
ujG3yUnGYkgR4ItOtP/ZlKZi8r/uIyI+ILFY00Ygf8D/wcYQh1bHlT0/2XanOB/n5YAIrd1wfpge
2DoN7vimoUMJ8X8iW+mHdUkKYmta1TtneQEYQWuuAP9nNfxQ5Lb1rsVtvGE3DZ68zyD+fPL5C76I
Cq8ZfzzQ6QrPvFUqUWs1nDMWWbB6K9b0AvsfAiXmGoOM4247jx1EwWYP8JCl2KSzUgtB5DIeIbrB
YVlqPNG8xj7GvU0hxN0itsZbVNTU7Qdff7KFp2Q8N/ZPpico9Z6r0SrivUb+9KhNKbrWQ6fQUOs1
qc5K4aOwvWg8q+m/3tZ5JTG9AJ1Sq9B0Ax39ohT0RvWc6wQU6vLROLrQ/in86gDt6Jb4F7CIk3nR
hFLPIw1bswRar+lJx/VhJ4WxdKACsKjzWHbJeDGaHvtPb7ZWvM3IrQSwJAhWcixAOvFLFNfvp1aZ
cjZ9Lvh+nrhjgQdzx1p8BHEf9btdmuSjrPU2dTu2qdECtHSZexDynZrAusfFDxx5GSQD5U1wV/zQ
cvKaWOFz2NQ1jJZLl2jT8ID0TkVTUBUQJtTrQz/4PDKw3fH9VXOsNo2L1zo8jQv7T19c1AhCiY09
qkLETQVjXHp+EUjAe6ziEzDW85vO/bqL3RF/OXpN0vEilar8IgmUMamxjlRiCCSvwgC8yYLYRLRq
vuBVz1mAUnoeDd58ic5fRmf4mmzrtQqz+UgbC3PBsHHlWoLHHEuOC/baecFGkUHowrxiiHoUfXEO
e+9YIrfoNqCfsCAtdL+rQZw9tFVcBxnmz+1Qem1p4wjLZR0NMKe78zrdLCuEzGYMGMqvIntFt0nJ
4vXCt89fLZFvk5r5DHybtzG4RllY+zFJXFsGmKpShyiT/SvwCCtGJAWnup/ttlSDonbOKeIcb4CH
9KMmNPHysz5UqpBHNp1K5bFXuEAI+OZvpBOTC3TZDi7aePL2NP1z0Gu1dkzpBQdo1FQa3Buxbh5L
u1U2+Hgzrpan76LWmH6qk98MTyXqqaALhS4XFYmG4tcy1Ry9uMCPxvRyPJUVkCIi7zzRKO1j2dQ5
/3tpoSvY2Fcz09tJ3Z1ZQzC1RFSn2+lW8DUWtUahhmkf7j4ySZNPXPrARkTNigO3ng1WtrKKLRIJ
hl6u+XBr0QtPSHZJU0KuZE9qta8tiGSA5N4jzJMywQKI8xaVi644SfkgEnJ1+9MRGEC8W1BoQfQg
VCJuzCODIDQh9QWSsBjOghGMo+s2E/Hij0YcxMMvGtEwaIXiECPcnBY6CHmtRWhOWQOcw46o/LVO
uxwOndVcxbjVHMJ3tiZy8jh5JKIIVsuDtXkPwNzlSQfNG/IqcP3BxTXJ84U19ZLGNP3FbbuY0rLc
sYtMGWG/IEeY3PRhNy2PRlWkB3xsOjD45ptEnGfJf2u6WjQlb0fR+7By+pasz0+iJT/YYxAI0iQQ
2gCipibLqbKF6xeklm364wc84VxzZo90XqA8yV55ybdMJeLSiMabwvFaRzAIBrfGLZNfeKrbpdA9
06XO6gSOyoNMneeP4EGawaAYFZk1fZ/wkbW+vTEooO+Si5mptXZavPgL9g0HJX+ojkVdRnyyuElT
lM7fPpS0Y0QlT9v7XLrsGtWq6N1i/48gdCaKFsuMAbpAkGwXdfdz+BtSWEqrr7D5xmhHYENm8Ajo
CqW+U6B7pidLKXuArU7A6yoMMyxDo+79USLtr59arGEzKUkNzYUCI86RaIjzAy7F9dNfuQvu+kww
vHFsFo+XIB1byKXZkEE0afAgLh0W9wWIRk3+7qvlIjOgUbq/fXIya7BhowFjlqiQgY2ogr7n3mFA
/DTedj0c3VM8LzPH1e8cckqToadpOi6L+Ae8/cm53aqeLg953+6UHjROQXk/YVnAEtWSuShSolej
oJ8gCfUUPeDQXF0trTpJMNmUXu9cjqfOhp3Hl8HCBg1pFDys/FsgcjzwqrK5mHyDd6iF44E6Bg1f
7XvChDiFoC95RpWlyVqwc93NG0pqjNhS1PbxOQMU30tdY9gPfKnQsM7CCrjFT0E3hock3T3ZcFmT
cFzpzdxQRAzxpAul17udN9kwXcAjtnnYRDY0dzmXexfVnJoXpUAhOmUqASt+MRU3wsLcN4+9Sy7N
J//liPudAfHUnGB1SP9It5v9s2U07hOyuV5ZZiV+sebDDKDvfCLwvmuGsErSyt3brjGubVmrMgPH
RMjQiDDd8Vp+30+e8VNkxjbcPmhRwSgkBAMxlG8VZ8XzVohJVf7Qm5qPPWdKGZtw0lCJeT3MifiB
cnsYWv2w7jvNQwhl+95HRAh6h1oHF8ydrVv2KpWelpj7RZwcSO4P/URVmaUnGp8iRHmrSop6DW2F
e5jyz+g6w9Dku6O+PGtpkUJrUEwaIzyjQFj+Y5E31s3tHDatGGGey49FG/Hga+WNC0GIQGg17oS5
jZmMCPpYDEB2w7MUHarGXeBwLsvGeZ9QKouPDm5atiE48vpKODBP2v0HlYraaWi8vy+XlgrI+6wn
Lk8ittV0bIifwJT6boBjRtbqszza6sg1LVdKghEBvPa0jA2eu2J9eyA3Psq+7dSKkw0rjUY5NgjU
8MzYEvsaWa0Om18C/De1YtZXjtiuOHjgZV8gSh7NREfAAiHQRFmCj1wkxWhM2q9Q4SVEeXzcCz+S
1gE5rxrifpG4CONgTUudzKZNd1Gn0IGzUNgBIpct3RCkPP2fQRyGEMelwcKYkd2h857hki86lXx1
0oC1lFHmyG151LpRg9eqpdtspZN4Jr1kiLRTeZtAgVSSJShnGbdRSPyPZE8CN2Vkn5oO31gOnlqx
BG2H6PQzgnooSfM9iA/V+7y6nZH2j49J/7k3DebrOTh9XHGjKCvVQq7vpbj/fG7DRpUYp+eTKjMG
jEVlaA202754j0PWtVSc1IBUdS166T/1KQpNJ0mojwtP6J1AleAlq8KRX6dLsE367bjZuD3XXBYi
yqiZ5V4fJKG4mTiI7dX+IrjjeZkcCwy+d3NQ7i0f8mQE0tBAYAxlornt/123OLmyUDrjtfKsZVrC
Zd40xcN0GoGYPthSHPCUCfAlCEG88qScCwMZZx6M9ncuaQ6wc92vYyZt0i/RSinuBwYsjJZAELVd
4iCQnO2gCMlkPkAieZ1YNHapjQgE2Dbj6ltwr3Yr8oSSPlQulML7rsTlCfIhG8TUfjdnUBgpL8zE
u437P5xx1KFn6YX6R3rbh/nuEajtAtMClcRPzn1NoV3ePqbYhqlI0/HQp+cawQsYVkDuyEeSXYja
WtZOIQza8peaNA995v05E4fbLeGhsLfApmwgw12KNDfFXCckZwtTXk3hZrYYmWmwJLwarJVJdvGM
XJpHZ/pJEuaHmJQw+LDSfzCV6rUMg5EtYKfljm42wiXH+hhNU2liFULKhmw3peBaqhokMkwV13I+
/TH5PjNFYxIPJOQCNNiAcw2Rz4vSdQdgEZPYEKalw2DJTBfQZlDmgx+cVOBzyq/gemWkvhIk5NMK
eaVNP3aHTLFygQi3iYxRjm7cuSURAk6G8xfvqt5V9UqHAa1pYY4uDDVfvnZHWqT3pVIiWIOgN2Rh
WDnbKS5ekghJUVIw1ZhUf5VfortR988um522qCAUrP7+TDhtZgGYFZPgdg0KOMoepiAZ2FaBlZ3u
PThWxJH14qZTJ0EXcEF8ZSFY4U1WjJbPKPTKjmMPeX/wWC1t6f6SVcuSyoJxX+GNc6e9C08JGF9l
Yd+PxlnpMl+v8hieG5srEAJ/mddF9uyW1Trpa29HqOQB3sQIFtCSFpf0JY7pCRh426tlfF5X+Zkp
4qe4pu0W0SuTM1HxQsIrDC2t//ofb+fqCzgJNMEPTc9+1AdBUtFq/lwjAXT0/gTLCIL0xWwC+tNu
bFbgC4lugewSsalxrL8Q/wMMXThZSUqZAEfFjmtDg6dDWpx0Wcr/xail01Na/YW7V0j5QgUkTK0y
RG/b05ipnO/RJY3dXuHhahBCuF7IE9LBCppt0GGjTnKgid3UvKXDDFvMb6TlNOrXajdNp1VPCWwd
zfL+ooZ+XETgi+9Undc13rpjRd/yOH6PQNFCasJ9pYlP2Vve0wY0Olnin5beoMf0Y6q7SoVpfqHM
Waa+SBnCOEz2vGxPDgf61mfGXqut2Nf1Ec3ajkgc/kiqXyjdEa/NQdK4rdz3jA7MrhEKLDbuF0+h
LXO7maPDWVykkCX+D1NKXOZe74FhvYWP19174Ote4JvUTeFfIGttBU8/0Chl4sc7V1FWNZe0dmyw
jsB6YINq63pCfm0x4ypa2ndex+H1c2DkxUWI/tlQeBROLLmepA6P9hNATgfVYeJaTbmaRMexrHgG
oLhW/sKEdzjMnoU5Np7r7oW0mIWH5rfnWuhM6NojAa7gy/4d67hoNHzq2/DqOQ9jvSeuHUTn74Ls
CaAffOboagbCB+3r2SXogovaQf+xsAZX0DLoZ0J4EgvxLsRorx0nHyYrkn4eQH7CVP2WDXHoaIv0
d59/cpyUCOy0G2oBvpExG0K7MCMJNQM5eYU0GQplQT5vqVJWCDgFZoJfYopV8I+h5jsVYyzNisLG
OH9xNMidvWCUXS0jZfV9/w48hB7EQfgHPl5D2qSDMr5gzaw42pxXfNk4I0HeKedT4uyxg1CyFK4R
C+xh7GlYwAoIehC3ksEXwSlOGm25qobgeFPksFeEgJ0hbBRg/OvOtdWWBxnD0IljhtgsHwmTbSS2
jsNlSHexad54UeVmsOeX7DeK8bfX+Hf0DI8GOx1Ojt3cSIKKvW0ZNzYYcVGvVGgzb66cvQX9zRwX
V72MyX24R7OAns9snuTlYVzCnTeImSLlXOXy8mOHwooLI0Rh9VmzQD4p2anP3LTTqarwLkiGLDZ0
1Zz0lqBoLEGcBy6Rputli0LO3QqS2Mkhb9mZETdQfhpDaKt63O6Yt38tjEbtwUAz/pzdw85CYY0G
KRoSiEpfaeHxbV3RvE6RgXxFI3LYk51ObD/7Es6TF3L6hjRsQv7u4WKqFVuH7jAI4HG/94vqmDkw
HGTgQ6TS8zlYmZECCeULZXl1UmWAs1pxGAPsOtr0yaHraJRb8noavfPoyUq9Q/vilXmfN34jlQAj
Y45DbvRs9qt0PLsX1qVFbZCv1qk3DwglRe7IL7QeUyvY9yYvDp+qUG0wfAwqKoWGuqM4KEwD9ezn
sLO2Q7NPztMlgXCMsdYCdkBc77LPgoRnXM0uU7Jqa4ogkbw/3jkJU1qXd5ZcWXxrghuzVRdngkER
6q9xWHRjJm3x4ZFIyc8n36t4hoYCSukrlcOFBgisVxoTESELJciGVsS+AK3EGIuvSILIx1Y1dyvK
5y195qXjUsvxGuQCsp1xXelbuXnwb/6i1bmNTtGekq++w5mxkqPknZHVcAiFxO2gTUSWnRUcEnXE
1/buqctyP4pA+i6pYpIaxnh0/A+ltRkozevbx3qJJAppq0bxtFhiyCM4x5Q2YV4EhK7GNRY+cwhK
K1JMRugtZtd2jwq4lZOi2r6hiQtV84dqWPRUVM82MZONl1hwL70xKk0lGDdXm/G3orypKIfAy7wq
Fcn4cdFKl0S31jmpOd1Nq2wdbR0SQIbj6MycBIXQHRBx3reesHt4Gf3WbYcliwBvPeD5jAGo3Bum
88Z1xIZJpmpaeTtkpvRTHjTN4jD/BH25i21MShKiSngbXxBZRE6xOWYFdllAkPHfkKih4wbhH/sH
7d2DAsesxG2NyQex75jh4kJaczQWinYc06tBJTBuwcSXVj4qc3fYskaB9pEakuQOlEvGWiCkL0hp
98POAqkB62G1xnoLsaiI6GPorWaiMp6nnqoWo4NAHfmVVrxjMoahvk0lohzV1IwM5J3WX/zOF7hg
Ii1RXzZEq3na5LAyAJCkIVmYqSu1RkMN0vmJaraI1A7jVjfdwa3/ROvjf3OPsVotRpyAF5CwxWyW
iZVE6wInGZJAzdcFDplKgRXM3TIbgEQhh/OLLXviX6c29I4AB9maXNX0WEtbzebjSHPUnMtqBPxP
zak9WQRedjRHotOo1uR7lxToDvJx2VYjCj2JX6inmJi+zDUHUo9lkayeapLSfis0xNBFBWIa9ci8
xWc01tVMXAPwhaoDQoG5ViqO2mpwxPWpt9zPkjKKhHojJo9v2uwtnvR5SB15u01Tt1d3eYJgw+HP
GqzRKt6fbRL7LjeNJGbE0VKdcIbSaeg4BOq1WMstVOI5P0Ra9NB5N9bhEoENVMHVzwYYvpG7wPEv
RzLqBnUyug9VVUrVIjx5SeWqrIvMmFbBC2KFxqzceOlEpEzrIgMjKNLys5zX8+2C1H7H6sH34JAg
k683asrdzQemdc2XUZwJRFUGrS04wdY4JOUrYDBCILV04wEvL4i2JLYvKSYX8EqVOTabLTl/t+wN
kIZLk3RZRN8+x6JBbIZ/RHM9hnCAmEmuXvATuD1bqYtzPfUSrinQsft6IaoAabhZW72ow1hfj791
PjriJGG6TJaESLlVWDXd+9l3PP6o4hGtMMUDlLcfATcZvvdnuG6b++WlsZbh8NQUh0BvdLDAYYnL
ZF3ezpizN2I34fHt4P5b9PfVenzDhJ8HOyEdGGbYAMXhj846kX20DPGXBurczlXJhnQTx+dqNH/b
a/qi3gJ+XYpX8HAr34SiXV7xXrNTRpX1LLZiw/y72pPRELYaWvIVTdqHcTT1yQ4MbKI/YuARxIXT
PCRyv89XhEyziSQ3Zcm7IqClX5nO8WEb6eiiTVwsFo+3g9nXin4mPWQGRAGyjxOxm77eIBAAbrjb
wW5UQuGqDr6KRuDiFJ31DH8flhisk2eI7u8IHAjotGNJ25xlduEJ35Iv72MK3bHRaj/xoPk9ECbC
yJ09QyPorfrnIeVOFHhpwH9aqhThhZ7FPYxVWwxnEosNhP/nbUPj3r06G7itBLS2x06jaAGXpK2F
rBExzCIlmUphdCmkRyPpIKgrp2kgZ8QQvlkFA4bPr7c2sU+L8vfI9R+mHgu4Qg/bV1xxnFE0ASKg
qh+Qbb6NMcTP1ofTtwNXuEWMMVES6NpKLr4zmlhWfvYxHEzOQ/RYRlljG11quAPGRBS+rtsKTNan
TCCG/k+Y6bUOC5whcA7lFpDFkGfNUxY15rq9uIhiYunbSQuux+59RJs3os47rTRcWW841Z/xqxNH
PHTl9KkYynwtlMS8k5Fm0C/nX+h4bWZC3DN/frfCTSxHLSuM69MFPnmTdGSO2TyU6kQ2nPL19CKh
HNykzEmxpDxGqrnMwYOJzEhrgoXV5EB2Je0GOUaNCjNH6Hnz1SM1xaPxSDYvafVsWE/MXNpG/B0H
CH4JFztrrMdRb48JzQQNPwYAjyXT/OGSJRvRo8LcB8FpCOutrEVJD0f0MI/1/PtAv4aa2xRg7CHD
hc/5rjJtwEhDwafrGvD/o1yQ/6k9pp2X/Eahku28wyudMQQNIOILWBI5aiWSFKXldwgTyGCIa5Cj
vKYzag1fXwSEYH1pgh1TsiUq83F0A4X5wruWQHxphSOI+pJEReIDXn3JFZrCxTg379qLotFbKJ5N
Vklh/ufUdhOQrIFK/KZXBXUrG+gqFJtsMuIF0O1kkbcijBZg/Y5HPz6QnavxSYTgDjNlRt/ynLYY
/g7t4MQuPJ4gx6v0Y/GFdw6gplj+52laVFWO3KjidenTu8nx5fZKT56QdXXM3GUtSt0mGlnKoczF
lDtoYYOgoVw/lXC8Mn9OhcBaV1S3XsUTCVcVb98D6HxGbQ/v3HFMboYNyDyEutUsIcwOl0du9fs6
w2NwhX+J3jYxGPpeKrcA4hKFGAQ6T03OtSeoENGbuj5pcQFpV1zH+cnEInXNEXNGy73o9I/nBYVO
0z1vCJdLZoa0hSNuKXmuDn2MNIj6lTE6qROcUmXubRJ0wMl3v5C7xHsaxo+ZsCAg754KlTWmXwg4
P7Bi6WZJ131yG2i5GyEsX++mL2iRjpxQJVX8+YXcKTo65KL8GZ6LL3g/FkoNJ4k7WDGM/Xsxv8Oi
8iXB8oM7MAnx0ma6pHoWRTpPaWNin0WIY3uo/aHi6rJdCvJVDIypaLWmC9cKnREgUyfPq9dOaJdX
+LvdOH4NpdKhIZvOo+/JP3pAlZ+sNIMCKeQVXb9Z9yLG81zNN3P+mjWfwp8YSXtCITkLOgmMFxLM
xXMXPwg6AelwKi1sr6uokj91HhDfQtvbG7lLvP3kU9EesE+Fn9D3G2hzG9WI5t+M3k1Z9WyAn64/
LbyLGZ8vuecD/3fyGB1CMdTkWG0zq3LAoDkD9BPlys0pved9UADlc9sPA3aTDoBzVSPm55zSWINL
kHSRVPqdwj9BeCOw1vnlKFsjuhYdKkpvaYJj5YQqQAWcjP/RNWOepVE5Q2YwDZggpkLg6KRXf4KD
pYQ9j1eFk4xokUvbmWC5+DsuBv1zXxdkMma5UfewYukZIgOOzzOZxe8gWELJlmNfpQMIz38FNenX
CYYYG9+jb0SJ2MGpGiBp86W5alpzUJAwXdtfjEvgg8rXQ5yZDvp9k49i/V6RRww7QDhbYqhuBIAG
5UmTV8wuDKsuPxzRNlKDuJAeADIdDKkNAhI0xkE1k+xXEB1iUDbcJTNrM4RpqeaH+K52jT2RSU2S
eseinOUOAEWI/3QGIzJFXZlqe9FfoL4jk/yps3cJjO92YQmjTotSnC54pFA28NekVMo7chWLhMuo
eXK6uYSCne5Wt+MptIiDI690rN5mUTS3r1Sg9iwUJhHtYy0nO+ALe5tk9cDpI7LRTcf/C+bloj2D
bgGO8dgdcaSdCPbczqE7+5NlXLtQPzvzqDtrWC4apl4QJJAcBFsq8kmCqOTdmVfx3wKD8qohdOiK
gkX3HGaJuCKxV1PX5sd//qkAvkcKKztmVoGgnKZ7nONoxmgwKuJqtR6yTc4BMKXPBmMQjNMmK9XM
lZHLJbGptKfthLAANW73LvfYMx7NyIqlHlvUFmKQ/ovUy3r6cGs4G3om8lRJH4zxq19Z47iBDa9T
qshAwfUO5PIEjEIBisbgqXUz3ZqzLbjENnY6s3y2yoiLIKhNR1/HeTTZD659EcVxh002CzI2LV6X
KhKvdmlyvXLKGcprUlOWe27Xho+Ruj5g/13gP4isLnWN3DwvvLaXzx89TrMtJIwyzmt0gVurmgxd
BViFniMoZOLMLlNMkH1d10wOxB9MvCfDPuBLsx7BCWCO+G8G+qT+jczdCSQW/F++yEcsRIyadfrL
YWrT6RdlHqaTgRddoZc8QBwf0Odh5Fy450w1FU8iqtE3rRNLZeFnJtHBhtldZ2EgiEiN8p3/MW1V
wt6hNxsjpJ5KAJk07ej52EvrqBJ2RlTFdNrJA+Q5B38aYqvXAqqH3esdzw9qN0xhVfjx5bPc0O06
8i6m7s95c2hQ9GTUfVBY+i4e22EhZlsr7FhEuWZMofgbBtUFDG1OvXrlLXIIvoKWb0vyBH/Dm6N7
nAh9JMp4BVZBG77kIKK5/fKDVIV7tKBhu85Dn7IVHmebtZcVEGUgt5BG0knNBx0BQPdBtoN/lsYp
5zBVs79zJ8ZL5APpcxpjObWdV++XaeTIf8Rm/0UXNbrtNmc0OAg6RMu0/OjUo0BChbAs25XRG2sV
7SzoCopMzS5ZOk/TPmN5y1bRkJkSR5flbHD8q/lsso0TZ0q/qs1HBCvuDt5UBYxu21pBc27FFPiz
TqmC7Y/ZsoKSkViWvOg26f0z1kN8Zgz++QdRpbrDTveObutHzKCYxpMxX3S3dWZT0xvIBxmxKKg6
Ggh7pIAJN/5+CIeahJB0mSG5wdNt2AS21PFOV9CgBdlWd/lNiPvedaPxpvXkEZJhcPket0XnAdFw
6Wx8Y073uEu/+F3C23IWCgx2nBqBwow8O2iT8niwA3vrEyAzt+Cn/H5opGNhDXqvhL2DLfiwe5Dm
4lnlZdvY3hy3DwWyqsdaHJBhLnxA/LuMRMXdiMz5H5m3K0fNFoestS2pXiauaAl51ZA9JXmznE4T
YislLhMot6Uq6YOTq7OjjumLlGJROypKSPeeQ3m53/A8DpwNo0v6KFffghZ60m9Z+osoz0K0cnCo
9dYQuCeOalSsMBbZtuMK4qZr26iJmmK30eleU67YVHssi9eWcetcg5KoQ7/DWa7GRKYMqznTwSeE
cAo5paqeBpAegRjKYpteC67G9SAoaNrk/QeeSYZba67yQaNuKjWbyLzJdVjCLDZlhPFNzdw7Ip5W
fyENwuczo1N0b2u2GELMTQN44SfUrwldz7jQg35D7GindIq1TBFNgDFzAgYJBkv6iR0QUqxd8rcJ
l3dFpvvyzi0OV0JSz91h9lrYJ0bKEUEXA5eTz1c6VxOnJOjzv9osuQY+OkC9x/pJ/i5mrEBp+JPI
eVjlP5Any0je2DPhvzshWlE4C7fwpI7Qku4TCIWlXXAm0QBmhYemO3cVVmuveYABDzpGN/Vjbg17
0fiYdm0rOmjNYjL94AftQQ4Ugn/EYWASusNXTHM0+W/EwHlNtJiQi2ledlxlbhz5wYby/eHX5mhV
VPgqi1/00gYJmJhd6LNmmvncV7gQL/SVqKspYNcYyZAoxalXvHQaFH86ErP6tNFO95Dy2DWCifpX
fQ+G1Ve4Tvq4RZXf3C9iAe+cH/D1svyyZc/tfMQ+ycaOwY8GpNqPxZk27XIECOX/qIIgmnNMTnR8
jK+0GmZJ1H4FxY5+c98+hkAEXOdlf+kdcGQBkXLCCRCdmQf1jPTs9t5DmO6gmR/Hul454gHIF9zq
vrQ7Rk51PkgsdU2VSwDQygRMIXyKJ79f79gpwQFxTY2oOIOwfMi9dmpLFmyf/yZYCMm5CIOghNKo
EQX7S2YQ+TVh4+i1fF6rwK+3GQkFEr+E8TtKSRAcww06jfL9ILyP1YRGx0tFEP6Plcj5FeRNtF7e
4/9hnf6N/ZEzZ5wbUFQFxH+lE6jd67HSbZm6tHSHyp3Kk/T0hmN/4D3CAgKwSmhq+womySO+DV6W
qZ+KXfNWdop7DxQlzmSqMzr+Ez0X6RFT8g3iA4SP1qs+npEichZR+pArIolmdJJxdD7e1OwLb8VJ
xvPGmmzDz9YIZ1s4hBr9qn9fv8YqxLEO7HjCEFAOgGVDeaU8mdqBaipttJqkN6/ffp8+ZAi1RVIX
KQIhkLthNrGnCHbliHffyQZK+jTqwlRYbXQCAaKCVWVrvd/zO/Smnb2KVgYVam0bWf/RAcfxxe3z
I5g2aBc6PjCjH9/Ne80nxOdxdbTHwgSSw0dtXfEvOCjXj5cBwPkTY8R3j7yEXpNbk/2047zN5CWV
hy20vM4+YsC3gxJ4QQMCBVLjDFzaUw4ewJppnJ14Ufgyhz4FC50LX0Aa/GEg4H3FVuECVVRUzG3D
vqLk5Ue4ZRJFblTLBkrvFSHB6Ce+X3rqv/0euJBSU9RCmjxIvz7+b1zH3lwLLdjy+ojOYbfYgNFB
wDZ195ZEqG6gCy8SAaj7LqMfwNq+6QzhpPm1A4eMnvhPtvBWUhP6sw63b9jgpyJ0P4JAmyvUNXPa
LoX9jzERWPX5Jvj5mWoLrV9CVw2p57RDW2r3RruYS/vcbJ41DDxgNb8Fy++nrid3AL9YknY9menZ
qaHdyZ5kshxfObKERkVciUHjdyzzaMrmDVubZBf9okSB0FwBWCb+ieKHrubkNFEe739teAtfSYvr
S4JqPGaTbKdTRKmSbGqnIaBnn7YzgEdBlqEam6O4NBtq2DSG3NO/RxiExxGfkrY6xaOCdqcDTpCZ
YNojRRWjRDuBfnuLDHx3wB2hYe8ruz2nOl0MGD3JN4lXJYipB5NyAZOJObFayVmW0eLDIt5XMn+8
si60CSGPccexVB/Jez3Zdu7UvJOQ9IOw125b37HsgJgnu2WhTdHUo4rSdk6US0c9ZP92/OL60dsC
43P3GFD9b7EwbjAD2C6ic3/Pn4ZKKXQ6t7S+0nVqvTp+f6tlDwM65AHxNgmp5QKP+3kQlaiFV5ub
3PzIUQb+aFhb9i/X1O3aoShTrrpZvS0IeWtnu+JzjFsFyzbjZKopfhzgcxlt1Pxt6AxVwUzRY0QK
AONG8eW5B8K4nY3bxwiDOfweOFLPkEKvM09pjWFISI4aBC+gbw9APcQ5rz/4NPzmu0wPWmCUTKvb
1MTNL6JTokwZGhg0GX24EFnklUQv4B5Y/o8Z9LKwJ4axWVQaZiD21ZqLj33YuI/zTouEFl5H3QkD
UOinCyisV34SMdZWR40/TyD5K/mTzMvocxBUWh2ANGXLiQ9OOwQ8m2+Ql5iN1QV09l2JGXNcUzSb
6wzx585t2bYP5kKYr+IJNnjN+6vchYdZTgardE0WbGaAz3rkbASFwsl+Kfpk9SJT8N4aUdSE0ZsF
dsp+Q1BEbL1WDH/ucG7V51YAy+XyRinkh3ubfFeraXTF5U6sWPt5fkwwuyP6v6Kw9g3fphOc5nEc
RmtDOA4quFf4oeHEtW2q9gs5cFSFaPMb10rLJuSy5BZ3eR81fxwj4pnx9EIXZX5Pt7mhUUFUDMAl
qUZgwDQVo3+eL5ITM+T5b98vBZJ9qThvBkzMziDOBzovfJnHIlPHKpkNyorC8pBYc26tpm0rNIYN
Q7RFCw1f0JgwgnL1ZSXVkKYF2Dayh26Y6qYwgjcpdDzmPd5eA9hhNX8NO9mUU38vDTA0Gd6/mBv+
ZX9MP+fz6gsZ8jJzzRRVj8r/NQnUIlH0p5g3OKi2KjVkgLZDwok+WNedClIZFiqIDkNgKA5wyg2v
4OsM58u9BuLyj5PsGIvsa+bmfBjZZB4r13l0OmnmGVfN+zinJtciKiElYedFoGUaJGhmOpZjik3R
+jwkOV9nmgilcyKI5EJEfb4ZV5MEKzqaGpwGOGLhkLujFuyVhHDfQg3Ds06G0jr0k63Gr/JBHQ/9
05lwM1CAIx74m23ACihoTDrgHabwO6QEDcNE8wmdTjpmQnGxiKx5JlmKvtWyrX9tZW3sjGQgX1Gd
CSoaH63bbxAwbSACSkM2rY2Lh2/mcrPOBK15egVQLw86mJVI82gijFIlOEWj1IMKR54J1BsI5vd8
xS8Hf8FXuc6Vk+Qvms3rVFfKcGqfYQbPZO3xZ2aDuTQBHtBkAtfg/CzphFRIaYH7EOukybUORcAn
GXlL7OKlmxhH75fTSBrgw31FZ0b58ZMjLpPywUEBP1lfP9sZZo9SYqH04PPbtG0HGjRZREJD4jQb
OA2P7jjxndnxe3BlW39rDDQLzpg1nMPaHQIjaB/GTL08qAH/RXd/ZVmXF7X3reqwVlYPy7Qnw/Oo
XAjueRwdFgX0nYkDLYq37VZUc5vkb/JblPsgAW+UJSZUuPTy9R1cgRr4VzZiYKEQ0A0gTICX2XSO
n6kNaVHC6Hw/8FrFAIQP2Oqsv/d0yTz90SL+QHfiTMSZziLpTzKdNtK4L4zqKaRPF1hvMfiWFlmT
3613LqpzGHzvngVI1k8gxKrftofU5TAqt8NXP5wkl3w3OPmX3EWFWzAmVU+QVlMMMXRVV5ntSMC9
oAnEG/Hk9Diu0PtoXT8O3vCL8bAlSQOKzRheHevtiEQ7VsLmPUssTC+1FR2jFLzJFrUl2nz0k8aw
CHKUacKSfhJEUjz/zoeoqtggNHviDsDk3DxSv19HimHIUHdFp0oidOuIOrIzA1akpSiqYNMXGn1H
8frkpriO/8YgQIoEpMsDgSZ41FKyud3UDJdtpUgscIxkRhP3L7QmV2ODKU8WzxKVPosNQyPoN6dX
4K4i4ugvkdfXgeqHjgWzRyB3etCchvZP1rF+Zvz13rgkl4oF3qnFUuAf9wxJzcxpVt2Oq9ZlKDZv
3EwBEKAhg1PWGI454Tc+Igq/VboU5zKtD1I0T81MNxr9nI+ksAJ1IijpZq2Kh3bRwtKWr15slfq4
d9dnas3e8KpiKtmoc968pv2bUXMK3pANvjiKRQ/9/pujfXT3MUSGgjp3zRggaEOoYGNclp+/IrcL
I4knEQS+6VY8JRf4ONhMBSMDrFlpZpLvxW1dxYm3E0ij7mu+5mj9B/RrPOljAdgi7f4DWLgWRind
qal1pGkD6MYHWdn7/nCX/eT6+zSf8OttD/3rSwzQ8AzV7erdw6Lq1hXO5/HwOwHyGuyLVxyJ0eEg
cbse42nk0Q5qwSqW/DKFErpNuolAuv33uuAOqQzLr24BaSezbQaSF9GLL19sgDHiLHeo4kn2rYeh
K8q7Cb5mvUF7kb/Ff3wKSNOqgSyTsyWj7e1JmLrnK3F9vs7kUkFSRMJqtj9Urbbd2MnsE8GuVx+P
OkqTMaayMj8AG/Sc8/wJUgjl/p8ttsm4OaYTAkE31p2Mo0h2NT3Va5Eae4qColskz4WKwQJzZRkK
OPZZU7NuzWkBvuiZU38d2ksqHaBTXzjvwN/dRwpASKs7vdk7yVwQpNfboGDfjaL2mPDm1A6y9Lc0
YTZhtpYxDhOmsyk0xS0AdKlvW6wnRrcbYSKXKREbjbJr+qU6FAcLMxHRVkiv/VsweN9BLhik3wVC
p2EY2juIuYT7siIUOW4vNsSSSmpFUdg7d/knRdWMdKVFfyOZiwpSy1UoMwpPGjifHh5rmvXsEpAs
Kl9CXHk7nD3YZow/rGqtXAQHkr04M0gZQKVQXXNKasECIzVeb9eHWNk6pmMbilm9PEoFKOE1zZb5
Cri51QbD9FnxMsemFy5JC2TyZ2PDzSHdBQONqd7tQVp881McxdkzLDKQ0YqyrosQvbPeYquEtLZV
EA3sPUIW0HEBVUlZJwgT1HJfu5VGW2LkVPIotp0EONPvoL/dK3V/kCli82s7HFFhByJXdYHJoAi4
FLAnqPp99LrPTWVX+7JTqHvb2Wy6A99TULLh4ipz5tFXPSJQRDVhKTrJzYlPqjYF0LJnx02fmYqL
p69+n58C23af6dDpCnwEnxfn6bzpIbbovlCAmhs35f3+b+LSxmujDjXvnlOAZ8g9GZ0NbvVuiprV
TxzaaVnK8lVw3NIGsATXaOK1o/ji8wnOcGeqgJBf33En0wsl7R0C0BiplN4KeyRx/w0xYi7ap8kE
X0XUxk2yA3nQwGzUwrGhgZkBQA1yU6meyY++DEKflvea4/Rd1jSLdyWwyBsfI7oJP45TqcJu54st
/A39w3yA7z0kVW7MZNqXdO1RCVVLvtQWL94Oeb42c1QSQXcFOzrkk4NApWlUg94oiu+MMCB0RC4e
t+qFx0s+Z3Xxsk4RS14ZudnU1gkJCc+RDlZW8hZsyviICNLMATtS+y4eMzAjqZBZFTgAWbHfgFui
E1rFRRgL1wHDlisJLuZrkVbT3qIdbvOfETcqGVdi+9vfCvT+ltRVrHZuoczibKsYKzDKD2sTTJiJ
/wru35j//+fKqUr9ONq+yW7dUvZKNSIzcHk+wEECdWE1Fi2gvqhczTDa0Vg3WVE6oPhqqzaxEH9q
tEuoGuSpw3dEjjyfb5oQr1tp5XjGzkIDeBthRQk+nGSXybdVbS2j6248XoypH8+/CJwA3a1UxZOS
4+0chnSjjyNvjJgO3s4qzfiGGEuLdd8qIaZkgpsSqR4bmHfw594F3UfVLagFHrWBZWhVhHFR4Asg
LaqqGuDS4VU4sBzSM/qz8WEwbB6Ci0YPMdeXmKcNdelnjbACyRTpUFX510akDad0m7JTIbKqxc3C
2rHtlsrXYLCzV4DG/IOHHCfPJnVtm93Qw6xg+J7InXCzaPUI7yRQSUJJtOcRlz6iWC0oVaY+Y4o7
HbIEsDlphMNbrvx0T8xVcjNC32VfsHV02di8MOV3bev0aEjlRhHLMbSsIEMXq0hgw+yVQbNmVCaG
fV3zYbnzAZ8UjS6MLtvlW2oSgp7fw7etBOIM7+xZ+QmfkK35STe4psu7VAiIaVuFrC+k3OngSZAM
HX9iNxgwbv8DUK/jkzeBB4uYujU3ZfeoCheFatLFAPMsMwF3oxa8N0KaSsCfwKj71wgTCuO9HrCe
Yeooh/SwDzsNT5lBNvjHjkJPNov8tj9XTzSNamdJelOkFV6m1jLS6z5UHRleCVPeoptux+43rPOg
/yBZXbHQiym0lQPfgUoxj0SFd2zw5z7q+89Xq1UUT/hg5fbD5eBWbF+T8/TItgzOQJm2YQzqYUin
VCWYurO6zMyk30UPlELyAQ1/XB1/MrnGr6WkxeonX/p+rnLLU0pHii32BPScrwDFWfcTi+bTtknA
5ppPdQ62L0bULENaxeFu+/tWXNGGzu8KZlC030hOF3XIhRJWz1yxEjKBpEgQ1te+/HtOBKSo4h4g
63ES76IcPVaUyeCMs0+u4MDq0Zs4cS6l+cAqBrsFH788rXgD0lKILe8G48Kz/L5jzbL4dB8K1/GQ
I5Bl5kd9XQD87XzohpMrRD8Pw29euXhdtkTDnkhhUhSm9V3OI5hhAFiWhWheN2XvCda9IIQOkELd
R5C/RbAcKhC21mInbN94XbocBISGmqOAHE3O3SRtfc+WXJgINxXCf8i+wC/ixXrH4uqE62SKxvwO
cS1kqHyZuQii6bEBreUu6F5yuXcw3Vzmgrp8q4rEdfNDz9sqQZgTgjMWfTwkTNSdiSBXHLBSSDFq
GHJKZS2xtgEP9y9b4hYnqdZcdkHg6ndB/bHcN6/EcVoIoKbDok8QkFYd/+MncE6U9lipFG93/g0o
ZkyIXMW7bBr1ncEK8joNVk38iqXaM6vq0dmjE7BJ4DqfnAGpmlRGLjYhVx/ZRm5ktuTRu3Y8chta
8vDFkqxQSlTnOjydamNH0gExezy+Hd6cJbpjsBMjim5oIG3to/SmagyjzePiX3/zfhehOmPk41sj
slfZ10CJRUIwLE9P5Mm5YF/LjULA5QgsupYV+FIHJE0uotZ3NGg6N1w3TRdQP5eMofc/OYfuiHND
/+L70l3B+DpIpFztBSdTiufkNtuM0mYzIDZHdpKGBaAUQD68OM2ITBH2VmZqb9aUPkdNbvtopc0U
S3I3mXJYT0/aWf2jYoP5+GJv2JV+LSB8VZTzAV4JXkiGmHBTRVwylW0nndA19Wx8VOrdXSMU/nKs
1rLjinP+FWvbnL8zCi0AoSQg7KMviurAH5CjhVn4lR5kUFXk9G+W/ez3jTeMUNuSph19m5R4dkIr
676AicG9OlrB9WWynxjrrvDjwA98TwS4u9nt2xBzBHGDDj+6ihjRn5ue7llCKwM6m68jSpjNUm/g
2cqZMZ6wbC1xEPaye9GwByPXdQgPd/YIx01focMbVyZz8DLkcGdMEng3mlN3IrHpE/6IBB4KNvO/
Mi2fqADkIVf1V/X6s53v2BTcFljLUy6QPlIRbm6UKDcamaz5B3tD+ofUUkpyFaq5u0F0C0UHVvcU
NpBK5ZnUsKj0bHDebFZaRzUSSAojKUj8N1VwpR5MqG72Gws2AjOX/GVPqXqH9fyznRVNepIFeXip
sdRZ675hDB9eFGejIhVla1scTimdwAhQhPM4Vhq+jgSeISipDUh0wJ+cuP46EW7LmjTyoAsaEbpE
8Sg5RJsrdQ6NmaVKTJW0tiej8go0P3eG2XAgI7pYUo3xOsQ60cjZSU6TdysAOugLFcA3kNJRplAQ
/yymDrSXXWlZC5ooK4AyNDPn6OKHkBDRB+phJ35YRSJd9xM2jkD74gMHeui8dxXkcGDD9FvojRlM
nHs4kwndjk1DLvu1Y8by5VBTMcYaKqxga2iWbEEel8qlLCChzokvqdMMrbc//K2rqffaKRQiquSM
slidrHwJRUrC7yQE3nJoqsYpBiKICQYt9Onu1ty6PTqM2SrIcuRMJb7k+IidDz5dVneiH49ewJyR
Mq6lFE/cJ6zdVUnyvzCgGiQwlqu8o5mkkR/3CfGSgbtYUF7qZaDxZZtytpW+cH1wSQm6w6pFMfx6
0R4A/CTLNTR2D3zgBP1KhxojGeb6I9cLHUWw2CudwCp5IsWU0Y1WAVlqeuF7gZQtzroH2UIvs9UB
1h5/eyLR8+ortNAkbJ+sjCH9IgeCh+DUKf/bv1Dnj36XVU9ZwiBBfVoFZ8WFPXT+fImFrCwRvzoA
0YvNVowEt1UVULuHvTOWrIzlBtSTLE8KSK6ZGppbnR4M/JIir6ApdOj7J7BtDpm94xDgUP72G8mq
OctPaTLhe6HoR2UZo98b0gZc095Dvgjvr+29t9ORnS/iXegabMuvYHmLX6ViiIGdVchrg7+PNaYb
LSz+HS2HheLYAFWtK+1e88MjChgODIzupW8haDLctJgSYVcaHKxX8Df+kn7dUzGdmQ1i50VHA6hY
bRYHR2yBCwuvdcFecv4jhNRupgMVj8LmZ7P374WmfMo/dCo/j/OPP1vZuE52SO++bl9rLId+8O7p
p+/f4UQtGeQtszvh5V+90qOuk40FgoPp/6X/oLMC6kSmROGon6lzn3mA05ZTBvwoEhTrB5CIHemW
gLfpZqcc9zShVSglNOKC6pYxFDxmtsjp22bO1rzgHseTsjtBSvlLLJUgebiFBWgq8sGoGZ2krjDp
Q9yog2AFTXYuB0W8NKdmat+HhFYYewftztiZK/P5P1bydSYp+ov9j29szTOVt7lmOXwAJVAq5qGj
tAP5KBVkGRkfY3BlL3tS+/1W9IktrfUtRCaDmrPitBdk4R68W8lAP4GjFo+P/4Krdt+KGs3lF9Dj
LNa2XWzW9ISKtt09594/MPtZq+reCrCDuTKg/e4wXGQpG6GgK9mv0hVwzG9l9/4GfloDAPKSgskl
Hd8mWBQ2j4zpze9kLxvKmpGmc1tM5zihF/WUJI46K9Fc1Ng2pKRqHpU40LpqUzxtSDv8wYlcN6U5
idNWP4i9Mo+T64KnVvohOenhdxyNiAO6iyPdDGBrvozNg92wrI2XJkLttMqutF+xFZBOX9jEbCui
P7cX4zVwb/nAaM+6On2j1ztuU4mdE6COEcX4eDjh/chU+M9atRvg8LHzY18oZZ10HOiBWHs6DZw6
C5JyY4gBPF8qN/U0OPYEwXiDwXKQwrmOWS5Tjc699fFMMvzshDodM5cGOZKdky1dOYo4fAeNPTXz
+FDjMxQoTTJS7dZsDANRY8xmWkKHywABct8+tL23hu2PRPdKnZhSMpj4AQhNdj2dFrD//WG+Vbnn
Ui+pglGPye5m2evg47A7dIFJCh5bsHWvD+qtv2PpQAaEiKVoW8AzfRI24EOF8PeJiIfSJ45xhAXT
LXZ/uA5mX5GOMIyw9Ar3K3CyGOFnwBqAp7b08X8THY4kvkL9mTnWrk9epAYEcr9mN2q4cM3+ndSq
uaIuaQFPY5X2eJhztL3M7wtDjdZMVimuuls48h+kgG+rGJeM3p5KKuO5+c0kkHOH3p40AwzCT7M5
hdPP17TgsacvJ0eDYNIzWyjHmrcIYEco62CNZ7eCo7DSo1GcQu3Yc4ZTGZ4QE6RquV6dNOTj6DS+
etcbY4w7nIg26t/n6/h/xWAR0G8zS8jyTkhWYH7tFQnGQy8ICZf3kRZcQuxPiHYMqg66pMqTXM0u
jtbvZIZR5DI9eae1smRX557bU/Itrh4TpWq3KSYFiwv6VY+LI6gdKtZy9PGMKP+p8FDfBOTRmXBi
KzlG8203K89+wUhHG4bebabOYJrflcsi1CW3OtJq/zy4+hB+aIfXI7rdIhF5XxMYOuSk9RMhpdWT
aFWmAH625nOpyBhxgMWRm1yKeKWXtB5+2BdICG476db5ZuYoalJgVQvp3ginggJ82M7g2n3/418o
QbkP1ZxNHO+UeMuoGECFTeYJRQE/oRjkI3ZLlcLUgf4sdf5OKlESeNDCTJy5Pl5MJlY8uxCBDQXv
oquoW+DAL+4g+ByC3tsMEUlWvVq73vCjiQ2p2D9LBSkVZecPgL0iSl21eiVUMO65tfNflSYLZYQY
+gnjXUTbaCk/8htlJf9DMYxiPEJb3zHMzOevSP+wbZMUYf9IoqrCEFPx3liV4ycLDr1yd9mk/TwH
hNqk/MMjEX26LctFPmvJ0ScwAyNCwNrsbObNXXp2u89htt0wxwhx89O/zLuQV8p8odkPrt0SGB15
CGKVVeAJy0ihr8/e4fJPUmZkli5LQYGf+1DFUTpQQFSrbmRkqZyVRn/7L2Cy7glkM3AiqiZtF98E
rkm8pmT28Fc25Ep+i3+vzqmE7gRT9TgStx+tiQakFRzGW+D5D0dI3ZO0iO7+tJex1JrVM23743oZ
hFWJV8eUvCL88FK2i4cDOMiWtcU2Zr+hL39fKV4WlE/i+BwSFhxLY+0MepP9fIcuFp2QscDIzsIb
97bdo5hbVCSHT5dUkvvK28ILAJ0gf3TXHT/FiClwZoKpkDCmBbVgdJJ++H7Ofw47gSoqvIfLgnpj
WaX6qGIZxXM/RN9rtHSkvUGnaiHNOShk+L7WTcvgXOYLoNpJQAi08Ad4Wb3wlEQAAg/DQCdTkkiE
zpLeL/2azO+g2on9Ni4g2L8zozSHgVDaK1Gr2D3Cfg/jpP7vfJBzJjwj1FsIrDDtGmogXbMD28Iu
b8cdpduK5BxJLg4i3ixUR8Kri0hQWwKrTFkBR6WksF/PDiqPIREK8aUSdwa/XupDM9pc/RjhHKqc
3NKxjr/alqsmNZDBb6ykN5WGyxRNlIGgqJT9PzU2a1RuHjoUamxgB6/5lOoR5pfr6pljYou5vguC
mDVABBLesX4Nw5auy/yPotuWRM59ADnZiLEUgjl7uvqTvBJh+jnhaxJc7Gwz85OI+gNTTzt6e1jL
IUNmRtlHNiWa8vviVRVVYDO65wf5yoDXeeWL92COFWhqow6zLdG2cvxUiMDaH+bxbXZQzhOqPOj2
1AKmGjT7ZTqKk/KU7zoDlQKpIyudPfnp/lKCfyGdACDYZfDrP4HMFU1I6wzsykQRHNXfLUyDCnyW
E0fT3pYQ0MLP7jysRAeX3EReLx/m5QEUVvtuVjsDTjIHuYOs2NyqpW01LIp0104s1/6Veg34cJqt
ew8Z+v6NH2IAeYacVIix4sZnRVzc+qok6+a5laoLPqS7VaBtE9soKKvsQ6vji8wrpxifhOhJsT5j
MSkwy6Y5/1u21q9/t9FkxD3FTaFXZ/kpSC3gGJcMpJ4ERWUJ9f/d0lOMPm6nrJJt6Vrwo9QXITru
/2w38HZqhYGZzSmGUPU4tNQT5wBZVQ7vFXRm3c/eEoG1unihg1NFOtrJUR35B1gFoicbNzIgELXL
yo957jVsyc08RFxedXaCeunJVu+0a4xKwtx0r8OPSFgkHbsoOtLaTp33nTEt3eEu0SIexUPFuAmL
iPmgMRN5vi7ea2wOjWQoAMCLZC5b0qFm9CW+9XV8DNIYV+xiJ9ftItjpocsUbCKPrO8WYKdTd/LE
F3Mu/zod06Bq3t5UYuHBuoohe7/SZ++WVSYXGATgCb78iTJ7DtvRpqdnhzJ/+SlgUww6d8ZejucO
9jo0fFp0DBKTWoFmBRt6r372yI1aOdupVLAHZ7AL6enb7GBUWM1Tde6PT6ziolkSXn17IvqQnJpu
+k2xECZtk6TG9AxI+jpjAmW5lfUef0k5SgowaxNtZEtEAAI9VqmdvO+dbUby/KeVn61uBizjGLOt
C9KOvJbHxSyq8GK9JRDC8FRfj/T5MAzvevnWzvJDA8oGHhStTeDpSKjKGSSmPpx2+7QJmcE0uGjZ
ZvN3BPENZlRkCoCvlzorV2FyHbGnTuNl/0MOslLwHpk24qOqBRmaugl3hQ6XqTZz3TBJINLKa1RI
TWxN2XnMGqbcHPN3JWneR6FCotKpkmU2VnSwG/oBmRQvEDUcONPEgSAnra9BDq+YUmEeNbOy19Cu
wdl1phkfAOZRIxF4/wQwYeNu2JoU+tbjJBqt8R5Re9wBygF1h6/+Ften9IDjVmEZt9jCzt3OqILR
dKuoC5atutLcML1R/bWSTxfbmyzjbj0+/IK4qocGjaRAaa6HAKfZCfFdzPQLaWLCuW9C7fvWTak5
/qaT/xOqxi+8xpuGLp1nU7OMf++vzoq7DJf+Q2QppNh316Qzh9+HikmDfDbtbb3VxCZ+ATUGmXS7
hlzutoXbwPzooynrKFhzy7Azzzvz8cbay1v2JWfLeVJFm7IBY8NxSZqYx6j6wk1oz5x3SXA01PPh
T6diMiPq+EyetVihlyRzHhsBVX3TPH8cTrqo2d+qk0/WZkKsV70KhEh+T+4VDEu74AzUOm8eUe2U
dV2CfwxhZ8V93Jh7Mz1EJOH0n69c6eLuehMJopNEhVMqYLZgt6sSWOQmDvBST/uuvS+k0QaNwDyf
45N1ThO/xRRuIjnyv1QP66NEspG+/BqIUXBZw6dVzrbCDrQJb3loku71i4PWHa/oPK3LrLxP4C84
VyJP97jpPfYi4TEoJEhUAT3d2KE7lDVMJqouM+LswzAvff5SP4aBba7cZLrMrdNMhSF8ZjH+r+q+
oeuAVDpBXJOrFhKg2QrzS/BkedCFjj5jFyqYuRu6mOZWdpYH+CFFITL6fmApe6sb824yLtFPLOl8
U9To0V6AjeCWEaMKcnbBzAAoIzyg6HGGyoQAErMAnHbLPhNyQKduE3AEiwTWwGfGOtMBK1D/op0q
KxtAgGm+0z23z/BaUXp9kmkBo6IrsHbrRnwT/oiiQsT8rR4XC6EOq8ZekVE7Zal2pEa7dl1+6Q5J
n29sE4WaztznTAgfJaRXCWX1jdrNWmmGXK/ODOiisgBMrXHbvsOLFYVb89BpK+xtw5wz6FdckG05
O9PNWcLq2h5/MaA/PZ1ZOka/nKGoi9rBUWbOv4Pbs7pZ6YX9806Qqe6qJE16opV70uUgJTix6827
ijRC4u0lDPBvvLaQ0TX/+0ltjTAtgMU72pIuCK8NQiwz3G9PcpPvFZbxeO7xvHo3cV4O2tLBmabb
m0bUOu8khoeXOyaFQ58ogTqIStvYsFD2hjV7RoD0ftTmTD4VdClG4ZdH9YNGn041SidqghOch8EE
cVtpfJ1YlQgyKgCu+u2SQhYfG0H8yvnYtxZNarpb43a7T9jGSXpT/KyIbro5JmvOWZgHhboGqQH4
2UQavFGt2wkZxATZls4FNShVzhm9rI/StouxGpzz4iyOe1SzYOvt6tNPqhwp0g2jTnFXQw9XFskn
IFd+ySm0+5Djoc3/6TukcYsNmNM+lt16mcZyzpxwklvav5euhaW99GESkXR9UyYHZry3DQd0kwT6
vIdgjwTHPFc5qEu2A6ai1RvirKSKs0yHWje2G/1iRFMzLisNwEtziwsDN9tyCwKMA6Gumg082AtJ
hvHDlnFMQ9TuW5RxjKk4TqTb1Zb8B8rxkyLHxCE+Y0dCCh2TE1tXrSuGFWtRNncdY5eJzoJGJC1w
VPu5RWptu1ym49QjtO3RUUfrIFJHDqLYPuZtwcVqzWM1moXrLNqq9Nij8BpX7XQO8Sq9bXx+70Cd
Z8gaT/OD6Mas1r3yb4Qw/pL1wJ0PN34LnhIu+0ntniB84x/FRxKKP5noRA8iN4AbSHhYRd4kT9eg
ZH8FmNx51IPYIVghrV1pMAchrkUQvEu+2p82W8u9a6oaQmzDrtWAuSa/EkisiU4x+WzPfZac+CyR
LiknWoAm8ddxqCQhHExaLS+fMNPRDU4qnwEgLHfgzGVeB4ic9fia2QPDRMzHsONRUUSS75QaMK2M
uN4ROtiKfGF+CSfu3+qwjOAVXvR4VV1KsQ6Jipb3jaoKDf3n+KuiuFzSXzWVWz5FN+yHxr3YwfrD
2MIaKSef6mNPiRjWQqa+LRUHFjNPiOw/q93r95asZ7yfb7xAtoRIL3z3fFpGgdw+sm2qhyoQoZBq
6Z911YBk7S56aZtsx0YTMvE/E/+iCeH+Qn7XtTtCKkSqNIvCifF4SHnP3q/0DY/C+DWvzFkvFruu
evfLVEmOmN6QCjGoGZDb0fovNJn8r6YPEU4aFPYBlZRlXC83cmO7ga1MfyALu1nnD3AnXo5uuTLx
oQXrUTUsbBuE9ZhRWCVMm65nSBMyTx3NA7O6xYKxr8TVqli5qOVbyEmWmfBNn76tKHBpdF3WcLev
/+p4ZLmJIumBPlNdChH7oYw2DXfysRDc0op6qXXy3F7xT5+8TtOoePZMGRKgRqgYE9Dob/YQnOId
RQcTynuri70II9NaRbr9sn/Q+Yej/ppc4TGeA+9sshohTOMs4MYUf1x1BEyvG3El82TZHn1lyEov
ALiwdV5N33dMDQVnlVWB/Q+WqFHdWa8mF6hgKHNyYywCIlY7LEMvn79LDxbA45wp7BgMvrSkm36B
SaBzqudTa7dtXFUb3QktABZmdIH38DjxlUjCrtDryQrox0ocIRnUR9K9hiUEQRYwqcFAw64vcbfJ
XdnHiF2JcKaA0uTyjsBPiM8o4lHSDw8VfcruAybHi8L5h3nRIT4WJ9TMvb4NVXvv71DrLuiOO09t
eHHEVbHg1R+oa89WAzFKND3LNuUy5wbRAfoZjDghx7Ctbla3WpZgZ7XC7GDE+GZl64PO9QEPl0m0
g1DDLvSAnfN3wLS09H2PLoL76jIJ5/u47ogFGn/qfHToBe6BpxTh5+J2x2CwVz9ZvJay6RHTcgy0
e+wY3FeRADaohpDN+qAtvxU/TC/hUodEnnq2AG4GqA74YLX6BDqUxlccySfz6EVdIFIrlDwOddcz
a/Umqne5G0dpuy16BXYC0uVEcgcylZcb6TvUSQQJro6+p1nOBl679vNMCYoWSofvmE+x0FxTUGog
ZUv5mTZkst6rBupxwCzlsorhAT9Noq2boaZ/X4FkfhNkKY+wjUEFu310qSDO+N7vu0yEh6Ol5QzF
8jLzYEfkUoznckv3b48A2cz7Ju8MsZkB+OFooEZzV8Agp+XyKCWK6xl4VOkLfNv/Ka1UjA+OgH0Z
OxPm8vl5uW46c5Sz8xhrjLo57C232UNkCLXyrupH3u6sB3jlgocADkJSL/S9AtdpfygFnlIZbSvL
6dJPeuMaeerGMdTZP/J/0mqSfUbdcYlMyjDZxfTXNznoH9jIWiNNts0ZpLtVNynqofd9bKxbVu3e
TPMAN5Ex9+FGVZIY80WA9FWxOhwEP3Uk712zVCz28uBEgZG/lez/eth+k1/DgqixklFiSKJ5G65+
IqwV8Rjel4c6xyGdDUUZMfDaSKLV2zrDFzyVxPF2cawVk3VEHSORR3NnFWDmDnY1hj3LEwToyqwl
gJ6YN4I9NKvBLB6uoLBHUNeAblWo3iyHH6g2fui2VEwHhKx6kFVZ8C2fgLs3zrmBlo52rofEKbQe
AW+KIFFWD0ha5unZtIKlx+hI51c5H5zYuid+g1aGKutkKduU83CKDkLosKsastVquWSuvGkmRBWV
UJVCu1aGTVofJ/bAkahejQiYHhRsfCyrN17PRZUSpEUuGQ3jUX5VYwgkZmABQfEBLZtWlU3u11ng
YDQh1IWved5Dt+AWqgdMQ1J0w7L/icnyZzQHFljTCOKp1i6XfRysk3WyvApFu0VoWB/nTCcwQ7LG
q5Z3NZC9FPYigbmVy9dcyEuGUye4GR2aPa+lQbBTw/LvidOIgY/spY7ZXArI1On3C6Pb/4LG7X6p
z3IDmNjfgWtLwPJQ7MYkMJs0mdQd4wVJBKNCzdqopv5GVrxGtUcnNUiHrQQ+0W/Bhm3L7RoCDMpV
fNe6wZhDQgnr8ZkQvaBz81XgcHQvIWL232PYXlez9A7LWRPfqmVxbIY4tGuyk18RQLJhFIb55Wix
ZDWD0uSQYa5zPvs6jkliueLxB2Co13v881fYbLyfMF8tq+5zbsaxeQO52cuUA4333bEDs++JE4jQ
s1zCjd4eHji9lb+WdGdA4urRUsnBUAX5L5/OvmyEtfzLA4HJzxL8hsgrPFKgFg9T4oiQ2mwiRkpM
wK6YThvASGijVzOlWCESHknBTI/VMjls0CiMaD1dfv0Wzz/mYxHIoON61DP0dQwTq9635Lu2Ed4i
b5rBa/VxWSanntFgcmi+KeAzY5QDpYAcKDcySHH9qc963aezWUtEkUq20TW4x++s+lPvhJefykWU
bjcGaHqjrVEvQHu/n1azI2AX+MdzceSZINVUyhuTqvp64sLbvW2YoF9F0QuPQR5tCM/okrjSo1BV
TTiRqo/Zzw5RZK2SB1Y8U4BCPf9kJCCO8AJa2oRFgnYUTFcg01zPsTfKWizPMrAHBLOnTqH1HHxJ
uXmf79IKGFErFHV99C8qxwc00LSFBsJ5c9b0sMj/uPU3rsVPAkXdFrTNCYCtOLumBNIWxRy6u4VI
1CmX6IxSgUnujef1B5D/BUwQI719oSbzUlF3lNdrK4SXTxRzFN2sWu6X9OMvyUzvWJmNf1IlRqfR
zohd+nFMC5mgMMu0nY/B8k+Ywk3CCDHZ0K0z/mXzUClIOvOH+Q11aMNifiYttAhQqbykUi67fLNx
a2pBHVaihMEdCLXSWWYKXv0sp/7vhjr+vz6G78uta6N9lSAXO/jSmG4sZacf5L2Wz3xZatRR0BGp
aicubVzd/ycm+VwAx48D7nXrOXBXAWC6dF+wQ3l9XocZ0a5JuuGUsH+D5BMgbZW881YTIoXBxfHY
bzYnt9SRkMB2s86pMQ2elpsrOPch4EFvc8FNh1B8wXBLqqVbHm0oNcdgHbRYiWt6LBJ+y/ku6Pa7
Du7+uAQcHtdjdmyxyiGPoCGVw7FFQKb3o6uiJUv+Wew6B+O98qfdxw46cCQawlaiYZiFVAnhff9h
LtzciOUwHy47yZPmSuKYun0Q7PLsLYBwEC+/4V5vmjMYE/Fs2xC6+gQsaJcuNXiMZlZgZ1mF5C+D
89bCrubLU2kZ1P6WxbfcwLshgMEds4a2YT8OM6mGFK5Q8F7EAZHkgz1rnrdCFMnZD8Wd9xSODJ2i
i9Cqy1nU8OXoxp8mcOGvC/AbhuLrWakmET75Y5V3Rr35TMGuBXDepVSnXmFFjZy3qyCF1QJimruj
pTJ1k02w9MV16PPbovlR0rk5eVq0pMBPSYA2EnA+BArwWRP9J7DyLzhInK62lKD7spunApdYoCT1
/IO8upwydXum9zTSg1k0GOUYMdMHYhFKDPM3oVyuiu4o98CHWvbzi6PLGD4BsOMHNo0QPrjREJlT
76BMsiRLuyV3J/snxH/5vkgAw8GlDp39BY5GatYI+T5eCeTPXq0hu4lKQEBL5z41Tl0glfgBOvlV
rvZ1GhVDuVIZwhXNWmbnbYUtDoMdCx7IHLxxY7Te+pXIcE5j0wUrLgep0XzGreDhijapdura51gZ
jgNro+JiHPoSOaSkR0MLBtg7GcM/HKY4uu4korWtxHfOGOjzi2ZDc55C61uzsSH2T7I2nm6gZ9Px
n/cHQ+SdmhKrKAdqbEMIdoA/wbiRjae9OiHFzbb6jV2rsGIRPjh4fIPk6mjSsOkBcMUAF9iYoeaD
/1LK/jaerHKWlP3an4qyFbPsWXQPn1yivFs7pZUj2PpUn314U+RgQEKTRvjvxV6lxN/nUjDevtH4
18qsMjATJalZ/m1x7O6T5DsZCmndWcOebPRD1KwEBy+vAE+ic1/UhRItfNuWc8q96LNrC2pCQQMq
ybMPzWtPuGTbXtDZ7Lr/siaj+ye13UAE58y8znb3OIWMio4kdRfnuJAx6eML+d9cXBmW4t0oFlbu
2gv8qk83yKmC29L9hboNRCzjCL4eOY1bilG3rOtevUV8UVxUdfMEg9qm6TFwJndZcQ059TQf/e1n
MjCE7FhHqqkgpd0aZzVGNSDCtK6sXvxvg8Q/h5qvfv1AVAv6hrGrPdEPhQrWNkSkxkocJfEJbVS+
gyoy4eQprC5KIkmeKZ3llPP2lBgG34HMwa7j4BKoze5dq7QP7c+Ab5vlRRcVeoinuWc3y4e5GMoh
www7ub6/lRurEdnTOPZA+Q2+qhv3BkW34Sx6VH8k97jZsavjyq68d/JY+jhIhVp6ArVuhNPWVaG2
LOgCJmTsAaICRisQ84FlS5eqAS5E4N2rhNuoVaeJqU1XGNYTnSsFe60+0Q8462HdcflP9zs3uOSm
Hh2J/3PsepYR3LyoTPCntsulIm75MhyAsDq+V67h1cuWnabrDigJH98rQfQQp5NOE8HEUzZvnxNh
7Rv7+vXuB/J02m/ceWjAKvG7sVwhtAd40G3Q+WIcF3QldgfI88mDRG5gEc3W+Qg4rPKxUdz6RtF7
L0uys/Mryn2z0adutR9WIZT70YlhYrbwym05CdBawQMcsZYuGOUWrCVi8d/eiuswdZI4pB5NhMhE
wswgV6by7MJE0eKy+B/SUupQGIsdaRa0NyhQcYiBT/+rHp8MtAUimgfpO/2hrhk/3png6mTIE3jv
RpL+1HV4+FMtlEaH879UOGfDMux0fswu6JqYHJyilPeVgfVXXUsd1Ul6ZjxmNz3VM6xljsvnML+j
77DPx/WyFoJkHfw6lVYinKJmTfgrQFq8w1EjjOgOgXLfq/hat4YSy0zGsTPB54IvV9c6Mr3p0rfk
GDQ0STLCMFYRIfJZQGhIuAC0gAmjV9XG9s3QRbxbd9pJqPge3P2Ja6clt/cn2bU8WKclHU0+Zi25
Xcb3EX1drpEAlWN5zcri17AeWupTm/aWy0flTDtTFJdBcuf1uUkc2O5b/t9jUSLCgm3T846Gwf34
+d5cUPhudZswvM1BPkxL/MbLrhkNlG+lfR4E1MDE3d74I1HwY3pYgNxU0C+RcpwCniesv9xe2tbd
I7RRTKA1MmGCNHYaA+F5AyOo8Pf6J7v0Nj/HU8aeJw1Q34eb/h6ksrbbERY6XxtIVqX6W51uFLtY
7QlASZR87h3vdlMCueIna1it1R3BhOO0Lq0zyfph1DngGvb1oPzZa6x7R7945z7cdF+e1zAk2wfx
2uVRw5SSXeAoXLiX36QfOsFeUIsMKIne9nCOPezrGBA30jugF+VEGabxMwboAp5Tp0qiAIjgmgo0
7Xg9zZtkJNHd0rKUJ0beH1Z1/NOu2bGPnwfBuFyq80V4S9+g5n9G5KKiPP0RvcHGitgbG1ne/hJR
ogdYBka3e7v1E1aFhZGzvRHW3ZbCXirYvCF96p1CXf0yb4hLzxTjWBzCi3p4iID8j8UWlbaC5Pme
oo78OEncbw1qrlc/l1tBpNa7VZtWf6hXxK4MvhLXIJUTpzBALHOg4b1jxLbOcbrodxoe3foYQhgk
ZqH5COt6AtNPG5G2C7RQjvMcpc4OdVexy6lZaUxWPQqQs0r/21LIwTnfB3bm6k6d9ncxWGL6WQTe
OsZaltK14vwByK1kDODlim5EO+zFDA2LIVZTwbflrZ3GB8cGNYEjyLTwo01l8rNk0D6tCJ/yUZi0
WtVrhBqWDQPc3IWUEvdr4PvoI3ZBYmxC2j5rvhYh3tnd+uf5JBqaEKzXtTBymSlsHerfH5uzXWsX
MPW4Q1YvcPOJEVofNiFKXXVOzGWyquB7qluQmD9eqmTkV1p6OhFPtZJe5jMgTZpSo0IUPDLdLDqf
J5QeCQFyFhbummCYzuXGt1IMU6ReORkj+t84JBzUkqr3cv0Yq0GhPLpfdrdl1uPzqSBJkG/eDMKg
ceroQ6v1aAQzvDO24cpptGoVFoDFaYnJL+RQMD218qqis+IKHQsBB4S/FVIraultovRUC2jVwKFd
UHmgEc+pLxTKe3UEr6CrnDMXVNfnHwiVureg1+zlAZFc1x7lwm1xW94V6708S8fKwyGhhJUNCXni
/DHRjhVAx1Ig949hq83WF5Jv+1qUd7ljURHDCnPV6PptmdIYaUy661QJvHUWIM6HmoqUf6We8RD3
7de7xSM22/5bvRknmRVd/ryMMdlXydpAX01V5/2iOmZTjrOItZhIaFZRNB+kQnzTX3N7G6ITSXZH
1DfQzIPwFBun/xoG/5mPqMqtbQ7ssklK79iX0m1j5MIXzsI5SZ2ezI1lMpN0JVlsRYSWSCAu/VFT
3OgoBHMC7v6RC0XnAnsxj1xXrNBx4uPVh35jGDN1I45OgvdETR7Hl53yGXou7oLUyd+A7PnYkstJ
aoGyubklha/GCsByogFVuEmuRK7BmW5v8SsGHyoPoUSuh9m4y7fkNV1eMKnXWYFHW5o8wjr2lv3M
vNcDpZT3GIDnC+dGhyjpeiWkU9i2MiwhzFNwl868R7+fIRVBXn02sjdLt+qr/SZM5DFOg8rpqoK6
pF8ggYqo9M68V/WfkQ+liHLQlS6LygegtrzdcDuFWIeZDF7Ptcazc3VT1pFNTfpCdQbv1DeSfODR
C+97f61SNGXRBUMtkwtGRLzw3JbpjU9AAHkViZLqZWZ3ePbTf8fckiSetuA89RipatrYYrosjTRC
gGZvHo2GAZtDE/xqOQjhEchx00oNFUCZwEKnqDf38Gp/HhrUZV5otqUcQnGW50dOxvXcRDBpprpM
IzHtERAId8akiusNgvRnSVs2pmHsR8erkQ/ea7sp1wdMGIr+1k4dztevJ6liT6Ic36wcv8fMxSDg
gpJ4sXtF+akZnbxJ1JynLdh7LHB2ZlXeo5ew58VUKLYIMC/tP0o+DxKjIh3b8Hg8RqxsBWea8DNh
3LmGenMbXO0GED89dHE02VOz2ALuJ2uwltnpZ+JtCvTrsYvymls8Dd8LjMTfs37l+8VN9v+uWNFy
dfDXWrEFwAv0D0R+9zXxFyrIn/biee8ETMT+IMHvvAdYbubDbQ2tW/37ITH96VIqQv+eXwGRFHGN
9FYa3y9OOm/EnVZCoGov7QghEb06EJS9wRv7jLlXJr+1OybDEzFC9NGKnD6HXguXB8Ej4Qt13yp5
S7DR+dBsvcnnxxht9Fku0FETvxTrVAZzv+nhpR1QVQK4Jy3VfskT9HDtJfvINt++v8PyN1AheERZ
U1XD83rAxMk3gaT0bUtHT6gIRhT9BfJ7MdIOXILGqAmrVXS4Pc/fM/Zlkt7mL75sqOqyCqyKzp12
1qfxBkt4F6B+FGw8+oGxLBMu9BqZ/PbeXehAzdhmVQ1zjngjb1nwu9WcbEMI5lWQbhFEuYLhimIT
9aTKnpa4ZN54Eg6glVp3oO/HhmYrS7ROtYt9g0lqEpwM3F4XnoPESL3zjFqpcUETMRmdsSqqMzPs
wSfYnb5igxs8KlWQY4NnEaYjI/r7WFGJ1PFOF+9GjyB9Gq5KhHPE8W/UrNyrvi8rls0Dl3SXDwtc
Eit48WHyLbsZ8VHSUblKbfSM0HMsHopLqZ3QjDvtZVqFmCjeLLk/g87KFMZAKOgZOVwsfnDsjdB7
GkxV15zd6mb8eqbqVpxFOq5UaPxGpun/NH8PRRDEseb7htepLS1GyOVRtNVC6/NwAVjR7ZjOH+Ks
5W5w1BXfmM402U0xnP0r1/reXbQk/W1B9rh+7N+wmH9FVVxPA8LLCvesNBZpuaUYLxoSnQXJsMCk
kh4ILjkFn1EBtELJhmcryg5HVeKnxNIPWlqq0191XRaKHzXU0Yr16uOLjVLK1ZM2jMapUeyjWO1s
d2B7Aps656nzKdHIt/YQSc7ezT1HWqS69BT9DNDVTTPQJtmgN4bhN0lDpru6or37k4XGQaAVZ35h
lbWaT5kwjby3ylFzKGt/4NBdx8rA1DJqSFi1a/geR1rCvVYTLNrItxFH2CaTZRdQ5yUOPS0PVDoh
twglYWza9KkY1fEiMXLAekGVRHXhAqjF0uL3YEcKD7b5YJa+T1aRY9LjPTevTHybaJ/Owlyw4lQf
JLGKch3comnY/U6AHpPPEV3vRzF1p5CkJsup0Q0ZkyyNn/LCtKv+HlbRWaSsp99BaWOISWg3YcUM
H4DhhjGnm1i6H5EgH981dqVe+J0mBUlVodIqKVqE7BPLGym+rYRKJ4bzkMb2+Qvq9gAnXaLMNi5h
Ce2vw0kpx4O96bnD3SAxHwkacL0K5EHpfKEhjQRY2mHSLp4SYvtLKLeUcKVlzSbRkB0rgfrK8AFd
X6u88YcSzsRt3IB0d0O6Cqsuq0VLrdbKpHNeqIMF0WggIVAJbR7I+2E68/ILL6Qfebse4cJ2cZ9u
OAEE+CHZlx97eaH0Rn/Lb4V6ynNQmylt8r0HCpd1HoPmYkFjjQ2Evs8P2eGuyL9mkWNN8GWZSpa7
gsx0gaN132O1S/zxEAp2xfatGrq1o7V+K+CMdcigaWxGsWVAzz1ozwNrVUWTprmbHt/P4rwPe9pI
eKC837Ksjd7MCT/V5dixTVfrYbSgWTlSA9CyTuQZKXKEwvxFEI75jaMogrv7lAoMticUlO18swuV
Cjbcx19PYJ7n2QFkuwAkGOoFKj64YdFterS3s575XpngV8GkF5FNaUIXI1KqmPMxfvEkbgxMjMIW
qL8Zp0eXr/c1GK76Hu+zTuoOEw8MfKYGCAlKDlF7oqGkXkvM2Ma9ob61YUo0tlHGeZ7y2baPCAEi
x//gSWAztPTWuP8TQAnsKbieiQ3jp5pr10bOW2gGfAz1TmF9F5KHnQxFCL4fNphE5BcIeDRXTqMT
ysL5Wz9aMBAY4ou5+58FOUFWoDf+tIe7fpkvtiAm3O6un1StibeIXHIERk5j0wE9Xd57oEzLNeuk
uNQPy49xGA3tr56cQ5k/kBonBwvOJxHNxKkE3+hhBYphgdvFd0Dqgr0yl3+kL59r5LvZloCkTeO9
l5Yz0eVtcCdxmCZ2TIif5sS0EaPofku+MbgitJMpaMsdek7ni+rjDExUcKzL8Xjibfl/oNWxMpfe
NJqww7Mix7zSF8Vugk4I8v667IwhD8XzPOmHlH2nnXyhzjnIsbqctULyNFj4g8II4XN+Z/auibVI
rea1UIX2mCdQKBvaOI6KFlofSgbWe9PzqiWW2nsumipghElpCQs/sTH8t9d3NVOvqxdoBHa71j2I
A9foGTTt4/ePsCDVrIAXs8VeUVH6Ba/YFaCAUx0s2iDtRoJG6eKkDLYApO/ImAFzxCDx/hURXsxy
rE4+51ziYJf3IeDOfP4a2kD/zcEt8Wb4JMLUFZuLQdQ73pZFIWCz5I5gNwMpEp3PUtcDkx68M6Xp
1CHG841iG7Tfo5IVDrFf94uYkpg0ZcpEDdAhi4wqy43+8gdKZKXc4h5dvGN0EnyhPKCSJL7eUa/x
gYYFkPEtwKEsXPDpF3azL/m07EAoHSW6j2WyoDBceUp5asGOUYTzwNiMYwk1O7HiXILl7KvHc1Jv
0FHRSJP6iTwh5wuOBl4JL8ZHa05JoChZ9Nfz7T4hdnPPOS8BpxgX2aW4ZqD7CMxSuMurJO3LMtXL
FWLn+1bWQjeux9UH/eiQDr8ftA1vnlh453kyS+JqGcC+4ymcmDZBuaXokTHo8DhVm6OrxwrdoJoI
7ZsawwXT2xnRmhDuoWMz/CY12Jd/V4hyfNh2iXXGfksw6NExiqKaPDqfoRkSIJAnXGq2ZnYU+jd9
NVKPHjU8k/8JW9F5/bIsz+OD/9PGOjvTtrU425UdRpkdvDGQegRsnKtG1JpNik/fmIPTrb5yLC+w
Y+7j1W79Ik3iGDaT819z9Q1GhriSmpjpMGepUz7Mg6XJ+YCh9atpZ939i9UXbzJmYXMGe78n+Nfb
DQCisHBJVWzoAtQyQ4kfjTEsrA5+rvIYU+hNw3EWS1VXSp7+f/7wNpGxIRgEHEPweeSjZcr/0WM7
DMXlA736RYjMxKaoNbKL9ud3rtE7YmJMoxjQ2xDGtaf3cefrNmKPtqjzU53OH1gYopD8GjGwQt11
H/jI30RR7l2CQw0KH+BdSrEArjSMsYW6/wZfHQrodA2b9AO3RV3At6jTMS+kWBOeM30WT+ME5xSC
O3iF28hbrrCJNnwy2CadcAk6zRZklAEv01J9JLSUsGYwlYYshMsMHzS1eyoy/1kIGsRuNtDWpQSD
uxf9B7+6g1/JdN6ct9VnN/JykEWdnxsU9mNB4XqWdYxficQtPeEYwSHMoGh6mNO8nYw1iiOdnfj1
DsA9xXwGUB1qnDY/1qdYQ3ct4s8c1xfJb3y3iL289ODKKOxdO0cUiE65pOovR+yN24zKI1kIWpg4
+t8cTpG3IwrSmKcWQ4lkAY1ffEXK2p1Uj9X8kO2mTS4y0Bg0IghiuOQvSvU0t9o1Ip0/paCvhq3i
FEEXcSo0Lr4vrtz1f8PRrhrm4k6EVQhI5YRCOYP2OFPcQ59filt+ZkSjidvABfvrjSxVOrULslA+
X6qTZ9y57tCfu5kEnvm2Dlb/Ex0yerLF3CVXCNYgd3pmfSTT58KxDp57Us8LWHB7p1FWMYzCB/88
BQbVxffIxZyusfseebeMIv4z2kvDhsoScxFS56ZI9WusF4FsJZ8IYWhHYhUE2B5Kg2ui3MQ7vj5N
yxgVEzraIiksApt/6ViFZZGcVdo9XLajWFsDLV4jHR8pgGfzJm2Ig72UCwhUtNZrlj0FKrbuAcul
mDRtJ1+MB0NSbSBmQt0DuS4SlQe/AldZjcSHqS5yBae2swdn/QdO4sJHx7FkOjC91FuQNkFuouxK
WZX4Te6sKL1uaaqUE1UMzG1fhuKylMIbI4A0M3h7YTa9j/ZO7HX69qV5s2DlJ3iz31AtrZnpEuJO
PCE0gdHkJAUSvLNqqF9PutDGVmexIEm+7E8xZSL1eZujDlE4wVbs0FLm4bPdCPa+aY0k19XtK4yU
+g9IclrsLkpyOEAfOmQsTXmaNnm9yJXBgfa9kjRo8SeprYwZth2c7D66vyHUCkvAsbjmoXS6OEDz
gO1wpwJHKbg4dP1pnKmDxdBjTdinYgA2swL3L/ANRq2eMIEiZhLNAfWqmq+k7GhRr9SWR8Onk179
4sIXOqjqpAQyQrjqmL3KiHwfgUpTV3KCAy2kXj79sGZOfry2Ca2S4KppekV+tpr1NnUfS7dljASW
/aaYyC6HhzCBgAp60umHDs0piGhYL3ZnOe2ugFmY8qPy9kabxsq6vZGaTHSllh77KnPU6uowcK6i
nvoZLcyVROgj3bqKGexUIX0ym91waFSlPuZ+HjtesOSKAZgcVH+FO7hPeqftmRYF0hHR9pmJeznP
4FCJxVxBTx6ZbyS/bZpVBwppKx8rHgMP6lMbxZI2pewnuQbv22lCP1YY6a108NOzx7Iybpb60ZKZ
VUVsoV9aGoMahaeZg0bVas/CVoc3OAvk4qyuDnBlJ0SP5F2tcMXApHzsI/s6Xg7P7JC/rDK4jp7W
vgGWdHoWQ/5Iz7nxTfWVtcOPPBlQqNJRvCiBP/YL7qZAA4AT4yrBo7+daVl3GqI+YjAVwleQPmFK
qN7HChUv+/cPRGgsjcA78yrre4g7+iwbMgLyM95PYCuWkf9B52BoNS3DL9oN3k5RKqSaZgv0bUbO
6s77MLrN1iAh7xi0gjvItgWWqmem9M0fBHe393GigJGhEKI3qDwkM7aaoMWLloYiqOvHfozXzdgR
sIfgMqgGw+2R9wj1vYUKxcjrSUyOy3yGPYSf8npcwG4GfYLGcoYdRU/h3Nmrtu5F1MSeOMkWLAhF
Myu0LSoz5rFnr3CDoxqjyQSyceVYE1wsuapM6iqfhZKm47E1/hZrrgpqS/prVAzyGvK9824b/bWM
3FOpm3R2N6WtMUf1a+xzGHe/fu2elSlxLW2AHQgSLZQ9gDseIwijLXSmDlKa6R1Gd9yhq9A1r/H2
C3gW9mBQaeUK+Pud3C66mFaMZF0uSgdmhSYqiO1nQqlJ7FbVyr+ZueP3Ehb5KJiOLj/RkLFsIt9w
dXC2uS0ucSTf9Gl8MKHrXOS372VnHT1bDwNUHOv1ix8VyKsFD2QKn6u0YHwpdnnhVw66MTlZewz9
Lp5+ZjRFFEySgUeLMrQUh6P0xBOmzRisoipSRvOGQYcdhjvakv8mRiSMOc8IH7Ciy/Rww9/uEE6p
RYEEYEmgUe9lTPcK4TXxQbqQfwfixBp/lCWq9m9nUUNZz8bM/ZauzH7OEWrdpbstiSPSnkFlvV0o
U349qAazLThPsHGEqHs1d+S0Ueg5VzI76QOHhBQjlrTuA1lbyy8qgzFfGU+fCA0Ob21msOr63AMz
knhHsOfscxMDTjk7rrqlet9fR2AZJUT9tiKYZRR7Lvu9bjdAzkRELcyv22/60rS2WQiV6Qql8kRw
mfASAGkz37Uf82uvFgBycq6lrW+jWQi6VTwS/r2/QxGXg3UyyG5aXHfrmSkq82I6gJ943mp9PeeD
tNXU8sr9xIrd5Nvqo5MlpBCaiLC5sN9Ufigit6qKe5Scf4CnrH2X7RvdYCdN6gpHJ7sO5YO10S+s
zoVBIx/HA+bBE/hmJSrzm8qvMnqQ4oJ7ad95HYP6uRSdvBabJE64Njchue4fKU1U3Bdgl60Xm6T1
d9AYeSt3XBjGLX1C3W5o8VWdgDx5Po9QUgvtp2+/N9icslV9skgISlYGlAvzG+MGljTBPBZM0BmW
qwUcTlSfmLBd7LVL8CrclbzfIuZVp0oCOs8mt3VJ1YZFHFXSL5LxY+gcyhAw5Ixff/ZniBoiDp/d
ZbLsHYi3Xlx/7oWLG6ysNA+8Rza3kfAX1qt+6fuCg14FTSlvJRmw/zCXEkI/JXGRTYwUJ/63O38D
TOv1Y7S7KEcskuvIdAyulyMt2vyF8n+/9gu+LUtAORQk9VcMIMlE5UBeoUsYqAsMy4U/WpDBnrYH
o/dX51MCQJkHl0G7OT3sKcJffEzrfUbY2srvMTWGt9aKjSGuS6LXtFO0nw1pvJznscmq+IABDDvU
UBB5K3mvKObQ3rVq5mzakhjOz9ZxRqwyge6AcKxqmR+BtpbHFMC22otBxwiBBTDic1RKXS9K2/Ag
TJBQeDKLBqzHRwup6ysfO6OkqnS4QLktpTqAcl1Z7jlfXFrQVCgGUKlrSz4tvDOqcIIFdo0Pnvjg
8yTvgDcgeI8sBWaDdgBhWw1z4re+rf0vMIyZXqcouk4gudyso82k26mVo28tqecT0pEMArN4Fq4y
BnxcjHJm96i0uBK6bYsmeZr50yk9wSRXqmQJoF3mtOyc4OwVDy9XU+GQodM+pSoABo9zLyyrzvXV
d+e/O725+q0KirokjPldmrKH8AABC/mFxp0PflVmR7FtuvWXGf6SoHDB80KNFVzGiHJjluVJvB/9
FckzqyX15ULmVMLldmQ3VGuYwUcez2+DdNMYWM9C0gmMVrKdhhxpXEOAJwvX8Uy8tjCxDrxe4vjK
Mh0JZetxR7CNA8eX1nsuLLJZERFdLZrqToIvGa7XEmlUYJOcfgydv7TdEIkyrdiLTZVWXFBQE/P2
ONsoXV0n/r8LXOaEsBjRgvbkCL6ZfC0l6t0kNC5zdPQkPdkOF84vt4XvNrgyXB+Zgad7UdNekAsi
MOUQqvkflX0E21phWkrAxSQ/NcO376KZ8Zc3r5Wnsky6M52YeBmHKq1q26pKeeJiLN7eyrSR3WP8
DXo3h3A8hnKNQ2k6rV4ywkWlO2Po+cBYKz7eLgODfUgX3iQqhJp9GT8O4c+79tYQm/IgCG7hluCU
KSw00bfgkbVZ+NVANOFYk72NYYSluQI7UdPgxhkUHmBHeT2eMvprAYIlVpT0B0rU9hQO1+Ev81kF
VsmJsCGJpoQwJeVTnsGwxs22B1aTuFnKcA5Dz20bsEZvZUfTwlMO+nE5R+6E+q3/t7eJMtBS0cpw
iImHYUbJ8KU2sWdysnd4+uib+N0ZxEmkOBUN8yZvq98av5U5U9/xXKtthSpJj8blyqaWw/3N6GY1
BvDrouHD53BuFCVw9EeLQ+pGgNV0JYZCBJVEh1OQ47qcytFch88DkPvWXnwB2XIWRXbRiUafd3Zg
eYlux0VCXtOYn5T9/q8S3xMeRA/KNyjtRy0W9xtUQOuFDmz1sBql2yW0cuCCFJ1jthEGS8sA+ijX
dgS1FVvWSu0v341k4Tnk+KMdor0xsRAtdDCNGR0fjGwhMGm8oksHzQK14UfpP9chvwB0iMIn4YVZ
m6cZO/9VdrURaAWUSZi8qA408MVvP8wa1w0FMgNFI2/ILzSCxD7yIw089v+Cl8aAXI6e1+CJz4bF
iUb3+FvvyGYElS0WeKettOpOWNsjW6iLeP8tAzLGXvrJV+Fk4MaSnAT8igIpewp/SeXRa27KDnh1
4aMmAjPYlOtw2ueyO+d1dgl0dea8ggilEKMjpxdIjQ4qZr9VozYKi/uBAuBx6gjF7BBGoO1QHptq
/W1nGTpQxSgyFr2NjA+Uz40WD2U4HBalbyu2YNjSgoX62+PBU8WMlmLkBoLP68LSFbp5yZIs/ETq
GuzI3CXRjQN46ZTHolM5Ep2LvvILy2UgYIBk0GtSTBMHETkLZIs+B0ehDbvPGyX9wMpCVErtmY7Y
PZ+9cnLnoqvVXyA8olrkl6XDOcJS8w0d8eRnJbN/xZESg5R5SHRnP+bh8cdFcyCzQ4aAmkbg2p0o
+hj/uQT7tTdUEI5HObITb3Ym0bc6hOihFVkRStM3g9nrvMkdUhp6eaSSRFFn+x2ltR+vwijTvXss
O/8EzIUeKaM8mhFTxkIEO2EA/S+DOqz+g9GaBLqem9Et/6iYuj3OtIHOHpm22DrmvquW29UXFAVv
f/p7WO+zT1qDuu0uhkaz0+eu0Hx9rH5Jrrp7Fh8gT+Fl/uHR9bEJBynMFr0xrPnK+N9AQcqVHRe+
/WpA4EdT9WiSK05LDk+O7YmRm2eWLhM0E9owo5b46trKYC/zipFzN47U3C5G/dDMokO5fwzqWN3s
hXP8XeXz7h4OvOqE3pLSlvV8sT5dH7MMVPwoyRYZayzcPlSPuaFXwxDahfYiYIMMKumF4hohfSbq
TJk/1GYExCxZAP9KGmG3j9ToI469hJhpWHtNGspgb/Je/5cbx3YnwIBjps38PaoKk7daCv0lCBsk
RMzkPCXABZg874INTrbpbjV16UI4a6ZVAwvEL360+di5gEQngzpfbo8hAcEFGIDBiV+6UBN3P87H
T1A5KD8KYjiYXig2QXrQdzt2WntW0zPlnXhfqXGqlJX7urt6L3/7HetzDyYP5vGgtVj+JsUDPUkL
sCOnDBH5K5oV7k6exESCECWn8bI0ueI660xYl2LXldF/1gswYR7HMF3fC1OtKnxZsiKMiwMOmuNg
kv53M1J/inzJfBJBKMwI8wZUUfi+Es/I7PFpKi0T63P85FVF0iqdBMGiAerGtrnBeLy8jY/VyqnH
oZD3QkLC0nI1QInjP5wUaiAkYaOsSRW0/g1vc/vscq8gVpRM5uRE4dLoothjC73KzX6ZXb2YLEhZ
K7Jgiq3amwsRXwfILA3oRt/xwh1H6yiERVk22HzzXZKwHqGy7A6qgg5efYVoYcNYgAIqaD+kTpLF
AedWAEuC1GHEcwpEoBtUe4klvKcoVOD0yJKBeht43FqGTBlVo6vAHlE9jyA4hJPMKFp7LOl+NYe8
cq0rSB45cxGfLniI39Xz/He9bNmJR2XwrVIkh8g7ZcKWX5rErakO5zCjAWVSb105QwvPIIYDU93I
l6V1OFyMQHJm9IwUwAwStDpU8ohPeIqTbPV3Oyq3eJ52Uzows1UWj9pTpnuSSSlPNid7TqlPP10V
qNwVw3g2RtiLJZFb2YYfCKHdmUJa373/W0ILGO8Aojx7GL696EP+dG0jZWqcvMPMgpC9mF+0KhiH
6p+9oe3ZqYKP+zz8CdlyRBjHi4iZGNWU8z3gRDEn8962oQyNrG5aGvLhcM1Z72NAXzt78MGpsTiY
pl8S4HcOwil1ZYV9GVIqmKlsYMoEDOSt1o9BKXy6D+kcwF+uFxl5E2EJ9zzq0ZbHU6psjubB3nfn
LkhQ26IS8XdB+64pU4hb8z0Et4L3Tl10WPglNHYXweyOjaieaKZAbKj0oBrbo5zMCVRajWx41FYk
Hj7Td3Iv4ef/2K3VX5q75A2fRy/kzBfnDZaZQLO+kORJ9mwZRPTN4SIIymeCLqHdQ/is3bJeiX6w
D9b+0MpLeGXdOeCTxlfIojfLmQyKYw+N/d0jbFTjAQVFeQtpWichjRQvE6FYVUKyOq1xsDlSIs12
n0o/i6lJ5NTIu+7lNYeZ0YB4qXuCLReM36ILSrff3+RMcJsrBgYSW47qJBmZPx6u+Wtt7vGSSqZ0
DTNdKqU+mIV6FhJzxwZRrXQ2aLzzeHVEz4gv++NG+R4Hv3hNxHAUpjeZTj07621swFewBWy2bgB2
ebhK/YCsBvKJEecDiKGmCzk1LYFiIcAIfqTffjkAGZ6jSW3YlXXvTA0jIL50ARFRfyC8quPctF+l
5Hg7DEthAsGn03e/ESNXrV441tl77tPdkI7tHDskugBfN/Y/PIx8gg5IpN1i+mzK+OJ8qd3Hdivk
DzF2+GROysbGHlxqNdz+N0hGOjxjC8M61HO7u1EezSb1TYkxcB2v8ySSfR7BCWoI/Oo0HKzUkD35
4xbq7jh0f51bh8W0ApS+P1qx3ooCGUuJOR1Y0luFnXb0LeHGYC9pJCFvrzHa5cAfnC7Z5IJBerGO
w+O7jz11bx8tcQxSWeXJospGdSTcf7gVFAj3pr70WZuU7rjWDoo0jYpxFoyeFqZC4t93JkEqRvIX
Fbm4/8mb8ipXZjYAK8UBRbD3h/29bv8g9q76+zdDJUV+bmuPRP3CvG5GYjwr/VKIFWHGbzu5cCGT
p9Ec4VQvJkmzzsvolTJ3SC1xyN9//mwfOiJjZ2ZbVYoiXJkQr+ZepG0SmlsDbEXG+KxaBTADytDU
+JdMEKIIJCoQzW/JHETORo4OPOyewY9VKZisY+Fo3Pf4ydEagimAjpPrha7GHpGleaai9QggxM1/
QwQ/tEbz+GsUcwM2ckYQvpLoL2UvOG3mfDbeqE5IHQGmPIycoAoeQ1WueraQSCzdnJooAM30BmCV
F8Ljg44DwsttSkaZjLFrN9dUCfhJdLOiPpNVO4Fi1xPF6p3IWqMFFZBJ8S6TFs2iaAhD8Jq5QfAj
l9sEra1zV//fj9amZ15+yL6XqwNSvoXiKQ/5nZTVf74TPWUi45oMcP7eCf0HTuDEODUst8BZdAip
BpG+5NNW8BL/grP6bWhoXVma0EDrSqWrH7LmuPX7FkJdhbcEr49bbzGGoM9AOlcqbMUG5LULZ5SB
eyoFpY82P5Dl2e7xFSOhMIYYO+ougch2FAij2sISmoUDRAKIEN9jEgOh2211rwB0bVGCi+x58rEp
tqV/idwdMOK6v09CW8Q9X9eJ1WVFUVAj9qLrYRCBjsCwez+6DZBloroPcSBnrvPH8ZLoFYTUetZT
eg4QC5OHsKT5S85eJuHJRDLTo71IRTe0YdaXwAa6LvKY3hevNrBhC5U52zH182JzlYa6g3XFJqez
iGiXKiDedIqTzimRGqbR6keUoJGYL0LlID1QyYC30yfIzeBOqHGGRq5LqLXVvqedQKqmoiuq65y4
1aL9p6Az92x5eZdnWlQPdw0+eblpbYYKrgJQe0e42vaZ5u8wDnXkSn/UxwzNR0xCICQXnAKn4iB8
UqD8P4LV6iomdVPODOGmZlfIDNMgxRWw29fL63ES1NTbve6kd6J7u7xJj4QmP36B92vp/0h+FWeU
oXrXYuq1KqTDP1gRz6DcaC/NOKJeV0APG5lPERDDUCkCmpTuGhWug3gHC0Gl1f81d4oMhPp3ZlfG
cf34g/5/mW01MG/mYFnAZzN6QWL7RTiOiam2hwR2a4Zu3WFWnjxm+4zTZ2gG3I01796hg6j1n4ze
lzOCaeSNsIrm5QfiMDBYROVjmGR08goGjoJefCE18eDg9EvFtE0tTdpWFMWd1YoN+7o3yudcoBT9
JmIOr096J0symESXWNx6URPOzSr5Ss6qvqTp/Xwykjop1baV7nthNHGyE47kxkdiriNEOOzCvQz1
UWTt+GdKwyH6oyRCYe+H4OibVs36amDFQNr4u1fyeTpjS0NG0OhXCB78kNJLzPEt2yhtg08kB/Et
4qbb6lf2t+CPpiLcyyc4tT7z938tjObYaeDO+FNYF2cSF/MDuK7vrCekq1X7JUBYBYkt7Ogd1ZuP
K4pqtx//xwxYsHUdngdujv3wjqJ4wV6IbMucfvoQU6rUHqz+1hFWKHTTwhJwmoYvhBepwepXweZP
IYnho+yVwJOg20lp/k43T+WM8ROAPkqF6uUMuUoaTKf/XsSubjhbFO1DTRaLqks9m5hUkcPmwDET
SIhXC9mzgoenLhfZrY6GpaBZxVZ0tkVEwNdBHDT7AnWeNfkPF1QWi06sgVA024ZUxtkvznPQilU2
I+MCglfZm1JNo3hD0RwJG/bTywtriL8P0ZFiQ/Qhez4Yqmq+7bDZ/9j752Tn/m1rUfkho22+pIaJ
nwpMo8hSlVOBoK7a+dgPrAvwtiaPXRAcGVJgrkZ2aq5lNgAHNQXki+v0j3M539PpijfLO1j7mWQI
NGMib1ayPlRRX+pYIuJiQrQldPGudtcx8+kygMz2ic+CD4nffm3rHNbArWxV61SuJEZKre6yhJ65
xWklgab5F8lEgCtLrFoOgt9SARrSrVpe/HHf7AdE7U5c0/ix4gOWHgeyaYa+eVWiafL6li1FLV3x
GhPBOFyHb0uKi/lca1xeUK+vf/cfY0W8Kmy2Mz9rKtvf8nUCSMJPn/4rpS7GW9D/aM7KhlxqObP/
fh0YrQ6RnWGeNRIFSJU6iy2kDSU2+iR/YES+rBKN0j7Rp4m29CjDe8fgBg62FjeqROVyzPaYV2OJ
v+x3SJDgZ9Pwb07pDFg1A0PT3HlYSpeDdz6MtM8t5W4bWz23leMlTSBJE1vxgwWjIgPfcGdZVqNF
oLEx1sy0+9b5idS7SGHyLRxWrotnzsflRiVExhJWe5U7TFJ0mvSGlIZ1UeC8Gfat0mJIXOPR7qgk
mmC1tZ8gETKvmXiKi3mk4iizSswNGbgmHWwgN8YXSML/aHslvvE+7tv81ynM80bGWOiIJgo5CdCZ
wxJwtlnjXlWLP8L7zaxquO0wK7f/UYq9gaLthr+yHZmbiLmqEjonlMPZD7VPAFhMQCWNyB9IDWgM
neFotRGrlzFquve7rs6JklnsEo6oWtzP0iALbuLV8la3TbISrUq74syb10Fzp8RdbqufUCy/6KBb
vozzb6DSeCyTKr2jn3bYPRT8DXZ+FbjdlKeZI89yZAWre4r0vbk3drxf9rQZJMYT+Y4VeDOdjBhC
lB3jdKvCoCqrvjYu+pBcglrru9UyiBh1AcYyc77Z/P3Cu7vDYE1iWumefz+ZiypbFQmwmvn/bZa6
5GDhcgL/ktwWqq6+WX4zOdJQAlSEdkalGrxj0LSQIp4AWO0Uas/DkL4wVFKFJAsjyy+kHlsIWrrh
XidYmM9t1r/ml1W0CF7ClzpDxNwLgSD86kXwkNveMvSPoMEFNkC6r/KrczslagyJHidWh/twIXtV
RdhwP0f9lj96bLLjFDP4ooXtaflwrZQKnKIMW3BGUra5WkkbD0LN5X2rOUy5tpYDR/bvIW/07Uzw
iNDiEdYdfMPdK62vcAiq2MlMuhCwDfdrpeVAiZiA8tp/n/TZ/MMaiCsRQQmS/kGy4PCFe+7S7P6c
+kEBdQd7tnP7WtjkBUHiH/SFE/k9OSdDSFyeQjLgVORf+kCLtVI/sMYw1y3zKgWa+ZyU+5WOfGlh
RiVimg3oNn5Yy8Rdt+Mo0gdkSIBomHna+oCkAcs67h3rcjvr/12Js/S8M5whgD0cyT2Ya+V87w/m
5NGROIlm7SGk8CW5D+HTp2nOTXAYjdKnigiFCWT99iE6nDZFLzG3gazVOyDD6YVEigBsgorLJSAY
obB0r9bavzRS6nQvRrIB4nJMaRKfFHC91XeCwA/GX4YqLZBdeEZtIVuC7EB3C3reSHQhLIoEIpz4
u0fXjxOItB2DGbHJr7fM4jxkid9kUWPpSEI8s5uKWuPRxSOd8TVL6E2hvyq4MENQkRjXkx+E+2SA
fcmdpKG8aBzQmwsEMxE9uTEf5lk/G4Be19st5beRur2jNZ7oOo/ZO8DntQTGG/l15osozbMbFvg7
B4nTXvZc/X84bsldoxo9pP5ZifuzM+1TFaUhpwhsiKFtRZP/h9xR+su+CUEbeObfhusrvHtvWDYL
52eb/JaEihIOd38g31U6gvKSi6UdKe/Ho58KApS1vrpfy58AS+YVXW0ZH1lAHwKYY7lSKLM/NsxJ
b6XRdAWBl8dtMETAN43PCtcgD5naDpYsyflbvtmTITPumi3O+wd3ex0eJw4uMgWYjvhvD5HZ2NWB
1qXaQ55rv14usIwaGZCDKgPVFt1PNTMFj/XVyMR9YPFb9w3edkHuxT3iaY956+WVnThQu2T1rXG8
mtdg4CNpyuzOmf592qg+jqSrUuiH6E2bWnghgvh+lpA/0C7Mq7gXCnplGYeXYEuD4eTIQdoyW2mi
i40iS+UpFp+Cj7Dldj590eaexpRsQ4Xyasp9Xqn+336yKQsmFWfOb085WNz9RxHcuM8ZBIsDsbxc
sCS4Qpw5TDO+mPFM/igTwwGgeBNmKHVBvnq+zhgEmdR1E33pQDH15j1pndJOjfFNM7StJB/5eZ5N
mGMn72dB9VLhbGdTgKg9XPvbxlEQsiBKD9o4xS5+LSj5WAMnvHe6zW86vQj1Zbl9oxBrGgzw963N
T4gBDH6Z11dWx30M81F5Oqy3wgkR1Uq1WJEfH+wQynTq2MSeo7PqSrSIiHsBjc2F6pVVrYOnPT0D
k5radr3awBaEHOM30eLgWJ3SzgnAQafm7cYeyDbYKUDRJbzTsxNii3GKsPIA6264D89KkO28/kBg
sJIFboixUR4UkXl9N6h+O1x2wbGI9vBWovnwfivyFzL2Z+Sof/F4LP8k/m5cCmfNRE35OttRtZ/P
T2dPHorCFM+yLxo0wOq4yXZIfqsIdnDW0FMWT531Pva1C7bPc+/wKvkiKyvcZfjREFPRNXPbeUOh
/B3wEDWhfv39qaONZTqNi7wyFvEGUdNQ522zjR01ECAJpjCoORzEoqTbyNQiZEacGOOYWJZsArJQ
CyGfs0Sn4vnKMNJ66Rfuti6g4ftx1pD3zSUvAp84Mr9la5UfWZRzJPAnKncjRyImOfujmsaKieJE
LfIQeYD2y21h0q/U0YiBdnEN7OJki3qpw6WuMSNBpJ9YFyIIWTD5rP99BzdnUf/U+T/5+MqgV33q
IMc3h93CRvW7Vf6Q9TpAriZTdLDzeYwpMWrReb/6XQY0+B1NoWOh3e0VpBEKE+cottcIcCJfjLmi
ohAdCaEMzu/EMivMjWvXYnE7CiIWKppHhGtp4/yXoZOvgZugHAbONagZBZROBb5Rxmi9LvzWSZp7
j/n7EompFYnYhyzuE/mGuDB3GXa24Xm53V04IZBNLJ16hhdqt4FIieaUV5P5z8uANHKiZw5KrXVt
fA+pRfeHBDqUq7aALk7zwc+mN7n1iaXabJfv8Th/xr1qwQztXJchSV+HpWArihRaWNCCZ8GUngQZ
lXRorBZFCqrfIxEVYRjE2rJWNMYgxaAzHBO5yMN2WJLfvm6B0f3tDWLpc+vvFzi9O9h7m+sUwsYq
j90JoJLkFIH7imRhXRb5psMF68Iisnx9ABleOwdcoZevGSEILPeCbhJxD+S4g3jEzYv21DhppO1H
t807ujkxev+PR3mdu7iCMbrjv+FoKhaKw6WbPsuClwFYGLl3QnZc1a9HhJlDrlrFKNSiEkZmKto6
/rDNkiTRPVuYCZcgWjHQk6L1o3xWG9vwB2OwpD65+cXC5Ou6izp8oYHSA9CPMaMgmSQSqWQm7uIF
emaLh2/qhHKZhvUAoc+nea23ZfBGeb63f+xpTbwRFBx24q/9pVb1oo1hTffY8HkBLgZZVNrRW4aK
a4b73e7txPwbF8U7+cn3HF8mc4DfPyVqVhyc0P+FC95NuixKGmNYXRzQou1y+RR9FWaLki0QWZUE
nvjyIWreuvUwVYaQ1BQUxUmQ862zm56AA6QDgCvmUcubm9yy11daE3PGay8dHHLJCg34oMSMF6jI
i+HXUcEoEIi0JaTjQN4fXzyBtA/MnXwHr+ICLJRGHW0ejDrRvqeke03A2s1wL+nnjXGcpcpA35eB
FfcaduiobBzwruLVv39sCkcVNXDvQ7SnrSMk+eZ/13N0IjgDTuw8OJbmGf+XxpSiQbJgy9v0XTvL
4TUZ79D0rbN3x7r/adhBwIGcTV6qoeVBuj5CxyEtISRLvnr+OLg/jiflxbHu1S7Vyqkgat03P6qK
dU8CALZEixiacIoallWHrKogcvKAj/AMiBYr605O9DKZgQ/dsZItjqrLk7aYQSz7yWvxDwlNX5e7
Uqxugzs9AXPMy+/LiQeDhQGWVp8lXt+pBKcI7ES2RERd7ycp6vSuXXvcp9eLcBLaitkMhrjGCMXj
6tDNjY5q6ny+uQ31nGkhkfRkEj+ShFCllAYniybuACfNMysnO7kCvmc9xdohYPWLm7/fHXfgut1Y
ewL3LLD1+mywCB/ysT7wQLteXdXuXmEluMMYDQeqgWAaEWChFdLq8AqQ3E0hCC3EPEpAc7hh/tIJ
GvKEX8ubq23AZtpXpZJNjVtRcGSfcxNPd8ESKv2yKDNJ3DdYKCYkHe4blNn8K2Oc8i/3Nk8VmANt
4lrjh98hb1P4UhLYs7ThOchvE+6jeCFdMyp5Zbfi8CoeMbiqpeZesI2V0vf/BrP8cay14tu8S/99
sgARa3hYjUIS8S/h5Q7v/crjrehWgci1qbCDd7peYS0GrZx12T5LO/Jw8OCaQ/MulR+1v2WdST+w
QHhLy1AwbNA9l3b6afLCQ6oK30AfyMzJ5ZWOAsAa62ceD3buS+Dy4Ry76nBqWX6oEXj0Oitva2kQ
Tj4PnT7buLBsl9Y7E/1GaYXA2c+lMSiauBLGJFMizRgdfG0o4ztjmtR3OQqThyDLxWGKrO43xuBB
p8EunSDlxOou5+4WAB7B+71gSiucCyeeVndeKSGHsdBZnnqO76WpS6c4gwURep6SL6NjLO0bE933
ooa7CRPvz0wj4PCJfndzn2/3uuAA1S3zNmiyhiCqV4D/o++15zweQ1j0oK+P0NqHRP+bBAcDarwu
XcxKJIZIRFctgNqUZWpqnaSTb4JbT9rlSIjEuj4YfCHf/UZhTMQPDrmvsLjBbOyb2hBmi+6D6EPA
Vo1uMlg3EICoWjOffV5I9u0ZQ96l2ZLkD0Bx5XdOgXcAQOl1egK+yhgCyMLPbqz1O6asHPisOnn6
F7nROVYXG7hvbcsnSwetQmJKPqECi86LbHxyw87LdoSYn6WtKD7kWqSbPQboNT6mFBsR0u5hkgpo
pBMmPHRftiaUy5/2BRyoq4q1eU5F0ggOdHgWSWXJ6PFE/LzRzxYnEVhnmr1wvz+ewGXs6KuLn9C7
lVMEs6nuktQcvYdjqxkHn4QbnlTJHPPlJ4mur8coAd726sJlb1XByZ6afbXJeBRZb5DBrBPK070Z
1+NlKLbaifKtvhQzlQWmnRz/C76cNWMZgI3wQ2aYFkUdphBt8twKWuXQVSN98wL2zEnUUkGyEsJq
Se5tdQKWU61cERmA54o/GmP4ip+hco2DrNYogqjqloqrs7JPvTzd5ubfdfVfT5tJeQ1Nw3BT9FV5
1AYWn+PUdg1+F7P0NWyXVeJGCxTynOqUooemq7rcGJD/tqBWDujjqKP8NIjmmhfGVNXV/F1w3gXE
MCIahyRt3s8tKynIpR7JfzbTE9GH687C1iph0mdIjzjw7geiEPnl/K4/mw2yf3TeK2Si6SWODuX8
W0h74jRGox6tnDKm1StQ8MPN2A6wG+1Isb4BYQLXEDyiNI5UXR7TOu5XQ+LBbcki3X2tCj5EuQ37
crS7kbbmF2QeSF/pXrp2CvfJTlwRlU6T5haIDRvTsgJDTdlShcngjt6yJrHHdNqJ2+Otg9zS+4ZD
uVicj+SLoVDIIUVmbv1KAQ51mRVyNq0Nm5gCBdjim/h4pucOPjsOULGHb1BpOWt9IHDPK9HgLQiH
zB5gVnMBYTwYHdtn0D1MeJUNU/H1uYQGEFfC0tfRz7h43klGoUzAYlHG5FRPE5yozNBjef19XIr0
cwpWQ1FhJ+DE98S+AwdYy5oBcEZ8WjVvLnUUoBmH62NGw60Xp4QhjounR4a8SpxirfP8/hnbBW+s
8MFYKH5rGIIrlRlOvTWxv5kVU23h3Iml7El9A7y73MKVEmielRMxRXs4iGqpFDGtWyx2k7QO8zsl
6SSFYGIC4vfB3v3tiB1BKI/GkgjeVzy+scyKfnWYeVAGS8p1mhGfz/qfxeN8wJs10aisGLvDE8HE
7ayn0fpBcULRUKeHXUiBHSDr1r9+jEtyHCT91hdnSqbl8ttma/arB25BMTxjMkkz2PUdodbyaMdK
G5fqubOmBugk3xr0PRsfAUpBBJlXy57nyhzVw39g7k2jsBNv9epAMZCZddyhEeTPEkww6+HmrhG/
ANeWrQS3aN5Eo1SqG+kJ1pD7HbsI/er+YVRPGS6HCPMc3sZLNdtw2nMBCtZsjr+8P3blocPWWSFo
7oTsgvZxwE+mQF9OeefCyp3n0Q7Bptv9mmjuyHqwVoFcsoOf2yy37ZgT8D8roR4GGUTrOjY9qrJG
d8rqYHNL/IuIxMJgwcdF5Up3ajj78wMQ4H7QtTDfNYZSDB7+5mBmqI6BP9EApDN63hNEvj0d1Dog
PtEuw+1ZUlx0Jz4XULjVYv3P/7AkRdv0TcnQ2TwsbAkR8tGytJPzZ1Rt1ITpgQ0lUpx8pUAlj68H
ECUBLhfbsJcfwcVNzt1C5JuFuQorqUIJ3/Kbl03MPG2eJD8+BB5t/8lGA7rrNKICNO2MWOMq2ReM
8plS/PDIfjNLoNZ+RdmcUdgbjeL5VF++H/uaArozwRERx3YWIJtDg0KQYwwKs/5/QG9QL5m7PGmM
mMoUGrP84LU8VX+83i+fv9WVhalVbJ8b6ihRLjXdspExbgSFirLKomj04cmW3/bzMjCyz9eKTO9v
3K70lXczAC+DFY/ZL7ODEsH5kReTKZwE6EzdvSYwhId3z1LHOW6F8knpcBnT+xnjXNsN9L0da5eu
RI3RVZ4GEYq/6l3fVlSiJxSdT/qXr0Of3oBG4MRNDAS39v809X4M12Q4aEjbuHr2cvmUnI55HPus
ORurIcoo02KrWsv4Tx32rlmhuh+NetoKPl4+cSu8fejAxZq2cSgHg1fdlnxnGAUw3ZMPdkI4Mje1
GRxj7Q9gtq5rMCjHSG6qVJn7I1rWadzYPmj36FskbAKoMlyET65yI8ehFMNhw1EO//7I8sfbymOR
lErsNabjXx+IA5Q+a1ZRU4kdwDtDXjB1vZ0p+ulqJW33PYBuCL56qMid2PD8iR4She/V681Lrpra
RpwxjIQSeYa1tcnI3EMfqNXL4QcTEYRuTb40WA9jx2hbrzfkyffUrGXsFie24lW1OcSezVoPtEXD
7VXOrNwV3Z67BlmT92KLT1u8wAcyVPJrUbomJ8odMMdSOcX+0KDwk+iVcgv1YB9YbEhcdJThjcXH
6YsmEktoRMifhqUTkHqs1fk5Hrq3cHZNju45YV92VZn71PeJKzqwISKIAa7T/LhwHZlrBsxLa4jx
bpee8o+uTBqL23yP0Use8GaVd9D+lOL5H6qAG1pXtWoXPPM/rtgwZUh3+9M8tC/EIcp09lxmBmbt
51ZWpb1M6qoTIzqjmiGjOFWqmAXoNhGPVha3dI3UJXnix3wgBnKP3N0xWesdUJYTXlyoFv5GLpYA
Fl+8hUn9OgwnIe36WH2aJXTeykgRkJ25BOaP6oAfiq0Ea7j+8cheW436DpVFiuhu/VY5GNTqVCZB
QebBW+sJRGclZL4OUITo7Ovcm+A7c+PzXuZI7Qn6DxrrLIxLLez9qbEWQ8petyD5Giev3BSx1VfW
fV2Qt2Bug+32ALO4wP3lEdtLMTxZgxYAM1tWI0DQhiKhcCFP9fyWXgbWhz2UcxvIb1GdAerGLJ+7
HTv04GphL2jOUrtzTERSK+YMhbXkUy342ItjaJfD0MyM6HRoxMLKUxF3E59+fVB+AznKJWK6Jv/S
PsJe8O084jvjo6qXxHSBdUGPDYVn89J7T71O8ulYZc5MkiaLT4XCndazZmRtxVuBBXa/ehx/Uhuu
bGwQuXvQ6e24SnScvUJMdPajJ1UEu2qbv/W2L3YtIdeMe3RPRTJsc4j1Cd/YyzxTm1KiH2cLy9Pa
AYuMoT5KeiT2or7DIXwc1OEfQrJSgOhxytzoL4VydNVymCrBP1wm12wVkgc0pmi8QlevHZ7802Bo
kkP8/g/TwwGvIgEXhKv/M8YkwiSYxxmPMlO00dm3oxj+5M2d7Mr5RpqYLoo8n34DMFAGLtcnp3q/
pB7qL3MJqKyoQI13ubF45Zyuo8748pIOn3O64zz2twR4HiCrYiwy30qQ/vDg2VsW9aJgQY8WsV2+
yx4mVjs0o0W6sNfGvuPhksVEVddk4HZ8INhCQQMKsiyf3BZg+mu9G0cg/Ii7rto0yoEvdshiI8CJ
8kYw2fgB328L6DvB4vS9MY0smr6QN8ZX+7jMH66Lxah4muu/BN+UGv4AY3oIo6FrlDefjUlAijRU
JDOUHOw8mtx6QBFb4iA+/wMKzoRm10ZY11MKPeIOFh8YDJiaKmLSQIzEBG8x9Wo7cSR3go+ZbVFD
Z3zFuHA1tbF5tHauflKUsQYNkyZqIR7Lke8SSmWXu/9R6IGWgR502QF2z8RKnamO/rymCUro2EY1
Z22Xk1hHc7GDYvji2sNrlSOmQTxwWRpX+qxUvT3pCSyLYrz+ZYO2DEgOa4fYYsy/793snMYl9VtV
YzEVfmhpLa6spo2lHIyp8oZt3oUqC5rKy0J9nfRyXc0tR/VXshETIM2WwlGR0+tD+T9RfUvwWU5o
dacepuMiGBfT6waabUMCZ0gp+FUavIwsz4pwlY2qPjmFB54zb0M+eA4RTfSQRxJ5JcuALGWK63h1
+mAT0hH2el1xC2LplTlOe4esH4oIZhj5ewg847dauGjnmkEjKVG1OdtdY5L5SOCqvj7srA02U/iE
YOwZupcOvtFez7g0gGfo3388sm1ttuN/N45RIo+ZLdM5mYoxYHs98vW2fyaz6xme2LlOmtdsYxW3
fcSZ+iZJq6LVwWj5PAH/3cZ3KZRftE6MiphWVN0k6369XHxC+lloKDRglgqE8JGd63ouLOYbRg8F
T0KnQNihi1Sp0D3AISk8A1a+U3A5cd+EHyUyp5oK+s8PglPbprjSU70GNsnFjFWMrmNJbieVZSNj
HaSc/ecDQDFfV2bvxwCFnA//HSU+1Va/iZbJrpgCqCO7RBMf/JYHIaP4Dd9inOIMr9Yd3hc8C/hb
j+VlrdZxJGwEVUokF9d8KBXiWf0v4EN7DH7yCtIx0OcBJeyJCUskk5ByZE55NhRb7pSte8V0d8vu
XiGkQ3B+2I6BWocgORAaUEEXaBEkoELruw6La85OCrd4ujUDXLGvn8RXfTpTniyv5h24aral0nok
kMgCKoCzJ+BMGgV6UXoZwpUBTkpYpSu69nFfHkaKhnBP8O86o3Tg0EzTIsd/VVgDMQL0Y/fM/a80
AyqNMxmPS/ML1sYgAm4dL92iIXRvGh78a9zw6z/cUi1i7CYiheM7o4p8wjfl0Q5mG/Qquhd3Eo+C
kGh4cbSmEujmELLn7GBb2M/KT/evrvaatjr7Outy8XWTu0CYJThhCsVLlcCcQoHZ/nYjlPSrIMXz
D9MVGTxL6YWe4xdjrrgK9gHPbET6uEAqV5R1eEQyKNTXnu4p3tbzzdILLhuxqh047c+6UjuI1n+q
SmxdxPbv52GYdKt+vpasjjLuvEmiYwbxR+InJf119I17eKtvNZo7Ut5aq27J+RP3nDQ4FnwGGXfV
jzI8yJtZLaa8kUcdxtT1JaA2a9E3kTB9qNgU+Q6YqbTh29PGG9WijDK5/UQOOE3QSpDPA7He6st5
MXXMoRWOMaVDm+4Z+4klxip2HlDDCJ8Mds5ZxxoznMwPgx9X32Q44LDg70wlz6BcSHSwFNLEDQJ8
duoNiMjstN6gjM/nlznqyfoTGWwXkMHXSZIbi9dZU/zvqG1tH6unMGlJ82vKuOzZzf7sn2OeGSol
d0Pn9eftGNx0d/kdkduwKQfCDiIXcIWJWAr8NdhRYpPt+Gf68ElSa+Q3CJ364I/tdEUMmd7fO9Up
2ZWWRdYt6Oa9/hzM/jI2ffBFh91tGDYNvpxhVdlOYWeMqMTfQy+yrbW5a6seQ1vOvQ853IcRxmoP
2dWIDFd1za8k6aXO4hlgQxTUeF5Koz0+wb6d6iE6hsZPuV7XvgZk4Knekd3AeQwM7e06n/BcbeXN
+zrzTwKs5JNkah0ahKjeEifDryYY1hlMR7X8eR900eRdghUQDOFFjkiBHHSa1xt20tepbYP89XxR
jFIJyGvHzG8d/YU4yMBaSnLIQ7kjcXoA3f3QMQP/YO8eLcWlGkIFK6HZinnNAOrfe/VKRsX35RYC
laq1RV3N8WmT/xOBGCNJONOo04yqefmjMC4EuQcc8/vscvqJzHAo4ruT+cPE7eRTN1bKpGA46+Ae
0uXtJ8r9FRkk4AlyEv/8Gi+djorCE/XMVc3gQxi33ngvLm3R7ZYtsQRCqnAmUJjtPIiDOK6SLktv
1acdbTj6IQawF5c9WkhPkzz5xO9ukhVXxd3FzPt+mJJgYWiMmQbp7hbGCzm302rLOKt8p60fLJ3b
jdRDCYJzrAZOiYxep2gpDCTfwlLD+YesIZSKA2/MRsk0CKI1969UlJE97Sk4URjeZk69TLBjo+EN
PsYod8AJngNuoB21wTiIXg6PKaCbwIu7OGkB7YnipsaYhzHpOD4J8KX/v1PpqFV7ESR+NjS73gdg
5M/47V/ISdS4Yyf2hFZFa5ACpRrZXYAv1y+Ghf4yrpmfjyFbK+gmGXti59N99y4uzJF3h37lEv8Y
D6/kNwUG66gx6UgcrxVvIZ0pS7dQNpDvirmeQJX59Sqgum8PZRPJuyW/3YPdn/5pfVLJWqwwOCOz
CvJv6ocJSJZBgh3rmE6icWti8T8D38VkHVGCs/cXxkVAmDZVlJ+JpszvegtRe96SdLDq67m+e30J
8pklX8JvhraiwjIgKqDUs2iQrOnw44HpHHvLxJeOPveALsEWUZ5uUR1RKgZu1LrGXKJK/8MVzMhw
brfLMMhVkBR/Gm4/9onp1M9xG+t+Q2rFxi+m3BIQpEJmEMzDg7jeKpDlimnzN5gHlLS+xYKjOo3u
H9/My6C0x7UfD3y5N9Fhz9t7akyKBubRQTdwz1oXFPAUj/dLsw4PkleCUcQKuqeZeom6c9uJ748e
Y99YjVgP2a2QEL+AEDd9qLQk92yl0ZHxZeaXGzASxUihT8qd3UBmN0s2Y/rvbCNgy/CHePuAkcb+
RF3bjTCvnKAFo431b1bkzXo1jJ9R0wCTzgvhqjl37KZMt8XoizxFtabyYwOzfTnRh8bGbL2hOLAU
KwaoR+JWoqKR0gmrkeubauWRo3PXPTponH0jg5+8+Q0MGjfdgh49luxnl25ZQN2Jadw7jr6nboze
e7YfTXY+ML418U8wDylOZ49iykr8d99DlTp/0dpnYc7WbwF8adCoXVHgY8q69IUuHZQYUAIYQW01
SIb3EsNgUx7HM2Cxtvu5kbwly8VeamQhPFTruLet7Z8DmaO7i1tnTiwojWpSGOnw5hUffOxvMRGj
DGQ8L/9sBFOm/t5zZZvrzCcKR+qJcrUyq3jcc5g9M+9FAwCe1+K4HVrJ8L0RmI/BdhAVAHqMPmuG
wzQrocF5bk3uJIXCuCV7HuTofiaBO10vK4lWCkadOnofdSQF5uSqukGEtNgUNBs4g8zH0DPe6MSP
W9n5w7yVr1qtiBykL67gu/3xDZgW1cioVyGSdW7rYj/vhp53F07FobUxxNkUb/CNxLf+MQEGydm4
CsmGjTe/xcqCtj2/QLBLiqrr7S6Vuu80X2qL0Mp8YrijmLx+02gfk8Yuqja1ph4nKX2vit6BJ1Lu
BeI1uNeyc64W71ctJL3FsWKUUAxti5U8930E+W00Ie4nOsbt09r4zMpBeYOVV+dELfwVTS1wAWwC
N9YkV8nFaIglfq1iNQ9Fi/P4mQFtcSKr9gzSFWiRkdnD3nU4AkQ/tTxnbHLDpXZ+14IZ04hdto6d
tzYEduSb/QDaHagLQThfEmbIRfmXmGxwfNxN8wC6W7TAU1cUxPj91uYta7DG/99zspci+TZwuTq9
53FJ59vVslw6isvmvcpDIxCahXUWtWPb+ZcXIM05Dpzvfn04oiziQSQF51yTUleF3B1Tsq0HfoEX
tQwiwtmQN9F9WpP3bn+amq0nghH6zqgtZ7l+4xU1Hehi05NxrZXyXbcCPOLCHdkYuRktfXfcxkrm
sBGGImH12jXv7pw6YM3POBIqHq2FYoDegwBCX69vcUuBBh6+X3oHzN5X+iHZl3BouzxQl7lu7DaK
fPfWNPPLyDs87MWtl/ZdXPULNsvOzuiQ3F0jXGTeWmWauMyko0zVmyTn7FStec4KjujugrcJarGZ
n0MVkB/DmSFXdSN8Cc1NotvM2J6i2Ju1vhemaqRhkdlNd8WVj6YLX6RiuWQYWA7KpFHF1ex9oUZi
eOmGrHfGOhH+Sw4Vp3ZXX5GfIM5CPWp4dBPvEGuSyVcrE+i06lMCNZRVJf7xQKi0UfdKtGxbALLU
toW2y2rocffXkGHlChyEMBEnbHesP0Pvs6nFWgV2Ftpk+jDNSkcTWIAHrh21bo0Huv6mhyN/wK9O
ydOR6YYsvVlu7QmgevcvevD1CUSINlnrO9St4qXij2V+iAiiVMVJF9+72gHVe8dM8/x7HStkKAuP
az2r8789pVKZe4Abk9RZDyCehrqCHbCVxg94LO5RYna9dzrYVkl/W7iEP2P1uHntl4ZlOeWE7Sn8
obS9QE5pOWNaXdDTRRN23Ft5rCitpGrTvGCN0JS8CNg4x0QFvOp4qG6OcuJL4pTzPOxJOCiT0zWw
oquVvKRWOEgIOFRsJN0f4ZiWRIaz6dFkbPvXlu+z7RklDpdu7IpHJ3K96kAvDEXWrl4TAz65tSB8
VhB1bJDBcjx+9EixvqTjDdpB09t3P+aZZPatqTsG2BGMZKPYY+C0azLVJnQ4lkeQShFjcub3XaKh
PBJAp9Tsh4kFDV3l/04jpVwEvmg+Pw5LAJwrd4p1pU5IEkhhZtu97GNCRK85DQp2iEW+Ab2SlHYm
hZOCtm4ZRIKqQF3n8o2qEDrxcHkr2c962TUCVMpX6hi5S2QWBeltVNoac35lvVUcQWNiYOKqs7fV
pGjIeaEyydpUaHN8ywXAXLVUCAzQVUEa/+c1wYZz2soUDcn2M/BazyCcjwFG/1AvWlhcFH46iQqB
H0/ATANyQXWcdjzmcJyz2L6vJotnpdnBB3sRsfWKW6o8oSukgwm+Ic/ZIFzFW1JdjDTN1CKmC6Uy
GRd9GdM8iUS1H00J0KSv3iOvGi5UyPDl6TtucwyUhVRWVzNgxGTx6BSg/d1eSQAOGeHE2ONA0uDP
wUh17oqs2KcUwzeweI+eJd1Z+71+Wf9kf4fyzsabx3Wr/Y4IFZm288c4m1rd29mQWi0RbtXgO+LR
SjLG9+Tx0zZGpY6HXOyepyqC4X9SHh2jOJbeszrd6n7u63WhXyVLiY78gudfbw+3CjsrGh3g90oF
W77FWJKrXvFYqQbBg7CTCEYY584Jnaow1sKbgUyPar+kkh/kzPlNcRTgQQjrbR948JJPU6KyNrU2
H+r+iEfUAszi8GdV9A+Tht7yomvXzf78zzp9wMji1RCVn1RiDGvQQyNhNFJ3ARzBFgm5jFRX5YGs
CyA/nnpF7XJ0CT/ALAs/1A8Nhraly1DVuG0qhdA1ZIohBNHPgz7A9cAkWFrdUuidRUYgsrgeK3Re
+rip8PSw8JwdemPn6QJDELeDqJC3iS0yE2YhYd8zF4fuZdAuOO6eO2xmOKUUFfqPM8uIvGJBHNd2
LHfwlxiodtUnvED+RO9iFEkGixLb1HHCnzffWFiKX4Bw0kP6VcV4wZucqRBRB0g20otxgNDp9vfM
jhMeiNJXyZ2whZGA2lHo2t/E1Xn6YtmyMRy+vPJ74dZ+YsH1iBQREKdO9JLMF6BFeBgQJPyDbbR3
kmfYAlI+TO3kHIX4wJeotKaDd2BwrMGRz3nxf8eY4JLPKvx0yA3nhe7wd+8cIzS23HYNkbLq9AyE
5KtYg2h3yQZKofrLoYDf/bz5P6+g8W6hWRw7H3TYvrIoQKaCuTAdIhXnEWChrqO0cty65c1T0aZR
ZOuoD11uwMxsL++7IkFPxLJkwOtgXtWoMHPF0/ML1n7PjfovogIb5jrpej8GI9PetBzebFpcUt1z
T/BJav8SUrb2PBQhHLFPr9E/P1cKAzBCYmfdOrZQPV2Snjh4VyrfPdL3MkQZBd4mfjfj8nbfRtCr
5bKopacjchcpfqSV9m1NsqamcYbnLiQxogGnEqU0JWi2yVvjGexkYjdIQ9aXFITV8Ybc+ZuZRExE
OuQJshnRRO+VcVYFBvyFOnGYXn7r7naPQEPp0Yw8wms+jw4WLrvDGytuP4hUD1St4/nRjmPzE+54
j02H/9hYiTiMCNVW7q3CPg5hgSWnjZXyMrP5nI0B7qszpXk6EfXOArAgAoHv13AozknL9SrjNLZp
fEVhbL5oIR9F7uzD4kzAEwa3tGFjb8Q4VeNQH4KEmYFEtIF0bOs13zuzDBKEjRJfcUMCYDHyjsgN
5W61hSAA4hFzw2wFweJyWcq/8rl3p90NppIs14c7Lh+/ohvgLDh0Wmd1udKRB1J1/eXYxpptiRf9
AFPzwopApWmQLwtnbcBuxO9UWVDTlVToDfUibIWc4+ZV28kpRP59rRrquWyA53Gxbq40Asx35+t/
D/4iOltJiJrW2oXYT/pm+bxayYukyuhNkv7fXx7hIhqaSYslAivr8kBlVEuyswc9A9L7K8/vGygT
5w1dafVHD3KBCUXzjwrxVjqqE2VwziC8j5jhbX78dDBywwRw+MceScGKEFsm5O5IrFT/Mo5rWp5F
JZ0Nk8PuhVI352zvveeiNSzq0anlh3SIBFQSpNeuj3D+uHClBtUsyt01WGWL+EFKpPfIqUtz+x3S
tQe61eXj88MTLWMSSKLbkhASv81RDPcmfWGqBeHXn7L78EqdGQGWuoIjPmBzYxykC4aQiVpRhJJj
q+UZe+HCgaXZrafxLTqW8BcothHImQ7Vmu4Ez9sZBJw/cE95gtsUNGMxq6Aduc4T2NarSEMeD6A8
81Lyi/7VWcZeacEgGi55vazXs/y9bbv2Sh/XdDXF0Pd/+WUOAwuWjJotMMbujEN6TtqltAi7ZTRQ
gxIPGiglwOvet6fOTmP7XKHILGgi3C8aMpzTI9j9uzDxu0ZMA8GuYpCcLqx+H5WPzZjRg14PY3zV
xi9agOdzjfRaYoVIGLQuzYnI7ccUE3uS2QTuItgU9hcD2A8UpZB6hkcjXkbBCBSRMHREwyo37Dd6
+zw33lHsfIT1FPBSb4kdFGMoNRk6g07AdK2BimFGvIgI+LgQujtxk9viZutrGilX2yJdPqA/Nbxg
TGh+Fm3+Chbmx6aSnVICZFKy0j7TjtvaZRf2o7qYSRfmm7GeL++uznuDz03CbSYymgLfCdoiXpMD
yg3omnHVNN4rjnFKX6+gPt8Ss9Etk00TRVN76PjIT1LA/wniKEhpUTo054ztHjtTIqIVe0LgSWUH
A1dOhdTv4uw8IQukqZeKIarTWzIbS3jmNQ9pgcIGyYElDtdu/6Wee0vyfh4nvPqnV2+aL+lmOZE2
Dn6M6SNZ0sGXvbQUuzSw/IMZDLSUmjoWIokmLD9vgY49GvOz+1ySs1v4hK18iq0mfmwjHNg+A5z2
txZeE7rK9GKRNwtj7TK3tnkRlybT7CLDJxB+cI4lEiLzh3HB9mrzUa2bDQtcdde64fCbspK/H+Mr
6VwykRybc/hOzfVgM+AZFsjfcG4Nul0V1KoJOihdXkHOnSbFC9Nf37PzI9sqTxnToGRKN1Edxn1u
fd9dF0xFF+tnwp9mhL4nuQwlffjbKTNZoeU6R22RH4KLyDrfdWKwuqzkA9JQJ9cnX6XccKOCmbis
2EU81eyH6yp1Bpd8nUZkEzTOdPwrCxl7+19S3eM1rK8Z5GIdm/OgRGBKlzS2wOjWGZNY5tWaSZIZ
SxGj960wIdGjvKck9tuOqDMDna+ELdrzrTzSpVVYv1rSHhTuTCaoORNiJvQrvIzSDpSlJSZIwMuT
Kdt8E3WBlDc5O6e/7wQjMD1Q8UAmgbxWr2uADyodTK+IYL6a+w93iMYEdrlQIEVcO4RrLYqbwPYV
i0gS4kpRQZxqDiH3G5Wa8RFHh9LhSKs9TOWdlY7x5KjC6izxrBHnIKZnzJ80cXXcnH/r7G0amgHO
b4Q+4mO3LFhqtqeFE3kVcGvFetRqivqDV03JlIBmulY4SCD5qbv1mtug4JehrsJ7NBoxGo+o4B5L
P+5u/JCFeH/qMiShJiXHYxG6XbjBghLt37YcbVzG/4lLkC0gRKEvHn9JVcLFVpOgrxw5zV0NcdJK
2vBslOp6ekaoIHCYQANB5lBc+jFeFCGnuzdSCSbFjkgPp+8mxVTCGokbK5/Rj+JJAoJSev+em+BW
7o14DgeHKHMZthwvW3UXC2JMpsQ35k0vmWQDykeSexlaFwV7n71i/y4FmrS/jqNLMMaxrQ4FTSeX
VD9wTrV7Xbr1iXKneP3sMPLGmcg2oefK4PIQomtjOYIrddGlbA0nov+OEQ6C342uYyJ6XfPx1bLM
QREKUFm+GL670bXXXQplf4fmMzlXVCGzbSszcdo1GVOWMvsm2bn7OcDWSu71R+JAP2x8GFzHYY4i
DMM1nRP2MkiMAjnzHgPOcMZjJIGGGSqfn/5RWXGmwT7IPiFrqpXe4JAt/lKlHa3jeUg/zM5HTt2H
BiiwcefqcUHCnkR9UlFJZwL9Mr/Y+SuQ10HR/V3VQfrpn4TrKdWbQHBAm29fH6XkIIHPfWV+20NP
y1RADXDcp1VZu1VUM5hJob0LK/0PARlPIyjzRsNLMuyNYgX9yPv7YfRwr36JUrFMZMZbkAzFSKmr
j79qzsKyyk+im/g5aa27l5YRQfTJcRHMegZRNjJ64WVJhA2kddHkDAsXR8EFe9xfO8STDmbMF2J3
S8maY0RqakS2JBdPma5cBZkaVVK2DLa5Dl1C9XwWhXUZ1unrg+fXiM05B5EYAzgyF2UskhzEqqgS
l8DtgSkC9t4au6VPnJMvyijONPSuBfBbS8GYf95uByNvK61orUJ8M10vgjYZc6Iskv8o+fNDGTfk
nIE3HcOwTs5dW/j8UMDwI1Qcnt5lVab/A2+dIClxO+COK6CEp7hyJH76oC2/E5Mn5f11K2A+1Zdu
sG1xF/jn5Sm/JBxm2qMc76gVRWtfGfgfbq2AulrpQXat/cK1KKIppuWHw6ZtIYUGmIWDx3zfMK2o
+AXFJRzKiCEYE8+o1WbGA4wQqk2mba2vu5w8OuYCZ227DUNE2C2lcKXEl3f5rsFLzKuySb2pIkNo
g/wfU1doJ9JlRuI5IGALZsnkQpTN5Jo/Vgi+Zxurp65gykm2F3uOb2TJgprKK+LuxhD/ZXt+YrY5
04DGtjofR2GIJq7YLsQaI8pMDWskKBVA01+SSx9La/mnV7xA+6HCv5ZvKKA08K86990qa4vM50K+
OiCunGgjLfc9CJ9HidACjSIRJjOoZQ5LEwoQxnx10/PJZBjfrc9jlykXQXPzfZeOHQZQNFi4dFG/
n8MG1nNhYcVG2ZPtmqx11NJ4pXL2sZsXdiCp+A7aEXOAxPmdyXUdrr6wenRaaS6oApmVhcrCNLg2
+Xl0ygv4evre24sWJHHGEubYeqOVGVRsavxhSaRO5OTz9n56rLdoyqH/n4skz2JQS3CXitBzKPbn
Zl4/gZ2KmYNXzDFsmTPodXdmeT4V8qBgHfo0IQ54ghevAd20iLr8gNoD1IeW9Rn6QjVUtYdu6SuV
Nl7r5WsyPTemK6/iVElsTchAK4or+W2hLl+loMvN0Ii0MUkLMZCLodyCmrZJuTPs4tbD4fZLFaoc
9hkiVs8o1fuC0VQUfAyBLGSwNSMXv0C7aoPnnWgH9JI2WuYIKcPNwaScsJgtQl5z5ADcRMTyqYAQ
LdtcLOiugBAe3CQmzQc1mO7jpfPu7NiXvSHMBYmS9fadXA2tq4bMvlIYpUtaybYDPqbQ9qhJKZ5G
aY3y8MLSsDL9OFjo0pgNTzEYRR3hbTIeVg7myCdde08Ec14KYfWlJKLk/j73gEVqr7PDYbv2IP74
oPBbGrPCpJR5vk6B/AyHLWp92DWxNfdzZ5sxYo3QCy1g/95/TWbO1g4KuwWkkPrA8mY3jOYc6XMa
1oneBZf1UTfM95wNuYs7b7aBPsLtX6JucolY1W8ECwq7BbZrRAsN8l+AB8Hvyl5EY938SRaYG0AP
rO4TAm0l6WKfnCqj4lvkqCU190qFHV6q2lu+Db0r4HPctJsjawqz4ISsOgYv17cAp9PtbSEZjDed
6XVeL+yogQackiFxl0nJXvrRW2fAQNMHr8D4yNldAXO5oI7KZWUUZkof2wbz/Dt0oSc8HwLppx2M
bXs+5MQuBVslvX1M5vpll+0kmMUK+g7YR4NHB/eeaPGGgwpG3wQ+jcUqh5ldESOOFucOkROfyVGy
MHUWoo+HfEXpG7CNGVcGNjq9BpZLwx2ufTSK4VZS3pNc+ZxdSERftp/vi+9obI7fD11mXL5x/R6H
OvSvZjLHkZX/49yqq+jWZ6iQYf/YfTJm/E4km9lN8xXxg0rSP1Sy3+Vm3S6G00xw/dOP0wITvs3T
xaAtF5M2HDU5J0QxLf4f4wIV6/AC4E6L3pgDQ854J1uV5U/NcLt2u/B2yX4nYNK9RViCTxOr0cq/
D59/sK63ODQ5n6gZh8sNt2PsoOwmqvPZVTECpblE8fJ+7aOBlr2ntP74veaamVSXNMf7DTJjkf2g
UXFoDIyhE3gMt2WJx/TpSnkq1LXuWbN32gsqaUmexHGafGlNaYF8fte2IA5RTw8ABwKoAxnUi3k6
+td5PB5VhvfNAo2SNOPby94BQEAYstO9r4nMiMo70mZxlscJxU9cITtE9pN8Hge4KRDY5dgMNe9x
/3Dc7JNMKQ85NSOLpfl+fa0hwkeBqDNsq6ruzpEkYVo6VMoRGkOk+YUVsylalY2hp653urxs21vP
6yhfdqjWqtBHORRKDHKkDBHqlQ5bnMgQ7FgBxPnh5QV9E1sNy6Gt5DfA/knYVOXrRN3Oni+GoUES
MMVik4lQW3/s5n3Ljn6rDMyRDRPDI8ii7KvPJcCgKPm4vi0F70eSgv/HvR692V5bFkmEWsUEj3iC
i4lPKv4AzrSK5zPKyLNJpNEpjKIp8Pces/Y/Wkw/7PerXHb60UnyboD7zj+IJuKUS7SB13u9T4M9
G12AITuvgNsKqCeIM/Ml4yx+JxBz30Hw2725Brb7M8YPBp/hk8s1ocrGqw0tCLdOG4GTFUosF748
rxHY4ylxnDJradgDrm9klldi6PToxJPUHQ7s7kV0eEZbmZ5P4prmeQXpxOQKbut7DELF5f+f9sfO
9BnqdpEoVMuERDKweYhEbsG9s98cvLuS+CzQnal3hnIM8XyjEWbVmgojww9yOQCOIDGAFT70FVpa
Hicza59pFtKl9/8QdGnqlHE1sP53M5M4FQ4bcWqnLMPskh/sh5glS4PsmIZ6gIxVvpuczctNMMZZ
FORMTD18KBzU2l9xyaUx84RZgjFUAKBaFpzRfnZqYGuw1Q9AyQm12C8CqXK2tH5EXZi/mBwGvCBf
NBUK8VlSkPvQm5UvqehTs5GRFwmurF5po/mN9eS028uv0K3FetRbgN+rJ1+WlOOA5W4Cnccfakql
Z2NVN4/AO14Obq6hXmkiV86iyHOsLGCxVN4VgPj2/IN4AMuJfsWnEsVcgvb64g6NvBQQbyJXY5Ch
6EzkEyc+l1meoUxuFvcDFJERyCULt8kq7ls5re26VF41zoUIT/zjO8ayxalASb8VFngNg5B1riJm
vH7StjXYHRe8idGFCS+PAl+3lJQIBYm120AAYC78yIW6RocRRUnGkOLN00AKznlBQIzyZlkeUjrg
4DjTIZ+0vbR6cZm3girhsFGoZmoxZvRv5IEoLbkDbQvY2Nj4DM2NMJmh2h6SRIZam3V3rluNYVtx
pw7BPHJhs2WnNOo2K5dXzRXMAvbFLoSPXXslZIojPX7n2cdtUe9Q3npHPc35AVM5ZoWCvUknVKQW
LTw/GSvLRq0wzfrq4js1fnyBd2uAYpvRw4En8eTn+beYbrqcm3bomnLDugBkLZb/zXfbd27ajrsH
OXFalN8vW8xC2T1pSqBeoM3omPPFdwtZuKpdiq6xjMrhCCQqvhyRHRtXDSVC0nYeOxjkkbjX5Z0b
xZjcnSV0u0uXNzVo+3KHl1he6vpzIxqUiNOtobJApyrJapUyiJYNpRs0BXB1idLe9qVS3/96tEb1
Rvt/tKN1ydTWf64U+bvfji4ouKy3tBmRQRhsc2QRdmW3J5RiTHxq/jDkUgNFJAX/YeJn9cbJUUuH
MjPGUTA1/DcVkjpey8puEY7VYfQs72uP8RNaisnjNcV1ju+zDmSxdfZ6B8ZUA61ypDfdZCSUMxAy
sDKZbIg8xipU9bxCaI6TQBEC8yNkvzgpnvFFK15BbFcVGxsgAWi0Qcbr8KZofo0H8foofuYPiBtS
gV4R0K5CWXQutWGFgs3lZTtfqFtSc+NpPwzXx1OYmVISK2FQSaJ1QBQ29/cuGamlCNMUhmDyIW+D
9lkp4P1l+46//8zMVjUa+WN1ZPA79JrodRYXylty8+Ra9H7v7DPMmyoDeL2qNIzi5JpDYtlHPPcg
oHF5kFaJOl8WZMyB3812WfQ+FjSGEkhW8nMFov0YzvqtwjSfrsRZqQ0bIApShL5QWF7apnVf6PDU
LvR0EZZWTg313i0y+YcobG5CO9t4HizShJD6lxDRdvpF40QhkExq18u2RLqY9Y2nP7GUdlgQSlp4
c5ryvoX9+AkdX3DfIfzqaGQK94GX1K4buTixTePhzJ01hIkVEbNtr7XZtb/7daBBLVX1pDh1rrIa
D+8goRyPJLR/He6Dw7Ellk3DrPgkzcPeYtylWFM7st+22HX81NLtFIBUJXMF92wH9aMDN4E/WzYL
vbnlfHYMtMWvTpxj375+FGpj1wHYTAVPtFVRANDYBH7K/jIyYMnPz94/dmNyTvS8020+CNM3x/3I
xua5IieDDwOYtZMMEe1G8zYAu9qmorHN2NoCZeAH7gttXDlvxP/qHDl1OMf4gd/piH4saWtrtLhz
FA8CktCDYbafr44kf6JNYo2jgULKF4r4DIpFNNwm8rtsOUkbrskL5JyoXdp1vfT8qw89+p3NJs2n
tFXzpOnzgkWy9karVBpQvQ7b9u67V7Pg2SQJoWwiFeTQKLf2V2ybWbDGRXYJBeZlJTExswHAjhIc
1C7lvT+cMTZ2WEts1UmYKUfqnlRbj2G6K/o71enC54GolcjbfQ2Jk6zsYmLtOCjSzNsxBskD7+oB
DVmLbJahjBpPssIwlyvkpVR42KtGQ2UEmAFGzj3hi2D+v/xnRkqm33Mv2jq5QeqBNGR8iDsHJRco
clEBrvfFnu4YVWgttRhrfuT0InSzljdIapPHdV8c58wxkshfi+96mXYW8Dn9oqbJYZ8XLW6lNM5M
dVsLZkHM6yqvuqw2Ytggg8rcIsBjAnjncHEvMX2iPC5IvhpMWpTIjYXr04FAt/GVQu/ujtuzMosP
ryp+auTLIo+6q2r4+3AgdNKgokPKNlataNoRPY7szpuuOi2lbCCCeBM8aYvfTIi11htjy+l3GylZ
zz03py7zZhSFTkHCwMVnRvhwhqGmW2zVZ0VD8M/CVTq3K1CgL0sHnN87CZlm4IuiEk2aZnJq9wHF
SAoI4wWFLVYC00CdOi+tFwJmNWuHP3v5IkHmm0uU6C0S7ef7GT0/F7fcEbkv4Qp8d+1/jyk7EoCP
N+il3zc9oGARAbcOpL2qIR64d0wRlyGRDbSNR1r7jaQ25H4bqGuBPeezloMWmxX872itAM8IWFFG
bB18t+DJF4JOvyhWvj3oXHSAIO1PzUAV9epCxTbjeyINnnuNsQxrXWFEnL0zFzeZDE5MCpbHUxz9
MJ5zLMv5+ziMPSEQ15jTochtsSfDfpRzNqKn7SaNVV5bUeMSTGnPD/Gpb3mnMZyWMiOmgEFnFCSW
xeZf7zVkswN0I06nRYodyPFZ8+vt7XAWlnUGgvIpy6t4FPe0Zo8JstYiMggTKea5YnT2jC085Cth
Y2a3QUXAnaDh6NTq7IQE/WonACRqQGNQl/+MP/BJdYnAhecD0wzvFuB+/6siOP8bTiqpmolTZw8N
RYrCzMWABoT1kI18mqdd3AGWBfoy+It3lLkDe16GJKOUNM142xGrOyVKGHAbmePyLAHpa6wySB94
dThEZQTjubiDtehIj2ReI4f0Z7TCrAa4MzqL9sDPWWYsssQ3B96VkIXWGO0053hO5ecjXknkPhS4
35qPQ/sNcNRSqxLMFgGvcfiI3bh4yrnpMn8I31CBExQWImMzuqc1eYQAKXgvWjFv4h2ZhaPg5E5z
LE+yM5O7p/3FF/3Vh9BX/eZoEfr3Xzx/GxWDqqYepVKuLiAMDqCtk+EUj4b5hK7d94p2rw58VuXK
1Zp+tjLeVcIqiGy+BDplJ83UMCDc99L6hyOqFsizUtlir7wudz00ERUdOvB4+eegEpYCnQl+hRH5
U6KcZIFT3q7ZlV1hqLvptoVU2uLtEZUcJKzWXRYwAXBvKPgAc1Qqc3Q1ba+MjHgh4hA7V6MY3par
Pa6fvyXM6z09wr/o4We2AvQCjMTMGMZ6FXKr9iZ9pgAraSLDxM7VwjxTdY6lIVJwYPODmM81cH4V
nhNVpwQiOreozIwcCqPIHQdvTAxQ/nip/gDkObcpVYJLDE3LIE94FdPYJJhPAAKBLVHFU3eEJQNW
8L0CloZ20GbTbaoes4T7NK4KnNmQrkL1LwoTsr1zsZhmDSKPKuhEJXSZxzExDZFpRmTHRyWmvYbK
cqmxrgmPij/rpNX1jmjRG3D1QchQTLkdERGYg4v9jvo9cBj3WaKZmg6hH8k8D3CehbboERDIXvgm
f+JOW5JuTjlwGOMSoDUMZtXQ8XqVL+taMYhumnS8zUGXM5hFlERDavBNQyDe18Y0Ns9DdL0MVros
CAy2uW8CUGd7NXS+wC0N6Io2apn7LWqAkv1TgNEeg92c/rXg96931aK34IoINoiBmpH6O3X+7Rnn
yOUHgGIk0XjugRhi2xWQK5fVRp1CRMZC1Gg27tiH4TiWFS9ovgjQeU3e+N1jnb8cYwFWZ3Vs8SFc
1y3N6lTkN0TWJV9wJlCLVr+ega1LQb4NciwchhcXPK2wMcF4ZXe9Utjd/o7d473Nyr+Bc0EDj0Kv
p7T0QRlKGyzGuTk67xZ1FuVngLc1TwzEKZXLEELVhJPneVACA9TSogLr9QYSc660mNhorkWwtOeL
bvXm0CKu7CAjicw8yLdBUHjZ5Jt6zHMpX7cyMU8FrOgfsX+fWu8kuuYEZpH1KUYg+3m8ouV259ZK
8DD7AuoK6n/JRQ/msRRAutV2xd7VhlyfKm+OBwReKeGJSLfw4ouZBteJhaSbce2m319/V6hRfZ4U
zveV+PXxfWc4nGV5lCFb8InWBcUmnaL+6hmrv7NPW5ntPpoGo3T0BiGyFmQgoyD3vao/lQEW0kA4
9vWqX5fWfc/ZA8xd8pWq8Nt00VEJRHWx94Y9l6A8nUMSk08YhdouNxNDXqc+MlM4x8YYknjpOC2B
ZyHde98JAz+haLw3FAVt/rNCx2nSnJ1t8Wc5STnUV+qXyJuyYpaHTHYguzlasaW5ngdZ4oeWrOvu
RXTYUHgdu91ToShX5sGAJXX7y3QKK6cxUnbQ6eM7yE9RlkTYIYvKUPW0USEarnufbQ2yrs0bOC7n
vt6oLFbXIjHWegujFvIj1wB2y5z5F/7z46on0jeDI6e+HVbqiGmnXWuf7JU7Bczy8KjqcUSaWQZw
N3aQpyNB05//IpSO2Z9bnpnpWHFawxNmRJk0Ox4r2LJQcN3So35QEgZn5WFc6cTPlYcADZjqkBhJ
k8SmO1vZLqwwu+48lTim4fYiaZ7K401Q4NcyPYRD2acqjcKLto/66m4uphdhaMv/pvJkxRHVeKrf
2u1aA92l/dhrV2hNQt9jIMNvmYqQvwXJ2TChRA2XYxj5pGfwBRc9sC6fDLmphifRu1KXSL0oY/Z4
ZwPsXcgNXbAhnx9qSvcF3z7sSNnatnvk4PwEh1kxsNkbLq6nnQBFxes4GUScWu+9bbstc0gKM/EV
07ANvJiSUmT/E6nRQ1HqEGfthQy5SQ24mehy8ggrmTejs/T0OoiOEWu/matrKUVxbt/e3cjTsoyM
qRUb472yTNLadxmVgjIAeGKSc1WjMFKFoVjAxcoSMokS3pod0RRUSpL1aNT+DS4aRcwFIdZZE8b4
Ia385bSgdOBEKtqRQIfmH/chLwjnDIQWoGgjSV5qdZjpmjSrr0A47gnJkf332ymdfiM9oAsOH+Dn
3sdgfZ2Wal9bPOcNS1a3OpHQKgGRfpzSZTbDN3TOLbBVGW4o0yw+J8X4C6wp9r07XWKQAO30fM+m
82BS4q/gkxOO7515A6NYR7DqNRfCPggRaapHvpi9U1DjSxZPal6hK2RvQqFY3YOR8aOl9+yXjGDb
cbrofSRlv3fPknZXA+AvWmbcck4FrbwdJCssdP5BztsiclD49zHBe60BoYDd2ITXDL9kiFYf/7on
0VmFkQFQAjTSNHi09TprFTj87gtUj8m3U2NODFeofi4jJVomaqulHqmRl2bN1+EdV5BoNKbtOlBf
fWl6c6AgwtyJdz46u6dbmga7GukJBkm1dupNCP6DLw3sHreOcWOgcdfdpPC+Mb2APrnb25EBV0nq
U8G4e6bn8antVhWy/VklK4moTiSjDbGhG/QppcPiXL+bq+wGDuJWzSuENUkisW/q0ttnMctdnVpD
GPcuBzsxcNiV38ND9zxqqQLcdHmzs78Q/+lMju8Uqs0kZKxmczJDMVi2ctJK9tclFc+McOPuP9/F
tOZ43Mmd6N0ILyt9L+45Jo/AJui+piXSZA690zy/PNZP6GfPYczYb6TllD6Q+td4v/ZdBDAx2ijH
e+md7LzSIq1v0yxT3Mpn2sRZeme+BR+5+5PMLD2NZkCeJ4PXpKt4okqNgwZrvYjw81NVl8yybJig
D/JHqYaVGSh1KlhwbBvwKH0rGnwM1+fr6pEct+FuQzM0pwLTEgUDSKZm77PpMvDLw9tk1qFOa+HT
p2PMYKiaVTGi5HyltQkR5uoEZADgYdCJgGZc71LrAwV+D2eR6PiaVDw8tNvxde53WTuhN+jqfRaC
aEBWm4Fr0MS0w0/fHLYH7VCNb9zKLxmHnKS4kTRWHxWG5X6RlJgWwdS/Kujjm79b/6dJhFrNHLOs
QwN5tYl+Cc/nKe3i7tdXhrlDN9CvUMGPHA2xpyyI0G4kwv53q8XV0602IwPQa/D2K+x+oO2/bMDu
wiCEMtth+WOco+ZESTlWkmIywPxgpdPbCRlOz28rtzqI9W2JX5V5CJsoUwyTYXbE46I6QMr7ywj0
rsJQXVw02hz3OKKj3Ov+2buoXBdIHKGKXQ0kqZ5lCrIp5kDnMKX02rIXYMDGvy5rwqc2zAgqqvEq
o9qMv6jZ06vXOXxq3X7NSCO9YLsMaz4Px6Yke8h/0+mDyacislL26sgwuMuZwRDMUdcnkSOlN5Nn
K0RlFhnmb76b/yjuZp6oS3LZihEz0vxHO7PraM1qGUVwtE2T199wFrLfZkETrNiJI9DRaAA6FF9b
6YM1pDBpiy2Sys7J4JUSL16nZAjritksmogLDzqYCBSg8GHrOHGDv/Ulj8yAkokHbSoxH95FW359
fejFegXGEiP0xQ7ncJM388flhyj4/tx/NE8pI+Su0pV9/DfIUQB6fpqE+rriQpncWV/EKJjTarbs
esdUuHmG2mEqDepN/6aRjTMdGvYvexPM+Ryu0QuB6ycgl6cThHvklmSgyQHO3MeOOk7CbCKclAdD
feNRTLbvtOAj90GPFdjBD8/VTBgFhiO1flPIKOH73kzmwHCvKc/CMMrwZSWThqGozdbJEw/oB1sC
GcjarktXnkyOyyR58QRJJus3F2iVIhsRCJd6DQBpPObXuszkDPepG0Rwze5ZQFNAehGDAMR33UVv
g0u5dQ8Ofu1vBjnVHdWB3y/x2e34VzTOgA2BYW4HbHZcCnClKoCZKNrMmWdWPhZVVIcknvI720SV
SvFvNWD9hNFwkbfslZZv/+45iYxSeinWCfkGV1cSxFFUCmILx7dI+vSukhQZPk0zytnKgFJNCy1O
h61VhWdOlqdpEoFaOlHrv+u/sRXKy8IgwBp2H0YPbLLIZwEJFrv97ERYTnzydtfkoNjc1+CdBX60
8ex9969eN2PnPB7TkjenKe8a75E+oiDCgmzDV1yHSwzy6EWdFEgEm/i678BcQ1+yGTN71vnJeH+1
F8Ukr3DK9h8jg80fC/R8priD5hU8nPHNW7PGDdsk9EoeFK00N2LuaejBmVAwrgO71uo5v8Jz022n
6t3SmwkRdsxQ1jleHXySS7jaA0ngAWN8AaeIdT/qcS6KZhU+7Eov/k4/rKW+hEYvPbXynTvC4rsX
Rc6EFiGYjWJM35DO23fLKLykED5HrE5bZjW40j1SN1YH/P5o6qLdP94gV1nRwvR2Vjo6FijMDAcU
GhFnT/3uYhtOn1iKWOPZQaZ8t2DC+/rh8WofKR69CtdqiP+YRAWrtkIRqHqow2Zaaaq0YuVIHBMo
AWH/+ZJJ9wBkBXsDeTIKkgbhr2BGF8Tu/fUT6bg0acYWzDeRHRLsDBoC8sydk5w9Nu3GF+eDcIC8
kWPQMpDItYjo+lYQhxhXlr9t7EmjyeMsuW+mi3t6ZaoS5y1E2AqRcVByLTZpJrsEGt8hJpEn+II1
TVd/AkdqJM9I/YJPW18gFr8sZ0yPdJowhbv2E5LDJkFUoqKh5ZuNNHdjAolCSUs/X6ZDNLiBW967
FBlF357M9Yxc/1ZTmcmC2ao2EEC+P8n+bV1hjGKpNJ+Vjw4feyD7qIiZ+5KggAzupFflaX1IgT6B
2w0b8TK6yBDzbfWEd1xxWpAnyWWpZ1PcdQ8SWLv/eSc0rzSC/MxvpKFNROuLxymifHX78Apy3CXh
VwLFsnO4cLDN65SDkf4r82uQhKI14caF03Ff7+aWSCA5Wp036qwPaEft1+tetmtPh1GKXYl5lwpD
eAVx/+6O7skFzSpN+9DRFxJRHM7STybwv/OINOfmY09liJh7CNUm1QJj2QHWPuXb8VGKraInIqsE
ebcnc8Q8uRKsItlbe5A/hJnWnfL4KQf0OuBIVAsaUGAN6mdf9lH+g9WmEgyKeh+h4k0V0j8iW1EJ
KCZHgRhZ1PFieOlI0VujHWR2Jm7+XsDeGmIZS2uF4j2d9vyOzPfoJI16mAlC557kBihEyupitCCv
b3MDc4Kc2taC62zX6IRKUCnGvyiDyPg70ke/uYJTEId9Ey2vZVoKtX3ERG9xk+ho76hqSixVlibD
s+vEmjs9PUEZmuBh67V0y50PH9phhdfiIIubFjJE2H01KgBb8WkRnYhR3T5aNMXpuP4SK14mafrs
jirhHikYNjaROtFhl4ZvWF4oQfVQMCmUxz58wkxXxGpsz6L0RPhzk77tDDeBjLYnCnbfklJQieO0
gF9Ig+eHgEh4fmYswdFP/r0C2wW0u7MXU5sH3jW8PNx2Ygjpfi1uPNc5vxdN+W5Rng2wvLJNdgH0
bNXKhcf4NMnR+MdOa5zBLxkWdykdOg33Dsi8TIqPjLlJQmFTc6Cqp2F7OEw0Lg4Y/W6XkcEjsVaG
TGYT65lKzrvn2IQIONuR4TPiJqifYd1VuSbYoX/2m6+iaq9DG1InmV+NAD05NVOvkVK56b/D/SZQ
62JAZrbBH762yeHzbKM2+E8oZ/MbpNSJXLbVD8YhQ3txtb+TXYOaYEEKeaL1uFgyOvnzOgN2NZ14
+ZMszoOg4K3qwjqp+Qqpa3ZohJBPSw46S+S5wHTLqN3Kpx75LOY01TdGYXAyKMK3ewJS1z+CPw/I
owG0XVjiU11UqOrFFTk3QxeH/wVduH8PTdvFqolPbZ6HakMNtkIMgVh/t73ihxV8dyl6KpMFuAcv
E9TaaIkOAPkI0P4DOGjPwiHEXmwDoLJB0Pv4XpBLlfYWnqMVusDehozIvU96dxW5RxvGyAwRFXNQ
rkHxOma5mEHD9rE7JMYYkE3Z7kId6A7u52EjTf3jQqi+dxwuUuNdJSVF4PkH+fbMY6+ggch2bUSR
PHXHe5BogxJkO+0LtGe61X7frEv0Kz1XsWxrseNUq8ap2jafJVyBZFW3lFRVlRFm6cG7Eyxis/Me
9V+R4Bw7ElUwAwYOpVyEetsKK8HqsH5DiB1UHnqWq15DgmGpRKfNCZ5GEfRb/jJhxhwoZF+T6h2i
btWwINO0EaHzBAU4ADov/hvYzJrtcsr8lj1u/x6HRLO7BxsT6gv/Pb1XwWOvxcW8Uh4zVbs+nqR1
f69EHx/urkvXdsVtBcU2oMDFxdCkg2c+8dQNt63paFie1P28T5aCk6MUBU5GLnAePs60CoyRMws7
QdwsPFwC2YYEKx//JYQt51J5Uk+MQzyi/k6jg7scJNKQLOHa/4AcDkAneW+CkfqMGoi8mfrueTQq
t6zafx2jHwggWpuG0PDdaNuQURJODTByQAD75Z0ur1g11ry1uv/brPQ83j0YTEmC51cdRbZZe+Jg
2aHoS2NhYEtZAqNlSMJPis3eGRj+Vw0pC2YKwTZY51RROx6aabtcQ1ltogePGmwJleEiPonmCF4Y
kwuSBQMAvYipMo3+qOCYBtmuRf5qNod/oOh5lq4EE2NUhCxa09EQQFfxAgIfjwCk1x97aUBM1A2C
nntaQnyY/Ue12Osg+FBKwNDYWxVJak6v6ry1+RQ/kWm878j+lRVisIIJu8YEib0ZiGzEB65J1pgJ
HmhMfUnNwTOoUBoqlQERkOimMlZb6ERoY/Es4xqGoTH03GozSSR+luB/0w8EC0cSMs/+/5/6qb2k
63snRNfzdPA0kAm/0KGIKCs/cB4b//F+OFVgL7Rc3cJ4Zpd91ngOsV6wXsBVB2HhTXRZVkVCi+PW
dcFlS1ugBdrAM6CG2AFlA98R0HXnZfzLomjY4sBiQvR8x/bgR3tnT1kYkgndy9PDiNCz3TsJRUnF
hkqUIhQGvR7aSJj0ut6v9daVODuRu61C72OHU4SNrxNdO2LWBD5RVbxLXU//nZbmJF2CUf5syzoZ
QSREBDLPKmRgaPp2c5Ag2YANCuLjf3iCdSc9eMBLiCwBps+S/z7CojvnotZLlUW6AUWOenzPBp48
SBdA7/40hH6gWgD1KRh53XpjEFgjS6XosinZNk1zpYQsRAEQUoRdeWE3P+b8vul0uZmeNRdbaYrR
o4F3ZvhTMp7VZ0BNJXfigBU6GbYhnUKUFqLeZQPhFyuW1D4Nv65LSJs4/5U2koF4yMNT7QoAerwb
ozx9ZM1UKqCVUhsvauvjsRpqvUM87D2Tw6pWIWr9mksHHsFdpXeJeikV0A6gFNj2UHJFRnIvjEMN
r3cISeoV/jP1yEJD8Ak1O5YQVRT3VDKN8XrsopAPSQ4VLp/sdmgKVi13VXLHJ5X5z99J1yFP2G5A
wQsaepeJEKefm0Oc/d8uEyvgGUBrETh7qUZW8Hpc13SvHICqYIKBRdU+jdAj+VkJf2ADv5ylrNT3
JDY9sG2edYUwBvHYqS56rQ+ITn7PCnqYGWAJL96TpuDQxXUmoz1oqaOUQXV1qzpBNiivZkgBRFM2
+H6Z+crJD7CWe10v1XYf2Ypx9KNhsm3DV+I8y++bj54WuNmPdLZAle4HhVWSLiUtLAG7jipfVgjF
GH3HzeTmok3baxjEEEDQEloNnnuANWbLjJaBXNjuGeIJg0iV/VBSkCIo6MzykclGuhabI1KwMYfo
y0oQwcSjSlRrY2YbgwVVq5F/C0eMZ1w2xG3VDxT7LDXFN4aFP99azvoZk+LGYnWRG+IFm/J7iXXk
+8fmjSoO2Ub3fmKbZA0DG6bciZREC9KaVaN9XVRCtzIAikFpyAUCTWIFDHu+GCMvndjMru/p/XMx
7TrqedHQWl4lEnsRrrcJg6mQ2FkXuD4YF2RfK8ficpzcfWLSRHptmDVisMBXtiHE3bHTapsOWqS+
Yn2iMnCqSc2pY252aTFt2EwGdC7lPywtF3Tr1kJt5fClCwY4w4etDRVxl0yxLeRO5evkSE+Od7ul
yz+P6b+GLUANg258cR+AHGnFzcFxPAkKzxSor2sGYUtaeQ/CN9iMvS1FjC4bzdk9RGDNsOUflP2Y
3Nb4LxvtCjTOoScnriAFfgrlnDjPYLUUx9R6mjw0gKwIJfJvFdXN/H3uG2eZ2OxljCYhR1yhC1Rq
58OjMYdQucwRNFegDr69T/C/XyCG24wrQo5U+rpybNtbdcVIQMnSweLhwKMsOBhJxvE92dxfie5Y
VJsohIg9k4lr0VYQgt/d/HbTNzgOE0xcwKy3QKiBaTvceY4ezdvuF3u3KBnuGZs7JlvnPldLCQ6I
xMp5SFYk34uMfyTxXBAOdab8pkRANuaRQWrg8UT46TEQrtkozvrbBt2LVCpsoy3M7FQxnCvtAiI8
AzdHlz0C09IvWA6oO4eEz/G0W2/UYsniE48XSAlHHLBx74jY6161mehZGwWdFfXV+XljV6Iwwq9V
+XiRY+PLmq+1iNog7QrpcEA4N1zw6XJ47ssg2yzrJWzkbr1dTYyUB7obKymfShKi7/dkAVKzeqjh
+P5aFSO7eQrxzkJ/Mob2Hj+0L3E0tlMnCP53Mpc1VMH+5uibB4ME1cJSIb1zA99XNrBHDY21m8M6
3dMFbIDbgtez75VRfRFQ+GQLKCLoIAI7rC4zoQP6ik3tv56+haSqAhLToOZZwxT5qd4UlQRJwuEZ
9k+C6aRw7egnZ2EGdRB5z22Mts+GGrI6/654INqURzslF4C0v9Zyzw82WjICDaaojptZnOkv/Ec9
xEc7vjnhAtB4u4RvHgRen8BuBXCzwgGvAok+op5ZgOPYaOIw+kTmX4kMf21DfQURKvRbpGevCpzv
od9LPtkgCVayqVsgESA3o/j31s6f8rX/+xKWfrKqyb3XvYguddz2/a8dIvAcSyuoXmCG2YXqTg47
zxLsJ83FeZWLYmK6tGFDLrKD+FPkbNElzqP5M9SHWEE/dQGl4VnLTS/8no6Bk8fIUaMRf6EFOmCS
OKDW7r5kW9CXBqBMGbf1YtV/I/Qhd8d+sIjmS6YMjo+CJ5TucmvD6B/NPN4b3XQBTdR7pzjPXP0i
1osaAxQkasJl95y/d/rZst/tNsp0XdkFKI2BXrBT1mhRfoJ6RJJFvnmWIfkodt1FXIFQcPx4sZg3
ZgKhsMG6hGo/IScEF09gdoeMPNJTXuKHa3CyTXtryQVObXoXDOVRwK9X+iJ1UEgTMtidlQYtL8fo
ubqilOOvhtb2u2aX1yUVtSQUyWXnaopGzwMoZ7HZ6r3hYHURcsyOlFLi7i2jXJ/UPKPzuLJasN2g
Y/p+u5urE+wzBuv40EnCtAAaSaQdgyd3oJW1rigX3Kqh88KdY44L3zDFVQqQoTZd5VXuD1op53Ly
ujpRxkhkgrUMsufk4G7pqCmsBsJUs9wKdtRASRfN2OvVceoOO9KlMUEh75wl3NpHYD6H0PMd6x8/
wfGWC/NbXe/pZoRAOnpxndwSaZ5pjrsyiBkk1PxApahZOtndQKErHjXXvLt1cf4ANxhsAPZqcBqW
+XQiSPt+c5561RHBdgmU+69Tf/idgXKFHGn4UdwRl16QIFHc36Y7mYhFoTQQTAWOrapuA0mKS4hv
K/YchGZ2MymY1dVaH4ObM3n8yUfdY5SYq/TatLu3ykOBuydCXXIk2pEwixu+n7lUuxpRJVPVOwA7
VZAJt45C0zEDb5oG/Cqes444E+TFuVi/5a9F2if+HQrXph6tm+7BxW+4MyqfuXHC/zdg8x4OYiKd
4gRRZ4bwhCYMJjExsYP1kN0JfToDIkPAwlW5fQRqagQHdghK5o3ucDzrjxixtkzcEqzVM/DnpLsf
NXik5nBy5I6CiVsPVa1tePOunuA8SiYPZlS7Csei2ui8yvmc7zTfwxCnImKwHjYmxujl5dItRQA1
gvcL+kYTvpr9vHnyDBkfMUdzVab1IkmT5TvyC8hYLVA5K0L9ePgMbBd+A2Tj/xyBotTskdC09d6H
B2VvFPZvy0rNkxtaFLqesqvpb8OM3Db4bsprzIBdayTTLfaYvhhGngIQHxOzG/DN16iTJrDhtkdS
uDSMjzg4GNbzaXHxHNzUgDOKfBeVRemL/trY6yWGXqr5uqbkWqNIs/oVd/Gytp0VjPdgWuBLuL8s
bWxDjIGI6GwS898/MfdRlu50nYV4vOKXuHzsE6wGmdGuNPKOg/6ctaU6Uf0zrfmjnT+RU+hYZFKr
8ecmEDj6vWgLH0WVdH5PbItv/xKjom7Yx/09s3tUAW6Y/xMSEGDN15wY/4QXdsGEFZlaEfmZjyxQ
3Yp1hh7VJGiYZ1Vvk3VpCJPpfWGfysiOUEW2n4gpQ+7kPy2yB9ZQZCOCdC7ND/ws2wKE4wLna1Wl
kS45oOiUyzat/5SRkll+QGJW9z4Io+QxuQ7VWp6SmnjIlw72p59PzgLGzEVaIOQyfVf+AQbY3V+H
L1puiBOLNh2RxyERiuxL7FFYFyAV+lpKMJq/6GNEiPrMfoIq6Rp7xToGwC9T6XyK2fAnUv2F8PT+
8QLz2IkGpAR+jv3vzRYxy8WVVu7TpEjyNZ45VXE12bM3c5DCMW/Z1DRz+z5Z4cCy3KKJGjN1mMGU
bLms/jcA1dnioRvi00JdH+OIIaYifNJICulYisca5lY5ayXuRXh2j3edydHiLSwUECYO46dtAY16
RHIJK5V7lG+B95dpU+/lJ4GZMo4g1duD2ZEJai7kXOXLWWmWYrjWC7zOlnjORFg23BuhBooFq/85
v3850xz36HbHpN3YiyQ9E9Eru0tM7PlxytaSrpAzuMR3T1sypjjICSVDBjQp0kLpsDRFQfr+fv0k
9yA11AkeaP6Hu5nmz1XfqX2jIv2CAkyrodKqDFfHU+wN+nR0AW7txnSdfHD4z5CFm9zo3SEUrUqd
m8uOR70zk5F3vQUy15zJq1yJJan/0I2CVrKVGGl1pHWCmuoszl+QxDzQJ9xQC933Ir2CFQZDyS74
mUkEd8Eigkv9BQaBKpabm0wFdYiRCin7E0PYKL2+BghEpss+I1ZbWPALE1XXcNHiKu5DyibiWZKA
NN4ZioSdIbRdQVKGfGdzfcVZ+V1mpU3x3RR9O03e5yQ0ciPJzVISR9NHIaMheZvLHaHmd4LVEn4w
VnrXz1c/P2E1huB3D3k+eVxq0RvRSiWrNU7QlnuCgRDvyUEc5oat9Z2cOln/q4cBga+zhlU6XQdD
6m+DZ4mMgUvwBuKMEvHdseaXczcqsrw85IUBKkcC4OopsapW95JfjiBViPbpJlNKlC8+7AljnART
/zHfsdurpeaZLK4ZudAwJEbytqfpr8gmv3e105iMKFMgwHF8bTAmEp27MrUHKtNvq9fwK2ALdan6
AgTEPJxvTmQijKmdUMLnckfifTQ/Ui3DngbG4VS36+T6VfDDKcn4jP4Gv57BHezYSxGpwHBCnULC
2f0PL6PfNVjW1qrbydO0kwSoF7De66iLv48D/i1vTNtaXUQ8FWKfHyaGfyD2BtWNiOGuFWx3licX
qyJLbNd88YFNuTMNqtEEfAGdgHf6lmLzr8W4/prXuGcNFvqlgocZoFounoieH2WffC/s605gJ8jY
s7llYPCBv/hCGdsPaKrwG0xu7uA4AJt2YWbXXfkTlqOPjItO0HBzONTSzMTrkS/y3T4l0yI0Gcci
vkw8MJW2HGq112+Wu10ZIWZ4M06joncDgtfXuAMDsixcLw+Rfq6YGFnGMJdHb335IE/cSZBC8FBG
pmLvfGnchS0NEPDsxPJsvdwCNxVk1128f9WNv0pbnFaEYG3rUA1orEQXXYLD1kkPfPCaIeZ6SiQ3
g/XDul7TxCnP6+7hAmvVZo20FZuAx9oRG7cR4/GV081EaIFc3tCAXZu8Vx4sb4ohMafbFRL5BBmk
BrqpLTGteRLpJIUeOjrJq2dswPhFg0d5u//905aKpIIQ27MQWrUDbMJEEA0mtmUJyIeNFN4eTksP
ckItooAM0Fs+8+w2sVN/LPdikPf12bUEfTWGkogyHLuGYKsrz1xuBs1SpAq9YEWMEGLjai6VPIgL
3BceoMpWqcy0KgIVnQwlEop/y7QpZRPLZ8OsZJ7UdMSWtBHUgLDfJf3qMWXAvqMlX1zhNq//oQD6
X6MFCc7gERNbJTKCxtXVflzguGSrLtEuuADktzC5gq/HwNvJ4aRKztaZkP7qRrp+AowyE1Bh8uYB
ownBxPGw/8mGCzpUYTYGIViG/0t0diCtxF9yZkcK+F5otoHyIY99jjLFXU+7IlUkHlet6jP3KGmR
JfvKlDTHSt/XTSBtbFgkjPX6Yuk8ku3zDsObusE+iGAVk3mnAOpoH0lJhAAueGcNBWaI7SZOO328
TJzjnZGvtZ1kxe6ugsKv6XNYuLj9V3bsv1FYYBzSr1yESM7dRWsFQXzZFeXT5wrD4loAHUwCHkaB
9DNAHu/wVCQPaaL57b49iu2A30igNIfzFnoI79G8/E6NARmv7gi8nFrdeB9KTe9tU/ZcYOup1vhg
huoNIklNYojkTRaa/WqVfiNfDYL4OQvVqBiAooOCRTXrWu7Akc3Gvjnrlp6zvx7mNm4z0GJYXh+b
01o2RdcXduxJRhlx641/xr6Ehgj8LYkhHqFPkdezZyZYBRBFf0Pavx7lHfclCgTjpvyvAfZ1XWu4
JI10m5JoObnh2VVJAxeOhLsztkTMQXgz/DhuTsqICFdYDSm1WcLAhD+3RO/Y+CSIR/jaRnVEx/Ju
o0nBFT/9PdA/Ds9V0QLemxhwF4xb7qW83uatqTk5mDpBBtghOHU/fmqWclFgrJY7tWkXIG3HLudR
FtnMhJaJAAJa6JS7Oh8onY3CYV3mCfBaClkIyhuSKu3Tr8SXjSreHB3jVdVLh6mopGxc3wxLsosy
ky704VKzqwugQ1mjgI94Mm+16Xv+SCRL9MuP9zB0e33pijbYkeZSKLcafK+DTvpVIUU7/Q3uOyBe
5TG+iWA/eL0QW8WKeAgg1WRztNwu4vcpVyrbUb3KW+Pu+x/1oJ8Zqy5nrI97LtD3CwpQBxawCpZ6
YOkqHdXp9Aeypggv8SOC++DzYtjGjjBg795VHKMpHNK4IIccIuVS4S7OhOgcQd2w6PXcnoDvWY2X
I3SfiBXsIVq5YZxRSDyqIMiKlzfjDyZONTnHmbyYMnK6eTc9vumh4Irgj8qnB75QqnGt6LWPjRTk
sQZQwLqhj0dbR+5gDPE+5gDoxN3RhoU7yhYOu9FRIXY289PEsJ+Bd9A6zf31Q1EPLFIe80rOI03R
M7AySjDOTVOldEjQ/1cQR82m7yz5/iLkisEwK9Qj24T5qMQZqQHfmMpPgFkjQomxYA+r5GiUJdF4
21QxwwX28VVBlJWFIatVrwJeEwHhvBkZVaQMLo6ccUfmutRG/iqaFxKaiaAqKjq8tXyq6Y0+ny5O
2wRXjN/0oQGsj9F/77yebHR3yyK5U/VspGYq59AWJZl42TgNdB+1ph4if04sRbroGA0zNNl81ioj
unIzQFPa+FsGWYt1ASOWUmtJflNlQyAucVK6kM+GSme/6x4BgYk4CoDzCz3OApnLT4lMzK6Tb+xL
KG9rW2R/e76RB9dS95WfETq8DXUMmfAej1w5rhcVYoP5FCAPj7+sbiC1NC9hb1DRXCcbqO91UBIh
27e6NvF5lTHvzIMeH42HnjgtSDLt7mNBxhL4si+24twgYiGb+jZaYaH+VXnn0YIIXql0PBbKOJyN
1fujui7t7exg4fdMAzL3kkOyzIzwTELMNa8toyaJODVn8Rck7ujF3k72va5X83EI4j01aSylGGbO
ux4RIYsh3OP/Oy28frVeqc23BIJhfwpZE9SX1LUxQXfK7tavCPwjxxLWtBMmhqvzFI60lc3MI6Z+
Ebq2mUzgxsB1+bg69rfXpCPAEwoRefry6ZyFVXttUFXNPqJgaPre6U45A0w/wLpyt6SRi0itEaBL
G5fOtWKURdBaSgocq3OO5UB3cHGDNCNtNZ3iWaERebNu61ljTxCu1jcO/tUum+ZndPHbMRmsrwRs
yGI21O0hk/vJrvir1TfDGMqY1ZGk+Twi+0YrpFMvpf1kicGdOfxpk/QMm/tJkTajSu34xwJkIhsc
7zf9dLKVBzPg/6Niik0REjd6lXLxWFcZfu7xJN6I5Ohz0j+DhlRrQIkZV1VVu0QdTLB28q1/cKvK
9WWCaWQJDcVPt7BgUpDgYBy1Jo8LXU5sA0GTD44NpVlErdL+lF5iwee7M3SJxq2/DgEovMPnt1Os
xUgDJ/mMQNdIHn92t3c7RruFKTw13tAp9sm39VTOGo55547CmGoYXL58iH/YDx54UD6upAo5UwvZ
e7FZ15UM0T9SUEdn7u69JJj6jrdCJXPhYj2nAcFoshDOE998Y42AMmU/ElfUSL0jktFxqkQNUWG6
BTnO9ZOGTauql+Iu0UvtLJmbsG3QgZrJjnnq3efKU7Xv0zm2K41LHi3fRIXAz/0vDtyvX3PNYajf
UiSFVFVIBmYR3K3Hxu+Rz5WyOrxLqR6IRL/+m2wUu++X0TIV2fJcyqFHRrua+s0FeOOL9b7ckYuh
6yZpngJuyHWzF/vIeYA57zswGj6uB/9oYlwDta4jYplJPV2nEiS4ompYKqFibkxypKcgMlR7NzxX
6ETYok3FWKYJMjYFQiD4jArxolvCXi9h/NyYQDdjreevoXL43pkCmrDFzkXXood7j5PgQxxGhfMJ
h3JqmXlXMXqFWDnJoA7SpqDRhGoeeLedYLczM2QttTaY/FS1FFLSACicrqKYZHfljum99opI5il8
xheYMilwSkSGSS0J+mj4ln2ALYA6uEnHOe3GBq95NUIJ2xZut0HRhQIp/yZfoQM+wDJxRdM6ge2X
XSGtimw/d+/1wtqo5Gvy9xuvLvEyyVsftw+f7TOAkwHs5m4ErafJnhKCgtmqdIn4UgAWPl1EW72Y
lGiL4Quw6g4RvNbQBEuwWUFYk1xmLdOdyhUSXVmLsSRJFulpTa1IMuian16F6acNTfr0PUlmeyOA
OoPngDvIjTPQYZCiyo8hP8pvh+fTwfBnHWfynnBWLyKmcOgq62Y8ed9dI+MPJv3RHq7jDRGhgfae
KFnOwhrtdIiqbh6g+yJBn6/aLqYax4xR4dBtW95TKNp5RVxl5Tpyp+TZEYtAXyEe9V51XrqaLfO7
orNpTsrfPJDxyBwDyqmQ9GYWsM5WiZ3r2JJJ7JJt/2FIyNoI6jHR5KqJVZ1zDPzPyCfTou8Iof5S
tDRMS1v63W7Q0KRWXC8gwzdJKbrHIApMbglI0rxakhcCVEOvXiicg6YHUG+12ypXpXiNR5ApYkVV
JggaE5/b2ZPGv7aPlB2yBIMFXH6FYOkbX/H+PQglZXLjfB0JgR3FQnsG5Jye5oadJ2r6cRZPzifv
z+e21MQzL3MQ4/X0Qolco5JhjHVLA7zQ+5zn3JXDR5jyQhb5QuQB7JdwSS9iaRiTLk/CU0PTdKa3
T4Fpk4OKV2BSE2tg1irT3F8pcxdBY0dF2Ab6/oHmqm/hOQjwMkdtr3aMkvxR9JN00cunLT0qsUS0
y+E4iTSNZKfW8fbSCxuHpB4Hy5JcSd9u76amgqmVFUdeFZs30WdtLYTF77ecKkJGpdHYU9SGcQRF
fN0H1b+/Nd4C2RIL1GyY62gKYmhyoeQoVMqWEhCmPwgsssVJQ+6Y7/azyecoK2AKeLk0p58HeVSA
FMxLQHPWk11X1ogarS2+CWtXcvDNlNTc2XZxi3D+BC13NSt4s2odCQAcbmb1zSK8ctUeDMzjjQFb
Rj31rYxK76ZdtAct5XBPTQaWIsNw+BFFui3687xZeNV8XsZ7/dgfJXCFSQhy7jDhm6+dUILRAb+A
ifQEf8GQVV8pp41TU6tudbxfBNweaey8BseVUpaJIYh4w7JxRG3EgdXu8nmefiBaL15MWidrEVJp
jFNvqMVZSH4c7SUCUuGWsGR4Pfj1lxUcJ6P0J42ahJ1rW1Mg0JD2YCyzVveSjlDSyr5n++jnSN2/
yGoSLahKoChxbBW8Urra+S+hRqr6PjgeFPu7OD7+YEH/8Fz8wdivqdWyw4lA/WLa6r7ju01VbDe/
mlI+2Od5VbodYt3J2giBZa/Y8w2D9HbLu5HHVSljj+5jTYuzF1e8UiSY3CZeZfJWEO8ega0jEz9L
xMPIUgL36rUWyckEuWxxXtfcc7RtsL/g+8v0YOkLerCjxAEKLNKO+Y5nMvJB/Pllz4r3c7xviYlj
Njfh8WKwpyKCooCq4LQLeLciTkrl/dittsrYbX9BKWXyb/ru6hO7GqGOEmSA8dpCLrhs6/JD4sHj
+F2tb0fjuambaut5npV0RdVSW+nEMz8sIPaQsGqUg3VDcUQkIajDmGNeCJMrjlKp59Cqjp5rLqpQ
SjKnna+rnZdEul+k+QvFfw4gmOo+IeeUiXM010jtNeeBGoqoXoLyyyhnqK3Zw6whAdGXPZiitoSx
oRG2SVe3rYJHwx+CgEUNWSvjvevUbDzUOdNLSghWUKDC2uITtYuIb6yaF8cd8e1HYp1gymU8yeHz
X4rOYm4ih0R9BNETVCgYlh8R8oKwv6tb9ZJRvvnYnJc0o6YKJY6295Yu4yPvzHGxp7oJHT4rC7ZU
bvJBV+b9xrv/5Upmq1B4TT5nmAkgqJup+AuDLUedz4onZJY2Uy3j1OV0IU13IZHQapvw4LXtow6q
hNXPgnFTCualZ3Mq6pgT46HXjqApBDNk0cajpWY4FevK8ljAdclJcVGHgkzbc5IZvBwO+pHG8W2h
DQufvDngfqWr6c9IGix6GkRFTzrOaU4REPVTuBGKz4TXeaXD7lc5mmubyj2vhzaNNJu5wjAgdD7M
U4jIDpAloO2fUhpTdfwAnrByBee5Rj+fizIpZQLhkjN7IwTMaSzE0oQsTj/Rpkieppsbuf4O+gXK
nP7YL6pPePwk7BHckxfHwpF3dpQvTSezvtTEmD7yfuCSUJ/P/tm8BkRWk2KXgAjzcFaVdEjYfuyW
pzfVndGHtt2dbA/NQmvsOnHf0Rm5Hoz65Daaj4aD0wjeW27kBtgy0AhwcVsk2ZbXBXB+ay5o7/If
4GdRjWOoVrJ4sVROgKCYhvDKUfmecUFWYqNoGqXkcf/WyjsPlHC/6oqIMhj1jes6Cm6/CWnJhgKr
v/xACwz1uckaEw85tsF2FgHEOCK+1ZJB6kYYnyXQK9X7Gs/83jlSkZ2PEjda3AleaZ68ISYDTYly
PwiPcqoZXJnQbXKunDHeGesJwpqhpM2FIbTZHvkjff2dQiuthiXFSen0GDThp4yDGyV4ZgFUoxPW
7bn4afZHqAECwLfRgMEHdBmjP4LHhNOj2Da29e2rW83jrmGLFpTutRbIDfSQtcVl6V3VX3HbklOk
OWZJyMRUgVgmnXIKcQiNBcyGMxCpvZFxhifJzZwnXGzp61L5s1iF/PwBw2yPPphj5uE0EjJ5PAQo
Fzc/t03r7unwHtw/hCTNfXqq4dm/8DRNC867PyZd1yAIL/2+vXekutLq0nZ6Q567YJQ3zcMia3rC
62AX9uLAGIHnR0aNIP426htQiNn5UCvUFOSrENrf918FNVfxyUIkQFqmM6CwV+TLyJHO/JaL4+64
e/AEiQc5H/PreY5t79GHpsokgCoECu5+VQSNz09ng3Jh6w9OM4Kr3Isxf/BXSmk7eyxGKu5jvjsK
BY4wI4mkCI/aWOrtrMAAm1akcgNOm5AR9AbOZ4pK6HDxHayKUJqgC7a6Z9J3UGqiGF8PeO9N/Bmb
rxUeSmff4xcPSeirX3gd6I/PyvgqlfTmMd2y++h5iqSCNyesvq07kEZdAcZQgCodSuGQRHhege3J
GTy+ix+sTmY0utIHALS9PTfJ3Peqm4v196BkkFGAqoFAq+4vWJUJ0f1ylG0Gr4A7aKkpSdde9D/T
kPPRr+mQBleRT/P/OZBE+Ddu1+oVqKNBzGv1HXmjjhn8tE5hK0B2VvN+Fat/snsdYuDZ2TF3mOiB
zsN4JngkySyyIZyJNSHDP2Gu4RXV2CMjX+68WGtqjTBHXnQcC0qpur7XJl3qghNn5XYseDGa/3c6
wTpier3LP4pEd9xCZ1yAVasasxYpru5da2zarNlz8vXtEUxQ0zoqZVddEvH1ASS+xZYzZ35+OUHI
5xJ19QnpZqF3rOXKC8BZXAjAabhHexJpDsLrxVGKuctI4jlZYrhs0ZATjMP9JdSXdHxJptoN0zGn
SZv0TRIt8wZWQUp/xLJk0dgBLxPX/iakd8gOIy6nl/WgN7q3ZoQk2QW641jRam5ec6u+jaThctFv
0bFsQpoou3aeYi7b/KYNe3gjfBSCifnXKj5OKQgZdJIb5efdPgoaXBHuwDGQ2BCHdNcsDSZBuYBL
ahYGQecLREebH67/eOUhI519jalknASbFlke2vyKIzfiW86TAGQQ4OlL0XNe5KDmJNVK6LKde44b
KLLXCDql/ALu+HhymnCeFOzr7wjWMc4H/z27XZfhSMPbrGPz6zJshcg3Hksb2F814iKkemCix7jA
rWTe2qdR55ieFKu8yVOcnW+8SM8JGa2r2wZTVL4GdYMPejwgAjDKkIW93+/VpdCrfdkMaOu8GBZ1
OCdkVoUq1iClGmcK5RLSqPNE8FCTTZsW0fHoQw8FRE5R9PcjXN7KV/Nm+S+Y92QQckiZ3Kej43Em
0srlL+xruNc8vtrckPwc/UCUJiuYmE00cTa1EEa4evGUe6VItAVNK2QJ/UKZpH6XL3g0SyYccpRO
EW9zw2Cf14i+JDBaIuPX7QB4NTjQJT583HQCCe6etBtdgWKsrt2LEHnRK1G1/PfqP7CtEJvit6nT
rGCAWJHdApMtyTnd2jY/6zmVp7JuaZxuC9oDC4YeSzy4MFyDyoqPH1q0VCxNRi1d+KU0JxiX6T2a
XyM5GyuPrq7fHHonhyerqkGNmGcG/ADdR1h4+P8YCaBM6XfWC8QQ/FHruF09NIqp9EL0VmzcCvQk
FJ7fuAFWWbEzUF3NKGefLycQWOzRf5yQn2Fq+atVFR9Z6iqOwV85MidLeWSc46vDVSjWoc8Sio65
fRLxlEIHNkcIP9IZhO1VTvqbOxXNNY54z/8oIEJPAv+Tt1eOR4x5j/yD7kzsArRp0LY121/lH/Kz
NLVURuob6PxzrcTDnzNIly+199kdEcESPiepZ0nURcrKK0yQDUWvISh7mRBUeP2xlPtJPoFCqpZ6
NeUacwASmp7Whr/w+zSHCpgP56GwIvyZ0HMmf8PRGaLq5i0s0ParmByWyl2GzfEh2F2s0p7ZTd3T
CjB+6Wfc5cC+AMRWmig4nTOUJCJyGkrrwBXTsrJwjooEhXEbn70VceLfYGjMgeST4iMqavSysmgg
DR98xKGqlE3v2IVJxkXHrkY0yaC9k/23X5DJIE8YISRm/V12Zh2QaOn+EuqSczUtOK+ik8IMaAAr
t453Z/I9E3ClcmTw9PtYnc3szv+A2pWaJoaPrsAnbgRFEZ78qVC1ACcC0CeKgoYcHdI0XdFg6L6o
Er5+ai1d3myfUNLlufcdZzpf5CaZC3j/e9jK8eq3qBExBNg1vkOVjjGSp8knSI9TQgu5VNNeVJQr
VEpb9qq3igvLzIhellw1IBsTqjbcqn7ziEylStKSILR8ijppm4D2w439UqzfBpbhRT4GlNqiEhDF
2qxflFHDd+Q/XRnzV9BtEhXGWa136nenwzQHvW+7+0p5kwHJrom3E+XXgOW3KlLc+2No0yPgxbaz
185P5p57SCbg/Z90gNBhsPNJcyPV24C48f3wXt6RVA/USfWln7cONWnuzKVkv1CqsYhEUJ0tBDVC
NyLIXgWJRh18NRwReCpdWYUncw/Bf59adEym3QNMcI5E4VKId+nvGKXIZjxBLf71txHgaC1IRFhr
AG7nk5HoUMFja3nLdxYaInIzrQDNzqEl/gGpRtpFZ9wBdumxlIlcHFWvKB572Vj7MQfAftdIxTOJ
ag5+XeYZwVt7nDtX9zlOMQJGiFZLsP3caoj/Q5n2yj05cjzmIm66Zvg04yQiz7KdeSxfw7VjwV5A
KkQPetWzV6OpTQ7jCnO0ncOTbUOFs/vt89g0KywGY0DxqkoUbLNol2LXmjTkzrEQixkFOMrZanQI
Ca5vwy6wyNJ/PuyG3eWpVuJw0z896pOKooQJZnRvA8/O8VXPLCJLmcD/78UVbfV99ikKtPIJFEDz
ALMPP1T1/eTLCJWg/fpHaFGe6EXery4gaZsMtyxIBZ9oMXYAAWZ21bTMeFPeRnZ4XZC/Pe7MGVZh
3o9qO6QN4URFdPLybOXpGH8hxvUOjExkPY1gMl8Z+KyCN/dalDitnezXrQmIBYKZxcfoHnvHE56G
iG/Il1IpamB9wDVPYdMUcs6MqwD3I8Jyg8rjqZZtA89VYk2RLsLiqIYDT4AT1OPEzYB5I1RDI4wH
ksVXFOyjQK36DQBiA9QeI2xCwYWxuaDH224/LkXqD/+IkRSuEvjAXOvsNhJekPIWwD2f/7E9hTPr
rkHYYowve90yzeKUmjC7A7cSSxRmId06Do6cPHjaLOKlp0QSjoBCtQ8fJZENwruPyVTalLp3GFS1
sTv4HClkFFGGvPEIsFC7zuzNpnqZo19tY4Fj1gxV1XkcOvbBbYXZtesPt4VYY2XVP+vLxIPRzpwv
QwbH2HWICvgX0PUxYo9yl9YZeKJCHwX/kZxRegzt4TEJZddko/dKRk4s2VBUefqMOrrl8LzF1yLI
AeZL/TpBuhX+0L/vETgl+DxhhWT+JuBJZWXurzsdZmo1bEijRZ9mjZCDAU252Y3bjNXiw8Jj1vxz
iEjas/sby1aqQ0bp2E7n80Tp+0BoVwLYHXMiqyJPskG7JsOLdk9KBSnCcQY0n0yV9wB+YI801axk
JSewX8pUHl1VZoJolpvGbDZywQTp5Xcn0pThOrA23gD5zC8e5tjQ+UIGPye2hHcZieXH9JG/1mV1
CAnwPOsga3Do+MuR2/PEYHh0TOR01oD/HC4NBYFcHgNL82P7IumdQ6oKma/FRvaUdSo2REIcsuos
MB1Ql3iPZ1Cg+QL1D2KfdTWwWAKanSdLl9VMrPHjZtvU3RdgQ439DR712u1mw01WZcxFzt9GXgvO
5Krkval0ci2JfjoOFp9x87Czru8Xi3IxONtO8y98ibyE+6FFO9nI7jcmV0loU6oMpcBiYSZ2Qt2+
zXee6Aaz2FPyyewCxJ48+T6mzKCjrDqcS5xxd7MMHlHbwhBengHsjDg+GoGoAtj2bR9toyu5gyep
pK2eUrCK6rnez52pq1O0IkSHQVkX92OyUfycgrJupDsoAZWKqz3BYwK7PIwpTAC6U3pgwJyFrljl
aAJYwqXm/67jwgPZIqflKcFaxU1i9hwViY35eWRTm8Zn8kXuEqduQ7/efx5/KaIbIy7l/QTHxeUf
9iGV38i5ZvddKGfLEvJw+L4cDYxuH+1sB6KYxhYNscvM6vuao6f9ugPVv4cgiXAU8jOzbshV3jtb
PPPn9R6yTKj/yDdo4rcwJySk2yQb5I6Iv7fkdu3Bg1s7pxnFs1LTxJKPO/OKDH3QiWDz9yp+1yOQ
gmFkF2lmblvS3eoHttkmxe6prQbsBMx3BIfSux1xnMwbCTGS3s60oRzTwqUe0FzMVIZIBJfpWh41
3A2/ze+UZzZB7rO3+VAI/C+r4udvbx+6Pu7eRHh+Z99z69Nq/0fa/eS3nnkiTQHU7q79UGcAiey4
bUEu0reDp+fyyVE2u3mRYCfG7VD/8lzyNM4HsU0k7+9bcrIiM+wfGcYyEP3zW2ZiT8CPiYd/wgbb
UGywZlpqWI2RsZ3s6jlDTEn7yjgCsQnZRbAN7X0R4wguv5TwO9hq3CmqhTiAgtofhfmp5Be1sJLQ
Z2DxHG0CrfXNWkibv04Ki+p4I6qVx2rumc+PRFioIkv0dFQ1rh7oBhCSVce+g5yn2vANZoWyQ7vi
N8YgT9xSk13tC/ismi49DC+eRqWte8BAwrbwij/t7kSEkOL8dOfbAK4iXPhwTgPN5PXkk69WnLsC
MdeLIPcUony2TfGyxW+0+0+LLJeiYdrdtGtZB5MMhopZ95DDk1r/QM+5p1D792/iPL2X/3S0BUVZ
mMTLXMbQVnUpnO97vowyVKrF/4ZpBcPIV0DDusCfJlR3ySjk1YXTrJcb4tyrUA0ERk+HDYLwH0bK
l9zYh9EMD4ssxBUMJCCA2EMfFohqPbs3zeSogbZ55dPT1DTKRpX7iqILMyX8NqQZiHJhkY3M9sMk
1zo9A2gFYMmg1h7HlR1FjZBmRZnpCDWGv7nGxfNmCUBPrYId6ApyD5Z6gjlvSyfskqHNy8KORFcF
YyNC8RkNYtgBvesJz3DoASftQ0SFRPPy3RoN25j8iyCzyyqLSRNo0KPXroDL9X10DaH5jQej8jyC
55RM+7ZiTCCY5QPAwSYMBa935sK3D/qy1LyLzq7BWEOnU3SfcTej7kL44nRv8sZLDr2m4ek/jdZR
e8MR0gQg1L1wCUZUnQm0tsZ64eORaaHSLTAxKADAWmQsPDZGFxEn9VljX61Y/E02UP9xNQLWVXNK
06K5cAgaeWvT8iiwu/A92ElZ8YNbZWJnRPo2ztKbCcclDGJ0jNAWliISAezBxexEZI7Uvx3kETsf
Cu5rirYhRt+yqgpnn0nJ2VVhZkIUauQkNhOdL+VVbpxM607QSfTTYcsmRedBCmKYXB8xHNrSrOCp
RHfmaUxwF5IySgVCdylX3rtUkbsIGokorIER8VP/q164erRG6BS9cIDm8ZwtRUp0XkDSk0oAEPVp
8Zn3Q4o0OX+gQmgwWZUzi4AlvJcOd07mU3JsYcwA5IutewppGgMAJ/81nilPVdv1hgg+0Y+h2AAB
o1XEcf+f/cWolJrGmWKcz5sTpZoiHWToE0p1UcAefeM04A3KF4yOpEbzP0PBrv1+bSw/j9/VJt+l
gXWCTG9J9D8QMV4wsEuRD7vmdfNEd3h945bG676dgBhdXjrrqXlxIsimoFnfZyIevJ7hNeroiVXJ
v6etTQ9JU2LWwpiXako0u0J/948AwiIyEor3HsRqYGdYCYiHzwB3AOyDOKghdkFNnUM/Vp6QrIMl
ixq+gBlIr26phe2M1Ui82H91kC9Hm4b4GtCQDpSFBRgo6WvZF+dOqn+POTGrouvk/6p0yHc8CI0m
f3H3dcjZwLD0h9JnzZBFh6j7WAM2qztXkfHfvKZU57FAxAD8VL10XB3E62JjwzewSlaDdnyM7nZp
XS3WpfiYj33jXZkkPQ7JFwYT18QfrzdGdexFdoy0IYgLtrQzLGbtyIi1zcnqlBEAWq557xfBGEKT
0XVlM9qBoriANiv8tSpUKhGx/PoTET7cpeLENqCnMDflEkuFCEdrcvQ60EXdwU3QG4OAQdxJ+ozs
REy3dr/KbESgicTglLDXqMOQxqTfrJsj24yKgP8F0O7xyzAvXvdPj8oqfMUfHRuD8gM5odQj7XZm
dHWeKRxwj08J5/a2w8Ckzd/PMFCVpNK8I/PXqMcPaqWWAH7FUzmEwi2MB1atYPGQhhDTzsZmINSQ
MxMvuh+AyhSurz0F8XxgSTbOGee7BauIMVYDt6Gesaen0nJW1FaIFLhJHQi2EU1G+PVwmmuSSmDt
VaA0kR2PpHpX+/2hBzh85vIYX+2850EF6lzB6D+gfy2Yo/2Fc1xCGGQBFBbUiDyKJ0yMVf8l8ZUv
6G/CcFFs8cCUqMDQnbVsHXkDLBSQkJpyt9P+mGfafc2O/8dl5HTGbjaKeTcz1UP9kDG+bafT6CJu
Zf8DwlWXuzpXYWlBw9pCRIa0SAKGq+xwZb4g3Ogheh7C9cUapjg5Ag8ZxKyA0EtUPpuLo8P5lI0o
VbdW2QA4yP51BQkQYTg4UBc0YIgKUsR5FcaJ6FPDAXL+4c6547OyfFAwRzH9FSqUogJOvH8tOM4O
hoNchkBkVLcwC3ul4CBbLIwOh7ODUQDVhwI+Ssf3VbnSIXtG36/bbZ2ntUeaqDs+l4TMGjPP4Zgu
ZJIibp1qAHJ/EVyEn/ydig74yq5ZCnESdQWaiJ1wod/Bw0zqdt8ZI/KQRfongIUKQH3LNv4P4Pnp
VAaGrLCj/NeIesBP2Z2UUnlw714wUi1CzWQ3/xQiZj806GdYSirV3UWQyB2hTrXiX8ShE1unnFiU
lC6VSbf2EuumaxRfrSeqgyWNyC231zjUgqcpCsWRSo059vw6Tw4tfPYNn2dxqZ+92/lynohWmACm
zPtbKWE1oxN6CBV9QAq8bFAtRt+L6bzO7lYZIicINjWNlPEQdTDLimy0YoyneiReSIOldFE+gpW4
J4RPSDrbM7zmbEK7LINuXCURl9JZjkH03lpFAqBbFUDN2PyKUC+WDqde3x2XPUMohjJgaZ7oFbsg
csjZ17IA3Sod9P/Z8Fjo2x0SbJHelj0sm2WQ2echVHk0Z47X2PaqWWwBzFGjWxRAWcsuKU6Y85yV
lGmDu7koOhjJZPHfU7JlWT2RHYTYVvjxXQ4j/+dEXKYCxYLh9eY4QM/znnZfAY0OInE2prqUgmUq
7KYSDDd3vYffZkcSZ8fgfEV+mbNsbYipnO2MIeHTlc6GjGwk22E7BTLf24tB2yN3yINFEiWBx3wN
fIg+iQN4zbyBbq2eXVkHEf1DY0qjVGq5fSzgwpa54a/bqyVblk9W9x3PnUYWErkpYAOOMX0uJGys
4WdUWyLmJ9iZKf/4b32MM1GCoCfRdzh5sXjxTuClzSAUz/GE2oHRza+PYsSZUxfOl0QocLDlqq4f
D2YwMA7t+ZcdLWSpxAq/8YXr8k+Fzd5R6dGT2dGR+XCTdxGb+i8+K3dQHAY2RzfoMkv2ZTZQs556
CmP0r3MgLjPOMhkNq7Gim3ZD1h1O8pPF32+3X5Pz0S45YJ5lhWLd0L4zbO5ZUFEzMiNq5yJxyHAO
OiYQzT8xul/VIYe6LoXt56Re1ck1fqz7PUJGAzWM5qMcvPpWzRuEbwgNd5RFNCXrwe/GnnTGkp/S
iwOfMchw8UrUu/AhS2jlBGOXeONAVAESX4Ku8mNcEDw32j4CrTw0kBlHwIJR57SIfWci4KRaJAR5
DOF2SYAVAHqwRAN78Jat1EeOGu2vKtWi3Rv8K9EcuWsNLaLdIpbJqboNQJYvmheFFiNlpmbr/7kM
NEbSNjN0C65MmOLl8xl5+AtnYBdGe1QVKA39bVBUHzjFRD1A5M5gVxHxAdANkMzKzj349Yaqj5Sn
A/MaWiiz3YfTs8lCcy2anpkTELKdHr1XnSGc7VJIrm/4xtL3yhNfmf2OvmMrgpPhTr9wNC1aaUzK
yzeRsooLHeG1vGUX5YBm/EI6/9/+m3tw5LLAqN5KfQaOR5l0lMW6OvMnyxpTAcP2jghCgm9dKuu4
HFseDM4XXMGV61sSJJHAG5th4B69QQo7DsFhadzti/QYMmH1nGUQKk+3AIaXrSI/yJ7DrqKU6r8+
bi9IKboML/bjOAIFU5CdcqmRotiH0of5ZV88p7mm9QnPmjvepgIBOzSZL5w/Lf1a4vwPvBMZXDNL
Pg9ehl6GKP4RmT6bauzFn8dND7kffbuSPxp0z/aYU+hWPcqHBbTaFm4hbE4LgOu4C32De3//+P20
vYTztEjGrdkv8mveOSRjx0ogZWmnK+Z14126pXgYEg3Io4OWt/XHtv95+N/EXi2u68R8AN4gCZ7C
u0QNnPrYUGG/8cPeWBu+y9t3pWBo+ck2DBonw/es/9sqsA3tL+p7joRFFPAXUkSSF8gbEwDFjvSn
3CiN1Uc1GyGzCBVsBYuwUzvkI29bxBg18OLrkoJW186BwNiztcaRY4cXs/V2aR5dYKTkPLbHuzmZ
dDXyYSAC6T10HL14qN4/b+K9VCyeU5xj4bSyVNNsbHmM8yB5B3Vow8eN2lL4d32SUbS7JOvCva9W
m0EzAmo8RteY1ZTk92vbTdRMjoeHG2yY2cA9B31UHg1QM/nRWFl9xOHNbVWEsTk9HQ8gTifVXB2t
h6IORYeHE4csGiQpNGax8l9TNKMyzPAThakhBYUFhWqJq6BNcp/AjXoWzbW/8PmP0bG+TQ/tRrno
3kA2YQkW2LSK2/BhbPXgQAHJ1jAlIHPKfObP6aGSqf7kwKD31TpEC+SmFHApfABYsCdN7qzbeVnj
MDypE8x8zTOTylUgVr+7DAPuhUBlQqU7uPjlrbLWVhJqof2MaZ1uMTGqx02+5JynXAR2vI80E29s
mz97YO0q1erseiv18Hq4ytrl1zwzBE6C61XfggQKOQ6DBIdwUhPvKpibOEnOVRAjXumKxDfwhmD3
0noeP48S7annSnNAcmuEX5XMjmanHTQUSBfuS6HRnB0LR+O+Ts4fHXk0ahneBLdSt3qvAko5H1Cv
nI3GbWjWPBbAWd7o24HxTe/TtMZTTj5Um5qoBsHBFD9vU0zvyUSahua4af+/aLwBu1bhGFvpDbh+
mgs6ma9B/d6Lq9C2H99+3SO+uaqYgY0vPKRt5vLF3wwG0qy5xXY1VkHK+CRssAwXRU8Ydx3VeVFJ
VIPQXAalPbU8po2kGXKa+teyhVDTCSiJlB7vS4c0iNP1YiS4dzLOvvG/KFpYm5gi25Say/uQNcu0
UYTMq1vpoK5+FhettULgu3s6PqgP1gaFI35fWoxQNbhzY/P2KA0IfZmvQnTO0Z0iINkT1yBpDuLn
eK3/YYomLE44F/b/Mn3P9beviSQF2FajhQw+zMrK+0PUX9GJdCl5YtukTYrd/+FhegN9dvWkWm0a
mfnNh6FPW/FmAt/GgR0g3tzwEC9e7GBfwKQEBZIffvWOop2FXcur2nOW+pnruMEM7+nLhSSwwKwI
6x9E9giHu2Z2NO6Bg+5jne5edKHHZzR0D/egDf6Og/BIPQq228pdDGwiZTp3+aX4rb09T8B7Cpul
TJiFc6KZ7KBdAlzzvX6b7wlbBpvu1e4Lp8t1zcrpIbch5AK6n5G6M+cUkbfJQrT/tlnpw5x+H43M
tFYQ1dEhZ/z5Y2t2pxC09gK+yQotVdHfwQCqzHdPqw6URVQ21PCc6wdn0eJuqlLoY+NXdngo0Mif
ULWsn4WvqMZyzd7/lKWgqiM8mEYuZBkDeFLquRwL6EJVmOvVPDJEzeBT77KKKJNEJ4Bmv9yPiR8m
KSIJzEgYX6PLj2r4LmEP4Z7aDv5C6TmvhkkspsRKj6go/sqr23xXu02EyL42EUlHxRnByHQGKL2n
gZEX/z2zLJN5J08SEP1V1U5bPihgPHzfHiiV54lnmjNePdV4XuhF0Kl25CWvxPRQXQXoLVD0Zi8R
xF4HKdmLoP2H5lukMYko5K0HsNqek0J/7IrQ6R0X+F2tG119o2f2WeLXeUgu0NDIhQ+souX5xYZJ
T32GzUUSs8mOJXjC1P3y6tOgLy8b6Xp658tKrGZjMoYWVyfWwvhFujoFVuN//8PdxQnuNugC2QP0
neGKeKYpyW/D5ufbuQNjLnDneEgCg2ycMFW+cXevHeetMSI/gctv+SLtxrWvMLo2p92Fe5h69rf/
u4RrPMko92pU49iRpV87UBUu3dbnYZ89dfWR5Gj/81n35hishxFDShKpUogVYdbqPgyM2ROa4dxD
Vzvd1atOTSYP02AAt+0AToMmDCNGeWB0XNPawa5u9s2LJaOcz6HyILxHw49toq9Xx3ldjkRiXPNJ
45z3WxloDaVMmss+bOEu7dehq7R3VdD6n8UD/HN30CbqBNnvwLzmuxEz4OxATPGkWSl9niee5KpR
bAbFMG05kAgYQLPMF051OWdvFcG/Qs7Fzwh5RsGUewC1+p6mKSnTnfAPAk5Nhx1bjMbipcmQcF9T
BzSNNfemlX1dPLYlQN9RJda3t7CgGiGSJbuSOXTZusDWbBDC1G5kpSNFv6k13TY5RaTkPLieBNBz
XLN8u9vjhTJu1p5b/MCrsxscdkwoPitsgvztn7kZm3nntajk6JNHi7Z3HKwX+k6i1OSoswynzgOb
P3y1tKSNUjAt8OLh26juxCgO96SZ6QzlTziVmejghXw5Z4V5WUeVO2lD7b3B5+ZgqSeusBR/Dql8
D9ZGXFJKsJvEGPiXIiILx8O62Frq9iSvzXRiNUDhHTqU4Jn6qaqL7EWDwmEe71TKz+rqE1vQVcav
keysiiewmf+3AS/8QO5Zkr6XYAr/WsZ2Z8Pjlqr//N7FXn/LQ9Jm81aLfnS6MMbB7AuNIHrnpCPm
F/leVk3AfC3Xv+Asni9F43rQYrLpaAQ0eDcw+/weL8oJ/Yym5cW5MJoI8JaWRPY0v3e+4xHG4f1+
IYv4n7It+j+YRV272n/AGsu1M8Svh7Q9shoGeuyYajThxI0CLbvwm2iB1lvLWUkD0d+xaPCUNCck
28pgwQIrDIWLJMPXkesHkEWv2iHHmvzIRxQCupG32LFreyrsnIUNBh8SLBgNJPTNj0b5/NoKhwzw
9SOCf6y1UTaC6aGXPciMSPMTmOHeJz4TlVGxio2DehjV5mSIIyQ55WGEdAlKOd5Os1Q4j6kndyIP
elah50e+5JI+ZNRfT8/bAfXDKSE/A+eonWygH6y27i7NRMsyO+WNaTubl+C8D2ORIQ1FGvB/NrQU
zYlByZmPxzgaoMjMRyAqLMpt+YPPQxv3817n1Qx5Y84PmMAV2pRtGDZcXrtFUPeKMmbPWkyLut1+
A2SsQfj55pGJCP/eAXXAdF68JE2OQg9r3Q8xWC8f49TP1YAao24sh/WQocT2qbvx9cU79cYJu4JT
S9fZe9sCKvjbvOa/OChQay7rNe7prc7LNOu27Rnm99cvCYY9hp/pMnRdSh1T8czSVFwKrciDfl3b
5iN/agJAffYE7hmTJ+hlq3FdPyTO8UY9YFYjP4HXCjjwZJytvARLE2+FiDg4a91AApgO8OlDIdgg
CtCn7oEODVewSI1kK4K1JJkV5IihBnYkQ87pA/Q+bQjDetTNrvOZeHAHEjYiB6T19BDf8a0IGApV
sBuXQaz0mzOvDHbJZox7Stwhdw/eImkiXUkN4YEh085vhceGJXL2yJVrxA+Cl8SUv/TaM2MQZqY+
JmzvNkvJlNMtYiVNGdL80pYd3x0NvgO+FkD7A/ATROJ/T7tELIJbgYcyCxUGQsZuMC20kXDcExly
CRXpEHKjFOFLPFitD4AkwBrHdj2sHJk3x/KB0d1ZCEmv6it9L8oSYm6YLQJug0/TAcWlMyoQ4fpj
RhbVZQAWP3+DNvfJ92HjaSb22ZhNymRfFmoaPSb6zWi89Q4zrWzZ0JtSbiXbZPwaa6B3ISE71wSB
8LJ3LjL+nuiv4lVF5Mu1zXAoNH+AxCQKFzkX0harI5Vd52BWXPGY5Nn3KhJ9pn7pIcEtgQ2WSUFN
tzbwtSuubWJW77VJvn5JcBYjvw6VVmFYGEhNv4jd+pZ/bA/lfcc1YDQOOGhO1gVnMf9jlyDhx8TA
E6MP4onEdkaEcZyn5M6Bu5behvN736SphijKQWOZt9eFV3m+Lk38zHh7mL9uNvdyUBDp3JczDTsM
dAHFnr7ORSYK/rdMP/9ApLgh1TmxzmAkhS7sLy2d1HEAcIItG3TXUjHTYqqxSc/2lsDosj4Ij1ot
zsk7wBGshfA87SWgUwu01cJ3rPGrRI4WAcCmyCG6yDY/w1cjkjRp5i61o7Lz+s1n9eWR10v/FFTp
JU2tpHJZuf16HOPM7t4x2+kJRrgkUUIXjND9VJ2rRt1HYqGCd6ITxtUf840Ugxt+oQHSyMab0b3j
1Cm/4y6wukhF25/nGLN5hu/gEYQdU9EnbwIiH3s6QCmQSk5MYOxnubFEt3xquRxS+IIWbpi02maF
6BS9Ii8GdfI6au7TBl/8f/eoT+l7SvXvzisE+a44Az38gIIwIIMYYAC7+IdkS3VOsdsty/ypg1uw
Q/M9mawJx5100rLrGG2kHuXtYJaQJZIsXSwz8urKu1pyoSHwDXS+mDaMCnJjB5e56WJauBNrLDka
V6NZCEoMzZx4fIKzzlt6ixWC/lmGv5Iq/EsEOfPflqB5Tbdxyv/fViy0TnVUC5oCOOn7ER3ovj/j
9twNsOFNGoc6Z0L5zOn4lrEgbLG/tTwWX/5+4VPltbFY4ciE2WJKE/4Eu9fLX1F7phteCxu/vyYn
E6+Z4rrX3p3gXLH4vx0kVNCcvQoSfo1EiTfNuN2RE70QD1+2D0zRWIRWyexU7FA8f4BCPYA4eRpH
ByynWIQmVgvfNBr8XTPzodqF8NUVbdpzDD1ChhrrQqFQ2hOmxBO1nYNUcPCN6x+DkRy6YwZgzNdm
kWpigmjai90x9UN9KLzydYT2PdAT/pcDfnYn3scSPh46ZH1H7EXOPn3x/1LgUDPH9H5I251Ck450
fMkvBnLAfZSylUClYIXSJ2d9Yrlwa0MDisN4hw6DhCBgFV1K54ETyL45wVeuwPUg3vQIb7nEwu3G
mEXgkLD1CdlK5trxJR38ErCOXfa9HJxVqITdNjO1YMRcBCNdV4v4iOpXlY1x4Hi8Rg9nPZUdIUpy
YQ9UNqouVY+8NMN0lhTL5nGFT0ZRIjKtseW4EQa9FTditIt6Dc8vY8xgaHzk7H4Orq2nOXnVGe2G
+6TSI6ITwGKAAC6VeQzSaLEDLIJHBrJ8Qso8muCmC/ui25fX3yIpCb8u2FtbhSxt6NtUKx2TjMmL
N4E03qm87gUR/zpR5/OyDeXQDNjG555M7el2vf5lsHzKenDNr00DehEJ+BOunERrIhcETNyi+mW2
X7xxRsyvfeGdlwln8b699RrxFDxZMrRthFadyucy9f89gEXoODOH3AnhQmtaHu8Vu1i8ez9P7psO
kfZd9bHYkycYJO5PpNHW4KXHi717zlwUNULUWkfMwTBZ9cGXtEBXjSAdqzLAvVMYD+MInuv9EMM3
KGRYS952Li+Qa18GBDczXcNZm+x5gBctbdFHANGtksVbRiW5o6dHKpDLATBRvkciymAlctkDGmoG
bb5YV2nUUKxecvDyB0k0kio/AyxlDh7FsDrulHWfPSUQgDI0AeCT5FtAAxFN6KDGOoankJxQIT+r
vdIG98Z75EiYC1jnGWeC6RntM6PZmJD9Cy13lXdST4+C1V1cliccp1aLKufJM8/drlDsa6Retl3Z
zRWbD6mfGfkB9SV9TuYCi0GJhPbTJ8S4msMkp61Oq3sgN0U4XhkkJBRgs9wD4/jweCY6RDljCXFI
zEqNLuCREv2jFDefqVnW6uctF/xrPYJXW4Hfv9qoiPhP2EZPvkUQP4pXPtIeSd3uVfCze/Xu1ODa
kRNOko75+U7NpfQValGABzT1MbmUdaG3bxmIAjzTe7gEeUovDTb1oP6wZvWs1WgIPOlcSwzPfQhO
n0rcuSqGWOHsUaXTf9OBqbWNz4L+ezML0hjYNfzsFGFGtWGFIDhxdMcvzUQhCb7lKUZnkVMjAckY
0TSs2HBG5KHc1pZPsxbhcqzNUY4XpNmoUtg8qxQ+zwMSzUdtM+yNL3ykD+gFGLjIh9i4EzKSFhoi
eB+ZcPNugHnAt5lIMiOAjjEnUBpKts1+E7GFcQ58PhSOPPYmqJKdIWdE2EMnaGsNBPqGsqVHN9bP
vxHyQ9B55fDDszcmZU/IPynaKMf90n63eHhTT/zW2j2D58zvS4Z/xmK+XZWeL7itEnatr5/00w2Y
FHpuHJADDCbuilVg9daiOXD6HRva52uLJj/3eOsQY91VKxUcAEpeIxYH2VU52cE0P72cnhQZStG+
sRo+qNKKDajhzCzGL2Zviwrh1sitaxFxcBJNLynG3WrDNiMfpfGonr1sEy02QbHOQwIX24MZFgNK
dNAt5DXgbTwlXcw6fCQ9ILrOf44Z+Az9VWXCvQYwsLwZoCyajCRyt1bSISR8Qtn/jTIkU4tC8edE
woi4ZA4j5T9LuKcbkCSNrSVyARNU7B8a454IYzGW0SgHvSxYXlYnZiCYJuZYEqsps5P8bKR+ZYGF
S9idfcRnFcIbp/blWvjW+TsPiQ0l+EGP1N+SI9pr9YvNa6PAWFtXIxtEfIbfZP8/Hx3+mlM1ulOR
jaV/6FWyGRQTpDfe7EFvdRqewYD3pCecWVMXwzThUdmfvHn0iOxmVTNlgVmidSqKqhIbe2cYcjmA
lvilVTaXjpfwIuqZzP58gIme+o1SUBvtvT2PUriFJ0nSPy/qsT4qRZUwQYC+RleI/yU/MDhqUUcb
Sc22FdimbHf8emuaGQKPzn+G8Lr31YVe6WIpJUYoFo6FS9qD8LKUxW+4EH3WZUS6IDyLNnISJNeX
gMRV7pDPOOHa5JkRAq6Q5jQQ9oucinxxBrWVjaEsdGkLj/BFgo10KhdwRIHaDXx9r9/4TyskP5wf
IwA5L9hliRdC0aVpyLbTXfhQmW5OtXHo6MQndHCQ3MTkjf8GT69J6QNQAYfSTRjW6dAUQyXIMYdB
CSMtkWjqptje+88Loi53OuHTWHkKcfJCBIIICHS60X/TXwGPZ3ryeSwmNdSel0l8S/tIV0HnVkYb
IjzdK2Yy0hAhae7mAYPrTgpQYrMudTvNzb2jqxgph/+SDZPgPwJjanUVxhiHm47tKA8qkfYEf2ak
DKmm05AJ3PS2Y37jW681tOjsMOqW+O9K71j0rDogjAkLgAojMh/7iEwdrmzSQ8B3EAS9gObE6k+T
0gyqhDvr2fAFy2BL/Ncbgcm1jSsr1bbeRzr/2pBWmR8XypWTDD3WatD0iPfvAeDGVavWSBAY1gP/
/Rl3kaHwyI5IYG5V6XF91Gx/ux3AdeSAGsvL7ClcT0oXl9cBhNAfL9KPEvTP3IvcjKcsGliga6fF
UNKaTi1AWUCUUHZ0NJxk33ZjzA8C6SweYcomnHlRkv4Pxp/pgMLMxssZ03XnavCM9qNdTACk9/2O
XEhmVoazQZFaCvTFm8ri9I17Qp16UWM5harcO0bizmcNEQtTjzUTYRq/xBBi4NUjPnCGRCNS0R4z
HL5Fzef0ZEZw9Oy96whJJK4zP7rebQZNkhUNj0BLocXB/MedRVBz75mrvbhQbQVKABcFbBp1gS/K
Sb0fGm8Q0Zma5Aa/Rwzpk7dgQ26TPnJSqKa3DKmLCjF3Pm8EdZI8RrHv/dMLyk68jafTaun0W7D8
uFQ9dAOhuLMprMh3hSsPD/IZgnuwON0OM1WbhCNfkVDr0IYGlt9s0RbTzvYHapRZ8hV2nn+gggSv
ZDjVSviifVldQk9zHAQAAk0fW8rTPIzn0dZsvfA0uLsw/Pf5I5rxZfM+r/+ji5egt4ZWsgypvEkA
thN+WSajuYtqJp9STBXpXQTgRfaMq/Ltc0MGdGXzAIAdd32ZBuhy2NcP2nKJ6l8IB9v9J84aJ+eK
xL+ieC1o2oFIwFmhOVXqxfp3/iUKV23xclZAx+uvfLUwGNiuUonpmvfePq4alpXRob0DDhpXPIog
hspAw+tPZBUBrMAPSnsMYNx+Lx5q872YevvFo4K8X4b0G2Mtcc2UpfVYtpyheEye5czbuAgcSCMF
EhCt/pV6vX7KHH/oWlxLfV1O+jN0XiYckoZILOJOKQum25xsM9qFSkqKj4N4Ya0bnqv4XGJUKCGv
0XAdCRI2J+vP3RqJ5132vGjvkMpUQ5vlmFYBRT04vbHRBF3zI3BqJjuJ5iZ16CXMDPv2TGwXjAJq
ZmKvtLA59jxIyD85SsHw9ueAh1H9vNumG9s8ibDwDBclSNyc6rf/U73EH5gfyyCuGMQze7v+OOay
+A81leY6ZfqtK07DjLyMPWkmESY3kCFc8exhhP6oEWTWie6p562Od5d5daDBTtYnwLDZAECG0MIv
NqwC7+ofrgQ2ptaBfRw0/HzynFdQMOQwNK7mmOLzI6rB0UIG0S2L5/foA0tqzRSvbR0pwZH+TVZ7
gYUcwi/RIsciQ0YcooXcdlzkbdgs1O0P4d7+VaVvZ/EDVA/wEskTlHHzExX+FKFisNvzWVXjLvxf
BWCndLiyC7FPF9WNXX6j8TuD4Q9Dy1KkyKq/w9TRPS7iIAVnqAM/rEu1kKXhSoHT0/HFVYNW7i5E
Ch2z8iF4WhLEojhOTwJr/sImJ7lPB6iKj1y4vGjGlvQB+ycZCRVXjREX4mkfsBi9aqe58f8IJkTD
XPZOowJcoBWkiViCLEj7un8EFnEoNqGxVxscGoHtbXYDOtB+iwfgah4iqS04Qj/bc3rYUhPMWO4L
43xZV2+917yBDcUWtdU0ROLvGUyXHKqnJ9lAH0ygTClkOKfjjmIECCDPA0zCs7gD4G0nQuh2PsRm
pjDyNCuKtojUTkqj8+qlSVDfb9jRkKZU4uQuHUqovcwHJeMkLiBnEvrdfrOzTbncrKVxBjnJmLGN
inD2I/oOW4KYJuNIzBxJBfbMB39jY/fmvvKzL40V1wQgsOtTFncOWLcghkTlOrboGfqjL8vIBRE1
/PwPCZTZKjtyU8aNdO/4jqa9szleyWrCdYhTFfH0NTcunb0qwptLFAsHKF0jglJO+tk9Fz1PhBeK
nSdeTuzJe4ygterEitZG6ZPa21NgSpiYb6JPAfgt9ah+xej5RJ7J/FBT0WWrB1zXu9CgvmbyCJB8
CXsROiKPp7F0KOyNtOhQUTq5T9EpTcShozA0ElfkcuX4unYRQYRP4H69wYZHXdUSyTOMesxcosg4
bkW2DB5wbTXIj4TK1tyZ7z2M99/RrnTfktKquScJMf7hoR443do+oWJJ6f2xm7JUlL+pN9jb74j3
U4WMntkbzthqL552fFQfCSL0JWNLTghVg32RcGc3Mr/Xm7QPXPK5R8oh/A5cPPa5AfF45dEg0LV7
YmsY/O6HuGqMzlc4TeP92Zn/skP6qO/j+xJZUSdWghMg4O0gWYajxhR+D83Hu4yHxBniVL4fuHJs
vgHM+TeDEGYCAo9lGbEUCUfnoQKhxtt2H5TmbZqPPpU4L+Aj5kTE1iLmYKpUvL2JtVwUlkwS1wij
LE9/eYLKVIbGFJNcqx1RFowmMl3fiKukKbuiR1pwjD8kiJFaG262FQGTAiAr+fMLFFyn+HpCIzN/
RUQVibYlfZw6+QX5wUB4avAG1H2Cx7YUXR0oAxOw5QBHJXrg7PHrPwKP0fNF5J3YOyj4lQKHoY0H
U2fHgud7yj6ZhYURe6RdrPc1TEo/uHBD0MpH++9zirAjhQI6OFxZ8wRdtocDmFnAMERD540zhQLn
DcKrk05gm5iYiqkCYWdEu0ejh76IwVJ0JTOmCZyHilSUIl8lh6w18J7Ll5VUyPkfplJ1dLSCx5QT
yjzTDsYrKk/lm0NyRlrs6CA29D+RHhJi8+EaPqm4A61NCD7m/TKTQDrFM9HUhp/C2/DKrH75yKmG
T+hy3VZz0Dw8sTxJr3UGLuV5L8PN5+FmVGlteo75ar+yn3gUXMCwBwfLI/r/fiuFf0HdBOOUjzF7
Twe0zW+SuX/esS19tecIGKinlRsjNcOw5xQ2m8OAH/97DaPu7eaCyiemTG4rKNFVzW3YnnjFjY4a
PszTSY5SmWvBqCWCQ4K2j2XC6tfb6qBivgnVLlpdAC35in4RcNmA2kU2mERTaSTK6+hGiK+o0Deg
f73ed89rNW1tpSrU8YbvENGPYIQf9Zu+81r9twQNXNIJZlk350uRNF8/fb8a+T4tyUwxX3osrL+R
/ly30FQR5nPKp7MGImv0n+xsJoRHguSmNjwT3kOrrXVt00zqIpXTpxt4MVl9+3SqqnqFuG6Yl0F4
ZsoMImqmiIY1Y5/thKlboDM7hN9tmcwhpSfRTmtct3BqOnaTxKOlwG5oD/kwO8wUkDEmluRfs2z/
/4Br/SmOAFh/JwfbKUqP/iJZNXGvRf6daxiPjN1F6gMT/DjCknOCSMJGvc0QBSXYIFfBdal2zwrg
Q7jE2RTDKwOvSx9nQ8HJ7wW/M94kQTKtbJJ7IsjJiLwePW7lE1QdgnCXBqIrlsUNcd5RWJtta5f9
twkHF+Vh8eWoW97eLxn4V4eg5wHba4Rkx/oW1yENeIKaLAvAjkf5dm5T+hND9el1f+wv0VYQ802Y
SKKf06TVmn3Uzr1kaxR9XrJ7ahhVxMD7tj2o/FMWT0IVb8tQ3GQHS4SRqcz7q0GpNYccGueEFkMq
PUHVL52LrZ6seDrMksM/v+K/Km8+Qn855wQfAxqN5Z2u8xAZ+4WwhH2N2knSSX4rISEbBr2cOXiU
R2HvemNXn71eRIVR1A+XenjO6j+CDXqe7+t0u8qxCf0n4EFoo63vyQ26Rg0zqXUbzcs73JSurRk/
zsIcPTgEqBHLPbI8v+iZ/fIlRLcCGmjXZZQvw3hwU3M/LHY8mFDjbNY50+A0g1NLufGZ1oXiHJad
R0E9nZWhesoVJsgYbH+ZqsLGAYnjCWyvmY72s3vUgw5R/LWywlUbabdCKkKimhGD0llixAXKuBGR
kGQ+gJHSEIl/WWxD/UguHXMqSjsw/EtXIQ6erk12h+QqcXadWvl29dQDIoxhFvLRBX2U77eDx/xz
JPNUzPOog7KiAHmeYVV2fKG58oAUwbs0XMdKxuF1QEKovuTVLQkq1goePs4yR0jWswWrrmMTw9iU
Sv1tlSHhwQZtJxRW4Bril4djCZ3epxVF7kqHeopyTMvf6FvlXnpEnwR5/AXdllqnylqPvVMYen09
nbBTeFOpyYr1JRpU5mFvQgq7pjsNtNvOljThCJZfiT44AvMu0LHsJEXMfZtIvpQpocE3MKct2yVa
A8JYgeOIv90SwOZLsrAU3IeKqckc3ufXV8UesZ4vR6zzziENI6O9WmXk80FDR8u2oSf6NS/UMnDw
Pm1zxGRhk1XfmdHxvl4cgc8YTzo8fNzMtKQKP5klHerixpiA/LCfPtk4P2MCHvadmBxvyDfwgHsT
2o8VPH2RQGqMe3dTL9Fms61lylXuZL9ADH0f5qMEfckukO5aBd60ZliR/cWK9ZkkE8BVlIbrNIGw
zg/SQc3kkVvyYXd+aH5KSZgK4isa2egKJ8zrvhky3z77uWlkuL6IdWKyB86xTZ7tlnMLPzUJ5ftK
OfdHXNjbGz3jvzSAK1t/mr+aBAfryJa7dCq5pifw4+KFbZIZr0FFGUhE3xg3kAzeYquZRG7EH+/D
FjXlk96MV+4+ig+LYtsXefTBJX9O9fRdyuNd4l7/B92R+T2Y65pPwFy7pyuKpzGGHzLNJb2kPlna
5E1QTWteYzqnWeg7Jxbc+oJIqwqq3zP+lWoyx1BcBg2MQxTEmMgkru6xKVBOA6N4FZ7+idDCyKA2
Jl7Ml4V+Cwgq143Q3izLPucBW35IDjy7TJaKWa2i39W+kY6DYtTfNAvjEAMZOwejUkppJzJcq50v
bKI1acCrHcTzjg8mgnHkZ5AYOwAecfrFR246fduOfmw0Bbbv+nWe4FLvKwPhpOJCcfjs+GlNVliH
gs/WQFHp4vaolDt7OkTBaGzxYheReOws80ojiT1LVrt0JowJAm1dIgvI3lFDMIM8FVTchl9n3Bsa
P/H77Qz5xyAddHVpjHwkxl/SwVFKxzkShrGETirRLmVAsAMbscUld9QQ+1AKiLWzq16S2qxLOunn
pZGMsjWxAzh/i+0Uhi8mYoca05DWcQiIpeBco17sZf95iyO9Z7NieL7Y6R2Z3MJdeCGsLMbhcQ+t
76GhtrubZFfba0iH6zPrI/Jr69s9b5AhDwgAnbaY7QJolM+wJYIg1+Qo1sCGF2ia9sphDYYjJuV4
Q+/p5pyim7enzmwUH88Ky3jA6Gc6srEiFkBvkBdftdK+DSWyByrbTDTEdYjLOwRSyhuKVY1x7JK9
CN+jcERA5GsLSIp9xTdB9uJkybszYC3fB/vF7a+V9pfTiLQFJpEP+kp9I3n/PhUUCtNTBH5+o5aQ
ak66TE3OXb8MVelSYVaEdjQTaYI2aWyikIJJVC2fUZXgtnKZqAnP+mWDuggCTf4mm71KoxEOtWyP
30rqPL+ULuH9wMct1nVEgvs0l/tj5+w+Sc/xrsEK4tLlVV0SfyP4g0d3kXYPzoZRWbcCcOsaumuG
yyIfLlUGImugJrAlMmptN+Bku3Upk0dUqq0mneczUSprhDzE0HF7gzC0Aju9EKlsfyJCHnjTvjZN
1JL5rrphPkwm0dtiQ/VwALA/q7AoXKM7MP39k9He4tsZPLshUBUHwI2/+eiJ0cWmHEWY14ov/gce
CzhsE/D8edcJXLwqg+IfhzTfPD8SRGw+QCtk4izuLcRsEEqsOgFCXolUggmo3ccIkGJzRPYkMoF6
R+j8TT1qeGoq2sSQsimMQdXH5mYaJKBIh9jnQ+VJZ6nFU68fSU5EhTEhgyOeBlXLCdaNuzWQgPkI
0tsc3h4VGu2W1LCLbWYI0x91mI2XkYb7KP9NtbUjQFvujMRKGndMdOosdYNWW0E4QMmBnQlFuwBY
Gm3SexjNNY5sCgLzHwHwKErIHbtk24JPsSEWZ5Nen1mdREcEX5iqRFFZJLzL90+ZTfLdp0v3tuSi
TYLmQR8LLT5+TpcF1nxFct/nT5E32hulw3h3GNXMR1NwX2YfVDbH/rhGgrNF6c4mcgBeYBt3M8+z
D7m8+rqw5T+lMg85Ax7WwCls/blU2kA4TUTweAJpyBvR0sszkZdA5xWWOgUS64d8yDGjtdrJOgS3
3x3Tqgb6qj68tP8V1qCoWaYvcNbWd0Uq42bC0UK7VOk8IbM2dsa6sYau0pkT1DYvn3o6WU4SWGkz
cw0vGJKNdql4D2dDlorCTosRWhIDuZF/RrfOxTIDT4gdydJe7bxRUOKTijKdfo0tfXoYnvK5SNnx
gMyimv1ILq2OgcMNwNTaz6lQAJsM7HLgmV0Z1M8WTpci/YNNI95cQxUj9M6ok5Vktnk7Ph2uvDuU
z0hE4Srqjlni1JvnUsYhweLPe04aRVUKicJ31DtKOPr5LmWtpUqLqOE+8qJJsNnQyBbcUj/vJ5w+
5mWdpwxtExbelhmRLJ17/QGyZzz4PEub10xEY8PZ2mftcHz2SOeO3yJvfulk2LFDvnkTx865vpb6
Iiw6ov14KSqoRH8ggbutUwmz21jsMyUAqMv4BVS7FLBtuwDG+rFdPvg677TP8y2Z0uWMm3KK/uH6
lxKJCermP03zHYfEHeuCewyRDC8nHJsDxDHs0tvW56GewNAPB993VLH8EvuRGBR0igv0BtE7P/AG
sf3j1vrF6dIyDw+txiGUZ/6/zjLIVsUv87RGyRpRfBGKZnuJa9sj/pn7BO511FYxtmBH+8XY/M1n
rBEoJMVKoRvWTUAgvTdzoiD1Zw+hI7gQfkKvLjnLGuEjGP5ols7dxX5tGkOXTQ2OmnIW5OnQhkRS
wNofbxxV6xc4qfdnolh2Y4V8vNS3rvKVXyQaSzh6kRJx/Saj+232S31nAQEi1CId8CRpuwfGHles
8XP8nqT91E2b7eiJ806ZK9F+7krHgjtv4yLvE7xHO0x6maiPYmxVi3ayXXhIK6MQGS5HGmHTU9Ic
JExAxdt6YkJsUF4VOhUX/GpteQBe3WxtAL11fBqOvytDSos9XPoLyEmXTBnP+gMQmn9y5g1ukWdQ
pehLq8GAtvDCS2eNG+iEbvI/5fGbXoTGonC3gsBTnV8acm/4iAR5VCp6vOWTywzPp26B8eWvl6V/
uLB5+NhgVitjRHmFBQzwnf+xUCBWNXgUSS7flntl8nyO2Z3aSvATN1BPDy33CeDgpOFgbPDWq9NK
kHoeqLbvccu0R0LvfAFuvj+Kd2G4OPwPt0C5+YM6kWiTf6cXpL0HmMBvZpPlIbz6XsCWuhrvcLfK
EqqX4EY97n48leK/bits9tGQ5mEAJMD2fDhvfZIziYS/djqVwVwQBkFH9ZYc+QAE2bVg5MsUDVKr
BWH9HfWVBAiLm4+nPzhpzeux4uV+g1KnHxo/F8kWC/K8AYZJMJn0/6jU6DPP5TIDeD49SEPotUgn
sKN7e27FozHgSRcyVrW/LWLaoPM/NIATTu21QVjyGAGYJdrW6AIYffxL0emItO/ULYB3ivqHcGCO
14a+BPZsNuFz/tzzxIUqGBEzXfEBg5KJYRQmm4k1Ks5BKpABVmpte0HNwFWqtPrueqmd36hBgbcs
v8aZJ9tlgX16dR2rEt+9kOjXkX2btnFKhk4yGkm5FH5J6R/lPtEYtoaSwfKsK3YmPjG6wCwhXQAf
DmXGJL3xie6HnC3vij8vZFIzpNWCb7kwjdPntO/lakSLjj0d25ubQSblAeHKyDnYe2bDVUOXHzQg
cwkw4nhkNHhlipTMnHCpVldITbP5dUXOwIaVvxMZUO6M8xyqkZCM3908yZyOAK7yYr7r3hb38vK6
KjAlLLudVcBvNGxmlarsqznvkj/WbMNyJOG0yDcNaoPAPlFtw8pj5gdeKpHG62TIK3LuqOTTf+Nb
mmUFAOkmqhBk4pNkoCW0wi3Xem4w193t/MfbnPjT5SHrHJMUMRn3+VxCaMoLdovUbT93kARCrYw2
tktbZ0cdgNek+9RRvr0O3QsA3pzZqkGkXMmPwW+KYrII0u7H1IBXOGHzD2HbAKODcEFLyBCX+W9C
yKk9yAsWKvSEHg4eyMH/kasMmpc51dZ13sgyyJ7Nt2XJVUuVXjfDCD/qphF5dWkpjWzi44zqoB/W
KmSh9HKOW8g49Qvvnri6VFerods63gDzkf7t0l2bKGiVr5CHgIOyitHdyDq4c67ZsRGakt0DhWaT
mS4jtYNSod/6PcPUFx8x2voT2M926e/Q8wf8CF2KmFE/5Cz0XoKwHbd3dGrMLLdZydW4nj+t3r2i
OXhvn5e5yV/qRocTySjqZmiHlg2zMRFw1cYh94lqLEozRaFCI16YW4TSrBZcaVVk85oDb1zemCeG
AUf2zkENot/JeP+s51gcTe+4L5T68kBay3N+BM13ZM4dUefX/sfchhqMlBZEh5ZJFpkmR3WYsC+t
XBPJL24Mhc4cKhZS4rI/SZUfsnpQCunN4/dyhs+ZgeV0ntvsA2jXoXWzQDvwBngCQv+A+Ee4H0p/
vjocKsNnMPjfcptkU1NiGk3SPcn+YQpynGSeoUtDUdIPReS28RNQn8RpGAaRoJ+KipoUYQZHjLlC
hkv45BhHAp+se4Hx3v9V7McOy8QR/uVpdAba8xlGu5HJpVGfE/CWGhYY6LP9uj7tZ/EXsqFbQtUs
K10SfFukI0GTa9IZtrFWlUz/ycNlq0QqMM0Ry0vX1hgbtrTT3xKit+aUkcJaEwhOBaKYmYjAST7S
1LvKUSyzDCAcUYlpipgtJGsTu68kWznMKaTKkGovEdPPDzWnvQVI/By4FX4JQcWq6NnBtdJitDva
Fhq9WEhxV3d6IXBzwkQ8G+cg4krQjScRSlEao/VJg1Eq7HN1/YdxrTCPPUwxAyr5RdZpMM7CcNnu
2/lsN6HFepxXwQDEjAUGL3Iy+8VW1NuzBrhYOwDzdvAuOBcUb92Myl2+34a2xMlzdoVBC+k1pNoJ
84uNE1z74uVprCXNK3hBPmTFfJTSAVuLC08EE9RIdzu9YfsAHGSYre/TC3SAt+4ZqSZqn93/9oPI
q/bHkgIhe4y7HvE+GFGa4+dNhlZdcwXnWPeaIpmmGPVBfQZIEvnMpEUU1Ywe5WYJ/xSCf2xi8G5W
nBf9rAqGcok+XkFbLA16aVXw3OFcg/rBSWIPAOnVT+Lu/8X6jj0IrC46jMGK5KgPxQezVRWlTE3W
b9RrkXOaslLJhb47U4RIqPjzBkfqqeZpgWfT1BbAP6NowdxxjWBb9E5wxLQ46h6dozjJdb3UmsPC
odPAPp7CaOmA20YA34cJMP4eyvublhdHns93F6liAtvtl37/+QQX9t3vM62gqwwgvk6zEgDS72/B
H5phmPGLs2+Rg6scHS04YjZjyGYUBs0XduCk1vNhi96WwSYhX158JS8nTlz7pJs7TvR4KPBqZ9uY
dthwIiAXMfu2xXSQhg/a8xrTXSglimes/sTDZu0+prlbQlgGzeMMzEUW7onOPijEjpck2CNGWmsn
FCANLiXeDbCQ18wyhpntXsC5cQFylNJp+5Hp8FUImov/z1xyBSsXmaVLSGyyTAePYvWvxLlZpPOm
kdURDCPKzNsbHPMtxCQ2BF7tkldO1Jl1J53ayDaXfkMuxnrseyEflPAHWl2Ah6NB7pRMTzIGJBBF
LsRyGuuXDj1hv0Jpm3npG2GpUPdQJoNEc8nxzBbLDzJynV5CLz0Izh1LuqRtLa4U+56y9liV6hwa
VNypC0EvbSXsoROuKvTMRfhIYYyRM9MnaUC5dP1d/Jgq8GiL474I8Khljrs/NE7uHkc+w/8hCCR+
oVC1cA+Wl4iysZaRInhCygq6Q8ek1sVzB5K3snJleMTECmwlUFtGS3aaGWHqNNjh1/co4swst0vl
r8hmeq5w2fdtJbbX0RAQS9vK0NXOTQnfS41sjVMPAEThuqoufFHJ0qpy7rQTZygjbpp0+foLg6Gq
al08Tt2YhzG+76zo/uvNbVpPsHbyzn93/NQi0TyJ5OpUyG62AiXY+gnrOXRXfH94Rjt8eWWxvfbV
YMZLCNg+cNoGu5pFmhDE4di0HbA2krepiRZqs3qPT2p6RV3wk8Bk8f9Q2aX+oxwL550vsKxfbkoI
9B95ON4Qy0dKfImiZqs1r9Ute8XDVBOzMBz3XwgdN9KAMVY2QNjxFw5/+ow8JSrlyOI+q43wkfxQ
LoklfisFbAQT6u47P5PFZMX04XoryVaKOJghPgrpJ7XS2Xx3oaT1aEB4RHNic/RVtOFBa4+dCU85
O0gkkoGoGLsWJZYChC/iEKD+p3MZB4+zJPf2KlJK5dw3GdJfk53JZb0tGV7qSww9wWzzHWZCuAQy
DBhjDCqBEEFqO5Hoj6to3iarlxZi7RJa1Aq2V6ur4ABP+gW8z2I68REemZZgwnPHQLeXCqhm0Jqm
/x/jUo4afc2Wdb+fMD/Yh+9PHR6SlPG5GcVz4yGA2gQaoLWbVProJ4gBlwecMUq/O6MrMEyky5Hc
J9ThD/NuvxiH8WQeavUS/QhO7vIuqut0WOMQY8YtPXEWVpAghDLheAjaOncDJidcWmeQMVJRUEap
qejMrRqI9QgKdmk9PYjUZ4iOIr40i0q2Oh9s7TM6ozaOcWSex73ptcpj3AZ6xEPEtJn0EHZTC/yF
GUjJHmQ+bSpZ8HtGKVZQNCJbuN091xK4yti+B76fuGspYT/BXfXI9oF7QSX23dO+BVa96BTS/Dtt
aIkGNdamOidH10mHbSN3mPArx8RnTrVnkDrirNf50ZUczAEo1OrMJVQWDCm2CvQxChBx2oQl7TyV
OgeEH9FL/mN8l9zq/GRW5tVenfoA48rb6l9G+LZRl8kYjQCWw9wIUwNRpMnWaWIwXdrL6x7WPglt
aM3XP1s9t0JQd1YZb/z8aJXMRVxxcOXhUdkxoladQMixDSmLdBbIVYatGwPxodkPSX2nnJM463DZ
lkR7YwmRVdzJR5sGaL92Mz1JiFpNFKgvbKGtgPCLJ9pp9VljqYJtzbTnU54h2RF7OfNSjXEekiFd
rm4L/5kQPulRZqtRDJdip2DQKopUPo3OMXU+oZ59kjVYecGf9N43uIH4dtu1Yb57SeU0EgpTT1Eo
JQtKtEtApwivz5IkawR0TOLz5Z5BeAcAoHNGy+6TFPlz/wLUrOVmNwlT663921PjuDKbyJCdvDxu
B7i/S85n8Ha3k1vntlkC7xnQcpo+ekO8gzt+lPH+uk8vV0u723wHO8ddkOgKceylSk6h5vF7qk7A
slJAcTf3P2GQmWM7QXQW9xY9kcKaLqX6mHWYemZkB5NL7E6QOtY/6Sfd75cDwgT5c9WOBeG45raO
oUcReoo05PX6s0TQ7X0Hm116cVJywvdZ4lUnRjQLduc7gDJyU1WMoX8Gr7NdjwATQPbZn5zNlcMw
92ngc5ibKVKNTsKs1rbGFMy1Z2xy7MJ4MVNBsd8U2hIq8XTMUQFJilLhxrKaembRjw2JxNIX24f+
U5snNwz3dofpCHtFMJ2T3VBPT+quXUARjDV2NlpT9XROnAGdl99uxaPSnpxlKX3fk0NgmAE4D5OH
F5Gwd6KNKjh9YAOFrqa0CaWuc6sCGE18mI/1tobo5kjJ6R+keSvhhdM9LqT4XL7MjNYiGYRbHbq3
/rw8JmvSCl4DmtU4PzwSOwA3lHQvsv9ZjvdmhYvXi+ALmW/Yz0856l0LFHDqsQl7GqC0D7gfNT6d
LthJvEbivMf8d6B3ledw/pKxzBWX1HQikTv1Wb1uDJePjaFRrtTQxXj6ongVMTVzt9CB4dJ7P6UB
99sFnazgYt2IuJnkax17YbSBQNyPBQM7ohvwXsJpgTmeSBeCWaPZ+8os+lHKKkiiWcKLAIU/eP0m
wZWy42VY2zWuE047rdy+W+ikLEeobPVWtq+H46sVl5lQeOyARLPSJxC8sCsPJ9YXVo6eU9dLF9aP
+w/kWbn0iPq6FzQuaixEDWoIF3Lc2v7i2JNkq2VRgTpYql6GSBhITOCLCuzAkwW5StpXv4tMr25W
wo6KOq5fkrKCY/sLHRiTfTb68bXt2/47iqkEWvuNect/B3YKBlYDNpaudb6r+q0sb6GgCtcPiK+G
lWE0UC36c7I76lZPv3YqWTBe6FKejTAxT2GcxGUK2nsm6q8D3+1YvdXTC7XSLQWqc9lflqODUlyS
BG08aeub74erW107sWj4vMVeqstvy8E+J7ZiGuboqKB+hpS3AALwlNV6Wsq4dpASgmzTrRUVsMMP
kmz2kAvY5ULJVhA5ViobR4jCH0yMHqdfXX/kHZ+IUUn+0TpYHSs8ivpRw1Jq0kUbQDEdIHrp0EQc
KkI3CUZhS8ZnR8WCVEaE+Fp8nm/FvYsT4tgefneSVNplr+DabaP2LVbY2NGbsrGdi2ZhONtTTqTO
VuSSf+UKQ+PyKQPwIW/IqYezJMQk/m9W8uyaL6V7oKpgFrfa4gYF66LKofEA/Ay4axbxyFz74UJC
ROawKQSyZVlGUzX3R3HmIekpdF9QuHekTM1b46iMTNCd6ybW6eL+buB63cBKVhZJu+xGO7uky9wP
LHb3qMlQaQ4mplz3oM6FVoImwbVutLV02uj8/S5Y2lgzZeshkNKm5G8F3cSE/oXP54bl3bRunkyA
K8LWMXT+SFRVBX/w+nbxVz/NoQHobH8PGtBlVs/upFkct7e2mo6mApI0mUNowrDWBHuEHvvSpZdB
8I/9gx88I7xmGcX8dDnMJdH951SpZBMeE8bOKtQfPUnvbRWdz6YwOH/2CAw2lg/UZwBig+4WvsSe
QeK0jucF5rarub+SmRS8cHzXcr+npt5ynHhMSLc9j/pDNcrHBreL2nvqn1Hc4wEC+gqrStHT4kqq
1CmCMXSNJJWj+USH0OSKWVmokyXbtmP9UBWtThi58trFs6ZAdxiqUB0f7+fVL8gF/0a83AHheFu3
UEJMTDAhAABowCzLMEQEXmZgWKJEyxu8exnzefNXSrjHF8WFpMaX856J2fk2FlYhNp69gSyaDatt
iWhvcZNBSA6vWgCMrcnAlstdy7aN5yftrjz8s+73lcxsCncAeYw8fZkg/p96zdgZrBBiLBM4kygU
NnOGLsvzS0VVYaq9bUe0Y49TrIzU3hrHk4kozqlLaTk2aQkREgQllVherqYECM0OTirmSf7g+0TG
bzp4SZZRfqgjmoJvjWALSoXOISttq1847nM7Y+uzd6nw0z9LyR/sVTligh5g+ygQMZAOsWSrrDiR
vI6d7Wp/BqUgPcPygX+q8EcK/cycp4MZcByFoS17OacjLmg6wrYBAdb9q7oEADITI0+XfzPk670U
BSKaxgoRWo8A/CqD3OiAUxrWG6RSok7uChdA2XI7/jd7yjEPbk8b+TpRJ/ILeXa0VIJrpQjxdZVA
5EGK7uWyPp7t9MeLVeRUm1dKvXKajdH5LctCoSVq0f3AvyGHGpcdAXhACfl/q97BVIY1Ra/rEUdp
+UXzIxIq9B8rp0NXeiG49fDLfCvcNsm0AlqVsUhRQX4Bm/Sx36kRlkBxt+idIKvKq5MYWFbUWsww
MeMJDYKCo1+2QipO1WdIDO2UNhuaHCJjRPguwHH01vpuE8RJEVhIpLmPRf3thuA+Bw5NDJMOeWuk
NWPpyiPA0Ex0xj1TxZmB3D/9ajmoNeZGy+mi0Fme6ig08rAKndTjaO2LekSYYfj1fRb4nYe6TeD8
ryVzbBEwGprwbnxdmkivssj3EmtDCmAaJHSNzpQa9nW60l9wn/vd0mSCSHhk3pTkFuMUW1Kf5Wmw
Kx8clT9uIKmctgDhyZcb5W+8dhORftNrWTdyazkNEZ/OfQHmCFrxXa7Yf1UpK+t2AIffLyhuYCA8
4rn76XF4MK0ahV6z4HVX++sb6TJoXkrk2qjyxrV2Va4+BispPbfhcCrw/WxreoG65aPt0+dom+tH
C4GND4Yh6ag3L2qKA1wfesGEn4Nr3j9JbB7E9M+n+giNnPGcbD4f98Ry/tiI9W+TzpmWXAec2De9
HgZcSQ/BdpgepMvmsoHSoDy8MM6qasFDtX+W2YbDnQBrhSXvq4EbZtndX93912bqWtGyRe/Mh/N1
nB0oCQ2NfnbDuykfr29vVyQH21BreB4Mi2MC0nDJYO5N/eKrGS3d/eL+ycbCzq6jOHTo/9qNkfBm
IoX3fgoRkR+Y3rSzSMqiUSpHdV07dyGMOWxqMy9nZ3/RzezCabxvPeTVzCYdmmLk1GQXkyv+xISs
uIObSroxu0g8a6RJA38WPennh9KrHthfoRRbCYESBxXHVCTt3PWJSHTP2cUdk6zmz14q+N4brcdF
rU3Htex3jhSjX0xPJSyb054UG+yuALG6Cmpxr4kiFNDNFV0JpRdzVTzMTH5w1KK01nHrgoDG/LGj
gdy9XjQBrSt+psn7GgNlzjwgFkUYc43Ug6UBJ5nf7hWSiHfJwHItmVDoIMQPqNfc0sYOAF1FKd+B
9Lxzt4o22GKMhEkmBnQpCAxx+npHnDOLxM6tZQyU9C0fyKDgMwWmLgUNSTmuqnfrbQFJwuGQOlKj
m8EmFLLI493hc/BUjp5Bg9p1bh555xnN+svZij783sRDX2xqfMOc9lJE3Rflhy+Hx8Bq8H1ThRC7
oCXZFLGSSZaic8jEOvoU+bsQx3kXz9Ke2r8eGY2vGPtxLvlefhRLy1NTFVuXuIcMP0WbThLH6Rwo
EEXkIZcAX+zmJtScbASaoqDWfC0NY5JxM1EoA8UybSp44txnQKJOhK0R3elDRfPfemtOj9Dg1/oc
OjgP3V5Bb2BHHY0H9aI7B66AdgdvZBBP3L2vxUlj1vAwZZP39djFCv251GphyWJusy3Ijv9Rqu3p
iKEkO9iSUrfBN0zFSk5gagexSABn6Clh8WNH0cM1UfUDf3vIlTayVt59Mihfq0JMLjR0VwtPTIxe
Qp01RFeZ/m9+cve3b+EdbhBG04QMH/u08DijR6FbXrwxe9BFxIiCXooYDbyxinyTENy8dmDxzYGD
aE/JNYAE1RkkjJTt5bpTTW52o+ipFgNrcBqvAFSPoOtMPF8YfxlFmHRdjpcpRQtCUR3qCqwvf3nA
Gj9EJHrbWtjzmKuVKzia/Kcy76xrg6OMAxT2JsvKBxEbGdeOTEN+gfApaWYmt0FCKoxtgkGC04Jo
Yi0aW5paZZAMtTFKF2Do4JBaY4epp3KU3UzrqpR1iqq/i5pqlEQeDWJ7d9DuDFooMojD4oLOGF9M
aZXFAPWZuRpNm2KQOArOK/KrPUyPjdZbQKBzT02TEFfdNR/8vdKtkde5Q+4HpA957GF5Nnb+UU11
4Y0+yRNYQlpcJGmdW+zFdqwp7DIBDVIoEY04d+cQctRE1ewr0lBO2op9CiceI9Sxfm7OF97/ByzF
muxCZ8dB2SSPO5V9gnoIFkL2UyWdsEyylghCFAjD25efplNR/mub/UnZMRZ3ImxmdG5gLgv29mmM
9GEK1WZHM3VLIR/Uv1yI+Ao/SgLfX7yajnI8PgcgFBNl0jhKUh8MHRGkLGfddOoOyBVhGRsg2LGQ
Vwiu8cAPo+8Gfaf/piSlWUxx1XxnM+cMKRZGd8KjIWVv2ZiJ3f8c1T0FD0ss4yINucK7lQl71yPh
Zgt8yt97UkUpXyimgpxo+jv5aTzoHujUAmsxfwDpaeIR+novMhgTgf/9zQG96ExUlD+c7CVD08f5
4eNtURN0ewbtgGZEWgv62VTw5c/Qy7DZdC/vjWDJ3QRgZ+7kTH+xjyyO7tWcfU/06yiyVnZi5sO9
pQYvSajIJRx766V6aM6qXoeYsuwXN3EgTFHBhSrSzVlmdx6WBcAEbxKmg0gL8zWsb8UyNoqQlUPe
dqi6hOBB2gSI+XKT7O8BCVBoi9sE68K48OQG8dAtcWPRFDFoh3uCLscthMfL6JkJnUeOVsVUYfey
bvYwjKElPSIp/VwcLpmEMCwP8Wdzzc4MmOGli+TgAkhssiRr4NiJzJegj0lDFBFpR1TVik83DBfA
HgC6Ag6Sh7yiwhCwBkZdGNK7eo/z31/hMDHWznjYWtHf412KrWqPTbONKZQUSBLyzBp+uOyvYwGI
rBsulEb7k+MjR7bcfqgRzL4Uft/oAFe4NpVczThijHs8+gSkxcfHf1aD7a/TNN66NtFlEZs/3jc1
T06vYY09fXhZYDI65aL4qmROa08rWopRwfMsh5baiEU4zO2YDVLlgyOGGFyo+JPymElrxZ5o3HDC
JQO0WO1prfX8PgZ1pzPe2jKBaysSR47PfO+r72GLhzbynkL3ukMDTRxOphJCyM1f3v/eVf0I0bM7
8IkJJlna40oDzBAqiqrJ2Dsxm5Mm9oZ1rt5TUf/Rk6bvp2UMfsnvuclZwosXYIki4E6m8Lf+mwbv
fn+051MYm2Lncm5QT51kiOeoY22AfTCfRJcdGpaknXxHxWnPfPoDkuxCM8W8XJ1BbGuGyT0jPAfj
JSlQGhzouw1++MqsiOzMEZj6yehlhkwL5lBpHJv88SDfUjjN1gDyI+HFb9tZn7z75n9jkYKHFj6d
pIYNVFRTvghBByw95MUDJCwkqUxj+TWFWc84NsNPmQWU5PbExSMJ0SGf/tfl0nwaNkM1RfHDdvqI
ET+eiWCxqiWiAoAfnL3XE0gVvizQudyejdfEfPhBUvOZWdgohvk0B924sdiZp6Ic7xhsu7YZyZc8
10xhEl9sZ5w4q5es/jr/NAierxiX/92zxqfmoA5ndP979tPjdVbjV028IgvRvFG+vRrthxTUu+sr
a4vD409VVDDR1sn9cQZcuxnZXpW93AGq4jV2hj++gnxSqGNSAN0U4OTk0hxxvk5PZU4czp00yH/9
kF0JkW+3JlEnZeZs+1cTmvc2k5a7w/xv7lLWlgUOv/81zPK1bsrw6VT2HksEUWDSoO05F1KFIIu8
QchyAWQ4FrkjDDNzgSz4sdIuln9h46hRykN1mQCUTsvQjrpEVEbYwUGmU2RUqu+qY3DYOeX6JtFs
HFe+21bKX1gRTCNxwbBBte6BnvNntJbA0P8XVfwgl2B45yUCDW6qmFNawJXXz7gRi9wDHC4uFYf3
GX3kIl8voiYPzCWO2DS/GFC31/wvnRUH/UN8tJqEwslIZywg7OPxsRJSJT4pJs5vHuIW+Hj6AvhT
Hl113nvm5yRdaji5p1a9XDlz2Dp8oiqgVhRgMIjkRRbECIlaXDnlTGEkdi5Q+vvSZVpLtxTyu+8D
D80xIVGCmwp6iQwX+19/+prSU+gj7YkhVwVTboQxKR3BOGIJXOpZsetQUzfcD3G5+VePrmaq/MOK
V6ASk287vHPcBxmoBOsM89j53Vc4NWnlIYlh5RgHnR8743J2+w/74oPzdD76YZDOyd189GjN357b
1sD1huy9XKYZieuGgUl5qHtIQ4K/AhKsFV7/1k++xO6RdKqitkhnQAyAhc8+IhT27vvGzhNymtaD
oVqLxjq8xTqMQ1sQd6xU7o8VIAfzrWA16JcZ+FDx9oNmqSQfSn6K0IvaD9GKvOEyw6nesQJIOZKj
ANOS3/0kFtTpGRIPW+knWC8aeyzRcm/INz211zEY6HGahYZYZhYmZiTYBQnCwdrQuz+EsiEItM7G
8ilAWx9sxhFLB1N6Yv+4NrpYulxtnxIuKqfp8VqtIeIdsM++Ae/YQ/iFNXXE5ZbPznB1WJ9XzfmM
5AgzStWqSxLY907LWiMmLTltvy4HngFr7AuAc4WOJOp2pLhVG09gZYUnn3ovjTxRg746WNP8Wtlt
ByyFgdb5RUOrV8mcjQhLiBQNO3Hi27bWTdDDGW8kS+oxosejOKQh3IONq9WNltVFuGHKyo8DEoYe
vr7H3D7lGJXPMK+4ZN5h3JDKGi9eRTgkWW5OtCXfnftdCjlSRrzGbCIilV3myuBrlGe8q4dlscTa
iKFlfn1fvVcW0xqJ5Di5QLoIa3ANt3GjfOuKWMcjdmQ9/0PeFdDWk3KALMOvjNMB1xlDco3/2nmq
pM3GyYIOAifxbXp6NKSndIR5eNKygQ492xbzVcMWvdXL2H7Ey/n0wqFVAS36ocXLKBhksJBdahED
5b+N+hQpMZ5rzHYdB36cZUTPuhNliyHxKxaFtsipYfK8Vw2xluJ3KSCDfWaLSWQSpjY+nInLu8T3
9Ey1lcJ73quF51e0Ac7J0s+Vbur+cKnJuCynIvsT8ewZ04ishSBmdQ8BGBGi11xHorx7voqzQPMz
DL2OIcJt1pDNCU1gWsIV3tId+2qiROWYKS9vTSJoB1IiDPUIOjikRZ9tsFu199xvqLQ+nGkQ8DXq
mdn4c7bBcxGA6WSPs1IPFRna14t0V2SC+PCrACJWQXdDwCvrD+tWpINN2fNKugczGKrIF8jZ3WR1
NMq3qbmo1b3Atk/GJliUoNydmLM7f+1ay1hprO3FOZys28mUiRE8o38V141jMsSMEHwMQNj8e7JH
OdFxZ987oF9w9MQKRH91ftY7yEI/h3x7oNQdZ2m6fjlP6sDUAie+cgT2vfnDFy0MdURrClLi20fp
qr+dN4zy7qMSEMeQfZtvLHFW5FFkmASy/ZPmz6wrQDWzcLIo4FNU0G7BNt6Su32ljF2qEAw3mTZm
2dlskJEu2LnMnCFMBERkCyyTf99J9oQWVSvoBAKO/9YBqg33aciroS235VfgATJB/wnXauyidd9z
ebF2us/rYyfET/nBWKThhnLCDct5flg+H40LQixp/D55LPe8uVoeT6rt8iJVIv6aJpi8kgWSuWiH
qd0+XecYTrxIKCzLryp+3hcktZpYACYjy/xRdpCGXH8D/JHXU+JcbCUoDNxxJVZuQZGVUBu+Hi/A
NnjcgkEGju5wtio8axYKc5FxqPMH90/YaD7r1Mbu0h+wfHrH4FsWqjvpHDxA4LxdFOpOzzHw7jwY
0R8EfNjV83q4gb7DEBkUt9S8nkuGU7dBzEqx/UWgR6YPg6Ob3Ab6eolG1tBALcx2Ud2k5JvEl7hC
Q7Id6LNNzKunflP31vGoNGqfLwY8hsUtLVBJNVEaacHXGTcTcEnDWFq/T8NDMTDqq7UDuXYMik2z
xbDkboz+G+eHKlFJXZA0oEyXn8yNAbqFM8ZvJs9qFqJWfufNapW8muSZ6qk3E6AU3krduerxtx6e
Z+GM3xYv3yNnkaDsWNIQksYjIYoYEeJZcVhhGKFrN/zquFpsK97Z8e+sBoZW70/N7X7agOomZgKf
nLmjzVT3d/25XMa+DSh7roFrKCncX5AHOJsva5xTIrHAfNSg7j1M5XiGXAtsZjJJlpaF9jIeC79H
BC0hIKvYDyG/6xMngje5sSxvRk5+qQLu4A5sGbZB58c8K++Yewy/PAzT57A51ta6eC67gV8i1ZJX
un9sLfifl2tjNVYz/2bf8DNhMnZfKcSYtVfMyLRgcovG2eu3vvSFpjXph9CscHBodUWFjtWxZnYk
z6NvnK/MlZUJQwTAAEBULcfM9vi8kP98240IQ/6VET+5c6Su8k9AxHyB7Zb26mrZJr73P2X88W5b
2OXNWynR+Vbd+4UVkiURy/M92MbysIiXWpOj7SBFSfsTmWPjV49a2zeprJF9OY6FZ2+2c+eEYys5
ZGmTHkEF7ZlvWqYu5T/PoAPr39SKT/C83Apd5aMn4IeO9GrSlKmeL5lfw8hpcp0+/KCA9QWlSkba
NlLrdf9BJ4jt73GMdGB19Gxco/bJI7/ZfikGI7broJcnJbrxMO1/PYJrcfDczHHyjORnLWXnWSHI
twyiHEJKI1qAM0RHrEMePX15Cs25cWOt9m2RH3yvbh1f7mJUYujytAKbzwAitYDESDzkT6SuxI/d
jTO+EhOcmPe+lTr7QGnAj8f0DCDqbj4uEKsOikWd2VaN2jDuZ1ldwARp69Otox1ah3Y6m00mngYj
B+WxX19M3vwkQIsvx53i4rYSpyAsaXdwSZh+ncR4oCZjjxhXT1LxDICJvAIsIT26ZLTn2T7nJNdy
6YolEdY4ln7rKBVEKZINWB76raI8st3wt0bA9eX0Oqlv6eNJrQg56Gw98gLNDzONaucUCVIE3A8H
0oMmiRgZuUnFkddh5M32MbMvLfxzDJw61ngR8S6XScPNKjwkTXbdNSMJhU7CZJuieU2a0hCynGSl
FbJW3fmk46M1KS8GOtqGzvguJnDDJ5D/+QNaQGK7hzR0v87R3kxWtCf2UkvIWW4r5dPx2pwZnTlh
Io2xVXBO+rUvadCDEeHRhmcCE6BYfSiLZjQW4/ZNjXY1pLTs0UZtVAz4DU3OSdoW8b0j5Cb8vKWv
BOCRij1ibCfyE5aCRztFhVvO0GQ9qS4YcCidDqYN21z2a0GyHP47irrdPDKyhKk/c9tw0bqD75ng
2QtedChO0MvZaMfv+82uGgvUPpTXAudjibv2DDMVoFwNaIoFZCwmAWKCCiTMAvcoB+JSgchd+qr5
tk3NcyTMr1ehoMPVPsOqsIFoB35T4nwQBt58Ss33hgkQvS0oNqPiKgRs4UNyl/Gcfp/hbBZatUZn
J1emV78aLUyT8S4+M/sgt0Wh6cp2wPObhkkoQb0Ro2Z0HGaZrZUzv60ZzDgw8d6cZHsyt5Kooa0q
/boxyqoHSb+6tPyBQ0SiRfAExUh1QH3nUI6/GXkgwiqyjTzZDv/mXEdL4DPE1KWJLdjoYaizdcJm
m4oPd+Pyl6zr531WwCpLH3eQMo0zNU0iiT3UaUSvkhG7wDhs/xQzkubC4xofI6BqOkZUkiJx2Ju/
4zD46t3h0WH3nNqsoBSD38CMTDCOnW6W3D4hG7OzHoiTPvCWvIY+0/rYLV/Ma8ZsZmhTQCcwNgbI
Lm6NaXnPEaka5N5T0n0yxjbYh2PMftKalz4MxujceNVcFF5V+5RnyWPpzD3a9aYv5EX7u61ze48b
scslj43FChCRDCiHPYTCnnt0IIlTSmxyBjpMQkPbgAF0kOjDrg/O4oequRmlFF7v+TyzWFy8RTIL
oSszpN2ehMm9lqb1mqissZRE8pskZAnMvx/YS5xafKLE4mTiRpYy78oDJPGO9YOIyphDP+WzQbur
Rjk5VM7KHrGvISxvJwulezIummEdOORUGzwWAC2Cgg5xwxLY5UjdXWSPp/bIpJdGspX9aiTzipcy
6TG5H+Zm78xelOPr/fJZj52bmQRdekKe0rzEbUMK2utFeJyKWkIFohQdXVV8T6uF26Fix89i2KrH
JQtsWGNgcYFygFFugEaDydLOcDLd/g5Q5zzgD8l6uo1JVbx8B1Z/vHAjxfkXlqC6anffaN6l3qyX
5z/W8aQUa0rQgDoLuJj1p/t/oA0sbfJL+JGzYzD+FSVpj4umVQ/XYG3Llemsigbeyt7a9HQBxUqI
eDZLt3CRcTiqRK4Ii0Em6xfWvzdM1sPCyG8dN/PKh9dY0beF8cRN06xTaOdQPf3Qv7PmN5MAEBYh
GMNBm9FLslvui7vhN33tdQWStvCgXstfkTVhMuQDEJn9inCIWOS8X+uQ/DOixoKxxMzS9KhXCW2t
RH1iBoaYE+WoxQwRok6x72RoWcrD9aLoZ+p3kb3bUL/W21Y+12WQ9k1S5lwF7OgTzmHd/YaOESCH
Dvsy9o9eFaBmqHD1mt6Nc3tPFf+ygrtEhmOkBlmltcMjrjPsYE3U5KmBm4/ZSPKvApTL93djNJ2g
/VinEBosxEI/1uvfM2RoU98IL8b+mpPmyIZ758YCn7szpZ1zkFSEm8qXfRifRHufAWfvahh9oGNX
yuwzlzinbQEBr6gBmWIT95Uj35elz03XhHEVw16z+YPeqOB8SOAhZ+vVH99LvXEVy1Wimk2N6t2c
XlcC5fPV+MADyhrYp72iPjLwKd90IC1tGSjAb6QcT7FWMUrxMxzBlk3O5U+QQtWjgdA9wPSZE99B
eydTV/OVRrwH5CJYf3Z9fRoulppSBXo62e8msFY/0pD9es7BdvYPRU4KWWFwWuAxkp/vDLdaZceC
zEBNdhfggMdOXZcNwgPinVf706soxCjQv0glU0+R+9QziQ2jEd4DEDAVvn0iiVrP5DpjJ7/fSXPj
YbIuEBl30SuhW8mqZKSK3b7bbJswBeH+lTrraimzEJ5IG+7P+RJ7ZzAKL0zh4CVEW6rbSPKTu78y
OsM5JRnisREdAy/ie9RdCNoRNVnw6ei/Hsf2z+QN3y9iopR+Pt7cTmE/mQV7p79c62IbDOSIPtVq
q5HDEo+xAal5KkAYqPhs9e7f69w4caZmpJkVWmNJ7jprPbNlIhfSw/AQP0UiZQf1Em3zxyPUxmox
TbVPm7TJO9HWCGxDMcSY/A1XRK56uYl8vZk1LGGa8MGw7dlj5tutRF2XqWRBiH7KpL8y14g1bm1D
jJbZ+AAFzsTUP3yXYJzmdz3N+3w/R7q1T1sBktl9P4XmwXrGBclHGH4qoRljB9pq1hdmrUXW8ozQ
6oDwLIg6PF7folddkT849nT1rMZU2pO8OnBUkQYhMgCCkhjk50fn4amQDnM42cXewhhd/T/XrwWl
3+ojrTBvfDYvz4CUBio3bj40j16GKEWM7FXfSPTFFMdakV5YahVi7MQKttM/75YdlkXmR/YaEFhA
BR0Vdpz4GykYgbBAC7xrVd09zeWL0e1PtKpM8T2Oa5JGCoea2/DOlUw61V1/AtXfMWqnkUXssWfF
RQHySlhzrgYpnXAwfVg9VfVhwqfQz7YdiWLy30VMVfBrf74IUlhISutgWNWkryvofRkmFHTI5xlN
u1ec0BcQxl2PoIonAxe2Yx1tcZjhvCnF99oxM0N8f1Q9EwCNeuckjMVUgOBMAQVbWKBcmMjJcmQb
QwN5Rnz7ZyXzLB+iclKiEII9mRlKKpAnPYs+RZD8ui/HTDP0eyjWWtLVM9fC6gJKb2WI/I26DB99
Xkyg+nuf0+otp+vOfIrXUmLNRCslfkV2oySMl9hGpb8XA246RhLytbVjvWNfq1Wz7hmnZKpUWDQv
/xkLBuO2v7sYOSwdk0/qGQ4lHdww0DCZ1XysoXLnLXAX3s+KVBfkxjENB66uj1KkLX72ItkMuzRQ
bfKsq5iJTCNlKD6/oevx60Eh9gWYggXZ0BAkfuq5JbTr2dWiEtXAwN1BqTH9gGlO73SiruzRj1A5
/l7fzt9xAlKF+jzGYhuGiLWzVuzYO1mFUlaaJ2KUBpCsnp999ZS/krKuwAxZ2/TKJlXE+DiKefWk
DKOoc6HbIqE5ZlMoVL2jNRQqJQxTi+LMddBbRjJpmSQ90wdBpnNuXyU0/Pg3OhQba+dCfSUzTJH+
MnEXnkLK15AfE0gYjGUwnmwpB/748/3DrTgu2VERBMWGD2DnG8zUvtL1MWjQ7wSzfgTN2Z5ZQlqs
6I16+TRTvBVz8V7j2zqINAU8eO44NKb3MixXXRFdBk5ICjjL+v22J4MlJcVh1InRG6lHPo8yXUA0
YPSsjkz3J6ZKAQNJ1tgg8+OnEWUHsz6NAtBgM2NBCX9eZIFTOb/SCl/x/9jLw+OFLRinpEDNGLYc
mJXq3U04NTWPHhQGVyF4q55Qxml2z1PA3SuwSLZ0KAf/fu5sgg2ysi1dmpXp7fC8YrpOg6tVbwKI
OvVEW443p9LzIk4Yu7o8an8RdyKnqZo2RxeKTWz7B/fc/zEhRJnrHYl0cWbUXvybu60JX4oPteeg
waNW8rrYx2YjlsjA06UVi3moNYMNu/iNphRxzizlA/L8Hvl6mvwbcb2CI8x6SSPxEx1dIw5gCxP2
9WL74A6F11e93/vK60/7/czbj95JA2hBl7jr6iil1TdsrEktOT8E0kGbV0hCNM6/4cej1eL7Mx8Q
khJFCV25PjAo/pTQ6rJQm1kkhcVAnKU+RHpwX6YdG1XJ6nxeZgTrum7clGx7/Q4zvE5dQzYmFiDo
dA15uH2nlKGgtnKqKgUL8TLrpnpquKO+UKE2zIOp8wiZv9hbM+vi3n2SFdPfJ/AI3U5WjuJ6ory8
H4vR1sAtyibSInXc6ZBtWqJ4IqRqAiuM7BRkhR3HjHjhG+Eo0CpVyjoDb2Goo5Gufs9yGTVKvntv
SzFTF4T5teJVesr5ZLkSHsS9q3zEbB3ozKz32lshfEWsqHoBHfZa5nHrGxjz5UYHMY1capMYkOOt
eAVzF3ZZWgJ8yBnMj6MvFnjH6nokVofixAFxCJSa+8bLp7kucSl1m6UMfWQvGN24n0flzGDqVqj/
UPs0CsZeUXu0gUAhPFDuHRbtQSXtrLEyACNTIXaHPtPu19/PJMN+3zRBzVvuLHES6+rlw4UialQk
z2cFsAPAwHhoBmKNpQp2QZ1dDR+9VsSk9p+0eIEEbsj2Wb0+ANwqb5a0yYvXurGSNBrCvjDh7iDa
mlSNm4t5DJlZTvu2uecBxaCka/Ne/Bifnm3yY02pZzelCJFqpvc4UabD1UjgRyJD0o4VqoA19c08
NQUEnHFz7af/mYAtdHo9u/NKdeHmRL5KfXzcI78VGjMN66QUzuO1pbl+dj+zx8H97nTvRIUER0A3
19v09IbfSWIKd2aMeTbrVgG28yyD9RyKaT/DJJBZGI7InzKtoZA/NG1EjrEYRSpni3ktDOVZNCcF
iq2XXYkr8OVVO25xbdwiWaLG4QW+0hy0YhrbTnt2s9Y7iV2dQLwAoBwTizKGDjDVhfAxbDRQcjYr
WgNHT8cmdnCSMeJ6ohTrIQ2+zJT9R5ZCeFV7pLSPXI+OmpqCajp5ZNPrlYClNgQYdTZ+NDMJJbaO
VmcuuKEqtmvHkxBAZhZSDHULH+So7eMjwF9C/2a9K9PPxPk8wAfhisZtagAYw2hIhIC28UnA/tJq
tZ6Bll2Ua2IQBhlt5pnmEQzprqWZKUc4r5HN+xxCyEe7BX5cEAcDxltRakrY8oKAZDSjYNypUVHs
7yj5r5cxKF68RXrzcWLPeOGOUu3UDQg4EutGp9t7Jpf+ISwWMQ3ANClBT/c5MVmYreByr5lTieid
vJrWopSPm7JnJ6SMQv2u6sTYTITLLk6j3chu2J7k4Mv0naseJ+WHQNrolTdqXCjEebtWEXzgbS8N
rktuNYTCpVqSMxUQJ3AjyGNt3pMTLJjVpcn0ogXeuRJoojta5ttDSfdQ4t3IXTsBb1HOaqMf67gM
EHRqQfGvBMo7M39jkt1vNNk4W9i2SUdj/1siv3FBI6wejN89RMgGrcTiZxlv9Jvgg9KE2xFkD4yM
QXqgUL6CD3c6fNstvSUSPPfm4R7S2Iax8wfnP4qb/W5tmg5v0tmLgahTUFTIuNXTlzDXk93uUWRa
//dD5RJzAYVMlRomo/LPd51HFhAxb/CSy5KQOTpZbPwJH1yW/ShE/OMl2nVEJ9JPavOVxFoviC1s
rVLeBieeSkhUuMTjqgUSUaYAaQIFhhX/X1IV4dUjAXG0j6n661Fq/HJbuqDWKcaC+gBXdWSwQ2RN
VwERviB4SHhz4OVG/nzlmeNIuSU0rV7RybSQEk5FKyubNNGUn2fF2xUw+kVInpIjXEXqFXsD1YWH
5JXfSAq+o1b5bZ+C752LiDlErE8Ce3Qz7NbDZwDA+eDfyVz+gfXPl1yoEJVFO6My4hEmJgdCh7iY
mFhVUPyEY0x4xnkoD+us1/Dc0Uskt/+TVbL9MM9ubSOfz4LpBSyVXCkAlXZhWUidZ4KzttEDH9OU
6cFCRYEFCQu4ybgWlpnzGHRF0RZurxfLDTfGKIwL71jVGCNPbmBp+0uD8fVNCkNms0VO/fYug5OK
O6ig3xZL8pony4dHTo9t5YQ2c6g8/ZK5v5bZtzR8mJ+5VDBfO/r7NX2GaPyv7BoDDaAaf8CstpaU
dgfZu5frFh/CPViB0fgEyS/RiPMueRQNeKbPfZRyNKzkPh14yYUSfqNV6ojhLvopdAQGguIN5o5S
Yz4BhQTlnThM/lK8Y2eScwASDRaxNBQrRJUR/0UYDnvR+moPDsC2lwv8DhxwoGx6LNJLxXAxPmku
WIaoeynisQctpyNEq/+g7irTuHgGIYGzFo3xz2GsM9vvXtq4FPgsmh7YGM12a2S2I3iMVRC8J3Ni
nDjVQLsS33UpmShMulFx1Gex77MaQH1RsObJH6CfYSUMQHyiXbRJjqXADc+ZLn5XdZjvfx3mW1Wu
8TVFyc4mkWbFRzRRJlmpRjlloSvK3hndTkjzCO0cH5LMfRXqozGX5DgiP5U8Vr7uZsJrE+Zx7DPT
NbjZn85XZhIqr7yECIfu9c5318oLMBHtKvkHpC5vdvTupb/VxwsciBwwqO9DBRNLSV/LbK9tTUrp
jbPnI9WoIEX67dLAVJFHV/lkEY1zGnxnPZU+FPEEgwoytI86qkiomtGCQgM7+jcuTB4SH8hBXqci
xx1eSdbZ8iz8HBwfId8oqEKmNiHkoUlyGwCvql49S7RqtGE2lnJtEPqecJzfwTefQa/MtatL+eOV
PmMNwcYvReZ+jh287zCA8zpzXaaGmShH+tepenDg+IE9nSDnjvttcVUdpiSRMQOxRmMvo5ewINzJ
rewRG8Im0tkJlYmPIgaHK4NQZSW1WHO/Rw1WcrS4rw4Pnj4Q3iPOh9B7HejmwrVukiKl0sUIL1fd
RILddLpHDxDcsConmLH1xDRYkyb71yhxNVVDXK7Iy/em8UeXm9Qd7M7c5I3uCpUi5ujixdgurVtT
ghLJZhu3taXiF8ckW7M0FW/Dp7+savAEbTGwf3Suga6OQXltwMkTKXx6kxXWN/Zi3NR8dt+FQD1I
twDEmknK71wSYKgvxVGl+AXno7c40HwVFuC05/OXl55Rj3xM1BsX2EbH++MmGiMREZwgxuTq6eIC
aLIaDoqYSmpqTvmcLOB4Qpxx+4oRvuqflTfxIVBEgVZq1BFFfHHWw8hkszIxvA8MfKllntj5TWSG
afF1uHagybnYAesiOOigaxRIkfgBxBJg4/UJ6Tc5j1Gx/rrs2Zi55kvkrtx+ebuioMrlL510OTSx
SfRsSDd9uMqTuCordq88+/PPduG5/7pSQdRHFysECrstBpbJbCvjWTRInkFHuhhaF5ufi53HMpQD
iZo8YUkmfscliKz44TEWbZTWwqBDdMqJjRMttFyHkrnchyQLwHE/QbFzuLLMHIU/3edi9UuRqcXa
fzczb6YU5bbKWKDeb8gPb/7syqE3UkMbwiJq+uBywMmNCb0hI1uYI2DCeynz3dZyQav6vJkwER+6
MgPeUKh31mzhgBSxB5XzD5YSgYYkN2LUoBBirH4uuQM7ApgTImvJo7fV3dyLT3ZMrHcJwY5FUOzG
nZ02+JAGdhymFbwSA3VjefMq0hhnyYP4aWUe/9Q4htkRSwr5wEm9QeuOMNq6enTHMbe5nyvXKoLn
ZP8RwAAWsZn5u3kL9zAyszqrXfeVPcDTVciPMmLV5duBkjjqe8nvK2c3/hJo/iB0dye1v/vhhro8
4InTpPZbf6EPa2e1RXrwYACFynDSlEIJUAySNqr3YGoGF2sXee/CVFhYv3SZrqr+hstLDWXJ2cD9
dOZy9Vh0ZRVqMVDAHabj0ZCG4IvUVKv7v1sXIbsomBy8gBtf7Jbg5WJac7Kj1anzefccZFeteZK5
6uTPCtMCwfiq0/t3e+W9XdWXPqSS9LRcdA7iWVpsTSGHpLt8lrTlqsze3CYlo9GsOdR5SxlqribT
qGoCnkDb8wne1kQDUSQI8g3iBLtBMYWIeg4l/biVx6UOAJ+CP8JGZSDQLku2e4L5KXAhczve0ZmY
1qn0Pc2rnv2mRZwacJZT2uikZ4RxDNOjn5o74NvxPIMJpvDVUazM4pFecC9+1n9DWAZFtMSMNCdE
xmqfcoxZ9aSGit38/lMaRCrkClE5yu7R4FgxpLvk7N4ooRSQc59/IcdAMR9SBLgxiD9erkpYiUTL
ynFmlFlNTTKRutKVnuOOra6dcm2VEfmpFkG/cSE5TzaqdTCzYXebAf6C7hycslcZrUeNs99NBeHj
O25ivzupFY2ruiVGghtJhwJbI/bOEDstcIg+lWdh5Ti65Hi7rMZnH7wq3Kx3ouMByP30UzbIkiJ9
OX2k/uQDM/195iCg7YuaPAeSCLFOol+MDpyFLB8Tj0H2XIhH7xNzn3IwTXo7VjMVZK2TH6wp/ZaM
ebLKkFn2kcDIq1beovAgwd7riEMZzJ2OdfIyIMb7ZiABeMHxEhBdMggNxlLmuJxdv+Y7rKBwe2K4
6+86c0zAUpwiPz33noo2Z27TcFDWRGqywyIgNoeYnAEdi+dGb1iR247DXZGl6ZQqCzWJGNciiHfc
tl58bAMhbtGp73W25xrY8wzdQ3d0EYbdpVxvUqsiSGivollnm8bCNV+Yd/3s7OAW6KnrMD7YfxYj
IJ56/jmG/xTEJjKORmnNIwseKpFhH4QHBV5TFJoCoXbCYddn6LC9rfIIuWUi/BDHb0OyyHMyia8e
rOB7D0NhhbB1MQAyTKtG6sutlA167M06gmdKxu6AO46cwl0Vz7jKOB9vDp6JZ3eI1ay+0lGIXhvw
Hzyho2xKPjSL3Ui23n6ReOmeKmaYVY5anJGZ+zVZELfcCERTSeHNQ0bHUZSy5iEZ6C90rqlR2oPo
nVxG+uCTNJ/gXbPgRTIEkJhHpDDC1UIBwUvyTbY0Gf4zClkaGDvwP+N1RePiMoTyuWetD1e0Taix
linMhA/cj4q15HeXCvmciW85qqKiqizzw2YUmMSiFkUnDmtORiUoxgz5SiaFdHvcB7pVsPMrgLN9
p3Q6ouF5mpywvvYqJESpe/Zd8fQoqtSxvUisx7/hv4/JaWVtZtULqAjcaD2+jFO36Eh2R9S7cqfc
SpDQo+I3ao7zIK4MKdSOwBXBua6Uaazj11hTz1A38xI+2bwbcu1MBckM28n4hpFowZfOfrU8on6k
qclixfw7FpSGWbgM9lttIzVFqnYuhikh+HwfVlnhTaqDg9wTH2G9PnJQj1sgmyrZwRnZ73D+gfBz
iKJbcpNCjpfm+Qibnu3igklX72vscxaNPVKVprCyHGe5nX+EYlH644FFU0pcYEpPDYNVB12b8D3/
zx72T0zZIGpibniCc2a3YQzvKaROkjZNFGQ1lGeU9QWa/W6cU+YxY03Bsla/3Q8Z6MaNoKPTBPWz
FYvOlRfYCc1U97si6YuYpd0vbipfVlmo4uLKw50Fog3QDuGyvF6VKs8g/lX/OKIVbKZOtK56DQsH
CcZnSEABqpkuiNVPelBXykVKN1FbSCrLiYMS7bgGJ7wNkWkwIHC87ONbh1r7JdVKrnvo2QlxaZNz
ArxryxM/LXuWwy5zkE4rOeJ+AyXsbWoqw2k2aQcRiWc83aEobMqLsLAB+LUi8vMwNN0kBd0wMtqj
QdY61XEdJLymk4apOb/aBfqCaSM+b5Z/AH3ir8tJDyCf4aGP2IEMWY0rO45XRohmPiWPEQNKa8mq
bXWTx7D2Hjtd2ZvJOGXO9dBt45RPJ0VhkKieHw8ahvBNy3ctrkmke5KEiT1VVZCZj+MJzt6Fm7Mn
x8BETTLY2yk1Iylg6G2q8r9kxzBYQeQnfcRUL7YPnxfTjavTpiDdmuiU9lvzCfyCCSYz/Jw9mdxV
jkbTr1Rwdf9HXkig5kHKQsKiQ5UYKRkg/dYC4VJ5kIdP5xZArYqfeA+k5zz8lAi2Ola+K0+RWD8r
5Deu0ewJfEwvnTaHoyTHV4Dx9LxcMCYlvGUKxTyFgCeVa0QYuabeb49k7Ql8BBPtGbz0KQ0yZ8dR
UX6v1WJQduxp912sFEF1JLic9ZNKbHE6ydzYCa4O6GAadfqdXgU5D0mR+9gvTH5K6qeLg/9ufz1F
G3EeuTMO3eFrYYgqELeoWujYbFY625/juOt0YsmqJTE15ejhKW9I7Y+C+nxRu2vcsdKifiopL4IX
hZY8N3zIErrcoxppPnnLLI4RlD4gIwGi4XjXaI+pjCm5lcpdij7jAeqRy8+XW85XehDJk+xv6pxD
AycmIn29XltNjvTqSLtWkbSxbHZxtU2EnoBvtJLUcV2WWf8DUJXVJASLtVTYOsiHaAZ3e2IKYsNr
JiCfYnTb3ATmCtgpZ8w0eLae6FN4+F1ilEbtbN1BBWtRAi4Punx6wC7CMpI+a053usgIA4tMHnZQ
Eglix0p0AJR6mlSukA1w5CkXwC7/L4LLKf0bpdDgxTkI9jqXR8yMw/4MMr9tVzP9UfhKabLGMWrn
vvwT2fzZrgB0OGTZV0muVDOHcB3+KS4qJo9H7YziMCMtOzCNeRu8IqszPBZKsSGL6cwxhIh4zKit
fQ8oQduUuM73mLEXjGbusp9QwXtLBkvcLITRb5XeZhyoRovS7XjW5nMZPOFtNgbdRkoYMHOCB9r9
+uK3/eW9Cswg8fM42J0pe1Sf1HlkIuomr9CXn7spXwlJucdswe3y46Zo/vCpW2eg9PeuELaiUyAa
WiiTw+fs5tbNgQrWYWWaEl4RZmnd9+op7PFTq6Ab+s9sQmld/KdfO6O8qfb9KcmP+RCXq8/+Tz9I
IO4S03d8xeYwetJO6X8FoWWk6Agk/S3oETh6EnWqmY8LcllPS31eLWIjYOXgljZ1MBoVpOWbuIJm
qdxO5MM5Pr3lZxRotHMqZHDmHbtq2ViKmDTP+ME8761tznAD4Hz/K5aXwvTJ3Iih50MZgrsvNxGA
lfkfWm+pmqOhSnJXZ3LNbapNDt8AEaWJHUNZbd04YBTuYKK1pEMKC2xDPawG8RAWdNFIW5/rygsY
3V5hKH1xCiog+J/onsx4mZrFnPuQ4UBq8ync5+SzFNIzS+Xz7NDIKCCG4wqaUmn0Gymq/j+w+lLA
zvyKWc+wR/qMYBQMcR7VLA4c9aljGXubtZBOd5rVpYE2KBFr+khonPT6rvCU9iFB0EPro62MUenU
Cs6Cn18MWC/knA0sg49ONo4zDYdJbWwGtKNk6X14CSXRe0wXo2iV7x+MXzUOI6+OMrdJG7EfnRh+
5R6HRxXRza87s95SDmbONtnIVhfrK4zdVPUbLvEDWKBAnXDpmeBqM1HF9CGSwZlt8zKTTpyQtmeu
eLCEsL+5YzBLH8U/ToO7AuHZKd1QiZo8PVIQt7y7IzNAkvCK66rH7PfsmOzO6CCLfaz7ApZNRy57
qxY0uBFNmx9smxTzUcLXHQl0A0SqFMNqZ0a1o0CHRCX1mPDJUEoXsfrRzRF7AWgvxfYl3xyyPWHB
TNxiF75OZPLXnUDCO0uEbjxfTB26cWEylMXkDxfHfAXX/DKb/8YfGRfHFAyb+J+hqDTDJNEjk6IU
oUMT/V/fVQPTeHC+YGcUzIHFH8tGxjZXQzk60MH8oHz1PB5Y4FHR9vfeAIa73CS3XeRfr5x9YLpe
sH7YhV81dQ+0LtX1GGVWF9lMpGzNtk1IMVbIcmvPrg0xCEg9UUhUFfSh3AOUTimBdKp4vtESniKC
cw8g6MdbcrDSpOSpdO0ZjjjQmuTpNDW3H5GBAdiVmFv+ouKqXoQ+9xM4v8mA41ABc7ZaanjVJFT9
XdgR/1nbJcJGbG+FwjPl6N8Ooljqzh1StYubDXAKV5BTxudQYUuvLB0NFaovkOYZWdfq8wTnsHj5
jJs+JI4a5sRYiRzQUmEJfxWLgGsT6TYMrcNUE+dRskorCwdHa1200CDOVnc60VCYVf6aSoYpl2Ul
pjVrsMitxnzJg+At4GCQt7cBSO6P5YLhBAAVCYWUbxA+goCe4EpHNi7evhtKUCcaiwqa1pjNXb1Q
yqm6E5z4YLkn9Ux214Bkr7E4cSA8Sohy1JqAEkgVVX/MD+7k1CncDsZR+o6KYVGz44Xw4VQfsjdf
0GUJrmmnDk6gPtLwTc5p/eBVbagYNWwWVdupw4WxYLNPF6uVy40ClMfvbATucawlZIwHNGsHb2WU
zNHtBwAg5bXpP8OQOLCEKtc9vrWu3RmuwYrqNv5BVsfw6dWzvIXso4Hvk3gVZrAyvtB0GgfEft6J
Bb293zimIHc8UwQWM8lTcmDrQgmo8/iNr04NDhFNG9bZ3/hfTK/tOY0ClX13msZT4vIVO6CcHsFD
lfhrd3aguBUk6h6GZSiMM3EvPB+cPotjZ/bM2xsqkfKF7QixCJ7w4tOP/Ns3vkfsb7Kd6X931xIZ
M/lXph8iySk7A2qX+M3MgQ6EXIaWpQqkd/dup6BtmGPoVcV5qFo1gv6BFOrc4auibQ1fuwSsVuy8
E7qw0TS7l7khfF5rlyM/aRYhglRxAxw+tGEWMjdEBdJniN0aFawWi+wVjyMuTQvz+zBMwznTbrHr
64u3TgvQ1dpvN4mXz0qeE8ArtL0dwbqnNC+TRONGYEj0caSH4NOgN42UK273hSfs90/+5aRvUjCS
agkd+3zPwS7QwVpTyeU6ZdkEkmVv9g50uFU/4kW85tTQQhqiKdSI7LBm6GlAQmzNx5ksjRt8nJYE
8IP+fG+O45HScRVbYx9QPIt9dcWaZoW2Vq/0Cf8Zfqj+1KU4LC1PZkUpqy95LI6p8dJ35PNWmoqJ
yY4HKHLLgtjzyErTjiszwmnyCzNvjn59TXSnqAK2I/h/0pmyTH2HzDzlN9F0gpGeun1gsLxcqF8b
KMNm55hFOfUoQznvsO9d9IrFd807YFtYy8cVJeE05yrV9Mqg4dbA8anXCYFDuqYto6kh7lrYYn+L
VYOho7du82iBkql0eLvv88pUsiAjdgA7hbGMV3RQQj4bJXH7KkrkW/gxYyY02tVu/LOQpGdHdWbq
Giyq8s8bJnOwavzEJ0Yb2KSXQ9TB78o5vYLN5OTOzOFjgfv0aOfsp0Z3D8YhLOYCx524GRVFQjLp
w+3fKeg+YzZitLZlptFRaoDAIvdmQNg61FS5Yo/43falj93Ir4qM2gqJQv59CJjvNk1OmUuE10wt
QmFfvB1l0/JQr8u5AeaWgSXmPY0TDNVXMStF7KynTGq+hAoJjFe2RkhRHszRbe43gY4a3S99JMb3
yDLo341RAPsJtwY4RWaailAQWLBZvoidc5yRDjQOhAd1oQh9sAeEzMV1nlaPnBMRupnjr+3bZDth
e4WlvFQ+CW1FUCMyn3KTjnKaiJ+DiMQQSJMr/ejIbJqwsbEJwcdstTvJLefJcPsJanBrKgYdVtBZ
EfF3NGTsGwRNCjP4Mtr/thHX+Qak8C9VTI/3eu8mPg/hca5dQsqvE7RlqVu7LdD4qDBhewsW16Ul
h6EsZnPz30yqU3aJwdMkMeO98WxKURJkt45OvfJJpFr13e681RhFlYiDoihoVFdEZEIJHCasaPkd
jPp28PKPGufA1QklVwRXAL2Lj6Ttf5DAlo6Cr5546M5HS1090jjFkt3OjUB/1HrxdLNk+y4ggUjz
9a4jmOuNfqMHWbsqdh+fJJuzjhDzs7kxr3DR5j2O+PTRmZzqN0Rb6PVTu3adVwgcaoImoXn0VilE
KJZFyrIJaXDGzFg6Gof4SdN8iZpxCludAPp4HXbRXw6b6YggngiaAGWAYJJFvjfM6MwwQ0NL8GuI
hYHBoil4RyqaYRphgTB2wc75Igb9/2OoRcguWIjTR6YN/JQCIs4ytQGPeCRh3UN4iK7X0xMr6Ljr
xHeJErznzA8YllHwNlOFTzzBs5wWVjDoK3/5FH173MEyS3K5lSWEIGlEYKiZMUHY+6B4b7A2rGGr
QafgefKqgQ4v1SNljK5Sih765tSvU9KalLAP1Do4iOnElbqiSy7iS7MoPPhWqqubaD2YMdPJm8sW
gJHGFHnXnHrjo4EPjtQ9RE44yc2zEiR01ROMjzTqZl4n8SyRxeW+0VpDnupfwSoyiCpbJtUdjSty
xbw0/iMU9iGH9QzNPHr1L57n3LJAFWxgxn7DMNOkz5yZD18OZnfhisiAIcnSFM1UXnIxXMffC23A
JX+VWpEMrRrNN50afbKM2TzmhLBaMRmtaSvgLI6jUiLkr/nXdBxPwTLk27Q0zkoKlR/RK31UaYLl
5Ag39S6KQiA+3DodmfgjMqVCdKLAEHTy/nBlrTzviv4Wrl0WFlHHfLWh5vOdeG+5q0qP1w0sfZkp
cZhbiWvLcYlPDbaEhpmA1x5LqBPzxyocg/DJxT8TBaegH7kviXQeVAPuE7xyrm1mwOufSyOQIdY7
n0zqwWioXck1t6OPQNLNLzmPoYkTFrv9KxX+vEF+ZBdTmoHAymaY9iSxQMloeNo51WbjZ5Xwd1jq
V55GATIbmCnAugDBwHPJyDKxaHHUEoDtjvHC1PlRh4P0fzcEjOLBNSQ6MAkr4ye7mDR171W+hCR2
I6RXGzKvuAisj74J5rHwJnU7qZXyLJaaQLXQ0cPKkmc5Ncgp15GXNzBu26jnFweYBP7OUT5UJhHP
y2FcahQW1Xt3NffpaXwC8+7tbTNKhDsycMs9GvgjjF/eQ8QRXhFYKhMyYoAe0PVCKMS3rf0Rhw2i
eLKxSajAhXo95yGmrkprLmKhNBefg+EcGR+4dAv99qBiq3ZuRa0F/asBsdbl+R9jPYtH0QQtv43t
m/63QT5J1IFWPZv2YynJSCThB+HfcpItvb5wvef4hwGtrmvb+QXVri0+0Qr9FrrVTJ1Xsgm+soK2
/E7mem1Yu6XGRSimGG8VVQRWtwifo8NCuClv3KYl09d+v+mgRYx5xmD7I11JiOCPtYt5u5QNd2Oy
2DCrhwv2PVJJzi6ijtFW5mE1T7tSVr95/cOp0/A4PtFlyg4Tn3pXgJFUgXOb2kUQ752KO0Vz1s1T
CXxyfEX6BiVvKA+lQeGq+0ZeeZeUT0w9SvaiM3fcBBouv4FvzrnCLrEV/lgSZkLHE5fLUBw1SfqD
+spEcG0Qey1rI8ZmKpmVgJYchCReAHlV+HKv4Cb/if+yyytA0IPUq4vAcCCSTTCxemG1eOeCqhED
95I8eSmnRyAJG16OF14IVhbbKK3oSkDcaaPpHtrupN18eVFX7m2gzTSE7A/VpTx1dwyPR/tMRDCn
DyoBm4ZG6y8+cI6FbA543531wzKn8zCX7bHBfEsOLng1R/Z4K71SGQkifc9WB5qel1VLGcZ0KhaX
RtIByUAB4RGcAxpFw40Du/X8mO+MCkE/GeqENvp/oVJrqSexqnsIO8rKCbbzdLZYURRhQf+wuBHw
yH+SEF8+nWq5AOs93I7FbCab+yWKWNKbOfRjv8kEok4AEsCDug33l7NDj7YlFcGEcsTpuCxyAkVb
2+k6PbG9QE4MnRkjJ6RJgGZg+QOGxJYxBc7bVS/smj+q/tgKsavcg9ve0FtXbwqacK40qe8qbi3H
/3jvdkKPBOpIHlzqlCaW9KDhLcVtDtO9UFYjD3jKAOOmOdfERzldo3mhcJzr3WDovEzswvaJnubl
ze5FYjR/Hg06z8Vt+GBiNFkTVwiCqhc85TZ9e05apDxtzZ7ESP7xMWSAJ9SKRgjSeceOzvFiQryI
KLgbFNLXlwF4MAEN1KsdVDeqGjdjpb9Pwj8DCNMv50zHfv+dbhqkeRwsq+f9orFKH+9cXqsfvNGI
iFyHcB7n7tMVpx0xHKbMiUIh5iA94q/t/HsdU9AufYIJ/yVdngq4JaRQP/YH3HjgLND5/iynsDzO
nyWz66PnHDZSqh0dDQjxC1Ok4sn29XL/8XBZoHLOnrVynMCOJCP3WZAXJk0trxou36CQ4FxT2LAD
J20RT3+11SA71SR8I9gHpFbsy9d3dhsA6fa9vLdNS4PykLaS+mmhsDETRnwqEmpLnvGxqftDjqCf
YPNFJs4dlF1ZIPqTj9/OxEjRzet4gho4gTBED6v3ADggFtv+BEhSNy+/xBv24QaV9+yehR4xNp3k
yEyDB7linsoaGCFRzltf+88dnpRdHkQWWyDDUuQsgpPJJTSsFRPxo6+jVDP2jXfH8TjDgJipZVqZ
fd8A9DZw41L9HQFLOPbu+weA6INB8lUe/AnSVi2/w6oQx7y/npLvX6F6JvKUtS8TlSWel7YLmfBE
LgzzJ5wUF3k7CpxI36oHdcVuZ8g1nrYqNq1KpdgRY8Ud8YuqfPPMMACZHzLYg6/5aq/sHznTV34c
LMFnVpMdO8E5TZ+hyp9oBYWnmwQnWGfsBLls2/p3RRVNkzDBRJsxAd4HROiQ9UV4tUUF5qjqL2HN
em9Ubp40oZ+CY9Yu20ovthkTr7Hl8Tuhi74Px3HXRtqavQk9T8D4J+aGpv1CAmJhTee3iyM5SSL9
lvdG22nrD7zcMFsw19Aep+5we1ABIrJ8CoEq3zvkkn/+tKnKe1lKUHpDiWFuw6zTVElMadCAfjL/
TGM6DJV5uUergi4BucZw3XISelUgeIMo4PyPwOHtAwOVaVop0Y9vavAVqjlr5twyk3Mu8BnrycpP
wo1NYTDNncttMQprBbdY5XAyrh/DCQWbdbQW2eTMQNijlMSyv1P0OqL9Szuw2/FJDyVB8mP9a4yY
lBq91ZO8RxpOjd0XXjJ+eo4pZbt8iA38qJpldf53PSmK5sT8S9cZgKMv5qsS3NDAtNaBdEdb/atq
hFMg48eFsa7mJmK3b98e81rgR7sIcIwmaD/QIAgxQW3y3qfccD1dvWqqJ9bd11Yzf9PEUDm7q2W7
MKo05wfGs2/+Xp67MJE6Rvx+TFaERW2n/2TselIkxaHrn1c0fT7WMk3bh/+uiQkQ3L4JrqomAbVh
ue+JCXmdP8UNXHTUBXaYO9S3FT7C96yyMl4hWxKW6ZjAlAfCtyhxrF/C4NKFniZJMrSiEHcfJjVN
GKagvMnGIQiB0kEXYx60Q327FoNwFeQSvYpR+aj0Bx3PdCluJDwWDw9tMxjvMersw8s7sNftO3kN
t7ZJp62Jc39evxMVbhLEJr6N4NgxdfGfHrL95LBtBb8jjF7Ns5FMP+sfnz56J0POem7C37auXlb4
53YNe6FH744mu0UYTpAiar+Muk2N4I01wDVNOfg4J4mkEoe7/qZnscfjy9Jp49gmNC/vfsNkzZ6o
Yj7QHUPF1b8M5wj1GfVckhFmyFumMx6A1qBuL9z8ZxQO9Wwe+VOvO214+1hXbct9irtJ3kSlPfjL
ehEI6yzP9E27ypFF/HT6jDkavk7XrdrR4vEs/4ofKaWeukiJT805hrMz+eIANYqUQMclYKVodDRZ
ysqoJL5vJPn69bTfBuOKsOcygQlem+PSEUthvc1KWvSfDZZjgrYl46s2vFXfq/KEsW41+SFgZGYU
kdOxWfYo5vTUHsYQlKvRSILk5bx/GHaNzgBwvTF4VhI37RLIHlWdjnGB53P82+ooEjI9JY6fHt23
4Glsdp0JkUaK2DdjEqlPYsaUBw8c611wO1ozQeuyZxas1g/+Tby+uI0P333npuRJy/bh+swtyR2c
IL04nMc3Q8MrlKc1QQo66cvtta25CI7vARNWQg1+G7T2K3xmCy3nrZkSw1HBlFzWt8ldc0yWeq8g
RnXWFjChLQeYYdGyC4fw2tArOI6JI3vjn7satDQ6lK+fBUT5i9wEZYsa1KY5pF+pQkuw1uVFzj1G
lSu4CvYZ0Cv1OyzS8eHNKtqjMnM/v8+4PEKvFy+NLKkXrSlFt43BWCuA9QdFrn1VNj4+aKZ9fcdw
WRKS4tNqi6PilzS8TFVAgmsLhG62AO24m2MBx1oV1qQjZqrYLLfpHIgvV8jUmqjS7bT/2pH6wGYl
lyvOhFFuXvW1m5RxuhdgMXGNigZmzDHYIoE/wt4K95pdmS1+i5uCJhQvwM05+u6dXGhqwl/wrcS5
k10tl3eSTGkBFLzwqeFWrMrKUXsN3RJl+ofSHnHkE4yIkhr995MPQpbOL3T00/GUdjvJWFSf016m
TQ6nj0h45MgvBZ/l5jnMpHvLprI0tJ/bhbEm6L97K3T6CScWz/122rrTNpCDu36LWLgYsFPmFizB
e9Vuc9TLAR7mCdbVwN2bqLtv9jh1oC90Jxx6iJa+Z1lwafrZIRmjzGcZL8us8my6mPg0n6WHspMD
Pc/qt7AQlE5HcCc4fJXwW9Agfv3mnG+DlRBaj3OEvegtPucaSVIs3R39EvhplmbhIBWS6kKmL38M
i5OU805/sKavZHfnnd6Xahl6K0oVka62OphYmqNgCPBGNfRbJrVpW3WhEPvkhc5++tmQDTNWOwBa
/CmO31r9Hv/qG6Lp6p5rkrkMxuX9/BBepIVU/0a5NMNSvXmEpesGU641Pz7nlCNNGHy0iEHugNYi
zRfVF/Qup8ze/wu8N4uhsrl6fBxqBHpFCvqLEQ2FHCh7CsPl4N8WCK9bSOqZkP63w00wFYJbJU5s
KbD7ogyvlvRbgbVtpYaq8r6N+ycpGribg4aUYXdFjybB/8EeE4dhbC8kfTXIvAaox57Dgp8ETbEP
rpsxG42quskDsDKynWOrmiN6X0b4ZQbPZ3aTw5sZwd4cu3qutGlIyB+4uT4u+XrdvwbB76GFies5
wkJjKwzZb5PUPR4SBQx0FWwirBUvb+OmDM/6wRemBymNE9oyBLf9hgS8UKxr1Fx9vagwroHf65gH
cBmTcRUG3ScQsp1ndAOYxCQa+4cCICBJGA8YS3h//6cXPMQPlV+PiE8bnTWsOe7DTcjqgpc2cp8h
Y4C7nA2tz4bBrdbDvC5e904sbN1uu5g8FMeSA1f14GhwDKWu6muEUBcV/U3tmSH9dzCH+A2DilOg
93qmVs4Z9t57TFNuaWT9UJ0SjezQN/+HWgTKApp0oZikpNLC7HsnPh70kAgytwj7E4vhoz2wdUmV
tg1P4TL1/CXkCMJJS4SfFaZRJj9jIwSSLQQPSMU9mXeem7DnhDWeD34O0HroDqt1Qt+tgIkaw/BU
3uSlhP+MMKYikojgMgH2f7aWwHvkhHoAaD+CYU+dJ29KfZv4oxek26Z/2SwEzkpluovxd2o42Ny3
DKNb+Ujqsjl6T4AThcSScuCt2UExtiA+EOo05O4mJ/cnUEi/rw2TJAZT5C7Kj8OlAtjBDB6Dn6zD
zl3r+yuXMzFMsy5O3t/Ly4MKmLy45nlBMzVSFGdtKxsZ/GWdL4ux7qjYmZRt8ZcMsa6/KaH32yz4
lyLutpg7hp0adpdjFq5JZbxJCK8xQcFFXti3yxH3BW6I26exCLhk7BymDLMred4gp4BGHWTz8abu
kfgI+MjyDIEpvK2tlKr8YdGB8awPZzW+tG8SZ88gWldO9bBmKjfT0fyBpYVASeoEe6q9TtfRMU50
hB8jl/aP3UhxmuM+8jgOueN/D/SU8+HxBW2MQIm1/jqMNusYFxhHmhZX1AJggwuNAJLJiJOazII4
h5fh4bOHdmR/HMU1xNnBCv0gcFY++Cr0GQsK5J4OinDdJPcZWB9sy7LFJa+pWvNuwRVlHybKydeD
0ljQ6H90qaXvZRuSlrvw8eJlUYswY66AFGuILmGTj6owL9UF/07XN6g8PthNmrFz17O1xxYyL8tx
OaNvvTpCI+l96QHzkzMdxxvuDbIq39vbC6f1lWU3rUCSGiyDNMOJdGUjYLhZ3eiHF5DOqLxQFRfG
HG9bL4hLKqEkN6PitM6d7CDk3XB+f3T9kMq0RHw3byxQ9ldRzbDpgBWdGas6SZGWmv7RM8CSwpfU
fUsT38lRbnL8D2U=
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
