`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0INbis6m4LNo5fuoc/7VtaFb6U
0+5fXdMnwe75smPOBFJPEC7G1jJjzTejAYkTl7IUTkgZKL+qPo9QsJV8bWnGHQsxi3gvlQOIaFQc
GeHAIu5kCH4qdG/Rd7Opht+51SV6MCUG+Jzw6T7NCWSvcK1kUSxl+7AIlS+WIYISlJ+EKHtGVS9i
EwJnDml+BfWpTB9xPafHkbwEu3i47lW0rm65AtBA0FQc0g9XjSdqF0izkDx71iLWtwdJ/ACCBQzi
xKC6WzfTWdQ3Z6BpsrivoZeePhjZfiujcnb6yLxIBbDA9WUfDsH0lPOU0oRQsKhh0luEFez/GPSP
rkrsGnuAIrs5fT7UjKbNKed8lyjY1EJzNW8aY0JUZ4dW5h1wqyiA7NGp31VIvio/YeQ2qkMt7y1H
NhiNZEi5Ptds5rQUWqcQZjnShxHqgVt7G7J+wbq4ADoyNgZEAcUH8oi6YKuFCVezzt901+ifefJC
XjV6lbkGKejjrMVmNN3l6w/7dqfMq9BAYoBtmfbYSJg6J3t0lTeYwexBuU2vvYv6Y5x8zbWaLmw9
tKevzAWPWzmP8JbxqsOkYFMrsxcNGwJUiXZ8PJOI9hfsmH0saXOEHgHRUccuwgHF1LGqyonLVTol
YBYixOFF3kBsD/3J6sdGSQv/gQXnzf+JbEomlT2pn3vRCks+IZK+0MqQeK91DaFJPxnYFYM1UZcf
1iax1/wgVprTnvZmGVd+O63wglzD81NFI8zsEZOhakbpxf2LZrNy3ePN6kD9xoZYldv3gkLNuhVx
RhSX5A8lLjnbfCi2VtD1hKCMblWNcRt1M0ArC2u7Jqhxaowtx7+oNFrsXc3dUDVQvlUaFa+wbZMZ
ifJzcB/j26GRUbmnH5H8SsZmUjmAxxWHQfx2AK/8Qdnwk1TSuQIXi34a0GRrhQTjH0YJcdZCLLKd
mUfrOmo9PW4NT9mVish54G+BwoJOQR9lMZd/tqKr7QDamIWD6inkxP5+zY7Q0gTgL66HSYA5MiSD
fpaRIpAUM+5IGwYgLdHV3k9GPGAnNa7bVS42s5L2oANZhGyAcNma5ruXeT7rEBYg/S86I3ydTdsA
qfghRQtBqDqb9rJ/oGKMCsO6/iCF7QDKZMMPjO7xryu5H2AbtXxh9pp9dfvVghHOee+wo0MlfoH2
IX0NTrmUTXM+xSmqa/0WsmnNP2Xo2/gNdwwLVdMZzXXfGx3zv5uYY33g6T8vsCGlpx5dUmdOJEmh
WDNZsuLTGu0d7/qzCssg/0p6diz09P3RU+nqrH6vo3q0976Ny/W2ZDSWSnAs0M5W9OjY1X6lTCUh
366NhnEciPevIbe+ypVtwjYtl88ObXb3N3p8e5vfLNAO0yTFb0nCIB904uZUPl6Cn7QykmEY00m7
AbdLfRUPAGDhl7og9GpDomj0lclBnQ0AgGXrUafAbgLUx1OkTOE5tNevscRD/6+6wXfKUr271UkC
vBwHL5F9iUm10cvomSteIen1igU4zpXmAGujk8N4GbyQaAauijZbmsk5l9b3WTNCfHzPXaPpRH2g
sT3YVwTQWi21yTANwWdKqofbtvhMChNqf5EWRSqDx6oGw1PTct7ree8UkSesIERpNezs38M3LC0U
PHGyMSeUoVEXR64PgpzlSC7ZzsulczhTTha/nCx+XTmSP1wcxKAk9JHi1gK7HCcxrM7t6QUEDIle
1gIs9G6M71MaKZteIy1QE7xawCWtaZynBWISJAmSsMPTLw0Yl03YpcJTY1pfBYeZ7YKK8NqD/Nnf
kPD6f04U1KzXZbZsq/iVyuEjF4nwOJceNAdo3ODN9wx/nMaAV5/J3PgYVEWEQTDmsYZYOPxPEUHs
eshxkwpPJitx94+usTKDAbIU0JzJiVCL8sf85sx6p7cx/f3ik9qRsjJ3rP7Jte7/P/9qhFJJeW47
U8EqfEyTDBTWJDvnXlymysGN6L8XG0BqwARF42aMb9Bi/weXGjZl7AGpDvlU/xR4PT6D2w21jvZh
DskIEcCG6KGjl8/+XppHIQ0J6VXb1vd6LFNAh+i2GZ5ZvjkG59VAIDfTRzLwiv6uRZ34EhUON+QU
KVT89KHqnlBwVe+vMajNXD5q/VBEI5flpOzdmnkYSGoyN6KiMcttAjF0ir4wJBo5c0dcFIZrkBaA
uc+OLGkSuhFhm1OEt7VG2Cutr2BKYE5bjm60+J5t7EEuermPDjUj0kwZfCUMBgYtDxVE8oXUvvHE
RBYlipamkUDljXMGbtJpPBXBopKdYCIMe5joFqB/MujCuD25LULZfixkurPsBf7Zwrcp9e0kzv6p
p857nBLbOUL9uALq2B39xw9KW1V/xHCmPcgp8HRo+MnHBE+DtiD4tv1qnKNIah2jukjHlUKkvIq/
IzZvR6qlhrsw3CBP/Mx1+GJ5MNTy9ui4lGG+9UcvWUQbHqjo4sFTRN0k60nUNivwMfoONXN6BQ9/
wh9YxkVgJ4Ip98fm+9hcu13jV8KRvVfkud72wX7066CWPg/aeG7gPbzDiidhClfCuaIOdhf5WIDT
yXu8hMi90AUdm+K5uP8J5GBzqxqSB2bHKhgK8WpVe3SCUUCW7vYc7Kmooa9P7MDTpRd79TNAa/JI
cBxTWQ8YyyGraHu5lv85qBnJ8pyRXpIX7raHhTD8GyGRP4DxKGE+LMBgDJX5FbpfHgCh0NgZfw7q
Ywr4Uj9wRJIFRN2d2gPDP7bIo2HcEvH1f3NwVoCA0thhQRBKrPJhA2jM/8XVFmpLn88p7thTAn/h
6jem5beTE3Vs2iWDqzp33GVPjZdPdH6Nt3sN5mVnJXApsUTn9tqdMHYlhG6FjYLj0eKvBONPAvud
csXv/fks+3JFYr96k8QRrwFD84QdjV2lHY1x5Vnm0bejeKZz7zq/VE2lO2Xzk8hPzfCez8gLiVO2
Psgx0LwAt9GGQ65LlS6lYP99Iq4/TY0wZ4oHEekRLWIs/f2VAf3nqyFJFDvkrpAUAwzXnulCvp30
jSp7DcpFt7kBx9+976KfSZuGLXXeDKEVOlz96NIHUcjIHb3nUc9X5seBaVHnKvCiYn1c+Cz43IGV
p2ccEJdnlMErHt7ZClt8DLq+O3ttqrj8X/e0dzSo6LUAOW+rlVtIjaCvUognr70nw0+myqu3v5Nz
wWU4VPUknHQ1LKwh7WdxMCvJl7OGXo9kOE1QnzpcMul6o3jR0sSS3o4o7SGz9xBmsMGey/tWc2xi
ZqxZy8lmQkJyhB6xTJMn6F6zLIpgiFlG1ZBCdEpP48Ukh9WlGsnXc44xRtfPs7SfejlLyEI4TyZX
MdnPlVGCYW4RORRi7Hy+B/YFHASHXtk1UvaJhlbjgPnb188KTeGjQGF9hPiz68Wk8HW9jFGuFJi8
fgVpeJxUUz6xAlF9LfLKm0B+bjCRGmx3nGMk76blkN97lAdpv2aAw+5WgJwBkfFLtfz1PP+WAFKZ
VgXXPeH3f3mBAqG8uo2gQz2uDqevDUOFbjYymNvHZ9BPoi0tBF8dNSuOvMPO0NwIWHwNIh3Mjc7x
9a5sB/xnx8XUsLJCD4BhzoFQzQaGJpsgOcijTmwnc1vzlngvCw5+tiG4WoSFSPBfM9nEM+A/Mzry
rfOOu/TnNNmjy81C1IgtWh3fJvtFFhvQSYnOss/rdGvYM9N09+an6gheh4YF39bGgPMlU3kOXxtV
AYEWG0XF6vMyrP/KJFhL58YrdDzghtUwGsVXAGS2yNaHDkl/S/NUIUUbCERRO8Ux8xL/zdgAUbSc
wjwHH26hDzzuQ7vcEgiDmJb2O1I5vG+NJM4u+fvP5a8XkRlQNa5EXL8sFKltTliHe6HlFuCRoiGJ
i3FNGsQskrA1PiVqK2K9UkLaayKpgH4YTSene4m08fBBoFHCld0dI8UHLu+7viQTHke5BaiUdELc
525kANo9DwBTGWudSprbFlj6H6wGPuSMvucUiuJV0mUw3qrioox57IM2A6KW/nZdYwXJSy4Tl4mB
ypdIhqtDXhJ9adQwxDLpShtDFnUdGjB9YdMEhbqj1SpWFRiEqHCgholIyQ8NAcynfSF+l6bOPePM
EzhQ9Twgway90VDnAs5b/tgNL2KuMeFVcvsP7e1RSf3bLOeYUG0JABb8XkDg3YbmgyC9kIufOQr8
Bek+e5Ot1eNRaGEWYNVJkSoA5mPCu8o5Fx+sZxBp6Wkhd3ZPW3JW0jldgkl1RbU7E4mD1fjdbWHE
AuRVhlKSTUlEgUmnSZbnfFwdP2EuKQVJfAyoIctRn4PlndXW0QRteKUeJrD2WyOBUPeTDRtBkuyl
/q8U826EQPthqq54CDoMO8dCH+7fewOA86MbVywQMUZLbvko8U1c56oKFDyQE3Q+QQHvY1JGKanO
CBkIx8h/kbou9RtEfdgzosGp5aWK3UwK3lZbCjRN1YW0WWk9HGt6dCQAzr4a2etomp58+E/PZgA6
ip2Vi7CF0VcyaOt7lr7q6KkOo2Ib8wMFj7fJiqyc1S1HrVqbLbPwTTqrnk5q3KEa9SFXe9QKTMb1
KZuYwfFi/YgWoxGb733CI3DR7idZYSZ+LyRnxeGv3NIlmsRBTZY9xTLFnguS9vUiIT9jp5G/0kLC
B5gtpdPW9Q9NCWaASAjPUtd2jOrxsp13ZKAfqUyCCrEdps+T9RcloU9ccpRp42Rhz8nzVPMEO2bS
whrgLP545fOKIixHiRY+moCh6lbNOyY/LBvnc2AYQuQ0SoLlZI2haSkG9uJ5Zz7Z8lMVosuRQoX4
XTHUNxXIOL8aeIFtvZ3JermfEGKDcHIQN77Lf1j+aViRQUE5t2yxGSu3fGWJkXO6CuisTQdyzzwZ
pS4cOBU0bsKxwe5tt0l6uwtXHL+/kZMFvUOGCm8jnea5NKu/fwDmBwDEO4IcyGqVVpAbTgv88BbL
D7B+SmGMTEu+21YOBoBHsKwPb9SpExZo3cF5Dmb3IG8hs29yanmDlKnMSLibzRs8oodn5ql0ejPf
fMtSz0OWg/Q3DYYfLHBbNondrP4L2Y+l1qAAkleLHlsAzI2Y1ZRfZU3NvoNu2NpKdOufkJO8V+09
JKCIaR53ZvCvQ+ak9l8mg6iYFej46nSyafqG7MCLiMFTnFAGkrjl5q93iUOr6nMdI257P0S3YeTy
VkYISnlIWQ7FfTHM49b3EsadhXQHWsc3sCjwpeu8LDtHYA0oggj4cqW5FSkEVTL8bnYA1+FFTaxk
UfFwpIyUqCiGnDCEblfuJ5JWUMgL9BVzMHeygODxh5BPVuzvFLS8HCEHUFo8xRwtfQNU9s8aBapL
gb2rki2UXtx9/viGmdpA4rmORukYmCLL6VK7NWB1YFE7r/we18c8ta9vVcAkhIw3PEsH0XFV/z/j
vOnEKV1CRrIdOBh6mqNjNJrSRY/TmYT0k6qhmtduW+gW5d8ttdtNOYNw7cGMfgPsYd6hREDpPy0c
6mAVqWi+DiZAgChzcyPI7tv/9o1HflAxy+XvuT/DPvQonmam2Wh4wSS4+k+xgsm83+CzaYZYKyAt
lriOiFVH00gkBl9d/mj11UbQeAAaE3+wsy7EoDh2OQx47jXuA5PB0i5Cgyh1EqciGeq4gwit+S+/
uJJya9yXnC4FqhFWetq+1GwF9tBjxWNPkuvYg1zk3STII4GrBW0KFT7OGOmZ+NjmiQreS3CmxcuJ
FeNy6xMqtgDQRm3brfC5kiIY2ufHQ0gSFL8RXsFqxKZ9uhq6ISc1vpeUCO/4GVakN12pfo6H9BRs
/3J6sT2rdFiNUKcSN0Rh4vkuvGXThQYEbj8d5+oZopwRtDzCcn4Kz4bM4IwEBYcCkHkre1kPdkrC
jJHuA9+fHaH9bPC7hHmMeDTPddv6z/wA8CVJcNgSJZOFsUzj9zkjH28waTcUiovxP/6YbISJ9NHh
6sTevJXyKjZ86B4NjqDz8DtadUOnFRFsCDLFbrNAqDO6sT+VaJlEJ2NLSytnO0f1KEmsVy7OTVhx
zz39ts2gOpcihzSWwA0zk1c1qI57flPB8mKfULSqWP6reoUzZ2TqAcPtKWgcXt/7XJZswlThzCCQ
ZxsEpXhsxnGSpY++FCC/auwf2Orij1Sm1Mm+vGZ/Fxh6/lUMRpd8XCi3JVNHuM/HEh2dGqg2mlbY
K/BLkNtcKjN2nko3NXVSmySI9KpUw1OGE/wo6MbjvN023Q5iRKujzFKhkSGGFMw5AJ1ItKE7Hz49
PjxBigbn+n/AgVSGC3RUHgoisQGajHvKzuvCzycnRVM5a+atdRGOafu9vJX1SBYfwqgZlTjAAGPa
Mmj7rEB9YNzTcjV/qJTImh/K6HGvSlHgSNVGEvJ3wr9UAg6kU83816vVfl7ZqL5ncYhyVVM2i764
ntv6UXeRcl/rC+m8cJ1b0Vvghj6W8pBCr/bZ5CWDxyobT5scnnA8aGOQDC3sUHYF8VhCU0xan/ar
6qrJTXZKqSVdJm5cUQ73FWFBorIAXszA2X+82S3Rj630mPFfnQr78rg5TABLvewqXH6e7syMtBf4
zifKDtynaOSMf8bgFGVjPGYWvFITWFkUxTz6k1oRRHsp4ZeqPoMrGhA8oAaqaQLtXHFcU7MvmoQA
5qdMhjpXsg4a+PSvl1EOM5RE3zMjbUoqMCnVIWdGr4Gjm3fpl1L1xUmZmYXs3Hqws8Pj5U1qfAW4
w8MKczD83/1uknk4vMsk4R6sBuE1a6aKZQXBSkilNcJr90vd/hu61qRX4ekbuFuOwtcxT+uFqu90
2aqKSjfhpr3ycCQ2rLXSvv3g4+OhDSa1zwwbpHYUaJOKCrYzW6YWw/0I4uXityap6gXIox+c5Oqh
+JQtrsqruUZGbuPzBCyBQml9CYCKaQYMKScVUQV+mNwAdc5SOVZqp5zOAi+IqgWX5KjouFmSBR0h
Ay4IOlunKQ2PNZBREntFZ5x+Dm7jjDvlKnk5D0y7Ok6Bl+eiDSo0h1GjqbsT6qPlMtHV4CkiKnlp
AI0zkEmGhUAEKUzH9XtBJ2zpTBenrw8/pTp4mcZY1L1YRSACJisIMJAcWlku6DzIMlBvNz4jBM7H
B4GzyiNlrirww9V3rbDQPoZx9YIEFXYbFsjcnOla3G9OwrO9HlAUOpO9CbGSfrvXJG/cSK4ajfjI
TUYoTSLAJFtUwUeMkf+lHajNdqKmJIjNxtvQ75hesXyZVL4owU+qD91N9wWEjIynKAyeopFM8fKq
Q5dbcb6Chjf9UJkPYrN9jWne9Afkh3rzyO03Tvx2bwxdl1JzeToJN36Q7vEbcrgfqCukKUHPRcmA
g8yrrO0rM67fS2Y+UHJ9+5FKKU0WXh3XMirJUYVZiUVNS6wb+jdvb+aGYdYJ4IGWA7k3lheaacTu
i/jS3rW5VfqnDPMFOx59G89hjIkBWuaM1QqGuQYIdJZCETSNm0F9H1pR08OsEImFYnrQdT5h4qj9
JgAz1XmfrGI4CJYwQM2HLnH6kUHkFF3PCMg/I5o5gWi518tyK0k3mt/5nIMwvV53sffz5V4Unbsy
VJaq08qaMtXI/wOAJvE5vtFea5H1LQkXxyDUyHKW5k5ywiu42cNGIcVpeNOzrGtWEbMEh7bVXpGD
Yf/0+oM7IQiQFhjMlZOu6iV1b3oSPWih5BvdQowF4yo6GlTndIrKHEfPAw3nc2XIRlNlhv6j4c0T
rU4OMXphac7E0robXw/KdasD9AshrslC6680y9/CpD2D46F66iF61OxNDEHbgYrTYtCAnoj+pMIH
qAu9V0By42Z5IAQ32XFVEXmxazLy6dmBW5kjr+dIpICx1N4C7udtbwM5FTlHzlVZL60R/4zc0uPY
7yAfV2DoKa9FbrsSsL6/NFK1MDP7rQCIg4zlyr7/Ebj0XNaPDmcC6NTkIFPLI87UFjR+fYHYcEcV
9BencqcMCN43BlACgIio1uQREeCHRXXcWuA7eMdOTeBhDhFxtrexucOsO5KpnqgoHrrjQd4M4pgA
wLRcFIBVI+3iqTGKoDlQa+Ikz6/wxLqHsbi0ncoPCEb9utKnQyNjjx/Lxx8csLBmkrm/6Q5IPOiT
dGHjHJSZS2mz5M2IdiU9MA6zwBPUNli4PzEg2aj3H89QR7SsV8pOYUrZhryz0ukMRiG3zrSmZAa6
Pi+z/M0frQqXTtTWC/Sin62giZjWoSEVZIIhPwoixC2j+V52Ol/1xte7sb189sHX9tCmuArFZX/p
xLPMZvbNeXxFGCp2KxLUzW/9r/b225qXEBCr/7985Y0GY0Enu7PpaY2Kx4KVknG2OQZJD75lbHwd
CA1pZwehG3j24cQchxUsfBPE7qTq0OA6hkfyD83bRbyTChodA0NgOglcooZgxpaIdDh0AfFju5Ri
3D76g9bi4RDbisrCg3JiJWiRko0k30bOsnmoIOAtzGI8dU39BVBrrbMbmSjHmOK7qpibNmBwJGcq
sBF3Wj+p5lN3u4maVv447ZLmOFcIrmFibgrtXrLJR7obko3Z2DwTwdQcaqYBpdzH5cmTisD7BzbH
LWPEFr5Eb37YJPfwMjtzzDCrf0izb7N3+Ic9rl1iK2J+NScNfpu/zgIOWV6Xnkm03K9CrUllMl7I
dFRFh1zCQ0KsLATO9MU8VNV0Suc91eYGs4mzMazg1poxljXBOp44/jg9U2csn0rupHC6I+nGT4cO
AqOWZN9YCZB2wpAasSPR8iRAkvm3VChSugEdt9lkxdGV7ZR1zQ8Yid4/bL8uWwAu5/vlmShphhQ1
ZW8OC6vK/0T0snH9BrB5Mu+loyeaimZ0GZ6VxilM+bfYtfosdofZjidDI3rUXaW1WkyD1tOMQaZR
tn3Q7bRBcK8gwyEGya4atx8sW89+bm2fLQuSmSM8yiH3UhQLp99D0M77feZkaCxcOKOVeBVnQsu7
AU1v4g3rqICJMJHZezP5CBYnqXOsLXrFUpM3MUwTjFYvHgcGnhxSINXkafmSTioi0Yheo/CS0C4c
auO80O6Nblag7dfAA0ln+pWyXDO9FqfAYz6pKN8dEW9pveAulX+yP1a/icos1KNrbL6cWYwFTYHi
lUl3HoCHqfOS8gUAwQY/dQYjDdj9hhs9BBGrDInmKEtjbDJAV2BHucz1fkZjOYzPxsFaOoA3LNSo
YuSuHQ/2WoEac9O9sL2rk6jgjyVsMcwOsCv3PqzUbnwXklCDz+CAJm4SzsgZqc+9aQ+7Qc/K6PFg
UM3QNAbaH2tE7uo/OSF3UU/Iq4ZZldMwDHM92LmMU/ADwbUE5ZpQyx8NW+SPXPnriyidTh8BNPJR
tabUwXYvI8Rme8YwBQjYMuQsewKCGr2J1it1iickFL8sKjLIOOd77Y8seyXOD28ZyTcXDhDSa7jG
G/toO9k5PoUUxtWxf3dw4I8u6VnOp114eFsbob1fvQGMOc013keshDbaEqCwfTABIrdL+29/e8Hu
18jpkdlbyVpwVEBL7HmTn/G4NZgQntqzc3MR3o52cG+2uRN5hvssjyqgzct03A7QJFPkfynLpR56
maAtwwHbSJvF7nZwZcsoPTEozjazGzrvy/wpZFVH2uu3niUJRHYI+bKdnYdEM5Gd5dgWVNezvM7u
mLyzAKwcXUtLO9OdfYBQ3NYS6FF9VRMqXduMi1Yx+rg/HbIG6WuF56aQ2DidZEUbUYhliaZHG1Zp
MK4XJSQ5C0kpsgYM31qAc6uSjnau0CYrMuZEzRyII9Ld3kijH0NN6HtWo+oH/xKz1/0x550Qs/Su
VE6dq4wgFDYP/YbX9ko2DYS4dhdNqx4T/DHc1ACMiGcQpEp5I604phurUi3wbnqI526Gy46+ZcKs
0/Adl2M0byyEa9LniM5yZi+OOwt6gUEJ+IrCeMA/SI7olaITJUKB2GlpXhI68btS/GGCbHMP/ZSE
HASjYJGqtsFSnQ+El0tNrSecKH1aAiw9pEX0F7k196vFLiie51eVqW8l8jLcTkzNTiz8NM5mhPdH
9lBIwt/Wgvtud3HzwVE91rAJqnulSY9751HqFFG1JZgP4bN6FKNh2AUGlm7wivUCoT18cxddTEhQ
wUbJJC66Q9fmZncmsvWDak5TjMp5ZHzzJhFNDbXojcem2kMdZ7XuFe8muv8CVxMLg0YEcARsWkmq
EetiFpiT/InXfOlT5DxZdh+t7NIZXDyeV4Fr7Heu72mABciMMpu+6KlpjpEIjswhZgie9xMtPY+T
r6hp4zLU1SnS2YssnWXgOnJtLBFg3/9u5Z9aywQCbAADRaDVcwjZd0XeHCIeRPL5YmWs5va5UMkz
Txheevq2sfJirTc6jp1Szg1lehDpSpW2mz/X4ttVZKjFcXnP32NrO2cX4nMH5bZvzqD87uDVbvl8
oQditzJT1zI2AyiSlmBvUoBrf3l58mfxNFn0bKwOmi72PUeSS56rOLi+8Lvmfn/Ek6TO5DTh0HAU
QMhNX5yXqVM24/PV5+Hkx0ETcZnADGfERIe/DZdKKCfX/3r0J1ye+A7cchwOA/cDLRP9wYs4wGDf
g5BdZux78C36gdKLJd+1BCtrkuDVP+lr5zaiWdEmo4tZNvcOtm0ZpZrvcGzscXpYFlJyQvkhVTtw
LtF6eUJ2/fEbW2hQPpFoYLdRUpFAGuCKKgkAZBRFPL/u6ug+nMkP1yYWT4/wQRbobI1ZQ5uvy9RF
iKpbJn5YmCNKYCg8WaI93T8SFtU3EejE/isGc3BeWQgr9WTJYfhYnuzRyD7FHqlTiFqY+7UpnFjw
8CAuHh3EwjnsTscJqwEwjE3oQ5SZhcx4R7U6jDEPRUzZFvelt7Qt/DvAzC5ICQ5sHtIU+rW3hQVR
udrxP+Z8c0Niwv+hDX2hRV38LxUHpPsli/LqDEuF7zpioq7ybxrsTvE1WIJUPG/fqlQp4ljdpY4k
JRukKe3f1cg7uuLcERkHlcM9dsg7xS3BttVA8XplhBi4a0498KHU85aSiDKon5ODxm55FnNGm3jU
YEbQJQfUSovpuDato9cCuSF0PRsBd99G6F1dFa9qU8nxz9LjIn9EueuWnaFh2Y1/OiwGBrZbNGfx
nfWeT9mJWBxSAVjydYvdTIDedpt2zt2ZAS7qFcDYP0lyMeC93zZjNSreUX2ry3iKjh5KuMdUUiqk
7ZG8aesR6NKoTTTRwFwbFnhd2Wp48Eta9PltgQxkQStuvqO1NwG5obirDa6hQBwCynDCBg0IPn9S
xSuVwd/VsYIlS4VLrankRzCy+wiVx8BObDAdXV4oFtAjsyvAV52o0WKI6tWZf7tCI6Zl3DXGtW5r
vs+o9xOfiCtBQDGq0dhcnyH3wYPqnZis6sIxCS73YdhK3DdmSFk1QdI/e6PZDOg9Eq/lSB2n2h9x
/+ZoUfJ8uKLpuCoFePnEZYmgppeYUYodwWUyGpR+3YDLqlZHa0cosN+w2+lxF/ROeMQELOtbJVL6
5P1PFZXIFlCLaF19KPDAhlRmoUymqPiIFXmzyeNTrsV1X8f03k93xfpJ6uVPTjZnDC3JX2s1z0EA
CEi7EjdJFO75BSH+jvLLumbwwTwMMoM80BMbHe9UylCEG44lG9ehuCeYx6BHSmZBA12h0p2fzHEa
KHxNtzLINca4hoqZ6Sf7tJXs0qJmWJlur3kl5yIcO0Q3gmy9vQvssgpGbFmIKVhYj93jUcClcx4S
GmX8UwiLILzJPTLLFrp6RiqVFo5gBGExbPG8OvYAK6nQI1CsukNoHJGu/q33GrmVGk8jGfxF7Gfd
m/2ZKumVUJs04Tw0vlnf1/tJZ5azK9CpbEIRsBZ3kJahCehGU2CUjo5lfRDpbUgnKc//TbbMlXUn
rh791ndni9jrrneWoqNIMLxzWDi7j0LJtEnrfPgAVooNTycYcF6+yphBv7zhZnMG05g+lJidZZay
Y/4pEGCYr90HwQGnA3Nvk4XSlWx/BNr8aECtVDWQPZonoV6Q7LbBMWc2GuQXNBT1MYxZTY2UZpg4
wgpr9Z2ZJ0pCgu8gvf/k2LW8fV0IPy7fWcJcscT0/nTBTC2T6RcwKwBj44DFQMpdQM1ASbVz7HtR
DIonclpKowFCNciyHfOAN/24Nhd/FY22ZAc4ZL4+fYwUfsheNw5bdXTaxkB4x4npNFJ6FGe+gibp
cxG2vi1FUiAwdq/ztTb82Orlizlv/FF4s0Q8i9jXpMN8VSkb92PuN5CtPMIrhx14iYsVE8LGSfL+
7SIMmfLwFh6uOCYXoiRWCZ0GgHkRYfwrG6tZM/NCeMsBLiTQIXMlHjXQsCKjHa0AkPjJ9l1Hu6Np
92ielOJ5nCflUdnDLnH4+fk9ar99aFFhu5SkZM4+02zpNA7NNKuBmKi81CuyDEL2pS65aAbet3Xl
TbjT/obOUGHG6Hc95YArlbNu+qxV/EKm6M259tAVp22GnByHQ32jziyXxOrwYKBsfoLjmjZytAga
LLo3+0Tl9w3/gY9PLfmacbSVqzwEAby1R0rMBi0azXnFo/9pcYdQ7uRANDJ/9x5DAW2kRfJ8+V+C
DXOPIJoUzZeApImsdhfyI9A8SiPztgGHjcUw/xGcUUqFsL/6dD9V5nzehPFc0VH14RFzbSadjQPA
h/D+ZzgP/AbpT9wNrMOw9aWRz56S2kP8/8z8Sw8fRGeil8GMctOJGbNe5g7vc25tNPPW8nMN3bv/
cKQF3eOTgEuz8KqK+4efjxWe1Ck6KPT7LKohiLh3suvVnoK1x5ms7GGBRgpH/AV5hGywHKA8EU7Y
9zi7SqZvd/3yTt0J8vPt6RU6jqufvq5bDQMlAreHQ01d1vMdktpj9FKyJDogYIsyHlSiDWuFVS+5
rrRih16LShbW1YJLRTX+8B/ThVAAQ0d7EAbUVq/8PwIsoVQG7iaUpnStWbrndDnVKfie0QOvLvvh
kmW/jJMEZYeH0lRR8hqmCNN1xwIC6UHDu6jg2OPy7XO8xkoI+rVAoW2Th2GEKE2/CSR0IOywpQof
2XWnPAC+iKfu4BeZWzxG+isP8d4rBc5LUnzqbQjdHzEKq2IKg31qK6bch61/rFipjwYlMa/bzUrH
qKo/DNFpHYjWD/8X5wH/abL5RArEy3RvcirwTaKTTG+tXPMkF1e5FN8XBSC9MWH+2LiQfc5aUeOc
EGK06srJALwbXy9zmMFQL9t5mzrIRxl4T91MXfNinbmzni3GXZSCVcoAI0EpWB581I6lxsR9hZPc
6ab8H/pcHZyO1QLu0HorlXfbZuGom7az3f76v/T0kMRExAmQhO0zzQfvnIukkdYGBf1UlHJogl7D
pYcmndCJbVxjBVj6FZCn+HHmXDVc1J8tB+5oUGfORCecnya6BCwogeSlx8U2hhAugm8/Itbrz8s9
pHHoVapUXN5TUkM8F2/KMINkmRRkgYx+i8SZ0qkBN6q7bA94DlZukgWJMYJaLGaLVZAk5bmlsmyf
bsLFFcjZi6xbfiYL2M/tIGI2F2x5a/Efi6gcZaVw0PLtJdwsjhcearj9mMemKDiliDVBcKCwOMWR
GvW5/qXJVnHflxQ9u+lW9yLiQjahxoYVpL/FPQj//43e/TM6qMV0QJ+Sr9lQV7HFoTbTvygo9bIh
HRGQfE0NG1D1LlD//l3u2MPf4XgsAvD1CkNdPeHy74Ibf373UZRSVqrG8GEJnCRu21BRK5x1wCq2
A8KJz0cL25px7ejFIC46lrXeFG5qmMU76qzjOVevelharfz0alCRrfK6xQZReT79mh1t9O8oIMYG
oQOURh0d4/ZcnypDr5/h+vplFGT8iwEsURyU49UFpUoQmFvwWgZMGicMaQyX5CxBHIL8q/HeOHnz
MGgVsxfnzB+VJfA/olT5Nydn8bkjJXwdQUvuYcCPwE4LvC0r667KY4DFLFfIT4Dd9ljNCfRvTexq
GTXhEGvIjRQaBcNSfcpA1jx3eGtYYPHn0pOagI+bBe8gER1gGRtv7Ye7udwNxwJ/I9dKe/8PdhQN
rx7wg8sG8yKu0XhkhsfoeeS6K67mwkkrPa7rkbF9IhJrhmA7rMvDFtMEBkWIO4w+SDwm2ms6YQBl
P0eO/djaSkjJpIrjpPImi7T8n24yMtHlSvQP0W6V6ZPpgEuv36sPjFQp5Kw784moHlrX6KmTqbos
QER19nifYn0wM5R2kYdfRIJiDrzdf3PStOxbmfJTYfeUnkEyZFCBdO8Ii5U/qEGfZenK1h8IcBuW
Pi8YCNPsNjJq2m23CYKGd4tdNxAf0WobfhfilfzP5jZ24zR+ulOyTg8oWYK1+zlhfuX4AI3yEOOt
ApoOlA4iCxkX4NK+gMgQ4xMZzbV71mvgvWm2lOzOh8KNglpzslG0YcfiAvyLR/bHoROrif3oKpNa
+7Xp6GK6jAiOpiaM+vzghd3Q6W1N5W7/9+Iy5qk5mUJtxkjfeuIyk1TYvc0w3iAuAR+dclHQMr66
pjsajabwHxLRqPnhaRl+EyBUaIt6FOGxXEnAU2leduCPW7VDEy76qh/0QgApbTYKqFU4o1KSPqPb
xCeK7GCTx1jSXzsDXx43zOZDqsRF+xT0K+6YSlH0kYWLhjuxKzu3YklJqqnuVeZ6lzAO6a+SKLtl
SNPTh+FthKuN1QW215yVkXIFgWe5ZlMU1+CxxuIoh5tKXIc6+ioaKVGrWpodBV8jxu4hkXnEwcDZ
GeT6KB2fz7Hx0cmD/v2fJlMBXV8z1D86+BDVHHXei5GPP+SL7RMibAooPXeF6LJb7neBdWID8Ptv
UhmUDYPWndAqDcXEn69gOfxrC35APlfVUJNCG/olbIrowxc0Ct92biqhftX41/LBVMlcn8ObZODQ
fj6+hNASwilbeG4+m1Y8Nb0ov4z1U0OCK5Ka7VEKR4qp8XzRC3W7Zl70ovo7OTAXJdveX+b9T/bb
VwxUR3cP7/DD45d6eO8mbGRdQtXjiCuqssoEt8x8MnpVs8SyrmF529svw+pKbfCS6+I3998ne7l4
79vwdNn1QTF8OEY7ViSHeKKdGT9pO69vneApUQapCxM9In1s6l//yyCPFYDonUszCwBG/c/XYG4N
ka+YucVyZN0JRuKv4SmwGqrCQWLbQ3hbr4+SNY/T2KEUlj3QniJPEyE372MVLFuz/waabZbuwbJk
xNLacFUPBA5V1UcYsI+ifXguj87+92Ta4ijC5lr+2ReEb8g5osfyPm2ZqoLCTpftw4/3cPyeI1qA
vZ8d5hwwOhU3F9FnprWA3o5zKmFOl0vX1i+DrE4skw/hstsV6AsJ/7A6GUnDny1NgeC57ACe+SxT
MZc90v4n6rsm8GTszxY3zhma5eRMMowxYy19Zm4vqE0GSTjM9n+T/xmnqDE6nGWOwkO4m1TbOegV
Yl1csSU9RoguwXG4c9S/89OxY+iEeKWWb6v/KDYgN3yWz99iDQSGnoz1+3f9riwRIAR6zfhMLZBX
GKRjOOShRP8Mtto7MSKi202AW5H1YToHQTKrb24JfJ01DZR/yIl7gS+dtsaMm5f/LCQ6U2ee4wKg
Bd/rO1qxjXuIVt9KrI3EfGoCor9IRtk2s7OqDr+fSCU21y1M1oFZ7NlGkIIaoP12PoH+PWMBiwy9
C8nWD0R4y18+TJ4RXGHjByfALm+dkgwbvPosGdOknuLWf89GR8jkZyO9VZW2YEwdQpb532rQABP7
H2N2vUg/kXJpAyI1CAuNS3Jf3KzMfLKdeXpGZ9padH1sEZT7kIVEkA9Xqk/T0oDXYjUoq4rw38BQ
jJCg7LslCXg9q70JebS2gULph9HMrz+Zu+1nK3WwG6Pj8kvupfSt0sqNpsU5wccvaZ7CBH+37vF/
20EVYZUU+rncnC4Cr/G8mH2/MUW1/CsQgvaj4dccFtcr3CD+ESvyxyqNdQuaYhh/XzRXj0pCB8F3
VTi9FRlSKDA9zKEr9A7F9i79x9JcPrG3ByW+CYJTHzYnYbGARVYiW/iaMBvXfR0T5G4QPYCv4YIS
0NVEmmJT97y/ST9stgpIHh/g0PeC6uLX979u10EGXl9R+FQNFoHoLRuO+KejhIBGMwbkuhfa6Y50
6zC8PLHdgAEoXYKDUtpjQ74adUDowhWum39NjlsjKgCi8y26S8c7N5eZt6TuCvyBotRnG6bYyKfx
dqkh5XSqi1mbJqXALX+LpnW9PDLmm7f7IG4oIm9nDiPgkue4YN6WQ6Ie22WQwrg/owBExqi9VV97
ur87Pnc92oAE3s9I7REmEfGcFBMrA95ePwJvqftPsmf/QwoctgjYrMpCT2jjhcmOasFpf1hHKwXN
QHOewLnHXKPMKCut+hQ1opaWPLI57CfZIw3Zzfs4IpwFU4RSKfIV2v89/Qcb69ISFR2s6ZXJhzpj
85rMtxuGpXTz49nkFACuRSl1kVzNmzrt0h2cd9xHiDIUoXbBhuZt38LexsEUw081zh5OrZh0HECa
7QP/sml74tKYRyvwlWhZl7OWz24oqXF92cgErUtaiYh3xG0otDm4euiDKKiHEZaLZP5DNbOFf3U5
1PDdJjsyk2LsT0v7FHZ7FN/Wh8ja4Ad0JJ2alVFbzLjhYnVjavylajCxv32CjxGrakY6pIZ5mPcq
FINv8BZTiptvzWkshMKrksfZUxzy42HfLj08BeKJmPkR/diGYWv68Xovba0Fi37CvfGWo5dtddOl
qP07vIN/5dPwiF45vpTyXFPT3UCl961iloFFJ9BFsR2e3VnbSWVUNvp5RGQnhsbDd4ayP38HTu8z
I+Coo9OtyynUemuvyna/Gd5Oofg7DPqngPEO8I2PJ2C5iVjvPqLWLiPePS/3m7j+2lNGv4CFYeU6
o7N0iFbz/3HS/uBMCSaHX/vkTw/Nt0RnEoda5Yg5jtRnKqf3XfE88h9ynBREWJtwBrr/0b5T0gsP
WTWT25X5Wxprf8d4tmoBsiQZPmrLS5AUfpWXEtrEFjhlSjSDl5kC4U9kC+OOH3KZCRA4WJ5YkSbC
wzbbT9ESb9uhhm0MaKUrdTJ+JFLsmjGzi6KvjHt5EJLxSMEdXXsNSpS+LcrzdPjb0Wbqe0Gz61u3
lSLs5zK+9A8JzDTMQ3Mg1yB/vjwXtl+ral/sUmyq3r3ExZSgBMobo4BRacMwHGd2cMxfKvtgoUI3
tTQX0LVQpCM6n3nnYl3Vh8xgwkCdY3MgQVr9b2/4f4TfxWN9B++JFx3kI5KjmD7nKAKOaymUpT1v
uy/lu8NieYg5qV5fxIOqsuD/2hxOjvOo8UXjErjjiXYiBlysrkKE7JmAIy/sbqwfMkU89qJX9qSM
ZJS7dt6ssfDSZ8ASQ8OqlODPA1+3MyJoIK/WY+9GB6mq64Qp0OXyrKEcqr0WFDsNSGti/dNqIUCw
pKs+bq68gesFN/qZQJhos72Ek2kIO6sVQgWAGTXL+p6l6ZRcVv49NzOPjcPfj1J9Zzayrc0p/ycY
YpsnYDmnh6idIky52k44PuddSRFeR92IwH1w2/PWh2Qozddf9wEfNYHUD3ZEQdrXtdz92sEyoF2R
9atiaZDoeGJUYDmjliFSqNYbLTC1ceY1bbBOmRZ+cGOqg/o7mo7NdVyuFc5FPJ4S5xBmZb1XRqO6
wOSvSjZPeCgimI/misg83DiujetSnzi9saVQP7Um6jmteJbAeVyENWwOj8ErNjqKIwmtcfSmMd45
bsu3RvvFfHjiFESZt+kotiw4vkMXbt+fXDdDzQ3xLuj4SYGVD6Jmg09NvoEHksSawk4QcIeTj8mP
djA4FSItvip3FXH5ZIjWpIs+2cUICKhDNEUB1JCb0lx5u8FGBP9/zah1QJdahYx589tLfe1b9G8O
+/DUQNzpmNjser6AQP8wx/napEq9z4Dnnq1tJZ/ppVTxE1yAETDBA1LiCAEaZVlMCVdP6GvQXMwW
5aLp6RPrZwKy4jW+jyTcUfcpUJIlEzl8Pf1NnEJd5jvleKVgmIEBcy/Itg111k/8flYgXAuVxA4m
UMezf7CRgTFih7MnT6ezI0CgiNpA1pVsd74Kpu3jmFRf9smcqJrcy2RYV+pULSImbRiGPq2s5yo0
jn9pCFGLqFcpZLmdcVjgOnAaSgJmG/lLfY3xiRl0q5gDq212RXGfrkt+TTMLI2KUmqaPMu4RRRve
zQC0aBYyJsSQp6ZVxb1epMU9ZB+UPPRqsPLM7xTsQ5loUiSJtB0FMQk8/ogUvZXyjIVxEMLQ7QWN
q0SX335PKwtpX8eP4awncdjJbwTvslKMgut2lVJ2vs6Ea+yAfmV0TnDgibUg+lJy3IICLuxz7ZF7
Vx1fM/X6rIqgt/vvj0qNl0LxhQrL3jt1eEwDg4ewvgeEHZaNMEuKyyi6J6AicWBbnHoT7XAZncvX
SKFqUAVhF+h17xmNuO7YyAXdD01xQI/fDdTHzMFk06cm2nQQaYf8hZD+RF/13H+yv6g63GBEWWzT
zI5tZXqUmb1g5SxgQTdKc3azOIS3SClv7dS00J8SLF++Z7gciMLE4Mp+sOHF6ZQ4cP6VoT7xMYcI
YkOuuh8/dNQUT3hiqhizi6DL2VM3eEs/2xQQaMJyPZKZYborNuz368P0mhdO4BgWHJ/9rxZP4fCx
H0tIAFzCFwo9P+tMzhmM9y3wRAZszkf+7w58jO+iutj1GQPcLSaMxQtx5Bx+PnpZApxrggU9ZiY7
q3w7ju3RffWPchXsotfxw+0SqlB+QWoXKSw/XjNUojU2Zv6UZRtKXU3VKkEBUk6Csrna1OQKF84V
Sl5PgP0Q/PjatpvABQKnMaZCFpQiOVfhiMFd0mdGvNHiCSQNa1SUfoLn9RKX2sCyKvPhFytpWFm0
Q+yfR7oDHJYEU+Nv1yHSL57QVNSLzEyST+becvspvQcUIwRqmaKYXVsCPtkCafj9JnIAdE4L0LIO
AbzObx5mcEgtz2yvzGXSPL1xNK8P1sJIBuzsxgjxO6H4RJ3QkPMOEYD1MFeGFAmRKmt81Pq4HDvH
Xvts7tZn3c9zQbotXtIhnZyTrQjwjhFlbaNfg6YvGjsJFGGta7ndlkFhO699hSIlp0mSxOCJGc8q
tqsM76FNqte2zyUSv5z2BWfEZyymie91Km+AwqSFVwv2tAWUlo1HrXLG97cbnz79dU89T/4UNGTi
sq1aU0a4US7YuzphFqr5NemTy9+XVHdEta70yP5N2Ec4N6LdyUCRHeDw1knxRxL7ab5N4oqnr/QP
tykG8+UWqsA7GEtV6Sw6jBsIInCNwdjnDmgIqRqf/xotmc/5zU70Suj5vcSdptZ3vkxBwkbfHTMq
Yszg96jUfoz/j/6Bd+SVdmeYqVOrEMoMEAQg+l1NOKNmqJQIjB58Q9ZRU413GXc+v2j7Varqho9i
Whi/OUc9w44xncMAdEXi0YbrYWPes8DnFvDHnfq9Nzr1bnmQ2F/y8xFR20a5FnhukVJjtBw4GZ2s
07YTl4dyz5lcMBSW283WyawnvLS61IOuc0FHzzgFPuR8s6VFvmllyrqluobOXCKmwYRvOJ+WZZqO
Kg+pQVsqedQ/YoEkW3hcHZemhUgld9cGTKhe/2g/BpQhHevnhuOo6CvCN4FaUZkM+Rs+G6Bt1woi
5lgROS2yEJlwAIgQjaVySY187npYbbLExdRN4MU78enlP1lUQDAXcipwOoC2SIPp6eR1EUM/oP+E
9gxrKCVr+bJgDb60QP0XBaJiHmnnZIMcORyz6V0gqXPkKKxjaR6B6Rm+Qpi94l+t+6B0/Db0rGyW
AmUkmb+++0sP5tTaklE1tED06VQy39qsCqERdP6TwsH218QSfDu2SLD5SZpWeGRDd8Ph/ju/XJrF
uBqConc0AfMwKOhbF0CPCSSZUSdpUhNscmx6Kz2uNbtotFCuNdQj2DPxH6zqAWn5AQXwH927QVhy
83dc6DuUTHbd2hdIU4K/BnFBuhYPQsgHR2NDk7/zlXGxaXwQtju43W8QoJajp5b+qrA5Fsq34nZ+
Ljy3qxsjDKWqtEqC07KWaqMIyBC4VnclG/zRlG+v1vKcGDOB8wJ4si3oZ3BKURRpTDfH3wBzeF79
w997uM6KdQbwV4zMKFW5ub9Wc8uQm906uw8g4iNiekUVTwv6UGascGnqTSocqQRngmaFUdLbqOA9
dlzsSGvHfwT1FEFnqFUt2kysqJSb2sGWs1maStSZhEHQ5ONksY/frSuHG+dOiBGk661theaClKgq
5wp+KsBjGJkjEx3qfO14SnsenlO5xxmULwEOyn2S9YTpm8XuMEzt8fP3r90Oe8UyXXTVsWEbvoPr
gu03Vg1xfpEWVk6+oJRHZI/JtJpUvu9yIMB6vWpEd/Qo2mQDeSdLRfXhF3y69z69uhnJEnG3XQRX
N/50GkS+V9aEkWQRokgPdiDR8fQW+iJH8t1J9/2AgynPGIaDxtfX3czZfzGOIcOsjGnQxQvU9L6v
ZLt+YzmBh903q8HKIMDocbVS5E1XecQlEbD2ulxItDj/0Azj/9rcVC1d9/7sCwIMpbS0ZsGx8CcG
L+NIlhw03U7siI9Z4gzDVSghHjBJxO/7Y3xzciAXy+ptYTF5m6dcmHrJY5KTMrUDq0zjca2nQVLi
pxL0TAd8sVa8lyAKIV9zPlrEZUWrFySTbhS9utyjbe5lT3gVQPW3UqjATT0tI4my0QBRG1ha/V6d
/DFV4NLywiJIVQoXeO9oJRzZ12/tE46zdT3yU1/3cvOa9mQIoYRd7GT+U4PZF4tDrD7JLMnD+N3P
SiFrArANx6su8vYAUzHMggVKq/g9MOmAekyv+ewEeUpsbd5coDWjthRBV/zCFKI38BEcUZQJFWcf
bV2uogp4Zt0IChzMwxH4ux3ovXg7fzt/JnDTSNJi1ugjkwsgYgVAjcULwEkdDfGIZLaBIIrNxit1
V12kqrH63brmAnXcBpJaYcqBEQaqI7EQerX/9g5qHbA/ZsGaaMYCQxHvUmtAvSS5swqsJhE+dDlO
UwaFR+BRcH1WCrqYSMPle0FhN1n+w/8GX/5wu7tx9hwVqV7rO7foMjUuHXAFD/b7cV/DbQwzkU2Y
z2JK1hJeAY82IZOJpUcxqFFL8zjH1JlBRaRP1gDJpWCeGfjly77v6JimntIlzB6ss2k4jyCkjXpP
kxIxIpzGAdyP5JlCp1VLFkOro4hv6Xy5bxOt6sUATJ3YE4o3FaPUp1itjxNm4fpJ9QUF+qeJlv/v
bfw16+5eFgCjb4vAgRfUMe2LyL2lAHxjRvEU+f8HTlWGyvl+L62xYkSCvzsuGUP5DratmHRtTL3t
slUlCbHt2GGkxour6pCCo03LAu2Tv8UuhB8jCxYxGMiZkhzfpGumzwF1cDLQhF+pe5b3AiN9UvXm
8faiIxzYhiQe2B7gf+iBYy4ttqE/bbWIJmjQs3BXXSaeHOx9EqIMroXqNz6LkIrC2BNbc/Uln6Oj
S6Rcln5Y+dEbSfwAnmY1iCQXnA6AFqLzJ7cahIjwbOo4SDDUo6UbD7yY0iG0k49c5e6iYHo3u3ik
xPRxq6n8Gz7tZT37JDkjwVtA9XcRE6buQBi045fgS2IuMasMWykw2+t4qnvbaYO+tsKvXIUA5wPb
vKcYJQDmQ5d9D1+kB6a07qziQQ7ExsrvOwDTuGTPHj5Pc6F6Rsi1hu3UyvhstQiZ3x8rOBW6f0o5
hvG4ATz560+91+xSjIrLk5EWXkz3AIza5R8i5SBKIiGwM6hySco/eyOTGDk8idwHWS6teyhGaTVg
Gzg6qMOnEhnxTwtl+AqrlKo8YXRN5tk/tJFnjQ1lVuhPkv+KfJZ7G+cYnPHlBiTazYUaTTIrNKqQ
+6v7JzA3jIcplbrN9Rlp9XIgxi42mNBAAJsw1vqt07NakIzlAs8S9kGuS3SImrY99TB+DMj39jAx
etP4EtXBlIxfno/4hRqfnq5VWpDjR/V2EVieD/1IckYDjviV5t3aXUqecDN3TktCJB7YE6IWmuJC
iEPgWxrFB9In2YOV7+7+x1PWoyyJ8GWKMuG1T1TVqJWpx0u0KmJUOwkA7tt8TxJVFo78GN19c70B
0CEygJW9Tv+lprnNHv2twlHYKGsIXeFlbFV7cjvwAvN7o15K4WktSCFF9nVrTEObv6OPZ8a29JWQ
ChjNm4OJgFpVTBbsfVPwHFEprRRq9E/hZYZqg4GvnV2zKMwfxPQapX6onN3efB3quhMJPcVysxRu
tV6pWVPhMB0+mcxS8C4rIPJjwhF8y4UBLtZaUfGxnz6Dv3dPCb/X2J8xw7u4hCDxkymWjlMfjRnB
lgZUSMrE8iWIW3H9TH3QmNqTtZ9wFAUBPgfgLvsiksuQbYz3nn/1jEqopvTMqah7R4G66ve0dQa0
sjRIMjhwf9QiNsRQQna4XGtixbt5Le3yyLems8EYVPuSbanzOkVk2l7bU6Tcm/nAD6oFrSpyzKPh
3zOmlEUSRv+Cp9imxJ1cNQbCFXRi5pw4T32DJ5Mls80MglekXetQ1M2+VIuZXu9t2lSx9RnIKdd9
HRUg4+Nq1VeHh6EUSjw7CrixZv+AFRK8K+Rjyn3olxSvbons/NM60vlsIBs1oadQKKM89R5XFvVg
JMMtsfLsMaCQ4tawgOs0d2TcOM98wIDhz9MZbpiqfzFrymoXcabyj6nps9fI85CgcC7zJAy9QNIo
7wST21HknDdIHoXfISP3o2InoD601EvkKy+r+SvCn2MPRG2UmzqHFMiU+ZMQgJkvYzF2cnnpHX7X
+8AGyINSE8qTs4YG4RMwW7sHHuDtDQB4v6ty6u308psIxHQMPgz4+1pJiedyUh0+WIX8sBwzoMMb
Ppi2eY7Abi+wFT3gPop4y9CIDE4H+nai5a3IzQ6O2566R51pPKVe9Kku6ddeDUqH+iC8RXxkcoLd
tfeCH3peaRXbhEIAXHw+QTqS5j/gBaGv46RvC47FX3Xy+dUfjbs2KqJPsmi1g4xAVk8SMxmZ2Wiv
+KhVtZAhRgU5aOLhZR6SPe4rc/cgU5DdojFh/AISvls5U+RXjskkYBJbHsTzTqNCnF/rm31YkxLx
Ft0xyk39372p0oC8TnukvAI1nmWnNwStj1T+fduxXU+KmUdery7HHoXa8vGfNg+HTDg/bQiJwen6
9UWUY6qLuJYO025NPRUDCAevG+4y1EIcisr8HfbxqCe2KJUg/1F6RCNOGgf53G4+2qshdR6YTa32
I1b9+erjq73GA/PWUGBO67jDZlOhHa0NNd+KVNdXwfBSNZzxAllle7m5zjZeqeugQbMHRWeNPrEp
EBXWrss6la2CL4C7s8BoRXbcoFzzzN6GxJ6qfIvB30MJRG5A59q0bPWFOrvtShqMs9eVYED3Lp/w
nAtIwl4qoLThhtYO4Ps4blojOCTQ+ZPuUaFo63IXkv1UaiF+P67EzDNt6C9nI28eqk3/oECkWM7K
O/KsJe/KwP6bKASNJivZCH62LlAyYhjtBm/ANAwVpvvp05o+LTRZs0SIDd9A8exDYWFMiCjoODEe
c7eGE4h+1axVR8p7As6pxNFDHLBXQ53O1myv4JOglwrRioU+DcyPFPOJROlLl2xgHDIhN5QigBsk
6gxy3zoTbh0Uhtcx/bCSq5NqT5XRYxRrh7kaYH7LVFcltTSapEhBylGYHPb5Z0vHnMNeHHvJV1Zc
NDbGmBKi/gktf6RsVSbPX++gKiZEEF1gm9Rpnu+9rKsYOBEn5h7zk0tHVtWxO0va+l7XQatcVyK6
OurPY2TvgLtaPMLIYjbJDxmAou11zg7/yZbFid2RI6Oc4WTOBw4oYWxxnE3ZULMnpDrN4+8pqxOw
kBymUpYwpXHAiZ6P6A4PP2/UfhofhS39RqUji4V2WouEpwk4tk4qGVt8sGU6jo8GVxIHiVmpvnak
tz6L6mDWFb2uEv3kmvzW/PH4Wzr/e3/nmvRZyAs4jY2/3nxx4hQcV0D/s4nAHHc2tSEaSD8IvzDd
evofLAlqHxdWnToJKDY/5ybLHluJ0pQOWWKeRUPzXr0OgNQ9kU+mMoiYKrnx7C7oLcB7YLwVhd9e
ug2fTMQOTOTyTP1lwm92px7wTW1B1Tp/h0GX/whgCdetjcM++2VDQ5CJsvg1zLTMc3T+/8kLKmJL
a84UP5+c/kgoBSuI3eRkVrciBdPVLzepOlQtF2kswUs5jynSyRFLEE9iJT38eGefwXZJaSYsFtZq
404inPHD+CkeDHc2cpRVdJ34NqA3eBPfNB6SHX69iE8BVmJzUgLrF3lEtxpPBReyGcMOVZ/BjAoO
k9dd+yITy2ogQE+Wsu4QPSUpNiAjtA/gM9/nr8osyY1NBcA7SHiy+cNX5rmipcM/AqKjBprrTwJV
7bUSRm0pIdZmQCzskX88hXuyYGBEyF0V/eYsjd+ARcA/EBy8f6EgROapk26QKHWv6NPyKN9uT0DT
di/z10OYvERS/ELOgH7mi6IYH2DNLMVD+8PnV8FJSaVoZDQO4lr3RDQWPy4cwU+Ac8b6JxDkIk3r
I/AzqGp9tZdxXN9w1pzmcVzXqUGcsaQBlx52ssJcT4Dzsc/7PSONA3PwFq64D2Ozgy14pbXLgSb/
wuFZI0M59+zY8XMPkaDAc4BHv5GH65/VYSPijD+DkSbTZOSfPWVoPF4OGhlvKcEpksef2Ul9GsZy
oFfBh5kUQLLo1LgvMpFKTQEo8WF1Yiw+MRmcFEXsUdFOMfbir+Vo2Kh90yagSE/WyfQ+np2xh8+0
4X4QN3+RXowdZou6j92Pmdn1tEvPP6eFoMwRIBbRk5Pssq33/H2ab/BhaSVGrghlIln4MqGfurjG
umo6RpCtWYds1Q7f2CrPkLDE0P1vPfCKjPFPdkfUx90+iY1M6VeobVvBxB2cX+PAIPbps6foCSb8
jz0iYV3Y+C0YocAr5K+WEHVl8lTIZx58tqRmQso4xQfmg3K4WRbeT46g+XrsrezAyO5tuXIGUHwM
U7LILx3OkDCwNLlfdudNSEzXgEoTrheQ5WdKaZEVWgiV7LCy2Y5ELFebWx06MnSq7yv6i4acXtBn
Oa8gL02m4i/KsllIXN0Fw8iiWnLNET8Lecqx5zEYhAZTG0Y19+Kb0MlTAWM73IWKHM725C3OrrSQ
7GMrW9qGvShN4hlaczB/MtlPPf/oh2tx0kl9LVeQYgkKcq2HUq8ZdTAyiB4Bgpvqm7CYLrXpPLPw
WyC1puAd/c/iS9D4ZMR3iEwFo9TsDrK+xvZpiyPjRzHUjd2wGBk6TODTN6EWdTftnGRaaRK2bngz
jVzxzaYxrHgzBv76I2dz5s2OJq8+6tzqbpKSqcZunvEc9B2VI9hh807ema0hIiAifJWukFMLFKcv
gLo0TTgOGwXVUxdoOLZUNlO+knLRZWoKF+Z+rXQUusPdj1muoTdbl19tuPitgyVRWj63IC9rjTKv
LqSphxAm9E6Txuw8DCeeVjxzU51l4ojIB6o6zyiCCyzYM6b5RvXEvX7IEzZAS7R6uFxqphYGePbZ
sudIAap4rUYiudvpQBovDpFdc7OkrtAt3QZAukNgRJsjhO3/uSPHmDIU11N2B4QiUmEsEvaDURML
uLSHeFjWU5VFawCsR2a2e35lscFXThger2DtNtCBb468Ij8vQUJYYtUKQ0kC1yXmFk+mnQ5C8Slr
z637fmmD+oiSZpzsEMd18te8PHJNE/aj1dKWDNykQMUmGiWUssxGfmYvF/GnEW2hqVHOGqueTP+u
ru61gRfo4cN6u+TTfgsK/xNSk3QkeMEwNOsNWH5AuUXPUsjGkc0lRgPvuew9Cv3KbiNulBseYMIt
QI+d7CX7QT0sVD1YU/sypNBiHVtVINIZU1I9I+ch2QQgaXfyE7O2iLBN9+BrEbhivLaqjqjASJdL
dWvBkgHPPSXMZngw4VIT6NYruFuav9sBjjm+U9S0uPVVpCr/HlM4J7Kyqn3SiQU43YvomIBy1eo9
DD6NszPjGzBljJ/EP/LyPUF/Z8bwYllEQCgSPyNnQAEySWl02oMjuS4skDrlBMNQabI32SrL2kqn
sBFhEfbdFC2dwGu7ccZ1lcz2PfEgTev4wGHD8IVFXHPPkwHeIJucy38QemxtTU1gRN5qqxL+be1V
9vRnKR13mgz/8ywkq/YVuZ7SyPYt9UyThVWT39m49BWCwlfK9tY3N/MHVT+EslN20iQLHk8JKqkR
31b/YAdEEQIc+hZayvk3tY2hWJrLfowS61wjHRrLYA7N0bkcycgc7jEpUDu8yOw1zS0b/WsVNQYc
+jztvtm6l+lxy7awB1qPxhuXJKT0EXtolt3d62JnB848P0Qzt+2aVUEy6UKHBDhNfoTXkYzWFRAX
V/+x6Ux5fvdEVPs/31A9NEUw7/xBAvP/TwwTqGiaCX6tpTaAX1WB4KxpVUkZbnDLdPtt780B040T
/hsfgO65n4pNDBECTwPE1fZ7NLwxHz3fljileNpOieN7vORO+Q2Yvxk4zgpLXBiiT9phTBJCcAOz
fef3wlI+k0Pk1cO9wwJQEpjimtayVOZfnpAOfgRBNw+kLi1ZH4p0rwlDDJrzkryWMgWa+fmwBwy1
oNAEA/6Jy3F62Bk6QWAivu0cB/z3MnjmvAURzNu3g5cBq0zVJNesGfJ4fdMYEi7J0w1kILfpAEfm
bs6U3ZjCgIS1o/KZZ59bV7iKzEA6Rl5EfYjLPHfYzuI8tj1f7ZxA6+n1k/5R1dPhSsDc9+oNDh/A
PxmN8JFTjQjfyivI7EJeTBp6EtTpvqaZ5zsMKbKg6iZj6+fpwVFGlYaTo0sgoqETw3OkZSZa1oKD
AM7GSMo5M2J9FRIFbzon9ThLAUnLYa8wxtfoWHbYdKqG++a3A6C33RtQ5lKqUzKgAfp19Yj90ugt
wFpBmm+0x3NWKNYl0CJI/jyLRy4dj0Rmw0b6BbquSO7XSs396SvP3Q4xqbEt/4nn4T8kIvjV3znT
hSoWfOjLnlY8+RbfeUHeNIkWvORpG5MkPLRs/KDpcrhMONo89l0fVNDk0AjITzW0VT86PbkFK0rT
n1dUzjS/nLUNNwOAchRdnXVstDzB8ebHV0Wgb0w7L3Nqnd1CTVG3P/2DdcObdg1UNKo9iQ938IHq
vNoT6a0oWRoI7diN7qXLPT1APmp47HmHQJWFNLKHiivmFATPrO6ddDOryatf8abhJ4MXUHULCTty
r/o8VTAPUlZV/2tzk2f3p4EmxGDIJs5zkiS6wbgskrCRVXmuhi2sRCN9uY9nQbgfYocWtKobSOHN
SD8bNxnZA7b8kdk4CMrqyS40Jg4kdYi9dLZ5kJKVb/67gfOclQiKfNILvmoAxEM9Ky8mFKbwSNAP
DCfxYSid+X+WeY/b4kVXmSD4wuouZyhyVpbmnnkX4Mxi0kcuMWOfUYSwIXgIV5PRrqPYy57rGrF1
SuXQeO+647ZzHbcYmpXmmhLlr3EeVbdFv11pFESV/c0RqPppDxLfkPqRN6hma80BOdzMtxzXUoW4
UzSkuZvhXom/UhouHMIWN63VJjirCUabCN5phbUByGMD0CERkgHgzqJbIMaOtL1hC+P0K1qzhKdH
qNBllqdyFz1Y3oAT7ep70NFUA3RjhiocmgXrhwSgF38u4DS8NEkvfvi2X/F79h5oIEp3lra6v/Yo
u5Ad/Emlkzra1hOMWURnYmYr210Uc3O7VtYIjPYBbgrKu7nIMc8GL48ujH5FfPExMjtDxCWehM0J
+zRtykPPnLqaVUBoArVTpvVZJ0DkpBXSn1lFAYH0lbrEo5bpBkTVjCHZSDCd41SSCeWHEv0cUXDa
7q/R8vfsoknLt2gGswbVHfjpWdr7BScHNe/1Ds8a+5BTl5LQCFpr4WMa9De8WziP74Gu3lQDd5AH
3ekuqBOrcKpAwarjg4V0zoU5pBDwga02sun6gRhMtUIF8TpBZEw5jUR9+1V5fDDm8mRLrzEB0IVq
6FtckA4fODpp/DfcnzPmDE2wyLJnBa0S3vnBcyzyx223xse4SbHqkgGX0gDwqT7RSUZBjtv5thYp
vO4y5dJyDj4TSggZvsxZBUAkIMJPG8jRBZImOoqOg11MVIp2bMi/uUwTjdiMxRoTXWpRTH4zbMVF
MN2kQcOVpFIEedd734+zuugxJho6rJ82Z79tvic2eGB/6iqRR5NyivE2UVUrZEO4W6NgnJr8EF3A
7pEK3+zL8UqbzoFEG6muc4naQNBQVclGtu8vtoCRrzophxpZK5H8z17fAnLiQjBl7ZCIU10Cxf+o
POC3YgCfxreDgB8uwS4tQf2ccMtkAES2QOPkE9y7KL1hdCrRT5EBcgORNhZzv8YhK47pmEsoW8Gt
BG3K+Cv578dt2LTMX/lO5cxDFsY4pqYzK42TULVqe7tMYTB7Ut4j8lq4yDNTteGku74CcKQY55cp
sa3D/BZOMF+bXoFaM+AiLfpp8zyPrWxnpaMHXrlrb8r3h2UZvmn4hBryEfV3KfS9wJZYyduMTLoY
00ZPAACCH62thLC3dUn1c3JguYE4ARm1g+zRE2f0K5fM6u2UfnpbN5w4nzTWSFMpt6ayzhr5Fw5h
hiaEnUXYtwrMHuRBakRbAU/c/QLh6pGzZGu/oeBzl9i8UPWrcoGatKBqBge0RwSK8ojsW79U+Jx7
Lqn2X0i6qSB+14ElNX5gB2ZX0zvmbgsGxH5TVm/9reRWTH6mwvS/NVl6b/LaTPeDJJNWzzpwFRf4
9gWIpBmFjOFFIFgoSF7Uyee3obBxWex9PlcYfzn/95PxX1+L8/gcimbiyU33xhHTmvBHlOVM/rkh
BuSTnYExiX93nLT8arQY6UrYWwIPczo7iacSMcueKs6sVaokPPGF38R40OMXA8gj9VezfpWcT3Wj
pVBruuzcGE4YRYH+7k9lAeHfv4u+zdMcvui3XsihEGt+HDQyetROdmp+MYZ2PRUBhnxnN5Lg1LCv
U1Awgplzm22msVsFWwbuDaycZB3Sjh+OlzbImNePimGL3WE+sgVsebm2AML7Dvg/mxSBWV9EbT3c
t9GvmcRaBWx4ob6niI0hCjOO1VEifZG048pEqKWt0Haifx2Eo8QZp7jch6bbwy7sWr4vGwYxQm+b
VBHofysAq780GYOJ7QLYfUd+NYF3F9Hg/xJsX0SCF9pwNdwazHpdnJOjJ0TUNZ0xADkN8nPJkFH1
yhqTpThtpOCAugzilqBlNwBSs2LL3fxRopJEV4c8XzoEHxTX8CL/RBjBLX8ulubyym1fRLhvUFeX
vQegdLdBQ8JIabN4bqjXr5KE3PM3rTL7XXfZ7IwDQnQxVovKgKsuih93wMpYnTDH0uVpl75c06tI
5+l0TBZr6v0iqF9O4pRpaDf7rS43hr/b86zZ7DP/PxDIqtEXJSGh/0XHyAjXKitBaUDMWoHfDFbe
N8N8u3TiQMIeY1W91maupSdAlZtrdn0phfuSFN61Fw7FDSfcRNjO/tWarpbRmvGK5eLAXfD7XQ9Y
XmWoJ8KY46IRgC1kxd98hoEbOt29nd0d+gKG8SCGuRnr2OSxy+uwu8wmCtJ/5GXtV4/PNAAbNDez
Wm1WxLoJbm154tH5WBXwxY6jej5hbSish8Spl8APw1c7WrZqH2kdZfyb3vh3ab9qrwLSIYq1zr8R
Eh+JsvA9pOyPF9BnHpCbYbowxlNcDAodB/y88gXkNUAHy/JC2oZ3hdxfO8u26pPQB7sqLUZZ29cI
kgcPmemfYgwPnLr/B5r2aAFJrjQL6QDqec/Ubp7V6hShIbsBD4W0jJw/Hl9nTkliGMbRMRp0xtq2
9Hkyo0123TgIDP7u528eAwpY6qa1tl/TSCEovpFJpGFZdsH4RpTo9NACnOLAETDA/ywMosP8xEH1
7PxUmAUeSJaBSruf2wu6ET4le6j173UCium6pWYv8IVn3+p7fFibrYF4RHJB0ahinNOWXLQSAFB2
voTaahqDTAYpCkXEBofErnl1G+LpkmVu9Yu/+d8PL81++ufHXJbCHi27iuhR68zp/X8M8G+QXnmI
pCBy46ZyDXs9h9NQ0o4FEg7AcUP1Nm6FmuiJgziiEXB7OdznNdiGLXdYOtF/7QNWiA6lpcnxXxC9
WW5AjG3VNKJeESo6LNCHMoqe3b5KI9VDYfegK75c1xHwsk+2DYak0vQmJsba1hHruh0A2LLcJSpX
PCxXu7qS++3Noq8ds41wv1wQak/fW7VkkasFJT5bbJRNMlXIbNt7tKzvtl/B2v9JESPRQ7kGbcfU
dSo6LFNsyWphjjCoPMB0zPpUBS1ocOElMvR4LljmsVX115TczT32XuumgPNwWuubQzbWOaCNzJPq
cYppnZ0474y2dSDGqHC8cNk4y4OiQE8jt8wjQUIaZpvUYZlzCIWoCUZV9AGuTtfdqkUesgBP3+4q
ru30CA7HyojaeMfORPzeVtnGDflaogUYEMVi3HCKBIK1lnkhP7nsATDNk3xZ7yg6gzG9hhDmivnj
1aSXclWaDkkr6FAbiOZc5ELQhQbZAQzdE6TBwnfsyEO/V21W5LER69VE++h5aBsa+azf1ewTwp50
FhxHMjUxG5KebTp8RQqkzXe59Ci91eHmEmoLGhQ8TwChfeMYY/59JacEN8UuvQFZ6rKKuIwOtnsn
QP9unM5xDLwxLlhzbu2DT3dypADj1ZFVKv5LehuihgIZV/SMRcYbPIkebfoYYoeqmy0z8YVLwEvt
6odz60d6vyWWYIaohLFdrt0PN6nKlK+lmWyImsczZVHT26Q/JAJjOMun+kPdsq0H3mt9O6MoW1Wq
B5VSK47NnNwnXBiZYAqkUYVDF3DKBETI43Ag8C+3wC+26/b/SP4mlj5QMngrGNkZC0hP5A74PPdN
m7Lw6VDpvUHFI7O8hlRgaN3UzBmJdq2q+6bJZcmQLTY0WkZKXNklf7L5i9a0EyjV9T/LJvHoFyIu
kyCLbNo2Ck+Qc3nLqflIUhnC3lopXbA4xIGu3NmffxzPvYF98qZFuIxI7Zy6OuesEZutLNjE9fZ3
2bmpXMIHKO5Q2q6VaxEw1TCt4qMk0QVZFuS/4QPy5PpUIsDYlGZnJickfYyFJau+h37VY5y4Cs8J
EatbvY19gz83o6uXAj5H5eoNzREi1onpKpXJm72KsmBDfgBl9+AzSA2ifzZ7dAiaSV1qJiIoBIvP
PryNSpnqzubaVXUL8WuSRNC+ylh0+tlZmcZdfByYvPcOG7aa8MB9EuEoloYkcxW4jtnSR19/bLO1
XTLnCydiYknoxdYOqUaqwam7gtxUgbMx5u3Osz5uYxYDboRb7SEICiGvelmUxDsFe3GrJRn37ThX
EoeOHqUll05unoReZEp4dgMMIXB0HNCLA8xc9k/41d7V01VRth/CYwyBqO/PZTzOdKnofBdUhO+B
G4II8+darKeLzxK6bpd5lkJ+pmAdv5GoJ1CPnQ+WBfVZFt00JN9CnmiZ2RYa/3EMubWso/9/anYD
2S7Q+rBk4uYcKaV7LbmED65xJPspV+aqKaIJmaIxJvyoZW6oBRrB4TR6nhZoF24HPGv+6BlWU8e1
p8VkXZ3QwRPVNh6z1EEMuu5wA1dQYbmwa1hdNLmDqP+5HXHaytAVL+sWDnwy/GogxM8HZE/XU0F9
KLkHdiWqchxz9BE7iEfk8kojH+lcvp5WlF5b1QCVlv65Gwjd04mWaNqnWcrxaVLezec4i2V+gIMK
VyZmEYYa/Zp3eT4bxMj816keXfV+7jR3N3K7jCkOVM7/RvDJg1rtG4Z27giCsGkxKsTEvb7uEym0
JGfWngnBkS+zGC5G2FYWL9GFP2BRiR9r8dm2o18ImTpCo+7V45SkrAs3pdMb/ypWcDdus5FWkXEW
S96iYqdTpdoglCWZFDYQ3dS+vChl9PByOpOpOAgcHoP30gMmyTMUCjB2nTmTxleORhCodoOeVVAG
RCElUMF0wOYapKRA5otn9zJRP5FgPBOGhrWCZsLchuBmLcT9vc/C/YKPyCZP0IiOwdSl1qsB/Ap0
YISgjLQfBB7OY0wHkZyp3ncb7JTXG+F3aS2m0EBr8Xal0lzqSgf/yZGoy34ZRCAwr9hhU1YugZm9
CbNO1E8KQ0VhhPt0SfA3ng10ZuN0RCBP0KGHdR3uX/TbJBUJ9KJXcimsDAyVwmSphdp465hXULxJ
k8enbEZl1gijLJ2+fTV9Kvu+9MbczdYMYmfg3PwfIXXqFqiXhrB6bPf9/zIvws5qFtCxYMdSf2HS
ODqyaWffldWipQrCBavzrd93/LeRTPUXvi52chT2dYDSZ/3Euq+B09IQh+kK0UsrYlt+QXTWlVny
pjllbzP71irDdzESnxEAWlg+7pqEDMIfKm76vXPeCHZ8XaihTA07njtRkUTGNXza4/0vJ7WI98w+
Sq8QKCn3zbb4CUX3YWKz9sFbP7cbDRDWNusp2VfTBBpB2k4HvQwruZupu3oGeVCJmNwGDps6Qabi
XqavnWLiZQ7u+ywaPSD/kZXSseB94MfEZQ5WlaLGUL5z+0kf+YufeZ0WdyTc9F4TsaIM1+4IU/Xz
CJ2OTVtRRDom0VTNUkJtu2+vH9wqSRfKqSgmiY8tmD+P1wSECEkMmpiWl3p94uwz48+Nnpq0AeEa
j76WxPZOXHYstgoxJAIPpqlIYXAZ9NKt8NkN5brgJfc52ghTQSW+lptR8VDgzX5EZuwAFcEa2MEW
yBrKX8dJOQnQ56QvbsPpeo8S1Bce0geBruRZe9IHWMa6IKRoUjEWCGVoSh6LI+ljjFCq0z2QX0Qb
dv+AqXv+5pBqlkgTFqR0qjBZMX4PLg7gwV7twrax6UPdR+oSZ7dfqwajRrdED3rCVPRzRAp/T2b+
OpcfPkRJcfak3uq/Z+EJ2dXk42rn19zQA06QBA3XY5ZNkQPb8SxUng2uk7fAO5JBJIN5kIqIUGeM
GLZS0sOjDdcxuxDvqSnfF87qQCXijyIUv0eT2GM2tZkAEM76qV81bw+Drs9xWpK4Qhi9VFcR6jbB
n1njfvrqulNgWVAMrFcDTVnIvLe0rSkLVcmFi7xjWdsMilbR0hbh9+HbZFBJtT3uNAWKqU/HxsKU
UyoGkXl3wABUVo4HNv2J+bMkfRo/cXEtZScMYux/SiOSAseKwlZaYHZRVG9E3IAHnIFr4QV6yX8d
wm9LwEwMhHIBSe78wyECO+LTmXN7xYyO9YoFjRWUCcxSnTyXVopXkNPYLxBgbzCxmXo+I4Mepb2f
ydcusIshJqybZHWTvWhwtSDl19/vVeb+McPM21bzlwwR85LqXGf3AVgXvJisNyfqUHlYbfgFHDwI
Cnw+LqCIE4CKxv4SKqdpPuy6kXjfqymW50KdUD0NjwH446Zj00/Vii+UEERTqGjDv550eGAptZWF
L1SJLD+5Ti2xyYBaD8gy8wIzPZUpcQ7xHreFAoN11t2WF4ygBP8pqwYwbQ0IwqNPKs9I/5qlrngn
MeEnzUwEeZAqDzX8HED9nUSBwjztxyyUGn3srFoccmJId5jpeoWIeKJHnKc+Lnl/cyhiX5cfUFEO
loDP7GPYBlTQKIOwqDp+93qRDOb8ZA4s+E60/AkE2a9f0MiLhhsbit90snxQhx+tTeguyOYhNuW+
hvAlTeBpNeUCGSC9Nqkn7sJF5bPWZpUb4vPEufxrRvXFtHLUd+hAg5yMZVpyMrQ022HuxUcjLlzB
kUHv8nMyeX1K3no125EPYqNR91GEWmOEki6veGJrIQdea0Uww3rgfYKXoRumY7Y+wL1qer+vktjZ
Bam9A8FKQymJre87/9Ybc6CNKca3OtIsjtPDjcj5YFNdtxSeSWFc8uzoo3mr3ZZM7oXP+sbbMTVo
iVO3E1Y8ZXwEoqkwQm+NhwavRZ3ABjlKQuie3iXi5bazqLjNkBawfoJadTOJ0eYpgNjhQPMVp3OM
62RG+DB1NcfaleH6ZEz06MigkpTSZkmc3AO3d/oJdl8U75f4jTeqVaV5KNKVij6GiVcUJJZAy0zs
QBC+iK9MoH5Ric5KpJY9MTtRZTJYZyPMknGk3Blxnz3KJQPewwA6jaDgB302hBz4qwzmJXwDFaKy
tBprCzmJQ7V0ebyCqtbIkxuFdBt0WIVvx4KNHwtyA8z9p2uDh5GkW24YyDYPIiLZT3jjphqM9u39
Rk96oSKU7fW1arOh314noPXWrdswMjUN3gdng/cvwmoMo/10rG3nlqJJ3XesQJgqaq03fpsGWFKr
K1fBpbJ7IX5MfNWk4jmJZzTCjdtLJcclWo70F14P86IvK4lodQBZYXS6qdlcdSFY2kTR7xEqdnQR
j/zH6foMwfAs8pEHftODFsk/ADLAue9A1lhCcUo+4NTatOcaX5Us7HfXGt9A2fQkhNQqtOd+rOCi
lzEqSaB/gX52fMtEsDX40SiCqrAQibfWwX72ZyVa+RfYDbD78SkOjOfMEdfcRrSzHfCX9xh7BEBt
+xy4g9ydO+eghINgXshFhdoCCbwapsqYaKc3pLy17DCqQJmOQ2r/lB6kJ1uPBgKc6lREAtJqvNUQ
ytR5jdqL1RYkvVeBlcV2BGTPzl8ucX3xbF1k9Gskeekw/a5hdmtccyjaDisVUfYYHKPgWjxM3DpP
qpTPS3iL7YTZyTrasLXFO/XSzmLC9b2bkrt/Aj4VMFWDovYr/8fT7XT7Xs9SrkFxpXFtFYrzGDu3
c1R3/r5ENPCVRz/7vwpUv+c/mcDNQYDXOKSxP1qCBFRV+bFIX+JCXoOhGikecs9dCevHYabzCNss
k+e3Fz9E1lTC0ldpLTdeB6BP23/ouP7wkckMvxXmR7B5RmLA/m3/TE5m3nAxMwXE39K2ms4YRFEi
odJ6ST966yeckqMo2EhFBq5MW0/vaZJORBiG+dIiJoYReUo+lcsQ1rWVZQcCELt/R2ZTr72+4xro
NaqnuxcXHB2rdPj4kEVf7UO2Xr33r+gIHZhwduIv8P9cI+9sFMUxtQXfs5E8z8jnSa1WpIFj32Ko
48vzwAc20zDABVEUTdAiPBvFkha1FK6+TbvqqdO3mMgrRWpBl6ji08vggwcTd6axllYikN/DEfEN
Ybl7ZaESmuAaPBqLvhHs0LQR+JysC5heqkME0yfY80YgAgYwMngQiERrCuLqu24OreHvSvBW+6ZW
ZWy6W5lSyLYw8S3O4hbv7QqFNS/PPXomF+T6FNCs92fVc+p5Pbr0rgf4Jtv+AdFNFnQLVq7XhQU4
jwPXrDQO8vqEUWzUgIupcAblCiDoOQZl/UdiEOI2L4uNyQNYac1HDHFquZtdbpLU1Dsbpy1lnzjb
V+ANKkprHSyR4LpDVDfPEROuUfehxLm5eRopZPR5NS5PaSQdBJVuHyg/bY2Z8/gSIuWhBDFGls+L
8pKFE/1nY9admSk3Uvn006CsweLRvugOh1IsQhpbUN+9QGp1qgVk6w1JDJDVcfS3Ad2lMPwlYuP1
hXUbGCCJ8G+sw9XBOY/42t8Mj2MN/zs5SgrKdgb45qNHFKZdvyyHyNR4rnJOs8yZb+feW9NcDDHz
V1Ja0GsztPDnI7n8TKv+4qgiH55q+JPh+0XDyZWq5sWSAc8hJceOAZiGC9bgXrKryaIT5Bracmjo
GiSco/09lR4qQ6k1iVxjlWbnuSya/oxqQMTw0uhA/BGOOlPzTrCysw53J+N+gE4rZdSqRs9KCnt7
ubqNAqS2HdMRc3GTFMNPACnW4NdDDYv6MPhEyo7RtSedCFyVq0+O5ykNaf3CfI3iRcSQtxCMQQb1
ypcbRrjQ6L2fDutCtu5TdTwEt9he2u+goza+mHxJVKsIq7o9kQYMOEU9vmnFPD5zU6oGLRmGdZ2/
xHbg2VKzzC7D883e9bTY6d4V5jEaivBWuvxG7etDvy7vX9Ji3LWXDdR34o9PsO2ezMKeKlz9yrjb
aI51GgJrIyh1Ki7gFSptNogcQyxriAFCb6MO5nz1K/2crPp/jzptfyAtAi+b0/HI7XZXYlrgi5zL
QJm74fNMOQqcNjNzdTc77vbXPdxR9UVL+ilG1c9pEE7tVj78zYCFv7DZEX3YQAsMXPg6602wKq38
wL26JbAHHIeEQnQ/IqOxAjSz5WzkeBI793s7lxh5IzfwrXHsNWx0JMDJ3uhuGtJL1OlSzY/i2vbu
zZrwyOdn+C4Wbkfj87iZ/omqUuUFM76Uy7lZvzY8/woMjcLBCFoWh2pCdflzxCARJgFt/xLcG7HF
O2rhYbSx/dISfM0dqHqy1LlsPunRpVTz+vM7ZhOkoUab/4gr1SrGn0Q3oFQxcICAwuSkYkjlgPj3
amXDUn63ijZHuxSY0/0crGg/i1P8O+6ZrfDq+tm5O4KI+njaXtqAMF1mBmW6K1t9n0m+giS4S3O+
YKp6tFjiqSVdGz4itrdmV4xwSzunF7vLSlyDkoUsaNqE42dabGZFgqoq17331DzaqiXXRQHJWG9B
R+duVVgwpEPAcUq/fZFDMBlLalH8sNrq+srOA180XJ+L3hn9hfjfJCRMdZC0gMEJ1BAOsIfA/jX6
ljMF37WcvSWvdrc4UyqeE4Sf/PSzSa6Ts0Csdhm3lh6wv+hXAmkgr6kfetFHJuRrCWOOjRFo6JMs
H2zrNuyvvy9WBLZmnLHL1kWrY+zRe+0lJUQBbUKzaSwh+kVj8CJhHKE0pq9fxrB1N6wGWGTKA4vf
tUJakJty88VrQ5ld3WfFqfzFNOihe/6Xlx114/dYsnNucTGZIsQuIkk9Jz9fVY0wn0SIyCoZkxl/
rrHPKg6HGZcsbzuJtmUcGr9VK+SpZ6JSutkX3obXSaBCIwEL8tg+E5jaz74Y5ZyXE3Hl9BDj5lLL
abx1x4CoCuPHutuLROjDJZ5Td2+/bmJiVAwbNBNvlNN9+geBnxyNFU/XFH7ECavh7pZhlPXf6XAp
+6beyNHfZJuywNVyEN5xiZQrWv3DPeB8ClO6OTSzP0taMwUXT0NgLQoSp2IhoIUxjNgGtUQb/CzE
E2IMFjkUsMpMfXfHMCccGogmE6PCMJ1s2b6MCC4MMSwegUdwI77wvsryIHoo05SdvU83wDDgXWzq
EBBIm5TxO3vSL0zKTP3b4wiUREldnTbMDnXVN+hxbWJNiMSMYPQh9d/L43uEyYf75egoAneCIdNd
eCgZNfA8Vlg/317nMVSRh9OGkD0tBbduj/JiTsozfUmkITkhmAOHBi5iVx050Z9pJ7SAyhNrbzfd
V84kTXyo4C9vrAChkmvcVkr/6iLFyUjG3ms0t8UWHUI7oIG2hWY1t2h7ALGAINHqmpCmr1HEefnd
2uwwXb41629E2IAqiweSw+sXVRMBj/J2wthVPCDCz7lCvk+JQF9vY7aL8vitxC7fOdrFkbuUd8UB
xgxNvRk3isALIac83nhd0uTxmjzXebtz1VKcYsBnWaMM9rxnKk1SWHfs+Lm7GQDZ7EtxRYZjpnPN
NWjNHZwBW919KDwA4Ul8MP+ofm27DNAlpjbvOktRMFTUgCa0f31xcIYkQdb9+Oxsd4s+XlDuindQ
Uee249VCYc9VYlGJUhyXWWjEzIGinV0EdCM6X+EVv35ZxyYAwyN7D6pJDr3jWpvD2MwZXcosMGPX
Yru10K/saQgp29j06RBPlC8P0MR514ySE7pWAc3xR9tIR/Sl/mjHcfxK1mh1PwwGIHIJTZ7WgePM
CbEnmICAFI8xYZwtALSN9BgQb/rdT+dvfFM2lpf5UUEJQxyjVBYLA9TG1s7Mw1COStLVAuyUZs4t
T5QNMShMJl8qLhxY8LINcDiQQza0dIiSikKaFLtXHARMkpQGrZCCYMNvvr/65OalU0zD2saIuPdz
5jGmPcsMzOnJQE1nr6Y4j+k64/HVfOgbUvEik4IStVD9i0Ylq/kDP28NEtrSpMujO2PSxVXfXlar
kcgBXnnyVDQ0LKrhmR/dWVtPr3NL2WA56dYNbQSsMsjl0i+4M9mvoSekLHshid/McUsX9l4ndojh
WGtS95r8xAH+A5mCc7eUPajR3Ls1FMXCACatLi+KbQt6Q9Wk/7VH7p9m2os+MsSjxWjlzTClZdu4
DYVamMxW2OGzC7Sh7gMGtaJD3iF3hjKSFl2f1RopBjjXbk2DADDW4hO6UWpF/04rw3mMQwV3fiMN
4/mNzfxiwNXHsAeiOyJOpQ8Hus5gNQblgdtVTu/tg6lbjsbqM1Iqm65/n+1pxqQPtSKcQI5yP8Hq
mCxAE5JTW8zxy7nn3KrWhittD0MCoemgFiBStyXw4Mvmd/51/ZnQc2LfttPClKHNEhefD4hhSuLB
EelOrQ42biNc4dV6FJfZlru0rRlncI0Ga5nZ3N5csPYrU0LO5y7U8gAhaVHGVsxarbVInolrnN6R
S2SHr3R5lB3DA43x59MjEDslrj/yLE0MIdd+8nGqLhOctuaqUKxNE96zBxnAV9GRakqxqZv+rXYB
sa1++lPW80qcACmYEome2/KMA/oFrAibofZaueJzwOLoZAwbHaASRsmXr6DLCSMgck0Lg9C2Xvwk
wjw+YicU3evPmMEwCxHXCqecjKEm7WNRMnFpp3nbOSNIIj/mgTJQ2mbnlFNU9FvyQAyHbfXiC3T9
vDND6cvYNV627S51I55474ssvCFx6fmwCSs2X7zwETlEN/XhgJ5CMQ05iF0frkjIrL0wbUCjGjbJ
UpHxfeC0g66t/o84Gl3BIvxBWBteH/QfoW55fpQX+2ZT0KWT5jTDzMotRiDB4t2ZVAseOWSFRcTi
BT2mV7lIaeQQahWtHEP7Uiys9MucE8A/XIqloQ2Ti9qwj4PDdjOs06FVI2KwYgpE75UILYku3PpB
WPrIp+bzXGT5O7YF1naeqzbpZBNlliGd5pZUNj/So3IEno7VVZy0V0d33RCAQMXSzdwP7tAadI71
KOXccHVq6lHC3dl+xgRN0iNOlJJ+GKb5pND+MVUl5GObVAGR47VLyLoAP3t+ASFBAGKcFo3j+s4V
yGdi8mUN6XJnEY467KaK/rODrlMTLpioG0jionZ8pdszfuWeI3Iwca13GnfUxNrZFeFMlZr8SfMw
DScQL1qNTS/hkMXgImJ9iYKo4kD290aVynUDIHtxdwX+DVNPbkje6oNjC24n5i43T3Z1u0xJ4mLK
gGs4D5Ot0+/8f72oQizGWFCEueee2MEFPA5xGjmSquDEbEm0Lw7xv3eCyBd2zwe6G32PsaZTNyBL
juTBfCYLIANKFR0vMlELhrwB/rw69H5t1bsckysPYiA++u84AByoz/qQjXapI9C+iii4yxSxaKc2
/IhOVOdwh8zCd5hZ9rLddwviycDejIS0Wuue54FFcJ5OfE+4i2Z8nYjnzIfYdluNr9C+dBy5cvDX
N5DLQzD2fwbIUIjuPT7bHRFr9FjIcCTT0XIypSSSicnK5IOYdnjY+p56MuQcRT3wJ8eRxrHG7Pda
zO11OQ2zMUD2EaPZlOR1PZY8fMgB3idpmBnVN6WAH2Yj3DPhmHGJjiTBssbdcNDsLLPu7TyWnm0P
qQ8lZrleOKz2rvN0p7+RlgpuuWIHXD+8WkBG8jDArW2ZVudh4+2tW7OXQEpxMNbn2Wb55ZGgwNkZ
07P1UWdvR80Yoe5ypPxO/QD4pA3JLve98cp77peaM9NlcLj5znVImS05zb9Fm88u0yOeupcZI/5E
u6d/4TMhjRWg57Piio3hMgQxEi4Bixp+rQbpHl6n/7o+74RpbME24gDTvzUM2C7/74QeFDlpEx6j
NygRUxGp7rr6bgddXr/ed3FldBHzWlcJuq90z367dLOSUkUywPSaAOOCDcxkFh9Z6nvIYrJL70YI
7OREvZ2DEJtGsAHo1MeeZnZ8hqRzXzd9+kKxiIRBYb9jufj8RpK3yCpWsgUCDVJyeCURysDePtxJ
299Zpmxv2IUGHQN14PhbP7vclG9X7vI560nc3uzAxStARHfJqdvkz57chTFcR4/YtZxJCQH9j1Jg
RCS+J5U12LSgGua7mGUxNVhiZtna9aeBuTC9x15K9bEW6aa2+a836jBUeuAsEa9bcaMYCfMTZFUe
NIHCQin77u0oqyL9Khnsoy9HE9PdBOZVgg55xtmsTtCV2lEoK5Zwzu6/DpNdfIi7gI7F+GHLr5gO
0YAA+uu3uCoNoCsg8qDQZrStVBrhEiZERhCfwPgKORpTdEvS/2eHo6zMEsPx3oZC87HnYddB05o+
knvS/KNm9H1BWqfKpZDleTcmoOG653gnaMj89iwowzOewgJqVshQbrhDOVEF8pPMFdkTEajHYz3x
+uEIcwEBgS4p7VrBlLdNJwRUB8k5VVGbTczp6kfiJrvCwUUtP6ECdhwRoYeiGRMLKbY/05gQlNWE
cHnx6D8FIt+9zaGo/RJWonPtsNljKilMe8DJbpVa3Saicwp312V/OErB7Jr32SpHLX3VN4sriFcd
5oB8acaKfOENNgtVhJQ/HezmaFwW14bjhBxpbieHrHPybEaq7ju3svK4eJezHFBe5mpN6wsktTlH
ZoOF4nDrzlEiP5gUxpHRCoeQwyQbhHz0VAh9ze6YDMkOe2h05RHwMBEAOv+Zd+1Jx3k7y5czYwcP
PkFI7p4/TGrWSwAUexJ8c6kMr3zK2YADjwwfxyAVymxakp84pH0a2vMPuO4t61eUn8vKbj/XPTI2
NchAtz02Fi8kr8WHjIqDiNpi9f7bhFWvnHu4pQdagsNGy3W54D7aG6L34ONzMzGhqGEK6WME4/L6
LGb+2vFXwk7HnH1oJxbflVNJtwbwkKMu/ch6huaTlnxPb0v/XHgFU5savEMcC1R/bnGaVY6bu9Jh
SIh4BbH3hPzCcWgp+w+jfeso7YPVvk8QLbPN9GuyKKrdJuOUD0XuVPKuL+9Z8tckhV17HnDCc3I2
P3lpoIZn0pqik/KPwny8Nnnj1LoZTVcJk5EOoBLUNNIFbaRalRp9h9h80LiJCL/JbknppKHJMGh5
bcztwOcRjqZVkjxddP3MfeUsmdfui1zic/LYIVG9gumxuxX0ycTW+qlrM3+u2i+QzrX80lsy2K/u
gh/omiJA2PjCVuQEmFlW2/b0sUldG785CfWi6/1S/BORFMTTmlSpf7S8p/qr8NAljk3rwIsxdUeG
z8qJ8BEoCWOm6lvlGq37OtDtrB1AS938pOwUQ9P5Z6oYrVsaOipP+xwur6DAnXtMZq/kkLWSi2dL
HRwTVYLqIGn3WKG+jRSu4U+BKqwFPhcoCSkDMZJItcsE1psct7MvpiclSIgA2xePZQYFo0mtmvge
OexS9tIKhSQNbuWA5iKqH9CIAEmNhwBlEudTHQikCx4v8mZtqGC1u9tGnPnRaiNOKic+Epyjt1cR
m6ghf+LSh2X70J+p5fulvYGURSK6gTwtgZesMIWLITCpK0sdpzG6GpyPWge/IVG7/t234MyBnZ5/
PCvjH5UQ/GOqHlX+SyunDBzLO+lY7Oz98IckgrrmgkWd0qGHWBv0rZHrLLEFaeTyE6d0S+pxAlTM
zggWwY+Oz1+vZlEQVCb/ZLOAhEfVfrBwFbHUdDcR9bM3D6LozZC6G2D9usQmXp6cDNAH3oruACO0
qEBem1J8MSltLYqVsNQv8UzQssPiHFBg9Lxkm/40fha+6ByryV8eqYUG4Iphikrn8AijJJ5GioyJ
QgkkHGFyl1skYpIwrgxXqHv+Z/L6vkPn/OQ54HTka/02syyLqt6qLH6KvQVCJZES3F9/F2yskBuJ
IgXYbY7s5VgnedWr1EbTv9Pr4r2twTSySVKEKZD5E7sK8AFNbjj42YqR+U4Wf9sadkDiMTkanuGy
6gMY7zxMusGyjHsgH2+5Bij6+s9id23ks9WcHW6oigpN0ZLS1dRY8wM2C4yErIsGdNjt1y0raXh3
az+x3dkC/WURHDlnGW2YcSURbLaJy8NraUKHX89/VEPuU2IGfiYmyyRfgHALvOiv6NDWnD3It/U1
F/zDtu4FdpaZ7Q0n+PyhuXFoALBozEks+oeZX2dtjXh6ppguuAfWmUJsSRyVDVPbfl376NJXBowA
HvQ1a2amZDVwj9dlv24m79c1LtQk7XWC6nttUaOGMgzX09Txoo58sZkHnQu/9NQ8Y6kga+ZW/c2u
ksfuZKiboiTvol3q5IDucHCSB93OBc4Ie4dE1xU3oMU7UcVAVK87cvdQdlnm4gpQvTXHps40DOIj
b9aa1rC9vrDc1B+l5VOzJaRabjSkMTFyOXXVtmuC9BcV365Dgoxs2dekcq/ytxdbXSf70t9Chu9+
32y6TyG/MmF/lXt8/VCjGxL6k3XPrSwHIA31W7PK4/KszrV+Q6YVlUmPSqpCmw7gheup1yQUnzkp
bHJLibh6ckovdpI++GB+WvevhKloW9FH83sU97tZPwkSP1jtBkizGiL4vp6U+bWIPSpAxJmnOyUn
euqNL2tKiSyy/CL4s59JmmTBf1g/kmrlkK46B6pal051sC2IFVXFSO26F5JlJj3ZRpKTs/p+LBjB
bpXjye2FlE6C/DPgqSVZCJQEtRgiyDV4+VgCzBG4YDr0Dr6TePP3U2FDUeCvBdohkVXTAoIAktVZ
VM7Wjef1i9EUiDA+tsyySQUUPfAsvr0gZtX3q3Oe+kyW/dPiOH/TG9p/wSSEaMYU6CovnYZDr0H/
Cp+gPHHBX70W+Sjq1lKkNy8TjqE7QuMRUg76yc+qUHKmoyZYljwdT4qlwl4+u36L8GcevcAu78sU
JaiISC3tqQUatTVLZJ8PRHJFdhx8KFU1KqMsMkTMkk3N5ECZUdXECNI/Ez8EHVd9cy6BOJlNFGC/
KCfVPkQVzC1dRCO9itOi44/8rOB3fnFFAP6zwyo7cNibMOPlEUxA+xyFxtu5LqOZMDtxUKKNDgMo
pHLhkdzg81QkEXcQ+mW3zi3LTM8qhD0graLKc7CMtd2h3d/Hy59B2EJZskvI5c7D/hRY83GeXU2f
lMEtgLK0aoEOZYlaa0qzzAccwwe+VH5fFdMXAUYb4Zd71yvMfHwN3CUezbiiR7no2i/l2OGjrigx
eceRfBuf7XDIDwal4oE6JfD7DwNG3a/+zLiqxz0uh8yKieb2riIzf2oipC5IjrFyPzhXAwZoOCXb
CS6cAYxbwXEyjd83mPMJypQ1KzWLTeBkr8ie/QyA+LisILZMBv7RJE/k7Sb3nOsfEHokC6LGvlJs
wH2arbssmocJfKGI7taOAcolH9z+oIyjYFrZfIr8ByugZiX6oUJr4++LU035kAph7JRjokONgHL1
51NtrnodWkJ5hSWfUo3hbxPUQ2v+WLgA/og8MMIM7iDd3GJgx+ID1qTGW3dQOR91pGWAKR9S2jwL
PbbKHXZrAQ7D0i0/Z1diqYQBiWvn4lC0xx9k3mXIj2vjiv7BaLJYwc1iPxn0Kpm2MceyKSQ01apc
3NVoezdNkv8ahCy0oHQk2xTDaJMdySzxNj0i/C7j4AtBBWS+Xim6Cg5xgTKdOosD5OHFpnwlOyWb
rIdxqNL63H2eQGJggeeCKpYtwJLmjgUMd4WQ6mJkEmJDc5/fS3RSBRDuhb7NLZ28b2HDG4xP1i0d
yeITMiRcC+6+anD6t8Wl/GIkHFI31uGwmYIJq8QkbMm5oI6K+FN5b9Q6HGRM/K55PKmCvSLYrd33
rb0oVhbGufrlKjs+EqxjXQLnF5TB2Kr63Klxre8D68u/q7BYjhlYfV4DR5dXYninKVK0ZEgWEcr7
J5sXQuvRk+j9t2Wve4FOQVjJB2WKnAqCA32hNefV7KrmFGpOsCx2JwO1VSfFOhrT1D3KVBp5BRtJ
ao+uxc8kvDSYrDgXDdrIWDGzFSyN8ZhHAUxlz2AfI2OpMbEVjNGGr6MhEAS6uY4F0B+1rPxHDOEO
K3lDWKN75VTaTw051h2BfIuscace/7V4GJv7r8mvTVM9mJMBT2XfTPaxytrYV8eXaDYebh4aTD15
u08ujHjHruyl4PqVilZ5O/kwRfzltY9qbjG5lfT9yTYoBy3FE1HFgSNTUbkSzvTCWjZbeak1n7WW
v4+kfh2mAWdQAPVU7Qelbl1hdh6fa6tphlEhR8cnxLXQHWuHCMW1qNZE5zgb9VrLzYTvonyS23DW
y3hz3RmShoCFBof8wSJQLVuVEe9228cjQVU2CzoXiiitcAB8KuLXdP/bidkFKkk18VwnXS+6kCB8
URpEq9ouduEVEokRrV6H/MquGq/gfhqgwn3c0Cu37v5qgNFVtILd2hL36ocyvP6jNj6ynlf1pql7
jLLikzSK9fEAf3l75yjlh10MZYEAo012Z8PXeVPnd/rGs6Aq0FS9ne7MJZlEeW1m2KXu7wW/6llY
6WoFgX+THfotEUPpDsiIMwI02eQbTJWITHEZ1YzQ8avIJGD2FoE/j69W3tCvRXEuUsQ155V3twFQ
9tIvRp7R7B+ccCvoJj7sJZzbFI0LdDwj42PKirUapvTCME5k3Cq2VIpNQtlIjLfxDfbikLHssWF3
CISAo8F1hUuC5jixoNcuZXQAfxBb/Inevz0Gsdi6wPcYTn6Cz3hvNQDGh6zn1Pc1ThmthziA3fxD
i5mxQUCsnkU882sI/2swNK7aq+9M0MAW0TOuMx1iFtSbyugQENMz7/05B93h+Oc2i4XEzYMyYqFG
sSZ9N3kYWaSyFGY0mkXOMrSKP998J8dn2AeO3YfGo0l/VfUIvaNp6yeEzHLwEEnSOGeu3AFsYGRC
sQDOg84BK1+6CN4L1ypnniEx7oqstKCr7a4DldTHxzT0fRjJThR3ogDI2aeJgSa5Aw4/8eLbDVZc
Xhuw1OFoTruVOsl9C20g8pm+pnecPzUhENHhX00jHFpOwsfSfVheFx7s635lGIe3Z+xpW8Yt55Tn
mWhGmXGXw1poqmw36es0y5xGCF7cPi93sQnl1Dvxmz2xgCZlEPk02oLmInE5RHsHR3WydvAAKOC2
nRkZDXm2vv9qRhtbq+QAcE6Nibx94y3AN2uJxVehF09zF7XZDN3/agS45+AWh9sS6FkrY/277bnC
6vTJgSbaDCLNtulC68MwUy1aAMO0BbOkbJ6u+ZvLDY8Jje+3GOnh0+82+xp5cwox/XuvF+i8iYd5
z4JQSd9B7E6duqYAvIcPb0gZ5sAh8rJV2K+xF0snJHuSGXjyP1M6gpzLHKZjR7uFPllkMYD3mAYN
ben4MUJrjlP/7QZ7p/WAqKaTeWxEMaPhlKew6jRhIUBEBnKkRt5WMupTFo8+gdmCNO8YI5ANS2z7
42fNulw4KnoSj4JsdDlxW778tNpfAPHyWTFtAHVBaLEZbyKdjgPcI9OrSfe0boGA6tJiwBBNoWRE
2ThZezEuvKUKjzuPw6vXc3gvUuuDn7K/FRe+wv/lh/Al6mF7H0tOhX6W5AEg5SDWW8Z41mYoQG2N
vujyHWZw3tU9aERJeJEnb3qUDnWUM2ohj+ohcdnLnUYWQMn5t0guSn40kq8CgpG0H23Z/ii/efvA
7+K/yXES/pffMtt06XQMOliNaIPVFNBM5ujVdkz+hK+Bp42aC9YvXaWFITyc4mpAgxPBXaBnD8VH
ptjNobgJblXJveNg8Pdg+aDkJLQ0FvLxebcGrO3cf3UjhAeSEP83E1X8BSIu5T4KXDhHssc0UMKQ
HCgsyW9HwGsFpo4Dca9twM5PhSsVt5zC0EJviDjgunb1xMjdCbX4wpHbo+YoRpHc/067MgdHK26e
N3hywNlkyGUcgkrjPIcTnh3WvnAtXe0CbMCz8SLvm5nyKDoO0xCaFqyaA8GO+d7TWczP4E0Obe6q
xCaOQEPHQPFocfcFMiMKnDKEaO55DqAPgS9Ae1gWoe+5KEMaOjZxM22jg7Gqc7GMZ0SoJLQCLdDS
vkG7sR6B/FUnDJHMe78reHpdyPPQrtWQaiFdNHKhL19CqmJGM1lDwiqWc968lYMhNbhJL5Xcwr1G
16qcK9NYZvjRitheDqfrWCbWNihy56GK5FznfqEZzuZ5h1et1nXBf0ik4TI6zYfDV+m6K8rpeKtq
AB6NfXKE+2joaaGR4MI5pbOaJAd/LIIXWLJfu2kEe1QV6AApaDEya6kQzHlncE7gr+j9yir+vyHb
6ovoEUn6rd7HlOd8YTyhazN9JUfUfFcHu+zPZELsY9/NsJtHrZpj54uatPoR9DRi1he3hG7tlSXy
OIjxfyqu+g7tkr+Yy+lE0DtGewUHI8GyO85zkcKdQBCW3czA/oJpWhUL9Nz6dsdCZ4sXpcLv66cH
ZxiZnQGsjz+rIse/YLvCH+NM76OXmEaglBClnUf1QBOV1+W1RMTb8WFcT8MCkYjYGYxV7ybYVzak
GMqwENqN/tkxpGat3EXd8DSkW7Ayhab7Ix5jOfD/Jctl3w7FEE2yyuqfxFIuJzqX09AdEn+7FIy7
6HdDZaXpkV1R2QVcZc9TPLi7UehnNfcRfEBdVx/SIIP8ZQu7xpHu9KZX/VeYgX48baG91adbImF4
9V+tGip8C2RrdZexSzN5N5hX1aBQu8zUnHxq76mIhF2DF7CrD7PoWo03sYj+EbuGvh5GFkTpIUEM
4HJP6N2S0UXX/2m2h+Z93IpY9WkmV2b5END3wqo+A8ZgVcM+lxGfsq8y2L2h6F1F3np0/nY3FgLy
SrHh3nivdn7ZpAEovrgl7f0dQBe3NMj8blsvmHn8yTSvcTNPhgQi0Tb5266xc6FQ2P/WGckHIWRu
olMnl0LOxtWGKbo0SPBGPVjwK+SdEzWDKGZY9zG459I1LfESuYpOy5WSZAactOdEBAuf5DWyPa1v
x8WtVG6r9XCaLrqRzgjCDUVHzkWmq/Ep9faVHwasFDvAYpe1+fE99XjqeufYenSU7hzU1D8mtxg8
0QtQ8f6wtxEnyZB2pSXTZI+sAqrlmOStPZKpJsOFvYASJmpzR/IaPFZ6Fu0Tx0aj5JBB/aD3i3u9
FQa8Q+yk7+dC6okCkHOEc9ZSLWth3jh8XGQDPtyV/DRi31B+FRbqZHvdHp8QltunKngo4WOvtP8z
hau+IXCV6uGzBlrEw3QvyiT6x/XvyLt3yKvLh0xG3qTG2XOu33QjYyNKbxXF67i94V/mZgLo2ME5
V8Ybqm+XZA8mb2KGJ7caULDwGHg0tZKStQC67xRxd8Sp/Uh4BSVeWrkbmJMkXK7kIBo5FCmFXXfF
qcEujyHz1IahNvTZux7dnZDRGzcBtj2dHinU4zEzVGOYIOKU5rKnhUvOYvPEzQdqTvCLoOStRy7V
8zP4RyKGPw97HolJtBGMepLyXZpjT1OTsQuK36Lnfc25lHfzb/jk/nRUOQNPgdK07UsK1hA00s8V
YJvhY/brpdSqsPziFLKZ1xO+oLY7pAmKv3UUt3H9wyT++vwufyL2DoVlOIEQwIfHU9bRIzDEejWE
oB5u1+CwvkmNrQqYTz9nqLvgrJmc7bxyOvOYLiPGzOjZgYbXHN/3mJs+PCwiFs/pJ/mAqAyIwQDc
E/ijJQJxzdfAgpazmSbVkH9p3GZefAnjarFNS73E3Xirtz2QjY/F7r77IL9gy7waPFaB4ptg/YWO
13xbEEY27R44hoopboH3+6boWuPXjV/iJJS8QjyRRVcoNdLel6NkgK9V6Them0+GkmuIFwhVj3Y9
XkPXk5WuUTN1wxIhOs3gBn0mV0lGzoVmoh4S7wcAG2BfbVKlmeNSpA9ge51t0+ZTBONPi23hYXDU
KGgNe3PkEELoIUYPk3yq1fsj2T1UoZd9Q5yAgGV2RRVqpl/fp4O3TxUA75UMet22hcXMYuKwEZ3Z
1P8LdxSS2EVOemgff8TlM1M8qE5kcYxK8fXVnqmcR3ul/1BE1jyatS/jw1f94FzAbeWcWLCxBoee
XNdIaJJptiaDewfAruIhCZpacI8kn2XSw3yoDeheRJMi4m+vWX/hC8zAv18Xz1ay1a/Z3D4hR9ec
0cHDCmWxUgtDXcEaORgKGVG+UilhD8opr2ULhGcAQ63Pl/vdgteR5mjn5/qF15cmkMpRYFBivRn3
icqpO7aCn7zYZ2WcskRtFPtldrPK0UG929ztelZch3TryH12V2oEMq0ufyK8YKqf01sPmA0an8vi
oOJBtx6ltd/fIr5Px9XpxQr6k19/RaHrEaZ8YKCc+7GzVdc/w7+Axut+mM8k9jj7/H3y9wypdjjo
mTYoUjyQcSbzKGWxZ9+h94nACJFyCkv7Xq3FNEoE+5Js+gmLWCYGuramZoNC1Bcd4LIHVogdsjfb
jMzpntWaejUKqghivmkXdjpg8ghV/IqfOLt3JyZSAk1aBF5pbR+rDkKeYjppWtLJuFWerqdSaaYl
VFX0PlUUHOeqQaWVR4ifVkJitAu1LjSA4ZoUWohiUcyzITfH324MATamUUrj+HSpLP1HFFvqonTE
btH+E3QSVUZnCvFqCa6r0u1YAUGAK7IeQbHhDz4ouygiFiur01z8VvCzEeAT6G4S2TJFqAjaY9u7
Slz1yROtgtnJ5xL+/c8Wg++I6nqkfwxHHB+XkZK6VUDFikANbTTwcvBzMYeYP0o+J0IfCv5H5N2x
zzLgvzkF55ySCofG2KTe+ePhCLnwJZPvpJrntP8IVtzNQpUzYrfB6Y1mlpPIUvsa6uwj+kotHzrb
Y8/gqvvF+FUxnmDXM8JtsEYa7HM3lYK4epVtbZrDKgylMsnvOq/NsrLBCyxzpAowWZ8RY+YqRLh7
BqI+bZg5QotZjHCDrZ3elZrDUq7yd2oM0B1gfRz+kV789dngLjgqmdKa/bKMt7slEqV621HD6fHj
6ePbvb4w8GBHHn6cz2GHk//vCzBAytarPZd43QPvn505DRcoMSRWnWXfs1Psceo3yqpo1gZmDZqS
j2Go+UIYN5/OWZYg8AttL2xtDtbveuwlca2eSZ/Ihwaf6r/BV0WXlUOndfHj1e0kRLQX7016hqvE
ObWBXVXTZopBeZHOAVhlmxW2POzcf3Qz5UXEGtbrRi0V3UegQsqwYdjoC3Yy9JiH+Gccxur96Au3
qjHlQf3p/k/ihpeq5l1x5V6M3xPC6fKFbUhNP/aYkHrzLlh+LxBIcdWXpI0t1ryqkvdssmgtgQ6w
IBg1hfn9r4/lI8W41ACEPJQqHpKEM34rNqJBWZEj2+eWjem8fEYEL7dhKYHEzKzbqSiHdcrYJWlm
1bGUDivRdfegPi8kDaJ/garDrsD4hJ8uywoFuC35kBIw2Z3LxGAVeiaVx2wbId2F0NBddcqrg0oP
AmzoTqLyUn2U+irkqkXHklCqYk+n3QFjP1g7M4B12TsigpRMD3VPMjv8pYvhLMSTktXzoKiUE350
sAoFVFAyRmeZ2VgrWSW1hEJwCUFNJEVhLYI+J9JAagO2n/9S3sOpEhWJfbICRHrX8AOUIL6r4P+L
mcYL0K1T+E92P5mYJPZejkuo0FO4x0nAp/5BesJJf60fCd2d/j5zhu/r/Jd/yutui0oA5BPQe7BW
h4mVIHeQfpqFj3Z7TaYc5GmfzDtppIa8VASwPVEN9qReIXpl1VSFFUMWN+L9lqSdxjbAwF7gf6eo
i+vVwkSrC1BivS1DMDgUw5Imb0dl3yE09MPLF+2nRoNXsl5LQrjYMlVaDapzNsQD5++6LZNyHc5Q
DpXwE1+7tOIGnoeMy1snwOg9cny3mgI1aPOLpMu7ekA33XPADlAhX2zYKLWHfR3vheivx0+NMN/Z
UAWPrWwoSuGZ3Kolqr/Nr902053i6ELZkAWquXd//lmOr2cO3WOBSDXRPvTrnMoxK09qUwPOqa2M
gT2a+Xay5a7B769vSMfr0GZcphklyOUsNQpBlRafVl8aECiyNhzk/77PQHvWyf6p5InHpPZaM36I
BR3ot+del9uo3akOzx6ZkRFtUyOLmgTENE3L/f05Az5CdpXjobsu7hxZpZFN4yrMeE9nxo6D+aXu
mGBRHd23dBhtXuErkE3wbZjdGYNW7Bers9Mi7CXnf0BVXDV6s0DZ7R9r5pt/+iBE3RLM3HtWPI1J
z+GoPNs/d7IsbTqsanL11X3aW+5BL0j2wh0tlhJ1fo6JEvje/MWWMLjdpn3XHEFEDh3n6rg6ug/j
ORSzS4qZtiMWgYwEQGrlKBub8zaSH6Lfd89U4/MmZ2gsNaF5ag/0Wg+oyCb7/NjjC40jaGRX5HWZ
/xzHW06d47noadN1vzMAXk9WUBSe5IGsJ9FPhau2RXLd2GjrGOkYKe1E57HzPq0sqg93VBgei+cT
4zatvQMugJbP1z2hCH9HtR3HpbRxkZADPWNvyjmGVhKjk8MlTFFOiqZw0StEqjrmkC4I6sLZr1TI
1nmdUrfarJFtHvO6CLo6uCkeIO8onfwI6hdd4JuzT873oxQWnt53RKU5zGsUPaajrKAhDQNyqGfA
LZGIAkA8hlkIwyJ+2nsSW8qOWcxOMM7R2KppRnfHbEO9/KBaS6Pusa/G2Ovj9eUbCxy34edBNLbk
V38yGKcoMEThoG7GjAe8fSUISavLrminNfWmkV6Nghrc3ZacZ1svyqdQ8gAsDfr0vlG/D2290zAx
hkg5acNMsus/rVv8HTIlQgNP5SRmT7Ekomyc0t9I9GRtrwkD5Qk3nku7+ZSBJc5v41pk4RkGu9Zz
F5dy24APn2RkPAlX4sAzfuQiZnbbJNCPAEo1e1UCx1nxWhd4TjmiWOuJufDsc/KDfPUi0IDhyw9V
50h3R40yJ0gc+XpM4fraRFJfwho0es1bRHAnsOE9XToF5Ga3lbR4/EaXiLFrt+MiirC1UOfhokoN
irlLNJGbYl3fyVIb1hskGEt7KMDaaV83S5lQNwl/QfzvMWeTvqauftjxR+ZNxcfh3/xLQPzac1tZ
6q/XQysYNYEVsnw/7Plv/VGKwlQH0jlQqG7fjwjGsYZ6GtTsRAWwi6U5NkvlLQaQiYq/D4opZ5Xi
vw52crMTBsJa95wglDZBb8pS3iStFTw2mavJAa2YWfLqEjkQt8jU5uxdt1M5UOQeKkESSQvcrzRp
evQNS+EMWcOMnvELmaU8woL/jqg96bKX2zw9CCR6PcALjSuMoxOVqPGEi8W/HDa5dMqGuE/TgUUy
I5NUR90GCm+luwzWTMJ+jIySTi3OUu+IX7mwgW/HvyQqqknNcFs3bp5opMo5MdtxytLk4JzHKHdC
+GHjjmGBips1nyIGsRL/ttTo8Ot8w02AFNWyZHo4z8UBiEePU/9+yLgBUToQrU18P3Qz0tjK8PPa
rm2nuDqzTTG3faFFngdWI5+GMPBvBC6y5wCiU6jx4Fv2Eg1b6MdOkVDuVYsVC1YeBj12jIZanxUv
2CYloAMsPWEHj1fzlNpqTaf3MUdjVtXE3DLjAf8ZrKEnE+ArxXjJbTnMxfn4XaH0ah9Q685IADo7
CjisGo2WjUV/R8ZloEnx3jkXP56WzLp3nhxBVsLU2zAfWck7mOTttyP+nzfUAoiqT+2s9DstL2Dw
QiHoQlw5oI0YN9yAOJ1x5YtMwYnQXUrmz15ExKFNm3dQO7sR7wpUHpRrJOAgY8pWOZ7PdJWAsygE
c7SUyLUGeTUlKk7ZEWZ96GOduq5qMQuEAaSvh9t6ITiMcWYEcnkBJ6lxKKUBqlx4+AorjpjLfvaa
Yfuztl07sbffFdJpc6PDAjys3E+phNA6tiZQp0O01QVdxv14w6CHjum7LjwhhKm+oWt93Iaozo6d
Ae6jeUAJ1YHcB2zI0Pgj2HjsW7f6xj8+wZ5dO8Pyj2IbRWe3F70OcLikcER/T4kVwJ2B5v1XFguy
Hqkea0fu/+WHsKbB5ARYjh3DKyi6ngruP25K6ZD5qd3005SyF6oRsYQwuOXMhiRWM5753OTrgn6d
fU/rszHuhP+3xSzRv7xkpdW7pM5S1SSMj6Ar+qDmY4mdbMBXHmP9J+HCupiGVahBNaRLaCQ9IBS2
c2lysEuOrYbnGCJF3vEvR3k+8GfzDXjJOtfK4dB5t5WB3CZrosF1SiKFKL0vDPR+xSfe5meyCY0/
NLk2Om033H2ORoC5aEXSJ6ZAXAjn4nXfT1i2m9oNfF1DlQCTd0+WHJPLQsaWwAjV5hEZJ9d6MF5J
sVWFVZULAO8Ll1T+MHos/1dUI821qWhsMaaBXVV9d/2HjrpM2Xm7QGnT5dZBZwSIsY0CzGHc16nh
fcX7pdKdv0o6zdtaivoLQRpOznmWqI6s/L3oUNMjDZTo5ydgtPtvjOON0z9A2U1mzRRXGI8e+s4R
Hoqm69yWHbLtYCkXRPd6NW0xgYHJVTGx6500ofcI/GjR3O8lJlSuvbCHW6b/j3JSiU7ovFlXsufx
gmclOTNSjIM2y4Nni2ZJnaPp2jTDTVVY+A0nTkrO8bzOJWGie9zQOz+4SK9xbcsRPO/7JlcW/JR4
r10ASZDcPLHsaYlTy3yUijk8EnwQano8Rrj8OukKVGgWfzCDg1qND23QpDihWH4a0Vc0UCeZX4ov
C0mVRKrn9PNoVZjiFSYOm7i27+oHQWVVWPlmfHjrIRuFEA+KgCdNraLd4pCFtqrKIsHivWx+PTmb
qlV8zVPi1ANpwjMx5p5J/5TIWHfOO6FYObrJRsHoCk7QD9G2c7OaJdCq07V1TiW1fJcMS8lplqQP
WNLrUKOooXwSO1jlLx5DDpKSKuGAzqOE6sXGWjnVWxWN2NgMosaWTL8jHz7TWWsYNBHmlfi5Jy5k
QaXU7P4mfDSmCbGIlqXmQSOdZC3IntY2babinG73g++WqOm85CF8ngvxrrY2AWWE6y4bKHmX8+PL
8yQv9JF4OKTz05JDnaZgzpswXF3BZPEzgvYbD1QaNI12c0Et1gMcEZ8WfLKkAAdzzvgMcv9ruftp
g3EKdVrWQoF3en9PQVPshylAvN8miCEg6H4y+17FrOOdTpaiUvgZjYEXpm8VeyeLIEZK7KUccrV8
Ug2YV4mZpD57XakQDJFEKU2k9K1QZGZlX9s8yk+LxJi6VHIymOuS38CstqylcVUKihPuKQh0Mc8B
rcQ7jSuxi1poAAO6pe36979GAEgttg72RRy/SDJ4fEWir8S5Q0CWp+tMXcBWJO9UR6gj6XZqXei2
w22GoxOIEvpx2EqooYaMKZejnfvZWPn0NXN2Cwa9eYC0Segig25LzWRSaNB9r9jXWoo7P3Xvrkk/
mN7iGmon7bqsabt+ci+Yht6DeMsB9a/ZWMNyDq7a4YwvlI5AoW41/+QLFeyRzO0ZKZYER9G3k8xH
QpZJMAd2s1w1OwcEHP67A5UtX5U3JSKTpZPfh5/3jgHSOxKmciZ0SJpsdOBumF3prdnBVCEBgAUm
B7Aaka62i/kaIHdFnQE9dcTktnwAOeHJwzszWkC9HXsInJVHutNe1GsTTfdvfGbl2Y98hmAcgZws
JHl626164ktnI0yB3vTQ5L/civaa1AtsHXFduy7RjHHVbTxj/keIRsJY7epOc78Irxz3dlk572x5
ZJsnttqeUUuGBkk/o3oVy1txAFIfLMHZBpxeLTMWN4lPehZSVUI2R2SsyPW7gssaGOduOZP814m4
+nW13l50EXBiiY4o13/03J1uzHaHR7q+4DhtSgd6J4fD7bhlaW368zq245yZ1lguAgh/ueSnXzQq
1VapvLQMgqd5+TwavIukHNk7WeAyEqepg8rh3vgAmUU42auMd6oRvat7GhouJxKLd4HxyVR5ZB/l
55m2rNud5ZWWoqJvWSCwTEzNrgk6iIh0afnlDfUDkt6KoeIDXoNOJMTdme031pi6oaIL0jyTCh9N
bgPPmDLKgoI29jb3yMXjJspPynlcG5O6lR3yTd8/cHbkQw34xk1oKxjOPbQx3oDljDDXQX+ToosD
0Ltt7ATNUNU5GO06uKfT
`pragma protect end_protected
