/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 307280)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPS7RKsNrJG6vRY21RDoLpZPtaLH86T8oxXnuLgYarUpoRy0InryH72+b9
yr2vxaOK8V5vxpiSz1hccrMuGg/euPIEFUn6YMxd2BaASByrzCnyotXpV/ggXdAaST49NpP+4UDa
V9vPHY8hctzbO3pJeM4j2SBTGCLJM7FzjhuN3y5+WgJjc0pC8yKlYctHOdFIKRPzegzQvfmx0ltL
05DBqrxHbwMxB/9Us1kSwWRRIEfkNWFCMUJCgdHljAOg4TIEl1WnLnuiNP0d6z1ripcY7zRQyKWv
gZhbO+UDesELW5oLsMKbXgS+y9OyRuscF5jnxmn9X/C/MdtGtSHQDOYgQcUJu/sSHtM7ZhhKPCwe
JmPlgXbNPoVbLDGZ0P5T2GVn+eq/8Wcen0WDUhliBR8iC/Hdyc4jy4eYzwbtZJvy3kE+cB9LaMx5
IUoXCaOXP3ltR2CBlOT0E3pDT3pWeCBdA3uLojv4AH6sRFelUjlMf8roSTwenmVAZY2hTtH/ApTU
iz5IAJtaLbraU5NWbue/Dk0YYPYzU7hWie/r+VQKgliUo6xjeJVXrFTdkJZYl7obvvPXoOUH6Zy+
ftb+KRHA70t16VD9xyN5XS/N8NfhmjJCaMfyibWu4EFSMlCVmNT+f8HQP3ZSCw0Wx7CDlx7C7r5F
07ONyLTt3Ug09GyfVtZP+9U9CjGmdEp3GvtqstT3GA+ONg7vKVlBtMzcph3l6kHmTWxoyITD9ea+
St2Eg13rH8BP/3dyDnsZiyd4m3wefN447OT5HVmuMW3y05GOW6hPTbYGE9ToJuvk6H/FuImwMqRJ
b7VIfDujTLv+iK8gNCbbhKZWhloLpnWj7/JNzjapjHK5odkcShdCOD1j7zjbwHqTUvTEFIV3uoba
WFeP20OaozwdbqV6JYgP+LSsQR86Op4EQftBJ7R9DYH/ct1Lj/hK3BAhQg4JGrRetI0BUXxnhDtL
JWTo+dQmKvu6x0zgOdxEVcbXaH43lQwab2xeVx2jQnQRrj9m1bt5ZUwXpbBKXtGOIWxNYZkfijmn
Jjs5ySRFdbYW6WBpiViUdpWhKdmWSiML7rSPTFe6H7nvXzNq3bvdbabF5ZgjFZxugKXJ8NklHKls
BtWMUaUGNzdE4BoKXpMBlpApLzQFy5rpoSwQ2iearvWTFOxDRt4cpeOZTTn1CiYtPQapLebtTOWK
GIWvDd6hwrZlLSj5twE4lpEFvc9e5c09pXWFr5VcQUIHUGRTYcm6iZMMJ4FY9Hk6IdgFFcrqs2Co
uKXgB66xiH5tHWEi+reUod/vlXGkpX5s2dwLkeOk9mD/T2acKWwa0EBGglN5Sc6GARSM8j5bcBqd
aH39yy476LtV2c2kS9VLI5fpkqiZLvs6eQxOB/+Jm2XoFASMYs/MXH72UbvDnXvoGYWxcoVM9IM7
ZMOuolTcx2oWKTYgKyIqV2F6+AmyFpUjZuCP2zqMD/areQw4D0hvC0GEpEvyCzI1+r1RqaOHHc9B
hkqTRN7LuGg/hFr10ZCl6PENhCdpp4h+B/cvPrI/u5q4s7xpCKeLScw7pj2NNLBWZVcLgvK7MCnl
20xd8vzOUfDx7i2DAvyIX81Kr8DbJs3cEFK0l8KdW326/jJZ4/cp/cRxwGIWM1Z40Du8nZkQ0/aT
+YbgJ72/pOh9XoPhrIc0nhMeWw0gULfCnu3VtnqQIv6+3FMbIeY5zmIVWN6+GGlf/noVeNxTOn+0
JE1HULbDlKUtk0+gZtGbNGUsTjpUK7XjCmclr0NpuWUPt9HqOp8vn5iHRE17i4gMUVzEuixY8XBQ
MHBlAC23ZduQgkokVcBVzHYBPusk7XvrqyRzysAOiiWiG1ZaenWCzQ90vJrL5p9Ax5x6v3U5JZCX
chv7p6D2aQ3gm8DLNfvNikRWm2BTcR4q8Ap9oTD0JpJIuAasS1Xazn9yBFxPXJc1qh5O/fSxzyga
7cpVJtco2moAVp6h9H8qjqOLWKMZUT9BMxGrbceiE1SO0H2C78n+fO2SspKfEsivlf7A4AXR/Xj2
axTVi8SKXcSVjo4YScOfpE5SY1hZ58r9xdQrwcIWTJ2WmttAQaX5tw+2jxpENUZsIFNLz+LMEEpr
yQ/nAPhpXgLiS/9A0oO6IL3z4d75d/3J1cLSQUxord4jsX/ghf8UaCoRNGFmL/1dnIzfCoPH76dD
wmiC2AreUL/POmo/zGUpnlsIRB1fPHVafnC2Ju9ASMRaDdG/QfUDsDUfkBRCzG7Mk0IPrX/OlGsL
maX4K9UJzXcQsWKp7ZPrTg77oQO8Ewqlej2qhk0Os2KBBLMxoHdlul/6+WuMVzGdAaLNUG+riP44
TNn0asMGF46Y5bw5mdyS1AX5GmmafyO64FEOKwXCmvORGSaGhJ/p5ZrzNxMPcZyi29znePbrCNxA
JbxEBrFpaYTSOC6dXBfrS33WuOjVUgUuwmpG+jKZJpOZ0Bh/FgI5p36SXs5YcR9wuKMH/21c53Oz
tJcoJY55am5t+mroV0Xu0JblNuH5kSWg6Jkkn5Zz5NHPe1QKLH+RZaKwRgKKUDcge8zjwTYPV+NS
zBPXvd0xFb1mJWFkyXKNXQfwpxoAPqTf6gP09CPnet7Eft1FYDpiQxcji9dMxV7nPughW2hHYkfi
NniqQa84vfKkATszM2fgujgNCpDgmE7HpbpB2ULWjKzj9m3UbzTZO4zkLgW7haHfTBobtXsUQiK3
l/HRgOXUtXR3mBMrH1wJIKIqENTc1/RAa/9OW7Y38z2ALj2q8GZr2PWPNyJu8rLcVbM6RovI2GLQ
rVOIwRGH4XznRWZZ6lbXCM3EmoU1XnqwDZgmD+uVe0M/LyBX8UJqyiavze5TRfhM99WNYwl6zezG
aGJhwBSb5mhfb/7OgzwexWGoOPlgmhcqxOJRVIoQa7PJKLJu1+1uQB0XL2dyw3R0TlWAN5IyZX+l
93KhMfZCKsNUiKh7VpEosMr9MbVX55Tw+gMZe4Byb4OG7icwnj1pKBTGhya9rrZwjZwIZuaaZMbw
12X/8kuNXKh20PfV7FxjkwZXDtz3EufB+JMHNEwUiOp7PqF1kXXogLXIACXuOqGjwHNRP31PbkNw
RY5LUpMb+vMx8+AgWD+jUqjLIS0isNvKl4iXs6yKnPCnt+qRcZhiQxc1n2rRZZSlTVRJaVAfhKhV
ir7yOIqv1o2NXHKdFFy8ptRrEVRiZOw9Jc13LXQ7K8/FIMMUeu6NEAtnpW92cYf0iMoGReDqZ/1Q
LUO8AcPfG597aTNPE5IgGA+ludhYhMSgEhpcBBxAhlcxfCFHY/tjXK7Ln+WeXj0ZdpHY7qL44bqx
E7DdeRtthIoljQGtyPdt2fFOB9hBuHLA+DX9/0GsKcBkRVs+TToYCn7kE8WdWVAhdvPOm1JrsNox
OkF0brZP78EgijCyk9bWSr6s1mt3NOO63n6Xe1ZApxfYahdgYeHI6tK2F35AZgy1IA5vtwqFVdON
y24RhCu47C/Mn7yLUSTk8f0n9i6bm15LrJagnH/xHXEjDwZ3H45WTJSHSDc5Q0LhKgW4kG/lYvqA
T3OOlZoj63gPaNYW3Zhxntw6mOCFQTkQLEhu1P/RxBGOxxl7UmJGYg+Wjs3SGpvj1YgUWuR4FyNR
NbqANhv01ag8jlQ4Wrfsi0gF9bV5+GZJKiCw3YuWlDWtH+FBccfTKmaMFYlsbHn0JBxzmDwIAoWZ
QjWpwutz+PIZPxSAHYBeFS8VXkQ+ExeOwPxsl3cCHyB3FT8EqqcWiwavAHUiDyPyMHDT2RT/BGOO
iDYJx0b9D2FNLVvQv5VP73afaAh0v80Hl1RtSqwMrvQo6R8n6wdMB8O3vv3nOsJ/yjhtjxFyEud2
IidcpFaO7jb6cHzZ8SfzgUmU1HYofQuNEL1f8sQ1+DGvbnum76hKcwbNdfSJ8m61+mo/nU79ztTO
dIagHP/vISQNO+jMFVGEZ+qot/U5/hn6ArbkUulWd3ejLCGqaPafyQd8jVqDLPT46fRDrgBOeSSs
JcB6ijRy0L09TpYDEMO3JdlHot0IQ+zwTd234YfXciFXDtB+K9hI62lZHJlbl6WpzQfuogkeFhw1
KB7NUuVX+4VuQMdRT/BRNQHu94vU0I0lPY9NkAy2H23FI8meQR2HW55CVdGAvdnRWhkBCD7Ke+zN
V5So/fkbEA7OIZuahX0Xd9U4Sxz3d66IZSkyjDHJ0PrlSNSl1QY0n93USHcFz1GfCgwwPGIwHzWh
cQJHq4wggdqZWdE7GOuK5oFRd5XPUSZ5GBXRfgYKyFXPx2GnehQXpQXP++ttQOR2imAw5T6U1H15
17S3fFLGz7XjEcjClnpZomekY6o41DbPBs80BmvAGSAMB3Bn+sx69O5onIaLb0ySBmHE6EmPbOlZ
06CX9Fk4Anc2ikEH1DqnHPyz6UUACHIkOLTZPnJY8ov/ZDLDoTcSx6mNz0u/RXFOTV7zvfb2iO0f
mj5+8KjnFpxpfGiSrPuBPSyPqadVABc740bt37ETbudxCU6O5e8mJ/89cbbJf2t3sgxz/C656jGK
pB9dgC5fEZLL9+zDI0bB6m52nrdvh9KA/LqtyU4KFU5pBckQVa9LZS2P1oYoDJiJ8cxEyUW+vRW/
wx5c8ng3W3nDW/Voc1ueW2Kh8f67AEDXQUCgXXfhx8fud5kJsxclqcjSNbQbJMlyDnsypfP6FJ6N
oxjT4hnFHKtcKlBEmBNmetBhdkyyAroDEEh3lsEYcOdxUzPtpilhE8mYSTKzyqaBI4yCS9YOJpQI
EQYG0nZ9EgCHogjfyB5Yx80BS1UfV+lHHD1LzNCWg10UT8P8Ac0uTaqUO7IXSP770VxikLII8EsF
qPgU9CGLHx5Lv6zzHK00b6GmLtjp4nF706oOtscsO/xGoYrp9VXuxLvuvE0E4qhR3xBtZZM9c/VS
/5ZkxkbUF9hHQo+xpS1WSXsCm7thpOdYnso53jg+T5JxZuF9tgukfxyBW9LaJjGElx7AsKvDINeG
KskuvvePGobmsSzrQVe/v9JCoPCZzpmSgBkm8JIIub6XvVuExI93WLXJv3KCS2Zj+ye9zJ1I6d+h
Ed4VX8Jt3r9fdJa73/LOYZHgogLVZ+tEZ+uw8oJK+QyHU8CBXHTbHkr9ejmDVMi83Q982U23xIAI
+sm5sq1yUphNtOZgUj6G/rI6P3ify7kMbR3RlvuCsj3LbOhUAFSJk2UUolr/kwmJH0sRnjtp+V5E
eTYoImsmboOO3hQyPh5F9Klb8CWPXYMUOenyx9KT3WStqLnqzl+OYij/rpVuaGOHqliuTzvasPu4
NA+Gw9LgaGluZlf03GUhhMnge4jiU9nQH0syXKfmW9W7pW2h64FRePjv4hAAWgT0kgtUewElo9WG
j1xeD+DxUCtaXH9ztrsZ07TebOU95RL3S2K6U53VSpmG3I85yKKfiSBCgqQZwBuMDnl7Y8P0jj/g
OhebKFRbye9GuI4rzD8CMlUz/Aod0LXeLyuUajelJMk9wZTXr0o3rYyjOKI8CLs/zlg8bPfAqoRq
0dlTvmIMYxekMLi5ykwfrPvgkxI/EMLMEWx+6DPJxoyrfHy9rZn3upR2acjBjec9VyaEzSB+2lWM
VQgbRM5WLQkh+RxQs0XEP6t9Y+QDxuNk2hLoi4n4dhfPT7IRuXYHgpqaZ4DWPguI96VnXmXexwyZ
VffZ854BhlO6sbNZrCjfPato3QL0o39E/vrZbVmcXjPOMkh0hmk1WZ+NkpPWI57AAaN8M9cHscXv
S3jAIsQWLhdM3o2TQRNBe3hkSPDj83M8z3e1euJmcifbK7H7u9RSuQMrraQ4hMShHKMjr5/tnuvA
eLEc1on0yCsEuTQia6PmK95+c9bIJGEwsrLehg7BHUeg/BWoAHNE7+zBPbztSGIqj58r26OygCih
kDL9ahqIiiMqIH08SrXLI4tkrbv/i9t8Z9jJXsJcRPYzM3EFPHfE3enrARtHs8lwTJ5fA039XFjg
v1Dgi0J6kRYptFT7ejgdV8SutwHrWyrEM6+KtpjcYD9CulpBPtOxpxHiBjJ4VC5zA1YfpdckQYXx
mh4Fu9nH7vNDQJyjzoucDO0fet//CycDXIPhb69ygaClx2cdJoE1VRUvPZp6bAb1ZRfpMk9ZZoJR
2mqBcXAoOZt+oWcDaBkFHPxGccXuqXMhKnn3c4haH9ei4x6oK04AwvHjUd05eD+ta93ZJuUhbf/L
UsgXt40Hr3klj0BSaK4HQdTn1Ja6168rvZmhbcl7CWMoR/VEGgyiLCERrGHx0NQoup8jKDiRGi1r
ZzmRIBGyThpO5QcOH7Vp5gd3sDSOWSHuQW9RSOvCVKCZQnp2MquWojjWxUaTMFV+vY683xackCP1
DJzoZ3X7LyTmnF4Qtv3LudfNnYNmNCXzFeHeR7/w+d+53UL9MHJ9iiwAW1T4lQYMcc6E0kUSBqCX
AhhFXbr9rXjYBAqvguW2dVkwFruB9L8MumEL7QIh1LUjb87mwumjmJVIZVCHALfvwtKcSDdrKqvH
f3jVyKU16YGXnKTb+N15fYHpQpx2dkSSQ3LtuXA/SqXdDOqSzo5nnE4gYpDKX+wAjHL60Y/FB+zC
iqbZKPsbiD0FzqdQVtEioXNW6egJl6dZcgrbaUNLjmzCw2IpizZ2bUq6Lob9P2UvwLr2ejxzchwn
80wEHRDRKD2UtO4O+zRZmG/+NbDbTVppDgp6Dv2aMKkr7oBFFVxuXKjXoIGXoojRBGcjo4ITeme4
GC9kUancONu2eBRn/ChJT5mhVik8xehX0iDosE0eFNgNZbAB0hKTSr03ruWksqmPOahDZ8J4aLIJ
YMkxdxXZBiOyBjfPB474ICy3GjHV4eJBsY0CzQB9Gd6IeZRb/DEyRUi6rLUK67c19S+zKV9XL3Zd
mJoZViv0s6+cQx6KV0qpsj5AMMt6hzk1wYPHGBV2EKyll9Fy7oyxZzS0jGN7+15GPCTAD8B6ob7D
PrDI6UyyyuTJFlDE1JAW+yNIXFNGMtz+m3nUw1h5tIZoFs/nvDLyH9N44ik9n5MRsJKwMjarxPqO
GyE1ltkdipRwkWz9rdPJOhVCB22LnkNTFLLhiB2GcOp4DI4yyZ3meDeGs/SkcVc/+n16Cim4CIFk
3VJ4CFDlFFqZQfEDsNwNhkgr8/0TKuSlU0CrfKap05exg+S9TWhTHornE9Icb+1nLoUOguhP+j4s
+OrnoCJgbiwGA6PMo75D/nO3VkJskB+1hDCS6ClpBMCIdLH4eMpRNklT82JBf2oXlzbqQB42j66U
1R8y+6qpQvOZY1oG0LpHVzVTPHMj59pINtNL6y1DHebfGegL0e/4YJi3l1njHhRyaZosXGgCNta4
W4urTmWz/v6tAC+A19FFiJhYpe4Dt757ntf1JrSiXoxphcpoYDSQimqyovCaFlwVEh+rJJuGTHlr
BLB9VjWk+rIx6/z7Qq1PQikRtzfGXKvVsiujjFgL7W6IlcaSimdYJipIF6PPT+9AUH0thhpHljzk
JYO64oUp3IWOkGpncMbwrqWMoVKE1jPigldagr1BU3wREpRDAo7dni+ufQK/MjRGIUOl3tQD6UAJ
wVv9PViPdLa537J+ev5ORFGSYFFFA6rHrFcYW9nKq2SJ3e0dMvdmIl3O3ZJs85el5dv7Qwhe4PZi
8fpAa29Gg6hdkSzUvcFMQ+371/6DWLvlQUynmymnLZsKUC156Lyr0mtBhW8TAsazDSQDxBXKh5DZ
FcyROdwUIHQN9f6lOPfaaJ2r5SzvVSG8BIhMKOeR9lhTHYS4kAg94/ns5oqfQ1x+zj7lW42QMkaY
SYuuhIYvrFqF0/958R9rhyfHKxGqbHzS3mmDXyFlA4Xr0vZLsmvaWI00CdTIXCOM0g1hWa6GZ2z4
7QQnFRUwUxlNJ+n6UtmoUCcV5gR3+CGAZPRCfTueJwySqo1UU5Q6d8kEChO9bgNl2/VTB/i01s2R
1MKOXrJsuzlmPlos2EQyttn1HCoLTycFB4uHn3iVenUiaBqyqyxA0Mc2aL7AQ/g2cGQa+RQ1T+7f
myF7SmU3Py691lQ2Q2iyO/qHQ/BJGuDnSQR8W70pfLoX2txVycGhIWCgcEm79JKHNnshOx3Iwnvg
UDXPqN7X4kqLuqRQgNmwP1448QRbggBmsu6X9JmsUJlcCbGSFFA3B1KQIHzmE1cqYDX/I8Q3qh7a
XCYM+bIqRZ2tJ+BSWofGliU4g4QgnhDrQUFdeONR2fVBiTV20qEwTv9y2TLErTm58is0CKYGPZ4w
efIIqkdFysrgGAetnLxetHHYX2kYVFQ0H0lIxQ/JKdfB9q8je46JHS5lUaf8gPUYJJMB8VY7xtE7
+ufFEN01ORuWpVT7WnvQOm3/j6D7JqIFRDIk0uM0Y0TLvCAP2dzuu6AjcoBZsQzdU/qMC9vcfuTj
/wZWQSvdYDZ/m3j0T9SijjKigTSD0eEEb1H9I2sMx3J1eIrmJRW0MAzASD25uLrbZlFqA2Yf/0PA
IHrjxQJK20GuJxeyWsoeLeyvgcTHez5/EZAUkmA6LeMq7ikCUJdq2AyQ9d4vC4fPACUSR3BKzBsu
+dtHOZjVyrUkgaI3iWA0nkzOkHAyfaJ8zckd+1Zfq5G+FSKElKsIRVLNj+8JJAI8bLC0rYueDLt1
82ArJd9kAHZsij03gUUsI80OT3Cv+li8+JDoFWpmGT8krj4ChrBPTj3ok/BPDR/EPiQlPTKHuXYk
Jyd+33f6w8raExnezM+XN2tgbYqBhBWN3YITudiRD5YCQTrK6RkRBOURTdoNUPqvF80OM0arKO73
H/BMOUulSw67Tun/06Ym5D8F0svSclqWU0TVybD82rqMM962h8gkK9M4o/84IC/U+OknBS3eX9wL
fLOL6b+EI+HKte3mAukn62HX+k8AXBPkzzTNz1Bbo+p+VSeBb3hFrsUIuYFDQWRTmHjstMrayyvb
uvi6RCnkNP/v6/9lK3QD9QJxvFQmlW9crU0fdmw/Id/xksOiq9jDizg6VQ1FkE/Cw7r+8FoSaAGe
k99cHw2rrnUTsV8BbC3mDZ93L+yDPqBgaiSqyhBpTzlbtT6XLSLRrcn9Nh9vQtTL1FC+o4Ag/oPs
ITBW6ovmbAppm87+8fQTUyxsxZdhXmg0lsmktj7rl+2nr7ZOS5lP0Q15/SuXujG2TsuNpfige7SP
v/8tJzD13Yi45Mv9+Voy2ShUIAvnWGSH4rqbsOvgRNg57MTZ+lhA+ZuD6OBctuA+NxPM/vDT3yjc
HeGVMsxvHBetecVk2PeWE/tM2A3zO+uyGF6rx5F8XpZ+5cz9uYA2ND1Yg+SpfufTbLiRdEV6/5Sy
Ok2aXyFSTBWDS5BYPdRexzYsbBrmQhj68Upwu0fcdQBzcaRvSjA7R/CHcRakWP2pOfuquq3+d++v
HsJgVAvqn2qRhzVyVdymcDWzvwExOtLq4vQACMrp2zNbNqvpaGPZIYBPmgJWefoWPzcqU5R/Ztha
8k1DJ1kr2b7VEfcfVhchwyMDjx4BiP5HgaVEvGfdPUanIj6zLc6VG21YZ7kPSKxb12zLYf69Skdp
NgW74KtBhI4D6tSIjfpn3vLw5TcZWZfBMxAbnj3r22H+7tBz05gPlqVacduT6/iMBi8rYTPS43bG
qQVz7iwc4iIasjVydqZszMsF27sPSpTHMzRlRbSZLI8lHC7PXwNoC9ceYzWysaovWUw9I+Zbb7un
NJj0X7BkafoEb6cgQA10vUHooZ6/CrckqFnsVRi0LwGxFSnQGZq9TZYxSbL9SVXGRlfs6+2YLVLJ
bzw+6U/NufFIY+AuXkEHFbCZoDqUifZ8MS0MQqe0+RSPdw/JEdEIPzjHcoJPXbL8t7AuEm1smM4A
yrTf8kHn7svTdTkEGvzzPBPSd1RNQ25oHIUchviccEpFXpTkKWav8qpl8Vewil+9uaOgO0XZHg3N
EYwCo7B3LDRSA+mFmuyxu9dDbV/lUKnnn+QEAR225o5eeAkmIFs9B6sCNXvV+U10C2Wd3KIqXFuH
5pu3x5aQilfRIK9M72yfYmhf4OtA3nejnml6qP69u+2su1LbX7a6q+HCt+MVLaLDUYF4A3wD/IwA
FfXYbAXOWfT3FA9MGrZ6Yx8hz4d5fvsr6AD2FQrYzUeaSdqzlYaRivW3MDaN/EHZku+xIqoqkAj6
HvErnX5rV44dFn2Y/OcFRoPI0JkBAJ8IxYmBQfasL/ny2WLW3AZPOufTtqv97Yt8UUC92xfs+xFt
qkxdsHs5oiVbLWcvzxKuERMaFNEJYyB2JigISD3tyWYXrSe9Fe6XwNJdfveklufL3PQj+/aiqBgj
Jw6dqy1DsDHoFGq15/CUHUWz0JeWMZJ5OpHfZnQ9SBHkO/xr96criM4DUM6XmAoFrfmKGZim79t6
iKb9RS3RIH6cPm6whORN/EBGYFq0hiWqymZFquCn1yE4BLVTJgUoMZcID8z58lIbeQ2a9A8Rgblq
h8vyv7gV/C823jNxTvWvq2UTVnuNPLZ6h+u6x/rY08gsZbehEiqr7zPRo8vS+tfdVs1tPzYZubew
yF5ziYThWO8LBpE6DlSB2cT2kuccXrz3rL370PXwL85cLt5R7f9gQjheTpIY6B0JE/njV+60LP9x
gYOuQF/+B0edJJ+xMZkfq2B3mCij/WBpLcyfQvY0gnZknrebtKoR5ntbxB66TBRpfIf44Cpl9gF/
T5K3Die7/2C+M8qme3pAbPr7tQcZQO/nKjbQuBEkhSRrwLHz10akO3UDrKHz5RyoJmTFkminJRA/
2fy6jyYf/o68u6Th1L5AyxxnBhuOtgLN9jLHUWfJnpVuGOjMAh+URPSJKGqsmhwdciiMVXGSVL4f
3wa28djQCQtQBsTmT0cUYDyXi86TvO+P9v65yBqvf1R/GQB+vfNaeFnT7kAxdW3emG//fdW6Z1X8
W/gRwrlZW6ql+32wojzVTDd0IVKp3Uix/imp6ulvJL9TOOU8FJRv5wOBkgNr/iXod++ebWADBM2v
Tm9wtVIVLNCFrgV7V9sp+GkgC438rx95HYFSHBwoW2CNz/urhhitYnB2QkboEA3/vzSiVe6Rmg0+
XEDkVWqMBSKzY6JUuVRZf4N+0HmvHjH3W/bENqADb5e8hASYqg5BhLwkIvrkXN8RFf8M0w02OreN
nSMFOX0BKNSVEqXTvrN7xTR/kGBi/tpjLszehY0T6Lk2+gBuSJcSn5KX4IKN0f37jGyLxt2uPeuM
b3+gDOkoKdwSDZGdHIKzYdx/EMPwXSLGUjb7lz+ZovRJFhH4fPOdXHDX+zR4WfuJk1/uF2NdQvz7
+XH5YyKQGFfPdDMZwZ3+5ivlstbizHA17PDQIuFzJSHxtYu1R+TxcUipAg2PWZm4C0wL5kAKEiUr
nR9mpUlxO1Knd7De0wyFBX2YpzcX3WbYx050DbP82GhW8RXXc4GIekIP5pYXaF2/zGSVdHH6busL
F884IBOxDD1EYIRn3rcDyCR+8uKiamy7EUnChCM84OQ1l9GmHhWGi9+TV/HGPItwmGqSxHbJt4D5
EO7QICUsJ5KgpFkjVjMon2zqPe2AanSlmaUstr+0KljK5f+KWm3lhhfHsaZqtn3zfw7kIdmCGxvp
isgImttnv0ol/3UUlHFQSoag34TTG/8IUspN3nKufKvHLOasayMVsygKxUCO7uakdvB+rrNPejjV
y8OhHTeJ/N2iptNyzu7/V573mLwCj5LyTRYkTtbgaH8xSfW6PZmy7gU7HJ1WKpBXtpRmBJM2uhW0
Sr49r4dUYYOgmJ2wcd6nrlAQp6Us0aCBNsTTrX6YrkvIUTXKDW7WIjFQnqWZrEKYB/3C+6fpMHYh
MnA8HEKpKNHGEnt/j5zs0Cfv9OyZkqKxgwnfybqmsnvYS0xEejbS3NcnmG9MZTGrNYmnZSx+8T3D
VOkUnBJJlHcvj5z9XRoqepajlvQXAxfHbTqAQSrIdIQ2btMQJ6AXwDxDZeM29vMUV8jPHugKcNKx
enIzWooTL5EtIBllYEo28p7FJgHDdNrPboOIKEJF5IOysApDCYNCUDDKYn3PiqkN5RWjfqQeEzIb
Y04MUUYsL3B55RQ2bN9F7/hG8SgzL1YoLKf2A281+CcovcLdHsuKF1FT3A5IP8qlliME/oD/FBHB
YyYlETqIqY4ycTtj4c04dk0pp4cKmnc253UB/yFFNZZHZcB0k8X2FtU+rhU9/uRF7yV/BOz9e2ke
MkUSYsLF+7F3QgwyCs/bYNJNLY1gG1hq3UKQAKqSvtosudEDfeaD/8qHxYOOXWv7iRnRCvnGXPby
6VvQIyd+RxPc9RNQ/Zn2xRpVEad3JsFzZjrdXFSLwmeY1LLMOxFB6KLZnFu1P6GSrESA3DvG+RNG
6ew+GINlVdaHERkN0AnimFXgyiplmImGf60sFmCpUhVzEGxXynR6kOZ3JT1fdBOBSIy4KwPVQ4ZO
+zsOUC0h2WEFquJGNSlpT4toaiyaBfFGFQwMp42MUhIfdNIT6bGwIXU+GoLthpV+9/U3dM8SviTq
0m/ywvY0d5xDZlBJGGlo4een4X6GyFY+7fj7GZX2algJ63BPtLBlbttJxTlueOe9qrybhHpymLBy
vqwT/NriZYKbzcuNzmuREQU4em+843YhMnFWeu8HM/YP4GPHrRPbzC/VCp3UPP+iH9FPUOGOf4Zx
uKoH5xphxOu6WxrQE76ThjIUu4zkdGHoO/4XFGVy5Au1AxXonEZFVMm2QAcL0T5g6GLCBwadg94W
XsiG2faEJR41ZFgtdJqvypZjEerh+ILvAuhnCv6P5hbY5FqKU+ebnTLxH8Hqjz7BiekAQpXkbVqb
g0m6S/XhyISp5639bkELs/fTiDtlxq0tzmc46z6KXJNOC2U5Ou/QvKrVvnu+peASZh2e7DkjmYrt
hWu70yy6niZlDAoNVfvwVlkeqU0M+T8lbmv4Ir3xaKaKq0yuPwq6tVAepCZl/qUY6CZDscACbfBT
BIDRsV76k7tOSldjaGr8DvqPBEmWjEYtERSDJL+SfKNWiSNx3cTP9hjKWhACsCEagolxJETyhwNo
fmVB3yWLIcgkItXKo16y6/+E015C2hFj18LoCMH993oZIXA5bVLPX9OE7hGNc4Ueoa2R1nk1C7+1
ujPC0+49lx/QrvahS0xq25YUdM8zbAqcngLZ2jJdyjbHXs7DrFv5MhEbwgjOEBTmodMET8iXk6Ki
T7rbADz/2Q5zbPRgq3FYb43k770z2q9CIVP86ZgioAbeuC+pyTyQ3M8WV5N3ZBbhd+zRxEjLAje8
JSxVzHeQjZexXHR6DcpsueFwEc1ZS7GyDc1hMkhYjd4fWrRTbK9dF4nHZiv2BW1S5mLBPHopWddL
fzU20OLpw+VxUWmtztAB9Ic7YGUkCbNckzYR0X/jyiFbp1y7ktD1OoQqvjuAHeInS2YWLWMo0cCm
fCMvfJyR0M2oCd/BWU8mKufhc5S+H9p24nXCMlxC4hkztxkDwXWw+/7svMI8FTjESsecyhPeL4FG
GiNWIaH/WvFs628FPeozKKWlRdFzMrb5hJgAouZ3wMZiSrBpDa0etyg93ANenzAUf1RQFVfjPi0v
cajcKE8HOVoc2DqMEey7H+PrxT0jV8Q+1qYYX62wFoBczmc2J4TZwCXKNmLhEvS2xgRjY3IXYtm6
P+gIQyNjzgjEH+Wq7eZNFdsZ/Fle/FUMbV91eXDdsD46VivXW+hXAVQCOLdwIFkgtp3KmxnhHRM4
RPEegudUX1X29bBxw/b1IMT6lohEEL3QNSHltIIJvMjzObyb6whX1QysSGChtC+ia7rzbRYyQZt4
RZ+aL49rZDL1ZKaHtQYG/nRFtaGC4hwmMl8LmA02lkHTysljEHgR0eO1Ayt+blLBCqRy6CoVkV6s
o/xNfdTquxHUihUds1R6um9XKxsurNhXbsZwvqdadIwIDtk3itUg/kjP04aX1OBRMk+W7LYnkOg0
pWJV9KduK5ngR+GmjieO+9s53TfUHfgY1RppQX7UVwAijW37U3569E3xErWuwHPaS6kRam4ErgCi
6acbVQI6TyTLfF9Elz5gM3MfaM9+4pECeikze1YXda5SASGzuDrlKf+x/lP1satNIYvD8MyJXkkO
AdFjUthG89XafnjkjSzWdj2fNRIHtVucnld4BLdaojzTnStcgJYA2wqAji7ZJ/Yd4GJ6PwSeUxG/
kkNzuDWahJf2E3bu+qC9DD1rZ/115mYfgtKbcw9NrdPcNhMHWg3+GBRI08EwfZ5DbKNfVA4H2y/4
ikCvC68lrjpn30u4Qgr+GE+Rp+xQCTvU/H+zNGI+niP2AjwTEW810pCtw1dOMiP5PbVT4Qn3coCP
otC5JwUgSgFOjjylsT/2ZT5+JPsC3wI4G/8EBpWzYBGHRMibtufDQIEHrBpDs0652oxmII0nZ/mC
2yuc2j/Ogl6CgI7SzMVz10vOdoG6OfVNrNXBDfc4/AGIDeP/ER2Mmy+tPZyY3W47vbKinrnqV8+J
/MfiGCvzeHGL3gtQq2zfW3uN3nPOu2W9Zdk/ZLwI2K1P7sg0rprEWVCJMBoJLxL1hfZBl0mjxN8D
booLaFncn9tfdlC6VPFA3BbHHFV+OuMnx6K1d4qslTuZsvtQ4sDJjrMlSH2JAsWL37eRdTGfkxbO
jOMaAIhc8iCg5wD3D5wQ2uQ5+ue4f9zyc7bZ1o9qEjfWVWF3MdP6oNBSYwxev88B7qW3Qnptbjzl
NCxKUXsyxrWMPERIki/C7XL+Z99Pqig4g5yUdzlVZxcTfAtbyg/NlOoaljMyNQE7zpC83MyPdL/Q
d5RPEVZvEF07f/c5NXqFfBOy3RUxdJP4y8w+yo0+B6Y+yaVLtg1V3TGJVJF2ujWLuy428a4xTdOC
F2JwFG0cBysxxnm7yu2uuk4CnDlmv7LNcf3DCTMIC95GrLbPX1hYPvhMSIUp4E3Z8ZfdBgbGPvKw
PG4nD7oeo1lqMQREDa/k8ZP8C3tU/BQF3+CyOkh09WnrNAZhdnjH4j9egY2Q6QihpZT069vEf1m2
vQaK8RAg6zRvqmYI9yrcPPit2LYQTzou9Fq+4iAjuxSaSwrZM6u1PIbfDtC9ItExb8HvhNkVf++q
tk/j6DK6rkvfdVvf5N1dZ4jnjH8Lytw+O+TYKsHUmjO5DjVNiHCeuGadHTbdcK5OoTZIkwZJI5Gs
2R0dW2r+NsgpdJ4pyyMM9LD6Zj6Y4csNYOd5NORdpl0XNSlAFVpVOBE968/fofgSenmciWmGKLT9
WeWPoWA/lkwxEXdqGuSrAoWCvhIkyeDZpJhAho0tXUEeOmhYpcjGaKuPBCjR3tsC08RmL30Kb8Wm
XNWFx0fatueT/ZUQ8YqQ6Ugl3GAkSmham8wIB1zMjY6ekDSWJb5+uuP5J+cuETIaVLrZLMK6Utzg
5VB7oACvHdeNQ6DqA7lhvGENfxq9YPGfBSUn4aAL1gPhfLALfghG6v2ZIbB9Q8AVMBclmNPpI7Gw
ZkyLpE50RuOkI/hQ+o2JtTQHPBmDn0g4y1SQxwlABDRFJCoU4eV8dpVEz4Uan2GoOBdV0LaOR0pU
gWJadurM1nB5ZVEJXg/GhnDAd4aP26X5ZVknLaPOxtUpDEZiQ3iLyXxw+V6pbt7wxu4+0ilHNbpJ
1csISCe34MO4m8UU2+fsvZHS6f3wWuXhHGi+G8JJ7yXiKDyyVoffuFxmZLOTZnbnl+53SmuBeaIJ
jrnEo9tvcSiOKSDYT4+KLimepYV3thyjdlnoJLgS7m24UucppmyI+R5L4/gwymbUjM9qKhMz9kUh
y3KIApy8jrLUGKDhL+Pe5nbqECrVjA3r44rKa9Q9PJf4Tg/VsumfSqZhPNqT2wZdAmBXJl24GRgH
TY1dbMb3/Xo5n82pnqLeCR2TW0Le/qFIfldYWkDmM0FEb2iCyk4Y9PejJcwXp292nVGMqml9FBdg
F+YNqUfsuZ21TmtD/gFgp284oM4XJBO8l43yBk1AuOWSxGfIXXVL0KxnkgZf1EALAFQJL2dOOMET
KKQ2uCLAzC+ElH3bi/8u1+JYnc1C92Vd+C2gE0bqJyC00g/rxBrEbwp4K/r9l3UGdHQdcQwSKeSu
WZ1PB2T0mttjal/7GyVrxe9jgERyn0lLdJtbbyOYQ+mkyCzYy7xVgbox3Sq66MESZZp0IkjEO9+p
tbZhm2b3SLKs6N2UsNQjKIrNCWB8WphEpmUwDw445g1fBhVmsdCt/llFOqSC5ukLl657E9iNha+R
ou4zEVBUFV/9pMwSZpYnN77wYOkn8VgrVZDbh1KJYZXikuPOfj0Ef4XEag3MDylCSuXD0UG2eADF
wu3YJp3jflgMIdd+W5nuruADT4akKjUpu2gkaJH6Hh1kJ9IpzllJne/v0AIStVw5G+xjrAtAP8ng
/R/Qe1oavn/wThypWtwSrXFprnC96LI4GMfmPpB0g57UmDu8M5I+AsynL9P75sPQLyfGRF55EF4u
qQ222WIE+Twd3/tZDzK1/Xed7lSSjX/KQjazORkS3Lzi7fcACN3+QZdaBJk6Vl3JyUJhxLbapAyf
co9fy4gXSYobdKkZ6X+OMi2JkDbeyHYN77PQ7RDFLbN1OpNGb+P4uGp6bdzu4bnTjMz55Iq+85AV
bsB5USei66+mYucxhpl5+iyPYH7gHhKXQUkgxXAs6ctJSaSqaKI+kRfOrfFGu9/+jJL3k4twCaRM
BeRrjmGJeObo+IQitV1nGrGUnya0bG+jU2NrWluvs2bKoSyhNBmyC+ILzvHBbI4IrFnjamqxqlxL
7tHXt3EpMuGNBvBHFhw83AcXatf2UIGsoDaSX2qhHt3TnXceKTbP+EbsgqvfwpHDtaqpNQFfZBi1
Ex3pz7SVZm3UKGklIyumruL3f17sOEaVNLK0VWBlFKQfDrWV5fAEqznr3vLXxBGcjVxk9LcsriWc
EGSp9aIP28Zc84uG1Oxxwib5TmnrR5yLFYK8UMhNVFjn56m2FXlJzxM93eVV/J/CBJJ7SClbiF1Z
+7JwKfPneKK5OPDyULdPl1OjrBArEnJQWKdL1rM+EWfnykLSjRvgN+MeUB7K1ouZHE5hwj1jJ6rK
YFHoSSZetQ4I47kMLGJHMZYtF4j40q02jV0fhZnKiT5enmvVRXa1MPf1t5GBHzN9Tfm8IpMhVbP0
MCf23rlw7Tb2/eWyOGgjze5xvRzI7xi6VDx4KpgP6v9WYF8RliT5+KM6yOCyektfgSydfRcfBhxI
f1lJtLPmEK1Z+R1sZj7jHLNs0B541VBRxQ2HOzhbr4cqEPpCriUB3ZvBybLHpwVRuf7Kn8m88HSR
NpAetrC/LhPMa0VqwYk1v1itwFwG88Q5cX0O7Mv5GidBzRIcnAzuEdu4eVyo+lBZLKrjoa5zGftq
d5hkUVYsvNP6/LqAOXWkkGOJ/P4AdNqCIT6qVtK2FZn5rEdp3o28F62DvgSHEqp50UA+80TF7JTD
aX5fcfJcaZQs2Tdg5y/XOpEhKcmhEM/ftjp684AyWkqDPDR8e87KfWXKVLBdN7RwgiGRSyOE4TNQ
zsQhYRplTCac0EdEW2oc1nF3Ll6+J0yVR+dWZI8bYQyFkv2HQHOuPKVrHOr/m8k1SoZ8R+1zEuon
g+1dwx90522+S5YbFoghcT7uIXZAtgYCiK9xxGRZGKyenaJLRUOgF15uWEI75QfJmxL+u4ObewTQ
yc/qg3LBAHY+MM7kvxE/sA/tgdV8CaKkTmFqJtQ9pHRh+uvTFfSEjGVPt9lucTLXo5WqLtBghU/b
AaTCnwL0X3YKnT58t5v1angWaugolPNRqOHHhqJnL5OY+SdntreDpE0DmuJAmUdsOWXgjSxN2zWu
28dRdO8Fcvf4UgsZe+ipk9D9eRi6u2WKPY51YTIm5saqE/zr6tsjZX9dh8zi61uUase6ll7EKtes
CIR51GTjarzCjkYS8xOdjPNoa9aymiCUKFWnVngQGcfRUmfs/G8Q43vlSArMe0gDrei04LWhNKvX
EodgfHLvKHTlpxC9zqWr7brzKyrfupOwUeT2xDMPsZyMUiZZNtg2LwXquAxttanunQTxIgVnZv2z
UGxBTNP4MRJI6bbNKk6cPCmhwpUgjws5JFYvqR4Hmbrky5wvO+Nd4Hp2LbTNYUodZsssmnq8SFNx
eWed2xjjSB4Q+q3Ue2YPzFrFnk+UAdaMs2lF52tszlNbRHEOAcM2DG0CfDQDN3L9bXJh3xYGRlk+
75fGPDDwewpsQ240CTyfzGpyS4bubbzyuUXcyNIzReoL+i/8Z5OrRJ53fBd30dgR2j7590RxEVso
cxSHfUCufD84E4FlY/or/CZSGKNnNXXHspeYH86X5q0DafnzemVoOjBNtKyTrxoug5JYJxoKoPKI
xc1AzZzIcwL/OfzJX62r8faBX84c6IP6Li/9plpXWtEwRaVhtJuREqHs2CuE4sSz1d4NZPcsnp0x
MfVxvD6TQkMudfzf/VSYmjC7b4Fhkaclsr2wIGo4ip/Ku1iWudyVcsziLGzRxAK8pIRAQC9GlJ/+
5/JD/6/KgsVxFnhx3ZPO7xcUtx9PY6X2A6mHu/i78vqaNBwd+0wYCynjqy9zDbd8SsFV2ePu+NPz
AHmpc1IbHOKigpOqeYDePUUDAKqiqNtyisivfwtQ5YCV4kEIWTviBNXb5LqF4HnRf+a8UaPpuz6U
26zpVLIW0L6bH0FvVMmQDzxnp+LIwyCDqukTpawyBDtepARiC2UG6R/sWHKdcJHgHIunhJceMU2Y
QDsVQOV/HCWzhS2OzqioDlC99vyajqbjNThvyJYWBCgURamIAmPj9yWUwW5Bs2NcGdk+e8FfztFz
JzfZVIA3slIxDxQTtmAVqmvK0ulPAHjRtBw+R8C/Sh9szMvI8g08D/UVIpnKx+JUar+FY8iuRE7J
7LoUEbuugFpi4vYDnFS2Do2iVepjTdxBuOVICjz2MLgCSUe046RyWRoDWgmcbXac+ZCnBHXMEDBj
F9OorZ9asKeLTQokkc3skcaDeg/FHkL7KCWpK9Crp41cqtmIOUiXX4qwXAeZ5q+NFLt+YY6Uzfdx
R3mdHX0836WW80NBzcEK01hKS9bpJRYEj4ovqVQ9apnGy3XtRSXsyuQMrIwORTIXi2xmLhKxlW6u
M3N5jt9aFQilFDrHzV+kdidR5Roy0Pw5qcPajIeUcPrUBHqFU8owFvaglt3PqN9XrfvB04lWCUQO
SDOIcZAj3Idxzj1kYOkKvx/m26rPIaiBPj+xycDYAuWAHPeSgjM0g9ijohezarZPKTUFpxT7Dys4
jRxk8qFkhKYYcyfROpbcVIhi2L9W4p+DOqNO+hHgQojNjMvQ3TGim6+NwAALBHER3YraqWvKgb2i
lXlTcrj2zBRtIv9yjrVb4oosx9EAxMzkeYfl7wSO8WE/EfCJtqX3T5G/67kShSFTmFLmfo7JZQLC
DFag0Ar0WRvWJDJhaPyeQxD4uV/y8YLuZayHZK/LcCFyXk3vrTZcr0GCURmy4SLyTlw2t+0oiIFu
VoRC6sHDoUY1kgew0EPbkd6WgrbPbT7ldY+o6XaZrHJjrkyVuCgD9ZHxZQZacDpmfJkJEgl0RVT0
2dr0o59LKmDk0e3zQ+uwDpN1HCLn6O87gwvP5Q10TnDIapeJzuJLOOyXuOVqfuwUyudEdvsdEsuP
GnXhavLVpoONA7/Pd8TSxkZhbKWLec6ClB6HIiIhI702J/KPFXfuPv1AH0wls+5OiwNFJCSuc988
lvGJ7O6qJ2J/ZKWLmE0tqld83DdiM8dNync0+hVI5JhlJuYpoSem5ZHzwN9yhVlBwPE6VJtGaETI
js8Qtl/73mIKOO5hwDuYExm7jT5ESMLeI9piAdG7BdhHFGoHRQ29+13b7tPXe4Hx2GUXcvLoF89h
v3Mm3hy/zUB0Nq5wbG0ZILHWSLaC67W+vMiHWuP+mm9aXSdG+z8F/S+YyuJhDKcFmlMzAsRvm3Nj
M0YjjfxPC/n/EtGvpPfVsToH6n4qYGGE3+D/JsW/FN7aB68tt6dX0GKTyUqX07cmJA4C9RJfHYKw
Au7TLC21uui7hWjWICOqPLraTmA8rlJau88Qg+qq76R1kHlgvsUjT+Zjyo3iphfe62E0bQIuvku0
l1CcbUd0VGivJJ6ULeOM+FDMYSxAYY44dkk6C+rN/PShnNNtk7gAfLSlPi44FfR8q0uSlI/G/Bn1
cCihYS3vKXdn9O3Gh9VsHPE/1R8Oc/i7+ddT/0G5RxM1+aowgQnXTSVNN18AZJ67cV9p2DrH9Ag6
zEeXBc3biHNQFhQT8XIvDtc8+ygoHQMxxrpevnoyDHkgGid80hC8RbPmwwPjWccSVuD3WV0/gtPA
lmKzNfh+M/gKW8rdbueCPp8eycg/d3JR+m4KSngMyfMXzlPELzMADqMhCpKry7qPid2ncS8LA9Lc
IP4L4T3ssB47vPXQByuWXE6FXfLxefTyHJfDqpBT7MzKhcwyw/r3hLOo0fMGCNylh5L22rLPHnE1
KydPwMe1JtfozUNBNxOB0bzPnpER0MwL/j82KmSTJAqQCTBzE5b8HBDL0eEC/onH9P6Cxo/8dYJu
dm9H3PHmDitztShLdN7ymMUNRD/eEQSTXF1MEwnRRNONPDR4irOwbIuhxGNFqEmOQa8Jsdhd+RxZ
wSjMOLUTyzdkwUYGGViu5B/JEsVr6HqA/g2QrJHxOiAnQ2lG5tu/4qL9h2tTmx8xkX4Jc2WPJQ4D
BRgCAH/+9ED/spXXmdYS+xwz7N9Uc4Nu9Pl6PUxi9dpPLEIWxmOJUvgPTCfv2IsBUkjDOzRcBdmY
1RA3qKjAY2WhK3PZzOFy0FYyQcAyOkfvoreD13gWIG2kVtrmf7FWLJo9lOB3s0ukA8rv2dObPQqJ
jCsHro3ijUTRWM7xp9vmSznexwnjjmub8rDA3o7WLo+PDVk6tygH0wgWr3dQjhBygPa68mA3nTG3
zfmH1hVo/oMEYYLAIBdgVKlNE6XNL7SW6iUfoVMDGOvZGQ6okL1uRVv2mgLy4NpXxFb1HfSpY0Kv
LK+orZxDHsJd/cDtmq4wuJKjCng5K1hTszKZWBslH/gYBXP1/svUjKU8oMDNha9mQYY2vKomubBx
+SFWYvTncNIAavCe6oggxD21VtGbjHb69/PO8Qke6D0O741gkLMmF7zijTlqNXNiGcUBTLa+NxPr
a2kWA5+OBQnttsvnYA0ok/ErGo32n3XtVoi2XcnN5g0Nc3Q6tapxqiYplwq7QeHjbBwex0IbZ7aW
amwau511sAJORpwboSDnbDrKbrQwc3zoVAW6BrhLAa+6FUGBy6lBYQS8l+JDBB2pgt20o/4yKhpA
nbRzMo0HMOTADPf6BkPXSfpI11e7baly6E8XPC50lqulSrXz19TsxarPPMkpbU/aCvivS6zbeCQS
12GqdivRFSBNRSwaYBwj+/A+r+ADdkRcXS5ocYZTdxqj6w/Q/+9dIcpaYqoAp3NlkIPZZ5rrokX9
Vt9qvqBQTwn56TBCwH0YROlTaDMP//DY52G16ruqghv6YwgXrKwIJx3vGuK3NwW7YY1LmhdFR2U7
sfO1mqFOYwe8ym4NcZLz7JGzLxF2w1mgglLml36NOnMQP8vIcguPh1q9TrEZeETFLtL7ofUBuijz
I+VzsqSjsm/jtENgXjwfeB6h0ZruuYhgAd0sK1YKbI6FeRW6F33x4zgQtZZy/EQrNo5pHVfIjkhV
Utk8YtXhjoHRXe1++Ll3cQCBpt6KEXSMesGAGEsoZp+Ofk5lhugneDozCmiWKAWLCc38b3FQ8orG
juKMm9MXYi6uqIS4N51aEG2wwasgWnnVD4wDrn1qFRHCyPnhREbyJ4ItMJBSgLaV8LF6Hg/iYjLd
OqxzeNXWvTWj1wc4M0U9s/hcKoOHxq2LT/7rdo5EvD5349wEqGa0pnhryZD4oTPrG3JxK6VMe6c8
HjJAAUwB2wd/EwVzNhu/lkW0KuGPAWBhO29ujTR9pTHlikW3TI2+fqhkXVo+ixgzp4iMwzYanbbg
kLQ8vOxoSwMOkT7cfEdocRfgeXZhRJnfYOpG44Cb3U1tC9PKnXRUMDSa3H9AUZYo0fmNnGlwooDd
ppAhMa8jsf+vU3gZU14WGqqd8Ctos+iRhDFt0PJJ5m9CiqsplHhH4A9636tb/sBWc0e+gUXjx6I4
cwB6D2benAL8kysqVHp449DA8A/dwRbtl4Jy3vilbWcb35ABLnh6Wrg0f02csPpBDKn8rxvy3zoX
5+A60SzgZeUc6W6iaU41pYyFLOECUXjhS4bZ7RaNyMOLg/2ARpeLEBvBfVI05osI5L1VTnrrcfSl
k2gq+UCdGL4NrqvADc7GJf4EgtlMZs1nFEwUByQXi1cgR0LzWf5STe5jLeVtBW/J7vC+Y3Ig2+o5
EcL5AhJourERq3YZ0rSWZzKsQVpVb1feVABBeHAzsQSrHFkq2UC91uZVJcYkozYaZBs/iwwgGOpP
wVLCFrYurhN/y5knievli2cdjfCiXGpGYF5JDsOC6P+XLvULGY9CfhOY/do+IOXXjb2W4Y+oc4Y1
E2nZXqNvrETihfa5hBVpF5dEBir9aSgmUhQBtVTejN0FtkiOzIXNp5wVrNidzZUyPHvZZGTswgKg
wJK0LGY5F/HaEUBXyP/f6rd2yyOqgfFcPdJ3FM4F+TURKngu409s62dfG8pWxzjrNbsFLwFyVLf3
H3Pkh5cLQC/Z1t+IsEG7VpKDHgxV+q3PkvG0x3nZOXP55K3nYIvIynP7sOMc81Yl/Fx1qlPEy5Al
55uFfEkQx+uO9gkUqEODaJYe3Sg6jbLdo3+70tPOXhyQe7DByFy4617Zk0Yf0AyGSObew+QLNtrC
woQjc6P8W9+bQC8INn8jy9Oxuv6HEfaauqSg3VCBAnQp5so25iIEtt483FQgkq/Pi9B8GpdLvVgo
FkGuJU9IuzmEFSB9hPU8t9LKgqs3XeL5GuvRCNNVK9ZvznohZxSSTcjdmHj8A185VzPCQCaYCW6c
eeBIowe62I9VbO2hJoYv4vCwXd9JspwEX9djwmWM+ebVk1VMdkmuIvpA/EFA8xzN1FCnOpSHMT0i
vPDxr9kap3ZEJXYNifWr9JGB9DyVzAVe/eWS1Ce3PtMU2AFJl580CbcQu9R9XpVxr+p5X0CYuydJ
uV/QA/zFAY0RY3DeR8Q5nYp4rxtc7z5VgP+G1WkVulU4bjFXCyLQgPReJJyS+v28oXMlrVMrf47X
vdEjFcBAAvButnKXxJsBBx+XrMRPE/EU/ssF5HjXc1W7E//uYLCDagMOHhD0/qaTcIFrcWtAz4rh
DmR171hDC6Kpuw/yW8ZRkumvjk2urhMyE7FWWUha4RU2SQMENKM8yBJJx2IemT0aPTr1pg/p7TNR
W99Qs2spNkURh3m2IbgNiMPKBwe/160xiYQED9JcmaXWrpbp6og1B8LbaHqU3d7t3o1nryJ35KOx
ZqhqVSulTXdVSjYgeuZQf7c3Pu5voiPJhczH8cx2FBu2WcYdSingZVPCVhslZp9Q3bCtI6F/yPd5
dKteaQ7zqdMKf4mNkKm4FTEZ45iqMiO7CaZbs+9DO1Isu3zcIwgiTIxDF2GOhvdFpw0yU2a3FpjQ
oTMDZtaaZ3tnpsZnfXRycDdRbFZKXlVf/ZGVcqJoSwAtr6tYPjsOH5mwd92GlxTgpeh04m/Vyb6P
Zu8izPEDwMmo2fJj67IwCAHnojk2Kugs7/m94eC/dCGxU0TxQoGglkmu5cDH3EpwqjS4qA69EfG8
LxTlbyt2RJGd/kKZ9vcihBehuHsh7Zcel8aKJJGTfPbmPTReqQH6qoxQsqRM6HDT3bAK9gIaZiIL
6G8F5AVy/BsmGqgZE53YaDFOAFdUuSDRvexl89kWBdXS8jKV81kwqaz6edvWxxfKuNpYvNl2lH2g
EU3TULcHgF9AGrh+nzpbPRtO6vepXdj00jK6jwWcGg3+ZZ6c0MTefxU5/FICrFNerOK4eIaRdAio
gjBJRyE/e2RCiSNDjOioOQwDtHKQjI3X4NxwaY7vJsfMkc2diK7P6X495t5lt5knSO08VZNg7HJk
/zEjX7165tnABMkboD/fmSfrON9Y7wHa5yLpMcsr5C7+m4NbJe9Ue2eSEkR5EJzXab//2fplWoTG
//NW1pKvcRvUC+af92pwjAi91IdiR1QmXPB0eU3DhlukodPGVQ4SX1mukdWhuXa3zTNIbvSHz1OR
U/zb0t/QkmggMlw1s3ds6h5l2s6Mdl9pJPPUz8c3bQHQf2ZYW4nvU/W6CHYvAD/TgoYEXBUfnRHf
WgMWK1Z6htboib4cOhP0IzCyLQ0XyBJ4NtipblmGo2Uir/3Eu/dM4hxIguS/TC+hsR8G+RA7s5+o
EO9QAENwOm2uO0oyGiYve1cRx02a+raNB8+6pCrL1eDD7RSk2/2g+o2+qXirr3ntMfPd0Xq3NkmV
M42skg0HEtb3Q5OKwEF/RJNYLuywYBeLhRCciKcem92Zvt+8yvgw6vQDHfu+FpOMBlxTpcwrxrsJ
KI6IBwQO8O9i0XKI3LgGhtNCo6JR28oHCGxtcsdT5I5TQbSNvxWf3kq81mCo/xHwjjRT8+udMJxQ
2dIyYWvwUlYbVqAH6aLbVyyNfUSQI8LkPnSZV7RJbSLVBBsu0fuoOkAengf5+CttOONi8X/jt9PR
1RYtSv7OsvceiTxZ1DLX44llvHqEQ7Utcc9jSmJtb4PxXWsZ5+X95NI2rPnV30kN2uWs4iYHthPH
LgSQdEaQpITcivpVC+EDWmMqLOnYHd++8H1LMd1ZItbEaQGz73A2TQ1Xofw3QZI3UW3a4sEPTIUu
2WpQuPqMIKtj3CTdsAZggZAKJX0fSC61XFIfrgmQKP8kQiZtdgEMA+wkAmfza1ri58IQzU7B6LWb
hGqRWmMOxRW3kL1HP4Tn6FPAOy4xBPCHc4ggyw7Zd2Da49ccyRWwfhOOHxkqDZWl7Ek9kGGWRVvS
EHUKtTdb3UxGgk6kRYfOJfTnEz0jbIvUlqukc/tWCiR3rvLbZvLin3f+Nf43fT4Nwk2dOKZlSSkg
YVRhJNq1ynl1d9XyjCRZg3lm7Kfp7XtqpZ605tDgKFLLHejAbkgGnirAECLGMp8q84WHh70XglyH
zpbzUj2RM8Z21sUtxW10AocTeMP1IhOzk4sfA1Z8/RTTQrpFN7aLwBW7eQFeO0pNM16V7+O7bWpr
knfke3L6nIkLcLDHGtdziRmvChVPbhjM2AS888aM7Os7lSBFTgHbcpISPMjM7YcZmZRGIOazgPIb
RlEXt6ufmpiGxEylyw2AuQ1iDbAsGarwu2dk1gsMoyVZKw7mV+m1ijDXLZh156XT5/k0yMlhuL0D
GZoS65Le41EXeJrDfk6mPzN06FFwQmNbvKf/kppRxkn7vVADk/UcaabdJMac5xQMkFgCEJgICule
VykGGvrp5P+WdrcSLZ4iU+Z7AxJwYRt6pDXUquE2WmyOv+1MsDULAYRA1mQDdrFoIGkI7jM5hJc1
Dzf0c4EnJgTGUYA0p1TsqA8bhYap2XZ1pgdXRVYIQuVUCgboEAIJVsaigr9GXuH9dwzSIttrG3my
WCWm0h+Dv0eyhAeI0hWBR42ruA6CbmOguatyO3LStAu1L3fQxg0MUjXUFyNFI/jF75vSgHchrgna
zJ/WSbNZ0/dE4QpOmQ6AzQnpRUfxOBedRWdhdhWs7JK8461xgcXuulcYS+MFyrbeyeYPyUTDIe0q
WBYbFfEBePzHA8pgI5RFl44JQMOQ61/WErtiPR+bhHtjyVeFdOsYV8DQtpIq1PTRY3QJ/DvRJnoD
7lE/veEXOByOpUiXmLtNHfWwp7ZiYQ1F/HNJeYAqADedkFw9nuaCyi5bIphuwbT7fcMInvUvCGCO
YfbfBqe6LlHdLIwZV5nM1E6ESUpKMHTX9WMN5/kI7pHbOkUkWLy1q4xe4tdNwD2KXyZVas4elKCu
7MuPQTjBGoWp0PGtxo2Avcm3+18M/02oUMr3M70HxGStSSB66Nm4pIhS31q3ZKkMClH+Ss4/32x8
CUbRSPmREp8+JAfUhZbcoGaqxMVXjvc7fs4uZkZn7M0cOy/QYD/dXgMyU4qkYU2/iYpM/8EYXkjl
l/GnoEx3AZTXyYy0DQ2CHflLMCYz8lRhHqXO3v/gyVF8BnByHbjMUGTIYPZNW0WWVj9PQa7U/sVA
7/FqQ46wPZLZy77umsNf2mwy0fL0N11obcDLkPD7ERVpMFedrj/ldmv6bg1aVaNVQ4zMNU+4GtPj
aHXO3112jDZrc2+KSY1mlN6pr9W4iMcAixbCGCYKg1vUVnecBWm1UXvdrAQXMhMG6fouhkD2H9GD
DZL2O+DdshalEqMSx05SvZYdKk+EaAMml3hcTfWRoD5Ccd7pYEwkRCENsZ6yYKIruNBrpeltrefy
gmbHKBQ3HntUuZiaULPPThG0easod3G5b5uOKwiACKWASJM6LCxFr1GuYQ+0cyDZZ+wpSUSt5Xwm
PlJyKNrswtqzwxZF0rTaRisxnKtoJSgVuJu33b+uhj8YrNDu58l9VMao1S3EFg/Rnll1Wb5uBVfT
PxB6xKTN7L09HWyCOP9nc5C8bcrFuRoo7vQCKchYqrKK3CC23XQzQTFrxcjJun72idYl0pD2kk/d
FQJGXfUw8f6pkZALOrWfexTSB6pLNI/iEwxQLsNvBzjVeuaCigWO1naULFPuV0sMbXG9GHMWd+Mv
cH3LrFpw05CSIX/xSCznn0vlmbasc47fxSFqNoj6Jh1x/8895kamkO7ptfspNTDXX5GXtEXMxdIP
m+YlIJmwR9GZB10QA/iM02KrCzlUjRrVRbGqbuJHBIlJ0pucpEu1x8RnkSa5QMmuwB4w7PfJ1nxD
NicM3OR7xPknjXbToJshMvYYITP+JCqe6vuiuhtb+x0Uk7Qs4Ir5e4qGxGMoWiK+AUy5Ta9+9ElX
BWRLcJb49h6VZRRo/2XIZfEhCPHpHJNdR//Hsq6ugfC9prQ23/7DA3QhTJ1oZLfXRwox7LH/WDft
VPA1cdcmm7GOLjtMpirrAO2cJZZ48EZkPITes9jy010sh6wxlB7JQsLtbBqlgICGFcTBKqardsYm
wFVa7ZH8Xu1E1SjOGfd+3C5TX9uKMU03EoTgfMDGtkB8WrM5L7kdAt/suphgsL1UIWR4U+tJVDvu
36Vt1lgjF9ax1hKfysnZdK5isSL2rH41V+01iJQ35SxP9NJnqhzVTucpZ6oRT/a3L5Y7D4zZriMu
d/EKz3wB5D/87KJYdKn1137m8ah9sKvwuSQSub8eGB0kPeYpZRlmAC4BqLpBXu9VZFzkGJvRz9F2
U9vcghntYFSFdQtai8FPfe9DnVG2TrZS3KGGXowLpv7wujvHztGhr+ZiWR8uvPQNEWkzQKKbZywo
LY6bzVdfk5KgfIvXJpxv4JoCNAyOrxImgFbooqF39N2dMUehvyR6gmy80VWi7o+19/dd0HK1nVQf
J40zx1TJ5fNm0douFiWN5krD9ab4A4I7hUQN5kzRCXiPfR+WbRVa+FO2bpb2l/pQTlZWjylpIufT
Z49iQFXFuSrnjtbfUQtM5d6BlbhT7oKZvGLOj5jXBNS4kLCk9aK3EdqPZ/VQ+ZsvgKebwOUwJVxR
jeno7VF43qLp7aU2xdGEgQUGSubKWW9WSdrR0BsEkCwwj7G43YJtIXP9yOrfA3bEUS01U6qa1CR+
eewF9LyFsHN/BmKlEbDGLUIiql+CEy3QNpzhZJuLgdeluAuOqTz3V7rDXIbZ2qD9Su+PoYi50bav
ZMMm32woTeMPKSzrGK4eqUBVP+ZCpSeJUegLpIyGLdCs+kCGXJjqgxgRsCMGU8m15bBOisgOi4mR
s70NE7Ft+WDZymzsp52hSXZRHXvLFvvvgdIDtonehX9pmCDbIKSsSN1hkQAONYfOmZMMfunFPGgt
qkVYhHoE9ren+ltp8P74PRCQJmfZD/5xTpBAM8XfRxRTKXE5oJrJjHVJLnSkr8UYJWIFqrqQ19F4
fBkVSxAn+IPVOoino+nyPA9+lXoWWu/BN74XFZ8Zw8+qX3k5gZnQ4age4cJbUHzMbYmYA25UcYx5
78Tj9L5pwqinN5zO8Zzq3K5bDwoDicK2adj3kfEzJOAfLlWGGLPFfeovIvslUlVJpokIHQsZVGX5
wlRL4iaJ5ngU71PqAyas2fIWAE2y42jmEKQVp0CHt1PvwZGaD9iSp511xP8Ij0I8lf2bLSogPC6n
Qt28IU/61tCdDgsDMaNAuXOK62s4qb2LmxKb6l/y5ehU3q+/EkyjmYoKwkwlwhKROjAYgTdT+omL
lyiF0Dyps9MzKehTLM+XeiuZBgsRPFYVnukZEGd1pkVbcaO4VhW0U0mleqlyT6l84Du4dHLud0mQ
BD6ijiFWTMEV6GSTfE6NRV3T6vjAqtcU1aL6ksbwX/sToxLB3uACQ92xJ+jzJksi/LAwbldrvi58
O+9r9tgaSBJQZgzlV/IauC7T7XlHEpULSceLQRgSIjASHsfdnuHugPemQaTvlzbZmXSiApI5PkBp
WBFG1sGkVk6oBfMbf6UPHFkW230gq7gcCACGOCWg06/cqyky/X+HECezp/+rWKpkayhMjuh7ncE0
XS9FsDjtUveGWGrjNNf5OEQ2j8hdcs6pgf82jU8d1TzYE5tnjeFOjI79/beD+y2x88OeiYhrT9yz
KDCbDOF+M9haLLl8neFjj7/i5HUQ9L5+aOE7r1NXfIs6Cfwdjnf3n3eVGSDGcFZX715DxKonfvsY
/Wdp83lWW1/9cOhH53i/U4rHFLjxhZ1V9vERflpOvzDpiPITzGpPqAB5+aHXsaUZ/MTzcOYD5q7y
FJr3DhAW1peEdbS67fxPJz1R9LYPfw16wDvYM4Y9o/U4E7o8rzTunTe1h+QXWHZE8fBZC8Hm52Sw
Bj9Irf9xxzPWcsiG3ZUQ24fJQu1Zs5tvs2QU+L2R9qSJ94f+f7NZb7oaq92bj9q/iHXjh5fs6bhs
L4rBPQEhtHwlAPaOEcDJ+YzuRDx7rVelWs2l1aUSsp2pYR8lJ3HUzaaN+ETJUdDcYMw/G9GD+LPw
fVSQzpGIfmEGXLn6ssynsPxyXBHzIJ1k61vcq7UIUHQXgI360ftiXgYFwf7GpnhCElvjHXis84Hw
a5OcavTlKTQIfymJRz/aoTgnnjBRgaz238gkyYCCh56b9lnDZWToDmIAumuP1QShOYoVtMh2hQfO
S521V558zt0lsuXDFpENjXhxkG5VYcsJjMG3PMnxbbzYwQsTNgA/sSJ79/7CxvQzeQhJgjcF1T0p
tWhQjDaM8I1dA+NuS7Hs1Hd8GhyCflGq8LKl90P+4J70pEKG7pyi8jG8iT3aN+w4O1RC4CaUFCkA
RhgV5NoquwWN3NmvnJ3ZIo99cSHH2JbYoTTKoXnLyyJKSLwayU7ghxgTjAQNn3g+fwyYUj7/cgLP
SKawGScmuPJj4PRxCFbbVNzFc8kHzt9TC/W2EWFdHyR5jSPKpOwWydgggadeh6eqS/4Hd7cX9Mcm
tUq2I0NMguzFjLsqW79Pj+wgEsVuSl1qqpSbAVEWXoUOqrAm+bF9qe1EJwkvU00JLWVPngLDAqfD
GFAleY0jMMh9rxCaVoJnfAY5I+k8b2Nqz4oX+iXpjfYqu0gBvfLtEvLi33UVI5cBJxwtZ75CUho7
0oTNpsFwL9Tp4UGmCkAJQyVmcte2AKx8qrjs9kza7XSXdjDRC/1GN64FYz0xBVUlVztuTosx27aJ
NDkfxog0bQN8hZ2C2FVm5JfDLBCDWZf52unjVkIu/Mq+ptVnyIf4BI1QGtIGMCljHcsSIha5tuxr
BVotihfdilB7aDf8lg8Ize7nKL21Od9L23gui8mwaS/pKOrPcpyDj2O8AorcxmiHFUH0zv3/+t3v
jrzHe8WoqSrRTRf1hQG9VD9MMGIp+LGo9t6jBf+8A314aNZ9zvEmA5RMx68lznPvTb06cCGEYgK4
1rwAymW8KlSLpTxgS1DMgIernTXropAh+zq97TLAEq/xqLDz9Lk1upBd6Nl3dd5FK3L5zvzcsbf1
ohNpOWFchnR1fsDFT4zVfMDTlJ89lAQ8CmEtLZ10P2wqIvQq6AVlZZBTQQI/y9Igw7C0WxnNgkKe
InCZwC3+SvArQh+ApfcbA9GwCssmlrk8n0fiLRjUUdZ66RiI7fn5EkVxT5BIwXiZ90nV25Jmcprl
tDOiGpLlBLOnVqpoDY1oBkKx36ppNk9Yr/L1CXz1bpRLC3+0s8SUbN72jMTRigmjUGqD1kX91jsR
SnRI+O+sMGqb+IksoNlUCdTGRJEGhLuyFhYm4lzmXM8f1A31q+3dk0xVLkS3T0xxjVJA2l7tNZy2
LlPGySYS2XgLO1btm1xTLrDPQFc+pHw66bbE5S4fV7jd7+WBPjWi3EXSLl7tIqI4gwLjnXBtZTC9
hRy60znxnznL0vAVrril2GHVRrDsY+PiN0A85tO0Z5IXx2n6NOWk0erQmlWfcFQY9cTvqzrUxNnd
ot7aw4/f3Y658XT0u2BoMz2CnZTzS8wGjxyadc12N+kslVEbI4rzrTINa9vgcWPWck6I5N/cBLwl
L7t37dFY3rJEo0cutoJNqs5wi1XwGhrt5ObafgSbgmDSS3eveM7+Ovl6jZht7uoaxe8WJUfQDHpy
bBbM0E7NZgW37JwuCqOsOWpNUFanKs3awMQOfaV6mZDFSPUwj7o9x25GHivsJr50yvHAvsMuKmGc
JudF/+pozWkQ+svoTPJQMD9wXvx11H5NX229d2L3G8AxqyrYOuexe2t/GYoU/a8qCdhgB4OYQjww
39isYQoEYPY76qaMtzgIzEkfPQ7xAyugG9AwYy+8MpekI27Wx5PyXJF12Lyg1xFKRI2mEmmaXEmh
CwLgvh9CaAxC+CgFMzkGt/c3bF/LF3JCJAULDTcpbEFotvPWZnksNLlSrgL6ufDXDBzeKsNjfdze
yK6VHfoyb5ALWhGaYETYfBQO/s5FGT/RvBWem6svlrZUX28tDg5R5+K3nZLVszKcdGihGWwLVQ1g
tZyPCapycEhHTtvwaRz7cLjQU8/ljUU05MNBQMWNP8HUgcQhh2exHOQe1DhXI39XdXNtWNXUT2EY
kjwIIkbwyNaYyQ3ZbXu7jlTqxsLuc9Ic8WFHcwxiI/eED+0JLxZwJNjLb38xHezKuqfufQVSAdLM
VY7m20rCNelVBGXYdEZlo/N2j9AHBGZj0/ZZvZgYvSXzz+OIqJEiSzaAEzRnGBveEqSNx6ohRLuG
tuuQ5jooWSAP4WlPVJ5Bv7g2Bwz29soUBuWdrh2GwQsCyvB39HZX6keBqVA58Q4dB844S9OW6gv6
5Tpj6zGCU+54Yo47r3JJeHyGOQgpMez2kv6jzLqrejO329XXA6mnw6Z+0jd8sRKqtksKr1FZIk1G
apPOwbz07qxNAcuLSqt1Z53ZrM2mBbfXXCacSF0teoaJe/SuUCeCqJKw7BkSupZdCYS/SWHSK5hz
BlTjozFQ84kQlHQ257HYNpFFlw//Ot6Mpjou/ZFhBqliKc7JbGCnPHr08YqUaPw7fBLd2VrbytEi
wivunruoSdvDiBsKgD+/ygeSZ7exuxXmuw5hQDPnIjegtUcVHTlTOx5HvmuKzmeuTUMTTXWXlTQY
vkeS+FUjZYaMtCTy4hhcq0EGD/3W+w8gw87+MQQsAJfPviKJjpN9mZbXBE2c4G+qivs2PSx5651Y
xYJp3WWfHX/QH2pzA3fiKNxKE6/tlSyXnbiglpGkQz7t5FTtbRHgiTORzf+YLK9geR14rbYB6cIP
8wXzA11bq3eQGV8o8H4R1OT9Q9VkLZv+yNfMOpnUeSka/vUXt0LG8uSqpHo+Yuziy0TZNA5AlCKB
GbdnsCmYZfCfcBCB65aaKVJh7nJja2EnkZ/y9GYu7SM+rmo/04UOHOx/LnS9SfXVjrCG4qMfV03a
tjrxlxoypJkRYNgUlrzjFrCeTSctu4qJqyu0j7YfHYdTXQE4SsqS3PrylEuUnixUFj0eIAv4GTUA
jkxfktwA0ZKA7pTQePKPG1EHMAeQC3zGh0DWelDizO6okumgoHUC31R7ZrYabBvfn2+GEz1QgrOI
8p36RP7OF7it9vHZweZUU0cmSO2WelC9RxCMfob5L4BulgXfV/Za1x2ckr+A/43YInsQnLxuB+An
nkavEq6bwAzs1V7UiBDgwW++6nlHMyzrN2NnA2Gvokr3a7ZcyiEhPnGblQuf27ilrjSODTS2tkr/
+9zx+FZIRKS0Q+dph6obvPKPkmudRJwilj+0lucWELTwejz+Oqv+qBIwJCJpDGk/pl3oGzzIsQTQ
oQbAnxHxD4LXcTcWIRoX13F2YAGvQ6/raCyC17m43yGI63KInOhVgYYjxJ+Evn9UkafBq1ITnxUu
f3RzAuiUtTDdc9QXsu7+bNY25JHhyPElNr/ge4P9N4WGhHb2HbU6SYbFld6hvfjZe2F0wjg8x1ig
DIcmclA+EJK1IuT8Mv95L+rR/p7tPNKPJl3AvPFEA2+z86c5sDqxjpcE5kuFSvPfk79gysx6zeFM
r1B83GRILOHYnNzIoeJQpm9YBAf0bT7hATSRz5nKTdLFbrAMv6BCBVZgGi2rRdsdNViJnfQaCw5d
wNId9k4DlYzWH4GE0BNxIq86ounllFWQeZpcP/scW992xIjXL0W5ePANlZTq0KnVhPrIq4zfn+5j
NUyrNe+6QnQkPkp5ZIMC9seZWh2U3o7QK5HPUQ4jfDKg6+Zlm1PbTJKf44JwlO0t68l917KKgbk+
29DYXwx5xvJkDNF5QdU5B4EW6EYbJfD3/I6H3JsxLUKxRyBr2gQ4+LAn8mcM5C6BUqAIVMd3kSEM
GEKVuytoJF0p7yyC6d/3n7tQt7VPf425q9ybfeI9vldBUl0a3CxV52DmbpjGLUfoIXz/GWGnNZXU
Ei5fjfYFT2wZePs7fZW+4E+dxh83ADGqo7sUQFTvMFSHAXxXhcGdBtp9bCiETALMY1U8VIu0S8Lu
vJnIDkEOmjymigMBdjrSUPesrlbdgnQYBwYFOMkkmbP2TmAEUYJ62juloc+yj1a/B1Uh/mfU+fi5
qEAj+k4gucbIwHOItSZx4GwUMtkYSDEjhTeEaJWjlriuYuhkA5G9hZJpChQshSNBvArodXhmrCpk
6d00LYr+f7aL/qghnuEvc3plDLn/Xq+Mf/O4K1+tGN/B1y+WSM8uhsxUwBdBqGWOutVEyfpFJ2cS
zYLi5mjOhOcbFagpx5awn8gi+1S2EaCzv7f+3GPgnpl8f4ZAy2vWzTL8rotiIfGdw18KK5a8Mp00
ygWUF+SLYEPAts5uVnEwr3/jr/TywTK0CUPecF7PyDvygTxZOP+k3nsA1A6TlU/z1N2z3ZrBSkAa
V8NdmKrew/PVyNmdpb7WKLrwDwuCExKnmH08KhSx6i4xm9tou+tQpCs2ymnrWKc26IakFqEnDB46
GCzsTV5fn54jAYJHL2Wrl7PTkDbSRmbKAx7gf4nntC67Br+2RuVWFwgIYsiQ5btFyxfkB+g3I1zv
Jm5tp51/4jIrYC9gkZiQrqjtnQWjFE3aoLLVVA39JHA29m9i+XaTp7+n7qd68B5SNn73HcMYNMs7
SC/cDMrCNmqrRGGSf3sn+YuYxw/44TzeK0v3ccK48YodtC1iI7dS2Mr1YIbA1+/0EYRQnokPt8oI
EJsFk9K5zpwv4XdsNticlD5I+EvLg05z83BFPjlWxyHodG8gUqFcpe5lEaR2lI6gVfkvRwbGqnOM
LhDDDROrj6owRmtEZ/C+29u9l8V9Z/vLFZHTWo+C1F5jsBA/U5eLwegMGrdjgqRIyg8hOb4EjeFf
YlfaNjlgVkWRtZSb+96NzKGzhEXv55hbFe1XFSVDk86RSPOeqmO4hnLmoEouD+whin4PArcrTxwp
WcoDN9ZOVMrH+Kw/NvO3E+gNsE1//UycirNCF8uYJcHB8IsaIWiq6iEH4NqbUL13TEbBO1QNMYfa
XzrTUVNCoRc+OkxqOchbgpPqsxb+j+ItCok5rRhED+2lWGr8Om5qgdImwfuE5qjoiuhjjh/XpzSX
5KQ1lij2i+kr8O23lA55KYtgF2JoE2mq4YWM9xHpdMtpC59Tlml+OMVcen9TIHldZ2unBsc6p2MF
/NnIB5PBvzET5utd5SZS17PdOtMGZUvKt0Idbv1wHwe9FepjS7kEqjsUKW3zwuzD6CA29ruhpHvy
8Hb9ZqpCN9soRKFZNcZaXd146hg7XcKk3XPvuln28IyuI3+nQ8UoSS7PKtCL/D0cydtYdPipwhwt
Ppdqkjg2iXZc+Ai0BfX3n+L0qeCFYhRpCZT+zZY8sGGn9/c3tAyVFDyZOeMclryJc4mceXdpVkbK
Oq5n7ubIO8xFQGvbrr4cgO4BR/2PsEIBRaKreAt1fJhYZvuEWlhbqV4gbobrFinwWOAJUOd5a91s
/iC050cGu1BVZaRg0gMePQRkYlo3b1tdCPt7lQbB+HiRNUakpZsydqTj9zqUKCw/9SG/c+1W+L/O
YgBaPnuSYUjFJkvCIrNmZCnvou/oEo+p0d/s2KAqa5knp499vITazY7l5GHtz7Im/D9IcGqfMX/b
dliwQp7RLBBjUfpwFZarIA9coFbRG01EOSrYP3QQ4CP7OLdMy0aqmvGPKY70ulFsPe4yZ67Y0ln9
QVTH/UieUjAlAnII+uVcbgpEZbX5cgBoGYpOwre4mBGkYjKDaJ1fzSDDbPhJaBPKCb4gLdUyduQE
/9XolIPJWy31kJAaYUEqzZDjQIf+IfDWulOBG9QOoBi7uwOeLSzRlM9iO+rcKJkGhVYgiKUgD1NK
6M9pea2oimaWQWgJimHJl+RDK3ZggDIQqT7gG5xsgk0NG+50gk3UQv/AczvrmKxuFAhchOWSd4Z5
gOdYWcU1WHq9BTO+pG7VqlqEbZpsdm64h3ID0gWAeFIc05+rC/ggX5AvxHQZjjJJUWPwJsC0QYe8
DXy6F3XMvDDQDrXO82Znfau7NZjAYllPdkm0Ky/6HEOGWmfPmqoos+citqFApMBWxfESyrFQS9WV
gtptMOeOrBrI4M7rl6e0DioaLs8cm1lVG0Kv0hWDuxS/CNLTp+n2x8Nnse5w2CcY/5Qw9IkDY4oy
GoNz/IZp+8D6OLF2UqZ5Tpq7Rm5z53yBO0xfyL5wHBa/aTB5HUON4tjr6d7zSADi09sPT/WCXMYU
2Bd/YpBq1LPLQHMvqy6reX8P3RRHhZV03Ka5laWqZOrNJxJx/dlVk/chTpZ5vF6ZtreBz5p1bt86
1Se5HCK42hLpCLaOc44GWuQC0igOePXwTj9rE+SK3q5fy6a7+cy5aa1mtCVALL+UzT8ctc4hOdmS
Y+ImRf0TTBJQPEws8u9u+GMGdbbQ2rvfqCNyeXksiV8oVQt04/NxgGYvSd/7WTllOd+2gWEOe1QQ
tdpqaSCPWzvpTaDEuX2cu1AV5aqLOCJg/KjEUmeDp6RbFQ+o/mAL0H/Cl4y60WArtgGSM41Tc2CU
prx1FHgX7slyBaXr40s1awIT5+GJSKcQBkyLA3I8QSEL7XfZTuCOcKiLvXwG0z+ucXPBfoJztsYU
cb/PL+Z3SVaG2fczLXK+iiAfZuOm+2Ahs48myGBFAaC9sLzTw7HORUTddlEMq4rxb4dP4DVmA0GQ
8LI4gAxGM7+iHiBFC92kBOnHlb6zZ3+m9jsG+j1y40OgvCjKZCCXveMakTK3O8q4BXvKXw3iBML3
XNhyxyDnqTYZtpPry7ehyBZaEzCGaVHRBnYd9mSzcd5UPdo504E56RKJDUQYrMsLyCz9e/eTF5Ga
aWOa8CMvgOdCdHrif9tktBhw9ov4oaSFTkiQe61b2G9WVgGPnx8KYmU4fPoG4x8KGrsFw+ffnGg/
FIfSbb0284JG9jfJCFJWdGBBVD5I2th/yxePrhyxePHvL7CNIG78yil7o61qef6II1CTXpT5NFiw
6JzDSZTwwG56m66byMdOJo/K7DQPR/7OdvVZ71fekJJ3pOVrNpjzF07CRTBfeZspCFXvh/R5Wkfz
jBlrYjrvid12uMXXma5DmJENMXqEhJHSyO1tpC9HS80Luy5Xz8NNr5nDERerYE/IZL67BBmV/AMW
81WFHt81hg3f/hThvzTI/STrssDEgoHcqWipTFH5nkchQiQyR7VQiHKzbRrUvjv+kjFaXT/0hhgf
Ql2o8CGEily9hjw4ygYIEQQDDPnYgsBopIdmjAjGureFA8qPTn0gtOfwAlTqolCLk3Ay/zEQNDKp
hXvcJbiJSMxcOjju6yrnFccC3lNTUbbsoPY9aBFdOYh5EZfXD/+w9eT84SpD+XUUiYH1hvaOqSmG
KaXlGCNOtrLADSPmU32zFJ/ha9SvEy6XWKVR9L4hEy3rq772Tf4KDWWC+0bTG5xytfmkbpqQsD/2
LFJyLyOlU/786N+R5lo0yuS/lCIuAractGsWQm2OJeVrxn7qolCNEXnbdgaS44Z9RMumc1d5XMCV
Kk92+wXqFFrXjbRsusM6dxTvAPHBjtFkhlruAs4Xdt8R8kCPRYxcSj5aWjpwFrd9JQMx6RYjh17U
HKOQhLVKsKMA4hPhs7ZD7HwU1Enh3YOpVSWguL9ioHmpwdiP9pfD3WAnqMWkFsFx5hQQSf9GqEST
WZ0vappu7sBkbLQJRS3/8pRWiLW5Z5Az+zPWvknYSwsVmhtLGgGx4omCxxxqe7whvhcmr+u47Pww
6ZgCSjHhNx/33VhUXDDQdecpkDgN+atcS22DuO2+qQRxzb4kVIYgjT5X5izCZbPYYvYon4jwTjHD
BGpzbGFGPFcZynzy7R/8EKWs+wXbXRW8N+EWHS9V7o3+IZqKFxqjmLMlEqNlIXHPpezUvuPzCtm9
Om7xYjBjtDMRF5JuNmmauZceFMQt9otFpV3LLkxwgqenuDNBy2UYGpxlzbGZeiAkm+bFwyxaTHJ3
TxWA+6GFgMWaHJOTQfaXMC9ZVzAenyhRFi+yUGBciOXBB8N6w4Hc0MeJpN4xiNB88HOY/4+TkgEk
MdadH2Yw/NQScTkxlTCgE/fJaNeyEOvdLwBqBViorOtXhIS7AhVgCBMtV6kEdz1IKdJJNJHmVyTM
EAMf4NMCnzFMNpkyhORQdkVZmg+TRvmTSNnxuuFENfPWIls8pr/ouJ6kkInHZD8RQGXeBJgYwiTq
i07Hk1UVMJgWSeSZUDwKu1e4TznHPfcorAA8K88/9hxuYAsuKnxpkni2zZaAaBdmPKfYGl9T6HT2
TT8EP4o+zOP500PqkBQpX47HU6y8EVa+5ov9IP/1PShYWBKtUboYKmmsd2gVaCMtrKG7iQeHXi3o
4VhyJTM4VP0w6R3ag4ue9Y2lx+OKd8EKOumNHcF1IP05Pi9R/ZkHagOrL1ItTnXPij4YIziUuvSk
EWbZc1L0SjvsJ1BgD/yvnUcK025C5WqiS4y7JpdcZWFI1uInS9VcUfjMwRJPXszPNUv8cn0uYzHC
nWzpTXtHkRPGYzpjSoXJ7WYQm3lJtuYG6CqKxpy97ZrICIK+HIFUNG9POXSIQnR8WzFZ/8aqwgqS
w9fNUOQbbZvtP2ibhGo8Wk7TVJMrvklXaH0kaaikdTwLNW+Iy/9uJjArHIrq4cqC3t/9Np+dZwAu
DocaC+Hb/uInXz9lbt/Z9Vi3SkczLM62N7ZMVbXuia1qC5rKuyVFbv2Ren5IbfPY5/sYWdqduwVN
5KD3ESqr348tMxRwG0C9XbNPUzJVoz/y1xlxBZsNatd66DyQlspeNfF5XUAPO04u82cyAwx/O5KZ
J1ByCKxUyK0aqTdJMZKoo/x85wzpWHCUD0Mad5J5NEbTba1Bkj7B3txSrecebwuO4xmohnWyLWGg
vr4FmnVHnhs778wZLoct1yh9GZzACpPW4hMbcJ0erTPWHmBdZuVXvfCm0viGuMVUBDzkM7HiO/j4
U6hrf0Ow+XJknQk1KgA9GK+49tcnmnBH1PgGglZmowONrgCDfQ8qggd8qXX2VqEv3WMmDsIpCbpV
KX0JJSExshNY10LtVKpY1nq2Xj9qppp+Aw4f5zFVD7bH8/vMf4lItU/bRxa0hTAqw+LXaWw3W5EA
86lol2lvKRVPB1gbtTB64u7PREieh2hbm+LVLAAy2Uc9aEBgGO38f/0RdbLpUYiyAQNN38/bsvAj
UxC0yJFKBb9zwI6Pv0gLybfXmgTfjQmfrQrWtczx0Mt3uCvwEnLcRFB4VkkSpmLw9aQFiTjr40o6
zeXbzhVYW+Z6TSTnE1hAncbUuKjZ1lYjchxKAXOWDuMCAqfq+0dUiWKvsnlM11SeyLzTlCPm3Vkz
pHWREP81aLloZkhbqQFBFKR+oJ/f7eRqAAkjuxCUf6SEwzcruf67v37EcCce/r08JEYYNIXVoQGA
SVOYkzVLxfBhtaBchvR4heh2HyYQga8WD+Xp65MwS7lLA4p5JRxavuDRntrfdKSj1rb35o1+1nTC
Ve2G9z85bDP1dPELPDql02fZU5sSUkU20X03DxqoRPRuQYP9WnheeBOobeGVnQgx0lEmOLgUCFGW
tJTxUyx+RF38Hrw6AQiUHk2bc8AOFYChKU5ravQrWkZmcxXr6LaeGR1baoFeZI3+vZ7+8nxvZUe0
cBTM772cVOOM30pyoOLJmKAz/2nl9+5BfC1Yel7B10VmYKECcq9gEPKMkk1YXFFS/Z+cAQ3bkNH4
9/S4/SAS2gNByWe0AInjVZlRWDQIDvXKX4LlxBoGpDzbo5fcd3YBigkTUL74YTUHdaEtGXh/c1q4
xAGo49+u2FswJ19nQq97jYlBz68yes06x7wrE9Sx2fm6r8/qDx+dZaMGWY8zU+BDn6GxJup/d8TZ
Wo/QjnNDUJBlBoAgm0FYkOmqpSYgtmDMNLRX5cHK4HwNB0vbW1cktR1vEQWu7tyqS9eHz4Uhml8Z
AnpjxT3M+Vfl+JoKw5qs4XpXomBeRNNzT02zLapdT4P7Q7r395QTe028tZ+z8DjmuYdCgZFkcWKC
MM7zNg960gUgAxh/YM8wW+7YlUVPyi5b0crBzxbURSIS1L65iv2eIVtYAtAVhisfTun7l1B5AYQP
xkNKx85+KVv0qXx8FI7Ffu1sbSVAjG61mdEfdTbrazzK/wAXVz5yZyEl/TLi572asrH+wErTsywM
6uilqDKlmsbqIBi7CmJgoC77mRuqxw2E7NoKSCDheblVMp+jwImAl57GtGr5tD3EUIP+qNPhTWgi
uvSZK7jsX8QzT9EnRsDOjgyclB2lDX0jgyFDXv3sbLyAqsExSt1BIwdlfHAaqOU/UmHEChd0P+WW
EZQNrrNQ/W29CI1dHbgjL6coDrG0ZiXnUUJEwSk2NLa/xbKvIdz8Wnjo8Iai5S2zz5yHjA0iloeZ
mEr8QsYPC1gbmKyRgwCOKvZg+wh/DyZ2gUM1JyZ5g5eByYaEdAjBG30MeEX2D7kQOF5G8KFxlUb9
1cL7vtqS5y+W/yBfMOC3V6/Nh4ATANQeyg3tyvnvlgl55VYfCNVNpBG+8P3TucaUaaBD0WEziwHi
Gm3iRRTYZYjHhZuUYGrmDeFUZ+5oa1CAX9vQfRlxp0T4hT6UvHWQK7LXZ8x5Wp2Nw1dxKGwib7/S
DGcLp2NF+esmWzRX5dblMwENlc8eEB7lRG/6HTMEQNwlPEPGoKDtwe2YNKF8UQO4EiurhaNlwJcs
ZRL2RVV5OeCaxtpbl44kL6Bdy73kBDLHarFhfuzFO1qEy+mi2fE/L70sM7M/5UZKozuZnocnNs3h
CgQ3awaTZbZ+9eBF9Q4TY++bwI4eHLQKDW5I3kzV8aKOAR8wNg873ptC49rMk43sS/QlqxcmXgSH
DIgPZQAgdB8SfF2cB3CAZD1JIKeDvGO0T0f+E/bVJXT5pXJ7hiTdyF/Kaj692RNrHmUQsI+kHpuE
WvyG6+IafOqvQVtNoaJ5bwAZjTMFfJ6or/iJyFugUpsIu30zDylgdP42kOBlAxMSg8NnWCOpGcjn
lLEZCynsXoqTwHX00aU5MjWKW9QwWq5MgLqYGammQcwRRFlwBVlw6VKYO2AlFTW+gLkfiV4VtG+4
mnX8UPRzHQbV5ChpH21N/HVjmCHKft1eaNY1CPkzn/WOrUxDZ596VXELxFcfP2T5XQGj6DwhvDX2
OBHhWTHhwQW0RIStQ7eml4/i2dZCKcl7qr0Em6uvqV+O2Xj81/knnSrR8NCAJDIgMyPDQZHKxPdu
8zwD6kEOAydwfK6wcFqVU0qM5Sb7mEIT/Ahm0XanINQr4RodoUVauA3Kvf32n90KMbguW1lHliC4
/7fNbbRmqfwh7U6YIrBuKGCUImn90UqRVz8UnGltCdaDPz9YyUjxgJO/dDe5AmrXxdQ1lDxvw1zP
PhtKxRUOv+DLumLLBkkoulprKRKTRAEJ1iz9PjtFpDyZh8Rm2rA07hDARvpjCdAh5lFmJ8P+rxTv
wF3xCI/PQM9nLlf6rBHb5lDdIYb4ePp56IgCc2DKrkwN/CjBvJLF8E2QIpJF872FNsBMKmoZAcVQ
hAFlZJs9PHbM52ZDn3YqcFiqbi0LbpH4s7Ze7z7J9aQxin+l6P/C/k6RfYlFuTHoOf+gcmTTxxJ6
fUbIU/J5nEPQSwoNGMpPwQh+bip5s7uEx9SEbIZZCdj3rFbfSdE3+ZRoW1eIPLF+cv/zVZHIyURC
grMSzAt5qhINbS8czdTRRDEVdhvr2jaIGZoRcohWU/MKZMURmFHyc9sgpOi1GHyBcWUXXcXNKAIi
/3vIK5KKqibjF54/UoStSOYvdbWV0JTajdd3VSuGaWnOytQOieEEhcQbDijuXQ2ntoECAWDWHxzh
KHxiovAGI+DGX1SaanHODTCpzUFcUiIU/IPHGEHCQpk95vTvXhuQt2FEJBU1PZNBHXDboP9n8si8
mKzmCT7kwn5gs0mEVORjKfxEbLPtr1QpRYf0vZf4HLmluhfuHZPNUhgG3CzZlKNgZM4aYstyuh7t
X9bjDHUXRW5LDVgxFD3ZrTGiKTTmBj/4D+jbyvS0Dv6dKPrTWgKTCYXKOhS4Qa+yjMWM1oSFXfvM
+AbMVMme/IKqaTWjjOGKTHbZxFP8Kc4M+Nft9+2MegjJjl5Fwj8IBmYrsfAiSorjJsYzGrb69ybT
4+vcO8UoC2INVKLYuHa4tQhCilMswAzB0TNQCrcCleeOYX3UBbdBiL3O3QvbLtRgmD3wyKi07jOp
Xu08/nVMYHMxXS3mFmr6ApfASbmR1dKA+veFJhL0qqDylev8qTPbjEhl5JhvQS1rA9Cc41MCucaB
caZaVj5qm8568og4QsJXv9FcdIRSkUYU4FSC+9HuoruMnSifa6uN98Fv7e5vWx+NlGLS3E0p1b6j
RHepksSKCVqWQwhQlVn5/j1TpibyuFQwxRp+nDpmoVYlC7xjvsDvHiniShbjt3YNn0mbjx1rgVTD
m3tUpVGShts2+VH9Q2tnGPl8HXr5zJk7knXmVKRjvnH19BMLJ5wnrOh9CGMETMkxtoilmbh/hzNJ
JnxFoGOPveM+xEHULCrmhO9leLd9WDb+yMMI314N1m/ed6j5HTvuGQF/7hQ8mE3M4LdMD8kM/Lvb
OS1TIiGXp+4hPiNYLIJe5tbxsOkn/sinqe8OqXV8kZhTQzw5BfsQ9XR2Ehco03yyECYd4qurWFaO
SBoOlo7RIafPetqxDGi92j2uxG/fHm1p4KufTeTnChpY6+4dTMwtj+1l+hCyGoonHp9qVplvfzn3
kc1A82plzqmW4CS/sx3kQ4e6M9W6Jx3yd5C0yzv/zuMkpCbdofnLK+/fLDvuyQRhIapyKipQ94KG
Df6CZVS44QKub9Jui3Drn+L89JhVZxWb11yQjxZTQAXN7J1Zr83NpYkFQ4Xh47LhvsmmxVh5aeW7
FrygOtynsavCHtigfJJjTnQKO2XKO2Zqd2roMe2zoRTjsSnhoKdajKYiDtWX6LdUiq0FyxBRQni3
9RfZdxzo0kD8kYKcEaA4xBVFt+AdETyN2DCDZQffjgfzOYtlJLS9gSyzw775uAIOfrQmXYfabbdX
MQhJ0unWMaZNZ7oseSKNWAhFodlWv5bhjtrYDx3IrG0z4mB4fQq2BD9L/b8T8y+LKjTQYFv5H9dt
6ZgLUvCds8zUSdMVaM2SP3HREcnzPxkzNuRbg0FxjZrfOwBtzTn38iDlc/7U3GdWRSgxqKUIhQSk
jBo7LsByh1aXAg6G3CjL7WDE93iAR92WHsnlxRu0Ww/PgJZQ6oMQhD1avJKwaTumNcCmzin6XdsX
WFNtiz3w+0pjjY6jSbFAh4IjusfU6QTrEGXWJr0CQpKUnwbMYBGZIXKJh8abFo2j2q/HJns74bMQ
tILrDVaax4NzG9NyEq7vmizNHwyr8EOmT41+qslswwRHmTTkD0Mg4zYVITRw/GQfO3xOXp14zE38
hJzjZwsEFyxabfCXzPd3ygTrAzMh3chErvFLy7ebdxMLQ6w6jqfheAHc3M19iWC39qZ1c7ARChmM
/3otHsHN9QkKGp3PM3cTUMVhKlky9PuYQWZ1s7wWVV4WRx7r1yvAcKkaN0S/kQlTT/Z7BlDp357w
vDFaFz49Cw3xla5RlvZDs89gP7PNSW+C4Ag7eBiEkk3cJFVhqXohIvSoSHLbYdjKWPlWpZOEYH8Q
v51VrSseu3Skj56eil1/PUBK8PVEmecHTvH+bNdcHIIMaFzdA4TH9WdIOh8UBpXEKnYDZtPFyD1B
c76Np47Pv6bLUK54+VXdGCQataXkA0YfuvLrmDhhrGBO/5/nl7Frn3N+NE056dbI94YazfWNriBH
rdRUrKgJZTOqCqvlRWuNxW9wI44XXQJ/0v0WzJWqa3rMaTQ+U3WGuGdlXNf1gGDfkawfmK6kpKDu
CfUWUGjnT26qRmxvjGbP8CSUTjN+3UfaPWjY5OXCqlobeywG5APS3fkrew66nin6ccfdUFuZ3vqm
P0KuiHbKPJ9UvbbLMhwIlNh8KR1IcNUSr39LrkxBalRQ3OutYnLqCoMp/pasWHu6MgMQu8kBwOVN
UAuwm/dVWlG8Iuxe2majYWPOLZvMHDKbVadVZ6jNMgNc4acj4H8kfSgvvpLQs4fDA0YXZOyvlgzX
e38GsGIMKPfSvPLg314vyXf3CMp99nm0uxv5E+gd07vs2UeMyld0gZ4iWVp5UO+/VYcBprvpNNmh
G0DWeUip6Z+zWDvCLldJpJgpzxrhH6UDS9ShTpFpJDG0kdbmRSj7AQF4zEK5cZBA2jcK6u99us7/
RLhCSrTs4x+d7rQ29j7nbDrRiZaXh7E/+gGPL2EXa6yzq9lTR+qOoxJENbll8mX9XLChzA1u9xlt
vj+6TGEAWQ7YPjbUHoBbIH0bBDGFjxMQsy2lUX0PzykWSXmqlWZKMAd97te7XKUd4CvFEKKAjVdW
Ar9Mb4v1vhJtd3AzapjaHdp8JlD7nAzmdqXnTUWQ6CIwBjhv9ij03Q8SdtGsLDgfIYKKjZhcrtk/
V/5KYVdag/5w5nA59d+5pZCo2dberqJ/F5xJ0SY5SwpHqEA7ZwQXdr+vOFLsbNFqQtF1PHHEaQUD
Z3QrE9G8vlOa3cwbX6Z2ioe+8kLFj64bW7NViOWpUDoJC7YCWU/djjYtRNQeNMbEJQCQTIvXwwb8
vyTyt4PHHwmhDF8j3FQSmUm3Pcp5CxL/+Yii7wHPgkO1NPlI33vzCI+5gEqkdfSOjTzaJ7W3Y5ej
/vOnj4UzqHtXH2O/QtV0Ez9hyyimedZisIPy6AadBm5F2gdfxWN9GXecjUUo9ExklakWBGTjt7Sn
xuO6U9VvFodkWnVt5eL1nl1q6AGgMBNjlFN5OmReuaBsMG4jaz67FhOFjNHaDcMnWAN6TsbeIr3t
sWyMN1bAyAryyXh6lV/4p4+EJ/ww9MnnJiizWnebQBYQ63lzvewVH6HPFlCpy2r+zMk29xj8Sqna
pPk+alj6hPA03mKDOaAQ12fyl+xAMwNjrYI+fG7J7yYZdzb9oF7LuPt+dRrMTJhZBpugy/KGBesP
uKSgYsXaGMffM6WFH5y6s92V2f+5GN/wjCWIe2oHAXahsHHTDwEcgoJyYHEe/KFmyKXVDsCXXx4Z
ph1KMdHMJMVdtwiP0lDkmAqMF4tdkY2saNqdL4J4Ikq9OGzAMsV7dj4VjYIbVmotK6i22DdyLJw9
GeaBFWE9aMsFfUv8soJ8d9KUgvlMSIsc8K47Tg7bFCW9hxE8L6RtiNqz4LHpa+M7Lex3V8fRSt3T
l1FJzicgupybbaUfX9iA8U4iDCxlX06xqg3zQsoYxxN8jvMNwRPx7eNAZLg2N0DhO9V/mj9amIBv
tnXUhnrHUOmrY2J4GPAqq0GpihrPYKd4vXHOwvvnjZTMMdQ7gm1MxP/2cQsnSF44mog4S439AsTh
w9aPEIZI6YZ4gs+7m/Ylq1dm7LuVflC1D4TC1Cd1ioEqFVZOKBEEeJIIWEwO/SegKiT6NRgWcQ5F
vHn+46GfsUQuo6Es1hCpuYXt3GX37uhdPYiP8SLz0S0Queu8wAT2HrEUZv8eGcqYgSawr1jD1V4K
QyaWd6acxkbukYxI+121iDMxrxljkUFx3lv8VznRMlxeuv1n2LPEBY08Ar1gpE6Z+Rfj711i6Wop
422+OQjSHEhTjIVYl7wRzo7Ms3KSQyj7tGW5Em1Gkwb2YohSm9dyRL/qvyi4HOwT++fW1uYHlCGM
EMiiVkJr/wXxGfYXDl6BmcxOnJ9QL0UUi3HP3CYoO8cdVSxjnQSjDVRxdhWj7rkQ8lDmQTgerb+o
yfFy1iM6NyPYP3wHQsgvthA7unR8csuwLJpJqpBMMsAa/TrUDJ/kderOBUsCVkZd5tBk1lwh6CE0
M/EYyuQ76W7zMg/f8UlPLU+3BapXP/YVi4R7gCy9K9cE8ErXAcEfHOHtRiqevMmYTzPD8xCwnI00
zwumhGCGrGTyC8O4waKFQpouYQbXZNBIUur9MKXMec2YNgXAwqJ5hZkZ+JxaewGqtTvgU3byCZkf
g/ejtnQlylywe+uIJOnARIE8fRWIrrzgloGrj0ENcEK2J4rdDnyqsdi0P/elsXteTocKvQgvmNx2
hqV5SBYyEoyH1g3Wvdz6QNSWJARh5Udn55yu6RZCyp2MUhjsUgU/YUeplcRaOgrTpMmOQo6rLIIS
bmcgCwF7EKh5NBhny3LF/HA/S5KDxZafGndtar0ly1gGBWlRlx/fz5fD7zYgh2vii6SopT1bmjf7
kXVgTtoWndGHooEzh0Bil8GF9rqf0IO58Usv3pBxJ7kjyoNWMaRjZGRrYK2YBD9bAw/87J+SWr9E
J0Jgb+MmTWKKF89D7g5pmTDgiWA691DHJali2/0FScr7B50Ikgyoa7K9huatFcKHQA/aD8YBG+bm
ag1L5FaWWE6nqH1uiwTBhgehKY2Sdrh+xdBmqWLEgaGYcQKuDRz0CCoDSGUQ2xQ9ex27Nv32Xwk1
E6YV/7DfVnD7YKbHVWzEFajys8NUFCIBBff2emc4yOumbBTn4fy1DaH1NelZj0+hu81BtdQhyMIe
dHOS6SbcTBE11aw/Oh1ZXfw9RyXR5pZDXMfJjUsl6hxxFWon2UGvPl03xKKkLERxxoBuvSMd2vDk
zm8ENuUrNxCWPPxBkiMZz1vfqD0Tpz0Kju1+XNu+TrM2G6maohbvBVkr93y/72vTtc2kTccEpFwR
LbQitsmqL3y8ztJn9vpX3mt9pufqGJU2O2kCclvv4YX531oLuDCgs4wPdXdGg+j3ADXZy4rAu1KG
5q0dOaLELZyVl0YOUkFcssCQGLnnJDvw3gflo2+UVxw++cqDGVTbYkIMgf6zI+T15Ye0dQHWQ7g2
hCWlwdxMopETUbR5IyzjMj24jJ9hOQDMnaJ6Vh45jC8FlVkyBrQQpW/21r9z8QNUJUo2IvQs+s7v
+B8b0tmzoEvcuz4nsJTwfUAAzWDRTZfjn4UmOgzUff8lEguFlO8b2MUVriwM3pxEBE/j2oGkQ17d
5yZHhUZQnPTcfCeIONFJu+miApPCBUGxXwmjTCiOOsZsFJyON+QDLj9J9pfRwCZ7DDY7JQZUFrLV
tuzl521yF7gV758+Sm0WxGsysqfHFinY1QcNRBR+ScDaLpxpCmqi3UICQH0rM/d+U+kNeL1MG9W/
zG/tm/zlQWxMnEEL4gvyUxvSMY+mCZ+h2yAuo40GkNazuupwOU8ugkm5qmsQWIuCobJpGxzhknZG
SlqyiGWF/O5FiZNOXXkLxB/G6CXA8sb+5pL58Ig8nkJ9JK/bTsv3X9jq+79xQryPv+Cu7JZmbLT3
1qab4ftvLnaox7v7eBA13mTpP8bv3YhZdh0H9jo8TZYS5ZEqXuPNLMav1vothvSNRJhDVqariBXg
SEK7qosjT8Yf73ta+YpxTUUmrcU0WsnBQE4SVnF7eVu7yjMqwtNilld3g76A2pnVMf2sCEzHPxei
s6nUDp2erNhQPqbEv5uE32yPB19ZqWjiVxTMFZczM+Ekhiggmraf1j2/jhP3todqijxL2LHG5SNX
1v3PaU2K4jnGc6IKDFa4mBv56GyAVqYmpxNkwd12/ii5cmggaUgNErwx/Q+arfx/o287zFT6TECF
SNcK8GJj51dvUisjK8K7z2Oi6vbCsFEFm6yWMmhWNSLmJuUEUOL8FkUes1LJ4d67z30zw3cAqBzd
eVHD17s0PyqiKssu0/aPWihXV9dYYlkpC2k2u3ZDxVB96U+Jsf1Y3b9EcDcslzYdCjiS7a3O3PrM
awgE+hX4LixWr7etelV1cvB2gj6imxWvjshcFWEawcIQt+O6K9T0a2kaqtO9OXU/nRGeHksups2J
T5xdXNahDc664wHW/x0mcc58znBCDmdsfqCl+OQgSjLHl6CKN3zpaXkY1ecvUI7guvVtRE7RtNWL
HoMzfR7WH5Wrh5WQHJihJnQVX1QfZK7bsgcBpeTXh0DcAI0Kj+m6e3+4p11I7u4s0glfR3dEcpHe
zkvSurUsDgsCrgfWMucjGLduyGTtMmNHeJWiD1rnY+FdFEPEHPmyo6XjPABQ12RPz+zxf5ImJXHB
GEyfvGyw7NZWObASwUhZpLZffEIH4SwMB0LO9mAG6rO3Cr7rl49ZNF5RSH+LOQZ5LVtNiDbn4ynR
Vpwe7NW3jI0JBBkciVS82muj0iFDTFkcysKMZpM22qgIQYYQYmrCGXyYsv3W750jZVIBZ2PrXfqF
2M6V6NGiUXreY80P/MsotHm1YdJSZaVi6db+Q521znB3rdc4rJtAIsCpVSCQ4pSpfp6ckWl1sPvY
bm70/7OjroZ2H81Owk04SeGZNS8YGg0hqkDXMXJe5DrgiEokdLIpGuPJgvv0xNR2Cy+jQAxCbmJA
Y1G3ht+l5iLG00VNNNUXrfGg9cUite7WIApC5hSYiztbrehcvjVy/fWU/lkhvBxM3HBmCEu3MgSm
EdV5GkEG2wLvkQwpuvh2/+CzY6S7OrmLo9/npgR93/yh2aVPRmMzwMbLWmuAitU3TN4pNgKHtm2s
UAHgN9O8NGJvTFaooxS+zX+srOLRV0Bwve0S9XTWn/JUAkOTj6zFk2sr1VuOEp7uYClB3MMKMDTr
eaQvYjkopeO8klJuT/4gk84vK8f+YYPv3zdcLlTCOHYTufxst9LNmpk+IrPXohw8H1Ej6dMQYoBl
Onb/51z2Hq8jF+A/doOFc0BkOjruYgDPNhuZnDTB1uHhVxslCu21ZK+LpDW3fmuEj85kxgT6SoAC
0Pe/ndpzM6AE6USjG2809MzN7RTO4UFGQNAvilSIGh08rg+uEtEGvBz6/xwIT+hAgI8xc27tWZ6F
/9q6bboDbl/3PEkgh3LBnygaG2pFjhZy+6WAJCoa8I/WoQn0SjDt8CGKkh4EdqnK/MVzbrEYV8Wl
2aDStBHXuYPx6pF4bsXzslv3pTjh4zTPFtrG3FyXQCZvwTsOUievbmLkp1I5hBNpQruaShfZ7pBo
5QMobhf/YECJwGRKIpLq+TrC697tkI4HfMOtqlOmY/pCxkCPl/McC/O2KhF4KzFoim9v9UbRUR2M
WWofuw/riGubeBX7t/xEs3VVpZEf51ppJNYNkRweBZtayZ1TfG6QvZzpNWQbDQv+K6txzFjy8MYy
uVdGW9ZQypQbi1RSR5udcj/D8Mz6uc8M1pFKza4P12ixKmCSWhRnorBLW+m9T8f7ZypyUjgZ+cIC
YBu59TZd69wwjRwrhP5OAADvF0qpcqr5oA3X++oLulICoZc/Q10Loys8x3N9EIhRirRuaiN6X5Wb
akzumkJypEvzJEwxJzZeWN+cQRLeoY/Gp2DFIMzzyoXaILnI8aI/bOzWts++GurPCt42LoZ+96SQ
nMeVX8BxYdUAVV4IMRzwOf5FMYr/b4wVgl+cC1axkM00yoJnwiWy/4BZfL8pUeA/jg0pCjqlsXr1
G85rH1JoScUVHTMOtGk0ausq/zuDyXbvCnCrJgm0Slia36hRgdQSfB01q+FLuQ9q3UeiBh0FIFuK
YYwlGtn0yc0ssOj9e6OXzwf54094SIOKRAAW0lB6kQb4IWguHFn8TQNf3MeXvPHAwmQadBMfPbq4
rtopS/7nQ93V5glaQCqeA9WOLQTDtowj8wbuR/yiqZF+xCy66ZhjosCh5+zzVauDGmK481witwXZ
rFFhmoOudrJrIrTG6tJgpIBDSR5ky2/T14V64pQ4C316mpodc8cMhuQrFoN2RNQHYStzV1ZNzXD7
/vlHQPX8PlU5Ty5Qn0R+y2cSNkjmjgsiy/N1/Aes/Kyfs8el012vxBZFoh50/rklgnDNW4il7aBX
DiBRAqtBSHGkQTgZ2KKWCtAis3afkaxW6ToL0HcZmq1qX+RGhep2EIJ2tdeb4AU3gncGkLOUhNLe
Jpuk/LYpXxDKXl9m4sgu/tsMo9bv2DWWMSqxbIrnlCUy7V4VPqw9Lrd6xjlxvQuCXpyRJHQszqyf
LDO9Crn1oZRD0I+drMfmujb0Vr+HlJK5RJb72KdyKqUDzP+dmznEak4/kA1Y3cCSoZgchHqTaA0z
VoJaVGdDR/z8M6ZBxVjVOeVXPoMzNjYOWMITL9C96O6Xp/isTIsl2j3DeQ/C+Xs2FDHknlxvnImz
20T6uZhDCApDWauMvMA5dTkMaCMlBYAzFS6/v6NgNWsVAswQnncvUaJKdSlxrRZRn8xY9yjWPBVn
1LIKyYtuH54s0N3kNzP8xXNAYnjuJCShzgEODhA6JoQXKqndTf30ftofHbOvuZ24V6B0yExyrzuW
nO4hXXFkOmpQTzay3oc96sA0jCPv8WVthmbXELCpOkWkgvzu3m/3B73cppY69/HfpttaiU9MBL0k
uiWbpLbwWK+Eq2hQ8vV/pvwhnVyEZ2jcrPyHiDQSU19efsEWPOTqLoWs/BWwpGqTyLEM9MwI3gz7
UDy9YOR55m5jOjx6Gqf0B05TVr6haqhQgdYMP3sqlnqywzHL6O/NKXcxXdF4KywPyMYw2Ryh1nQ7
sqRBKztgvOxFQWvGlbRcTWdRk99a59uSLH7934Xjt+/+X4LJ3LNz+hgSwj4Voxz8weQiCqVFOBAu
X7bSaxj/UPHmJQ7GkGFLTKPXHuuKc6k9QiC9ZOcK5INYACkLFVAHajdCJm2eYK90S2733mvcaJci
s1XGmeX7SArNyZNJlZE8WgivHVJjBJ6efFOAh+2QgZvv3PJ74WqzU+KI0eE6H12JJM238CP5RIoc
J0YSkyU/jYWKZjBxt1Sk3ZjlKeRo7MRYy2zBD8tMq3myd0tQMAB8Tui+s0Est5mrhikPHlwNRILj
CoV+/77qDg0ucsxUQjpyuzPZYVhbQrbkuyyRRuH86SUUXrGrAtbm2A9YoXkmJOU2uUzunGiGUrr0
+GRlUSwon3u1tgZ5RLjGSnNjKNo+Lvqf0+atEuIF8Kk7mnapEiP8+gDnhpx7587Jhz0XptJbQTff
lPQC1d3aHrACYPExPA3yRHhy2TGRXWXuRJclKbcgkr4Urh5sI8/bCJVfqJwTnVRikoAiPOudBKcU
jEEb+dM5m1U4KPX0SBwwgAwFsRsB/YWoHRA82fELc9XR0r444g5Dlamr+He6S/1h85r/wkGUtkQD
IxNJQgt1jCUTA0tNiCDmmAOebcMzkfeHh7ezNn8tc1MQcBmx+bHOXWJCxNbbK8tOIPobpQUxhkYP
LsPnRUYi5rcfGYMRaobRsht047uDGbXIjiqqL/edCS+JY88F3i1bB2XEBwlkpkP9kKd4dSZgROwg
ERlyMEFfxRlJGD0gGuNzutAGkPBm1pZeZTnLImdSJN1h0bdkm5L6+fxA7L9PziL3WUokrr2g+yBg
R9kT12OL/vDWSMTM9ye35ZMzixYOueZxpTxsFK4Ulo2BiFI6402W/HwPsWCBT9kMLQc/Rkw+sarR
GSIN2PsMn7Wd1cm2OdEP/Mpqqsmj2GP2hwFL5vVk0CE/g9IRvOBsCoRZ8ROy2FJVG7fjKRsUsEnV
HJi9MDcflQusAvSi95rfIfZ5kPxHWkA0Mar5cOg5hjgGvPctSYIFdmN8L9/pRJB8D5J+LpoGDQUq
ucwUN7vt0Y2VDvwtfjP1LQaCULvGITf+bNTcfhpjN0ht6yBDtwXNCXmR4XPhsPkVyygZQn4zWGxu
/oLCqs/6ysJnX92+xgwGGWtjUB8S3h+YJaIlcS05x9RCO3AySFfs/mh5UctwnS6nwIMai+ap6oY8
2ykUXlVZcLSsZ88O2OTslkNmzmvQFounbbRVuXRaurP6fNymUw15uTrUoBObQrGaZ8Ls2RkUkl99
a6Stc+bizbwdab9cG7i+yPeyTz5iPrFJiJD0bp1Af2U+/zYgCQ36mepXM73/XcemKcaexTbuYqHG
9zTEYwbPzuPnM+67JxCe3OuNTZDjUGBZ/XubDEUMwvbW55kdyhj874LI4WZJK4uDNvYjZmNsGdEx
ZmHcnTrok59GXdsIPlPGfu75ZIIvBOpyLtd328OcEiVUIcyqQJTRD/WDIzvChvKdbeA2xfMbyW8m
66KE5evmWFOPvHn2PjUFUvF8lULeFRb0lwzW2BQ12D+OP5gYTm44gjAw+zW3EeGZ3tQ78j8StyET
KPf+Tbh2eofxe+yz1NdqlsT6wX1ZTF5iMvFWsKO7TDdTa8ACpeMtZoQCJVSn13/r/WXFs0tkpCNh
pyb867TlPQINjOykiW1KR769UU8abH/a+Br9IdxG9W+qHFsuAf6nCbPRf5BILx5a72vHs0mZpWJV
/yJQVr5mpzv3VE+OOsEOOidWsq9UchrhNLZDmPvq5plOynt3u/xVSk2feQ+DjZQuU7yaPSuyHqZP
d34x2sc6md2HX9X2ozadh8rIX5YPhp3NwUncW2y7mWoS75TsvW7mjMPOXHIa5u7TqGxGTcKv/MGk
E9UJG81OtQ5Eyg0nULSHaCSjIYFRM+0j5yIq9yALRHxm32fQetHPK1izj2G5/j97/o+q9Ki9Mtyx
yCJhjWd34LtLkNW52ge1OZGCvrimN2QygpO8B2Hss+KmSmbt3oGRnlN2KjbAetA/5Fg9NQMfhpJt
CfS+M8rqZGEZqvLZhMGFs6rZSjjveN2MsGbnFJEiMW4zT/ZD2y2pdIoL2QHwNkNP5TvdsQey53KQ
WlTNKDcuoL4cr/vkjc1tZwOss8fCcqn2S/3KwhKxy+5bKts87kvyQ+wQC+HuxhSEfixhPgxUqguQ
QNKR0rdc/KvelIiqXXShHIKJdrfpPGLB7d1xglsju/jiMXKmXTlw2bF5wVoa+DXN66J/qey9g2JH
QsjrBKrzA9KAY1yKvYscuxQb1AzlFUV72k9CDVXKm/yy3WrwqyH84bGSdNKfoSUNyuyqHUUt4VL0
VdTRI7iykPG0sKMq3Vi7rbPUFTkEX5+7WxOuBLP/RnVDlq/amiEHDZgdIbn40GlN9ROf87M7KYBy
iDtwkc1zneKol4PDX7wwSxIr9/XzG/Cj3PcqNGQLJapmZBSJ9aCQzd+SUpYwDfWS6VjEUIjq/chM
9j9l4LAIDkGMJVa9CexrH5M1nXLjJ0rLB+OdBAema/BUI2IJMeZ5ksqfnoTxTwTPBKkJF+qJuYQB
mO71kYBBfPQnQbMvXu6Cj6eHS5hx7/nJCJ2J4Gmgd/bQTyu38KvbJZdlChUwVZVGJL9JghbS57Pr
qBjvOfNT+Mk3YsfCRj9FuQsIwYIdPfDWs8t/S8oyTKugVKdfQOBFi1wo4MOK8LAsFS2+7gBAEejt
1D9ZkEavjA3wNFwmH6djPKvEyOllJpXjFCXs+2m2//Y6p71LXlrWtKl3khu1cPPZJsO5ZVW7rIi4
7AJAq5CV4Hc7exhhIHMOPxBqi5cUoTuqkM8sJMD2oxnpjqCA/JKjuq06xySnMeiInXRmZ6Z5vJ3B
JfAKXGQMW5rMdfIr9KoTdvWec1YdMC+19dzXTJuCsfAcmoJ++0dxt1tfXId6nt4EfxrpxkTXnCW0
jr2L08cUV/5PRavmcMr6toa3XuCU8mMviwSQDKAvJwKVEHjfYRGJen4rQsrjbiJgCvFZSBy/z4r7
Cnb69vDCjAdsmyGFeEYXluqJPPd8UP/lvpkH5q+57NVIuFMI1P9u/lcL7RkXtQxMItyuEn9j3xVg
Web1BPdAik0ENIK8nJxTuxfB2Wiw1vfcFaE+dPkOLGhm7I0ZllbLtlTIDnzu2EcCTaWSYIq0UT+D
BHbtrxBJ/P0qlGQalXpGkIxprYq1k16tXninG6NRdVRXadhWs5IDU3DBh1bwR1sOjkhA/+Yb/2UC
SZuHV8tj5ZyPmpQ66XXw17HlAnl/TDs8WrvlyKT16RVTxNc/GiRJ975syEjb4Y4v8emN3eJNlzHF
xKNwRTGmd5inz36M7+/0IzVGNYiisl8bViKOZNfzs0xdKFNrZfft7R2O6U7j5gJW/E9ICmWXuou1
n1E9MBnAayZ9lecctDlzNRZLBN4uLh8Ic6Z9MVZWOQuN9Za8cTg8xVcPT4KHrmj2vL5VkW0ptWKH
ynZdbvxVk6WErVcU/QkeFrfX2qHU0Ak6UZ10SVWF+gBFia9bKplwhqlCXzjqPLg5C3EGTXV0PZiu
Gyv7KXqTGkxNZaqltbOlIR0GHPEtocfOImI0CngkwITWZ08//F1nMF2l/ZWTxEPPiM4ygISKHiuZ
QFGWrpbWxbO7Em7XkKNWq94tMttpMt1VV4Jy7lwqtg6AmT7G4LDTryIU1sET5RHmxRwRW120jf4/
U4c/FduSH0asF7xvw3CAlk39393MAdqHCd6nONEd0P3GQKrxRF5d/nrgbUrlviRz1czpEo+wUEK5
D+ikW6kKbkOGt+xikcT7J2YsmV+zpNix0V0vzcfu/RHsy0olCSwWtU/VEZ6jcuHjhW2+3yFd3lhK
xeN7qosNAc18zJtJ23vrQOOJjlHgkYEkI7sKIO8WXAf7E4N6pnWKrPGBNlgCO9vLV/Bpu3bCAouO
Dx/0071eklalIPKiLvz+UeFqUL4wZK4lCNrrGMmG0OwzHdKmDRNMdKNE9wZaBEENekjFVYo5MagI
m5LbDTVgEWCWYNNshCa3Kgi4ZfWvlkI5FZMYxwuiyJWBXWJaAHQ2LdtAuO0SmN6KVerXlfiL6kFK
SLSsqQ0/n10/hpcuy/4ee2eGIPYsrxC9kG7exVK1J110Mvd96g+kTnQ7BIe4GTZV4TslT9M/9cOt
1+CbmeLXyAXgxvKk/S/BjJQQ2Xe/HFAud82SPpvoEk41vQPY03VEsMZmPVAZaqvW0oYf21bH4tJB
3TxsbLZL6FhLXnueJCOtuaNnwGlEBWZa8bzaoRYupc3mLvxqxJCdrizJU2pjWhIoAtwhvAfGOhPM
zUWUtzlkC4OduqgTEUxSESuwOccgL95c/FjObnpQHDe/MFSvMqResA+PHFGGdSdDQnm9rqQoy024
zomLgwI5StokNC8dx2RZPO0szqYAWYsJSLMRUmUSrv6b2LnUvWcDHZN5k3E2OzbgQLNmnUmJuuPn
+XuWBEuxyKhqFZIlC8n0IxTj6VZucOrWPN0jzbwADG+8lJlOXIEUYRBlTz7C/tGY4R9mjXkTQ33T
AjH+g/ub5Iboltmype4E1FeB3++tCYwE2qdYznQsiDKUjK/8p09mujqoHM4BMLyQcGPn2VJTTCgb
cNHBivHsklrURJol/uZrrnfuWsMh6jnaF4rLn731hxGlvJV8lW5ZhktAFUZR4jfoXLxV9mBJuLHl
1aAiFUFmM62b0hIvy0kgKewtl+LA4yxWMacyu5VTIN2upi8YR/t27087DI2yAJkMPj6nb8zGana8
7ZE0PzHKtTOOc1Y/aE/bgI4yHTtMIplVXBxn3mbe60X2VzSmsfrFPXXoXuHHXQAj+b0aE2M7PTKv
e/+zA7OY5XB42z85gpvrejRW609KGl2dy7qf6dYW1/dBXg4LlpbvAUg96E+cjaevPob2TMYdhJSn
FpSW6anF2l1TYn78iN10Nqy50z+yxSo45CdNHPhmOJJPB90T26W9Hll1TdFhKg8OZBMt5zJs88HW
k/5ywAJIgKw9wcrY4ZH5LzxV3ZE1BCMUCqFLsOPdncSQbl7/j73Igj9XI0LIPpzbwApbz8BdHDJ6
7fMLP8HhMAZ0jQ2ncHhIMPIYPM4Dmtbi50JsNw2KzZpRIAdtXwwlwBtNtEiJ+tTorTtEcH4Bi1ug
0vMYTtpXyoEe5p+CRF60KQ71qmMXiNl1uIGcCuNk7M+CxSCHzvbt9Hs0bAqdE+G4yeVXrB35OfhF
hv/h1NCgz7NhUhOvNU+1PpqA+wjoHNCtRiU7dRqP0+LSzXceZaN1pExW5HJOWIDjlQBT6x5IS8dG
FcPfAbK+Q10IYNzJYVpt2fFohbjIOENIZMOfzlpDR2M+HtZH/yNgcv95sS99u+UXmOrF3WXSWS0x
4S19aF8mWCXlyIjs8YHwShu582vUP0GyUZCUm8IvhZiFtbtNtC9R0CeKjdfQ65svI9CU/4lUbB/K
fQ+jbSI1mhEYByByhChKGc1DgEIfbAwjiVsIzMSfm5F43pciwgEwhywjqPvZBohdF8V1wr6ntQp1
8LTmaj0HS567sQv7N8gv25dTGa0Axg7VNO0HdM2JRRDnNnTvIJ3DIiHP74uLZPlhVeVURwnWynBU
v5c5rCthS6QVw22EdADaSQBwy1pTM+pN/Uyg+6fWQZObfYqbU/ps0l9YQMfseXLguNQG+hejHaru
wavCimJ+xYFYsgb5L8jH0hHMLFLHpKphkNKYqHU9vq8Z8ip6BH2yTZmm6rAtESyDCr+Be2lXnmPb
13NBmdD/fOMLXxbjHjVf4SOVjadeA2HO073W3Yp97JnXvtzku9+VIAkfHOHaq/l1CfzexYNUclYS
o2RLRXfyOy58iFQ8dhz7XLZFc3gv/sHZMXNTNSsrW9vKsFjbPLZpEXaqU6FRZuvB4mDLG7J7OK73
GAulqtBWSk3ppm9msOtIoIuZCEjW7PXPhARWE/G4HpQdrK2K+VJAnHHrZga74JKEu/3mopHnglJa
wE9Wwsne9/1CEH1Z1bGDQO/nrTpXrJDHQi/4ov7HrT7CSK5XbnWBkVyJy9xhr4x/11TmiUzq8Fq1
nDjgzrCSY3tSRF2r2xLicx9TFG78KNGZTzOe6bE8SGFpviZ7UY5quSFjUIDL9bcEuLdrD/gwB3IC
Og5iRQj/NYhhNLwJMQtf5Ul+aYQIk0XKmWvbaQ3kAV1pwh2co4s2w+kJQAnMi6aa/0qmRUdPS0eo
e2pUt6NDX/k+M+TM5m8mnIu/QWlvGmuKvhhAF4FA9d/i/N5TjDmfJaKzcoIpkxaIAEpp+uF2Rtmp
3amw8EHjgADmISId43YsO+hhfjMJ6VO5d6zo0vfGUkhoCYdOR+1WuCWzxFztzTpm5C7wzSn7QvpE
PiJBdlnTfA4TWkovF4f4z7mcKIlkNm9rFT+/BoO4ZYgOTMHIl5BeTggDaYgVn4MIJbJfEDSWcyr6
IizWXXIpiZh6Qr+kDG3W0uXVvueLbvvej9Jn2g+S4LSIA1m+rS+vwSNygo9996iYkFdQvrCGTSyT
WsqjB9vBrZqBjCLMsYN5gw0NU2WoQtrRowR/j04AeeD6iDhqmg+rAVJFCF03bvyM9yNjmvhBQDHm
RmA0ZzMhSXSPmL8gULcUYZYQKidmtgHHqCpCLBJ5RdpIKXRWpBHwCWL6sktMIyTQeKYGSQWDWt++
z5RO6eR6fcYY6Er0QbbK5IFD4UrPwZI0WE1f3e/JnCXt/C0WtaiQ6GjRGLqaDnRfK3VCI38hOG+5
RlJBr9L+eamAlTlDgSoJefGysXh/dt+0UJd+OoGAiCPBMx+N4h5jxRVvlRHtp5ZxJIeWvkyVD6pY
yh+u0cSHvLhcF7J5OGKuuKNTXvoJaT7vYS1KmzgkHR072e+0howrk/S2WkiGOEJZCsFnrHrYZBBD
h5HQr3d6jcI+oI4gDdK5tk0mj7pdrKAJtyUlvKBc29lAXG0SBu14i73vHQ52S8LhQTLfhu8iEeUU
nmoz4DuP13Jcc8hdAm/yE9RIT2TxlxoqTwYDJI5h3d5ipBbVHTysmvN8+XKbEMG28piOnNrX64NK
09OIxV5911c7sdcEISgTda49gL4b6AFWxKyeUpFbHcSKzt7P8QNC1uxONZrbmGdoZxyOtpXrxBH6
YBlXKsYPhJIsALqGNdtML4B8P01SVEHPSu00gaa9FAZUBWjGkSQBRt/K6OMZAIai5HuR56NNL5HJ
SAmN60UkPMpYUhCoIWVqiVIN7yoA6hID5NaFQNbWGBjz++39w5FGXF5qJZlbrVSsvhvO5hK6Wz6r
fQnLYIvIbxQMb1mrzzNiNMT5jdXHTzbs7fsmJqq5LJ9ORERx3PhAjX3bkbYYqLBAYvLpmlKJbVj2
8s4kGFrxB9+C7DVs6oA7xhljgEJ1dtI1MUjlpIJMr4dUTAhdLJlRvw91mb5Arm3veiZGLLM5Eq41
R+Zdz8D8v3WNtD74aqmhJw2pL2GF5Vbb03w6W22ePT2bESrRL07HP2wJusiDimZHT+E5A1cQAmP+
Fd/uadQ9u+eLhMlcjz/uf7gubWJznw83KVmpRhcjiCECr/I0OLF98Q1jP++VO7q/gNqSjZmNwXo7
6uQ7My8+pZzA6ewQWLG4zqFziAYAebyH64jblju0v2I+C/JpI2F1lRw3hF+6J3PDdLdmmX7W0BX3
kH17jYYwB2k0J2oIbZGgkcFFVInzs51mwVXtrYoB5A9zOtj5fSZMKE4lbGmag0LtRridGupSA3Nz
epD3XzQiiXU8wNtA1yYUjF5imnNorfPjKgYw9L3sozyUQRw8/Ls31mTItRkQR04Bx5TnuAooSbzu
52OKCfjP/plPqU7CGiZQx9GPPUmQQnjqwHhsmSyyucOvCIZwkvGybb3SRs25GFZOOKPgUTqVcFn2
Fz+uv5utXoFztUV6FNfj0D4o8HVuxGOwYWfhC/W9U6Y0mb0NbwIpTVpJ9xLwXlzImai8yoAHgobp
snUNUa59PUDDOlEI/ZVTz+ET3aTsA5bO8MSuZ7LBP3LD1HAmbBqgRt8JohwzWb3QsaEeIMYdu2Tm
ua3ivfPejsuv1RizIRciBi3WbMXrMOyTXcokTxTaDSFxbE1lgAWSL4m1TicieMtbYelqxV42djJk
U0C7NaqkBQJXih9McQMKXWx6DUhZ9CWft9Tv4BqknrYtYxLKxTIdiQe3OqV6OT08y1iWXBqKoOCH
Ia11t5Ulyyf3EKjk+CQ0FYJwHTqqgphwtFdvOFdpNXECICzjJGPoy3b9vqNgd/4SIi97aBkTe4b/
EQRHAMLipivLzWEclpYPgcN3DbBAfviQuG50ykn32tDmE2PwPiH0Jx/9wMWe7c1LRsVi4r1h+NQG
Js0CSaiphakWWm7vgSORbH9tZVBdIwsw4m+UtZ/FpGI2jMeHMpiKdzKEiY9SGvax16hV26z5O6GW
9NQhkkFnFPULOZNOVtvE80RTln8byld/PefC0oUR032Fd/xrUiUyGK8aS1HVjZ03A0bdVgsoPsjI
LvKotwI7ETQnfuhl69lHI466axddUWcprOhyXTkJm13HG6SPiMejCQZ+VXQH6cl84XOS7RvtsCbC
KD0NM+FyAvQFV9LBEt2gQuu31SAz+CLzIgGwtjBfxav8GrVpOaDCHruQfboz7N/SJZxFsxNea1PH
v4ntuWeMarJyrVvxcqnLEESqZBkoaLepUF7M1L47N5CSAMVjwFVaEBK2qoKteLb0ODFqz0/FPEuZ
0yIro3uXEZmgzmxEcVVzK2fYxifOgt4YeM1dAENlIdctJ0SIojeHiPrXIaX1wwBXgL36yH0YpDGJ
PsEJypTLJXzVOaMr7JHCqW4wd83U8YofqKFLM/w9pAhBUFaG2lEUXxmZ0yhnpCR28QBYjKQ/ijRO
6bfPIK7qCJHqWaECoz8pusXwZwm1xXS95FP9ppJfFdn9h6Yzms1b//7AELi9y0raH8IKhah/5Gfn
gwE1zfhdvwuRT7p2IEtQZaJhmomOXKQmrUnakIpVclP1hZFUYyYtKpx6qf8ljBlnSV7v7C5IzLSd
kdsM2AdK4kV5b5rGICoxIfURYoVNoiTcn3lUPPREAGXnu/PaMDu9LQ0gHAKhwhIvkPNBhQax8Oxp
nTdhAmHtPdOFzvV6b7Aw9SjfMEhrghS2jnGt5LvnA9q5EwkuZNgKNsklwrji6f1noK1wHt0cbRzJ
6yOKWF+Wkz67/zNcF/7JIw+/pDZ80GjFla+kT6yZpwu7C/dLfYSiyfob9I1BrhdxgM2fO9QT1f5z
wQa2kAyMC5iCUXlqJYLNPLKpBV7QOcwrVH/DVOSrMhP6tDaW8QWSTNE1XMJ+OnmRjaV2iGMFUFyD
V/p8pkTaRwC4Af3kFOgcUziiWOz0VYKGc6hqBfVax8iR1XVg2yLpMGZL4ye93aglNyobncoWGzyn
BMtrmg6TLNHiDUnEAQmTTD6PeUUwlf9+ogSuEdkwSMlIFBnqGGifWSXI4O0TDlh7X0CzoeRVlJG5
VRpXTUYCDE0p1Gdddkkqrg0BKkXgs7y80o50KinIVzPu+h5sDNnmGgGQPxH0hpqXclHxqjPrDnmf
1aUhM6NGEqVowHGiNYmYrBOXuQpmWPSN9HT6Zd+OQ3Y/59A9ILYRukfCi2LBIF8/2C7S+M+8PzcP
AYzIf1Jm1cBqjEnNBxT8YfU1Tq56W6EKvewGjIf6ATi23exKJOs+kYeOZtGSuSL612GWqb9ASrbm
fe3pk3SwMIucuuBEDjgUB6fyjErdKz9mKHbmVVgtDTvTG7Y+noVN2LwqppubxEY6/iZiyXH3HJ/C
x5BsPXKqyBMIQUgzCdJCAvoti3uwmdsD0GonemWCLrBji2LNQnk8iU3wKiLs+3c2kH+pvtxaPPkw
D3d6joQ8pRQokuLq+SGtbYLlNNxftPpQVzsPDx2m7O3icXjcWPjfXLe0Y9/nVudDu/XLZ9sgu8eL
j9sixo2BPy7lMQJ+b16iIavMgN5l9d/yVWrhFJk+rqxL7ZHu7IwOVTC4upe73oKV9mj5CBEAnHRC
yWd859o8kiyBxM7fK14c4WrC3yFU0ltAM9uvuiZ1YqyLsMOOnsTKTTmIh4fGDOls/qLK+fwhS56n
nU6RIZoRostYALYwQ+IP7Wp3dVZGzuCNkj5kWdKI1H4HVWUBZaMs11Hg6degsewanvENo7Bxca8g
FKvmgNqJeRM+rABTAlw/cRpSXN/bY0DrndcH1h101Za2ra2M3tQ651a+GXULb6qS62V/xKmqwxw/
+WQOcPOeZIXk34NKxzpYxbFETfWmTXK0m6P4SOfJyHoSkY88+TOyrD+5pVllI05/8Qo/GiCH5XMF
ThWG7qBgIbaF+IHO8/RvMquGR3kKw5O70mIVxyzhpvqfCsRltZTZKMTqBsP4NLQ2wTnTXTsRKNIf
9lIXSgltrr9nzx5ZCsQmoChFJSbJbeGklF3wltI0TnJn4F7rkgpNZbaO49D6MdY0Oo+dxlTI9HQA
ybo76ibIiZMsrBG5LO7u3lHmeCSVNbBjdVZu1896zK461Sa4XaNo8eX4iFmUB2SYOy0hf64w+6yH
RjqtrAvbMtoJ+LbqF7MfFyVq/ArzIF5QdmEwf+kXOcG+aU1nY/fDs4Y0Ajf9TdDzIL80QTpiyyA3
30Cpn59YOpXixCOga1DP2EBBD8/96NTHw/X57A3+QoCJQMnim4pmYtm5LzO0bQn0AdyLwngv5p+R
Yxlcv3ovYQZ3Q16k/RuY7iV/CI0XzTlUjEWnqonRILTACEEBr4jUcr9/VIaevML11iE//0rI0R/P
HSOU1B59PFP6incIl4x7b9F+C5bBJxVTeD4xfYN23KnMvqdltHMiR/BiMx3I8Exgh/jpSBA0LptB
RWXt+BCNBAIY+AwyhtIRtU+wKab6BBWpqQ6Adp8371msqlACNg8m8Wf9N3UU1EQxLTULMh6VwbkU
1lrK1P2XBvxxn4rsJ0lxkE5VYYGSzVmJkQf9qBMsMPM/yFL9quPwq8mrj6lR8YnmHdilJ4i57L3y
W2c1EIkWGaLixdDapOwl/TauuxUOEQIlMUTfULQPQ/QBPmon6t4YgDGX/6BalOPAZcbt6TcpzovR
JatPtTZv0cLErhKQBxGamurL82CNDLiXc6IIlgCFDA2gkvctreex5cywIOqCK0wqG8nzw3BtQezh
ENh6AuaIl/e2OJ8DIdsYgYoFCgeLUXGnidSsf/npqRaKU3+G5RCku360I44qS9Jvv7q61mwTcY4D
mvFibiZRebkrS9hBNvTJMYCfHAnQysVacZzSKBQyrUqWGgLIxQ/lI8lefNAgOz0zdUwN+MwiOiid
mnX4jW3OvO2K4WlyJoBF0vTUSHCK3fWygXCp1BXBUfmdHrZZIyw+xu5A1ASPr/cMDB/tMsH37zvg
VmaS8HtNdMKE2aMdlWnz7FDZG8l24H+9ubDVHxOUANz90LnbCGmFfBwQAw/pRENCfHu13ru47ybT
GNwvaqJaK3OIU06qoXx2nIebJrkUcotvUsKAydpuMaXBMrD88UctUuHEu3T/eUfKrENsxmiZkwKL
R5ThRHXC5SBYND8EZqmhYVx0zs2wxK8mV4Ch+3XQPm33DQN9IIKcDd9nn9Zu4S0YxsJGPJ3E0CE0
vllUVQgDMqyuZm/+u7avZr41nhaoTfrdvYKhOMyGXnVfBbennxlmQPEKNZlAX+bklOU0f3tCRfXe
HEdFVLjUCs/H9X/W4OFesNhSIRZTX4mM2EBhUK61wCOdOaJy6nKhRS8uN7SJLW8fEEzRAMlCbse5
ftWnIMjsw8hdcSV8QyfhkRW2kquwqMh0OM3ZgdTzWKwMtIVF1w1qJRxusckmAZAAPeX3Lp6TaQFG
tlvy1V/KtcQmzMAqnJL1goMkpTDCygPL7XLcuBC3wGsigLuU9oO/GzQ040W9AVbeRefGWp+naGt1
AWYpqXY39MmXvu5H3pVX1oygfHI+bMLe95zoAclYHTmeGFFhAZEb9V4d94x3V54gftaiBxRLHk/q
Kt7k2TuCd0aGfJaqTjZqbXXRGe+LiFyvrxsCM8/ZHuKQFiH1eWmd4H96+DhOHugffcG/mgLhItTR
coN2vWTax0hyr9ns2zwh/I3YTxNZZuHV6cMQubWiJNcoGOOJS0i/l1NT4syUHpe7KLZ0lkzIKnrY
39aUFM3sxuWoZriBdESB2LDpy51Wj1RoZA/W50ZzYpZKp5dr8vmJjQNiv+07FOWAQoa/Um07XoTp
hA4snk+fD/0FKIYmM65gnjFqlVClbMDUSHqC44tL537rFY9K6l0TOsRJudh5twDRcMZ2xK9fbxSV
v4XeiIXMQX/XHLRJSSYos869HuPcDAzc3xvwj7VwvQ6BwcHBCo/aYBR9113s7WNq6SDYmEBPSx4z
r4J9ja+F2Z7ckOPM8YClS5hSX70eLb+bV6uVeyldlZajDOhPWqMJQ3Z44aTOm117mne08sZ/iWb/
j6Y0A04US/1gtrHduVVB4vyw+fdAsam1gMBhkCQi7N/fPn6Jf0/OK8gExfQi2DVFotQEmdbH0j99
C1bb+QHvrWWRUP3INXhaHaDeT4Y7ahWrJm5/gfUFaTK2bCHWXh9UUCmFlnIjD6ZbXORSRQOaM86e
p6lXUj2TOATsqTjPn+bNYAusPyQ1qvTBm7ihENewAkmfsJWYKlDuljt2kNVw1Ke2k9/2eLE7ziYo
n/Vk5JREXNmXpcXjX3rDJnVcQuvZ1+eEQHsXZopNRpmACtS6/2CHivM5PAooPH0TTuozpitoyPP8
+r8cA6zTlkxNNBqx2Q7MLdv23/8K1DXPqsW3k5UVdh66DlqN8VeW9VPD/5hQl/wg3X8RMYbnJw43
wXIyfEyRUe10qU4CsqNCpQSOmylXwotU0or9c39SXuN5qWD+hvmljB6CwnrdGk0ksD170fqyOWAz
tXqiMWxY89opryq1h7Hq1IDbjPpq9Xj0NkKFj2bo/RzLELYcauVKhxpD+pMOzlrIIvax6UjUmEGZ
u5vN/mkjsIh2dEg4/pXlggujTREe8waD+/ZtlRirRMjJr5Lu3rVxkPyIWDF6E8WBtOez34S15jCn
iaQ79c4BLi4I9uC+0wPs4EneV8EEeWmKcvH6Da1fNOVeVcCTzjTHJS2wmREe78S01UB6e2+FRGUt
PJ62tqNuEdK5W6SoGSoCTqmsVNiTC4Dgs/p5kwALfX+RpIE/rsBETUX73Y1ny23dmAcILeCdfavj
CkqX/9W1eUjUC+/D6Z8uNBQeqSnrlyxkrNzWThjKlK9cRy0Hy/scbi2Pv8RM0VVAhnVreMszVoPR
ULv2ONnpv//xagRUGf1XA2IJJFCTfMxQC8rnn9xOffLIiRMVZBCR85mduPaLR2Lek++4s0w6QLBX
5uOqQY2Kt+AbM42QsLu0aJRB/RvhxtkNDs7SMtKscbaqdwyUEOWUkxzG7dWCJ4Gai6i4MYrpvJW4
54gBvm8cV7upXgLC5vFFMuIhuD1bcm7piLxFeIQza6VCekc0cBI8r1BIHrEsVmb3NawBfnz0Nzd9
7utuVXUdpKvnI9hT4jMBUTXLeppeIeSajmrn8BwPXmc8GKWmPuoKlYybK2I5KktJfNBn21o+iFdq
TfTA5IESiX8A8CjiCXI/vfXrqY3vctjknvWd5vF4O2UpaAKBKPt9tC7ZE0pZKoOig/d/+zedZoqU
tzGFTOerutBkESHrDHKHNDppJnbDsHhJQfK6fzhx7x5OrD4lMmHULK8v+lUenRMD5dKQDSawYh1i
zvi8qOSS9X1TQSsudsnx7U3PKqDY5AEMjatQS1v5fc9gIog/a2P3zVgUUzx9jaCFZyqhFYkN3he6
5eYuFteFnTTek09XqXk/EcWjsgH91UUJCNktXGG2n81Y5WMjLjVGN1aqRETD/IeaW574I9rFzjIk
aK1G0VemKF3PZu0BH8uyaae62+H+nVBmFXOh1oyKsyQHR+M+R23FwryzhH48ioSMm57P9FxSEOV2
9xPCGDg5jWCyIG4RiiHXnmJ2WnbM+X/UPey9YraVX+BXcs8Af6fn97490pLGiQh5XEmPO3BS9UoA
QL8IZpWw2ZP/VHrK5Tc4+BnpqAUctRooYtEeaspWY02rntn4BGDszBMpymNp90NjfuJR2/cAbXk+
pJLLLTjkYRs/+vapWDXVh1IjoKMDojfjDCFIyQjYVyS0+FzveuW+kRUrgld9ne4rTVtRU01p6sPT
UAzqIzIJqRrkFvcScSzQFvCuWX/6tD594Awr4vdfnNUzDs8v+ZiufLilpAND2OqmJMoIcIQQMlrH
o3J6wIKwCehnhVYcYC7I1E7ofjCHvEoZTglhdixIL52ZHzOS7mfFz9Zxt/uT23qvshHuABA4Q4uA
g4T7bNlrLjHOMpxw2AP95krpQaQ5VFe/lK2Im0rxGSwL75nGFFCuXxFlqAwGbWooy3F9uSuPy9Y5
lqRkRDmqKO0kA3j4rIp2eXxEqdsHRxk6RzVA0Ta/N+bqYNahMNfIQBLAV8J9M/A4JfzUmiLOvNPC
K4fOoMqU2L6s2O2fVdENsJ3OFXvHdQjB8pCdOzdW45TzHQYPH808DQjLOkBDK2Lwzc5N6PWh4fYh
7YV8NGA9lrQGdtFHxZ1ltSSigvo5D3ztyBxXuWyxRowMTquAXYZzNNNhjf17szrqsfpwHIbcSbh+
Q4sIGprCFrhk5I840OxJOVevmKpROLuwIJJGBu+0ixCpV2fUOxtiLGeoVbIOuiH26M22D+ZbaScE
Al4qATNhY/eeV6eJ3Ky8Quz7mjFbNVqVatX9WGVh2WoSSuLgWQXEDzjjeKEcN0EAGwB5q7Ohk5MW
aZFymBemozJAqTtwPZWMRBvTfIFu9MGV01bpYU7Z0KzT7zZIhUbASzjbR+4yJDKCb41uU2+TwwT+
u3aEyHTDdY0oK2f4kyAoAFWsR1UOommvmDyebziUJN7E9R4yf0lNcHu1ryahYKXhfzCfEg5OlS9J
69JPfnqis+hsxEYf5n7CQoZWxbbs55yGL2hC/TVgyKLCjHrtF5kaDnpG9+c7+dByfzRgF3yi5MV3
yWrxbyKIqEO3TSBQW6RTQ4S64YbwJD3XIeH0NFwIp25ylfsewK3M70pNFvTYxjo4p5Odwg40I2t7
CVvHyDGTuYIrmScPnDcmcCev72GrOyq1ufQyOVKwKqdp5JYinntmR2cXmafvKTAgUl7HXHJOBhAs
6d1rd24izDgK608XJt2M9350SxZQB14b8dUO6DqCTLCoeoIidqQ5aH6W9wWRlqa1hb7XIEFGNuz4
/zYKDESwS8GUujXuBcujM+o/x9dVLY+Js1ThimTa17epG/4rhkHSSY1jMY+kIu37uIgUv1DkRxfi
da1b8F9NG89szOLtbwozJ03qSEq9MejvN8jZTnU7PKdkq667hZYSLsz0ZCw9ejykDflYvGNgEVbt
LOARitCn9ZWQPhVqti4jzJZBVje4VDTH6IElAWgkB/LsnAZ4ydDkiDyFpuuKsv3FRAJAXFaKZKGv
wgQhkraKCJulGxL1RU/VgwEBO7WJO2B5EYxwNoaUmrzklhAm+AYzULCBtWoDSvu/Eyj1D+/c+tHk
sH/rLJG3KMiZ7txe+BFw1FyIYlNTYVp4eEe9Rrql+omZBfYI2hIXwPDFDUvOPaIRN/xT8h4Ycv8I
bp/mEZGNi/sra7pqgITZpILAWQj/w6kMHo+xQ7pnY1kcw9axApVhOMpogFdKl2x0C5+umkKuvp0j
2H1mNKOksD5MIWciH2BiNIWQE848vPaOP4+gDi7LxdnfavAp0B4XFk0i1hjM4FTnnCKZsrkDWlit
JLgmCgHJf+KK4OMgmHjFBkKSx1fbP7qolHqUGPRfTiYkFfTHmwjou6XpJIMzX3bXRUw6z8HBtvnW
iKJVhOpGq/naCYXHDz+zUgdECu0y5jBia9Jt4rxDmZxr9LR1AGh4Kg4Zn/6pnMfBKgmLDphLg8Mb
kdxS/WRg3eBvbUCiZxwnu+Eh4Q15MldnAG/0+5cxGLQiDnpONTQuDS++Mt49hlZ0G29SFwIQPJOC
OOXTsOzjGZ0RUI6kNZrkvhyQ1WfkEZW+pDImajKA6xGjsQk5kU/ZFibjSB5J1U8kz2nvkW2TNIXh
js6dAfD0RsTNTfoLpC4VzjdExQNCSOQaqxYW5JBLRXastT2Qy6bZ4Ti3UnIi3AtyIRjBooE/xbFY
JhevahqkuhVjDmnS7+PaObPtszRulyZulrdIw2i1UpiOgne6hjrbuQ2U8459tVCuOMxiSBqSavgZ
6YJtuUvbwJuUy+6MBQ7yzq48PVhr+p+dAKmY5CiKNA1owsrk6WaYeT3xSM4UkqMv6iAMJfv4Ce84
BAhlM/O/JwKgHqX8LBO1TobFrrgu0/IDzssjydwxl7vXbT5NkvoH6WsTJZPB9CoucNRlUvQseRC/
oF/NSX7quAP4XXdS1l8pjCRrR7aPP6y5X3KP7MVzInqELiUqPU/zjZG4Dy15NcCSiqZTupEicM0s
T56iIhKxod58vzvaZAQ1QWad0ZjkHrwNlIBtcB2X5wVH1+nKtF0riXGYd/wexV9OB+mvqWzE0jmO
53kOeZ0MhpxeLo/xEAtuB/bEGQyQ5QJH6bD8gRga/Uctaytd+IcKSMl0klOThUHCBh1SGpzVmqwk
bABtcMkZ3+2jD84zjh7nX+xkpyUbqkrMpxJCknZR9yn2vU5We/GTVxFatTvWRhFN9k/m/B0BETsa
fdAtl9bVY28dSyS1GC/JDxFiQNLWGU0Z/W+AJZwPS35aahmYVRj6JBPm/ZC7CFtd+Arb0KNXDKk6
Zmp07jLyS4WrDCdnS39HfUdwEx8feCrXvhn+X2mkdm0eKrLyctiFaCC11t7TZQWhiivWIoEBlcnG
XJ0OhPUHNEy6vphjqfUQ1rtaJURrhsWeRXOtezoN6BwzVKUkuaZlCky864fXi1G7xihIQNGQ5IEL
fIZjGyLoEY2yH5uEcMVCmvtfCvyi7MjcJr1dTCZJPvsemOiFtXsCvFbPu/GW03uX/rpXPAGb6ui3
uYyTVn7vKlJ4tpPPfRHUzgPYOVKHYd/DdmBUbbJM+tmsHG22i+3Aq/vK67TVho/Jda/RvbL2izSC
ovaj+QKMwY0uZPNWhyEUEBM523YPNJKBJfL0pzTuSYLu36ZFCenGWD9ZggBBhTZu4KmpUeRuYUCe
8K0B5u7XiMrydVnaqDWJrXTJ0H2i5wBIZG5qNwow21CvROBkBFtuVVW6bcaCXm1Bs+KaACcmD++5
0ubnK0B8EFvqsg12vXg75C5fWxBgtgCsldGIhHFzjKFCBB5/FNLgewJa5Mb+ewy4bjbm3h5yf/ga
M6q+i42XTqLlChwBSQfncldHHhGgDMvVGp78zEAphBQdrEeqIdPrFsj37e/WkKcLFMChaSev1M98
6/6Xp9Yf8Flomi7KUOc0u86SJUzPypWYnFlTlsqhoTTxLZn+ucUOXybdJn6Nilnrh/aXsbZVQzCl
ICc43Ju1Pl+bVDdEAxSnZqKKoelBadTGsh/PVwQMTFwVtDfKbPR0fx6dmMC4a7/spZYiykiVXmna
JFE2wuYL2hl6IKwwDWs+jqsTjOa56cWPyiGDGDqFGiB2A1Nfyh1Zk4cx0ma/kYTsnvpqA3mhmHVe
r5Qs3RKbMBO+fG4Je6Mo6R3rCgqU6L6Vwp9g7ZPaFs030dkBt7XRU3muoV+UMrhjoxSwnt8M4QWK
SaJ8JYCsXrXloddtPENFBQKxV9qdyhJ65ISTbm/9tiJzHXtV0gQgn7WCw3msoOrT/JAXmU9Y9ZWn
6RbAmKyniZlGBaHzqSO48mZMNoDI1niLNbqZiqaDDvqxewK1SMgE/zUE0Stbguqj+XSo6exd2EtS
Znv1rDuiTdUxRm8+pIC50Lr5jHFU/NxsPx4idOOPyVZKIwGDllj1CdGv0iT0dm4feJUfOOtlbXVo
Oy4fLY6/A8tPThumWTuqiUJ5oH7uRbrbtQ/9dBm3ctTn99x14E77jJlfKULojX0kai+lW2LXm+MY
gEoZIcNwWvF9ByCwCLXguAvQolyuxr0gbtSoUs7klVOc3Ocr4bI+YOXtvDsjSCSj3nJTQhZ6EKOz
ZAacZNPW9es7IsLikU4+gRC3e6XOzFBOuMC6sd4UUMvQWyD/CrKsg5b/O+E2U9ncuYSf1NpHeXfw
FCdFJxi5QyPoYoFtB+0W9TaQUkEfI5TDN+WpeJTwQ6k+AAW+0q7DxIbO0m+RFbW2ZEg+k12YQXRU
KDQ8glaq2R6934Z856JtLT6VKom8ZnkKLqUew8WGr1HIXfL8RmPty4RMJPfFPiffDhgI8SC+mI2U
GUQsLdCg0mtK7AUNFNkcNxl3rdEcKoBBebj5GmZ82fHlqaafzVP4WkfkzIM2ysPRIb5ojbTHDjzf
dTi77a8SpkXeHnDA5rRekkZvwssIz7d2cOJu4LkexNYP6s/IPBUyjcjSeBZ9v/miwyheSPFPm67l
HI8HbWHDmohzuZem45z4hpNeKCr/tkupZKhr/yO4wFM93ioWHbS5HR20lidmWka40kvzFtxIVJpA
hmVT+PAAHMBDF8HQxAXM6eEdYfy3T5x+hlyWSquq+ZTv8xEc3A7dfPqO2nl+QZBm3N5gQ96nlCPK
1PZiC4w+hMW3lXSuGQj7GikuT3UgzSpRkcykmQiAkoPN5b+CcEST0fdf48FD3IcgptHapv5ckL56
iug4c1qJ7LaJU79zlLC22ij6ppor2+L6HDdIyVqIaJ6b5QysJ1wMij5+5sn9xNFD6wZhpdzbUMTA
GNqgNR+nMfZQjaRfhHSOCwQUYjnSRHqTFTUVweuJjnhYS1nzTUdnyoS3nVMcMGC6ikMlK5Ktl7Kk
PSn+HzaS9nwIeYUo/g1eO2d6dENJ5I4+ZDZPL28mi7hw2IeR2Nzxj83h0TDvQa1PzY0OjDC9ooGR
6Z2njy4wNaPGy9uFCTkV0eOc+VA4UrYuM1eXSidWrIlVpzEbriv/KQj7qd+VJ4a8NOmqX+yRKpkN
fQNPL7v9KVJ0NhTwxbbe/rGxshu3vBCUKAI8i89E5NKsYRdSDVMwG0E2F5ZgnQ9UM0gdUpSXijCL
FSkowoJo+PbTvO5DXR5AXmqIAOr9oJv4tlwbAr0oc/tTf6tpgoo2OekcWYEcDAj2jx+3cjn/+4Ql
IKyf0hsOiNku0NQ/Z6wl4ezmCRfO/267VV61GadywDhRi84O9Im741D7WppEdedPwzMhi9v96WqR
L3GULidLcDiBya8guNmAnYkf95QLz7GHT5ikBAdh3e4HAb4+FWDhskyU0w9CL4hy32caVHjEj51I
aCNj8JJYeLHz3ypxtJQdlyyvpMDO/AfBQBqxsuYHOam1lx/9QS2RBCPhBx0AbJ52JvnoP+3sYokK
sH/z4EWV3nqnjH9t9Z4NtnbIaQGcNkMuTDxUzIAQc8dtUU6r1i4JwoR19pHXZZFuH4RZDjVX2I/x
CX6SxenWYxaDGZif097MfPbwkhUS0Qz6W8bkuKbbjjhOJbbsJWkmXEXK718GVPSm4e8XT2Po+hk5
IWR6Nh6ZdgoFUi6d74cSzG3zid5AQ1a7el05w7tE83rJHqmClGGohbbmIZIafXrOssNTkv5LtsH0
MvSZtginLtaHhtFiZ5ad+YRf7Ed5skUjrguHtyQxAZx/9W16ldxhyK3Wj3pWloBj2dyZOv6a5dK3
bSuu74zDRawhOpFB6qe3ObIDtFyrm661nKcUfi/egKdhW2OOxpUzuY/osB0abjUWEsbpfWcYUSkJ
eTn1krXKZ1puI2ZsJs7mfzMpupwKoVoVH99QJ85sjKjEA0vRixvVz0Dy8/P/gOTJoIOPO2GU3tO3
tteSjnao+YnrXcAy32FaInDJePhdTB1XW2yuwaumFp+5tYbrUGWHjEmHZVyt4eZTzWelWMZl7iGy
D8G/nethOxBb1QMa2HEF4dz8823G+hQrDL1IgnXJMfB6ibGncYWwkBvqfXfZ+mBfqYrpehf9Gtxz
tTgdQ0Jnr0nr0IFCovH4D59E35YdmT0aapbkFzxCCE1xgtSbmt+S1tXIv1JjsOY7zVEaIOhv/iJf
hLZ5BEtPjgFiCSLyrXdlRKbpNJAykSjis9lM9JkQZalvpt2YyQpP8k/VdFyg1BfOTjmGXOknczN+
cqtdaPhPE7tpnORFJdu6qH4/I7pXL5dZWPTelW8LxQDGWDQBrZAQHiWw11hokUj2NlqvtwFzHyqD
wULDoOgZPXpmFN0gn41QNByzkdv8EEXKSG76LFrXMimKAsTkvyp0Zo9lDIiYpX3BT/jUjLJxpN03
rwQvB+jx9R+sVibApJtVQqO4N323RPU1Ct7Xk+TYgFTmWksW+XYEsj5zCwX5ok4nB9wTKdxujE3B
BgRdAZTy1W2VOjoKDkiUfA8W4DQ+uFARFL0FG4sBSh+0JpcW4K+6mdsp3Dzfqa7lHzXshEEwb571
kA6PXHDX+bmNR4iSA5epyk0zdx5Aqk8GoSxI09MgKUM/EnpwkWhBcR32j6ukSy+ysNgq/fZyWMpr
5cTgQUg1UTS99CSIyNaJQfF+ZlrHkc2Hxvj+5Elg4YNtNYPPTcuzSAmvI4BbS9ySMGKQoCUwqGCL
3PGRmXRxd19nHHujBAgYWfWOczy4IoaSP/oSiQOBI7qEXAC8S4iMXpCw77ME/rQgZR3VrzpFLFEP
5V0g62F03P3Ts/ruVHAP0duJTcw10KTdd/aZRbyYUagq77pRro7MDNw5lUh4U9H+Et5yvUrkv28f
pUL9hDVLnS93eFL0IhaniiaG6J4u3wDZoWC8X/Q38c66orFib/F4ZvS0SBzIZd97ilULukrC4Zpy
X15+UBWs/9yif6EA7/gTNkXeh7frKVuux5iAXRyEvlZ1wyeIhN3HoVv/YAX7sIdgF5YrPrmQ7Pzm
0Z/FkoAmjCP2tcrQ7/j7CmPAHYdF1QNNEyginE00hzEW5KLEIjH7pVRZbaze3v1rT3sy6IjP0iM9
mdWBab8tulJDgZvej2OkV73SP3Sx+1S6mhonxP7kdIYHSUzF3I6EQjvVVDCK5J7SMMJ16M4au8k7
594+1oSAaHErH8R3ws/nY8LxQb/AQGRmvrcYoL2GuZ/HlI6rbELkMQDbRDWQOryijgAEUAgeXGZN
EsKE88SQghFsuRuozBZP8+whBxctsl7+fStatEBzKxO9J4rftdnK7GbXm2y9/HcP2OxrAJdui9MY
F8R9aZoBk0P8ktChWM1DQxlKMDG82kXJUIg5LCAVRoC+X5ulafwfS/OZRX79f7Z1IS1jfWJPPbTY
xixJiUmgUhXtkiQmSWGkh2kGf2CKJL8ZjL7TFjQcgkFAAII0ljMIecfHva7LKXbmEykT6h8+hsDB
i5Ix1atpQ3wrK/Sth3OhynCz0/t/zYGhm0hxlLtBFKW2FBf+W9TJmNeg0plAViowdtuJXogr3Lip
c/ApNnSxhmnaFdB40wtC4YQ/64NH9wRGF729iiCOV/C9B0d+rCPfasLUvg7iaXnOLE7qtFTid4sN
cgg9+2Edp+ehekJG9f3fDLFruyxncWanWtWhDSf3Q+xWOenyFl207Zv4unq/t9i9ersg/TNVdGYv
x6as94eJI60ESehVK1rA1+0x6KVQ5DItZzHbGFYugtjNhHE0heUCZksP0Sa9cAx+VEKN+hcS4PwU
3lSbzjQn7OVrEJNTBDTCMI9hGqfUiAxsF2lu8wl7aiUDduSCbxLTc5sETnkq82UKD7a7ppYTDf2f
4Jw/sp/4PqMd1rI0vdP2h3A5MFUXox3Bch7h88SCCdya824vggxsuACdrBvNgwtzBrjkbQSJ4WFh
VEf41jHhPiOzDSkGoYPlycyK6q/xgrqRf4MPEjA4cZzXPcZqwfOLmvmb6vsnvZW+ZTMA3jauUrW/
Onj/M8LM3yUZois3URDXgarhBsE7kaG8mneUVn0ULwUZbwSAeTm8h23KlRc9+H4Sbej86yONSIMp
EQgMjVvWYbeU6hKwscGlt0L43qB2EKS8iQi+to5aiPm0Y1gxXBv3JXC+Hp7Wu/5vM5rJEULq3HnP
8kG+ZRVpoUYzr9JkbOmBrI0oSK74wHptmO9Mmtn/6GpLTNQLIyUqoJonxwOAr0N8DzOo17ZDBZPn
W/rgr52ZMUqcTONyouqfNS+kwcDR1BBxK/Im29JaFahZRTL6JDzwm1V2x/5pBbHf3cMaIP2S3TuF
/8wJXlEO8XutsARj9BSOSXNt1q/y2eOsdhl+p7xsBIZeTVwZW77ulFNG/xX/zRr/NiVr4c3jHYAU
4EfBcnVcXsZfKDlsNaWQA++AMynryUffNe9xuEfKeD59ykbffjvk87Zn9DuS5QuxjreHWvRfXwHY
JDBoU73FPQy4lnXQR71zh6IPZU4TkmLe0yDW/2FDpFFd45dtKT0Y18fMsLdMatI/R+yMlERIcLl5
3Wks6nqKxcU0VD87DF8BvfjaA4BEBlJYP/2GUAc2Zh7+quwcQtsND6f/VX5WuDqBdi50zzvBJN8H
SImaABfxu2IQomcvINv+PvulZDoBkmepHs6BTTGvaDZ91utJdl4o9ycgoLVQQw2hU1BRfgcie64l
U+k38E1CFOKZwM8rNZ/nhuF0taJy/EKMhyq7MbAoPHGI6+Tc3gu4ztHsqRF5VZJmu+xQ/YjdzNvY
0Ruc0JhDKRcUyM2gm5fRlDGZ9KG2/Ggxz1LsOE+WZ7gkvdGwSWOXj034hark+UHnVfiIjRq3QTq7
M3ZuCZt3uFh/DI78gckkjXosF5Tve4azd0OBCykEME59GzhryxG6lvBHkCWhBLJl6Dnku2pxHkAO
MGsfVqJk9Zg+QajoxyXgVD7GltuRWGrnPI3aSPNAAolDrnfTITd5jOp6Hh+tj4e5HQOydksGWzg+
ijiMr/ZjVB1/3gVxIbxG0829tYNwzcVKGkeqC4YO2N8o5qvTiWmDv94slNzZkPyIEoR0qWLzDCTb
exOXAhC+9jR8dNCgjTzMOKLEsanYRvXRAO+klOl/s5b/ryTbVrKMS4XUU0WUbY54Eb74ZuA64/yO
dL95NbsIODp+yW1+yTLQigDyJPLaEYpB+5JfGZELGCXcAhn+x/VP2YCmk9UxLUkrXYGD2mjcYFwe
+QWBD4uSk4VON3mWOUchE0t/vrLMSjAhOHC65dva9+69bPskk9U3diaAxTBn5jqU0nmJBGiNmoM5
cohqP5WwlHF2g8fiG7KAh2D8F59/PlAqlzn00m4QATAfNulzDP+O41Lrr3KdK5OzTyTMK9cw8pDg
kHWkNtl33PiXeefhIOT6kA6ohDjps9di1oEHC36S3xordoEcdzuEFsUukz1EaD0KiSbCT07sOeuq
gnDyLOwYYU5v6D9ShMo4MhKV6EweBltRlqpD3D+VTHKwxV0v1fUeEvPNn5SFMzDD1im+4FbsbY0G
DXv0k9aXFD1kuP3R2JGMuRJItusLCO7wx2g75n9d2rvclsH/Tj3XiA7suKQ+5xs/gvCj1QRZrUmq
JJ4s8Qu2B1VxDptCzxbt5jqZ911Xy8IEGjXDahq9WsMEkRWh/Y+AfZ/DnZLfQBjsGb7/SBSgOPjk
SZI6mXwKGp0wlT3arbozkZzvqf1AviOQO9J3OGhT/NjhjOVC/3X+xt1SiyKDK/P/x7QVgFyO6PJq
HsxbZaTGkAI5u1axenkhSuWmz2MU/eVOwTz3fkyji9SAu1J47VeoqglycPTJdwwvbmrvRtbgEDqf
qLaPy06rgzdn/z9ImJhxRWrrU8Q+KkxtJniv/hwPkI5cOcEeMF2L/8Q0csj+yJQXr7cG1GLs/Aw6
ZM40iFHFj2iixq63pp2hm9SfoUAWujPRJvaENi/uCvlUAUdHaYZ6w5boo+bTOfSaMQrFLdl33ECb
pY7EOjTzWwCh8n877zqBvuFfKmpEcoARYMou6vGmDvuocB36oKxbvy8tFR2N5tB+QfF+dQVoge9b
m12EgxyzurVPFEia7HX+hRhnrCkoNqkhUjWuR91HJbvsLIJf87ATpGsNQzf+rNhmPDSUaNgCUYFt
B/uXIPsevw5Y87daM1ae7/r/sqPWamjAelfhA375tmeTBxSDQVJ9AWhouniZXBasoW5RPpbRtZDT
cnpfD7qui6VL+bBC04zMNJJdy9IBy3LymSnQEsQgM/RIBHmOYLD+TO1luDhRBgu/0hHE8GeHSCwt
ZSEdaW1gJ/qWKyO+4ND3cvTJxhiaFfrZjORdrtanqw0BU+3/TnmPeL/q+jmlwL8cQBPNUfyG/MYE
aReNr6yYokTLhGHS2uPAkabCjPDnlEEl+VnDRmCE4gm46jFK0lbMwnQfAkabNIm5zNZ9zYOyjPtF
ldC8SJC9I/7HYPDTcKPMF5Lr9NdhPd8S+oXzfSV8pM5nqznl8QUhzMH0WGS1erQwyDXY39ThPvNZ
birVhJktQAcKyrveqocvPBfQsp93M3s41fvalK1LkNGZRL6/4QhTFPN25bra4uhdlI/ZBkJCxCM0
JftygdOqVabFIexqYfwYqizYPOoMZwEyRJhxwxypWBsjkApbWz3qp5q/W+m4K7xL3ldllqZb9Oly
ABqgXPmXlven7yFMPKIHF9NChngpuN5cgZMLXFPIuWwSKqTQPiB0yAMEHYm0zqqVw6x7LIsPZJBP
ABcwZAXnfZ4wMg7HQXLUR8sIrLDNysJILzM60ECXPGUDp1+B1nM4gMPxw32DY+eKsGaOyOHvzScn
a8dakvHLBcvo0BGGlCq+CKZdgtcCAxFsTPPW6UBd7tLmGQyCylEDYeodHtWd10QXEGR5YqhAEZMB
HGdawT5JmfqVeRxq+bhHOt1rDp/kMXXyF2z4D5N3ouwobKX8VVTYQX5vMmSlvOvKa9rgCInX0TZy
U1gg0oOe1n0upsCvxUO4CL0/q5vl7a9Ejt4mI66aAaArGudlKaFRFOXJgU3sAHiYAs9uC/lj7wpu
/c31Ep9UtDrUA9WLis4bwU1pdyoJhKTSHZR5OdYFGDZtO9dT49Ib8niFr6AamHJq4jRqKWqYFRaz
dCkqNUdRAnZNmS7HOsEXLyd/8jM6HSCxYfnmAR4pYzuc7LClYiPfJOOJIXWHQm9zbrHYNygc+HT0
oW/DxHxFwQt/y8mvdy66IslLm73vMBv51vIRIeyaWkWpll0sMKuM+oUzzVMxJHgyFhWe8jo2dbd1
15yItyhgwaaQD6BHIYo7H7K/jaqxasYSbyt1+nD2snIEcc/RexEC7mTlezcQgeWYa/zFdwkiaoyx
l8bdcqeRkm0T5naiRVW41lUysiKqkBajZ9LYDJpCjxd9Grhb/QDfzX44A8hbdcPhVJUQImfPYMD5
n4/IrqyJknDTRMCLywNmJsYOrPwDbJCO3TZhctZdjTDGVKA2aOkAH8OsA48Dcm/3+JSero01nLBR
hV+wvyoFaKgWZdwx2jpWI9uWDgM0OaurFgDJt43wcOln5NhNONPiQHbIOvfwyU5oB7pu18fa/Txy
XZrJqsbrcIl+K1r6v8isHZkO+Y5BU4ofiCZbnvh+CJr9Fw+Y5ZlfxI7pokf75+fRZMW5grd7ZK0R
UJWcnCSJZGJ4Jnzxk7oFDh6Jp2cek+SA3eqiPJSFV5dz0xYTHi+atuDz3HFwDGJxlsN9UE+7PNXu
xJRWOgbechoeq1tqTdBWMdoVTwWGR4ZAAn88Om09XVR++EvQ9l2aNGNjst8038zCWnTnbShKI1sg
ybLMTry5V/vuyXhuEHCyGtgf7LAbSv6QIDO2ampmCoPyke5E0//1kxBneEnYITzaC1BVJYtq9nmU
y7k03v7IfAGde2A0auvkCI5qNTk+JBg7uPdUdBXKoPHW51iuHLVfuc4tb0m0cNLGr8psMelPjHOm
uTBJdk+iKzTzCMUFO63ebjBAqf+EV110NHHMT1Rx966UB/YG2a38wpGg3jul6MWC1sPgKpDUFdcP
gBuERbZxK9jYkY4+siaiIfh/v5pcqpZjWDPu1FWRR4+4xrDRlC2/9U2f2AL3Es5XxQ6gsM0avqSN
pSw2MkgZGoqt8OQ/V3PQyAc+2XkgOS2TR5Ang+kBZWQh2euuPacRTb0PhaAZgS5FaYxGElcKlSsU
tUo4s9wEX+l1v4WfdepZfIZYwDIsGTi+73qI47zFwLgie2IXhFyV66u33cGcpiIaxeZaAWbN5V6q
fYpqokrYnt94qbAj9vFzfbV4sTz+TC9cJRUVNgUa4vKquZBuTyibyAM2maTLLWtcBkCT7IPLhfN6
b6PbmU/aDSLjkB8cBDM2gsh/bKiKm33WyBL90xtvbMHShHJogFmhJHKdy0vrOpLWIv411MhU0AKU
LvG/TmE5MKnZcva3K3BQwHW9SFwuR1tcTmfJ0KQyFbpl6Mtt1V1DMEiYVaJeYf5bv0Wf06qHP3Ec
YYEczh8PG3Ah/PYhSLZDBIp62rPjrgNDzraWOf+ObcYCFreZdCPFLu2JE4c19AhfpDyn4D37/AK8
j23I1Yks1SoLxmONfuaHDkq48ObEk9aomRWYju+uvSXssz/+Y12TWrvcZXm8yHFZPBTOGDQx72kz
/Md+vVkFxmDjULGT+fDdqrJCbghfu78LSvuoKoOjrTq2CifKKhW/L002RDci7OL1vE43kgt28YWJ
9TdOpxlzNh/ywGohCpilyQ/nSNM4xKk9N+pbVOaKuphIk+W/EqvZFJeebKz6v4KD2PAcqUwgL9cO
dqGuZqpEEONQPJeL2aGqbmJWi374wexXPq9jJfp0RIEYKWoROfweThOirxWSwrO26BRZkHiOnt9z
mWVPS/DDSzgjTumehMEqUZl3LABbBR3+eUb4Ml9d9qpOPrfnmXZ96uW9Gmdq1HzAyZR4wI5Os24z
uryxMmRVkgoU7d3X51MfFvNxWcZNIhaZv2PLzEq/rFd6zMSVKiXO8ULrLngVGF+WYRYgBZ5G1eiw
5F2RlO1fNR5CP7MZlu6chpaTV0yI36z/S/c6KQ6uOgxQ9FWusLXGtEj5rjDNAzf3Lejc42yK0LHK
HU+FZ3mhf40xpHJUf1Cc/LbAaoHpJxRu3wEK5eWjLkF5fhw9eQAGFGPr9iM3SDhwHkY3EESRrAA9
KjdiUKzGdxpIdUUNNUSpje454LB9AWxXStkvJBloqTdZDSpjrex3GpfW++Kfi12lzKtPNgAlL11X
lh7A+5cEu1QpAS7yqI95cpY1GzAekBkD0XYR5cbz3U+/QACfjXUQRcUu1kFDuI/teRbrihpZEXVY
z6OiBJCeQYezGdruWwrELCMmFkbJ+/aeFSXiw1a/fTygVM/BF2lPGARsfN1B+tXgvHRIOq4ZvADk
Czd5uddTQYqeB01FLRPwUAkHT8pm14Sy122nPYzDGcQFltffThCGc0vLDnhYMtYfy+5RxTzF1Fj/
xRXkmZzBNkoEG1JveQbGV3Szosx7jHF9+iCBNMWmCAKneFd4TMz1Sd0NmVIDBbOrVhg/HPtRwGm6
W011ndbkQXvS+1gaKMURgEhPTVhP+Oyi7bnPyqnDgHkm5YQF5yeHDow+raTx5Pi9cJq1LYVffegb
qQCLBjyCr1a2wLRe4jf8Rh/Y4ZNV5UNechulEXV7rsnOXouiOER56HarKaeDAqxoJA7um3VkwcIx
3eRHpQaFQq5p44zcXvdHjDmS5ZNZPk0Ef8BofQawJ4ceGimJEwztsco9iYsszizo892R4Q+ut0Tv
tViMmbKPaXbGzcKOiPeYt86wFQvaNBBUXIOMdqic276pCqfcQs/PhZ0ykQaSQovKXE9qkmXApd4J
jgLf+vt9LcPksdju5wiXFhkhAog1MF7Aqsxix/Ub9vAlP+inTIRb9WQpjScjtAM1ITSHZZixKEF1
/HalmPLsXykYR/fps5D0wyAOb2MHANFDY3/D7q9ezPNGPPSnznOgXNXT2a7EQHJM/AgMb0SXN0iw
4x5qUn2DDoYLvpBxCYJCDAYUzN+qLws3l6BFjmq+06amkJNjizFvGINg6UC8+c3UoDPdJ47UNJew
oczif2C6k5EDnmcPlUtgaRqbpERXf9O+4VzQM4tfkMf4UrO79acl6G9Av0Fahmow+pwYKhzUD2/z
ZpBSwdz5s/BpDop5JN/aTZ0ASyjKrEZcZ6FNO7JSk3dLnYWIzHX+wjpZ0w534aqEAMHRJBmxOT8G
c7B97ksYwEImQR8iUPZbuo5e3Tnv+gf53+6yoPDoV4AZwyvBfNc/2wPdkm+G7wJvldt0RNh8Ker4
ocxpRjOgXnzJs3J8lJ6nDTQWzavnXhP6/gMkcyzKse5qPUprYdf/f2r4UwCvq4ugknymLppJ4/nt
xUl3ly9Mhsic8m+InPRBC9V7HoBh9dpVmMJ4rmnrcrvGmxfOnJKRboSAn2dNTvpGc/5sCNHydzp2
qlZxF770T0LGzPEbJdeTs/AhVNpGwGXkO7ZJswHEeAxzIkVqkUrDDsma/1MOah46y6YgljQBYPvE
ViRpFWXqnwqVuG3thMTa8vMYzgDf58rZiJDNIUoafvMc/2Rm/pNccw+K3XdiDBra9U4lMoedqZlE
LFUf6yNo2nH1aZu2brReuMPWLdJfEhhqe96e16pC5lPy8dHAeGLaNG+P50o6C/P2SdFSZCs4m7nZ
30akP+d6IIvzOdg/beJf+yS8dL5qr8gM8k9dgSNHAXIla72XxEWrzJ1dxqSnOZbbbgsrI5yl/B5V
98GqDRC+iiQNLLF7MKLEkvfe/GI7mZnqmEgaMp04+ShcncgQh+7SVajs1qGuUg5iaO51Mnnhg2Nb
jzDsxq3l68PIZlyzOGbK/xWv4+EoFmbR1sFQ3GhysgtiNjfxMF9yjqH2tgdDYaMo5IiAtEyCbth4
qxvw3bIaCPkqOudRD1rW2+HpanWpSK0l+dEtYgTbDLuHjyERg3aeSCdTJJfhBchvClPwzvNLCjEa
uziKGpnX9Fut74Tqeqrz5Qv0AYFDbaDwXSBXMKQFtzrD3KLv9ykMLk933bX8Nm3T45opQS50FYLG
Xpkl1WBBBMeccokomgiC8nyYb8EnSwed9yGYoPB+T0bVVRfDDIu++Kh1zoBD66gl8NkNZxDxRnSf
wQ3f35IPMZlLDgSNhhuweW0iSFgutdxwQljsMYKkEwtLhAiv5fPIyhnJ4aTtw1qh3g4YINmD7odx
JzwUq3m/pyz9qvc+WFKEb+jkDWnmP8VeyE+Rbdi14/6rHYuX5vchtjM0VEsJvuKT72rRaOJIityP
5IKk1Dvr2xumsHKftcbiRY1Dtk+EBpiBzSM8Fq/a0I+5i+SLCkj56fsA6lJf5bpml8cyg0rmVzGw
iVcuNgPSufKlIIFKBZrc3mZcig11Jd+rVw+jj5BG+6Ty73N2BmTR4oeOfJ+Mx32wBATyESvDi9FQ
pbs93CKcvLPlSaUIfKmeSf3tODAu98siUbMG0gtzBmtXMXsdL5PyxQXIwjU9c6P84LDWI5msr0EW
VWTKDKuIG+q2HP3GevUOqIDsitzYKlQ4PtaKVCM5GSd4eg77UCzgW0a+Swz17qSSedStz6QUALOI
/rCZTI3UAdebt6PGTHIAeDtAShLo9/P4MS9WkOaNZpaPGwjrO4hR+uqC1VAUsBcoqBCHxGeWI6As
A/1U9VjtrDXl3js8pdk+21dKUqGt7lQCWc38I6B1Q0jppVQKrayh0cJ5fllOY/oC8tQ4+6pjh3IA
XUSDAZKaqak5KQ1ihNmrNi8/tCm1WHa2bmuey12Mpis15xs53Vag8mNSkPU8NZGNHrAl6PQ0W2TU
X6Lc5v9aza1KcsfipQYtj+eRsC5T54Z7pLPu8wUFWUwO3lyfTDEJikMEZnkh+1saxZAJmXdpx4Vs
cB+sJnK22V/ibIG5fxSU7Ib4locKLlVrTwucsPwzmIj34bEmFgcekVedTDWBhyru9nt2lc+yhK52
/2NB4CRv4kkkS/KsDTc8pR186m/NhSkOUsvZnTTcXk0gK0MC1i5tvREPHeUknt/tjYLx8cjJD/l8
EqMzELKrJ0pIi06kvW6OnY0BxFJo3ugvHWOAH5axQxURqGd2hjqRJocTaafDz/6i6ibMYqXTMDiA
MUfiKX81sSrkLS2dET6WGTqY5+CC3iri/doNHkTTKcT1ytzLqKpFR+qfZeYkOn58DmI+1U+Ok2Sp
UVFNIx6ZDieldIF5ppOTSETP68Mk6v2YgBsCLD9NclgY6CPt9sdfbV8NYT0dcY2IGrVcRRGp1ZPr
OjShmGDVRYkQE+yiUw5QUKM8o2hA6A0NGJ0t2Y8wYHpsPxyFmhKI0ddJHfFHEf83ju21GUOCxW4g
Gy/NfVv67FbJfBzzmtwe7hKn3RPfEFEu75FPsiEx0Wi5WxyxZspu4J34AUMqXvn5LwAS7UUGkhV7
+6wDXyvTZz6roqA1BgBgpa6xzho+uVW/c0FpsWe7REt60FnEAsOuReZ7NSg6DLTAf0SxLtmPGvNx
rXTX/GXl2jL6P+mF1U6zfozL3sk9enD6SbIKj8G/AMOxcPGI3gTZPmxLQlpe9HVvMeHcID6/hiLi
BxmEtVPXfe83/0RIVoq6a4S+WetHdeGGNTYZ6zL27h+bm469rPhACdp0WXSBZOQ9zGxprxbvUfo/
ekQAglFKNeyYZhRieuIqjNYHQJi9S/5gNnKebPIywH8BhZZVVGz1jDv8LV7f1imwZ8we9lP/I8BH
3G8i+Gwbp86SAXgrammApgMob0yDfBfYw73uAEpLxqR5WxW4T5aBvqCqdkgr1Yt6ZnoXJL5NklAa
eGu+91ktdX5iYEWDQ89Fw2f+S9qPvTCk4GugOV+xGc80Pvi9Sr01tSal34x6mUiTUUY59C160QC9
FPEct1ytRU0Si9pqUN24IVnxl9otJi9bQbai32ZI0KD8gQMO10HqoCSmwc5kBZaSvkrPYCJID6+i
baHoou1kicYvmrIaJN37aUyXtd+BdLJiGQyUzcJ8t90PTb2thTz3lBJarWcN16OM+lLPmjqJY0Sh
f5ogUKdl5gDFav8l9ogw8otY2MlyXoyCmasASGRPIgnGEpORw3RUhwsALu+vMNt+WVdWt7Lurdry
owK+QhUFZp1XOxNfdK2KxDKulPl2WMZ5x2pu0Bf23/s5xRu9GPP5Y07xSR5eeQsmyp5KJ/VVPayt
xJg4yLuA1eMuh62VqR9fPuW+qAqkLbdx29sud5bB96fzsDpUfdMq7Cow3TuFynmebj6+5Zh9qGr3
YVCfjsbpHckXbsa+4BleJVCKIKBConfpB3vR6+v03vx3GmSVk9x5IVeYhIDob0hDzi3R3X2lkJH0
kGwLVu4NaLNkR093FKZpY9uN/LHFRvXq/R/tc/TDCG3IqsK7JBBBzZxmUctcpn57T3gXS42jqF0T
Nqh1QBZv3vbhgtXuOqpsKKThHjRhuMaUbzXo4+vD/DxCCnRaVFCL6U82LL2SapFQriBbCmhS7jUq
vwLGA1O94bhF4xrNvVMqu4g5ChLtjWojy1RA0dne2QqPBUciFGgMk6Dgl77JBUHt1pA0uHF0JwpC
zbIg/OiqnQOR53djI87LIV3wIqLTnQsCV0fA6rmzkIV/cualfQbdbjpFSiG4g4qvUvNZ0wQbUYu6
o/PkkFzPainy1uEwXGwLRS2qgGtS4gP0MxDeOmX1s3cvGMbKBjKNbHkda187YdVSuGmOBnAg7Rv/
K96Y23Xa6xSAQ7tS4a5RQ+i24I11GSA4Wnfc1N5MGZV6a0G0dinux7AwfVZsH6sY4NpMmzIXb3hh
SzdwJ124Fy6pggXe2r7gRFe5udiVU2YacOldGejZefXT/6m95U1m8trBP/RtKx/YC74QQXW3HkkN
lGiVpr8GX6BV5k0Me2EqKYq0pHGw0+iXpT4SXzrc67T0A+IT6ApfNNdqxc1ZPZv3wcCwJ8JojvT6
jSYFktgEnMAgaiLj1ljbJHdm9eWOxueg3vzPxsbW+LMPWdIYT0HwReoZz9/l8qM2Py4ynP4Au6GJ
O2aj/qbMIjy4252hewmPxOTDg4kitujzQhumne6C0FpgoNFP5r9Cvf2OyOD3iVpIBLOw+goLfKhr
Jpgi6uJ/+H3qK2TOHSCBNyKkAhR5/ShDXeXHDyqY38yb7JTlexuVc3Z+5mIpEkw6ZoM+EZ+67Efj
Ut4isY0M4HZcjY4Q8+s47xAi770pjoZypc5es9tS932dUHZRyKeDb1IlxWWuyqQ4S7ncr8sjuP+d
b+Peq/BeE7sNxMjBSYXJJfLezrWKMiRqwoMP1bmpb2th7KtPCZjiwHQQBHf08/llxZHhqBRyHOVO
/LOmqlQ4tUeldjB9ZRPKdE8HCSOtth2BmyaJrXWSgmVS2RBF4fsJa0mZrGGMp47wumDyNKQo7HmC
FLLgQIZHaaeDJu3i1LKlpeK2DQVC2dH54PJTeJf4a/j5eiQDkkaX0pMj+O0Na7WvTIhPplf9WYqB
TpDBTkB6yNP0zTnOQOsYjkOvQsOQIgyTEKVFP2dIvhu0blx2EXHSQFCDthCk8uD0IYv5JOCiM3Eb
iwOmcWFIGD93NiAf9zhjuvAaiF3M+i09TRChem8iCF0HPxTRivhfrkP5Pq/wdzjlSZWgZwXmi9MN
9TpqOVkFgt31b2O01mQZ7pgL693O1jCIbU5wK2mYG47Z1gxUvP/6hyV4RVSCAG+3A8w+odk1XASL
XEmTkgATrmubIjV5ifkQBQQPB1SojDEVM/Wvk9EO4VYhwBFT6lwglRIDXWpI1rM0Y7ho4oaCWKyY
hGNAOQNDlwXMI6zJbjlEFtjO3LeYD1zvNmj18LXUunfRPvQ8Tl3CLctf2tCxgss6IIYTrCbzPji8
3TitSPMtpvLrL8jfR4iBaPV+e4epvzjAf5Lod7n3s2wPxtgRjvSrZ0LGkk74UTbDrrJhII8BUvFM
Blmllb4pUG4vv4YQoqqLDJ7ZT0pusKls0Ohn/PrjW8SltboOC4KBbZn6VAt7BG+NKcXjZMcIEfZy
x/EfoLE87y3xfdVh25aoitaC7w/MlXJ0qBNSUBuElkrOH0EXdlj59TUq5DxJ9A7GtcLjq6KrwM8x
SORnlLjSXjWlS+CX6SpeWUtfD/fg4MG6DRfvrl++i8HUJKgMHfLnOn4YT0QxXv12cJ2tkC6tKRDp
0nJ84VbaQwKYQCcj9C0DNY1XUHDhBl8p/xuHFuyWlOQFMUyfG9NVJjltliobIObxqUj2cK6lKaH0
VYdsflE40JlIqPpoLV2geV4OUjZMyUDNkK+uUlMjqvPWVosctLXdPjYRuDQ2tXgxxLgSyrMaGG++
zDnSZhrpX9bGn15U+Epg5zLjlcdO3GNb56m/WreFiQJSrg59ddbSUzpCVRUMtF1wXnJV1YLwkb4m
LqhOb4qLjiRVhGWPC+oMry67H96/L33z1tSeGadtKP7G+xkdRMiGQHqcj+3kbx3ISAoSja7z8JfE
18Slq+QAX59YXCTgBrc2PYV8L3InN4xisbmJwaTJYNJ+ECE7kT+quxSa6mZTo2Uc0yV4QAK4A2JZ
6xp6m+Zf/+KQfq8IG0tFz60P7PPzhHxG4F1g0GmZsStgv9rexwmATwl5G+Mu72UhcFbm+xTewFf2
d7HkRtfX+t1/QqWwiFukKM5GNhTChWH4/wiaRDjCjJ1X9xHtpPmwH/MIdIag2sqDbRSu2xEpcort
AvUbW1c4KW1+4eF3JyWvKM8b91pEImnHhihS2sBb8kr62ChHnVSn4+zcXf/Rxo2XnhDf4gTXlhPH
KNvxMrEqStLGoVVVrG0IXUIm6Y/265cvIdoBw8jaBOS0hxZ4UhbB1mu80693j/znwcll6dDZqOUk
C1/VIolBsNRd+6jtqdxCDshmSmi3YGI0nSDUu1JTITo33DDw/o45oVYGAIJa5H2G3wIGVBmkg8Wy
bCprWiRuqvgGU4hg9AAFNUm8waVken0/NAL2jWhhhS8qrp8wd6ecuxC0FqV+OkDDomTG/6l6SX/M
gAwcLVRxHfmGVAIbMzB8SnL12pOX0cL4ZSqqGiUhtbHsGune+bv1pCz6Q7Xp2McWjvJmWhh+tFDb
FqcdPqK0Wj3LrhvgJa0wIrlPfes9/+4S/9Ki9ggjEqkXVU+VHPMOoRzFt+3NTKjPmCzIu0X9HvzE
v04KIIeLIjqQP8T7X/B/lxLqvuXjbc1xEP0ojJ8lJtZ6uY8kW2JF7D5ZoQXUC17yp0G8AzA3CUM3
mQCUIKFDUB2AlmmT4SPk0u2GmBdGU8UJBPDsh4zQngv/o8zK+/WFu4d1Yhtmz7Dd7nHxVetLwh16
40KIm2ID3oulnYtL8yi2lemwfmrqydO6wuX293AUUeTfIoo90vjzE0IkWv4KCOD+j9AqHoTozMlj
ry3FAyhEsOKbTpK4itWJ24TXYgEKV9wWCNHr++XRkMwdfXQSqW+SefHFjRWMxXd+kfoRnppEdyKV
qN9/QEc4P4X0ICZCaCZfwxKO2PGyJVIgnCMF+PutiL6UNznz/qTkUWi8JuI6I9kny5nvpBsx9vm+
yPsV8irT8EI1VGxHtZyJ22Q4mlkwVys4blggA80uplaqf2B9BaSTYbcgmj+wgKoMojqnntIlDQlj
UyEhcQrzeLsrhCEoIc5ru+OB24l3vMfuWWTZDbcOvefaskofSivC5GCFtyd3NBC6bicIjpEzQ6lm
LHrrlnRbPMPW5b4/LYX10u+ZTo5uh/DKXN6m9OsX4inxXapuJWjJK2E9AJxhUK+0HhAfMrFDhTKk
DzWSvS3fhWiupfmSUM+3vF6ljNVJ4MLVNyYHq9ntUDMAwPFV2cIM4UXV4HE5IY1Wk8LeNOTfF1Gz
rakYnjWg63e7YJ9tjcdK2kkibCEz0Zx1rgGLaZhdEusBjHFDn7eR/0nsApZI0LE66UrQWjLMaG9f
CCrZGREmsDtNjMH8DRmbnTvNP/0904qs9r75UKebYnOWp0uHfR5TnmAHZa4tyAbkK1Iw1JRSaKFy
4eQ2463HgnigpNuJpUCm79GMfDrepanexLbVHDtOcCf6Da4EF2CAxdDuEkpRMiMlPcETjaYfXhDV
idJioNUxDXhoVtxcXPFeOKXYF/9qBcFmOjA711ZXEc+tgMocSM6akDsWW+Pqz29feQydZWePc4OP
PIahemZEjQe1Bb65Q77Bu448cyOKLbeyOUkWEn5T6LMbg/AGnY8rfqiSSVyTcpnlEFIpyoP6gxgE
mU6NXLqdi4xf8UybuvL+f7ROecRkfMNV7OiVBidnvx4p2Rvu8JRGhEfNJvkKooYZaffjmtbimvk6
JSmNDJLFeSkLULTOH1Vb67hrjNRSEcBAzj9C3uSL5UQSPWf0KOPPBMRIubUHJCZW4TZcX7y/S4T1
fzHwvX5MlwlKM5mK0Gyb9N+5MMexkT1+9MR734b9ZztCkvH5koivBqNuJC7iZmIrtF9NWsZwSYD2
20QVmPCFBaoJn+nbULZD7xRU4e9qZFmeOXoYpHZ0BfHfp+rXk8cWq83ujzk82mkjp+rmBH9hJ4xI
rp1nfzUzKfKhOr8nm4acfpqfpZSwYJU1jywwQK2LLCAqiaVBsW+1bcSCGqjXD1rDntGVLxfcKFYK
gcXZKTNv4h90QRvB7zoOz9NdQnkObc/CeXUA3dtb/cwFWBGJ2mLtFzmjqe+Lz1Tx4fZHlHPWZLC4
ARwRN5hvZkiL8SuiGS/zO7oyt2pC5esh5abb1vyBnRBA0kyYbeCK0cFn8UQhkGTBZTvG/5uBc631
LSiGGRCKKZiI1pPDqlHI9jqDdWPxBe5ecL5wCSJCvxhAxQuTpnD81bWtpXaaI1mFQa9VO+BuhnT+
KRtPhw7b+ZHKAFeZkr4AHCIFufHZFw/pSyifUsab1TRQnuV9A3xWtio2Ka9GF+AK7uJ21kOx5JKX
8i8zlOwtTScgO18RnGNJ85T8Tif+Kf/JezV9S4gJS3Eu7XUJfA3wZhkNBYMVopzNZKcn9ck9UV6S
tfXYotayZbiQKUUYQ2ymUIuQ18vc8eQS3FMRbf1QvK0BVvKztXmE+quaLsi7F14CHpqGnF8BUeCs
0WRLXudqEEKWCgNsFe10HPKxMSW5fGgD6N9F8Gl0Qc5eyYsXk+b31c30hhh52X9+sRZBvko6CGfQ
+R8vnkg8trc5dqIhLbXlMnWapHXR9aGrGQtybT2TA2rgxc4O1noR7naT3KiSGeaTLE0KJw/auE+v
m9R3/MH/mR2JhCOzkAPLSq7M/Vjo/cQ2xbPlgWzxSxsJpQc26hjJLOr20GqfQ3r3THi1DH03O8vD
EiNMdz/YRWwvOHaeQYdxlDN61e6l2l5HqDPi0TExvbCIBc8gwcfxHnTBoX5TRe5xdpMoF1BGAj2o
gTHJFojz+jls4oC1Qcv4NBOotscQdULJTvhqv+Sdannoq1WQgCVx8/Yz0K9j22qdO5rVxA8nRvqP
0ri9SxmVwMvpPYZDv9iDrYILrRlaLgRdFppmt1mbdG7bl+AyU3l58am9tVWnwuWglRbVoYyzM7F8
4XnTdMqmxgQGVGFmejk1R1ituWweVdbEMIfUxVtFi76XR1aCZALvQXO0qjxhXYV3ozBuQb7Z1wnS
6Bac90+nA9S063S3yrmuCzDG9oUSa01lJYwzziyanffxPhaMSel9cIPjFHTwykSALq0KTsJGNfVL
StsaND8NnCYOWsd0P2q/tfTbEbKanrYW/3si4EHn6Wbr7LYpWBHstWFq1Y3Q71KQnqHwUCtvi4aI
H8sOz0D+EOmBp5egKpCBTyMTNTH0ohmFquLmFQngmtLbeyr/vY6t8IBobtNKnd/+2yvfUnhWfY4x
iEYbz4TRVK/AQyS26ra7UMleoioRyJbaZJoQsT+eWzZNBKJOeePmRYXumFR6pBri/IkS6BqaOdhr
oVAaQQKBS5/AdP4Ex+5enqxwPKZsTW/snUkIU5qgvVVG/yNUBu8txEFfpadSJhfJbYET3ZmnHwQI
/mOgGUi5iJZZda6J4YYc+krQvoCCYJjT0YcWuXovrqqKrADG38WF9ALvE3KokSuxmqkmIGcBU4ZW
lPtS9FQGGfymWBITmWPaj8c/j2o9AEwKBdjhdGs88Bqw1ai1UER7EUN6ClCPeHYGsaXxedzT7Q6G
hhROv5s7a7yUZga1N7BeS8rMQoTqn3Q38/gs8U3jYG6w6GSoftIanAVd277GGdfAgjf2C5rsBbsv
P/qt+Ee28JBH0gCgwBzcr8pQgrI5n0xy0qCTfBCWG5R1LPgWnTj9oPaoH/pCme02fpWGLW9ylYFH
Edqzkt5eMncXjgV6cwxdm3HInzano2IAQPz8TddNBC8tQcGcjzHfTmf0wbKZQSLUbCrljXPp8Pfd
gdnnhSNTaRN/H4aNfTFphgW4XCTDjd5d4i87T+R/H2YFoSrgrlks0JfHria/A2rPuGqh9FYzJJqS
3vTQSNkGkJSZxRCgUO+EkBYJxFFcZh6QSPcejcBcXXkVRAGaOp4Kfni1qoTtrqcma01tIXF0zh3w
EBxDNwS4bAll3fYmFgPUqVu/Ai5z6Gf7JD4nOHOZStiyf7qwBrVgKrCJHCWCiVo/S12ITn64icPp
e0LKD5PHFuFz1xd/W59Hs6uUGR9PiRwwxuS1GMKUm9kOcQMcI1m8FDDlBvmu3Krmi+6r/TdQ4SFS
qSlnR6Dni7sVZOOzYd/h8WUKBUdGjCN1xFP2RsPN6Bygh16VW4Rn6/Tyt2TP4t1dnfgmHWS2E6Wo
nBcZa5UUzI7lQbbwqCNADUejRUqiw4l042L0sLhsaGdcV7cQlsEcL6LsDAio1y/vU2Lewa4Koiq7
PoFvWLA7yhULDP9TPMuXe4R/SbNDoB/zuLRqHDulroItcsPTOeK5ODq1dBVVidBxDvCwbrWpS/b8
ug/hsJ5/8741k0cqIsesI4nMy385HMS+63aUzmwM/KlvH8ayhEQSxMuanRD+Ob92mSatHDSu4m03
mvlIo0JlhGi+yo3AXYVwsG97gaKFGxV6Mi8onhi62toQ4iY//GOq4aryN7AciqaDUhTwf04Vg2hx
lTul5tFESMIJZaKagGUB/MIF0cjpIlEQXGrAjtDatRIFdN/12swBXFQPLjV1otDFrUvdfkeD+BjH
qKDPlhV8RJT/pbH4/xbtO04N+0rs1IIiakYMVWWf2dobsAJ7EJj6ULZK0Ke2TMR6PrXpi3WBDwVb
FZGEMV6u5T2WKLt2BbJu4Hl7G0GbgOlI+jg2t2Mli9PaBf8ZDqEvrMTdhannL4O5iLXE83hxlMZ/
B22GJGnvbVgR3f2+oQ08ZoFn9KC6WubxcGWIveHYfVGSYt1YA5ibo1KceCZAETvoDtoEETaaHNVx
jxfixNznaghbL6E9U5jWtz9/v3eKxps8YLi/CoyaYJxXaWiOkLfuupOqwZvguB66gYpEHaN6cFML
Ugtm9Os0Jlmy4Z+gP0Ei6r9BpyeEmmCOah7nxy8taak/xHW1IBLhI0KTwC7hxF8PWJETwI6h6CdU
ahZBlWCxgzFSo1WhHvFJ5g5u+sZA6x4dO5UowfLQE9tbgXaSw2U7I9iUlYAFWaQsiXA9aOSX0Uwx
PNwBeZs3voyX4RAW/c5zGFehf9Xs0T1EMIBQ3UDd7VFMw9OTv/V+qTUjUeTCc0CoYYpUW3jNK8JN
eT3nYU5WIK5kCsVM9gVO6lvKT4m/6EobnUtaKuzSVMk2ylcei9SUC193Cl/MNa4CbPlmkIGwDyhP
dKkRXT2z7hX7ttHsrHp2UHTWUxEbdP8cYN1GdhC9v7wLoF2L7Ry0gfE/nUu2NDn52vi926bMYCK9
UryXSj63URzomBntsV8iQNV9uCfIhoN7pr0sHWdE8uMnsVBywHCQW9Z+p882xLs4+08qdYEBc0yX
UKV8O177v+VYTAquHIxoj1lzKQT87TN6VpsMUY9Zf3Jj46e7BPVo83oMEnk7cv5zXjaUb08mecOU
5T32Epj6Y4rZXpturjetSbnuqSO2XYqeGyrFZwykCaQxSVWMKWmUliwBC5ljKCHQQm1+3o9eXypz
meMApXFwMlkLwD2UX5THOKIhFKO9+cByBUdF7REwkSldJ5qr8fkzH7UXfODWF4fVyKbUF2X7awm0
hjpVLD+0qzMlGCdz3QeNN2MKrk3Z3wOIDc1YbFCUf56icsoauHyAD3F1dzaPNInkZToUOruKeuHI
SDgnF5Z90ROmh5fTlm52dWjIMJOkC3ocVErY6phEfx9uvP1IshBldMRTH+rOm6C5UscPZOR9HSTe
cY78DKjdjXMQGFaCowlwPBYFE0mEFaM/G+NCC28d5NxvIHFlZxX/len8z1XXCokwPO3BQwfHl7v3
WZ3ORGc+XAAf8IltocPG2fRmAs9XgkNbtALPjct6IblBCXV9wy1Dp3J7jogHDzca6tJkDELzmnxT
DFFmwaQ8bSbJkMPu6R7ZmibAIujXG9sxiBE2I/Zob5Fuol2gj/BB21c2m2Sz9XmoOYKSHqvD5HyL
/OG1WomwnlWJLELFPwYywZbnGjsuKnYNCV8j6GcIkfpNXWPwZKQ4KrDmp6Hj9lT9FfiRcJ0pI00P
Axhq7ARihu+yYKXXUVk15m5KTEWhMqGaOWA0NTMcBbPwac/0ivPRaW/q/r/CrNQZ2jKE1QsthdzD
t5bD/kt4TKFzAAhdLikDvOnWezgCsClGJ5Y1RZJdHZrHqjrIAHSyxICD3tS4M4xP326EV/ObgD72
QJS1QFNRXfGBAUe/TMuQA6W8hwBp0P7WCMX91JihFf29WIFQ+HN6rShCKVgo3QA0otY6GJEhuhPk
2C5phMQP93ztGBw5mhs/o1vL25Y4YSdlA+k+P+oU2VJeI93YOi6gL/ufHEGwhm6VzyrLOrgpVvIT
+hfsuVxm1PPjBxQIv14BBAhCZks4/0xE2YqskGSR+8+9JeUk/1QtRXNmpcNNwc+jYgzrE5XR/otE
JupZ+aCaM7ilmc4s/WMNkOxpslEyCu5dB8p/lPCLZD4tE52xbK+oFDfeVlS1k4P6x5e1qD+i45bv
LwL4mf3FPtD/nZERZ2MAfKh1kRigydIYYhvr034Rf1WsmgKX3cpIIcTiNuZSYg00mFrVPFJZwXTo
ZLFFO7roOxLSc5WehdRBB5flOFugu1Gyf9ZJrDW7hx2TgtYAsEVxy6nSkAxihkh8WHluX0bKcRY0
a164qEVxPniMSTnMX2BKbtbb1KVfD9i2FmrkfIEqZTiol3LVUTCD+jOD1NpT0I9aAaANfYrkYluD
JLCDsTxgj8lwxvj0cym80PfVeGabdz3UzD6if5rM8lBikjxv1gVbgbCTVG4ItpLnhO4D6Pp7NlSp
E7lIUK8tOy2oneZbMcaK8xnUWXWbvOeScHhqflSysVyf6Vu1elCZ8CDnssKXkCqTwLxOetJar2y/
oU6+82ob1uN/wCyxsndp3a1T+Oywnj2x9j1H/uEHx5dbPBvSuvxpQZe+yftYrwc6K/9RxpBV7aYI
Omx9UKetUQIG/4nHtTKjWFY4+DojyTlje7oYn3GYwUmOpyBh/tBx7agDllI7ggfYqqi55Z7BzMIB
/4AXAtBzqTFL2fcqJY8dg0f3ntV9bImOkPwsXOpsA710n/ntCjQLDr15wZaBPY5Vhux9Vpz9I/H4
lPQj17D95efRBVMoPZsqeSP6ROY5V6519GRj41BDKFh+TW/ubTx46kaCXVkwBkD650usrUYYr6rz
+7Ozk3IpAHkhEhfgWsfTvDydRfvtX6nzgeiHMLvX4vZ2/3TAT3NjviB8X/E8DrYyLUFdzONq30JE
traHimn/HWX0VG9MaP3vg0Pkx4slnypZl3L2NhmG41rpihxjlqgLEiC4am2Y/ltA3Bg/f7bcMApK
Lj9BhYanXn9o2GC7dPgQTioEwtERema1cA2ebzWR6Q7Y/er2EaQBD1CYiNUUzxaVvkBu6EcM47QW
K0TLw95HCnqOJhF3TEejTvmaMEvh3rP6hVvrkG5zrMbPKVW5+/Ug4aXf/4Dkd7pxKjab1WVCoXBw
mLVKUUqhwb0oF9V7+Cis0cLrOQaYJyOZIxX0HiAq2vftVJrZSeizP0VAe+N6ky8BwwpJYH7NZpCy
6AlmUhJYf73wcgfEvvcO443+9F/RsrB/s6UVbKhn2AVB3ad8Nee48D3qlTMs8w1KbpAhAHfFzA33
ClRPM85th0cOI0cbILHoBqrvyrAaaenUSb/xkrmF9DJj93xLjMNVXKqnfH2tO/oYbdItBXgNppcf
JWtIeauj/ZI3VqejkGmf7iVVhSiwI+QjNaffIm+wtzCI9/zNCOcADD+npgAxF9/6Se1h00bj28Pr
77Tqh6nuqE+6rVbYuzose3RWzbUNIcN97GoOyHTCOt+NKrUI3VERsl9fIJeVfvkGV9W/MQVy7I2o
/eH61ZvUDhJMfB3RDn7i4z1QWJcGu8ZIVMMGpDJczRaDuaeN2JxaOe3tRaJ5kMQcj+ZhPK/gyMaR
DCzu/ShivSpzU61cdVxi1Ns96hKAcJB38FPCUcs+bq7qRHojYhUgXX0/GuOj3KcjUVNadtb5R9sj
aIM408aQK91OsjFvafBU/jDqV9yWR3T0Vvh3Ql9BNACos9+55+5nZDrMUya3JBp89S4qUDY139lg
wGDyW/N8OI1E+sIGK5fVbFSy9yKs/0MCOrIWW5kT5wPTbgxrLPD+pkJtuVzDzUUOdelEQ9B+LeGC
KVRjrxFGy4Rao1Og668yAqqgwkMe4Z/oYk2r3DBPmEJIA38pGIagmDeivWsrpFJHm4kk9aWc4Mtx
zg7dOcCy8OaAFUHPXuX0yshMV9FoJPTKh49P2g0a6/4iFcubiGuBXGBjS6Khifg6wcerd5Dt4fan
dalRztExZTLwo//OZb6ettDCgoaACNGf+7BCUQlrWS2OgVDdQf7uVSl/Jg3TvVnWq3Nsmq/eazwF
pz9bxBt729qNxYdi+hjlQR2S7iKjK0eLB6k/zqcIPK5uK/IdZn12qeBNQZBBR8f2GLTfT5o2XgtG
LI+N9jAeJqU74m0z/v9lvfvJM42MFEEOzpQ/Oid72vKI+5fNAcXJb0/WlneE4Lf1gA1eBAUMHcC0
Id19BpQZe98aN6n6IRgfVclKRlA/HmAZag4K5FceZ7TT7N4xBgS2f6Iyl3Bi8fdxoucwr9vb7yYY
rBaH8aaLoMwZrMf12TxBQC8vcF5BmSJY9cIWgf8vqSewAo9oPFZXBCwh5dzSMYZkHKo0EbPwVnWi
BU5UPZikeRm9+HWd9TZdIT5a9D8DC8rGrkiMizyiYeW/LRcdaJFbu+Lzz2N/Eg15eTk1Mw7hYTVr
H7kXcUhVClYqLdzP0i1mni5lcH/upi+rE4tEH/brBmoDhYEiAdOhMgWVUpUyC70CHpNSxOmc5ykn
0eE+ow1biV0EsjR2kT8j21BItKB1lnxpsTedSykqaNIS/IEMGe4vEYmcWIvyST/A0Iuubq5W8p/E
0pAWcbaR9e+gZSOreY8sLc2s2tUG43/VfjCzHBrlpZ3fAoxXyIlUyyDEHSRsjW7rp8SXehxTKNmX
z2m8AryMgzdArMTqlAOeF57L6n15TMecE+DUxthqYdLQbRLUQRBjBLcR+RGN1VHp4TmwO0Hs78H2
g35w1BEtbY60S9GTNENZXc9uHEoUqqxcw7McTVwmvaLinCQvZ8A2nVgX8bPaJemQQGA6/TIuszit
BOSI6wpt/e1q+zD4T9AkyOqsu6/ty/pBWLJgZ2SXEwdxSpIFLZhnNjBK+9T4G3hKeVayN2qRSBec
vblV2zYZSchgm0mJf8Xjgc7cvkvEg7dslbMoEELt8iBM+r8ptMH62tM+3BWJbbG9qjSchy63znT/
QCqrNyGqOxvmHV8n1x40w7LL4TxMjg33w17G3XqXJdPmIoTwlufYxWt3TSSaieUmQHwyovuqM225
BRgvHXmCAMhuxQIg4U2y9pZhybBNZvdewx2KULITZ8/+pLDmpVGlqemkr/WhA26MPk9a/acaUkuR
CsL2xTTlBj6ocjFYVxukA1Ka2logVL4lSj9SWjOFLbOGQKIfFCs90uxNYEKlZJofmxkvIxSJJbld
ao6gAQyDiVPgyM1+g4s+SRZZZ+3gzqfsZuUyqdY/bWc+WGvBf7xP0vTX87kjyIHdg6HC6N+bG6FC
F+O/A4+ky9PJjldTVSDEQT1AFaByevnEABe6ehWnD6aodFMCOIVULS1kB3VXFBp8lXKJV+F0UKti
l19WWXMJc46+veSf2yokzP7eSsduRn9RejvWNhF2iPSD3mD/R2EvOzqUk6JhahkAH34FnFCg4zzP
lsDEw2LvtBXWlB4KwJ6isXKgbprvxKUXorGNLuCrJ9bov6qERVIk10h9WKdlwt31EtbkBKY1KuVD
hiPc+Vz5L+WxgzZr0oPpRBpI18Fz0hH4JF21eLji8fay0AB+Yd40echx4TGDMKxivpoecjZVUTYr
uF9zy4hnhoqc7KvQkY8yspMkjMjJKLeefvMdeSelx3/DkG4m0jMkRlLjlTveaX0T0YYimbnP/1ih
qluSNLEYGM/XI382/moaZWrp3gDQQJWPox4Q0qescoTYPg2rt7KZYzLQqZFiJqt3yH+auYTOcMZi
DrGlTpYF6qh5Ic/MKnq37zf2/JWTx/Aa7mtaTEPzFjYOPc5IB+c2MpaLu7xojmn83Hw9qzJScbPM
F1SSk1qUnn63Ifh749jcPsEAzV2Wc2aH2gatFoJo58mZvQx4n0BiZgjNnGnOexwYu2Keh/JPFQqS
GEr7xrgBP/rItoDwfI4Vdy4D/6wh3xHgRYuUDj60vkOHidbQcWbSan+CbJRu/qrj5FvXS6VquO+o
IgSqikGKlIVgIcdaac8dFdA+4bHv9nZzaF0Akc/fYp7pxPzQt8JytbJ2IVXM4n0uuyXciFvSXV5a
Ho0stYOqCXN8hNmrnBB3CZhFGlllk5F6E/TPD+LGaOWKF/E15F1pM2jRZA+Lx3l+0iI5ktJGV39z
PuV1F4dGvx9XXeepUM7L4H/2xBKRni0i4soreVxQ7w5AAjyuGqNR9LFIZVqTiH/k1d0HcZ21fPbb
d+fylbJtUqWXbQq+ufvZxLEH06LAj/5+KJ/kegWzGGWcJ3URSly2btOySIZVQI5G/ZTxohuXCuP1
HKyIHJ3mz4d1SW4YUqO0eJ/TZOawWidUv2OauIM/xbhXXZwGwd7CV9i4/UONI3Gaf0LAjBAAkSWy
skk37Ebijciv16svSB+uQTmpJs+5qtHE9/HDm6LMe+pq7NPiCXymJSmKpL1OJRKspqw8RQr+PGyr
tswa0Srv/KEPByLrm0UQY9OCsdVmHlMPlRCWWJZR7V/BVq1QVZsPrMy5oWgbarMJo27sH3F235SE
NfdwEByyISuJ1yEKxlaNHb49PpUfI2wWRKvt555j/JhetwNGMsFpASHcftxzM5OPwv/+xc4a95zi
KG5AEWaUZeLdtcK5a1kr9ylda0ghrZwZ+5MYWgYopo7AiY4Gv5pxxJ5hCc1mI5vS9q8+y5ANVq80
bCeN3sP2jtsL8HyrX+V6OYPMi4loq7RhCe2gZgF1/K9g//OhAPI66a4OglRUKQam1MorUfrgUF7K
KExaFt6zjsKBsrT8hfc2nbcaSyw5VXFXqRC0X4H/0avZX94MF1dcPJEHR6nPZybO01XjdBqQOpfE
dAseTORqk0WrnVVpurpIR5tzTYND9B4jP8y/CQv74P1nRLv5pfpjFgujADRweMeliI56pEEkWLB7
uG7KZuzt/ymLFTYmm1IQVubMQMuqnfdt97A563dBuG6mNSlXasJ6og2wetPIVxgy+y5+kCrqVJ0E
Xym0zcvhYp+FifQCOzU2Qv2AR9MpT/cu3f0jj1QQoJF2tRWrZW34qBuoHp7YYBDOFZEzS6C+ya4b
UeXIwI/5/jEw5TiqWjbp4+dRwXU31smoDz2nZ9TfVMdgsUiDaQC3351CC9hrlguqdELtb7B0v/LP
26SOLp4bcx57lCXwcp9usX83Erzv6OtyVv1HL6JVc/J6Zt8io0QYNO59ue0WQf71N2PcoRBbpa5C
Siexf/FIc2QfaEWhQw13Y0yatNduD+v6W5AYR/ZARWSNkrxgWI8qmQIjbyHMc0GUnBg5JqW0nQna
OFkiWZcPfSFFGkaL0+QRTCBSMXu1eL2wAgK/8/P7FONnBS+mW1axyqIAc/sw00gLe6eMcyxut8Ti
e81tn6pyL+z/sSdUdW6zHpy5WuFOXI0PMzONYk5BHIEaQPCkniBq48VWv8F9/xvGhxaTp7SZu7JA
a+WvRYYoNUTQP/+dcDmMoQ48tq/U7gNZroQYWGleuyO2g8/+5V6w0rqAf4e76AnF231Vn5WmTs09
ckLmjEZUmgWfhSkBBc2SfIdwd2WzMVtrNtS1ORpQRxr0l8GxjP90vkWC7jwf9ymLy+olNN1Ra6QL
0N5tJn49zOvXDWu4M0ywN4z1DNYMylNFbnQ4bvroVHV8XshdBpc4cpOCAEA1r82iaR9rSD69DaQb
p1tq5utMdruX6RnLzoRM90ACLuEcA+xpxA3UVLVFOjESL5cqv66jHQHr5Ttpq9nl/OHF9fM9Cypm
Kf1ZVdT4zvNddDsyxnNhUXWZwjtg5KHa9yPdF2ml5+RMTFFdoXfcGel0m/4UVMiv9F6+JNXaI7f4
M05CxpO8qEskF2Y/BCE5gM9705G4zjdwy4XX1nFLOVp4t7jWwmTigsFlX6Awz8hbE3DpUqsCM2bF
N+bhJuSIie6ZNdYHJsk8Y7pKcptWDreauvSJm8aAUUVxbL7NmfvDcEjIWS+Rzr9OfiA6qCn91GW3
aeqmvRQYCiGcU9C33tvHtgN4o68512DHQ+r/4iRaRd4LnbW3aJV6SbttTTCD8NJe1PxkwD74Z4Sc
gCxyYNYqEIZ3d7OEtbUzorV7HmojfO9Bd+PT+9GqH1+OGxfDseigYl4rcllgvlrPqWUqDbHmERR/
cfzxbF+LKAfx2Bf8bj3UcDV/Yx+j9iJp7+rTP9xsEfPKsEwFyYgrhzq0AsmzKfyENcDRPn5MUyxi
s7/rMRe3zkhX9atM/DAizetVG9YYGa/9+mLoSTm+XCEZg9xXm1T1T92bmQQTNweWNK98PAQWAa/x
LCbNGYtfwth0yYBwNquM86d9Jj3+PfNn13m+SvGozinqSIMtrK4+NAckq+4D6E4EacgpTIjrKCMd
TUDbqg0NGWK0lejBxs6Y4Wp1UzqX2chwEbLp9VahhikXP18fy/9H8tz0A+sZAng0HdvHeLf1xurS
7xEZpDWQ6CK8oJByBDWeFdjQB07k/qAIUm3F5AJu9ewNIszqWqHWJ0zN75naIj2vlJW/PSb0As1j
2TI+Hp4N+bVUO4TUugkztFkvUZVLFrv2cRevPVYd50n3aP8MJZI9vHBco2KmTYAImI6u2BGoQKZa
3C8j/Yto/lBh+Jn/Zjzah3GJ+0+unEvLLcI/NKNbRuxJ3nGy5d8VEmd2zQZLOSi47nmeoL14gbsJ
JUNHRkfuzHnkrk02gCmiOe5FCCczB8V19H8iYDxJoK6UlxMvE6zOq0gzUl6AGjRzmmClOhP7NEpU
A5qG+ZzD5mSf0B8i25ihzkOBa06x5LRUohNWqPIzaGOWag69mjGFhnMsbOoyGVo1fXiBgoZNUtb/
uklh8iKZmeuVjQMLpDuCUns/uRZK7t3urF8Jf6xwJ0vtTk4dpDtmGBvhD+ed6GtNQ9V0EfMdu7SX
1K44dj5vmywe8l+04s+85GRXPeskd+CSXrjkXcCEa686vjPHYhrED6j2JMimYRpMoSaoD6EwP8RO
Hs3gT933ueP3AuhRU0/KCrCczNruQ2RQbSbVgF25aSWD8HlPdXqwBq7XJ9wKWKZaCLWLZOwoPMcW
WSnI2ydMwghv7KcR8BCoB6u6PITsVtd739W8t3L30KoCe6nbC55EXSlFJucZcZFkINpDPVqYrhT+
A0di1sd169HWH9zFXd3DpPxvL9UPItbxAhB9kPm0UP8mGdMYkV7n6bVI04uolkBa96X++jJ7WGhe
zXjB77+QsCLIJAWBJzEWh0MOjYmsQ1jtXVx6/GOGQT2ipMs5eOiMmPptniNYVeg1BV3sAZxYLKW5
tNW8+ZhgIptISMelQxQoyXyf9bkBavYjzObBMoQLMTxUnP8sOZmjg2n2X8crwutteMQAWQh5ZW/p
0Gh04sdcT3P1yoAql3vAelFU5sRIjg+IB57iGjuZn/V8YIvxVsNoXk0Zwv2vwbR5thyiMyTTW//y
7uiQAZIigUCOsX72h1Z0OYY8zKqxpwAF5CtFHznuUoODSRR/XmHjegmJfws1F/zGdRu4lpR8Xwzw
tSz+C9ncg4d4uxvmDUdge7GtM/xzLX76py6edvHTx9/mH1Xjct+OTGYGmvoT7fQPxYGJznyxJLOM
6gjT9OG0Wa/eeXouHwZrFXGrcXcOOcl6m3TUktKsAoGUkRtLgwTZ126jwhojhaeSu4bhhoMW1h+r
rfq5yrsG8kUYszoUfj8/fJsEwjDbY0BJqdutQvqAUFfdXyVzZ1W6MC/Ar1/BPxVG19hJqwSB+8ZT
gob9+9vKJEqqEsWIoSoGBsBIicZLbBNEK2lZpJdDeSNNGyDPYNRe3cYOyToTCfnc2DE7cmSWqhdt
ckgRVFIZMflIRHfu7HFabCcQvONXTW5vcO4hzh0jFeqhSBgvYv07hMdp2XRdWROsizIv1Z5Hkpqx
NqYxg4rBA2ZNjalcy97znH64BzzYHd6VUDNosd5Yf6W75eB/t2kzgIFYWeLQlWfXhHSDp1Os2Xvu
IC1S9S/7S3kJFjwlZCQgusRdlbU0ylabc59v2PJkUmG6sE1zU/Pn4pCMx/y/8lV4YK2vEogoU9Cv
0vCQvz+9tc5APXSCoylfrP0RmXO5b/Reu3RkacC4JYt1y24cGarZRD9T+LEmM1Rn+giutlrP8DIV
HcZ09EwITg+cDFFC51wToMdsKBxNdNNjHGZRPueTWHRF6bfHB9vIuN1vJP+NmuSuIuzTyWCVHKKW
pkF7vT2oOdVd082UNatUSiK3Bd6gO8IFMwv+4hQRs5zR/3dIOdN4tYd0pNwRFa1ZF0hL9LHAWzvM
Rx9swy7PynmHLbILO0clFbEBnOU+yjIOQENsecZJMz0s8tTLKQeTZvBFAljjc0QRMhcxkUS4+NJw
lAnmMMyEyRALp//DHNr9tGX8BrU+lCidYZ5c5Er1zInIwN+sV3YNTYbDBWJda2IH6u/DKlpGgLUa
Di/mpTnXiVfvwWNneZJSuPt1qXJ2KcuA5TRZN1esGAt8u0cKGa6inmR/xmvYNqBL6kT8AmlMc2QH
iFSe0F0JqkGY9hGGT8tLJjgRdrRiscQj3mvlgIo3AE8ByRgn+SBnhiahRV5632G1M9Un++9d7ph2
jqdV1tKe8WPeMUkK/Vh+URhGl2oii9ts7wj5mGJb7busWdIq2rhTz5GXofF4OB+uVY85hottUqlE
d5/MDJi1b8yhKSvx5gcIc7o2jCXWYbOjV/2f6srjSOfCBkfiMenMT2zuMlh5nCalQklitb+RYI8o
cTKJpHXzQpqK5Lk6wz1dKu88m7pzd3phenp2IFBHMTH8jupmvguuYo9DhvyzVwSDlSpuvo56+Vbf
eiP99vGPSJ+TSmOeUGXzbYBUvSqEd2baK1w46g+2zdY/QPuHZzhjPdyhnaxB07VHZMLkLMwZOUTr
x8p1O3mmBUMsjw0koZpBZO213f0q5cWfeAmLDQhUnlIf0M3aPCfWFSXWz2gQzUQAUlpTEKMKczvJ
E8UL5ywC2uK4Omks/U7o8Ncm9l2GjrHxRrg/VfxiLEOs/MKhLJRLg/b9YaNhYwK+iV62gItcFkAo
tE3YZXYOxGGm9kmlrg3Hguk7szH2b4ergsdQYeIpSvaYHEPXxvIa1lfi0tq4M7P6IaYvc0J6WEsN
TNxznbSYSJnJNny/7AVNUWpeZuaigloUEtvwvV1ffDboFK8Gp5ZXMnv3/ZwYTq6sBpLS2qru+4d5
aSeR17yKoSn4GeyHhZOXX/sEm79b/pDDsz+hb4GEsxa6mEs8guUgqHS4yWahqBj+Bx7FL3FoJ+KU
zHtirv6IKJpr2PUPHwTCMtw8EgyP8TiFuqese5e1Aks6kc+33I10y8iOO4cTC1N6sWIcRAiB2ok6
rBPmm1/qFqOHTFBk5cyrZz3iZ3RUYTEq/IBVY8S/z2wFGj//Vtwv9DXNTzKy5YrUC5M8+qFz+1Ba
eft7BjM+w4pdz96FgIyww1sQB8ycPS13J8ypn/6HIpkTzoE40vmBouxNN8qeO+19KxptMDWnMaYt
+f9omOv6O7PLs/kcF0XPBDMcYCG+hZZZeTJxeC9Xj9VqTEKeyufr0G2fLjwCcpeR7PicZVbr0du8
Jqi508yGTUE/raFKjXK24YjlOdeM8Z5copcnYR6YbPsEj17ih09G0Q+Vo9cE8EyGKqd/rPHZeZMN
rBFA1jWs0Okz3pmmeIzcNoJ29FlZKrHd2GFEq+vA0t6pdO0egR9cFDKx6biSeiPgLIKPJOVrtIAR
ClohgP8V7FiO4VDremqceeIDdusF8PR1NKUUSStpcfSwzRCsihtJ8qUWRkoV16z70P4v7Q4nab3/
9AhV9yvNoS9ZdcDbSNJf5zXiC1qIQaVz4OJNlV9RZxP8h1nCdBLXOI5dX2GXyb51P5SDOgvov+VZ
osiE52GutiGhat1ZjLy7bWxwAtgSEOYJvz6EQUNlhUvFgHbfVzy53bAIcCTmGWG8xfoM96yqR6L4
dR8044LuU3oqamozV3BzdVgSnw1UZOqUoXk1WSeBMJ/PdFL7dElYiRqySTaz2J8TDTCSTMXoKiAM
EqIAGx/i2aX/V73pgvOvBhDY40gMG9rJCmaIkTVZPUmQBbGQa5iDm8oOtH4gHI06s0bsphfbhGyf
2PZ0Nq93PPGlQpNB66bfPHfJX0ukqeTng618K+/yVNhqP7FuJV77EB2H45WBd0DOJ9L5BrQr+GBD
xeL5x7qWxMcb2OR63oUTAI5OeOUTF1qmN7hrXHytnDOoKvNt6nVrr3oO7M66ZOff4NrsI0mA4JtD
H4xejD6m3JjxKS3CNEbSxdjwRVT9iYb1eYkMyRV0tkVwQOkRerMcFzO3H/MCaOEmzCAumuNKK+ty
r+j0u6y2jGBzNNaR0e74KCNjYDBM9NfmTGRhaT6Oyh55l6NpWM4YHE4uo5pmcSyeo9KuD7dwqKMX
n3ZtIBilhttEhl+Mgj0/ztAU5B6llQ8GH3PSgonzXiOD+WCB6C+DMWgsVF+L050MPkh0FiNWeRAX
ggK2+uPWW0xBlvvCoZSCImW/v2x5Ty9v5IeBunuVsudNiLZclULr63uRvcXMl1zjpoGyNN/kiGrT
hxux9S+ENIhIijmEBRKRBQvxIVU+3juRAA34Ij0f1dTQl94kjBrz0GFaKSs/99ruuNQzoprGOYMI
InFclTNOPx0GrYRKe9yMhZcKmTX4cDPp+xrr6qo21Y+LRfIVkg5LvSrLYoja3DtA4+qUj2m4H38q
lB+QjJU1lMjYAzfBRYZ4h7BE/wQ/KxoKdX903yzEGw7kRvROHe+zKYYWO/+2/1JBdELGl9HOA8t3
+hrqyL0vlagadeVlNY7qea75dfrbmw/RvS1ga6kqCCkQ/JIbjBJVOvyhhRiq63KZT0SGtVWqgPu9
h8eagrfovRsiatPgsUoZdhZM2rUvn6/kdeWGccLHrDcu2KDr8PA+S2Opss5wCeTc3YuhKAVTVnl0
sF0UC4fhKecjttLP9chTxy4+NtWdjH98lUYXp+QXTRvPSpfSBFvkms8UvDhofgnaMiPnrE+f1ln9
dmeZUuNeHOHJ4fmcb29pPLBu8+MkJ/aV31X8jHXwQ+ZsVWFMNRcBvaacYmMfc7zxyU5ffVCvP1jT
+v/5Z0vz1inSmlImGfXgbXvAmLoQdCmPT3KVvJoUhV2LgzGY/AQHgLyuGFBFs0hg4pIJtUEHzRuK
IG52L2foslvuR0U6yqTR6xFr1tI/YuBOziYBDKczIQ7T6wU7L5As/W2jcdZteu45ruCO7Yw24/ka
KEanefrr+N2kLEQa/tS81Taag70T7LRF9x6hOFHQOau6rRzfgTnnFDeokHfAuvpo8kexzVykhLfL
f+lJE9I020MRzE3cWhI7uw7jfDO+M9aIyNwI/MZ9lbxC7Cv5DaZ1laQtYTIR/WExKA65f297wHx9
IyS+kigwIMLiEG2RiKD8Y/LDL6OUPhzSg06+bOpo5Mq309+TF7PevGDFtb1DYdQBa43Py2pYPRt5
YKU2A8Elub4TgsdYCLQ0wOmlA+i8WEa53/KV/7d7/rkNcHJPZcx9HT0sOQVrxLrCUHtnTTzPhafq
4t8uXacxIekn2R5S+fM48kmCb6BU7b4bjL0a/TpXSc8TRWqLPNdUpriIta6nnC4b7pupdgcyzlGf
QuTcgkyygxY8+ZNpgeWUNitAxeMOOdyrbom296nSPPTkFfqnYPjxmS/RSqIZRZw2eJbm9EldLB/j
8bhlclBVaruw6It5sPqjWdF/s4eEZukE/4okgSxAAuQlUXfFyyVoATYUJDQmJSQuOPtGZ1WySl8L
xR6fd8GFOAJ/vQRLbdz1oYJK8QMREJXEfEWCs1wI3R7bja2sHdHLnsG1rEUadqhunaM0HkBJ5wjy
rksnizrHvBwAnKG9htarXEEQW9mGUTcwvdQOdN69lz5NPvTECsuPJZMHvxL88ixCswiNxOIzGrMC
3kAW5NfmzXj+Yyidd83WyCkLxbKgj0t2xp1tjxdSy9+4S/8g9OaDtGANk6j0wnaqustF/PpnPOyf
WvE5tQoWNI8gejifip55mtM0ZrEoeiyyPXX3MGIrU0+O0BWj1WKIh1N0v7Q+Cl2+7UofNa02GdGV
kKRTgLBbwfxpr6ocoujYtqfalJ2Ft/d55FaDm19AZzbCh0u+TAPZcAvAAr3z7HhO6UYy9kyRavzr
2ET4xLm/2DClgaryp2dnqw9R509/dvtpiNBMXzwH1cKxTru8tRBisEkM53jX9nuAgkb20RiAihL3
qGglWs1mHLDFjezkONn8YoYX4Mx1LeREoy5gtlVz2T5b2kNgB58sfXKC+uyBMdPHhTmp0G8ydokA
3UKVFWrJJIogm5veWyj/loRnqeegODCEvoAmNX+KoGiNErmUMyPOFnQUV0adqWRGZD82MMPPZdJL
mNyPs9U9i4O0dyKYcf0eFa4MSLUoiDdXYRjJUfB/anzjYdcCNAcPcPKvagiNXYhaG+9ueDrfUZBD
CVLrlKN7/FkJ9F/70l2N+2rG3OFF4bNmXVSnjIO3iX5f8piieAMMObhelWhgJOC73c+sKhXsvfcj
Sd5UROoG4yorbsqRoV0s4tYuTcv5zYGp7SeeqmNrACF6DAy/djMJkhU1PyS94m4E7eO8dYqDmZQm
chwxGzO0LZ3yocqUH2aCEVm3ZPR4wcVcwnXEJjW7fEgohn7xWq3SCg9QI61c6bkDKNRHIzt1KVC6
Eam+PYlGnLR8tWWJE5MCPjJl7uPiooJw+AnyF5j76ANDKtwsZIauJc3h6KxF60y7hrWR1pTQBUAS
7n0TVauWWKkjC0Uja68vneXz/jmbDxSVLQIzQgh7Ae4EmlNOolEESaRdUtjLpWOIsAqJGvGyvBbi
+7nfsSr7uGPYO6Ep36BN1i0qKY6ZRCdRjQjBcoB7jR2ZONbvz/YMm0lFpbSn9Dtv/kYKPhyiOUlk
WunoUdjcNbcIqzjsW+EcBzga8yH/O0QdTxRii33MFtglwDhtFB+vaw/Qn5b0uCNzcbDCU8t1a/Vo
dPsbDNtBQsk3WGy7SiAQpjJ53Bbk0pN86azFtbpRyWeTYceDVkTmU79tNl/L1D3ztFWVo8mzjbcr
myEXb6PrIAMqFVeXVoYvgMFbAQyzuibciKNTZ6h+TwEQQsEj/lPf3pmGm11itx6poDQjwQi3XL3y
wmrsL3p33N+Cpfy0Q2+ZDIugk6efuQhFJ1mj0FrZsDd4uWc2RXJFK224UqBwsAJGzaHbiJ+wT5Zb
EHnvotJIPCu2WCn29bthz515VPS4pvS/s4Q1vrP97nsMvmBsqoHbhW8DrA4OcFG+W/EV2AN21tV2
IhoRM7ioXhfQSLSVbHigEmzfEesv0q7zpGHvDlfUHykFATX5gtYgem43tryIVLqto5GrxT3luFp2
dsemVXppez/qi2Z0vHvHwK52XUDJjrAKAskVAoL/G6CS4CGn86W81JhsV3rhg+AMANjWlJ36/sk/
Io/EklfTIrZLeeHy3CZp/afEeeXmBY1anh61aXghoaRb5SKZi/GkmvxpIeyvnUAbuuV/H/L7fhPs
Ed+Oz7H1pquPiKqysb9EYZ4jeBE+hAaHOXVtCfnFZVW+MiWKcouQS7lQtdU7WQfNHdQgpfTtTSW1
BNM6a2eU7w0zoRt2T5VaEDzL16IFlgcD8ApvFX9rwOv1j8kMBOM8RCS1/U3dBNYSh/tJ1vKVqM9f
XANDXVl/lE5A7Gggt3RVhbtZ2uadPBe7C3w6EFbtwT1I48eIPR2v8vMgoLs/jXM6Ckv8e862Yi0D
g2ery9R7XfCvwM0VSmDcCyT4p6hWZddYOjjoRXcXMGQcSlnddM3OAgrpIzGbaFOQfPQH2xHRzi1C
+/2yAHj/Jbatha/yPq6ErLW9RUvnKB+FNQuCA1seRa4PL6S+rRcBK+dM0Jg6eCAujuPdWsm6gtXn
KdNDYnaspcAniYDcgDQqf6ZdUdVnho88edF0JI3BOUlBCPWW8c4Hn0K7kS41Tv/x8isdSGrICanR
WBipRAwln0Qpg8f2lLHHc9vtFESEkgQXexH7nql0tfg2F8bdtrLd5og/LdGFcgVQso7rL9Milure
im4DMFug9b6Bfa43dE5pMTCHdfVRfnGZdZ4biCvdQiJJAdbSfmEWo9kZoUXs4vs2pdz83A6XTNEV
YEbxMzVPTAeBuPZv4akmLHfvMq9klc2DfvIfNyt3XwvbU5EUlxVkCUYdNjx4z+YPxatP+0UAwjg0
nM+a+bw5natY09u7ZTymUyinFbOj9O1530oFRNdU38Bldumz9NVXVYQQHkWLoC8u9yigUIuuFXJr
yjbh2kbYDTuEpV4OFsOv8mQW3TQhSqqNVCcxaYMcYCFB5y8pZyt0f7j1tazhUU/BiUjgZ7T2BdDv
TNrdZnSticuYGsZCB4Jum7RTEfXZkO0fluTrafhI9FO1pVrcBNzgZCIgbtstGCCbOeTfQETdp0Jw
Bsy5s4UbsW0GxuOlVFo+y4zs6ZGXJm6mJEza1+bpwv/C+L2r7FZFp+75OicdO6XmgEnd49myfcuS
KEMMHeqjG7BxAqsJTe0ua4xXHohPQNTCjEZ7ASxAWvet3EUVFypCIh5f2Hu6RR5ZyFRKcPlvKhh8
hvKq+jwzbCywsVRUfu9WtrW2jLd11yxnbMe5UJHJm+18MWt/XwbVNH5hK/ZAWLSMA52/CVMl15vg
oWMS2f7hFqMgJiuU7Q8/abvmvTAoOrMexPQg9OhUeBIOhYYtMq0pyLa4B5L9mlisk3LBdTSzCauP
0IP3OBtEaCfR3I5Vp/Idpp65xonXvsuETXrsW2xa2DorxoraPt+F6Oaf1IgyssP/V/9aoq2TkziC
2B4grOJet9PQjZjHqcojBwXuXwGKGFhuowTnnyg4tKQXnLoQj6GNFCxLdRXI7jUVNaFOPH129hd+
ZeWysRT9bFnG9Pzf9VTvipwybuLJkt6Rl7hDybM4WDK8194qV+SwZ7Nt+5vnOkbZWj0+/al5smMz
sBF1yt1G6oxkBAEyqosiqze4LNPaJtlDqEIAP05pbcwPsA2D7+Xc/vf4ysfphjc5mNgxhJIkUN6r
onF7aOXcjuJKeHX0UhJXj82pGgi95BTMtlD8BYuheHPJm6knEFPxY1yynW/ExIUwUdobI8DBFNEu
XNNPYMHOsMKnlHQ2QtNLkws7ppyBYGGFoEFwOK61Fb/Bs1gvUefIPn1gZuvIkIM5641+rPQvQPhr
VZCfVGLW2TmXr7NHTJ42kSQhRnqBs6AX4jELKtIU5rqZQ5rKC0opouq4UE0NCYfBHvjLczEGP9ot
UPUeq/U79yWk4KT69OOjL4PAdF9GaClxKC1LoLEeu3a47em1b2TZERMbB5SjMdJUnsoSzdnBOveM
Q0JsY481ZupIamQ4os0KKhEd7pik1Z15ySCUCerwvIC8Kl16isyzrIgD2aSZJFP5luM3wUdCdkh0
FGdrsDypQC6kTQdTnf56QIErY1iyaRefRsM19vuE7Mc2VTjGJh64rPs6dPgylZq+TklqR1hC8yJq
4SPt1jKiH1T6X0lLvNNAXLMsgI/Qc43gqGgAufuq4EcH/slvoY060U2z+9XVSWponuAwJIIiBU+H
/mcmj8C+PV60am1jL8k2QKRRkcfwv5csWO5z0n+Wudd3WZLwmr0zh0UUhotYrkTqOTl4Md4LDvFl
C3D/ute5UwsAyxBf9Q1pgDLE2sGY2X65hQ9Y+v91Ca8CbEx7K4VEiEhVBz/YsoOQB6TTyEqyhnqU
8sX/3E6soTUnivxhxz0w7w6vVNGX9zebY76+bXOL/Ee6adAebz7So9W2MAsB2KfAsqHP/lLrChGC
c+aITlXpoQU4WYQktXPyjcI3q3CoWJaWUpxKqvcmynEbWLzKprBP+PMjHQfaiLIYnV0kSw7oeitV
EiMcA9pZlo4uxuqbBbRRyUs/PHE19DqbC64dbsGhBkIN1PVguLGBbP1lbQUN0dsqO/Qbm8IHoIKu
trw9xaJca2LlHsvsX9xyWSRT+NlAr76+STvvfoZ9cc5qlce4T2sMwOgEvsdYb9jNnm/os1OeOfII
9yWmzlg3DamJkiqIPDVK/35KvvqUHk4WQ84jSvt5FRO/8B+xkJ3odtbdEwJnDu8pqPfcLz7lucsm
EiAv86iit/9/jq81W/AZ0fuzEIH43YlPLY1loNx3BR7koqa7Q55YuzRtkfS4eml+nvLX6QbPltTP
9/Apg8BLuGsniqWXS27jIIA79Qf6z7fqJ8iPqn26iVasKfniIeHYFXwEACoNWNLqNQDhff7KcYOn
u7S7XxWl2fumFAfBbKfCSa4SK/xfoCc589q3IEAfjmvekPYPazjtN1LEZqyX/La8aZe3pkIl/4ri
A+xUgM1pTWfgXMsDeb6JluXTIvuLeH5735egzvRvM0q/p3bIfNVBJ8Fz1s8PKwU2qtqaysxJpCia
6e5NnSGGqZYz0gsyUG1THNGG0OmQmDPweqx+YRMYA692uF1QrRdimdrykQBNpYcNPVRpFBKH7+V5
zjNX4uGq2N+QDHuqPoF7JEne9SzAGguxgb+HBt9Sh7YuezikfZC+wc8syIY4qLEFj2yH0Pj5TV0y
lXxIxdbJRkBAZ08EwgYcHisLMHU6SkuR97M6xqikGKO4Xxy0xLSMurxFKU+5WOGCZsotBanB9WTg
rGPVDyp9Xe2XrmrxjLvPavZiFPwInXpv4+p39rVYU1j+qfdGMNI2hmcrY/ci0V9YAPb/ejMVXgIh
ymNlNFcwtXx8kkNV7cewgJurCR08fCsx2ZEMGYT4l/Nh0G/IVd4t0PumnVHpuSqVsoj9B7AoiH09
YZZ5IulKdjfEnsuAmYj3KVcqV1vWn7Oxm772kvI5jblaXF68AgwKHfFSUeP5bfN9Zc+82hG3Bjtd
qOKwNGEwYA2Af3SMVMfH47LPcTXxG9PkqR5tuwYq0e0wqWFUKnF7DZGhLnHjDp9pua0Vv2q5Dmwf
H6tR3pkm8qE/QjEHxyUWYt5Fb3PtuKGgiNz1jEEJ/t55MYW1DUgZyXOrJQ49wpymzgQf8Nwck5SA
RQEDP9cJTYrpfu29LiwlZzYSPT88MpHWYrxms+MP3+PWs0m/Xa3HQnkuiVjQWVMsZKzmBuKbKlgD
AfDFPRx8IM6chnZWO6+sfu1O66nhSlPvpfvLKmXjCcFDUZLpLn2uYYxGQ+6tZaz4QUxZSUTua+ke
G+u3ECAzDSrdWqgztQADa6CghQgHQ+QWxjmLAsbIOl8quzDMkeCOmILZVl4Pvt4yBOLiHIP3pe+6
AiIvNDeag2vJPRl5ZLt9uc6/YHsNwPtlU31t7v7/ZCJMzRiA6teZMPo0jTabwWRGNEhPVKBn1wPY
DjyYBxwIR/8y9m2/QMNAu4sBsVsdQsjg3fO5mP8/wUoaAnFlzE0wZBx4FmiRFC/GF5RNFKMKFKPr
RcUP9Dz1FGRBef9Tb4+pEfe0GfcO0lUYkjAIxHAGMNxcYG8dA2rMbfNUWFLs+bkYJ9uuCcDfhZWS
ic0AYbTnPkt+Ze1rFVchHYEJGUL+UyjHa7D672zrOwddvWW0vAvZmGSN3Uze8IoHvk+a4YrJdj63
Ng2jDpmTiUpb1NaFUJziBbAGPG/v5Xsm85RwO/4yR9sKWkREHgB9hhH+zXTF41WjDl0PICWXWfm+
b2tu4DP+UPwhld9K8jBIyVHyr2xn9WNkxJawbO3Jq+lC1U8yoI+YaQFHRtOGkXf2uMSD4ZTnPrZd
RVfrYcNArzPtm685FHpWt7XamLeKdD2JUXn3jndmC5p5+S/LTFp9U1ec29iBtaCJUzrlDX6RGgbw
cLruhQqDiPJ9/5BgplTN5rUGuCzxRqEk2ig2n3r4EbveblC7vbf5N+O0l4gjFNawanW1qaVTcHYc
G2PyF5YpiKeZ/wlSpnl8ccRXLJ/IH1gAtEmRMhorXlZFXkOk/zxouY9XCnALU1nBeUEu8r4c8AKx
q2V/CzGxjzYcHID2rsMckveGdMMbepMhpFjykM4KMx9HdCPyJ9bohhXipNY3M4JiQflYGJXA1R9J
1nMtlKaPDvGi/k4/YmykTakwAAxCpERhfK7qDYPty3xIOuXLzG9rDKkFlPCa9orHyybhkKJzF/Z3
7mBinvsGdrVLgi88+AETDgqxC1WL+2OQueuGaJx5dl2nQLY4ACzlTZI8B90UgWUOlH4yRXjvljiN
JWeXjTqtygG4uGC1X2LYikC/7z2ouzqeTm0lwoTEusxeLPj/1hur6pnYWIKpZ67TaSeRvbKs9Bsp
lMcIS0AmpCz3JKqrwoSAYoUyLwYGcQUjmXQBsPyd0w0/aN6DoAqQIsuxqF7KfYOVh6X35wJs9avK
epS+P9w9NAp1gQJRq9Yd14J9v4A0IZFsKUJNsh4i/gTbT2NfTjBh21JGR6nnHc+4KkNDb/qNcEkA
mdS6WW3wClgrn2GL7sKqPtYYCtx9TNtoZ/zCFEPLrNt17j1KSjG1aZgETI7u4Y98ZLVXAz5vyVBy
0DVLQSZlsIaAvklE/zIMg210UoNDY2Qa81A6IT+Jycrbrycjd79qhiBxYRwhwh9Bv9z0aFS6A+GL
BACd8PZcR2lXyhQSNYnX9LbY0hhIjRlLgAga6TF7ejq8pJBK2uH1qwM5ZJKekccrE9EdWyzl1xIG
XQQ2hJYEaLGoXcpzUxmZsLCt75MPynbjRl3Y1gkyoJQgtqFY3dZiuZbMv7dsO25GEO08KwUL8X84
MGYKQDbQSlcSGO94d8DnbNd0X52C9bWYSMMKlfOVjCeOkYjPhJIrhBqTheezlDnNgLc9jlkkeq2W
Wh3+jshKK+Q6cx8mjXLAlxPZhgeoYbFx9yznNvGJva+HUX/JDspS+FO7Oj8olGLvfpQQxr1ChgoS
RGZp7DOiObxVs1tqpEm2RYFu8YdAGsNPMx4M5cJUyyQ9Rp9qYpP2NCOu7wUX+VmrKuMB2EdfolBd
qJOKugiu66D40wkKOu15fLsp7nhkE/MFQyVLkxy9NxcgahTC5Gck8NPFaGN72e2EHuTJ8RIraLxd
HpcLVV89Z+I4ZncevPgfdTWZ61Z9XzPi9Bf8bOh5nXNuvDZAm6iG0Nv9kB1usVfenh4vO7E0vJA6
uvMMLvAp5zbvqhFRN940myw5ni7m5l2oqia9T+PoYDEo/Aw0uZZ3bmi7mzzTRT0iPK+OwEbBP10L
WRi+t93m0/MU/LvyWydCdUvYB2RwBgOFK37a8p8J6dG5Mg5LoesZG+xjT5zH4m1fR/ckT/dAOeB8
eQwg64zAmIGXCSEYO2K4bqnG2Gbn4R2WjvFtaEfBRub/gknJPfOWKKUjOCXji4frztcY7C2dt1jE
ikAjosUqmfaaaJGg1WqNwJ+Tl3wYDcJLz5+Ol1ZB2Eb7wtwaPFFBuUX0jJH4BAPEy3DFg+aQKLjL
f1Lh11hvtErzC1GQvXodhJRXhS2qbbvtiPHQkt75MK26+UT5XP6jbHPnc0o6f3hvRlUfbAHWWNZR
zDq762bUgeAS5zqZvjfOAVHbt2d/u5dc5VxOWVIgQ5V68Lxf344H57PPmbgm2LuCNMANX+DaLqPa
zRj5dIPYtXMErAEwqdOphbRip1Y//4sj2xjbUe+qTTgCetWe9ywIiXzRnfXEW8QGF2s1PmDkYcqA
bUS7fOVwaqwIIrrX8mmBP7EW5Wfwi5eAytj6wlsn9UyJV67I1+eZxyfzfjSt5PA/+xJ6FsEUNI8h
INZbw9h8nh4I1oQqc6SMHNteaMV8aZ15bDaMKmK9+mkuX2LhLBq5NND1U0++NZXDmNg2UWoiQOys
E+Hbv9NcuTaubIwmTP7mpWVxAoNLlMEmRfh81RDzhosV1uC+p3ra5blSY6dMANSnKE6J1SWEqlP/
j1e73zPWHr9Otyaoz0wvlmv7Fxm4JdTNx0nByRHTPNUIEUvEgoONvOsZE3pSlOzht1ZVOFAFRbiv
4lSt9mUrvawL1qXvBBv4n0zc+cMGvHmOzQ/7deBZW4PUWAAcV7a9nh/SzuV0y6ym3ggavj2reHo+
PnlmOmvjPXblKZsqKsOWTkJgRiCPHKa64Qv8WRnzQnvnEO18BkSR1Vq8v3ABYwyLBPrthRjS7x5i
BskVoJPJuYygUp/9Q9/qbcIBrCT2CJrXw9IHlEnXbcZLgUoEkFjompqPAMrQSn5dKATRHfcaB9ys
cDjP7Q5euUFewPlh7RLFX1uA2kxbq9JNuxtMfpwiNqfhFNu+DDm7fyke6eOBJuQnPZPxfS9SR3pM
x2MfiqEIreH7QNvIO8CJ6bFLcIR9HbZ6pZCkpoAH9KxCj+XI3asptJKU/bsW/lLrbdg0QUiaz1hC
471MYr5ygUjaC+I/alZwukcbetCv6ZEjDruRamwMNytZ1ZUVVsjaPQaOCG7iJ7ZNcWtAMul9NTXv
m8a2VopHuL5AiMMKQ15ORuynLTqb3y7RL+qVnmy9Bw9XtNU3ylfBuGEBulcLoPdFuNrESfxJBHsT
pbs5SXk8eqtHgdIbqU+bdR9z04kivvfA1OBIZ7cM+5q6OA5ZXk14M6v/mtvyMz32Y7b2lCvw/tTF
yulSqkCYPQpZ2erbxg+zdtO5+eagf+C6JWe7dEQw7M6hFFWjPb+jLqHtOO9FVSx9mYNwOGP5+9xs
lzXvjV0PjHLkciUZBo5ir4nCyCrm6zzM9ZNE/W9iVOosVgDksDMm7DmLlxymToWqUTpIm+LbQPEL
EumdR6a4SNQVUSluU+LkclUdVBPA5cgL1GshQ9Xqr/Lde+CYIE49YEsH+m1bDK07uRmhZwj+k1pn
rrJjXp1ScYoqJy5+JcGC4IO/bPssJxWLwvYLSwDUFSlU4uJ7F2aj5ziEYRyh5rABvqMedh1cVaQy
gir6odhMby53+TgGcPkvCitG/3oPlIuU715guAgfdceOnmZZu2gTWJ6xfDxp0JnokSY/kK/C52Ij
GzE7MBbLKhlRkyALmjrqcWVQv8cC+EgK0AIClQ5iFQEFyk3SMQ6r9fHuEsSn0Ha7FHGtV6GQdVFu
vNM7qnYypSEkP2ELHP7Ne9rF2OJtKVcSO7qo1s8dRaoD9qmsg3G4x5grAT/gSAcJ2Fsbf1i0KgYt
GHNnstIaB2/9V6jiDGBmzVYQ3YLHsasoP51tSM+KgxXH077zh+O4wn3LTwv8jym3ol19edehkH6p
/NYG7jY5xfTTXlm1YKIQbE8gXmAPP2qmSE1PGz2+fIAVeBPLqqWMydaqnhqCvaiOh1IPnUYHFB+V
o76B203fXTtXBesVaxOxtjXjaNHgKVb3v+uKNMs+0dbe+daRvZpav5Y/+ZdthN7PoMVJIMQttV/g
5aHNcNSeZtkVrlduHJfhWOlBK3vKgWFC9o6NUG3bs8P+SY3vd1lc0ESbFMao//UXR2DClj9v+QPR
F9QfQTIivxehAxrp2g3EjfE/ve+7a2w8s7WmWfsJk7QwTQwYdn+PooRzJ7wmq3s/lR23zgEXaSq4
/jI1nJ5BuGIMgs0L0hcNgMhhSJny27lFuYlGVYZO5LHqKQ0azayx9oOGGIpvWtwsVFB5ELFSK2SL
STImTpblGWuvbTtS2sMZ6tiOt3TdJOM7cA9zkugGy6w+vvyDrqfljVvfeE3Pq4/ClUqGuLcv3yVu
4bAwB+vBYdvu0v5tWj0xBonpExXvz5A8NL5Pi5GyQ7gRgLF9LpsBD2O3+hxqHf6zDoxm4xI5VCSy
rIvgd9BQPYUe18jtiBuot8jQ/e61SiWLNzb4MIygWt2ej+Pgb0w3AEpTQ5b3SPdONMP7+3muvBWk
jUCDg7PralBzg81lQcNvFDTpDea9H6isGgnW0V8Xf7p94+N+DKK9c1BMdJmLaYj3UDSoYU1FUk78
ntAuaVkGA0/+AUVsY52kY+8uy9+0AaoeFzVrmp0IH35/v3Vqy2+olOxrNaXlH6p4Lt1BcBs7k9Gu
LsGfLAa78w0FG+dpyXPAZq4G/YpHULQf+gkvXRm72EFeScHRNdXoV4G3IPHLCvPIBk2mCOTmq1n8
nsZetzkDfkU/ia3m19/P395adnbBUlrMDE2ZKCyqVwp0fLiUsQWt7qmgNAy87GmGTO+K+lMfoOux
WxUXvs9oPHuDRVzYpXv2cuAbZemODImaXlJk6D++iiFDPFKvaBYpxjNoYBWTA7RDSfoKe01YvjPD
xAOdUslydSNbAVNmq0k2YK76GdJnNKCii+rOs7HSoJbf7WDMyoRqJf9Pv/E0r7D9nkhClQIXEWEL
T4TzxSQ1kalPfH/kUni4Q4xaTyL2RjSqsdGUX5+TKGO5CRmo32xwqgBoanIkNeJ2OXYMy53bGwaZ
rMcjG4aLrojI5vMCsXizMaLgaVf4n7vmWCJQY9KD7E/6J2RcQ97T9gb8PP29FDEg6nPecvy2OG9c
GDKHaFyR8FVpzAjz3RjbIogMSTuDoOekAuE8m6phkN+/jsj3EC2RfhLsqtVyoI+zQrdhAeScEu2C
rGXmrGZrCWuiVaa6rxMy9xce0ifQnj7dfaN4fDkjuTbV+qPzdoF85V3UMr/vfi2gretPJ3yFixa9
pluQM0fC1AzWbRV76wmMHXLw/xoc9ooH0TCxkfe0pF3sLbc7DRjyKCNSaK39JpZPgDOFkJO3HFnJ
y8k38x5+Y4lRudTYG7f6UNiAoEcmFc+j/BkbQWi5yE+hP2iLpvr2wp7SFS4r7NwLkAMYo5IfzQzx
NtFjY6eGExrIz6eZPxBrpfiT5BQLkRvkKGAEZavfg/8L6eCIhlhs13qGBLK/kO0AHhVgDza+S2Jw
6k6F+4PmmGOscNZ4kSXbOuiPjYEB6EdDXt5issygp28eT6SgUVIYgBKsh7K1lbkrSjuf8uPQTr7J
HB9g94MN3BZ4pm1RJCKqb1TyBMjYyOZkjxtYHN7UaLGyx9n+BHFyTpnjzw7lznVfRiK8/Paoh+xe
xsAI7VjEma1kw7szGBmEnKeYnv25ptRMW29Fn8jCI6+ZtzM9iQemsmLQKdOnAbCu0PfhzbrnZt/C
UqbrAVv7EEXbbDp/vvWGGMRoIsKOLu8SsSfyrN1ksGio1Jsj3tM6/pA3mjzgpBcJqHLLFpm+kKB1
zbMWVcMsr4F2TPJyPKYk5ealNTtMAu7IgHdR6Xe9tzwTw2hNyRqHVODDVGV2VYU8orbmDo8voTTo
dRAAd0Mj3KzfmDW1IMw3yO1TMZznjQ3jWtY5s/b9GcRCrbRWtxRnS1dxQXoQv0Ur1Npez5mJGDLN
88d0mSQiK96TYG0LXkGzmFeyRirCfEdOFwYUhun6py5sblXuerCXN7Ea4WahedNGX3V4+ykGEgoO
w8+zQNfWYub7uHwnQkK7UAzVaYRFGrVqJVo97+A7velLVG4WmMffkMd5ntV2boqJfAEGDVOxWHRn
dop5xGKPsmUm5PPvkL/rZGeOhSu53VupKYRcj3R+vKNaFCMWJ/N5FjKfMHAnsmSUWf5UV2WQkF5b
lIyd1ioYGdDwr4PZCvStrksWWkbNxDIjJkJ68VkcAJnr4trN0O0sogFPII27Hk3WL/bQhrhu8IFC
YjwIjB7F7IUz5TU0rzx0OC7uJK5k4Alx27CZW7cw3V3s0H65JFd6BIoMJOCVgHwn5SNCyTCWg1z3
lV/xlZRzYE89Jq032AVEmnBAR82RS8QSu42QPRr9+6ntcwblHJqVCrA5CDRwlvkvhqmrKsfnoot5
aBUa9v3yPeZNNqpQyMWpRA4iOoi5JJTSJWcXCW6a+gv2zScFd79HeF/+CnMHMIKgtURzj/x4n1yw
rWDThYSSj10Yh/RUjf6tl7yRxyZRD9APotcgRgXq7/PT1QN/Q5aFQJ7dIErUsaWmjyS6QRJXsfsr
JImELgO2en4aYxu4CGE7+c6/yH6b5ydvt7vn8QNdloab0ffYOvXwgip7m0ip3EMLH69/iWRpWyPM
8X36hgmgYwnVDi8TUTviB41+cZ715SBoN5alrvupq8FZ/EbgEL2abxnoMv9OPCEeBiTK7F0Eh3tT
xOWqgo2KigpTS6wILWXM34Ik/VkQSVSbXeJidpO3iesQl4H7JSweP9FcC375/w7qQFmpsi+iN9Q5
h+0tERl4AnUKBEh0ufTNXa7fx7NAnn6qeAm3uKOxc3Fob3+SIFKlSJ+06ZAoZZcqNwvY4GaSGreh
KAWw/nuZcZeXfWfeGfFan2huh5m4W75kOqvqej8CNu/VgQqDpKZ9T6wVoz4eqtzI7FAb3yPA/4QO
C4XLWAQWK6pWKghivJy14mOV/cXkWLPgmpCieh+ShvUUnJWQpGWrk9FNllzZ66Eu2Ttt+TvSzpnv
y2uBfPucLgo1GelGiQaP/HB+u2BQSZ+l857g+A9BpdAUI789NJiOav7MqIBFhASBH7W3+tW9sHNW
mTQFww8zKxmkCe/hGNTOnjtg47WjlwmFbcKtO/uOXmjYJNzkEiIdnmzbC+JbfJWs+16MSpuNYAy0
xoyGqzJGNJ5PFSg+aDhtf41U8wxQTaxj34bGY6dE2/m9gPU12mn6hsbpiXi9uPc7RKq2Pco3FQMy
WUv/U1jun94nsZ/XUmc+boDe88WUSwpaF2uN5cVs3JxcJ806Nu+eVhNOS1JHYzhKOvurplWctQVE
3H/I+LuhMS/MyCzxfKqiuH30ATO39GcSBmGO/LUcpFKDOoG8R0NY0xQxUCXEBZXaHxjoxMnreo5F
0G0PDsValE6rnC9yT6tnRP8z7nlxPV8R+UHNT3RuCT621tFetpCDBBobBQ7pRyrAvpyH65HMtwpi
TGwnQtqVLUN8JXr9JVipVSlcdyZkoyontg1y8vgjrQzsbjKhEoCUsohECqRxSyw0Dwg3WB+n3Ab3
rDEKPkR6vMu7aJ68HXADNdDyGQ8EWhKM9wT7300SCE7cHYCRBnGyUWktDqYbwW523DrUEFf8lD77
f3xZjHQrIZeDPthIl2FNrj5GwzAczbMnYj8+kUhiFeZocrQCvuPhKmhbCknaPr2K+FtM/gvGT3Xq
BtCR3anf3G1M0JMmHvQN1SDoSeUd3+6I0UIjWXEKMs7Zy7xUzknE+noF/snD9NYSAYKEeHdpCDPe
T9XNvDahjJ6UumXflS2/HKY0FzJqE9gXOIoRePGPWYS8PPjRJBId7hb+PpBpHVRpW5fPAMIdXgV3
rbwGzoqB6woZT27p6t7Rj3rx63YgPVNVslcbyQ4Ad8Mq6M0TfWo1ZP0WV7Tub9EQr6eHMahQsa/F
DZ7wJMME+ZNV96ROO4r4f12dfYRswEpfsyuUAQTQx1KkOdGZlhhE4KregdZDjp4Zj8ynaiyWCr/W
MToLggrZtpENbXT553pyaqQ1PzJCiT7kr6G6ihXcQnv0JV2z7hkH9M1er/yAE42N0tjupNK5uRRU
zxn1sw62Hx4zXh2zrz4oYXF5BS80BfQOibtvYX9qi0IQb68IEyYNjC478VoPvmjrZl4il7vYnGW8
Oq7b2V74sXk4Ve+MMa0/oWAIZlw5AOSI88O+dOA6hk/k3S60pPjJY/nGFUTCO7flaaHsxKfEefh6
RoRO500ev4Dk7WMnCHmUxEtXsjANvIrZjzRXZSEMzdfyQAEU99Z9cgCj8zuXkwV5zSIfrz9tz90M
/xYnSwkjKGmAgRMHi/VGiTMAIR/PXJJLHl+IKbwCoCW+m4z4lAYnMfPMts7YAWsPPkbRRHyyNPq3
KV5ZZGEMo6gFfnelmXlSHRoqdvDFTXf4BAvXx4X2kK1xCYi8YLDLQ0edUXsokqay9rbERDFHMaGq
Bvreh9LfIyqoADPDEQ98MDs43SYs/0k0B2/vKeFpRD01PcwnXPlKlsbW2lKLwrJBJZ9pLJ1tgWUW
zfIrdKFX/ap3hWVxixAiD5AMTkbxTsOSD6BRCA3GnYuusWeHSDnoH/qx2Q9jRcaBqWel/BA5tjql
Oc9KZzYmL36a2v0IcfICA+GNpxptZgFjgoiW4oCt4VFS2Z4sYL7dJ19LZj6FBctTZgrj2ZvAPWGy
lGQM8cZL6zdmzljtKuISFiS4MTl0WT4SiMMjXOWmZPmLubE5WgEfmmbrT237mCFChpPLzcIU1gOF
YXn30AcOj6p/GnTq+xKKAQbKt0sD8X1dI/HainmOlrGjSNp7wGnLuToG7dQGix67t36tRZd+Ie0m
JBpWGuXCQBhz+dFj2Df2CI3QSUF3ZwGNQ+wV6MKy8WmpGp2a+pQLUWoyIJP+wB4u6RQ/y0VO5LTb
9XlPCg1CMFh2HIzyvgXune6P0Jq34Ol97SaouSzGNUsLF0/NRkKHrkaTKvLKfWmELFAQO/RGQ80D
VxST0lKVLcLTQxNgzBKxlvP5lS8hqRGpSfk48ZxAEPVTb+iCtiXPnF7q8rcAErmIowlWrHLEwd2w
DRGryOwGYSkbqtNz0y5X5FjTE/3UgBCXSM26AuAYoXfkGlBBY1BYMqXsojbh93udwk8HKEd9bAfF
LW54BYVaju8764V08AAhiDUo6nrrtixx8um1d/AsFRtIvJmUKTAqkhxAxngCplOU5zNO9X2o0ych
XybSdnzuY9PC70u/BFmjhbumG502FrucxXQy9nw1tk2OCHnwRmooMU2gS6bON5ExC9Wp/MDrh2d5
cKSuLMQJSxrdlP5auNKyBF0Jv6j7IhAXCc7eDzIzjYsrp6mpMLv6O9Pc8M7rBj1ffTurP8LLQM0L
kstLIuAkRp+1lb9dEN3eeiu0M2i9GZuYgMIliSQytHY5ahtH1aXGfVWo80+I3FEFMtcbE7BJu7Aq
GFw01GUbnrfyqaxJ1EfwrpP0+I4HE+GJDXHNF+PebgJSugu87WTrexvp+BKAIEv2tzVmrQZASAoi
kKdtzEvHFjbil8482gy4gLAWVSlPkqfHz2sPEBLcacASoR/t7V7IS0OD22wOaoeqTEZQUaC3Vxhb
jh/WuyhiY0Q/G6SKTPaF+OBTVmNHSA/rHO97uq1AXTXMePQNF5OM8U1iVYGS/AQus89AYQe+Vter
0jIV4yDyVKbVft0z8txe7rt3mbTRoguMfGy2U+VsGUVbH2h2WYUyOsGlNTFsSTYPAFGoSGT/WFs6
WX6xvc2FESZSSw7IA5yLRUTueTQ/WMQZJPcMKr9w+nTx8rRsI6wOF4cD/GQM2KfDbr1qxPVYua3P
GKFTPcOWHNzSbSCxiqT6zTUh8Tgn6O6VH6YqQJFsVLxkefvJbib8DUfeyqZ7VfayALdpXW1CnLvG
uJD55pl0Sc5Fmw789ri5kkeQrCeJksCkABS22cnIyVZwmeLMu9BG1v4DEGlEPStF/OWc+zKCiM4q
j9yJAkNEui/s7Ix2vzAheH+gOeJeRHnXPPwS+wzYxNRpgj5Cs2Lr/6zeX1ekc2/S9YBS99M/rv4k
h89RBwaIP2q/TU1MaRiciwWvzCOpI588AqS5czZe5Hj3gpxfV3XD0NzsMj3WosrtY1xnjEgYEWRi
zceJh7mOkCo5rCLj74Sycisx3eDq58Ar6hTgZFv5GItpyXDUle/YYsnbrcfxdAxUM4YPnRQCZL45
nh6k3bpPPACiMKO77NaTFWJ3YV4YQgFlz/fLD8IdYn/2bxdEBinaKNIOW7RIwzGfSqqxLpjv3sGQ
QiD1CHX0G58/SNdrxq1vXq03xZb18OrNpIb6JjCBXuQmJhOA6wwWFsPGkjlsWLpqW7KzFzXtl12h
faIyXi/TehLJwqwx+5GbghF/wpZQxJxF/xVeLsTm4oykyrMaY6+YuaaVpwD4TwCirPiDqifSmXcO
V7WIf1wcMwFw2a8yEJaF+N1lXeU0JnLKJ6hvpUkBp1ri4Dq437/l21wsDVxvbWyAUanbvN5RmeVZ
j7vB0W88b6Pl7LmlH6v69KN+cHSCDg4z4gGjnCztUfJYzaH4cP+86ZxQ87e5U4k96xOaFim+liT6
lZ1FqXqDYlqCVu5JIg8pqbgcgDxrOGnqCDOzQ6PhipFXtWfdK2HzjzPP7FcBsAAUNmXTq7MexMB9
Yymr5rUKaA5jBn1Alf9VxIl6A5LWNILqer1eFccpvxxz1NadZaMAg+pslyrBAqRLq8/qz60auj3d
elyI7lXDH9wNv16A/tOyOet0XSLvWUBfQnxWPdpwPfvplWsmluyUkZK9exUHuNWE24cKNv+Qcef+
eQK08ebbv6WIPsQ0F6Az5ptXheL62Lb3l6vvbo0zGadZHcCRQuwj4XKT+HqJrINJTDSvRunwxajH
MUvUy0DjNtXDY/m0Y9V6/R2ncr6hiTL5KhcOvuhCzIkmBWUhVOSxXwvdYOaujAOlvjxkU4vPdU/U
yJtCCrvhBAyvi2OOVuOrk6vgq+4L8xYkbUigAruWzGKq8oUkuFP/FYVpHk+eNmIrjTiaXlgbcfC+
UOui3161GSXBZEkPWuEqBS1SlpwK5QbVfq3KR5jN0ccj0tTRd5O0GvNICQJnMhgrY+EGH8nCkn5n
FNXudBLy5Bn8ly3Mm/6BBCPQkuN1crKz1ObDFYClSlhUz1dQfeEEUuHJt0P0ITr+Aja+McofwESk
eWXbuEOidaG1xeblHZ9790UKlg6hk1tUpHYRdsqg5ezWcPgugmcPaBCnt+Y/ZxAz+4NW4jANKUAK
Um1qOaU5eNIcXYzNWb9SByjcJPZi6I3xx6mfYAGtT2AgdE7tVofr74XLqHrJ7DOTdms/yKum3JeO
NNhzY2b8EC6T3Yc0kbiIFNssh/VTFeSuNuk3T/heO+A6MgMbFi06oI6lGaAwoUJo4jJh2diQQS24
fMhe/WZ43tzwM/oSBvDel78cWYMTf9YnLOSe6Jyfs7m0h8dW64K1fcUFtLgmTmwY7pIxAhSYqEIX
K28soVK17Gm15qESWtzfwtJ2Fp/K3TGFj2ZqsAkZPABKAXE7yIincGdrwAkesZzRGIYpDMmrgxJ4
eI/w7YS8w8/OxF1QBOEcATnFZ3QN9DXLoEs7X9zknCVW5YvYepnbdUratNPJAWd8MQpHgsKrj/ut
hzrW37V2rohg+iVqm/wZq/Db5tylLpXJku6sDDBedZeTIDDVWh2NLdirBHyfvr9IWjh3QY64agwu
MJPzqLKxEowzmhhKZmuVgTjjeswbvWyfdZrP8NbsUw51dEofuUElZ5xBNhRNJV2625gisjBRET9c
C/OOt510MzXsaRlOFZkxOi/kSE9bIRXB8cakVqrWulHhcLyPKqILHfpCVX6QJu6vkASrk8qJvcHX
TTURb6teDiUFUSqpMnDM7xkmt7rQvUAoBtkLtrDsjhXMqZeUkLWYfiZpBopOIZt6WD0bkeYMxMOA
WZDdYw1FrZfJW6IAGqqTDojQg/hIeBZVSsiyd3tZqgEV3WI8G0tfQHwHzbZSZUQuOdieEh1yqqox
rRsv8zsQxd4Tr2CoBAZ2BxNKpiCVcTh+127f9s1z7VGbrHCmDGQat9ouAgXffYVHHdbV/OBTpr1I
i93drXDFue8XQAVUebCLsMOamdLzYBRcpGiRu5Fg2hyZT1zK9x2+S75R+kj1SHrEj7mfFhKmIbls
nOnVpx5oQMb0Tld/FhC89H46hP3NncBKbaJA/RezdoD5iNfXAKMEACL0DrlWKycZEHAQH/i8Yu44
ZY/crr3AKNHn1n9HOrcG8eZBctnW+q9miee0U8Znblu5DzcyRBYvV00uLb6vZjxE7PaUQVLwpkuW
qgXWGoWBkYLaxvCCDdPd8r1m4AaURuu1ASfYgW6BYPh697AFDdyayatQyFBbg6Sjn0kCfOjdKCST
Ks4gH8xamx9D2ezr4IE331nY2xMdmBJHI5Pt2o2XajoWQbsvB6/ENOSoBbE+BZMAMtFaPN+Yh4vA
q4HZkk6AmrZH+KRl8DNZSC7GUCl2pAQskBpexm0nxFJ8Wytyjm0RPIGelzVR52xCy8rV8WkSn+MC
EeF027BYwJCEGGqqFzGATo1gNfFNXVmSktw3GEtOQX26ioyzZBpTOgNGIuzxVT7imzCq6vFdtydx
vupA4u77h+eHA0/AjtlEwdrS79eGCHS3bmZlwSem0/xcilzYCtD9sJaNN9ZWO05QNJKHlIvTZ4wL
DIbrDvRYvvvumq604xLWTnarlYN2t87zhIfuXuTMGCZnrR2wN8W85qC9Lz6MF+9yw0Bqen13F1E0
wxOKx5kNAP4uL8SO2Xx+oXseSApMBKvrZkNHLWgZIasYQ5Z9Yedugb76EH9Fk1SmWQfFQXgIGbXo
LMORpsndX+zGiX5afNsuOPdzVz7Hq8tP9cYAdBEwCJ3MD7/pmi2XJGEQDwXPH+DSFZPC17ADe5xC
oS46iKwJbL/3uNbpDKNj88//pqpXvYociw8QV3f6lRd9Re1ue377BT1fpNbAzRL+PV75KWGp998Q
wuDaNGxZtzQVc+gxmAsMUxXsdpP8j4O5Ol9OJLhBK8/+mkH/WinGBV9RCy8aEkb8vPn8IkuZwnum
oPbBBoP+BT+53dKkLFmmh9BPeDTYwwvIYJKC2cWm1UPykDd70vTCPoZSSmZYYifsmxRK+7s3VAry
8uEhilWMfMh176WsQbNJM8bGM/V+Lxwn+iQI7oNWB823+m3HiansYkQhXmF6tHBtzcjePAC9hwNs
7f0XERlv/E7V7M0pQ7un5tNKz5K5iXDrKd5xU/uU/NvSf3N3R5a5IEVyZow+dx/sIW7VFPusSHoJ
KJVrz5tLM1hh4V66/PevaXgqi7TD/IUGnCkGc18QhZK+YouGGOQndOVtD56z6emJGWfMogqK2APu
SWSUk/z91iSIeWe8GrM/L2scbiXSk/BodN9/Nvj8tMWOGAQ3qCixd0KXi5h2LNkFRXzJHmjmbEy7
27dDpkDuOei/DnANGYPSC9LGTTeO3zaLqFqieV8YY3cLjBkjUbRAt0bYDYMcxNOUVoQDV6UNHiAh
wz25HTJBq9dPA5WUOc73A1eQ8QXfpqCq56fYuUsXJ0FGuaaPkNJ5WM3zBWdLbsx/SKd83srsmPS5
+Q0Icxd2VUNaAT7H61zpmj8K+FaIM5RmmQrd+u1zGCFlvKNOxiOnBBaBqkmxpEHhbxbPAYI2vsKj
XosNWz9juHemC2xhxHfQDpq83keD5oBeHsABErFEkfW+UhfUIuS7DYmqTqisLWypkaqAB6+CDjLq
an6N0Yr2RT2d+oZaX8Kg14oSy7+mLKbl36Gj1vT5ikGLTHpPrvSJmk7Ac7NOoKkc8FmBzTd+7NRx
xZSrEdnnShv4LOzTvV15ooHshA6EH0PIc0NoDrSRwIuIHz2OMan2P8ZsWoC6IsPFASXH8O+Goqsg
+yYtRzvL9yx7mBQfbFs/VhkEPQaTk3Vfn5esCttoDjWJFU0NM9/vb1sOYgNYzpjlDf0Hh3uJp90u
TwLr+zjoi7mHsoNFDx1d86ur3OO7zh/wWwlBfaXuS4rWJNi+6Ml4pgQRgQ3SL5sGFry8tzcJi4BC
hGdfSJ+Iwnmg/FqGmQYN5FMMiqQXH3QpiN5Ar3ZUMIAkK30dpIc2Cl760nz9wMksv+OGikKoYOWv
GJ9R+CiA2U24nk56JSMI5dS1ofHJXO67PFxqMa47FqOAdX4O84ku7+nnI2FIQnROXx3fZMMcP69t
5URRvgvMb7tS0uM689CpMpljMxQ9doojF2nZjP7ZuEYIP7YdR6isfPp4Qoa2DCe2cj9p+JSH4aGW
NUpoOaJ2rBm/Wfu4D3BnuLPtw4LM9Z0MESy856jWWwYtxakWRHjTIoiIvkJ58V5kkxaXOwn0/nuj
G0kGmpjTsm/HjEHSURtMX+Vo8AT4AE2dRdMemZC6D+LMdtCUEyp42NcIGkzlSVrMlUJ64GfEIWkC
LMdPDkcwplu2Kkc4BQ9GwjmbW2kZi7gLzoKUYx9OQeyc7DkkYtB6i0QVszLkT2XEA6pzEL8fXGUh
OXE02f941mGzcloUF6mcr3UF1xfq1ELkwKVAP3Pk1zJ30jQN2C4L9+nm7WilozMe2jNu5COKhfBc
14U46G6Zfra7UlcrPSxivI8RLUmId/63DCjcaaFY/QpqM+59TcewNXt8ZO9XgCA0dLK4XFlNjx8D
Qi9nyZ3czyNVuFJRlpLyhnXLkCjT3ts47TcE82/8DcMF6mCfkAqNi1qqHRBMjzM4fRksnEwyRrwC
aScMi6b5YTCbDKbj948k+3slj1K6rJJrgjRUFv9pITqbjNomotQQTKvAaEvQPN1mOSKAFWSM+YfN
8wzocgaiZ3/YLk7gTWZx2Llstxsgg9a/V9UPKTDVkEOqyEQkNLpUpRWgY4DFJK137BCH/1japrdK
YLpd89wX8CvsUopwr/h4DK+b/o+rs7I58YB9G2YPTIMjUI4EGwcFVztv1oTpZyqS0lfi85g/fVFx
bhkaI8EXvm2lQW0K3NdxPvquw9iHHRo8EhtG0fKcv6bSh0LOHM0sWVibvqAfvHsUwGSgSGcnk3Vz
uBHrF5ZoxNP+t6S2PP1jhuUySqHL/VFfwVaQziy0Y7FKjXfTnWMUegnZkXV4GTcJZir8KqrMczzZ
PAUQr7lha+hcNpnoMyUm3ac/qmu8bZOCkb0lG9ngWyu8ksH68dJ7t4xfUz7lc4eNZYSLgGq73Hew
L0O6UbRuOTbNVgRHs7sdmvz+ZUJq7Ss7XYapMoq0/kjgUGpJs/G2hI142ynHkD6cNtC3Jlx4hZLk
j9CqgL379QCIduFHd6qymdPBnxnLBwjwr+4n3KC6KSq/bj10K3a4Y40iHMi5TuB6Et6NLuBAoERD
7E4okNByS2HSzhkQeBrmW3PMQT1lsbt2bdc6PaPqsA6dy+/IRCxiwy5FpDRHOS9OWXtbET3Eye0Z
Ra5T1+I4DNMpJ6/M4ldC8prMY3oRO4YxiYoHZltxgSkDZDISgjgxClSY6HvXtnSyKOUbry40QTb3
mjXYzObPLiJt8fOgMs87ZDiHOtWMpuyDqzg3WdXLbO6ldq/pKqgwN1YHvrQlc5XgDcGCkdiWwu35
6o7pZmMIjYeUqUsPoCEvTHsLJsKWYP0YkHxrd0eRU6+lM22NygWg1cf3OaOtkEnocTyt4Rxw6Du+
9EpR59tLPchRZQiGOJqUa1jpDgqwI/T2QZNlJsI2X7bFvWl7zaNBUNRyixgwMb1kA4behwLxkd+k
5UijRCfVhP/oTqOFtHDzhAYebtnfYC/5VeaPprqNvm8G07XA/3iU1gIYFQ4I7gekyt45dZH+StUV
KcqqN2rYENeHdhZaLU3ZcuhDSAP80eml3t+mqOdW4Zy9g1BogbudECWNW3Dp4YSg6ZQZ4dyqiK7o
UyyIfbRP9lHra5AtN2k2BkFHOKugjjEGQvoW+7HipTOKEUgIyFPkL2npGPhWmjlK7T3WPf8FIhj+
jAug/JQd8n6N/ZLX13AQTT8B1Z9G0iPixvYazaoxcBqtY17xKlf4G/lppwYTsIyqeiwdY+g4Ys17
DroO83RssfNEOOJNZcELu6ZSB3dGGk5pejAebhdqB/0DnnNZWUCFI/3W6EvN1/tkP/1w5LmBobJ7
FxJm3D4t2X1yWMuniI7UOAhH8I0S6/zfOV6iiLulWlu/ITDgR7+Q9dtP2VSR9ZDeCAtk4nEXAzds
zb/Vqyuf+lPcVQn0bWbSS+kD7Ymc72J5LSttn+8eAm9jvYuatdw1kalXrNFtf+kWfuovp/QYyYAz
/UPj5+cXCWoUc4m9+3bPdzcJ3bPCV61oxhJrIaAOg/oNnK4UUvIOmgX84TCgWCXYC8nyOyduG+kp
UYWxW9912fBJ1XB69mX6Ur5Of9Bm367k6nij760SYqw3LYA4LSarZzoVoO0oSVa2oReW73ogwU+/
DCTdBmFH74r3BRvlZ0V+wTODVxw6wyWACfVl8NfI7STxi7nnMpHnZcm0uhoxQoRAD8HXhj+Du92w
E35wkZqpjIPFyR6SRBmCG6yx20i0qYMiWDbkWSmUGaRFiK+3LpsBV0NbCIozVFFl1ho9K5TIbwrh
1F6eemUIon6fhaCB5YllOXGcifgwtZKiSuCJQr/87f0CzXR58olWqeAFzWTTecgn/CwwkNYF09rm
rbjWAck+F0vBuc9XkpZWNrox1nrdeUWiSMQwt0S/4mYTmv51OE3t2IGF14d/26K5NigO9JDpXWmn
wZb0YrlP+Y5xA7rABXqCISd0uWq1p9nV79lgekJjUN+mowc6z03xiuADolEQ+lC7ggVKJmLoaWSA
UxT6dIsIm80k1zPpsV12HX6BD9HkwVFmtNGVK8TvIbjat+aYhkWHZiRQamD+bSFEaSIuhaQaJ3SF
Rryg5PDllrzic7RLctOBUKL1JnMUlkNnhN0YREKnZFusGN87QolQJlKm1JTvNRYeBQ9thSLkU6Wx
nuPnYuz1s9jco1x4ptdy44JYjV+cVJr2pPn5lOTZxNir4Mucu9cwf945S5eYUaciv8hFalU4IQJK
2aEUzsftPRXSpvB0Cy0a1zVkO+hhRMsNYppkpkUCsshZ4GoikOPalSrZzq/tTcZh1jlAO2jYMtVp
6VFaEuBAXE5+Y/Pn8hUgl5LyevVG2CF7OZ5jo3YUi8sAYUYQvX6HUK8wcKd2k7qrd6qQV9YkP/na
xz3tB6Bod5kVt7wCuNx4fk3LoEHVwcs4Cw1zmLdhT7p128+6WsXBMJPKnk8rQnxil60KaSkjV/t/
QOyrDx1VJaS+e47AcreXmPaOR1OZ1IbBlDpy8hXG+Tg91UcTU0JgOQSFswqpPeASv5bblTxSEMJ4
y7VkP5r7S+5tfbocM92wgyl1ocJCHVKE1YaQSNsKND32/7I56ZH9e7xuYQtmce9TZQtFUB+mFd+q
cNfCJY1oNiZgIr3Bntfxi7zRHUl/U6ZU7wht/e+K+lwPZJHYveLoRPeLEI8IeBLOVLsDGmx8Vukg
Cseqf01ezK0SAhjBxKM9+dp23j3bzmBEkZVxzCxsMbb+AoR7R01Wu0GNKdzWZrABJGlJZqJpxxkT
KolpCJUpC3kmbb62SGmmglqSJ4EagkJLHCDMOo9YMhVzbkBHTX76cxnvU4sSGwFtpFrdOTEirm9i
msfOVnfsODjtjdUa2J2PhM0gIA8Zbputja8rI8gFPIuwgB/X+Y+ACAy9XrpRHIREzxetyHvA6sh5
Mq95IrVHH+WVBB0Um5NxjCWccxtVPIcrKi9V8B+O99oHjZs5IMtI0pEJPBFmy9GphW4w4t0DgtD2
uVNVN6ztgKPgRnAJDvcAaAj2j/fF9IURzk5NgFuoV4i5vpT1K8VavrrkPnpgkkP5aRbVCTAwWdYO
18oS6/TGy8avqS3Vw9EBV3UIbQOadXtsF3aIMfPbugeu5dxuS2iyvZ7u8Ny6/f5RUpsHy0qPV4ud
lLxg/0NHRNQvRuklz3mWGbjvgEAay5BCti49+MTWn/TzPR4Bl+hirPlB3KHdkjOFrkamcHQ4JT1a
IuCeD9LombDyBQNDQDUJyd1USKGE6bMDUgOeUgrj+ZaVXPrV7QG48mtK1XhCBrzgURUQgk/qOhr3
huL0vnUaDtgqQmGjgNtyD6xnhHFhxjQlhCW64QDxRCiB5lMM38fvuuawyCjqVsANgujaIB89fr5d
bZruGPfzCQK5F6xMNM+MQq5n5MnXwCCUoiJXbdvYOGpqT+vy8iEaDP6YRm+uQlMq9HcHHHY6RsHJ
6fBw7eFr7sF9PYZG9pj6+YhLj+WOVtgF8djszoFPEHmvae9bnTT5RQipd0d/nE8dc1swXdakZfl/
40sFLK5N136OaoMJTMYTEheQccDYoFe+IH3kpyTWpCNrLELd7AofyHTF30h05AmBVpMr0K8aj3SC
cDcfPJZZonTdbNomqlbNRhYPuwOCg4DpnUcicuY+GfepkCU4ndCg8m3gfa47Eaw3ZzaPR2Izx4rm
d2rXlM4iDVmGzM+nWH7E9LFZ6PWog94RM5/nrJFhndaQBnT9y4LOwKD+yfJ92eoVr8QgRUnB0fTC
8kMHVjjcx7pcTsRX59Q4UmD/2lt+pYRN9DUTXTC0XW8lnt+nkFj4fWeIrdAmEOPBKfPHO0a1aTaD
6I3FAgW9AJ1IccAe0FOx07HRC7zsR6N86cjbIIuVY7EdPHOmpfzs52z395S8mc4Un/ZTReeoarva
bTgUN3huKoK9IAfE0gOUPQ/A3K6ODVQqZIkS6ZqHIlzIXc9uWaQ/LVyJd8FOM3KzW9ZUZ4H6SeCL
4R3ynC83bRg99ZiNTI03RhAWbk5PykYNocCqSMqB/PQvjN+W9CzAYsgnSgMGSp2dXyMXOUVpM7LO
+fWOIdK6PYuV/WrL+nztKz7F9jdei/+Sh8CWOlT7ND7WKQkIDvyutZErXJroxamxmvttBh2sI8tQ
ZS21Ujua3to4KRNh+3l03OYj+doy7XCsZbXdAvFrdeFpTEgRCPhTc/QIZxAN3HxNr8XANDBMkLd/
d3ukfLy7Tf11HmINl1pvt1lni/Hn6FTy0noLxfz+BGVbtJxO9mNN8vWRXtlD9r8e8jHs54EESrR/
wx/nJ5Y+KZSTUPW1DsVFvrql+w779GnHQkVqF3a5KTVdOANvwRmGB0rRNm/Px5B0+7nKu1C0HLK1
VC7Z2QJECLuwtyUjl0EKEVmcftG89iqktr4faCwKipDpuYD1Yd5VyglR2x7G0n2J7QsW8xY8xBQh
HZIxPV15KvoKQY5cipdttBf5Xs1QIMh3fULSOQLX2l4ErvCC9s9NDv1WdJ63M5lRVuC6qk2iqzV5
A/ZDTEGIdTdaCkovvFNaQpWgE2z2IJOjcx6WNJJqoVaf1sHq7EuJjT1kzsQV9V3BXCATfEDnf0RN
sy1kUikN15i8r8dVBaM3GmCIvk6dA1/1W+NvvTDmbH8hpqXUlvlE59xXL62Zad8rT6ViFMeo/qcP
allAoSpZJIOYKHPwUZkmeHTLLw12GCbE8z2+O73jkCrTt4kwJaTS2FYBwBeriP3S3pNIuIz38F6s
f2lXOGYE/wCFFw78i8etVWLLb2F2Ztj7IaJdfVqxvxqPhAkCs2KfCKomK68Ev658UPzgqNoJmKXY
LnBwTEgEsSEjmD9TOdz9OIIfWSkUo1wNX1DtVlDrtfzQLCwYSNdx3zAYyPN5wcUjw+yTV4ZOXyyT
9FZ38miJ5PNNOUiBZJAmFX6tCFiKm7B6kdZHSuS7mtaOc8RwKheoChUMFfFGrH36H8NBEEbC9mW/
TlOYVrV29V6j5G8H9yx4Nh0pveuF4Xh3mvGW2N7P6Inbist+VNCgE9DviEHujJbK8NEG1JIG+rCS
QZcenqfonk11X1IXPpyCx+z8CYDAI9X2tkNrjJVl2FMAquDaBjbHXgLQDT08JtcH9fsqg6VkuLg2
5Xsy4cJnHP8uEut3IMO7f6cyWZM1IZhwBl1coBLp4yIohR87avAdIr1HBMIH2AawK1CQ6XnFMiTx
wyKzsdrVoytNPZdWNRbT427EBx8p3PdfMUmQub0c46IiShsaDndG2xRUOfaPO8MBxSXO1SRwFpRC
o2fwtKrmV8UQFFSu/3MYDmgjqWHMKQ2i3JHo4w9y9UlCuk6xX/6TG1lRp5iq9YTlvVOqAazV3bs5
g2Hn0t/ASLPFj0qTv5BcW0vs8Ky8RyoPnV08+Mq8MMUuwlB62waxpXt5EXl6zapDJyimG4WL67Qn
4KIRlnXj3qQ12YwONMerkuVMmPpnHWOvdOuMjpmWGLQQCoMxu+g6mZ9DXNofi3pUJgUTaxgrClEY
V2RWyVBxWqGXfjYn3w32UpPXeBDJGtDzcFoFXQcsYy1Zvap9xKU7iScvcPyitPZRLXf2qu2pLdy+
e5verJDl4J8x9PPBax8eaQ0nTtfGn3Fay4t+4/ItpOdKS3IMc+tSX9QLb7d1uXezCq7RNVglHGpM
ISTKfqgiqc7qIuuZ4HkYjtM6aJNHf5PDGu+Dov6CVPMAeYHXhK/ieCuFzcX+DVLt+hkaph3YMSz4
qCWvonX0QwSWl4hywtZMPX+1KA8P81o6lSGrW/cICIvOyWagmoyk6imKWt3tSZLtovgKG/NW3QxA
FaRZDslwj8rQ5bD1Vpvqa3dQER9fkmxB4PlN2Z5/+BQ5hfAoCmtyN7wha2GoRaSnf8r2IJvmS3rj
UJm4NO+Spt/JVqIxoJMJhvUej4clGV0v+EY2iH2Zi2Od6E38ir3BbNA4h2u0NgGy2VLxdxEPByV9
xqg3QakgbZctldZe1hlWRFkGnB66ldd59h+OK53mLVGWI7lwK4ThQGCYcH4L0+5eL+aaVDMALSoL
kzYxNRBBrzA/x8UnyTpJrMMIrEahKT0dDtg5Jzo9b5zzUox3UzyatYSR+NLn4bTz9FalGX+XsS/C
YdRHa3hD4chbPdoJbW4yCwQOnL7gse/PVVmB4xv3ZsQT+Al5zhDUaISTxFrDvv/5YTLWcoPFMoz9
UQBZmL9RyYcVNYeNDaywvqjDJDPIr5DwLOp0uiBMr9ak01xKosmkYODnA71CICAosF16MSVMsn6Q
myHu30QIuZoFIaDU83gxMz2lMu45truUpqPfp8SE+pHP6ylHUj7u91xIBRa3P9E4D1i5vl1SZLzy
RT8t9bWuibOUHv6rtmx9VZTu6R0fgXgzAoso7fpyuGRJnCeW0uvWfMk7PlVCa1L5OttsDQg5TJF+
9mLEVhaiBrdBNFMyP9x9xcbXuW2vvtfnF2reC8rRmrVAnvZ/5Keki1qhAKh+RBK+K3qEuyj6GXjM
sgzd+Wc7JyTU51f2ye2MZIpyYPA/STIFETqfcWY16rFBh8wm3Wr91f5n7VREYzuxoIZgAQxHjuam
QdWR5M/srPRoC2Ypz4g/ximF7BMleWHtPkAgGWXiQK3PdaXYXUMXQ2UJH3odybYMb7mVMAuRajVW
IJ6TjwsNu5OQOvYt04o9uQyTndwMxKoxuM+H3NWSude612pNy0ruZMxdDWy+yckf2nG9nrbuqdnx
LhmhNMyB2NggGueLAvTVJDvbuPtpyslvpI53XneDmMDc696+xmrvFTtuwLk7qZ1kJSx7Ha41HkRZ
f83F99xn5687NYGD9HORYYeSS0UOQuDaMngMLJYFA/5WbgSREqsXwBlnoW66VkcdVwqzuwhYW5G1
hp3ts+F9zotaikWiduT+iX632XLAfkJ+IC2k/ZG56UNyaud1a0+HcAg1qJVfkDeBm4k2bIjjEUdh
J0VLs/K6Z1AwSQcUDNK9YxT6VsJyhwkOcxUXcLwIpdY66NZEXJR2x0R3hQnO+YETCOFKFDXsZYEz
xpwEKB7FEvQYVeLoNFHCT/Pj+2PNwpdzq1uzrn6DZor1okc91sS8Ozh6wClyHkZMhd5cEnHYp27S
G+pqy0FTalAXIN7lZlw2id9uKdMLPmgZyhwIIU4Hw3zXXR33BP42eoFAtaWNU+7in889lWjl55iA
62LuwAxV1A212CqFg46Dw9q6DyoCfS1c6NF4orm5t9JY9Jix7xAw2Fw4Bs0QIodcxfNtnYdm2Jqo
VQ90rEFdtBuIZHWlL+aIk5jOvCignkoID61Q9QkwQMTY4OoKOTIYE3Bu+f0s3vG5EXEcIpgR76D/
nsKwk5ohDxVG6f/U2ZQNYI/4rvVwb8UsZFpYefcyXU/+Yptrup1tpl0E9qFrMjG6AIvdaGUe2MdB
o7V7+OPfxbwlIyb0/2+ngDr0sWbohGey+Dn2R4XUCzbhcl18RCITHPh0e1Joz+DMlzQNgLg8Ltpl
ObdY0ZrTNJ7BhyWXapDNWx7rbIVUNj3XPJgXetJOLIx7i6NV3beGLpCMyLYf4Gqu4RjnvaSisiJH
CYghfKf+TnhoJINjNjv5y/3pivM2sMriMEDOSLBxvnUvxuZIJF59sZS0ZAeQIDIIGCSIae59t84F
ZmCW5qh9v6GeT6iTiBJc48bU4Dkuyx732FnO+zN23QqmcK+j8sA2vFAu11PGhzL9zIG1Cg/nOMuu
vOcJxON1fCa9j8Sb5v8+8HC8Ugn74JURbCNDemZ+2j05gh/qJegIFhnmF3aUVkqEikPu4bL+AMhK
+6/hFXw6vUjGz0+RfcLFpeI18szARjpLYuiYXi/U9/WG7w0otdleKf2QwGTROQwCXASIZ1/bRQkZ
scRcqlIQY1BmKc9AMnwO5okonerFj9zIEQwpPOFWMN0Zs0e8lz5DgMHnmuaLywzHbgCZWC7F4yo/
Qz02msY6U0DAJTR0XiZKKY6z37ZZcHLWARpdTIPAWZcyim7R3BnjYwNExFHEKFb3/lFYg3LxTkR1
Kjw0mB/kszQDZBobDlvPab3On92KhPoSxGU9WVpTryYA3Xb9aKjgdyvYyi2EvdGv8MMlCedk1QI4
rpClVUCItCuSjlHqdZZzm8ADgPTsv8BBCOKDfTpZf0hUde/PTRwJa9wliVbyyQPx2a2D0vPpaqp0
3S8ReR5rOh6HEjz+ACOUodMQXvh2v1Tg7PLwafVJgK7BHId49YHabNPHwIKmKLtA+VmuaaJv/z20
vRfGLEI083kABTg4OFWm2eK41nT8rqhUKeh1IeQ5IpGun2cToIcrqVrdgaEwqE+7nf1EM3BRFIvp
YhuEJuAomp4O9BFmy836EOx7RAtzxnjwJy8a8A6CxGf4b/QcqEAu0sxXW42lLbleJ6mngQSgDlh9
kFf2t0fA9Fh8Mxd/Cfcq9KMNKkcAIGKnS9ilgacTGKidVyMrDvrWhFryhLP4e8JxmOTTFG13EdxO
GFaIbfBaVZd8DssZDYmU+41uaIe1z3qDELayfr3ZUbSTE+VWKFomcMBoUa79VEk3kv+22ySqc3+a
MOcdaO25OPv2JcY2iLPqqGUUL0w8SqzquhRezU71dGQzJuyia162wENH7uXPHP2jL9LJRezOXnBq
lCG/LZ6z3lXI1AyT7V8jl17MYLmUU5q7N5ued6Psyil7YUh2GPWtTbvPcj2qkPnWA9gr7KT/N+hE
mud8Vktebh10bVKod4+3EH1i7EufuMbYpxsUtue1dipr+WKi0DeVtGsj88SyVaJQRNSJ4rGmyrED
T+UCoaU94pr5eZhdorPgCMsAg25e+teqlgh/CJYkJej/FaqmVitLCUCFHBXuCfAw3Ms7jbyFaAZw
CpSC+dl+sHWVL9D0P/8lcac0tgMNtSs7u/s0q3OhnfFysaAqK2YBb+vb4KrNv9czvRbTx26VczlL
VDr/StoomjQHD+M6VVpHJugbmgLoCrop2y/H8a0ZCaTylGxIYXEhSLtO7GGBzaUYioFcdUv7S3gH
t/TSspT2oQ1UnWLAgwcvD/AHfvCTUAKc+rfA9YGpXCfGvrNQ+7NVKTMMNIlTwX1kGbEmW6s4Xc3S
5GESpZU7jlh67yCkqznKWI9pM7WWew9YvwVPAnaBxvTYFpqHAQyvqgzXh+HjuhXj5tanSD/Cbf/Q
hqj992T6lBo/5SpplN99jbxUAYMdur3hCHu/qbLS4HgeRH9tJsQQ+qrQ8mrx1RE55KK4Lvi0WOnF
Oeg1URZwLPh37cBdmxq2Vb9WwHxKHEz7VtsdgJbv4erYol2o8aPqVQn+2FW4AiDtAyyt+I4TTk7D
+5ZUpp8BPTcZ57l64FsXsFoOu1FsfBK0hCv3ieB2qShwL20EYky161y8GE8/5ppSofEY8P8o7cT5
5IM66yfeNWR/H3R6iyrVG28fOOM0tmAIdzO7aXoIBtDGnBomY4f1jBzU/ovsvavj7NscKwZjvAbJ
5GwXZyJG64vKa83Cj6iMvuUtRE9rui8gcEeWk1JA3MfZcZ9E37MBrjylU87O/7Ofmqkq+ofFuCd0
r+h+8k0GgNBlAZBGv/hrV9C3Z2YeqNpqgv6UlgUCTZwC3fzJDFwnsY3Jgt2ZSZ+TUf9iDbEP0RVg
4CN+Q8JlkWepeBcMEnjPijgv2zJ1Y3UHvEYgnKGRrriQ0JM8ggw4CzQLHlsB0+WPl/LQ+6sNTE/f
ZS56aK/JyMT377zz00wK90TOFcURewLaHuBEw/sPGyC4U0yXlfl9olQ9psBZ9f4KaYLkjy1qfDPG
JSg7XR2qd1fpD31ZNLSRV78FElNo/Yl7HnyWiJokFNtsWQMglfkF/Yv/pA07tg1xElERP5nJeMg5
mO7YlX2YD/CkPsmGqMyI4OYuEM3L1HmDtEz82ObA14Ba18EtkEUhPU7Jgxr/gpBqDFmUH3RfQIYn
fjl/ZTJYD3H14zxxrXyaFvit4L0s39X649OT6ryAd1Wh+UR1Alzfpx/Bd4ArTSgJWrR6jOcGx6Jp
MYIlFZWkrhWyLFYqdjnq9BskDD2N0ZYyrUxTWOQLpaCsccaboJnH2cTU+uxsiOGxvhATr3Awc2Dm
aMckRMYGpGjOfaI8ejhZWvmlMaCaW0xOL5BeDu72uzL85LpC6OtRh1mUTxISPePJJQiz6D/j8oQp
M/UuGKabI9DEZGxDHDVuYeBf6i2obg/l1tG5sbgh7VmetzrxitETcoq2+zpxjXNN/TovCqc/dlHl
4svCHaif66ThzuDJ6Uqzi6dMe5BCDRdceivvZqckAUYCflcFNk9uk8pPX4zMgC6lfRJIka/n4Nrr
GKQy5ykA5sV/F/wAxCBHTwVpw+8HqFo7rbihGbr5WmItYTTfp6N6GknylCXHUD/Ea1xkv5kR3uVr
e0+qFb8ndEL9MsKlXus5Ph+gRnbtX+iFcOrV5+2quY1PcUIFJ6kCXmejtlpkMCfNtTVM140lR8Io
UWUcJYdmzB6fun2UoMhWsUgezhzqqV0fcaHLB1ETkdYoZsQSo3PFVjM+OrIAl7HY3K1lp8UJ8fMZ
7yMAjvBLgSHDqi96vKW0wEhvEBnxduws/CBGWHj/nP2C6AUNqVImB05kwEJ3yQ8Jfh7Y6/2h0T66
fzlJhG0njB35lSMzCHwqc1Rn554r6nfhovD1NENenJ+fVKp+Vcd90Rq6oOd2rCyxFF7TPmCw1A0a
PISb5tR0YJ3UsiAodpt8uWXu+yykBDsAmHCCRt1OEMtf2VFpA6GtUTAdKP8JZAyUesAbesBeAMvy
OUsy/9UyYe7fmzkA2Y2WuR/d2IiwRQkaVduEFKY8GqkjQFfv9bTb/RE97QFdgNtke1htic3poBMe
B2olg+9u7cjVElcZU9QmXyPY1Eex8BrIm9TIiktIL+T2HhEmlXtzSzjVPdosPomorCjU5Fi1G039
lkY3oKiqFuR+IE/X6VSYRT0TA202PlovVD0BKQy5mM5U+9WRX6+5Hn0R+uY8N6vLCOOYjy3ZGci8
O+/g0d3BNAVysvB37GlDUEHNAuwqsrriesXrtCgOxgMfE7jKyCELWrNP9n0CNzFUwcagajX/wb0L
M/qkseBnP96u4VEoxGk7UNxmstfO5EhX25wvUa0xscCWKlWEHsaeLQprPGNVpmJ98qfhWwBgcsNv
E9gbzfyknXgTH12b/A6repjd8ggz62fRcarnYaDktoDKc5XmmnSEAhYuYkdrnyBQRur+gIv6e8Rh
7yf8TcHbfwD6W0IQLI/wIjx11/sHCg65Vhv8+j92IHDcjhlo0hWwMsCe5HN4QQl3Xk9VwXZFHxTp
SdOdHz9SRFziijSfuEkFe2LofeAsyefdPwAyTBqTj7Uyvx/+YX1QKUW99mxjopSllX1/asbhrlF2
baLoQLS1JAlp3PSw/LR/Iy+4i1MkETzObHiWu8Eug3LEn7VxRziAK81x7H/TousighYwoUDtj84e
TtEJRsSbqTIiwkAarASATDHtEMzJUL8JOQzTrUdxaLJSPD0HVmV+E6Q4enMCIb10/80k7V8hT2rO
nnE9NWMk+rAYgE3nCa599RedyGWNvOnw73kedKVuwGa0YHtxqmEsbmfGrJkw2HM9yPWRbjhM018/
IbORUwP/kBQwlURUAfpLriPYdN0RubXqWtgoIa8ShLB4jSJ3cVpxBn9j6gPKj/Msv74BsOe9gmlz
1ohVDeW/x3WUjJwUz+QYXgtADrt1ZeRjI1yTBslfss0jEwpjz+F7PEUZiFofAQHhIQnOiOF/Ihx2
ofkNaHGUf++1CoghboLMA+lRTLQWRvd0ZpXC8vMcEgYngvWTuRRIG84sQIJtq85/sTS5gFFznY38
Ys3ZZ35jaQlav/kneIkTDdAr3GuX0VbkhWO0yi8/orq3wRIHc5Y3qgSaMwHyxDHd/9XADfQrwwTq
1uLUurxQ/gYUB7RlqLXKk0WHNvrVM/PYXqI0KxB+xapIa373cTS0u5vf6yx42yQ4c5M9pRjgWKdd
KNNnueYtjEAeWVV5QiPz39HXBR3QMrVTeYCFhDLADKkGTq+NHyFGyGAoXVRh6UkNuzKAdFbbAFj3
YWrlafj9+v+dWtUusGx5JVtUDCpRfjsAQztBQGBVcUmi1TQu5aTCugN3IubuLWV/1qVql12NhnZF
xQ3DK1NwFEWNTW1hp52KxxzweCHhP9PxTGv/Sv6X9PmtMiITAjzVTRCyr3kccCqhgC2XGLY/xQz+
qHdwf7K4m37X/zJGxZP+mYBPeTMIZJNtx3hJey/tL/FbqWJJLDP9cdoJWn+aFI14CbAKWn8bBXVl
94vzL/PisfbBVHcXs7K0Eu5paWHUDsSRC4K0WCPk7I1thG2XyWdnSDcLozg9/7KUQRqEathXgwli
axm5grrsjh/vuNAi7Z89Lha5WZex+3Suip/xlzRuodx+pWcZ3IFEmcyC7yB1ze0+7iw48zMNUA7t
XIwXugSx1ypmtHmGsdMiLiAocLOyTcjyvsHepM32Wh2AQpA/Bpc5ri2xWz5wI2qAh2m9Zlwe8rWZ
8BLCDOIeKRdKF4Xx2iuAnn3PAxcXGjDbuLq3bbrEE58kU9aK7xz0Mai2nF+mbNW94jK4LLJDzFXO
UCd9MjvcskiwGoSjX38tyCbFiMBIi1QsB8hi29/lbV+LYNqMfirz22PA3KO2NpYrgQ/p5fwAGIHw
uTHdSY4j4ZOZsODkx2PNqMYB/1m5AXDys6U+9dkiu2FBlnRiyUaN93JaAZn4AINaymJvdHYn4x99
WmVvaCCRIlnjQYlrvstL7s9ydNDoBYTZjIMheyo9yyFZYPZCjrlnhp1rRhMi37IBYxBKWh7TCipR
PVQpJqdEBbydH/HVbcMUe4rqiaw3Ngs7uhWU86I4O1jc1cs7+4ZAQpJ+3k9DjFHsvUd/rYWrrd/l
RMBtMhP566smtATtj3hgC9QJvOaPhFq7Fyz4wm74NKFejEEPry+vcqZKracu5vqR+Zaw8QuNiDei
9OczSzUIwR2xTA5mjHSt5SXknSLzuTPKPqi5jc/MHfbOcJRO8D+vLBfIIUfCmDm/Od9tRbprzTP+
jeZKp2Z04epdDqMwQVPhJvimRcQoggn9x3XczFTFaUSYqyPm7QxhP96s873Lr3wyxf/H27UMMcdY
4xe1ug9YNCL/a/nIU6wVyst8CjakKBVdkaW8pSPgQ/lU0yqAT0RNbeKa6lKOY4fu54C14EXC3CnX
NbxF4vZj0yj+XX0zy2tKH2Olp9i20exkHkq9Ne2t2psrLB/p5bo1YwlpCK2pkB1BEvggHFsILmpQ
BhuzcdXDFfLcUJwly0OQQN/G94azJfuHm7Du6dajwAOEGs3ZLpIuER13yWsbgRklZl4Djd7RtksF
WNdljPXgLblo6loUF3t1w2u3i8YntW2uOdukaeakVf7hGbFzIne8+vvBq9/ciuTs6HT23m0ZuWwL
mTtmsHFlSbfXNf5hs2NzQlwZj+sqE6Mcz9718FIApKG/HvWjK5rFacMyapCiYNCaWWZg5/9POkmw
ObDGwUTE1wQcBeqKi8z/KaDBFihc5XPeOiN9jFl+3MI8GIJjeScE1C+kbPZk+NKN331/Q288TNU2
0wYsidgBWzmU1yK9I+aH4TQcycsCEqb9GXkvl6OtvJEjFBaIypv1ZUOS0tGmjqcW2NuC5q6SMN2O
CXqLdMehhRyMAyLobrXsjDA3u7afNR3ZfmmNy8PdgZCg1NoNL9wxKl+DzIWlHzqy4kwx7fSRiVGH
G11gtmBs902b+j1GcGCBsOPEpJittNLcgsAhSrpWyoesz0HNod5kPRGCHCqkdq3CVDek/TXHc7DB
Bi4em8De0F4Cwwpa+cjuXFBUv4scH5iJGCNSnKzKM0PAZRMcUZDUjW078TuUDmvd5t0H6jgF4vkR
LfeANt+IKUiq/IBI/tgSldD+SdPCFDPte4e5pedKjfEswuko6l8lx6Kvsf83abGmpbZjQfaSuF9M
EdzrFWzaqc/hF5PUDpJR6vrtMDLIxPo+6hahrrQfYcehQ/dKVSMMmULKVqbWqneT9oI/L5lefSjB
1uvxaPusMAe49ubAbUcmqp/NBFyLjB9Xw9dYsToQ7xvbwq/6haNclxQAMn8l/3Q+MLgif405gkRI
F0dA5jUpWMyR1jjfW2mfD1F9gqPUJXrfOiyDUgonserxheUvgF1Jb5fVlpD/2bd66UISkgvbKcdX
OYvAHLkBx6YDq/mOAZBEdX0cAq2pwdRrreRw0QdrsBNcn9mFXJmKbGN5GyZHzq10QzTAMgTNs1v5
+DMwtnrRJsiI/CSBx3DN0HoXKMezJQyozmNcOXAM2Xm14QlNE58gM3tlnhKtqX0IeJx7RT9KjNG8
BUPj22E+26/GkAXEzgBfAv71elQdPGRIzYoRcchIvxxaSgY6IbWdaRKshiuw+02214dS8OFqCjjp
3UI6ECV4zSvrRCMy5+D41heseDrMfTQJE9OQNhwUF4y8Qo1WQxqq+XX0TuLnb693lhHEXwrH5b38
se6NhGQfNg3Ckt+qAQQn1bRmTsK1ZYWDL2AFQmPPiYNluJ1Qtof0qe4u4UNS6Ajs9poepJZwiCfH
2MeVXbWO+r/wUaEhDCZ9y3VqZ1FflSVTVBzn5pLYACj6Re26xJNXqQF694vLJe6BpXnTGPLBCshH
sxvob7KsVXr0bSP70w1u/glNAWjj1NfFBTlhAoXbXEYGHDJKh/f2uvPsOmVQyA3uXLZadxmhetW2
jufTBNJutOJS9gzbl4y1p0U3npC+eDf50a296ywt7uPHB7sr9r3LUOvxS28CN602vmTi0ZZzlh6u
IptlJhFvks37SM875KGn/brTPuD1t4p/fGDxTz6ID9ZaS3GAmDgmWZ288iCmERHVDS4/3HVo9Fxs
67KhJcKNoXnd6dmNnWu77JFlR8VL1gOXwOp+qLb4VfN1ikDZc0eFBklwXwTV2DIZRDBKd4qiYSC1
7lhF+jNthnsGMIwCcyw33LjjEdLZwJWFWMFD/WBEE8ujnN8qf3Ia0FAiqs7XDX/GdP61Ps3ukWRu
Ls7CCjT3+u1RoKve3nAsd722fxCPu094VFsIMLMQrO+1fHH5E4ryAZXtk8W2yK7eBhgPGaHXbHkT
T3RzYz9T80VF1OaYDssiCrYNU3zNE66ZL3EKiWefFP1dS1omZjoApF2E3chD5myIfjxruRfYfaBP
u0rEKrVOwXt9k+wJeg36nUlLDLb6vVmQAJenF8d4ZAwjRJue2S6bHs0cwSCg+Lv4hu6d7rOPIRp3
qjsijFD1JZ22/s+dc107pC24JoWfr2BweuBV+3+75Pj9kfyp5QLdo4CJioo3bPp3E/WhpUaucAEu
7rijM94le25gmZJZLvQrVda50WghjynqfFoY9YjB/BesV1Wf1HjX/perU6Ouo94FS5ypQbA+sfgo
6etDsV6QLMoM79PWsTwLMpQ8zTXKt2cebsC2LA52h5R7vxr8yYXwWKwg4fPxq2+lT4UQkSNw93+c
KSMXXpF65svwSXmF01vL2MG3VpPwWFB5obT5IvB0Uo2t1V6fWRU7PH1kI+fhVLAc7Y7fnT8HdSxg
+HWgm9RMR4rD+MFa56jmspO+5MlNTJYIOBA/WMuZ4kZQIC3ww4n7XbO9hh3K0vApWG1BTktvSsB1
qgntYGJ9Md0SFHpBdaiz3efpYRErU7TQlxbD6L9rAWcxC2NMoLsHsTydsiHJvfDMWRrSvzHmVfvP
i8kUAhVdB5jzEbhKYNeg5DZgYJ9gpAJZpFZaEcPPWw+g3kxFAi7Mabzba3FqlkOYUPem2xAQjRnS
+Uy2UUCk+QrShhQFIjbZXQ6ep5v36+9W0BFpaMNBImE3LrL93rIPTtwHXjhL8+ekd50Q5rw0rD1j
6dg7sXxKe003QJlFSmhV59dRL4Slszxmz7kIWYVmg8Q+6SbnXad9xrRO0vKx1pK466y2ffqG+x4l
j6aptiawVV1vfrc+2uS/XFz8IevvrYeQotJc9YDC+WLSOgbn9ALFU7hUmWPQOusXdmg8ej/vOkLs
nP0pkNKIDwtAJF3Kq139uNZ2/GNhRiHVrAOTpRcFY0naOPAaixp33m66e9Cy4+bmq5RkA4rY3A++
XRAs1W9TzvS+yKgLa7Iy6Y4oIRbPWCLUJZH8foWnGWaj1d/IQzzejT7SrsjIOUG6ULhdBPvYUi77
mdOdpXXnfcH/AcIr1tv+SD1nPHxvxBHSPnQ/thfEm+4JmIxssX9BPSUnTHVc7JPTMloOow0vaCT0
LL9lUbo9CtzK/du0lcHZqa4+PNr4h5mbIVybZ0pz8sUdHWw5BLl12003hdeMxV9nfaWUzNw2fAky
I8HlqFbp+Kb2ExYaErMCKnjgBm0bTRESoPUeJJZTGC9bSDPiLOal2z8Yw5Z9kU9eRF1MbgLCqeFn
hAP0nr7JClXm5R8NED6Ao1zIQ7i+y+JVdwP/PLWP39ct3aluH/l6VUae/kzs0J5KHkUeKDjg2l1D
rR/Y6uA70b0Mhd08tvAIZe5diiKwYhzgoXHdRjGiVVszml3J+gxEXfO8AA2MiP9dGcWRzNnZv5oy
TMKopwzVdbgqkNEl1BTJlg1pWrnmwL+aZfO3GXWu08udvwyQc0PZ7cUByFQo42/9iN3VV3ldZfF1
d4n769QViWEIEcUr9Y3PG+f66CvHkm4jj/TQP0t0W747lEfIejlyygg/jlTAw4xbKnCp+V7FCCe4
Rty3Qp3+4RkKtJD6MmZPhaI6CDUtPEdMR8z3YhqUa5yn4h54Hfegd54TUV2EgCUiJBDv6WTK/DGW
RHANpvnqIOO6M6Y1a/NXMzbIxe+BYwro0OZzKOJQT1yJrVxsBkxWwygor2BuOovwYbUM+QPuqlrS
8oEh7NSBj8U5vuvji6vSYaIGJQrx9pST+4UiT61o+TnVET9ngpKKwi/PPXSmeYNb+zswkFCeDzHA
yYmywa0DjmJnv8flNhp6T5uaT+irb5pMeT3whf0/RIXrhN6WsrA7i6eB7eqqPpLHoZFBRorij4ww
RLyhjjCucioVtIfRuJ4Eylr5tLK3nUs6w9fbBW3PZ0q3l8fi0LsdSubXL1ZZUoPLLy2Dbo8sd/Hn
8J96/wHcnZdtRBhVVia5xcTt4sUxDOMPWm0hnaiExE2V7RHKir6PxgIHmueOfx7yVVjXnxY2dTFY
+n5Hhz4axZyCIkrhqu26Ie+mRS33NPAnFX5gFP2cOUwlnQpO4l6h8hGy7/3LTwexSKpphsLylCXb
uMsPHcA+lYuB//8OhRcM8iy7wBpofNB54WXU1txd4RiHyqPnjrwrjpYbl0cc8u70mtiOJvXse88G
roUNrHlFd4qAmbjSqAxy3pcJ8SsSm3KX+XjzwDO31UXiY+1vMPcycTDD+YRCfMH6d2+8TLI5ICun
rRNr0pPX6dEcZQfax/95jYvr6D9w+1lWXAHPs5Pp/py7CBFR+fUMkxuo0Fn8bz30A6P3NbDb94rP
75C5ZIkgv13vYnL8HWzxX9LqYeuw95TzCyukLmkYFelBK34vL69o3JSEYGp9puEudvIGoqHtCVaQ
5kWlRUSVLgaKeXtp6nPlYj+/tSvwaVaMUNqlNfgKkqkHzyXucgkzDZyNtBAcBJmmKtx3sKETEiRX
mkFLZ6Y3A/XG/ANeSAYirXAGDEEUZQSFtMCnx/2uB8bmfEZTwMA/TmNWDnjp9lj60nby5EigNWfs
2L2Wx46UBYbSMOm8CWvOrXLma3ClzgYChu/foVgo+FJb6WVMYQ0Tye60Ux+vWv+wtBlF3KTl/JCW
OY/C8W7VYbL9UXlAaTZCGxrMiLaQHa/npBxHqk4hdwMq5A1Vf5XV6P6NtUfU0dj20N12FqGXg1lx
edtrnI46iWDRUnwYyl100/lGXUlxzUvpZBmVy4hrWNRSLRkGx9J8KquY978U1dbDUkJMDlCHHZFB
XYnYMHjdQaBKAE20HMnU6VWQrHvSJd2oqngMg7e9AZ4S2c7Nm+t5ECO4YEwORNYGZRIK16CDq1su
aAZVxIx84kjW1YW5pbVqx1JvDutKkYcQch43fP8/Uygrq/RW7VDBBB6PBzf8GFS2QkaQQCd1WIrq
uHFQ44XbXFF9ZmNvRPb46zHQsQ4z3dBHUEGugIh9wGETqTSr8mEhRyee19XYbOpJrl7mQfeEwKmB
mVB0DaAaMC46fLyP7RDmTEVw5varRWKOufZhOky2mg4BvnPsHY3tXyjBKEYkCOEDlkE/ecOozJUG
JbPdB+htmPbV7/7BA7tNMcenqjEX03fvpodbMcxaS1X3fxaCwDsikfJvy5UYHZl5sBnrXAo6DLk2
XyBlbqBxNu9fsyo21/+Z7hf63URUR4xXToI8waky2w//bcKyWLCJtLiHtG8BEDPkvrcH2wnwihEU
4x0F+3eUdoRfr+yzvOsilQ79DI1WOBLtlbndAh66eqyTY+Gsdi0Ytq51s296jhK4ss/+PdBTdG+4
icq+U8vBJM3F0qcV67gTrzsC6w4aDRFLuPIgxfwgPBEkvDIHEdX7C6BORlbg0HdiRva5pcurnLx4
3S6FTbsOgyb8JOYWCndWNTyn4oBwk6Pw/zTepwGBWqmjtmIjMF9BX9SQCL1cU8KD2APjgA5PwlI7
N8J6gF/Ws6FP0bA89YyXFb5om4h5YQhg4ntpD8WGpvq2YvribMZNJEK/OvqxP9T2UrGtuGchSlCj
VHp0rufsJUZJhgYaBZQg+TdSbsaOrPEV9owpeZG3YugvNgf0ZHNapvVUS/B51Ca9Ug58ioLWP+uE
5LPi33d0yQuoSl19KYwqO5SJKB0pljrvhdotuR6yHso2HkDskx8F183HpYyjnUOjzqpqqAUxBp79
e/TfNNaWKgl0tCQ2guisC/O2l6t7FrRc6nD7hzBxvw5XFmZig4GXrgFZbnLVLETX5g0CHCqMUO7v
duG7jHyF6NKQpJ03viBFc5p1zWglDibiXUtqe5h+lLFQh5/HyR+yf5eeNH05ElF1qyZy36tccsYM
Sok8SRentB2ACEboX2SmZyda1OxLccl1suriB8dEYjK1x7aA5yOotjpm/8Mhz749119q9ZrAl/PA
scVC7vU5GWkbNVgs4Oj77nWWdyZc9azme0ic61Pkg4w/nw/tSNEEX1M6Is+Z74cEdl5d5PgcNw3/
GU92Gi19+g5Hci48Iy40i0hS1VrQII0+cVX3XA7X4pL54K+UpCiybqo0KQoY+IXHZC6JY2yzpyA2
2zSCrKP6vkBbvFCGE/l7uwbXkmAI+CJ9ktAx3Cu2oHzqgLDDIT9BHbFJIRiQ04ioH6udi8YlrLcQ
E7PpvV4113/ioHm5M3ZqylPm23NLD3I4sXqILKyO6b47oVPVV7w5IFPheqp3IxtQHjEqoicVuPWh
N+9tTnSnfQfApK3CmBuDOPKQdSURIIIKDDzJNsEg++uOe1aBI1lzTIkEfZilmRpJrEAjWz55qBzs
Q1F8haQP08y8Y8UDQVJo9S0XnLUng8ZRg2PqlZESqvmR76cE8x55e7XGf2noApWQ6LKfYxFkhnyO
CoKZhdXHX7lSwrmZaNieC6QPSWhSEn8EvU83qWjbCEVhdQ4PMklunqt/VPBwoXeW+aoCPPnEg04X
uZrL3GImLvuamytkZgLCyp1I6c44AH5hpXcsgrQHMtioYGD/fZ9EnQ3eMFTAQ8VvgalO4Zjc4sA3
XpXP0/0Ns6DEjAls8TIAKCaMEl05t5Ps0EIT05WxB5kVLXI2VG5BnuHoKHfPfkbnwCd2BeNJ8xta
rnRDY4vz8fU6cDMTTbjl1QnLWSBkuhlq0ZTxZNbk1hvsnyzsy4MoFi++AeN8QG2t8Z5IHrVajEW3
y+8lrGSsfjaIjstHC/H0a8KpWxXL7+WIgcIrvRi5Y8ecxS0dVDyzsnXk1hBaBJfdsgyUBWISkOVC
huQaiy1+Q/dnB/98LkoYlYSXiXvNaz3XQQF1nE8dQqMvcFauOvpoEwHcVYhCYzZPi0WPnmKv5aeU
lFlAd06RelFOgbpSmeKm9AAMJvWpsTx9BXTiixe+DyURbM8Oq38UxJ3M8bwI23IPNXw1X81LQNeY
oCshzYbZJNnd0UxZPiJhD3hooDPU9V35InFBwVpuu/RCqc1vvmG+eI1belA2R6I4iPpYLNy0Z1HY
yRyc4r8ApU7crxWhEYW+uSyN+Niq7y2DkixgT4h6zlhKqdKa7PdZysOMes3dt3wm2mHClUEIwsjG
TRmgP0z0MW3GbTBR/QpI03PSszt8BT82wgnc66pC5Ke2ju4lgSdV7ylancpSt9W/KadFIyr/QIzG
kgko9/Nx4vzc7H+QI7WebCepT+QjEReMX+BbGjf9Q9Y8R6BRimXywCzK6GzM43gAAIx7TpUBS0/M
MnsdjDF5+QGO4+V7+joUXjHJvp6yoPRzrnbn2WGQClI4Y2ylUFxDtkjLA1hcjmy5MKHpfdhEkjOd
cxUJzoJaYBoidR/CZ+UW3WcBoCWd2+FMz+QeNAcT3iavaHRO7A0EwKTcULUN5C55aihE/vWd8RP9
osKetd5eIpwurUQs/aOPZE4XQZ7qN+9WsGCSNtjunqQAh2h2X9VZbt7opaSgdOSVVkt9jBZqMAjT
IUecWxv8uq+lwEMPk8p+ymRTCW6E16UU1CeDPEVGcSUy4Rjm/pOlmMaakIwy8PpWUj5STib2vZ1n
k9pOaimQeTFXjRtPBePwVnoPiJfT+qRVbXHPAt/J6YPSgP+6fZsEN4IP/A10g57kLfvkNTKh/bSn
9TdXgtsg0aEL0f4367F6MlJEZY0A1xjwiqFPx2mbfcqiFu63efqcGJ2+FkcZZzJwwE5pI0pImV0d
AAfGKmVVBuJcrs3jPVS6chQcaYIi9C0jKctN+K651HcYYwdvp4uBuiu0mwI5n5XTCJs83iHIMyY0
7Z9xe/2/n4X1IBDluuitQHVXAAQa8sMcLtoxnE+UZD7LHwTRah9a9tET49COj6e614L1oEwc/mtM
vAgZF2IcT85XMRO67FqDtdDmJWmcsAovAauRQawKqFTXACtCa/rt055COnbJlxAalwVM2RcIddRh
UqsrGZ/IeXIpitIGTj9wWSOfkBMdGWwlstXsSEHfiBCrxoXbK8vEUhryC8BK+jQKzJUPhpTPZqnI
lThBqjBGmVp1/nU6ZTzLum2Xi/A0DpdWm3upYVGiFlrzyCoMKcJKs0APeonPkkiKXtcTMLO9A3zA
1lKwNNDCOTj2EU95j8lnXULcpW2BjhGHrTbTU1Mvd3+t/NTKiMqnIxI+MYvH+w7qCxbljdcj7jnX
IwDP9uFFAW0sp9oyIVgQfe3CB7NLtwht4wzfAJw6z1LXv+3aRaYtyyCnOoq5XHg043ORU892Hyv3
z2kkTgoie5q+7nO3IICijGinvzBauuzPNc+DEYw1hw0zuPB80fdENs4LnAEfg4V4iqQTWKf33NJH
HSXGsGBijE4zdCU4rIQMqP5dChEd1cDCIsZ6Lc2nDhr0MZqJ6NiJ7PwwsSuF6T+hDUR2Tbyqp7gj
nhzByY36d6MIxZ12NKgy7yg/BYKglzlokd1JcSJWDGWm2+09/A9kDBib/tlV4Vj8W6IK+sud1Yk4
deZswIGO2Gc3Itp/7sBo4iAzOegCa/49blIZrsVORj2cPJu4qQHVXTWnjrEfwy7kfTN5t3HnW14R
9yYRzFZv1sOtBJVQ41/GUO44pSL5w6qBiRjoUWjjDmWN7Exz4v6uvo2u3Erkdaxd09Yvs3N6T4NP
S/8jto53B0/cZjFSsopnSTPJu7M/VqGUfYMEGPPj3KGJoAJWPlcIaPbDhYfAfEfiDNbAn6inAeRE
ZFVUYxGcUc+Ou0CWA1cLBo+Z9UCTJW66OO21a99/tWonWrUKRvGu1Qw/7MR0ZX/cVCm8Lf/vKxbF
NUTuUBUw5GNg9leLnpspDAQLz2xQmtDyDNq3qvYpfHumL7QqKSaC3ErSVOUVgMrbHKwCPkJ9xW+/
BFa3q46KxfqK1A7uo664d1P51FHKxGSG6z+nHguUuPfnuUXO0rlQz9RFct/uq3G2eJlXyZgjtv1H
B/CjeGcpl24hCzaiVuCeSv3tW0wKugLcC4qzZggzMCe2Xk4NcNmCnOwr9F3YvnWZmV7bTdBL3/4a
QeKyUu0K48opQLQyopEWNHI+uoSvk3LcD+8+/+jc7t/Kt2dQM2Fx1pBKYrt6qtbpD49cQo5qWRpZ
fyx0QEdTUN8LMMKxPtKFJlAUHlo7d/ORnSkRSCW8dwMbl+VNyKCzuHMqvfnfU4dwDdqi5b3A5BUo
spQNJ4H2orfw2TSdDNmqVj6OmUQ4g22id50dqb/3orU+7X2atEDrAM2SYqkzKMBxaTbCU+H4U1fQ
HHFawujtCkb3Vwv6NF6heGOdQh1GHQErcy9QY8O9+dFigyYnLYrfRlskqc8Tn852izDM0m3DJAdV
zWY34WyaxBCi8gqZWdFCt05zRwZJX0h5NIVyaYVIkaSmsD4xxMIPsKPtLsndsD+uZTp4ZSvu19yA
3fZoIKNM86uHbYzGsM2genMeDA7cbR3gnD8Tjq+R1PrGDTfHGC7DOmR6o5Knor7UH9DRGvEUeRhf
QFCMpqbuLQufT+BOj+yJx3Ukk7KYrrGUStB2WMthYsgrDYXbhwQZ6G0EXgstk7BqE8oUtr/GABJ8
2PJEZKPhGXFOyTj3xlXeGhWZUeGg735yCZ0cCeqJFmJKflgWRGRiceaIVoCDRXmlBHwO/7R/JMlN
ObxDTeTXImozH7fIdzCK8GVhHFgK3ODLglStsQiA5Y4ahrvVXNGZahOG5oH6gcl5HYDeVVQ43Coa
UAc/DNUzmNMbz3gaZjklXazr3Ap4HIdI2ehj42lcMtgQrOh5eq0D8XVauh9rQ8Q7wU0Q6TGNXFPv
oxa8zZI/3LDfNXibN+Y5pLWn59KvzQLhEfmKNJCVPbWhQsHFjBOq9l96A9PwT5JqlCIalWKrsudN
gNwJ4vWyDJNVa8dIELhDvv+o/lqRVgH5swsKGdD0plQ6vyVCsOagj2bwXssYJxm0oGNAQS1cQuKR
uvR2lw7n5R3qsvHKbAKMwhgWpSLnm9lqcNQroKb9AlLmOjqPC78YFc9VBP7nEt9GdWLCeSJOgcUj
nSTdyzh74hZBxcIeiMJsY0YBeoJPbj1GijVNDhgb8liMDmOK5QU4Fxf1CH1AQEtYgj5eblvKyNrH
xK2OshaCLiUgFTh68t4XUDIBd2PqFjNxV3TFtU4l90dCW3dpya8Hd1/0i+a9uotfLNkdq9jpPyM+
FIx2OmJ3RrRrt2s9+vZfyoQOvjdL9cz26P+dra27Q+8q30lH74iPSXhZnnCt5ia2tJ+XUopI24q9
+YTyYWiVGt6sVs9QdoP17vV/CGvFHK2MDRa+GxsznEmQL6rPqf1pOPzAJOkCWVqhszNcO+UohY5+
k4Pp3ZPzv+SHGf8R2zWHm70iToZwCnCPaSqX1oBaQ90T731czpc4pO9IPFTuUDBcNlmET+TYvtoM
jW4JF933ylmsGznaWcxWAkv0lhS6EmbqllGXUeuJ0DVKMCje+5+acsKVVH6MTSfvRQEWsnKd9/Tr
HjRH4oLG8HDaI9bW97QaCtVdYo4upCis2TdkZttznY0+UEkbA1rtg2UzzosiNTCYDuWL9Zp6uhYX
cKr6k8HXG15b82vOyiLRkI/MzlaO1ePs0frlwTl7M3c3LKuYtB1874SzuAQItnYu6Num7BlJFSX/
r6/ezDBY4oPO3cSj6IYCMDrwRfMDh/uTC1wyQyGSqSmXjvrfu13n0VSfYETZDxYVBZ0I31ZKOdxN
dzfaifn4bvizVlgqLOlPVMFs9RUCohZuNNPqKVB3qknGqhYYEBEgrCIbAhxyUbG8FjSNdOibBZDC
n0HLiLCGR8Ilq+LzQpI/N7DZtpA9XVn8MHwp90RJLzvL7nNV4MktEX4sl9T/uD8sYnUcj7vQCB4d
QoU3rnvv25plGeLvz5SF5iFCHwG4mOtAXcqZmXPWBjxDiWGRhumKkipHY40zago+pT3zwmOin0Gj
It8bBHF0zQEt3IF06f/60/LAqhcHyekGYiO/tI87tbYDy27yUwr/vSaqyJr7BJJ3Sabijtm+g2Z0
fo1bOZisIsVhO0l/5+lgPX0hoGW3HL0NO4RBtlSdEXl3njZa8/b2VoRLqfUog51Kul0k7vc/KCQD
2vQwoquPAUkPpw64FTlYJimKE6+kxP87/8dMRcR9nFyw0ze2g9OrDVrgx65KmYXWNevFf9eD/4pi
Usm4ztNHrLffunudUl6jN5DONny0VxMQy58EsjjvmPtSFR+sTT9YDdA6ZvNC1m4Fux01Toj8r2D1
lMdYH7+TT/4Aa+CAMUSsjqNQXB6Iuc0NplSRwTTHzN2Yz2xLiVCF/cRiH/6SD7LDCW5lFAROO0Vv
49wslT6zsSpH3F+9LlwDdSbunASLuVXx8aGTuhnU86wEZJ2JoesIDocVLMrBOVWjbOKfU2HAAN0N
fA33rfh/HqGtzM8NRQNSy/5O1pYcdhj+jqJ0MeN8qfCiuqZlUckT0xAAVcx0EtmgPThWaVJDGIsi
glckaYn/nAabFxdFvUsxDGZb0GkQB98Z12+cqZS6y4ip6jC5zVJTYo6Vr3aSPYxRv39eXsRhaWhR
IS+jaODaeE974nBJqu2dorSwUXxG9PeCIVpseGvHll1bijHasAuGkrV84aZr/e0X5SXxJ/luHy5s
XqfsUleMTUoqPcmtEn2DzKLWY+nJe38MHjOCYho2LETXYKB9JpqxNukffM3C1SHjgPg/viIRVUqT
3E9hhrEsy72m3i0i/aRARtDgd195QZTH/RREIASt7g/uEBHpxnV/NwJ0LvkYc47fTHPhQy+WZeBH
7XohbgwwTX2flavP9Q28hug9+wi3OWZrk2/DICkuZBmOULMX2h9nO2CTTTiuCGb7WZLQ4cLu6R7W
9hE0+KqXTHypCMRizyhT//mekbQtkQQsyW0jiXwIYHVxh1zT850cItFchsP7/h2lXYA3tgPOS5qj
ydLnEWN5vtfKA46IGizW6/sZr/2+sr65Qwxc8s1UG+am97R8rsa9o3bkXt7U/FqkpTpn7PJbY96P
Rc3eGF/4O7oAGQvgDwuCk3uta97bu5vLg2B5sGb3DhBhxSIzbdECwGCBDPgFSzgBfH05ip/hLq2f
HSxdTkcxAuCQzJ5cZK5ivINeEq70Ed1Sl6rxQ3bDhgw16rK3ny+6fvO6/MyVPBFbFX0GbSjR0b8B
dtGiNGWUAojJIHAfqo1QMlcHCoLaOj80Kfjjk0nHzgbwXTpxiruXtIX6+ifdwlWivIWxbtgguH3n
k+ltaTh2gUwBaG1FaIirrRmnzC7waQ57z8tjkWlQkt8wpoc2EaD8/QFlw9vRXVypupwzMnZ+7Kp7
a8VN+zFWPsZ7Sc1a4HaV2lThcDR07zSKZhm8QNGDEbrHZHt2ec+LnyLhG2BVdXNYIRMphftyM4FI
ktnyXpjBcjS5j/GobuN1BvArfu04RuhNiztv9S4PZlCnnH/tfmq/vGwbZQDCJbFR+nYCld+q/D76
XYLX69asBy0v4WFLQgdDAB+HXRSrWbHz12i+1KjCDpyUGqDVIK+Vt6GyWyRaFE+0ldYp98mMJ17X
DHq8a45ZsJmdRSPjGqPe3UgQPTpjcyxZFX9mjkA9+aEDDb/NJCwfe2YUpO52Sq5y7+WfnXPcnZmW
vcjQckeFbOr/ikkpsKiuxifRcvWRxj6fjGrtPAQgOoKLwHBLHi+YTKF8AdR9DI6mKcBMU1gj2F32
uAfWI8bMN6CX00c7i6KYxOMeogpSaB5/nHm9geComZ4W76X9aslyy7PSqcGmJe5TFBxEP34V9PML
jiH7G7YV4LjzV6fp6bjmtEvNG7hnyJxlpeCFGecEAm0VQWjHuSXnS1PxC6hVF4qJBIJbpJx8EXtC
lRWjTbhE9dNjvKRgFg9mPUQqOjn6nbbswKdP4xsu9yVhach5b/qsxP2HmcyILKpnRZB1BsPlzSqC
oyJdnjJrS3ipyo0ARneMpgdaoIlzL9ZAqjBXDeDeYw5bxl+n0ZEYsZhmPldFMouvjufhFHWBgbwt
G+V6omfMOYUjEHLn2RGDtDzf2Ix9DQXB/d1iYxJHR8TZ9G7FvGyUrAVbHPhKNbB3NwNHkJsxlJjQ
7618Y+zLxZVn2MGQ840qKQE03XSMl6C5c7pGg1f5is/mSblIdHGa7ltshw6sBtBPSZbaL+d4t64o
HQ7oa9aaeIY9CZRm1/8NQaPW3hrqWbssZuJ8vVSfbnKsiQX7oo6C2ce4+dktMxaGtB/vCM6Tcnwj
k8ppTiP2Ux4BRPkSlxZ48IeKDARys/Mfft5LXew6anvOXDJghgBt7DTwsDDAi47cYlcLLAZbIN3I
xSrwAEs82oL1BMbl/vXOrZlEmaf2j/ZB8oR/Kkb53vmcGEdz8oxPq4V0i4ntWXMv2iW95vWNIPPe
1iuqSap+40EPV4a2qnqGJp6pb8m421H18XRHahqpLhCT4vmNYbfE82TjRobCQjjaA9iDSRZgv0mX
+cat9xjXFqp5ddYiOrTr+LzZ9FI+KrSquCj/JQtimqRH4NZ+O90QOsrNviIbyA3h0rV8KzwQiCsa
P1OXDUEDAOh8A5S/Z5ZL6VYlrJdEMeWv9C7YWsMbg0UPYMPzU0prR2kU9ub1WpNxFFOwASDN/yxC
kF1YWAjpViU4BO4YzRT1FgnN8S026ZMQNabj3n4O991neDZ1APzHdFDCXPPwjKRkFiv+IqKi8dNp
LzwmeeCl/9knaDxqnJjsC8Rya17+Jp5zeW16s5Ph2v8B0t+6VWQrBTeXf3WmNGr9DCzw5cgu2og7
U8jGjYEFm+EQCQ4Nhnpu9GZn86jMyLjtEI/LBtZO4JuLBwwatZfOJZVQ6e7eZeYSh0xt7l6Qewrz
R5zyNQhptfmz7zPygvyZEYxU/dF57fIiLp2NFr9pTU/v06Ji7B6Aw+FaPqgkx4cc1jz8fNq3sSQs
hV5P65CuPZlncV0O4jOudXkW7Djqji+TSCFW5KYd6TitRHIHAt48CifkLEhBfeWPFyXiI7mADGnJ
E2jC+vvHEQPF33y59u/oD37uR4SBXezAJe+y1cZEoqlLhLBFl02vxeskfG6U0XxPSMZL5ddEZ7a+
Bb6AxjdTHCI9LKgDliyrDmuJ2+Jj4ZtrCg6q//i/DWvsHJqn8ocVbmaUjpiHKFtMzyrJazONAYH6
6jFRifGb6rsGOmPmGUxOtERGanZzM/rVKIYStrIkvLgsqswaexKpY8W80lTX77mM0tNi9yr0mwhI
29iC3yzTtMYGRJyIP+AnWQfW6qBQMSumRSGG35iptXc8VTgNOd57lepPZAiQNMLtGJOrLQ/mmbsT
UV9UPvXfrLQQQAKUm4qW7f84MIdwrcLnAeJ1lzMicX+3tDuOV3bKiPxOsqs/ZK7AdWYByQMtG2af
kmVsJcrCJWuPYOfw7XBqDmO+Vs5/AkSEfnLky6CE08hqPcczIv7HRaakV9YJqa2g5/0/dvNIQ6r6
g2sMbBr4CpN+qCWOLTdFnKrjU0WhYD47IVIrVbsF2L34wBEX4vfjs51tkflcVETNOCsaovswFlEB
kWJBFmLqb5uzX+ewmpGW/LWOLlXEaHstJmGHr1tgqS3nDGsNpRxFWWM37I40Sc2nkVrBWi+lp6rJ
nAKckQVZR0CGMIMQhM5b/ruWEzvwCGQduAQQ36KBffx8T2Sa1Sseus5g4cGX56Bxbb4fIlm7ykff
uNwhMaJUYSxRuGWfo1XI31SBt2YeVfQFgOHVJSXOlNIL3ijUAn238O+t7TeqNHKWBIdNyLtVzlAT
iv8oyI5LtNrnWSh+gsMC19y/S4fc6tm+SywiA6HKmMrbKTxAxKoPbyY+iN1XJNqfXhshqH3aCV0v
f1xzKVyn/BAeqt1YeU7wtv3lQls+NJX8angfYSm7cdY36yV0nGm2vbJ7pgHaBQs6xbhG0k9Q6KzX
7T2sOxf2/rNlV7oO0g7zEqGUMiTRoC0pAeTkhdZzpYhPfrwDrzo3teVWwrG6cJeRDnGW9DwwKBhf
VQGy4k52TSoecmgUL7GWR57X91UShVV/2UVXziF5kMYIu1s9umnBPgiSCZBHeGuJfrjg60DV6nAR
cuBLxXRbUzYQb6OL7uOfxOY2YNtJpJIcWay6inpvzXxOWl8OkJUxWTpQwhJZGjlLgX8o+ipvMU5a
4shTxKmVsbaAuhpY6O2jZa89b85tHBGokE1FnDMbd3MoA6V7QQ9trCBMp3bCBQE2FyvZmLxk+yRH
BFLoQyfKXQivY2EXO20gzultvWEUqgF8hvTkxqaqpaG0sDNAhA0B0rbIh5G2XyVfBIawibywFPLv
vXgiCXOpynaDhN/rfsxIBwPl7lNG1D1X8lHVpmZ/IDLlUClTVZXjhE2RMfLtaDWZ+ZefewbRCseb
Z8j67urdkISzses9fLGzZJF+2zLrgm6MPpJ67kpZvki00okGKvmavBemI2wgoEUvSe7wb0vbGQu1
RIuaEEaBJ/xlSbmCoixJScmqto5HF5LVMqSNP0B3RiXEZulW9xAlRYhiGh7AN5K0KaAfT5yEdiCp
lhr9LFBYsokQ63/KpxflUVYWcKcQ7UVlIZuvfFk8qT5TFVCj4NrNNawtXFS4MpZjTZAm7bbD95Vb
emz3zxGN5h6JNa/EwLGi5RXaTbEXE7/FtuANVYnIL4sYcluoZleQYXhRSUmHDLzyZzdkpGxKhoJU
jWRjTuVFj9AcJumEsbTj/YYWl2OD1FL4P/0OoF7YHijNo18Gg2ULhQv4tm8GK/1Wg8AVfQy19ebZ
InYrXRJwmCmiuGDeAJoUB0dDhJsnh6fb3VfqhfsfZLi/wfgu2yDndEyw/Mqvvti6kNzLOQVf9wjg
P9vGeNl+UVS3uNvjq3iCxVrI+ViMsg+HVlryxsdi8XcSg5iTOenwY2l6pZOUxasC4xSM4QMB1EDw
FrWxlAtbx59KCWjId2z1D6NMSaWX8bK8DAUNuxmjaFOt0NR2vkOqvTaprqkQQR3BgyZkcOxfED14
Bzt9chXhiOp9M8P2rd9MJL1zXQ+QCcypWWO2fCCrmnL1Vc7+WeUu/JeK+q16pzQCnInbCW02PlG3
kjH6sRo8qEOwakCsRff5IilVhm4iCAyfhPqrru8c3DzjuR48RMy0EH9LsrbJW+0km4dzkEl8rihG
giAInzsp3KLkiqHssVgtwCu9SoNrb/Eqffty++uqYvV2fr5s7LIk70enrStO95WJSDG837Kjga2r
+sGD31ANiUSRFzmmBHTPNLDf2m7OIikdfk3/OShVhOdNFnsP8naR3WiDGoW/6ftJ8E16pAwU/EaP
xhbQ4SYegTXppXCPe+uYAJbmWEIITnPBmjxX3mpJsxc72KiF1bCGTsagOBomWrnfirNJdMrLRomQ
AN7myWfen4Q2RiLvjwkrYLDaOGddpXJnHwYIEuH/MhXh469h/upN49QtGuSNSzpdXdnk5cUkIogC
c2pUPWBoMsCka9q5+UePiKaswfdumAyek8frvkF9U4tTxPvdA5q21Tao80wL5pAL89HR/0xxljeu
SYIQmEUeTwd1xFK2FdkVbXWGbtAgcPTukWZ+8EPc+Km8KAEM/Vj0NsBS2Wq+Y5ETtIc2HSSXjd80
RKmus89e7yeEdhqdMJ/DcjILugIxQFnpH5078dXgU0TE4f94yUXQVFlxiwWs8g7PVUeBRhtkmkVk
96cRUV+DK1a3esKWYpheqi2glL04THTA9nT9s8tNJX4YwOqT26/pCLVjmNwju0pycKTieutXU4Rs
sgPRxGZcabYHxu+eeFOiV172HIZOr7awdCQNgoVBfgSxCkuww8VRLXL7UFbfyPXz4md9ZzfbKtne
bfHH4MULOKpO5C5jBPs3Xe/54zAKIIEao9Amagltc5MRWzUf60dF6NmbUw1Njuox3x1vnj1SgGMu
7U7neAdpSAqf/ntbCE06qZ84ucqvTq9WCP65uoGDxQ1UkjwyWdSKEkDLqkdf8ec4DBMs036biGEL
45K6EkDGwjulogWaQLkck5VvadAhsFZxDAottJBsvNdZ+nCkVIUNEXlFDl3yeDRLCrK/bX8E55Hh
uXkBDmUIqx8e+LvozO4UhwEEAYjrBEPBjaQ8TUlDebTR0ROuXb4IeiH0UCtMJe608rs40V6mqIYJ
UqfQPjyOE4JI+gDc6x8VUN3fTPblgnz7EMSd8biPIVndcRaQtZ8wg6MJVphst13PZZKhNAlXr6VB
nVQ8XNeSMDvoLK1fjwNOERUvHj0aOADbcp7gzDVtyLkMeVnnFvzfNL5LYnMNvdeVxfnMCVDYiYI6
noZKx2SWBadJJB/Z1PjJEFw8eQkgqBzFYcJKH2ozLSB0OGel4/gM4G57uPpdJ/F8bBAB4+aBGXs/
jnxeyAdUGzCWxffnxBw2iSQFI3nC9K2xfCdKYPgpp+kK32u0ztSb3OuUgVKV6F9vM/T9iwOP3pHb
IeYLvc3Jrq25g9oLQjQsqX8Bj94juU/nkxe/srJLHjQ22zEfBqEvLTxO5HE9FRmbJ6i+dqDM9xUL
R4tyMv0hyd8zTwVccsuDx2ta+CrX9wKQLkBRsNRkmfufEzr6T8Ott0ePfHI98S6lf/aWiWGZysDM
TgLl9X5sfCXpFRhH/9k+SKNL3i+X7J8enEGYwtQvjsc/wcS1jyrjWsAA/4mn4YpGhz7Ey4Bi3cMY
6DqbA6bpBbUQ1W1681krq95qxXMZTiw/axButGQdtPmYKV2G+7GG6faSdbTosShfC77xtA4dqORy
AyuyZ0cUQhbIvxsGFKKOKxRpZEBg6atyxQdT7tkbq+nkvl5e6oumDUORZiV1nANhOEXn+YJ+vo/q
lxqmFD8aW7TOrxobuGI1roWdsY+TyEM8ul2nR72ofX4f+p5FxYXqRZ265u/avKQYpHEw3jhEoep9
XhO61uGwph6Rxg12RMJMAtYnfyIKOr+U/jb2nUAjK6LDudif7CkkIMC6g46ds7XuZvIiDowrjxuh
XAMIJ80M37wA905ZmaCga7zZrRvzdeI36w/zUhWmzeLFiRNOqlZAwGeVWFljnqlzUwqJCk8/LnAs
9cCbTxFkfMNqf2Pc9JhEovw8kPBVFjwCzKHqgTghRTxF4k50tQZCtrq3hh8VWVuhxsiZJf5wo99N
vd+/4EoeYE+i+uugzRrxfxUcf608SEk2XmblIdmXUcS+zNdzqjPA2eBLiKEAIjBEbH2IxW6Z9Ecz
NtyUzTzmH0i/t8NmIzWJ6xHvgpMCi8zRsaUPlDLtCUv0m8pP7FN4MYoviutuWQK+GhkgN9CfnB/2
+fpDV9ajRgLTM5412//PJRa03zx9ryuIVHLRmEb9AeZ+A3xNlxxHWzAs0N+L+ugfbnIOQTZNYvrv
EdRQVazm7OJtEloL+6Y5EEVJg0WvGocKXboXxKPlxiOo8pEZEOZbboAlUYzPmyhcc1UfY5mz66mr
KXi4nU5yMmUA2t1PrfijGPwK9wEXKx2Gxz2z9QZ8sDKTCj4hQvHEmXGcjruAR21cjMHEgoGoh1gi
D64Z5TX2HkRyBU45KfD0GtQOOWhdVroGVnWmT+BL4F1UaIGY+9AMXvRJ0IlCsQzGtBZR8uhoe7gX
FiVVJD8UCFQOp1Swbcjhrw34Nn5iCQjG2/t54D5gB9C1oadV6QPLDe9W0HeIVwVNs8BBqYhHFHuS
nt2tOUWTvu9kEL3bZvLoQ4FIDKsXBE7AhXtXBJYHPcK09sifErA1XPa04w2cKBLM/KLCnJ/7syPg
AR4TjDYRP/igPc16wmF586V92y3xehme1+bjELU6OY2mnBri8cJgG1yfFT4ABXfTFQYL3xcyTSjJ
09frxzE4EI+zFj2K673UPZxvIi8CVI1cpiOwDxWSQ17oM6+wcxIfuvYc0uxLHTfYyHJdCufQW/nm
X3BJ016vBY++fsm7UXwH8zlCrK+HsihMkWq9Zwaf+VgydVj2ToJFHPFQ/rKVkg9A4gyNBWkzpWUq
9IK5I5rR8lwKdV02hWlwrbrp2RVESOdDa7lqut12qt7iSzMDXwUH4iE/R/bZzrUoBFh34ceVMTMV
6RLBODZyU/onMenVC4D9WTTUV/n6hLKW5rgqk3X5ZtlKjJfMvyVI6FAtaKvgJvyZ6wr9mO3cCMn4
JRHZay8X56iOdfbdKx+kuygW4HztZreynYHkayK0p3Zx5eYoZZ3ugzVPHvTBbi5oZSZc5M6sRjgb
nTFupZm9gUidfZ/U1pN6cDnFsZ4LDUuRdQtLbAeysLAB6yAZ9S92h8YFDs6puKIqFuKW7BfGgFlU
S7dXY4nsPkqRpMdz/mPFCLksaBhiorfrII8vuCkFXkNKAEKsK+Ov8mGiZeDjgSQQHUjr1zrNfPNj
kHbBehZqKQXcOU1Xynns7wh90eTk9HSxRBY+Xzxy5FZ6kPJu/399WkXVs4B7WS5J6xNZizW0qm1P
tgMYeb2KqZ4kLFTeAItrN4Bsu2Z0KcMBouFIVa4I6rm7++ynikWvLgNbmTppZfnF9TxCSkH7ykIa
V4b+1J5Dbg9qfGrm79YHrt9Piy0mUBWkJy+6ETmfJlTytJ3oaYedHYRwpVyrHXTUyDmRaL8ozXqA
rRPleg0JqgvkLidoXpPgRKLTuSWL6hhqfRv93v7nWb3kgVas28gpTvkZPMM57cBTir9ElwPrIqFD
IGYzVhs0EC8wxz1NPEvWFEWEsiIVdo2u9FppLp1yBPXEqCL/H6dQm/jEpC4mx2tu3Scqh7WF51Ho
TpyGWR70/YJ5gMabw+7BY1pnpYCcC/5M8UGRS+v/2drjZ+8dhrwxNT+tmXXVrBJ38l+GWMBi2h0p
O/Adb/j6jJakX878NhVuNc2Yc1tb5ucmLfaHuswdm1xiuriuUo5MJZKkjou5DdHq5kqvGcYF3yKg
D2n5pEDIx5EhqX3bc2BsY5RLUG5eY+mIo0E1pIhNAsQaNkb8sNVYg66JX3GwsSCLR7RYwolYmKlD
kYncGVT5mNNXck6kT7E4pehzoLhRkaPUYWhlP/GxTT6jJGJ4B3g4uLUClo2L8+JCDQ7nYfy1tCJP
r4V9qH/Uo2eT6J/zl0FP8ywp6fbkcWiD0rpHrtOCaUSHDDKE2RjnUqqXYZpo+G06GkXxCB35VSCE
i73DZReHKz0l8O4qHMD8OxbiCl8zwcBE7pnHA3lnAy6khgNjziNM+1fwsoxkYyvuziARSZKE17An
NpcjSKxPO24EKvgQmOBCeRPD4Y+qRohgqqTRwDS7zlLBqAOJOOz5J8a72qs/MCyt5xXDjeyIOLvP
Ago1D8/pNtFlG8fFgOvuL4oiTGMXNNlh5ZzWSZFHUHFiTah3gNwKc6RsqD9aaa08HvrZjtiBs+Qo
IB0+vM2Gn3Xst48ysafTRHoDUbaF9nbU2GzS36ebISAkf1cm3mmJL9qkVBnju0iXZTjOvr0bkzkZ
/Pf6L5XyCpa4mn9zHKywfzNb3mqZgAzhi91f33SzdypW1G5GfCmLz5to5aQPiVrlgNuG+Xvwke6q
/pI/rPfeCg80LXnhOtSZImea70MXnGdef9l+jsT6dGR/iX0Q/Fbi5nAFJYBu2en0l3SpweLnXGya
ycKzN8V8HPRiZgxZQTYOU2Hnim2ks3En4s8K3j3a/5vXwgkzIe4IryCGxt+pYXQzbjH8vceF5hAg
ZclpxZyB70+/Ej0AsYKHPoZXYUJGPQpczkujHe+iXPT0wsiA6j9qrF6wcyNAmQETAx1A/4eGPQr9
tteIr54FsUpxIcZ8jJq9uYwhv2O7sTgUQvBAz9BgLhdRt/CqkWiy0gZWa+5vKt/Vvg+9ONAPsod3
nYoduwd4JiT8YVrz8NtGxxZS+vGtY15InLJGnrDn63e3BhAB1zCRfp6bD90HNK7UoQAuWgS4iOIr
dYgls2RRzgBJtcvugrepZ0FwMyXkLysN0jwLGc6G1YHszcaM0INGwvNpbUsKMkhKfVGz8rXoZlCj
+kS10PPsjAd/2Ow0xZL8XIwURwnA9G2Dr5eFXTfMoh9kIytBhNJz5ARYYL16mJBOCZfryeX8OwrO
f6XMCItJmKJ0LctETY7JROu6canoZVsC6D5ZctY+cm0+pJruJvwu2RAdCxr65F4B1U4KSvh6DjN1
yKHYvENpDv9fQlrepEdMSs+uFOfvRah3ajAg1k738cdOKDrwnGrHavcldf/nEa8jB+7PBgioD9Yp
F5GiJIhU7n++V6aqhp2NcBt3RmQgS9ctSf84GD3NUpwFE6SJgsetr/BAGnNFsdQnp+1RAzjgiCLL
s+SebCtijrTdEOToe8TNzHaQYAllaiEpT5lxoyV1E8CwW+3Ul7FC3avTM5AhctCv5qXD0JzempIt
JnunelpSqqHrOaPXKC6krJiyMsOW22wYXC91tPHABFcC8xj8Exz7sZuyvWu/fFNJtJ7lgqvhZWGv
vf4mGNNSKm5BdzNF77rt8GJAT+5Yz+jdBAMa2iRYC+VEtQfJ3hBz7ocDcdZiJs2jR57YLf1l9BQh
9SXkR6z857qmoe4Eg3VWLYEau1+PkVBi2ZpZ2XNt1z5FlL00LeOeUIVDWSRWhjgWRJySX5ax6HZH
e8Ri09K1ozQtaOGA97oTKfdM/8sHSyyiE0pIQ+TTaikH0xHJxJoxiu6gcLZ4Gr7YRBbugMZ5venT
L+5dNhwnNuDESzt9yxlZhJSNvkLbSqsCKlCXB3d0ldE5909qALYsYBO/2rE80iIPRse1ar5mfOen
wnYudvMeNhbg3HU6lN5/hWAo+o6cRcN0qPwVzt9pbEkkVQ5nYzPIHwRuUUq9YXzQX0V2VdGDItSP
WN8sgGl6a+w0LGz8VVjTBSXk1foTRnzw1weeweElAryxGeY5wtmCsecuPIIEA4+azPYSrHlTy/4h
6qG+eVIwYCQpONpJjA8CkA1FSpf6Lv+VS2nlsF+OknNQ0QdHDvWud99b5o2LUYOrkkX6MZqaAfmB
Lr4s9KxaRaT/6yescHRTZnUAw6PFAlyy7bXfh87nC1hP6bPsB9/Vk8F/87TiIXPLosxmxBgpE6gZ
tJktoA5ZlG3At+c15cAtiFF77B2vYWxEgf2pJMvnF/+nwKmTeNanniloYTDo+Sddk8GaDaRsIKEp
NHWDmIc6zM7S+0pgtIvzrZRFAHFTA8DYe23efPwla7iNnmQa7h8rlWZnAaw15IXNgIKjMqX4whhm
9C2arhElwqObPMkeS83mzcFJn8c3m1zPWZdAzU0M7V12yAT3CfZNJnU3w2dUGilEVHY/q6xhlLsd
iPSA/EN2DhXmPGfV2LlYaFrnCfN6bozg230ry36qv0iV0gCBB8s6PHG1ukjrjlPbsfquvPUeu+SF
tKYFveyAO9LWA/rCeWylJe3zyzLrs1/C+7UneeSS/UkD4/DMrAIiFeRFTxBKxzbM1OGhA3vcwmu4
I0meSqTSw1pLAdPrPz8uaK9DaqObvJagd2Bjy8rxXqQ5ijeTveWcFO2ktaWkPgxPGAcbFLBtQbyU
HNCzkKRSRuYlqxBXZ8FI8Cx63Tr9b/8VqmUK+IBb8/Cyg1GLxQlv01nY9czVpgXKGGtWdugOo2l6
ZAkIHUFzS8dO/VAUwBIexErkrLEOVkosAE9RPmh+s1iOVdPFdtMIFi59N75Xp2aXI0kpZDJtknwy
T1SqB8zpztXX4ORUtoc2e/bQayaoBamhDup2E1rmJRTt2O2ng6lmE6Zh7q0OcUTN2aHWwcjxoYcy
cqpznNDnzbwzYr5kp2HcfbrFdg1c+Wa5WiijqchF7Fp83zhLrNNtNAfPtNIHl6SBI62Pqde68Scf
hJXfkHBiFprJM8kZhtHG+jrJ1jXZyHMshJPx/2CkfosuijkdaZMNDYRxCRJnh7fsuwNTXR2qpGar
xikLBHOn/EQy2Og7CICneSb8n1fbkvHXzvylF7hKpdGJyZHAJkAvmxBYziatWZ+YwOw1Wa94lunu
fHknauJH8p/GhIR80ln4WcpPVy1rDfFE9coPNOQOZtq418YrQhyXjh4mAsa1yjQoYb2Xh+AJsWZv
MZ8BbTwv6qUcNfhD+mOoDhqysQr6jPRNb+8gim51Q2YCLDAj28TqJob60p2S7GbmjUOm2tzO4qvW
RsZSHFpTSxIwRfxindgo63hP0ZPO0CrZqx35RCHRZThOsyTFYSpEjTeQaUyRTtR8PEeWI3GHLV+w
EcwEtzw1PUPAXG6p5qIa7lR83/ZUGrUatPXjU8rvWYokQSzdwqP9tbjUYDLFkhLg9zWG8AHh2Tpp
TSMSz8ZqyLbS2siNVF0ez98eyygN6J6MRdwyqIncFdx05Z11GwFMETiMskTnJ+RftFtqq5/BAH0Z
TBmVlWq24BsVhxekJ9dtxL0r82+/GnV8f6MUX+RA4tKpfwjmeNixL1cXdKyQ/OgP2YRdjf1rYXNA
dxqxjEsTnFRFO//el8UiuPLFebUjOfzAjweWYY9JoQtQGrJFOahMGOR981jxTGpJT8auEdtcCm1Z
qIBWp+Kv2cb/eLrFO/YXZojdKGSKfAvQvpXxOBVnc5ybleYxtp1oFO5B5HaJRcreuNBfhEUW0Goi
tvt+nHmEQdkiGOiNsQxq5ARbLOZGW7hBbPEhczNEYkxvTE+mO1qWlfHIliSRDKlKVBXi6YziG0mn
WU+ZKhDhdB/+ACxd5n0AcMl3ErCwyxqZuLTXOpsjJ+XyEjjOXQZZJevk/tkqTgdyIPoPLp/7uKEK
iFjsWBPvHo7sOWUGwyeiNVAXhP7vWuqwR9aEe3xPDfTnQ414dZThD2rpvhsaWiwfcDFnfSUtGdNb
UXTuSikc//ICF75WQcdoadZ/whlj+mZpzOqZaZhFwqKdfFMfl/GHIQAp+tZ6WxIxkbUzK5RvYjsW
qjuDC2dRZ2U86Ttn2JpwZl2+az2OgIz+Cr6DHiUhX6v2FymSeqraPKfeLONwcRR4gOY7xn0qKwwA
19x2g4YASwYL9Admll8We9J2VlNbPr9CHNJBub8hv3e3n5l0b84WEAmsO2+1axsmHXLyygdrTfnH
oEZ7xKHUrqu6DoEO5ErJP9j0CbuufNNC/vXDN33UGGnOQ/TnCKOEK0/aguQOwMPqzXDxNXevTUeN
OWlxQH8ByzkBEAD3q13UQw9KGEwwM7uh6437qNr9xK2YjR3S9GuwGMNyLB7yHUHWJJAHbVoyGfcj
NzzMvgYJQd7JWo3gAE0WxCIOIrY1wjYKYjZrjCOyZlr1+ITO46YDTJzW11NAUZfrQNSzKuN2fwhn
WMYa0AyF1tZNsuycBR9xkwhhnEk6rB8f6DvpUqXpxmuwbFynNN6Hk3qjnAIKiagmCjOJsy4nJZDv
xtbRS87NlD3BSHyL4YWh63zaRU2NDJZuO3yJhYWFPQ9JzITlqEAw1rAftHEdW8bkfGJvemm5XbAa
z9JBZitNcz1aLN2h1b8lJ7Srdzxl87zz61xCe7rKeRm+jka4unyDGlDdnPYoiulBineL+X1r6oIw
i5wRQRWR2ly+DPQq4GR8PVFmoAoDfQdp8/XdkA0M0RTzv1ijfv6zOfZjimoRdsIL4ipxtAiwwNLi
WyVMMAYA8+bVsAL66KfW/oC470kI8rL4E4McAn44hf+aUHPQqBppS7yUxzjEoOdjzrluFXX1AEl8
Z+sub5o3S8/AtnUpN9pDkaXkVSGunW3Qq9R+4IzmSHtkaK627aPPjYvnBe7nS38YqHa63sYbuKEP
sc1ra7ZfGcAR8rHliUrnlNaRoJdAKlCwPXTQz/ufWytOI0WE1WwNYvh6N0unRAGM482z1bXa05Gz
kJ+KdlOrjsT80p7JhOn48IUYZ6RHJraZ+xIppMnQZ3xKD0W1lUlg7hPeb95j+ADzHwgqBHgU/RCT
DSs5f2+ZhHJZA/5fOlcJ8Nz7KAJRkiFejgA9WFhNs2/TBJszmIcq9XLl4ji+55GscUFg/g1xf1mo
ZY+fIxP0R+t3CP+tFDEeWkpALA0WfMXlm2gI/po9b02AfFHLZ3Mn0IkQ0k40slLAYNKyCTpDGwxW
rlXc+inaSR0ZVJDqigIME54ITcrjil1KlIZLlDERQjvOuAeLBRPHWmru/bHXeWXc2MAyYyYIiFeD
gWcGnN04VdVuXTBMNwWySoRXwgODeXtAf7BjpNpGBwdPouU2VAgvp94/91IrZjHtF+hH8qx+4XGY
MxAvzL+i+xJrdcGZQ1fY4cFmKTrbmxxEOOWJb5MXjH6QAz9YpuDfD74klb4c0JFqf2PZsc8e5ElR
gzy8HqBsmrTypDBGS3U5xCY7zAmWsKZD7xHfHhWBOIAmw7KSUNxmvAo/v7+zSCIHX99eQDVO2Zla
wK5HxOLkbCy0ptcewUf6Sm7y2rZCARra8hxuSjcRKemAU8iM6gp4lclwYVYHcp1mdCONbfHuNTDI
VZQS+tlxsXdo1EndZJCHl45klos54fHTgRVVOE0Wc5VQjwuvKUAKfZp41KfZ+Tph7T7H4UR4Pyt4
t1fFC8UFpQk8p08DCSHXBH6X4RUy/ePVsFGOFIm25ovuHxZnylgOpeZ4oANuln5heOWGTHaEo9Nl
E1aaAzi44xGRZutfql/GkrSZL2+k9o5/aidBAGSNfd0yKl6sss+2p6KYIZ/OeIPowNTmeNSv2+4w
dg0ITYfbFAf1XS6+VoEYwnDj8X4FYUJ5fAqgIfG74gED9cvTnxmYF8CGmdSXW9byCmeTGHrKejfd
7rsYSQQaEZwlUGGpmDKlJILXUwfyp1zs3fSv63GnVyivjnQ2IYArWnoZOBEWBaFgPpUUIgq017wG
wd2lbNaEyZv79/kr5fHo6lZbPgq/VV/kcOU2NGBrI1HKBLSwhQST0NHZag/B4/RHBMkzBcF/xp65
K2SD2waGOqkDcEsP7U/pR1+1na4vjTWY05qX/GBh5skSLzuS5Po1U2oCpbol/pjF9vM0W8094MIP
ppQ+iraAqDDbtecHbDZjTQSYmMbIzjT0+2SGhAEfqgE41hbb695cdB+1xR8ooIYBKBXHy8fvMf58
W/qNKpcrcBd0IXnIBc1qyfOUBtO3yZeqDnd+dpMRFxjgWyU8lbhklYP8RIu1dv7UD8FNpXiFfLQA
zi6VZTFjfcbganoeqbBmy4bxtG0+0UyRjFm6ojRogJ8uthMR0lV6TGeZ5l4tHbACQDEGs6qv6iis
4KoanzPXcYMkaJZYQBbiqV+uwXLyAJngPI8Rlw2HGiyY5qF9oXt31p2Hc8yWzIkQ8/J2d6IuOPN2
BQceHnqs02z67wIqogo70/52x0lRBjroeAe6cEIO5x0oxiLJQSZnUR/G0cUOc7gCe3OOWziwHTTB
xyPnLx4LpS/Ez3l/12LE/tVz0R47znoZxhWLNHrRveNnW4aH2kAfCn3q9HoaG7yoBh73kF6i6v54
zG7H4/VSYHcOZc60erAZwODrhA5ExB4ykCg6BoF6i7rBESerJ6IJpqwgIYjmr/TJn/UQmk+DILJq
21u5xYB2mS0qI5H3A+a3Ym93Xdv14p81cTL2ZKs0pMhXLuoXzjFEB8ESlsOHcUUn9+mU4sT4lCdN
6VEQ07E6O07eI4bjftPpKmDazeFaH7ghWXaxdTHQe01xmbSmuw+6Ul79gpHLRCM5pk/yBQ4h0JMf
1TdXU4bljySVaHtEX2633f9bHq6JBUDKjByB7eQxi8eNAP5c5Kw2cdMYWy3qlLTs2Wa2tZDVs/7w
mEhtc3g3/+Bovhm4XSxKIbVi25vBGKyj/X0u5lDGOnl0CjQ6K2ZpUx+mSre6iLXvQUAWcIhKZYRh
8R5TLSxPDkwPqEMhPUzNsUuPvz6qOqfLWYtxKGvGjd8bG+M1XBxB5Y6PqylC/KnbZHMUgQuYOKXZ
mkYYYQMoE+o+BPq3TZYEV/8c+EXK1XFqGEE7ybpmk/+vnCaMLZjWtRTC8qH/PQs/ytAJsP5YSAzl
FlFzAnuIixKuezBgGsstAsJV5/WSJPO3X1iq0dl/4NrY9qvJAPrxACy9oqW1zi+xwjqPKcMxWEsz
3pNpGtALCRXrfcrsHhJXa1ggAmt9ZEitDSifDAdgoB9FYcBD4sgbaqE2xf9jQZ+zDkN8s7v+NB4+
veUXKhr8u2tW2/9hF/8Uq5jiHW1URwTm8YNPTVA2ZkbLXxVK5mOuXsnwY8YSF/9G4pEmntLuBEDW
7vrhe+q9foqQerCU9CXv4i+fPd5s5Qxcgrazl9opBx7Ig37vg2NkXHqf/9I3YLSY4RkIrig+sYcn
oqC3cxCvHCw0oD5q/kf/j8OrTKDxiIIXkB0D61EH7TUZI7AJNuzn265BSULoomk9lJ1b/i1XbESc
bn4mZ2DgXpzhaXjQH/3ttjAjlh/Bt5I09lBWl0vJVSUBnEE2NrCSVmUbdFNaVuVc9sAc/EaHg0rr
wQ7OC3rvZ/2B3kQ5Qvl7YUeB4BceU5Fj2aq7Vz5Z3geGksICncFYqeTYvwwa+trktmilZA0Z3kXp
aoLdaDXga9EgZpOODIeVeS2TkcXhr1oeTly0qvlTXXqzMD53LSBFSVlZynlqCwI29ccALthOl2Ak
HYB9Hu1QUXKiSMmcNJmtdGAxhQfdQtGoM7hjek4uhXpXaGVdXbJywn3cuoVItqfV8LqGywLoQ/9+
f4bIm2wd8pmpP83u73mRwie68eBQhZlDGxkmHInhlkip5sLARjfBnIcQY4vwzP889IllksdeVbrp
symvWhKz5M4QukyyZ+TuKmeNSn+YT7MycUYod9BTLBtf1nDuK0acQZsDbf3VHrHx0JI7PIgu4oMY
LLzFzUx6fX4Jfbqg3LUrS9LYCRVeAOaTaiNDm3iAZp3CzdaJz6VuKP77ulHnHQcMx2clzO18Z7Eo
g875QhnbPN90GHTV9oP30obKw4/N0Kdfai6pHheLLEPho/kZPbacIgDpIxlCII2AeygdCySZh3Z7
NcYNQgvNZKTQClL2Jo/bey0pupRtt/Nz3H9cO1/k+Qf4EdMf/KUGwzZjmLbULk6f+USJNSmurr5n
3vzpf3mz5iG7M049eux+DfKQ2Ypqg2/EkYHGqyTPRKyuE38v1S7OSs3mssPVPczexZHRjC6cXkKI
pFPdz/SR3gMLtY5UDvHjNnYurmsErXt8KemymuNRLkzbuCXAO5CcnZ06l7dvpQhj5Qj6J5explpD
PP5vKugcZnKYDBZGNEo/W7QaNMCfwcnI9SIOVd3jNascxohU/X/e4D+DLy9f1w/7V2nPyW8/x/nh
ruDCZGebI9MK2dfzO43wtseO+rpfv+6IyKTrMiJPEc75WFAKleTm5x8UL5+7O2Kc1BGASH4+E7gt
T9CakXqPMiENx7QD2CEAhqhnqPGyuE0yixwVhdl4GF2GlTG9aXKdRusEr3ZnLn4LjPrFRz7JLGf1
R+diQ4oM2+El2tjDBvjNKl67pXiUeBg8s00GIHRvqKbYKn/+FsI4NTSGkjZbdNkeqfPjL7kBKmld
XSpnIuaN7mXhXqfwNPlZTSbqtdzoEdUIFDc421K88VaGyETRwLxp6sy3mI2lOvbRP0rISYkVGmD6
7Zxy73asGjL14gPY9wl8VpO9omb+KRBiqvDWfLELlmZGAYi8Kx4xPUUAocrb4FODxZVKB0CCYuwa
CuEfVT5RCuY9be3vy0lAh0MNPfuIcHYzy1LuapfaQjqsFoRjnuPGsCBjT8YrJN4Vy1dNph1AeGVo
7qujhmbLUsKciIHRmA9bupihabAcXPNCxlcNVbxXeYTvut/tInyt4bDJnBJ4rCENT31A1VTxLqO6
/ZAdjxp1pzM/8E8wIqpfLicEhnQJn1tHTRjmA/EO08CCpfr7ZcKjDvtFttGR/XKbw8qtYK/I1Ddn
X1V66qDJaX4IzNPsWddLFRaxtUzJ3YqxbW2zYjENElPD2pe5p084hTXU9/EFwdvqjQeI29ijzmC2
ESPeNzxlM2G8sDQBuDjaHHnj/X0oMP04kMQhm0VKKDuGt80C0bfB06KCzjlAsZ3APYeHT+wn0dzL
C7vPWWJd+38tngvQvuDRAHCkcs1pg3nv7q8zvXWcpcj4VE46nTuyFOCZSQ8J2AiemzQ989rzCDDP
jUtA38mQfWehH9fpL6k2Twk0Pco/Vujcsyq+a0sAoYDD28Xm9hd7DMFHbIZHT5dJqSHoYTaQawdL
o2ly/rjNbUB7PWQikiKpEUtylasbwUa95tX2hYY6D3A/0rZDLPZZG9Da0AeS8SpzgklGZzLAdJ0E
CsME0Zg7ZPm82U/t2dRmHVqpI4O3rw8YOtaxyvPXugTGeIWoQfySnOU/JPTxIkODhz0S7ybcTQXv
6W9fN2wXTgTP65q1F2xKSZYKRmjZv1IwCjY75qub3Ck+2tOefu69uBm5STw1RMnrome1NBMa4Ug/
ZgVem1NyAGTwtvztV4I2wMTJ2eXOajyqw4jfQDE5uHjMWt9pSSO69UZMD6ofynStPbBNQE9kPIDb
h+H67OFV62wqgXeAd/cuAqZO363WgF24GTdD4zK0ohn4RtB1zMMwMljONzaJTnlS/ezKNfimnYQz
ebWvu7Kma0DF7L4i2O9pg8as0GeMkLT2KVGfAE1PdrXEdE7ucYiFcnkujksLYiIwARyDj+pDix1w
ej+s2pLh+UxelBEIqBIQHfUgQDb8X9TCkn3c+FwNxDLxE4jXNYfd4h2Lhw87RTwLQZ+kN4Hrscwu
f0M8IwXHJaqhBwx9DS5rQVFp2ibRhvB0pypN+nwmkvBsvLfn8YkMcOLqN0yLqkVKlZW6RWPJeZ2x
NFFv0+NSZqA92FcbnaFkgz8HYZlCb0+eVi/waRkFLOMcHUY3iyDQvSTDtsh2WPASpnoMtI/gQdQs
OjVZ1pYOwcIExlTCvBXBw5lOX9mcpSu1cGQzWQKABr0OA1wugGEv2E7R7MHN4hpk0FEaGFrI3Z/d
XCJQinwNdZFReyaBeIUxlWBrwRGKpCfeARrSL11GTLaMBJ3tns2inGPCdXGZ+PGiaqaUJBeWpBM/
R0f1WhgQ6TZsVvxaS6q6ysVR06HOGKyBP6eZJhTq41QkpdL8aR+1WM5b3F+sBo2i3XD7G7GOQgjr
9j+XRjelAWV5EZz/2/MQnQo6M5RF1UVNIQmu3vbQD/fjuD+fmWyd9a2TfCPgsxlsf8uY7fUawkJ6
Ao8fbNoFTaecW3HcRmQ05417rYHxlf3PphcUHP8ARl6Rx8g1zm1rp/o7918PQRBP0uWcGdmQlEwG
fDM25WjnCJVmp8UsMhTN4Suyk75k3NXyXT9YSQh5bl9FBzazsblRCwpssqFYdiS7uZWWAGRVx+gB
Dr0yRSzu3GfS8fh5Zpp08DVfuBwWLl5EA3hW7oe+QitO1pcqdF2fEsiiTwW0Fr8JZt4oSx09O5g2
cRzxpDe8biXDybWteRg0M99RxzfUEfcwVVsy6muxyvYRKCgSeWF0O8HsJ7K+JiNyg+egQV/5fx2H
KWGzDoeuAYwKDq4T5WcGukCDC6S83bCZzuqDNgswN/OysVghf347K9pWSST7cPgh/eRsDKk8V93g
WcNKRbqMi8MzEOfosZ7YhtjpfEkosp4BfppkrSOfuiaHw83NgHQJA/M5PgTFtsthwS8syPipTkEd
Mf3ogXa/dHUhubKjLpYh1zd8Zeosqa+8VqQxOsCP+vjGa2dzEuOFZ2Nk/HWuWmwmSEutkKB/gbtN
VkZflIf451PVxPyjmS9mz3rI58sTgqIIkluNXPonns3xrohG4ib7r/6/MfN1XsKhrUzLx1iBe9NO
fAX4Nh5vFBisK4MqXIjYnYbtFUyKD3vIvzPpcbmv+xeXtBQs7MduU5MLAFuXNOa1gDOvN6oT/fuI
zky+0+kiiliOM5CcLD3xKpiGorYLdKrJ4QsuYH6EIIbvROKW0z0mHijOgHLBtbFElEViwmA4nXFt
vZxGcH/w0sU2ixbnqw2zvm7ohSFgwkxn1SLrFQpiCLOqb/hvo9EIS4Yb6V0rSMlW0UExmhAV2bp3
fYiFBdyxT+q2uwA3livVBiI6xFbP002od5jTjnAJGByUeRj25vKBptCxrZr3xiOQbgFkT6EuhKGt
Pkc2EEb8xWt0IEdecGExO3Hhjdlw6n9uCqfG2yOY2uA+4q5LV5jis6Ghcd3nYT21q9Qj2rwi8voO
nyNzR2xyspNm3NZxhfGIw+6AgzKqhx5T5vLLDYNPF8ppI34Gf6Xv7yFTYEayXZ6gsZudoTY4+OST
xANvkgIwv9Qb7Zd4U12fh09Z0eyu560DTCYy/YkXnru2DfwI39DA+REeflY5oHZ0eRtoK1j6cr/f
GjiwaBa8eWB2nJ5AuTNCd9ripA0UzWILd6uhpEIMwRoTQulCi64pIn/0aqik12mxa2rXcDAVu1xX
506b6Tgk/rznmkCRRdasjzKfbzll+NSU1nelE1D1gGNBonIjqHfwIUMtd9PI//e/OHDjR4EY3MbB
A++D3KWJZMRbOewSb7rGP+GVRJFVZ0zdGhOikaKKx1d+uQ2QDp2slHUwhN6WFjF6FgBg+RQvY1ED
caNgMN2IiMeqoRQ/Nhzru/HWxa/H47ugJsAOe5sjDzTSDN6Jv3XFhSzJCZt56tG1liZKL3ZmFc3+
DQmbl9+w8OLU4y85OputZaWFDqGVcFcamaDOKaQCAXnjktkQLbaOICHRAtQ0BnJwKnz4CUrzfZNq
wjV0u3ebQfXSnUL/2O6AMDVKs2KcJxgM63IuCrnkY+jioFM1mWrC+Art1iSdZh7aNjlQzfey0N56
N7HRF3zqTnXnx5pY3tOsfnCwUTBBcD9mjwHeQkU596DC/uTfDjs3iL6TTejW1vy7jdT5eAJy78gV
jDFh1MPLLqAPMqcTSKuMC3DcOF2AniG0k0ewiiwx0fWf/DIk+t96B5p8LdaVUZHxqooa4Xnkv6Cq
a+hnvsy6DXeIFKv7fLAYC3r/VRUKTU5njY5OprqQ6O8qb9OeC8qFaHOgVDJEaJMYsTBezLDjqxnG
s7VIiWWiSHQ+EAI9hsGgDaXh1Od3Dnz7XSss4LgQOA9FpjPeVggWd8GK43HrNA/HPbGJ44DUHRWM
MBPsaDhPjlvc4nVLBrUPIkmfv9v4nDNTrYu0iomTREKDDXYHH8iUyn5MuitaxAk71yW+kYFhaibs
F8RFy+CSLODT341qZRNdD8aPIiOOTicmf2jVFY87RfccjjpLWGyZdD94jfb9LrphjJxKce+5qTdn
eUBBw0rHDEOwifDRfHermiVrK7g1JIf3oHt7IpX60Svjc38DhbwnC6oIxqXqcflgX3ymm4e9GiTI
eU3bw79FlRvq3itjWushvLBrSUniFPoV/x4hr3nAsgale6lAFbLH9sYbhDG8XhBF5GFY0uzxajtH
6pXIkP3KWVFWvZfGfSuMQC3oXRrZq7RIQy7cxXiDrpcfT/9uDWwsO3JOXjBuUWSVKHSjhDX7ZbuB
bDgL+LtUfoULdsHtsJefihtJMpDRwJ69cfuNJy8M9lgqOafMNEKhtpLjlqAVY4BTJYrMxcwFDT+M
LqynLm8LQAKJaAZF/Y9qLCwiJ8Hsz1GDeh4DEisIRJJ6z6/cv8lo/PaN88vm9Ez81DlmueeCnYeK
dbsnmhj8UKpRijnT4selfEZmDEudM+cm4jRMtrUT/rJBJu9BeNxlbTsxm/eLCzXE+l0UuLBxUNl4
OVkxihfqnVTOPqz+0qY7GjSyanJnXLXJVvABPqsPWVaF+/41nrKy7rm3sxt3Ycbx1Hngv0nfywqG
1b07v/dB366wUsPwmg0ovt3iiby3IxiOyAfYiDpU296cOYJLD0sFmZLtxe9pBdB77H9x5K0jXB9y
iRIKO467Z5CK4T90RV91f7s2DukIZSwqxzcLhHF20WZXErxab/+vHrXXL/PdFJShRWYsBZTQeNAx
pxJpiZxV/K1jVHyGmvTN4m4nDxNCOnWcpVI3YcQaDo+OzrCwc2yzl9xaVFby/L82vvsuXbwXNEgM
YZfqN6+j4uVEj0Oe/QurvbJRnFIlsHuDHZZoeWr3R9L4rGDuAHu9B8S0apc8nWL+E3CqEJOWIKHN
TW99Qt0z//S8xclAKEmaPm2pL6ppA/SxTTPw4c6RKWupusjUQsdH5T5Q12XE5Wvs8C57B5LRB0ji
DPm/Ra7oIsSZWFCLAnPtQwDErnVHvDzA5qTdscfjrKRLtn8Ynuwz2sP1qU43I1+IXcSd56HVVCaN
27s2rfLKfcoHY64H1+JcPCwrkV7jXWq/s00Df74NPHiRFi2yde47mHsUIIYGj+DToMLxzo+N9dU9
mom73ORvdEngFJ6qLJe0ce6xqzBmIeY0pqkLx0Kd9rn3qLjaFitNz7kUJJvIiPbzzkOdO6TxLW/z
XX7TOcfUDPu2x0flOlJF7TMXU1Ps7pkU/I8Ds6670nhAG1UjvPvE2HWprW6kfrVlH0YPe+23lTKG
L49pqjeiShoUCTD9LxUi8z7djNp4bEVIHFV4pRXNkNjzxaxkGQ3sYuTBOS/FpXNBoYDAx3cerZdc
9CYXTyIuqPrpBW+nbJK8tv+RAeQ/JJ8dDlw2Mef0OXeBBKT5AAVdAWdHTV9H3YRJ3207nJf76uyg
8f9TxMR1PBUBs64y9tQFI+zVWIKFNG4vO71SefWDMgYF4e6S7yt8KqCNEkJDlqkyGiiDC5yRgrkd
iw1765rT58onTwQWaTFFwjlu//QrOKJCOmPSGboV2G6vt7pmqLt6oBHX6ygPl+IHBb3z5ASu+eTJ
sNsjPzn8rQ15n1uLkujbjbk3fjwGNu7pCNgsQ1C+bjkYK1h/XdH/hj5eYmzYRPf1RDJX4MWx6AGo
q9tMpkFI0KswKQSbrddcGzJP3hHhJlMW39Ch2oZsPSUL+nNqGY6zeOlRHR8Eq4zsuAb3f5UlqqF+
dAU0r84LMT8Ai7nSkV2DMt0wHpXaGGllSe8Vt69fCp0ojIYmg0OKvHMWfKZnAGJIMZCe1lvg5Dxf
8A/BEGBrbt20smgfyRHHFR8/UdOvU1/72+8lJrFHPcPLtWUuFkH2jdi3oYGGI+w9zaQ9KoebsJaw
129kU+1YOT7BttMNi099D2FGyQdKjYWfXhGf+vpC8LVo8+VBarEK5Udk8Ex7f1/i3uTba+FbaVHS
ugMQ4Ev73vlXRgWsTAFHh4Fw2F5Nl39jn+PAO6CnN4MRKzWOq1lI+QoSiFbWCxRuE++M0UzVNswo
J23Gn4F/YhclUqiFhmVXa2X7OcoOhYu4rWh2bcHpmlXt/Ec+mKqZuPPCrYGTdhu1BHd9CfD1dKSl
PQ65DJKRKRzUKrf3OYUMi6zk1nfuvpv4sVMLGr8tDSFLnDXaHV7GGmgTCGBHafjr9ZNf41rn3sU8
/ngIB4t8VpAPn/Md6GDobVWFp060Fp97AiUPXwDGzg2cAMVhYrFagROsPYDMX59Vim1UjlSLtd0A
chnxtHPZkE21zEa2gSWh6HL0kruOU35cHJoealCajxtk5u+obrQPK8qFWrKNGIEGLZAmQIKr+Ex4
+8MY+uuDtAnhFxfAGWegMOxcWMU+m2DZQ83+L0A9QHVbZ9UL6jFXShX2bP4YTsWw4chtfVhaxj0H
9/3oGFYv5bRucu90TT2c9V7stK+VV1zpo+h29QDm7TaRHf052pig9iI60zDZ93R1xUxRhfSB0hiB
lvReLLONAVf0wv/IeW5T5RwPIQl1O7ITL0udxCATqcrJnshITTpz69gEDAi0HNrLAu37L6kI/FEi
S9gqQsTEVXB+lb4yH3lbr5cufQuqWVVpuo127tqslEM1PHHwy4NMSs9Tf0Yp2qezWcY381lcEU/B
wML5why8OGb7uO3wjYnK1q8LT9WpU8IjCIxuYNBoDDIwBLiqcB4ubQvoeGgiP1nC8wAoblOY01Y+
IC/DIAg+19r7Nv8jY2HaeE9ZDN31HxuDMGjI9Yslp5KPzvaxLSPY1mE5m+Yomll72j4Pe5R3nORu
q0SlNl1U1Gvv5WTLwEFqsmyYW9go9hwkblxctK1OEr5uZuUItaCteNPdkJFmnwnq4v8yMXkf3QoG
Btv2NsXiK/9LSX2Wt2qyT5lrTknD25R0U5Wu/3VoBPDNvutVrJ5LHavbESZlI18VcKJJ4Of6TzD+
J4fHwpl0gdwMJz0X9of0xT9M0JaMQZnSh8gIauEZx1G66uSmLuV27C7JSlnRpjMLRuY98WJxJrT9
1qeAaC5vFuMAf2NsjBudOTuQ2sX9ajTz30F4U8cpcfEFhNZ8K5YLdLwxDASVxJx6arVNSOHfTOzQ
yqw76tUF/9SFzG8+hIGxw3P5QVQjkymbLQmeQdBdUzzWV9wMrF3t0sS1bvYH36Lu+9kvTHOdgjo7
DJEUVzGyKig7TQstXJ4NxDeNiNOiBURms+zXaME9rNUc/tCQSp/AHVgCc96fjQSaDETjZ18lG/q8
3UBLQItdbI2I/ZifI8segO2d2+ivrtzOof2JYtcAzp6t076BMc02rGMAMOvxiKY26xE9qoDWsXTG
On9PqWMg2xNl0pli0qghBdQ7xqwO+VF23P6s8Bj0lnxu47St7W/bgZzFsUAW2/PNDfiMA/PKbHF6
YpXB4Naple7tF8UcuVEFRqw1HkWqf50+8t5GOqKfoL0jG9W/2EKJPi+DBDsRgF31IMXETjbe3/Iy
uv9Hq6+7M+KwFQ3PSh58fP045j99BcUrUiuNj1/r1a/6tUpt4zDVxxj2xp0MOzmrCX0eMlj30ul1
ReBF+KINjrM0KLkG7v5Mtl5b3Qak/nKnrIUcBRg7g4DtwPbXcvbs3lVTMIOtaCLmrMRRWwNLXuDj
jvBU5lI31G3qz5C1lxf6jEkZssvfw4/mP3zPgdLw4FZ4iTR9kxRJtrv5akYxW56AThVQ1DbYsHv2
0f7+R6pRJziJ5UmeVpfjHCYIjwe8oEc2/pdS/QViw9l3z//7AhmvRxs5IPIhBC0ERQ69Arx3MHLE
aRjPa4jcLpfmt3XVlDcWaCROKxcWqQrhynTSYN/4GgD0tweyrvSKopHAMn6G3YwuP5KMGN/WxLfv
FIOvXTyOrNWXxirTcJyCxY+zJ6ZXngsg8l9dByy1kIVZT7LPzHAfUGWPX/M2g6LUp39AKXOrliMv
vpATgY1YHEyWa1oy0e87g55VtXhDo29Lv9iQQbHv8S9TREmQ2aDSOT0Z+pbLaWbVZ6lYLLf+6fqa
rrhfMkZnQZhOmdDB9+hSzBvb0NnRIa8kkrRIekjAvcgY3+11V3ZcfSNMQsjwyt+/MCCh7gRkrqtx
RpysBaKtkcTn1RR2k9VMNR6atk8iM9qbDWzQZi9yz2hwVCL16exg+o2Gx4WGTng4upVfShuUoxJS
PAo9YJ0Gyq9maFwUtQysGG+hIZtjU2KjJbSOAbSp+TjZLUMxi2sDUE+zEzJ9D+7lyOSfYC/of+Lp
Y7f4w07JRjbx1cNFrbKZSsJnCiriakaQNVZ6qwqjcDIPnobF03OOv/MtsEwBdMo37OeY/2Q8+JM2
Xi35QCZpqPj9DO3woG5WhLQGZ/mYKkgFD+9mG+Y5cV93VZ/Aop42cp5VpQ8GPx3ytfXGruM+rB4k
GzLue0ELO/ypl2fWBxhFMAKN1LW4c5optc5ggPH3PNL9mQsXkniA5TA3WXchye+87oXP2nnKW+LN
NHaSch41jvEXYoJuBQVP5i02ZxbhlvhQPqjpBPYCi+vCHigqLInNt76ZnOzjGeXBrFOujXB8sKxk
13ulztgzWhoKiSaXFpDM2nRSc6RomEl46/Fn9S8pWm4PxDnCHH8+7IvYuBAsbCsEy0tOokTK6eP+
otXlCPQWZpgtVI9zFAbaQpWmG4vlNYxGmTNRtb+T9ngTdDTo585eHAJwA5dtrKqTeKRb2NMHoP32
v7pMsbzBF8LMoY7k9ZEWuV1UPwZjRmRXggcvjs4KT/6gnPYLOdQML7l021RKHAP+sU4gmCMzPw/f
1f/yWVStPQTH8GSx3hU6+9iBrwRB8SHonAUBLHP+ndFfVrSlt++ND3rMNoBewoohagOt5o86p1Dl
VzNUcHiP0vOjTMfDTmH6hi2bE7Y7AFxpV3X9sivct4Mb0LVLeTJfLmZTlpyNN7jZZDvSav65ecsh
7YoWrB/g/3PNUe7V/6/HYduau1Xsl+yks22STwVhEVSDasAaUrq2GX0PybESeVNoYRFF/lDQ7HTB
VWyeFx3VDxrWcq65320SoRJlLgHwy/U84A5W26S0Kg5H07Goz/cowqBZxqY9LFwv/ndhCbXR1dLX
aIRJxiP3GlSB7jGU7hmUidDI0YknLHwkSQXP6qmxy+TsvaMwfiFjomFA3a1cn8YTKca5jyEV5awo
898wLwmCNmO4c45FMcWqbdfxrict+LQU11tkyj5lbIuGkSQ6lZsay4a1R/CtbqUazDw9RP0LNSOC
KHjC3v7HSRk+OawLtwjCMZfaKcNKTTC8nrt2BmZ+rTWSajmkB2p9ZeRwI+0Lk4yvWimy8OVhML8N
8yLOxoBoVIHF/+y4XjQMIPuGxu5DDEQKw+mOY+vsdmSrIW5aXtu+szNCMqBR5BShevnivM1TBTNX
8INEN8OxVjWjaGdih2LOynBs4CP4Mi1LgcFQlLng6RZIL5/wJhd8oEYQcUx594V21dvYnXnJDjWa
k7bch5KvB5+bCsnnlCon7QxdNAjIyrFM5r4fJqhw+dVvbhex4GwCuC7plTxcFmfPNHxMS6UPJhaV
la6Fk9pOiLj79xZ6wFBunDnrMqJxA/jth87bciJ0I915y1IGA0E+LfGqbIFmyvBhuEPbM5nk/qpe
0+rp1VbOLY3ffxwyyHBjIIDi2hQzErbdeSwfRmlRiEmT9zu1s5/CBamFNQAR1YHkNWOtPQxl2OXg
efymS6S3zfKavg1+GM8Z3C4ddt7NtqIgBSnTqkAyuAF8qfLOkdhyU9+Lq2Ct0Kxnrq/1V6C8q2nc
821aKcpQyZHGiERoS7H2ORzXJv8z2L9dR4vFbQfgxsmA+5fMlSH1nWppF/XJbOrIJ3yxevXWDOft
ZIkA08cz3LemBcXLRWE069OTJfxuuT9pHnIqliXow/MpMAp/jd/wLl8oMDJQTYZ1B7FaLpP2ox0v
2sManczMcsXMx8JueUDUVQ0TXDL9bxcNySG4KTy/RaY2PiiBolN8mR3VmO3fyYZvcWRLFJJPvyjX
fsF74X7YFSePO6VdzqzS4R5L2DfiXA1moO8wPnTRLSCWpOmFRzbG5rkk9C4vfn6EN0CEybxaOtMT
fipG3pkNlU8GeWM3IRM7zXGpkq3fCpiC3FtO+dOYKQFZylY757e6GfyoEMXm/EzQVdsEb+N3Oifu
CpFZ9u/IdQhpg+xncgsbp68B5sdUquo6PWBNI/YOLkm/4JnMy/377SdHIdyPaUYe7RNZGJ+/z9UZ
FIZAuRufeqTdmXFb1X5J/XrcU7M1XavSglXPq3zdTUE0pC2rZ88AYgmhT2U4s9Idk0DvEgp2nMaz
+uKRbNH64xMGd8XaR/0el5jHhbzNurc5TsiTKP+bSOSzXyub7/ej/SZCN99ziR5rUFX390dHzQN2
iumTtD2AplJR5JaFudFuaScUaTbbUpQInlS6jO2jxaic9wL2FGO3+uEnhe/bL57ABCMTgINpLE5f
RXTOH9d2N5NdvAJB4qa7JDTsy/e4OE3Q9M04eNeK5ligVIjizxtPeQj5pHvibFdkcB7aO0cstoxL
yyuyPndqYmiIpDJf8iOMwnoDgW00yoh7BTtle5MD2tBgdEfeKSFVL8IQT6G4+qwLOjBQfzFxf5o0
Lldl2BCCCi8eiyE7YkkIfsMhDUAglMdjdtMc9Ij/bdCyXu4f377TlIFhHHF0O0wmZt299vz5qR4y
VmL1mrIHQXdWBVNzCUQ8Syi1FxFJHiyD5hzzxMAfFArabTE96J01pkfSFTLMhH7OmRxZzZP5YedQ
vDFuLCosodEojI2v4jYz9HzuwYD1MO44gw71B7SnmKS6hDxnghJEvkNXeZBiebP97R4PS9ISgk3E
2j4rZ8zq7AHKKnTgHED5uelgQDvLNnykPa77/FH4am3GhRxF173wNlj2rctBkUiQtCqjMLxKUCmv
K5hWapBnokf+zQhmw1SLIJ4vVI9I/A735vDEQcQ6AiGa/fKtURh7ousxchtwR3gBwzjVDc1c8ZQ7
YUpeO1wJBCpBE5Irpl4EQRup401yVgu7UD3C/aIyWQvTfXoEnyTvC8yHuO/H2C7ZYD3VKSae0UyW
e1XQLaeHrdHFgZiNPMlSMfzNY2jd4A784dhNNCqo0mm55L2Jkt1VtBg9N4pGMoyWCWW22q+qnxL1
JkGSKcHO3WxcXgs7vzBbHhj15mVMXKygJ4K1hf7Eij4Y9TqmChYcroelhyMgmYTefcyvEvjIeU4H
qv8QzGkVmp3yymjX9JFQ8Wq/gWZU28mOGD9aOC5f2H0QzworoywpzJSDzC1dEMsi3/tohYfYW8CX
sUyMRF4CpXiGj7u51y7LFdKGqJCeetTjcUV40YHtfqasBY569IktU4N4xmoPEWwD39030vIgxhlm
4OfxnPbb3rzP4HHMpaXoAdYiye3hGU3s9tSqMH+DmkJPpvtn7rt0n8F0y1/t+wd6uYlOunHjM6R1
yjYPLKk87Q46i59UI18k0krEL/NmzkVmAGA4ZhDbJHhboxbTmbiFgv2fuSQF8ukHiZP69g4c8QXE
Vf0D97mBqriMOpxMb24r0BaAoKpPzA/4OAK6TU76MH3NpC06pn3zsGtMqeB93XUhEi5HOVLo4NFR
6h1IfbznwdmKxicA+7Ybi4WbZVqqdliCF8Bw9NXLhh5cM+68d3r66kFScJ1U79SrRAWlIZhJ2OOS
HUOx8zw2BJqol8L5U26GXGS6GoR2LhdtjsbznyV7isT1vvffugymfj3LuZZyY7OTA9eFWXu1DtwO
jccxYn3EE+oVopzeO3yaFaYEB9shsqonN/a+N9Ydnm41VW9bOKqWYMXUx7qacme6lJwAh0NySwjy
WVDKmL8tEAZaJBGh6hrIe6YTlXco118pWvicwbeUT5gS9TghmrXLOdYqpkuKDulnDeSjexJQYROF
FOB+Azu210YHnaPwivBKwqVxVGhJfbyarXUZTG2x94aUFoactzc077bNZn7RczgB3krtRqmo5GWi
JcpnDE2gq7y9gcw8fzFomUXil4HmfdZMMISS4tjXZOpnwjXzgvskOY7RVG4tNvu0DgFnrkGTjLlZ
jIndVaGbehsnEw0sQonA+baVekRRFleJ9k2qDdw61WgyTG4/1a0iXklX2UBiyL8O7z9zux84A294
NwxNe/wgSjiIAwNz+5cqY6tbFMTUouzqjvkvwzAB+EGshaNwZhmL0Uehob//zGmwo7FBSfQP/2Dh
xXgkfzmiECUpd2atjQsI+14VgXbrHtdViRSNJYIKhErIgdIXdDVMjmP4iaMddOTsRQjh0LNrS5j4
336nawnFCN32uyN12BW7I7Ua5Hb6ySMeZS62TRjYa+br6Q7rq+ZYLHWuEDeIVKTC4gus26GKyPWW
0TR2R3+q9hMDSds4irh6sl36k3icqww/7xgczlvMJY5htvJG1HWDym72LPawcBtWavJZRgu+oEi8
faRmtPOWeNnFTLlZ6VmppiISsBAl/Nkg3BHNm9xod/D0RMz7viOTXXTbfxuvfzZ26WQdYkniaNID
YwSCmAj16micWzDbx+rr4/WdUpdSzMxcQ9qkkCaRGKWQNm/vOM3MZ7hkpH/+ddKJiMTWWXHTSImJ
89nrw1x4k6EZv4PV1OPx1f0eUXl7hQDY0JPCM+l7OfxGHW/euVi/X8wTRBR6pRNsGiELlJOxztnm
V2ePSu/T7Y1C3VYP953Ms7V85DQLuBj2mPjvWLgw5NdMppaT2igrU+v5gqiCybSeRlDv2gEFDEoN
XYyq1bOBnkqi49jAIQwZ9qk7ZMUFhsic++A0eDhhHd5sA4WokXxnTkEGXsCInA/qz0V3YouVLHsk
o4d2rS8RUhTbDY1xmUO8frz8wNE1P/j43zaLcoR/PyJ9UEdNbwCwUiwoIL5LuWZhEe2njOHGv6zC
cuAChKwumNb+EG0SDgtbdfEMsA938WuENYgfalYXCJLuZpM4cWJzAjSCo4zkSeiQRDiJhopRT3Uh
jwcpcE1h1JCwf9GUmiR2vhUAHXMgkUsKKRw4lTiOtZgGvu748n8aQNDXwKjixQ1OgSXQoLJ9vZ7a
wexQF1huOMZA2j5mKcRKEYf7inC5Yf4m9EiyEK9ArtWmIEWmv+vXjrXRoo54Wgba0C5Gk9aebBeE
1jJANYP7WrVWreC7fLjQtR56xuSPcOZhxvpKh+h1Jpr1E0H7/gCKD/Ghid8TVbbR7ZgllLE2Anbz
wEPfn/XCr716T6xcRgLKakslyy1mCJgxklWVLzdHDTKGPphPnMrIu3vbPIa25lYPBWe9w20J1lfE
7P2H+jm2fsCjnbZd0yKqoDQkiNAKhlpH1Xeq/uCgHKgDIbhQoUKwdMSbbSEIZ+hIUetrupskzAtt
XVfb/mBgCo0/yTJPYmrJ4HVaYQgtGe/EGqoB18YcFu3A1/rnrjsCIKEsD2WLGiUTDHdaH3b19eDq
FHXiJlqJKQLZJgdist79FshBs3LTsmG4iraLX5j0r0hpsWaOTmdntzcMIYUF3A5tMhHb4il3q7Dy
n28YHj0Y+GqXgDGwX9ubfbb2zm84//fW3xwrneXDZ43+t6+QiMNlFD0/JJRY/D2xQMQH7PGFr1yN
iRyvGIZQNJd74LrURxC2MAoYvyyRAqhZGpVMURVjpRAIrzxhypGl5xG+1ZjN3M0tOe0+D1DD+RhT
PCtlWxzklmrSsQUC49HvNNlNUA7w9UbPxbctp/nRRV8kAF2bOyv82UTv3Hw0Tw6RpT7k+QwIRNzJ
U/o9ObtFuBWvO8Am+8B5VZd6zb5QJiof8SLKwHqz645GVtyNZWL/T4yVfuY8p9IwLsnI/JXmuBGU
EwL1zwHnIVB24WnBmQ6Q5++cZzQeW9si7DJV+oVYyGHTWdhAj/lJ4ujzUF8qMmPZ58hLJSNhm6Xl
2Pb7kZWiG+DuYDC72QMw92kQaQ0KWmN6wfZrlVjYi4jtP6hi8F9JW6x5Xea5CU2zdoWe2R2kyrNo
KdjR/2JuePLY++ZAa7g3/nyC+Fb4VZ1v+lBUTNbOt38IfT1IL1FUwEWzBdlhg9jxsLbCbZMG0yr9
CsMOSMuQTgDIq0N01w87vx0tb/fumEhuq7VfXr/i7opSX44Nho2auKKh07oiz0sw7M7iU5WGrI91
r0akDXBAPrSPx4ip7fF9WWdIzLhE01AxSn8FjrJIYb9nOpPebAShApr8196C9J5MgLUXGe+fNY+b
Gaa15NnLr/MRaCNR9P8NC2LnGumrgGjuOFPoAo8CUjL5OiWH6QsF6NFEl7LFDbEP09HeWYZrgFgV
a+xbVRk6r+EM/IDS2dShh1bz/WDXCmdu24ABFoPcWwhRV+DHGKwSM9PKtk+cWZyRLLVM/rHVmfxw
GqYxXBeqAF/kh1IuzjOgZ5b1PoS/CbjdmQpdOjcF350WC3qKS2L4vj1Ge/FiXh5mGXYUmmkBDmc+
VLlhxfOeb6ygWZDRPenl/lUIV00Es9pWlkRU2Uzq4Wtr+vzt8XNmBUIXLMWgR1bRYgBRTt1VhvLi
8V6wW3prpBQ4j1VU7zbROtLiBwp3iWIF11Z4aDSmx9VHQzYcX8Lx7xE/exJNRsfAjDKd9jANk1Nq
GJuzSFoSul5SVcp3dIAwgwn5CEVDmQ12rcN2e9O0KerLHmeDbnSLYnqRNt/AVHXy9wZS1kBRp9jX
AlOgaSlJO887AD7FU7jY8VMPAhM+NHnA3r4q95H7aGbzA1wY1DDsQfpE6u44e/n0kSb32n0K/gsQ
SK+UpJ5HDH9AqPyD0l9mfGGddzE2N6vN6pO9y6xbeBVbZtE0Tn3373W5it+KDsJCDg9VDtmj1hf+
YzJ4tkansbjdWLMy8aUnhXgJduxmGe2z7c1VVlS+AOZGj8qeLfcvBNY+ZjB6lbX2vU58FwGO51Pn
OVUaRJiKWmKnE5tv9TKKztoOU4L9+iGEY8nFlvljfNJT9w6GIKmEuuYd6PsKaE+OBBjMPFEkJdG+
2BSbZz21DCth0zh5gZ+lLvkCMbyUymiIm1SGmAjTLy8WUC2Sytjr+iOSjXM7EuC/ElI1Jym5OZRU
4zYXqAQlYHzQ4kHS58rCbVLQ93Q164FPkWF0RFbcJjuNEBAnl93DVHIoO1PzNrS0Z3764yT3VQhQ
LLp8GSKgKwUrc3FjYDyqkZbhJfAyfBWyjH6GCnPoeVXATq7BiBhQOI3j6udHlD56GKHSBvWjzjpl
/RIxbHZYuITmhGyBlCeOIUafWiOT4R1d0uDzAzCCazSYZIUxhY2DiMUnzgXJY6w7LdGzPN8LzAy9
9jZyhgMdYmJYAnc6avnP+7b0DTVN9Zv1cmKRENhUIVnNDHFP9Q4otVaXAqjvxOzDnz6Ka9kFAv6j
n+h/sw90Xd47N1bFXQH+EgxuIQ1zbroX5oSex8yyMJkdPBSeoXN5zNy7WbYNUGECaL6DgEETM6kA
3z8t6d0MC2+LZKzF1KUaJ2C7Fk2xrZItAcPLPEuqG/vlWx4rJ+fjEBIKDjRya7K1xexp1TwCdVih
s4+WW2V54NxBAHUyBXJ7ppeFxUFPMePkpjhcjRTnRVY3K8LtIiLyOL9LmP6HOos9kQQogt1d7eik
JRloOjP+DG2vLmEtnDO5CoZEUMGssu9nKageOjoTM9Ek9MhVIqqgCBu5NY/aOR8pZTVvkh3VuTJO
MNqo8gNonQ+DuE/TMv01hk65yCC1TqS7wXUtpTKKZrXjncosCzTicSNxsl5DfCXr4Rul4WdS4JTl
LYYc2OyNcTZGL7nc9Q1AiujR00TSBjUVKwKuu2uxpdMkIqz7mZsMh7wpfJ+SwVNXbzL7UDvpcZc2
tr+iohyw55mBaiz1+oiskOxVFC8hzlAuvqvCy7PWmWyIdIPeFQD4VXjDjqT5/KgM0216QhqXVLZ3
VW+fENk4jLNfAWW+9so8Kb8YQCqzMB5MQWgJ6S0By9qFvAMnEHettDPtmMm1vnjhby70nnezyUSa
zm8bHf5SifAuUcWk9HwjXW68f5pGtI1qhHt5s5gr9UTyGRkxnl38ckdg45E0fkQUBh4owZoOb8o4
HjYrvOe1H+YwOVhgbyfR8q3dNcjb7Ou1rS07mN+JN0eig4T8RxcG3U7st/KmZDY5SjHAmWXTcBPM
isTy2pWOqqyYx1fu5oldZELMB/uQ5eZIgIJYe8BxxaE7s9mlhxv/rwcPsYvlsqh9nNCmda+1lXaZ
m+0qn4us1kjwDSjavuXQ+qs7HTC3oIYWLsw2nwf1daIE9m23k5Gbej6vL5iGqwpvREC4WMYvk9S4
7TY2Ctj7NqMV0t+yMJvsnLkYEvlTxMoYf/lDPI/MJT9lNlzp2z/V4kPKyj22AXPsLrGlk0JBYGZp
gZ38Qew0bkLY0FDecGJdxgn8YRzW1kxtsvAa06DBML+e2fdTLgAaXm+EyqLr7YOyAqarCQbnEgE2
HYeR00bQJFkBY57pEy6zOY8el73srRsLYZKspaVqDYcSOsn1A3+rau5rL1dEVqNkY3MyImcSoCv+
2bTJ9BEKPtnYAS9TZ2AXr5Rml/RG+039FazZCyVwYGODEXmMpEt8rvZkGMtC3NpVGsr5T/wjupo3
3i1lOfe+RC6XHkoo4ILsggM+VvPfq5b/rvRsaem3p9GYz1JAT2fHRwarMm9KPE23yY01iMWYsR2x
UTALifTBhN6AR5zR1ut9LD2z6H2cwHTVewSRVYP/j4aeIvsagzAsg4dZdVwQ6eV2kzwbL7kBgJOl
f2kjAYbZdT2GBUYZiAoJ0Kupl135tHdXlSksVxDN6ois/EWCaF+NP+KRstqcaYJyTWxJk0TCAMVk
Zb+xPl6huaQey280JHFiKxAqYNYK/4N+rNQTdBd+fSbSFKWKZ0Lwm7h2fX7fNZcFw4zPXkiXn0oO
1qFmLHGsvs5A2hcFdw9VcOZ0FC5/2Aky4k50X0ziX3LA86K9I2DuG9k/jMIT6HnxsqyTnkMj6MMY
l29oHZ/Ge6kENTVdXGCm6fMLlUuLAI2T0CzjdzmyxunYKNrNfIYWXTO2hloCgDGmczIKCZT1aA+f
7bGYH91yOD8uN87g8m4Skn4Yqami4TyXdY0gv9pAXhHAyXk3+shtCeJ0KKrWvmfvtloxpeDvKtyD
T8M4y6BPm5YVOfXC9l6pYoebnZPGsE6CkOymVqntxI77G8WW1cQpOqy3gptXQ5iSx8qmnZkbERu4
xi+HQ3Xcv7ct9BgAdQUqj8F12VcDi49ugEXo0Ra49uVlE9/fXKoBSMutrIAZ6ipMVlFQoTT4Pz3x
y7Hk97FGDveD9WXIKDnoON9eW0ECz+uzDa7q/RAaAzRzzZhYglnWwRaxikXNgptrNsi/1QUyOfAg
Ems/8OTrJZ5KP8bAUpJJzuovsslz++FapLX42l3AxMi+mmS70kXh94/pwuQoqT6+/ADBM8PcipTj
pGqUzlhxkjuvkYG9r8b/DGoUTnHidQhfsn/IKmZHB/XhoMSZItBUmoSIJ8Z7b4/CWjnblsTKxEsa
34e/GWRhx+R+m7WUNXr2EO6LhoetAPvXk1Fzrn08ZLxZmlw6fpsN0kcSAMPg5fG8BXv4e74xpBcZ
2i/Kt24Qs5tnE0LZLgn09eY5xyDvLDK9tRiYzUGZknsJUDF57/r7AtiCVvfm3LGcPcnUn+zMYAGk
qipIxkNSbv9elI34iyz9ZoXRS3vIZjgmUSvB+KH4UlA5IJiqxSot+IfM2XoMsCmbCu1IMMWiG1Vr
g7DmGi5iyXtX9GHC/mskcbfcQvm1B87UH1patJ08YYWI+p8GI2NSf/V9rXGuh5utcNxQc5Dyy56I
EAbQw+GzcVtvLIoytzfKOPzwUogpgtzWYj+hKiJeCgzNggBKwWAsF48nxIbTTmjHbK9GHuf81IJv
pIo9iFP0HWzSytz72vhRBg9crHqy6hym/ZnSV3pXhODd9lNUp1mwgaLYW7yM3EaxCupariCsW+g0
N5aR/1mbA+P2AQSPccycVaF07hdttTPrkKuzDdS9+XpsYPQiv5ri9qXhp69jpv/QjCihOKmLkyOG
/DBw7GNQGyMxdh3bJpXYx5p0IJnqSNMMmDvCv1Z1bLe/9DqjcQAtub/QdV2Bc5HjeWhMj8Z7zyeX
z+q2995miLWHfNzn+eQUH6w9/3yuk9Mnlh0W2EOlteQ3t9yvnbLa16ZzjS9BXjK3fMF5n6S/8PKE
NhJ4tkFJoFW9WSXke7UDQjjPmxcZkEbu4sHCtTDRHCtuTLbpyK0wz7gxF1bhxSrd1owEibWT0L9H
9JgCmivBCjF9FDhlJLs6d55gPLFZDfIixsRdGs8Xxxz8THTWstSfkDWqiaVWKnsYgd2lj2h62f3x
98oIe0Y2xZIPjYdE6F3yOq0Lrrnj2xRKh8kMgHjKgj4mzP7nZDMHtyQ56z8dDPajk0G9IQuPAPdB
/dk9iP3B/DllcPWzhBGv4X6ocF9Ro79sfFGzTXOCvoeZAwm1hXymDSiBGvjXc2cNJjkrdnVfSGuF
/f4LHEDGnEkQerb3IS8imQP2RFXqE3X8LXJ4p4H1sVPVudhl7t99AC64BhLGgGPFBJ7OuTvPeAg5
ReYJcLfzPBH2N3g/KRuGxHRB7jb68HTMcXtVXYgm5lT8z7+E5zxwGWWhq2YdTgOggSH1YPiYtdbu
FzrTv1mFnoZbeZQpAU/Y6cHeU1mZDqXiMJtl9x+EhQsc28PFZOAFuL2rnreKPfFc5JYYPXHxYgGI
nH86E+EpMIpacrWPeLgAP4BBqTEJWWIkeAbFR+NHlWy5Nlm3cp+x2iHqWAgmEZgjOwbNRR3BtVm5
uZQ0plW9BvSy+er0ZXNxj4UzDc832fMGoC2MZr4lxpuGw9G/InJ1IHyeAAMR5ZwL4JrJ3W0b5h29
NXbSDoFYOT3YZSnNqOM3b2CQYgT1e7ruF7JhnEKJtI1v3635S8ZpS59OFmFW4fZnFEBHcmjjxJCW
EXJyYJyH4OU1INgeuwkrXoiHn1oVl3mOdqJL8AwxHi55+dDCJZFms8WhvHnUazFAIXd43BJCBeGx
uXqzV1Ggxp9LinnA3febLE4BX0e8+N0vOH7dqY89sXAcY3E47lBR+1dB3dRGABKFYGFPe/EmJcbW
CRjxDCa/cGxDNVuxETWwaHxOk38k2+CvGeyS0QQPRXVXs8WYK4iC/PZESw4YCZ2xS61mBqZuarmX
PkvbNK1B5XbyMEtL3oe03wccYPh5JLyCftabRzGFQXeUhQfc6zySGWTa37eevfKReGm1lL7WyEwR
UWG3YK+3Advm1TPPWzUtRrqigcKjkjI3hnuInNz8t4jJ92CLYkv8hlo7pi612PcE+lb2V7UaWjDM
H2qeI5IIAN4opPgf/RWm2aYLY8XXQdTsgYTxghxI5mVjeevBpK3MaBULyqi268gOLDbcSzpBfuWU
NnsYy9d7xHKVwY0uoDkIJIdVn1wIfhq42qUg08RUXULLlW9YiIkPrZgcEXth+Q6deIs3s+sUtAox
NDfuB6dGYsYzLUZGNP2Yjo9kB9UCLaqLCdE9KXYGen1SUiQi76y83eBRihF10pV5sj5fBWdXjVc0
PvOZEdeHL3CTv5Sgsv2CW8a/zzfifiQX6F/nUG3Zau7WDM9Bhc1I/ymF9AeRHb94fZWiwJ6z2suV
7esmU0XE7QCKka4FJjT8ySKTvqnQtDoECuJ1LguEcQpirYR3BWnZM6TIaxnsEp0BTVT/Zu/ZhQzY
FuiTB15BYVbI0a2t5LBh33u64nRwHdelpGy54PPxwzIFoqrf5bwE0418h6I2rSpQCclGFPDcKTt7
lwzoa9Jk5+H1wq9drBZ04WwM8O73jZ5KkcCLRa20JJzW/gk+V8c2gP1FPx0pj3li2a25nALIqVyM
GF3nM766WL2Nu7VOfkeezfV6KZ7ehRgFJY+uJv27Fy4UU/Y8NjAkG3ObjfKQ/r6rmag0MLASj7jN
36feZazSQks9W158MO3Vc0YahUG+jRv2OUYdgErYUuxXaJuRtdDXjvdOplAKOxRhpCsQcsj2ncGS
vL9ux5+mEgoQNeWrYFIEImlCvT7IwML8XzjToOfKqa1K0Mb6x3UFUCQLHrU56Dk07bEug/0Nob8u
loEyCfB8LBH+aBlGq2iYXjCg1764AoM8hYgd9r+8rxlYiVyib68mxcop+t5bXrmh63zZp1OtIWd8
bz2W5DtcU1f0zW7TpK8xp3H0PdFCdKT7MxJ4gYpFFlQOuBQzre8Qr+wvF57SCrxli9Vc19anCvul
3QvftumLhbAfJUKS7DbOpT5KWWIJZgCrHpdq8VfX6mS/diz+SUHszG9YyNX0s/sFrisya3C4B1TN
ASAsFv4nzyfau6UQFRwa4UDoLw5GR3/x9k7m3gq85w2Pv32Wy1EFslCSURCdZquL5zL+fssZjL7f
CEysbf3n831jOGMOF8/tRMs/80GlTFrf5isvI1DsTcq8dQpMSdmxhAaik6GHr2tppxvqtH2lCvr2
hAcRqB1zrY36xoyY7i7k7RrLu0s7dfvrwfuu35ZQNLZn6kE/FMcMb1NT8kwv4+jSeLl8buo95htM
U+/ick0kBDeevCSgcHnxF7v02RUV3j6ryxo3GSux4f65z2drVP3pDAp74+sLEM3NZ6OpSvuINM+a
Iiie6HDFIMyosOrI3U7uDfE9d4SjcThcM+xOz+q6rn3zNH8F/IuUB459FD6AjkxweSzlzmFvjq0x
3aBl84PMifXztT92aCrhwBkthD/GzNyGtmEib/odD7Tpp4nGQV4OydZqX1fYZ8RRvyiNZAchNujI
uzZac1bWW1sH06Plp8PVb1Ejmpc4W6WsrqqPlDfAlywxVZne2wMlHZ+KFsSsT2tc7DKsj7j1ZL1q
y3DRbl+dE+V4pf26YdzupjKZTCCscss48AD826dLEukPpXwWQ2S0nbkql+aoT+XxYPDTJHNpBHZg
JEqa7uy13ztcpR5XUaoHY4uGJTGRGNtmRCHYiLRokh05rFuIsvhNQ92PdlZkAWScMni7cghsuzx8
DIgNL+kxEPa++8Bj8PRKn8NyND/xHpKtehO1/2BrLvgMhvLeUXA275bYLO5tvHAq/fzd1h4ME615
rLJItuVwesUlj8goXw2oAOY4rWLdAgKC1/NZxQJGf1OhmCw7iHESnbzfI0Sxz4SvKCbsgJG7ckmy
C+GObc6HkKa1HGYj5hTqK336rf0GZO+/1UJ40ONiIWJOfTvdrNdnzXy+q0Dn3ENX3jjLQp5W+9JM
/fEcHuMXdRb7q7v2QtEhKPs0qYriuyOe6o29rHDM5pjI13An3i9pZSlLlTBNBoY/Lso8/j+/f9Es
C77RsIgupnG89ardwtvbtEc4PqSJDutYEdGC5rE6vQaJfVWNzJIupltj7SacyJhjYWdvNiTc6K5d
ZiAVdFaidmg70PJtHJV/Rs4GsnYxcyz2hqkCwRNcZrMFr2l7Wm8AW/r02XJKXhqyxb/VjiQw+uIT
x8yNoYXdK+AuuthZ46hbKUr9WZc+op4bvi0MF+oxk5Oqxx2NKgm46BTj9B77copxZ3Ka3y9Z+9Na
P9WmVtQN8u/4McnGZ+rpMq1KokXp47UoIKjtCNAD8F0E6G7NWs/b48m7tCtnAGS6kXWaE5rSZiwM
aIf3KAkOtnXCcEKLrGRoCKX3aDyVl5amH5fsPuPLogblj180kxX7/gh9bRZjtyE0RkdDhSDoOk9V
F0UvMfNV75hThNtadiOKbSAYz39VnS6RRtTi5ky8fED51zuHQMRz22CzZSpD+YnDhwG/ZbDU2pki
EhlLoAm9PCVDe5v2XT/zbX1G1be8OIOx4Vzh8FSMjFTqprwWbmT3itaOgQrkaBWTjag6KllAp4jQ
BT/4S0r+irni/2ag8SLBKJzqih8/CrL8d74yTYIvunoML0TBo8iMtPPwvHs1e6mkQmxgZmbfREOV
5aWBz01m9trLCdZUAaN8wjUBXP/fJXTtKyTu0bEQwDap/ZEaG6nW+ysaFkVPdCEX0tAMg9wk8fFA
Soc9FrPjP9euQKqS9CTYkdlvoz2ZbM8P3qgfh8ebWNdxQvVqzUvP8Z8r65vKAmRcPr/jXolcuWJV
cGAhhYr2tMNoEIjgtrGb3+lLMOqBzUC8FGVoQNgFF4BfQ5N6SSLZLjat+y8HowT2Ob1Y6RQli5HC
jKDsgRBY522PK8l06sP6xXOeObfWst3e3bkKjToS32klEgqWlQrFd4fvgf3uLTn6IQZqZ4sJFSbW
OydF5TRDVpcePzz9flRgv2HJDybekFx+CrcWn6xQvdc7O6zk5YZ55/DqUtvI6Su65Ry/CLfwJUUJ
WEsJc0bHwPBGAwgHy5JKIJFdNeu9hbSYMVmpakU14o2I0tcVTXSnsne9/PygTzFQ3XOpV29vDmj4
cDKWTyUfdhZNVpmtj7XabgdN7+z04PoGYikkUdhG6muQ/qJHxUvi5mTUWsMv/8XBccyvRAEn5JhV
zoe6GYF7/DVPElxptzj0F4t/q2lghLlCaXSkZDNrdUDAeIJIUttoO40jD5jGz3GVNwBwZdIQoOI6
RuC8llh5kz/wTpc/9Fo13AQuMj/oFXrSXhts15OO7JVW9vPZlaIjaEZRJznH6CdCgiF5E4FTlBYF
10CnIeWKbqsd0DdUI1MNmi6LPqxNNO9PYAza6QWMNeOfE1edxaFIcU7gQlLVYcBttAi9mGSukUOb
Ph/U+bXNu0r7WLetxqwojwxyQgItVpW85Yx5Ej2iKQRI+DIHutsQd7FXQXAExf273IvF9bxClYUN
6sn8Cy72/YTs0OJGSRVBaEn4KsdhfFk2/ttYWhiTyyBsNfEInE+KESaKepsNP7HdiwC6EYRsbP1D
d1TOZQj7ZR5KpDoTwujMBel85C4Grc2dKlOgemQt2fhACeBkRZfKzRcLzgMYm7S9EPQsND3biw4L
Qb/aGJwk84jdVZrpb+FJ/ttmkrot0UP1fOVjMF1/a0a+Ea//NDySC1G5JIMKZQ0JGY0FM5N8sRm6
ynw8W4XZOZGQmIArC1wIUetMgIKYHsfB7hWOTNN+OSytA2GGYLMpBRFBf2iDCTVb6sjqhdEQ2gfS
iMQ7HZFF7YMiirq5wdqaznfue/RPUX34z0FdG3XaM8Tmbw9WDygKlGBa/i0fCiVqh91i38Fiv71s
oomHkHw8oan/9G6zEvKI7KbEtdR4gAj4/VjMNrsVHpU6pvW3M8DyvuW070nueueImCeJyyNMLhUu
BBZMG5caNOQjTSAnhCEWUfht2VGuj4KjgYU9ZyJj0yWy0rizPErPbc6ZfsNG+WKECOfS96aumPHF
TGDI46BIXRS/vRjMnVJ/QkMW5iHxyOMXuNfAUMDEoVinm4OvWVT7rz51qOwrMQfbvoKsfLSBC5sC
LO3I6aBLOdGSI3jRaxW7gMzCsjvBjRdd09UfatqiCDFCdjCL2Cb666expGTAJ4ISJU4b04UP0xi7
HZSzFrhjMyK0HNYfh7KEBun+TwPk128aCbBBwVAjC31N4YJUyYmqAxRz6nD6ROLqxR00DE8Q50Mt
AcTCLnUc9UWMmhVdDaD9bOLstpt+/B3LjBtSiUnXEo0n0g+/OuNlAtOw+yPvZ89aAzkEkVJ0sAfj
WE0pkZ7WPoYCTKkHxYgq9Lo3j99hBkahb5qrZshmToM3hYfV8X2aP6XxAt+7aVVqIMBw+sEAF1Yg
SNh3jC7nf/Urdb8vwVZOyWUvnlql/mvSVcIMHNcr/QU+SdvJZvTVyGebV1VLR/SaI2SWZ34rggQL
bgwaBDoUPNSWTBsRtwN0bvJVMC9skBmpcCOkWx0wvcUfNRkbGf0zwzGKwi2iPDwEYm4RW8KPJTr2
YBuFknUcNVaDWwjku0gqtlHZVqcSDLNnkeOotnaqJAOACv0toqe1rRvq32tsML6XFjCg+7/WK4xz
63j3CVh9wbEFrEYowKyh1IhZ4XWGWbTcjaM7zKc9o52a8c65MtfQpr8y7vWpRupak/UPQu/P+O5h
rIr7WggeCBpyUV2gYl4QEp1t8tXELErnO3w1DzNL6GMxTPAKYf+AA09kTZTlXAX6NsDW4lFndVgm
WMVlYiE2piAOut6zpYPLtHV8JhVFXQBARk/Yi7yv5i7zYC+IeVzNShUZFzGfUS8nsMHBZaK+Npkr
vsQ976QpBVChKhATItXifotPEqQY7b4g6MN5dpk4Gl07t1fd60xA8Up8tzEdRnAUatkb35eD9M1r
61zVmRKTuHbePohjH+/EhSt2rJgWEs6/kFfnO/a7fpcteIlaxHps/3mj8dmrR/CVGSGVMgRYsOcN
W3NvGIlo7uDw6wjEjf42Vacu3BAYpZ3pXzKxVF7Fl57TI0upIdvaqTEMJVe/3xpaI/D5D2eyJAGd
EzTEP5enghWsPnxgu3iZ2Mqo8RIJE1Z7a8CjwHlgcJ+H3H8eV/kxvW2JFdi/pCmzsNYfZ2VoGOyG
IxMNaQVZQDUeHPVxp+HhGnJl0H8UXtXzzw4xXzNb1ZLV9uwLLNwBZat1fR96s0ecgd6T0ocLzlxZ
6sWkkYUTGjxhm25yG29Z1I78G1tXcERgn03i3Avygffg7bBuPglv2LLS4whWc5nBqQGaqQKw09Ei
kE8BLKn+D9/P4bJ+w5rUo6dS0JVr75dHPK5QOFyG6Qw4Da4iWDNn2EUXARKRFIifQ+EBCawZSwoA
AiyNycFaWlwzGXUtz5DORRoyNM9nIvvIOI5bb3s6n4PcYxJbSmQKQ7PVeMjno+rAUP/8slrH9fQC
U031kv/0ZSx+CcTFrlSyfeBNOE5O6n/NsOQMtBdDJlIBtMt23X4J6Ds8qhEjSdqbT4LpkW3cGAem
VOepRD/phgofe4cPk+u1/h61wtu8CeEC7d0wTdyRk2s5PNU50JRpqglMSP02a7x6aCG08zi7fMnP
HCAEQOy/2rmDDqU01bwTwCARK7gV0YuIZoWSjm8vfplBxkEy2HhQm05tpwAxAiozdyIW3x++l2RO
/eevPR1D7ma8oEZtez3ggZa8hn65lAhai6gXQ0xdwDsi2Ea2bVgARf9Q1as5jf9MLP4EQjcLOpJy
5ofynJH4HMTQCbd32I0G4xt7W6/LcZTWOfwevDzYCbQ8JYw5I0PJs8AH9VXWeFxUnkwQNVbpyCgS
QHjunGJ4uULlGvLhHW0j5++TPAtTHWo3YeNIaPBqgNfjiXwFgzpDvIcxXfD5Qy7o/XAyM22UMjw7
IhLXrzOWKBdSsJNmKbVH/Q4SfvyaTGofXrQT+epTgjSZuEdUqg3SZpcOJGa+pPb4IkbeS0lpwlyr
aqjA/rH81qVpv9KnWf0h3RFANJLPIuxbr3YvIoRwtL0lbtHZnq8lcAcUaagiBRZ3cuTvorFMYekq
ISmnezKtktTlVa5LvAIPYNacJMDeI30KwIIAsxkhrj1OWYIxSSOOzrK1A2eBIxTx35H7QHkXTeCy
2AQJZAHrJE5fSFHsHZE0TVxFfohvsPGCDhmKeo+rbeVWCe0cbmPn64vsujJo2pXzHvdhUh+imYMh
lR/k1Op0Y3mncXoudGdsl2oEejxNqT/gN8TkYyvVVKhIx4MrZ3EbsrvOyGzTUUG7msCLHg2msNsQ
vt+6S9ctAVv6AGcQQ6FpQYgkVlvTwN/bhx4AdgqapSY5SAyz4wJUtMBrp1pEOu0+VXXk0uAupAxZ
oAP5daAsfC6xMG/euVkXCBaw3vBC2lX5UpJLjg1AVSgdCnu221n47IUvWUOlVOmJvY+8mTUb0m/u
xSM5v7cxodIExYkjNGNhJM7IaFMJTCTr777k/PskPHETCLKGxV/uWSJkhBxpECqjRUVFakEhGF8F
seSbyg4qX/zTyQlidJSsHag6vU4FXDcfIf1JIV/6GwNon4q6DPv3BSR5W3zCgNRqXOL1YsCfE5cq
lS6r/+HfWqLVEH1x2WbyUavNjTWbF2qCFqJpQqhOo8Orr66h5b0LBvJuFbC/6xd6dlslRgYU0Ffv
ynRji9VELdpvWF+fENWNBbMjAKlOZVWNJbcEoSkeovQcRbGA9l2hRIvSJlHtg66LwNzNmhkjCPnJ
eQBAZ28pLTYoktmiCJNCJakQsx+CMdBYJ0KqCKzxKXIFThYSiWN1Dq1YSSfHNiY1t8b+IxYjEk0b
Hvu1LOnaRyuP4zuOhdVVKMViqthrElQomwE8HIjsjefcdpA6lB3D3m6J/yG1nst2RhdhpIZGrg6R
tNm7wB57BAHRnnjufMTb3Tcn8EFyAmZKYw/TlNdROGiCHkp2CtxtUpuOVNvSJLYZwEJzzDbKskW7
xifPOU3HnBoti4XHoW068ZTU+d6zy156/WoRQnzLy/i0qR3XJo+EIUmBBYxW6swZJB9eYNQwgpM7
+G7Mi42GL08TC/IVmCNRK/7q5gOr9vs3tIzSlo7rvMU9DxBWkwnFDfVoIOJIqXi9QyEBX8JVkkpx
ORgWIaZNbUsf1tuk2JvbnK9lzacszI41U0gwq2F1ry3k4458tACzWjr+xupvpHKrUTw308aibUJC
I1S/DBEegXbty7fj+DNFG3cYoCYZ9pVmHTr0Ol/VzJaWVew6txha457440bn0wv+fMEavnEKlHHh
UPmHFo5yghoctOHueFo8kUrNM525PVOQkdqhdeKwa4fqjLxJp+a1XS7HHCsrN2Tscz2XVBD5WPFT
q84iyueJpzAAdRgD9+GEeZeEG8g3xaR+Rd0yzq/2AuQzeQQG3WZD6Jx0+UReGwSD0RnOY37D56i+
Sn8iHHW6tvUqsaKyPigUa9jG0qtMW+JHMekbUl+rqUiXv8/vo+oihQ5tWqowIIMtUgU6fcIUiMVX
iYUAVb62EQrWNBwwchTUJd6hYsnvfyhP5n4P7NC/PqbkGD/bhkabb2B93poKj80ePr8TzNHvTuc6
pXpLQ2+NB9DPgsW514XcOYQE8Q/YQ+AWRdWZYRmj2pcQRy9r/p/A73gvKTvcKVDhLoROV/s+dWg6
p0dbysl6ebAbTNYgVMZvFVKcCqQWzjzbhZy7SSYQ+lT/b+EaSfmVoK/g5ZK37LbzIM8wtMgT2P3s
6CsKO+x98iSqbewqDNHkpVD6vGbWjOexna7r56+UbkGtuvZT860HJcGWNsLmkfd8XBxpIqzNJ17D
spBHROZnYA7NcmRyJIJ77APv3Aip/U9OlAg1gK08GzogoskohTj/X6ltwcZA2UwXja0bjeHnVwmX
N66ZUEremBbgFT2yewonhcAFVOclaVXkqGlzZP3SuEmOadhrHiQVs7TYMF2PbnSBm5yM/XzxDz3Q
6QgOx9seGMMwgaGuXM30dZNWMdZl8rtqGzpgF1NFYxm1yi0FR9Dj1kLTFFvAMeRQ80d1FYkBfu+c
C3Rat23gE3NusXoYKmX4P+jT53j/OxN5JYQj41lYNL4k/yx4z0ms2hnrosuHy5kc+LNi3Ylche+Q
+QgnrIDHiL05XKC9FkL+6uSSUn+bGiJGpaDWFZL7f2x5ysOoSWe36sT9AUE2TOjjsTMFjZdeWBfo
1OgAQyhpR7Vaew+QfCSznrIz1VC3hf0jKaVxK5h1H40SLdQ+OFnaOqdswiptt5PAuvCJv+ddm5mB
r396nmWff9l5rTc6GCKJu9UGJUZ/BExQTBYnfdKHKNKcKsu4j3UaIwJi8V54xJIlc+y04SVs6due
4eyBw6hYb+3eaBuqM3yBbrsQ6uyz7j2uyB/ptxQdqBx0ZExXijJxvexMhZ9U6y6lrO38Vo1kH4qd
Cx4VGhg6UVlkIw/jQKcy4NGe64J12y+iVK/jKGWhxXowlsLxwkvyrA80PmPRm3bdw5jdtWvZSdtl
4QbObgYh+lmE1xBqNZS28Lz4IDSnS1WT2MQUWsy1x/MXOvJz6PX9pcIVL0Mt5nQ79y5hSlbmk598
mTNBClnU8FI8MORrP9E2FVDYUQsdju42K4c9ELYRXJ2wctM5H9sTiajrAY98hK9Liz2hNEUETeHa
+/k2J1Z83/ONAUK4ALIBaRVrZM0Q/a+oeKMDVFH8aIumCI6x5+npJs9H8lnQe8zmdZPUf4TlNygQ
cgERSIrD706sOSneUOsmEfhyCODwqYdxpXZg+4aOvnoTfkODnGIw0cxGlw4gQRgBhiliEa7yvxOr
5q+icxdKNW4eZ58AoMRGzYV5LzWiMqFDEMcr+8ts5kaENNZWi9cy9C62F0jXhEUfzRv2gzWXadzX
DiIV0d7hcBOIc0bKt7ieTXfXhbInSAbxEMjcGJQa3o7bN4vqmQ6PEbF1dybBfiZ6biMwidlY1NVK
q2cOQs84KJpOiGIvS6G0xV4wneSjaRvlQ2b68FJpjRR8UIFRamdEctmCN3QMkLbeipX5sxgvylyd
nl6S3kwIH1hXYm4IVrJ+uHw8kddFT3oscLC909Qy1xXlDF4z2Jrfek+p7yZEF/2qwCWlfTMm2jCH
xdw84U//d40/kLghyvzLsVOc+DT13zR3xelEyPn8AkxLMoayldAINeJm/KesBpVV30H/j54qm9My
qO5nQTZl+Kqr3sZ+69RCkMskjpHqkCiDxuzWS8N9SxeEtHarfkAl9PXdLu+tIxY/uGv5s9gd+M4L
tcGAJySyxOWlPQqrft1rdX9hasb0EP1sdNF3rv2zMxJ6LeuGKBclQstlvs4a4B0M8Dy6pmlU0pD5
BidgIQRn4CsVMspvvO+CDoyW4LR6/EBmMzDo+frWnrkZM9H36sdiu1M55qXN6nc6JPVHWBPfCNNj
X+nGtcCswm2rkxdUEbT6onCaBzmLc1dLsFUu0OWZXw0f379WJsTZJvuKFND7N3JKU/JkhC6qAxHC
JrPC1I+Nj2se/Bzbbw5gJ3gBhdPNJog2sg2urGx4bFGIF9ObEq/GObAigfMKp1K46LA9yuP7aLNK
F+NMPVvajhkE287dEmz5bi/aUj8ZIjwx5BDrOr1b4vuiTuT/YfNGUmkHU12TCkL5Tkcsh8WnYgK+
d0kcu8ab4HJw1zqmvtCeCtILz8Spetkor6648ZzGpLVTfsu6bFKQ996VmT0dd4WIsU8T0G7USQff
vmXfw3UtUmNERDoO7ApaEDOfFZqp7KBqcD74sv8wjDxF+RAfa+pLMPFwFtPjjsL8akyBgKezK4LC
2kiUopuu7Mk++Ck/2Gum3bVGSav94okhkXS6OLWIqTG7GYSXxxtfTVa5QiH67tg5UIm+OAxbKF3g
QG6Jq+hzK5m46YmBc4ugn5THXdlH1p4iJ8nbZR947dT9lUfFUp2h+sTsPa/sUCh3cs3Ln7HbeMeu
G4V57KEbsq3BS4nsqNnT0WvK4nC+nxaacZmCdkj3Fu6jvMqh4pc0sefcyzxOmHiU5DueEfA5Pg9d
Vl0mAUxEys6wMKSgVH9vVKQ/81mNLxw00QnBE3DO5WTOtwLH9BFl87TLELAJn4dp75cr3A/XuUDA
nPiCwYFPNE7svP7+Npa+jCblWVfurpvpK4BrkHwJfxujhH6ABjKEyqdjs0SkyNbCq6MUr2WGdhzf
KqA9m3aUUTjp6R139vUm110kKPIIpFlCMayQv5P49OBy35bhhSVUW7Fxali2EnraPYMdcEquV6Vw
op1HqZN8sCeHjv5FinJjRPglI+9+0cO60rMx/TIjxeKBqDcBgEkBwJQPblJLHJ1u2FA7LYo2N/6N
wOfLS2V4iFWmXNZYKmQ5telL3u7pQxHXNGyU26LOD6RTuCVzI04hcCmRpM1KLil07nwt0ynNympF
atDiPtv3rrW434csio9btFTszHno/aIaDqPNh065R0X0crqOPM/BStdtwyuiscTpq2ZUWNk2OvZJ
pUcHzm4KFMynNHdVRKxNAckcIQCV0Q2zmAGIvlYiVZKGkU1PPvwaEePMhu+zb8AJRvSSGxTgHCvq
cz8amfoDonDGZfz8m3CLuhmFYIYw8H9kri5HzdK5lCFLcfQz33hkpEHjLl7Lu1lgVAzYtUbhUTnr
h6HAT7YQLjDmig5USLEmzfvYRZy4rW1w7JUfgwHaybxCzRVKCrz0YYqiZFFO6WQF55jE/J8LkNrI
KwmL2e7d7ksjwoFeczobMMxhgtpwGAExwLCc+Zzq17YHGquh+gn7gt5stKaxB/8nLLaep2ATTzF3
cIC8sWvDGqgyrf23+mbCVMdK/LxXPMgxIqV1lnPk2cMoGJUklBlil3NwkecaakNbmIgYIo8xCfoA
gHDdPIzLoArWrJcqjeqfOiZaDG0qOc7FGj1NOXImuOpuIq1embiCFFy2dn+HMarC9pQ2qTlJFSWh
bnFn6+R5GPGR49QCMWLMgQ5/w9bKtaFmEtayX8469XFqGTDgKGgC+clQBZpiHtpW+XDtdSHzSgtY
OBHBdzG/iRaUWWcc3anYH81tdRarEKZDKAYaifPlxsp8/HkCgWKMU8FEY+M+KrIkF3dGrEmnfraL
z/8TeZjT2hf/tw2EvhPvfmWeQIUfj5C2dAYSyBuf1zlGlWnDfELdhI406nCoQIIkHxnOCkpw+7Jl
1xlZmkkZNVJuVaDzaqnaSzCtMNpfYL2fx74wsB6shMSeBSFiEnbBscWCrzbY8Z++CVGyPK8X1RjB
eauv4nZF0GqO8CYrITorH2+qBOFDD0YSS/xg8pqrAfZ3xFWYm1B/8DGVLwWT+dNs5BwtyLxzjpBn
65vl9XMKM+NlleM0ebMTd2iSVF1cZAgdd4Wpirc9YFoHHQmJYYi7GLz2Cs9Hj6JMgAQ/uWWz9dme
NyC+lxOp+qpuI4SKfIZ1cSy76wDrEvi9IKfWaSXSGech+V7i2yPb8SxYhNJEFKI3OXcY56qDb3XG
ipwXNEjMMYVABt+NujYcqH51doZa2phaFIphsc+3Wj/kiQsXDUK6xhv/r3dPQnkk9Uw1kfaegvsO
yk9DW+LyMVw6X4EqeIpDmm9rejrf7kCZJxYZuKzRNf8ccmpXGYXPWvlQlpO+GqF7JfQKRWCwCvWw
EFT1o6YKjlNGb2uQEkav6BPI45B5y4ZB/bhEcyqpnv8RBp9rAQDxS0W176iJkQ5oVx9SSBcATluf
PLRrvUkwXwHW7f05W1uW39pdGVQBTH+fP9bX/cnTMRg35fUgEKSSfjlwiJm42xS288Ay4devmUGY
XvyIl3vHcjZQKW35jD1i4cW4/Um52lIMCGqKvYSaFj5LrnTgkTYIwbUyHiwtyFa9c3j9BD596/s/
zJkes2gkRYZb582OD5tx9GEe2Gco08Be/J2rJQx/Z7pkmLY4D1QY0kDJOusnpEdyfD9oiV6pshAY
+QkGo7Ee5tetHFeX/saET4vothpjiVjbjYPy+buH8P4/lhz8hfyRMAZX33H3GUVmeYSvkbGu881Y
pgwENHLKHd6Ln1KMBma8a1w5wW/S3QZGexLKCyLno2PP/DEj6GMHIJ6CbVPTYFiSwII7tcL5idXV
eZ4o2yk3MgtGngbcB7pDLVPVmDAlULFyItBvj4qWdOCubRHU1DQ2H1ieQoYelkmMpvwFcBcnb2JN
R2SWmZE1FH8dPJB01/HMzOSBNkLOc8co2peEm+Vawo0FUbFHSWYJf52SffjC+pgH36uj8x+aw7/Q
U0fUEKSha4s7Clgf78SVxXkdMTM8paU1sVg2y30AlvcjAM+FqCD1/7943iXRSgXXMJk1BExXxqx2
xpNW9Udc0QeiNP95zmnZmGzEVcb02QgOw7uoYxhA0j4BYFFg/9YEw68tMcktB3LnuDcKyKXj8ORX
CoKFLpMF3rti6ZDzLVz1aWiaOrXpPtnTfiutNSs5Iau6AzglkPxUcBk3Ij68Pe3KCYOrLQ5e1xy5
yxRqRCQ8HES8zxmLPZO9IpEf13Bsc3LMm1OgPmghAgw2WUx6+BP3GfpRXiIbIN4NWjDyezLwiP1s
Sb3yGCXmAR7gsNIO2NdvfFuIWzuMgwM+FB6PMlqelTLSYX1Y7tQmdOpvQkwLIUW6+aK3pma5g+z/
quoa04VGBb5VU5HdWHElm4um0/q9JLnxecoVeAzZafUN8UjJu518IgQZHdFK1+wMwT9lsIx/O5q+
2eI8/9aIibZYtKacrJtqdJ+enLTA9r/TPrR56B46sO6/PM9ddwyb4LDcri2Hewfrlh+7Ka1SduCY
BdjUhzvPV18qOsUD4ayKSGJ5YeAAG7Hk1R4Gu64J3Jy3LvzHD378GdUol/wLK1rh9DD8YM/QFGTb
S0ZxNWVWy8/2BDudlk6kkhf3MsHdxOZvS15VmkreUdgyNo3p/ECZzEUZihNXacUWJ39C4JBwUdeI
rvBfaUqJGAYrrC1wDmlFn2XKpAnDSj4ghvcWad7OUOZlpOn7zUihwpsnpkCF9shtkwG+VsItYHFa
zSqtD/lhPvgb+35BSSrsdUDLIQcq0789tYQQ9WU0cadu9Tk16w96P1oUlf6mLS4+mq3azEbZEnyc
2GTqvdX0DJrciOT7ea2+fGnv2Ou/hQW21A29KJPbrY3qqzIMWSO0xPSup/CeorKCezPSplA69AQF
SmfNKP0ybq8TIqhFiSektfJHx8/YAVGBR2TTbFLD20Q2f9JSMsaLs3vJC5AWrQpkxQNGywVu2Sg4
7G3EZnyemb0CGnGQZGXhEq3QnVKDxyYN4zRM1rZbrCCRBRuUXy16XaNXdzssvreGVXR5PUf5NHgc
1DBfZQxnVfYmx9gHutHB5QD6ix4umy4JONSdRul9nzy2phP+OClyqf7/tutaQJbYoQHegddhq45T
eguFaGjOPbsrBAyTeUoK/aRchs2dV9VcTDtkbC1s4cnG8TOCbGZhwypkD7aOoVuaRrRStqVUNnQW
f8Pvj1VTmwL5crMBj4hderrDPZwc1WIkzAI4qNlfkI+O4uOJ/N7FksQ1k4qSE9cdz4Y/wY5nCSsM
8ENmXpypxO01uWFVuwyUc5fF7mjwnJrqQQY6ZEyXNe9pGaDXRVwnLz6PMVzNQrBgpM1INKFg3x2c
BeeeTSysVWvyx8wKUmZ0xO3iRzmPKyq6UIivtlHe1L7BV4wUNiH40yz3mP1pd89JZpdzZ+j5BIeK
ZnQ0FoUjxMMVIePdpTrq0/sjuCG3bujpghJTSP+QcDW6iJSmO+G1V+BNrTHAilwpzaLN8Jy2DBeT
tZEYmaW1v/Wl3+mR7IJnsDXCWxMZSbGQr7D6ri5Wfl1Su4lJRB5pBuS9VziEekXObgXid1vK+tSI
ILZxazN+5d3N8xkrQGuuiQytXF0PaAAlvXgF9kKG+yI3H2vo/H3MlBXoziPBIFlkpZRpmLyIXLmp
WjjjtLPA56WPeCR9kbpEoxUUTYJ+MVt7X3Sb78rvUM5DZARMP5QOITiULlBBVtOMIOdxqI2VrorZ
4jPTZTA0mWFvxPlKsNT4Fyp8bw4jHoUcVr+jPOJh70lVpq6Vvgd2p3De8ieJ+YrmgWlpsXaWim2b
1l7C0W6oTMJrncwYjJdbgZKeovlH/NBteqUxSsipp9IVwU5N4XzVAQwHImDfcpJDQIuBHQT2s2+W
Ivd5IqSw5TKWgzmFgPYX7bZuMrFmWM9EClwjE5z2gXJHMZvuyy8dGvchxrNAXMssPM+Apak4YK3E
ioQ9M+I5lftmepk2h9cmEa2Z3QwT8L5AEL8lTjgcpctQPSYkqMtirati26yQYwr6vrhY91ZakEdz
LDCIr35A+a7nGQBBpQJ7XNDxZfhyMBVvIOlMGbZA73zYGCEQD22JDLQQyuizOekpxQ9VKiq6Tuou
jjs3aNySaMBg42WHLLUdSl+x49PdCxJrntIoHMMQQzbrIH1Gx66S5OXcZJ1WrTvWaOr9FFt7xOmG
m6a3pxOR62tAaEwK9U3Pe4I18fswK17vGCkP/jKL0Jv3pu5gHJyYWhYvFmyM7QeOUKegWboqYgxY
ZeIPSFygxfvH+nsCXR22ZCDADiwFv9frUfbrFqJu2fLN99vQwHfCr4W+N8C3wZJB9W722TturSxj
C2siWonAykTpKr2WW5FY6uINThZyCdecxiassg6YMU9owP9uEtF3PN8ZIBiSSv7UXa96OmNtoBpc
tlmRbvNT5NT0o4faNQdvlZF7kiBdnNcwtyb2bm1Sg93v9jS1FVpTeUCQvU1FkLxTlH4RdInHxrFa
+A/qodgG8ogztJb6qeBCwzAZHaX6apfSK23eFqG07JsePSygkm5A6IXVIUDToJRRdmJZP6mXFyAO
fAMjCizxRFtWLMojCnj32J/mK7DGlqN1JLe/CjYMIxsE1uemGubQhg0lm0fq51tpVncSV3w7y2Y8
dotvCaRK2FUXzVkmwo20uDN/EIrLUtDQrlwGCmvwi6MWBQrKMLPHK0MhRWG3LqOimSMmfYQVKdV6
xXRkPQ1c4hVnBlC3y8Xh4948UKmSl/EpPNSNs28L7ArH5XFdRPIhA9iUsT/hMbwZJoB+mwUz8/z/
DBPvrhIAmyfpgOpL5e4MHycmg6eKMuVm9JTXRO+FMwL9c7nPmNy72Tt4mQyVHRB5cYk3g903h4gJ
+geZ8ayg5ePFqNaYZNjlLhwAaSrKdbB9tuKb4XxO0cpU3g42VA1f4Z1WgONzRZThCEQ6XdRETT9r
/5vodjN66Rng6E5H1L0eUjXYUclU7Mgj2nb4EreQ2/mPG/Q7Vo923oFSj+TshWtLDvInCX9alRXs
htVldIGG6W/70PxwCAvQSicbJfKwK+k8tVNBwR03/DuwKDpiGT/LZ6YLyYmzYmtmJ5RUa1YFmj5k
JJmnqLCFlvGCBzTp7TEE3zobbygREcOBmn62Ze+pDGmRp/svPFRyVd9PxRP6UPV62qot06feg16w
IUQIYs9KwQkmSuhLbUtqnEcQz/doIHutasOeu3aGlVdVbjTxsiRPAJ0KyDaD/Z+nNXmva5v6wj6P
w3eZC5AshwQetjTERoxjT2I7FAF4TqNyrnrJLy8hevCybWMmrQZNGtQVK6gyrPIW/9g6Bwbz5MYN
WTX621S0ekVRDEA67zUjexl+yCwToPXnhRIVO4ZLvr/tRvqU4+74T+J7igxIc15HLErvkGRrUAan
pELmve3hWi5ZRDdQmx2IAIGT2J2n4O3wInnqEITZzQkZegga3+mHAv+j7j40sJ64M061z4u7/rOA
n4X+8i7eqOUHzQH37PLf3hqiBgRuPvcpneYXy0er62zIgIg3a68H5oO9cV2DlFTV6NuV50ihdux0
eUVio0KCiXEACGdQkRB/NH+3zjtXEy/4hJKBA8+aekOPzmheY/4Zb2qMQ1bK4dfrIoZKAN/eDgQT
HivFci8z5APTSRTFaPk3ZWhno/+PLmKcx5JHX53KM8i46/9W7nBZjS+yoOpZNwMrD86hkUBtqmyr
V9M26vZyfEHWpOIArIHwpRzsXxXLyXlFp6VJw36ctqDVX7jLVX9T012owmvm++I9qno3g/Yrhndt
h2nvllkkGiYpXtO9e2qbyKxvC0xs35u0nCytoBK2oOFMKmFgzvA3YbTCpivkocjEw6E3SAjNqyWi
d71PiUEdkELrjOzPQo0wzXXK4SuYxagNM5Swl7818DOB+b6skVynkTgFmtsBSQ8XFCk5shT2Gqh3
qQdVuGr3hUaV3QqluSol+0TG6h/VU+9GDe8NQ3aI0Bji49ONfWG6oL6IiYw2iM5sXdxcYD55Pgac
WIdnJKpdGTlTUj6hMIpeYyftKH/yMWg8Y7pnxYLQU+6xfGXHqsk6TCb9H1YKWdwj60Aas1zk5lvm
xl3eOmc/vGm9ShTFJzB51w60hD58KYKo8eaBszcd60HgFCWeqrLIdn8iWgf6fCvUm0c4Gdm3IA/c
70YXKlaIz+AMYjzCgriAg7eVmbQ9AxialZVSFFmFuV58VOk3SV1M7SmD0hL/5D0NL7SfPg2O/APw
RRxWeKywT/ZP91i+rh3PbZrpkuNsAzFgxlFCeDbIu0xucaVgOAE8NPXoEBvwVZqHGXRLQAWXrjXx
fMKdqdQKI7qhloNhn5txDOpvVXvVUM+Qm5fDKvWwPK5uBZyDezK5tKMD70wHOdMnODsHXvOiEYq/
FV236q0pisSLeWcd2z6HPGokw6JQIbuAa4AARgxh7fDUa2DCZzcZ9688bJshE6t8f+uMTwgUfRDd
1Nf/CXEIv7ej34KDZUXke6+D4VF7VqeCVuaxCyh/hz4IpqWEFa7lzk7UWKmIqNL18stQicVTo/pF
F3Mi1Iko0RWSI4Ithmu3RqO8K08CtB1jElNxGghPHho3k8fOTuVMwRvt+R/wLiNhUE10AyfTYnIW
YEwy+P9gCcFJFgqzKDeKCkA/XfBW378jxg86jkwxgPD10nDNfTFQQNEUUUMKgRmcYiCBoRFS5jR9
utNv3vfa5Bq7cJ6vNCJHkPeU4jkz0tbwztiRJPZZExmiepwnTd0sCb30neFXbzltBTv1XN2FOfGX
PHH8cwbeTb7piTzJbz+LHgqjm8Y48Hunjx61XnAeEV9xf+4bRW502NlvFpqAapHiSvBl9B09EsW/
Q73qWwVy+bhpbLkkSN5U3FmMW7quZxeIz8qtYBQp/IauGHVx7Xc8pWWRTGWLuKv64JI/CQfGq0Gk
2p1Cw2EWAsc9lgnhl3Zw5mpleU/Zjm8RQCyYZBE6RbeHduQLFVAbp0Kfgixy+FRxsDepPkhRq0Pb
CyKcn90TXaK5Y8ubJgA90rw3kBepHb/k1xrddwQU5vmwJOfoH6O2NB4XZMJk//9p35vNOuMQCBPf
/GiCrv/rLaUfevCDJFJQwGI7xCQWJZ5dOaWTsOOdhyCJ1si9bUxNGT1JavBIAktSgDVI/v/B9SMq
L9NWjVqx3fbGXt/pGFmLDACaoTwywreaFFQCNDVyLFuWSGGXASLWB8f9AhSURyfitvAJQnbRjYUj
x0SnfrLc6cxc0lErYtoHmdCKID6dSKhh47jsNhcr0vByEOY9QK1wMgzuaE114l3p9S1oEpM1QF/W
0wma6CJMj87yL1BqGqOSIRVHIpa4sVRCmKPgdfpiplECwUIADjHh4T/Rmlo8nb9geTxgZ7T0Xy3w
vaP0gCEiGnEJyaCywzCzOUkmB4DvMCTxaIeGoedi3Q+DpxEQA58Ualx32d7exmdscg8UYHF2UNmb
oTvWBltv5Y7CbbqcfG14My0qI0NFwZoowNm/tiJs0hTLGezzWeNMLHfTEgARyVAbBYbMDS5GRhTT
aS/fjfnVnDyj/YbZ3bPw8O353Ib8/sCGkJMGKnGxZfSUJI0dQ1Z9nkth21tpAsLGCOs/QQPmd0uR
0aCK13NBEjWYs41+8a/k1SsyCv8DCw2lY+YQIg27c5W/adhqnSXEl1L2xR7RJSFtXt1hlm7AgLcF
FmsA9jX4t3yVmwEN3K/1AMuSBZsH5U1wVEOkQYFFRNM16QPa/KSBpYefdcdXI7cNNUfnsvS5J7vG
dXDfhIKQjBHIeUm27y8I/vRDs1GfbFHevdSdcxjE/cisqVmTPPimdP78R9Fm5Vd9SFLtNxsNvh1w
5Vc9hdiOcNjrJluFHHiYTNsMF15+dgMVYFpciF69uiOrfOHvQ6g50EW1FjZJMM2w5z0QHFMfuj0l
rRpuw6eAJugJ9CgdVVTUVKro/F0igs6jsWt6wz+2kANzwC1/HsSEibmUq/vzNpHuTX+c22Qzr8io
JVgt7DrsmF3n07BAI12qKdQD+hz3smPooVDNLnZ7v80Sbvdmqn/fO6TTKrSrpZ4VHRq6iOAL3BG/
uUDKCgHg+yDziRwa3otWQzKvibkefYqzdFFWPpGsQ3T8/RBppGwuZIpEvMX1/laXwpWkN/C8OWHS
Qn0VbmhR+wO/tNwiGSMuxYslpH5WzD09AKlPXg1B2xwXo3kErPH54s/gNWwVfN/K1a8Ib9rSB8li
PCoNG150hYLpcBzLyB+7pKh9ApZlDTkwQntRdVxTjEPSecmRUILSP49MqlbDhMQvEvgz0B2dpef1
wIVGX1CZWPHD3I0Fnb+eM0F9lp9JRldArJSJuGq3W96q29ahEIGCU/vX55Em4FJtXmb4XOGOAY2i
szof0tk1Eem9lHW5HP2PMpyrin+ee4HH3aG2IXCOkuW+DVFjI9Zb1CpAkwmm1Jtc/vskcdSEpqV8
3d4xggjWzAX6NnfhvRX9SCAds1aIYKD+LqqThFD4GOp0PlSJNWHfGaooM332/BaI21f5dg0ypPpQ
YFpvWWjNMSLk8Q+SEriYse7C5jyLDoSSwxSlbCUYkdFaQ9KZjjiZJTjI1Vt73zfMNJfjZeal9OZ0
90VlGhGtsbe4SWTY3E+sJ5CI+m8tuFbH11ER5RVT6OhiD1aYcFiN1w9GKH01FSfwrK0foZkLntuY
ApZOKNXDJvzDfjKwaa03IoDS1gj6P1t19H3YWeirqRu32eBVhTThJXwX6qEzT/cI9zo5/bBPwhQf
Rc6GzVYXptgNLflDRz4akr3eQzPD1XXT7n+GbdGn27yzq+Ex6zr/xjoRoc1NJIaeP0Apq3IXGnfG
4O0DOJHLSO58FlQVdPfoUp8p6bE4+hgsTEDksi0iLOiEo+T7QFbrLrPhT+Vy015M3KKclgL5nmED
P0x/4fNu/fJ1UUBHJrLk4bsOCEuksyv8U383lOKWWjp0+IYjbOEHtdYVhHKQqbGaNJyA0+2qnYks
Ciyi+UOcTdExv4JQMNfLsM5ws/ckamENTAy+6pn66JFZts5/sf4FjLeL3Ky5y15rduxMg7h09yp+
pGQI6/6SwGPogSGuwX1GhTRvnpEaGulhFRfEVVsAJinKZlASkEGFNMApLJmAHF7jpBtwygTjduL/
KkQz0GxKSTG2fhcm+604/nlinF5uDuRc6A+VOuumFz3QuUf+OL16Um4q5DIPvGRB5uLkVKng+qzy
CDU/TXjxOozlIatGxhhlh91yMlmsqg+lGmFROIfLhfPXJlCAlDFDyqL2lZMFDY8bSpQKNt/U+EPq
lybr/hZnhjhOoASg9Tqwqmn2nXQuuWNuM70ux83rtsRjgQMSDw2sIzt7v2Efkv9u5vhVtDCMOHJ4
jznsyzozHAGRk47SWx6PREwsjlo6TYE6SEmQvN/p5fP50KZYEITQDtIp1mxze+zN4fuUeJRoCdhM
zyNAiP0F9E2UZFzMHlJpgUpChd9Q6gOXTeBSXBABlP+QvsN3H5eEZnKjs0WINxkspOK1AfZERNf7
NlWxEJd4BDG8Rx/rxF7uCywO+ulq8DTRluzX6/BLU49F6ppugvehDnFhZYjsLRnLwb6RqGpDJYCv
6hzxzKYUJkBEBd/lnR+hDftT6IJre0lZCLB6+X3YEB/1YybQUTKo13eeJM5eFOU72gTzTnN2mIgV
Fc3drjWQXSvtRmSoX7rH0UdSsvH5/JWwdZ/f/YsJn8z/Ty1jBYEAMyKM7Z4s05RiJ66UzBVAy3BR
VzsUH4mRZuGhCndk0/h9/ELvSaLvvGEi/fQBaVWvTlzbUKaTfjwog+Ap6rbb/6q1cnWXLixAeWKi
bNXZJLzTLQdwPU9TSI6iYEEXXfQmCabbSzGYlx7BitDFUX4d0Sv5vOTLgxKMpvBD9x5R+gqg/HeZ
n+VKKYCmifRfhRCFDDlexODU2xLp006TdYdhSPrfFAN2dXr2DqAaFA76seQIhNJr7+7Sy1MJZuVf
XvPYvXHEw/STapFWBuJ9esB7PCKZkcuTJBN7jz6O7QvVWR/YMvB0YkVH5EpUPRS+Pou89IpSqlG9
BFlfnaNCGH/E5vFWco7MOdPfDS/fHg+dk6j+f4X5ZMLWLybSgmPXA7sEKgnYf8jdjUi1ehOUX5V5
zrRgt1cN4JW/06QWbTyps/dQexzU/ED7lA7c9AXZuTj5yCygDJPuv8gabwezKkrMPUihmLWOC4s7
BV9NWGicptKrHdXAI0sBUJ7PCYWPCAoB1yoLKG12yIbXWksDhTHzjGvX7wLwH9m7FFRheRWm0gLh
rxEKfPasbNyEDIEF2sTz02AI7vbyNf2T3mYtNTiJ1KGQqSkw046DDVP7/ewyvmi7wn+qpWyBx5cd
KcOsDozcoTUGFnP6IdC3H10l76XY2m2iPAoXfKB25+qwh60Hm4OQ08Vw1w3BUu+MEGyEX+l3Jn0v
ybtrGlrrkm4wT/t5xaeZTEFZHAvOMPforHm+9naLrZpvaTzE3CNtp3bp27H19WkSD1pJblXBpOhq
sj4cjQobaBFMiTc3Lv+8awIF8jAzKSKjEOAb9ay/K5R2hdSggD2+49BBZLwiO0KNqJ5L1nkHzRe/
X54Q1tn16kFXNUjOgf5Ew+cs/uFJxLAbe0eb7Gu7njw75gnTZts/qQNfnVwaGrxatNiuP/IIgvtJ
K0wvLSadqNNIUxah3votsE5PpW7EWt+HrDm2Ry9gR9V3I59DD5BHeBoc48FeYkyEw6TN1uBxT5Hj
W6WZgcYKAa3eUcjKny4jgqO68/XQWnu0pynnMnjCz+1geDbZ0eBa6NQb6P+6MX5cOHkDb38wa9/P
4+MtHTWQvj+BrBDSazFxR/sT7iTJkiQIYPw0HSGqmpbbr4+q6UKg+mbVVDxDzl+mw2Wd183eDWBE
GCuff9ntvD+fhcxM/k1BBm6RNt3lVIhzIgdaGgrpTfd9usBmiP0aWDm/87lGBVrYTP7WxwpZt+bk
q2HFaRv29feUX6SANXK15E/xRwty5FtSQR+krjSjXoi3cwe4DTXRFtC3LFdMd4btGA63HQbjxZqm
DeyOqp0G+up7LOl5QlEw2xTqVPw4vDTgfFczZ+I9BiVZu3Ytkry1vBWzMLiXb5Y5D8cPe2s7qHCk
Q7ojOX/PXqwD2N31+inCMKeUciyMzzzSWbOVVW4fogLWKBFRWZJGkXQnKszOhZHCo06xfidaUtEC
sUxlcUISQ+/JTHam6ICOZOJengjk2di2jUv8Xg3bYkC5ceDWoCYfQRtlD7/ibOx3RERVGQsjGT0e
kYErQ4U3EJpuVPX4lQlOPB+2e9vn5agx6/bxSALKS2uF7ydcINvLi1nCMd+qBZ9heSU2pNv+y+0m
BtSPMm9pJVyZ22JXcQfVUCLgTHcYIG6wG+cWwa6bEf93P+iKCOFMWb0xvlPt2fVngX5grP9YsJw7
caQSvpNYChNaub4fJ5gumYdvBStswBz5M6oCoBY+DSXPeVTREmY3iyAFsCXjmc/RjHUzv199oIxn
+DAhsQb7V9MeNmiPk6/Xto2Fch0106/NOqB749kMkMQ5wA00jnU/6/oa4Oh2D2QSYvS2ldFBGsuk
fDYZn4SxtEdk1j88hTRHdwWi4xqXdQTtlwEm2xHmtu3WEwyOSQYHxLE5T666FWz2Z5KApC6uMpSa
Pl2letYEMcLt8/WIhpvqICNpFgx2az81AoUdjO4QgCowX2p9UVJRJ1FQsD6JecU0FLAP1gyiD5fC
aFyuB7U1gJL63MWV3zj9FLJIvDMqyssHyccg2WoIZMS4I8ML/hnHdXl/oZaISKa0iepK1IBCUVaN
nPd5B0CEnPbD2PpocokYcXI6iwY0CKcldbBjPRRSGdfyKyfhIbZ2IKp9hvL0HzXrNEv1rv1qt0mY
3xC+7vN8Sr7NwM3knxiuMQMZizzQ0necSt/tPR2ww6lRJABnF+7lDlf/hHE9VymB5ffOPGrR4Ozr
2stAymcoakS0NJ+uybgw7vdC1ss+EDyZVqsoIgauRZaCJkxaPzkGVv+Ba18VoguiN38RLO8QRAbb
UwZeeOnrmTjM5cjrysu6GW8DEd9ocuoaMS9cRqpMbpQHAhSNDQEQFfTs2P8XTgChC0COk/x2xaL9
GBOhMB7ni5lBJmPG7PR3pMl4YlvJlXufi49FFsJl3QI2wKCCNdYqM1PeOHP+ZF8Hd++4SBRACheL
Ma4VDqDNbrVXliDRP2MG2ZS/BtgRIoBcuCm/fWafYTVaeZeMvJ9PlLjTheC+U3DwqUMqMNUwM0X0
xNTCLNZh6d6WWir49s00Ssr9Nxuf1IhvJEB5Mm8w9pniOvuHydpauG7wCh3wKUSP+xFXIeKhKS0b
BzavcDbwnXz0xavKkZvyCF5VY5fNzRKmuzhCOCvRr2AJrcAaEJZRHJloeuPov+OGxW7i2Y3s24VD
ImPwmAZRPr9iodpf1jT93+3I+PZ9T5T3SCuMJYR0CfHHOOXUpFtOWdEomIIJivsMtptF+SOm7py6
BvzzT5DUEJnyWUiTn+fKM05+WKLSSEGgOMnvx76NDgWlJ4oMzEK78Z51wGe//SzN/fqot4GHrKry
YR/xDLpaYPdrSbETcqhWljM4xoqcYMiRKez8NJ2WdbW1OX1sPv/5FQWf+Qik/CnDQvAbC5ocZDPk
kDC9nrtzsFeNMzlPrO2KDgoEVCO1LQ9K1SL3klPnXx/Xuo+KtJj9cuzgD2YgR7GXaKDTA469jnv2
KGVAVHQGrCCagClUH+jxAbuMnM3s9lm2zZjoZwUFSNw+62aM/CK26z+980R7xch38E2JCUkIMEOD
Srb7rc8oqwvNZE3CgY56WhJsuxbe5TZjJUCggW0Z5gjFT08zUJRzYQvHpBJ/jK0DNWE11Na2Zhq5
8E4CJE8vaFb/H+T8KAy2hAISMPpOE9pLS3ZYim3+X4sl1Di/k/nKPcwHh3TttdXR2RZ5RysJQr7J
uvMebk2DSydWSNNm7NAQfDVQ/SCsoqrQMi6wjrqCaiEFD34OTVn9fTgeeC+xVTpe+ZCGlXcharf3
9jRGnMx6/GU6LLFldwqfvqQIIUzPs+sr/atoRSm9dd34Uc8G2t+HYA9/Ko1yRCQtIneOikXp4Lcf
1duoqW4EMOtC/Tk4Ye2jM/ogDJx5hVkAKGfTrm+mepC4CQKC+rAIm2cpQ6LGl2Roi4C1LPtqc0gU
jyi0mR2wIEI/x+Gj60Ko2+B1FBx3+QpQkUezPajgktzHMghya236iXDXolehHumT5Jh2WM0d7Xmm
SyYwPmRKrGmVLqPAvlwMLxB3VjpvFyaOzAjHAvS3ro67Fl+d72ZoyzxAbLYb8ISbU/rphSYiHZjV
b+JbWiW8XtmFh2Sue14xWVvM4yQsDBkKZwaAQAM+AroWJ6w7xgekf2N+Uo48qF6vkhtPT31I4yip
jsAuv+td0kpt9a2cKWsezNlu3E4JqBRiqDLcSHTfAbFAhZUXm+b2RBCJg6cwN1k6W/ElBGNTkDZg
XhmsDqJ/63aonSOorUIdNbhUuwWDIX3a9iw7yIGwRHS+pCUMKV8TK8wa/XAf8OIXIkqSFAIgHtG3
6+CN3QFPsqXab/l4uuxmJZWu6hR07oWWgzMG49onKXMOBGboiqbxU2xf3vRehNWFVSEJJsLNcx6a
Ifz7ujMdVTtviC8WGD20Jo9JVMJrW0RDI05ef5MQWNSTIXPCZabZ01NlUxj+NQGIuWN+69Y3oDX3
FA/E0XCcY8jNWfLkOppBdoofDuh1XlC88e2hhzJiZaManv8ypvh0jJaWuXPvUhkn4fv+TMEepads
9D3zmRDdzOLseu9Z2Rp9qGMEIs9BAVsNGjQ2ujFs5HnnN0tnxfRnODTH32dfYoDMa/CkzuEiKOQ+
gKvMqYveNBBJp0SkK/l4m0ieGa2TpHw8bc4TVL5s9dF5iSgcV1uTTIYcWPAxu/cyOXWqMDGasb5i
s3K5samszAysk7/RJ3251kUqH9sLHP6C3BgNlpldip+W9ZjqlGhnZrUg5OB3UcqywbiGTGwXk/m8
qHg6LBg6+bKNAeU0gSkJ82weKS8/18INzy4siWm2nMdqdjz22ltr6qlq5ydSkpZY/USGnyNGYTNN
3QcI9qotBMfOnV+aY3j9s/RhUC1MhZFUb/+VnvWGSSJ2cwwiGTJXmGHKKoKsroCB2yJpBd+ZX7Bi
5IL9bLQHYLrgHN20SFoHLKvelwVvqQE7PiHTRvPsW8Q1nw0nZuZD62yq+WYZaTbvByUc0ZQiFeRB
/YL3NZB6uRVMSVw6DAfVUpZFM9dWgpNM3lBbiJoU+raGTTYeysSGtLsqEk6TCmfvCQ2ApJWlIrw4
qvBo4/7YwOsXv+zdUG7l/3pUX02ge9gITVBETgTCOkdCPnCD6QOO/f3EQxw+N/px6lcgbIzQkN03
4VlJks/7yP0+IZQpdhg7McjysQ9YZT4YXSwbJSoEQ97NNKzHO1l1YOJ+PJp51tw7VhV98nEcQnRj
I/szIMrJbC7+mfjNNEl8tiWxmihUi66jSiGRsps/XxF2lsZP2qyMAuIKG1wdZixykRZ+DpxDrJBL
+FMWjphyg+oMWXZOPT27Z0k5sJijQXWaw0Av/2wkitBVx9uVgb4k5KySDmA2SUPSO8vm0YvRQz+1
Hv+U2OghyxPRyAS0UWYHPdOMpeGtiPHc77VtbAXDPDmaRnW4Ium/zmPnF+YNeCvLXSuOvHaenjv4
G0nNAaHreVHuBTyuv58Ogo26rSJrh7hJh2kzUJD2E/KLKJXT6tMKR3ziu4GW+fNFOhgOUl1flz3K
d+EaV7wbSY6TfhbkvQHGOtU9d6BnWrlyls5ZOb+ppFkfrm/+MuGPLCRnQr1mtouU6TfziAaeW1eb
ud0L/A0P5wcqomq7vnc00a8fzWOHLp+M2xYf2GMEXHlmCngZIhR11K8sPTcCQbH8ZGcuOnSGT/8I
juXKm/2JEtHiPbZ4w2vYFDiObli3x6a3xzyUZgp43WVH+M7pb5LFjur3JHhablgYwY4NFDuqmj1M
qn4t+cHJJ+pKFn6HfPIlH9LIHwJ9T31afrz7qT0tNsy5N+5mqKWznE8RCQ88wJ9ZWofjPlE3GKpA
pvj9244KFZiD67jMO+IbRYOhMNttvjkbjmuZUbl1eoCPT2xfbz7MQYLRomfCutN26xk5nSGyeMqA
SQFVizHmVcOVFDxePcvlXYY7JWJLgWRjN/SpG7NubZEB4xKN9MZc/Dd2bOZNJWnc17SXWCTYwdJz
HsE/NW9Au4BixdBD8ggbwtxz7bNnDPYCShZpbVv+hDT0sJW4jiI29i401h23VjZqwBV1cLr0WHbn
UNVOgef+/s0htokoAM/UJsrcckm+9GmPT3nweVRLX1irh4Y7ZNg6FBlyRwbBMIV/gGQcTOL3NJGh
C8Cyf1SNSBW+4V1SchJp3p7hXw4wVySdm1jbWwtHa9wR+kDomPmZM3zBeTdysUvbVwMIYBsVPwGL
v0ijT+BC81I/mM2lnpKjL/hZtgruNybVJSOwQGX7aEYBy+wif5tQj10lvNUqW5jLM6jB4/9AML26
1b4m/SGi23dYEnAj/egv9d7RuojazW540cFQtxKgHhIfdPUhL0n+J1Toj3qnLNy+tlGkxzDAUPh3
7KZTzBA//ZrY0aY4E7Wz63g0zMUedG4ZBCFmuJV9v+HHI7SnC28RYKDjUdH//YIlIIp/KZXWNVgJ
1RbvLNZepaE4IvVe2VmqcOY7ldaDS6MtnPWymnX7MpmtgyGcNzhpx4WWRBiOtSUrYB3JSwW7V1SN
7/JHm71f89Gr+Iirul/NBzZWhd231K7ZPfMSNrWSFDh/bgSPJ1qw3ochVocABs+MLEJ862UDbPKd
unaow2BZyExpakve+DmshiIxyHXBXFOBOW9g6IrXF+8bVChyHJT+Psbm5tz2mXMelvuuEn9Yrxq7
sTGYNdFmylbpOIpt5e1krHjdk1jaRhiXNohbJkhYT2Ng1WKgQr9TwkzsFWxhKR1+s2/7SpC908lG
KAJkH2+xDRAgKHYD4MBC/djglcV8Q6MqI6OOGI65jK6NqSy0T1BGCJOtAN1f7ggWfwv2a8Xn0zq9
hQhYKVHO5u3ZFRGVqrRQjFgboaz703MXaKkDNOJ+0JVYLraxm9/RbqwTF3cRXVmGpO3OjdJAud/y
q86XW9ufty9uD6uBbmufenKCjQZewpgq3ttT15vMZCLt7NsZ7jasmn7AFMYcLLcK2CBdsIQxKTgm
+8YPIRCxoslL83WoqA5qXfqNrLoSXQgdSF1hbQT+71mF+cQoJLikWMQ1k6Z+/uqGDz+k4BwuxlB+
fUfCyEe/7CS1tJOke6EjQy+Oq9yg/xF+d62YmETj9qlk1WEWY9/0L9q2CRu1a25KRrSrPzosSFxC
FZcDR2uoJqG17GFvh8vROfMfJRv6uZyxdUH+/DzHWcAmRca+JEyYF9k8RuNzgN3Oj7XD095SfZGd
PEMy2L3omv3fIIEu8cHJgMouR24RhzWHy/B/MJdraf9+XW5ZzyLHtgmZmflp/4V+kewFJKMplsEa
nU212KBhmHnv3q/ZbzFHRwl2ZfOshyiaqnEBqCHw4ppZ1Dy5yCP6Cqyl3She//xPzluBTUIqTg4V
M4PRg5TkC73nfbP4MAn2OQTwZEgbKKRFAKOuYPQ7KNmpTDyrsoF8AVxKneLe6uRSagFVCdQHjRW8
c6OelwQF5iZ3A9DeQllv2PLwELLvsQpQbzFROUlhEGWBnAV80H9tN9uLdM1rP9DCxB5g5gXcy/Gq
KY0mx7FlHx0Lw0yo3s6ocVY0GLfbyQ9T4IngdlYrBQPBJ4Hy+/97LmZA0pu12Bbel20OWPi2eBXu
lINdkTyOalXfbNVjYk+b538a45/NPysIjgOyDrjW5x687fcVAZu/Vd+urKQgtulQsWHS/v/zE0+K
jdg9lFbxrElAX/gagjVhtMPDRIJ9QjAmgZ9WpcWFO7CNy9PhzJ1hOFqEfR5f7201QlaQKMLOt2JM
vTzR5m6E/OCsWQ0r+A0gk+DwHauWuUS3vmy9+GnslYR8fbsM0Wh2w/ch1jy/82wGUZnN0cAIK4Ox
6f39KNf+Jha4yJEZVpWK5ll+yTYQkphPy4UGqxSoqypZ5g867rIui3IpD8KbmaFw9blj6hY1O23H
isTxTM8/r/1U0orGkrQlY1cs7OSKIyPQ9yIZatqOhdelTEPcZC3+It3+8zbvDt17CY06tgR/cMK3
h2WJoBRMf/ZxJQ9ZT+kDN48YuK2NcWy1xJOJZarjFo72IaM1fD5cWTM5Cnx1YmxjD3n1wiRynHAt
ZwW5PBEv2JSzZcCc5yUZNn45b364pJFJqqXjCGQRfzuy0+9chAO4Q/j4nsaIdZWb4wZ55mAqjVif
0CTPIBiAVtFhdxrEhtF1XMO9+eAD2APxf6TCcptUoFAG7a44vvXteV/jYAF/pBfsj+qgZruQVKxb
u1hjjmMoaDJ0ec+XAJi1CPC+XGn4CrkX1bkWGlO/g3z4+1VlC7MBb88hD2XQ8Z4Ip3acwk+NdjW6
oiEVTci9Pa2WuHol1Yx5JRz3jhQpCtpNFiRHFtoKPWSj2XPFtILbLe+EudhlLC07sy3lPkGQIRWE
4b8lhuZgxDAWCXr3zxlExW0S5i4A3gNu1F5iajWGRJAxIpEkXHw2UTsQ8BBAQN//D5Do/hpkLr8O
5ofcmbNLeFGaf8N48wpphrlqlL4wq7b0k7mJV0d3GZxnKNelRbWDMQwVoU93er6zFd2fCbd7OhSp
F6oFpABkyeXqYzcF7jZbLXoNl4Ek4hzSsZhEg+2gJ0pq3c0sSQRPxmMVyXvv7kEm3AnbUTFy/xX8
9FbbU0JKZZqDVE5o/2370NJj/keAHcC5gx0BwJfa43Vax3qeHgUEOrtWC6x6WF9ZHq9pu778pwfx
ABAbhJbRFPw8NlVh92+8ZeZi+mE4/JMkrqxry6xU2kn4ajlY8xAKLSljyMqXcspmUQ46PvRg/xYn
YO60jW5dWCIx6x8/kEzDd95PUmg8LkbsmSZRszpzn/oYaB0eVYmYDgXYKaoKErKUDo7p/J9tXaVg
ck6p2VSD/WB+q1kYWij2c6QBKEfz88/F4+gr5WXvFju7mWgSjkhkkURDzytSgxbbRkjTb08OI0Hb
NUvqCl2rRVk8ZUj/Gn4/tdc1ZPIcnQfT8eXwNvjtEnWjziDzmWEMqzMOP37xwupfM+mQuoOaAGjd
YKHK+Sml2fIGveJuOZWHfOy0QAcBY0grGOEEj+v++5gTdIgq2NHK9t6bNAAx2L2pKuxM+DHih5k3
5X4xVrzAU1PIkN78q89QxYdxrWJWroVingayv+A5lcFzCHBYjwU7IG3DHO2LExYdIf/b6a18DCK2
15+/SawtYq4J+3dy4oI+uV0RRHHQ1sOmeuNsM4+PrY78ToTQMxZLKGrePVA6JqMuGsKTBhRALsmv
3c/PiI+iRQsX+4c+9Uchd0QvCXQc5j1nt6cjuMIDuJ7U2DPUZgork0O704IW25UKufmZZ7QDtSB1
ARKm6KE+oqZtyOkJKh4PNG0fe5oleIJgN2aSdZvNkoH0S2sR700u91+R9zy7dFT6VZ+wYPTIkfGw
fS+UbUtyDyGKHicbJVEACIebiI/E8+mjC6QGa471J3627+sYtZ+Gi/L3VSR7DGQT/mex+tLlSRLx
nTnPoVVktQJofTC0BtMyCqkl0pDe8FZ3Dxjr4F4cGi7Ozmv8WQTAol9GBjZJ+H9OFXcqrkymTFlu
7L08JLa/HHbAqPzuKVDNzDiFv/JNQU2Ec/dJ//z+yo35Um2/VyY8r6iY52hyaGNIOAAIZDRZOHu6
1ueAm0YfEfv+1gGMaYgz1h3YtCWX/YksJN75TGu67HCBv5SgxcbhBa9eGL/e6BhlBm2lX/Qq971b
sEbdrPO+7afzXKDXvlaseCntpovO+Lo3kFJx0kYdVtm2tr/U7dBD9Th4FB3Hq8gr5OwjJBEN+gK+
zUsU8cmy0ql6/ejgVQCxLJuchFwGWZ3C2ToIsPgQP1byRVBvZaokpglm/U2h1lMcVp/SsFuIis2q
6XXugIQ2Lc6u3DE9jZBHIlZ+fpBO75VgYMOlGWAjo/l5guR00Y5xyky7cxTvIVFgG5ujJTA30DJe
ObNqZ4BN8A5++rOSYQR8ewcnXUE8GUcFVhnVctNR1sh+aDAaHKN/YIB60npOxLQ1bGpRcT2gsiNK
x3juL3kX7J5v8xKeyTSmHvCDK0VsVe4qM/5Yn9NVta6OvqlAVY4USyZpkIFr8oknMPhzWuTB6+gZ
bjgLwNXnXbpxAFWtQUxXzX40VLqxogn9aBXTMA51+gc9VsAo9prZgrWAoKZS7B1s5HN12OHpM7Oe
tXHNice45hyoXkZM9kHcn/vggiCHq98ZazSZtg78VR+siZk7ik9yl95VOj/i+H/OBqloqMVqEBFy
YUSaFYLbF+/yFwmAttFzz6qfFzYVxa9OkQ9/QLSTpM3L4dGWkAcDy1Mw9cSU9X0Ule6QTOnI+Amj
fLfAV1bPhLr1cdM2nkIfLtzOY5sDbtkCPZJqeREKRWaC/h6hQ8+I72nsY0McThR2at673EQKewsR
Qt82VAfBAwQgZbJVJvtD8s/qr2f6MUlWosCdkAk1Hk0+jwWMUykt2XfoIlMVUQO48T42KKvUBWxf
Os/VUG1HhFpTGzCV0O8tQoJLom/KqcdBihTD6xoROBRttLE9qmq/F0uBktCfjpazPyHAaSb9QAhT
JqPJZeDglDvWfoLyGawIkK0h0R/JHY39QdxrYkndlcWIeBt70t/Oxj+Kxq3Iw6AViD3fIUQdTmAx
rj5+78pa3EpCbMx+NhiX46Y9v1b9F4SsdOt+M+RtOj/vKmy7i+qEmo/WzF6ydgw8XzprYa+VHFkg
gfQULXJGbQN8Y5r4RHDlUawmyqjCKfMQTK5rscZufFsQlJ+B45RyUIcZN2mqgwzqbF445R3NnaJT
SpJj+ujw49/AdLT2LL2EWUBzr7ygITu1wZE6ewBSakrh9tl6LAJr5BN7pN9oPSM+nWnn+CpniIKp
8jfYzoDg7JxaG45AoEiYS9cAX4yLNYV0nXPie1p7F6Isq/GuUgvHWLthfjt9TWWRYxONlio8OpbR
NUve4q1bsnF7uQTIbI2vdKPtudtJKG4eTLmHkBqTtsIs/Xc/wLQsn/ZHR9kbTTbEEwZaY02BRw4i
wBSdzbzZJ99nHZ502ak1IVqn8wwbmps9jSnrL7HNtgiVMKh2YYYWZj3BmZKerL7jgmHzSJGNqwNp
QXbQG+BVw+/Mwn8rKfkwUiHs0AhA1DUgdOAYG+5rfxEgAhQ3srRZ1wSLQ4pjzXdVTBwKWGCwHWcF
YaPOGCabKIOqkUVRMWzqFG1N0u1yRmFbxlIdJC+9V5VG/AjFBibliZrdDRU/xHH1AJotfUvGuXQG
MFSfxElWKQ4PfZnq90Y2gse87Vah2iVmJmByi1hR7IyZn+kDVErnLz5Zjj0/RssXPGlEQJuHZZpn
Vxr8JisvvlErtfrW6LfHBgZ74sXdAKle0/OSTX/hagGka0pGcctPq4cpKyMGngK7OPj3AbNDC2Ht
DxrcTgCNtEeNU4uikiH1LWDY8KqLD7OuWz/MLdpwl/NAgZu58RhgsYMmm9j6euG8jTOeFbmSk+r9
pZoP1KjPIMGEY2OzDvSFPMPpFH6eXtoVTxwwKEZXVifpgC4usLit/+KTof6FHG0HFSnb5+GiFC/n
l/ZVTzCA+R7sfYDocbnWtnzQBzzoPZgn8HbkY5YMGmXAN/94LznOsKNH8FGA4izfYKbQd/zk5rc7
gkP+ciOfkASnAXI3UihZfPVfbuqG6gxBCU6Vlzxk5ITlYhI+7+bJNUDZldbuU0aFg6KglKbE2KRy
YRT41wNZjYwtpHNQwBSMVTABsGfcCcAHPLe6fFyCd0Ieow5elC1BbPWu69QS+hBI2WtV0JctCTWz
EJXmXYQ1aNzd1PWjY71pySGgyz9W3qgCTrZ1lqtegI2x2H0RnjCa7OnJMT1R2OR9xdQUTIxGs01G
oKbrXTEVtlQyWDZDEr/Z2LMDQ7EfTuoTj2Y9X8u9qb+bcCzRC4sqCEgUap3E166q9oFjhQEzAwSR
xTncsAm7/jjq4/MJUh8UXUjY4mmhklt5ruXbfYV8atRGcNLn8vu9L8GPPnaYFXetd3VN7fZ/I8RH
ZH9CVmwbgpopficc/pOMJeLneXrY8NhUfmHazqJIJ/Fehrw2Ah3ij46bUN/1763zYnTtyfSgGpcA
sCDmXocxAq5ASDM7bG/UtKWWLLurJfK1isBC0xGpwp6KXAdWvD1sg54MWW3lXOQkrjlpPagzOYiF
v46rub9bI5fy54q3IKkZq5/jSvPvxd2ImSEoveV1lsNrT8Oqo5wXzG9plCyJqz8BB6HoZ265Wojz
HXF2RIa1YM+n/VH3xA4Y3QkmthZCWXZvbrsTMEQK3M3uvfPbiHYgW1AfmgOYW4L+Tq0I3g/VkJu9
acQ5CvqT7BRHDedCRax+BOojUO7aRxkK8lN1xK8ZRG+gzxC9tD3zYWX2WR12SoYXiOnHAkU+u0yx
4ot7iEPP+2MjpqiRz10GXKCedGpm1DuqMZkeF5n5QhrVm7tikU8K2qEeZ4PISEHK73nTyqhdKjpf
KXL1EBGTjVjD8bv7Bttfl6Y+sCocCVAny8hrwVHFpv4bwoflr8TIvnEP1w+lvkfmbaFDIhCcI9ix
byXUeMYZt+AqvYlyJvaqHD1gmCb+0wMs+tld3OjaKBXXoU5pLinb3XOKTo2bSI/zIkNLyinAHKes
LKK1ihtgATXOHvSBdrn75RFhAKaW3yJv2diECJQYzdjMwsiNgB39tuEmAy1Cxj2lhXXdGEQS36FX
BL0X5ypzK7XI7nQk/WdYQBA5YXBuddzrf9CB0Vr4mkf6nC+bLhRNW3C6uWOg1jceLFzpF7FZTb8e
MvH2J5ufiGQw3yIvoq1Gv0BbiERKhuXCuhQy+emUuPXRNGw29B8ylKhRHkOrPP32mkCJMCd6fz+b
KEHgy6k7fitGwg8wcnyngVH2fhGyRsmIhIAwBRzvTHM7BCe/cGmY5PiJdmeI23ANVCULVt3BjDSF
NplQLI2Ag27fo4KIkNsrtN4ycUK54drx/ZkYAD4y390U8sqtVeOnPRzbPSDJMqYNqFo+1kppptTm
WYDaNOIvWyjJ7ZqlcoTAJnh35v2R+e0fXfXIbLE6B2EVMC7Lt+lym2aGNans8juNtsd4p6UO9SYc
r3GGKmM+14Ut1yMqL+LF6w29hrv8025RPTNiNIsKtgqmE/mfgwDWDmr+M8odqsiZ+FQw9iptxU7f
HMu46QDKUST3m2YxyP6cINvV0ZCMVoS4miSwczZBooqWYOyGQGH5Cf7s7XEp6qhMOe7z0d/JPAy2
Xln8ntzIoj/JLHIogpfN3lwhp4IkBbyDcDfWyROKe7tVR5EFD5/abKRfE/Dz0QUgocpiGkMpiw/a
xzKEc6FpZiE/30RQUcVIjKFSgjExHos2ItaXMvZu4gQioycvfY9xs64Fkk2I/Bdib0aF398VWV+Z
pX1jGzSwHUwp395NCd2xgDXnbBMhrRQxfmDTabJIKXehjq7Lxrn9KfBmQcgnhnktiGJ84mEq2/Kv
Fs5/nZkHg2oU46W0SZ3fZZqFoUT1KIpk+j74I5emgLcdd2mxxPfe6hYSpKq51cblJuBZWcmpwGFy
R07hJ+jja+EZVs1yb/bIjEa4zBzfqXsPSJDRYIjTtz7FLUfYD0uwKqqDiJr9OS9t+hsYW+piGBQU
dHvJaq5F184OJicw8uKVnRVHcMPRHcmpptwid4PyRPu6WTQA2k9PQGV40tFWvSgFnoLbmchDKvpU
iWtjo1FVWB6rqDZzEX38nntWWuOMMw96zzrBL42LR5dH1TiwiEQCK1hC6D/YMPWUVXcA0gMUgGRH
/2mT8o7ANPswirEj4ulJgJBOGQPN3/Ep3Bjmo1RsYcaKgVcbJkMwElBNJYt/mmEymB0CKkAzzOze
s2CAu3HxcxybbHB+Rwb1uTBhjdilDGePmvYv7QURYWENx/oAxCpjMFsxerxQ/3bT0UaC3WXmHWv9
qjEt9TxbaCDIZl/s/QObxWwq8TLIGPyGE0NbB5lamqRbG4u1f+5JQiKOSmWfJ9j9mGRMbo6dEgKB
kUcOFmAtXS+HSoXArTy5ntzLYzxxcA9a2i84E0X3p//WSZI9tGfqTfLS4XPXY0nL99VA455k5FBI
Fmc+bdFhrMfoPvG4khj6VTCBICotNN6IaaWpEkXmHCMpyBy26NSXnT5gBQRYbtNOGi6zryVcHLjy
leLS6mTos+2Vv8LdpYBvgqUzw8Q6VqATgkeaPFi6kwUR27fKV3//+UjyLHcC8c44rLQbDbX1rccZ
nYZ559+sADDsgLbzkfZIv3OGUpMW8iD7sei61pB3iiyBLuCrSDBK+vp/rdEgR6d3fgiIbcjs5zCq
BR1U+JBp0eIeps7f5eG5Yh3i1RclcAjTSjjN9posDD+2n8Hv1QIvjdVfQ3ZFSu1fHUgixZn85yDJ
CiWKGPzM0b4pzLvOkF8bP9DmS3IPlE3tjvBdZgsG8DDS2ZFCas4l+1Q4cD/gimtTLZVvSdBpST/f
9eM6I6Q9mAu1NgrZnm0l+1k/LeztfDrx4faPaGDXvPzDLfOSz0Jlg3YIa4G0W7Vn66naW+9sZCDY
VbiwO5TEYP9SN5SQbKRxuGrllE1r9ddBTxufk1G4HpkfuZWH0WroyE7SG9VGjMeYnxG57OagrujE
pPJeCasaRObDxRbm2B8ElalykdIcBKemmN3x0Eyh/Jt1rVO+n8HNV7EAqSol20r8dV21JJhFcv+d
aOPOFL9F+liw/8u6qiYrPrapT9gJ7irYzlnEmC0F6Ti1Su9keH9tBmnGZl10Sw82Omu7ypytffMs
H01YT+wfiaAbOUbP8Ep8zJ70pKr1F5ksr6IkxI9gyTg9YxF8xVYikOAzu11ap67Ft6+BTO82azYT
+993QYyCrvsvufXYqNnbKvCsiIa1w+YZfA42JwjGspohFZ/5NBO7BE5SHfLrAe48o9iOOYjGovTD
tPFJPefveRTQiiRsElqUjOrSIa/hjjkKNErr23nmIiJ+cf4njLUdkQG0FW/nE84hxeVIDTeVqGF7
NLAjdsaY7EMqIFfDdPkCmFegwRT+ZbSfobH8lW27ljtrGTerBPaMGPj4cDE9Jd2MVrwA/++PCxet
Ws0n6jIITF1zbs0M1YdbS16Qn937GqrRBiDgnBkNGZ0G7YL1Ln/CDQYYszrg+fWasxl3vWF4/QdW
Z+MFy9zEcxW5AXx2zgSyxpdWbow9J9HqK/hui5wCi1cIA9ucg36ti44OmBA2LOD+5XVsnip6kmfz
xdKhnh83RlyqVhkwe1B+DAOSFUE8BMMb8FTTTwX1gD25jbtUWgoi1L5C7OkUmLnTTR6K3jBhQL7D
t4DVitG3u08T8KREGMQhmpPo7MyEDHmvv0A32LHwarunIjn7HR7f5w8ch3zlOBpbuB8T9W3LNtmq
XuSLDPR7HXA9hMidDOKzwOhl3miSyyCrSdsCXxERCRt4pKBBKnIwlWdikZgvD4IZe5bVsLbluknY
3iqgI+wh/hvbjj0c7d9QBZozORnPKwtZokyZywlR3smB6UHl0qCEnPhNUf76lSUqytoGCK5uThdH
NNr0780BeVKtMYxcvwFeDUEkRifBLTRZMsa4DxKCDHmgJyHy29wkl0zhfZxeTjdp6kHI1Ej5Vqi+
umRT3K/4nqDCYebb+7jWcWPKAfGFbKN36ViXksEaqV2xMpU9cI5Q1s28HWEIKDmLFXwlFk7HsqE9
mvydUlYT3hBXjmN72xUn3XvAyTwP7I0SLmq7dXbCm0U1i35bXSBad0Okysb5G/yitX/NjaFj8S5s
BAor03tVsBreUssNDXT+deQXZqfPNH3MvuiqplRxzgkkpCxhEVvCW1iyBTJSbmOWS7mwfmd3xtgf
9cMEP84BS02L21QTpp74qSFm3VMY2C+O8CqdvIc3QwOjSzw2ldZeYBSSbu+4jWd7jgSbk7jCdjh4
lB6UNhc+ujSa0xBNy8lJe25AJtArhMTqaazUlnwiewt/Qed5dRnmAgBC/S5/czGGGpoZaEm4w1Nu
4xQVRqjhozvyQXnQok/EW0LAMFejX6m+wkRte0Sehs9tf9p6zS7TAE+60h9jRBCLfWSRLVyMT4Nw
xlnqFRwgk3mBRazKMByKJPxhCLZn0YnQN1Cwsm7SavP8VbeoHP0Ec7tsFw1mrPi2JrJeD+UOxwHa
ZglcIPS4fAfFe5gmUDjcK1IL4EY9kN3wbrVvNUfnlVRfpbXpf2J5VQbhnesU348jbp8Ar1yc7SNQ
inQaq7ljnBSaJ7qRd8IJ2XDn0V5dv/O2Suy//3ggf4M2cmVMbS01S/AhLb0xesCUb6QuHsphC6Xg
561OChAuW8pGckkrLCsUEBf+I0qqcWmUYWkfT5E2o2ONVkGAo0U/bfanJpP6CloS7+efQi/zug3O
0ZEBHOz4TDp7DsaGfsJg9ou8BsXUAKz8v0c3Q27OYTkYIciOWeV1pc1uxRFk/vZhl0NbJCKlC19X
qp5s/aN31QoLYqsHyP3UAnnZLtNXfnKpipS46poeCLGZ1PUw7bctT0dJvIoKQG3VoTuwTUedv0Ou
Kvn0nweSJYZicvI6JWPSCEzPNkPAh8AQiSifbcVnEXUhIXV1x51L6aMa9BN2bs3qlGENvSwef2db
VcSB7uj5Noj2wMixrDaQnviTb44SzjAD7PR+uqJgiAHKiNvHRM8njmSvPgVvaAzUGssT3iS+fOH4
RITO2S7ajlqitInkY/QGNaC6QsqHoPpiRrUAh7GuBIYjD9g6lhedT+qIQf6UjesVCtzY3kgWVOsf
6X7Mi4kAZ3LjJTxdbEFj93iSXQdA2QWD+zRw61RvA6+R9wS4phLQ3QXfDS24iUyH/PO+5DX8Pzha
URql859bWTKgzG/GAI00hGUZxvF85G3/js+EZwrfARTIZCzluUBdmz+oMHuUNplJIXvnCx0v74Eb
S1ND4qWeZfmu01dOQvDJPUqwSMoJf7GZ7zy9bB7Bn1upz5c0bJxOiab5oDgcKGB66dd6PWuuhqUm
dEAuot0uDfO5SkIBHiB3d/wfxQNZKLXPUBOz2ZO7m3pj2ndezQ4qGIyI9AKRIC72R0twabyZsDVl
bskFsd5sRb80CzAqGlW2pWbZ7J9MrrImT9BTHaQYyiybNBXCka8Y8ROXrZTHgOpU6cqJv0rPQOxx
q3TiW5KWJQwc+DFn8543ioN3Q0np2Q61vVhUyE/IW78XnSfK8m4spPgLgv5/4GmeyvCg6f/Eayi6
LhVpkPsGtmsLVDeLtaVkX10epBMOWdFhrGcBoNi4aK3p5ss96aZr5dbDGgY0TFuJR7A5HkWnOQO3
hYML537NrUh7bDFEq07zAvutQt3LcWTYLniYN/rd2zs0eH0ODi1Sa+keoPf4oydfXOfoN0NsSRrw
exU6+ilFJPJaDnAyYUICATnbsADrtEWBchoL18Z98YK5bpCXA5ZXxZvzv5YmBwM8bMqW3mVZxgUb
hZK2aPB88/1oMQd730AxlTAFhCAiOjjVMXMc1abSmlH70Sa8zOmCO2/ccLigiua3LckoI4F+Varz
zp6PJe04jkG5DIl4BNzbD1GZ6Df5ugDnpwUl+aPwU+5uuD4CqqjGfHvxUUMClhBKmqqItdAVVqLA
SJMuV9nV5hovrsNajnt37vbCbfltI4NbcgkaJP/Myz1SVvTQlVhE1TOGYyWAPz+Olz3bHvWPlvlR
DkFFbZKT/OIqXYttvsuOUoPZKDPjEJnrgWBaWyYOaZM6yfyj1le979jmG9rIUTKRmLynUSwUIErJ
DIDI6WDIASuY+k+RtDobU8c7FA5MSvxLO1r+Fkr1ZH+UawhvNMEkj80wio6oH9UT/qeofAzZxLAB
HY3SD8cKupqTIEzHJjAcvwXYIHtzmay3HTwtcOea+ivqJCJDRip6lKHS9xizbXCn40WAlNdEvTUb
mUVrXZN3zhY+F50bq+Ey2U/m1Pye7zZX5IjnnMiEimA9niqGKvr6X3yrIH5q/Xqfj8RNMM/gQHnx
IZLcSfeFp0xvPoQTdvQTZ9gN2DUh5ZNOtJ1idrjM7UKtXZc3Kg1gJBh11Vjtp8CaHFOWwqLjTGJz
Z8vSnN9EAmALIDae19fR2h9j0w4uhWGmvCGD9d7LPHWgnwAiY0wEPTz+tlx2mFbgtqzojgHDGeoH
AZa9A280BDqfmWZgsO8/EMvsdfaOduempQa15jI6EBPYk55tYpICNK6MwK8fBk+P2UhOE/FYsQHv
I1niLJ+dSoYYAeZeCso0URas5scMLgPswifM+TBFC6uXSC1hLS8bv8r4ArtANKXWC+0oqYl7Qzgg
JHOYwxuJZiAsLIR1E4e/ZlGnNW5Zm1LhuzqPcXvxrt7tZQqG3yNejVUXvenpTRn5+DOzleIfs+d7
XpGVoI2btM/KDcMgryy0/Frsc5oJdi/7w1vJrEO5no24I0EA+SXMu9CTQUZcQv5I6cAqaMJ/ii9F
+RyC+I3K8sIhWFr+NDeJWRIzydbBBdJrYWNqoShqazPEPU//WmHXcjxmXsOuyAijY9p3THCkxvSm
wxV6LNOWlpAR4O1eonX5jDhfRfm1Z0alP0UfndI63T2xlw4MMoM50JbO9BXOMiLIylbJBVTdxRe3
R0pQ0sGWjFdhSdUPvvQsHiuI+GPcpN6zp4XwF0GE0/ItlMVS/cCwzLe/AUBwLzAA6x+IqoPZ27t9
QqILX+M2IF2eb+VFFLvdMFlAOuYzjfJZiRv2bwazWdR04RW2BHK7oI3/G3VVk1m9e+42x0dOds3R
01i1BU6VTPOFbaboK+3RfllEWspfqfKUgfZnLljZ76uZp/eadXk3zk07eUzq2QTtb604yCvGpzfa
Bk3qXZfdBOJU+GK7HEaSVIA7cSNk4ah3gWAnrjuQ+QLXCJ6efzL9bnOKA34cLsYgU1MsYu98VVdz
T6pDySi+iwomFKEsZwj7uNBpgVhWXf7BJeYgj8WZpIpxI4gLsuAeodxAWIS48Ze1MCMxclNdQPN+
N16NkUNY2+nD/41kza5DSxHX4r7Xlhpw/i1TeGBxWo3l+ddTq0zdC2Rrj6XzzSK6E5TBVBdH8uh7
QztZyqsGBiagLyOjTqi76b488Y6iGONGyG+iLuIONnvAPWUwp9R5eKeqVL5zx68dF9gwupQnLCRY
mnpAa4KwxbRtMPRMoPx2SVYqi5Z8JAm/gDgmc/haaLK6Sf7xCH+g2rV+2GvL1DMkXkUI73dWxWOc
XbwGd2lDiqAjaM8eRkPTEfxYQGJNu5TtEDICG9B1IFzNqN57usXdr/ufIjwEUZKXXvp9siGkgH0K
evNbLGb+/hHx3fj6ljN3i9Nl9jVFd7QecQlqSnA+V/kWzHd2cn8FfnZE/1aMzOfO/wNfuGo+C1u+
4f206wPNgUpYW0Q6nUGOQ63uTI6vGtesNf3yCb4L4yTL8R5P6OOCbjObmOevmxghLVyr0ZTksLuH
Cy1G1ESD4X6+i04k2r9sr+p8PptE9aF3XCLuYH+ZRMFXsiBs313kAnJAx0qkdyGatQZeT5OL9Zbb
UX3nVB0MdtYvAxq5P30VOvfwgAmIFxoI0uKHIS/Ggwy3YHO2d3Z5sQaQ5wes+dxjCdGIfuITY3oR
UKibbpEZmVbhnZnRROAf+CteNM4CC8cudcO0Yl1lN+AKqSHPTBYXjOt2qlvImp/BmHs+FvL+v/Et
9YOvziMrKhgk4TFnDmfQn/mRxNptC5mu+35LniBuFqgFFxnNbbKl1JWVI2d+UUCRfyJdvVUl5+vQ
RwN+AlNJIGuZWjOvcEBLOdNRbqD43UuX7IMOoL/bviM/8CUoxYFV8cnNQ1VNAMJDtMyqum9UY1j7
YWnq8nMB431WqoSNMwdpfMSMKwyGAb8fdxWgy2weDnSQBLU+uUq2TGNv5rCY7rSVTdNu+TEAoOr2
byodYEjds/Z++FZjJd7AgJ+51IecLPI6oeIYUoWfpc1rTdiKN+4AuneQIVoo8s0J/MJIHvN/mpF/
h8mkq+Ar0U3xSz/d3IGCYEPSh48dzlzVB6aGqocBo5vU/Krn7yD0jKCrrdzmtF07P4BgOQSZ9Rex
z5m9HBl73SPk73Hi6fgpIDb63khlDNr4abI4Tb5ZNWvQgGFFZD7w87IUyx+AZpXtDazugXz798pK
R0XjThjNeWCPvypuW20l8m5vuE8RwAFPO2ggRYjhvy1BnoD+Kr4uoVP07r4US2BHkWXO8XcoXOkL
zSdEvrKC1AiiT4BqOwa8BaufWkkbPTPwhXpAjci0kAT+3lq7DoL8NIuB+918sgNrVegPDo5fhTaR
kvodQQYWS1Akk86gGui8rzyv54qUYkiB6bLXH9ug6qFwv+OEqF5gG2+OREHudv2Pq6DhNRhY3zlu
wYtSA2Np7NJZqsvBHs/5GlAVXt2xkorPakENHrvK5FMu2zz2ZbkFlGv7mqrZHuqXc8NR9z7WBqFD
l4PgBpY+BbkFDnv0TAg9qho2dRzEUI/+qvd7AV4dT85UX8eq3EwZWojhiRfmmi0uYFhIH/36hYZv
NKolCVjXWNBrnLGLC2OQEDScVzo+WMt2fsd8rayqbaaT8/fpVy/1dgw1vUBUznAGNHu7j1cXMp90
JRdPsx9SsvCesNPLGS1SjJQxPbyIEhJeW467S4HDsswNePkmtVOndOq7zf2kZHlb7BoTL6fQ1TMa
hg9M/pHwRgTo7y380QPauc8KyIZd1fxFb3Q86yRAgotQk/F2FxNqmAUH6C1gi5eXektEMjtegGnE
EzXYtOIdOcJFMvpNLdxD4gT0gRkuF+ZX83tbWi9qFGChTarDIYjvr9Rd6nzfBRODJljcckXhvAhU
qZRx53HAJcC8F3ZNx/JaGt97KzufTXkH5Sje3wdkTT+DhdV3XyVRcDxJmq8CltpVvvJk1riOswZo
Rlvbf7cqhoom3+uHgm4q9KhZpPHGkaA3BIAXn7mRxjIlwudfeho99T5t/vw8MMr0/On4rq8S6d9v
hQxIwE2HaWZQ91EyusYJ5NCJxAoWI4FwGYVslm5En2eq0TTdwCvMWjv4vfwYwWT/kX1ZVkOgyw3V
xtcHMBLZ53Z541L8pSIdlxGgB8MmLm2JbpQjUyNNnwt3Jm3FMv+QY4/moOzUayTpue5pkz07vqWi
hE9r359VFZQ3WqyOp8duB3gDchXn96Q5gy4BgqK9VEKnkYB0fWAO/FlnCwKhzL1IWK0n+z2v9AJh
lIOUFqk9nYwVISDm6Tyq0cLhIjo2O15Lf9jmCrQiNaSjz13VrEE6KUeLp53V2FUdiYauGYejAxI8
oOH9Z+XACPTn/642Gq2VueHwDouFJSXW/5oQ9WbEgJFUq09BlI+EwafH2YS6wpXChyyCUuTmLg2G
kyoSywISCdvl65CvOhB9+wwYxK+huVSkzTLCuRzuq4USlHHqLmJFhsQlzVsgqXFafVL2gBY3wLyq
6fbicUsqgKxPlHzMPpqrjZXaOlzGV/GYVaywTVK3OvkzonvfCBvXyDpnNQMNFjMWqINGl96hedfM
swGMmVRQ5FX/sB5ra/aa6XmfxqVAYvwSUqkTNDH0kJm3aIbrUjO9ul9m37mM9toUzEckJ5e2Fw/b
V/uZVnhPlC3TuBwuimWA+dlGiHVhct9jq/DqXGySh4og6cEKBdgXfhIlm9pmYBJxF6h0fMdeRW51
2nL6ScMlw1guFPOiSR92hE5u2aSKdVvyUAwdtgf6Oepj71kf++ALs8Z1lV1K6IdkCTrXHmYltTJ0
5TV4EtoLwdSFGjd0DJF/K7+sUGr8kXyeIROJG1iHsjT24LBLMR5Qr0A/HQQx/idZ8LY+wFgFUFEv
w7sSX/33SLND2kw1q28qyddekCd0F2HTh8LCyRySbi7MvTFgw5J9VkKo8mgw767GCr21p1jVKkci
VPdLNQuX0eEyS+uhPqF2jjt36TSAva5LTLm42OV/HD+cKCBuxB1LsroCduPB0oNFH4kdUeJ4wUgY
KmVoA9dTTW05g2cMcBEwC9wXOdnT9kOxXwbfiL6I56XINcuSRIsUqVqhIkKfyq83t3nVj7ntcWlN
I1SIXEtz6hXS42m455ANP7AH5O88lkMK9eL/9i3SZK/H2/8W7hQ4rG33TOyI+v0I3FPHEH6guSa9
z2U9RPc3RbSJZ8030EyaV5mxJFUccxcXZrmRO0PwGFyBTlo3vsyR6NGFa/GLshJEKWdPjXqDLw4D
sO8AQUS7bg2OLxdNRdMS2MT11+voInFuEBYlo+TX/LYqWlqMq1ey1DR585UQqkuKJDi8NNILItch
Xi2CEwSCkwXLvxKBc5jWUrfuq/qgmxvGc7BbfSexoT6f876e3UMWl99HPhBOKbh79ks5Wi3ZGMKe
exxfYQ8+/BbpSnwqRHmg+ybie5nMmMyYRjW9mlQVu3Wy6dD1ERqeJBOFww2sKMmBl/49n9no2rco
9QAoNC/1OfQT126LqQt3EQ9H9LdJ0zChJLdxShaVkfB/rcQ6i5/wiqOHi4TwMV1zVRvKo2chdE/8
Cgi36USi1t7zKqPivmPHOUZrQj5huTXVD3VatkJoYfHRUTU7ZinWukJf18FwT1zI7ZeN4ci21ZKG
ExbaAsesEMokjffvRGMaNPxY0G2rk6my9zEdZz4R5Uy+msXBOwdT8rXckRX/5yOM7gfyrg7eVmT2
YIWr/qNmiBR1s+BJcHwFfIYcQtAckttyiXzZAkp5Ml5lgPdvDZJZnGA4cAyAI9S0tLoQv4NKqmy1
E5A24rQHuSGnty/PPrDWPwHFw+UYThB//RE/cA5tbIG/j+YikoEu8hSVfeAytXuxFY9p0y6189ve
Y8LK/qiXGfac3g1WVYXTXEjPm0IfSkN15cS3R/1HHhxy5fj5AqCuWR0HZo8S12YXUnGUCe1U9qWb
Z/c41eVB9CZOkcZWW7m34ZXmRG2EgkQWFsvEnS3cXvgDciS69wRRX2muYU/JT1DNK7yjj5mXOu7G
ByyIOA5msS55WfbDFN7zyJVX09tu+UwmakiAN1ijx2G15oRjXkP6obTOb97Vg8ai0HR2sQYSYupO
sio5ECgdQvwCV1aNmBUqXj6TZz1WzeEoCzlKcmq5UBeKrzeKMZZu5QahyILjja4YsMx5Q7KkzryW
2f7aG+X8FiwyNwfrGZ6I8EKi5QtdcynlNP2qSoD0C4wNRATaQP89tIRaHN4sO7fjRKxLXnMbux14
gv9mPzkSpliBLdYWJiP4dQ8+TX9ARXCG4TKTKOwjKlHcYEdwG9SRZGhejnfVs+UIyJct+ge4hlFF
a1eKXDx1o+eDvWRGdYzXL9kVaE/KrTASRN5cgXMrln8SzhdIR2hOZbFkI7Rb+YiT5o74dfpeB7rb
69ed7xAh21DdwJtHxCi/ogdj3BteH1V4mv2QD+CGdaS+h/IjQTZ3eSJLS2s7fHvcz/5EYkOgzBRn
vE8kJHEOsXsD+YQuZ3lEM2nFkCrovBq7A6mJYQdImCQBCjzZujkMyjz9u6Wk1LX7WqS5oMi4V1g4
CHsxuiXwjMPM895VRyXu/o0CC98xpYH+FCJd4kJMRVpDIFrNxgNKnTJsEpJjqkNWWNulIM6dTXk4
qYYwqFO0YtNIA1ePwfUUdvMZvndT0R0JrMrwPLlMpyy+5TtaTSgpJetYEHNjLsYGyJTx4xR2wTF8
Fsbvprlec1ONjhWLJaQEYZX24yjmMXF5Gn+INkqcOgq60QEnSyZ5i7eTEg/1HvFckAS/ItYJrtF8
q+2uq01xPh9EKCwzc4LIqUkqed1DMZQC1A/I5w29sNABCafpQN9ZCeeKS1VCelhaMt4tM5jvosuv
wq6sKKZai6JiY+OfQAIqfUjORKlXDa5U/9R7FD4ELopv1tEsjdJufsNGM+aJA9CBn+5ON3IOAFnX
jQ03uH5RoRA2QS2HsuZqhEtMNdcMi3PPJhMK2hU0sk3W5KJ0bRktxxtvOeATgw8AQhXVoN0XpgYG
eEocBwFybpbn2xnSlfom5GDsHFl6k3rcWsPwFObFeLVE4J76KdJAqiax2WissM+nKgIfxL44gpwR
FaaFeOHRLm/rqd5ywToz0KJ1L58JXUYsKKspKu4Wt4DSh6NNENHV1TBLVR+Msg7sxxRdgJbURZFB
8T+bGQKhhVejU0tdiuxZOiU4Jjzmh5TzODNmVGc3H/88n41fYcDzF4fYvSWQeDsXJYDK10YsiH45
ExVyobiCjPi1VKFIOP6wjQCtRvOSRHFbmT0u51eNkSfvfGnxPEm+bLkbrofO9gor3tSU2iVc7es3
eh2COnhjM4wJhs1QpqnqLz2nDS2vVcIkgpQqHQ+jS8Bp2cAMXnOPfCefRLq6bKQ1k/cu/ZPJIACy
KZ60V3FPvJa6j7nDgMXHmlZ+cx3N909reE/wBwm05lsr7q7T+TxKV6iJ1cR4UnQCiIbyOtP89AfI
881DJ3VLKDlOcgBnqEUv3raRId2gT8jPft56hMehGtvqf7W1CRfa7OHC3HVVnbIsA+q7HwFI+opf
KVx/kCrIUI2V7bgpjUfqgz2ikwFerZq05vEf1/bj6fepsymH9uqfU8S+pkG1DT6AJK8Pl1lmziGF
BGOQ8ntT9rC8q2aQMFl/5/x5qyPqRbe80C0EepXgYJhgrxrj31Dij/aEHm7TWDT5MVUUDFeIf0Ob
R4zFroYlWvoOZzCP9Gv+vXMrwYJPjQLr44M9fE+R7mM6ikVlDfp9UPL1V/04YxY1hCkhuwhqKchQ
eu4WxUdGUyaYxnb7XEN5lnQZ8Y+eGK+UNaDJE4YAHss0kfdiHRYZxtquULtJeMV57osIWi+1+bO4
9zVaSFusyqjxwJgsvPDaHwzd/Yup6hvtPgvH1l7vKhYwRN3YrahglVQdD91ny33jXm8w/b15ViGs
NBym+ogLXm9sVqhpN4yD4E4bb4w2is87FyyvQQ3WeI59ViJAYjOZOtIcNrAyyTtvy41rtLPLwHIQ
0by7owbAZsnOMuSQC0rxuci7DoLGKmpHDKBgNfESLMhXiM2bzXDSPmEQQ1AMt4hXHWTzsNSGW8sI
MBNVZ8jG5bCTgtwPNT5e9W/cTGHGezzKtpHpHGkb5CwL5gqA/4QabdJ+KWJH01PZmvV1tgKnazsZ
jXx6t5fis77bXzfkwUhsE6JUgDANcYcWh9j8aS8MowwO6FhODCZs2KLTDNXsOE5CMNnbS3IRb6Ba
ciegrZhhqXSSShR995keQful4/rnwe/GnYcktes+a1K3Su8qaGnx3mXyRtOzmbYLSVuBTG/ShJpO
XPIwWWIdBUX67XMhBa+czUuU3gGLpEFhx7dbndbf+Y1peA3UBN/sPmi5Eq4TDEsVCKK1yD/oLz+H
A0qcB4U2lQVBew5GhMA4KjbP11GiLXJCfOvL1K2mOOzT75kJYsOtvZpnwYffE/+Rk8uv12whq8kn
b/9bW34WQxUGEaZ4tZZaxdCrYbdU65uONC8VEjkyOlDDNHEmfCmVormD4vCIoYmwlFVIIkFE9DBA
q4BvT5G6v+36AQKIN26vkJEjVKsEa4gfpGsDANOk5j5t8IL2NkY5ID/kEUpb7csADDU8osjntt6/
+TdplMREOjN6hhDuvtFOVyD3nKA8NO+cRv/LBwodoM1jc5CAkI2+KQbovLROwZ2bVR0/CY/SezLA
WXJZJ5E+EGoBku7zjA2M9HeKKlwSIDHwKNeMjMaG0xxwHIhaTGDjTQzYtNqT82ODZsqaJBe4UPVj
Q1DZS1Tlu5DldTumtFYYPMs4rIdVHz+EaH/hRf/2PboXuzEHrzd4btir04p4AttJ6g82zzpfn4KK
kx/IkjrcxlReC9yLJWEhkkqPqF+Gt1yh+CaP+CTxbGhkVW4MIUBZxdwcULny0jhK7w3atq+k7OGZ
Qcec3H2H0wlboJepvNQOcaMvfqIBYh2k7xhNyQ9vkbfLTiRgEppS/ladZv5QSRvPPZkZ+4KatrH6
VisgZgkFcpTubjL0IxhlxGsQbs14swX8SSylOZp3asBQepbMS5y3ngZ3L/Vkc6PCFfQTSlk4NRmy
xxtcJ2iM5jzoorOs7lvPFAR/ok5ylcN0RN6RWpmzmoSCo5R40DHw1NNY5tKAs0r+VlzQKhGZqydF
isGXHoIUm3UvPyziFjK/qF4jUexu/ghhjv647suOMGhbYL/yPuWGjEK2RhMvyZZcnVZMkNIxNbNV
jc4K6GszEBKsEPCpXTtLaTHf19g+zr24hACP0e5UnpbHWHXgGrVw0K2g/43rddRd7itdcpyy47jr
+BL7oHYs9tufEQqup+I0EyFxi7mcSH0pwZSX5XXR7Y8s9qUcy6b+ccOtfJsY8F2AtjCGx44b07Y9
Pr2uDWbpgFh9/Wdt5ZsgWcYCaVIJoP9PhtvBg0BSiaxHDe0i23xPndUMCZd4BjZXOPX60XtM8PO9
L10ML/gpAu55b7CIztwyjbD7DJgBtaOK7jwX/y+rt8+p9xxBrZxXWRPqL8OOzXdklO+Oo1ZKip1+
BcakdgyCrZAZtsOiPBSDfFsbcjjsShV2DVtgEPahtZwqDLeNq6eWP9VQsY7MfPKoceVVfVHcVvui
n/U5A/ePCegdbnjviDNwcYRSlWlKn48Du0fpKRhODbG+JVyo70Z+byeKhudaKTnKm5wWUrOacgIC
YKjF34CginI2Sls6JSjnv6xPa63os31WQ2k8ndRx/tk+xaWqbua2m6Eaz0dUrpT79Y8xZ2N0FHLq
ZQQHqRzMfwXLSorAJFhSI9U/WEDi7bDa1SKwpkTHYyodJ4fgFz6uC1S58ZmGqFqkhJNtcbFP8dyo
AnIOXnnmzohWsZbUbijF2lo9Sj1sPoR0g65+tmO6Vvz4lOH3P1Y16lgkn8yWRezKGlkOHU5Aa141
FABB59FIEs/WNlk5nXvRjirQE6oQBzLJSGzHldS0HHOfFIehdGwGUFKut6gCyEFplnCIahCi2D3P
ZLAS6BQ2qg/8Y8H8CoWO0nsYc1CZHxozJoB9YUFkNF2s9wUqe3+Tt/XnbKOHOC/cehIQ0wXMRKn5
mLYZNlGyX5WpBBiI5IkhdF74Gu4iUpHUk/AJQUP/68T1zdLphxOgpudz+IVRK9V0ffie9oIG9zwp
yUOqraTMRrOKq8OVO2x+KhP5Msr8SiqgPRsu9Xn3LdGBar7PALAjmC30Dt0IFPBSTO/akQX3SXH1
0UfnOVa07raW/J9E02JuOtQ+2RjzddypYCNJhnHtqVEhUw/vxajoi566WS0TXY1500WL96nGaqXU
qFEOKcxPHGjgXYJzyP/dRrMssIbPorDNSpLfdZRbREF/ZgZRTxDvK7kGarbHIjsuBsJBIDkKtZty
eaRKx8hmUcCt9e8w20xq3XmKIPRYq+lOG00bM8BTo8LWhY7hK+YjuNv1Z1pni/UnM6OJRb2CxNK+
HCfedg9kzYobpUIV1HpBIiP50R9URgnYrf9trN6sl1YnhfH0NJLbwuEvE7W++i0QXxFWVwoV3F63
JqYMpKLm2tuzhyWzR8U81gwUEbmmYi9Ir6IAKgy3Qr1dwVHoC4Jzhn1pDDGB+6a+v35kH4gsEC6b
jEzsw2CF9QAiUF5isb42i/2bJn7y6/m07V0xLsIWNU+55eso58FzwrYkhqYPTTp6rOmfRVgyVCOQ
svTg1BLv6nJVUfzapQiyFKVdv4jDIcroOs5WFJ7cwIjyWy9F+7eNy/7XbH3arZ6WaK4X0CYpKoc5
uE1aKPyeCJm4DAEB43t97NTqAiFJlFaPScC5zi0KVDWuCWNgrjptKxxVL1CjG5CqRds4qy9ohqqm
VD7yT9NCRTIMTrzMD5bFrl4iiqMyVMakzq+G3cMgoP1GiHP6HFsZnUMLIb4/cCpP36lozCmqobyR
/in/XmFpBPIcjtMcRiahHJQQZfN6rCGVoxZuInJjOFhOaz0bL/9Dj1OApbCupEkamJGs0aiuHnX5
irS6ebiodiLPTm6x4GKHndTapmRQcmS24ZCvVv49TiZ+Z8Ms8CpgSH6gQvs/o0KT2PvANndM/16d
ArTaAPIbo1ImcJDJvf19XL1D02nobOpEYqNeaAWzGix6lDtT5+bufss3mS2wkO5mcY7IaOsHbSki
EBBU0nwOAhPqVUpbqm9nx5qNJUf0Z0nidjW8ZBUxGGh0EuBqSxeNYv0MPqR8umIqvO9gmBuecZqC
mh/8BXSRf5gH80RnqoascTNXquuseJFVST8vwtmfmcFlUZZG6LJV3QTuqA5v0PGvir8U7EnujmSc
YqpFECBtOWLbh9f+GykDiZY+glwfdwGiLuAlbhyfZ+oNSSrXpy8FlJcXbj1PO5DJpeG1Q9UY0uLC
4iN/61ZmCrwE9EPmmIxYyMvi4PEjm0TXq+m21lcAV0SUgSRjVbZ3TEMS6+8XopSY9AW2N+mWXgLr
Ye2x0AnjuMcwVPjlo372Y6+MP8fEOfk0RJwHPdBnlILCgVc222XbWhZpKPuLoQ9zSfRKKYBI+M3R
uZPbUjVttZ+eUW87zIER7RMl6wtQU9Lk1Lr+TQr1UbKkV4deMXgucPX0nPRg5+uoEOv1DgXqCt25
tF6HF/yWujK2TN3stuQZ1fKrVElh2EHTjeT5q95rvx6tms+lVgNsVb157krbXlmoQb4giaRWh2+l
a9cEmjobinwwvrW4+BYMdz5aueY0IPRa1FdI/8MUM2A302psKz52UGgLLDAdGMG5Ld5eivshI+8r
swVXDpq0eambR8SEmCi2z0FD+oPJw8uNyVL1FDR9gZ9SKHNPH0Y+0bdbMY2eLZ5zsM8I0dsu5hNI
uDApgSNRRD914/Ezot6RM8gae03wTYoU3+o/teeTXHdZYStqKCp3MLkFaHl9YjArFZuOi0GeItjl
4HS6mXubfNcHGk9oyDDnwo6Rn8aXDKEqd/FVER5a9w7C+mtZmaufnZg5MrAqSiyfUg3cHlPsR5if
N+HFGkPvqMCPGeUfEJSBqcJxLHvDGJ5Gfh/vEswcJZILt/OPPNzRnOqYPNBzohFzbXhn4ggcw+e5
G4kai89VkKwvt7zzJl+jyauOoOD6xJYhFouD56msOkgYN9khhK5WmNLxecbVfpk0GKk9+YRTKZOT
ctmymgonXjpvIqMYGwxw7CdgH5w0AK0/xQdOG4TlqULg4MNr9Qo7Gj2USuujiTawXKXJVsPlLp4c
IdT5TeVW7mHpF/K0hV1EcYEOm1/ta8/9LTqSdGBnhSmNNqV8VBuDAawqorMS38PInHjPyjkm4+qt
nGZtqBBJih4eHhpdXDMPl7R5JhhSjR7sKn6xgYtwPa3xluTaWtWuR4w5I3/WCam7DHlc6OaNmMYk
4RW809ZlUeejNCljM5c4HiSiMxXVT2esB6o0SCVcPx3kWUsoRKk2ZDPWMMTE3asQxIjDVrPkGwxc
znelvcedcalD0pik466Mh39FODTJxjdz8BtwUoR6n9eQj9dhyFe+bz1qkWzJDm9Dk6uMb8AkyPNI
GUIkzoaBCcelo0UMDnj8XGW7VVSZrEcg67YgYBpBVBj5iSBUiFUKJ0L7OHFnagiDyeB6/7kbp1VY
qqu5RI5cvEBYsGvCzTHiAHUZX1Jg1zigb/r/GtaudmBmoUnwUpP8UOAiMcTHW4bWO1pE7k9jvLLr
zznIrl0Q4RWEG9amyyfJU4DknMQx4Zxj+ChRNtvkDUBzcnh1e7KHIoqT79n8OlKVPQqaVCEwb/u5
pkIiLYkeNHB6zsY4hY9tJoRQ+bA1SElFBjkK2vMdmTSkBbgFkGwTcEOEWdpUhytJUpmnpiuKejWY
gewpp9SyuJTMYXg7Gt6TALL95assTE6y2v05dMUe7Tq7bpbE/jesMD3YTKfYHVtd4T2vUxrCIjZw
1CWuBaf9bIlxRRCtLqwPS59/cS0dJcI2GBUaHIj+SScCR+/VUO+EgojZw19faYUk2wVaCjF55sTN
f8MVavOOZitG0tYt8c/sHvOEFtKMjVYWDUne1m7D0I7qf6flhviIm9REFB37VaaBRwIrQZzPOgSh
HTKCcNzaDq15BYJG6Lhf63KTzAvTK6wqqUvp3wVUfu+SqxShwX6mdZUSIJZDQJ2kexAbiwVgbjck
cwuqxAw6RNO+5RpEBrhJNRkYGw4r3U0OPTlWsEu8Hj9iDHJQe0mroKVCTph6JPG2DKPmJihBrzGz
apsJ287tYhSqejRezMCsuaInQxkkRTAoo7sl6wRrWOL48LyjzDfN5BtAn+uJUaNXv7s0sRazSB68
hKLGWTZCUUZAugT6dSsWVA2/lBHU9xaLgaKTnWKbc0YS14GrAvRp7tBD5lDStZb5/oKQKRP3t+dR
ur7U9g08MnDqxKMlWh3Y9y4NgmDHwxG5iAnU44uQjfroFa4lpzoRhq75W5T4KujAMtSV618r2FSa
N/XMBnZpspIuP/A91co+WTALjUUxj2r4bBaaQeYZYSd1bCU9hydC7talQWxeiKupVdi0OojD2IVb
CgSCMG+tJkv9JvEJqpGI4yJlBVJYgkGjLqQ0sTLSI3Wn1oe0NuHA1A2/6EtORVwsFrG4MJW4g/+S
h4AYKta19RLUMS7Ob/TYgwkq2TA67PXarn2mNAWYHa6F5EnxI/D144rvz58duKwmoabpb7ewfsJ+
WYpSyQRlilN8GplTybJdoa7eR1Zsyf9+bZqOeAysFR4vlGtC20Zj4BPBu9qZX05hUqxw4CRLxXTz
XYhSAWcCMjYrLOjYn2DxPBCi1zohdnTsAFbSyBQtPZNj342vSehjppU3G+nyO8+4iiwmyv+KglMF
9/E4PJXNWCPAEQHco2HzoiVRXt4sMdUkypzKPHePG3umySXSracnlWnK4P4WtLrTl1Jv31A7/MdS
uH3xgU84zCloAVzj3P89D+1RXoetEPoVlmDAGn6I7t123kCiO46hK6RNRjxwdM5eKgEbxW2LqznT
jiRA9YvCcQE0gyvXm44chx9pyL+O7bTEoRbuCOz0ZbMFd9w1ZUQteF9q1ErNcHrIjgClqN1VfRF2
z3sy/XTaWqKe5O72+RvoXNemppwlnfMh6uSV9s7+STSLYHW0lEdnOPK0Cn+lpq+/MLTntlXGOV2r
zisFXQxpYRSQHbZda8cyYBs43BtY5nqPss/ouEDXzeaEBK/NAv1XpUJTykB2SAGPUdl39gKA83ZG
/KMh4gqj3xsHTJ8DaodJZTw2M0/ElRVpsxQU0ezZ33BOV9RbStTaEgAw4AWqgIm+3N1RPwX+MlPt
wvXSRFMNcQl/LupSrvZe2Yc/icm4XVkD5tG1wH2HSGzfWeyblyTmKmR4aQ1iZcf6yMatcADF28oo
a785fYkKCwih72zhklL8UTOqVPUkpVrGyxagEWRGkqaPoAgz20Tu2KYOqhhbr/BwTZoZc9KJ7ANZ
7ut/TuiELwMfu9WwLsjxuklN7q1DewQsud+XXYEHKm60c2FeXwHPc5YJ6jxJr87VfXIW2K4kudTx
89CqCerhe8xkEOiPbeuhO5jJEEqZu8QonRy8RdiiyxPF5nFS0AvomBpIWI0LO1uiOslzRjr1/TlN
rVCBBLRsodJcE4qlWmjxAlidrv4rfUGBHdgxqe2ANc42ZaDLTkGWLFaofsVziJfknfs/oek90F84
F5tuL3kkjLtMMoHupVjQxKMsB8zkEE3PTeVNI2GJbuXQhTLKI1aEAf8XkDDOvLw27f/ZtWICWoAr
taqkAvIXqFTgVNYoQgk/c8UcB97kBNHNZ7RVpxzHyK2Hs5EcHzux5tG/cIskqo/MUXA9Cw2AkfTz
X1UYGWKqAyhUhPtqNkIWvH7BtMkybr177D6skf6WDWYfpBKWx0F/VvTmxMoWlvmg/HU2PMCmz7kX
GdC3gbRs0bZL23QR7/1DFhtWJN4p1RxKsVOBQbt9y07dBKDBUE0Tz7NGnOg8unt/nX105WpZKLb/
EMuozkeeeSTClco+Zn1CB4uTC+4yiRatx4a9wEHNCqGyM9lbqurxr9oFm6Ce33IvPDboKxUbKjd1
F88a99XjyQIMD4COJs7ofJl90JGza4C99gitkxEJdyZNIuBUMixaiN/JCJ92QH2avX9BE3TusVtb
zGnjj+qiZQsaHU8fdSMVETj2gcIPlHB2DXZkPgGHZw+X1TAsCCuGsSk3VDTNZ/JpAAkfj19JrZ7x
+4iRoNTEXLklo1DY5NZl7/LZ9vAxhVSIZAv6++hpOB0FWVNh/bNdKV1/hlmSfezHyKe4upsW9WCb
Ew1yG4xacDFttD6LcE3msswRd3ZZcS614Pu+4iqClWQ7CQLWj1+M7xryXx4CxNC8T0jgGkj6YXc2
EezARj3iHjLzaMtSFqc2lOqGLa5p6ntfQGSS6XN0obf/KlxE9qLKrlKQIT2Jq/gQAdNXtEahwZJC
nwdwICe8yAxqhwb8qjVUEW+0YgzxgZkl/NEyGZQH+n9EjE+Lh03ONMO3HfKjuRUdxepHFSwIej7m
ou1UeVKAgCT1c3RfypVCTzjqr9KHDJBCoFflu4chb9+oOY5RtuIwbMDgXcV+SoWMBytFOBdsOKzj
YS2CEru3NshGEC+hN8ctDWDKgk4RPXoxNbZzu53uPU2sH70RHL0/lwIxFZky7HlzlSVntEWv4mhO
+JUdDjmn4kL5OyQfsN3OX5sZdiipgQAYwCaU2APr96dooUD9rdCLMRk01DCrW5BRbYNDTJoq0tsA
QMDVwK37VxkfCFuWcoQOn7eDBFMUp0EE2EIwNxza/M9pYHgFzrIyo4Ktsg1dTZgBRSczAbXZE+Kl
qUYmvKBdQEGjAB2N9JpKm9MyGYJdStIAl7oFQH8DTim4a3bgcnkaGD19cvnF5rgXX1m80VPDNk35
7RPpNp+VUJqafnydlFcjXaoLIb8tQf1cTiITdKcF9oeTU3KS9tzQSA/Zy1glWHEgYEWWR+bCQOeK
KE7blvIA/Ltbf/pdgsD73SMR6b52DsmEl4OwfHw6O4zDdwKAN4W1PixNoaXpJIfbipNea+bXPgXi
TotoV24E1kfOpd453M9SsZBHF1JCS+DjtTAJPPFncKNxLacmG0I1uUMgSxoq/lSElpWja5YBDxYI
GF4k1+yTdC8NoQl/pO8O11KKkqPgdOZQ0DJKOaITy0P5P+PhYSRprKEuv6P04Xs/sqChczYpda1+
MZ+NH05xNr1Gkik5Z82Ja7upGmY0/vOLPhnM4oIiGYqkPpc5b+d4iGjm+u+wfQD/0t7JHI2YzCXP
mv4xEVNMfCdEuu8rbroNoUu8GFAUBKTFFlm9eXm3jhwhrG0Zx+q+avznIFTdPSF6N5aacG2VMPte
/btxIQNbusrxn69+yJ1/59nSCa48zNijYwEIuzqGiZTB+I0uVHNeP18ollQvONKk7LjB9il1S0Ha
zNMgAzTcQq/IjviPJhxKAOwziZlLtwi9BTXRVOIt8QT6Th+sDYuLfJGY1omnmpJlIYIzEOCCUNDz
ww1sGow84iOhxoxuBGk3QgA6vyFCs/8DzZwQ4p9dF0xNIyH8zc7II8HgV5MPkf7mdi5++Yv+PRMa
JrkKZGyZ7H4jq9H5b196lkc6Ts5ABy1AzRGSWQ5/CxW7tgGs0bvULsJeqtMicWVeGIRP9rGTPgWe
nW6GRV6vCc1pewewL6wZBOaYgfv2GGqkbE0SioeIHpuW5xXw2GdUAnZQatlvY3REi7meOjna/xDp
pEk/r3OG3T7Z1UlRG7MEqDBgKDbstVP1uU98COCmQPPxf7noDAwXtIqgJOoa8I4zK8ayGwIIN5iJ
aZa6vy0tDPSz7/W229ogn2KLp0DnjRx/d1jpBBYgrutyU5QWX7uK/KHB8lYb2IX1t9Cg8KnxhaZD
6ITU9ihMkpUuq4zd9BYGDcUJm1zUVqshXs5Jz9Sut5SN2/UxQzwUowp1eUyrI9/1f8eTnhTKgyhK
9FkrkojU6M+kxseLgoMF/kt2FzJ/Ip7BTiDMPipDqfM6bDUJ3sDjkglKBcjZC9Q4MCjHI19fC9sc
BJVKmj/+MUKv88XhNmL4E4noeRwA8Ou+r+0rqwHjV6V762fAmy0hjy/0fKIq6lHakujgxwmcZOhe
uSehAIbXbHUG3VRdR//0fcTmumfw8GcD1CmGBnUAW2+MRK/jDP5UY8mBAi466PZ7w202BOf2nwA1
Ps4FHzrvmDqnI/85QSNu/9HkASHRrbsErBngV5uAELZZ0QYFUUfHNxCyFhs81r93C40d2MMVrpqv
g5fb8p/EZ0DLc1VMsHwfWE5ClptAu2BcImmh+povh4ybHO6gHwZCMUtgpXH1Ap870eM8+OBIRsaN
4nC7aFMinH+tfyCottlZuZwFkVeqU7o++AKAeId/i4VuPTfn81YaPoS7UL32rS1IUchGN3fBLE9X
APB4QFlueCXiQ90O2syKysEZQy9DU1Y8+/1lu24aiPQSJyTURkvOsdfnSYsV82zXyiWmHywt7OVo
MMXb7So771HPrhbdt097PUJpB/fnkjrHNDekwi0WDAiZRP6NZU1PJ4wvHStgCQUXmNwUIgtra523
wZmLU65+ylAhvER4WpPKXqQzifAtIzDYw+huX/zhHs6ExnWe5pKKfFdcLu2Tpd9f4aGt3BkS68Zj
vUSf5X9nfjr78vgX0YVBXU3AQ0FgnFK5gJUNpD20lay3ZpuB1o3yiwMhb9Ivu8skbTIr8qPhnsXn
Gk1pljIY8QVLOFpOkRFYmmzvvQfrwubg9+EISU1sIOsRogzKoCLTIw+3wVHyWMZzNfcszVZkYyrn
iIrFE/THI2fdCbsdOtH3+xazjZnvAscjO8MXGv/EQizdnaKQx8IKXtD6ic1DcKy67yU7UcjDayI1
GPBtg5WG5JyS4ICTAD5RGYLuIjd8UK5N0IfMzGaJb8V4lIfZEzBnSuYlsIFUf2bvW9M/FdYdUMb4
ppiOqVPqaKf1x2lm2LfJA9f5gUDBTreQXmGW/hgEr/O7Sk31auuShm4hDBJqZxWXTxH2PMTlJKZS
NMJ2yDfjOi7HNXGkqtUazO1vj00N8HeCDSpjSu/yPyasHkoVXXRRMlEqt/5UOaRk1mMGFp2tMUVv
0V4S1x25KYpb7k6dVwlHgZr9FqsVi8b1hFuRQnQyAp+w3jqMhPXFYZZt++8sG4SQAPmCK/tgVKZ4
waoq0el0meHuhWWifyjpbNLxwe4fTxVzm3ew9Fe9oCnSOjJwu1a26BA8zGfFbtDnzPgkql3mvenY
wRiO+fpJ82LsLEVjiodhJCVxv9b1zKx704Pfi1bvSQyw78bKj1ymrgw6+dPHxDimx5S6plDgz4F2
ABv2y0V2tWCAAgfpYz+orjtgTvDFbURHi/4CVqYmmQO05XjW7aATidoVGX+AzCIAg5wdYpS4SxBc
QSSkDutpZSj9zZqi2VxF9k1qeuEN/ZAaDW/4L8rgs0HY90RWSyhMQQdY6/fpHr3VRbOU/+CbQ0P1
IRQL8/1wkhttn7h53fBhK62WSGrk8HIWKAF4wqsD/bfCD5n8WhwePZ+NHZ/GK2YUEET8x1kk84/h
TxVElhXCDdoPDnwDq86CQek00f74SS+Ju/dsJfi5MQCDQ6SUGnXS16kweNw5niK6y1QAXeKDYEAA
EGBXIcdCC+BGNuRAKBJT9DdC8Go4OeUwFFzzvShm3uQg30f2rmm80J4a/rqGsqrY9YmJ7AdGXtXj
OrGUn/plX+sl1QVZsAYktCsDR4/lHCt+jam/g3qu47G/Q4cU5sfWDzJV0CRKoJ5UTYlHRBJOAXOP
SRWLp3uLcHofRF1kQTT2LWx6fgZShgVlaDaBodW2VvLgzqwCcZ0qJihEVczb3lSdYS1U96mdATKx
+Fz6/0+OliJrAdQx611Wdj+ALZX7DryimXP3IvNwktlwOLNlCWGOGhihSs/w1R4DBhErfv1x8gSS
pMFj3YKqlH9jR+WiPv9euJSLXTpybEZeoccEKr/40iR2oQv5mCuklG5/x3KeBqkiuPisvSMUU7M7
/oRXz4Ds+ToVv1jCuASTtBrMJV6HaPAbOMKjgC2YcqQVHza6POWiB/q1I5mQFa+DmLzlPa4AYTML
oqS5GwbMsdx4KXdnBJiTptI6hvZ/V5JMmbJdTj0pAC5q+kf+ZPOuDGsJEi14H9E3u4foMVriiR8w
udKLMK/mPmAWdJHk57Ps66On7qk6SNKxOF7+uD1288GERVstxeYDrRIKWlpciPmLvEqc3r0TzDjk
AcN3sA32DNZisf2WY6JaZv78CheQNxCR5vUqye8Jyc79YVOS/y3i4rOCZ4r9i+RqUarAtCg4sbfN
d7MkidFbdbd7aGCHiqlEbY06qpkxOmUQg+c7cEk3IqNiGHIE+DDjaXkOKCCtg0DCvwdAZq03FLO4
VPy1sXFaLxF3DRT+gbxsw9G+mhZBQlgUCZ0TEMrHCNP+0g8Ql7YguynGOOYCVm8LovcTL44Oe0+J
DBWzSePMbzK2tVhr/hdu8UovL6Rl+zX9HuKxG9Zo8zDal5fD8kqtzUrbfyWev3rNnSbGormI9WpG
f69NUs1DLUKgg3X09oIiLM5H98GvBUEU0ID5RMZAo7NhyDAQ+yRUbhc6zw5cbn2+erbQHKNjwD9T
BYxE9ItsElp+EvaK7tJMFrhYCfgqU3gFliEIv+TfJcrl+5A+KE0MvmOr9Y6Zitljb1o7upndrGTZ
dLenRirQjxyfzAZFwF/skRUrw+uk10NZtqKqrVaIEdTbM5fGl7Wr1tldemdonbxV/W491zcbghhp
FPbQIz0iLNKcl4+MHJBVs5h4Ff2qKuHiFWkgEzOoYqCSOt8vKvONhj1LlXQ6IWSlq/Lw69Rr9t6z
Dh2O28cCZC1HtXFpNmHtmpQ3jY4nz+HWGQNoAE1biZh+pHACz0DHVfBfpVZq62u8im7QrQTLKrCO
XMTJmqxvqIm29t7NRZpwft3A68JLqhyO3G7tsGocXXvDxCXx0IjRJq2XnTBvp6fn27mJFL6O4+PH
76EckesGKKlO9POgBTBaN1UEiWhdrO366C47yJG5K2W+aoS51nlZSFtgUnpFMEoCZfldn9qJcVJh
iuf8VbQB5H7xn7ggDGBRDrtODBraWmVc9gRKD9yQhXwM8qqPIu7YsZTzE+WG2Gt1ShjnTs3dOkml
oFOUGaw2JWgmZuffpu3odiq7cuNQyKuHOZ44ZDKoVXAPR6HtFIRleodMW/nVChkrqmRr3U6xh67i
VCqR7k2OdJJ87BlYih+zyyILYwc+nFZISX7LfGU10qgDMSSQ8g/X4KkF9bbn0HWcBZSZmeOK1Z4U
ziS0oL9uH0AgsC5/m2M1ZTLzKYGELG0W4t3NiONqp3utTfxGiVy4ucWKzxYuiHB6AlOtJ4lDhB14
elw59dYt2obLhPycR2G0K/RJzVsd41y0Z4fNJ7JDOOVYx56ukCe9jp1pvK8FFNYZLtIcU6YS+QJ0
/IvmSrmaGqZLoe0EVaEmDidpp+FPF9YiZjTNyH/XBu27UuJlXvYa9eQ2EAUI68V9uiBHprim+4pn
nQNOOAprSSTd3wVmguWN5mTb09uiHwsSo/t7uOTWVNj1BAsKJ4006zM8majofyqIzwL1zO8u+NpX
SEwojMnuX6ro6BhCjt+nlvnbxAlNb05wv+4oIjw7hlKxmopnuOSfVwZOlY4gTFvJeivgtatJZR/x
UAPsVRIg7RvXEMyYMQIXTcfhUTRSnhUD0Mvyl374261UxwvV4iRcoyaUwkf0LolIU+luYlJx0B9n
t0A1tIJDmGv4f/xhX1UGgYHBPLwV66wlfkB6Thfw5Do/Taz1/6wAe79JqG8wdY+yjbP/VnZPG9BS
iQm6u+itKGVJi1blbojp+wUyo4tTaVzvR731CdRWvDsI3jkhz5AX+IgZibI1PhSarYhWrUhQGFjS
LFyuKcDkEv1qSjPvaKqHXpmY6iyaWtPkH6DTg5TxWxl6FZuXpDCAorndjFvo5tIByYDKSQjH5e7D
TOQyYbf+DD+qWTw64AJntAu6pGhhKYuyL6+QpRVN+EuVV3zcXhbXy9oXzYrLpUWFUlnpG1Dek4oU
nKqMg7Ca14femtQEJGq/uEtFpZcA3t7ezde8yUhI/35m+JJCMMNEKuPA2xDkwYJJr64yLrNgJuKm
3J5MjfMkVKAu2AdNR0zJfXhiQrTt/9jdnQqjT32de6M0Shgc51SdIS+BZGPpjMHVEG9AhXyHWKYz
B9ienBrerQtrPvEHSdu1h6UaIZRjojigvLSTWrF1Ok3Q//IgAU/3uHws3WdOw6+JDFDkJpIeV3yG
60ENnC4KpQ0NYUtPCNjEfrbZQw3YthshJN40wIX48ZRuun7h36DH2B2Nbn8ZERskKU7ylTjZEGen
j7y/BmOjv+/jWQwTEqanQYR+qGAZZ3+4brhXiTvj/AtigWrztNpVr7dulFQXT4fnjK42rUdGSS/Y
EL/75odVRON2ZJAmgnFvgLAXeRkEXdBdyXk2bBLxIIS7Z0grDOSt3NiHcWpDpUwnWkazOx57rrY1
FRuwNEdY7tedtVBiffSqwq4pTw/6iFaWAFUrp1A3UF51w3gLjYTDdQBdKcPaxsIsnuHaws1gawbZ
aei2yx8RCHiZLGQQdZ8ec2ckOjViP73WnW6W8WaNa4hoFs6XDT0K1dW5V4Qxvj/yt4qwX4MVO3U4
V9a6eQGFKK5iTb3ljNPa+YJNrtXpJqQifhA0lsH8ecuslUBwh0GOx9zKjQMr/WxNzOFA5eiid3P9
PcSIuQGa+DyBlQ2UyJ+ZDioxkfpGa3zy8Yer+EHc5SOIdH4xPYjnmNGZuN8XpyPUzF7uLN9oWxsg
keoiOhbbyz0gW25xdZrQSCvTVCoRTNcOefrj51rtkfSZYP1Q84l5aawYpmKosG8oMvnJlmYNiE+5
caFVafBwSKWCuAqiQVU3q5D/d8N6Z0SH6TC78amJ965Tz8MFeAmb9OsZZRQeyGgYhUVhLlygs+05
uvcadUwfbWJf2fNT2BWFjmTuODQRct040JiOW4QeAGEzEduNsHAXczOQ6dKTp9rgVkc04wQaD/C7
IwK+WwvFuESThDNmhMO8KmqPMCwBSsyC2uBNFtnxYXGY1Yf8tcVkVbd2Aa++gfTn+83wtuamzkdM
m2elwqAFqstQllDeWizOWMhyUVZg+AXdO1hfKQdHhcuJ0cFjUOGimiyBJk8nqlDS8YfGbgRoqDBA
S0gcGH7qhZxxT3k+YyhMSzwGlpd88HcZhlAEHHcSUpkwtKTRZSWLsbPMi+dI6tKSnHURcpdE/Zct
4b13zqYmAblio9coOtl7A2SUEj6//DUZZqORCO6TMgvS9yYxymOl0OBQYHROAg1Kj8cjH6+iRF8c
Y2xWoweCLpVWbYmM06hmvLj19+XH0oM38bt/Y4rpzNy/ugLUuky+L6YYPjpJdquy5sLBPpyF3MKi
sqrxDAkjzAXnswdRgSneH0/fFq+oemqSeC5fAHCtw9h72Q9AwV/wegT25GKRAqspK+hdKkOVmLCo
XET7DHCBKpwlK3uKyULXhKw65DPFR/cOJhYPwI/i9BSC5q3t9PoL6Wyt8AApZTTFMM9xHGD52Qp2
wyM8p1A7/3L38F9ZiTQ0l684U3+y+cVZuGdujyuZ909eI2YrsBWdv2wNYHG4feyw4uqEtDfzpXLr
pb9WO7Tsbyg7Rw0a7ODnXKGuAhNV1dndSrzvQAg89kQwhrV1e1TbQrBXRtlGDp9PIMwCprrr5MwT
IqMeoZvCf3CIyusCI47wurM6kbN6wA1PnmBmFFzlDSqxPo+YQ6pWFjzqrVyjTbRkgZ3JC5LhYRbz
MiorKknmiAoBwT2YKDG9h1LL7nikqVxOXAKuCRR6ytBkGdyzTXFsHqranXed0rROCG3bd6OChbaQ
ND3wEw7q7CBXRz5uelUDi2T+1lXBYHl/MAhaD/oqFI5Tq4NxVoxcJUCOqWD4eLfN7nvx/4Dv+Q5/
jU9sQ0KaWpAAaJHwff+dNY4aXteAfeazyCglUvZKuz6COpGDL9v7CkC7ZKRaqtD/0ogmVApnd8Mw
JWwrLEwnR1Go1ZSp1elCfVZ0mlE6bYiU+h9+RPptVSs4LvdKbOgX3yL8YaJK7/onFEuRb2COjjpT
f9Tc++pO/PeEkPos7FTjxxYGKawtfjhAjFOOdw5iPaX9yuH/8XuNOshKM8fDY25b09MvOBVONVX6
0IqIT6qnufF/h8rWGK+6aOaot50P1qbjNuNqRSN63J7WHyhb/VUC4qRB145By0xuVn+QMHsK16lr
Fy69+mIEj7orURBZc24CXCPbr/TCkH3uv7dSk69jtE793i93ljut9bZ7fNwhh1PGZZPeMpnUM53e
It4VJsmo0zCovVtWaQj60fsrxyCesrPXsHPGOFr8CEJFB211pWFPOxxHuKQr2xMVj/Q5VPjN90jf
aeuS+jZQPG9aiwZdGwpPg2vNkIwcmBVEM3VtXtKaMm0rinjQ9TJwL55GFrJxPWBz4rXAoK87bAvT
VWhq8hcCIiY3F+YWCw7xZwVhcHw8/xQ34NHu28SzAhiMK1N9uMkA9ALTJ1Chkge/IjovSU087+RC
uN0k8G7Bgmm3DijKvE0oYUIANHIuCzmXhHNg1nHKh9L2pCiS2yM55tN85FtHJycvDPSn8ro3hhk6
/pQoAILxBgtnW/dMoMhkSKdemZeECiLRkIjQFtf5L8ZMefj5moS3aR2u3VaV26OJyFosLH7G/VRq
yPtc/1VAxVk7UuRY5O7211CpkZyw4zyttNuDPzc78UaxyccQEynoyrzDMA9KusevEXUr9bOzn7lB
akQXQSbC4/JnrtzK6Jtsl1lifu/AnLgSDGMtfnGvA1qzWhQB14+U2QMZkZVkXj0aHvQ7ue9h3hMQ
LZVCy6ws5+eTojUf33c8/iYOLHR8ssq1cmihHyi0W0UAhyHzQ6LubfBFfvX9dBC3Hb40Q2uD5lsV
v+ynp9G3ardosyCQ6MMXPHKXySfpHHpChjoEp5s+GX1IfYNKLitaCxLZ7jEiB6oCsZ4AbPxLbzE4
7VksH/hEVrQIBSSILfcfAMHxmW3wntJMM6xp1GJO1ATNJWUVMa66SpV3FB+HOQ+pBQQwpkvfVShB
HCMBEJsHbAiDqRra16qrC13czN1SWQfKMLJTC2NiRbw0zI6s7dQvNqxR+K6q0eYrnvmr8D8SCBoO
bfMrVSiGcddACFnTw0uDIchMFWbHMScxcoKOK5/hRsOKWBV/kxKdNJVVFYUpjD1H4+UtE2Q2GJJc
EPOo9QKYBHHoyRgmsQEdm/VpkT+TLXN9gOnOsusps3W0Zx4/8N9VwLMaktFAKRiJ//pc1F8Mpinl
x52e09l6+FhHze9uieK3sFG5lmjStbDztTosYxa/Kj4CGmNefXmJeAZDCqX9tmO0M1yiOFhUuRN+
1gf822abiSpbOhyZ3NWFl47Px2VtGeYBRsavKy1qwB+C9d8wkW4G6BfadhlXhNw31PtWQGbDEua0
6idiMjUFLb52GkqdP1p4p/NDuo0X/HgfYg0hKL8M3L3IHtetzuflBDWYTpHdS+BxSaSjmbBGmpM0
FtfttCMRIG3liz1kO6UGZNwrtyCQMkX8O1B/zB1JtccueoABlwVfwIXpo1/NV5yurnEW2BXtBSem
s375SuYigzixyPSZi592gBVWy6FerDP6nzIdGZYmda1us3qAgHzXqUZg20fzPPEo/Th2h/e94lAg
nqpYdBPIgKX6kBvn2qHXk4x0a8JCwmD8/5y4a1ljas6q99YA7jMAcn8AzwCXGudKmjgi0G6LAZ2/
/s+eq8TcnauRLd/2+yFgCb2MpkMeHZOp43/CKtk2Nf72DaK33nYM79SEba28NwipGx+yf1WsG+U5
fCgArTIEmKTDnn/nYJG7T7pO5CD6rZvsFYzHIOUUspTLbfNE2HTPPsKw30JCyCrZE7x4Lyn/Dzbx
E4Yt6qlvSITur8nkHrZTfCDud5HsPoaHFNROkHyxS0LXzCEIRw93P7+Zfh/u4F1A32A7LEQLE+ZO
VjpFR3aYYaFC8Ntb4TaH95opiJoyfyDk2lTJntSeMsTEgkK5FxCrWSQ3dpwTzWDvRPfyZbWW6Pfr
55Y2eJSwTYpqprpVYzRQaHfTQJ4yQI/2pmV3IdMtg/SNGxBt5itNHqEKPbXlsaup6Y3hKsL+4ZJv
mirdla9VdDIaQWy/Z83+L29ItJwsx1J5t+fnJRyKzreaGsp/VlxIXEZP8BSb8bz/rALeTEebtHZW
BjAqU1LW+VlE917CuGbwVfmRhIwiFMpoIZpK0Ka+ocMU8nkD4jYyR1FpqDUaTCQjyj6yrhK4ag0q
XU+TVQVuej2ay//CijZse/+eY09tcu5L4ix5WkS7glJh4+T1o1tt19F9WJ21N066HCA493CTzeGe
YF7bMvSyUWcnDZoVN1270+bNkVO/Rw5Gh5ArrNZv3MBcKES7TuDquWd8w2Vh8zlKzNtN2rA6cf8K
Xw1EH/jOB5bAIccl5u7vcMI+sEfcnewwlA3QCOU9rN7gSD5u+2Fuabqqo+xtvfEZe6+52ouE5Kw0
+ntS5GiLtUCvAB4FvQvXeEDLuTU/CTgBo0hkTrwc2te99pL57u8Oqe5RV4OMfFzUK+5NEIVc7S3o
BNfpHv4vvLN7VaNywH2WbfJ5jHYtGex1epMqEet5QWaAlqiVIznz1kgZ/v78cXbDvI7SRyXmPCvw
sSx3d2jvaTcWfwpA6EPM/G7ONf3z3725lzd+LrKDi54y6N0dgmgP6A8EEf6GgKo78nRfAHdlVGrv
8pkRMooy3rYfUjC84q8Vxdgwne7SNWpaAedEosm+IumqWCI88/yCR5pqxsmtHTF/YXfGckvd0BUM
dokVgyUVxaWdUV2CRJYvLesVMgYDI9zSFzKq++n3cFCZhCtgzk8PP2lRfgR+XlfVe9fiKiL7uZhP
YNL3jOxIlxEFedimwVF5JMZYkYiU5RCrhs2fEbvmFhH6mKJ78j96AARv4SVzdykDctr9YtHSXVrh
PYUdqbINHPoFfpD3m28ApYavEJx3971n8MS6k8EbEmp5rFlmrSUmJdI4Ntoo14+ZNxExJFC5QADU
WOnm8/7RRLPbvuoGVW9ZdmZinZNqx2HXRKJTsg3DQgA/Hub88KOq2TI/hyqXMvNEAjIEfGtRClHF
teNW+bI0uo046XbFVyvlGdibNhSHaMW8LHGu/C4nEX4yDUHiHExvoBs5dRsiLYRf8XTRIXOf8bCC
oJInq8w5wnlVDl2NpPcG+5TH9sspcTZrFDwijjh/xyAXu0DsfvYT72XETaxvtK45gmXHZ/ob7oBJ
woWnJX1Nd4zxIXgXN45MylgAv6phNYEs0H1L1FxIgU7coISQDHP0RjFq2nYxts3TljJLTocwwChL
EiWGwFkpPETcnMibPJ69WoOZjRk4GBGjjdXkkHiZhn1eTZtKb4ON5sisjtHw4Plp28POrkI8hJ7b
q9C3YPBqCqsiCHh0fEGWlb2KAiJLsDSWu/qytXa3ufLFeWP8OGhJFW4Dzt2E7O7OAe3NlGrENTiV
sECFV+Vkg15jFY7yO7hr0lyBbJWSwZd4zqg3n1aZ7HHoA/tIeaI/asTDGR9JzC9jA252i6T0V2P8
NhS0lV4Fthm6TSixSE7nzs/dKpIIcHohRAy76AoZ4RiXIeaL0eM1+x6YLytxjkAjrDlNSv47BYoo
xB1CD7hxM+CYWTdtu5HDK+Ii5yyMjt5u+J//IuYtkizCvjAAhi9vOsPCRs4aKRrmesQpDpOdgT0d
4FUCBWdOBjlx7Gs37f7NHxhfZHq+HPhtv0JSEccCqRk8b9LoNvmL+mTAYCaWYFVkz31O1L88dn5T
HzcCVUaNnbLh5BP0+P1jZ0qwEDOEl8XRsngYVYP3PGixXDpvyxOovFPW3lee9uGW2EljhFkvue4H
Am+TAj6BIQHNp7OZFjHWN4i3yp+nB35rYLxSUB3sTaeMC0/giZ7UFtcvNXlJcLvXM+K3dpEYzhor
d9F2Sg9Run8W+Hk2BFk27MOl7dSKYdFxuDx4q8G5aP4joGx0uOuD4s9EpO9iC7YNQf1EptYUkBPb
WCkgLb26ZTqcpt0c7omgrTSuNtxWNwjxveiTVYOIEK9cWK2ECQXeMl+36pA/hYIRpibpRIR2PsPg
EOGNN9ugTj/X0Gho766WpWiTdQnyVEOPDRYCjTabE+MM+ZZxWNSYdrhmdVExQ5HtM5NMQftdZ/PN
ZswuoN30a6vyFzwYlqut9FhiWDqARVlKx1tm1Cr5oMFPvHDyeMUKrD2qCaE5IulRA4FrPD6vTCYc
bbOr3c5FD3CAqKoQgc1ydiqIqvwzqlDxwstmhx8Pf/jFBNJV0lFcTltDF0lH6pqBqAkkjZo/5wLI
5sn6hXp5YTwrupGplTttUXMlyndTtOvWfnIsknnFrJFHbvaCiFPWR9rolhFDp+SUOQxx2P7V5wP6
W6NQpBPDW7FGXYPgQhbqkQF1HZC7HJmJksQOuOmfito+0YE8ATe26hWYHuSd+KEztqszpIBKGBB8
1oZI28xsfGzBvpCm4a++8JytGXIx3ps20KFsvyvLSTfG3HXZiYlGwn7vJy6FYhlruXmCPKNIZOsW
6xlRnvHIgYwPgCk3ZzQSJm4lTwrW0smBI40TXmcm5cD81Ik9h/eBrGG5yS3fi1NLxcpakucxl9Nh
t1SAuX5tQpRr3O5iGjHDOV9p3TNxYp2D2bXY1JDbaADlcsrLZ2rp146HL8TobqqKCUeAU7oW6SBX
uj0QFNrZ5MzRVosv9tkuAA1yLmZSZ8gsMhn90ppqESoQSA47tBtGFnWKnwpQeo89xsBYnV0O9bSl
kIGf112SEQoeeoJUuAZ0LJXgf1yG2p6p9cgIaCKS9UOwZl9Bpi7bg8rWVlh6gRnLIoIuP+pjJT3M
K/Z0Hts0jHsI6E8PPuZ65TjYNF58x3Vrywe3x6VCpvEGUUpSlub26oAdr4owKeoBuo8mrfBa0lmm
tR/CpZPd71k1aZHBRGzJlSqsXbi6OyCMhg9Rbq7tJ+PFT5ora+dd/1UChg2G1Xurx/vukxgO32KL
2izuqUreT1DeDeT68Jw9QYj24khoP+jl7sP95r0Qb8+WPG68ZS2qOpO0f3hEzeentYr9+mVBiMRJ
Ck0l/2EgaQDMD2IA7A82YWNoRl62Q2Nm8LtCPLShhdy95KT/ePYa3vrVADOtbHVdYEMVV0RvPC/U
htwoCddvkbYDYdVFBY4lZ39QyvdhBBX5Ez1uxfkkOncvz0+dEFfJO3+yEwm3AHMKfJBI8vUAzazl
YGnLSNbKQPoZNJf30Cfc2YxhaL+2elhXnsIcZDG9tQCNKpVoaHUnEZMlrwhEtXjKBNzZ6B6U1Wa9
AHY9Xx7S9neJqKNa3ExOfTeG+9KM9b6HiYMJM2fkRRO+rGGoviuHYSyUfD7jrpXum6ahAlr64Rb9
+oOSYsx98pur7E2qCYUVPqnA0ocxsqhENp4MPTlqLH/mMO8MJ5BVzQyU1u06eR+wmCtGiMs9vgIP
F6vIUItaKR7fJnIBYYfYpQ0MjDIRJG83+Vp3U3+uB2toGJxI80gw8fdygfSIXTyd5wUEzJHB3hBj
Fd1MXvZVD/DxTNhEngr0l968cOVIof4ufizesLvpCjWC0rkNXDc+aNtdHpSqG2BGrHXe8ObzFk7F
RX6pUX5sABd0QweOt0pGAYfY15QEiGW2T+jvXhrna/t5CI+j/89JilEQSiKQi5M/nkBmf7e7nyBo
+kHnnnbPOlDv+bloMMOw8X7oPWfx1tRX2ol8x1jJz6t8cg9kF7Vq0jBC4Rv7ArfojnklNEz3PJte
Vecsb468CztUMJKvGgFVtwpcTObAZBtLBzsPB+cDjeVEHUdumidS9cdo4KoZnXSIqd1qIbpq4ez4
4kBhuUV8MvBsyBrF6ZC/um31W9qhXxFZNa6MbjTSRjo/9clpSUk0ytVHVGIX1eaqUPQYMStblpOm
+Un8DuWCWPaGHtjtd4oKTU7syZ7B2dnijebo7MBfFL72WWM0Uy++F3ZiPM/yaqMh4PG+gbz6Tetc
Kf52rUt0skKnLIqDv+5znH3QjKltCfo+8w0PHF3eDQRn/Gpsgry5WXIbYntZcr+F63mctPx1l80Y
GW8m+I68oRgcfDi+wB1PweMKZ+HvIXhfs2rrJhYrp6AKXGSk/58i9rg/ZO4oqzZUrheRNLLfSNW2
MVRx9UNEMT4R9Wip0yWSRTUbjlvN6wdLGexWqgqIlXhJAt+gz9CEKBOwt6JV0YwP+GMrt+VdTnnr
hljv6rQg0L2hlxSpkXL4D2jwC2aLcRetTSIUBrn/6L8qi058out7LX7cb67XvRMF4BY388CnhK0z
rdp40tF8U5fzClbu3/LQJiF2uaMxpdTeBe4iDkHbrCebcEluhzg4R5pcjxfEA4CtSAGEhnxm4XYJ
lSiqttJKvsdZdtUFkXxJS2O8ZS0C7B2r4iPhf5Xlt793PdcTXecujS0gQ+z6ey1G8dWBR02YM+Tc
orbx03TrveCYmWsFiunRH6aTs+6xTT0EUw+1DO16ljSsh3hJb8sPY7Ye2B5KWFSWCWuVVamqmkAI
kPJJle/yyL9RROXxzvr3mfCQLhwMhY1QOcNNCsp/iRv7vm06H6OohrOtC+nhSSNQG9eo+C55k7fu
SPndRvyEDE/xwcYPYQ57yV8v+idaxys9GjrNeuLOTiel9VtOG2D8WU4bBpEIu+8NVm6mGLJzVc42
IG3OU/5XnWqa2/DNHcwmtywkYjrazWZWzWvaflcd4Eb0NRB4wubbaajkRcM3LKOMZz+Rr2Y1UNyj
qeVh4+pV9SeJswiNknS0qy6M4LVBv6I/ryerwD4c5xtsLlSIpLSRuzzexc76diecRflIk72Kc976
Mi2eu6Jmr8UE0H7dc7gmcnKCwE2qmVjS8XaKrgeJArYxo0JHSo/AUc88M7Pz2hQD/NaWpWZl0VyF
eO8u8lqt5weVp33oo3uxHMG7WOmjy2oLizHo3/pbNh5PcMT745zDz9rNI7HY39pIFC3f3npYwUPq
r8UnzV1b+r8Ezyh0EpPfHl3anpFj5wfXc4bjnGrMJ66dctzoyS721Ra5gTqWMjXa5mPY9KiIg3cU
fNdeMzodcSB+9AFvQEXXSTrda8fTCp21s5wkKNDYGQQMUDspRFMclfQNhMMSnAHSgo6An9COSRqy
wAsabav36mLaq8NI5koW9COlRPZU15olsTklvUUWIPPlwab3USX2dYURV2scbs25tzWDdmQMsDtT
nnwFYb93/q9E7DJB6xffknASXrDNaw5AF3/+AWSDBq/KTdwkD56xGGJsKCOeumO7anhhgzPrv7y0
HMjIWc17up0+AuQu2FjYQrO+Tp1PwxqoOC7rP4GrrREjkJZNrs96aMxojWx0ilyLJUYW+KeeR0dR
PL7FjPVAGsiaUSGKZV096WHJ4mJYy7WjWiIDNWaW/b4GKF7T+Hofnb9HymNqgb5W1GezOFP/x5RA
VhPGdz0SYRaP4FENENCr3mMNuQZtjMXJHW9pTNj3p0vkosWaFdX4ecyzW+52gXNRTH1lnKFaax+8
HWKDfnMammPy336T08RlgS7A0JpsQg2DyMmya7q4TMxq/9tyY82vLY5KOF6bVoX8Fy+yio8hWGDh
z/fb9c0eRI6sgqTWWd5E8Ib0Ncjvs0Jr09aA2I/n8c+547fOCDx5GwAnwkgwRcwZRza9JcVbXemL
g+m6ZwgJUfh9Ne0YHXKWctUPyFcR5upRgVthrDTPXVmsrQU3IXNPnPMI/YnhwP/qmEyCHLcIqgZ0
3lzKKl5bs4aFpO3N/oIA4XxANLnglcTmkJYg0wJ9EAM2REPNsEcAR4H1Iusyb16HKrAFZAR2eID5
/0OYsprhO9I0wRO+byzf9Gc0E2ldiiwUisUxTUwTGcmgZZ9dDfUl+UkL955z62NlrwO+aMw7UiBG
brAUYZJOXccyMTVZnSNQs1ihAUGZQGeqfOChWTgZbHh9eK97AZ4kJbzcK5kSSA1+/KdWiFoLMdnk
hEx2cA26/8zJ1S7rKOyJrUtuPlVsk+BChiAKThzdpK9RK0bV7gGSLLUwQblH3HSQMdAD5MvFyhLQ
GjKKr8ZmGp5P/cKQ1EkLUHHtMhT0gWanzRHetpiUVoI+WTA1Eq8+KTNUZ1Ma5mq/X81DnsmRLAgZ
tLL0LYt3nO4y63pwwDQl7GFgkJ5Ri2JBuOEYR/2YM6vPQAPzQ9Sm15xkmrxi7A43FsZMMc34OVgh
ym6sI8zbH4Z2cU0v4QohUGGJjOzafIemvKDrSPIqbKgAx8jfOx8owq4EqsoO4rnq46vW4+9N8uvO
ZirELhvM8W2vaxTQFotGXrnqd5ROb9NDg13cnDs0icqVcoXJbBBMZLACWM82Ndf1Lbd/U3o7Gfsz
iYatNsIA7jdJLoayQY/pIGKmtEcf8ITSYv3iJ4AW3PwahoY9A/RovRAO/jCR5+S0i4ZQbEcAtmbK
iIlxCa7VjNsvtl+vOmWNr+5nfHhIXoHyJN4WDtPqRzId8dtNQTv6zlRi44xq9DCRxrMyhHd4Almm
3acsxlonk4ulNMe3JQ4qPIoXsGWaHuzBG1asyDPPAkL976nIldYm45v5x8T96r9U8PJGsDqUK0rE
zd+TQz4gTx3U6lsCgtJdm8m7XxQrrp3s/paryJ8XiOavOWoh4p3KofYfOIRUFzgiDeaknTvJRlVO
0hwEInJKtVdw89uc1SdyFcRhpmKV7GYLp2Ib4a6GjNm+y1JNHdiJS6kq5vGJnlNac3Ny0yV2xK+6
VTKHN+rfbwHPiJEJziksPGDzfYb/0XQ70msBgbhpfUahytWbSxvkJjueJx5AiSgR5/GmCEMycJad
A8R1hn0UN6eyzIdN0+PIjPF4SCDWaeIeWBjUUwEgRBqyl7k8bbYUB/yvZProADN6SpesfXMb39xH
5qpnHX1JYzFW3Hjo/JgWCFeUzhLAG89ISweRYBzzV96BtT3rSHtDHkDZ/5C8gCMI6pLAeQ4L6iU5
cPoWRvj++Z46HfU5KcIVFtFrMJZpjmMhA6m69AL+FHU3mBBvTmZXGQ0nSLJnXj7ry0xd2x8vJCTf
y3KCfJ3wPhLUw5Rtwbw4RnyLc7roNRte3QziFq/HCxLyQQc/dUC/vrA/kL1Dp9ZQUBDdxbRatiJk
jK1AECcMssOvyS7l+t6MMbTQznADtiHDistAQ1xr9YONzW/sj09onv0YEcTEF4ANcq/+81OYlrAl
7YUqs3GV4oB81173+QztLrEp0ZmKBx0YpkxwX1z1xvxPS3YHNpNb6OsOnKpog5eYOYyfUTAfv9Ns
oaQXPwyjlw6SBdGpzzgWgRlYyUV+MMPymIkpX++pGEGy6G/aCxLCSCldNHm9JIrm6DVTBnHwvRwV
i9hWQWYNLWG3LEDTHJXZ9PVROsV0V+RcrDneZK33tklxTgWRRfDFzb877+LyP5Y25Aoc6Bf86ghX
9RCRHF0T0gb80BjG5WsKNIXH+TZttItfSRPH2ij/iBEJOv27GaF5+T7kb9oUOvDxvbFTsK2og+Fx
eVwTpAL08njf+mgQeXPaKMIFZI6I/lYyJA4OhuO61bnL90E6RMYu3RZiBblAaV2GoSGpaJ1AUtM8
9BK2FVzEgORbpLPgU4O/z4UZWCmdCUxZ3d2R0hd71a8Bv7HWdWQVueOlFMm1PzPeUH7KdLKAEDw7
qG9V06weT00BNTQhNM9btDI8XIJeYe/bWSUXxvxFOJVz3WHKsB0t1J92dUMMs5M7/fRkdJUfOuPd
4o75me4DWSg8I/MP6GUaph1YXhEb0ZkrDhT/XjaOFgLsGBQpZjtVduiTRlKVmRErEwRwVVh6/yAt
YmgDnfzvfz1DC4m7qUy0C8FnWUTCxV+y4xWx8JOj7nOdH3aRsHw6QN2SFpuG+6qnJ0AMJtEJfHSB
IWOb4/MhLQ5beoiwELeBdjEbIU4Tan7IYMvzZAksDlHYYU/ymaJqbPBGVjwfHi2XGc/3WhYvxq9u
A6/i3EI7XA/ZHX7zHOVXcOuziIbCZzKjAcGk/yCTl8Zshv8ayz3uKN7MS2PO5lJYXd7wYNbuGmEI
ucTfdXS9OcHQeJRXwmlph0rklsAd/hyyHxKFGAN/walLDFnOSsa8eDFS+6yVuOGvEhHRbMEbKr43
fWPW/v3mIHCaham/UgJcRQob6LmsI6YZcdHKQ3Wv5dqRr1unzgCHhZLrJjCKakMox1qWXFdGqQYI
9c712/8aVxfXlSkrPlQgb/57YrFnxz5sjkuFFuTjl5o5WtzaZE9hoNjjFBJFwfMNAwMsPUpra+Ny
xtiERyiOXvkLiA38iw0ZgML3+9c+TPdgkm+mbX0GPgX8axKcZIAssWIqi7CIUBabZMdS6CJF/e1S
pr4Bf5GfGaImLQ4lPzZbcObZeq1MAZ+R6ica1EZyH2XhWSouY4acf6tMU2Ca2W4a8Y0JwYXaVwyy
i9aZ+A6+BmZFj9x9/AWkNGuE7Wfh3xz3B4IKTGm0UgLtF6h6GzDaADjBYc5KCK62NXrN3bOyPGhd
mBkJ1p0wUDQOslQ4WHwS2S2caWHxYyHOUsD1Ga+9kRrB6W7yH5r5ba1iYvgJUIRuORS6LSkphLRa
zkFJOFvf587HaQPhzTXME2Vuba8JJhp4uls8UzyF3ZoNXakqMk3nvQ0Ozj98t9B/Ml8+bgXDeNwA
xEqlHX2Kjbguux7GDH3MVkCWMYhfokw+rqmyuWGnnprWpsHbGaYNIRduyCYX4E9UqERBKvb1lX4z
Z0UAiPcCd88U6p6bG9PTB1t86x68JU9s8BgMJDGLd8lZ7a5TyeUDcY9K2DsSjeeDG+3BMTnysdDi
AZmaUXGTAGhq/5cE0PF06ltLFbng+sImzPfnHB06KvvJjttAv8F8WGDrIGXT/C742ze1Fh7ZTmfa
6d9eQ8ROvQ/jgwqq3bNB7znNwuBVAH8rHxOruaeFRcSDx3/shYnO8KECF3EYe3A/iKYjtYmx0zWb
mZKywOZ9gqaT5x97HCEOZtiiAtgAIDJJg93xr1VL8r84Yjj/T3o8RcuXrdhImDF/s1TkhNHXj0el
dGN3a/p3s0B8t5oZEhEZCEGST0Kmuhox8/CJAbqod1Lx1xWqddkb2CM/HxEmdmMggwSCqReQRCOb
nmu5TQRrqtGChmlOhTel8gnQN62Ub87nJxif4V0BtJ8K99cue54FvLBAeppVt9R3mVt4TTRYncqU
fUoHQO+ZKA+snvn9dAPdz1fnAFcpgPkLHO7bwHXwPskRvaEv2WuktqhAF8g5K4MzjfV6IWKjmI31
xJ+kklPHbRNdkUGOdfnjk/Ge2ZaH66HbcQd4KXxDGI4pRRjKpcHGRzcNsFH2STDeZ88PPoTUY4sK
fzvTf5RypZnovynTLnlcpD2eQ0uVSzoOuIbhthiY4tRxAfjadiYk/Nei9bK8ILSrXZT2TB0I8ix2
dqde4ZR6EAV6+AWh6Va/DvcM2nYJmPwc3mnHJ5rVDl1wvb/VUt40u6xK0XOC8glxSGd3xp7Rh0DD
Le99xeBgN5/04RHImG1NK4acOki+6g9L/JuNabZqTTi2oBZHo9dEg047vGkN5+7tVoqkQ992rF9p
tTUyF0X7Gm3hFpCaNHGaJFj5a07g36asLp4vzlVuB0b3qNeQgIrurzHQfdtGSQdjqur/pjrxwfca
IChlLWMibYDW9cYXmuTdsdzvRPr4Bmp6QLGuisG+ww+wjDjJPja+dIQwto531/01QMEIMR5vdvFw
76ht9CX6fWCsNDcdP1TNkDOHsmDIrJEgSrLiZJy+/9/kM7np83yzp3bs+RQr1WqrIWeG5VP2kyMI
j0LuYT6tltjdRTpn07o82lmA9pXDRn9ndQfadNLCF70RtUZdWmwFZbbR4nN950ImttYefi9lp1QM
cpkQlbRzYnlr45H27yZIxCd1LHHlrmZJtl1uFvRXJ/Uwrn6qcSpTXHBLD9Du7mheUX8OpcDAUPML
Dc7JUjAejiOa5rNAzd267uzghSjIdz3dmPea/wn4tw1RfWrm+meQsQ6bA3I/96jSvaoupEMc4ESX
7+ewJb0Yj/s7OlJGZBLgdmz4OK4FHfBws2k34EZ4IQHIpQx8/Hq33+AaQd6ztxkD7iNie8vuhKZr
d4ZSgiCFRW3OdLgWO0jaoO/LNF0bEZt/V89aHGDwXDbJj45ou/Eb/6sQxPKCMP8YagQi3dGQ2/Mx
HVTf45yGZtEBynlROt0erPZqJzem06KFJjqyFUex0LFm3D4kaC6ZSRknaOSa/7dC0J1XOO+m5VJD
vfz5UDJ5I3nRQR5b0d0Hkq5yEPiwl1Y3aYS0k7MngzRcltXAc8R+xB4kWZYw6KJ0Qok184iSjLTn
46tNdonsrBM0/oDZozLfoy5HRr4VvBJcKkUPBPwBPCT7x3mPdsWzviXyMm03X9ga5aCQnBFj/hc9
EAEB0tIEN3giCO3Qx/rPqmKvauzPek+Aznel9TqKAekvSOcnxCYJqXlFHpsdnl4OWD6KtHdgiRKF
Jyj5vtKe+CaAjOoy+/AuvXECPWOsEa8S8AwWFVDT+vO21vCc3iWTO+v0jEiLPE0sZCI3gWDbt6TR
a8bbKXoNtFHWK2Ehjenmw5MR+GHE2mUwy7Nl7qGh09rJZ0C+HDtgQqyFTD0UY1cfiDAP1cGa9Iqw
3eDz1DOjZt5sWDKtDW7bUYVHb9g6t0cqH4roFBC31M1sGv1wCB4HBinFqWdku7B6uUYPWLR7OBWD
xahY12AaMjbeAs75w+hkmynrPZORTjy6DMQMHyU2WqLi1g22WYFMFKYn6zqWIY3ENZZ4tzYF+I0U
Nzvt87qEFy/Kxmeymksa9cyTGuDMzb5yzQ04nJJ6zJxppBDKvmV6vCFDDTiegx8dJGyO4xOfoL/b
XuXqn8C/sSm7m5qgmCVMwAFMZfJbACpablfmhpbqA2DKqtu+SyLJAOP/MjNyaXjzw6AiF/e097Oe
dO3ShAYp436NNzDSdn39098k2aPWbi5+h1cOM6wvafcWG5i5Ys6QQFXNTpoZ4vESwiU1ktZWJgG5
ebKlyrkpeDR8n9gcY8q917heG6fcfLkZNfdKwC5dmca7zMsF5A7Ch71Lo9+Br3q93S1UTqFhDg13
+8HoMAXEM116aK9CJFfw0suUwvaO4oxpGJ/Zqch52gTvC4rOjxDLe00UB9hKn2te96izaukgmHRn
jfzT1tfA54thz1zZaEIEWDxcuwOhN+V256leGt0ym6869yJun0XmNvksoGzsDvsqr06MCqMTY63E
2L7f+3kxLzazQoA2Z2WOAT3dMcIGYCyJvVaML8PT96MaGr3eel0ifrSNwgrZxd81RaTggauEMa32
ZESMKEDGnT5QjvVkzFOBlY1M/ZbEC3/PirXltPhKnE+HDOr/Y4zHimfCP4BBE9o0doOa3DWQU9pt
vD8Ygg+pgva1zgArfcSUJXU7GXuhy42rGe98WQz36iEuFtlot0rb9nv7XJ5xKeNeT5dXj0axm070
t9C/21Ca5LPDjfoph48zhT/f5kPR1tmD44Gy85ZJoy9sTRR/26RrBi8Sy96j0cylxqouR72f4zPv
crRkUIcY+Xm4cVHKFgGltuxvQDP0sAEbpzPoN7oQ3HhaFgzR6yOSETbkJ1eNl5wip5ujoU30N+aH
hQmq/ZgGYFVXKv5viV0ffwoVrA3gnDnj0IWFiPjRowmcr7S4rn/6Hv+QHLpwbITKOU89uHzKtsPy
gzvqk4QCMqUCtJpuNULIIZw3bZqQw8U4IO5JpjK9Rv2QXu+2eQTP1T60TRpsYzdjOdRyyTuAHc6Y
NMNQTO7RmpdG92l7hXfx0kTAA1jp6I9evp6UkVpIoHvQn9/Diypg0+78UrgNR9rvok9OGEKfBM5L
fSMd3DTZO7UTmT2UCN74dCgeLdEVjtocA1U7e+4DvDX7aUDBIkpSeizBqVNL5FwLL4GdSWsKxJ6k
VvGNwdI8Mi1InwJpuESrElQfp5xQ83Bfn9/P6YLFehr2YABc5T2kBzRMvjCxzGXfInqQbB+4c6y/
zwZvGBpuFde9GbJkFqMrIDuVP7wPXcPxR6/HJVPlgATkp+yXjI+WGac3JYUXsO6s0VwuBY7cUYjg
Qx1wO4gAAhNuvlUJs0rZU+FIx9GCoUATqgeEJ9voHinDk4L/c5Dk5lVeYX50JUZZGC32cfnUJB7j
6Z+8RNvDp80G4TiW/KNXPLM0AkjItcCe8n5r88eryHehT0Ti7WhyAc7E+aytqIWmX5daQrz+oifR
lzS/hMV269i9BSeRXwI8IHbdxLBpf/9mmNmnP3AGPKmisRSqhsz3eGvwluzZs17naIUK37xGh7NE
UrgjpUxgU3t4fcrWA8XNdzOW0Ue5iIAQIBAaxDjH1ZUUeu6tvXtMaix63d1TMggaBDs/JzvjSUxO
F/2yNB6R6zFMedFB/5zj7nLpoRpOSnPupIvm3i5YRylNxntvbY1NhYKpUPld75pErdXJQAlHbq8W
jOien4zi+dVUr7KjEfVUzob0w5bsxGHi9WzeKtuHOkZIA0FmgFsRbNz5m4c/JYOqVZ3h2Y5dE3Ri
ic7Q11tNTfGQsHnx9n4AnwpYbJQdnf3VvcsDAOeBOTN5+3WvNIbfM373+rHTPolpbuQsghER+1gD
41e+FVLzo1Bxzii3eMNVS13GnW/FKp3lmSt4YrJsM78EHgvGLFELhR0tNFyUAqvTlMA/sb/dFRez
UwrrxL2RoCJmeXyfCgffL/AChC+TOkBYSz5r9iYF+a+aaDPO9siVqPT9m+JtY/hHDznnjwTet1in
mns+b3XbWG5um18fjXpWTJVqDGzn+jZ/snfe4Lk1wCds7zjsQt2SotpiPQ+2+sA5MPBDZZMMWUZY
DGjTiPvOBiHJ8HB/arCZZsD7kUYxPhd0T8Wu9vOn2sKUhxlcYra7XnWYUErz6B7AfeeU0EZCLe4u
2UniZn3/1/6jIVLQpUk4d8GNTgLncYx1B8bGacWql7RGHNCYSt7D4Hs9g3/wteLcke2DErzHEI2N
UE3Ie2vpDIec816zVblLWF0H9wBkDWi3jJcFawIWCuZNHp/SZKJImH0STnekf/l1u2h/Ti/CLoq0
4/TbBwBqVbfQp52eEZKs4iJPhAt0uMSGspnKuROir5VhoNzlAAQVXlIWknx6sik/ROb4p1yBIP2C
UbnPdgwqbI7Y3oXefJR2AMAiJDgI/110R5xBZWbqYI49ayo//Sl5otUogteE62M5I+y2W9dAgxwM
nmQqNZwKCNL8vm6hOwqRo7llEollKjB96iqYeZSTlAKu7dK2xaNxW4AVjXRxecHduDwbnGIkGxZE
HxYhnnTD8H1aOu8rgFD6cD55ojlGtgGGK7GGd8ou5TV+JnpwpxYAninuDq4LzD5DKE6yZsdNPRAo
8U/XFRyH0e/+edvljnpra+fG9fp/bjRhvSVVHhQ75LwccxAgYM92+ymfdavARK9nFJwMr1jS1rgg
rYfyoge0JaK4iOgxNcnMe/TkQ834+2Rux10ucjaOGPK6T7XVUtEQzCT5EqOCjmBcn1A7FEX0sfnv
l4JcBwpnufIxMrnGYtJXzJ/GIfcDoNhmjO5h9/wy70ekSV9XVoUeHDpHvBU33w8R7j3UsKb3nG2s
k6a0XckCe1HyCedyF5dUQ/APoPHvrUgyAVU7KPBMSbfRMXv2Rqmf2bZal2JRZPsUqEB5/1AMDGgW
J5K8TijKtkkBOjs5oQ/t4YaDcKoR5SfGmNA5TYP33Q2etxeFJ2cqugrQdwHbCfEXk9HqgDIcPaXr
jBVh15MftteOn13NA6Q4UnhR7Uv5b1iHCSxDQby2DUswtN1pPaKQBTxfzym6sOi/g1ewh0ydieaa
q2G1bPNytNZFyc1AvQq5meyJcjEzPJ3mX8aqdUNPYx4kVeaHFZ3XnTodYZPZw3T26cth5kkXfEMK
GHKqahHD99345oJ0TXwfPTonAwkLutbsQxCALNCMBhNq3UIqrHNJYcdhFDkMOkuEQ0VCf/Z4jGjk
2IPjAykn6uKX9HYyhU0N7i1sBdGD0DXP5LuO9u3Wmn1gk+xZV7mUb9RFDgcDrE3JxV662KWW17Wj
ri5E+cEx/IymydIgDgMecLhNtAKbvImtoMdemlymFI0g8MzNpEVQNP7lcHSdJlqtbshxDeIaY6/g
AgbRTMo/YGdzx7eAj2TKR+xUmmP/FznAKioAJZeoUf8Z6pCx7MF4UgE4maE7c07TKIYD6gHUk2HR
p5atlWCMAB31skFZ4z9OijNqt2m1jk7yFhGmxkPXkwRhsH5CR59lHttmfUuCyNkHnJVxBAK761lL
RxgwfSOBSpGyzYbHfqJyFwMr7kk99Ke41xTUqK8+dYvLgle1jTizL/ZDDpDCXXy9DhRTemOJ7kS3
AwzyMlovQnbQnOUi74q3xizs3q/N3/uC14lTlR867Y8iiTgnmaH8A3Z9oCq6EwcMMFOWGcPTkXnz
Zwv8yFgDjfGSxcWMnCQWu6N4Bopg/7vrTp2QDpmTl1ex2ghV924ZgoLR6YOZwH1gzfx6F7spvniS
/TLn8e6ffJE3goHyfFQFWPcRyFPGzYS3HKgWnvm/meDfzfqVsV+eL4lrqX02jmGlIimO/DWOIYyH
TuTaRTEEwNWGRYJxYLuutkqnpiFvR34skEINWeWFAybI2g2ktTKqcvYkZKGlQHtMkM5fDeV5MP1i
RxpghZJU327CuiWxRIFx95H9nFa1H8wHwaIFlp3H3c/LDD3eZ0L50eCDFX3vUXm9PZw2yuN0nBjw
OBgfHOgJ29yq0WQJJ3iJ6SAhx3vY4oiEy2Y3huJ6iRoKc/fZRa4sQy4n4xMAZPOz7QbDBbsp2PbO
5yyfTkLLFre/eZa6H7YMNTtgUVkhZfhjq339eC7XnR+5D9sjv90+Cn3zU9IE3cSZ9D8hjqmBEd57
otl6bZeHmLOgZ5/LTQsB0zOVnibIx8qLRNtYr8RiuLLcyJelbzbSJ0gK73t7Cj4gxoHiVzioxk8e
Cgrc6UjJTaki2HvUQ7D4BoSupBWzQuEFDma1P0bPSHS1cxZYhd0/t7qv5lMfhSRDH76OYpM4v2xg
FYny0BaOi0KTAvXEAezagNusmeoVpLzC0zWqJ9lRRxeFFdw6G2BdhtDFWfJlZx+k9gmsu9kr0UfM
rtSqxKKNLZeTDaVn54LssMQXR7Wta2TE30DzQna5cQBBgiifDqXvXnEDJhOGCNGDjEKEny00/vTp
DvdiakKxfuJiQXNbjKtCB/efkaTwVR6FhfOPA3O+pijShBeW39hwKJcLVNHoqtZoFOZRwS114TR7
6PPQM+myYprWja9Gl7Ygr3OpPXU98N9kU7BG8ewLC34+/bUe/hnm/zir6q3X0WSGDDzcwVTnFnN4
iBXscYJQoV0zMapQ4Rr3O5Jc6zqZVCtmVVTXfNVtOOF1iWrnO0h4nqoE4rYngXxHnkkSJ0YLQlCn
/icPxxca+Lrj1lOlPt9Cvnfft2rpHluN0zm4tbmjfUt98rNHuXpVNqwplN++2byIi3/WYbbFzO1p
Kn7zivThFQCjrskYjfhPAjuwlJhtPeWxjUvoFFGWuPgpYZOfBYWn2dw1T5O1xaYa5XZy89thn99K
LULXU22PjHwOxdXU+l0Fiv9pyLDNciLmt4G2opOQcI+VyJThCJUlKhv7Es8HM7ug+WnJYrPRWhLQ
hlhym6XgQGDnaA4mVT2ufqRDQaNYewAADVOkwZj7mONBrqFpLBMeXniycGnrhlYr0o1kPJTF1JYm
OM+EojdwfVy/XFq/b5oCr9tKjR2P3TDDJrvusWgBlQ5ItRw1cuYyQrTh+pXPloYb1beDIctHDryz
axzjP+CVEK0TXf8PyQ80fZE9FrVjdgG7TyhhBAjZ84N3sd50pFa6tzEf7zhXa6pYbuZ+uu7wugxr
+zIch3w82ZdYoHlld5T6IeYgE6fbH8U8daQ05ZTjCIaizK2WO4vzIgth7T5mmTCh0shPMFo1DS5n
XrvndBeATvIVjqTqqZa41LAWJb/WP8BDgV7FZPg87SBYK1z/m4uYVM8nOkfCKM0U13hEYKe85kww
kIEqqsdh7sjvdcdq+tWnD4U6s3YYjgu4TC/qSMZgWFItll3bxxkIZCun0JWUL1Kl1MliAKvvPnDB
oDmMAaXnmmXT8btGAnp9HIxQXDNsQdWbiQ+eIV3hek9gGyFcVk8TvN6wavel0L2yhtbTlynxNgm9
7GfqKR2FNXpHuOjWJY96oCGYtudUapHbV1ltY03ggCt1ANtEvA3pV8VLjqENu8mOoyGQ9SOWdarK
O2eK8Wf9rokAm7R4ZA9QRdTIP4nji0zHXpV9DZgFhsGefiXpS4z4e42RRGw6SSaZSps9C8c+0OWh
vp93BQGbf8ts1MaN3cOX6bJ81u4lWVPcXFXcd3phyugc7iVOpywO2gm9Bbuix8lk8hrODPDIq3gI
hJgKviDZk4120Ku1Rp4NMCtnc3eD7SjZiuIN0vneN6zwNqPGnkNr0ZZ5nBVhDyMGgQSvQI6lSJCt
M3ykiH8NrYKCwnfnf6y4vKRuUdkUx9DtEj7XCXwlaowAxCXAMQLzLQS93U9fSXY/Sx1FTz3/nFx1
f1lhNDP3MyDskpZ3TmbIssFKtAHpz566K2/qZDoLUNZxU/LnzHydmR5uTi4a5PJLwyzO1nFyv73/
xqwrwa21+dn+JD5pYmMz4ewKkBJtAE7PMZWoTrybrxPp9PnE4zVeG+5Jp1nDK+WNDcFa7QcaHkFB
JJ+kyo0yw2QG2kgeHS3sPoEc1ULK1f6NEDD63b+rkLBfhP/xjGnZpAoCGF7ADDJnVPsIrrEijxBY
b3HRhm6stTKdQKlI2b6VVwSaYHB2UIBjo34Lf+zhIFDiOJRoy0I66zv5uSyjhi6yIxkwKny5TWps
/uba0Otm7ChHshRMUGUSsMA9/CLYG/J/A6rilcb2xUl4hE64SnrQik/r8Y3xAgN0A1hyIyuyIyqL
o0Ck3smfioXebYVut+GvhcARF2xsKQuxuQL9naKL8Zm2lhXSOKCKU/Euj68YwABDPGj0lWKcLRLQ
kxj6REHRiRZqMag//wcnARzuRfZ6wCN2ly85A7kw1NgJul1Q/lxdqgPd4n8K8ZiWVNEGXNiNel83
27t3h/g1bVIEycE5ElsrvTTZ5giupeBQi3kAfcGMT1Zde2zNaOJ5inR/vCOmVyCvCSPUQp7AzJq1
qg/jPRI19bAYGt9KCZ7Z1qEKcPOxIaBfUTBDCyW3I7Osb7tQVWpX49KUbXqQnjoM+g9EmA+Olqhh
krNCCorAxT+zwhCGpCB0KbF8b/o5LfHJbW0i7WcDJ5hPtfwhQHolGKig4j47TsXuFQogKoRAfYnP
cpch6wS36VUpiw47cyLhYwr9Dknf9Lz6KVddQXYRb6rxvnECgnwo4NA1jGK16gRa/SquA3IRIt0C
8o/XD4MVxlKoN+ptxwSIWh1dXsA4ILP2PZ90mnaiiYFxaatISLLsTMpNEt2l1R7N7D2ntpBPcnSr
NZhNbTCoebmimcs+sGOdva79CvFvbIXkONdsZXQyVKKhBCngzDbfDZbJPnWAv+Lxl5papomlt6LS
xuiK9yom+ir2MPnd024kWluNaCKjTC8qXbilHPNVJTgSbYwbwYs745jv2YRF54ihKLNB4vY4u7Fp
X6NTFKtOJ3nQ/RuMWb6+m7eV8+PKolb/8zdhEL3DAwHU5ho/I9pIaMjiNqwDKR5Tfarozwe2eQLx
Af9GFej8NhLIDo9c8v+Vtt3ogYw5gdQ2LuxQedpR2EPyuhiJtkppTlz4xmEamm9guaXxqcA05L5s
MjyjlFL4NrcEteUHmDtiaobyyAxAPPwok6CfXGQVl/xHY+9h+AZBemzVafa0n4moJm9Xt5ooxj/l
VSKxFFuB8SAb71+UgTFxiBfgi3xanHFn24lljrTPcHZ2Akb53z1jb7q7qAhvJ7mTA5Ih58cVbHPA
z54CfXj0n6kFYf1zBTtwyqHcwGExfrLO9a6uX4KHaDTf/c2OJU/CdBDbyAdxRxcov+/YYB5mkDmZ
gDPRxN9qDOx9W6Ijr4V5Wo+eO0wCMTWmIpw1IBZYa/l3QyRzqSApPf+QB6rid1gszlGWdZ725ul/
6RXbNqdzVtubQ8XbkyVdaSuY/Jl3XZVLZULaTlX0rknEuw3WAKBfR1nM93PoJq77ppIODudFLP5M
XMFTFfn4BCURyKVTysBBLI4Gcx0Zli4z3/ROuSZEPMYh3e/icRb0q1AthS9ZPvhzd2IYr0M3dHsG
AsTBiJSHW/ISwBOYYpicqFeNXBPm9P+7kGlOpaKrDdrcy3V7iV2fkioToz9+JCQvaJzBaYYbplJT
8N5T4lk+j41PgGZkc6V3oul03f/b9/YkPhM99szGbLNKjs3cP/mYFqDAUz2HvqQfDlmcilJJUPEA
f/bmCnomKjxTkO7h/yAQ2HTcEdLhZAf/Y3Cn6EE3qKJ53zjqhqFOLiD75oKlgt+TvIUqS88Tm74X
4GFVRpacWKq10EhN4sABs87UyzpdEqg0b8mtqLGO/v5tIKtyboyWVjS9V28zPUCtoH9ztJgSMrjE
S1NALYmd0mAjmFPGBtS2yGkkCEBSid8oLxj2UDdrE5oWjAJ/3e6xn2tVc+T4pRkVqd93rHf8m7tR
5avYiKSe6SATDlFq1EDCCghvudfzu1hvHueMHy8lZjr/VTSXbOMbGKCg60lvk6vF6ZoNi/iDZlep
SJLef1Tsc0bcBZW5dyMpNvWf0eFaQPyYIN9EV/xg6xBRgxxUlTw2vIGRNKDn/kyLQrmtOgqo1d5P
HisqbQNGYJ/HCLhWzJc9O2rmMMYN/erQr6I58envNdW24VE2AXR14ErqnV3smzsbjTJjZi1gLV16
oNt3kUPVnGiXo9WPQALbVpaIEtzrM4ULFoVdqqKMROB3fKF60A7c0GgScBc7seqTRbDfsCL1wYDI
X1UPmXhQ8tSjgUAZJUih5s/2jHc6JoRt/o2ILOzuQax+tkEVYHcBu/sPMmSLXtP1akN7Ac3M45lw
h8Hv3VsdOnYFX5W910aYjF7xCxDutbNTy+o8JGYEXM0RmieNhiHITP2Z8b0uguXArz7BR2IKOzD/
blM9jXQ/dZgnUg2IIOhGIs2c8BunTz2gbhNPB9CiPOXKQMpIxkgTtcGChgBSNy7SJJLV9BI36Ff3
M98xjQsAXLtBwkTBNXGxGaQkYu8JyAguWY2pXrebvmyzh5+EmAl/gyZcwU1YByju60vmKi1FXmx7
Hzqtipx68r9wi/lGsbesfsjqXAY9ewEMyUEb5D7+AzTeiDL7VRvAmJdbZRxs/pEeIkbmvn5989AH
/SOjoHaSePW2geUe1SpuJhkLdEOd+S2jTa+N2Y/UryGmDBaFmFQUFmgTACi0jfZt9N0e2s5CUwxG
lFNfOTuqAwdREMKKqaI784bZAIhzbXG4OJ5SuA3F4rWZM9nn6GTNVhaLtc0gdT6Sc4OwiIxHdkTX
ll8qQJhJ+XwAZ6ck/VdV0Snq5EjWcabWV3SrwHhlVAeQo8CQxR8EN+clZKqMJZU9neAfRjcLi48q
3q7PolT49hkGCtWmo46MycU6XpYzfIuXsnhfW67ILjbOHGK2b0iCd8UZPkC09YG8KPQGn1G6Nwey
DhDZp0Bgx0lUyVDoghO+dOLAuSvD6+wkKk/eGmfwnvO9LgpJ00hHDGQK7DADIaELzHtPd83x2fwY
6jQcl7WyrseXsuwKpvZPeZuUwq4C8+724Dom3gbewuqejTx5YBvfei596MMt1H0bL1RFNcRgj0gf
bW9QQ3HncWLYO8BYYNRxBGFXLZGZ95GpxtmoQVMvNbR7S9m7kK08oV548uJnMMeyMY6hEUX+D1QD
HEKAyWxt0ZIlpaGCZlzS9PKBZ6YMajJflNollcLEGMY4N71NF6Mb8o4qhVINqWQLDnOV0RIIX7mq
FKpmKYODlFhUh5cdnNMSIn9cXX5Caeg5RCAT3fbRXN+8Y0cRPah59vH2knho5fUueQbpaVcZHNGp
k9g+bX9fEWku1kSH4pHgeze87XrdPzide8p6q1vnPnlfd37nlmlx8+VHrvFsW8FbF8lGA1nlf+6Y
TP1jT4jYf6p9jcD7pEraDxWpxv9z3uT0c4faGeqmczq55fDm+e9GylUC6PjO/7Qeys+nR8Y02nWL
MzQ3nYQhyoOiEzpwpya6Y4fEi5+xHLMCPlC6JWFe5QfVcSIeNZDPScfqCsHuKOPiZ9GfhLKctK2H
nEt53xSIIByzQfXpZA2BfXOY5rsLN8TDlAOx49OTd/Xdm8BPQeqydw0o4ufjD/2XTS9GSRHAKU2V
1CTjiXvwqIu5RDAaoc9ys5ZdmeXzQZGY8t8Kv+F2bT4JmxRexwm4PmLCoQVP3gNRFcYEo9TSqDQD
X4AxmprbS8haA8lKkYgPXDelLQ39AlrLpUCzElvdS44ca5IChZKWp08wrj++IztagVeaDv4r/Qqo
8oFjsuV+E82jFM4rzUhpThI25vgZLl7H8QXH0gpKPo1cZSYjpu+1nJk8UPJKRar0So2yJjgA9Q2G
hTPEL+54wASdHjFYNyXnPdDzT39bku0oIuZu8hQrTno+veF+R0qTZXlUlqNvagwT9o3bzUrn6pMp
3C1NdxrnEq/osXpNt9k1MxbNsqrRdmlgKJJTOwbXGp/D/kXaF40ROAZZkH03SAbNT53SLNmQo+L6
jNFNdQSMlDZ9KZf2Q9VqJ6nXNTkQ2lZUUIBLt4jScYN15F8Cnnp0PLYnaDp9sgH9ULRV91yAIV2b
LCsIrWorbbx+PNF9mZhaflAc6g9hc2wzJ3OFSk4Q1pxV7nOHvPKb6J3WYmkKpClvi0uhvOKTcFcJ
2uVsjxerFoSmG9WJ+1oxLNSYQHQbc883oeOMP12oIJSuKS+1I/uTbdjqLS8nN32o5eo4EmtH2EnO
49VMb+28b1UzfeVX47imO3r8y0yuA0ELUfkKuYaJwhYTPc9C8O93A+MSyPTII3cZwhTyKaROzLbu
yWIQkqlGtlO6vXZlMVbItg+XD9QFZ12TsjeeyQlxNoi/MBfz+pykRXEQvmUxOTrmZ65/Hrn6Qcd5
dZ1PV4QNzgxROZxoTet+YSXx4zHxnPJUdUEQxUvkQr+iBzWNoPLSQ9Bm/BuEdf48Aswdv5jDnI1u
w81Ct3CJkkahj/Ct2fJKyTnoNWQMW+4ZVlDUOYHCwgDOABTPSREF+Kh5hQ3tbq3tAoNyNSFTNJbd
O+XSO9QcbC8uAumequRExnDvhrg+Tfimw4w1XpDv63FiuXMnpW9fPG4jJmNovbLId1ShW+Lb5K4C
w5ifj7ykUdlfilXb/twSvngDgcLAR8Qv17ZBjA2Uj5l2Pq0hgrUvci27jG9abQvqelmqc9+hx99y
Nl7PPUxD3jG1idL9yP8R81dKvp/RGgmvlePbKPIiCQ0NqlSCKGtrBGR8USKnEj1hlv72CTgow8Dg
/o++QsuMJ9BleIr5Ii+2Es0fFqAUTKvaWKKDhUKNW/empkLHkqJKvqyn4se1/+oRvBblbexbJBaa
HbKqdtq77oPyUHt9Z2wdmc/akgJ5vCVEhklhNMVA+pWLIDYDvdK1nhEy2+DptstAzg8dZ9HolnR1
kcbHOt4DVR5xCuIuPBHzI8en6g/xDUEdZt+vL+IczZU5R4rL8KLRKx8fQKYiNffYrS1oHrXCCpB5
tgQx0IW4J6bVZFe4QP4Nj3frhoXUkhQIBVK6j5Znfei72cuYvKd3DsD0CVpS17cBnA0LYzHvf0by
jm7p6K/597UGMF3nwINh8x+k4cxpTyCrSNqC1ypdZygPmWpY47Zo8HJymcPzikf9BTZxvogQfx13
t0x9hi/yxtF4tnr1V4ubmoQ3m+BhWwOBwGg3n9hQzXGx/lR0+mqlaNOUer7j7oKN/D4qB/6dkWc+
E/FXAwbrLe3KqJEPNj9m/VdKTKg4ZLnTdF+4CGdR5mT5v3F3blCMFxKcRO/Mcw3QzBZRxjUhyO0Q
+zj26ig+S95f5kL/IqsGwckgxruzJX3xq0RbzlrkH2IIDMG+2ZQXYsoAZ8nLLRNexLR1WxvVhlOs
Q0ItZsQfUaB5MZVwjOFLj5tTog56k8PGYp+htpMbyFdzNTCVlEb7+HDjZ3gGlso9OFUM6Z8pgtni
ozhUS+BavAmxqhTqKFlaP4tAJrm8vih2B8RYC0MkPG0GkPll+hpqHVudFFpzlfFKkBigVH4ZISDM
SgTHBRUy7hCxxnER88kI792kgyJO2J5A5CDH94QPTP513NNuD/BMUq4APwXg4orZ588ZBncJdCw1
sr57/qQBvOaehFXhkxTL9cv3G0f9fQdsXArrzWVGOG/2EDJaTcDpcZo0I4DujC9JQPlhEmibqbJB
Ce1CSFPLSdRavCbZUmSFeN1A8LLGWb2yyPchBxKhcfMd8lxAKs+b3B6EeSE4PArDbXmnTlNBNPXT
a4cE3l1XJj4rwwSvsR5/fFmp4noNJofvemyMVovL8N8JIvzP0SIAexCAHS8fj4h8J5m2gAQVy77u
2UNtVdqnw9VljyW9ieS1Xoekl4xKcnRBXupQ8KxrcFYQA8A9Q3lCKoUpun5iVf1oy5UXBwMOvtim
e30WcM3w3tpH9qoCgC0LK9r7a5XUoxsi+TnCJo9x/ZaNcEBopZKH3Q/+BdUm5JVQY8az/o9lTjBU
FXd409n58h0UlEa1T0aI5TFKeY7jJ98wzrcf9ZwLEOP2UlidGYkfkLPH4wkb22UEytBsVDfUi4E1
rIIAPXyD67NcRobHEehx025E52Jqxavrll26YbMI+Wn39gT85+FtJZcPDohP1Yh4Bi/za7wRCwUH
SttYwyOumeRJueDUhNQ4gThlnADrYKwdzIGgyVHXHfQHC/G9wjeSPPgMdkNf8BuS7q9GLcUZgUtQ
6s0k6XHyXQcUUqPFLtHVZtXqMb11whFTRN5rq1x0IO4YVCh3LnHmi5c5NcRsKDO8fSVrwGL3yc4l
s7aij/zDU1J0tSt9ghh7gxaAyrLfqcAgyq1T8ALT0smfiESq6BWRfjbfGlS8vqWbvY4BoXcJGCDB
lUPDmqCOsk42uRT25OsyWH6MnLkFvu+vLq663j5RjAxt1+SL5+xOKdxVLLmqhMfuXQk7G17ixXVB
TLhpPuo34E+qoY4MeDpk7FREidtV3wrRrcDv4M6FBa2KHpjJ0gqZ9PQ1VzqGgI8W1f/a0B/XmOwA
XzAh96TNQsJ8jN1S5z9hybN0oAJxXOTJdFG+THeeC1WuTVF4B8nZq+/QmBmnNuAc0QT/jospmdwS
pWDM+RyvgI6bJZuBHaZGV0k83UvGaC9kcYfZGMPedUVl2cKwlJs8V3l2em6KwG8OOjJ3FnadlAWM
eH+uZdicbS7MVEfd6XaDScSluOHWKiwpWUxKRxZDzI36LBEqwcOF/p7ES51RLLy47eyPE8ZPt+X6
EBDysKVOKtX48oZlysWWME+UJAtqXr2nVc2LiCeh5BaRng0JLLEo/rgcnB6U5QCEUlKbSISD4LoJ
WBNtaOQ6BA7GyOB1BZfgAYo+3ddja7/w++j+zh6N699BKSQhpmvWFQFFG5cFr4OJhZG8A3ZD2eiV
NKKdfO/1qf/qDOoif3o4R2s0HR7HI7FyX8QOOX9GwjuSZbnwELsble4mG3quNGQg5T4G2dcMYfSs
RcFYsEl/UMXJ68dZm7yT4kw3e27LxrrMgrRKjL5RlUL5qd2X/KOX4/zzkOTHMAqHXgqAcvSonUOb
NkFxEmONLHjrhVI3D0cvDbxijkBX9fY3fDfQSW8ht3QLMZ88ogJeVP2GOXiinRxzYWDRjUd6HR/Q
WICox0irprDcdJG5UOt1BKzsJF9gzA8/20a9ttCGq8Yz/mu52/sodHvndxw1vG9KJGNYNxKHzJdh
Nle0ToearZd8Tw3KQbdwj/1pVecyA63ZgomwJ7AsXLflo4TcnJFHmd7aYWpCaaKmYMaswfldj1h7
RfsZtvjTEJb9u6mqnxgDFJUTXkygyotz3zmzEyNiw+3VgZc6BlZMJ4npGgck80sJ2q7+yo+8tQ9y
jE3a37ecS8gKPBPE7UwxQuG9O2yvbpXY1Ajg5ttaHhi6CQ4x1qNvNynd2JVNQeZCJBhZ63TiRSBa
uMRxz1hz0X+0XbqH3A2Ddu+NmKOxzOlp3yoVoTSYHrFelWZ7wqTqRQ6IcTFy9WVcoePFxUDlhqhi
4PVNU7t5gBp18deVeY6S+XxoNPhGK1iyUPOI5i1Ks2hxdXseckz7XY3uCj7qA+npY0iECbgxfPRY
E1JmtwMmG7kYH7HyFgVReZesMEbggzOaR7/mgIx9ASqbT2/cppqM4NXDSqH8tN6zbsiKQ0ckCF85
4jWt4zEcbv92htMTzCNGYTL4NLgeYkZco66KS0KQSM1A4RCoUCAKnjFuZkLIDwau5kWkC8EbOmVV
gsErUgxCSJDSeIGgf4A4P7vnfmf68/G7TI+mPweB/nKT5NFSEXWRRh1lpFTZH9o3WKPzSPzurb94
s9gVNYQ8KqqbtnCP5yo2LVUMFdHowOUCjUB9k9Y+oIUQHlf4mrMkXqqQJVQMLObewntGGoFh0bJX
N6WQdI7Mw+bcBCyZrH09E+n+XwOMFogzO+ZxNK37/8uTCQVQd6nRv6A/5qW8Yo/VZrxqMkyFsN3x
BhIjQtRSs/whd1qK50tq3ENGsNQ72iuNLnQjeaopVy+picLvN+GxMDaTStSXHYmEGXoLzRURDYJz
zmR6tsOJV2eR0tZqlJ/Q6WvtoGitpaq53QecxYbHaVaCKbTyGdBqZElVBSEbkTRC97YqS9iCRVnl
IQxNb8C8xWiUCAxNS0ZE/GJ7r5Jc9QAertSsl6X+AvgUCRBk0rKxlDXgpxKffCtUApooKXetpU78
IO5nVx+RkPFUFb6I/uMm6pMKoi8bUN3/NXx+GlBXcOhRfSe7BFUrfm7IO7xyJjC6LImEDbXqLz3Z
c5wWDVZ7P9e1xQD5ooe35vGUw1B0Tx99io4dZ02PawOUs1rZUewbLdi4p1v9pVfPua+17+OpJRyg
cND9Mk1S3ErFGdIyY0kV8Mu5kPfPiffzfB6lAJBinT06Jdcj2iN92bH4IgFjZEbBg+CG29BIJIe+
yOk2eH3K5ctQvdJ3erdn82oR6Un6IJaJxoACwuDFeS9hA5RVcAuXCy3g2vWQYMhd4Wy9EdYK5cSP
uXopRLdjS4sjGbeQ7Fprd9FUHJyz+zdm6c0/wWgMDlbBHy0AbjyIm9QjzrKE9EbG1x8bYvef8CMS
OnZCLwYoCtbLAF92rTYLc4J3OoCBSD1IPsOrCuI9PVgpvRfaU6JsgHvs2c+1KGVcfEkaWxhsqEZH
LUu1txHdqxRzRL7K8CWQGQ6O1NezA6TM+5MnOtOmluUjCyt4lmKxAQHZA4usTwKlWsBMfiWNp9FQ
ztdV7BEhkyiHynzg3aPDAx3gFFlZ9c4uC5h5oU9hbrgPeu79GMfkmavsrvrQL5jxuYOVcbiaTVM4
ClJA5ijGnI00pykhGRavFp0U01zb6R0SzL8xToJDP+Pbvi50gT0CwPT8vlRrYNqE9vat5ul7+lpd
FkKi6ie7MSrFLhAaqJ7Y+LOxTW1WYVRjXlr+b2IjOyfsQ5UzhzgLDkRg0R1WN5Y0+OSfziOXwLLk
/S7e1bwEsNEgn8p2w56P/zhzK2csPkbab/+dvoTvAgJzVwFc0RZFJV0xNnCmBX1dw0tbhkdolPMZ
1LrVa0SiIYFSI3ndMXnHYBrnJHUwl2gsAKbi3uhORUTFR0t7uNVMhIaDCLMyvSGmaYPR56dVtVw2
x32Rh1SxK0rQGO4nnymBiv4DzQHrm5nUZBUk31nGV/JricLv+GatIV4k5zWD7rhOw950JaokfPXo
p+fUUk5oaUET+uPEIjxH2KfyDq5MiJ1V28nPtg+agPWgZ9XrtEHW4nT9kyudQgFjmhauWjF0lc9w
MZi/vDBcFuNXHQq3uw2+4ZqrhpXqHU+eGKbxzg5z0Plz4+k5RRpyMtHg5Z7hXXcsbNvC/PuZT/6z
bXV5cSH5ijx/luirRukdIznRNN+rC/EOApNGsRzUJowhIbIJuVsmqWcAZOUor5qTvRSqxU3dsw/Y
UdkU/xfy01EseHcPI8kYPZH+f7EjyTfdXzYzsu60RrvWz1iHWeG1sSRBZc/tl6W5ulkfohjnJu+a
C/dXkKyZjpZ7+o0/B1hz63xKIjYqJCtCeDlqLeYS6Qh+8WcPIixS5DQj0TTlpTTzWxkk2fTeB1mn
zPmjfnbpfXAa0q089MxwTfwoSdPWsJ/JCzkmonQQAecC3YjjGn6Y9GPJdAOFIBt6/ZIu/fNyLb9N
OwhWD3s0b/nysTHGeWdrVYGPkvP9f3U/qiho9bmXq3BXoh8DevfZ1XtmeGGys1UaTCsKeFDxS56z
aB5OjA19rkQTaPTd+s7xukLPRUypF1yf3isYLMZMW12Ju1e41uuKrgecVE7iWh3KVqcflUEtngBL
e22WA7YFa73ppw5MICBCfApvIKshKvwRzb0ic13ECc13EcSXT64kxXtBeVzOYfrCzHcPP/vC6k0B
0OGVIvfINcjr4bIWb7DlDFQhlLcZeGBhmevV4KHaON+TBU7Npj+Lprau3GZYeTY+3UtG2iMEKVvY
4E8jMsah9+g/C1E8lKqoZ+Mfcl0gBj2pXfCdh+x957xy9vFNdn0coFWUFGUJLhjT6yFCjakb32pw
os9sJBpztRGqUM7InavBuPDEWKrYViPojQ195s/1br593hcCWTnyocxst7ExNLpVnMpjEQjvIDmF
RcR1Ncyw++EnUFCPpdDtZszY5tL/hrKTYxF5otfiev8lmfT6qGqUdE384KONRs5J7jd2tV/K7JhW
0LtBd8obCsKEQdXuPBFbXe0u+SwRWyLYpHeh2U7m5Hjzum+VWHCou22TFQ720PIiBjVb+oAKzO62
lR6im5IX9CRInp1PJTx2XrLtSIadBjmeBYaNo3iXyPyCYD+H7NvB5aosToIf12FOGwDTGMR+/hF9
2Rw2Cj+0AOb5stSjxMWXP3VgYx35692VmFsNTiC3mlaWDJEy5pBCsHXRV6YKVbQh4dlnHt8ni7hH
UhNkSQjg35M73TE3RiNXnsdsFBcpRjMb3e4xU5BctHgU6KvFyd6uxZMyliCt0v5IuFI3tDdl7l03
onzynis5zTG8XdUy3Z+OJcroGTEO5EPtWcDx5bYapTfDZ/OStwyEAeAvOMpbs7Obd2ie6rHUIcWd
Xg60nXm9Oj+Nx+3c6dwxPkBErm5/KaNwbaEWzCWm89bwrD3CGX7m3ziho/9zgK4VzBE7pSGC4dpz
0mDdIMIh3axr/l/3QDqUZN1vy0FM/b0MqiNGl4r5P8/83s8CU/mNvSFtVIoXjgs5ngDClk42Ehjy
XRzEYJgBaX91s65Qm+60aoPlorHceabQtH9Z70y0U4UAcaEf4rwLOrj8n99wD+Wg6DU54YORjODG
aZu1owXi+TPetOunyWnfjP3H/1zDSN7LcY3QM57ZxJm8wpNCO4KSjjgCQyFX6/IWi2s8/edMkYSV
K6off9pKZxdAOtWagBvxcyl6ObZkRBOhLzF3hXv/GrdrcAEjpdj3QEg05pcMddtK6WHZd8vxN2SP
mubt0BCNd579iGvLBb0GugC/Ge0agd9dUXKUSKsN+MBPT8zKWOcT+ie0l9SV5AtPwgmKH183Sso4
qjya3q/sKYl32xTPt4grauWj3sDOx1DMFL7cg2wJ6jc+7IUyzSWggzBvvAL+R0UvU7i/ItrBQ9Yr
ILRWu1cnsHrhKJruyfDE9U4EQ1GDk+L0o0FBaAK8O/pXy0NAUPoej4XbgkMvNc/rkxp8+ax4a/kK
XDjclyx9xMvdCcB3H2+bcziVCRq0mG5NePaW+OGnnzy8dfhx5xG6GfotYB6PnShrhvPvVd80c5DY
eDk7UW46LjeYUHf1c29IZHx55m+RowqC27/Y73Q0nM9CbcnPveWSbf1GoybDrx87O8yzd1RvVayO
KtK6xUGL0LG6pXL+eL0uOPHQazUmnyHGYwfsEz/a1E3ahxSLCO/ShvORcP+GFXbyjXnBJTwabSj1
7axPfdPB1adeDE/+2ggJFNmEY/VlE8dAs4Y3LjFJQP/gjwmDPLZWCfGhhi1lu75S1Dywvog4+WRS
G0g+JgDtdbEdzT8U6e/O6Z8BdsoxqML53EdABnfrwVXKYavJU/1KYNiMJqngGO2tkHPL3bpNVU7K
WOwo4o+EAqcQ62cERCtxP8Vbk937nyi1X9gh+zmF8aJMkzvwOnUHuvLW8OvPzBdnzrki1IYmRSc9
qTP7+eXsAHxjvi71CAqpzMuzjAL/gAuDw2Iv+60RYTFUbouR6F5J5Q+rtJ8kRUuNNynfHOgCEMzc
B9UiEuo3TOhrTXQYeo2NuP56+Sbhk4vmV/Vc70RJDqLVCWgXSBe9kAFNMC+dZkAUAG3HqnrIAouc
riXfpSbcd0KDAc3LZkZYOlq/h2OY0n0J34U5TVUxxVDLo0K5CFag6trXM5nfAGEVZbwzHITVIHuy
wHtE27qZH6H1Mi3m4Qn5gwSozpgp4ImXpNvyBrxrJStmuM3g4Eis6RJUvU+1S/+QJ9TQzby9kumc
lyd9GiVvJGGJ3BJo4yHf6Tv9BdPEa2tf8rkcZ3HXiUucLhcJmofa2o9eWzj1Han8FlgMGZpYE88a
xuLWZ/5wJk/GOv81fCJXKIJRiefxmJl5NV7c4k9FgnYW9R3eAjYOXOiibzCRLBIHbrwvmsqkjcrL
JKyltl+hU5aRdD4ehpCgEYpsOK3iOYSFztUM9+Fs28Mj80y5kSpbYwPD5b9MF420lp8vTspcEkzR
TLIkxaKzuwhHbKMj63WmDXuAfcN5uuRBPq3VV/ESPu9rvguvRyNSuqgcoUIjbZongNxXHtJMiGMu
iVgDhE+Sw+NqTf5jHJWFvFBsp6kxrDtNhgVzj0oEOT9ZagEbfb5ThRxrl+rcQiRx1EGM0w8qmu+z
nnIlSiJ47xdNtVwOg/YLhgiFJzrE5qPI/Sq961Vt0NJ+eGXP+ovIhYy6Ji3RyQBJYmRISJnaATW5
z1+IQNim4bJoSDdDpG8XmJPCNWFJ4dPmSGi9nsb1Ikdvi9ewQEeFSDYe6iHL02YsVEqbi/RmsyEz
GYzLVG5zNxhrMpA/iXUa3UmjrldvVNqBiI1jwoV3iwR7RWYd6rmwecwF1064yVmaRSRPrccaUL8d
+RUTzp0/LMR0iKulSlYXIyY4+WyfIzejQj/32bfWkNyw0FmH62322645RnELHv59YtC/wpz0Jfjl
081K1vUKqLE3B8g93AAyFw5QJYmH15u+ZOY4BMZ/yQRHMadg275z5eMO5czwJ2HvBz/ieBTmybW3
QaQjC2XUkbfB6Q7/x1AeL0V9dvb3G1OIewOfRdcadzsn4CfJzT4oRuk/Uc8Z8x3ENbDRmxV7x5oe
E71tzVMCVPU8qUVfa3p4zKn1r2SYVJopVknNLQj42C1cq9DZuDLZhj+sJsFy34F2pAVVR18SAhYr
zaDaruAZQIzHoRYqx/x2TfhElAG5ZPbT3gvQDIcsDX6SA+dY8WlcIg4CBF9KB7fG/BSRlFqA50Dq
fhftGby38jbu2YfPChxkGe2TJJmLIN/4IS3bOf5QQ11h00hzZAJ/x3jbFO4lfV92yiIpwZ4ueCtx
jksa/Whj1+qobMHxi2OOzNzAYqfWPdadjdHQMdCpCBSe9u+0gXdzRAPNfXK1YRdt06oOOpd1LgX0
H+iPveh5yJkneLo8JLhisPxgmHcsTobnaKc1FsbON48X+CsvHXxiGqTM2pV7tFCRIjQvQHgguOWW
jWgQvVWwxYnRbWEcpWRD9j43egLx2RGgj7RhAe04sbtwEOE8+/dOHFBx3QZdLGK0E+AZTMtT5U0y
ltwf9BzIpIuE8INIeb5g93F9mhS6dlehe0cvZtrYqnHKjPMAFn+e1VltCEsSi0dGVjejLBuek4/J
A23D6o9af1BB1zl3Ga05pwKub17lM9yubIJd1AzR5CIw7Kjy2Jsev/tIZK0DbJinbGil18WSwlV2
u+cIBOaF5a3KVAm4YcZcAY0utjDGStN8cO7cqftjaD3OZGUZlhUJd6PZLKjzVx1wstDJF5CqFCta
lFyUer6OQVMR+4ax+4UeVF7fdqurOlNdCYrmixRSQX/KwTCYLB/sV13L3LUmYYpoaHTvt5Hcvzc6
s1N4NymQZ0PYdpeSlF5snonlQr2MsSJPjh/tu4wYaJMqSlnUQ+cXvrx6ctJSSF+i1Js9o40nYCHc
VUyaRFjsc/XxgDE+H7wAS6gBV6q31VI0GSkmG2N8sOhIeyorHAYubxUgrczEb9hGqRojnVG6Phsm
n396NTEMfgR7/v7d92OA3x+cacU/geG3gtmk93S/FajcLhTXZqgtt5iP5p7s81YEDDWdjj1j6GR9
ONSGS+VmfAYrElIFqiwuc0ujUi6oogT0m23H0RdRy1j8irIwB6qVHv+eZViDdqccwZojr/w1OJdH
oy8RK+ACLMnVimQz1ZRQNeEpX0Fm2rw+ZNIwJo3VNNEpWvQ1biavpVg9aBCBf+B7/aGF4TtJBUfF
Lm4M4OaMOY1R8EO6OTjLvWjxPETlrAyqnWNPjwGKufvN91RTS7IB7ENgMEsQ5UfgVGNctinXR14m
cCmyw5NM/pzMhvPUI+Pp0iD9Iz3CFNPD6aoiPQRHfFxwPoOGOqjRPshktHVDidO+9cEmlqiuNKN1
erQhGf2U/gNvpos93yI4hJBOK1aZ4TpnoG1HdZl7s5nnmL02HgJo0ueu9pT2C78+MgMuN3U9TgZ9
k9sHJu3hvapdJP+M+MioNl8AoAWM8Elg+COmIHdlSMvYODAOXvqOqcD2j08YZ0GPaXg9t9euwEUe
xj988iw+3VasYnYmfHLpxwwJ2rnIwaq2u7rAyt5UYc0/sf/RQrlV0MLVnrZ+40dUIDMlpzG8REX9
3oLrGkfNLVakuBoiwthidaHXz7FQDm2XFxxjHBwFnBz7aBAW8lciliKUhWOjEfwbx0ho7SgNq57p
hZfFE1UafNJ35SjANq2maUUeccPzt77vFnIfICUTuRwV0alH5TObMEgZbY2sbGAyXbsaGoycNguE
1ikaG3eFN5eSis8OdeaAwjnLqVaFExB8Qes4Dz0+LopxUJjHQbK0Flxofw9xlKjogO0aqI9kXC0N
fKtsB+b7FMJB6YvNx7TaOPTzImvX0W7BbVY2FjhTPOmQgs2ALUjq694bWu34YoE0ix+BGeGpETuD
mw3BIpv3sSygwXTujWCVeB3zkphfzZmCKR9es56yneXj5ssGunPmf3S3Nd1MBiDnypPIlLaE72PA
220aVD2iYFDz7WysVLv3DnviDIxgwdU7B7Xi0wX5IC/adl/fW2clT7pzYSY6KhTw8ulvJZjCVf50
Zk2dLb++u4dFHZT8tMGJ0GpC+7rjjCTvFeXsUDeprePQo4NekftrsOezk7CtP7XAOiwH8Dx4bJSh
5wyzO8XQNeyJhq2r2NORK2TlUK9WrQTtWOaGuEKi15de6hX1zQ6GbsWUAez83tQmo7S3C1nW0riw
CQiLwhbpeOuk7o3P1+HLjuSWDZUNpqHAXxOphMDONZAbQNsyJJ94V5B+9ecOgJlI5XhJmNEirduJ
f23RQSJpKt2w8kfZjjR+xpIFduTUteoG/HMQkkRduMAkeqQ9jWgGP568wnyc9O5IxQkB1oJd5uaT
2A7GD2gq3P6l2uHsCkYVR7fVSj7/HdJKRGJW2foySbe71nP3fqqEELFVH9U9+OBnU1FYpAnWPpjG
10HyyypqC/wylRaf5WoC2uAUzU5PukLuXPtr1m2A3wxwn3QaaVDQfwA4BOCwNdDIIo+ePCYEuvmT
HmnpO4ZpWgYI6DSApmKFW2Qvbnakj/mlg+tl4cAKoOEG9SUl+vsVF4q/KTZdZGxT62IAtxVjZSsJ
wLFfpyPOIab1DutAE+dMgEcXR32i7JQF64h8YrA0Zm9Jx18oupUaNX+9plTDnacqiLdIYLnx03MR
zIaGdqmFG/eggoiKxaVGkYH12fDirk76AZvQGCEN83Yn2e8uUMoDmAR6LBmiJYH4EORz1VkPvneu
+/bGiQu7VOn8kPuHZ0Zac1ZvDE6uvFSxyEe3ag/UITB8DUgCV4EyPRw7JUvDkZ+k6ESdXbN5cSYh
9kVTcXK+R8ydKJ5QNsAE412nBkZr0+PKrt44YfyFtVVUIgKSZXuEevqoTBgKkNtq3D7sEbwhd+xE
2SqA2rs8yu8ygIkBDWlA0equHZLqt5LHxTY4QFCLMz4RdBUIPWyBh1yXDpOa6rqaDoY7nK/Hp8yn
gk7UQb3Tf58CZ1fska+x6er9r1u+ze5NeKLZURHvMR1L8+xBGyHajpAk9MRnoK0sL/M/9DozBkxD
FCa38WP4z7uY+sFvCaqB6tKFKLF6CfjU2/BXuNRtspmp6iZMpHOTpLs+yhUh4rlueBXj/sfWiK4+
EEn9pO4YHsHu4v31DqDzIGiP3rl9ErA0CxuxWD4OfJsWkB6gSRKlYletQuVu2TO2s6Wm9Rw6inT3
AP52xJ5/7unw1VdkwE5M1rNJsFEhIkVPkLKkU36x7JveCVWB8vLQzmyK+qzx3H6pgReKbqimLSt8
u3/QUgg816smBqlhGmBx6Zvr+Tvrnl/An7T7H8KgoouGu3u+MbbqYvHZjCJUEp02Bk522fd7ZI93
3/wga1Ntf5TkegJq7x1k9y3MVnhiMFQ5HG1lRw9mkNk8/vRdyxj5ycUS0jLHrYbOjnv1y7m1TQzP
2wioL3Sm2O+ZMg4f7nDesvLgT9us2zbGi3ih7fXfTaa+/9KvNHwCfTolPvbRIY7eWvi7hebHagKT
aoxdiXsGHmlDtzjqzT6TGwqGhtERdESuh7bj+pvDzj4YZol20P7C+FQLtDwlxflW6MukldUTHnyM
5QOwnnT3yf9LxFDUb6GzQ/LxcJo2kkaMeMrx2l53OPB/RrXRBEmqGLnnZh+NF1Np89ki8xJpuQci
jb6tYs/02fc0QdMOz3rU6cdvtzMAM/QLHL2X0SYPLqW9K17LolPL6HIlyMYmuDHfW/u5FMf3/NnS
8uA4Fh65Z4EAOCdrV//IpbsnkKk4alFliGwH4+rfhiAvJMVDWDtsrkPF/pCUZ8PF4sQm2pCwi0ao
e5C0pCDwUVRfVl3uo1lI23ThapDeW866TuvX0rY9czB+DLdjL1BJPeBZMAc1CqYRgKtx/0Twlj6J
VED0TdQcc5n78vyRNavwiewxE1cXizIM5uyxfbmuNdHdBZ2g5aRtFXq8Rw3Z8A3gfpJ7T9ZMr8oF
d4172KcEEcm4jydzNypjChZUWwYun3fRD4NVMHWcRGXTp7W8fdysHYE13dkssbnMlJbaYwgGepuU
dkAzaap17QfyqRv8EEfzMwCVL4vCUIRj3cDRlD4loKzpVdFprcAGIwQgQ8mKVeGe8GvgMPQz7aSc
c/+avmczCyL80ngIdedBEKlKEBeHvdOHgofr5Td/VA5SgFiwdM9Qsi3xVEsItjgv9U0BGYyTioNg
yu/jPO8LwTsg8ahimKBUOWdM1rMkBZQWFv6epoSGeKcNfPLlkAZN13WtIsmWj0FthH8UX+6pFneu
NvFp194gz7/SLL77maFuG568jLEXfsXBjLB5wcB5etzQ33fJaEpwzmWZV/MPhrjlAIWSiz0Tn0j4
0pSjntZ0DSApjD5uIUnWgnRhgckTTPsZG6PlgwGERZROILXyJkM7ik1Do5hLrl+sn5ZRQgls0sz0
EFQK1Vw9LpQgCxxAMfQ9WRP3pluMFl/EwVJpid0Tzm/LYdfMTmxsVFNDIRn39RYZF3BiaJAwXa8b
Y5V8MysW3HiKy6qFpWpSNTehY/T1P4Ujk1xvGg2gDBfkAelrLwJ25gsRwwFmtoqhqyyTx3rgEIoY
JiRN60+JusjVhKS75L/4D41Sz2souZ+GpVcdNaYjmlpKPhr+pw9LOsxK4uHWbzXGxu+3TwFMkiie
9RgNNtEXJpi3vanoIkPxEhyr4kgbNVVA5qEuvquXLgu0ynQ8ukXQ37jXyqefxvih3ZVjTTsYZQbA
vuK1xCC2l4dHyKqV96PNPqRsg4obgbCvIQykEBCD3m0PHGNiutXp/GFqnS/F1dm9Eg1gS/YVHKDb
Dzxd/0bK8hNbZnjlmvF+JdDx44FY6U+RX1cEDpSpuExVXxIDQ+cef/c04gaJy9xvgGhoCDSUjHHP
jp0V3Km55x9OS+qaoOSxKKecd8aTAbhHeNzFtvRcKC34zz/oj+DG7ZzOAyJuF48pfq21eeIpiZnC
MB7b0GSfJBBiDLHVzGJCiljg4vabiF24N9exKYJzsRFD5YmhOx+wqH9rPkrV1XUeUW4AzgI87UoZ
W7xuCyFIiBsnLJCFoLR7oZlYRzdav7WUSeGI4HTK/d1Mb/D3N8O6Mdgq2DK4O4thQIvlkcmjY/Qu
Ez8JQDSHSAKLKaWnWTHgnj49KkUjub0MzxwqR0J74z9/2bfUtRtvGv2qhKbw4SAtwPlltikEtzzr
D/m/yt/EPdlRmomGltCuOsnj/kK6qXay3a8ePQK0S+D2Rx8BomDcZ4R6khf1v+Za4Wz/EmS7HjLH
WAjiveCvMsguOk5WPU+Gpsz6VMq+dovDza99q8TURsBi0UMKjnoIJIhk5C5Lv0SREqBEiDhB8bd+
5aRp99fu/SfC6ipDDxqtx9crDqryWX+a4+xPV4k0n2LN9lArip5/RDF3t0cPfpkSkr941sZuOCaO
hw+sK8CxsaUgaubpH1aZZOw+HR5kvsaFcfJYtNSSMVQSNrCdPZlF9SLzYaATmq/EsXYLxNj50nW6
GeZYQvmWY7F3dICChfAxm63BVoQ6bvc+xTMiVlpDKhP8/vduDUW/7qTeinY5GmnsWMI2S8V+2YGC
iC0ipSIIZLpX7C6Fg6JB26vvM690LvJ0/PhUxZXq0/WDzBCESoyy5ChcaAQDChE7vaES7QVTs5ET
jQYTGQG9BMviaCwzUm8dyouPjN1v4V0gWrlcmk7+zLKKBe+uit0g70Ta+OlqVvQpWLTuIzjuYB4O
WlIU2j8vb84SbLinJ4fwxqyS4o6DpV9evUmjI5vxQ+dqkUEhkDoEKyNnijgh7HTuk7z768OSL/U6
Rj69KZFG//0az+pEkTDRUsD7KwbVQSZ2UUVOnNVYXmK+HaDAVISG4pz7TeVXVxfmJxxrHZ8ta1uM
IwgxqwqfD/R/DbX43WBRI2hHLQpAajQefsGC0wzbhkXWFhIxkLAlf6Vdi79s9CnYqJBuj1jcmhlf
BxjfA9cj/20Nll8SM6Ove6liS4aLq/t2lbpVQXz1K5z0Tbg9zhjWgQFxd6jRxFdqMY8WmCN1jkM5
HG1U+nz6T/kT1WnX+69xgH74nzZaM4lDJKgpAezJJLhzOdS6QByu2aeabqKCUyrXAkP13ITnpKbn
XDBg6rrUjnedhospdbrGQGdXnIs9g7CLkSOdOYILEXevd+H0YYDs+oSiO4k73QP9LtftNwbKNzRL
8SArQXeqqP0cj4/Cly3FMF/jYd4VTypeIFm4pzdlvqFTacZ7LhZ8wxuYQ/S6mUVyRwQFg5LX0BAM
SmEGu+PYEY/7oZvZR6/0OdVXKPF+QEpmDRV2bh1VOkOAi9Ene5RP7ED+OQMHONVl13QDv6a4kBNN
Zi0talv+LrXpJA6q1RlzMw4ETDsMjEsRMnYmpy4akfVwSXXm3Q0d3cAPNzgc3Djg5GwD+7+m6hTC
s1uPBHiW6ieYrmLB7cgSq8zng9V1NSPTb60gAPPGibig5DVH/Y5fBxG3mp+vgMbN4DXSveZ8fc8I
x7SgQ2tOWc6Sx71rMcxm7Z8fifXKRVK9M1IYjQ/CUQJvZcYReDBlq7y3+HY5LyH9a6dp0KTnUJOn
K1mtXAxe+Q4VZ5ySdofPKHKae0tcWxcabaiOaM15v3MzAfVUR/Fwy4oXJebkZEPJoscmEaZgxQ0Q
KhGR1smKofB5A/pXehVUYNCDZuC8rsGzL/AlzRwSrnEjukkUbrXsZJq6Hh22yDfa/QfEB3guWIZf
n2Kh1pq80oXMxEdA6Oehv1rWrt3WaVN2qidOk3Qvjdy1QFWcbYHjQEKxySBC6wq+i+VkN1CJm5YX
k155pbHiwhcmrNTfNeex/dhTaJTucQuJkyzMiRvMGTU0E62IictMIn8wlP3w/jNBpKuRRP5VJAs7
j0aNeke5JSLunvHfnX2AXNJ32KRRRnNrgII0447u9xJL7epvYFBgLpPhElqlcEOX4QMFZKJn7CV6
GPrMuG37I+Q/yg5u59I9+nXme3oXuJdyoKytc42TRSir7XpVJF/daJewczWwRLy9DnHdwufl6M4K
VtpTvkR20j8UjHSvPgwg92wqT2LeTaJS4ffNwcL5suzGFuYiA6ngO7ySO3DFFav3DyutSZi7mk9i
KLXPW9EWdLVosQKGkk3YItiBgohvbmnjo1y4syZDQX/Bi5Ux8lE/BfVL44ns78QEXK0V/l5roBfw
53JJZnGZ1hEayFkwnhN/AFHYRwHZe0YxNhby3UlXpGAFh1M/dJYz9mksSVkvUa7Ip+SdA7kSVfR6
D5YO59qDa0JXoyJtEChrfFLmDdcgQuapc18HaDD1vnhrf9fXws8KTNpdtjaGveNY3dT2aKaKm33f
zNetoB3U7L+6TS3MaDiseJE2IZVygk6i6p8D8d/7GDcREfx8mdESU0KalUYPNrP+ktc8gh6H8rTw
LPazqnCIOtRJEJs46S+61nsPPXr7pCmudR3D1rfAxgKBgiiUr+yJdISGCuol4Kt8etevAT5knypq
HBBYESniOieZOxVFPzFptnyDK6uKSjrsOQzwuXfwqKcKZHzLB6/Xtg7fdzn3q4watx2TFUo6ip96
9o2UJK5AAx8Ifjw0XGNgqMP+4Hn9iKBWlcG88poDrxxFwKNMVfewngEDkNKPqyO0TrC5NvfwOkv8
BFXMhjfyED65aIMNPayp5mKKup8vF8gVWGZbdcHjVB9nreY87tVO/BKeHp6tBas/tSO2rPW682A+
fkL7QAatu0seoZKWmWio/HM/0ksPoawt/zLdAIHFpHrnrWZNgAC98PCaEWqpZjTdw2fYtIlmT375
qgB9jE/SFmxgtKJF/antjTYZZXRCBsIKUbVWvLfuK0xtqGb7up6dBAApgNU+Oun9Iu3IQhKSfp22
EeMnVXWslX8irLpHLFOQnFUPGvAbsv0QhrjzlzF/SjC14HkOq1wsSTuN5RoBAd6rNri/7DQ3OaRH
F86t0KuH+kzBUtMO5xZ8OKf5hjnbLCJ9DwPQ9U434cB4z+2UcllTQh+i4iBkkxL/hOqpFzZcihvj
umDVkt/x1WFbQCiK0T1jielxK2bwvEy+Hv9fdd/zj3wQfO+jXTcprwfw2G8XazCg/MrKaMpt3b4L
DY16MJApFMOtvn0LyzRveRn3N3VK+XyYaOLKRVVqc3Xzb2YyebPpoIuF8qwnu+Rf9dYx3klOvX6I
VD4ayyUzQ2WR7F3gb98yUNY5F/lf9jD17S+Z231O8mZ0wnPg39Q7OAb0Awl50tc9DcCrN+b0jeZR
hfI3z5vsf7Eew4g+PXiycFoXwjo+UXl7xS2CsS+bJm95looWSnykHi4qJ3t3+E5G+PiFcx855gFe
ZynuJq99O+iaTGy5YbmnJaj+jrOBkMt6hXtZSLWy2kQDo3R9YVzobwhACQt9pb/olYAZSSo8PWF+
9nLvaKzxD8Wh2G+iHn7VvRaV3vmeOOxdblmd7Ieml5/pbdLyu8j7axdJJPKgez4JKbMdn4LStE+N
G9Rm2UHvYBiK1kZg9RkVWJef/ps8Tbq155EVtF+ry9wIVM+XFV0x4oidxzKwM96ujBvhku4X3/N1
WLBKKT1Duevx4V1iejtd5D3EMPFKeH0cWLjliQNz0I9KIm9kiT0Ns9Z/tVvd+DZFs8Q/PpJCabnV
kzSR0i6JYYt+WSf0l0TWfs5zAF67JvHoj/V3Qluc+QXasC/t4o8BS5f4IQy6CgHxfGelBaWSUZhZ
EJErg9mRdjwVqJn6/mFO6enKWveFIPDE11nnI6PgtHssAfySNT+z4J+7RY0pPUtIcwjByyUEYz1C
UW3eDCZsFCAaXKnYlKA/3pffa0LZKuasDT0q4akvAyxq472QyAubCwU1PMAQgAYlpS71HcUpgRqe
4zLGKOfg23U6cFelJPp7Q3WIwV4UBSUGcyT7od1ljhbWZrXNFCsWoFZzs8CoTPcZ+3e93Ry5zxp4
sI7f9S20wQZzmIv4vVrGbNCPuuqlGBdvsDZeM9wk7JZBD4rrnerFDiumZIUhk4Q+BmvpdOZU95GG
3wfCrH06FgecV7Ujz+sASSSfQhWFGlRUheZCODe53Nq3VEUJEN3p32RtgFsqMYQucla4/l8Y/R2w
5MW1jh2OtscVW6c8+rLkqlY/qCrwSmBuP1CCbzHMnmxCq9Jl5J+NKxmil+uFPktJFQvKLRXxN/yj
GoN/7x2d/glhck74uUTdqYoIGTw/2eiT8OUocKvJFn2941K0QCjOA0J/eQGy51ogv6QNJjz5efZV
L7e92AZ2j/UTIV0l0MEFsncFI6vYb+/CTZ4Hg+KxsWSlJ166hHh+MX8qVcFIEVdNrN3L+thogJv4
EpftWGwNcOnlfz3BmGd4eXhF4tPlcrrD4HhaWmVwsiLQQLBhTxDk+/xAI4jSGAW48OCPGRsmggjP
rttOi/DOhTv845KJKRtM0UIa+AZE7UcHrtt9cG446AB6J7XRW1H7mQp4LGHfdYyJoMM2sqX67bve
xlz1eI1iLI9pwBJ8xFkVbrCh1tPQfcRGRy6tg5w/1lr2sfAqnCMzjXtxoOR0UgPFAe6ZFisaczaL
iljGHvUH7ze6n/qQ+d/sD1+qKzQBEfuzdIeispbJ4pBMwNPh0Guc5npudvxZyjWq0KcN/zXrF92k
6D2PyorRbSGsbFq8vMaRQNNfO92OCXJ7BL04H1U0jq495ZliEq5FFeb8WDrG1YNLMm99INYAKvPO
cL0Z71bO555jvRuQR7xnDTuzsRM4PfZPdzPACvG9SH5rdlP7YATvPg7ubevrw06KPsHfMgUkt1CS
chKM6uYD4TYpnNtflsAlzLtQB55kmbsAJ+m7SM0oys29o0+l9GGctAVAK6Bsd+XKx6l1Gr/oRt0U
idQhRp1NMMpONZGKa3flRHesIa7XAlb42n9TXwn2aX6AJFx2J55h0AG2RJcARVS5VADlWP189Wv8
w/Yzr+b0Dzk1Hf7FcBhnyQw2cr9bm+VD2sEgHaSEmvBLKjBzHv2oYVkW6F/Kz6JvoOADUA+zsCMZ
bJrmM113+E7HJRpH1nfXgAMvIRLZ8vWl1grzYqfKC7+Cs/oCHNwvZjdLd9mbuV5EDQThaFqn/NCw
9Zwnb6QbT6k7wbqzT9LxZAS2mubpsCXdXB4ing0cRM7BP1YKteWEbilu0vGhB9GVDyA/yw9pVTXO
xanVQq7GPRT8CAcNxCBNS+2LqtRCKbVCKa/1I+ScNGxGWAXo/Iwmhn2cx7hQYrQffVzzggl88DAl
8bot1eTBArH+O3tChy9Z+Y3JxhHRrfRpkBTgLkvw2Blksfp1i33RU3IE93svzkGCeJW1eNWiNSwz
+jeox7/U+o1dnz2iaBbpKbRN29h8UE+GlnHgtY/DGAMFVEtStkJaT5SyPNpFI4lY9lRcXbVHjfmJ
qaCvecaCl1b3aNi5r4JfrxlwKbz3PQf1zFoH9pvd3jFc+iYHDe10idnLlYWWliTB8syYwGhugiBo
NLIl4D/il3iek8u+5UQ21mO3UE1V+q1aeVPYUy428+YzOk+LuhVq9wxLo+etmCZyBQbK2EWfmmd/
+u4GjPt7kfEI2OGGber6LRRhL2uO+G2j5TLb6pNVKcvNdbLKLUuuEserWoYDI7b0YS4gklMxucIF
D6g5XHzdV4RVpGCHWaZmpIHeSPhd+jhChFzcr5YCEVVZbenQoEU9Jhi4a63uPcav81lT23MVb1i9
B/dg+2UynVlTQIDqiU/iRSsQCOFDC1EPiZYk1ocHjHo4Q+iusFJPlk1N5oCI7kcJAEuYdcuUqPPQ
pVWMDWerkISL+LKe+gQ+HwkAEfRVM2u/IfIsuPxzRgW4ko508IAGl4Qe6naqsb22DtSkQlaJ3uHu
6v5g2NMCLJsCm3rUMldrRxCwULeljhLt7Kc31BxTg1tafIcuQAxN9qML8RdV4zE/DeR2LB7jBF7J
It6BuFeTQbMTp7AmKnUCzP027zn2am2/8gWLrC12zRH9/41lSc/gMVPPrwDEJ2mQ1E7pc/22XoXi
J21jc49delLD1K4YRXMFgqwG0QA6yufCKzaiRSg0p6ia5uwudmq+LIqnrUZ4jGWlffpOJTEOgdPV
aMCSi6nc3tfEWA3DmewZvv3UmfGk00IBssz1YRQzI5CYkb7H/jqCiE4AvQ6WyAMxnl/XOs7abrzZ
uKYgClJLcNFDXfXp9mA7UTqgE1U6yCiaStDg5CPxah9/IVVKIQyLKVKzqwPlv1X8lhHt6qu/GZ6S
u8bz/k/DK7+0yxEijpUhBT+NvFIPOwq6BqTDC0bFKPw+eQwKZ9lLtuGnGEewZpXCWPJSwiaB1MHs
rCsU+Woz52yYPFtdU7GBLR2IhS48fVpj3qAMOvRLnBwbf3COQ4zmSmo2q6iVUwdGSOeA1qVmzlkG
MrG762BarsSpiLXhZ3UhwRIMnpSJYeRYWtTneCYMcsqxjoKCPHHFxmNNaMnDDGlIiKH2ll5JoHYP
Y0d+sQG89WnkbrHnPmejWkYbxsJCy5SzEHko+NYHfmFZexqGiPWMRxKKjJlbd4f9Cq2dZQhMei5i
4iDquYhGoGAKCbulJbmlIp0FjGfrsHA1QBo3oI5VqY+QV3VGMVgE7/x/cF4aAVf54uR3fI5GRvfw
lgc9IstEDrND5JOw+rqmNhI+v4rulogCwqhUE6FP9eAfCz50U503m0jIAZIhz3L/+1O1BOIvadUN
RXJlCZfkiuxqlODxOTve+s53j8JT4bpdL0x6A5ubUxq9p5SC03fQOW1gh+bWBWKLT5m12pHc93NW
46K7aJmbEZw2I9zupKKZpatSLiJzNdTf6ii+2WPprA0V1zYw0UoHLgmWo6Dqnx3YFWqQOTiL6btG
tpeQobnHLd2ZL1HO56dTxFBX71hS4I5e6voSCST/nw/FhXTqi2i3sy8vnEm64PdC560G0W9eUhyY
0B5a2uzU8ntYlUjrZmHUpQJ1Wu43E8FpKXoBgvisOW/rmKzbqaPSMPuizYdrzt8++RwhwARGIwAR
Bz9GJ/gjpvG++p3BnbFzcW060ulL6o90SQztGQfSEtQlhYcxFgrMx1A3goEZisNdOie4AtH4qqXI
CP0PRlRW4/Sc8I6ZyTdguSwOzPHm8rRIQBnAx1FOT8+utsa6Nx9pbY5cBAgR3o5CGwohEdhe8Cer
O7zdLY7hng9dhXPR+rG4prHc+0SaStGhDAzxgeVLIv/M1gual1ZG1SuU9q6++iH44imYDTDqUjVW
+3rXttP+Z/U6uSCbHDELn6gOkxZ/kSKAtqxri8XGsJmCe8j24FQh/wICSV5oiC4hZnfCAYmeodXz
J3iERvzXp4USRl8BrSok4WRyAId6MBcZ56P/w7HNhnK6YW9EEVBxTwAaV1U1tCCdK69BNEc6lWLM
sq0AKYZT5ci9L3Szj3e1iPruXEhGrwdXGxrnLJx4WF6e3GRKQYoygv3XdtfesONeh6lkeyX4spv1
WqBLbLCdXdcg6ZNplVQH4CAKevBoCJUwd9rb//4X4XlFgHsX1kHnFQxMYpeleO/5Fv2a9E6DacfG
2zG0RRsyi11pFKF6kFrzQm8oJPZOhut1+YyOpY9CtLs/hA5VTLckUlLEKNP2khUIaihVKmNc+R/T
UsAeBWFFoDXbrXuJal8Q0eTLTZlhL8jiNbcxxLmu1tDk0YDt98OrFq6FEKsVzikse9HNmuu9TgJb
20UtUrD5MXsd2y6RzuVzqHcXtMGXkcmLjOQg94a2bkuySU9Opi0O3bQlAaSjEQYLR5o1zszJbw+X
IxjnNnitoxFr8gLO4DJv4JnytEt7c9cGEI/R5ph/yz6MIls+f3D0dCdTH0nml3yvY4MeV/EgGTZ/
M3ZQFGOJ4rP5laX+KW2HU4hpONiVXVvKo16VeUTlkSwtkcuYKKuWkBxBsIYA0dbidVbbLWMFJk5+
lYeYzHG8L8ztH8Ri4pJHcUy0cUMFkzRvyRGHFGerVPsEOHr0Y5fA4SaPt7OBz9g7CN4mMM1b+MGN
sroQMFzwKVzl18eWqI3Zk4zm2/EY8Xqb0IuKRtbOXjMcSofn0hMTum0CeVCqSLFIjiP9HuLjFLC7
shPXvVkcDUYanG3bkvU4iphIe9JJJXfEu0iIu8fYUX7lEpv4do/EAs62WRBPP2M85yA+mjVXKpmM
B3GuGIw+sGHy1hzocFDCgPkcf/6NtmKZoPcCmVPkE7sf01pZOSiCB2tfmAR/AN1Q9AF4Y43b5SOu
MCbIgpew03tB3JT8SPXxn2Q9AIa7cWz7a1trEIUuBl+rRplmOKiISrfVv7fYu/+QEg2nAAry5Gop
JxZvFunwPjS7NRrQSjR0F6ocHJXLXmmj9gJQ9QFK19tJZo87BKRkTAfBc/Y4Wqv8eDVqri9W5DUW
lsYWVvaitVPCrhVQpLvUy23LTcg19jmdNA1vTQO95vgF1KMqtWtTQX5SYv5ovCzkBkuX8+MaHCML
WLnXzzm+E2DcOaP0rCZ41deUSD1U3Usv8Zjywx3Jk6aHg6q3Okw1t+fgcjQixHDLVc8BAm1Xj/IH
CRd3e+ibDOCvdN04hTMLFuxQJPo4aa7GLUngI+twj6zhCmsGCi52K8P2zlysx/GkRXqoA9gjItko
+u5W4mahU5jzKTlnfPB+gtIGzGCH6m4TApNiDfJigkX6ILmXMIHRJcJC1GD9Cye3zFbRQ3aceFho
XfuP2jRbNO2W/6zFg5xAUxHa8SwVCk5e3RhFVlKb4z7e5SqrBOmbNs0RTMzJa7OPIxWE/UkClgxm
9y03+k5svSBKVNyCafjxd863EZyXKNTnlHbRu6C2lOJ4WKA9yibFBMKKJr2+i1+4s1jx57Dpjq/Y
0MbsZuHQQlRGzDZFNqi3zUqhDXaLlftYS+zDPMuBYycSso0VhoY1WgdNBtqGBL9hesTjarpPwqHe
thSugNMHF0LRHHKWfu5fmrCrkLAa6Upr/AcUbYFbWtPqtZzwljeRp5cONzXdPoa3g3Mckwa+tTMp
UNbOepGZgL46+WdUEhnLrYRW/U1YXs3h+/uXW23ysXwCjmk5OJpHKXdr0CMkvuRG1BFkfyPjbryW
mPUFMe7qC185+3CPVi7Q4RTPJHMW2NUEH1NyDbeTjZWI6EgEm4k2kIIHa7GSZdxcTB6GrL+8Q7hX
ZZfyxRy+/IobfP2E9ERh4CHHfsDrVMo0impDa+KxdVDn+LbeY63LrJWF2J0H3JgwSaYKcW7Ur6Q1
NBgEVsw1kKEF+l19lYpJSJp4OAqiAYEo2dC9OWa3PTqNE345eSVhQxJbCI/oiDWObj6uUyrYuukW
R3UmRsR+HRUrv6Sok3idv7dup96BiF/6YKHlsRlnBqyh6n/FIcGlZLlS9J0LVkBdhfXavjUtuTF4
dOzkrYl8O7SGGNstPmoY2zjej6OP8Gsfm9/bbu9W+FjSTzNlH95KExdVICMm/cBjfGpiBemRDSLE
DlNVp5pNLa/W36eu2HxEQfGVAbBqQAghuMJO87PgOaoN0TCsEGcR8ZTqxTJSXKf4EuT53/vl24YP
9kILXdQePGxzp0UXVuPbvR3xaXahfjl4mSoCR2wa/P8i7IQMGqs1oP5W2mRqgvH4NYJTAGk1mR0y
28YAIGM4HuGqwHpkOfBHwnklIGfMW+iF41RuPowup9Q0+dd0hz6vjw5f/DwODtVf0SMAMWbSW7h2
erLK5V/51YIvyhFhTsKcQhmZOo/6fxtNsxKR6jCU1XvineTvxyUlHEOgRR/7jc1p463wRWBZXCBj
PmjKTbIrfFYRgpFZtGY18GrFHoh68BVbogkzvEqzkuVQ8ErTSTZuNk9DJDHYrDW76tViXspuQskp
Q5Uz237RzJE0xfe3mw+lrAD6762vaOtPimVBXiFczDaSpCxkzg6sKLEbzytel5QoPMl0uV5MNyZp
QUTXRHBOPgLCPR/xWojCveH0hn17EuNGBm1wIO4TvZKONdLKk98dO/tKfe0Ywvqf4gBcPh6Z6fW1
5DeS5mcAolV0rZ3NE4X0wbiWP8o77tH5YmPziTHb2U09BkIG0zYvsRXAWCwt5X2scas5Qg/DN0Vt
5RQxATQZiL8qUkNCdP2tEyIrF3DDlA83Ud5NRnUSSvOc6u2CBCmU3m+JX4CxQWNi6cgpZ7SZLN0N
dC8Ia30R4sgKHpxmzfmUapYeqcNVzM+LkvFPzHAhsi4JNi2NRaPwBKz/HhJG3cDFwt/56kzaWYnG
P7gzwd0qbCMLi7sx8HoKXyIAYo+XY1uKlxLsgnu/DklTXhyoco990FbZ4JVmpyL8GuH0Sx4kfejI
V7lQU+mjjfzBF+05ggfdMtP6zpcE1eO7fEpQg51X6VgULxHuvhcR2rkuP2v8uvtWgYUlWftblOJ2
xn2upMMT5TGEoYw9Sx7/Zs/IMnIpr/e9Y/n2uMnQB+oam7CdvyQoWAvfN3j/TIU6Jx/2brFoU8mH
kI52kE472p9MZ/tL0D9Fmksm66pX13hrB8BU0vwDnbV3i13T7mvm8O11dV6kXOlVNxPCAqNXiZsQ
3Dn3S81hQeHmcNgytUmicn7YNu0379CLaOPQ4rOBbXzHirzT/Y62NkIugWQRArIOMpevH4F+Lm/z
lRjv32CSF/VR299V7+Sdw9ZaCQdodkKllvlMwR4wGPatycOIDK4iwyvxB2s4sOVMGl92mh1Mkfjd
KqihzDlCbp2lzPHZVMypm5zyhuo3DD697l6fk7edPGhmHt3DRYcgcyyONYBPiH6Eb5w3ZUICa8J4
tS0Bs40WEeRiVHrK/cj/5PdOWebD4dkrWYLg3cMcWi3qAGdNMbMJqfk/HJj12nzVJKJjK1K5usBT
t8wzYdxKzIBZ0V4Ok/MqRLa8k1hNXoTYWtEdQtcv2KpcgeouasBOcaQ3i6lWzGZzSBHYD0dL4E7s
u/41fufQq4xoOiwX8c3+ecOMbxWU7rOvcGoQGQWCYkQnuSYnarM10rebkk/GW0rQ8KKoGbOF7qqJ
QLiuI6B+ewc0wwKBx/JgOq/2Dort3XJ/oEf4zadu6H/Atv3YT/4WM95jN3ey7qu51JtqI0/LLk2z
0GArpN1L+OB6X5g/yfIjpgd4dWep0NOa5WtSb/Hk8bd6cP5h68omuhlNtHEroHsM8A7JwrT3hjxB
OOm67c0R3vuuqRt2i85MdsdZ25jyEzw1gWQOU4WOhcnUowCfK6RgKM51WKVUeZ8Job2tcgZHZyGn
R1+BDd9jS7IXL1by9eKXBeVhSljLeXB+abbDMRtrDZBifMYZf5X5+n6mabzhbb1iOSy4iMd49Wj7
8YRqmb2RW484Age1H55OglKG2gM+1SUqybsj9O4WHCAtNoBoyhXPS+/lMePiLA3hN2bHBLD/GG7w
PmxD7R0Cs43SgaNeKkEVORxH9ZW1T/GapXfjjroFZ9/fRcLKdf46o3GisYBXdXscpD/uyYUPvLF3
AyHdHjUaQCq/Q4X8uQOqQXbwgouNT1XVQ6I+r5B0Nh+8ORC2oMW1w+eRwJ2WZlTyan8zFu3Hfu1V
IVP7oAB+kQi/uCUm8PnPfj1PTs9sRnNaDwFcQjvUMRulIkAZFy2FNNGgrX39F5+3Kd61Fz7OGHzG
LuBksS6de2Lo5oa0XZfHzxw/y3VsKyGqXNaWgPoseB36rasYyA1ZbwBREXr1nVBSvJsoiE2jkc/2
FUhN6iNHrZbdmlv1TTONNaE16Sm3XFYoRPCS9V4qsCX3qSCPg8pVCR25bDgZ2uC2AGrNwrQv+psY
CfC35rmEGcropsD3jnEaH+IuuaHI24Ub5s58Avkt9T1DJvCsKsFC0w2Dg4r+gakjOGt+xQZpRt9A
OfE6qocAz+zh+j64gLA6WYUnCif3Kpj6WZ9pwsfLdjlHeR86qZPKPJLw4ivXH6fW1fPLk341tWkp
eTOnDsOJMiPYVVPqh4Zx1K+EvSCJXxDl2IlX+aJJHSE2dKT7+aM9I4IToPnMP7aLp8t2o6Wlbpe2
VBdGVTA8dDCq+4GeGQ2n5RkS/e9OspSRddMg7GF62n3C+ikAFB3A2DNlivSkASDbYu1eiDiHzFIG
0ghSxzkYTDSV+BRl7r6nJNFn2VVZNyv7WcM95V04IHBkPiVDQ66qan8RQ+Diy7Mj8YcAmV6TogIT
9FF3+8JKres0HKRb2kGX3pWQyeXpw9txyb03J6wGkDpACM8KR3vTe3bWlQ3YKf7fhwZqaWbQZNWj
Vkr54jIYIlW1qAH/LabfT01iP1KYY5Fh1yN5fvWd2V40zuQ76ETL+YD9o4MSXViTLkZqIY9MlGjQ
Kb42ydS1TgcubJA8QLkZCDM1nideFnEUws32Oo4D6/bPWMtTObAs4TR1sJTi8XjaZ/wUx5DwR6wn
WVzIY7+xYWTtS5tJ9opG/I7skcZSkwDLx2TlVQDKJgYE3Dft6dIOQyGghYAWqjJ7PmYc4JMRUz9A
LbuVvooGvi6TIYMySygC3Z4McTCgIvmH0g73efMDsLoWpQlGB0zxzp3oAcPiGxoLlCJSWV/Shv4y
3inpmiijl3iBm7yniW7aw41LnjiXcPxV7Mq0sDOvi995BLpi+kJ4lSIxOCRoQvr3IuXG5FvTsw04
e1iS01mPDTndxQ1TaHzo/PehVaO4IePDegIL59OZmNynedPPeGjlrRmD+IBQBDCNCp2LKPbyfFre
aLrtf1YVapKHzUGumdd45DY/kPkfAxo6cktyOX0sVRkV7PjJ/FGedy/K2EaK9tx3W4zYMf01LfEK
wxHqrDB7EAZWP3bcZY0JLuhkXI7PtlKH5VM9fv7b37e1kEHqy7UUDGKRRBIPOFRfeS1Jafj3dhRG
elCC21Yh6AQTIi1p52xW0LMMFCBku6QR3kyGyNDclPZ0Ryio5bkzPDsoYeh/ZDrFdUcC+C+Dh9y5
ziwI0aSYd24BWWhIkxVJ4lcvqmErSH4m+tBNmi6u+TrqWVCUQlGZgJaoGheMYuhm6B07fcCVdYH9
4h6rVzHiyHIs57GdEpC5mcBoWWlDNDjxfrH5Y+f+wjmnk7qaFeOhkNluorkmJulzNBfY8byzQA7c
ww2Q/sNdy+DUlzNb1+olqs4PwraPYwrt3a5If326qcrc09F4YfXUrNv4njDFUe7B64QNMUfED/uz
nFmGgd0gWdNoQv/zI/MziSGnS8Ax6EHZIF3wlEJyfejm1K00XdJQAW/3yJO/U6Rs8iKH3e11Fvds
OnWadSQHayJfvNlxK4JV4V4DowcENJO9i4QvMy6pNKju6X5xOMFYDYKKPSXFQXwsnbwDFDPJocRi
zJvgvbk2FN3bSb6R0HymK7N5ZpTi+cUeebVwiULWb06sZXM/QygnvnjZ1GFH6d6DojduZySnK1tv
AigVRPTr19g09ZlKSnn28g3nbOL/VG7y8tWk22oCNO4pWRs8czr8Jfnc0bEStzDr88x68Dx6b8Gi
DCaNN9jMaRkvQxze27aFkFok/CVd1qruIE5nVD1Rd6stOIYdSXBgrNmA0XfM95SaVIHqqusJ1fM1
DywSsMCroOixj/hldaABIx3R5WJAWtpav2X21NrITw5KDE4j/01U8cQ0hST+Lo1ckRpg7VPsJtOp
uNjaklX2kLg7VjfC5Cv835I2hoPGIhNg4Nd4iwNaiNnRC2PvwL9PMsjiCOHKM/I9/s4iy/KbuiFT
e4U904ETrHNS081NzL6IXAai7XurHclugIdHlAK8Tkm7nq86tjPni8YuRKk+S29grpGH7ioc+cmp
FfOu0o24GrSNrkenaesuMlZF7yca0AWtXYhKkx3jYgGhpOK+sEUian+bd6kD4BaVUBbFwVMqXKbL
4uJrEpWCcEKFYwjCIg3npXgeEfPrxfM56dM2AJ7h+jHtOs8NaahthlHOExaUxVeUu6KD8qtz36Sa
jlBHGYTs2Ry4F3rGUd82wT8iKgH0uz8ZLkUsEGyteXtBhWuQrSFxqvBqTYLFkWxUr5xLryEi3oql
DY3gtodTo2/wdEBig1GRr7w6KpfuIRaBR31GeQhkRf+ULGl/diCiqlwJSwtdqZ2n5NBtyy1fI5lS
9tXuSVT216zuvKDrlWRaTrL+ZdgBDtGtjKheY7FiweDw2pV4xuTSCAfDpet8UPajH6f95UrL5ZI5
tMkSQ6AUt+w4G6wetsOVK7hXiMqnO3WSk2kd8VQWOq+4AH8ZkPNbqCj+yX/tArrODmjCU4TUy7YX
ZBumW5E909txHp0O64cgoGiOpJTtpqt4taJMYPWqONh3YRidhTQGYZfZuCcdcD3FvJCls/QRqUOB
aLabFADe9XvlweELTUncNw2KX4SceIHiLYqzlBCHBvK5ONneeDqOqv21nH/JGBeoH0EF3hD+BxpE
7WRuxCceqZCwQU8K9lFxEj8HUl5PPJhqR/7ixMk422+CYnA+hjkrqooNEJ7xR23jD4HvfRd3/UP5
PFMlfI+8inopPFujVP3BlPJvvrs0cpt/ZT7kmQDiu0hn0fXYEsx69kPnMD8bY1PIwqnXjbm+HNax
kAfAOgvQoKnkXkAJerYGTEEaEpz7lsBCntdbROvPaNFFcdtFgOgqIIs1/nv8pRJqb6zCPauQVLIa
LN/aoI9xmHoM3+JvryF2/ll1fxfUsR61G1psPPWJtGWgfBaYjuo+ofdINo6OZlLYvAzou7IylWbd
QG3+jEwJP0xwenL+2nc/6vR7myXzrpHQajGFUOJa/8PlHWZPdSEDQMOPpMHgcnUJP8dqFjITbrn0
vruSD2Pjg7WWYPcRi9Lik48DwrIKTsAxGteOYAqUzuE6EaOglKwzp05mWTKSWm9XWuP1HhPfMrG+
vJaMPY1/5rBvykj+DKK9LuPr8ew/0wjfhGMo6+74VsEfdyhQpzOVSnE9NX6BYWh6VcS/6AyYEbWZ
xynQTHD2YWzWGl5Mhx4Sq3tY+TzYmvIQ2B2HqvxoD1jtfUlkHXdEqF/53J4FpT0q3qPtnXjO76lf
QCfvELkMX9Uiqrux76sIDfPtmjFO5bTZG/A7XgZol9H9NngU40jvGvDUbKQ5YjpW4QoibuHIvTMb
Dm/CauAKgZI+8UgEpxifpSEmnoJch+fF8XWVC4b4gMyPCJiAGi0ZI3XvHeeI6hH+JO1pSAJOGTDL
zGkXLT/yZ2l1sfWFVhC2yHQuDoaCQTRzDqXjfG7GmnTWd+2liCovZPjOVQGNnrNiuypOfXKAOofX
o+w8ApFZikDBJjKI9XEm+0QfmvXXrMlOTAizhA3j0BhpDKWvv1HO62mVgbn5GF/+JBA+o4zEIt2H
W2FfIVNXa5wQeHCjb5cZMnn4tEhbNfHl9xKbtvb2zrCQ3wavDclTYbwcHQRVhNdjAnZf/sdjKeLT
Vl3SuE4GeYul8+ODTdnOnJZNJW0AZGLhYrnSuZYmFIYMnSglTIQkg9dnqcjM1QQxtXVPHESYF21v
I6DjqBj/Bk8HjIULNEEuZPhLBKy4+/5Za+rgkK2P4S3E9JqTNU+jSV9zyEvt4Z+it8EVssdVKluV
ha9pnfy9epiyIx4Hbf6hC2zrUcz/WzmivERt3SZHEgTMC6K7xlspkWPHlAZAkTnI2rmELGRpv3Z/
I6buXQJfb6w3ev3blM4GzOrNUUirFcjwuxVkJA+YweUiMuXZnSVTnMM+hm8tGw3fcDGNivgj/+pg
RiZQvv28Bs3djDSbXMrnQzr/d3aeCkIhGPlr1fwSjjahbnE9VrPq7nxqSfISbb7otvFbnDWW/379
x/pOPqRAHzVdvuIEzty3Xov4RMOIrDiXNw49t3Se5ojFlIgQh6xqFaeN8+tUn/jVjjg7vCUPxCQA
yMv9nq1WB7Ws0XRK5swjdmUXQE8aCWF8s6t22MItDyPBEbb3NxV0nx1QoXLj7C2FtpMiDX0/0gO/
FGZ08frpOT/s1pr+Z4r+jIN3wcfu4bcOHx9/Zc7SNBxu1wqjjQ80LzJqhnkdmw1NOSjqYL+5Svxg
rnJwoiYx8NwTTTi9pd5ZpWtor+kYXi+sRPYe89W1+2jAGBs7+5Ldl5AlAHyd/0mpM9/R2p+rYOJD
YSMZRd98ZvfM6PtL3DvVSwlfPT1ZMePaZ1w8D6m4A8G07uQDwT2fZ+NuzMEZi41wyPmm3RQTluVT
ex0+XmcuAKDg8SYiisgcEVcMa46/hkbjNC48N0ckhx3KWGlfdvBcRnMSzOZQI2r7xYo/Ut9sorJb
m11WiR9FxVHU4eyPCugnjyJoYZOUzSTTRWr0ho1TqeewsR1jlCNPQoVj8yp/7F+nZRxkB4uizVff
3Bv8BqYwl9rHHb7ldc4DCTkK+lFR16rZSAJP17yGjcuovk9ub10yn6mp0dXIrd0pvT8hIXGXKQIa
ymPYOsQiQIClAF6wh4EqGhv8bQoqE1w8Pkts5ZoGQQmAZSJteBePNKVboRaP36+zgvWielo9j1B0
kUDNPi4oZCfrv7wzxjBH4M7qbyGkJuGs19DyURwD6bFRSOFkVmoB8RJkRMf3pWd1zTe8HBNR6175
sekXFjkfhLM7xonGjXIiSCdfqy5I0CzkYYklpLBYNpZNt59rsN7O20amwCaUMEMv6kFkxrcIP7P9
QNszzUbxx2MZkgZjraGp77o7AHDQczHPgzFZbwLzfUshwdaNU1hpH8c4S68ZUue32vPLAG9yBiWC
ngc2+fse90koNELd0yMs+FfHJZrYwpjnrzMWmT52ZuB3TumYFNq1CsXePou/bF5VPIiNdW2/mylk
4wZ8hGx5bk5v0s1/+nwfvUCuGv4hf9KGStxQT8sbm0jEu5HpHLqsnA/bJG/MEQwO4btDYR5lWeFG
HV8wUwazP8w5YT7lZ9O/i4knMWmu92eJLy69HoC7KBUTxRM6Ou1OCb7Zd4O0eoOJe5bXaB2b0NAB
Eo8kdhy3RU3EQgugboxcnH/oYu+nfSoX1v8d3xXIBTXJRzxLy8rcGU2qQUknhns9fNQICL+KK9ye
HPBFE5aQ1s3Bjb6rvML9HE2DZl7Rx3j5p8v1YghIazu9IcQvsFcHi5DVnaykesJYdgXdBvUw/WSL
OHHLDbqsW9kTtgD79xmw+vueLnfrs5XZ0A9VYUJGTiMD/451snpihmdfFZxEewGsYoLySgIez07p
NzRVSry04gEP7yQy1YG0kD6j82WyZ1DIj9pToX8Zfi7UiNC3ESNWQOlVK7KFo5QluTpZ8T87C5UT
3zVG8909V9bZiF6AKu2HW+ioN4APRkkllE5Ke8QU3lrYrwEdfL6WfGQELOYfNvokEpDCEDwCVlvH
RJ8rHpy/7Ve/e/zNIrWQpH6Gghmk0zWb6Rd0FD0Ruc80SkgCbebILjPZSO4aSuRgXQ9R2fFaia9I
Vw/AWOSFinSgKmkm3UenLWXepLEhFL3AXnMJTbjq8Mss8EAStEE94iAza5Q59Gs5vhCuv/VvZOO0
eXR9qeND/n5Bw+45szTbdLItY91kx3Ep9hUqc5x7lGmCm+zr9WkgNwrLHBbM9O7kCjixwr/oHEtN
lFpVmuyfVUdtq5oGBUaCSrb9n/+drhbdTgAacqcp34B/c8nwEHiwEt02s6HkOVIFWnqFqUlfyzAg
4xlQmGHRPC5NSw67TkDaovxGjwD9nY8Om82QGzjJWdJMABKhaXmWtcc2/oIt3dvFik7kJBLPIvx/
jRXE9ULRkumgOJGQtt5Kb1gVZTYasd2Vkco42DH9pNo/PfAvPXXILftkjePzsEUi1R5qGdgAZcqY
I/KRMDNmItjJqFIRKgikOWV/l5PEDDXQaJiD55vGLsI1IzhuugpawZ96UyKcxbGQ+JgFqapZGX38
j2JP+5rKBVdirGC4itsrMGXUL0nFsR4JN0Ha1U36yi2oSZofhKBKY/yRU5MN/AtCqU5VVuW+GPBB
ObUZSESa9wlbK3je/+Ot6WAknf/kA3fy5TaFZEUEultB/pmG0vS+e9oXszq+4r4+mOHPcj4NZRcL
Vp5Bu2GPcx55vNqnHSoKRaVW1PwCjHQXde2iN69762hN1EyrMZpswAcsybz7tOp5r1UoChw2x7AH
Y0pHJDYE8ziaY0oBDHJO5vUmro/1A8qufQvD90kdjr5u8aCQqVAC6bm+N6I6/XnmBDXI/kXWlPxN
YZZv8heYdjCmD/uAbCBMi+GkpU8MENr1M0HQjFL7Ggaw4nPwPE1CHIqouNEKd22ko5MdaCjoWe+i
Z68TKN7y9wEfltiiU3ujjs6ExSwoq4BjCuyM05x8Pc3dVO/gF7U6ZGaev8D0PN7sba0nvzNQYqo4
yjuB/smg6uPPmsAkcCXCmK0H8oAbOCNET3GaBd1g2hl2BiS4WCjSybaxdaH2CDzVYxcU+tXoOi2m
OxgKj5CUSfLmJwObL7Mm3auWOSo55ng7AahKs52wyHp+A2jjPq1+yPrWPQe0jTa1goikywSxERI1
CcADZ4yMWlfiQRwr9RufQpkBiL4MFuZKQRC0pDycR2cvnBA6Be0A6+ilxTkIc9TprBEOkXRskt42
G9lZljbfmLx/AgXjk8vzICPpzS66RXc78OsZHKbp7vHn8YdzRiYkQAWZQhwg2Y/HtH0649Mw3F7A
JUENlaNGxdvFeC7ZWwGrrzzND8svicvd/xZ+z7wa4PO+pAB1af0p5OZwA8BbJfjtnZV+C47ipkwo
dLZ0E0vfz3fK4rtt4ECUWc1SbLP4xkGEJnTyoLXJBV3iba3nje778sXmlFyZXC3q1/cfYh6lK0Zp
1NCPAC7lpl4rmQE/dIzC2MuOZ9M4kMRCsDA20OXXgMe1L/+ntGBf9DdG3EH/erRGNnevVbNKwt5l
h7jqaOr7saAqfgx3gP2tnsR2Ogropjw8j563zadZo+pXDpjoCt99034IrpQyCYjqKGuVIENuUsfK
xtglq1reeIK1HshWhCofDxWw+9oyD87+nIjwy4bjkyrMtHFA5Ae3wrdwqgrjd4vRA7dwIEBkSHbr
kgcUfoNrjZLD9VTyvLbsuvFoLwSfZ48FoMApNU1IQuPbAGCwzFocaBT6/LAG/TYXHo0CDBs8ei3r
2hWkeDbw6jUoo3uLY1qQ98evilYWws2DKf2qQfTJTL/x2Bq6OyJl9IFd1vihJlh56w8Ky0QM6YDk
1Jq5j1rhN10eeIvl+sgkDftZ4zsdHsJC0vUkRr871mmr3vasjmIRpT+QcWtAvK0IkpqbFSroWfx7
7YlD9oduXi6ll6NkX/o7W/G2uHYfRDIgRbHU9w9XC0crXzzCAd05x+STykyEgFQ1YaGEXwbm/Sls
dDW4QhUq32ZLh8Gcf+cTGqXEIn19QCGxU7n5mhZYO3T1Nt6tTB6t6QoIuMVcuOlwoqBsU3ZpEPB2
mDjI177rAl6jISBKMjxQchYRGRINRiKDRH59zGcTAJyuytGC05H+1YOUUYrNwadf4IgGpmkf49KT
8OSd3vUcGjqAfdW8Djon54uqVXUXYcSJqyPyrHGzaS54redgye+pAszdeKt5geUlIeJsgh7QVumR
MLaohWtWaxPINYlpfHsNDxHkpgrAJp5aa15DhK4Wv28+LxMPxuKds8T4iC4ooMdF5UUeA6CjrNXq
cXesH2retHwSWKKy7/k4XVs5rMlBvgqI6O8InrsDWKd/aSjCzRhTbN1gX2xU5h4BZF9e1Ta+jaTo
45FnkXxCu32SeVP8sNhgoJtq81kB3WATolSDy/EuGUCjHlmvUz36XnGJClniYBkjeG0MFGNNw1OX
o6IKWEIxOcUYfZEp4e4004beB2eweyztW7TOBNX5R7kY7LnMATLlmAIV6ot7pG+s5qreVxTTNpxx
YWIgN+CmOmuv0EImevFuUEaute5nMeSsESiMXlP4StVbCrx/0vjnnDBaCsD6ctDlV8ZtmdHWyq+6
LI+UuP/nzj5BPk1Ej7dK85ljDjandY7mNyWxcKQkP2u1Ts+5HWhiGpWcxtGox4sGDJBdyizq9d/W
WybVh1NYPS5ixisSmeb+P8iUIzyuzY04YWAiJQozj3w/Ly2JZ8BJfzrmgjLHZLt2VwU1FxH7Ied/
dXUM0dhNdP/O27Q4RQl6+yUrBG9jR3272Iz91RSIpkyduDlU74p9iwNNMQyxU73oRnzL3SkT8Xk2
XIwODZjwgXluCy1npqz/L7Xd7NpWBiZQRPy6SwlXQX+Ib+hzDHn4f4eSKQZqdSgb+FYMUmwndgno
ssRqjGBaBd/Uu65zppA3UdWAcVjDjCiEDPMNMt+PAF23SqVtiu+x9hL+xjp7nlF3fBNcaQ3eFUeE
0Rbx5WCRJnxQ/h431HWYkhmkL9ACD52eaY3gIHm99uiuCHCIrPh8L2NwFFyA/3NL2P4k8hpS7lnM
vYQzlFx4EBs+zpXKlfTlmbwHJEFUTV6vMG/gmU3ZUQ80UKw7ASngQbjivXnhUmE2aE+BrbwYg7Lu
oZ+Jj9a8dKDU4T+yV7EGHl3pVIMV/GGi7mvNkmLfLk8zk3LrPgfXU7Lx5aEOjOt17KbHm6mNzgY1
sgV7vFLunRNmHkII9brguIY5Wg0lYJStNwZ0hLMQJpBupHQXso947LHE1QQqi+PLQ19J1qdMGYH5
U8IhpqOMYySxWA1aEE5nVdeV0RJX8bJF8Cedv3OPIQqspkc0pNRfPURGmUkUppFflPnxfpVYXvqe
qkmRGhcfOEaDF+LUiDHcbnM/ghgEA/meOBqxSeI+zIE6RtDwDR09ZFB4PgyDLCu+3q/TiPiy8+/O
F+49XuIVsU68VsCe4Qtv0mzYm4XaEaE2DAIOTWVGZBiL1FRDdj9SOtLmsySvJL/zQL+Z08Av+E5V
yCxCn5niXmpGEOnQDCWBxmAYKq0SS1EXfdtOQOIHn+REDDrdYEB5bmd+W8arXk0xmJt9oFPy2iTg
pKu6YW3LNE5hZQeUMeFgLraDQ6uk8Jjgc6OAoBugS8d0EHuOt2zTh3iGm1hJVLgKwOVkdyho5YFz
zSEOtBLl932rraXlVS2NjLgHoge5N2jA0icspsdGigB4NI36TyvQ5EKF0Vg5rBSwuS9bO2t1hvJh
eSiJcmuLHUI8uOQAAT2lBby9JUxlOWUZVtmWesoyxwp/fIyCV838XHOwxlDyLYt+qmIwWRx6g62O
LqX7htKlFNUvrT86mzVP8Fl1j+n/onLmq+0F8nUM/r6YWyleJIdjq4i+tddHUaAKRO2fNRGp9AT9
w54WKl7/Vq5UHyr1D2tgZZJTASxIdomaePw8oRVv3mE6yf8NTV2Vk+i77lqgX6lQEcZLnoc5ayjq
EAcEEqELUVk7UISfVp6NNU2pwiDCk5fZVMAa+3osg+yyAUmCEXwZ3knIm6JFlMa0NbaOnd2nUHuf
fGhPKrKwJ6LVK/sZO0X6LQb/udqbw4utHQdgLJ/7MgGiO3bZ5ue62w8jBC9Xqfwxfn0UgNDXmGRI
qlt3F98ByJw/a6KmmSbpgrzZzXyX9crreW/1OQlYNp0bgBcpDExA2QGlPVf+Xqd1R0ZnloZPfEkd
VElEYIhIBwJXH9Kzq0dnbdrTnf7klsK5n7tEdJ6roAjdSYxapKlVzAzR8jEHhL4KZwmDy2VPQOGf
tT5nRP4KKNy4K58EIxvsgTi670m5dJ5fjf/J6ayvNBicus8wmFwlZCuJEYHzWyF+aRMBbswWX/3s
Wag0I1F6GWorBqXXclzvL3O2Re3fPuoagNeN0kpwQ6zvUhp+VjrfuTUtaAWcflnJpxElHdeK5PrL
wwsXURwm3BJu+gyXiFxiBMN2Q37uNeDRIcu4NutcvvofLVNNDIP5irXRAhyI0JSvRiFkT14eiIn+
2SxOjKIldbKx3Y73ZLAE3AUwCdjg42ch/WD8UFQPbgj+ybOv92RCI+duwlN93lfCNRG0a2OoTEys
APVwOuTetVnUefEAXS2VFDrv+kJ55iWSIMY/tpViXHAX9XybvJu7TtGUPM8/8saVY/hhuVeF08TU
GJXVP91gE6dwcSlUNmQD9yswzTL2zICfgPNHXZP/gUdz30fCXG2SCil1OmeHoOHXaz9ku2StVI8v
3rzcHpDzR5iUGmpYS7N9I79L2G2XiQ6FWLOqMmhrCJmmzpM10t7CLM6yhXdnTCr6IyvRXUl620Qo
9WJK8G4UEVIbT680xwCWBSKjb3j9oiHxV2JDJwvu90zZLk6I3nfRrrjQoULxK8PSUxWEAniQix5B
Ta8hUxQ2d6fHtKfUt2SwkiEaIOGdLKWvBWYC5eyo8eI86ZnFMc3F63l/Sz2yTq4PX7b59hgWy13I
VfBTyaniuHpDOMch3x4edLufACA0OnNo1oAKdN8GO2AKMMr8Qftu8Ir0A7uWf0h+XbDLySfo7Y0O
8wC1LYEkfkrUusXtyfpz+vgHDgG9EtwsBtZ6XY+iKO1jzLbd/puq30nRtcNECrzbY3bwsDWcngLk
6M9KwASBYXzDwG7mwuGaQ0wEc+g5/ZCrcj3RuXcJeGhXLG8Ypc+RWBtLmP20BmVsNEL9Rjbdtqu7
T/6tP7N4CA2IJ991SyI2R2MgajxFai97d/NA+C+2iTUgYegp+chPhPh28pBFZHghno6FZOl5I5zI
NND6nkNZSgK3F7CGFuO/qbhoHpQt9V38urmjgxhDtGcOVJT6JhlxPxdZ/Q0uMGRcEeljRoTG1VcK
cdqf3n+i45dcvfxmVkE4B65+MMzkeoJXkxus4659MdyLngEc/YT7BXLAHJCfMqVK1EQZ7Z06GeLS
OQTmzHFquPMKA6WUoekXYIZk8iVJbJV3MTxDUyDscxb9qcxepOxn3xk1thIAlN+CVDvCRWWrLlXH
IIXZPabDugRbAg0pnvym9b5CLZIqsAYw+Kofy2VmwAP4/Sa0s3bMnQBZlEH8vWdnuZSuQUNzNNOF
KxsP6MqUsajoiQW0fqmGRqOAUsFjLQv3fp3AgPBVTavUhufc3iHL9hDndhF3BD0erhXfQD2WnFfa
dj0nSODuxX1PcZiFer9JzZDmTZnULH7q1MIddCDnPWg8s06EXplyvm437lngF45qZ7SlL8WWt+d/
9nmyLYysS9zdBRlqsB3vmCMbfEPUgQr7ChcciFGpVUC/Dva60uqhpZTqLv7O2NdRoMv8FRo0nkLe
R9TVW4vRfNLYpEWIvJ1VvyE1lYmzJAn2Ckuqz8SiYDabTY0L5XS+MT5pTfEWHjnsjEIGxyZfexu3
fBqzX6eeoEBjchLlmTt1ow7VGLQMs5mi9UBGSGiKvcdw43oXterCz5DxVJx3EvBisnxx6EWTQH87
viZskOEVo65npEuN9rTa+EIC2YRL1OrNbtghLKXFLEsPPD1hr19slRuvXeXDq6Nm7DiTbjA2ahUN
mDbbIIL7OlB4qfR9ylU8fM5r5VpL6Ts/CQgoqdXj5F1Xz4GS3+rtq51imE2aExwAjA8+DYYRzQxG
uRe80u7Sc9mvqthuPwPeT4FADmUS+N7TK8evpWGVzQG29xXWAyxhB+amwLCa6Pndw9Zk87sKdt/V
BTMgnNT/eXCldOdaaAu7xcoWNJ0Dzedgc+87U7SBLRbT8B24gj6jfKHEQ06Xg7ofjr4qTXjINI9v
t0e38DcuLqvYPB/E7ao+/RVN2glVVNxPwv6tRyaRdbjkHAc+MsTKaXwj1gtlD8lqI+NFfdUeg4ye
2BXrn+2KSDpWQCvEzBYfNr9ZvVAGnbGvpSldnHcFN5ezHnj01TZNqiCtabJWtUlaHoDbuu6hXUvA
lwBVytg+ICfQ4FhWouAI+iGa909JX20Jnethv8U6KU36f0o5vlBIx+Hhb7mwoH/eqtZ39xNeBElJ
mZn1PgvEgcXSBfPk1bSoZEQpoq/rlP3ONvyqWDO5whPYg8Id86Mv7G1IRjPcQrdZjScsVGiYvFrD
Rr7em7Vp0UmYmIci4El3tem8/5vEIuIsg9g1TyEVZx2Q7TBNZBQIc2AO/DI3+V3LVA1EmoUTn5Oa
FWr9zdENzynkPZKpQrqlkxETCGC0tAeYZ9Ch8p2q+2bKtwLsegkf9KuoQt3f3DkmRETztKL0MTQG
yUcNSIztbRUs9qyV8mJP5LXqIkFcx9+9AZZeBgbMJ8JqpHwLdBuo/mRVXkJ15BukWc/xLjZ5PSuz
yXuYdhbKjvHOlu2VfRGnWb61zmc/IB6hVk483MrBlFvDqHuyy/JHUI8nddDShoq5/sODCLkTlu+Z
DErQfc7Ys5wZgzdQhKqb2s5BD6FllXE0xx2yQ8PvcJ5heUZWFFNrH1EgMaxyc4u/IkAYAcXNWbn/
NpFllJc/R8TGuIya/ubtogWT4ZJa77fJ74TwLY6OifCDSF5MU++IO0UuwC4J0hAZyP0WQ6bwy5fU
h62Cwq7hprpN1bpKQRRZ1IQ/CeaoikCpBMXEHvq8yWbqSDTjPx5x8RRcOit44DaYj7n5Tmt/lScV
+uzUjhXPhQ4dWMPIZBVnWTZ5mjBXTpUYcY2PlIk1L9vP6l5FHyF2HIBf3+OoRmDVbPl3PbbMVaU5
lsXCa5xDEzdJQGi8eAgSlxLWyBSyMnaMZnP6kdPeeMw5PBTu/woe69E2DRam18ntzlpAsz8mM/8A
VtNiL3ffmyIqkBAZVixTf9Un+Mzr+AJjY+He2MBLn4deRj4fNbg6BH3RMpG9VpquJz6DeIKwJNyz
vtcnH3dpnDkCXTMKqRsy0wIMobM638eeg3/h4TIGkXQ52w/Fl1uDAdrtW35EqPAi54dEMv6Psai1
AY66v/NyjI9ihLiLgYhHGymXfxDEvlKOoWOB+QCS+zLb9cg6iTTu5qJaA3Qdahbek6MnS2q417SD
URnQtezTPryzWn/N96LofEBBT6o0KKl3tMeWkVKRXlccEOAFE1tuDpcgB0byJjb6zgfCdG3NQSW2
r4fxpVoNfQdQY3ecUXYZYGEIzAOECQXDHTU9orW08Tcx3GyTsuFsLEafNbX6LIuyOT0rFRZ2YV/e
+jvuNGYcxZhSsftTCHW7+1hMEdiAwueHknP1FlgFmIpIhzdpOBGnC9WzHpKkmo5Z7OC+fPBsWyGg
dG0+LcP7ns644Hu7j5JoM7OrUXXTyu3xKyK7fdtoJSD1TiwMR/WSKApwYOIeSyyI/Ci5/6W+vnNY
W4XIEUuDjhN2+Oubzh2zKZnluseEZ/7ZHUNKQ5dWsiFI1bFeHJxymHCiIAWn/izwXv2nW/TosJYk
2TsOs5kzMasxnGwto/bWeCVMWFuN1BK5BDccC5WGnJVOYvq6c7kPdvxx694MeP3vGiMj3FAqEX9a
CDbNKjSo1nUEW//r9E6AKVuT+9UjZTwa1PGBnqp9UFqZ/ADg2Yjjnh+MpGVF32M77qQoT6cZBAPY
+mjhGgHWEOEzcoVSG7TM3DGjfxFtHLYF1Pb9nxmRT7b9nXkMt+Qr/ZIMETmcCWRckRNKr2RUxtGC
yZav0ChGZc8xDPMUOsXOVRxNBkqWdMRfl7Hpwd4elzfBKKoAeFIr0YiqtgXtMZY+gA3m7vbSSGBq
afioiLqvWGntMrIZOkWiVzcMErxIBOSyBblHdrua9+O12vL5PN2CT8sTSCSaPe9D7uCcmMjQL2rZ
gfoVGN/q3KE/EsWFGTEwL5rXJdze/Mmx91qOYHESj/1OOuOvx8mvWlEc+mwJEALwR2Ggk0VkxzEE
C00+u9IvmFPXMoWbZ16Vt5mfWRxbTRYkPCb/Yt4pTE6r+Rl/qABDbP7Vy8fzeNQvZf+VheCN55Nj
sWuT3Ig9Ic0vLvd6fA8mGee1EKr6JXjLxJMQZ0GIAbhUgyXHeOMkwVLkJu1QPemC9kLab9evU2s2
EcQdZp6nsEofntQ0eG5Ff8T7NHrulRDe5StpVUIllDSVEMtfT64Dg9x9wThK1W7Q6r0a6LqKFUm9
Qck3TsmCNFmFbUZoPuD+30nUZlsFSIshisZ4baIy/9xGiE5PYclTdx3yqcHYboRPScSRJvayrm0E
YCSmkQ6p3c4gzgYOzZWAP/wOeIBAEDDB609HykgQSqLOaQXPqPUaagLGrF8AcET9p46Rvyib8VVl
C85QRU+7BM6/qN49r3AsUgEBqfeGdGsbgM1QJv8b+GuV0Eq/IJUuib5C9z/JoEhdQjQrpVMdfJi5
6qMmMQAudihJv2dHVysTvnpx0MA1r77M+qDmq1WOicg2kMGrXmzlNj3oTupstkGbct3+byb3A7Mt
GELPb6U1+HSQOIni2JUxOgBQ7gYiInNpIRxeEplf4gSOnpTEg8zondysUCB7UuhoQVaoDPNIy8n9
sjN0/s98b0fJF3wCyCfqO7zzrGYxN0Lc3E0EXhjkfXFRNqFVjM9PBJ6wvknJLN937Op6tXi7qP67
nQ/JxwUiLFvG1kslhz5ESZNPSmQMlwLidLD0rCU2DwHIH4MxH99K4nPYZGDGDuklMrE/nIcFoCB8
7x1kSYMgKAvJia621/KhhP2IPDT8a1CfbKZ3fO1tUyfGnTTKfa/CrnHIUiqIEIl2NxS9sUCqVwju
PObeCylMl+9tTqoK4x0t5yXgLx4Dnf255WZhutuX8C2pBE44BTwQxYGQBgK1ZH/+QKI+a9z+7mhx
zs9LIM/SyrLI/AcUhwZu11Hkqtgu06B15ax2fQUmGs2GqCeTSs+Fc9Pbl09wmCYA+5SdoQGm68NI
+34Az7AbOT/wTbzoICFPCvAwxJsuYgpfMgnKOd8TaeGylb5tfZnYyRUWhbBAgCovpEwpnLGI+uRH
6dFFlVfwn7qUCcrAVOKoO8+kJZOpfEUrtiRzA8YdzivOP21uzJ7GziK0sMxxVPdS7iyhDNcAGmNL
uz6tFj8vfE9sSPUFtKY2TsK4t9vd7ZiVXLQjQwjNYLZGeEDIf14Qz3sR87JOy+qFuVw8sVdr7OfE
u5n/1JlfIlg1cl/VWgF8Ao7fLFOgv9guEZjx2OAxoWMGXahb6ScYyaOIj0OdaRZ1NL/o/act97jc
xavaYOLW74naiCp9DfpN4DDO1YdzbPDYWss+QlOUJbEynoMSN3U0aRYAQ02wE8m1+B/MaDVihS6P
zPrfK4lPG0c03p64EA2VvUGzLmKU2ioiz3wzs9jZonJi+6bxVh+ChSWgXWp5ODDSZexGgmv4zybx
WdIUdzXy+4WLf2PC6kJ/FqGd99VkJH1YDuW9r/ftjk6oJOkxQt62MEK+OzQozfw+M35e8lma+pQH
dBCEIf3ZUAvY7eQa0Rx+Pd9PgPcps8GNdhfpCFT8uEJQs9Ah4JeD/cs9kACDzLa2GiWVEM7JDDaV
cyqOQcJZjEQ+qsMvKvFMBcOL3DBgFnCg/gr/Zwu8XiTLm2JTjhzWuxJhHtqmSNdVcVp2K/Gs6pv1
aqHO8dVYd03fr6vPV4qiSTRdpjtUvLmkxWlXBuC8MLa1u0YFcGGbMhGg0sua+CWgFO1ioz0rKm6q
5UD8TNKB+EzqdVPlja1v++Rhl8B4rXd/4Y+HPVm7NMQRPe4/j7I6nZCcfIPosq48PT4y0LX5eWpk
tNDvLmTbKFDc0NP58C1XGqRHM7J2r6n9mFrbHNz3J9IJgMmMcC0fLFxa4sl3xCHLK0ZRzjz62jGl
jA6jkgKFzQ66y0ynVkN3UH5C8H5kkrI1JZWcaITR+Q2KloP4aa3cEPSkwLzd4xoHOkTsPWQ3Ety6
ua+9D0JdwO5QWkkgaxW8/gZAUMrWeo7Bkcbf0GD+RhVvlm/r6LJ2/wpEYBgP7PYpesi2MVZ/GGCo
CYCZe7w02TZMhCLRy7qf9Rwd0N4PNVyE1NZf3g8F+TI30iwvubk2aZAGeut0iZjZAtldGp0ANdqD
18t5qa+RC1mdqKwNrp8jEpdSEDEPrAYmWF1FVVNwBuvAY3YzKJEIlt2OHTHMO1lc/m9XcX4DQ3RD
G5QN9Ov3Za/rkDCei0wSWodQAKvTStPnJF9rc0WU80IpfqaM3Gk4JpQsHzcPPecEtKfp1eAm4cwT
HYcFcMWk07v3/XH5qRGsabuQhESePFHemQLvUL4MCtCdcsRTILWC2MkX2ZEQtbOG+TbeQ+XgPl00
IH147WAo+w9h+NkMDFdmaQ/MairJZ3nY6d8IlP0Nb871aBxvBc2CLAbG1JjCKzSraWy4TBDDiZPk
agyDD5ALrirulv+5KlNwErjJSpoF7dvDKpnoVJMcxSYhQJlo3K3cdFOOt8iI+ywoVngVeJLds9cT
BUPO2zLCspD6lOiJYwMLWEu2zlQ6X256CWg9xrOZUURSZS92vddAjal/OZmDC2AntH74QKHqhd4L
Z+K47j1amxGYWJX2nNh0mCCm7Yo5GtE06BhwuHghd22qykK7UxxhmOqOZGmf6qO+MdAhEzkIaqjF
LCGNZQrayvnZHQde5GHksbXiXEzCpEjRvxUN9MvMDW0Cw24Dxxk4u+OhIxoGCrf/wW/PfBHe+6IX
iwb69fc890Smh09xgEnbQ1qSA9t/saaz1CfK6qf+Q9aCTNvZWEQicrNuYltFKq11cVqcHFr0F0JO
bHS/r/mVPybWPXAyoFUKB4rfx1EglK7WWugnzs7MEYKZ4HJ2kDMRqhGWDBsJArgyQ2TCW8Hv8KWo
OkPqtSzL9f1volng0FBwvJkSoHEAd/0c/gdoiVQzD87HuAHDgI0qmHcGV64oqglPXa9NPXFv61cx
xHIUo4ipwra3Kyf1043paXh2RPvyqy1eP2+Mk9k9iY4kjtWo03Igk0CUMpSMF8oBudamuiIBSI96
Gu/4AiEvnUdB6o1UME+wZUxUuNhu4qb0X1dH0mNcxC0/+2N/FzEt/C0PzDH4GkjRN0vGGuJwVRx7
aO/zZGBDdVt8K0D9NF4aelmFi5UlIulE9KKS6UooKAxKjaheSZbQj7efxp5uUau7TKa0zzhovljC
Tn5QSGbjxGkZh1VoPfF2yK8F8ci6QgaPhESYWS1BMsGQr9YJtwijAf7/8VqHgmA19cHvYUbHG87j
tkXa7wEuANN2U6wCB77MmrvQPICjPGMYAg7iZHS/Wkpr6ZIaGzuDVMCgoPhAE7N1bfJvzxlUU0P+
LMoyzmKXlcv3LGOUmw788htGyeGnqrHrAJSqtJitUoEMY9Ab98c0ZFVI9WnCZ3DMccAOfAnUwV3w
To7rFwhOyLNqnkz3aWv7udeVA+SO1aDN3skT8Onuq1KrYYkKP6LB1ITkwn44Y+TCb/jG3ta6ppVG
Vslk7cmycUEzmG8aNdIDJQBm89G9fUG9jdLHctwBX/i4NULKz8yWbufJI0IucFM90d/tMJUWHT1b
9ue6TNljzNUn2ziK4p1oMWcjyRKzAj3CTHeomZ6OvSUDuXvKYGrFO2B0QJtHH6CKpe2QXCNz+ryj
OPFwnekqyWY36mVZFgwzOJHA1H0cxFIUpLv8a9f/K1nvqQFM5fdFvwbNCFtzUW9ex6uZuaNMht32
EK57G3mB+Ot8tMWsohEmhySRPh8bzFVy0MdJaJO2Ac2CEZiWneEa8RTz54ETUFvPn9sULAD5xwbc
FRD5ikQ2HlWhIXnlTtBIyTxy5puwtCL4OqRcK3DHCVNUdjrrcqUWciSLuYDOGMrNtC7OmaSexkJP
ei84VjI7NjsXMDxsAvwRHEUxSXS+hijcrjvrzQoXRH0ev2FwCrf1kEy6/AjvgLz/507txWWjhnRK
4WTkDUnfERpS6fMXWR6bd2FIx3/3Rls4AFMC1LXJL+81TJ1kzCwOfTvPocQh17kGGqxpHIT5G0Zh
5fGOGDYj4EpSlFKbD1FEnG7Vsb+MIq6MxhGLs0uTByMxu8GiB/klkl2hEuC9jlHIL6DNmS6xpecE
KLRiMdZtYx0rHzmdefPde7j0ldQ+pakXTx+BAIP28yR24yiW4jcBRpInQrJrbFrRYn4jQ1NeYoUh
w5ATomioP8CkLHwzNS6IaAflpGn9/UhqgVw+Wt8rWwGV/ocPPbdZL0sFdBcunXS2Pv4wSsDHGDSk
qw/Kza4mgIQYHC/b6LrJ2nhahywxaofcprsl/4lUErMIhJvlUKpzip8NtARPE01N+DNKZYzsZB6g
6+eVb+OrRmfLyKmpIwsMN4cUZVTWHXmcvEWH6Jg2xDtFy9WmXxWdmePhACNpPdmUOIdGpPUfZhcY
mbcPg1IKjohKNtNi/NqNYkOD8KtyhxMcqpknuZofOFqN3v2hil/BgEzMAFbvM6WJveYtANZd3mkA
3SDE2o1moODQPGhO68N2gedBj1g7BEK9V7wJhMmbZJ7wgXG6+bcSjzgJ8gFX7IC1ho4lD5HTzfIO
OEcgtp9q9CLialKJjwu31LDPe44A++WCtgh891d0lav8IqdJf4+qiGN+oeCC/4mLk1GPb7NaZMDW
0zjGc0oWwdTY2TOKZd1Jwz7b/jfcVD5q21Vn9gcfXclDwuBRhJasxybdw5vpkTWbhkpLaiFQ4QY7
Ay3Qzt6ksbboB/kFGoTRI5otTxxd6MKKAyLfZOhEQmotI4jgHCbCmvaAcDm20dtfErgduAS8tHiG
JaB7gIoNWbt1B5umIVmIei5+xIIsSr+KOgsCbPW1T/wJV3Eh7lPUnicyEtHYBQtfos3US2433OVH
YMRt4PmO2qFctglbzFu9atqsoUxb4wqXGhOSRZBLVAsmFQgiHLcri+h26/9DMJtxOl0x5Ak7DdiY
gPPaUf1TmfCoS0doXmdFn81A7YQJ2d4La9pz1g9W8TqSb65Ubw747b1RYKfLVJ+vqWb0nEfq/S8k
YBQBFlsqtNnldgiAoJPpnIOdGOd1wUP8+YGPp61+DCtoZj9hFt02lpgLjlxkesSIi4fIyHYH3zI4
1JB3ysGPuccDSNfHuQEMPpv8XtOtsIS1xaImwXbnB+oscKKD/vE+M/8HbXwg+tQ5t/HcnDeR+EGD
QFyqpYoBYXXLw9klbXcioG/cnCJyCSK7ejT7V0iOLermmWgVzDIQBiKtOHYaN33xk9g+BZySLZlD
HNPuN1ZUr0XENpIvvxk0oCgfGQpMn6TE49mSiqiV5HoFbK0nZR1Q94X1SYBCWG9jGR6wUYf35QfA
BCSCbl51m5OTQrxMmXeRR9SHkHeEQbVHTlhOhLjWMluSBgMGP6u187ML/GFckmBT2f9mht0svCLm
020JUU4NGKuI7IisQOSlJJL88C+Rat4VelPZxdROW/ojCzw2cAmgbbtmz6e1lN/pQfIa2Ttrxp8E
8eiPQbq4nHYRamPAkHlwLdT1drQN/8KWV9dpEBJsanucZ2biu/+X+w2MlqxAe4hkas1s7fpffEW2
sRk5B6fBLgzkQtoD5ukbBu9czJ1NeeZQYnbqBwrMG63hf/IPz1K0jf6P5aos8cpGz7bZ0NzWWbhf
lHtDMW32cpO0sj4e10BYleDk3gl8jU69KdC1xewmXJEYs8FlZpMJLvlpCga1tEXhtZSB8MLEln1K
ilBgS/F82Fhsqewp8dppr4MvUs+H4TF7aNuG53Xj1tJ9bSdZKwLXLb76c4CkQGPLDhkfwx1NrGO0
MSEhtGW71pgGeE2EZY9a9lN4sBwDa0ujKTjDmNPTRk0Lzwl9BGU6Q0L1lizWXtKLOmBi+nkl/mD9
pjMb31yzSLZ+D76x4zYKA4J4quYyfa4YTIfkAUdgMWmIjLirJ5yD+1oIpIc166LhKYtO8gAWnkUb
S4ne/LJY3m/Po49rgi2bpIZxF2KARvQ9eWCu8ddMw48Sqi6OGAa2hytqLVqFR//IAJEk+oFChM1e
oUVvGaEumaXpbw5YRnq5CcFy8JLIn4TCe2sWIeu1oJ9+G8ta7RHufbu4jG/QnGOo8huzxNZJbo5g
WZRjDzTpAMB6+vDrSDCglZ83zjfthKvK/ex5DWtR+fF902h48ilR+CerqRFrIqTY5L2P2/VWkP3G
FwQCnJqDM0T3mxh+4v00Wv4LDPuZH/0yPcXhDDrS1RMUTm7SlvmJGhBpcl9X5cTwc5vsDr7kK3mS
dhRaCMXjK/wDH6oHKrg6wREOvlRtA1Mfzvk/R1E7mbj0HHzMXt+dYY5EfynKJKiu8h9RZkPrgAZR
P8sJ7f0qVoJZq/QPafcRZoJW1f9LQ4Z4xhIBc+UX/CkUIhPdOJke3tOMN7txIKStzI/3LXSFHBXi
9d7sor/1NMbZ8Zd2UFD6Jwbje6cax8FeK7XcVLeFaBlpvAoQdP0oAA0y/quJ129zL6CSvtU53fLa
6zXCyNFWOU0Oz5tlzwGllT6UQIEy5S5BsA9AvLM5UnYfS4XlVl2c20P7pAIWZmACyFFBx3nprTLr
t/U0DQxkncJVvk2q3UgqsZslUo5Kyzk9X+X1O7vG/a/Z/5YYw3BKUbc7AxdX9/4kGrU6KvxlGP99
GepElWzqaoa4gVdfe3Vy7sYczbVTPzwkjnQLz7z+25rPBJk20c0Wrfyh8UU+mpptBgm3kp6xRupI
hpt/yJ8cYvTNkkkuIkCiTpXDZEbYAi12kVP6LKe5isIwmxINTrDacKJGUgeNOp7+7sfL7V0w3tKH
LCOwcyI6018ipODRGketdAWIL0PaWbwMHvdfkguTqFL80SdjmWM5akePcVZvdTDSxSrIWam2RjqE
MvMQjRaJ8HTKbNNjpNeh1q4bAgyw+AVrCpn1BnCIZ0REatnE5nflsynjnNSJkp3+9UDQ5k3sGXxF
n0AUvyG5Cqld1ueVpTWXluvhGBmDi9uiwzEnP4eJgtfsQfMhnIcwhtG1TPSHoby+hpJTHeJNo/+1
KXuDDENt1PiPOnCeSWi6N7A0hWiQEAgx286CYcIsL2HsJcOW0iI8vFKmfla44IPAARSxSON4zgsY
SVM71kVNa6ehoXF7Fx0fhrCTmd80AVMi9yqVKe2bWLfVvTkBxpPY1QwetAN45Kj6Lp/f1+UemQ1J
XvkAtiNJU8JvqIhnaJxigGbL7c8HrQpM79Qdfo5AGlxifNuIA9i+hPHsovmVShipT6kRrKBc1ivz
gMwLuYC1rhwBjRhpU5cSv4IpCbRT+lQPX/GM5w8RCQzk1KzefafVjNoLevVc1FhmwLsaYsoX+FOt
oVF06yySdcqurzRThbu1R5Z+7u9ZAjzXnW+vPQ0Y4UxpswTdze9s7LxERmqhjh4SbdVaQ9239U2K
hfVCvGNK/GyXdtlEQj670xaa3cAs6y9on1zUel9zEGNrDiJ0D8wIqiXxLnAuvfSOsEoHML7xF2SD
7QsP77YMyDxIhP4vYC6Jj0d37nsGjAN5h9dThTqimzyzbiHf51WCGX05xzDH6BXevrENm1hym/ZO
nogU69Pxj3B0JY4/Kot5yRblkkY6TuTEMz6hdFgttI3slJYZ3v1vFuT1j6BzAkwt3Bcbqheh+2vD
62D2v2n1w6f/RXZi9EfDI4BEYtqoaga5CipwQ7B/vpYiARkKjoeFtRME+/huCOoHNI+s8lbPv9EV
dMzzXsBxGngUNG0lZD94ciJd90YlZOyLx2k6ZtuUi8GBnn3BQo22pxzMfc49iCs/hi3PlBdxkJtq
QVvZdmmiEtx+wR1LrsXcQhZTnGC3WvFRhw2CW4u1BRSgeg0OnA7n7+lXjz7eCGB+Y6gjD+D5GkEY
OH/FXlqtCEgYpW3+zx8pDarbw8BdCAPZnY+ikXAigdIdmsGSkxMkbXLOGP6J9wTtsZ2ez7qmcSdP
sF6YmFIYxXczz7PTG8RjP29VX6ojm+8EI1l548kkTS6tJN1+Yy6IqFXX5nPCX8EVxVdILiv/kM4T
BwZ2yE8d5qz6U92Mjp9MvY6nUHcIcouQnCtw0TgNl7BfT6fHCSd3LI9VIQEK3sEwj/8FH9hn7qO/
mzapny7yM+gPj2UhljssVylGUSdMjdrL6o2hvM4OLAHi+h+DnOBOd5wl7OfAhlJxkqleu8mIXmm2
XCEXjCm6RSMXki0mz7QKEbrza8rwQPPwCsUQ8DcmolO6OZ8iSvRV/sp8jvxnoaAm+C0x6p+zrElP
tksnYu53Jij7QIcDXiXCwfgXLRwPnciNV1kbTzPS90Sh2bfWvAez2h6e3ETPrSg3cWP8xNA10+1f
BsT90n5kXQTRzPPBbY4NHw86awwhVF3sNohiauosTiBdFMLoXXNUVSQ5egLW/G3D8mL0aEV8M4XD
jnP+FgBt22Qh2x46vHLs7C75XZCc242e2Ev3QKJ6GpQaEhCqwY0QSd3iK+a3EtlDOOg1VulX+Db1
28nwhrQQiBteg/aVi4QrOJMYoK/DgouHszIJT+REEgRBqEQjkITHINhIbSBRF2NXgyLstTRvNrU5
vHtKHxijluaFn2VTu8xTqRbWpF5lX6USBdgo4+s+3xAq54MI0ozKYn+X0JxSDEC4UfWz/R0Bl3DG
0hStcn4HraWoc+WeFk4+7Sb0/LbJIqkC5LV1vzPArIMkhLfdNruDL+JcQIiYNLG2TlLq6Vghn4FT
zjeizWYzLJGZHcO7qHdCIALRCJsbpmxHFVlxQwehRp9ZaLTb476urz503EWxHMv569sye2jVmsdN
SFl54LgLwMG0BFmV1wqWollzLt89mPFiZSvLhRmbkdKFZcNfQj6Ezw6Rbfg1SV8kBD/a0kQVAWWn
pwk1TGYg2PpjCGJoJ8QEGA7eJPi/iZg9s/jbZ60tyiRlGtWcrvvmF7I0EEV0fQJJIBdmv4elxP0J
oM6GrrUcGsvo1oIGK7IJU6uSiS+b+gLco8MiJWqor8RX7c+WzzMP9zc8CSiHEi3SnPEMEk0meB/1
I0XkKtcua/HekLSK0VFf4+55OLo5EI3N+mUYgGQ3PPEwby0Shu73+q5QQdFt36GPSmaNwvkhUocX
AvmxTNoZ7pGicGVXC4zw3QsLothy6i6pgsgOklJYydtg4pKcbOodyNbucxbjdH7cmaSo77DhnJXA
NMoA3JCDjmPCtdMI7j9Nois0AKukn9dBTl6uAdD52+QKf8+/4nKNkb3TxtugpHs/WsDfAkoUsAgC
1isiipUNfDuJRVoRisYV5zQvp0ZZ8jAIrUWFAG3co1I+0x3L4rRxx6btq49aMV5X74U2E1BQp5gb
Xhroy/lb79Du49ToqoDnfNfIGIdIo0x1P/dBjwsc7CsTQp72N/qih6FFLzCEBpAgVFG1RNugY7ag
+qnq4BQhAYEmpwdB85JDhInexeKZgTHQBTZvchdab6GXBml/NibexMp1kbjWChz7rnySxm3r+pOG
UGUoLU+MV5XwNVhFjiX1alXjkzm/NdE00hAbJtE0tPcfZG6DwZ50cSxAlFOf5u6kgwb8B7DV77B0
2sk+m2ylkq2XqUlAxNsNlwiY+OMNAvbgO4R0rXKAVxuflbsdUM00uFPDuAGTmFBYH5lPNFG3kMCd
ywNYJDCAK1jqO9+Z+WHUj1M1tEo6+pWQGx2+T7aKERQveUJta7SkOkRSwh+naW+X1H4sEX16Okrg
FHM+VFv1Tgu+Dda+sVhme+gwY+7GIOUaTn4H10fAech49PozPlRhgKNRYZwNCk0If2bkAqvP5X/5
sKeIgSo0GamL8U5xDO00PVpkBntOQtfXy7+74iw4GkOBdY6QOpRbsO1LdBBfCBvyAmbb9PyTl9c/
6dr82yD19FZm2p7ViXd59FLkLWMYpmvfesjBRrJZh2XvzF7sHYyOjQF8oN4iD8qmcgGzMyTgbpKm
KdyhnA2QIl9WtSFdIbPE9v6ZavXVP+dzPdBrrJF9Q2nv5cwXoSTgsocwaffxX84IC8gPJomTEOnM
ByFYx3hAFlF9NOQoLrWugWAe2cohQQbedQIyS3V+1jroek3ilnMI9J0A9xe9G7dTH/6/glHAaMj4
Gqg1CMqV5MHAgFry/Cmimx6bxwN6G5kQkxGjORC7D1k8qmViGwwmvc5dKmzVzNHqH89m76XWbFhj
p7NG/cfONugsnHhblZmoBu1eHrTV4RFNbiXsC1qpwIKMhzBKEln6iAxVBjJsnpLJPzR1ds4qVNo3
GCHJl6+pnadJaAGI8VIrDzflPGbBKH8fo1Zfwk+UsiUeyE9/AGd5V3p1DRFG0xon/5lMYtbMIWiF
uaHFZmcnhqHZd5zDLwz+Vegr51JG3CA4Ke1xsqBQkS2J7/Zy4Rd7TvT5qD7/yFNDeQZiz14GNUB5
NNJfK8LtaUK3R/p3xLtKLre44yoBYRxOhRTiAlC3xR1V3Os6bP7j7ThEdHe25MZaWE28t7PAemvN
uJt5eUV3TDR8JlWhIJ0CQO5ogzjTjPRuOaJxwgN82wuKtsJf9414QtH6GStyy0Qmzhi5zrZWDySo
qG7xPP2YytohkT5e7tLZ1vG8hPUkO8b2bZHx+7icGxQGQxkepKXxm6XzFz3X332xbocY688izY3j
Qll0eJKda7jgzmtjl8u3mrtEm12rg11TIukAsxF6rbCrw8WcdjL4Y9anKSNfLoe4dQKw3WSANfVr
DL8z+5hpO/1aeBZyajbpDFNQGsGm1IBR1sxqtcLiT68pqlSX5QtLbnRE/hfZ8O4VR1yyVe1g2c2c
5oPdUl+pwiS8fpZzxIkAoqn46vPPf7V+IkXQF3Ns/khGGntR6CBaMZ9XYMYTQMqVQgoLd6htY9SF
c7IfCj+MnSmz1l1oggERelM7ZFM3WddOvVW+o0lVuy2FHtUQON48dq0j7bM+yHRWNMiMciMsvAFj
IIqD4xYRH6N0R5dZc1x7uPF/Eu+Z8x9OHcs2HR7uwZxlL4VnXsmD6EHqQ5LS1EtTH4KdZtm2snz6
pyKK9g3shwOxg4JIFkTRKFHkP7m7rWgVaDWIeyi+tGQdPt7e6NkgL/ioRnhbwtFLKjCL8s/L5LJJ
E25e1+ufhJ0tbxrvTiqPvk10T9ia/Kuh4nCxl2Hk37tjO280kPiYG+uW7CQWCZ+A3MfPlXs2ZIw1
we1ZSMFaJgE5lKC5xr93GTXHQVde4kcBAo0T4GCTfmgb0Hk3w9nTMX2O+ci2Qu7T/Q1xoLMbH0tF
iHzWnc6l6juyNFc3nYffDz0qEsZRFiSsEBZC4vEJW/A5ncjKfHkp3uPlZs+oMk+JyC+h8WlHSBTx
4LM/7np0rwOmu0hd8T+MuJq3FPpby3zf5Pm1kCjLOcxEFwvpTIlEMbtovwTQ2r64diPQuWRzr+bH
tX/pjqdNTj9zMH9WdyssK7kYS+5PY8Hk08S52tTGsqoHaDlyKNe/69jO1uVehyF6mH9lrnY+jbdB
xiOM69Ghh1HW45U8IfSjyBAR0s+wIkOwwY4NtVahuw31qbG1PUYZfDoK3CY+0xJBaAdE64O+sjYY
uybgIu0NuScRYgawFb1YgUgHdvdhs9NthHTgQlUDQkmeof2KPL+F2t1ktZ0DnCBCua7NR6Cv76K/
siQw6N/n7dk72qXx3tUonTg1sUE8CjWEA/qCuoXLFxeeUkOD1Z3I/hA/swgC2SpBVzaSoS+Pl8uB
orLCASXiK8iLEo317IwSCLX3P4MRzEb9ALOkAKc6So7Z14Q9xWzKixkjaaD79a/iiBICRw/oq6vl
RTlOiK6ow6l3vcmHf4mWnZQLBsbfx5pDU6xGL4HkXZ7pNL4kqzKvCAZ6nvashqdTKeNGxhNgOUSt
bTNczPP7BWkGZYE8lC55mguP9h9Ilsgeop+PzzpSCKJIdctOSKEU5pRRldxsMUtk0EjheBS5O68n
eg5mUuNFjhooO4RR0CcXAxNOUZSpmyvO4vFCS6qzvQomCbblCnz+T67U0jQrlQX/LNIAcL0TtU5z
RE3yI9cj0JOLAIJH8vtWgcoFadiwZo29bVaSrwGLotmaae8yuIuz4FVyG7K6jgKG0EY/iMoroHI/
1MbkpmF0LmnF0F3zAIggz2UK6RXkMSEoCPVfcjdWuxqQhTEiU3Nnvgm8BEMqAHKKsBD0Lnm/EvVX
M30p2JeW5Z9UZFf2yDDkb8qfI9MxSMBcXevoA5y087Vq7cy7VPVNy3Egq+fi9ovNyhfFTB1+YVS1
T8vw6parETioxlYFefA7AXIfiiRE5OfFIhBDj+ze85Irf7yUSz9m7oPF+/B5Vxxbru68OUAfxR2w
MeIiRJ7FEHVNGjJy652TGYLSsE4a8mVoO3T0tq865unTuL6bcl3nIxDgev/MRYw+XLniV4A/WvPH
hQPm1vxEvyOOSXCfdQVBbq7IhJCDenpfYc5fdD81sjHaibS3Q65WFM3qsCAMRT2dBXyuqjz0Hcgv
Uqa8rHmWr+6fEne1a90UMt3cJ/+FPH943XB0lsm0PoA0cICVDHGzUK9SPqO27G90SqAZ5VAzfpdy
6YXQoC2ElkhMb43BswN0/AbxRTs86PPhP+Tzm6udG4QsE+1lv6y5oAF/X9hlKlUPiSbuWvYrLF4u
sXBIYzA02obtdGZXTL8C3p3VTXd+Gb/+IPLZ8lVoVoHY5AoGz4AXhlbJeSekFyYL1j68nhdkuF5b
9TfChHLI8gpd2btGRl66B0FjlL9HU870Soyvc+CnEq3KBnRKd8YZuoodBcSIkCfAG8zwjNOWPIEB
lW2EQw6lwCO2FqhYdxMITKBc4EtcrRFxWhpJ6KhSqWfvuITsILr1MDHCV3E6BCGwq84iIwNWmrL9
tIYQAPEr52mhlp/IXKyz+ZuSjITOyZiqvhovNWOtQ05q46RY6czAHKgLjzPB48VjVJYvR4wGbmTD
uNo2405cN5F78HJN2lMac6JbkqMHuFQm6h1csrX9V94DDOxlpaL5fB1o98uQ1dpKWkhrBsUtodpd
lEQ+s7RTB2bt1UW7UygWW8MMWaxw+SGtQekLcVJFlgu9vYUeId7tJrp4E5YlegMNV+2EaT4wOc/4
wDTq1VIkG711T5/pQnwPQI5N5ZTnrCSrUH+y+zbBTW73w/RQZQDvGJ0GBMLslhf38SkBgrTmMolh
To9y7Kab9+y7qfOzAAAvolOLCjyV9+5XXXRAYqO173DjlM7Sb2KPytJXBKnCbAoqw5DmxNdoZVUa
APwQHOEPR2WirPil/cNJ6kKURhKDVABHdZWzEadWQYqHIxZ65jLQcXOn6alyB1+zZWJphIT7TWxV
sZjxSNfnqE8zN/mmpNCNyoj2TkNdT9h7KahH33EfPITONlgUuZvK99iprKUteLgcZ1MiKMsO1VM5
8vPbUj8rUYlEPBG0XcpQknTY71UbLTj6TWbtFr5GXL/AcRtATDEzN9fkjYG3rKqxNjz3HP+l9fSH
TeEqD++YM4blUr0eotVeLVZvPJmNA/+gjs+ebtaCUQyZtS7pCO7MR5pbOEprbig4XmwoTBTv7xvy
KaoOciZr00HJJ2TAtLC8DWtpCATlyeLuk+DJqVwiXKg/mPSakxboIjtk3jGl3pcJP6ao0RGyCs1u
Bw0WTbm63/0as4fHJ4lrcKGUyy2DX/fROUVBiGDe55y9Cq/fXSD/t+bVisWE2JkVLFtwBElFjjf/
E+MvM4cg+S38Jk96r4f5yrhHn59WR9YH66Jde4R5MSpSH3vV8BMAH7reZ1XvvFqmZnP2h0T0kwrg
w5Z0oc9drgF+0JJradPD1gxg7L1ddkHEKTOfCOvQjpFbGRlUW3Q7CMXCMyVqBedQF1TN6oasKEQV
fIcOCJz5+XMExh3ub4oO3pr4/2Zjp4JKmiJmBkZ3VCT5ZzG0EVeZhdcUZkDrOu+1R1akQd9dOXLS
HoeT1f2jORjMe4KHaSQmwnil9jJsJc1PC7jFNqIHUDxtsxeEdWjtd+6zVOQ9J6RT1GXsYhLczDtT
hNCP5mpQtNxmU29v4aC7BVJZe0u3wVQ4LuC2VVkkKyzY/zw8cQwliIx5OEL8ZywnuZuEzb2l/O0a
EoMb38CEJ/j7XgVsIJvpzIFi4LmxTW8lBoGxIBIslRLGYPqSeqhG1gR98c+JQEl3Rijne3leB23/
W+76+Dby0WaN0aTczq2+GVkwydKoIY5FjTgD4Kroh5kWbGYScbVCaZZcNb79TlBVUoB7KmFuGIi2
aP8BCqICMdFbVhb44/skscu9/PCLTUn9RK6hpcqUNCEL8Z4byqsmqNkutiNtBp53eBt1HA8fHJUR
KFmuuhZ4cNy0yZKcNtGINRdriPEwVJwy68EeZaoExvVyCEHMxMK+3+9C6eBSMDg9j9k8pAFBpOXU
PSKAZqVcO1iR+/c+ubrDO7Ecy5UbxZRkxm1Fkb1CTUDU7cSPYsrR7n36kKhV7UeC+8f1QGZm/BGW
ZwMIzWyo2WY0n7vRQ4raZalGYK91SiO9w08pQ8GRQd2D7t1TUMECHCHHz9aF6TCDAPNORISCVTZF
laBgaEh0N/0FP5Wxt4CMqHLdsKZD+QJyNqe64QJ7nW+Pqqm+3koENfp2Cam3QfaL2GuKKOog9JKD
2Q2gyg640b3zKzaBoFzrTUGrAjj50WAK5M6AdHWXuuvsbD7sCI1h4KjQVtAYBJk2RnI1bhLV8j+e
SGG81Eo95uTlE5powSXNOnpOgGhj+tEIZAOWoBAuNIzdI/QfkspTFbgvevBLK0L0CD6Q63kY2msW
XQnxuy7QMlnSFTIWyqBRlbwVCA8IMvfiQUxNFXFzzijX/csxYdHdu86+VPRzo8A8eB7Wxq8vRVMT
5AIwb0iMYi+xA+cRNGzhDWOZhlvMt0jdKeD3RP0jXkE0wPxWJ3E2b31fzFSwxSDrlPC+UB9LcJTV
IY88vVwFffImzt8Q9JCQkxq0eO7wKjLnayOrsEmefKi09n3B+rzJRMcLJ7VlyiqKbCI1NJ3kzeGJ
9I0CrabNK6uE80NgCuBiXVvm1VVxzPVsM84cDBTwNt/fHB+5latwQvZfj/qkcl6vYcUo4P0VizPy
NB7k3g2FjMHjLHUvnBZZ+Hus+iKZViiGWIWWFJoYecqLNSc6rc++vUxgIinJ5dD+55LDlHKgt7D7
FLHApSQ7SCnB+A70AfmiKeWlZviD+TJvHN6+ofNjhVoffW0aeA24PYqKV4t6Z0iAF8B21vhyPtVD
5NYFrtwxEQVtqoJLLnGbmErv9jbTROub8XW8Cx4cP9rQRn/55ZhZmODlgB4XwoFK24kB0RkVclxt
kOAiQsZIPEfHRCGg+0t4apK3upIFoNUSu6fN29JgfZr2eSAS/K5bGRi8YluROhbeTSqfnuGpprlg
ElfWhaZwC5/oBKepG/OFu/DxJpoqmi2AXFPLZbRPppRviDoe1Jm6rUzF1ouTx7NNUCXFt9pFpyC6
Dwj9jn+IwEJ5bR/mKGEoYubeJV6Fqsgzf91dSlknfdi8zz2SuT8tUMdW15kSY1bdBTfudNtJI6VG
9+Kf4N7YTrLom5pSusY4KckASd3aIDwBXFrLpfDvAHFBT91B15ckuWzTyyZ/K/4yTKwAVasolFHs
ZzE1wbU9TtnuCt+6Fd93C9uNuyBhVdfKfdDXOzjVB6AmnclB6L0bG2IPTVKTI1XJ7cXh6G3ugfiG
5MVKSlXbFTvsrjZOa+nXA0zj2eTinwkSrNxJgm6/UWBup8K2ec+QTyRpLDmxOKQ6Y1+BrGMwMLis
qCAUpZZ2nybhBqDyZmOqmdBXevnqhgOutOAuCJ3Zgz0xo6PqGjY2AzWVPUsq07ufNnxzjB10tEfk
EI1vMjXm4N3MDuc3OOI/wdFmrE4QMwFE2RUDjp1sfUXOxilwtv37Ac2EgHfNZXPUGX2LWTQpxxa1
QOxzySL3OvockefwJmF58SFBD8NZ4ymCFO/YV3XalolCjbC53UnpDluJsTEZw5xIdoToLQMkdCZh
JZH02rNaKltZA1gUWM606MjAVzcxeGGF8zimKanEMV3NAnHusDMHG2sox+jTrwFmIFgaUQw85oIs
+cC/Uhx0Gk4fNvFB2ECIrYzYfD/dqfoUnNxu5Aq1kg8oYnaN/WpP97Exy6PtYTftBepjRqIyjpAs
052lW7qD26tUBVPk/SjbmE2Jdgd6QX8NbeZ+RNmSSpPfvP6lUF7T2Tl43TSU0d+BAU35wMChtsyk
6X0H4H6qYUlRjMD9goSye3KvBTGUica115KXvt8qKwXmZ/ZuBknQcMCdw52bKTwaJ97EIeQ2opnB
iQrjQE+QZLBuv7tgQr9wjP3niYDZaWF6MEPiFX+FMbC32mN1ND3DZh8PSpcWC5JjYEX8XavTstu2
gP2+UyA3ZplnA0aAmZaZmxTGYRP++wYfFev+1EPnWBEZ/xnSqSN0TLbxkMajmxH2Pqa9d60sCdfH
3eKdQYO1d+686RIL4da6OD7msQjq8IixKi0VDBIHHo9ln5N+ytZPpHyxEzA5CX2Fn50BdNUjXEaO
zEYG31fcNrbYmy8Zd1cipj+o96d7aGWqHBFe+FHTo+7DCB3QFgbXIH4LDIljDWMKwN4zvOxtmcMh
dct3cqeOe+DjFM2+CVYoiTaQX5rTwwAkpvLxsKGGVepWdwae5PyUGAJxcwQA/lKhx+Bh3ihbu71u
VYdGaXZba1414g1nT1k9kwwgwhA2JJIdc7wtQihkCnJsKpAOaGP/aNzIj9BQbgDPhvefnpHjdfWV
/gYfylTUYTW5msmslh/Ak8nP3A37Hwb8vCsWp/zgfyZFnzjbnr0XVtxqbEIH4UcHwBivfNoQhd9/
DFAPSQ4eXYVvdUekkhYIXGEKXgkwRmmm6+TbbI9HCxooe4GDUIUvymFkHrufm2Da372urRPzaioR
Cwf+bWo83qqhrQTyafXg71sYZjGvGDrs6nmUNJi6UNuSIiUtTvh/mYmy5fj7pHk0JAUNEEtmb9c3
xjL/+/SfRZQ0m6v6jmONb6/dGj8yFW+Pega8ppaEhA8k8Y7wNujo1Eu1V5upHzDm0/bJL+p+r/wB
0o73B8pb0kU34g21dfXW4G++Ru6uuGQcRZwjtmck0Z7mRShaX8FQ9WZZ2zSvk4k9x0o5hsn/pSQR
Hyrc70eDkVs/Ig/enFIgECd2Sz+8iMewYmjnwqqL7rFEJmmr7SZZfztoVV7IklXb+LcW7d7ilVdd
XPjeBVGdDhC+2TkXGZ5zQ2xyBGBxY9Gbwss+s1ovj8vmjjMl625c8c1dzGZe1EU67Vo7Mh9rtwid
4y/iAAI+C5AJA4k4kirgY+lpjtIu2Gee5nxlID1Jcj6QT7/hfX+Of1l5/xQmT9qlpKCX2keBM314
uXE7IKcRCxc90h+dP01Pv41hdc7FZI0CzPrd5sRHQrURZlP2ENepEyOid+KP30V6zmWNqHVbiuOD
pbM9bMV34k13IUjfwvBXPWQqAAcf1XO5yFWlPJRcKOK548yhuRFsopP09VXPSTAoM5dW5W5ynP0A
ZOWmPudpJwY48T6Op+vwwxAw3eJvGG3NyQA3n0HBsIktNzmVLIjWyM/ajZ8czmizFlhqQOt6G6oc
WFqoM0qPCeYdXMSzXh6tAnVMoutu3lk6mdyPmA2R3OErWhheL3SMj4qwW3pMlKe0cjwv5v9FvEyr
Bzl8UZlCsLYt3CNCf5JZaofOoLHVxbDeBNjaqGJStZtNL+6oeCSTvZ2mkoiUOENlyTND0zpiPk+d
lrfc4T9RG2mL33PVjD3t1v8MMXD/+/u0ragE3f3GlbbHHUUEH0A169sYDWp6KOCmbmyhiwEJuQ0A
adxz0ATHmDGA8iPr8y94rVUFYGu1yv4X9E/OGkLxFBahea3C8nrLcfhiokm9fffCkseSaTbkQEr7
UcfZYC3+tt2J6rGAkf7WtllhrQZxpHO9o3/3/l0dhsM9v3lRpQmMvwxpGs9RtlK/5BqmLk8JkjVS
/yH2PRgBXjtztqinaUFO/wgr2U4fwF5un3E+iRWFOxEIpmRTiMDs+xJb8lhzKIqonFkYNyYOzT4N
PN78RbFIXxHkrqaklK961aYgEQKk7agMSZIREQzxRDhbzGXRxwDhJtmrmeSbsA5Z3tlo1pzVWJ3x
JU3By69Qupnv5ZEJO+kwNAW5xt1mLyPwwI9hUEIZnKeH3ARkvs5BjxRRmC7YUeFjcCe/XU2AC8PY
gK6k+6HkSomIJu29XyQvo7kjKcRNt/pMX8U1/qzFaKrBHUnXKIaDlgntsM5vbr9V5Q6Edqh5iMmf
BbaFq31ZDI/otSEaX2gFtQ+HzWIEhlLVrbaS+SB33aPxmS69aWKC+hazGqDk5YhhV/J9OP6w279k
omwzH3wYT6nf+ESHGCY7RFpgVpZgGxQHBmktavoKraWAUoPaDcJZGhNRX/Czh3CRp6pypIu2VB3+
dbO0fF6jc9sOjMb1FuqW+MgRzXo/aDONi4/2ikpsVXiHqNznVZ8zrdga31TcusQeEgFxW+PK3Pez
MWCUv0koXr0/gk7gaf3P0OFxTaCjTMRszTqFgUNs2ivDl4Oy/8xYv0SkpKtTnBS6OgYQaaKUtwGM
yHh39QqElaRgk0K2J4fv93KMyLPPAgr3pA6dfNTdWpQw86kSvjpdYkJ5L/naK9GRUyp+UiLTxCfD
6ylp9BvoIx+vevIYTqtRg9vZGZZkz6G8NeUIzhrcDhCcSzgJA+beS7t3onPmvc6CcC/NIICuOZal
KcgrD3IE4ZvKLt2QQJIymhjLEj5jnY13NYd9OVCdD8ZKw0PSp7wmaXMSm0JlyVnjzHUyQ4fcaIvK
LN+YRz1gyNtdWPWKlyfohlbfSzeFEJxopDguwZ289U0FkUH11xEEFmJGqrwFgoPP07MWSBaS11vK
O3g9IZHjdf4X1d5JX8/hdaEjQiYqj2MfqxcAuDzOFWYWLfSOvFP3HW/OSN0D3Np5trVY8pQRI5MP
ELnhWK2a4OOdTHwsXoGpJRtjgOVQmK2GC7G37dh75iwcSMFcOjuTQrp8PMnsytkMjXdkQmZbWAE1
y/nFYF4yHTTpHmOGWVMg9roaYnNLks0DRsd1DkTKOrSmnRU3pCgmpF8gdV0u8LWQnFhZUZscrYGu
cGWvyHGnJe/XSdmtT5oadVNfoi6EODs+xV0LmEZRloe7TPeqKlKG74q9br3DZRNKHfiXB7FlWgff
52hQTdnbcBtXyeMWgS2cgZQLcH+nsjVytKT6djEwwvbQKFYpu8ay75uODRklXpb2SI6BWbVmecVd
EYpM1X6WxredrZuklZKZ6D2YRMvN0iYMeH/2vPyfv7drQUsY5JOoxF5n0X0flgPGcOXtabRlc4r3
iFoTklqUcV/s2LfEgmCCDn7YddRePblxymKuBbutQpOs78phPOEWtWtLXr7i8BnFh9MJsVrHfpHa
AFd6Gt47CX3bCM9GO2D/f8+6W/0HLsPB0SH8gAuGYNJCaPUDzsi440wt+KegTxTh0cWtZmUvYs1U
RYptJhsf+4Pl1qsezNFbQiikHs9TUtCcSoNdSN80s7V8d9A6P4hrIPyCX/5PTIFOGq6MLBdMeHl+
JcyJwDs0xdBZowxMDwL6Q3kuenIrUkVdVxq753X8rdLJBwbgB0RJsDCziMm+YlOe96p4PB8TqJDc
3wjVWjQF/dTIVmg7xp1wwIr1f38GKNRi/tO7cQvDm9+tj8zSXHDCI1etVIUNlh/aba1RGJsywIdx
kdM7zodaLLM52vRo9pfql+dk5uC0YCKwqifsOmTKIU3mB+w2lhm8QNJJyqR3ZnltWzZLqJ6FZ2Rw
1z9R3+BjNlqKpn89YQMoYwWBsLSYxW1e8tMwU4slrXT2ANwwcAm5uyvmrH1V9QrAUmBKyY19IiS6
4sYd32Ylxa0S3aMdJEF1MjmhCZHJRBaoT2TGyZqgXfpoEjm+Cj8p5Jh/FY08Tit27FTODcmRyERS
dP2AqZZbHrfqhjnh8A+ldoqXaiYd/YU9p61t6EfEl1Ov6WbtuVb8FUQvnYgt70eFQ4qfD3TCRFqL
m29rWPo8B0pRYv7H+aj/trgCG+u5DLWlVrt9FqFhhZse4iDlVMXUIJjBeGXCitPxMYJtP1yIwlo8
oGN7cTLHyk0/Bsfcw8d51MCDm6HpIAHnnc7/IA7ETZtwaa1L8zxnvr/wSSJRS6zCQxQ6bDMBUR2k
bMtIA/aI5ilg3LK6RegshJj7bDLRXVoujsMufsdmAcIvqzV3ujb6OK15IsDeL/aN4yZXsb4zHgg6
sjczWI9lg8hyTyGVi23RsY+flfN+keLz2D4gVzwhoPup9nh4INfUlGRDuDwIUYyBT/vb0FzSPUHl
WJR4xS6y7N1QLQEGWR2/pUHf1jHwB9hFYtFzHZch/gl8WzFWvEsG/SlWfSlBvxTJ3bQjTlrdVEBT
mIMKIkqghwn/SMEH231u1z53XGPsJYpsf+FdD0YUbjih50tvBL2soEv05iRYSD+rLMYvTKd90lz0
WhNyFOUHf1xLdpmDP7/7PnukM95C7YyiC0pEOBhSAZ5SIwmtAP+ShxYahVFVjmRxK4rd50F9i7ZU
v9T07U/pt1ekPgAp2t43vouKocCIZqjtEXxnH/XTe51inzMYtmzjKIqSdzF4Edx6AT6MImocxiZm
gjhE2xP9rwS8IRVr7s1mE2IJK7JrtDWbTQ26nnpQwYlwIf0kp1ZEAOETo/K7us0ssSuwvCJaCLiG
vZIOTHyaSUUDplEiqcxLlIGUWNSHpFrcizR0NNmMGDKn0CcRBmCqK+98NtMB/mh9ZC7d+i4Qy3/A
EBUYu7LEBSaL1jVj1Rx80d5qBSUkbITZoCLkVqu+1gKVivOALb7BIAD+Od0s5A7uaRBWQUKLGmqi
WPetv1neUn9ozLz6G2DNwFJ1wA6GVMfIyAAt62gPapEC5VT27ZDPSd0MEUXEgNNeNYFvGiesuC48
+30CZu2XJEd82RbED0nN3iE+gCLQo95L3BgdnumtisK5p3IvHIjyxlS0OwQFAoKNWNVxeN8mp466
wmZ66XJMB3NWtat3sB2GXi/OBtS+1l6th2LtNOD9zcFzjduoqr35fQs2xSo0T4V0H3eCcrTCx0jv
x/8AoCoLO/Q6J5lJl2u42ml0Z1/LiUt0wwMLkBqpMBOuwFP8vGiSlPFQCsrKZNCWKuwshcNkbkQN
MHM6NM/NafXBxIge5ZCKRgd1zheysFruY/JNSiftlXEIlR4uN9IK+AJwUEsTPESYKB1M/RmhnIcU
qX8dm8AT4Kh7xmY2ShViZAS33Ee9LePdqmrOJMzpueSqIMJ+xvV4dJwC/gCs2IMYU4Q5OPsnju0u
REQUFKJZAeViomIaKr7IKXa9ySLhdrp0dsZ84I1dXVBbzaenk0eL99IS4GralztH0uPCoU81AO8H
H2wTKcl0rdcxlSfuDw39D5nBHTyMWSTNP46gbhiXdikonc4hIlCf1Mv2FG/jr4nOscbRvmZ+tPKh
aBcq7ektCbbidXh3xUURlgu54le+o6BRHc2crMWrh2jSgcDNX89dmA2sfK00apJ+23mbDYl63tIK
dSWaSxHmcZZYRqkVcNE9k7Bp2a8fwjfgzUyuJUwIM1RUbdKpjHLmhnq9pimTZIds+uvgbyKSwH4d
7swsl9QkynTe48whjRMaoFIBu0Wq246ZutRDlDGN/1D5YZ1PoRcwunpfDvV5vZG6UXDGULTfOm/9
Ap9OZcTKCRmPLe5TTzyC1WACw0TDotrkfP11anJsHdg0WBfkH50djKE4ZrzPnl6pg1w1GIwRASAC
bFv+XaCgcO5iMGnpeMldojUO6LpOSHCgckFlIDou0/s20pKynz5c24ouHaEpZP8cKPzGEUrvw2vX
Jgn9xrODWPPrHnOUqZx1kbfbiho8Q92LXNgB6f5jC7ckqYjE9dd+OMkcw+KbgEqbTJzci10U3QKX
1+hqideKBjiZFcK8q+g/SWyUFbo352E6f+DqnnaR4uPzHaD+HVZbxb+8vyGxPA4JI+LUmKJYBOYY
nFrjZqOlsa4n16EtNG/rgl+bboO8zdX+2xXyojTFoa/7b5ULMpgPqFHRrK348aOnebHS7xyP/rcz
ybBwgzt9Ak5XFInnakV8SwPEWAB5QgcOJbrz2mYDcFa2CLjw7SZ9QjSU+ZkWeDW041xJZKV07w6B
Q9w995uCoOpQWIoJ1R1xypvFMB6kRa2XZH6SFk68ZDhyqSwADuMKyMOYPyAFkO9V83vz54M9Xr4+
MEsU6vj99CfnrBTUqjIv/nhowDuGoOGVoeaN/lpVOshKrbhNKL0+CNx5QXvkRnXq0gwbPNu882QU
Vca3cjqBOiyN+PBSgNHXWeBKSBe+Dr6g9fGv+YGgOgMFuhYbqBPP1EzRIfyydgAkavfM2bJiAIjD
WEhKNHF1/tAYye0ay3bMlwHfCZ7rExUVn065HZ9n828eGdN7bpeSMKLJ9+GozXoGibxb2KK2MuEh
tJlWVdgavoxuvHLvYNYc3o0y9YcWkGQfUcteT6HYsLq6UYYAT06mtI/8n6dEHVBwEykoS1ELsXmn
gBv+02FAvx0Y4ABCpnt1ic1BUjV0pbQfNQiB2WGPGx1vWFIDetthfhh9qQihfdoHyPSRor5YaCt9
kb+YsJE/JLTJTPPanKpsi3PRBBfTRQ2W//bw7RtDvP0ymaEfGEfsog7vK+OqTNIMigbZEbRA0rqD
jC1Q3TR8wxGEY4mIRwJDmAPdyJVNrIn5pZJBGKn37h2AHS/sDjSpM/0nkGvCuMTzlMe31Q4h6ZSk
T0+lCBQeHNKmoTsqio9SUaBVrHOVF5QH7Xg9zdxjRFpaOEcJXHf8I0ULtsEfl0RpKwPUHDI3As+t
c2MDcTqWfoIOCv1VXhdT5BE/J2kZxIrmKABu2PgE5oUdehFsAPeDzm3nAUoJbJkGwL6lPZRGph7Q
ekJju7TXsEB/R8dN3pMDpDOVQsx8UK+RiQhgR8nVg0MS3+YMf0T2gDwXDCpxXWy3DDmZ8Jo3mJ9t
SWfdXxeRqFgJt4qT1LcGxztffgjDlEeRhkaW/zy2i4bkT1FCpKim7PGx86/GgiXoQdLz4w8ay5Pp
QpedmdIy6fRzMfP8SfadvDCo3a5yvmGLMxzYGUxqduHnfOpSQVoHEq2CAo+ifCXISdo015MVz/BG
vPGa91Dw14WsUgpfZYo8LTg4aoJ8b1O14Lo0ucvR8fx4W4tDOYBZyb7y1PMR4qToO/QxSjP6vEfy
jwMEcWqM7q+oCTB4+ws07Yw/IcMf20eqXLPkCK67f2hnHvGN4SXrlDqMJp1jxWWd2Rf6wwVqvumG
drU54HW/8TEKWkewBOHflDVHQtFbFVckofynigvO0KPNwOkrKCHnC0OANcejUtIHR284z0ZdJ+7+
BkX/ReTWvVHCH9jg5t6TbSh/bnNv9UpBCglP+7Myq8slgcB5AnoKXHoqugtR0lPjdsT+rRuDVL6J
cehAeXdqaK/0bR1AmS0wS37z1m7de26UWoDLc6eEuapw8s6lqjOSA2NiShL+pklc1RePeIsZ5/Zv
elo8l9PbB04N2c2RdO7ii1ypYAagvyAeKcsJrT/ur2sBUHjkYjytame3O/OuR0HiceRfs121se3u
zy7qnXX6bNY3wRj8LHfCGpXjzTm8GJiBrjt6jvVC9q6+Hb4wsc0c1nIj2Nb4xyvf3HbTOY9ViU/J
l3BwFapziT6vrmiZD2NFSANoPsS+lT60/4OtgdkF79AHSmMHOEdaYai4Jp+cbV4csGOpbJol8bnE
Ltcg8eAOR06zvPJGXhpMzFb8Bn2ZR3722U954X9EhuFUjNI/rdyPkwIkJiCJolciL6L/Eu3ICMOO
XxIvX3ggoCq1HECTJd3ChAuwOgkN9/XjyDfcA/qQmEOytWTDCUO2DGskQRMWRIgjuH6ZFdzdzvpY
OA9f1QNtd9FLgwWS0CV7g4x0XtF6Oi/MomZHuhkQR7zAK8/TAWNfhzaD/EIDZe86gwV4HwuWk3sX
WYZo3wTiTTpItm558FTFOXeTvCG1bQ6dfPPB3KYoOVGoCSl6HD8xCVFSkMwKKt6yOTIoNuvynZpk
vIyNUTAztE/NoGEWTTBv5f1XyHqZX3mKbT9Sm+1NCitXG95vhlCUv9NLTdnbZe9lHiLg7P9d6bYD
fhXeAi6bvZ7q8BfOVyzo3Ks9Oys9v/m5APi7cuXnOUkth5msyxaOLqR08WZ1Swb4FB0xArrV0pHA
aa8L/4N3fv0zwARsb8fJ48Vxsh1GnCqDkB36nbSPXq3ArEvZqnam0BvJrzyhS+XqFUKx47xSfaaZ
2NObFAeZYtvDGThH2yb8j0vtgnqP4jYA2fOAJuVrK3X+b9gcWmkqAl52CkcrCp/mp4LbcsUspqdu
nJIq5PVknZDrpymgcz1Rn864KMCBkTAgNhLFpXmTwldDi1pUZb3DxNoPPfiow1rZ72OULhVqWcV4
iS9OpPEUp7tJH6g5fSjjmOZxZVi43NCCQ12/s8TzZFEBj42ru5zhf2xsRtnhnN+J7tUScAfkVCg5
S4U0aoSzBqpyYuKCOML+QJgDTxyynG4VfEoiyiH8Cx+YT2iPWjxLsIHOkRa340PksFOlXRZcG6r3
Es8clof3yG7IWhviymqVbZrHkgbyk1adRw00kj0fdkpJMQxyrFy1OuGutlcdcJZkLu2KmBtHkHir
GbWpgb7KtNHDmurEmdEynSnH/KvvRw2PYxRr7Dd8F+cFQK3yxyui3Y38/+yHoTXVDgWPRZFA8rxH
zCscvpMQx2zDOueLAYKOg687j4/HQ0nroxFK0/37z7TKVRWMw+/9T7Z7imxxulkI2mv+aYmCBSuT
HHYvYqP4ueU9Zd2qX03GiEIoIEJQhISBaIMU9OdsgTk+iGVk/kQ4Trdrpj+qVRkyb2wFKNJOka8K
MwuQATbpk7gT80jFcUyWmGER3WJOkLboduZE/YbcKiaeOWbQ7ZJkOo139X8Qv2QuN7mJbXtLYBUL
ibrlBZw8LwoOqsIE/gxBHLHnhrvA2R8Hz14yGh9K0d0JZnP3oTtWFEhQyM+fhAKI7VrOveOoHOYc
kb5E9QGoGBiiGSmvT/qE7EI6pUjq7vqZLvaf4941EgMPxEmVeIKeyIBn3W/YHLetXczifq+YGC30
UjqdN5UCTNmstr1VRZCGT4b6dWBhqsTn0/c81cMSmOKRBGrj6rUocsL/vQ4ZUu0MzfoafvSuynK0
mA+fWzqS463qxg0AmuhvXx8pVYgdaibDQEKue0l9YPEvPhrY4GfbkKbe0igQHdqloO5nAl6jFSgY
yvq8tZhqqJ9CvU/lqFCNiyCq2D/Nx3IZIzQhMVKmaTUmJ6NA3lUrxd+VYjhewSu4oGYRspDGMWSS
DCUKca1HcOrLjQttkKyjnAucNnq6ofQTJrDOsuH2WRITrO3xSwfpQIDWzL1pPMnlOSjh47pH2ect
rsMwPO7SmHMmftvm3hW4Qy7Gthh/hRCE8/39IrGNaxxGMmZT0rA7TTQ8KUFuhA1PKHUTy44TBzmW
nNjpxAhpJLXOTRBRMIrZMJFnQmNAs6fyagTRoSdJv4zp5GUKnMjruE/pBnonqdiM8uyXnP6NgVM2
3w6rINFKtD18bnz5qllDYGXXG2kkaeajGbEQ+JEus4d8pbkL/2oDf7OU8UGNY7vBSHFdk+himL8m
dLZTb2euUM5flAOfQBYNufuBzAsjZd7VvKg0ThY9ChS5KRce6xsT4qFZCqI1is4mjYQ+FaMCVZhj
dTTYGJFL2cfFw4VhTKy02b8A17wBeNpfW/fQyfTVeDAFfrC45c2BX3PZobO3EDUAio9vOacOzP7f
2fAK3N45JpTYNAzqRrQAJ9ct26XwY/JtC+iax7R8sjKLD62zB+8q2zN1x126Cw0TEWPmRhJNtquR
FdMhw3241dg1wiIUODc8x7O840CYleCSkOwXxQHnRELokLuLMhG+okaz+ZnZGRWyOhLFCWIaV4zI
IqU7pr/GIXcEXJk6FBVNl/I7nKueGzT8Sek5rMtGto4GEqm2W3DZRm6kDLXgsE8BBKLhP6sJk7lG
xHfueefm204HOcOxveBM0IPoiIudRJx+ZIReMUcyVxXJTFi/gZidR8Gzjo29FvqqrIHsciQHU1X1
jkBLNR9NcYKKo9+5muWJpg8ZBdueVKBm8x88dC3bd2MB48Ujc64H4eseKFIXv2yFnTpAbmKWIDl3
cw9Lmnf4dfNUPPGBYfwir41+fTgiJbTLw4135IYo1nJN1dUvIFl4MadniFFx+h0kgukuRCCfby7i
PpPiwpiBn2qH7koVQlE4AV95skOxex1O77ReNkNvMC1YxVyZLUiZI3QGSvYkYSMuxZLThABh7bjd
fTC6oYgqSXAal4UxTcEyR2hHF+bP+FAAj44wlJm27Om+tF/Gu2ML9Gs/OAD8JDoPq4rTTieih2Db
nxjG7xMpLOlIIg63EHAkNHs18UXD6PeOQ/gnF6rNzO0glRB5pqkBDoIsKA5NSFqPlIzv8OGEb18w
BKGYFZ+842yvxg8mWOq2qhHfmmVt51rsVAvcWPWEinMUNVnEaFUto61NBJ+lgFKsklK54FrHGa9q
SY0pMx8+gRf35nX3ulNxrENKRcmsYq7Kgl/h77BSzUMpBnAZYCTof9xojNAk4WzdjQxUWWnPjJjN
SaBpuJaUiAcmGUbdKWz8KhIwTfk6PEw9HN/a/W8ZT9M32ic07B4xfXF+E0HMKw89DfesgnG5RLrN
IXvuLBMnVOXHszvmEppRrSrdabx+rpntWquXKSnxfmx+7TO33dvypv4ScOwHx/DDMAcHtYrnFNPw
i/fOjQLzVR3NEDFP8TC5BJh4VaZGlrZJpOhWJmqzzqdJ2BfBCV5ip121fgi9BsbM32zYaRHPbJY2
i4Go0CcXakS75Kp8uKIKIl4R6tMnAN8YPsp6TltN59T1uHXnZ+qsh8jEVjst3BRgM2tyqfNkd3fX
Oq6FgQIhDUrKxyxVt38O8sXs4pObLrmlNcB9og9LeYBuMQIDSu2McwM//9HlstrxqqRaTRzVFkyq
xRR1hI4uWVUfNklMXWOQl1yvx0YNuyl4kDcSyyeAZzI1+8Fu8SkGxAqAEZlmo+iZhz63yRsoHVfQ
igfve7FiRUYPKgFzA1rufmvr0lU6zcrmv9rxdCo0FZ1SOx2nxU2PL29HUVpp2W3NKBJNEK3r1VRu
KSndnwWLdycjPQ3vlZtjeAI++VpKU96J27Xs/i/LRiBDhQdhuJ1LvPG9gyIXaukbNnItBwRuqJFm
xABgE8Qzg6jJqX/AoUo681V5/IQHsKeJoCpAN2YpJRRQlBCPlz7j+9RlGmT1bYunBYy1UKWyKAsb
/TvJEqeG+a4LT/K6NVI4uFMwsvXvLsiW7yNojkKiq2PwjP0mbRKBR3CCNosw3gGUjMghz85t+4eV
b+KxGgAMYuqcLrre0WvnKayO4bNzMLmf2AjLZuax6Ev2OFGlUIOt4YdaodWjTMKEt6Jne2dyNYtA
eVW+szBiD4ex7z8lW4awwUtcyeFjTeZPtyAuVluAkxLVATa06msWqfUdeMqK7MiBM2OLEx4dT2r+
GZPyULoHHNLEsOCuiy/lnzWlRRjNqBkZc3xKWFRWMbusCMpEoTWT/NINaClygA2ZxQlYj/CxMU7P
w5SljRx4SCmTqKBxkI+Qlss1DFPT6JQT8QsVspr7PrxhYfF+QVqmdh91AgpLCr+cxCIgES9t0czO
o4cPYG84BQSKn8k2FMw4ujYaD3z52D3VseJuJHms3/59dnXMrejar8NwAjYN9HLVOMjkGHETxwYP
UO2HC/tVmOEmsy9kRHUCF0DX7njZHOPakf1a9ZCkWh5yv/g5aqu6FG3kXDWJoULDTZW/xOjsuxtx
U1fRvnSA2s8Q9j5LsbfiALrO+xPleFdtIiedlMjIH0a3WamhnCQINBDDDp5le5pUzKX2jf79nIgN
fgw2mYySjurXJl5apSNgejQK5PlMG4xszoK6v7zWcQtxps2RtWqGk5UBzWE297P00r0CjLKzJPiQ
i2gDjl6aI6kBrTzeFwNoox74BpmMjKpgI9twL0zVSXD8WBqFX0oYI+w+ls0Y6rZba39SeRZEw78D
L0HJl6m8g+ez1o6GicRXDMWy2XAxQa0Vk61pBAv7fsMNplm95hKb8wbiD0TBDyLRDD9aFdVa0dwa
itzy77Bpe2M4oCn55JkkJj/gPRgvOvQFq4XA5E2eItoyCmTWPUBGU55sxSCxjf3rKQJ+6NTaDPwF
Sl8TamNgFBX3aYE9OFggZfYp3hjO+kLrE5XY6WfmEy/wQwjyWp6xw4Z9tV8Fg5b4H83Dp29MRfSP
akzD3s2E7q7P5gMFM9/tLs4OX9+wQMpFTLCc4AOsXLFbKfr/0GQwF6A82y4XwfpgIVHAZRSo+ZJ2
nS212h65rlLK9ysk+x3ohLbTSaOLn2u/TbgPEQACsUCxY/ibTTaJA6mnfrjNZfcmxoF/frxGD3th
dHkAwDmT34i5c/rDGuuEoIgCYjMcHsxoogEbsVXq7wL8/iOFde5S8DyDFdPW6cEefikEZAGWbMzW
+O/cYSrbB+9b67D3aZNnsW1p50p6S6maiP0go0iyq0YV6d/ma/h0PxZBfm7yado2xOGoKVbTO+1D
GfFdZyEgGf6uvySVGF1czhI6YUGMKg6Lm5Y2KAZWpAhyFlg57fg++5B/2t9VlD8StwZqyAdIyVHv
TKZXT3szTkkN9Ff8Qbu6mhH2TWngITTxsUJGRomi9nNIevK0x8L1wibeLaIuieeqVKrh6DlyOWKz
mnhXJf3zouFC8/PLIkjhTyaowwgALHkw1ElvDQEmEydPg0Jhr4YhIR4x6iKTG2yDjD+oi4kuuP9V
mSnv/ghsxXr61i1071o8FgfO8cqPB8oJXP3APArcnN0Etp4+I0ekkGHbydEfurZxRmNoKvXwkG5w
TeRtyqDGqjmwl6Dhqj/8pyu+MFJzggYbBwrdX8leD/0zC/O/6uUI1l49JVBlWhb2+RqnHZGbKVJ9
yG8Th/ocJeNqrASYKxjHJhNykua0ZXxERuuIaoyaGsnXthKWWHGwYO/IdBqpMy6JLSZ4DVlSlIAG
JKGiIA5L3t6SDqQ2GFG9nfjm0/cxQp76mYp7JG9eUYT7sxPggVzipCTYyk90Croad39+lCZMPgeH
CbEm9HgGBNK1EU1dTqKEJxedE/qWD1iM4c0lU5HkQiWtjYhOaFCY677wd2jQBvtWP116t3SD7hqz
UfNII7FvcS7XAmr9jFv4YOKdVFHDZTYu8jE5c//1cHKRUoxxGi9trePlSH+/dMdWiOyXc3aoTlhd
F8VscrZeMygmU7B6J2NEJGYOH9yO8jtJK8KpYBwLunb/xOQdRfZbjTcPT8NUDWE9x7PyAtvWYv/t
Un2bWXzTtnsGvMzPPofVDc1JTEXF4hDAXsql6zSaR/wNWjvBVPPTYNS8og6qhJ1/KC8hm3lzkU9n
V5BMkiK5Rdbk8CsP/+8xL/n5TJtHHXUVwBnJ/zIZVMxT9SBQcdOEg3szuT3dbf2kYgpFuQ4ss18y
p1H4bw796eqIm7ahXLyhzQityO1NrbefCYlNcGJ2xyWuHB7bD2M/YzWcZvKGrY/FSartJuZCgd67
SYTD2M45Utmnpe8gyxUA/RnjCvNyOx+L5AFwtrdEA042f3jGtqcZ+zFCA28FZg838VO2nxCYhiH0
TvH6K8OFJNyIl27S4+bDp2EBIkGiLk2btOedOnnZk4nYqGwoqUzfxgBmLNzRx2Tg2gXmtW30LF/C
45qx5+l6257VOrkR3xAHY5SpRLQOXyHlfSNAAcyilHntEr8vlExThquVRciIhLeSNwNN+1Oe+GRD
XqbI5HpDj+7hCzw1Mq+L+FjM6Sw5+HJIOGmdJ7f8gwEsihyeM7oX/aBESeAD7jeFVswC7HCbQMEh
hSl+OIybJJZ2mIbd9Irkk5AwjHJMGiFWlzwwwpJF5D28V6guWVrr+8qcusBdSW1Q0luiZ+b2hH9e
j9KI65AzOOO5UtUR1SMG5hp2w64PNcBNZkucoP+pJqlFDUesw63i4hkDaEm2tUglRWRiLiG/ndwR
OSy9rGWNBoNf8O8fzJuJcan8K9B8YI8Ix/y8J7XogYsPRuGK0vlRG+drIwqDcKYDyr2E6TyqwDu9
m4TmPojqkfTgwd7szg/DZ+e5UvXHz8pJndHEaQwgpz0PF5CKHHnJRyD8O5kP2mrfPOQOJKToudgz
3+oVhAQ5Des1803vrCrDN9MNWu2mdOSVwnDchu91g0imAlEPB5nZgMjvIkcf8aiMv0fSvd+vjWBI
cj+WgtYBfuIKF+ERv4YidFIbqunEZgx+DNan43kxVxwdLmJwNXr3opAWAu0LdXG/zJvO2w5tMQaF
kaVpHHRUPFDjgvNSMx40SkGmIiqVOKeditsK1qZI5owlqLwNcqLlR6vw0+xs6dCAX3urxp8t8scQ
NyJTw3B2nAwruF5h3sO/NCxpoa782tLPVA7llC/1StQEcwGeFo2kGnFnpX5/IDND7aRZzm5urErw
jmrJC33XTiwjM7UrMcGj39X7x4FO9V4qkTTLoEw3G7mgIskmu1O3g4HnX9sHRDEKRmIYnagxXA0R
XTCxAf0UhpMC70jX+pfdg6sl3O7KmH+i07ElDs3i6XtERmX42nNipLpVJ5Keax5afUrahwQq9Byv
7p5rN++PsQ0fo4GMGCxyhtxf3VdFRUctWZgbFd8jRdfjJoTJg3Zqw5wxEmVCjV0hYZYRWxIyoO6E
p4xhpXfLEQ1spGtqulID/DRWj1JyhQf8Mu6EXFHwvP6u8lLTf8GFf1IBnZOfyDMuJp2bXUr9qpPN
b17KzaZPNxUt0FoM1uS8+/Qo+No8xV4IYtbUj37tLqahqu2L0uhMKlr4k4VbqAdcieLKdOZ27Z4x
h0wDWhuXkjjz1uXVMzbpBBEBsp4La14DOwD5ahpnQqTt3m3cYMJoqNys/XgfATNYbVpp6lyqnFFp
IPJtViKH2PZDF6Wm02QmyxaO6s2HZij/UAflWLNg1i4Ar2pCfkrhreE7C1uzaSZSF/8fVqOq0Gcy
5L8nSbZVk95k6f1fMfykoAviNuPsNKo+W3f+DX5QJCzkZgFQ54YmwJfGUZ/ZTYgOKvzYVayrOJQo
z2HA/vFhpDPw3Ld9WceWd5NYmJ/ilQjSqJ81rCsmzNKH+bA9ZfBDLM90Qa256NnJvIuBcfeeh6mS
KaArJPLnBk/RbNM+a7b5k6/4Aho0y0b994hTdYZhiv7M/+abrQsWApcOirYMAFth3GaKkKwYPCAQ
HQZMpA6mPHHu9k71zLK/vc4ILUwO1eE6H1fxi9JTmXT1xt5lqSG4u6PtV3MJywagWdLupwmrzCyu
fpn8GV1bc2MtRtWK2x9hF403eZXOGN8lo/q9/8iCm5HzCvwH6hZHeMwS7aYLF5ZULW5AygenexLm
Zh7iA3YPZXfkk6oGM9D8pQwUjEXYE97yMRGwiJM/u7q7M0I3q9fhpPvP2HIdfeC9uKXQhYtvrrwk
XCLTMdZRS05tN/E0zV4mkQ5j1xS+tpKU/o7S9BI53AE33inyRCqz1lpfNfLCy34ty+7Neq/sDuc0
BYQIa4m3WZGsfaqeiJRK/gP3HOBXEyIg7BHdOBsS0ryS5UdrzkUFair1zCCwQj+G6tpL/JrEuat9
qmI3r6Fs67I3TRTXFw6IknNEFXibuoL8yz+JmGJi+90wubpQblqpnwt5SUGToa0oXeAWfLbzbkee
KzdsfQdb5RqkC6LRI5Sgzip/Tm/iWZL0VOEJRRHAKqZA5ATrC+4L8yD5qYOt6kXQDC7PaQPgkGeU
w0znUxACvrITy1mZfQkn/Z9DgDLusCdR7+yJwutAbY6EGztSjJcTYTs4wG5LRnJo/3/Ffpt0+TmM
KAF1zK3MJ17yN/Cv2Z9FA6yxxyUJtcrDQSOZs0NGXgRRxUhT5VG9eWpkXBTXkwz0AsBIaHAv6oWV
XAYcsa2rMxjAFE7h6UL+mnPJ76Cvqmbp2tSc/IY1ZJegla4JlxcKnen+zRB9HFJ9OTjtQZUXVXSs
Q4KDuV4WuzpcUqFQnvy9Yp4wYCeJySPQm/SpZnCSq7zsBI6JjvA6CP1q7mFD1b6On1tKqw4NornW
vCA4IhHBItGpt8qF+Dlvq+9ZT5kMFz6DQi+BCcbUKsw6ThM1nNHQJMd5w+ax7GMD1gaquC2MzPaS
il8U1PyS80GUr4Ms2tLN51q4GmT2u1v89AyeYESgJSMeDjD3LbecNHYozSxd8IAANUZyd1Ju75HB
TmTk4OTHn7doA91j53otiV9QCIhR9dcTesYrhEn7irIqKo0ygkl9kYxt1bNyb/SQhOdp8oErxXeK
bee4pcPn8+YyQt6bCiJ7cdpKLapTtzwWm2kAnRSNEAs89hjgWzTRKLlbPq1NFXJSMfj+xC17YtmI
yBAnu0Ej/zmGtF7dT5znJEeOoi+9P6G/+n6gO/cN4raKEgE/wvwkugmztBny8qDGvBaJmVSN9GpZ
m/pSz7Pf9ERElR4+GWkAZQKpQdXwnCc1iEqomiLyEf3BJgZOrqapuHAPe5Jftz0wlgpbj+5gG8nH
G/2Z0WpOItfij4skyuu8Bn6IWDELtGJrQsmPwgKbI9i5WPGH70yRkWrk+V1qerDSQECAawrlo7Nz
IWPiMzx4TILeIOH1FaLlssOl3rONKncoiNMF0ttSEkaZlvxXGqKSrMO/t9t9iQKOg3/2vefqSgS5
U6G8FtiWDp5g5fo551GBqfJjVAepLUu1X77roXA5NAUVnsWkQrqVMjhsCky1AOVEwljp6akVPtxv
wynFfHr2XdDfgzTNaV+fJQw11EQuW7nE4iG39XhF+8U0FDIU/50xqupxEldPfFe7uiPBKpDbsM/P
+hSS1h44Ht1xiPLOYpANe4tQ6Qfv+/HIkjfZ5OZF+YDsSLHnQXbllfRv3+cYb6KL0yacRn0D5L9b
IOGZre4jpgv8vFHlwaxFDk6Ms+vwwGhp+tXAOcCUSVmcQQztWB8PyYAchXU2DxwTx+V3smNRcrlu
VmaeWSnOh72qW6ctHrHrlONARi4WIpoP+OjLoR0kQFSxF8U/OvALtM8KoFgK9t1btL/FzbtfjwbC
ssonQ7G/bqI9K988CiPgu2WMDz881zRVZMSIhOChwdKUy6D9e6FXl/S1FguEq5QuMFI8tiBkiCb2
ljMgeCqMLtIp0LN4Tazx7G9K0kn3hOHJb4hMjiN/GEba7fQ3RPYIc9PMoXGlcfLgWLqkXRZZ2DXF
NvH8i6x0hMMomiQV9XCv1P8y7adWsWiV5MjoB17lU2Vjom6KI5PLWDZfY78O3e6YhGYEViOvxf0U
n5bOEamyfdvyZmujTRNNgyRn6GPJyvKTVt1E/Qj+hFUA5UCvhzfyKMMzUaGUsfAHLP4EDGox22UG
inWHNl0bD4p2oWkoe7Z7Pu8hgsKadLXiDn5G+7zq7LWxWnCm5WMcvAERMWIy2SJ4mMry7XKnbiep
tH/1Nic6jzWIjsQwFO7nww5NE4orFKLrClt7ryUu6QOj6O8G0eeXNclOKRWbZv7FYvcNldwE4iek
H0JtojStElPXLIZvcEmSZv3qFnf6w4PbTJEnAO95CwOgYULFuvXgL0Ofn7lIO0ozUfb2+ol4cmF7
uIt3jQMvUVyKJtK+u7Nfzqauh2mmKKXnlLW/qjpSxNCRhmmotZoHQVbXRlINynQK4HzbpTKRqHZc
3xr3JebLEFeHlN/LC2OydG/obXy5twXo1OUMMjSWArIQ7F/0oh6h4qXyMof1a7nn1hZfZVxE32jG
ZPPvp0h6L1n/Yultrf/LwPPk6/1shmPlxmS9r6D13ZlVe+UzCEio6B8MAoWJ8hpHzrZqtAKsSTY1
EztVatgVR/ixFYhutjEqvbpowkrh41buEKL03qxzzNTwJ/9wSzF72Lmw+k2wCeLcG9l2f2vxBZQK
3elIu5QYTw80KveRMiTQ1WjtO42DfXc+EM3StKkLixdlgTq7pHFMXQ38MO66ROZIbS9WqsSMeIaC
XY5+rVLzawtJfsZSw3pRy8t12oHfKE+JWHdlQ0qu+OgRBy5ungXJvOq5AIaXuht83Kfa37npoUss
0f7MGh5gwdBvAooxyGSSd/2OZGLw+lq5l6qJxeIlv5K9TaQD/viaRgOjHaGhWn/AVuVpmszgckZr
qOUh9vlKEt2m39boX72P8q6Ql+fAXCoC5iizDWbT0SJAWKas2YxmxiNKU6SyQchx973Om0s7PssM
Vu3MfbD606eU/CRyXlLz55TdzYynbNC3+h7jbxxai3VJpBqzatIdRH5k5uCCUSVAtrDf0rXejnvm
Ibe/RDWmXTpIAGMUDKqyMivNCHSrKbs8VbRhaOhPKNBYUAh24oiwwbBV5VD7lnuC53O9ZF6kDugL
n5EwdSj2KvmXMuCDqhl0jo1xZLXizGXnkUUPAb8mgA3DjCvDp+K83s2Rd8QclMGwLj9V5DQc+OPN
6DN1Oa5mYPH3WTUBb3cOAqI7ximjG44IJr8L5MdoQZnFqzLSMcaMzafNl+8UycRuYCJLs6LK+os6
ZE8f1kl3x+lUOs6XlW2kKz2X1ayKX84NKpBJfhMm3Jp4FLisKpk3pbDEC4YFtAK+PxJ/ggj4Enli
ie/2O5shrUeAhYu0KSyU1GMzu2kvkOnFHTevwXU/YAyqBpOVeFd5FLFkjfzPkL/uGVaSER4hsauh
mbX/7gAYtmzQeU8jDGcCbbToMkDwE9/PpbDGGRccYLEZFgNPGE+SaVMvpuuTY6TZD6nwBgXN+wW/
FCyl2iYXq/b5+oow6lhakoJL+MLpEzlNsiDW7cB1YcsVflj1NryI2+oZIIB4iCePtQLvGQE0GW7b
4NFRBq7XWa4sz26CH6mfyTKwvuyiTIDvvtQPQDtw65tkVZf61ZMAIg2Frtt3GJgU5XWDwIBxHvk0
7TpZmGT6ElSO6leSqzfoHZIdwbBF+9Qp9+v/XsXZpm49Vn1DDNPPevVD8dnR9JQY+fpqwp/RCQSI
qNAAw3v/qDtn4NT53E7vQ0C894Gs15AdH+q/M4Kr2yu7u0zvbZJsPro7s93tVveEo256FCr6NRZx
WicKgNkAuIISRcQ48MXxBu4umNaV3ifMAVOCig3kbfdiroPciFtJioaIEQDHyIgZFItQOPJ9iS3f
onDT64U/E1htW7EMfwaXRBJ9Nsf3nKIbiZ1LYDuN3MpUU1DWWNKMHfVmPQwPxt63xbGitt44Vvqe
E6t63acevDUl7K+WxLFNN+lDv0D1vbB1nTfjj5akbg3Ws+ZJRffXXCWctFTQLpWdfWWr5q2twsBu
IDyHkFoKadl0Nnso9Nr84f3ly8CN+su9mEPgWZPOCWAqf0f2pKEZqiCJbJCLxIerscQTGNJKHyXK
cNI98BZ0Ekyvl99H9C2aO7aqH9t9r0IDuIQnD1fbEA06tm7onO2iExm0kAgUQ/So1lFtLH8uHPjJ
s4A5aCsUce4tlek3GmiiR9ZX0pi62RKkYXQJtUNdo6nzRisyo1wnc5XoVHSt09uyGmCDlJf87p1w
5Eg2nOEeO+F2eTMilO9E1EkOGUTA74wv5HYZYUaZys95OJ+Jwt0uIu/cSUdvIKJstQBQ0onP9SmB
wMu5Hqj7eR3o00YEG+vefqF7//r51YsZywIV5RTVWUfDNLf4/17nlCHVDJMNCDYX9JTLMmvPL4Q6
WNb0rTzdDvKuPCxuXcS62RqO0GCSXOmnpo3AFtSYa777LW24onymmw0S2Cn2RVmpDVfBk3ez0K0J
zU8lamfKJUYAxNvBwSz9Ravq7N7t5LAm0rvUMEoQM0EWIi+dWtvmoOEJr+/hYLji/EExU9kCbqaa
9LlnvCEd6MkDQeLrF0+wbp9GfPsOq6EGHjL6Hs2WVt7rVVBS572k0DBNa32oldSqGLMHR3raanKa
A1uQTUuFC7Bo0G1kWX3fcv/Xf/ZcqHkasMNrfpSyI5Nyu8fD0XjFFQlnIMPo4fSsvjIfChifO9S3
s4BmIQCzjoYNUDbuSD7tu63NIU3FTAxAY95SN5VLCeMaF4oHW9sbKuVGNU5IjoKjz4Dl9tOC1Dsp
+kxet31grABT0qUdXrT80cLPrF3JsuPigjz1ADqkAhElOeCjsL7T00oc8lW5uBIEpeg8kHuFw+JA
M8XsfoWOxFWb135qhFcrMxX3EkR2SGdDVlEf4LR/bOlUmvOTXyc00jrOCDpYDrH29RftzG3XGeAg
/xN6XxqOG76L7pyftp3WMxofbKhQNPaUmXXKrHUO/rLlW5L1oDIDnrLUxeqfBclbmlGMSohYFZ+a
6AL7EwEZge6UKT6h8D3SIZzrFb+JodwsMNj4p6brryH3YVhIX9ncwooGnzCIIUkpuVIvxmWSzr00
ZiC0kNOPKfF9asQoVpue8LY0E3S3Sl0coTftr1vCGL2jV6qm8cfDHiHVvCo9cLpWHSp6uszAKE3s
THxlRVHVUIcOvfYttQ5PUkp305rtar1gNGm6GT0SWz4JnOjOM37TSrwmfUFsOBmraAWJhSs/vv7j
Kfo0ODiE6Z8X1vCkSetqzHNvf9410KOP5jKZRerjKf99IzXoYskfIN+afgDuzZXIAB1KsYZt/zuD
HByfG7t34GmcBbFTMERqXZatdxjcXp/A+GvjZq0Pfl0dEigVKdhzHQj1U/uWnLVJggY1a/peJao5
BEnaEkqDfPHpoRE6MyI2hTnDF8G2k7E34eIoiuSqc84VEpq50zOoqM38Dr5WP92q8mhNE845MBWV
c5egOAqbavcg/uVfmsylnMd32nLNyT4sXS5TH3GkhJ2MOZO+Dqd+d9IX+OwudDZ/37fzjgwdDdMF
NfP09P52jdvSPA3YCwHdvy6kKm+lUSR3zgEGZTzhxqQp1cjSpaonqyiFcfB7crKRz+VRKoDlH4kU
uVazuWtflOFFsYrIpcsHRNGp0/TNbfQYUSGlq/JCoRt7keuwMpOKgbZCD9esFluDhDm19ZwcQygq
Mwslk7CxYzbzQrR9TSyYSHC5qMavrGV21Ft0OXh4LT+0EyNWwTIJYsyMy9XjddbTTcgDB1A1wntq
0yMc34+6kjXe0wemBPwAPxcsBH5Eu48Or2frd7WAlWBb7hUZJGLX2RW/NnXBMTRKLSQnhGH+6XW+
d8M7Vavl8dssmVrjukCuZkU08GG66NksNVcnr65Z4jK+rTUslwGLINOgIkDjQFZ7eEWD8nBra7LA
Wrpm0XlbxHrM2L4lJVIxKEWgE3V1X1U8vvv0iQ2NB1Fv/jxYVaRnxZqL02r8NWce3rt/4uTLnIxt
5hD4YYTOM2rFwqnl1v+0AjZe1D9ID3AEd8OhQmuSWJq/AjUsp8haTH0oC9NZXYYl8W8GcLw7x4T2
VtLlgcG7ywK36CDH8EKTwxN9tCm5gsGUIt30xlrQ0C9IL1sV7VKCqgSQmmnEnrttXRrh2zh1u03B
NCLM3N38IHdaTTPsmHQDHl4WLIfE7U64MVwbIkuAVMVkbvbpxeBdX2JbY4Et/zq8LQjgYSqrJD30
tCpwBwUPh/+sTvzwsJQhd/RAa2Up6A4TMkmqoyIG3/WGuJeHuoxahUmdo74E3BCQiH6qsNhij8IQ
2lOLU8OewS07mHRjKxg3OCTcmRiWdNbFOK274jyTuh4ICR969iAeclelcw6SmWaDSlGIfHNfkTn/
XEFqL3P5z5I1TM6YfyObrIackfhu9ADjJjaOC+bpnZFZUXJ4o2332WdzMDqMC+9HuVAC9Xjurzwa
xWa+ErAZ71+7VDRfBfJG4RfYKFoaddefAPohjkbWDnKkVIt+lOybK3VXyPFQeAAXFqkYPq+4vYKg
uI5Py/D4CRony3Z4ogi8MKRUvBRxSvgegudA1KeoXDHigxVHspgJMyYcJfnOWwZ1TB8Ema5JHlkt
T00CixJ/1OnQzEgMpbTYSFuyr8B0FxjjD//ZURMJxenvINlohWwdOG81LWJ0XuAHJc69trsyIO/i
f4jY3WPtyUE/l3jU06w09uP4h/rNaBb0b6/fdC+YeXIDqlMzq2b/kvM6CdyZ630u20VQ7u7Zodkp
jHoE22QHeV5IpPx7Bfo5CvnYog3yahXS0zCJBtkthavDpg11l3+Mm8yyZO3LicmBW31W6uSu2rT0
DOb24kBtqpLC/eBY8LKA2PRjp0abEj0CXVI8ULfEQnG8dBVRAKbFwRbYWxyCmDx0dScFlVBQ04hu
O2bBdwWEviB8BDUOAlZ4cQ2R2MRWqhhz/qwoYzyiygervQNBNyDJzrFySviSlJBES+YNmwLq+XQc
EIN5ZFn2ILfJB0D0A94ftXNnFWLfCQ5OBqS2UXrHYgM1e0p5i+VM96adJ2V2EO59xrheQSNiEmON
/KitB4ypOQTVweNVsxEb6O90xzYqfAUQRr+C6YfkzHHrD/lGH1XSX1D78ya2Wjaec+yapQB7NaxD
AQPDwOMh8FwbUIlupBGNER5j6wcMjz8A/+UYOp/tjkLaEZr5wf4kmzTh6TNjndtQ9RNn5ECY3pX6
ODQz3xU4m8QIkYxBZ8ksPNPpWTb7H88wruYp4hxGRuxJYJkOtsVT130VkX/Cl8UBkJ1IK7hP2FnR
8DOgBKXljrussFU1CB3MMKTSw59A3UKKHgQTX5QcFy9Bq5yW1GiFZqk9TiX8j6MwOX3hx734nIh6
Sao5tTTHyaQ2zU8PHf7eYuJh2oRT3MTItCwQWNfH2OfOrr2qP2KRIKqNE4TkiLfxmVpQbWahI/sG
rU2C15UybT5NcSch0DZ0nOu2Bxbjcs48mR8MNpa8lYIgA/UrdvEsLQDurHd25XL0j92M9PcP+sK4
a56f/hFQs1pdflVp50HGGYsia7a9CNG8777gG1CWpUZ91o+iWoXXrp+RXrdXuYkO6AUYYz28sgPs
5kpX3gA/qWvsnRMTPa6VS71HnQ3SGBXUuBrHecxUAcn3VOGTtvxjRWxF109B78k5dY76I2Czw3y6
NmMZsuUWnxoGAxhFLasgFsGCLPgP4PsoMG3W8sWxtC0ER9BVPNMo+h3QKSXikYHk4M/SE84C59Ks
kER8Nrhy5s8bkz28MnIMQuf/l8oMc4+SwXWX+N1MStDZ7xWT4ayuKc/DHxusUXQj4XFMBeSyMQ+Y
G7mHXq5APz/nZI6Q5n/bCLSxuHKVKTLpibWWzMrdFTcdpFUyh1+2eyENHnm7ay9WNeTOzxs8Nhbo
aeyNGeljxPw3Fp96u2Ooq358ZJvyMuKVmnfNX+W0KVMsRE9RKsvPsDnSHe+Oh/+LNkFf0w9W4CLs
8eBKi6YHzg8UyVH+tk50IcA2snHkzY5wKpLJTeFHMTyr6h3rowrbrUeBi7NZE8dd7UrezikSLDLO
ngqqCNj5yxqQgy2f23UrhD5loKi/h1oxhK5pXtbLvvfClSNofqS+Bq6TeYIPrjzkSZ0TYpOI0LFi
xkg6M5yPdtRspEMHTR++pBa3ISZV4keGwGo5jo2LMpMhVULpB+euenxdtmQb5Wg4k6n93czPbwNh
/VlLfLxV9zHPVhXk8tAvJNUEsxgmCHX1mwrymE+p6uI7SXzfKbgwKHhqEKcyFrSojwhm+Rz4ZQpG
+W3RonIXdvlMfGU0bEXugL0LKFzqvaWroMz+AS03l+q4TA1yBKzvIebSXrO7LqBqYgOdAStbczRd
c/STLOouRGREMj61JoiGZ8QHLGpV5W5n6ixUmnwpPRc8EpDwpS+zc6dkM90od9oLs7RLmqETptWs
Pjo7aWSxRRc3Ij//giZwgPB3CG2NZR7sFMo38aOwUdmOv107l599U6F/Snw4iqpnkLlH3fCvb5fo
V4Kgl61Wts394JJhT5tJzgZdqjcqfGUAf2gyUrdOtJIvSnYdN1A40KzhstdTeSyVilloPRqgVt0E
8Ju9mCUBNTXn6uhdnpix+AS5AEYiTh7GsIW73RKzu0Po/y0Wyd5y38vxQodJICnLzkou2iyReY4O
sg9VkUSvK6b4HQ6NPI8uZBvOFUqVHED7HbXNIIbS9hfQXj+d2F+V7XtXiopbW8Av+unYf2rnXXMX
0UOnSvzJ7sQnqBppLjzVG1K4ZcrUyNokO4Kh7Ed+Jduenfc7u/ZmuQrJvoaU+XRe+LjfmjRvgyby
iuNGoKMto+FRn9RgSelqfeEtckIg2M6wlzPf7SUbH5ijMZ7iruatTcrCxq2EJs7nntiOcIg9kew6
08h8npOegKRVpcEWJy/hDk0f6TmK+PAQdouu1aUYVPqQ9BzclyloG6aaJU60jLmoDnLaNa4Fqftm
sN+4i9KnVBjNt8/qnFUDM+1gtylgUYWIt2sF2iCdNrR64KV5b2eYy4XA4F4a4miOFrCdbBzPbNoM
EQ2mUcm+M5acj76MQqDzoVGGV447YZlZRzMGi1+yICbGNhJrQwDGke3yyMWV/GeBamFzfc+CZwBL
WR0oVh7dovNkeDPUEinoTHRVQzAy98YupqYiSdoAolQ5YXdqnKROYN4m/PEqwtC2Gj/NTlYWw+Ip
XIXNvQ36DQ6cuIeiLXjo6RDAqJuVlZfAsLM0Rkm0d7ZX3oWKRRMOr9suCHpMpx9d/DhUL/7TCE25
iDh3oqWHB8FBIh7CZxdRRLuV2WLMN5hGqjyxRdI6d8Bjvb0hFlwZ6DZYuw/4wK2LOrj2s2uVNfFP
YY3iNso1Qg37lf91oZn0rs8Ssur3d0duHEyjBmdIyPvgGleP69bFExm7DcELzAZMMh9TmqMc6j4p
HjKcUqrBdJgNEIR/pjgTLujGXIH4sOmlLCuRpDBQZTZjQ4UI4Eds/nb5OmyDxwx6kHW/85OU/ifj
MyKZJy8hLQFQGKkgEurKRDS4gT3eiY1GqzH+7aq/K/Ad6+KQ+WYTwxfDdUUQG/v1NksPizO5vOZr
0aoaRI7p8MbfVN/TrmsmGOyqtfyxxZd01qZwJNL/1twHlPqDZTkvAb4o5yUCaZfM/D6RZ+gwyWvP
WYwq0zd8Wlw/jTkmu4GdFHyOmkxfKgK1rtdENsGkYch3coPEFTL/V4XBwzIAgfqnuwpL6QqQg4RG
YWzO/DO0kCAhyunohsR170mo04V7DcITFlUxBYZ/NTSKLXMZYThi3uPqjszq0/JQoIeiSyLnc8At
fA3v7aN7zurP8LLxBi6JeQTS6Tclna05LvkAWpxsAvFXeDDAAiFCl+BAV/Iwy9U8UK6PumqrsjXj
ngTpaUKVzmuv599cUtgBJFqz9dGqFt//wKU/58nTeu6hMDJ3p7CnJKPa+ptfpE5SnQqbDW0aQpot
3eB1ENAfilAChajqA2K3mLaw58yGGFs3wy6qviHgnQcr3AxyiMY9VHzcSwjkxzsYHSeApG92Hrqx
fR1qzCNaemhCx0DAJIRSf+FRGD16ibn9lQsMXQdwG8YEKtFFurMTxIHd3xFFTvujYvrQiRF4sHw+
rW01KXSDN27GXIPzLssl7zup5hF+7ZyHLXlMWuPdA28fdC6g8rD9sf9nUBMYYwS+48NVA3jrVUXD
no5C6jsPKgPYam9ZGzYnsSGx/QAKcNnuqNlU8rJDTOIANrvCksHD2+ZblKB5plXxaPfYZjEIKN1E
YFc7+3VUKqyLtEBR+sx3GU/s1OQvsAaUwyKncx4gtUiiAGG3j0tJ3DzPgPKuaI0hw4omu9lbOB9A
TAmjx/iKFC8RrM9S0VFDUZUnUJEm2tdJdYgrR7yPNReiLVg7GqhZlwUCF7EHH9X4yf7y5z9fqIeY
aKYc7eeyvfBwP8E4J4Klq5lH6KWvXGqn7y6DEMIk/4cNXw/1J8Y0FXVS79eh0D+ZEV2310doNxo3
Q5GO6VH7N+OdUH3Zdc5AnMJvlv6kvYbLqFuUIDyovZyjrMB9cSc55kz6kQ+ZcmN1IH9qJy9fh8xO
SBS5BxEIeGcRhPT17AwbJ8xBI2/UpKa+Ka7DNji4E4McByOulkBua+0y5rIO9dld/vj89em5WM90
ySksJPhdPog2bKgJSgCAcKZEtrjX9w8jsujcDrXf6H4jVB5S/+7vt12ulIsMC+Wk/7/hTobGM6mL
pjvrrvlNRxRt4WgZKPSqehkTTodWk/wp8nDP37NtD+ZS10eftnA+VjalNmp4rgH93o1pADEKVszu
T8h7f6sLIPhupHSxgTr8uOKnbxiQLemu0Ecwj8NKehS7EuYNkLaAs3AGKn1XmCsjIot2jv0ahQAB
dTISRfuGS+OjTDNAH23RsAoYxk7KIcuyVxGadUmOSuwRzYXGGtKhwNhDwR3i2y4MF6tALEUrXJjx
nYuBA7YGW4psmnLGU9z/WmM8uf4EiYLIMWInPZ4fGVkunheQn5QepwNj+JiiepVpcDxAifI3ZPq+
7BC4d7aa0QrNLaH3KtARYjw7VjtaoQVPRIHQRyDvOYXcHRJVwzxTT1gwLFDfcIN4/nY9mb1o5XZg
vPRyIIguNihewz90LDsSJLc6zdIIxUGlK3heUrOCbRmZKkartvRq+91G9Sh2qXjX8TV06B+U1wYC
GVjPy75er8Rxua1gV/elwc2GGaEB90cUzB80ud90TNnah1jc3aDK5r4gcW5E0qqVbjTxcYOi3o4P
Vu1IfRv+qMFsatPFqC1zFesSTLJzgYISHhLBwEPonewsY5KpE+Vc7mRL8k0YwRSDdHVQLJD5sxh5
frdd8KqfD+d3aeyCcvs/gCK74ZMVy5ZRW1Zy63RQ1cDji64cXKn+BCGutBvv7ksxq2sPGVHR5OxH
+SBIU6r9vFTEf7BT9Zh7hcWoggB5cStiNTHRSfE/k3dm5xALkJng399FD5Gj2j6HabycURLNydPx
H9hsRURtBAk9Ik1DAK1Tr5p2KHQkYWSrc/OnvsXFwq8fSQQTWeBGwM9mtI/3EFM6N8R71v7IMiVb
zAfg90indp7ce5fis5W8vy4evYO+CO2EOf5HMzFY+hl/OUl9ap/GXmZEJsNU7VoZrXTqqUGm2gd7
WsdqK6gAKMhxSeFNatzscya3IkasyDn9IUmLqA6RpCLND2VbisjgfuUro5UyjttrEvAUTVdN+VGS
rXJwtw+j8ZyMSRqqUbmft2TkuXmauQKjHunDgF7I8H8Li9oJzvEMTdZ8mXWjm5ru9mSPLBcPtEVA
ZLb2HhGSYKgCCpexJDol/P/pEW/EeZGkd7HpjP06MohnR3iPETPSNaab3HsL3FRs8V9vdAoXnOR7
KMfLNSCvYtIBY8KNR7x0ih3cLxbC/tk2kDSD3ZZwT2EH7fR7Sc1+XxQQ8cUvWXGV5g/CgSPyD7R8
cz+2YgZYwqHmiSg6gFSRUOfRa5/w3wfHSfngDdK3YMVqxvU4QVDsEAjGnbz/Eahi6YtqUJ9OTgkA
whwqKIqRXK4099AFFD8ddQSh2QkMjiHbI6I0cdy8TsxBuKKAYheHMtPlSaAGRDuVFNNQjfc77dVQ
1JctLZF+ylKEU3kaFp5seV6tmWDstMZj1URPXgHvjVzQmble69fYmPnvfHg0/TCBjxbCw2SFRzTc
jzgptE3zgr2Xx0I0gqWEtpQyCP3br1HC99tSWpgL97VXXjZEqeechcShq5aM8hdJ9nFsNeTxRN9c
z1Awx8zrxTTzvCPiTNihWXJR0FK+hxrT6pfONPs8JeNdThQRDrJrl09/Df90vBPc/YvdntCDgwyC
KuQi9MlQKkhpyG93KWjFI9i+TYjLXUp+O4s0/RcLktvzlTFA0LgM0lZ1UGnAshD/44ZrkbvwAgHY
lHkU4pakZcPdtiHJBqUhLUmWp7nmB9Co++hgTMkKkQQqqjiExsD1EeZtsPR4t3i/qhAXZ+Dc8Dqy
fR5HXz1SSU3g07xEDWs9IcGw6zZUmVyEw4jetHWXxB3lpUroL9FaUk5pWqD0dmlJ8SRjGTWWHnii
5s/LCnTjHo7Smhxk7NhjQarK4VstVbbvUAm7ZCeP8zhY2UNTXa/bv1YD9hTlP5NO699cq9pih+CV
chgXLL8lLOUWTDLhK3QrmkOcujiUYdt25b+fnXwlxgizEWKh1RWbZExVJ+6roe+i4iCXX7q0ER0U
w5V0ftv0QXv15qIvGf/QnUwPT5G9GvqsOa7YnLVtfAN01oCPGDCPBpvzF9jIANicrNbqH1LuNU9o
inxELTC2M55NK2eJ3L0nYqPd7Z4rIzUvToQYjFyVyBf0LwhA5TupN6edInqhD01XpAgMLtMDoKYh
5kdz06FcOO1T1S31HIwL0rjkhuvgwqXEqBnCq7bK1GK+ZXApA4AJm+EUIoWgarq9IibC/72su34f
dLBlj/o6RVMQvG+4Y03xYx7oHtBI9n2zIxXKRlkTDi6qkuRR7eDF9amb8f/NFquZYu1qMVb9m4Q4
uc4iJujCF9cYetHXqwkrjvwgDBLsv9cYN951w3TbJXo4Od2vO4dcRfL0Tzq5HGHg1N3aUjlzsM5B
zsjAWMrw/nnqqiq6h0gMloMeEn8Da2uD5DRnpf0csmklsCXAuy9Sz5DPYr0OmcCh6lqZl48TduUL
oTWyit9hGY+moDW4BSgUrd0Q7+2VMvGC1QWIGR83PoKPU+LElPR9eHUb848w4pfHr0tQmb0UH+UN
MZ5nTpiod9Y4Dj0rcjL2f4NBpD6wv2oY7LYYmUlQuW6UC/dPQCZymtmgXCzden8t/eBTlFx/A5Ga
PELbpUhQEkvk6ExHyZl2Sz0T1A93sqDQ5paucCJMWnR44Jxo0WYuumLm81vE1tgIZuts/eeUEaGH
mru7Zjt2ZDHpmaYYdh92rvtL9Y62B95KlEeVw44THufqSnztn6oC5V09MWiwcZU6A/LA878Pf9lX
Um6xHiT/9UXEM/x9bjqLWg07kdg+Q84Kxbckk0UAVcSu2266UNfEj/hYJyMcP4doH00zan8BI2ow
vNST2pVVvisFtqNyl9wmrjoHyvF+qbxydUjEh2oZQjEFuORWyfEEwVzh3mx+XTEWX7L0qeaMIazU
4SV9LXsGhw+coOp1jykhVsGC6BUVUBYPkEezkTjFl6T83T783tc+Dptpi2N+u1tZkSQcYXv1ICof
r1eTCC2o82FzimT5XVTPgB//mtwUPXH1jcTP5yfJ0iv0JW2udmadZ+vHf7cQgTghIcCf/QiCXFqS
ylOz/kfpFDnRNnZm+X4EwgX9kE9N52pp+0pZmDnCT7zkK5m2QBdl58Q1KMdIU8yvJRUIzgbSsG99
3yXAhyhG/NsmWHXUY8BLD9Vwy/HaowW8wWhDdtzSsOT+ivPiKsclWqEwWKAoBMRD+VIYGAczYBXV
UoDkqcJaE+w1ftBOUhI9Y8JJqz/H5Ix1pXKkShdK0zDD1jORpznvAcHB1Y1//m7iRm3RKpAvzn5Y
C+kUUqTkB6UfLHUsGq+LEht/0MVYuJMaWJy42VUj6FXmJUhIZZIKz+BesLFOD9vp4wQq7asZlmEg
3uniCnH58UdxZ+RfdL/WZRR5Ex/EZzstdPCD9jT89VIfrOAtmrBaHBwuRrRgRdfM7+o+5/oetrX9
/L4SDdV+eQOL5zOEr6HSlh3SEMVL53vpJ/XLuD+Zx8BULziA8/iRjY1oxDDL5evyea/8hxkEASsO
M60C7HuqNCG+x9HGMpK+fXvMM/cPuwXGPjm5oLM/X+bkqea2krkyHaEaN3YB97sOzxbOh6wg1P16
g4zf1gsuXQf7QeCdlUeLc6Hi0nLV9pJGfNKoAVvD2/nWMOha8HZxXSFxQEshOb7F/+ZIfiw4U6gP
eihC9ljNXJfpPBpSFqPpI9EgH+/cihFaFSu2iAdjveTr3p++x2H0Ffn3Svw+W2pAYElFGwjVfbgW
4i1k4Tob586NWPZcdWhNz9srZzs2piTahSUxvi6ucnI+mKzyJXnt3z2SJDGzzuzE0WVQ92rXJNzU
EOhTLYhwLtKUzWpJh67silSuSjI2cGEpbwPF2jwHRSQskgYvdRDYQtNJqCmRv+DZ0Jucl2ZJIbXc
BCCreDZDAm07gRzG7XUskD7ww0KOQHiEkt7KyJU/JNwd9r36jtPHlPNj/5zKm2IfdzBy9UirkFFJ
JOH6fGwvzjUfpNqBM8auW6poVYVobmv7tNIptMI1+/8akG0uhmqqPkVAX+wfCvRVztt/OXzTBDdF
WM4E4Mg2reb1buIvt/2LvzaPUa6gEc2u6wqQekMKAKoCzktnxw8zcE6Kkkj7UW/K/X+HMsX8fHGs
ojiO2iWighLiL68TubL3jshj2cFnaYg1Kf0XW9GBjOMZNwihSwq50+dyrwKnMiFwMa9xzI+bomTT
uMfCqx5/QC9qcFPhIHR6hsmCbzxe/6KQjaPZFB5KPDNda/J1kqKb+PkfleA+gjMD9lpcV+l9Mywm
bzrURbIxO3B5yTAzXvkRuC2JFBDd6VWk1mRtYCsVw+9pWPRMzB4R2S2YOVnplcbiJewes4rxHyMx
QOUlcr71lsRkrMrMeMzWVy2k1vt0x/hs6V6vI21RcHhgdCGVe+c6wAt3oX3HlqiIfCwrz57uNRlC
B+QpnJ2iTHhZCS9K6kdAg7Wty0b08W9XiejZQ9QH3/sUKbkioBNDD7TPRMUg3F3VwJjWSkBFyLNd
1WCYmNe00dN9oOFVC4oWbOXCA8rI4d3iJdP+U6lfmU37RCHkOpyMRLeWlwuQEg1qeBkXHgcbPj4N
2j53dzIe08SIaIche34g8YGLoeZRT40jdkhIfQXHpyNlherGXXYlSgPSDhUwE/TGv7uR85VpMqyz
x5G4ktXE234SH2S8N6GWOaLG9y56H0l+PP8XTr2EudZun4StuzheA9d1bh+3q8m5xKjj4jsWghPB
ZSi3QabvJ4wJhOSvoYcqNgnfH0mmAn4Y0udmSK723U8JLDYBjBo1kBM00dAPwinT0MR5dBCdig2y
3Q5mYfsMAOogqEpEvuMsYnoZKNTPY3HaE31/T/+Q11yLbAt6RkoBdLirKnhqm765aYlDYm4/Kcg1
NDNYBAIn8iLOpHBO61FbTqOge+4bqr0Qw/Ae5/mm7GdJl4feFUsx4l5S3quhGhgc54dHPNHf5INA
PpaJlRfZGlHSq8/Y6VJ0Eaoqndom79JCf18v/fXL6H3jJ4jIPxk6AK6epZOnMVb+qQIZIofi22Du
pSpwbVCHGMlpHX0ungUj4ZSF9XjUdfpYkRXZhl6ziI21v/oLk70xRFx5MIYGsYDWUBaYlW0xsD6F
FzENiy3ei72Nn9IzlaS35hy1KoRCu04JdhVsBggrGrwVM6KRdxyeY4gDGg5VRD/ydJ57jX0a7Y//
4ihBj3375xjEosJxnWRi7yqQ6m47ztS7jGn+jpAb1g1r4ZSbPXRCZHrxggm6rfu76KCn15Ee7aeD
QLwCkntpBW4lOcgDGgusXIMBXvuY7ByIa13fldHFUOwbfi7lfailFDFl+7eJQdv+FO37kZ90a2xP
/10biq90rSfIIb/f+2o/zg63/beyUlwKp35f0QdhzC8HwTvwr2idf4Jzyzgb10WKGAXj0luaHEw2
36RBBqgR5nSkSf79KRnhVfoudzRQfRINynQX2kmUZYdbAjQPnE7HYlBA1HVhvU1TJKStoVVQR/b4
3HjIKGg8caB0xisETJw5zAu3/DhKpVTszp92Ni9i5Du3JwcSw5sDWfZNgbXZ7Rm/+x15nrzOZK4C
0LhTxqG/kGly1k1blWQdKarNCxPxvPB7nZDBMIDthHVdqzw/DafFP3B9A0Q2l2hamRrKPi/EbyjL
k6vwLw893f+aXRGrV4hMlAZ9qCxbRyViOjgXaiEM5/ZnwGTXEvk213rxbK5DFoLRK48DqYo7J+B5
mm3QiNMBVE0HkSIvwr06T+sj/C3DLGr3gG+UbXDFXJ/oS2SjNbclGIZ1UdlPMbRCx45dSyICyj6F
yHCR2BBaZDCWX4k13fgf/NSvi9VCJUP8vEOY0sXeUdYP1NoFkuBJSK273DuMZuVdt2WFnk5FaHxY
E5MTo2jKV5lC3Pa3kASOalLLM+tYyp3SHW1GYUn+qDno8hedU0gXaSYWDkOAAorL3IZxu2QfLZDx
Sg0k75P18OK80csT9KLUitSTBcjywOpwHT+s4Ty9Jybf4CF1NniZZ4aqwk3SodLU6sNMo4jkKSpF
iaYoIFBjvx47GaryOcOhZ2zWDNdgwYWjh6We8zr1doY9u3cr5rRfXPT6YOf8uOs2TWtUJ8LTyner
4TcK7F3WSVlCAbOpZHzJHOziVwnMurft2IPWBp8LJAA9VYj7bCd1Hw5iqQdq/qTSz9GUW6vx4I78
P5DKaeyk36EI9IaUqptvkE7xc7oI2w+Gn5OE+ypXk2TxFddCyjmmxaHPKE9MVX0ZCcPGT+cWb4bu
9Gw8I7A2z3YBk1lJ4xDJBToC7Eo31M/lJoL3g/uTD+kF7OjgThGcuxdLhhBpiTCrBrX12WXXPiUB
Zpnc9t09iMhiyZgqwqxW0m8uARITfkdyv3uRN3IKAs+YriipJnPeygq10cqGv1RePKQDmZ068er8
ZPDvksmvrNaZd8/i9vrJnlqQZmPJQWvLVuyTdeH/0otwdn6ZJF4cIMd1xZ9UGki9/3bzmpCFs8DO
KLOhmnPVFQTCXdtLiqXli9V6WDwZybdQ2GZDvvmdwx9sllKEHAc2cSb1P+hwE8a03q+5eqqwaw5+
2plP79SAg0EKHy0YwMCWW/co/f2NU+TGClUD4p54ZdmD/CMnWDplza9Ibn2JdJ8UySCoL4P0vAXY
3UERk4UMsYoCVG0TBN7LzMMLfq+2py/wHMJc9BnnyEDyfII7TLfG9gS006+cT6JlsLb24goeKCTU
kXHDH/jHfl+8C/lvpw2Leq16ZxokA342xYuQZWsnofvYJwosasvhajYUqgTPPQEqU2qI5/qEzmmq
nf9szjETIjFcw8FPPwR4/gd1uPmIGaCqRwrpRfg2mX7Z2mH1pbOKK/CRHNaUdJVM/2HG0eil3YBG
e4nNCBe1ufYNnOKMj+8qT3yAdrKY3xarqRLZrsVnsmZb6y+es9vLa9GJc1H+yUXCPAvJ9p+naZ2D
wzQLT91XpMA+jA0wNytxs/p6imQ1X3Gr7IHM88AtLVrdYYeGzuSB9s+YhHvh7dElfonDyEleZLvf
mqF4pDf3hQ9gneGEeCbYKwFibxBdw9AGZ2Z1YQR1CVTGmJFOVyJcpwddLIyjKhE3zoMYhGwGeH+t
jifIBPapeaxLnnMwmNLvZ7fWAUnCRVE6nzK+nhY+5+39PcI+ZxSHglNlrk9V/siDBbBmhyHs1gqK
mD/SUVdLp08C3Uytv2+7vh33P/N/sgjdO7nz1dLtPRNLnJKMTQGjegeFpzwOXl7VzjEbgHxEUN0q
hVIZuum6WIZnBtkBhmUpBiNrgbUvDPzSDjVEhGWJ1ZY/FXiH8FNpvBz9zvLFPLhR/IipJR0JAh4v
fRZWRq2wxNp6QaMsES7RSh93X7IZKthGFbYj+CoT+dHs9FYl+blac2ZyATcVmC3VyPblZIynyHH0
YVMFCAxWAvt9N0MlHyFTVNvF3iR4RM3RR9DEPvB3U/FrgyIuVGOwFhO2Y1OVDlSOrlcogqBvK0Ew
4xnA4+USuyMnF/jOe/82gPjQhpbTgVQizwWrrNjSc+OdtunXWc7fpUjeje47U5NpHUuvGdSnoIaT
eI55b5DFsvDuYHsS+6rCF62uiRdEpxzaMzPk2wI1xLkwaR1IEC0ArEA4q2eQA2lMFaiDvA5Zfi+H
/gHVg0+L6RziPQj7FTPVtnYkHOEU7Q226fbr5hEbjIciYJiWabsQMw5cv9zkvI/84P5ubo9q3qWA
r+flb0bvDf2sNJSRhceLgCILdRXtkrjJDw4SuNME+GB2usomTmyhVwmkPYxnDtXs4xj2xFzSTT7v
hMlT99YHC8jKTmuXfb6BYXIhfuzQcnUrMNCvhokcYIQiHURYaXK2l6YBaSCP9HU22DiwRek69AU2
MCMd3adrZ2yw59jUbgKNhjUj8WCo66tFWD6ABQHrde0MI2LFgW3o1zuN2A6PjH9HhFpc0e0+IdTu
JV20Hz14Ybl2Amyv8Pkt9mhYQ7rQ1wrkitLry201Ha50Fm+1wjJAZlNrGIt7pPRZA7OdKQoalb/U
F+tVvkmBLdErw0sBglaSG7WL20ZQZN4Yx0k7X30TvSs+dVqWoft36EnFUT84QiZRatAgstJ5g8Va
zLLjY3zrfuU6esaKAJrJiAovldzqvVFfSJruNivmqWtO+m2+IR9DJpgFFst6P9eDRYMCFMhJvIni
vdBe6G+QnbCetIebUAiARzaxhV6B0tDqDyC5Pz1RxhNtDvObO4WIhkiOH8jFVgDRRFHN1oZSKP/a
TT2nRbm7iKNvh/1G6w8/hrRoh2b+DDI8kx3Eh13ekMlGbidJ9atjFDU+/dL5FBp0g6E/7D8GgA1g
wy/LSD2UDV06c/AHGTFDOdqC6SWEFCcsYtQOilk848CmiU9fLmSAnCVWp2QHzEfEI7zJYQKI1Rq/
iCE3alEWM7FwHMuXK8M5CjjmO5HefOVsCTCbkzMFiJJ9y0M1jVK4i7ajOkq6Wqn2fb9hFzDK+blu
29Hrr+DQxreJhdKUH/wqpM2D8A1ZMq/kRFLotbjOy7zQF1AWaFTtT75xgp3lQt83TLKpY79VBiaG
v1IfOSw9l8J8wXNx4agX1K2UNNtD04jKuyc6ePhgLEUO/gnAT9Q0WPa2D9ffbCi75FxRw7JzhXWx
6Vpen4c+w3pZ5dyMkT672M7MB0pow0bXoIIdhhLqJyyCGcjA5HZJqgA2S16a1rUvND2AB6dQd8pL
ZLGMOM423FyBB/UJLM8tmOdQOkvSI3rWIX9I/MaJ7P4qfsDtziEliOZPEfIOCU3/T3L+05tiYfwB
MQrcwLm10GmBZKpiqBgVVaIKt5P3QY/9hnVjEKPl6CNB/QwiH2byEvCzlUfzQEQ4fSVh1WfULogB
zQXAxnsk4Xf9sQYu2l7d5CITvFkyCTXdoL6v0PLyj9ocnFvpHwf06T63X2FmVZUQLvU8BxLxtmSr
tGArDRAslTd5gLiEs7IFNOMse7DmKQzqRQ6EIrmJpwg7hLMCunHAQybvrwJEoCkzRmh5B94lWYGG
fLQOIuqAAer/nbRQYM0kKJx0oOjo98V+Ehnd8jN7huyFbT2pLwjawa71nNd3d2RAtM6k4wTqNrNw
15+h/JJfmB2bsKfIgHT3vuGxaG19Q/ep+Pdfmm/46UcI9TkkT2p5o7ZfXOqkTXP0RJvc91dE6V07
t7sW/vX4JzY9b/E9fiQFccxDVb4NWaT39VOEIom+asTO8nhvlvM7QPkuGNH9QPxA3zxDwRrSTR06
u9qEYwj1M98zs9vjjqT5VNTkuyE/tGCq+ajEs1MKjPr9C4trlVRqyrRHbbYRsddBzNZG0axfDFPr
hge/mKhxUKRtmPkrKmP5DzUW/batxhpcRTFhk28mxbB2WZrWn5I8dOr21Yc9/8nVvjMDyjmw1ejo
XiXdC3l5QJ5cK9Hw3YGkuY8SJ1wuswfhbsWpX4re0TcXQOdeowTJHyZSHxs7skx+yrSNrM33dJAj
/U2Nld00KHIs2OH2TadXA7LsoOQ9BMdehnVgIQLJlckbCu60YJmuJ4KvD7DYRAsLeq1aTMAj8d4U
GP+ZKed2Q88yPFn09F0ToxgJX/86pd5hRtEeBoHyf+P5Uq2UBU9OLjPcD+LYQirY3NEfHtBrDFvj
uYKSqaxgqblFagpWLFu5rYlbm9kzAZurjwKbFBjdiCxaIRzfJ6Pu1HfC1dsXWkCipGL45Ht4uacV
a0nciuxxumw0usLxbv4NebAdRHrFc/4Wg5//9t6j97AD+5IhQbBwD6uujEpYCTCs03ZLv/ILYLYp
Q5rWqFb9h36kOcY/M/+IloDB+b//fcbHgFYYCUsaEE9tgbDRM420O+9mYzgG3hbGwD+edPO2yx8q
4pQbC4FgAkUoq3qqkN1XxwQs3I/gQ5rpyjIyonWhjpswl0qafn79m0FXyQchw47G0fKtZafZmy46
k28Sef+cDhIr4SXcg0kX8rIEz6xfrMGc5zdd45EuX5tVNtQIwo19syRkjZkWK6v/eahVNHOTGeV9
Z+D5f0suuXF71xBa52eIk65BvJg09r4yCQry96onrKWhzOfz/UH8uWO8pGgQls8j2cQVpewLRfOk
d8GIUZ+J0LsmJAiq70sMENiSxECRFmmpj3pnEF6qqFAQ98KTbYUyX/TdTOLWkOZ2IYADDpedGJyX
/ULdKsXaVixN7lzvlo96djduf6Fu7TxEiomLDBIla+fsLUa7JZLkdGcgpAZWetpc6lkMX1aHDYw+
D1qKILNyuMo1u6+llD3PWkMKmWCuZh8w3OtLx1VW6WbAVCtssn82Dtdlh1WtkeV4PMyUWBui65Ke
TvyLsT+qadGFhYYFPMiqMQj+BlgvO/kv+vplpyqoG5pFYENFsoprhonnhyQMq1FF8cK6DHRdPk/R
L8N6UAqZ4eKIywN6dsp5fPlNysiloeoZkeBix0S+QamtWKqxbfxsceAxHaw5TNr+5rKq8fjal1lZ
qZY+SuLPxSgN8kgr9ZqWCJfvUyINFBMRUGfCPymaiVyPWVL7ovcNjbLS3TD+IAKscPIFCUW11QAl
KHFW5NneK/S0NbkiXl5dJIU8nuwuni5NAgSyz2NC9ZcpNINewfARDBXB8RSB13za0FeG6GfRT8e2
vG+zh9pG+hKBt/0NllPb5uoSUuovNjxA50GHkWjrxIvNKB0AAX+jcIsrQW3ebcwFFdkL6jF1rcdV
qZ2jYHJ1ayWmYz4TUURgyONPQaC75SRp3hR3RZQwXRN7zSJMwLlVl65U7Hxzh3QiDEJBD0aLNYS0
0R3+/1Irkh9Ll6DCUlKf3UK/uYsEsoOUmmCUN9DLu+FapgD6AXYjlsE7B1rFYbb/hTxCtkCEWMaO
KVZk5NxvNnRQo8orbgCoWSQMCRVvShk5jjeoXxZeTmk4ZbBF9wEX006cCNcBLN3J8xxvgrqVg/cQ
7HPiBzck7ZNvsNnbd9eEzrhXssOS0wDvFhAU7AOT8o08XULbF+hyRSj0LrzpTnqf18E/1n1C2cU8
FG9PiurBJ14uspTLGsz6cM1a6avgjeeSZkwMWlfgZXl/skRXcTstd5cBEgouFd2MKD+HRPnQZv7J
doruAtG1RHO+XGNX3pZGCwXg2zOCgF31e7R+hv37xTNw/OUrWLadxmupyjz9YBTXrLfl7FPoOG1t
cbFCntvhhv1jFzOTMaFSvbbMm0/Y43fVZHsSOixWfP/CMt0Mod+nMgJR+Cun+QsjWc3Mm4O+g0ov
ZqYoVEwSvl0FLLsym90mFtPgjn2Af4BNmz35InpBsfVqzxcMZFsRmBaeT0+2Az9aAPfHPD40GDGt
G4OBOe+av05IEV9cu68xQGMmXbfWymbPCJp8MEcYu38GUOuzI82KBK/1a++gfC7hGI96rW8UySpX
qql+rIjTlWt3OKBzU3VdVJlg6ZMzkkCntwBrCo491fEgowidcnni5HoMMWDI7i8Sfq8Lkg2PpgXT
WFG5QiJZxluv9oxkOaLJhkZWdoaUSfQmdPY9IQdaBcCIW+hi4LsX+LghPf3ipk/vfySZF+YiGNfn
LMWjyFYyHuungwGo1VYCCVRfgNSldCPx/1zr1nfHy2aeYey487UD0974Xsfn9rJDzO2+zVb1PycG
B4ivNBTgTKNIWqvXhRuVNpoMTV5/LaZJq5rkcER5X6Nw3fN4GEzMbGXGCx7i272FQW76YLR15/8H
D8BTRowD1Pa8X/GJBQyY3nEHYY1nqzlrtN9RtuJ7euPGaEhMFJTD2r14J8L+d2wPwsYMVcf3Oi0P
bywXtJAnYBEW3SSTTgowdHMIa0NWWQ5pvLbta3R+SBnh6a0EC31RC+xMbNTJrbHWFU33Kn/O+ti8
JomHV9Wp0iP6Ddse4ukEwIcX4CI/6dyNdv+CTfO+olLZW+mbFNjxzdx9gDcCSvJMHmdV7eIRmCAE
qyPx2mqYAyDvXRxts+STDI84MBa10AeVyeTLjOOCvz38lvKs/U/4oIYwSBJLvtJ4/tnKcBFbry9G
Xkd3kS7sgWhox25LQHxqcZFQGxkdaiPJVKPsuoDHvAkIxda0b2km/eO5fCNOoBTiIA+f17c4ePrr
VduSNKxrgVnJx66OE8tNAgWtNKhnNcoMpBu13fHzizoHOPuy46vKE64t+cvCdrnoB46rLlxH3n7Z
g6wnWl3gQxZCetUGaTjXd07HXz90WlBblF4lBi82ayVrbhaCyxTqxZd7akvKVtIQkrZyWaKJ/3DV
05GyVFC8cVhFnynib0Ypew8hht+mmL7CFpPNJjm0HgiXq0c354FboZJzs1Sq0Bb7saQ3ql9NxIkw
j6BZvUyNCxE/cpcJUljFsgZGRJuhz4yD2JEtXz6uMXidssLxFJW7Ypkaqr1v5MAOmBaBrvnfWYlv
JhX1we32hmujDYgyKR2R3U16pHGSp6Ruj9XxxXATVjfQlC45+mqbSCzivfWQGXnkPPz0XJWeUkjQ
lBpIv2vJqEI1c9QUvFplxxGoEMrdSQA3eAL5d8gzxfQr/sbvcNe6LsQsFJiSa1BK9j3fndGeyspM
STYpwOnt/DddYbzhz8t89j6OtYSxQFTfcs5m4+cmSuiHvt/nAKuEFOtZMYgnbJAQMv+gSLujR5nP
vehyRvO0FLmJeJUK27kjZfxe3r0pvVEC/pr0zQ0QSSA7EwWuYWRLNqOSICYo71025Xs0tOPMSsDJ
jp8l2jSYs2EgxmpNtqtjI/5W2jxIom/sV8vt6R6HgfBCR+ZuW0t3PqvdbMnbJkdr9JcVEXlpBMvc
bw+FFbzqdAeDw1AVc3RvoqMZqagJ9VfQAQbGWjHFLLmoebY/vI5TeUfNELnl8Z/u5WftWwGoghXT
O1tmmQ5JgIdIYPTz357EAkxeutXsr/JkhNJq96o25fRpSOmZ2QnNkh/8kUeFTPLM8QsqIl0ELF3R
OK7B70tj/uExrdAbRz56XTeV5MYnv3CkvIJ5rNhUQlZn5Bdf/4v0LrLbX8KzTviP+4a5dLKQ5b+C
0fjhi+HmSA7No3+lLqMZItGEzPEY9hwMgMOuaMqDOXhnd3Ij50Uwa1pKApVHE1/3oD+2Ta3sYD5V
/0mPNSnQtkO91Ob2mkXkXkUEtCJdAtF8Yv75r59aSoWEGmoi0La/7K4byH1lrYLg+SbWXk9zn57c
+YwRkihAOK8+iWn3VOA4unusNbH16/4JAXgemEVR66U62zoxPc61mbzXu6FjE1xqHT2lYEmp3e9g
9cRguzTy4qdbN+hrLEIjMCNRVR8giUZ9RCqr6Os+bpJlkjWZxV7dZ9oV0vAwkkCYnL8ownldenFr
XEeoPDq+54NB0ZwTyPGpj/fJqxysIJMliuHUibz4iwkn5flMV2I6zPmmBKLUA8+8K0C/E9MDpkRn
7t3lSucNh9uUSfbLGRSgfK2+kW4dRkgZH0mLc62PIn5907u1TXNAl8DyjXWNXtCJxYWuBFrP7pNk
A9sa4Jn3NIoUCD2D5C+YVd55abmTHomxL3wa4+Dd2qofVl/TQgzK+X0tYQWrDMqznul1P0mcIi4g
APoJYqmo48oKrJU99gO0tl56rkI3C7LolAs9cqWO2dt1u0sF6V4uEwnmZIY9TADcmEmAcWB3jUHF
S5tXaE6Q41rYQwQ2oHBiaryjHgSswuPw29t3ZeC3cxYjylmO61k4ylsCKEBY1H8jLTgOpX0g7aXi
D27OC5bZoujag/LfF98L7ds9gh3j2OR9CuM8PVqOyMgDpp0UQ9z9Uhj2doMu8S65d8GvLbtsCVol
SEyzWDhZ74Nv+Vwg2J5xTMtUJmoM9qBdOkiBLZDUE1C9My40mt0zDK2OXXwHF+DuQiNdIpd8y6cp
G8j7DxFPYP7f6yK90gT6XZt4KEPuMVO3rCZ9GKbLy93kqFdiWT5ZevNiRyY732wKWJgEPdVDiOwc
5eQf3HzcOrSs/XXzX5cgb3yJ6/kGBtufIcUkHdgLbZKABcKDlbx/+yVstvil1zMZmxEYR+PAfEFC
UZvw776XAZ8JG8HhhF8jy8TCh+miVlkQqpZ5kXQ31dCeFqV3cu234OsAC0OAMHArrSvW1fEKK3vY
N1mDZ38IMSidogCdMwV0aThVKS6oLmzgLdDpvY9O30gJK/C70TEggXHAP6cFRL2nT9792geIjd14
koguT8vLlxyqxUoXZhPdVFfkomNrFdqMWGq9QOuNE3Bb3DmOhHbuezAFZaZ7UGv8tnoUlwXF3KCP
fcAH4KSTClcoPSe+XKtWmRg6I6tzTdeZ6uIpiGvBVlo5QY20szyWhNvKUkUTNvxFUKJN8OKVC6zH
VdngjV6Io6+bV5zkoC9jlYNzEC18vPs9ubO3C37TKpQ5mf6aFW0/S08ntUQwv/qXJWfoiK95noWC
zQtAYSbmWP78ejeZP5n4yFhAg75Se+h8/aPiF9vP5VMRuvoAytgOktOdXg0pTjGsPBLF4GVn/GxZ
An7bCaK9LB1e1jnFlx/GM6wIbzg69/gbDHzbJKRIOU/lWahrPDaJ5vKCUVry8+NZyK+XiMQxRXIy
spGp934nElZQQbINiFcQ6Mc55DYQdE3WmCwMRhO9RQaBDuJsHanrlaPKU628k+lWoQuZBx5wujZt
8D/2tYn+03q6XMfUSMfkLmEzWu/CaQNbnJauhsVbSeO7hbYESK6MwcwwrtyFeaF7QybCXGo487ur
dSn1DcxdWq8s0Y9PdTz5HFYnNoC2Ejl7c6/ZQmykZrmHgWiSt5L9WGo9Gcnl2bdvUvp2Ho6Tdpb4
rU05UEcFZldiKhg8TCKbmT84fnfkinkQu5OkR+zM2ZWCUWCGQV/6Mnf+y5dnMVeG4y5llFj1BKfC
QwD5YiU6KRkgVV6zARiBHzbbtXgYnwQvH/WZia8EHEPASu6ZxhdtBizBtTJHjB4QG7i5DFt5HM2q
WBLe9Q7MGMkUwrcuv8t1Ec8ImplLQXWIa46SDMUWPXlHi4rYfbbnH+vYJgY/inAsJoOPHeHoW26I
ftIJ7RHdfj6oBcoveChczAWr4nSuuYFaeXFSbAhCo+/bvYteUp4joneOJtnCvIniypZ04bCoco36
c+CJudM8gw7wY9YOM/+X43y8lIf68aWoRV0EKyW5ueT85lsC0gEqqKtfBguixZ65EbxQIDi/n0SB
VFq8ytEiYewNaYprnaM9ZknGOX3iIBuFCd5k/ew1+KHhpnrTk9xdceQGcqn/QqLRigbNFQDl+6XA
Qh6BM9vWk2dduJW0kd9PX/zvU2v8KF6uFtYaDeBZ05Ladb36/4hqdoPY0Ubq5M1XKVHl3ZSg8lw1
xKeor4IvUq2L/Fj2IriMJnD7t6yqEXWFhqNVlq0aEQwVEstFrWvsnj9omcLftD1uv8n2esKI5sWH
/Ta/o+lyTdQQyHBuJrnePkEgfIGDVK9LgI3xaIAUfyjnw4WiCRp2Lh+qtAGHUaFP0nJLkfLDMljN
nwHBV9somNTMAyIUaCGkOYkxj0TgK7+NfksvAEuMRY/GXsxMQRxtJUEg0C7j33YRgEALkl/dRheg
HQ1Z/+MVntIrWCJFb8hmnc3p6QCLOKT10E7M5kpfuQ3FvUJ8Bxi4G6Lt6eV72TrZ5V34r2qj2Zq/
OfqQxy8TfUpWXCr35S2NSHTpRAQASkXPWTeFz1sgxzA+TZ2gDj0L0e8Th5/KoMIjIWaakCR8gVKL
Xku9oYeoP310FMnLMQGfHltv0pr/jzsA/fjqrGQiZJ1tb/tWwotCNqgY5CbfJATJFCjO+XmJ1QfN
dkUhtmAPiJ/e/R5FqjfqBiHMgj2ZGsa4Ih5DB0gUY66QUL8C9Cu7c6bps/XQPHere752GvH3X64x
pS1oKhL/Vg5o4nGObLk2WECZQR74K1SKc2Qi2r7wRbPPECbR/+QAh2AFePfa1UJWGfHQ3WlsCFup
Kd9Umem8Mkfzrxgx5yp2/YMxu3X9Ces8s2BvuuYIhUrL4aaeZCBalCrY4VZKf6bsf8GZZav6W4gX
ArIvjKCKvkQyc9vqwT15IHKiGPRtCH05D/UzkZYyLCBc8oJpm0bBzWGm1wEm2yRFq+2fvWP8bp3f
WijEK91bljb3auyZlQ6Tkp/840RYT3um/t+j5MNdDuXGV+s9Xrs06E33FNF+HiapKfLEvEisfGVm
6NgNlh/b5jzQ+x/oI3yXDhCBTdh9q679+4OrMPSOIGLq44DY2lnFU0NS4puZjayFEimZtQFXa6pl
Awyp/cb2rYjYy5yDP/xvEqFeIOtAnSXK1tw/MByL/qHZSYU6xHI4r4rx8bCN0heJ6LqmLLhyV2LG
V8HM1jzgbipswHlRKyfPNiOamMpXNAIHRpfEApYFVDSG8bqmOr6II5vR2jYc9lJhN5yVsQHioFj5
63TyiYTTnpfZsZDdroTj3VrEZDlw8XZK0wIswcZhVHn0PjCW/xAMhUwu4ceE1DnO7so2QrxgLE4c
elFG8KUTqGtAoETuQXyXxwPhSlL13atMaY1lvQeSS6J/BKwhqLH27JJ7opvPqOB6LnqshqL0htMb
R0yR7aaD6UFP8BBQ3Rk3CF8CFEaD2JTAXzHBPC7ztRB447omBiurPfycZpodhPXyfqgFvobxjPUE
9KDz0RaDkfeSSNzSDERkStRfYHrPlQ30++ZhR9BwHnEWIDYVE+7RbYkLV8ReqlCNrR9LvJnRuzgm
sHBFH33SazUVA2lD4/U7aIRpDmg4mxCwBpNlRLAR0/4vP5eFsRmS0RvjU0sU9wLnBz2jepLlTSNU
ZgIPnVFHuJRKF9/4jM0jI/zHSvdR6UZTfjeB1hcxcorSyFVOJCJccCQ/A7fdR/SmL7C/DdbPYoNI
xfticfoSJpXwKWTUAnixi+k1iFagxfSNqUudT5KKqWqsZyFgrO7csIYkfT6PhZ4yNtJA+3Iz1SMY
5mgg+5O76Pfc+MnhmUXP/uNK9hfRRvBH3ixkdx6KAFAMAa+i8CJikWDgJziTnE8+1UO5hROTM7BM
bFs3zTs4iBruaJYNhtLsHTnga1GEIbWbMuxpC6qmXba4oGsmPm32TV6EzPl+KxmMsXPBgwZDccNk
cycmZmr+Kfa2Kc9aG78p09e3RgrfrBD1NnZpZ/TKpKM1OehGmScHeFOYHeZnFussqeRiBkrS/Kz6
MAzzapABDU+yudrdhBD8YLI/H6UDCnEbbprWgxHtXJZg7ruNP+sflZRWSG6pymUPBB8zNdK1zI4E
G0gJoA4460X2vaIw5eYKl24yTGPgMuHw1Pu1g95K8XppNu0ZZxpFtHEpq9WaG9LoYbMgelWy8cl6
TYQ6MF6S7Wrb6MJdKwY8LheNQsYOxjtS902A401buMiuukeNCoAB4UZdAcYGtt1zFRGNiNY+6Ybb
4qqNt4Fm7rqaDffNjU4jVoFkvNbY82HQOGJx9BYP5jsugnN+tRmOzUikpgKaa8VLRbG1C3F3yCRA
KVfwYPCVjh5/zQwRAPlxXTyC0krsq1puf5d1XF7bAkssMudxII6YodCmA8URaIMV/jV0xHZQ0nj6
50fMpS+dF1BYiOPzKI6e+T1g9S8XTCWRSC6TxuJj1LLo8S/09oACw5OEKVhcQ6BzdigoiBVi1PRH
phjfsPudfDeV2HxlOsYqYKfVB9AKfC54YiH4SuBPqiIQNav0Q/BQnlQwkSOJoFFftS6AOHhE2FkP
tLcYtAU3eGSWqT85mCZEkjUwdx94An427cyMty84dvIfxLLPXn9NN3BAdp8/9Qw0uQ130VAFWFbp
rOt0DQKdiaPDb0E02DfGtHjP3Rd4mgV6VrBYccnfsl7CCXocyKQ7puzY2TJU2zC7EAoGUAMsgSmt
Bz1qydx4idZHllRsmI+SnLJ/Bn5qAkkgj4mCAXjxCDtvqD8CStAaio8QSrEfFWwSE00cNkinycPr
BShJsTA/SgewH1mxdDmIC5jdyAsXTRXOnTTcbS0OzUIy/6jwhqacAbEP1Xo9EqAjncReOCMXRq03
V1iUZwD5dyeVXRRJevBkQg9V/KUm0Md8+JdCs/pXqC/4YjCX1qMljKOX+hs/8lEtOk5oktgdFXgy
34Ki/M02JihOC/zlNhGBtdhcH/MknLrfRUJGLYghnJ80CmIvm+K8cfExEgsBBK0yS3mgUDddEI6T
7hiD+ULfro28hPLACEeRHmXcf5TRzAu1oZm39kTmxfwkZHom+FtjGFa01/S6zcXUdXuznZ6hcTVg
lee5h1SpFpeBhs2gBz9jCY2+eq4yVIif5Y9phkQXFyNvjWXY0a5rW8MtFM7+WHiZ1fX+UelP57Eo
SeXjhB1TmZt8h3mLVLfoIigukrBFm4IfxuIrTOIjdTdhGXorofm7n7XlsAfzunw6LA4TlyOklU4C
L9giKKifJQDiIvHeTX4p+hu2lMewAbMFxnvIIxpF7R+LsNI3L5lloDbiOlEzF9rZlEMJ+FsrAbfh
6uduZvIUJxBtiWs+HJL6NaSdSr3yLwem5dj5IItXTWLfjI2URK80mndtqxUYW+oQ25W+nIjCzpYb
SA/Wg1SPXCw9UMD3f01ghtlmrNi8cvw0Pd+cLnhWEw5f/cKtqljjwXCX/KrB+gislR6prLz3bjYM
5n+fFSU/iiLXH7dinmc7iYz4OsPwCpVaFb4RFzK7FQHb9f3yeS+fajVWCBy5hnZwkG3eDMJCa/Od
Zev+fXqx0HQhdhgmfWWWIpnWj8YhQUe/Qp0aUPkBTFlNT+3T1sArbCkhSnOg9cRoApHD6UYMqvIj
pf2MTenYo4LiLlXE318Vy0gUnJHJb+tPEdWz2ND0TR/TUuo10u9f23wUbSW1IfJUjwOP4eEWFvs0
msIiy5l3wFrX/fWIeCbTJMO+FPUtcYaO/j9Q+hkGY/8/5xcDkyMJDXvB3gTZZZhluVaeKUPTES4R
dKs9BgwCXjuzCPOdckcsvt7my6q3azMtpwVlSLCKPyF7kGFeXeN5+RtoDSP5EdSeas4g8eDRsN3j
dhOOBa6sfgi8JlGLFjXc9HEWFYbLegWoUYv88RNzF3qPQxA3gJQyfH2ih+U+5eNG4ivYVcZwpdkd
QN3OKUju0nfzSEa2EBXFnsFSY8unbtOmUFKZHOQfT6tYnZx7RJVGBYTgcBnh/LPiU++rL2MtY6Eo
4NbXHPq019lvTavEV6zTCYoZ2BKE8cqPoBPW3jszbqAF53PWPbAqIwfLge3CpbWo6D1r6AwS3/n3
uc7KSh72mf/tykWGH+/zCG+/sk1SWw3/IrwALdcrVp/c916+4VTGTt+Y22hnBrlq6EEoFPter5r1
L1rsHVA+FLb2FaKERBywlzIkEqM6iI6OcESx/13YmsQhyd7I/ERMeVzd3Q/NmwxPvuryY6WbTIgP
3gmaZu+82tfHqc26MuXLaCmNbyrauT89SmbSukh09ITm4l/hyALqcIlTYTk/p8kVuzSXltAw/TEG
0GORenX5MYf5bZnmN3BCrpsmmB18WbfRL5sf9hy+Uj/ATJp/yKqYwhi1BysvXiEtXVxsw+M56KIj
VIBagcUIXA9Bbk+iObHacH4Y11nUHnjiVYEFAH3OijzImmMQKnulkS6lMB1iuw89AJFfbtOmvoXK
tQe6CgWS3mL56Zsa3QWb1LLXRpi49n8e901zpGNjC28suqj7H3fQiCc+UywcFwHOqXsX6nWLs6oU
cXr1Q3AE65/lyWgRloSspHPDxHYeJU/f5UfZjKKJLoO8f+51fpA21WNE/X4kQle3X0hy9Y4gq4Pl
vhx46jy1ozh72tYcOEYNJDEMPxXal44hpvy0CG9ObN1N1MxR+WstgtEYChf1nM+teZO8DIi8c1a+
xxf08hypJl2y6CsEa6/Fifp7hNaMaY1JyD8zj/urevycVaqf9m+eb4wKWrfWMK81MWR8iVizroIi
zK5CnQXR/uC96+ASgaspOvr++IGulgPg5iHRouNoARD2P5hcp8vlfPKrvYzakHro/4RmVKAVTFw+
fCnyEO+7lK5EoVM/OCfxN3F7Kwi/e6l+Eop024UW6exTM+2I5Im9dwaJx5/PQh4AlTPcpzfD70Yy
EfEch6fTo3hvChBHH5NHb+e7GwWLfioxXifTxF6FRmZDoxdmBwd+x6oz8JGRSvBZzg5Ho6wck/9p
HMvpGzC3Vin5b2Ix/21YxBA/qktNi3S+8pwSI9OIBOKoy7tihKfwhsWO5gwaV/KHUZAoUiwJzjKO
r1B6Y02Cwrq+BVG4qKX9tSHmEfCCaKsaC/0oWJKKkhQOr9EEXACZef+UsPlUFAYAX7kyEdLZH/Aj
P6T8Zuih5c8k7RCsuvLpkmz6bGEyQmLPgRLNQCa6Y4OJ3LDXDLR6OL9rqIkeWgQQtDYyO+zeWZw9
JcFhopv0jUE3RwYsGE55LpKvv0avWIwuOTv3MGnFQsiNbUYZum5tBlrvU8VXFYLHFc4YU5GbkARm
LX5iZHR/ksT+4ciaRpLYRWKU2BhJM33zMpjICNx3fIIwu2m8N3rPTILBx9lnnUQqmgmgqxKIIiaO
Ku8CpfaYHLy9g6zmIxho//2Kf4Om29MXXWspy6VbcWCoVHTwxtdX/oP3N3zIkTawjAU7Pl15sSfc
J/FftQRzXeCOEEZ/sa6aq8emCsqU58DsERCNSAn8VJMgdmTmZBp/bj6Uj4vyvOihR6ZNmrhuFoIf
pQ/Cd81gyw0Ix4uJj8UAQEdV0HrMwrNb+fzxvIrp3P7r8jiMRWYR80JvhFIglrhAfajmgHB5srn4
XLF/B/EGIDGOdEpLxU0KoTjaBJ31cZFQdd44LHjuC5oIw2qZax+ikAxlzKGVKzkoVbcgJDGq5Ldw
V6lFjS7x7QMOuuwS/z3Lr+f3J5BRYheClr7EmesTsFu+4bjRBqUAUdWFBfTHWMFfTqtvyCuX3QLy
Gf+c3lnbBV64SeZ2qt/whqZ1jbjDCTIUMg/giGYN/bTGSuZWyeoaNmf86tOhAppRiXDlzcZ0qD+H
JvU+s+ofNG+vF3vTbBnj+GTpPVWt6rBeA7/mG8yTY1rVC+4VdVBEB7+UOLn+qmPXw/2awLWnWm1C
alA9AnDJwRO2fBJCVIc/LEhC0yG8UtDKGLTwqkCHp1hTaX2WcdL2ZwX5jxxwO9S9FLu7r0FIKzSP
Il2mPYXSnWSSMcoiS9+XdVyFbHXexbZepFJ9XFwT1jmXtzbxfC50hbzW+yEJgfzipjBcpBlx7hU+
/j/1SRsPyQNdFS7i3W1DvLEDTs4tW7fN+poP9JWmUj7hffNsLGne7HHh1F0+pMkjAt04taGgbaTT
twIuzLFo7YPK9zA5BCspocA5ArP8uv+osw5dUBUoU++tqQkmTiR0bPB3Tkp/UTFZWOxUU67pudxa
nHToE+QAh5fhUuGNGF5kpAXXgLEoJiQrNIdU/WANSyDIiFxptiDIIXV69qjxlsH58/OwW/yTKnZa
qBkkfPCBYqU9H+gmT5nspJwbpMBHBue5WRXvVkknaPFnJy5HZQVvptGxrRm0aC1nvgybkc/4gZut
kGfDQs+ynMTndBZOsUskZ/zu81Hzp9J0I/l05J6MDNx0S5xYHo1q3ggBZ3ZjNSm0kZn3a9WuqiQH
OofL5lHmn/tLyHaPRxBar542yKIPWAoNW0uQqBvHLBCsu8jiDJuYqFLnjTaAC8sl2Slh8xQ7zqS0
z1+4P3VpbB7mW2JYzWYs1w/Rm2zjdCdbBYd9EtDenmqArhVC47z+5EpJnS7dfxrL/h1YR/3QRYCJ
pFSLIEgtnzpB9sq6juE3CYyyDd2G/dp34Bsgbsc0Z2jblJbXm5hxnuYJacAbBGa/JM3awMf0YR71
rhPhUVnZ2g1Aqp5an11o6xEjCm/ETcuD6bwlgHGMc7wmwL7SFUaGqr4P1K4r9HxDkBYGzU+SeGdm
oPe9+kaOvX8RlaAF3WqDi0oPyeIsGz8ARJx63tTiVHx5xInZ2RXCWcwajpz0KHmTbU3iBVaoMmqK
cHlfw3Vk3UHE7AMEOsEcCRmjhonGvH90HOA6W5MU8NoPqpildBXBH3/MiDLgmi+zKd4k0JiCiSDZ
HTcZEzzZ5NxK8aBb+zDr6NIdUR01xOWwj7vbIKTnO9yMYBRRwAMdVhu1oVwfpi8wJ4MLa73FJOoN
vPvw6fLY7ODc6DA5sKKhMnHyGzOeRSIwTLkUqNlXY1sU6XOOg6y9XpXtFJtLq4zKr69cAbKfB26c
Tnz0HWB7xyt17kq9xpcTx8R5qRy7SsdjSbVamgiu+SMqbWUs0OJLTEhfzRr4Oi5I1x5gkZcLEnoO
zeorrYCToOt0/gKnXTVvFhBiKgBuPuHig4iEeTMW807LjAU2EZ3yZk6SXFG7NtvIPMoG4HJj90ko
OZR6GxIQ/RAIaOrDJNIbVNDEFvulwLeb7Byv5og/OFTmZFE5PCdKuHIPqKEbyDWGlHU66rULrWTQ
FZzWaljkjn8jVk82sb5MPymNPLj23nDuTRi3TLrznBuOEmK0xSTz8OTjQM3vPGNaOrD4hOvEuBUL
Orxwr68nmnTtoTKcJI+cX9XK4+bLMMfBlFMsNL4g0fl48f1AtplN001SRz4lgpTr3g8G/Cq2bbG1
w/9pZXNZIu4LZJXHpytIXrjX28L08EPm33mLhw1JfCM/39y7H+j3UBq14/2E8LizzP6Env2r/oe9
bSC1yZooPQAKCl9BVwd4EgV8d7VNsk6J2CbPqVsWmQJDnz00RBTCvqfdPB4/vo7p6oK7Kci46Qzl
mY3Es8Srh+ge+1NEVK8kOVBzK8A7a7pVT/6wW4qrbAFLI9fldyNAJfb6LVUu9qD1XoSeoxPX1pzH
9xEB99kKBiZrKFzUqQQAdcp8CxBkjbUkiLgtVAR8WOG9FqcZGVS22WKTE/eR3DV7xsUdHazbf9V6
flGQUBKe5ri5giaVHh9Y3gNObS3DZlNmCcdKcogcJaHJq54+9yRYqVMS5etHctWiL71Hr6nnaLhY
iyXJXQ988UBCHaebSX1o8KgTe0hHgNTF8SVx7ngjRXKv+QgiFKtc7uxsw8lLZfvBF+9zmhB9fC5R
ZIKvfe7cZ/V9OGtOTiitnqSotTtgjG0lfjS0N8HcIMAtu0wTWkPSBtiSVRJTh20NlohoeIdoDLlz
FV+XnEHlmj+bdztO6LbWyf17cZ5xRl2faMN5Y/EwM6nQmKn5n3VAXfyxFsWwAWWEx5XxN9cUGagK
HvV5uV4zhaigdS6pZo4l0XnKyKGc5VkhfJc9G8RQHjGgEXTSx/64N96+VffZ5d3qoUnEPyRbJ33I
WBOj9DNNrpwcsj/WifeFo3bYiheIXWKPAo8889Z72rmvQtJ4cTDn++GQG4oT2p/OyUv8G3Wbs9X2
UNbYlZOP3i/7kv1rywhwb7fEoXfmTKHQTle4yTAXTGG/FbLE66PzaDp5z9AkQv1n+yfctY0F2bFC
AFV4endZ9dgwkCcFMPH6RfLtZibf0jKzjih5gwNQPIN+P+jRzSh0PCuulDx7Qu6ucfKDG+JrDqSj
8m3CJGxldBIVk+v6AiaMlpnrWlLfwl7F3KATDxzMv4EHyB9ZlzHrocE2yZ8w9sHitRavBFRhtfKW
cI5Qxu4UzrVi2e1LHeaImDNHpkiGeyYYDVmFBVaugSF5b4XsJDVbK7nXI1BWNe/uarQ6HX8oKxSl
BuYD0a9kWLpDy9TgHnGHsk4WBmm4+5ijx89ig7N1GL2A+gZ+9A2Vz6sD1u76uDDxuGO7e9XJRsTy
rg3j4wjRHn88ZzTOheRtRYRKnfLi3zp/ZwJvWm62AJjtizZpuVEB+JGtuMPt/uZEoGODTyXHnbKu
JFRpID62Ta11DWnT+pWd0yvC8mQ4vSOA7Px0DlSO/PWnwkpVFL/y7zJnBdEumGljPEJ964Il5BTR
yJ5BTI32W4wfBvtu9DoGrBVozaPRvpRqYLoHw71xswjktVlJH3p6mvrYvG/ieTICBWnkHykbAY8S
wQnJgxoUZbah/tiGaGDyHpKKVkhro2/wlTerXbK0FXbkk3o595S/gpOvQ4PezDb8yQMdQA2G/0oG
5Mcdw1/RCycn9leT6p+5Wg/Bk2187lUbKAb0Cx5RrKvtSZvT8aO6GTCFjyXdhlZ30GcwhSFzu0lm
tXrHN/qmIqmfhmn09gerRwfeowtmUSA0/BETX21vg//5f1nJ/7IdG9PciG3pH8PBn2SYS9aBX8yv
6IDEIn4I40QmMhh7ZKbnOLZORQHUQ45zeehRYN+GUOiCc9Tgc2fVQnG+nKvUr0NG6XcdWBbxhfFR
NXVqR3naZQiA/3dwvD7X7hgf0gGNm37nughP2gDLv2e9KjaDd1fExrcGTrGl4n8mY58j0GvzG2uq
QOJeYmdjX9V8yrRnRINN1B+icbaDIxLaJVUo1J4Q8lVelYhm+m7E9NLGRsm6yad/m6KBrwcJc3yX
14vocICARNs02KV3rtsp3g69wlU3ZS+rWt6g16CFGuzRRrlIUZ6PmDRwtgryJZvMXIi05I5eQlWl
GP5Rg3Y7obzNAayNGqHWCbvopfaJmEsmeM4dRJshG9OGvHV1WBcYd06Ln6w8MbB0HXFylnPDvlp9
/O/RRwSgCYw8h2DexqKgEvOo2LHKps7C7M2nJkOsi41wLOWH/KzLGXfEmXr2dGGtSLLB7Mz37hBA
NbIvo2xpVhAqblDXybWboRP4etkvcdO8SWXfN9lZ6drh49a2QI3lcniw01qIFUeMpg2YoFwfm0kH
HSfgQkTkgTv1v/WWjWQXuCuDSrtcKHUEUn2AMhNfe81AqApujnddL2wVS9buPziLoNVE3Y8hF2XL
OGVlLhwa5TqQxOKuYH5k6ealSzBEMQLnVbal+cc3U4QbWyklfh1QhZDHJVl6jsndm7t8uFEeGzAM
A+XSZq7j47LdV+fl3lVNWO+qq5GvqhU7VrXueYQFtNDTryRjwUJoTpwYlQhbDCcIxfCpPxShDS/e
s58O1ZFiXGEPJ1Vu6dUN3VXygvBx2QEsg/PtO9nzg+rKLKAVH3QZ4Wyhh1OkFAt3zwVm19CycZid
1zJbWc9bQrR5hRucxDz/dVnK+fTyg4lCFfd3qFDr+ExQIo5CTgOWPZbbnGvRovB5wf6pIETkyPnR
4yUiK57DooAnlBRyYpVfwQ6JjZtNqBNSljuKI5SwAc7vVtrcYXjgxcsdWq6NAvdIduWSB++zfAh4
kogEsctAwFp5FVpAUFb8nd8gG6lIPEawJXePyM69vfXSNpNuDqrE+WIPN61+t2dZmHytAx+uYFPs
Wr8UggkkQBQfDiHPVnHFMxhTo1heP1XPFPxguY6lLkIYATn8rwPZ3fBlhLRJRr4ZgH2H38QIWfCJ
K0u+M/Gnwr+LFGuRzLY+ur76Y3vzowOuK5a4LE76VMvHMp2FB14watz0LVd+cY41jJ4ygxdn9aS9
StdYf37UO3kumQoNc0xyLumtd5zNc7prm3VWRdltObaavsJAOvd1KZSbl+5Z0zXtFlv2CjToY5ks
5yZMkfiiJEADLYN2TrTb18Br3VjeJcgjjM6bB60NObJsjdp4RM9BtY9I1sWIIIAO0v28pu8UR8+7
A6U6hUdMmRHgJzW21yZrcK7GQHDuZgVtmMYOVeTXBB97XEf4Thaf5TbuPiWaiPAPTqCO+UzhwzRw
u91jKTFwvoBrnhgB0s04gqao0Dv6U+i7k+y2rplBLl3mCjccup9eKJjkFji7iOOjWOikIv8hnraV
ILjj8yc48E4Sa+O5MJ//P8RvWrX25dcXWQjNMv6VlkPOnoajXJaQx65QObI9hHGJ0qPQKZnqlay3
zze0EjochP4zLNv7wbY/W4gUVVX07XVFRiYlXutkENe/MFFc2peed80JaPIGfICT8A1Dp9ForDqp
IPlxSXjV9Orf5a60lhy9QUgVTsqQrPTBlGObCl4sAomKe9CUczUnoV+rl8Y0fNfcxOoH0BsVR1a3
yORVWP9mxlElzmDZStwWpwu1f0Ox6lnCbmiUHr/pv4qR6a7X2viZcyV8GGzDZfIpMhJpAxFOV3cY
hsFSN+gypWkwEOVqzFP4V5NDCfjMiFi4qTmTjv+d1wX3hKuM1RJufiRrxfCuIzDWTW5mKJhlJvye
kNTWz9c+g/ZD0EWGWvrOiu8YVyAfZ+yPio4PeEzjpw5X50ovWgTdZmILQdE9oPlxS1ukOvLkip/J
Y+r/vICvQEI/THNNu7fob2ZbddDPv1kictfDw+3XcH/wS0JpwhMjZaZGfW5hN50HF6x/qZs/825M
riGWvhUCYBX/3VoxJQ5cCVxPTiUWHRs3h9pJAXQ+S+5BFKIhIeorE9Sz2KsyrKE2/nNs9CJGGU2U
3mvbGhnRKc4CopqSYiqxIAGtlBjYw02h95Bw5+hNsHuy2fU0/cQnRbzri7Tss8ECcJVGbNz+3xHN
ArL/4nx1QEiABvUAqgPxosgtZ8rTER26V1RmUwBb2RhCVOgiWssR4YlnbGwRsM3ZVm5vzGVF5c6i
mzxQ+nysC1G6QMaWOztNcPO9HmkqDwoOpmLcgP2k3FvIqP746S/RE5ztWJAglAN2Cb3i/l8hvl06
qLQ3I3SCNw21qAnDRjfbE3HlztV63SgMN8hvfw41XhYMlwIz/KzQbR8x/GaGouKO2Mr/l2U9nj7p
jKlmIu9Mp7yTMUq7DIOc3nm729DFfAbbOrMa9Wk7jBWxyJZLI9WuQ1PAGGTGgVYiMNYvlWHKrzeB
4PKaTqayzUpIGJEJk/jgfI47QjXmnMoWqAqjyhscNTUP8unYEbPtoy07bugYY5WM0hULU7R6wyM/
fZXhiww9tGoEPEzp1z6C209KmSP+C/yVckKLpq6en4Wzy4+ncTOKFuAsPXBdjPh+Q7d6+rzDD+Ka
FjWRe76t+GauM4z+1FyzC378c3ZtWbOkry/o23qn73VNAa/hsh7IzdWvKuuvrtaPF17vnIEucrA0
hYHdCGvE6PwrdT49UvcNclb/aGe7ccxlDa0/gpLajM4rZhlNd+7w9JxFGcYpMrH2ewWhLo8a1h2t
AdINCRrtOCXq1tSGXPSkOs86GK9Nx1+8RIs+w0IFSdGNqTEB2y5/J6QqKdNYlp6Ts5FkwcLG/dN6
+XfwdfIglZ1qAMOY++0YvdnCTjVEj9e9coxpLZRibadqUkc4MsdEgSvCP+vvBntPjwIbB7SXB6lf
pRIvpbJpNH6d1mPIgxvkh0ExpSBpNTSbBHpoHU/EWtfpdSK/obX2SdjNM/l9ZBHjgSoZWxOsdh8Y
CLUkSG6dwQb3bxvSdiUXgDv3rK6XjQzpBgZrrz3oyKwjiRgZMBQtXUQ6cBFaFaWWg/A+H/dMO6Vz
d7Rrz10t4PaYbliq6wW/E2yob0PHOKWQpulGCJS9DDL2e11rLR2AOY9gsNHyXLI3JAuYFhG1qiWM
LAtXgnkrXQEXhfcmLzaD1b0dpjQcRu0pZ31ih3pv4O0ljuFVM012heN1R2W7+J/YaZZOqZSGCFE8
NachOx/ibqNfx0lXQ6J1HVPNatT9ZRg+bOKyALvYKw6C4loy6GECcRBzCIg83jzPv0zvBGIhhRH2
Z9PT3jAXXHNdCS6HT2IiZFE4k2S37lyuh7HbYGJKsRGgyMI1E6vgXiXPmvAQR9aCL2+dKdqghDx7
J8/5E0N4cXUReCAHXLvUEDF4Xe8TR+F4nHp9NX9ldhNeXcRKu6tXeWD/D2WHPexAt19rsJbWI+di
KfMWEAJ7pu7jPE6nv8QlZIiK+x3XaDNaWzU82ru1+HQr4S0ZK1WR4psi7U1ZS56zd+wJmOdD2zMc
rQbYbB5Y92zHHFLknWiGTFL2D75tKlxXUI5MSEhLK4rSkgm0sHIC2ke4jIFtK5abe161N1s+ukSw
4p3EEY0WcZc+ddhG62lIS9+9e9d4SS7Mth1CIZWfEsrQbjSlIa+2NUiiLO8SNrtp6cJd+vg4B+aX
rSpkVe3wjbhQ4lplUb961QuZimYV+1pIXUUmqwYxt+HTB2a6clEDG0R7gCRJwon96WwfngEP6hhp
5022YZUz5wR5kox7wGeDkT35Yt1EpP6INdnmtKkg5zBpGuAtxDtqh58FW5TfXIjA/SH92wEBl2VO
K7RKKuNgcSh0uAq/6c3xhzexNnpXbMAAAFGOrCWGyacaW4BkZPv9inM2644WOEAG9tfiL8cGEOxy
9XcMPJzrxNezoHFrj887hf6+oYCCamZURm+mCCGr86hfu4HM/3wpZUwoNFaKudZuCjkZoJvX3BF+
XKLSgP1lOEF2ioPFgm7ZO9Xghpvag37ymQZPnptqHb912YsLojXVPaQc9pbmlbTLa2x14CI0iGBK
/YBjrnhiCq2edTDez7aNvjIkqDVDEzhpL/nc40dQwbe41qljUdjJKpO4Vk4lfK/Yqcx877iSkj+q
Egtuuvz4/IWV5JDvZi5aFA+TTBoLbWITRkpNYtgzYi/J6/sgdmShWRt4ZHA03xKpTz5CYZRM0+JP
0DbY871surkyKv4HU8Su+FVPl1fNpijUc+JsA9DfaVb345/YpaJbg/7bs4cTtwwYlMRIK19SEpBE
7N2s7S2+n3bf1yyhh4OagbtyEKkhA8xzAn+lVqwxdGsMYEL39ONdvYuwmWYkw441knyqt8QaSXCM
DSHInvz0VvJHv5htjJMt7KLoIODcgLfvT1qPqLK+4K2qBxx+EfKBF4tRoYYo/5e6MX7VED92aTDV
KZxche+a3DEMwTdil72BokE6bXmiLzyXkSvEABuEx7YXqf/kMtdgmV4UML4t4mvFvlJmuKGSdLOU
lTesmrdk90X7ZDOMPeBD7vaNODh8FA9mf7qbVSUlgv33rcQfGXQSgQtkxBchJUGWe1JyUd8lt7Af
nmqneDhPz/ZoBTPHtmH68lPNDnL8WRliY1F1tA0vNN6hZSr/QySfFIL4Anynr9woCSspIW6zrIbn
pAt/y/MhYdzO47Z7SP0W5s1LHqOfC6UEWKnhIFfzZA7zrViwmdbZAIY0R6Xq0m+DAVE5Trm6MTNe
I5hhQGxKWsECggSb4fAHmVW511GMf4id5maPvd5fbq2Ojj/6BLoz+wA9YVCPrvKyjJ7c1r83+0zs
NNlTPpCJvM+YlRP7yN75XMmjnhjkm1KsZ8+LERGUHb5guzqWjPVTjXzGZ7FyR+uhHQMHAj7/622K
gT1c9uf9+P3tNVFiBe3aCLRoZWrSp8R2ndpKsUscDbxGMAL4deCvC/faxeY2H8NjYgCscIvUKoas
+9sxUzGvS7AwbWNbkoh1UlD4MmdktwVWjGVMHmZjNNi40hkk7X4+RxkyGaO3TZkGhP5sUVFtACMj
P8+B1Nh8YnPkXt5n5XX0zSmzi6p/J/QJ+kqo7Qq4Idk4HTqgwlanMMhqKF6KRboUMYZ4zzRAyLP7
MZpinQAkCUWomYgpy3nj2NVg+8UIx2oovluDRAMNDigRyH2wIg4gk15K11ruhChc4q/W9paQVj5Y
PRr6iY6YDixWh64QbvR/82oajpaE2SPaotqNQAnIYZDV7GoYDbKFL3Wl30Mr1EB+t5E2ZLX5LMEU
3Qb8ks3+fDKCuTcgOj8sDl8xrX59Caos+vwD6tiyxrp/Yp9ybEG+tUJhUBOOqZN8Zi4rH92Sniqb
P7LblXTVl5Rse4DAf6NFYrqyi0y/QxVdNA8k42gCKzDwT5fNVwW0HYn4dproBCn6CxiK5FtLXVm5
v7EmTcvVwDeDwSBVDY30ihMULxzfWnmA84JGrKuQ4+V9ozD8WUkZ/U+zmkw/03ZNsNYhiYCkq2kw
OTMKNIaBrpqmVGjib4xfqexVccM61vKZfxn1x9QxIsPBu4smk1aKlPYDpQhOIsQfau/i/F+btf0Z
6tNrsuOn+YNCyGWzoa4SOqE0LampLufCkIsl1cedkePOdBf/kRSgFIeXGOFg5y7vzDYhFrSTBha7
sll9pI/e7uun/i1H6G+kIjzX4eF/SH/JTf/ny2H9ZFQR7j6sg2HHelrViI8ge5uqUmY6PdomPcgm
ihVinIPauFkQ0FlA8dmpBGg3RLk3xCO/samVQvIuusoBNKvTAgKPd/sbeO+WErBTwUxosukMM4Wy
EgpMcADW2L+NpLd2R3wzkMgg2XPs0JFZ2MtDf7O5NYNxIzZtWuy0Zko+knlc8aOj2es3fc35GHV3
/ywzx92Ay6N3M2WFsdoOqWieHpyLGC2yXYSNRWtPAg5zrZq9lfvjL7+y+3rbLiF79Lk0WMJO/rpa
tOy0LFW6A5SvansSkHItwH30RZygIEkO0u/0ZrT1jSvz8VQTqpUSoczqQoBKMg9qPRvEzT3LRNgu
7id49rglFYIpDbszjXmetS7wplwWZNZMESwo/SuxkBG1LhWhNUzPPrp5J7u5GQK8ufL7pRa3fCXl
gTRhC4OzCKxn1wm8AcnBCwajoC//LCHAD46o3tVzY5oQWpvD9/Vs9gVrzXV9dBvN3PzZwdRCA52w
e0vfC6Gucj/LAGiqgL6taz7QhfuexnheXE2QZnpH3aYHm8UFu+ChT12/s+dwHvskIdKZjRAy8kXi
HjXD3IdgW+O+gW2DdDMEOcf25teZUeO6gk/BxsNGy9T+SE15xrTIYm3ISGp5RCGFUcQpPZiKX5tF
OKsXobFzRHyvNeJ4YkZ40VlyusHZYdAJxqJveQJ5hQ8PjroiyDoHI56fdocpgztXKePK+2yKUq3B
98KDgaMAKHrmAAygxVIUoNM1NCTbnbGWyhzntaSUihGh28WfOaL2vY88tAeyrmJffJdV9gkGe88h
iVVgU+Bqt380V8rmYzXLVG0dgA4mKziswrM7Km2V0cZqPKAq4fyRFDAnJGoVJQLS39Gz0s+82tu8
kn0wzMRiaebmz4ACJktX+yZtkwZIhPdSpScJL2s1s5lLqgDVZnT3JyFDCliz2k9caZTPLQ2tEcZ2
D/aqLfS6+uHWzFsZhtSn0PhD5ZPNqYRhcKMvLcpwezEXNp1NpNJCgBz60S1BVbcuPtrChRfXzyKM
LbAHH9kZdOzuZnNMPjQ6VMiIPlOcpiXTi4wbt1IH9T6YMr1LaxwAEO5GFpzl11HvMjLyun/RNul0
GUWeqQKp4NiKbeLwuUn/AdyZvlpiPUdHZ8aSH99T4TEoEhjF7fhQ2V35+xLtB1KfKuDUqm/Uwq7C
Yg0O57MQh98orEBazsp4bdOm/c/xoEZ7ffO/uYkMwUc7GG6lYb8FDMXGn+3KavcuoMv8wn/Ttrri
DtY2aX5gmWEtIu3qBHgqp5ppdePNudVOIs0Fvu7OFKbsKHvyge0056rT7cQ3etJ2e7/+B3EX5744
Bnt35kUzFT4ERQBuRTcmtrcUHRcUTxNpmQT7OFsdbvBWPJzYHzjS6cUuyhxgKXCEvr30KgEkkhZg
INN2Yda0YZXBdV/0DAvUci5dGMNXIOD52CpT6Al7lAMSec5JO9zgltSxGT0f83vC/iiesZRkG/LC
8gkc8TZIYTwV5meYRm0xdKwmn+ViMPV2Ue8I4qSaQPmsbp/Du8zizxWhRaRwdy9nk4/iBGVpX42m
gp+zKm0B1sCJCl6xhuzsdUIeSE+2OML6yM7e+2hdilgMqDL78ixSosUtF+6r123nib7Jr7Pkfl28
r5gtTqJmEWUe1nHOZBj1J9TlTOBPNc2qsE7GW4bTQFa8sbY4m2KcVPp++XawN6DA1wRCn0QayjwE
DlpsekC+b+JUK8j3DGljrbce4KyjH6wbfI7u7JRHIb6uzidN8LO/+eJgiaOKD88phOnE2+l2vRUt
Zg9U0kUrQdBW657naz1JqPtLlilGeYKBQUQp5bRasvJXxP1p8Oo9gjV7CNoIurBz66QC9ofLuR01
xxdI28jFXBoy9oTd6rkWx8s9B3sNNBsUQaMZYw9Liw7S/Omwd3Q7eX4A8894UmTExYnDLqR/u8Yl
tktf8cOvlgZrBr3GPTSRr+fZFkwxy816nvEvatlr3zz4sWm4MHLNhf9Tb4ydJAOSWVMBqllLIz11
SfN4xPXSneVenZHlA0AkNQfuMyxixaHq+yxVVnlmIXmMJZPyojvHi4xP23NEh6BsXLIelBb2QdOG
NYVqd8uiJzP6MgGIa1mWAOL9BVrjLY6oCZOxhm6FJg+u8zGfQ2amotiYVIg2iwgwTKNXovB7U2Dj
40rPMmLTf3xeasqhK0NxWdBg4Ob+yyCGwDV0iAN6afdj9612plZZliu6rS++H3XrfLR9z97xytPT
Ne7UXWWlMQeg3NEETYjbz1UzphGRbS+oUi2BbiOWG78+typM2BQ+FzyXQ7R8S6xLyNjdTaMprdV/
Rf3eS6x9BKg0a6R2v+Q15inL7li6/lGXczmcZSlKnIIbYMi0LI2H9IoPu/f/ZhieIS9JrrbsWVk6
IC1Q0vlIOBn6ON0No+5CeueIugl04FGJsTnHKqGBsWajxwG2JvYYEioYVStLF6jtazZqTa0e/3ES
t4cEvD4+okJEBKbHOAvbxUgYCrD8ShcyPRz5PHNoecDDfhY4elVG+/A0MpPjnL1BZClrgUq1ZYf9
3E/FwaXSl24am0oPRtn38USKmpTf2f7sFs7TWr2KSkUpa48apD20T+dyKxmQa1C47xc9FkK5bUS+
OIoht1LQI9cN34uhImb5+ichG6bQSX04Fkk8G7B4Hsoeu5wfynXzBKGltC5cfvE9iLX+0869pYJr
uCjNBuz0AAas8uZi0WgJtiA9eZY+b7IWsT/DstiCUs4Z/q+rbjY3d2HPKaQD+ALELpRR72DeAVjA
lqh7Ryel4MsJQwrrEpzae5ZKM4DQ/2InOYWd1U5NaytMlnFf0WSh1HiykAyIcbjEijmzAyLJIZ1+
hZLJMyDmVMvrZ/9bcRHSV4076TKsmZw0OCm/YTT0sKusBCQXkBp+Q8QIOJnRUodI+gv+L2L/TKC6
IEER+heqIc4ytW8J3oVdzSF0Ks6t7wkTZ/+/n2jT2FwAuu3wdfgKUChYEGBW1eOY8nBFwS4hn8q4
rQJeHxA68tP78qDNNCri90Ahw+SGS0Xjvi8P2RfJNcdtSxOlY4DXlZZfZh+77LcHsc8xcC5y2zlk
YlDNem3Vpd8ZDS7yhLFcoQxyrhJOes2uAfs9TM/qoG6xWOotABowyATExuXDjeC3x+/2FtoF3PDL
HZlbs/Tb9qP5wgjAwi6jAWt/rMKtkkonQAuuHYqXSxLgjYYnk8Rlzvkq44KyjnUMBOG7/+SoIShg
iAOQa4IyXchl65jhouvCAWVqFF8l2ygOAXtyeEV5QpUXUV0TqlFR9Y3zrrP9EPQJSPY/fW0zD+HR
oLUgzPye2rT1QJHV4ov7ov8dnijmo6LJ6vjXYjohPa5JEKCJWUj/DyL698zhFEtXKtpO4d3lxb8T
SkzwLzL1E1Pkqv9BlVWRwah154EovZhULCsWiOgryDRNbaLb5Jnh+aBQRBwWKhmFeKKiaStfWdmU
cQZU3mHICYlcJeL0qp8V9/JA27fgezYKu8AOyUC9aT1j9lo/ahcMzgMp2uovuV4YMLyPqmDSFxt+
eok2pMmFEILZX0NRZ2b/rQH2sZ/nHSt0qg3SxlbvJXeEGoyBShxxfqJBaeQOB9CmdWtDKJUwCEUn
CcGTxFljJ6FMIbRrB7xMMYnXa7Pbr9+YQynFOwRgT5QZsM3y4zsbykQ+N7BqauDllNe9PDBV93lF
cuC+c/YqbtI9MzyK8FieLu520CTcB3rL+C8tKet4D0wfaFud4x/qED93qQGtn1wkYYjAWTU/lQ03
cdub5RLqNuBLsss2nfb5bA0zPRZD7N+CavhAP92f6hQhUXxM7OuyyMreUIyf8dnA7pKCI3x9GWUE
TmgIXTFYqqP9UpWM0/Qc/R2c2tQk9oIV5LaqzkZwMRQn3/yEtk2hFOl8f6KHJZ/0j+m6dCs/PFAG
2qp011KPg808iqSz9ghOaI+JFMYPuhF8JK+A9DkUhu+2PSeZZ6CqG/nRMLsfqum8mPPKSowoqFuy
jcOASWFiE9ooTT0uRtQx9szhosIa1Qi9kDlJoRTfkEn30GD0r5FSpvtLEZHudA+WtNmW/dkHbgZ8
Nc6LQus8YfouCuDI/pgqoq9l29If3BCK6TpWqygc0I+Xf2KZFzLCX5uDof4tKGIYqA8aCjar4cxg
32Iq26wAnAO+j1IoKBRhz47/KQ6mgiqqfRh8qdYQ0l/jJ0KRTbRoFZd+drz9Nze1S1KdLEincCgh
/G3KnMzzqlUFzt3dkQ6enwIhdmIVZQj+szpdZTbDOyO2VGrrrs6TUZj7x+jELmf0dfwebsYMcDlB
7rtgOBiizxQfvCYPjJ3Eocni76XPFbpT5KvsyPVkTNN6XapeyLmUAT9/oRQ1xbSDiJkRZBDPn2bb
KWLWvpFx7kLb2xa0Dp9c8+pexGWeR0obZZVh4iqYgytb/5neiQisx55LvZB2ZUHkMJ/cPcYC0w20
hN9kdaLadY1FZUlPDgZFtlLzX1FoArQChiK6utGrTZvuRJfoVxhJZzw3p5QXbTfEnIkpMDsgDVyT
t/+EucxxFPQ1W4lLcQvP9biHz48+yCejmLglyU93rEdtUefMnieoNxc+pqhVOzUPAKf4A5qtz1Df
CCflqI/nPE50IU+/tWm7KyfKffoPGdAnM27V6fGED5WqlNloIjizMWnvo42ubL0mKFA46a9Mb6hl
KS391Tz2I7mAHomMewMr/NvU+JlKk8Ypz2m4gK8IneI2Efs3fqPRqTZrxuo1omuej9awOLk8Dsh/
ocJYYiUW4Jcu8t4y2JaAN9IYARzrkV75TnA7jUUqhmVDFnnhG8bWIhduJhEDCRXL/PmNf5Xd+jCQ
SsDmWjnqtO9cCZEQb5J736NkWtdEH8PvPFlUd4uJprrs688kkK1Xn/pcajoLEgvr5HtktiTRcLus
pAT0w6TRcdTlgL97hBNG5OgG/s3lHW5Q0+JNf+RzdLzA6Z4lKQdaGRJLHSX8pYR/C14XcM8k5bqh
W/9LiPAOoJwc43w+ANLVs4Oi6qC/vOE/EYVNLVAjH8RwRVGzyXH612haMu8ZvL8eVRfeYWpHMX48
zSOk9BsB0NJIuuAmZV8F3DUKp8HOLk75NX0fvEkeTDWfH1tjiZ/SSYY64Uz0h824yujo5kY0hIlq
UPfrufL7nwyzDXamkNW0W4MG4zP+TiUfCzQR+ySgKKAEI/hpwojVwhQB1XFb4YtqVWwh8GfwFuCe
jCgacfKOEURob7sx8J6VDD5enR+FJt0ZkiPQukjjUwAT/nY61+//eYVtNts9HSrSrtMwtQ4BRs+r
SPKTNFpefYJpnfTQd62yzt5B6eHrqUbU1JoGnnBjREuELsz8xCUk9mg4ikpzhNs/7Lo7pbFC/z9l
eXcIOBlW1Y1+TB1Bl4N3fEKgHCHvRiUfwFVDNjQwiu8qLadpZAxWbSxkmdxsV8nPAwjRwyZwX8ed
1hWXKhf8IZWDE6pRpdiNIZBSQpBlEIjF0+h25XkV8ay4VfhYg1T1niYF0Hk8yB2Jj1Tlmjkl6qQs
a4pUc3gglOAhhlhepwbIZjc9lQQGJhUU5qkU9nGoY+dPfLG4ZKbPwrrYbgGSTRWAIJqBbd9g41rX
2wp1CPi8Fvbl2yvZj34+NbxMlx9wBK5fsqd4qyrJJDoglx8vV0agfmer6Ug8mL8q/flQ56ycJVVs
7sdEAWbMHHBQIapu6N1DbcKdC46pnYX8auV7LKXpNDps0MH1ZG+ULCeLCctvE4PRrp2Q7pl942/N
jPnwRqcKac5X1TrF+DwiFd6zB7zxQGv0qLsQpa8xyJBoI7XDOSLg2vRmmLLSqe5wZk36Y5zy6bnE
IhaQRInBuJivJzljR9LLagqAWTDWOWoCg4SwU3ZOCYlip9TFqYZaRi1ScDS495SjqADzG1fK8gGm
zvH+/bo3I9Eg2HhmMmxmD9OdqHfw1QLU7TVY3oDbA4IF4bGqMPc6jPPTS4HYnbFQfXx+HWX+pDbw
oegdl16z2PQk6skQIOJSohsDdLuwK/3oZJlCnNSmRaH02T/54DfbYIhLkz9LepB6KdWSi7pLM8TQ
19AqmRNkafDNPaVe/OCUlgP39kXbbCMBtFhSBbGtwTJ7BSNLDhpYPRyGSBVGfvOcwuMa61rLyXIV
LSDjKvUg//HeFwjIiDRacuuirfBLGy+/7cIJ2zPgClx2+ucUipnxLLCeDiP0T/eHdqErqF0BMnhh
qcKMIGgZcf4QF36MAU8frVV7aNjQBhknoQ52r/lRAy1RnukbOagY4x55wqrF75SToA9a/Qk52yOO
e7KGwj7l0tD+SYl5ejAABYGLSpFuLLiFfCM+KaYTDXPhfwScpQVA5zde2lzHislaVbeGTH2hgm0+
wYvBE3KeenOFrEfX/NLGW43KjQPM8H5N1I7Rwc/t79M0heDPlCz5PfimUgwBAerLupGCKoZplcw/
NlecACTSjqDgwDboHVophsLqH5p1dm0tLPWtB4o93QfaE/21T5uBQRbuEGIRWgkb1IUh2I2hrKco
+sRk9QUGKv8aVmwKr8+jScR2bFWaxZdpcSojw5INTRSBx7KSBw2ilZFFjsHwWnIaClvlSKJUwoaU
F3HmZDSDA1bNmICw6QnWUTqDeW8NQGLUm1F/txQSXShDxlGIR1/ZtM/F5kw/J+/y9r8eIXvcwKsf
NyyFRaqIOrjB+PsO0bfkWdO4Rd7aHEgpUb1n4lsPc+oMgk+1N+ETX1zfcZS3CKSuqIOn90IWd3Qh
pg21AXoKngbM0NzdbrV9IhC5BvtL7bMbr75ZXmX1Y1pO6Bm4WTRB16aX6+SUPI1XIthCjjKSYtrv
qAo1Sx1sbpkBzro9E/s1okDdvE9okZOV5Msj8FTkDq/fiYz0d94V4q3IX5XiHVg6l/6+SsSbVSsQ
QG2+BHNSJyKtq3m6PWwD1k9KKDSXVmaweeQ9n3K+pLHNBS4JL1qcZqLRFL+qlG1bxVGrUUjhDwpe
PavAIPYWj3AGxWmtYLDYmiFzRdnjy+DF905dcu+nuJABoDpOEnRamVDVuXUac5wH2dfniBTLW6m2
m2480G22qH9vi4+yWii4H++Q09QxwymW7/uj+e2EkZh9HH4ZvcNmP6qxcvob06z0HXMs0Vmx9P7l
pH3o3VRboWffKrO3HzD8vfoAsILpKSUN7y5eFl9iW0dUum6TFrIlGmPeCBcZD4ZnVp2IlAk4YqRg
T8WXe2BL7f2tKG7+Gcwlyv8v6wWByX/jHSlMvTm8O7fQIZC3gz0dtTsZODKbnkP3p9mFUC//4BPX
8iZG1t24e74INNmiEdZAF/jHawvun8z7MPOCPBmGsMw4cXRuiW7RvRX/A/XPHsrbzj8D6+sOMDY6
DqK7RnggZqsMyMWIJGnJD2LCrse4BYWDmy+DQpdQBVShXbzYhbB0tWzQ4OWEdSK8nvyLvQE54qW9
B4uu4Q5+NmcggNdOmzmJZV/orKSTStQ0/+nkMLAOOUb6zMJcifedL+nbCATJj9C8Pp3jwHVIlN5B
75sTpWXobHfF2KNb7DB3Yvrmj5AcPtCkYxX67vR/znYI192mphDNvSvIA2jYba8npN57aoM/5G0a
YOMn7ZoGDlwmmQ3PUVklO50HTg/OZrXowDt4Bna+2KoUpLHPuQSweXlBDY+qS1k8z15bgI9y/PTt
6s48A3VazcxrTl4QBd5ZfDUa/YPovBK99pc+vKWZi6jEeup37y8gNaV/xlT/zRZC6QYhB2CTpwc8
a4ConhKkR2ESvMEfqCtxoaErbZ3uALXJBUAYDa2RFVg++cM3tLKhX/MzrI0uPwGo7V/An8v7Ws/P
ShObtbOkKHo35qLrNLHR+Kp36I1/TSWD83l9jEQBbhh1KIiiFRc1qT177t3C0KhpkAXEjW7MTdw7
3deZmdWMmYP0sx1YRHxc3IU3JeqtDTvCGSDgLpIX3riZfrHizJFNfbCY0nSRILykN7QB+pz5CNyE
dOOD4HYOUtOqj19NYHrZzVtob/Dqi82T/w/nQMJSCS/KQyPeZF4uH7rN5rh6WdqkxaO7OC5H0W3G
ZuReIWcTN5YJ9NefBbeYcJ5stjzpUvvOXm52sTQrI2x/5LLJNxNF0w7NnDYCVO7CJTAHKGxsx7j3
chDijBeTU04izROmno0nuvXHB1al9sc0V+pbZVIAwDN2LlyKK9rrbpRCYWvAhK5fVIvpIoFa9eBk
p6t0wXc/AirSZ35TorCsCHbmuqsOo57pajbdriRKkXAamd4AeX9mIY8zIAZHd3jeZA/KgZsmJGjL
1WDlPjcjoqbYdiwCRtaKccLUjq6Molblb8vzmumLOjImnmZODainMSPrdYp0oOUlZVkfXIWrrPIw
+01AgUpoN6zD1caGOkN3lcaQADdCver1JT8qlY2AIj9KJ120eqRsG3fWYVZ50pfEM4UctAtIUz3U
aoT8kDiAm94R/b3jUFYER8DAMn3wmYPfmv8EjfnYeKSq+0A5iVwZTIZu6/ukfqW0oy3xTlgGp/QW
70yzB/s46n9P5LKyHOeJgsgpb4eQHyccZ4/Yxnjwg1j/I/s7iPOSNwMuh4HREnZcJCa2QFF0WXID
diq8AJWv4sUFzi0LH92GbPEAJEqymjSW0XSuwXbzFKnmOPVYLY1gk92Xce0H4HY+iMwctRMIwKHP
EwoF9UKGFcDhEdi4DEdrhwwNRBSzU/E8J1gZhuC52CyT2xq0QprYer+/UP+dAv3kbomz20xrDA4O
YNbblTsgBg/eaQgumrWFObw4h7Czlg9Zor+VDM4MDnM4NlaBRoUG32/1/M1oQtydBhlEWLqVE/2G
zaQ/6twXQJ+ovPB/LJMDtT+qRODvYJ791u+1znkc2/dxFRjIMAmRlfuY2wR8dln2m8k7kjTtBSTC
up7fjVTZfcSpEwv1ahTi4xBm2KsAPSwMRtFfvdN/y2AJPM5EoZdpMl78CCghYw3l3iTO5bIeb8ia
zCUGzbqn7ib6HQNSZmUm3rRQXAmjDsp/gnlqvVk3n6+kBkswetdHE4Pxelf4PiRFQCGOE6tN4x7+
UcLQ57UAr5H7jk+WBmNrU4rX2Qdrq+6Z058+QRPrcHuS374KQsPwsD0StYB03ZlFdQDd9t+Lp9KO
x/RW4A1CUvZ8o6JnBARsWr931Mv1rfwlGgYcPvMCF77b9YoTG/E9Yv7JqLZf4Q3QfOwzdqoR7GNZ
YMdxFpc1bIQHCUW7sO+d4VWKMeuMDYcbslZyIXj5xKzK3De247r09UdUgNXVtxsnRXDm3Fsp0H2s
24GV5NL/3y5p85sFqIwwKd/I+3nlUghNp5ZGAoClblXSRb7Ah6KAsMuKoOHw+xvCWwhdcLOBKQm4
TWe89Fa4rrYY7nsnNOWoiCRO4+9MYMqLIX6/xwZwX3GkvsujR0HilHJVJDEwaTVFGkdXw3tXQ+JM
0OOudG5extAnCsrix93Mtqr2dKGR4p8jLExIw2tgcIwQwZfFGTWk00RtlGvBYZDpSysLniYSC/NX
Qt+QT40ZLsaDg5rtSjcan2Oa/FJMF5LFB/HK79e3cs4Nd50DueMkZtf4nXLD+KJfa3QR7gZ6Sy/v
Pavpw2N7qZQcCHNs8U2DUKEOxK+krrP9RDvZNOfTeIVJGE+/tflC+dzFaaFehP+/THIQBjUGyfJL
eRnkzHLM3UGWLm+jexdQ5efRvdce54QzofjKGSeG6hmld/IZDUSWvsr5mongtMtJkana+33P9sAK
bit6gVwRMkfhfgMc1nbyJDEj/VDv7Fdw16qNzgYz7G1S/E+Hy3AofcO+HcMp9UZAXbXYKV+f/+TZ
82ncLsM65ouMOcAKvNKOVBwaBUiYExxX8acU7/rKuYAWqt7ji/Jm825kumfrAFfv87KFGHoLv6pL
M7li7t7iVcOmnVdXc8CYquMlZqZg74CIf2Dtb8RqS9cQgW058aH9S/ATPnH0FwyvcEFioilODg/w
y+OlEVjrB0CHEGOiuuZkXFLrkLS+Ozb9+MXBjPvKRiWFfChwcLYHpVbnnZKe+1SdLfKbVyH1/dAg
BhEcTeicVsGhby7tX9U/FxjSC/efu6c8ETQv/DdzB4Rq2WfzZIRsYCsN9YtIk/slPqDe7Wrp1zbj
MYu//zDG8Lp920qBeTuXA+VZvgEXeGGqWfzgE/AtYauubCB+06EObTBLkbKyD+toK6Bd3MBB01jh
onvKLDd0hMrVJsMvuE1ogG0utRf6Qann0nOsidM0d1svShfaY9+9UKHExeakLVJ+SaJykBl7+LF/
T0h+ZEd6h7oW6ns28c8tzW/Pp0riRXjFdpUGV7CzLEBTjXbS0aMpi7JKltg9WX423VC5zrrlzPwn
emowsP0H3nNRwj2NH+fJk8J+93NjArTxaZTa4YJaa5g6AgKn8NWz0T6mTwW3CkDL+kfubOFpUzV2
DMJiB8lR63rFLYrfN0Vo62RBZtgzvXJoSNCXLsdCROQqOWv+eClnMwmAQpmhOzPNZV8D/DIv0ua+
ZQt+kZv12fLyDYNurfBBgoey8t1CocTnm/LSVbytf3a3l/iOmUFQ8mQCCZ5a1lvkjgjwpnJN9lx0
3W1QxZVjJPbgfQTMF1SBNRqvYHtVtDERhva2tA3lXz9m5ZCuvRKNN54v8Tg+Mb5dEMVv7BAg7yD6
SKo/ESWcgIzJpCTPSq7yN91Up5FVXXdzquy01RbYO2tuUv88n5/r3y0FNSKmmj3mlA+03N7+gxbs
VNoJbEZoMl9rCEDPtLZTvDcfNfFoue9878jJy0gUu7ZuEjlEik0/M6YdQwaF9/We3bF27FoDlr+J
zDs2DLMElpVZJkNpbErtFe51JGRiOHsc3FhZB3PR8DwpXLWBRzAxPd/cs/GswVMhEgDkCliSOkoQ
VmoPLdfItXzzWxuj313kbyNTjYewUmWMsWDpCL/KGCTEKOCDgedHy+0YpaIvWUCsANRGDcDHgsCW
c6ThKKTrzMMTwIZmwnwfa9K+bfErT5UzF9rWE4+iGSUILxQrKTeE0Isur+Z88byLuNeYEgdgehUj
pNkZVMiwl7W/bEWCFkDBTtarEI9PG1dx60+Cz66VRPvBoacoYPMCav0UPa0kNhmgbNTZLEcmLhXY
SwLHkRvdiKiTibMAwObAkfLpreRCJKRYQliYvDpDmKkhObnO6avV+IVPBCHz5bAYMcxrt/WsybiT
xLQuDsazy+q8UoYtyWD47Eip/2THBq4KU4IBzMJNVvAWgui0pX0YpRBA/vvcVwwy81//6yHEeSVt
KpBdg5uYWyh7NUA9nYPWnguYHsaj6uq+AU9a+YiBOmrBgD2csRYAO8w/4iy3vby43A9FSLrA5s7p
Ka3XKV06V032QFzzYivUswfHtpKAcIr/aGxb3R6vprUheYc66Vd/Am/fQkx2PnJIKY0ZcMJlSJsc
8Fwi0ai1uXZDMrchV9CFw1r6qaD03Kc/hIVfkPlVDVZXni6Yko6j+4KjQ6IELwU5xpcgQQtI/Mne
/bJzdKiEE/dj3SCMgCwvWnt8nKyVVtH2SLcy/E8Q7iwQFuNqvEWWkXEMD5HftKceH0V9LEg4qFKk
SZIMdtFfWC7VvWg5bfCSOXQ1P1qDCkI5w6hcnm4HUo1ua32w9a5ZL7MVO6GoX32TM/bqs4atskUf
/kpTXk/6tG52xVv+gZ8JAsYlkUxefBCdrXixwlb6mXYUflhuT1uGQCxnQZIuWaI0BdpUVL1Y2U7A
S4S81dfvIPEJihy5Jvs4qwMPAGeK6b7JlR+RFiRsq6B6KMxpqWq/lo92Y33yXgDr/mMWZ10tOhcf
ThrSlD4pQvDHznD/pFxNi5MTi1yKxHL2OztvD2oxz17wvRvZqMeaBLxqhIwRff7dPOIGtyDTVKAj
9cF4/XhA5q91i94nn8D+ggekSc2NHEQx/rwrO3j3C8aU/WxkbMkVYDwQh3AYS8e8YGUPHuLrYcTy
kGIl5v3LYK3KOw0eaO+K+eEdnhcwaUboU3qvdfEBSPAecB98ZI2eBTHff/bpi+IOOYOYkbgcT5i2
PiLXU+weWY6/Ew2+G/2BClgLBfVlArreA4c67GmAsNjp3AP5CbfaZuZVQ8jwPMn3cKWIkwi8uZDW
GCJ8Iz9EO9wtUZvc2EWdHdfcReE2HLvD19FCsLzhmxtjMczrvjX+zorjVcFEszU0EYMNPT2I73J+
UPp6UaAkw85s6+pz4AEluSRIEkKTD0pWFkFs3M7kU6dK+a3kmZsgZQPUT7wqBg9HCMxLKpy7m66u
W6S3rMUeWEM2IzeevTo5ZdCdGH95kFIBL7BR90+noLL8MVeWllNacfI7NzRJV6mQk5wLyR6vD8rN
Q16Vwm5h9ONV47n66eb7o4NJsXNZBpFSF73hRxtRKzpRMKPTGQCDtn3WxM0LBJLZNPyQ/P2kcMiA
vBhwJ0QeWghw/nIsQKxmeNyysi8bu4SUYsLEA8y4seD2eJHNxwiIvQvu4KMiNpNn2ylDgjwqgdHf
hvOlN1qG9prLlspzdcFKrdkXtYQ4qDQuj5lZL7geDMqMNasR6rGXRIF7dnMZOxOuAhuVatpOOj3m
EdTppBBUpeDSQHMRnUSqGlXd5z0EqllrpXc85JtQnqQdxSMrOhxth9M+xkWt7wRq2UQodP/idfmG
gsSfzttA6aEK2gizIiod0gbZBoZjUfR1IRTYKCUC1Cvsyv5dYZqQ4RY7B/qAKG8Nj8zC/OsI65jy
nhM+9sjNOnl8q/PU6o00ITkYPaC2Pp0qkwn3DAim0aNYr4071UsD0lzodzyhGldVmH0D4XcO8uOX
NVk6E8YZbTUmmGk+/oTzym3Yhn7KZB4helGKdHpL/enKFnAJm7tIj7xjJLS6SQr5UsCAF8fr5jEj
XlDSj+J/IHhwRaca/Wk+kGmjaHqE6lzmjkC6G5IGSii2upwDoG5lt/YdEcKlNW0L3GK5asPIIvHP
1sb4DXW/qx4c1HSQdMNEDXFPgOxRIIicWmcchoUZKAo9VnBwaidsSNBX5v8U7n1YpS7fcOORj8l4
V3idytLQdxRKLjcd3j2OXE9SOgQTqwBuQDCzrfqvePLNecbW/nye6Mt7CJBGtPBBcAzkL3QgCuYX
1J8yD0idpIzNutArQVokK+9cTl9/F4z1zoarnRkXx1anuqH1+r2zwrr12M7rrio2sX2CDOxq2nDD
oSyoPi+cYyGJ0b/8c/5x/4BtDv6hbBvXCKVrjWVhWepkN4vvrCnbmVMCb0OajlQmcB3x1sjn4A0T
VC+9B0sPh6xxcAzdEy3pzY7MTiHOtawSD3n800GUzkxQTTiAQV/UTa2v/dhaVuwmHiaAp1fIe3DR
Bugi36i8g76MPcGyhiu5iyQvF1Y4i14IuojfafIaVaxEItUNsX9FMrdnTUvqsmrHnTGMAAwuGaf6
76WC8r3SWycczvMBJzNt4UiLiOzpNRgq+mTfyzlOV9EiNa5tosuLYddN4aO3o6/Qmr4crTVxbfb1
2jwfh2Tr5F2cK+I8+9M+XIN5cIgmfHQbzwWIkJ7vP/xiscypbYkg9U+AldhTsxckxmI1l0gcs9az
11/TSvPLnVdMEEKA/A+2o2hF59i+JV99VmzEdS4zvR1/AwAaxWIHIhUO75WhVNBLeY7myI3z85T6
BmDDMUhqvTm3/jsXuv/QTVuKeB47vxKWkH5edNKQibe3ox2WonjEZNROZUQnYcz9BKgfbJPjVu6B
fUA++IeqmDrDqDg02bx4+sEtJRs8GXETWc23/wQDtFKgGGXerRYw70JPhdesBJq+Ura9Y9cigCGg
TfHLOMj1eHOWtAqp8Orlv6Zr9x87zQ519PzLiy28SnkZcnuc2ZPQgICwZ5BGzfmCj9TkqPuEsi9f
BXptmEGBNbUWANCCzeMJajRhkShlgCEeRwEtzcyDzbencSOsf2KCWK2mWLRPPiZzX+iOas9AWtss
m7iDTwUmc/SyFdHyg8LgrH/dU0kaRyeiS0iI5LgJ8W92+DEyCU83F2tkIuwh8nctaP5Il0+spSgA
BwxD4JJqR/+oUxKv2YR4VkLeF10nKCwl+5LqazDV9cOx9GD1G+xbT1reu8rcNnIIVKxHLIgRKq+J
qVb2qXu7BbI0thQrZYDzH904AZLMFDESVy5LSdT4moTetLsnZqSyvgtlDtK9OayeaM+z2TslzLKo
OQUp4sxjO6CPu8/5NXD3srHS4b0njz/ptmbZ4mxkD60N4/JZKjI9ZFw77uLGEDAAHUuklOMvGJwi
aasvsca2erZOOVuWm7x+GqY4kMnpwwtwiFCbNbqiMZ8kKgmB3q+zzcCoBqOHvorxMC2ckGmmlyVq
6F1xTQcKiSsPsM0f98Q4QBIH9pcnk4+dAoUf0BFRNuRw2MCvDR0NQSwbgOqjxmHgnopKBp90xCtc
PlXudMIeX0Km/Rg/empbDZxyhPZqkMJek6S9D51Ghbe4j0OKiaoPueIRZ00fOQCwoZYmG0klmlyy
UU44aTouJb25XjU7iQ70t2+sux0DNQdz5m80uy0oBzp7m3ZgH4xBRyJp7/VVKzpQTLSSlVz7QorG
27IYdm9DFgJQYnRjJCA0cysGnnP1Lc/G8nrkIj5dj0VyuIHMjx81903G9GFRzGv+yPSq/XXW3WSj
3eB4anuvBV3XHo7INP/wWG0b2Ont3rXev6GYfEmRq8T+ma4mjioNfjbvVKsdppbevHuS5cb5EfLz
rkenZp3V2HSevq6k2NgHXsiCcQf1qGadQ94Yy5Tf9nH65O7S35NfomE4/z7y0+4wh8RUaDUmmMig
NDk3XWP3lMRLBBwj+JIN0oXQ52lrnYjnuUbTnoyo9v/JEZU7cSMuwGQ76sM8hUOkbvA7tuAeOKHj
zPq9wIB5RLKlbdN47BtprER4O/UWdNykmO0DUGMGO0A9biPa60MWzk9MIKuk4t0AX70GYamwENtt
irDKjhg0WfdxYcRwuXzgq/F7zn+3+xuZ9Kr76/ShHcYzQYOeRgYQbAG/O5hhQClFaQfs+rkzAE24
WjPN6F6hg1UHdQQUyc1kmvj7cFXFYK5Oq2cZmGOzWiyYRqaukpKeNvSK8P4Shw18cd8dTodfE4Lg
YX0C0h8XLsWqK887KDZ3rXNSp8Eyiz3zB7O80KKDtJkcKr7c7t/+afGUKppmXx1IEkpwMPGL6Wwg
iDNUYYY7Nw6eTttW8oRnLwCDxaL3Oe+qO87bFt3hU2tbh2AacuaGROitUXAz6vrQ9sin96fvrD1f
1lMo+EAQxPapt0GAiLm+jWY4Jp8C/5bWZsL7sS2EneQFXEBrPdO7KwCDVOnKf5qomUr38CgPzACb
vOdITG8kTPRzYb3r+BNEjBYoonB1pwzxhInB59f9eK+VooGnS6ZFyF58o/vgCA89mh98qembEGAe
OuFVgDV/HbtvFwgWDLuuv5ND4Cld29sB3tRe1HFSEaI+No1Y8kNNfE9IrsIOSFzoRvO2jpvB2mYL
3YX29wSmC7PcDSH+CGWA9Q2RS4AQ6zdmF0omwUL58JUXca6IY/T4rp9ZHp4HOjGzT8qNNH4Wnc5V
8bJAk0AaniYLwlEGLqW67eEc8GooQhI43NAh9mTSfnfvh8iaLsuw4QIwKjEw+x06CSdomBMJ9Z4c
c7tXlb+F/DSaQAVHO/6hOMD2iSAt0p0QUgq8r2JHmWYT2TASZpuSkIV48axJT2Dh8GpfyxbIQw8U
VlZQwnXRZSnboPLAFDZZIP7iQPfKj3Sf91BhhRd1oCWae9ddb8dbBHmydaD+s3zdqJIOKW8kX04p
8t4t5jn4SVnLhRhqyG3iQe8EabnfYaOhIyrm9qlU+dsU0IM47jq5Wn//x1LoWNV+jIm8gqHDOaXv
RBidATAxGk95ycGMxsIFHqgl2ThkV6e9o6uMimB9iAeA4aizS0KSFn4oo0yzY5A7ffG8bhn7RKBg
eeOrhyOSw6TCrPVhRtTSDvXrV8G6mNI8FmJA5h/ASo4p2a0Y8N1fjewdggwIPPTfkGyP1MaLMjTi
D3NBihAj2Um+xdY83BfPxWyNwUxZrF8aQ/mq228nKbU0d1xLDP9WWLJ8oRiBoszj1goslwsbESNd
Nq0B7B/aXvUt8qQaYVXOKkM3MSkpyCiWu3FIhfxvR4Th6Q85KVR5w2Pg/J9lzmlPuoIm3BaKzQbv
ujTz7ALvyeQukx7XrDnZdozj6TjTBhZ8AVQZMBlqFWzLgHky7QQP+qu1K08gBo9KDUPgaYJlW3lp
XOJMEEyz7fV1WDeRNmEk010CKc35/O3UFtL8ZmMzQG9iWj2vJyOp0dDD2k6ouu7H+bryHbUHQz2w
rn3psFbkPQpJC+aYQ7s4InO+xEtjtEKd+3KQTqojs7e1zna6G+a2kfAsjDSVEDsl77OrcPr+ZLmI
ztIk1R2ZVeeMNoa8qGC3Mtt+AhmKot7/AI9LKt9Zv7FRoHOEfJo7j3rtHFX3CDs79blJ75lNBnKi
hL+uBAtWWt75oPSUTvz1hR/RjQm2c9r5gsyGlIpi3MlyvKJrX3yxFYMsWCCh/BBbc7YZwUEMB4AJ
tULlJGLE7IqK77h6W09cM+WwVrGzRlW1VUIAM3H4KNklmTyW6FuMU/zLYni7lbwAjEwV0F/1bH27
oWfx1WADRzWS+JF6K8sabSp/q9LCTaLwmlxr7rDWQoEjwQKGwoYJE8mqQH75hchVA31bKbeMmXGf
qXcSlIfOCwY0LFlMAXOLn8W0qkVxfIfq/Ra09Ho6pLt4SN2uSQWl/JZie3xPQuiddcOsV1V0eyvj
LjXqC8uSWGk1WfqPeJPeOnr/SmUlFkQV7MKBj0/Y3a5R0PgeDIs6gG7A6K09RqMKRm5QewHMTuTC
RSc3hL9r+5K+mgGTSyCf8LWHXpRbtpxFpdak0z+BhOB0UvMVWabpP0vnF/yj8X2N4eD2fGUXXMni
9zPENyAVq3GWu2Xjd57IsJVCE0F48+T+G00maInDJQJNHW/IHHh9uVROrX5kYvtcNKYNoOhq2nCL
1O3vCmZZ72qEneX/eGzoitaQ37e8V2n0oxBRc/rZUfNMoaQqiRL6gL7YiJczt22W+3mvNjr27FKm
JBzJSlvnFgtDIHQVf104FqN5Q/7MoEsb2fe/sQfhCA53hq7LhzYPLnVmi9IC0423htADLIJmPf19
4lIYGtWoOsHG/sW+SHMCgekwOxkZA3gueeq0iV2eV8DBwpNas09KegwD/yCJVaFZwv4IdXurjQTe
TLlfMi3o5hBDRzIv1RZbwQ7unjcAOqQS0K+JwOi+yd+k+NT22cv8T+5rnpPDse0NhgMxvU8NHxGy
7Q5GOkYr29r3MKopHh3/xooSwYyQ1+dRfsmcNrYzM3UKnGWO2zbmFd8N8/wNqcBb3ez6TYbbRjId
WOfhryuGg0xwbpULkkwwbqnhaZpeusoF1NQWMm10mMOxvZ7Juv45SMGILKdXXTI2TPiKb+LWXvNQ
JKQWAZH9+kKT68yVrGXL77b3UPalAk6chhv/eLd46BChZgVbKm2+kPk+4/qkTQgfLuKENUYQYdue
BLfuGrPa4sDPRdg7yqoc8festaZl89JFaubFyKnybOvOU6YVVG3RXqC/iM+rX9jZH01QSdyrFgGU
bdMQdMFOzS6RcAlpbJrTvcEzpJmQdfbidbU1Ny/xjbTKYCf+xLuDF957keATLzWkk81kBGnsTqMl
IuYY2pC8lQYiFN2EwC7FmuhMYgqfgz7czkQzRcnRroakkjBKyEfiTm9A+aOhCwsliUaxAkwRFRhq
c60jZ046W4d15hd8Yukq3RsSVJB/I/Rq/7WxqnAO7vTvQacEC3aVUwdtOZjsL7rZJ6SMaGDlfPgZ
2abdhzHw1Abw0qJlu67MztFwcnWvbbuSSF0XctJ+Jw8zK/lk+o4AMI3Y+/OY3Y6vvVaL+DGGLWRp
pz0cOkROpqpBJdNJEWPjv9+1HwdgeVmS/IYo4PUc4aMFvggmoOley2Xz9O2jyhtV64sHsysINvg5
MAJ9ux+zX7YcvAAsHhuYFeOqN5rXWCr9eC7R+UKi+jV8tAXilp8K46UsCZUhjDyXMz7Z+GvOkYU5
yAKsyQDd5SK/5M7bktwpacqV6N6AvjqWYvA6Ufi1GOLoBlZpoHkWdcGqy4YPPmx3QNQeQ2hAmnR3
MUOGVATn7X8JdjI+WBOJQcDuTJ89enGPVYJk9Ggz18RoIdmIori4CKKSw+VooJYeL4L7wIAN4ydI
nFsYF+HcqjTEMQ8OftQ+1z5Reo2unsZ4nFIitClzUFVLr7qH9dzY2B1dqpWVoMQGW8RI3NcPFJPc
5vfXVi7JCuqVI3B70pQLfJL7fTCiVBBqKN79RYl3San5DFFuayTob0EonxT0V6oWB4DLszfohgiW
zg8xOr2lz5oQi48Av1UlFCtLFp0POnFmfR2bwTDcbCASmXBdPuIQU1EKC0LPUrQIHCbno+ol9FH6
fQ+6jdmZrsu/0QgRabvP9/DBeF8Na6c09NI8VI1t5llsQTKQjNNXzl6YC63CKaQI9W6GWJ3NxQz2
1bb2eUzPnBeOauBBizNNWa6cLbkaxFeGx3WqubLC8MY7zLW4RFm1ocm/dvF+xx4RxASSgE4AYOVb
bVViND7kfANr7mKMHcG/WJVNpXZQtwPX+yG1G2qsr0AXFQ3pV0YVhXwW/spxSRkutIT6e7WJ6Z6J
zRtvSFQ1a39/YMylMQCnihp4wuwUnBFP4oflXtAr6pzPWrZz1bll5l5dY1UnamEQ90Y+3gBasziw
mUnNxlEP7mc6NSjR5QxS1+KBq+2cR4HmQEqoZYhxJBV6s2nQVRX/4kAGbcCzaB965TYdK736yxih
fbs5e4q9wA+7zKNfO+8DleMKO/SIJRw8fnOBnlHfeaPn1EmG2BN1F0XWfnyDYM3tND79+gvXgV39
GhM9rYIE/3EcwiJ0B4AQM8Oeg/FFHFNmweDaKexPf0DaGtmywsWO9boxqi/HDjQI5WJZBGaWqb6/
SdSkOHB+BuDaDn/k8WRyq5ssolDROvAA0bjnnM/O3l8iC4OK+LbyYnj9wd75wi7iCYLHLwRaIm6S
m1QLh6L0wlOg4tEW6spJVFG0Hf4mhB6jj3N4uXi83Z1klquxJi6gC/V32UXBzeG/OfYZ8YDU8UEB
bykpDvFlsjicC3UXHZo3dXz5lK1VPQt5IC+e04cSSd8nka140cMjXHrxUG2karVoGNETlvevyFWA
l1VXSrgRUUXpq7SEnEVHXI46Vmu9z2eAAfblEmer8goVWvLD209UVjwaORQkmdYPwIEFldePi3Oa
Gu1pDdi+nRgfg3RHtK1EMoZw8PFHBn20O6BIJAfHjM+dRbXGFNowAbeEuRnVXm5O7n6Uzyx58U1q
T0IqwqImO0vHer8uPv4hCYI+Q5xtx2kztgqcxDMtGxeNPYqtmSYR+jjazwZN1LCvUYLT/PTJdvVF
QCLpYrQrmEEqFfH/1IuDTIXbeNZKkApgIGMADYd0W8Cqq66y8LcddU5ZbIr3g/8NFqffOjenMYsC
+Azv1lZuiCPBpmwMCorwLXlWG2o/rvAzPOpLVIaQrkUQduTHEBu2G/t0eNgjRyvD228QXD3rm2Xz
2ormPqMqbFLml2a/VgyG4beJAdC59LR0MZDkQRo2mBG1mzQmq44u/GYka8GPr3B6xSffMswZrAQB
i0QiK4pAcn0tuVcqX69ms6TmoLxbjWgNNqPGkvBYvRalnGPc9DwWjvlj6/8GA5E2Uhz/8RZjYjAc
0QMMfC2bNt3xmCGKy+cbErI0u4xXBUo0zf22m1M6XzBhTrzil0PxEGWdBmS0XQO5FcRmDAr4IO8A
owhPTXqSLLSYxjMLXX8rDO5mwqefnk9858+MjJvpu57zOP+HY2KUwhERbtx5pS3JXN7GFZYm3Rxl
aWgO7NVfgpt+3Llpd3wJILxbTpSQbNtObj3zIWfO7cboGwOx1sGeSmArOoaq8lVml0GTK13lcoeg
iwQCstjgk99jIFczxxHHDeS+jE6+6lRkJlvkfO6WqO5FMsKQB/uMi1GvKIotZBQBLvw16CWkM5bH
/+fjVtqhfcgJDFcd668kzGfdkqt5zqmlVIzTRGHJznCqerG5nqYr43dGEsNI8YKLi1pb5YwYqdAd
5oziBXuvzd+mt/tY1jJMcM68XGPkdSRzkyKBqWUnec2VQkGS7PmBqJTdZ0VBgHShUCHN/+fx2kj8
2rCJkqyYZBcGNih7XkSij9vABDsRqhYPJAtGWrUIqoG8u/HrvsrZ8XFgw3Ymojq1Ngan0QbbtvjM
scQCfnti1AtJOll01cGQC/PrbL/ZphlBlM5YvDEE8P7E3S3KmJwIWliW9/5FMP9VitGsT6W4ThQj
k2zww34JcnsCsOfVGZefRzJzWQGt6oCDEMfEsfJa/YQZdh0lK99de8UiYE128SR1Z/lRuENlBHMF
gMRBZeGmBlDSs/YGqOPEvxUUGBlp/Lmg8kI2m45qo+MScbDiKuHHfboQmfAI6C3MuUY45CtBIi9p
quYEZCK+CCEois8kOL2+O2Iid+eLL8ZMqNvi3M76vl2WSF2yxFJiRWwaXk9ohNKpdaw4muCy7RUN
Lh2VQ2JRYEOz1qQi74PKZ3lyiZoTxcpSVVslGwgH92G0HBKB+Pu74eQfZ7xbOcm/oYgptz0BvY1v
UHaI2v9KIgfXpGprLpii43JxPFJ5Tce7CStqj4FBx9CEYuHiNiWT+BicVD9RICHMDgWzDDrgkNb5
udCUPPan49xvDJ9sGHtyJnVDB1eBncmF/IfpVXjN+bS14mc4Dq0AnOj9XGb1oj9Eeqj6NuAymJd/
c17PtyxD9QLWlmVbE1+Z6BE/j9QOTUPBocRlepUZc4h47SfWP+LiboG5GS5cQXuJ4H8jNmw2LCdP
lxbMEEfGwR0g8qAC40Hb/uzn9jUvKor9gGbCDjD/nlU/WncaRD14M4zVarqcyBjG3bWyDTf3Ltsq
+0rOtFY3D7MIQZanJY6UnU37g0COLLcIJbY8MRGU1jupbDGYCy3M02EREemT0gUW0Aly2gZs+frb
jL6Qij8Udd0+79cg+VrM9UaOJUzUrR6VYzLIE175KIEJ1jTmKXD3xPFJTwRSLp5eGcim9T+VrwrW
JjegUjGcpjD0n9xl9KRxr01fww8fNAbxYU87Eo5HSfTWnbsrXGxIoHQWLRNSeogee2Xp10DsrH1+
wpKb3aP5gWs8f/GhIoO35Q/fMmCaWNaoV9kRCDRr8Vo3n0p4bS0lo3cyykJ1lG5oZkAtF1gFxZjQ
LazD/K3A/84mpr/KOZvidvgyTKHUe5VyFRZZHLS5lRUyhzJ/H48stgSkoptNZky6M/HfI/YxnSbk
311y5dn2MXVGlnJSs8ihBc27PaGUM2I+QGasNuAAcEE6LWO9EqTIC9+fubDOlwoIoKqE06gZN/HQ
kUy3BxD2LHAxJ53cn4wWaSVbgMYdMgdDlWLkFN7+GA0JtguMCcP9d0yaHBgGCB9CIV0kYbR84/dI
J4L5GnUPGE9fOWL78KGKYwYjBz+P4XAiyADh/HXJDybxPYt/Bd45FyWeSNTyflN9H0ohFpqbmdCB
u2/U8hgXZTygF/Zv4rQfcSMGI7wfGX+HrJqAph9connuhcZeW1rBUS99uE3wdNFvW07OQpCgv49A
HimAA9+oo+yJTjYMV4dUX/+SKxREeL53zOGhlxiB5T2096xAnSGwjVd4g7iBhi4Or/+h9F8p6Lr6
gi7J+0G/PTxMRBcGkNjJX/VfM52+0uxQ+tiVmq0z7fHCmMEWrpkX6g/EVsUhlMNLTZx2iz7nz6w7
6Quo9PLqTeTMVdexH5hFPdTfNcvKScgUsHm78os/k5lsx7rA3IyM+sXuWhUK1VapxIxQt2vW1q6N
auzkbbjMw/ghBqRxHX5qXBB9XIqlBmZmLaN5oU5x+9Y/w3nUbZe+cqSZhT1s99KxFRi2cwS4aqU9
8H8yHoQgI7ox+YTbp/eRLkPcu9nPs57QboXcyS5kNYWZN/9wMxuII3UQYMIDqwL1j7yevrzEhrW3
uPUss1JBtVb5pE783I/ZeF1wn5yofNniDfIpa4tfb4g7sEEUce7pRoOIqNkbUqVQAxxcyFxgXNoI
NVFH4E3ycOYgLLDQo3OoiSfOxls9bH6U95VZO25mZEzlO57AI9AAPUwKVfJRMYjlKW8CNdNpXCtk
/XV67lNx9TJ9LztZE5SnkflIbH60vhuZKkLGlTMdtzjwsdzEj2/TR8mVg0JsbbDQ7jaH3w+zqLtn
CYDaLAb9jtZ6QlDaY1XsJcor9KsQcyy0TE31nBuhQM4hRFOa2DFs+lUl1FPv5ViMTSpgvXYxcCDV
aLYgQvaHCWLMSPvw8fdXRRtkpvLlsh9XKbpgyp6WZOf9Gu1XAw7LHBoeRN9Oz6vuSUn9i0sI8+y6
r1A+D1fFeNkmvbOkiQHIFUOOlGOf6tH4SZwU4E3zZ3vsAZz+WVwvrT3DFSY8UyVInw33Y2uodrtN
gPoYbI2FkAIq9/xBTn0pAGvjoyRpX9jNW44xgTNARqbYBMTi8dGqynRVe1bu/Yk7aRhldyH2xoVo
fN2/Zt1ST2P2TsCOGJgXo4gTGcByt8XRdK7Ak47Wcx97qhonuEwXjpPs4wAinvRo51guRKxxfCen
Fc/FLAoLsvPpyh5+TdL4/JE1q8cMGgiS7PEyGoKvHjZA57A9OtogwnSKjNsV24D8b10gCxXIXdaA
Aw8et/CH5gYMfMJbdUB+6ZKjxnL1gxEtlCCWVamlGUNYSStC+qd4ApsiXYe0uQgKz+Zh9F+vfMJ+
XvfhrAH0cVB0PTTUT3H0FZpJ9tbIuCx0sXNTANvE+xW+IkwKNIcOuE7bAxKMtd9VgMB46SyyTJ88
q9159BVI5CHYO0g7ST0NQdz+zg51q7RR2VzIh/BhcBdR98FBerhWi+gWw2dV/otyEewMSNigC5m+
l6ZhVitKBNevpG7lR0xZkzn6sKEcGPOQ4g3Wngs22o0/7AWDM2Ef+nclK4f1neqzhjPfkHv0BrjI
bcQSiisBRkoMlaJSnYXOwkaZsrhn5u62mn2Ujn9shgEtW9geVFoZHiKq78pG8XP9cL/XrgHqrT8x
ESETOK9Z7PAM8lgYaPnOba1iEnpajhWrWL8lt7oSJ0D86k1z7NGUnUA80nQ0R6CbLkLZMJ34rgRe
GSPiGBckSqBnD/3LXg3f31E14eysSvAd5LDRBWMjOAj/CrRfxRuBwZvUulr+axxa1aMVPfidmk76
RRdp7MXVcJt+k4+ZEF+wfDz2RKLxcJOzA3pMNz7/A9JvEJOoQqWN0aagMFitwVerVmCVJy8atpoz
Djao0x0XuZUi9SKHGfqUWXZhAFlJREtawmn1lEP46v7+yp+Qpe4eOmN6Q7Wh/lLl3Ri2heg1X08V
f8/GVGM0oHxVC+7E2PX7Riczgv7wqlNk+4zi1GpklzSqy/i4rp/aG9wPrmKtTcA/M9J/PaY8dCpG
VEl1S3lwSoB2VBD9M68950vGwznR6ifuTWBVzwciuOIod2IgA0qVX1v7tj7ozMUDGdO4c3iWM5+z
St6YmToepPsiFejI7FmO1KNuw+a6tnCCHy11N8OEFo2gq3drF4dFyud6BtBuszN+57sGPjCBNiVY
eDwc9SDksk71QWvmnia7XbigiAfUl3SVWfda8d77fkio+wCs3Ife8F2SkuDMQCMpvSjuG18oM3Ad
QAJKrx6mBh3peoUU0loM4ooXKkJLEqFRxJioTn5w203q/r3rs7EWA/OdADtZmTLTX/16OhEUQMrT
+r2KiBHzyTsDUCICIvTsetM2IQZaVOgcbKR+GaHopYI4CCwRaB09nTla1WM7eLubc8d8XD6p7SQr
ps18tVjg5P3sYfOIQo1TX5H3ms3mdK4xoTQZTOPuWy9n3780d2AGTEbLI1x+JvgwoGChwOETa8JU
ypc8T8PWSt/QvLbt4/Lp1p1ITbaJKUSXoMkMwV4DRjaecRsCGQpqwENplyuzlYmU6q6ROnADFMPe
etXC+Dyayk/9H4XneFJKSj8LKgDvq0aEdrbGqBeXZNwCZBRRxpf1eW+/amxDXomylz/8au32ngkP
UXwe3QjtgCbrDCJ7um7oFz3qfRXaAniUK6rqfBqp3a4UTXCt7pS2AuaNGmAFaL8+F2TIJvzkxv+p
5JpqMae7Jy73ykAc4fjY0w+jcTaTEBBy9nQJIujKvO3UEi8klVovk7UTMBq4TXy5iqnNf3+1ICPB
+OCQFz+8V/VJ4jNk2m+RQJGqQRtc2wvUOJeH4XUbq2xdQenVMZDXQD2wpU1xVCve2iX/f1cfn4ph
aBvkXamSFbef98q78T5RLobubd9r3j9iT7ny9OZy3YJInyBH5O5MwhiWC7GNpoC9tupBwt3FG2fF
8SkRM4WTD95MrCk215DzHNJk34tGu4uVO+wr8Hn6rWPUHmIjMbApj6g4sheHrvGYoud906pIL5Nv
RqimTAS61fJdCl1bxd3DPFeaBkaGu5RoGpQiQA7MLQu3h/hb3YQLFsqfdGz2P28PLvB/U8P1IUc4
q6wcK5gKOivYWD30wZjnmhxaa1yYs+2aXrQ5sZ7/XuFdLqrs8C34RgcpznQux3suP/JIvO9/FLhp
q7JhbofpmkeJn7h08M/udL8nfmKmiUnBopHd3rSkp8w+ADbm01AD/7hCnygMBjWr0HbsiJfmmI1M
/aIjFf6o3S91jOv8//dU579QQ06Oq7dnV76wX9R78UlIFn8mba1ZOVLfjgekPcNA0e8yXsVhMAU9
0oeV66KmKV/Rt/WZniprS9FjZ5+TWX/+MILhC3yMPJZ1ts7t0e8xjiMaes4+uwRMK3viR+ebRyLf
erh1x+CpWBzh3fhb5HjkpGr/8pVgzs3UNiyDGgqnyhiNkCyDIQolVBFmsjleDNnTHU1aUH1nmQRf
0XDc/gprwyBK6UsIsqJCD5NmDl+EH3Xv4FYhUntcPsm+SEqjHZHcuJyjJfKUTnGW+18iQPKUajI+
xoUAyhEhgB8YM4T3t1lFR0iVrnpnNjZta/Py4TQ3KheMhn1OKBdauG1UshWk9XwV/2D+XraFhxaS
pFYydPmKMBV4fmAHbh0NuJMqPlma0VFOue0MNRAgaEY7TielKD8xetBcBcJOF66QJ0fCgAR6QYon
snIlzeLQjdz6mnmrlgyD2qIwcnak28tY/vPOUFh4Ptk3r/wtXRJgn5vSBFhq07giKe0R1GMoQE/G
NMyw0QAK9KBC7P6u94nYAWGXafVPDJhHnCuPNWxCr63vKeVv6jTOmljLZUNQuEaPjhILK3W7+VkQ
focXxZqQ0yli67vsKjCKAuFodhyPGWzvH5Af91cV/+7hrZCsIfeUKvNqOQYsTEahnPfmJF6fu0Ry
Rot9BjulCFxalr6Qzq0NBHmmR4HzzPyq+sehUyhmvhQk8YI/KdinHIuBmab4vUmZrkMTVWIu6N5B
zMMAc9bg9GiE8EM9OAn5dZIpFfuQYaGiwQQd33p21yRGfapXjg2HGL/Wk+Z1jMfALBm2KF/YRCnG
sVxjULfyjPtd8ls8GJO9ywPJNcZ6Mz3Xe8B9EwM/rabGe8hb3KNEJvQU9o2J8Vu7uhQhyxnUkE2t
FTk25zdN+4nnDZnXIDmKIWamHFyzmp3hh4BlNFH2isSbgLmFqdqKjhpxFoRltT4anuzQERJQa3BU
a74CCwJ++B4jS9IDH7pfk8+8pUMxeUGCQa1zNRzoE4FH8M/dBDP7egQhDEYicrKKnOAr9IWfb9Ke
XR4xBo/bFyu3/UimpWQJjcQhkyXVAmnqv8NpJkGH6olB2xfQmW4KfdEz/6AGg/AGQWA/aqPAi2bS
cageRyFPGO/QGrrQ0PHfw8QaLeE3Yt0Ry7gz0+6C969YhdYoBFZMnrRpk9/lwMoOB2FjFxbYNJEa
qr0QZ19EZ79G6odsCWFE4gaoFfKCgw/LrBYbgbw7ffBqJNXKWTKhuBLFI3gTdPvuG8keRrd9K93/
5+UbBwhv9B2RQgzhniu925Z6e4UXJWpcYmoIkFx16XJOUyXjQ2PeXTtBZz1bHxQ3AS5WxjP4qdV8
g4XzWKU2bGwx+Lk2LvghGc26zfvnpYiVqLAQ6HpDo24G9w96sBkMB0CrW0ohXCF7oShSsORSxVjl
lPRJ5Ub8Z0kWhmAuhye0WeLqRyI/5bdVeZ0ikpxL4Ez9A3dpjXL4vjkzmUiT7Dgg5KIU/HJ3igl5
53GJoC83FDbGU2b/HbYTk9SFvvi/PLrgfiYkdZYEQroIB9NAWHCndeMFZjMU0gGokoBFgIeYyzSY
ZJK9GFHTJ8ze0DWnUt28Eu806A3tyI6zTQSVOfhG5HjOIhIko1g7EFCtZrmfVPt9T/ahaUiYh/e9
NAU9eaGKy+s/Ehmus9aydI1+SelimCE6HG0LFsQ4hdpMmIfBjD8AMusi6oQcNl/fS+EmHKlk2jNg
pTHWXaf7W48PVRD/vG5mt4sKQasQipgsncxhCL0ZuPBW9Xmo246IHTzxszimDhAmoVIMy0iV62TX
y2WkL6o5KOcDY7RImXAdBRg29FXoZ0LvyA3oznoWyJWYK/zegTrdiCKWdD5boshPzHj1iVBG4TjY
G7tl4ywQL2Lz2EBj270Vy5goyp0RIu0wo7ozb7J/kgmEZTLoupmYc7NYJrU6EhL8MJ6oIqCORWZq
4ZBxgB21rcjGvyNZNWuUsXSmneqJVpV71LkJMfhi0qLoknlz0KCdInD3otipBC72ESpUeegCJAKh
B8H78aocclaCiRL0cwO0q+SwIN+P9oAQspkPukDUdZwu6X+cQIpNo1IamHICLW90O3iHzEKB40J+
sz/ybduESkX7qd8TcCxLskDc/Y/6+C3xZScjvxKa4+GTIamL7zXFmB68bLCRs9D5J2pKNKfZrYkT
owu6NlvrBCNWhjVFeZ13xc5RYeJ7wGJ6AlSk76lA0vH1Syx0ailKc4xuBtttgEorrTyBWpf7Ms6x
1qvQ7IRcF9TvE7oetKePL7U3oCqRMF1V+2eJhYBzA+XHav1pFWyYXzzNbADNbqJUBhimf3I7nlfE
gdJX9t/dcphJS+cIFjEvh9ocTRLdjqecaZ9ESW6XjdGfuEgenq/0zeEumsobrr9iSBwlFZjPwVTh
Btq0W6yaGfn/3rO+Ek43W8cIBdiA+0IwMi606qL9HbkLUaj1gdui3o+3o9Eef9EFvAoG6+YM03FL
+94pbVwSN3ymDKbsRJQoKGK21Jw95t4UnlrMukq0wkSsEVUiXXDgHrJnZfubwARQSUyikSGPepKe
6TMs6pZp9AUn7jX7MCMEB76AprfmJCVQcCg1M0xFLBnXJ2OFjdvmqzoJmENMnFbXG4iLXwmp1Aic
uXwPMDkBJ7DADUsu089ckmVDqH8vts74eJb4OUM9mnVgaDcwbY5q44XTS/kDsbEysPqeG1iodxz1
/+JirCgnyoMXUSwFfqcZYXJcKmblRqzN35gPSZggeXWhCl4ru9yFujtxr7g7uDrIq16IuO6hR6sO
xcuK4i22aq8vatYjvyQ6lk2J8zOGoxrkEd57MccPr859fDZgxESO18BtgJ4lsNIxmf+0xFshgTg6
p43znAv+wmWINqFwfEjXAg1IZmrtv+qELu4XXdHGA0M7aPYEqi699anQkppKTXImkNvqi/+qUgCk
VZIk7OnAY5NBwP/UIfmII/ydeKE/+bQFDet5VWgwONVoMRh4HTFCYzcnlAZLl6JXA+ou2Bhuv+4N
jFaGePqMhjvpvdR7OcHhXdbxaybKvjBnbPwz02cW5CKb/nMcSfkVOBmLAl93MNlIv8/sGSY75rWd
IYwcN6acrfLvOyJi9zxBxQ8Tt+e/k01VmkbcfZk1MQVMu4uLLzH1aJHh6X9iMmCA63EK38MhMin5
4cNZaXyMQHPpZsBQUn7YgA2bSJITaSRMiEchVHysfar3fRbqklWtq7k26g8tqg1RoSFUQ5W3MfvZ
wbA/hNvjur69r33fYQy1G1fSwZTBaj6dgoREOu3JqPk0ANvRM3i5/sL/LC7QGBO9CaM8tgQPPZGQ
C1JLssPGS1dThkb2rfoQL04JyLmdrbDjux113zFZAqk/vAPkQ33vp5oHXPUplXgawAMtRgnlIS8l
PngaZl3mv3XhTVHDx5806qlM8yMH5FOLG4RDP15eTalaN8UMAs5ZCxZUqZ1zNYw3NVcIkbI1v1YG
AIoVa2dvUftrDxDvLrKuNpZc440c0k0MDxEycPDqx0Lg1BbXWPOs/MPxaMBC0XfFaRkx+G6FTuC2
ijEflUTzgz91Cp9eg02cW2dfUeaC4DkrrVu0Xg+TbUKo34i8mW632bVLLGjZpM7qUrWBElPrePnC
aeRLScSBfDas+x7EG8Pt0XLkrrgHPQqBijHgMC0fet2WYphfaCiT6ZlbmovqYmV/vBTqpqn6mt/C
oDAjOglWN5dBQy4PIdh6QKFa9lItCIPmq0xLD24EbCj4wVGJPiy/jJwtWtqylVZBjcYcpzS9J2O5
cE2LGOrKdYLkTlL9UuGuTA3kErOCPnI+4UcvWgmBOEaIQP+uSdCJiRwv6DW/8zpaCRGGgTGWDaYI
qaBwsAx1LFxAQ+Z2soQQH0n0ChHCO8yOlvn+JOXdxsFipwLLwIq/xfumM5o/iBWh/ZUmdBz2BAYB
dVP59vwpyQ8Hg4N7/VdWCoPOlbKHxE2OBISErhXn9hmZv0Sai3EklL3Z8YS3HIM7LBWGvgU+CmO9
BAwWIct5olxJZjBmJ8kfnX2mxRQB2A2gipk4kLd0XAqcx9MFgx1PFqY/zlqdEA9wBHZswVBTQv9Z
gxFxp6jTT9UE8RJbVPbqWuE83uPpTHdv22DA9KqVUo1Pjtv3CfQy9aZOl2Fb4Gq0kjF68DKsBEVM
iwN+3HUfwfv8qUho1dkzDjnjoqOK4zhoHvhUOwk+OmzvsLb8xl0Tn80QK355DBYY8iT2aiZ/54NJ
1vGSogxnEXOhdf4kS7BhnQ7/BII64LItIod249UsZp8MARkUJTTH5w0l+rAwpsls6E/4buA5b1R+
kaUPrL03QLGXKgDn7oO98y+BUn1whZfaPpxPiGP0iJhED4tkC4SNOpGDtAQUNpZf5bYmFeQRSVNZ
xRJd6tRNwEMA7sVeNUCKSWuEaARwBZnpHho0FfdinElNfLBMQIw3Jk2tttq1uBv+o0kk3y/R9C6M
zgXbSrQacoLoDs+u8iRotEPHVsUDy6wvXpaOMdIJJlLqkxWsCj3JivEfbnZAKglAg3mc13PqlrBs
yR7LVXPoEaPcJRyETSiSeJEOJiNSawchdzXbz6JB7MRrNwGW8rtwGHjpBFABddAZVGWNPws+NwjM
8JmFN6o4BCEc8KIABLMB0PgMUF4RbnOpFL6aqtX3mISl6/qAOKFpUFJBidyOIBuKkTQ9IZZ9JMHg
e9sLoPs/nrC/tUy3ozrYVB1r2mAsuhJCZPsb7IAdaRoBOLXDdALMsdB8ohROrL34EOINtDpW+ucU
RSuiXwtNJjG6yxJ4TOiqgpjltewYM9htXMs002hgnvfqQWjRpNt5gC6RSXQ8GjSswRczHUDluoAe
qJ2Jyq+eNWVpwZKxHlFXeaLHC/lWmO/B7ZuTTXA7sefGF1pSArSBBVMkfGYYit3uvU+7On138lmx
GoNbgFk0LV046bGIid31rmqX8ZzFntsMH0o1EMQ//bQB19/nxm7V1U8GrK1OuujxRl7m14Lkc/Cc
zkQ31g8FRGInHa+9uqWCQXC6BXaW9LrOD82M8uRz+L72QWdVij5M3FdE2yN8NY1XyG/mSkZn+OVd
AraTt5xkvDQGQ3CVgd3T0rNa60DF7djCPLHHFjzMo07ZOgyFC5lsV72+7sNs41TVWH+t4e4u7Z0e
RNrE0zWJcPkX86NwmmgKtw8PqkQQIMB0SR2TECdtBgMTjM+C5V2m+rd65HReAj2BkISEqpvnrI/w
5WGminXscmmm6T6bHHwj8X9VDqMmHGZ0LgpUajYJWBY0x1Wcg/dGLCeb41sgojL9pF4M4VayrThc
Ws8QOQ7ceqVlBAohupc4SwMpy73iIjW4Lfrc/f04ycUjH9D7CKl0JRg/AM91n9luEWcpW8wQ10lw
VPjQvtSEbx4jk5BfXtPbYjfTUm60sUNg3KtMG/ImPRVd8ZAntNR+WHZSXPv/YPMKjG9FCv/3c5Dk
cvlznGQ5oEW3FA4sAqIBgeU096kUA//4WWsh1V7hT/1hmj1LR9iP+fKTNGsfB+CmJNWEvDcd7Ntv
AVePVjuAgIf3R+rfJudPL1umzfgKLzpsYA7wYPBCeNj+G1bVZjCcWUieKqmorQDrNpIWwer/i3+R
MQHrShDeMtgXPsDSSp2Wa20RoqZDPPZJydD/diGWECwtECqk2hsxdf2Amkp1WtcgrF2trtCU8+BJ
Y3medWKZKWpM5DDVVqpIE83iHXfbOgiXwDcnORQNMHuFmDGxO0hQnsfWFmlAE0XdZNhn9VGDjgv2
uEevB2t6yxT9sOBXYFc0fLq871StBfpGyoUE83RjMrIyWweKdd63cSDtWl+zpT/UnyQ7IJpfVsoe
boBHYhTjmmKnsICeR00B8vkGJq1oxY08z8HUyCuwipdeZ8hLgPWEmrE0bI88oWgmf29Vx4B2/qb4
BeY4aOeuyEQxAVi/DQdcQK95LTRi4tRl3o0S9Apx0hNx78hYOFDaLhjhKWr7WRu82uXeilZICWgM
7GziYZH3X1dGJvZqJTL8jZUfnlCo+IAcykZfHelS1RLZaiV1R87eXoOKHhL9DcCgVJI/PHOJW7e5
cHKYMANhNmD2YxYwDy+abpd4WaZKpXRFIpzDFdTfrpCCms8VfsiTy4evGFw+4xnA+2dwQg0bwXjZ
1SArbrVsI7bJIu8TOG8W53rpT1xvCObDjWSYFT74x6oRgmFlhj3Wn9SX3YY57hRK+RQ0mhhMFKZf
EOpneFWdMdMFp/6ELZyjVFEG/bgl00fDPW1R0vxC0krcdO/cYUsIvf8XnjxITgnOPmPIEI1AJoHz
Qhu5gLZpkKjGIfHWa3HiBnzRA35tnlyXimqsT9243plNupPIn7qtbS9yQuG+iOJVeFRVu3/FUaTV
x9EWDM4ONnWWp+3J/EUvi0AuIZisQilxfPw3W9LxKC0UgNdxlRUMquWGBAF1l4i7z7ZNlytHby/H
kQ6GU1MmhSCgBYlQqnmUUKt8Q49FHY2e15kbjKldLQeMTYainsqx972wRvJxZ1HA9KmXhQURxiBl
sOU8CymfjHv+r9SHNgnlN+YLZc/IaxVuWQP5TzU2Bm0wV2k3zBc4yQDBthXYagqlEK/QTZWIKUiz
N5zlDE3jftZ3Tn+ZOTqNXZIIc01gmpMCqFkgjj2R+nuZIgcKe8StqB0Z1tQUmlaSq/xnAnzPgxbW
rRF+GfKHZwnsYknmzNdrldoKR9qFKmOoK/lQjujp1aLP2ZSXMH4UMvwZVkV18sV7d/xhsOaygoSH
LP9V5qDjLujY7Xg5bJoDi3p7PsaD4tUSN+EICb4uBAwEWfjkwQa2QDpjghKPKyJP9DtqxuZVXMVL
MC1VIfYJjinTd1YXCpmJ3K5OeKIiYk+BQzfa0nuzacusGNA3hOGXoHO8qT4Ev6ZgAlkb9HXVhY1F
j9tlkj4NcIOmh7rEbmjr+MRYYjh8AikD2jyUo+BrP9pFjVaJeeWtdpPM71k+QhaipG6i57dkhODZ
shu+AU6lIuxjUF0+WI8AROW7oan5wKywuxRSl4+Pnc10H85ixWjQvo6vGVdQSUpEIAe+2zlvwFo8
JllzUFIa6qZbzyYY8yBEZuM4v43XmH7pRFoRCEeYayqpK55VtRqj017Cg2WZEiXmkdP2qNeiJ8bO
XTTgwPzWSb5xXdH2QA85XtEU3UOGeaMmTTdPGcQc4nTsBWS8PtpRZ5jLpIL5jCiPFFWzKf0XZ/Z1
txtk3oehxnDJZce9QffbWHPnSQQnIbVlnOM32bKC6wS1oNcC+biPZ3xGgmPZnZOX/IIy/DLykoop
2wGHtHUNBwPmOLm70nJmSNH8oSN7EE5XFUATw8UQa3HX/wNhaSrDcMyQC4vSWQNVB8Tb4dqGJjbT
5W6dLg45+jeLAiWoLhsPe/sFIZX/dAZDpwiPutO3bbAh01fQnbGAIkLZB+F6l8e4fg23LpA94rhh
pLLHW4sLpZeuCgQ5h9qKZ1j2gRDMv1GOPiZmKs04Vpex/yvk7Qq3KN0BQztjbt6XoLsQkM9hksai
IbeNSgPTEx9hX2g/XMI+eNBdr5Rlqth/po6P/uEObdZ+JW2LlfFse4WQz4b30ZT0JNCv/IWrZtq9
pHsgYldQbRE/QOE3Rn+UzbVOGuD23BH1b2YG0oxLAyu/qF4tcm2qT8mX0AxHC05vccolqSwSrB3X
oiCSaMtJlOJOQJ1N7QpMlxdQiQOhYLeDab5ouY+jB6+jaBYyP20s5ZLBayzdg+tyIkjgVPNsoxT0
4svUYNYBPbH2U7vzkrYfOR6yDleL34kRrh5iYT7k7oy0d2/Ml0svCQWbmjCOm1+RjyrPHimKJbnu
ouxh3DTAu78u9ijZ5heXK1SwiNzq2cg37vN+TUrvoaUw+9s96V8cRcatjpFXJJ5KIKflOI09inp1
WcSymoOlVhGZ00sMZdAz50qKDe7IKnUP+NzIz/cykHWPJn4HqBBaaUCFmSU8yP4zaG7vLybk+ZXL
uMU07AN948GSk9pPRngWKM4MDLX76qJr2vaRZHf1BkKOjZStsI0V+ATw33gNtPH9hvffJd3UojW5
MF3W/qBsMMxbdxEKmHTxaf2Win/tv/DxOqkliN6dCA76LW/xR20NH0MAgwmthu9qwtjoAA2RvYva
S8u9dZxdI7EgxTXtjdjvvTdIJUP+Ay4iRfBKhtuTkX7FhoyvZumq9xk4+TkeXljxWIewtzt3/ruG
HabZxiBa8cdpKxftSy/lKnHr7o82K1Y8aaWzS6qa9xwvZ44E9v2iZ0gvXXlVoegbRYfOc464HQn0
McqZAim2mVLAEcVHtUQqPjyQ93vYYijEBs6OEhXpAnCcJtW5onc9dIiYOH6tXV2TJ53V88UHOSJV
vhx1ZsRWRHWz58h150E+bUPIDHLPzCq6FVLofzBScRN7bjXD25a8R+CfpQPKbtoZSIfkiJ/5hqzm
YHw6urk1Z+iOPB3DaTFSfKQaRAmVnI5ycUSwiyTpSJ0tVPMbilD/JzPxInDAjyyat/c7ouMeV6bx
Tmqd4VSpZT6NgYFwEPy3GQTOMemmPG1b3MD4t3P+56adiPtMndjPBu14GkcGTTEw/AqEiR1o2IhE
7maRtRjCqCZvonkqN0FCXQIzKb241f53vIXT1BLhst8beSqOX0w71Zsrm037A3O9o4L6SabcOpeJ
R32HDcqwBNCsA6H3d8+cj5RVGBPhk96nJn5G3qYjD6NdncFdYKBcgLrYJkWFcmtfsCLNXL/8GBAZ
o8piif8MZazJPbH0xDv4t/hnJc+3NgESHPOSbevUDv+M+uIWKHbspVcJgTMcoJGQLJuJFhqs+cf8
aUDP28Hbmy8OZLi1wRFe3lADBjLk5WoKBEgVOTbRjOleJI1vT8QCOhjm3v2icGm8kWEvuqkPbe/s
M89sUNxTz9qh7p8A3ZeP7duudyCk5Tcgpo0p0G3vSKYTHJJc7rAWiPWeOF20kqPoEuv7ZFKcuqcQ
OtIinN23R49clgZLUJVLBMg+zcW1lRFi8xYmo1Tn5QsdZKDSTEsPlco0Hu6uzrrw9fxsxIOF/LYL
jYgN6AohIoxmpFe5mVyP0FZcKKJ9sRHh7v5agGWyPouTdrqIGtPdPFRRkKrlWdBjXF9+srAF/la2
98N4ylZQWf1k6rGDkR1gXYF1n34F9lHG+Q7Abvj7X84D9gAdRbG7TjimU5aK8y+dXJUuMPDS58aw
KuAdOKq9M7EFxA8L76Ca1xu9I4n2AcmSftvis4A47yZGpGcZutzw5Jt/NCxkpUWiXa7pxGRJzymK
LuN0JIhWXjyxAV+WE2JYY8LUJ261zVB3K5Ylbb58sPWebciQ5/j8Gm2HGskLXpy7li1iYG7lzX2A
iu7cbiIR+IA15MMKdiH4T1QgcG2psq5zA/ppQp+q9g2tPTdJ/ieXYIN57OXZAUl4vw9CLDDWPnG+
aMRN5lH4A/TnLBDOT5OPCfIFl7WzAYzki4RqHcBeBdqBH5SnS8CfpIOoHNgy9F/3pPKFA/0yJWdD
lt0VVViEHKbXna+KTCCWchommDCMqx8Y5X9OqTMeGCOxWJBCf6UaecEcEFi/ZIjtdWNoCrBdxFSx
7yGziMUVi076haQs0s/AgeK5x3bZDDcR7rNvmaQZXDZRAIcoRg7UcWx6qoEw4PE01VVsSfnONYSX
/jNhP3HWGd0sar3jtSGe18JgJtwRiTfMdZ4xCUAENauN7saKJxkbwM/pa8N7N5owlAwNllvHA0h0
kIvSFSyHH7nq0HHWNpO3VJWzceSQpcCqJqMWtM4VHokhDnpr0N1g24IVh8P8X2UVVt+PysrEKkcz
dFIF0a9iEtu3aOEBFcWGT/dfSLkTnpVeqpU1i+y1FiZpV43vYa3IZMmPoJbQtjTiuupZivEPayIn
+Kq8b5gctJEpKGnekPCMMqtoD0f4RSlW9AaGX3oB+xl8iHK2HbbLpdjF4YCBqHNfsYzdhOoizxW/
NRfnFg1ICrNmrWlJbh/ttrzjhfP6TMs4RMrCODFXq8Ti2Vc85OIqj7PwmHv/hetg2e1wjqA5nDI8
K/g3KA3Wqw+TuBXtZH7tj1Wky66kxmt5TrP/CYQjEfSMIj297+WwZHnj0ZVcc+ihFy1aPd4oJ50O
jFBofcAk+gOp3vXtA/RuRf8QHCtL+jGpUs2tgUKUf5mKaQ7rXipkcR6OtV6shLPABLefkCor0zUB
htouHqPjMbvX0xuj7oyyXxg6Pndf/yc+zUOVd5qqJqWklM1Xvodl8PVDgFblzwPmSgDoAkrFo1Cg
LE5CPqUtScjQL6aRp5n1dXySMg10m/1IoT6/rdWwk1LrsvGK0Z+S21DvsUfKYCR+NIBbzDPuQwuh
DE5hk2Za5/KA4kPahncpDirOBXMnVDW9t5AMoKyZUkMSECeVeVhHlZLGsyXgAWMDoAKGJpvPljXA
33YW4Z8fogYQxP511Wp41/tb2EzhZ3wV70wv2HwIq/mI1UqvFPp7msX/nTzK8g838Yd4gHy2fAGi
IFxsoKPtcs0N7DMgV4JHN/2yRMlHJdzT1vehAXVhKycAmy3s57M8/mNezXHEGY1W64b8RJ2z2r77
P349RPwv8FSMUbEzOrkGojUbMHxdW8LUhLAxU4bj4i4McCPDkz3eCtYi1Wc+HQjf50rw5e2XHa2c
jEI0aHxaykV7/BaSoftUyUORkYCFZ9QputVIMtpwnWDvtTURT4SNXWaDlwOBSplZ+wOxWkxO5RrI
NHDtNE7rtBL7029+aZqt2E7y+dDL5GSfxa2FfAXCxc4KCHIlWZ8j8J4CMk0AC0L664GvN8ud7oOj
SzWoL4Mn+fj1yq6MbC82NJ8rDu2anxP19vG3xc60zSAv75QE/RXAp5CWFuM8Xgi0e0lglu1vSFAG
aP/fbY8KBwjN4dX+5s7UTz4qbdXwKiy8VvnUoquYW1+xkS5HOfNmXkTf/n7jlykvt7JMCeUdw6T/
MhdImsDtZHMHIjsij5biCFFAGEuFWwCPJMd/jeTMWUCg46Ut6U3MZstnKfBwkjxd8I9Uvn/A/hlg
1eVDubyPc2njQ231bq6ce4c2aKVDLkeI038/VgAyfdKIukocWh40rSVK8rsOOw3qi6g=
`pragma protect end_protected

// 
