`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3824)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPajJBURzf9QNBnvkEwdAEowuDbvjI6JZaE8weHIgbUb6Y7Vo/NnHA/Qi+
UBuliUL5EXfjlmXcrmNchzY0agtBpr8ubW7lI4HtXa1PGgLcPnA0ObrsFaMGhIC05Hgy5Hr+n27o
9LjDxpgofdf6rHk1BOqV92v1UaM8NHOpIM7/U7EgRBGNtth4v1FWxT2gdMMghvFx+x4k5HL8zqwS
0hjbqf8op37WdRvtFUSLuRpL0P1cWX/hzb1NdRRdiy1K4RLXBpCh9VKK9yBEtiQ5UUWshSEPufPH
3ubmXwB51rVLZkjbBgZmdB862BUnlNlMGRUh+Otj30JulYsc++5ZaoPqz1wb111rSLiubHZohrCq
eoNYIL8BbB/IL63KCBquwEkIMc8STHI231NKNRxWMls+wnxPQkrRZJXJ5oIMO9cMqeDfohtVOVaR
EOAZzvMhml3rbXpEmPTaDSym6N+l+BAntClpA4GoTSbc0/qHP5v/uWi60xyq6rMtCT8voh3qmF/t
rsdolvFUvgO1Khe+nS1E5lb/7PJSEHMkkBhEBKiRDxdZL5jAT608OBNLr4nqhIAMu3/hq2IoUI1h
bujmsaMGVp1p66VJcNmaJLigWMJOXK4q1Yv4k5Xp7QldgDoA/OXncwo11zGCiH1O4Jl2t6hG2euA
zVWtq3AXkkwxMwCqrYoudD08ROUB7Z9wYHBBfxSliQBEXB2s3X25gUHDrJm0qoM3xInYLoroNfqJ
dP4SJ4I/x2tsKt/vxP2rVl9T+w6eCPxrqQJRHrrKhpbbPRmuKOkgnwesuBCuKRuqOsGPa6s6G0Wr
fnKxBbR09xTUPoleZwfsciXejmDAHlqFCEKbTisaNBkUdHsJ8lfV4Vsn0qnhZjBXNVimXVWDkhOU
oGsHgj1HxQO1BTHv/exnj2Vf6ZkRW7N1oFgVngjpc3D0uXwhFZ9dWIyC5Ugg8bTWH9HnfWiUxbSM
4Rra26FUdYQV2923D6dDzrIz5q2xJ6MAwVMvauW1PL+xuVwgj0znNLRohmVLrDbPy32elEWbVxfU
cZtwAk3WrqJn/Mse+XhH4rHLMLP2ct7MrZMgyG1Js4V8r8APL09E/FKQqvmDKRFt1UbIb+vBdZqP
7RfBejiYjRw96LEb/WjhkjJC1BdanWTjzGwua4ec+aX9HCzuX3ehVgiu0GyzpsJXDeotBWrm3cmJ
fgJ3ZWebY3I8WrAjBBtlqlhynYCDLT+87j8dXZyr3iO0uor3NmLJ1ZfU0T3rcGXkrgae1HWd+LRk
c9QoZXAjTso/0F34n/XB4NpJLqxBaC3SR27Y5Pp5CBgSQhFLhopNsJbU5vBD9w9iWrHnNgFtO4E3
IqE2P7vEVJBDHg6iCWK8abxeKiKornCAhJM3YKLaWWDzEC9MZp30Wr2ZoVUmeVC1r591ENglZHOr
vQrlxU4iKkXdzWdGFm8ymZ3Kgz08V1qLG1LPMqQta1ozaBE+vl8dIRyd/iTEUU1vGnTFY0RgCwOZ
knlvm456MBG6kmjUJauW0OoMW/virDmZb9vKth5zS8mvDR6xOuZYzJHnvO9RpAlSPggqeavKAJhT
vl66+PwGieZ4bbXethzJyqez01qK8st2uwHvB7ap6VDQYdfqrB9gsFoYpEeumNp4tQTwVwnr+jz6
3gUyWJfLDXv3Oh7Eb+M7PbUVYffgj3t421iFAud20vwR+MPywl5SThHeE8+2teFL6eB7VbxhmosB
s2D+tCsF3H1KQql1nRTd5Del9sOwRpuSc8v3BQTwekOMSRBqq19VsoZzhpCaQAqzHQk3k/KqGPGl
yuScE1AjUNEPCujLacOE8NXM5slp7rcgAqSOUi2mMbVqbq0vUo0kE6+GgHyZErjcs80tlMq1I2yb
NRuNFHZzAdH9rehXRkpdVxS9HjfeZ3HXupublgkdK//4RaKLlMhSVGS/NqBjkAn4RJK1v7ZtdI1F
jnqEW8cuQWQBVJBny/g6PRMQpSSycs3cmgm+1pq22eutCacDhSz2Aeukc0mLyqQqDklbyeBq1fo/
n47g4WZihSxtoZRLh32d1us+lzUk/DecN39SYqdLWpLZzuSQ7AJ7HPAIYMwqPX7FFwFTC1NXQv/l
s9eIVjNMC6Tz02ksAWbSkO+/0y88bm/5IXTEszrDtZkzgnwnY835OevsSN05A4tqRX66hZSldJ/n
eNwx3RbZMYQ5f4fAGr9Cez4LH8Fuy7q0obdhxlVdppb2D8UlyD2E/1jI1nJabY6qlerb3/BDZPQr
tlPeqEQU6s4YtkVjft9UL1SWwkkyvs1nBnFKjyt9eatxyrVgfF6qe6bWz7dnTBw02a7aux6JgaZJ
Q68A5XAvSCit3HB5OehBELDGCcK0kq9rqmYjhbaCskx1slraJmpyFfhY3PWAZuLQDXOyUs1+/41N
LLQLGfr2Jj3qQ6ynC1DMcn2mrH75+fxu3piZVAuhGKmHSnms4V/khbw/Nk70vgUUxz6f4VypKjos
naaURGVyHBRBZOILkAn81OCknovxHH2ZCOXQ2xknx9EbdlXnGwbEV93OOfSXhQtxSZ+FoB3ufRpZ
jycTHvyUPp+KVuAMxWAoS3qVjWoALoE66ak3F+OTjvdfwAvp9389bdNichfE+NBdAl/ltD1hkbGM
33WAfVWw6spWkXms9a2P9gQFhsi9ukG5PQI/2vfVVojv9+XHFZfHIva0BcxJCr+xBXfR7C37wYYY
Jmt8Gs8UlChXO+7pXEjfXfpUnf6lnIm1XVHR39ORAPwZmi3zYHwe6/z5p3Q6ufRIFNbnGWbPHkOg
X+YgJ6JWslHe8hjYxEE8vBp9b9yUt1/F8HzeS3By6PPU7hexJEcQny35kS7wZbSy4dYbicPlDKa9
2qANkRr+gFCUwzLZSkAi/pHOXDAM8VADgbCxQ20sqFNgmPL6eojgF8Ldy89YxSEipimNONzKPtvh
PsF2pcCi5vRkf6WBgfTkKyOcCwkAzivxBEm8brxRq1ZeA8CVmb0Vxd7K1UC0R3kJno4mCXLesQ8D
4Tj9fyVDCqCmCNxhQC02lAfThdZ4VIRyerKkOo4Ez0DEClt3nlB1m2udVKukrGVc1ut2tG4lFCPw
w5kaN7LcdcH2zKG0DfHeFWILn1KAWHpTeW4ZpDxKc5g8LxgPRQCa2YsUyzyahm/LATroqKdaAjhk
eXt9TPfsF0PQ8CX8d27fF7d8QX7NK21OBzQZx5SfMqx6CFwh3U7u0t4+FC/RDgjtnpVOs4AA2RJV
tse1woOt0I/zRr/RdpFFCzig4JOqGVfbYDV/Doren96CScF2de2k88eeC8a2sKZGilszHG5S3473
yACbgOLT9x7pAi+JiM4JskuJXQt+dSgQ143UiirCh/3MRipXaSFTFA6tw81ffv3034AXX/qXfJfG
7M2wasi9bQ1pshg5IIoPQYmJxvI+lDk5rYah9GjMV/XgKyTDSMN8H3WC3VS1hmDlvouL9gWmDmPw
xtGbxVloecB5Y+qugXmHoNmieImrexczW+rEmcXGmAHERTBnXx83sUnE7Bd64HlCnTd8IqjQyXWE
hZpqwXp32PgR+iPqj6FLtkX4mTEbd/jyj4MO2trGlmnKkotcWMr1YY6SUhch+I/6/f9Zwv/5+IsP
X36TLdsqEYgrE3RxWhE5rT1KpiDe6FJZv8ETkPmrbVdqaDulKh1i0Ua8jLUkaOE5kWX0ww4qDscz
vppRiNBl2LYelOQpFzZouKHHb0Sc0MA0hqBXEhT6dXbkY/EayKLB53IYfZ8VZtwiXJN89bJ7tg77
sf8Qu52a0cMxfG3ku8BoLmzgSdQQw5nTWSoZSeuzy7b/4WNH9+SNUqRz57ezNPwV3iWUpjx+u9k7
l+CsrlCmBl6jn4oTIq7bP2+/oMJJdB6mM5KNWHj0A3GOhzF6owhxdRr85KnDc0DyxwbXPoUiG/hh
3vTkvipFP2jI80jRpUKCUHOg6sw4pka/8aVimNm/i/u52LtdkqtXhc714Ff1k1Yruz72EZjyiEQA
Hfx465FFHRhuG3QA8768/TpRnTYlce8nmRwKhOl5sJUuoqbITPrmYEN0BJvOHZBG+6RE1RLmQ7Di
qj3Cc7PzWJrAj2TQHViwBnIF372o5L7pAeaQlV8SixEJlpYHqwyEWHw3NE1Iuu3gh+AU+P6fDyUp
wR0yUNeKm3Q9ARL2j75rgO2ykAZYl+h/u6k2VT7448ZxcgcfNMv7K+LqUacxhMu+SsN3pWuF2gRW
vIqaaqc3PEfHKIddQ0iFY7cQIYJz3qf2ebBK39mKbUUl+AAW3KKzf9hEQGPLWkS3cs5FOCv1oMFY
0kf6X/IHY9euBHkvGuSGJ4DEo5PgRPQvGnNtZlK7PYLFL1KHuAe6Qro9oOkLYw0SbE6/nAxdnVCL
HveybtH9i5XnOHYqySAzncQawB2ImD2OZksLD6DS1K1iy0JEOSieMpyWybQV4lA5/7Wj8SKu6c5n
1oaT1RovGj5s/ktvxNyApsibXJmTfBSr5ehkaxI0AvrlZlZIMGNXpqiQyjrs45BWA7U0u0Sy2gUN
sNXL2NUZzCe6jS7msxFC2DTlKICb+qBnyQtapPJUDFq+9uE+EmzftNWrugE197wjRKO5NopHBi8w
xlKnhkzXVCmj98aOb0LVy3l0fGHqlca+P9eS83C0sbu+SiyzYpaDKvMKn9do64YDkfEg8kMFKeB5
vYAxHiYi9d5cWrd+GKkCJTF6HOrA/M0FbMJ0PmOCj4V0Yypr/NuFPpPP/AM9OJYlHfUpCjjx8XXA
KVAsmuEBjkrl+gD1FquWtDz7CXdPWmA0sNFav+J9G6M9EgSc8c373I03gztqd0RqiI8wXjHaQXWO
NBO36aaIXa0bjyE+Me7Se2oDf0wACE368w5Ov08tBnTguqFJzV1PuR6pozkIxv/2DjmRkTfThTpt
IoiQ/Ek3IuHokiUD7rxH+dHs67sMt6J3HeTv/9vVbo9TRZGNFQklT+uuEe9vV5VPLW0E3UmsbneX
he57LJDzH5w8gMEtDxu3PBfFiHlbQKaN61itmsjs/aD1AMjgJ7b7sK6ltgi90iEKtI+VMQkUnBBk
7bH025g=
`pragma protect end_protected
