/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
s/EpkaZ5Esr7MVCzZEwOnIbHE00zL1gAu7GyDpn5ZES5Rq5iT1997rhg3P+2y3RuQKGkS+hbEgHQ
AbFLDTarYDqtmVlQq21+Q5xHrJp/tPypJ1CIEuDdv0JZvU9OvDqVo427vSSf7i9dwUBEXHMQCUUO
FRqkUjJN932YQ+jGze4li3CyKb3ZAvxjVXKYRRxmKpawa1ctnccaL+cLJMVEnhal0WGVloNWbkea
Al2W/r8ImaNwMN2pB3LOmUJS4nR1j+sIdGQZsc7p9CmzmOYhUdJK7ZVr9L0rmIlEWEMEiufh5U2n
hPNkLyeb+2rUlLHd2em65xC6njRVqOEUU1mu+Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="tBdlzVdTlQudNhqUNZo99dMs8f4bAb8hL10OvFfzUAk="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 303856)
`pragma protect data_block
k+eUtgvNJkI6TbcYnLUxbHD4B0k2IM5rwtjSyw1EFkrIC1yuT9QGatQOzVcnS9hqwbWDsgACdoph
piZc33KFai5blSQBdlNgBmEhOERL0F1uvjei/aGrG/HxOoo94qn6rIJxJwtcyhcQoZqLFnVFQmLJ
MsYGnncSEq9XLxPha5qsAN1WG9bXq4nX+4Lo/KoJRxO9mhqtdUJ8mxcPpJ3Niggg1R3AH3BBKYr0
7pPTpvquOtIls3WT58y/VhSGS4ZAmOFq484sgnEK3ShO91PaEifX4VQAMQRIq+8PdoY8YbW47Vo8
BZ/jNjuXZGaag5QU56BlUypaB3QQZ8cIveQeDcHUcqJDwOGtpj0IEiVqYKag3+W87UIOI7/vczUJ
F4wg06/pGa9vJ0INyE+iCr4n+qxucrK6ZW+OWtMVYgCyUghQbqZWkkvi833QNv+moj9oWc1MyXJh
SnePSe1eftkXZrgdt9hFhW0mz65GvPuaFbFd5aWWwrE1Eel5icxHGgfMPrwtTdeQjgJmsGPD8AB3
qEXNIGSDfWB4YOGcGM6ij9+aa7C5A4GyqrAJrxWYl1AiRswCy+mwlonQ5BROQ3hbM3aIXKy27tgN
v+5qj7Q853roBnUaymjeLEk9a7uoP9y9cYJPv7C2MF+sHO29Dn0rOYR0VbxZifdGk0OVp+TUi6hh
c0edc4lc/lAApXRQ9nyZIPtE9bZAJhQ1MwNTEjklyEVwEn7CYdlMpbP5jI97yCD9Au2OmqWkpyTq
wAX96achNEcmoddQkdgPJTN5ZM8JSL/hIRJxtyyc2JVqGTKM4xBaclDwMtpR2lZlMdBZ+Lp0Eg6K
0jXDRcXLQ44w2UV3tUwHgBVGhag+Apf24et+1EUhRqEeoBPx6XNFhg5FJskP2r8L22MEnu/kINru
OzMN2yCBAbUW3KF3Oab7d60psX15C8fjA3rLGYctsIfjDwUqB3ANuU7e90X9tF1+6DqawPHdI3I5
XLmwJ7G+bJ99D65Ct5nMSHmlW/90QWLpMccjPUSEYbBUXgqcayYwan06YShPtBGcjasiT2ZuzGS/
LZv2JV8tN18Zc9tUUFcm0pGxjpHVyR77eBK5lyh8Q+6dhJmYSV30TOExDBXP3E/+0TbIIReBqMj4
a4e5MOzEOFNzN8W/x5NYFEVUoq7sE5iT7k8xGpaaZ9abjUR5YoolvPJCLSGmXyze6X+IyktwJXt/
CsXfD8RSo+PxYUC2T2iNBWcxEN7jrBV4Vfdh+8s0AyWBGOv5VvNRXpXNh+GGttm3sHZp6g9a/Dds
SsxLuvezXE0y8zzj/PXizyZjAwiwhvNzzE7WX7g5fpVXlvOiifw1S9IDep2rAY84OifinUb3LGrs
TBDUO8yl8FijpK13W0y7pHImLXjdP/l9cKgYXVDUKPE344WIAneBJdVp0kw1VM6W8Aw08D6+ac8k
VxS2i4aTGhvVVRobhSqCjMfKwT4ry9TH9cWZRMArUMiC+CDtDwKvt4Sn2ieHjYxcCjZQpC7S+peL
y5sYcgSVxuZFh6DP4ALltdFA0CP07LztjjMukT8iZHpyeEsZjWOSi43qOBdR75T9P2WDCOdELSbj
tBwke4TiVzXSRHKu/aoia7EX2IUhVGBEbtuUinbcDis/+QvUifh7OH1YiaoNr3IdYrROkX4hjZIL
IMQFhhSUCjtpswL2VtIuDLWzx61GoQabctuLs0zbALdsx7IrGbh69CK0WzHIZCjGg4enntQ8Ayq2
az4ffBkSBjHxx9Jd5JO94p7GwL1AZjAq7pLmoKWuWK5rVd+66pimpWi5YjYKwTU7m2GmPTvxZora
20/chwIuD0K//G4KPxgMy7uPw7ffVwe2CccjFEV4+WYeLk42HM4kZfnnzxbSpmHpfKMdWe2IKpp+
PH/ZZrGJg9wnnGBgXSG4ZvFv4RwfoZrNBQBko7xFuL0m/4lOolySFjzAOTo6SxPl/Ng4HEK6VErk
4I31ZFeFI+k4uqVZ1wXQpaSrnW9XEqI3BFDXGM2/I7mM9YY+ADvNG0sofa9n/n7KSbekZnrVSsRK
Q3pQz94vksGR3XUZK2zq6PtwTSQYeI3VPxPjZZk4WYqMM9tpW4V6Wm1I/qic/hJIbORr70yBfcwu
k1oUzTQ20d6+NMNiqhon8mRMIuR/2Nfouamyc2ZDqEtWEvlBzg9pcf6RwfzjeU2UNX5Bqeq5xXlm
xt/UyqaOKvbiX0b7i6WK0ME357ErOJ6Tpfusi3YRVvv+hsuci60+k2A5kWhu2f29H1x5ung57qC3
gLJht4KLOC3L7iJoywbzE5WvrTgJXTZVdZ5DmI0WP8iVT0ESfd+rrZiBahgYHlUhKAOskwBuchv4
qXHRctO1WRd2+L5IgyxlO4JCcFTjpIa3/5ag3B0CbwJKEu99jeWsFeBHeu/sxmUcmuEZ+kFPDzET
h76QRtz1na5mZhyFWu4EXwbKYRukCs/OSZgkvAoXCl+znns8MOWBwmz8W9Bn2exwxx9hBS1HZGvr
/AF06TdyBmDZ/fFVYz6WO8BzPtBZi9yK0YPuE13mXg9oNwxSmYSXXvQfXHTxKiQYnZfj/iJzyqoh
zPurNS90R6mw3uG9C0wowQmdb9CJrnVBSzLOm7W5QwfYepZ/7tnBLtEyX1HwjBIRRQ13keqqvsVy
I6mBN5kw5/JbTc0Ct6Ebt9ycnDmD6VbAkP087NVKBVVYXl5YaQMpkHAY/KFHEvNcIxxnmrJ/HsB/
yjK5pO+H7Wgn6ztQaN44eVKnRjPWFSzb/ylcU+TkWlGnCPZC7A+czgR2VTNr/wGEU9aGibuSduVU
u0H9pquJosgfRMPI4Yd+KlmVhRclQOYZQ8lEvgRWH8uizcG6H1DCck37a0mLfZX5q6vtHz7uVCWE
z7VJhDP0DuPytnRxXu20TCOrCnD13sUougPQu9gwisLn5ZBnfIXC+Ln1ENnSF+dqYIudg1UwANAS
qGf48BlIEsGjNZGCu88N88ln8Puwi90PrEF6cPaCMDMKXIBYDyLsVRvKFF4dunnWcbOY62idMsSL
0CRbrGestoQCHfOKDztdjr5UCcbyfz7+QOLrv9ZjEBljoTkRK00vk7c45qgyhU3oWwgsvmmSDT7C
vE+45TjQ/S8rIAw7TCyoAKAn3UJ8/jQcW+TMH68j7vxsCnRts8ZOTQXSmn/nlQ7y0sSxb47GWHpX
dQaB8P25rVUeC9lZr9rBKMYNxM5q4g5RxTeU1oLH/lkaF9HELmi4CaijWWoWF8y+Gv04NpVPtsLV
TD75XIJntCyvprGWjaTWjAe4KX2EB5hblknFZFaR74gzd2zYZDGhVqY2uU+VuvzjlyzYcph8n1St
B/newBlCruE1uVTYppXmpglpepcsCrsNA1P9nwuboSNUz2qlyLvBFybSfHqmoycw5KyB1KRfSIcn
e7yiz2t8lR4ith/YnU4aT/GnqkozYNYSgpApDV51wIHYpnNAbfXaeajAx+b22hf1TrmNhTjFXpBL
+b//Cs1ta+cAoVFpLgOLgNNS/29MbLaVXQ64vybk4Wk6t5SZG9Re0bLUjMH0h1PPl4p8nqRnjIj9
1lBnhA3x3TdwwU5rsqJ54OfVJjEhPsco2CAYulw6J1steP9vSopJfwfLdj2+YalhEg+W82SQqCab
bER9GbjvJqhguhHR3BrRAHChIdDDmTELesAJV8AqNPGvC1axq//PpOFuNfumOtyE4iDwOuXyDyu6
hW0G2UZFmc3JwiT09E6iOkoMv16ulXMkGH90n2mc5IrAlLEkeuMS/tAvu7lqxK9Rj1wqTffleZFx
Xk8TF7+DQZ4QhychKGTuh4D8kIwjHJwxQ1IJyPRZvUBbcM/qMaHFzo4S4U5IyTsvUb2+W3kcBkXG
XHe7EqOlCZ4sLETxezN5swFhV1A4Z6VBC51sG5zigNnex6UVXicuYMLBxQOykEfQfyHzXWkYyHNQ
NDcOin2VNUHpuV/qnU6A/0FwEyNaGP4qJnGfDFyDGlanoUpzwGs3SxYDJGLbHS7MKbrVYWGmVmwo
90m+kaoXgoVgEJM6ICCcMHheTQTIW4aGNKq34/sknm91JK0yA1aXS+fHo1GtR4Pr2g9anoqYLdOr
TrSYXBCiULLQYEiYQNP6PxkeYOv7znNXRbqvl3mx6MAFxikQNJixhFjtB6xG/SsK2IhZw8lgvE+m
jTzYAID45xmae0nGRiMVJK75FwIkNSi6yIc4BOdebu8xLTHEXgP75ooSHYiE7gitHtoGInNLCwHW
mpnxYcQGRYeCE7HK8nUajvNE0twpaqd1XMU9Lq5MuKsTNh35yRTZkPLznVENpT+xM1/aXNqoXeMt
g3oPNvLHo4k63m2RguZEA1gF7JIRvpDa9Yo8JHn+wviLAiROoIsZbc/E0W2V0VKKQuX2MlSwcGNa
1Y6i6WWx3poaJEBHK93oY7fB29Qbx/jDCLEQpvmaLjm+p5MkgI7VicbjlaLGp3qlUAOy/0pxFj5g
Mct7Ax60bb2OQgUvLGr8PZsD7xl3ETqPbfSRrW2vyfrxi2OXsJZ8B0s95suYyJvvq9nnAxTuwcYq
MV8UHdLVHAfwVKo4C8k6NY3RJCnkMJPX4GaHKEEOnIPXFdDZZoehPRbW0PjNp8xZceNicvtIAb+6
KhJ0I6tamKKzloDCOxLlGqOgGuYpdszcvSBxWyAIaEaPNN713hcvglYa5IjWhoodX2iyMWDWLmjN
9cC8YxPeRcBYZ6GXDtDgj1EqhVmmoY1zfkqTqaWI917gTvrTLBOXPO4i0XDr8QW+OEtKhYqNsodZ
2ilal5pKtLDAmQZspW9bkl4rJHNtsnk++9UXwQ2C4pynUCX7Y+wSn2wKAmIXRY6rUKFx4iIv7fS6
h44bFJT0rbeKdxNvJEY/U5biypBWVcVw9kb0HDv0pvqrPWzGeq6YOceXCLgy2MfMp6uQzNl96CiT
s8pl/IVxauhS4TuyJjsUmrM/TO8AbM2gAKdCeuNygqGrtcU3RCu0oD8RMgCVKKV63ksFdqzuehxN
fuCScH5DENcKiz38swv5RY7d20j2YQ5xXpujvM/3VDnC+530wVRt3uuI/dgWyxrcU0lCJUbtch+K
8YK/FvOhe6kshy/ROTsKjSx1yzQj/0OlSlXH6ssj02rlV7DKa77vg40Vrh0Vb76CVjAf2wzeq0FJ
H0cRZLOiXHZU/AVNY75Hv1G6MWdMvuzIZ0QtnPF9gr0E3NCmfG4LslBdu1h1v/nzenpkMZILCdEh
mJcpn8nVmWAnOz0Q1rtg51WubvvMsHiSP+VRhKuUYzWvam47Ye76zA1eFsnqR3DZ7sdxUbnywbzt
9VsTvcxryHVbRVKDRBXONbSzOE7ZxG36O5Xolt/DyefFx/oG52isHGngD94Z96YPor50bKRAvUMS
iKF0uC/1uc7RQvcTzW2aXCcy3U1mtlD5B6In1PEdm05juNlph1Cx3MTDXZfMhxvn1sZ8pDwxg6kb
cboS96dQMwLqkr35/nktwKnPyOAkG/oSHScbKmFvQZLcAu8nk/X5AgADr21MdDxxXZNYSOVZCZps
NCo+L9vKfNVCT3RawBpCtTUuzqNXd831dmGedVtALegm1ccRXhPoOuXeEQYQRy5B/UBsSlwJXEpo
sqJYLBQd3okTQlBXw/pHkf6T9R5VZ2JG3rFrPsSwuirZ2u6uNaXYsXJ+nqhhGlNYmtXm1vNWZmQO
AR9ikshf2Aj/wCHo2OnOv9k+ktRKlJt/QkeHG2HeG2jM1gEyOV/87c9T8Cb0ya6IVQydwXH8chZU
P0KOwb98b77p5EfIGCBmauu/BRToFEquKpoCfKoNvdjJhjmi4zEx+I7oIIuFiNNrBKUGg/X26iFW
Va8ieCl4WBWe0NfmStf7GRYOFnbx+VVswC3yFTg/ZznavSjW1RCWLwtXRHiYV8WsuXFI2K0dcp/X
MXL3UOdrtHPyiomrWJSUmXhlnhu0T7tzHWd8pNGKpTegnJwczHHA9QzE3wFO7Koq1m2FChTjENbj
XBY70xs/9INGQ96WBIAi/5GHsYyTOASjZXwH7LGorCR+y8DDMO4n33gP2iQ4lAh2/ldnvXQiquRz
ETcYa8bOzH+LGSwexi2KCjXvdlSmrAypgxWW8Nyb3vNSJPdPMSUmR06GmY0/Vf15y2X3V0BbxdpZ
PoACGepg5E25+EpCq5hSKa1LY8HpiF3YHyISsWisSo7nfWPshQztSsvqu4C248EWd7QZZEcyQCjL
fM6kCyNvwC/rVDpc0fazjJz+zEBmmRoPQG1KsJSOOgG5MmoPTR3xiRY/2+h1U4UpGnqvdFX/nPMs
+Dk9aiMj2hQq/6XE0UkRIJQMvEcCXEircPT2BnQcAbLsmvFwOn8dLoqef6c6RcpJUKtTvqhoxOoH
9gEK8RShlZ+A7L7I0exbe4RUV3UmvTHWIwyr43Q6SmN/10n0or0zkxKqPnme3sWPe86+EHjZ8JC5
n0gXkRqXGbzqw9y7oDVn7CYtmcawPvAfzxhODRhvQlRi8h3nSXUBuqVg7mU39e3Cd1/ojMPGs2Vb
G+m8+30iYqYMj0OKwNOeL4WFLeS8+U820Pwy4cEc6P25TDWVsrtdsmuBJEaiR9QIQRHGXYmZbbSk
sMIQ00kFWPRYJ7qN7JZNYgb16IGUcLp2nZx3s/uc3pJ+c4xki/k6rlkyCD3npc6Ju37Zh8QFpBx+
24gfeQqoMLQ4rQ9yQcmzs08wrNfbjlO+vYI1CVHJ62oCNkunDK2uimiPd9WJibyJScHIUUx2Yixk
wAR27ZaUhWUuH/gJWli6gC7APSwMkCx9CKdPxmRqQSk905Us0KUFLitmV4dtL1ZHVIzt4yjUcWVZ
zTvhqshvh98faTEOZnoPXvq5aresYqpq+hJki4iicJuVtTY8AbwFV3Znan9zuPjJ9JBXur6TyUjf
b++XenzW2g6y8wN4O6KzU4RsN5gBcIkwv1cgEOMbRetNu+m9cqPnCptKHfYKLwmxIZvXnKaV5RcB
pPamnqZtI7aKkfEpYtL2J2xhe8HO8YTdAwLLXyx0EvMwR3No0FLHlJTGpgWfPABG+zDFSMiLS24n
c7568xw1FY13Us0SW+sR3K0oCt3lOV536ahx4mM9q17diTnOrDy+/dY+Q4IHrF22ZFj6d0SRRGf+
07MWDIWxEKdvRktK8DWXh5R9bwIxALqCCN3pM7mDlJcCrMlZmoUYcJ+42qoL3z4n8XSzi2iByG59
6nJ0ARkdsXa00YOQ+n0lTTZFTsKlNXW3qw7VgOXqIVnypksxVNr6L75gqSlXoDU9R9YAfSfOvpEO
N2VyRzDvCriCLYUDBwLL3SF7ztUKeWr2ANc8pt0/6ADWPkQSicn5iWJGrbb4v3sOHSoM3HXrtbnX
7ar8v6VQUcZYFVKvrGRw1ah8siKk4FPAPACCNLJ3WkjPwY/xYujQC5MoOO9mqUneQ7PuMm6OK7Nm
8+f+AfYFTBulDdfODwuUsjkQmYE7kAZhP2a3+Dc3J9hNP5hv/rVIXKAY13BKUb65xAgk5uQrz7vW
LoR/rycku2ZfYL8xF4+uUmZ3cjMfzAkmpxZdl2BryZ4pmHSb5i7tsvqzU1b5FjI1ymShnqzzV5dr
z58QbMbNcYxnJKOWbbNi9ATz3UWp+Kd39GhxAIp8r7rUGkimVH1V1QLXYSXod9IwNMVa2DQ/NBDN
Oy6X0TX+bmRIrzrl1j7wEzsBmy4xv+MDKmRdKHBWfkMUoIymSc69eZDIYN8r7siKCMs4qT3ECIR1
1wMUmuCpnpTnpPd7+lUWUr6gZuqaj2GmUhleJyVcBsK+I/4b5ClYZaHx3NDKn1a500xAczIYPl6H
zOgHmCm73FDI0mjpVw0Nw7ZSFomeSl/oUGcJbfRzu853SKahuT6HrPGeppS2n2276zYQrt39wF/y
OF8BXrKSW9z038M2XqvuTI0N7xUpqHB0RoVrjKf5niKIkB0TLzkOukjSA+s73NovlM5jCxL9sZ/2
F2uEJIj56xeCMfYNCfQXQqteikNOnHWMNqYe9alYk/vDH4lzNhgsMQc3Bhqh6cOtMcnKwNlCL+k1
8T/wTf4ykP/6F1i3M4F+0YrNrJ2WqqzJN8k1Y+zQ3kWu6L04DC1aM/KuQWouZ4NI+5nsznRUTNL1
k8lCy05X7IhCCU0GuhSvdC4xwu8vQ25fXLcMity0Y9YEmcS/XfBMPcrfunjwl0E4uTvIByJHsJKs
MF/1fXSQC85iT5fCzE+gpxr+SdhGSn8ExltoWkWGvqwR5AYE3S5X+TxRYUsmvaQE9+ciHiuk0/yI
BuHI2cDZqsD+8Y8nXDBoyVwZ4ZMRNDZHRGHgQASejdT2RvZYMeVyUwjVv75un2AORKcu4M2+TBB3
XquBHyEnD3H+7nesq9OtwYKBiasX9mrwDisBtnwcHJBu3cDVATJF0l9mhHj/rgRwKmc8YmJPTQpU
s3WTKCiN1zzqzKP/pcEtp2Hmg92UjUiLvfND0aHzi/BnWz2QeA4r9UP+z0zb0l5OIo4cjLD/7Y81
kwIIPzDMbs5DIm7wTENRwvkGucDAegROdwm/Gw/XNDWZ5Es72QnIe5cRobapcVMev75/+EI+lYkU
8to7Dzd4niII3NbRoQ6YMJ9l1rq3/S4H+jAp5qiyKR8pA3MxOFAn18GwRZ/zLSWmMiVLqhRTvE6q
xigiun4hJ5ukwuOFAKSk8IvvKcYa6XwBmwp3KGewYNoV7BYb1DDor3QWMM0Qj5Fv0V86Na+KYQJQ
g5YBl+rJdbFBxwLQewqRNOZEq7Qr94hUZerY9888Ipai3B2mt788khltVMenv1zwMFaOGg+nOkzQ
WHTF1CVNQipbNGr6JWnyNYHVgsZh592The0fbQTLrXyK6NYgh3DQt61gha5J67/WSFTSV/PvL6xV
Q94s9Jf5wHKqMVOVP4V2adCjWBYm+dEpohnXWyPlfRWrpktKigfZbaFk6aHIQw0HQCgg10/dGAgp
8YMxvLTlIcq7/ls1lOMtOHM23JFVasYrx5C9knz1svxLIXok6Zvqfql21SNjM7NfRvw434+++mWq
1FhuYVjllSdfzURnfTWlGzWzdhQPEAZ7hGJ3R1ln+E+bkDwy98AuqnBpcV4ITsOh2qDHwdedqscg
Bvhkyo9IriBthpCv6JraurXDn1j0jhBNEfmNTBQwWE5ehF3kr4RpvrrkFHuXR+82efqsTCzTuA+Q
FSO3ukOanE3gOI8EjMNW84D98EIM3xRH5b4EPWVel9mEbyt26zMMH1TV0ji0jZ1/uQCIAB+B9Nyb
Pf4kJvKL5bRpFvaHJX0cbTE8atVN1XFR6jzwQfCoOnV9NZ0uJPQzIEkmPHxewnk4uSriztPlKz8A
qQn27NkiflFGo2A4RSguUDRbLzxfsoveNmmCuynpA2irHkSVizYkZa/1Z5Nb3Wg92y9NobonbEcw
XLxXMUnk/7kdHwXKHGb71Q5bQ2i2q8t4Pny4ymzcVX2+9wSnFSBtFaAl/HrYuD50OqBehGM5IUlo
jqFDqCFx0dmiRg8dgje9tCDl97c9Uh0dJPzu8VTDAC/FcJHzKY+pXTipDK2xhjuvGSJr0sZ4/b1o
KOw0n4BRxvd2X0g+2N2FOSMWRt9PCa28j2eCNYRpjUzNYmwVQOlHrNeLG3JhKzsMnOm+QjFZh2mf
v11UFPjckAqL1Xd3sqnIR3KGFnllGbywhhvBHzYjw6Wz3jHJ/ky9qQdTSBUni2GR919Iojwrzdzz
a3aHQ/L+N9oKmd84Xdjo+WjhHe6vNVYPTsSb7XZE3fDj12FUVFeB75W8YQd9bMNiDREm6OfwdZrm
sRrlEVTwsJv0iKhhxY9p4ifzya3scO8LNs4RGpkwz8OGdA4z/bZJHuycNIrKdnt9sla1Tf/WI9ty
pg3aiBX0kR+lzsFk5gWZMNF7HbpXzRImPm0F8gi2hubgYJvPBFTSyYOocFg87xFs3JuVdXsTr+2N
BX3QVGt+swNIEnqYfDCCn4LSoLL83QqWArqnasaSMByItfu+0Z/2fBcYJQ9M+s2UA5cbYmbeyhCS
lqGpWl/56A+LoECSB56FHet0FmMWmQJJ7JYDZH+2hBVN7YBS706A1ctAVeDd52rN3mIJQ5I8PG0v
qYFz1QVVFsgVOxYFCA/swaIPewOM9GosTnENmC2XnCGpRuuvo69SelAcIDpAWNeZxYQsg0FvsNiK
lIJceLRpaK8ZZVpK4kUy2gI1/1JaTowfp7vDNNXBzOX1vBDdIXwPwaUidhLZRvL9ULWa4L/dljcX
bSqsqqLnvi+1Ukn5igld3njdf8Z8WXB8UH5ilQOOGcY967becGvwSbwfkWw7afKAkzv/kYWhGIM/
51pi58P6ArC0Z0XUaTzh9qW+howL9rwEppAmzyBe8MLR4miGwkRsGEu87g1ZW8KF7DSyk+BTpb2b
SQdXkes8K8nV5UrQMbUH2wBit339pOd3zrO/GBsxVxR3lYou52P+rJGq2+IHXNlNttyzv33G8t2X
cNGQ5TmVZdwimDhIYZMCi5YWM072g0meNeN1206u66N5B++jyWpFSStJ/qQBSChy4FgcDa+zBp7N
lPQF6xBJA/6lrQ6rDJXMPzKuYDAmstlv379ZjFgf23mdez1CY4EHY5LMwybha/T8cJdyPxNNRWst
HfgYvOe3I8JfcW2SQqtSFDneImMWzpY48/je6vYcmFF7YPRNr4SLLGtAIUbkw4kbgb03pkAE9UA/
yYfzbNYk56NkzYqUaBj4iEsVD2nqEQ9dObRmoSCy3abarFEAOclASdZ0X07/V8c289kcme2xZJrF
HzjlbHQxcNuOmwktc8g5P98E4W/SPwB7hbijpVUzfVBPSXQpNN3TgyDySPNSHxkg+GV2VtEgVrVD
k4lpGaJNiyIcmrXe9UcAAcoM5ub1MehwOOb0Bt+4f9/hYMJ7dzMsmcfnPWw6LGMzvn4LqjmuVzFw
/xZJSeuPBsOXkavUxPNc7aBGcEQkQUuL/UeEcGkYd+JYy4Ew5akd8SjHelvUIjA0rGQcRVgUsmU4
+JQHC4DOVVfJACDSoWsBjuHaq+vdnKl6VfrmsKcV4LOsY1iTzP2moFxVkFMk/OKZr/N3Bw3itQ6S
rB3q3mV1QXa0cocpNBQoOcSVGg3muYbUm0/pqPNfOxk6HGLS2kz3oWu7xUCF8vvjXyiuwfynIXuO
K6wqZC+wnrdE6fiIqAnvbzIyZ3L6B1R0XYpHSNJ7RGhulqoNmMF5IIzB6SzgPkPcdkUoWpFqRbHh
Kre5y3s+RLGOC2jht3pi3FIJC0vlP5k8nm6DXAYuM3LQHOZbI/TjnJhnZpY9+uUCy/BXp+P5jBuV
qIDiqLlxko68If+dwgvxbqhyH9GvP0wvtygxElCYnFaG/PYeLjelEpRq+QLI2NfF3KaqSwk56DTU
d3Hp3sftLweICFyQeivvcCgw61+ZUAuXjo/CPo38v1bNcFbuu/8lwXg7qG+126u0SjADDKRgXRxX
OaMsoaewB3tMdwwO1rOhG8cYH860jBI/PvnTBWvchXzPDlHb57iLX89inpt/C2o4pvrKFeWJEnqA
Wl1HJyGKDAt6WKYhfThcUsYgbHSJQMj5W343eUKF86hvrDNbAWb6JExP5GPbwPLPFmx0P04Eft5C
Ct+gzUcNsWu2Mlh653yOiWWUPX4n5S3foTxCk+94dIJu2QBTkvQDrdRgiSop8FsL5um/8+2QmhIH
9BUZxL79DC8TEw3Aeyfji3PPyj0iI8derIRL8V75HmQ7ueGX2ao/LB7rzA5lhBfoNCfE9iz6rOvg
X7W5odDQ1+3Stj6jrJfS3ybr20cTwmOG5NSHmax/hefb5eb7LlMriTjG9uxYiYkUcEn2h0xFLcvX
JXQwFCPORFztMfYf9X32OAP/RuRXkCFUi13v0PFX2ZXivNmi6W96/5UnLQTt6S1R1MrGQZmC4lWo
oa4GOlv+A6NXkYTWTmZwuMyd9HmfwKijR1jpiyQFCmnqw0Pz/YoLa06Y63Sc9i270npe3vS5zR59
34NObq1PhQExRDv2XAyakwb7aMn83HwKabp8Y3oDMDoSe2mum3tzYLPvN8Xbwpyias3OsmlfU/sl
uCvePQOVHFzViM3PUoyHPyQWZqeI7gUONW0S4eTRpj5Q5NbwEu3qRBvJvpn0Z+V7yqYOosX+MLNt
a9w2BuXjHfUu+RH08VOehvB56x6yBi33t0skWfx1qnAoqVMKqa5zA/RGM3SFhs2uDURckM6h8xLz
PvWgB8dNZl4YQGnrIB8cxQFDLSTn/+rS2xdZWiGTKb/f3WeoWBZfFxh48C/jKXDaxLLP83AO1RsO
Gak/E0yEgfIJCpWN4QViW+sOfP9fZiWlLDGNSrXjYHSB8/m7rZUCYhzd2waewlbdJGINzHt2KoAk
2ZSJ9wIryZZMDKvq62JHoyOlwbueAohkeLuW08V3JpIPMtTpP52JEeK1rxaa8BN5D/V/M185pjcn
qEa8kLrANeSiOO2g0Q7mQyWYOUfbpNC1hXA+WFEP2zutmSkt+9zNoF5GvAUh7IoSim9CTgibUPxx
bgXAi+u2zHw65Q1+6uFb50mFCW9UQiOlPzaDShGbDKVMtAJa48CMedVFR9Legj0IDyjYK2Dltbsb
uJN0BuJt03qT9nVLHLlkcLlP2PK/N/7e418FuRWuv/gB8RbX+owLVlkRIQs6ATYzTnyaAbB1ncsT
Xt6mqFHXkJIGph+Oz1VaqJ1KXyGwtWlKRxTb1YejaI3sAcS6AWJ29/HFUSZlmMmHmu+k95LO1OnD
JTRpShapPB4+UYtPPBz5toIQTx7Bfuo1kuQSqxncaEOzml2Iu5yXRFM3QkYsfrZs0yc/zhLp0r6w
39SfRB6lqAxo4hyvJ5fNBlbCLg9yojqlvWDtwAQe+IGr2i6qiWI5Z07U0P0U7lk40BqxuH+PqfSi
7/30iRWu4LxfMIEDLbAYdhww0HO7R5aL5tDMZDewkLQXLVFkJNKm0B3DDyHMfRyIgK4zPFpQevxh
V0bE6ud8nEH6VGH47Vev3QqGwX4vruvj1nHeVXhePKCHwVZ0iZiYJiYWwl5KLSWkCsre+euxVcrH
BHrgfuS7iTpLaP/YZ5ttiVfdjhdd5dS1zvjEkyOudqBhkK0GnzfoCrP7TRSdojGo2uSqRbNOcrDu
jMkaJMqnC63UgZ4lJ069U8ZA+nuB0OFxW4XELC2/fJpMCp/hH+PFMvmipgEWrAcSJJ4DaWVEFHoB
ELAjfEG0eXdgEzdNwzzM8MgX9Na8pJFAtB8v3z15Ojy2E5dlF6CYPoz9D2jkeYG4XJSfL5RlqvE9
9QjuqKnYptTn301oFFOquVk1BN+QJ8YmIa607DS7w4/5mxtRXRyb0R/zsOFxfAdgPax/snVLvqyZ
FXzRjmP1yM20HG+F5mfOE+9P/OyTe6EFweIM2RLfqTk8k39fDmUbepJtpi81Hd+IT+IvN9Hk+6xm
bGBPW+ltmsuqhnjjXnfBjGmWZ6ojcEjcGHMYwjxBMBh+DQvaDiP2sAElgVmo0eQD+nv9iUe5IbLk
10PeprY1LWzJx02o7kXsynRP7+Mf+odEtILnschvaHj8Q2qvBzLELZK09TI7fdJArJY3liVuSgw+
WYEXy9bRBgva4GwcODRVwq01sQXiZ3ehrnVXZneq+HcC+mjcmiNKDkdkSSi2Yg9ihFBGxRZjsDOx
d5kModLSqxSreenN4qpAZZ/dgAHU8DgOJE6wTPgA5DSz7CwJxCXkWbdigvuXPoj1elgTkNFrtV9C
NEI2rkWnwfays4iVv1dfTR7wFUsXY/AWwFcnHUn90P6a4CLQ2L/M4LwV7sneVzK3BTmYkD+0xNHV
INtNRKgUMPmynXudGqovaXqJCyMS9W+oozeeM+3dZ6JQd8r8mFIeKaDm56OR8XB4wrShtGkUVXu/
HISywT/fSFe8GJtVAHvqKdvbTyyaEj9Rh9pmVqJtc23M5vGo4g8wMJurQSDfEWj+D1DR7mXXE2XG
8gORbcbSyPpMKkdZaRd3S/3ytUIEmuG9DZ6jP62hd0rwPiLB7HmFxypv4ARCMuyFR9bZ2s9VlnKQ
bWFOpR51C+/8ShRwj+bd32SUYoyt6ciqytHBFYRrABmOcwBD6px7JHhBP+zlgGrDjlO+wryMBaqK
WsmXWFRzWejAwwkKpGdqFjjWFZzysHgzgY7d+dWD2VXTSpQDVg5L2Izjgfo1v/62WyqeExQI4AQ5
HZ+Wye7MJd71UX80xyyYdY8Th3s1ncgEzt1VJNRFZn1rqDKBaaeHUj0y+zKBdkVfytR21DAoQaPU
wwXMjIo1+r2GWx8RyS9p42mdUAKtULqi6dDWNlBnmZY+IYBC4kf22vpbY16P+/ds8NU3swdfdRB9
RlrwXaYHvRKkQyDmJim5c+Wzf3rmCOlsLi2ju5+AE+0VxfK2ycdsNrBed234D6mEFcAVKre7c7WM
pwq9DRTHUQP/E9WpxqCQ+ulU/OF2ipF2mSCWgsU7AgplFpacKKNx+ITccjwdemoFJ/RVoqr0C1xe
vfEiIRqBHCYDIEYIIf67FkjRKJSqx0XCW2RP7S8x35Vdw7Mz3pUCFS97MQdubVLBNLiKedxRK9xF
60buvhtZhH30gHeU97mWukKTdNLlun1kX4T+ugqwF//scZ6Dq2q7XOuLF/nuGrNStcQJff+asn+0
9rTaqrS0g9kBGqMp71zNO9rk8EBNdcA24bNaAKggv2yQy5sgRNXlAHqaS2AHr++HtkkNMm4s1Odv
38xnypDOHZxsEgENQ0ZEENntn2b7skXBQBTc8aTI5DkcPKrhKtJtzMZZIWz1Z8+qu0QoYEVfRjL6
b112Rvt/okZ1hlFenpPMl+JmU6SV874jGB2fBHZCPtNCtApGTEnhiIeK+M+z0H/HUMHDPq4ibOqC
zDfUdg4b9JJy3Rxq4wOsmJDo5xW8ictceUxftuBkVilL9bsy1quff3O2thwZLp8nEgnxLJhfm/hY
GRS9HX+qsHgpYCvTLgcpPUauVDVeKFttcS2ZuW3xts9KXCY6v+G706eQOym4U5oVxLyNjoEiDW6s
av4O0LAcdPZ3/qXQXaxwsDa8UIT3ckSmZJ2YDrjiBFcAiLeHgxs7+E1Yrp8wBvcmd+QKQkQxOthe
zPoCvBt0DW+wM5oeNpdbmx9A4UUd23qX1Yk3sGma2h7iGP2qvDFrs3bOU+YwnjbyoKmhyH7Aus57
BQ0xHLUd4yITawDD1P62Od67GghYFA/ezfmhFxAIjhvREOAFmFxaQ0BDVLLXxUFFaBEv5QGmmNjP
nVGJEQEG/qEDYIFpp8fnqzzbdDaBsFOaZ+rFulIhd+mxWWHhH20ZrcaVcvCXNgEXrHRX3DrlgEc1
wEQiSa2J7I6QxdUFRAolEAleT1lpiVJHfQIL9xkteH3aPMLIWBwUwNIHL2o91YoLM73Mi113nO9b
qI5IxDNFGnTRQPDJxRjgaffzMDlWVJBnPeJ01yqokR6M3qrvDgVSSz6ooJQiHPDGMSgGDDU5UUBT
SV6nXTjogKVbRKzJ81GZ5ge30DBEIMUafnHOQBL4IRVYVxjYu0I5aatz8wTfN2cS457DtA74Kh+S
YbnvUw5sxFbLXQXltSQviyY1yQ1VacZlnlw4CllbwJecLZ4sFqdsRKFyCNcYmjaDygsEMv35kCrP
siJnGwRBV3JNw5cB/TDHRUPTlxgkjtS9qib7AULlRonMRCUy9fEx1QQ6K8ThbW7uTEyVgxsCI/Ic
QbEjBHoe+AmON4ktizbZEeVvsonrkFNSZPrfP0PnhQGgg72yk0fvPKILnkLsIu4C7Ut3aikQTC9W
hJrM1pFH5me+I0XU9vOzQ+rFVwDrqxvNbdT8iBpQSqaBIxw0TWyyJkjDLlc/b+SGdWj9DCwT5ZaR
aKmHhbd6BDiISRS8fFI1ODgcEgZwqM1NyapvJ6dobLmZPFHpRGouzdH2sZdsG5subU9SSRjHI64D
Oj+NPC+1jMXou4C+QRSeG15ikpuex47Ipwnok0y5xI+FrxEX2ultSTifu6PlID6sD4D0qz5ngVi/
Vi+fgCQs6UF5kQKzJJHElzdL7GkKBkQfmWV/ap1A8I/JtARrhn/KIbFUOgFoC61z3v3LQL4g4eUg
ijN1NBoSTMFPERDNEeZj8dFJ1P/1eAQmSobs0OCGsT+u53EUwkN+/GlPIp+HZzqFIKJ4dwtCr27Z
NPSIvbt7Fk/omZu7ZuKj0hZYrbc8nf6cHhueQsJAImmt35s5xye6RbuVN0WF9nR6Jh0lNGQWIoya
u3vH+amiM2oCap610n8wIGTmK7K5Tz4dezEuFmQUcrn82lPrbaf9cyxWdWhmxVnldljNPxurll3R
lpVUtawW1XiD1aG5rgGbkWL+d4I84AF7buL33YwVFxVV0WTRl3bEAmvlTJZEccdLYxAYqsJmceZ6
rPtxg9xHrNaC26CcvFxuAfsUtya4lSukOzNvSMbdgxQSIbXUUfkAuuz/3KKQDxYeWW2fSq9oVY5/
7TxyYZAkIhWnKZZ7SnpFdfwdY6Ou5hNsQ6Z/g05AX458P5af0BbTf4SniMemULjLKsoOTU2z00NM
Ka4aPwNtJQBLrdMF9mnx3OaA/eSo9tkvcQovOSzseVd59DTyigmz+cGiXQQ5i3b9Wi6LgjZ31FTT
oqnyur4C/cBv7GenQ4kmqHrQL00Q6jfUJNQC4YmmjpljUgtarO7XVduIBEeO+lF5/f7cdMWe82CM
qH11pohgSNy4IztNAOYAYlM7587C1fvABKxqdjyGhlALsg6MJ0YK2qLJPXvICQcoMcL+pAJJU0ws
KvrkebRRuMUe4C2nkdtPUb/b8jHz8jsxdmEDxUYlBLi/DFWrSyj9jGtR7N20uJ6+eUIJa8qtndDp
TI3OwhWob3hod+NS04BbDUqIV+n661ni2kfzAPzY8fMZXJXYy5g0gsP23LGB/8bHEEKav2oy0xta
+w+xRv0buJHmxqTZwrV0hvI2jmggzJLHmFH7NYLkte9dk/PyYnfZGfDpKW9LbCmMqJ+oWj1mQon8
948/TbwYUjSuXXMdMNCPIgcC6bixAC0RTvkmlcAGGgmjqYV+htGP0TzwjlVumb3Y9L3RoD27hxQ+
2MP2OlIIb3cPq/oAiM0LWEIsZS3bbcy97V/cfOrNhi3nxjVArOMQ4kaE74cbi2BVHmpgolyylZz+
IVwmIXkVwT7/RJ7SnOzfstloVKAhG5SkyncxN7cCOOvGduXzjMGs49REQzVI15SkMY+wRIfP2hQy
41ZvdORbY6t8qAnZ72HHqWCAlzbP7WWyTKBf5JeE9gIZA7JdFTnF/R+UE1dok1fUZnm9iBpCjgXw
ri5nV9T0A1SntRMh/TO48FzWL4X4H8OGATR8Q15fahTScEmOieHH1PYQJNY5+N27JtrY9GYWkoKf
jmPItkPqISmVPsmsCc90DN62xbz3ktbNXl591Q2+vapi3DUnRmg4RDthwsinw1tSnHHxYnpoGGda
oAzozndicIe7fUXDQLm8avnhPdYX/FwaIbOW4pxw834Aqe0gXBEa4O4BOCrhvYGZu4AMqPKAn2bt
Q25GMTJ0mvu2yGKMAAALE49+eYjSeOTp5UQUYQV3UyVYHDVUBH+bLPoWZKQxJigm7+bzbOB+nsvA
G3oLaz9NZ0qBd62/C6TL1n3jVndjBgWS2/ZUQescM+oE/LLunB4S7FHitAt5lKi/kkgONNGDFVDn
pklr+ZYbwEiQU81fda2KjlbmRCwEmtbX09AzSNEYF2fHQ9aq5x1MstltAIVk+ZlfE7acWue3QeIW
8FFeOOa6/KCRXDtU1UwM1lEcEo4ppd3770iblGRAfhiJxf7ICKEfTrpSrCcVMhRBmYI3C+b5ETcz
rkJnkYZq6qdmZkJUZKgop1IBXU2jOpp+ogunjZ54iU9AaL97NWJjv08nGh3VyGt4fVh0F2cmj05P
UdxWA3619uy1CqQlDYWFJe/tyPkyhxqJCss5/hrUZ2G+OQQIUTs1LarT2lSJzU4m/QJnYcZPkkN8
t1w0TjJdYPBeX01UwYBJh0aQF95oEJ8vI0GP8iNvEGfJKxBJDnEc8fW30YaAdmqKFExDdXL/Kprt
8jSRx7HOyxmqVfCIaNS+k2X/AFbhHJc1aw89IRXuWTzpt+9c4pcRIH25UK/iLhXNFtHkizT/avXU
K0aIWv/UIX6Br2JquATMKxNaW7OxrLF3u3J3XamPelac6t9h39A+noHPYqbi2xQRUtif4ofv9bK+
qybVDvUvijuJhTSbE+gYXnBTJ4sPcd5BohImnqw/3Q1qfvefiIPzspEyiiqG9UwRlSi4VAPNXzxd
vfkXUZLdnYxQWm2+qile9QQ8KlRKVaA+iPSqB2GXCbJsJeW5WOP1vvLLqROcx9No5GnR+zjV1xmr
SvJJtXi+Dr8WTdjlKPwnNZP1EPpSvG8HnbfG/xRJGKJuEeBy4Ozz9yg/cC68S+zO921PkVXTyBy8
YL6QB26a4VRZLPgtMYJN5Ygdw1Kot1rMhVRluCiGADnv8ku7cOvM7Sg30syNLPYBx/B73Oyn7Ihs
KAODVrDV+Xjlxb6UxHdZsXNb5JPdM8PHxq4zN/BdczW62daOidn/jfoATl1uHF5X01N9E4rLWJX+
3go8GgPNkBgMYdBF5BD2rOQLqYEnC1txKyeZ8ABbWf8YtuQi2SEAX0f0ZzDbECkdqR3pq9aUaYe3
ELeW9JHeHekxAsibAjYrYMtvD3NM5j9pEi8fzugT3jGKs3lLYg73JpdCCsnQ1y8rfLVQf7Uk5DK3
MRo1ac6TqFoOdaD10hWuzxmmkNYsFxLSDQdSTCnKFJuy+4fcmgGhXdiSUU1o32xol8CihPpJ3XW7
hoZbhMHY0GVnoo1lWHMLW2BEXloF+1Q6ag+gkZPYkjnz5EbRtqowqyEd/tkSKY8/ociAm6Gzw8TF
xDYlFXtb5IHLRF4phb0Tyox1sjPkGXwLLiAtQHljT3F4bLH60LaAfyJ98lo8X0mrD9SN51RkdRY1
9A9QZzi1cCebKutbZ+B7/UGv7n4fv0QmIkNs4F3JQok/IfDH+zh8aC2KZ8oG7YCRx0KIYFAUTNZC
q3c0cyEy3Yn33PEb8lBigEUmj5nXxcsu65JRCCBZ6vXSg9MWoXxmjYo6l4zuFjyXxtlppHlSMO8U
lNzPhGCLiizyxyD4yOaPXF8EWdY/WRhalFBu4AQxdvDEtJLANqeBv1V5xqs4kesMfH7URNpgK1Mm
mjjFR77md9Ads5JF5nRe7YjByYlbFdOsO7QDAUoFguLR8Ab/rI7nwAYPf7HRi8wTzbIoytBt7oUT
UfLJNnoKJ9shcS3Wuy2t2tLdex8iklaCgwumKdb2b/05BowHDyuE/qzw5lxYrR4pmM4fRBpIhthj
+rCqOaMcC8lc0ZtUrpgzPWVatuW/AzD7t4lgb/Rh8OEKapX9Ajnp4th31gWNXHTdiP+dse+ENd8O
67ZvUTrQTaSyqO0QQahFt8E2yZ5cHlPdj5N01UsCp0ZmkOb33KnBduloPioOdpbA1DpnXM7BspTK
Twf8QYPpzJFETsSYjZpBlarfkf0hB7YyHznZfO50L3fUa8n8CK0lOC2EfymtbcNnQMxe7cTuZZvW
+ywid2N2ZLVxJWQXqJkfnN17olmmwcSaguU4e3hCvoQT7LcjGHY/Ye7XghaNWCkmsZahA/RcWhpV
O6H1g3iMW7SJHF4junSES1nVvPoOgc5xydT6SX/yxDrp2hYbIpeuzFoWTeKPB5nZhUec8Tgi7Qtr
mnKtH3pJUlAxKGYZKQk3uy1JHzekpgEQagp80chSkT4+R0WlOv8MFQ3fGKhsOJE7Bd6uKpOe1OgY
fn4tnDDaI3je+yYVbodELNf6COkPYYmChLmN95wLpH6FSPnziWrmftM6iuTmNL91CCHS9kqEKABp
y7811mt58vwcXizU5P06RQH8MhOPMOJQjjo0box9EeRMnzzAbPud7b6sPVsJebGnL/793IDr+c6u
5F3EN4cQp73xNyJOO6XKihfka023XT/a9jVpS///XoBZ6Mxmpq9XaW/GIBxDP0xkKbuoRo8p3QKm
L2zuoZajjRb76404P4xemaqzb9lng/qdxmkjF5Eb8nSWnJSihCCSAtxxIPIVTSy145KwKn8Au/K+
3Soj3aYWvDA43DAlLogU1X3E5Hl4sPFJn0Wl2o/39mLWdU42R3aE914aZR2fVPjdoAqvpe0tSnW2
Q6lrzFSfKGDIIysZlvO+3hQB0/dBrEK7T6+/CzqPJ4jUOKA56P7wtwXhjq5CiANgezBm48IKHTYS
x59Qusb7DqMXb4s5hDIVzoFw+VvyAmrpLPxI/4fSmdC+jX8FubZakDBnhMJdy9F6uv2iklZDOxww
uRzmgdDdS2uI3st+P4cZiHDRRETW0v6QXGfdSkytR34Jm9R4DtZ0C6rB2vO0NjGk/D+V981jmwxD
MN/gwrxrley3b6MghIb24YoOuJw7TbDxVoR6TXe+lDSPBiDHrFm+8xgQd1L0SeldDHwrDES4UCd5
mWCeRK1uVqye27GlZSZ54EKWd8gKieXG9Mu3JDvb28tqMPIBKtMTeB4iGtm7k8ZwGv8+5Q6P4Pup
iTbNmuBVbYcYN1v3DJUom64fyweiobADHbs0CYsabbpYxjK5CVc6wxsFVyOx2oJzfV5dWiNz5dHT
dz1nyMnsu/L9/t8H+NUUGDff2/QcwDho+SQj3NvGKGXEgdL5YnCclS8mJ0Z4SJG6qx1bC9B2u2HR
+wRECp/Z1shlu653g2g6bJx3Gp7wjtjFPDCCkzOdygRYXXCcLIohIZ+/ieHC3lagJ2UijJ+zMVkQ
B445XfW1Wzo3OWJIzl8z+kkgTSVnc/kUZSLre7wroRmE5fPfwiAPzLD7/+nZGvFEvcQtGhTix4ni
zz5c3AynJwfFReLtmYtF8gN4rSPreRkcmRh6kc94ZjhM6yEh1PJXBRZb3hHzDoq4TBh/MgWdo90E
HjG+Gh9rXmGqaprlXyAuOlCC7RyS1m+3JglaCSltIbjmYRDXOREzh34+cO6pPmiLocbAASzolzyy
cp0wa8UxSCC+52IX/+0VlkR+uB7MQUn8q/nuBnayhCHHxPlT4f7rKCRG6QMh46m3zQUYhsT/z9V7
EJII/XRGAhp5mMThjrgWDO/uMIs54Ix1o6XzUvIOe4szSShcUKKAa8N3LIBIX5MdizUP955BrvOP
cQCiDHAGbl575XzvEJZBmGy1/w9jv+KVLAbu3OfovjD7R2GKVZuo6fcgQWGZjjR+7AQWRsBTqbwI
v1TZxAVDv3vLh2VeiKV7KlF0wXOMXISuyvXYFo5cLLeunKY7e2/DaoeZgP6scD0meXURwjiF9I0L
vvgdvxuPx7i0HwpW04v0D8+GkdpbRT/LGc5BEj3BGGeSQGF3iAm97YCzR15N7ZdlWEODWbF46Pme
g351t/xWNPTizVCe9PMhzRxWjLmu37ULC1B1KK1pT0vquL2kW1aG6Y32wOfCwdUz65qfbUsq/LUb
f/fd1F1cOadc6SYPwhhksomx5viiqlVkZVqtNrXa08LZKTv2mlW7oN8Tb0GurUF0okGTKSS8rJxI
0FjqBMwPKKFPnt4kj2kHlyaCKQ0YW8mqYEF9/VBGLoRXFylO2ocg/16Idt5yYiEYQaj73I8XxU2q
H7pTIct0+4rIKPmmyjbHDijdsXuIMdzy+R5MUjv9y3w0qu+n+wU3uCxOHhR7RM8IfgNBkt7HnMhV
Q6opJY0aMXxk1xkWJjJ5Ce9arNY7EyMtLByrvqm1+ZMTWxab9PV36C2YaPu5wCCDTSTH8I3Iu357
RNK8Vcsx8IivFKESiT5bJsK7nIfYSPw58mfqzc3mzCj+P9qMPMmE4teP2CqiGNkEncLqc/cloR5J
kDnLo0VYx+YrSZDqbCxiwFwIgWM3Zlgqr5nGux8skZNhw4ITeEsQLiStK9iU95mGeCtINasA1sQS
nMsVKf1NWpQZmTJk2IsGGI/CywsihPJeKvwTLz0HkudFxizAYVWvLgG8xrO/k85iLl4HpBwFh/sR
Xz4nEeqxE4vsLQM31Rx4BS8DEmVkRodC51A9Q5xqM1cQLuEu0htTNBLRgurmAfrXL+KJkvYWHodn
hs0mSZ3KDRw67c3TYujhCIv0PvrVK4OJA4SUBcT3K6H/D/hRvME/CBv7+9yClRgThjTalyZwpTWI
6aumvdpIrUu3GdKda/HSMzSDiZTomTcPenk2UkB53VJST3pdIax3BU+41Z51Fngd7v0bbPJAp+09
w6YWaaDlyFsS9+6e3lQaxi7ALFjkVo5jsTcaU+fJFrOzUB3N5ro3KehEQq012Vv1Ma8YuwcwL2pd
lN0DQI+kiBM20Vg+DmOKpFVmhru/VkUSag7DTTOVvSm5MOZAq8WO9ToVsKlHm/eA3MAR5KNKIlC9
/UsLWTz3rSTVzTiSdBYHgl84/qhUXsnI6GqdgJ23qMaHExRChsl+kL6DYCvdiDdkrCTSngntDjkX
uFt6nSePlh8T1Qdu8EWqSxWhNaPxHbNovom/cPVlrkPHduqhaF4tWpkmgcAAMbSSiCyMLL+cBwu3
K8/1txVE6xRnWz/v6QloB7PpfeBiUcDX1fAVUHbvcm6/By/ksmx4LiR2hUhmda+oa9geJQ38vsQN
eiGnbfZcg6LpdM9qIE0xQXc6ku4elZMqqX1rv3d3jGExHk04nAl4aHeJDHxr3O2FMKrUepD43j/N
M+fzy9YQX+fWkMiEohVDn7VuwSCfFqheDYkc2OIKokNvU/6nTsZh7Xgpne5jyP+JYVu8+oyjXFho
FFBY3C0m1e4cwdJphzBWT2mH1nqEBq58F+d2V6R/IlcHo/1pqstOQYD8yYMyCWi7PhwP+q0toPnJ
IM5oeb279q4OSose3kyz1MCMX4/Gr/5yxONOqgjwuqqrY6ZPB7ZXiGgNL9a4iW9/BkmGD7rSj2da
28aCFnXBY/ObpOtGUVE5EjFuH0nzmNEPjqHmvao7ws2VHs20uyf7+p35l15sYhiGZr/IKyMD16YA
Vbk5sERz+BHWcWQ/YB1XUUS1y69xHyx+gA1+PaeEczmJ6tRSKOT1ITBxMe+f+B9b6vARO9Rd95uf
ATo55R0B1zdXtktYuKPrrT5iuGMguQPgm4vQ5xsTJCdicfIVC51QaK9hWWzkZUR7YgOvvBuJd5B2
3KBRnLLN8ZVJ5e22PKxMeVhcFrYpaspSAd6AuM1JIke1IsWL96AnLXv+OoDBVdllpa6s9fCyRwSi
3M/jqFaN0nerL+BdAuMMET9q0cvWuFDIFW9ei3tQVE8bjDJnRvGP8P4URZKHid5jDW3HAqNx3YAP
EECfYPfbzsl4CvSk7xkccZ83K41bXf5VI39thMQD4mgC8WoUhP7tT0/FQTsqqQ34lpG5hzGjJX8N
ynkHoROt+d02CpCqbcRdp4WuhQzTVW2DQZuVC6iN9BWv6GZNMWvqYY8KxHFFQjy9KQKOee+rK9AQ
LqMlJhJyFh26Txr8BNWm111P/aOvtvbEhUiVjf2dTUjcEdtxXJ3lU3nKj8x7bb8rW6FpVfVzv45N
xDFv8HeSSggsY0r9zkHibExRE2sP8xmhLdSYywRPaax2D09qkVXHx4911kjg6BUvT8mDyfrFzBa6
e/IfxazQnRy9e4OEnmukVrl1EUvYO50vTyJIf2qn4hrhA8wkoUBe4eDLx4zH0cK11jIDMddca6gY
qCa0qD3nn5vad6/YT1V8O4r2Lq4BkcQnPf+QDjDzVGwm7CqssRwx2D7oAMnF/aqgU1wAk1t8Xp4C
bi3HU2jzq9ShEzEvVzNUCjRqTItE/dZsJ1PYXB2rqcEeqK5+S4gxDulcH6znyWpF4tJy8Ii+PFgn
5lsfxDzqc3R6O+GA9KhXTM1ZD48dTQ2mogetH3BnIBYHZkIZw0eNbhevGT9c7Rug7TineeQ7htHW
Cv+I7dnSla35YSv57WfefiypaSZprJQoDQMPaAi6Z3JyUsyG2BGsxBFNy2EH5UVy8I4/cQrJ9pWc
rNi/j9jhOMrEqxixRYQvelrHEMPKcdzp2obWdLDVQI0eo5bS79rc7VsR0AdnOgjW6A9pPD2ybBCW
LFR/xEi1rkPEXj0TMJLMhVE7BwS7cl836EOJAuaBVE/LuhH+Q7RLeg7stEd4sL5Lj1IrbGvId7bB
Dpv0sWvXoYUFS19zZh7siKbwagLkTSQYRiI5Dwpnb9sjCfwoF4dD1rnNrrOECJwgRZP7f0jxiSRZ
QnQLBksJQYTwkB9IV0cLwlafw/s5jGV/2TkYxUoTfzyyeZ8vbAFBcTZTexBO3fsZirSK31CZraPh
OC6c6Mh6g14TGPAL7/K7Vw7r223BEZYZsDVXCl2XezFkBsP2a8DsdICq/A6vMUv+5NblhTk0/X3m
x7p9rbwDcCIaZbCiTpbm3SwRn8NNfCoLyGL8V265SBMmdettlxyVjzD33Xs8SgwQj6XHhgIRZhaW
OUkCX98aqudkmyGwC2GnOguJPU6NilX1RlQTjVoKojlPahyLucqM4kGt28osKb7eGsytppTBOhcO
+mwe4rUsZnOFcuvEGR4Plz8qQkXRTLjLS9G+mj191C6OjBj/glIxTCf8PL1KC3Q3oUNHpVFep2IY
MEWxDIcMwGhTTH6obalMTkCJkAgXjQ+rcpGkTSLEoH1/9g4wM0w6thpzLyOGYc6bqR2g48plwBMC
QiXz6xNhdxXF6INP+tfgkuWonI7rz7LB+qjjasYPkeq14j8BSsoEm/p/hb1CJHeoHsfkSZiew1n0
zTvLEUkRYz6uNAImAJ3lVaPduHH0/cLegy5ljMQebgiYT/FJRhfaow+D+gDhHYQxAD+LIFiBWn2j
6dDTvpX3rTvE5yjxOk7+IKko4I4d+NpMdprOXwSKKqnfNeQ+2d0UGas/b3ypzeZEExfLZhj+Wyc3
Io5P71lLzAxbKR/xiNkPEMGQf8FDpESVRL5cV5MR5W+mJmIjnf6tBlylelZF89VFirtoRvUxMuPa
j5vQKzq5EdYgcwUr7QV5VaaoemydjyzBcH2l49MTNTEPaf5e38tB+9W6+eeObk/nipnTaJx2vrJM
rolLEqU8lVCKKGO7NjFjjXoQsHnLFLwJnE2MMXAhilZIBcjXVwayb6nal9of1E9FKzboR/vQnmiC
YRyMQOYLRWrTuvd1yeujdQ5Z0sUivWbZW7xxaJtqAxFocYqCl4BmegsuBcfEDAHv48mz2NVQKsNx
GIevp9z/2k324E1lAA/geFHxH2Veo1nEv+Zc8DQ6ZPKrxXKYpA1HgNa0QLswLwCLbgbvZi8tweFN
cEQ94dpthbGW4WdlbaecIIxpCyAjBlRJLayTAXrMFJZYaKmiZAz3ef0uWNfTW2ot6gfGZ1k57a36
D73usRFRriI7Iz1UNV1pEs+/dvMEn6kbXCX6x4pJZVfGgYf4e7uqEg42CSIkb0ll1zi6w/gycX7+
QH3Kbave187BxOgI0MklA5NdsgATop6gHXWKRw4z1qm2K4bMByt7KdO6nPC9bSbgcAMqeS82qrnb
QpBMbmakmLC2Sq28OUOjD19+nS1fNPfaHooIpmpO4yFTSTa5pejRdsG5mmW1VU04LvyMjKy4XG1l
iV1u7bNUcXMn+JehmX7Zns3Uv7MqWWD2KBOT1Z3oryGK8X4uj7Yks+UzPS5Q1fdSNjoiFoi3qySn
c07nzk+8T+jqC3PXs/pOj9j1xTlamvzgaFtvbUJl0rS0o0KTVwwhz3wFqqyT39VpTYEUTpjdxi59
1gyNfIa4lG2HVyVdKqPtk3O+zaNa5bEviExHxbt0pjQAwNqleX9uVVNbl2C81QtcDffFIOO1XlOa
7iXwYpJn2azoXF8Qyu3l6LJat0Ijx37tux+97hnu5QeHQmzuJakKXgxJGMzv8vEMppeVCvt11JYK
Eh7n8CEg13FVlYICKzGWFLLR8+zlt4JRiIvKvJIr3+J6P1cEqfbtvEiNWLCepKKRhtdpqDb65WTq
77JbTzjJG5c9OJQ5nMhs1CBffAmVCCInBdKrP1UIV65wNjFrgXxQTqzZB7tSu7WarhYpU8xQox0e
Fz/laMo7Q5BeReZpPAFgIebsvSuHCjjq1i1k8MvjdEX/Ij5O6fi1XRZ0g8VmnFWnTv0KsYPbdaSW
aBbWDQeGkLAfmP+fiFuByr5j2EhyVUWMIlWBCN5m/5ZE1IJCZnZcjipWRnpQDAzkFmcVWLk8eLXr
erQhCDGFFL3covhc1S4w7PnsRVnd+29/JvSErX5IndeZoWKorbcx4/FUoLonHUFGNIpKrLEOUudH
rEdyygTJHV2O0X3mlby8unT8B8l9WNTXxyhyqg6hA/j5UGtS/Zq3dNLglRT5ny5boM4DDUK39P/5
TX4sXHPyWgXOOWaMypJf4qNpK8G++BvY8DUidtEUAGxeW/Rc19UfCwrUdANlZNNb5hO9keGNvXlC
pHu1wggTc7L++RSILbDdCvhPwVFNkQ26bGztuAoxvA2/D+XIonXY73NsEGoORMdigp+Jttslj560
gInN1S3otXxwpCRTacFuItxUqzk97REeUFig3snHSDbXRPvXcYfcAe/hMen2+zUd9TUhpctM4Zxl
ed3SWmco4tDcE3wAt2w5HwG1k6SehSkhKnwwKKCXBo4cDikEH5JvMuInEbLOYchhrgs20QIppE+b
ri3WVpSMOZnrOxmcYAueQ4ao/mwQLnVFKnAPJ7pf/AF5zRjFDMKuScJwPP47TqTJAqIkNXQ5VbXW
QZNbAlimKWB3z4IEk7LWgECnhUtusNKw0adznU5zXF2MpE0TJJfRLm5Bxehd6bZ/hke0/ikkZUTD
wVqG6PrZS/HhMs5XR3udPZ4u6GbvXMSnuP9SosArFfQmoq3oC13Xh0ZGYGJ37G6RCLX531oW9XHg
AVkNoGyGp3KhkdA0l+6FQ6vA73jogpDDKgej4vwzxaADX/8ejqT6VPOdKE539+Ew/shSmbkwM+Is
5LipXOhXoXiSEmjmhpmob46wSFWkssk1QABbKV6J6jIG587XjO7vVK4larl1DErBhcvSDm91MmzD
+Cttt0aOPdjSjIXhoWhGGwwKe2byvjz1Yf61PYflOnjqVRP05WEttaN/w8zCdY3JttO3TV2NFEr2
7wEUKdgxH1MFFGsBZotAGHWqZ59s+dVPzbEOuILSUJmB1RXqox3mMs86lPhNg55Uuf4TdsH9etk+
P3HdC0/xikbJCcfC3YW1A6IdTUMSIWXtUtWlz8qbb0kPPFG6txVpbe9NQdUdTAFbtUspkEYAObfM
CzWD8mUFgkMYhkFWpGDkFZyGrPFC2lmCfvEGvj52mJQG0/A2joYIGStaR+sxQPTlRPm4M1X9zRvy
QFpznfbR0AAVLj2MHMrohO5js5wTXggWiFu50chXGbpDBnp4jRt0j9JDxURyWcEgz4av3j8VY2UU
yylQCe9Kg2JABp3w7W0rXlojLeLroJP8zo6hhg2Zs5X5ldzaPyODRzHytLL1twjaY3ZJttHIwbzD
yp4H6DhDL1g+2pu8hTH+u8rAz2NjWdQTRCdsi1vM9IZcKmihK4b0pLMGlVuyVLwWqmTAHz/fybBg
fMZKb26cM2LtGRL5qYKYqNcMBgq+kJVJOJvhhRrcFPhEGKHE9uFCUiFabKt5VvT11PCJeS3v7puY
4KO8Em6fk2+sJUay8b1N78Hfn5csWCLkuF21ksO/eqJHwxXLsDUvklrbIv8YyIArfFCitXRCzLfJ
Ywi1bRktM3Xqy5mY0aE3kDAIVtadUSZlMTibXll15SXoY/H1KdTijS77xu93Tw72xz0mqeUefWw/
BmmVWuVEcFxWIlZLw0l1ByBNmqFC7JqnDqbriaXTJdbl23rS/6e2HnTfC3QvsVyekeURKjOsX5oA
HTIxEfZs9taSua2HcLGervjt6dvfJ0+OaoQNpCckYIcWvE9Z6YuiVIfUD8dggvHAxoLP3tk1Ft5B
Q24qE5tVm4uwk9Eg3toFDTGLM0wZVtOr0AOiTjBSTF50KXL5YmoNm5sxIHACABpYUNLyP/zodcSj
dznMAZj8q79sxU76yyXX0uuhEXABnzMc1kGFE9lcTsCa3W8i+99W1jNozsANiOnrz3MocK00u+ka
Mg9LvcLtaYcYtULrbDzUTOEGxj9oAtcFZZGzpQcXNq/N5Ml53h8RZXAGreFEAb9dExflW9RT+J5O
MMDfoRYlfjVXsWiVsUBzNRSvXj323BfsQzJqs8f8Rp02TkWoZyIZ1uOho3tSibSAWSCUXVHJnVmf
HYmzP0U4cXZ2bCcORxr+SMkxru8EZ3wG/t8Hz1uddvCG4r5gl9kgQ/rPzQasxCcDHH/PjCDKOybA
BApTMgKmuSDLnHV1lTRe2QvvY4nL8bAoxMRBk4DmsqCZeysD6ZFFTMifM1bYR2hZCK4BDBHvqgnt
R/9WsYPHGNJDNL0YSSzN811adKyWw0Rdpdu6kequBAHXhbGgrtUoY0uwI7s9ZrIeWmLnYLnmd7Ai
wlyu5LinNuuIV7b08Q8aiaGAsd/Rth/vkbngXNmF7v6EkqFU8ahl0P7Cdn4Fz3XLDgkIjUdBiiEa
+VFmMDBQ3Otf6VVNuDigZ8IjnQMHA42j8scoUBoAsV//GVawgDrJYylTj+Z9SgJKVL0Pdb1nf+1U
XgqQvZ72pA1MeRWx+J6rYTZLCm1vsiRsjJ/gxhMYtdwGhr3o2DBgQ0HprznrDZQbNSUZr07NY/wy
IErWtxZ+5YpU/Xs69As06vRdwg+UUvIUb/HReA0otx1oMUBmajYWugR0OU4L0XEUH/mUjcONe1Hs
8Jse2AfWpqme7/WzizlYJLOGkCaAyCg94jvZvQg8QZ8xltXgoUzgEfoywMPeWMsHBCdk7/NtFGQB
KARjTuLgTVJ1iy3nyQNFDnBaqy43qJ2DF8FENcOCJvgasDTbP06PLTj15fV9cojE8vWFxfpYQqfw
U7tZ4FOfuLMcjBmr9o+y71lJfog5a+sn0vzuT8ywBiHQZHO9WDM+hmCA1ZRK77mofanFRekdlP4i
GuFtqt2LgvZ/JbkZfwwvsrsDtI1r/fI2qDyFocysdI/CbbOu9QWK84ucmTo0C1WksLb4yo8+sfTO
43HDkREUQ0LZki4xUqzJlxGAOAxhbmCk2WgP8O9tix1q9s0pngyQ/NU7Ht2633XztWzhcFXmPW2K
GCCYBZKXhv8Kung3u+IOmt6vZwzGAOMgIzJFz4ibDimYFOxno41bo3CYAMTpZfsiSUKlUZcU5FXk
1xco4F6tUhdMRvjtIy4Cu95hmrZgS1jL3GCiebfAMBDycbRYSAGZH6VcSOWtlTfHOGxtx9oB8qGA
e8YfAhTQ6U1fqK22D10aZ+mxgogrg3wHupd3RdW+DEBkxOXwtrEvirIWR7IofFJd8Ze6GtB8fIxP
xiiAc8hkTiABmhWwydhFXk3U6y6mBABviIiVJ6UShmsZy35v4Rttf7d9GVoT/4IWSakripCgTx/A
f7LsuY+rAXuMtMNhhxVaj4TbtORIUzS+7/lQ5SGFIK4B6IHWhg7nKfr1q747xYzJcLcG/qsPEPbY
wm4hnotn/txgRNThMKJyKgM+8I7JFFC/yMwbQe+ifDmFdsgKXAxQbFdNhZ5kFKn4YetzCejYmJxz
Duggg/LpftO4nPYYGjLEOfZ5tHVyB/KqSmEsNJptPNERjJcQkCD9xe/z8vW533h81WplnoJYey8Y
8eiH+6yBwbWnfOueGZdGTKIRmt5LrRV5QHLWyoSI5ljr13RPcBCu2p7q+rborqu0dRk+AT3m8g0t
NBBq0CTG3t3PYHO+LkGW5ODAv5KlYGPlYfLZ7WvUdvS6AOznZqfBM5CCrKMcBGBkwRLdJy112g8g
HGLtnPUeQVXZSAXUoZ7yVAD0SvOCEgf10Ebqu+Xrvanrlisla+e0hQ2W7HgRoItYYvDtHIfmzSNa
Fp8JcHQFUgU/qNo3PBqpGRUozMQ4AEHj9JJk0B3gRtUuzO2Z+uT6/nD7+HCvC2H0Ht+ulSSX2JNw
1Q2byhbaAmK5KUmQf8NmEeD5oB8XhfGj2zJPfPkRNOwR9GSsp4BmvqvI9b6G09d/rCcOv/8c3uNB
b+RJ/Da7l9JBj+8Td3TWFSL0i5+lqAFqzIYqSxatzYK3N/7gkKzxBoGVb3CV68FxHneG7xNvPNt1
ZKUXE9few5XDS9HPZauRWHQYyY85ZkQy/CD4smsMIlQHhIMrFNVAIgCoESSKfWLNOudzbAXUQzM0
APRrSl57VxNSCTTAl4M88bdV+I8zBloMAhk1DtG0qhZDMXwWrMDUI+w8cD2Th+cRZiMS2O0hLhsp
Bwoun177UNDjrvlrr/Y5ns2dIt2ONzDR2YQsXsLKkOdv7os7H32FI8B/7VOQQfQN6BhdtWlwUT3l
ARavUX6LqIWMJ8BsrEJRhsrvGjQIhkY+G7TQddXA0pDcLt2Z/d6ynp/cUFqIuEbxa/npzzMBpYMl
DMJb2kZnhH4w2XB26lzFhjVUufUoj/ZynuTLq0J5oRDqAHXFnjPRmCO1o43wgRv/hyhLGhaENUi8
5jiaPctreJAvCBJZh9GKRbR1GbDF/7kg/Qce2YcGHi2ybM4qe8NxGMZci2eRMmPdRgtpngQEIRpX
R7bA5REkcdWhZ/CTJ2hKoiXCVc45BVNSpP8/6dvcjzIwTK99SToZoyz6yB+lZztSSKr3kLjARgTp
qEorUgBC0A+KyruGq3JPbW5QNXJrZml56gTcngBM7iahv7oEp1EtqZ5VtGdQpvAVjYmKcYdzZtXK
vNaCCYEK4rAZJQrawNJGFFzJzJqSAr+v5CArwNGhasdzJ7SQ7/Hnnczp+OE6Ml7DDXTwnAqDvMbI
Jqr7oTGy/vZ3O+biHi3tXHyFSbW/JCXMDl7ifu7Vbbvf4oy29WIbb/sp9leRnqEo9khaHsMGxMo8
USOQo85hDRArN/6PXG3B0mP8j0HdK4arN0rPJ6otsd5EBkmhf7Av4vARUeVklbC+LiQ9YNc+h0N+
Z1Xl4fbdlgg4GF5W4FhKmZkrNDbdtM28/5Q1x8/D6id354Ss0zQpe5JEGxvg29LVw2ub5MAsVAch
cx/G8WFhHu33jq4nMcxEGwwucrwjNX54lNqbzSmC+7pJ3/E1lwKaSvsNhEsh+JzEzND+xLSlELkU
QsJvEfHGaDTuAoyKwB4Z9q1mM0trNmIlyaXVnbHNzuPs+LCGuTICGt7L/jl5GMqjzusXnFbP+X+n
C8MY21L8sy2ByolfNziXNpEzSRKZQWQH6DNIS8IFqZh5+4Yai2L/6f1/rqJCsDn5z0jfBI8zTCxs
GuNCJx7BQKsC/ckkMQnHwlP7PpzPs3M5yEZghdbhMeSq035c9K6cTZ61m3zCBOinOhfhIwHeOLEN
+Rn20KgwhoGXoDGniNUBCkyFc5Kaj43xb2swpDtFTne7l7/ve0DbS9f4Z8oXD3aZhX+cRNxnSt3l
RBsvKS77GSQ1vGS3wjGbLsA2qtdf/br3UtaEk5aEn5hQHamUMBB8/rNOvt8sjRaNrz4RkYexVnuk
QSChvosg228Fl0X0bJniXACifH75BGf1t7kWlK+bvKB5e04tMkTUKkLw5+h/sHuOX4tSfycC300O
f65xLhXw+/jN1JjA1vGHiwnpnS71O95ECvOQaaLn3iyEZ0cKkgGsp4yPWiT0IUV9/7Gajl9r6jfS
erCIjyO7IVYpy5CQ3z42bLw+722laTugaU6H8Jac4Rlc586dYnMcnWgyPg7FRnDy86ckyEAROBTj
Obt4W4Bj0udf6fQG9Q3zBBwzoCTiAVVHuz/tqE74MKl1rO3YBUpgwpzEwecCQIOY6yQeMPw4Ul7O
iu1HIPZlwG3MeAiN45LMRfNwb3TPTe6njYI45pAUQ9Tw1eupd3N0g802kmJUjDyt9I4S5rRC9pEl
r5+qNKpWad6G26VH/06pnXb2Fu3qeub38YjJxSZIrs9NFGMWDn6p/H5+hHT6eRh6dQ8hf19Tctxj
asD2OB50tDnOVk/p5F8tD5cR3Q1sTfiV2GTkcE0o9ty/1kPe/ydKyrgadXG8ju4a2T22aZx2JI76
TFs9Bejgn27tu0N0cKxU5XKVyELCRRTU8vtqv61r9SvULKeSBkN8dUarp76zlBmsC3w8sr8sbwGv
afJj6D4G1h+N3f5HcNll2KIP+hMxzR708n23f4g430mk4welEdY0kyh0GXu4YmHbByZ2U57tXkHf
wcdHwUKZ+j+9VYhe/lehsrSz/UUncS9aUqx09BBLJUb4cNt3+JJN6l0BWsv2bIWEi9hW4alao4sL
r/L19kkkPfSp0Hf3dALZAbOCjBqU6FMByaQjaIK6fwaccMJIAtqX9CoxZfbZS5dmIa10NS0nU5e4
PRQB/7vDKT58/3314ayaQ/IBpLMHqCs0F2zU0yT9/fiANNc564iPnsQq6nlyO8qyS4OoX3Wrkw3o
PRonoxPHLMVA48cPDXyflwZi+ggS8vCf8rpEzeyOmz74S6Q+IU5FGn8Idt9ee6s6WUfL6R/r3bGJ
ZDLHyfxY/nrDOFLyEyW/FgoIZJ523KcugIX9daP8FEIcV4XdnVNyYlDj7wjve3sK7iuGnurG6WjE
DwvgPgl1p/HBYdu0SkIG8SrLf9IKVZLpcRJt6NX9j+n7CF7U1RGvZexcZV+Z6Ec7mbZjh8jvEWFt
lRXU7bgvXa0eks3rmBaCbfr0jokj2V09rVDiOumXX9AwWMgNbrD/YEUtANj9gBglL8gxwKfEm9F+
94xUt7VfXInaUyRDzN34IWYdIWFXlauMefeWcISxLTw0I08gzAie1RczJhcqsmfQMYwHKVZBoeRn
uI0X7a6OhfQnhCBo49+oYlgFPHNeO7frzWw7fZhPgXxL3xA6JtmBBaqkwjbcD56EJnfY9wo1MkAh
NzYgMbxEF3Z7n2nfKf26vfxRZimEOwbPVc/OaWIB6aBrAp3wzQaHqeuyVlf4xpBY/kC58ScuKoVp
t+ruS/ipQjZJQDXuJrSK1AWNFIt1GbwYlLlbfrSO1bLuyFpQkOpz2QG8/+CNd96BQ73ECLqkEN3q
EiYZyUQX1yS919wn8BPlololduP3ppqYFbQNGQMXA73orL9ocwf7iWA91ioX/IMmlEnyJ7/4WQ3Z
9ChFx9u8nDxScWSOwJ3wsyc1yvEw1XdJSKz1dQDpaYGrJwAQEw9KZmVxuBSmNwsfXlHNFkxpvYM/
J477zTprB8hajDOZs6gbTRP3ELc6uZ64KYBYRKGgMvfN5I0zh1WMwBit2ZSu3BXdG2b3aGZLUC+z
7kBx9Rny/vh41vE0DtKRrBiMTSMADrSryMwvIZVH8kMDeSbt2QCURfMXeNiAISGImX4HSL9cBIAx
/U/6KNOoiddoNOAiv+1eO8cwp3ek11YZjr/hbFarizsCqd93wPAN3dZ7GY8JQw/zedw8yhh+NIyt
lKD/rBGS11LDNuHKti5kGDTJksSIFhj8yokz/QObM3b4JzumeQ312BmGm+Co5HZcHaovoM4equS3
NN3LKD5qOTL81FSGPJYzvPRYw/CV1TzdWYOpg2sCGhoiAP19FDuU4A7LaX16RjeMRL8lHK/9zCWg
LitfMawbn4Hba0ApL7+qdlZwIq7n4amQ+EioW7w4lVl1+gDnEXNRRjVWnrnEEtjyg2qkyloSXzZs
ShUO6I/ZMJbsxSDoHPtaNIdTwKbOUKDhbWF7CHJlb8A+tvbadHvrKsEGBIHgnZOa18Xzqz6lHPPn
xT2bchkny3eiOXS2w/Hk0oVK2mBfk/pap1n2WyE+0+B6GWk5KUJrGNnEJYJM3Lf22q25h1tsD+mZ
5M/Sy7D37jV3+7NAV6msgEwoaVQza1v5G+Zd7oWefOoavJLUcTfsgzT/Ln22YPZQYpa+bI92LBnH
6VoTVmERNlwig3TskvI1V+fnE5aGNgrt+3mpOr4wAI9ZgWcPVfLmzZYqJsj07UCM2ZM6nC8iwrNl
DWrU/Z8LRvB0vLxjPTDzJYqcPVaIhIuq0mU4wVDmg6RBIyPbmAmAWkpod15BaMVFWNxsEo4yLg/3
4Biw0FVq48Ed4mP6aetuQ4AUKCpxnQ2DGs23QmFE0JgyB0lmuvMQZADOenjDkKHOTYtSnZdg+dJS
uxA3O8XW8Ux6qqPEfr7lR4CKuOGtjM9a50/iL2g78W5ngVOP7eytvr1Z0RT71wvr5cQJuJeN8HH+
+KA9Gtt/uSYvL9ctr0UMCz72fRESVAFAp9QnQv7NG0uUCSJL5hKXnYfD4GSDMXDkNFW6UqrTvDkP
o+09YerOFXMIxwu0V8CRWF0Lj0wv62+r0Kn/jCPJoGkT5T9KPEM9xBrlTFLh5W4908fPPDHqgr6I
oHXfYputTZVD0ZXdNo83CsSSe0ghloriUhFsy33oodiq6fbtt9j9DSDOkPUWTZg/uBgYyLmcGr6p
yD2lRj3IK6r8mzZc067Y0uImhXtvDz0Fq0PwCG49Emfrb4NbOLLwxxSbPE0vjq3pWMybilixdame
ueQ6fGbjeR5Eea5O9kM+9lQhMIR5s/UhWDljPLT5DsWN1265aqQiTBnZEQAuEsgPI5X0z7IBdhDA
oBZ7eta2c6EGv1EhmfvxDSorbv/j+fXwSAbYBGCUVsXkVTWYnqu5ec8BWhxdQ1fuyGbmXDcvcORN
8ToDgZK2yFbN/neblUzEKb3mCxqN/BD6voPchtyjVBTY9EwEkCG2rkvx1LedcWHXh4UDPzhtyt6h
cH2AmQAimR9AfA9AFUIAqUOEkdv9s5AhFOh1aoPeArqLVMVcCLKEPWGVbADdDYxHgyOV7/DK60BL
5dtQPK8noII0fSzZ734NJ73+f9PeDdSKdY/W/gRjWraHMzofS3DpkTzhPQnAXgkBSiZR245LUrwe
hBSUC7hyzprw9NJq4VnjlXlaHrV2qmyWhgor91kGFRXQBncdnytlkKSxMXDbR+oiI0ymOQg8deC9
8TCH1/VtOJu1tHeWby43sPXgPnIgYWgRz+i+9t0c1WOgUU/r+SdFzCAzcQHSgOgIEQY9WOYQWYQE
1oWOv17hM/6aY5bgXSDLAjDcEMqZM7jivrQahEE45xohihFiShhEIuG2J46M/D9jBdGFLTaVUUhe
VQX4flF8tiLs6KNjU75WqwYLI8qEXALOPdW90aigTebtMyDfY+dhmbT6wDYXUEwDyibJc2eqV5KT
kaNv24BFVQIHDdFqyc5TJ9v4/MISikfNuGYr0Rsg1Kv4kpYBLN/P1QvPTGf+5QR7vAKnsnku4vb3
hhz9m3BNHJn6No6T9PHWkaCL1L01UHIi3ROtGsVhXl2YqbpssZ7Pf9E1WeGP5LfAXkqd0Hpz2GnD
P9QcL296CAogrEQlrIw1KH/2WfPmTvZtShzf0+EN8f3F0lTS/tbuzYpW8Cr75T425ZzPee9LvJNM
NyaEqDoFBUGzcKMH+rsJfi83I27MfKpGT+B0+MjGdDDokqsQuzIlKOT3+YytARjyfIninCqvxz4P
/Bzp8sv9S/6L7h3BQSYthICn4BLlTYFmUam3J97pXUr9NGfP3tszeVorF8HcmQ8u13bkZ+a74PfN
16a4ebD8p13ymdWK5asWnpScxaaKWZpkSMkd03Ti9ENLP2NLO0374Br4puRqBB2M2NiDP3eCUrrS
Nc096wqLjyOIqfQTLYxBY6y0HbMK4W6n2mXhU7HrQT3+s36gY8jmCE5+ieO9tu7QgHWAXI5S1VKZ
ayV8+vvUwUBOLIPr/fGaMgQhZXnhTWviPQISyzQR0zF4za0Z/yL4cLu0304zxM/Ozqkn7oRmzNDs
+KPJDW2Ns7Tl8qVNhL/lH+DgXgyjeWCLsLmYSyxVWlAnLu29vRJCXhKNuCoiRnfwJltulg1NdArD
DetjCh5x4Zh0ejt3mmWBnWK9rCaqTjM3h4P91IBCw9n7VFftzhdomfy/4VN0Z87g0GsQuGOlUCh5
G8DA6b3F/+e9R/zC8rFmM85TTkE/Ho5pGBAxCId2thgWlxIYSWfKdJ43grkMcFwrB25/Sn/Kcn1J
RwE9NwwtBSE28SysR1SKDQ2PCl9Ic3EIz1Ajixh3LNLDDquyhAM3tzBWXd8DjifO5iFGKGNGin6R
jEHW1Sd81tbhaMjELDFsBBxYUQDrR99x2O4c0DhFsDBQo2FT6s6v5B+0hI3cIz4HKryhf7zX0+q8
kLkoTE9FsMn36F3yBcUz7/7xuEMHj3SY7OI/V39bX/fMn5q3BU2C3pBwvEEwha/PONLTXkwU/4fL
lE990kA5A0KorbO5+7dXHH+LXMZdD+rNXdNUQcDprnXaPkiHrStmtNK2hbkDl0La7LIQPPRDC5ky
rMH4X4y1jn0vxZrvNNg9ggDorXYUK8iGbMnwIX6V2YYU1QfrQWM1Y+LXj+g9sLVRWftJYihhTH6/
lEysbJrvnBSpUIYehsO4gRaZiAKD6i/njCGlcS8kmQAwTeyoa7OuQ1kP9ik7R9yLs/AwKtrTqYUN
fE/Hl6yP0n5Z2P+W1rS+Tbh08nLYjzr7epIWhjxCfNzUys/6Ze6q42R+UGiyZhpfWAu4kI3s3BZ/
PxN5oVOo32i6amnSCO4x471Oxu2fOr/PRaecDJ0tcol4eldRVFxMdTATgKXNi8rxQli+32VF2krX
kJufGq/pRhwWTE65LKj0rfgHFVy22lh4+cPlmCsBEkiDKR56h5brO7YMvxruRoOUtfDYQnB5CMgV
xccTokYrSaw3wp50PRmY7QlpGHrAZtE+JvmWumkf1dXKkWLE2ht8+uRVtQGdNUvGV4gM//G8nPaz
uD10x6xNM+kZp1gYsh0sDx109CLZVQQ8BI+jkTW7QnHoFNAM2GgywvFthS/ZQ8hkhZhpmWugjlPX
0n+1PWRB7DTHJexBk93ggm1dpVIC0cp65zli8h/Vq73JMcj+FhrgQp/czvX1YJCR1q81D9JYcalr
O4Ix2mhHzPnlkXoqjqNZNKQQqM1f/Z3JrB2zAqGWmeDKQAWGGDSOf+f2+ojZTp1FibND3SnoyOdM
pKn3ty1fKn12AJgIokd5lCPKlm7Xqy4MNLPZbeyoFfCUcTt0JIuQ1bURFmjaJYz0JEj+y3xVUjws
S+mZNKrO7ILOg+/KpTIv5BLRuyJrHiatrqzhWYX+oqGVyXAm6ZC+LABbhyXU9sxE+ZraIEThHubz
ZdYqstA7Z6AIjJCUu2YcSxJiWOwhYF9eiO/xK9OaESDNEHW6J2IT7lP+87JZsrsaWighfOKgKKlU
/ln+vlQiyVT8rzx7qZnahTJyMJ1ntwtX0KBMUyz6BKoxIlE4TaY4dASPo11rwMnwEAKrKsYfgYb7
yIFUdbJGI4S78qMEbYsfo+onwFHmiRXoMtH8jIFzf+ZJFa1lUNkfyQkSAHDGSxZFEfNl6aWwlHoh
0QbS2+lioEOQjK9cerX8vWaHFqZQ8wzw2+uQQ6ZNLDF57yFr6diD6IdfXXs87T/6fQjWgeilmenN
TfDEMoStsO7oDilwHloNqQnprvu9pQnzUFnoeBaiSJ54yU2yvU142/0dEtzoINTD1zJIplZD7CG9
566O3v+D+8JzzT0IGTGJ5OrOHTRtG2j6uPyRXha31aqSptd6HiQvc/Q4rw7qEk+s17mESlYQ6Iuy
UEkh7/ZZiPzUaRtPgpF/X3KxduYmPz8pIn4wcEfNyc+TAQftMpOsImzo3DAXmmbC1wveXV3ELzvT
sOFUZrrltR6whcTqfNTVoXm8PDXvpj2Lt6Tu91a9ukVGyLY3nKr/DszqNCRiptStMWXkJg2d7Vo3
uFRwzWE77IVeQyfTmB3EPxE8mBCHTb9C02NdUkJ4x/mNDu4lA5mXasbuTsJ6daQ9c6f/DZOdfr4U
BBWoLFTQWg8a+xG1RK/wRJAMQnqWULHHi0r78/DMjkF/RVoBp84GYwCDeNJOKmX6XgpG8h6GHOrN
SOfPRhukbSJVu+u9OaqVWYaqrDnxTSXv9/gBVSFJvpgMg5kXYPgKWQ4KqaPHFklVOl6TDzLPNJGG
qgiGQqrSHmoo+WnYyB7Hly0UsG8mjKz1ev4bFdPUbX0BjGAaNx3o91+1iahhusOOkkzd/yQ5w34a
+byF+lpiKgrtLQMWMw/G3jZRKjts/MkKxR4sy8dCRWV4Nr1nVQ7QP33oJQhQincWxI1Qsl/l8lfv
GBtI07qL7y8m8A+YJ88IkuRBfV4oXL42YAqM0kEYzakP7+UV4c+Kn81ugtLBNFiagYet0Ypcudxu
Jww3J9VC4rX3lzAfqvL7++Er9B72m4t7M7FHUWCgMkPKPdzgdBWBVNLECzndwWoDkqzyBWnslRvW
CU8nGKiyLm3/hFz6YmijT201pcrBA8m3ghYJA7u47jb1J9G4cMp3waBLc+tCz2Nd0vGsM/7YyvSx
oNz/MWmc62AsX63h1TeDKg4rQmHG6Fp8iQbYQx9tXJEW/z3ulklVpik3TvJyeqy29PY/4Q9Lc9mV
A5UUbx70SGzEp0Jl/ycvvdrDUHCucyMA9SI0OVXErucIx66x1a7CDMPqav3XPpt9BU6WxBFdBfqv
Tt/rHsfg9JPEaDvi+I+IpFvibCwR/JCgDCReLnY6LHU/N3FoVvwm+X1GC5pog4sH81mfBRck50/X
wYcqmHGe2/fwlGzskJ/24nxHQoTnexCdHhIW/JYe4LzNp49TxgwUXMUa2KXPmrFczZURs5FMD59k
AKLHAGENYqSZpSF1O54PpKVgRoDOepmA0a0KOORtTGtP6P82cVC+If0XDPDXo2kgYenL5ftHfGd8
GCVVqdYm21pytb90CS5s+cAUDBBbG5EtoTy9kmGn5/XtDNgO8v6WLFmQQqlacrFcwb5KUQB61k9B
j3ofVM6laGtPZGg8LRDpwtB91vHu1NqVJ3WX+/u6M7j2rt+y8xijt5rBaG+x0Rdv+uZiL4Md50VQ
YZzYO9a9PsHEhYiX3n49YLlrV74LIwE5Pswo8xRk6QOwI9Ad7JneCn4apFfg87kGgsXjLYckUpYC
3P7jYPv4Wh5aeYfaxMiiU/tt5axAqkuy3HeHiSXK4E4flnQVMfHT6QgGkDuIlOil4apnRkbj5/7I
KfQG/iadFbxAS5aWTPie1PoNfToVtz3KPvn/hW0joyyq0LWNv5CujNmv95708zUwQNxzKzJ8Vz28
RZ2stT39bf3PU8H7ELe2zJnyx767A4dcAr1OmPyePln5BiikwTAI1Dkp2tOWaftKLT5Gd8LdXl7X
1GckW4Z7qCnhatnhG7yXClcVRTX7Eb1TxDoyHBWNZP1zZC1+dlMNxw3isAAOGbN+k4oPvIpl9xmM
GoeVkVsdSjuddP2nX/iXfG6N1aQfXVunMPHrzDEoIG704/fq7unlCyF/tk84f6l7FtyPC9hM4s4H
0PYyL4bIMgaafP8rtEammas6SoK4xeoOCckNrr8Dw2WI2puJxOVPe58Ys9M6cqBjkeDXXAblJldm
nlNPJsJJiQbcsuhtm21cnFiXbsyxJtezyXu9gVE99w36Qn/78DvlcqnfssDu3G1fDQoLdHgbvyNT
F2KDSGgRUBWIVDW+wkcmhhnSSITQLCzHx9OnJS9J5OEOu7FmCKlzu4MWedghX30lKLxOZHbbQ8Mf
L6A4OJ9JAK9Xdr/ZXV1LdOYnDoEf4U3/gjjDn87U9ZdUMrCdFOtrVCX38fJt8Zymd8zIcTvqpgz8
0TYOhpaPk5KuDK43plws1bFKWhoFtGXvoziyKn+0iXl7lYHpGMUuhGWx84paCf6cbfpNCvhDkKuV
zPu+LeCsmhpbzVQLqAN438cfEot+mY2lAQGvzvYu7xx6h+WTWo3V0LlVKLNc1grGVsbgSDbzyjVv
EkDP//gfhDkEFUsj1Cx5nwBywPG4kFz0MccA9ZSl97xmTznURv5xAbscwC6T7WwcpTJaZVeCYIH/
yBE7ErpuEsRXybzDBum9smtWYbmZQir6JZs5xfzaCsnUfvy1FA6Y/8zPX0yf0hccPbnkRkRBYzok
2CpXH2NTlzwjmc7N5d1XC4y02KEj/NqB/9K4TzBGvEWuIB/WXbYvkfEUVXXQSbjDezJWlTIolgrq
Y67r41zmCh1HySzRBn6rCZ63Az7lK66cyW/V6ZIjUxPalhX3dxYnLQLk/RfiZhYjcCxZXA3+GTjR
k/t8161n1g1oOT4FkJPo15ScL8sNhYIvfzaLbSm5kh4ll1BY90RAmXy9VRzqsUoXUE/gpSYTHRUp
GpJFARdYnSDIXXoiUb8HSxVUauqpi+jcjBJlEMpTrGfrjSLLqns9+ZgrvWRByThtU/N+2SAov8jy
iTJvZK9jVWbSZiQApujHQ+a9FrZr0rWKuOVhZSe/euyq7eovImNJFZ9OJlSVxw/I+3kY6+RLS1pB
dxyriSmRctng6jbnxvOG85xgG3IN6m7L0PYI2htRHfKMklNMFjGgXrC233W3TV9QtYRy87Av7IHV
I1CRpwVucAdfo/BnSlxpmG2JkUHZhH+iEvOwhAk6kI8DSMeVeTaGbtIo7Jtp7s6P/f+gf5K4vCiK
U6oNXH3Gxr4ONF1xFIKb49rnc3NRzT5tbWOnn81LHVeVP0QP74JR1VNVAL2+D4q+rL33ZEy6KVnk
+TOU9JiAYauHclZYfHUg0p1YXZ2+l7vM9kko1Nj3FeJT7rvgjO7OICkaMseXoFUbpNOxwl88cK2S
7BK3Tn6DAz/j+/ocqg1wRSMlbBBYYWFKRAvJ1Ip/X/Rivz7VLU9nGJ7Oy+4hIfi/t9PshUs+g6CC
QxUZi4u4PemXfYYxonFFfZTEjps0QurIesSE2G1XnsRy0MMiH7BABdQ9xGoHWwPUlV7t0g5ZePXK
ofdR+sYWqj+qYf3WAQfhMVBD4iJHOJXn+5/EG4moWTHb5HgAnaUGyIvXcNNdCSK5udlXVZJlu5zV
nB30JhwyAWrQ7IvWHna/uW7MBEEiD8meE9yV5wttz1v8iocui4klJmDcCT8gXCr9lHTdQcCIAEiU
263kmJRrObA+Ykv3KZ+ArDo7/r61w3OSJ/p3RwN2snBMq3uyaDt4Pzurp73HXCM2Jj/+SHWxsBop
CLSLDVM+lZ+fPNFE6Ggm37GFNSltKLKqyn+2bHxh2ALAxlhPRrm916zU1LDjIFe1BY/w0mMSSbxK
brKB9fIVriSuOciuZKe6GmtHSFkOxOFgAQRCjJcu5dHogHsImAvirq0HXULTTMsUTO9IWemwL5zJ
POLYUN28emWYqrhw4Mp1B2RaQ1MBedg5gdW0K9Rk0SwrpYzI9QodE8MScH7ETav5AUaXoA+6UVYc
Yn8wo38b3X6VZ7YGAauyKuUf//mQeh9qBrq4K/bBlPs2flX3Cb0KkiTobvOiwc/f7VsRTfyurU3Y
hqKz5YrtwvjLpE/TR1lGyEpEP3d3P5QIkCGCvwhNU9w976cOYSipKpWRpEXrz4NJL5E+wi4cjy0X
c0T1Q+3ucVc416oFvLLhoH3SyPm2eq3YnYKZKpZ6gd19WT3iNI9upn87bjjBuVIlYc3qp8taZx/l
BZhXswt9IIniH59scsabPoVBw1yBw1Vok6ntzB70cT78ZFLmI/4VzcC1l6/PsaYBvB7ynGU0EMQn
wPfrmjB7xUtNkMNrh/yVH2C3NAlnVfmBvaz3HqpO5PIoyBOE9/xnDQJNSu4jksESodLGtOB1AA8L
O0+ltlsNPNXVck1KmkLBMEpItqo3qqLU6DKWmeO8WNmrPGWuJn8bHTgxOrhQZd9r/khx53E3wMwR
uRxiGgK7Jw778tDALD3nXTluXO8cZ9KZAqQUFqGjD9amgCfvq7OxTjq0hGVXOaGwj1LH2weA4JF8
pQAdziEX0qCwHUsepwsSfSje7QkQC1+MjDCX++F6Eib8pB95Txs9tOSJrmFWywNuWY99h9PzzKWm
4ruvmDuTJDeExAcXvR6l5UE0oK3hsSBjwtdBLjg30kxIr89KtIaXrFwJvrqN2hsvR8ZML1Rtqdle
Ckp6w+ykV00Ajwl2KzjS9Cl4DNd5jRkak5qtg1phEALsYthy5m1MGbUnXTzvVpqGrTdfEwSxsAHW
gEebZXVXjh2HvoTUw7cysjq69VFa7W3uvpApgHmbTZZv40MBt+jypEmp3FEGiC+emPoAADgsMbvL
dE5uJoo5Byg9fCB9c2ycXWU2oNyx8t1Wr/wHiMglVkEm+0+22w0P36l9RJNQemsJKcaUPxqI0wri
BThl5ve2d9Q/hkam5/ynLbcJc8VWt7eA0iRKV3wBtlCtUO8u+VEm5YiJuMXOPIHF1Bwc311Kdx7L
uyUpfpA/NL5HWX6IWN1Qa9qUPW9r6ge+9HZaVNTWp1TFZoPriPc8pGzBxOyVIJhp94rL5/f2rwWT
d6uXOXjv6IxNpgWRmuS3sUv4RX5uPZVKLuLqyT0ltFJrYA3KZR8WSBezsfvFmZr56mAoOUIXlat2
UlQid2egylRs/V3GwnMQ/1F06aM0YO2CmOEnzTz1o6echMbpf3gq94sjX2mLm3tbaLXU3STKDNIw
EbmDP0Db3BaTD3YLSzorqX+6iRclVlLOyqkzA64a33myoshjXrR6xj0aEbwEceJNNK6FCTKx0HqA
vasBo0KLJGZeEAii/I95c9zFpISnceUtVPDBCIe/fAP9pnn4iWIcOrBskUPWhz+1zKFSpJ+46Qbk
9dTFErR9uE00Jxgrx70P5QpVTmonSIF26nRD9egN7PvR4ZpWdJjOJJfx7/XlaJ30A3ST6lnEI8Uv
nDoiQBCM9BNUYqmY+Gr92taoBU3fGU4b5qW9O8gjlDBgAu6Tp1fTIa8gTsdyiZVb/gvSbzaPhoc8
d9xIIUnG1x85ObArZBz2Xp3RoECxmsPa6+DRaY+RdwXrDNvcet0psqxNuG24H0DGffb6vS3Ljwtz
yIQdDNGCGeLbgkiwX1QlEMvXmUX2g1sZd2yATjdlbwHiX8J70nzCFh96O+sTdLXMF1E0QjcRvt4O
98RUOlFDfP7F0bZIz0aV1vQItGl/7cNONpakfwDnOca07jPUfxOVvhCdB0alnFycWah/lMxt8LdU
s7VnGHMc/oLFHoiKQwhCCuRsGsi3FARO12yEccseWq1gjA0ESJxjOGjKab2geWRmIC71Hl/mZIIG
j6NROOGqsZMoPpqJELiLlaByeyP4TJZS+WOgI5KbZoa3QcSqCJfJpoV1BoemzN820rWijyHEWI0X
sfsLICWVZJlLiTjFC0x/Ma+uHrISf17QEdHJoshChjAp4OnpnWhYp13OT8EuWQBaQlaOKJxpNtjl
EQNTBeSd91RsAvhUG1wWdWJibe0Nk/D8JIao4yRLY8owlvNzrDZq9jUpVVfi5u5jUEItyQMBXIN0
+8qgRivPIWwlqlfZy0nbLYvXpWozFoAeBB+jUtRQ/Jttzl++l4uY8TKluu8jD9gsaufLFlnVU0D+
rW/x7cbaGvPBMBGc04Q8iGzgCVZo4IVr+goAZcPBLYPrA+xKE4NF08DQyh80b5D1dqIzesrfLdCj
ce2ZVQVYIoHP2gCofME2XV2xs4x+nA0R3BupMu2xayocxEPWaHg3snse9FmoEtdGrR9e9/xYjnKa
/mkB1oJyufOr5QdfOB56q/yAhMQuqahwCLK/9VXOSZU3/o7qpcRZiaMNI+Zbk4+KF4+CpwhnalmA
9IiD2AiBLiBYFBtYvrscMZG6f4EZfCFjLNk1nrX1OkNjkEzsgNXHXboxxlnYw37qHGR5WJE+5Eog
pPGoN8zrJ51lV3bXyTPvE30K3Dpw1kNYnqOdC0g018PT0WeujMlac6xspbHxNWdHFma3jZEAWRur
UJ9EH4/RHT6iooK4dpDoyrud+UPKWeEP4yzeofQE1WnvMHS/etKV95G6ipGHneI7bu5I4bxlZJkS
jHcCY3HB9LBhuPw8kPPJkpf3rZukDqexiOn9dzrsUfh+WdQg8AXRmN+g0jPe8UwSWXETw7DZscXg
rTUJlXH9u6t0pHOSyjKwRf3Y4MKwnglOk/xM6FdqCZePK/CB19YgVoVTSmRiMpsSGSQuwY2Cf/5J
BvkRvZ9qaFxFuffNBUE+qtQuAS+IeMeQ3uph1SEc/+qs6YGSo6yFBbnUCtijxVLK6bMY0X36ZNYO
vhgvJF2Pvn/L1DYSQIFo9stI1FmxPP5LTCd6cw5cmj5wZh2/R1aRvmGSNeTrcXHq9ZqxcDPyI7Ar
Hyl5t2Hf0fKFferfQnYhxywsD5a0ZQfpqc0Aa4SuUbVTv43N0ZQbuQ+089LYx/baOlmS9kJDc+aE
wkGdd0p6PmpJWOlR9ZDywmu0CyRQqVlTjcrLe2QI1RvNM49yLI3IT2GqYng3ltE77t134OaoKBNC
/odLeMDP2Dto7ZSJZgRRC57a9owcQUmIQJBpVTWz+YS5hyPG4Uv+ppP9KeFhQCVodpdN1QEhbNdF
9an+mDI+NyG9v6Y+t/AgiS8KrekqKtij2JYQk3PTHhxcsOKU4HJKCmL+QDgVccmwPhFaVer2WJkL
tWfEtrYhhTndzkDQCkIkA7SMYvdl3nEqzgm8ZfYruSY3J8AI20cgPGoE1XOT34APOSVWxpwkqLui
ai9tKlxp4C60BLsGy+IvDDzq9as+zta1v/xYOnB74qg9UVop0/RK8Wl+m2QasMrGgChWPEOhb4Cz
QlvoFOvZHtKANNfW9k6BnX+qpD8EkRaYjzuVSfAUBI57w8Mfj+ou96n8sVWXaTwt+PFlI07euMHM
/SHkFUO0wuYUNWlgfzZmpc0Z+vgU82kAhk6i94twrGbYEj3RdTcCpxZowat2kIy8+vhTiZ2Tm50v
nuoWP6Nee5WeQcAwe/Q0ZJr6pKiflkeNDmI7dvZrPljpPNr0mezVTkK99uO9cRXSUIvx3d6BXepQ
4J2ARIssFFVy7Qz87mvlIAgVNZ+LwlOB1MtVf10tI83ty38jrXmeo4K4CZDQUHnlVI1zf7yCEtyB
dwiXfFgOkkIkI+cYqxD0k2YGuYcbXCfkFt8pg1fvdQVeu/mHyOZ84fV/Er248C6bO+fnNgVOyRzH
jQJpw6md6bXVfYtKCcxDW/rXJ9qbb4cOC6YVWGtD6D11+sK+O9NF6X6i9yzdTHvqwTpxFIk2N3Ib
4XevwRU4zyxi6UKe6HVSvhXWIR8o+GHByzE7qKienVkf+2wjCtUjVNdKIz4EjhvT4doPvg3ixonp
ssZ2E+QpsRsFU10H2Jz9G6H0bv3Gpq8IwpWYZAofKozntkjtKm0VvkIDVbU8nZP8mG4xZSoXpdnM
2aBcq35em7zkWCRGF/Jvu+f1WGbLkyq+G5D+qAu5Nwf9hxSowQFxxIRzgVWV19HaBs4mfz/cX5L+
6ZO+U2OAaX2QYTh2AfW5ZI5rmNpPvfxMNv1BJ2IvMI2jZUId8y481pTL6JZQ/DeEw0HaExQyL2vc
+uVTsH9aQqLOLonG4G03fW0aHeSp+sENeWmT8umySZtxs2zfS8A9zvC6oi06NmZf8VGVQEt/8r5P
1vgLJKGYR58lX+M+4Rb/bvS2eVv51WgVj50bFGdObTvxG2wa2jWi3iwl9aiwP/0CDda20IKBmPw6
8ZIY0NgK0P/zDFBIMPUfGuhBPh5cpflOBqyIvDuYv+Ll+rHZ6JdWWY6FdxT4mMHwNEMAb3EFO5KW
NW5uzrVW6QourLRMUuN8iokeyHR0uIUKqnDExrggk1CeXtYu//AXIFO2BKtoB6ZJNK6HGhd90MD8
TGpj3hUC0bMLTUsQJ20Mro8IeLHN/kfOEpkedFrMHz3aR5AY/rbJjC5aN8ZBueOO1diCzErcKVyO
Qk0y7Sj7na8qrvmsVTMowB8kCljwCw42QYaQ8s9pLzGZNZvHkf4BA50ASHxz6EnrOo/obTUGrgeE
wAjYDIbZ9yU6o0+VTXimQBSMAMpZj5vUIBP8tGnMTkPb5zRgAGEiibcUnmWL/s7amLrvEmUruhb/
YnxLnj5jsO5W9Q/e783hK3nJddaYy7eOfntG3GIAScBLEgT94rtMo4M0KHJyYmmAUOBCO4vXjJut
uk8BB9YRcalDIQQ474JwaGe4YySVU9O72tAATo3tQm5of9NOKkOyhHaJue2UF7TXj02zCqq4cZnj
CgumVjTVpA4iSa6/FsQuADk/OEVfPoyfMadQgFCe+gwLaNxUya3ebBFbDJnbJOYZ8o5wxlzUJ5Cq
DTiFZeZ5EOqAO1YLJVyZ6VfuXhMzTmDt/TGvdaDnjloH+YeYNdesoveSTCvCOVbBik/WE8WfT6+/
0qiJrprVkoodfkFAEr6pRWIXyhNIN9HFQDcl/LJRVDi4Phn/58Rc4zCPF1Zdr6trc0EnLAlbUANT
3ICSqwOMXwQc2Wkk3vdYPwWnrZhdqYemm8UpjfWPiwUypF6ALWKyXR+gCAqJbStji87voddaplRD
gh/5e/v/yDJR0jPMLcD8zoWNNguo+9xzc9Mj77R/l/QqQwuh9Bigxv18ixupOAPocM5Lb0eSdtoI
Ymmz1WvMktI7n4q2ieiiMZ2t14HzluF4TwLhSqwemRr5Gi5qbmfMEn1K7tZWGcDheysS0O/mficW
h3ssRzJQSdSbjX56Iz9l62f9KPtseZQClxqlTK9oFo4oox3r8H+DCWiKPdCrzJiqwc+NVjxFKDMz
1l41qgNZ4CHs15EhJzPzR5uK7/6D6Y79/bl+fOgr7SJdLaNtPch4IFQ4sya1nD1WDQfOEsLGQIH1
YZ2slABftBkzrJ6rKCqelTt8yRWaCSvbCA9ks0W797u7G1WfoUureIwyQXWJLbqgWdQ8tm7BPAgl
iaVxVf7rqiFYYUfwLY1AaCqCKPvMAySOyDYFPZ8uPVI0bQjRk5CIMGslPZ74PKtJ+ZozX/QbgvJg
ChVLmOc/piOu25zuM0usFy94wcgbRB+R2Ep+g+fne7ry4DKLLnDUvKczflzTuZyBNdU6G+vNAceX
Te9XAdDcjfD6PKYdiPpQ/wdWrwq71MeKsf/C8hmzU7lgI8HDmMA7IDEAS0xWkT2QaA+eH8Zempn3
hX5FxGihX+/8Cjkd5EJdIol+mF2Z9RN0lYZ+qgQVsBEMWgi/HAeM5M8ZOoBaGhkqkrpb21gTOZ4j
gRZ/YMWr/+h2Oo+gKHaU96r48ryDAnyWPBbSVeB50+r0hljjEyNwKz6esPltg7URZ+PnKI1a8f4J
7qYImFUufnP9smH5oC8E7xlD5w4l0xJLcuGfJRfHONB+3n2RuB1/TSZzFAEOEwj7BdSTON/l5HUH
9Tta2746yfFFOdRDQOUSWp/JPrc8SBeq46NYSILYB9iHCS/i4zryrDEne1TdO8FNKKpUnIsJSp6M
J831npwZ6ji8/5mgdNKps6ZjWvWLIEHBpLAn04kdsB5H/yEUHz/BLnq48C/nUz4iC5DGdBCM9tlx
K6InVB6i3wku12FxlbDuLzGICTWFGgkDYZV4cwygjr2Htm1/v/JPOhGR35x4uKw27spXl+Hecx7l
pjHAUQ/71EFqU0kI6nPd+WK4gmbN326ixzSWXy6DZtuwgXveiN8SDA1WL8gJbYxlO8QmmbDYVCbq
2+glhbZDZ2cpYoacH009eutRF8wSw4WpG/7w2r+CMQuNz2TsndnlApZAnH2lE4NSaIKiRch8UD32
+HjfDkiy4XGfURyeKTKZCqCH34QsfNEe226vyAagkwWliBpEnlUzN9yedTlrh2LbefXTXTmykwza
f4Q8WxBH+ygQZD43f8X4ln+JcWhcUh4l87j40kQG3r36z00s4eLnF8r8+WjCeFNtsM5wfXSYSMK/
WVBcFEqZwz0j/7vZTFJSkCu+T/1p7lFr3iTbC/bKhcy9vBTj8z0YkYsz3wfC9/WwnqKfa6jwpoGE
TKVaUfMi+fEdGJA9nKXCG/r2u8o4JpialPBzRElmH/3ctZAFxJ3fIpKtnPcTE39E9UrQEJY3Fkus
V5WvjTB3ttF+OZp1nHbqgMtpPEmZwPWRzrHXMV61hwnBb8Z1qgQDEVbYBVHyUxEdd3gZjHJqzz8X
VtkHYa2VVF6PbmiZfktqnioo8CjXUJf5za9sgeVeMP14mtThOwfAG2PPefIT+kqJjYik3oUP8x6v
2ijdQcZueVPP8NHKE/PiOerUeQGbl/FIat0G1yhjUnBTYtSdWhI4/6FcBnAI5idcnhF6Qoyrq9a+
y8fBi3Lr6EkEcoVeJ2rfmi73zmADov2qUpYmxAs5eBjhrG7untFaDJo4LSkgtHzxWI8JqTlmNnau
qQNYfxI8+yH0REwUsHiYONlYbCQoXi4fo8tmsPaIxL4804Q162fuNgF1ax4qEFmihiGYIS1eC2xU
P7F2fvNmaD9pyiMSuVlRbm6v9R3hqPxgxwijTByq+/eFehW4pTDV0Qi24Kv21R/sLCWB4oCCdL8Q
tNUbdaoS/qcHvPNcRso3J3ZsHEsDsqJynFsQz+FyOsPYMwQ4Lrxq0mjbkmR+JtcKHfwmekueFASs
OchIaY7pDrFiu/pNgdL8T181H3En3T8zOArwDQRMhvGbUNkjLbd+C2f3ipDPKF4UDbz9P4TdmPQc
oHAnbJXJqaiTgkEAWsvVDYQoiinWhp6zAB0DiAjpterOQW2leyQuI980mXov0IUafWp+RmT0h4cb
AvS4De8Xxa7Ru3HG2WIFDeETNS8IYNOYayDE5yYGi5q1gkqKmjmJpsgA/OV21oPC6XMPqS9Bu0pO
Fnbsl6vRu2OBcWN/yVE3+PClU1WP2jfGyH3OTKTNC4dS7HrDGCDSdGL+Ch8fAV2TXv9AyhjUAQPn
7H/pug1P8NIv8k9lxlw7Z1Udzodf7NjmKw5tpFehE4qs/jZRmeD3bSDlD+Dko1JgUtX2QslwA5Zu
A3yE+YhOTIYKTMsc02NktdnnWvxGYj1iaCINKSALhthcPGTCw1/VBNWfQnAkM0uCyMGjzRSBtoEa
zxkFP3e8lX/5pKSNndLsmpJDEkNuPinp7rC+g5JWSdt6Su3k+gSK5O35v769Yw9kLOF4MXj/kqrE
CqxTa5Be2TI+Jf09pht7xjdt6cUTd9GKCnS1pK/MhmNcomS35dE32PAKqjQLPHAA35nYxU2uM7A0
K2WER6acbLrkPjz3jVnKoa3mRn5jqAMDyEjubS0NlCT7lWgWutFkM4cPm/3OC/B5rWk6ngr0eD73
a09uEdJOzECr0qe7rSXWNPnVWR/QaDGo1jtVx2jtKbOfDj5tQioziSxw86EsueKlhtQjiKvQ/U9u
EXFFQjRXxCT5zRettNmjMjYi4xCs55++PpCIcpiaeI6hhTu2SoyeRpIUxp1Wqld65c2tExjjTOBA
cYGnzproE5fyN1Z5CtRqa1qygKCP3mThQ/wlGryq3bzZ1dxhUcuDEqWLDHGU6kNf7vcVvNCkCKoj
qAvEvmDi3RzKXYW3OW3kW3b/oDS+xJUGqdjuWdCTM1x0FVaerjdtGxfxtbfloxNqVmTmrmvw7l91
c3YbX3WOUkDbjgM+wuCDOCLiSufPN7sJn1Y+FLt6qp/NROd+8OC4QJWg966tQliy+Cqg/oIlCs0H
qDqcTX9Bv+6aHWC+s55xiCGUJmGi6jPGAjLOKGWmVqlKZ5nR7fkuijzLl5mIjuyZEJK9AHVXbvMM
WRH1pfgIUcCPJfQS44vtVHtboO1Uf9D6GpqKAp2zVNEcRrKRIz3Yd5fscZRV1fjVq9FnCX0btCmQ
4vgdVSiv2ibsbsqdBildn5rXZU2XkOFQwMHVQdRa6d3ZZNGtkVz47GJPK5FkP5DY0L3+aBo8E15k
BrVDlsjyFacQG/Lldlfv3GMCIsZKwhgUeS3Z7/UtrQPVBoz/D1nRHpBP4is3DWDdF48QdtAxuGxm
j5lO6W/FYt1PQ5MTkiNBPSypPG2PucAPjx/0fC5iYqRzrMxY8pnDxV8Lxj7uh69c0St57losMFEF
xkv0lqx+HmnjCLOexbjRfOKVAUMKBa8eIZnlh7xCGGcdXkGUMkYYDBc1l1vn4ybB6zhiCHuR+SFA
ihv4V0FpPdMVHx0Zceog6IsbSvYdPDJOHQj8Saa0A3Or4VUz3+RBMz+skG4RzrkdTmn8jMqnyY2X
PY4iwVhQBHm1P/MlHZxmLVo4CVBnfoEw63ml1rrMnh1YzAOAT7lPQLI5ZUhYg/pbm0WDdx/Ys986
apJvCdDVz63Vh2WEO+xUKIGLQXLjhq66GvyT+YQj/2GZlqwoqEDHAQKzoJuMK0um/Z5IPpdeOaZP
IbAn/Pbw9rSkm4NpXyzO4A3sxHqo3OE29pGUvcMzmUSJj0a8AaIM0AyfLcrNcXKeKDcohECyaBvJ
+EXINQPV1rb6V4JmDcXGtueNEyIwLsS3bFfOIyvX/GNOG/nHqgBE1vHRCHD2QZV+qJUJkQQCrF07
jEmrm9yYQd37RpY/AZk1dmxTM125oPpPuQk08YVjX2UNYZJK2GCBpNHpO3L2G5k4IAo4ZjGVinN9
s2BUGZG6pGvLFJqVYk3378PoHSovEdt2zI4WPBXWgLCGTTLT/Xsu4mDExmtaDZX95sPabiJaElHP
x17eiEAPvRFi3jY41+woh5vnQTSL5XDMH55VMIaiGCOxZ8MD2CKuHwBBWYdbgVBvcRIt5PRr+HkL
0Nyj8vmaRoasqIInMWz86opAMYxvO+SGXARCrmH8KxTCiHKNG9wY49jtYancGQPQKzzMl8zf3cbf
Fn/6EV6N8BD0eRTy/WHMVeOiDevCHQ40k7Hv+TQ9KryQnf6AJDEv0mj6Ex87YbfidE9C4Kem1v3B
F5htqEWj0P6ZuyIJwB/UkorRpN1Goy8Gr6lx4wgR3pH0KsYQJ7GRMsOVU5CS0HNoqVVlTiVIOFYd
W2U2bEaU2nFiin/byG8hgfHMkZ72WMkHSaLX+UTXrQ3tVQRO4hV0WJzDKDuBE0ggzYB0Dj4VxXuM
A4/q6T63ZvQItWMLQUzPSUOeJwydNYMH6bcDjPAOLaTGnmksj6rulhHCXSi9yp7U+RxM4HcFUtkX
Vne2RsnsN0byw5uNvck8TaAXPdl/d2KMQ4fuscFsB06PtkHSNLPm0qmLTGR1rfG0qzQoQAjeEiCV
dYgE7fZ2VdOb6rEmTCIRUT3lM6MwAKIZzltzlY8otWrVhVxO8GlfJJ1EVJi+HCGxZRyJ31K81tzt
9hKryeCsEvoaANRUEU5nb1SJdrM0NUwO+SKCN0cUExL9waRgvI3y3VJPbCuz0B6sRqDRHbPsSWVA
/A68ehweuHis/KxzQPb38h3Xp6ytrhpoe2SP5ktdPV4gXCoefAXgu7SmYc2fFJ9+eeF8EJICu7AN
bwdCrzm3pAvlsxias3YWSuDekvQtljDch8wLWNGKb2a4FVfsD59faRKtHp+0YHGoct8PYgt9nsYi
coNWTg3xoxLorITNt+0tXaylQWLRKp/Y/To+J2HeqGOoCS81RLZzUPMmv8SEDMd6Et5Fbo5er6b0
6FJbJbNeb3bYLZlGoGT4KnHUAgNzan7qpSUIQ06W86ZC5Ecr5+VLU9Oa9yKdWa+HQ4VZ81RfFMPC
xf1jliRQX2VQDzIUYaRCdckJRswXrXY+BhSlonPRSa69ZvkGN0FbvijPJxjE7T047XPrm+R4b33t
p5bDxj/7Azt+X3RUNBgTXkUlBiyYZjhVKRfwnfPHkFusvZ4jBiMthf5irKDm+iNd+ksZVP22E/uh
PqIMzJEtnNt5kT54o5LG3CjZ5Aji7UccX2mHng0q/tE6/o/MBygNtRv2QdFrskQ/EH7SnepAibzy
bamP7zHYGJhmnCkf5IEf2V3OUwGEC9ziHNi0Fyv0yvTkoK839ZXdPHya3vfEkK7SdQiVhRrCUpHA
1H4ORw4GEJeinM+EauoPUcmyz4W1GNrRIqm/uJ7yeT/iCry+VRZd2q5hHELMHfJduavXgYk8ybsC
JWQ0FcnksExhBAZ0Nt3Vk/e5nFjwBkxJLqTY5pBU39Af+1CRTqymgih0GmiVILTOHJoF2aTo+qTd
fq/oCculcEQO/JBoHgQgoIaRumpUqZPpqX+bSbo91BS7OQEk1lSodKdkHY9Uk4LuQ0VtgY+KIsHU
n8DB10zVbLX+5HsgBosOJi86KaGWr4hTmZ7uOuF+mH5F0u4YG+fSDj7PodobAxydUyiLcK490TAQ
evvJTaTSjpcCwtDijhpC8SQ6pqioqUIDeuoQH8VEaQ7Q79Ga5IVugi61t6lA7cGuzPlIQ+59Mqc6
jEvTptqRgX/n/ZmBy/+XKADzhyhTRWgZRtI8wZZ0R7pgbemlfxK1RR7pAcECETQJ9Pr6QWHDmw1b
6FCAcEpklXaYDdwKqdLl4rXnRtbh6Qy/6tkkN4A/15paZIwzg5lLzQXCvsuJaAvl/EnjAknxpyyv
Cn72aoLGC3q/p4UFI37u0NF9KfcD6rWG6JAanvdWJrY/Whg6ACelHkc/ZTob5a/U78CcxKxgwfyX
UqE1pNC0gNrMd5NwmjvjjFKtfWwqnZY24l/GmyaZKyuy9FoJwd9pPpYe03oGYUcCDQJm31zoL3Vb
0Jk+LY8q6ZTgKmrbP0d/MXD70YXI1Dvku1p/Oy3z+i0qTg1KPZO5rYHJ5AgCZmrR83tD6solnOjf
R/efe/pYK7u4MeRwUTobiDMLKFc42H4N679R93kYFmYr5+qJdV0/3m502hPUFVxJjw9zSjFMwhMI
KckzBu72MwW0MqntDJX8iSUp81bEQSXkOsaHqsJpP0e9kW5xe2/nxkSsit72ZlcFg2FU5hytckgi
7IR0HLV/Znwrjmz2O4We+p50XE/CG1oJlNHXWeCnuklzkFOf4D93PRJbKSZLTKPwm/XBoqCa2Hpg
pHWHIHdTIc4TcxMBAokyJNZHMWeokNVBtVbyja+3bchqIPvm/WGDyTbFWzrYoPV59gxGQvkoW81Q
4Yt7vsXajW2JZ4wC0fVAaf0J/TTuPDYDRZ2DYQl/aDtv94CAUck7Yh6OAn2PFeZAzyDHyL8Q3cK7
tCBhZ0oh7XdoF/zpyMSMFVnglB+bM27ZYT4q5zdu6x1DEcOow33QyC5qAfTk8HGYO1w84dW+p166
nr4yBoHPXTTU39GETl3/wT0aSRcw15A0L+6p+QiwLyEviUyS1wh4R2/QMd0c4TXCCmyN1woVNTPh
sSBqTj/fWyDSTB3EC22UahQCH2Xutj1KGFcvRsB5zUXdTP5KIv0CXGBidAlcensr30KPr2U1lKwJ
mfjyRzaGaHoqKfTQBLln59vv0YgJD721zCJR6WrtJi3I0FiMAbulCeHv9fpcT4snt2PNWOV1lDOT
tbcFZe+1pguedbK53nu7jdIeAG6aslt+GqKTnBHtrk5EZ5/nMhhQfqmlPAqtFsuK3YFEPCj/FEt0
p47wL2iLHOCZmwpxDG9b6Z4Y+XSkeTHrrDyKx/OCIf/jzVY5I5yvkP/aKjqc6nG+QcUezJEiyP33
C4yvJbygN6keDNkJvl6R98lWk2WvGO3nI5KO2k30CF3GKT3o14fDqXNB+kbu1sveq7XN735dHFTz
rLZlreA8Ta7HjzTpcH9Q9IS4GYN/JBiQIrycBMBqvhPblPeh3wdDJhNVgJqXhQLws548nbIcM1zW
wbaa3Q+X6ostAN3CtyHXNLnBGv5pwCXqW5M9KEbzeJ9+L+mC18db8XBkVWIUpXNG78O8fhKgyScn
Z8b8Pq6/FXJwXQExWj3jSvL5+h/lA9pyvquPEb3Vzk7kwtpFixFCZwkzkGZEQdcvXLaprA7sD64C
2NaoHfioxbky7DGpkG4L1w97SdNsv0+g/GcCrKlJrSguk7qZOe7xAhu5PJpZACDEqcKBJkDsIdFK
8/VWDNPoD6C+kTUDtK8wMFndWoYDQWhqgYMKz9wZJRPcL6KMAam2snD6SU6cnjTBji3jbi8mZVx6
6rhXyIrS1NvnykZ3L6yR+hndyiyffq6wbuAZFb6POg7CdgbOmerERSXWPTC8wmKUuY6xkWO6KVu9
nD17I1ZKeQnWadvhRly1tfUVMRupeUGOyTrCcKg0RcuK/KhZBN7WDvr9wiArH8AMj1/Q/mJeINCw
7uUEkDFAPmy9a3rgtg3VuZNI5OWTwtslif8sMrUpmuM0d3CzclGo8YbX0O15/6NPR0rM3toDHY+E
p0/Y08XKEUbJhpJH+rGF3g6aBljPanAwaubPxQnBni3AshNvWWDz8CvEuv9M+HyRIcazIEhv6w1O
hqziLeFHOAMUxAop8VqU+JJv5MDPezPB1aCbdLnBktva3uMumQHxyMcNXML8wRi3LrVqgQumANWA
i1754YqfQ5r4C4DrZusne1NR6UBGqzb7AOx6172DYnTT0IE5o6obwkst5A2SB13EWZfChxALvlRa
I4pbsDUtl9L1UHRMLxP8ThHeenNZsQ04EISbM9NbldkiYgKyn8SLNaSWyqC7UZnSjZMsqYBvT+u3
j5lDBqDnEntrre6/Qo+o+qeXEoul4z6P/REXE2Yadr1xNVieTkG2IH+JGj8kanNn00fW7hNy7Tdr
fFA1GR9hXvRnQtsJtSD+GJ61evD6YqB2c+rGC98WAg82lVvJZqdpB0heR0qcDGvxCI/YIRvyj88/
rupv8uq4oWPv0CzbtzS9JKJ5xMu5b6rcD2ZB4sjbOvDCywEyE2KQJ+0G4mm+ktLM24mdwjJjKmSD
vwbg2aN+zazmh06YYutjBvjykpH200NlzrSor8uUxAjNIO0/1bOKnl9WS9rebkqb+nYJ4J9RcGnS
Sa3GpZiiAaWUk+C6tru0eheAI/gitZpxWgPdFfptlosUQbgB+E+C1NwmFFvx1o4jgmqndT8VillG
6meotB8ehQBiKywYCi/ZcDLZkG9THAXzo8lpbT9aQSxXr2G10vsb7XidD6DYNvCNFy2WwgzsFV2Y
IDaVP/Eir4b4/s5mIP4f1v+nX+i+czzIv6AppfPD/I6Sq27bDriVwpO5TP10obH2gCIqGU8lFSMX
ScKnATbzNB1JM/sFKbZs9ouDnkGZ6S72VOeIUVN8awKAR7EEn8dOhCcXKGa/XZItz0XzIGv8PVCT
fJXNj8pMK6Rga7xtXGDf/iB2sdk6KGCNpZeGOzf6NtB/cOWKbtmXkDCpnYg0I16Z8WoUnNMhWTgF
DbDej9jsyKffOu+9rqGTCbD795aibvq+qpO7m4Dor3+d24Yy3/GZ8fNyZKfR5XdUG7Ex+TxfwCqe
ZpvdmVMzPXF7JRhKCa0LtIGkoTvdE3KysEdAglTNB6YoJgwwtXcRyitKDZVbc/BlcQ5W82hholK0
GBpwGvr81l8NtNLk+C+z9AOzlu9T7h+IhIhQjzjwhQSJ3Qr1WlXTQHRMgL8pz5uN3HaLN8/lU4VU
LfOq9LjZgAvs8I2e+pIxKBa2M6z+btAhW349uK2gGhunAAu+E4lhSd29TE8SFxfWnAJZAQliqUJs
6OggoYeOOal70r+q/UriQUm7FoH5K6wDD7FRWXug245i1j92wyoJZwYLKBH3qhIeLYC+0j7q09eF
9TWg0ExnqNaz10KLNuT3fdyyaLg9F62idgzmd8pErkCJy2PdQasJDw3FWkcA7hql6EJKtiXab3Qh
14+C0TBxiMjIXgwrgNgqPckwXN0YQzvKIUIPyef6GMYFqeQgSIWmKLPrs8n0hrU9js1WLU+EzGWo
iqNiqN1lkPaVxTMTuaeF/LSwCMsMPSTxPxBbKW1hslzct0OoWO43J4FsB68quehXB2BYudDNq7FX
Fs22zN2HcRMzDmXiganqIIyXS6yLytO562MRGjhGh6iTtojcY1bQTzs0oPpl/i1rj0GPmdZnq48W
bGq79BmVaTBiqUtMyet3WM1eRLtpONLPjjgKkIu8HU7FYI8Ef59W5VgYfXA9WDtLithfmLGoARqx
xioQwfwR5840DO6/IOKWAJHispZRiyKn2W8rSslY1Vx0QNEgNNlwKiOKyJlnSsIK/1K7ayE7Puow
jw9zUvKrH/jXMJhJPMoOKco5J4y5WMMeL8LbyRYgnhhTk/DWMXdZ96Vf+rO5tQtEV+9/d6aqD/zG
Na+EbmD2mgFatsOjlFCmO6fcUXMfWBcAu6ER/kuPbDWZIXIlAv/TYQceL1kf8mRF8fYvWSW9+br/
UqUH3FhQd32cQDCLkSdlFE3TAxiFDsqT5H7NvpYMZtwn1rCL9JLDkhsaoqlYCvKPY5nMygRpQ7ew
y34lKgCNJZy4me0UjUtGL4NnpOov8OmPxHkSbejI5R+AvUgGiWeWNXUqfPAZVQEHE1STMxafD4s6
KHr3kRmeZLOOnPW+voELF04+kKRl7SfYfcYXnILPN5Cg/eH4HEDLplkPwKULqAAfWWiyi0INCJx3
17OQa8pB98JfyzUgoAp4IkXi898ZLJBst9UA4SgA+8/TFifJOECz/qOmYQ/dTj0hsTVDuW/GzM7p
zqZn+qKM7qfr1+jDgT3XKhu7wm6khzY/gDYtjPsxImu7fyrX/8SqZ9WExF1wZ/DWwzdKVBBaWcFo
QLbAeKZOawnkkmv9YNvKFn+9RpF9u1VSiK5yE57sr4r1OP8sUHLSNX74eSCZN43EQcdMuai8X3iG
GwkRue6nnOaT4JMFWDbjYG+K2d8YPUfS0EQ7Kl2/uZEZw5tzO7VKeeyyFGJeFxXHvUe8+7741CgC
MwRXQ41XMvRm3Unjrt1n2M7pKZInu2RQ9qOU/OjtWJ4mnBye5/IT/ZqwoXPQbbCESByA3N+ICA5x
p8IR2JRNlo1IHrLIFzGORsdc1ugdnyTRCRVUVVsRmaxCGUGq6Ps6Oo9r/3vsOkfJoPRH2Ujj++Xi
gwhgc0bxz8DAW/3h/WuWkUs3d4E/nJAmWrnbxqqqFaIV0kzsxuh0GRDwXDYbo0bn+sEHw6V/+gEh
5pp5IAYTlb8S1lZkO/NGWMvoKRtutqzv2QuW9mwci3Mz060xaUz7euCYgS7EHNyLxoSbIAJnq3uz
pkQY+dFf80LTKlDu3WWDbKllaC19kIhWLRfR0RJEZB3YmJAIhiNp+gQ89SfhaFEaVFfCn4dF26pK
IMPm0mVlUDE6WF9j75lyZdyLYh4YY4rKCrXDQd26a8aqS5yrgmprl/xTBaZ+dF/bcqjNh1CYQz4Z
upcWEl02qPpG1qw5OZJR5Q4JAwykmy4ogS/N8IVFQWhR4rAFewW0sDxDJ73noxuoOJ32e9Ju77l6
o/noocFIoply2crvpSQuPEZ69UhMUBh1dVrVStM8unqB2sA3sipAfQhWb+CKw8PSD6UEs5scG4jr
ClhwmqlErDc4SavzSjpO1G86fcSgdHS+V7wawyg4AgA59l7MfeKWInTFjxRZMA01sCP7RrIKwt9H
NS0R1Osh+rjMqFwjcDBcAf1NBHSoYG70IG9xNtxdiM1s9fXNN9s+f9SbGIWqCE0wWFydB2Jb1gwP
I7m9Ld7I+fql70v1zMTI+ceG5QfWFKgDdPchKo10X3NWPEpI9OU4ykPXS/kyzZn/MoRHUmV0Ifrn
hIj3ddHJwGYcn56A1U7DnCdsPWVT4ZOAXG7ACPQANznbCFLPiFEKxfCFHHKnRPe2E+pESXBsTi6b
2+vMmjq6nT6u02czeBh6wo73fX0sqimPDkEieIR665ntsSG+crjKKNrvQjvn0TREmasZm5DE/7vN
r1oRiH1TGG9WCb24YUu00pQeTNqnBEmMdRUzY6/fYCXgrbVgVMDIMb1ZlPJgylzOOUaqacVloV0D
crp+NehS1jm7bdYY2N4Fj1lTzUqTlukwamj53Gy/l10ckOrCdbL6cjON4juNs69meDHxSJ0f5u6E
A+0W9K9cYxwhQ7sO4akwCjJqF7GONs0SJh1nVOVJDR+/+7Fxx656gIPof6H6NYR5BUjMZ60ROF3d
ItCxC6Wi/4onTS83aRGouWIwzlA8SL1LSju6wDxx2px/YdrNa2llICYeIkhuCioqLBYUc9TOiHpE
kyzLP4KI4hpCPHKc0NvQ7th9J0Rnbc2gVX36R6zSfuDWus5bU1Zd7wSoKeF2NyR2hJLTcqP3OD2o
v6jsSahv4xM6D9MOwE1qohWtofJ1S3nWgtNOyqPp9s6zC0psJ3rh7lYeXrwKXMJmGxxmg+2huaX4
7NN3/XR4p0mVNAflEjkXr7biLNp9l/QXvAg9xQ05st2LZfbdmHiKIa6UysnCf8b5f4Lr69bJEexO
4Vsdv/vkCxO8vR8PFsdjNX6vo1vmqZiv/JkEYcXCyBQ1R+Pdto3KNgczKfc5OTeJCW7k24FvK6Qi
qgr4xlAX/kPA1bCu+ru2CJwIzNipjIJUkNBxeitB34cG1NL3oYuMAzWq879w6dM2/rV7vmsgMZKS
tjbwL7DxEE51oi1WRtCd736zJB9WQXvpjKqN5qnazzd6ir/ntZL9AQhERkbIIAdoYLicsw0Km0L+
J8YdPedy/2v2cOMC4Eh4kj+YBwauX2S008Jko2+ek/dRVKfn8t1X/goYUWHoI8HFmDO34dDLTv6k
CuV4zwU1XyDJvT+E472oy5m8rtGOk3EoXAZm9gyRIkn4eLKhOlveobZwwdvO6Gh+IGQuJhXbwRfA
Ous+PBfOk9vMwobKrCeoOhx9QwUb4O95gvtXg6k2I/J5oLtyWyBHr9wDxSfy66QVIv9iutQQckYN
seo7mq5EwrmGPLV7cMljZUGrkcaN9TT7WUofMuIO4JRwHADIZY/7Ay8uR0MkIxMMUF/btNoz7FaR
DEEE9eV5ZaayKKFEpcDmbSK8x522Y2p7wwl0I+dv7Uov9/WmUs1T3gGgMSUyLvxaD3Vojnve99NY
nzKevx5WJLH+/m0gQIMvXRIbW2w6fyd3obHyt6gmhPGLxv5J4wdobCATB/Hx5tEPof/RjIqzYl6S
IrDuct7K7MkboFu4C834BTDvfejeqBZhRk0tBKFmraMy9+5nS2ZPbQvFzHg/7JWYHkQIqLspNTV+
I5hD4NVuz49O/Xfi1XIEdh2f1Z8qQPiLImvOkdV3wVLfKLhoYZbnZZLADnolMKyLA67k+LhbJ3C4
oKIqkVrT5Y3L6WAuow4wuUIwcbRBIhmgHaB4u7BCE+g8JwYEEI26Wbkf4MYdnxDtR1CRV7wP2PTF
o5jyKmPJHEBxdBksfPtOiPRFegfOeiA37jUDdxfssORJTemzd5eCtktxhNVXE1T6C4mQwuhMZZu3
yeHZkhgNYTS53rwtMgm3i3qCA6zVAIQ1Ru792t/OLVFJuwNDEZ76ZSeGtnA7vJ5IYWqpFZ7YbY6O
gUY7OCiZKuR4IuPU2audHclXfaaik6oOCRV+qC+0pX7BVepj2znMNi8Xrf1XBj62ITTFiqE6abr9
kG9IXjjVRoCSchVK6NTn7ATEqpq0XTKTev0+ZA13YwV/K1AkaOLU7GbKfnF/mjDb4kv9ltLgdW42
ReIceW+x4djcWk9RgY051XErxkvF5YNAolcBGRIh67pwliDBeGubIo5NRHnZvxl/PPdNuGD+4wer
di6RIX5L/miXf2bXDVO5iuPsZkEIrfDodYduxD+aeyx9C61VBVa5IrCkPhCNKLOzpQzAcCbRwMM6
j34+Qhfdv8QOBqKfmHBJRTN8vp4qpeTM3OX62OOvFNVo3IWkGsD6TLrHiUeY8npCPbfIJJwqdiyP
aJ2vI2stz9M6ddZefGyaEVia5ZByGniRkKVlGai6vEi08uiSOvL9rMikSFFjos5DF6vgZ864MjYv
EBDnLzIQi/HHzBuV0kmO9mI49pG0jSVbJQ0ymS6ILnyw+4MXxqDzWfLtOzAEAvDKC4yU08ebYzev
ECWNCiTQDidOlneIx/nDJvv8tpYqDtb7+OUvmpkF27Jj6y8+UmSJs2NrXgF8aXSNz1lEdRchvgFQ
TOS04rwZaBslKCSLMF2vIB1C+FNtdKNN7GYdkQhcjwkU+p1iifjcxms/eQRYbtrane1dRDuMk/yC
dOwEXE5Fn1Yx1N+dUBi8XNE9IKNJMj6ovdjDPu/Hi+heaDJjyp2AnYWiJd9cv4vCfSKO3x5p7xWO
GStTlUwc3NK1PMs97cWKKpfyh3KsBP2dMyVoqamfpy5JbtPryZ8UrWlGnQlCsUCgbSHt11meiYst
Qn8ErdAEl7eFrBW+jAACL5k7vBsYV79Cw/kWqpOVGRA8tQNCD6cVSxmR7IEVW8kBZwTABG0PbOzc
nM2gvDVGUDSTi0+zWwECQBvlZIqkq1oGMIhT2a5EQTU/IzRH6Zin9irZu2v/GGheywzMLdEJ+x5F
VqU0nFqHYPBiou67BjXVhv2GCgnko8+AwDHDmAoINH/bzhcDckVeJyVHlVY8Jc2wJD2JCN84p5wC
hj85GzPR6ujrHMcK/e6QyflbF0h9tzXUgPh5bsCgSckIjcl7GS8X4TFhSovKbKmpTbZppZzgFbk8
SAgxfUriyLUE+SthDhUhAJqGnu9JtYWU5ThGn8OSmpILqqxKoZyxU8Vbbx1yOlaVFBxajslC0tCF
Bg4PmiFt2h9Kvv9K9uUDXoDljHceuUemdbymFSYiR1H4QUJbC49vamDaTCTXNHImnCx/qEgw6fQu
0y5TepwtTeHMckheHiYfGwJMCZmbxXVNd/onAQCuFanIPbTKepySMIqyCugDil/fNv1mHiZjqwcM
BH0hHf+RIV7vmiDUXuC12SdzvtQCGZCdNJiLCHXu3e6e4QfDuSe7YxAwZCuOfdhxTWPwp9iq/G5y
N6s23g20Kmnuid9odlsEGBuDUaZ5EnkUV4CgfF6veASZKEkuF474Qz9OZ2XCQ1UJeh6lS9klbH7z
J9CCTB+ayPTr8kw3/0ejgPRfMzRcSCcSwWTbkbIXiKkcjNolSsB+Q0iYW3KxZTvWJqpGIWMYpFQ1
egNwF+jNBPGhiQaxXitWrb9ez7/INiVyN2euxZjiKYAD1ToTGmjlSp3gepdvBgaIPTbK8awTeMNb
FtSnPkObfDxHhe0+XAjTTgbQ0y1kKoOp39epVSINQxER3258YVtrPJ52BzNgJZXGpY7g9ChGGm/J
PN9TJiIE5QmejhYWcdyJ8oBQmBwRsoy7yIwUX6Wx0qZ2WdIoTH6ve3FHUFIoLkq2w5LHFR0IT1bh
iDZQNyfd2xN9duHeRLB3ImwgiEWv88EG14IWrcCSARt+XPNbeaVZ6cBk7INUDl96szftJjrpHGH8
/m6DtCiQZcQ66JAWLogd3v5rrXEbRh2u//R13HNnb9KHcnHsJcmX4U6HhvQ7TnBaVmmuRpm0Yctc
qnDj3jfbBmVjRTh9J6xgp2F+b9rivBjfc4BEAIhIejmN1YdmdmMBxv2ReRYDQpQKvHXou+HoOBD/
W5y8nramtA48PTd4PxWyvyE6tDQUXYUy1AqrnhAeIsMKXgL3ZLDK5PUUaVZL12vG9z7OkdAVbsKF
xrgf6DDwChm7KZehqo7BNE3tYvU2Usn1MdtH9Jh4el/QrmzHnmYbKnNYLdYN5sav4lZDgWPMKLpM
cviAls4QIpXCxXa5unoRocYrZ9g36/wBeq9zRm2b9X2+mhEIwqwAHRf+Pn8J3S1ZRUJC9EFPbbAg
XB9qmQ6xzy6v6OkG2RsKBGcqJL3Ig7fUNk6+xpErb+6jhx27H3fPAxAf7TVlRdNykHDocszfzjW7
0/CvZjTrD45EOsc585Xl2p/U8p/Abpx3UW+UnGlnmzAFAUFzua51Jvatkkq73xY3Bouh8bvnudFU
0VJa2M4K3IWWfWWqm984N1v3AycILI6Cn38dnnXy7A7UYywwsIO54erfqd6Uez6JZMx2od2XqJ6G
kGWVNmyzlg8bgGu+Xsp2S+LyWzxsFzVLB0Szu3nAp5Ur2OD+tg3w+iXbQk5l/ObCOSr2Wi7ryXSf
I+b1100pq0dpX5IPtwCKZISSFnKfmiqw06qAiAEA459bmh0bG7zjP9Mh/hAeNMwhFrYkSR2CVgxL
UoxIOJwdMGAHgpca+FEyjZrzDOOaGpwa7Pg7sHppxGlAUlKZEGWEmG+uZftQqgDErKQMRV1UVfgu
3SNDlLsU12QmmgSCpWByDUv7UEjj+qdrbtyomYiCNEUhrWJbbes/Nq2l5KKAKosqNS1rmak/BOnD
xz5KVBjg4DeRo96wTdmW7LCoDjAbRLCApAcRLNBAb1Xb/wgkaSnyGtK3e5orBj+a12Ei7mMd9eyf
Tt1/gHbwWt0MHLWWyMGPtjIluhYKDKuRynTsieO+SA0Bh0cVfpIymsRPWoA9XwYWr1T8gd3qjwBe
a7cM7RmFswr7QgConu3LqgOFgsbeENqp7QR1dQPG3KDWKEtQe2mNL8SrNbhCiqEQBQPA5cyKr4kt
UInmYtwgzGqYbseKhubjZcJisNJsvIZ3NVcG/dOpyza9e7FHkbBjgi5JsmS3N9CFt0xFuLBU4Eu0
Lecsp/mxe7FCAQzc4DUvf7bz27Q76yC/Lq2B8qEyFmEhNty49zlwvPh7xijBoUx8kHKvpeh8mrAl
kP0OqYqB8p1Z9Pl9l0aSLOQBKMcBRe8USi88ZqNDAnoADD/uYUii/ArsiWaSmU8EeXv3boY1gBLu
6UXa1j0i9uL20RB3KXIIVU2iw+8bIGVLFp7AEhSvfNZYvHgtCXgCLAIcVElsI87iH00J9M7Y31p+
y1Hgn51zfy3MAbuVvDCSyq4ZTF0IGsqtH7CS4i1SK3xy1DB1MWrOIYlBJrYjgCiocuAZ9kLF96Co
QVmfz2pNUaGsvJ+s3x+Hx0NVaEDJVIz2nS53W08+iTHIGe3G12KXHgu8YgmBkrh/sAw/vDGOqpBH
Tv6741YD6Zp4jIfuru7NVwhQWwgz1pMhMhGjnlqGx8THHlXD/l9lvEu0Zn4K+hmq4PTWgyaCWq9Z
ajbDOeS/02irMeDqOa+YIZH9DehSG//bMgNwXh4agCm6cS1I6Xwmnednt947SmTB+OtHngIXueoW
sOYq/M2oU1B6NUw/0XyHqr+aonyqBj8QFj4tpXPtGfdKMAKpuzSpQ9sWcsdIAsFr2WlNT8n0zjpx
Q0I3tPbaQO7szZeliniF2iMc0CHyoPRIsg3eBOE8D9wFwe6AqHJZhZpXuDhzU673C/UV6AQCheH6
QkbYHkSVlL3STVhIiDlL/Iv6e3sMDQ/JFY9BdOZT3G8uodGwj1xmuchLt3hqDxWaND5HAh3PRvG9
QZC44l/jXXAVAsg5F03X+7EG2/9ID1UMy1pUGiyQem6QgpYYM0MS7akQ/IPeS6OBleKEGlhilMVc
gn8mml7MxraNcp+TobEOyhLOSy1JJvQkMXmvUVlA+a6Ic1qEO4g8m/2oSiE0eQwWg0k1IadcmIAa
w6MKV7ScErQ2bF62EFANIM2kzj2CzdGBJSRhJN+xxMYZ9hG5t+iBJIkhON/XmDmv2OU2GKhUte8j
rRyHXZKh4hGfjfuQXQKIT3oT+22feSBw1NjcbPQgiiL2BkMxKC+LW3VqiwkUZhxx7ND8FBje9wbR
hO68p+34gV8tRsMu932v9dqMUuqqV5dxT70wG2+4QjYMSj8VUO2kL8yG4r6rS2A/M41BuTRxcaBg
2F40J/vbn3MYkOyKscEpdWeJujXEZIbjivjGzN5P7kHzHc62w1qhUW5TgItMn/Mdsledi4X0uAwf
dBlBohscNk4NlK6cPFC6pOaajm347u53hxgbG1x9efgZHQCFXQQj2jHZoj8L771c9AUVSe4yHinH
IgllkKGgphq27AtwXA0MAXkxUR7HlkuX46A8dbGmcgPYrk8bLyaA5iheJd0dltbm+cLtbBzK5HCs
J31XRSoMtN2KaJbYUQWzvS5IJd5Sy6+RvM4PK/LhakXs21yBR4/afXrywJJn/FW8H260j4awF1By
/0frlouD+HsGOxW8GUCtF4xTJ/rweGKtU2f3WuVYpe4v3hmXHnt8feuee+pyCpeLpEk8StOZ1PBW
wCakQqbaIRP7xZDMkb0zd3BdyCpQkzdeIomwYUjPNn2GRoVzIBAsm4SqAFWqBvTgN52EIXPoN8VD
zkUbkFD/uqWndHcNz+926FTq+CIFWleCQDTo0QFIkiCJKP995c9fgmtM9m1U0X7REjiaVKAZCvvB
DdIO8QowvHOoxPXSDnK4AY04aiKBfjxfg2fY3fyW+LDcmSEWutuh/u8wi02rE95rB0XMvl7NNZ4S
pg9uqmzou1zlNWlrOlGj5dOjFLJNRDszofLNs2OdqXq1w7OII1jBx3hMehjTXnIBEm8cCGzXEZ7I
lnrCOEfdWRQD1D8lSMdSJdBUqUYLs1wNX+Z5+UvXBXTcJCpL5fIVJgcz6lzbZFgPGwe/2ZvQ7r7i
YWuLDu7ZdDsaJMFGh33P7Q8140ojtkrzMCYfTvPYkZOxZNtin38aiVs3E+VVqZoIH8fRXt9OImmM
6aWU9ibAa2RJHSWoo6QsWRAHgsCSCAtj2CENrAN0Ajsr2b4DJR/Mz9cBf65zMRRMCtTd/uL88yXn
xPsdD7SMXlGPJF+c9TCzgZUdmDJKj6QmXesT8ezBlVpESjQaHDGbAtiorApEPeBRB16AuirL6oZb
eyA1ghaxBMPNzQXv5Cx0ntuKyB5wUDJU4ieWv+FDll7Gt6ys4Od4QIJTDPksSTfDBgnx41ZSuAj4
/P+IF3mP0oVitM9PzeyDh4gr7gFK5vdylixSjruQSFyYv9bS/9LVPUEJVYUQgDgdSUXfgEJtA1kY
nFjBcqISA+jk0kitA75VBsWvc26xFuX1SsrAfeGQ8muPGVyLnK/zDWtAxN+tYAq0k4oXXdYqNexc
3l82DjJmfmM0iyvz7QC2mYZhZy2c8NtE4KfKnf92LfM+8Rk7Gbpd5+TTfrzcgi3wt+kxheyrvXsY
mo+Yd4NCwkU4E8pNuXYSGY9bhBrVFTP+/4X8L6oV2aAxrPQJHXQY8mGlkiwxuKP0KhW5cYwzPi6a
mwHWA6CxnkMun3/TfD119WZXeh2zLvN/YKz1sRt6GmU/rlcw/6OS8Bt57xiq83+dyWn/oJ9GjPgm
H8cwXa+62tv9DAMDXkcx4ODkyOLHGmJPydHARHHf/xhX5Bfs0U04KsgtZxji+kYkUg3iHxXNx7/d
EOhOOBOFjup3NNxdyP3rrcLtECztWfAnOv2J18vb7MQrE/4fcZ4PTyvLbtjcCABGqD5k8JqWb5Ck
KU+Ecd8WYszI3a6FL+3racbeG2rlW1j+5UsBlj6CAxmWUo6aVRPtaYrfPk0/rpn//0oPhdXJVDLq
WR82/E5CpGpnwP+bz9mJOZcoaenR8UUEeCOsTv2oTIz/iDI7r8phtMzD2eIYBGJIp36fBeiD3gEA
AaQUjT7huN1hTCSx8vSuc5sX1BNZtuXO8YQMtcia1DStcNAXTgYjmRPwtbEFkZ7nFhVjm0UnWUkq
3zhAIL1zKcVbSkSglSLoZUvIcF0i4ExV1hZIIXbsaOLXs4R8ZQIeN78Ip1OuJxWmYQl6UvEER3d2
ow3WKnfGAQm1IW4wX5OZUaWIc5EicKoWOSBJ/VP1gDa66NkAGft+4RgJlkzaIU1CX8Fk9531aOnp
Pj8s+DmO45Dsxzkib5X0+FuqaieGhrQaSS5EZE0PtNiOi9rZOLYwk6P1qFhmEJiXt3U3sxL9dg+y
GezbrDjfdpqxxCTGgGVdmR8QA06TzjTIxhNUzSJZqUQYucWCD2DeSyn5jACoDq42YRIQRaY0HCVz
R1+M2qxF7WHM1UhXOvlGrsBw7PitP/V/m1HwXd7ifuvbbHbYt5OxDp7RSYAIZaOHa0WlhoBwkUIW
+RZ0q/b6vlpVoRNjytaEs8x3MXcRy8mTQLRdYx3AA8YvBR2/3lJhE/qAHQdfbVu7jmborRwkVIJ6
AMxii2UStrWEZLSA3nKa/fAl19X8t6H0bi1tqrU1uOye4tp0wnNJ3aCTULyy95vXbdnAHuhTS1lf
aAgm0PJ72oOnDNLXfKMko3LpYSQkuUTKFa+z69PExm3QrWBuQj5e6bxgRmK4lrn3q0/6pcYf3sJT
seDXfoklGAain3bjmGv5Hoc4B86GQAOQKIX404e4Ctjtw9AkvAtIcHeS6WmAYJd9cfiJjWMp3SJ1
Qw/bRtatF46FvQ4bl4hFlFBioKB6z5lFxvT2dG7UtXKw6Af9P1n9VEZN6A/iCFrWmJxHAcxHIbBJ
4ZnuFWqJqKZ81a1dTQUeCulf/Nuldq/sKojGeR0Tz5oC5IeZNiSq9mlwVRwFg9JpTcdS4pWz5D1b
PPtpVnYeVr+vXB27deG01m//G8ygGUVtK+Ui+tHchvo/gCBtCvYTV3iPJgBY658YEw0RTru452+l
xyooN63qK3lgcFEf6QYaERBHmDGmYMEDW9ZbSXfs9JiEx7TZnsl35eb7wJ0I76MvFQzEKxVvV8hu
4tpdBYMm2QbkwNU/4SHssZg1iDra7hEphOpXt8vw9xcCGn7XStbWwqafhyRRMmwGoXhHJzEq8ZMs
8GE6Vt9EddUCgM/8/3IgElJ8ZeuvO6eNnMKgvSP/Xowlk+sxIaMVCJVku2CBghvBeZD7Y9ZzGbCV
YPmodkecGxXdYnPyyCGjk2mANibOBae2T4aLGNSadMaTeUl3C3bqrf3hsCMprurNwpjHSxByJBV+
D1kDcARoiaOj2zwI41Z5I6qznaPCYhy16zVYoMgi6W39Vj8kfOHNC4PLAnCieUAcPpN209xAOhUD
7ohcant30lp1QDZ00OP9LdHVRGgJhP7WlT7CwniTsIBjRRx2u9pv7oRkk6SW6ARjgIPKz25UJfIr
MfS6Ed5espS4UuNQmiYBPghnFo+9/KM9fa9FtqQ81YN2pluYJTbBzdNQgzsOddkjNIr1YNWZLCOr
EcFhg0aEiObHO9aMcNP5JEqIINdwZzdismFQK43QX8vxy/IZQs7n8OF3q9svItpRpsK+Ro6QOGg8
FnAlLafoY9IlLJvhzkVS3RGdk/cyTFjiT8UaBq9qCCZr3sCVdXGF8c3zBfYylVm45ESUewj10Zyv
KYTcSWTbE2mUZH/YpnraU54QuhmZHQ87FkmjUSZ2tmhDouUl1wCoC9j52wgIDeeaIJX88WE8HrNI
w++XE+zEanzGJ9rSezpJUKh2tSEjrbI3g/vohcBpTuS6tXr+pzmonE+FOrpjjskx3+MRHu0zhOuo
IhKMIitZhKKT+IJHfxZrCFDAREo3n2qL97KL0SAOi+C3CwJD0mYNz5ILm02dQV0Gx6iAh69C1Rjb
nHIVPOxJUu/QWPYBRHc10KR9e2fqAKIde3bWVKrnwpxCtwhbqShR6Og+E2edZ/2qonLmFWTw1F+v
L8FVxvbjGNqoZmv3kT4ATBm8RWBeqMd9SqF/cwbpmwE1esYdPuNZnnS4o/ePvcO/fj8Fpk3oxmNw
V1RoLLZ/n8gUg1z+VnYDJ32HAtclawQD7bXs5Ukg21IANeajkHsctamlOCQBcVif6fri2rneKAN6
8tjWFHV8PacN2Grrt8J43WjBl/ecS6WWLcEubB1oNZ9ZnpY6KYMhiqZeoWk9jlM/Kk9Ysu8P/t2Y
3xnMExtxRVMdvQmo8ZqyNOV9YyscZkLXCdGfYWbn/2Uh06YLD9hkvuh55y9lHZ4YcxPqkFK84xO0
O09+KpZaOccwpaB7CIBxgODTfkVMHEoJJL2q8G8wAmGl8u8S0pa6Be9YXR3niysFF2j6YXRhwT31
E7KCbkF+g9lKuWb6BtoVQIqM6jO8hvlMF3KyIhUNvDfhqrMuJnxpgI7gV8e/qBkUf9oVgOYsWi5I
yfvfeA0SMnkcB5zz3f2xB1i9IGrHeaqjmzpK/YeNU8xHYz5BJENlYcbwM7Fk9sl5jVaeMzG5GPsl
/9CX0XIsODmCW2cnrSeux0Vs5zmUVBf0oIuadMf1IWXtu503NpNzgQ9nsY7VOS5VhgPdZ/xrBQQR
lurzF7vtZa+fvZrwPc14dtgsPZnmkaANQ81YhY8AT6JIrmj+DNRqTUt+B8CtCkjMtXPMNhmQ792m
WNHPfD4FUGtpwTol8+0sT061jx2hu32jL26pKIdJahLVsG8dWM86x2Yx26NRlHM/YmY4gxlPnWsH
y4rd3/DS5sRiDqWOtUpZ2J7aOZNqE3mWIJvUk2BFkGNcLFihbwgLrqlUmtm8zFvZ3jIIDkNnkfGq
Ys4o3ZzdgzGf5GHczXvd0cc4tksvkrhQnD4V6bcAm42uuAhcHwUwAHFVn98dhlczTN7Rc4oo1/AD
olGOw7VGDz+diuL18P2Gvm0+QtpQCjTrPT2aaRFarhjiUI5VGXxECXHHxzwsmy6nj962wPTWlxbg
6Pq8uFaCKvf4fR4KyNd1yfA0pN/bupOGnEKt/vu/Y+NAV7jgPK9FoRiFwu2xcGx9AUb8K86oOjrR
NNZvf8AkVxCwIfh6/auj8soclo7ZgZKDkV4eh5l1YClK9hxtT7qwpO4sqVSI9ZPXFhtICxCDbR5Z
kYJXt9AgYcjzbzvSollMWovQSc5w65ziSZFj69Xz/3wXxmkEwE529UE22SX0xQO8nZl7doVzHnj4
z606dITazWJlU0BJ33HBzB9wldOmcDzI6bzC20XV8vvVfOMNkwWNbIcmDx8prdbXo8bfv7w8HVQV
WaiideQVPPjTEE/GB1LuzC1r2yWxSjjZONvCMN6l0LLYHUhurDTZ8rZhqwuSepxLaHggDH9AZKVc
nRXzGbIWcWTvA2p2FB5PnExoZGFaQOyva2ruZiNZ5UrtSUvKLDzYK7NnhqsCduLinmTZfxWnJtnY
77Ug6EHUQsuDMMMDB5k8VbCPV4DFyABxMdqCBPbh3yrOeJNxyCqzUCP+GUftgJNIA133m+bGEDN8
5/VzhebYg3aXWWU2TAcfHLpEAge8A6K7PpDzjAKvTacRXueMyQ226/ii7jIswy4lW19yXyULdRlG
SlwseDEwdhPjHqL1O95okT3vqkVEXgnpLsIJkP75YWT1be+M+IO6kgjabgtb68D115Om7lDMiL4m
woXK/5OPRiJIYlIv2Ydcz90qCn0LIqUjeVAtRT8mt0TBvZjACZ8CA4tFQiR/GhBjffY0cB8g5d5a
qw2l5BERMPrkqaH2ZSZKvR0IXzaJS4pbyQ89Xbsm4+Av/ctqeSPXk8xUVoNg1ttm4/iECPoZ3o/5
T/m8zUORhXLKlnd23yfQhG0AmHrXGWgOCZ0XUS03Yc4uTGG38OnR5NPvF/vJtJQcHBg0qDSjeMPQ
OVhs96u3VyN7eN/1ChOtOVJievGHFILma+Ji/0FmGkI0OFyOG1XIRfhaOCWq2M8FQ65dxOEPNcYt
Gg7mtaKsUuXNv/AEb5ayafWcT7l6fQEu52iwmyFQj5HK19/kTCZcruVGeaqRW1iocT4ZHCcYR27d
z/HzEOJmCVamvf7HZ0K5ZBXuBFDp3h0lUP6/6TazF4z2T6R41Jjr9PS9VMhC3UIPrcGflplFJXHG
/ADQsb0ewGPOpccCYVQgHQ0TqNv+KnUyrz/Y3wIQ6gEvU08BGitrC5yfLD4lgLIOT36ODa6INW7U
+PUkbSkq5uFU6pDaScSOsLc/BYJdfnZ/zdbLSX6SdPJdl7zJcWPXEBvPpKLw8CMZHHss3Jijmojt
GbKaWXc0262aiXazpNjePGT7XU7FnkIuQzABaqStwxxqeaJL4y1hhYMUOosi+I5SRARCgbTlgE3S
4ya/n8Eay9aoCHYZmFHyd93qaKs1ShjZ9soy1bGx7l14YIPlVklRZ9q8hsdTzNYk5QxP/Y186DvL
+58IxWmF3ERTlGNn8VxZbwX6htf/5+wDt7sXwQKiSVVHwdKvWVNxGf1yNEkiAB7a8ygMH1sSOV8S
zBFrxnXZloOECtjCeWSRFPbphyUgIXdO3UyKuZrUiBDUZzeth6O3LLyViFeqHcWzkvcRb5CHNVxM
RSpVgycN9FFkM/vgSCbwkzzYn9C9ry8QmHsemde652vNjZet2wlLyQH+J470kqDararfvBqB+Rqn
wGHZhhIObPvGHkJbYuxzEHRttXv/HhZF8251/Y9zg9fqmqzYjW4G6QqYmNscFlIVDxc83/XqKEt9
rYvPb2BJpu/u+ORZyFy6U18qKeJG673GnixbExH+RLpBxGxSWsetPhfs42/00exE6GgItE5EiGHP
/yOsigIhU0jAXWHJbt/8AFaWlJJnXoRXUCBDJx9HfCJEqTIqruq8Jni9h3SlWCVTVXxL9yfWM8FM
6zyaLNsP32aEyt0a1e/bW9qESnXKqSL6rN/SPDwlSuuz7oBu1iWeZisNvP2r/OU5brLB8ZRWXEAE
4SpppH1H6vasJc8+eRSUsTmW+5m3ohN2hHhsZh+McyeC0eqpThTlYgcqZvn5CHXxpMZnWWmvl9IV
jjABn3/VEHw3rdwJYKucZ9dFV4c2015p8dDvakM/p7SC669yeK6TBpekbAaUFy8mZXZ7AzkpT3oG
KPc40qN08OZLpF02/T6jAfVPLp6Z5xakwTE/fpKW/9je3jNOHZ/9p/l93/9BpTZ3VPNA48EW9zay
BuKWcwedLAv6gNLT6Pwj/3saO1Jr5o29UgLkdQA7H4Fy66eheWIeOa/ErI8O6gRrzrKmSf1Z7CwZ
XsERoq+/FDHT/RdvBwL8Jmb1itIDURXgrSH1v7RwN8Yj65wBLIlC2kLz85WlEUm0CtINcPTORMgP
32NnTVU/1Vx0wOm3cwj8AwvkEH/GMp7MMYWuq/haWsSsGCaWZU6doZmdsBfevKS0nlt/5oM1N7i7
vbeHrF9QkEKZjZUWeD54gIrN9p9EMNadK1VXBveFPfRu7fmXTUeV+oZqCtIa0dEJbJ9er5c9ZO4J
1w6h5QILSM/OdkgmzwdpqHKYERVMmBx1Q2jf5DyXQLKYi3C70dunGMCKULZqFBaMX/Yj7L6nOcEt
T1uCNWz8zRctTfru+kH9b0l5xRnhg8N42v3FJhIs7x5gfJC+8RdX8EZreFPhK6akPB4+zn6aSjfu
QnEiqiZo6xNmCCMeWlHWsQK3pilZWHddVMmZjoVCMYjYpeiFVE/G2ZOW1mZoaikgeTYq1ohWOcrp
GWpBGaxdgUxFOkh4Aw2ML0N861IzEi382nn+4nVOYKysEBsoX8GrcTqzaBGtFUmABiKB2V2gd26r
ymjR1/l3Wrc8KeSJd5gSAuDxQPe9Ks1LIAe4Ssv39rOc5iqxj6r/7i8HHCeKEk+LNBNVwFWQhp8y
ZEjyC/aswKyjXckwNRc0NyXQyB0eR2cFZVZMVMwuQcKbjwSYvkW3BEMR0M3WTYNFGgobLQ9sUNen
qC25lT1+3icb6dR7pBG1t/j9P8Pn4Ai9eFvppg/lLq8X3m/fdo64wFcmNqMtXpYIMI4Tj1M0B/Ib
5UYeU/5QAZCtV1QqeEVZ65+Wi+coP0AmHjV13vp715UQftdeONT8F1S73Xlb5FC6Wh9WW0I83UGn
hMg0z5QQ7rMdgTH18UPYzX9xdVGAPMiFbCO9OrBdDWd2VSHQq9JHGUXvHv7SxwFMAvenxWnILVVb
30jKtOvgw/EoSKGVTGCxBPDagqgKqO5Gpem0GEB8Ej6N9yF/XEABs2W7RUxSyB0ShB9cznYOHx/9
cPf2aU9p5RKzgYaGflZcxfr30j7ZyIRwjwokvqXV9BgG3mN7/68n3EOHjPd3WnRVViXzkWj7aUKi
TshQmt/xQauSmbI0Cx6zjQZrSYBxJHgxSk2wsuHQRjG18gJmLnpSfqJ7U6OpOVP0TcfoabTgPeOw
F3fieRHA6ZP74AjRopCbiNHLwu4piuwCRBrSkf+gDz+9p21C+dUn3Zbog0AAAgz4JltTicbjrBM2
YyTTWtXIGB1+esEC6wE/zfNRMUl5ZlFvzEzySWB5VjzAKPzioI5cLByqwZ1guhYwNHViV2A7MPQX
DrPwBGJJBoslVXdjD2gts1KIXtz4df025afYamjNK+aCAy+nF67hIVt2I9rkdZ3xOrIJk1sdPXSb
B0UJNhy+jCSAHfdRpX5JGHQxG/xB+xK73dwlXcUZUwzRpBav0Ci3H0by2Y925BeYu2MH1uPIKcN/
bPzCGG+G+hzi2+J0CHKVWGKzwMt+N7rtEH/qLltTzng+X7/xmk6GNW2gwKPjW9ueR2yhHaZuWp8O
U8d7ZH7mhpvT7T66AraFhIKCIr54FVmT+eYhcvTEvLWqs28o/1SsgPrtQTUVcPZJCthqgrpc7IwH
KOJFydYGEA25G3O1fK6cT/lyuBHSGpMUjCr8Y9UXpXJpvqUOFkh8npfV14fSvry632N6kAWqoHrb
X2EHkUduCUcSvqbu9V171LeDBrePVPsgJXwE2mA2R2oG+0Ts2Bi6BQnDfLc488Waq7bL4bzz6umM
FxmueJVws0y5wwXMPf7sDLnxfe9SMem04Yh5eCCAqhZdh5n9kEAczuqIq3X7kzNT/68SQQoqYqSw
fulqBzeCNSjBK080e7YUcnjsaKeoRwpmX0QoOPCAWRJXwAwTQ2zuAtoZS8UtrDH4c6YLsRj/0FpB
kKZvDwmkNyIA7Nz63fpDnISU0bspQpEqUlJLpH8ajheIYbb8nxxIfqLPSz1Cj7/KV6MKGwUKhErN
g+Uc5uEaQpPBkqR+PJcn3yWIUJ6fZdB1C4qP3X0EkjZCIb2XpzrgkZcn0jhavgR2CFqPPg3mFaDq
0Ie9dXU7K0GBuqsgnMS94f3K7OmoTBz52Mu3dZY2sPI1U5A3TW9RyuvHZwvtIVZhzNpvylrdChLX
hD2APazqV0vzY4/OleXwES43Pe+nxmG6b8wgDwJL/fGuAlbf8CPmjOdD0AtyFHFLNEnbSqz7RqHC
frUIlvkrhE1ZnHNFA19etiAjfCg6CJq2AVf5ZZAN7HcOpZVbPEUP8MQWx1uNCTzHn8ypg9dDqLRg
gLltGO/FGZGaIVdSWU6xt/JbsDERRHBOiJZTJc1Gn4SNDc644ce8kH4Z/m82IrTjGL91lN7OxBLF
eLLEXcmvidElZJwkWBNXFczPuuFAvDBPondvskiYgER9LdRi3cJJtMSjDRU41xRLLDQPQu3CG1nb
lkPWIEVEcY2jkpWpFbkCrG54RJn1txo+JEmVLyuMANeKMDHW08q62t8oij2mAPYM8UwGbozOEbSq
UGQ97QlhnZVgUKBUhv2mNbTkOy8fsIJvU6ChI8DNNrJlLcAfjjIKPC/L83Bc5WMIF7++b8XWyOne
sbFnEs2KgVGLLjb9rL8fQ2cTslJEPP8CjnytzoW/MaIB1Ow+M+WmgOfNGjkJOmRd8rAaRCLPsGjk
Zth4oE7eysAR+3ORLK5+JOdp2NW2Qx8VKFHgmt5Ij73/hvaG+D62x3e2bgWRgyu//uDDFFJsujfQ
s00gK86igNb73hSvyazy/6mukVgoBhatrAsLEoYR98mLQJT2B4vMz01cH4u6d+tEIRK57mSjK45z
B04S0Re7OVlVzyR8ljLCEMyOI0oAPxyf8jTSdCX1voV4MCmD8Q+ICHxzaVywLrkYNCrAO/yL3rJJ
2HN1UdApJoFJMMgwE+Tb2hYqy2WCdogJ9qHN9eS2vbzbphnApF09NMCmLpfxqiwtNO97vPJiQIMX
8BNGTcgOERGWgPU8bVzrimPg2y09Op5bk3rKuJWFA14B0Z0oDq2YDg/Ann7uVRLxsEoHAu7gw4ll
BjHM/7h4HOkzMPNTA9M+6D9jtuNGH0SuFMisKm07uePkgvNFdTWx/d+8mltx9czlhLI7lmIbscA9
bkuwOXkTS83HkVQBu6vMk2OOHOFj07H67K39SL+XIULdhmGBZbd0X0nWdZOkf1E+hlo0AzLAC9H+
W2aew+rSnHiA51S2+uvYOYMBLSf0mHFdyKwYDFg3nQIyXPNKzd+vlECflK5a5iQeHLd2KRlun3ky
WQy2Uy5N5N6FzDBIR7au4B3Tb0wBfHDQxMYVnhu1bxL3JoNcUiSgfpVLUDBppAfGFcKL/Or1mmSg
03ykg5bdU/ue6oDqA7hGjvi7pz2RFyTO/fmi0h23FTOYQdX8g/Rq1+ThdK/LaCoDf/zs7xFrL/zd
lRfKmkgOdUKa3G6XT/HRjyDV+oYKMYCU7Itj/rWi7+DLgixkhzpg4U/5BEkLX76YIrtZYnhh8lWD
HtXZ0rFpJ99/f+Ul/e/axN7A8/hqdpwm8bx9rYBwh/XdWKtzIJgzRhozZubazaQYoKWw0QB02Nd/
tpvoKHr4gEh5/FAWnsNqLCkA801dYdkOVnyRtoaZsCHwiLe+EhL3mOylTPRFMBUgRCooVA+E5Ijm
yfdpuwtdFaGZ8XTdO7zN4USpXgG6BRd7gsn5kB894PDAdd3qv37wrIxZsmkVDltNlAO7i2a/of7S
7pdVkmo3ujiyeKDtzMMd+tbgI71WpMxQpSH1cH+hmSG/HUw0dAVd5Wg5BNB+HB4xg1Ds2rUFUarY
ImJykXOquTTcSDRMh09JkRHdX+rTDXhqWibWL40U5wF/794t8QGnWFcDF/XOwh9/pmMDaPjuKlMA
CcTiovb55XRLawY8rkKtHE1Okmp4JU9qrtNqNmGsMGe2ONS798SCX+qleMwOqWlpPDPnH3NzmvfK
fklmpWenWhMHX1mndng4qCvuiz1ET/4Y57Dvy4wjQs5Wfz+vWs+TPIIbxpn27uUlCfNjMh1DJO+l
liZk2bkQWKun4w8a0rUKrDF0TDQkCLYS7nDaY5N8hgI9t7DJdgAH/2v1V1Qg32hRFburNl0xKVbg
h0hmtNUa/HNUKxx9FBDVYKWuTBUjIZbvJ0AJmugxQ3zIKkh573rXZqCkLV7jLnygjCZK8OBw3OfV
Z48WbkHPRWYFxbQpi650qCf2piz+N4RHAHK0fmM7yWkH2ctv6VvJZTgm+q3yUbeEVCJExQiepd2D
PSnF0TFyYstW9VZ93NB+Hx75m6N2mzpKRNVxGLhMLqROji0CbiLppWhFU8NzxneS9+rJMUevjypP
KU37tgRIARA2wKS7UqHMqjh3tBqPSAoSqWib748MILPVrTV4RuNMPH9VMCKaY0RR+OKRXm36SyPu
GcWpiCOkON/axiz05M+A6zmcdPLgL0peRUKhfkevCDqCEa0GjnoC9Tz5wPWjDh1wv4LaI+rO6Jx6
ELROPVWu+8bKXMjMsD2+JcQRla1pF1DSKZ1sT28w719UsnUszuNJRmTl7AJkEA7qCWJrOeiRLyMi
fieTzEaGVzs4F2fG4Ly2Dad/hIdZCyEOxsjIRnPu225bZoj9UeLPzBD3wcXD03B1rollxt8uHS9Y
sLWfGnK0SCdnJRKrftQZb29JEoSAWhXWxSZrO1FllOU7pE2NSfzWXshVhchs/pFzleA+i+88s87L
BUDZ75PbP/jde6m/WRHpnZZ8sMt6RMd1LmOm52PvBSOAc5YZRc7HJEm2noXDUFKlEST6chUOZqDh
qrd9RlHIiMNuqsIhYiwJszWAdCJd28NLt3x0onaB7TCwZdCaoZUS/GRNBhCF+4kd4TWwME31OZcv
Nq2EM1Yx24sYowMsEbeMU1Z8KYYBLrMfUoq4ArIUqDGf8zUtcIfe4NletY7V3lkAYDcO6nbuGFsv
JU9bgA08iZWMKd84DYZAOGeZ2JhifSl0ldUpYAq3tjUr1SDDrYNMOv+tAB7SdS56UkaDuPkUlXf5
+kHpGAxh0L4EjkHyezw1CFrcsPMuij/ne5xa8thx3YlkgXlxyGk4FV9vsSJnk5Pctf1utST2Nyx/
td+ajFNO8x4U5VJrOVqm205kADRsisPHSj4BI5zPbgoff2aJBVAzx+Lpg1a4+hfmcnObMDFuyyIp
wb+VED/kOjM7gHaUZYoc8rKXOlbh2aHPyQmrSCt7iSbdlzZ5uCExlO3Xycx6jQLecDn1yMGJ2btP
ODn7/5p8dSu0R1hZfCiFZGiyqygCmj7fJDXs/nLrdAknUeHu8yXrssmzqpY5FR3dqp2ImERBuhYF
JCDul2VOsqEJ6aH3seJtecGGRjkvKHhyiy/X70x53PxE9r++4+Y3lwjnyIwrkW/OPlGXsjUB45GI
yBZ8py1InSl1GArbDFI5lWlBb7y6T65fIhGzguiHq/vVgTHENERjSs+IjfVnPxSkR8pLx5EPWguu
r1sAZVLyVOJV82EhBcmvPPqanX1tFLCtMRWp5H6rnx1iumkHPFt7AQ527zAHAE29paXl6kGgGzN2
um9O0+mLvO1NrCs16asm1eY4ZkUaib8bga0ZyAiWyvbDE9Pxu25YpaJ7DOhLl0aZcu51Q9+YkuFC
K+MQDqkUxaZn1PUJNK72+xUWTGJRC31wbbRKf3D/uuXf0I9JsiofyS/KQsvbLkajsqMEWaym3waE
VhI6+8H8LspbyufuCLeWzScG3hAB0w3bP/YEJj04SiQXNcsWy1xkCGdFkhsdzuhd1jlNkSBGdi89
KVpyYlb2b4D9Yj6u4WsGeW/vO0LM6TRsz+kpC9t8TOx/M0InTdGG0E4AxKsuruZ53vIMD6lRibyV
ovzqy6gTIdcqW8u8ageSnvi1y1lmHfhBIxNHKCk21IYaXKy47XdlrzBlrPxf4d3VFX1DlSLYiEdP
1lXLaugcXOrLlM3ddGx2F/xNBE/2e1L7aTVk2fzT/pN3BJLaV+02TMdiKj4fItOyG/AUVrqFmooX
6RpXd7Wz8xvNM8A3hZEqR2oOY4zIZ5A5pqo+2irmCe4FpESknHPD633D8NbhFKsVEl6oUesLutGP
fVaCkMpm4KFPN5kwMH9CFtRYlZHVmjjNerstZoc6liSPbMnmcSKW2adtZS+1urN1eEik21FBKgZ+
buM4sSlFqK18dWj57fANlCE6QGsjaYmIWaQfE+SKfyRUPkMEXnJdoa2jzB5xEodbOztt58WnZc1T
5St2SkMMOYF3jTdD7fPAPgw0ypHjz9F4gOFqGS/oicM0ln597yOG4j5whmm0/bhd3mZ/xfOtJKiW
cKClmQ1d5sERX7d5K2m/yb8pJUiOM21kNyTUh/bUgN09xpKNWnmwyY14w1qPFQ7KEoeadIyc5wNM
OHCsxXZ/5/yf4yOgogxNnT3QaR1i/ILEaU2AMrK56kVYyJCxXT87WALB9K7y29yJ5QSHzsj9/a4d
rdE7Mmw88s1/1SlBlgZnPOawF7xZPGWwdV7kRTRPVmSTw2zqt9rdg7Hza2IfuArifsmC+6WwwyPK
tRzZIY+ECTNhLN/XSrl+xyn3x0ZK9QMfjA6ozGbZrw1Qdii6DXRU6p6bMZxGJV5lkLE7If8lcWix
e3nYVIs4xsO9JIAu2CXB5abwkLuk8b0NqmjJlVUc0iwz3qtK/93fmUcvvML8AC3lscG8RpZjEFOE
Pj/cANUKVviY/IxHcOUWEw9ZJPlzPOWXWFDZO5sTA5kQ4HDbiw0io314kGO6+abbZpCAogoJpQCN
iQlRgSsOrzHp2p+Qfw6AXqcCwvP8Y4wzNGkFp5eg8LiPRBAMWOSv++bkbvB+5BnTDBeSMiFL1y01
lpqtPD4Nhz9rcm8W7m8yH3La1O5x+KRIsXnY2rwOj3sCI/NOOHy7fG5z3YY4tftw6B6vDwweAjoU
v1MdjNT9PPFHs5O6geQyhq6zAP5V5KLCFl1rowx+RdRc/CJgLXHKj23J0vFAZp7drX4vnfNYhFET
LMODk2Jyo+d3FHn/ZKnZfQBP4YGomaIGjOHKqv8JKc92FEnBEI1Pf+nyRw+ip41fIPpngM+DkCyM
3E5/JRjel4l7+wfnvkhuTUu2A1FqnV23lGFYOsU5nxURUnRGd0HF1dwaQ/QmFqTBJ+WsYWegmg0r
iku+wRP1rttlhVApItMbkRlPvKph1eryprJ2dvcpxKsEeMeAjVqTPqEd2nXCSOaYDEm80OLhOswp
fuLrVQwexYwn5b+t8ew032ZToSCVcRDBUtim8vrbCALKP6qZjQR/4ANptcmOOOjFak8TKSnF0bU6
Ed3QyLZG1/Ko12zvPML/8dhogpZkdH7a2zLfH8qxc9aLKRHt76JVGJbeq2wJjHCUoiWdRYLBKM16
V7TvFzDfRWNqs7Veli8+v228ufIG85GZ0CIpzmLjUyJmxRYkoRfBQpBAWjtmqbF3Fi5fFOj+ErLY
11v/a2kTGeXTSPZprBl3VwphoV9tYEd88Jwq1pb6wmYiFtDQbZvX6U3C2+XWjc0kf7AK6IRQHQAI
rBEsH6R+Q2jGk2lce/b1AnOgwU1lXQH5CLbxxgVXtYQaW1flRDh32ANa+JAdQoNxdExPON1XEXjP
/CLPrI8PL5TlKKXanKP8LpwlU8axwtu2cy2rQiTxTpTeZ7eZmnxfqaSsU8yMY8FnQU2SXSd0hhy+
7BV/p6pkbPtKiEwgEED7SP1OpFPL2nNB+yYUAKnlPtEg0nq118KKOdIziYwYGrPAH5zTQci1ludf
voYi8tFlJSzepW9MOiH2tJkkqL/0B00GAEiMK0MkyRUv38XIg9WxFU4LO1DPPd5gvgwUFtooiOzH
tXuPR1THqg4bF0giMdBzxIxlcTHSaDn01oHetBG0hh8AlG42E9waMUu33ioOropl7pmXdgTY+BaW
GhgvUQ+A7n2yMmTKGuLA7u1ZWDpeawhz8Lw95UW8ifV4/6m4KAoFHbCEg1cCvlb8+a7OpMNkJr+S
HZcZUM4V7y2VM40mP7OoHrXs9YstrrA/tHRBo/4j7lGJ7dPWNvZWFHm3dgytv+MDzLXuTp5T41R+
MXt3s5rrERHYl5SjbB5QkmPsegR0cyha0B16Z9gJA5n4+7EtXNnvTFFfc1wjxaBJY1NtL0flBpsg
cotRYU0uzu1AIMqZuOSUhiaPQn6Njh835NynNu8SxN/SX6eWl83tBZhOkfTELs/xwE4GsHniybUK
GghKEFJ+wvH7OeeHXwXwS1z8IPNVRB1Egn3jHVj4T3FcauGe1oYVn+r3Xpu7y59aW0K2PRgQPUle
MoXMDyPGBiCxA0H2IH1kAB/swm+aDoLqE3QTIfLHtPTFghIooenjCRNfDTzWox89Y6oeP9uAIFxi
DBeTKLx/xxxxzHK9xlptXb54yfxAzwDRBbcMvnld5f+BKMq9Rl7Ja3UYtqUp6ZtA2YFteUl1TLVx
yj8zo4X1I0ilZxE2fvltCTFmlur/5fD1xWPrJWMBymsSfMJhHm+Qx2Ox2ny2vvo8Pxd+IhZS4hmc
xMdXQhzzm3u+WtjFCw+TYPsCg/V2kFu0x5t7zl9gC/LiEq4tSAoYz1l0SGaWPyFicCBK2+FR+z2d
NhonlND09xURXnexns1Tofo0T+PMjgYaypXE8x/fTUqD1KD4Bb284yMRWeGMVj9efM3Wn+pd6Ig9
BGW/uqbQr1i7MpnbAHjy2kPtgfsalQ2JsvfgeCscXy2o9VJ6jKFflFbDvHl5S8pR6uFJeBy/rvO6
6gtIvqiuZHvshtxXuWkOrIO+V/vmX3oP5BVLpYSGizrd+5x7VKLLsVqF+IklaPTAbiwCG2BHMf+d
UObQd4BrrCGeTer7UcLADSrQlKOXRwQET39GMFW9mRJ6Wi4YzJH4USFJiHTkYPp7ho1IcaHeXHFU
2jBGDh2fZ3eMmZ3RZ3Q6RqMbXvv+Mzb4VLFciYN0bz7c8BSjCe7503s80lxnXSmFL7KUjf6kk2EM
x4Ty4lZzMXb0AKyi8ecpKxUkcSaz4VkNT7xdJLVFkRiGw5G8M18RY+hNlyI70GQB+g0Yp2QdlAGX
pVN5gXpIb5hBWkb9TtjHcLyMBpXIw8baZRumGRCYq1A7G9+1tTGj2+cFxPTEBEUEzCvOTb8bUrkJ
j8d7CgsOtevz+TVfsFxQQ7tR+IlfIbggavOOT8LiYOtsybmBjrmnoF7BL95/1d/hJrj/F95425kV
QoOZfNXZGWFDtW91cxx/mg1R0qHzLRIZHZFRCWjeVoCunwYkj9h90nAyuK8JJE2yBqmez12ICL2Z
SD9S21BElNuBpsdej/NNT4eMYLuO2IQw/k+XBkAaI8y+DCcj/VigLjiBqLW7HfJwaS3pOOTWFsN0
AuMFcJfhKxI3Y1jhpwCfhfvYlZwkIaz0II7PzEspMHtB3x2myib7JPs+eOgzTz8qr9W2jFQ9WGpx
wZVo7gydlu5wWgekJo8SmfEwbrUeluBgDeKLG6PliSijj2igh4ixb1Ii4aoIqYCKDVaH4VuxILkj
DivSWyWtC0VnbLQ4TWSrVbtCKnpj8rZod1tn4k9L98v0devpUVkJcEIclyjqFDZ1ncEhdijLUCIJ
xVTu87asoTI0AqMpPqYeMOVKb6AbUkyuqi4bagQmAtQJ10FwOPEq0qi9HJPvFD0l3vcSdqZ+iT6Y
JB0S1ZFD5I0Uj/5HCWrH9I7ltCGVGSanJ7BjrZMm1xx8hztKwzbdjQZgXy6RpNxFghnuSxlFHqwn
mbXh6xtHPuAcE3A7FYOEM1eeFn+eKedSMiPyYNtQZCyGbdQxEeOqjG7rq1bdaXj0BXNSrhxt1JWm
SJ/KKRGsuyt8BTOCbgdKJ+oXUZeuM8+JH72QbPS8a9ZetMTFROjlJiWz+AS+W2qTqc4KXh57YR2Q
BIq+vhnWCiWpkkmIgPtkRzUNzLMS3aZFEcox9+/6BFt8qpT7uCyYSgfSsyuuChRXVDVqSz5szJ2R
9anw8XL25JfsZz0SA1GU4wImHiPzIuPJSHuTRRxln1rGwH1gciviVcDuOcX9pV/fCrLELtfVgXkf
rk5oegHi2IhF5ZMXCFEXsza4s4uT1ZQGmig8LgSF0kP/kftJxTpMq084EQ84l20UfjAlGELlk784
QoIB300wVud9LjoSko6RwAdJk5GV+8t5gq1dz4VDxZS+44XBT8k0qGJzsPr9xK4SWCPNKrcUgYpZ
s5QlU38Nod0/AsniHfAMWrqT9kzDEK1dRtmt3YQAROgYgf71BANoenqS7vE0Q8iJleTlRYYb6jdc
RU0K6xrBDwdrnbKRJAemByiyjFe8zf+xMzhEfyoB0nqz6qxDexPe1LgSnyTH8ieGhx57MmUcXrCB
rz0F5GqOj//GdRQy50lhxwVMVntEEqn98HYP3iVWyFFsE6lS2m5kNvYjUHiO/rCgvouHu817wKK6
WLMtwFIfoyYctvE2jrObpUTvapidBabytR6Uo1mi0kMDPxHEJFBRnkjEc/gQUjrozwQ531hahl7F
fu+Q26fUN0pgdA10IAZPpfOqcifUiMqy470y5ROO9rqZxKVEQiQlz1ZJ4P5bO8gbHV95+ptZlaD+
GBZAMalLL+txxp/0JE0NqtQQ7FMr5lZ3kJERNomliPgFjO8RZYWc+vnvq4SYB/UK2KTxJnIAwI3S
6hkFW53de0s0BodXhRitVH5HxJ01VaYWQOnAUG0RrAdkX3BNjC/TlcCiDoXItRWoDJ1+O7yzBwtJ
MMN/L8JjyaoiC14JUbKh+dM9RpYkWQbDEVu1PVVRrM8VXf+UgXD77q7wWaWnX/g8PDqswWHBGY+U
nNEoL6DTi+ZOUaktmuWVZfAklqncOZ2QGuXr9PiwsBx2gNAObMlWVdV4F9AY0nvBzI/OaE7qrbQ6
fWenTXL5t3bAUlQxEyN9avCL1EglmVZ0kRyeovkbmLf3DWp+JBJkcH+A+KFc6ZOmnPR7cGmw3pfE
uv7mxW8yXfWEG3dIm1hIeMGMtLeUVmpBFY/hYQTpN0DBDQiEsoDkxcriqVKGpmBSahogMKbl30e0
endv0QdaobK0ZS9QtfGZA6shveIwCm0a8qz2guHRThYQ8saaRjsdeD7vchEoNVu6x6Mp3AdkH+7H
ffNAwJFdlfyaZLVc3FASGG1DL5Crjxw+QTjOh/ryImRgRbDembfVbkq75PvfnYRLTQE87qoI7XZP
rQeh26+JX/oS9uxOnNbSJPWK82T457y1MOfiMGNVMrZs6qNa3ZGsShdWXLAO1xb0UKcmu0Bt3fUu
M8WvvQd4NlM8jvAbQZ77TqJ+aeJ5a/v1vPoZSDq43Kyu9DexEQ2RCOtr641REmqKoKZ5GJZzqcp2
uKM45MiosW+u/tWBKMAhmwaM1EUPRVhCK2AMvNgWU0yK6m4h0Hx4vEsaQnj/Z/Rw5InIc+oZa6C6
XtA3RWTZjOEoKUwi2k30urt4+IQTaA0x4LEPFWkFPomJHyAia7Rs/7hnhGzSBWllCyZw7MBzPq9P
mNflk0LSSsAsNqL3kGjZ6L/EL4HYciJHDVk4Rb41hlCtQQ04S3LBzHMLgpfq5LJwgFT3Empyiqrq
2O+vqRjrY6VVD9cV7RZHYobRy9LW0AN59D8d/+dmykpKd1bxqLjTD0JONzNmJ48YZE5jO+bVRwpQ
rqHG7uD/Nm4uuG7BLXB/wzUvg4dVBDHzInP8D0l6TgSodb488t19+bK4L6gZFk5wuxn2SSg+pUlA
PNnVbUDLbZSUlWJvVIBcRymX5ym4qeivNP5wjsAnWcL3l6I88NmwWj0cjIYCxgaTEXjzXNWm6tsz
MoHvohXKaA1BzpnGRZbAGoEuL2XTqMiD8faDYZY3Fr7/3ycbnGuRslDur0tLI3HF4TV5zUEMQ2N6
4GIYlX+J+E2oYrMcEtRCNkUTEBLq3E3cucEIFdf3PN8cQqWJnmk+01KQgQSkifUIH+2L/9ApAEy3
NtEDuVXgg3avNEPTevRi12dzo2iI7lPW2hjNJd/TtA5DtsG8BtIouuXfQveyZ2yK77cmusEgOxGz
tls3PMA2P2FuxaZ7ETr5+YeigJJ9YcnpY8wnyVTSA4+v1Vuxjd+axrWspIeRXyQrk54gzQFss8Cc
iU3fWuzBFk5MNuOj5dg2Zk9iFLgf9GvPANyhy2JWdnVp3hqTEu9Xvdwtt5EAChMPEAw9ixi5msD6
cQnKI3yeWByVfcD0nTZuJHN8+yoZiqZgU44iROUeklziemjy8T4hH35n6EGi4ZOvQfx74PnkLlva
uNvN+m7MoXd1If/g8Tu5kXf04M5AfLUsMqpWTXKhqqjGGvynELi59W4XsqgwBVpDS7qCWnzd8BWj
ZfaTRpqg7DFSgKQVLPb//eQdyXDYPU9xqVFxJvL1wcT4KKN8SRGLoC5AtxtKWRf9JpoF07y8BAMH
hkBMVi/l2VkBKSRSXe/d7wpRtp1GV1ucj+dLHLIDDdyEV+SP/zx2KxqKTU4TOxjTZKulwGp05e/a
hI6sw5qEfsVdBC3pGynrpjLB40HNEyAUQ6QYKV8INgHrt7hHkDS3IL3KOp5hXkY4WQZh9tJx1ha0
kn8nJxyiOhdtvZx1tFA4lfkpxrTmE1zOzrmH7tuQnl36ZEiPtWArPt8BkTWPb6pW+YvUxCsA0bFS
xmioobdUJa1Ekb7cyGGz9w88gAZvgVC5uYPbkTQEDSsLgPcaUtoM1YAih5q234fZgolS19j1Ymgh
6GmTNikOI6oSGj8tjn9IcJYVgoe+AYKKpJDFj5/uu0stkYhkLXGFSwst+NxjDHo4BDr7Uk0vqYPi
j72nIc6Lo13ouqr8Y1kthjtsj+/T52gFRSlWJznQnvyAbyA+OfzZCRC8WPH3zt3+iefuTPxmq0jP
P0VJd0Dww5X9YgQ+kYzhUL+24iZQEfwFtL9BwRo3RBaU1smOQytgu+nZDDY/TvtD0RngxPz3nYiW
XiB+39bACOUgWMYM+SpFnsOR2YjbYY/9Q74I6pyeoO2Yi97u0A/JqcfCI1Nxtr00wfptgJNj7SMv
e0FyasNqMq6yDV9lrXaPdt//BsXMBgT7xqrqkgYixNYSK6SxdMxmNsrzW/ARyMeMbaYlPoblMBrF
i8nK/s1ZFeBAeFNhNto0N/aXEMjVyVAm6hDCjP77aDp4LO5eWelHHRmSpvG+Ztn3qriQyA8HplrF
PuA9sfqK8fbJdilqSqpbJuVnPO3Q3Jo1StAYjjHUqRzyrmlsfLCfDNt0wd7ymBja0+2UZQXeh559
sBm4zSTuOzuUA0O6WDlyL0Z1zHOvJPV68kXVBewZwVMIPgt8IcrZkbnYHf4pHTR4ytmyIW/5b8IP
uDD+rLhiCmUOC9nLELq0agCFiSqK8jN2mFWvxI5xHgzYrkps/TwN6oYA1EzVO7PR6WNPyr5J9xnD
MfG4jqlziQMBovmp7TAB2bHRIIa0h1iewqdtRPWrO2oFy8fjoJX1I73gZpdqZCZxpnjPPUTgm3Rr
Woa6kKTq7FufR1gGG5rp9K+pVdeLk1n75EtgZbhYfCWCuSPVDYfle8BLUD7Auc0dDeLI+vWz3tSH
D/SutSCry4JbPZXP42IRGq0V7dGDlxEvPuxJ529urcLB/B6tQpOYKDRvbFDGO6l+liGzsXZeME4w
BWzy6Ff1MnIZJhqNu06WtwzWud+lMv+vAsLx2y3IVqiBZQbsATk9KZiQozS+gkgyEbr+sHfIynOX
+bBmLoyR1yMWOBO0ZmRPdf5EfBA97prtl7X7qwKhI2oBMwLvC3Fqq3mOp9R9aBzv/ratUEwFUTPL
PqKDwd35WUegC0ITl4Hd8pBckDnzC4vQRVD/RfKuy7ke+lXKiCFiId+fwIxc382XmKaasDj3HFq8
k24E/2D3fpUK8p8+DbzZp7sk1j1kotEERS6xl9b/tGEBxtxaYoj2gfmKVHJZHPhhQ0QsA26Vdzqz
3SyNie6RdDxLcEX3wIw9FOuqRwDVP0RF9ZTbzgQ5bVyTFCtRhlhWNzulyrVKdfHanQW24O3sv3C7
+ptwLe4Q/kni1T0FkQuQL3+BX0BueOu74jeC/56Pp1VikSK+hRVzApH1bXsiw4AoSK7wF/RQi+6u
/4Kbum3hQ+DPk1u0ipvmKPpLghewq4YarZMyD8h7wL/uU8vpouW4STcbCy0mO2KzTiq88Cw/eCuL
jD4TSr1xwUlUWu3Vh/OzFJm/RGk5MESSQvgNDQ3vDX8kn57ICch81VDEKkeEF30pTm3HSkObTQSt
w1/W5srcXTtaHUa9yGxz9qmUCR7WtV1cQWEsiws4+6e1I+m68XxWudzvahr7RhD777RjxJrjE43O
qSQ+bImqonRnGGRjuSSItz85nXWsAGEdrSjlXIVvuqNctEWUd7NvId5+J7hF4iaZP1x1WFwFJz6T
hlJdpNEymubWu6TpqBWdSqwy4+bGsd8xgVSQdB8P4RaSlQ4L7LiXBC0XQlGV+nzCZs08F0qqq7gK
k3IGwAvd96wt5LtzLs1AIOcdNqW+iLda3jixw0hiSLVfe+DfbYjHrRtfWrL5u7TOWE1I22AAVPu/
TTBsOIkIHx9StfyLx+wvsopK/qwm/RdxXepa+f7Y9/FR5imssMQTUr79Bi6A6o98QHRD3SnOwBnH
fBwjOwrdOKShauJWAVj0uanTex+VohmQ1DtZmg3KElT8r2FLZ2+T6UywJ02ZFwGswpnUrLx93VFZ
qbdf5P78XnySBXE4aoDkIHRAfWTQLldscvKGTQCmrlkb9rL631woOkvEiThti5y1Z7HDlx6CvnKS
m7zcRgiLokzFXXMS73BPTLa0Aih0f9U0bPDG5q3ZZfjlX9UQIX921YdWKwPpG2qlUxJ4BGEOYHWI
WOVcc+RA3IlKmJlRqbwyHffnmhLCNCuqDjAggtwzA3Y/K+OAtphkWI8mE4ZOnJlJ6li1TrluDYRF
uZVBfWt4eEJS8rytn86/O9E0aZJOAuibyJjP5bMPhsQbyxPtmTCyL5w+bPIEPtEsc0JDaQxPkvoc
87FogYecYnmg+lg88nIQ5ED+lwbpC/jnWpnnpa4rotKrjexIuXe5XB8DyLKbKyHnNexo1rG92pJW
dHCb58woiaQKHkujHR9ybo4OY2cDmpuTaOcBVP1DYbQAxNdo6vlLgjLupzHsV1fFyGNQ72toSMgW
3RDFwt2yExQiKWhdWgUP2YHu9wPh02gCcl6qxpt5tW/rVISPQYOi9R+6T4OHCcWsPNk8amrHcVQx
42k5qzULFq7zBDa/uSI49L5sxP4pEzIza25kG8V5W2PpMveX4W//NGgTibvZnQOg1zj9UPrv+Tqp
TjyitNEr39UPzBeLwOUi7oAcwjmMTq3MDqHAoAtnHTv8Kd9pPNujw46ZfVo4RchVi+50Q1YojKhN
hrZTJWdnfdiG2tdBA1eKq0K4kL0cELE7ahLi13nI+Dj+ViwYwJ/tvy53cThfq73kAj/FzlvzIqIE
1Bk2t8ClTqevnU7X10FNEnSbgccJ26TYz+RZOiYwIEiako9kbff4ZJYoMyggJwvJKaWqzqsCzjdO
k3FARhuHheYz1RFFDVORuifiwkBDN63PgEdtRpsBlL3GASerC1pOGRT1Jyy9y89jixk77Zw5c0AO
s7dq8Fr50Y4CR/4yoOfa4oWsdOhTfA4D+s0YfEroI21wd0uI7juOKWXEC237OLwChqYVDaik/zdt
YRoyqg7Yia567xZ6kcsM7lQDgpqhsK2HINnnuCwOmkoeKhAzdp77Ev5x7dShfx5DGmgbPLK7+/n2
aNstUkIBlOqGASWCq9wN/fHkGYOJePtVpCXoEnTru+6QzyoEtBZnyudn9oGrgAK8gkjrtAwvEA9J
PEzOQw6ASASvh2bQQTXURfAzrhiKhvZGVM93Le9ssPFFAZ8GBqb1Yq+7/5rSNGfg6ej/NE7XLCDM
yfxdsN0XtrOpWjqM8pJXKsnroBxjOh5jf+GaN+tU0Rh2DEYZNvtvFGUcPMshitMHNLkYJuPk7MYH
sWakPLVEgESAgHAr+aezFEQ8R0hJqFdc6ri1FcYRFg/x1ExWrL2xGgRhv6WbxzqUjP/WuPIx++Fs
Kp7SdBwbPn42vxPwD/PzkHc+sZ9yS+7/5OaFgIlwvr+Z2SQZ1RSL/doJDrqxr9qB8ympvW3CgpdZ
XeR7xfqtOXyEUaTWcXo2tBpQEW15cw5DItJbOI6NUGbzoNLd2UlRoRgg2WzqX4BtgomqV23M9bnz
ODHkX4M0VTHV68UHnOS2xbrKVhSwb2TyxBFXTKryQ6LPopW/QHzV3Sy+WvMDK5Oi6uW7JhmzZ+Si
hFpa1pjsFEyROc/Vj1sdRJmBxzT0jSw4zKn83dQENeOO1yn2bQDrCO5WRdO5SH7XCR8IQkurCcSF
uRbP7gQAq9d1479ge64xX8X5lqPdQzx5+P8s3tcs2+nd34qJ6pJUCHQz+dmhlStOLVcdbTWhfs+s
ZAHeyAmlJB+IIW/KUHPcwaLCVSEfoCbObgs7P7bO1O3sx5CO9/mnQ3LLrMfy1Q49gQBWW4osdQzT
eL719cMtlKyrKKPjbWAkqhBxeNbvMQ6bIaxXawoVk4egvOEN7EGiinADOIE6rlONa9s5xqIHRZ0t
hdOZMK21dZRZN3LThgWoWqp6wFQuystxwae2sFT9HmTnve+8QuO4fMK0o1RuGhme+1WZvcKXKlP+
w2Xn/bWevoLGZv1FF+S4wL4qIOcnJPjOh5hOtULs2AC8SkeF1Dbv+yvqE9O23TLM1zBqw1W3/znB
V+h6b75Qhoz5M+IdZ/9hK2ujqgr9smiJveWXzwnvJivmY2qe0iyr68Xgt3kH+4/WAYRQAzpm8wVa
LINyEPoRtlNyea6S9YTtFWhQ6nr7C6rvOqshb9JtUbxsOToT4Jv3HQPaetVXp9mwYs0STAgJPwS4
WsRMHBCvvbxbVqNJ/CbwTWtHA9g928H9NB4Zn1cLYzUMMEJPjnurGKlipH5TzDTxLsCt4jdvbb/g
jksQ+YIAbT5n/LS1b1Sur4876p7AiE7NvWaYeYdRjPslhcnrv2cah9lzBGQNgj2OBHQ+LEp2srYU
8k3kXXqXKZr6Bw9RCDwKA9UcU7aBUso3/Bc9EEAApDaNqkTKZj3Uv733DTf2zqFl+fXSlM7R7opz
dq4kJiG66GXuhUU1gxwtSalMF7VmVCrkD7qlsdCiEI4ij54+tALPPIUT61BMGXCX6Bn3i5SllkAu
+F25DGW6UUunUzyL+4Flrn3ZUwnRkk1xXvquAAXWwdB63wKAFLgwYHtsgwQe8BKpI8Hceb4chGfs
JPPb0WBJHCP1OwNLCtbhECDa/wilQtllXvV5+T4tJa22p197tpIpJv+a8S/DTSGJaIkler+SLfvU
58PyrXe7NKlC719FSScpJL2FE0I6iTqa2X/O0xoSVYWztG/3N0esti+mDoKBBsk9+tz1/vPM99Zq
JlgD9gA9do3zIVqizfls+bodTJfODDEShQUToDGQc1Ag4f14HMmU/n8f+Uy4DhENwmZNHF4HPIIk
JBuJsCmGHMWoRXssQMe5o1NKx3DzpMay11ldk6h8eH+9gPqr4If/KnfCxB9Fh1mKoRDCuFFi0Pnc
eZ/tpD1b16U+nmy4nbTh1fjFmMliIvjEejfQdantc9jWdTbU8IBawlUtPnUUqcPKrmu96bbqyNIp
nIdHFzTyZfK5QDiZBMgzwin8RukjwQeyzIKL6zEKHPtPTFd5B8lUuZR6A6cMHDassZ1RmmvLcut8
eHkeEnl9qGUlSypXL1eh293UltMRYDK56bjTbWfY+bXpVH6Gh1p+HhsCHsNtKyOlxT26/mTOjYsc
FAw+6eDzTtK4IRzZZEBeTYtGQsdfDmHHOen8ezmr8bSXAphgCL0c6amdbpYwWP7dXfTlXkVNTPdW
g3RFS4Okiq8qanIiblDDT0W7TRjyaTOxu9G5pIuPebqDWaFfN9WGtohdcFEPMb+BLrLJAD4J+Dv+
82jwajq0RdnpudVohaGIV/yDMlGTxC9jWem9c9QoLntqQJzb4eFgOa8ZtSEl5PKDdn1HfXkqrxdM
vqE1X01vi0IQ7CxKI4O4ElFZkfsFwuMBDb6gkKkZcXqsMEBVYE0v9WXnc30fziefWPOnkyIz6bnl
TmsRhAYglEVJqsF8MTjG4AjPqOaOr7nq1OuUsBa7ghoepeqig+8qOW/ug7XTruHUqNEyyWfZUjb3
DUmhI8x8oDt2bMYZVTPeXAqcXKC25pV2+ZpdqqhuLbH1AaDZeUU1vsylKeYj25xtYxdohGL8EKwW
ZecdJATwIdNk20vYaLXq4ASBCbtdSBL7JVMS0ldsj06+WUhxwaIbBpHcyb4ELNJEx0fRloCR/7J3
Rv1++kirkbyz333gIKmI/ZSzpqfcc201HQzWB4PpFz05K+GgMzCHpNOURV1IHQjWf8L8e+lGa+ym
Cb/87wLZncL68+zFavttnBM/Rg+8HGLAVLEJqY/ruT2ptmjxpjrjhqmMd0IYKk02X8YHLx2k2mdZ
z8CMgTX8PsHkDwnrrY4SqiLlymm6PwxzcpyYAVcpS1GFEIgWX7hxKjwDMp51ciTIWVOKl9CuTxus
woO3Fr6RJNWsRMmtmwCntckf6f6qXZ9OmWSNzwZD2U8/oAstYmddueotS0lEC6T82W6a78Oqt22m
Xn5wwcB0BYSFHSW/i7rYbTR9CIM62OOJtfCmzNZe7NaAn7z4S4PaZndJHlxvlZIfaDEi/SvU+HX7
+iuNIRdalZ/zpGjm6jNW0PrnzwP/QL7mwMcOVuEEM0jSd7v4koZ71xMFKZpq4aZda1n7NKU1KOHL
Lcjgx7oHxl+snl96Fqlgq5wJqXRavhFzZYVUB37JdFHhn9iKNkUbRON75yxf609Cjv5UC4+GkiWC
oWf12pRqYticnfiP6wF4LGgOxPmxBQKYKQ25aSs25sIirOcem+q9jQZRw0rWc89ZkFyAG3ADNou/
tps9vIuQMG3pJbRFp/T3zyzLbbcym2t0P5Vy2DTE8VtF9Ey8TuhUg+M6lhhQNQKhUCJ4xxyVFNB8
7uQNorIiJSdoqxTZuAMNnoALI0Tw8ucJWZGeF3M23cX+Lc22LBpQct2fYLL1auaWWQk7ss5pajoj
0tMBIp6EU/Zr37R2Qzl4vRJSYJiz4v6VM42Q46A457Cpc8MJIXmGjlIO5zwTQU2lghsuxgNYEVSS
d8tTZ9zt+Qj6rM0fSMCL7yYpnKFNcXkUSD4FJXotbc6Rhx6wW5j5iMpzIbOLBZhJAGK0Ly+vQylL
Npfc2AlPMxBPP/XVtMhVvpT9nYQ6b2u3fH2RufmQik+fWbX3vsUQEZIyLbNwKAJ+6tOfU8VzPWJy
7lEB1KqsV9MDVzOXam0k8o6x11+HmagZgoSl2bRZGphqnlrKckAmUPYojqpfk13mLmjU2qASJjFb
Z89rUJCGB1cQ/bT03boj4JDwpljmJtvDyZi1ygm/EO16mLLmQ2hq4vD5XZz4+3BUdmfn1XaHRVxn
Yn7X0TT6XDw/qi/oxmziE0zQ86EFnPwLAZO3zweqbhgZXp5fQVBTN57+IL4z129Y5mdxvAUlKuN2
hDl6IotW7qXiIpZ8sE/BK1zw6mLiVwHMPDV36MOl2iQMn/e5PiejW8jvg9NcYCsqgTlxY52M1nbF
PvaVChTsS7a9E8dfHUcyRVBrPtiXCg295mryCbWlgZQnw58dTvkYJ8ai2lH5bmwkWDZ0WMbhqjI/
xqbyNKeVY5V/z3RzpMI4Gzg/S7VP+W1S6hT1udc5qnRgE8V0aHTheV9ypGuDDA3XhLfci+Tg2kFs
tpHeNjYyBfkFcsY6qH1Q5BZuUJ6GS9Ik+E3tl97HZsEEgnFMpfGRgwt2VlN1KVNvLcvD8vwlhTyu
tEfD/qi1rehFZns4LrKECE8UYU4lSbOLNCa6FaVtPOOd/+TIcxjiOiqt9d8sONOYj6BsFxqLGAgF
Nr2+iNrrtXA2AoWOfO0xwOi4WdQmY/wCx350mw0PpVmKWRxLy9Fb0CrrRaiHCTbrpVY7pJ5XrUlI
vAdRA9dg7GMkQ0ROLi2ncagOLENssb/qsBAiCI1Y3WQFTv717Xn+zdRnE62p1RRGR1sunJhLVmqo
mjmLg7D79DrO+jVO6E0NOHhOmSNiILODFya/p6xqpgExlTcKOpwjVd66Ke98iaFJW8hA4rrNLn1z
my2S/p/xUvUZjlFyYdZwZZPuIuZkHjgit+YAl+XdLKMQGJ2k4dYOJDlrX8f/aFz/nxukcQ6wuIs/
nj5yH/non8vkMowwPPNdEW6T4iRQS8btqRnrkADNO7J+9JiZaNePtNBj9lEBaEfA+aG2u6han3vp
+3Ob64hoptNDqj9rAtRRSUmqwRlMFMDErQTCrC6yuvTfLDNbEM3GlC3fRznHB61Mk5AvgXZQg2Ov
7ijiQh14bty7VLtq32Is0AEmB/ehfVSbXn1OvZ1zriBMP7K6ATZVxpRx1CqSzGeMa721ink2TpAt
qx1SebHBIqEqBv4X3K8p4DFkQeYNYtrGgH/8SpGwL+f9/R29zQzh/uDUxovmH83ZbkVRMyJIINlk
pe5Da70pz8VVUdynJ/2v4rYsZEOQ70ISkMGqVqoOayPhVcXLyxmXLn5l5s35jCTPC1UL9HBQdbG1
y5ZRaTrqOrDl328C+4l/3ajfx31o+Hp11IPBg+d5nrP+w7ao8O2ckPun6HlD/QEVoIYuiCcD/kv+
O6tuhQfotoqei+W2/vET0Xwstg7pMY/jIe+eT5UzSeHVRiXjIuPa4tE/Okkl3eZ2U4bL0eAOFzto
8W3cpgTDynII0yce93OlacPbeCIfghxCotDqWoTOK/JFlWaX6vi3a22dvhM9NOQ32cfCfRvHekHY
wpWp8Ic66xyVsATbfGgJ+xmAgOoIGL46gg8zSsHtMxxLiHUnVnxgBV+i6G6CebP9e1/DtV9e/cx7
1u8h8uLU9s6kZlRrqLBi/b8+/TRYZUaeqmUofruPuwq2i8DmdtiDRYYrgXJx/THVVDKRyH4buQKs
meAJdla52/g0lHttcRC5Cni1Zv8lc37V6WF20aTHbeM2yIYmUt5FjPXiEDHmBQ7DToY14eFA79Bm
LtHmIIuCbuyKgXwzXEBMbK2ev2QRWXNdjyL9BOFtoEHFWw0KzXcoPZurfiKyAxu1jqlGrWd7PEDe
kSnaBpDtJMNpdYi+xUn53XFLfR7t3n16AwUqi9wHlyEqYMpSidtkVZRtDIMjuarmVSov0E5hb+IW
v4OJ20Iqo2OJ6YinZMDLwaRHI6mQ4vKi7T1zuT9PTOr/i0oVeJgfJW2wlTt5DoX1HQW5+PpDp4IV
eX7Ooxra2tytwCfUx4YaoQWfcrzgPkRL2Tyvhv3OhEpgtDxBYn01cNLQmF07FH02TaBWxIBCttOu
ZE6M53p0aeTJxiJ+IwMcm7DkCJvab45g1nrD8iUGbYCH9mJIxWM4lAnAb5u9zE161wUXgHrwGq5v
w1xjRo9CP7JBbWggssG7vRJR1HdFk8a84vMbNC8y0VCcu8cHYLTlkePxOrWGrAUycjXkF/mgTPC4
zQRj4CGaQYTEBQUb9DQvgs4FX8xQcm4btSNHGRijmGEZNxXE5uGMkxXC/ZuPrXVk16HOCAozvbxL
+EKVmefy77XKAz6ipzk+kC71pznlTdxcA3qVIjiYVrkgVtJSkoV9+HD836/EPpsN1BlM/Izgc3L6
ZebTVBFP9bONgwfzZtcHr72+ss6aBavkkE55Pi+yqlAskqzkIVtrtkgQDrpTiHyEGu+ZDEa8Dwqh
fHOFgKyt4c9stC3y/qAo5HYMfVR9LXsacmxJO6ikBXeFfFxB/dIC+7IAw1T13x1lPnbVJxfkUKrq
cp9iaPNMwOpRcWlyamnx3qtUA48ckQVN6Cltd9j+gC7D+ljBED5KO9fZEwkdk4LlgY04mBfgnoxN
bION74uswUPqqXG/TSvDsuJsQgZr3THQv/uAeWvHpRj390hbjG7eDIk3787exsAchlACkmSiPgCT
9IHX12utZ3rLB839PqSeiLPiU+69YxomcHQ3tvTq5tH0NGPHQaRLp77GqsCcx2Hocstxko1HI9hc
puQGgzp8oYVTrFcyNPsn10thewAsYc4aqCzSeXY52vv801tMv4NhdmGqRGEruHR2iWFJ7XG/lit7
WvfRF5OsNaFDSBjviIt5f0WnUBIOB4kv5RIw/2vVYW30lz2/vOz5GTzGa1pK8hSpHXPvZ0Q/p79C
pOsGIN7qBoP6PDZ1pcs1fsARullBaprVMvPHCZcqCuAQnt5y+mlkNgn81UKPC9RIajQhzNuFzbJy
tpBN1WJ79EFKAzfF1CPQ3f7xJ3n+nEDbPfcjY4k5yhXNP6PwQxRNmQeei9uq+L3gyHiOpwzoC2wS
ZEx4o39yXQtLrPm3zFMiHTT2zHPasfSTu6WWz3y7wk45r50Arcce/vOFVDLOssgu70gfnBIS628O
csOmNHAocLs8s5UbptkFO5C+mThOHTFwfggs29t7sTzw0BdaCwRsOv5e598lddzTjKa8niJLdP+G
UjDBgUsWW/7lfiG0+SNoqujAF03YygLJwNCglPalfEgNSC7C4TIZh1PtouVnAxscz0jrjkgDwvc+
PtrYGQ5kKLi5CWNUoU6ymkKKbYUe7BJRrb6lF6J10tVrnmbLU5Hp3S/q+fuaPswDoOd9WMoQXkCb
NY7SdnXnCAvBaLffqk3vWnRrm0Y7ddM3/iV8oP0aGrwj3/SVCoWsIAyRGHkFGV3YiqYet99fA7Ic
a4wMADoHJA9vqskIULYlN0JYvsMhukxv/lY9pJvxV+N74Ue6HDeTy86xQgiQ2F7TDBGm+6E/RmLX
UAnY05UPDAbB3gDROm6mv7PtjhOPzqqoymLXF8+h6fYT3g4/eVpB7PVmp8sKhhL4YON8/0gux+MJ
2eCLPGYL7zQhF18pl1n19m36CUycyYhIQyA5fj8UeClOwaZ0umyE93rhKo+kpINI29nrToB383mj
6ipl1/IgHR8VMK/KVi1+j4vWVv3WvWYyELRnW6l4IuzBt1A/bQRF2EljQCIzapkRht6Ldsip6Y3O
CfeYsBH1WXnw5pcPzHOrM30VhGNyS0ITLkS7FIqMTdfGwkx6fLxNrzNTvVOfPxpBLKs0naIadckh
vmiOyR1pwNoPL1hkMAi9M2xMEsYtHkGboTDZhKX7dpQ3z4yr4oM8MhGe+l4ayT9m4IQGTwJnORoJ
M5l1ttnCEX9zs4kK8W+OhMyUvH5kS+FinjbekGSRqs9jjoLbhFg4g8h25sMHjc617w5cqihNXOrs
+ENx6Ax9w8uvX3BoLXDWNXFjceGcg+0gAVB0zJXC56PWNPZzAHZF45Fwpi4dd1Wgng2HRituo7MU
hk9Fz83bmTIxlTkjooqA7/71snfXSCP7OaVFhzxpRgO+q8IySQmIFXRaMV388KSZmEZHtRTUw3ub
YHYa9B2mK4ZhWqWr6jx1E2zzKzl1ysqVQBS3MdWgjFa87Ii4ATsOqRvp1RKyvYI0Xav8XOz9bYzS
D6aswnpzawE4IJlTYlkOyGR2XQpznNgL5vFjaYl2x1KITvuZciro5vUhOg9rx2MuYgafLtT7yroF
6jl1LbxdCTYs741A+raw9PCpJUJH9f9+Dkpv5CkeGByoHro0VfTt4u01xpl1BvYmaZMFy5AAbXbY
C90CmmOlfIFLNACA33XTve2MMjYUE9IKK7ULlHX+64uZ6bLQe+f3oDjK+y33jSto+FvbP+NAkheo
FWFV6Oo4veGltYVfiynn9SWkXr5rq+EQY1wH0/W//XXRhKrLKPr6XQRUNWPO8P44jwIGfcnXs8J6
vYq7fEwRiaBp3H3o14U9oQ92RN6Qvfb+ONbt/jclLkU4JzOZKXuc+nicEEYH+rr7daRlgDIoJM4D
axXZNRCJi1k+D10/8VtVo+VsnPFkKH+YKTmgDcQ7og7+0wBHYscEB40jqjpjyE0zNyZzJ4sOnPay
12nYzwAF5QPRk8QT5Yc+kixVVfo66UaqBU9cq1Sabb7WkICMeUabFPHjL1uWT0hwlRY3sZWfgYdQ
tdpf/y6uaANcwjpTpp6l0HjHq+rtBcPt0FDPC5VXO3uvh1HKPS46JsId8qgWG7QdCIrBbKYttKAz
til1CfZLrqVHmvsWwTszTQlJQeIyPnpR4x70HEhulPhhbtO08YLsZ06DvU8U+O6TwH0MLTxR762J
AaYIsGjG5jCr886lgMuZj55fNgHuX1fc8FHUPtKd6jqPnqHGSu87s7f+QUoGlu+6kJhV3pQea5Yj
IqR0+bTeEsM7wUOMhiwd+ZRac2EaDPG5OYSUYjSei9Z/3cg78qwXoBW8EsASfqOXPV1CvArJToDP
r7ldG1IfjLpjPu3I/JZMLbWDtyGd/p/sMXJj9OuJzQWOBse/sOg5OozREBTfRlOaZTk4xCoSHfaS
p5v/ml8WCKaq/xaNj5aRJ8bmAQyilrHfyjn9b62eTZ0LCffud8ub2CXL2P+/mnFNqUuo6DoZlFv/
j236p/0/o8H9jL0w7JW9keTQ5+P4/vZWQhrkDUOhe35wjbGCU4KZ8lql1R6lNz9Is/Mb3sQpaWnN
RmBii9qlFu3AvwxlLHqRAu0brvAQzDKqPxCDWqpeFJsvLOfp2ktpjN+oLKwd/1LhdrfPmvHQ6oda
EthrVnOpCEbqnpKirXc13y/GTMQw7M2Nh/OWancld1wfiHLo0QfHMJMWwJRMY992cwaRpTz8E3DN
EJm1K9YfCDyXQDsMvXFrZD+TkZ11+sG/Kn6f69MZf4F8nT3tSBdJn03KvaUYzn6gORUuDQ4uw/yF
KmuDfR3DrsAKuZod/BL4WDwMcJ0fYq1tN3/kVrhVAqm+sX/piLP/OQYwc2+hf/Uvmho4vhJcoiVQ
hUG20dZLlZ3SEHmYhm/zCEg1C2h2w6YqDJ9nd5C0RyeCwzgg92EAhNpxDWFY3sQdCT+VHnbw7Btm
Alja6Ar8NM5QZ5MJgpUez6W3AqXC7RgFQV0TwtzLpK8l4j0BQi2Rxdz2T8kGMf64QMeIth/PhbtT
dFnikR0BXzHefwjW62y1BFWLZV9hjhoKIVeHRrRhzA1AuEPfV5Yd9TBXLzptL6rQAKeEba/ylqYX
ju2eF1h0o9nXz9E+szLTlJJiKFS2daRg1vgcClDbiLlZ7mbkWhTPxI/6S9UNqTrkcNWLJjqY0tSd
2XTv8jyn9EiyXbvLAilOrbm97VDonwi6yLpuIHTxzl9vK2Fyd5M5dmJgTHI2fEuDXPBW3c7yyMbx
mVQ+QzLoRpQ9BoX0Dcptp+HfV3ZTF+HyPNK+kY1vfX1BE4UJguTlhnE1VS7otLNeIMrdkW7efGn4
7CTNO4sbjQyt2faIx0tNb1MLMLTzxs7TKUdDA80r2uMGfTmtx1V9BzyAL3RKsYLChzPfvefK95OO
QVvkyB64D8RJsbTuzH2WLHLNnbflXuT053e1aaAYPUDVfWoldbopx1XshEusem7Dz4ODntFdBPzM
0898YrSfvxrUneSXNpD0iLWPafM77kaC2uCuLwxJ7qxkHZF/E4D2U0+qS78w3rqLhbY/uMG48j2A
Q659aUF9eDe6hxUAu6fsI1/Dq7dcFTFDf9N0F1czIHMJIuurmwDcXyHDCSeudg+F6ZjqkTxKCupl
ozSN6X9Je4uieKyNj2fI7ZA/4cTRCqOL5+9sHFDdo+6elZEq9pca8dOSvuwMv3ZafmGApRfAu61g
ZttQa3SPfAR8rlnSrR8QnrzufqRB0NQ/9RQEwpHBjjir1BsavOwpB6uVH83bG+HnKu6CZnOLt7uI
ECLt2KIb6l11Np4QdQgYCvTEIRjqbd2OS9Q7p3K0Sul6eTakSwOq7HEQYF7nkrvkEDtCFcoANoAt
pY4Svr8M3CyrSViJ4HPaUzxRajc0LlWoYIKggg3mxuDj25Md1Xp0lLK0WsYNtTEnmHBEi0qrAiGb
+xD1NX+vxZumjSpzNaNgUmvbbT2YdxbKG1xfOdItA99MfHCMjd2ciDcrDfjsGq7xIHxNcKIGlFeo
HvVMWPdIQXv1sQRBngmif/aJ1j4OgOs62y/zzzFGFLsUSFSxPgmoL4pBjTNFuT2dn1zAEZOU1Lp2
S7g+Ch/Wm+F2vOeK/FBD+kgSX9XWwolWYL6XEnNaECDOg0ie/xlm4/QyjI6NEb5CYnSYMPPEj3+N
++7MwcJQDq7E3RQSZSgEmZAweUQ/94vFgD38+Wi9n8Ud1KhHhfr5VJgQla72waqDUsesySrtKFlp
VZrvilwOyxnB2p8VfAKhuOKZMxbugF7TaS8/0mC3vo7U3FeUbZiRC3CE43cVRySSIS4Bb+X47Yw0
ClxrjmJpl/nQUY93CEReQcYQPQjU82vEd1Smvnv3er9ZLnp/xgO7LV/ob4It6s2y3BbTjucMHaGw
XTf96SQl+1zBL5ziVy1zm4/47CsRs9oPNhgXYIix68ke9AROhAIUZJKID4fgx1J3BD++QzkPOchW
0bLTfc/NknoMrl29nD1OI2wVqz7q26TGotLbi9aCbxfkSK8oe7HPGhIwGT8IF+Jo4Eo6PHnmxjg6
tgmEd8GiZ6MreXOwKmgarFb+XVEakRUnx4ovTFXth3atyua9q1Za/V6HF6ywhcE5sZ0JgFU29LWI
EXEA7FRKBoOAQ7HYra8bobSmb7dvFu0XzdzQgdROpbmoiUbZ+nXh9EVTpnbADZLjEBxKd4CSNJoT
ff5PShX9cakRZHb0hWlliAWiyYVxXlGOGBFziwYAdUu2rzzO55s/yM1owmwGXNUX/usFem6YCrVd
A/Yhn0gWU/fL9EEPRzhFm+4DJy004P7fqgxI62nr1caZZc49hnDxMS681SgY4eb+RRbcj283p4X4
ICLtNSmdYnHXYL/3pFDmlH7QKcExHgKwFZWHgLMH/SHtwtwxzIjaf8RrcNDPhj49+ez01IaCHxwD
S5HI5sG1V41UZ5XMnls7IN3vDEm9rX2Qa+MAaF/NHLn+cuQ79S2APcz7lHWKZj5XxwmEJ4we02NN
kRT5gPQHS/RpGQgucJlyq+5vyC2/ByoTYu2jckOvsm4n8Pft76iwX5wmtuAmg7vY1aYfwD4yvcDE
/6IgQG18XWthGNtcQowL4taTtSudUv7IAB2+EgsSyMGfew8I2hswQ1DD/rV72nZINwSDUUv4McUN
BbtrQP138t7o496Pw/g79Rx0t8N9f7cm8ggsewg77BG2Urre0/8+5jT9wZM2He4FfnjTW02xcnRm
6O1N10L1Z40ZkO3BG1s6MnRvqb63+xanvEtnvc4+v8SJJRg+FPJxdZNCbgY19Y9gurHLAn0u0YBV
5Gfm01GQK84JM72PO0742dIS8n2x1P9+jriMF/CFYZqeEJiNQcvIWEBjd/HN3XB8Yw5F7GYHE3cI
mVQIqKg4AaJzZbuwRH5tBI8VRHUmD0o22vhZ8Ni5AjPMVzJZ71V5ThLheZEE72A9bd8VeE5+OZUf
fKMVFOjbgTrWuFMORKEOSwZrBO0z1Qm+mVOP0KxCS2xKNhogUt75PdwN3pc/nKigEeye4DVy8skn
YxbrX7P5q5pNoR7GfFMXc7KNShzG6o/+6M6t53Yh0a/YGa/0h33DZ+IH9tFotX+T8MFZqJH2pYOY
b6gdbVucQK7+WzA0ga/Lw8tSuEPCDIbEG6/9j9HnQ/x+XMBdVe+uxRdZzkXdaaIkLB6Em3eG2uU4
Wp34oL3cDEemsVPV4sY0DZSDTtqzKzIbyVCdUHcPPXhm7oWYtrySqA/3fEtsfLyTQWh1ZvJAa3jF
AKzID6EC/W9q674vsjzz8g4D+OVWYXuTRIwhD61XGhtnGcvekW68+hlv8zjJ3LIRrlrvuWl4eUoJ
udi1fijY3wr4bJGv5zi7En4kFhZwv2IZkRAKKqNoumBleDrCUIl9Fr13XSqIDGNxdRrgriWwYsOR
WfahqtBYxe/qSHn5uETSTfBHLXfUn7/NzD1CNvTfEASIv81nOwvJ0/42iU+LA7R9cIuSlw9YVxDJ
gMXL6La3QxmcM/ocAEmpeBI6LlJoyoNcUFb4PvWOhOHymlztv8f0Ma+zHouxjG0142rMbRT3rjOm
mdkwgqZ7LdQJpcWxjhhQhJ22j4LMS+j5gVXsFxx9m9WoG9x4cEJkPYOMBTI0wr9bjOKUHEW+7r5l
Zd5I/5rpdLoD5WkivSIr8NN3tWpTzwwTxHe+vYJoO7Q6Ll4Me9AJmcFy91Q87guIBtS9easKaJI3
vSeg8VUFyHDN8OxvULHQ5VObw9hqeQAOB7PgErpBlI3GZlXR+MMB3/PbsZAqGXiVH0WT4LGmEkne
c+qpGC1sK2WdVG9CIuvwz0PVMNUOXpDbc/Zo4BdOEHFdZvFNYozge1zjxSiGgX0nUBV1nY/c4+VX
p9MWDcPippd+FKf1zOij2E4Z1+ePFwg7IM956uYFg794FrZO52UF+Md6xMWwXt26JI07W62SAfwV
R2xgcU+6vOO6X+NEZQ9lyfUBDzFq6ipIFoLwfe4zsQqofnv7cLRG/05cLyi6LPeOL38Qr/d/c42p
xvn0cy69UQMxXfKmi01ZRQgJLGRy5Mqmx7hreLOVYPuncxWURHW7Kan6jC57z0BjO8FscmvA3wRi
JAwIlmp5DJcvPj30cxA0jZ3UTNgzw/EDpGOsAodM3jNhpNx1nKgqiMIWFOzOFKUH50SKahe+Oq27
zXVWVQcMklhdewtuPOvAKIcZBSFf0XCioV1hkzd4z6wRLIMEYwV9PootB4R3nYogplj07UDHTv+I
F/PjEnw3pxQdB+naeoa7b63+Irgf3JiNz7X8JiT6duxkNayyfufCZGBP54iYbuZbAcR/gjPMl26Z
nBnptMF4KMgpbNlELlp42JpWh/+hZRcET6XTgtzlqMnMRN+cZCk4sK5ee9AH0lIziPzZCWLo/Nn4
OQZ1OktAL9BKngJKrNYPeSKXbaalFklvHX95CNh9vSR0XmUIR+T/DGNk8HyghDxcGa+OOfAecnCk
FaRSb5js3bCIqrt1zhwjMIayDVGACo/8iFPg886aseBXjBt627KaAVdJrKNthW46HMAYCUgBYWjd
dql8V4K+shIf3+k/YOaHFtcJmuv/DWzPlVkEI7UI0i5MwSdXrASlxbbOW7pajAQ45pzlwJ1d0RyH
GbP7wl7WBOU3yO+S0v2uSBwAzlOuxQeYePgGIZd3umu53MrHszaJbTX257dFqj93QPje82zc4giy
xnM6yDcS/boROSYOVtVSzAVGe8R6GZQMSDz77HUOI+dyVLAk4ZmiT7WZZ6d5ilpNgybJS3ZGFRnt
Hir7HP4rmYGpHdzORsMUoRbuV4PGaUwNyqiEIsQ8Alledp0h5QBzgCm0WmWiT8fQY+QHqcQPFkZt
uwb2L9jj6jOXrtEla7tMgiXZYeKi6XqHqx1a/ZQQrOtoXLGOt2MEwpWuH2F+RMetEAZNGo2hD4sx
eiWjJZL4I7SS9XhZWsEJ+YIQVSBJfedQNh52TXsskBRXmqklnM/NhQ68K60m7ZAWt322+kvPDisy
sLGC9YM7u++k1rHltddwi60Dxo17i1AJ3VopiZ8tVK41Oh5T/cpIAH4VrsCTg3J1+OmKNR4wAWEd
pe4K1vIaQayieNs+a8eTRjtimSA7sM0tFgr5+46pio0I+aMO1d8cLsQuC81ly1HQBw+fzlY4ZCDy
cb49DhE0ZK3r8dzaLsdAQFLE6Lh1uU8tfjhZCLFwa1n0LSMbG/SoAl5JrA8sEBRs2k0gl3FY7PGi
2s5yqP6IDge/CUc1HmO5jfyxTTGBIhChQsGloZJO63PyYF7hXNicTvsAruOXScjHKMZ6p5SCKhbQ
7RlFxJi19XublfZ+lpIkbJqe47Vef5XK33gLbQ2CaPMVyq8zf+leILet3R15CfJgSWmE6uf4P6fU
9RuE9dXrRHnIEcySJHXdScjA6CcjWIQMdNZ3+lsoREI5QVvfi+LAP5TmjlRLu3AKWcD3jRMiltbA
pRGmbJFJpXySz/liqCzmmkHZZ1vA2sEwhqNn5crGFX5xxF43DY3TosDVsYKpCb0Gj/XeczFKi6rx
netfTps3/yte08ir/gqQzxTNapFa709/frKthiHlBJJQ3lecIyhxpIOH7Vw8xBvug4WIHta4270T
7QZHrv17oTMZQFlFMzLB/SRNzuBHt0+Zpeybrye6waUrDX6DE7P4q8SaiRT5Gew0xDYlCo93MmU6
LMCcVdIcelm8YzAPOazdY2Fx+ZBXTETMd80tSCJizKJkY49U+gtr+3hHpwk8kBNeCIuk18pETosk
MQc4pIJxte4shw6/cNDhRhL5K1xsoor6yZg0n3u/7Zfla64dRa2CUFGQuSAKKc3iJD8X5As0D1vj
Irklm++Tn/uH4sEvPV0qbRZAm3+NC991vyrM+QHxI7NCjBLC2ppNaPep+e9rxYxG5Mr3moyF/e5I
DS8vIR7eBp3VZweqamGOqEKCX+pViefzU2u88CtRE7n7aXdfWZ7ahJtK5Sy8HmSuPX+Cz+kb8h9w
3EsOrQFnKTyYp89zXR2Pw6hAawWVMsTd2jVfrLpWghYQgi6hmk9rFFjiN/7E4GArYmHhtUs7g8e/
lbzOWjUl3gd+/8GfQC4gPZ6yWvfcab9E1O9QHS3g/WTkCg349X/vie0DxZAlpGzzjQV0F7bo0MVX
GTlQME9PsRrnIaA8YzesuOcCkQT0P20kMckGz+5VImn+r5EfY1mouPctUq7fTTXdMlfkCQhsQCB2
dvMTmnHhVexA3Qsl5WlSgxUfX86IEsSgi4LNpx13zf8Amf3Zz9rVCUvOfwqxd/HNUyHLE9VzneE+
gP3su8ALjOkvcLdOoII6ktDndAsiJTvwA6j4rMQmSDD1wdwEBw4S+4NSbuK81BRT/hxWHT/g70MZ
ze1PJZv4E195o5mYxVIPsXKbBaa9011MRwlSnpQIYuUb4DNYhALvd51mmdatmNn1UmfTG6eAlmyj
T/iJbXwpmzDnLP5OA73ADH7ApnvB+4tVW4jAtJIwCyZ5HfI0zoVRT9JaDM3lmlOvboft8JBRhLeE
qtLFBPxIz1rDoF3XvTmdSgWHm+3U0CHssd7/DUma8hq5B2qd8QbEoC/NEC3dw3LKRZduldGl+7gG
kT32SoA/+L3U+nwTZWNJWojfP11F+jlbYPRDY8LLIPtxZeuyy+Ur2k58v/mHvSVT4I2/n25pNgdZ
qoY/lOdPQrns2PgNIDfBZnjgiWZJ5yuQDQ0DnNjWS2cNcQloDUz7IlVga6C/d9R0TNPoMv0yiF2D
xxfZH+buh14CeOljwG7kqTCcYZygFsUWbZsZ+e8rSeHLuWISoTxPBl62xw8O37ipl9Ee17oRyw2V
CMXfi8jxHQN4TQj02M0EAkzgOEkJjBen8jD7SUcSQ19WZ93JDiOsI1PF47nMrfjVGtHycHlfc14r
0tAq17uv+ZF2/ehZ50IozRgtBFHzONM/x/uEckvaA4+EzdCVwSD6ScY41717y6KZ3p2TQTiutOux
qDzau5cEZ0+Hko+KjPSLgU31cdZzJsh8ue1qEmm0dVjl9g3Xzi3bjgOwv9SYbkW5demGPHglOFR0
lkDEaqArLGYwGwCLy0jKvCNsWxcwsAtnprJspJog5M9+ScvWv1xXl+oCdKJ135RXzT8f/jBFXnBF
TSY35s3ngrsZHdM6d6arVBdg51nUzKn5K7MFwO3tddqumOapSXkOTP+N1A2ryA0oX1ydDp2CvQP8
CG/rI/swIsK++vN6p/CmSi82frxOKbU1GuuaFWG4qx+OZLao3/s9/vf3khIZwS8+BvCBimeTAun5
JKPRp2/aC8LoEAS/c2dARcDP/qcsJyOHiJVzxzKh4yLvmcki6N27xl2LHZ9jObNQqvd+JiL9yrt4
1CINpOlPN2DJB8nqYrMOuYO9uKyWoehDGCqTqUubLgF/nPeOWb8dIU+chwjfCtBJ5n/3NCdJfqck
oSNMdhG+eSRtddkO8QlaJJH1oRuEaU19otmp5LiEEITEN6p3nLYxxj2jfOT9Xl4luPmWQzZp6WP3
vH1iIoJwz+J8sHyziKU2GAAiq+SEctI8t7+ogzlTCF4rZqAn/iE+7wkI1sjbSn8wePB6ETv2e0fv
xgz6mD3McBFieZXkKWvbAg+biB2DEyitKwWS/pK/M2gY4yFc4nTp8VJgZ7BtTbWZRuD2i66PLNMW
BS8Xss9E6aBp3Zg/RnNajZI2XCjovaXXZJO0eejHPmYFCMAMapQnhIyyC653dPlaUkW/Av+URZ3d
+0zMBntO2uEbC5KMZPujIlTJ9pP51bk4SOKTxIPTs+d86QLZWGiL9m9tzACkBKQWIf2+PzvS07B3
hNMQHWWiLu8G7odoFYoC6wDhaRg2OJlPRao7GImPu9AfK2z/Wj0SHQ/5o9CGxAy81sIDLd5ABZY1
F1phelbGnTiU13bZiC77CZ3LDh6C1Dfi4QyxVZtsN6EAHyocCyBSQgQBoxobmbdIEsH45LHks5l4
hwwhS1R2RQLHcM85f+odoY7PhxJpJIcpClYzRIUZ4fEjx57l0mtqapfvVTfZFHpUTkuxoF1rmxEJ
onyl5njjMdYncTwYg+kOOZ10eZJkMIQOI/GYL1mfGV53u8kqI0VFnjI5QFyLtld/tpdRg3Cv2jvN
ZjjgfSBYplrqoT0OaSfiqAQh25FH7EB4WbDGXOrFYXG1JCHanLAzOwy+nw1xpHY0CZMzUl7/zkAV
Aib0lAmfH4KYqzxrf8WG+myhyVE7SG9YXZWYPeaclXMgrvXw2CHKTm6MXhc9jeD/AiR7HRRy5XJB
an5cAcSHpXltrDyHhWFEEo+m3/RSUVkJo9M0EHLZKJmB7vAACREkAR4ksrCT6zu8nWC/LY+Qjul5
hboE3327tuWTsQCaSbHS2wiomDj2ANIouYEl8fiBKNf6nLvXWVNzmRCkwoWnmuOh++3xV3uFvkeY
+D88qs8IwJ3DPmOs9NvubNeqYTC0xP0zfnctgDI1I9gDLOooWatDUlm2pcHc4K/xK+V+Ym+aYNfY
wWFpcicXZDzm+8WF3FMj2g6VHEOvhdSLyQBF3yfSlDzjnSJDENi+KnZyVjzgrXF2nNlXEumZRayN
X2QGRPQrzrGKzP5FJME0d0A8biNSNx6dEWLbc9Mkd677zQqYqaFJLKshkAS+kf0ZFuJAgeBXbQP+
zWvV8jLorIZjs1IpY8ZfKraw7LiELoOth+luC1vSrLwpxK5vH/2QMJRLL4cFLp16x6DR+W+3mBWj
3qfeICifeNFSk6DTeUhbqWZom5NnIuKCYRXLb62uEMPRWqfGWAsxEXtYbBOZ4PC2bZNqKhS6Puqv
Noc+U4MC0moS23cUGIw5rgrpoQivWvwoiabVbHfZIu0rxNG81ZZCML6GWzsBNhESdXOaBMaP+oRF
jnrRwZ6bkof8RCQhVx9cNnyoW21r6N9dWogtfT14DAt8ieFvLH8Bu8V0XL/hTCzDtfY/R2glUSOw
y8ktq7flZk/7EJ06C2xHLYOlW2FE1Xi9DTHr8Bi5hCIi9R9PZcqxKxAyHs8BXBoON9aHL1Nv/9A+
6QLjhnn95Qyvrlr5vr84qkoe4FBdftIri4RrEqJf8u8UJnDBNh+HgOZOGseeDse7ZIexop+OMFqB
BXaXQuU1tpHXvFLbxQ/T7pBbIaFwOB1EgD9GnCB3EnqomBlzAxd2+3vzPQlCBYu0w37K2nASWhGl
TQDZ2lO3FarWOl5prd1oo0DsjhJ/SSdxu7rdyZzfEfLhO4e/+21IsNpFyYswlfSMjVVwfW+Et7dr
jEPQUKzv42ngHTLGprL/Ig8NqOgxatjexwupBlayNo9GzDxvLZSJgTVfDnASqrzIQw6uwwCvJNoA
JmLuXm9+Lj1RM8/XnNKArKT3UOlo4FjTD2CjRmBW1g/YIkdGzF+BKvHa3uIxpFrS2HxtrNNsy/40
HJ1eyL0uKdFEo57zX/nGE5g3eRDJYaWj45vbl2f3nsARW3K3eZSyw1RQ3KDKwVzNGomGxXrUDpFN
phx4l6JqK6OV+3mnumkG9bCO+9iAb9W30D7/1vyk1QdhqjGpCxmNN0Vjzez8kWBHnXOQa/Le5/jS
yvXt17wuqgBHF5q9X0+Ip1i4VqbUDCIxm+Z725NBrVyKaBDgukgHYkw2xEflxzWJfs480wc4dkoZ
ek6bZfiYBkUAK1cbICIjvSOPCnfHZeP9KfQhS76DUbTqV7DNyfJ2mJhd0FgAqoIVS4sQRIiSI4MZ
cqcg5VmokGJgJHCkYbiYuEayqUEjf0XqWGPYIoAQv2mjibDqdMooRouL/fzYY2jTIhvqcChhtVVZ
8Ndx2FEMv7ontKyH8I0b9n6pYiesq9WnzPGxRoZIi5O7y2ybEmczVFB6ABjtzbhfxcJb94jiHn/4
Ed51ysyc1WxvSncf1vIZ8OwBl4eQU9f1LQ6JNVOAMTCM90iZg5cS7AuSHymXzQ+pOp1zTZTgacx2
I0TpnaVSryb0kkLF+HpOUAk9EGKlQVMkg7+AqXtZZzJ9YpjQx6lyZ1U6ZOxGWg2aoBXyO8KkAPZO
YK4bJNlMe1TYmIqWREiaSRYK+bthTpgWk2tN0mybVykTYJ2Ff5uVAycgUVsdp0LzxKJyceBodnOD
RkD0HZ+phO1l86Hk9zCKA8ilLZ20fQFgYnIcTf6CzOrRCMjEpNHkHwPR1Mq3sC0JFh3EuaG2srNB
vcaHp63H2+VcICSj9farzFFPHjULqrPB4yZdMD9BYWGcmOMNCr0CRDOqsp34TUoRBsVMgevaynWC
6CWeJoR4QEZ7JFqD2m0sW+YJQACPY1oyhBYfj0fAJxiTCt8sqXBlgpDhBrqyBtNU8jBWC8KQC+AU
vGNnzP3x1/X3VOAFZD90imv2+P7kLMNtAQQVn1GWQMABisveZi5Ik9laboB0SOJYlUpszlvecPBC
bdN+SbYJrfbzgZKPmstirjDUpn0ZshFcr29wDf3yd9YF85oJHTu4g3Xtz9/ptTMaleTmiP/FMuOe
rayPbP1pTeU9wJm6RhGw6GEbV+sd50B3SkPShl61YyDPOiY4fl3PEJQW/6tH4KBoNbv3jsFQu3ic
0/hfASQJn0hHD/E/WbmkVDZoGbynhIJ1mP4bYm/Oa3EO3HJPA9JxcYVspV3Lm8s/iXLMIFAyhGpH
blc9j6lC+5q7q4YntKPlOzKh0o8VMHCAG9Mdi/RuMiOlQoFbKfMuP4P0Ki3nrSdgT8M3QJliIK7L
tCBja7c9TDl7mQxi5Q6LCH1OJ2ApzwVRecIdl0gAAuVRNxQUMoCWSAv1Z3sCX1Ht/daL6zTF3P4w
/ugZaaI/gNkU09Xl2/1HR5Jvmlau71IgWlChOCRND5Mua/6SA2PllLj3MsuaKb0jzkRVSQVmQ2J/
RNCaJeHzZ99YStOG02sCt7aatD2ETsq7buAp1FB7VFebXGThqWREO5ruDs1Y1dSyF9mt1hdFiRI/
OsJvtTi9A+aSreOEBVYkYnSxxDLj4QkbNY6UYHukqlLPOJxYYPddx/nvN6RJSnJeyDCoI7F94FAc
9dRO+eFL9ZnNIRV+gcuOG5Mj9QZpmdDSmuNQPfgem4WLWogC3l/kAMb48W9Ft994oFni52GDr8ei
GTR7vzpZtB9irejikejxpRgS2VpHsD0ckktUakcy2y7kMSFUU0Z4gtHFocKtHuNNrTk49nvRcqCD
3L1+kqmmS1Gv/f3w79LoYqNgG/u1dBDTMcsjyH07HRrAAEbEHtMBVKT6q2Csb6P+RgrOnpjRjzWw
FRqO/a3Me8GabnCJS3ZLaUxCXlaC8pWKILx//cl67ARJs9qX8nJZi2o7U0x4tEKSF8p15iih4zqV
wUyO6GQAvuJEVXRuNUNoC+eQA6EMvStkbV1uxJATOsrshiMgoZX95hya3G+Aiwqw+n4UjzpBkD9t
EVFfAgh3DKK1B//Nay0H16MKEuGNhAYRu8D3nSA/qmMhdoSIL80EjNbmWNpMS2LAHr+0n8cLhEUz
50brBozCWRAVHRFxxRteUgwFt+qQyPrBv0ZClwneWpWBKMv5U4upIjPWyBD6nOyKdlM1+4Cf9jzf
D8ZAflCzEj8+zyJz17zj4j/73IhuO6i1u8oTMmMS1jzxsY4uMYeswnmIg7iosp6ndkSjRxCyP/aY
nhUmxDhNj2cSc/r727dBLH7Nvia0+e3Dq60acE/2hjxfAMS+D5H+xXeMjXpZ5BsOjfMGlwSga9KA
ekGJ7vG7Bbxa8g6sYLpEkGNvVr4zhIxN3yg0C8N6JRh3pCpaFZa53+eMJk3/d4JqG6pWoLYdJbBC
BR7h8iyPWET3o/GqZBCTKXxkHQeyYI2V9c/ePTToAST+iecwzkac+ZOUD9OG26MVfVd+somEHWbQ
dyX0/YTYw/Qrq8jE0fPv559PyE6nfkZiNcIwL7V68kixXYf0dtuXVVLyK9Negpi7N/UCHD2dmg4y
GYVNH0JUCcSf3ZXkhl+0xSrpSwRt0+IolxhvGAuRZZVJpCXvT+uR2pZRM9J36stBsY+HHXzxaDEu
MBA5uktZtXkZn4nyqIZGeln/KzS8eZcMDH4mHK3CWRkuzaytW4M7F0dQSZ6ntMPLFcDzJsMFuIqS
+XvWN+29t9J3xfnSdkyMCy+UedtNV9tkb4x+hWn14sCpo2IimMwFQatCYHNhpb0lPd49jwEgFNwm
GWTb9dPr1MqbmeqKsrEBgBPrxbt7iq/Iywl9U64H94OtvkMKTrgTi1irC9KRv/Qk0DCkHl3Sa0W/
ap4JZdjfEMmjkUW+X6YW8H/s4BIpnIeieRmH7/NKi+sugM8dtprInYMvBEZ3/BjF3QjiD5vANZ//
N8IkpVjkqSv5tqodTmtNbhbOdbRrjrNGTgBRG2+YQoiM36SCkTUVpv1lgaICx4cBrF6S3cevsuQz
x85DWHx8rsA+30vyMMzlgOZ54xoNry8N27L+9TkEYpL7ffQePNzS9uk4rzwwFiF0v7QKeMf3z9N+
05Ng+bObKTDXaGCln4mJStyGXdnrG8uK0oV1GvRwOGCB/dPIrQbattXQncw2jPSvuoFt/ACoBk/9
n9JC7if83A6BUZ/UcbvQ66i0iviefSA2ScebtHoHyVgL9EzcLXZefhbtxzqJXLQzngB9A/R4cSsY
4/0BAbKAMZYqWjhPSQuLwgbpQHhN+/ZW6V4866vknKZO8ZJCe+wserOUVWfRq6E9oie38elgp50W
1Ji8lFEErq2J1mstOF2HWLuR2KzTjCtE1QWZemkkmUFEK9cFtWzL9a5JLqUvSkYW51BC3b4f/q2a
Z7svLCDvAF1zhZylc+iTpJMkRcafm8UatQpVptpBzT9XuK/d3pGyiEE024F4G1UCC2/2gqSAJJpc
8/IMHrB30CuXZw1xvYQEgaweUNBXAufWG7Z96FCtT1oAEMu5H2/4nDiqhu6VedPaueWY5bLPlzkH
GfSfjlQNGsbGNmFagFmo9Z7vttLoWvdydxR5TLMEu7JgTEanCfKyfabS9ZDnHJt42GLzyUU2+yWh
Ys7LV7vlJuq5BplK9njetsXLs/565K+otSoP8y8jhNRqJyRrcrmUjmVaaBCoO1RgNhORNWJ50q6U
bnw6sbJq752QG/ri7PJ5Rw1SKrOk/g2ZTI3OqGKKULClIPT6cJNc1LccNEY+WUvgtQZH83XvVtTS
zKAluW341wnuEbppAmBl7cYpZr+5KArfiFMFsN1qymSQhjNcJUZJYrNKnTpsDnS/IK6tiDmWFKjr
VYbBqwa0E96hwUmPtzvdW0Rs7NCBba6fdre9y2tPaZ4/y50stqhtC423YAZSQHzwLpQICr26iJLO
mF9CQLW1uWr8Qnr1YyOkBvaR6raSNlWWyQcL74014nlpjKzWfDotfvjw2e8nUeBj/hkyB2C/bz6q
1U8PeccudgCVoRI7xcg+kQKU6vvnFFL4/YSud57pdW2ZGVHj4NPvL8Kuc2G1xVkRGHpmvbppWwq/
+33k3gwMmjPVY6HHpIDb480LcyH16Mz/k6gMGHjbhD+K9+uLNjPGLuI3dQCzYp8piwe84OgSpL88
SXF0zhS/r0KwSK/TOV8RoTdbZ9W8ia3uS9WAIP8tNuAN83MPTmPEITMdORPIXhooEynFEGzH6UBA
LEOBn8qtI3B75W50pVqNf8YUwamMCZfuViA6CE3bvQIbHNXqD0YpB62SdjFKqXIE+qUBfEaYpf2V
asEln4+B0PzrwukHWD+p3n7Ekj09CfRYY5Werh4hayGdMNNTXc3NnvhaxzLO0vBnbKbs1m8mmS55
waR5zBR5KfO0pKsZdzNzWb+UuDmFSVZf3PKNzU+n6sU11Ke4JVuuIm/MSKHpKapre1uCw48P3YRk
NNdOujefCzeltMALAc2PuA4SQLxE8YmtsNSB1SYbjZ+i9/fuEkYfy2RhBN3r1z+bpcNIpQXas7ln
mB/A0feGhHREQ3odN/Hl3yMYMuQiCYLxSo3MykzJU1hkHl42yGIum4UCNC1YLXrY/bFzhxpTBRts
C1Z5dE78XFvXenAkerHhvUxQeL+zT+Ze45iTFwbEkR4XBlNJLXFIlBvVIW2KONH5iccjj0Lvuhbz
LzRSj3Azb0LUZrrxrH4LtP55nPu6YZxRL7WLpMRfvJFTXvd2xgATrSbXmM1iN+qfQLSp+Mv4z1ZQ
BO12SFt8K6UGcRgkoKk/cK/kpwysWWxK1H+En1HtXILljldk5bnNirtPrUR8HPb0IBnHvEYXREZc
ryRZRw8xptJ5gXbZTVhd2M7gqCRuy1IlnJkvRQswfAvhfb9aru+uOLlaE26exhsUJwo0F4aVVGK8
WdNa8yHNc5QzlFljCQp31k1GSmykGjKfbLKixLIKUsW5fdcpNhuH50MbRprZmjI2qJDhFUqQQtVz
OSNPgEnX9puQBiehVKG5f01bo9Jd5MDxk57UJ2Di5FIR+Ogg+klb5mARDomIloG79Lutdnfn9fIv
nkk8noRPjmig4c90sHuYJ54iPmzYrOV1kWi3HoDLe5AHk3NAGsoR14raXiXQKBfHU2UF2hsv33+G
QYt6dPB1qulo/w5ckrUWuKUklIsHS51B2/j5scXeN7Go7x9Bx1jEUBR5MHM6uKs1PLA31ANu6Uwg
b2zuVvknsUWXArQK8u+QJrfZL6frweTyY4WWjPEg7yC/QSKeB/jkMeyPt315uzEADX9LW+E0RJk5
TRMocN0EszZ/OHXwrDCtTR3UuyPdECYFY+rnZJbk5svUF6ltwa7bdmSKp7XfEPWARxO0bRyhPRUn
HTzKmRtaK3jyjThEsb0NBBFy4O9SbdX2lYnqW6IlM9rIL+dGkoIFzp+u68+dsOrgsBOiUG6t/XuP
a3dbkx5+3ak/0gTeiqC9ioIGKP2xhqGlo+d9L6ChaPydc8Rls2gvgvUxzJI9lonFMGNVv/9cAtu4
2PtglamD6K40yj+bzKS6fdRX99czBzKcCUid2Zkiho5IYv7Gz4DWVewZFvnsOxNtiPo2DIgsbqxK
ijmEER15KQOQpVWjQHZCkKdvyFBK8Hw5z5ndbciIr/il2/MyHsEMpFjHk7/DRpsqkZOJ7kTh8TpJ
25TAAHR15VsRzXvSuvcy+FILryBf/YrytSqqECFd4WlJwiM5mRtMLJXbgUl9nInZQM90FBce86/U
OXRQTvR97BWU2dsaaSXF5ked0SgO9ga7as+Mm1ZnyrPxjHVAvSBbGUcJo4ZjcDbJugIntSCD2wRT
9PeFaS+64rA5QEoHivQiaOWXsb4QtyTpv5oDe7BT3JTa2StreNajZK77nGntI0VrEVpvALBT1szq
ZqphDPNwGqv9LUOVpFsSeG89l21p/lDt3Uj5GYCPnMUiFpwwGZmOt5IyeG7/xF5hCUirRow+1Avh
JmKFwfcA/vs2Z9B+Z5tUUMV7tC5PiuOBbklIrbph0ZRogUx8DibNn9LjWmQaINVvCq1ZO8Fxcz2Y
o9FiMiTJbXSc1cryeNEywgb7Lyke0H3yCSTmSFuZ8K3GPDurwSzSr0PxifAw6FihdB6Pp77PiM5p
Aeo5676z75pLYRwz7D8JsGpoJzZw+FelBFcFGnVB3t4WXnLkYRms857g0yZAM+FWG3SZ1cssqGAp
Vv+BC9xaXI+R54PfOFFdhuqD0YWDjuyWFN77/HfJO5sIrRIAeqFVQikgmuJnbgOME9EnJMZavCCN
HGXfjFkcvOVqUSgrHwAJRJZ43TU18YaBubqQqv2TozU0qfVoOEBstLcYhDPUXCD9nxc7FfKmrwX1
M3zeh0XeGXD3OUx9K7vHRdfq/Ez/TQeE7xHGhBT4lTBRviVUQ2JtoMvZjnuOqj5XeV1azPxeGdgv
5r4PjtmKWQ0GiPhPTZR8C8fW2oDLpRbQeL2oaiWi+k0SzMocppMff6VdK0LStRkD5VNrF84nA1rR
U9iTXHqYrhDzKSLVR28Oe9mmkANApC+Kam0A9kj/ULWCfxkR0V7tUVzOCqRDfJB44HswWCtrK2mW
LgCdCXCKvGGtyHl0FoPATaTxRMpdW/sjt+HItPtYM7hlF5Kd7v18rcNAnVp9CllDUpRvRkNhdbdE
Ua0PyXmhzuqpqEMMLG5gKwAnpKpNSQuH2g12YTChbJhTSFj2Di+/kpgfmYUx6hZ9F4td8Lvn2ajL
nKFxuK0BNtILZ7r6phGcB3P+1GWbV/hFIYNvx1WYtJ85bjW69I9nddfFqAC5MiosWVP3j/IecvTY
cf5VbDMAp1SXoPMLmUOKriUi3r7jJC+83MXnkr2NijWVeFoLO/+sP3/KDbUPKzmyhkdMN2OKfgse
pXc4wBhlIF9FB3RE1bzypjCY+RM8tzPzHd1Ns+Hw2yYtdVfD3BYe7wpMM7GDHNWO2+Fh2KPfzhDb
kvGtElAHKVu+G/gxmwweLrwZt1iT34gN871/KZTrgqxya6hCEYCdis2s7A0H5CK7658pqelP53UN
LqTb75JkWskOOG9BQ0H9W7F9aVDy5LgdOmAVtqxS8eVsxpXFvI7k7OpB2fDg/L7JjYiPry12OxGp
1GjjgCAt4VXEueLKTVD+ddOVts2267PhLxy//DBSgqSRuFem7Bjaz+I678j5rRJ/qz9tB4LI14qO
PAo+cuk5ltHCnc9jbw2kF9Ac5G+La/GAwgjWTQGQRHL3asEeU6t/CZlC/voPIcrmw5JzHE+pGaiX
M9KvxqGmVHMeKiMdPcVzQrnN90cU8v73QwJlh7EQUrhudD1yzxIFfIE1GFm2tKUBCFUTtICz5WDV
UgcTfdlNNS8LiSLna2C9VzD5EDtGD4wPG7S7qPJIMhRuoEuc/5pScvLa2trZDMnqeMh10Mre9L1O
/4FT+dm1KQgeag1Gwgib/BaZJStdAWymGgQCtfVj7fajVj5pdhWK0Sy+/Ky4hG6hJB770jy9w7zt
xEt2V4sShWQMc5tcOP7HJwsz5F5TFKona28kNmzJlv47+aO0xr2IZtfHRqGW1yNxLuzEK6eK7LDT
m5S5QXZlW1waZMlGSpwbA9TJfiTDGqgBPGrCZQ7SU16j09gXsZNNFkhZgTlWfWXaCtCQA9u1TgNc
wxlpiT/y43wIj4C8xkiy/bENoPY8HLsGZL4o8tdzxknalI/FUKgHuNLe0B9wdeh7R6YWV1PTNoZa
gs4gzbXTDa7t5nWDdd20H2IazZMXrOWC4dMM7rsDXTo1w26TVliYow7UtBU8Ei3ZhLrBHpbxMx8Y
3ZbdKmyZ54JgA9LpkomkOUlGr7zEbYn20wXxLpMfgCTWQ45i1z9KwujgkgzsQDZZSFxJJljdqADE
mJ2CbmM12EN3bkxydTB2F1U1TOrOdqsj0tL7KBTGN1RqR21Lg1P1ARMTyguI+tXOoNRkJbGLRlZO
azxhBGRbWtUa/5OuULEYlj9MHf0ocb82AUcCAc03aeJLSqdbtdgwSHZIN+UE1VnWJlsMtUatBfXO
Xuczd0YG7k8s3PER8FAjEXkMbhe/2MCRZfQr85NTBNRrGXT/BxrSwLY+2T3Qo2tmlcViqdNsdJM+
/tEJdsPrwqw+LE15+U+jGKN45I7bn1ENrWf3nJBKJPFCa4QWHyl1d2eqQmlSeU1JJX9hoWIqmmLH
UwWQQ7hdlretCUkoPJnXEXMUyNaBmmMNkYI2bnJlQXZ3DXdh/aCH+QUoJBoYtNYZHBcyQPCRtCLa
Y0qh3UDbcGCDJAsu+X2fjWlDmuJ/NwT6URogu3ySJ/4f1Sn1VOFczdBKhu6MlH+gaQl+IhYW2zpI
D4vP/AelXGIgLP0sLUf2DOO7QBaiadE43CrCOkZlGdGIQaL78lFU2FJEn1Rf3m/fUOlEH+tGwIS1
L3lwnAxwcNZA4ChfmBRwhk27cKB6KsgJVFh7dKXPUwNUy5/b4lfilzLZ972b+GeXu4WQzt+heong
x7EqQr+gO9hcAGc4g9A/zie0oBYNOsMpX3AEILJbnG6AHakYlbKp6sVg5vruA04y9OXLdwJlMtBs
ZRngGtRtmSoAURBSgOvPyyUBGXSfKzAd/xwGiB/yyAJxHIHlhsz+bxmnVof3xGdMvgKEQ1GCN/yy
Y5pAZ/CNcOOyGur0hSbP/4ipiEAR/dAoJY00UhPBhTu/rewleBhJet+2XQXE4C8IFsegbn+PFHwA
hSi6RhEVRvZGyLkHa8zHukzByTN6HFkoIQmh+zNBE2hogsiYtgAbxWbgZrpGkog7wkarU6vi9HmX
Vh4PskXdVowbrxyxEhPjsWuUMdm5/rOApjsIZFaifko3WEo1dwjRbdOemi+S75uKNmDrwP2uANf1
um2M+DniALWaHr1iG+ZuwqIcPK92Sa7FCN9AQS+YbiE03XnqnxUWyCfB4TdpQRBfA7vSV4c0BiYI
x/mGsMrdncpiZKE9iDoJM7dCNZTmr/aHbw3VzeH3O/Hb+/W1z7OyOb9TFWwp+aQxXuUMnPuQNUd/
2lTCAUZHVWqNPMWxV9i7Nv7HRBK9Gxzft7ArXqvMiwiY7Co13CTho0+/LkBVD0PjCMf2f9OS4aMz
tMXFKZH+WxjubMWW3rPGpSRnuyTUvhxL7Fn/2fo549ExJy+MlLq7On/gI2lkI/acxASIQfgRgMBI
fn+fIN6pOarvR4VazF+8NMSPO1GNYByATixeV5L1e68LTeeOcROOqyaidw5GbtRLTjW/HLHVkK05
upNTSdWeteBAzb9fRmNXmPkuCi0vuC2FqV8to9UekYdunV9/R2+NT9NA5q9mLllEXeVjoRqNLlFb
PS49VVfXFO+wuqjA9Hc/HmGWu7F5wdjecM5tdJ9SQwnB7Sh9okwenT5ER+GAd/zfl418AFnqOGmY
xy0zYOBOsXGpcXgDC94Fm2AAlFCiKN+yYlriPhz1cfO+pRi/O29dmUTTuzotDk1XegOarj2TlaPd
1jUc3opM5tUgwrgcEbhchNI3iZYizUtatQRny1tp0EtyhHXHtHXX4ymjht+q6IVemynFS+wwtDVb
BAwtgD4CNFiL0HtSyGON9dJ39L+LgQLgjne/oczUcBVogBE6PG31Iv5GhQQp5TJ4CS5NjWFM5wBG
wDTo1/rqLKv85C8wtWi3HFUcDDvvY48jagdGzPNTCWx3lQdiLAVpDNtTm9sicF+1O2m4x0WzYZ03
Vkxdc1ElANy+/mIx7EVAQaZegTf/8iB9R5Av8w5iv+ZybBtCOlCpOIRvL/XI7QF+VcroQN7oJWye
DguP01XhOkhGhQjoEDnuWiKl7Nl/iO9WyKXSdk/Rljw8eHN5eF+8/7+/BZ1PecYvCKWQHQdzOgZq
7SKsOWDPvj5UHmY76T4MMfMbC6vwXXdFwD2exwLWGKUb6TFodAcJ/CzDvr8Dd8snJZPl5hR4GjaS
KS0PJpd6Fi0qdO3yme0wWSlei4K0Gy4Vc2yxwWi7GZb+7NYjzFs5+djZUXjS41CbCqNrx0nl0PXz
rxJ/aZuxr8GtmYf3SQwAmsSB2lnO8XGi5MuwEATuG6QU1fOTDVhFp5QV1jTiC+RLBbJIE1c99TLL
jy4bsU2xvqeJfM2ikI45QltYVlXP6zq6U4ZZth1l1cjWd86M28FVUi3x4WZEy4owe4pZFnrCS852
USLPJVBjjXXTOiOSJ4f1bw8TrMZqt/sflvnFpdsPMXkzlL+P7xXJjYTAuTvQUfodZjXy4Yg3578U
Av0b4FfNmbDF5Jd1WxC72i7pDP632cMBP0WEVFPiJ7hMu/BeK5qpgP7u4rG4DF4Ae9PYJdZMIJ/Y
mmtGRTNvMeY7v/hEkkr7tmj3RxX4d//3jfmIsYR1OK4XdHSWrHPuzy0lCLj2IKXAT3QOFy9Y9MbG
BJQpwQTtX3g3RR81hf0Tz1e/vZwdVym7MsDw0OE+A6p8RHN6rK5GapgFAObS95bWa/nRUZjSArB0
lrK9EjemRXjJl/m9Gokwjs17/rzXCXUxruVkHDx2deH6LR6P1T5ob3VyrsVZKt4413P0R+B9hBh2
0/gxkDeCXvWw4JDHbmEubZnkOdH+x37sKk4Rd0+kogFwKVf3o5KPnYowN6qJFdg048VRnPvEl8A6
B4lGPPlV7MD82ewaxnojhnmcvC91vySTxLHPjxl/S7nYeTvvHP/i0vKwYsY8NwWlF6/HDll7qV4u
KsY2UFxyCpRr62b7XlzLTr1uIsK4Kwo6r6W5xes1ecVETxBcBkDxdsxZuG5bFotcDUNOZBI21/fn
xCBqCMX2NgXkkCW1MUNGYHPDuOIBOLhu2bE6hENlI1xn2cxgdydhWCQ4cS6WpGk9JSwb3TH23gPH
LaGnnHvROWCu+5Qc2n7nMUGK/m5/ZW3wi4yFvqYwoR5BmdmoH34hFQo6FtAn21L1VpfT3o9j5PPP
sslLbZTGTIeiBBBghkt+aGwLNt6lPAwr5QJOhorRiYcWDHKR1MitGolP3co11croyFtB4c4v7e5W
SeuN4ZF33sUKmN8Th1XMSZ9XZatdJBvdORxgQqd+z91OQ6VahdNKN7HxNPAWUNlT7lV310HKApkf
fyXZus56YublJRahv763eed/eBaFLoSzigMZg3sAyXRq1eMFMje/eOWE2FbZV6A+5Ps+/ySiIzaO
ZQzEVy5EK4fpyO4EdJW7p1dmzrh9j8yI+YfC2/ySizEbpP3cE36qGwXYau2bcd9ms5DVKKiu1RN/
E4L4UrogxpulK7CcH17vHr4iLNLDxUt9OAP2Q0BqUpt+MNOEm82duoUnPc7Eq8kg96kCONzb5BDU
mvaktL7aDEncuTOr66RVXpEdEfgqwXR2ii3IVF6tv3ZNCc3d92t91DTp4mhcHqNPhXHZUNHiGO3k
Z4IMrZTKCvME03JbJsqTCIBcMgyL4wtc66rC0VKY9G5BqLM0FnRz5H5qLPUhk2z2cnwewydUqxp0
d8XOo83PrnqdsSjPqM+lhlatvNVpJViHPsHN2Dm+53Ynagm5VjtK3QdMx9K6NX7PhKTykWQSub/t
9GCzFSsV8lHhWLVPuidx5JdAwjipmBrRBr44IN6F5S+KlX8Mri+gjC6u6rUJxOmLZePDYB2FElaf
a7rGV52PH82RA6W7cC8/ntoT20QC0r00iPQ6xG8hWvGmmfPttIyqHsnHOPgd/OprE+7QPekYMmxL
GRkoTuiurHdcNWyA+TOTC6SF1CEO/jUe/dWwo1P+VNbbcTKd4d2oyQ5ox2e1TWH+wCixsJT5P985
+uDPUPtjq0kbb4CJ1xQ4bSHUWZjLAzYOkIHBWMv/E/syU8Rm6GdMUbGfk12N5LAsQGHKHmnRB4KB
QG1yuzQe/QTEp6bgsQXj/Cvnu6LBhdQimAEwX7G0bnV5R1DsUNHGDMkiQ27/tWI4lQZwBEIPF8ZT
0eRyWgHxIMwbZK7He0H1i/otLy40gkZ8NA/9pGeF5XcDweKlJLAGxR/VuuAZ79nCOznghafJwenV
DkLdwUfuX+OmJ05aiivD1aZp4poOxhVkD6YsIsZcnX3mEmoNc/LNhD2sod2+OSG0GlAzfcwGcu1i
+OQ9G7+yjBa4WCMwKDOmiIpDQgfVTlULqWg16+MZX81UZt15DKGflpQIP7SnLftfDuIBlq4eEE3I
+NRMYXnZNIgPkzQocLSlSJL/udclFuz1HsFXPij9GWddMRla4y9ueSMqUpV48ZIU1bsHafsqFzVB
m686dzHjak7MWKdfunml6jbyteaYCLuGBjzSm31Ca/A9GZCVKSqAlp7zYkO+DW304nOxIBBwO2kR
yIbWeTVvyvcmyawE2PKuER+vIY5UF0hgJh2dDrrRhCCyci7EnKCmTNbkuSmHUA7ahUo+4OVvLsp9
mGhoILGZy7UeSFBgc1+ucq42UBNa4ki6hZ14EGBIk//hjxFRnK6Mgg/X/jRH8kUekY8VoHayhJy6
q9ngTPtP9m9rwArCASH+wNg+Fm7Q8Ryoh+eXpWOeb20fexZhsBpYZ5J3Gn1M0Ue30WAGIK1vLbG6
vd+9cZVrC9uSq7yQxHiWj0F5lmCgJoFgPYfWh1+fQKyZj0rvi7oC5/wnHvfG2j+F2ekkPsc/Tv80
49j/sGXzePQqHBtZeUoZ2LqlGwPr/RVpvf2FpZCA2LzCDNSW1u98+8UKtNL18cRpgZjpA3msafrA
yPZTD2C8tYtsaOFr39gDLaAyoagrZ3xlNiYXetZOKiVvPB0wa6QM0MVA8iRDSSLhYTyHcZQlrwz1
0eV1Dtczvwe59ZPOTENM3q9ubkk15xoiru/eesCeLiO1RFxPtd+3ClIejWyl0kaW7ePiCr6mtwIw
/DdncTkdHYOEy6lHoeMxZ14DBn8OXegU55KSir2YgbsDpiZLKmNO6CWZUZSbh3nIJymntYqkD0UO
j70hwymuLrZZtmiDArRDDEPEtUyLoaYJoB1fcQ+h4cDOVcFGPR2flamlrzpS5j6QtrD4r26ObSKZ
EKoJp29SqypnBhfa02xwwfNWtyYWuJpZJmrlNpsg3IHhwlf21iF5HKvMlIURmXpBz+sG/oqVcwDE
Py2uugIb4hAvjhnta5ATVSm+y9lmCxdrroRvepvR+mEYM0+UXNvgi5FMqJP+HjP6KfMKAheVYRV6
SUmcJphrVt9KCN8wXgq6Wgi1wFxH+t7a3b2nDV7ZCCjK4xl3m96/sPew+YkXxqTuANUswzKaSYkk
B/wesfTEZQJ/Z4zfQPEJEP0JF5/cRVt4V8CRWu1wt4HDXq+iQ727/HY7scZOxcxO2LWj4r3aFPmY
qjvvrJoW33lE+x6j0qRmH2LEa4v9kR3CQygV1ZrW7v+4CZ+tn4GsDXUhn0R1STGDRRKUlBiJqNCM
xhsYnAY6eIK+QSZi1Z70snC8JRRT6PQ2wHz+vknEcFVB5WE5QGptKZNkKWdLxsYYcHg6HDTY4XMJ
07080z/iYssT/xjKLpt9P77lnbBJhA9AMcNR0y7Z3Kh+dfjAOzfxCUz9gJ86R16rSameHTQL9Asj
3msDYVab201dJ9+bRKrXWuNahbVUAh5RGdKhLY+4Zfg5DwiTSgkd/vCP7O3+SOThloBJYGbavvUy
2Mz72BPCQgCWhnU5vJqP90oEGliVH9HEfjCz5cafIuh9K08JuDqcVRYTl9Hb9d47H0epi2H3HEbg
KU39UbSQV4erzOwetfIf5GHRZyKQtZtOAdIQPYi6Oqh//sS83y+yIGknoOgwcXut4fjtpoSU9nRk
V2+6VZ0GSWVpvkoYM3GWYDMZMPBLeMm7zI200xAiuxBWOBZ5PQOm42WeUGDIIY28q0FofbdeVH2t
DVp1yVbOfuqkZmtFhz1AoudJPXGJA6H3AXqk+sBCsjNm/ukZz/9wA8DbBcyUxyYlvlJZ/V66CfH6
gaEbvJg2nTND1CX2ZDNjxupRnK28YXVVeMa8Jo2OWsSrbQ/mvCL6sT1KWMdqqv8+wpkzJSQuol7I
opx7LHiM/dCrw5m12pizScMpUuwkszTl/vHAZVdIfx2QTjFY7YKquUYQuQbqB73WZ2aIRRffktPg
k1zZAwzBgKCEJMojT06nvanXNe9aRSiWpkyZWqyvVaUSn854bgrc8Dn2J34x8nReZJbxPRj/bGzL
PuB+7uYMWrmy2HY6SR7R41dDBtqMCysNa8xI9g5sAmpmpPL3b8Z/G9JUFChqli3gslwJCNo/85rq
YEn5SHtnM+e09wWTZWs9kH2rU6GXi4HQEtHQjT0IoYUEQPVbFQ+eQ+ZmYMxlXuMDmXJW2VBbejyo
wHOiQL0Q0ZOY+UW2V9MvI7QaVcFAK7+VZIjSkhn+zaKdNXKvemNO4arZjyTEwhfp/nNHt0JfK8Wc
UUsxQBTxnE1smUV9DrjcrbqsoUFlsG/UalqxZvwBlzuIyPosDaYEPN5NzOy93MLyyWvtvXItwCoL
ftkSvzHADLWR5YhV5PD8ntTx9Lahdt+PVsCBxKxWqxFRbu1z95R42sOQpnV/vUTNGwpBi9uxPqHd
ykd1x7GiGpkiH1E9q65VzXSB8vUshgkN67OR5f7AH9sfpmnIGPQCfgZRjTsIxeUdZuRz6nHcqddc
bOEiiAU63HfmEBZx7y6EY43wu9UECZGYBD6pKzWKpiaVXIgoxPUcTDP2mva5+ZqkNepoTihB6wga
ATNKjWK350MMJ8uWvFrvfrWftSfkHGvav4Ee0gVNB4jKu00pB6FdwICFFBSfG95F4RLstyLC1RHf
drVGYoJ7A4eO0N3P+NPhaBBE9s20hzSc9GdUS01cxQbKEVKxoYTrIShE2wLUMC/9g3hMZgskvsAe
ax6OZ1t7x0iDsKFESVYyBV/eHwCtEZpGQVlzhVq8vmbwTgmT7uNrFHd0Wix0J6HMOkSO+Dtla72s
wvojewnPyUQmySq5TFEcUoXf1P/k38FUO+gJzlFgVt1XSPG4y59L5HfsNprN9dXXToJam4kKu+vF
ayc2RMSJ1paJodsSNZXeSGlY2InRvSlD2pKwKk092XJp8qU4kue9SrkV3SmIPGthuSV1tE9eOhO6
3Znod49nRmqsTZVESON/so0dD0hUM1EloY2rmoVbWWLtFHMBH6LY97+8MBkRv08NR+IcPP5ufWBi
ZWN6L/RgoPcSym9hTQ7SNr5F2WIiJATdN/cD5gxNq2jv+ws2/+b7kt59kDqvpZP8LWY2HryLNhue
pdVVmWZM/ylJKBRfWhJ2k1tJU7GDOhnWklJ1eaIxeXIHNoh+w2LiaFZ0ns0I4k9drdp6PzQJGW0y
XQ65xX33W8KZ9x16XJCc6Fg42xfA0i+4Z/Bq5yuWSpx3Lv4DauhhV4bYOQvjXs+qk8vANmrWgnZd
R5Tg1zCXKwqg9XMxdg5TVgtl6Fzvpcv1bIqK+nMmeC5LMGY0xqMuLtcQkpaB2vklpTww4WhajBji
msPDbY028mY5hK0CQbzgfOpIePW3OOIb6BDBTfLLMEjKyYw2QS/yIPb526gDW14NsXXERx6QSuD6
qBMbi73APJKknLT1/lICBisbMEfV3V84+5FWTcrkmh3uSh75V0skA6MCmDvjdDSVeCfPWThxCk72
QUO9xyxaTTBnknHa+/CV01QZ8sP7EA0g5+8vgqqg6Tf19n0Kyv/O3ohvyCfJsM6F8R1W0RoXapCp
x/WQCLteYMzXE8+lCVPJnuh013l/kxosXy06ex7fd9qgymmHUGQS39Uo3xYHZgC7a2nLBglaNEub
KYaussNBBSGxGvfuS9fBiQEXozw3S4bEcd8Ab4+ru6O9+SdDjbMKqswRAmow/PYdArGyfr/1ZzHH
n0sslUzxXlFhF3Dl8eaDV83KATKsGT7hGCqmmrwO/aG65Hsb2wBT6FQE3C7h3lyW9bZgZO28nhC6
tNCXDahFFvIPdjb2ZWr+V3E5rMEcLSu/Adq7fqIskYPot8lZzp9MXmRT03bjN4FJPhkKJ8S/Gvyw
XuCHEdZ5oMDgZKOpXtRUWyBUXi8+tJwMoqAEhbSfIyp3s38/I8O036S16e0kfZprpOUBq/jOboMT
pLxS9h+UZGs9GmjzSNyLnrrKbFQCFqgEbo6SVHYAFxjihwlpaKo6uYUYES/RHSFWOTvzm4nmypkO
n91SBKEXpkT/DjoXLsvl1pZ3HiDOw6NENYwehb2E1RX9fAeozmmnZzx7fyiueYSj6QQXYjrH95Xm
tvazCvtcc4VdyY+StnGDg48ArxPsjKtze4LjdxM8We9ryxXL51kyJn0Joz03imBVN+qbOZo2P4N9
pHa9OvxMaf80fXdKIvogaotm3jbFE3p+Wwxq+b4Docr1tTZFOb5kmklkhV2JZNMaIIyIo4AjUyl1
SDJbJIt1SFtL39sGcxQFe47QscutaB+sU48f03YY9InwFwF4dRHTmBxk3SLotgKAIuauBbzwtAnt
65tnK1EPz6kUkat2SC3Uxy5kjKJAaQWi4hmc0cgkUcIoBlfu1l8sECFPpDFNx/uyeU6ieTTybjqc
KhpJLHjfvGmdWcQr+L8XvuMD/2CCk1OFITTU8ElbIaARd2vl1kSFCquryQ3mUT7vrQkI6vI7LNxt
GzubL5A/dTTK/q13PqPNVNUnk2MW6hE3sz0GovFEfC4j4JS8rA2UU12BLu8T+CuIX/k24A4Jdxej
NY5oz/GIHEe5Lg4jwWaFfhSXVhMtuKaqqGIIw6s9aeSnrTmp7yHNwAPqaW4lDyUtlFR092zHwxC+
JnQi/EoumbGdeiRDuXFp77ilkfVjkeVNsjC1CV77EPJ942EK5vBw5pQldBKqxZnJx5pIS82t5BlM
Xmx3iCCSJDLvVZVLmMR0QvtGX5LnIyIfXcMiKM8OZQbdo5v9IP9wRUVgVeA4jkoV5mzhxozcnEvX
AWyRGB/f9WibLyMWD18BVr9qNpn+bAYMkKUythlOqmztD7NnJpi0e+RY9T9bdMsmodkNSJZDeuce
a4VIO8wzOt31snjNkKwzeO4tBO7WM9EiA+4QILjn+9fk1Cn+wpECBgcFyx8hKCTiCkRRUtPZotwo
HYxfASALcYevIJpNBDPfMgSthD1Plpumspw6zAgrVUmlunwXI0XwyV7TU2ZrO54H3gE3HKL0x61t
q1x3bbRYHVXxAZ/6xWF+JiVqSoxDWJOBlWy7Q+7fB23/eS8NfKYAtgzDM7pQyPj21T3K0uIzitR4
LDiATHv3OvwJ//rTjxSsOzCeEuPjVo2850ttfaGOR3k4i5ibGs6Dodb6cBriba0y5YaBl+v29L35
k2DNKHGeZMYyJ9KDH8ESbvK5MxY8ID+8NCOpyHRasQ5D8rCJj2NE5RxKC2x2DOB2BBzOKsEzNhEr
NN1tyneJEgXaes+02zprmsP+d8hJEuRudjA4di2IWT9iTU1eCcHoEqohBdAlcBN96Y2MM+iQh2oz
HeVs0TSZoO6HuYHP85KczN5LTP+n9dUdTOJgK7HHwZHTavTyndvk2P5FVi+Fg0XQcn8+yU6hsnxU
GC3LLN1+7Ksi4o2zqpCOI9bpR3slZ+M+WLcdQUV2cRwBDDG/srh6iziPvWehvEHaiXq3bfQWGsRz
3UYotZxqTLQkamuFoW2d9k2wkFzi/MRruP9n4/CfxrZ3546UEWflYJEjEKc2S7tn98XUADaDM63r
xHbiY2voHb4Myc632PRyELN+IhB/h98GsGmOiAyVaCAPPfAohba+syYU5sZWJz7rPXbTpDTxZCmI
X07m8YaOAF5XeA3ZyLFW0d0vq6RlI/Y1BgMw39vTYNiI7Oo9q9r6dI71UHmVRP2Pxsy1kcGlRWre
BMGqfEPKLF30qvKhU0Y6N4kypar12NM+KUJoA+CMjWcGofGm6fS0I88UTLGdJ5UK6q6chghlMTXw
eQzpqy2+EROZ30hcSx9EemS7HBDDJdZGG3PWosp3fbhr5G/6zaQUNsGuzAWdW45n7ggb2alcbX9f
na/Wthijv5Pq6gixwh2F2nIn2VBzjXj9SgaON1pkqZn7/QOyH3CcjzfitkWu1QC/uWgaiQt6ULbC
BUS/f3JgjX0RjnU0+qflwiurryGaBChEHyu5vsmLWcK06O2mKEHRqmFCUmttoeboN2QwdwbeWQ0n
VTm5JnL91Io9nXHeOxGEWUprmPobXfpeaUbN+uMQjLeqrORQT8+hJ2DRTDmougiCc3LIOt6SIXot
mcK16hmlAEvskTemBxgoYskQLsFarp9A4Y/UVJ+gIUHS9cs7dx2DwWJQEH3Z78wOUwX0cz6wcomN
jWQVOOsc6K8g9jxkc3T2soocOL5VwXftPU/T7q/GhicqYJOKmlhtUoHFaAf7xfJ1a9WLZnArf2bk
Btp60SSLOkcQtM+7/fS6wpgndjXarR3sth6JAhhGJBuggWy10Cpz7EHkP4ckStW6X53YSniTeVzR
04Le5K8M+LpRKQcSpM+FlLrnim9ilK0qb+KzXKxab7ZjEy7FRBmyJtuSL3wMj2bOcjo3Xjw/sHF+
zLd2beJonxu8XPKIur48utz9hi2HxDc0rq0ZHw0RIV7O72zkLyknKnQ+GtbehvTde/wK2QAI+dSi
ueNlOIF1yUHQFV1zaIuGuT/OD0ZXmnOF9dI9n6JWMNQAsuYvwPIDD5qPe1mzD6eSWt7qM2VYsCnA
Yq2ZQYhMQijwE5ZVLBwqne4xbOX7x7xNxcd9AzaApL0p1MLez9P/ysNE+NX/XovXI/G/M6/C8z9H
ME+C/A9rONu5ZdcSLoygcQ/oC22P+zgn/6PAT5tZQlXqHm6xQsVhwg397XxNGKXrzABfXPU3ERc8
4IvnTKwW1NWiWaaRU7D1LDR5scXV4T9xi8KytVWf3LX2lIqp+8JAdG5jgLiVuqh/MERx9IjDWQTC
I/UhcwA31IObxb9ArEmjvcw7KW26l0+9VsP9T9y81BBydwOY7raeA9GEjJiJx3HylxrEeirrTiGo
vI1jU+DtLD9uCnP1PNuffsc2Oo3HgTc9xAe4nOR4R7Jdrq3WvZ98FWdb0UzUwbOnTp3zHbBaCiPq
NPvG81XgI0RCiKw/n/XEAZEVp22Nf7ir/QFSFqjsKsEopGXD/8KnOqNHZLEhcJHezqdmhp+SOK63
pZJXRIV4rTT5DzWX6QEmA7c/QmLQ6KGBkBDzj8nqWj9WmvSUsK+9QIVn+5TF1dA59P19Huoq9rli
D7/P3mehq+1mG/9s61dPVZdpVGJm0IxLslgJoU+EDk+N66688DXclmyHepRid6PBZcZOZM2J4FnA
f+DRp1uMS9MAORSHTKBLfJ7gXPXMuqWZ0tNyEJyNvdAZNdbyZZRh5uVw7pNOBqHJ4p9pVJwLy7NU
bZU3QrIVxsuYjhrWKR9lF7WpoNlhuKPD0qZA6R0S25H7Sb7veXwDse/M5jNUVwSfAzVnIiO7JfFC
trqPAm9I6bBTyy+jA/2HDSCFnya+HsZ7eqWhlqAAilShdqxJtUoDJtPDZFCzGIpWYbKyqZY6em4B
8YchSz4Fhat91y7VzgHRbjITodVmgzQPLsJA6iSEwYNtSeAOEYkg16JIYhbNkRjezsKZO+h3lmL/
pSPPuQHLbAjq5ynZerZbqpbN+eazu9fs5K6NgAuWTjlvNjSIjjf5k23CcYXnzDRbWI5tDNE2PkAq
DcKBnjyKynz2mddaZpMIzA9zuUpyhOLzVCEBE8jGLz6wHWmztF1AIcJAN3pkJSJjPQi5HPFBacdk
8qIfg4aPZUUqPIgrDVku6jFEWvOjSqHGymHa732IKIKtL0repkGhQvwGlW/Z+FIgyWKw6wuhOdxR
F4XMJyNh7sggFcRcfFJwajJ7KA/JrNkaygydFPpFUjNNvTAb1zWzwxT4+trWKIFtsaQ4PSrKmwo0
OGbmYNtXTCTDclJEiysjxssmgWMthSuOijzt79dG+FiEu9QY2m2ZNigo8g66TujgEeHBsOkb1IoX
wIDocZEaFpH3D5Cf6flh6QR8AFnL1DKciENeGoFVwgUA8fHDVpO2Trg2wAv5YrqgEdeeA9KFqr1S
87aHSEfSvn24FRtkSkF1DuWjaXevJBZtbMHRqxwqnUFMZPROJ04hNfq14v63mWwFpcUAhxHQdjiX
/WSdRwfoz/o4wdSQlpVCwPgkJLTuLShjBhaB+838T84U7DX1elJcOyZilU4MYt09n54h2AveJYbq
MlAQC3Y42T8SrG42pYqvmDCmN8xgrk3BCIs3OT9FZToygOdsoMtlqYUvUhrKPWlPJ8WfGb8vc0wx
jgli2U/hKECuafppm0CzIl/1g/ZL96WuPI+D2nF2Cc06OvbiOptk0XH8PHbztHEXg+TPUKnJlRsT
3KfP91LNrYiThJ/vSHhunhZP5DDNBqnNNaEeWwlXoeVVvJl5u/vE+ZefvUGqUUddrTiUNq+pqM6b
mGmeTuFRAumBFH+RMp27Qk9FEW6MeyK1nw27XoYMlMI83K2zwzP5pErfKkWBsSnni078jh1CQzs1
hYELq2+D7oImc6cgzLtyOPaAgATHV9vODZ0Du9gZWnR7iwv8Qi9ZuApZXh8oemwGBr7MTZUQT6v7
ARU6KiVZKG9DSZLFeYwthBSI2hKv2bnvm4EdwGSUJzUJ4/34F2RtFK+EKAAf++bpWOL22SMT30Pm
5jINWG1nDtlMuPqPuifKiUM1Lll3aXUrIU7UrK2Rhj6GR+gY0XwHKI0hypBLzCsXEtBqPkKvBKvd
wF20Mzao6DOXSQaHr5JG1Se5PaalRZL12K269+Ejj329IQ3StoaTeBYDu7irfDY0TFdb1thPf4hg
wBHsbEH0n1EuEMl3wzhWC06CaDFHaxxZuow08tD8c44FXQ5WaQpHH9fih96G2Xr01MOYUx4cpN+u
G1pm1l5sskL3Tu/eMVCVPs3knGu80086t3lpYkTmS1fIff3rBmPtH4Mjbz2axptaqAznba+h6D7B
PjlTzNrAC5H+cCwYb0r0tGTfu14tOF9Pqge9wxSJ7NapYOmu1E2amMbW/7aNGatPyChLlKr2AwTY
r6gOaX6qJM5eoV8CxZbFZh5YZSK2qjQMBl2/M2+KRhq/qxo2a3EeaStpVs/z47oO9YvZWhjYCf4U
7kfHDrLV877gOXy6LNPRC0c1j03eSbA+JcpNAsjGzBQz5SgMViQLkhLhp5YccV/EtvlTXjU15EXQ
9bnB0yhBskjhM2sgEKd9yn7w+Xl6mvXQdIBj6Tf81ihk21aUL+d4SnkpwYYetV5L6SeGTxRwypnN
wXBZkruP2LMOxtZAxoIJWQBKZywBwuJyhy5RfqF67CMFPk7G31/EOMlcnZcFIUUNjDmE6qDA+K0F
jRzR3rdPBqre8ZlDL4ryV550bmDA0PUmBi81kHxm7+VyrWLNQWE6SyG4F9BXTY/93KN5qesAk5d0
5+9F0yKT8Pvpp2CR3nIsekB6aCIHRhZTNJ99/RanAcjuxzq24mmvde9pLrsSyX2cx/BhwLfEg1gd
bgV8o2Z8k4QjbHgSyLj4OJ86Fl/I/TR1P2KgGX9Bsi9oObgYnlL0TA5yzb91+LtDrIRSK3vVRZ6U
KQqLIUKPo3CEUa56xXhq1y87QRULhRV2ZCb9+1T6bLFE2eyYajPfpMZ3rpM/ZJq6a5RmT3j5/Pjq
8SVe0JJoCViZRWj8DFWECx+1umb0c9Vw0tgIOU2ELyEb0WwHVSyXmy/gaFNTMAm9ROf621Fz/5Ow
d1t3ljguv3Gr2xpkNBXfD6iDaz1hlHke7qUqFhdAnkuYUOul7I497cQ5knXQ+opAf2m3q0VCSRo7
3N7c4qr1LJkFVWXfffScPTs5g/KAKcJAp6LWynsyviVFZBW0cV5jO4RlIIi4LvFIjaUrje1xnoCF
KDXFe2+dQFXhqgJU67mKnsXg5c7LiIcpQS4QBzMqhBeLi6gdw39uIj0Cx3kluwSl5TxpHmfW+g8A
1fPzJ8pM7MCCKVxw1/gzMj5QvQBazEYJleqzYbrgnNs1T3jEnDvAqlwZ7MDchGLkoJA5iroqDhha
L3XQHnIEozGHq/WkEsgOStTCRR7Zf27fz3oXSN5WVixqijdVi2NHoe56qYYIyhaBr1vZq/NwH8rR
1xxl+DBlUpzaHsdV4BEhOhy1jh0q6h3NHPiXv9F+tr/tdGO+TcHH4E4v4kOIeCvTAV5ZRv+7t74w
LAq48nYqVsdefXt9Y5oezt7fF5m6fOSai6DMIwAIpN1A8EpSSWG7t/T8/wTedDhrIbkhh9Zochp7
B4P8Yx7GIYjg9iFpr3ezej9Xc/qCqttOm2ZGuNFKKhmTcMezeVsr3c7Fuj60vGnoEazsH7NzSieO
5uGebrEr5BfY3y6CMSzY9GZp67oMp4ExZyri1+yur8CLD7Ra9eR6E0hEFwLgS6xAHCAFsylLATse
nAoOjEE1yYBDj5fo+pDZLL1Z/99xOO1JKtqNW8Xi0LSAJHsAlzORs6LMxRS6F8POdQO6Pkyp/dwO
djyEs3aZ1EwMBSGFp1NQVU84U4TImjms6SmK7TCe8BU0Pa4hT/OyQZlxjZq3FHePHshxRqtoX38M
Yq4MUxiI0LL8+VbgZqzpRHeAV9ppuA2yavRF0jlj5LEaxNUEWb13QsuodXj9NcOAC63YXpcUxgc1
4TZc431VTwCXXtdpxbH4Pf5LKSGWY1rUVaSXzjL2jcz4hlD6Xcp3WR44qjPC6v+hojypD4n+t+sa
4IVdpKd2GKYlICmKwyHkM6V4CsKFH1XYfnPQqI3X/nkPH1NLDTBsi0GurWpjTCCIAkVFBlaMQrdK
X7BcQNoWRZgS8gFByNm0kToMaBrcR6OEzafF5Ayq/7+76ZnqFIxuTE6WSWjKMbMxUBYyb3gL4Xm+
MV0Phv2YnS2ZpxZz5ZIcJOc9j/A2Z0haYMKfayMR9LiIUaYuFNVvucxEMdSYfwjmesDbKp/fHTNL
vxovsbLhfcogm941nd4el3YaRSFgzf1pMZHXALR/qQ8cCNyyrbVCei6CxIYOs+a1mHLPsH+ZS1wO
rjeAjLgJAWKZNWcGgPf238nAcmlKSbMKKJN3nDndhjvKwSflsWRvGPKqRqtqS5ZuP74jALLXB49c
VfGDeS4iaaM5/OSZuNgZx+5odvX8OT/Gp5/GHBtxX3q0IOWfEO2ANGKLwFwEOAqnC4y24MQyq7XK
ABUtjwzOK8w2fAoPdauY3GHGd+PgplHK8caqADDtHci1qT2OC6JUHYpjMVXko/v2vcPEzFvQ2AOT
GTydSJCn6R3fTAfzIfX+jKIrsd9K9w9MVpy1RvOf6/WHDBBxw9UfgdAsQBJ/mzQIDXUutuPtROR8
BFA6e2gStmS4NW6aTI0ykaw6zwOolXGJvt1kicnMvrP51APxbURMv9QkU7VufSBMF40NMluXHLY6
X0tu5Tk8VfFSuQBEzESGXWgU4TZDABLDbO7hIjK9d6lx0JRyqU3sJXNantRkpD2s6y9OvMNF5ALA
NLiOThKxqe2wD7b9UsrcRg/3jsIUhhu6D7J3ZB7iZbFUhvqVCKk8lrwrkxw8PzLJV8qcC5qBBDu5
zcgf8pSLuFZDaQhsZ9YJ03NEe2ZbqtnTtY9H99B0KKDmv5bT5yQ/RCsAFMd+X0ffcf1BWKaL/Wfa
qDMpyfFuiaGjdYErj8ca7KvtkErUwCm+OB1rnN5r4KqNSkpGbhdNF/09UGXNTycnxJjbRcpYp7Hu
0RSPwl1XP2Xc+9tt5LJAstavSTprnym03DEA4DqgNVUaMOw5g+fpubn/gD3mJvg0g829+vKDZ/+B
3O+t5dGWBGGqIy8wF7wxXnQNrbKy8W8ORjsS/EtOcQ0vZ8wZUmk6KJH+DWlijXIVso7YZ6OKw7AO
HUKHsNC7mhK5BRF13CWmVSz0gX08lL/UcCm857ux4HWYHqmnUOM6ZXn7l2fAEIph7gErNay7XR/m
FDCW+FQSJAnv9+qsnR7g99M1vsHwd/gwcPZys3aLCoQgQkOxN7BjFPa5kcVBsEUE+AJIc7wj8Ve1
wzqYGrAjVhpgDtRaAg1+e8QdQqFl4Rm5bYAD15vTTObcETk/xPcuTrg9Q6vAMWrqOvROsnL5tblt
8TdDUmxBnKe2qBZs7uFrl+QpadKbf5puJnazspj8LOanZ8nn/0v5eRRYduF4cRE98LC0TO8cBGA4
eHyG/Yw71Blm7Iy2AzGR8TtoVZvVi4what6z4MBF+Ty/yuGPFXMjQhnkyDx56viA47qUoph3rFY3
n9mdDKHYrol3Zo5ySAWbsGofFSp/ch+JXBg8tE0a3ulsD/idsW6BNTUq3TuyMJPlw1rsS4k3ip/W
pJm+o520U9zNzThH/oPg1gnVHAseLtgIExMo3jdtcHznJvXl+cYM4NujXv1xYuX4ZtE0jyjt+VK9
+CD51wwicp/kL5LbZHHz9LUM7q2+8ZHLsK9E1uFv7dtLq/BzvYE662lvmu3R75VUK6Ms3qxyd9B+
/0HQpnOOZ+bogCcg897Zw+xB0KzecfGewfSxAleSgdhwvyvRF9tFX+YMb4TemPWJzNziL8yzXo+E
8L3lj5AxyJimYrv/ES3dw2Gri8j5rQq50KeviZs1s1VqkD+WyJgKQA1xf5rdm3wQFr9tFX2nZX54
jQx6DPprNXo/zDLKyLCdtBzAFnC7cVDFzAUtOtnbkfEFEOMxQGx7aa/bIK5BcdCYQKF1QwdLxQDz
IGHrwsZW7T1xkgEcgANGALLv3jWxI8ll007l4m/K0lu7Iradn48wvxbaMDFl6Q/qd7szUBBRv/Tu
p3rHhRL15wT0IZfDxKCtgbRGUcjUA+uQAuEtc+din1oIMzu//hEKbqdeZDoJIe9ZfnHlg11Yxz9x
ngAOnvptM+P9YJ0WE0w2R48jfUbbGWqj8vCkPiKpOS4WVpXIRbCCWbK/NncHU2QOXG+YQOxKGSHJ
8q1qN6KZ0ehvf5AXKk1UH4x1gRGAhyQSSnLlWOMauuLT286xE6gyE+zIG294h9n1tIn2bz19OVSz
SjxOtcTfk8Lf4XrXpl/PHphhBF+7ZXBly5gYdBH7Bk1hnDNrxn5B2KsVpWlWWzndjf/ir679UGEh
t0osxTtelt3oXxYy83gbwfN/RC4gyDaX5NTxqYw6OHsb0YQPAQixptzIM0fMjWRcglmADLDgV8go
2C+jS06Rj4BvDkFHSOiRfcajis8h9ws9GB2r+QNGw5iw6HpaIjbX3jrpYuSjH72qkWuc4mfZNJMD
L3X1DIZ+sq3nZgDT+ZyNoJDm14zpO9JbexknCdcgUnDyAWTrg7o9Hk/RsTQT+cVp7KDoC2nYL1FQ
O9gCTYFA4Kk9IkxkRzaH71oxuZ0w+cUbq1UWfX8C5gT1oGzzfn0BV0h8e31ieZk6WRXCseAhweBe
knSCsCzuDAuMjxA1/IY06s01OT/Cvi4xX881i7YGFENWxD1mkfhXYvY314FusZLvcGrWETA/GKl+
Z0IuapHZ2qPZuJ/eEhCBEL1mFDgi5sHwO+xVS4qjJaDh3YPdY+gUK8h3h6bsVlDtGOfGBHsiULf5
IOj4jWtnFAjYQRNCZON9zLQuZp6DE68lfssFX6dNc6+t4/xIqG/dckBNoZltCqZGEIH8l1owzqRh
UQrIOrrtWcFfY/1IZFOxN4V1MCf+Y344zpmWn38uQ7UeOBAYoPjwXkR8he7/MpHEPcQJw9iGpJWI
Y72zTwbODqAkOb14gOY3arO8tAqR4886wcSdn2LXkQQddJf8YgcM1c3xICesMDXFedIHTpN2wUDV
6UZKCpfw0bBYqosMhwhVLTNFcjZvNtIj97GVerOx5BEIC3ZmFc5WXEFg0vPpcCo/WJW8ZwExEjCH
lhrhuDRPPglpUk3wyaR+3ZZ+Vs1DMHbOHT2813pRHlX5GcMoG4d62sgEfbz6we73Ev6AMW5NU3Rq
NTzwkxKsdRwSGaUB4EpznCn2R9CwBPUcsvrrpHZ//DPNLcfd1gzgQp250XqiErFNMjhGVC8XhvDa
sKBuQEj0laDM60CxA4dr9Gc37ckJSf2FMm26X6SPG+KAttq2DNar7iVd1ndZInKQqLlixUe8EDDt
Pzj/VBUVU+JALjG9TYsObw7G6ps4Dz1LbniqYQa4mb+Wu2alnOJdiw1iKR7jk3Yg9KnAw9pfSAFi
q9py4LqsBYfOtMv01OS2xZDH6HmVB28381+r8bOcIn3/X+URhtyjTrQAE8Whm74rxVR7FJs7jX8w
trOaiEzYnxRl5IFRdUk5ogfXsdqBp5z9blD4D1+m8YRPxAH0DKVdPHqmaEo7S4LexFP8hV0qb3xv
Pz/RY+4+SnRFTHfo3MTwruL9a4QT0CfQX+eex50uas4Y0dbAY0wCg2YHZ7qOj8S69h7e00IB0dRX
YDk59rRFHvaNK3yQHFkqS5U6GNpmQUkH+MWZEi8HS2h3DFdpixj0kvOmWS2PqH6+mdzN5Lee+mCZ
lB9pyoDhGOBmkzpwSEphu7Ho5x9JFLLDuPOo4Kp13ZXlNwh9cgH2VSGhAeQ1e29O+0kCvu8IHt7w
TwdVUh2pIVbX4OIPXfkBWVURLqGokXamdcZeP8aPE57NcxZWFoJC2ihYjvigbvISuOGBm9Mekhz6
5tLWuuuPGuaDJCNwCbeKJa3j2JRjmdmx8VfudjwYQX9YnsqLGQPdO9tsrQG62KsskWFoFgYdWx00
IbjcInHS3eWVi6Awp72jPuLa/lNf8AlfnUgmdj7bGJyNAZKMUm4skS+aONyiOK0vajSYRToN0A/8
Ka3hKMUoW6EUxQzZlq/u23o1U6GexOjrXGnZvSVWOHS+nPbTmAhFboWzdR8Kei1FUoflLxzPTD2o
Vn87abIcT3wxCCA2GitQFbTAdXps4GpF5aIFAxZ/MsI0MOa9KCGzz5eBqh76TX9BgO4yX4IK58T0
4CWHmT+6jD4HcsWO4vFWGeIu0WL9iAYMtX0yc9uw4fPcilUSXH7B9OT4/Q/bZNhj/o0i/I6Q3enc
DvojKzE7+yH2w6ccosA7rZUAIsIdqzBxZhqXMw/MYZM5iby6/YeBzLSDlnwxYCuaoSVc/WhwvwOn
djzryj2feeGd92A7pJ028fGD1pg4oqtbNaVHwiyrBM/J5FjRRQc/LI0Hj9OLrXDh2L2xWnpULofD
/e7QGM+BgecyGu2gC0OoeW/uPCrTDBrzzNOhYHY/M44xCQ6aiunaTO+iS47MkpJxLrmUgtG6Y2En
UciFDn5+qrVkdb4BpzlaSQ0auKaEkeSPieqYyQmaUvnrkbrQ95zk+QlF2HCo8B/81o8dC9cJW27u
U7VeeDZ2JTFFv1SanYRHqKlxLk2uQ52I0qtp6987ekZ0jIN1dgCsGNS4iOY3L+xcDlW/ip0wkZ7b
47LsZkrdIX7CyGh5ZUYrs+1gfzQAwO3f49NyB5fdidFHqHr0ebFHz8UjtB17azsYw17Kg486guVu
x55Z0hwZphqp4du2g1gxpJ/0GrznQuo0R3NUS23oe5bD1OaS8ENLR4DX5ZpZL8ZLEVpW5Dqn7aHz
ka2UZPgZ5oQHJbmbK5XBB7ghLUrzBXtYYAkhXNpH3PqkHOpUqtPIpWKQeEvzP1n1izfkazBP8LJD
uXaNrwvf+ssD8/3Okah3/IgiBUHweJb6i+tmW/O0hv2qWOY94IfAn64I134jRHFyFseZUlzUoivL
jG8PspZd/STP+TcUB4UGdTTVP2it/QVBH1cybdc4igdswdP49XHJFASTwtW8o8oBVNvSqHl++kVZ
1Ecl+RsKjsJv6OrqZQkdbNAIk4vXJrQgBMtP3aErAS7T821kRbjIxmBgUuulXteSEcWpLEfZA8bX
oFJvE5Z8Shf2Q25eOLq9twthWOK1Zl2EiFPfHdiB4uqEbUcdEdfuQt+HAr0SCLguL87SbAG3vmuA
dJwmV4iGdh54/lP6Do3kG9bcMrizxKD8sE8w7R374fxtU7sMwVN8EDR1bU/mhgtOl0CJmSrkhE1q
0ZwdZSL861RwGMWNJsZUhv68p3oPs9WBjsJdwe3PNMIAFojEWChvwl/yTCcwJ3Sj1WOUGaJfOBVP
LHJmBUqVOc3L5ygG9yJ4ZzQEPu44L01U0jr2Df+vZkmB4OHjvuhZ6fEXGdofuDXc+yanorp+kS2u
GtSQClkr/trJ0KU8PtaUsfrGhrP4VTaRmBK+NE7FXdvzRzP/oPrC/egUqbVRhxwUClXUrlgnJ/Rm
1JYs4v5/8QqavtEB5vXUmp4jBtwEteLvhePuIvVOoTuVwFXRJo22uKiaR0jOsu4deJwRWc6FFr8d
9ls0HlAn7nYkXS8vyLmJ2qpyD9vi/Uvwl+ZGGSUN59DpxTPHP3195j3YG/8/KutPyZCLen6FO9Fk
gZNj4n6hf5xQmqg291gyf4l7WBG2L57YSK08Z4eevs+EbGiQL/Pv07VNPrZGf+wXmZfYKFvOeZJV
ISu7Gaus/RHUXHv+PRTdMMyN/XBHlDlOt19990FPUHwTj5sxEccy1hh9xOflnPbGpmmC1dzS6WXu
dBH7zIIVAZbFhX+QK1rR0nolHRoqPSMyHEdXLFkUi9j35Ufkdexl5Nmhbsnk2XVj8rSBV+H8ScIn
TpGo7i66yValh3LSfEUkVe2qfrs85f00DpJrQoIMbLRLa8uyoEzYd1QuKGsoWu/YPNYxVzmn1Ss2
ULcjRlAdBmRbPyD7MWsfTDMKqSGPi2GBNL5r0TH1OPXuFmbECXnIoyXRlfkcI4SWJF4kCLZNdZYP
Yq0hVbjZt1iwzAvL2jgyv/tSE66/mimNUmRc3uoVDiu6KlEz2144/IJbxDzwrZ3WoNlLFfxkG6r7
bP01MTtbmH1OGLgCMGAibnMryAe2n1uvCiy13AzHN5bgbNGrnSa/4CTgh9KYL8AAoohGICNZXhbe
3i77IF/5LUMR2swfk6m805ED+2/cuCjP0ZzABJsRdzQlhJp9Y9TQoTWhB5PXC2xir25TqKDgys+r
yPAcZV9JyCh+smzQsqg+6eqGLxyO4Xf6FKlkTNLVdI5dEolFbaLaXzi6R9pUMUFeX02fj2cK+bmg
KvrbbELeRfA4sH7rYxVL3cSNa4NZZuNqQ7Y/DiWxZ5vkstfDVedWskuIcRq8EytRAI2LRqSYVFj3
6sifgnhf54ndK2nBeT5XofItG2V6GrA6Rk5XKJvzst6xp0U9S8fQADtcgHI2BS6qxmL+/OsLAZZb
LWtaqw49HXeDuhVuZyU42sZkmzCMImpObeQPMcQwHdl9CJocC5YsxOo9lwP0GAhICrIlqETp1G3u
7/yKDLPoKdVzaS2wfMiKVQv9cPUX559/bq8ZQpC0oQZoKy+vS/IjMZX+FmIcXsa1CHWoyjzLGtuW
3WNg45DdUxACUiLS6rjQGYorooOp1xLLEyqWNt6xH9CDnK5YFMfH71AoSssCZQA6vuwWKOk3bn44
R+PLZ/cHpR2OejlB9x0m3BH1xcJw9tWSTgfkggOGn1OG6v0rHx9seHH64O0XJ7u9KVBfWXch5Ym3
zGVB7tIfr43/RHtzQPpP9+3/t7Tluk1XSQ1rx7p1tGLFLxEiOaXCcXX6pqyHYIUTGT6P/slU1lZ0
gaYq72gE4iM7XS4/Nldj6makeCUX4Q0oQIe9Ubddmfa8u0/u0XqOj9oNlLRKEeXyG9/Zo9C46E9I
njNoxxtNQgbmt4nz58SP3++m04morWnF6Ef0uUwQ6ggvzvbZd5pXr4jrEszJEvlg39fUJXgEumhR
LoPOXfMPoaryW+BHul7JiDjdzANsm7Sogv+mb1zO0wLx4/nAqTfy01oTMoa0aAx8d4OX5Fnb6Bkg
jGYAlPcndu7BRtBBXMntZymafkVDaZhGOZm1RntbKrHF3YVHtJBa2iGxhNGamCHIZ3++W1W+mfZl
Oaq+PwShHl+L/2f1PjgXJb/s9lomk8Bx8a2kGB6las5CfJh4NsyKvL8dSgU8m1g6HZsqoUKL7jYM
wgEnnI6UxGYCDQFV82xU08WBL2OB5eBawpSL4Mkla/bdJ9COC9Q65RdwzbL/7xNZgrDv+S8B0wSs
AojmuhBSUaY88qdgYZ+ZyJX1CWSlzKbJ9+2X6EiJCKTaXAUE1KVkN3DFDejcQSbeeGFRCftv8MJk
YfuRQS8kyikhIWErivVeTBdqcC2rYZQjkvqZoSajxynv0D/8LOtwMzUCril8iqmwYVVDs325b9A+
Vz0Lq9LiIGUFxotbTbQWmasqLxudFGCdTOhVm1R0zI9Hyrdr+/XbfkmpS0Nn1x+7L0O4vw3R/xhg
hXwV6ozl4Di2L12C5j6DdaS1Q2ihCgtRQuDkAIJp7Dk7hy7X8L/4w/nonjBtwojmWA5+0KoY7gPm
/YXPuJJsXoSGI20Gb9axzFSuR6YKo3HM5hpbM+5v9uonbGleX3AhkLjhfp45L7J12I0sk9exojzW
C16UgNDaFfRSvNCWFTO6y8g06uaLHzkDCIh97YGf2TL3cAR27m2T02bnY7/3LMt42flJP5IKTGDL
2bjbnnH4XJ1jVl2yEAQtetxwNBUNpj8ltU2cktvDbb8/iFVisD83nPRbynnYvDTu2/ck5uVNbtuD
+kG9TpvXCiFyuNXQMzt37oUYBkWIqe2MHfxzJ5BGIqQSkroxBnRZD+vd16E1xzl0Z9RHR85JodH9
CXaxPav83cuLLMTBuiI8dEotSKN7axNeVUqe+KCd1hqUCx4yLGuwbOKjyEas7EMqTQzJOB7YA2r1
Z6gZvqRUhEo6JJTTKepVBcdocUgYU0aYlAJ3BS1Mgc9Gj4Aas6iVULqTmTU1EBavvsP3eYhxjfQ6
KdYqHSLGR5KifxSgIjks5NrfTjXttJMS80CjseXxfdb59OrmJlTKQ6Y8ra0M4I3mcVOVM9h6LX2K
hv5WixCXBowsN6qG+ljenHX7KPgm/D/QElme2jL1IDtQHIEg0JfTNfAV2ob9SpwECO5pKhNIBmCJ
yTXe5wOJiIITKFLYZeZ3VHIdmotcKre8ZM3B/JWUNWPqSoVRbK4y9HcvFtRQJ8aoxPIq/TDr/1FU
k4l7H16x3WxVvLsLNDrheZ51DiJ37Yuef70TFkyYLwxLxzv+qd9rotLxg6iw0EvOdM4GCCckOlp9
FjEyDQXz8gFpCt+Qi5CqeMr0uk5zWERSr4u+5yR71BlSFiWdFkzTyiNtdC8vAIZt3+EZcmWxxauH
nW5dK7AwD99SBFWeW++Yl/gEhJ46RfTn/5Xf7xt8+enDBW/LG/MrrQYB7A/YU53ybmptkcrTdsMV
X5WtnQnTqUnGW6J3lYgytHGylVxELDMGHSHoQiRMooCBCTjCiXAGAQvaBQSRaRYCyMjeNfkbxobs
StrTNtQSBzsHpjhs9Invu/7FiLLtDI00kHeD797Y4gIKVe6otLI5jSY3uYpO4EQwaZF/FaoDcY9S
CxvERut/tKM7UtAVI6Sql/fukQPmKZur71jIT5gS9Ft4Eziq4QcNw8hoEVdF00e9QacfjuwOz3fq
taCSmISQ/u8Q/QeyIsZdksngKjGg4ZQyDPzfiZC8qYAPVsT9mpMgdVfzi8yvvy39VHkmQVai+M9n
GZkVJMP6CMXBKRyer4TYC9EjQWYccF8VTp8L7a5q+Uk9mbRsjaupR2pxWxhJAgipWOoMEzXtRchD
hTBUjMjGfEZ4npCwLLaBiAkyUyNGrw1CKLRp3ZbcXdYhx3DwOqAeBOGYJm6CM9Dd9Pgv8Wbl35cp
vsCLBUnXanyQDZw/B7tQnfnlObWdgvX3O65cQfDYDiF0eyCU3ES0ILGt7sJqOx8WYOH+xjJ0Liz0
6kb9jNZ/Ps7GWNKqyut4nlSAkmRwMvSfxlYWU6dD1z8tB/mLCon6HGowJhjiUNhrsmRazo49kBsO
7Xefg8I9F545BTT7D6wwsl5r6VedFy9VzrWqpsJ6kXpB8n2PC2fvk0CMWQz+Wu695uMhEqw+tDiz
xgbUD3iXDMoP1J5drtKNqPnQgEMGiVY7NmcRF1V+ICXMjEmdyZdEJRpnLd736Kv3mRR1qpNG3MoX
9LKIeF2xUe6AK3uiIl46GCSQm3LZFERq25K90S54y9GXJvUkUK3Qlr558fZC4X7mw/JaHxNQ1iQ7
5HhzYq2bSsYQr3YtYAwGpzwljjIMkX1hBStsCZRvpxCNCZGYqL2Waj+ICDfjpPd9ymsAnDjKVHUl
mmoRnA3IbExoroxOnl5ReXdpDibQruJ0VbbIkPHP9dN84r5wJmVw8LcarKXnhpkyNPawU/h6SUbN
cz1fccjUwE+/xNUsFHQ6CDlhZWMInZbYJ8siiUZFCODFLm2ts/hvMhkprlMuCEhLeoP4i7epxk1S
z1wxb1Au0GvYqQDkH/3Y3oQ06jq9veHlohGN/SRtPHpBA6y+9iHeChtlFe8aOqLLRIA5XXilu/+s
GVHpMTcHerwuQx6heJ7Ke5BVkkREE0wyhzU8dVkiyt01EyCnJWVAmKQF6udcxJ9WeQD+lL/ZYBK9
8bViKLmSTtjZDxmbmfu4/jsLRU7yEo5iJPfjQe2zCBQfDCrWR6MtEC7w4uhhh0/zbWyvc2F26Vef
b+J6vpAaPlHhx0+sioCuwtDyhU0IWMHU07CBF2BIt5Xmuz7Ut74opKsmjSWsvKtvvCMwieyCNna3
ijGfq/fJVcm+L71GIo1IkJPcHiXaKphbrSlPlmJJwQnd0pto5bdwYoW0I1XNKs3wRIwWTRxJjK01
r7ODR/KwVMWJtR/QFDXv1KHZbtmjejHseGzXzT3PAxr20M1BG4N2+LUTnLcdt5NsYEPv1MfUIeXu
Ct9/bwY3ou6bxOUwOtm0F9dc03ed2lNa8cxwPa0SypHbgMLQGnRgnD0vEl8NIWp4c5CZaiSczufS
FUfAsrB8N3LptE03aeIFslmGGwiBEepdhe5EDg7tmzZ4U2ZveErS0Q4uhDCV/bYijAX/rpGLocV2
eor5nV5nNsgt5ulK42wee3VkeL+ni7q405vckaP3/qwUcti8iyTKs0d0g/xNknyPaPbNNACPL9xl
rsxq5PwT42jk7bAgVBS7P59YJUhDSKFBh8a9ECzPqH4VsDY9ErGPuD4FBZcm+ilaGX0HO+iEmSFw
rjoywhgzP35rVc35sVfmau17SaTB57+3SpLkFdp1/U9ZQbpL7CPs5o5Ay2JNCjXJnk0AJbKh9zdF
OVAj2fPQdKZoJIDZOG+h5su5p2i4i0zthUa90b3vjIs8O6DKEedHYV9SO/IYWl9qxFAWrYCkvBsj
M3iCKIUCziVqwfND+LfUZXzGVlPVlb9PeaN5WUH+j3VxdNq3hpEijkL6I0h+q0Awue3B8NFBkCla
x5JOUWv2ba+znmtyMfdfk0AYLUqJItl3pzoKFI2Bh7SvhwTwdpsy2snfhe3gXdmAlvYw0bJUiF2I
0/vYTH/WMfrCwiVyFs6BikYexbUU76Qf4wtxml3SICrMJbZGJ6MGTeclYzCMNThdUGNikJr0zbCa
hHzT6bSEkGUgQZRD4VSF6mA8X5c6CmADNEdeayfJyeLrgOoWJbR6rYk82IwosUE+mKBGBth+BbbW
xkvwU1dBP7oiWo3rW/AM+YMAMUKHFyV2Mj/fdrWDMzBLKM2RLt9/ABL2joP1T3hj1yxVQJbIndQ8
0qHPnBn3Fd2jckjObpfaZsYwQnf/Ken0Q+6wVKMwdTbBq+Pmdg2PUW1IbsWcsmASyWKacsK6yeBu
iWBkHsVlmimBQfjyJwTEm89uh3GybaAX/Dj2lZEjWZTT3DVUEXnQfWOmRfaMEgENdP0B31USsjv2
saNtj4o8j6JEXIUkswUlgVg8lPGRUFt5AuAqc/6SKuRyxBa+gt5j5OcLoXGjmQr216PzdQF+oPtq
JpPtib9kpPkAF/JuCugVgXIxeiC+XD/F4YxztHrZOhop20aNpoRMXOE58hzgpkiyG9ntsnNwoT3c
7IwBEo6Hj0kTWbVIdOsWOvaDW2yS7azWX/oe7OJ5EyPWyr1vIOsw262QsNniIZVNuMvHS08lRJHv
Av+2AlpNhx2+Pw2SloJyoucX7G6iTe6mp7AFEVAORft9QHnyw9brkeAt+C9gV/qTrLfQY+OSQAeF
H+eY35arVoGizb9GF2zrW7WKiJo12+mDXhksGJDIROcvjHHcCV19RLUrO5OYgRQHH6P3A8rix5Tp
TECzR3X2giN4CdTvSDhXMIR9CasM28dHRs3RUpRhtx/oKBIHUKiE26bRUXKFv8O4wAhv3NA6++i+
DHRXGvhfoH2/HDn4uqROA3dXHET65ekaHVxQt5b72RzqtlO6r4YOKN5mDu7Yan492PmmwpUFZW7P
Mkc5ezdxafy2f5kvYiYGqjb7zKQgWiye8DdI5e1L6lnMVtqgzDRY2UaHzxVQs4T1SS0AFg26P+YN
77G1euE6p217L/evzGpJYh5p4sNYX+EZMfhjqjYLgCVr5U/OtXiVUY9SY1zRelB4gCpSl74cEDjx
FcK79snDLBTM0zJ++PJdO96AQ+wrY4dpKbSrL8/A5nvuntVtSlo4n5th4O6x5WUplPJFedpBD12J
Q23TOvfIdwFnt23BFk8KxYBpYlTswnyO7QidqOS04y2KKSgYob3YOu3QPBr5kz190zVvq76pi5wV
6PTS/i9vpdP6sq4D/4DLJc8yTAijP15SAkRDRmS9ugvuxiBH0vV+Hv7WwpgvpyESw55NSla1MGF7
ldmjRXADvLzhf4LCfrc/cEtTyBjAe3KogmCbw8cOB2R5BVpXWCrqNPNE3dSN+ur2ZCOMi/YzHJxZ
Wk2M01TnFqhLJ6+IpOZoFvL5Mj5pfxZ9Qk+k6e3nH+KwKbPVD3rKRJPmJ21aqgkkYDJl+nTbsTFN
mnAb0rpzHf7l4mXsRiw6NKy8pKGwt9RdYrmuNcMZ+DfY/mZxfO40GJqSWvQc0bPZNfkQpP6RVS8d
OCUUr7FjYUyxpdBfmhuhcEChbsXFB0eEGtudV5YP2cxWZ7lr2JxK6HELpimg59+OrSFrRJXWpP4t
DoMe4UCNmMtBvRRDBzx0H1yaJHrqLcvDIVyuIoQXkkrNMUX8DWF+V+Z7i5WBo5Tf+5czR3JGUNlq
Vvm88iUusDHGJnDsN+mAxkbdCLQ2/uJcD0yEwOFToPr9+8olPMySIWiqCHQGNptISguXAe370+Qf
1EG0rjvfO5xQ9TKwtdqdcS4i93hYtcQtyVqvikGaU9oj+97Pf/e8cd+og+bVF0UMQA3+prNX2Ezl
pIs5Lrm5XlQtgqMHahTp7hyNiTI6A2/figTtjMipwK/y7GBAUsAsrw73sTHmjHvTHEtdIiuiBeUO
45g3Isb2n9ohKVjlXtfBHq7zLPYMNnG5wsISNNMsaZoUdl7G9Uo881QKdnOqu3i2sMfe7KgIXPpj
sz/u0y+Pp/QULOu6mGnfg5cmpuDboBWNflrUKuJ4shcam5O8OYegiesNg5FLtfDKdEC2JcgCb5LZ
Gm0vNE8Yr3nBbhDHXPsDmCe6kZtLDR4Vubvjq4bULhpkxDqUhPMlPeHaPUZshR28CP81J19qX5pp
EYkzdpmulmqcagcitEcVT3svDk0qrDB+/Xk/ZSxJghZAAaWHU1HN9dLOItzztNOHDcV6XIBZMicu
4S8NrPLVwO7G/4kCApaUvgXV4IBOlgMBSOSC2mybGW9Qi926VTqPcpIvdaWvvCicsZ0FBxaC6cmf
lrg8juDWRph89FBD3UUEY9Aeh/IwFpqLhNFBep40oz0AnL2vb67+f4p2OonfAPv4Q8YHPpLj5S5k
+1dG2+42Tl8X3R9N9fkwJX2zSDHe7NKSEH+QY5UxfmJID4kUaRswZrCYTVafo7CCQM7VtTbrDbyT
9XWmW4896ECSrP6/JN313zyQ02kBSDEO9k6nGt0SX1CGkU+JzWccR+Q8BmZAnzJ869RCW7lM+vag
/lO0ECg9SyUMCndWyLtyqY3SfoPlqSlUHZPMlqRIjYiRxjxW7HnzV0cCXCN5cbPur+wTHINrqg5t
c9IGcaz37Dz/+z0khlIGxa/cC2fHovBdxm34KCqJrtexcLDBVsGCyOCk9BXGhy0kZZnsGluGkJEK
ZAcaqsSkOC3lZ/TBZSWr4mXtPVcnuWnOr9hmnPiGncGxBmV7ssG0ge/9dHW3Xu0t4YrsltpmC4lN
gIKsnoTLH/AifU4SY7PgR64C6XQtHxXvfeOt87z6BSxQHDD/u7IEtHoJlxVsQ84OGOv3XBRtAZH2
EeVR2k91Ea+7eUYCZeexI9xMwY+3Iqv+eXYwLPW6NaT5Nbdlzy/tbvUiPhb2B0dH7gm+uybOZOT/
9BMRrmxtoUTbxxmfhcSgM56S70ZNKB0uovxhxqvQUGUk/r2vGADIJ4rDGTjc+GczYQgo9u4PeRRV
w0iGogCfzkVjfs0yF76KKTBPLdrGTGafsgu05RkmhWMlzeVTtWHMMr6xa+g1NL6rlO9I7tpvAyWq
TWlVhW348PO4bBgU7Ufglx5Pn0jc88YjfFQP5CyoD0jymkiSMTBVs/Ft+dXbAsjqu4UKKOtMGNd7
a+nNBtf5ligI8vOjQYXJSbDJL3YmGAV1p5ig/VcX57vfFkRjU5zSRMfqx5B2QlGxl/fWr8Le208F
2SsNR6gnvbHyscGpCPxEoKqxSNKZVjxS0orJwiILg3fpPFV1jRkIGakvvukacTYUX6LzS0qlWmFH
jnxnAu4mrUdS7F0C67g3me2NXBVwv86yNx1fJMhe0AiHftnv12nYUQ2gIkzil4TNFljdKGfFjMgm
PhtYoAm9qYAxqdPXVUSQ8kBy7/FdtXwWt7f2aeoBabkGE7b5+rPjOs/iS6dlrHpp8YCIQn2t2NHD
anld7X9GrOKE2EhdITracOIn7qB1RyJOVXwua06Jf6gSG/eouZzxKfcnX32XPEJBlHIAPH/R7d68
fOijd8lAY9cp7BpGO14QFAtKcRzFQPDMRv85K+dJPAa6K4q7XcrB7+ODQMAGQKEprmliZEQPdVT2
EacofrQA17KVEj8w8UNj0i/6j7ArMzeDstvP0Xzbke5c70cLF4RINBCDukTJGqnBogvVHFnR2a89
hZwW6BmXQsjvgJzFBIiBzHwt+gUeuuFoFYisjVd1RPWZZ0e3WWiIux44Z0kbzqWR8BpEIduNJy3Z
fWsw+EhXyEd8VR/7rxgOb2nHXeAuNJLUbYBoF/J6fhBfmBljJwI2liSEZmQzLq/bWVH0FI72ZOpA
8jSCb4Lv0JIe1wATQ/5z0ssPgszbxrc5SF51n8GE5oxlutXy8RvuNrwsnhvRiXywMJ6SITXdrqBe
asycoRRSRjloudg5f6O9HvwPV3nplJ3v646ZN3T60rf3OvwU9pP1dLj432Ly6JEOQvWdwT9iC9lN
V/celzBN5iuMi6SKtDhhIJQjjQZ1ZsPzn2WCQM8RHq8W4Kzw8iOlYyLpbRF3d+wgQ0ku2WSnKb25
M6/rfY4TnkUBf2ik/q2QrDuCLFsrhrwYvAsfTc5QxRLkvRD4MuBpidWvNnL4Out/YLeG7HXvHuoX
lOQqnA/Zro+THddsTyJcb9Vj7DxE63Dz6mPLsjeN1OU0VAj1MTBeMQDVobj395t+0uoJpnkD1XgK
dXmibjMfMbDMLTAXb8+j8mggq0XO8raB2Pu73TGESZuhWC/Y2vhRJw9HBquYD24M3ohYWgbNZd3u
WH+zedkp+wXjT3bAHJdRHQK9XbUZ+aCnVPivLZ3AsmbBPtJIffgNZxbpEam/AXGXUSxJioyV4/uF
Iyfh9HGoFW0iy4++iP7Uw+r5gmKs9FwgFSDxFFV0avmgCnAOMQ+Z9Yo0HeLL2c/iza+xLhfl+QJx
eflhY7x7uHF00O4FXCO9HX2/HCgv0zP91oR4MgzwDYo3PeeikOIV1JqZpj4DkK4OavMV5QxUnyIn
XcIAX1RIUoFjz+aExF+fmuite1S4Fo5eZWBvXUMF2oqwfPUG16y8dhmKhYf4xm+tn1H5/XZ/zFgS
2ciiWgu6akKQ8QN/7mjtsNrQ5VTOhCC+BkYp93RXlC7Mr3x3jxsv1AkFp5b3dMXIW/C3AOL5yRLZ
w1JW0nSfxRLrw33tD6R7xxm3gu5LMukxCR3owjS5VoIlKblx/5hKJP6ZQYvM07bwWgaUKPSga5AZ
7iFf7YNjfYATPbgsaAL/OVbzHXBqN7t8FmEqQw8GFt14F8dqB5LtTPc7Y+I1cW1Pv5EYe0uEIv0R
Z8RVnzfQ5RcXNkozJVp6zTbcYg5Q9s8dWHAG644Lhz23TAnLDk2PMhkhiIqM98+9neg1e9kH7tJ6
dOKq2rkVcQJ5Bllz3Q2rKkwaHQq/0K0T6zBlyXhVWXCuw1VAbvVZPdGn64gSSR9Ipx8jfZJ3mSu5
WQ4g5FPBnSZ3fdj+qOEBaF2L6d44F2yWZC0Jhtga8VYh1K89k1xu2RxTGl83a4rp0B+b6X5Ftg9Y
h/Z0ipf1WLUEfPucgQDjPsrDb7cZ65bf64Gzq9fJKq1XD/sQkns5/aAmsE2yoGmbcEhZDGQc+Tgq
W4rnj45VWIAlIaNI7AJvPUZThQe7hoK8gJ7ixQqniB0rr8E8r/eUm4mPHxJGslM5z1sSWHNtbL0O
YIZWUWQm2pkNAt7Bfc7sOQIxvUUga7zIEMK1BvGzV3b7WThIOmSKQV4fz6AR9e8+HpajNdd8b5Ki
UNs8Zz5dQjWEIhC/BAIZWXSSpYtDK5omUoR3VpkyEizda0om4zYTL69DrEgi51R7As2NdvXwzi/V
NFA8IktUlcM1D0peH4g21FI8aazJCnyqj6VL702SvY3e5kOVy93CYDmOuaiBebt4NFXQ22cJWr6F
LBSHQ5Ij9BXN5+b1QCjduO9Vzhe7poSsZkL4YhOeVAxSFZiqVpvTuTzgBQb6InYUqm9lz2C6AVWh
jShBjhW5QIze0jXf7423+8765S1TiaOTX5JfK7nY2MnJ80FrKuDOenvYSHrakutwkGbJ4EvBOhPE
5U9OD+aSTGYdviVJTuqxKGPFDwPPpgXMYUtyX8yZvlEUWMGAyYY3Ml7d3iXmFUkIA81tD+sUMBwG
mNeXeqJclrf1Z8Ns3a5jzGPnEBkVFYKbPXgwC703nq4oWgekc0o6hdsf1TLOqj6jUK7zg7GSenuL
6HwhWg/7R1WXW5ls3FHBr7ZbhJfE8GmY0cYGc1+R9jYEPhHh1KvAeoV8u/xIqlahtZpBNW/EzQFC
g0pHMO9LQc1lAQsb+Gv0+C6LlmQBfYKksQ9RFTZksSGdKmZB0epLxwwfUYioQNA70H0+9QxSWwHl
yZprWStzRB/n59i4kMZcS9g5EYeYEE+0JlRVzi09/k7zRpGjMlN+kYqJXawtFi0Zq5sPYpxA/gFv
PFDt9Dp46lpkcfiQU5HMo3q/orekVsdYorjwZVzNP1JnlKNRpHlfUgso3KTTwLXlBpml0QeSG9g8
D9vQp1NL9eYwZwyJSHnzP17FEGDqIq4bLWtEZEMdAJ+cGgDgnsjedMoMNtBpNjzaz1os4m2rdYK5
AESowCUI/atzwE7lrp1KmO+lNAxgZHyer2V/IpRPVXPeuoiRYJHM2Tp3DP3RLr5BNwo3tp5sTUtu
qF8V0ftITA42rZ23TyE+OKyOqeEpuvxA1I5FOFIYs6T1Ejh6wavn1T0Un3v0ghM80h+Bq6+ceFSJ
LAkN6d9ry39AerSsqg1KR0XDgHq8lHdnifN6ZMaFWJ7ATVgmUfmACum6Csc28aaGmAfhbdHb6ui3
P3CEygpHmvc7xA3Y693UFFTcmwSyvo1tN/EYEmpCCpkQJ34Hm0qUqlxZ3vErUD8JzL7QZlseNBn5
29qZLZXO1X4sQ9KCDL+fMH5lhd9KZVLbgFEbREVZUPjESL5FCdj0EUX86s40wB49JO+c0wy9dLuI
elp4gaC+k2BonwOkDGnAzqB13H+55C0GqTIvvj9Gb5vF/9AMg1JTjqong3KTnOMh2QG/tqUrq7gF
BToql877hQ7v0rMGohtGGcF5iGcWjjRWzBg73mqBMSAorXxrEqP8TWf7NV0qjcM0v1nKYvtFMb93
D00wjAHxaiQ62kqphtrv9Db1jobi/fU5epMD9pd0wUeOUH7PKP5oEvRu22uDnGwPuKtrNOhF32rO
n5M0gB8fhZMF9k0NYhUmg82rsvyuCMR9yAq6VLRTUdg2Snv+ll5Ui5twV5ezyCcahfcX8Q4w5qXt
KB9yl9FXNLg5XNVL3xg+jovz1930+g6f1s1fA4NxzA5FMU2fM0sLej3OhawZ0V7t2iihQDivIsL0
K1QpRbV+XR0W67LKj5uqHkpTs+5HraeQhpSs4TC822/wNjYtvEMIJ+22UQwRTM2ij7UgZ0fKIEOm
N7mERKv+lzmAgse+qptI7p88QPJ86XirbwneYmVGzxm5pBV3av2MTH8blWUaEVdcz82oZPVDyk2j
FJOgVZIJxRwcbaV3lt/OKlxm2cyv6DDJMLxBVP6ogOU9uhhbh3w/pRvBruHeEKJnmsVk7KtP+rk2
3jKGJ9Kh5Nu5AVTprrlVtGf9XLI8KZof3tz9HmXs1XGZoxqWVvCQFWnBAdYcNmG/mUXfBDWrEU1P
4fgGw2rIoVqdEOkroNWgPGLI+Fpxo2yv48N0hNTRfjRj000c7P8/O9wDnnC7+IVjoAG5payi/7cg
d+tD4PvCtfgx8bgnwSPI0TQPF1GAq7DKjkJuB9XBRb0nR2J3BfiDaOsRfKC00T+p/zjLPSt8nt4D
V15iaNn+LI7SsAz4wAmPjbsdOHce6LI9xyPAqfKOJq+E/FdR/cDHkikJi7KWMyOFi/7GIXYCF6kD
+TtX6X+Zhk/ZJEIMer7MG5MxrVLrt/RvTXGbTiuEXDdXZpPLkw0RChRLo2AXsy50Qxd8yfOqduNG
BeDAT79NpFjwsVGJ34ue/ighudnrb9SLc5Do7QohTv+O8jMzPuh3frOM7ZzoRyQ5tIIkgzx6UP7G
x1KjSxDOEEBSB2Y1Hipyd9aAVgJY3Ltx3s5hfrgiWh9mlHaavVjxDFw7rEJm9/6MRY40zK9W4TkY
PeCuHJvqeJ/bApCCdDmn7jBiw0wrScSL/SHcFEieRM+KG2dJPXV08N6NXTsae3NhCU8n28npUGdm
YiNnfbwo6lN1QdlbZ48uNfqde1huxrsJhZveSiRNnyYLNMwP/pnE0vV18iCCfV1svteTJv8H499m
Wd833t5VLsLAc4E1tMaBD7MXPMZbsbNgEZf9siHscbuan/X+aEbbQy4W59R1JR7KTBlpXHsXDfaW
Sv+TYHw7VedzF8V1nEHD/xUmSMRUlE/CkvuVqdGUGbJeInbLwsyoMSxh7J4MhI2NBbtsxqGgL5WQ
KgOkLXMx4fNVFVh8QKe3qiMYv/w8zFKhVZ6Tkt+QabLxavzoahDw1sYHSIZshFtkoEX1NQIbebzP
6yMuFZ35NTO3Xb82sv/c+Qb0LXq/z6FsxXcneGBf2P4HX4/zEYKGkwbtx8ovj2EFL7k8x2SOKScK
1olDDD5oR6b5KhNoVi7ro0lwKzbQWDZVuJcg65TjN8sTkX/YNTYJaegyA+bpaYg6dNvXhgUEXgCE
nqMgYug3QmQyb7dVV5hrZ+hylFQgn2FzLF3AqtTzjX48uJUn4jRsBpHe9/k6SoET6w4t+cEhkSWP
n9VLA3jI4G7EuN8KUU/zRMGnvyB3H5CB469SUaIg5LP5wUVcRqXOoE4aKkZtTLEWvSzM8gcGhIDl
EkfmWgrtgDKlpvxpGj4x8zyOItNm3m7rL9nJpFO32w08RS4i5XmtMoBFKRenYlqh5zKGOkDl0aYt
iIfrllQpqKDq3Czq/Tsb1sBI2CTT6ipWd6spuJR4elB67qZNTbc5YOO/2PmoIJs7Tu4e43WN8O1C
2+mniRhoMwSPAExJZT4LHpHCcwqEzPrVPkl3otipxMFQ8owMSWAq6OEAdpSPIUIcHmITrdwPhlBV
QOEZV5y/6NZ5wuXVU1+kbQ/S5lYPalAH35mDkwbB3Joepizq0FchGNa2iWuvraBtdj7UikBW872a
3FbXZzo3pb4lpo7WaIC7pYzdRs02SRvAu+/1+GyqtO1F/mnjROmgMMs8CGVFynBqd7NVUCBkShKL
kGAInIMqnXmvHY4oQatnkY9VeSmYltHG4tBY/WsAN90vsiKf1s114ml4wsmZluqZikXnPPOXvs1R
DdGl8UELvnNDtCSUtaQEPX8XyMz5UFdMn1JAW7DkEwrzY1Pz3ndJ4+j2tWjq7F/+bzQtcHJtgwty
D7sO88LyV16F4PJtxaYOrwNxmdshXE2+hW03jRe9jSK5gQhZChVAC8gniPIT26gXzyfGgq/huuvK
mC8vcCbcp11YqTaFXQyDLqjx1EWHhTUBHwyi2vCocEuLXUy+Ab1mWIrKgvEjJe6o4j9gUVBSOV1X
lSjfov5ZVTLof2CJaU8rcbVqW36v08CQGkJiHQH9k0we3XiCebA0zj84f68OfAPXXnllkQEtfV3J
G62JH1N/fiq6UJBYQ/x/+Pcu8kyID1Ev4w602ofhzpee2YA4/2c1wEbY4ax5j1biwD8lUPt4ZG7X
g1rW4fDu7QQpUDmHpN+zNMMs+vNLxkFpEBnHF5HCQN3/zivQdCZA0XWN7SLvglUQncmq7lkrHzKF
vrKkplwH1SgcyGE6AogmlJaLBpRwe92P6Fnhy/ZKKHVJpIc0NZ+rkZM1VSz/AUKpfhpRpLgTjbnp
27CMiQOE7iR5Zr+9z5+4Jav9P2ZvDkvXe5i8Qb4SriKEQ2OkK66VlxQ90Nuoj/FyyQySlTu+wTuh
KoBvDqlnJPb6kSz3SAytLxwXaJ8oXlLwUqbe2ST1A8vH4qxfrJ3bgDFaCTAkYTrRKwgzWRCtIGwO
NhZ3kx/LsdAuHg//OfyT5dFG1uEdGDAVxE2ldGrWaGHTLHDtFVRYts8hLnp0aNpwVJl+ut/55nse
6eY2NvuFs5j/e4crT/6bw1P2JfSfjxC1uhVDdcQtYwIsmGuKq37j/lnF7QDkTmuHIUyWu95/yRsb
QPwJOdfhQ7Q5Kf9CXDBObxHpRYDixsYrX+1W34J+vd5tkp88PlIviamRG4paYe2ye2jUphroHxza
lUMRF2jm966HHNF6SHRVah3ZH2bugwNG1EW/DfBH7rvttPPbiHBxasSYzr8B41ZwTW3WRZknWRI3
RIXMAucf0jmhYIRlbnHY0SQZfHWH4VHohGUATQPxQyW9IwPLpE1DjQFya0RP7XfLz4C+ZEjMwMJs
WRasdJ1l9ADTC6pCJoEQmqFcYo5/MRADiRll4VvPcJABEVCtH8mMeD6cz4p2b8//QYzh3yApFRKq
e5os8Jvh+3f6BXCWQsqQHRCQ03doI1XUDRGOqn/GVTsClvzZQp3jMQzDx5311+Ity4hXNhkq8JFh
YmtsnT2+jWrVXeZlafy1OyIRWZkalppMP0A/Qig5s4Fs3qKZaPIeMCrUS9CgyibGj8JXWR4fsHOR
0hA5HTDxE8PFxpWduc/BGDwNNSWw9RgC69RyRSRH/TIHyKVBmAsEKienn7EWQivmRkEpZ1nwAYxP
rT1DHFlTFu0uykMU1tJGibrRAxYhHM1iQK3ZHwqY+Qm3Bw/+9b0jX4fw0vOfr5SxWGNLLzd9Zgn2
GNh0kMsAv3EV0ZDwezGEhFI3N9BXrNewjYXFBl7AiYF/5fEGf/w/nkQyvRzEfThiLl38AQCCS9/l
nEi5S0LXa4yTWRU6v/ckgoulqlO3uGXbpynVKY2op/kb87U+8qHuILwf9K7Vec0DPc5ZOxD3JvEL
NzG5pou8nT/UPAYZyOHOh9npNUDn6v/Nr8YFd6Ky6hnrht917EHwMIejpLx+3q6tO1Gb/y/mVywH
dHjuz4j9kJ8ygqrLKfhxJwdq+LgI07M+pPdhl2A6v+nGm0kTqdbTOEfDYCrgSgFFQq1TNlzhwTO1
cDzah40+z4fGNdEEfDuWYMfhyakRNHw22ri9JD+PAdOxSVoZVj20FF4FUN4QSOmmLLV2bSCS0cPG
SaCwisbPZEv8RFFrOUfmlNGNjSYcn43T/SPqX9BwpviHQ2igHC105nQlhaV7LGWqc/7U6peUd4Q/
+DZfcgCDtjuxgiSfuleQxlvwWIhDCIF8ayPqjwQKU9SacFnFtCZ52TmDNlyLEZz+wNdUP3PO/kAM
CMxNfyW9ba1gbq0YagsDDJhmgkLW3xqaewu9YYAikC0tKWlgAQmwfoqzGo+FT+tlerSIlq58mPZb
9UvnVwJKO+htzv5HaDsXAU6NwdooffsTDL1Ld5hUCu9uld8++v+ObH5VuDOL6Dx0qmtBFfM6jqSY
rQjJ417AK1ArMHWLQNKrnjcziR9EM2yiK2s2/LsSIbmBgiQqT9eCbzVNq0YWlzd02ncNW5CO1W1S
BvIxZITCwZIQGsOP4/DLuNt2DBkCFEob1F9PWaO8vzZlv7/BdVmc99dXWdyFxi0eIA2Pjel71HsI
aXsMOp6b6HBIwr37vlqXdJjrOR5B9ERwOZJWJq8YimjSm8YNEgpRbhpLQcH5cs8gK6BHmpPVK3ku
aXJxawt35xaGhU1AcAOjar2QFctm0CFbmIBz3P4vSNs8rhrhM+rb47OFH7HHMzUjtf0ta1ruqZZv
HWB3jmZUvMkh8NV+tucSmsPieD/XOGoqK55R0M7QkLRxw7STyUoNX6t+RrOgu8I+KbQdbwhbLXYh
8gkC+e8HLoubloMo0Rc1kbTJXmXPtYc+IueDnDNOkP3uowG0slVB11MNEuICcrSPLLngCHXKi+lZ
ra1FqhxxqsZwlkILYp+/bVGd0q7s57Xnm4WrpfpDDyGkB2+oaYNpETBOiL/xG3IruTa3+EALt7K6
gV0NSuSBC3IEqjZ+jbX29tFbINT9oPeQplwRLyV6YefluHzroAYRuW0N8CRBmMQsPRmD51dE3ORW
rrR2mKl6F9nrMfzwNfVeGDyMUwauTUO4SlrWz5RAd6khr0ZgxEnhPrernliaGseMtgvWCuDTa2+G
pI7EHDNKspT5BXbZe7VarZzBxznhrDZwEWt1lYm9mHpRw+TsbIaC/dXEtWbNwBbCT8uqdaX34KQa
YXsUNP1Zq9xE0WBbNEbyKl8F45F6bmVMvaoadyCPVFKNHZXjVGhrGwxl4sDRcimCs1mBFRpM0TIF
gJQwgbx02Ew5QHKVnKgYisQ/dud71NSWxWjNAOX4Sf1T7FfAINeDSUpKv4Mi4zMPCO1vue8At9v/
Kf4Kt0+gbJqF+VxqeFmh3alKb5gL3wr+lrUaK51OnPoOK74fyf+pSBMQQ8TX06/Sbxkk5h52L9T6
N2/KH+NgUNo4+VGkXtlZCKCRSYJPAyZakiMzJOyWo+OobYErU+K59UERYVBnw8sL+1xpXofT2HhH
ohS6y35+ViFjFUR91vcyRiG+xaPXi/2B67zh6WG+6qYnJQyl6STHWJC/6QB+OSjrF4XwgLp8XKtj
LUtps1l6DR3/cIwa8q8vMAAIaWG36+iRbp6a2P/obIMnYEaNag0ieZuiPwcu8JZ6t/8FFszZpb/d
I47sTjS8W4Y+WvuLZJbrlBIo0r00nIhij2I8vTSW85wXmv4GJpkWJPEW+H5rhqyo/hCfawnQXrpj
Suqkzb9FzhZmIwBV1aeSyfvsRmBL9r6iv7VGVb+B4c3hJ1xmYCDjfRcWXSff/Q5OWgEWoXLuXj/D
dfpyiG9sjczaPJU1WI9b22nKHQf9JPUN6g4moDMDTkcXk2ZCpHKrp6JriMpisdkkB1FGClPVWhrV
IQDxat+l8nx0eTpR2hM8pG3Y7hJz+5n0nwQvgatijw+8+yGCkl/y28dUEGlpbJRzjJh7PVlPFhW7
qaOfsdURo/PP5/k8hyzD3gcdWtESzeGWjWNFfSjcq/KoQe40LmNz4KbpixAXK9SoZaVFXc450hY2
J51QgZrgftX0jPVU2x9IUOu2ijvjEl+mDOwwGj4SlQOMUgjxNVD7YM97hClG/TjrvSZKp/+7B5VS
KOh6pMAlRJFCpTW4yv3M/BIK/5qlTIKutsB8vHHqzyS5FOlbhD6B8V245WuNVumZrxoBQCYqswWB
+Au2RtnUQ6pVqW2VAQTR79BG+5PV+LPvWwxsjcZeLk/ToD/vIHphfM7/dWtKNARprAtmMGKTN1Q+
ODkPUpdoFrdMQMqAUTZjTdpNGQBYkSQIayE4GN2JHGfEWyZJKUrQnWIheKjGDNxXS7/k/EEYbU++
nkXu27sgtfuOerJlVuLVpnV9sFgfqNfpw+xHs344u4Fz5uba15XSx9phB9EFrgV+sUBl8qrUZLis
FUHmFeHqncrZlu2QwAqAnyinc32i6YAvNcifyaomqPj8qwSSyA0PYjn3jtUChJ1SuFQ+yH8GBYuK
i0Rl6qpmmG8PjoIDgbweeJysH0rQCKarWh+u7Mhyj44hX3++h6TNnWtY41eH3wE6YgJbEl28Hpxf
oD6kkpVyxQZDyUlPnVV/04c3/Ouf1nlWQhCLRlWau1TNxQGXA878sKRazW3QSEjBedz9MjLbsjQu
1igTfF1SblU87gLBInQBSTqXfDEyRkckuK86Jww4DF73mY550DBt11gtFD8Et/n0NFhOvHnt1ghL
dBNKc28BRSPJfxW6yaD8wkSTKY5Ltfne8mG+t/vNX6jq9EwVG6+FqrOIsFQtE7rYDQdTxDKiBjc9
KiuSpjE1j0vPo/MjfmWKB31OM5+m8FfAUT6SLtRuFIgLqMTTDB2WfO1SyWV4k+U6czje8xCVevUt
xRqfZSTkds8njBCdhy/0qrhNjYimj6eO91mlnwC8h3PCJK/Ge7son7lre494w9m47B8SSJ2v8f+A
j2mem+GqJkRd6jIKSvKIyt7dxElhMk0HoYtYott1PN6Fj9c669gk+4RLqtlCtW2HBmQ0oK/HzNsB
6u0A30BumC/bVh8dEenjFHDQK5QKZJct9UE6F+EktGiVE7VAhFOm22xbuX3JDBIxfZMnqFcxiWHJ
6WrQeOvY+Nlw2Gb0IgU31o5spH3uZEw0qfXTu+NCL3N673mlvmjiOiWuOY6/JMvyj9cWwYcoJI5s
LX6vEFEqDFFgrIhJwDJqqm4s4ktOfmWdFjHrciqJNqeIM9Wg9Ed0mSDrGOB+eUPLnPWOcFlsnuAs
r8L6AkPxJ6x4vtMSWpG2Cq5r38WlvK0NbvVBtQbNP3UvW4hAoQqBPpnxo+cYtiWonW3o0lmvQiCR
AOXcz54qxbxVG8wkIJBIrtZbdN+kEnfhB/a4DrzoH0I0ojlCBl+/OwvasBvT7IbZgDEOBJfMeiwK
ZBNgJ7yf6+WcCVrd4kQVbILWVNSNdEFdQa2/hTyHBDdxxEKFoSbEwWuqfp86ILD5JorE3o8te0y/
0Hd1gzlgsypIbLI4uyWun+3n3TKxRhEeP0colwnRDE7rCDLRBq0LmTnnHRXX0hW3lIYOOJ2DiXOj
SKnqxNh5cXzw08V8wImGuisrUhwi9ztVctZYVfutpUoZCBYk6azAnYVhZpbw3qDOeI4I6EtLCgkE
ZgJED0iZuJXCXR2UF6FL7YXf2s3v6JzSKzVArexrvQErSfl3AMvyKHbGAxvKKIZUMx8hfUrEvAnA
ImYB7eXMC9QPqgGE9Xa59M2bQnu0AiDlpIQDw/jcDXFHQ11Qy22toCO4RIHfcWj7h8wv7I4twMZ8
LqCJruY9yKgDe55bIMTsa5wnfdqanetZRHFpRNDcP2CBBmganZdm9mAiLSlKwudtZ3e0aflGmnfm
k/3vFqqM/AeoBO6z2A4bY2k/UDJuCayKkA4jcaeT74P9tTu5Uy3cH9UBsRC2iKInrCLHbufKbeIc
wCfOfl+UNVL97FTxkUJV5omNz4SwHzBX0p0IHXyz5O35Am3Uu4YatTS8fNFDmkvALVty6hBZNJZ6
g4Tl7PCMyqnKMQYIUYJL48+tBR6bYgeVNspf13G1Cg6Cjokdlf/Y1j01ITBRAUzgh+kjVC6v0uTc
ERiEah9VyuCmSAhuRcviqYCYynRASiVdjtbhtCgE8+k359VbuAXHqw/SN++vySz/nH4vufbUufql
0OLRaLKPywhVXsXhY3bor/sRNcdGLmd8vAxpeK6sKh27l7Ov02gT9L3JeDUZjw4O3VgYOpqkQeVl
+rHmMspK+kqkWoyFhBTveqo819KK8Qp3MUL7iu8qcT2QEIHoSVZtJgAFrFoVIfVUN7Z/akCvC6qM
Kyfnh5ZrSCX22nHbhN/dImavQ5S4CigzzpHGhCE+1sF9zdHGcXNJ2Tw0c2So2ypEnNn8BH2EOjCa
0Mbm//WMx9ibKePkTfW+FQ46V6zsi73tjPOQ5Bk0Iyn/WEAo6Kl5z7bTAsXZw+0aH2w6F5jhE7c+
HEfb70Ji6pt5aQOTN8KxxuQia4m4OCYGbMJ21EN114y4uMPddm7/qY9hJodKnh1vzGkuRqlTq8+H
+Sihvna4+O9IyxWv7fQQXmGkXChZEsAb80kFd9iDXICBBV6N4Hps/xQmfYu0HFTJFD4247KjbL1a
Xwh7APX0VpKLHt0Vu6DfV8uxClhqrSbRFeG8wswBZejKh/k9H2G8qeRfkYqUT5ULrdyqE9kpNqSY
qjywuXQ/AY9oHVt8jyJaVz3XSv454nhwk7k5G5Y63U+NNXlIYTjO35HMbJNl8aFV+XjJ2U085Dnl
1qRh9ZfqHTx56MUyeNlX9cafGf/SDZtInkhsSiHMnSxKyCK/dhClxxdyTW5xpCIj38ppZ1BaDj5s
yLJK8z234Ms1ke2uUvOhDi2FOmcfOjBX/aV+Pwh/keUfjLV3p7SgMXWaEBCkF7WTsNCTnZOEQJIp
JxKELLDVf3sLrUcGMUVBXAPCchRqRv0LT4tvQNivORK6QD7QUEaNGE5f8eUssy3tizEZIpo1bLXa
aYgJNShmVd7hSm70cI9Q+HIS/uNm0rtS2lRKkrnm4GboaeOdlCs8L7Z4SIgweDJqggFGvwmSBO7L
iD8Tn4MVrxir4vxDASzK4+Y0c6GX5zLEtp9aMDfvnIqeI2ISo7Q4vJH2iotLxiI0x3MP3PD5dH2K
NrgIZU74lGN7Kzi14SgWzAc9a0DcWC1NkGjEOV7Dc6DXEbJvgYdvOXFQ059ydzlj6sPI98bFz38z
poQXd8MP7zvUme/ST22Tl6b7aFc09UY/zsICrD+mGtKU5iGxXw2Prltqj+an+zBbMZJrtNfRoUsr
ZeSa+oXCO+DyXACD9pzAfJYHcrhQDxjLnHgWZKAtVIyuG1vVjqndOi0xlkamJwqPbl7ABv80fZ0L
/5m/Zwz0aG0nr6tZCve5b+jArZOaCynYR2+kJb0vqhJD0Rg0zpJJOCurpTwv4e6bGaPICijKFnUU
PlpJ0wnBm48eaBSBwSiQLNnK8YzIK5/E2cvYdlSga/IZN+DsBQW78mbppAVROb73GAtg2099eep+
rtbhVWLawJH5qRhv4pijSEUhE3FxfPnyPQUME8dDNZzdQnDwmC5mFkCcVvjfObS2ToqVqQtmW6vw
AbVlin6WyEHLlcDNCX/siyf8qCyQ4ohIgAi+gjyWqhg9sYhTKjucZqtE2A9YUAZN0oEkrphT4MvP
WqBzV6elYro8KZsZ84XuWs8Z+gLNNWQn6SUKzvnBX39xqMXneCmDLQqTPhlDOWeLTsz07B2bqH6H
82B5lBbDJZkQHxoch0bkSLCLuPqfxpbMub+01Hcvsnno6BWRbSUWhhtTCSNLQHp2halbjGFdARxG
9ALwGrUpXDL41hdvM1TDwAqqAHGsDfdT0Kmaz3KX0g3Y59yNiMNc9xPBhkgCKV97G7d8ecdYlC3y
/rj7mWl/UfpG98GJ3m7gL2mw+2F7k5k+Zd95vxSXokYyqk9SQfA9yZZVzGNyslND2JxmOyttpJTD
BzbDKZHrtz8VHUKlQw1dfJFC+F6cz+1Zo8hHOAcLKl8a1pEpukiCQynHrrImmUXYps6LhJ3JiYBc
DPmz4CxxQ/aWmjDoKZE+ix8C6Sj3sIlCtKvGl9VCkgq4HeYQdtb/TU54jpUk05vqvmxxGopf904k
AWzO5IFlEn3YuP1awywahrFUSNIB2usMGRUZ48OL24zTjzff6WDvkax6cf6IfotAaYiBmsnlTBt6
izc8kRQtXBPiZiqciUgaUHsHC9AoaOueteghPNB6C6Xuzhm5N3HDj81Jmy4s8CLvWapUoENRhnHc
wZv8zfBI/U+/uohFVqVOzQt9Wjc0HP5dWgGGZyUai/Xi8m89h0yjoAxx8ndnUv/Crt/jEK8i48WV
pjdBVL7nmyfgdrBftnNfTm5L8NeT7l0Y5VCdrVyrfeVAHvxi0AyIaM/SsvEWdZGBE73SMe+O/RHV
U8sabugQPkTT0gpuG4mg8yRvsTrvIj0nG2iOUiofPRuWYBZxFmhKKwmrJ2pIUoNjwUMUBVThKItr
LH3q2IuJib7lCnXxGbEkHsjhXaDwAR+H9vzwdPEtih6a+aRSR2yuS+YlLSsUB5BWhlQQzAcuWF43
0YYxqHo5nhohGSNB0BiqJ/KUa7nzRAaMQVxzhCJ2U9dYXPgOrspBQK1ZOARtXyfQfbSan0tfTFiM
78YQ4kf993aJ2lReftOUBoEvfZogCt9IXsdsdjAjlIeG2HMD2KtCWltsfTBwbZTT1vwwGXwPnFtd
L1yeNKIPVZ/9phqrav8JT9GN2Jyp2wFb9wG9iZNR/+2/9UUP8Iwye7IkF/ePvA077QOG0UQwSzeB
i9nFY0ifspmDRGanzHMP/MqszWlTRClD4S5hJL7NZ6KYJo9LRkylhhrJk+usVrV8bOuQkOE+3Tts
9eLjg1OsZdD0GdihQMVb/Ik/mc8tjg760p92i697DUbP7zdBWnfkRo6LqORJh0SpLpJbvAtouzxB
w5//IMZ0NTbAnCOQy6afZNc9SUys7eRtjUMzekmVkVRz6MKW8PesHh+5885WEMk8rmPsznZQPujc
5wBkYZtAQQuWm8gof+iQAWAfcJ74NyCHfa9HrHV8SHC5WXO1W43FHndOpoAUOntPl9QIwgMS63Jj
iQykp8UP75NS3BqFzOQYSrIJQRUjh9bZEBh3Aaw8h//eKSoq9uUJUsq3HM9GcUn3ukPLsZTmZgDh
n/C4mSv0TPrOXnfoVWBQcBxqIky/0vdsgWl2j1OcQejoi2CbE9G1s9EQVCFoPNHO9JLOQwl14eGJ
s/yeRHsi5QEJqmqv0u/iBSmHmqHzLjfVB1i/JOEWzQ4IuuqVFo4CUTovqhyMS2uJauffM3xkvpHt
FyJbCyPmFzuNwkxVnXyTQUIx0B3fSiNfO0ZZu+zzTHdQXOU5kICZs6U3uaZOE0VPEhJtdB4EZpUz
RQgFjhWO9opiEtD7PjD0VEXcAI6EMvpcPYrDIjkC6gbOtpHvBf4CJ2VOGlNf4hf1iwv4yJbfRk/s
94gaRLvnIa8RGQH+d92UAlTGj+2xtcMaSnTZWcJN6T865uE9gUhlGSnwGBwaPH0GZokF7/rcY+h2
7zhIx7wLLkS+rcO5yOUz+HN9bsoI0V6K+JrszV0JGcevw+O19PaQoBww3WCRyy8OgEXPzCjE6HwM
tnztzTi3ZrP7sXaPx+aqN4VdOxnLFMyNANvX/bDkGGFf5oPxf/v/zoUu47xUvzK19DKzIrlUe08a
2Wuc0QDTd1hh9/w+xiSuPY7TgmzE19rlyijpnaR7bTa9uK+1DY3RAhzcGfL3mi0zwD/X3XQhzfd9
rRbZhHZrOwuVEGGdFSK9S4pK2/yrIPoSMR3vSuz4a8ILZoRG7gJUS9/Yfn6xDR97SCGwpTgwDpRs
0PPpfs4Z05xOFADEbR6h+WLHiMXsAG/QlCjq5yLYuIOxwJyyLpYGZwjhpRgm5ZM3VO4oNmE12GrN
hF3Nji/+N2aPlstQ+P+yDiACn6szCUSuanQIq1Nf9rowZQ1s2IzCGnylJn7M8XZ4KOf8GAjzBpKE
oHIEk2a9nlGm8U7I9wUdi2Tazg4PK/WQ8nGJ3jE985vmZVp0uYjlqH2EKh4V30CA309v+asxkEuy
oFoYBgfwu0CzktQ0NoxOhmRaXoukdaSLnN6eiQmIMa69mb+gXxHHDkACB/O9D/yiMb6pc4uMnAQE
rPQ+iw7lP4SAFtSbsfUL0sllWNhTxWOoYzS4Es66ski2EZ9YG0t7L0F++xqLhO6gLKHCKpwn4j88
GYm+AZvVUOyWY1bqcGlw2XHRlpmVPBhie4eJi5G2MkLUVdpFOA11EyY/THiL3xYtApmyyUrTiwi0
JKO+1vTE5b5wn0rBUE6QdmA3H+FXPGLNd+xsIaVTD0BsIOHssCopX6F1PMnrKWv/DBU8F2umWH5a
9lTgD/hXH404Yx3l1yB9YA2qH6Z+xL2ZEXggncA6dAZnadbVBeo4FokAqoWrlMLNSwD8/pFYDKB8
AmqBUxKwDkAdSe7IkUUdHnJS8BZuxVtEI87kFfMKDjZR62pcEE4+E1avO242AOapNgj28cmT/rYN
b6m1ED4ORkKu7RRwGsbLXWOXYudfxpvpFbMciKHmXnUGHNg7oZWGdSAE+D4hH8c6aGBrd7cibiUo
rNOKsCSACusUEITuRjIbIpzn4UEN7li5c0fxOV5lMPUve+mQS04NoMtVVZgPMvVaWxuftHDoMSzg
AzPx670LudnIaHWb8Ny1pryPYSIfn/0zEwYz5KUVvwAnb6oxRd+qVBXuBAIc8LwQyRydPRs631vi
89RUUejv/JAp72UK8vQQYdwC95ZQXtDoQi/hb1bhZAThAOoUVGbtZ+mra1nHWgfMGXaNCPFVY2iV
ZZyGcxH8aJBR9bEqnIaZ5vaeyI2Ei1rwSl22clnOt7TzNrU1GDS+G98DiJUk44x3i+mPq/tVEz+z
4sKzZItguFNiHuZFVbhG6wtoFaTgFDyNBSh6XSm43OlZ8ThFhc+0sA0W4RSvsIeCZ2TtYFeMclbv
zAENtvwez0qeea6TrHjjCqQlcj+j5Csdiy1i9opY4LVrec7Hn5cnJF1YtvnFdQeZwDHyHhg8wNjI
3evu+Qcu2DOtOLl4f5TEfpTivrbSqn4e+IcPtpw4NNQXJmszFLJDFH3nUVLTT/TwfUrgc7VmdKdM
oipiv5VarDjhJcEId2/y4lc1xYMWRyGO72xEfAFPRTFbFtGX+oakHLwOeR3nkeYNswDPCTDFWft5
kYoOgpHO53uAHY9ug5apdmtQ9tAWsBWzodHwDXpYb9r4kOXpIiKvxEf+q4DnVrpNH9YwQlNz5m9L
7rzRK3MuO60l5Eu0x9FowWR18ArYkDF7xFCrqbIQx90Ug6REGrvMRKG/QHpGOipKrg++YhMPTyM5
nLWVU3N6XWx628VwTuoZEfh/uPQK65Nd8Au+oW1Iq2OYDgzbc2lPFN9Dy/yqc/+PYsgSgOftTxlf
pU36rHZG5dcDgmnFwGZma11hB/cr3zjTmrwj6WDv5D/BepVLU2xRitfuysoq6Tm5DiqwWDhL8ulo
WY8V46qkgXf1xiNKarI6EHTDDUPR5HcYMzKep4jaNk0vcuD7RLQfkPfRTK8rcKzBLlCZN+8U1JqR
eaaf60Yc/feqNHTfd/rL/qv3EIDRTpgTWuPl19SHpA8WusoP5TcCo44zQhUSN9qhrSYiLnbovDHT
Pm3PiJgIF4cXuis3ViaUPOKr2JQp6lRI/z8Nr/gDnTRnzbqxiydRyfhlvG2aBJEiJhc59Wr8srRU
5gqEyfbjE3iIlbJBeejNEX8uy0aPKdFt3uVmJlRSwoN22VNwcfHLBBFQt9CadHsf9MU2d4eZoB18
mYdLntkDkwYqBkW+SDRW9Htu7y/jxTlpcYC0Bj47+AYebmQZ2YyopFNi9kPxKIlmbjXtnPchsAER
rC8d4hhUcWS4ukglkN25h1lpbcCCvbv2lPMrAnTUF+UXjJKF/PLKzXDu0xrg0Du+IiOf1RMpFglI
7US7jhUwkyZt7FWBStXxVTpQ9DWUFbpttDRtWJbycbjANKOtSjTBaO0QPT0gN0lLvw1vv5rCgsHM
CxGnHg6pOrYQYKquybjad4PgV9rL3yudVeK6213/VtmKF5Xm6IPJD/ohICcrPmze+9LzFbjhCbol
r7KRdxJMj2mKzpNsJW4hxueHcDeNy/YbcptsZFu+7XY1phFBzq7quz/AVFFo/eYN5z52Kx8YuubE
7BetQ7TIyk5LG0UHenwm0z0e12+D6fJzGp8vNTPuQ86d4SPpvJNv2HX3gfREPXwXj2zxhchHYZdi
kNIsxtgW2HBce0VYDN+5/HUNY7OLi9NIx5zwp8ojU3to41x7fu39LBhu1TVz4Oo1spXPzTTIPOWT
u1+SFKK50OXIFR5BfmVtrAMvsBdqRNzV8McXEMUOAYdPb5EomOU26GXv+51y879Wr4ctdvlXmiV7
JUY0NO0OzYXsGz3GswVXN0K5MHNlUfWzWg5MSCf9Ka0wm3m9odhE4XOf0CiMdwI9yQGWODenVEIq
Toju2m9PV0DYg2y7xUQB1WV8UrsUbIBorFJzYrDU1VN51tQmc6C1BHO3oP8Pn7IZ19n1+VfCZrn1
kUvf0SM3LYzaUWLx6jZ5O3hS54BZ9StOy9N8L+wO8HiVTcNGafVmt9QUPpE0Bco871DmpZLqJbju
McNeXAai62W7kgGU6hEsvMRCgkzFj1CYoGa500rqcZP2cqcjpUQeN6byXCR4k/ZAUBE28wEGRc4q
CXxtUaBeSuFc+qhPbBi5gt+U0fY1HLzbvg7aSS8ivMsCkjZnLLckdA5D9EOX+NmiuME88LemsIIK
OfHdWO6e3dvGBro15Wzrt2/Q9B4dXigeEJAUQok5c2+xhcDhH8Kryx1xhlv1ZLILlguRa/zNAf5r
/COk2jkHJc5r1UjU3rlCulC6sv/T4WDjk7LNSmavMWPcCubCbwY1scfS2JGFdrgIXk+F7vMdPZ2Z
rXdpv8sEiFpTvS0qMwL1xLpXpT21rX5lkisFnS8xifwrXxf8LPE5xeY28bl6C//IPzO1HxMnRtGD
g3Rymr5bLjumD0uaPs+r0LOg0SWRGSGsUmj5hDU/P0nn50xFnPpue0U4+BuBg6ihCuiMdW70eHQT
WNgRrmeOzudRkphXlo/W7dyZuZQcmLESHuiEUnt1q8edaqFIl7qHq0Tk/IjVoJwEoKFpRTXno0vQ
RGYr5M8I6Z4Qlt9EjeOs4y+/PEPUqddk9Qi+iDC3Gr7fQ7Vv1eSrLFhTq6T2l7cDujZdEjC8yFxG
zhTSH3kbeZvn7ks1sq8TejzKnCDELsVUOsQx4czOEcqQDb3J3R6DEAvS1jkka7Di5YzyA6NDGO9Z
GrsslW8XTVCbPILl3Wba76RxEcSGWPblTwHknuW99kZuw+G2ugWcqk6eJWdifC6JI2WRMg4OJ8ex
epM4Z7rvWnkGzj8Rjrc6J2vIDXNfJRIeOk4SCZnQTFvu0t22f9Oz1oa9ZDV0HSeEqc4ygKdV/hGE
GTnjtTfi2NPmpz+gHdo42lu6B6uxRG9tM84A4v9r7a8l9q2/Hi9jIxyPDze8C4Xj6e3RThthfCUr
Km7tqtJ4+5yxsue5W4Wcazf/s+hhfbSQ/hJZWNV2c+0od+AYntcll59wlSPaXHce3+IBRQTySiOe
L82B79T2vjFho/3j4ljQsXCKm0KeBRO0SnjsMh5j6ytkqt2hhaj4OWsuK8rjD4ogaUBUSWGo9J4N
OMPOEHWDdA0XM82zdwpmSUGGrGgyAOImq+0vmS57nCnpThVyXyZ8guKkYZSliR0q5VnIfpTcbPKF
1/dYbjUQVgu8U/OAm4oMZc1+vdDVO8emzADmt1+o8EfKwJBSM9MbK4zK1kZeJ4vZWRG5EJYGHrzz
KyxvM6XItA1h0wvNgDW46zSRanWGyvvZaLFT2VzJv/1ggODQ5fkc1zRfQ7skox7O+JjtMmzEn+xL
NFIfsY51sPlw/hoRKF0oz4g+cW/LXaA7yAgkbYUJJML2Kj0AWk+oz0cYctqzM2r6evJGgV8OCRfr
1GeOOhy7jjVdzJec4wr83s0kqvLmvXbC/8vMnQT5s2g6TjzVivKlG8N2SyHmMBb+kl7Pq4iyhFr5
ecxJA4RqxNBrpLkXqGKcUQ5estaECi7KzmnOQlySHzZ0SF8Z7hCJTO9ULn4iaitdqo8np8pWnGAY
Tj8Ymx0escLrJwCUQmAvjxS2jC0xAUslN83kJV1VezwjpS4YduGmh8xwPJjGRkrdwu+E2A2PG1Tn
djvOLFbl1Gf9Og0DWVRZTs/XnMaEsQMPLVfIhu38IxChHT+noiVaY03micZFEQ5zlQ0l38oM0Bbj
1buQ5kXJnUgFSpkX8PkrQe3KmjJrhVZwYN2RuG+lX2cihwHwVz2MUnsnCjcG2ss3s+YPfpJWpeWX
zoL5m+Xyykat2GzcTLlzCMHUjyvQIKEbg4v4ut/4xULRpUK7XVdyfaLu4JlrjX8Ky2BiP223n5h1
273eOMKew5w143383mNZtRxKsDdryC7AYbEGT2GQlCDwlecHgB+LvKPW74hEiBPFmbNaQuMMnCSu
Q8OXuI/jy8IPFfDu3lozAhGTzM97hrzGx8FvYmxIhReIlOa7BEiM0EeXf+Q3iIDg1lL7uY6tEZZ4
5T0yUcpeXhhpfUug9FyShzyH1Re9bbFaQnSL8zj5shcDizl3Oz6qL/ebmrGp1EHaBmjZqg7+7EuJ
9aMHwM7a7s5jZNfHVbiKSsP2YXVOBMlwcjv0tj54hd5IIWreZg2Dq1Hj7djeqRsv7GwGeNdDtZ/8
8c/vOOxd1M7fdOLV4R5NJRvZjBHE/R69tl+KCfYTmMtw0GSOfg11qz5fXoF2VayZUqda9VjSuEc+
MU4J4tL1gP2Cv3neVvNvepIfbBYBjt8iGLKin5LZrdR3wJml2gquTXxd06IqJz+hFUG3Zg5qA7PC
9rlVKT4fO9u1CpyYb60cob5m56FDRkkzVN+yL9dYkvJplh8DUQY3bdflDvN6aKlZI+EwyEZQ9AvG
PBfDKfGaHxAyvZ5wak4TpDBGLNMxS9iCEb7ue95wwISGLkGQ95TeGvb7VBLyH3uCDTJnyuW0/HbG
tlqfD7oGUSE489cUAWpp1bVZupNJJ62r6soYcBFSXxGSfD29MHaSjfZ556I9QzvaD2QYJ+8I5p+Y
4FDtqDydfJ39N85xrKpYbevMTWcDC7XAl5kAOimXmjCRvt521q59fh6wXXso5l6WIi8gAPikdQST
PQ2kzj/2K6ldrNImF+J/HyiBOqayqmsl23uE4A9yonfz3ZHCoHYVTrpnC27XjxQnuRdhLOhuqE9l
aOBGzfZDFZH7K/uHo7Ffc5gBEMj5QOFWfkGDa7SuxYfqt9bBFQeAUX1WQT6zx/OfQj5pJQLc9efI
qk/RvcwWYpuIPot05kMfNiqjU9yRDG13vxwERxbeycLMPiZ2RNMJK4tBCHaA7FkGGDIdNls8MsJn
zHgeBF9IMhfh3H6H5pAERrPrSVDsZMwzTiV30Ped41cJwSAycZ3x2y1DQELaVz5kZWlWYhVldEfS
WCDim7AjqJG6f5nN9fCbDcRJSSqLyWi6ergt3v15ER0+XskcT176CL00f5trlFGWOYZkK0X8XOZ4
dQI4CwmfsOxc2r5jwGzO/97tMJNGjwiIXOVp5vNEuH00h+2LUmhwPzZf8EHpfFvb2LGo82aYyQpX
7GLgr7mxaaJ4r3QkBnEWsrqkvpftIA85YgHhAALxDXPaz16Q/FNuCZMYxLY1wuWfpNfNocKQO3cF
DIH9SOmsvKuovQRP2uTCodLFJc4Oq7lNPBb/scJ4EtT+qSNMWRvagiQ9OV7IEa+coAg0/oX/cuuj
j2u2oipCEklTeMBCDV+U+NHHs30kXqER7Z26KbBH4gw4hu9AekrsJhT5GnfwNvBEowRq+5LTHiXb
EvM5WNn7VuTyYcy+wQEuRMuUv+xLZdFf3oKGvINgYJD6DKOfflBbnOj4Vd1nvIrc3WlqZq9uZoX8
n9F5wkzWZa82vvD04SNbHY6sXh32jbku0R4y286Lq+XjVnILYj1NwkyqerDu+7wc5aExTPYfFaOz
H5y7Uzm5wbvQD/U2Xo5R7dtZ4I7OCaGGZ7bM0BEy0F6WYTKCYJw/RvAsPLeHBclHtMbZ0NgYvybI
JYTxbUF9Wzjis9OG1PTeBK4P8cSSjjL66owasx0a2ivadZKC4inQOkmkouSucOw5lZDlFSrkqOkr
lR2nAxKMd2vCuHwKstWekHlm+kadJ/VCpCcrkdBRTFjUOg65UTdOcEcmLnu6ETTREFkkrHtzflhd
Ckekh2/t8oZA5+2gjvYDnLuicbKvqSWpvt+UkJxZlAvshoXqVNxcB0qc5l4u/htDNCr7Ix73rYyt
mj/ASEcN+Hx3kc8sbk0wwGYyNEOkXbgVDXWqVvtLGKKz3ysI6OH0bLr84gFuPrwph3SHnulJ9PN+
pTE4sEm1cptaZjivfDFxlyyO4S8o00QMKVh00Mk8Uwe+WVlgXqgx3pU6xljnvnbaQjzrxPGtpnIr
Wi2F6EB4sEUIlsdrMiv+COsSI938rMotClL+/35YxdKLtrgxLqp1SPGI97lI3zzwsTvv5CutN6e7
6eablNWYCIBX5R3X4OIB4IuAVOgEH8VmqMSIX65XQO5Qa5fO6FlspMIn/AZz4Jzg911ZwlbJ5xst
veeB1ccOsTV/mq4KsZXfYMoWA6AujLhOaF01hIp0O03y0RyNdyzVrvCb+LAQtGUbqiurjJWXkiPt
xpyHIpG1YZL3PJ5kI34Zy/8EAxbX0Lfh1cp/Qj9NvmmtsskWbhumjnK2cKNAG2+otRxxbmUWa1Tm
kXF1j+l/fNvAohii6zdvX2OnaUJ3FUNBAJ0aF5cQCNEpOOpW6A9b1hiCjFAbLVglGwD+3ezhR3c7
5NFrsGkcNpNqcW+N1hYfu9yjmIK83UCkcTNasHuFcvVJqxiocfDFm6MbZpaTRrUbwxdsZE8o+ezY
gQo8zNnlNK0IdqpBxJmQ+tddzaxwyt0tLekXPMn4s8Nyw6qoPZ6wDth0W34DbrpklNlFINltc5W9
bo1X14E1xxEdVpsPqayzKb64x+XRY73POFbPlmRoHM+iQ6YwQRrP0XsIRKRNpngHWR6WtI8xafZg
83sUIi1WjBI9Ia/0bUq4Rcbqrhp7b+DckaAcgnWafk6x8dq8x0mPyjrKaif3Mm8yzdMxIoyHFyqx
2Wp2PullTyVs9EZyp6DZoVDlPAaqjBQppvAn3UKeb0StrAMxAevmXBPtjiN+tLs1bIbh/KlO1oCI
0ElGl4EUuso79juYSx9njjTGA+bxjSFKgvBxaCDAMTC28TP/KJZoIfFsqk0dK9/4SsHVMeGoIpg2
Sipczi3O/4RhzGBn9+wX4FZfiRRede6P/RTMQkaCi0O6jBzOP5O6pWzFgyVMUVkcxwZrw79xYeSw
cJoQlI7VU2YMYfwSdGNc6M9G0u8/M5SQyd4WIZA2hzGnepeizTHKErUdQNc4UBtHRVj9pxBZ/Vi2
7e2I/PfyLFHh35XGLCCyaQmJimZjMVo8ZYZ2QqUn2qSReSoyd056iSe80cDy3Tv/2liP2cNtv5PK
kwwRGZw6wXgjZ8KdQ1Zg/Kg7S7eem5i7/lvVMkJ+5JWw3aMAAJ2L/vOksxc2LWqV+VQw0fHDMP9y
FVJXzaTuUSmLKo4x5WH3VJzUE08vs1xXCSKGOWIMmTE+8tvdsLEOjLOdQrdA4XQoG08ZaDIMBTHf
Q6INF8hLIBz0AZv5ilT+SvtBGm9D+Bd5r5n1WEDSRDvFEwmA3fK2zSGOO74gDS5RYygOawGf2ZDB
PhLu4dExnrHpRs3LqOl748qdxf8gt1KAXmdXsnMkbvbMNb73cb7+fHAD5UxzI9ZgVin9wEuiOVls
qAOLSqhbNg+kYFmewB+Pff9inlTLjEMoDOpiKGqThs1+aeQ9wrxZQockrq9oPaZRubyhXH+Urmrz
yJbkvGIuH7kHWc1AqO0Mh9AfhKQm4V3rDnPSMJihtKftF4uunbsaWml9xC+xq82hkK1kvowHad2q
pcEF7MmSrN2Il059A/QOVZUkKUHQimu487/X+P+QP7ksP028ruJk7mF03v7NX96k2Tk8Hdr57S6B
Tc+0J9eVTJtbg5G4/4gj3OYG3owf1dBY8MD0YK/etyDr2I7vUoysvw6i6IEVrc54BQwzScj0shbc
p8nTxIArRDTcUmd9SLek6alv95Cerg6m33CsuAS6XM1U76xeEE2OFT3LT6QFN/on10ONIDd/YRu4
uWcin5w6WoMaJlYtnhfVOtfizmJytsj5eshQzhLe7NOtIR1PraZY9NMZtKMXiR+kZVEnSYpjaw6m
Znq5xyqOG/ZmxEKfSa+++wgHItX0983PXxUXkwV260yQWZpRp0i/ZnN3rHQjJWzr8GPwhes0Zzjd
XcM5Zr9gwJcWDFl74PONjvdDP9BqDpMLGNAkjzlDXkqQbbpqQdaJ4MYdtOXMt3Otj91UvxetQLUG
B9ZI6+v3IV9fSbvNqKqOyCFRYOjR7zdFNR9qheyQz09+rvSm2PlGLF6+wa0PGI5Q0xUNpX74SRhx
2izlm9C4xDrgqCMaEv+zM0TJVHQUlVMik/VjmRg1JfWERzaEkuik+30LchlJ64mCRiEEHafTYZ70
VkTBKJOF705anIHx25lA63J0YKVKj27tgzXNAyVDHh9ZVgL3hdRUieDEaQeLe2dQjbj0++2/qufS
R3tLd8+xUEZOjIpCjhi/KFEhV5cv/5etpWaGUnbsBZIHmPptZjUfK0mEBSjXO+DW2pJbijGXBfm5
OAf0RIGX9Zmsmjbk97K9kbO55ZexUBf2vp7LVZVkjiKfhrWkcmJDTg0UaDfYBBMo8TDH7nxKd8kr
QzfgavsRf+fiC5bXPpgrBpUkIV7yiZE58xafiaJPFJbrMtXNnra2oW6wtl2wCWihT5+roumHEJ7v
MWAm29aL1e3MEYhsHE2Mew8vzijb6PIAk3WQJ1z1V+lnWZpwofqaHa+3FH0b8tA73oAYrHavk87L
xat6JTulZ3xbpF76kfIuAcs+S6wRoVkXd3fESfGywQlCXMdISLMIlSyKy9JlZA+7nixZpMHT8zaU
QunZAtucNu6AuOK0WCBrVVZU6CTYveTlRx/72GwVHDXjFLb2MePipSTJtQNHOoFsLu3oEO/yKg9m
jSNnb291TN9xyrttsxWeOymLbRHZ0KSXQq8iQ7lHc5ZTZ4LnWQFtNLB0UUC23EtofVFtrYLWQM+s
EAWCuq7by9/Ws5xvz9fNb2rq19QwqIqPgdzESNHFQ6NzS7xFtkSIc48YEXlRPwwE//MmaA1TiOU3
YkG9c6XBKt6hNufC15nk0XuFi6kQ9QXssnrcfgLi7PilglrzbhzwYc4pnauhzwiBN68/E1bXvsFe
loVfXyhNUNzOrH8kuTx/wgQvhTRm2uUQCwCB02rHmPbKSTIe52wA9QUmgBpa6LwGpjTH1sf+h4x+
z/GmuNTTjK6m9QjSPPBdl/0l7Boo9BVif0kHM06/RhnW1tYMbhm2hTk0xVeNDEQuwXiOne/w2moz
ruWLB15jKHoBHK3MGp+fNJxZUkiiWUQo/YFYjXWp7YhGofLBx8XJFQQuMzW27JCgkIU/YfvWfoZr
ADEqTI7CdZi8gOETcf3W2qTDxezOAkEnxCU2gA/OMvD25jk4eU5igsfkVoToZWstr2NcrUrkSsFP
oXMxn/eMWRoVnR1pbA6J9UpbH365Pa1cE+ufVSjSGn1anmY9FiCwWSCVdVmrZAdBuWvXSYPad7a5
LOhoL6GgMPYSN/vMafD/MUibDUH/yC/MzuzHSw94mRaOKnIcxy4Kcd5JcY0xa1Oe8nxBeg7CrGCf
O3fwWdhjmc1pg1ewP4G/f6/jnG1G+DYvJFjONh03qLSbETgaPX+VbbrhqlZD3yj4M7V8lCiSwlp7
TYoGoV30I67vrTrOgmAy8p5xWzjrWfmwwqCw7gggjzFflCtFalg+AS4roeuQlV4abNmyO2kRr21L
l/oGJpPfeWjlvmZH8+rEG7EWk5ONMavKWXeyjXXZu7ubaJDgwjk7Ev3q6OY5rpLKzM/bma8UUByu
ZGx9LsDioK0cTD7V+fTNSM+bB7n9VjFKQ9Lg/eh1Q3l2BBNhLEwGZD4b8YIsGLh3SfRx/2BRz3Ds
F0iEOJX8H45yg9iCWHKGUhO1QSqr+T9PFfA0MSD1iGlCQPEnYkAl+uRC4PXtjZH++RBjNaRrevRL
9uRhKF57LEiWTR8DtpR+B/mgABEyRY7PzNc8P4P4wZA5Q9DPFmwnnp//GWz1+GnlCPiBV8javm8B
XnUz518cfH69MwkzyXjmE0TRYF3s18SLx4mjcavclJCGnB1sHlzv07ZVbdA8AXRQZwCLHb+elBHm
EIrkz48DTnuk1eeybebR7Gu15fOYpjDLEoOqjhCskkJg2NKDDYefj+ibmzup8gV6T4+JmnQ+StpD
iGT+qV4TWQOjoWIgx/AiZD82Aox1BlqfjumKAxJ+4BvnzbGw7i0JQOlLMGKDmdRIORaM3VzqkWW5
q1vF5CmzCX5QambgYRozMyxbykbNw8e5u8cVvybgjeBkj1ihqegUdmUBLwV/g+cl7gZhhwAIrxze
GLV4Dookw9n6b2EzY/JmDhByEA4ESQET/cbB3cuMhg/+PRmeWGOw0gElS5kd8Qkcnbh1jT+QmmEx
w9ghueIKb7hF3eq0+CvKDTVew9KKoc/6ZcQYDruq/OY+I3spMak5RRTuDrN8zAXAbBpNm9Ei0x6S
bUfn8TKw+i6hRgH1dJCzXNgnJx4vzghdqajz0fP94h1RP2Uj1HPyeUfc55SnNlWFR8/PirZN9EDw
ZVQjGeO1VT3FQhQ4kQ03aeomPxHSm2H7MTxGFlAmQk7ARzkYYNFd4yoOx1l+uRaluvW55yCbz8M2
V7yq3HT3+kDB1fSuxBICZw3cfHIDLxlZmK8j1H4cyjXghmGzJrUyb7fHqzKphoTBKxqM6IkWzKtq
km9cpjZb75MXnfP3iXui4z53EsBev8MpaOgRqljampgCnureZxaQowXN1Hg+hk3V5tZDLof1PO7A
5TasCHGZjtpvdQD/E0pNY9zWg9QMFfJG7Z6UmQ8WCzqo4CNEtzPmtaspmxDkeZfl+J5YTfj3CfND
JNvtKNI7G0Bl4860KFeHeFKhtk/E6ATbTZcFCYaI9o5EwC07OoCbDQpFwFnaX1yBkuzJNPjxwtdC
g33CYZZmxN040inm0QuF2ScmVGcrtP3TAjJMqyBGu11UG4OP38w1ltVmOoTsQfrRVW3Pao3xCsil
qF/cX5wl/8V9A6NnPU8Kw45+XRh5BkGbytw5B3xP5Y5PSg2loJJ6Go10L5GUcYvApeI8JNUZV4Lz
iN99/sFL39h/DX2+bfgsA+MdA6RuY+QFYriPjT1+ICF87PqPBoBHXsTzgMrx/fOyHKf3E68qBy/J
830ZSsx0XOHutjWmqVRhjBPYdSvWOvG584nHrLWndziNeyPcfd6vDkxyPraGR8lnPij6iyHdeM08
IkSVj1HWdcQYab/Ni3hlT14V0iBYT6+27gQXPkYzl9Hfut4KAJzLRIAcS3OCcDLtAqXz2isnvtLz
2WRJYiWu9umTPEeD8+eziXDRgaQXHmBoGjcEyFpY+u3y8vnlzJhJ16pm29cB66sG6M4hceIp+GEb
5tB7TNe2a+bPp7rnZQaG/Hw9KyoRQUpkv6VWGLNmlCrU/LAPgM6sPg/oYdmbTsy9GvJTxbcqhMiq
ke7EnfRWgFmI+6mrd4SS/lG6r5QJxK9kztxOnMbAIj5K1iIZsX0L0GPju9RVaPwHRhcQFMfuARIf
h5d6Ef7tKVGW4GVrqbsi/nWe/BrJd43VTD9wB+00UFYD/G4FNkGUIROMe3ioJLsaSw78d+vbtoh+
Mfd9LyvEvtkEq61+6HWSrN5xz3zKvfQurvlYDzTfseVk/0SQpKp5aaeap4x804b9W8mq/KDg/V6v
MVW331bMfFE7cx5JgB20sebY54vCJmbU9XvI1JcCCdrBjS54/k3aA76MVgIN8YN52WVkjPZxcstT
ulwVMYI6nNElk2ztS/JFt6uO1qZtvXDLLF7OzujKBKQ0xMvON5yO1upLr3wu3QY2PsmlBoDPQepM
pD1YrDqIB5N0+qLfuVAab+AwdzQsaRjAIJTPCfMxFfIaf+tcycZu7ApQM+mjhmnbHAsk7YECFeE0
EO87WIlkw/viEPjNX/ICNKGf40rB6xePe2WeYDNHaybUnTCRYSffvo8zWJ9AvNdtYRedu+sBUXdx
NCUTP7tLHINhiQS6Fhjl62iYVcSK0qLcz2BURDYGGDnOu8OYfQaMg/0UxrWyTNMm/AKu9+xasojq
E1E3/QU0xfocrsCDjXIdWeutx3MqKvM8AwCQHfXJXtcVXDwZZ/E22KaO2KdDM3Dp/RXrFNIhPalo
H1zcXB85jGlK8DjxXk80L6pYP3SDQx4j7XRyrvfnhI7t6FcN1s6kNk7hQBJs8wf2H6aLGjNzDRbT
PSE/mNsLBwpQhSjxp9lELLpGoPAlaGzLYWSMyHrwRWstdgf3pi9PaRnINT9qqytR3qS8t/fpnB5A
RH/yIrexBV88FfGM+X/xx4zVdxJuaT9jY82FTXW78Y94zG+UrWe1nrwci1FkMOseHhQWTgNx0C/G
XurOHi+S0FP48vMso0MK+mcYlcobC2RhSnLk1qZhgZnmvwBeMbnYL32Lo79SSf2a0Y+4KKHZv9OI
c742VVc1atgpnfjRFgjAbnQNIJwu8FbC5ZnyRIN8sYlgKA+8aDlhWkcdHTCtq2XqFwtFp/Dju9cL
eHThhCodloFCxdTN1/mkuRqJuhIUignlduPfH4yb/AEqMtFyYCN+mBxv3AFA3qt0FoMxw9f+9Yuw
Deauh1NlUXQKJ6zJQBHnI7bXz1WwYFBH0ESzWf7hj69FiaS5+VSCeF2qwQ+YGef5vsgluUCyrg4d
zRpXa06AvEl45UanbmAJirtnq/SBKYAK2GOHaKfRy+/P6zBVohjwmY8zUtZ2PUbD9fxk/aESuxj8
sZ+V+IwzEE4Kui+ZfyFHteZIdZp/BY37lnBIr0tTogZ95LnQk1nBppT5x2lebrJl6sZ6r5uLFpZh
03UGTooE0d2Cyk6ICxh8GsrcfuM6n4AjzOHvAiWusNc75+ZOv5w1o9iTqWsGjgn94Ov0+6vRBmR2
F/NUCrob51B+P6kYFdm5oZepN1FaHUazjQLpJIcFcE4LNAL9uk8pbGZvxx7cix3iduN1By5PdiKM
FnoQCfe2m0MELrUuGcbT+JR4eVayUcHGP1g1nVonDOku8GCmXaEkMSPB1np3aEwznL0tZjfnub5M
I1tMmsGGaWJ/t7uR+Y6If7uOJMIOR1cmGha+Fk9icwcYa9wtFVIfgr5DtdIbRtoA3/z1NDFGumPf
g7Mj++NKj3mcFGX8+xt7x17pSz+zyJdQ+nyzfwQ9qyhKNfkXPfgw/a+RK1pAD5N1y+Z8Diwczyw5
xkEj6bi5+AF+JlC0RZJCYiJX0FNBMd4QA78oP7+muDmc/Ue+0LUIe7NxcNYAdfchMKyJxq+Q0H21
wJ6TO9qKw/m4rkVp/Zg0hfdmyCpiu0/ErAQH4mJ7Z98g8/Pk0KoAEq9vLVHDr47o1V6CuezaNAJi
MvEHvmbAJuBqb5gcbK7Vdqf6EqnkCpww6A2mvos3OC/yIELY1q4T4e9hnPeS5pp/dH6raYjn5ZJG
xB+odHmKy+gXEpMm8Dy62JtAmNBeDK2a16hEY1NS0HO9RPVtaqy8rWfMjLOQAOiuFeZLN79MGhFy
MT9TPiWfvcQuEsEYkaHKK+VLb+KpUuG4qmdRo7bi4KdGscA1BM0WJzgoDmjYfVK4rvN1LqCMevln
P9ydEcWX7Bu5EnPznRM6Ek3dkJAe+z33i1KqJcdBbofNRpg8Zmb7BhMkrnBRA8yy6XGf+H4W6/vY
3KprQjsJyrjifxAP/bqb4zJBNbrMyIJ9nfGZrKTN2QYYluaQL9DMOT4jpB874rbzNZk/2YLWi9PV
wYJpiFmwzqcLN4/hzO0IFel/Y8vvGEHW4mWUoXqgePPeGBNhJPEmg9V/Uomjk3/5JEAJQRE6beVg
EBg8MDVIT/JiPolIcJwBJpkjGpsd4QUdYhoA9c4b1gQJu6aa/d5E070rYPvorSm/1Hdj8t05lNML
mXP26zHFUSBV2F166rWNPERgrTZYf7fk5cyOtWXW4iq3hILxM8gZxwoA0b7vLiRtBx3ZnYpfqvWj
LeBiwuAp7uvAk7k+PuoUr3k8Gud+B1OZYV/Xjs5GBLJlgjvu+uFiLwohLT2xbI56/QNNpaXr+Q0W
xS+czpHEo7a/noOYqjHkE3+nEZQD7Ly5vqmVFDOu2uPZ3FAac8hUXfV5ttCtiMoIZCtM6I2JMs51
2GHybDFP8yVoHAHSl0/pFYlJMU+bHsZNqU2w7KqHeJ2feVqgTOwMm6hRT7lW8KTQzXX7DQXOrgu1
kzH5qcbx+TUN0GQElwGVxvgDkwiXq5xlEHO08GlC+qDFCVIdngF0rYCTM7HyQDTEHsDFWb64OSwa
QgBvWInNv7Rof7iYnIDD0rf68thJWoDa1c+1DZ2EfUkiUCl+LEnZIojDU3lUnUmUcMTOlO4yKPuI
kFNvJZAhWlsuJjzfQDzrb7R/DdRSsfDFPgwNOfTGYn5rOVZ80kqZJUsGZfYcfiUqRUHgyqrXZrxF
sxvhb8HkTaSFnsbnZ5Z30O6lUasDhbsKnH+ZKXAlnWA6Am1kbOdLIEcnj0dAxp7D26w+Ogx+iPzJ
LUEQe/6cPW5btf/vNiFryf+2YRe4P2JHt09z/VeSlbNmtosQHh6isxZfC4XwnzB8iuvlgPR5ogju
g/qDbFbST77dhUGHy7DcbbIhktQ2frmTD8kaDnRTcWdTVD2tk5w4qRCTbelYhFyo0mHFq9Se0py9
EtfMEECXN4zyv3OfPLTdbpGmwcy7VOGB0WzxJeeCSQ3YASVsz3YiMGDeueHi76LqSRTgDkmiPp27
AwATuR3oS2ztoOm/1ZobCeRjc1nr5UG3nQxJcCJ/SED0x1rqY+yPkdRVLYfXI0xgYa39kL1a4Jtx
twyaNxs7W035O5uiBZmCstCwhlMDgEAP5O3+a/sRDgUf2/3KcUsqIwT0j+5pFMt6FebdVRI1pZpa
gzDuJO4I8whqSZCxpRwZrfwyN0/TQHq5iP9BcVDLlTc3W+Om4+r50VGV+AKU4T6aqfWP7WMudSLa
20jLib1+BdnbHoYGvybykzzaKb2geAMZ4BWCYB+CE0Bh6Ih9hxhia7kpxeuwCD3b8xSiIha/6x5k
6oxajDUfhvEgBMDGZMofHp+ONB5gx7XE3TLjK19ExVmHa4bCCCRe3403y32M+SBfuv8ateTcu0zv
OXZ7eBF/gAqQBBd/EwPIfosP0gxhuh2tgaS0Yd7OS6/Bih2ZyuybXD27i+Xm/JNnW8nfS8z1MlR1
qTxhy8HD3QqIhCqkkMqcX4asZOkmUDJudhqPzlOA8hRGry2Wxav4zVHmSVOJiMDc6Gw3h3hQtUqW
8/bYm+HasBzATM6qiiAzWSOmE9qhFfV9Pi0vzcOvmBz0PwvoYEB5f/rEklc/+xB8bCnM3GmQUAGk
AhiTErK8VSsOxBrzYEdP1v6fvHq7edyG7yUro/xrt6Hf2mcUTlTQB8zyOV+l1OqNzvllxXhq6jb+
kGmeR52RtmHTYqEKHJfMvFzFzLxXdFVdTuMVlvoPiMJyEf4eKg9YeQxrV7vZuur/vwinpGX/Xfm0
G6EijD6s1GuvDk67ocHPNjxaqwIK5fms+LlHJbDJ6MPI6h9oZHY75yt6dniRlF63UFmZ4qPfHLTF
VwfvCyWac6v/aN1BT/WFoslfT9k3QlUm2Rpe66LvdBbwo+HN78WHp2/k47yxWR4VBDMXVlxRVD/2
WazAPkgUwncCY/KoUTQJuY3mtGRuxy//G4IgNqChDhXlqiQe8xVSzc8m9ReAHcXB1aXeD1U7nm2v
6ifvnLye8btKv3AcQ05HKvQePMdMcjdgKUvN5WRWhp5TKsI1oTWrzaLe/DiGjELQxNnpUxnAUkEc
DpbHjpwwupgBWrsMmSvC0eXBxx4tae/HY9xVudwg6Q3kOHYcw/c6x13St7XxnSG8c1AAJPT0oxvW
xAo2/ntWdw7WPxSlLXJn69wKy30SqlFov5HCCNp90cnzUc7NXmtFfLTX9xKf5I1X99e/n+EHjdN1
lPc+YTVnKkWVlwKv4TPYo9//gn41CBw2Zjvt3YZaW4f1uN6dsobG3Z9h+cxar2Z8ZXPMkJAX+rGO
D7yOpEDWnMXvEno/WtikG3IeV2v2B+80OHoOFFZ51lzJKd8uN/96SjzcS7/KJOvdKtc1zd2qOuV3
Xwft0Bs5pSzVjAy2sa46hl/TBSY9EXQghHE6Vw4YPlHiTeS2bhASMoacYl5JiWcveJHPiHrydEo7
ouvmKByJuNkLprbsKCCtHOk7BJ/TdpeX9K9OxSBoGgRN4xk8b/89lzrC4MMcDoOF4xU/oP1Ug/Ns
+7tJbvxP2rbFNuZsSI4vVxQZxMFPVl7WiYp3fzgbKkJTKgrMLjea1KwIIgvG60YKUv1D5FKoA2Bm
0a1QxnHwRw6kM1hKZA7675IaaTYUqNMx0p3nHO6lVPz02qXlg2Ra3JyhY+Kq9gDYi86lG/Q5RM+o
RPN9CBHXVChY1mLQohGAXYH7rHzmMU1kSWD2xvaFWicg9OdL85WGVc8vCPW1szt0DjcX9CXMuZK/
l5M/1JFqo9KxsbrQfaJEDCyOfwkZ6s+DePkDZlFIv0kZ71TeDcHrRmbMtwRsoDgXjYfpv6xt7bYd
BdPahAMFty84RGMszKJ1m13BUy/X4X14Cj2No21VLiQQiNtL/nGhPqX17KC+KKTov32gSvwJ4fA3
75IKzvSY/nw3Fn104NV7WvawFw83CQKr8Hed7l/gbkG1He2LAeyCPF5jBkSLQtMd0S9x4yunDmic
6bvTCpGq7LN5XzFTWsugmypYPpJoh/axCvYLK37s7UAkUd0s5RqIA3EgPcTJbKwBbWpYReEkqee5
XKDMWW54ncGEmEmEG7mTipbQfP2L6zxT2lcFQuf3EN2JvVXfWXMGvTwvgO7E4IQgUA7RabvkQ/mS
N0Z/ojppPOAwRFTdoI8XeJzTPHT1bvrY/LLv9y49md7tRDoJ9MilCIMvZlp9AdyhyMlyeVPfPfmR
oz06SsQwiJiXRDheVUPpIDCTYihR7LyRtdKzcSPaMTNuTnu9wiy2yzMZxEg0FlrGAW7XyJzBSfcV
MJRgVK/MiKO83qKafWmphs4716nOlE8vKR4iXzVKbTHp8FkifNRs64ijf4Bdp2mc31jz+7iyXzPG
0UG8EzG4iNtASXpJ1AU3jFmlVFnIrZkELmT41AUd9hiBPhbpm/85XA9f+8COpzUr2gLUeRiwvpCJ
jJWtwbXfRicI5lTzUdA4rG1zwRi4PgWt0QVVcUiaARgCFImhOUOCD2sdjcmaazmPVd/XZSwmteNU
JzEmk36CrYSYjmlmOHQjieraKACTUZvSvIqT/8JzMZJ/43OJ3gy3E12p2EWjjb3CKvOZHjDRZdsX
YiadwFZ4ez21frPWQ9vU0ZGKHH2G2d37Nnciqh0ZxvQ7OCRSxG4gtQh8ycEVV+bhIf3AIY2u0a4n
B/+4yseHRQsAS0e+Va9Hw//naBp49ZxXRgM72PzlUiyZsQmeLWJwzTn06A2d/2GorQeSKytwI7ZH
U8xitPOnMF9rmnMGV6lJxDiv0ur/HfhKxlapdG3Z9a8stz1Jz5IMO6pX6IszE20YG1IFJQG/pl9t
IBupI7TpI4ShuZgTYSFCbNz6f9/nE9lLq/t5Ze4fhlCpRiucxhfpjTqdZ2j+9bogD3haTPO9rwDs
r7djzfOOdyqvt5O9oYTQ4L516ogBg/H1nhIANMstg+R7rShGogo/9K+8fSc3x4LbnQ3yPv1cfWSF
yj7mnS3UWw2VK/VXACyyFdUfPxdEraVm2ooLjY8CHaAJKa9qPIqcMKXQMTBpLcAU6Mz1mwU8LoEV
O5zDYaOL8ZqxmChmnIHZRf1q0CBJJww5Bp1VugLhX0Go57tX0mt7ZUFdG7QgN96MXLfhtDrGy3XW
sOJd0SkD48w4dzoTIpqcoZ/WeP4u3LW+PtQWOppb8NeSha8y5LAfOM0glx2Fz21GGUfQlQ6Fhadz
ldQg8ACRZqXssRzHTVny9avSBdDv/Ziq3an2jLM8ZSWaJNDL+Tagbl7Ll6Wkw64Qc86dRmPEzEwa
FNY/gl+rbCOTbl+xtcWW2N9Bg0kwUKuYFTICKHdGNOtaPZctCnuT1viWTYtz1XOXd9E5qW6O7Fka
lewMj2pCKWT4E25Ulw2G7QN3Z7wRm/gpvN1jk0VdWms6OW3UseZkGIwepm4ZEqTGTpwhc1qMB/ku
hOxpwhKxraCh4NwHp1K9jWdaXuo5GGH/3KT+V5LbYcGHm+BVg1KUezzB6+QkAR5CMsuzYqmvlvJf
b9ZuBVtkJgTGMGcLtDYJEZAFUOT3bu5GC/cYMPNhkVUBzdmwW3zGSuga8vX/skCOiLbQLNL8bvm8
PICwcEFLMaq0y6wKC2+OP2JQbD4IBwBKdnjV0Dmhfqy80WI0wSFRty10HUq6unxkqJDTXgaEJ2wx
1eiCglO7bkJfTkoMrOgXsVyhsv78I/DPmSi9ZdnmgrPjwAfsEK22zs0KB3tA8DS3v+TePxnrpySX
rm7rbygUjh8gKtoZNTGt+FnwdF+yKvu5yOs9doebYslFz9lT4vqhMrne1GZOuEzreqWl6whPdUDj
iy4FtHMFBFDY5JoQZWPPbsPUCPX1g3qkG/pvlar+BJPgkZlHC75BKfdTItltqhdlDSFOy2TRCHBI
XltN41EgIV65txaXzuo0myHTG8CoNIvW7dYGpUHtbBXjco6fpHexocn8EuMPrLOKqM8GUHMhcr4d
CLsOQCVqeykCmH5C7Hi9w9B6fCiS2czbY1iAwKrfRoNK6wCu9uzmYFkX/s41VvVI9BoPhPtwUGLk
SB8pqcDqUlyQlkcKGtfnUrIpzH/bviThINzzI83dJ1cHp/cQK4zeY8wxvQ3YoSV36v2HSlGoRugT
wPDhQR6HHCAmPrSy/KWotBEC5sw8V1D2KoEiUIQ9FVuEs35hzZr3W2KWddJlF0sK9yIL9RbQC8Jc
7hAhxivpfaGU9SV0pynHMEDxTCCGrzNXermoQt7KtsFPRgeUP5pHrNWqrEHeFlKahzkOdN5T6roC
i/maa6MnUnzDOWKKVKh/MiSIZjHHM/VO8QmBX5sxGS6OUzngkB5awS9PP3mWABwTBq7Xfz1t+q/x
vr4BiMXPxquZ4vPP6MLTPen9GExE4OIo8Nzt0s4kEI2OFRoGey815sVaUQN4SpIA9XltoyBltJwf
dgKbeRp7XxjnEq1dDuKzBiysMyVzkDLf1VmY3v4ZEDrpziqEF42n3lntf6Bj0b8Sq2Z5MpBUd6GH
Eat8+1FzQyHSj+TQddB3HpwVfLCwtUx7l8/0MozvOlnSetlJM9HNh+wgLPa9L6DfVrZd0bbce8JU
nZPfUJBNspCoptD2aqPkpLdm1yA8PU28GQV1BUchoceVLvvi0LmzsvD+DTMNTOJ8tUK3pkR0+7MU
gwVGnPi1c53H9Vl//TZy2yTSJrKvVVIUrYhO79SpG3GiWKugT4t3Duh/RFPsowM7hITqCd2a43f4
XTZDbayhOVHM5h+YY0Dc/lU6P9gTf8UetBalmL7JrIKTgxgm39mxTPxxjPTVYGUHMRtuFmPQy++4
Ng1y0MZg9zMeLsx80dxozcVkJJaFdGVm2b7dvEBT5fnlA6tkOpcMKGogYDhDJTnbSWEWb+ZKR7tY
9Jtw2wsw78M4C/uVpFa08hsSBWToZXEIV5loiYgpEbvXLaR2gwk90MN70cOAEsHCuIWt2mOZa3JD
5cENacLRRaNSir/YfccMMBl4HPx0pjIJuaH3nKvRQiBhjVEH4BhTb4rWl30yUsNOgj0JaPA0BgM1
bbsi7EyxxeSNPMesPqB5Dsd3i7ahZB7EnF9xgVJ6pp9NPtNU/V0nXykWQ/hoaScylKXvJr7r2qLy
X7D/UamCVfzm63pUdEvSAEaK+jmJGpof17yc0PwzWlvB1Bd5C8Hj6Y6s4TwmbYWnKCIEBLnNgXQ7
q1dWJqsNPHzIKA2pfH7NYEgTD5i2BhPT/URossrp4LUVSeQlSDu9Ppa/Mni2Bw1E/guXETeuqT/q
4Eo+nH2XR00x6tbKNE0/TbodnXfOQp/OvG3xDw8Ok8xC8kBD6P3TBQK7EFVXzawL0gcBcUik4z5q
sHmgP1+gqN5MV0BcEmD5iciIeMP3hQXczghsdYCYKx2c8gqFpkWrEtDt2oGQma0/usIqwbPUVvBm
QissN2940v/JDDRxWmbXRtpkgFXKcuC5c0jawoea9HdXzbrd4Kz0SuxBNqrrTJY3VMHpbl9zxMit
LdarW/fNh2Syr4fsNX+vL9rQdp2hiqzIL2CA0OQF9N9bePW5Z8qp6f5DnsB8t5LWM5kmnMZlv2DW
S7/3taTGspW1KkHF4Cgios8FIEkLUKWHHWui42iC6NbFDnFU+LbiEmLD56OeDDvEywUjxzjGng9a
pKoEWOVIPVHfLeE5nrqNGGOsSS9Np3LWFQw0CJM25qqkWm3gFiGbBPlOXc+/nRbnYLcEZE8yYqLJ
yiM4m/X//sspxAgh28EkoMTAfdHuExipqD8vPAqT4yuXpglR+UBPsyrRH7x7Bb+DctGhBGbFGMEk
pRmYTNlTGZ1c8ANsNM9Iyfz8sK6dXn2uHQmz/bQEXBquijzu9TeoAZ1B0jH4qORnCFVzM8geJ9dj
2+Wd2bSqn5Qe6jdbZgCCHGwraYY8PEL3/n2MzKphsyYL++ksmzPm2/3xiQKdtw2J161K5UezRoj4
xtDbAbsgeKGakeppC5ZPoYj1yZYr+//H0i/RPhInyCuW5rTGgugmUVtn7ec33gv+xdq29a1Q1Tvm
gV3w5kitaHn0Bnk9kHzwQ5ZQD59h4C3SgSqwcNHvKJViwAYkQ+D8xecwSgxuarQa9AgMcyMLESsl
Dukoe0Dz521iKm9pcS5NO97GYtdsO1QE8yL26lrenTyovuT54CwOQ4ihBjVETVBEBJqIJ/kg2kc0
p8vmlzm5UrX7Qj7eodDXZmiEM1zxVi6EJhI4gZrk6d1isY3tKoConRjehz+8iaDh5oV/FPiXPfAn
XjnFAr/oiE/b5DCCRmXdvoYR6JSZp35KwTxD2zL9l9qjMDjbZLCrIbbR07inpE8ywu2nYSTUFJcn
PCEP7fz/9tOyat5EEGhrSDIviOx6zIMeZpbXHmYM/zqiBqdSXHHoZuNwX7O2nuGCBBOsHWRBunpT
/VPW+szbIY6PDXSmykQnv3swh/tmgI1u0rl7BGRZJKlCzrw08XSqqjPUmRRbxMey/8KkT0XtKuTU
BAZmxAIwU3OgMixwTyc7mjXBBF2hvy1/2+kSNbyVGgqiD8ZH4URDVF8vx4CAQeJ1Sg7+PgjDavAX
oZ0LcS5qItZgODAuMuk4nagSg7slzFkmMMPhj9CO0uKIJRpeXTzUlSDa/rmGeKKqAdxLafkhXDrz
W36scn/Jf9jLPo+Z9TJAijIjeLxZ9KEJms/nU2M9lYEWlUjAO0CmelcJ80SV4sTGO3mMCPdPndE8
DCLJr53Y6zh0UBGWKkIvGJl2a8fdf2zISWp1e0IBhLyziDibrdpSmN4NviZz4jcTh5b4OAFyXMOc
7SKaYPpW43gmDG2Sfx0BXiA1ff29WkR43AvSPxbu/DS9lFy2FFhgMPUVP+mQydE54F9dFoKrfGkn
UcIorQe6T1eZQg8KuEWf/NEqJAuH3dQ+JD+/sl+V/p5g1FRJfs+8CxwD2Aj6Az3yisecrnWu34hK
s+xzUD2OtWYgXmww/1yhZtnNNv53EZgMTR3H+KcXqflLSnVyoF2m2IhJ5g/EuLOR8vFZWpNhh07P
lS17hV6kbVcQle8JFpnMZgqyCUZd/vBnj7jhdNy/okPawSWT2tWetVGNITi9h5jalEar2SwjjBx+
gAAHwMwTNMJS9uLtvFqz9q4N/AY11W0fhC5iVW19Q37+ytYnd11KC5KgZq1FNFZFS0rbS8Q8lMM9
S2E5As540iBP7SkXIxnt8yOqWG/sazLgnE98/1swosbluMRFiKX6qlIJzPmZZgWl3atjHH5ckHN8
UTRUpWJ9BAzLGrpLtIrhVJRMbO+YNsDBhsbe/zvof/Ik0zEyHgz6WORUvT7Rz3CYtT/pyJHwwRUo
Of5oDSb23dqhFGakrCoZJ8oNBHpAc4OPxetV+vjelwbGHv59zCajU9oQkomzUXnS8SMWfaRgMfDi
Tj/u59qrFVM0p7SqiObRDIAeZ4fInojq01vF8QSBzhrHWEPpe0LT6qfbDz8isgbldhYvpac3r4hi
A2hyF9FPCesxvcw10lve9C5lnCl3pHJmFhUEh+GKj4RLct40Dgeg1SOCpC7L+cxpT1DfixwrFhZN
kKOGWBvwE2oBqVtQyASvHTGN7GXdu/Rq/FinrjuIw27ClY6qq2aRTVfruU8dagjd0c/yo18Xy2cz
7W5C4vARaKHPw3a5/OZG6aIv6rfhtHOBqRZonjq/WDXOeqCYkFdt/xrY1urQPdZaJHa3XBzb8KcW
+rnkOvlTXTQ8DNY1Ge1qawO9IFcUp6J6DBuZtZQXknohCZMBdjOhA7FhS7Z4mNSeGcN520gWYjtA
r902+Pn7Dgtb7zkI2UFtOUogIjT8Ye8TF985cOZaWYZRVPBbhWGbCrmTvDauIfXGlMncHefeQhwa
ls7jnmMN7gtB9qr5GK0FRynYWBBhpRH1+Lz9/EV32QQczVDdAE0hxB24iYEm87I+DcCC+BuXLJ1G
uFeV8lcdN7YbQeSKkg200+n4gZGshl+9Y15+MzPhWVmjyCVH74HN1kwyNG0itBQLK4AZPVN//+RK
f4O7L1ZUSfFme3tFr9FxNtM9geebmFq8K53AmJU5BmgYM7WevB62f3ewlVgGLIKVeh+N8AiDAlU5
/bfjb45x+TzfwRIraFsPCAOb4pgdR6WcorvtO0TP5Sid9ytd+drA6CYA/PzerBKLrbp7Txem2d6e
YpthMjDYAecVJKLLPRYnZW7mluh3EZlIFgsjVU+FGnYPU4O4QjmP9VkEYUTdUInOVQio55Y7s9Fu
VT8RlcBOL8MFlxm5oUDdDwdZfF5z6ckuFECJ5x/MntdO7bqIk/JF1ocwnSaBIDi94zufweyIJEhg
fAP9dsHgvmmA6Ftv69wpxyX5G1Ppue6lxUJl4Xv7Fn+I/Gm3VLFQp/E8EBiLqqc5jRyML8+aB32Y
egj2IeSpkXwMzzM4APux9BqhFYD7TyR9qcMUyDPCnhhBbbbJSWmAIUv2cND5sHaKpAOsx2eTp1XZ
vK5cjhyjt6V4DHG6yLYbWDj6WoRq5TwWQF4OtR0zIOmo7+e55KwmBUVhlRbki3lKgCiPYEBmhPYp
u8+OTf+K29RECltBBn8qPtb++79UMnEFYt8krUm7VRyrCPSiTw2uxhfowfQFDRSGpjD5Ufj13cqx
3zZOu/xfByTAOlBRgOOETcYPajTvmOTl4iFo2zUKIyDUZX5oTz64G2zk1o4q7hO8tSHebQom58OG
5IO4YyM0O7oWEFl7Wg/kwUiReMcww1wjow6uFC2wUsXsN2JZlwAf2IGoAgnawRj4RDGEIg43PMv9
siSdchN0h7wkFGEuR2QWH63jPn+U8Pmy4uVBOkbbpHf2z5C7XEZ6EjCAT4VbphJleEldp+dlAnaV
d7e67zhqaqQMZzo7TdTz1h9lp5iR57Kh+z618LEvkmPOGXlf7n8EgO8Lkm6sgGYE/fMeruUH2R1P
7LSVLbQtij5gQ2OdjRx27d2fmaj5FDP/b5M5b6k4XOSHMEKWubJqKgZozkabWT3oCNtTad0q9I1b
fW41PfIukYYWHqlRQGfOnUs8YQ2cG3paVUiQmZHRdZuCf6iRr0hZAL5UMlJylcVsJSLlH1Z+29kB
pOpgbZlhDUOxPJmZs2S4IC4ijtDBkSknoX2P7jQSgiWiq31BZ4cm9YwbhjayYoo+FaB8rVDIaCzt
8XsZT2bTa78hm7k1M6lPNV4UXky9bgxX6NUQcZ4v+Bb3BZMtQ6suZcuYDsFfc31OLcpW2WMi0ZhC
qaJzMcF1su6NKWuRT7B0kYhqS26xXu3LUC9rYBgnmzIxPnOEWjYvSlcQsqUD/qB9rI9S7z3ei7FR
MuRwYRnRjGAzLiNR9RCB0CrwsuaX8wm9h/jbRJX0arcQ4jtXAK33IdcV5I/BcnSWlh7ch3HDXSbF
jG7hz+2aYE8nfQ+jhSDKOOwIT9jFGEvrWImOA7JrxdiZb8zr5vDy0JW12A5p9DPNZwCg4ep2v3Vf
QY8HILwjK29bZ05AHyJyXcypV9NbJdnFRMGCAayCmDbiadQMmsNs27xgoPSwNw3J3Z1VkrRxpmiP
LUKjMVWUltBLxwEWuJRE+a/AH1nCemGQB2FZbxha7AMBzxgzVGH1zsbY/NI8bXPDfYMkdwJwbBZn
bcFW9XwaMVkWRtlUlKBcCCyMh4ASkJX8x5yBcUP8NmJ5leq3wZbU/YP1xBung5jOcfatiRO10U23
QBj6YPK0Hk97KpWcMyYiETeRXoLYne7/WG9dHl9f/35+5TcKexgjta3iGUub7Lnrv8SvYWxu3aHz
OpwLkO25Ndc8ylcy85hqKn3+FLUAtfE6kf/D8O1TrdRe1kqy3llzxEhxsdD+9Lf3Rdk2Cc37RnEx
uRDWWsFfW2Ejuw9AfOKlhf5w/Ap2R8hiM8QWsLHPDQUGrPHtlWS6YN2Cen/LyEz65z+D0DYhcgkW
+6SOfhfGeFKabEBUwa8shpKH29INNGnoKtE81tzzNdSwjDYTw/esLBe1iDYUmzLpEDHoiUDIpRqR
yeyDN8w7uRPAdDW29jQg6YNpK/NytKcIobPv+V7f0o5UKYap0v0XPNwxJz1yTiIsBtuCCrx6rE6/
V064rXbvnKYVxx0c0PoK6MRmD/1pJW4Fy+PNhmLgdHCge4F7KACAqc64XWSiKBrsMtP8JsyZfJDU
+mz6qkKc8sggYo8thJdfMx9qoz1GmMCLWxb53FANU6IpmuL1iB/0zNVPIxNS7/iWidWYIXWjwXo8
trpPkVP7Hq/sztXUeEAju6dOhv1x3rUehkSRnvtTNPYz8P1RtBRiacrPem97ZAO2E0lR1471PuGY
mBT0JrplM36QE/Nt2ZCFDtacSaO0tQrx6TtY7xuUHTG66X/8D0TuL0KXa9CLMfnwAU5+wUTyaRkc
2As8PMIuX1OIZMWsKHeQKbjeJ8sRdc5Kmy5MLcbhlqAA6ja5oYjaITejxHTUR0vynLbnKpTfslL3
kDu+BOw6izMQ3BXfJAFAoTOPS20FV99s6WO2MRi5NhM5T4hYpXGuKOppqAlTmFa9Tg0M4fJRtH1u
qiOouoEuX5XuhWEGPw21ul83amDL/rfS9nGA+3c5Sv/QYG/3XM0rp23Hw2P51ZfsHvXbbPhpVBbJ
xNQusL7qrdrGrHzYijCMxc5BVOImMc7+6Jd7sXpdGSM4nqq5Ct/fJUs5b7A7a211G05aRPt0q9oU
b/FGlgZvO3qhp9O3RXRtBfBZKi44GLizX/rNrkVuPWj1Or3bmiIqI8rvB7Ch+n6Wq1MU9Zz/eCGr
BqvqrIxCJCrnIKZljORetXiHGl7o2khe4JSvHE0SRXlt5X7vDr1z+hnjWGEKzLnTxxabNblNxyLd
vAnik8KJc1V4ek/4fl4KThXIM18joAtTF8OFXMdw1Mm/OsJp8qu1uzpVeziAyMyLnvH1Pmg6ygEF
adRPA1v0k+fYzsHSwmZENgLdLoBWYhSqEPUtqTl5BUmwpyhH3G6VeuG1qo9Teq3RqsRKB17oTtPA
rhGufyo87GFXqOizZ6FSyzQRTd8ak4AjqcKq52dppG5+aMd/ESAncVK4MQKDbClexjaTxCFZxZS0
kxneEz5Yscu9HwA6hUUHUWFI7lESo7gAQkzz8j26fqztnulbGq+/T5Z7rHeZMuRkA0N3vmaJWhga
2eWtpkyzeUZfc6XLIZVKosxL6PoFpAt3+WnLI/U2rWRaGIJLkuChLJjgFVbAXEm6JL4aVa1nZeEZ
/Z/28/UWjA6mSzJTbyTWf+6pO5sHToLoPk14RzfJTApwvCNhX08WmqUl/imx6dgRd/33joajm6aE
FZ2dXmfBPyyt0OBRf6a0jTZ9ruaIN7SpLJExUH2J64ageWwMMIafgGb3eQF/tzgDwsjqOEREzVKk
Okm2Zr9IYzyzauKNxTtkLer22p6lHUbBezm1mPADVqNPRCSncFhm5cVs5J8/RWL8eu7P8dPWrYpM
eC1H63OPIK71S7uW5Ve0PtA5W+Yr0HCMAXoRhSdBu9bzNdhjbzWVd2UOF6ji7I5XnFqbr8o8JOTf
cXOwSaINu1EANqwEVfkxlE1GgvMNSAYzm19zEJOrH7R7wpzoVXo1GOgBZ95WP9/nqM7+TcxDOJ4j
vnGlX7NiW5/A7gXwd6ydgr3PhQG+/loYvXsIezRaH2xW+v0rWSquyB9+lsSzJ+m/JqcHAor+WBwW
zozftVoz1JO4PLb3aB1nur5HF2huYg6xaVPWaV2Okq07Xc0Kq+Cmb04nr3kXiL7FJkFTJnk7oSJm
V0hxg2LjH1FS0h4ilVn7hh1albZMBmZB4688m4NO9LlF+KjMmQ90l/Tv5+pD4SBsHid/PWRLy0fE
KoT50ZKGdqLwMBTOeqCNMLsIPy8eHazhmbr2laCfi5wy9nrmUZhma7EqphumAxHTLfcfkt5ws7oV
aoOkS4DiptfDKheYjCLv0fqVhcrbmHIHKRVaaZxlCdd7dsxGSJZNhXCH8smrSrsO7k2JLYWxwnd8
DoaJH7AeaH9dG0pVXzbxA1lUOMb060CX0zyucP7bWGMyupS4WWJogTm9YxAgddjBEZqmBnAz2N9y
IiygOkha1E/1CK364S+bEsAKgaAP3IEh3hAkOdcaWuVJS78g/mSfbmMtlAW7hQyTx5mto29QonGQ
SA5B9H9nv7F9NWHhR2n/yl1DVIJ5RwPgEcjXsMGS51hD6rogZvdPu5PrLrn02ZWkT2EsPTewSbYR
OHy/bJvc7rdqamdZmKS95eUWr34NgxUsutMk3pfIgcWACl7yByTVHr5W1sqrTGfoIejO8Kts0OkY
dFXKM4joAowkaZn3GW9uOZE+uUTlpX1VRoeOoocfeoIJEmJoOf0QYn+ZPERual+adLieuFk9TjO6
HO/SlkU7atKRrqkF9ZnlKq9EqssVsf7UOd/CALT08HvDiJiWtCj0Jd1GnubXDsG2TIm4ifPVP0PJ
LknDhj4SHQJWaSCkXJHXR5t8u/Htq1bH01fGSXtXMxFMkl4ZXq25hCJjdgUOSGfOZ/Y0h4wSS/4p
Gp+zXZPuKjJrlt12K5qZ6G3EBJgpRdw3tplWQpPB3VtODkVuY6rDh//6xCC+YHc8EJyRWYKtQdR1
b4/KIysKFfzDjdcQJc91Ot39n1YrNwm0ncEBHuB7DUoB00QoZ3QNfeEYrzi4IjmowpfxK5NTEvhe
NZiuyxRvtflRfgi35RCwdverGAKfAy/Bt92LN2DG+q9VCjZuBzAvZPi+663AfYdp2gu/uR8VwEpL
rkHC2kG3xKhWhWwpx40llyOdiBQiQZiXEj8DwOUSTangz0pwEwelSxjediws7Cr+/g7GOfLLOPkl
CfBkZsljTliA8OF5j1MJeBxBnH0sOVwjns5JjmhNNjCpEZg3y1J82lppRlCgO6UyXq1T17k/ABxU
m0TC3L6LrRo32tHZoSex00fPXDEb272qX2c7H5QZH6rdM0RUb2td9U7OPgm+dDaNGc5yy1mk60y5
IC7SJYxPySuNXydybE0pAgLAA2oH+rRaMG0Ul7Z/HxZD6r67R1Q62893ka/DOjUCIJ498b/p1kzE
eonTVZcbK20n3w5FD5wWLmiPkuQe2spKdLG2r0uhA9dXJ9QK4oA01JgJyoY8IP1KhNvL2jIvpTwG
ySaNTc7QhfSBH2TGAWOGuxX0o20Eb7HkPgLC3n1q4KL9tt4tuhlepOABXYeUUxgFC4NTyHq3NvEr
mbLZUaekk7eZ9AYS5e7LeAab1sw0VCWZzOojAWotLQuOioa/RI6MRmQkYIP/tEuBgIQRyJ7llmuA
DGR/3OT2AivLRKayZWCSxgvdNMb5y+lU7f7f87SXVbMlhFBYucGQt94L6OcqduUoiZNez2RPtvk/
hAsgTqjQMO72qNB9Qb6olgCqzHBls9Wg7v91VrTZZ9OmUN0GQfGIJ0dPG9+dMhr4WqNr2dd9jje6
1nyKOMrBlaBKoDK1AiutlJzVJf7/X8s7MFHbs6NZylivAmr82s8jl8MbyqwyWcTHjnc0SIszCdwH
OCJhVCSCsZGaYnK8OeAO6CMNT82ieUeoTykZgQzJU0azleDDYCgvha3hXrVbhL67uPomTiahqmMn
c0WqLxzgIz8k+0sjAFPtFqpffLVeq6aI4NaqA5PAgdY2HmgXGROYU8fJQUV9ZYftmvW91ET2jPJx
UHVMmgcamFynGjiyu200jKcVx8JC5t5XvM0eUUuNjKUgVQ1uGfuZ6LDRCL+7ts67ntpMwv/xeexw
Kg93SGcF4pGNu6C5KXPRoKQBHQoWGQ5YLX9xZ6BcKRNGYI2H+kXZMNdvOQXPcLQrOzsoM1j9Rwra
OyOfaspLo1+6xacQBLJOYsOe8XscVDA5Yc3aAVHJ9diWQXLtgENadVHvW7cA6w7ZkxLCeTPoc0Pm
cj4nfgJJmb7uNyABaKNQkMxKNjYu+uANfeGMZYiyphIqitpBWhPIJoTdk5rZcuYp2JqXiuC0G/Wj
SJe1HVvsDColW2H16bZtCTSFBdNQXmz6+oSh9C/kJ1+T2CUUU0UoSSHktr4YDCxRwaTfxH6CdWos
rgov8b2knyZZmFWEEOy8KY/hxneaejMWoQD+vl/enjXZ8t4oYgg54ywVycJnWZvtOYEn1qkxCaQZ
/2pnB8vOu/zOiknqM4l7PFV9CJEAn72VFLXIlaA9Pw2rJsAYbT7cOLE4pE+BAmqGiF7csrXquJfz
xefE1MWl8hk7fBwtAB1PMUj01pmLuo8Rmd+fQNNVWWQAsiTzcInjv49nJCywIHMwfOcmZNLQ0TiG
H0xtQvM6ngR95NZDaaNuJ5Qsgf7VTRPCfkLdJ6baFmYxn065/6zoOqDIlQe1PsMmjjxay3YWJFlr
6fnw0xmF1wZvBWt59d8yibHSDifH4bCLTkRVIpnVdiczGwTemzlcRWhgCTUmyvbW6FYt2c+wYkPq
2JifPTSiez5GZySJ5TaqaXteQ5/5yrPbSBvor5d0b4rxkwplTaCP40WMIkpywGRejV1QgLOKnuXD
vlq5+uGkIfICFUupV4mWfYOIrNfPJONGsR74mLxo2JPSDPIJLdUQmtEOE45E8VyOw/g4ZJBuWnQG
WpENaXtl1TsSK3dFuPXyVyyt5G9Jbo2w9nrnMQsHYH/6pLQ1smK9uvYjC0Ab2+Gzddh0fqICNRyc
1k9eYh2PVr6/KpGRoWF74Y3++9zfxwMaa9iTz5lqTXUmcx6wrRDTBLhK/VYdQFyUFjTMcwY13u9p
TEDM+h8E3A75JiA1S95cN+zJqpW8sT0u2JCT6t2R1u8YzqGAQ5myshLAQ9hCEDj2fARIIeihL2QS
GWd7EwHAaH8ZlybYS+nXJ4fcY0+GyO70waG3kbaurtqvCCSFRApln0aCILBmM7+4beorpdYyaaXv
15I1hRqgzbLqKa+n4MyozJPlmImG97ElNpKhMcvHSGgp9nwePxcHC1BnpRWAiudvMtyxo0m+R17z
kUX2x1zCptJXZkO4kO2dMzGQRxTlzlheVdS4VTYRqJfeZsO/sWnhvwOdDHj0MlfyX1dezXegdYp2
5+VnjyZBTlx4tiusf4cSox98gSYQRPJZsHa2yjjEJS0fdQtfFmGuQVsl4tDYzZ53N8xzp2b7fWr0
Xme1hvXTXIl0E3MPzmQ50WktQPD/seSFs+JtdTkbSIM/1aUxez3eQ11VaTH1ab49CcylZ+ZDHx71
j95i8IvwNtfDPdCMjaDUqPe0FMRpa0vRfIdO+mBbF4XLDYLuA1xRDr1FZJ4VMHrFrawaJqksTPu0
gQHrrditRe2k4hZvV2k1RPCAJrdojq1+TCZVP6H9Mxq8Qlcg830lZ9C9D7jidSnNSpDQQDGFBqDY
2tHJyjZtTDMxpJv/zdgzvvOzhb869NrAKvYgsIgmiSvZ+zOd+P55WLpHXadsX38a2owSJK9sDO7V
XdY0BZqIb2swzRat5P/iCFbYAZmIZa0AvykxiV0/1Ta0NaJydJxwViNfM7VWQg0XTO+CvpuIHPRU
DDF2UBav+9aGQl5406quOq8QAwuckRuWMkRQAKq4UJ6vX9OTfedeRJA23OllV9KGtJIPW5HklVVB
itpOl2Pm6USx3P4CvSgFTUizZaCAM+YoLLybXa4kxVAoaAljoJkcuEQe6GTd1/bWppjVPutNJRbv
itHuRPqaAmp/WI/F5i0X6Vt+Mrd9zlRhnySvWiZEJP8I+RsUx3ezpNjDw3MZkPmnHS32VQLsuUIX
ooJcf4jleHWIdatR9fTpeEJJIgeuOOWgs2x0ZWypwUpPvRg8yM/NYU+WRX8AbUmjrwuXgLF/YSO9
j8XM2SQ0puaLI4QOylJ8OuYxLyzCZT/DQvQD7NbMIFJyAFHbnZHpwn0KDBJjdSrVZtVb8tCDH5fq
g5t/I9s3I45+y6g+iXY52nan7N6u0ezSz4iqbvgOfaRmcqCzIwvA2dmLUo0GNB227DIx8lLpK6Af
dMUJafWDZOIXOpjO0AfKz3vcno3+EkWLKZ33lYORtnG9bLhBUtHux5fVkPGeoRfQyJ8LAOEBeNRE
rbGqOrDnm4B8t5vo+tEgjSh1OeRzON+KkUCgv8COLtzfDwItJ3r7elHnQ4CCZ3ooOktUja3CprAh
laM0nIZW5i6LJ90DSl/vUf8MvXGNAGYLeWxDwUhTQKm8lt8WJ6hr1UUe4kK0dFWD+N57OA5A7f8W
Qrm5dZ63E0+A6AEb59nkZ5aRA9a9UkG2Qxt+Y9dfybec82enYF0mBO9D/K0likfa/4Q+eWheLYDz
/xAgwRq6SdMmaFgML3p/j+u0TiFGPsvd65/9zIEj/aZiSDHEgMVRWpjAVaWHplSTuHLLxrs4awYw
vv1JE012P6488UPnK3A270YZFz6icmoXGAATO9QLnW6bqDaWwlUDRAqJU72gokbhf2gICkvIZeIl
L4M5AmULdE93FiSp49kQ8ljrOWU6sN7QldSJYA1FF1QpI81xcNkpvbg9kLoGX44cv7pRJkDY+yt1
zkcDxbP2wP+38AePdDdn5t5o7RrHNy70UkxTx4omU8Y6gOGA3uK39odDOH+FassLxrevJCmvGfVT
PurXMmRgBayJbPTzeEhzPSbxIGsA3HsN/9TT7LpqCTIJQXhw0PUBmgyDmCoqe3325FrEqYmABGcK
wtMxzoxEBc1buIkWdnCuqAbLuuE488jm04OY9gii2nqPV0XpN6s4UONVxQ6TqcHfdMX7/DHhxswY
eCIGnkx9wYYXSmoPNGxpLxd4KzlkYcyKm8k2uNBydd6fnsPHQLXh6f1kpfG5XxNGb7mzwrnU3foY
mRLJspwpoGw1PxZxyakhAaMajxLJvjDVYs1kbNW8zbRpAvRuejV1BEN9uLZ/5B71RkwrZqTWw0Ny
gCo1iuGn9VEmC+WOhmWVMckYzSgbewvAcfNkmYWnEZsdiSVo9OSZ6nK0k9pzLDxQcrlXKrnok/bF
GXRtv9r367JtIa3UpMGt+bk4OCkfq85yPgAdGj35ZwWNflkafazIHG8F9Qrc891KapHFhDyufxQ+
2ty5fWGLQkpSKs9IbUSkMEy0HnQDIZbDeZF2z/KMijJ1yyh5VhMTKq1jGfnsvup886KctCN1fAXQ
LKxDgtPdoNA8M4LhWnTkgMAJAax+d81PYGduOCJ23uN0IdmNI/1uOTu8rhW2IVaZmIFa/psTV+UH
GNh1+t3c1ceUl/RtNxkAfpfBZpUXaZenasgO74v4l8wANGizpWgLJrtAZwkR4SUtZnSKVi1PbCNj
7FszV4xiJ4YSa2Z2xcc2NxzOK19FHqv6l1l9Uslx9nIUfALyezK8amVeT5dLgFaEPIam+QIo/w+8
rXgF4I0Uj0ohoXg/BuErjRfp8aZHjmmVe/+JBFaosoEKrRRZ/oDzyivcvoI/XDnsD3/0i9JHaXeH
1Ixnfn5NSI91PTVfBRlJa1tfxH01ZKuha1J68UwQk4aV/RgxiH7Gyce6vgyzydndo2qu8uGxXGqG
GSwcQMyHwW6TrsY1Fo0a5m344ojTq1VATSWFwmYHHzmhah73cm4MPQ7QtjRfS9GIsUc6qPmVYb47
T/QMf2gK/D2yJdmufTD0vKZIYN8fPEiewavNS6Y25Qc+UiHque0QCNzPEQhC5uYJodHLU1ayxZjp
gr3yZX19F7j74313tVYBmd0HL4Qhu/f3yLSTaDYBdPf8rdJDSG0nNyjJ/S/kccZaPv0NMxjdcJlG
8Jl5j30dNkORuCrWbaizXmEWDArO/4k/tTSL6XMftes3w6YNLyIifrlDgIoVwLcedqOgXqrcPqgH
fKIJxhV4uesRQE7o6bz9l75EUG3teiZ4Jibkgn1gdSfuJ72T/eGystsYr2YCvPDjfTGOsKH7ej6N
eiWr9jIWEXNr+YCtQUD+WqwYMOnayEESW3XVhKfktu/sGqayEuSX+h0BRqFjMCG1NqmFjI5uXzN6
WaJbgTM23FA5CsA19VR76aQyy7RaBw57KGEXq6E8aorVGKHc4Oz7ewiuolMV0G/bRk/dgNOQOqxC
zWb0hmO51O+Y2aA41NxgUvcePy4EwhZg0aBT0W8WoRdG3fgTPTciINO/zBBf8eshfKgadzu/b/0M
Okg68ZoiWUaNCCJZ+wYf9AY0egeiiZl5jrpm7zQAzri0j1N2PlXgi14Krk1xfDKrwRlGBVIuWw30
jfFpr4dmKW3oRA6XRgbYBSfJgWp19pUPRDKMPuvPplIadlFJP85X0hsOZxlCyzrf7D77usGH2uNx
FYyjDTRoNL1aZwt6F+VFeiEXoAQnefdyk4BAsPP/pj5WB4iBJJcIyaAih+oTTKThisqeHVCMVhNS
2fxz3iXYQBRAD6RTNpoZzNwz90dRB6YBYBbV9E3PPwl3xMwxBmU/kTe5zVdkbyGka5oB7dHNjVLo
c0TvOqGRac5E40nqWNSRF6BV0HrIb72w2g7VMY/K7vK4vs13341n9/QnroyKG5ElLCCTFF/n1YBf
SRZt/sPNV0avTd/teSr+nYACejCkXuMar4Yhch5D/qdY7BUF9pcNSQoz35HkZ8xZcd/idldErPwR
LiYqmT9VdCufoZA4UNghr5x7ApHeGID4lfBD5FifKuqx7e551r+G7BRcyCJeUItz6ayhnUljV41x
ujSJvxbh1Ryw1z/ObK93YuQJ2C+oQAJH+UbPXyPv/uJqRqG2LaWjfMyhYBykMENaREnvuqGhtaS7
0nx1gCnAn2BtBjr+Af7/dmrGxq6gyk1sALrYS0nIUITznNqgtGLN+fjOF3ZpAuoGOiK3m2rXYTMO
MzK/qN9AjaBUQZ7Wm4KQ04CoeSBwh0OcKpE2/usF5ZGHQhG7WPTnSXqZ6lS3nPLWT/IW6fich7WX
mceomCShFjEd/YWp1WsRVhivshT4YWkY59x9ceIjG1tK2dBSloxdI02bXq0bvR6LdcQ8EavZnOKT
ss2CfHaA2FpzWDX/htfdTWoIE7B9bJ1F9NpLn6YX1YIjKS5NqwtVNwKQNQ9SMMKFtfUYQBcUpVtE
0qFXjvLt6SGyU8gK9dNA1nvciMeTi8aQWnGMVkJ6FnLd0ApWSpIbRV/W38QmTBPJpV6YMT/kGo16
QLFeOZDPczXq/6UTpzv4mGXtKeFaZcOcihZO5Wzi515Kj9mDKriySRIU9xOdT5jtuw8Qyapyi1wC
p5phWGKa1P9ciWJP6KPg6AoSGdv4AHGPbatgv0PAUcc5PShvjdejZyIzVblleROd+Hs6kBJ8lLxA
CjTBqkUmZW12uN3NH4bOK5KTvQP0vC6igY6fst1CldYcZBWdi6fYHC0sRYQi+c+WpDhdNw7mJFs0
HmDiC7Z5+jdgeqhRQEEzRNXFsEexe+wtyooFtDYytduIzq7M1QlIhvDC+hvZAXMHi8ay+C7hKz1V
ItXJtEXtrSvZxqEKQbdXRbv/pFkHpwSX1yffbvKIdwZzYGy5qCAGZ6D8GRXxLjyxjZU/cVO9Sawm
SfUUwVwzSlh7mSJEYPXMiTV4mH1XeQGRUvQQLFvsXY2vpQuSAbkrlO0Lge80moWKkzVfxQkos3TP
KM22Qx2nNmlibXVPmDhABbEsqu3GYxyXz4B55xt9XvRb4vsx0ie5jsTU3AkqRlz7bqDyt0NyCyh7
JFZKDvcMaI4JGsZLX3RG/Jxa6MFz1CUK6DpgEQnPHtu6IgZYvlS9Aa2wopFT8YNyWx/5e+862ow6
Grltd96UQrNVnPBZ1vUnT1b8dzii1sXA5KQos9VGnpSO07xyOhqksUvCYUTo74/UdbRFF5Wm1vC3
dlaaqDD9ZeUunxaic1c5rqifIK/jZ8tIeUVRmCXaLkLgBMe9JhEVb+nXuZArEMtwdVfD1vCVDM8E
q+xdGSyQPHr9bSfXxMwx6Cp1ooqY3NPhQdtmfCGFPYwEMwJAWyWEDbtJ2Vrlu3v4PET1SPUmlJ28
YSJPNowsxFNCXtXiC8lMQGZyWSZbrkKSlZdHc9rwBZghlszRQR6B7HSSDFwZ3/Nx+q9R2iLHU5WV
9ESkbKFYtEHJ19e1v5ulkuXhJapyH5J5lPKYP3OKqJiPN/zQZTlXSovD+i9oqV9iWjZv/1rn6Jfa
tkCv1Wo1PVjnhMjYPJrNEtfOVZadhG0lQrG0ZYFD8Cpzec3kEmdZ8odXEr+W8Fd6G04eaBZuvVYH
y/INmGMmvu+kvqmI0Q0qS9tZ99xpT9BXZgDjYv4s82fsUKokF79PhX1Dp8TJFvxpI2vBan8gXsrR
wTQ0XLy+LZALK/+5JuC8dn5kNMqgyYqxxKdtY3iySAq1FPWmcbU1djM8iDSwEJ98pp1Yjf+bhjTo
r/1j3fKrYwEh0MW8sFQZM3D7STgSSZW+k+xxQNQUzreO+AxIGj+u3xVpyW407NO6/i/CNj5LK+RR
VfvabGLVSAig7TiO5odaFSwZUgrfhSuUOL8hZJ5hwlvE5JujxbJbE3aTI6Rv1Q10phHMupgs85XB
gAVwtcWJfywZHYLiai7YfwLjT8ubueEcmKyMiYfuRMzskoUq0kPuX/WcE6sg7OIcRKddhPYOCtlc
e9zenev8go5wJSBed54qcNuXuissLd/i+9wNiQw6IquhOLWEGJauhzQbiYhQeiRzEG826DW87pT2
PSk5g6QE/jqNuVvpFLy/RKKywujxtYfWdYt2feswn6bSjjXq7SVRlfxc+xbaI+DeQe7iW82SHb9y
3uTWM3X4aMjjaCtimTeHwTBTB8S4DLBanJ1NoTrMWN6eVOIXw7UdAVtC3FdLeXn5SeT59LtES/1r
ZOpEJHm6chif6VAQXZTIUWPYl6BLVUapnv33x7COBHMvlXTJBpEmuNRs3otnFxCdiRnpYr9mRxHJ
OtVhoUqQKvJfUHOK2QLkvWFq7qaZ+/nnTLZJXPVEOFxH9eeXDyhuWvQ+4owqbugHGy7ddLAdAdih
b+iG8HLsg8XG5hMfGzSAEqWsAYZWAeEf/D3oGlSrYoM0CbFUQM7o58T9rM3FIdWckAAMweICPAo6
0eTCy5u/pSJHvz2eLQEVcphdiAUBnyznfrQWiVr4YIuPQDro8cfMEHzFq1KhOoddCzRvXXOoYPDM
0tSXfn5rnke405aynq3BQI06N1HpX8Bqi6RD4Ygg92z3cMg+A0zMibNohckgxU7F6DTk7gDFxy40
1bn+2UDojtlQDWWM+OcwTezCcUp67elEuI+3dq4VcVxeYPhiDUsJhOfYRFYfD6/Ri4oMOJmOrnjM
vFkwDSvUcKoZmM2oDkIplljPnevuySaB5gD2daAEslvVludM9P8vn3pPYXaJVO1S2DfKfYxJPh2n
5TBakPvY4TYrz2XD58nUZyeURRgnO+8cQdI5hr6H++bWOKrSmNnoGRP2j4YXYg81FcAk/Ej48sAV
QHgqdNWRg4Lqspyl89Y75qDzqoVENbpBQRONzaQgKg3PQh4eBL1HlOALmNVJN79iTtuEyWki451x
o01+3XGHeSltlZWLwR6LrRjJPi166tY7Wr2b2/2JqaPR+QhrmS2zHQUgLyGl6WyGjvd4z3rUjDB9
FidA28dZBgvZAbtY8utM4xkXH9nPLXooFIZm2AxC8bAh/L3+VOWCvJ7s+S2q/Ue6/TygnAFdDRQn
GiEauYfrGx2smYR1ufYxvNysju5BvIejTG+vwnBJelobnSxhrdZ2RzkEJLifFwwFpiMzrHeuEknl
LQAtQkwyNbGU4cvUvhx2gnfEzHQzuoxQD9TFbM6IIIcjB9IzVe1y9C/abd4PdTZIzDowR/IEyzQv
kNInGhKAHjQCVzZqjFqPHHW5RECYXOooq0FJGb97fqr4SnQnSAe6ILsAJFhM7HZq8Fi20JlAq6BR
QYJ2cx6hQwugHJXww9gOBbhqdnQy99araFGMcW2hah2Lmx8WJT2hdSb47zLzwm5ri9fDApVu3YiT
d/jq1QfmGHQhkZ1b9vP5vgTYxFZSaOjXF2H4Y6yZoQ013aH1cNErVVuV62fpAmh+HIyc5sdAvjbB
Mmsk98hwciNsWv6luE6IdkuUFxinAW3Wh1EEkRGHP++1urunYosleytRxF87XsbRR+eMHxfmVf2k
xwPuTTfckxuCHvRqnZhvzS0MxEqx6uv1HTaJ9ODezO1CceQzE7+lK3gD1p/wKYGvensY114w3AAO
tGNjKfhidTZo7wNgor8em5IQGldM+OjvujXnCewkZdCHiZI/4TxSSeCwxuTSgPd6AEfpqgyqRB5k
8zl84cm4AJWyn8OxQlrpwLhI9N1hJFuRsho+LU1ARuyuc2ZFa4D3mFWvIVi9flVHzGB7gmPfhfHZ
Dexo2diKhdgoyymxlE/waCQn/uZtBcZUebvI5pnmaKeQTPIxAutlWSn8i+3sZ8I4IiKFpd4e/i45
B1/G4ey90/HAurnbh5k66cb00BYLhAQV7ej9RnyHHZKLGih9LoPrP2NzwrK5kCWnlaWhKvvpTTsn
caA2yLB6mWjduJvfPL+84FQnNPCm9R7a3R0v1OFoy8HrN8Ulv+ymTQWyqHnDT7yEV3/YJhzokdM8
ztSpvqHkPwyBPq2YOzLQLiXJm+QVsRBMhNstSP81p5ifrcQVgJZqum1CDTjziSfnPbPM6hSC6uff
Q5r5qbzFmTyOhG7YQik8f1Iuq9QrhPlFiX4Oax+LW/h6QSW4eZScx0fJeC/TLl/VYbij5zdg7B2J
jW/NNtGfftQiumt84Vjmi1rlUVX5n5dimBviizi6Z+Fg6CWbTOlLuRQ04jMIsCLNtat6eoTfs6DY
LFqKvvJ7ehXIgylkKquD7UorlCUGnnEyK5JQoE61UI7BwGDdt4yKzORXk51o1yCx0Su2yQY0/Ozm
hupXWVSMMJ8ocS3w4o3BRaE66kuN9S3eTGh4I3OvViFKry5hIbSjpMFyoLwxRby5NaTerJg4FZCT
6Xu3r+OvGiRAAAa3KA93oQSXr7bKLfjWE7ciPfRzmeVu7MofulIXCIvO4+nnh1RzyNgsnaDFo3cY
mAboYNGCJAhhJtW7m+ojJl+OUTkQxJRKD5B0QVVQElIlrL6cVkkUibOTnKMEj7P8Tbs0o+ml+BBe
5sYo9E2C23ZtPgAYLVBIfnttc5iqGFa9EJspm9YDmls82unVYOXEV13KEFpZZhD89sWd2P2AINxT
xBTItTWWvm5R2qWg9Wuq1mLN8xOsAGatVbZ8eQMEFpwU+V1n//Eqc3RJGcPhWffEbxoJewyPQrG8
o6yA53SCmtJrxpH/jhBeZTe+x74mtvChNllkvtG2OfPxW7W79OZ1r9vTvyZ5hOpW/yHhskjuloBM
hs88RZcLacBWwX5iMxc+gCEBrfXca2XMMSAEk//k7hoK3F2KKNPXGbD23+oaf7Al201Lw8VpXo3W
TT6BI0VHGpEIEBAQRAuillERk1ieTARWuc4IOHF0Uf9NJ9DPVKf73FpA/aB2DWSy29Yd+PcihO0r
qZFCklG4PG42YBnZfewDnNfMgtCRNDrQJASScbYYbF9Yrk0uBXuUEiBz7uUE4su/n6BY1R3+ME4L
DpfNJTXajZYvOxtbW1eV70eJlST945T8QoI6k+V2GpCuvYbnHX0zJfVWodC1d2jWlqNFEEqTtBwD
dalyUjo83dDcYNRP55UGoewu/qb5cCVHkJhO3D9cpT03gYbbxZiqk/YLHUUjIbyoakFO3BvobjiK
h78dDtJduothUJ3UqvYQutCZy6PZdluxxjJQfHShmQmqTDMdPyum0ca2HpuxY2ZTlOJKcwWrPAjG
8y40vNRiaAL3flLXKFnSm+DTT/ofUpc3QOy8QS/MO7+kpXemLEduRRJEyKAAGHBiK6Cf1MT85trl
uwa/42D5oyON3iBjJ4UN4jKeBsFLNr5ZHzWNNZCPEfTPYg0kG7QaMler36Ql3V5aSudXmyQu9OWg
C8TOWlkzeXwIIIpYm1BMOl76+mibB0qbapvMTu+sioF85FbykkY+z/SHaKytcL9LHWmLI3puXTUs
ZGyJwE44naddw+lv74mn6l6NjT/KAjy7pBXdtAwyXCLAFUPs2GMQvZcqCUHTmevA+i2fQjWNWkcn
1ThVZgEDmJ11/o3q4wZDlachLJel+eDSO17nYCB1rmJcxYuEjfjo3e/oAj5LinjMZY2EMnN017fp
dTUjuiEQx8zDGup1ozeJ776TPlVagxjKhlplMyNP9B4sDJLFQ/I+oZxUB+kGSAp89/ohqTe+1ank
ADpBjtFSw4qOdj1vvtvOB2FgsV3TxKvAzgtgAWShgcVxaB0y6DuOMhUC8ozbyVcBhBceoX30wjKg
V/QefM7LzUU65uPt5ppSxJL9ez04KkzzWbOALH9I+Ru5PWSM/gH26B8JNlRyYQetBcAfQTFOkwjA
Np/UTOxWcRyi8NNIRwEyxph/tGE5F4iTiu3luDpiiTNp5mWUjmEDmGM5eyRUWw4haSy7IdMgpgSa
xEEX0XSfslAdk9/+BnQnY8JlI/l2alSftSEDm++wLM/a2Zd5nOJr95dPtsNHBhY/EyDB5TmPJ4ir
mSUv+1b3y/T32EuhpESyIYkzT5AynRImUQoE3DYB4SQtRz1sRZSfChw3z5QBjRtjiChBiQx2Rax5
vL9/eTgHyT8BZf5JqUY8KWZquZnooUZNuauB80JV4bEHjiZDFD3WcfSzUrjx8OsWAhsFYnfVsZee
QbZrEDo2+58sIZBdcD89vcB4qyLHyF7OuX5h01GKgvh3JpaJJA5RWtWo0xVCLCXTQSlGrwA87VKi
RIhBbruUBbaFH6xi/VlQymicjCTDEU2pe1tJ/IxG7JMZbKMt6VvgbZeflzoM+wbNHQRJ9T7xAmmk
pE2Qqtp6xk4bTdARygJYlhvdarRONIUshCM2GZXqSxCeSyNnxe1VZSaf01GlaUvCpYpeawgntrY0
nYoBNzMxhCNoFSxgEJvwdgstnsgNeJjhYDDswepmMFZeEsVx6vTHYwVwNPUKyhC09k1eXNrQfM2W
EGZsWxS4kq2IrU4nEhMdwyCyYyou78VR+u42M4n1XjRD1ItBhlJXLuj5BeMUmP+x94zeofzT/md8
3EvMvPxUSOYdPSkLCYXE4bmpsABW7AG36lKa19bEW+bUPj+Vv9L+WZZgy+lHLQWZsFJI78HPEuES
k7KOPL920ErCERtn2Myt6WjwvO4SUvrD7XZP9/F9yPFFbERAHSx4QnsZqM8ot9+7PxdkyvAdwrGI
N+r/Gaa8BsqflZhgi+1yDAkosDU8IZlynPed6kHPl6jMdLp4emD/aalvMHW/1Zg4WPtmRl9gV2GS
NKx+b5Rne6HFra9E22Zle8aVYhVph2IGuBG4B9byG7GZ/PzeeuEML4b/ZV4XBcB0kd6uLaHjj7ar
17PGGfsB7ZXjm3s78nZcAVPrBrFvcIQSIqtgBOyEt4ecN7qXcAEKolWzzslhkZjU15TFb4tfD/zj
uWBujIyzmg8jmd0Ucw1GKniiKKkj6uySiooBux8qsyzRUzCjFbWcWF0nDnnkHlwc3WOebLQSA+NA
mHMRW9xLPq1pk5uc4/N59StRs2LaJQ6UfCJmHQmTYHGsnq28v6OH8R3GhOyiuY0V/Y+KmHZa5isf
qWZEXNgQWne57eE5KV3joc0vVSrpKwURukiiZ6xp8n/AF5K5cqjtbr4CCteQsx9unwN67QJ5lM7e
6dE/LhB9lXzkJuAWOzInd2xWumf45rbRVEBWmknDUCGDrKMizug0HVCYI0XBnQ/mACNXsw1oZ9z3
P2vr3phFnCXtge757YTS6nYTlGQXfaTAB57Z2QqPO6n4Rhg8YK5nxeB1LnWz5g7tst1jEY/3r+1B
4673V0ixL4yi26b8NWJxqMek2xsHMsiDztxdamn71oWfvQtxIGfKS3W3hOuo34MjyNGNSXUAwDCI
vTgYVEptmfxwWcvm40swikVCSoXJiSH2sWMmFhyI6ZhQVLSePp5B8+Rn8t29L/ZuKsIWX0xZW/rl
OIaSLgB4C/XOUeEv0yIbo7CUTmQyVyNNU474ZXq4XLyYQqasqQwHBjqUwvGsVVsm169N/xDIZw8p
AlYnH/f6sFPkYwFLQNWwTBRqkqC2UQvio0EhBnibFHTUOYdqi6uMORy/x8r4tXglW7v1dU0ub/Zt
xTbCCPXeM3fJaBS5y4tmBlrKLWlQUsZ27PEYNx+97m0Gxro6vFUE5G4DNcEne7EpduoAE4j2ighx
3z0IGoXgJ8zaE0y/XDSGZ12o5agi+AOHBkmZ5XxvV8DWh7GHvkfblMsqRYGl7Xa6JB7+CbA98/M/
ulsp24ppVyFr4njvuPc6T/UnoeUh1/kTKUqqNPZgkhknsTDBVujLpzuPxU08oRdQhYZTljhy3gs+
DM1rcFf2tQus0C8tssbwwi7LRj8ofKYIQzB34FsKqo94VRPJpir89LojBOT6727+YCt1YD2tGDZX
Cp4Ifirt538ra1oT9U+hw9uTjouCbF3aTsj5YQPVzv+RnfrgHr1lf3P4bC4jZyOIkAb5xwm9qgwl
ea3Knu2d9EWV3diLpDMCZ0l2Zhh7W96dtV1F2STZJNCpNtRBotO9vfqjmWJ/eCIIvDoKse4VxEve
gCizhJO6hh7fVZeqo4yjZz/0QnaK5wzQeKtXiZXqw2nXlB71txQtsiyExcP0Fj+tNaH+EbfI6wcU
cjCn2pPHJNsJ0bds5LqQVgwHJMR1CQohTq0mZQro5FwVRweytoHZ3IJ++nwmdzNLdxmoA4u0vQLI
6LOkXae+Y/g7YpsT1c7L6JtzVvkGWHqZ58PJXQKoC/xkrtszEllNJ8FsaUbG/mzZkIJTc17yPpI8
klMM7tvymgY+jqLBb6iQ2ODOLna7v6Z+da7ZC/zR5gK2uSe69gME478Coo1ZYt/53pQjQUz8C4Ag
V3UPgFVlJEGzavG4pZ6/EdNaO7uX5ECXeMclg/iBqS+DosVVvqrmopB3gfO6ocBmO1lgahU0RGnt
QfF5QvRRxRfzzsq0c6fmdKiEBfUoDBjGcs0cdIjWb98VZmuvVlQrD6O3NZTqgwXoeziXt9gvoPbK
L9XbQW3QOPBXLZRy3Ysb2q+XdZmanXd6pGpOIUExk6VMU26X/t7ppHpiW/i5UFiQdFGMrbsWHJoq
T7Kx6XrvDKbYDKoR03soZuWmV2NexdtfJ0U+4dBkuPY4fir12nDhMDyt5nQf6UoXtb0HWFOA6ijN
3arpcgUmQl5/Cfe/cPIQhVawH3rE1e92fr7Lp20qf1qTauGPNLPw7hkxCa/k1l8bculXHiHvWdGN
r/WSllGt9V9StJnjl5LeuH6kVD77Q1fj3i/zF/8K8GYww7WgDod9I28yxO9ZLuXcTiYamHZDjskr
eqL2TQPI5db8Ux3OQ4VwV0YYG7k3QLZpxAZjyS9VCiSd9on6i4EY5YyF15yZuANxLQ3DVF6qG3L1
lHj5ve7w74U/aOGdMJDPyCETlXzETk9EXYTn5nSXzvdleXkO5/ASQrhGRSi4/stRxVmPTgIx7XO3
vhGY+XbN6BCqEyRg4oPPdmbblknvp5nDTWHXQTiD3EKfOQniR3f7NJml6qXQoVwRRkl0b/9lgCEQ
h/W3iGfPj5tlTf/j2mtw27kQ2n1hMOr7NwdqvWfBZTfqqjFHgeoeq7IDlqsqadPH56aYm1G7KBYA
Uf10iA59PdtgEVPBM2YCNyyH/WIK/h5Ig4yupsA1JRxCBfFsvSSf4lVObJVYoZhI7k43D5AnNMX2
oDT191zD0MEcUNK5U7yf6cOMVOARZEBhJCo68VwzKgZyxaIguOcEorfdD4W9jrpjZkr0nod5arSI
21V0RUkioiLPa/zekxsgFhiDwjawwv0+RC8V+fKk4/kNbPYMRoVyrJQd0PJ1DAAI878LcOKFQdH5
1TbeCX6uF2zUT4Ht2D1yUzJHx03FrgMGyE+ebq6+RQJP7kUf2i9BHZj9By/LYNQ/4UBZpetFkHuh
nCb4CkWN9JO6eGtQL34R8Z3Gk69xB9S9QQOfPuhhp7kVxYqBwNYwo0HIsLE7SlDwSsAM4n5RNA94
m6hvdF8YAzdNO44lNcbGAHvqmU++RRKAESs5IYtrjhdQDlpfOZTeuEIOSY4J/qThn7zM3CoX5ONI
sDXzyDk7psunm4q50go+Ekt8/fgB2QTPqis9zqTdTV4XhYl68MAi6vaPkexsySe0T/23K61PNeZI
hRt1EnzMh+2UuGozsHi2wlDAWl4DGowpB3V9Ymfccc1u8yZec8GWRc3UG4lUYg4hFQOl9JcUrA/l
v+DzA+kvSOnpvdhAxeajtb5WKMhuCbsTPHb3dE4rXpXJD5ffqNWN6x6jHAbE5LpRn8G3znJDRYV9
T1MzIPisd8wqCXxWSwUqO25gwHcvHFFpUVxR7PkDNr/pRCHQWJtAnimF6TVNGaPSvhVyJ0871ibs
zeSJlYRLIsH1JNy1YXPhPkgEBOkorop/CEHk8/vjhoFqN9SB0LGYQcbpZwbDKSQTykC3KQr9kkrL
am1X8xvSrbifARWoZQaJYMRTahNHmOrgKAo/o+R81CDxW4Ts+K8A6B0NnvAmnqZox/FYwNnsbU/0
HS7tBjYCVvPCN13yllqi2FpcBXG027EeqkXBFWExDyT6P8/AgluPuipDFTvzrB2ppn3k8jaK+9oi
ouqKk7/aIl1Z6QPdpEXDSnVfP51V6VOIprPwpG5Fumli74xQ3QvU7tjszGdazMgQp1OEqQgyv0Xg
rJPqY1h1EPQ9oY+QMCFjAXkQA/JBwpDQhCiSvSbRf4Pr/ny3itogBrMjGQ+Go6GW2nneHIbjiOJi
MFLSGNSyJxHl56wv4PRcRT25M3dkFZLa8adEKrN7WUyilagEl0/M8MM8ypTVaI5Io+tsmdf60CoG
UrMEpmfEelGW/mvGqJCt2E6FnvFPLsNi2ILYGXOfsh8VMbW+INlwDKcNz9wGizrxHUlPknT4k+Xh
qcQ8co2xTHBWI83wHN6/AGKcArfuIrJIl4jKWFW310SzswfqRMuKhimwumG+IWI2USpyTuK+N3lO
LAaGRgj/hqgBsjjWrF+ZAN1yI5u0X+AFUh6l2qI2bgmlRvxcGkQ/bV6eFr521f7V/2TbkZcJ4b/W
YIOuqmWpzQKPYvtL5V33n6MTDbSotbMw8ZZ1gzqDQoGMPUuB5yWfZSsH5nDPYtorayrFolIBKohY
XICH+1DqdPZMITtOthJwAUoFI4yZ6VXqg11iinSXD831gpGn4aruK5HYqixa5N3GtxNHVuU+RPOc
frVVF+0oZf2fF59nOKsEw3xnsX0GOlyIGleyW6KlW84nUJVUaF0GlA07nrl99n2H8UTfF2ZEco4L
L2i3Me1BJJGPcvnnOW3HqtrFsf/2K5v9fKT0F/tvTQW0MO4BCvs9hsUXhsfzDg0KGgvm7U9FfNmL
4tqD/byu8Pu12vq5NCCbvdkGiOyWqB703itCBlFJBJtWw/Lu27X3I1gb6FSN1wupFDuQlqA3E/8o
28HSQYtBvdmHQD+AI5C3doA5x4ssQXQacSUuetAvDgrsjltWNz5EBLELXBP5EjM+B3QrTIjXnOoX
NVrGe2LDln4qMZk2JMvpAar1vqI0BfO94RGKKfg8MT4L4ZPAcjqOWlpCognewnJHS5ATZ6VrmGTA
S/wxaqkps5mC/lSGdMkh7RUEjq2FcY4urXg52OfuXALi+3PDgE864bsdRwFgJBrQM0B5CGuWpzHI
HRnAPp2yThy0M3Gicw0pqT1qRQ52Pzt6FdnWk0UAHbdGhbzzVaG6UHXLDIKDefjp5IWXsGc7OBDv
cDqN1wu38L6IrC6CrQD+CjmEdFKH9bDgKNbHswm9XHyOXD70UjXG/vVBYjbrYtaa3FnFTbRpzUtA
FLsjxQrDr6vXCCkVTY63b1c27ZXvPaaBwKttYOVFivN2VBLX+zKGpX6U1U40EE5zcbItAaUwr/ky
3CZ5FtS95Lxm12Uv8oalwoaL6LxpvTIiz1v6GuQ3EqEvutqABRgp1RLgIXpKLgZkPCxDhe8LW+qD
VXBSvLYTdzZaZHJlDoyfQPBPNcWRtw9vwmFMmec7RS88/VsAvYkwZh9xsyZtNuxdg0FbQvhW2MK+
SVal8TnrgzUbBtga7bP9plaFUfmTaV2mwXTDkZ/LH6hpVE9ym9GPboN7D+Wt1Ocft4URvFoWdHWq
qZy7vvYznLvkGOWSIUZMEIr/Jk2VSbJzeJfbHTKQDL/kx2XLJjZNxlmEeAJjez82cvTqwW17SWqf
jtGRInDOtD7X3P5V1jJlfAglkKsfycwDhIxGmrRIDJKAP4v1DZkjFl3XbOjbcAcLQkSfiaJukOuC
icCYyWsAfK58TGbB2WH6yWLw534Is7tr6I6x/DyRRvb84GNRLksAS+pbG2mrlhKWCUhmChDuJsLS
2pdlv0rqzpMqHCFm6B/m0M12rJOEQXdgfhFeW4/RvMRmz6ukS3VjRrb4RbyPG/GQKyxAMPZrjqfY
SwcFf7wcOXAV8hELBnBDsd5UREymA/nhllBiWOqYcwpw4Cj1q3sb88ZMsAImyX9aR5Imzl65eVUH
7L+rc3RdLMxl+25Ym+ipvqu6MwO/K/80wvBR7r35ayDxQBPo1jwxwLrITloALf+bFLcEyo4RC/82
T+F0CLL3lqV4j4wrUY9wZ5SP1Ahnj2MnVjVeG0GkX27dJtwRCThRku3vZG9yKF0glTMCL+yoW9S9
KHjJodydSjRvywZZ/epXjpkBEc5INU6qHDACuFQ3GdXzCotk0iEl0ReRhFgb69MNsU+BukA2kkO8
LLoN6UplcVJ4NT3oWIZCIgGjSExBZfNwRx6Cm7L99BHKelp7ObG6b0y7ZA5FwGKWWwlxJEFg7EO/
7n1/7nFpZmjoBArnJw26+XzLZjdnafRrJ4bbNUkCgYIMnGb3yCNPbirSMQKUqgRN9Lp7ioFxBRNG
CDCa/QuV8DuDVmxoyjkPZhug6evJY4qT9frT5gMZCxdyX22mvlICG1mySp7Mc5ekfzCJilLh8ImT
lFvaYuyxE6ns6vp6nq4Lgg5NrmC7fZtYdfd0zVG8wutNN0XtlcBx9SqLbNaW9lSSLhsd2DCIMClN
zioz4cY27WQV4eN12XcM8qpfIY/grQinEpLx98SqN4/vzGc722UbwzkEoutazweq7/yAosjSbni2
R3qfsvsXYrQ/2iYj/OLaWDEaWy6Y5IGhg2rDXGzGfbj/qHYRNWe2vTDz5qU39z9PIDS+tlK1d6Vk
8CajdJrbhH/BCCgEjIHwpragS3IGponIsI0ycTl7O58z8yZZIghxhRTmHts30VfMoQCTAZn5lV1D
9CbV5PrDxXfI4+ogws9UPWzydu8YVqlCr+McaF2GWrPhmJbwDDxpdQ8hjVUcCcvjoCmTKXDB1MHg
OZsxEmtLFqtWwEcCw6/D1z+66Z2ULGwcdqthltZmliUv8V/7Pp+ChTlxh4XLIr8HmB5u/qGei6hX
eFhEHqUwKjkkmRp+6DAWNAhz19BX7if/rAzl5CcgxpQPGWpIEGVruXAgbwQL1f5gnzGz7IwmF+sA
CNDg7JV80JJ79WWyWPfDgfQsw+cxqHw0BWa7Y/9Ttor0mMX/IUVViEFul3mXWNfMJ9GVLXcFuPQS
jSt6feNUgqcpwOs4ouSwEyU2+9D/9XRHxvwuhOt2CDvhNqNM6+duc62WZIgB4Bw//hagn1CPVUGy
SURxvgTxmVPkQJOuNin2SjdZu/JQz4o8SJgm3MF2DZNRnoMysPX53+lE0uOVE6v8WtDab/qoVdtZ
29+qCa1yUqoHtVecdjCtpSYEmtGv7oorHJEHj59+F6RaBqzhQqU2OJ0pxAwFtd76hroj3H4sXc/B
SncHGYMjY4M2VZl+WOkPnAzt/w5SxvxSxHHtB50d/uxyaSVQQM20PGbz9n+UpjNPunWJTq3mL1Nx
Hr9NkaJAdA7QMPwqXffXSoalx0bVRGF9kI4m7gUcSQVTHn08p5pdMvtZpzngI8A9YtcOuwqlBJCM
AGmV/7qkNzoG2LQtD5daAzRZhe45fabbSvrwIMoNnHBxQPoILmvd/hD3bGTpomnFWzk/kSoEFgvG
kTzfrtAQd6V6dk73ew9t4m6FN929pI6fqN+dqCvQJ8Vb+r6S784vBFYs58fJ9NoidHM9IM2KXq7f
MiOVMfMd5CZM3tu2OLzVBL9RHBAwD/GycbqnFr27aHNfvqAhRanc/GpMVzzF/oq/oxnnEG4acz1Z
uFWyNw6v0Btlu0K2OR0rDRhjoKe4B76JFw4N5qSp4o+sr+Ctudfc2r6xkH+V6YfMOqmrOapd9WhB
1+qdzeeeNRSGJEt7XI7M79HKq7azoTOCiNTJA1gfdhd+bmM07vGiPD/CNjQmL1OHu8moKrW0/NIW
DS+lS/CdjuCcyol+Og5XFtEeZybvRsB4suAQGbb7hwmGNmRbNjq/DQw7EwtQWzxkFHx7l6eivAWu
Fkr4U0RxHkNqR+Y5CpZXfLsVbt9CSAv5L2ZEIeQg6Vye+enIE3RF9KMbUJ31Lo44UP3Ql8S2SKtx
f96mgggW6CeUFgggL4Ss2gHJbxSa1HVTHnnj5QXHaVQUoRC7zcssJUKdQT+aNlejunsDZtEWX8r+
fha1bT8j+BNx3XxxHMhqxaqlY53/7tUeaHU2akDtLme2aaRwvmvI1aLpWkb8VROdfqKsbtVVmY/B
P70ebt/f5qQ3nYMR3IfSoxYohTvRR/GP4d/hgl9B2KC/QQs1l1NnVqacspTVH39AjH28ZFfqnXrL
w3XCYR00tRz0LkMXn8WMc2Su+q21IFcGbYTMO769hohkNOjeCTAfXRmnjX8yJQeaTU+KcHXw5DDs
zNKPqDJ/7gTYSFu0WAoLgbZBtyzHoAdSgeAgKoEGRWYown9yachpqvPfFBX9vPLC3HMiXDgQ0H0i
9RvVOfin9RTer1SJ+CuEAjNxyQWQnn6ksEmi7sTv81L4FjQUlf7MpCBnZjvZNklCvezhddxACtOX
B5aHL9S7SunTx3Imq1gS3i6U7OfJ9rrRSqk7tU+rjoh3/3WIZP4b2QN4npiswvkrjogbZp8SwHZ3
yoAO/fB9ORT/0Td3fnWYFPvN/wlB9izqcVyKpytzu6WmN4/jpXqANuPp7277xZhai40IJ+sT3oyn
+kULQ13tlFqA5XsndBW+5XJDg7yuXeQLEcuKdpGGlvOmflUORDCynOHfuHOa2DdCWjBOs95CrCbS
wgtjSD4dGvYjEz9ziAe0GIcsO9ekzfhZ0c5SZ9iZ9r2qaBjv+O4GgzAtaV1Bj7kvMmB5vP9B3H31
3AvftKTvqNw+4aAZfO300mjEADSksE0Qf6Aivz6wi+lFh2QIIvPRIN/wjp4nS5DFy31xHwcRTf0r
+u2LEJlV4xo3HcXRlOd9Xq7/enwByVwGXQ86vqQn9JGD76Y6NlNXXIT7+dV8o+7hmivOhLSPP2tf
Blb4IZqMqA6ISI7kET5CM+bkhTMkwTiTLAM6sFpVbi3LFqs2sN+yUSPujrbpozm0ZT2gPeVBuQtL
jkCvvjrandJ+vBHtgu8USXnY+YCS1hTFS4Kr63Gwy0qoUCI67dqP3YEc0Jx1uAMW1L7TTralYHTR
3PYsFQWauAwUcaPdSsmjIgMyKOm2R3Lk8qY+Clr4llE3EFFfdppLCPRgS5soNrmtjubCSe0MivG1
qsqAHCrVSUW1CCulFSn+p7f1OeRPb+J/BCYvk5Yv/ItO848EODrIHS2p8KT1oFZwjiOplNpJMMEo
+lxIjLrKt0HBC33N7wQ+WBdoAaqFzeH8d5YV8c+t4qjFwl40+weQyah2Pq9IA2UpDO6KpoRtKYVJ
5DiYSzCchyzG9Ixs182zh9pIAINPgxDmO9qlYsxyUy12oohJJo+wgOnH3ka/5d3aBQsO6NS60pbg
tnxndHAAMp9Uu7MBCwq59/u1V5aLvjxDstN4LkxMtoKK0yRhKKV4YKrDS97CzK+UQp7wESj5dtk+
VbkQOkdnmhKeC6g97r4UhQtxCzfmZlqwbln1eQDJxOSeo9RUKdrKE7ASH1ZpYOrAnWVbLWiui0/R
50wiWi5+Nhy0LyAx5yKH6xFomSwfWH+VrH5Cf8xBzl3//Xl/jfmEsDMYzkom42MwEp2IuCDhrUc8
R8SJ66mDgDELr0cXA+ceH0L2y+9rUhxow7GgalkXY2JCTM5WZ208svGDZ9xRJU+9SrEHNW+QRwQG
VfnCvEbrp2niUd4ywtF63Bj0gByBSPuSiigNtWEWIBl8Ad3O1doAtUwbQ3khUWVjsxJZ8dNvJtDC
Pa1c9xp7OMD1SwNBHRFKgiYfEMMWiW1AqxzBXjiLB1VxGoIeSfP8WVDy30WGsVQtwEa9Fvo8T/Dg
8O9hSnJCG5Qu4prm/8tqLeiW2PkBVKnqoy1GfcqoxXDjCgdxqua1GvnaqWy/SNoSZ7Z72FwW6Aez
l7LaKHIA/I7l4dz7qvAOmkQCF8Ws2ss64ZEs9Ftl4/k5diyWVGTJVJvr0b8NPjWooAUqxfdTWXTa
wRxyiqO5Z58lFVlnrptAeMoBk8pdwhz8wtsNH1nUr5Yybt1gmXV71Hp90wDhyhs9OpA2e4pRrig1
IZa2HsIFotghBYE5ef6Fk4ISuOBE+B2cplP/PChmUb4mxdPYe/pfqL+7WQSha9gpCWiVBzW7K3cf
Sjm6v61oyX5tPIb7p8xqg+Uvka78bECCc1B40teGt+YhcXPYEdZsxmhXlvrNlmqYOmJVy1hAanI2
xIX0CxViX1II47IW029ENnSHn+GTGo46rYFrkOA596m5+YGeTnUwBaJZJA/bNpcP3cgiFC8bCeM7
SVmhhDtpCs1m4kBHgPme36aeSNz/+yT1fm8qZ6dZd1jL3ZmwLksapR4T+ONoIT4AHnnwNDrMF8os
cO3hSScAwqZcoH4J2sPdw4F4p5CukgDXuekt5QQkmCkMo3hXbWnRRdkk82d04db3ry+HBJVUfmsX
CGzs7W0xbsmRKY5VnnAyOgoqkbYIkwXeodszwKnWy9gH6MfhR4S1Fq9/eUkA9Sjn4Z6SH5jsGP1e
9T2grR9saTEzxz+cxrmW2p4WqglWLkLdMaolkO3cGxo+TCn+x1JZoueiU54T+iMwiMnIGeMpCce4
muHRu3WdXMeql3EXd0erFeKP15NUj/Quydbmthn9FKT9F9HetJG1jvo/M6x1+sn+a7lqS5Itf4ek
u9kEOe3azvEn2EHRqkJ8E7p/0MVaV1QXC47H8KeGZHbwK/uuQ1dAOuvhTib8qaYuWoTurYHf2I3Z
zN/jfxbpiZFsnda2Tfua0xT3/Ui9RjdU0AG3rzfO5BfPumRmlHk24mnfHGxVvMdfnHPf41RRpH4m
dG+ABKUQiltjSZZOn6E/OKMU7NM/DpWFis0gombv/rcnau2F7hN1rPlKdoujS1G3KVL54FUIIGj5
wijXvEa93zabc7hRUPB2v+GLHdryw3vDvJ150Lf8mJFGRQXsGkhxLJESYGMlAiDBtV4EvuS2ayyf
xJ9ehO0KRItBwVO3068KbxTY4ZDIuPKKc2CVdX9JFWqR0I8kMf7ot4Nu+GZMLaYYLqRZQdbNodzK
eS89ztI7F8beb1/wFJKe5F5UYzcsbAXY+lprqpOjtGL+3+lXr+J7c0xv7fnpH0i3bXEpt1LMZXqf
zsdw3pHkFQNG6VhBr57M5XYpNA8DWRTrHJCXrNiZropY7o+4CNByomKEdKfgCEpo86MS0XdEcAR1
6Eey33a7NISK1BCqDG+05zo91Ik40pqVxiSvhYUZ3eQw76ixFEz6EhMVRrXQ8+sh64UtdaQnRbSx
4BI47OYhyhrUTQtlh2WtgV7yFTZmMAyLoTirJLUbacxEwPyiHSzqC8vBAW23P3kWmRuwcaaTjGK9
/yBw48xQJftiNkwKq4wyPGGhMTCMeqdXhRUNsA9k7rYxQj4xZBILImna4Bq9IV5fdhG073GY+so5
n6JhjlJVIC9qjIiISorP2DZjCQWXJnVH6Cqy2CEFNWCOFik697MXn6QGA3VO0t4kNPLNcM+Iu+Xx
5hDqRABiZkHlz0RrkiqdacNw3lkp083/tl/BW3xnXlYPPuXM4ddrYjP+ifBfA5QRwWQG9Y/9Koqu
2XtuXMjuGB2tpF+jqwpVugDHlMnNrw6syVm8tyRjL+fw3JLBCmX5soET1nP7l6N3/Sgc8gfuaak4
a8h307VyVFDhjWr2SD62Fxs4VoK8FVyED/84Zsv5aESoR4UTjLPjyZpoKJy8xi2UqusktzaQj4+y
s6J1njJeeqcXooZa3z6aYG68a83fGYEBNQmtUMUv+6Q1xT4lMbDlf3etP/+0ELVK6FdBy77VJEPE
7h42xtBThZ84xSz4jjkIrf5VyixZ1pW/OfuNo0ONr4/P5WCkG/wi3L1Ms7lIwud3RxKvQD8egZWl
jPQ52FQ4ZNx1haUnzsAoE9UkiTLEllU6BxE/AOYMxTyLHqUdzwVQaqMYX8PxtRlXOaqfE1hhfVt5
jadYhAOU9Qnrd4EajXBHPReEZSSMayCb+2N/dSlCRVtSCw1gRFTjynzHPM1VKgKbAfulTnUm2Ikx
F6yS834RHvaXh5MX6tpQ4B1qiYXLPyKweT8IfR6I+jDiHZhrG2YAw1Hvxtdr9xHb8JDB2hDEGR8+
QQhh0DsvzM0mbfNKgBXBnb918Um6S6SEhEA8q76IGtz3aLrCsk+b96B95mwbRW/TIq2rwuC9lCfb
4gg4LaDTTbK6iavvWaKQNLOaOXJJyGqJEtDsAtpBam8wydulvTShhVkgA8dNB6rvfUKdzp70FPcQ
ofEpb1bJXAOYn/8QmGgOCidUErJEMwLL9FwS48c+uElbcDLk9jSZhTyFBR+41Z81KmEcloqgAniC
S6wmq0Q6b29oQCK/YvNVX7X5898G1TrYib/lNZl/eyIwaN3NSrcJx+4ZSwZ9tW0LzSHx8K0/WhR/
gVvur4NchvhYikYkBEVu9Z/7QKkVklsmHGe3Uk0CYvyvQfpCBbR4sQbq5BLprcqOlLxC0OO/CkVE
WkqJX7PFohCWKZzuCXlQGZv9FmKbNG4OVvNagJkswZ2YwiY54VO8ShAslC+GVHDyevFBelgcUkEb
8FJpUWDNRdYgLYwlL7q0qYiCy2T83TfNRK0j5u7gYtL3gzgHdnpSGp6RteF3jG9KJi5+KES3eNti
jBJKXrTTbUx0lu9oEVAblq/EAWMZU5JTg/sPp0c6AVYSVv0Yoh9IX13V5u6yiR4FX/PHGhp129VP
YkAGyNKSP2S04FWaekq/fNDdhEiSYc5EzxJbKk/kgH+7iB+pHEcY1wUha2hlf5COaGedPRXKScAw
gORnJwXGSwrJurJvnPp+W42zUGJfzDRMWkSMvVtdFXoqQKDrXRk1+MgWpow3xmXZI+KEoQXHqcP3
cDoJj3vkKruJuoBQPJUG/0gRW7691WzmpRh00sYSQv1fpCQ+t07xQgzXhwjatn8lJXsx6enLSqT3
tKMYC2CqFbOwfkX+w9JAXdtEbKPpeyJHqFPCEWE6tj6IkXO3eP7FQSc+Kl6QiFS6PUOI602ID3/Z
uZGbBnAwYhZ9IFt0Y8WMyVJuTSBfycWS5v1JSixqNSZ4pCRqjFpUelSLPwqlutbW+2VwNvttK/pE
IXtz3M3nT1v+8qiAESnFPMmM8REgzeBwDF0mYDW+LiqhpZUDo8ZswlrsA19v0Ba9WSFN3kYeOnZS
VcHWmVssUwKw41s7GR0AlJxr/6nee8KW2eg3OQpCm8LTPUGtrO6IeatdVHi8F0Z9djKUkZdSzZaq
5SVOVnllA+rzrLYoqfLSfyplBTSpapfAxmYaRkO1pRrS2a4GQ08bpLel7iNp3/0X8yNe2wsFyN71
V0UJHCtWgFlrcMNhIRIPK/tauqGFAUs1mzqIX5YZdcjWWZS+74hAUDt19uCTRIvcNdCe0/KOqUMH
o0R9GtQ/envmCjrgNbOGLRypnxP+f1XMuebaJ9BWhv7aW1RSeTqg2plU682IMKpZYVQ3tAvcwQbw
UVG+OmOZScddit1vgWq/rUdmjPPDXbDSnKvcTmO0lHvXTy5wMonglq1wgaCSIc6Vr7mkUD+IlpWN
nlmC/RBkE1WU4rUbDmjbJMuFrkIclZ8yTuzaohuTxRAyU1BSSGAIH2rRL+z24muVBrt9EXr4gc2E
L64CJLJuZOEmFlDs8489sbnbxoJvjARO8wR0R2vpEH61x9H5y2GrT3AY8W0xjU7P8RDbTMJdX9gt
SJ1NUicoBbaxqMHu0u8SXPRXqTpiumUkzhhWpgthYeqOSnHwh0cVytUDaScABALbs3EUhV/W0xOB
ccBcu8rJlX2HZNNtfz/tfelvDnqfO2S6wrnIhrm7Ef/JFcZ45q29X+Lz0GPfbe9i6wPhQRcg+jfd
Jp/mEdiPlqoZajxJWrKJkY4Zv5/z6d+hZJA5JMfob4vDxktLkIT9uaympuaz+3L0QH/9ADbxXajX
/vYC6v7WYtJY7HNUfpzHpaXt09o8dGfyNSNS0NoCThXkMrewHvoXNOr4XnN72fRkx4KLl2/qoj3e
Ze303ukYlnDu/tJD/mdmzJSkDo4TYSeorQbFactDKMO7jM63dyLZxXjVl8jvpqL47t9nctDsif4U
SIICxZ1NCd0iM8ycW0H+P8d4iPeRFTztMGwp9B97/hxZ1nKhtGdoKBrynpde4PvuK6rebUVeyNQD
nyWZtKkjXtapGLBFhl1GyTbuAI7cUQ8PAAGFL+KBsQ7IjXNwRRUrn7n/vfxoEuIC32KYoR1k7aFa
3NRShRhWJDSizm/x9tLyzdXdaHcXwvWXbIHKI4w+ttVEGOnZkT6QBwgtHaGintJtkvI5nGWkdHq7
VkVv8hPS/q1aRXegg7le0//5jthwYrSObeqM2yNlknxEAcy2hBWleFO4SltRietseVDnQ9OGKOo/
bb5uRlN6DEhN8ZBrndDNZp7R3HpGdwMuPCVYWjgOTFNl8OmIfrqz67+XNmigMthx1krjy0BMhMqe
dVIXT1MzlIr8wSEO0vk58OLiBQwPt1P+zckxXm+agha1irtt8v7XTmg/XzSjsVERt/ay6ZpRxiAp
b2ZoAYEHaWvZFYEtBuwWTlIt7E4Py7XwfaG0eBTRR2pRcSfTXcDKlnAiI5B5ENhGL/BCMp8s4+Yd
f++BPfBNowZssO11+oWchJAdZ8uMZE0cVIYDaovflpfixuQUn9Tfd3jMKGG8r+btC59l4qBFw4dJ
QAbNxEIxQEbqVZRk4RLAondnFn2t3Yqac8L9oWDKVzcM74S+klUx3thy7+xOnMK/6JXvxzqowSxL
/4MCM63lbiupfONENgaZzF4Jynn0djpP2UeW35hqRMaZ0iPj9FsTSLR2MC4x9bUietBuhHBP3Dpq
KoIcYGtMuHyrPoW/c8ZbYY/diTYJjPDxON/wG8ojFECgJI/DJJwXVAslOk5x3SIppU9FjqvcjupR
KopkNdKkyKNKWf9+ZZhvo4CTY30kZZPd9pdHMmJiaazJu1Gz9gV76sOpZsLZ6jBLiVcyI9CU7d+R
ozoRyqDYuPkskNHmcXt0UGZLspQfZy6oFjyG2CUTLFVll4gtQARdpTZh1r2nRiuqRyAnsAECnxt0
P9+MMvDpgXiNQyp3CK9mQUL//hSOia30rtlcrT2L174JfpVkBrqY2keq0scKQp1OlFclHW1zqENr
ixcyeaNhth1TCH9ovXWx2KB5zyNjtNy61Whw3/IXnZuie1TKKrQcl4KAhSqLmPECnO4P60qPv6HB
P/hp21jufts8MOKOOCxM44k4EGlm2v7sW+hHbSbNZ16R+fLzo7lgYGVJjeCmj/3kHq/PMx2WuW1M
CJa0hHxO0td31EJN/8Nkh1VjJIaV6XRiHADqGFXEl5lrq7lpVNG7ujfQfhRq4wSGCZRpXOXwXw6u
jEv39A1t4YxygEBCFDtYlGX+iqMVgOboC/H+f+TBm5IviFTE0HlQxMAYPHz0Ag+kBJh2P5tlP1sA
C02QiePhL2a02lQGiEbosKMH8TZuUoxC3rXKf0nOsJEhKx1j2nIlksYIanKg/f31EeIMybk5ztbJ
h11fRl7knN0dty4IEUTMrdXWGpAI+AiKYwsIUcBGVc43q/qfugWsl1P5AhGQTeVC476kMq8Yi/kr
uCwinwarsT3oc5uycWZH6oCnEzsPkQFq+ar5jh/3TC2hOBMEj6z1aUaMdGn4SyP2a/bUMe3Wx5T8
Jyt7SiY1O0/HZXUyPPmkL0OkBz8K4YAWVmGkl8ARW2lngGgg+iYs95IhC23rsiyQWQ0HunktRgdy
jcUqUypLiV7FzTy3P/FMiCWwb1egvPmXFuMi2BOW7Y1DG2JROedNnc7yhqTaBerjl9Y/Dy7QLu3m
/2/GUN/7fpHbNyC1c0YkRs5mnLfylIdVoCEAAlrwQ34wkPRa33rRniwkJPPD5HPn5P05ys3+jIr4
zdK8Wff4l73K8ao94//qFTd+mtMaUlHGmlTiqfidQ1RvQS5BOse0UlOo6UOYtpUEbU3kYD81DXiF
y9cJKFDfQfNZeqo1rmDUE7CHccZXsm20VVdSSZt0pZ5T9VGR712+nI380hCccA8qtmYrmBIvZ5ch
qArvsEnNaBBeWQB7xgYfQsGoWtHEf2iGquLdx/5C5EGfCF5PXXvJcXMUxKVttA058RwG3ktzFoqk
d+jj8trxViA6OnwpgBcPqTv43aXvCy8fFg17cDxdTl3ik8IhIaJXH4zSiIKduZOS7E7mwmknFy/q
oQG1Ij6vICGvuZKbI1JrLz4eXewSlsi+PF16rtCiuuZGvIcy8oxJsPMeN+9wcp9Ysss5OKs5ikHy
IaUiKPdhAvK8s5ZJflnrExFM948oKco+0Owpt/jBz1gCX35Qba4U/dH/RTLQTDpvmTd4FsV3MjNp
buOC389h/PJLyDu5VV0hSHxFvsuf8y8eZnfa7F7vf/jwWT/g79wk5FLZNTtE5WlXHGDztvke5X04
xQL2JgUvMRZHRCnfdfGls6e8BH8QQetEf/vyHdlpn/tJCSSU6LPpEiY21axG8QXnL5rTv0NdvakB
/ohbzDGeaHVqXv35hHYPe4RRIY880AacADb8L+ayki4RdGHpepZiqX8fWABfMQKo0ARtO3cP4ZBU
j36p7DxQTrGpxKv0Kif0i57Lsv0XmuCcnUvNTKrrCx1Ym0GoiEcuKExrb1l4h3uws4taS/MxKdQ3
o9XsqdK/bEipCHsSwbUKuDKZb6Skll5DfFPRSROGd6tBtxg9quDtYR9/DBJcWU1Nix6kBepe3hhK
7AYhM1dtUKc5Se35o+/Z+VaaNCRMZXzl4uuF/4rN90kJolkVQtiD+4aOTF83xZlEapreyWLdJEOi
+3wPVnEy1d++jLXqcgN3s9KSwYZ0D9VLVzkE/dF54u8Bxcq6bUKiPnb3jCPnCNWkH4UIcM9bTHkH
7grf21LOQKyFAnrQDdALV+rfaJzjb3ahDsaaWGed+wv7BOF1BXfcc0owOI0DSUZrlQzzoty5HwBK
SapOZF6ZtFUM0aZoDZkPtyvccw4nJvG9gmDbhN+CSBqWwHHqzNjFFbTkOw2Db+5E16HvHWSMnloe
2Ga5TaC3oj1o9kJXIEd8be9hK1hPKkYng3JQfcBPs1TFtD4FNGN2qPCw3uO94pBTdsaX/4xLdqyi
O8zNuYQNBAb4pCji82gr0f5Ow4JbJgyz9A/iREuefGhDqW1Vm5zjeyC6j9nsqY5bNZjW2KBlQeW3
cwqQL4hfLKJwmgXplRjpt1oGBjrixBJ51dVCqWOw67Jb6YTkNr1sN31HFCVpfjPF8zHxl6ix0q6A
9wYEbZdHweiD0z2ESS22u5Uh+muXkmL8FO9fQKKvNGayKMKURfXFNT0dMw9vMdRK3GYPwxcXaQ52
qmyrPxQugxctIAKSH4vCT7ykNk8w2gY/9sXwhWzMKhNhKCBFmSrYeZ4DPmOrXo6hKJB2VTD6b6Jd
mZyO9RUV+qJ1DfK0E+TdkxxuNWPbL0Y1JIdU1AxZ5NdztAceRxffcsCXBG0ypX0/W2gGkefTLDoN
lF5igfTopjXZTA9YSf24DsyskeK7TiYabr27hEXFN1vJRTkXqjPThOxWIzdQkMFZLvP/V89D1JlO
tqBQ7q5wIGxrPAvyG02p/P/iPXi9vuRLFINLHiHYpdavlv7XPng0cv8BdWHT78LpgkFlBq+N4wC3
7tHQpQYgOeAjx/JNV2nG7AxYliMosR7478dmD1l6dPFzc53AL3rI8YibbKcdNaY6XTYHIKTHXxcT
fz5sz6mQGbCNs2AbJzRtT7c/9dTr5AtP3vdgv7elPTHMbV3F8Ptwq0N0gYisuxw8H538wzyAWFfV
1YPVqAa61m8S6flzQtVk/ZvL27ope67MCQNOowzntrYsxDR94IevRYSqcqre/sGrJlp+foMKIbhl
7o5q/cNlpkDFRagMo/FeogZWMcmz76LutZ9QZzvJUrZKU7XKIjjIdBeUsK6iABYatR1lRUttO74k
ywH1shUHf3sX2Tkiry6lxoibXsRg5fFb2l4jPXFE7n2GZ/orUly+YZN2eKgQCSYcPo+9Cnu5Iqkg
3LFyZclMKmrtOTxOptRqsr9J1N6ETPOGR8n37/6/MosQKzEC6V9y99hHUPi8a21iTn7aycAYZN3/
VXD/tGVi5JdoStkRFX5Tt9D5fObOAQ6rAqWPzMq5+bJvSrcEurYA0aN96cX1qo9ZH454I+xyFNVL
GOSm0hdbx/0n+TUEwQTRVKpTiWI222+hOD5AWQYLYhNt+NtFSKtlX9tvItumlC46WMiFn7P866Jc
I88gMQTcRl2qq0gwbWS9gDyUae8b/eqBN7hn+1qS49Qe44qvOpEH5Y2R2z9u75H2nqvJh9ccjZ0D
NZ9/6uGWAaBVGm8LIoNeOihc9q4CADhFIrV3QrdDvRRIEWOUDw/P8x45OB8pcJpeKzj7zxBn6xKO
hvUC2ItXbA2o2HNY00oRxOx/YK3XPa+e+pz+TODF9nHIJZbhITPAaf2rWbEkr56qHJ7HWcGFUlxM
SsJhhlKXgvV+jmJFFmxukr+6K+9PW5c2cYPUXOMxX9/ienayfvoSJNNDRPRPkyCi78IVvOg2M+ZH
w6VuR8ZJ+r8o8G4h73jicZQ6Dh6rRU5+Bc0NZaSAuCLtZsffT/T4SmTUA1PWidVlcwz0X+zujvFX
0CXdYnFQ0NKl/4ExBDPUp7DAR3LYIQrFV6zgS2TGuDwJV/l+DvFj/yyPXYJiqBu6LN/zIcM1CYQj
WIV8tVpBNBdqtc2YRe+v6Jrwd8vkzHWikzgNpaQJgCX2476u2vkdeBbGKhzFVelw9yrKZ3NDtmUb
Xv3M7w9yUpqcwmkz0+aQw4rlvJQjb4Ahx9BsLM+tTLayM7mOvQtVk6WnZYW1xzMf8mOX7WwDVI2I
TbETngC3kqrlumUVa6aUaOgqsjr+XW5Wf9pTzdk7cp0wnhpA+hkAu4PyTHR2OqgWP4JPrMzgN/pL
Jy8n8IA/I4FGqYCtHDurtuIbVhp7m30q2q8Y+vdJW+8F7nCBnsFSOk//M0YxfHVFzx0Tgp+TYw/Z
u4oEARkVuqbcP5hxQS1Yiujnk/nCAHKcP5OZNyOggXhXuLxy1SgLtA6c32nLbde6RgFqIU7p7r1t
IQvG8AXIKXoZjuOSiq4dlXdMkAQE4LKS3spQG4pPXxPUJ/39eMntRkmgkqE6aAudIpufJT50fkoG
dqZ82ggEw4M7IaArXW+56K85bIYZwveDQH+pGLJUfAk6IqXPAC5s6vbSZnJ3PqUKX5Yd0fW1vrNF
l1ONmO4doqR9TeRNHXmWuup2l7YxgWi3QD0ZStf7ltlsoFaqYqaAqZxgS5P7nG0fvRThMMbN59/h
b5rr3GWB04CS3snBAMOnSsu2DHU4g4UaQH8EtYI73SzgDbNw5c82eDjx73WljXyJXxAzsvjie+dZ
1XUy5Giro4fmWogD9aL01KGx+Pfse7PFSdr5OQ/4LZ3bXyg/sC2yeHSrk3zLt0mtK8wTVOrUsp81
sln6uuejP3yK2gj+8t/EnsQ4Q1I5L+yG+H9xsKd9MhWX4KlO/wJWCCea2Mb4jisK8uJbKSX0FMee
vi0yuxv8Rge2xWekQ2fe9M41/IFY7g2FnzmPnITk2SMWVhyjYfo+kkK2plsx6qoQ/yTCnE4l0kbM
NnYDKMBy/e2YJb7iEdp+FaJyWl++xZc4rQ+6lkRSAp9TCgmlsosAMlqCT3pI9PHWXe4o4097K6gs
zGmYd2UZlGd5VRbVIncWBhAciKbAqRTWV23lMOaA+cHNfu/sOgbzrhsHTRngM+7uYN9sveb/7e0x
1d4+ICRGU6xR10zjjkOnpIgj1ZdEu7ngxTE87uKsYTaGM2uV8XE42W5b8FxQWacnhfv8OGrtvUGp
hbDtIOuRbIM5DpRwBzJ9cVDV+mh59Eg/Rmsm2qVc5NlDF9UlENPighPqq+PyJXFezNoiRh1NjbHL
KHpHLkIeIK7yugOMjdS500H1AMMfTqnFiHEty53I+iRp0TURnNRwysG3YQ3gCoPKYLTkFibcT8W/
e+M6D/1XN0wsplWGZn/irSBeHLKILnw+G1WPcYzCBimMiR+IhoHAev4PsVOIVJC6lP4Avovd1TF8
bjkmXzIwyjNaicfdI42AvxN5Sy7jFxtMv7IBkBJGVGPzO3p2Tg4AmDIaWGhOZSMxBZJjKiGtC84u
L+6EbkDdZc8x9uxGGosrlu9hUDpTUCHKnk24JZwaz9P7RWOUk2kmpyxXWYfF7JFW6f1hq9jyMc4N
ZBp1p8QNkJ57CIqjNVKDZQcd79n9vf7Y0PbRn39PvnQJUtQxRk07pUQhLx63Ti0Fkg57rFaRfdXc
MR31yQjod4h52l3BxGIoMgmoJvN2Hg+L3gedZQbUvCXSAkjEhhH+yNmJbx62v4Js8Z25ef91GSpR
skIM2TxSrBFT1lEgLWu8IqE/bISJmRL4KJox1U3Wx2zvXvkebjTOeTtVVpACvBFKZ1PjCEted2eF
YwpZnuTRH68tiIr8eD5cjy+A64fz0Rbgu+TvvdF2Ux2uaqK+KR9cQmBlK/L6trr5Ye8mBSb16Rg5
HRMcIP/3OUM8KOinNLImFUdyFaUq5y9NKiIBCH/ZGArnUl5bJPamIjLR03jGazNJON6BfLSGyYhM
cD6AI2tCgGZve+3TqQKiKGlerasrhJDtNsBYKt+TPdxiPr93W5NDqFOsptD2Qu7Ue3IRWe6WhRsL
dcaxKPQguwyQ5hQk+ja5Dr2Py4ksMD55ugLbRxYZHR/M3L4ETfxPTwMIVSRPIn4N78cjUgYkm9h5
wgq5v4FQ9Mt54VfF5e/UirDISqQSDMwj8I07jCHfm030Sx8jrJR5UHWilwhl0JwrEAd+tHe108/d
JFqzTvl1ieqgeSzacBtqf21cX12zdSzFjnFCl26Cgd/JBRFH64TDjDfPUzrh/bc/52YsF+4hIIvh
ZMKjx+xGBpF2ViKM6hUIpc0CErVvQ+jVNLcYWiFBlZ50QyNlcBtR4r1U9ssbAxPxVHkYXWDSeDRS
aMfEpWLa4Zj0Wc+zNS6KKUp/EIKNw7MBo3Rh3oPGFTvGEqTRcPiT4AIlDlde5g5kpiIyD1HCVYMo
7ZlCyc8arbYYAbiEHVUI3eqkxLsIMw1U4KxYMXeUFH/H+LTDuBZ0Ug+cLyT/Rq75wKHkyqKsnmef
rhh/iIqlxGKWiEmxBeJNbo4YzBhwEhTYdRssAHBf1Obtwo9u4ysCU/iISZEpdDW4r/NxaOXaiiGT
PmOB64m+ft3W2fYUSAPpX9GASt9oJFhUfm5PFagWKCr3f19kzOiSkkKYJKHzt2VeHxKttRLFXR4n
Fxj5CfI+NB7lVrhyAHn6fh4bT14IImiInT8GpG6RDIeDIY18gKlaX65JtTbFN1htwNBWi9JCVtUn
pF5KKt4mJXeseB3R2EysGcXhwEc0WGOQPo76J1jcpaZ1mmpARxO74w8nPCYGpL0+RDFlkLqJvn2K
Ze6OtErISPY3ab16Gq0iBKpfpj5gjBjxRl5Esq/0fvCNIQR+VVo1w9j8lQpEZ8SGy5OIhloItmgD
8VdfPv3ZkkCutcvSTXb/nWNVw4sS65Z1uwUAQV3KWhLWg93lLMiu73xVufrtIeRFPwiHey/zvM4J
LP5zzgHBIf1lsUotWNc4QV90GwoyPWOREu271U1XiL3eKldx6u9RyJW6+z8l5r/yh9q0QQXSRNwn
XuzKecBLYrchrs8zEpCQFBvxArU1Yt/tHiMEt7QKOW684PwlvBd1r7cjevOXMLX35u7EO2IFu1qO
XxCKx0cVy+39o6ALTNEUHxXbAW6QCrc6iGEL2x4qxDBTP/ceQb/2TjwqaFHTBPViXOVDly/ZaImu
QEdD33Kh6woPMS6QsX6BmI2zBPpaUV+zHBhrAb/Qaky+rh9pkWtr7VaJ8YKA3NQz7XXhUocQaUEU
YvwvYN+mjjL1kZvA/XP+uNgq2u3JL7frzhHEmozLxXoF/eWbMHd7iBiBzu0Mw7FvvphTtBpK6czB
OrhcgMUuD+iAw36faHXjtXblfzOmWhNy3klglUbtqsZgDXFTvee4N2TpnMlMr5f9Iw6L+sRj3+SP
Ia7zN9fsJvaD8q2sec8knWkGGFq+uVS4lnmBmCZnu7S2A7IUVrb44Om5jirAQ3/85nEYENym7GHj
LGyTtSDx64nL6IqrsDRjJcsddbH4IxQXruNffknTjpuFHRp0rxaQRu33X+XFuB9tUfAjkWsxib5+
3mfvv2KtEQ+pGNjT4UDZJBZqyin1dYukOAPsDv4kkLgAGpsOg+wCPYZcOmu5eSibAEOJ9oDXUlvw
Z05wtWTFd3JOHPEorveUHZeOspy5PYmvUo+SJR7E73ptzDoFAuQROFSy2sW5ireleMdOA2gCdcAN
Xtv8YmO3HhetjrGVW4lRLIuBkiEvKXm8lgE2ar8x4FcMrJRZDh82w2cMAIdjk+ILsX42Wep5EJKq
U71N9H28OKP4gHVr6oH51BR58BUQABT1CXswi6mpLNzbRT9eijs+aIq1Lh3pEVfRFMAs0m9070mn
tdQjpIvusP7kQHpT+HD+2YgB+HM57AtjWhNMUWdRDEx+Yre+YqJOINwuypQTgfxdpXHQ27tnpcJ5
yoT+JtRIrRQuSTT3YcoQow+SlYGPIqJOja2HJQoPGepmpeAsrOIPeS5QDZkWMiF9NE8vJMnbkaZw
C6BbouP/IrJ0Zx/e1DRsyYx+Mv0BOLNc3I0HcyTzsiObZFDX5ajgi6QHV8bIZxrKw04nmTyfZxJy
BQSWDewP7vO2UHXFo3jRQj9QACeis+Id8H5JzcAwFT0Sq5sZG7sYA1ab2scpZvLOVAJtn0JlTP7s
fZ1iewaxRjZZxcf04MELFezZ3k0PeHaPBP/HN6kgwRp6fYqxi1GLb12sLjS8NS2NpCQDES9FZXG9
yPOA6putPJV8FyqCf6mWdf4i31NQgsqqQK6+jFcefRnDc2ZiZGeJQ0MDkm1yfmjrsqFePe4rihRM
D52mhufGfy/s7guF3zdd6wyEeK8mcjbW37QQuRLskiVgtv75aRWIIvzrkoaJHO7dB6NUy0jAJ7j6
Gx9Rwsdo13hXxOF7GC69Qb9XcV+G7Uor4MeZxRS1HWuFa8tOXHg4AjaBGIyu8gUu21AfJ6Y1wjAj
oZkSZD2n/0BgyzZQ8XVUpYd8geMNIm43LCIFVtEKXhwypmc70fdHHuNCI4w0Mn/WGD4cHjNQC9Tl
HmnfwFx11bawsLfH1ct5GQnkVvKKP1Lf5h5B7ci+6/ZhLQTfAiBsGB2Sc9nyUY6YJpVjj6zRxKGm
rDn6h/4iWkpCk+nElk56Gx959/tgsWtdhJFM9YxJwLuGZc+1fKDo+ubwgDiwDoRyESgDw5k3fDpK
9EKjFoGB2TVtftzsBwNKnCe5CN1Bgye1YdQMOA4SyTnYQ95ULb8lWixtQB1Y5TAT9eVIAx9X+qOd
7JjtTjDGiAfWhJuDcGN85+uXoGSN2LY6fVVvxW68FpHr/nfmHlWPjZw0Xog0P3I0MCUJFpRFdtOb
JhIcfBlj7lMpCOdBoU3OVBVbP2vDzq/IeQw4nybIem8azvl+1R8acpeZ/3IJQGLMuNKdE/cEDvHS
EodqEE+0bQMt7b8UrqHTfHP+wOdHS9nXRlwuuuC886mnEJEAvzdixGZj3dgdFWZVHmsYJ41LIl9D
oNGAb4BdpHkNTzEnK7ZDpJibE/SKiZQwB025NFmuXPpkM2VSrsxge0UlkZmFNKQ/ob0KiL+VQQEZ
NmuN2ZIOL0Kh9SAV/xnwTnBz5455ZhpuGszWQEpiVO/fMFhjqAfQ0GRTDlAbZAPBu1GiB6OSOxue
hSckXZBWsV8c5+UD6wTQLXsXhLhLM9/MLiuO5K+sOzHFOamnza7jpGjZuI4MYytkI1pG13J/Kq5K
mPHlW27oD9own/jqJHpI//rYV+j1j5y5CoAhnoSpvQrVVvwbOyJFCcaXsstFh35U/M/4iM+B3uxJ
U05Zx2iAcFppTFlgXpFuZToJl+L9ij0nkfgIMGw3fYTHMtmlLfDELbMEz9AOhS8V6Kn4tBQlaYU7
c23+I6IWg0E1rTlItkLLhNDdI0jZmR/u8Dsy0+z+i66qbGfadyCTOK0Te32G6d8unemfYQ42mKT9
MjuTjVIYievHrSHViztk0Y/dlAkJjDKyzp6WolVwRb0pB8P448NMBb8ZMOx9th81lVQtDbfq13Uf
hPjx4ucfQVXCnD8o1W3hIGdFKI1HPJrjZtafS54f8sFQQcH/X/WNU/iyhDz+f1loTghOpZmeLdlF
pc67REJ/g/2wYpH/SiFq5MEviYPYsnUIb/MmPil0wIv2vcuWLc8PD2jSMHevP6ZxIUIl5ZZo1eyR
kROKachy6nyGlc7TcoFYV4xUmatXMcdconqtGmg9EL4rPi3lz0O8WdCCLNdEHLWCr2DvjrdQkeAH
bDjkaKpcdDW3OqJIBz43Yj5wtReDnL6r6X7B2pZjUI40xD55TBoW5C9i8lvRAlVAEy1xoetjXkBW
hbGQ1ZBwU9ltNR117yyYpqZep5Im65UYG4UJ6rIi8DkFJUmdqhmY66O376QlmRlPbxn7fDusGeYu
8j1e6Aalq9R38BYLYYUb1sgAtcs5itvq88zAG9oJH+BMpwn815gedTQryuENwwjGDxsee9h9NKNt
Dmtc2mYKhhD/oeTPqyn8AhT2lDeUNod75AxpTiNXvvYA5u203B+Q9osO+6Pg8liW/x91u1BPaXyg
pziQ01prmjNeitcL+7Y8jLP/wf9r6w+bf1yJvQoyfUBxJxIF8F+iP5P3wWTnBE28ThrB900hlCwR
ZS/Kh+mUKSbUskg1s9PAQ/5xmnKp4EpoMS+zSzK63k9koGM738m3JN1jzcZASXiQ8qW/9nyu9qxS
CFBdxwaJxoQJbihwACB/8dF/gcEzJkV0gw6shN5M91os7HUfH4/S8OMKlnST6r++2cuY6Ge2NsVz
DT55G/fPAb3Vp7hM1YFDjzhgaGGQZFyNPy/Ip61vEBFFXiTpYFTNgShL56Lvn0dueFRJb+sjKCkx
vpcnJ5vqS8Zg38y/KPj9EicDbO86b94iAdj5WA26ulFJSCu2jtpVbJ6lCQPyckjQ2hJux4a8ZBPJ
7TAOnzJdrOojwSyT0fxtkKilT30GUc8Ucx/0IDSkV1gH6MX1Hrg3DV1xGHaEDfq72VQgQW/9j+xZ
F//WboUhBO8Ni8SiHlJGdcEi4+NRX9QL0mVjo6lLJSOQAGKisEHDjOhRNgx8NARNOw6FS0sb1Ie1
hXRHrcKZ1Ts4uVignNDjQKRbl9EVrxL4qF5P/AuaLCEl8jGzn9H04yWGC4StGpDzKtGB/L5fZD1L
pWddIV3hDMQc7zWhQhnUVuT10raf8usGMBxxIuSAuoHUR4BnDJonnVDBne5TPy3alNN3z2CpWgWn
8LRpl6ym+gYY9cKrddDTuLtyew/0ppYzXbwyU2vtp5E02zgDmSiqyoc9aaNuqtK0Ze+09tRZF0Uf
TjUii2Dfds6ff7OThwhAOgDGPd5CcE5egOLOdc7nos0EtsmVfg8/3JTMcDuWYSsrknvoIHBGYaRE
6eYEfKAJFX4GhyADyvPNbmriTjAkU5QTGzlIfXj7l/KncjvcKdSVBgvVO/p7GnfFzmGs+YNEvfSE
EefrDLSaRRU+fSKZnuBqlRKcRwSMJdBdgVLgC62PpjVq/gykfLPILvxVzJ8JFGbY2dSK3Unal+Dv
Hvy9fjNK7cmRNBIKOyTBUSb8s0r0qKqzVpzVbWbGDSQ7tPN+1hEprcWO/nUfZW8f3IOv8a1SHxxD
1y8QKTxDYzxkVVlkZaTE6lQpymBvU6iMWTAknAmkujS+jY/QwUMrFTOz6Jnh9iJsLXncsRM/yd3o
CxlTB0vedRcg0wGI/fVfRsDypXTanXOi24wsZZySYLJUkqhyUY4P36vn+2/kQns3t0C4D007otjm
KhqXeJxIEGlBJAQ+lkZN2CUIFYwNdxZreAVuea13WhqRbhnZgNzly4gD17oSR+pIeZQ8TgHVgDHX
fgiUwjAi8gZjVOd7izrWPm/x5gpEkJcMb/A/zsrU2R7Ta2NuJpmQ/hPV+bn0Yl05iGhkkOhCYiJ6
Zs0E5QjECaxW23uyHPD8FXFHOHDagbmvSt+jSQkukrp3YLnYEW9GxHg8kQTLmg114ueod1PoQKAE
7yJLAi1JGWwX/A7EGgagSRaznbxiwZoR/5rrE09Im2XJtIdLeu72KC6MLWxGNTMc4v51JwgdlmZH
5vp5EU/zlTwbowpxoG5VoQYl5nEEZSnbLuJmJyHFwOZ6xOQjnLdI4VWmB6HOh/6Rs4fuc1y7IfvU
g7WBQj0Tjnxa1yPLvZZrjZXtm8Mv7flErJAhcHVySMTnoyDYJgQY+keeNR6PO+I3XNJ10oPuoa+6
MMK+ZH9Ewc823dXZcsYnSpuwsVxYyXYe/OhWbCPUUVNACKpNvO4kR/YWIlNVlbt03bzK2jV79bsf
eT2NvvYImEoBYzC9CLWXMFUqBeYybWFSiL0IN8e1Kt5ZjkLz9Dqtr8MoohdfB5pXg6fRR/DpTAa4
myQ6w150Akdj1spupgc7UoG2Nk82/xQw3fM98yGL7vEa2ofFvIQAHc3OAMrGSSWeUx+LVnW+06r4
gLhr8R/WXRrzuTv+dEy/Q462Wfk/WO0Sz8nqZje9ePlZP/XQwvpmNvkELvZWT3hcvNr990s0NUhR
dKJX38a0ww/B4ujO7ShEXW5NI7hH2AX5NG2+y0kUaNv87guY2z/I1AiIq2SpDNMZt9T6tcXA7Aos
Ig9vJvvrkYI0cJ2wWObs1OBWj/WTBxJaQylEbYZAPGwJumpgQZbX0KApPQIE3AYJuuLsyQSgFyCD
dMv5N3le2Yhs8Rr1fICPQ72aYLl5ZiwQFYIApaGNiMAHLBL7TKci2j5g9DSzmcctxTyc1X6e0K1t
hZCZdtXhDlgqqdxV7Vc4sM/g4jP1qiO0uB0KGk5reQcNTjT2y4msZ3EIWr0EOgfuMVqyl99VL7ry
I+ZUrFZFgvnjSW8vVom5lMZrauCL51Z25ygxEFeQjpmjEVuMy/F/CkRbodiqfEeNeok3V2TgPetL
lwuxFGKY6Y1r8nmQZ0fwo611Zk15WMls1uRNb45hbo9Q0jwHS0lrYBEUOOyPHj3OVU5cJS47flx2
H49k6DSa09dCF41CNfOowOcNUJQbKLMEjRH+jyUcPQuXitQn4dCa6yEmYcDo66YeZOTbkgOyhGCV
hBSMv2ghCaYXLKVe/hODC2ySp4QSKZFdNUb/M/B2dTNMieRHa5i+sf5O5n2S62LzcXHbOuf5PZIz
kKC/w2/C0GbOD4GKSGwWhdE3Kjzfia39PxxRv28YhyhQOQOo8MduGg4E6mbjqcM+6mUNfgBfrvog
sDq5mOnhfMvhdqv81pAcb+Iva8cE+l65KIWJdj/dqgjFnbclAZDxTgSfYb+n/fWxztSaulhUVf5o
P/9JHNOqOgmp1rgYamqcZLqjISCy8tGVthCMa9zwKqlFB4AQnFcs/sIn6BC8tzpzjvZ1c4qE+blc
I4UWcq7DXwNuqUMzrQeVnLa5AnWUEdlF3wjISBLZeUt3YZYiEZv5Ipwd+OlEABs8pwuhD+ot27uf
LeTfyFChAWMME4ID3Z5eVX2wn48cr5TubmI1lttNxkUptbPsIV4UPiPT00Hn01ljwrJOamqs/ON7
5pOai6csK9y8WHLv9QRtznGxKZkwsIcgUGZBk3ZFRwHqKSIMcEjIITPB/j4Bd+PgkVAUSSJE/2+f
XY6zqzV9RmLXjpU+XXdgfwFXY+Z/iw/wrPSM/sfFwITryPHPPF8s6R2DCXW5hMhA1OQkwTI2u4gJ
ORwBUBa3a72BUq6Y/r3dswh2g9+fMAWyrsBukF+UgW89a3KAhZgGqewbWROGWD0nYbpzqEze7Jni
uwPP3u6IKfhzbNzPYZ+0bmVLfPZcS6Il4XGoUFFxb/NO8+PNJWkOvnn8lqMlpqEZnVOG1Ro1rlms
Tkt/WCXBzAwnl/cF9ejriaEtYcAH3L95Ht7Hg82YSdRbeCWRTQfNBYk74/QSg2rhkqretrvWgJY7
T/q5i0FaQgEC1Kwx8a2kpXqLponcKpQC1PV3DRAZhVggGamwOiQ3aklpSltq9vTwvaRHvMJuvgoe
CpX4r0RxTWzS450DJaMKQq5k39cgtbY3VQJNj3KQxx4PrPHYcw+BuxZYrOE4vSPeUT85kU9Ns2WB
vS2f+winexsmong5wKai0YGl7HIXOP7AYRHqWrxXkE5nc9QbQFSwLp6ra/WIKxpnj0FAZKRxFx9H
5si36gd5vx8wkXbt1Qa6ZMasacH0GghIfejsvnNVW1AcM5HbQ95n3r+/GHi5+cWpsbBJusBpolwA
cxIQNHrtdkwrufCuKMPpTs6kjhlXytIBmKF1FcYcCY2v02ZMRTmCEv7C7crL9xf/tAxAfsj8P2+v
NQ+s/xT6Ki5z2MmEVJA1biHhcmJWwVBDj70OkmKgTt4xJK0jKMdlCXmB7g/cPwrtWpSjafzLWyKf
E8s22dm0Vu9XXFMqXEXYoe+HOuXpu52zPUHtn7UsTUrWrFzP+AU15SWHZ7fcRDH2BZK+1SaGHFc4
NZqtihmpF3zf1lJudOzaAl4JyauBIGa5PMQ4vMaYkr8nIdBp0V5Ysp5FQBGzVYEa0bIf04t0kHQS
7TNvoNwK8It6Y0rbm6yobI0C0do65xCOeslVOZx3sTcu84wtdnPsHzZeiI/OMYNjFK3Mctojp35b
PU4F3sFyjerKDaVDUyC+//Y7CmMZYefvxvMIkYPF9yyeV6ZqI4sQhmUQVuJyPFYkhGqOvQhjHoTB
a5tAIdDUWSGY9s5ay1kvrOncl3XIZBFyrcvJLur1tsgHl41SEBKOHwSD+7FVRJlvPNTdWR/PUlVF
daj+3uBoZzCR5+6VMiq7WZ9/KJb2T1Slj5cLNFW+/mHTL9ut5zmLbOEdy34TpRugQb/c3nxVQWhg
DCLe0Dq6eL0SWLw0jnUdJHlYjiGxYaSQL0C3u3ktauYblKfLHwVmIpSDERtxQLi20yY1UiUx/2iu
EvECuHSHQwwAglqaJE2/r6OBWAS+XjtWHIAIBZNPb5cENcrHkuL08ut1LaCe7NxBqrWQ139IBs1q
OyfvkIGuvIDmulyJ6YPYhUxEE5BsFiD6+9JOLQn4kjkEhd48TDQFcnXWTyCg31joDfV0TcHVG2Qe
przD/P4JLATARzynHillhBwFw/JBTU/Ey6hCGyr6s+iEyuCZfkNUTZetALSCBB53MkKGtMQ2Mbx8
qkLN0VDQiHiW4PPCFjJVq09cOHLnttDFlduryeDbhnbg+7rlAmkYwAKuaV2FSY/4Kw+48Q0JrUk4
Rpq/icOMXnOTd65XfyoQ0yO9vrp7jy3a1SjHXGNkd+icY2eK40De9EaQCpMrEL/b/EwyYMrbiACK
CXQFWT4ULV6lh50roJI9GIyFDekLb6j+lWJERbKSIgsGDR/61/OJSQ5MDFA9yjVE5cIgBfjQvoB1
PsmmYfMhRotNjuCdtgpSZjF2njz4fdWOeQA+e/UK8NkGVVfB9bgUyAZokA4rf31H7tzUvx1Ua+zK
lrBqZ4dxh522RvE/flpz5B2Hj0yIzIU8Ghd955r47Z+GvnFTGUT6VnwD0kksANKdt341cjSVAS7v
R7F9nFD1ODcP+xHcW/OxZRLyngEqF2hMQ6ycPbOCVfrtsntUBq1Cqv9drOBMGuDuCUT5jx+Jz53u
ot12afPxm/XpUAoGq6CnkEpCtNTI9hwxkXWIXAdm3jsfz6kV4VARjnXAQgb0PlGBqNtkpiIc5u/z
p/RbUxFh8YCuUFC0PVWIlFYWeLxfkWKtSUAhJcyx8nGfsikedFk9GAVhxWunN3oJ1h+lWOi1zMln
1uNEtPOIO19hb1nm+y7SF82G3GwPkqBK0CDuwVh3EbHvuneG3kHJpwqXgEmrN8JzQFBhNcndLCA3
YFc3sn9ch4/sOyaWjjAVU13q6WxLMIl1i2QrPWyQ449pMiechRw3tKIBBKIa770choitMSyDBzTP
/if3Gohg2VaX2nwE0khxT0FM3d+o/ZWGV75R5NNsIJdL+eXx4dJSyI1qFB6YK+br3N5Z5x2/1gDr
FsPhNHuHD1EFuBKqgSZDxJWat+Mr0JIJHfl2VyOt7zKBAZBQfP6vooDNq5pxRMDCYlc7IdLtEeYs
OawYwDkvjmkp9LK+zTbUztPcJwIX9t9yMNIpCywWRYx7+4IP+TzoiSlJqFp9tDkp1mMo6qlc1Gx/
ktEkmUizzUFL4jlOWle/eKc2frzGKSMnB8wj/VjgzOnXpRsonLt9X2qLf6dTyq/i1Vabq+wk34Ny
3dQaHnsKVdumHrSXPgnHmO4pSOfPl3OWomMNHF53dWLHAzA1vADQTQCTXZ/sWQz3hcW2XbJTno8+
4OVApip9xQ400aKwy+NwHVPl3sRouqpgtTO/l9I1jdV6HzG7j05A9KL8l4pdYAZVGXpFZp4a9t2E
rHy2nR7cMcBV1KiAi/oN81OO7b6YU9XVv9UM4J0XJCWzM6AO8AOO7dZL13kD9w+npxEJXkuG2J78
X7D3WRXinWz/2wcvnCG+TpB5aCMCmVAeQRL8xz2dDOmdQLeSlK6qeeJtDUBnCjuE4U3cy3bjd1Ue
kJCr12X9yxtSTNwJz6n4MQ1vTF1coCVrTViQ2KVaR8gsP0gSAVDMCUNWakGK+eNu5nTA0TGq6Ovk
/Jl+z7pde88TNkW8OKoSHk7Mqo1bUgquKaMvkczvRqr6VzFBfE/40g9Hi2Xr0rJEmoB3af26vya6
BLLkvdV3gLDJHn0jRJDQDzY2GQ2uWhk55+BRYNATAm+IkGfdQEDxCKWAH9cl3XzvcEy51AFXwI83
7pkcEVCoqN3187hMYlKfBvEE8qqdmJoMA2vZeszHvHNqPB9UY4RpmlZFHe0MXFBGMG83oIkEHDeV
2PiyVhXVGKF2n2Xh6WJbD/cWrJp8YD2zj9dey+hQAEDSu2GoTudIgxby3j/4n6iWf0IX2MUgc4Jd
gGrT/QTiZZVoZjVJFiCiKQGrQmOkkfINSvvIDnvzCl+4+OciK+V2lt5xQhXAA6AcHthVYQHIU+py
pdOrrBVR+TqVvECnMHvbsPz3WWVIyDOxlYXwO8UhJ6d0yPT84ifx005AeC0PS0cWsCweSMEKdFbF
xOyh+LGUuUbH6tAfjbX5FsSoMVNhZvfw4qrjUNDDFvG7eyG27gyzxGRNub4bEIs91FP76/FgrDQK
oYSK/DPwWJup3oH52oGPg28Iwk3AD33i6OKGe7z+fGs/CyWGFUlzypDaeegfzSlHpIWfm/ezdI1/
So+ck5tFcGPtcISiL3Hs8wXPVMqvxnvmAFte23tt+qPmdf1DlhfiAN8KzgdJwfqxnOQ/qxs/VFXG
SmLcyaT7o4zNjuKkhxuX+KJsuLM6R4pFuDgvBgwa1Tc/rUYeWrC3ZJ0R63qK+0LnBVKKkB0HHrOT
BZpx4gEeaxT38/YrWvLrE1i7M7zNE8lBWdQ4IYsBqt+WTf73oX2u/gH0XDLW0ftpPwTBIMYFte7t
3nj7aOSX/eh0RQIhVmZFDgiWIRmYYDfF9tMNXeKlq4JS3h/LcpUsJaDBlzmO1NgCuxaOivDpwvdc
AirWuCziYMWO5iWbHMTByy6JESdawXl1h2vbPcxBrCnl9djXPCRkvmzsHJFnKHNoa3v8b8+21tRh
PCcaPeOrTxg0dlyzHe7nCPSYv145n8LjjiWYq9elxxJLJwQOLuP7L90wzQibtx6TU/zp8Sn7smxh
6R2/m7zQFTe5O69JvLUyRKWfDcSraG3VnUw87sD1Vc5NBQ3r/KufvtKkH3IY4W64Sk2e2O7aQR4w
9hh3W1sCkKV8PXhICdDPocRtiMjBes210VdfdTzlwNlzIIh060LWFrPVKFkoTCa6X+Ryj1O2adRp
mqlC9OIPzrHxntlDtSyQoaydczyu7QOAERiny9sgq9EQbueJkZ7v26OoutXwpahIc8VHx6fo2TFe
jNdczZ040BoREovJPPO5sOvDva9ZDFgjFQZh+8eTdRUHVgcaiCaRaJtahvnc6jMcYyqfqDodmMy7
xfw+ZMF8DfwsWc1m9ZOYeZUz6NOv6jvXoejrzbyC1JnkTbTRuMOsbrPpy2emIAojCgvIgToDc1lE
pmToxKit/u7pkUJtOfY6/SAW7QoL/A/cFFVeYLEker53kMXdtOaYShG/qsxeZgxWSrmxAfMRCT3y
cBIDRlzKuKpu+zGzZoDVaee87ihNIDiwpK42D8lpF420MFTSrR0W6CKxJX0VHeLSVJ7fA1fq/1fF
0sb0ajvdarE6i35ycc3bHV3k12A4LdVR4oIfffvW4L/MfmaJ+6gqdy3z0MB/l4wC2YZU68pLvWLh
iYNVXG+ZlEcDBE0/SfOXKnWI9Jz4unvuu1mRhbmJ7mf56TQ/cicrIGscxTqGMdtGpIOtOiUF6ifr
xQL8cZB92MlxVkp/XhrkAig0pgC/CGBln9gWKl5/RSTSOcWmOXU8m0z80LNS3MUkiY3pHAEy4K8W
OoDCP59oPO1Er49Sbw1bOkE13yfRiOihLbDliJdvr3BR+oyNEvRAVoBOe4Jlitc3GnCt9JgwyJZL
ChumL91I7Jvqlspi2JennBuJYXpdgW9wiz98TsuleijDAoTxsaoP8mkSJ+8afhlSr65ifrzfrrPk
kdJo/E38K8NZjkq6reQQk0OwFFs/+arwWX2/h09haTvtfig37ZnJE0CrRU82CavMYSn6xCZ41Lmy
OyOIQyOD+uyc10PtLBrA8qHQSBA/V4Rbb+fpr6ctmVIdfQwDQVrWNaRj4rnfC7iso6l94ri4GRpS
ELkWxkuaK5PCJYS6oTf0Tja3Kb3dP038IrWYnlc406gscXaEN6XQHXHiUz6NnaaLYPKxd3wSD2BO
FoQHuo9mGeKB1wUztqYE7irVZQ4mv0rVaqI76GvXMueFLllVQlRnj8HdRRCr8cjCnKnFGb1OdH4/
PnR8M8gFEjelK20IYO5eFJvm9k1r8goIZKjlu1p9CsJNlg7l7jvy1+tyryB+LnL3sOUiT3y/icdX
+DPzIZNTTJkFwhFG9MccltAz9kIs4KD0lh8IupQROz/l5qWR4GpuLxrNXZRtnCXWnjZYR5Hdpxbj
xw6EUk+LYVXJqP4yKfoXwmQx40ns2MirWjS27K/CH00pKz8SNg52IZrwmnYuIM9xc649jCunDSsG
72VAOycRoYFbTGRQB2A+de9M7j6UXl0KShf7V4RFtcNBlZyJdjvysGxIRnXmWxGyU4eR+GQD5SQP
WvcEzzZB27dCio3lRTq5zeuJNRD7kyvoc41el6KVx4VFZcEYqdg66NtloZWSm7gs6dkmfBbJaug+
w+g498OcejCSrYoUKnrnioGCEarBpj9Eh9GYoV3tOPnu+vpePx79rYrITQv9QOpnlzUIlpCdbw1J
b7ejnvvyTLkMeqfUQgh0YI7XdsefwF5J3VP++BVggJe0uS1o7Ldqdk8nrx9GXY33L9PrFBat37Kg
xx6z5+TA0EpdRWUqP6g0sJrYIgGpHfpngdipY1EFJFQM55S75ZUBweTVRk5kP//kQJJWDcEOAvE5
ha5NIYdbCU2shqYoBAfmcmEXeWOHK+WMPiMniJOa7fNK9m4UXQkVSaVGYftj0d5MFT8s1GdZ6syK
3Rz9/EZok68IWKPDNJhGTR0pGe1YAiqnBYEmq6Ds+8Z6G43mXkszMWOlgKV7Z+n/MugAR7/UDyWe
M6+bxm9/D16l4cp2qbPzPVIHi/2TFDrLhDaV3YKxDbHZVnhQyUHjbqSDLZA5ELgUrBqO/g3MRBgU
8RuXLE/xLvlFKmC7xKVv5c0+qXp2VdC7IMs1DUbKYemVxtzMpXALzIdO6HnUMZ9j7etE7+BXpK6H
oldOg9LYrVzrhu+lBUHxpRPqIZzIK/+hqbNKpsAhPWx8T/cr2gXqGKJ8Zc7ImaCTOf9fOGyeG8Rn
lcVxBWTc2WJxenkzs32o0GWqSCeeAbxNF7bMmjbtoqX5NqODfKK5e63kOUdnpj7kS/LkYyMq5PfO
YwsznTH6wmHhPviDUsRtDI467di0+FC6/S8xjEuzi3aWwtbFbEp9Xa8X9C2ERI0NesqkPzhPyK4T
wz/q2acqL62wBfXFE61rQFuap65NouQMFiLayB9ju+61qaUXgEmAWO6QYk91uCFuH1a8LkvbJErc
NUhk+pEbAuRQzCNqMmd2OBGAj988O9T+Kx54MAlkA0vbCAHqYdAOicOrli3E10UU1OgTC1KLV+SO
lmWrrr6JP4JzAprGIFsH9btVNYzPCiLGn0GltVboLgdtUPXWGwvFus4m7u83gRXJTiUkxUt+5029
sazP4bG0cZE4eozuE5Y9o2OkPBIVdrX6M+WLM0hqKQqbaIARlTOn6bVUlSuj0S62+r/jJyfjutI0
lT9a2NwVbBpnL0zGr130wbag9p2IdoL89ewfqsBKxyOBxBFwh84tQqvE0DVlZpWrd4kxcriat5QM
edP8ISkuiQZNZc0xEQ+PE1z5cCj45E44THZTCxiPcoj0jIMgPEUJZCHwTS8YrThcrFp5nmbm+BKQ
w9O7xPxokKh4QlF5J00cG0EguZ27HjOF/YUXIJe7OYuurLU8lhD43FYEC5569RL/jC96O+wz0LER
svQhdJCQwel3Dv7URfIRiNhunZ37feeKgtWdvmzMIws2MOmyP5owE4Ugv+QDrWhpiGIj7w8SQ5i1
musEjgDQIsZO4MSnP1YxTSdEiToDPviTJX+LCVqfVKXgMlhrS+BTpGAV1EbrsqDDBPCEUelNHh4J
+t4H7HGSgtz+b5ans4l7u3rTj8P7eUeRvapByypcueaiIkzoLYLX1Qzsufhk+BqdaQV4Hljt+Vke
UmofMWuorZmW5hucG64yIu6CXJUZBxFuHyxWKHGmDtFh160uBX9bWvCBuWcBhLy7iDkRsU/tIngZ
V+AiDYQZ0vWY1bocZ490HpkDGe0M60OaOg1kwB8l+BDuS7VoQ8y5dxUVHSV5PIEwBfRjX0ozxH2I
F9ESQaYtxzZzplZUfoXYT2mVg/AxaMPe6jOUF9hw76FxzhXyyWfIx+oHAeBO6gQJZK6j9OsApFTW
Z+05R0Q/Mma0cwFZ2xCr2QYEAy0ic7JOKudbK6aXr8PD224Qmr6MMdy7Z0wrYbyFl1HahsSdlUhO
wbLcyvo5ulSZCzDa1XnzmUGU/dRqA2rZFY0pn6ep0D+BB0mJuKUrA4rSnKF58xbJ2rreRr4/qfat
E+8+1SjlDHpAxxFIYXnLBz/EwUDzpoTLrm8hzOgv058mmPGpp2ThEXcK8bDoDRyYMOpLtlBAFHp9
6XR8dG6WYhPurj8cwK6/J0vyZe23Y1Rnfr8XqQ5wc9tdgQx5eSSMEJnAIs6BQxNJlqj1wfYAelLb
sW++auIkoeTiOBDKjycqABua49eyMYYyhYAVI9Ur24D5OjuPvlBWa6eCxDwDBLgsLdO2MxacIpnq
Goe8wZvfD4KxI1lZ9jwqyppGzvBi15QhCoExXG0qu/3iTnMGujcDCxupNIM/FdXDMY/ZysspNqY+
ueoGG/jHBUf5pkThtXwu4/HcKK5KTctBKS2zjJAOYoat/RwWIQREfUxi99X2XfLTsaWdTMGKQLbH
yuEEDHUTzo5RxiUATmaecGuN+LbIGpjRmI3F7WRE/sXHuRENPI3nOczNeCCGRoooV6/atGcAq7fj
ITkNDp4g+xrsvnXcCvonTwPUpnCQEdUACfBtOXIGgnucGuN6s4/QG0293QgAz4rOW+TyjWmgNsC4
IllHP1qeDg60OwR8u+EZAQr4nkPIvSZgzLmcGsnJuMa5yG98mVz/lTuhPFGXAuBXY6PvV+GKv0C4
6Nm51gEgPao38FL4G84M+ipcfgJ3KRpibx983uiST8xPRSJE+B5Hq+S/IeF9O7Wm1N6VE4/bJAax
JwapDdnV1DkHuBdRmX8ExlxJLE4TkPVQ7vsA6ZfWbZxgVyvbgDrDYLJsez0S7CwC2W4KPW7GPcZ5
gCsvAyc1aiK32fRb9yJUBaOIX+1jgLBxQliHKh+jhm33DvpbKpyAwO50b4h1OtUmEeHYQTOfWliR
VkWzHEve+EMyS+o66QFeK6KqhQ7Q5EEz9Wettl533CKj912SY3pYfQjjZwDpFUJu3lkagP05ipIW
e21/QPrsS9y0HOZytgMyrkF8y/2Q9DHoQ8zfLrW5HfmDAXOJqTXnqQAn3UTnv7YojNTxFC2nRPkd
wWj5wEawpJ9Wig31VkI9ptysXfmM183Bf7P8TfaSNGjpTum/tHvluSWzU/rX1qrs/r+mOnHTKQ6l
PUVA8vMCoYY1NRE/0o50IHOphqcHQT0fF9mE8eiILjK6uIE7FSryh68z6UHihg4HfyL/c3JOzUij
HOxV7ORr7tYd4M07sfWEHrSfvUc+nNzDiguiqmNJcPPMA+T6WEiYVnPDQxBwIqB/NWuGCzhOpDhA
ZML0Rfc7xKM+GX7cdjslfJZH+Q4d2EeBfEtrbAQr2EN8X2wXIdognGZlEwBgBlTmVTavz8TOEvSW
0YdqarcIEFYOYKk9x9ccggfN5HYYNr3FjZtvpSXxUU1xVP1op6rme/ZXyHlBGeH3iJlnpRADv5j4
HzVEGYaXCLvFeGFxVOnH15m/+BdKcIeuFweToHP/jh1G3DiJKNr6YEGXZuCyZUQOxUi76GTZ5FKA
yJlCvjTjKmBBtgBae/vySYqJGTBQ5hvRgKt+0u5R8D6F+Cw0M5GoMO6ppLMoFuVs146DVKxb0gS0
N/ga+9oXfuZU2sxCCAwV+W0b88F1GaXnNY2KBTQIes3p5UYRPBoHExMlrb97TOY+xyKshx2ER2f2
tIvHpF1gyC3vdtdzJhcV5nomo3xke3s1sePb7gIdHagAS6j+Lhqf++c7zn2hLRjDZq7ZOHdX8aNw
CzvSzF8JwjPN38C9ISpBTC2G0jArTCg7xPmilr5IzKwqkz3VBywEb6Xy174qjdJl5PtivLbJ1h5+
pUMeF0z29nbf6dJgQarjewoqXVj6lKc617ShZwUgghtti/TXlq2zlhK5SM3ZC4rNPTpYR9x4qlDK
/odEIXkeppEDiELpcua4me0EVZUAubeWFr106hX7KXRDn7whB10SJOh77dwfXg80ylgtY452Rybv
3KsPzUqL3/ZpGpVPkE1VIk15hT8DIisjV89hvYF6VUJjjoXYHu8ZVBqIDUngKueC3xRw0JrerscX
GNJncwd/Zo+s4JuTwGG67slcLFpg17HsfXVkZjucXJYPkK95PuXdATUj4iXvugFJnPDyp6zA479S
vwUJs1dm+LeyLPKa2jQ0nnkjQYvCJmvYZ2LU8MMSz4f2MDFaMmVks00CkHPnLQEeEAos45CZMifK
xlZkksjRLFGT4UFYopqTPEW+O0zH8IDkEyHNOvYNh+1WVokQ5k53SFm3r/TaL7KonxosZ/EPz+70
Sh+W9YULGEm6k4/quMAhGmLjRYlquyWryHDExyFTZXX11aPgI+msTxORi/275dpU4OIzViQIkurX
Bme0SPUU1+g9dM2ZVbqeEvNNv+6zkOwJwjSCIbKnu8V0qNFM/9T5HjPQ1LHeUAzTHi5QAJIgEFir
eQgsiAxaeYNaIzb0/+ePXKTfCNBRwkiqHVXOjKWyy/s1E+wdMxF+JgFaPypw7s5dmOirqorsLLMs
tAptUHVROcgMFDf61Xd1pwXSiTqfCrSOY1TDCvJD2u8ui0SBT91zBH3LS7pzuKrzKLNNjsdlMf8V
ao4KKYk4O8wAaDTcbUtnQXcO7WvG7ZFGoL9WGHr2/VlLUs83mIK93xMNJJ85o+/njvZ4EM+lu6PB
kkh0MB61MpDm82QGhYsCIKift1qFrpsg0kiwUJVRcwlQmQ7vyv71xoAkS2q71D6TzzPRTwfvRiia
/f8mrTKzQ/erdwVfFcQV9B/3TMoitOwu33leB7QPmQU1ySsvnCYhh7o4Ro93B/aClXcrUdS8pkWB
jbTAosriZ1Wmu1AHdYcWBQdFhNOwlRCFVulchk5GtqPbPlWVA7+b4HP/ZlgTz722fvg3QyqjDzwx
u3680itjcjppa3vKGXG74IEVH2eoShqP0Jya5d0JFJt+P4K/+pRmx0RjzOTFWXFnaKBFsF2IdJg3
NZ8x6GAXBGRcjFTdc9yl+kx11k7CeEFthZ1As2K1EMv07x/4xowlnvyyNZMeWlZ54ioX2x7kvHYL
bgmjvW24pdBI+b3ydGWSbqYrHg/R+bpk4gGSuZBID6o8IosHVHFbKwYSf/HZoXL42sdLhbcE1y3B
CtfLvVlOfbjPQ6pbmkjl9pEfGj1hs7gyqMz8zpJYJ5SM5jaQvJx2bzWo9FWH5Gwf4h3T7Du4Zi72
ij+wK3cxqCmkjM/FGfS5FHWEXnWnTXqRnYFLHy0PnP97lolYkkUP+cxhSba3BSsgi6pM9cAHh4Y5
4it27hMCIyYybdL5ps8KyqHJvWbgHsN62slqfdwW67dwGOlVSxcRccrromxXjkkqXU9NwQCWB5Js
4pR7tXedw3UvHInKdoaEgBAE0TZvcF5IE4AW8vwWLRIyVXIhYmJv2U2tvWCLQ3F0O/3Q40Lny1ei
f94esADuBEAqdSyNXneC0Cg64pfGJXwaq3+XkzCM/qlkL8jDNtObVQDrAj39NoByPI1jBdvjKuyu
Zg/w3oIL2gqX7uemqcXqEy/N7rEFMaWBLMCuspEY2VYrwI1z4QM9jAQo3km/KBGOB4y9PwYEy7vw
LEhM+WXAhcGwQuo5Vh88YGrk/hSQzCE9L1UP66R8VCSMW32TXCkD2Z+dnd3hR4Ek2AXRsXCG4eUO
QsshjDBF31QdASrIV1QaZz/3xbv5R/EpM1+5z8B96S2MpAmwQ4RmRunK6Tj39hTMTntK0Nl2kc3B
JjibzJxyI6BhMMXGi8wJP1gdwLqe4xJQWy+NdIFDeY/cJPHHcfmFaumW46omsvEhb3L9f3gg1uJh
o8DGm0hJ7JsVFEBMnfq5W4jaRcS3NkKV/iNavw1YCI61VNvNzt/B4zpCh6Zn/Ds+LUd4HsXIXOQj
ihTeak8UGD5187HKVdoAqmw5pNGFOJvvjG9P3m/Ou5WLw86Z/3o7Ue5SwcInmP1QJfOx6/uHG4J6
6WcmzB/AW6XI6SLkz5aamaa8QQUIszFlEyPSXHJQObUWmItFyuPb5yzPOkbyxQrzclSUgQCAveJc
nzaIbjvr6r1aXPcHCItzk/ProSxkZmwBylrG8ehGNhcOcUvGS7ATX6t4xpLEyj5jljXwp2xfvGH0
jm8Rgjl+H2qtt0DcrgH2ovL4kA/cvwDtvYUWEB9go2PhJqfPfrc5dhO/VIAETDBjgfAC4iqzlSAD
U8xfWGG/oPV8KFW12h0zA3MScYX7UlNKoUxM4rijOeZi7CKRzEWJsuRKmu/ewDLfvvsagSIWPyQx
KsCNiaDwcCp6AXC5jpkmqMp1GNgEAfJ/jZZisVhYYX5+nxBlaNs4nSx8WmQunNhmRJ3yloN0Kyra
PZQrN/H9+QroSqTjcvUPe1Vm7YqVfb0ZFWOTzhDljuw27VITzLEV58Rz+qm0/w9Rm/RURUnw+Ae6
IhmFXVAOtLGDAqpJ8wSZVEd0pmclc0lmoMp5FLgmrVYdF1bdB5wZjcl2eM2KE/b9dVnwZcUwyloF
Pm//eOvURZ6PQDZlnIpfQMIGOBVGX3ShX8oNbIQ1ZwtODRfQVrwvQY0Ma8eWzWENPenjnglAZY/K
zMcyOlt7XLBsFiRKdR9ffL71AeTNLhLRW9fjIILz8F5hq7H844wijtS4EiiaCJ08C/4r5VbBBi38
v30xvIdPZLDgjgHPK6d629f8dSav0nKevecVoxQJN8bHkJ967afCWkNPcThPqTDAATGHbO3C/neh
gfqbd7f7EWaqT7FTcXLblVpPCR6+2MPrWqQZeXjGmKyE8ASuN76iVNWl4SsVzL/XF5Bha7OtJlvW
sSLRUv++HPuxgcfwqSaeHRuETVVAZ4VY01lWliVl01bBliRXWw/NFfE8idYAP3HdUiJoCJUi/qQZ
CeW7PlrYV9lgnJcXXLB8ZRpb4qTMz/pdwLZvYjwwPPMtzd1ApeH/VcADdrkp84JRhARpl1pMuXOl
9prvX88TP4P1e/PByTy/N//0Zq8WiECBUomf1FkXF4yRuFnIOncGuvF3gx9lTN/dj5PTafBdW6V9
3SqLu/UVQeXc2diI/eL7t8OV1ZSFOcsOEdJ0QuiehsneQRZydDdoGCUPgjbbvhlkP4Aq1pFCAmsz
cQ6Szkvbv72C7wyDIauogrc+9O2jBi1sMW/xKl6TPREoCfOnNpMRRDBiUurVQLR8NeJZuXvC3ljk
QiLKjyUy5BAe6YriLIsWeHCv1nOKSrWzvpHS7Yrioh8zPD4/i6D20/JMsp07ns7MT69QXfBC/iDs
NHwZ7Rpq8eICvViEki7JXGuJEc/V/pX75TaZgBGF7UBcuQmoM9Rb7eXAGMS3cPqLG7gkW/om7KVU
nd/XQH2YNTkSuoMox8566r0/jNFInU+GuOqzdpZ1EjcFVyIMoDM5RVKR0AuGBdmxHZ4ETmHFUAGY
ybEuVDF6xJwogElUkCwRvuqlrYPz06QBhTRNzS/mKtIopcskDsJbj0DkoF9zdwX2KpRGM8Roz2cC
xDv4I8R8GOrQ2ULHoaKLKG2cWEQfihSpDZthL/1ZHsxSkEou2bZxgeofwxLZ/xVYB+tlp/ir1ysa
MqITWvSmEXmvYdSkgn406iIiltx7WPdb7fIyHta6n7WrdU6ffz3FGyOOlWmoLdS87vSoVtYfRYBV
+TOxTfS5N+PQszPcYMAGlYbFQsV0uIDV6/A8Z9KN56lyHT+kbZNhFdPtWToz8WBjgjbU9CGP2K1R
/jxDUy3iqs0n2ap5pZKr/ZegnXsRG7fgOIzSa1x0d9JiAH5xY7z3Q3ICgd0sipe59nB7ioLTdm8R
Pjfoa69vxOLwAsO3PGlYh6ht/1FKim00C8Ia2sCL9HTcDzsGlnR7WrOjaH7r78BG5AKM9TsSbnBi
j8oN/DV7r2s1osixNfSFQQqrqKoBIWp7g9+q2txah8VMaV04wgiEb+fkegxxgpqCNLySml6s7yUz
gsxm6jmaPRLXPAdnbXADcQRCPp7prFlxBgr0sLuvkc0w1RPRguLQLzGnvsqGHhBJH6QwrdC99Wxv
H0jLW9ff4lD1a4jpW2KNWk6BYYqc4HoZlSnlSM/qphn8kv+FXP/eJm44L7Kvos66sfJgr4dihV6N
P/WNWOdljquaE2CwybSD2MF5BD7pQzFOOBVGuHzT368F4qOiyOSMOUf8eYZq+WMrkL4q+QIn0Wck
xlSdkRENHuo/qEP+/gFRTheuzcUMWNizBX1ndg5MSplnq0YFp3t2PbNstbIJpAexXu85PoA+PSZJ
0T/BQO58ocpXWQ0LLwvWlLqX12BkNvFp1i0aJfn1z6RyfFdx+wYMQm+NvYVn1W3nBD0MTug7KxqR
pqgs2NWsjjCaUYOWFFqm9xcThxJ4b+KsXJEwuCmLFG+twxSGMSx49Mlw/6AHcKjrW+bQwqIROxSW
FFpMk5NeJgI8oaWb7EhZJRJW+L2F4Y2nfpIP68XVZI2QEd0HRD4krsbcvY+XxeuVFBgdIpNXVC7U
LEYt+z9MqCiYfokJyCOfily5KzTkolHrdWrHsyiekMaqJ5sWSETQMEEGL8Tvyek7L0bXbDtFgRZE
se1WkWH+SCX0JzRXn1OcTuGT2+zTlQZZBrM6UjWdIULpUoqCaiTHi78nefIfNZNkZBOvauzosDRs
/OlJgi+ioUykTlYEokWENOi8LgAXnStlDvCVrIo+xsS5fsM/qvg+J6c0zq74UTS8SgxRyvHfrcWh
RcnQoOQ16aUzS05+CS4DjoTbZWJbFdVEFblyWZJB9OclH/jd1v5jW/wyiKq5hpJSsqC/PfkR6nQ+
Wfg0tKtwSHUqaS7DtmPKltHVOtwYvYvoiRfLG6do9nkiYsA2da2C8LdF/EQM7sSsPvFt3C6r1nbk
uDHSnkQxFQ0Cu7vennlUKNU0MeFvRomZ47EftPT4OahKG684UWCKgqe0wiJcd5PJLkBC2TP6tbjD
TUxOiv2N6OP76/QWG5J+9WHPuQ7FFxrpCYAE503iL2C6diLKq+tihx4NORkV0JgDV3JHq6lvUM+s
ieGLwEtbFEbuiIV0OpUFDdX9llFONIW7Zk6shJnKQAzdqS+Q7S3cxJIj9t2mNtGEEAYOuLpeG++J
bvr9cljRSdbw++KmQgVdGGVqZBJrokpB3j4wUr9o5jzxw6zsaWgJ6jAlXRfb8xLOUyTJ2iyzQEoH
dwl2CnPJZRw2TKtFJ8VoR9t0Slwc/6+0iPCjBWVTsjBrhgwyVcvXmPsqxKV2W0LNluaflNDT18vF
tGPBGGq3mqa+qmhARzp9uyclg3dncKv8XU8eyXec/q1XLtVTM2bFfcmcyrl3zGy6fTJXeV0/NtRW
W1z0zVbtDoaUAUqwJaLadyRePQ8ZfPaYNNq67HgeB4Hw8K/7DsI7Bfr7oPs19aHQLDK/b0EioM6o
G1pV93hPiexRqjG5Ts3Eur+a+H3RyOv2sBZcF/VTYK+Ee/JBS92Ncd+WLqhOZPFzRdqDe6gR8z3+
RwZi796tG7EnJR1CYEYxmGTmBRPaK70ykKHaKtn6MW/+keDAeOC7Xa8U8fX+J+/jd5YdDvqpAmd+
tMRK220BAtmhotaGI3KSria38odA3JcnmXmQ+fpRRabApJTzr2oPI63S6l2U2X4wG75j64JUIW2c
11I0Ja2ZTseYBfFN04WSOvZFMOaUVNE+xiuvceSLTRdqADqQvO7y6UP9l9XUUGHU7JRbV/U2fXKT
1zbLR7h4mzq24mngBQf6kqCO8ximEHcoD0aSaCtp3CtAVD6PaB9VzcCTEPXPRoz2EJttMLLhdBXH
G19c+fIBFBSl4U+KXdU6pnt+ggEJjiADSo6eECbqauRufd1qVxaXEirC7TeDGMtMSqnbupKD9g8J
Q6KTnSppD0oYJPudL0K3qdX9XjqGMves/unJ6kDnhP34smj3T/LzFlVKHxUq+ySMFkTgyUawPOJ8
48W03G2DAFRGl+HjWqi6yxOrAnVPCxWnksAYRQin4f8b4TvL66a5VR/xbQTjq0dBUR//tizQ1qqa
0F84DVjmsUekE+EEld3z5Q2/+iNCPQ5R7xuNSZBYavfRKIfO5jfLSXtKHWJjb0GNwd52aVRX9Xsg
ppdlur+OF8vAov6QsF74/kRrETxw33a1WEgitcniuqpIOVn+xkn8czBsnDmqdRxMEx0LXpZsJhBk
/10IUKAiNAMnGrh4jJg3JIAhjKTEklkajVFLAUEqecS4Pj17w2rMqO/fMcCYVjgx7hDU9FSIdNCt
3DqNpg3gdQNkHCTy7at5sKN2TMEIb2izdJPtUOqKvFQ1i3EjsUDUlhHWUN4R3j9lWCKeQjSufWhi
KCxtAcD0eKLWu/Zdv1lMtVxS2U6CguYipel12B+3huS0MSxcUp2stoGhYKPpV/u3OxcI9mk4hRHe
oUA1BMM6vumZSjMK1KTLIdeoG5cU2DSTvBWT9tLu0L1ehMj2rDllfMV45jKlA9mJFlQ1LLXmE4zM
j5TJUj9eyzhBWlqMMBjKGeKekSi3ZiDtQQN5PK9uvf1WpVQnC/cTxRzz28A07m2oqxrgmPzF/o7S
jg+Co4zouNyQDK/17uZ3/kdJYC6n60bOmtUXhMJvVfmTCjFEHd6rywMFe/GZ8HwqZm8M6gWNNrhd
ksJ31YhZJhucMrMMro3osgRRat13hr57LgXiKmv2kKTK4yseZQnSbYfmSEHBRxOYovnrDaTu9yuq
/+lyYvV34GJ6udwKmQ9nqCdCI7psp0PXE3wyT0AwJkl2kQKmlAX60Rhia3/K95t1TmLIinfXaCpT
+zow0R8Mqbnxfy4Hiq+cjQiWSq5LRCB5yq1Z2DUeozRqmEdGXIuN9ZuxHZ9J2ZgtF/xE//OaDMZf
f8DduiSN1IN3xZyYAImFCiyuriZha1u+psiUPUo/jTMk1It4F7XPZfI1RSrvf3oHZRPURU5ppTcW
O3GV24nSDwMgUp7J1sWmWTLeRje1rQMTywAdPvCy7XwD579L97LVNdJfA2oQSjTnz3+tJdJIKhU/
Ji9m3aEzx/sup7HiRFSx+AyYxtNMorJ1essZvxDIg6pKBJPBhfNOlBjNN6DRTHUJBlKLp1tBmEKz
M5PyjgnO9d1CBBoObWYNzflQyeVcjlFwiPMwHCj80HIT3RQl4i9MuJt9mEOxeQUZqrPgOn4ZNguz
DM38RjcsE0XwT4aXJfdwz2k2BPvfrWMuwHLwG6y6y5ZljjHDjK9PwVRLyUEqA2FwtyptTsMKPAu7
DDGgI1eO9qfuu8+VtFd8KoSLopNfxwXwwk5NvX8Q+ioiPcbsZKK/6KrR6EfLx9p72KqqKcxxu6YX
iOO4qSAdX4g+6eRdeEbn8sU7ad805myQ4HhizrzBgA63ldFvtOjm0mJz5aEn1AUhP8GEl1xkuGE9
tWPIeySJspK062Lgz4wSaaFzLPdYANlQE2vY1Ti/sMQpP2yE9FQS979ISe1HU4SZMQOuMLQbZh7o
Bn8xqlVYHnGiXLB8ShtWAM4G4Oc9DH8d9ep1lyQeEPDmr3aOVostAlQm74K3CQ4BrHRFNEd/3XTG
w4mcNXYfZrp26wUEkfJctr3ynu5aXgCwbocu0ZRLIDBmtdKRBikZefcD9BB+G0E36rSCuDohZms2
o4IpAX4Ku0PHOECZ5SunI9NSrs17SDZq9WZISOHegv8bKsenjaGqdF356/UK9xrdn+cGWNj3g6/L
bMjzOHDMxA5GwZ4Opb2F87wpe4yp0kBY+Qbow57AZpIQPyjSX6ojQEWqWHPgarFQdQu8hpFIEE8K
ZRLsUzO63GC95VRUCP81c6v9RYsajqAbHiXO9tehcc+6KIhQBBwLHYxT50LJtd3BNBAhQ/tMgo+j
p3gkgb5mWOAEFLAxl2dTZ7KMwmO+OWkKJt8p0FHQ6eDnDabk/Nyy52k4dNVQ3ZLo0R64lorIY120
z3XNXeIICEmwd2lO/VYChSowt9dEKwzlilCdBLjJ+8n1r7HInVoBY+V5JjoaackReBtxsusx5dLq
5bx7p6Dr5nqhvkNuEnUuHvRnJjop3K/ddAeqGudiFcyWtJI8CIc5JRA+j3GoXMG7qDLYnR4GTcrr
ystpVxx/b801ceLPoLRFS2hxj644B+uwXlwtkEZ2G7JAIAdXhWXIvKdOiuN/OCt4DrmuwebxiqpV
nJ3doZR7+uE0PJjtCifAOvK+WlDIqPt/TKQA6ss3mffy9AD4A8+0dADbXoyPkQJrdpQ55aMfUV+K
h//sXpmBfNpCqHmk993G7VnqkMl95JVrH8sLzmJhOUU4s6TXsYyTw2T4x1iCXQNXZrPIhG++ZTHH
+AW5PlQtZXZzPGVYf013PxQpImDZ6DjwfplY9KtLFVOtpIUgrHLlubUJ7yD1gqZKQVQMWZQukVyo
n2WalXLnW3sgdvsm3sPPfgx3CMQASsjx+YzxGH7dDY3I2U7ESM+inZ1tyh0uE3Gv6femUIhXMSSf
YxwJ9rFm76TZVckeO6GihTqU206CQOfIoA4XwhpsLFQD1kF2G8r5dlFSxV4EbLHNatkJw1QxVZv0
OgJZeIReIfknXsc7CqtYiR+J0Mzo7TBWK9AZDbeR/FPQHGP8Cqss1vzhdZjmJ0WBYhCGUmYLCsko
8r83QU8ksUmLEXcVBNJNCCMA0JyzaUjhc53VTtWt8PtsVvLQLlORDbonXGZLS+bKp3ut7vDsjs9g
TAXm9RDGUqd4CNMg4STiogpoTJJSoq2lcspcPA+QceZKu0BPITNHNEu8vbUJD6R8gZorB5wiP41K
IlQhLfGkAvcyranw0/borUmGVqUbBEfkWGMI7wgajHQQVf9pU9q6iXGcTHmAoLFxp30hCwIxmLQV
bD5DtlFWrPo6dW6RJtfc78qcYtogEALL/Q+906UD4fVmmCfxO63q9vcL2JHg4+ZbOObFYlLajW7h
I+Fb3m6MbySf66PBTiCi3OcC6lW16rXwt2biKohklWWhvet2LmZ/NVJA10tCQPhl3JHG6ZKn1AzB
Fvgt4ZGx+Yt4o5s5QLln5Y4AYEzLq+VC/BGksIn/Y17qtBgxGPfMleH57e9lXoMjXnDuSJQLOiLq
utGnWx0SyLWP3rbreo+MwRXhbHUjj8ssTXlMY15xH60PCzpPmn6x6fWj5YIyQuWkObv+bgur1AJo
4TDUNP5zHI2buDt+CCU5PnDT+sGZQSnp36VsrqaONlLFW1zSAHFiGo+nhCRjVyMrTJbCqL0VWGgm
ENLkrWFbrGxngeQsyAtgAMEzJjaLFk02wUHIpLCpNwT0r7ypuumuORFZjGBpAaSx57llaY0jE52J
MIl745l/F9sW2aoaYRvjnM91/TCrL467Cz9T+Dtfa4eHIQB3cQTwVui62+wYBPXqsW6e2D1fbKnU
Y+8Ssm8Z+3YjrcBEbtHuCNSckn7cp2VfVe7GQwc11I+Uu/8vxVqIVlOXQj60LhwdsOtS0wmOf/9A
BHcKe2I8+ComnZz60LuD2cLti0+XGY6cwDwVPS0TQ+Hjo9g9Ko6c2Q1IPjlaP1IAtFIQQKDlRQL8
5fUS3avEJeJgsUaL7z2EANz20VaH4LLL/XKEDCm8mdrNLdvOYq0DPWO8SqJN7X98WgWWu9TRvG8I
OjpMU3pFWlbHwM2Vc04dBGjeZCUoty6WdaeXFlQXry9zorvdzqK8tLC20YfMpt95iX4f0QSUh+Hx
pgtCw5hndNCTgaI3CrjzT29JwxtkN8H52jsgfbswolC65m2fuFXBqyd9JsFWOU458uiM03sBLFKN
qyUJlTjuk23THP7+6Czl5zaOEwVTVyt7qd3XFJWd5MwbgxtQWNL6aKnYcUOFcpAHDNiU4cyDp7Sc
efYfTNvUuJ9V7RSvz6afzSIV65LhTRcq6Y/HsQde3nNyUvpbbjYEAVCo3MXMExuB6fXjhfJ5hD5v
cLkDq4+BQnkoM8tFnqAsoxJT0HYk9zhFa2WU/0+qShnKXOndhGHSP6kaA3QObUD9COhQNgCQt48/
9bxN+TO89HI4oKx9SDjR1BtM1BnkPFO9MWk/74DwpOTpfKB6BFyrIolU74QkgJdqD8SSALyzTqmo
icEN4ukDdBg5FNrADjNswJZk5qpcIojGDFTii1F2gKA+hohHWS5E27Rce/dfXllzT0C5rzZpuB+7
6E3YS2tLN4sOMnu3ahyyrRQACxF9hmKrWW+ioQaTiiq8KzaxatF+Ug4vGr5jqBsPOVxeNjtIeb/I
32l/pvf3Jkw8fl4FfYRmdE2ni7zotXrCCTlIFgstrcqHcy+0vGog3H/HYGpYhW5wPjJoCJygeveP
QjxTHaLGJqJIPPuVa1UCXNKoABMzbxe+zL2B8hTeYV+vZI5fwZL9WPAc+vFlFqG8ixoQfi7FnuYS
lR5bPoUlpRJuD49me9GaZwAb1oPBEvZYysBMjazeKD3DlUBjlahNcyUIM3BUtre6wsqOKeln23bB
e34+Kjvf3VuHPnDPoFWImaz7Pk0FSKxVbjCty3BQguzmwHbNUPsSU/RqZyfAvacK61QtlsUoMIAd
vYiwiSghVlowfMKqYW+CRImhozbnYDujVmpINkfYyuHwZHwW92TJzb4hbbjjKZM+YJgh608pSH6g
rkuq0IspLhLyXb7PBAG/7bvavl09mAnuqQRmMsafLjeJ+v8tmtNSLE3aNxrKfZIp3M679sQfiGn8
44eXW87gmaCYCAbpHCqvZ5ipo9jpV8abrtoR6O/byMBNmgiPVNr8u1vsH837lBvoCHhOJLpf2ooU
DWlYawgvyrrQ8EkTunyrGXe6q0tE+rUyCa9L9ynyq/z1HO8eMgNJootpD2Qi/RsJ0rGcvL/spoI2
zoGZKvKJ6/pCg+sWHqzAeLHVuAPdC2Wcn0BfmLisnA15JNNcA2uwLl5vrDYLL8g9E4fFpa44Lv/b
3Ruhi+XpXrzFaKGPNXU4W2diLkCATq1LvrEVb716DuLBRXDrQ59Um9e7YeNcb8Y43kYDfpFDgULO
cdW7INNqiTns6ef3MX+03DhqrM19SBWeqsOH4srMTCA9hB8VJiBPTzDTxQ3D9CZMt+0jvIRL1cRH
e0yH5s71iKvA8DfjywAsdVRzpSfVfMtCdw0laLS2odXQSp56aeHxbS6qlcceSA7nkIZLnn0G1TKx
5ecgV7b7z5lTMEhYnAiGc570hq8ZfJGoB2kQ3kt/a0kwuLdGr1GVEJFjwbmFNhjvlEkE4xdnuLhL
yYgNmDe0nqe+o5qPvffNilYvYAvrRDwj1lsfCajdgfs+36/AwVOBc3NGF3tUK3XVbiOYk7DwvzwQ
C1qgnFTX4m5h9QhNnr8LBqQU9+De8Ju0+SA4FtcBiqi8KxI2A2ZJVglLSgbv5uw0C/KX+k9ar1X2
G7u8vNDNvYRSYyM8GubxzgIf4OHxxpwEpYiupJpsYht7uxH/YnG1z1eOtF9/XO7Z0Ss0dj9INTqz
GZLGQX9Siq7NEhZVQ42ccR7/+Ypw8JBq7RVCE2AfgrotuIsSw1AjonkO4l6VahOYZxYE76NGUVzr
hYMZrlGqWhUOsxylB2ee3QfkStE/tT0cEGn9NoVcPEUwitbN7RQ9ijKUd0rI/7V5QGGkoQpEsg2U
POYYdRJDn89K11yNabvBwe5jTDQtLkCeqNxAkJnDk932wM1VN+iLNJ2NoizquEOpyV/2s/Cv+t7B
xIgcY7+Zr7krZy9dNEgVo5aAp3hwTbHXPTnWaHJOqbeDqmWiNP9GwO9f6oIbW7HBC9+vbjV6/1F/
148Qa16OJ/Fb0sBcD4CGd2qg8eHrDAet5y0elo1mKU3N/BagTjspJUm4bXNgYPKcfBf2ngjGm6m7
26zYDFwl5Uk3a0kM3AZnuCgbyFuoM1hp15zDeevf9xfT3PWmgbrogpsvQg0B9ZTSTx3ZnWpddmol
s27z2Iz2H9Nec8O9NHKoyAg9yG2bx/ESLnkgKJhl77mtUgQi424mKfXEH+IfvJrnZ0JeJLPIDPO4
KM2et6CLoCodeNA1HsvNSKPn86tiuQRCntyvNnQdkV5L1rB7iJmjZJf3I3ZEuEsCEbW/NnT+Bdrz
FAs5KxxeziTP1ylWh26SPsLOSqQ1pnrosOj1+KhP6Bo4MrbvXHoZZqspWBFQ9/D1OpUih1VSoup0
b0WTwTBmYiioQzSX+gTVPF7NZKxHsze9GloM/y/i+6XsVTXpOTMz4KBBAPu/ZVe8yL+4++2dqTq2
XUyGW1m3joyeOGeRNhxAjFEW348k+ZYah3oIPuWLLeScfHJGWmx7cJMsMhmMFZ1jZ9k1rh5uV2gz
K5WUm1tYFp9PipIBbwJLGgJFUFloq073geNZWbqvapSD0VrX/v9x7b+W0PhPcsecZRLrafR1SQxJ
wX6TKqTbf5NLal5FYqx1E6OIOaLZsb/hk5sMQf6sHIHzh9NasUYbrWIfb++RsPttrhT9XCZFau5R
vQIEXsgfE8y5vXeo0GoPgmwgtTfp6dTO1EBDRsNEq3dKXDwUTglhMNapj5R/a1sfWLX2HeuTnC4H
wzy+p3l4LiMaOkfSe6Ox8B/oSpdE1CgsPRqE8u+cexMWbg73vTlAd6howuOAJsc3Fcu0lGqMY9pq
wZ0iLuKzOQM0sRIKgMA1DBtoEP5/Njq8ctLAVIPDsT/DyfYQK5JWn66dmnueGQ2ABuKgii8YGsrh
i8aXUO/2Qitf+SewIpNJrbtlbPDiFXskUNj73IH4JcsNvophmezZaCEJ4zzwLM+si8cLWTx4rJ5C
Vd7NTq8TBEs8S97pfSxP7JKwDFLedJ0hODA7ZB7CAhCTrN1u952cdnI4mSi3I6z8Dax1bnksUoDM
J/YMFHc2X+EGjyBn7HvRzp45P1CDQ8sbPdMF9XSmktgFQBCD+tSE08GvnDUC7Zc/ykqmZfnQ5g+B
IqZCG6PQQgcw3MoHvH3x++st7zw3T6E4rBHJLVliEsxHuFaf5lLb1PsoJlXsZzgN0ZbFBOPxiE4k
DH5EFdfY04gTcnEOaj3MCSQE+5O7BRlSdapQx2I/ABKVmnVDnoAqMiWfnraL7FUJ6g2oA4QSecbV
ThJbN/x2g55iUetIrv2lbcpF0h+c9CpdsDqeH8wVuolPPKLywRXftMClVNbm22EfYRQHL4Dce5rQ
vlBZZkV1omBgfupnI/JkBEXm/qRwceSf/snEEC+SKzW7V5D9rzW6TG/F5LBA79SC46BodKKJ5yc4
U0xbO3jR2ekfcllfHJWYF0ikGcoQ1oVQgHmW/Msc41cyRcxNCFDXUOiYXhD38+1AGCnpFtuRo3lf
9KvKv9zH+N6XdT/nY9H9aQzcHorNjdeVjlc9VbkZlx2tZjZO+WjpuN68YrwEDqevjHG6KmzKDDiR
Cvt7KxjBHR//Utfds0iFmJrmsNEcDZQR33a0FOhywxdLFH6zko4kkY2rI3pZuyk0WoO6GkpBY4nt
juluz2zlOQMhrmvKkATGaaj6jyLNd57FGLgdIp5jpMVbYlqgCOPgxOOoe6zUopHVSvBR68PU+jz3
hIC7mm4WP5suP4WgtPqjeKvhZ5KoPKbjKjqAJ0RfmlObR9gfRmLcaQ/nNgsv78y0w8gXt8KgYfub
6fxv1P1+CKAnIqWaxhmhIrHgSbLlku/yjC4MmnqUrqQYqQsAq0QXRdOcfmZtSHpCFtvei341BQRV
RTWhW6KTPtWO1hyjdnhGcintSP6Nw2OdePKNqsJj/sVy+xUCLrlXHLR0/kraNMfOaRb0Tpr4UWIY
XMSzhmHMIrQFpLuMqwE7WaQrjZXRPeF68T8t9CdSFoTQZzmuSXQvkvZZ80KN037j/comNqH8fTAU
Xgo0I4d1b9hAGmUnENogYgJjdsZyZ5q9oBwLhotpLlS3rnw8ZgWA99CH8irju4yk6w2tJkbTvFPJ
qKu0nj9RMsZzNaJ0WoDVdBY1pQbl7z+2OxXMZMdCRwM3TvuGwcvbR5GeToAscXjhozhiLp2cXsTw
EghOTV7om8HfCt+9Zqmz6CwSx7fjHgjZBRkXfMNQGL5BZTJH0vjM+iJZFJUa0HAqCek8avMnt1BO
flTM+TRjgs4v95BV2Hzldee+V2TIzpo69sS9wWIk7l3WiAm3HnmNrwpCMIT0y1M+Qbnf98fWqAG/
7DQr/g1qwWaFff9NansFaT17G0sU52j4AvRTfxFjLZm0+zTbFXuWsZzkyfACo5W9fzZ+L6VWxvPR
vrA2TyRGXE93fHGzFSOX/2Zul3pV0v++Ej/aDd4D1e5nhk5LggSMcVSGT0wGpQGqICq9ueUT5ieM
OL+EHPNERkRBHNgLqDRjXglfOkKOEFXkdtaR8XPgHvWgIvQtLsUStduUo6g1Akfvx5MrNjv/6Fp+
XjUIQOYVIZG9TJpIPY5cr6ixhdMq9Nwp737ayGfgu6g4NzSSp0m65LLo3Y38mU/BgqLRlOeWkAfQ
deIvqAwa2N2R8xcnw/E1E7z3sDauK2QPsZHv7T5a6xYWQxeLQz9WxGgBwXzSBP1vuKN6D5WqPu80
kRVDTb7IlUBfgTXyOmWTXT8ZHy2YPsAjAuhKzlFFTvvYFWasJpw6Mmsb0fe+8MuZ/qytx/OmNheE
WGrf7bL2RKp5PzmRII9nAnDebz9AkgN7QAqy4CODO6AapEpiIHTgaIHKyUY0EbizoBTWUNhvw7t9
MJFCg4cVh73n4GEu8X+eLdC8G5cvrEVTPkfuhcRto8HsDzaHeIqgKBsiAql7pmq3AqhouuxQ2mgL
mUvJIi/3GPbwlxiaOXvHFcZxi53HeHiOMhaoFl5RA+IPgmSiLtHH9Enh7H6Fu4WKg0r6EYdYSLlZ
1SX8kQKmWcQhwAhPehTLQ7q2ltqi1fkyAzniqT1TyDv156VYWktjtkt9ZyTtJYT0vfHyWeM+nOZL
fla/CsEXgcVezKrFW/qlsBfOCTGzYTiHfYiEplDCYhLB+Q+81EQ1m0V4xIaAVOApkZrDI10o5ftU
cFkrPxpHx1EWp1cVikjcyreafzSmrSmZNa1YdLLKSfqICM+5/O0ZrbgnUpAj2qmvreLQsDNdv9g3
DC1U8Zw0tLsZd9GcueR9wEEdbdA99TsnMbh/jfgEAHbJV2OSX5LpN2SyrsosTQbdwrp94bnmp1tW
o36INQclCdnrs52tX0qWsjqkcEen822Lhx9zf6uqFYxLL9T4//N3FHxkF6Ac3pDoZtYFiySEMDCo
TqmRdaesD/+7fgSI2QPN4NUfDzj04t9HIingttp+845VXW139OMZGV045IvK0xkU3EV0SnopYRXM
wrQBoczDJsrGzL5d9jiXOfZksTMQ3yFeCs5TUdLGDzOCXho6iGlun3kiQpLzJPin4KXpBqULzyub
l4pJkVPIAMboPlYLDyU9KhZ1TsWM161qdeWOXhD/wUVG6bcaE0BmWJ8ZRpCcV1sxDDFHBz3IL/Sd
A0GbydLvA3xmL1DLb/38GKV1PpxuWcm0NoXhpfw3AQhjHF+Y8L4yER3TLihaqCGDhb6TYIVSCGED
noWUaBrAGpaz6jGRy1keJptmWvhi3R3XYw7Rex2M+51EDsTRo8fAOP6rNN18oNQN7avjHfupgWki
s3MUe/wbby5bf1DBSh4UdltYCteM7H3/xBm41XgMMylwzukm2anVghWnDFfal6VkwrR1mp1l/iOj
QiJADwIbCg4FU0sEg9XbkOxQ+sm88SpXvbUgIN6KB+h1CuHtJGk5FFCos0OFT1X0z1X2KhXanojD
ZYGLx7LolavJ8wynjL4oMmydKHsmylP57rsNtKlQKI3vPG81KASxqfIl+GrLpO7P121bzG2UfsDX
jgY7nCFGFmtFxqaL4m+q8Zl1PzyGxdZUsYZW7xvybxNI3KTujTcTcztNAGqYP3f6iW5tT8o6ltkW
3B7j8bU1QLZYhQBJu9EMjt9zBHeqNIYXKgVFIoRwwd4Dw33Vvy/6LyFwuh8YztMGUP9jWxFN6ZXF
QZIr/h63v0HNE0osU1nO6y1bc5t2nrdsOw5787w17Hplq4XiQuq+OEFgp1Yto5bmjgOexsloiLCK
2IMprI0iTaQNRes45WzhdamlZIvmcK/zpnISkYnFmmAuQeQh+G84xUEeWyRdJ1mWLrtqk6LzDd4Y
TSBbImR05hX1A89foVr26c0AWPfrQGWdX1QgHHNsQ9FzrqTMXRl7waMMJ3YUr1XMTRZI7o1NImEe
0xVhz/iwbrcleideXef87rr6TbzN8AepKJefqUxaZafLYLLB5Rb4XmHa9RqpYYW4pzOD79EzdnQK
qIg33rakW8xahZI9pYXELvZD60Fa7d2ZNNJ3m5CjhEae8GGGrHwqFucJRtx4BeLZqlRbdg+aBEdI
DONB6ZcH0Rhyxh7EGP329eELh3PCu3Y423Km70eKKLaDceFyU3raVd9jOLqAKisGSrjodiCHAaEb
A/yeq0QEESVDRy7esijhk1eZ9GTMXiWSlfbonuAmfZqiltysuoetAbtm1s3qfgeWrD5Te6kjmUTy
XUkULOo608s2J7ECgvfRNZ5+M/uP341+HcVIyalmCGIP8YVssmcK55WnjUosqT8xSeBygdptxlkr
Qpt21WXLj5NND3ZMl3+yLEDX5vXem91MVO9lkZpLEwbUTjLYSQSn8IMGpwwOhmOzqsDeC6uwLQBt
yQ8cleq1YSA6pBkv+rARFxYQeE7+9JVt9ha3FSeaB2ZkeOhsqp7dvmmk7tYr84S8obOJ7t8UL1cq
yL5sFaWqVYhdA7sykB+yfYNygr/scL/4nNPPy6e7oc1ayUkerqkyf1WJaZeUphSlOlJspCBDvscl
4R+OfHBWM78a1ASSMeTNeGRv5vbsEaw1r94WSv/Ks7Pda9Sty0y5TxKmZmOpwDzCp+iipgrQLhJ2
UP+WBS/ot7e+Jk6pndKJiX6l42d1WAE9hmB/FWNl5WvhSuw/QuozApGuZoN3JyKaK5GS2a5w76VO
DpZbPLsqLdaEtPAG1laInILn1pslOHQgyBFo0JsGiuxo1Xfc6nnxdJNdsE6X2RBQh3gAsPH+4hdq
o2PAC1bVWLZreJiLxr0CXL9tqddChtcFvRYxe28b1Hu96eZBP4ISz8VN613FOCeG6X/MG9FApL+7
/2t7JkMLDm2kgFWR6g2WdiqyCoW0lWao5bUwEleo3xid7nUf9pjHDeGQ3n0zk8gmSFzr8UBFOMXi
DSUqjoeQTNFqwFxiUS/RJkZWbT3Ztjq//60TuMbnQmPrrm7ItH3lOZdVtck2yFWfHZ9rb0hnYcgO
91F91AYgTjZJr3DeiBQbSWTgCG9vjUs9jcQtD0OlsWaUOPqbZS1EW34joP03eGkwR73Q7CHMj80f
v2s2rNeR9vT5rqKBTdR14ZE/5KPMd54miuV1XoiWjDA2Coz5RgVQJpSGsbbNAseqlf0eVhvZqdS8
G+0BC/JPkWi7kTQdzJG5Aalx3wXyKoZJ2u7oEj79OKv1DfRKttiUa1cEdFpB5Jw4g1MxYAdkbqjD
N6JtMqAwPXqXpYpgTmj9Qoaa3AkFlHs207B2BH2gqd9RjNHUerrtESf2UdAQGZ2qk+3u1ebEgyD4
jonxDEJMdwu1EMRqd9Lh6Bn3QAU5ZYedUrg1MlQi4x1fXvQr/gHBiNCD22yPiB9lMs+THVJAPKq+
XU5WrSXpO4qnvWR667npqGqehjFAxk8UddQy4cuXxHa6RFR/kyjp/lFqVas8XV9n/VbpOE1seInK
X7sdhXwoPxEtdUoXcAwlccBbnhGwnxm1w2dNMVk6gH6oEeAJO9qkRxBsE4w52uSQLJzMLn/GRfYF
KzHvheLCC6eGBAUk9MTfdKAw9RkQmPPrMUYiigMTHc7UQ7l5k9+LdHlBZZi+3lGvMd6/izUuEW11
bJmZJZ1QW30DwheN7kD2gh3JEIencWr6zzTUr0Ku8DZmlPz1Ut29qsO3oaQL1vXWmp8pP6cPJRQq
lP/PVJkgFHsFgbbqqsC+lqR5T2ZaGOjMVT/wfJ3upauSo0GhKBgYRpMHWVYiwNtXZWZugzE4dt7y
Sm4Rn3pTfFz9BpaJTI+kL/Op9rPWRqSZRfDcNXGz3GDy/0C7tEXZfKouVYw2M7mMAKm/5SbfhWZe
8Zc1a0EGHoeP9tQPc/3z6ymKaZD1KZUFeANYsITEVLNSy5sZLo+O4HwPN2MTWzrB3u0yIUm+/+HB
TbcnRhU+r+qj4EMU1OOPnPDvi2R4DUy5g8fqP3NPBR3qTwilkeL7e8a+K6U+jtvWaWHgsJrzvKTf
mMfVTNOI3uTU1cqByu00yK5j8UeHtswGYoZpN+i7ixvPRfKT36/2h6SQtxtKOTp4VTAC7I/zIOhp
j8vmXmGauH35Fh9224uwzGRjdPDLr07pDoTUirS7C/qLLDHA0vNRkrqJdst7vGMBdLLLA3FD8C+6
znHAlTFTdeAf17XlVi2GpC0o/UbU6SiN+/cpiDtln4EWLx4VTSDKBEKt3TIXgnW/vFag8qiADKHz
e6jMAj2JCloLS7ydxhzwJVgKF8eqFUyHzc2PIcCLLw+Z10BWOLshrIb53idpmdogKGemDE+URnPP
Wobg+C9tCpO0mEsHDdpguc4Bmxc9ChjZG4TL/OJ7EzgpznCL4TJvr0zhBo/NXKjGjcrL7edARNzt
XdxKVCb/AH3Q2P4AoHW9XE3uTPgzuzIj1l2IN4hgBVDcEhdqEl9CMcuclPtnPBFtjdlsbKmyppV/
oKW9SeiUyWfHZh5eKy5000DJv8GiCAUpW1ClIemIkMjPGEyRuApgb3QenBCIIXB6p9YCZMVq6yJO
/crClTv8smWcyE4gjmlk81AQ9+5x/+FixexC9Odj1CJ2dp4z0TYEKhTsZyf8CHRI+Idy6Ttd5hWs
lBXxciFcdfbTujt6XxyGBhaQqC8nOGF+vnxn2bIbSAhjVLNQqWmoERylC7bamfcCGkEnfBPh9Nv3
NU9hMeTkkc8+yoazLWTyNtG6WqlkyjAIz590VYQ0vVcsFM8YbxEp51KMfpOHEZXnvTfWiMhia5/k
tX+sdM4Nlq5XfQPLy7sUrtTedYVFwN9i1lFJeicgvEzs+LiPsms9hpkGzDwcL5uKOKuo/9BAH4mr
UYMEmql0L0ZE4EuB8+A2xsOWdGlg1tslsgmmU9aZkprm4Ng8mYx5isqMu9y8c8Ffz6/ofgXvl5/P
POtZGt389ZnGLaoEBDkAOlTjL/Es/Bri6PGZhejz71pvbDc15v9bViZAW/sJ3Guv8TKJr1G9lZmQ
W6sF36WHmNPRqjHug0QBHFKVj2h7IDUQqL9Q/8jm0Z9QsdVud9px9ftorvdBsJdJfFu4j3F1R0I0
zzQhOypBNS2DQT3Tw/SvSufS7CX443KREyoCeqQmgyy8OGp+MuYY+acq7lxVVN+Tm5SdoAVEZrmw
wRvNDwDjs8rQoyE8U6Dp+FdxZ6QVkxUwVnYDczlvZad5gQ574VkgxfNSIDNiiPnPoSRohVfykjw/
FpO+zH3okvvk8XpVjZIcqfIFYxFuZYluRBiA4R2NSCKM54ZObRwHDCFcw2zsCcwDQ9/XaH6l/iSx
f5VsdTjUD74EB28UhTv+lGvQpp6jxnhToAXklpG8moKap94a0NpBqlB1IzX+uBRShcfDfEFRgTQs
bI1anf1WK8CUMxYxJNA8H3Gv/BBcT57CIShu9ZcGfDHdW+wkycg/0d8QblU1mfdM03N4oimk0kV4
9LSThpuXpY9kdQs8gRV7Tl1MPvamOu7Dk1kApTSDtjHMhyTKIWCy/axVO4vUSkKU/Y0TCTqiCUO1
5e6uiE5e89IjR9XPahhNHOTyHlFAs2Fz7lfbnMtBe5heTMT/azl3wCRW+Bd3hZyj16grASt0nwIs
hTVKn2Y9syB/sKvojSZlmg8aq9WgLEQAaRVl4HwFn+1ea+jkqpDBJ/x8vwP4tEGPbc79LuOe9BJ7
XgFijITm9qSzTIPwfsZ033v84EmtlBuce+XDP1JQGlCNvCRFnKftpxmYwZ8v4vI/h0dmx7poL9Y2
ZFxXaWiOYAAjXg1nPBcgPoqavEC4I+QlBTAvmpuBhPnU6273xH1f1MckoCnHA0Zu16wypHnXdwm7
pDKImxrjxj1dY93SNnyeJXuMrnBDRoM+8scMG3qxF+wJBcLEOE73Pkj3UxVDKhEJEUi+w8+lqZY3
eRig8iNTfaRDnlPSE2gnuLgTPBKPYgGAs+393+e9+5n0l4ro6hQyoC8iDU7gWIf3aW0fL2n4xzpt
o3mbhT8lg1mJXMrfMD5AUjXEkGfKiH1qsDawK55dCQfZaZebW1VaRiHgNEHL7HoRRdt3dWlwpvCU
ccVKZaFb7a2ONo5OvR0W2YFvvHmd62v/mWTdo5wDR/rpN+ST8Mu8PdUzIEW8DydO3mJmCZWqv2ZD
NFosdFfkyk2hY5F4YY7HtW/FRF+lbZsSCNp/Ej3bOqL9ygF3XE9BPf4XZ3m5FYeMvsafRyJ4Kz10
Q1SC8JL7ujGFs1BgG+Fa0+t2EEN8QtUnqvAQYHGHattFDTnzrP/YLxtFxO7Pd3CZqw+ivJD7OXEc
Emi/f8PH4ZSJzmEIp6Vj6Ox6P5uR6d5O6MGuCCFVDvqJ6TUjB8SO7Fm7wEYoDdW5CU3u5n22L1hd
TZpS0IH1T7AtxUyGDhUsE0hTDQt4Ljma9spsD9jwxCwtPXjkAoR70Gh1lrw2N9C8x6YnO//BX2m2
+IVvbKJFoHmx6ncw3j1LHtr/9psIoGCYrKPFVFL8svFoylDNWl6y53WxAnss27ZcsAtupkz65Z3L
uNRa9z3aN7wGnSoeiwX09wPqf5PVmgQ/lr9DUxSsKMi5HjfyB3f79XyDwKDZea/RaRQ6G225d6Xo
1GbeBBazn05/kz4mLm0ocm3l9yCp1AprOr8gZHR4OFDDvXcpdlPnd1XdPiK3OcG4mYBBW+15o3Ag
/VqlzeHilxesEInYoalG56V0wLc2C/Okv/hE0IIPAd4qAxmV0R6+AvLkVsM5dUwlEdDFd4+lkcJP
1iiz9VCrtQP+wrWSv3c2v7dcGf2K/SfN7U3Qx87OW+yyI/GfSnNKMd48VWnnGRaSzaShz/Ti22bn
NOLl9vU5kYblcRxHxJjtBTzkQtWF3mjyvPvxbl8NV2uWiyHn2gzn+DX8WlS4/Nh/kwZyb1uIBIM2
Qas1AaAvkWCAYzIWrLZKzi5L6fIiT8zFmQElZM4EZM7wjPB/yvHadRQVaKm+YKqgOG/hH4/XrXcH
hHn644c5d/khCuVFBYUF64pn5oK/aFUeCa0G/A3OywP+8fQccMou6IlE7lochd5pAj3JJBVeN5Sj
crQ3U/5rZ7ByfEh+OiZ4HvtPdbPFOIT+AXWgcA3Fe1RO3N/vtFRI4CPQTxGukzTkeKlmhzYzucAx
gQq//7W3//4iJs71YtRJZAqOgFAvUvs+1QF0wylOo56OFhH9rJx/G1nNbEp2t6zXv1iCnDtmZonB
pMfczdUP+dahHSQNfiaGMPzl0hEFmsR2XOPC44Xv8xtYAbpcOkygG/qa2Ubjbx2M5E/wYC0DFwPX
wd4xjoBLl+/vyO3jOoOFCjR+liPuV4fARJLUiuhN03oyBsqsiVsGP01OVCASMJQIlX31fox1rQtZ
7N1uxgWx4RvtfJ+kiLb1TURQjPLGMY7DVP0MgkYsKF+HbXVglbTx0dmgHKR71z/zLuaevoLe25Gi
QDrK0Z9QcH7FoaxeY4onKwduoTSbL2iu3f0TD8eABXlMjVqO6oaE60GGUfVu4vGmxmie7vZzVUEI
36WELz/4/LVh7MQjIFwCfmHCou9OMeGSFjJJDmpmGUON7cSRURudb7qLi7KNS2P7W5eB17mEUy5/
70JIxj5UtpZXSxNm08OAdFhtjbQXGkvQYPFAqZo63U9TsYOLeMeDDBwPQ/ATjhkF+JBRfnEb+eQg
ftfQNxUsX++ThiEUTgv2cKBs6d4FZa4pR8FEpBAnXalzVfBbu+uSe0s5dPgDWs2PQi/+BvxA+ibD
USPTshAYSt8yv/udtIJnzW8+Fkx2GZFnI7Ln75TfutG4Dwmn+IgnLRYhOi8SWiLOoIPSdL8A72x9
G8GFHUqVeYxx22ZcsB+POjHz9D0Bjc4AVnr+o0tFfkOLazK5nPlr7uECnZshWrUIq5j+/hhgq+oq
b5nohOUi5Zb5mBYk6qz04DcyFuOp5/CL4hQmyhFB0XivGlQFyXBvamwow1v4dXe76szSIXZp7zcj
w2tIJVMGkGCRxngO6TFe8E+M9dAaz6cA/rAD7Np2gGxylFe5/XF+sKl+Gyt61yi7+3Wz168vnZr8
4lEGfDuV+e2/AMHmmwkOb+ctTNAYfVGuMpDCd4fAhhPNUp9soCId6xoSeYFFFUSC8jV2yEVNGWTB
DRcWsKqkM5ocSLd/momAbGHAaIdd/tWuejqfYmYo0/PimSttf3lUwHQmv+Bf15YYin0dINcwaJ8C
thga+pAdUmp+3Tgfl9Wo7O/H3jrzAaAOtvQwR++AGPhFINX4oTOsn0KLFhg3RluQv6IHz+yF4121
e13C22q0hex8prp0UfdySfhmk6zSrpvwxBIQe1LSAxEUpwVAupIZaF+vsA8hsa/10s3tBq89Zpz4
YJjQ1cmZCWT2PFqA32rss/TUPrLzOVbPiqE9jshgSXaMRM82i2wU8Z4lumAFlmDA63b8JFHPYFmU
ljpa/foePNNIAt7Hup9WHdXJrvCAP0U3uw8T3s7vUTw5Uj2JgGiX1+f5MPTe1Bwh5/mNG19F/+/T
c6pBTks2GIxacC+XtxtkG25tlwRDtYMHpBUo9d+CQ2lTscfBW3W+LpyqIPUOhOI/LLObJkGu+tLu
wbuzg47FCBOdEswkDmMkFHdlU4dP+w1tVcGkKEcGQyHjhXPudnp424Fz3We5xi7665w4zJT1R4xb
kKMWctnNkhl5Dq4sOPy7j778sVHeg/9qFmB+GpXfOYxDfKZan5ejHdLCtAjpKFwlNijxOMJ7vEHH
/Kgqs0ROWey+JFLIj6OZ+6836nwYj4Rkf+8Kx4VDQFM1nG1Ta9iXh+xGYT056SehYN7Ftrms4san
FRR2wJ05n2ZtP4j8Go3yl0M3Ahpd13VgdTsUbdrrEiYX7djJgHuFCgWgzAzoiCGF/ADXVdUv4R/q
e2jmqLqfvfXn4V603YwOzgooBmCx4ECla6tnstxZ2Y2OfhiEO4KNY2fSaRTXfhJ6HrKr/SKNmNbB
qXHNqZhUhW1gwP52KatG3AuFhuDCyvwawV9jAz8bMqhUwC7Nn6tYj1q0qgyhEgyPyJcc3ySOa3gj
dI6PtJ6ubzWWdg3jtClAKYPq2l89/CpRKLBECvrH/fm5wBD/4F/6CQkTW4Z4iiC2fkF5n5+PX/Lj
+MPqzLEO5wjP3f0dlmKmUxRcRtUVpK6dr8iyQxyTt6VMI/CeJOlpWzYu2dzWYsz6wb5oId/kKu2D
j8R1PZXW/ET3NkFtO70LlJdiPkmnr/l2VwpfpVrXhZqWBYL0eUadIebDmGVQ+wtRUH8nLG2eq3cr
SfC83iPD+eM9POat2pe5swY+hTbDyxOylb7KPMi+qlpZLZhOVztYe9LbdUMq7rKhSRE4Wsjo8ykJ
G7nydZUxgZw8QkPneHVCQHMTBwd1azXPEDan3xnlc/clf/EY4GUgLu2fQvHYTo6BAxKuxC8jXU6j
PzpPCgSyYAoolNbg6GQb7W2fqUTBd9XAM7lcz06hoMvdbTCWkDmJijV/7HtYqUywr+s0MPdCi5zY
1howTLF71eOghMTLicU9TZqJgOcKeNl9UWSThvFxGFGDPFxgF7GV7YQctlqLlGizuJnqhFWbKJiR
OOy7IfBw+OWCBL5j6JewnXVZO5qXKSo5zmuW5dB49530ugo0zIkWRJdprkFLPPPjNcSmYOgbVdQ0
6ratZw8VzBRO/+CQhVNGLksC0E547tzX/6bBhbfGNhGcYbLuRlGHLLVpTbJRZrjK+xjlBa7JOwKf
mwTZCBGvwM7QduxMnM+qnNCq9Xz+Jmqhfoqtt1v8eZjNg+PfWaE+MyO/wqz+KaYhbZpLXQy6uKAP
d9p58jpBNUYI4RPV1qQtZAiQlaCkfVRgtsa8fu8sXcFRgR5p085KFyH0aZZF3btvXi1NKRGI0kgw
/+N0yJFjjq0WKsdvw1P0PUxZIRXpq+TcL40huVClwtJlVtuxLgKhdikTNeLIQOpys4A8krQoCVmA
iUwQv4zE34vk82CH71dgJF4qT2wHz+SHPaR5wfwOu00ffOB/uaCgRzAml4PnSp+guGYPiGFaZyim
5chwSVrF6mS1NcAl3lfDwkRIK0k1iAM7vmXsR10LHaNfEjxNbWRc4o3eXvfeb0K3gq38MkTTu3WL
54RRruGolvt5dTRHOGChPr6Veojw6828MmK2/1PApMD8tcJvd8KnfEw6ZhP9XaE1Ua5ZE5/G2gAB
JA/V8wrD6T266dQA6FRs4/xDWIXm7S7+2Y2IZiszGHxalx7k0yioa9DIiKg9+WgkIiMt5cDwpDRO
1arpHCPjLEcRfQqi5aByy5shSa7XM5IE57WR9aLzse4OExCLd0DbGwHRBP4fgJFrHhPWWtW4HV52
OlAG/X/rd4QaSyAnxJj0KBC2Zbs5qXB8JV6R1Xz8Pw0XOnwCArOEJHG1L/vX9f1N6TEyhJgzmJ/o
w7XentZoQjucUwpuv3JsYIwd19wVlT9ECyuHQGomXamWKX1sRZM8Ej5baYRPKdAV/A35FhIYe8yB
c/j1ZhQYJKezSNi/UaNQDU2+9HmoNOzeiYi710dtLF+ERIu9t3iz38yZrkEiKZJmZzPtg3hqmww/
d2NxZFacF33mAeKiPjHoGCHwt7a1ISR5/ieX6wfk3BTTI6tIVHNAqHjw/ew25VohSyUTuxwQG0/n
MewFI5k1wo+mAn79M8fXMW7hfqSIqhIo1GDPwKAYni4eYyRVJr+mY0zpKSHhRWeqwopOyhcdseNp
lIRrBZgfnYrGQ5fvHXhvB5EbBC99GtKPd27OfYdbALxutx/SxDn4anHnnjcCJi6JbEU5UlrQaEFs
51ClAVqMaIuM1loqsDAhz8s3FG0WDkGW/KTpUXK+m2htoO0OpX8Bt/xsoqy4IXNCDCTiAc+NRTH1
dY0436QsYjn7CpaURoMk41sQiFhQLmgmFmLV+KGS4CNY0aDtCZDz1nruKjGYiXTWNOMgGrdiGjRt
j3XroYH8M1lX7pKoJKdaRPGD0pcaWksafBcmBHiqFGBCx4aZezdVf4aScU2ymd+Dm3rwgX2+waB5
/df+e+sMEifIxcxEwCtkLnnNtOdqE8IxKrM+nIRA6CoHKDM9Wt8p/IYLvLqO4pBlwGmmhOW5RByp
VT46tHUel7vl1d5zMy9qMUR7LQAWdynEQO2OFWZPB6IhPKb1ueap+Zvks3L2Ymdtol/9hOKSbCs3
Yu05x28xF+PgGqlrAwrp1QMSN2RAv61zzslTJCRqPfp/Mr52a2J57aw/W+JbDw7qJZdU231AmJxU
qE8B0+z2ZOo6xNwvzEYZlGdpvi8/L6WMAh38QajJgq3AiNPH8Ktzug7FjQAoeAbjHWM/aBFItO5B
1f5W/1fnwdJ8LxNc53afpM3t+RK7GhJ+BP+EdDXJlFnqFmSmAkVFK4Yyt4pT4Zx77UtHkk8rnLcc
r2iN7yJqeSdSn1QnHthvoE2hFM3WG5edDzP3oc2ozAlWGWkBnqAqBd6RDSKdDTY+vGDzSbyRxwOT
RiFFX/XGCO8wpdJPtfigw6CloHBlKvBbTcuwkmOfaXRxpylqgYCyNm+8+E9HlwBS7G5hXiNAQU1y
uupRj7vQhytCiOzpDzDjcROWblp6VvGsYs3a5C8eKKDclr9pxjMbfp2RmCfECwl/JzHNwfHqJzmK
VSOotbO3fxCmxjuWHkIW8lfoks4WatddIkBJlY32Mdr6EuYX0Li70SaboGzbxeeaYsLoUB2HgkO9
e1yr35qPU+wb9VH7Q04E+SpOZmPM/M7ZjEVrti4Cw67UYJZZc5q9AFxJDGzwMeMMaeyk18quf8Ht
jock3VlYtZ6LFiUnWbaU5HsqgluVsVCS/ji22cYoEeAHGBFWjqYqo1T5udpG+IoedLlHnf5scHy1
k6AcBe1EUNpCwwI0nEeIWWdb9OVhc0f7DGvdrW6/SMzzHmS4JbHhAWQurdy+pOrOtiajyZbY+z/s
n5Hx4YKTPHWUvyJa31KkfQDlYnoeWHoNyEkMWIqVHx4k/9YMLosQ9aQNyqInH5hiM0tDubEKEgti
SRBaDUzc49Az40o9wr8c3I/yRgQXmOG6Nmdm4fFMQHnJnXr668wlGH4yBUuCKK61Dy7DU2zGTxst
fiouxwzn9vHsLQydi5s3qDZotFKSJ74DrvQsRlZ/+Mx7oxE/h2JInjWgZv+oitODjPQ/72YBatE8
IXekSKC8c9Nc5I/h9btXlcEEQMrpOEQuTiBe7L3ye5nm+HGadZBJ59UFi8x/R48X0UZ9cs5/Rc2E
qCuwqamk0Y4sH51r47W5E+H7P9jvQaJ4r1Xcu0j6U0wQ2DkxnRDol6OY76wsUfgM/rkScttoo8Du
ih2pLEAf7z5NvOXfIVorSgNKoXsLlXDBNYBPbDYRGZDQMi5LREfA6UH7SYwR4xByfeuzwlmggtDD
8Oy0Cav1ejWwt0lxUiO/1ybLU/p0tKpFR1NG77RqZqSxoVWh29W6ECWvlDXiF+TAmF0+m5DkWIHo
ljNtbzTydHPiXg5a4d5FlIS8R4NH6X34U278JsY9UhpW5biUgE1dKkwM4umOQKSO7l8qTk8ZrvkD
vxqM/AhOkkd3dbyR5auZejTwGuu2inrcKaFDGP5F0Bx0AxVyS6BOptugU+7icYJx3r0An2vQQ4bj
GykqTZSbkG0+o3/gxpKVATSII0GIkaChcf5LfyTf/NshVfGMx5iRukA+LojwhRuKgu57Gq5gEXAd
C3wVh6SZpPTQaV4AdW/ta0KQhy7KAMiU7PnEr2r2S7NHrdjQd3Gl0elG9aLIHreW0DhmS+6WyMmO
uh/fQmkESBqfDX7IvDIylTFDeleRdTR4voiRgA+OFmT+4nuLa4eb2uz/fFm4tbL9OQE31wc52Aky
3Hgpz4YAQ4B3Jc+hsDVyisrlNtGwV173eNC+Gxv4BW3k779PhX90H/sto4xW0m0/MDuQMNhq5cn9
+rUSMJ74FKlhTqNjQpIcntVoMqz7cbD0KtvOhDOFRgBaOLqcovIsM72OP6rVogpoJpdJlZ6GAlYG
Cy2gBe9O9++X2o8e7NgPmmgbTG8umDhau3im/U3pzZVdgsGrN5y2AigVcXXTuibsIBs25ubQ3Eek
O7e5l7B0VDi2TG8HnBKtqJAMAh9JV+taNLVzl2H/R7Q4FCIgVfApDiZcu2HI2ZdB72lclqycSPZL
CW8axfWb/7XWDewA+gOVstzGkOPMiFOXWc2c00BhSYd92YgAUoAoYFwtnTMkZiqWnlVo+GL3IVGL
osTLP1qvt0X/JQe84qo+9ISWiiH45ulO8IcHMbCeMvRYYdmlv2IY48l3vdIPI3QSrH7k9z61wxHI
V0ondLWSZ5nt1cvv+jc/Wwbd5BUsm4Qyl3yOwTDaFYXKnbhLV2YL2vge4Ayua4xYcl9VleEqrhPc
+BA8PNcfDgixZmSBRsvv6xqsz5tlAX3QbV5J0LlUbqMMp5vXSybZWERo2CALAyaX8FjdJHrwS2Yp
RaZW14nf5wZO8jMfLd3mzDI3CXgqnX8UrvEE2xMZYNW1V0DBkB4ZqjeO4E5ZbwXkg0TVSCeLFpB8
uQmXoiypSQFEjOBLz1hBdwE8Z8lRr/ByZKvsvhmSq2LaVjsByN9YqvX578AA0OV/f+2UWOoRX30E
9T84LpQL5ZisMn3syknOOF0eqx75fr04ncQGbU78O9Kf7cQhuv73MELdbJCR6fSV34sAYUblJxLt
IPj2t5zj8gwpsakUVAQa3DNFK5/n3Tgkkk0f6r3OHVpM5E9wdg5PparB/5tG9S7TyaOrGo1Qp8O4
aGfGEiTwl1VuZUw60Xj3TzmfOiodaqD7Qk0q12N+DnGTn4NaNyLG1nHVSYpE8OTCULmbGVCkCAUM
eoxpoTQdczrZutmA6xPTgrqUNSXmmo7cJkWLIEz1T81wbAa1UpbdDkgyo0bmDhxCBEasK9xjTrj6
xOGb4OL4yAcwWNusrCW4JhCWxjXh1VJUBOxRYRBgwLTr/CAPJl7OzFRxKSS0Y4T7UERuckWOYeca
uj9UymbpdjHYcEkq+5sYhjG4ECyGPFKej3Te1TSaR83LMHdLSbL02pA40qgf7ZRVo7BprOmhVag+
aHWhRnNbTplq1SkUwrzWCcit4GimBrRxItfzCeq1Y0hh7sEmOgi8dNBmclpekcw2MSKH5l6rn8Xq
y/wPqO0ganbNSa42fhD8+BttgOXcJ4wHcS1+D+z+4riqyrCtv8fjv/2c2f2ajP+IZ8OKt3UEqAn1
GtpTrzTT9UMNzAboIH9qUPEB9Huf2RQg45vZB5p1ecL84Uq+QasLPx7KTzDSTG3aa5jO3NrPUWGa
+yZp4ZzkAofSuJblnHJejeenMki3BcbiUb3PwefMFg3LUXBqQkL2tN4DCwZiv0ryRJ8pvKIB0C7Z
uyCoKOrrc4P8MtWirJHSwfrXRabGq5Y4Ba979BrPq5OXR33zDA2dtbM1eGsFI07DRnz4t4N5Z5Xx
6bkAO26M5e1ZcYWTWkGEGg9xzY3jSDB4yGwymfutm36P/loyiGdiHsXLqsBJ4E8wiSow/ZYpRKVV
Mu75sz5S8gIhbFQ6Yz2Q+tv8mjyUXa7vhuF1mqCytkYSZT5gaeXAlnJ6TdyOQ3KxwdYHO0TsmfCi
Rg4+iL0PThhtSMA1uOOlQ8ADDRHfsMdj6jIdIeftE+8V8dfkH+pnklTBmXpvw7XIhxYemmdwCfPo
uhH/wjySlawjcj/aAciXQkgAqbcy74HSudqwZgMI7aJ4BRA4SMje+ITE4XFwooiRQ68dpSOZjoqQ
DksAHY6K/+/bdiOj5AbC52aGqQKCCk5TlNlFnrMmB5O4kA9sF9Gl1XKIZP9UrINE6HooLeB2A4EJ
C4Fjm8/9NA8DDoZOrE6kXgMAEdvo4u/611iX8y4DsYlQJ3gR5M31iLJ79h4Xxon+l6cPCJQE4Fy9
APoRrgAzhcDXGbsfAAuQKSXhkh/IhqzAhXI6h0tV/3INNSKtbnRQWusEVdY+Y9eoC5FKp9Ba5AnF
GPRsQ+9CHe6Dme5KKHRZWa9e9VxLsTKTrH4Fhc9luYyO9AinsoDkjKpuhL5RiDEvhS8/+si6S5St
9Kcd+Kdy+QZd1BCl8VZSHlq3Ubm0WWtdMHdAwq2LOcTZVaX6qalbWdqj+z3BQOWkBkjQv4AnJ0A9
xvm1gEnFVJJiBxWTuYd+PRHuBLq5FcAj0zfDNVp2ZV7JbRmIdA3kcmy/oY+KU8fR0bhA2Izr/3HU
PeAwZIYFTyh6gfbZnD+kcz4jlm/9ZORX+JpQjjZbwpkg6EKtiafs21uyLTPept4t3+xnUI2AWFcq
hVFWsCWJBltwxMZVVXnHg//iu3AZo2xLyYifybOE/sWdfgTMeqKmnfhx5feKXUb2J1pfV4bB1Ap0
H1tN9sc9B/7P7TV9WDejzYA6YBLSc/rU2Ag+Cs8DB5lhy5oh26jYzS1Sul1nM/3KkDKPJu1w7dxN
TOrQnwjcplZw8S3hYl6etUHzgT2pPw/nNPLR95mtXlVy9VaSkJ7E6AZe+3plrisYQt0rR6jxgczo
3M2XnB9CTqoG21ND3vYGkcdY70V4/uXtB2ixS1MjxzeP+CI8j7dN9IxrQSSRBYpSjacKG4cQupUb
XeE3E4xT1yJUwQpK78snKEbIZK6jCx1H5gGdA3SwcV3zsw8HoolGKtzCLLuP4iXTq6ti2w3bzmKL
5kxu1vmW9b8ka/oXvqPTep2H0ius6J4/tm+AnyouH4di5TWZGesV+/5bMm2x4NOtK7Fru8VzfXFb
6F3TKSDnhYz5fz2rXxUtV4o98DBTIZH2R77j+vh1bOgg8lttmnb53XkRsufSbJRw9SHw67B2Nit0
nCa7uEvWC6q3OIQuOLCRjhQT/QZa6AYVC6amuwy/NgLER87AoZlIWiKrR+ks5Pnaa3ur6fxcHzzM
L3awC04vW7N7e7dQMOwHXQA30BejG0rJ6oAaztmRY8njgJU2UNeF4SBKlPmPSDtv+ZbgPaHdyvI8
e4s71ypcN+uO+LuXYHEH9HAxJX+/Ag69vsaKJoRG43j6vG2071OWsSXdjQrdjeZFmgtcOZZAUcGe
XRt2jXKBgsf3nXKGFA3rR7AjSHBPrkywsW/RhN1kUoQaXd2igS6vgE0WUZs5KFYQaCDnc7Me6Kzd
joP3iEHV+piAIj+s2cjBznQLCT9ZiW5E3vKMS9PYXyzFplUG048mOMRvICXmMs+cX4XVRHMu3P2f
mwBEIdjF7fyBIxcjl17jMtLJh3cCVwVDNXSZAVpXMXdHOpIpVGmM7O0gIP0Z1yd52PGpS56Iql/L
TGiQ4ESQhb5xTLC4tV2U47dfUwHKzMzGU0hNNDOahCxeziLjtulVPYa3M2vZsnK3P32mqh3tfvMH
hZVNyzNL/o3kRAS40i0pZFdB4KwCABgb+d0zaMHQthJlsuz6KbU2MX/4wUnSPVoFrgGP+YCku3eO
Eq2+tyYV2RXzD4EQc6iuI8o9U6vWtd0rhTbUo6BQHrv+Hn8LpWugENYgx8OFI+lq46q7arycvFvq
h7ff/UqvGIL6Sq48LMXD3DKr7b/Ye2ZMAfSn1aStj7oLKCSrxqI+25BjVLqxiFOaMNO65kBNQ752
+4uFezgivg0jWxvQiCHi1XVeApqvjY4+cxBRg5CgJ1HTsGLQrgT1kf1jrbR5Zlp9pR+7T8TceISx
AcKNsFbI3zuPm1wgT44PF0MNrDlc7ipEEcXT9u89g18CmgEq7uiUd2b8LmAIhR/EyFeRb6OV3hJm
P8Ze7u3W2QXQ0UYxLL1t4uGTZJfconz+snQHizjzriUr7tQj6O47Ng7Y5XN6bN+ZI73TjPLZ04G5
kXBLsxwmqR/Nvegn2NYhjRaGxGXpCpE1ZtvWDgjwgKGpAd2Pt7E3XdXHtKTfPQUgAZZ2nssAAXJW
EGjh/nud7ysOtoD08tgPTiq3K1fLH+qCHjOgekEEqzKRSu70etN5LwCvZrB1KgkkzloMTohQyxj1
8/jdutfa1fbIp8/NJrZIYxorp9++RIbN1e9mDz8bBeTapWCnw8RpGiux26ES4yFK3bmYxtCHP/v+
GgWLoGBzn9dKXoE3NnDeulyU7h/CcbFq2Z3iTlZxd9Ew/xklzSAwa05+dnsXogYSDQbDN4PXm4jr
nw1u82zZQpIwfBqOQ01xwVNO+K2Plx6vw+ubdrCT1Hel9v1TP/bID8z34mhlCHqU52mQNh3+3Zsz
6q9u502UTWLQa+6kchrHK6M972RJ5WgUrYT9Op6+BWq4Fuz85NiRiXGRQR94M5UUyeDyd6ziaNYq
5nwN3ehxd+HgYqe/OcO/4LXqQMG5IUa3RGEWKuE5I++Rwd5fCV3+H3Y8HVWKienfOdRxJ/yAmTeQ
5RFgPr6KFeEyc4w4fEHSIw1/j9r0A0D+3FgiJ4Vfdu36Dao0/FDMQQ3TjQGwlB39je0j2wVJK0e7
bVMt8gMD3prbgpFBANmmhr8t3TTLNWO1j9YAGrNoUlcOFClcb2aarqntuOjZ3RubZCwge615myGn
eQsH3E6+T1gGkcoHVlpyBNA+/VVIl4sJe0pve59MU/Zrw8Erm4j7cblyL2vnM/kU9q3o9XFyUt+V
IpLP5Xp9rvikg+ZLg/4BHAS0lpREUr7mI49WcHMq4Nq1aC0TI3w8cOgrVzUkvbfyTcMnNNIfEA/b
7BN/neRlHLP9vCF0KV7LQHWDZUfZsTDn3TJcTLyHAK0tEML2kHcw/1dO6RHYps4iMJw+TsnWV43u
AtqBSy1GWo9VGQVFdksWbjFtPCM/qylYWHOUoIBjeGHt5GhNUIpw8Mqqb3mAXWaKKD6nZJreDs0E
HxavWfT8tj/3bJo02ADbvfGhrZXxZtduCACpUxb1qbf50J2F6N8zFvyC7DNmRzrAw6DjiEpFrL8y
YqV4cIkbq2a7tdNCp4gkqCZeqVxp89Tof7q0HNu3cAE0/ycclPcscWNNt0J3ZOdpVRRUBgwfmzgZ
q4xZB/KLH23onkqVexyPH+TmAuBNzitwMbwik5/xDv99A/bHEk/EbR9cmDq/O96TjzuiZfLDL7bM
4Nys8xFgTdqR5l8ehZIbO2oPX9HR4IvDYBL9+Bw/gbVAAbqtYBSVfWxHfJ2DVuIcLUHZ6GEbgVbw
DWd0i+/2Y/nGydRnQ872Wel8aDpvj8rO8T0QOXuAy7aIdlYt++53NrYcC3RKM7cODhYS8gEMsPD4
Y8p3E7x3zQ2kkTb2M+PNMILXqiP/dBDmA5q69SVtMCKBMSGzsLNa4FIrvSljjljVMFOz/jyR1fdG
0Ef/8ue6Tg7xM4gasjvE8VE6pHJH1vHkKXwY/N9kQSf2BWGq3J7w1nmxiuLhcHU3URef/1s3bSuA
KoSCw0MNmnGexHIbdxC/3WxPSieCyjjZZ1vz4j9m4BJy2faUZfyL7fkBrFi1ehNXKCDgLlWH6jcA
90ZXOjuTeUPeDHn46fXMMG4cyuEH6O1AJKbP5cGeuvXJ0fU2K372xbVncEyL6xW1qjsZeua5aFj9
W82rSz2ESvfEsDP0lhfILspSpLiALQjqZQnj7vSljMzh63T7TMupvqJMjcEBo3uF5/8dNcNrN4M6
reBw5/VT6cSz82NbMdAX/w1Xi9CoH9cmKY78Km0r6ODY6Qoux3ooZ+PGf62iGOJsGRGid7g4pGvi
FKNW1XwGaIMpnKUNEzZ0MTthxaoQGLCfHzT7Wux7/gHLbxyJc8ts4F2I3UdnXnI+Tq6d8uS0wozY
uZT5zn+Gkyjpl396lVdR+58szpzTKGFmeDsvOEyYuwm1ZUXA9IYWiP/MABRdotfFrtaz3ptpVUJA
XyngyZSCrqT65sqRShP1PSpTX69ZL/WxqLmBVDyg1KxopXDG7dMwKheaeBLukZnd/LM/2EnfpJk6
c0WGAe+EPHiteD4RRs/xG75UlhGeeG2nR2XP233/2Ja3FDpDVLknu0kQZbL51ZPL7hWEaBqqVRSg
MzOKLc3X/r7VyuwIhxXf0VBSLiv9bbpP4xZtMcSbCPsCXOR+vrqJTG/iHdaklUA0UXc0JST4iJdd
Lb8JpjIAVIOtEXdNtEkI9uM7nnKBGVXqyPDmo64si7gkbJXUcjtQv6+tazz0EA7WENi9vyvxjlzt
+yMvojHAeygvIYcRxsxBUq8nnjwudrghfyF4S+P7H26S18BNBAIrDFaN0Yy4Q0kicL+aF3sZM3RH
x79OOt9v3TAuOluWVY/v10baw2QGX+DdLm0J0tARnGAlEmF6rPg/7EEaV4M7IyHqGwdO6dE/rOz2
+qBSwFxNysLqU5elgBIYzua2jQZeJ7dgy0b4HE3UP5aPkiteueuj/hJ/aIpHH13SmOHUrqb7a0mF
JWiIm94bqpLUJXlEqysXvKKogHHXL/jWhvi/QkeJorje7CXhCcgXYasyNsM2vUfTezMFknIGcdCv
zwVrW+Zx2hr+PLMGVUJYjOs1is9AC2pmyJmbykL+NxM8iiH+13EdA0EPw0EMNOzhxOXm1O06z0Y8
R8QtLxZS5OuLlEB6w9dMEKsjaqlpflZ0vmMx0NfK0q+Ic1p30ROHtlv2fuuT6+xetWOQqfG7fQek
69RGPqNb5kG1KfdX0/LfiSJr/ZOOh9s+1f2NxR6JTZPxvicdTUWkSkgikktqdDOtb53poTBd3NvF
+JneiAzBSddhwKRsOopYyjrmfObIyp2ognDhc+NDVUL87sDFcqeSxe0CAQqiArhFbj81g88lZX4y
znZ3II6vGapXZQqk2c6Si7SzpWPye9IQM7aI9OmMg+sfu9um5ysPtZyMxdkptefJDbCSIWwAJtlt
S6KeygF9LwDbtb6QZTfWLevMtSLYzUk7GhXI+NMSKW9vQVVhfeAC9rVIAPotpbTnKBk9GY+okQqe
+Vm+hsTgNgNBPA/9qGMFzgADlgF19ajN44NiM1OZIdsvPjZ9CrHBXw9bdv8JsKazpcUn7QfMTAdZ
ZMhC1jwDVPTkA9eipqlWp6OAhv55Qe4jRTpcHJVwKBunBnYbpG706sYjmiGeqztWszS0qRsiRAGK
lFgnldmRXzyceXLZJhaEE69E0ets16lidHf251rjTYRrzOr5mSVOx3wy3vwUlrF51LUWriKXX4A8
/hbyODT9rRl8+QbKVJzpOTYfFZoKxcctZU+nP0Nif1q7mOENAJKS25ySscDDPvzS3VqYwrgUZaT8
X2ki7HO5JCm5FmgW/wjQlsJg1bMLsOXDnlvrDSRezknaM3akRNpEiqhxaUGHIBEVI1Yzoe6gchJB
7kgKT4kCG5AhLqpQkL0jefus84vPm6TEERXahvHVKWNQHjUnJxzwbtxYsYztrBN6jOLUTE++FSow
9vwi/+3NKrj5y1IY8ZfBb4974hlOqF2SN+UNJROTuQ6YpcLbLRBFYyrQrFbMcSAEZ5C78Z+xvICl
K0aZT3oUkFqpCJ3Np4zY2AR17yYXJtyTV+2ZGQfsp23YO/pfKK1Qei7+IjFKc7LESlKCdk5FUggL
KppNeOegwtE6pxndqYtpZZgf0gKVfHV6h0VOgRwdLo1FKPZrZVXRoS0kWf6SJP+2uMZvHSBQVd/N
I/aUVU23Hy1x6SD6aEGjRgJ5eGNipXdRi8YykLFlS/ytIIdJyneZqLOnd/mpEW6ohWuati/ZrRdi
hvZA35NUYDo3c7dLTBekRYelNnx+AMmLVF3qNApboKjlslgz0lIMaZ00aN2MnboTriC4HRVj8cCV
nVa/sjBZG9FgQnk7hw+CZc8EEoZus3O1QckdA5sWKujiFF9SIQWTio3NwEHzvIlnfz44KbnAHDFR
VfJGJMTmDBhxnrRYRzkdBfQmCbkN4I7ixW2zXRG3lSh2QXFWFLiw361CADm0w/cxtTD+nXjIgfJ5
wPuzUAfn5vooZO+iGhbqZuEj2Tef1rPrbHYBKT65hWJDZxR4c6yV5QOd/cnYlhwUbYAl3CoAMtRy
KBLbILF/Zq7rHo0asD+dkHO/aW7yTNPjpeiIJ/+pJWMIIRcXh+9axOX1gtUSyzZAYiR6kJvFWadZ
C//XglgzL7Ug18wau+59xJxQYujbhhqTj3QNB4k7drEHqGT4NoxBEGNVM8j8LZlaV2mg24JYBFMj
/Ju4Ke3dpDEFerVf67eJSaatqniHyJTZwBB5UDDsRb3NBWqGpeQZVjy7wDLWnnMF5p5BTiR77PsD
28F/CwsaNUcY9IdddOGATQGfGjEv0N4RK8svjnYO/dpUIGB+NRxvmXStsejuCVhULIwfT0XSVxFL
2A9EnFfhhp4EvEi0Z5XjYDyZgriuF8poelOaQMCaYKm4wn8/KwdnHTYDfBMneVeobiVIdCpJ91qT
MpzNkcxZ2oOV7/5Th8f1cUYHi4GYSnukwpN/dbkZua+0+0j/GNwQGIslBCcJFya8rPgAeFrXixqM
1bS7y0yFQsIx+IeSzpdTJomhvheSmsQEzLcs8ET2cSawmdUE6LBMC2lgb6J2bghfepElWlD6M3pr
SHlCO4bWewzZotWIHtoWr2nlhJpbHUcriOlBAZFXNTcVa3jnu3DqYTfxMfQhNgEE6CSJrvGNV7iL
jJ+6ORJOXPpW/es0l/snOnpecGNCBxYFWHQ57Pq46mSTWpxdFGu3mjk2ipCGHXWDJ0Z9yZTrnh65
PTlhIBCE4YX6IQhCu+I979OBnHbcF85N+nzYUPTnegFKzOB/wXC13Bi91UnKOWiUO0Vv+sQ6OiKn
wHpxJTEgy3Mvft9cpiOefQYJkZeeE0OwYgKWlDU1qhg5AKkzEuc5X7+Ktj4N7K5S7JRzoKFU0NVS
rJyFlttDiO/S3UBdF2LVb1vplcQKupigPSbEggVdUrb7c0KFRePxJ7OqRc2Tz50R4Ng133q/alFb
U1ci+82C4jWmyR8acIzgksAwIWDlyMt5RtYNOsTaiwOV26cIuiSAjFKb9HVuorvvVKdVL4r+KJuj
qOEIucOPBIi64MpD178qzUZTEOHpg0tdWSANu70L8hl9iP1fkPcM824M+xfZ8jZHpHqal1fV2mhG
Lnspzyeo8eNCVkQXufmkv9B3I84O/SHJyj3B1XvwzLSbDugS+QTEy/nlhuZk0+kz8OyKZIMW0M7N
4FybxQG6Fis244FQi9IJcVVzGb0uly6HFdhUDYtb00L9agTvXNMwofFX2PpT7/0mpSzWwXHyJlUI
FBb6fPNTp/n1Lf6j7RF5CeV+SbugYIE1GqFNQjpq6a2BgYqc0QgSYIc/a9qYVs2gCwdRcsl0XDxf
TkTxjp++uHOaZdY39fFuX+UZw+JwlqiKYlM10GvuFdOu+EKjFuNwdN9EmMM5Pv54H3/hxEhkqkpM
5u1siZeSxjyeo+Qv3d2hoDjMI5Bvhv9o8p1jEsrn/20B/8ERdyMwvxerZuXbe9mmSCzRtPjlVn86
+PdumAdNUhvw0nSd2IUvqboYiIBOXjqe4XGl5eZGma5612Q46hvmy23GIN4nEs3pgzCcHA0DPeyz
8p+S1EGWuyghhmg/ipDUhGolQaMa5Pl4zCOZzK4RO/Ma+K/Gesd4uqCNbJHO5cs9FInZF675GGo8
xzpgzz5wbceQgAcUM8Egvf2eRTtn7TNgjkXmAnlx+FBXqwnPC4EzxV4HgApZrO2UQyx3c6jYA3Sf
GEUTWb0LeIxvEkoWC1V2ikC57uVjA1awPv7SF/5ERsDj5J7BPjy+6qiw1516yvUB0rULuE6Typp+
4eyMqsdV3O/XMn63ZEt8BRfgKUSEjkW2YXrMBkLcDv/RMC8Evrq0ExGpLp/lvMC/IH6IQJMfwYUE
jbxznZqFuyn0SiNkEkZC+xXGLp9NBvXbwmtT3s0bcOxZo57c3hHtBeWzWgfGDV+nIT06pEt4hWrR
XkDPbt3ghLPq6YNhLVrc6eUgoVToSdQP8flsfiZv49XH2r8PysVH/YsrDUpFFPr44mgXm3hH7nu6
mjmg4yeR8D8mB5pvRZvIXsA0rl6gMEw3ZYnNn9DLOZ5D8/OJ0mwjN8OGSJC0Dcq3EjtNAHEtsskM
ObA+v1if/wqgbfygBJfTcybKHXYCYotn4myzOuvWpSxpRFPmpx5KafSo63OkdbTrKehOgfJkhd+J
QYtZ/Ud2phWJEiOEIihS8Gjz6xX2mTtihPVdI/GzAcuS68CTxhCu1KRTO7Dmo/u1P3P6g3dWfZWm
EK2yhNpe6rPfSIwLFjg+4GdQ9a4djkvEF3x8x2KcL8x1fW2d6NkWBzT6ApeWCNWrLmkBpmw1B/Qn
F3anKi4MW1lgq29548ykIl8M6gO0fqScl/tlxJVOE148S0zx8p8b6p2aWbwjd5km4XQaIfuMVvAx
/nHQpO+tARsCaGCSpMlk4UJjZWcS+4LzIayS6FlewUkLOSODL4sD0Kf43+1eXf7katZaAeLEwIcC
0bqKl7MyECbImU58mQPc0uAo+2iod5TBikfw7L1qwxsdEgomrpwSCDGa2o0UGhziOKoihEFwjFuP
KB0u9HAmagxz5M5GkJnFXkwqr2HfQ5O3ldBl+yQ9d5bDzd+KzDgKf4RzGVdT9dBjkNWC7FdGuLjE
YXzEujOnvMNh6QY3aLf5eiKprJ421/WhM4NHnSe/Ar3bQTMWGfl8bSmnjUT4i0TqxHElVBCWKSG8
R1MLObsGpq9kq8lrhVj2GUD50TzyUm6Uu2jNjBSPBwsySAyAPNMy1lEcz8SLEY5V2Vpx4Sii1PHJ
ePRIxVdJx/tTqKmvFaU5MB0Dma+5xgL1CGEq4WtI/Jx7pe5uPJYgUNg4NbIjWXrD8y/X1qRSiQG/
7T23mDzNCOUS0hZCpIts9DyB/8wxDBCuZb9ndojwL7Ar6aNL9BcXlItBbvjFAR0z62AalcfDX+kk
xFmPdHFJI1jWnnraMQtr2Wcdg3KgyDOri8m4UrnF5Iq1onfvzeQuUdeAfDy7AdqjhdxKdkCxJTGD
qe5lhe2BvCC0DWKjjSd8rmDzlE7qwHYIkgJOa6h2HDVnsED3Ur/04fy5pyS8v7oPQZzNlEduY1kc
U7j4ilsOhI3bFFBMHvjhsPFuuPFD/aiNbDkiGbiCm552CYQXoiEfw1GzT37OGlPwdE8atCHB3lut
xx7DA3Z8QucnfT83vIuG9B512gWMq20N7/oB34AfkGRw165/z4P4F4nmwapK9eqQzIRPHwpxI/rw
jbzfLYeeWCPdsP75J5MQXK6AB/gslMobHTCm+95b6ZrHdQOgYo8wBsAfEunQEVviyVtbqcrEh98m
9H5DlU7cc8/MrvH9YnokxQLUfLtWM9Kr2U7m2Q8pvs/sBiavLiTfcqaAVLJM9Wcqhflwqi+xZ59f
W6Nu7ntdXva6j2xfBC9zfGOiwpNR3SXl7QPZpdWB9S9kxv9gkMRIGELG/Q3Qo+JgcsQdOTL2z/mw
XxMqP1OuFWqtY48XiWzqUORTz1r6+UZmDsiH9Nhy++DVbpL6WDQLfA9zxyhFkqEYAsDP25f9WFQB
C+5Zbl+kzOGIcELkyyvbkCnjKt5OCNhaO8RUbyn1sSF+mCenZO+43eZRkEbNmsuZKae5sfoyI5Pv
7y9IZfLLRVMPj4y4G+cIrEs1yDTgg43poVFtVcNfGpIqYTSjvlHRDh846mSlmTG5noSWWq+D0z4c
daeaw0QieVaX1r2sFqgv1LXM5BGt3KYhkaKIdMpJ+271GklgF8To/SY0Km0SYU2Kl5usmiohuroY
SBEn/4TsbhnX/v6su85+sc1M6i4gptc6GygXW+81Fg0DXMcyUgoUxiStaXSNqhFOeiechuDq+O2m
vLnmlEdPhdJuqrepBOv4P1qbKhFsD/5+PZng+g5ERp1SXA4ayFlMVq7yaPliSZrhthOu4mewkmif
g/hWqT8ueBPxWu+OB1sqoIt4XQNBVXtM592+XPsxXDUB2QcGgpw34y/+KXvpbi7Y+/8LosQNs8Kh
i/R+xLYk9ZFjE6nFOhlbIJlU9FxnOL12Snqz/PE+mdTnHSuW+Uo9wP4slMcb5zQIA9o3ZcJHUO+M
dhPF1MS8HIxV8bGZYS1HGum5Pa4x2E8/8/Q13M6lGrMO6OJ+ejlILYyjtaBAkmGsMpC+UOhPuW0z
HOCngWELmDH3v3CT6mSvIYOFL2YQP7vU8xFfIjYIiJJhyKgqZApAsX9j37uMh4+7i9efmJiz03LC
RVzIk1tUh+t3YzGoM396wCAAMQzqvSpF+7FaZ/rSdGSOm8NgrO+Zpk2X4mq7BlVaWqPONh9DNGxU
aF/8UpzqRuieFMEjHS5Gbk30QAeMyB5L8W8HnDqynqnU6JNPSDuBaTFZwjvYiQSXtREEx525fHmh
AS8/giMqk0uYUc4Jz/Tn4oEEKgfattHHj3OsBjUAZJb8bDg21CoD1dbqSgEcri5t0RSOmMN9lmwe
suj4uSQhWMIW/82zQe9pwmOxPOsyjSG4J5aNuQ0MrZAoqIib/nMSrhhVbjTHuJQh4Wpeu/qnI0NW
xFJl3iEKrUL1UYczFHe6Jrz95u42EI6fYhjiJVt+MBXY5aarxEos1bCBA+GN6VsIS8Hd1Lhnkcmj
aY6oF/5cCB7CTvSwWTN6yq9dpfo2OFUBcT3dzs7IJr/DCrypxmdOetslq3PXyBAGaoQO4lHcgjCV
KJe4A4wlDpHuHvCCf5mTKxE5xaWYbZIVAvmt8Z6hQHqhOk8OzaMw6vDUFLLunRNlsp/xp2OiabSd
OXqNX1kMrG9j//8yUqMzMv1+4iHzx5/1LNdT7MYmkT/rNlrxfgBejZgUSoXKDdHUUsObYuSVP/NY
IK3lMJRxMfaQ7iz2eJlXRUldlm1X0brMvsnMija3hXt3jZkRtuJ9HLR7kuyj8veOSldZKSqSU/au
JmdHxiWzuPWLt0fLXLgB1000HVRRbvX/hK8rYvgK+oGvN0hps/YplMxs3H+C6pxMpxzR9E3TjhzQ
4kB/pe4tGbT7SHFw+BN3t25XJVVMzQH8xR4fdz01hsWyKbe8ZfJBki/zk2aIB3A7KykycDCDkoFX
UwRh2W0xssqG/gzu9vvTSH8utY272UVK82qPEdZN6ZGt7d8tWwY39bH5805qjDS/eUE7Ch2DbrJQ
61U9aiuEAB8G4A4JXQFpiF3BQF9VMiY0P8qkj3xllioZkG2hortuQEzD5vx5uJ29otz9nVDnp326
jEDfPy4SlmsCtNIEdmzW6PVuhM9hsw+xroJ03ApdtUayMt4Ykz+Nz8k2PA3H93yE6vJ3qD4Lhrk7
rxMB/csVzwdao5JgvKD4HVclyY5EcWx1jfdNhhvykJgpSMBXPqkAs5j3Hm6ia29T8ib9fgnTvdqX
bllWXKK/bmWFAeaz9EF0Nwqx5p8xVoMFwuKzMVLpbYFRof6lAgORFG56DzO3Uv18ECFLRodt2fS6
AKyQQFm+CYTC4pVs9fNDxp+A1kYwKa/Tl7HOlLun8hyo3OSMOvrLLvB+9xnve1Xm+JE3O13qViTm
K4Rqni+hF3Bn0QK+LSAMkL8IrJej7y8sh9c4EWrJ8NZCcTYItyjmCRWjej4uO6o3f8F1MvzIcthl
vq1T3QwCXyeiaDc3cKN7qpQkBrM1QWYuCvIxPYU6amx2HqGzrPhb4AefzuxrlXNmB9c2flvSXSa+
s5vw8caqHYRu7xPmQmdu1AUKd0E7VG7Vcliobv1QK7uNnq9oGyJ/EdCu/I33xtl1SSAMb3Hajc5+
HgnLYXUlBjIMRvJG467qvKH6yR2lRmof/iZuoDWUnu88gTnmJys1k3UR3Pke8lWkEt9YOiFGpg5F
xMGbJd/5Ms9fCSTsKFoaZNXPbCTrE4R2FXZkiziH+o4nPa36hHW5X6TZpHL3oS6Hr3gNuQ4UQrnT
DHBj71AhuEsUWGYtmiUHpFXJ4ruw+DDYgZI9yKvY7JC2C2frcJba8kaeMK+KU7MsDC4NOd8mVhBh
2oMIzO1mcxc+GR89saCSU+PqYWKFLOxiCvcWafACCngJR/Y9XI/PzK6PH2mhUzAGOSVvzKGiDR4G
bLkE+aQ+k44UwqQ9QREkeCS+onpZnZr0FpfIWXXkdTLwBkZect7u1kGoTxXaahZaMDcXUD/FLZRA
o2TxFJ8Z0DA4yFOPFl1KQrcfRrSRZhQ4AChiguHmslbnxkzD95XaBDPjHb9qofyKThp5DbMg+Hi5
Otxf4WUYIlfCri36VIjwFlLI77tGlk5tRIE2ux21scHW1ZhDKEY2z052a5Lm/DsjOgzoI4YOgni1
/wt1aVYZY/8XU9lxpyA2t7kouPGGTEXJXyv1/7X4tvIgf84m0ZIvAJFNNV9XnZKlpAkrWyKTts4Q
/IqirJsiu489Qzb4RxbIuGnMk9PjR7UPpHXtk/gUqCzOLdNlCYJR4IMz9jvcPUySoGvovPpLumNN
2MSqJYtQEY1pVq/ZR81x4uMTV24RYXAP27oBC2gEuwRwVRIjDmC1ocUzfy+4e1izmrIBbMBryMDF
hyS3HaR3bsTvb/k2j6GYnYARhIm7YRgqHBb/lE/SyK2d5qqtVLpDtZHh2umlN27jKEvgmMGL4p9l
JNVDbvL5ywCbwmOzke+WSukDGQK6SEA1AaDqA7tt2dglhjGDMmsEoj+OXqqEChTOzSZq9nJ7hWq/
usmYJLLizTqP5vHJqVz1GdUZ1rJc/k374lAXjiVhe8YQhJP1s3kz1ReCDGbPVhgBDJoN0r2xlV2m
5oCi6xIcvu5YrFgdAmi8CQ+pz/v6yF8XRSUF5YB4cJaI3zb6MrKX7POjSpO4T1IlvGZjg5vMCRiv
253veBK7HbJWWMK2TQjYSRvugz70ZuPb59XMGqtct/ntZV2N9+NrDtpptAp1ow0+N6opLumSAh3g
45xyf0pyipISDGwLf1Faef0TQjuhU4bz0OeH0Tt3s4HkxF51glh/eMnRDBIkm6XLySDqHxpYHYoG
cGxS+VPZsXDfT3S5d1j+kpxJGISsInmAUYulxAtcw+RNnlySZd4jkn55f0Sk37p0YGI33Ol7xUbw
d6W6Ilea4HGXwhwlA/FqC7aq9UYsLzDnZPOTSgJ5/NnVtigG8JsPLd+V4CvoatpM+21+QtaeugAy
EFN5DDuCSeKWjrIfoOK5u1nGjRrCSVgzbQpTs6opE2THqTIR26pGqxjK19qSm4SzFUSEnAOMclul
eTwX7EJ2j5iCqBCE7EJupkVrW/3pULeXD0RFqis4eBYlmsKvBj6hsphoaquFJVZmqnxO7nZQp/Ez
y2eThE46uvQHHn76ugmndr5NonwcUP9oPGqiKTagFdHsIVG3FTqMawEjzu3GT+O2bOwIRQLSO1/I
aWsT98BSg9SNpsG9U2IAqTdtEOTuBpO6fawhUfzoBnZLRwdXByX7I64yMIZsxu/fbCuZpttA3s5v
R8IA0nUnBGmXkHik0dDDpp3AdSO67rvG/e+iJvxQObQJKoOg0hFtyOBPp4GXuo9wOEvzjc6P29X3
8hK+ennyA5pJql1SITVS81i+GYqFPQWws4jI0TYBt+KmYdxyH1phDZu+aVbG275cEgLellBSK0eE
S0WJpoquNvENvfZltl6d3grk5zWE5boU7C7waa03DjNSyGt7TeWxEDNHFGzoogEykkCk6V0WDcIU
iYOQTnivD7qMQ5qVHKN2kLoTJHUFbwib78BqyZiJZDkTv5LyfUlRA3Adr+mSQz3p543SjWYJmr34
dyjKhZSyxB1o/bkjC/Yu129RU5daiprTN6JYIyvzDXZFjl6X7iFzoLVdkpCWoxLpgrx+StFfUQAi
w9HLV+fR1i0VHPUUUzdnT4JP40ZvSgPQplq3WrWzxKQ7a3wTwgoMf+ENKV6u5D2qsb9W0Eto1OXY
E31pOpOoGxp5c5+D0woK7LN5mbUd0URWWrpI91OLiCsceECIw9k8BP9XxyYgnoxmsSaZRANqmhwz
X5HQRGDSrcq3k3vsExGbzS/VPGO+oGx9lH3uulAVu0dOQXXgIwj50a3RuQVozSMs0RSvVHL9A/7n
TQMSQepUglLwMgnfB8LJYvu089ovnKQD2JZHDqy0HsBGmqrgtTQZ1sFZJsVkLE9d047WLf4zv/3/
5PJju70c+bMKdkx5U1vELTXmNlNbYHxj5llTzRc9S2FbNeKYKuhhEV6K1M+Yhk8kafO/2kI4daDc
rn9yLF90OD2lJIXdrQyyhfQ27iYti7oD0BkKJjLOLGDZeTrXEvQpAzSq3URsFiVU6qayU0qric2n
NxM4YNAaHaHczDiIWhdatM8F+JcSv47Tcb9iRzWoJ/bX5KxiCBDg6nL2EnSAr7vUsr+fNdCZw62D
RRkglulxcjEOMeHloeMEpeUZcyjUj6xkI/l5XIMXf+9tKLM9vlWUPOazT8Y74LjNvkyt9DwYbPZq
QCqy3EC0kRTgexxQSD9LHdGdLupa1HV+pfZdwUSVgDMPZscIeLreZFRm6+uvvVZPwags8NLL9xdG
xkPjiWPX6GdpQTwfoPgnlwI4tZDQz1kmItLFsf/ASgeimxRzV9EQhA8HhIGyozkxIy7rWmhTOPaj
tCdDxqJvC3wWoRM1kyl0MdNCnv8lrC2t4mBe/UEkiBVve9TdEnOdZ9uNSgCEUM1WyL2YyKZQt6of
4n764OZgqlm0kAdPjpFyz56kUBCaIg32b539Cokj3kEi03/7TJSINB25AJrvS4D8nD25la6eXs+t
nKTc4APEdqYL/Uj7YtqAuaVH2IqauQ394mhgljM9jgS+MCCXjXWHniUmDwwepbFFl8gmV+NuFzWv
xIjqxtCQhOoPgpEu9vIbp1LSqSqybV/jhDd43G0Razne02Ql5s73zgt0AbUAHqO9a6Tn3589sf3g
fclxMoIAHHF/SVu+HaWC2eTJUbU8Ycf7E2ZnhtFBz7OKitC/vauOiO05/dFZr7gg/Fuw28Y888JM
QYJVIRgA9q9ls+fowozYWOl3Sslghz/JdbvryyfKNHS14HmG1PGxq2awbv7SKNKBY4ZfqlYBTHnO
fcVFsnw1RKVOfQLZ1rd41zA8wxbPpYXu7RrP5Bna/oKEDBVU7miZusl6gGCJ+oeqFya+JPcO5j78
YsznFYH53uyfvlIX2hj4J3hhm7uZCSwMEXzY1gAHXKmLOuV9a79ZM6CbnhVCaikRKTgs36eXqR0Z
aqB1JCbL92hyTw8Slk+7VraZ/p1sMYGIs9UrsB/YRr0QS3aCnNj6NgnW+z/jGekjiNO5Ofve1V7X
N5soemoI46/0o+0/L3YDq5nKzbkvNsDaNFjv2lWvpYKin48vofaeXVzSWccxoiZirrF+dh1DFIyo
Vbf09RGlANtpxkUYdnDVx8JfuMOh/Yx0kMGA22Qs1WNgOumnfsSgIQmm7Z3WMUGE+ShmWt0XOV/B
gXuQLTccgYzLoN50cp7HAYnYD1bAsBoUfootCmTwVjzhIMn0BbxBT5VX5s9v1C4YzEsJX46HCZ4P
RjW9GO9it9k9MqOuIUfu6ySyTYWnIRJNNXJcMyFE0atEMvmWgLHOuckAyQhw6Eh37zUhjCiQAzaj
40SEvkz+6iwzxVTRzuZrLfwo08EXHafP5PWtDeAlvlHpijg0OTfXkUFNcFbrQgcWfKtZShkXbu1d
Fdrm6UJkoN/PrcPyziYe6qH5n40JQkr2QiPmu4IMdnJjbF+wHXdQWDy8z3Lr1rl/jYRQkwGM31c5
wvzS2a5DVue3tRP3Pcof4uHkVabnHgssc3A/oCwCHVcTGiVDui3sV8gBiNBayTDaGSib6BVdmEEc
XIeriOkpxofUfqq8QDRJigxupq8HcQKtxJuBXzU5+ntbJjr6PXgh5NqAQLGZRQvz6xlSKvMCF6GA
ihw4qKItIgyzZhRO1j7bClwIl+ZCAUzFIIoa6+TmROnMiJKLBtgXjWl50KZuUB4QqH1+tyMqBQ0q
AW16SpZeVMaQhXo6wuPrbDpJTTdYIcMxn3ASnXJZoa/DWJlNQnhtLtwTljvH0FXf6p0Rgk2VeH/q
nQL3c4Z2GtEQZHUw922jQPui0XkM9PUjwTOggGrA919WeKBujKRG6fUjv0RGMnl2IIgXdIf96JQ8
5Vbr83XBkNTd6LV45JlITiO4vkLs91B6Jyt19x2hJSHmkR6XH7hxcFHFqIBZBjAu8PX/nyJW6Yyk
U8VD0JTMBENgq0OVhfphL7olSLB5qFsETrpqWfPjoHRP0yFkRUr+9FgMhCHLCzDxU00auB/7UFPX
5zGsny8elCaMS8E/aelUfnrXmvicEyEr3tH+omeaItKHKsEX5qZeeWP+clESkJHDoc9O+ZDnzEmL
0qt3vt1W+lODPLGb8PXleZm6msSC33GWqYSvn8QjZu7wFJFIHNEmiO+TRpDDzEmpV+eGAF0Bd/Wi
LitFWyzcFuiz/FOBbCrri32mCTtCcjk5IJMMHQP+W3lH3Vr6mXpprGwL6vVT7UvetUj4Ny/7Uyns
Ljgu+22d4L18M/fAoJp4jOuXY5K3FLR4776YNQZOn7U5N+a/+bFLwzU5mq/STTTscf9XVFG05CKi
eU0bI4vWqp+cdis2EPNGhv37HOSpXyVIVtlWpt8hcAq/qQMMS5kG0sRZfRUpa9gwbjPZGdsmQMj6
OvwN8DD3JV8BU3ucmzMJ07UqNtJ4Ov4nt8TLfQjKk3GtGubPmkMbps7+Oa0b2op2jeztAgTSyuvz
sDQVkHY/LBKL8i8s1CFcVYT9CojCrxus8wiX/RgyNjhEgBNjeYdwt5TYqiWdLLCEWro0pfBR8KOw
V2zyd/GLH2UQ/xEwKk1i63xexjCvqOluChn0hRPXoRmgdUILFp4uibPbLqvfd9a0+Si64ZzjJ4F1
nF6dr2MSFK3jx+ZT7os7ccoPSid6AGXur/4dRor9N3GsCq3mht4WnGd4909XUHym4g6ZV+FnwtYg
yKVoHe9ZnOyXnUA8quvquIQeflsv+7egtWxWnLwqSgcw1xaO6+ID8kmx8Nm1Z+SaTV5aAhP/xSoP
hLDO22ez6QdgNlQrLE/Sh5R7P/yPiVlN+TxT5rNDqR6gQ+H9XxRkuExk0LvOGs4mAsli28LD8h6J
pRYXd2s1PeLXZDV1CXfBqXkMNbG5YQIuVORRW1gvmxOTsz35kL/d2VhDj2v7zJnOnw9jF6hVn7KZ
4YcLEjPFPddQHJOU8pyb0ljA7pgbeJV6zAEAPAogWTDDzFHreJWBmDKv3rlxsZAPiDLWjJw2cvwr
PpUH452KYw8Q+0QgLqV5XPprX7yWk0O4jdxb/OrjlsJPGPiX31R7m0fMGALS36YFWih32xmDsnDE
UlMmb4b3fovGTgbbX8tkPFg5BbAywBvTtaxQQ2sakyoYzasUC94qjQg84oKeoO6mrhqSYURXfyi3
GRtYEUIL2xwFHXIVp4dYbrUrgmAbXQzIZSnttdhGwXTGLEZ6oyyb8ouL1DkHHp3dJ4VljPSLmQPG
UbjFISZwF13C9DJkz5H/wDbe0YDNCFA16CkFIffm9/vdMgWApOB40kLQFivkyXPUct/nDET1iicH
2eYZprpHsSabBqHO9RZQ6IxebvTJV7w1g0vDlQNRT+4Xidw5qb9FWZ3e3mcRm0SB+RzIhUiwd7YI
HwxRazKOVu8uYwXIVnfk/65UlqlPAYPRcXlYP7ZOJ54cYsofUyGG2gmV+k6Kksp7gcbgUYAxCTyr
iVqTI/kO3ixIbLV15G6rSALeU+xIFze6EHnvqlWiSSJWFkJba+gXjjq9wrV9xlRe7DIu8pTGEWwP
0pBkBJpdWcTwS3SxgDDln45pi1PL3d8WFRwylXcrMqy1HnVLOJFWdn0NV+Yt80bN5shKNcK+/F08
1jRn4XtBrJE52pDI50y/D6pv6KhyR4D8OuCizA/M6+isL6/J6wstdaQ7ylXgc1Qasfduh7EPAFxA
6afvUxR9yS5lOAXml4+93x2CQyzUHpOFsnY5zbup8b5ROKTvSdy2tPanPivgjtu9f3oxlVsu74rH
aSuskuXkXycVEfXdoZ3TRWy+9ez3vYLo7YjzhXiDwU96d57IsvFADLYfVzoECp0Z8taUIFNCWzhG
vIvCmDMfZt2evk20AHKGRsOEH/8tbeesdUcOU3Y1UFiUEDMv0I6HA6Ub6AwtdqYxQ0mHwE8qr/NA
4H+4ufr7XGgFwQ2wR5sKXGcROPYQI4h+rzs0L9FBWGlnlE402MNzqnYpp5T3E7vAbfHX47mpkOXk
uxYDh9owfAqs2kGE3/2Usa2Gsxz3rJm+fB2CovJf4HY7BbX4LYV7aUyOb/0YKYYgwWedw/vBdqP/
dzbfCkVA7CrImbosA921jOy2dcdzbzx4Q0PoVy2ol9J2oc3GZaXlABk9GocAYrGlKArh2zgj1Cfp
/3OQaM7YnsnTJCGZQQBTgfV1irzhg6soQ6UsJTS1+96Cjd5T68NFzHEBr3Wew3MEUX4011I+LCHs
VUTFqQjRxp4DC9bBX7Cm+xXJSlDrYOlnBMTI83aBtGkAo+ZuipkTG6Ikr6fD3jpasGcHmsE6KnHi
oSQ09O/QyhKRZs64q702XaZOoe5Cq1ddOZU0G6pQvCjsfIktLveHZ0Tnb6TRRB+rWYL4raxgA+el
zIY0ipXTFRHbZEH8tVyX8YA7cZwnS8QPAUfaSPWawmt8IFNz63HPCQyNO5D4cK+WbjhqBcOx1NCP
J02sttQxxpPEvjgZLXBrCAIftRTT8ieMa10lGHFBQfVTQHvh2h4J/cXotVxwOFozJe1lSX09wih4
kv+QOjzjURCqEsEs4cZcKFqooiertXOI4S0Gbh7R5sfX9Eu8tWsp9wZYx+F1pRiTBw7bPhHGpLNt
FEfqpEgrBd44dV39Urag0LqYTmf0Q/nX0wzyifxED9FTv2zd1VTUHLK61Me2UMAy9KyxsVUM5uP3
2NRkaiX18Ra7I4vn6nnr2KC3JzyNDRMtnpPAfPcvTpEjXdkDoud0bc9jsV3yECajQfjT+pJvO9s+
B9/kurRCVmSNHmXNmNSOG3riUxpNPkGpmt695irOVkJXjWyTdgMQtoxmt6GCJOOVibTcenGwL4T4
XLqi8/fbjRt2uvMgyidKXjf9ZO6NpE4i2t4vKEpZUMKgV/F/OVjvsVG+dmBefIvUpYZzuUGvh5im
eer/r3RarfxXoa1YvRLdSGldEVld+LVp1/3iC145zK0KKxWahpQhAR50vvqeCrKeNRVN38gk83K8
of4D9FfIFfOhBWfU2wmkoZhabDU3idaghfu7/d0L/ljcmY1s4WaotE2ZbfpxeCWMLzPqydx8qBOC
ZC1k9oGFuwhl2KXiAFe4cUOahCDhGqzD/bdQxVI+vEMOc09Gm6ujF8r5FEEQChRbl33j6z8pUynT
yT/GvcNQtPIvR7JyQWF5X+WkzOArNNlN1P311BN9oW4M8uj6NGlPBOwtPvVyXw0RZ5mX5v4nUVRZ
52uDOhi9KichzyjZmHIH6zXdUCXOTBrwT0KKVmnsYTEiAJ1TdAbsJKDyatZB48sy8PCsYNZrku9D
v5Fs4PmaVl7N30lZBgNBdWEUQu73UBHaLWMMw8Bt0VK0TmOaPtmsCLx7qAkz7ShYB4Mi9tV42QL6
R4wSXS67EDJEJ/P9FNJHEY3pTYBZWwsIY6jZbvOTjQ4jCWNRxHFDBrLjgX3UBoSz9m/ghflHPlbs
5HrYUBU8KVu7RYfdfAjLTJshEbi8OQJGsL04rwVMS0YwN40GEPaLS55OGrYgA/WIoZ8WcdHLxJ8k
sl0PxZR064hlUrSaQQe9WfnpgGyxBsfmfW9VUp0JQGzEqNxXYLHlxbz1GEWAyi2lL/x5sJPNQtRg
aDz91h2WGrV/PzvvBTjQg/LcNjK+4NEVda6OBXXAPe/IMnK/cGRNTRu07oxYE/kZNOeLFF2AhGeV
ZKYOAN5Sf05mUsC7q3lMB+QRnnFkYahw8rja4Jqtcq+3vLd4rJscvfgb/k8sjypQcisVgtn84OcR
RxyyKaWcukDjFOuYYI/VFCtz0DB8Zhl2ohC4fk3bWrnaY7QkcWgRgeRsZROA6QYW9woiGZGtsMQ7
i6UQirD2n1k7KYFZNhJFFEoXI4Im+DkLHkQTRzbAQcbZnBZO2RLmkt5jDmpRZlCpPvPF336wKdDp
glYkDUmqWuFLTD1hReHHhD0gniFIGrCNHsD/gwXNq1BSszC+k24froS/ADkihfdVTZtIJNYGu3v2
bi+xC7keMBC3hfzx3PdvMqrQmRR+uZP129zF9sNXFjxMtwHqMwEFDnsE628ti7MRUH0Di7DTvPIK
OdO7ayEHFpoij2eCBbG1sTnJyGP2I88wrZs5Syokxy9HwA2Gz9DuZVPu9hARpzIf0fc+f5zycYzy
LSjQxyQOyxHw0gdJYxI9oIv5VnXEjwvXk35csDNRZhdDUc+Bd1yeapJ/UYF3F4F32Xq19QnS9Ei5
D5RudQx2bjQHCb/Knq4JC3LEiTNsj5x0JR/lT39m6jPB+3daXvFQJfQg9XjJ37lsCGdZaTNkYe/c
WsmLAWNsoSvKShkTFrLV275RpPqiaQxMS3if0m//kN159MOvp+As3sSTdatlqcEJmHOH9rKVVS2g
vxGbexbbI89VV3J8x7cykqxmTcBtapJVfHTkKKhW5hy2nfQcJDPpyyfD/DqNOL0GzN9YdadyAZ7I
bH0X3aWiBdGraWDfIPUEZ3OhiUOagpQvZ7jphkTkfG0C0yrvoysavcxvfU+LCZp6mAXJ4NZCKrGg
h5uaYswetwM5zpUZjaRvtcWEUFkoQgT20dM8/DvppRGZNo573MjfuN6L8vwMERa1Nw17+d8A700M
ignzNtY5k/DN22Jr0TAs66mCICYe8hmeHx1Fa5yujzaQFd4QCyiQ53kyuv1HPv96YF+u4EZDgM7o
1L+pj+B+bAamMF1OYYhuz7myaYkk5L7MBfb3LKjzC9tuiMzrRvUFBqz6V/KgA3lN5RLGOvIVJXLB
j68GqDeZ6k0rzx7K0J/V0JvYecZSlS3DKQRHxudYMzinszyp+cbSFpdpIUwO6JxThtKyBRzvQ1HO
6DrU7dDKq7SlMoyIDOom3YSnII1mDiO8/zPOFMW/JntXabFILQ59oX6LYeMo8TI9nqZlxbnlMq8k
q0Ef1JL/xW/n/5NsJSR0ai7dqCgufi5FVVQUnHAQmFeEbTwn4dzeMCwdGisnzTJHTWKNXYcPf49g
W1PlAHFHuXIzI6ljgmgIpSlsiyGaJs96e4UhJuBf/vt/nLcXZtfduYoI23dv8+35+c37KgllPPHI
GfbKPF86dkhJafE/Wa3q/um7KFdlBOaqU0GHK2u/bnz63On/o43+U/eP5lss5zP093LZMswQ4oGY
7kxvdpW3LZ6YtDwui2r4G+zpTfGdWuaxhS6CpIRl9iKOanRQQ9weffnp4QxOJmj65d+wMM/VXT2R
K2GCrPMR+Hx2rZBO9VSZxV05WLVAkh41oihLFkFMbFSN3GqWiecGsBaa+H51uvecxVvbi00i70Dj
RmlymDSuCk9ABfKauuQBGwVZ6XXmp1y9/g8042+wGNyTiK1m/VwQAFwtMORFweHCBHKZHesGl1Qx
ZF863gJ5pa3WzscXgf2Jeefth5ZfWPYaTGz0At+LZtS5Uvs84nmYZx4YF9KOIFwqRmr66TQZ4/JH
ioRxfDuTi6hgtH1vCcCz4xX9wBnFAdzVBtbb96kdHi49NQ+BmJsThpNLLHMq9dGFDJERnV9wuW0H
OobsJI/YicuLgrN1eWRba+CFI5q7My13UmnlSO68a/zRoLKRmOHDGPgX12XJWjuHBC3hoN1t5aND
F+EocGdLjSLcHhXG2yFVp8oCTTpyfdw/BuC+VILxVTMYXs/1ePrqD+tq417rzg1YXzcybC5ecwTc
5Ddh4Jatt0+nzPZKnndOw8X2onfJZRTiicAnHGLkD2x8uknRI+DK7Ltt32XDD3bNTGEm3tRgD9jV
5uouF5nOAOJhRynavNIY59n6APRDjD+DjuzEcs3hfvmTE+121jhIpS6vRkf9ptSPcZhkbkvtIwky
s1poboPR5Q992N8WDTlgaRzRzF1f0Ri544S1i8+Eds/8a+lbMjR6k2LvnktQfHbMCn5DydoCqbf9
3implj8Fu7MJ+CqnC62O5s1APKnHPwcARqMA1JuNdY+xSaC00u5zxDvTqqcXdRk4brU0mSH3G5bp
nUYCs8mCBZGhm5Z7kUy07igXdqboTghyeFyDpX5NK6sGdseQ2AsIy+4BvS0qbpEPySqPy2YZaLxs
7h0QgK2rVuc4mcsywalPGw3zMBJHFpyd8hPKmDDf8zTjYRBJ1DVvCyu84Jn4ejw44ma3K/Ke7xaj
GDnxAx/e1E0I9+POlOJ/U0/jnTtzlp9KkgsD/EEXS1wxHU1ZmTOchzGuOSFpU33MXCgZtAzAu44N
og913cy6tgzwVNDm6TRaazCl2qm737im6en6FUvICn3PKh8Bxx0p9cAmurGrHYE05WDZcae8sw/u
s85QZH9/soAMe8CBNBvTZ6FEAZ3ExbW0hE2XjCBP5I4BlhjsqqYGhns5vIYENhOkLMN1YC65+dqa
NNuifNfdHm921bZIMY2XNUbzmjj6NiTGZWK1MHvVZWgeIcFZ/zi1ti6kexnlUZ70GhX1OwiqJjay
ajdXCiRx3tXFRDslOvmVKBSJQ12E+FqQaOzeSySJgRWO1D8u+h66TfSgipHu0vO432bSq8gdaeOb
sRJe56Mrk9KA3w44leskvtOzB/+yIcZRQLDIgvF45VCKrOqJfguY707XScei4BJhwQYDXtxIfR03
3c9rC9p4qXUbyRlfXR8JvRA8Z+upp3oguYdGbWHKJ73MDez6/VMeY97PS8Gs+R43ae46f08SMY0P
8/rVrn0LujSVRNXh/82OjZOgoQVTgfNG1vTQrEhPoLhwswuPIlJuR9mdXu7bBWfXvAxt95TJnn4k
0N1MMdjf52NaJrZyCmp1sX3jC5B3a7Hh55a7n34fTdIr7gxajmt0QmBakrGxazYJw/gr4wXp7kov
w6Ib4mowA/TEwX2lnmac297QJ+O/AqTxjUAHEp/mtORTadZ4Jv1yBioLGjv+imtWdx5iucR2UAvw
ep10aDI4L+1+bKSv+29khakqY0O4tTqeNMTHO4aGUFX/CoxzJxXAEeQ0n8w01IpAJiM0C7UbDV4Y
31653yebF+sq5AnwB3z46V3npNBF30Fq8v974ypl1tbDgdiOyleXBzzfvfVSrqtTEg1RepXzkQAV
bR/CfJlciZX8H3aTJP7KbIzuSGaP13Hk4tpOSo7bzkPjnUK0FkQkVJ4Vq+XXrW6mh1U3+O714qFr
4W7u9pRHW3Cqcn2yHjnUDNKa537LLk9iBYpEyK4j5funt9+KfbEZl3sLrmv9hBuUj7xLZkPj26ks
/GO2PC8ef1Ec3pa+gJCBRJkCt9Cp2zzNOoBbH+Ny8w/n/yqFoEdqLjd7ScBQL+JLYEEwXNdv9JxZ
rDMu0v4CwfsOA5WKR/uVILgV6XeKOCKq/tQ77hB/qW+zn9XnyxPVTOuDVrN0ZDjmOmfD5suYZsW+
M6TDQpRziwrgMvTNd3n/SQx1/u3heIrSVF8b9VFh+jp4kNrCTShLgV3VW1OBrA1JI8qthGi245tN
VEILlVswzW+TVinoJRpREbvFRz1lC/9QY65tchjwqLQGNBs41Nlcu4XfqA7XuGI8djHT9BlljakN
R92Jghk4JJ8ClEUqGs2Q8erUaDKfsxmAUp6pYB3nJShHZimt1X9YS35Ye8qKgf57D4q4B7fSkD7x
++vO4UlpF7nEER50eF/H9Mdyk9ieiMR+/r+ZBPcDRcKoAfjASVNfbemTzvmldmxlFd4lpVA9hyVv
SNrkT4k8KIwMS7c8uwspdd9i5IZ5uCPOO4G3Yl4y7Oj6UBq08YhNDAvJOdy0Zyw0HqC/MdEU/1BX
5usI+EB1OfcUJuojuhPiIWSsJD9k+eg1AtDPbNbwmRJ8Nu4lmfsiTEUSmXis3u9hxCk1nmxq6eLC
aSOGbig0JPEX5fYu4rYqqsghhXDiNS/8mE38huxxJpmOHf0hDPbk8ldeKsJ5djq69VouqEEapld6
kVZ9L5TVbWklWKqlWa8wpjwrwPfnH46jX/3bF71UgiGtwqyci6II7faLbMdSpcnzu32wfYidKup+
d8CSGEO8dYUtGohc2yUDFNTyuiQKK74CFs9EZ+YamgpNYrncRH2VOraDaTSsKCJGHp2kkRGCOf7k
66YWMUMGx+E9ojKNWJQybWALJKKkqK4s9PE+NJZ9m7zaQZJnzOsU3CYCPiAN14Hg75PSJl9Ajn++
KHaaUn5zUG048B+PVyce85+nWoRFIGS7AdEwTKmohVrf9VyC46RvUuQabeMWw+9jwjzbGIjkgqpZ
dEKqo89l7zOVqDIytFhZLWqiNabgiA78d6URqdh2Y/u+tGx3qML11pLZuvBoDxj1SPVax7Q6YS1R
v5JCDFBHZp65nkz2erzYRUzqxCV7sI1GMoS3KOU4tM9dlBoO3ULKCAc40gMUE/NjdopmNriB3T4D
7Zc/SO8Mctt1BfJRYd+AZ4aEvqgy+mXqThxC+YYszFJfpY0Iz6ds22d5jZ/pXEeap5bUuxB8LdFE
1ZSb9PSZEYcYY0Gf133fsmXiNxN5/g07bhgtRqB8SEbaN43bCrEL+MGmfLnOHQ2nmLIcxI9grrAs
UxC9CHnAXCCIBxrSYZas8NMxbS+wQIdXjqXp/vES9zUmoFO//kU5lLtFJKApYL4owCyeY3ktsSyP
95lv5HMz1usQVXygpVafl1qRczN1lg4XDmVsr6tdE5XlGpUHLAmVMT3SLQBW1pITyYpcIlVTduwi
kOTU1b1FAIIS2TGbwv6Pv01ofZy+hjhCfIMRRSUzJShm4oI0wOg7cttC9M3oco7dDb8BusHbgILr
nnaN0lo74yuY+wOE6butTRqaJHqq5g99U3MxDZiZwi16ueomt67eTtD4TsuKzoHeYOT9nNMHGFX6
+KITWjEhduR+xycLJs4cmF7aNeULyXqhw9eUSqp0QKLjYpZq9gCW81heenvPWI2SKJbQReAft33o
FJTbkylkLirbdqmRtPwD7R7tOByAldY+RleTicdf35JOzAIIPYZRZXl/Fg6V1PqasAlzdEEaFxcT
d/rUZlzHG7fcwyDh8eKhgjUkf5nNfVInZ/EjuHPezRg8K1aHAuXIMYiy6jt5IblVsG0PIDf1Mio/
HiGWIodBFQ9AUj6skaPw7smd8irrLnWRPLehXUtPWuz3tfQ9EKQcbyKCADlNiLBaa9M9uw4n/+rQ
HpbEFsJFeYwihiF9vkChBp9N1cfYd3i3J8UTHKByy2psijPltoCMILDFfNVlQ2kSVzwWIqaNBzGg
fduUBY+OAYsc0xY3uc067p3YXXklG6Y5w/DUnhyP6qxPbXL2J7ENZ4d9Hf1fai8L6JTaATroinPI
xjWEX64eyvmPuQS4iPb5DSIwHL7IITOscY1eBeJbIqh5KRwiID+dU82pnPOTNtSYKtxSetTA91nm
IkB/0vuBuvt9Ehzv0JNSHqtu7qiEYXCEK6KWh6pPoB5RhnPgG4xO+gK+ib4idqbi0t2XQS9hA8I0
hyrA+5LhkDhgtZKH4GjmOVJteoYph3kpkbwh/TxvfSo8TpYa32TBfZW2KrdSm/uWH7l9D/6p6ht9
aPutj7HmMtyOKs8bICqR0IIyyyRuk5B/FBHSdFbOpn+WNm1D3vcAHTbBIt+17DzRCY1SKr9Wrr8g
ZjoPfODgqOXKJPda92ZNC/8v1avVZx4ZP903mMmRZe8HYdEmhZ2quX7BrZGaatoaCe5HdnGgXUj7
OKrkCT4zhzy/6nSjNpAVX4Thp4XLHA6CoeW87cenFR/alvgBNI6Mtz92pP8ISdlqV8pF02REFUPU
YTB6hTegtfkCaA9gv452BH8XEgzANhpAKBL+4t+Pw/XATr4O/5X/t9X7z8tO8qxU4elfSnnXH4th
mbOQP+7lECcwaUY2u8Jh6I3VWZ1Z1KDAqIV4aL+PaXCISM/o6P2c/T3X+53HhFgVHXfKyN9jO9mf
PMYMIo/C7lXX9SW1w1hAQ23KaiEF+lFd8jRREatt33D8U19EggqivLPr+y5+sT2Trv29FSfGWfd5
SPupWjpg+1BKcfua22mRZ/sfd7es6EakfAy/i6xkVFhVhyQWhZhExoyOMafOjo1JYb9dA7kmXRxY
9RcWtonSuXhudkErx4I8afc0cdPEv7oa3VsfWkV3yscR1yZ8EyHGYI8T/3g4QczF3TP1Fh4va9e2
bAeP0gp7/7h/fYHUzfRdHD/xgUdIQP0NRNX6bzLErnno7N1i5AuhiYfX3eQHgAsAr60ss3QGcGaF
KQubXUOGuKOT2KvVjahfhwpip7/gB25Q0J1Osw+REC2oSL3TEqzse86iXwHmbAvtLJ//BR7OVpc3
1vxF4o2snnIvYyVQxSmnhKOXhwa4n422mZMYC7RYQlUl9T+D0M/x0rfs/KsE+jyuyk/zwW9cZ7wU
V4XXPyNhPV6BcnzD9xSprhA/Ne+6w8cIY7UK6D0TkQvW348G5TEa/SUIYv+iLoc3+yZwLYf/hxjD
o3eZb6P5uXQTlhArckYLNMgDmW/4dTVx+3ht5dK0wkLtTA/AOBrjXruwtSEVu4ltGAHiVivQQd2H
l99DKGFKpH8AjSH613iVm8SwO2CSfcKP9+GetfLyetcW9fm1e3xNGlabK7ETMrhefmPJaI8kh2nW
si87aAjnnFdJ5h2g7aEYlK8T7YjVd2gaeboacH3BNu25Ug7XaMKY4NUycicje0yrloUHAHyXi9aw
V0TphPr+zw/1pkAZ/eO3eVu3uuPuRlKjHcqKDDLJD76A3Z5CZuRXDbLFp0i3Dv2Qm0H+QxwdFIbv
FQAYXWWrAYtTRUU67uI0w8zmYjZkx0tD/vAvTxWCeNy5KcHs4Buy4VPlHRmKm7MQC1Tu+jxfYvl6
2Ce163BUyxLeEa0Cq2llqd/pUoo7YXyWwckgM9I8qo2oB3FgOPC0vhhDOVHscDIvtBMJogGRiySe
N+OO7JAFA6KdV9Sp4U6L3yT0mew9DA8JhG6sk8djd4TKXlK8Zt7ls2l0MSrk/W06F1ZLasPNFq8Z
jKoGQsGpyN9djlNc5yBJ8rooRtFEnzEcY5Hzi5/x6yLAi9b+Ubr0A1VQkrp7lRgoIgRJZawD14i0
kjialFQ5JvbQfHe1d+AJDrd6KhiIqGoWk8UtQtwejD/fWhZ0WB+DcTtapOc2X5CcSqN+waNVxN6R
Dn71wxwxkDH0SFleebXWIfLvy6FJBNxlIoALPF/v2O2kqq6z6k1CTj04nGtjpveKaeB0Z26dFHBW
NgA4dLpouDLzYpyX+y3uLWvuQrAOYGww/WavKDKJ2BrwHQQrYwln+7biGt0P7XJxLck2KaY5MVst
4tbm1Zj3g+OlL9CA8yiY5w/PAWKeIgWktJtAIxDeVEnH64Qu+tfYx0xHn2A6DfRnOtvLngXclKAR
Rd1egwOty9DVZhwEYtPpiufQDwZ4mSJi48oqHkCFx0Jc2P9A3eMNaIvN88G8LSqAGTYVf0qK41sr
IkvkFZuLxbmRU5U0LvaB9P0uyGqFWpv8myGccEqwZMt//SatXtSTYc3Bl2umn+gHt519XGjr/G/X
AIjROnivNUfH1vWa/G70fk8sZd1AiytaW8IRkilzE9z2UbsiUjww4jZ5B9QLbOIDdI2/29DxTPvu
hgI1B+HekupGO9tcg9zENQeVfyxoMe3Yp2x5uPQHwo2cDK2KsnPpvR9nqWlK8UvJYsOj34b/jAWc
lGiIbrFeUaD/o3vYN0JrEi8K+N2MM8tC/9Umi78u+Xdq4mQ45kd/Sm2VDbeAFuya0JbI9Mtth4is
yv0u3xyJdVUxrinbi9fv7airyTCicsj/oCq4p21fz8/+qRIXu8DwJcbJgyC+OKDMNQtVPh3DMokU
5telOY3m4f9GAHACWM7nQUkPBW6sOmWQzWhhNPRQehr6/UExkifB1B70fPdMbHtRrVmzo/rM3bxi
OZCXqxsOTi8rGlp5i25vC/3og9tihLm408oXUGeck7M6RNUzUO87Jp8YqgsyFszLpN0QCxpPL6Nl
y0pi6O/9/NIAVUQ1TkSUm8AjqUaOJjcd/dylK/k996VCi3HMQnhqfI99agcsfKCucZ2FJnSdSXpI
9NPGxFScjpPDF7wy1McFroyPf8x3uFJBXyBbFpQ8K/m6U9wDA+ES7A0a0jIV15YRYjNIXILA4VXW
eDBD0Zu2SJVyMAlGeSD8jr1SVtAMBVQuD77wSR5UrAgH8C0zo8abYjxUTnpasjNjkAqX2cyGPLIa
i8dBQUFBDp891zkia/Szo7FiFA7iHwOJuqEH2WpwdXbSovnYGjy9OgfPxm0WDutlm04nKcMPZiiQ
KqGirJ9s6cjUFi+P5qYb3KYKFPgJTHuGne4E9lQ660qxW3J3jcmo1rxwu9lVAt9QHHC1Vur/fQAl
uBcKruIVKXSzn6GXEY+EQoDr4yx3b6k24ybyxvvx1m0PARLrc99Y9m3ykzVYaLbeHAH2dwKhwnnz
c+GmPGV4zR+Kn7mUATYexGcUgfjRqu8qYEUj32FPjsc2UQVQRVuOma/f3ykmYhhJMUCeCEDrco+T
BSqTNSytTC+ym9KF7/40/j2LVVrVNusM/O+W91sSrpkfiInc/BRjvLyFySd/e5kqxEGJ7OnEbd9s
DChqq2nvafg7YKXK243krFVPILLWr/Kb0JaCeL5Q1HqhxFi+8VDd3iY8wNkJuJ4ul86QLqCCf6Hv
kHW2AGJGcBuPkyJKHdTnSYI+FddEMV4arXeVLXPikUCG+zVP5Ory/zrn2YqbxJFlnGWbiW9FrVjJ
Ch9NDIpVUa2hwxGSCqfoD8xnYIpmxwUJxSe7kx6xeYyeKEomm++5v7VQcmhG/QMCttYKfMzX8w0q
UrJz88NiyG6p9F6YhVVaBLF/Ket6hsmfL5Sk0B0G9CnGSM7oXh8WrR0UflOptRa13v0NckTrXeeF
9wy7GrjNi+6eRctpuemP0QHVWzxIJcxAd1ytIe9T2wrcTgaiHcSI3T5RRb6IeZO5JtVOkcMaMe9i
rIgRAfGaQ0Zh2vvF6u+vJnLqWw94iYsi2RhEompxI7vmvLpUa4VvVN9+PAU6k3Azx/4//nr4dtPH
+R0Wg6/Yvf/WQlyLqSM7+RpVgKaGJyEtvfIfQZNgzvY2jP8kGAEH042Vo33gvTXZ4rctOLg1ECXK
XKse0wcn2trm1hWbVRBcqzp2/Vs+Iuo3XRaxJEXtZHasyv48j0y2EQPtmAdtBwl48plaYvInstMl
uuU/2hR0w3KXCDVx91o534HGJCtD6k4fb/VQWhSouDYhI1tdUNr+06U6TaTPmk8zh074WNCT0FW6
jLyWh6APiCl5ewWa8udQSwbCBnwoBTP3RubBii+ZELggqgQOV5euLzzVrDvdjNVEzBZQ1YvM324J
6ydkmMysX4x19L7r88M91nhKv2oP1srS6OG0F2hZg5vrvz6sKSvZxZqHH2OBz24W+P9Pe5Ddguvx
leox0Q9sgoytumEuZ18byUT4ytVz0mVgf+IZyu9L0ZXNQWfDbuTcAhbV6u/Pxoz78eNUe9lWH7I/
aVU6Jb+S7w/rj4Llsal7WwWdSawb/H+aIW/WsVyK3WslNkWxlhSyM3HspWWpmDMpVWxXWFFna8CA
dseEjmienGDVSO4zf9O0JGsn13r2vU4JiSmcI93WjNF4NGkWdcgxHT+Z+u0Cvld0Q/g2Gthp1Eu+
XUNFxDUh618hLUSuK2rM1ZSUvEbnB7fis3jxl3ufe7BlS9b5FTcu1fX9byl5edpyUmbBc80gLwbx
x0tQv0PKnHqfkpd1N2jG6+UPa8+HPN8n6bFwZ0S7raGYdBLReG5NP+GFWjF409dov1wSMwwGsgmd
mOQcJqV0xA4xvWUrrf4M2jtS/ewWtzH1W+7HMHEThXGQ1c82bibI4VuX7wL/mlcqQtqyNduU7kV1
LdX5La++ejGtX/E8XSf8yzJ+Vg1vibFHFS2BOYmBe5r8i5LCSRN1tTfhhVuwkpkOvZPeWvC0urhF
7VDZJ2v/Kxld2SiYHGgRNkoRP3uIzHR6s7xWs9bginx28lfxiuNZPr4ib4PwccfKnx+mYDzhumPG
WKVwR/N31+CL5YdzxmDRDdE+mP5cHdiQUF3umgy3XsxVCAY7O6z6axlCXIaryebo5wQUGymd1ElG
V2XMeIgw8al22a2i35p0OdeGi+A3txkQts+sfQPc/lvi9JG+7J0H1vnActqNHw6afMVzwDU64u3Z
eHt5krGNvkS8kMW9/FG3xsjuTWUPdYj//yIqnrr2KU3F9Wci2pLFptBtXhwIQ0K8XUIkrxcTus63
t0FKMygXHGhRcZRlScJ3O6loSXbj80nanUPJ3XbgDk9fYkPEQK1FPocQjqIctPCFFSelGwOXtrzD
y4Lc2iVZg7AGnCqqf8qYGyeCyr4sWR2ZX8TiWq8aC10shL4NkW4MoLf5LhrrmwaWbQaItQgtpesq
7/fZ3OZiBg9xTBYago+aVQxL3FGsJ3LgMsofXbBZFvbtJQG8tXNs8rwX2I8LuajP3DDfE8o2CSrx
D9KG4VxxsCkirqXxNFPKFrsz6gdReoQVl1enOuL4AZcqXNVxTomZKNUr7SxGVq5/XOPHlXrR4o4H
MzMAqcXhoU/NPu0jNKxr7g96ngYlYQxXwcB64Rx0iSJxamQUB3AJh4JA8C2HWuFzWyJ7iXxLUHa6
0EsVqSfLP4BX1bXOCTIbekFQOs+eyCKgz7PLe/kDVoDXDrc0f42B/8cQiXuKXN/M97BXXUcuNuxG
fosS4P6WO3SvxqgiHLqTvmApFdGiFEH8LbbasLuMN37qUUIkbsdhaU+51MLYxAvqFfgQ3PSsfRP4
+cZfI46p0Ha9fZF6zzyedHahkbzgpzZdi/e8RAQ5NegviM/W+tfmLKPoqcUuDDRfVFBEysyoXyF+
j9ix4vlPw9MfCuJ78aF0i05VLSAIcm5FVEOE4ZZKmQLac3qiAQxVPURceKvBSNkm7DByIIEBpksj
mepn+X/ZqSWaIlUDYAT9HS6gO1Uypm4sXbzuzKcQgWk1JMaXasnqavUGdGFM+ayb1Q1/JuuNfmR8
catDZNRWJ757MhtjbO8VE4egWploqi5RjJaa14aLM200555dXifgwXsPE6Y14YiyM8nb+Ivk/Lkm
02IO+0RStYmc9ALpfEXKNewuoVs3EBj3gGeZtyPXg/xW7aJDImACGqggXLmxwV3ntU8zdFyh0355
1P0+RnWyhH8RHK15QiRhGxJbYWP4XTpzHEod/M7GwJ+b0ro9EbDqVlNqVAPaATz7m4hqvS8QS2DP
l4xpoz7hWb4EjzqXJYWw5q9nHnPTGHrdeAsMtH9OeZWqGIDZP0ptvqu1anE4OG3+3PHv0BB1sWZi
VAZtPvvqjKGkV6wny9wLChjn1L1K5YY0Vo4KlMH4pGnLdf+cX031KzLmxUdQ3S3aEFgAThG/G04M
NLfxx6/N/kWRROSqZfuCOEYWnKN9EHwFZRbP6TR73Jovjt2q55kxEUol1pqYEi3+3jjvdrC5X1f6
Fd0ladQDd/mXtSmtMfbo8ZPAVfjCETwsWWsj/1bjT6my24Ps0Q1MSZizYHqc+CrJ5m995zrvpN+v
ueNc7U5dD2sQKiwDQN8ZGyWrUMFutZoSKJWcvKdoNIUBZY+jr8gz2epLLv64ozcgEKkl0xiM62BH
zpd37A3NEgQLr3LeWSp1KNThZ3oDw4A1D+mMVx7jRT3y8I/JPivEHgDi39paBsy6pSpeBwduef+j
ZYI12zfPKmDti1T9EWRP2sPXRZD0lVZcwUHtRAjdz0tkj1aPYItdJ6fdnDToZJ3rnpVyJqECnwly
g3ct1Wrt+HzDctfBnlAYH/mZ/8sXUN1wtKiuC/O5U+xsA9yRk/odnPF5/D2q8CBhAccpm8lhwWa5
LndKnFjRj5TsgZk9n1BDDatgBU9pkNVG/V3L/M5SL/63YBhk8yxQJVnmG/EfKTPr8Aox0cewc25V
Jb1F8lLZIz6UIEfbZtqn4cRStV0L+ZfMDzDBkKOQ43I38QyGwRueggmJy2EAE2nW31cInfCVkfNw
0OSnV/0WFosKvess8DYev2lRWOlGQTJ4XmVUuXZdn5AFTdOS3HtwnROc2AP8aBlyQ8Pzv/xBH4lk
xHXGHSqsr5O1YWD7hvMlv+dx2lh6K7P49M4ATn0xnyf3SboeJLC9uwBlObZa7JLHwaTZhJm/QZEJ
awfgbFLSiBl8O/aoSLE/+wkoxQGjAfHNtdxun5Lid9cKsGcqkYYTnns25BHlZPchqKDtZW9Xp6Lz
bqbLwtklvrmzM9JB6GSjEL1dXUt/HxCeN/PgDDFuIq4c81pc2vl/n+1dbDoJwfgSpxv3tNiXqstZ
hlXIffAx8+ASZi2My6jG4Kxd9reaTvqsiiapsQFGoUTh8p8dzUqh6inODg0im+FYrGZ2RS7VY+CS
gqHhvMf6zbvYA2GZA2+Kre5XOPj4uYu3vPy9NeZcdSbr9txxiRViV1i1TpqxrjKd3MPFfpp2hdYt
ICD0NYQD1No2BtFT990znrf7a8LpGavoa30qspp7k4R6vhGsWcpOKVcOibLg1MZ4UCYaeJ9Oe+rg
TwHCuWzuKJZIFQPYXa0ADW5Wxc71eHJ/JRzR5BMnN5MAlVmuEK39G9IdkFItjii+u1086T5uldvP
gUpmJ3BVWzedn9ZD10BbcVpTAqKiVCAsZJfBARv503oIbZOwYW+uj/7wUHQoFGU3ZMRhFF/W0f04
dersZx+zWplm1rmug4xHU2R9rX+Q7HdHm4bKSDBnAntsDs8J/efo2CO4ZjOjrAWs8aPrYAOkRhCV
coC/1wj1kaUpwSHcbt88eUA4lvDtqA+t8Bf/Kg6DMJzMI8DIahsyfC61a2KGISWg/7ucyCXSGKBZ
Npw0m9F/2epPoE8/VBjSx6zzlNsqKih9PeZsoa5oUiGcZE2cyvMnyQ3NQRP1fK3Aa68rzOH7KrqS
LA0ICXiMLaV+AJbm1jOq5ufnkyumxh6Y3fd/4SVWLmKQy+wIWZScXyOi64dJP66eC0XNckKK6kr6
ZFswoGWycCDrZzDDIW6RNEUWMqDzeQxUliJdeO4EM77VZo1Fuu/0t5nQxWAczkoDhkgRNOxN7vBu
xOFZmJnkiWc7P8Sc7Y96aDP7JsmnPbGEFdVbOtkVjdELCpox81N7q+FpMmwGJv25fRsd1nNAiL1w
LX3rPYGMwWBoKLyGzD5TNDfuWbVcvAow70a5VfhdmsVnP2kgGXY5/860gZMeEuIFxqcyreNynxC8
oGAzCM3kyMXdkv6ewYu5NRJExl4M2whAVXMfi3beChQcSmezHdnpotDJLkaF/msObgW+1mQYyFeV
WuJuE6pLGVNR6xvraVvcADkr0kO77ENTdEoIhrdnyKR3G/OZCabb/MkAbSfFjIhV3SGFB2vrEX+a
BYMFDW+FXhgtbIat1bP8iNl4yk2Ui5Pakb3ZYVhE8xICsjnWmCVfD4vZzNW6raC+Pg7NzErYNIIy
4GnLOs0pkoiRjgpjENaRDy4I+ISwGgb+uuSiRXdyCbPoOLR6bKnCWs4VF2X91uORk0lsy5SF0AuS
2OtsFN5gv/1n42EoXQ0SA+n0z9+ILk9NgmpP4wOKO34zP7O1rysiwmS3uM+Cqt42sCL9+iSR/+NW
xsP0i7AQgFCFhqF6+yT+hp7FapI7vCKczKD2pj2e8nGgIHbVuxvh+X4emTu0H08W/HZpc4JpasqW
bqln3cvLpYZLiDPHGN5IyIbRG1oWwRUgR4wgPhfUSQJa9MQYJv+5KMwYvYZkfEGnovs0EXnOG/z5
grxobIlrRssX+He2NkbOdWzBb282BdRx2V9ALPRsuqnt+YWXvniO/60BsanlbRlzJ7xK3MdY7cuV
SZRlju9K9kkFeQaO0P9dumTZMmT59tWN2+4iJhZ0vrCbjNAdLn01LLkKCW1chkvGOCZ6Vh3fj/NC
K9Dv1ji12V3DEozFrYtex/TQijwsI8fnG9qEdhwCt5Bwv/9TbrlJMnB+F16hsCC71SlNweZa/mLd
N0zIRQS2ZeRcGtdKwUGGxb1cCsm1HSKom92inZNdWY63N6foFMYES9OPxsEVTkqfw++NLtkPYhNM
4DkHnmWuRAMaarJefdSsqFc6L3JkS/ckDyeWHgwY/dwWgT3buvq7cnt9z5r2ElBrp3BG4JrXkrsa
sght4FIaxbNzmymA0Y0clPIvJdqo6pryi8GSE8qlLMsygK+Wcp4bG3waW01jKWrQ1mZmtyfHAmpN
879mYviGUZo5m358BgIbsUwvZvM4emS+x6z7TYY4UhkI9rA/Dltj9GsDpiIdDHMMlcpMLDjpfdN0
FjHedgqFbKoI5VW6qPVWO9M6afmWQ4uupuCss9Sx8yIMtYLOENeZyiQi+fAWqvuxr7e47LvS2Y07
wrYO0PujyYL3roJG0aZEYusNxSa/Zv8VeRUhi9KiiXMLoaxh0Sl8k/v7fDsYGJriQB74tTefzGts
JFs7iZkqdeTogFf3WjVYudvoRO8mIl7meg9Y1CG9qmdD9s9g/wHnP3WS+leyxWGYGsc7TL5Core8
yfJVTJ0DRZ4uW0vXPYRuSVeiKYbJpD05y6M6fUipX0qDKEBzNJyj6FDpcdd0enucIdpm3CSDgkUk
Mo+vVfGsyHFxGgVkiD661Uj+p69jCFrmUsx9qdGprj5j7Dq3MMIc7HL2dk9hrOWw3teaEJF1a+B3
gRhS8Xv7UeWPajKDC3Nw/hak1EkcP7B6xzp7dt4RA2YZJS9wE/cq2f19r3ZXHSB7zUiO6Vy3t7KW
SPFv9IFS4T3x8Rdq8v6a3e3qJzla+I/g/aSD0j53XgqyJve32Fv3o9qd5OuxRMOUaLlGUzVmDO1h
9Beq3fbYRCSsVFV5bwfz4Qezc75FyjU7uFgVkbcnV1Vl0Y3QthOrMLlF5r+TdiKGe2Y5eJ4uyVGK
NKr0lHZpxUIJFGWqRNu32SgbT7Q9hYMPXXBZXw7/DMPY/s0qqfWxWQxS/Xv23+dOo+oBDXH2jaD3
8JxOQUWrCi/VGP2niaQN1O00Vv0Jww0MxkWqLD/1RX0lABT7fUNhlQ2RPzui6eqNwB7+xetUZESB
B3s8vmjEQOYtRGmugNxICxK/5oEzFpSdbUVxKf10bwc8wjyc5rrkxts3kOpDYJu+l4o2SWVojCv3
8cjS4mUjB9gsK4QTa5Gc24nDHz9awtpPsNcwRpV4UKLUUQ45OFe4Ubpvu8p1lI96aWGtnII9ik9r
dXhoHRhjt9XuY20IurjqPvbznLCmAe7md9MH7Tu0xMMrvBYtDD7/a/+2ha3ywnEv+19qOW1Jns+x
mL9tUyPZc/nYesRaICdrjYFvfYqOBudY8ilXhD3gmUZSnLfcxhgtVE1OW921k1GVsyqGaW+xT7wq
IkJ2G0tORLZHC2uFGL24CK8C6tRJ/po2wmAuueJn7x3HYgZm31BJ6iPCLNC5HZz6f6IdJHV93bh+
ar1XG4vPZR7TrURweob2pTdK0hXCWC7Rg53krEorUmvPpye7aoDKXo9ZzrfnHu9KeRP9lQF1S9kG
9recwoteNAwHiNYFlPfPujwKfWH6KSEICreB9Xl4PVf+Z/KWes5Ck5jp6pXsbQdQ2yvaZvsfLDbH
/4l3VVFX4tq53gtt3dGC9NHUGZXiDYC5x/ws1fiw1UuaBhOWQ0pewPbG9uODGFa7E2vBaHuQpY0v
EOgLig43K7rGRoAJjcCkyuuMbWqb5i1fI3K10KQnDwpOiUXL33FMYgbfZ5RS1OUnHvd3dfE1Fzdy
tSJJTj6dpDAb3NGQS5AgY4GXwZrf+2AxKzh5U9O76DUWIt4hskw0kdEcuIaHIWMIZ7AdQ/l9h0Aa
Ss3/HmonYleVQ/OzWAuwjQf6qXaapnObDDOxejXM3WAu8ICdQbIiBpzC54L0id+AzE67Ha7eFk17
+JznCT1R5te84Ma0TAqVBf6N07lt9SZLcHd4ouaYlfPOGg44AIaaTQCnVmpJjoo+snECGSZ/TRF9
BnbVRMoiZaX/wQRKayF6xZTFr4sEblWq2jF0aimhxTwgcuUn4T3vKygtdlaru8iSi9WrbwPCmt3L
sdi6yMcwqh6poSGbvCdt4yF00ANGMAQWxUdIpZZ9zUl8mksDqVLwQKsC1YC10e3STtQ3lSWJ1BeO
jLfyNimVIvGG8ZSGoC1OgaeaS+soSYy0PdIXpf5qjcJ2gi/JHsi1j/42V+hKV5bunDf8Vh4jv3Lt
xxrH86XNmeen6U4nCTqID3JFDx7kC8HFvUI+L+WvLQIq3NAB2DI/nAiaxXnNCSTyMW2KRIc07He9
BN9F5uk0vuEwuHthB1T9ZtwtW5PSIYC27Uo+GuIr67vkrfuY5pef0qnwf42dnzoPeKdbL5yuTmi1
FajzUl8SjI533KFXUW7t0c+SDR2C0nPzaJeGhGxJX1AOjAtHa8EKTDa3gUidLpsTSk+kpRUHA0Zx
3hBKyPLRB8YJmXPyfZg/7Z7xvu/aRTJmJlpnGMTAQaCT+Ja+NRkVuunWbk5Wj4y4QyGwQYSS4B54
PpeKaDWl6+ZSGqlmPiIWo0NDR3JUprcGLD3Z6mOwzbfABZzB+q5yLZ9Xqxg9eaL2Nf/egYFUObKx
CMQevJGp60QxLpzmUL9rVq33PuyzQ5I2Ye08jrwzdWqed8Z8aPYFVriNyDJW+25u4Wmzp54zI5hs
FDb+tuXsFOLr/0+imkR3dvJn6aFp1RlL+dmGS6UGxf93NeipcoGv662hl6pETp2AbcaXaJKiPiwU
Y+NklFSFx6j0JxSWc4noQr2QRQsnum7sm0x8ODcj4K7QjJxdSiBjdqczU9dljKDCD3mBR5uopAHR
uIh7Ib+Tmge63zMQ7bOg2fj2qW09QgQqX0/TLSY8hM2grAiLXmun23h0FdtU2nNs0/htxYammxAD
vmnAnRKm8s6buGRF9dCWLfZxVEGJSoO0hmFtHe8HGJgeorfwqyQkxPjihW1UAVUch2CqoQosCmTi
pc3SBvAnuqlTXXT9t3ZhmcsFVUm4TAmJDGQ3OuLBABap4IAcMJK+W1tSADxdm+TehQMKeGFG1p/3
NgKuCh702HOX1ZhiDIklBbysMZFZcIwf4Nk7qpQQLXUW8XJUhlh7nylPRr3XIuY6oXszX31fvi7a
g+s6Pv5UwbdUOt9cKG7l8hHCTDWS1PU3WJuoMPeUtJJLqxRrW183+P1K7ceP80hYxsaTqr0dL4Hc
BzqT+W6xq90YXSoNtOA2/oU55BE/A5NXLwCsfcW3PpfOmFNFlRADhrn4KbyXgpTvPzGqL4GwxGzA
lXzeRxyye+Ef2FEIrQ7bGsBSgGoxoEi1Tc81Ch/BD4fblHyUptXmbITToxETyGznn1qw9Ph78eAU
o1FIsHRPKNdw6kKqZOi+rGobeZE4hW9YWAEPM8Vhmd2ywkp2VAGpZkfNfBk1cuHtRfNR4IAJjFaG
57oQ+z/8vHzNN4znaCtlIBgHXGzHSmE0hweVQIacukchH8JKOTaYMCpyr+328fPcVIb3/KIpfIft
gs8IpFgPFgAWfJ4odPke6yF1WWrd2aeYKnXYy/l1NhluK6tJu/MzWONqtBnoi8WC+VVD7NtLdu9q
lgTt88IaOSQDFPuszHJRwJFTazrlxpcYRZYpMIJsQwSLJblA+PvMmutH/hab+xtexTkrolkIL7hD
YaYb77YEKlzCQoJn1fVMArS4wu2haF1IrskUuw210BR8ePFOgA0dXeyPukYbqHt7OLv7HtNGVlw8
7Ym5X//OWXG5drZeEqRUS6vWsecywRoFS8FlsmzgeUNwvO1fDjYCy/SdjMdRSexBCvBPpyfrEFVR
l3BqTZKeJuSum1K4gE3MMeY9prlrpuHACsqosZnNWJ5z2eAKdOhFDnDYpj/6c+gbkRFiG4JUpyUR
nrBrCf4yEL3BaC4IHFkxWHv2aglserVhf+mIh9UD0MaVrW8vLxTxSZfFmx+5oJRlgHLd+5ESq+90
Ok9T3xPPs86dT7AOUtV/xZgXe2CDodE6v6XRyBvWf9uhx/ZywlpfBI1kh2C3trnx/OZ8wjgUHUIu
F5zMqNZg082yAVR+rm8rEl6Cj07nOnAlnLrwRJv6eUGOWabWphJ3kS4hPdhHMXCfIm+bhOnRHzon
q+lXPDh7KwO+lnlZQbmKDDFYNQewXVQnLGVyoW2qWTufr2aoVEwXwUom3pK3DeRlC2R2HrS0F1Ou
oz5FODuEpdU64j+y8Zajc4iHEq96uE6LKsWB5LY7dAbgAjViwWeNB/OU7AMMLuKyJDuzOxtfDTAS
6dmzcuFfxs/yQyX5lbJ5jKcjT2cxRlsddlZkvcCBoISwUJrwEX/hs/QSgMi0I7NMVbDFoHoQPSEX
FF69ltpGLVeGRUuZ/74IU1vxkDElTZmRO7jbPoNUZP86ZvC0UR3oeoNL3H0OFL4vR1avvbouO5Zm
zfd5Lf82AUaxuFC92dum26LcagLhrygH2MtHdOquMJkC1ZEoQpytLX2MrT0a895fTniP1sO+gDty
AYQicqtrb45E00nK20rnnK8O6ZEv5Qy34so0tkw0oSm7YcOikDC1Fw6meT7E9swNXg/FhHu4sWon
9hplk/nNHVddsA2NbTBvawIGxBsAqJmQzwc+wgAsbsV6eIONB/pHh/uiBCKvvA5SIDw72fo3pKZY
G1m3cQQ6/kr5Ob6eLBGM29PKD5O/7nYsSyeMXmLrhg1ex+qgNdoQ+JyaMdlgCfx+I5m5D2Kua22M
+rEtDrmc5ygidvqKGbN0IboB6jDVE35DQFCfQqIB8jURr39dZLqvnbot1jl9cGs0j9ImBt6l3ZqQ
0+ttfNHbtQQzYXe+kFkk/0bOLAecA7yDP8QbTm3JLRFc01VOr6sa+LfR84GmBmPEoe9FIT3mi2G2
WO5kB3ICoXKLbmdPIjkO3xI/gpZYn2jjEoaMsBywurSp73+q2FdBSdXEQcSwFlkzy3WePpHW0Wnl
LVJYHhcKQDD6W9SvzJJkv5waba/pF64tNf46nX2HglYlRGAzj6LVwpiNnouA9yuwuN/dHaxF2Ki3
Az72tk+qGRim3Ac+Hzh8qwbnxgzgkp5mJBPKr+36BCR+zWUGvkeMOIbjGbWrais3AvQK9uvhZcm4
ifgzdbT+pIt+rExjIWHyUepFaLb3qqHrtOMBJjSHHDbVU8NCC6PxEsSYXyFRlbbv+LSVxrkHPJF+
xYVgziHJqlCUkye0044jQz7iAbiQOsYz+kejV8qWunJYwgPYCCX1Bv23w73wLFcUxHdIXhE3Ovzo
kUgeCuDQ/TczDMVLb19OESqMd8bGkS6IXZRV2jB6CMLhnhsk6iqpkpLOOXrGduQgTBPT/hg7ETYM
Ih3x4RqGLXKjbzRxUcobVU4CXNM81NuRAr2ajvyt8tacfAbM4rCZuwcKRBMwGafVmWPWX/MfM98I
KLPhAGOXPUNRiiXRCbYcTQOI2GqIF1HtQ+eVr51DH93TakLGgaa4VVe0hsduH8sXzxiR5o9gfc2l
u5IE4wwlqAIrBYadzof5gXGn11wrKOdes/15J4dLN1GZjOPXkG5oH7m8KFxTa9JKkcx6TQ2qjwPn
mleodfmK3TLTDyLBeYz358jcwpmvJWZz/hlNex+b2YcMk4yAsz2pZrgLZtgUzgbWZKQG0L8dcIIH
/dqCpYi4KbMpvOhEFk18JowLkhUOLER7NZTSk2IM/AuD9SrJ2nPKZMux2PXLr9Wfu99NlHPOpfFa
cXvJ+wW1khfkZgTluPEtlTfBeLjKPkhsJZXzgse8uFS64bO8EvWRShRYI+N4pt36/E5w7vNrdGzd
g38Ld+ADRh0vXlRFv7Z5byJGTxLqLpyaJp13lC8kicaSdWboAsqYVU23LxYNWSBcjvCb07lb5V7X
BSLnxHWX0nXc5bdTBx+DwpkLHuq3U2BJcznCOD/IKqyPiNnomHrqLQS0QoFxIjm1FnYs52llndbI
TDK2M5pEbLr7pZYhjzLrNWsJIgsW/dZX5LpEOlgOQ80Ov5SWu9eVIPxvFclMKhZxYmjxSgPAbM+S
EWLpnVPePpryVp0NxdWQuqGhRYCDNOmPIPPCHrVrOAES48x3Ql3imMZhQw+6NT/X4HtcDWX8MdME
iDwsJ9vqmT5a76UgdshTnv+v3qQDzBNMFJXN/5DkMpXVvs6e5tgpNm8VzFc9QdxaxKGVcSGiWfIY
hG1xxCUrRHdvVrpZ2p7yRgoIlNso5LUkwpmnkj7xfwgmV8rNK8L2btkUwar/e1Pxh9VIqykdlMz6
SJhFSHgetr2tTtGfEtzEISj2dLNCfqNhZMQjECiuJez7PzFehcfCUORW100nUBtvyjNtRIV+hz0N
L3P4Y8PB/tqpdculNySJLcOsauLhHN8GqyCYW0cb2x8dlJ2vpJDxnMtxpu0YhzsU+qH577/9+lBy
qSRV2Yxo4+p4w+2MbHLaGn53uvbp5smwgpLtJxUQTltaFkx2VYmn4fF1WHBSRfEvgIRmksvv4DiB
ox8sGcvO/OCFfADpaXLGZJP8jmV7ISp6OygefVSJxgH35B7XtUfeB7kfuhiv52K3Dzkc5sBWGUub
wkGx3kZKTk14xmseF3EvurKPXehCkvLn0DBTJOhfxkNwV9Ojg8ut6FUdmLbgsd+7qvQGnwwKIMPH
5LVjGLA3VuyH/3P1pjCf2iQ6s8IszLPnuNl1BAuePEiX3eEHMKHHleAHUxZZd+1fc3H/8lT1shoW
zWkBqYuB1Bgedb5lAjsZyXnTGJgfinkMtGAYeWEsl0yEfdSpq8lbinrC0dhVSPE255rlJNpoKQlu
gXKJkkDwv1H+MezJmwVtuo+PxN1VjKNjcEiu7jy40YVaFO9RNUiQt5EJoE/QwE+wyj0bpJ+7gy8K
KkphEi6aJ8yN+RkeUrihTJSua8pLPhzRgCGboRnlMlUqD4klby6drptzslytigVrYhQ81LLodZPI
vkTVlYGtXgb5bKjUQhmFV1DlOmP4XDVlNSPbnzq//sO5cHYq4qyEfA4znp5uGrpuWjX+LwHFweo5
io6tjFGyi9HrBXh0I5nEgxE7gEWB5A5/paQcYIWt4imkL/hPQgM8ASaXp7/KJ/WgHIvZKMpY5mon
zBMr8BCZK8vsw4MFM2lWx+iPafhDld0j6NKrQWo1yM8n8AnwcEIQTNshw76HhnvPhGyL8VO853/o
YavmioAI3UzTmQIOUEymeyPWORKImIxyqGU5Pr0vpuBlk8BkRgOZlbcpBcCedQKiKUoCRDVAEIDq
uA7CR/I+EE0Zt7WzVoL2QPKwjw51+JFGa1i5xuB3rlrAoGZY2ngYyVHnJ/Z8+AhBlqPbstm3BLGS
Sx5hhU522o9vRYymgH6OjIJulgQ5OWfH3ihBETkbj2nX2oB8zwFTscjn2qVqJf0X5WkNBfz7wudw
zDIpHs+o5HxWEwd1xPj3JH5CzJkYFDkVffQXe+80PD0nFdj/uuLq9TaAAwn3Z+9gpJBYN4oXCXqD
CKy/vZZJi70vJvpOcFtnqAeCNuDeI2ulzjD1frB+yI6hvOW+Cehq9Pb/kZgo9p1Cn6mqxQXyjzaz
N6OjsyKqfKm464iCgJE9MhOUciB7wY2MbNM9Rr87sVrK9OJcmG49VyL7QVkq2+Nk49qBytTU6+dF
zCIifccGStNNzDujVPHkFNxjrIpjRSL4IcTSKI+dIiXKzzTzIdbYpP86GlmI2rec9QUyXWQ5mFV2
S7Rf0sMCKYpjHMY1UM65EEyedXVveV8Thdr4dUl4YsqMmu32q40oa59yLuOBGY3cBAPKODtkXf3w
hY/gz9Y020DtlQckWfgjKEaJmxuMKkz906YoEGJkj/VUfCcYp680m9TIBEu1WkszdWkGVbWm4PbA
iouwV/NfwFLZcXWROpU9qR7G4hWhyAPwxX4pYsXBErNfX1U9L6ccx24ZPug0O+uzshR9hVUoT7oK
q9GF47Ta5FtZ7xajzxaZOnk6AeRncr4yOAcW+6AcOJvc3BEcfPV0aeICEfoBknQA+ozu5yiGINqU
RGvIrG70vL1RmUYte/NNVQ30Jeser2Q0fHcC+buUi8SSM6gNYiOAXJCbrOEPVMomMnBeBP5HPzkD
BzoWzgRYRyhSyM148iyneXsq+xcdKYeCmtVmFSnoBRx+m/TRXFD6Jtm7ksZvBdKQZAo26aJBaeHk
SrJmFTscDpTV6RGDO9McsOz5cg3y8krfAubzadLVFQXoslMR+vcKhyYmpyRxWmGfSMk57URVVLM9
uHcE2SnRNSr1rEa0h8DT+Vzl5DPVijOpb9fQXgcuWlKa01FyUeKeDTUuXXMaLQpPxUWfsk917zad
NmNB7KgFNdDKL5QMIrZoue7VxkTIoDWye3grw+s2AL/UDoRDQfKtywz6eZ2ZSfOTtrtydPQmgJAd
smnJpS6wv/M4o3hFISqelVH1QvQ/I1JG3GZo+cACUAnl2ia7kMED5nHDZ3QdaXIfO3/A3D0qbGLY
Z0cObVJKL+wqR6ftBG+vhvV0YllfYLbsqSUSAaHQNbB19VBst+tVQI4ztdd1OJEILwjvMVhqTDIr
UrB7XDo4Dt397KQ8NmL7HSM43xnIFYH+lHxTHoVO9BsvKBCKe5lG2biL4l/kF43kKb0JyUDHXn1+
bRo9JBKRi34aoqGm6R1qTtPzVg0nBxAF6nwssIRudooJArvu/CB/FodhRi3KjNp0YxompHJ6MqE/
hQIYEiHG8AslNqWUXL6EPOndr+qSbcq03UDOhJMh35wuAI5gRVjZ6Q5INPeDeV1S2wy2f3BMPTvx
ApLSMd7clrQzF6eXKge16OZllXr6Hn49jDL7yh87ugNENq/3qUX7XDIuYvoap4CU2fqn5yigt/Kp
MDLnaaivYwOTV7R3cTLk3L3hV7Lb0d7uVZKmgCVphjrmlmUl7IzwnD+RpgyDs6DgyJX10EoEABjf
bmTGPt6unhK8UmMaNv7miyxMHz66u2YfHRjqlX2uGO8bbIbeFAJoYfQa0wUeUTdAakZMav0NBzyZ
fryHN59cJwXWvY6ZqtfFXB7qMUdX7GTIkZDZueGXbChKZ6twI2L0nfpNQgGCNpp/XLF2gd0Be2ex
gSEG/wCAYYnDblCfnQwoh8v5A2Zg0dhtf/PaYx0a988IqLvonaBaKLZf/B6sIZ4xVPGIPO/a0xW9
/KcLNJJIOwCNgOzLt5aUxg1KMyRpB1lzebqpQFowFGJn/9yUjJb14stsoZYE0T/81LpVEblO2pdR
XXGb83uGwT7/cK072jmd/jRZGGVaCt6KEn+yC+3+jSD17qUM65vFzXIeaIGr0RTCBBc4wBA/89pf
SaGuugTVVM0PRdN9LJTtElkTLEBOPbjslwRgfSxTSWrSbydsc81hghFMCYr5uq/Van2DLnLDXdeq
0ECDqz+2/yRTqB6PYr6j0QF3PUw5VYOWIZh6hDZkefKyAkglnniK7ncIVoW9H5mZawR5uqIxfCgT
uLXevTd3P7Elk0u9+S3pywLGafo+A3AO7+hTgKuVWrq925pnxuwZO6OQDV4AhSKvCCk+gGyKqUbe
b3OUC5OG7NbC2dOZLi81NPlPZGmN7ZYUtjBZQoajUyjumCJi2xWvtSkSaJOHOUCkp4pfKc44PIg1
kJjmIQkso3Piuw93+kULobnVOMZfPrptW0e3Pe5XpPxBW56nDEB+TfBqgOoq/bAqxTg2w7KgWEJD
4u2uSnYWmaq5lFNCUU7T4OP5gjN5sS+XlAoYU5TYKujhWMqsof9Hc7DmJHQj95z3gqgXETmt5bhM
/Wqv6b4TWJNbFEoYdRkETfCSNm4QvOuGIQYKZe+psGvqfz+kI+W2pNWVyckMHUQp86tnoRjd5McK
c75G+R9NTwjn+uXOWR8l2vewbKTmFsSvEsuDnU8QkDby2koao8MUVKQbMXU6BB0ZmeIW5ryFjQQg
x5CxL3vqtAXTHmR8//kliuHD9ejx1256CYKYetIewhmusEUs5RxsFEuGBhqiYVbRw8oPlagcPnUK
Usiz5uoaNCB0IO389Nr0ebKN+qwehnjBQNfM+8H788O6NqskTjHFJqb3PLQfsWcW/znrrcD00DMh
nhOWohwkkEp0s493yRlRN6bPbOOnASTAr0nw5D1XB9ak9Z/pi3fKLTRozatO5zcyDhaWZgR1NhhR
OlCqL1W7VQLbmJUO5FDh7vUTjuZSQINuBHIy3yIrY2ln6wlPNGEXgq8X7hD4Uvb0RKuaTDDuP7tb
V6THdr2i/Xr1vP8DVlfl2XJlWEH98DN4Yehpe6fC5H+EKusbUCReIKpuE1eq6qVFmVWh9EvnNm+2
lBRrDJKVezIR59+ZzSa/bAUi8WFY+gEXOzVhpEWYuGqDroHbFLe9mc6z5vyaUYaRUVkQnfCU0cZ8
Xv7fPbpHJTY/JJCfAtdlKj8mWXumsTF36V4alE9YYm38jd0lSs2DJaGOut/45F71HoqG4MTn9Yvf
WcSKDCZyHSB10oq3txbOWeB9Y94GdKP0LpOnZ4fxVMAIND9nm94n8GW7jPCvFjHkNMB2dUs9/Sxr
q4Sss6q2qA7Td/IFmygFZvSotIk8pLWev3BS+Hyb5Y3EFJNHL/X797tE27hwqmr6fZe5Mb6Z6ZLu
6mlH68YrsAs1Y/8HV2/m4HaM4MglhgQSUu3VGl0XXRie1e6u8qPRpsYTD6XAUveVA2YybLnNyYkF
TkShHz7xEaFPXm0tP5OAwlhwocrz37pR2XhzCYecRmn4Pn7xPsMM6NWqXL1C3Jt45W5ldtA7TpdN
phBgau6kJFO4plILPRTNh8FmuSJ198vn3XQsSk4hCyXt24r9N6t3FlRc5Y5a3jNLvI4try0Ox5YD
YMUsmD7eCn7s9CtB8BdbpIBQQ0olaDlT3Cj8ALyMrCj++h1JcVgGNHSY5QlZwQq+uOU+NvTNAhUG
6VdI+u1ENJaKafM8EXTNkhCcV972J/tTPqeZorj9QzD/5MJg1+5TjadFYzESmVCNeiPMDtyNwFhs
w3UAQFYlpZzhNPRgdvwz3K/Pow4VttlZqSajW71QEQ9tjxG2BREfIJ0uWhIwoV8LGyT41CUnVPVj
Cbv+nsCVc1xg6pqBZsmyad0X9CTKFp6USpCxxjcVzx3yv0r2UADw85IdcbWifo20a/tzYsr/KBmA
428h72k5wHItdlaqOpMo/17SgRTY9jAGx9Y29Ft9hjhPa/8fv+f5uv6jkQG3aDSabP3O7S6LkRZh
7I5UqJSPyo4/fGSqZXkcOOUHCdlp8nZ+mzcVp2dkzIarM4wBympU1HaTSXDwlFH3n9Z2N3WlCW8U
9g/SvPQqpyAKFCoTmR3b6JOIFmdn+qLG++IaU0ARo0J7yPNsrEAFHqbXIYGredV3Ax8u/ZLvUyAL
vz6Mby8Sah6rmJPoXSkLn8ZX9TLVfiXTrqE9EXMYpe+SWDQaSJihaGxaP5u84lGurQoiiZLWdwgq
JYG3iqgw1b+qTxd4G16nhMCUvI2vVTqiCoSQXWmKmvUglVPHtEKBfs1VZYsm474RU4Z40/fh63dv
00km3RPVd0DjRaoJg6qg3nY4VXMU8qGmxiwGqpGaAUMHLVATzVn/VzAs1JUf8iUg9pDHQsANhwQr
zb6YCcU9rC4mfrKvIcukfgkaEps4HRyoWgMXtIMGbcRizedH2TxijlwbMIAP34yvR+T7/Imxauwm
joZcNReYEf/jgF+QSv899JSkfU+2NJXyKQ+ui57sUYejuzrzqR4tA3/Hyz4yIZI9NQeaYnsPwAti
5N5j7FdR3MoqlKDpoqfBuAQ7iAllB5H2gUu/gZ16n3AP8eXCjTdjPjw0InpPa3YHvRZHgjiMxBL3
XBRVSPeZNmJWeXjDWJJN3UBUDUFvPMeDJGJiZrEHY+v/DJcMJwll3vDzm56mWta+5FeIrbVU6sSG
RG5Vpuyi5+SiNdCKqT1ljsMpfw/jqKal42VQ9zFEyTV0RGjmyyNxfQNQZ0enXzKulE6dHzl0OE4N
KHSA+8oPoVln4qFSyk0bRGdJMHEPpNnHMSyghv7u2SRR0/7HD4ZIGrdK7G0ZAJCxK3a7J7Cu/HK/
rACc9M04Eu+yKtaiNd+W3k3O9gPklwQsv9jLOe1/0Bo0GvCpVc1zbERphFo2MmgpUgPG+FomhZB4
RNgBEQLglFTC25xVUBRSJfKN34lgb7xdziZhyChGZSYeI5YarvMoMWhg5I8dFVAKm62zDRHAlqNG
tioeikkyIgtcq9W4LCP3A1Rg5kyibufrMIZuWTHudT24deieLxmYM++IwTYy20lyp6uNCzQYRZFz
fuprZC0k26l5vxMbq649ucZwDQBwZi9FAvAqMWmfhZFbYeznEfnxEOpRyNsPEhqn8JGDZRy7z/nh
0qThhVuiY+ttuKUlSq4Tg9ddxO3OSYjHYg9lmIOAkJ4cj49zUFj4yRqiTwHIzWByTyDykb4danvW
xDGaS1HmJLo0JULgkqoCMbbiVi6u9Y6yNTD/0rmF5hu+nms1JNoENpAPkuEBO9/0vlA1RRmnmOmQ
rLhhAgFf+qQZPo77SyYfVdibt32UEpz9bL7me+QqYUNrsp3SU/129z760SoI29kozMJqmlkm/2rF
oOGTz/EZnlxc1lLSLzmV/5VopLaopeCfcAM/2vmrpNXPDVaBSf0FjIXV1bzkg0FG/aANXJMwpXWS
qVNcUT82EYmlLd/pUW5Sa9qi4FHTkKpfr0iXPyPxbAf+ofByoC+MjKmTsVbiGnpltJnul3mt15th
78zWEGJsSbSiacNtfkV1/gsWFdYBU0QcI3jBcs2GJLNbpROEXYqkGNY+Z4472YfgB4I2NvfihYfk
L3b3tXabPZUeHtL4FAS13UqbECJlaIOhelBN2hRKsXVKUFvZLR1I0zYqL39fBWYYNpX74tEbK/xi
W0n7pC7338eGnnKwozAsIsEBkaf1cX4jMXmyUt5x10OjYC6rh7ntEjIZizW8BuFuigL9rCTdobHV
sFtx25RStoZ6RYiJ6xpBM8vHWCoHED2dGTE5WeuDmVS1lQ8lJMx8B5ce/LvnKOC5zyCKIpYHbzVC
VvOa71lF9a/j0UtpaUVzG+Y63LxrMDy7YBn3uEQKEuo3c/CcgYwQHUe+fh7J0ZnM7AxTL91eX1wF
ZDqsWhWuZwdA1BYFsXLb4a3Zbj/twAnfQxxG1dqYWl7ht38HzZkUEHh6wEWOJ4x1ZVCY4wnhuz9O
wBUV4JjIyI057dQ/ev3JKishRujHy3T5N6tPL9wEVFyeg7zOzrzYvzqcVxU+bO/ut6MJmZTYl1YM
EPYH0diQeAreFXWAMekY5Eeyg+jXwEfvmO+3Efcrb3iNl+u8f5N9O/f/H++TsnQzMgwuFPu2801O
yyH2R7bAchy2XFDZpzQtRKVsTZpZY4GzMo/yKLUPPRa9vz2M92yeELRTO2CtZLqOsfK0I5JOpLDx
E87N0liesVDJCff8EyI789QSQ5EUvyz6QFj4U4SAOYwCcMpo4fxYoh/zyim0wWi5ymJS4+SVwzHH
DJkfTRWjmynkJ8pwoXyMjnMOFfjcC0t2LsZ5AkS0r5WAnTpG+C45QD32XYEU0pOvh9pr6Vv3c+JW
OOWSNAxtKq0BOszauu317CFWoksz/wjNNpUqzC7lmMBjuxuQPXlXV7QofKtzhMP2IUlMaVZB8EUi
Scqp7+djXnmJE7EJiJCM3F150FoRs/fqqp1kOWYiPHTvWFA66YW2l1UAxbJwbLsnHBi6bxwQHiWW
wzoGhaYcYg5lzeh4HZKeSDcwJbpisNppOZej9yPAwjrdKtGjWVGGKg1CQrkY8/SwMeuXdIAvh2q+
2gxWvjCByNJ2FATWTaAq5cefCy/mFGznmoyf0WHi6O7ky6RWzuEzt1r6LCc10AW10AUYjkfZmfbl
FXISV2eu+evpRpjNjp3mGm5mUGamIPtR9VCaXYF4CugrW4fGh9qEapeQp+egCT+VqBWsf+NS+2Dj
J155PFBNEwJ2KUBFa0cZNa0WMMLlVGDVjbXxOXVkuMld6+GYZlw8ysdMGQpLspRaCD3l3yMV8cwX
kF+xVqDTr1TjfYKogI9/2PMpF9gSaIDpiIUFK7TZq2UT8PtNW6z3DnuV8jkt/y6itbl/aMLLEHv1
bnW3dMZvURrC1fkJ/sIckJH10SzYOea8f/eTyMBMRbEtt759DZsx2cx2riKMana7rXR/LQNRhzg0
xy/AZeBuSZko++6varQFskRkPWBqn+kvm4tyw5ifOaz26wNQEL+upDZVM8fBUEyzF5QdAB0tuiGT
juhiYdtIf7tiO+Bw2MtANBrrP2ZxEaLAS2bN1Rl3yNcIhnRyEaRYlKvJqAtcNaG0HEJghJcmzxmV
IjDja0q2lIhrQpsgR/yJkoJsK0r08gJnR3pVAgLej/Ut9TY8wwtu5BIxdZXk+2AWdY09A1thgwNt
xg8ljdnPiexhktNizfM6eW1sLjZJCf7woaCsYv1dZZdH7M9ycieZUvZLdu/EVN33c5QNiEAdWz9d
3NZorWuAg5I0VxhNdVzPB8Am5nBFB9JhzqfaZBa3yBqluTS5AOps2derghYXcluw55nz+MzOX/cX
M1S+u8cVxdbYeVVu+5KKzBMM7vtpozhLvKPpa3KPvhesvO3HqVVrOjz6Fgn8lvcDYVoOF2wpBBs0
5gAQ+ecJAUGjAEx8ych/TDwAuFq4BQzSoa7a1u5B+qi/6+dV5hJaacr/Li97ztBORgnhJIsHrSA1
jLYC8775g5rYhmxg7G2+LqFBOFGIGRuMRqFiD1urZ8UxMfjgHiXL/AgM4dA3TWj2HZWUhnvL5/UE
dYpL/fR5U4G0y0s/8GhABd5tp8jsBuS1HPDwl9t9ZthwNfxNEj5fG+1FdL93NbkTLhWbgISbJR5k
n3yc1Duyjxb3PsAxkfce/b304+V6RXvP2HTlxilis7H0jvNjhF4CiyQ9zX5QEIgA+SFEMGOC5sLQ
B49hT3KUdrqAYDHXa+I0a/rF+j9WJvdc23ZuSqQTwKLjPMcvojAv13LdbkUj/XcyOK2b7C6EtpLa
A0/YRRV2NpuKrMkfzP5ROECKVW6ZIA8ipX5q5iL3oDXPOWctYbt7t0Y3C5jVkiYSaB2m71pHJ47n
H2e/Mc+L4CsNDJ/w40LmrYrmMlYMUHKVRSRgBepLWmdvh6+65kmOGcvipl10x27xOi15zaIPq/hi
bkwGcp/FABZONgsnTF4N3nEMy8MzIB9D3qX7F/BQChgA3Mk3VeN05rmIl7TigqEuk2ivoNOcyQfl
LxKLk7HEYoGUQ9/XoKFAxTv2Z+XRzrbugHJfIK8tjndfajVXggAj5LNFVYIuUtO7P6J9EpxZuTk3
lq3Dmk8UzqXeeYJJLvMa2KCLhS/8/4lvh1Q1uRT42xyxb4GQFZu133I9JJq+9fe27W2v5wawdrV9
wX9ucBMZF6YliPty/UpogxLSM46LDhYiDTOGB5IvHraeeFYs46JopQzA1tilpmKSd28lWuQaAgkZ
ImCi7UJ/TZfR5QD2cjv3yOM1lD6qfPqRr4L/sMmUgynAUdyLkJpCsZagYHW+JyeWprc+/9HISir1
zqQSnA8lKSBii6OmbHElfRQmEdsH/TslR304nN8Mgb083Uh3SA8LxsW0Ub/wspan0HqSB6ONWs/7
GA4eHFXa0RRm/E7Haw4k1g4221hwhh8bgHsPvWoAvZlcfoRRb4pu2bb2Sfms8j0yV60ovGHEYh3V
UChVvws2Xb621VzcV7eayM429m1rnK3YL7JK6suf0S8FdxpNnFPcZV5SWVvLCU+snMZkY6j+tz9Z
HTnhiF8E0qQ0lyvQmjO/ljpu9fCPY6U/HbgrvTQVHdfbCERR1u60aVwJMreNAxO7FFuyahGTWEHM
4iinAbMre4SIb+RNvum1byv+wxHFY6IY5VZrpunOOOaQUeKhg+ZlBgZ9xqXPqwBoyb1QDdwM6Cfp
HCR95oiqozRVLIZLpzPe3ebAZZFmom0XsygJ4Y9hYUgpv65L5fdrXjcBrCZURr9vW429NBNF47iL
kFcj+ZeO4SaFc25RUFp62/obSa2c5wgPfUViHXFUYwckYoZ1n7jS/KoksiiheVxAXs16J22sYH4d
lYvJ1yPgl0P+IsCcUlNgaNZm2B4Kljn1MooN2AeMi6vDUUUzhMWI3sVHXeBUM1tdWhKlRV6tbCF1
Mp62kMHEZtiu8jCxmk2BbSLTk4ZdR5TjHHOgy4oKEgMcKPW0XowN2jJegRqUsu3GbW5Lm2VP8sPp
NYWwlkCQSsoUXF2qcS7GYyTTe1DgPcP09duzos+p8x5fGUBMyNqijdJEx92P2AE5mQlyJl+o0Qpz
e4Ptl2dCADOkdSUxW3ll6B9hvO7uqLp8OGoLpj2lcrEMkmQsIYmgNxcdVdgFIQhu5A0+Kvcw+iba
I5GSNxZnHgZb4nt7d8PH66n2CpkRw1lB91DSlHlSVtdhX5h0dauDUVJAsHfBizDXZazBhYBa9UuV
ktGCtBu4hVcEmrGe0jveJAu15cd8HRWKaDzDjB1Naf3r+K8gCORmlFcETx39Py/agUcP5bnUldBM
MWIoDk6fnS9ABYRKjdt0FIqcarAcCUGQcS4FuiLw/hH0A25HKt/sWLJhYpCdasU7KRnB21MvxcT0
Ya7VwuXJyDG9OSEyMEHS846Nhgk3t3OUKTE1KINxneyQzEIYNyvHz9pv3f01eenM7lSBYueTFXvj
Ikj2+m0qMyLftSk8yFMsRjNw0QqE+e860njs65v3Gdj8Mfnn2+24H0K8fH8nGi2zoGOFggsJ3aAL
nJY3do67FMum2wSTJbP/m41VD/ut3u92i7O33BRVM2pGRqgCQ49oitrtiPdDMb8irAF8Qcqb70YC
m8hGM/8BN0qzfInJek4OraWGA4SIRX/OcpOls/+2mA9EJ/YhMdL7Xkuoy5qEJKKXsnCIEwJsmP4m
T2Oosdmngk0TxsHjvjLfqtlAq2OE/cYsWMm0SYPq3YLnsTPwSqFOJlREZknkFd2gx5a+DlHi/dWZ
TvivrhbvMGOn1Q5XEQnLX9fc+UQDGPfQECHowAAbVFbAqqN3sFIMtWSTKqVtahJq06UnCaeclf6v
a2XnTwY8LoWcHeb++rlstsy1vOnUf8UYLeFRZNnrPVgamIQpvkUSfSidUBbcdRQMOMJC7o1YKlir
R1yvZcD0hRBiBwRhTJK7Ejp3xSA1R4SwSEOrJVWoeR36XXkpnX4A4dY7pVOYDYpB1ZgdTzrnQTTN
mH/36Abb17Z8Ts4RwUQ0P5EHaA9sTuWMSLO1HKXjjNMMNFIoAgZr2apFO0htdByPD3GbX6UWpTqJ
XMo9kFKWnGtfJ4V6udTma8BjWqod7FBlpLsNnQDbYthWpZhE7e4kf0nYy46qrARj1pZfIqytHXjL
A0f9hDxjkCEJe1VRbQQAXG3Lkz7f6j9J5O4QAMeMb+NU4F/MxQje+IpV+3cT/pL4yRJ1QAMG7m2P
R5k+wRnBbBZX9XMl+UAzje8oTT0oefoLGi+fjJ4KvX9KhVsy3a3uuJXAvfW7omXS+MbzXjIqeLtY
iY9KKwQcnOta7IdkIFK4tpVRfEEsilkUgA/RDizgpQ3fbqedi2WOVxXperSsR+8zICgnR+BxiRh5
eIxoRwhRyxndCanAwCJIruHV9S28ZkN/4yshSoYMeXfrMuYi22oUi7AzR/D+jO8Sa/jVAlelLs2K
GQ9blHCpQT8JBl4JQN6asXeo/xgCoYr9vlVAwwJIlTMSEejoWfHtSMzDPMXBPGnZU3T/1TU/zgoM
hnwskr1eZwn7EUNjIMhy44+0pUZ6IYlHbVTY50f4cu1c/jZ+Mq+5N+G4AW/i7gfoP+EuHKyiU+hQ
XOTJR5HjuESSQvmKnc9IeEinUWnPPhZriCv1oMGWdlZDVJEsrCpqlI0GxiB8fnl96KQVhLLmBKTL
byJUHBniIbC4bsVOd3U/2wAUsSmQlZlFjDxi6g+EiOUZ5ZdiIlnVNVP81POMSMf1deTpdSHJntMl
P04KWfCBI9ljdQGq4cfOxajnxBbSyaaWakKvg1SqlCz2WYwshJgfjiUnHWELrxVsneQJoIJOgIp8
OoGP0r/lLStS3iLrPXiuh4D9u/6MYO8EklyDnRknG9vKVAqg1pszvh6BqTqenRlnAotHL0ivun3K
9hAPYHJZYpc+0Sc3s9DhltiCk7i7tVAHV3HkbjTi5u46I9ffLS0JbdF2aT0zd+05LOWRpx26Oglj
Yro65Wu1rTbpp9qa7dHwRzmiZdbLjEhntMA67os5iJL3PBLEv8+dtNn8vErolh50FD25NoQY7Uc3
CqbBJB0WNc/mHR+lzD9AOKVHv+E3aISxQIQsAcCDM85XowUVrdVa8CRE9oX5pZeVW5lHAasELWfI
+lEy/qdG1xV8njYvN+mMQHgufmjAyKWDTncON/WanPHsrfreCP24MOjxR/Pn9F4K4zA4sRmsDpqW
4fh92nY4ehbrvmJCEGWQH9LVw1i9KgfsaqIR8cpNY/Ts9oB9O76BfMNHEXJlF1plMIcG3+R2mjOh
0vP3ECvLw6SKAqgzIIOc1n/S3g6H4tafdLB901tW1wOVISMGDdjVsRre8aDSDqdBtwrqhQ5OpwkB
zBBVhtj8KJD+WXeP1OqN2hojv/65+Hka5ikCI4EFg/OD+9VASsFP7iovCzegJnB6dW9KMsII5f68
58ItUWFDZy1XR/9ERTgXUKH9BlHgBT4lScDz1uJwFrqTooOTa1KsbWWNo+epGKLLmM1TqzwMkU5B
wZXGCtzZ1d855jKAskfrj/XAaFmQ92hU1Nhw6S4kkfiKQSW8C3zFYIwVYmMnXiJJaFY+PF6gKTFD
HhcLC0ZRzxp5fXKhliwLt8p/P/Fpg2s8Pc4x6eFXGWJ7K8WpcWOdA9pmY6qKPBWNHCFLX++uCrNz
75UNxsnbKyE3ZQyACRJN7b+LK2LF6f2R3rguYlpBBQKLHqnHYp60BUUQGBmBWCF9gvd9YRqwDAcu
X86cBvM2t3Le0g6OfnSOoFIzOnnLvAwg2Dk6eyqnbC3pqsgRmYOq3AmPIdqOzIan2AcmBnm9zkqr
2114hEwSGZIqi/JZQPhAhbWz9sZkbz1vTJMXP0NTo+fNh/zz78IP0/CkmB+qKN5AaPJmKf4ABpmu
lHfJ5rmhwIs4BEKoah+NM1vQwAtO3dtZoVC3/8dmGtDmg9yDf1RTZhgML5dLPR2h3TQ23+QCx0wZ
h80LLzI2r1YBUrP4aXYfQHQpNUz+/6xBaiT0MTwRCHFAacHxbpUE4CGcBQm6P0shbjwDd5JsqEBw
TMBjCvBT3eu2ii3+Fw2Kd0MJcyQkyirNk60ubWLuN9L6uzpEbmrSZrmfmeJGdFEzeiiBVHxjucSG
gjNjT6w652L5ecfFuCcPD3sI9jjCPMDWhCTjwKvc5mbPKQPs+4/w9CSNMm7FldfDb33Vx8IFrkg7
6AJNTdcyHDO7v9uc8HGnp8hB/HAB+3cPIJGvPs4XBdhTyJAJOoBE6+PU0xo4CBmT0/U4Rb3ci7Q8
FT/WpiJq73FOtveboeRbSefw+dp2zqo9wBhDtEWPzvwtAM6Ac2IgVNk/E5kw8KBEAWahW3uG2bOP
LLNbgrI72Bv1+1hF9Yod+gICri0HGVTEwpjVv5VA74lALjuQokyiNdqwXAvjSWscVj/X/aAH4/9W
9G9DwmqqSxJ79AX6xIRtNYKHCo7oKYvhY2hp0V1OVN7LuIABwZ5ux9mHBR/9mKSB43BURzV6A4Pv
/oHJNq0wHC+aLOdVHIpYlENGK6smHEDsraGEg7nIhhu3pHo4nuwL+MKM8Qcn0J7j6GBmTDyoykR/
to8ri22ulJZA+IDn2izq96jbpVSRUkjCbmKDXUh/UJj3a2/VxbC2kPuMDMctadrcUUxuvfKcBj0s
bzwxG6P2AtELOjQ8f69MOXWWMoQgYupz5ztnGa5jLab9yp0NmLqNR+JOqlk2uu9d72zWxonHdkxY
dbKIUjvmUUu3dEU0Gk8FA4Ao8HZVVwODVQzefrHudgj6Q8wG1ezC35URkGmwUoWGMESgErkJjk7p
5JT4y6Wpgae9Y58KZx8GAzRrpbbSrke1XwfwbdustOoqffUcoZ1pJUXgoXQSNrP+ZILwhOa3pfAH
3VynqXc7MjJDl7vADOy0c0PIGxzZKw8d6O1+k3tjoa8FQfKkDh/M33P/AwdHi7NTSKz2Q1uUn0O7
pO8sk+ecDEA2xNgTstuxy8BmeCiGf/MISu5vrMVy7vkoM1Q7gv/HyKHLqSPlyKZGLz6y3dF7HG+t
JsipFXwMBvLoc5/NdO+uWR6ZXIOTQx7S9+SahSFUW8ZIyS7gul3lmPEFsNOpsM8AC+YULUHGAyKL
tsSXvOEGbTW+ktVZPXnq3f0YY49tM/EGUYuLDECFK3WwEYq8jy1sWYzhacU1981dsY6/UuSUfbgf
rbXwYSxb77dzw8XNfsDyPFxEzUBRf1TiQoetCBHTJNI5X8aL9eyzgjXOBwFA2wFyqg92MHINOZUn
oZaE/64MXwerb29xqSW7qI6OBrsZVrSLWda1J1pB4QOSq8gxEQWHLglTvasHWTKGS8nfRoZ6IP3H
DgOcKvbXumBYc2kDiGRScL+va1bhD/qnT4VUQJZDoZX6leTQHxlvA4bnvbZuuloIytKLJ11SgPqU
UNBurocP4Ux1SuSLM2aajXpJPkvBogpEBbooWv0OUwZTSP3Ha6iw9kvNlkhlBUCZ5r/mRPCbiCKn
gSUAzAgzJ2t5q9hsLp4D2bBTRf6aecX0pnX1V6zztphFkql5fanQKxJshKSKogJAVK0QlmgXnAhM
IRQ6klAVqHu4fo+jpm8V2RefKTIRhIvm2HJGLSnoqwLT3+W6jHsD8tnpINYhjyt6X7kq8HrafJZA
6h5MLSmMiMKoE6Xi2QNp/FiHdD91KgO3Mw+V4BYhvu04DZ6yQxfivEFYumdo6AMwd67nULbVgAof
cIZn9hi5iG/esQNu6LsGlPhgiN7PpGRN+BIIYshwB+y1M93i+Awn6hZH1NbcJPVhzlbr/niLgyS7
+NHccvVEmYDIyMoT8a/dMiGxGlTAEnU2u9MuGmXm/fVnpgXt8j0fIx8dXeHX91F99nlY+uT+1lSC
f5D0w5BR4XumDGIBVn4NBJOhZOty89/Z7X0ijxFDfRYIxxUFzjEVNyKS3O79OAod4yfli28h36q0
2djO+thH6BOsVl/KfGEKKx2lvR0EGebxX8CmrRY1R+rgGGQZBaxKyTlpNu4FmrTzEVfHyggjkLRH
N2eWQrdeGf27bybBK5bhcaHGqfIqwO1P4Mm4fvipNWhOzYKAG5BAiG0xOTpGmT1eWwIGuu9pnI39
SOEvVP8+u48rawgYPRl6eO7Al1AesbEYO6FqxLJOYMD/SeINepXlSxd37dODgremVn5Wmorox1T/
S8kDFrgOYg/ppwJ3jgGXZcrOWsXoIm0KeEUoqSs9a87fbAP6PIWKmHJgGFMEHCLvyz8DJdayWIGz
LVoy5e11c1ayaJZrJ9kDIo2RqhBCq0MsAt9HBAC4+xhA0ubh0+G7NYu6OGvac5LZhbjwfW8dd95O
qLKfJF9maUWs00UHqwnIBXr3IDXmutAK/mAvNyMozl7lWAx4QJ6ZpH2ywOik4RrfJHuTERPoO8jy
H3G1KEnk1c03wkH0d/mttyhhB2pKbHgFrb4MuplLEOSRGSG13OKbW2HBUXTCa+Tod71A+p2sp21U
Q28NFuXyId3GvfovP9+OuacG/9Lx0mTNcbbhXvXRXV1UMXcll8kdBSCp3Rmew4kq6S9vOETr9Nr0
Tn/b9nWZh+YpfyoqBFVg6sfumaG355KwPh6lpYnsScOXqPqU31UTq5fYyutOPhwp0oQT7nDlrx3Z
1VMbNh/6aJv3c9pCng5+9mJpSBMMVDnslbLjbTD+6yctI+8Bmb2CpGNQWrL5Hda6mTUpeWk+IlXU
9IM9h8KQuF00c67Q1QPAcRycnIn3vCSJL3smp/1ALZhL/NQepfQBGOEkpQ9xIjbD4HU6HjZ1rDL0
HeXOfzSkEjsFAsZdTRRp+nLl3zpzX+OsAzlNv652RAkPBswvtZzQeeTu9rwCiZpdEUpjRY5ciHOk
PWP2f+Ra4ufLIV1tqwpz7/XWrhnpD62wYIEcUMsrd24LMCULq60q2x/XlgXkdeBwRoqIVmHKA0ta
8fiYq6LkzMIksIsFhOdl7mTJrLU/2U4d/7FiNCYBiwh+fywaYwP/lgcS43EAcRRlaneaCpJo5fTU
O3y2Oke1svB/VnrG5kuifJ+Z7Z/z/E1iYzb2BnDy5u8vNDwPpEEDlyUSf7XftU5ifh27aEQRwiFT
5ECh2L2AjHKAl5MqTh/kptRG7k+gQp5/IwKwStvlqcCNx5z6oCIRxLicoog0VkTPgU6y7ABeToDy
xbMu9FnLENuovZ6qWxn/7k401U6iugk8Y+MdYDWcoHIf14vZ/tAOyYU6D9SZXxU4nj5VbqRDLrFo
DsaKm6j9hU3vXNKivcUmybdBOgCplBLw//avE2Vvvs5f+4erwKmlKJrkUtTvFpfhs0oW6OGeqFIl
YZ+RVeyLMztYBLZeghUjISHNJddiaslAvsU48gFgXM++pG2UIWlhn+Ae5PRK4xc+JdaQ+iDMvgoe
KkSPUYI0HGU/nEGV8PRiPEfIRAy5bSWEdFL56g1cyPr1uflKib3E4qhhtnmW+jXO97A1WnVs1Ibf
kn4yjeQ1OIKobaRKMMHfJHsPkKNPNH/bnxn3Ejv+/UZOf97ShnWY3Hw7SG1+namqjcSE2Q01yr1y
n/DrJ1ftCZ7+b567eAa71rDCbQCKIXr61PxFzoqgYf+A3FUvHE2CQBQLgN1bYhFQPHRzl5flGejO
X3BvwcgSAQtfnf+XhAPNV5gz/+cFMx9jLVF4yjsg9WmWJ85tABk+0c8Wg4tL9uVqpMcR+oGeqAuy
01ZRX4puBLGgiam5bASPQl5BsikwaSy92OGpt7JVq9qvKW1TDMKGdeHt4uZssnyDXiJYLYvQtlQL
Vmp/Bk7uj/dC8hMsGDTVWaEesdgClF7pMci0J9L0sGKd/NEW4EDhFRFhKIJLZDumh7St5GFR/tm+
8vKarZvYlkVVtIw35R0A0bvFirXnvjlZGdCFO5AG1hpa4zocKRtPrgnlzOwajCSaczYriq3HmZOw
AA35Gv7JhkmqT/GhQxoWUunPh9c+XdjqE21FZeWgU8zfv5Emja5P11CgAlayhEg3Zx9qBdoPcLxQ
mBvPBW1nGGfG3vn6qM1l/O4Fvyde6MaJ+5w9Dx14Lr8wAaiRpyw66NAXNh4Mk6WvFL0trfQaXgMt
XvBlNDIV41yQ/93ip0DIdZvK6xvTeOUScdHkwAeEoSOI2naZCtaVAUbRlzHvB+KGLI9kOv/SDP4M
R1CqvdLuXhcq/GdASF8a+rSlRb0HUoBhhl4PoZUztdtE4QnAm2hIBNyzT7IpD8FnyPeoAQB+oTaT
ycRNQkgNQ8wpXx/YPAsrMK6W6J/3M2FTeVBmEAoPWY+x+1NxdZ8fyDrFOn9fLC5pX6tGG3vrQeEf
8HQV262K9YPPgqGHv1yccRS6zWtCSQamlM3/fz9eZ9c7UAF55sUU+mN6ID9HB99r3HOySLDbIfLz
t8xPVaHGt+CY0qPE6y2KRc+/0LQXpfTsdehJHon0omNujffJNhnjQ3WsPgH4Vhixzos23UlDCV7U
58nSlcSTvdwLtJWbqi/5/EKIcVRMdC8imlNBA0X87tyDGJkIJvAsGSmkKAgOnNHdFZgftDpbIknp
gaj9a6qBnxjMd9C9UEg72r0O1talVLD3MvgGThJP7BpeaaI4mhUyQs8s34IYqS04rMlyox4FyKGi
waBImnNy8wDBPJRsMzm+8fPco/qXUUGqFWmXeCEpg/trY5jKkCZ3cZt2pVBZ7nqwbGAtTBCe0FI1
OjZJFxV6AlhLOgNGZLYDSH/YHyZXFDKNGRo6GDn8SNXInTOh3RPD/pwjxfVYw09ODM1bfz37C1jM
F09xftWVWOwsG4KdG9A1JdxWYuLvd69GED6VIRUK95IV/RA6cr4SdXzmHlUxi7Yi3nWklT0NsR49
uJZNN3URWoPCYKm2zhtgUz2W/euOiu5Xm2eAJEkpEijQwxaUFJ+tvkvNPxMi/IibdgR+WiGALbgv
et3HdDeAJ65WAeraeSQOHxCPKUOtBRHp+zY5RmQE7fAfwwbSii/cNj/PhjGcOWi2qXcI0yJCInxq
w3IAt1GeXDdJA5uu2BgBGOdWDH+zCk6cGjVOL6a+7jRvyFFfU4PMDSi0oVrmyUlpstITWvtVXlH+
knPbZzJtc0SQVrAIS6M6FJ29SVF1ZKYHRuGK81pfi7dA/CaoIl9eC/uK+sq0uM/ox88GMtxRjP6W
CbR15c1reyhXIuZiGbWhb+Jg0waK7mEwnz8SG5Yaed1l1us3PmltSVizGns304ngfkJ8EnJw74l/
Kxsgsvoh2uKWZtp+QjSUnr6+cm+mVoC/8tbfcWuxnkdAr+F1ax34O6rQmswbT3Hl3hM9Q4ply/EY
Z8wooCtd4VY6I9GPojYP7pEB4VHv1k1zQZ/jtZpYvRTkGAQst+FNCO+vaHeu50PfGvyuKN+v5PbP
JIF+tIybRZ0fymKFmINuH6YJaaP0HYIPfiaiXJMqa8jwKwi1zR6R6HkSc2thNJEJuXcDAH0keBvt
WBcpDDTwscR3z9/FGs7EEpZVSrB7kTvusPlRgbOwfnuSfFir9mSepNqq18Rr4TsCYDVHehBZ/Ayw
2lFVr6egZpNym7UpJdT5x6tdwqcnB6B4YnLyOxB16EkNN4ohlr/0dIpuITXZoZdTNL8T3Ht+ypqQ
QJLp+TKr2GbuD3eu88DOxrwDW90o54gfr7fGNZtCztFkz4stJiZ93hKDAQBgC+Do6sNm00MgcoZL
UHzWRgjv4saOvUHjGg79abiHVrdzfKiayRz/wGB7VqawZ8b28if3jOTD0D6nNmeP3+wc1fSqIRV2
3+f5+VjTZHuzwWbCS3J61N+dlHHpyMqo5J5SNjzoG/p4Fvj7boVtDAzmR2+eCiP1EEmvBenC9B/G
4lm+LCUW6ToorWYqvHvCOMRde4fHpMOqsOq4wRRaU5td4R1+Y2LQdWKZ0OagCjZtw7W4M3GibfZx
4R5zxTg3nyq5Rl2U08NJwwGaMFWeqSxP8p9BI0Du0+UFL9n+0lY+oGzIl2PdKo7PISmv4TIMqWTZ
/Qa51Bib/StTHhs5uE3WlhtcDm88ayhV9r0poqY1XLLGXVO7r1oj0mwZRaPdumuYohPUAW0dhUsY
Dt3V72QD2YzqNXhCsnBewXlZoPprzEvQnSkYWjl9UcnDYhuzC/0yqzdAriHHOTZHRtc2BWCWinXY
QaECZ84QK4k5I6c2UeanU+MQHgOnSwP2Ic7BtDL1Wu8RamCs+7TdQifOzSaH7fkFLH8f+kYUAqJi
7X464ANhcSyenCeFiFqVt967quA0JNG98Wkp1n4zxH9csx7dvNOtkTfFecTCLmf3xBCnx/h8aoTa
guBfj/xTshIZ67bXXxXIZYC2Dxxi5HFnM+oY/TLBkAT62MNNTDRXMsZDZY/l83aZGogmoQ0befzd
gZC/NY6PrCgSezYEujnLJK1mUdh2aUQn1bqK/KgYhpLeinIWIO2w7RZv32wHFV3rspKhlL0UA4si
Q9fUjzGD+lPJGNVmPHQXOcNRC+0o7iDOhyzadeunb32vM0htr7y1AO7JLsYx4b4TUkHxLYWfP3jz
IE5v9Ppcbbneunbfxn1km3vwzI8Xa3FwTfSNv6nMUmFSc4T77J0V3xQYOHZB4CcDDUypd3GBzu37
R+xdZhedICTuqCxZN5IhCR/miLuZJu5N93TqCeIguPI663TrHvL8kswG+md8+dGHVH4+1pGyPuZH
2K1IRsfSjwB/9BIURmv3p4/R3ruKwaIOQyKbsUt2cPYyFIBhk1sM8ShzS8ysNTRMiDJ/7B3x91Gf
cppmJoSLDIKiLnbLWLtDLNacpiw+VBnNFqdNK9smD/RqPBI/dy2TUg/s8Scb4uODSaX41x//L/a3
jyLw+I/SdpgFW9Qm78IqmZuRJEVPA7cQvmwsCfvHiKB77jjBh62XaR/wdVQazGFA4OAuaS97MICM
JmO9JYSOl5gckOfMxRIO898orxFwFgpBJFMmnezhSKmzhPS1HCLTuJyWP8MQX2whqJ0g+Bc5lCvE
vp37tdDqCwWDGd3lh2DMssqEsGngeK+tfl/ldw+vTY7FQDcrZBDi3nEP5pXQsCjrHmoXfUwqA5ZW
L9QLTfCQ08fvB9vQYgh2s6GaQdy2EubCLGKJfvaTYv+xdiC33L6eEJwqBx1lFGWgc8/ePG7WBkng
kmBLemM/xnIKe266Y0TlniWUly307V+KOyBFjVFnXyfpgEGWQCim9MOolLLpJuC8/PrRctDhf54S
lmx0m+0z0aMrBeTc8XHN9eTLA0QCtsUblFqsq3+NNGvMOi94N0aQgIGR+yHWEdsqt2UMILgrWpHS
fBz5M5MP5I5w+ZixfelsR+3v7MEljxQCcm2ki/C/qvaCzGBo6Xifn8dlRIwRCwvyR9sfDMOAxB3Q
AO8S/DMYoKN+d4LiMXtK0b2pG+ezj6TQT8/pcrf0oVcRjCOJZm5lePIE43M+8G6//tu5tiq0eEhj
GwCdO6/yYAhbm72WTNWXnO6m5Rfm/zhDb58SktDP/5+8Be/L2S/wLCfVchdQmxVRq4TRy5a5Sg3i
GSFG7KxKyM1tHP67ByiKClynYikKSoK51VCWbuS7PL/eNxJdlKosD0Qyq+UQmwaprB9hI6hh15p6
kYr43+/STXgDELxDI+xrarFjBSQPxdyhhZP3alKRjf7vb+NTC0YRy7pm8Qtaf+iSXeF7+XqeLFZD
eqXhTaoNeOQR3kFoAxXFYnGLsJU//JtMfNAaXM5QUMfCOerF351ABsGe/GsKEK3JeBDmzGHtGc8W
j1an+IYv1+E3ljcicjXAlJ+lkv+g+tdNU9yHIDjQf3mh5SwdMqKO2o3BzJ5eTXMuZ9NBYOqWgmuX
yT/JdTrs0F1naxUk1XJu9hviw/eiz8gP4D/XhxDT2HfcCc+zwdW/7rUY0qfirvng06ilsH/Yoh0o
2dpSJpwhbNfcZnerhyjV6CByE3SeB++bRpKUhvAJ+CL4Aeb6cnGLCRpck1X16+2ebIPYrNkwqdMN
+BJAFOecvh1ksfc1qIVa2u+MzCXl12xdLMYHhbPEtO/cFI9k6bSNngOaodq9NEP65SWK/6BOFQEh
XZ6gU16hRTGkQfVTimc955NzAS56SeGPklMxSEjrpMoPUPelmqCJjrGUT2GxQJChouL6ThIim/iD
rqiSvpMV2so2aDdwsqDVVLZ9oYysaUo+l/Gc7/ZAbk4/fqU8B+yYodEbGQ95BR7ZE1cWjIqWdIx8
ybI+fP6iKgOfAfp4dWWsDmav94Hgq84alHYUy30gsfgQzhAZgEP2sVoDv56sTCXylXE90SIiwBiA
l4gRWokbMnMeVPWNpltSSwe42s2a2MnyXtS4L8k1SkGK+GW4NJhabQiMwRkNEmTP9P7pAAHz1tpa
3JhoXEXSRrsHGrfOuEG93mkAgXNR+YfuDVJIv6oDE2AzQuy0jW7Z7euZVgiGeyz6EMu1WSuZv5b6
cFVg+NzeOsqr5XgS+sFQOwfM+nBIkwtEU9I0U2n9mImpyyDhzDuUEP1ROJukJbLJVsPDMuLcbTdx
cecY0Kxkjbz7B4SKBTBpO2SdV7oywgxAtg3/yrGWvOjcEGCoSJIrNXtb41HBXaG56ML/rDY0DWoS
qZ62Kjcnf2Y35+Exgnzq9BQyXsdekBYxwkzPdEX2rlybWfKJA21Y72IH83zEu11EBi+peuXuUK/c
uoHj3QEasQ3pzARXRNKGMvRhzejr9M7rFJxoL/WdC0B59SViGYWld3WM3f9JhFjOuNSHJy5FHsPi
t+JuDrJznQTMxUrqHIPMCqln5MprjDunkqATouehUjR3vB7DT1CT5RNb2Y/fTJu7IJLmayHIlE9M
zoOkW+ZRBBO7xniMoN464yhlDRhLVfIDhhuDb2li03bIB8KjLGdg3gNM8SDCYwSxVaYaU+kW/cJC
m7ZyxZNhQlgwwmqJxGzuFo1z/6tj6dSH2B/rvQf/d6UwnChT2xcSj4xIE0hVXClN1XbiczL1Zkwp
buTP9PuaKvUniOofbU7Q+Q4Ut59LRAe8dSXr15FmbzgyNBNIv3gMrg8/8cf10OrBSdWfRLtOrxHp
0hAVzJTc6CTS+iBpxPdksmIg1dy4paqzq2g74B1Nq9+498+SaPvdvMT3Q0JxGRwpECuZ1BeYPfkp
/2Vfve+uIb1TAWsB4vcM0WyZp5Uvsjih76dmhUVmGvVknZ1S0jQfRz6l6caDvDfFWMPQtDP7YDVv
GAqabxYryV6/5c5UozzKzL1V+xHgwXrZhjXb2ksm4ahlwvPQZk/z90noc2LIHT2yTAFbqEfwwKnf
LPoHGf538/sAsmhRY67YzxmV9oLqxFAfn5sHf1IhzCY+LKdCNymiywYgDEMwBp8TITZtwkTxspXT
foPfLLuZzzeXq68VYg/Qqiq3vW4smMWUV3P936U+7A6BVfHHm8rctBj4qh++eFgMD9+54LxDfB2O
y3r74TmNo0hXpGeXTNLIhkihz259Lzvfo4uf5LKBWWMMEKwVMYvg4L92UKcfUZoZvivLrkxQK33d
wehp6z8zrMOdPkIF9qyDghAHDjmrz72PmkhnJ8OV2HMh9ElqDkUSwqUunqx1GACa9ivB40xpmj8y
3/rncJLGihTs0MeJIOAFazNnNdtTg23fmGRyX0/HyHjXXDBVp7yxBZERDv4HFfVw41r9ze3Ryqpi
yGA9go0tTyLK2fV5QooDI7SmicMb1zbHqWySNcstJ2plgpzO5m7+iv9FZzp5W+l39JL714qG9TfF
2tw+Gv/0N5Arl6S8krG9wnlo/nXLHNkV1tsDZtBmmZ8rcKDIuWfmzgzFljv/qM+hZSuKsDgsQsUJ
k6g+uohRH2q0tbYxXDcHHYvXApqSqxZfw5p1D2H0Zv/6CZ8f515OPG4P3eFUsZd3UDqm5/hTyBxz
KVXE4yYqpcGQiFN2PXY48eZ7RTqdJHvR8XJh1JsD83TmUQ/oHvHQf1moCmx8jLo9n/sqCr+FduAL
+taCN7nh/hdXf1vd+GXAS/gDXbv5jtGWyd1ob8YrXYngvGYf0zdkpthkJnNOeSJliEPcsQFEhG57
6lONcC5iz2gMhF5pgzrj/QFXCSOxdgfbImf1C7M8T1C6DiCNkYLbEyoDUK9V6A7MarIfohD6yaMS
4nvrVcvmc+oUj+YPyRj1JU68wE4305UAtvh5zJw7xApd3ZJiIsSOzGj3LxDLq7CH+oqzrTpaYGye
XmO/VgNp2BmBroAhIEo356BoMctCgw7JSYHnb52SBvIHctPd2aGG2r05/rMkqCYz1do7TeTqS4qS
c479vNRo8tB5oL48w5oad3ArolfU6BtZGYvlEfW0eOhop/FigDPuAPNcFFfepcOET8ScLvVpfa7N
VFCm/rKm/Q0H9Wemrlb2jtlRx09rpNBF8myeYBJ5JuQQhdOuS3JNgIRHXrlL4nBNFo2cI4IJEr56
WcAOoETKfFOucQR6d76AR+gRWR/i5FwgXXHfmG5zc8Yqr4xd7gTu2WpyaQdk9xzPdbz0igOAwi67
ZAaAwyG5oVse+jEnDGoIhRL0FV9n7KvIUzN+bWBJYP2dYpMVlFVYk417glwyucyA5Kg9MGDsO0Ct
1SqoOttZ+YSR/VZfzZlmu7ZCfpSftpcyLpZK5O25qXa/fWP0b4pLX32EiJhKhXzkgV0K57ZgxMcI
Zi69oLL71f0w+x0aYXtggAXOmn2MrmYkYplLoPk02Tx2q4QCQNRxxcif2UiLRlwjItqIUIMa55ID
gjMzjH4tZpcGP9vL1jA+PtP9ldRt8Fdzli90LsI9g7bynly0SPqkDOkfvEA8YF/UbLvSanwbPvGN
3qphYzWkuTBIJ4+KMYwcycwaoggU+a2s7KjblmslYzCIZjkc2Pw4b8IkuPt9cMs7m2GVjZyQ9xSx
oBjmEFJ7PhJIYh6Tfd6rcEjG+cSK0pbKgmhbJSDiqavuN2f57J9+UtqdmRml6wilAdsvRkP4VnPf
axaatgbyV4M7RWhLPw2ZKe3dMy04ak7lMK9OrupRXEA+LMTQ3Wzn9Or1z9iAoECzk94+xTVaSkd8
7hzTydf1Mw1bZi4aGTc2zFw8tWpTFOy2YufGBskDOMMkd1uyelFLndaSNtOIygkOIfHcPm9vW8DY
6IaF/EbGxuVmJLookuQeMGTnMKDpBm3E7S2bofvkGoox4mK1bz3J/t+5J9D48X47KaY3kPGzYw2w
tBd0rQpGRLpE5Umf9vsieq8+UVppBAW2U0Xno3YVbyd1miS4RRgJ5TFd528HY0XfFzF2kgvN5jSy
SkwYHG8hsOs1huVLYVXdY87mUgKG2sN0a6Fn3+9IxqCu8xS/IOcHQ3soS7+QKXdloFqK3S5YpFze
yED4fwL3bs7PPhDAj5CI2wv83LrvnDd7vW+v4fNkby9WgZ35wU5lVy/Ilxzh7pUq9Ob0JUCWMpEM
C2LXogujqaOd7NHOs6yzARgeh5VYtDMEd+95/k37gkrXVmD3+n8TwU1v0l4rWrvUqlKEHmC/2nRu
J9zZHpMYYFo0BEQlbRD+ZCuwUhLMZd0OoDYLcRQ5V7F7Fla8qpqqoIT4cATDwOVwnqEHvpwbFpWX
FMRoh5fYAIgNaNEPo9AVh9AKbH5PqEgv0IKR/LmxuT7UlOZUM3ouDW+Inyrfta0YgzZJQkVTp5QP
tBmq8IsuV9uqcHyqF4LPj41pYa8vjPcTpkCBlF8KMwlbCGoGtV2M4KMQaUb/bWycUJhubth4cqCa
/AWoXOuYlk7JGZpHlKutLPetB7r5Chk5aVqkYjw3E+AVQVJSzmvboG2aOFj1taf89hq1FVjPHvnE
K8ycN5hP6zztl7YLE70HTi7SUiP7xChYGGMktqdSwtyPUyH+nqKfPvdAm90TJV1Zu6XiJyzu+iwq
ErGydvIms9OVeqjn6GsEH9P6OGv/PvkUgD5Sxh3vtMUk5kWP3nbPbe23LDcPc4y90Bx8DmHxsI9T
dqxOKqiY2rk8wXSvuHroZywEtxnx0tCCu8/+SOu5MpZf54OVPZcjNbjLzkns9gXgOZe+4ah20DLW
5SMlyY8Pv4kPeNFX70TAcqzKPWlSJzCR2nTcuyL1rNPsGB82BEpzOjk9yyw3rHL4CBNv30fwACs6
42/tUNUHLu+gJRKb1Dwbgg4vwx5OUUBVQ5f9PQa2XKqfY231FFFEi/plCRriMDbgHL73USvaoSr9
MkRdE3ROLpntYwdl3rhruyP5Qq9r3dUmOHcPdFZQg/TO3saIwmD+OH+pZoBYi2iQ2aUN0R1KHXP+
UtJlOjpAubJuxCgUvX5kqBstkKakvkpVFW/7Li8pTq1nBFRlJqX1M5iSyAL3CBzPG2IJQpGWo5c0
5r9MlQCPYcNvTDQQM9niKW6g3AD4w/RS07le+1HmF/FoRPLgHmKltN4wm8QidOOrg8NJ5Arw4c84
BrEFy94Q0scF6/++QXsyF22C4BKLUPJxZHCfXyMF7WXdkA0FSSLGsmv8xmOpI1L83urJxlBXLH0i
tvg+sbc4awkihGt/keQFdrkgK5J/+Bbm3QJx/NJkF2+P/RDJWD4dbbhJdTJXOGW1zRkpqitBNSR2
cD41BzDxB0I2LqIhQqgmQHZ68ICW85W793HY4Mj0lqdQeSXtOzTxZiekdihFWPfS0I/vskyMlBbN
sw3s/FKBgUjf2ds9n61O43FbRV6w65alIz2PmZkQDirtqy6YO5fSYS4XkSo3tohZruXGKPrM+fP7
BQj5NSvBemuoTrOeDd4lDWYH7u2hN1nGLzq/vmhrjvBdRRrhkROhy9RTl9VXhB2HgdFJW9uFOmRt
x2++tfZ8ApBKRMAH2luRUBwerOxyxOKhm2sNS8aYytJG7V2t+j/ZnrZasfI0/4+l2fbu23p7F7GT
mFPsKvwQLlo1C6k10ICPVQ6vuewgk/b7VHRzg9VPlgH0I0dqxNipxEob4jbnZ4BstuZGFV3f4cBG
1+Hl42lOF5ERss/0v1bD1fdq/hPNOF9Pk8MGX7BfqIiYWVNPG/U8iOq3zGOih0GxILp779uJEQas
QGmP0OAF76E36OCw3JxC5b359YzTCEsrgk76TtcgP1MwoZjc+IKA4vXUwT7/HFHAMDJjjKt37omA
zkKK1BbLRR0eGsRVlQ7DEiUJzHenDpYV0SM89aEzyv5jahxVWk3UnM2p5FssiDqHJ/CMXqXPhtu+
Ntrw/EOYc27CnoprnRSyDNGWvCrwQd3bvYvr9R5y9rSLmvDdQUP8NGtnglZdgxoT/Ker6LEutXSr
t33Z4bISQVm4hHE0C/fvR3EqIO/lCiE9DL6PmGj7RSHRLLZSp5lstCX49eyoqmB+NdTXDv9YA4gF
kAYhTkZEw79+kSWoStAKX4tkEAkj9mmODQHh77EbX+y+sGisp1AwsSBpKiJ+rj86wxklAsl4YtaI
AQdFPFXFXeioSTYt2VkS96ZI6EvHjlvFwrN1ASevKvUOIys21hJ7lI4DoymjxupsvKMJ1aBPbBWP
7rnAUudrjlhVxYqc98gTROTZFO/rTCjlckhrimrZlnM5w6LnrO7YD14/P+3je06ulRMrgFO7wHDz
3vX1ighHtMB7d2FE7XkhVoPRx8Qq/Iae2XVOKHmp6hBHWq4seh/p1ks3X91HPDdeFbUIBE4dam7r
mND1rdu0KXgcKEcazmS8b7OYZ5XZtxnXx/iLDULl+SJqZek0HL5SmfZ8Eq9JtR3zeC1KrYZlqgPN
sdujrU5e/iPln7G9yISBTaetwVIDLfpawZMGWRAlse0tfbcySYj/e46i3jEhPv/NV0fOLZKUO2BY
1iF27AA4K1540s/PigFq4q1OuXkobKbJwSH8rVDmO5LDfP94tpZ5eI1riJ3aDy7nUBxNagARtKbo
w9UT4dzHSt/dFESlD8KEnNxlhrRDS9zX9iiJjo6DUqPo3bye8RLJD1AwRgyyFR3K3VIsBWsH20YT
6JW+w36d25WOTDaZBgw41fuDqzx7VO157d7TkAqBhx8h5lI2xFiBWUpUIzlPxUtGMhdsr3pT8p37
6Wkpg7eBIsPECANg5QX3jTdHCXDzIklox43yxtEbWN0Q8NAImrGetjm3kF3Q2JUhFc0PZz4Y8n3V
rOgpaITU1vwN7WOvLy+E0o4/92ldL8lLKjQ20fvecOZBDXXAxIP7k0k9HrgbKliuNrzX6RYrQIHU
Zq7y4FHmo4KaWQKx39YjUooSPyqtZ6vSShzJCVqujj/9T4bJHS1wBsxD6fUpxSToUfDsXZ4LBoNn
R9cy/gUxTWs8NLFq4MFz0J4KalADannimwK4AwLzASaRLVMm/tjgcEi3YNWIy3etCageukdt0QHP
FfX1owpkopAhLptvWnjSUdLhok/oryKw2z+ETD0rMKbom8fzDNYsv0oDOHQN2BUlDUjXC5hdrU3m
lLIGdTVhPuvH/7HOW6zoWGaLsxQ12ZYImw916p5FP2D84Cn0j3wX1vcqZ3icUdhvXU2cJb29cX19
nAyICefpT5OiAGYCGOl8GDnfFJzD3DDkZuLlR8RdGe8NLtS0gw62gIwuAgcoFbgZ6IFmZYXSuNHC
t5vNkCgisAESl8q7tp4NvXM8PrXSL9vKRahHfQ1YAVSeMo1O/70nu6sJyCzArVFpT6rW/59ECI4q
YBhGPC0oLSxBp2l2lk+PWKqYfvNdgkeN6grnDc5E/rmlzZieu2c933ZIegaG9heBAvF/bwkSoaZ0
VgmZNYoLnF73ibT6QO315MMt3Uuvzxy0yTcwZ2Xf/GYYvd9Irl3K+X+f7+ighUlqmVSIhJaMI920
KO049iMdXXdXcgAqMBrEobWlf7lvd8kapaXbpJwezgCkDN+M+IDUz4XRCGZnGGINQk7wU4kPUebS
kEH9ofZDWRjcYSakykSxbbC1ouqqFtSQPy7yThuQhTUQW94usNLAecM9m1pKf8hvlfTe057RPwKd
67s3L4F6iMD0pki4MwnQ7r0DeuptRKARLyBCaTAM9GQk8w+a9eow2DBvpbWbuCBvDLbKwixeUGVB
NFpCavkuZko5tiqnlJaG4xrfIAdIA22Y9/K65vAh42w16/O1EMiE0RXEN1rdTH7DktsvgCisyDQB
DvrxbAc7j06eKqk8TBHcCKqqeijk2OJIv9uo2VuB4CovAxwQN7yl8+MXyYBDW1EOErovd83+FTzC
zsiasH97+YVpR4+UyywHdXuHV77Xy7t/KN0nDoQ8YgBf3pahAYnjFyMdR6sgPmWGFOhQoMmRnn+O
Fgk4kwJxEjxIbyzu/gI0TX1yfCM+PDQnqlv2CXjkxqbsr7EZU0yTjrRA8eYlcSb+Qqud7MmVeGN7
Ma/XwW+41rVcmOBSXpJcm5iD9nxHWv9oFPsZ2tP8jhEI3tJvaUEdAnXx8qSXcQm8HOln8XQ0sjSY
zQIcz6tPl14w135t+0njCwyzqQ0sfCL6miNty16lpN0O93fsCZe4vBoG+w3RqZ3oIl3CkHBSo1Ri
DeNE3/m/FDOYr6rFA3hHyhAEwtUNtYdbGmXlKaoNloAtSm0mMViFwY0hrPuR1rbjWJFsBa0hbOcr
08hxs2z8nPTJQkh6hDUNNZylf1q4V35ccAnuEXBn7Yiyx77kekQzS5P1qzXwIdkL7xCjK9OHQmdO
1lHBALBk8HBgrsWLKwRy2pLdSaRCDSM6T47iDwSEOm8x54iAuec/Iha1sruqEVj8E51ItePB5+D/
ytNkS/pIMRjx6IitCSx9l79T6n99rEX4y2MULaL8jh7CO+nUrOeds2bjrGNAGwSmpjoIKAWM2zjF
DdgtrGEgEbOW9ng6zG3ScjDl5dOImEG8W79PeU+yF2rNp+zRHGUacKDA5HP4EX8pgi/7UcGF0F4P
Hh9C25pzbi8hkLNJoJpav7XtUWV8KJzUZPwcIXGjBV4FfOsYcrO76RBVbPWY7ZM+SsmYI1OuXboe
v9FMwY1gEOmSgytSTvfv9aUGN+xlsyd8BCsVO5bd/kGNrF1RlXTUaE9qn6RJyxuH+M6QQLPvLujK
N/n6SBeB3XURC7ULLWduV2WyVrHpnEz/1r8GvUwrD2W2QYkup2TILhlxc3g2GqbGoe22DJUEZdgm
3xxSPb5edrSrSf9ZBR78eG3HjNDUowlluNn0Hq1U5xfURkgik7G6U9ywYftgtbUdyJvaMs+IdUFM
5lDE4P3QBDTNj6Mwir59somwRNzKsDSWra3Nmo1mvw7pLCFNrAnsFce1V1VGx7YWG5SZlmkX0Aco
DpNo5QcQ4UyVo3V6jlwwM5BDQgPN8oiZVsejCRINprCi1O5ImfTCbd9n9NQIJtc7UCiC+nG5Bssd
hiqcetWh/XL+TD9RpErKm/ClImry3z3ayjApx2uPohFtz+Tp+KEZz9GLvpm2R1qIbPY65V7Uj/lF
P8OUjTb8l9aVcZKXs0AegtWB5jMdKnhJP43Ut8PcsaSXR1qDbfuDGiLYdMkDQkv9JYBw/YYP5qa4
cO0B0LL4b+H52Es0BqD6iZov9bYSMymPfr04m+95OSDFKH2jA6YwWgEmLNo/HrcEOaHH0Vcp0fvv
vGCVlaGzJ6x1gp9obH8S3UyLr6FRGg9DUUloziftZOsrb4kpcWyhd0OsL0w8IBh11qnIjHmDE/V+
4mjJDE8fbL8YU2cUd/ifThCNBSofpdBiOmt7mDT79KjXbzQ62DGB6oJ6tZVpDQOoN0eQrAykjitP
UoQwQWastVcEWUfv15gHSaevRpeZl0D2sOjEbNAcQHqD2devdDBcnGkqiKKaYPwcKRivEJ+QxxpD
LWcjWujsnNuaw3oyz5gEnoeWdKz4pNovCUPvivmvPZvsH3hys1VfhO3flAtxtAL/8SVZhBvCgFjG
BWv5k7qZxMD+o5l3Hk9LE+n46nKdhlSZ9w4m+1NC5Ghm1Q4fpPqpUcjA4AjHjkdrAttvd5953tWT
NJmVwkgoLg0PpVCqxWxsuqHZJHjl0/BacpIyhtMAegbBp/RGFIGjVF4qbRXKurQYDvBX4NwbGPUk
Qq6msG5VmBL6TttbuMnIy1bMNVS6z5KbzY3icry+b6Yhtpp23DvOSo0x/UhUzXuz1csS2sHlYqcK
hmBP3S8/t8Iko94nNmhe+Fea22M9bJGeiGCNkfaMNthKX5eby4RJJfV5eaxkbQSM6spWDL+m5TWR
9+ZbEV+/nvV4twoqnkrtjFRZ7VXUAQDvHw+zURRSGSFCl501eSe0hPgv7JyIJZXFZYhNk7L16jdq
023zq1tvCeeeDBbHTwciq2WjuZAUgKgH/smjvjH6Xy7u6RuZ9j5WMmHU0qqNoSm0GW9Bruf0a+qU
M7FDpYych651p3beMZu8vHNcA+QaXAHyxN78IG4eOLkn1z34EgWXC1/T+qtFdsyvUeEOdGsWFv9H
lM2xvvfeCeOZ+7k+kiqsj9ZtKS+Jlib11otzbPc0IDTjepvtOfsO5/GCbw9zmERKHvrrlMVL7hMP
MpXoaDKbjphKburjhMlsFdPPEvPquVdnDkv5v57vXctGZL0w/zxxSUVolPFs8jJSNSv60pPe3a+z
5yO95b1uFM5ow5YrVAjIvIBhjJr17K3bNwtynU+0VbMac32BBza9VhSBuu5rFMp38fCtCTMorfHf
2SrgJlQuoaqXPv+UIsbqc8qLZRyGynZNhidOF2/Nr/66lTnQCEMeIk1iOBAFs1pCNBCr9xQngvn5
ld+uuKvMcFhS0Pf4X7TDbvii2bTl/YJJ6zh2hHJmrnS7BZczyl6/i7FWdGDPa6VNz1DnAwSL24Ty
aHTopjG8IrCex1OfBV+i2yTVNynAaxiSR7/cagLXASvbgzX3XAtYMlh3/wS7CvDzS3bc4pF+soDd
s5VkLofLvd+ToJbUBK9LPUhmop6QgJF1TpV3CqJ4xQXoK1j8wdzOHuXj3/+qhFgwqDZECJEUAJ+d
M1oeSSoVe9oCQPR/rMxOog5p8jybZpYYebwzs+hsok6LN0tQpdsQTsSrg+Frhy9PFOgRh0bKd/eT
wVMB1OmtP/5t2ymEGV5Xf2u/lWH6M0RmQFWjFfvVcB6TWrSiSK3rnW7GVTMKkdsWN34xQvxrP5Z3
CB79Zt5bBObd/P0vgAWM7kYsdCJIh4b+XBuWeiY9KbQZlqln39efi6rKK3kgbdTf7SpEMG40V887
SPOHUmrWEVCYow08ipHG8GY4D2XUk/MJPww3pdKsXOFolzuwQp0ffCpzqo0+8wPkk2QevhUOAPMt
NcL7DBHAz1+EazbDtFsP9mVk/zgBqMY5CksOPCwRbghk5FPWx/Zi/RN62r1DpxJd+OHYr8XDD0YB
0KBx27Xap6v8C+jgMMnoCGLkYpeE0v/ajoys+tghjs2ZNcGLmyanK8+kSeKwWAfnHUE47+3wMDNO
2n+2MeEO72uIORHeXVdjRaToQ+/HeODRkMSCL9HX3utErnjYlucqY7ZZfU5opaqmSIutD7e8zgi6
VGrLQy53AkdXvLJ6xh989UzDlM9No66wsxv8jHKxlk82ue6B16lseyFvRDGRLAY/0BvRzMSC0t7o
29qC26Vt0STEznprUuz+5MZV2fiDK7maw3s5KjtzVmchlxOJGDqivr34KEdltuO0kkIjH7B2w/v8
dgE+nuRn0l2JfMelZOvbxQX0nNYsxV0Lq96yAEVcgkKqPmqEw7yKvmZb1jIDMzkqm/sOo817TOIq
5uOWSWBolwXTe7b2cUHoZ0zmRZDTSTuXnGerItz3NlQ9QQiAEzcGv3feAhiOBsfPXPOBzlBf3XGi
M88PeNZb323bqJU/Ap4scDOotHG17CkAS6ayFlojSiffCDg4D+q74mt221Cp2QLRQPsOzdL5pfmT
9HGgqBsHS8j/ipk4d2TWBBOq8ZyvTySbyCcYWeuu8oMGADrVKLlUtTqb6XmTpK7g8x1mz5C5SI3n
ZhafzMPZPn3V/eH0eGkvibyCUMdsSIXSnOSYQahWeKXOkDcGRNCx9InK06nxQYW/B50DEj+XQV5V
xHV3TAJEOu2PwWCtYq50CbhWoMxpl3c/S1i+hGTqkdJ6Xm4nlSxEqGZhRI1VbL8cSJQ15tgIZgjd
l4FX+U9a6EwdLnTzKMDz4SvrJBtbP5AoGUigCVZ+Tw+Wa45e6nMMWnQfPbFEDforYptsvVSmdrd7
Lp4BTZfkkOgQFulZi+wBKHsYCfBb0hngaSMszzRI5N3N3RyycgA+BzUh693WrkdKw4hOGWWP6pNh
fTm3fkAMBkKARdO9t/38ryKLpaqxnzWwkKaRTNVtHJZtocB4ghFwnfXNzIvUrqfzWzGJpXDir7uc
tW59zdW5EpqzfKv56OtOpWxMrjLWANAEBkcWPz0TqrbKG57XmWdTXd8zmvlFuZj7H/MXP6czWl/8
ExKv9cH5i7LK6IhWXHGh65bDUfeKRYxMR6JtmeXNEGoNRjiFt6xKJIV2Hw//O5l0d3uCiekfoL2k
o+HabYVl0jhlJ4qy+iwevqlIYUVZR1XJKyt6eJCEjy5g3rWrxdYWWfVvEXgfYpOQP4YuNdP5Sqzo
JPQ6zjKjp7jBJG8TFVhNRFq4/5kdLJLtvDVOSZLW5jkeCPbgcscQck0ikKV1AA1jSlMMRGkqQ5ik
EX5zl0lGSgjuLD0k8VmJThZz74ZdY/OJNR2TtFlM+GLhvPzXhDjtIJ14SrYIhl8KAuu39GgWbpDk
yqpaKH9Eiif2ylWoWhgdT8jqEWWmVO87p2jPNtx9KB7UWbPVfdbFoBSkXQfcFFQ6qYUozlP8fj+V
xs/BmFU5/4vNRoMjbpS45q87b3rwDMwnn+KNg1tblRanuWDI+l/u0+78UV7ryjPWI+QcZoa/bWDe
YkOfC+Tyxw9Cz9xr1WWFpmHqVLe/uaBJhgygG8NYNeqoZmaR/76GF+gnf0hEY8FknoA01Qyr56by
ITOUxlKbGKhEtiEZjFagHj3qsmugHS8jm2wQ8dGKbk6g80ospkAZE+dZQoXOfA4zB6oyefjTC0As
2qa0KCkYVSW7DXj+saICLZ3SJRzWI7atJ+0skmBSk2jM0eV4fOMzi10kQduMGrzfIyIZKyWYIplJ
3JFdVkx3Hc0WqzeNHHplPXAT82N8FeyA5d36hayh1JVdEtIOjSLOIWIfcCqSyBzibCfeZWR/f28d
8MUKaEtx8QYvYa6O7mparuhVqH0aZBR3WSKGBxJQCGoQ6iSgFEL/5TLpfhXlzSoVmblu4zvZ9CZT
xCbyv+Vz78jHsjEYN+JxO4RXPFO2odSISr31WqSxK1cA6yQmAV8Pc/d/OD0rfd7U5Kqj+A9gFHJT
GgtulZJiYNXUJdWN/7FUbYXhQVsqqsI8JXzZa6uUgnk064myq441FXNFsneWGi7jXwGjPUwI/bNM
W+crBANMYTqjETLko7ilFtu83LpeL/AeLOVFDbNzH6KlvcKJRyfGtaUfl2a2ssd9u10VczwbFnpt
a7R5rq7hm/HSILVxTNAGCrn0KH+8bhntlBaqGBlpSu+0oYpLx4VMnhd0eUp0EZ6/3RXnpAjgE0Ks
e2FREYp2QksGLnkFyeIncqIshMQxIIaMiy7E8oXWjZcrZ8fTKI+CQeFC11UId0DDX7t9A7C1f263
jxMjnbnIFgpqo0qxdNC3sDqVZjb8W7KmYA00JANVeNDABMpNJsLiw3Sjuu/PtKe2AsSGkkEkQHgi
oM8hWkEh0PwBbSC6L5gKm4P1dTdWxq9ayXzq0Ff0LxGnSUxSZ5GGtrulOyexNYex4e6n3y0Bi5+5
qKP2421DXsY5WGu7FTGJmWXoSiFfBNpZJp/KEPMA7Wj7q0K3U50zBWc5EN/nbyGtqiVvWHP7G+sj
U2xBnTcoR8o2KcOlcb0z2DYx9e1izTxqP3SzzCbNKZzbR2rjG+Uynn/BxF0OTgIZAppRZ63aFSoy
+3/noCSO/qNP6bYOzEevXolmjeCE6+m2Zzol0R8xA4SsvQm/KQS3aM3bjciFldKpDIYr70K1iuKP
kdzhxQfXspnVU/zl8Zu8XpCRRM51Ai1fCe60In+Kav8bFnUcAQdHLcjiQMPITaweF8mial38/bUp
PYP+x9ddZxA/jEoZLqqoL+MYhqj2FvQDzdLJxDoUmPNGdta/jBcKGS8XduFXIZNQa4TErvfEOhhB
iHMfZ+oLtMkPqnOlvcT93g7tXB8nonZR9L2SIpI8WKDb+D1xqouQJAhRUFOqppnrmL6TF5ovQD/Q
6vFQAZcIM4GuXY4iMFNIUqCd1Xl7XY7aVR444AVolWFWM2gqaBicBud0+yy2sACSIa3qpujlH9vV
swDbdMk0ceFUTsK8NX7t6xpP7gdrWuPeGMIU5nfj0zahKSkk2vXYOPNNABpkjPgVbbi8tS7mToZg
uXvj9p3j5WeqESOBZFSQkpVkttzmy9wdzlUdKej6I+D+Hnd+t6M6RV73padu1Z2UGzDI+e9we+or
ak5KyO20tG45aiR4GivL7Z0E6xnx8Am0XwtnbEkL/pqAzNyjSU8GCf2antzmDMZWZmEJg3e+CXfe
0obUYtKWHNP3oQ7sNMUED0P2jCMGDlsGrS8oRLBk7ZXOGpRrn5oU+ao0vaMJGXR2tqgZwNSUM0bJ
GNxLH1hV06V4jQ8lTrrWgmMKbAlXm9oeTMwM3J07hZAgx98uRQvZUlf5G6ZRZIJxH+mYgjJDPvjj
FhuA36Im7uj4JBI4d9U2JB73DGjJuXNZmnI+HA44KK46IGGMzZ2bUE8zV9hDIBRy1uVKfhbSLlPR
IJe4acm7gm5UX+PcoSoCA//VlunbXINdcwVLucKy4O7IzdG0NaYC130YGJvE/G6MNNhWSWQKMTF4
xGuZ3h4QuDUx+YUADtafx7WuwladOlAIjh2PDRzRRA7cbxtAH1FBBtC0AdXIOosVi3Mko1zDW4Q6
KlEDqLv72HnBIOfZc1IF4cvDOcXgwMu6TJNym7Vq+E0pc8ORXoB/3LFbk60CbKtB15iChDLZbM7F
Uf0zWhwXm+N8H2h2FZbqYKZze7KzhYOqgQE44SY0PtjY5PBZpuobN7jHYsmdU2/PK/cfAf+3QsOC
GYQibqvi1NnhOk1m3d5udh4LX3jAkIoJUM0KeOdgcfIdqwVuaOim+pNFEl31fGZHJFyEMlNy1jPW
ySVuBFgwEv8CQDgPeA/Hre9C+ollV/eDdcLTJNL6em38B92eMe9XNXflGY1FZeO+cEpSryBsSIgl
pO6D/U/kaidtDV7pqJhj9X/OMrrCzCUletf5YdW0vxI8JZj1gD2im6Ws+3jfwcDOAsfqtX8RIGLz
fq9/k6D4pysMGWHGeJPR6c5BAnNsb8RxvcbL/ys+HrQjTM3Y68mXzLY73vOOr6+pt9ltbLeqcMyY
YBdoUHR+vSAitiSGylT/u5flPfEwrP19YIJefm2ce+buOFsuWPPtS/EhhCIzYm+r/w9Kfg028DnU
RWhClZl3Cdt9Ym0psvXbTFZ+R9tos1PKm53+XPpDK4CNxTE2IhdlpxSjlPclKlNDUa1n3vWa3pYL
xCHmy7iHuzKxRWFG9jHhF6+uqPwAcHbHNsw1xJDS0QepI/I3viVDW/eZAzz+ur+3zLAzl4/yQuLU
dlQTU/l7+7V9E+JlC/WutSO7i+hARu1Yo0E6m2a+HBV9BKryk3UhYCb/QPCyk6S0gEkufo7MuTQS
Hi6StlWwuUX/PEK4+RjjIZO1cZrLZLxQ0Y1VZ6Ah91T3lfmn1UxmSwTgADjZ1OOc2K7nJOn6yAsg
pYfRfKwCqmTvCOg2E9uOLYtPfzqicWFJJlP6lr/9AhHV9E2cWAP8PhVDiS4Ho64Z0WtfPbARt5VW
9s5wJALOF3OQN5JqGPeOI2cVdkcNwmYXXVjVk19Fv5dFhxlJKmzBtX1MXDRdcgTMsyGXBQqeItQ1
Dtp9gCUoXsTK7FKyB/BdWJtrACtSgEm9dw/COOWRlzugBALzsXOSGpnQuAyvo2gi+JQnnUQJUMlK
4zUigFHJsfDFNY8cu/UYb9fEy8f+Tosa0NHARf7QV2/ozB5JMOX9uQuLLzHkm7R8SgVySUxfQxhU
KD4uVyPXWn6wWsaJZGeh4T51aGNpp7mvLwYk56lOxX5oC6DplElj9+4x4hVNfHyjcV5RhSrwhRQd
jvXsouKjRGMPvkQY4IyZzhnie+lUKQX8etBN5WPrHJEOulVppCb9Rjnwr+gjcWSj2miTMe/wzpvi
6xc4KSs7SSnqhlw+yXXjSGxijwdfmc08bJyvOlGwhHDZP8OEh7asapi/Tb+Cku715YMSGkPyD6go
/x8iSD4X18eINf6mbWjPGdonDQLEg2gT4ZbYP/cH1zyXOTB7J+HC2c57Ix+AeRHPn3rxT2IADVi+
5EkmCHgQW8iuw4dcf6dwutVVHwqt8xq5FLaS8MbdmHBvU0HezST8C8/CetHLdcc+NBhsBcqI2Whe
4XylQv4QqN0nsJYyqjxeagaVNvzrKml0favoB9BXo1SD5SI+kH7YvwM3FVeX7nx0iRDKJtwfdbi8
iygrDzS6b1T+/WpSbR/Ow99wqb9qERywYTSzrVtMHD3aegyJjU2jEJVzXVIOG/HLnK9+3PB5nS44
fJhBw5W7fiFd+dAB+yQWWXljIMyIXNRX65idxM7L0k8JjXCzdZcbxAagwAtdtC2b+6oZrXuLyMyR
Q9h6bdYrUCqz5zwEE0SPiBbywTUNiz17ArU6eZ1x4Rie3pcD3z17Br81aQbFiUx4wd3vfErXQmi4
gRJAMiqaLqXFzKGVocKHTmfN27qtd+IC5BrT8pCqDjo8N9GeLP8QwEoz8vq7t7SEUZiD8ig69svZ
mMMxN1nNNlF8TxRdZwa0OTe4IfgKiAZErHqxD3whyLTYw4pBUEzQfovQr2ZXqKdMQ/0LD8kQXSBZ
FaH8sDtlCoLOfaPZ3UPARhs6dCcB90Gek6WoqBvUGgmYsr6LBYSYe9hKWYBs1u2Lh65sWB7F3Ww3
o7ZKYQkdLwk6aWgPNOHIwgKNUmHSQDKhymzcFMZ2bXseyuXfMSnHJSIDs6WZbub91rQjOjau8j9A
TQGSPhEwIcbf9RIagMSZJk1w8HLaLWX6aJpnSt0JXybUCesFSQVcpP5sntgW0pYyEeWM/aKc/95r
YB7J1Vi4KP6l2Lv1uzw5LIB+EoDhDILewStyPMXw3QU6DUjMIYF+HZPUBaY5BLxVUVKDkMZAh87e
7gNJSKreZjAXkNodAfHbkL4S3VLdV8JFlsJ2uGaAWbaLS4TpRhUPn/kFLV5KyLwjl5hOman26r9u
gtkWJTWRRer/IP/WoA3q8A7GXuopgHqNPIhnICblucbzRztz8RaX11yywyr+vR54SCgiYccdOG9n
xus5gPhneTl0GwTfIZ2c87jVqo3RjjD38PcSl9Eu+ndX7w9l36b7u+/AqFfJbtS1bZb4enRwKQ52
WYAjR6fb9WZcSdLtEvGjIbzOt2q92LBexoT5hRLSdknj2ymEUeKxAulE6+R7SQV470TWZHTZBVrC
OuKmQmDXkSuQSVRNIIxomSbVP+f0G6L+gBK2i9gy50/1hryMz3Ouj+QYRD0SSOrT6dt0b15782Sn
Pj+Zdk66SQDuMFX08vIk8nk29sdEIgmffstqqMhpoqFtjhOO7Nyx6p0q3yllk/W6ZTMWxc87uq3v
moBVONaygexK6b3bLNavvKi0QuCT75MHmfTI+t1ItMdk6iqBn1IN04aDUou8mhgoOc1+eplhQEkk
IJcCQFu7E4TMtYiVNvInQg2GMtSN77ciXELM2CyyXF334iTTfwQmibDT6FsqfAWq4gYd+9b6sWwl
UfcejM55zX0OES2KL0DXtC6R9k2KOVEEh4yFKI58bw8xBKZneMGums6e27Jkuju22YEiUvmxO+IJ
vkddDY7THBpVGvsh/3yFQrGTez9hyoX+ciGDD80jgwTbOJ/mnDpqdUJcvJ3cjx4kkyw6gVgoBwfW
kwh2R9kW2eRrE+kS25p7Fn4sizNa5X5ksSv3HBrdmnrL3SvNmXmsnjgknOLSw6s8+U7kPT6sUUxX
oV9tVSWVt+aRbtolrRcKiDnYAvPSAlFbieraOlZaA13u3bNKgJt3NRUKUh1Of1p19GXy+G2obJHY
NTOI+hIir6L8QxJSLfUIGlkqk1f3kb1LmsUzl8XO6+gdIx5XWbxtjNPHFfyyo7MKwKqc0vD1x7cJ
EudRSu9oRTLjAO6pXyNNPTLSxSvZZgIsHnnWx7zJaTIlWKFEUBJ76QPuqL2B4Llc7kJYz4vCAbBs
fGc5lTkx+9NQVmsZgSQIYYAsqSaqV59tgj33dEZbZtT6tv1hRB4hXiWu1jrDKXEoRUwGTHRKSOyI
UUkKAvZjFUlBoF0nUh3CK/lYCGw2x8VFF7W/BtG56GFqp1zZkvXywLdZ2OHgwuYFAwCHLn0qhTmc
ojK5PwQf9GmhIz+5Id2tfK9l0xLF/QWCIklIxl/wh+wGxGTCdhfCeB1HI8LwgxrC7abdU4p6GQgU
V9cobqat8LOAyqsOfopsGmVfrmjyVJEx8cNPE5G4AY0WNlTyGtiKcQFtfvoh/G0aG+lT11Hv4AJ1
mlTsvNqvshAJBwA3MKr3YB/OB2/fMFT9HvHi5PVDTG7TYuS6H92qHWc3S80nMppYGTgiUDXBLG3k
fPED4ZugrU/pGfqSYSt8BU3hrSM+9adE+Gzg+tBI1WYftFwpd4nv5YwC8FVnPIJdSOh1vV4sbn3P
SWUAs0lfbRsu405hVbk7eeS0uMq4F7EEauS5gUgSuIi7+X0SjdhkXdOrghrjR92Ze04dSwtksnhD
HR6CJsvIrO7TL2B39gmd4tSTtMtladTnGRo8DN/Z+MyuHpRm/AQcxLZSiJ6zjvrFeVEwgt5QrRY0
R4Hf6RBXbk8OOvXBSlwY/4dMflvAtoD+2QbNljs67JWuuR5IV5X3VfDedhUaz2eXtRHuWXkMMk+o
98V/o+uDHswh7WA5+AH3H+y0mlO1s/Bq0X/WhaPwf8E8PmZmyzDpbZyUV+pwoLEoapQEE0cbxaQK
OWvN17y83vjZcfQ78Hk/Bwa0EABtZuEeGiAKfh1iMWeI5LThefajrXeRDsAHt4zv9iCQNJKa5VPT
0dEvqjQxeRDdOou633HO/4kCt1oyfkX4zOfuguIOVa9iCMLut8wQacc+g8PBS2loH89azcXpnQZz
Gwdm3IG+4jhWdUmeEcUR7o1ODvaA8GdsY7NRIhTkus70eWSK736u21SBtbToMZxqcU8eMsc3CFJi
IZkawxv0WojSbKaLgIThoPKgfU+Z2fNzRxa18pSlS9LI2X8ghEGQ6F4uLnSyBvZYFVDOEzmZPEge
6tQwuPeWxWV7cVLtHDqWfNDL9iz9qv6Rz1UmGIRA2zmRsc0WKxnoc0fVXPcJG86IyAGKgf2tUsub
JyitmR3SQWoPGyB74AeOGYz3OR87u/j2bYa6bt7i8X1EqAthF/rH0PRtL37MX7jakVhZW9ds8R1p
RyFMD1OOP4PGyTgFJgeG4kUkK2ngDc/j5nealqOFNytvSvypLWDT+PX4Jh2fauY/X5ApjAiN2XNn
1GFZq++WDpfq1WXP//AewfWPRPWuhH6KZkOH0LdbPN/pZ1Su8s1zS2KOJr+v+7QnBFS3H3IBoMGK
LhuIUO0pqohSMLhkewuJu1GDLAhWNSJrwgGpBeIZHEYaZGmPkpGwerO+Jv74aGBLkMbyedcFqSkN
9N+4kDse3Cr+xuvFlrqXzYtrrPUEjyZApqMQkTRyRLTNbmUpmGjSXGz/DwH0snHPRKp2F63Qk2pB
oDlEqxjTidzVVshvQWXyvlgBi1+zaVe6rnHluIwcvcbZd4CLKldC31R8vY/C8/h+uOmX0XlhNkDt
tL4SvwXXDMRktr1uUfm9R6rZJlU3uPGlReAoCAOGSi8ebG4HVr5y44mlxy2hkbnAxcKKewxTup+X
IXNVVyPCoUrMqhmb4E0z90bthcX+kpJZGKwHlUyicb/+V47vTfW7PU822K6Q0ZfebUAiWggA6wUA
B8jhb+Ccpj6VKSKoQ919DiPDsam/xbmfBDo+QfwXdNxrvE3UE8qU5wXm8T5QGhjXHFRIYSt28h4Z
mDCbaPc9vI9bXUSRX4keSrDaX1O8NiS0qNx2yBU+IpcgPp2efpVBE7oJLD91/yweS6UPakHHrpny
I4O/w0QtSAs9Oy4wXUc2FWCNTPBX0wwx6AYtAj/1SGqFwXSdRbFYTcnUbrnd8rWajomxTjrbVY3L
d7oxKhqGca0HGHhn9SqO/bU8ff8Zn+wezsoji7GTV0M/91mAtsbPPHeVhsAxUiaxKS+IF/oo9RBG
9gNWgDY8zPX63nGTjH/FOf/zQwT0DouM1ee1NHuyVxz7qeDBIaRsHVeVPDwyjzfdnsi0dmZ7FeXd
ugSfWdhnuq+biNxQHkv/JZ58FqlnuAenPfqIIoTwrqKs/c8XpapqF2q8tsIdmTkNZpd7dNPnDEvv
JQfzrBuISFcCuFQ4wNMD30Y7/qQJfzv2/6mkN/1Q60uTqKecVa+4IjL1YCdtImDuFm0HqHgb57AZ
cIpdjwO1lv8c7Huju1npM12r6TxIiOaUwQt5VFpkyq97yWnKXBDdia3sZf2qn9xK87GCxJdrnN+h
EuOMzX7FpXbt0PnqK5N6wLQho7oRNdWAcIzfhl/RNauUlYcR0nuYWjQ5mznjLMjMQbGLL7Ue3d92
VFPT1dTEt9OxrSR+YZYxJhRBpSp6QG2WUTK0qxQDw9pnMXjz4UVN6eLRqPOt15kE1Or6MEUIyPY3
iPp7AJbnomtEQgQ1gJCPNf81ZtFz9ci2NwXULN9lnOiU8SxT+v0S2qyrR1xE+H0Tj8o2qzlRVgY2
R9XgKxMSWHULKbY4+d+Va4s9JImCCqDssumUUFHxKRt1V7q5CugMf1nC6qecykghOJaZMSfGsBRv
/bp8CtXBpcA+iOJzFk5YXVX2tlmj8G8VyHDyN4dSDZtPjP7uoN/Q7DuC4nCXjKPZxfMH8bH277kj
H97aA96LdcTAUoTlocsKpVCjIodfqIn06FFCKyL6daMBCa/3LruNY/RvzT+LCQsn5jpUC4j4CO9s
7Hn7msEYJstzvWY3CHEPuPp08//a2QuNwsYTgvNdrN+5xkh5xutGSSN0FZgNumcl8wSiWDs2UQjX
XBuxEijKRBvoD6/Mkyr8bRsN5l6+vilmNqix2EyKoImOspo1uHllhRFYJ6xvywG7uKebs6XHBjBe
sdntQkJ5dAAjKGaJF1R1tkANnzVY7XnbQsGn/WAVoghcVDMbhy+Ja3hIii2fnWbJuvW+ImmofbQ6
SefdPYMKPgUn6jWScLHIqaHmSy5Fn9JsMmE50MCu1W0UUJXip5Oiip+kBQJOV7TiwQ1vDDheGBi/
PG3b7/xIRJNTnEUhp/s1Q+GHqX6pjbFD9MTJfUgB2oMotF6fYRKVJbZZVqajMksyevMxfdQ01m+1
U2uTWL7tyT8bYlAWb9z1ECOIGB2Xr7mA1HUWUZnvPDWb9rhOWdFtkNsu0WuJGdeiL00lecYlASdB
TIOrcaKhiocsXaVggddAJtcF64mWht2VLwM/+IvhWfBqK+9aeAynLOdZqWsO+4j60VO7Phv9KnAd
M46qLzm6yXJvCS/DYaJOqGMXjSV7B1rFIs+/WK+8ovyZK6B4rNpJ7jOSQfO/VjexXED+U1v8bHen
ZDUmun6zWCK6kTbyGDXF+KXDevuI57Y98FTJ4NcEgDmMStie+5ivKFsdUzqAeegL12hOYMh7T5j7
9NuEmd9wTCsb9TF94pBhpjSMqJ1Jfgx9wDFbXeSen+O5gyLMRa0x8pFnbwWBWfSSXX0evoo3SdqR
aU+Y3DaGokIx9VlKCuR7nrh1DXF6KSC+JXtbPjaDodNEJzu7R7GVBWf3s4P+TvpBQlRtswbya1Kz
eEZcL/ISZl3R3d2bv0TjFWehmb+besOFf0MuJ/aE3bxPNaJV26QopUehbJI49lpmyRCKvzdlf7Zn
msHNUCHwfUyFJ2QdzHIRkXM1LYe9G8BdZ7u2/lI8RzUJjVoDG9dBQiw9eYwNVsjtFdLFZUZweQES
eLMK/dy5jimtVI4muSuUA7RirBb0TMhBPMB9/y6mJXI/n0oL3B9ZsMu+9XUZnlruldFYVCzZ5NPi
qp0Km1ICWSijnDXjeg/Q3v+914ZeRHQk1V3DKqGyi1Hb2CJTh1ASeUSXIR815uZxWRNJLLLtVZsE
dXKIvoJoFDTJEzrRsfXLLo4wAMa27pWPAOyxUd0q8neXWe/39T8jUqmrK3PzXjNV47NC8+Wi8w30
rAPGqm5rypNAafNXUzzcl0rwy00SKiFO50oWzoLgHO/Db4rn5sUXvbzfBVIectiyqsbIg3viADZr
+uy9YC+uzeRBSeqJf0IZtW577OAJtwI+KZoK5oSB7E2eu+MIilzJ0iw2LeM/ntNaZMHKIkxnJ6OJ
HU/u2CH32UeAe9Rj/jGnTnBFbjS4lc8ApM5Gp4b+kQKeDyQZpa/CYLOi9oxw8cf/dvv0+p8DilSE
dviE6bBSQaaIp/qRr0ewZxhDP54q/xjkG6DGefmnB4qdrxUj5wd5SJRmG7XXB0qyt+0Ol+HQlrWH
UltN4DQ+xAs3wZCH+EEWSbJAkqC7uPz+rLFKDTiOIGq6ToQjFUTcjGy+L8nfas3mMP1SF11AbZ/8
ZidWY5btw/0Un5np74bhPX7l8c6G6gM9AQCWZugJ6Z1wn0mPyo90j1yoFzM32aD5pXlslIWo/D3V
5mqzdMVVzwlHJHtDFf5KLLLsoK9jkQwuC582toCRGSuYbP9Z1EZfxJHKQrt7vwv171i8gZETTlML
vioipDckIvSXkT4fca0EKe8KkWY3OU9HlNSTIigDcYcglCx+qFYZAQ6jiyeZQAI1qjBYyJO+GlZn
8AqEmpy12DT5y9nUXitRiZhnANyOI7pab9qrPPSRu8wEDEPWCP428xcE/dqM1oaVuloEh1qWJkM9
IckFt8SM2NZnmIbUXcPvSU8LueQ3UK18iBoSp9gYMnGpBwx5IXPRkBwmJNyIjgR+x0rdrjZ2z212
PzHOqo0Oglbl2eSfyFwlGM14bMYTY8Io9EyFLCMj47C3vXuXqsobhiVcNq26s6kZhUuBGZOZ30Xa
CQYLf5MNmQCLgVwwrin0fZ6IzEF6fKGK4TC1t3VsOF0bmKeVGgZXTGZkKPvXy72TN3rZ0B3JVfZV
VQtyDtOy3IkitQmQZdzmBx7U+Cj7bMr+dg9TfgvBL3wM0uXYawP0m0eUW2Nmo0+32nxZ+ftVX4Xv
AWi5nlEELQsUu12u+Z8rFzif966duD39Q5rTKWxwB5TKgXf/5GeLoLyAhQj8kg+0/BErpx3oJBXL
2qEkZtanoPHovJr3iWp51MHejG8RB3OcuvAIzzLSkh17VcdUBC55YbYD2DRMMs94CK2SkzQN1Hj/
h+dFkDdt1NSdpd87SVyHENYPopEbXCjbeJJCweDsJDnXXnI9qRQYPzuoqnRCxdvf/BLsJY307DSv
mkSznjT5SKbqcwpEJXWbqEw+iAqrgEaOHcHU5WqxITUXdVC7IJvQLGk0NYXBe6wov3sIxAa31/vL
ki8M/9G0lUtoX2V/fpnd88/LGd9hjqGNsJYAlvNniXpqjGhXchrHrukM/sVprjo1r8My9RevCpF/
Vt/bTw6Crphsi2WTVIOzJ8hwkS6W497xu1KXt480EX47xxaX/I3AvkqhGSIN4aRhHbZ3aEm3kpxR
jGF5vwRH6G7pdE8Jhilr2U930FmGiTziFUSr5gaCKJTB4c/VQWvYrSeNmqilSURhtX7xkwFYUQO3
woOxN7huYTDnIic5CIf5LfDxBaouiCca+kFPRbNFBK2edfpxKIj6+sYcAH6sdZIN0vV5J515o8dQ
s05Qe/wNnTVgSZKU//ChgZ8ojqsMICGnJqj4ELyutUq2uXFem2GFpf/yAMw6q1zWmkjMsaBzrJ2A
YICwC3dw0JbD8U0CHN/ZhdYL4SADz7Ss1Ki6/fHwJy2kuDmVUNCLNqIVrT0gSqA+x3DIFApK9Sej
xfQe9A0fngriIM55Wr1EDUJ5wOqBCT4Qf42dxTQ/BwVgcKuX/4ei8M8M9A0AlHLp09g4O+JYgUj0
hnVCVTO9NfeIh21fTTcbPgI+02B3wdnGgrtR/BCBuk85jYfKrocEREzDvBejlvwLyv8yrSDP5yKG
DsArwT3yQKT74YOCrl5WV/d3y2qdQEj/N25mdBtCGrE529EzkyhDfHZk2hm6t2DcC54T7IDMwKI0
ARhvGb73tcDFbnP1pMxW7N8QAdQ1yWtKIxnGC1elNr76og7QZbW8IPj6+LTUBv8tinIrNSLCezQG
cQ+L+5yQzGej9K3AgL7yJbtTdawx7Id+9wuurHJ4o6VqisqrphWEicrxhejJ0a/PMp4ANtWTvMPu
yS5UpiCgqrKB1V/Bi467gWGscjR4X1GwD8cmWU4jvt4HZpHW+dZXrneuuR9Kl8fr76T9o3gNXCgV
HN3PIBFQrNupfaeaPAADwYnPTt0LtglBm6MEQprKTJm8HZopSPeEUqnaeM1id2ubht3RiySz8dSu
7DhUaRzLDlx8jpLbB3jvXxS6uTAP1ny3s9IQwJ+fIiwf8a0R+h4uq4QGF1p2cAfkVkDb9tn4Sqml
ELU82IQHG8URpQ4AlfRYOamVTjrhxR+QwEkBQfIdq9ADQgHfo9HKx6RK/vCdVaGV7I5LD9hXvA/6
UECCkMY6jjBsq4tBoCg4Uvh/H7FHxqAF/oNjfZVdequaHEQaXU7sLb1yujRwMtzlWq9nlr4ULD21
EiL+YQNY2lzITreEYglmAoISixIS5fQ7HLrgj2HVhnnHKb5HemrZ32HuXnmh3m+GeHxn9X92LYMi
ved954tZwKxwujvTc3rjmFUznvAaGlWUu2KwcR4sstISWeGaB/2uA1vEJuypgUqx/gxe44EL9NRx
EF3veFVAYgAWoNaOMMzPx09hUoG6NRgHNix69F814gdqmMzCajy4auZx8K6QGbGe2xmLkllqatZC
mAnViaqS1Y6yUhj79c34NztBcmWmf14WH+hhLxL2Z4ZBT9IUYbE9chL4fw7pLew+/0LDiT5PIW0b
C4gdoq4Y7ItHPnBEZb4D/ONps+CRKQ2Agwkr5jFXP5R8rQ54h2+hAyefaEksVbdMgEs9+Lw0BMDi
d31Sl3L92E3KgECItEV0yXlwCpccqf/5M2nOgkyEjm5vFOElaNz+tVC4CINUZ1NpkhQjAkD+MaS5
eB2hKzWGQA3+TySgBf7nvArmJm72J1AJC6SltBfEeij5DnULjla2Ki5EFvfj5MjFy97AAiwx98yT
GKaNQ3+8y6V3V+isIT42WWZjj0I98vJTxz5mZPomNQdWPQHExW0pxip3NJ0cjLMFBBcYfr4kyaKQ
SiCzM4yhcmhGGEZS8LTQleGozwWsbxH6uZ9un7VFWDsRDLH9FeszfrObUavev670GT6uPKK1y9Go
FDz5m+P+NvdlZiW7GykqZ3Bs1ALbcTwImPT+mh0bsf8+nT38p8w9eLLSb7CTja2TBi0apv6dZTzy
RAYGqh1Zn+ihn+K1znfX59G/ndBGC1dqiDJoEI6sogiT4DGRm0AABaZKLV0dOV99WE5heuGO33XC
h7MUydS8k4fMziBRY1TR2LXLyxnp+bIV1CxZfOQ5Prkp619O++MEBPrWtfBSeZNNT0CsB5d3zxft
oLYdUteeCJSncAYVrodDvwJWhWvTHGiTCdWFxM7z5CG8OLxJuDgoxJuUAWdZmw+RsEwlTc3b9hGM
zeGdq0QJQs2f/GrT3gkbCP+itB7pUxsoi3jKo/kXo03pwvIVDGixuCmJdm4DurX5Zy1Wf+1564v+
AjjOVJXL2b1aIO8IY85L2d1qn/bNdU1zYW+gsNqOjkesRNp1f+iGdsc8ee4MnLLVJfCPKzphTTwk
dWUDUjgYm+i7MqxxBFGhcwKDqbDmTtqInaZa/kHPKXAW0EQ/kEdRc8D94wpk+tqo25fLIwcr5aC8
vtPr8SNinaUB45pXFeKeQPpjSB/fOTXJvzqCXy/Facw3BPjvJ3IEdzem4YkBJ77o486vqNBArG21
Wz5eGt6poE/gbry79kZhR0tvqvkCPeEPq1r54A4yKNP5NSDlyExxXPhIbyRi1Gxrqi6LlNt0gPlf
Swlfej9ZCf1Rdk6cs3Fkqoc+VR7+Dq7nODW9dGh9nYzewl0Qq/LW9lGy2hwVE5bCqSgwKJ5WHsSd
JpZt/KSVRDTAAkIIz63F02Ay/JeWpk0psb7jcmdTIvy2Qtwd6uyqMPW1hy4kSNHlAC2O2+SZIwqU
7b33K0B/C3yVqLgrLqPUHNqsuMMGvBT1UR44iThWybq1clL5YH5haU+tnFxwC2MNZQWiV+KhE7vB
pD2B8NiamgjLOi69O4vNweTjUFJNFZwfWsLghZtFAOoHzA4MvXyOJdCUOSKCHiQtAaMAagrFfztZ
zzbZkBaWztj212Vaq/jVZ11SLsHeqhlnaMe1mSV+UVICqBXWDESHxQDUgoK4GiNt0yZQ7Rf6Xxqg
195D2Ic5yqHPHFWGzlCKkBqAtEH+zH9sK9LaVC5K/obmxZvk698gTT4kw5aAvySHQQ+ct8Wp/CTf
OtMZfGecZCWuQnXzwMiwC2FxJeseXe9Oo1b30QSTZL6ZKfJWN1PK6K665dEPfP34Z5s9Uz3xVZB9
clFhazVtBJRjeGCt9it09Gyj0O6fsbujMT/WWoe+7Xuwylo0pN14m8Qi2O1bafpAnuXqAMAqBFcx
RnnNrQVMUChvXePPdtNjP1PWQDk1R7HvdLZ852NWODyvmGo3bwOwA6pVz5N28UcXg3rkarjDMdAx
WQ5cvhwUqO+YHwOaETLcTiROQVs6LTb5mx06PLP5piuPHolxe2cg/bBZ6M4+nXwjgFIA2u9B7jf8
iNJ3Xju+XpW21E5mobqpqE9zSZrI1i30i2SXzjDxfvoTNYfTS7G3UFf+PmlXIbVtJ/y8dX24wauM
X7L0NJ0Dk9gVrhny0B2SsS7A94RsfdjIo1YFnLAf7Mww90GK0S9iN8Zxzq8e2vsrosJvkOuFzf+6
zpCLYpUojVy02G6F9+oF61azoDJKjehmCgJE+Ccj8D7iSSw5GVu8Z1ABfFEVewtK3lNCjxR26ZEu
o9C4OUfXDFzhE4ifZsV4BpyYgb2Po9x8qodF0a7xaKkYfSK7Y3eTcQFcvEHSw8gpwW1mojdBhy1e
ADJ6ObE1FnaBeZ6LWDooZyx6rgqktlN7RvmS8+vbRFPlgtg2wv2xXBUpSLqVDwOYs9304W6yOzMG
MqRffyI6YdG86bC7DUbPPING46Ox4upg4ESgclc57rOP8tA5hUlOvOHHUcmVEM4nBp1eAmDDiY/c
LshXytKiZKdrySQjwbxy0rGk2j9dAJ3VHeuN8LB/7O15G0kX/grXEGPdnkNkpjC74S23DKZHEadR
Z+dA7lPlZ/8lDlvoA249BIktDGwIDvdu8HY1d/R4YU8kGGSZnylxEIHrdB6BgMm0Go7nOwr62o9u
/ZFc6M2ydkXCdk60VwVnXqPgIlehvncJMScccCwPWsa5O3zKCyxF3MqZAoKgML78jMU7a4NsHtxf
pSqnSSCA9y5p4ACUBbFnw8hK7MxYwy6TNwFhycdsV3jLFbHm1TVDXboIKpB45OOScku730BYHVgg
ZeCLds/xTB2fzcKd7yJVNvqpOCheDEo6JoQOusHbHf2FJ2I2jCTCxGnka4nASj4M0JXD4ojYtgNZ
WdoTHsvn7vn/6nkaQ6NoVfXm5f9W9R0iJR2WKTMKJDzD63LB0gufRpPVapC9mnUtZYrZhubkwKvN
bzOz8JvEwtk3YkSGlo63n/ctdKYg+mzOqj32XwdqHvZDsKyfqMiPzP+fXCarzgv7ff7xb2YNF/fJ
7j4iKFpDQZvoQ7M56SKh25ss7g3zSsnhGsS0K3V/NgwktnMkuh9wOGTgxBF2K74pR1n9Y6vl93Lp
kwh9u1QnmUlU5BtobEu4UiDqw9sWKkgcopHnPbkDYJO6U0I4EW7HgyAG7sc0C1U42KfB7EM65m3O
/wNAe4/3xW1BZt5lGtLC1AbrCnDyqIS4SxAPWARGtTEYddFHp0317DAzRitJXNbgaO/v98usGLkK
2nuTwNHu5/rzhh2ZUkeZ2GzNxn6cRKAi+O+SEkPzI+oc5vRwENmL/UsLvlsifRNv3j2dKtJw3XPK
/uXeDdY2qFrMQ/vCizs6zgvWI978fN69e7I5IGhOZ7MMnss7IoRovWlMDFGmOeJIwSCc++UuojS0
q7XO5cGCRIVsysuHv/pDdgVyi/Qt4kCZOb2RNLVYUNSr7jPP9Dtx44KgKqCmtuheJ4Wj9LWRW5mH
UpEw2/eE9kuFvEtXvZknorHst6df2+LrPugX0mpZBjNL3ptDENLaZH71wgVefzkDVwvOLGw1wyLW
dlFb2ESYonNwxKFcs8EdRHiXgooPtl5X2y6rmBcTx/oBgBjIe87yO2oEbh/pn2MzGhBV6aCSoeB/
z3BIKG23c0HNVsBAwlPu+kng9U1jKzPiz6hy6Fz2QuIz/GPp/ULUPBY/z2xZgRwV39jbLDwt+Uac
N8+6g+F8MadavYGUHz5UydFtX2PQ6O7Rwm18BhSoWOjH0jMWyLYKSSkFy9yzZmPqnMiN8cbb1xEm
fsYulW7VgsdX5rVJf1+Z/uryYM05poX8MXNQ28TtRWS28EqgsYkfPbmz4Pl21I/e7hTO0Ik4MGIf
ste1fD3iixsuTNWLvZn5Ypvw2NrNwlpN+v95QaaGUORTCc+FnMaZcn/e2+4YtvjbU7NDA+/s8Ka2
+QocVfIKawgTxtTStHaQLKdk/lCi8h4rOr/MpxkaiMwlLQihcBdmyo4J2h1B5NM1nJYQgxb4F1A4
tSmv98V87+C8m4kkhQWk+whuWT6aQpyGPCo+pFDpksclrz7X7BKvLE8TWaYO7lYepaU+S+rSeh9Q
KZHFdAi5RWkhwZCE2deDLKE2odSwptzcbkYoaW25wFQPHmUHNcrsUXKY2ALszx2A/ySLAsk9YWUZ
i/U2gOsZNvheBuPwqm8Y2OAeVL9CKdjHzIBMdA4vKETr23eB3lwZgjOkwUzp6uLOsiTA3aDAmFFD
IFtGpQZs/pJq9WCe4wAYEihDynxAd15LnijxFFTLF4BPRJ9p2VvqZkQ/3blFUt+eOstyIIHhzdp6
I/OpLm5gDaL7OekAHhWtY2ZgGf4+fOdVnBRaJSWTY0ilmWXsPlXYmSvM9o0dDtm6RlBeUbS8qhFA
nVOjXh+h3jPKI0eUPQ4iDJMWSJ5sdi6KxE9mNAOfqRcFCiIFLHlezsUaTIqfDsSon+ro2bfplEbj
aqfN8BYWjlPmsrtqWEJl218d78QxQMsJNm0FGwcxVOZVnxfN8cXbSrrxBZy+4AGOX/fPr6YQ+KtV
PkOvP8Mn5d/FxM6+WJ5FkSFAgORA8suyTgBSmcSFeo9qHV8YQ1wM/MDG7A80m19B2afll/BApM4S
bjoCbArWb9+FlqNN62wrNixNPdumdkN4XSCZ3tfUVpdGa1o1cbR5MyHBwhPpBVMzZEg5TCWyryEq
BKVL2JuoQahTC5iYa+fNbvDoqVNdqKvtMERwR4zjNPfCpjU2Ob4+I30kJFYJ6chHqjNSVHdjpqkp
vVwhWh29C4h8XNep6G9MywP+HnxyAWYPpsWRtGoX8qexTVq+vjkmYISu0wq3YhV18j1qeVybplvW
R/B+u23qLjn18i24kkit+ErUe/QKzv70a2TwhC5l1RZpL3eKQ2jdo86wGCajF7ioV24QOgRrxjAB
BeTWcALKv8Q0Fk3sBw+61zxM2BnU+hJWAStWT5y35+6D72cbMHpN5ecHSr5ZNuB38u1Kc3RYMyr+
+WWCpsJAZGRSXlYD53z02IYbNoPjl+U5o0YSDjy8aREASpKf1vxUNTYidcNR2+pg4u8aYgs7/KiQ
XJ3WIQbD9Ov7aaADUzy0a7u3Otcf49SlbecePhBg1J9aoxdYvA4bjSC8IAF+MmRndWeqjIz7uCsg
GUFmssUNlLCX1v2J8Znmzc9WZYeDwXsF/ZPALCCT63qSTnwY77aK9DK/I+5C5/KHRRiMtdgR8lqO
jvyJZCH53WEj8ScdDvkNL1LdZbb37D5D4oxzcuEG6zrgEyzbl8rPKTu8gwCv9om06Xkz5bqkQVck
sudSFKRh/uTc+Mhj72q3CwXBpQD3VKpEUZyfG+XH18gqCuyRvQfPp0pNO1aRYbO5gy2eCCW3reEO
gkCR+nDTobKvPkQmyyz84/y1HAMNBZlW/c8Z6QbVFzGGvDaVcccWjtQ+Fusa8G1knFKoLPr+SP64
LhEGJBYBXU9KS/E+S+76oUkN4RqBEprzKLI75nb7Pjgu4unBaNUEq5CIKTE5B3J/Q339m2BIfDtN
fqUBKhIpIYn0WuAQif17tzu2g6p8/nzj+XAAUeJG/gIbAU9+ADHMnHRz2xS2KR6Bvq/00/atBdbn
/oCwi7hlXvvjrNjGepbyu8V3xyjnINyF/0L168mmqnRCsr8rznshlayTNf/iArqXOPVPu68ASF/r
RLo5n+4bMxPszCyGXIAVw5BEyGa0/gknmgzsnHnDD7lxO4WhcGPpvAUsM/YIdfP8ZbHTJD9U2zKE
LLg6hRiQX2tz3nhFYst3hc+Q5MJxt3YIBEv25chWVCncVAokdkcD2svy7+u2IVTAxeDtBL9OQs/V
9Ckk1OZUs2fpW/YQ1HqehsxoOG1fX4Mz/EntgyzkTcM9J6dx134cvN9a18ZazM6a7vdvCwUjnGem
fImXQaR4MDYGAFCbPpZJjDKWQX91sI9L3lLXsGS3AKtLmyDoenqIBNtZzRTkmeSzqzS4C9BrlupA
TO+WpMkY0T02b+oh9RZwqkv2f5wjy8ImQQsDlNFudi1P30Tiw+daE8QS2K6EDS4iP3auG2HtzhZe
DOW9XSo5/kPNowjVMHJa9jMmUz+zLU9yHEy9nafwf2eNYe6TdTShQIzoV5/e9HE7hiFXHlj5vTEo
FHO2AmpJ05iSP+WSjbybn5BOnVLoECy8UCTFHqmeeQcTFwuv/4XQD5X89qDY9xsmqJejB7KbFIhk
BaqLE7K+hhMkG9VIu5u27axwOXe6SwyZ3dYosvbHzUrqp5epubEjod9+Vyw84GUk1U+xy9d2MPna
OHmmkDDxfegQ8jYpxeYj4SooRHlEcesQgqbevBC3XRrtFk7hJrspmEY6+4DrrCdkacc1Z3x5VIm0
MvyKrrz0rhBCbjAavTdh8s/STfS7zs69Em+/Qpc8Mrzj/GKxwPOOSNfKKdgVNfKEjt0DE3u1AbBd
hd5bPGz/G4u0HXZ4g58zD9ySukw6wJaZsVYuCsdRT+6ZnoYMgkNHJdNDmSSyfsviSmTt2F2SIlKn
MdbST/A/9k7iydt2M6ISNaZqQwdyQK/nrfpP5K/ymQ2qjb5eAgl09AT4xTfx/HVe2B5ud/Yt3tvn
MiX8gQChnF3RTl0lHnwsPvY40itSyiNIgvwtXbndIphOV1TheX1BDG0C9yutgfePwbkHX4gnPEgY
IFJ1rMDS0DCdJhqsxNZfsJpkMN1uVD+9HlrWPjEgUxuafEXtrEflGx8nwlVXFy+IVshc7K01zJ2I
W2ShYAL/YF30AYnXIIDV0bomqfCBbidZi/EUlkgLEhdDVD5jWltrzxmINyCYn5tWBfCmBqNRaomH
rspHUobfaz63Oetenv6K6gzP/UhinKALpUgWV68XZQB5HmrDlSVoDCB9ptlpjlqcWf71MO9/c2jL
4iUis/Ijzp2REulR5ZuRn1317Et94WIrBXqV7iYGT36/ySv+pHElLJczZxPm60dAk8pxkZuRcwQg
fhNS/Qcx+dyxtMhNw0KnReO6QYF4MI7QadfrEMna/amvn/s7z87LsbUrLdlE4bDKQdRekc9OLYLE
fUJmQeg30MRgTNpo8tWQ+isTdbCJS9q4T6jdhLZJ/dq6SfaLp4ywJHpUkLAmjjF52U+a4X1JqyUn
0kOfAsNmaGRWY3BC6n8JrdPJ4ZklJAKmjWxDu+Pmlc+vVTU4M6NY2WhdCHo6hOanPhfcMhvmugC5
4XJ8QUwNWdYzSpnIPjof3ru92LUgC01ne/7/HBopfy4Rj+pE8HKHQog35YSurhyw4QqO3kl+t8dE
P5CM3Mn1JfI4o9lqbc7rW+inCJlbjdky+G6VZzPZ45VfC+FpLqDsFyGhroQlRHnZcp90vcYx8qK6
4xt/Z9hWKY45z+57RnCajn0OJnOxAPsR9WuRJzcXKR5wi7Vszsb8PzUGTG4hxCEEHunRGC9N8yhv
T2mj0Yxs7gON6m/A1E6U//RzMmR7sDBnntVPY2yPdqMLm01OlzedzAcvzpp1kau8KeEBHgXd30io
dSUUBeCR1DKzIIQ1FQAH0tpjQMISTdCXppm/eOpoHL8GTGRJzYg2brT0Dr2TC54fyzY79v1Y7fmA
qmZ+bdXFFYkhrgttEH5e/KXd9pWyDtZEYHAAb5V97wbdinYezqUha2T6b8kApZTXJKGadpuv5exR
WTEJN/nJPuS0lzS1NM6b/Lb6wKqsjTd/VJazb8MhRR+bFF3gasyaO6SkpK+GvOvG4YRkgyyziJZf
KrJCooTSxZxTg2l2UTuurCdlgK+ldHVKBaRx2dAqpQgL3ABPJjhxxjtvsXipCyhoouyBXvOxCKvx
UCAn9jShxXCaKIaKVaIFElbIKD0VuO42ygodn9OaCA4FtxylnUY3V5m+XK9grZMeh8QI7O7+pmKl
bd6d8N15sLSKbeSnmwcXznuPZ6FW5lO+3LM4DEOK4SFmGK9aLi/38v1U9/7SGv0D/WuF2gegA9j8
uENdebHiZRTxGyos2fj6RL8xtqkOtLpJw0Zbn9nUhnMfrtOtTyxbfHw7WAHDHYDyxF/s2e9iQMku
KwflvdS9K3o2p1+Zw3edjPPrFrIGLKgrsX2JRrxK5gK4g4+cb6Qrg60UG8SQY178GSA6sfjp91pI
SSiZPsekGBavqIKq5+CqW1E91E/NykWH7QCgzRh7C9wIoLB89cCYbsXCri5iCgCwpJyu89C2QFJg
+JUEDAxJdCkoMaz3rWKgqb2X9YU9eMgp1hWmgwuOiXUzSTTpNrSakAO5zyuLtwSDOF5rBhUXP83h
mS+4oGu+85p4qXHHN/6BDAhzS65/doojqWiKa8HxKGOmvRqHqLO7qJC38x33IqD1m87vUunjMExB
P2CSAungmFHc+bDTFw9jCXXKw+Dm5zXzTzT4wK41LDQHflD7yBta6VeS3L0mkGEPwrsvIp+44Qo+
x5XvCNxyMgo2O3ZO9qtBP/tOcdhsOat0gIdqAf+O8jTg/zfJbY6CDacfpoyaqjPW2Rs+dkXBLrnk
3piSzGIOuq4v6M8jkv+fER9FAyXheuoP9FRvlaX1GFbVbReVsbG1Dxct+IXLPq5I5nU/n7qTOuCm
wwMYQJdHQyOTUuMTiBo4jUWIner87vTWeMCovXtsiiysvr4oQxcyWappTcDmNwD1dL4SYam27I2t
9lHSryhVsdQeNgrbbnO1niQ/nAWKhIGlA9aV9mmuMxZZr15mjzv1Zr9ZwEjPUuBgFVugMm2Ek6s4
JhhFOVlqQ4E8K4GHx+Qk+eM/eCejd+pOIJvzdpLgzTV37HJm+S8bKUOv6RlJmNsg2zCUEBEkvt9r
jQiuo32bhhnE1/eDTTKy8WV5cf5Uz9KrMBaUzckxvVWbQiAKjj9uhwyGxLDgp+YoA6B5hnYKnJk2
m8SgvnEIf0tFEIM5ev9ZYemFnDrNCAcUkc/c57HE+uxINCnM6AbpbxLasAxZZ2gWN9W1o4Xk5cDo
aPN8/j3PksWro+Sw6GIMPZUaoHbAS+iaj3LuarH7zul9wMZNYc1YbbRHfH3m6Coh3lLLZVW8IY5G
JyWzo+DCa8Ai3Kx6DRNRET8nzDMtpqhkxFsdlPT8f6Nb8J6hToPCiKIiMkOrBp1KsB4Pq2Z8H8Tm
MvZrtusA3q00vIkcjGUhXLoiDBM3LGkH2bCUNG1PPB97cTWK9LiniO/CtjPommgoNJFBIO3Sks4f
7n4NjqbxBZBvWZ4dSpgEw3gmwWyTRraFr1FNukSJuHErhYRfx+TmWjuKsOVenLUDq6tf1dEtWNlB
ynGG2TNpJ5aZ16h9uLy2FADuEHwzHxamALeVm6Gg/yeRsqV65DQYRI8Cf3cgQ/4cG5ESvVf8tNly
C4OsjkCtmo9xXWKPWYqFgnVFADHw/NiJSU1Imo2b5ikztqaiK6mAtC21Zqyt9Ss0x4ckIkQWj7up
siNB7N6NqlDsDu0mv6hsdlUnVCJOJ25sQHpKPnu5fzd0jw9J/371fHYJ9bXXHiFy/5n7skp+gONo
J8YtyBeV73Lf+xg0oYr3pNHLGfK3dRu/7o/g5K5yOpe9tKQOasUJz/onlraEyKf4/HIE8P33Q4BS
swhl2pA6AHqPWSfRowu46uXPucL+OK5uuUjWMyugWZRm0IqZQdh1QDFCfYxxkySPpQpXCwsoiTtr
Kg04DEA3lI/v4K3mHMw1FmXYxIrUd9YoIvh8eALWT3QrZg1B6UuGBFus81Zr5sS4QZAiUNccZkGb
7Fcxz92zwnJEb/bckS3mAo4JvuNrOMVd8o+bEhcq5uf15ZTdIYh+q4qaCFmIhScZhBzhVuOcSAZT
cApxyhcipjvRlGJDT4WiV5ia2YYeHChc0/dyeLELluSC86d1NLmnceCZjsBNQAAwNZv0Z3XuKWUP
ALNMyBj8OP+9B6YMupVo9z8U1DTz2pyRIkWD3dPVwEfNgxbBpd3JYwfdhDbrGdHpkah3O09FVd6e
npT/2g5GRQcLyJH4fknJWVDjjFaP+sHOcNEuO+1FAokEIyOUh6cuOkQJsDat+YamJl/Sx790XfAU
K7Yy/bANyqePvKEsbWM39OPewVyZ3spwOmTd8buIsjAtA3yAJAP0KwuXObP9ApWPgmoEdY+hpJzA
Hri2QzJE9mmxWA5P25u/lUGTmg6yqIN8iSUb4OB9IYzRcK5aQTG892hKa91HtZt8L3wIqhIZQgXr
eDAWjsZKZ6uuPYuKcy65jc1ia98GG+0AQzB6utUVeiPylVtei6bnyjhB6Lc4zxohxBixuM01jua6
+mmOtaTCnH7REt6qARy5LTJAMq2I8whOXfb6BGYuheAHItxLlX1/SSpwAC4u6KDxs3xE7GeUDnkB
0mSXhN2SHNXDLxLdDHycSalACJiQ/Xq0E6PH1vbtzRAO9OspCesWhogBRGsUa7ALbj0dSZdHcHj7
9jZhXRJpccDE844xmXcyKnf6N5T7C//8rmtaytEOiEs/4apTbdvWaaRefP1Qhe7G6cE4nHgz+35C
o5zgv6G5SoHhsGaRElXo1ByJ1Y/KBmfR9k/cfodbYhtVtoSJsDfmBXGc9EQyZhkMMY8dCYlDsreZ
yC7VWOx9aBRLH2N/cnOmCluCsxBIh/cJgMsohgTfoA2BNYbsn9VauiBo8B6eWloTIWjWuJh2IvSj
N9yjVAwpifop6X2vsYyHFEN0r0JiYn7zNtguZp80YiCGJiCdBWjW3oQzJEqsQ1TfWAuKriP/oT0H
RURDcg87R7x8VmPG9/dR2BU+8QCD51TDns3Ca3ylnA+GpslJjDVTM1r9R7e9VMEDICxcMWKgSSZw
xFrVtoJ5fH9GFd5Da/F4EdXp5Q5HMLgMB4uk5A8VrtO1CQeaPvC+5e5bX/ZQ+ZDW0XM+vK0FAKhU
kzH+LB6D5qela7gkx7f634cS+jw6ReN/UquMZczLy7Gqd7jO9ElK9Y7cXs5O9/hKlQ+fgYl2HH2L
6aDgEVvNtoxDfy3GNSl5BQYmTiiEZePtjcXonbZGG43+RihNwD+mmjd0D9hc4eAOkBVtPEg8CNRH
NO/hNKD7H7nuHxBj//tdoHpgWyye12t2ysraYdITer67RMSwgNWT3shQIxX50qjvaPxUheUJv9Fb
3QFY4Bi9EZbVnA9mNQqzrZMxfIxRjSKbTyL/5EJHpHV1lmpn5+HoiKxIQJTAeq/N7HMl8nh47bIj
F1SU0Q7gaehXNLGPryeoZ2FpQY3l3yapiKvKX9wO2fMsDC3MxALBzr3rtsb+1Gp1tVtNIszoEJ4T
MVDKp2Ilpsa6cj/Y+vWziifhzbFFQLl5M/RboCXgjp1RgoWHcoS9Tg4nfX/OF8XhG+NdvWL5y1LZ
XCwdKQI4BE8fxjzWd/Ye5cutoi+FMVzFEvDnlJ7fw6SKcxdDod4avx5p8gdcpuMs4RlQOMYopb6Z
Al+30uotDmaYluk6SnMOcJuEyEKYW5vLV06pCSv1JchOlSm18tvAsVGxwT6zV68MSRx/8+kYW/gU
TApGntMEjsIGWt04UW7OyVeRAeiY1UYjXV02GTdz+U9fikpKH24ZlSQVKQxmm/iL96fjD7lkktN6
vl1BGsRMu/97d5Cy/5Ua9wWUrGMS4EPdZVhgGASNMWKuCOl/n+8fIMdS2HNuykJUlvfcnPCYW1pA
HgS/jpnAJF6kQAs7PPAf41jvqapqC/V1//9MNlVrlAN/eZemrMHaFEwFV0Jd0sLH3qTbyZcIuxpe
02sqmFcb7anH5aOiFeFXVbKmpiCYrsTVrYIHuMRQ5M5Jl0x3xzxELEii1u7FB9HXFKca3VoU1ZDt
eiJ0TUNCQtQXXID7ZEaHJuoGUrj5NS3T/oy+506/keG9u7Y4H2iSeTiOGc42zhklfvf7u05r0c/p
J1FPouWaLerFMFlO0BirAvH/DXJl1RBx5GU4r2R/YCkfoLoWszuqi9+mVsB0yTEPu+VHL4Dfq0PL
1CA54uf22EyKT7s5oUjWqCKV9agiaF9FMgJf20orF9/0MhoPnb6f8Tf6CPYt3qHJd6p4wdIMPFN4
SB3R0/rR1cWo+dp+hkBH9GMb/v6pi8NkLKwsNzAOSQc4sKtEnw7e/E4aCl1XulM9fgHwd04c/bus
kTO//UtxV5Wi8b324WjeE/3gOsa0Kbj9Fsbxyhh7QQ6DNW9ZXxjZWS7gAnJrtlBzBvZI2FoXm0E9
2GQfpgUPgPmeyC8st2q60y4tsiRMI+83Bl93wDscmgwwpmwcPeKPR3sbQxTpHN/gp6BsMnkx5JIR
cK61FqCYmQkr77ACWPRftxTea22p2Tsc6g0j0j5E3Sc/N14akxS/J7FhnklXpASz2c1FiyZ9Q2LP
+JCQp8g2EwZ3STuTl/OgVWRkLvEy1ItEU9IdV9s+SQVriVrMGQqUBqo+Tv+eJVrorRRpHHIo8+cu
t/iwXeqp5bUKOibTrdN2fHj4ixf5ui0lWLOJXhPqdETLafRDiwnlgVAqaaH824RREKs+c/Gf9YU3
ztyDqVzz/9TvwzKlB+hwcSaCtvf1YGkQntkSh/potEzi7D+kdmYXip+A6yT+fB82rj+eI2iACfKW
uTE1aofdHF1NQwmMnFie6UF8dwZ50QPFuI/b+x5IjYY9Jy3yHWVvqd/e1ow+G5q2uWzH45wFRtC0
8NnEQca/FTILWbQU4Jr+raBQsIAJN8VQiG0CHvybTlKI7HsWgnpymKOLV3bXt4jAi2SnWehGDKjP
I3yWAiSHHGMFzflgdh8QdmjaK2acnTlyqs8y5+jPic3xgn34sKmX8+5wil510rU9/4QfXi1fDMrL
nDSduS73B0Z/6PUMIYpQwHtnlaUNXOMjq6q1wXjkI1ir6fWsX54i4O9Hmu5gLOZMCNafAOerwDIT
cVpsJIvDB7fCACgUXfr0aZOxkKnKywQPnuNAuzcqQrjShbGueLjTF95IjPiKfJacEOo9Ff8xCxYY
HkzvG6c4hJnPBQf7KwusMY5TzK6Fsfwj5ZcBPtRsoe7siuYT5e3EimGzTagfbliSkqC9pKLM7gkj
3a8/8OVSOSybZCtx04n+/gaK6l9AQ4M5+8yMH8dhqaaRgdn0NKZWr1rEnBKm1syVuiGEV+Kzyo/G
Hm0NlbqvFrv3DERmMGVy7WNO+1b6RsYE6VLgA3gl9dXqMInX+w4jCSJiYzS5T4WoPIgEaPoxrxxR
DVRSlEfvzh1qx6sDKG/j9hqBBAR0ph9lNmZWi1qn3nwTxojuwcl3ngrPI7nLIPXfvl8U+73NLi9A
Kdaf/DzrL+cBAksCI49R29bHUMmDOFw2zH3ZsoHSvoDXr2RqcGNhzoY0wbw6A3EcUt1F4/O82JxC
fMB5wQeGzJdDyQzIBU6SdgoijdMzLSJtDIwOtazQFFXxpShfmiJpnLuDLqKKZQVGnBOQ1uklnYAi
DyzQZ6tlql84waPEZsaFPwsZibA3OIXc/IDORCaw8+3xH2PfI4o0PbJWlpNr+P1omDhABQDZw6eT
OQ375K+yJ9iEOwIdEYnjGgRhHI6FLOXq8O4Klnt4q5MMq9QF63GfK44QDVf5RYBZwvohV56grPBD
G5AKHxzd+4O0QVnocIwG1QJOskrlGbgf5Amx8abG1Klu2Ph7xZYE27fkWsB/nYV8Oc0RHRM8C+w2
StpswH2bIZh4UtD74mq4cYF/BTvV3SGjhuYBYUsMQxbU/eZDEFK0/CfNcbtNX/cFrNBeo99lu5ww
n0jRqhMZ3UwY4A1vgXrJzcTScbWf6Zs6ufojBfs0hbk5j2eL+t+AsN2LuRWuAv/kywii3fiBUDa+
uvBlkjnrp29hKD7ceRq37nygJPaqnrKPWBHG3mBfs9/9aU8wiWL1jLSsPQwGudAkPLWtLYV3gOTI
eYiSWUEujtZbBqYGbN6+7iXfqR23kf+nb97//aKG89YhhexVNSkM1IrVdDRAs8MXiI+Q7XZM5pdz
0fhdTYmEeAJgDFrvSRiv9dA+plH6aec/ZDxOMgYUyLXcU05V4OA45uGy5fGA/HWSA3p23uH13l8m
2rpCxsZO58HFl7EfV89H9LV1VYUGtKTLIJlne7Ijj+Ij+yZ3oqLSBiycQfVlvmXxPE79IGXOksPZ
L3mZISaSEt/EJu9VSb0PfypG0ozMBL/zHFQj6eYv6Jtk46WjM+kU9QXNWvQJgA3pi14S5j5wd3im
Q9LSR0WJFi+wp3HtD8NaQINxkT3C3jSvI8ryTWd9u20EoAPp1iYO6In9xAcKAGuW0nhCR9Q7bcTq
rgJdMY7GEc6duMtI7A3VCGBISXN2IrA2hteIBkFCymuNAm7IQtPKUKuiuvGY/txau/mVxmRQZtMD
f1B+4momBv4XoXBG/xM42iAJX6rFXu0DjUH86Y7i0w6BArLsl3RiwnC91joEKlIBMTLIZmugUjmu
TtX4ZitIVvv2B56+gnD0iz6Rb2Bz+nDqO7MXqVtaxIHds03LViz50sz+cCwRt0L0C26qaGYfrYsY
nfzCiwip0bQlplatQ0AUmNFZzMy5EuSUvN+SXMMfYuKM60IDEZh5w1WJ/YmF5sGDLhIkLdR8rJkJ
kCEJGCSS927LPrBClZwceDY4gXq7dnNIeVyDFFIqZy6Rc9Xt3wvfwgxGGcFdcb6cjIVZ4djy/Atr
Ausf6Wt8gDV1d0PYmHdg4kIr8a2yhSca6EqtfcuYIo5BAnIut+YBo/7Q11okxYATSKInxmPZrOTZ
m3pP6MhReQdLj+TQMeEGhRspPlG2EiA/q6ucLVnju/22FM8AwVAigpHfESWi8DBnXKcijpGxzEiM
To5h/Z5Jt3rHB+umL80va7Cv0YJwjF0/JtLggrWIFXb8WF1cB7izt5pWZCZy0gbeIplqPF3/QTha
1mqDSjfUNj0QDT7oMQ5H08FxaNNNKBlLxsosrKtYC21Kx7kuaDe6K3ObPv839zJeqTzgJxuWVeXJ
Q09MgPKOgeimFLtfnI54Gc6lOs2bR7RJ2mYczQpS1ZTNt6eMEHyFIaHcFb5FY8LxCx/Kxo3pl1SC
BIYHnN4QONk0nvZ60W7+1DJZDB7z7YRJPsPwv4WclBpdsUFgEqMCTlD08QmmiNsX4WsRNAnZBq3P
2kA1W+0c+4e8jf7vSkFDLwiWZONwHWFdpVoZzaUoLIWsTmGHkVlJv+nBCkTfFky1jYURfevra1Pj
tsLIwBo6lKTdLBdTmXEuIdzL+bNBuQHdQFAVNMfIwtXvtyw5J15Tn+O36CUPoUmKo1UuugAbEJ6P
zyv7kD1rWaEyU1AiqCEv5t9T6gBNKCQ7AAuhEMk+SuBRuMMUyVOe6rG4oqItGLuLHmVZyNnyAVMK
OdvmEU+5oCrRdVVKqncKoj9wxSyhA4s4cKrcKc8nVfgTEKqlWAB2s6dPhTHUCGIgubSePPjyOghE
0GcZ3fbAQE8bByYES0G5eQBT4znVtF/BERyO9Z3GkTeZq3fG6BRfMO9MqQcZ+g8IxMco5Cf5JM77
Md46aiMgTZv9upr9ANLGGRNVRb7v+TOlq4y8JxU9GNKaLikd0BAh4S/K3l4wsvViaGfQ/ZMtl8mc
PrtRf96ADzNLp7VnogwyemUhGON46RHGPfgRz0fIIe0/HqK3cuqARIesi0JDy25KhVSeK7m1F8Rq
QUYnrQggpgWcUIRvtYKaO0TY+uSth5Rzi7C9mcthy4ToKavHO7e7TElk+HPyIN71wXE8xtMGY/05
lxjxElscg2l/VdBUUZtiHqmCKkLNdEzBfM4D3K36UdXX7rw5Fk247MVRjErIIQLUHtvxBHleqcey
ihiDUiy/M8Rpuuo+uXXj/aXwmCHWug9We19R0Fi1rr84ZpmTKU6RwlwakSh5BNKVXQJjtz5VlJgJ
u2wUDfhiefxn9BuylsNxNRh8ppSv21jkz73TzV8o2c6bF5Fd4K0yssbrJZm3NXSOSkZohjDawTjw
pck7wyl9/bOW4zTfqBQ7bjdJodwO1JugcDS20I9FE65ur/0a2gnXxBiBqeKIDOvljatNcr0PCw0g
7nKivzcbc5sahRmxgEHBn1uQgX3LxMX/FBifHnu+kbeqSg5oSHWRHvDk7FJiR/5FCDSfFexL0JLJ
CUz5p7UgFSPpddz/DIe+JkCP5snosHCF+K5gLPM63+0XmJoCO7SlxiBvu3mFb4CVcYvrwCwg/r3C
De7gtD9ZhEFt67nJSXm4J5bCr8rbLL7FDgbUtJyLIYW/3r6PA0RK0nSVHsfa+GA/u//Dr2xY7jm6
ld4jVF1T5vbVq1yCvDPopIcWUHqRBDGqTnbMWN7nkphrWId3HwLrK7boVm2BNcHfpKAYsjKDUS0g
VcaZjlCwUR9rL5IopvB5Xg4WjHhcurdgRlmobYa99eETu85XcQQVq7tnkpBWUOg80TnpDFo66Tkb
EiXZLcjNuXgQ5kGLfbMFBc43Eqg9X3NNxNx5TMb5adKBP828lK7cazzyE7jpBWrrNK3njdoqs6cT
TjebV9beVHYh+kGLA7zjH8rAHOVWJ9y0IhxiIvMZBuSSfat9mtCbOV0Xc0bljFV5W9W/UMqGR+32
T1CYUmj6W+q6bfQcGSsinkdd3eunA+F4bPUkJXJSzIxSIr1FnzbnQpfWE32KiWnSATDRLgXw1j6O
lEtHHeYqAJezVeLT63ih7yioXZJxe4RCn5czi31Hi/PCkRNdHD0BpnRl9kb7FhRlgIb9BuThHByk
QOLjhnEoZQs0NQWrVXXjYAs3iRuLX7AmjR1QiXvdqvbGxiam44MwGKtfB9BZj05Bp+Z2Hw0Ywepe
HrfeCYVoHedh+liO6ibpCo0ZUMYlRRodQylce+nOgPu9qmOb7YWfGJsHi4fKeo3uvq41PGMS/bnS
K1TNzfCMHTiMGn0wgKYXwaUkXUSXMHhymEBJ8gNswzC0sU3J1SFYJKupUUByeb2v8J5BcunUqhjE
Mn7jzAWuWGouQmGEqWohD56T2K9D6CWS1UPPbKzskEDkiUnO5r5R/jxd3lnGhWg+4wXPG4RNZrSe
AIIwN68XGY0rNonLFGkp1EqhsNhaw7e4Bxu8jCcrxS+vJORUz3RNSQl2/H27M4VvDSNETgaM+D86
dJHw/AdFvTPbssr5OcesaVoaH5l09QRWj71X74HY79iLsoEplg1TBbRsZ9ZTxyUMZuj2oYdKpL4y
QtT90MvnBMxWJrKDnctbCEixO6vvmyTiq5aRF9tN+Z1RzZuVtRZ9NZqe8VvrADXAKU3FbD44eEcg
Lcov7g453+j/31BMB83NF3O/V2nd8X/2qd91ABQXuLBT4ar5toqeZ8OfOzxmuSvAu3Hb3ulivpwA
jbkYRC8++7wHdqxKyZb/S7jmbSrpAQhaJ5BLJsfXfCOvWyj7c3ClrE5dfRqhSYUO8LLuIJsQtgoa
ol0yd/Mo+i6DwKWFhxvABzpuSOA8YeaJKRAOd/r2WNctvOhOKXFcD4lAXDxLQlXzOx7IY0dUO/Ed
9f31Kyj5Ivg24QnOWRBbueF1ldW1BfsxACtW2i5XxtPlTkrHNFfX9ZytBBJgB5A04dN0v/cGa7T9
2PoLIwjw/Lrk7aQxu4ZhZR4/wWk3nk2fESGbEukcNgSm22SvWGuuM0BM/dliDveIJlkanjYj3eZs
azFgovKj69DSvmzNLlaEZQ+0LaxyO0uzTPrUHnnyswotj3t1WHglJJqo5YoGtm7PoAqay3Rl+TQH
gr8vqfGw9QJKs/x7vRdY0DcireoytC3WPbCDclxk3C474Xm4AIiWA7CjXZyr+J215JGdjY8htCSn
UVyJSM5mRY41izOkWrKYPFpIjF/RNlW7uWoxC7Srmbdig5LczZYHkPASsWYSJD2nqmYjJ/uHhQy1
O9G3Yih/IXsnBloGdfPtruzk9HxYtM3NHacVQWSeWpeUe/PteKZ0AAKeV3DNOrKAXkTkcOqivUvm
ovtijsrEdZGiDZALNjFm6zOBUkeJSeAuIlyKjkebL2m86vkuBtlnERC7egR7yjEm7rm/UwKzyI+h
45KTVAikGJ5Iil+EyVrZZGJQdo4SI6qH0oZvDWnJBywcyNCjXyeR8pfn/wU2P0AuO1XgHksh5wsC
SSc7g14mRWXa1gBVm0ecqcWYrCgXw3MJcmcw7pJqP+1aoWV8YRcoZSSYvAffhyhForEvNqe8XRNn
fBINnKjI77gqmLoEQ84AN5xNRBTqXP5J4qTkqzI+Dj2bd8SNx6WVaRt/CHcWO5MWUxjy8FzkVDj0
CPj+3AqE4Yezyo+7B9q6URnLlYyIX6ZnrPOpw9kddujuhSUVXdtDsIMBNhQrdO51pu7TDaP2c53n
4utQLKHuT7+wdk572OWxd9W0M6+zdoE50peZyCz695JnZVS8S7tsviKuL2on8VIjqc+bg60iLjsT
pFGkychLCx3q9NbZEDLzs3bCKngc8iOdViggJDEV56LOtyn63JaCs2Mt3lyMS+V1/Fow4AUl90Lj
UKUJ//AeQ6XdZbodiQgDBXlf+VWNBeHOXcoekxXldcKrc3kO1RiH5J2Vwzz5n41YIf6/gb+q1v//
Uu3Cle2ceeNPk3/rwxv4DmQj61x0UsUGcqwiDuBL5A03UY7L5JuLS9Y13DA5lRxAPQ+RnZHGFCsS
daWF67Q3BWZpmqe5T2vYZWfwfdAD0D35DWMMcnqSBJ7UKfzR2Ia4EwUq8YcolCUB4lEzdDIYRwcq
PWaU5xyM7zTMj4E2l3MvAGtiDVHwgb78rjQmlyzyd732uOi+nXqnaS6WW5Lk6CgdDRqj3NuMjcbW
xIv5WJpMNEz5FRdBJzKaFKdStK42HOPqg1CNzg2YNDS+IVVY0b4WUO2QfFmR6sHf9dbXl1vVN+uu
fTug9im5Lh9iEDfavFQAuXsa/qp4dK54iW3wPnaSu95La7gN+UQDibYqGlNO2nIN2KwuVE/VJ7nz
jBbj4IaZwewEYpqx+yMMSFU7vZK+t0ThjT5QYcNXlFGDC6WRuw17k5cHPY0IcYgpspyy5NPVilDo
gIoDiYYQ87u5xQLbU22KpF1jbtRynljEOJieY3n1uHF/3FJYUWyH/xR3vei+/A4zQMqjnw315uAd
TZyXaVNcGWQAexO2vQtoh0yT7OxUK9MGuMQZGLl0lQUxlj/RY1YqFL1uQpPQlmsFkqx7vem3xSC/
bM0JKtWUyuhpddOilYbjCdCKNlTZuUMdzn8751j+iaImqv/l83IRZELzlP8TdjmrYbC53QYelDKy
GGIkyxHWaECsHVeYrCdTjyPNOkKgaouHrHFQGFG3G6YMDCkCrCikMzYBZ7gTqIUuVDfgQ3yHaDdB
b766KeXVQrHXevhZPPAlKMNE6mCVUyEmg/c7HB2a9n4fuj2cEPTGIokxcOY+XRybm0Gn8HLZyKMT
KN9T/TJ8YA/akGRTVrIIA2UGfp6VFmTmccLObO4jvghsGXBcU9j1HA5q7tLV3ByVq/Yww6DLwwJh
uaI+ERrbSrVHr0LJQ7JnFsZvQIP+HyBh/gJqDDY4Y1c5pJo5QHwEeWhe1D21CEyka8CXzjsVfzF/
ZoMCNGmuqp4phtkIOOkhb6uYh2NS5EOhkYeI3Ybksd33Zg3TdgSd4+YXa3zTRVAxOZmGklEq2smA
pIYIgjzPW0BFrhIpKeNDvZ1COKOonTWktnsQKV1WdTqPjg+AmNWqr1Mibo6Cjeg+PL89F1RCGgPW
bTFM/i8H/ovrfF8GMSd/gK4BxmVIM43mvUS/v26Usx5wx1pGbDqGtc6jPs/gyd++doosSFRLBB1K
9e+9nXDssolIOlQHJ/k4ahal9P33n9/cBzKmm+6+c6ecIiZzV7hgU4bRa9dF8bCjPh4B4Dm7u4Kx
8bDlGDgLuqCso2z2iIs5072AaB6WSAbP8Jr2zFX4qCQGZRdslej+I0Lgiy24QDgAarlXNWscemDS
JNFUyH0zNxtfzuQZo5brEVpqgZs5PzwNaFWw0OWs8TDW8sTxMw3483olECHO5iMbKOhNQeWIwji2
pYSJgkdgW2PGKSKYdTq20apHltui1WW3iqbQnBm+hKYmZfGYryCDGml2tnRo3AVikqI3Yr/wk/PS
wdY3zlw7Jkegbfd1pvcqGK+JrnDyvZQ+OU2wiWBwImfPaCTOfshuAgYuVvra10I+Arg1kO1BUYBC
VJLHPPmPlAeehGnQAI/LAAkp6S/zIVH5xVLTj/zeg88soNnsLvYPX8SxzfGfXvNikUvaBrTKGNrd
oloQBVdocW6fudE0C9kxsNOk3/pjtG+/sOR1ssFvbA251r6iqb9gehsMJS9P1hUzTpGdncyvkWSC
wBzU6i9AYQzPN2PJlV7kmfgQnoQyNXe9Mrsa6gAcN/p/keUEYK0FpBB0W4wXwDPcN0cZ+90noNKn
uCKHUN5o+OsezGiWTUR+gICQ927CTb9ktp2XyWhI69mE4Fv4GXKGhJkYIbVS9CFVfO6IibHS9oWE
lO69PQwXhH4r8YphB4y/YNXi6369wTe6VXrS4HNNIK6HlJZ5/L3DmsdZdE/SRLO955CFtVbtRna0
igCHFrFH+Fx630zjoXA2zE7O0zPbLZc9nVPsswdhqCOHKpse1M6Qf3TXgz919fxUahNtxFHNVtJW
3chzC+H7Pv5fV9lKwB69sXsqOqh1XXLMHwXPGYWZk9KFnsXcw9THbWek4RZurV4WiUIk6J45s0Rv
GANvYjph7gaaw1UQAME92uGtJz1KE8MPHO6eVRK+2Jrfg9Hhjb+q5AgJeUF0hKuU955sCvNGEOfN
D28yqYsa+UV2zb4tEDH4ckXaFZC5DwgmNq48KdGXp4ItlC33ppHuU1nY+RnSn3HzxHys7X5/FQfE
TPJxznDb/xTVJ7uIp9rT44kN4tzjAkMHX0vd0gnJxEYWITfX2EV1Uljc1WMQ3sr6Wuu9q4VSt7ZP
5CncV40k0TZ3bjH56rlcP8PB7Q1zZ8KQjeRZkBFwFVeCUDD8QxmLHP/7jtFQmP8K0Fu3+7bTXXM6
mYh6ALae2qWnk+ZPt8/c9qpb/NupgfQ6BzaT15Ae6kRboCCIxSxRnfFb61/TAbiC2OtoMQw2+vil
WSmwel0bzfKKqSMNWa11u8W82LJcphWWkrQTGygBIZRMOU0952r7vHK99EXz6SqVKehajLelzRbf
pisFW15tjMNYyCqovMGbSrr90PM2GUTlu7ekwxJDwEH/W54smWWWXav+p/rgKljmkBb8adRObrcb
R5SIZRBXvDejKfraahPkvCBJEsz0AQ7PQZ7JZZQzCHcNxE7B0GPgTtwC3rES0sTtmtLzEV8/2ynY
noJPck7S3qzze/UlZ/7hPEY80ZbDdGWuKi85UTqNCUdWNRTc0DPmhqXyCOo+P5mdbvHEoNjrz3ID
TLK3EPRubz/32PJAzhBloyePx3+Ow5GeUR8mj9Zw0CK/BmrgKZ2RLvbDyQZU6ZeEraPP4WHK6it+
agIZK8tH8RLVl8muaIDC5YpCRF+EGDM0TuLK22oU5ETAUJq74psmT2TZmrXQ+quPw4UEdCWQUSx7
KjX8aD80uCxgvxVlBRlIoEgktY6V3NCrs3Y1nnNQlcIY8bC+VtIVnh1JrY9abRwLStGgLjM0Zzul
ss4msEqOKSbs8KCiz6t/lwfGccIX8ENQ1wxUtiTx7zjzW+vwkN5o0lZ6Id/7RmKlZIG+l+mlH7YN
9YKulTgtWE8sD+ruypYql7S/mo8iiCKKDO5uYSKzwsGTI0cWy420TVGRb0K1cfXXPoySwzsHC4JT
pK9wnhEBQyqkhSVtbXS85hl+o4UhhGyElHg5A7V0fTH77Cl/73HkLDz5T16uCpr+sUA859tv5UJ3
zsAuMMrCECCXNDDdXg6gB3bZ81cknCIOhBfN29nMMf1Bz9eX47vo2X2fwTK1nC8sIAeMkEIPfk7B
MusNxao1DdLd4N7iyrUJ9OeFIvB3WclZxvKIa2aS4L9X33Ayn0vlSwEzL2JYtIvusrdkRcX1OTjO
zd54C1yZJ6SHwQDsZadMZvSr/mDdHmiPS0X9TTTN1jDXOcF8gFhwig6UnCH4uyy3eBPy6yxR7jAm
S2GGwxevl1atlEBgDLjlVJM39YvsemWKHOduG79iSQjRn6tnhxXduIPGn8iBCgANKmL2yF1FshsS
lJHsyN4VYVVZISwQJRgW/T4aqRtqxqHYsFPeWZGgsfTe6L12glnwRyelGxYylRNlBpTFCsS/rTvs
9lpDoO8kf8wx4t/rGw4rAzM81vS8TP0FY/bshum0li2RN/PiIlyfWSOCKiwSXdREpg+ZxtOV+yUd
jsQWaxuH/G2ojklPIvW3JPsJYRooPoVEhAum/5JQ63nCs60j2QMOeXauOvGyfsOLOR9/o78wzS1S
FjdTy1Qi7hDY931DegFJp1xAI85eZns5qsew2JGITpl+Z3oe4kVqzlrdRAPpucM35myV5Ki+o2uw
vUIU1LWW/x0O0BMFayymQJHNMlL2kO1lyseU0PyFyqXcR9UgvXbttNH0rLmLemwvZgVJ8DjZzoQ4
q++zSAjuCccjgYvxBNjr6rJcA5Q7PMz8YgCYvEtyFQVfoDFflwJ7uJycO/iGaPJFfFxbMFN3TRuV
ZR44u89HCDLSAHyTbNDaPyEruofg7HagSGX//AI9gz/c8wVageTyJSDNm1KbLIzjrFVglxAxhNBa
DdLN/RHUM4ry0QtXWqe/AKZ7Kff4gt/cdDT8fDnry6IqGhHlLd1T75JGc2nZfK5rxa3y5x5AK3Sl
jWNejgS9VpRn8pXHbIIOmI2swcLyFQbQKyKbjbICY7xhoc2SbiqSIJqyHM0mSXSisDFv7zwBj2gx
KAv4xXUtmwdzoCIeGsAm897yG3wyCJrSJ7/AlLht+mVFIKmfBzMdOBgmTLaY7jP0cLPt8FVviGJh
Y8D0BEE0RRYT641ptSkAGTGErH7j+S9idMDWsXtsFx3dkPqXFxIFYp8FbIr/aC2x8X4WpS1askly
3kF/+M3twTfZiWw7Tgec9yqcVTJxZ/g9/VhUC4PHFQo0piitFA46w+nJOaW70ExVPxvQdxUA9paq
6o4owU5sQwpF6AoD1+9Un3HFdKxVHFp4x/sELJAVtHKrC+SnU0VPde3YPCxZBeKN04xgbcckbwk0
x4YsOin82arHlfc56NDckGHO9Ck/9Xn8Hlzq3hJ4M6nY1BZtQugm0UQ/8PrYd0GA07abLyg8gbEk
yPmIqKOEvmcs/0tvwUVGmOuJkfy73D7htbQzdGM7zNYjmHNwS9YnnmTJQ0+eFpdyJ0uEKb46Bvp7
snLzLd80Zesa7pSJ9/oIny4UY2EHHsQVYpu4VWsFht9pjbN6sOHi0XPZqPHA+YJPToD9dh1syp/+
wlRYk1iIF1blMQbkL3FE+aacQZStgA8+Tzy+Yy/XW64y1ZOaR0O1J5BQGkM224UBbfJkzuGDzvZp
oLvNcV5T8tOPRzlaTxEhWIkDp7cvHnIVeDpIj1YBxv3qwm3drudIcjI5ugldJ1uv+C300D/HjEhh
95fJ6KdzsjwvWDwokcfUGWW61XAL7dMpzEJrUGdkWO32UvCqA7sa2Py/Ng9dCEwyYLj2fhQao6S9
rwjay79p9nb+GqKlbfAlpFu2pklUMDUt3m0HezryilI9BU9+NRITdUCb5eKzCL4dAoE+h+X9PTeq
UYRfZ+acsimG2t543ztM4wAKMJDjaDnC4ByfzxTESF+OE/xTedYysfQOZEi+LvkuxgKEHkvd5kVW
Yjk0O7DTiucETywUps8tyn31TseiveoR1iOWIPIwS9U2+V1B/z7Z1tuQ1e5RtlokEBxT7Lzr92kU
pxANk4uGAudKMkVXGABEipwB28ZFToZ5QroRiNHzeu4I9jROuUrk5QU3Gh5yWy55lMJUFimWvb9S
2HHCXWpd7MczxISVtWZJFFCGNE/caImpOJtX7qzH3US36TsJtitkGLE3tYOqOswnTDyKH8tvGAkG
upjLpr09LuepkDrwN664QJz6nPrQDOoMfy2R4+ObScmK04E3bw+/X+W4eMrG+XzvZI3LDy6Dmoh0
3bKMQAsMSTaS06SSndoT5Rq+tCSOG7WBTNZEhrpb9y3cBqgi1heU2IIiJHDgm2gBrnIylNls6eaS
gkDn7UUhQWnKPVXZ9GAWoRMZJ86hSCVgXr5glspNK+vIBCD4Br8gorQXA7o0Kc/UNpPSlqT3o2sN
3a+fbAfS8ZJgI+Hs9rXg+iFO9j49fG4b+NtIyHCxdjUeZW0TLCdq+xuBqmsEA0uGCPcewqjlNCd2
5qrFoTXJvjGRr4/DWiKEKGg3CTNbncHD/j1KKHwAt7QFZJnHU0NX48N5gd1S5T6iYCGUD5Eaphac
wAqA507H8aMDklMZtJP/M6sAzq5PaI4lE56r17LKJ9h/rR4790p/40ZEOPhF6A40g+oCnwnn1qLC
XsT8XDqqHOaTpzcNv99UZFck2j+fccEZ9DOJxmQsDZForSWYccgWzTQ6wCEp5KyJxTw7y6bgkUWd
OdUjueD2aGBLWv1TJHLgUYTVcx9D/YR1ibZ3vPNqioqzQ2wkOqOnXaM0y7NhkhBMYzXeAqIT3UA6
udO/nFDzDg6EhoNN8sSH2O/Nj9Zi1WT5VCP1BCHlz3zUBvXvTpKcyvoVSH40B1blioR/HO4NNFIf
DC/9jxPX8EXyPvzYm8EOKgHeRaQUKmUkhnzqxOawZaTkheqsfGzTMthDqDc9du+KM1P5U8sebvD4
EG9nfrHdYZnpJ8TysXyWI1sjnTpi89s6SrjzCzrnOLQfpDAyOtS6ublQyMkjkjO3TXl5Z/w342Cu
y9vBgHJ4gy6MELGXhUHQa72mH+HHLkcbxzwTqAVsIb5UJbQaalKdJ8jwj6VdHEiX2hBzlgcwaVka
VOHYVClGq7CegKFbb+XSXP13p6b4XMFJZ/Yoanqmgdf2i4VJjrZ/CSofgFO7piLwe9IyAiyHHWLi
IXODmIltqyrYJD2s8mKe1xvnFKP3hh4FJKQ0K57aMYwFrtpANjKQNBwn8+5PIeGA+8XL8fY92ub0
dOyXVK6EHyqtPRcHCEaSSDdVclcugdE5MzsDD0kbD0u8NeUulJu6pAYX4vhRM+WdaceAKlNBzlGZ
narl5mz1wCu5bu8GRj9Z0JoJJuq3zqMZuSauHJ5Hy6mz1HyQFi7F8JC1Ingy4i7+Y7TtT3umJWa2
iFJJ0ZxQXr8wpFKz/QD1wUS1jlLpNnNgdwmLR+IjqRyIVsSSLWLECRqTur7+kFuMzHy7vxdHoMYq
JYFsGhAMncrZ0mTrcfwoNVjJnCJbTFMkBgo+TSHQO39SdTjBWYkJDX6QUZThJKfXVoReGXEhTeRI
LgG7RwJtSnuwo7VjlzYIdxz1jXcW7Jct9+IkiqfAMzEj2ueRyaXiSk/krA4cCOUqx1Pn4Pz/qfjI
apDIUd9Csz76kqIgXbx08SnpAFvIFBHVNG7VOvhacEWZSL3kJLp3qAtgqVGVaQhlzH5A6IC8mJzL
fY3RhzAscF3esjb+aLz/vpNs11uIlfczZ2wpP0Us1aO6JYKzOUANOz6kr2gj/IwvkYeZXY0C+WnN
ZpQzYCZ88JcoP8Z7uLAHFimtWNseE1rjud8S/PzcQ5Jzpzu9nEXVPH0CvPyG3nwK5/xp/UwjC167
aUO6feh1W0CaxuKgdiaA1IkuMg5pysjetjUy+eAngURn0HU13NVl+DWyTiYNJwUAryTDyCP1K/bV
xHs1OtzGJkDhom2crByakY+4+n3/DY0ELdzyGco1qB6967twAAfu6DYoOnHz/uaLy8GZza033/np
64hI8ZIPhwYjrQfmBkB4rmJ5F7m6POY+wUdrsyNPX+vnt2bzRSQI5NNV0hQfhBRL9rWBlRiiNIOM
1+TyrcouFaDHbP8G/AiEOcIeWfqApzAqhfoUEBLal2mKsRe1apK+zujrI32PJEE6FEnGS6I6HgkN
JrqGrgyYg/U4CgOPxPxkFeBMnElj7tZf0M/rW5h9dOJ980qaDr8jH+AoH/oTaPZrg90/uhtXaYaB
4JnMv/IVNIlPS12z+otITHVJw6Ts8rcwMs1j519GAZaWtujkzhUQLeHBj7J2RBvIwZZrMMhDYmEW
G3Wo1XEYgFvE2je63DxZA7N8j6PQ7+IzlvWPckbhv3Eb3BiTrjzp/0nL6Hqc79n98fR49v6WiW8G
n64pSRLerdwtZoo2unb/LfNDAMDb8IOMfk4LK+isZsaioU+sVJ23yjGdA0UjuNHGPScw+wWq3md3
aBiNaM/KzkbOvtsd/+XRjF3pizJxoyL1cemMBcdryxgjOj8d/MyqX/XcQLyWfqH80To+E5lxPaOb
M0H0WmZx0stabh0FE0c0STaLDrWTovrV4AOz+frvYPzjf77iXoFhFN4t3Ewe50ZbksjbLRoY4UTn
bj4z9SPc69XdiIUAQjZrKnKZmJSaB/QMSsBnzzy/476pH670UH3UMTGSo24jCyWjpvB9zB/zqVQL
9zI9WrUx0e9gP9bLweSgs+HBM80oYdpreeHPKujZ6rJAZtQZwUS/J+2FBB4OwQzsoYfrSLK/caR4
UJP84qgDerAefaZESE2T2WZjnugWwhjs7CuU3Sb9Qw4NbtUSClPfFtY4d/9pzQbJzIesmX4v+YYc
ShIxdZ2M3TGnyjngJNkmU4hr2dFvDpTnc9TKFr9DJdkll3nxbTJml7t8OR5gAwXvAvb9IMIAwVTV
/pCWETMiKSDmdX7vJLUjo+IPiXCuJzQ45ikUEbtB+fk+V4XWB7UNAe5e3Cj9jq4aKfomm/6G0DPK
4cF5rgiA9sTrP8WY1tIQqqbquxu6UU4JJpxP0qbXNGH3hrolYQRIhUFHVZesApvcEo05mb5zYOn5
BYZT/Dg/xwrCsD1wuBKFuMV06IxK48D0cT3YbTW47sxBKeNh92nYCMiaL3sMkHl8VdrH7hDNQS1k
zW+r9jUFQ9xbuc4dBYy9rDxJqR3/LL0ROvUoJBl/FUyIbZNy6odRslC8kGezy3jRPKokQt9BcDrt
EcpNF65fIvMQ/fsdBkekrxs9Njo2RsWfcc34FJKJ439ud9weSO/vPVAg76Rca8MOrhdOCM7uV0+8
nHrq0KiGA1WRZD7BimO5ReIkmxICmaxzgbgqVfRWcZ56r6LYTUj/aGbW1g+Dr/ZWmS1Jd/JUQGjD
54Flg7FOdZoVdl47fDJBBnyraj/nLHyOQcLh3Zhl7AiQopQunjhvXhWkzBkjdfmnzPJq+imqR/PZ
pLw6dgXkgPrvCoe+tCyq18LEqha3CZhAgjpch5R148AcvLTYqD1xSfHz9c3AbT3Qz8g4PiOgn4gz
yGA/pGGHgfbn4Bs4Gd3t6N+OQ+PrDLcNJqng4oiwwiTZO31CqRsqtZdVn9fhygjiLYq6QTntzc8x
1WrMeJEaPnMmjAzEEI3ldPsR7SiN3CR6uuft6K0wo2xutvM9W6HS+IiaPSDUu3Zd18/IP994lCDj
a6YG9RG91fxyq0nLTRXL+bftGgSkqUJDkuEry8qRiYq65qXjKPlslDNuZsIDBge/C/G5NVUI2beg
KAvbfpRXTOyILaWMjjDzuuTBJKP7zJkd1SmkjUMgEpB7WJyc9gqud4//xL8NdWxHPy+miQB9M4+9
bwOa7BJqg01Ut3tJa9diwCAh8/A5lUQMCR2+VH1nrFTXiIkWBsV0L46H8GrAe8xDDtZQ5hMVUWom
nwcFWsS+SBoaMt/iqCqjDV4q7slhds6iMfntp+rcFJnQoHhgJPrPXoiak3XLH6DZxznV0cBmGaEO
GfHXL20laQenczTEN4OOuef4KP/gMjrZ6S3QFqzVIPFspmotEYOQll0yUlA5+T/t3xbehOtd2tDF
v3FiXqRJ57CEeDJD3aK9BI2vwganp1G6ZbW8u1uXEmiwIDjkEWskvd4zt1l5hSIR8yeGgdSrFceX
Cny7Ng2zVxAJ4SowyG0NV6oLm6IgnZnbICZHTkvVbjwtoWwP+oHnSOmtUH6l6ZFRdI+lMbSjfn0A
AchSDz0qhf7uo8emYgJJyaRDpEedI+c0tI+Q86Xh/zRveuAvRGLasxMxfLa/hKwkBoUluOqwjGxa
vtgIMnHjWYwKgFlj/l9p39pmb+1TUAf49NkWyg6JKVv9hANMehgN9ay4jgUrdNTwu4lbpwRwGowZ
wwKNaDahHHFyVUXNtqM7J/Nzs+0DBRM8bN1MRDAYgSzL+AwjsuUNaV0jPmk9tLiI4oY7xK0fcvbY
AO6WAQfZjl432qFNEkAommwbfGrocR6mBkXxRapsEj3VziAbU3EFdsOto2DBGrPUh8W1cR5Q9pKL
ypVjtIkXRSPqkl/rqPwmtcin2uZlIShEyW58obSovJr4h8NKf2YSg1kuokEdndKx87xn3XRikmHy
E8vwTzw5SUHSm/Qmo3xBAB0eH2b3jap6N0hZfiG9aO2uzsksQr1uxLgvPQPn//JIrg5I5vlVpjSv
SQLaKZwEtXjcatGiC0Kwb394Je9jEKAE4xMxeoSvaP3WFJCWaPoD/VDCibmr4HJ69/Q/iv5vHF0c
YCEZrIDjX3e49GQgTu5aycTaNtPT9tpbUP3vQZib0GxkjvI0Oj1A3HW7vQPm2Rq3475PMQZSfU9p
xxqp43qH3SPOKDVjE2LyGx60ck7xfYY18DvM8BP8a0FNavnPWT2O0yP4zDAB48VBpyC4m0c4jUen
N8liAgtKsaHoTDxxhPO4Nwv78YLvpIXBl8ztjvcbpZbth/mPeAfg/HGrzNmM0TeCYN8+egLbPM6B
tm83SsYOmWAOlT0JoAgMzLBMcUVrSDJj9rTqbQVRa4q3AFy13KakblSaOng8xE7Eo1RYbQG4fEOW
eqvP8gYKP+RoKZOALVmBHM929FTRFABE8ARuspZ8IgA7TTbUfO8YlC2nMVYaSJzUdUMwPLTDY1iF
EmuWBh4+TAT0kVau75rGJGaRyNfVSaUcsOuYScW3o/EVTl4g3rYM9WPTGDVREpb/kryXCxrV4v2j
fsoeg4EgM9yZOfsDUki1LhSEgO2nwF6LXUsyqHOBzLOyHdQo/wY5huoFZC1oyTQ46ian40+2RGSA
F5c/iSYWrjydOgg6YnIkCqj6NFw6ypxx5UWH1lPPB3+Zm/gJFjH5qaiSVVvidC3yoYySy/xsCONq
F+F/JMxfihwtWTzbeV04FkhWOrET0toN13ombiiORXH5XVk4DKTg2Q62A7VY4LTlhVsTW7FPHFLM
cIJIcZF+MvpsNw6A4wVsfei7WxnXJyXr3EsM7qfriFRL+f5th9uh8CsBDVPchvxSbQ0tJm2dldNK
K8wQHTyKDSquk8AiWmTWlrjvrJZsWCo4h0KMyPDG5wlkUNDuIAqyejvpP+h3EjITxZMWJ7f+MVI+
zLTmpJEFPhmPzta+YSB6Kg1qILWYSWHolgkC0tmvE417GfAbN46RN+MheoLZET20f5GD62lc6MUY
xv4eEsQHnlgvQqX5IPBuXje9P5AjH+IoDAL8RGVyq6xcLpMLLZn7kZ0I0dEQwscx8VOoSsAd9KCd
IePSQvRBzJTLx/JsOah+z77E6nYL3zEsf3qyhFycMeWXpKQu4DpIyltVo/D4kc+2pabpEbAZjqd6
14OwfeS2eeQ+AN5TY/ImWbSKUezyNUsvHGGXKWObtqjSDt/ZS+naRvmcyOABeJnfN30pxiTNs945
yQKOMb8TeyzPmZSqKTF3LjAue/96yhoqZIxW1xZS0vP0g9fe+vUB7p4SVD30c91l6inMfUURRQQM
mxdLnmf0dApi5vrG/dyeK84R5g9mbPVphV7x3A6tZOkxD7h32GVu4PASzCT2vGFG2N8Q6rEJh34P
EFgXpxDjbT1QOiZPOV05ACnCuU81azuZ74ODYKE+TYMMZxX9YIwcQafXAGo1772y6j6AmRcBWCEp
+Z32JD8Dgyi4/NZOsEUfFvkV7v5c1s+mDKDls6qrQ/VljwUwhW3YgIdIHcXbE34n0YT5qsTokJmS
uBKTzfUiilvc44p6G39b72QcH0PFTcCmOHcvJDYC+4C4hDW7VqYuX4u0TFlf7xcE0CxgwejhWA8w
CRalY4jK9pkdN3uSlpjWbFnfESCkLJcIA0RSE7gkjkLfVM0fKaWZH2ppg5H7kLKMJBnkf1qY1Dmr
uxNsa7GOlUY3eBHscwvp+0UC8RGiR730xvhZ/5HqkKIaZvIrX9/qWYsHS/IYN8HNYJGd2n3WVO+G
Rvdru+26j3dcZZCWdTViTgheotm9QGpHRcvScWlZ5mxVXY4j6zr4by/Xd/M7R2nf0Zy3RWuwVwAP
KCdGqaPC51FOUAuwVSV2D9zLBaIn4PnlQpeoEvkgL4HqMJUhB9WquzuimEvNE2PnVC2C+Y7i6S3j
5zPZWSmPKMxtvnqrO4GIl5ovZTVGHdRN2kR8GNBqoNNSzBjDS47rbcWEqNpaK2fHqBrTsXCID/w3
2zBhBmJi0makvN28TmqSDz8g7hsvnCnc136snq1oruJTEsajtXRJ8O8S83P45YqZejAIPV8udNXC
AtVvEptHlnTPoWx75ntocgExFWcLmRJw18G1HmeTppN+m3+ce6OuFEHD5V//Dmi1vskMommwfzBh
dfeEv4PXBeVp290OmrMFPd/B+6v2wFA18VLQh6KhnNGY3ZOjkLBDSjsjkJxA+yloyQ9aGugOlbGW
RvVQ+/Ipg0v7UeHSLnm77pppQNmQW4dCJ59mLPlenWiEuwhkOpZRuqwVSPK7b+LfnLkVuDqO9K5N
/HV3d3GNKAsqsIfbiMjKJvz6xykDjJTGyuDj0kLjMXLSbvNUxRG5B6867NfGIsIyMmBimmFEyZZb
3A0DQw1st7qH8RG4MAK6+BWDWYu42L495YAlftJou3eRB5e8x6NRvavUMSkTeZU16dXC5mWp/JaZ
xgIzlTKyTi0UEawLciuuxBdZUt7KiIyGSkyGnsFNVZYPWHJtNbG37kzHoIF29vJQLw+Y6NPUeOry
s4fRWG9KAmcb2AUQ/sVTIWBRaiSpVaDhtx4s0d1IhY3q5+T0Z3j4KrS7knTYkaxGGaTvuIz7rcuO
vqA/vLxzYSUQ18DAinWLDSZPnjyMVrkGPROyuI+g31/b4ycX0qSkXhluPa2o+muQgj02Z2+Ay4NE
czpnDorXod0v2tQVS/KPjZ41fkspLvi65UucNSlqSj6PpUY0M59ZjR/bAxagaonho+ZSXdCfAx4i
oAGHfXqIuGlbzU7MQ2O2DXXl4H/QKMUZaUhO569DOkfAzOqC0zKFPQHsjJTmSiV5Se79MRJM+frO
Z0NlDcKIoBBuPgfgXMjTqxDrRUTlrJOMnRnBmCGI5wqajY+u3tJTDzLHRthT1E9oDR3B9zs65JBf
UZ9wttTIAQAmU4JroYVjfxh0SnuQtjLkIEFfVmFAvHtaD7Nf4xFrFbGvziJpCGNirQrL0wwEj5cZ
T79kMsTKQekPsz4KKBcm1T9kkWkJWuzk7x6A3cHDc4TMJ7TFi2Jc2W2OzbifpOhrdLtxysx4t5G6
9ghCWevGHkQKPKJKoyGaiwL0Ad2t0Pd5nNjAIb40lCnecv2mLIWuE6VJKUg/UZFxfiOT+TrU0IOb
146lLBB/C3oU1WZJO6+Ia9BnuCUiQmvxHgFlSOf/RB42uzoMBdWM9pUEDD+buN5JHhnMs/T1/Akv
Z9L3g37mHxZC2tFqHpmZCSklf6eviO0v/E/p7D9vXfbnVEdFAJ26KkqljzJRaKypv1i+LJ5PXg3E
ekuHeORuajmgtgS72YRIrQcafWyYaT5euWbzgPWWsDbPLxM3AFd3GskEDUwur1MB85OZcswzuIHc
lRQPzryVGeA+dDEB+96qoyxG2bWpNG8wtBcz9KMh4/yvBlcwNk/hqhdmC7NMfMTgoT1HHgO+a9GH
72d9NB8ONO2Tre3QRCzbC/CD0kGv4QHMRh6TbTGrJqxnvTTWJ3O6qU7eHkQBQ0ub6eL6H6EXttiM
Rys4SP9rl71xTmh8p6G4XMlJb+iHMScZwbC47j5AzUi8hYoNbWIar2pPv4c/R/KbwyxN3m6soAdZ
jY2xlr18zTcnj8q5B+WQn2/8qD2j/GH5xRPD9DIhqB8rC5fcpc54+11Cc6ytFsxXsk70qqTkX58Z
KVC7R27Bd6pl6D+Y8vecFUd7ad67pqnBk+/FKDXN6qnY780OQAS2woKr/auw5h8K9uo4PYcP5J+U
9sClW5Ll6/LwD+nWRqGO+/mY3tImuDjLRm+EHqDRxP2KHwF+KuYPFK0JnKLh2d95RFVLPRoWNALB
m+jTcX5kc2BwagHxp7WLNuYLaLQo8eSzU1YlYrQiMcj1cGvwFys9mbgEHkbOz+tdpv2iiFBgpmua
FFeXb8I38JRj2tyQqkjiBEMZgg/Y6I7AS5rrP0qGCBy1eflAGw9dVEQwhCQr4xOWOummDzGHQz+f
TuOBMhs83c1SvyJIs5kY7+Ih5632Ds8Ss5WlK95084hrj/AMhdF32cpX/E37UrJfgDzbvhQKCkhP
Mtxxyer9qnvTditSd+55WDt4S5hpTJHSHKo9JxzhDh1p8uv2ehwiQPkTNC1lDJgnlqeWBA/beePA
lygmW4mbjBYaeinqKCwRyNKEkynMtlh/s1nXXxF9dRVtuK61zuOLK40JjGd1V1nDnU/j5nyqjS+P
zAXo4cGmM7DnBrtVOyHppncgT8ap9hGQEx2BsnDjV0/uzNxSY6PSQR5OnIRHBJvMi5DxwirhF5t2
LGyHZ1W8XKVLlmN/d3TUeiRv0kkVRVFpp0EuIFuHBVGZqxQrxJROVQVNWbm5gWFeFg9m18eQX+1t
r+6wON6zoZc90QjWrOL0dj9unMmfmblErWNtWR8QDf87Dpx9kQx7FUdsdcj9HRpHswtvspZTwk7T
dhRxzEUTo8152cF6BEN7/skmYfGBKjyl2U7cfQIqfQo6s+M+6DU0gmdY9rNwiwPdSa57VmAajFe9
3z9m/1B9l+3f4UligIDxcdoHWv30Gh7Pmz1QW2Iony9gIklZ+XpHb20TV4uSkLAVbEucFf6MBOJF
xv1NqQRKNK16y69pl97ZEmwxYptAurYet5YNVhM0hf1tUvkgyFffTFStLmFbyvh+pkEYENYFqhaK
i1sQ0itZoxKgL+s/H4Qew30Ok25iDNJ/nDJHUVwFktfYy0REjW87zJ8qsgBRGo28ZEQVx9RRF+fo
CbVVS7q+ZBJthpiifmtEqcElZkS6Fzs0bzWnLjIixw4Sk1ErJr5U+mn1eRyqDGGa2tCT9Uuv7tin
pFs1ow7BBr+vMucJX4Qgj5EjWX15i8MHjlLafiFBERF+DzHn/7a6CpIChsjTRZ/QzhDM+3e7QeSD
L2jrCEnmab8dbJTYEakaqzydzWPZl1PqUZoinLo0tNtgyZ8ltZwhFhI+lSJQ6CAzPxy7VfAbwaMY
LM7LdTUNm5LTvHgvON02V5ds8qnQiPZV5PaUpn3cQROWsa0TFBOdqwkaHzv2Gt5eZIgqPGGemRYQ
lAqjd7S/bd0hyuySvEN2WthnEahVL+tP0lOUlMgfXBhNgbJ1vOd357sMyJIrjetW1KCJOMff8Iuh
pI0YQUVMWoYtMJEdhnN059+JiU0FxxdricsB6FdHO1Omn469uXervbNYoTc1y1NDaE9e/YAmwm6h
eCu90oviM5Ec2zUpBvBkDJQHey5LnSWw+dcvHjwe/lcRN9Vo9uBDGl5U7rV+NHa9ZCRqFmmhizqX
/I4OPogmrUmyBXYeZD4a2JLbIAw07wrLPR0AL31BLgT3duGkcjjbf0mkJsg2y5XmG4+B4SEePEUL
8w6jbdrZJ+COe0pXHE78RbocxOSEAzKZx/cmQ7Ey70Rwat53yZXA1aDNMr1NHx6VYKPhrRA9lGHB
eh3BahBO2Pb56W8Lv45SOJfIEZdC30+f191Szm7XOch9i6PoDIN8Q8bUOC6vEGH6h44VbkUrM4Ff
6jfAUaEPGEPix4pCudVeXDOYb5WUZ3vtjif6ZIowqYJLfIzedeXjcB5Ob9UTdROxqgcO7lAc7NFJ
9+icwNVKPqczPpcctMT78q2I7H1vVVNpmaSfRsP7fIxTnRmT+HVJf9yr5GuYQqCsx0yX4athpnZM
LdZOyXClDdAdI+g8p/iPwAkWwIl1V1Oxzg+TuXTq6lqjjzs+HsQCTRKUDyeRMTaK+qH01Es+rUB6
Ptr+pz/BqmGS2iPiFSeBcbCVHJSRodJOBx1k0/4FzZZsdcekuL8VkT8aCggBoVzDfjnkKbW7tYFI
QvMYP4wGwfryZU1qdEsxzVDCVX/YnhiKkJwNdXAUbxFJCErDHr62/7xG7J5X1Z2F65gKXyPhOkSr
WLA/XUZww/UH8fucxwUlLrsrizwaiomp/j9ULVy8mmAQwmqDm/PYvVUU5AnL/3r0ZYwSaGbQz+W7
9bq6yk8OHt5uRU+Zz3YIrmZxPm2NMEs1gOAJ1YaSo7zjLtrIaAHkYu7IyuTelVDX5bZK+WkLld8d
TFCZxv+j7TmjbUotUeHxEjrg7xuTcN8QelwPZ3cTYy9aVrkRxZJAhWmRVsl3mOd3rUz3lzllcZmH
is50kczg1Wo8cdnP5Ch+XLS6DYdYQ5GCS6YmzU4dMZFGvTNCggZr93CBV03mh5xtXb4uoXNwc4yu
bEnYOr9TshabseA56DaLZWP+48PBuNf/kwKnfXiGQXb2jG29M3PPbL6H0L6An2GCYUDeQb24ZNqu
V2Po0eRsyWpt6exnXu+E46bH0fX3uO/uWITovpKq7AWfp3ReJsodRPLNAPdpwVXLoh0aPkY0D+nE
p9e6+Sc22AGRt+L4stW2yCk+UdABntDba4ZKAgAyR1427MKdbJP6ldF7fqtwc5f5SsV8TbEcf5TY
zKMzkXMGfBD4Ai/WlqHIBiXuM45xWZTyLhDH0qD2P+GufWaEK4wrpOEqVoHBPmSccX6FiJIEWQiY
CdPSd9X4jDLc0WgR9BbbpqDM+mcLiJg3LCkkVImGUxb8+cvvYxhbeLwzvsUXZYtOFcLYgZF4RBMg
CsT/HO3TvU/x+v97Ag8R8tT716yKNAAuvCQgz4sDA28uSPf6PH05GhDcl83PHZRXaGS3ODybXLXh
ubm1aVn9OKFRtsPAU0d6Joc3qGoJ8iIAzRQ87rbTOBgN7NJv9/YFpT1CygUjCDGwBkk61dLtyKwS
es4dlX1hKGq8px88eFBKlAcWZ4FMhBKIea3jTjX860wYk9woCSsHzM1vRh7u0oAzZYZtWFU1BJhw
bwuhegHetxFL7NPqbX7FdHFMeNc5QPZM5geDYFq7i1WsFmNrH1V9r8QNZq+xAXlj0btOuMhL8iQf
/L7SaObDU6eKN1Ky+Bo39M1X/1zpOvqG/jy5ZXzsJYIc2SM8dy3nFlfjVzSmsdaxoSn7cHCfal6V
hoRdWEIoowHvtHHkm+E4aJKD8aOaQ1919Gckd+Z5FQBJr9UJSu4aJt1048faBm+fvojIC7rwklEK
6TjH1oMpSi/OUK/Gcz78OzPDgNXzyweGm1mXpE6hNBp9HSe8GujbgJ36MtSmQBAH/BiExb2eJgQw
fKhy1C/oiBu3XNIsa6b4TE47lC6NK/QzEHXerw/i/r6wxBA57JSZALEMLUtO+Ex1DHrD15D+mOJZ
f7p9aj1PCW0scxRwZZmxEI+DO86flP92AQzLzNGcc6oEkiYsGYWoNFdMFmpkDYuGGVP3fmXQiyBD
8WptF5eUudLGxX/eVFmaat5PYRBpoaWSAVplBpVVaIteyMY5urDr9uZYk2Hh9jFHnAzADD0XbmuW
0NoSXHnJSa2pjHL2OraR5fHiWGRXvroXkXRut6XVAGO3k4LtHLv9YtemdzzQxphljZObV8XIwvW0
4y77fQ67ptsGh8eKTjkHbrU6iZtlASgt86gRg3ypzAv3hKuhNzlCoeJmt1AIOLl1zRNl9T2kC65V
LiJv+FndAcKG10LX5b2RWZciR3FMZIIfJsjOWPcAwOk8INShL35u4PGv10viHVAr/wnoJbUydDPk
1/cc1jfxTHo429SA48lwB36ao34WfKQgCR+FPEPohJ+Ez/vPlfq0/YsUx6Hz4kzFcyRbdJNl+rUI
MF+nXYCbb2umB4XC7tDpTOpIHsMlBISZj/efF6U/SwXjl2sDHkH2CMBiWxnXEpu7fB8z5DU3kXVf
AHN7fWc16ZsQuVNsaTZnMGpL/0LMiIVwQKsg/4zd8TD/oyxgEmPMKkXUtNraH2cT0SyUGRbE3Qzv
PWBx55PclujhhETpX6QpQ3lP2hK/Vy6jAAXNsJ6Q2CLJbnFbpFgy8uX0Ha1DFYBcACvqXYjx+nra
KdPW6owhLRG0Q0ohGXxhBB+V257mvjQRodRzeur840OQ8r7DZxAqdVyDtSuYFhBvh6IyLI4KVk56
Ps1m/MF51FS39qoh/FkSGv4fIlV24eWLJg/GPHYcw85dRqXwonOurTxN11QnCkJl4uamBRyobki9
SceZEgcm3xF5VtwIZfo8v9XODNBKWXHvGcdNJtjXLIpkOIzoOHzx5Y1WnDNbs7HhO0Kuv+bPuwYX
Qsb92EjT2JXrOoynwLQ2abgy49/ecuZoBirJKfmsBxfwuKb3IhOyIiH5ypLK1okZdTkONlTL8B4e
50LtV79FGwQmOicNkk2R42I46NMuvLAdf5HogHHGQwcZe74cM8V1jB9EVGKtIR7mXWbxvMW14zCx
5nf5RD8Ye3T2ZsFN36xfLg0qqWpXcrWjoa0bH/zvUuNyRN/fhiGJ+iCZEUgE6cCbYa88FAgIOyek
M6TpHCpcjj78Fqdn7xyWhh4kcCtAFutp7igOrP/nGIVsPxn2LP0/U8DauqXHST73+hcnmcBUZpKt
ZmJSUv4RZf3TE+pufpiixwEiboOJ8E56aQxMJqJGWVebTb6Xe2ze5ZmXe2jeyoP3d5AWjiyQ07Cz
AFiSOcYQuOM+CFWSL4pahPuzfzT16W/O5yqNmHozpfZyhYB4m+6qHLDC7ngWw22mgz5dvEboyY+/
gSCfCqhJTLrVMHmxJ0AFX7wrCozk+hMC+FhPdvshou78bRjiZAIDyzpaBTa9a7lSOEpJaurh8+qz
VZJ3/iwsr4KOQDOFz9Rt0Jn5k1Y9mgy9vF5lzbAg+quDzkAId+3K+2mZxv7fErSvByP9OqEPO/aY
ZWpeVlughPIlcPJXVuCDywIl0lYRkFYhvNREUul2j65qVOQEf0MHugbLPOA4G7DVESOXHp7mH8v0
D0DEL9WkxpuY4mwLqYvUcnvhjK95p8VXgxp5rAIyLG/yoVNeYym6OGI1HruOXUQq1ZPl0NK6rL9q
viOWQCigePSqImvS0v0hGkMuaK0CiD401kgSEXp10p7gcir1oWIDxvDqALFGszUC7Yf4g6+LLYXy
ujs+hp5ec4v0pv9Y9qa3FxYbKPuEzr1cDwiUd3eP/zFrtKr9EXvVaE83GU453xjXGwur6akLqpJ5
f+9xnVBSI7R/NSOHB6SUckTQDypCwWaXQkavosW+ETtlhmSQlXMJYmorktGgl7p+0urm/UaS57+l
TU2MTeSzsIjyWG5knmUOQ7FND6t8Qv0laTCDkRdbF4aze8chSqBKuMJt9DbID8lqGl4zR6xV6bOP
N08YH4/R9+aDhLLxgI0zewffpF8gu6p6rNSprQhMSlIGN2yQ8OeZc6AVm4FcV1UNxUx8Q87lW1EE
+qJAP5Gy0VKQZsAqos0CFUepFNCSTQo1FTGwja7++tdh3NVOjDd6/kpyS86IBA8ZdoGAXnqzjHcL
PJesFO4FSzT25g4Ge07HWGI3aXIaxaXIOixKbrElvMHaOPANHjnkYXa+KzIXl7dnhafELEbCVxWi
bzVNPdDKp1kLd1yrDs5l9LC+0KKKoAn9j/zyPTQ1fFLPH19B0k10b+mUP63YAUy9CsYjyZKtI6jV
8xb3fnNbaSQpmqFaDmn8Kols4o7Sf/W4lIT7Emu3lbDoMDDjDpGZLuT0ktVHnSqD8Gwu9VysIlRb
BeSax9AIF7guDL1LOMr5k+wkRmfvf6VgVmYk3Vy6SZVUdPmiULWS+VxqOfHnGkwu5K9TnXlH1Is5
eVz1hpwKxmyTgfn2gX1vDW7DmeY88pZK6NCZ2UJRAYx1PwVQ6iwP6mqrEr3kCpcGp7YX4r749yEy
dvtGwZ39BdBtJMTK19mySB084nw4pRYTm2rr0ng85sJEHXIxuiD3wMkeIwTLM4Nq1vMXVwVOhC38
KuTjpI/gtxvSgLYcMgr2gVj4L7aIWCI4oJorzj5nr0fyvgm/lemvHsEZuziPWnZEbKziLY5tut+c
szdku8Fo1X9kuiAaRMwhVlgaisblStRPakUGCnuzaBCDjNCW6t/67FUY8ZTQqbIf2McHvfunen3O
TYoV04CdUq7qc2KCFRtYq18+YC2maKkHJPCtrX3GbLzJh9bQ2iohB+fTYLJRhfBGT3NbBDCYjNBi
xsZf2LM/gMUb6v5juR9MC4OjDFARSKaNAN4uhX2PiLwpCRWrV1cVzeA+rtYm/VOFbGiwrt4I17Ym
6rUsgnT/0Ad06K6GhCLmdHWerdm1pQdre+AQRdDhMPzM3hh0+wpaBo9ov0J9xFEgg4qKC0cJgY6u
Exe3O0CYRvhh0or7DSGEgAj8etYChl+b0eD3r723ncaOEE600HS0+aqJ0jXEfWQ7k3TbFcb36NK6
5a2p1vbHEAcbkLhGqjJIyp+A+wcE2PYTkn0oq2yMn/9rg02DR1f6NF9Md9QKdjIKL2vReCcS4ChO
XXzElfI5U8Ra55wkLF4+u8M4QeKBCT2swey7qxsniw86LofmnxG1rl+ENkoz3QM9VdV8AsnzMcYK
ZEMsy7RRvbNzqxxjjWohm19vNAIyPvWYiAABoNhoM54ykIE+l+2/luYVPZeO1l/gE3vCfzz4FYkT
gbseskhAZRJuJ13/l+wxdXduAoTOj/uBncnkMwuVDxLD2oB6AaNpBRewZzlNp9kgIs6cd9I76L2j
ZmJeJLZs7nMQTSdTemWlIbgp1QSELETTTUCKenicWcKbnsrchRT7LVOiqrcJl/juev0Rx68gx4AY
9S5KMnxhlxaPG3FuMbgMCwz4AIQ0yzm8/ar+5i5h26mq2VNqEWLZD3sTqQn4F0cHRX/gv1YbqHLb
PWbgtwHMoZo8K8wQzclw+0Vj0e0TwM+MPSnuxrToyM+g74letENG2vedv/Z3KnuXUjZZNHPJ6N5n
HWjlCnXLOIEmRe59/tEhO3k3vFK5/DtqqquDRxrqNacKepEyXWmmLlcLiWUYrO93IeiCiZIiicO5
kIp1DlSxDmnyUXDAgRii0tNjjP4FH6eAZx0cBrlnLox2cgArFnvzLXb3zo2Z2twwaaGDjJv+xln1
PxQqcNOwVM6AZmHWovjaYm5XCUkn7lHJiJCsZC9wncD3RqKHTEJg9lbqR7MTVJ5HpoTG9seSFsLg
31xg7+lgk7Em5+tWMnZ9bBtGiGd43ALRa1WMWyeEwcX+HAkWDSZMfdhj3i1xS6jfm4IyzfH9cdSw
JoN7yi5GP4FMkdQP1xGFK57VIjnXkQiMuE2AQQLtpd6xr2SrJ5AF5RYWu0MuVr5pHIAECoIMD4po
5AxnV7RW5iwNjfDNEjI/HBzCzmFoPyQbXD9C7AkDMjY1eoRKa/Qilumt90zqunCF3G+QWDgqlP3k
glUryJoyQn50RaRw1m9IWrkiHvepe5QasQNfwvJi0IaujJ9Z0FiXza1BGw/3u4mVAvYBNaPybdhD
sVl/y2VjsB9kO9DCV2iZyYSWWdCBfZYiYGL2t3UAZKGa7/d41ijBXV26+YnzdBmi0xUgqtqVgTwK
nKBvNfawVGqjdN+fIXO4D1megrEpqxLQH+fkiyNELPsN6n9zihtIjW9MTn7ZxyLX4r1Azz3sqBAG
JfZnNfPjsi8IKC9K1+iCRxTAv5hE99xJPc30VhY5IvRuNLvTCaMZeNj93Ak6RWNF24TBFoE8L4l1
Eo9X9vs00anoyPQngvfCLSMw+hk5aljiTXDLa4jStFOVtE/Vj7j2i+bYRtnkJTYa3Vjda1XALkCh
49NZTLyUwkAaPSjpMEyTixJ4h3DJeITYUKorUbPg05YtzghXm9rL1lTDhqE1BZqFJ6b+SLbNbNSi
syvGz7GdWizyQFShe5YsFyITwXtprqKb4mwakhep/mQmNj3YMIbtXlH4HVOOvfcMhwaReYQpIuMn
7dQZSeK9TbNVBeHchXIQVHqJ3h+OAujBrzWcg7qOWqz9fCeffKkWtb6ZuEphbt2dUFad5dx5GBE4
rvTiY/DS/KfRy5k96/PLFLhrApvTlily28niVK+bYOn3948MFsBprVUk/eYGrRQajT1ZhHfkZYYw
mbzb3mynfDNWc6AuvIHCP5qoh0mhl19LCt15eEhrJMBIPKFkW+ZKLeQ4Y//P4TUZIkhm8UVzhYTW
SJc2RmTcnB25vXzYbyg1HghbBFrWnIuEbpzUNtCJ9rAsAMCbHwv90ltMJrQdjItwIKwfqNBbdzwT
IDU98Nk/GhZmPh+4IFIHWuZYJ86lQNCmNVJqsIpxMfUKT8fvJ9fh1Nf0wp4EBypNS0kpVD49t6DR
JpDrCKrlOFODJN23hAy2HnGoX/hhBkiAHXneeEoDN+mVAU4O6400MmOXAS6wD1MPL5lvDVPv/DEk
miCaVW1CZHhJvxcD/KmPyBFmj8yin4crt6M6GuPUvmC8+TY3JQeIB7q2Af6mYgjCUMdEg9oKnoJI
YJUA1MYVeA9n0uRcLYdlSyVZvZ/uta6hUGb4GB9l9CBFkgVFTHLqeL98TPlWVxkQVmzhl8yv1bFO
d5CgPSYxn0xji+I+uVIqvU1EQS3VFbOMMv/gTxhzQ8qgE5ixrZY6BiqTvjMas1OX9LVm3bqSpr33
JrULUevM5v/1ntbxqx7fUUT2/KujYZW8+DSa8dYnh/rMYzFw0VFUnYfgMpqMcxcsxIjVx7lxtKhL
n6fPEBhXn5A9vwsKez1v4ds07gyDvfqf1ip9kTFsXvzeP4ynrOT+dM76lcWUQ2UDcy+r3ZNZAqo/
J17v5SR2PTizufpokYDO86yRKJv6zbTdKZqz+2sx1O9yXdXdP506S4JJyvwA7i3FCos6E7I4wbrq
EM6qpCAk19r/uILYiwJKULvRBD/LBkNhx33xCtUJx3znQAsWHYM1RcPurBcKDkgSPRlznbjOWqUf
A/hzivbubZFauoHw9mfZtV1s5JQiA02uAl0D8thVqWv4US1DzVk66/eo0KqPvG8v/L89ouZDcRFq
/VO2m1GXRcZKlEWhvKIDgIKbLMqvMoynG7j+XvDazZWAgDqAUWax2CWreZ1N9mYYnMWnrea+ZNKa
RTQyloEmUjy6uqUjBRYyv6kidI30wBDO+7d7V9igAEEtZHkBH9/fIE92XoTJMAFWx3X96D+RXzim
2PuDtSu1iqaAshuDWohfX/AuHatVCrRqfIgJY9bEpTNn8vEMl0Z4I3Gtld94wab2Bm3liSeJ8Q0x
JLMLKEeWk1K4ocS3k52ldeooYMUeIX8SgU1agCoQYWno3x1oat2MH4yvW+bdo+59HDWYdFkDe5Fg
rU6VxEcpyqt49yOThK+BCjrjKh7P63tmb1+aa3mOBw/ZIG4FuxK3oh0R1m7byv5SaCNIClrrQmOt
/3WjurjHm0x7QSo863Q8DFZDZaVelbs/w6WU00HggV4SqNVs8mgAYcN7yMCnS1pOPfZ+9ZK+Iqt8
Dsk0jTs/tSQnXPGfb6m1Bfwa/LABBQ0+WseXXYeQpLDgSh6QV6x59qx3ikK2JOCp85zZM8bEqOoj
HYwZ7EemWbxyw+l+ScnF7KTkj0HT7izWcvMaMvzuSjhUMxMaNZIAWr/R56vOhBxO+OaBVPohuff+
wVKLTq4UPbTAw72ONrcn3NpfABfYg4flemt40r7wMleXE9OPz6ZlA6akiXtsYht2nnnc6mYVeSIM
e1UgrSGRoCiH/Gxf/XWhlh9wjfPrFMUJAqqRjgGrcXNvfTWuP7B8hiUfrqPxmlOgj0LEAqPWd9dW
Skogx4aj16TArmFXmcMO4c+kmNPf+hcoNal6FV9dL2AiV9ILTpdezFsBKEpSXB1hzbDwvm0//GEP
+VwcgR8hdPwoPX1mtXBTCsquSLiKMu7/e3NqnD4a5kE+09DV1a2wLKM1MuiBCKuRgIATFKNM5hmI
ZaXFyIetiFzTIYOe/w30Z6goAGCh/KCooh1aXVig9xLIpP/0ee82+r/HL0TqUb8uQbTd4AdUqbfO
uK9XYwp+VXRfwPgladjY2q3aiakZt7iEFy+q2jWM8O+LJl8RdHhpAjWC8+X6YYstZn2fPWB1Z0qG
8Gy8wS6brzAnyQAQtOR13RNY6rcQItIei2+va9Ydbk/7Ch1crvJViUTcfu8SZcr7wXaF8M392jBl
ITP8Gpw4xZj2LhHb1Wbfr86wyz9sOT9hRh/6BUBvhIFfgXftzeqSbJh5ytSNVPJyl4C6GJuIWGLv
VKEyqdDe2QqG2PzaslcdktlZl1Gd2AWujMOGRKCt9/fbRANi3UdEzDWjBP70aTdsTgTJ7aG593bB
9dpiyDsYM/Q2TEkYIencgcw9Gndbeypet+x20EJeSRT3IrntjLBfntLNBKa3YpeeqH8VDf3ZC3/U
3a3jzFUCLGGfz0UcCuILQz8mLV3y+Pv44psPLlPFQN1ch8Vum5uZiiEFWSqBY/ZxlrlWBJ9ejFqC
+ct48fEjhYiJsRHmpHK1/2xs0cSM2aIOhiN9gJnzxn2X5R08SNLi5DGVeShIDYnsY6HVY3iU0SVW
GpfQH/HPg0W0uGwkU6QvZh8JuC7CVW7o7mQdH8hf54RvDXZCRaeqvLp3h5PehUAWU4U6ItRH6euQ
CQMraiSIV0OEl+1WqRW/pcFZ1XKrJPcmzRtQJusSvXIp7l4zLFi2KKbyCucjfSUhaZjCha+mYWHg
ZNcqDik+T3N//K1DWh+lv6zeq9+8AENvxwok1nKmfL82npxZ1S7R+923GPOXYDVmfi8GH3j17KJ3
yoyJvcj7K+S7rin+8oOyUeJbaxv/6WxL9Y1maC0wqzYBVMt7PQnfqFt5tHwDKFIkiTS0461Vwreu
MQTcjH7lJWtxucx5IHFmcP8D5+dBwFvGCtUVq6LsbxJqsFa34EaxNKAzjuwrJYK/b+5K2hOJYVqU
Rz+FqB6CW+iIuJen41mjsqEvnIBtHXF4hpFGT9M83Jwb4ZD/M27WvNYVSAlXNOeUv8I4BMXukw/8
tSSzFrJ8TPeHzaq1L/JomxG/Z5x2rFeOCi8iRKJzTdp8Z7DnSj5gTzbqRsIUEzQ7SVmvpeg5tLMi
sFe1sLTQzuOyP8jfQqc8KSwVntrSTgY+/z9LIs+MI9LrkfQsEEXDm0fbX38Q07bjlqKB+v5uy5zA
Ns6FeHktJKwHkOJbYf2baoAHJBusJSHZsWl0ZbqhTWGH5C3F68ONsTNTEIgHT29JvV1KMMaCRzKB
Cov1T6HotnQdSxJ8NkJ+R3Lbupsyn2j6vbVqsMDHkPNz8Xq3rTDvUSTjgYmYbPR77Q5cEN/CVu0/
FLXoSAb+xuFCtzgLWQULk3ci3eOCrEeMSyfxgzz0w2a1gFCxt4/+aLRgmUzUl9LnaQrRc94guPun
QbsF4fltDjVtcia2kvJp5DUeh01Au+yRtrq67ANmGRjkSuNLmhHvIHFca4szs4qMqPVbUoLGgDCI
UtfHBkhJ6O5AR1EzBT5S7YUf9TwFMUX4yBZswnLY50siVbF5u4pbXUP1VMwp/ffPKbikmhpY04/S
Bp+gjb8ZgXguSrmK7qYvM8aW8McKmFTWsvAuHXE9M6b6Zab4pMtwUbkAphdRImpZKbvTQ6vt6gCr
4VGP69Z9qqUVIFifPbeezJwKR9Nto7XfsGA+McL3tKD6DyVD5JVQ+mvD5CC77oySZR2ctsOE3eYs
/83tldn3O8xWDhT4tZTFRxVSdS8E7C3bfZQ0LCXD+GumtfEKCidkaTqkb2Pj/OOchsjclupWWe4I
tUGleAmkIvxfEuorZSKs28KZS8FFeDCcv9DyjZBUlZa8cqLg4tIg5PrhU+NfTJdvThwYug6HYGFe
038aX1j72X1fa3n7x4cH0siX8TTJoWo99D3Mj5r5nORiobqlRbEjxe+bF+QTU/af1UjPEa862Itv
xugKLF+R+ZG0b1pvYItJM2u0D1xbmjXP9GTY5MQeNw3eXAkFWpS42Hj0/hkEfSHXkISkBXSNa86Y
aLZtQpQaaaYnUZbxQDQ4rmrq2fI4HHobot0eeCdV54o5+KzT5XU7CafYcpGC/YD6JiUlnxxT8Wk/
6Hyot1Xlx3ZS2o92DswQp0hso3x1bennqFCCZg3w4Hf3bqAA6OHK1qRhjQymgJyKY5q8cjdawUVk
d5KPUP8tch7JSjLBWfQ5iypjbA59Ju07ZkV7ZQnrV1u7zbbfDgguM58lkT8HijH4b5Tl5Udl2ZYC
qXE/H4R/I5YS7JRUXan06BY5smMkN5mzIPycEwstXEQiCyO3h+lyiVTagPfkknHz2dDkbmAJ+4aE
ZEJJR40bjB3rurjB/VALhrqxft52dUfVn3Zlp2PYGyFwmuL+EZKggOfnx9hPKbbuWTKLDwGAXRfa
NySHAHs5enQ76xqJ2y9DuFFotvlo2nwrLx6cbTjiLKJuggBUuh41yMyT4W/6MRL+ixT9F9FlhwPp
svUHsuzlyH8XYBInXbg1jIh4dUHuxum3xsDbl0MSiGcPnwsNdbeH/4gdtQaBLgK6TX2KfMLr2vMD
1tpLSFvPAtJkfqjONpwIpnFPtE8zoaNgWU7x/R27RPKSpCdYygg8fkZ2EJ8XQIAbS6JYplDrJbu/
bzbFPTkdK8yt4KWIXHgNUaO1iJWJegqeXnOc4sfReyV5E7X0DDaS5JvbdV5NK7mcxE3V/63c+vPD
NdEZA42zaDOcH5mWNnD0VxHETMFZs0hw98ZVQxwtK5s2W98PiAR7FL8sGRNW7Hc1kXc/ObvBF0D5
Z5pu7uUJIumsWz+ugRSe52mdyWBcCpMJ57OZZFRKa+6Gft6sQC8ZbEJZh6mLhEc+j6/X17PIh13j
q2fHDZhlrIPn3AyOpFy7nUNul+ZFxmrOKKIlbrWn/hJ1cpkSn1LZ25/QF+D3vkXV0BQyBtw8oWI0
aMiTvyfkwIVbgbdXQb/HddFG3asw2VGBTTD4NNnIwJ4ZOhpsTop0bdllc0+150+JpliqJzlczbZi
wRkDNeBp4GzOgBEXcKSdZdiyhcr9N3DZLDSP+Rt3kgFsjFYyx4xkqMshZin89KwETk/IjPKX/vvb
ezkZKKAwkbWvT5C2rkjjLaOCINEFuyeN3oxRuRdfi42bJRxjaryDOSZ8UszRryRRaRbvNdarsi4T
TsX7e21H1yFKIRBTSpfkVZqZDawg1XLThNYOnLN0/OchZiEcw+U6w7C/e6L59LTV3SCX3bIC/TUB
sJ6Wohd2m8hdzovnLJNGbleVoOzeQUYCwaqAiji4FF94QGrBaRHjjZE2qjX42/cQJmplzPg/3/Nz
F78t8fNS33z6rFOl8uV8qNDOZ5BvWuQKY2n51tRNQjM9pFQzGcfDpQuXpdr4zqlIkS3vpwVmRhzf
xxiL/bLG9GvacmndQjkWOFpksDWWTUZCSNWQhsxOUqkDGlrm+rWZW7brIvhPDa8enO3FgJImmQOb
50FCYMrv7UOaKZ/PSU7qL/EMVPeHdXtxngAypwC5tGB6M75lo6cj9brw9DOJjgxgcNbEhSwC9ADP
xQ5dNuvyZuJ4LqbPf5TOixnS22SNekW+QbImyghSzP9bgrLyRs49lZxQ/zaGeNZ3hqwjPh0wF9Go
PflrTjkmwMp54zadRl4pX9pioLWO7ybuyW72hbHkTxPYEV0Z+2VHx3wAkAZ20tVubtEt09q+d0tw
CIX75yJFTq+SN0fg6TdOVRJIwrSLcLpsPYxa27cMHeXOYany1Wxkj+BWnkRy6I0dduAipmhhqV++
byvKnxYM/me4y/hA3OrbsEMGXGMgHnfANHKTHfiTLZT+6g3cJ2+/l5OEoVzdY0Cs0SmZdn4596AV
R8Hb06XwX7PFyQPOFXGG7lODP55lHLazI4y+PtHtuiGOR/hz9Nf1gHNm4MuJ1ZMeHTZv8CuNWUGC
qfLb5QD2mDU6Q7YdVbIqP0P/Il+0Q3AVItHNIeMamfnYriGfejKyOyjaCPr6eVo43F3Bs76lFNqw
PtwdimVZ0/lNmwKoFaMicCDc6K/kjEan96ZezKvSUDL51xZMlH3ca2S5YWpExvk1OcnePgtaswOq
DC4+weC8BuzUwT10GvWyZx29AIaE0Y1aO59g+crrqvPKg7fwjX+4r3ztCZgs8ih4HGwMaPInwW9B
Re7Gu+61mcCVNIceCpvaI5+tOO7esfN+3QXf1JTRVtsPAw/z3Jz+oALlck0Zt63GyLS2zNz3m1lh
aLhnGTvHScciKuNbVjhzErubrohsHUCNQK9CPT5k8MZQaweM1EWMqDmLz53v8d4jTmc70gFMoxCw
l7j+DRW/GL1C4k1GN+DY+OqssyhPvokUYweVDqRIcHewiz8k6tJJW3p3m88VAcTcRe6ZqHAoiWQj
VpB5ZL++c+L29YLzevDJUMjnzt7GKSdAxNhMxtvE3QjYdYEDOloGBRpHI7OKDXWrXDRgfpH2lvSO
slgwTZexAIGkqslE3O28bmY9Fza/VSsuJlatZPKtP9gXA3h2aRnLAFDtCaOMEVqSUvLPXp6Qkr3L
NbXsTQz9wtdJ2yrWeqSryrhj0SuWZFs5aUJNgG5WCbTdJvFE3v1AdxJw5J0moThFdNDtFwH1Kuce
itjVmOH+2yCg0Ve2qu5ghYpwE3mdsae94C3FubEuZ8mSp73Auah4B7x5qL2FwTC+wndSMxqLpsAf
ikKNwmfuj1NkNE3ijBFM2s8zjESpUE2TDPddoRw/1dodrUPoCuoMPYwW2+vV2s+VOjzId4Pc4b6o
T/Q5eJ6MguANbsRmiB5y0KtTjuzkCvv9NzcptHG5XCo+2vwpeNYQYpAtNy3KYaNplmb7+AUs/2oy
sWgT4QgSgVrqCZdfkemJUlt1UIBXM0Uhue8IYA1BiQezuhSLLFpMsbTHq2GhVq1a9RybDxLB+LoB
8Dddu8ojZhPSDyDE0lknbInu/zPivLoV86pTSnkGTCkbYpmWtfHZqryyWN47Sf8gwtMtxS7/KjUD
6GO5NIh8fmq7B3r2ZEF6MHtL4MFPLaREHdvZOPVRIyZv8fjWiku6+C17sx5tV2acnjsDnbfACoaa
E3I9BetCa1cUxpdTuiFJj5D5EybeTOyj4YHv5uiZ02lJAaefX3oblZ2zFcgzZ0bznhidETYO5Tze
jSkj4ELW9PWr+DwYX3kUzEmLclHJ6FcCY8Im9W88Xoqe3GlSwJfznmGi7PfX3WI4Tq6NCd6C4TNz
z/W6mUtRxYKCMCXPof8mrr6CXcp+F/Eh5PBBtc3jzH+7aD8R+tZso2zdPJFkh8LEhn+lybifO/Tl
iag1AVEDNBZnl7hrmujJ+Qw2q/XMpg0B3B3CTKjVdIkn4mn1xJTzWPaYzIOUN8PDFB/Ed1jUyWBf
1doOM2I1GmEIzpU931fdydQODRzeSC5ZioQ+b8EpoeAJG1sTtaKzAcSzbDdGM8fPvn0ElYTttUew
zcpxRWlpgRs55xHxuFSET+KccviATtzYUWfPavNDPpvOtcPLhNC9MAA88+oy6KHP0jo5M1mzZ1vr
h/xZWDOuNbtO2ZKGVBCoNGkWEaRsDxeb7RvBpAxfiA+stnHFb0ybu8Q8BtOVOTKrG1zMJv2dVsVW
fRE9wzLh5QgsSD6agOtiS1/ltx2zyvmgx0K9NQmqm1tPcbxAcjTNOAvRnvOffPIgT3G3mUyBXydM
1F5XEkMaFyktdg4istKCJ8yRmWxHBXNwWLvxdiia6zHtk84WA3bYOQ2twnW0ZxXPDZPT3mMINPQY
ItQl0JAG9m0LYiMmKtwejpXidvS8iZikZjbxaxGEe5g7eVapSlFE4X9jGLN4+KPFMnJ0Y612WchX
jvF52wpro1eVj7UBR62yHqfAYmxgHI+jkGsxuhClcv7JVaVHt0rdeD2psYZXOvYjkn9Rioby+/V9
VM/C/w+3NkFAyTU4OEsrXnHrOXbm1hFX/qoED/j1L44kF6JNDHI25+7+tw/N6xOk7fLhLoC4KJ3J
Q25Wipq85r63fR3810zJm/YrU4pS9H6E5a1y2rN/t72jhyd+IFrJxwhCkEfgNLVfP8lSuRXURNro
fnIXWZFdphgO7fISwhYi5klh+qy3FA0rYv3Jh3EcjsU9ACwHXTVB9rp70B6BCSDt9Yab1Obkazvt
J1SAg89r1+1NCpVu5vzi6uD4M1lAcDY1c+Jrt0s34hB+9nghW6O8Yw/Lo6U2c5UAoKmE5MZlaRsY
As/GlnvLPKwWnWgbpDFM6TDAjaeSN4QCIXIGheumTblwzW+Wn174RcWBBJuY/Obc44stMgw0l2+l
Om70grc7X17+O2JfVhNrRDbyGPAfIZv4m8hLkhIxMSPGQVKie7MYe8pU012pWPORCpo8DpQZQA5E
SqzwY2aSadh5xUhumQUltaFw/RL8E/ZFL3NF3QaISGmbKyDRcEuO5uXAWE78tgBbcOfeakEFeDnL
hTqAAZ28O06o45fL+3Ih3LrXqAeLXWkh/gtjXAKg33y6bsXv/GdOOClj/pJOQ2wyfQ7d0uMF2vjd
plb0TCaVNeqE1o7WCG2pNg3WMEYCdQe0lrzWN6NO/WBUKafcOmEko8RDNflE3SmhmscH6ilFmfGF
eeXZserJ4RSwyxX68O0GIUEaUwab73YMkWe4zfy7JUg4cpTpsRRCLsKI9CL8FcdvY9arITSue57Z
Q302ygmut0uk/HEP0dMbqaQrLvOBChYTmK2ftgkNqXJue8YaMifA+dDsTO7HxAj9PrKsfbxThL5s
wfYOvUpbXaOAv/TC5koj1mRpGCuOLL81tUJFtkf3DG9jNn0gDMUvweIArq5+SIRXW5KUhhqA/J61
vnRVEvK49B2k5QGLETYYjs/1iT5g1iF+tWUhDFZudIKf2dYYf5BiejUrcSUS/b4o60rf2vjmWw2d
S8GRk+fVQRDDUs3fNC8/TtsHfPfgMp1bfnftCCGW80/FNcttwTFifhOjlBoWPvx++4cTW50NpAZe
rbvZsL3FBOENrwa168TC5vqOWFdc++S3WU65EHY80Xs7PwQ20sbvtT67g/vM+ZYGoUzBz5DAdi59
H7WYgKoT1Jqn3EZn0F4i6ALKbZ2cBoYEvcs9WMqlaLVLsp8rhEaKMh4WttdF8HES7BRicXgWKM1j
JmthB0DJq5Z3PxyvPwxtdPn2sjML9ohuM2EhNJVRDFuvp/OPTWCLSIXxnin0eLnRBUWFxdoDbyA5
azMEahtHpyrS99lZF776LECZ8bgYlbSbNrnttdzM+PHTYj1d3yKUlUoSsdRAna1q9G76cyxzH9yK
v3vQdKJ+4phwmc60t4Au5XbvJBkYIOL/3RX8W4A77btvNmIbibQuvZ/GzcobwW1GO+v5O39vA847
o2r1weuhLbKWu3tvw4yb3e9WrHEho7iTa18dP9s5CnQXdF8eRGUILchlw0D2UBFrtfTDXBug+vEN
kJ3Q951/y6UQrPjC++K/ZJh09+n3d+AfpNsfq38TaQT7oImkC7o6wXcfuqO9INMIMMwxmg+I9foW
gshuujpo1XWrOFNbcmpgx0JnMxDfmyv24giNwbavcFuLPReLN6RV4R37slQ4rRcu3w4Gc2Sqk5/C
qnRzWrK6FZI+XZVrCnFoOXZu2rYvSIUw6vnXv6/me3zSUl1LLQhvykpC8Lp5qJbn8xO4QOv16MWm
Uj+I0kPifWez2B69EtdIPqbfO/i4PtcVtM2hN06WKLjI6KeNB1eKurYOErLWjNOmal95zbw9WyGj
q+wDwGGUIrXbOAcgsBwCT18zJUW2z1bBrkJaMnUnec5l4gxIHFhlJ0+PQIWCqeZnckqPDuty3rhr
KCz6E1P7yMYFtFYuchdvUGN3BbOP/xsmHYQeQaTDf62KEyMGAkXzV8ACGCin6t+yuisK/QfMdTCC
nIimbantHvxoJc8jurFWY07MtxzOOCZMtearWOGtA2RXRhK0C88w7yxLUw3O98pc1NNYSTXp+hfp
P3cGMuLQoD3yUdlVoQYZmOTVyro3JaG9Q6HK6nzv9hE8jWcRS7MiwaULeO3iSAtakvMQz0Hhk2XB
xvvIG1Ol9UixFlGU1NWkVq+N+nmDFvClq7IJjXzaZ0kUyS3KNBXhBzvIxSWEJhe2P5OcoSh9JL9f
1wS2QuFUzvjZPhePTaHtQAg2v2MSwAlvFIc+VkCKBoJb+lPLgF55kr8VbfbuL9Qh6whXMlQs4KUU
AS4SLMSeeNgf6fbm9BFIrFkkNI29+ieV7gf+QRAI4+8d5aPA8LMELYbLbR4Z8TFGXdfAd1fdqI75
YRBK/WJc7LzMowq3l4X+cy5zgQ+B1N740burs76/Fb8kRAeacd+I9CM/UbzlliNoFKvaTDcob7LD
ALNjuE/IYCCMsS8M9UgBsxS6IRR+KUOny1LBPekVRHKRfa5pi/9oHL+5mTuSW3ju5647l/SGf3Yf
xw8Fo/ozPWskaKEM3+QtX0LdsiIB81EiesJrMquJ2yYFeEMB/Z5QLHMLteqjiVca1x/lRZ5XjA78
pNm54yF5+rPWXPEQBNeiupgXxtGnOJBSsVNWvd16TSGjKrXK15WVv23wZX61VaZp3MEcJ8MroNGJ
l0ZVQJbhG6bqwKojZFq15YiBeg+UAo50PYPOjbATxJZ4YZwK40KOa7SVbfzqSoOnMjqeJZkNYn8m
qkkHPx4NZ8/YxfMycYFNkoKD62T8ovh3veMjnB7HL73o/+r5nUelj3hzrMbvYEfCpW9bAooYWHJJ
+uc2DZAhx7Gls2/IAQQVFokL7rRLrwC1bKT15NULskudIn9AMB3uuAmseWcyKQ4MDs/Rv824lxdK
Obz+hwRCdCV5YDkyr9pYvJmtSVdF53yGqXL0EmhvCgR8k9wRrVNAJ/6Be380O32ATcav54wpnkzo
ekzCubMeSpoQ0oZJfSNnTdHAOhVv1ncTwZN2oqB7C4Ovpp1sJ+Kjb0aIT56UaipNfxJCERDdSNHQ
xAqnZcXN4VBqM6BwcCg4r2wJklj+Bey6USr3nEH9dtlFgOU7kEC7IJdUKIhvnahs+ofVD0y7D+HK
duVJcKvPF4ZnN3dKO1ex1yth/AdTEweFyJhGiSDhwQ3uoi0cP2K4usa2ykVmskZN8EKutpLnF2zt
uztYYbvDGcSaG213By9lPUFxGGrn19mN7unrYsP046q5MKaQCRqCBBueeDKJcZC2fmiyRxZnEWoK
xffe8wDQe5v4f6DRkcLVIWgcrjh3MRLS54GpCvxSCUvVpJOVTbwCQUHQBOdZxl2f3lhsBZIS5g9i
xxuk229Xp336ivj1Xz4yTGJTSZgm0l0SV6gXn+lz/jD/ta0/AHof2YpSmq9djyHn59ZyDwA3UPcl
ZngP49ynvNqntgX7eGOq8/sbLvV3f9mpX+WsyyD8kQOoGVL3MPAWwhIzqPAAVECUO6Y7pq/tg7dW
+I3M4Px7974rnSbmFb8OkmGxoB84NOrqmPlHulqktOpHYcWQd+Rn6wKrh8b8ENhmtLNW550JvtN6
AYR/Mg2OJj2oDBHGc5XcZiOfaVEih7D+7iSMLAZO42C4oIHXjhq1JP2EpsWsheN0DjlRMxuRbYlz
8PI2hOQCnyj3wBWY4CiF7grajZSUpGchAI5dPr9sW6W2BVQBvyB9I/pgClVKciQinjhBZ1IxGbJY
Ji3P9P8D3UcozZZcvD2MhCOKddfLRxejrkzXrfV+G5Hv8EMhi4GIK9xWtkXny9h9W49mtap5xC8A
mictwHxwPuzGmJqmi8pFbE0n1xcX+1yGwVbqUzKo+BUAkT1a8eovNZ+NT3C4Yyzn16pPcNmAeDPo
WFp8iXcRw6+ed0InOrz0pSxQd0tYiudEz7N9SVcYHhFucxlTSyXvUVWA/cZrjvvPS/lgGcqwVlGR
USrM8P3n+vVJMgA59AstvDTz3dXoOwSUx5mmcIQdxSyhP4km0k6jttSOZfVzFju9uvU0iVD4Up1d
ckjzRQg2eTDInrzfeZl467wkYJ/HmfFFeW2sVYLqhGTldNGdqp8w6wFXoMbQSO29NJdG9KKTVWDf
Ik27v04oNWCb/NqwSJMZiv983jqKauwMZMHp2VqQvwcn5x4GJ/pdoh2S9hBatcV9yCWhpdVlTUfz
vYVjSom/vykrUZW/1j7vYt5YLkW9osG/cxzHnqh9PAjXUZ1y4uTDrWqF86DTqcxiHrF3Z4lebU/m
zBTXRncXFQAyD55GoCyu9g9Levj87LTa4ooZKFxIpFq/jvq8ZXO9zqQPEiRAcABp/RH9/m80eI9F
qe9V6ywF315y2roDqEQ+CMod9pVCXOfkVVoOKlPSjcuVB0y4lehysaXmqmSSHn4ZFnjtinWXSfLK
JDkSjJz+VSPQbYjn1odmJ4iICTxiB2mbavefALoCGY9E8+ophSjYRU0uQm3YrQtdv6rJK3NhOdHB
bNLda2RvkEGK+YBphIH392OMPFAT19CcG9VEMduLdOQf3FOvRk7gaC7bvyjcJucqXT65teoMWrOg
SpSmGW+EX6w5pWCJHwS/jTLFGuBVy6YfLJdAbbv9ENJihBdggATBoA7wJqCljCtNHc8QDYnITuLh
v+8rJPY06XQaLnDnrpMiZczx4zDOgugNxsj8zY/lnDYn3Be8idz5+54cyNBeHoMWKPEuGyvuYAv1
0xNR7dPYCpqguJUr7rBVIT/dc+PObwnIjeqQgfVRpaTPWfqDNNKUMb7T8CswRxWQcP73nOFzaTB+
EFLdvro95dU8/++q2k16E41Qm8Iw7RXwzN8MAgsIbNcnv4AU8PXNfE7yJ+WovV5LaUOfBtwRZsam
56Oko8BJo0cI7Mn6ofmdYnbG6CBAKPdRgJikQ7VW3pinje0WnU1KR6ExNOa8HOnBpQs4CRxEHR0s
oN3z6sLeVj1oW+7BVyT2+bciHPySTzyHizoE5QcSYzMain8jFjh/GZRrLkUUVVjtEHsdBN4nGRN2
YT77x96gR6svRbJquyspUcRSttz8NY59ah9CLWbUGA1iuiMn5aTlXlzzCi2yiddpvf0EYv2aC4q2
9OhxtsWBQKRhWhIOovUozH4novIoO2cYNb9vTh4hTpiB5l/zI/JT58LCJwAr+9oTT5GlZynR7EkW
Jgn2TZMQlTdyjVbdeEPbzT4gujCbF50AjLRQnABJRDJumj6N9x+frxiWnAShLrig/qIsX4QxNCFs
ILAmVNZyowycCedwTdoQU/bMUaVSBB89UFDatCb2drDyoYhE5jW27hF1ovWDkya4+wgHjZ7rkG3z
GuLkppA7ljIvj48HI/PBa68Xud8HrsIg1zM03HMojs2mIGDlT0U/iSSkJg7Qg3CmIFLS7V4xLwwX
IV0F0MB9/p8anG6j1M8d0z/vErEojDA1274uY45TnEFecoPeMKc5N6+3AASFVTUTIi7f5F1aGMcE
KY+5uG5t2JxZ9NKZOMECCUSnZtvm+hl9flIPzvJNPlj7oEkXmxUoaT9v4CmT68Dm00gCe2Uw0w1U
e2EQW7l2SfpFJyhvPxU7Vyo0JW6JCiOQVTcV67+f7u9EbzR8ibqIs27cs6vHug1TWoXc73K9HcHF
8W1JDcMuQDluSBC0eiP3uyEbQ8LWi5grTPEKjLK2a0IzkQzS5FqvMiQFSeA+g25p9tXjaroAu3KK
KWe8TBqPjhLHJNYgy8VfFRvLRl1f72H3jl9gVCcmysJ4rA0TLexHhuRWvwQF5Fq+Le4yycaVrd2P
2nKgNjHmWV+vtyT1/JVa3tyGPfltecOlf/yf2MIaHASMAT+iQZZOa6JIMa2dgGtUTsDEOfzDJI11
RyhRiVw0NdE1wXhf+Dwk89ZAddzVyFOoCAXMHAWzKncotMBv/GOGteYEj+crVwQMBIEpdy25/qlO
bNFQept2EXbbe9kLPvL1e7H8lf+n93sM65fXJ2rsrDMdnwOZVLweAL/pYzorQseMz01oVWaBydl9
36EfCpHO7S6uKBVWhgiF49o+a3G+wTr73YyByUEvAnd2dhgXl1IZT+or482VqMQIZYFxuAMv2RIj
BJX/WD9VEbfZZJR6P5YjmbVgexYXtUTxyKdArVVU9/MHMcWIJDxK9eXWkAZK833deyQZMxUJDCvl
35fLWPmkpcFY+TdRevTeWet1/SS3XYMmT2Y0L1m+9afigZfpfVVlh9R0uRhnQ32ddVb+wFFFMJwo
gJjrkj2NW4aXny01E/0ft4THXnMK1ZqCLuLOlMGbtQoeRsprAAUFh7oDHkREvN70yPClKDyxqEMv
h8371k8xk3UidE6Hk4kfbSrNZr76DXMQrGAjDzLV5/iF6ArObFLxh3khDpREA8SXaKPFMLQVYH+9
u4MnpiyLyxdjA8HtFjK+obVFlyaQdNUQxUDH1YjdC22aPxhDAse2xdesItjoOOjSb85wpGiHfvcx
uJmo6PpEnxoTbVSlquyUWSG0d6oSfk92VpRJIVq6HTc1gTFrmg9nTJzvOE3cb6B/G8aBmI3HGxHW
r5dYhWkTer04pYHP0BlXYGNJCqsUGV6W1+dmRIM2z2HPogaQEXwtJadWqYBa+4Uz4SRAjQA0b+Br
Eqw+VDGP6mpXRvvxFcRvrR3a1VktVnqADS4pEn5frEKxl9ZT5odUz33OecvqD28k1t0SannyPEmJ
L7qh5UzLxrmw/fr9Ksk62JKLFCHanCCOEalrJu5vX024bf3jcwfuuuU3f5KnHXqPGZsKiO/fS2Ai
ovn+qf59sA5VQsvsSoplH871u4hvIsTi/g8NcMNrp7sgKFboS7gVhu0JM5VnTg94hYpoJXASMQuA
/HFwmBexV0nZZgahQfd65L8tqbhYg8BN2PX7wJt56DhRbDm+eHvo5jMwtRGkzO261gVnDoRgY9nt
KFAguyXrK2fHaTL/l/JBm80LGKny1o1HKl6rEfjfy1bwDSLAa5h4o3edjL5n8OduEowZx0TMYWb8
8h1UgYHaypl+IEyvahAyhbUvvaydj5OgZIQBA7wfaxjrELzd7XEow9VyrB7ThImdvFt/iyDoCTRm
x7PYv9GQX8/C2DELqZ8TbhlY65FHhfCzAXUP6t/F/YcQMJyAMG4bfQMBCGh77HOBQ6vOHxw36NQm
rZXjedJj+kZ2pdn4TNdl9BKmeKfEFDX706BHCiaO+JLuDEW/jDxyaPXIoKDy3Jv0dqojuJHTWOkJ
nAQO9fM/RishYQvQN8/tUQGUr2CiPzP0XdmgJy7ARPYfWD/JJYyZYFqiqLwrqFrnmNpKczNjt3gD
LBa8g0UjxGiElcvYlH9y0GZ/aXSpK+3wzlb6fTCSP4PsH1sZ+23OBfTB/Fn1gP6Q8id3g83wcxzo
jdNaAv0dX+wKWINVQpOhTNgeDGFHCOWSIHLu9YlBp6sLOLtlNWKE3QDDLhx/KkOOHKl166OGWPUy
/keEKerUpwsWI4xNtTVkn8DwtxxnIhfwX+UXx7xGvmtSxaepBnBIMBHE+xw+SLnmpK7JhGWqT/1Z
2NiiDN/z5m7zawNx0CwLR3tspz9kZDSEuKgl4olS9+g9o2uDOAssG+MIeM2T5w49g8uMS6KmlL4s
IwAK/kC8GjPHjWQVp1vxdCY7ZBT2+K0vdmcRd50HuWhvRYrgZmhvcLrBGV4HbrFxYwTEhik2lsNp
7GnLMq0ALzEIxDWvybO0ibX+zbvaoj8kuHeGxxaOMg86xRoj+ofDfFr5++brCXcO66yEP0lr7teT
5ogCzmXhTX9WfbH0iytZRV0lfQaj7jE3GpPBWZoahLAdoHd+vpXju1ygoG3VTlF3XowQ6zlkTCiA
NdhF5vCPv744Q9oG9lnYEs0oCucCBAya/84864enjdmcx9VVqAbmm/Q6dnisWHDviE/SXlKa3PPv
G/TiczBmhnahleC9BprEZkQ/T64tLyBljjOTkUuUTczgaFTMaSt/5kyXBEB4J5eoLzvb4dErCQEG
IEoCaUCTh+2OR6B4UoJLEcwqRz67syeeL5zAFx5O6v5c/VVrMOoW/POkBR2r71mUTsctldi64NGV
boPc2dpFoDrLu6OcqDTX9SAbgTLbPpPQuqWq9ki6MqXxjZM2LwN30EmqLoI288xLs6PBFJompYTU
zF1jgTwA8eDAFOIZjxdqSuHwOgdRt+0J0JNmv/y7WMHCD0EDHzI1PLvmIbinV0PcE1j7e7nvi8ac
G5dLN9wd1CgZsjedkZAe8dy7nQwpPzYitPHArUL3QJpQgNSZBXZUe8b7Njljo2ExJKxRRwU7q866
hksxNsS7BTdarPTf2PQseFbrbjCWGRP1BXBnF7+7w6ApGcMjHHLBVM5FAx4cW6b5tVzH2gZUijtz
6Wl7XlCBz25rfVQH91c7kLKERoAxLeEiJlbdNkLTGoV+rsMU0xfYJq/xXQAmSG/Zbm8vTiok22BG
9rvmce9HKNxZzuivxE33Ikgm65wGUvlXtGAFG9p4FT/bIGbHzEUt0+Ks9XkFMW5hEeJKVCBoS05L
bflVw2WtkFzaRP85vtvxA7oAQcAPKQ0I8K0VnOZlmt9AypPDFUGSBBwiPMcvraawGcYjEBvCbbcP
kTHYZWP3PoO5e04enoQ+3+sTBQtvMXL+7iLMCBJSSMkjXoQjcbKO8mTWedunzr26kGKi78QrNSRW
Se+fXuyl1pS85eLHYfup1RgeECqRRrqVuYGo/kcAtt2to1LalNVybCi1FbaxBQM+5MQEjFD+J+Wh
79ETwIOe/6laSoKcEa8Fs8SUM75m+nqKoOjQn0UKlLdMuA+wELYkLg7xNMMPovyMYcIHvcyEIJiu
FoSosYsvhtec1+AmNuwU24yJsJNfCMpdf+9drXRvv6ZhyaQhrXweVa58p/5Vi4uAejuP5Lm1pP6H
ajkd56l3wYQvgafTrvrn6wbLURU7BTP1adUO5WZdjRUzj76/kNIp4ysWHFj2ZpQtiMz3Hi6YV5Eu
Y0ORYDYoTC73xvmemXj2EusZ0Xti2PQ/FOp7ps7pC2DuVl1f9cc+iHCJ6VwDwkLnrrdRxU343YuE
tGhyD7eKGVroVmtWx7Ukj3EcYLZKh2EWnKq03VYuiuOBWaaU8j1knyZRGl4P2IqIW7LleSPHDlVM
MbN/hJst0+9itDAHmZb1wXX+ny5PLvp/UCXYZJ6/190nSTcJITVVoyNNbKvr0Hvo97XiQpczZIlB
Xhen/P+BapcjGRuRGPEVT+ecK/Lw0C11vvop6wzZ0OFE4CXWlGjCkiQLtmpOUGHS/Phe947f35xB
+2qOv4wSBBXnN0zWKA4LwcNR7iTlqNT/tQUTZx4w9iDkJgvJ+pf9h/yJ8RBW4Pc1f8UDS7JeL9WF
tZc7fh7d+LIB4ukHPVBQpFi+8x2aqB8vji7cNWApSIpgrPLtbWkp9aw7EphMB4dUG2oqf5QNFPEC
VmSHzF8Gq9ECBqWRNHTST63sLM6/pTRJcBCDqoKeuMfG2FC9YwUQvRbNgGH5p/ZBbYa74lTDrydJ
khVf0KXPgCgHKLa34++MXqxeEujR/dxmk+6o2xzqd+7IOASZFH7DJvmJ3i8uq+eMtJLwhdHzQCum
oG2YempyO5zEtzdafUqIRESCFbSDiQM/gsSEJ4IIjcU4+eNBaXlSz0iBLXO1R1kl5ZdQTV+6tplc
TMZ4bU/X8tx3yDM1zqN2LRXU0QlCUOI+lQRTGffC+EzKTnpfTF0Z9aFGhVIw1xlEcybxt2lM1pQ5
gv3UzAG6uHBkvw+QGiK32BLW39sXdXHQRKI0LMr3NkLOmr8lFsKx7vQcSJTdfVRjLSnQIjY+J4P2
unBPT8SMaHwX879OCH4VM2A/4HJu38vXYO+ApcRI+WadvAYbedG0SL14cupPG4S+1LW4/TXiteqK
yiV5p3U58/Zb/V3cRqDd45oRuAd4u6Zo5lOLTf1cVLi7mgbMR2vcKHNsibn45p+OrfN4I9WEzZV/
xEjylmHT5Z2+MAZ+LNPm3lc7LePwpi5Eq9u6+n352Jwun5zw1HkZ7T0TLAu+d+mTpWmdixCzZpu1
ov8CGITEE9kmRBEGFViLAruCZG/i48ZFRlmonDLNeI9RKBZaypA5AZ9KRqQPCImh6rtwoJmCZm0n
gB5grdvee2a1Z/ED0jekF2On4f1DlkcX7H0kTQdGh4oNish7tAjjQMpIU94ysZLid9NPZLgwD2jk
fxmFL9fkr+mJASzvfKscsOjGJYVuKMWQja+uj6ef8FChDkt1815xgO7NAG5IXsn1A7fmpUKwxvme
V7ngHjz9zlIWbq1OHP8ZJqb9Uj53QH+AdwAoV3WYTaBcxEvz7vzJ0Op1KcaGBM+nXl+n98G+KVDJ
Hf1qDjUuV9803iuZ56geL4339AM53QqMv48V9etIR5jMlmtzCrwh/98ifHtWwC7umBLnMc5byaac
qibxE+zEFKqUznyUcLSdPOcqspjOUlPHg8xGdnMTHGU7y+5QTcWHjpxsKjpO/j4BxgwSAw0QOpqc
WXbLhp89XrTn88vci9g1FXP0oVxlu8nBw2NCsCVkVtHshekJAjW5R2o9cp8iFQHzfbe+ijAVXwWy
klqNQfJfJE0Soc+Wq/AxWjNXWGfVCflfvx+btBCe9idssZ8ub++hNr1SnmdfGg==
`pragma protect end_protected

// 
