/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
YULis2yomg/kzjFgzOdPLWCb8hrAhUhK45ViEVLTPnp18MjTTmAMM2+I1/rlC1Ev4I1pj9QnujWh
m39etpBwRlS+aTX7hc+VhhAyZvXM2DZ+//Sndik2DdCY+PoosSQZrDjRhqeC56M6tvG1/iHFmLX4
wYfLo4c12b0Ht65dwcJK5COfOnxDnqDfSuZUsKjQUaVd+Wf3ERz7RS5uzA8yo0ZDybtjtZhNTdDF
dr+nJpP3kGw9+QOZ+hk8LCAwpgkPWQInSQYkR48tPcmAjrp1bBGqrLAB3UTT574+5Zs63JZWTOUi
FHz3gvl87LFRg3pbLvTzIMlfqmXdG4Wy/MJdqw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="M84hzKro2ZXjH3LMUxD/XumzYV1S/vm8jkqX7oQeRN0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 848)
`pragma protect data_block
wknJWhNPnGnPPHAFxd9m/1dz3A9Q88xlQ07Q/+NG//++TEGfirAWviyPuLsj+uuYB/or0aBICFDH
BUKQhZk9RtEENxtvA1mJ2tnZrTNqSzOoWBez9l3ftHEB4tb839CkjL/6htBLEp9pD6JqbvdIlIMy
pDK0l3gNEX4a1IMt5XLz37XToPG20f6oDwJcKLvKqz9M7Ycj1AzzEac9NYUcxwSxmkOHfYwRV5hX
aEge8ZK94xkqajwAMyk3DauUdH+18lDrsu1+oXol8cwyzpBS48t9FvI4bcideRTP2cEDL/fbc4Nc
lm7k58A0POUs7Q+xPxLWZly+CpvfITXvnML5emUrYrNoAD6xBAoj1P7Qy3clV91Dqz2Yu1bpVCJx
T2r/wNvXUt3ylNTtvaRLR7UU+wL4NTJD+ztCBsfR4IU/lDi/i8rg5ejzE+sPJFGWvf5L0DhwKs1g
Gu5TzwUlF4y9I/Btd/JTt6Ust4mJJWbO9utLeQUyJLrpuRTZbSd41XtUUOHhZefrFjY5d5zNBdmB
BgYcRqZ8VXfC6zBqteY9aBlV0714Zry3SvR3GYpj0ziWbp1Ty8KZSJt/hRM9OMNRZ6lCMJ58//S2
vbGrl/DFXWRY9AtrRYWS4pliSYcWVXWBDKPe42u1Z7vkKpn0ME+DoJLkxnre6KrlJXpkJeWv1RKZ
4KCcMeYJ6TQVLB2sXGuHVOE7kHwV6ldrzb+X8KMPyAexzNRlkuN4QoEosxcDag1S85NK9nJNjF5E
rw/gxp/GPLRYaQDdLUrr1rpPZP7VYPBMPFix6snXTd+sbjU/c+HL8IG54j2MhB318BqNrQObOpy5
eQijKXIRMcqGfG4OQ7lQ+tDAGYHTnXrYqAXHtplXMkxMHUA2SilziAZ0HebT8IamB7NITqmC9ps9
WhXXl8Vl3ivHBDKJtU+LRp3NaFf+nhVrHS2FSLcRGYbpo6VdNRiADZFk84WvzJT9al4CogjP43t3
76pZK9p//DKSRC9kdIoxc3CCZoHY9yb0WjTlCZDCwCbPRAR6rOG1l7BqJnJwrAJJv4fGT5IMx+vF
W2d1TUx2xiWWWsMWAk50eWeRicFnb/SkaQ3Eghkk6b6dQ6OTAWMWxPdZ9qMXq4LEPL0=
`pragma protect end_protected

// 41d051e7f991c9dacbe8d368b85f57380b272bd2d7dc26e6c472a2d06e70908e
