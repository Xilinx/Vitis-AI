`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47024)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPamfPOr+rPAO7s8fOE7DMw165NnF4LypmOhpB1U+tn6mBjDcdv1/Cf9F+5K6DVtyOku56qtj
3eukJyq/kFYbJzVPjoYEB1s7gpnM1l7Iyi3CTXedBGMY3QfcPyi8sq/Hll3lpHnWHJ4XV01aqigS
v26MBpI3skmydkp9iSaDD8+KSrbPUfEwqFY5myfIZRMkU4wvF9XNtBjgqIMOTFH/JoTiqcGHNn1+
7K4ONA4Zu2VbGK90BdZzJdD3Xopen94KvA/wmuCAGbD/KtMFO3ix+uQFytXRTjxdV0miq4Hecv9p
vlm5d96sDldxYe4AoAyFJlz9jUtghRTpQl3b//7SZs+Yipkvv3vKZXFsEagT6/GQhoYTRE9cKI+6
jS98Onv6HZzqc7CfV0k+MLxh/qbWqJJfgM5+sl3j+bIltue5OO2pZ7T520d0hKc4g1ekvh1/1crH
1SK8+I+RrjYIHExQCIz+QG0C1B+lkAkUCT6iBtR1oNHzwpQ6M05mVLGYFKMWUYH7FX2q+bmAL5uW
cfnzybqJRCetcrKCcrcKX9CQ1BBmmmX4Rrog3noUprVReYp0EYJxmTIs1H0SO7H6LS5sie3JTBLz
sF0r/mlfPJKQ20uJuuafhD3CHExxgE4+D2vH1en4YA/f2a4vZceR5A4BQVVLgZELBsgJ7Hjz9lky
w0JgKwEa27aWdvihMlPDDaaFJ84JTrBpQgWYJ/Bz2jsULW+E+QCh2cWNMRnhBnEaibnyKiGs4qet
alQGG6wcUKjMPQpeSnnUCQt800qyr8Wa9Kayw29xJrpFGBk6kIqG+e/UwiTROQpJp5AKsFYGhRIK
C3B4x5Md5yu6yMhSDkI41xdNH8mmh2O01iZqHTaVOZIvoEVSg5ojQFxgYv8fekpvf7jJ44v6dZqf
K34R2Ag260aCDv8delz53KStKvpNAhDbeXbTAKtiloD2VF5JIEzahgoxH3Do1rz6MEsss69YqriI
dPkRN5rzMziUpaVlZbet/WwvmSaTJNaUaMMjtqokltKKqS91z8MYs6lnbK4JaLvD6V4jBOpWz9Zz
XvSWuGoNpclWLlvs+CXjv9veWSpFrvNpyz3i/kOCa7MJNgJCXLu4EUvJdKHzu7nrU5qcrGOu6CBM
UzPOUcJA2E8t+yUjyS1zRe5XmfW1bhcIe7giW87la1yK9bdugJbqVZ7fWUNRrUcLp+LqF7tfEDSv
mewk/vnkxi1cAXqdaPflM6iFVzg11peZyuNyaiq4h7+Pfedu5suYW+2wzkVh3xXauAzGCPb3SpqV
xXnc3L/LTifNKbmU2XXx4lXF1nkndZQbInEQ6wj+XnDc32UiMXNCijc8n9qM+ZjOvv68bOzJE7ZA
9UDxJdOrEnnmNNLntPDcDnK/NiSXO78NpG3wIcaRsmqVWLYw61XKM2R69lbJLeM4hYMxPus7PjEl
Gp4Tuk50gfNjmfsMxBvm8LUdFZQCDmjfQFW5j63E1OykHJn4RFMiaY4+kjcaZEFyc+0mskLGwwid
1jcVjjFvABKa7TCgkIRLihezYJ8a4fHVorCHN1/wCXTidMO4P1omJkHGMqfrfEy6RROBW9iatFkv
TbQ1PBNIJ2ndZRbZFv+NJn8Dn1QLI22s436fg/NJLXZtiUypSl8u7GwetPjujo12AK6wc4bVFN0y
CKkY+WXIuTMWc7V/aiiQz4G2nqu48M3bCjQVCFAUlkoHfvM4lwdg6nI9Vyn4ibw7gdMUbA2faTVD
7Uv4yw0A/m93uYLhqh3remeWGgyhobLyivz7qXQxtJtXKo20oHrkP1SWp2431fcqXgR9gvDO/rJR
oNFECPDPNChuavbpdxDPDgVddKOIiCIOF6bLMn7yWCAVeqIy43BtZEuyciy3PZpWHx1f+reZI/UI
JrEhNgr30zZw6U0ngnZSPUCZlHiUvdJ140CdaaBtVdl6QsIMIv6MxRX6yfo/P2CcfSfFxBLsZvp2
IAJ112ZlC6sf8URP+cTfvtcCO/1/GzKmmi3fP4g7SpIQPVT1RN0vABQErwMTETK3GBcnE2x0LlM/
d5jO9eXdS25JW7mtJC8/pt6RMDSt5+HD57Ckd1bve8dh5joGZM1YuWKWg5N6wrwLbIXPvfQsWObc
pWK5B5oDk5Fo/bqGBwPCODGc7HERnQ7Zd02DtDx/Suc1sQHt7daoKKbaOZXDclqslUphXaBzrZQ3
6klBdvIShedYorieE/xBFkoybpaJ3mDDxdx6xJ6qNBnaS8DA1cmLvTOJaCGJfJJ/KH529IIiNKnb
C0y2DpcsR+KYLl+j5lgygxo2g6xBKnN0kxqiTxVQDFWGdn/9Cwu3Rz2oeF6r9z3UpQPF762InPqS
e2Pl+TkFeuP5A0k4tutZcPNsUNzujLN/6NPOXwGITDlEJRlVmbK6GFeM0CNgtTdBgogSiipv7CuE
w8A2eadWvjK2Eny/D0pAieRLpGzSMb87uBhgfLt/d7NFrIv3dx9IzJPwQV53xmBtTVx3gr3plsv+
zgjAs494M0A2MYgoLJDe4E/At4MxrTO4VnrnXLYChJlIjxf2oqFL00gzqv1Tzhy2xw2bOSj+2sC/
u3lTm5FEC1kSspxvWQ4uP9SzkvdCfe2c7Y9tZtnitSM3y2QDjHWnYtBWsq8HiRuMKQx9XSo+K3H6
+zoer+2P1KhXnaM+yQ4TFAx0UnzYmp8xlqyMPZ1Olcz+b8v55W+74uAWGPKZ0iMXcjytermTD3M9
diA/23vh69sCWqzlrsYbhPM9AADEFITg6dddz/iV8l6GMH5MPmmE7N7rt+xZqzFxLf9EknB1h154
Us6wVx2JOlL3w/YSjCYebQ4XaS7O5IRtMY/IE4BRzkc8Ty+NLjhKaR4F9haSvQaBuZym3xVCIT1P
aKDtJorPtDYVh3v3AYB/Lss+ZK7GQ4bXFxICaoJsJ21L+9iC+1mVrMK8g6xa+0lX7ComCOk9YQzm
e8nWrgA0hHCluw8SyhPnBaUxfOGxDmQRvo22/szoxi44aPYry8CtPu6dybO8R0tYA7BrBCSxX9W8
R5qaTks2ucIwCeop25s8+RleGAV6sIk9923rDR68xyBFvJbI7RotlN++nYIBOxVu9U1+1A0Pgyp4
VpF4aoHGemAyr3p0h9Ec0xBJ37M9IYskBF3m8NNnjCwgkITIB8z4fFGwymSJZ6TqgWjmfK2a/sYs
xEYaKX81GN3AszAlr/Vc416sRrBSYEGo021Pd3CTXR7u7L2rZt0DAThXlH7uiDUYlyIQqnDu0/CS
1I2EZex0eQgXAuQFgPQTKEcZo2zc2+L1ZLX/86KAjvlpSnGOZySKvKqWJJrqFCBmPl6DoMzoA3Sy
x9F8BvIQOE3xs31JOUA5hT+UZcIJJ0erVp9TsiiwaY4UFAI6XjgCdp4FyibROZwcHwasN7cn6uvz
KfwL1qiMTFGlHBmpecLWjhYzk1HtWf9iFpDhyt04uUmQMVvGg+fuKwhUOa9s8mpTqa6/tIdYzQEl
Bol3md7Ebf+eIdSP07o5y4/KHOUIUenLLZw08MJb9bQ94nNFG8cQYU7+v+SS0DHwytZi6Yqq7Xf3
SzBVelW6X0yO70bbyVupuVkYGc8HrjkFRD0pG4/C8AIGfXwfdf+d9bru/yYve8Lgeuvh9vHtVRUe
tcK1+E1efbs8VwNJxsLSKJJ9ldGnqS12BvT3HlpEhPXVSoN1UaabJ7/rC/Rz9CZ/Z0AG/65UuW4l
dJ56iXPntFV1IgfUvqt7jSzWT5S9R1bd/hAhRqlZySN9YsdrU8BwWLoaqOLvbIDUMvGv+ve9KkRl
GtgZf5dbfxFmF66HiPy2EKmzvDn60LKbphDA/Cll0j4AyACURUs3PvxyQV/HXZ522ad7xj+cu/RC
AGlXVcjhO8T0Wn5e/u/Ym7EHkBJglaOOl9Q6GOorP2YgCqxiiSfgBIRyy2xMB1tAlINhjrXV/S2n
P0ZBNEho7Hv5xIeZJvpq3AhTvf0jjPJnVuqAmLFB+aoyCZkPXctWJYHPpM71GMnjXQozgEW6/cdd
c409fKPmiqJMfC2MYx0mBQZgeKbR1WI2FSTM+zHk6oAH39lY+1Ju6jURcJYBDfAAkP8CnZLR1hzF
PgTLXyCXp/Ws3u71LPCsAr5TrFCuCdhCMvJFxqBhyPkyPjwpsxDpZbHv2OKbOeeQH2r8wgOTNRSF
fL7YLD0RMddSxyvTyd92Z0HXksVINTd50Gf+5H7cWAMkFFNG03A/1AOGzwaCWAeMlyYc5MJAPr07
dcygS7zWItjDruOSOJx3JY6t2efKkY4rjpgAQ/3bftTUwNdHg20BSQsglb1OpY8apVToHGgli+CL
jtynwcfvuGwLLbTRYJi1mEFR7QY583fwArzMDUErDyuGmuJMuApXNifJyI8VTtEiH7NY3OsJ3wj0
0PCNC1H+jNMhsYnEB8qN1skAEXR6OCeLCqoO+/AadINFea53R7VFLKG9bQ8ASB3Zo1oJSiXPwdAY
d9ZGDmXbfT+17AfFmd6Jd58wd2mEL7popt0pUVW735TBRKbThM4hiCT071vd/0kJeNFbPxQiIbCW
g85Va9rf+L7LPoDMFoYa08zEf8TkQGpUPIXqTCw4E2YzWPhfNrLV3D0Il5aDlpcqpO7ULczSlOk7
uNHP54y8skk3G1VJkADjvCREh77qS9nWe+Tmk1kqGl5HKahQe+a7Kuhz/ebFR+Gs9ZAyPrIHSSnT
pdbOYKc7ycC1EGSzHJL74dCZNhQPorsxawnoJsBB32XrNgIwh5CCn9lG0aTlv57zUWHjfaAzlNFE
3HPkNnWL3DQUSjIsSaRwVOyIF/FTmpn+Bpg7QofAjg9HWXihOMPrzF6M8FwEW0tpbeIAg3c9tHU7
ZVM0zBUbxB+V4JahTVJaDBTBZ1ITSGj1KfOgQGxhcGqAOFmX1vaXe4R0YKr7GH36vi7GSCaX68tI
iEzcKxSzSJEKweatpsVS6my0ya3hHTOBubd9NwJ8vtUssqpVzZgnOHAHb+AF27nD3LsaSzi27DzQ
bAbSHt+qjBCw/X917Z68tEYbysH8M4fOMqjT0z17fB5RoXgM1O3ajHTvANtsBAyuOFUUq8WRc8n7
SGK8Vl4cJNuJeBtOX4+8eBNjoPUDCjf8EVzoVg8dTI2LQxwxjZ2yJl9ZIctzBTMpjjhNTjOVVFC9
DayQb97XqS7/RYAVNGRyYHwAE1Qv2FxZHhZZ11FBFql4lGNCX5u+TkzBVGGoanOOqy5hBBH81Uwx
WPCrDFPn/IXwwDO4aEMCalH1fbAXF0902rTvxgM3cTVo8FeERDMGrMzXY2LIHDJvbrcPM6dXhzOQ
y+icT31rcS8bJPdPNyIFDJuI6H1AC1eim9ca7wUhS5ufp9LLkVZEs478aclLZ4WxgDJwuDeJIHza
Y85Sh+VuDa5M1wl72ttJ7bGLTcxJcRpb7RthYru1nbcb56FKbB/dXjk/DP/NFp0Ow3gIOpqdhv3P
p1C+A7HF2Rv3B44HNy6zO8zunkTWTRm2W1HX0JOmXt+7R903FGTo/5koJH+ri4Y1axbN6N4MFWHe
JHMKuSiFHLgRKYoCOXHU9L8EMx+jB3H2DLye14BKtIhiAALuEW05t6yixx5+5JA1F5b666js4PEx
aLUaQLSWj2wd24iBuff3E0hMifppEpCzZoInpwBXH8H37i240RKBC0fj+IL0hi/BYYWpxdAnDHQa
eBBy8mfSPYJ5PMEq+sqBuFmXZWwR1zN6cTgrfVyxpKUzJafFhLSymH2JLy5TNcDAD41OK3mL1zGA
mkCHEZbQOY650gMmxA0moBqCbpJoH197/KK3tfSVhyEPG8V0yKChKXKqq2JlqxF9ZP3DBDX/g1lP
iXZ5PuMXvnyrUeuFyQvj4/ZuFWpnU31HYjCfFqgF5Z/oa3oWcNMxnztNfgbfLL/B4J1bJTsAkIur
ifPO6XCVXNxnnjmL39+m0gY728gPB39CrVAEhXD79L/gmZ5rE+6NSdk87VgfsJzxXwWQA6XF1J5l
bXaqTS4Nh1HWYijKbPBwKXfIWRK/7euOZQu6Fk4lIbFtGPHG63ll7ElYXvv7csRf/R5pDSSESOc1
YRK1VByZtSIP7RrG3u8pyV4FhI+dpO/NXDDFcT1+vfuu9qzSwurA1c3HywW/DdjfiRV0CBx8Xd+R
QER6gdRc5iogN+iLWgQYuImxuDp3g1nR1MhXxJijJqwcCdPs3bIbheYIEUzqhlUQw5IFFbSbLmvX
v8cGeIyjj4ZtgXpz5euduGaUJtYeX6Tle2UrKrTk9p55zBIb71sIaweefiJh1UGUBAMrXjnGRBfR
KZ5WmaLhDxNXIw+qAs8LWdlKEhgQubOHOOf8YPfTCpsR0OXbdK+99Qaz5O4Vb0Lk+/msAsLCzCBh
oYTTGveblV6+YvNnpARi4uqkLOGz1BqXjZ4zo7B1VmEd1sZNhDE3exNjhiE7nOu47YoxYSwmHMwu
bCe+4jjvYm+kQKZII+dsLpYc3tOwcfCWqWA+nVcvUhhxyUT9FCWNVdSn/7QY4dWvsGmv/3aIInNu
umP4P4cACh23nr6/lkR4Fr2LyG8gQlbZX5sACnyUbYD3Z0e2e9k0uWnJl8aCI2M3iWBT4p71atyr
IOlQhFE7LHwdWu+fYO/TRhe330+56/AayC3HET80aPcOz6VMm7nedVVEOdlqJE2dw/1WpzqrL90G
qZO3/f71kO4xSdpaAREatQwBG3U1x1zjGGUimc3+CiyLPOOGKxlctN2EEQtpS2jihQwuX4xr059a
n+c4QsQ3t9b5e5i6dFK1Y1kzlX8fmQHvNDnVhZ832xnvIDOGIIVNK2+TjrPqLiwb4Vcmfa33h0z9
UzM4lmEqe/7wvPSZUbi9ctonYlbWzeMcjIrz3Gq7gtBtGIfBjyPE3vXJ6G2Wcl474LHtjQuxhIuQ
JDJe/5rn5MXdOiASFdlEKwUWUdDGHeQe2Db9rkLlXRracFFBLpC0KBBqzOI6/pBHMoIWIKXaOPgT
LMtiea40a/9R+dhT3XP48/1bDXmAhdfvdEYC/ubgx2oBlFlMie7VLsNk7hA4pyaoPVff8krdr8Wd
xRjz3Ltit7zLC8hRU7pngxIcVbpm1tV76NZwrdgp5T63uJKMXuOwj/0g9B1wUVjS00YlAsMPb58x
Y8IBSXrYRE8waNM75uqVpPPtLQVWyLqvi985sdItqyRhnGlwAiIzUwLuLtB8o6LM1z4p/xVVOdz3
GOKA5xjoHt6qNn/Qeq07lm2+m1VOejzpNIgSj+w89vab2vk6/etRcljaU0y4OskpsMBl+1xEQ82s
2vv2/2PMSNNvbRv09NnWa2wqbGPX0MY944lj/iOqdkhNJk5kRAVGjDObBubg2IrxOaGYTL8KYswT
HDHUS5bp6hFDl+0lxq3TMQGw3OxqyxMwUkVQF4dhcjo8TyKWwuwG5ye53v/RCyN4OUYFkwHyNgze
yVK4JmUvvbyZUTl+6PEdhXfT3cT0n9I/PhZ1Mo+waOysE/EFrtgOvQlroHslYjbD3CC+IUOO5D/j
M2m2ieyfNrxS8P3hFMQZhIJtvJBPMe5kBIOd41SRCKQ/PrKEnw8eH+I83cLxVWGVLPg5DlQUnmfv
6cFlJgybrpt14h4S8/ycL5mHg/Nu1ow+sMZp4jgp07EIpJ3GXlm8I+EacWsILFZzNJGHmnCCdQ3v
x9AlnEtLXC656Gy/FcOnYIDSZkGpJF+0HVxui9CCTXDk+eyV7tADm+ESTLRI3q6JW6F0J7lNXAUO
QbJdWVCs61W+JRf4J4CNR05UYCKcQXri/EA+GBzsWCMWrXAmNgUE7e5UFs+jGAMzAdkXConANJ+W
Ch4zUnpiz0YUPzjU6DlU0ADOf6W3fZFodwF36w/TZuMR1yeauD7VMsfmt4Gka8p1LMQMkFOzwAHZ
OB5gFDBWKmXODWnH5pYgB0MkvoNNBQdszeyvq10GwxRxmMa7KrcWg8H452oQL4IgZ5bx6maPpWfy
QO0ssgBj+4gHyFH08BRgr8JJzR0xec5T47tuPdERcFR3DpLjQnuLfyhc7lPsjXUwwuHNP3o5RXzS
RWZaHZgTZDME9TjU/XAYCAe5mUDb0N80iztoSPyUlVgldYYZUBZwRzObB2pUPJnACNbcXupw9hIs
6OGElgjqGgKd5rCFBdJ7Vb23U62HjFDSDNjwFJJI/TN/P/8kriIh2U3IPIOfpuP32f7DEKbet1cN
EckRYY3mQ8xPuObS/EpqtFD1ZY8bkQRpo/AaOv3iJrVUSlPig//4si7uffFC+WY3FlhukjMJlj1R
QJ1a8Ocfz2lsSywgGsC4R6TmRA1JxywjD8TP55rBNk6X4heemgpTM+tAmCVsSM1nFnVMkjm33SwC
AQZ+DhxZwLAIQZVCU80thxh82gLH81vofSPO1+pCC49Ntcc06WMZv5GCDdIjCr+RvxBqzGEqx6s2
nEr6Cxirixq4tX0lt1gy9Atgbe5tdh7D1Aw+C1EtzLgsoJzp7vYG6pJgX/RT1AzZ1RpAUBzA87gT
EFUPOKKeXFDL/Y/oJJmzMMpzPuZERh15z7Mz9aj0qpa/CTYP9UxcLlQvnU6NKzMobhFqp3yNuTm9
FzYtrv1kRbWiXCQsh0t2du+TIIX8V5nZUNBsErlF5aTHGF9wzmmKSmVIU+jfuSJG1G+fnJQs2C80
z5rFghR3g2zcBL8zo7WTPRF1BpQD6rAArmpUJhY1zEHeMrYGqbxugSbW789VMHcBVtDhaOCosnwg
wmf28CiNbZn4YY89bMYVUWiZJTXIjqMpBcaNE3WEAsdf7zamBHOcVAnehpHXLYRMHkIEYFXjFp4J
g3J5pspRvk7Ca4rvW5Vg+g+sf6I4OUj2SVnH+YUsoE1D3z2Ev3/+0TnbcqxiexoVGaLrCP4EAw2k
g+HyVNRQTV5/vUI/hPx9iexiUdgF4TMjs8//1bDxBd2OT4GyywokwCK4o6uNlEsiYbHyorRNQD9A
BTUdUeFxvHLrTDMpY+yvd4xAcyTwt28fqjZE8fkc/kj7a5u9RBmvY7iFIErdlcxCoZQJN7FbYMbw
uV7CBsTdZnVCfyJGDGDswWG8ilMGlPOPvmur8bR0cCnX4R8TbQPmKGMQg34HD4TQ9NunB3F0wAiC
hc5QfibMEqWQTSoG3/hzjEreD/FKevPpns54WmUXORfiECt8ue4KF2oEr6Q0xV7fuzvaVICCHvwo
7d3NcjboE3gnVup0RGeSvU8i+wjgD3Cz9jaT2AflyHqIE5fP05zU38L31A+jelnHFFegrOCqS7mt
h24rmjiFgIDGTKPg7WTd3OUb+5XhAdbUxU4jM0Cb7oOMebfHgHyf+X+AuiVJS2jUE1qw3LD9ExI5
kolzb4GGbSOtHxdSbpfXdBoDdAGd9fxkp+YMNjQGsgorHhTxjkmZAXhLbOO8IoHrKMCuDEM8C+6u
sh0WqG6EHhBf2ieCbM7PczZ4zBmY2cio2V8Zwr4F/H2rIo7Lnw/gF2Ky0uZ5pu3fUW08n4t1buJE
t3KEpW9HONdwhi/jeXFpX2U7lsmp2ON5Bfu/FlbrLfbd97nSDa4Uv/gR9QewbdXK5p1WjJYK9SO4
TgtRGnOAJ1+fVOBLAxCUVzUdEB81QQicIew5nW026alumcBJcY08mLNU1KcDn+4idiYSB1UuyzY2
RxOsV6UQiHD+gOMKOMgCwYQVQTlpYvUTpBkBG5RDtw5NZahtoBP6WAQ4f164Rn5fIL4n/BwfaM3u
RLBz4kiXRlRrOHS18ZDBe0f4IRHBFMUgRyhV8xy/nDuoZ1xiKEa2fL5zEl36E3F6spN+HgKeV3Z/
Bxm1pgzfJgAVSylyvxXEzudN3xOvsWF82h/gNj6qxn3pYNYOmvTxCCLfL6pfvd13zKwOXq52Ci+z
5HewsyfzNmMMIQ2VYnjOeqPGO+EJBz1Whm8ST4kb0/I3Q4Ufa0lcO3h8KOTSVizA+X9+CJbJBLGm
TjSpYX0gj3o6h+1emttQmINVpPPFu1+SJgU+l3TixI0RXFcqQ+aodGD8fOyPfGkUo5zkchEmhS4D
SjF81TTB3tgxZlMX0UmURYfol2wyRaMbsQTRqltg7jVCtRKxNPZP6x6N+JiH0EQ1XFZ2W2Cie7Qd
WDYObYFhZk2NmSYAxCA7T/J9/4SiBNfxzJZblB7d/N3hz2XaRYrnlh4DV3McDClchjnGFOgZGIDB
UTora6lYINJBdhIXF4TqcQSYj5I95s5itH0JzDFHTHcaa4DZlBTZu9zXVgJfs3UXvu+ioVizt3qn
nqwpsU2uERKzxVMxYJ4zFPrQ0izfz5NIKLAMKczpwysYvhtGYPcUOseJEafkXOmY715CuBuBuN39
yQLfoamnJQmvRo4HZOSCBxER74QjYitWhZaMhEtF/7vtnTA8aUP8PrDDa5P1Arbu9oIx+bx/P18y
NOTUlLTNUmP0hkB4qbDfEdMA/8zqq0+5etklEkIi6HPU1qE9IH3xjU+qzBxAr3ZbJILBHBQoLulq
p2oZ/Q3tHGUSKn/5b9LoA0QIzKxv0g4kIv1v3tXWL/7wiVNObm3KBf7VpUi09Lr410oAZ/nsZT0m
fK6Ky1nbCu6b/UgJw6VcOSSUa+9skd79WQKlQsUY0Ee1kUEtFOKCf4HHpjNxKOc8xH1SzZppsfwR
te5quVrOfx13a7+jh/Ul3M8+yv6YcynOxSeTfpSAl4P0d1KI2nN2kfsMjW18dXKPrwOeVXzosuFo
Xs0TCUuQq2PLa4Le5vobCFxMWclOVbLlKKth2rdfu4lq8eIwDPYQ4nQl0AaT08wkFmWTGDFZZwnc
vaBnZA5m73f30t7YKW8eVKlIs/7qOOOyBw68tYeiBg5effO4CLGydAMXMVukRGXMwJiWz4B/I0So
RSLEFpCEGSmj0PUEyZiGeyCmwYFCqEseMjdbcqZw+UQXdG4otrgQE5tiuSL40BBCONA+aseoRxHW
BV/xGeIUQqrEuXr2iK/9F9Ctc8OeiUj2nVwigS4t2v7Ic51r9D+8TDTIeOwSbKjLvxD8+J7pZrYb
BjXx0kvJoxjROzNxkYCI6WtSKfbOjuaoXhnc9B1T9I/0MHappy/Kzm1JVglpAKoAoGLPLGdLfMgB
RdsnZofAe3wbIS4spPT2l87EI2Z/9t4I3LIzslSEogkvi7s3T35iX4EdGpmMCDcK34ZUwScYWbhp
tQSJgZOVGPdzrsUGfpCp+P6/U1cawfuMN6J4o7eB1EXyqpkUp0Gun0TfS6bkyjJhImj5wCanPkQy
gED3cbkKLP7SbKZvf1CiXKda/A1/0weSxQ8DRAPIZ8oYACvfXOpPivRRThUsMZxyoUyQ1UC3yra2
A/e3T/TG3/xoyoJonX2ykW84cH1ZjDJczHuYp5+vWS2OveS+1+yPgvcQme/jpbrYK+sNV0bV3IcX
AKllINKZuPfgrrIxj58JH5+Ll1ocJqwRRFftfGk84uIOyqbGHaULS5FkzSCBixjtJ8SdO5I8jXEh
Wy4Lj8bFQdw+diqcSkq7p9uClasSG+ec1MleOfoBx3K923mahQEZ57WoxjYnBuoPguaFobeq31vz
gWy/5yk9srS4tVrXZWBuZzYaxRa2aRze9hwFDBn5uWPqmvpz8aRIqMAWDsRQOMaYW/gfNEX2nWkm
aOiXAlJ706TnsAB1Hk9YORh7SyMHujYopr2pCinVA98OandQJ8Dq9VxQ1fJ5hRR8mDc/QPYO6OdR
sskyFowUTi5yjRyWQJ7gQl39U5k1cdS5zA8IOMDJ8ZcGU13PgWHmw33LokNSUoe/zSi7i2kWlFrI
+H18M9BKCweWAokC6e1CZbh+18/CmDNUQiM1KNORmn9VEYdVA2s07HSYcCfloDx6LSeLj5KEz7oI
H0bRnBTmVGzGnz+URXI9/klyDcXwcwR7pSfB5QpLZTm1CD1JLR7vativ/3P3X0BIISDSHI6lOL1Y
mRl0CIyKv9uCU5S/pC8H1kLsjvZ/uEqSAXH7dFuydyA/bvG5t2IRHclJCQY+/aRYvr3U6T6tDcOb
R4YVZXoIQLDhVUR2jGeiebcnFDaTbuqKUtECVsY+bzFcO5e9o+SE7/B2fMxdcBvu/2A5EdzHZflO
azS/0mi22SfmnZr+iWx0LA9TBQul5DiFCv1/AQaQfDy5WJK3Ra/I0jdtK8JC5l1UJ4bLbHpBOGg3
IDydvCD5yaV5FLvM7MKVjenSTeYEtaDUm907mUC8G0+F4d8/U2HS8/W0iOZJ33CS/LLm6Qo1QZlf
E9WgPqRFT5tqbhIbxadJTn5lFce+M4b4eA7WcF9ZOgoJhltrfijmQ2kiLwkhu6/HDJ5twEiFL3rQ
21PUx2FBNdCZX9wlhGyU4xHrYTSDcvxHlV1tN7HVkBn0ioPgj8Rrlyk1OeOK9VIjIzlc/QprQ1y6
TJA4n767Swqdv+czB2qSBSj82npIbv2T0jhXumG9SXgsr/4/SgnzHjJGWpWK8s8n6xsNgfJFGjpL
47Zj67yDzRPUUhA4WdWjxbGbZ5rYNyxJef1G5TKSPfQnQ/VrWJZLDUyjfnin6zdyIAsBMLURFRXJ
0Wn1HNiWPDJoPg/0C8AYWDsH/WZ2A67nVCfB8wYxEnH4blMKPYZsgGuxNAjndKR6RxazLzYQJ8oo
Svp7m68WDvcvFvJ2JRvNEdzmJgF4tetN0b6gU7o966kCIri1uQOKOy1M6aXgC5R+lsesTpi1F5yY
DPI6WPj91huRSGhALdj+yXngf1gY64m+dJ1GFli1BXcoue/H1AZJ+qvlxZIUaDvn9fOD6GIdDKE/
HBf/tnIJWuebJ/LFIrh6E6EmP/mWZkxpZNOUs7fDpHuKBS6D6iJcf7K5AeFT011GagZn+/wRS2+c
g4LXV+Z78WZBLZG5uc0MS+6pUGvHb91jh9sYB8/+m0BDKQrFKh0PkMG4vMOiMOthr8EeHkMwasUL
ayNEq4KEk3QJ2edoDKffuG+nCIOb1QCWWOAvefjzM9zxwyTXe6DUmTkW/xSYnoyNYwpbiCI+/pB4
P3VVb520j5geywwKJDHsS8SQOjzcaiaouVWv90QQoitAD24Pgle1XRV3H2U82LmaU34IRZhrRsE6
FMqaruxVCQ4ieN2mK5zKkCPPHgUO2sm6qmCvKzakR14Ifa0IaqCTATALy0eECt5vfz1MG58OO+IL
2tZ14Fl+KCo4wZcn5xOLOzBbXrH/3DrVvMV/vHJHEdn9Ec5cdh160Yz1e+vtTssg9qhuwixJuQ/B
+A6kviHMHQpWcbGM04otMj8wRuoB/fv7F2u/22oqWfgVjSTJRREPcQVgw1QpTkpAKnLAki4G0tuH
eBzV5+Ck9zBA8SZ1SQr8UiQ6pmBl9pmLW3vJ24xpmYRIRdoeEO0XY3/FUu19bYe047ePVlNbpZy7
bmeoEoXhwCdGN2gsoG3XTUQqGn9soRPhSIDEEA1Rnj89d2vTyiOtpjhtC2e6EtKUNxhTNM7VlkUW
87btrQnrbbKcXwrj92gY57cO12dMAr3tRTWb3PPQ2k+RSiSKNykvuzBHVLsaF3mITt4yXOMZNx4a
VV26ig4Fuwc+GWXAXnILF8K4xju0o8a+QJiwt+Hnlnn80PMxaxDhdU9wJUQ+cEDQiY9RJoEhBU13
PD5TvWXaC8QFgtpbX0GhjDvNA3mQI91BMHEqBxKjDepDXumYfTmEA03CWx0/JfC3186Y5P++sfng
u+DXZ5q6YpD3u+aeIgWddt4/SB4XDiJHmbzNoqJktUGofxixtUou71sTiVGf68lJJ9MCn4AQeCvU
S+G+SNg7H7hyPlS0/LraRBM1HjGn0AgR4e0XLqHz1AG50i25xJSTlxpIgCOZapLAyrJBI09M009j
rpeOgJ186Gp6FP/gfmZeR3su44ifQzl5BDfIn5bz4+6FX3TyPCamxQaKRngMNUuFvMv6tv0HKDwd
yN3TcCXgWehz6Kcg8RNj+ov85UcAB3UtZ3hNkyB6duf8vSSC0pWkv4N5SBpLdmjo/Bth4/Kfeqx6
yAkqaSLcMNuOutYnRqSy2QRcZaEkOuQLA1P9bT0q9LbAKu6QnmeLUA/e5oI19VYp4L6W9JnC08bQ
IQOP3JBf5E7W+WCV5MbsS3n4iqGsycbQleDUAVjVkMORQilMYI4LqO31HVnMD6ac6mMc1DT7ikUd
U8Qg6QrDPDSUIhQ533LXPkYbZtKYCyYwmtqZe+g5QOATBaHMC4HTNQ+2RgamglWNxHHm5oRI75nR
oG7QvZgcOj6SrlYYUyoU4/ej5LAPhtDszouS8XkRpJpflfo6xYS9FxBYZfT1/OLBKsFLDioO/T2+
3L+A06jKaRCY5wzRR++I37MhX4yaiTFTRBJVVgMzgLRxjZOwG5DBXXuPgKK/v7BafFM5Qev3PzYv
24DrdfQrpiqCaajztH+E/fqitJNI7XyzGsoVjo96Vt8vGg1B2Z6lWiwU99ZdxwvGQ6QnRtuAKj6Q
kJSzU8DjKC5JeFjhgkaASFGnQWpflquWXwISzOtSaCbSdSDh9U8wOPMvW3Lfx3U/6Cyih7BSIZCR
qy/FFqy6h8A7FjHbkhsdXl1HmvBzVyqiTTheBk5B0enIkE0eUStMi8Ffo5+sRzjpArLZ9MdV/PS4
kRrZn5hLPGGEkuWgwriMRN24t7hcddI5FqzncDSOczJ7JpEJeoulNfE2Obzqp8xjfcevTMTXUu3q
J5rreqEBGWun3rC5YUVQNUZe+AZlfgpY3mEynQAvrI5c0Ct6/QQfVgIUIm1CJwZBdBdXmrorF0vA
R/6QPaGx99RjPbYQWiXmOI6VfeUJ1AADd+s9JGIHd6ivaWjSncNGsu9JkbdzHqTSiEINqenXYY0T
j/19RWyXHfrrqgZ8eljSPmKukwq5gZ9k7JQeYghfcXRBQ62saaHah2AorXBDvJsZlZGDxrmeeE6+
Yay71UyXH2x5quZAFemb925cDWokErPIwslOc7vJHbgSoCZjUIITFPUzL1MIsnncX2oBI970pSJj
wpCwRXOpozhUX+lQ5EVCDdt9Abbd3IW/VDWk1zQaNNQ/kbKDblEtODtpNSj8Yisk9UpLxBiKYs4x
1Cz2S5oadPa7/44VX7gXVUDZPhaBN4qSbOXOnlgR8cSJLuBeoLTJmMcRt3PuP4flWCI4sts7FsGc
AN1yOrMQTJVzC1n3YCWUDaAPRDC4o+yCS5vrfBxSqoprHlzZ453kdITavSBxl6bVvWxa0jpGpiB7
2jCGfoYxnN05c7+smTkFd0O711T5uGkE0pjyubWi2uoB49P88b9WibW3CKqolv5Ol0zBYKwHx2mP
fjLos7cSu7FxNpPurE3uPEfNybnKbqf4JtnBSlm+J2joIULn+3UCo87btwt6WADWWGHLX2iv3OIj
pGhZgWNxZINqQEVcgokmjdzjYJ8sz28dn8e2sLn/wubGsTKxrtnEjumZ/sGLYBJhVHE2xDkfYFHs
bMdC8KowR0sf/K8ANstq7/PYyCnDhRxG1mIBzFMatb9ZUdf7Qi+M8u3yXQksaYhovyDZ/hCLsud9
IUH4EyUZ7SSVLSXLH3+X05Z7Qw+U5qANm9ZHkOIczdCKGERAQz/U4vmisYSm5NLNjRuHXQqAyhTV
zPNXGlWqQmpEKvowszsUHjTw/4ZhIOUUy7jwuXfOgZOZiswUHtP50geIEXHj4axVPrM6C5Wpkfvl
g2BGJE4505fFrHkhdbYqTWdaUVRYzCHKF7ZyoIyAXh772EHT7TstDJtc/WzXFwq8VHOXwIl1bs7r
5ix35CetjiEV+AiZCw79zH9O9C1f1eHJBnXy1ecEpstyudoXB8wTivjfezqGvqknOCkv1GNT2DZk
RlaoyI2Zp8JKSOVlJN6jyLj15OocWj4JogGNLCGoToOLZsXc7R25wONpEjlSkjxck9ehZXDFeRKA
iOONsrPPGqmcP+eCsnpoECwKV2B+2zeZRj1S8kHChz8hCHfb201lD+WvHcUYdyRrSEiP1OQbMhdV
yZuDOIeYs5hYu9mDCycEYW9/hzMBi+qJ+IkGrObmHgLuj4fHlXiEmWCO4AunUYi1U5G/7UImMtwp
lDzO+jjcBEjzopw0G/Ml32mWDRAahJ/we7Jdfy3qTxw04zHH89DocncxYyp0jChgIAenw3uFuh1X
c9QR00zSgToBVlLbq1o1uqrZ2VXax5qwup30yTEjK2a6wzcUtwhHALacQilOC02wIoIoxKUX1iGR
arPsFfBWG4EZjM9RseK6FTg3RtIosQkj+YIyYnf/eGTLKE3KB9FOs/hJHbFw+w3CG+XVaET3GKR2
/pSOFRzBkKN2iMzPa8Wygn05AGRCIby5asHAwSNn2qdjPg4SKT21yzNH9pGffgyDWAFdABnm76KD
d8ITqTaMUrX6go1SKw/fwBEmwkL5X3hxbFYnogxMQLOC8/evIUCZCeNflUUTT7glkmLhrR7ndkGg
S9MvvKWuw96O+oOJmDSimgC5NA3+DjsD/agP+gIz7rabKHHQl+4shMKjqTC1iJ+YrhMljVYnyi/C
irrSh8XQop5Y5Bc6ACwKuhHYS8iyZvT7xJgp65v13U8zpWlrLdovhQpWiRbUB45h4h2ciaAx6Y77
ZUaDu/Jmoa/e1tzsnI205KW+z5K3F/TeHoLLLp/KsERM/4sauBZB6dMisRdrUGMkZhKudORM5Lvw
5zMt5qGPuTjBh2Zjv0vtFsFR9+XyU/s8ccduSqyP8ivMXBZXs4LMMdQ62jnWZg3H3TRoG098p6Lz
Xj262I0xt2Z6zNvuCFFhUKFwT3ct+XQ0FIIDQjgzwt35LaDv9xkI8sHV5zEVaxCTABRpw9O82eC9
MLhzpxeBTKMT3S71Nq9C72qBzYavJvS68bfNeVX/SxVC93nugehhu0V0SGCdF1CDu6TFrN13vm4Q
+bahXPdCplmUKrZTyc8IbcYBHrm5YQm+GLGot1WhBJKwuWxDzeEcL2tq5lZ5tGzY9pyyvzmOUm+i
ws9ckOIw7MMx3zo4wWrXr47Q83DHpss1PKdJkwZMYD/4th3f+vxT//ZEMMCsoN5bCI1EmD9VFY4/
9ymM/69nvUAN9SrjkAH0I5ksQOVbYxf9eveVn4HIadOLYHF4RxHbtpOW4eGzo1toDlJF4/JpAH79
+hdrbS5c7iiFo4aMohJFqMJNR1RgtKBP/KbmZhCLQkC0lyUeV/axKfurf2QTdKwGp76c6GDvvPUr
weJSHiqXIv3Dpc2J2lFPj6H9DaLlaF1rDFaYWM+BHn5MlOPSfH2S32HnokQT6DrUPE5m5hfgFpwf
jJCiJorb56RIA4i+29GDcfgSROE98V0LJieh8nk5HPQwHrLKTRKtvYSp1xHHQzdhsZKpFqFpOntF
r8A2t1PcnVZExj7GaYv+5IyQ2iJab3tCVNLNZsOKN5Ss5Lc/Et/sQdshr9gQQ21Cmb1addZR/SRg
e0ajAJc3KWMBFrWy4frr+VlqWrKkomH4x5TqM0V4RiDSxh818F03J8rE8cw48ZdQTYLDI0QtGpON
3peMqtvYiyYDA+dBP+7yPXSzck/IC8qo/uN7aamXxlwnay9ijEQ+k1VG34eI32yYifiLBkjI1pBV
oWbTBrGmvvOx5uqj7fcO+LLZeoTIji0jXmtNfOmfiHD5/TpHJNHQo0vAW1UEzfkbZsWnkrcvK0vM
oNTKA0UtnG6mL10qp4sXcpffKVRyQcfq0jyGeKHhtglqEOzENSHzCy94JArLLWBVCPS0/X07HDeG
/L8poj15YwgC+WVcsMQo7kQebZH+wELu4Vxihkqw6g/uE6RrJF5CEBBCSeHT/D31ABSNyWxvMxD0
Oc3d0McdXTUlzear+/gO5W40qwPJTpaTFrknN0yxG+19FjAfXK/7cIouvH8DJLdF9HiQv/ZHkGbH
ItC+dwexGYp9FpjXl52THKFDkZ8ADEPXSzALRwHqeqTf2LmEBFehO7wf6UFB63x7t1erP7OW3xui
oiDhqy8bDn704QZRBqJwYLDfdT2oDrgTZ80nfjSEhn+VjzDQlK4fu9R0iQVNNfC3VacMYz2m1JKX
/v7cdd1Q0gY+QH57Qg2d56efFzCgs7emkExZLcj3iU22jSx4Qf5VJnDF+aR0VCzPP/qTpw7M5w+a
rMY5RxbN0SgoW7J2rNGkUufhNqPv5cuQThItGJLvNFSRGLThPqjLqP6K1SgLauxus04lgU7xQDd2
Qm8yjNRAhw/SXMn/3MUkGptDD58wQTZSUgsXvmSB4PV6OBfdMHXPtP9uuXSVpAQKgbb7zc9Gr2XW
rndlUQRQWRc17UwKw7+hLSbZCNXgJXz7msQbgoHR4ga+7EP4C4hyGuQEkEsIf31ZMMgQjL2Qak1A
+0AQK7+7Mxgcm+Ezf5WtY4YcLbsz6F77aTgziPHNzRIMFivnKpzrA2mFIkJ4+isx4da7EU9UbUzn
RvyTvbi/eyPw/Jdd6rPoQkocBsf9imi3OuwHfYVBlbZ3104KiSM6hY5UQmTgXWUIvCRdR1jSLc4b
932k9kF9enc+Hy+9Ao2CRapbxazxKWy1E3E3tuI8naNaNOm8qG5fo0nUFlItv7DFpTBxO32ZPuLg
+GZRKXx9EWViIYZGB0pDjK8+tt9vNfAqr1Y5ORiWVULROHHtr33zVOEVZbq1wdJKKCrZ5mvyLkCO
pnDW2Fh1KbxoELj8E3Uj0L11opHVzBvbiu0r/hMhzOPe5nqapKp1AuoWxi1kxuNgcG4jsGWhKXJy
SklcEqKboxeCzyZRsXpTfZivaN/9HnIABR3yxJXEFi7fDus+N0NjHshOIAjBkIhpeJzfPZnGSfw+
EG48r7PpBCLbXw6ICNiws+BJfZD8tFV4I/CGj8U2ozTUdHhvL7KkVIwYMQkh84TEOmJbuST/R6dU
y3xZcZKi8SDScScEHIXBQeZPAUifAO9qmTsrUYgpNLvZnZTnKrfhWE2s/2cY6qL1mlhW3GzYYjDo
erS0oI/cqHnp6MpaO2LbKHiRuLgi+DuUfzDI587i0MXU6clHjvZos4G9VsSVDDnUBRjjB9DyeObA
KEdVNdJnqV8kDa0Zk7uuAhYNN3FkhqkeFxBze1zNAbQmXuod7X3RM1yiusyFc3cmF5SRQP6pSvG9
xxUZdQealP5pfzJKZK1mbEmmsTe0sEK28I5Se6s3ljL3Vc0M7hihqF0HS4W4wlwFzZL96B6+KBst
8H0pN7/CxTB3gnXVPk2GkVxFcRUoW8Ur6Bh8FJQR3W9mJwcCw5/5Ffu4UvwUXJRsmzr2O/A6rNZz
0P3IM23hX3paCctirZkiMdHHS4v7kgHC5CazI1E0zClnr+BKUA0n/56JBct3bDBS5B9ApYJeKSDM
ssbb4QPmPDlnj+sJkj95+2BlFmYGdqCMFPlEzWzKFDQiY4P8dpFtDV+PbxViS8GyIxu2zTonTLv1
mkn/RpAzONfBVRghi09lvUV5+AeGmNsoo4QWvLs9Er3ceWl1+CkKfxcwkXRcW8ze+75TLAlXHOHw
3ELLpDee15VEVAwEdfRrhO8UkIpfNP8htQoFJPBdQZxEwpw9h8GwVqOlpIen6jSDtCQHzr8/3fkV
kuKfws5YVyUi+7xy5XK/JC/+60+3wqgQ+ZbfYI4UGY2xVThVHShXpfA0FqHelG+nldp6r67zywZX
LjWY5jGmPgIXsRjaV6xYvcCGBUMMIzqb0FSuucCE9A71l55ki0Xc4hIOiP0RYggpiSf0ZKKoNXt/
DFPUD7GxlQ6+9tQyNgqw4+HG2YEH7TJ0AVUHCij8s83G2EVyAK6/UUpukZUzLaUQ36qyESWZuidI
I+svmv214H+YyN5rmnUpamAo6MJpYMv42d2MopYdkvm2+XDnfhMI2wJVHl0HBjsaWXknAnTxNIOg
7r4BDUS8ftmcs3IUOOXRDA57dd9YeaNY05xwMBLsh5PlvIPQg3XDiLTvLb0IXstYGUhG4eFF0+ey
Xuvtpeg6D3pzg/tDP07d5dVoWbsHY4PE/sLzC09A+SxUakSaojOy03WAtYwl4HV6uh/hxjfEwN9P
H+TM/idCqgTFOE/1B04TF8ACJdYLLCnNHPnE9rA9l+0WDyZjR16X2qPGF4bPN2UD2+C5oRBLD1ru
JFafvQ1irY8o9SDxZC9Qqc0x8dFrLQuwZPJLKOxKLOFtclBr2PR7P3y1XN/nK4IuSwIeif2hKjbT
VHU1XxM6yhDGBlcRsTXGdRq+3q4MGt2KdfKucGEFwlBWrn1gDykDJyrV2SKBRKGtZZvVp5a5pRM+
QoApEY0KpWQbPkomsnE3NZfLb/R5goBcgeFSpf5udddjwKTFyDjz07b6OAqk0WfB3rfX2RKEYzKV
dwGXGHIYxIeMTlshhQGaB1Qzs+HLX3hEZkWzWKT27RNhtJtpqy/xftJRrNEowvasBlZz7OGmJeFj
fZF91P6L4CVUnvLIvQVX8ArDh9JlmDwFuMtIanaO2yOeaLeKUEA/llZVUy68JcNsElWTGTUKVXjw
f0cXrSYnFBq7dVH4i/r6IqRyJgUXfB0k+P21dbWc7XRymywTdkPKAGTe0xLI7moBjbWEQWNK2CLg
Bk7pYx5FUQOLMfwtOSY9Y+TQIebm5MwVMcmx7e5P2WDnbsSvezApKhUiSB50BP7WbVobQCYCXpS7
wEXogKtsodr18yipYTsammqlT+ChwGMk+w3ZHlbkprViK8nwehiLIiP3gJ0BnVU6pOAZPBfjUj1X
f20k0qIaErX2/7iRKh3eF+VHPh+hs/ZG9VdgQLrInXbrZUa5pz4ImPl2J8685iVxWXmarRgpi/iM
tEfZOC5MbGbBXDsfzRqxf7U7KQNAG5ONRG3KGNZ9mmCFDZ38Nktf1Afbfdmt/oDyrsZlPhYmYdJm
OAhsVA3YKh9HCB/pMlQ329V+FiUgR7txFVVVHfQHg+uASui+jTJuJjCaBNaiVs+od+iXx4PgDgSz
n0gQTOyaE60w1bqZ7jwEy7PxStxBiM2Vzt8vm7aFKiWJODITzcMoCQRSeugeGQLKU61EwMzOcOtd
D/IJZEctExB3Iyz2s7veuH8t6G94CSTww4wHdfetAPiVJvDSxAc3pcV9aHpcrdqQiNvJ2iIUtefC
y5z2HQak1r9dsTYIL4RzB3wu0WMCa4Dg0b2f9jX9CliHIjJ2vlrDI3iJ8EFB/H3/GuFOPiaNpJKs
Zhhmo05+O6kX1EMRPE7fKn4pnodRlGTbHlsHOCUzcLXNrSDJOk8RrMGjUDK/NOUe/AOWDzYjI2JV
EkfmPsFbiPIH+xWU9OOphhCS7cA9LImhNGHFLlNkXkv7XgKtrWwBk3+HeOZvWc9OVgaGTxPw7h8o
K801OcAPav6DgmtArxGR1NecY2EZrYRqmpvUNqe6O9D09IuhyrqkdicAUEDwnWAcZEwE/dlk7+Dq
+GrjC+SQSWPEFG0rZUW9n2mTlEyERQnNfpD601S3AcY3n+Kr0QGVK2W5XBM2UB8mfXa3XE2fWGy3
LNVc4VJQXwCf2VElN1UnE88RtBygVJnBAvfxYQcs9a+BFf9AZc1tH1IX5/Wmj9/97ArJyUerXCdB
Hcbg4IdeXEGNWF20AFztJRg1BAf8jAI8BIrDEl5k9wdRnqe8Zif5acRifua2tOqyiRUW6viHVtY0
wZzqV1Gs/PP6ddWgKRM4fpnBahair47g1vO5KOA7ZDHNDxcYxNohNoIwbmjtfcB7xQeXCgd9JEHO
0jovToXkKaliZ7hUQNF6t3HXkzq8JqkxZogoSvNsk2pgTeuK0SID6XLUB1kX6NkZQdNVhrj25Uxx
6WtEaI9UVU5VkwefDjYe5Cf6e5pNGy7H7Pi6FiaKW6zTmR/xdHNcjrGYZfk8X16O2hdMPvCaXrjc
uKD59eNQZEF8zhq0rm3BY4Bxi36+dDDFuEPTjWyh9ZNDIsu8zbXDEjNd0YbFs2tIvIncU8B5Fu6z
MkHWQlqyh5xc6jQ3Im6mQC8MyewIHFtufaZ5/A1MGVnbqoMrZkH4QxvYD0Z0MAIqGfTHzbcPXEQL
QA4Q95K6ku5TK6sZQL24XUx3ZdwO3P+m0WagRjNwesdfF3dIEoHs/tNIiAU0sAyHl53jv/3wytlr
q1Hecg0/hF0Xc0vkvg2ZEeHY6w1UWwlEsqIc/2m9QPjku+BWqqpq0AGRHN5/s2v6x0k5Px4AYyW1
HkOgWJRWpCqD9j56PAFIcEKz3mxVYsWYHR+FC8NMpgaLOEYfZDnXc7gjP+nXKj6sL/rlgeu53zET
RiLOjz3wzWYCL5mf7juzUhuNNUwi68EeICGX36H2kUdUJzpc9Hr111K2aclKMU/xEJPU+amY1EfR
k7t0Bno2Hxk8c63znf9qhQ/sQZ155tafLApUvIr82z9337accD2BCcVwky7idCFLjzeVxH3p5nYV
IFlg5jlVFOgxOtF39oKXxnOm+qSdsBy6qJvuMBRMp7o1EXt8r6IKRv4kLkrsEqv0TjqERriwVbxH
5u78Du7fj7HxV/ocxcDkYf8B0bjkqf7mRe/PnmYgvJAMyCfBDkTTKVp1/k5Z6abwpz7L3n7W5Sji
d3hrn0mUlhFCYM+39RPS8GREWBo8ORGfHOJUHqVaLBimN4Q3oSs++sPz86ywr4EDI4f2JKzyeiOH
0pZitIS8xTXV9gFu5mCT5ViqxpugJHdPOA6HZe0YfNdEyUPuvXHBiLz0L8xZxES9467lCPSjGgOu
3Po1RaSQerGav4p2RrbDR7IydZY0mnSrtnCVI3DuOZCyl1JiD+DFom4pA6z2XMOMHy+nDtk2fZI5
+B7lUH6j0eP0n+xusWD4YI1H62SXEhhituIWdIG1Ruz64zNmdgsIrEo69jPgj07dg2j6m/6WLalx
KncEm9OoN81ZcHSXA306R9jf+DiTi5uByP+sKWUiLDOa3wmstYzkZbsKD9RTv9jseTtlmSzH4hrf
Tj1BdXtHMetG0rZ5RFr/BNppM+iqbWFYg5K9kFJYLkCJ5wo46g+OdPEJH3COEubZkSp5hHJBLeBe
t/YWFRMGpzt+YPVer+C1aYUHYVuFsR5MT3vtY7Yj6aXaMjlllp86pnPxGDyHGLLSpfU2Rr1eE95s
cMS5fcxiscb0hZ05r9I/Txg6wQuPrWbSee63TmyXkcPaWz/EOxqQ/dilSfZO+wJZggkX17zk1Klr
nUVKmDJNDHW9qz9QUEA7rXOT1QFY/+LgARr6PBE8yLM/ngWHk1ubMPVSqKGhofKJ1+H0g+QVNb0u
SYKVB5FGy4BIB26qTdXsGE2su0q1N4mA6kkP10uI2tLqSEop0NE4IMSFGduTmovhUcgf3XwDlxK1
YqhxmHSgqRrXCrEHOx+qQ4L0FfUD2ICPoegwpa6E/ffsg4ZD0hPNU9xQxYPRny+2dOdHnonGroEH
Ze96ESzezMb6MfGEKD3yXkzYfOExL83NNBIgkh3CVFMvujcBoJDVyqM5JMc/5I72vsDP4V5rgwjG
XVc79f5nzMnD6fi9aWwzjTCr3wXDi3xQ5HRzrgBSwTgKdd4oUsK9G0yAinjRMDTtn31wLvrrRIvY
u0ry+VG/jr/OJF93cWjPEuOrF3+uQBIlpAV+tddvt020FZPR5pPw4Ghwc8h2w6weRGiJTtJumniE
YLky0bQoE4HGq91XJ9U6jGr7paZP9plCYfNpUATT/TKL+Q97wFHkKHRj4MHLoCCU36YeUGJFkfRJ
21aoxOBZxOI92sH4/6/yqR7qlraLjhYyKcIUhnN6SD6UR//TM/dLMKFO0eKOHZg4HwF5ZmmzQ7z4
OgQ86pZ8nUVs3a8zArN/RK8/j34R7ZXDLJDrVUoIpKC8bbL3t4ZtSXvhm0FQj00TKswGmAefamq/
IgCcbazYkM421AKB5102M1dJ/1/kHqpVY82fKJz76nka2O9wLsvK5/taJ4cgmEmEmPqwFTQh1uGN
eHt8rqwo+JMrrTdo1CqlrHaN77tGmEP+vDOlDNedW5sA2V2WYec9tsghI44wHpJvgkwZ44yFTN6v
SZfJWTfBEcF2o/nvPutL13Km/8Yvd4U7BL45y+uLJM0ZSNHSaG3GgCKN2GGMa8ubvtJmfCH2L6M1
RQFPeeDCmoii7plkKdo10HzBUshOSIccURAwUlYuefsBjKxQ1c0CEauPct/J2Do/zUnKFjL1zPrV
O9YkOmRfZ49RXOHNRc2FezgYrvDVDHQK1A3EhK68z3TWJApboC1+/qCoHJuRzeD0YIiEr0LcyGN8
uQPVjMyBUw+lXDeN6Aj4qZAI8oo71K53njBqy9FtGinDLifdd/a9vtD/DG7ufjNrWPjPXuyvf1qA
gkkjWPn0Mt2e37sRTWiAaoDCOXgWD8cEgF4zPCkgUiirbRHLFiqn6YAZX8rHV8T9eyUYPokyvJ2B
MRoFhl6Xo6d8+Ry8enermtFByVfexH0JskDCRcWhJuxo71kmlyjO0+o4691fbl3gOtLkXz97F/BX
b5MTJ60zocuUxVd9bAE4SP2xgntlpVMyHbHObXNMGXjsz4+53u0rJ5QQjj5q5JDiKs3wBTHG0UKn
tLSjAqyS8DiK7fY93zuRNw/+ghqKEoWxwqxDL9nFgzMhqrMuHSZdcYbfysITLyfy98xm73bY1A1/
uNA7zp71rMQ11No0HMzAhT8ofjG6PCIIbBPIuy5mP37viXvocNvJ+65zEd0gDw4Z3TCkx9ddwVtH
P/CXC1b8ptbyqw8i6/b6dEfEueYJYLctZwk1NOMCiQFHCmz/YkjyJYKs69WbrmU7jNT8DjZjpwpr
c6VPuxmcfPKo9+3RaWW1BUSfD2Dpb7JPmCdcO9mLSvqwiGn+nz1RqngaGMvP4OHLoi5BOK95+vig
6dZLRlZYm0xERGvsouZA/ncd3H0m8QcYeUtsGIOjhVBV2mqpleh63VfSmvOH1NWQYwM6l6VnB3tP
0qXV6qO5kX0X7gULbUgBuG4LNMXgZsffGpd8kKMGWFofGzkgg25/G8PwCMQlIPE4Y3i9WS+s7rGN
ehC+v1wPrgD48w6vbIWWloulnfHTnlpnqfhQh3G1YLKeRTgWU+m7FWsXiDXWOcf0CGlUnPvyEv4A
zq80rP4L/aSKXhQoTtSGvwvp1o2VNbhdspxw0/hsm8M2b3cFPOPgoyv0VHshIddeZWw4TcZ7MMIQ
bmin9kTCWvW4uQ+gJ2dUkPJR73fyPihmJrgrSUnr+8JAkjk8NlDOhyqdnllh1J6H3oYVX0kW69qI
1C2UU+4598u6G66vYRRve7lz96IoLH+Ze3hhDS0s+CurFaEtmbZoi1D4dTArQCQp0YCRjwsbdX4u
PhJ0xlRS21Dqp7v58VPBp083vrt0EFrvhDGE817kUy+oR8NVrEdLPsPZ/820oYsL8zeuZwsJoSNm
r4rWytjjNExlOIGjdrZsoLEBFUe7vwvBZjqZ+HXeyya7EH8e8yP0t+imGzZdUZr7H0MlWQqDmG0Q
YpWR0W6/L79caQDlhsFDyoJ7tss+5QLwmDKEPEduC4RjBlp1W2fCIEMOPPtGRZJvOim4GI51FHTa
or6F9kgA0JJp+jw29Qgx/r9gfv01b2M5GmZIgr/cXN4qspipqyt6RLnnpZhMxKIt0sM4HTvRwvR9
/kiV3Phy3eA5sxZ0u4QQc1QkM7fDcQzRQ+bLPmc4TYrPsJ7+/HtOqQB/pr5KGVf4Rj7uG6AQYU/A
KWGf0KnHJKjQ25xA+R9wMBtzrQ53DUPwdK1TO4cm9F3kyNDoa7LblVYYBQk5EQx2iNIitFHIzS4O
7vy/jJS7/39ihC/KSutOXjwo1tiUacAnaXsCSxrd7j8cSnYSAneKqVd0oMb1LsBsLLbXyvAErua2
kba2jUSOH1OZwY9E1jutq7DnFyA2oFPpiadySOJ15zJUZmpunSTcRl5uU+mcw6UIWPZJdxJaV8Uk
doBgqvyhaUZCnF8qkLnXSvcapZNbD2Pcc6GEyMT3PezCOzphN5UdpsHtOU6mj6BxDjmnsujgOkhx
oiEfGRuGUdGKqjyNLQhAjNFrgtIuxiMXWoC3CLQ2kCgRXzszEbu9C3K5KdTW6j1cIiiUDvRNWlsm
fAW60xELWumoFKb9WwLHO6Cw1jhOMvnLnO34/78UHlc2GpuWjej1Efl7sHpFW2lC8eMlb/bkc50o
tAKjC0qhvEETxJFDv5drMl2+Q07tFDAQ/1Ib8oGMtb9RQcrqjhROzRguU10r2nVjFuKdRAn3thru
B+3XJG3aaf32gkTO64vXX3AsQyK+rh446GQTyFQGfJGOGOo8J2kiGRdDt+0zNsIqvDnEWLWCQV4X
dYNQ6fkf+aLQI6dGuxy1OcIdLB+GYSG1SJ8fw/LtsnKjpdYcrw5DmGMdgRRlW5r3wJ//UN64boAw
E1AkSrgkHsji++TdQ1+Ay4gt2T7uGZtdVdPCtZ42Nfck/Mmci9UQ2UNNU48fXGhLEbTNe5qCUI/B
MxO+j/b3DPFkjEz9RGDacRC0Gms9Amg2R8yLOP4xHMfAXnVR1E6HFQ05yy4yii5SQ0N87GsWF889
pOfmrkvMzM/MnD6kds0vzwkVL8aFMnZAmbxU4E3wGp/zEfejCBl18TTrXRp3toLTNZkgfycVg1W2
g44ddIdDX34YgklTPncXdD7eds09onPixXWKIjBu6Wsp/uOKXbMxiuRDXENRUMkmMcnjlnbiG35/
PGO30C5a9oIt0hPkf6o9xyEU1HqKjX/qPQ7knEIkRePa/kLEW7gmQfw2SXHgteYQuzRx0nU5sONG
ilYkP+KRcpfDx1lt/6gx+IxeDc/uHujz/Jg5TiuflVNM0ONDkXfr2ZESXltVRcbJULn4wPC/OTsX
up2kBqV3KaZrOaaBLO0cjetVYZPjtve9vNAzg/mfOpuoT46pKq8zHN0DnoQRlE1ifKnU4LWZmKhq
Y01HzH7Es1pN83KYqjv1S2RDMHkmTVDyYmcTOjLGar3tGdrPpLCXD841GjReZoyKttEXCi/thqZZ
Vjz/BybLXO2axJa2g2lE7nE5s75KRmOrzbWO+VO3PBxlZh6XjKWKO4pPxwa6P2aove+hlBOt9XDX
MYbtcJvYVisemQa7NpuPCyOIciEZxX40qyBo9jJG9AMCroXDKdVs86zq7/xayDywOd4FY2JhxRKY
XPFFiXQEGsyAFs+WHJGFib86JJbjqgyVw96FQ0NMAzQwN+nvq9tN0rcBMLdxuiAaWBsJ78nlQxkS
EE7OSIA9ioT0L+bJ7/nM5z79LCnLtCGryq8DO3I+Hfihv0EV/ki8SqhM/9HM8ymef3gnBO3z+jj8
/u4FtEoobjO7jTmTrLg4JjtfdNKgjVXf0ig1NUiAoa7YS94BaxCDX19TEzCSvSD3ob/EBwyCKnNP
Olne1wUaJaxmCkKQOuZzHdCEFOtgo16CYlv9RekWXQflrgtPigSoPR9QOjnk0DxDKWcmqNsY054B
fICQdWjYytLhveTS+Gfoo2WmOHR28iN+xgc9LwxBTgCjhyOMxAoxe5cy+eIL/9kpvGZzu+Aqj4eQ
rK4LfR+eA5jcsQrH9comrX//9AV6yaV4jv5ce4A3XZOEDEYQ+WdpcZ/if/AOMFnzA3p5LkIhSRWv
72cSZFiqRASuDbsy9nGy1UT4rsUmU4P4xZRmX8PLS7ebOxq2vTqpiA7tHRBkRfJHCDtmcVLkY6n5
zLRqE5xFkaLaGBgiTSEPyeLi+M514HJFUGqi45AoXMyPDbRX61m6xv8g0IG0qTqFktOAIgG73fYV
+YPsCy10Qz3OAIjAl3mGZ4rmB5iWHxbrHI3dXc8/143YdI9YxYaLxyYf6ImW2SznR25reESwD/ul
9A60Gw5i5Ut7yaJy7Cy0IaNnRiRThtvtsqBcrFUgRxkIK/fHXua4mWfN9NxuZopmL8u86iOkh2Zl
wT2qYlci1ahgFAfAPGguL7uyHjOvRd8VfDa6SQ1I0d5wn6IlPGD5vF1lNVlmYXQ/rY9X/589b3YH
TyAsgofswQVNITEinxbcK05SiRm3O5e4XVYUfKtI4tvI8QvrqVrM4cRnmIYImZ70YZbLV5sJpXp3
ADpMJaP+xppNeISNGetBhwd8QbVXfh+Q2aB9RwHvMM4Eukq7Lqxh5HjETrIaBx5rN3yWoPdk9o1v
j7RHIk3oW9JQsBm0OVVCvn0GiprSBA6DqeFY9DhmJxPtOcYV6IcBxjDibtNCS81Sru3kUitvy1fM
LB0LfqGiwyqsFz7ILTr83tYD3APPrTW/X+Nb049lhzbpskKUF43TBJl4y36hcctpTwkCOwtKP93U
yDZfznOUZqMl6P/6BZv3BpsdBXKRUwC5A6x0QokUSlBVKAtrj4jLa7CNXcnyJAm7DW5rbxk1ZIWZ
8InxcGCb+/uHCE8FzShDwVy6ifzQepzYsvt8zw+IQkf6WZ3x0J6yQhOxUALQ6187ymtK+hKIA3mQ
VNHwzZ5BxMS99LA9zz7/Yt77dMQqlx2vr1fsNesKY87wIe1dI9hFcPV3MYfhZsVS4SU5DCoc1Fx1
CA7cNgwb8IDzNQq2AKFSpCMX8l6388vNVjAdiC/8eM/pNv/X543HgRgkMYKBJwMNpgp9FtqVS0+a
Tm4lhi7xYa5Z55EzN8g5qI9PfEswB4GxyEDpwUTOHkN1UK4F0R9zkrfke+YZpmvoAQG/ZStZlUna
T3yHrrUjxsAYhoECEKV+z1hLecS3cN0iT2vnAQ9MLV9LVNwQxN1pt/WhUmpUw3A2kKysIhPgBxDX
x555q1JKYCR39t8wqq+qQ0EIgGQ5d6XKpKEl/w8oVql7Wp83bKzoSW4OK92C9JGYiZleh81jnCd9
IenWKhrBaaMiNjHO9ngFkrgl41HqkoCoWnbmSI9iS1Qj7hAwx2GME+7Qb+L6eyvLXDPmeWoL6qZY
4IvTt2btGCk5AaboXbxntPbgWJbqkoErt1w5kK9ckPo0aGcy3Wnw5Ftf0iGjulEwfNsvEdzfMAxf
rRXqEls1q9CGEgzNlRa52yazDbwU101JR/1YCph6m9FLgfXt5IIYUZOEY3IoNEpAMdRdjtu7ck9Y
cB/CUcZCxKWg4B/x9ffNcrS9+Lu/UBQW1W6Nxi62zCODSuiBPY0jpWPpKwUthnPNEbtXRpiCO294
tgNztV9dXpgwMdwcQCm9HBnYTjRelDZsd6H7FkfyWUTph/I3cCjyAmVPqgGlERFXegj6TBtI7IhB
RdVqT4VyBlS032wottDS8X67NHed609tdykp56kg0oTpCKK8CapHOaoOdtRiGRMxj/ozOb6YEqTB
0zuWV8rbrI/+JNAlzEbfDqzO2YEfhSnA9Z6UkD5VvNQeTQYFydEkfHzK5OLILqm878ImtmPqLcX3
GsN5smsJNxFial8zXc3QmxLyGj8ykhF2AHB+mHRNtgwECPvmioUOD0eSHJ9Q/HiYVhVcmNCMTUgL
eA3nhaL0u0aF7wsN5EFWKv3JVV6dpa1jWRKMd+1RRIW14yBmV5DJAo22WUQfIRqwBqWHCDtBY1md
+4GSHaoY8Wr4EiNrLxK4pR6HgBEU+QofzeSNPagrEegSRJ4g/m+xUvap3EuNsF0qIX6mk1KDEbWN
4t7nT1qDMK59O3sxBXkW1O4gQF+uukXOeJRR3X5Cl/ZcXlZ4LERfbIti/aKyFYypnfDR6CN7Go/E
f9AM4GTCFdTq9kztEpz6Q3gobwADOJ+T9vj+If3ZcdhDtmVhKlm5J3fCT13bMwFQYIsj7JUVOKmJ
4D74gcOz3VEd+vLNAVNOdvb6dJACSoj921xEVw4hP2YSCBlSovuvb0OQ0iIWnIeXYR4wb24hRmbA
OsLx7rzRZkniIYa0HeTtvR1DeUN+HHADzPFq8XEx1H9zxvPBDeXcEJrJlm7GThSy8uFuA3C0Bxen
ctSjkSMYTRMGTBGZl5PUoWtUyod9fGb6OGofJb+gFiL94WIxJAofKO4CkJo1Vk0zl64JdRw3ZPQc
2ab3upCZu8twnIibSrJlH7cka8KUAPUAgOu6P3c8QFTM4hm987nsLBmUBYLQsyfpS76fLb1zjYfF
3wQn3xNjMHHWXl9tsJYgpu6Lnl4kz0UgtITvMGCd0FzZ9uCko/nZ+2dEYJwmR1Wu0tplTesRaS56
alhuQ79lzBHnXcrj/pjwM74CKnA5CDyrWjfW3wwMVCCL8fqZqNb5XZHmS7pPjXEinpgogoffZOEQ
N8piI63/TRyGEsRdL/y97fjL6mf9bPVblfg4CS/+o2wyL1l73RHkSgjmX6l9EVnKJjR5E5fzVaB7
Sjsla+53HJzc8le2Avrc0N98Tx+FNoFO2tXJFvJ5ROIBPeiL4LdBc8+jO+I+P6aHbztY/pByeIFV
0tOQ+Lw+T/53mfaCcMQYQp3Zq+mug5stFgoxYXjtqMWQrzBEZHXL9UzhS4nuNArJ19wbHPQy6FLY
OIcIVITJk4q7QeYbaEIs9qLoknteo5y1ROqXTR/XtJI2pApr19S/9m8gHNly/RXlCW8isWCjenDI
VCpNbc3tUXB4j0EoWQRUTR2xooYdBZuOyuZIaRD61Wrlj37VsOWZZcXd6V4gm4tzmD6vdBHBNpPh
0N4RvpVXn74jacFtHJTqPX2bjt4MEOVR6mfJWDbSGcnYYCUy7hVQuaEhgDdhtRXZEQrWQbFC9667
8/7I0AL0EKKAjehFXjZfa82c9FIn3NVSrzXVsYI9cFnOgweX1KdHct1XMIMA6FRLGmfvdmY5Ipkc
SqZUZUUYGTon8YXkiNvL4jR/wisCS5eYuaLAFEfm7eRBh57npYBT9pBqaGzDJi8wIBfVwiR0C8jM
QTqCNoJ3fk77UKLOJxFi+FZTeK6HgnxcaAylAc3QVbX3ezJCeW8E36+TjpHvDghwgpZUXK2yfR9R
UP9QxZMpFoXh09eI4Lb6K7Jc8cGLNxkhD74lHaKzVGxBydKN5oVn43fN2JoOV1qEbY8UR4fH0mO3
crokXfdqMx9eoag4lzTU1rDHaeU+06A22XsPHkUynQfEzCLR2QAj6P8m76UvzUx7gvnoxkRuJTzO
0iAhdohsuLTorlojvqgDSLCABFe6BwIgH5xuVD0+qBmvNuxN5CZ6Kts1u0Isy1aMHbF9f0A/f6R9
je4+7VrSmhvM93aPZXeGx1kYSP+9yCAXL06hYzXL3avMEsfdljt+tfiCFd8ZXEJRX4UTv7nRJzqr
YOwNyDqCG7z3eOoLMUqE78TDiPQWdi2bePKEzQ1W2errv4dfIYgklhbKa8tLAHvP9ZTEPsdOIp0c
2DHkgsxSAwbGMJN1Tp8hi73h6qpaQyUxdaBRN1STniTBtLT2+FK3Mk8GIGkwEyyVYwM6UQnY/Rca
maVXs7Ic04jRbJvWKSBAWEuDPkUYZTQKaVCsleB885+Zy7NERD/TZ9p9bvEjhc0Z3g+zloNF4Xrq
DtYGHiOAIf6wvknu8G7rPD0Dkkeqbt4N0sKa8VNw7NcWJUgzmRpbai3dzyViW9llJzrLDwWvege8
EW181WBnTDUdp2MvSOgZkkMFu8AFKmuonrhnecUTTO/Lrs8vfq6c9MQLt82YQ9nrbzPbI2jImRR6
EWHbYqIflgCxgKswmrO+BWZkmbzt05BqduyIh2kh/rA8NkEY/gFpSJPTRUUyz+tl7vJ+ZNWhjAL6
6uJqp9kEm4+wkSpQ4rcxTMjBVqC501bXRX//PCiF5s0ZSl/LUqEbxoYTZVRDmH6UrK+hb1cuu9O2
Afe/u+xwdrxRBC7LZm1FpTdaaVjKCN0/3fE+/gRKk/qphiuxw70w/+E/U9X0xaVEmzWkUMJK9vnE
fLYce1sONuaY/CEqZwiSaBcqMD6g1NEg7Ec3G7UqWbyppBqHKSxn50a/jurhoPloIeDcF3zvRnED
tHP0RAHAb3JlTUsLsBjysgRu+PuXdKzRvsoerstTvCfKc0a5RwsMVRsu6WZxp30lp41LKaTRI9Jq
NRBTOw4qH40fE5ND+IxY96TMzHjNT02aCKgtv4/7E/bB5LvH0tS9FaUJBZQrJAJ2nslkoHKTf422
lVR66EOeb12L6Bq9HPsz95adnDQDfmnneFsxM7D5OVJDXSephbHDLLZt3imFbEhtJsvJjEg6eP54
z5xzlDWzV9FEFDWtTBelTP2sny0qneYMm0QWqF0qgdKQnQVRRIFU7PqP7GfbP4aXLXOi9nIWUQCN
GRlEUa0bpE/NmkV6sK2QnuGAU00mt5l/KAnq12aGRvbpQ/8mU4MjkZzcQQ5TAroJyFu8+t5RaIE8
i9XibOcUe/3rEZw0/k3xNr0Vxfai+z0fESnDdSrGa5jjQSOmSOGmt6IAbolN6AmyNOyWd+zlJDmJ
2Z3yQxwJvHNm8B+voot/hC9p/tv2zjSXapPoP7BGiGQgPNZsB9egofnSBZYKCCbHdRYoW5N9wyNQ
9JwgqvIN5l4DDjbdVinn8NUPT/QC1eXjHVsBvZ9bdXJSiwVq0acIoSGRbn6z+pD832HBPvjYc30l
AOhVcBgqb4TrSlbZnVSrAHHMM9KK8/aDYZzG1CIlAywkwaUeujIcU3J9jOIVzLbQXwU57P7x8lwm
0bdnbz01sNxocIgDlR0osC02FBe+a1q/tnYiD4I+2ilvBP8o4t+0XQiwDSrAelFdA0xcqXiHCEmG
oC8piYD81GE4iHS+OGQsV8YqUeQSm1psYDaJxuCji2Qpd/0jhE1XTqNezKsM7jb/ubza7khDsbsR
IbPDrj8s1TvwytmybkWEUjjwyJIx5bhgyN97rzdr4wOyIKWQHQoCaNlRA2U0U9OnjQISkKiN0OCt
wRbYBVw2f4GuaF1G57bfVM5xqz2AZiJ8ihuI0XOe1gzLkRNJoeP9mFaG+AwTdCY479pPc3JHRlQS
3gU+/t7ioU3nmexK0LBz2eTnvyr5w8c3LoDyP65+DWvxRvSSoznDbCzK1Nwv6QhqxsTzi47IuBuS
Zo5XmH8NUBARq6tt8nrY0P8uR75pNiYuu6x9tctZOiO9n4YND6yEMUpJMX7cExp4k97npxUAX2Ts
82wazQUXIqo+oOsH3Hbx3eMQf4C1otkokKHM41CqkigDyYuo7U2jotu3+3RJiDPKe/sDZGJ5wzpJ
xIP9PM71yS6YJ/Zv5c14G4xEPkg43WewfijwDWZ6S4ll/t4pUWL3LNCkDVPvx3CP8AX0Je2C7r7K
q+8MM4ikbEjKDqG8gY9LquOgiLepvsCxRbTYQRhFvt3M9zu0SgbUBtTdBNwoicCD5AtRfMq7yPdZ
kn4O90wI8o2HUbDcCdbJ324DpvA4jPYIjR54K4xhDUN+E+qZpSnbmY5y2Obc8wCdVHUKuMDUegUP
wLJ2YJt0avtRa5EceUqW/iM+RCynLSvjNmgXXvyfTQZ5SxQYipfkq+JOPUN23ETXldolUKeCgiyq
Qnx/jKR8rmmktOjLUODQKbhFWpxZoBt20ixPzRQaB0W7zirjpzffxvT67pUenhMsCk6naOvRky5P
j+11I9H5kH+YrB7ktzt+n3ZczWWB7zwQIlajZWmTi12PIhGdLSuL9LrSmmOQy4zIgpSY5fFTMurH
h1EsltXHtNTTtb0IioGqttQYU3BZc2Y1hY9Y/sIEKTbbexGz+x9dO1ko1ePyYfppzBNJn8nxVWwZ
5dPTeK3nm2Y1lXdroYioosOAH1RXaro0iw7lnfbsHF14nylSsIyfza4TrTsO6E+MMIPWqg+nuNdq
MVLSxNZ+qqzrHnaI3oBNeWM9wze30l9LwnXhyd0DcbnTnEEpYHGgB5j0drO/g+2qXO9lGGzU9WxZ
Pql2hKlxerZJu0x13noVIJ96okAr+wXVkuTRBy1yR5XoeG16O2NvIP87toqg85okmOsdzNR6DqLc
tyc7UCOnw6qryi/injejmqdNSDvo6Ay9hIxuYe3KAUYVyz73x7KPHowINmI3u3SGOKPOepwFSLia
yPt/5iAGLz+eeybZG5jAMn0eeqE4cBMSASLYGdGiTEKQqzXlGSDElSSanbJRBOGZf/7CcOJrl/XP
mll8J+iggTKviuGRaAe9kijCaXXLEacB9WLCqI2RpAQrIjIYE4Lsi5nlBWtoN7zcLYayh4DSnJKI
z8oCwUaYc4oWovwbnpHZb2x7+F+qfes3uHpycSG8vAEP6ixGXvqabqItCpOw5EQPwYi1io1EPMIz
QbOm1uERFW9lZlEMTMEmSSs44z7GlPm9kb457LMC847P9/mo/4/TA6xmOwS+2Hq2HzaR7IQf0TVu
JbT3P1jKJWUy18QURfF50ZUNzwspGvECiBw9s6VJItMvPuJze7ql2JlCke4Zy3xMG4SdPQD6m91x
JrShB2QMNNK4nCbn3fDWjRrZcdqUAPTj3Z4q7kCPoNEYCg4HnWpX92eUVHujOAyHfPM7MpXlMdLE
t9dPBxPcseVw1t9sbUAe3GP98MsAry4/u2GYmtf6MkBb9/EVotaCb80NRvdk1DT6AiPxD+wBHv4B
gB+4/qVd1rNI+8gY0kEwpe6b9eqHp9NW3THIjTVK6ZL/WAODXyVjuTQbH7PHDetyCyPL5vLQL7uR
XUFVzc1r+1CRPGE9CiEgTVhwD+JeG/Cfjxn7Y29BwBY9Bsz0YSwdPANY5pHtAX0PBXDJ+4RDRj2m
a3wSE+dMW/9GhWDYm3TGiy26JVZeWJ8TheL9gMRPY+0/spRqDFSQDijwRHXoOqG0+uf9Bd3raLG5
cHcFydfxjRY0NJ4KRmHFtggcOyeoZAWoYNJMTqqz9aatDQT6RH4muO3PCpvJHXDY3RHj7QhiZ/HK
CmKsDTxerc164tqRm1JTMOTTdrx6c3PKxb8MkRb6HUg5podV4jA6E1TrIZ37p98aVArPaQ7mWYe6
u7K5SvEu34qyetDvvOJqy6fG9O2pp8jmXoSIDHa446yxuiMGkao8gOwPx4+0P9XsdGmG4XQsVJOe
SVfE9hD7Z6fJBn6ly8jOdS58SDm8z5mEAp9QkM0pslhLMvVwhfWjIO/qdSIqalCorhtHgDZ5eQ6o
MzH6aBekbk8KnolAzd7XPOrYKgeBp66vXxhLEHYsVQS8gDFlfLKvvxKcEAjkZtnNKkXL37nguGSe
p3xwN8WIZxVx+2fvp/ItJ6t8wU2Fib2ORsJOR4KHfc1GG82pZPitfR7jYjLHfGnnqrEzdWT0jZ/h
bgY6O1lZE/ccv2ZCgqPrH4AyXbkXg5rVBRjhPg42QkCFxlzBTiWtt6Gv/FSYh28G0IWD+49e1trF
QqDZZfMixnvj4umOQ4GDQSTNzyHHpncGhyeYcgCdQUPgYK447vR7u/ZbO+LmsboFRdEjM/n32YUa
w49n9n+ODGKfGMst7nEtsF0oI6orYCJZwajmZ0NGLx0998bDEiJ+ba8ueOE+nRk6+gOYsHoV60Bb
3/bnUmRNC2uxkW04g46jW8QW7NR61YmWfaSP0c/QaNy1X8wKqag+BdJ5EhTdFZbH57rayxgO1CXn
5SokGplKFsVGhw+wfJa7ZHHUdShzI2E9Hyjd0NayxvH5YnQWGLMWJpjnUCW+tJ4LAXF4KGd1PtXo
XCMsaXTb4zTiZEjR+qLasqOEZHfdCEdu9odIsjn2hD1Mk+kbk4cASykPNDNRdz8LkVOz3CAPCy9V
u/iBLUaTsG2bIeTABo7cASpM5DDqi7SBDOTgLmAjFG/1+iXw+FNV0YRpvEZjfEEl9lYSxCLCbA/1
HnP5H6lCtdUtqNN6kKaJwfh2pBh41IadEj0HkrDWixyfXyD316ckHrexEtHI2hv0/aaDpDSBFs7N
j7MFSzZ0wGLrWNpuNA8dHd2VZYDQewqLLZEz2ikcak81gmAHSPqN9AZf1O6AY2DSO98IZ0KCnssu
YUipI6GgU5QZIN/Ku6j3Ag1FqLmXWnbotilMVO2m9R8gXaZvo9W9BjJ2jHDxxPZ03UvBGl4gKsfZ
pWQDNwzqD7PdiTpkT90iEzoHaOrluSqbnue/Yaa1gUD4DHkjOM+jbLjLGUTypZ/9tZpe9L32dg4H
T/q8dE1oN/OtwK7N8T4NbbhbWU+Ju7hkZO9sA/d4v11RFUDG7gBZ6AGDUvQb1RGmdi2xXAT+1v8t
NOja59/Nbb+PKSfoHjT/uzD46LsuHvAucH0E7zPaXrCIWWGQe1w0goEE4vOsmriw+n9hVw2XmCzE
Q5MRiuXi+SJczAc4JhbqW0spzpTN+fJKKA2W+CeucghL15KS9oNGOy+m/u9tCN2LRmEb6wWasAWf
Ga3hERI7mwRGeXbHN84hOyEvpwN7J6025v5LhqmfdBHSejP7FkGdfrFaaWhkknz9oZhB/lHxWuft
HwzZ7u7YY33RXcpqopetW8rEdHFh9al9eJcgldJFbDV69BqH/81tf20AiAteUEkuFwZLSSzqcZBc
Eb0UbOHqU+j9zhtE7PgOCGAiDcvlfLOduZUwG9UvgHbR8HF7E3vEY+WFuMTSlDqf1ZVFLmbBfaev
+zs9QCIUfpd6K98Xxznhhv/NBGqFhhZsR+Ps3opS/Yr/YeQs75/CL/kFOt87CjKHC1q4+XyJun0U
HvYbln87x16n23y1uRKidNfOY1/DE/+YXEjKV6Fx21iGnILxo2Qenac4E8lOjjnfqCB1kjrqGm8e
o6lIKM4O8NyqlYcJDSCvOSZlvVE0BRq/MqJGZn3Ujb2RZdy9kRuSknVKfgQR3jxUZNVGAiG+v826
pwuYvwJjw5Ya0/8+T5phESx196aXoE3D43E5S7949yJBC6S9wsyJ1NjP59sFyvCxNEiePVXGGsvs
FYGlSDNamakBACcyFV9o671cAk1uOlSlC9BU5ZeGSTP/V5FZvun9aoxNheuHf0NGeGJqDvXb7Oi6
O2PFEcDOHhOqHw5i3Mc0ZzTFJUFRzQM7fu/EVv5hSVglEnFuTYb6fnWBYaJWDAkUxPvFMCXrBeOs
PlmmUY7z5IQup1XWV2d8Og6lBk6/1mcbTaFj/M6Poe89mtVUuLiO28C9McJ269waNrx+PP8ubA5y
vWcZU1x0aI8C4QVWForh2nQpi35b2QwKSrXLPYPORp/HEsdR7Nsg1ZEIJmdXB4XZz51VMx89b5mo
OlVedftcmxJv4RldBwgAWxY+LpEpUoRo64JXgrt63ebrDX3czlVJFJHOVCbQNp5vzKmEmVYdRB/U
mYxaCQ4ZRqsmcNortwwToBrbv/aP/MYduBHkuYHIxbo2ddc82doRu0YmWKDGsmwjCSxubfY/svBR
QmZwJxiJRIdNnAJ9M8FPme4BJnfqG3+2D6BCjezBNrVjYQtnMfXHyCWJYeICHnRAYjC4YYnsBR8v
x5pR/YVXawfWp6JTvgZS7VDGjxqz18ORMbXVuujQ2+HPUjwwlVjCeGBeBNNv58Qt04BHsKwANAaG
Fns/JQbPiixVe/3pIzkDfbXWhdXWQw+fgvsyI0qlSLBicJFkGlH0dUgbSPqMgTxvHm3WY/ojg2Fb
egSlaerneMvl1M3uMmjiYMSpPatXpRvWLUHpT/1u5WoXBeW/oj+DysmLIIJwJzUuPDtccJYwHCBO
ZSiQ0CmvbdsSQFNzhaBAMJc9gHq0EMv77CUv8u1PEPgUS0YIDE+xmm8smUj3ha5ScLb25Or96ehS
Bg7X24bFGRKcVl1t15ZMsfgqqyMvshHbBtbxTWY9zyISAwnfxoh6QLACWkgT81DveLaKgXsjGDSk
3Ex5UaaoqKM7TxXHdyzFSDc2Oh3pT9ga0WJKgjA56qGtFz20MwOX+NZGigKgBc0smUhNi5wdx5RY
lcj6Tbe86EWN+humrT2TbxF9LBSX3uMdFf76snpCmnjeSTIjMbNsbXlLYV+3P4hnGtwdA8QrgYyI
rlkh1B1xwX0wEcArjavRLJc9lk7EiUrpf/pzbD+y4p6XtQL8zMwVdEKxUYCM2Tkc3pvEyo9tLYuW
jhZV+sljZ6qfE68gveL0/fmcDPZBY80y94wFNiOtajStscmohBVouBHtCAPMJxp4tsDSTTQD4I1T
lfMfLyGnwYti2ORPzt5GVd+SCznLeJxLSDyb5m/VTK/cpUqY3EWXpUB/7t201KPnKX32uB9yChXE
GzizPYjRmACcfjrEzjpJEQi8PuXlQBvizf2KsHIOAAh96M5YRVbfMoMk1pG3xzs3CwuZ/kWGAmof
UBE0tllqEykeZ5+PdSxJExvLADml6D3XASCaLhYIlrN0A85fE+5oZ6CXfsxD14Y0RGC+LYBusfcd
EUAn13XhXmiDag9J7mVZg3Vz2ct3fZomCXyrr+qaGkSyjN42beRkYn51xIP2Hm9iWgKy/NpFiA/V
pi4YGBF/tsNQ1oWtn+oq6c+pJ4Sj9pcEQacPgxty6qXP8dilchzvbcioizE1UVJzJtzW2rnRMNS6
ph3IIRrpteSTJu/tXdupriVRBhqQhjJZ7he7K6+UHfyunPGmfwmQ7/EDADOhd9skfiK6EzvtrQaX
tgyX6aIZy5uxoODmlnX7ZnxTXl2zLQfQWgRdfH+/3EGGXDe7y5/WRWrRBd1np+gT2Ke/WWT3Eire
vJG8YyfGfcW18g4314hQ8rMQ0PBK8Oz3r0GFV9InkGQYQ3A95gt4/XvAh9m3q9vsiMgD72Lgx32p
CCb3VzpnYQOAzTVqiPehAAPX/+e2Z3nuXqqMk7WIAOyNwr/rDDlBN0CX7KLb2K8JQt+n6j3bJMG6
6rsbJRN8BDWMLnpHTgWX6GY0HgAvmggWsMw2fSLLYdEH8ClBrd5zo3PFs4lUvEOf/TmnWhh4TDwi
vobRNFvEq53UAfuNMubN9nFxKD72E/+oQLc584+e2n0/v3YapypBFBFXLNa2WVmDhM0jr3CpyoOP
V1TQLJrse/NCaM+LQuwhIhdDgLCdkr+NaI98oyLQi20u5OJ54R7c8PWfNN7DS8Tqv0o+Q9Heq93T
Kn2jSEYLEUUs/W8AbaD7XRsZuZhiQFMGvNkNpcRcDoVzKl03pV7tm0M2RcNwMODXY6JsFbJJG7H0
VkeBVyl2Y0q4ZVBVLa8bBh9348ZMDA5kmWqVI6xj/rywwmikz8a4N8xpVfr/nUvC5+JWIh/U3A9M
NqA14Pav8HQiGGGaqJcjUJHWvtKfOyYV6x9DM/3ALJ26SMMenssG69df3jfsfHGAMyASWhqD0GaX
DSbhqVe86kJZDQ44VntegukFc789mqZuoAnt/uHQ0Zkh5JaErFQ01IaN2pljAYppfzs6NSkhJvhl
+Z0699TxAMHPhWBW7P0iQN6xg+frOr88ey3F7l07T5wVXmjX+eep7xU3m1hX2+tnsHJNhtpeCEbo
rKafx/2gPPz9+wPctVI1TJnNyNuWCS0ZM+Nl7/9EzYpfb78vKiP8UbTt3gwlqxv/kejZf0KraXJs
gkpYxPb9+zhyWIGubo7UuDttgnGh2nW6hl7er7139BOEO3NOtUCROPOFoyy4OrywF2ZwvsiiR48r
a+1qb/rrB+uNHRHJbcgRrxxAgF9TUs/ZKftJ6mCrbMnWluwIkHMntBvWAQFYXbZRLS4lnBVqMExK
A7PwefSWf0Gv7wyO1QotT/uFVylGM6k0Xkiyb9pBE3GD7YnpfULh+naMu39WvtBmPw/o5f9L0+uw
GhiEswfa9NABz90dk8iFl6DWkJRNeazWpiLBeU54SAZagUC3p2N9eAIOJdkN2M1PVeHqnK6JCFnO
tuu4e7lOdJ/h8/jbh3S2N3BAEBrOjBH8KV4J3xbu3QZ/QFdOHpztwTPvMDXj8UN6+T6b4LolO7cN
hveQm0GD43ATPmjBxRXr9QGhEZrL1saXbgyV1SYAWahom27dcWchC2qoIsxSO86FhD3Ah8GxsUw6
I5NYAAZHPIz9bOdImMD6pCNp+XhkbzrdVK62Za6d7RvTHFVP8RqHJmbkbOL2Z+0CLkDDSZOZoHLJ
/DXXUfOyLUTz4HBIr7quHk4u4K89Y7dpSIQyEnWYMf3f/4cyrBsGbLTAi7fAdp5n/XT1AcOHF+YN
qj/dxav2AORFgqnunePoxkC6qtjmwp2u9HNmy1ov+Je9Jp9zS7D/feuFs2jGq5+HITlu9zYeGoFH
AxHwwNVgXV+JMggQQThPclePGSgcFkPN7Y4I/pPmO62q4M5DIdN4VWbETUirOCyq5+S1LoxutvhX
iv3h25LlCXgWkQFr1Qo5ZhHKPC4ii//Y8c7m9gD74XyajoiYjrvQPDiokZLW+roP2HNTu7RAarv8
H90KTp0pLp3dXuWKr6YdqBtqpZmT7ZydEiWFjQMj8GgqH01vjLDPskTUB4/C2j5xI89HfVuVVSOF
tIGx+YDqIDQYXkZW3gcvOwIcaOCMd5HOB5t74R1ClSRfzDs+E3Rg0tqB5S1y87xtBCyrjj1h8bLf
ir850NDyxYWhBvhY0AIxrsnv6fp0IV88VoKIaZM+KyADApKdmUGo/RF1dTjK7mcn0t+XZskNl8T7
2cwx9Dm8z8+wtKHmvAfBzsuUrJqK5s6vehurKGjpZVqiEZwWQP8lxd4aMAwb3yXsq5Meuy+SUXUq
WYlvLnHAtbWiCCQnMLWp4s9WI2LAJVL9Uy7XdI6hzm1ZgTExTvviPyj2LqRF0UXICJLeJ4qgkmY6
8p50bZ4yhOgdGBwLi2FxqdpTXWfzhS/3yV2PCzLuDYomOh9j+AsLUfsO+TKoRu0gIM/hETygEkhB
5EW7Agxjy24PQeYRcBkMR7F9o3gb2JPQ1reSyFgdx+U0FpkAyekOLPBiw9cFtEPj08fOWEIj7pME
XnDsGTZzwHQAj0LonYSk+GPBSWDzn7VkdApwFoTYdJWfALuCnY21pJDDgHAXrOpdNMSLMOZZ+mWc
EWBE5f86R+wUW8XEOgmhynZ95ZMZElGTI2wJIReZi6z/NcBMOrqjLpBS7x6gGluLJlrJ1BYhH9Xf
62qYymCJYXSbyxZveKE26Kpf7DIt8OZMp3b0hP5w02ZlOh4HtjEhVZx+wSGUywVczZl35oQgVec7
qSX2iLEsmkMAg++CGWUW7XHSFizCC/QgRdqKzMZCCeQdNCbLukcWuisHDVhwSuSFXEnOBR34Q1/L
xI+NMx4vsI3eLO8TmD2sB07bOzgmVfGhOvfaXn6LpHaKQQxqgOS48qSNLA3p6De9xkKPH+i7JyW9
95JEWSxYBX8Owku6bM9HmWlgIEY32SzDfWyGozZtpaTgZWH2Gddv9wB/pvl+qlddtOCSxU4ogOwY
JiXGVoCRP718JEaXJEri6CoD8ORUUsTJcsP2/FnHslnP8RrA386NBn2vioCMKICHjRkEawqToDo+
Ot7tycIcJA0wqxaIEPFkxqVHrHSPnUWM46Xpr79ZlTnCo+iZqEdBwN7tp9T8HdigmbaiX+OTftqo
3IDo1xa0istrawZCneGILaBSGwCOdBZ1VjYorjLsz/agKMQzQ6B1x39+P1W7agmbS4jB6Z/oeVsr
/O5atsw+4Ssnfh+GkhrrWUxK/1+Zf7Sm+tjREd4nwNqhQE8wLHcjA6+2hfnNc3Acvib+FPDvnYnL
Nwq4L2jGz2Fqu5tRimGqnmZiQujAdqX3JjzWTRbM1Cw/384DhM0W4BQkow48M1HZ4SxFKDSDV/FO
I4nGNzH7aiv1dVX9a2yCbX638WwfBKXoR71XGeFz4x4UkzMbgUVQWMXRDIo4DXYHW5fkS5I8/Uh9
OeCSofptvAF9XE1b1TSFqxj7nciRBTvuYHwC44dg0BN0Gw3bWOEb6XUZBcpSJjp0f0VWDQjktGXo
P5LAFM8lGio4kGMfVdSUbgqMrmtSffgjR2QXo6owO5rCZEVfwk/lOr7ShZ3x9ZzN2yo20gHOQcdh
r0n5LaESjICeqoj+5cXIBHbppVFwyuIVcxPb7E1BpTDNASBtWtjc1/lVwz8hvsP13M+/E13iaFTV
Z7JbbXJcSFym6WZ/Odi/2VJmkZzSLFqzCN75taQ4PHebhHCp+4IdxtI2UpbzoCMnAX6v0iavimSw
9tc190daHKzIAWpgCnL9QKmKnQ5osHLW0tfBAIaEAQgNZsGvclVy+iXJACmICrq6LI+/BOqTM3TS
Z0MU0Dcs5ksbcE683eUzngCjgn1w4OOVio7Ts8x9xuDh3KcIk+bfMVAuLb/U6Wfftiti7mQ9yFDb
hs9Tar/0kgqyGzLFCotbecD5Ku1uvlGxVRuVTOjjYXe0WP9qLaCEd6VaKFSudy1cXMJz8S3vcDlc
tO52HWY8DDnatHG/S+q7vTpANeD7bt96d8tmROY0GZUJKahSWJs4wgVDMIVD7ndHuAbPlWsuaYdF
+0jJt6xTq6Tfi+TP3NhJdjpmwCn/89SEV812XN8coNQ37VsK18LWwRuZ13yrfMwNJxbb8783AhVX
35hOiQPQp4wFIoleMJMPduT8VoyQiopmTBls5d2djYmqzqjeyKYGAz7DjkKVm9oRzpFdnme2PxNT
7+ALaRm2BuBfxCeZTky8U6hf+UK4Ti9EWovGTqYb0QVnSkiNyctfBk7i47pP6a9ne1LZ+/pQSBZO
p49ZHANowwJBxSFpgjMFW6sVa7KuWHQYM3ccABFQS1b2ytdR4ioctqVmEteXDvagmposldfR3Noz
IJKuNi7HukLZUzA29rwhhyPR5eNp5SWKM2uY352oQilzGzT3SXgC+bx5kygkuMCO6v8/B8TbDmwT
Of9O9Wha+zsh8ybCYcI0r1a+02sFmBcca/kdXLWL9zcHO1uAhRAP2fJLjRuhAKNPMOItmw0XpIk/
dNE7RGGsrpgPfjky/5WJwXzD3FZyDLkqWsqvgggDXHnfsdc5GBKLLkK++l/4uwAyxbNabK6Is4hz
hKaecMUqhwi9QDGuRyAYTJGvWIbimsEFE1YHbx/1jEosEW/UisTmaT5RmrjFJIDbbmtje1szVk2l
Pv9E6nBak9OAvIGvRcwy8RmlLfV4i1Rbf58YCU0GwQqHTEfhI0Xe226PVsx2Q+641eL3YbGOUud6
sEQs2IqNbf08WdRM14012525TSma0oB0cMtp2EmrE3zPGQVvm+vHizYj+kXMxx2wgqfkj+7vkcl6
jW1tAhZYHJ3X1S5XWrZhoh7n13kizjdrKQYPtBqm4pj3e4EW0zmY8Sgg/XLXeGU0rw+S8Cn0pHLr
iQUbu0M+Sdov0+Opc2ZtFBJrpcCQZrXto3k5r6pNlWSv+ZwpXK3fmO1x7zEF03lmH8wwZ4lXnR3y
qwVc7Xy9gWS51N2Y8gR6lU7yQkawBkITDRg+1IidMGrEKuOl7WGt9yysYyFVqWFwq/uRuxpLZngl
IrGnNMk+uDYY1N0R9STYW26QIfGItz1xks729dt9LSBivajYL77rneQysjh2AbHaFpEKRJLZH6eQ
jdLse7rQNpcUTnQuOkxd/djifR7lBHkmf5Vbzgsdvh7HJb9mVSQla58mPUAi/1juxjZs+oezP7Tg
xpKg8QiIgko4DSgOuidE6Hsq9/dQultNokUGxAbxgVvJw7VNFK44NGzFJVs9FUCc+rNh4PwaK2+g
AQtxvXPZHJ/OErzUXGqEeAgvigs51Ta0WnOiLz2N19TiB5mBOaPD2Brq6L64lnJJ5zWbpc3tuNRu
tGl3Rqt9szjzz3ykU4VqjaBBCJOLZALLAyDdoeD9J+S/hs/k0BQTJcSYJUYLn1KXaRDsrUT5lkOj
LBTM/tNNHppdaYn5+X44HyJtNdS8deFvYK55SqEWAjfEFQt82ILEHsnPNkAAiF58c7kiO84BvnRA
PB6IL9uE0g7g8xvkjzeo1KkNqMbKSonPMOofMhTZJRVKXNA1nF+SAGCICmqJ46nTXON59VvdDPdh
6aVwCkcd1g7dI17O6y1R+nAZ5zr+ds+7jCuQZsfymJPtFoq9+txg8Hti/2s2lE/6PJgYVKfqr114
4smmd6aiG1vFnY5am44ub1zcModxIT14JeVyYU5t1Y/LI5LD4My+gF7PiLOdEDabEJeISrqHws+W
CYZD9fZZt9Nm6koHVbOtW/Ew9pcxVbHR4KJ9D8rGNJoKpz5i82+tKRrNlAQRV7YF7eDPNlbDRczO
7/fsun4gVM0NEKbtJnwq/x4f/WXM9xc1JAI/YVifpE7gjaWMxFozi52K2jwIzKVODXX5PIdB2MDJ
MkA7u6CB7dms24hrYuXzMzBT0LJYn187PnlpEcyW5lDSIrJ1klVVRgIFLi+9VIVD+OfqSJIpHj6d
kU2CG6IcOarG3QKKlYFL3QDpLsjfEiL9qRqy6MQEyUI222xd7BNCVHEvITpKIpxoC6R82bYsO4Wy
rmi70phh8TAFxDxF1xcsx44E1f12ZolntOUuPE5emX+tVfCptq/yKNrPGFQpUsMpV1tIWLIk34yl
/BAE6CcJ04PryqKpbapO6m5xwBDWfZapMrGcvrA5iYVW819x2E8OssdsoSHQWKpo9WRrzLV9NbII
agpC2qwhLgCBb7Af4yB3CwqhRcqiRvujuy8qojA7k2vrOml+fMCZYiWCCxrHFBXuQsruLorepH3H
lTOC9uvV3qIVDwgTuyjTy0goWuuuWjsIQFyqhzhYQkAQrxRI+6zUtGhIq0IDvNNiHRjX9SvpJWqM
skJu3r1C5oS3F35A85hW59K8yuIGga1Yz2wnpp3ycjLnXXda/0QMBMNhiDjhSRnQVsBQWJGhxLs4
F0OOcibbVNJZvD3Of+YK4lwhbzd5eJkaPd4bAqMNZSprCpGCdVNsjz+wp7BegaZ1Ys/+u5pITZLE
h+D7IWnXYyBy7mJVz7Tw/f8QYn9hdIGTWBm/BjaH532+0SaBYSO2aOp945oN/IwO0SxstnKIgjgT
P2wd1T4FGmq3PGwMZhryfz1SP2qaGjXz7IoVCXqzF28CvX/hejlC+NRgOa4vHVwUs/O+uj7gYp6r
0RtFRYGFQ2BdIDxuowPchmQfgwHJfwmOyiiJVFbQxE+N4bgalrP6ggr7xfaV9u941UqMzE4yKFJD
JgvH7Z7LSnQvsTfJeVCPVL3RWUPEcIyZpXYjYlJ0pLlFW2I28luTFsdh0fZaTs2hS//oiMSKYkZ0
ZHFLv3mLW0zPjCIDQgX/4E49JCIM5Of8xyqpAtFcK7A0pvrXMdXjUI7fudhri/Lp5Vs1xybguIcH
AQL6cLqHcU7GX/Rwd6L/V0AEwrMeZbJsxj8WJ5/JCK+BMXw74oy3iqeqdYBApzT5FCTVWL5AtuAY
/iuERRj9bZa4Nni3hfNOAIb9CLlXGLuvF1EZqvKuYAn+5B9fxUMcQHf6g+n8iDWC7s5ybKiXpOe4
FdwuSyaBiPf5k9u2RVdKzLzYZLcEMxqOxExr3AANNI+0ecZezBPzRKnqwWx0hdI9Q6t9BB9+UgaX
Ejzju8jPCCDor4TEMs48qiZ1CaZXLp1EGQMApeAqMER87IWPZJlmDUgiT4XV3fUiYhE7AnZqxiFr
3PTGYOHFUnSvdHXX5uvUts/9oJA9ZSDLCP73bt5xvnw+IpERltVhC+Us39Aq3mac2NDD4H/FxkHj
nR5UdPQIJML27JcZc86kMVV0SoSdJLTyszMZOT8RTyzhmr+DlE6FCy8gT4TdmEqdIhm6bW6YNpLI
GeWCpaXW/iGLP7eRY8ZHKADpB0xk9ekzbya/bDV1C/DQhw9FU1fM3r2Jpb1YnCD65Ej+ixkmRZtu
zDmqR0NYYeAukXXp0G2ydHuBLueVIwq6wNBX3dMeAH8XgPJwH1G0rJ/xQ7e5kaloSb0V7T0rfmlL
m6cnVOD0aTATsGf5kjcshxZdPURFQigi6p4QczaLAJGbhf6zSUDuenNAmgb1MVxjukloZMz50ipo
EkK4I/zFXZi4SXBd+HEi1HJX3B7ebfbX0mVS+peaPBjNzk+itGSrCoZ72YJ1nldJKkO+JZ9//7BJ
9P8NvSslYhof+YhCdPX8A8M1m+L6ciq+Ib987N7ezY5xx1AW22BipStWI4rl3w98QLlmiJ2GNVNx
1Rm+Gt3muQam5xxCaYSShNFG5/XHSINWkjYA0QYZLXsmIzi6ZCBGs558iFbeKNVIdB2Ywkjhw+hF
vgtLufhntd0ivshb0KfeO/va+5eZRUcoghhZeVryP0cQ7pxQtJcogZOYETNdKBrWKFYDy7LHVLFm
dcGAQH4vJ4PQgYfCkDX+S/RTfGL6TtVu0URbBF+juTjCNhAvhr7yXcp60EoIcIWHIYfAN2YiuJq4
54q+2t/thKTqzBQPZQUNUe11m+exS9cW+chcETbwqgB7ZyPijeE56/VqVd8oKhFRR4fb8v3JGkFG
SGpqKctk0Yiw6PUXjbH1lPGVDBrkJUh61bUeApFbS5wa/KYPENR2eexDbE9tShRtsxTeOYeezqoh
scXuOcmGdTOWJod5PhlQOHrFUQn8zQM4gx1pkCQ9qB3NWmWNySQkO22s5LvWMfsRzYJDA8YP8bhF
yKycQUKqWcgvSzySHuY2RcBLGLBR/LBvdVSyuhn5upKyw4m5AI0P+/iQFNAP6L8ZQSySJK25OrHn
y6pQPjheYO2ddzDtfHWr/apDdQJSvlKMpkF8VJgIF78g5gVY59B4BIfFc5nzRhW9b1Kh/QbKXUzA
lxHrfAaJ1nMayA4VxYxnrEFOhzjEW/IWJRw5NTW1LlnOI6yCDvLbMqeTMB+YnbzT1ajevadrRKiX
eSZYdTy1850i5z8zoOUbmza5Zbha59W7bnOVQT5EmoPdhLLL8suexlxzbFK9IYJclzUOe2WHQNGE
SFaz61f3SYjc0vD/pWVkP9gETre/zmwWx5oWv+pYR8qa7j13fptlprqG2oU6VhNL3/pcT5x5qyNX
9XX+3F/gSkfzOYRvVFydnqsUsNNcB5YdII4kFudQM+FZE9vzE5BNBG6Fa/Ub4ayho154qG1BXKEq
/e4eB1gdq/byObVnOxm46HqWew84FNzIKZDBv2VXO6BjIw0C2/kLRapxJc4ajXPIl9xVBLO4PRZG
/YUG+QUu+ednXJdV64KVIVMpSZ9AYBQwkaNlE2PRgN7qJTgsyVhwlCLQACMtkXCEJ6gjO+JAOl5k
Z52LiVG39O5/oHO0JZdT/UM+RquyDjeJf2HEti1K8Jf+kRoeN/THHh5EYYOsv+i1fCAEGi3HbB67
8kNog/W6y8uGaf8iWUvQWKLCyppGr/JGgIc9EMmLcLf1JepTNHVYXLO1y+nWHn1xl3KwG3vdF7Ju
96A4YXLNBgsUqORUQLbJtK6dR0dFMtKamS7wVW4TPfImnBVGW1LHQAnS1af+7bqAVHBeLfjczhCW
sf9YhEWy5l9BJazKWPpJxGCQ2aX3qdZpYKZoBx0JrAAiwm/oDkJiKsFYFVBzoRk1whxmiJf7jNid
ffQqnTCAGc56duZ20frPVBagxX/VIRCf4Q2DreIGPpx8aOI0Q2wGrNpqzahyoOQ5brLulkX0Xz8M
nG2lBZBcww9HyK8SBw6wpXl+6XbLS17a5X9tv3GY/EvpQaJim+/ksCuouDZdb5YBpiQSC5YJooDN
BMFs4bIf+AgzQxJOcoUzHkWQUMTvt6Katb8E2ddE4b5fyHx7g9JHr+76tOnISw48YG/jK6e358e5
JEqbU14yD/bthJLIbV7O+OVwkH11qBRnAtRD3wcki/nb2Wupyy0cClpVOfo0DY9GPBLYK0z49HXJ
pK0e2O1gvFCmP33SieiJwWuQRP5ClhT+bLocccRrZCPOaL+2rN15nOnjyjxgUdgYv6CIFJwg1HXR
xSjNXmLSIDP103kKgxHetPV5bHTM4D1BHR+6XrpE19YfmsLjONXBAw5BD2oNUVxQtH6PpQTj368P
xIdPUJwQo4hup/gGTqvIw7LWBFvrSkFujmAWjylPAAZZWLTnokBWEUznV6//HRaCBaOpVdwepYQf
4dHqqyEIC5wBQ8KcDomoYDDZt2I1oXxU98bsjJvFOz5+iVtRWSTj1LbjA/QBw8ROo3R1Yx6ptrLV
CdLzw/F9XE6UgOfi+mAHIJKTPzxP2ykz1LkZhigSsCxcynUkfFzuY5mpRJDlVoyXMbSK1H/pEHMb
9F1HYhwEGNGwqYYR4OtDlU6DnbbO7yGU1aRddJMcg4yVGjIvKsgkekrsQzCCUSF6UJUDhdn1I2gM
z+nMWY0bhO2AlqSg2XHTWx6X02czr6AbaSoD7Ik1nDqmVVnh3D/sQ8R+D/hGXFmupxGuDUxfEBfv
L1q53dy9StD17HoTU3bp9NyIjX8YyatF6Pr9i03Q/For7I8KcAr3qg5W1CG42YlFaVkGN1/qZk+K
v30bjwTzEdJXpbypoLU0DKcwNaLdMLGpPdTwpYoDKyaQ5okW5zSz4WOZ6Qhle2OgemOkIlfbD16v
oCw+zJoHidXc0e6yNQtqM3utm+F9wd2gHfD9NgkYMou9SKOcuiXhs4V4YYDZZX6DCLSjkA3GABjP
6OlQgWGq5lZkEQaG1Xyb7iAy5k+3BKqiMhe0MYe2zeOPnxnjFZcA2ULM8wKBXixb/xXwSo0hlieS
t3EOgtZVkJXmwrojWeZ89Z5Prwjpn9R5HjD8WA9GqyCisEr+1ladidhvb4ZVZLPEuw3J0TjDagu7
QZ0w7lI140NDhns/emJJ/vr6JSdZphljbu9bvBAaL4TJkoPzTsmYbdKjLXSFXkQi9Mcb63AaEgri
9T1XDQhF4xrz1+SAZAX2BP7l9QJS641Ffd6UnJRUPVeX+DJq7zMma4/6NjmoIjHzk1MfHgWfuWC9
kp3QFZNSBDo+EMzX8OLoPV3NYfedaMOyNuS4dwmnf8SQLyhJf0Xf/QGqd7OYrYVQtB5wZSHgdw2H
J0fpXOLLYjyEVqauNiD7z0pYaCFs3Q1WkMnPXdoKgFQYOHrXZwzJ5L64MfEalXeOJL1TK0eT0pB3
L6U/oF7eAVqNN+ZR0tPkHlqc0dc4EpuXhsD/KgZNFN0FVCi1M7sNyFO9Vr7GhmFkTM0d7ID36wUp
PYC+f7WKnLd6Tqjbf45/ybp9g7QEHpIZ8kGrTSzK6so6TpBNaz1FZgpXphyZ9WZnQppbb+/l3QyU
6kZPGXX5Vf6dqFIFR2pW5GFw+ZdtwhhawF/SomG5E6+KpQaVpxMX8kG024BOWHTBfCE/1bFBVgLp
5GngupO0O+i3CRmfiHNXKXMZE5tpVIRrEWXg2ypcygaLhUzarajqaPXl9u/umz70RvCMEOw5rlOZ
MqK3v/wjddjQskpKaiSgDSgv9ggsg5MEPVd9lRW9dzUHLSZM1fRE2jEiTqAOUQFU3jAAaeBEo5F+
q2Fh/9nEbQk2VEmV84JO40DxnQBCCwkXA7fspxQwe9JbS1eiJwOyzXDOCpqVZs6FAGjM3JZi7AOi
w8dIgd0NHqUUQixlEiyNwmLIjZWGySDzBuhuCnV/cgI1EB1RxTkmEgWDfEJW1vVmOPTpL/EzoLXE
4vAQDDQIfvkT0pVt443I5ewO1Wz6oweyGjICtJVbctWtsW2KsecwSyGrVhDELpEsehC7tIXfQN6Y
zpLT1rENiH++ukDfoPXJfjMRHSplDVefExQDhKkCwSO73W5W66LuYzlW2MBeuIKdn/51pPY8z7wI
BZ68Hds+A2ZYyT1op0ErqPgFJcvxs8Nrp5kV86VNoQW9rPQV/z9DvaaZECwusoLZ8dPX2j6HlXAG
3vv1tvNPz3zj3JYi1w9Ahx1Up2Ru3eBUNkfNTeSs6eV6L0/iW1mJvdk/56FgVtOtR4c6j0QuQIsn
+/H4dk7MllmQ3s53iy1tIoFbNSst028jI7qIM8tWLVUranHQGitTHr46PfVSIyDWZeKpQtfAyP3k
dLZ57O3YXdrFVSGMIzwhL9pgOFo06xYFBn9f+EKF6/yA3yKTYuEODQxG8rq1j5xpNEQJdQPr+4LY
0BXrkhbN2g5GtZVKRKvJrtVeb4JzcArH5eQq066QuY8wvSA5OICboCcha/hAFIUbCu2Eg7tbdiOz
FYmVi94Uwb6yzMBvyu6WsUmZkle7n/qSVcQGwJl1IflA2HICS2E0NSSY577Bwy8rYjELZ32BrBn5
+zPN8nMCmj2VVXedJjH3qsmAzbZTMZzcFDI4LJ3rVrV+IXn/aZ5Z1K6DdScfQyNBH7hXJJzmTb9Y
KH4/DdgJ6jx9eTcfGW5AQ/0e0HBK6xc1YFT00PIbYtuAhuzz8CyVBIWifUfIu9JMH9xUwlTUQf9B
nOx0aFBD4wmb6+v5wv5TrB54t7W6gJdhhZgMbskEK54SRUFmKN9QkNv1KQAEgCZq4PbPZipw55vD
1ewG/9XeEEvFcAg3sTwICpMI8TxjaoEZI7jUVcSVsFvjQqxvX1qVxBC6FLLN7d7N7qFG3Irm5+H9
Dzv+wqNNVkbhz/lkxkmg0tWrTayOoGQHg9aVByHZcJQlRwYzLpVQAh8Ncqt4SXZ4f7GUmc73L+WS
oD6gckOmE7/VHqMU4s3GNjOt+uB/q0ocLJSgQ4D/jqniHqR7nHHGInqXd6dJJA45qtELjHro4pzM
6Fhy+/b7bL7QC4BmXfaRKdXdGKjTsC4pDLGw2TODyVFlO80gap3mRKnnEoN1RpaxTOf73Z7DwkLc
2hrN3UMYR1cmWjxtIzZQSwRVnE273UfL7CygMAo9D1vTplSETwh18QnEV18g2zU3Go7vwKDDc2WJ
NHEv2fEkxLA1XmNmGuwTDhVFCHdXaoLJP2TbOGh/HWEZdVSkBdb4azJ6RTh+gX3qKdCabRW9wjOG
7QflErA0t1RGzPNRk8mG0h+luYx4Gia0Qrq5RL/E4yRw4Cv8/fSkuPU3K6rCZUAu5W8B2owcPR6d
1WLAHov9Phvl/m9pLqT8E3/qjG3aT+g/X5i8JkfcS8Z6yQYr4HIZny1IFXmB52AY6+yzwKaRevmb
ZhdySfeMWly9wX9JCvY38i4Ft7rJbz0Gu+DgHd5+JTl8LGN3f+j0Pwm0WeRx8KJ/xbMwRfLpSBdy
xMi/Uk9AJaXRVZl62abJpST/PsgrPNBWF6ZZPsm6iKC0QgnO/zo70uVRtOUHSOCJjAQjYKseYrhS
VRvv9y2rtC0jyCNHgU90Ge1K44WUP2oKFU/OXYLgGiVDCcnAyn2kmmykxdRvJ8SgtwEflN044wC0
H+1vcZTd2bXhdSkUU/dVCFlpu1GKQWhrDLoeahcLouTl753ZYnZpiT1BTPaIdvsuXihtvla1g28H
ajFzzP4/SbRirKkEg24YPrYuk+JZ6HXvNV7a69lymvfbuEgG151SInMqwu85+EDRITwW0+YmQcs/
EQSfxZ6m+VNkaGnB679VrqljnkU5elYELYptnKWRSenLKXs4+0HIucCw79kQ1Iou/DdXTOxfH38N
NRiP/pomKZSXVORDp2mJGjaL87YrYH2/OfWy6vAb951EEuphVKA3Vaz4VSSl6ZtNSbQ2i4e0Sa4D
qeQgExnnKR+wTlY1sphZfJ0PZG91ClQvxIVZdVjzEB+Lh1VRBLv/mUylinjjvZ/uJczCh0hW+2FG
hv5JnhbxOkJXCo8fgAzKDg8lT6wh1JBroo4kfEtdFglOpmbWiHsrY6raqRRaU9zKb/YSLfMDCeZI
eAlAsx53T+X3Lu1/IM2DNMhN5gixu6FPFIpYj4PZZhdeyz5xikCPQXhyrX/BQm9SXWpt39r75wy/
j1qpx4gAJv470U9Po+aN9uZQcsDrebyoPIEWJdTYKNbDjd0ksWYB28j2nFVUOBV9yqvMZy7S+fRB
ydVMmk/5jR6//BJ8d/jpuQW5MDy4zvO+dvvHFoFMr+KYwnRbyfMqZkjFDnyzpYLa3RvIvbQAGqPC
k11PoWtGakpvCTHIhsP5yEGjoB2XE9WKWt/cShHoZCy2gKnpH19Gp7UFHSK/2LSOJw8vIB99mt07
o724lUbu18k32gcxAmTMpJdgF2AHD19qoTJazDk0QCQiqtAGgOJHp8TQrBfuL+WwJliwpdyu6YsO
EFVBg1OS3Qz3cMIbLe5JfKDZjQbeWMPEoEZ2RddzRtOz3OJ6DVPFBz2t1JK4vklPsoepoP7r5fsD
ldBmTbNKyfQXaMaMTAYvkw/Rk7RVrRJyMeXNb8IKmtVasry2sDoebirbuYDlISIop32MozY2O26T
Sl7BRCZbINqKDog5qCCMkdRCvRUJezeBCaKeUFNLvnEW0YqAyQvGet+AowgOs3cVOLjqgmQxRUnm
23mDf4wMqJRYXVbGfP1sCrb3Z+OpvfMjtuIURYIqPilbdYu8hS3PCcl9zqoSfejVDq8GzDKqxgMB
pzyMgBzrfGbDYopTEZRfxJsBU0EbwrUKeWjsb1hnuu226NLe3qMfvDznf9iqukUaHgzTfsOtEXZ8
UfId6fsh5hgHPK2+4JLo8dKN+XR+XK4Lhh/IenfRWP3VqVjbRJYMeQSAAE5nZNmpy9IkKu6Htb1e
hnq4Jx/R3FpU19ZyRw/dxPWnQQuOBLm5MdFloWUouMD5BHdiHCF/T6c+Ve+tf7jJUMq/bhmLjprW
l8qePQ4pvRWEaGkjshlhsnTgezBsqphSgIlmoBZZt79HRwnwJyUaUW4jXC2i/vvnrT30TkGd5jkC
kXOsiJ88Cafver7Ptxb9mrEShodlHmP6mbji2lgVNURMaiseDIg12QfHBhaQcteGfdi+wy/QWtl1
I9zM/iDh1dYKk9m+QrDEX2UKVF6WOwPzrmrmmuafVAuanVhQwO2yF/JefuYQmqVGqSIVIBqmKzkp
9cUQlQfq/U0dgYBe/ovIgfbqkbKkJNddC2JRt+UGoiNxFQ4QqxYeQ0+FD9yDaqduFHBd+3rEr54y
RXqnl402O/GphGF1lmcX5SyTjvxa5XbBNmD9LENO6e+LTMD6V40NxelQ8AbZNQwMOKD2wkP3jMRp
5unWDiSFZj4d9lF55aPTiUeS4lpEC3WniJv4Xe8kMfP/w7ovZipWDzda2ntZOGhNEe74SZ2CzsbQ
y2uT28WnCU9WqRLkXHq8oyi5FAzsT3NLoYG+n7vaV96X5oXwfbvmQjqYxvJB4iAL/euP1QdP8f/I
6d2X6ofNTuDLP4QMpiwGtYhCzeL57NFQaIEtTFwVKQ+tpDOFoi0cEgtmVHy4KDHaDurXn9wvdrpR
/zdLcXe/wpaeGMRlIHpUIIFZCU9GeD/qMJi7xRbF+EBeVCmizK+XMxMVkVBBcp2RF9pq8UqyN4d2
y3zmK0JxQKHmLHXJnczQF+HcFYRvF96vkpvFnosZZw6olLTEp6wA3qlgwmsgAfUdVsUCcJKdsCxU
9vFMA9tdzz69HQDJk5bL1pKiJVR/EpqQfn3qKAKYDk7K3tmr3sMl679ZNQ2eEbooKarsdd7rp6xF
xChhu/h7q4of+En12byqGQKH0VGSKE8sksA0YhrXf8hSpgN3vm7VZx1kMLDYkptsfs3XmJop808+
QDCwhXVVws+EdeRy0dZT0yxBmZnC0wwxZn/VGjKumnVOKP3kFgYLCNZPHP4Ro5jZ+txHVhOVtxLq
J3oLNcwhp/naoFnSdNo7ZtU3BgoXLkGo+AtGzofSgVMjpOaQdyZ/U8dweq7nHqP6Rf0eMsMbzbnl
qbvbS+VdB8vTxlArJthAIOo/s6/INP30cLaaskWuTPaQl+3MVIwpWeHRTYxBpFL5fGDKYZdJuBDy
sd2n0lYarNryTuO4OVY6KFlewsY9u/Po2NEQmrS+jPfTOB5qf3+SkPXwEUG3DEJwEmSzkIfygnGc
x36w0mRxI3yQADfCDQu8jorpqH39CXPnxZ1QDQeb79fWbJ815DHtyrHLyXK32DAY9ZVNj0q7GHZP
buPG33E5NfA8h0P17Ovq10U0kSwpRpmkKeObrMYryOrrLzjF6t9CmX81a96+F9+LJw/kaCzLhKGo
PNHRm3MYn4KnuZz0f1NN9Rxp7X6WTHokq4Y25kgxncDsjUNGqW7Xos8vXW3owI2E22lxZY04COS1
GWSCmL5I42crL1x0n6UmKprfETDWmcKklrOytZNVr9ll2tNF9kIZlvGNvcXWfCt6sV1D4HrZf9Ns
HMXuK6ACdhLDF5rST2kIho3qnmq50fCNA+vtpA5r24fSu0ktiZbP/RAs4e+5mdau2ZpNalKckETi
a7Ge3UG6VDJWSsSZp7Crx8P5QNO0Nl+w0H9g83abuqAgNmEkV2/cs+CyAG2YQqeWLL2mUgebfm0P
kcTE7kczaHkGE5qkofdGPPB1Kzzo8ehpB5ooVxxabSiA3MYdq9BNDsxAw2yz+Oip6lrER6fZnGPv
qjRrkcF9Z1LjDgrku6Bwnn6IJfKtuttmPRLiZibyKpfCf/ZwP37jCGJZgSN5BHk3l5HWSXVXxsNw
hmW3U7ETWmbyAfoXAI2mGyyZLSum7s4/5HiVywzY4kuXXDD6g6I1B0Ae74WBTyRzrzTs86i4yyvm
LhBrZbIV3li4pGvwg9Uilv43izn9hyRIEQJ9SVVJX1X5zsOP7XKbo5kSBC7ZuDCxqhxZJDuqtyQ7
dT7dd05hzch5sLYT/zp78g2C84n637ub9SeESSv7YaDpB6La98Q4xy/zkgqG1XRPUI7kHxNTUvbc
0oaZixOnfpfQOZtfA64gdrM6GAIrr7Ddpdoc114QD+PWaXkWI5o3LAcbIYSpGtUskrIImv98hcct
X0b94aAFJgCnBUmmoO9Xg+h3LayfUAiCeECzb5XmuA/L34uZjqmCXxq0Eg8We/O9aFhiib7mOkeQ
wt7hj19nCVeIavoqElYbgoHpDsiz4ZfguHJT4OFBmRpgAwE9OLFU8t4UIHXx/dxUOgJR4HMPHAc8
kmyqXJ6dyVHt7isGx8dO9Aw77YO0CTnTnfWHq1TzuBp5mf1ibb2ZesUfdyNL/FBARH45wXhyY/3r
LyJFvSN57sammc11blAsC/BT0TosOVHY13RYfX5R7wghQWttKIzoFps1ZxlUl7OGsjFc2cIgSIND
/Nn+8jACuo/6ghv00ARoM6Na4mvXXldQoTQpCypkmSB1041d1x78JzgqfOg4/DxNrMIEcmGdB6YF
GOEm9EmmVyPz+S1ZyBM4Zz8fLaaROuSSgb2F0wo150EkL5GQKt3zITmPRY37rUiB7vM2Hip3Gmg2
iTEKWajJj6dWJjZaXPnbgBHp3wu3ehMGYNoJcuwfghqq6i3o+8F4/4/Zw9yB6G0YWCfmuAqoPdIi
sFwE8jj0hg69VdaROnhVH8HzWR0C4CY1BJqE9CfOaj7uG3MBVNtO2qVPRIYBF3N2tp73tWo+jqnd
1cVVpdS0L8kEqkdyAtLQGQ/8Nk0lW8sNKedfeztcB4eNAvqHkzRrf7n4agKGBACKUl8wPGocTZGQ
z9Oob95Dyg/NoNQN2jx7t5Aul1L8at1p0F7AUq3E+woDu2dELdwykLwdCQa4kqtv+L/3vpMT4xA1
bI48oyh6a3idFU81zmrEbdtYwGa/7iRjpcR4NQbHddxohzd7I4r8PJREnQghWoIGrx/5TTJkm1kz
ngHyMFpC6HZwXyBV0BLzH8KEUlX4ph0ADo7xSAifLJkZCLNXz13GArd9/BGRggdVeeYwYidXZmyG
3YM4i5RCBvTEG7geHBGLlaUhZZDd40U1HF2h2gtH2sC18gPApir8Lauh0SUbQxrWJAJNl0fnXZ8l
d1X+oC8tMSm2pZrDSfbRy5y16MBN0PO8zSimEXGG/eYIBfxMIadDWkF3IRDhSMnfqSjxgcNjYDhh
BsrSTs2RyvRPMB5ac4Qm9TyM2CewzLkE885PcTxJx0eO+b1mQoZOvxY61yNXG6CP7dm8cWFdA5z5
5ROB1GODsCbrey8CVBZ4CdqRIWS+578as/IoKC8WyWAhAh4BBp1/EWegXJdJydETr+nQrWGL9DJs
GuPkIcR1v4LQ9c8RkIya4Duh5objSthw/ulQ94DCYaxTkTPUmOesUypejsr60oKaRKhf33ZDlBxK
q+v3hChwWJPnXrhB7l6Bj4qr1Kp8UoaEvAV3/VNs57pYPm5sD7/FX76fzGcT/DRI4QYR9SfK4tHq
aH807bTcp/VaW/skyWRE/elq1rAo6SFPtWcZSEpvf/ZGmkaDUTRjJQmSjzZjzNruyIenbF20WYca
Oswl9xB0nhqZegABAc/UTUtFZg7AwJlhfi5aWRwGiJTNWrJlv+DLdTF+aj5heQ5cgIMajl4uM4kE
MrzcAxf+p2bEitbv6Ryw4tPJjPWZY/ssvUz5pa9KiW87pikC7ryhI19lSFBnPab9oWIqSLhQlTu6
dSd1WpOwZJbzo7vfpzLYrkRJagvGSEquS9hrUuA/rHGhXT61h4N8J/PS+jCpZI1yG5Ccmgh888hn
IXyZuWoKNiF361mCi8sV3YKpXzbwEe7rzL4O8k7+2zJpwDIxp/6Mlj1JMoOuEs6e9lpaPjtygaH2
kzZn+XEAamtSwLWObWJaGNoVDf7qOoicpU1rTdEdVGPx/iZnarwnROhGl/Yy2VCynX5zFck4A9PO
R0XmLQGfE0wUNA4LM7DELnhCIZGJrry+j6LKuZuELC00GTazKJSPDI65Y+RN1n7dvwe6NzlR0UPd
g8PMJOxBaN+GThX/EBQZ8xhQQH43AC/7vRWLN2fUz+mV6cL5l2g460sxneNsS7CcID1N12JDt8DG
XxI93Z0fXIOPqJ5m1mrHj87Db3Aidw+tu/kc4y70CN31FKPyprBWPv46l8BfDIdNdnbeELV5olTC
4Aq4n72nLcfPRx1yr1KhBcT7EsNtyKxrg4F524PSU/yKK6tGnIQ/aA6Il2ft4z0Bu567BdS6suyx
vy7iWAjuO8fqP0dPjhucqTFQy8EwKrCKjhJPciPQCzBv7wEaL7XBJt3rMu6yDCR6QQhBjxs4Vb7F
dEqETJO49b0Gdl57cnbUTxi0Wl1rhFd8GBgb9ydiu8u4TKYl9HnAlsOq8xk1jEbNi8UxAZ6LnXoV
n6QDHaztcZeWyxRmk3/3z9A+AJ77u8zXl5Zcgu8fqz9jWrUw5f00OTf6CFHzdMpXEFvQi8l2UEj2
CzHT+doIUZhytec1Rz/IjHekNfaG3W0K1liJBI/eavoNzvQTtuJbixRpXNlxu3wQ4fXuA2NojFuG
bG4LSQCQA3A4cD4+3GwbAFoze3VZ/w1FHSZ7xRkFoqoVVODfxXA0+opSc9tQ2iXBB85C19yWTiRe
wfV80m6c+BuPOflnpLQXhoUaqwiRtN0MmVhV8ZhUjoVma4hs8e2zf3hePQ1fhl7TaB108M79+i46
owFMp46LrrVTxwJkGU8rGArN/OAXRIkpnzyoUO/jlNnhSchTtDbfgsxGpJcXghbiXc8BdqEcnREq
22FQTPyFSuHInk2VsklCBlNqhTDdsBe98h814PoH+1LNd/AYf2DvaGms2kG3su/1Ev+MkimzFhIx
PRX7Q+MNaBjjwJ1cmMKgrS3+6j8QGOHaxxsWliKVbDuV4B8uIEBw+SNvAYU9uXiE+XeWdPWOnC/w
EGKovYSCNtda9dBWuXLksw04up1APhtIEkGiyaCJagTf0dyP8qFS+qQZ5VGgdIipfBqundcDbHFR
K8rpPV+76ZOioCkBLzEvaxV9wt43iu2hxv4Ql1qnsEi0CtD5PjGD0oYOy37Qt7LntYtshPAji19r
sNPQkXDTfMzgnWRQjoC3aYfUh4mavSFZbNmmgZO2sDQBQTtX8Hn4jr+wpAOfBjC3dKM5Oafc5JxH
PbkKHBpOWMwcVnSwdvyyKJ+MTmf+3KbHNEhXb++F++2CAYkxVTSp8XsmOZfE+BCca6mdw5xqyOv6
LjdNCbZ4TPGch5r0UC0oEqUVGj3JVx+Rnk0mpIoLNSCQRjm09lMCrQ3WFpZkHk+znaIxDdKckbSG
8eEbeK3mO8q7Qd5OGmxwb/sTFSGh8IWpP37/KvyRzVYhBi9KGcFPjy7LR8JQeM9J3cpyVoL+IXBg
zieWVOkA9y3tHzxHR8x9zN7+NitNcGvyvRAJYASPec1BCsPeogDLOqdhCbDIfw8GwfbRYTKkQZgl
Xpo4vjuC4vWrmOC1r06cL+FQcvlGf9JN4mAfz0tjJ4hu0d8CHsT+uVSRgmILrndKJYvFwqjXTU/B
hI7E6H+RWFfElqjSpCCMmfoont2BQoYYTv5fCXZTzI/6R4JvEenYmxO0TXviQAPI3vD0abRhGZum
MTCxzpg18EJzHtrI0kserXrRSoPoijXlkY/fdXQQ3svKE18a3w3VJl2egcGoPLawreBCWO1laRX5
TCqMgML6psrqncq172UARW4Fst6ho7b6Gbd0Do+08rJgh2X4FXnkjbL/l18ADTZo6nIXk9Zn6OcM
wJUTYv0sz8JkjAIXMn9/jV28MkPU2CRBEhTQAxhjQce+gEESychRHRRDVc/beAYISKUxSztGt3ws
GoSubctxLkzoRY5WCjaFhl+A83jZzzjbAHHyNIhMpUyDVVtsZ+dkxnFTLXOc7zlPVKNw6K6wNpF8
+Dg6OdzIR/iiJB1gj8dZBP/8b6HC1czZ1kePIu3PdXLYql6EBhGbkTlvf6MbLJ0WSzK45tFGq/GV
QnOoKkeL712o0C08XSpDHBJLzie5W8LMUk+e8+RhE/PQABBmaITbuIo92iUd5IAB38NMfhGj6z6/
dsAxQ0D2SbCf4g1DsjYxzPgwK7h/NZi7sPJPpRvlH6X+LCskOVzQElwhnr5qlx5ILo2jEbIGqg/H
FKgRYh5OlpV5mqCL1H1BmIa2E9BWA+O+oKH3r0tTACutE46QWvSyWGWwjnq/nKnKqFqg5aGW8mHz
65L98KKSXW5Lr6kWct38oDHsMquKxU4lnuSDcshp9dXmAF8MlX60nP1p/8rJYFMZR3QJlD+Qfe+L
dTipExMYey4klC3xb2KSk9p2lHBDlYlSm65N8wa7i5ywLKeohmuOUZNXEkt1+BwSb+bM4n9OOrNX
5hXkEpHESzK9OpP4JlNcLNGWu2bZK3ogARaKMFR3GUdOeHoYkko+yAYUOIqKUjyaQ5bwOc8VBXKp
Ufb49F/JRttaSj9CfcGVuAMfeGydh2Ppc3yVSp5ObrvJfjf8DFk5bFhjQzHSoI9LdjQRTKmopj4N
exoPixaf/zNujj+rkKt8P/nvQQ4lt70jVmMKhy/fIHzc50dtzKpomOOdQSHIPRGtF2MjavZiHk+b
2z+ZCQQjb8vn4+CZToXw0f3LRKbRyz3PX1FVlbgwGfYibk937S7MJxV/AZVuVlxpNxSPBmVyCqLT
Frf4eGol3lnM0WoluuJJKdhfIP/8G4ygqolnpyAztjGfbHNfrChT2tc7PmDrxnfGc7XUljZus+As
0oyhHt4UTpXQIej5KICiP9DGsO6N4im32Kofy/bpUFL1LsvPCgB1Ap1dVdptpgah6fc53r1cX5i1
Lk8gK0EQbR+Ffy8pZy5nD2Ki497h0H53E0rCI9gDTIkuXc+lVR/14M5ILTdO+PMhTy8W+KIm11b/
D5Wj5eseDQlujjqk/5oQ1SQtmL9y976WBOviW9ylQFNrDxe12LntoIJfM+/8VqprHINLHCa22xmN
9I4jSEnQ5CzKJvbT4QmJlbY4sL4w93dfypJYg2fhgmtlWForAhnlo86ZEWWZPJv+K3PPJjYfyeDQ
9yUEICIlMM5LVKdE/v7iqunWD3K5LfLQZL1OvTP8Hh013mSZN2Hp0Y0/BhT7BR0rNKUqphwHbRYs
Hk6Yx+ZmNqEANVeCVI2ovyYbm7TtT1cROQ43CWCjmtUvWjT1Ran376/ReS71uK76atatuLpp//Y8
IzGVZwhzVFFru8GJzGoxnKyiWyvTwku8DyC/DxAbtPFo7pScDmqSOmOljIf6+dOpFExjX7WY87wm
HFrYHdmZLbBh53OfB7XTCzLa8kfLz1xkVqHydYQZrY1MpuLDGGfX7VKNjM94itTSD+LfZRVOqd2f
qia12em5AiGwrBjqerzZCQZinCF5FV55ps1mAGFFDkC2iJXSlL9Trv40HzUQubceUX+ohVfWooSs
a62TkgAB1jZVZ4nwK7YjUfUwsjif3EdDI00oZWw0DoZMEgL8EBdnQKIWte7QO/xvDdTU39VzYpic
B6DCKiXEy3Bj2qZ++UoGN5ft+08cr7rZayqizGKaAl8kaw3hTEReXo22onbeQjvGjmluZihs1bds
j47RTUCB9zSN+2xDNG7BW5XL6F82RSTsKITvj6ZIMG677qzXqw69UOlDNiZ7VZ3w5uu8IXDi0vAG
L7/l+miazfNWumJ7ucwarL2BN+SmGwJ04uRMUEiVTAiSFz8As9Zfeuq5GzyfH/3DZWGI3jhK6Tbq
qsZ4CIb0SS81w6RQPTtE5h75GKo7/0zyuvXn13XcPT8AWDoIzNOHun1HdhLlAVy4gEfyzgiefTTi
1CVgLbV4EkQ+pAoVsUraM+S8mwg78mnVBmktt/X3/XpRoxT0JxJHkgzSSAzreaOxvAjjrJCeVy13
W0meD0xd132BNbZgkjjn4rhRrnNJ/oXE9rr2ccDmqy+eCyo3F/5/duSTghDrcS1e327PP4adsCM2
2jJumGUbMJC/NSWEq4OsJ/kH4aQ5sZMXcisIoO19dGVPVYto5p10RJWJqx++aFiTKvepsoTfxWGo
cuBTqxt3I88Wuzy8MqZcGwd6kUbHYD1rT/XZgavVF9ljq8OZxgmwi+WYsxg2p+NRUsLNvaEh2EBH
ohH7mLIisDV1TD6Abi6+cD0q/+Ia9hydRtL6+NIQJnQV8JLkVB7DEULDM562p5gJivjVc5hiAp9q
dyP/DZ068mZsP6dVM4ir6dZaPwsgwdgzKIiiSG9ZLwGRB8l9xD6AedzTRdV7XI5mrgMCAagC42VI
sLdaGzs/SQtglQmIU6GvHtRDBFg+UV6lKpxfdUxlGIWGU5zWfEpn+JznEyK4r2GWRC/+fuOdZcRQ
U+eRCZO3BVXudI6rT7FL5tV1Ync+IdrONWd8WOjVsGqXkXm2zKtLKqEzjh15wDceKigpW/WFpIst
bch/9KSEu9gB1CTvrs3U7QE1baVib1UtMejRuIs75/72FCnn8IKEKB1NevrgmeloTR0VL+EbwxPb
ICi/oDlmlWtSZnB/sGYIBZnCcMD+RZ7iwN/2KXl+d5QE/F7ClPCscS56Ak0Vc6DaDK/D+vG+Juvn
ze0/AWPrKRAWo0ZfecdzZbf6I/hy+0IFLGHqzAzNeTTNyo8wFSU57+IqOUdGRxtfNygprFPSV+x/
/yMFPVVZmUCOFB981ha+iF6iS7zlVjI55FP8cQH1205436FkZ6PRaXnTzdyEcV0GU0B3e2KiZCDd
C8/K9B9bRe7IbcetGEU+iPoEdrC98eo+R7BQDsGCRRrnt8YLR3H0Z4RUBsAc3eAbhYqgxYciHoTd
WoQcUaV1K1aOsjoAQBIfU5dq+Ppyj3AQiHHT5sN9DGA+b/cw894o6E49y4MtLSxhRJEjsltLK9CE
nz0qfwM/f1PYmli05CZ3QWcyFkywevjrjwGjwswO+TFfG1AXUopylLH3mAdgf73C69/I1f7vcjmN
hldobVJTXUuwCMGy4ttQq4tfugf9TRlvNnq4H0SCpvacOz+kWZNhZNQyOaX9rocJolS2S/CwWtZ2
hNbU5/9lHOQuXwsD2zRf/LezdMSyT3l+TyyhyCVFsrA56HgaBruStzhVz7/1v7BMH5X+YxKxfxlx
4NAZPW/QLD2ehgwxONSlGWtQ3U9rL8iraieAWNWC+jO0wJw0Uu6628eBF1cbtK4HGpWvyUw8SkvJ
51WMPiIuhdMFgwYhUP5Sn+4c+B0Fd+XxIfJSx9tcqEQiNg7MOapa//VavVftRo/vUEcAOkrDgAKw
ACB4Gb4/TqNUCvFdvoSr8MH8dnFjRE/jpdKvpyAa9cCrLJwo7VytoOI2PNulQj5lJ8wM5vZhD1Mf
B7LooFxiZOJ7kmCWYS7YofOs1UXZT+zE1ywhmDe8CuDoSFeEDEyK9AIC4hG+mkSmMg0SPKWvGX3t
mrQIGcVTpkUNSmYFL6LO3iLxjMcOwHSSM0eMcB+HEFn05y+ubysHvYtM2WfEauknH/16zZoZ4NF4
K75Dth184aialX8der08aHda4FRI/z3EmxgpqNX8pbZ4hvdWJpxZShIcpi8iBzKxjNvyaiAlYq66
kgyCyY1sf0qPGkSGN5eX9YCfHwiDseSV0OYhtQlnXHu1aoGsWeMFJSnstrvlbZKexRq/ypKUwqjV
0MNaK53vzfRuUHmdLdLi7yOHoBqLy0UfudUXoWcVMRmgegWE6ETESWmzoeU5pq7e8nuKMbPhRQgr
TEd/9x6UpgnxivdVJLfHaUYq1X8UPEF6KReeNQyGgJku4llatgb/xLgULngML/mf6rucp/FpIZLM
2Y6p2wF1HytBAgJ3vE4noW3yRxWsWQkyNtMIBY4r/TTOghGOrgfnG/aWGsSVxeu70r3FjmLZZ39x
4Ymzd01zvtBL5EbBrffpzgO3D3+pWr2ei8pdbTX7NgHzzxQRgPIFne8zWgwCrUJd3NGIXZA12jI2
V9fLQy/pepWaQSjA8IP/9T1/gLTbxRlpt3bcKM5/aUUoY5W5r0GsSn0PyommhoLu8VvR+U46cwE7
wx1OQKlSxa3gpReP4nxt6U5ADXz2tyONFvJm1ApywdGiJmZYUgBhh/Y/iqZwjNLUPZXF34aK1RTW
p6dSY+XMMnMsiuv680/JN0HNeSbt6E5StNzPGUc9HpFWL0MPjfMS/uEDmBaqS5YwaYvDDPuM1OKQ
GQ8tAsLllcD9awYWKKUFQXEojqqhwyYU3YwfJRa7K+hu8qIm/SuqHd9vDz5nShsahKSrkTbkQ/o=
`pragma protect end_protected
